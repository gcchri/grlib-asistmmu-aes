`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hjZ9hwpeTYLF3ZYYjB6zFaHm6hTDnNxGKW6HJWsxGmGXXtLSdTYAXgm5800TBiDF
PakjxseqC8l8VT+te1i+E8Y2gGzXiPlvpdvWOlQNXXLG1FQ8+M5FtRvFZJ+VOUYX
Pzy/jZpM410H1Un0vfWOKUYzusQbqUaLoOeIvzXxsYD54C82Ha++aUka9zKxmLOe
VTIrag7Pq7+knyhB9KcNpeJr5wiQVvBpYYm66tkVYamps4Gp4YAty3sgO4w/zZeb
N5Ic4WY5WbexCnazjDer6J5pRwydLnaJQBdYGTfbm+WK/1Sphf37jPVl6l3S42mv
RisoZ1+b1vMHF+VFNV1zi4L0Etzhd8oyg14QyKMLYaw9C+57/+Mc9I2RCT6e97MY
RXIt5wX++rqSCUaIpaTOuPDPEcPJKLQHkROKGI0R4MQpQ+dZO5qzuRISzgbsXDgv
PuBxARlh9IvrwDr/XQ58prUN8asniwraoC8Lk4IfJC9Ho0eDRfA1mNNH6jhUmECs
XhwAcB5ibrdMfjzGd6fE0Ih8hhVKss6g2YCUOybkc4nAx+3a+ObnBgma4mTF/Xov
46Xv8bstOpa9jbEEHV1YBqcLPp2WLUzCp+7NeW1bcvcfXVmRl+7GAPpgFZoETNxP
HhZCOrAx2PGD70j8JbvSx+gZhGcvlmoQ1VaiJgHHMm40Qi0ADPuYfEn4Ij4kJ5+4
UlSYaLYUjtq7pquVNmA+TcNkHp6+vFtnDxhBrQ1Hu3Rxj9iF+Fqku3S05Y6of06v
EO3AMV33Jr5kqyj+Bixvzw7l/CN8qegq35Ys7elK0LoMUmNmLj31JhrKlgAWnE5B
kLYIdIjNo34kQ9NZbmc5WjkeZFxNIf4C9XybZ9xhBBXjbemFlvGr2r1z612LuLkK
ViBAmHEtZ4YdjxgvgitlbhLNXDICa+aeoLfNLP3twcdf8cL+E0PmpGSfZNdQitCv
rJ1zlEjSvwQtjao795D+bbQK9c9p2JuNoeFGx0altzd0fXuIs3Z8LxPYSfnaO0Kt
czEWb3yz8xrDtTRnxV2dibkWTzDCFU7+MUTNn85w1k7MJdbpQghm6F7hkSrzA1/x
GxshGGKO34kFoCohKTTHehBoAFY/CMWrR4AC3lW/0JWojWjDWw03INvFEO9oQcwp
7zIjDS8B52DLf2UbdDus8kfLVeLNLOPn7Pxl3XgPcdwyZu4Q20gbe6jo45hvf0cH
aWJvjv2BE6hFa48tKzSql5DTW43Jw+7trhiFSYnNmpvoic1b+qMnwsb61GAEjp8w
6BaB23zqk/qG8bbREacccqhMb3/hNxNqFfEY8B3JtpqX9DrjL6tk72+HVjT6Xn0d
cHP6JR5G5HQcjXyWJ5Adx6ePhFmW9NhCvh4sSukVfGAo2v/tRl87YrdhBmQ1DL9S
dBQzB+C+ClpE3YlDo7ZCYBZU61hbPPEQwWDKXXel9F7pZYccHJJqUaA09o9Yhhaa
EcTzKhgcwL+Z6W5N/Wb2vSl8skEv4qOFW0s/A3aV0kjgoIsPNlZYnM7cwvbHZrdm
g1m0mxg3W47l5OnBVKp2+1d4AJXKdjqD2y+hWkGvrZrD5mILf9VC5JR0nYtoIwu8
RWv8eL40P/DCyGdCodD5Bh4Sz6xZvkTv/vjp3Dns3mP++/Inj4tuQgc9cfUiH65u
znBg9lgMU2jgK92+2VxaXKJ9DxNSGoGymm68d0kGvU4Dx2Btzhm8oWXuN2LNwGiW
9jTCX/MSNYaWXkaXVXRw+FARtr/zgp8QTWmcrl9sS0myM1k3I1yfTDmZck5Ham77
4CFAijbiF3F5qciA6RnKgke0rQDoqTI6zzop0R5SVaImnOnR8386pIAk6Zua8GYE
wMraILGiZIS8EcjE8TX4CHP2W/2FlruwHqU2GUcn1z9aQHVtv8OUOwCPCfZF9aGJ
Pic7ef0vahkC5WFNg4DZwY+NpB8wr7/ljgBHVhXI4XJz3DyQyAvqbE0biUGctZmg
96cLfjrhForOIGu7TgrjkTnWhkJpLVSBeVEgWCvyhUXEuJ8YM090HEYSAF9YT4p7
21rGA+8CslPw2i2+KOKSIoUk4V3/zwa1937jmGre2q6wgjRbIkRCbks74bf31Mn0
J1oimpSHZtepZsYOvww7j5VOLTWTeFFSX68YKruyw62MjrUJ9rc+xLFv1PE2cuZK
D4VXQJupNZAtRmRIuwcdSGtMFhAKf/zoPCqAKKOwKDYeurnM8jqaOReclsUJ+vIg
3coIUh7POTBQt9GwMrUF2N+2svEsKbYixt01VGuJgd+rA1x/MLNYjSf7oqcQSydQ
klr3LYbmlDqBR1bw5f70o6iwu0S9lgushoDJ1HlXMD+c3zTZZwMCsJkYT+zyqTmW
0Sv9GrwV9T4goeNY+YiysPejEMCpi1842iRGipYpvIbNp2hgQBVFcjOSdzHhoOBH
CBwxydtyCYf8Yl4fvhJeBkvPdn7Uoxu1bRkREGaLx2PVARap3X4Li+V/0QYetTPX
vHZ5r65eBVt6KPcJk8dB/fvdTfkQiU/BvTbKfej9ZT2TN+pR/RZ6+Fan1KJx0Uh5
cg2JWGw85IPmJgevj7QXBRlSiv1HIE3FkeTlbMK/Ch9IiLsn6uY+LiIlQft5RVKm
TdzC2kJzjmE55eWmEJNV60niVIyFedGM/AvYEquKqbzjv4/kbYwxboI67+TrtewW
a1DpaEKC5RGpE8J7loqyVf8emouP1azkjGyMBesnpBlyOZY1Ov7Qd9VMQG/bEgMB
/jWEKo1AfdGQAKvJTImd0ZaIie3BK2TuqUXk2mzZUe638DEpULCqshRF0LZIhuqF
Fkzv2GU2J1OzrqF8UAu6xYiywrlM6/Gh2V17CGhbnWKr/UaIJr1IkTzksu/N4MCY
lr0hp1qzbGsB0w7euOl2O7EbDKQRFB17qjCVjUvW5bcxEp6Uh4LRMkfn95QEikGQ
MK9av03x5J5QiN3IsSYH8CZnHD1qoJ11y8efyYvaoaj+D3Z6YZCo7upTLW297eI+
Go/YYQEL4fI61gcfzvMJwR7t6on+5+2pe/RZCjED9ZD3SLtfGve/8G/NyIi3W4mg
7iqY0Pth67aaRYGhbWEf+D8F3adEblV45yzYePah26Lx/i7fH8xVsnibagYQ5UwD
Ddr3CouN+/5wSaCBvyUGyKa0OW5+WzH+vXaEHN7VvciPhQHnPiwEq3re6AKiEZlw
mWF0zGUeEwkxxdPjN5B88GqKMIrHHdnVqDN6foHyyO6ic17smEiNc5gXpxYhWRPU
afHrZJUTS3B+bGSNxI+9DVd0ZonQfzofj82y9KzVVyzQtwNBet3khzY1a/i+oE7T
Shr/6l2r5MlHcKVGKqq7ShAv9r7hM0FPpmoCCHFI/uGDtEzNHF/Y4KtUGitEW6qE
fPOipGWe6EUV5Jz9/4PsNewLlIQJSryL2axIQGQloE+nWTTYZ2dqeIjKFSVsK+Mx
K5n48YP1/8uuFTOHsWAqRaPFGKhoWU9l6DNbKpi/ALiSPJVKQTZkA0Q58p6t5FQB
qijIALy4JHSCfZWunpT2otJZmXrdVWodhf0cDimrRISPGtOADdZRsYe+pG/YkqYv
oNITO1TiZi74U1id08mU2LY8hsAXzKdfWRHspL4uIhGcz8PuQWdsqRggz7p0zCYY
0J4nkXKxFrrCX3AzWB0zkw3IVSPO1sKiKj8bVAgCER4bsCS6hc8dV8TY2wazLWAl
kzl5MsPnvANzV8VAbmg/nfrtvLU/K1kprivItj6xbjLxmBoAwGMKp6dZYYeW1WV9
O6VEuLLVBLfkZvW81JOJwYkI+QqBfxHgG2AUKosYCyP7Jbgxntno/+78ptn+TAox
AUaQlCwQUOIpVgPBw19J2nwkd9bSbcD/7FcgkqEr81cdWgQjrf9uDQX5IgoNDyT3
pu0TcGaXNrIir88/DV5/MKv/DtdizuxSbdRbFfiDsIN8jmXHeCCygAEmQDNkSYx7
l68S3+ZYaZuSZ8XkBJ0og5kJqTbOZNIdCZbN56D2GKues0L7oELgd1rEGLw4+GNL
4IXMWZ/1n4/9fpb/j4rZaE6UuJMDle/0pWI/uzXP9io70Oktb47sk6tphO+OH9Kf
+JLmm87hjFQzcbF74FL2Vy8LSmZ2K4joVfvvktY3aj6p01b/BGdGfjHszsoKIsd6
KDAmj8MTOhUFfZVXaAvv2mJr82pcvGnu8gOHNqEAwqIYS+/5BDWO9immRil64JsH
bIVfRxFYK+HZXyDpUALw3Yl6cI3Hapj/gxllR54CrNzpbgT64NV31N3iq33bZlxm
CYHmwdv0V5VpCx8HCWCRSrfUYTRW2kxUcxASafnQkkkY9r6lU24fCjcJBu0ugphn
tyq/I7N9QIAxQ9NFiMT7rktffneHgpYGhMo8jHVyjlms8DE0aL/f6t516kadNWi0
SiTzdIi9OxaaXLAW4MEDIv0tSVipZXV89CeEPrz+NWFbjP7grv/1RJRkXxu28gIs
mruLoj9toGzCtYxBEuba2m/LSxH1NT4JVoX6hOm7Bsi+aAvrEANACq/+Jn7uvlfx
7px1KTKPWOyj8/0B3NKXis7vsKuBSZL0/egVGyF2pBI4wuAvvE6NJ4X4ZJF2FxBZ
FUO50FozGsPIg4iKAAIhdfyDW5tk/lAaDb1rLuqXdNht7UaZfjJlY7WTiZdz74NC
YYO41SIviFXffUbWJatHGLgtRfDevqpS8z/tf6NVwXvQuiKmBcMA/Q70jUeWPH7b
umoEKIz7i/jTPHulEnDoZFMZeKSALDbdrfz+DW6dsFKx2C6ytuuKubwMXUVu/L7/
ZJHGoh9BFXwlpWiA/bJa14Rgry+kH3p8O7CurI46IiDACzFjsgV72sw3t8thAV2h
+HpDOf4Pp7reiaCZSbMX0WtdBAkD1XpBT/mtGWu2HO27DnrgYS1pjZiNDZi1H9vg
w2jxeMaV41nS4vIzWT/tCFr8aq0n68m52aIUShiIW8RogQVt2ywtDsmZ08lhZ28b
mmYpOBpBOrvJ/YzhlC6mw3WGh78vFV68DZcJcDw83wXDygLKV7Mp0+gN04Iaw1S7
L4YrQOodNOxd3GGSM/IFveiK6CkmsvtfwlVNR3wgGx7QjHenbHCQlIpogJcsmfTR
u5IyZhqaszAfo5JWduJJTdYWTuPCOq7GYToNYK1Ban/2vSKhX6DD03i0LpTxWVQP
TpJZVlAgjMTfolPOPdegD322cEM1nYEC57AyqzWa8xfjiLUuspb3H5j8189glg7q
Uf3fjjwpaj65MOqoxh4Gy9izysN4FvwYbhCNQRooAk0PEBJ9bQC1Lm0dlZ9BLWNi
20OxB+U6i2/SHM4lWZrJkSaJ6If3RIGpc33d/iuLzdBReqy5RqHYP3M0qpMHMZDJ
i9FvqwlmnptOOWUcFMXyNLS9cL3cf+Icslfomv4LwcekBjQnaoW1LsGgQaFriHT7
agvSIk8HufthKdMo8hwNa52Sj6YT11XzIGPMBT6KlxsAwDLckR5RQfJAeTZEMl+0
w7g97FjH3hC5CB4WkClpnhIMZhn8JVb9uRYgMPpVJUocRUe6hQfrzDSW4P3nxtZX
CscTHR/5VcNSOVAJIo9bcRN0wfLshg3KJbgm7wtJ8yOUzKZ3CDUi1DEqVXQNTcL6
MIDywBOa24vR758DUTJJF8PAK4eSP0dpyD01vjI5RFfij9k5ecW0Gt3xUjEKIxQt
qessEEOD4fhOaQBuwD68fR+P1scE++2ffC0lq7XoA6KX/CRHbiLMeak49PxpLXNK
4WHhTjM+HOC+GG/M33YcmSG06RPj9F23VyFFqlUERWolagoUsL8en8qjwb9V5jnB
OlZvumpRLGNBS8joP89nFrBSaU2LDnOcSm5EAohOv+ipb450XYrS3qpGw/a4EC7U
Qli5r7ffMnJ3fc0W9IjZpNtq63TeVAIP6gBJW8PN3bacJ53m6K+BkvdAtPYaKL+d
RMcvd2tsZs564iLx6PikFBOZbuiuiWsGNKUtrhT1NPMSaA21LoLTpSz5/mgh+JKN
2PL1oydoDv53LwVvvD22ERmwRir/njVEHTobwQ1raqvMUmzMnBvSXbVEKRlHTIxT
LfYnW7dv6m2MKLuSw0KCYOzc/Ln3p1MbSGDwYSS+4o3ZcxYs19DijKf9ybI1Vynb
S0GBEZuBoQqZf0JJqwl/1+lZU4tv2JYXbaQrlj0wjMMjUJ4W/IfkKXx20x3wyHu5
oXQd65Ein6CSrPBzKxonHBP8r8UmNUl/ThzdTNoKdJSfeXTVO89xlGtxN9r60jMa
zOcrES6DM6ZLO9x7m8TPxofeDOqD4lEG3zzFm38q4gsl33/qsqtLBcWF8bAayV17
SRV/p7WKF93GknxToJiswudS74EdjpUScW/XSDDEyuoclTK++3IpI3L5rreD8IYu
6a5RwwmAG9im+2GnoXcbr3NrdeLyEvap7KRemmSx2bTNll4tnpDE3KzmlkfAhPWx
mM8V/2XVR2PBJF5xCjAOsJm6kL/QZZPN4bqqplzJz4a/HwXpPnXEshQGlxc50xZR
WAZpDYDbr8AjdMEUGN7Sq743tAsl0mktU6kbRgvBmbvLTJfNqgLOAlAGIAA2dY0O
prVHrz6q/ZZQhsT/tkVWF2yRIkZtqmIk5fsyKX6KEQiks27Um7+gnM1fxHrp/p0/
3bmyjMZlUc13Wx5cW+nS5v/7eoshz/g3peYORzG9l8WdvVkWcPFUrHOLsLTqmNiX
0qIiEM/9lz/OnT7Tc6O9++strT5MLDbnS0TE2SAbKa2MsKazvd9pbDXCihkgh25o
PQ49Hd4InaaWp2lxKMi70vLOBColEhsipVO451E1MFOZ2joYfxA2ZF/f5EcYVrtL
kisTYNcavgmk276Gh+TqxQARLZkrEgSuQ9w8gR0CMojLHeyXZjXa5wPjZid0H1ro
elpf7TkFKZ+knwX6wNyI5mvTTtUeBV8tz/KYpGOeIElFcWQLZBjhqXpV6IT6vtT7
R9b7klX/JKwxtOLvxzpYWIfwI6BeXhQlfj02tUx7LSnPzwjolTQjQDZUsnheqHbs
tmy97eo5whsyBON31LQrLUkU9oYVRdrJ38xDDeZYk7MnVxfLxobulogVcVhXqa1D
lXac5v/yYLxAxU7rmJsukLYSBGPwdOb2IDzMzmFyGe5SqYis0W5hrKj/jfPHlZrn
qs8Fkk2DfBSmL0kMmTw5G+OOW5DCxho44KYwKp3HusODT2GKiT9d6jUY0xLblS5T
Suw19ZgkS9LtfWWmYByJ19J+6TMfA+4SJPE/Kz9tb0PMZjXXyFYUGg6Yz5R1NP9G
T/4U3PconObNcMQEe01PMoAMo6p/5AsblJUS4ainJL/0YeipSnxUF7QXWj38yVW9
aFMpcEJ4MzR8mz0xJqnJaZdJ9KjXD7s9TEf5oBrIhpdp8ijPsCz0PfxFZ+sdNcDY
VEMA/8eO1msmmXUGYY63QoK+sOPhfbosP+O+Z9OXP+a8Ixi49jLEpI08ESJg7fhd
Xra7Az6iPGPteH8XF+LRbcSqEcUIBB/HVNOgcjSpClgsr+CvgAdv724bRy1k4mLm
sIKxXtXcLFRQzZTitQ6PXObbM0BxFUEzhWgl6KQt/uTcgRvRDOkf1QnmnShQoT+j
+oQSJ0+PbzEp3M6pa8C4n4Kbd5w/sdIKPBVb+lTf9u/FQGOJDA7WAS7I8uCUN8om
ffQYmZpPbuFByiwzix2p1ram6SmhIpJlcOvMyuWjiDyI2ElT0G5BUzoWzqgZGnCv
HnLevx9dnVFfrVOzVV7quX4ggVDo15ISU4h/WeWHss3zRsf0InrEfddxGyv98lRX
fYFe+ZzJu3cKkbh5WcJNbW08qb/IEzhZBnfrdm7J3BFIXsabVsVASjLPAPOOsoRz
BahMHi7W5OwgjYx0Gq/Gj35gqxIGraa8KJGxxFUnRSRTR/aIMchaL7ta4EyhadGa
3gAzflZa2vMmEm/Zsh8TonAEUoRgkkf6j6tqcNR1LZVB+f6WWeswX7RfUg2FGXGB
2Yc2PnrRkpXlLRWKfk+tQ90UrS0z/rix5l5Nz9HA4h8pXkv5gGdi0+OLDDfRFkwF
wmu6eZmmufMGj56QlghkeITXuWLdtpbtq/1VOJiKCmpDk52n5I9EtL2SKMVKIuMB
2YgqUj5pLRVvatGHTVYKVB8OPoLAKSry6XLoy9prYegr3S1jhGWk/ISKW7dCIPSD
yLyn4cVJeKHOLNFag4REr3y08kJUy04KNFvBsrQLyoYrCHT+2Hrpldw3977YlBok
EPTiRisPon1ZAe08hglFg9aR7fIgkXcUi0GIl6B+0LBFecnXIS6N3dUvsHD3FFtn
78VyoT81XVyzOKOuM/63Gc23978fsRV+sSPUpY1VHYhR5+wkNva5g8GsWnxjKJTX
0heommsdj+IkKzH3R2p29s19jXiVVhZfNb/i2seN34KG48uNDGu31A4knRtrpP+F
plqrGnOi2ug2Js61lyzphhCODK6JQGLWrvns8X1hi7wEB1+pID2LvEMHZkTNv810
g+KpEyRZb/6CxEyuWE0YeJGSoH47u5P6D5OXTuOymii3Uw1mnXWKLD+hy0uNnc2H
QXvv6Kw53kykFywYv7nXBCEx2652142epni+/dQ5NaJlGAxRde126Nz/RUXcGfd0
yyHA63Ew6arUcyFsBOsv4g8JY0couq8MJmbOqY3CFc7CWpywU7JtD0JXobGpDF0+
1YtewiPJ8s85Dvce/Zuzk65suJqmfwADTfLTfsosuW/TtZu2SIAS3gucLYduUDFK
lA1DcbrqKr57ZVSbLRFfcr4Nt7JQDqUlbYXjuS5jOBiU30X0kMf7biAihIbIzV80
z62CriMbFJx2mwUfY/TccSwL0kvTwOFjGwmWCW7PUfeKFwKqtsFAGQ+1tJ/52yk4
JEn+g11pYxe5IE7hsrhi2cHi3B6lOFRrQi0z71qli/9a/D1+hZ+T0uDq11l0pgnh
GwpvhOTmHsAKgqOFX7JH2lvWcRNPjgsYRiIBG2pGwVNjPQLexTxeR6Xq9PqDwxTK
Ha+9TUBSWTyXddrVwsumRb5VhHyJwoEwtJNLuIUK2yt6tCN70VtNe+x4xK1P/y8y
Yp1yJF95PDTJSM+eWmlxEU0GY3pFbkkyA4CMtqzJlpwlRhLX9JUUHhOLm1aKK4iS
i5/Vcm2e1f/PgKKQzvHuRP3DZA7ex1Uryzz5CzOHUeQIGpIXlSWQ8CtfJTfsGtJd
8i9vnhL0sc+UI1ECj6xaij5Ep4RbqDoiKNxpP80QC0uajeBdyq+1zTN8ETXvnoWw
ANgnPLPVDQHSnHeeElviRDV5F+Lq5pzS6x7qiS3M59sY1Z5VNOglC8lZmJ9Q+QMg
QmlezqKhZWp8ZnS9k7QcxTpSEqRFNm5Nl2v2rrVX8ocPb3MaxQ5p/apbp9qNh07b
U7PZ1aTWjAbvq5RUEf9RFqiYW4YskuT4Oc7eW2FLecrfN8y9SmWORxSH7FP8bY3m
Mc4hUZaK9ZXSWdpwDeAmqg5ZO7CB3LelQjqBvqWwDUBTiqMrz/oDs4aeK0onq5c/
l8frKsNXX3CQaAhM0GHenS4a27aDgZxDzhm8W2+9R/ak4iWldrelcYpjbQfd8ZeS
3Kgcp8s+PuxYMRb2HEjgERooVteSklxPGiPxxAHtFL/3Sd3u1KEiZMKWTFJz4G2B
9vFbblTIhKngjY3gYF35qWM3SGd513MZvdC6b2Ac7kqR3oofbwVp54Gqc8iVzRQY
1GK8HIFtUtdKFaFGj89ujV55Lf9doSH/ZWVAKNfVqI+f4PW97NTYOLfCQOczex4y
CBL+Oj2ABgJhNJIDfdT1vCYpvRefJNdTKhcbiAo6E4eK1KAwBx1k+XvDYViV2ZD6
SpLMW7CV9VE1FFACnYbmVA0J8rfRStVI4T2xst5Bsxu44ZL96Sj5EY27puyUxjmY
3nL0tpTxlAcbgU6aHtToPpKPvR9UDnglQRRjarB8POqh935wB+axi6uUqbtADHr7
Qxun7ht071M1OJsDJmi4AiH9oGBnd5MQxzC/XR/tYKpF6zufFQTfDGE2uQxi9G3J
9M0Sa0GL2UWftDCF+vS7KWwngcrM8ELgmYlROxgcTgpPo6PNkmSOXrLoTToEnjFj
waxKEHXkTc4qwyBvZKwL8LtZzdcIczc2yTu8bQbJTfKBXCdLgvQN9LrsRWnt0cvL
sBtY77rIA/QPLG+07OyzePbd4K8U1k5gg4HrnbMCSuusCWCjqbnz/Zsvnpqw+3ox
gv4CXO5hpKSLCphn6uAL3vahnAGwoIVw3qDKdrdgT8GR6Hnroby4CgnRk8HkQDbz
D5m2qg5ZbYBfCB8Oju0Yozba5Ackhr3xjUQ1et6/UokT8e0Nh2wvDEEdOY5H3pzx
oNG6jxa8ySt+i0kNi11YzkM1LBVxp8dNdIrXgAtI8TynFi6nY9ENd7djLoU1mqIF
/t8BJqZlR5mURLw176BIa0GABwhngsJ0eqNhIaeBzFe87/vxsk79tmS0bKoGlTsD
9N2x4QUTLboTTGMGO2MyxRaGDBKFmvrK9fcBaHroaZuT4oN8ccAYzyVkd5Ezh2YW
dgxgBJEOXNNSufk/iKoC0Ob3c6Jp920Oplxfoz/ofQWpkLkhFYqhSBMBGSqOa+/r
uQMrBF1NYwt5bv7NcKuyAl7x4HDihNJRv7/JyjM+ahnouwquVDHEZBrXQRBvEKYH
WJ3E5e5YIMoHq5AKjV4ZFOCc78nSlPiyArdoVU9oHR+SC096ud2l0gAWYCk4egur
qkYcPjivhF8qI//A92Z8/AgXEA9fMh2ws/1+Ql6a1+lSqwgCpaHOpZIuaOn6tO8/
HoSXRp2NTz/uvW8OdBl+3ACCejEcqVzV6PKsaLxIURloy3pxSZCNqbON80ra3UJl
huHfBKPmdc7eM8K7WAa9h6MlHeD13UPtQYuZkWVP5ZOge9bzwbZFBBy889a/AKkD
+VD2VmckXwHI+y4IY02zBe3hV7vQeCMMyfxc/VSXfjKtuTI4a5N4YkTROnsBYgFu
m3EqT09BP/q+h3vdyKP8Rop/QHaKnLz2zx5NXasIUfuGhSiIWlPdQOBmJYUykPjE
WMWoMahJyOcI6rMfUgXoyyNVRJEThRhE8N5fUqkMHY8muraiUQ2KzjgWXsUu3jJs
+wRccrH660afT/NFIJtVtNZFn1C0RqkcS5WnCudZCRte2fiAl4GGHeeG2vkUDAVi
kazkl7UqZ0+tcgk7vui3Qj9NU34lbirjowzeiM+qNNu8qNi3LEn21e6TQPLsS6cZ
9qSU30wgEdckBXN+2lSkGdn5DOKssijIkxGQayjtvMj4lyv0ZWq6XvE1HaWnjYdN
OL1pQHv+FempijpB4I8NCUm5xCm4S97Qklnz3n4fk+OfjvS6DE0Wk1vUtHkCnGsK
5Uz3rXvG6w4TcYuhSiQ5EV11w/BmevM9rMe+Rfn4ZnwrzHUylix653DAvkgfmfdt
Zchoj8Gk+Y7L/BmM3VO5RM984vUDOSuw5Kjyj+LJezujRuD1Whm0lC5QGK4xMH8E
ClsnooWnt+D5RDQIM6oyO7AnFYmJ3RIbXXz3rptsBA1sC/7L6pC6iXs5pio2pnYr
ymXO2YpN65o/WGAFaX/vXUvIo8vGwHcl3lbLS1y5zDgMMTTFoXmmNthfHDTf2bsf
mqmGaflrrWCWnfNqqe/QaBII7SSmjbz8NVCoCz8rFVwcs7dlMdHWQm6Y1s+r43yV
J7z7d1zlssHqxaw+PaDDlGYLRpIFUOv4kMXD05r5yg8lTBN10CAQJHCqPIaxaWFI
DgCG8TLmw3+uiyn/gKmdNsopZgnbRpdFypHWhykOp53tZJ9F4KYtqMGcMmWO9dEW
xtaJiF7tBJTLJSH2kyny6bXEY+vA16qEimsuK4j/FYmaCftLweAnpsPvHDcofMxK
I+W+eqzjt+yMBsUpE5Jor8q6ksVq2jQMomZTR4FXUVa4XAiZh/VmpXjL4Xtx2kfM
8IomSzSDcz81siqyh0vh4MqpEGRFNVGq4VYbTLW1tFU5kk3hakD7O3c9+zFOlXOP
6IqMXGL2PH9fGntw9lIzmnDDmvhQ3o6OujvhFxjsSrYd/x/nfIFSS8I5w1307qFD
xR/i8eUH0Ya/zAfsU4N3/9Zad5lrnSlqsshfS3TSB4DvnoWm7Eq+RwG0U471q3AQ
hLgAQmJZpZp+v4wROuhxTJOAfwc92yUMZNrdUlWmLriI4ONZ+qGRaeATytzviHF6
LCKjbir5wqskoXHwWPZP1M8rHSSFg7zB0zF7GsR//owJUqROvG1MWJpFccQxfc8V
8Fs9th6wuRpxPIUzwuIS1JiwK5gRZXJUsw4353E3QL6cJuS9DbaZ3qbkOLMtMoRF
JK/96PUHyhBzkUGSf6r+v3GwfRRLf5D5sCvS3hKd1cA1QMCWKnS6XcArjdwkQmJJ
x/zBYFVS6uoASresBR5ORg2cHF9bnlifjp0VA5UIrodH0nbXwjw3BZOyi8OVjcAm
9d7X/SWDMNN2YdY+z7AfXmJ3TlrBuQX1U26mf4K2LjHsovi6XPU5zW38+ZUzkbbW
qeLPVDO9Qv8jPse/tx3XQ/xtTEoEGFb/X0Au/rmE5kbuFrarRfKCd4aFzMR6TWYL
b3dzXhIsnyfP/2AcbXoBdZOpPB7IhB9Bei5P0vc5lvPhG7PD1G8xSFLuH5BPjK4l
VoLJS9jwjXxrLfAbPxVWexo8qYbkecuo1dmOrj5di9VjpoZjgppAP4l825BPNqZ1
d0DMm05qThlDFTaE3K/KlBXIHR9IjJsqS6QsL1qRcRRX9rzz6Eco3X4pnoAqHB3U
KHLI4Q4dwMdHWJFlONdso8w3Ol4jOJka8XyDBVG/IvkKHLxiB6hxMttNdMWOUQbi
iXMEn3HnkBVW0DwjqlHBLo38TTDWtNPnLlMPleYy/rD7tWNa26HYjkd75NxGkqAE
f+nsKm9IeDfQv39JQCeJdPMk22q8OCUEljHsVfBl9Xc4OQs6Pkme1+hxBgOgRspl
pZoS3pqg1Z9nlb59ZJ/4su3xH2i0EYBmK84/nAGgl4Rn+yvW/1PdontQZY9QKWuU
PtIa4S01zHuHtf7BnKtRM7nlJ3AHKYJ+bgEEo6K9JeJqMz4oOgdWbvmg4uyG/f8q
qVJkTlOt0t0BNUhksEUKSiq8uX6FQda8CZ1Q9DykvzQnKuDFF8ptD/Vq7JZM4F7h
HGlz6+GoYu4SfpvFHjJvEgkrfWNk9BTLZgU+Bp8GUGKbBhqAipHx624QTWnD5pUs
Skajqj+w5nel7TV277YdzSS8hP2YsvnO8fBpOdpb8IEJ+dfjtmpFOR//oWGvfSo+
KBDaP99sE/tgaNOBJ4BVuz6xTegtOR7Z+q7MHCjcrl9DrYVo1XdWAWIFEh+at/mI
9W3U8vBmAZKRZu2Ca3vU0p2CFMTdtXxbWfkJNK2hHcUu23VBH8HkFNyHSP7Gbocm
9Jda990xYfIUA1c9TASnCwdDQDgv7S+FzttJwbTljJ6ug7vnqr08Z/RNjSCh8iZZ
ZP9Z7v+G774EiCv5pjlvycIG6g4gFg0iflX/mpr8+2cg2JZ2d8+KxWyMI6bAOy4O
2BW3w5EsM08ChvKk2mbJRkNiXFdqYeUHBPezOnPLvC57D4uFrxyTEZRscY5ZVuLA
0bYlU2XidojNCk+2A/OPopMEUh5HB9O75qZccd5cIJDPHi+5V9vboDCUE6BYDOmL
PUmdSJhCasP4HbwHQutKjCtc/8iAfjcryOCR3fgC2gLWUWqFR6Y51AViHnrcfoFS
TCTYhKkEYQsM351if9hS9QgGkwXTzrvDgapYYWoPKQ+U9SS14WcsRNb0rxuOa+nE
opH0b7u3a1QZVLJfbj3FzN/p3HcPJx3AUN7XbN9aRx24G5jue+kZfg9XJ9Yj1sWv
4c/iNbN08Zd2unmy6TaMmqNhOhJM3BVvme/72MyZ6A5oWTUnZqpboeRV0wMT2mZ6
A+Y3NUZzOZWdcubHCvy84y2H6ccflTMN9lHuBtwHrXq+0lYbopT2SRDIy/kEdulS
1ueJDxAYLINdQpTsBpIMhJhWqEYpMa+o4nQpy3p/jJ2VOUR0rxfsyPcxThyJkiRc
Mlne676HN6a6bRQG7ra+FzvtGOpHZ2P/xvMDS3tLuWwFgGcZthkq7jI97H8CS02N
RFDF0MsFaUkDXEbHPXl6gyUQsZNFliTyE+Yo8kEaZF+AB7lzxVdQe55hBTwghm06
gjOcJLbT5El200qn9LvU5rqpBAaVXnFIe2uEs5ai345Ol7OvclR/SGq7+VNmwxfo
QioS8dgF/KW+P2FsBPkmq1scnAlH4GVc0pd3tc/ZYQWYM8f0kDkdvdIshxe+wPPe
lHblcRe5xs7TiEMrfA4PwCJOFD6o0qtr2KTixzkanNxq20+4MHaBpj0Q4y7B2yFN
Ch6ScjCOV6ScEdh56J8enO7Bbi1n0qhkgvRzyweSoSOtdTLi7BbkiForCHa30RVg
KI6Pn6ahwH2nCGCi3gtVCi8ufZ4576HrIqmqYD1YtlGJkNlMbIKIOOsHsEiH+lBJ
OoxCp82eLn90Yj1R1wUQiP0yUYIXGm381fLxF/XLJmyIgkErLjwnUiI5pk/+GwX/
XqnHA+D/kXf2EkASKbGT2s/9tU2DvcjbtKIgT6hIytPTIpzMnZ0FS6TYyy+tMUG/
1vvgtWmGvleq35wBypUK2tQkT6VDlBaxUh1EPQOfIiZFps2Q9FCe+JS5ciuKbsnt
qLqNig5KmWG1wwIgPgf7CSoXtO5wX0kWkFR4cpd/OvXIKdwz6xab/f5ot72QlRia
Gk6HcEAo7CnjyVTgnTfuHO97J42Y0NsEiid4ay9wvgVJc9GIEWU82j5bw8rcdoEC
mJQYCM79nqcgyaxRhyMJkRsioMiWEeXe3r7DrIW6tQEmxPujOyd+TnJLgFKXLC0Z
4FKUDOTxS3Ysa+UqMgPiHfiy+bQqH/dKk3JvwX4IQDxZ9Yev65vRC0XZ4yVzruTX
0F9krccYM6v/ZTW9niWhAWpVLaSFq7QeDyLUEYRrINPb3eUyhjDZnsZUzwRtQuHi
80zsPmn2LLyZsaV85cxhKhiJ6V6n4i+zKefvuCwOjbLyp7krwvAAJRHI51ZZJViZ
IpJndFh0HcpglfeBNu3giwxukSu3dhea7fHzHhF4w8X61vzpHQjsAU4c9RDaaP+o
LsQ5lW9qoJr7Y60WfBo5HKWdyLMzMwY+kFwiIroylVTgJOeAKHkUsRxVF5U4Hgmz
Z/F3Az/zPXN80M6R4aZuEG6znLh6JhxlzJYvQBIKnDA4U6d6/b6Lm+NbCB2zwpTz
rD1QP1Rm9VZbtKy1HHmJh8k76D3dIk/85DrsL2pzAnH5OjBUGiEF22IaeUdji64d
8oxNM5DlidxEaVduzUcM6dur5uuuv0rqTfHzxZtxlzzSvFsU1ogAM55M2NSLQ3LX
3OY0NxIjNrQY1MDLHc/mW05b31X/ToX1I5CmOIgMubB18eqAIZLowpQpQd6dRxPj
QWcaidV4f3mqjdVbfdI+s5YNAz+zzBMIERmO/RIqfmDNA9FE58IXFjhA9pQMiMYe
HYTEw3hXoh5tQh/93CrfKm8CfuQHAGrS9nbHeqkEqzsKUUXz8+CMF4YbaNzPBfk6
CvidD66QASNPy3sE+h2rb961tyMgcP2J6ORSvcxlmtvmWEWLPFFLvhRi03BH6xvV
KJgJHmfLhCcmcYp+Xa2bnxga4e+zPsi9S53oMO+Ac2NYs5fWN7fmtPuzGR3szMmr
VNWaweHETp3Ttg2RCJ62Nf4zf/df7hkgW53NvQeAeeM9R58edLdfyqYLYHlQdrGj
HV2azYcwn6OhuAeKYb3n2DOShU40Dmz6JnNiHuPvV0nyEB3KYSsDIRQfAbB0hZLK
0mX5Cgo21VUxIJFkkZCs+7v4/Jz0puyUaXfVM3UPidY+H9MLd4Oa7zZ8HUZ82lUh
BRmV6Lkq4LIOkcCUUsWrdbkbx8p8QbDUaDESQVT7WtIGp5gkEkRE0Vuk+J9+pcF0
/MPu30SJyA3guS44d/rQOWxSiXCl8ZX0itF4BgfOeKjmWBVsvB3SbyLqsSRhzG8M
HJ3S/K0Ygwt3kpdrsj7kvrEBum7+JHYzQYQ6SpiYGrN1M2Y9e+2K6jyRtDY0qxqP
75hYo1+WFQoYk+AUZEpCzXbWL1b/cJKFqXYC9dUWECxdProlbQLC7ocwO7gYRF9R
FluV/ACLpiUhCwzg7MtKNG6B8il0gAq8CNMwpvvswfuke8Bpf4yA9qi/OhSqBLS3
X4JgF1/HZPZHd5ullxTCwtQj85uo/Fkyf7Xp8VpFke17Fl+BihxoCNl2fH66pm70
VtGUUoFXu+IyWaqmnlfVhNfv+cgmS/bvVOgMW8TrBffmEVn0GwhPMzKbXBGmwEan
YVU3hDh/NG/L7tNV0XNIJPvP1NX+M6yGWg+obDTHbtObZkQq68k9IeIoV8ZtKnB5
05fnu9MdFa/NdJM/Yra8AW/gPOF/efdX/bLw1ukxAI1ansgRA81fFZaT9b7wEWHD
GhoaK0Myj1uu0yAn1TU/fFl3EBhXcjGl0GEgokCn5NKt4R+Dg7PZqYxQSqyZiJe9
BmswwGqKZHRGff9j9NNimuLQXZWS73Z6UqJEM3zV9acCWQwxoh4yzo92hMN/ioud
Hl4fLi6LIPFcOiJwxeywnMYiPd5toIoLJPTEUusSCACeymhj7RusHk8qYJ/7z8LD
Jrh0hdRneF/pnHBrthZK0MZFz2kbtauv8qnm2BTD4XegPtknBW4wcqsTtCARlDLA
Wty9l51JXNrWKP9r12evFw1p6MEyf1SL37CkP1oxxdKAP8Mu97VAsXfrFzMZK2ZG
c424q78rSMeeS17gwdoa/L1yg7fXZT2iVfSatP35OPddy421dM+XGhsKF6CAfIb2
dj8lmRxBQlBmMy/kZ9XE8exlc/0i+9ryyIhZYLC1DOfrqLJC7hkqlioAdu1wr8Q6
uFJPSU0sppms4XPvoUOubFUQhis5qOOAUJm6Q49+Mzyvg4VqW9kVgeQxLJoYTqgB
eBdeC5ngCVBczpGa3wtrgkdhH6uaw9WzHFWV3+q+rqMeDUavZl2GqgEj/mpHB1C2
jOZRPiJBTTYR0m8A3YHYmAGLcpncVJbEOftIrS3TLfg76u9JNBYClzC6IP5KFwPP
OzW2fBU0aOTwxcya6QYIfE3nucUq7TzFR7moJtqheL6405ZtX3oxCUJlkNXkUEPB
em3w3Id1KLWu31ukG8ngJ0MIzZQ4XA1fyoqRFJqL+vYKjLtIyapc9Hy4OuAu2uO3
+R/XKX/MnqCnXYjF+nvQoogm8QCaA2qOCAlx/vZC0tPKspGRhpRZdXJyRMRqPfVX
FvodolJIGaw53sVM+c+9IJBUruaA8u9CPgy285TVxYtgnOk9aAuU7jtuquv4TVM7
lFUROYexApWbRUiPrI3YFhfewgD1V59Flym8pl2+kuVTBf1zKvFZjZDzsgLWARTc
IGhD2yHOpX9RgzhV1cUgRkhQdt/6x8l1Xc6xWq9+FxlctEvHCMb+q9B8q92N+uC6
5aH6so/eZM0+lupEJaXiHtJisAmiI5xFLW3BBK5QcrzujMkClcIsVrv7HD0giQcQ
EkmsIEhM0qSkNasXj0A3h8G681uYsFoFE5/GcCT80j5KHRe/f+HjVQW9pNgA6uuz
mWPmHT4L61UKXdJdjYbJhfGz9ULQgKPAPH0owTW5EJneHnnDgm563426keEIwcGg
iiDCIBK5B36EFzCMju/9Bce5rlFHJMY3QBSPp7xOy2hX33REMFhD0jFfYOeSh63Y
BZUydUMolImJbHPK3TV20CRtYM49Qv8/KwsRb5SudRD7NU9yx6StyM1aVeuGsu4p
KCgKA+O8M+SMEYhAat8MyNa6WyfgtJhRY/MgJAdJLkeZyhS3zyBFiRDps7grAr3R
z9l3bm+rvAlsRFWKTWvAf/voyI67wwQ5hMSi7vgmxgvxYFpP18te+MscA8D7S1me
7LyTty8/vNtRLSWwcywruRqWnmXBl896roz2CxHcOhnbgz75okLXWUi+/Wx++ebO
8nZ7ref3jwAOnXD6qeMBoD8LsHCCeXkkEX9KlkL0C/0tiLMfKT8r57N0Y0JLuGns
9MQh/xlQ6ZjFwcS0XIftG9ck/2NJFAwkuxE4pU1Ynk3FmTB+KzuH/Yh8hK+EGHTL
32PTBArlNcDConYXzEQyBtqApJPZy1SkZxL3nblFtjAnB/yahoYa0pxdNBhIWkLr
7poxl8LIWjd3c72tYr1ncEBOKl57xC/9H1EuGKlvzMSR5wqpJpB1eYFfzELmhNy/
HGrDEnhVDCZc2nITZDDdstyZL/VGge8HEdFdBeCsx78dpENxsrs78ybgVxCcy0hW
YSIgVM9f36fXhqkRMjPFm7G+6hmivip5m89+4xmJojr3VezUUJaAJCL7Kc/NC9AS
ozjzKBoMESMcMSGObqS++2U4yR/q44EquiIZv7ECrIeuc30xQK/7cmvz4L6+0gm2
t8CRlfdNiosJshWlyt3Lr5aBMcYtyx8PjZ8kepflDnSYQ694PK5nFXWAIyA0HuWW
Z4Kd9v86jOdPD+knv6BsuxK0ph/9mH0vUCA/KmXwsS78qXHbXkP791nCqWTWbCL6
VamsKZH027dqz0M9LCJDlUBZbmVvzwVEV3vhMRzW1yQsBHoMmRxK+5ZN1JqZ/NLW
H/ZHiL0AuJioSXErJK7G+UD8GoXFLXREF8aU26VMy7SMnAeuxXdJ+gDYTuiH/B5n
UH3P5xFosU3m/e2SDt7hKUapsq6M4yMMjy1vbl5ageOMzK5PDVkfdqvRYmlzAveP
mZUafLWwQeh+jNhPkVNL1ZJ22lH9B3H2mC8qgCaen7VQ+wzxOxzAbD1awmn/f0iK
LuP1dSa6mI2unCz9HDdD1+hQjb8EhJCGBJERbNtnBOMndcNQfalXl8361kuKfMK6
N2prtX93f8wzHCFRgyknikv2E1XM3cf54zs+RmLYu1apHo5a94rG0up92M8dpuxU
0bKhyEO/CM4r4mjVNVMJ48aoy5YpitOWnI4DC+oRLcVZn1m/AQjqK/kOEccj/dDx
zqU4+53sCU35402SsinM6dGCEaThhyLBzGfAMjIj1fbv7FunZDrn8qvQebrBjiFF
x80zx2VoTQ2LpW3WUbU2Z3zlKn0Gf/nVN6fIiWfEDbJQ2WRgyQVMNuDms/WBq1mV
vXxO/IpPfkf8sDGfq+ZGKUXu/fS/nzAdvX9+DtDbrtlpLZYL826ZGwZDs26rhUwP
NHPPw0a5XX4LsXJzwFqrwb+6wJnRAIY0MzFTxmOhp8lCNdjtMBbA9xb3GFXooqiq
pn521cOOOEB0Oyb6fKGGmBC9Ey93jKEu9PeO1NTOWmYyP4lZyJjYouJK4w/fBHkR
AMHsyF6tgc86PP1Ic4bgmEbPEtl0dMbKf0f3cAElMKl1BYMiAra4rjOedfey/ZuY
5XlsQf0pNwQw/FHYeZHTOhhWPf3qct/bENv1V35uxJkpZwx/fuYUHBDRMUFXCPfD
wt9NQnsBkqRvf9Nyv/VJ7udsKX/jcC6H6zQU6if27jOMogwv0FAMYBRyP7KNl50P
BhDyQIL9s4chDEiZq6sM+mzaFPnw52hWzclkoNs4GOXa8+F2MZCTHiOeoxkitxk/
SsN9bh5e4VTl+GuXlLeikKeJzddat7jkHkv+uQl9MW08JRRegezuiyVYqg//s0fm
qtjpbx+ql3e0+X+zTqEVpjb+Po3123D3NUXBfp9cke4hrcYlBpMsgBGCcKQC9IUx
RRLKVD5SqCWl6CnCjUniDlBXmw0FXWzWp6lRYvdYXr2bs/R+MXuq6C1NzgaeT9P9
D/aDH2bEyOQIh4eJc/8qDgKLvkWV+7ZXVi90zf18jAC3Eprn7c/mQer8pto5gOXc
yHakfoxXTSLT4QcnwQYgrHikXS4lB2MYpxi5DEytMW1LP3tOSxthhRqwFQFxuqeO
+7HM2dsLh9pwvSGCSJdLVHHvV1XF2s2VaBMZec5U7ZEiIDoMTmSKhfqkyHGrkdyR
Ibqh3WBplj0L78MA8GQwkevpUBKbeWUgHA0ypqpicIuMqlTG/4EaoRSbJ7bZaIFA
mPRK6ZBKrtcqwdlTqFDXfy7EoRsRZIHrp76gIjwNYEwNRzwSAOi7tVAuye/f5NX9
dh7EYmEbEyRwMaqSYmJ1W4Nu0CallmHgodCYk/3QXfCIrqg90ODufYT/Ggmt/FYv
yzc+LIFazvNusayT1ya/xorjEqMqX4X2rN7hVR/zr5q+QeXWVv6rI/tIPSeHZ6iT
mSm0W2AXIy8EZVq5cTiqzJAbzndfqnFab2QyEnhXJtzTKz8bRv6LLGXqH+FLHZDt
ndAB+i9foNMNmGG5fi0u8MeYdPzoqZK3LDjnV1thCCJ/Qj9a3LyG2rM/7j+Iq+2d
yDGet6WEHSFeARd7hQl1H4MkcbICBWFBwq/2JC7Yj3++vHWQ2MwjH5TH12xv6CwM
lpdPpBAYi8n69V+2SUpya5VkjKVXw0up/BMxR7+sYxJY9u1yIMWdZyTwoFTKMjZZ
SjPbLWSEsWwREHEx9uPAWXsr+Kgd/JJhBF8WUOZOYrm0oM4Iepwju6GrGzHa64p/
dOXHJ3IT5eOrirnyELN0ayJdHT5Ba6b5EPUd3wtkjqttwfUd2W7I5V+TX0/yBNy8
drurXJFUQxjpxDXIXaFzNwesv6vY3+iBQjtut2UIWHQA0q8GgOFUNv040bE7+cgM
pIWeJCuq0PvOV42oWVhIk6CG4hNtg8fSmS+lQw+gjuefX1HqaXWxaXOT6SFuM78V
oUWwleUwZqAc/P8aJr95+uFrz8zfbznNeUHcQz8EUMggl+FJt2lgfNZfmuUby9nC
auVBtsjbkKD9B/1qwoZiXKseLTIYmC38gUg1e7B8zZ5rM6M8q9+8IywKlhiEydND
U2SmdNI8QpYq4tMtrVLYvGEPoxf24LufSkg0twQL0QgoNEbNEoW+bRS5hNbQ+DL2
LtAqRXqTQsb3HONNSx8PyuUuSB3fS9yYa3BhVmr6lt9sNh5w5KDsTlUZsu210ZQF
5IvgEbEy+eS9SuqIIPxTC0nN/El8h1ThKDHhelZ5noODAaYBe1RnuDWrxJPNWyeN
6rw0JbPLtxX3AEDLZ1fm8nb3U7YU0BR3A+407vB7YP9FD0gbBoYeMxjcIOYq8B+F
CXjrK+Qh4yRHvMUVZXL4CVy0nGiMigvpAEIN+h9lH8ATVIUcvHpLKgWF7iJ0U1an
5mIVTUeziyqXxDosFPhfnF3TtoFzcROmh75bgqrv0UT1j5+9A9n9LIsFZpZQFrFw
B938qJUk5xaIKgtad6y/Jb7RC9/ku2GMWYgBAI80P5v9HKCDqDJzO+PJgv60KYfn
QJVDPyMBdAbUp1rW0EKf/bWacMcu+OpJXSx4NAq3fi8q3qTTgFCmjDiV/5NOhgZF
XrqBiOwFtWr0lHqCG4Wp4ip/H8dKc9ylX2fLEHzV06nzmJOw3zR/M0TDd+lz9YuG
1dPPLRdOcMJ3QAmm/IEeYdLHhD2IkolMKc2/mUr0c+dG6YOpu1Pnv6OgWPlFgLQZ
HY2YLV2Jm62r60uR4nkwVDC6wxnfWA8ou+RgBdGYfvrtOrbccfQ3Al+R+VKxfyVq
yUPCPQB40tMqPj3n8QYfiT4Gl0pkXICkS+g+SoCvBjJSfbXhn+cOA+lCMl/202H7
UGPnOlEgZkiKk9HenfSyaa2S4wqcRWBDMTyWvW1Dbfig3dnMzSRXBNEw7EjhpSbu
MuFjeRq+t+xlJxbVx7Uja0tCwtOsNxrfgrDfkbWA2n20nqv/b5YM8bkEMIkaTFzJ
jsMUXamUdJo7QQcwTIkE/gdcfREtj3PyBc4FPx8u8bB3PWnJMmzrCs/FlVOZsprJ
O2o7BQWlb/UoDPD+21fujTQP354oWS16v9nowOmaHwZqKgSHsS/YSQ5gL+thkr17
ojvit8O5fRtUCTM2LvkXaPBH9cGAxCLhiFOgxjzZKGjafAChIpNQ7V/gPc9CHeNx
FhFa6ISFPUKbxkCDsdEZd/ExMJ0bY+IYeMAbqF4apaFqL6ibGGPo6vj7FmUEapVR
Q8lci0s1tbzRHL0SA80Mh712nMd9Dy11H3TowDsURqbJsWLvRTtzyo/UtiIEBMj3
KX3fdUxuzcTF5whXCFVdrJuS0YIp6gcT9Pr0tTYCcffp2pr+IExweMn3+3Djeh7H
597Qo7mtNIFQKw53SCOs9hRgbEpYjXTdRanMuXgfCwzFmKKZk+n3Yft4SGjZVAYz
nzC/kvL3BMVF+eLQ5mfzXSATCgUGFsSQK2yw9K3FcGq8M/I3cfOBiafpuUM90RFe
jbogiAwO2owYTAFdMJTxI6T7hzYePQ5Te/0C/U4gvuTq3OWompz8bUOtuaUbKeDN
94m0aq5b7IGkzQLV5DS1obqTt2iWmbNEuDTMtAIYCTaIKNhJycC4wbFrABCuPG2g
rR5Mm8uRWtlsBDI6z3N+hiVA9Owih5HjB2WjoRfWlD+1EYOVxyRIRIazaE0+3vA8
vLxnPbLnoyKkzbRAky2z+lAWFh4kboTWG0y5X0gA7vtYOdRlj8aLWwxLSttJdWYJ
j6lDmEGSdIDoJJ39r1WCpTszvqkhuhBPsxtWrDdwK1hF81h9joCj+pC0iVC+jrGW
8PwFIK0bJdKGB1+ln/jf2MubJVLaRZq3iknnxC69eECsLqwmX3m+kdODNtXb/PTb
QTSTWz73I2Qt5vzzIz8yAF7zAG90r2fiqij6clxslfI3enhqZuvz/Bu0vB+e0LbR
7UGKxye7J4trkSQJtj147EFtmo++UR5VaDtNh8FtGexFsq5I0NTG7APxofml5xEE
KSUjXOSPIFvIq1ZZTPmD4KXjTCk8BW/xrE9LmNiKvwTzsV7kO3G7vlmq16ro2GvW
JYV08lLE93J4Nnu7zsAHVtGPFXIEtPNt2BooEhmEUBgEHJyF40tKVmOOIPiQLwUd
sWHfFAoznVxco4d902oE8CaKVvr+YREVDaWjqhYHyW5TOZW5Qs69w2Z2wl1vQEaU
WJaeEg/EzbaaqGBmv53BGXfJruYiYiqsVCyxW/sKBngfBCb618BDqJKqmWve+Z8N
nP3BeAMFGA5sT0iI12F7Ib0EgBeUsx44tmnmqYKCEVRhTf3697r2rIiNCPYLBkxC
+g/cEFoL/qdORNWGnjC5oJzDmirJ7WM9AG9uLJt2Nd3Q3PmXC+b0OBFCPqPQS/+0
fHOXLXCBBrlnoZP1GaBW6vL6aUJ0S6hG2AycVZYVcM5e5FIkswhvvrqKFLerD3QQ
wLiCW+SNUV63P+/KrUhV8//f1OBibkTZx0Wtwr3M1HtDGREyagHjRNGayJzfBFM3
NmYDKj2fCkn9se8GtJqASda/lP9YdNg/02HZpmGl8ziaL2aElVEg2xxst56logWj
qeVCAGchgnqTiy2EC6nqE9pyjzoXbrne1/BtCvU2K0dHzSfFKEgP8cpDvS4ovCUg
8PDofp+aN2czBR4d+3tT9p1AySrxeK/jo3Kd2sGv4E7s1H9R24A70MaJUv1yyoik
z26QDLKmMi8b7jllI1JzMS1j/1+4jkyOclUGUfF5iTMiIOgfL8V74EaPgGyODnvf
pTYI6/f7hk+j6kREM90nmhfpzOzu5EtymSBoUXJ8oA71R7nYPB58uDHKDbVE0D9u
kEEKZPBRzxqJrgUn7FW6gEFC18W5hS+ugQA5XZD7sLKXi03m+ai/aclBg4A3sOtc
0QLmbJrRMhVKSZ7O3TfrxiIeBO3dw+ZiKS1tZn+EPWyzlHMB+HYipZlBnZevxCXO
BN/CUXHXnxqKXZ9PWOHfM6Y6ubuYKwRUQzAA/iWSBSRXnTIudp7UlgMj4lJ199Tl
+bEoGUeW51gmKOpaao25FiMB+ORcEAOBsoPL+zOsisaehgZuQoWw4OkV4ew0nwWY
3mR/d62VIhwq42QrmOBFVEeGXPCOkvwJvVRgAuMGld9zSmsgdPM3EWS7qwjFzswM
rVHbBZZiNXJahlkLPA5BTGcc0CIUYM2YtgrLjkgDJw2hQMevP4uPPQAkPSOM3AzW
0CvIRi4fFSjjSmxf+3eQU+QxDVv388vK/eKJBXgUB/tUvcQtYmVtppONh6IINztS
GhzBlYFL2+w5tGp8wejz4C61S6/qwArvnWfyIyvn2j8w3UnagFehSyER47svChtr
Q7tENHbhy3K5TJK9cTe7K7RzMQBTi+y8CQULfSuOOuH3H9wETjTYAwSBBhmqJbnM
sPMGT8tS7D7Un0wNKQg1oJ+1kcksI0RyIuuDCJN39cRZTCreIfeacujVJ7zA0cI9
B3QL6puxAiJjDgGF31didEOiXGKblBY4VJpLmEMfXTPtIz5uOIPUo72lAV230f7N
XVRwcwKqn2LZlAxu7U/VGA1uN3oPKaJQcR/3K5wWgHWawmXTDiNondlnUdFo43V9
ZuhsROvd8UrJs8/ffJKsKSO+/Q4Rb1sr3G//6dwJYyKxjvEp26ne+E/kpTgsG7Yk
AdT5U2ijUxRnot+BoMVv0ZTUd2EZkpfP1/M3e3Y1XbY8txwx2RlXMkPjytBcFj41
TVT3uvS8aksJ+jhhaRNlgrBlTh2+wI/4hiNQBSyGbUpnjTSSWlLdS5CJtnDRnVMN
saxPOnfbJ4PRdu54lUwpG76vc657rf7InfG0lPHqA6LFjX9tGE/6R6b5YDeEt2JK
9eyLlyEJyuC/BQfk0QO7OAEVrztmJz+PjcjNBv2N/bpIRIANltq/OreK0Smb1AIv
BefrLRtti2Va5qZVne0Djj49lyhFDXv4bXCVGWdh5SkWAc0W34MTmK20vc7f/VEo
U/1y6CrEgu2/Atx1y/yKypdTU87TaQG+C1tOxDfwj/0OON33rwJxodWLQANKC0QV
JDU/jWH3X1poENyt5KLF1l9ymbExKa9NjQXXbJP9Q3IDTmha1hTQj0NuBsyXQ7Ip
XmMll6omvmvfkqSHtyFaniNedp+kZMphBcnNAM3BP7WJJZGiMLM9ARKgFONwQ2DI
iaTlxjcnKempq2073jhluCkZTlWc5eJdxUhYZzUa/PJVrVlSyLOqS/PAeoKoY5Sk
xWIlMAunOcKwO4KHGwcfNQsli979yuhlYTKalRh1iUA9CxqDMj6as4uhuacI8Xh6
vcNUjpmkJjgPlKMXMCRmVkjwI0zgaBNtr4LPq/mVbEsVhunPw5bvs3CJpXYhUoJi
4A+abENOHh49LYp2rQmwHm0PVR/W69k/Wq+lyJQiG2qt7dx/9Z+qxH2YxJhEXyNy
oXfaxZrnIikwk1qqlSbPMnKC5KjG7J5mEZexL7ZHfWUsuNEvEunojkJ/YNBywG4F
8VyszVq3E4xiEPhyKlT/5i+MIo0gtYB9dBu36pYTFtY3Hco/3z8UWulJXO2eeqMH
9VJOhQ1D90jxoIxIlqXhYB/cVLpG2Mb0fJus9nw7ObjPHnT3jbdZO3Jr14hQchqy
4DsAxymix8tygL2brjW/RFqw8hcdpJ8MnTZoqBRY0nAlVLL2VAbBWAnwXInUJiJi
FW/Htzm5My3i6ClGOtJeWAMsg/2zF6ISMzxmdaILYpiKemID/t8oFreFNBqEJJdd
MyBwQnvJY+T6b/bvWMZWt/ILPP9M09NAhi60ZFaPKPi/aSkwm1Rqf9ggGRJ6xgpd
Ibxwkgy98y0BqMa3kzLw/ImYy0qOfAEqNl2QIb5Ji56BAe2j3o1I8ZTHYSGOc/5g
uP5SWxB+D5XO5QIoBCgBuuBDthB9oxDahShOHNrWsH3W9CgVtfjeKOhc4wZEzFZX
iVerbEYiJOU+gEOPjUrevurGFv/Z21YUhwMtxL3em4ev25s9IoSa019+G53tqaAC
NHYe52EkwuQ1cjFLiqk6xsHHPOAIx4XiNjwcI0WZX47u4wcGogGjcksYowOBpFI2
rG5eiby7FA/8syia2DJP5ubfhq+vNuIsjs4Mm4mbZGGMxE7zf0ZsgzPkRmNs8BY5
N0hQ9vAjQBxlP4onhjdejY5DAuYoNdWBi6UevIRQcP0COfKVfcjbY+O5vsYGz1h9
rFUFuENMWBYfnTeng4i3TDHI9i6GfIvP9EZUgtAS7Z5k1Bqio6BreOLOXntrQykE
JNJzJYSX3F3ajXSAe9OxnDYZhncZ16fDXzRpMTHUz3YDgRYPlbStgMKd9yboxBO/
olT7lS2KC4OPvZJdbZtu2mV9ZNBW31itGIA+ZK31uyCdVhH6iXDXzVYm/XXWyyJ+
qvV0yvYQ/3eOdOqIvTHewI9PQzkMN6XCsQBgW6zBJhwoDeEmKUKQJZ2HzyQOI2Jr
cIf5lkPqMTFvk6/e2eLGwPdZlRJsfCCN6pIzvoP+hMjd120aVSN4RKDiwM5E1AAv
/RCqCJVv7WaG6I1flYqed4xsoFtwi2++TyorGJjvDRvAtlxc4XxHUNgw83sUApSn
QsbTE2Qfjnhsf98sSIfQbp0qdqrv1gF/I+nnzFdbP8NFPUlc331RwtnIuTsp5YuN
QUzGge3Vy8JTwyuk8nM9SfrfbfHdtb/ggeZJBNJhCXgCp1AnqiBVzqoiihIjnU59
gPH39ge/p8dTYb/NbTHe5df6Y9jKtaGGpqLRC8yvZ1Yi5ySnahCgzhV8VpHJ4w7T
8KE+lENJff/ny4Qk7kIgxG45+zFt+fPU28sed2CZslkgVf2eqOIXlM1/uSVNyiJW
Kd4oXYJilhHHZ+IY/vFPXVYZiUxfq3iOiY6/mAVRYCTolzZ4EiO71tX7ymC6MKB0
zaz38UyEzTM/a62daZqGLXc6aubOiNDg0ydms0Bp9AUey0yc86P/CZjZzvN/+yBn
dU5+veWg/FNFqtg5IsQMxPqD2Y92zHPw7iB7w9njnK+BZqP9Eq3FK3kBA9Qn8OPD
PzMyugxNStx0wahUt0sD1+MZJZg44J5QgLFoQtKDZPUt713YiqLpCmMaNzaKogto
dYx9TWEFa+Zu9m9dFGkZVFLitFiqX1o46zxDtLz6/s86ACjGf4PtnPFypnRmR1tI
OuFFhlWH4bsRRUNF0XkZ/9vzBhZbI8Kk9pQInSQXAQcHjkUnSlzGM+2nAf/LmW/U
L84pghoCUEf2nLk3cKXBWdRog2bsJCXngLdJQ85m/3IGepUHQF7eSV0dBqYeuPPS
/ISADepX3YdEtPQIJap+zEiDLjRR3vhc3h1sQhS5vu2/6JPK0UgdTRlmS+Kunitj
Co6bfnM+nR/bNqkLgXJmSMe2c+5dqX34DddzYHvAfNeASXNEqfBrqm0yHC9HyoLT
wudyYkCoPw3BgF5G5kE0vS4NWMwqLmQczD13ft3U456GYkqdPu+tD0jQFRPWnDH2
7l7vps3qssJO2+sEZrPQXXcL8aU4GEs52AzWn+rNmcS54ANpx+rFQiH1QgoSU+/n
kKP+yLn2qKdsomKgxkWJUM5m/1ZrMNoFpF/UmmoHbHdVc+DIe6CtvSjJ/cxnCI9D
Noex9kBw0UL2aHJhzg4jRAqyEUYNk1l3V2giiFFP/3AqVv91sAE66oLUb95b0L7j
LsGzoUz2CL4qQTQdcZXA+Zr7JRYj7yCpj/zmAHqH8xSAemreymoLivDy4OgNtYpI
jR7aU85Q86/l/yJeYfuYC3LssmmR51DXElV8AZAeDtZBrVGKJc99qLfRp9/HnrXx
50qepASmreSkvpZ6O7iqSgYcl4AvJvFNHl18jHLwOI5QBj1bIsRudyHEMtTU5soE
P47xd3SfMgjmUmDU0hW0VqUkghop6Cme1Cn49QRC8GeSoPzZC5tE9rK5wvm5Yh5+
jQkYpyCwDGKo4pKVrLKil+EEPs+WPQuKppaIeeZCRO4KDAFEtsYjcD+oE+qUj3uM
gIMuMYJKa7BvXVD8uFxh9u3mcoZhY17g2rBEaRNwl5kha6lVQECEVOpxzvDRkYcE
2VKWlGXbwh0zhhcufPqnhwNdInZYH6MYutq7cDiMWiP02UMM+feqFDUCy/xg4yY6
KXOMvJFx7alZcp7gPbJEUDcGDYZ2aIN+PS1leKEm6cjOlxKXrQOmpGBnpRqJWm/z
ZHUSGhVz0eCxJ9jsDc326Ms0WSiDLTYVHhr0wiuUnISLn1SdWS0I0Iqh3Xh0H2NA
ZpNpB8KRDnkwsYw8paa4LZbnz0/WxUMK0XPCyjHkpqSxguaEgBsbebwnlTZ9clw7
wnXAOsEXEWnKbDrbJzcpEerqsS6roKVnJ2IHxeYxd0By5a+AH5cAOAe7s4DzTdgS
y034mOxRNbHhzH8CHIA6ebT5Tr3uSUO82qwGTEy08plU7cRD7OqExKA4Fy5N3rF/
UrlELC9o7WcGsyLlKc93AQfLfvlDvtDkLIJAF14pVkOPXXRxY70C8cq6qzxI4yQZ
2b1Ix2vm0kYD5CyJGHVUMwmu2etZ7N5MrR2emkU41KFnxSe3ratk1wyNsPjzkuyP
V2VE5Lpj+dgal4Ozwmp8IMatZ9utWWsy85SGGSpaOHkm0DPUrRhu9PaXGF9DduY3
Bz02FWttFZxzmD7zJQyIWaLzk7PhDQbdwI1f9bFovKDQFyk4PbHBf1TMzDCAwEit
OtAajEYc27ofFKgSsggcjXDSjc0tyvhJgmM3xs7LgmTTXmk7+nH6JNoQGBtMZB4P
O+QNvYtb++M2uy/Ico0wAoEsHmZZVPa4BOZR/zUxSygQ1ClS7bWbB/oJ9ug3/oLq
BwJrYHZftK/RZYgVnV9HVL9xf2iqV709hpbaXrzja2LdvpKgeMEzvGg1XjnWYknb
XOAqTzYF+flPGtcJtcfYPRdIyGmDEGtWV30EaBmx9SG3cUDrNvpIxYZgdbdNTnle
IatgTQ1r4XOQrpR0T9QcALqBiv3DOVeWJN2XyFjmC+Zu0bhsvdUvobGOy5JsdSVb
fRwfZfofi1wMqfvIM4lJfwu+c0r5jOMw69aImTpPn46EUCqeorLeyvdiVjZbkMYq
ueCfO0VGFHU+oZXAH/cwSgRtVwTJ20lK/fS0c/Pj6qb3Dc7GnJETx8nmh6A6C1vZ
O7EQnXLG0/jNbJSqDYDCECRVZ/ULMdTx4bbUZpsx86gFZYIJlfecH1oyVfS/venk
ar/D1hzxmLCcG0tBztSAdFrAc1y0hnRiZJajOzJp5C2RRbc6ZN89UIuZz4YEsc2+
0xm3xeKxUiQcZldEGnqLXtS5QtuyZkMH5ivcYt42myGwf1A/TEpKZr3+MLlVkv8T
Xv2pANU3uqcpUM01VKDj3GlqV5yjhMnF+/zSKwQHXsmtpUx/yvWaVhaDCOo2Ev/C
eGYJGJnZc3H4zVV3KdBTF0Hwm572D87r87N6QZEW/waGmGLlijfdDSqsVe/Cssom
4wnTaTiLFp9b83RkC3/tAQ+oqEiVf/kouiTe31BXMFslCEHZqjtinUeio6902Kro
RVepKi3EDMIqej5bPAtKSFfp8XW4or9arww0GUDMYEt2KFvsrYb2yoRVYh/mi3+q
82h61hSx8Ag/2M8VXiMA7uX1SbT/8cbBj3jVy0hJrW1UEaZEqRP2d1WOpJO5wovt
Z8oF/RS5tSk/tY9a1ou4amOXWSuW4IS65cH0m0RKzJBTZC3IgJ+oIcFlmlpRDWuj
8whjCfzjRkb1H6sfgX0GTtU8ZCv4FEGpRwlJ72EEXo1825MqPuJS9y55qpkozU38
uIHDAIRDbXJ2kYa0itGI6wi+ejnnf/vo+kGYLTUs5S1g+MwggKKVnOeH6BnfsHHn
PYfDOkgXotdaWtqasKKn3IXZCDUR8+zlqiuYDgVyGIdGFMf9TIk7I7CgsYwZq7L2
oa3Zos24RVnXHJ6pGzCyECiemRG1pghLBScdBQX32pX2LSkpUqWf48s2EAFyKr4Z
nlgjVnePo+YeLX6PWQi5b5qIoLOZqXd0lktWlow1ZD+MqKZMLPhYeUMHjHZQlAM4
ONjNSKVHzgIfPK32MpXalPUPrhtME+4UwFMiKAMyYX+xJLm1V+3BwB1d3JaERjXi
hOYCoSPQQHB9VpuHdWBhkf0Sn4KIIMz10tg096qFqVjCfs5Sd1asWgDCXq2/FPpM
zZmj0mokcXL0zPxPoJN6+WksQzM4wk0czjdPpVFU4TDbCaTNJG2T2XP/hl/3N/5D
kDcIdFKY+yYPIukaFTZ2D1cz1AJ3mtqg0spIxex4mS/HYoa2mJS0iuh6qNqsmZTL
di+L/nEXtoMGgM9HRcKmj9VNVXSivE3yZWNaI2GcLGAYKUq0BwCMlZF7EJ1hpmF6
DfaVQaii3qfGs5H116gb1LGrJdrMn0wQfhfZxFPpy60QdvT2dCGYlr8ftaZ3RG5B
4QdE7WBuhHE9EqE3EVAjORxHXnNlB/WqCEaJTUiAHSwyUfincDMZ/xdFbaRovqId
3YlSVxfqxlELzKHstcVpjNHtdUH971gPqZx1s8k/tylRRxe22UWB4gDJ6rsLc7LR
0MFJSfuZdRkxifqmatGr53k2bbnacOBHARqGTy260tYC/vYyraZNNrvOXfeiH7ZX
F/QW8vumVLcnhWUFd2V4cFqgfBm6pqQVb9OLeN2OfCi/ZH4+GhSkcHz2+fvEI1M8
AUk3dtIV+wyDvazpkEc9v2px3aShYKdGjW4/4HmSd06dfVb43R95vLlc+jyLNjPe
+X2u9b27dlxIMOEixtZLW3BNDsWz1+O8WREVTQXrftSKY33BEN2d4SAdZqNNmHRX
nmxBSNT3vDvZqrC4N6aKc0AgcqVzgIPPfHWB7gBQut+3zHedycQz/azjHas6aQzh
+Zltb0NWOY4CV19q94mf4+OnySoKksyzk1rxfzLl9GKwCFN5uVDWgP42f8lV76zx
lobTzRx5htyevaQbWkIc8UA6Tpq+i4tQJBve0o5ghNWynR0rIEq6aAIj1cqTe+yO
7u9DFviDELR7MGDEchxT1PmM8EUywYZv1BUep2N4Njq03Cl+SRUT+2ifhu66R+bK
SQBfHL7NBjum7Hse0RX98uonGR+TlY13FD5zWb3cSpSAJ+BFMnhvDnchaAWKD54n
+NPlo8dhTPSo7eA5ULgB733lx51HOSG9Yp/uTaXW7geG3DrWWHjytm0PDM71o1Aq
cX56h9HOdfYXrKxOxxi41hzObOD1b2fKjqTePMf6i071xpyxqUatR4YKKC7GsWMW
ee5nez+Q/V20WqL3UI9WVwZXyQspSn9HplZTKOffFZhuJFBZIGOtOGhI2QEOL1IS
/1AszC2J9YfXnbTul3Mvz/1q+sZZSS3OZMgaicx9x6eJVIbP7JwSRBRoY2FTrjPU
lCEUIsl9at9oIdcSw7CttwSqYl0uhzSHqwQsqtZ4cAsbyyC2wQHJ/87EUhkLWCUA
oQINja2txzCyB+HCadi2gsTAwCJnYDoWXD3Q1k/ty5GMgZ6uTPkVEINb85/MsoAl
5cklaz28zpUKPTctcAdyciqNrXTj+re4dXv9NEUtJh/yQ6CZHyfR4igACcdajFI2
cCANhbpZAYNZAqq6FkqgxNht21iF6cjKGv6KJzw46fbzTsJenNjdNsa8Eqqn8Jmp
nzNUfdGY5Zi9KvPu4pDKqiOnTfECZEU9AFRBKBYwOtUx1k8XLYmH3pYm00cg58Kk
TopHoO2HO55tiPOuNg/8997AWT92TdrtvQY4HhKmPoz1X2JrDPXfIZIc59xRa9PO
B35JcV9JKZTRJrF3T6MPlC7xfq+f7HKpBQTYkTjN+kY23ThzJBYpbU45rwx83f+Z
W+3H6P/55r2KK+pHrPSrMUITU19vXk+eBS8e0U7VgR3cCzkIes89qVzpte+4X+4k
Lu86PkUKcSimCYbWp1uo0tIFCXFHR1GWK6hVGFiDVmNK5jtV7XQvS7d4KRwzEEmQ
wgTf4kPn2Tw16vKeM05lMO8CE8UiOs6Gn5VDpIjBtaFM4CCNFLs2gDYBdxUd9DV5
9fH65ijpGxbVAtXCL8A8VVYKHJfYaJV547mRAjRKyXGkIic1gxOEt4JEOrzpK5NL
dqUmAA+q2nh6MQJqu2ZJ5LkNg+mR+8eHC8q9edVEhhWHzMG+QG4mbh3drWDT+Ftf
Dpre0uo/i160hn/+Uj8kBwpqYhqI+pOLp9LFTRJmpDAIe6KCI6vc3DKO+KjV3EMd
D+Oe1krfEbV8y5VIEhlXopQVwg1IngqTvjdDpXPHXH8hbROdZ/uBkYeCompmA7hQ
nhrt7fnyRaatSbJfPq6Tr7YN4q92r+0HO8Km0WvDwA/S6e6/5Yqt8efrQDyHp7O8
LW7jzckazwDWqpFRacsk6MtxfAjVUNCTiKv4/JBiC09iwUY7bw1ChZIusvFZlYfr
2KP1EBEvw8+IURgJOAauTsBk9zYbEerVne8p7cw+LO2yDzGJ6ic5W7WmG2EtdaA2
O1AieS3MvPIeynIczXILVP4so0CPdSpii4r/JsLZwDFD3qWVJHvHRX1hMtVNl5XU
Hyj4ESNtUOGhwp6IeptNVo6Hd/Yg6bApPBxAH3Mlqva8IuLIIRPvMGCG0TZhpREJ
fQMBxmadnbSC+P05ZH5/h68IDb39x0wdVd+2R59qHCEhizCo9T0W6WDjqIA9cNQs
Vyt/QwkHMWC4T2wxzULueUB21vzM8dVqlV+RGfcPDsUj0oUnsNfPOQIVHylrwrdz
hs9P5mCpgWbbg6C2aeONuxcPQKtpvnBsV0mmnNI8qC0/WBAO6c3Ja2p3Bj9hd6Xv
MseSr206gfS0MfL7tKGY18B6wtJRndvDbT51RfTOD8KoQI1QP5OcEsPSVc/5k7Jo
3dgQEXMw64v+ZQUPACL5VPa9mO5RPiEjFH3Xoaz5PI+5B18IuRVP7Gn2bK2U5YyO
bbylFWjvjLEmgwG/SkKVcCu7vDc+9Orstw1/J8hVDz5zfW7uWWP8DiaqLnUnCKf7
kClwslJOrJirPxx0olEJ81RXcr3eTlU71pQQESScLyu/ZbkneuifZXe0fLS+kEdq
t3oOX0UpgQueQTxTAKavdu9Amsd58Z27Sv5F74gCBhUNE2bddQ9S8hpLyBReHJwH
xU+Up1SvNOXB7NuMjq6ZM+s5M2UkmEzNyOqEI8E0M2GXUB2nfZdZpcs+J0QkJnJV
cqD5kk6lvT6Qj4maIZjAaGLV4aisuta86jjwPDoWz6lwaDAiMLPmueJYEQGO6Ysn
FxHvA6MuPdCt/B4PLwZePGw0JEqrf7Rxex3paOwzUjewHUqDAiQvDlNlDuJakf6g
3iTbUG/93gh4LeIaWG8Uk5DSK9nZCcfLRhNt4692wn24OkrAbe3Ws2ExGqLcRN3F
ao6bmY3rTtdpiZXgSpmliQCuwm12GAK/6si9Q6gQG1A7NslcfJfRDLZ1ibe2svUf
rn3jragzf8UKfULX5UWwQ2gGtb80lvJDOZFHNa15T16pP8C0Q2VJyEcrI7hOnXwm
nyS3Ckp5OzrKG5arSgP0rO317xHrU/pU0lNiObssHeboPLnjw6WFCQZtrtlyhMdN
Emb85fNC+hWKv/i1GQjqDYru6VGK9hk05GBxYXVXUDsB0ROF0rE6QY58lKl2f2+a
ezYJDV9867NnaZeutPRaeSgRS8RSS6kxRHPNHNbyKZcJlid2pXI/RvodW593Wgso
dyBqdyUMz7U0LjUiO2gHpvB7HSQXfCBmIM2x7ikdUwrm0fa2wbLAEUXjYfBglken
M7uRm5QMj0Q4wRpBT2clr7OR0JqBOuh7Rz+OGkARre+92cEv2lIBet1oLoNVMlOg
t8ZRoOslZtAGZm398gIZ29NtonQ77F/VkdvrAqR2rprvld7FiR2RmS3t/DcKmX/I
sRu7PWLHGz8Q0YIRAECvL+otyQXaxdfUasaBpCiw54WEGx4fo8JR7WxcV5wFmReQ
bh9i/6epX7jaCfS7aH7DQAheF43NYxvo4KLdUs5t/QKxlK1kLqj7zF4gU3h6oTV2
IB8rGD1XWW0uVhadejBy7NSZ6RBXFMC1piTj1dw9BnhsgUBVnJouGiq3O5uwB8AQ
W2CQBGERWDdUQgjSwLla2YOpjf8LgwMf0FBFWYxPe+B3khpNh4JnLmvpLAj5G8W7
XJAhbISPTm+XjmKe07cnSlag9/mWGuhY6tBu9/v7uPhwF0nFCrRrAzY3USIRENyX
bUl0ik+lTZZr1j3dNPxL4JKx7n7flGHk8qEmVDb2wRostjJ7pqa9oEK8adXWRZs8
mVVc5HVC69ekoYfpKhV2rHEiY06ULieOvUefTRImnepYoWsWTwTWiI8CwMX3GhLR
iNkoGbF2He4eZ0L/A7+kzzu/DoucW3kN0eY+WzxqTxUPmECRvAaRG7DGpcZqfmFm
8aauDMFN0AEFHlV2RHElkH5+9hDfvJo+Gv6ZhLJN68GZ3tiD/MdLbMQ2WH4bPerY
o2o4KIiWLUwRWzEYOfFjL4KW6i+VUxpyWGXTYdRZ1nIj+//R8R0lly6JPMpK8mrh
2tC3gTn+QOc+sTw8Y5uik6DLcCQ62/2q/kPpraVBfLH7ZErjvvm0fdWiln1aYYtW
9pyTPHmowCvs9rOOeTJibfzkokiuWoPg13NCXXx5XKyMNnD1zN3mXOv7rY+oN9fU
FI69mkQtLSWGD9l61qtyU8raW89aQlsIoPvWZQZ/us6px7S5om9J5AutNzf2VMW7
5mVXZYakc3651ImE0XtciZa0Jc2Iw6iZONfhzNjdgcgGtF55/i4SF659+VfsZsrf
G3TiSu8Azk8JCW1KyMJ1Ly224uwP3dG0LSAkZv5R4f3kOuspbMRt4bJHUX/kqf+V
KlXZ362lSkB8PoD+E4tLSwQZUJgHhCZXn4W8xuzXTuxQjKA0pfhs+DhXbC2c2QMG
G6zQWV+kX14671XjgVX+Tu9BCaHpcRTv28u32RjqQFiYtmITckQORkZUWU/1XNgF
Szqz3fS0JfDa5wyCWYjhync1h5l8ErOEfMmU1DtWeCREoZxoJnyj3xsyH7LFz1oB
bWIssiCe7ZJwm+tBUQN3oMC/FDbzcKBG5SaDFZwe63DW6+qOec+pFJO22cHgJmXK
w/Jo2WVAl58b2oCT6yD2k3ixiTBGWJmzDknFx3iBpN6opAgHHY6PxbKUSSiT3ouV
S1o6/vKhJYXqT6XOsMb2tNIoG9/jd97HBdbwrHDa1Wokz7AjLNuR+ManIEJYopCY
Vvrk3tsS5pbhOyHQslG12XnOveQjTC8SFzhLpMxQGcDKI7lxQCbr0FPZlQAdALAN
am2Hz6E86B3Qq1esJjknl3egpqOF+99soQkCEnLX73CIcwkKmPoW5gYtXXe+PxkG
jn8PfQ69t5h2EqgvcUMpJ0iRAHXgu1lLMvMqqMl5c8Mn03bx487vacbEMpIZph4s
Hsl2+pGm9zpGjkLkcI7AOlwg9p3Wz0h/0750FKy53uefIm/1WtfyawYKPi/zIOqI
8uBem88TcUaFvuNekeBj3/aJLonhl/SxSkeyBmKTN/AADBOg9mZypzwoLdmL7DJr
59c5LiX8qWAE1mv6K+6hRvs7UAyqexFo0rRMsjU+6dD75CatdVNEl5oJFTyopNt0
ca2kOkVsZY3d+rquo07dFau/7XGTRdgRkk3IvejGDUROcnNy6hGmFiVDw0Bvhd2K
gKsLhOlMTFzD3+SH0cAtycHa0OIVjB6s4qoIi5xk5QfqGIBfXAXoCFfN3XEkEJdl
Q4KIjNTgmlCOal7LgPgM9300+HR80ehn2esKR9ZDMsrZPiLaLyvXO1iGDvupmdrt
vYIc2NA6ALuhNdjrx2AND0XJkoOFw5GkLdzp3GbxR3/lCgqw1iSlkkIy/Y4wxMJn
Ufgruxhh1q3D/cKppoTAQbXiRuSLQ9Eo+YCNvqtaXARJExFuha03bnjI/1PD8iEs
ZbPSwGa7ZjB5KTi45pJDk/tAH2w263qKCviY3ahYtsq6pDSOR61xYXskM9E4pMt5
uu522KKBPi6c5l1MJcxjz4r0JALLQ4EfeIaSOrrlpXdy3o14BoVE1427ohY7zsyy
OAwSFfl/kZZCVOYJTjlmhIFbv76MhufH1egYU0gZ2sV2ujcj1r8emB3OQa+/kVr3
w9ipVvN0lp2d23ulNPgAKUmvJJ9TguyTiVTGt2q7DmeZ4BsVyVFOyLTOU7a5hcYt
FyOo6wuKNlWiuRXHG9v5+8XGWgsYpOcVOqmLgVLGy/zb3fIRMA9cqKW3+J9q3WHI
FnxGPSvpoJdJtNc5aqTOYu+oQrHjknqM1Q4KtZFKR+qsz1lXAqquRDStavnn0/dB
xFvWv8QeoUwSU6sqTPtvAPWS+e4kwYWJwpCvLQOpdk9bULFywlcQdUEGuEc5dyJp
Dx0z+zbafQiCoPqgriJAw4/GSsgg+OQZOEFaFfZj/FFkA5WnUq765WlNN1EVrpRA
o8eiR+xyChiHOFm+SSIbFp/lx/14JuDne23IcU3gxCgS7KPzZzSmuh4Ti8UzvbWp
zGoyqsQrmPYtgqR5YhQQ/plxysZ0+JVJ8R4DbSUl8YCIF5DSq170qFXCDc5VJAnz
AgW9ortoOIjNYuNyq8PygE4UywiU2EPZehcm6eetwVbcycbsFlXBDzrvHzapvPrm
t3nYPWYghAGlgak74ALuGPz5jGR7S9MBjeAKgtrfRX480X5wZxH0b9JNJ6cV0GXx
SU4LVg9mqXjkr8Y44ZyUCiv+znhPuGKkTwZsQSEOci4B4kMuvFbr1T9PfnzQmMxf
EfwC4CypLh00SWV0ys4OiNoxZqXYni/HJuu6wwyP2A6wSZ/nNEVeh1cxU5w5tLfb
Uo0MZx6ircwrIQdpRSq+ZbB+R38a8H3gjDw7h+mirXt8xuxbBWfeX8ZAiazrazHT
KCKy2dxH4YtHo/cjNzzOyMLjsy7fEjkqTtdo6IR5WIvcArsH75IWeNmhV++I/PVm
ZGGhlTKIEN/zTpfLtFtpmnu2ca3xxukzymAeacDt+6kVFUQdSKBEaJHkebr6cvsS
9AGzI8sRESZRVy9S6OgEKxi5IPeHSFRupFg5U9PrlBjpgJnCYtZiO/VIvuQ3/IbO
vj/okf3w6zDUPPaDY7Wd9igZ3dEVLZeIqfzgFpgh0dFKtmv+EfIC9pEsgxv4njuh
tGAWeOL2gFXvSoE2EArW3+OISePeOWJo6oVJEAD6HMqg2KGgcX6hik6S/e+sU2lB
w+K88cTOc0faHwniV2zsGtWInYvZPCeurDZcNCnuzjXMYY1r4LqIxkl+ttxTBlZ3
y3FbD5A2IhetBluL4TfPS/9qDggH7Uv6ACHu23x+xAvQFscSyEhDSAXPhsRGQhVD
X0ALWLjn4ATjnWMpZ46Iv3f/2Qvxi3s9OGGeURFKqwdlJrHfbGf0LoRHDQYNnOVy
ZpM+5j02ZcsuPMAQYZlg2TBhtUfRh5msUvxYg3A6tZPOb9LOdNSP4E9hUZpXAoi0
9CqPiviUkXnDLsqaZtOYPEUor872LmO8sHsrTCuVtzQuM+AFUErqG9zD2uiUjvvy
jKAljOr/xqtOZZqfcYpMoBgxydpb/lFIoQcBOy0Q8S4dll3cayIZ5soTzlcwNkZ+
5NlOx9rBmOPzHhFeukhk7O7sHaIFFS7cDXadsKzBJG6VNIXfZc3w1fOoptb+Nj+V
byztxdlrQsw40yCO5NKEjbPEpscszALQ5Q9y5B0VxgPwqOLQgVs84okOdo3zedRU
ErfeFYVn17UZPu5NoEZnEmWOYrSBOS/7Q2aFFs653K2GxMbxPz5s6MeiVZ+SDY7q
epuFIO8azPiyh8sV+ygU/exQxxIdK7Z8/97yZK+SeLetNFDZJSe1JZaE36uEF82Z
+kNYmXkzK9eKRPLnabPXjy8T8XzHMPskoZMZCgZr958PKK7TGMuPLoFN1xKqkAV3
fTzsuAwTNKRYTZmZCrNDCWdGgvV1rtpxiOpr5t67M+J8+UnaMcLYR0lnCMnaQDno
EAKcQjE7JsD1pfJ8FqXrojnyyL9DDCRTU2FDBKdVcQ55ZKoPQa6wQgdGKX84tfvn
exrn6nEMx5s9+rqdVQpsGtZizVigUCIfdJqm0ix5bACg+xjrDJb0VocpRDV1/7rL
pxq2E1n5rZ8M09AjZGXp5Kk0u5IenvTUVW6KYuSlpriVB5R3Klvtrr1taAoYLZMV
wvxIfPBythX1ftgh9Ia6OK9BecLWl4oTkoS/BvxV0eaDHYqYSvllIhZ2Y6D+1Jcz
ZqKP23MRNmVWSnfbjVGKIodZLlj0iHSRjBFpi5+wkMnoTkMcQkmvmM8WJpHvDf1B
5N60OJTe8/uZZLO/FnkvfY4qrGb/KoGAGya0UYCMg4+9D/4i0pE3Rfo/ivqFlJGf
XGMuvHndoWRq5/G4D4OGK/jU85V9e5mAhg/l08XqiK0XroRXdM2nV6x0cMDek8/g
m061GGD1jTpvwzF1ggoJiNWwXTHx0FaujraqL5RSKQrPOeqlhgyIkvv3+fLawNsu
4GW9GFVwVjVjLKTIjb5w6NnIaAw9eTk0AvHDYE85QZo1PrzLlBE4kR6wzrEIdknb
CygPGNAyzUnSKweJWjiM5oGUmtEk7tj+c+kngBhLcGsh6L796sx1dBRYLJHt/4DG
cIEiwtSeMKSy/GNXQU/vpiGA6WCImMsfB3nunwxiTsFdWTjFAGMczRvamdbj78un
/GKJjluPPYHofocbfj+16ZS5h/8pGtBk/r4RAsdmg7DwawxPB2Aj/6IrwTGB8vkJ
D6F+VZF7PO4Mag7gtkT+Pu6FJ20JLAYNqdhQyIPRhveudsMlkxPyRiqIPrf0H+gj
7IY8cR1XFGs3X1vhd/dA8BOX3gP8waqU5tqzItExrdWwF3L++QU2AyWYCG+T0yuG
rTy4ho2VFmzZ3X2S41JQtvbywRuHCOZjlSNLimeqJXnFxjBbywGw2THa8++/aFnr
HBXzNuzMzNkRhUg7h+jCh77DIPrvRDqHrJzxumPruEkrHXqjIdd7bmuuLbFWeLHp
633XnLjPSEhsbda6Sz5u9vw3ol427rHlH/SBscJkhmZqpmKxntgat0d7HegLz/HS
UzykoJf77eoevF1DgBnBDMNjmwhqcfN8HDzt1FFgg1cka/O+mbED0utchFEmse5G
KrAnt4vPlcf2RdeNAj3JUlMthSJPvkO9vRpj3jqp5mjH6VXJTUYvnKDE3z5RS2Af
xMzNIOWylhrHOYmrgr3v3QlrVWazvZYoZoafETjiFYFkHpdsEOtRzuSqTp01up+X
MeyBI1VMGjABtjX/RwwnumXy5yKpG8ZurI5I7pnR3J82/zqrIB9N4Tw5mapQyg5H
4RXbi1XadK0TNFwYJmPrmDSPa+xFcXFH7GTtcnRGhMaWGoLNA5vFmJVRqAgC9O1H
2jqB6R+VQA7y5oTJ09puSBxysgjeqFOedbOpdWCowadlzoygcfseDMnfwrhwa6g2
5BbmVW5qiNqz1f1cfVN7thGtP3QtdkjyYHt4aCL8Zfsy1WPOVIq37ECxgovIVz+D
t7jThae9OXd0RKw8v7OeX0OVqvJPpg4NyEKJlJhdbw1I6kBezIObrizpJSTpCoIa
LrlXIbtaGUh/C84MIcKqCGzr/pjpIBt76h6jyiNQqtCqDVgu+8s2UEgeUNmN3tXB
wEvZG3QPWXtDmMM+/3BzGVC8x5P1zlMNx9dyNRUyx5chXtsWheIxn0pgbgKwBQoE
tyORvRUuy5Og4xT4X5JEQRB6v2tt/gVZp1phCdi5Ybhexr1tAxspnjrIvff4Fq2H
tpQH4eOIDr+b2e+nn6HdGlpuNOuT1pQQncrLhFzVFsaIJs5AKvr2Ua+mszCgDzKP
LYJush37qYQIf74/7xwuvPrbH6PBarSrxrykKfxdq+N8RdvLLwZf/Dgl1eoPhf+e
6IN7ez7ScuI4xlWvhRM22HO7LJxue3iw4pRjWaIjz+Gb0xuzyznCxz+E29JXJ2lh
3/xNk8fjlIQkopvdpNqo7IToA3RiDXPeSF8RyueElucvA6mFqd32Nt5kJPwLxRR5
A0XNnRYeS/Uf40K4Wj+oFlboOx6aLW/u8K4UJD0ggB3AcZzxWwdjJR7PICfYsI/u
kRNBIzSwYKQhahNPYvxVG2XtzYcgo6g+m9nFrP4R5W35hhF0Kg4iq+I8tL+J5xGK
SZikPq58AyE2ckcVO2NqU62CCc57KWvBPxybHjqM97a2c5orkr0HYIoIU62IQatc
dWKHM6yrbKQDOnf2Wir9MNQvBbolpdRnHfvwaFEG+CugCbQLlSukN+g6DdXfqy7S
A8B7U+RoCCSkfGrtZ2+wJMVCMT0dc7GunNDN3QrPLmX42XXkyhmo/HliVCzpTIAp
dE5WheQOGKjjelb1xs+GGWSJFlrFKVplHxSMCAKf7YZ0RFUZxiECOVXDXne61RW8
jbWHPOIGIuLjLThMDiYWJyTTtKn9LK8LZnUdEAH7l7Gi8+7Mct0I/7l55/ec3wpJ
OmStUy3Oz1Hs0CO9CHnPdQdSFDwyKbiaZYdFAjDcTW9Pkb6F2snKq/ckANBg0/ux
mEnGr1Om9mzYSdMZV/WUiPLeBaFUPeXzxLpgJxC+7LG+8tgOytTdzFt4vr97CafB
eco2g6RWd6IWhxe2gYlTqFnrrrPtDCV0abRzrc0jKhIa2HmyabAraIhdoz07lz5C
fY8gXOo8HU/l9S5YwVap3Q5tJ2PNBgvc0rixI6vdTgTmwJ9bVboPLFiF78plLToK
9scxAl/6fUHYtMaCE4sPxGZiF8CxhR0YP2dN23WIKiauCncY5C12DrgW+3zb+lU2
RMXy4B9PIU/CmME9I1uB2EXpjJUsgIl/+zYM4itug61Gan9eFFkITiiebBB11FhB
iSgRrIosg8DNA03FzJ8htU+nM2QxklTOYEyW3kRzVzWp3KCnFb/Zq60gXb5nOFLf
SmQYpGG7z2d81kifzAOJAJyEABpUFQ3Acd07b9foKneKH6uXaDN6kLq85S5wKTaJ
vGqvIzq4vnz+Ef4StwLO76aI1XJDBJ4WVzSibX5yB168BKcxwSG3J08v30si6UEN
lmCNHbl64lxSN+ounL1X/f2YF02kPoTd55RtXS94YYHO29XEiC137bIYpzsOvdeX
iiiqUTFPdJFsf4NcgefqtsY4+PeHqJ3F0GtunzXm6tuu+4pw2mUK2sx42rrlNNIg
wUphseep8jTMsk+q9O+csjjWrj0EGOQx7LB1xb7M3rb4ewp02JQe09ef+7B29mb0
x1csNeZj14uBF+VIJ6tUFORA2Cuth3wwYMzSpYPqbupmqarWvIkrynoyrYbASXRl
h+R2fRM9UVt4h5iZ3Xco/mbrvl4WfEHfJGNLiUF0jP5Poeox711XQ1JAXKL/9Ttq
GnEpP14zGusklLJJJnKV8QI8caz9bMb2WNMfEeAAxZhpMdMqPIyVRU7dgcYnEVXU
jZYb/pJMXK3ZGTaWMlk52rg9L+GKjluNazVg/cX2hNJN8yoo1dk4IITy4L7eFFfr
r8w0b6z1T8LKVs7q0KzWB7ecUXyDhAmUWQf1XMy/0TWjIEn29hazevTSRQK69t0v
WGFmoML2b06dDckAIdCPCTrcm63xgV8PRE7C7lGZfjr+5Dbu6iYEkvoG5jkdmAl5
3snhmkpRyTRnpxrzvKtKEcUDLb9qRdgXpe7DwBRgmbidftd1/BsKGbepnwGa4bKc
D7CTkGEMt6UCImSUtt+5vaTOXk1R50gvkrb61VUcQyDTXUsJHwF2kOul7FwNdoXN
guKpcjCYDq6YPCVE9mQ66o/VEgoC7ND3g/z++J1TvYt9hsJcUZvm6pOTq3OoNGpE
nyOGHspEzbEQ8Ce8BqwMvWawS1Nb0Uoqc92KtY6lqyTwV7BhaGgqB5IIWKTU7IwV
+JokBzhFDiD8q14Oq3FWeOAw4fEWniErVQfIudX4d2ZqyRRPrM13EF0vsW592VTd
C5/eWQx0g6K8+rUN+u7pQROMi56Q+xLA783xxtyNye0vj7wIdc2yCFwpJ1Jv6SKb
As7HyNx1TMcIln82d+nOT+xMJMYHQZx1pa3qk89gyJhCSaSML8eLct+DP/2ksnxu
oc5Re9nRPAqUMQpW4uegocf/q2v2628p6bBUWP8x36DeaA61kbp+T4uvhemFGtQb
hU7D98RoSrGVm513TCZL/2uzzdIm1Ezh74s7uT0jKxI9qD926lNp2seGYSyAbctM
LfK07RcMiVFFKJMGFCZDAJpZvO1fyS8ns+Se7VtsMAhonRc/fs+qcu4kZvCfGugo
q5trghhRp1EEmiyqHK5jY5U6zXAZ2Y9EORgENdrSTjfPwWMdlAD4YR8LaAUd89x4
mYQBdErr/s1WqVfIdM8QhGIp8nIzBLd4kkCYcFmOVWjltBVnermiadm6XsEVksiB
aJRKQxhD0NF7oVMLLXHAiwcAzW8/lZm4RKxx8kWiEWxDa8HhX7cXsSXwifHdK4PG
u2L8AAXfLgybDDkLUiVB4e5cyAiYTt+hvYlWaVxJvXj0ForqLMWmbrypQB9wT9M4
WvihM/s4rTFJPcmW1Su0tPq+HYxD3/UasoKgHXYvFDXEKmyDm0JpD5m5Frpl3iD9
Xzh8XtsyG4dztN+lMn+toJcu+FoL4nxv3GKa3ovrcooECv7OeEYxkRs9mJM5D2eN
qqOYsIbBL+FWpcYrlSWgCte6C5FsHOpD+TIOzYNTuKu6XlChy6efVl7naLC7eJ6e
QMKOa4WQ7vPXPf/JPB8OSl2ZB4nQhOECiTAtWrfhxL1qJ77KtB9aGE4Ue22B/uR5
+ao7iNjU5W/EjSew6N1etOhfmJWkCeSxFewKAo42lEpuYG4ZTaNkRoOvSSMx6kXi
Ic4VJrn8Rj8fLMk3j5MNmi1j3b823e8fXO4jzGXnXgLB5tU5QUiSvEGxWKyqwVLX
nTFzYRmq0xqupyPFfCg9XqxYj6Q8OAFv+J5O7DSuWHMxrlXP606lyxtduWtg0IYj
Zw3GRJt0ryHRjLMByzzNXixXsKLqVMN1sEYae5fxIu4HIv/1amDOej5crED+O4WP
SSTK3eB3ALcgJgb0DXQkkF874ddwj0pMaLXZkz1gYrP1uhGig4EauskTH5293J2F
BMHqlQOfnwxM0VnkywgDpZDjAoYtIUTmMmiWeynnLFuzzOKzVmv8159+hJ1cd7GH
yCuHYabFQhDSFWYpzEEsI81wB+milHyBWwW/LT0NqVxdfhc3gO1+lgopZwFdrMUX
IsMCAK4WzEPENRRM5Ep71XfuUiwv1sf/UBWwgyc0duPqoFvJ44dCHU/b00ys1roT
TKzMeGc0G/0aO8p1fNgTU6x1qiezduu/8nvBeA2WNCNYKqXjF//fd3zwd07BnuHE
4vYGCtu5E6nRFARVyOrQL/7b31DxhR2pMFvTCASqNgO9UZXq+siCvTD9RDBZ30IR
ftFYCmIMXWwl0fbGGOJkYSEG37c3w54f5sgfPlJcuZbAW0KnPPr4xvSiBz1GIPbr
0r4zuFmGUs7avYLD8bAE/tcbsVnTvgNbEziV0zm2jLOOuupXshMPUPKbsRrqtoA+
AbhxXs6rX13wPvaCHvmPbeolKMcYmkjty4tKStOE1SvoDL0F1reCZgHIk+4ugaJl
k8IFd4+jYvskKEXPlG/YTg9xsihGehrYLEgeECdH5dTNaXZR1Ih9wbNJWhaREDHe
xK39SPgKQ0QfQt2PJjp/lK7YUI3JxodxIsrVLH6JXc2Xo4RRmYMzglHO0Ul45vfQ
AHCxW4jadBNMx0Hrd3xJJlcnt/ag97oBXR1zu82Az4pH55DWKSBOxiCg1nyn3Ypv
RciryX5QV5An3XGMLUK4njG5H5aI1w2FUKKk3IsBeAzQIDInvGT5aBOOZAfD2rcE
n63Ytrt1719aY5MdE6VXDp8OcIe/4bZW/uK/8qHtPQ2CTqRTBdPsx36CCXoCvu56
Fmn8iXw1GzWjWVLreWSZN4A+Iraf4dwCoSuJEkhzbPe3Z2KdDNCtKzjISS2wcPK2
EgiBi4ROUQCnnwCdyBEucWyqZ65hcOo0GF6dVfraT6lyqyO5/3NmkCP+m7Q1V9mG
3gOc23uLwenv4LqdEopV9dp0O1NrVK+iargVUeI3OpmyDOzspx211ap4LDAGY6EO
MY+sZawvC7AA3tPrxOaruySzkM/XlHIw8aqPlUv/BvT1pIW6LkPOXFmo6MGj9IkW
qEnQNZhma/+22WG2xlaw1VPm/GMJXECu6X1lwwE0t2l5wB0hL69LvYnV7lKMoaCV
VEZvg49PxaA7EYxaOuxHIHigsUSh2HQUFN6tTnx7jbDnOaZNnZnc5yY1Cnvc36D/
Ob5Wh6GqOx+PU8L09pQJ/234A9zPUgfif1YK5U/3JmmMr3QAgnMXhDVERPlKdXig
PFz8zIdnf9/Dtlg2J2ZyaIPb6Dl9i8LY1WGqcKwViEDGlC8Oko+MCY5Yo+/a5nVW
Efpmrm4s65dL7VAa94Zz0J9KZa6UN+xwHYrFs8D2TgkTQwHJwVNcDbkTa6AmLupP
GvCjmhEqt8ngpwq0WD6+T0wACoM9srFIRJn+czWQL73v7m1EbYgfuZeuFeUjvCXo
qtJ44xWdbOCCXEOoXgsGOlkTLeoVF5EXLGwgJaJ1135m60EIVH8ZBPK1txy2i2Dn
2xxMGT5+pBnZK+Eey+foHKxqhfA0rhV7HFwByZfgTeAE79HvNufxYsvblQuRCCPI
kutQle1lVmaIjTAVTe5qQPULP3qcNhMZ5GfX5+XNDxM+jBUHiYex5KLMcxf0XRr4
boeMMzpvbLSTpgLn//wgjJ2p8Ba4ZSseM+K2/Sb/xLELBQrOxpCC50r9mY7ZWhrk
tWCM6hzx43SbSJJ1UTiRmnsMpl1VQ7RNNhJwG8/+mD1jfCelsoiSrci9fxQcBM0D
00pijYQbPOlH+sX1aA+t+QHMt1/8bgyqvkEBdzMG4+E0EmoIKVvZYCwzPARxqpaS
4Qs10yKRCt3fyK2NSY0e0tBED2wm930dSKpOZVrLRjYuwqZyJEbBc4wzY0ZZEjoA
VM5yLm8/jAuMeCnBeev1LFY66jNrpXU6TUy2cZe1wwHcJOKNrTKxssb9khhRQXpQ
UYfTgHC4ANzpsKVpVuZIkHOTyRt+iWGKxoAALx2aMm3qrRRfH9EEKIHwlcB3arfK
2Jl/pohLFXz19fPkLbUasVuFuyj+UqzvUjToJHBf7rfHkXW9g4vbyI/VjraPylSr
z9wIu8NJ9RXWURLtABYYvjn/LHuanc/TYkhE3SxrTJocd2Ys7d6wwhuGMGc16qMG
In1YHrvnkQTyT5SFAQAHLcpKlhL+oTRbfCuvhtsrkEjQHTfniFefujJDazBYNxEx
Gc5pD1xZQ93X/wrOKdct5fgdnIGqiqXKxx3MCY/ffKP9NuNwlKC1WgfYH53vScNj
1fVF9wrajYt0/7D5fdEDsT59NMGG0C7KphTL6UATB4G74eJmVLgZ02aAgdWM7PDP
c10EBrdpg8FnNlJbbrfSJQoDzLZ47xoPuhg+hTdJY2N3Ibe/FMgJL1DaVrNLVcAj
gRnVoRLaRwxhVaMmPQvPR9fucC4VQgnRfMFT8CcdA8Kygp9+RzLUkFLChe0uAlnP
eeDzpAH7MZyKAnQdRwI5iYmIKBnYneZXplvo+5BYVDC0VxbmVTy7FOazpcJIq7le
/cyGTOJf+IFmKwgjlWgkisPMdDQrJA38KVcCtO53IYt9okDUdbchyemUd+vTPJhx
PyrVevF0VgixxBLLWFO7eRcLH9PbmVheHrzqARipBPEUaM0nHPCnOU4mEy+jiXmr
wqgm05JG4Ad2eomrQsqIRA0Vg5B+zPZMktCxgPyHa66Ey9LlpC2F8Toc4ZtQxezL
x1VTh+OhvbSv/JMO9+btxerCftti/n3XRt3vRTwo7heLrAM8JJTrPNbQPkOewynQ
SD4O1fV1p5bjz6QrZk3Lbl4c+E5Htl/NrQSemaMtTkTiiOTUrQQWONmG/zHt4gpa
Aq+F8EVmhzXvDqgmpxFbayaiKp/Hj5DJ+tZ6YtyqpPbPpCDqmUpw4Nv2TmTfiGyz
r3Gf05jX0+L0q4iFhI4LzmPPcykFvZH0Kzp3U5qXiCb2hottmpXDDA+MG2EzzRMm
Isy+TreFIgcaAvyqa7cspXopbEgFCWVr5JmKTizR6H0NQWp7C+Pk+WWL2qm+QE/U
8Ggv76K/5F2XWcKX824eeSNLg/AK50wHEeWeZne5gZvfB7mHES369zTfByiIRb/f
suE+QyJEIr/PUUGPyKCdOb90cWiR0Zb2qYbPO1lFRiexGBR1iXUxG3rv0HDL0vKy
TejMUeXkyyiv1cL3cDnw9EcjPm5ENsl5GdwnqCEXuSFc6A84/flrqkNIx2LQWJU+
jnw3EbqknYJ82vz86dPWBJsn7/ni3giHUD04ZhJTWMslwDTe6aSSFfetTmbmCOmu
ccl0S9fn+EcoDh1JFj8nYfSm9zUUHlbCrrEjNlJPEm+ofvYucwiBMHzxSEDbeTHA
PaShWjbr+LPr9li3Rrty7946SJAonSOeSqs2KVEdA+dBwbzYHVLqRB1wF9+SFrFu
qCvoWqi3v2X4sEER/WT3wSn064+4mpeDq4TdLOgwSoEH1Ui6tZa8/2nDeViEESYg
sXww1mS3QzvfdqGGML25bRjHKWsW+aqJkry0cbeZ+rPnAJ7wCxwIBxLDdKWX4aBC
ny3tLc+AaJHaacDyvljloHcNm867E1LsyVk1n7JAp8SXkTHZVGTqyDWgKa9Hhr0z
2hIydNpOaTaGW28LUhcCSMPxyQtqTeHIGbDggkBCp+UHn/qcF28OMJzbeGnHBOvi
GbBYp/ev4xqvo+EcNxx4jymxMeLFDEsQiklZz32nXNKo0pIcrQLULDTmJtSb62id
ywkoe5RVId2Px8ad9i2Y6h3naOwCKE2mwJtkLzMB/sdj2D2202w+4ALCGy5zUXRf
6X8yxMi62AtfaD2VNc/nNtjcTfa5UHWRhJiiFVhcFwDTBW6mL3jTdOboRnMgXhW9
kxmA+UTwvbkAIixuahnqexi4znFNdGl0BzlkgbQqK8chGsvncRmACXILAs+E2hLd
TE+xwZiPBTY4qNoy/auaRkAqwtg4gRNuAwhIqS31UDzSjWpm5G27AHNXlagZwB/i
skGCwmhB57hnl0vscPZu6Tkrxh5GMsfLOEcUjFNTAekyplRLpHb3F9lBh9D9N5LX
VxvsA7KxKf4u9aonDykfunfWi+XXTjSdYI6JMhXZv7trpXuff0pnPCmteQTXwwUZ
3sYrG0wBLmdZp/xH9uYsrA/uuef12+ui3v/qkCqIv2Uk6ijusJmn0fk9rPa0IVa/
ZHtoUX/ROcTcxPxQAyhtbUA7DojNFCQsX/eH/S1KWA3C2fJzGKbRfZEoJD3TtMuN
MzjhXvy9OKdxyMukTyqk+LRqr5ZMdY9LPBVGQNEaOtAbb7xASfe/PkGOHcC/+LKD
rJ0ggtS+2rLU3Q7Whef9pt0cfvs9Fvou3nD+CMJseqnBWGo4rGLnNhozZbUYlcln
nNQsIrm4CZ8DOCyrXcy8vOEDd+DdjZOKYTg5nduyI42EOqf5ktShDdmMNdl4THwZ
fG8iaZ9gjTSAl0FHPjA3H7OyfJPw/Q22s8KSNnI3A90cKKdSr3LnGSt1500iGgl8
vwRwgmxmTJMTuONhCttKfNGSDezhTPXApkod7EaMoGLxX6VokRDGaQZQ3J+DExVi
d/T/frpL5gm84A1BcPwVHq01AZycz4+TZ3TfNFtApqS/28UgYuGSozgDTdm6rDC9
ypFGCA9xLd2t7tkZsxPZXvN96EQOSpCVYn1q4pnLJDhmb8gAUPwWjZ3CTvrTP+zi
hEb9eMiBod/nPe2DDL/DysBzbLedNTRXx8IZw03rcuVyZ6WwQ2JUAnXJSTOuR6JM
7Uc5v2nsqVjBTDF0LSZbLp6McVAyMBUxO4XRz4wIkdfvexhJBoZ7WwyN7omM2w2O
1TpZINVrP4rJy1bHv4U2RCQj16ZaD7TpEmEa+2kfyh9d7Z6euV1pURoU2i7OmC+k
f53BSSCkBulMRcaPOxsF7E1g1JpBmAlhJzK7zSVfEaeRO8xHYSRVj4y4alougCPF
IHcK7kTh4bbuwrPlt5iQ9lQp+AYNc+8RcUpOAIvmC7fRwQk4wpAkwsZyum394Wyl
4/M9OcNg3SPQA1+Pa91PUJsP/kSi2ZjLEGdxgvAya5N1bpXm/Mgn4I/zanhRY4Bp
VS2nNnmCGv9QQwkmN0q2uJFEaAmrfqXYjmXNM/nBRxVs6qmyDsh12kFrNz3NfCPf
jc7gAObRSqDscuTv+se2puJlFyCmQwNeLq5Xud9ex8JcpYCnvnDGlhUeGDBMxF0s
ZbHiwmqYqdGvfdhRQANEzGMNjh9hDmtK6nfQhLhAN80UYPj8WwnQEVRcxeeewL1I
k8tGYngLrm3uoauKefeIjFfFc/jrQ1sl6BHIzHmbwpFoQdTRZrhx0vERUaCtS5zH
uRT4HtfyQ717Ihizcs358+mfFYuyP4cCY3XwwlXylKkq16gTJVRGSBvrnM2Rsjxs
smutPAevbE0ScjiT60pA5sImEYNtEmFQYLXgybv33aguNToDMkFfPTBMsv9RT3M1
UMABarGhU0ORVg3548/EX57Ujx757/SJyvMCQqabwhD4y/c/QAxjRHzo35alL0vL
DJMUz+omzX56JdO3IGR2THB5jYU80bVC3vnRL+3KOUoucvIWLJF5rKe5Y1BtcPoO
StbOJoch1NJVSdG7HH9mksOXx8isYh8Y/WVxx/6eNioeM01oug2m+6d55L0wo+zi
C4XpLRnBAR0Ob/sGxgW4SoCDFkW9gLwT40j/0OcDR6KlwY4UYTsIXf3k3hdjuOul
cnfR3rOXtWY1bT/eTxlBcaoDsRRRw4QYKffjOQgDLMbjxKp8rKHkCKmhTRat1t2k
rBQfzpir4e2ho5gdR40MgKTzzm4UZNYVL8DUwNu+PQBUyh3kYIdwkjrQQ+fEXy8W
81UxgwjL44BeKKHvOuZkq9walZ3jNMgdKKGsx/FHYP52ReiIaZnmRoJ7lkLmLbho
cJWDv0DDgAOt3qJxUKUMpldnnN/RhVAX0lxqQ3iiwuwKooRQA8ZVEdrSuIqcYEmh
9N98BPtuTCiGBgE3KQHHzkfsSrYxdVmoBkPHQq6VeHA4npGQ4Vjdad1apLoVjSvD
2pmBMw76PJjXGv/bTGdmmVzD1C6KoecfdgKnCnpUxRKM8faT3D2pRtmaA7lXJsnE
Ly/Fq0W4fA0A7/csmiplfFFFHArBdhmJUuvYAHJAp0NiHE2AMhfEfADa13ucPmuo
teZ7nRJ8fwCkN6Doq5AjNKqqZKT6cLTfBG8pswGOmVeiVo3h18oRdH+A3TPlY8WQ
2xKoaEgvIboRkLElQAVkTxE7kE98vO1Zhp6QhVZ4jG00ONSpMuhIZht2Vlyc061g
r5mlpYpW4gGEjLj600KHbGh73btIR5AmkiaNiIcVqd737ZeC8jI68QtFqidSV4eC
gXOW0QKUtrcCMIVEnPeHHGb+AL+JIraQ0tmeFKlU4qZTMMVgCAgJ8iydKCTsjOQi
eg+qJzxcD2GSNu822sUhCWWepa/WlgyDKh2Q14PjtnxpwCCUBdlbXtsxG8++YOit
ZCTFz2Ab6xFCPd6vtlPdxXVC6df9K2TX6gW+nk4mff+A7MspEgP0z7NUS7/5C3qI
V7t8mW87J3XbSt/QzaaI/IFv0orQ75etC4ewQ2+72frdVEf2YrJB+YOZD5kMD0Cy
ItyvzDVcyjBIMYNdIPPnU8d4bdEULbgTCC97i+VxoYQ0XBKxoWGib8hSPjFS2AEJ
V+jMKcMV+JHimH7LC0sT7sZDrFmShFudDjoNAryutHqLHvQIMJas6sPt6YYc6gHB
6iQX2GS7tqt/NZglVeXO/DdyGPLVS4AjnDPQMQlMOBVtO9HxZIdi6AsM5kpBwsCx
Mfk6gNZOzvx29moFJW8+w+xXBpgsogEIUwHuqrU4Pj+HBsCs+UP06ZsC8i8W7gmg
hxnziZw0N1+Q7e9RM0HWCYP3qY0taIP4wlSwjxTJD8OH5PYhCy95FhNbMyLc68DF
JbTtdjURTAUwpC5lL4OnC+R9JDKz2Yx4/OmJ7/QG8uOSS0cNfHKWZct2lSuZMXMB
bL84XyFsS/ghZ2UzsKSrRiIFgQvW7lx/t3pIeDsJcLPYy1+n3eX1Hn/Sgx2mGhgk
+CGuK43JrGqqk3UTKHi/X6LT/EDEDaVhHH4YhTVK30y43YwlWA7qY5rSH3bNUiwK
tmXb/Ai8qYjuV1X6UTef+tWND9plbyz3bGEzxcJroXeP3G4eZBWm3o+eWH2R0fqt
ow2KOKdnkkIqVC3WNSDO5IIk3hYWw4JeirwafU02jzokve3j3Ect5D71dn0qSBBv
PCX7qWlUpKp004qinuSksFfwwamv8EQfuUNeDHFCQgagAooTUB9J2x1APmcLGf0T
0msgPH2N8fKG44BN6N14iaoR1E/el2SAEP1pfMjnOvcctQe6nT40t+cfMfTCAVOL
aMDWzXRRkf9wS6L/P4t7WXTVIUdgLxMLEhz0YQShIox61yMkcSi/pGY0jH1xzY6r
nyH+LkwJb0FH5reZZQ6+UQhWQHHUbyQl7JF9jKAFWSFuCcgWCA1qVIW4eSXS00zb
fo01I4A6LEY+q4vrvlghxbWmW5WuRXVKxYHBuRLgZVsgeajVAOeJGiCwk95D6ZcO
16kMR7FVTbdle5QXWmYtm+DdrsvxwPO1ffnAv9FR7tAHBCIawslotrsDDqv9xk40
uS52tmhizaidPF5+jDpugqnrX/Txm4Bz92aOeyqo+qL2dsTZdcvF423lpMJHWvaP
mDmCIgE2QZRkNhemLi9Xs6ygdUAIAeT824juqCnQJ3dzIJ5TuqjSxxC3exj2deVu
/TB7pSc68shhNFklvPuw2QjUbMzYnwChk/XB+XKPW2qkAofKG1Wp4ET69ckM31xR
AdyR9/EZCR+puOUFg4xzO/fATrza68aHQpTIO6g/Gm6KJWEuVQd+FIcZSCBKBNaX
kLW70GykUJHq717ADgnTD5NpFHKy7PM+Jpb+5Y5pnpzq64R7crEtac0CXO6b0ygT
+ZHk+8LNbXVdu0YI5ImmiuxsOTHeUMEIzxs317ij5j9TfCCSZrb8wiiWLR6DBBUT
vlN5Kl2s/i/SYXTGaZnkmCv0eAhChX+XwFpp/R3y/9/q1HR27OIYU46NEsmJ/1ZW
io1YVI5MP1RNb/jy/4uOZcELQPi9iarA3vDGX/4W0ujb2uzbTPN7B3k5qS9RjKcF
ifEFAUHb9RMrnc9PSAhXLdfDFF8/4PmHC/WsKC7OLvvwIAi5Cdvkg3k2ElIVj0Gz
311DL1fKZ1KifmlPz8p7T4DGKzEeAYcJFTpuUVVCf7nExQCEUCc+NC2jhX3pGuYY
VBlJ2QeKek+vzAB02+asubOM3ddBrog0cJBHp7hwTFEdFtyWolu/t6J8z91FlhFQ
6EltxL7PTq20tV6BPlPc1W/EoIJ7SsPGunDz7URGhBcAkJaq/TCxJ+btNXrSLKOn
+/prShCo7x8rCo0yAQQ/ndl23NkVvf6hCuEsYqLHnArWkTNzCVhGz84Qr5sQhXlj
ziTE7eURh/y0F9ZCR1CLZtMdym+s+Mq84MxQ6VsV0xl13WWHJnibVxm8AJF9/s4Z
sAKbRpCd/n/cEO0ytwFQB9MCM4dJ7z0VZkkQWCyYI8Yn9hwzhqYQJ1FyDNg4cXIt
EPD8S8Atb74ndQ1T/FM8I+lEadTZo/mKB4e79dbVfsHLjxFFYHdv0PeqSMjc0nqt
jvOBQ47WfBghg3SDr4aa9bx3b4EKbRTz0vmRFeop1ItWjQgSN0RYnc0BoHM0RmZt
68/AMel/LgUHEzbuhBmqCC1/AgtK8KQyC54DJrpUcHp3y+j8zfpcM/nhcJ8XF9VH
CWf++5lHk0pX/5q3o2oXM0S4GsvdxBgKz1ntMK7WLblLkNYVQqq4sDhjie1t50wL
YaudqjItaBQv9kle8OObX+VYk12IbZvNnlhvl5sbgQDX4/E6Dw2UW/RsoIspJRsV
AgV4OkYX1RAR3zbOD9Zui3mge3ivgp2SA+QTqvhHm97P9jWeW5xZhGp6BEAK7Np3
eeIN0LxYyfmcCP9dqq9n9ST8jvKPUdVIzagikiLkGeJ5EoHrL8CKWCSkxxGyq4bC
EQ2TX0YaDLIgT5hWSSq/rsU5Gs2vwV7zcCWOtUu0Gp7ORwsLF2pYrlBtjswpDDN7
z/g6B0FZ2+/6jR2jhcAiAyXmfm22Uz0q1SjjVuBFGoJ0ToQY6Ou7hIFbBwtPzQ5N
KQP7zE2QIhunBNKQIjd2s4gInxd4gZ8GGGMCsNKEB+Jq8yuOj3QXuTpbLDq20O4O
ixD1wn0dZh+Zqz8SIXPOXDoHQ8bafKY4lPjj461xi9G9ePMQlFjZZo9vAaJrEh3C
iDr7HC5V6l5KihXuizm4tBzWMK5TdtrrZI6dugDDByHUByzNYEB73W8k1W0WEZDw
e405OIUCLrZHuAiwkyhh8xO6ZencBhU0b8mmmWKmx+TTbGHPq1Id4BeTDSfd+5+t
xj/lkl/IrZnGrsn7SBfWrTR4NzYB2RsapR4be0knocEMa5a3yHjwRY5N63wqhuIE
xG14MwXjStHFFa+sbj/dOBPTOYVquqOEtcoKOWtiaUeHPYrXOgOjPWlD2gla+eA8
dS4Dhg0TC0Ytqs2mJ5YORMjwwPt9qUnW11/1Iptc5d24MtbFuDYqx1DByA0xrFab
XqJx9FHFM9nzz4Q70UjcNcx/5MmCWnG6bxWbuuXdQ8NvEtRZLJXyq4wZvyfHTgfW
1NJl54jNm6t0AisjzZBLgFZsfswgZx3CRMqv7ZWDKadLgT5dTHayJ7Sn21Y0YC/D
Rbz3rVO2+Ns+Ozftr9tfVoaDivaj+uqpazPdFoN3whb9MJ3xZU5HB5nBFPYOHCK+
MHMReLLImOvgFXmXGYLyDOsByQkfvLTyB2egMsuyg1ipnT89BjsCzLHRMBkxXu5f
Ef3zXm7NJ0o6oSrOPJjcIgQCqa0gKHJB7aiTXF/tcBq6aI/feqF4kP5vHdZdH5L0
VYgLlnke6CLXswcXSAWSx+6vOsyHfgVPgpxZC5gwPwFwEYBe9z66PiLgf5X99gyi
hx/nz2qB+Eh3oK0XKrxN1nOEqiYDK4qmndfxIfxChDiquEJI+ewscvDBWmSZ5XCU
3tquCbLEpqPuuuQjJvNtLa9Kf01crzKLKc5Kt9qQbHcLIc21WDbFiJhEaprTz4by
UMtMPBGJTT6Ki1gulXiHNamQgEqJRei5avS+nhZhIIEM3M0hzMRHDJTZkcSDK8Xx
Q8PSUA+66/Zo6DuXWGVNBooSZ9T502qBeCSAHglStkqsT9/JJwhFnHAzyCj3LeER
dPBNxLFwmh/6I6fxUcSj03I3oFF2LOOJOyLQpE66AT3M+L05Qhr/pxFJWQf+Z33n
1sStpsFFloc7BFf9uxezc4Ao+e61kMuqnIjKvykjV+dFId08eomEDb9zjyiopvZH
W9HNgW0kWgFd3CwSH83O7v6IUUrms89PpaNikemqYYYYpA6BUpHmlHMlBMUMt4N8
F3ooN6G3aj6p9IgJGpymDwBlx0x33zKx1HJnungUCwV36Ask1GrKigMo+DxT93m+
w1/ntvyGJQn7aJ6DxfHySmwVgwkHRas98ksNp1+qTDWumTdA7M1/xjs8qiPmIBfe
KiO6awltxQqm9Frl4VItGJUu/lLp998n2jz6Y3yQZPDWEFYzjXtsnNgvy4gRn7Aw
BAhs5FkEr+sEWolJ3Bm42Cl2s/VMv/GZMLNxyq6KrM+/D5C35i3W8rg2ZBKcubF1
tke7dZwdxtqbzfMpDmBlwutJEztXwHh05mMB8d+N0oOaO4ajclBkMY8H0z1ke7M6
GQF2GIvfSIRunfhzbOM9i9hCCTvD8JoJST+pvTkvz+pFvaNzXarrW83Z/+BqMNXH
RML46kZciLAy/6je8vpHetCfEg29FcGQvnyjBlEwBdWt21t5AltjA0iZG4OL7ns/
tZDg6l3R9hWopHUKV+zBUpUi6tMCPF3ezk/JddpC2U7LjIhrxVmlUwuGWcsh1OS4
Fu6+Tqcf4Lp/vfeOzZZfgia3LH6RgCLrScMRYzJfiTv+ZbGmAxscOcMFscgB+q/h
nfYe0VQY8xuFXIJlTrFdjolcfT1Gvo2kjc69CkNSNXDIFgJzU2t5LIMTUXnLHt42
ZUZurlm3bbdPsrfBvYfBYB8tME2/wQlyfNjsuXGXCkDuGN0kxbT0zath4eFmTnA+
0WRIPkf6MpP2pzL4ruRsHTcsPsjnwNp9V3RJJDE9uO4VLkksJ011Xc6PohHBw0yB
MLc+QnUkeFcuxYJYIEGrkD0EWTa8uzGxqCgYVMmGtQq5x5+WygNAW8qQnOBondh5
s3tbwexGB9qPlubT/eZISFouzmzoLpZON4iGnomRGdbOtH0jYCnVWATxCEFzNZTo
cgC65lXKSwIrX+3ZCw9vA5yBbb4n74S6yEsDUfKBP7JFMQJl41YAPJCsSJh6zW0Z
kUzn2uGM4ByF1x/fmYjoa15Wlv8DML7eXXbcCq/DG7Rby4WpiMdVNKBDemVzLKHP
S74kMwh6hmGUGhMbt8bUIbLIrcbYZ4j5Nv4ff7Iybb3T5zq55P9V4z6LC9p7pee4
gZ8Zb+RIWLcA2xRfXHNYzGZ06a7VhCJEEi2BmqFcopmpyKCGEB2+JCw64M42q4/0
a6BX5jq1U2Vr5yevc3qnKEIzmGnwDVTiJ1D/aLPeJdgfUzGwMmBq5pjHgTBH/AKx
J1xj7HodUMtid7n22blCZ9j2Ne0kMaMrPXjad6olxO5kwu4wxp4zDFcYcVo37KSG
y8f30IAWejWaLFMUKNo9o4/mlc6qxFnx658tXur0NPVib0uEpP60R5EK4kwO1g7a
SmlCN5witHgpufdv7JHXGToxJlXz2iFRhnKcMYB01gAARVCICdV4ugiAjS3sLlma
94yR0xxsz8vZ/T7scvkro+Oct01UXWZWIl30Rh39N5QhU6fiH59bY2RtyLKhVWuS
upln3jNvQ1+0ySP43CfPjTzuXfQX3D8KO0wgINTnB546HJ/stf56SNbYPXud8Kh9
mDSfvUasQ1RN9rT/WKV92H9ESUacPXweJGUHgCx0AoIim06eAGH9BgqGoZuhBkAL
mEIWa36lQFpK/ulXr46sfl3wFa3+1oEJBc4RDk8g+bAsIIZxWAKWWw8gsdsACH8L
MFftSerfEhmzyHu623yei1EzhlXwu7gE85eXAOEJCylQnEoGP7LA029GHSulbpWG
zr/+eKgqW6Y1Xky+gSdBkr8IE+wWeT7amiZXtciYqql0Km0CfAL2KsVbt3YOLXnk
Md6iofs7kWDBksNnJ5cPWYR61hioiu0H7LYrsWFoa+X+uxAFXqycl9huaaYyjOyy
gtjtfNLGxOtosRlz/TG4Nyr2Cq0Vsnft9bdfm2R/e+CrfJc+Tvu2cv1q1/1guTkF
ZHjdPhgmZ7aN77uQ8NI5leGjUMpCKVn9iMJt6puFm0+qlMNKET0rT3hyDAge/LXo
L/Vo5h6vaUAwPvEGRbj3qgAe9Mcisomi2p1uymGRouRS91oOt4wSZwodziMEZrMy
roXsBgi3aE/clmshrZ2wJR5NSy9OOJkNd37qXEIsuQRESh7QDVZhiy2MSzLYSSGW
1YOgGpZ1aT3nufhXfYf3kF6HkxQmnbxDn1aOWW28q1zVYq7PtXRJS0MKrbE9vzez
jFx62vrnxfrRkhinUrHiEO7uPQKJFOIqIAwgHm5K2IBtJIlKkoCMpg1zkmBacUp+
sGEGhdABHIfBQRlmAqMypZL3bNA+rPVKCQNRoZ9XQTvvDFpueTBQ0Ca54QoXQOF5
sVh/T6UzWWAILyEQHZxWZs3MjSBYlcYKgnAHCpsAI9gwtScHGRl4p1jrk4tOyzO0
jxHr8RrSe0L4eeLgJEAEsoV+lYEznFUVooYLddLTIUpwT68NB9urItDItO3XT8XO
OoldDRg1FVD5kDwfkuNx5jJhM5IdEE2QWAWido7XvwOnRQSLCGigLzy8cl+zWpV3
p8S63J8QmQZuKYjf/U9n6OVu6xVFIKFAYV/NcApqJpc/g1SUX0/Hr8Rh2euXx8Dt
/8yrCpEKsbf3O+Icvk7j7De/Tp6cg0Ws0UD6E3oTPgCJ8LSVnCcCmQLbEWubzI3W
CdbzCmTXUEkngCpCZHW/fRo01KL67thoWVhvImnL418Uhuzv2ABWWN9AUSaNfmCk
h8E3H0pG1x3xWr9edSIOOLFmKX4Bi5C0aP4IMh+C8FFhBxViQCA++0fMkpxXDcP1
57QgyYW4exAtgc1IQipz08N1q17awZHxxKfSkVkOFLJ1leP7qOzbag8v24pr2WYI
8dZ3m0dDgf7EW+UCeecNAREs8FPMLvnl0WxzsiKwWcZIT09NFkAYGFe6efo/yaWf
A6bXfPkQsyJKH4oHRWx2jMkxa3bX1PrPH+ewKD65o6IK6+DhyTaLSjbUIeg6pzbN
nJg3KntC1ddfP7mjcortxtPFEzBXm3m6/13MalalohrEayxHhbSPSFGpgexvifWk
sILeKPSqmwvo89h0uyZeRbF7GSp5zj5fu9c9EYFtO892z3Sv5ODRhyMy3FC8hJ0Y
449//QtWm8C8nAS7IqUu8leMCU7w9mhh9Th6RSzpVVTpPvEn+Fjuun0R4OuI5Qjw
6ySpUroBlnao5PIs+Cy2tfz6YTO26dJq2c9ikQyqFiZVAyhv0bi2pB1Sh2ApvTk1
k42zL25VzZ+4HtYP2+ZYFq4pfoY4CLB0/L12JthGNE4Tg1uxe3KaFznNF7MnWumq
BYrKuJcaqTyZTbd68qw9pcMTEH96gQMa5PLV3uSbgUCxJxO9qZncH8S4E0y1narx
ZR0mCGHSM0ZAvZDVTzNWdwvyfpgKw1eSRPlWHBRv809uRnl8v8ih9FRH+IecvkIS
6DeWXvpCDnCc53BiQeibcsSDxlG/N1p+NrUayOLtSa5SD+pbSo1xl3eUqs1n/W9z
EiSn9xB2e05p2pr51I3afKTfzLAWBEz47IZ6peROcoMyC5hLj7Tg8yTFIyh3MGsN
KjcCvynRD+BzJfPerY/H8P5D2uqvaU+Sp1njAIEc1ano0eXgCfRcLWAnRu6cMgbT
4DPJvJmTVT9jrswyL7wxpsBfn+uk0r0c7ybQW8X3owbBF1NFmcb0rfD3AjXpkua7
PoxYPJv35Pez/MR9G5dr0pHGdzoTJQK8b6yEEiZRT7CbAnfr4WEUih7taPS6etlH
cobeBvi9gHPXc0FbYW3mabCu51mLTpqBSi4rnhyrbFbCFsCox9L39p9rx+8YE1BE
QYMDu1MIfulgMIozY1ZNEOL73Pnlxir6J9B5cvqLo64OXvfKH5/wvvztgOIplPsm
dlpr/G8pCmOuoMtvWXOmUyGVHpBTbDPXW5zUI+/x21eIJafVTihft2aSlQZ6Z+s0
b3sdXsZNQcFVwZdOIkrU++IRftIKSPfQsFFnlnQ2GOeE3pGO0pz3uRAE+gjPsLuo
qjeYpXyPdBwbYkf3Qwb4Ksnu7SBy0UM8cSxPtPfjhqR/+eHjmSzoaUphLl8Pc080
+d0iqWYcAuXH6JtG+WmZz13VPLke28QnZloj5O+q6c1WDj58CJ9UDRjufYI2qiUe
6MXmVo+OXkKvwnVt7hMJjJfMN1hCzxGvzws04QF4UJHwinYE4MGaNuGmhxzfsqip
SzROTHzQJ/gd36UgV4ZZ87iaF3DRb6AD34SZoFQIAuo4ogvGuHisDOaSBT20St5a
8LQS5KqqSBe4szt8BSR7URxYDpKxB5ginScctYaPXdI1sHGl3GQShI9tvotlZBJD
fPHdurfYp6BrK4ScZc/+URgKDBzEUvJCKaziILtqQ+YlN09Kn7pQPxTNq3Nh6StS
xTOpLtK5QfhKM6U2FzredvgA7gFvDKqX8wsAnTFunkl9f8/5ZsG29lvSRuUm4bQf
BDlC9gElb/YdLRxUr8JwoCWG2aGeRd8iae6cdQNduPoS4a3ozZEwLIzAAcSO3yaw
2MxGjyepCsYK6025iVunFIdLH2Oy1cNEmvqvlgWZCQ1SZafVNT5y1DRKfhfBV/hW
bYR1g2RA9xMngGrnAB3o9SnzwI3nEy64324ATLdunwM0yonzbDOECDraJ7TjBBnF
6yBvoDLS5uQNAv/k9Bel3HoMUOQIwlrt+sMHYxxKhQahuGfNS8pahEMAVISOImuG
n2W7szq+aKgDUL3k/GTV4rGTjbEoKOzJeOrT5TqoepXNKlhjr2z9OkLbAvdOlb7X
q135clVsOqm4++Z06LDZJEwbA1fONv3DPG64H1+X+903Nsi63oMC0P92DJMx8ZJo
eevP3+BurWIoiEQhfGGJYZh+37hPfcu2ldKK2YTlcD3oDFPsSmLGd5zspWfkns18
8rLIjQCHBzvs5kgInWoFBwx+U11uBShJFv/F3SaeKRZFWOSJIscwfpkzZZGc/pmr
cwEG5N0NnPO+c5ZcWQtHajF546MliPEO0Hc3Socev1OWQZho+qkPC9nAaU+JXLg9
TQ9L6r+VEQZqeywLguMRByqHKuZWmVWq18TSNxiMqdjl8nubR/ndFTcyt7pwbIlW
S746PM6kwsOOqlCF+BdJMzgarQXFl0HXnbXvr3xfVNpygtysJCTjUm8soRmEaJXa
LOQXdTcAwDUNwM1/G4ozP95DPmrnXArTwp73XCZeuNXGxHuIq2HT64y73M9AV0fZ
fMeD8wbAPG0rFQMpm3mLj9bI0TxWtod04NzwUo9JgtbVP1f1j2PmkaUQP0QILLSy
p1wEZzkq0NVWZm4qFN0mjy1SpaoN9y4VqkOPdosyFIjQl1QkoZRp6evvJC8ipIDv
Jx47L5VwcbCSVWa9XzVvNXdsYNfc5LOqz9++eo2ybGdGGB+O6wjk9pKLW7se2y8I
PxzUyPtdFLGr4tyFb8LnjcbhXsm8esnJaOi10E0Ok8PEyWD9ej6T+4OHoRrEzNDa
2rEiUMIEg9GXVqNYVLhRRkF4genpzvTeePgiqMv/EJN8nDbBO9EReWUsle1uJhYL
yH2WFVSCyDKK9ya+q7wWeZ7ge3/zmuFvxwdhiOqXiSBUvnsMJGu/aNiyK4aNZTwJ
7C0CNBu2mvXCVfvi4QBZrPyGffRwzhxodYXXvpb3E7LW6zt5j4iTFgBWvt5x6vtp
/SJy7wtQ1Izv8c9qZf1NeYmqmftg6/UxGhuGtJa6YAVsbggUt0J2PeoUCaMa+wiF
eKwJk/ZW0SoaX8SQsdSTytiA8HOzTEnA8OdCQ9KM0EBP1WWG0xsEt5gO/HJvSj4Z
ciqOpSUyTDi9hD4z+KogsFCNjdg2EgyRzVKCtIViQwOVlMToQ9E2nok1VBEZvRra
DwaXWB94X7BoVdyjMuVCzDx5jxF1IydgfPsDgIwnAC9gN5qHBnGyGX+JRf34kGh5
D3bMxFpfkBslrDhh6dCPPz8RtGB0a8ryB3PU/WFOLTiDB8/5LN213gdQoabR362+
Z0us0tX+Ex10gf2qqa0muHvjUsWX3MwfxHz0QG1smv/s8cmtl0mWcofEMG9KJj91
ddl3jf4c4PlryUzA2lq4rbbxXiXinJTneM6mugYLYjxxVuIQF77vAGpNEFR/GRgA
3Ltbu4C7LL84WqbdrtJjHjWEi+D8xtRcI+QVGyX3olZQjwsgZfINEq7DG+n6uAFN
iCWLszct3cOGu08pv0Q9tmhCaLBxVfHwUEOYx5/GW8fTtTDPLlH4gLas3udC1ENl
O5kx+ATTGEm8Gswusd/NCZl+cMxoQF71zpS/VqDrLaEVFDXaCjFcEKD0wHej6Eou
Qr6IcCBYx9iGx9m/U3kULBLSSCvdzYf6vipWBPepbOmoHYE9VYELIKB3oVaLmuWf
/sypbuFnerftMwvYBpEqxOzHtaVCL2JLWNfqC9SLt4wnTzAgCJNjDk2YGI3x4E8e
QvBa1GaJWccxCbZOEiF8sbi6vFE9oDflEzhjkxhkdRjma2LM0i8kaUwqT5Y9BGhg
+ihEPliXILd+cpR+EJPOYHIhp/VwrDw3VBveQq0fPkECg+k9VuEqTJyf+MLySQmN
VZh58iZrsr6XjhREEQWMdYAowAGYPnYu8Ak0wQYRmklK3bEz8HpgZoO04LgjJy0I
iEobxAhqAdqgSVKdHrDZyRiXzdZvmAqYNS9daWTKw0o2+Cq+tibbaPocXpUw+H/0
/bbBfi/+3yjH1lhPJAOo0e73l0gi00+7nO63qhGeiTDqkTELvMdTS31OCtKQQtvV
/oAqx95umi8X4kgn8J/tUZcsQ2U2Cr89pgvRsyWetLIm9yTxWP/6bghGeSvViPv+
4pBhPBuivj2HwWT7hia/OEq5TTrrssh1VJUZ4rlWr25G2cAOhc0l81uRzEs++6SN
PdM+ps0b/cPirDezkHj1T5qu+yJ/UsBAzUYfsV9qNkM5o4XCJL1o8vOdWDlYUVsb
QKUOQiMgRMIuwQRGnkbrIiK7qP2JSyzT527lhKbUZvWhUGr4Aj3C2MIN6ePiYdCu
rhOOr04A8g9o4de66xiF2KBkhMJgHi0u6j//XVEE+9O3x++pt57xmqHGW1fq1GPo
RN2mG2d7ht36WJSFNa7dARGinTOYsGYkGSs8KOTUu6Z9tsS0qOIwBSgZw35mh9Zx
GA+0AyeHIK5AOFKTad/9jL3FLi/43keBpYjiJm/TL8hxemX0mE6y1DCWf7+USaSc
Xyprnch+nTlfnmNgCb1iLTbMDIr1W3Bv7t7J8lY3BQWVssJPjz1skhsoMfuMn+Of
1ws5fxlVQJW+2f9zp4npX5b5vTUOJmRDWrnc7evgay/C0bQtsVAcbfLlefoaPOiV
OD3dwuzSIrEcs9WFlFjxTU2RNPf1mt04CAyTFLI6mg5uFfn61/aX7Wcx1ZMEhMfl
TKRjw7UXgy/T+bWBGe+zZSQavE6IxCP9PD2a0N5LfweihbzYd8jt3ciNVomtch/v
CK1Draqx+ceUMuT48e01j4YAzI6Kyn14a6176I2jqOfDkJPSirK6zKrnH5uZXkDD
HJzhcU1sf9rob10KsFdXWS24Qy+BswKDdX3LFWXXiBrl+/LtUzCCorsyEBsn0jK5
x1vsb4G11lJurKYYm0Z01btmmcMWFzIaTLphQvFWvqMT3VRBq1Gn2Uii4iKcJjUu
uDNll/rwHzb7aZWnfExL9fIOAEHgLFBWtOW+WLy3gWaMJUdFjv3s6eaDAavFahwC
+g1q3LWk2pqTjnfD/jM38AH5kbWAogj0NegZAthNETjp2UB13T03xvRcYw3whrCY
TN+KBCnf4raEnMaYrmhDCXbwCKMRNsWhForr4ROq+Cg/aAmWH3evJ8HeVNGSfiXu
OHzO0NwttRIIBrTjMsaaQNh6b+Kp5u4BATa6Z5DDyzHnUP/gXJR7SOUp0J17H3/+
YDI4VVlN5A3shTJHoz1pAVEfh3KAQzztmA9P0+7EIqWGaHledTtU5WvbT3qamhRg
XX0kl/fgOkQwjpEOPPBNpGkEf1vhJGz/iFU966Yv46vZqpqWM+03j2fQB8addvO9
s1VVGmE/YAmqNn4/dnH1osMktbSvUXVl3MQlMCb8hFnSTSYz8bO9bxSI+daNppct
ho9FOUubb7Kd+DJD8IY9Xud9mOLv54f+U8480qsAkVI6B0hRA29ba1vNf0DSYQ+U
fujB24cCaiZOhiiA2MNiu+ZWsp7/FlqGOWD4Bfa17GUMJOHZ6oB6Kb0SNPh+N5gW
OKCPBfzJ26zM5VMf+hvm6vqsnfRLX5IfXt/+fmbTydMv5KjfAJZgSysaBmfFrUhu
FSPyzIM7c2FIAWvklMYy+rKF8ppII+dgsh9+MDPOHDhFFnz/B7lBxMbW3A6FIch8
zdz4y8DO4Q4TW9SoS4N1uueWHfnrykZGdLxXt3YdJrvqt/YRHXv8JmGAdIoRqnjr
H1I6f596KKwatRjfFs2Gu1hZGP5gx1ajPloM6Q65zKutoXPyhN5CrRxSHtIWpLst
KA6DNv47nb+OeJxFqR3ktdrRA4GHVqDVZPNt0q242mG6elcd4z1+gAomzTnG3hDo
IBNMsR/s2FvzRSQFmlvnDiZs9otOJIEjw3yH0x1EBMbeMkYicenlr/gpPB4+ml9I
+8dAEqCnN3D0kpeQZ9wHbSuDI/7tN7QZ+4QS+b8jEApdvxcJ+1Oqgb1wcvnnLndb
+DrU21N5VaP+j6hDxOpCcOUtrijeUp69Cli1qvcbMyFbNlVPM22yVKZDn1z7D5z/
Fym18wZlBQmrfmV6mDlsvmdnh12elWrQ2fdZxmDx+nOg4Rr+WJfzF4bX+woUQNlF
gSLyJutHTnjoJXA9xwwRBkTxQQRicOOs0SbidEm3R3tGEuVyoHYlvry660qdMNSG
IW8eDQsJ7q7kVNB68D3ts15lWnE601NPcNGEHP8SOXjr7oBav8JQ3U14vMwWJyUQ
XNF3UtWB6qKAD1wbWsHpACI91Z7XboLa8Ctdy2NvCsJrjBVU4ieVtRorplHHOUad
wAoxqg8cYGoklpLwjxems2ZLzJZD8hf8CirP4j+i0vVg3jCKdp+c2KMnhCaNcnqs
cf3yvabNmCEXN9o3kNMh8FzpddN/JnFsppKUB+TXAeLq4dsYowykoxGvFZ5uyy5I
CJa2+4c5BFxuhqaBQVJHfxxQg99GzvPSPC6FFTec7WJUYz1Qo4Vn+ufU/9ngPJ2+
uof3qZajV2yXcIa0Xo98y6J1tFqXi2XBoLrYVSC6MBiIVN7E3s1TkkWsJZmbCPFW
aC/BiY2f6EM4c1KS2TkFo6MuNmUjfR+DN1iQy2AXDWfasV5cs0zeWPsL0kADjZFJ
O4AxIh3KlpyJPRYDc+pSjqHrUJYQDbq7M1BsUCHiodVSs9QgAFS6ZpoH96Bs97Xf
QLA+bYJC4ZTqGcwgraGVvBt63W47fgvX8WNMZM7hbk3h7XaVYVN3pK13E2F5zfhK
aJ9ubjeQZqgdMumrpHeHX3V6iAzSzpU164R/8qkqEBNTjl0+RSrnXVgyAsJjK2iY
1HE95AoEK0bSClXuQ3Y3X9zvitBQ4uhS0Xjuh2G4bWUKVXEJtlcX3M/Rlpvykybl
wEK8kGUmUeSlSfW+9DgKa95K8DKHZx5YDnEB7v9zr5mBPjOEeTkaoh21l20+QYkb
yWfTHmFzyOGr/T8vPhPTKZ4ONf0eNWFwRAvbE3jxiOR9MQnwsHJycqAyDOZDpbgq
BkUH4FzCYR2X7smL3GYeeFLtckQptMXkIY9v+qcXwsa+aTzdONBrwV4ztQ/eYKxP
B1+wV4OtOWbWe+0AMpCrTy5U+S5jeGqPyxpDrBJHDSuX11ui7a0qM+5FoChyvd3u
ZIjK4ypLdIpXTYePfGL+PFdiYJI4LHitiX9ES6haFEPphCgivJpmM54OkSBKEXis
9UimjYvlxylJjAbLtvKnRbOyT9OULhT0CstTWt4wLbqyg2JU1I/8KjpOgMyKfrG+
kglQLrmrI7m3X0D7j0cE6cnEWlFGPF/Nhe2+iJbDTXyzNF/KROhehIxx06KFI9g7
lPkW+zGjIGB1fb3NVL7DfdkEqe9PZdniovbvv3h6+KacZVxhApcWxR8h82LR1OmO
bOhyorn81zSHch50ejO2i0queRj1DYo+YSHz5MEuGXucxHHuBypUjnV532sjAXO0
NVELetRr+zCXDiqyg7r6R7+C8iSvqrLNKaNna2eeqNS2eSFQCrnIEA2yDR2wfrGp
N4Otj0uUSoTvLNEe/ZEZtrFeN4mBtGfLMc7NF+FRABS1BCzbvTbThPkCN783IzmO
xjzEHnp+B4iUTVjYmRGL2bTsWAKLPvo/iksPDAu1eps5k5SOED1Z3skbN+wtXPGg
MrZNk1uTXMD8FCKUQuJCkseIo3ek4/9U5PKZuM00DhDt59jYrAtr8jlnxdAhRhsl
/oLCBA5Hc7Y3nZfmcA/gRcX+nJdeKNaL30H0rf3/YEHibQM76unq/sSZZMJZbdOm
LTcLKUXVSoy7coNAwi3mOJ74xCAqIYxS0voglLXhm8ZJmHPjGOwuDCtksqCjvP6n
3W5IPRlcsuAZcUZNLb3OvGIqS+WBYN6SrVWv4M4avZ3s76sHZeYX9lKYkN4Yr23s
i2qG+VLbM+jsi42qRV5wCZnTcF8W6XOZ/tTyu1/ulNlJffy1+vjWFokmqkyx1X9w
FyEpnAdNJuF3RLa25iQpIvgrvGJ3igYGoKcDqgvhDFZlukxuiJFRHmwNPrVN8A3X
N7Ea8Ly4N6W1vIkpTSgukOzBeoo9PVRtQNxtxezZYyboFixOq11nwLoWS0f0v0da
MmS1NZZvReiy7wx+rrg+BLI300H1kWnUArzcpDdye9OuLziJqgxn5HJXFf6zukUP
yWTLCwTqO2QBZDiOCiqM8ZJ04km41MSQ1UE0gDaNmodGzNYgWhWnxypdb6rUy1L6
vbMAu+8jp2GwdfPoON9Z9nTgBaCieMG7pgUZWIGFRnaO8qwPAZaj3mADYr96/jEw
cKknDO/jGdb6XTnRn9Af/66ju5v6+v8JUhhc5jjKMYYGeHVpfLEsXHPeN2CN3A2a
DfFfOAf6F9uL0bpsJnOFq2bkL+BWm64NITHrTCn8cMuC70QBauf5gQnTitBI37XJ
xjmvNbymP7w5viODC9ItDV/JHr4bWIWInlmOdY653ZXLM55YJCCFNWH4EQdi4IML
5elRShqOg3WTzxyoApAPBEdaLCnr6mMt58ZLkqY8QVvXuwySi1UpyqArMCiE7X7c
5pJGifV9Hb1ETaQtA1Y6LiuEFhISsyJo/UyONoYIZYTryr9AZyW/m8LiFz3gn7Hk
SCnJfua+PbZ4MRoyL/Wu4COE8Kl4L377j/+5VRDZzK3ekVgHC7O5F/yLFXipCqNp
5IUTIDnSc8mmkT1VIrTWfIRf5QCiE94GlLymLMWtxzkAOu9aWHsi/aSAPPnJV4e1
WEbYR90h8Q8I0NNt1BpWQSqZTfp4SZviWOfaMiltN08PEiVJcFU2qNoeCShiiCim
4Zs8T6ajKdugYB4EcyjsX8XOLtiw/deCCdVvpd9s8XN76V0Bjg3tSnTPgRdLpZag
i5ZjL8jRlcRMmdrZL41heHs9xM7ut8A+l8M+V1mfqhy8WMnTGLCXkLQg5pe20rJo
kaSEW7AGA7yocL1s17aoPGPJEvkLAZxzzBcrsRgd0neCzka0CmIVOi/HrvHFqCvn
kkc+mvZWdGcDSjz2x3Gfesixmj4gj29LGohGtIXNFflSWxuYWON5I0fZz0NSHOPh
Zqdkr+FVwgvJ5HDJ3HUwsB0MhgJAGlHTKQr97p2V4GWYQsNyVVb6YEhCEJe/TEco
ChaqmfTAxwB2cFSfgyro8ebZTMfqOZFpYFF/F6LGPWLELa624JPs26glGdE/KEpL
1AcEBz/aGNh5rs/2KPS8vyExrmQKhQtuQmn/H/r7vpJ6QknRJ2u6to0yKUAfiiMy
7lndoA1Dq8LzZj7a9r8TwM6rxbmnd+qg9Ojs9/cKFuu0QOf57RrKTj4L71QNJ/vX
eZZvudRQBm3ogPghyM6/AUEINiihlRRfjH6DMaXQJwxeTxV4vcrCzZ5ZqXH2qsfR
vI4xJb30BYvvJBNvfWjNls+BitIc1CxSlt8VylS/rxTTQzMHGKktnOlxn9YGqVre
vtfAmdoIAqx67ne+Jm8X1yRdtQLQF9nQuIx4ybjMHiZdRiCt/NssnFIQRrUBFBlv
PBgUNTjG+16H/CjCeimq16Ajs687J+9qZRUq7qVfTrqvx7OLzPYV0ZuY7KxQIawV
OUKg4BlGk3eM2Ti3oN7QQzKKATPN5zuK+zltoqlt2bJ8DCdbIc5OnaD5saYjMAcP
/XWSw5i8HByY7ka0f9TyHSIZDorTothEff6bBbgpR5R2tnP/eTA4aBvW4VUSeZdS
5oEeVQ8rEo+AyUUbh4NTvj9oXKrCCLtZdq0BnNb5XMmhAXmQb/tj/MzgMrASZd5W
jA8Na2NXllNHSMKlgCw6Gq0tIliInaA6mbQNiCQmO1xRHBZAe9YJoMX8ywXcME30
Sf1++2ts0qI+x8TfvNq7OrXDpJJicw6Goe3sRbug/QOWhmwX4SzJhTgKl9OxjSu6
TaNXgWtJObemhcoZJTaAyw3SkdUBe8OQnMwXLyaD0RAhEml2nxZXes/WTbqlAGdO
qnSZhPnGFx1MTRhKrRoT7yhDPmF4aEKLg4m2ADyMjWuCqku3Dgv1TJkpuMmmhryz
S3qQWqJfCa7ju+eo0V2XxlGOoYgsLbFH5ZzNrQgRB6TjklW0hG40kJn+sH2Tm3Nv
HpRrm+9Kdig2JWzVReDZ6GXi+v4W4hULxEUtzgl3mjrYAKARc/8H8W0xFO+Amxu+
AWhxn7d7ez6Ze+F6UELb84Krp4dYK8SwoVnkS5nuF6RvIIH7gr0qnLvqRUmUyJ0y
9hjRBYVEudNhCIXenjglRtAHVJMIoAE+hwY7XNjesvJ/4q0XspPAU43dSEySDD8+
0borpE4/yo8lgMivz+A9Oy1CkqVizF6nURdBfdVb+PbU3cc+4RYO0Iyj68GiEuMe
asNb3U2Dfi+Hcdom2T2NB+lUNt/U8DZOYNi0v2ucsPTGazyTQfwD6M3SOuiPdANy
PEn4ekK541jHOnw1zDENJ1dWl78AwyNwQx5f5J2yAHpXjJgXLhfHRL+Ndf62TGv8
QOrV1bGJLO9r0ijvmaggP2Qsn+hwUO9P0ofPCbHwSQ0XUPvnmopi0MP86OCqOMaM
mT+WzFG1BYbWCPQu+xh7gVJaHExfi9yyd4ZOKGl8ReSeefJfDwNphyyMxrjhcyrR
5dZB2ChrLgQax2Kk3In5ID+5EtI9sWx2JnyVvE9Gq1IrrsTLxbqm7inYP8KgXOJK
9DGa1fqJYDCrnTnOzgePZlhUJiS+vTxiK11SBu+punMmJBKGXs7lJnm2ZMNeQKSC
/h0BQZ19JB3sakjGMm+y7rrEXfdD03NjyktWx8eum+9RE0+LkPwXRB/X9R19oaR1
vPcg7rtjlnmlI/Q84Bkwyc1kIeMio5O2e+6HuXY3daM3QTRYFCD7D+zQ0IAJPjX0
/+tfmDhrLFpGR6/HwASWeW6Vd4GoJXYid3wxKFqexXV46/IxCdDdD2hLMtfogeqs
2O10pItljxUV39FrcqCQwUJDaE3eHtg8zEpe6n9s/Ge1coninTj9pALGruunOXcS
pd1zJEQPbrfJkhULWvzdc5kW9GmbB0lVRPl020HBOzUVtu1q/H+zYVXXhsJ6kGdN
TIgS+ubCQ7uLnQPl79M/UxyTcNDIL9ZRIUMGhS26557oUH2ln4ZxBDSyER77e7Dp
iSi+xFQEb67HZEtH6qkpgQmKeS1v6eim92IQrg9YJxVZ8DBcPPx9CWK+Lf5jxR4h
LOzQJHmzrO3gS9Z+OEFxPjYd1MRyVyY5yba3Z11so3Km8A+rLDYLJwekxGy7Wlxa
NfqUMwNzYOBJbZtRDcLpkesq69zIdBxgfBH3XKBn9iL0kER6hdF+53+aVZFDR9f2
ZUfv7A7wlMBxtjcSr+F/rnHiP7oW/sixX+TBd6V5xfGOPK6AkNJScp9//k5ik2WZ
7amNdE7vjcYI8Wxtprzu7pupB+SYLgkq9ZXiLs5c+jT2Hbaug8RFj3s6lJTYDLl0
bQEfigy8ngFlm0POgFwF6FLxGtHRBX8gKV6zzc+TWulStfKW7AeaY+lQuPduF1Dc
YZ64fOugRSEAXZ7MobaooPk897gG0ZU88ussqdflfuVacJew+KuQjG7gaDKxA22Y
1tYELrGid7ragZMCwGnWPvqK2XC4sv9Lp5zkw3yz2B9vp1v9ueZ+0N+/nwVU3Nov
gOiRdgNVJhLIq3TaIM8vZcTNMz2fjsqw58/woyLOsTSXGb9omfnzHJkNj/4lh8Jl
oBvRutKk2QecbxVksOt55s5nmu0OQG8cgP02KnjThn+AwuJRjgbAPB43UqlNFT0Z
B79tHYIK3FYO57dG+T2nQH2KxabmEqOF10ByOIlvhZ6dMm5X0K2JU9L96MfI356p
oNlfRhGH7UaD162s7H/kn4yERq18h8yRnlt/GkKOpFw7kQtzJS2XGgDN0DC1sUdt
RsV7iyNBpH29PrTkfx5bw77mQXxvR0PsOBtuvOtF5s3iMKLlv4G4VH29NdHgKtxo
z/oEAm4YbQx+p/d7RfDa3zOa5BM/mpRlLY235we4tm2ah2Njm5gJmvJ4v9kdnxe/
9wzeTn8tDFUZitL3q/E8jEIOsr/w/LAi0uMIC4NHXIG/8WfCtmkXBqoCNE15GQlZ
+FMs3pRqHMbA084ff6SMOy4nkSwWlsqq8YjCQ0J/mCBXYc7ba7vGtWjQlSqk+zVY
Jnlozocziet3fSS9CpCsp1cixTP3O2XtjOVZ+XJO1OxXE4YooLtA0L4guE2iMNaT
dQDgT7L4TfidcRM0I+sqq5o3LPrvz4mtaohm7QMxZ4ReQo0pnODuTbP0+MeebWIv
qh7GmbmwY3wkpM+7rECrZutlQfAce0Gct/AU6ASCh8MPZ5qb9QvzhmhGnAtJSr4Z
LZd0rcUT2XFQhLKZQzQky715BEwkVeCwK7u0UDDdSofI0Yx176PKh/KgJimpvceB
pYO0E48Mt6MlwfslakQCxn3Eh3GVlMYvb+mUoq2wOfKCFbJ4n8HbWEWaNIGH6rmK
4ht4Vp+uENhwATzEWNqjaHRDKnFAglWAFb+lk/NUV/+NJbiqf97Ek/Zet76HgWqM
LRRx5TNU3OhrJ0Fo3Db8jaEq99LhQGaeJDwgpCyvVUn5W3Yr+NvoYMkejWv/y1xx
GVQWPvQ+M8aKKgAhmtTbdeeUHEr+EUxJp+o2GtktR8RTgcQP7WSqYP0xyIpPK2Cs
R3ppODm3N0paWmJvhfBzPaBuaVdKSJB5hOwPNhBrwdsd6q47E4jwTzA2H3bPg39x
EqU0cKcycADO1TBzWW0XaKKanKrx61lTzF37sMaZUYtwzwvbWU1mJLWVA/VdgFP8
EiDlolhbxMIgaG+pnqNSiZOK25vnwxtvWzJeWaZuKx6jQxW1JRVyh1bJ4yUYzcak
omcAweDF8PAikDd/LoBDhzNcqY1gN7fGri5BMZgEAUYvtUQirBqy5D9a7YxkWCvK
PHSvlsVvteKOK1uIrxbxCPhn/nqyNDA6zHl80hoP5I3Gqa0b7VrlJmHXKup76xGG
h7RBPmVTCZ6kLBVhD6ICliKBlKG8UZpxfbEuOCHKOSLol2f3IHc0oXmH2+I6gk4T
7uVTlbLmgSUGKVwLM/RCULQcby/1PaYkXjKvp7H1rlSgd+V0mrgnuMfWTFPnlfq3
EVE1ScBoh0bpS9TnOxbc9BcA+Ar4koCV/YLaviNjuVYJ85hf3UBDQ4zkukzbez1C
pyMrQxnbrkTBj6Y/nDouWbRh+6oq+Dmd55Nqio872K8Gzf3s6TNF3wJWkwGseUmj
a4FL7uZtlcYmqzbNrkEJ9RbiPwV0B4lwQd8cf7OM2i1W68ePhSJQ/XZqO0E2a1Jl
UPXli1OIeX2bIQjPhA7hPLe3124HWlZoGnmHy1qmp52pZfM0PVgGzOKZIU0+JiNu
Ch+Mj6tTI2/WaavAEj35MZLOxwtSMw2+E05fpqTghQhcUkdAcAuIvmXtsURCz40G
05TyGKQmCebxdwzizUM/PQJcqa9GGKbkpOVXGjpIowCjwyf345jucs0embkpOKan
MdVEf420w5MlUF/8AiiJ4yH2Rh4UarHTQD4wkhz/JMYKV2p7qkzHNs15ujdKRJ9m
jELnANUxVNMTYAdxL83nFZkY+dDzsq+RfzJUsFTscJVaQ85xxmVmeh/yb8ppbXRm
XQx3cvhmtGOwPIZYaOkalP8fXkkZAHaFPQ3h6JYZAKhUjrrjCiyB4Td4N0NEIjUT
E/ZYJrXJAFYgXgo+ky1jdmGV4ggFkT/+EfxGYutyqB4vlRn1E97Sa2cO8FMT55M5
NBilYr07Pu3eUQdJ8b03nKfkgaOGgxXYMSlZCz98EOC5Hq5mdI2AyaYjfdlGD52n
EJWg2jCAx+SCjJLZ6GIFcvvxDexNsVGO5sa00Hotq4e/cKue0WeTeJWYGRjmetVQ
2qH8dNtEP+b0hHq6n0ww4aDnnA/RjJsUfYFk8G6DrgLLaqrxFxr2gNV47opOuVQa
Ed5s2KJI0TctvHJTfSo9WflvEyWoL8QXo4I/kuhWPFEXFpyxAX1fjzFnrVQ4uj8J
q4LpnTYar6ROZSHrJPWqcCK0d73DyR+y8mm1e+A57VoGGj8YaDn66FnQly/J6/Tp
wXwuIHLpapY8t5Rl4TV+ZE4LERKojxJQ4GB0rXyMQdU5sec7epDCr4gQlazqewjZ
TqeVE2nL83Kcw6KThn7CWZycD4PFHW0YzxFq5WGwCbHEDeauvTQgZUmSYXd+ghgt
rlLaqVYlIQGR5r+5BUmDrWNKM/VunY7rTnMvrsBwhPBE+Vrc5y08/d3qq8UFhN6Z
A+7qmt8SLn0PN6MDMlsB5HzkVQhSco0Z5/KPVi5zwkA2jnHcn9a6sBg0U4Pc2gC3
lodkPQdjpb/lcvyVPUjzuDRzdLHlToxX/PHI+zVbRGm86N4g9zzst33Uq2WyEffG
2sHd6qZoNV4VxM9pKP3v/HVJLsOMUhd4m4cTI2dMttQxuz5QVJfal5KPMbcGOyiN
LQdio077igPQL1VHH5b9eN+e2c1N1Sy4Aw+Q6/WxEBfvWzj3wBItViRP1gigtvda
Rak0ToaR0fJQcGKr1SLoq8XIwYLbmYywszXOEw8aKIs03O+dHeaGNlS50yDAuaD0
9T6nnY7MbrTj4myjnp5AboBhPgnlVDkHGtHhIiMjJm5XIwIHgVgRCBgwLI1moppm
pz3rG4bQFKwJbkbmNGJqXY+XIbqrweJYbWrHFA75sy3ygPm4NpfVfZzzGqMkxgin
y9lDiFK9B6MbL3DbFo1EhbxoYyQ+rdYLR7xiIVca7v/L31yJ6JHOqDCQ3/DFLZL4
wDHeCZo4HPcBWc7wxNnouVRzPnU0fvKI2cAOq4gKUMtsXifqW+AYsfIcWNH4XF0S
xfbs45ADXvUB5UMZKGw4QOyPtybdZ0XxvVqU8ZhQThJah7JWF1MFk37hpbE5HKqx
kesE5eAVO0ZGw3cIrmiAICwMEMWgbNJljWj3jATl687/suuD0A0oewWR/bzRkZLs
Xnu+d7Wklf80ULgmpXIsmsmDm9t3RedLq2d2a6t/CLjyd6xE/ICqmrj2bO6aOSlS
7H/kHR3MuaTbbEyJ6wX+y4jdivZdE8WDdI5H5pvbAl03T/ORiNuxjf1mONIAtvmo
sKQ81zXW2gDfBAmN37qoyvLW6MXesu3ZbeFEcHhV+s/j20Sq0y+uy44AnIAmnNDe
KhzxcQ9NT4kMydjL2tny6JTLTX6uEWeiWPNXQ93IZgPS+CKENsck+HAvyUySm+g6
MksIhuLJ7+aMvd+iDv6IpcCfCFfA6CDy3Mt83c0HmIgdlZ5YOZ1HhPkgYLLi2o1M
oh0mKu+da+qnTZgJupmga/vvhTNB4QxjxlkvDvdc1aWGxA2dMRI0LpNdXzC1ensp
iGVyh7hkm1E42uUVaRdRSQiRNwHfpVldKMAahNjJy56nfVSgJkEuXODjvcb3LIeg
9kvOnlAcxBBWWl+d3Fjlwf80vMafBtGqJe/SvPAROXl85yJEB/4jTWyhsfVNVFDl
6rVuFnk+QUefby1Bf7HGxeD+XiXatiLCuFKtGfG4hAeWCTILVqdcBtgyEXtId0rl
GaAvbsvklM5iH1WF6zZAohIfMo0FZovO/7xuvCPd4QH3F6qIa6TdJOyXfgK6/vn8
BIV88GsJphjKsX29VsBbZVRBCBqgd3ArS6lX77SAsIia+3X7E4LuF+uERz3qJwpw
VqSPDtN9uHiyLESrtgiLTfk/HOVb7+4O1U4FvPlamyiL54Bj9Lc5YQccF7D/tw7F
wf0PQX64fOkaKWure0BIsEXNaA8q+XwxOdWXmCb+yl4sin51yFfZcaBnz8Iy21ID
RgWfkm0yEyqmuYmCs+5xcM4wRnzZVr3eX4DBPAOVRI3WfILgukg9kXySsyvCYBBW
g6dSsYQ8MUnYZql7dYR5ZuT5XgMwm4RCxUFupx8PO+rXDmbg5fwK5gkz1jFTxqL2
GG0DGl7uFbAEkdjRctwfPQEysgoCveSmZwil+Idlt8fD/C0WHlzO5wo609hEcefs
ASFyQQn6Qj7cvOrudON5O0XtXk1hlHdtqUpH7OGpLN1ALhxIT0EDYDDSjcx+leVU
rgcr5+2wArBrBl6CvHujHFjTaRKycVyjYjj75SC7Vlfj6Pqytq4V+MqLHAwfWisQ
u5UEo88yY0XtcA3dDm4oHzAoPka7yq4n683qjUzkf1U5mctTrV5cInVaLLuw/MNZ
sAl5rF+3iYP0ouiYL96bZqbVUfs3RBUbdxJ4Qkd+2DIk8Wso5I1NGaBAo9Z+6EhK
KGeHbOn7yMl3FmjMZwdQnHhnUEqCr7mBX57kEObwcaCtJZbBAqhXmn33rcPJibMv
v1aZNDTzAO/36Nki7YzIKmgU32xdlE4Bs31GnA36KKu9ypkQ2F5dLrJEk8zrqYZw
2MLKTOL4gHONI4GF3R5dJI+PVKs0hB8LYGGqrWPRWessmbCZXlPAjM467WPNu/SY
EjuS+P8OiRISYl3E68PpgVYmwGDwJoxsfFc+lCI0OTF+Pbafae2cZ7tYp077/FOn
+0P8/2DKc8KuHr9ovfHOvyZda6cRxNBQyFhH1elo6uyU1VAhFtDXuCQNPFJfoM4M
oOTnp7ReC3q81GByLhhzKDdaR+fcp9cRnLs7C82QUjaoAuv6m+hE//byuwlxGN59
osxsfWMi8wclyS3QVrrPibGKYIMujkL8LMylSLiA69KNcu4+6pL+ne5Vco8T+H+C
yLcCtvaeoK1azXysCyEKM88g+LId4J7uKuNExaTDTXxmijPVsIaNMXoiH/CY3tz6
n6pUhF8BNgPkOj4npWs8BVctYJW5NdjgdF4maRABhaNdfTiU28JoMWWw+YdIWuxz
OZQFyCJFhnxhdWIguVvNP1S/QWDIlo3xHDIpdUEJrG0OgjhacuNRob0NxLqn7Tkx
0POKERlQXEYflPRYfBFvJI2a2TF3gpp7+pd1XgfYxxWAafVlJnGXw2r6WyGdNxiG
zGptgRdgQTab36ulrPNkJytLLLavMLu4MrfE0Yz7UhDEDCY6sCBVUw3aVX/iACz9
JF2IRC8H4R+bh6sQe9ulSI+yXv3XlqrYTK1j3C1Fnaq8rL+zL8HjJDxF4oZ2fL9m
mGjWvGADWheJo2gwHHFA1iQ313Dn5kIXCOOUAnow6L4nFEjfLd0JG4spPsXAPP5k
ySwCgjMUBfc2pETyWZJNmRvsrV93o+t3hMQBQZge8jzewrXcEeRL0zDwPO9st537
1Q0VbsafRwkiM73rJqY79BY9jQa55hrIz0FoZ356nNx75bozAF0clOBQRiNqUgEw
cW+/wWm/wnRDoHQ/phoRRcbLC6NEs8M/eqq2CGDVHLtt2Fpx0ABnsJpeyVW8FSLn
e9V9nXiOsL/zVpOI2ktkdHa8RPF6LrTGjDs92U+fQUuYAKl07NY3zjXNr3TZoKpa
DeY0kvOhzEE/a577zCmZZoIfBhvZrnAuFRvrN5D9f/4esCzILNQLbT5K+xh6Z82R
lykysgH2ZfpPxERs9xWy0H0f3Rv2RCPsgFfuGZ194az4KNAMkNJuuHeUFAWYmMLa
LHRaHPFTuJfZYmiTCeN348i0boDwCBRMnKRtumj4m2CqmOqE6Xdld10z8D6uugbt
HfSY4FAzQm6CtT+Win4IXOxz6Ea0lYxJYId3BVLnwct02yYB0TQcCp15cxhsCf6T
u/HpTKugFBGZuwxTLYjdX/0X3pEW2yZJpS0juHa4zdTALvrtxfe88aX+PfZ0EEzI
Iv3w9MZBVVumNbWSvMOV93phsn+9M6BwIij5ZXB5xUJhMBhq1xzFuyLubewyYVdO
BH/niInsmdYnWFTiqLFW1Fb/zRmu3MiBJpv23KdyhqFY3XCSp6hAP7qZUkHz1fXh
PTdkZGSychTYT+L4gPknuZ18dYiKZIs9rdZ1eoZwXqISx/xk+7ITDj3cDY1wATQy
ucfkmrwB//pDKxwaaZJJmO2XXY4N78vKtdyxnPncMSFGQWQBAC/PHCIvG3yrIaVT
QftD1OZxZWD/AbwZpjdZQnbxNI1j+pbdtenXAY1LfWRhkoVC8KTNqrhS4qKc8uve
LqCOd2tilW+Be1hcaN5aD3OIdIY8H0qgMvmhyEJCJ+obhWgFebUC1QlJd73KcAfQ
+0JsqnEn0jzFPOKrcMdakMq+2WuFYBWdD7BZnpG3VX/LGDEuM87yWZUaX5DoK1rf
Nd6wNwdIN0OOXWNGXRJQfLZWN7B4Emj8bh9tulg0FUCw2OEBNhv5IYjmMg/GMhKS
I3vbF5gHPfYSrW2/wqS/59l7B1M+QRI7ZIVjAmO2s2TwbNQzqvR+kDudGla+YmF2
7vIjXIZ86H1FY282NP3PpQiVoP3Vgp02rjVDbywa9e5DMdHwQonlo120wc/nY6Sy
unz+I+wa15sADdO2Hvoon4kb6NSIE/4vNe28wT0r6P+XOCr2R9a3eUVg/iS5THRu
j2ks3RcMd+GYaPAgaRgy1/NA7CrzzvUFL/8iPZxlX6j8OeMzZ+afTcuodcuwWAEY
miWKfj29tzxhOeaqrIM06BlVLK7soZIgV0rMG+sXaMCxgbhrs+UgYCLGMj4IE7xt
PHvhCQyl3cFwFqpwE0uww2gKD8FBIuHNqiY2Hpp8yPy95gy2CtjMBQ5ssVjnxS6z
wqM+QMkd6NV4nisBhqH+Yoz23Aj3sa82oFOkot84EOX7r44eipOX/69v/MIyeZEp
cIijd0ABhB3GF+OOj/8kAqc7NQck8/ZciwS1eezDydaytk8T7bB+PQwYX0kPle4z
32Z+VWOCDYPRMUnTMtFwEgi0kfnRHGcpoWjMHyuQCu5lXN5q5nTxzVjy/rvpd9EB
gaZMOVTbArL7E10pTImGJ4aiSer7+Z5xRrRqdsluaFjiduQacbDxLKOXJ4LN1rnE
A9Z9GCmtyixwIWvWgaG6A5eJrtrHbwZCzWGmdTNz+qLuMCqTir+cZfvAbYzGrkPX
O8Zz9QWkrc9ZXSO0L2VlHzvPhOASr3MPAJFuBgo/mM6EQyqFT6sRX/XvNsTRD7s7
6eADJIcmcWVqdul9RtiHbB0Cr9VAvaBz6jR+UHTI5MteBBCts+QUBQRIuVbWzx6f
UBPkTShPW6cyUO1EYKHsj4C5rSmYHMatZKW0jicHAAo+cbE0TisT9+b1SIc35LCZ
tRyTv7qJFIq85PhhAiloG/HGFg9WOet/ZBBesFykTzczBiCmetKLv6D6UdrcUnre
4UJWzZWlpQHTRfvpD1tepYoZDKtSprNZD98Yuimd3yegp4bagFxYceUqEnN3dNaB
kY7VCEwc/isN850U9jelOtyoa97LIQZZ8t3es+PQDPmPHQue41hNcxaRHrszXmrN
TcGzjp/LW1OcwNbLITzitGHrWhv+Oi4R3OaVU9dr3l0l/79zzdYxiYAKppuE6UXl
A6yVfqkwBNQ64HViVfsr88r80YNZZGZodVut2RIDQhEFy7ljrVv0ksQ+afnnuQUS
Ivgukavl63ZteU75WfuhW74F49VKG0mh3qX+rBkHp0W1RKUCw/0FUw8S5xntqdPg
nrzLbHNIXqm2kxhYX/weGwiZGqRm5kPMaRjfsEnSfiKM6wO9mgIcUL+1S0GN4zUO
tcgzyos0vlVga5g1ADOJRCM2jB3Kchd4nTANb3eODVfFRenEfM7ECmrXdH+wVq7l
TqV07Pe9gJZSkfUHmLCkGrBfSxkE9DIvHhvM08mGh+GHwLl45hO+PD7T6aEHHmPw
t426d36b1vopixjrCzHkR9VxQYgvGeiaA3gzorTEX9CGPSykSRJeix6FbGIUgAlk
JBdIs8r75CSRpKQJJZuAoLKOEnFvRZtlRvKiSg92Ok59qfDiEkyLyOPs3V1+SCtz
3MSI5iJVFufsOhBqmvdkFVNX7bOZqrt6fzmDQQNA2w09/0G9GGUkIKKn1iWBJ99c
Pglvo+jXyVYe8KRRHH7LoZCnx0RrRnDcc7NT3UkyRqA9Q/q5JQ7bU/0wpkiJzCL9
40XUWHxKptD4Mb7Bzdb1qEQVwB9tG0qQ9FOfzD+qdU0qvScainwdOtEEhPlLY6In
NfjdxuWsMvkMv8JH/nC7DpajyWi8usJ7LPWgG307EmdWb833Jj/hcEAkE6YhRpQ3
6kqBcLcvktVYvhx/xVk9Uiy3Xurdf4x5BJw3XNyyW0cKDEvPIh2v+To/0PNcpyWa
p2FLhrvrsZZnjCWl8ZhZa48FHxbrZYwEzoILwtvMAaWUJ1m7Q4papKiCUGRgLmjL
IoitUuI05THYCnFggJpFqI0xrRHrCvl8p27f3yRpu0PfEFxVPJWrD07Zx84DQ+WV
4sg5JuFiHt5w9FJBFuFURu5CZ++rDv/5s97MzP3Vpz3aoBwrhw8dN84cYMCh6v54
Yq0FPwbmj66sZWy1JyObEnGfG/tbTi3AqNkIYfH1JU2THL7izll2MUqARtDVIX16
MpAMC9MbPvtWcw3A0YxVuudHBRLfQ9o4Y2cnDkhMCzASOJMTgeht1HXcvHq0HbcI
Q7Oa/g1h1p2eBkt5gN2P6mQecgBvDzA+9qj13+VkZx7cNdu6Uq/ojkU0lLZlB3L9
hw9t5k5kD42FQbG1t1l2fhgESYG9T7J5kBe2v01BMhcpdUf0n11zAnz037GqoQOU
xnPnuPhgSvULeNJVnALWCkr7vRnkm+inmNcUgSK4udgfqktMtS+L3Jrbp1qU1Ftd
uNIUjuRZY4VVr37OF3QPf9/TojsqSn0FI7Ja7MjjptIT/BfL2G354JpZ3UEEM/e8
PpG4ly6fY08RsPvFqw6ovU5Nk/tpJDxgbbJSoPVhiTPpxl7LSghIcC77wT3Tozoa
2cxUpjoB4bEOKNg6+QUz+nE0Z2CrQkk0oeJPF6HmLRuADyWSqx9CbZKwgVrgI958
2bD0hsz1Z+6wRF6AfYHfQ0dDdLK/BBOG1J+SfTBF2kosBT4EbZilWaEucGHiqtw1
dORUXd+yymQmWH4se/2VU6sQyJzc3LCto7Ge2uP8UDdhxtKBbySqxdQZypXjcCdn
wtDW8oViAT/BsTN1HFnpXy+85tnoZRgWfr3z8mR60oRZ8Cs0FZu3ADr5MLPjHW3l
k1b+0GPy7p1Ax4MA6Jojbvr7MefBq2/tvTEKo/iMm8TspCUjLlqhYRUh/z8P9wEO
ngO0Ci+V+nlC5hzH5qWOEGjzqHfHYk7qOmvD8SdMnsuKD3D8RDQu3i+sxSoeYLrE
xgUxBc66Yo4+MAPYH5eBQ1pPR1Ab+tIOXthCQ8BSca7jwMm6Fw5Bu9mDDSBlD0wQ
1+hm/Bf3W1QMTkVisCU6gm7LfmHHSNKnGJCX1CAAJ5dDlXrZDO65dE0LwA9n6eDE
xnCuSmB6t8yhWtGS+EvMQ64B9SrWR16z005tU1u0Da4dDxWDFlk+yyNQWqBlaF+l
u/1WIxHew57+0EK/laUfSH/08lS5L19NVdxu+WQ/B0UVwZLjmlpB0ZTsl9vC0WDg
pLQflephkZ6GcslnU/KdPEdU51FUZeD0nJ/SxeOz+N643CFGByCPNXl3ZVcsTBne
4V7dJOrqsoRWBjK/3OOKoIPqTmHEZ3YMZQ69628fKlw00eeCPLu+34KtS+0a2MMI
sSOFqA4MHEI7rnRemHP9yOb5ZLI9qylazsG+hKcHrZVeJWWNJL3ayJLh9soQhar6
JyHwTmRGaFc7MnpAAMkk6Nxk3eWCxB1ktYTgFWNtUy/CEgYCYv4onHHpn5CCsidO
5fuOrGhs+VuC7SmiQJzaOGmgh2/ziB0njazAqUe39aqB9jeqykr5PMtU3quTySGA
CcUObPPwCOVOJ762vgeF0znbsCdGsdQviaW/bEB4SbSGWAC9LfBzkFuElzddeZg4
daxv5xHt79GzK+4XZO5clsgDJ/Pt4OOLvAsiN0S8TdMLYdLBNqvOMAxlUipwa+px
JpTMiNBZcoFYo6LdRtv6Bf+dDQbVVpTJTPTRn4rI3iwvCdMFwJ268f1osxAMr30e
kJpSh1V1pS4ajjRb1toObYVK6Q1g/kTUTJuyBvb9f1gC4LHXfMefw9InQC6KlUyd
exmW0eRnDmNCOv5SMmlY9GQhVBg3iMxJGtw7Mjtebezxh2wQzhfDoU5L60NYUWhC
SXbJyhLM8WHwuxEYEuSlhT0YlA35bm3GJfFusxdGYT3p9UGyxBe/+BJA/+iW3NRJ
D3fPdQn9RuMD+Yzv4o15TxhTHCsxCefIhFqViv5widYlHPSA5ZsBYfbO1xRJMnYn
ky36LwBAmyJlUZk7zYvwNlatqljbPbmoz5Ws8TRGb7+QB0XShaGsNFsTcilOqEB5
5l2gXYNizQS1hslbCijqekYI4x0CesPkltRiSue6M7xt/fC8rFy5qCPOilyR8kqa
86gZ6dIo20OjqhWAnUM/IEqSTiKpgf8G+qSz0Ikbk0NMj909VnqOqdnavi1CqwVK
jVvvYuQxjQyy+900PCiCxm0+gITFynrz2z5OrdOJdCgZf5rtHxn8Tfo7oj4wbtym
ioHsMPNF2fUX9ovfEg2NY98ERHNlcgQvFZ5SvrCTyFDf2rAraWnVVnj5dxKtKPqd
ZMV0EKrAER8mViK8ZbHFyi2/7ttOsHqcL+oPP+kaPPOCSi7WLOF6SpWNEIz/bRXC
tv++pP85k9wQBG38PvMBm3Vj7oCYlS71h+x/yQxy82NXN05szAfiNyMRNqho6h/R
fn4uxc0CPKQt0mJBFRo3A3A9qmQPzjm6oEY3IZhTU8ty2IDRpKM4I2rEsozMKAQK
PwbXOZapzPjNyO+VP5XxlsJkm/IKHjm8YapW0RBvrQ5S/WqaR27T01oDtzVGkh0C
6xX57yT2OWpcwd0nIOWh/p/knNAzM+zbS5HWvw8p60W7141IzsUmwc1htfmSFck9
htHUoFPcKJb5nureu0cSheT9UjSGMA8MRT0QUD+/tkc9dClBA4q5LRD4+j+mM+mD
aGh8m4qcUDtt+BNo6hmNp3BrPC8R4Jqfi5/P8z0zLOsrr6t0QtwjGupWJphgYkjE
F2+iHWnvgKnuUfptwUgDnt0gAQSfA8pDtD2i0JmA4AhZ+ahAWbREfXue/y8WNWPz
USS+djrkiljNC+awwyCW9soHUoNbCc9Cmev30Y2A9y1T39d4ilITZjV4Nkp5iGaN
FtEq19D2WhzH3y9zNTEh1MnAV41I2CfqGspPfSgevwuSFyGer4dp8eCjIO2si7GB
sdw01hBh+T2pJOjcJwTvQeBh3nZnOfyyfafDflrOO1Jho/iaa6xhWY0+3aos3TKI
uJ9f679yieCJPj0waUupCg2BIwRuyia38X6swwUwm/DPMMAJ03Bdv1N2nDTYRZPJ
v9mDdAmYT1kkjbHCW/Zo/HNQat6niYlu8RDyO44n8oJcsmu/+e3Q4WRYZbowi4h5
Zz689hA7u2n4YNu3BfOSKyauwi8zJ6I1omk53jfqngkC2hrrMwCj/RbYQTzijn1Y
khdJ8UiNNVYC8oo00Zq0T7xkIeWwIvFpBHleMJcbkZ01OhF/DbhVh59Hdn05SUmd
APlAUi7G1Dv6rQUd7H0HD4uy1OLvfzn51vvLRU+CoBKLNc4xG/QKAoZNKYYC+/Qx
LyshKdi74aKLD3EaDjqrs7AIhv+vEO/jrYeTTi64QBeHd2Y9iQRk4va92+vvpran
sh0ihBST6BPoSWYgY/0kSGcwXvLN7g7wXVlL1hawNwFHi34cCvmZ0507t9qficNG
GKWOmDzBIdCi/LnnDs/84+uFLsGuZoz3kVRN7L43AMSmGlow7liK9n0PnsL/X5w+
OjoRq7VowBKIC/qCwy4lf6b8FolrPm2fZQyjI94ux4WWgzKCgkcZD5lVGvKFIH/f
L+d8nYX5rnkC6TFCj2WRq0yuVL1B3d4KPYWF658bKjuVJfM+BsGC5T/Tv5E/Pc06
J8NNxzxto2PLJDOHrMjlwqdxZnQf/8QTNiXhH4SuYeW73u/T+jRdekwsSPnKj6Sm
02QwdgGH4+QosyQi0CXxdR5ROTBVUNfns+Cz00wid/Y0qldViYKCc5SpfYbx++jC
SPeFCNNyJ69dhct5+rZOO9/HF5dLkPpS8fiEHdX1YzJ7o/84C+wJDE7QmvyPdh1u
Y02CZTrkIbyx9+Mm9tAfQB6huJgatHit5nf4H23nDmI/6gznC5CnwXS6oXfdLoCi
DmXLoB01qVXxR1JizFcDF6J6LvYTQlGxFQUXeqjvMrZB7hPgInhTt+wMJ6KAEdva
eom1kUnBbBU+z8nuRLWpSGdsVsepJtWddX8kzDho1Hm0JARv4OvjhmSj9KmQMBe/
R48ukKKacbtsW5W9Gx/gIZZi+wUlzRcoYbFDtj45MVDNiJQr2YQY6jEJ3+i+kpXm
ASHw+Xx03AIgvqshlU4WPajR3aZJv/bXZFA54i/939vI7zqnaZqRjcqS+DhjKbNi
0Jrl63fBSgAmGU2o4JBZdai9xvPJiz/4lwPDKYFH+P8fEy2C2Kzb7aBJ3wy9qG2p
bkItFEnFmoxqvdyAzS6EJtVf5K+tvVJHT/nVn1VB4X95D4oX9v5VCSq+l5MwZiY0
zAM4BPLGTNiLOiarAkCY9zLcZjUZ+GQ/Pa9WU61tfoA3rWgtU7OjNttGTFzEwaBJ
iWdiDYDC8GwsRcyAaPa6C4dq0ItTn2PwMRjiw1QJaTYMxQDfkS6xuQxhHUGjbGRg
Lawjvf8+Hhp4RAKsxZGmzxUrFI5jtOkhOYxtBHyRtL323YLeTPGt0WQ6nMexIvL8
3QHZV0eSNyozLqlIlsIjpIkll68pz3iJcIVI4bjjWYX7jAseD01ua0+KSe4gTfWP
gWNGG0FYHzUNHvl2+5PXklONbscD9gv3A+X8bCp0EO7F8eq4SrWiBbBE/YHYB3fL
LXf7Jkzaof/SSsiYXzFt4ekLzO9mzJLD1/b7KxS68FrMn4rQBagd6GaTtt7rbGlC
4Lrs8EcGhIAXrvm3X4PSArMT04WmSEYkopg58efBLIf+Wp1Z5Xhcq7Y9pbP3aqk5
z/xZzRHXBb3qqbMd0yDQg3+5MOyHTlqJY6oNtDk0+DXxbHKWPAcouq76ypJlj1/n
V+2YTTiSyIDHMcqssv9W4vk05sMaMgr7zD/ROmgY4DSl/l7e4KmJWqCIxBuMxG+V
ijhZpfgm8BUwwxecu8EdXvXUhLbG1Q8ErS2X0dw2Mjh/RiwtCnS40QkAvJyYXs8R
ThogPs9z1NoFek1b736L+1q6ndpjRs9PRuq1a2C1XYa2ObM7sNl0aoHyci6zLpJA
+fT6VzKpG4VrNQqvUsarPJmW0cXIk5krayizammeFKZ0ojug5H6zCdvVfG/GMwqZ
DBrdnuqlTFoQdp40HvoRlgjLoBjcATQJjaJ7fkIzlbaj84BryNMU8wVVivMImIyE
5tGqEzG4ybVTMFSlduthMSg/vmGjvGWnf9+pG0hPqI9YlTBkTYXegWun3X647ezs
NvkJrMD/YGegH+vu4CI44G4iqfzCYzCKlAwwzxk5+f6Fm9/RWTztZryXm1n+VQzF
ceB6m6cryjb0NfHSTQeMDP7AFc1v4/lmAr+VMUqy0scfXGjfTQpUmvQrKfTX4p69
9b6/pi/uQdn7K3Sa+XvMqDtWo/QnTBghu4axdKhKdetLo9qdpyooOi7233fz9MSZ
13xUsOgt2ZoWBJ4RS3auk4StmB75nFmskKH1GSANcy+ULqZcBLAqbea+K27PtcS3
TGi3Iq6BYW+u6PnEvepkDxrRu1EgJYeqFAdD4GI+TWs3Fj/M97DY7+3Yl4fi2B5V
VfMx3nyps1gtMNkGfzwyM7DUTp+W+809TrTTsZ+g31t8CS6ZXaUYQdCt2H4fg3/E
gP04X7PcF5QX1X922VZ1IHdT6nKT7OBOQS8Rd3fKnxYDRDbLiPSXpdwddqx67imH
LsKEp1O2+cyvcEJJU8YWO9Gpedy0WUE/Z3HJIRiPN0bNSxiF7y2KXpSA2EVugm7v
iYrUjKK2YLM53t85m3TaSxI1j9fQl6pPyXgP1gBxogitJ6lGeg5m9N76GI6e5lEj
SNyoKAHfS9MVFHjVRZU475mwl8eP+hdWSSKI468MmVageJxlQ9vERFCm/gTWUOB/
Ypusssq9ZQ0KWBsD+vLkHbr2S274Km7WJDPJvJVVnF6RyGHUsJk38MG3PQ/AkrcZ
VIA49tLfp2zI//EeiECSpjKa0ota8Axvl8XMjEiAwpEHQXChJYrZ2NNvUwsjpTdH
yp36FFA+2BCGJyyd0Q5BFZodcXI6Xyx1Krfe/zHk4ifKVJzUchD47n3HkFSJb91R
A1ReuCKbzXuEVG/Ribc4sUKMDmzQQ5XS4JkdqRcEXEVmBL2DSwTSmheiGxyq1Xyw
eZI9POKps8dTX5mbU/nwxdY2FrGzS/pInc8TIQ82EZUI8Zs0Lex7+futeefAx9EK
nljDoTF89Qm/G/TSDPv/9AxBa7W2lAV5dmUp930qwV7Z3NTpNhbkEmr6DFiKNeFK
fmabtq7lJ3Nv6BOgMd/m3EQBfEFy53Pm+94TL8IeJtDyCW7ktjWnsHidMd67cM8n
coDpun7xfUAmjM+/emq+/JRsmS7WAwviVHX1G9tNzsWX5zExcfd2u4yUZa36wz5K
zqSf5Xyji1/BD0T5HdcljEXU73pJbqtaapeOQlMAOjTTlsTz7UFQZFEKQFy9gXx7
x3+LtzjMpnwbGGCJaUmPBPQhG5mn8CoVR2qdcRyO0SjMoK8zrCMAC9h3PAF1i1ku
iYu7xOqHn1ZH4pgHGumU08e/qnyRldRKpMWIQ2GRrxMLhAj2oClUMl9xPTgva36k
Iiaq2tifl/Rg+p3OZJw/mznC/YG1WvaAmD49q4iaR5rygCU6j0UOaWCKYmNf7sQH
2MdyCHDHQ2Q+iK0TgYpRvSJbohlqlv0nrffyaCuMI9lnE4SuPRPpIjSCf3k/Upkb
Hn2R+FL/WrhZFOzjcc/ZelE+/eyeTDACz1ycJS8PcFVPyEIu3GvRx97fY+mRlnQ+
IdEJrnE14kMz1M0UZ9UibtqAz9JJbCHT/ZvPYh7bQv/eP1qjfC284+a2Zr8CRIGb
FGvyZMIr0rt5zLkon3bGtbWWtWorx4BDxVR+poLBKZXsDiQXmlRTPYbcirv8oTgu
2hwemhd6OTxc/JHckRfh9+V0sI9WIdkjY0DMt/2jZO8gKXXkUYcBR7gZDA9KM0qT
6H+1w0tn3fDySLzfWxUYZLgcfhadxzW7O+5QduHCp1bqALtjxf40AnIjVX15VJ5E
uVXxy9hVqVUNnInXXntlTdUTU0KcB9sbCKGgR2tm7mWgR4WSP9Dn1fMxj7SrwNaA
SZSVhJm9MUvgRX3Fglfd8ww/cBozHQ8K2qpJ862rKiySm/n0dRHwG/4qWHxKW7wh
e87v4DbQnETFR0ixWru52oh2vMBBNPTpLE3/IGZmnvJptz/SBVzEQZWCw1tWWQb0
M/5/Ba5RGLOAxDxcPdymmJwEqKeJ1pN8+0g8BwADAFjGnWdCKX/BKiiF2Ra/1jth
cCufdB2TtuNK88OZOS73yCjwIrq8rJGtErFsjsuvI5wKvppZmxBQhuBnNxJNsfya
OYVkA6EFQF6d4FogOxPDhV9dCTjEucfjKg55GzdmKUkWwxU4bU9ZydqA4HU+3EPv
Fvp+cAt+aBtYsS82KFAWfFmPzqvzOdCLMb2KwrrklRXkArvme+PxppLk+FQ3Jsyv
Z3+KHmnOwi5O5Y/J+TBDjKmtoeAS2CnBVp/4RDBidW8TemR6/JUQ6wwwHWh3JlMr
kqDytNt/AqFE/P3eTifcI4z15ndJOYwZN6yjq6NIotcWdMR1SidRQ+qAMeGBHOjE
S+cZHoWSrfedSy1oonjVREEbav55ji1zbj3wRkuJK6hk289LxMurhwLQPJD6qZ+D
KwsgiCcXbvJCgiiSbqYyq/tlS163x2LFf5oTpAP797NEeZ64fybIMtXzvHF3GmDu
kstXd3+b0SkRrTGiKeGjncylS/qYbxH3/JsuNPIvVP/QKjXF3P4vxdkTIyT7cW2P
BF2u8wgifX12L/z+TypD0o92OWQ/M1/3otfv2bPb1tm30tKHgMI5WtsjmFcSdcPz
wdUvg29PFzXswGOpmnXVyk40mrMMfZ4qFEdrvyJO6sJM9uDe5NGJndW6WXXswKZ6
kOfOaqKKMULwZeKaRq2H9RG96eVQdlxlBASZxPRYQ0rc0bcA1b1ZBRTc9IZp3BMS
tr3S8wJQE4ssWwAGpUl5ZQ4DkO7OFr7fGV56KLDQteYpvbO3Orn2oY4GQi4VPbpc
cV5Eh9nN0XstWho/dUO00UZ3nZKDpDgeutuhRspRYoaRMI7VluIjgzEh2E2Mh3rt
BCA3KZ6zUEquZikkrJ8/nQOqa1/ILnd31Fdkkmt8PwLMmgiy9zssDLgMoyVASg4G
BXGBCnEYnOZtDpvBfiG7qRVVk9FbMd2aCIbZSNrB1RXgD5Ruuv9iMpb0vM6qnBiI
K2nJIo2TYI+eeKBPFMeycuG+l7Uxc9xNi7t4qwGTFuIP0LQ3Pn8bmRmv7w6bDTe8
NwgbxSsdHZmm+XVOesDblbNjy0jalg9h8IJdlKMzf2slyN8vHlGh8kPdKHHgUSQQ
BeZqTylbEsX096gsRqWmoA1Fx4HctUL1SDro86QudHcTvSsBt05oZkELImoS6qSQ
15OEyVI/4tmFGGihElvjWn+Iurifa1lhphqpGvBBJnpAvrEXE6bocDobz3udqjQ6
pBr9Lt7rGx8xPeUTA0jmp3RiBVvSChOzZw1ktJdmpgr6ZNYApl1G2Y3c+9lgKBrf
DkPG+1mOBBzur/e/PetK7rpKPqXBiB/gXqzGqAqokbeSn8Z65wWg4gJzhpopEsch
9XiKQDAQJV4S9/R/779W3aO2AISxfrgTQYqMrUmzM+0PW9gxHiDRBHFwkAyKZUxN
RpWOyTl8q+Pw+tp1XnleO0kKlx8hOZefB6cqMMFvR1zvMZXDKHy7d+QD4ei/5EXn
IAOJXjiNgF8WvAqkO6feSH43eRvlg26ZloCNJbwXew9FJ/oHe+Ss0hw/brAVgRnq
PUNeh6Ra3Krl/d8BOcSJcj/6he+KIVw59h3wBmD6QWNFn7oIb3Wz5fM0jTE1ni/C
bISCe70pm9bTAf+fYlYvIiLIr/VK5gHJslvtgyW0bT0qoZNH5ZP9+3uUygA1p2vA
mqUHeAgGvnPY1TIKSvCd/vVLHi5BLlGlRQIlrYtTXE8EJZmhDeTHeceEUkaBblcv
fX0aUWhknYAIsf2Yx7XD2K7PD+vSTSKBcRdZwr7vSdj/PL2ofxyiWr5vmbBthdF8
S+6B+Du+McS5s6im2ap3CUychKv/Qtr/iHnKctt1aMfvEcjLotvAqOjXVG12xvtz
ZPoNRol99yLLHFmEbhkkgixgBrYN+dYJRuldTVKSEmtnatSBCdl/uc7qR19sAcW+
wqQhP3TufP4RgxDPsP7tXO9hfEfuwtk5SPJ+G0pPTjzjoAbEh3NhH53gEBRQkgn3
7gcsp+JjIA5b1RIAt5RJ3O3gQZDFUwsR0qWbqOnEwxRMkckfE9xez6bCWjAN/l5u
zi8q+JV8r/x77pfHNYaY7Uxe+QZrtJlIulpU70oi+F7yoBAbDw+8hvHBjBIueb/i
R++Qurl+xPfgE9gmWc2b7YQEiVCU68RVYJZG85E79H/wpsT8RSl9HOuM53uT44EO
DVzWaVURM7zEbyPuSE7UsE9RTpjuSBRCJ3GGiAWmlPcGYWrq2LbAc9ND2mkwNF7V
sE876XchEdHQwu+jp/Tx3MJCJ8sObDRkpW72G18ahwvNFJxbWvB3OdrIIw4EMWTV
Zi18X1p4S6fTx+UgwTMD2ZTk2hf2DSbZD6TV+2h73f+ogfCfsHpkYnZgVPsUxtU/
SxpbEBe0YXDRCHmhVhXBefKhOmNslD8eA6Sdx0J7glYDVzJOEBAnl7rs0VDw818V
yySIZXibMcJWTb79NQ+CBfpF5EBh5eGjk1qf3Mgz9VEz3WhaYjob1L9NHnPhVrBq
4qHosrPLN6uLa+Tcj8IQ1FazxVt4+tuAGjKrxnFcNeKG/p8WKfgThfn1pIde0uf7
mjXZTGaPiTBrGXfA0RHkbSBzbhR0KyaOIPu7bgWyUQNnuQ9ThQwZYtsvnj+hQFbm
R9rAn/xVDbF9tN+U8lIGIgbzRwsZBKQVWYZL+geKBfKiE7wDWaZJBGOgjdFh97nu
iEP/PKQqeAA2Q5doeVlQrLvrg/ftW/RazBqPeliw3F8/qZ++vXV3UDwh/v1e8xjy
Wba1NAkY9scMO9mfytVjp3F54Q4dCe7raAQBFwCoVXH2/ek2neg+xgO0RDEMmx+c
wT+TGoEliS9JQT1gLbQ+OKnOBo1SJQS3eUSzNhMxf4tYf/eTSQWmuws3uUuKvX/x
E9BepP4RnHM89+wlcJ21pNNRwsZsQmkjFkG3FsEeVgNFi1XKocDRmWuwMXggQT2C
eGHq3qsci3RF/Hl9mTZCPY3ma/ZFqi+DG3ZKvGeTeF7YmmSthBkmT2Oe3UMrdSaw
HDOcFoNsScT3HEvOqXvU21frhOshuvw2hXlk1glF+B3PvzrGvbLCDJrcEIGJnMWz
FB8ITfn8G5FV6nBmyZ4ym0dB4fzoW4hWrsFY/fhbBHA6GHDks1LbjL/3omF2nubH
e5eugJlvrrB3+w2yl4hj5wgLqR770rM/YhzOEFQfdNhIud5WH/HHj8KEZeXmCPJg
MBMhyy0r+GbL28WEkEdvACgnxMrpnOZL/TrQhavDzdJHiF7qSGggQ43GtxpTxA/U
gExVUJTXyLv/dDhvu428G2T7KHXod7Jcz5cMOZRSPybCIkeWxSyuXy0U7IK2ibWa
kklI6811yZEhpX6uwvnJpiocKdDxHyPfGOwQmdktqW+7IMabdGb/F6XvgsC8GcxY
QKVEDbw5pRYbFjS4Lk0WuWb9isKTmMkBBoPc6Ei5l8THYaywQXubP3+jtdg2ydpi
nyfiedSAMTwrS2VLFr1Jlutb9pv99gOWZYXhcMtJL4h+7Zj54IjRtzMUXD+aDpRx
tBV+2MnKEH0Aoiv7ieZySxJ3B75/YQXFKqpY7dRyVJoz+Rs1TZF0nrX9oxSrCucB
LXpwk0uoPur/uQEI45yN0YtdxQvmCeiCUOMbAsLlsKtQhK5oazX6v9Rhvl9aMAJP
wTrmgZob0SCp7T+/CVLoatSlF966Dn9Xa464UVZMKa1ch+wXG7OIUr1y5q1PapsQ
7vlIdJlmI5j557uWHxVjkZ/agFk9ZqOUAO2sAZXNt+8SFmq2bRsmiB/TC4rm7lPC
017Dz2c2jotxlG8mYFw7tnBO8L/0arTReHKeXdEy2wqt4RrAj+qqzQOv8URe/p8D
VS5+m9nzKofRhKIu/k9InchIW//xVdHZPBHrhHVIAyayhLYjrgc5+c/zdp1d4Xph
f1gGxDHo4g35JZ5EkoWcfR2APTL0x+xdn61ylIZUAKrwXy0TD3w9Fh6i4uUYFfxt
hAUnFNZWzDy9Yr1y2cjUHiZKVAUSMQN8osHg1R24FoZdZ1Y8HsvkrXloozKHBf0V
LFjd2vastbPc7TCfmJK+pWTjM6YEEyDSRxwgjH26vDfFGB2iC9jx9r6ADgnW2lsS
TfisHnJEU9yeI9I4NX/l3VBtIPb5E8QjV9DfMD/hQTbnvaeOLYUTVh/kQ/h3JS5I
hdMX8U/iG5tsFu1JHqrDuqLACbDwdP39vaB6kFWTXTtIOSVSiGj7zReg1EwJXsvf
WITBlMkdzPtQnEuD+z51M44qq/7n336Rf2Xtc4hEPrShFb9qVQ0AnnKPu5cLhdNg
nYuK3fo3R8lT6Lh3Z1E9ErVhjjPLYwSWGHfVf+iiXExA6SpzmQL0XEPCYN7C+O9+
P8zQBPxMGMTa41Bi6/nMtmRODFp5HjcIOt9kkQvkAHxn3pooRC6exyODohEZXdQR
d+OQ8PCjceIdZb/aRtR4emRfDYU5VJZgE2ObfyHBc1crmHT8AQXdHb/Bo66LTjr/
byo+f6NaV7BA4exYDgmkLZynrNu017h6AwpESHx9cxE0b7Tti9rl1kz6D6VcCfhx
U6ZDfFi5w6AffOi4oVBXznycAq3XjnplZaTmTqYoBq/S6PKHWp0yeDragqanUzBA
BGNogmZsOJ3rJs0EY0ofQ44msB5YRI3z1++XXlaU0omqxXREUf4Aw0HAxzgNr9Zo
OkubBkNfpnSL9hmoHFf5XfiTD8eFMnwINnLqOiMlSGxp3DFleg9zizmM57aL1DAy
+FS+VAAp2PpF358+AEAd9bt5EwKSE9zRKRk+SVSmx20pFOSBpJ7x9c8NZNlFAHS0
f5CwwhTui3ocBQOVhiXIa+6JZKxiamtiLYCtqMMEbxqlAFTKHxCU5Ie0OEb/kGL5
OWUVmJSo27iJ7DEeAh8uDwC5XOs+LOrgKjRJmkEyXDJT0RDk/kDFGVJ3cx0i0Eqh
/0CY8+xW8u2+X71xHz6csDE/mFcfCaL9TPWZy5COjlKPWy9ESgRaMEMYeYWXDpsD
BPr/tcszKZDqJ9g3xoddv7Dgvv0xIAW6gVc9uLbDICyTa8SWJc0v/zqRHsg+qfw2
p3tgsfaTf6LBcq2UB7p/ai252TK4jvYusr6CAxbQZWUxnkr5/XcpvyeNN1flhl+i
3LCGv3YVbg//ul7g3Hj6eZZ+6BJQazuyxEz5QPzvwoTD4FnMqVCfmy9NS6Kc7LC5
tCJpEapOb3BzwV/SyNg0OEveLjPnpAMOwq4jKKRGBKmbQ4ztbhV+9uEcq6KsioQt
0SikWFcVTjXFkh2N/wzSjPxFI7MvPgzgcwVWdw1e8W0C+3tjOROe3akQGJM73ni1
Cm86MQAfpIedIm8EFLRp0ELpqKppaCyEV2t3MR5fNubVrS/JWzzh4Lec9k+I2jGx
xm3byAcGaxeJ9n7l7zgI6NKcg7tKoVVpcJ+AP5ZiPMAlLrWKfhrvqPcy30slIfn+
jC53D+GpUNcy4sXcek4GKbt4H8O5BWmKTtZrrCtVUuwmoWREmnwzf1GSwUH8pPMR
HOw8x1O+J8m2kDKuOvIXhpEAPwzS7eXPa677XsBU3nhRl0I0xFbLrG4TnfGFnyA0
wpQIA/T7Wcz80mxD+pKTRtQAMLG0Hf03FVp/B97g9y38NgWW2Yeelk2BM7Om990R
6k70DSbl5KCAUTHtqSlu8kxNvXBO5LwlBaDnat45TMllwNGSX8HmNXRIqS3e/sR5
x1Rku49cxvjnR6Tm1qZODz6E2ajyyxhFKVsz2v4UIGqhy0ig4gVQxXUug9umzWq1
Kxie6hG2MIt07jNiDjySnJ7GrPfDbVx21FgbOWc2kMn+eSD9vINPd4ejSgG9QWJw
RnXP0AlVIZQWbMIglnrcmjPEwxr8wpwJYSlQwdLsXo2DLNhcID1xQ0yW7L+vJiae
is61E0an0kWpCh5eYvAESl52WgxkyoydjoX9EsSSGNT0nDX1TSXqXRwITKFKYj5w
Gw6lUn/3Msb4zPoczYycKYI8rYN7XxK07o6e/wxo8Tj3mANxoYplTkd96dO+K/Sh
t6z9tKaM9Ez1Vn2DRwarkQKz/aDCCY4cLmDH6KN0+9yeEuoqti65jbWj4/0DR2xf
bqSF+HEcuusXR9kHU1FGj73W3LLbOEjYOhP3d5eEg+Zoh0fm0+dqvnnArLV9utt7
uiFPPmFSSg7/XqyWLfjIgsQy4douyZRCSHgVr8YSixo5Ydy0MjzoUKoAb4VqSt10
nfqrcFMOMLeueoK4kmI8pJA9v0zGGpTaUlQXB4xpiUVJcDpSKe3RMoZ5c6xkv1Dr
OH4Nu0ZX2w3YJ1uJNpka9MVM25PhbFgGWqdBFyy5wwGyag8NRDn+l15Cxd2xfITH
5WCGn1rqUxA663w73gojrAZqZzhQthN0QKuNa7IC/zqk+Zj9LSH+r7tWCfL/Apop
3DZyuaUu51HztzwYPTgab/4lbZh/urqGYGQNIaXt3wykpruocT4ZFA+wu/D0qPV/
cKrzaaiFHPZ0VhhjjfNFFk1HQ6soZfHy2QBpFWZuUmYX/J5l8qUAjDz9eCwSO8zi
c8mLNNWWhYc87SczfSDGK41iLIVKuFUqJJHfl3RSnRFVEbNgj8wZS6vk35202rCA
0qyeWajJMicP3tMigUcV6NjdM3k9ky5tCGft7p1yyrjQpR4JbBI8arDvewh/y4UR
Or7jNV8MLevu/OurJm4TX7xPDDey8il8DYldWzvbXVBRmKrz66tG5znQIS/bmhXZ
XzpgajqYvqG/QymlpF9Dl9hVRAMrAG8A1fh+mqG5mUiD0bgQSQSb34wI9d1aFoyS
rcKq9myo213xxOqcwdpibGBccyaC2+lcWsrD44IaUutxdBWBCw1xRbPKv7PZkezp
jBKJsPZqqiCWJ5bh2p8j4Fh/DZn2dvFJgb+ee6OX1GWhXCOTffh8mO8Nql8b7X8a
BSQxb1O3osHh4e7YpattoHV3TJQThVgmdrFE967QRm8MOt6pWnW6GP/hVyceJkfT
T6D6RiG5uJY4w8BZUZQithphkKQenoX1q1pYymk5+FnypEA7+kw8v3clr3pvOR/2
MEx6a7zruECa3so7sR8kM8uneXaNDiScq4rOkhgTcyiZKNp+YSd8Qp12bh0rqNby
BS7eDKHQIMY6u9VNDV24hIzVbfbdVmmkUKVHPkR8KmbfKxY+3NezUfc/t4LWZVky
x6hH+aTcmk6FTphkDd/MYzxd4Bhe0ECXuVV6mbqt6KUx2DJUNgpvMEeiQJ9qTzYf
xEjd8DBWObdh7qlUSVqElvf/HiF6XTWf1LZISB2HnvedIURgNL8uL8LM1v9cuG4o
MCiIbT1rd5PiZh8o0lIdELAWXGY1y42wogVXd08tTagbmjyf5yZpSC84iRrgU3Pj
pYH0+cEX5tGtiRdfmfUEdu8GodwPHOlOVREViv1tLqc5qSj+v/AocsilYCYEbzQd
VpDYK9HAwID0zmRrj0U2jdBlE7g2XNmiMd2N3xGENAXhRNKu9ia4Zs42gDDgyQvQ
KOMHQ9z7DgZgwHASX7aegPmLi10Qb6wbWrUy9jthJtMACZKceEtzKEnOVcmVfR6p
zoTOflxoE+DFX+/MIiUZskm+I01DK6AFuxIDLyi1HauMwplO2kHYV801AvKrC2Rc
El4aI88Jh0ASndh9zR1JLOtGGwHuevd49PWhsDMU145o1FGLKalEiUdkV+06qqRc
MoLlS2fMVWziAOZYVJwbYivcPLwK/5qqqWkH2WJvcasOMIBN5yZNLmJH0UwDLa6b
9wRJnsd5Ddq2FGGv3PQWfyEjWhBLzITpmhkyJrVyPMdOG/eCA2D33MWOupXsAuFC
fkX1Fuw7bOCIjMpdnI7zBKj2Lgd9b1RVgWivP3R16Rw29lF2SK1dbMO0PgQCFSvC
Hj9YifTVQ7goa5WTXPbUVpmpHEBn23atYRP9CyFswW+FgMv+xSNgEtmQ8rtsXIP0
5RoIn71Gxo6U7X5NBQOPMLHs9mU/CWlUvy9IHh1qrnOR1+BomxHYyYx/UKS1RNHt
FIHeHhTR1yTjMqjPBBQC4FFoEIWNWvOc7QkIuWPJ2afHtBK++oPbSS3ngAxfRQn1
HUOtMYQvOiWhsD24PXFjki/7KHAUZjybgalZN04WLxWsyVFq04PgLvnbdYJSzYUx
nUg35O20aQ6mqhmCCwye4T1NFk0xn6K8NR5nLL5H8MXjMQOiFZ9/hWwbEdiIKVUV
NieuftP7Io4c94Bk3ZFZXVA3WEbohaP71gr+jhINT7xD5qVRdlrbrolkQmgPPWTE
Kon3umflJs0IHPlt4iQKftPM961tSndpCmivDx+gcp+mWL3YDbr5G36KjKLid2U6
F6N6uS9iDM4LZT8iNgT4NBlUPn5uQ6eCgscUBYB226CP5ghKmAxgWYFeQdr1g77E
USSbzQFVJJI9QAoi5K8L5i+NsPTXUhQk65jVjqDla8nLdcTPiiGZ4WievNsii2Hg
xkkIacNVAQwYx3B2WbUbL77nc7HTjo46ZtmqenNkT22jtwaC50NGZqpFmG84n318
ClUOTeLQEYaSbbNhqyGvmJx8vhqt8PRygy7KNGp1gGrH78KAQyG5pCcQyfFALFPN
isMFpldm90NjS7LKV8X7uKAsXHMXYFLCThVu9w4NvCx/W3id1uEREK42OM/C9uDV
zo7nCeim6KQcNEPkX9XA4+JGROliWx9+9INQH7VaPb2kgofNrm1d8E7hPJS5erVe
GsA/XqQ5UstWGt5FRYVvjNoX5smChyT+65tvtuaJuzCCVHCDpSjqhtTxgPrdauQM
higXfeD1K1dRg83gFiUtSKR1O7kX9im/VCP6SR+Y6sgE8xHiAcxjTFscgNpgcIza
/Z1FTCxby191UXPkSh5WUtWbj39IEsX9q580tfeOLH+4VSgXxY8UXa8qkvieUec9
IHfWJ5VDwWg8MyU2ieuGwrEK3w8RVwGjig+lmRvTrQpAkQzdNbE/6Wcs0F5UlmQO
8LuT7Ryfp9JpqRgB7Cbd62+c4a+480yqceBwg2RsMr3hsBQYVc1Kmg6qAXEImvg5
ys9Cc6pUIcOQAGIZheAzffEZPe4YvYUtWGtw/IAbMHZx48t20HoSvAaR+obouzAf
218vdWSEEWk382rWw4pcY3OsJowzixijwRMUCnBhXZjg+Cl92MRRAqLM11NikGUF
3t0uqNBKDc/4ncTl21XO8kZloj8VxWOfhL5CrGcs+JUue+VUGI3w3D18HI6tKUQ2
y+lMwp+WpLnz0jk40oqd8evetJlb1dJ6nokZtiBCzMGcawNqjR3crrnBJkxo+mqe
+DzCkFYkrn5Z9eSRQifAoLS91depetpopMLtZhUzUjuEsJ1fd8DPOsvi7fWYhKxH
YJSCdSeqEC0xNOeg8T/A6w7yeSeI2rm9dHyiNXNFASbrarRipu5YHNYg3Oa3yj1U
tMrdze7zx5y6gRG392KfQ6DEINW2iWIyUrguYHUUqTgFGOwfWo0kQ1n86Z0nFV5K
gRc0h+1XTJaGbz3ZD7cbnNpKpoWuT6PPMhmsvJc9ieWU85YMYojU09oHkyVAAtA0
+dPlVLGMj7jhykbiV5UpLrLD4Dsj7RI9Ajk6jmTyyDNiWWnTxW9svyf+KPAEC7Ct
tjNqhLceF1zYnczBwnMppM3b3N/EAqaW5SRaXd9lJ9ASLTu9kD2plv+1q3QZL88C
MHtgi7G5Rmy0xFQahJDjM0P5JNzvCUL0AkJ9ALjgcN2XaQl6/9zpAahVeVlG8eub
JrrfNz/+2BiSQmKBYV7jtLWj29jeQZdcymJFdDEyTASbXgfshcDGpFHlNI/skq7o
oWXYpTEN8Jqee1fjlc662ohkvnJOOs3on+y51yV7/qpTTzALiwztOO8XgXusEFEt
mPWIZitpmCcS5tTJg2fysm8masUF3YVIRNAfWOIXWD7y0r0kfl5idrxdvIjCjqXz
IvmFA7g0q6GTSKq9vjIYa0o0Ylebs+eWj9qH8c9pOamTOnLjL1TbJQPVB6m87EOn
hij90F0EQbV8hjuWvif/cjQKMYN099Lz95BhFdvq9bDucfnkLkI1tencdskjvSk3
/HZHKdVMBr0wouXOLti0isrvAjOKWHwThxdB4xOTzpSIqHobja2L6m6kPVHfxHWX
zOebV0mKlcOtY2wesGMtOY6EawRfg/OtQpWNVbo1Q6I8dcqRlawpRXiD2FLLommP
tB4uTusaN7Vad2UFH+/vbRp7ehYga2F3ani+7qOiqQxXgahjTdXpeffImpJq2Avf
rrOZW01wZ4y++r4WvYoY5fQDE3TugY6wqbDwkfu7aQ1ynO/wYdHq0yWbz9ONvs02
8tXIsQZdNccattmpQFmh8IVbbzOswULpHZdOMyyXl85Re/HkxzVsAQmUn7Z4lNH6
x37JSZTe9fhSNoQ6M1hKUZ/JhdfpHYFVqtdiABBtTVucZ74kjNEIx+LRw51HSzRZ
NMAB4z1xrAY11gkFVy9uFSYNB2ZuOffEn8mxGx6gnxcLdBoGu+tYBJTNeQexsCAZ
q9BvP0ENzZD5VsepW5ldwPs/wBu7/P6gnl9Ae6gDZvcA3lstNUPviw9+JsJYT7K7
SNHa/FvYXIclWFHmZZ2WLulzK4/nzkWQukAXKW6bVidyfMQcJDA0PLNGzqnOPFv/
Q7WxdQJy713cs0GSnqOUqNtHwFe2rK8pe2b6c/NaffLsA3dE7cwjyutCQmeezadc
M6vS5mWa6+lFchcQrTkVu1mmQGD5sY8hG2VNLYC/5mI9Mc5kQtwayxKaRHZ1yDRF
a9SPv1oJ89gl1LwnLO4n6wtPrzKSYTw2M9pMLvd9EnBhjj+v5wEYa9EPIHyOUx/X
Ti4ik/er9xYZeIBk97cO5pynXE6Y1QQ+6w8gY1pbPMqDaCNXxEYMIKyydIJUrZm9
qeP7nk89hk5Jud59ihq4luVDmK2RXu947GznsK5Vu7S5TF4xyViEBuFbgAl1/Qgh
JGVqaL1hlxe9uhD803lcb5JaT7z0K7L/wTJCMClqCIojTbtRtFryVxJevDtODhU1
iKJbNiWaEF6sqPMerqBD+YZUK+ZAVXoOxda9V4kTI3d+9+PgTalVc3+fgJ2bL6IN
4fYjGBf5TxJdeWjqOAl0EmKVlCh/t42+OmUcre+8yLqNPh8FFPpMljvIepzXDG93
CeCk5Gj8YcpLRqV4TEl42Wu6MkFsiOGtD2ep5B8TG5G+zamn+YCTNxS71tu8Z5D2
jU8dDSwv9sGE2nDc6gHphoyHh74O1/q5kfSjGM+kEF+vVE7TMLGZfdkeLszTc+Hu
ykcnM8mbShWeZnlEViLcVuIDGGTYgEQ2WWcAVGeC2IPThAeSF9oiuDzH8Op222Sr
MQmWq/GpUJe/splGKu8T7GVvHAUW7n4Oaji9sIODDRZAbvfMOcqlolYRqAEQNDVq
OY8sXeExIxISPLlT/mkJ0uQO+LmCzi8IVpkY6SHAu3TudeKPwiRKcvQXe6yXjqfY
1r6jcOZeI+B4y1KXm0fxIu8gBjBQmqteBUEpJc5z1t03oVSiluQJYRgE5ZofYBVa
ILOSrQZPJSZPpKFnkSTPVL9sz0Upx1TEgYldNl9k/ad3UFAsbon7WlHXcJAN9S/w
z6ZXTA22naffUgG+IEECDyP23Me62F50IvQBmkUws3o/ud2BKpg1SStJ/9E7aeZd
wtJcNvF3JzxVGCvVVptNPmQIJpBYsEYoD8VBt6ByhuaulkOTWFGVn4HlvXbcls/Y
WkIrWiVN2JEB5XcGgqE2i0iYkDIhAhbKawBrXhucLeboF2Q44FwfMRoqgK7+J9k/
DBuCoQF+BTqGMxyqOZXEFNggUgaKA+HmPDSIsnRPgr1hqQxwlDwClfRVr7TWcZGq
bJR9AYofdGaqshxoOsGDH7FhK7mcObra1pn1DTk6qSqG49UF068lUwsR62lEyou8
UtX9utEz9fsZwA77sNKtyINgThyam20oAg0hbDnZeqqfhxB55VNexRW8tslGZsKy
wURivyPVx6nmYI3uRtQMDie7dO59ZKWjdUiq1HCtShc/wVHYyIZqrzfcTEgHi1X7
FdPzQ2RHK1moo2GcsLPd240/qc3oXpxuDrpYu9LCuM8a5xb4vCRtjDD8rJkbWWUp
9dFtvslHp+7h7/BXhMn3iLAtMk1dS0Jz45oPDC/d/s93WC8gIsjJSv6nFx7g86ug
vXZn7vY2lYNF59mFbeI0ZrKFpfT5fDAGbWtxMkq/u/wnrvfezUvlxlJCR4V+3eUS
ONAt+0dgXCoMih7Xs2WitIWp3v/q3oanj0w2OuHocCkXGGIGD2R2zb6w/HPbHpTp
gnuWwQA7SoPtIjH+ZcEAILanX+FY72Zx0oKIa0Rylyyo1x+UMP/WiDkUSwj1a8DR
7J7XN/dM5aT0w5dmDQ6E3IhFAW+DyuoRFdh6faD3ErTH8cLj2tainVDfPL7mPMyQ
j1NPp8wvmuKTwBZPZ9LDHdU2cHIp9emnkCsDqf9AdkXgTxApTCsgblMjf7DYINqr
d3OWutsX1Dtvrm7klORAtRn5HrKIFQT/swrpoGr2tZ4Zhsm35PcPRdcxDf1xChtA
AA1i8Il6blW+7TF4/2i8Zd1SLfP6D5Xx4jSxffoLLVhLuj+wl2+802k9riKVHfC5
qGwMrO4PD6jmCgFHiS5ME12/MjdZnsw8VMIQUCnKMfrAeVLqVlrZywW00/sece5i
EP8FvAAQ7COjijB5MMvtq8dExJ2GftX0uJUYw/Y0MFVD5WxU24H7ngr0zVgcoJbP
Ujc+sXO42d3bN7lOvoIbJnoh0oFPc+ksMEk2SBA2WY+XbXlBVJuLn7+bJ5My+jFW
cnoNvWFZVWp9RXzPuH/g+RxK+/P0wScUuypE8GFOJo5ZA5gPrPc6zHs7kqYXipKE
VepM9NOSHFtZ8iB4d7d+4xBHlqU7zWLYvKNSd/T2C0tjc9M8h24Ab8o5MP9wjvYg
E2KyuIyulUTLU7kEHU/DyOA2JO6giUgk2NDIN+TvAn0mS6loHMeuHJ4zvwhsejEy
eccH4dt/V8qG5tvHNkl8UW31o7O+qQVURRoelY9hRCRjmdsfe1eOMd+AJhJcPuaA
bfAg+2j4imuOF5jwPLrovojXOOVAS1bSJQHRRqatcnIbwwCqtyJzz5p9+LAkKqMw
he/z1e7ptd36AnYz+Fq2Cek47VdKqU8qgDgPFmtv6Q5w8XwEpNERlfBY0qRnZi3E
uv6YpXLqnzi3v1/3xg2eQ05SjcxpAcxOmB6wkNygn/vq6QrxyjTaT4um9u4k13Vi
s5NukHtZEO/3VV0mLUmGFe37KtBddpnQ7kmvnprCjuDVXLN+XPxt6Mi2g+1xhgal
XxcXAdPUiPUhvhIW08yN0YZjF9SoHcZS0s5gpR1kaMdRnF3sf+7We+0EBh4ioutb
Tj9c0daIx1gia3GMeEf2eVo7YP/LtcQXQcCbUrn1AGWuPg98Nxsx52/caIbxk/8s
o1DJq6Ie8uDmlpAcuHtItW9CX0ELchdshlO7rekEz35wM21kbJ3dvR2RVMuOQmFd
wtY9SyzuixErohJzPkSMlASfNFX8FvaoTOU+3kVn5H3gmUiopboOM5ZjW9MXodfP
nA9EgaQm4qI09+bVQFefWX3ToqApKQLE8e5ZwQHyRjIwp0CEMtWOMGBefGFb4Hac
ZtI52iX+eBqDpbQU5tNCvXBPP3wiXqmiq1wiKoDz7dCUjlkfIpHh9kBuX9ZE6ObG
CA0Wv+ZZd9ZkomDChuTlyKm2j5RC370ub6Yv5q82MSU27Prs3tKeDtMU2jpXayUU
Ubh5m834SfBSTCDYvpN0+3tYjYNJlQ6zIUzjNp0iAFHq57K3bA7EPRSxMpnV/Ixb
afhBEIybZUVaIZiTZCJqVdfJoBMmBcb1LvHI6a9IvzDYevQxfK7oBuhV3ENSfXUp
zD0kkMOPXA4/hvDTgnQKbCseRe/PKdu8XT6YI9CMZBVS7fa+cOSAadphUourUWBW
z7jg1YJxmmt/AeZ89weV24l9kA4HOghKvaMglJC03m14reJIYb+pnkB5qHOS4vcl
xgyTslDrSZqQsgD6xVAfaHYzUxmJ4xGpTQOESRE6R7+QUMMy/4uqLBg7gcdzHtSD
0KY5nIapLq6KjoxOcXHBHryTqyCuA1298x3qHd8W/EL+3fxDdPkQgt/d7VtnkSfJ
PKIUFufHgOBp91biqhb8m7ywCCqsGOeACHq8jUAiH+1SNgXObT00wCtPdjRHOKyq
NiLR9vSvGlkMZ7oYBg7xHQ==
`protect END_PROTECTED
