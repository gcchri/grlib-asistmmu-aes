`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1fr5AqdM29PmPzX74E7AMdTtf1dhxHiSXZcCclb6Qw6juV+/uibxZBvUSnzzTKaB
2Oi6TWWfKAX6Lng6gvMseG2cjZUwu0QL4I9Dw1EscL+e4p4s2KMV2Sr4QtXLxJ1u
ICQ2zsf/UJ1vJhFNG0Ul/zfg+11RLH9HnNYwinaqQc8IMBwhSwpPmsNITzBTyjpp
DE6VB7c0LigttE2yQiuB82T5tKmth/BL+lTFRnQVWoWyD/aEkLaTMuwQ5oTisJck
VXvwZ7Ffq7MI5ZnLLA7y6sU4Q9+kyb9PUgTTlyIrlXFhL2n8X7r7sZVSCQuMXDKw
xYhaDVB1rbFuyY1SftJkYBGtJvcQWpOfus8BXcVzr77uGrZXd4v80PLNAqPB3c/x
S6HlveJYVgKKuvv3cSb15Gbn0stOjUYeEkEi9KU+i+wy5Jm8FToGSG/BKMfwxD8/
AbWWkSPLrH7pbyXS7cYq9kuwuQu+ei1dRepI9gCN+ddCb3RZGGlKc9ldtN+y9Ic8
nPZabhnXULlUyiaoflIIAPr8Rpti3mkWuNrhblHDCD4uU4hZYdmaxI0ewW3ag+hm
/3oNM6KtipCU5RuxrHUJPIAoOspBefIARn+yA/vFzRl7ELTiqzgwUjeqB7K/6dIR
mSRuJfngnnnRON34wXB+800QdZQKdtX7p5dEoMN3o9mckgXyja8RhoRSklcsUket
m82qe2dM2Nf9N4PONe5WvZjadFUJS1JPk5GmXT/u9jAkNJHmshhiwsQPOewzBEPf
b+tpU7WAQVuxXuHzrKN/GWAv23K6gdLQx3tvb+6/F+QgoyNkHws2JG5qT5wq70Hy
rIEWdsK8bPCEbtrCCXfAFbpE/UZbxFNzJgHyntpWB8X0hWHtcMfygVs8m/2/QMIt
mhUVcaz01GZfuhTtxKWS0kQy07sMQ9gA8Sf8Y/OaEYi/0no5XxcVEiPtgBSlol+Z
yueGawzf9l244uVVQqhK157sCrVCiwWBtYvn9PqIU6oURlNjLqlHVh6IL/OJ8tpB
rfjM5bwCAPZ3PSSSuzEIIw/o3av3i0KytUS0U+Bfp9Fbo5r6niXk6znV5MLnis2b
3BtkRcbbmUTqc4aLYFDNs+mhw7DCNaQ7jddwBF3buGqWN2SA1VocmGIsh73pjSnb
Mwd4th/8lU/ViJaMBIPNf0AA3+Itc1Cv0lccmdqiu9xkt/mbffXnZ7Bez//oO+LO
S7YZ9W9OwKDqlffJ/IYhz08GIiKQlK3ANw1q39IAO3v/oWMHSlpFAxL5mj0/BKmU
moVhftkzThDILoZY5Sxg99T56jfaa+09uXPXVK+PjKjQEV5SY0749Dt3lVtqWVM9
`protect END_PROTECTED
