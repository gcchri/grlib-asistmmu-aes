`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H7BX+eBSxUimWqo73eZD+rR8P8OZknWJotBy70Q6on8mztPhNJT5cXhg5Yy0tgB8
1ER3ZM33IeFfzXuk1hBbvBnnw8B25JjGkm41luI/bzAmNlCKRajIEpBaat9o4tPd
JDhNi0Ql/Ga8u6ea9IlITImpQSdo6pQSj1bz+TwAn18PlhE7FlLoSY7P8NGXnYwh
m+Jbd4qMdAHw8wn5qXlbuBADGJzfxJDJiBKPz07GQvpFcC/5QmRLQGYLW7RfhEFl
Rskc7gM21zOmwrokAVccAEEyTgK4LSv8+79qir0nEw4tJVIBYR5sJbbj9D5YN8pC
MudU0eh3Gn7gP9ho4oBI57XHFWPpw4f8Yc8yB1zGpaxWmkArTu/47ypuJmUh0dW4
V0x7fd9HTbhbvdEOSPmt0kwiZ/LMPj2ct6cXDum8QzJNFHGIJj9beYqmOiuHGgCo
`protect END_PROTECTED
