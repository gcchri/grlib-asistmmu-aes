`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZN8V2DgFtqz9+3KMoYvHRppHroWoxyxeGSuyKoBrJgcTSVA5cIcTpQTL3CmIetvI
M0gcWax3HnTJBEA0n05A2tGtj/05TzFj9bfnUhuDFrzowoaB0MCEjoJIf6wKRC4W
pWRsPnFSQOCIt2F3x/I+d0T8GEHR7UroMIbIzk6QLEeXSjRaxvjpeRvmbyzjDWAT
m9UtdXzFV4odRnU4hH+R1WLW9tZqySyLxjC/JZprGiXgYPX+0mgG7sQfmOeSkUfs
DFduX2ov92A1cbgNO+XsvPbrbiQuOquWGx32j+gHfoiSqvTN3BTIMkwE6+0oURTB
`protect END_PROTECTED
