`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DCbp7Y60ckNxpHtSbC0MDdhP2LFotIhmNH0iMDVqR5EpomxpjoiGzNuqRU3yaDrs
Pk0WqyYFDZxYhUZh6FLBS8SNg+6edYrWw2GzkWZAPJH7/ccB4R/uoBXl7M+kz7Oq
WXfGrMd0TrSv5h8dRjiHpDtX/VvIDnXOQ/AgrRPm+l0Yn3MrrpeNhk6oYxQwHiLh
bjF8ZrRcqe12q8g3sGpXHDA9rEPvJtOJNRqBQlQMVpoM/CXJi9KnbirKT5nIddA/
hVCOT2aULsz68KTlLiK0OA==
`protect END_PROTECTED
