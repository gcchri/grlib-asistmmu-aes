`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O59caidJ5SUQ9uEYdT8QR2TKgDe4rCNbSYaMPeyGdiYb7Ibppxr8taw47aN8kcvS
B3LDBSi5NKJH4fuBUmL8OXTXKR9vHl6V7And+41qhfRabInSpC8RP2lKgCA1/eiU
zni/5k+xLDaEtgKewva8Iunu3mrAriCrw4dIj4EScB2QaEsgBEmOtTf1qq7i5Bnh
7EKMlZqydesQIhwoog4/3YM5Iw+Mt38w46Zks2QY7uvb05eiP0undLJ1Z4/jkRih
sIsZlxe3rQAS/LsOdyoAQxsJG8/VtwLWQ189GBBAp048ZrYcHQUwMG6nwFd/rNqP
KodYoUBQWgLYn5szWtxghlr+9Ed8HszuNb5Pcwt+xnjtlKija/q5bX6jhB9+mdxJ
kugmPVP9++ThI/BwEKdy2WHTP1R4/xkmbwO4OLmOJ9pWV+P4YeD4msjHX5Lzjm5G
Qdj+H3HYUpP5DRxMUA6H20EUeVSHzIovJDHunDdqc+1uGzHiaBU4gVm3C3QIkDAe
eOoFssVetYK9CHAgYaEyr4flwe1ufyrjG33EWH8Vs1ev5x3LFpI86jl9CuPqlKIo
z3r6CHWqZKes21bRFK2zU2HCVBX4f/4m5j4vesXIRhbyiNQE9+mN1jBWMOIR8LV8
Aixv0N61N7rWfhnCtIM3vq8NFn7FUDrtVSOzzwOWzVCCmrgEhW9IhTptnpbPIwcW
fBCk6lxOS3e26gZD///VODGS049xbLSjKmngFcRVlYs=
`protect END_PROTECTED
