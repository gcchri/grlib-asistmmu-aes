`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wwx3dXbBtmHX6Wvhv2tH4rF+cbQi62WFA6ffOmtJHvF14EAOZA06fdEEyXdlshZH
f3cFvs/N7kEHE6Gwm3fzAbmrBkgmUD5e+AtEIY/K4kSNtbvKwfGwbLtYlKo6a1Vb
1mXiZ4aF8m2rEfv1mruoSFSFVziuWi5mn0rzNALr52tg65DyCxwZVrdcJtim3c+F
8hsu+pNJXdspmoflZR2l6u2X1MMI7ryy2nola2Cnsy4PWuLkYht7oNyWAo332UbP
B7Uhe+IlyHMiEBGyEEIMjIjRHZfBfZ8LIoKuoDWCNmPD6U8f1GzQUHbPbAL/28xK
NKBwadFpKgpX20iVh5oix7r3Wsih+gXerDYZu18V/PjlR4/zdb7UecB2+tzDbMKo
jVOp85ozKxA8f4P+UckpEaXY6H5cLYSImHzVpPx8cvMq1mtUsDyS27Lee8RB4iHP
nwENDBLRH+39DL4LxKAYhLGgt34DDirmDByHMemfSLJPho5YOmSi9e1sPRQk21Wl
PIMnGbiME9+JziKbdRhRwppVVmWoXc2+Jq6+FQxa3ICdnsuzptLXIYpJVo3VnlrO
ZPeF4qxEvZSGulNKR+LKJnaZvai/XWuITNFlCqFFxpPLYZbQeBQq2hjCpX0bVk+e
D+8dA6QHXhN0FtnD0fQRNinrv1TBokAmc9/8qdbZd6NHIX5f3KZTHf6JxG9brLz7
FdV9Q0j2V7FBhdyG+DDiIF/6p45VjnyTRhUbtvTqs9p8HAN/KyJLM8Zaq/SAh99o
2Kuf0386jzDEz+1tyTJaMQq5TdzLie0XE+EJOcaHX8LlcQFTKcuv4mL9TVf1QvIe
HYZq8BYQhVhe1k//4dnCDtgJH0Rd7+No11TwDEHKA2JUOcWq0S2ycqatQgS7UwKr
F3uyPv8CffrdbIiFLWNrLQqbEPl4iT0U/6pnAi+2IF9sKMaCz6ldURQ2UMOPUQQt
NGURxDu6ajv263PvS1W1RBYI9FlWALIUC1p+CTgWszI=
`protect END_PROTECTED
