`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FJFmt4/Oykmz/KLk25YN4CpT0QmZPjZ6bGc0AUh5c72+XSckKTwAwEKPwXHk4x/d
f5uGeixk/nY3AuT+1anfySvo6gKsZBUgXpL0mDBbuNpKKYv2v6yelrMTT1S+eFqA
iPDEXu7r9OXAdpOrLTMwkbNv1DpK0ieGphapdKjUTZGnjJP/3zqDHtUY/IlxSHLi
NO4CKpwYtf6+VVuf2DzF3SB/YbBoUj1jIZL4Xx68tpGY/JgB06c9CMzWJyraLKje
MLks1uLPdjIxY6Z90BbHK9DJXi724xtTMkZa2dxHe7zflOH0w12og7dYtpe30Afw
06YeTHkaL3/uwaxBw535qppGepSQHj3YhvP2E2BgIyion9W2wuYJVZMccQXw7J63
+7JkOJq1AdQA4p7nSbj8eUbu/4c+Tr0Lll4DNaV1HoaJ1T1Uf/UhlwICc5mdC2PC
xj2Zwh04rit6hcsHKOgQsJ5TCRWNzK2MZd2wYcmLpUf92QBtPfSvW6RDKoqzknjQ
CtcVG2qgkWX/Z9x2Ku5fWtsIF386WbUhJ7knzc3E9yOozOS7shMksrJIUgThptKk
xETHzTHWqFt5kKP6rQ413TC4rwhX+CVDkQcR1SaWzmWmO2kDU86suKJ+oPUwdpAT
OULSbhxLQNOEEViiUGxsQOqBfBfvEqtdDk+VoQ36rJUQBZDkRZDpQ3nDg/J/Fdr+
FS9uYf9iaDj0M7VlOF9VSzBb6QHbz8vpEtr7vYnOe9a9uV1omvoaFROZDpIcI2W3
kBlngqrpT/QHF/CzJho6IR3E1m7Bz2SnUtMJgSEN6YksKXXH8FkKsSx1uzkA2OLq
VCVl+hyIfHEtfOF4mb4JVJi0o4hIRX15DaTuyi7FXfOx1Db6cFCs+AJWr2egWCi5
OpLKfd0rtC3mQHXaEathqObcEUY21v/9o+XR4DbCAPDum3hTX+NXz+UM/6pOGPXv
wpuwaInCZHs+S31ocN8pTWIacZR9WH8tBxWFQ/Qe3bSB9bqNy/X0Os5E0UNUAy1x
aaHFNRGkWzrdhP46C2XX98eCfcg4fnItr6nEixEOb2cshrYI8QdyRpm6MNbefe/d
U6QJQcKNqkTYaTAih3PCx3F+q0oV2aapRHwM8MBiHaj0o6KMS2NXvyQZOdT68zhv
VEIkAf7NLmrdBZaSFVYQWY7aRN0i+kUyvaP3Hail+ApMpIlLxPFjivLWDuF82XKj
mHUdwFg3p/1LhGMwfOSwC4YOesj4BxFhQrzh7QMljaJwc0kkJF7NyWK5BWAJsufc
gBpsF5r3MiJAJSASqjmdIAgx9nhUcHD/Zy9rfeq9nnWiFfm2aNi1hE5zyoTMycAK
2G3F9T2qM7cEuMWIGr2itvQ7QEXUOPZDiI44z4XvbGyXXomdwOmjnZYbx1e3xA5w
A2DLAqXL98e/VR1UJ6ajFfifM8Omsz/K3Mz5at4bk+gC98/UABJOufXognPA8Pb2
/pdX1B/9Ryafq388gYlxiFAUP0bP4FU3CnZOx7wqpJuyQyMSd/+5L2CRQSOXzbUJ
cWxEoHtDG+NscFBIxgSfaYRdjAtz1C+xHNsnEBk9V2l75tEPzLPbMyOWBoXppJ9Y
J0Zd3kk9xxanaz3kmT2wLhPNMA7gFPm1q3/EPb4qQs2633wlZvkzVlVPFUn5bf8J
Oi21IzuAwQc5Wrl5QHOP0JMLYheqmVW9kZNOKOxcz4ULmWVfegxzentPX0ytHjIh
Y9d7OtuK1e8jNURn6GbZ8K6TlvHJbYn4aK86hksSU2FLszKWZjFhVnjYnk3AafWG
BqMQZo9/yiTyn4EeDF6sT8XhpWJimeLQkCvC5kgxks2e2zA8Jo9P+O4Qc3KI72CA
oEFeXbtVGGDbX4ijSn6Z/l2lWaBMDXUUXIocVfGLFj1e7W/OiToY1Gbll1nzEcju
QlyDov4ZcPJNDhzSY+0Jyhjy1AhekmwY70EFEQC+kNEbMXsJdrRIwX+7STswRec8
znbYb5Zv8tZSRUTnVtHhhGnKE/72GVbIA5SNqIL91k6fd6T5VYtPrwGU60UoZEvL
SSmrX61+ENU0dTAJyWXQdmEX2977hDRpYDn6fgyEfbp5htnpU57w3AO5ILE+WsZ7
vFY0evP/8nAQ/3GIT+ZjFXZSIm75ymD/mquevLyCXkTkD7yYASQYd28vOtOFdiVP
E3trQTNBUyIVoWg0eKk7e5S/Crrq3DUQ93/R7tIcPtXyc00e/ttXqQnC9Dpv3CKQ
TxjBSFwx5vMa+gUpWV3nk9w48KFze8WwRVqvNLl0+BPuGiMaKW0qdsY0UKsNftn/
vKGZvOz4tls44Xk+rXmT9ZriZ70KuczvYybZGyLyrm/+4ZU4JAorHLwDGGO+U9hl
pqgCPNBw5XJ9uHy1L7z20WgT+VtIMhCSOne3knshPTCBdShK2E+S7C2Ae5Z5Okrk
pCpYSkJtoxlBnh8LlIP8F3w/1I7LefCieqPkGFa/BcssHNHVGyitE5IZAu9LF6xc
3b8/k4Vr6nMtGw/oFCXDBuN+eG9dyt5WA2Lia08GZPE=
`protect END_PROTECTED
