`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tuoFUWaSi7lPrw+6BDJXMJFekK+59hgMUHsumAeRg3fnL7Tg/VmS6gswMhtTQRhr
Dg8BUMOiUo5lsvVw2MQUQZ7GcYqRvu9Htofr2HhnwyW0FzS2oZxvL3Mn8yXPPgux
TRxI+qg6IvoCfa/7iyz4KzIL2wIrPFDxWXYd279vFI5SuNtb8JN9eL9qbLAVROPf
7VgckZfNf7elrNGDTISa/TOic8YErr+1dkmKCU+ctP7fY7TdDIv0qEhZbvJBh2Xd
/0iWkh1xrZZJaTwoxvB81Y48JJoJRix5uvlHvkLHRLlQ9+omJT99suglZR67/URo
iFNs8uXhX64HUwpedQkSvqtH+94lAsdfhkGW9H9KlDHJbBFQvjWRRMT3ikZ+fbsh
g8NOEENDtzJ6e6QMMfSpL93AWdF8UenxGedG5YpWmlffpOssp8pPLBHIWtOx73bd
`protect END_PROTECTED
