`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NK4zhR8PhcUbAPdiJHb+0AhsDjrbQ7F6TNsoYjmGi13QzOHWpV0HAExMZln1ZgvW
/qKvT8ZfxXJC3297/rgK90kVKbm7WhHP5AGCULgMDYp/69SyrF5BxefcwzWp78Ve
aFOIkHKZVQRzyo972ulXui3J0dtgT+GlBojswJ17P33N7T863Ru7s4I+IHVDqyq5
xJBc5xfuawLdARGATbRQPevu3GKyfoGAjs90H/dnO+pjoKjLGhZUP9v7IxDvv80J
yDBLNeLRFmkLDuPHtDWcqlt3nL8aV+j4yd5kmSRYCD7B0xMNGIRp9qXz4TjJ+5Fi
igUl7UCvpUhK5T7d8koRF3VZZsvMd0mxrflh/oB5SfC8OfGzxynIivIGVfnxolmv
+NZ7fTC568MXDcLeeAsMuGT0nEBJwqJ7eCa4DZKQ1sTyZUXIenbs4ezgVmToPxL/
4MOAp7FkKWtmfLKWSPg9km3AQNK0VmXh+GMij3mwMJ9Kr7DgFlynAg3fMhnIj/6j
7rqappEPW03v/Psunlmegb6Zr/onmgG7Ge7pdbQdFP8rZC7cEU9UoKGd43XNwpiz
SWwFySWEdyiLqpFoe4yHKuMK9xp8dzBUUYw6NpJMSVyaoOPLVN3gUJgPyVMTC1az
+K9CdXo6UGVlM/z2pj7+8uKn6jXbgUaEgX4iBvDnk+jZwWdf58qjXA0aeFPHpwpu
uiKRiKEUNjS+sfNMX+iQxLFQ+Rznsktbv4NV0v8ablrHQ4GpaXM0nMypRAsrc1fs
WSfSDVF0Si369oCeUVFGvL6qkc14z2cmwq0Y//YbuGPYmg42QMRJ5bwbwKU9o6F8
IvwYS8gykrfSgx0dbtCp11i9cs08f6AV9s3RZ4kFqr5ZzxfB/oNOc951ZqVV5N6j
YPps3X1U1SnEAex3d+AsWJiK1UgZ2tTVJYQtmfyzLLIoKwOrAsZ1m6JP6Io8yMTm
7iHWRFh5ZNJKpc6L/NABVmUJ9ULT0flcaEEPWVmHdgwOMjSTOTkuKVuc0XiIh1a+
`protect END_PROTECTED
