`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+rKeTXiCkU+7fwXhathAbIlPfwKobASUMHSdA+ii7XVYX25JOIQCzGtUvlDyRNZ8
l+j5uGNgWatv7pnUWmlqK5eli0J2l3B7AbJjCre+hxW8gVcfgOcRvophcwEnB5/6
rLH9smMJefZZq6JGhHtPa6C+sMcYIynF02yPKgojHpBpUBY7c0FZTeii259QVrUr
9IZZbnXWVIrQcrsbgAoTrMOPTfm460DhwahDWPt5ZyXyecD/pKW/fLIeDtzu+Bon
vtxfJ7nksmc6TySLB5C6zdqAzOIrq2p0hhOJEnAIuI2wUGZnRdu3axhI0yPLvbq5
ErkcmxIthcVN9pPGjs7RZZS+oIw5i6qYx0/JPTe9v/395VpR5sgHolYz348vq83N
VgncFHwAy/lOUY45NPGov0zvErLzFbskkEsi46nyBsU=
`protect END_PROTECTED
