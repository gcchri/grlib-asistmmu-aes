`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xf4OZxi4TqqFf17vOrp1UPjCWxO1CteqX9guCxjkBlQX9BDHvZrR+THpAquEAFgt
aiLA6KdMIjqfDY9hVrHjiRoTcicBrQSN/Q90MzhM+7pcgho/qkjwas+xaPc2YRn2
MeBh7b6GK+BmK6K+FRy8E02pH3/dRVmW4z/yVKcnChDaGeIJ+OlBbHlo9aV+XIdc
la/M3AzEV4xtQX2C0X6WUGfjs0Jv48088RDSSZkhWDlwyGtDlEaUrjelhgIeP77e
RlMEt1Cx78LidaqIqNXiVfIBErjlqqt3RAdwSfbIFbiXx+yefjPrVobKCbBG9G3m
EWJ4kNnoQS847chM8qaL5lHvqIPbn/vMn2nOgXKqEk7jMEErRC+xWKwG9X9vyCUm
Zz31HWhW+wrLrzkd2xrxYjYLiHNeL1dDSxuDMfaeyR/f8BK0Y6/unyIiII5u/ijc
`protect END_PROTECTED
