`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z9HILNJ3L2iRt9lIF0u13e1QkCX3XC631vtnzbcZu1/aqUBRTHoS0+c+Y5Z6HrqW
Q0aPBN8oXnU8lGuUpkesX8Ialez/5oAozIDzXJTxH7vCNPodQc4IAy49ZBXl98io
dW5b00NHb8KS/CnzTb1KQQQJeqc9hMqVTfwNp4hJbO3WndpcZYeBojhB7ZIT6eUL
yI8A8JOSY47LUy6A08pAj2GCyJK7nILoSSyTRsDmJO9d6mD12nJ/bWUNeDa862uk
7vWOlfi3fjzf+J7iCIxqTQ8hQWouggSPbqRCQXpQ6AFcsFtPn1YxMjE8fLelsb05
UnaVeCFsKO40362gLwkuXTIi9low8z6QEPOMWlUrQFwTpbNlE5UXqoEXApcsA3G1
kFgneMhBGbDpdsURgLWX3U782bKAH1aM5v5qoAf6GSXyx3St9KXaRslwFFYTOW+3
RCLiTxFK2551vNrSb4RYK3Qh6xHRCgSo5Ebvigz2OeVY37KqY2j5o6gpWX+hqF8T
oPOUykDrGdZJlTGhemKOXKcoeqHBVv3cIzUh2zAkV8nKyOoLsDVBjzo1iVMaGnkY
qjwhjTmXVlIpTidFiqZmIZZl0+eiFG+dSUA5hYGw3Osc7wQuOKUZiWdzKirh4ZTt
LNJectrQfkDSkGOM7ef88umX+FUVrLv3pzreTxJ9qpemPwx4eD+GwR4ySlr3lqse
WuVF4ZfEkfSXbc9Xqhks2ntyqxWFD/gHJHwAHSIUHpUXGO0FxZK/7muxUlTSL6NR
NMDwIvUC1H6wyOG+YaLJVpFQjZp3z2qVhfl/xdqIDUhPIq4mCxUSc3bAmBQSMLZN
AalIpI0wOMgZy7WjawFOUIRQJMjKKKTeNzO4S9QdslTmRaM/zsenfoeZJQeM9EBK
aswBH1bqYeGYE9gszsQg1NuEVNNF0lel4VN+kORIl0QR+qI9j0xcUBHAGSSkMYaW
lm+Ahf+MDcqG9wh7Lkg95p0LKrYVMhIgkc1IfL6or3xS3pyVcdie3/llwHi5GwiZ
Hne71ccmkPu3HagyhQiZSb+XDWRiwQ4I9kNA3wfVaHYxTsJxqqfLwnF6wdJxd3KD
ShP4anC6QrGdXj0RtopHWOTItIzeUVHT2ZNueVpliSfruOsg9cU/bkVWqUH2yzJm
IlZ9ay7HNLz2rg4gyYo4JXuEmVqFClAdU95RsLk0rlYdVFZX2Vfsuz8lJeyn/02o
W2jM7Tc4xxab5x+sUkVID2193T9di9/MGRw0/9RR9NbGh0MigOyaqjEcj46VJ9IU
uRyD54VDG9euXxjw0lrVKhQUlG6486y14dZUTQ28zjPFOtNXD7/WrF//RGG+QKcY
B6iZRAFx7fi0EchVT33YiLph0GQxs1ko4EYttm6Ed9RiB3d2bbUiV6/fqX3ioa0s
vTOv/zwc0hYCfx8OS/Fyb65pRthiG1vhL+eoDezTVP0xqT7HIqgz7pJXP0vyYOn2
cj3AH08glWLUfxJpgaiTYjrG4KEnJg4Aqy0SDHcC7HrMYK0FJMKeFGXM5aeejHsu
f7QwcmWj6TOD3vAl/vRqADJrfaInPZc6q0ZKDSWOBuiQ+aviNZvNlxJs/8THnokd
dFMeqidNxu5bhDlC2fs/0uSrkI6U54kKIEoqfovlKAP9TtYVvX5AVcrsKleBObCK
HlVBB+oTHX8kGWp4d/R8GLKJj308rCCBj6N9P3KXSSJQKZEpUQWdEoUik1dFOgF/
IqLoj2BVgJ+Ijtrjv9PVNUmXn/Yc+CO17moJ+qJYWbEq+MluTLLl4geJg0Ee3jRT
RXkCAwOJi5DckrLnpP5j0KRYZxxxZTZz1prFY7B2U4KkQHNAY5DM+9GDi/Ut+utB
FH4pd22z9HGE+rSUFoZiSr3TuFchz2Pp2Zg/ZJSw3ejrM3NbfAW0AUqRsWRRpR4l
lDjfIw0SNEwXN8UDUbjLPIJGVMopvl1SQeKLz0TiDxs1JvfKUsUyZ043Cc7Sm/Dt
iLJ7qV01pCEsj9jbAge9CF3eMTnMaPx+SUNDEPzc6ewaZUXGVqkrsZ0Umv70eQfD
EceaAjfua1CiQZfeMLpwXqGJhTnlyxL9zHafLZ+TXA3sZjKCyEk0Ln478BOsqkXY
uFVvor2oBLZQvHUTQyUeUe5OB4SnJZd7nLovkE96BmDDeuCeIxBWc4iDxAaY5G5Y
DG3Db6GnTnyoenv1fQjQIMHg28oODqMGGdZ8Ese0OGA9LxY8amcTF77GXYT2zqOy
uEOkiFn1nVBZtG7yPL0C085u+N0wdw7Ony0o2WjkGLwnJyWxT9XBgNDIX/2j48n8
1SW3MfTbF6flrlFJvWR9MY+L5g25Ukkl61omIQUX+02PsE1AXo+Q4PlX7cwTJw5R
8ZrD5oYcc2SX03f4TZq10JMXjP5xHo2sJOkak+wBCmzw2NhZbcj+uY8GmZEnTgqj
3Hy5Qua12lacnn+hoBM4sK5BiTqriTBDP0V23qMj1kc=
`protect END_PROTECTED
