`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W++9WPm4eo8oG5xLQNKPCVJVRm/ko+x8GyYa7UfCvrn1893i3wUdfsSdRNHHuXgB
XCgsRWTP1UXB+l/E41uGcZfbtJjlRgHRZ8fjxCTqa8kqzuVhW1/3B+1cp39PeNQ2
BgugLwfzcv0bLuHcp41xOniTrUUy2gFzCn34RdThCdFlhMAaHxMqL4bZhkXcNZF2
3zAx2cSyLb9C4hnaOlmF91SfYDN6lIAn+6KWkkartYLDni6VdDtIElx7MiooLBSJ
nesBJZV3uirhK6h5F5buqO54VRUHxGxjVdkd0NXyMVCARS7smBMnNxRVsdCRE32D
30d1+r/ewqXzGnPQdBu75V3p2YjqHOcg5ZXyeWwQy+XWqw3GEdOHHWQ5UMIRdyD5
SYjZ2nmKJSu/xexYCRteFWjyZKPcFVm5NiVq67DtFbSuX/lH/RXVEYlMcZaqP0fb
BNDn6HpfQw8+cfvvamzITwjmK/ivxTTeOwMYdxNS8w05+AJ2gsdAfP8YDLN4q3Ep
`protect END_PROTECTED
