`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
36ZxuQeXQtL5zsqlt8Pxdqz0NrL6g3gYOTA/XrTc7xqqNQ3l8695yOMv6mjeEDMo
Mf9MYRIg29qPv+xk51UrXgNN9zCCJZxJLUotpuH4sqzfqXTyWL9N0xzK7P5n3vtU
c8agqH6QLvwZnDdXhpGgG2wjwqF+TzWuAGrKk6p7ofjo2jqwxhILSCtk0AZRkJ6Z
ZI5JwE6RITh3wPx5hVMlqY86FihPn/r09nPAV4cw9Lk5lCpPlsf1PDYZOuUAMmUc
fBQCsK0RNP22MR6bESt+ZB8G4ZjFvGCk4vgZ5R2zIPowKG4bWAIjxsBkt1S0ezvI
bD0yN9db2i+AAYuLi80j/Zgy4GzbcSnlMAPGNc64fUIy9IkZFqO364ccWtYS5yqL
QhgZ+mIm951AKF+q9E9E0K5cBZAnE8RUR0TuO3TSovvBVASnMH8v57Dx1KkuBkjN
pPxPQxc4MjGhMykJxHiJqUR+MOKxPULghyMMyXL5CIoWM/XbcQmSqkJRx/7ChUr3
a1pLdQdYxf1itp7hz0sT4bmB4SgA5tlRsUGPgzoOwU5xL6dtQkBSxTKTFXSU/kX6
8hdyN8h60R28gDpsZ5bGqEpFX33LqpRAf/S0Az0/131udKpVAZ0hXJ6+scZN7yfo
dNkQIAwJ55lSGFLzi3OdrXP36yhl1Aq86Qg3s5axH3PV7hZyo7EijRcn2YPGTvJt
kIXl0sNCTXVY4G3FbQWSnj77NfbcI2VmN1nBKZGiONwzNlDbDQ1PdsoSp7d8Lvuv
8AXIIZHenB0Kr7RPhMcl4l4U+1AgYY5O9+IFnVltSRLBHowcIbTGb9VDifIkA0sn
nZNMJRFQpt5CP+beMrWitN3lv0vJjG2kWvsAWUaLdknOUHGWTVacS90EAxnay05w
QH6Gatd723YnSdNrM3+QKaU+GxnX/pmIXM+F4IU6m8FBYaWNWU5wFcVdoHlPXk5F
BTW38J29MUlBzVXrxdxnzbXMcCc2O3LK5GOF22CLR2in4T639QwPtuPxCG8dqcWm
IMLQfwM+Q5AfDj+WRpR3Tam7bZphE+nhfBkh73smLK3E64+8SS29WNjtRX2EUM6w
CAZCFGsFfhHD1c5JXugEfSFupscYkW6vCSk411Qz9vk22vO1oO6ibNF4d3Hg9OXf
/v0Hk5IXGtewg0uoGWbp0tjNe3zviGgu7SO5oDfhNSlanV09i+7BCOCRvFwIGDfW
nSHlVWbwNUemZYYUiPCOEE/N51vsnEee3smL6xyRbLPNHh10ibjt60Ona65Rp3BO
liOnD8BH+ojQvt3Bc5yTEG4JHIRHZR/do7IMm9IW5BEbhHiIg1vnbVUivPSg9azs
UCFi96yi+PY1W+wdKFB/ijDLWOGPrJHhYo8BaVipzygcmWaceDLU6fj2uvej7lx3
/9X9JDlWjsg/J53oiM0jwxE8mXW2iFGB1D6ev/TgBiAfkTmIZa276m/EI++fsddo
97FFvAHFq0+C0eVjr0RwPSxRt2+cPHfsyGo1t8z8nGpWatc6YD8xwdiSZTRhw13c
WVCRWGBWCoJm9tA3Xn8Nh/hUZ8XYo4Zs+jiCDKngpicWDaz2FdjORmofaFynuMFL
QbVoq79ma8IgzyEBJe7pc0yi+ChODXx7TlGfNWsQ+VHg/U2agxtGfDwEldBwueQa
IfZo3i3NkS9inh/CfSlNIu51YGITlGM3qBCHO4YMjhoQIa3s+23D6uDertIGfuUk
n7bv3f/fc0RVUtj1+NGwc+2F66zC8+d8vt+OiDnkOiv327QakG5yXzTY6QWbCBEA
D8g4UpmvjFNwGzdmlHj6/Ezy1fwDouqPquVVhR6ioEH7uhF+17bFfKzEdY0A9uq6
zNxFMAFDftIQwqOdoXwne5KSDZFiI+aZnrjPKDFlaLMrlS1M6k+sUBQWSe9CiNQ4
KGlJN2WOSDoa6IuDru5dvgioUDLT3O/grGiMtyeAuu9iPvrFd9UU/STw3vdJnw/b
LgJ57RoZm16c9sSEImnH8UeShl5uBgYpXL+uHaKg5NPVT9Ah8Z1BqeCUQWRZcwot
9Bk8RBwgxDBVjDQ4AObJPyzQxD1OSylfvRb9fR+vjvdR2+DwDxYeuWU7gJLrofyF
qLNvKkDdBPrUwXkW42mldIHep/ZkRMVTdIOyJK/acda1X1AsBm2eQ8FuCci4EnNo
d/rYZJjTWXp1CpO98KQSDLThjvH/WiGsG3Q4+55ohgg2/xWpDFXeeEDAi7JyR6HS
/bHOm++MNwBPwzproqiU12LaKifTbeRl0lwbVginVjD5d+hZHeeJUi5YpcWwYx5G
YWpMc6tKfeuiBQlYg1J/rm2iTB9PP2zeEw/Ch+jQgHQCMpY5KVQR2H/uUWgULatV
Apx8R+7b0fXg1Zt0r1J921JU4CcL/j+s3wtwbb6WlvTpme60DmkUSXo9QclUMalW
pFwnFtEJXpCm6lYBBub8tIwDffUL5jNmmG6bXsg/Vxkv0AUpW0VFmUv/2eJurORK
16dUTyO/i9+VWVfJAiMDqbDo0rfThXE2dDKYIF9kCHIieYpHjQxtkGv906iPvQ2w
zaoHPuRQtRs9x87wwATZDAa/S+m4cDEbjSiEhBlNxztMGy4e6HpUU1++n2B3l8fr
GbjCpwyMpLDKc2mpZ1PKpDlZoS1YvhNbf/VUH+kdbSUlV5YqPvdkaPFQCzKrjqDF
35K0RFtYNDAYXDDBc5b+FLrfwooAmtYMqM+EYzp/09MQTi9yRkJQKK7Bagpg61R8
KKkJxYROEVA66S3jDle7Rsf3kdvpmOqO6y8GPorduHhVVwFjkW6dx7eFqJMk96bb
3mSN20nJR00EN1tfrx3fiBNZfgwTj4btj5hUs+Pn/TsKJ0sA1l7+0qsmVZ9VimUn
Mv+Jtrbl1f2xpGrNps+W0UV9kVcm4/WZE7iVzdzlZ+a2EhfFdhFVhZDzBPZhzr7C
1CmVJR2FUWu/uABb4uulJD6tGvKPy4xG2VOylI6jh/DXTiB2c1KV4G6AD7YZHA+y
6a2iH39/V8E2ExxPcPwg8zS3phNavhGQ6Zd3eKP9gCdjWcfewTP4oh4Rv7gyoEcv
JUpvnetrZykuW7BaMAu1F1NoyUl+WATW0+hAnQOgUiKImH/x4+VQg7FxSJulFVBf
HoMFbQ4NADl979N6chCFcxU9mjt3rq11e5dzuriooz6hb1J0Li73YJ2k8vkmxxkT
dhoUBckcbGxJbBowjbfLwPncVS0qinN8aYA4jhqzHIDkncXikB0+wveUenKSM9WJ
QJGIEug35d2+FJ0NU4EWAU8v+dgKVfYad9nldQL3bqrDJFP+Bl+FAYr6tnxsuC01
vnBVwDF9AGNRswXE6QAuwJ/igLY6G80xJ+Vm0rjhproG+JfU/kUVyo0jTcZkxL4T
WetmdViBlY62u7cAA5zkcstCBhhVN6Y1vPK5dacCtCFMEuvzT0xzm0lL7j08ICBZ
IfbBb2/lGFywc7Mdc83DEOWnxpA6GIwDBInyotkI07NJYQhP3NVrX+5TaRA9fDcE
0OU6d4VPbgSW2sC70OxKf5yFA4EW936GkpWo3zODdQ6F50zWHC1O2u+EToncM3wk
pGkTCabg01zjsb2GY0ayvhqQNIj8yNgbgzxWsIkGlTKFth9kPAeYQaiTaL5+tiZU
eAoLcQtSZyh+ATbQ307JTWUHhj4d8HvTFf/697giOV/V5fOWqDk6HyT3tKcw0wRn
9lbSpT/OzZveDk88cUINvUBsjTzBC6hHnkU/5RjJet6tBWkVDbo2LMJrEcsOZYVu
BNZ8WM7vs7zqkxoqUR0FZpXGS4Cv7T8LFXXD+UwRnESVYBF4E34C1gd2tXEtF8sU
8vQtO2LyuUwDc0JoPriex6Dl64oDqffBIehVEXnNPnNd1c0XOkfSJDa1eDsAp+LC
ymCHAyzNsdtku0XDNr1z7flNg7e+dyICLvx1G7sq//KqeH+s4WIIK+NY4661yiCH
ZfmHOZRZGCovNF4MsOEB9K6xO8mwCv7Aj77638RfW8bsqo/ZJtZO5+1Y21OFCnIN
vbIEeUCRdbLs1hTLR5BqmI4nfLID4eflaW9iCJu8nsCyuJC3IhVeXINsC7OQI4vZ
/y0T4bck1D8GLaYYjpFM6QP8Sc7JBPVA3y1A6TdusUuX+jePn6GYJMGVUO1Debe0
`protect END_PROTECTED
