`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i0HTCGJeyoEiKabDByIZ/7SrZgSd7xTvRCjk+bSFTinmdpnnT0BMIUmQAC1h/CD+
joFWj1IacUUIyzoOM59zyK3QsSJzXJTd26zWBxmrl31a3/NkepBtjnDOkxF3entH
7CvQ41R5FUoDCWKZ6ZCuiRZgE937fV5jwxRRF9HobDBJIGiY37CG4M11cSXTBS3S
PgB6zZQe+fT2qeF37Trmdeir/s4TISlpkbuzQtnQfvi5AXT41a4PEiFTHXz2sbLc
WFtJgZkXAIFDupu/uF25IpNH2SwSjWqbv5qVyvP/3/J9r7mykxeyBS6ExoIKTPLX
PTh1L+i2Y2zAYzaGZrD7yFx9bwB3OLbXuMQbDygHZGnRJzjws0VNxET4WnYJStkF
X6rItuZMv3OOTGgL4l66RafzcRKrZwoJ3iR/U+x7oUnddmpg43Lv7veSK4/UNnOj
zYhC8AJcMpaXeIUrEF8IWV+yHIaLiyml+HtMSjp/OGoOfX86jXxxElGMBK128/cu
GAE8kUpffrJWk+euRiCBuIuGGeq6nkYVJZSFozeA0S5iNb6zyshrMZeRi1+j7Meu
krLNCrAr/6u/SZ+EScZ5aur8I+GF7x1n/LMd3l6gQ5j4IYLO1Xu3lW0Hzv9JrNcY
vwL4YRLjutheRWt883W/wH+v6DBc/PvSOK9xSGnWYR82OweMgRrHuEyP6jCJJb2l
vCGUBRpfUXFmT9I5K9jn6A==
`protect END_PROTECTED
