`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bQMqjTBw5qV0oZvXZSNP+Obu7j8RhjBsCypi+C06/z+AMqnw88c9SSn4ZAm3hgfS
jG2vBRle5lzHrWnGE8K4Cd2C48Ol29JKWPpq84f/31WArNeQCiuwmOPLXuIq3nxY
AKceVuWGyJJOAkAxoZCxzqC7N9LnBCQ8dIDOrLe/ufqrPL+eMmCW8930W889qArJ
c6WNMfrL7E65V8x6dZN+qrSJ1ypdKQDu4UlyGov3WbcT7qZThTXcgO8UuDkTOCk5
5mz/ExX7QbbkAWOc6gI30qHo75Jjaxk71yTmeEpwsTMJoiRr+QP/aw0MfDj+xhC/
qK0UrqWLYEEeRquHDfUdtBqMmuTsCoJum4O5JeLKkJ60VXyNcR/BpeBskR3kxcCA
0cfSnt2boupIMgBEAv63EKRoLF+gPpG59B9Ol07opMBuVlksyRVVp4aFw02UfJYV
oo9ubDUENFmxwtr/frbuPNl5MfoFppmeWxqoGto6eeyBTJVIxunb9+1xhhlAz/q9
E/cCeRJLefa82t0XxYCjYiE2F9nUVmbLImxXtT/3ImmlDTh7OMReNW7PJZ2WLW1Y
OHqDckUepg1ZCLWi1T8YdK0np7fhGBUzjZR4ysm0TlLzMcK+5Hul6jKRMAilXKIm
xqqH9Dxl1+TuvqSAsctjFlDbwoBMhgtkJ7uY9zMviBws0D8eXJf2eP4/kuAVuCKq
UnI1fwnpiaqBriHlq5m2+LFk9vAGpO6WKSMqv6qsG8s=
`protect END_PROTECTED
