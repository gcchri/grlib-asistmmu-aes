`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Wb5wohJt/pZ43HfMNxFPcuEaxr8R4ADYZ5yPhxYOiLTt80D8wS7nZR7Dh4JozvP
eIoDhZm53edwJMTYsrmlG2LjOxRM1BADeRybqL/pL/fRv0Zkbdl3olR1lMaKClPx
tpK0Sas63WpwTUXtBQczwpnZtl2+Aw1EMxO+WooNDTXlAF+UEwzMG9w3vNAx8JtH
7FZdoqqMp3z4YRYe8sbDT+yXNcm6rDM+F1x19rohA5Lg4H775TuGlyYyYirPM9qY
YIu9VmBPVrnusPtOGslACXZaVl4IWvDut6rlfsrfmvpGBa6IWKEztzWgwv+jgnmG
6ufPyLEIZ8MLqDDvZOvuj6C9zJ/yFyQXXlaHviCE+swbjr1mTlnoFHb4tBfh4CHw
jnmQBziE13r4bRtUC4C8ed3gf/SwizbPrFPtE2x0czN/MyfQhpQR6NYmST0kbpAK
b5BSityNNlWAL9rKV+mn6k5t+N8NwCzvIdBzh6rJYpA+uXDTHRSbeYww2IXqkJkV
t5utu9fnPwJAOis1ywofnSuizRrOVW2WVB43Ad2wVNvfNV8W40cfA24Zk/KGCZz0
GBlbo92OomdgjqU8e3Cnaj2y4hKgpttENh2qFPaIZqE=
`protect END_PROTECTED
