`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XCbp2dn17Ya9GAiFr5pjMA9znJ2QlbWUQRmHaOgHpscFcgjrS3/Bw2TT4EuZve5+
TWrJHLMsvuHqjoNr+al5MU21FvutpmxZwQj7V0S0vP8avYXKOTWAYaLl+FCv/PC5
ptnJWPQmYzLI6dZ/n9BuYDiMgiX9yuH6qP86eBUX6QjqANLev6Dh4i1s/rJzZesW
FrOQL5pAbU+tLT0tAV8whbJhxBWPXWtUG0+HlG0pYspzusPT/YbHfJ5xCjCwdm4m
gWh1R5GFfmlfo7VYpjRREBG7eSED1dRMuczNNQQB266Ocz6PKT9yXKGq5zVOs8zn
NW6D17YsYUt4jUMF0C1VPVE4aTCwokvPi+LK7JnXm1Y=
`protect END_PROTECTED
