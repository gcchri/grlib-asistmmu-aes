`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xMx5ENj36k1dgUBfr9lIx3GClxNIrxVIt44NTHKNBLWoxgO+jfroQsU39Hw4uybT
vd74/Y9h9xLo+4O7K51uGRXCNSayBqV5/WVAMnS6vN/ObsDdm7ikopG9o6KJcKCg
BauIAShRwX7TCA+AjNkXpBZAgblE0pe4rikhb70ehQA6dVkN6hg6eNeZAM7vETl8
FBmoDSVqHVnrv63NUPwTMjgcuDnghSuHCSKZuPOovSW274xI0ur3Lw71bk3+9QVr
H1uq22ATy6vNMdhcXZgFNCB/2/+LRz+A1Aot8S3B/QKdzx82IVDajbM9jZwYJWP9
4bQsgtzyeuzTeZEHJck1c3Ny32nvRQjunK0AEJklPf7azo8d8Co8oURqbopWbOPy
9uVXhxCTc1wnSPnjmPjEBZN9BNfH8H3Ghc1fqVz9f5/YX/x7CFRq3Jzp2JDcq+/C
Mbn8NO6HM5i9ZSAwbBmb2UjPTl0ZwIwEaq9r87PyUCE/PN2xr2iqhiVBZjCkeCzk
1sO2CcxJZTPt9iDTHCid5SDcNStUfVBNeYk98jiuMmU7xkS/bE/z/RTy5DmvzQtF
uEBUSDzUfGT8hKc/8NAL6IlcELfDAHaqpHUENenhMYPEZt+hFrvYnKHUsofWqhan
d/m/wwEbO9E7X5k9B3FkWdaAzPqTgmdNEjnJ5dJNN974QIv4+nXYYLTgSf3YxNy6
zJV8NoZENsiDORLBC4dajkT370IqGMXfWMdL2kRwKvsn9XGymRToTharix+1yrep
cGsEbLpcRCQ/wU+JilY1w39yzjq5NHw4c2mpAgwJ6EEVBEyt6MyvygzFuHm5ssVq
XTW+/4JyoAQqDcThZ64HPxz/uZyfzeQ+z7S2l3PsqrlPO7bdO6IJr3DmA/1FJa1q
taujCBpMHu2pgbWAyuRTy5z//ie65yUJR30849TviYzchSvNXsKmcuq6EeFSisXA
jxdCmSrGNYDY4oblSfqcalf/JkK9Rt57ic9djLJkNabIv/lGZbZmPXits0MyBDtE
6idOFA+/IcmC3YcvGr8u5Z28U81lGn1isT9wQkv9+f1ZGvoDTuw3+Z9S+UAaiOzX
+pOE+56VHBazOkaCUoiDgKF+3U438X630mhhpTkyAL/gpD8JMcwIdUZdKJYS90/B
rdntdNtY/gKfLY3cdJm0vKWxcoNX76pl5JcOGR+zVdT4a3s+WFyt5haWesJqeXpH
d7BRxrz9emaaGG0X1/Z7MKsUzk3X9sV+9vNMTCkf4AZBucYfSJHvzFr99ZI4lrns
Kv8wv38/LOU/GsEnA98cuqnVDEOziethfJqNeBgZ9xNrCTBdMcWn+6bInvQeFIqU
enQc3isCTCcw4CXqvNLiZ49kKp1N9FokPcZo3f4siKS3nNR/0LKkilKEAxp53KQ6
8WU0GT1rtrtMjd+igaDSClnASV2QXWX7WVG6r/qSM//D1/zdRPACedL0dA6KeUtq
KN4SFI9C4pEN0p1ubMXXVVABiSJqjBUhI8tnX0DFQkjmEXtN5wFZsFhxlOhYM0jL
LLoimxezsCFXm5HGvj68w6/ZeElrsCYKLHnRfG+r+CcYxKqFR94Ux4eHWcCx0mXB
YDP5ac6DkzK2GBJEVyr2czv2DtvRjsHdjuYK9ve0aU0EO652Sk2Qp94/3nOFxBHC
TsjjRXVqlfLqbbBVOwWDm+eiXHu2ki8xcnN9dl/7c8yJlhrU6o9NHCFdJAHZVsAO
FNC2IIG+cvF5ygVVLiC4abWYK2xaWp7GJ5wOHJJk9Stkuevjku44x2RmN37EOfhK
7OzCTeKHU6JD8dRT5zAK/4wLgXjFmqJhmeXkO9qCcGVLT1V3w1S4jeUFSXUaPI4W
3JOaQ/hPlX3jFlXnUlnM5YaoEfeEk7TtQ/w4+mb9XlBRfxnqSUxNA6DIVV5FDU0x
MD0SWgUAldgju48QrnAMC0kUBKJJ0LRN8Flo3FRe5T1tRtEA63q46WzWgZLuBM4f
3mQ9O5xRdQVILZsgTIUPtHBnJ0Akm52x+4YV+GTD7WIR3EZL22RCQ5Gp2vIFbKKt
1OAVsJ6CF9W563cXdM03GuV6Yd6tSoNvpGolidnGfHc1TsQQymmErcrNgmRW8zr6
q2R+ERtZKOyhXl6VwYE0qjOjroI5Slptgk4rJv1WGA5ivJdLY96TJI0WouaTpx7f
cz/8oVfxFwSywiXWhiG9A+gTcDxX1fRKwCS0A4ZLswURBLGqELb2jF+0AJsfTLnH
LrsPsb1dZ12iOj47DqVYeffT0O0RQS9HB9GyAa8Me2CdVuEnLJmm+hVBjLQQ6JRX
B6DJIDkblHOwiJYcC4KSrfcn80w2IqkliCrPDNy0NCMl6mNZDEjOQVBKKLN9LuRi
Pr5fdoAdvxS97V66GIk/+w5GQI5jrhWB0Ac7sUoZWFmfsryVG5W6x7ZAF6XqtLsJ
lbJQmocLjyst/MgQOX7w7oM7nBYaMhHhMq5GhCG7wj+cJekBLia4Pmi0X/XixfX6
aEoJATWA5xFEwdFwjgvWKvqkUhP7EO8+cTu2Edy3nP8WFDnlrO94zoJzQR5dZmk3
Bbt54dU9Ub+MQBwa1y3ny1xQxof/nGFNbh+UwVVbJh4BJVhVOMlo8fbsDNNJCKSb
APxbzZyQPVLnaZ8s4u4uTmrTM2Oe2wl15sOhWR2HU/OhebaAwvThsaEjD2fmJck0
Q4dd/1hKS9NYwbhDb+HXR3VFqcxTcL0XYgTeLytG5W/A35UZq3VGn6+V1YtOuCGT
gpTpZI+yDCXM+jsyPEt+Ow55LCnh85KJvHWPRIlCbd7aNHwX6C+84cXjXp72+zFz
m6ZIR++kKPseX8atna+oHj7BxiGY6wfGW6118p1OHjdGMo/ULqhzXUPE6VboQoKx
ZVF4ZK2/Vo+cSntSq2PA78gB5VsTEm/+lyhk4Cb2fpQQ5FcvzkK8MAhdSbhGdtup
W9Z1wJ3UYH76KE824OPSIdvVtsS0ML/jqhmllnWZLeZUM95Oo0YS1ep/3pB1Ayft
WOy1ygXBjUKfrosd4ZgYo/dEMACF03Uzhr3xAiPZRSjkpvflPwknKweJWddr9Lo8
XfzqQ2K0QwLNdqvmclQE/aukAJGeLI+k/lMFHZ+kKLnK3sCmUywS53hmtxo/5ycG
Vo7AKGfX0FKdQCbwiXpAXoEAh1Px60m5XL6u5stmK4uDCljcXzZIx9UPt9Bh+jYC
KC9gNj24NASsPNU9hb9Wc5i5Qu3TQ9R8SlV76OTNxpQDAe6NRaQM9dR7Sh1mKYi3
aCKGsQ5TGZHksH5lkc092nNqAtfg+6cOH220rLHwR5aAFvQR/uuhc/dG92pmhPHr
QpoFCvzzNq04Ytns+hePaqXZaElPV/Y33vdGcxaqaVy/GI6Iagflh1+xjmKGZXwc
+mfV9J3TWqN0OHyn993csclk3Jm9R7EBJJCjB5ZDHxqwgDYLa9lA/tyPWp9LstuS
V9+cKq3/DaPXiG59Qv8xskHh/aFWbsPfj6ItLJGHuifg5XURX38T/Eoa7HsP9t81
PUf7Wsqjz2HMgk+kMeP7zYT8xSeNVugrvCNdKC6Tim2WHMIkv1vUfykUXdOO2TWm
tYrW9ZhDgv5Q4b19YIN2Frsp8TYxJtfCq9Y/+7BLKqF4f5P+0bSwx6CgdgztbDY0
WNeYIKX7yI234Kd6StcO073cZWvdulTT31aKDsmHiF392Y5k/jw7z2BZhRfuYWG2
9EJZBBZkkMi24A487I8lJzuZVMtPBFTtdlQvEAkLcvIMCj2sx1BZgkIRRkgSJ6G9
kxFavwp8kJDphPz6MvukDXRsJURZEgdmjnd4Oz2jE8B9WycWuWJFoYQbCAfymwhC
sx7O5qdIX0bLloZw0c9Vk086LjU4xcBg3H6q6aWy1vzaWwUjXuBWf2whvFGvoLMu
LImlcBJzpK5QVtkaT+x4Lmp/myJ9OFWw5BtZExFGR1Yrgdi3Tmf8YXDJT5EZlvpa
Ml/o64NDPHbJ42AFf0MLVjmtb3kjrE1m3sfmJqFW3iuAqpt30LRXhWLgEhypGuZU
FOyF1voqhotZV6FpGVe4RwjbqrLXirKZXH5+xrpnC5THBreCj/tvn4Vy7aaftRW0
B1J7kMu2TqXVkMljhOEVXHijNuVZstaPwquw/5req2xfGcOCbeTspxsgKne8LSOn
+VbjTgW3x5ACxYjW3LGkjC7wrUYdkYZqqvJ6JcEu1BtHe1FAtjx08PtfIjuNxnIB
BHN7KfsmkJj1skyM/+Yij5sl4hp9ZodlmHMVog4uO9Xii9sU689JfVE8T3fwWgWb
okEwVjt+nfiDUdHFQfPqBjhGsFXfpPBYUJlGPzYULJofesWHsOBYM5ZjaczyuFKV
KBuP2SK9rZLk+yC8+fO8tSfu4cT5C964opCAOWF4dodh5tXc3PO2YaI7RbqkUdtj
2E6CC1ZsL06iA8NejM11s29mTDc35vdEIfQLs7rl36BZ4sQtanzpzqBgVV2nerUw
g4KIey7BRyMoY5KHnZDzH7Eu2TngLAqJrkqtxRSbRdCIGxwnV1LByY69XhmsD3Vq
lcur1Jw14zERBZdUxSOEUpda6ojVp1/5siCiq/5qOWPW4fcD4kEHb2wMXlgJ8Y4c
ZUzAwtwYIiJICT8zRS97LlKSYawCzRbj3WIU7kfsD9fynl7EZ9PtepgApnVU7wgA
rb+T/XfVBXNG21KQmkGXWg1A+ZNolD7xpBAVvXaJ4IXpqLUgUc0qq3FASVb0CgNZ
YHtfUWKiiAXWqEcM0RayoTxExZZe5IGvvp69uwR0j6+JoN4YS/vzdGHBnk7PRCkG
Iu03zr31TOiwsfyF02hMPwKs3jAZLelBUqNkDOxKOzPfjP/7pvrqaJguYy3czx/Q
z9cUhL1LSgwA8vj8klwRb7ckBr0AuSIPwKY+xT/19KfVdBFzmiW1t0rtUbv7NhnY
WfEWsATWTiyjr5OpAYRO8kU0dYCdFJxPgpRd/i8UcPKU9yz8xmdNm5Gmix+ZJP94
rdyeK3O8DhyMqTEjMf5mi3tKFVuhPcX4uoPDZB2v3M4gL+m+dpq7sOBtUFd+3sNw
c862sElPUHgAZxBlfKr/C0OVxyXDW/wm+nSdS7l3aaZgAaKXeJPU+N0HSrFhwjuW
SfUlxjTqBQ9tVaGy2HLLBcQFGvohz3qkxHdL5pdSx9nVmeTc3hx1qSxPfn943VaO
bIjlUh9KWftB/sF/qk7/sWQtp+eypX3OQzW3bsHg9U5XijYPMss3EaujDxrCwZgf
Ff+wkKCx05D2beqW1lm5JvDFOj6Bnmvb41+3Yw7Bq6dKhnNmBynOUZnQUAuRbK47
VWnPOl5m04XuF83RjbD+7urUxBs/SYQWWzC27NgsCfH6moKqBY1bzYWfYQL9mNMb
MoGCUFlB/7ufm8DATb0ZFP7TKH9AOkJxsZnDEuh4FGvZmE2woHuqLTc3/mS3YCiB
gsLJyWlBZETTZjXObTkdF1nfCgy2vl34qINKwSKpP49i+HzIrZIa0Kc32plepTEO
THlgF4qjTTm0Gt6sD1pbpApzo+ysN6V9cJVeUNcwNHEDaKOr3Y4dcAa6SeNXWpPm
SH+rlI7oBiqONhjILX4zWKUF/LB4IWt+7591d0+dIeQg7yqgFsKCrdcpl5qxJV2m
VnbCjUs0FJhao3/7KIkE/7A+kfZ54m4NR/YyNU7qapK6oDwGfGInQUVjExHLbonD
/iw7klsCie7G1Qd085ZkHTS84EeNngNDSzl0vtRe2N9/qCXiunc+rTPQplYBqOWZ
1L2kA68PIP14D9cmHKl7qTKTM4wgOB+THtuuv7JR2dnANB7MFNt/imcTVH6Ck9i/
6ABPWKF63pD6xzy7oHtixJoTfwSYOwDKQ4WCJ2QYmo4aGV6HGHFQKPeM+XrG215+
gvsHxd8nPbqU16WXfYtd0r24Lbgtjg0PEMSSU+dHi00qI+wKOMHE94LmHKARk6/c
dIc3577rmOVGp8Echgugn/aaEl98Ai9cqkmosSXdu36OVsXQ6yztztxiM0TPy4aK
oBrhK2oZurERu1ViLq/3MttPIywYWxTph1ErOGwepN4w6tDvJFeHlQDLYoWtbit+
QULJnyZ78zGJBEr0FVd3vjVAn3ZaYv81ZAu1tZaOlMdkKcBFOO1tO2QhHcm92hZ4
1VsLpywm95n17RJh1H9q8c1RgkRZdVEH1jpQOWJFzGT6yInavsC/XpiMVP3MIDHE
8+oVyn4x2kqqjFcn+7XsRTFTDgOLZmE3uzbmgLrKAwT2PpkNRzY4G+iXHLniwzre
aybf41b3FEkpYlJJlWf4h8Z7IL/6NcPkwVsOeF/LLKFZNLPdEDJOno+f4/s6kTe5
h/9Fy/9KjmDIcF7f/ZxgvdVIH8NntWKamFhgHp4r3KdI88BKVdrtGS3IEj7PRLpy
DQbep6wTqTqlfMbBaTwBXvNLoKyuBQqCL/r/9sKQkBS7oZS646sAQfbpXzSfpTrE
heH9NAXFF5kivrorx9LVqarUYJfu5Ljh+I841q15QNXQSmGxVISVK0NGjHDKO6kE
dW+2lq+xzf47j3ikd1u15ln+ZBcZKXsv0FqAon+hYEcTZuq0RwmoteGLa/ghq48q
akjTYjPVua8oEtDkySBmPhntkrQmFuOGxBbUMeEvPvmB+D4LJ/9KFak8TC+39AUK
3/DOTz0pVYFKhQIEgSCyxPW4gqn2aIhMqOntplOMdD47mCeHxnqdRJZUWx1QXziF
lkxZ/cJScinScxhvmRyCX/c59NT7AK8MBq7Lo5l9vYujBwC9l/ggQo9C+NjLFR3S
KXWNSEC1zLCFd79VOhl0IAOyCG1NUiRVOgpU96I4yV2lBcbuI1Gre3YVfF8QHP4M
NorAHKXPtZRB1WiH5rOp0CO5Bt9FizCpJq69v1Zx8FcyH2JhNalWaxds8BXJcbyo
gJusdfyRkqys1htjIzc9UkVFKJf/j2A/8Ax3i8YniVAzImxa6sgN3klADT5MAs2K
exZhO19AbBEx2ArK4Dqzqj11m7R7pqQbSy0qk6TVATFcGj8AFcfg4oRRGXoMG+YZ
B2ZP+vXkaflFj0ayRaxA+l9B3AyxdUM3tCYpGzf/6DCec7UVT19aO8ctI2F1GZiJ
Md4pAtNDjQSj5Kl0rbju0tjDXgjop7S924lS+JCVQu/9pre9iDEzbD68m16nDKWt
GC3JWiH8+sqCskSJT4XsQuzGf5RBCSYE+opgL73ISfIFCt+tDVQ97fIoiVGsXc0A
P+trab3rNjLcK+p792kX/toCrY6HFc3qtcewbLvYXes8yO0oBNMjeaUIahh95f9q
36B0mX5cuVwuFq5VV9VnQ617R27soigqTzrEBxM6QBhYBfs6N+Io76ed8MRsBOKN
HbW6XI+277yL7Xh5vXq8iiHMc+bTcbDsKtc/ZcPjc5bXiz4AMf9ibWZM+T/MeZ0Z
SFnP4SoLPA+A2qlJQE/JvRWcCq84PvGZ1yYEYrH6w9DpsAJu6Ghi4dalHS7bl8uz
oaB54Xo0U7afVp2009GXvm3zy4L34p2DM2QrGO8azN3jbCq9u2rh+nEYBYd9PUz9
LFk7kjdkfwfZ7vDMxXDH53ypZQnJeCS1uk1nVauwrs32dgcO+6FHPpX3a4tPKDn7
vYtcGLsy0jc0qSdqfU9p8mOeGkkLMOftgkc7cn4v9SLuUwL7ku5JMfrZ/QQwJYZL
dp26lslCZJPPw7WJQzZ5KDsRVvWGKTi+eWtD60vOr6SE0RmpzgC2CjVUK14qbQ25
OWyS5YWGwIOdzh35v8q6yMav/AkayRUuvHyrgqj+ICGfSF1uizrw5/DOhDUylP8Z
FeOEe/N7gSslWqd1kM1bDIXwyiHyuECIycfU2XmZ1E/jmRDfYBecHfKcPRMA//mf
O7r8U66OUue7JAtXDE/gvLdKqcuY145KFg+YWs54ua6/NRjP9p10amC8/rJ0yAYW
acnbfzVyFm5IB+SucKMxj7LF9kiJaBYr0NJe7ZY1qcqZqK7chTgYyb+1cuhIZnka
GL+kIs8urysIFPsNKcyiK1p+IcPJBHyGbKYPRDuq7I++HfKXhlNjWMJuC5NXvy8k
p5c6MxtXzsxK0/29As8+Mp0tEKl0sKZK9eGNgOebpxcKMztFFkh2ucWZ51666u2P
77VYisaZpMmPeD+yyQ+VwK85ZXdTbh1dkK4EU894M61zbI6WZTSKyn1GnllB01Oe
1LnJ4Jc+sau7S8qiTcizC+q04NxoPm6N4XgJrE4E+fGNTLZ9muamLB0fJBGxBdoN
ivjs1drXNHbeuSiAxxBo7Z3Y3EJZDLtvYIMH/xLqA2/AjY992hCynjUxPmWXzijO
KEdHakxuWpDJFC3wughOfEeLpfGBmCHuqYG/xYncYo7CRDiNjxFGjZ8u8LPj2u3Y
5fLc0Bz3rl6TjOOtUmXFvOasTORfqsif509rVpcFAsKBOmsyeRO4wPW7V5Yj+knF
ckhsMglh6NAuKNTuVY3sOnO1tm7IuxeZdN4CNekeHTzuCjzD25puFSDbOVaubudN
zm07wSySBNiohFFwfatkF7oe9p9W58nxspTr8mKUydvT3Slt7vNkmgI1pEDw6ArM
VdTl6/b4thi6f3BI/ytGiVdArLmOX96tpMrQSdMoUU7BlBNddWEmp8ieM/B44KdK
ydP9e+VEGoMg1GsX2ZD+D3bOtRJrZV3P2rRbHlLWRTaIDnWphawAHsFO6vo0f3ta
KBG402J5fT5ANw1yVjLYV+jMzDpo+yi4Z1nVRTfvBiSigsLkoEV8y/PPP3o4DiHD
lRkzqe2QVyKORynK/ATx2Ouc7iyDVqkGsMEmCfnhN8e63rF5i3qvu/3kGbWUMfxY
EK0i2690iE2mHIaoG3nokt7SX+CeP0ktYmJ8EuM3Xm1H5mIva525EEYWYrygXWcS
P0xUeCyte5adZFw9FtA/0ll4bVxmPse+lDbi0hm4MlwbrDeNBic4HSJN6f4kV54m
Mjnb47gMR+ZIKVjhg6IaSb/H5eNufa3fsi0RWkkIEqPnioAPqQjM70Or3+hx6Suh
iDWi7Zf5hp8m7f2HsAl13OIoMkwSTLnQ3KJrWV9jIHFwyOlHzO05fTkMWgl1cpzq
7MIURy7ynl713+jNZxvmuGDCPvBsDwstPsFZQUYaGS2W5gYq80fKU4y4zLIHEE8W
YkSwItHPzfVHmessCjZ8xvGqwdF66BePsjGMi/8YVTEXCcAtCNmLFsLko0itedAI
qd0Kn7hrnsXPWUxMZ+X07CRixNLWNhcwi8RnJYxXSrL3X1PTUT0G2NzsYVe1TWu7
JSX1JF9oJv/WljYhPgyQ2QCr3okhvQDt7uHZ80r80vukNC6z4heFbmUpthp7fePr
XWxvFXCsNh6g0uhF1yHhK1MJ6i3b6mMNyuLGHDjDnvo/HofTha0ak36dW1kj9GQZ
YFn4k8zZfow4EdehgsGsEjW2NaOG/2DaL4XDFNhWmiYUSesj5ywqw1YzdfW4SH3n
NGQuS/K3RWGSEAy1Mciw/LZ+lqNulM+QJn+C7cXjtQPymuDHLLzr5Tkyd19NP69U
wgz1AmRJ7E/tgM8fjnsF60TPV3ThWZgCpKcBTzYtXdk=
`protect END_PROTECTED
