`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JY0lTZ8jWqldL6Yz9gBY2Ehms+DqTd61PUgHDdY2MPYoXSjmMnMX25W2DmERkE/G
ATCLFRzkUG3OjZECyMwYD+TQNMlLx171Lz9w4MLENk3emjQ6qZ7W2LIM58quWbPw
k4kYFePAzw1aTvU15LizHjTa7rg/B18+Th/R8OmKhU+tKnRDD/Z783KZK2GHR2fJ
lr87RC8zbqsGI92Vkd19ASbzdeo9q/v+i3bK4YSIlyStJCiWfkVc4d1PCRl2s0Dr
NEu5cb0PhqZjbIkjutf7+mMS4N7pEDx2JewKqDI6OqXFTpznbNszLY1xo+VS+BC3
qJJbKtKM1PwSx7pM+OIu9Q==
`protect END_PROTECTED
