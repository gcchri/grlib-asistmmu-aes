`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2SpfsRxBFubxurm6ocBwsI8hxqfDDuQIPnW7i183AO6XkkOw9pinY+VrGA1frZl4
nGemTgWSTX0Vl6ThZce5uieOuMmFSoc6XBRxeTeBe28H7tzVW7i/kZ+LV9ia4Qf+
zJHcFIZwRVkgDwxOwD9aq6KRL0PaIULPdd0h21KQpLGoixsLZrqCPz3K4tZQAmJ0
Cb/K3GskkkBkgIFOC4sZTiATL7vPg1gIRnhj31s9ISAW2b6esMemZOc7BCjDfMl4
qgrfZfe9StksYckjh551871iwaNrIjdcviF7VqQa4q9eTw+5wDf1L/BCXslXIKj8
gQYh6TH4U9P1bW7Ot87UNw==
`protect END_PROTECTED
