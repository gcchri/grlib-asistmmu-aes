`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+MvwfJ7hNUdPvzcaeOrC3Kb+yuhbSGeYHWuNiGRLE8cg+pGQ1k67sG808oTB5Ky+
y2p/jTA5l62t77yeIfSeU/yOeK0w0vlcPhXUVyaBWn51kDeF+l5hFSagLkx2RB34
1BjsXAdA+msiYEK9kZ/7lQcHnVr5FUk3DlOVi2UMCTjldtB06nOg8qG4L7s24zIw
l+i/Z1QUE+DR12LKPI3gA6l28TWu6SGCcoEG//s9EWOxzvqmyeP2F8V3xkMk4rpz
`protect END_PROTECTED
