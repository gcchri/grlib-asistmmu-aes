`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n4n3lnERlzNGAIgMIttqzAC4Y4Ygc6OcaYlgB1QzoFgmQc7dTUeNRWF1aYl7SZQF
oGwwWXY13/cJhigjMg0TQ1r9jKacS9L3/j36hM3YlqkjLSk+PifMyiiPQ5WyRZ8k
2gKzPy0MSwCbNSDNMWb51dUFtCKhwmmLgW6rvrojwvgg1YiSr0scLJxKtfmbK2Vh
U/X6WVo222d2tImdEzdKPrQi9oh3OTfEqdqys0PG8OfBolD6MaqvV3n/EjM+pMPh
pTvVmAEEM1UDexNRG+XkXHlashPcvj4Y5St3RK/kNa3kLx8iq9OI4rKrTel4Yk0/
Sj4AIov2VyoONz/AuxzlnZSZ4NIp1XxXBdH/z2GEItk4vaed4WmBvNfBzFl/sjB/
ziwQWXcrJ6NXWBuZFhokqSiFX41SWcLAmpA/7Z9mj530LSsSrhd4OO9ugnXc9VLP
PJ+HJNudzr1IUrxdximxE/S+OlJrypTRoSVFczuL51mY3Ch9yqq2mEBvRjFjZxRj
v9uZhhc7NXLcxsAGAffJxoeDjmn02gox5+3UjODpsFqmd5iuS5/vZ40Ns0f/khVx
2eCYbbr/U0uzV6DQ2e6IY2lq+V7Gnx4UtgV4cuFcC/dnVrA5iW9ogdEQ13Po+qOs
z0ADRuprzCF1hnsjSjOzSoYmkzwxnKDJbHKoZnU3ZZY8n0T4UsMJFDps6BgTseh0
exlipamvxchcSMqehjphij4lek9Mus0vf4EcnPuMy+dY1vEUZdjL/gFV4FDGrXQb
j5APBQfExifHyS3ultdlLlhQZix6uZJsUBI3mVaeVCeXrS4Xcxmq+247rQC5XcR/
qDj9mf2Tli7nCuBpBa1gdrfjNiK4QPgpveCaxAXUYXMC5tiaRxKA/nGdmgO132zC
RmQV2/2SawmeGrquoykj9xQIUOlQ8e/JSULca+YFpNyDNiVUUnQY9tR3FLK4dNRi
sfWHaSlt06KXLe1+DbKSwGue1CIspGLHqrI/offnpeifI9OAEKfmMCTm+mOmcnDJ
5wP66qrqpnCFicHePvY/8Z2b4ZWRi1dlPtQd6cDaPaSjZLfVYHfkmelbiJ9ujhCr
jcy6Tyutzv1xD1N2fn3ozddsCVTGvI1pT8Hpo3TK+Kdr+K3fYmmu81i9iVFMyBmX
9xorqaU1LdurQnGZHiuMm23eD2I9NZEv5H4ImadXBdl6XYv1TNQkhQBGRVlG376E
0bRZ384kfAc0zKWDA3jNkTAyghT5j+cMTo2agmAUQ3BbCSTZrYE16Y3zolFSmr2v
hoIh3kraD2G75aeoWD0mY28IMcNxHVNhiusGdPNpczQAgZQ+ddehBBicUUCMzBf+
jTr7ADUl4fU0QeOO+XrNVkJCuqCDvl6BjVGqST82EbBfmKC31Gj28wh55lhTWClZ
vL5nkBuBYV5g7m23mZvB5MK3cmVNrd/bhD/bdYX4IxiTb32AT76JBKNuxoYkZxzn
ow0XS3rVhVOmrgT6AcwO4IUse1OD3FIbJCPI0MeApZYcbLKDGeqmCQQ6HKrIrloO
mavUOoVozQSEy6+1uGqLe386lD7EdXit1EaqaRBxJSfuALb4hrFDD3uld3UdRUCH
GPosVxiKPh58lX3WwAPmwBx/H+VLic0w0T9s5hWSbvEAFtfhkOyKWvjuq4bOY7rE
JjwFMvwbihzZJFV+4jGb/RcN2eNf55nmm/RQ16JRlo5Ngbx8j4RmAKxpdUTE8ib7
CnOTrQitzHZ/kbXmD1mlVx82o0S6KJQjAgutGd8TlGPCuK61X6CixtZIAtoEBeSZ
PbOcgJCd58k/m63O6WBp35CZWQrh62JcOdBnUi2jktWPF74AukyK+2YZu1q1iELU
Y1e9QmxkIKv+U7FsDmg1IlwWr3WixFaE8LpvYO41Wd1aXLGz+0gFUhdCIs7EoSf0
P7+XWcBubf4F28CQZyVxgyWlSVlcx3Rll0c18zQr0UlvUof3gbEePFrp5QwnNWzG
P++GEKDa/nbMB4leJp/078rit4qJQC6/XR3mWgwYMIsj09L2JUjaYJ+VoPfBmSJe
zH5P7QchdvSo2ijZfr32XbQ6hTWUjRaD40u4CU7/cT0tjK1p2Jh5ZXViI7706X9j
sXPViEtidjUSUwS8cFt2iT1nIVlwhU1LXd0alEfzEvd+t3OG4k8HJ2oVwwYiJKLE
PD0WOROpCBU5RTHGKBzz3eosYZ7rPRNPvVFmvumg7J+wpCoEuqSXtnMj1YU9FLp7
C9qLWBDy7nqYERc8iDiHcaop/YwRjTYGtawQBmoHDN/3NQLB+U8lB216Ibe+m420
eQrTElTJ5sBItuKr7qxSO95iiiS1TpMgzUHR49sbm6vNe/19rhkCxRb6HcJpRMJf
VrVRsg4gsI04CtiUrzviFraB7EQmhZjC6TriGCNkmx2aLaEU4a95RcDnWL6gS8n8
e74VPNTYi8siigua+9XPnn0bj7+qf0r4jRvz56hMvXdP1oquQiPObVAXkV1T3NNF
EoRvW0XVQoAFMbJlDsHuK+j9YUdVP//GMiJ/GWLUr4gRwGvM2U0AjEqZbg/4Zy6T
7QVKS5VIYEH6Rf0knqdK7hcjlXT2EfO1Es6766NVQMSYUjcwr79AlTjl8Kge7HmL
32M8AhzDokFmDy6hbpJfEavzZmaochFcYDz+FyHJvc+wUFrrd2lRP/ebO9wVuzyD
tIrwBg8HmHgZle8TwqGgBm1DRs5RmzJ4lV63DYcSqYBuDY9Vwkh7JJ3OK3kQ5WQT
NWAY37bfmxY5A8pJfEdUnKX7tS5aGPXJUiRG1d9BXazRkpORTWfnIXByxrlqze7k
ahbxflUdoNXKwLFS6cHGWnyd1vuFHw7Gx1AcfUU8FU65q3OQULyd0/O/D9vjVrc6
gguQ5VjlWyxckb7ptj+hoUUttVLJPeH457/MgHWNkA/Tc7tuPNMBzGCZiqHPc2BU
td/LFgjLH7ldm6RIQnn84YftkmtMYG/n2Apodv3koBVV4mjt9antjbvAxNlmgjSE
zYDO2RRtHS7gqI8DoBz0Hd9YnWoUYXA1pvMU8ZSwBl08avczYrQjGlwp/nZIU6ak
BULL96D3kBrln61IrNPgcwdmX0E5BktmmMXEwA+LcfMJCQRwXClcTRkQSbtHDktY
Rzn8Em65F7GIukfHmLH0jdgPfuV4mAMkonZP3fjqGancfnC7coYSfwFCoAf9YmyF
Tgn3cqUbYSJCJYxtRbUQeJxgMx8+qe8ojl2z9t8QnYcVl6rkhhqA+lGIhcAh+TBD
aO0QAz6bUlDqumaRqgAjZi0jeRSWQgZ1eop2efaBrk2FigsgaghhXzQKaFSUq+G3
t0D/1BloLn/jV+3kKHoXLPMfTlqB1kFzP2Xcdr5qYExBxzWQtKiTo4r8dEHxsT6o
hVZyOFXXttS2pkz2lXi2R/3WQiepRfSbAkuCaTgv6nPqm3w9/4j2vCOqzh+mVTRA
oPwfru9ljCZJy0vVTP7eAiCNJQqtBSTb0x9aJAfAHCRzZeQknFSJMFylTeAbVKQi
Sv3YMqIhIdN+RlKz64ucTmGdoJAUqV47m0ItARYp42EoaICXNy5UPgx7stAG3nL9
6KWm/sVbHO7YaWX4a3OAc1uEydyDs0AKeKu4TdnHbaEYGiBUXyXbpOuA0Y8QBNXo
qIAKLXHUU4P8cI5K/mDXrH9+8cS6FtAagXWA23GWHfpNjYt57VvQf8KucXOUuhRQ
SU6P9ZgEiDoyd+G1ttJZjh8cFEAjKqZ46axK6IwVwiWDF+9M46QUUFf008EsA+iE
lCZGQugUu91qrPY9MhC/yDapEuEfjDo56p25JZLNRzrL/8JL+LGiLoa9y5z+6dQ4
UswHi/3DPKdJQL1689KWaxA7F4H1Jv8Y2LbaUJfiqA5+hW1+0ACLXbEkLTNP/K+M
WiBrCqR0avtAaOdtFpSEMuefObjW8twT2a8KV5t3FU+TRjByARVTph4FddWFYR3C
GOf04z2sz2LwUB7pjCaTk0C4KRMy43st/ih7Kam4d7yxTacB/KXF4rJeJCddTdSw
8+VoQZW2/wsPy2kG5fxDcOVk3PNbGsL/ZbXQgK1vb/OykG2G4eRjCEXH8MU/vQsR
DnSrM26Qwg8xjjdG7vf7S7dKj9qmVxQnuGIWfkO/aFpRp5slvYMstpc4EGbnnQSX
eByaIfYhCjNSFsKcBf+6XF0wbNZN27Ig0Yem4sMuLbzDx8qlyH/fHy/UHirRL51m
1fuTCVCI9832CpF3ibEoDLgza87V8pyB4ipVbscWRx2wqHPJezmHrOn7BbWF4U4c
x0YRA6Q0pakd8ZQ/OJk0UL1GEwGi5C1xi0H6ah2/ZpNn1M0DO3uacWy2wDj66Fwt
us7IFQgF+0i9QWvN2tnAXK+xK5NR8htPnZI1VBY8Gr06AN+nCgk5I1DLaRSIwdjh
Jz63Cg/wurds4u16LdNKUlfr6N/goJc3954TDTY9WL0EaUAO1W39KXye2m4uC0rS
vVU45DdLQhZiDN36cndTsdD5oVEXhvwHqPMEcgAoV3j69uGER9lTxGbcVwcgLgnm
wz4IT7pKCMxlMNmYgbSvEm/2IXfJsVFAoKAwmOQ+yElfvLUXhsUG9TQHndumlyXf
i9O3O9jMkmP8Ypiz48sLP2X7kZycUB2N9P/Qdm1cb/TmoYgVwTfJkuf3a2ql0iGQ
dP1zxWX4w1FK8PuFxleqxC+56BbO4X5EW7VyoGA3fDRkHRp5wRSUfKJP+HzwuH6t
BPicOnLPymoJqdTkfQw0pFPctcV3UFrSY/Tpiq+QPaZCse6leDE4yZaiCZf85xPK
BYv2rkkVaXsIahr3jjgoczkJviUydeMWfsWfXzGGpRUezDs/yv7k+NnGz2p+50I0
dEGcLlJqljsYFQ1juyudP3odmgpSor/UMP7wpXFErfP9FqxEhfwk/mykhAqap7DN
bvFKxMjpOBQz51pUPfnAm3NS8vbGGadGRFA/U5X3WYXVmONU8OU6YRKapSiqMukD
M8TA3Z4hNSLjywBxaDxmKRyo2Lk4Rtt+X+A7LbQ+Hgci8uHUm55t9WZk/ztSPGHh
Apj4dSzM/6l0j+UPUUIQY9LUUtLeHimuzZbzafwM+3QyvrloT32lB4yLlG7h8ztO
KhjAUYi3livYvdFjQn0wl2iLYNhwqZUM2nTE1TeVTufzqlbWrZvJC42xghD01gw4
1kMVjeV6+BTo/t1C/qgGCOqGaFIzucaheVhKuWFRwl2DyGO9to4ooC4zPBbucrZD
Az3CYI+EoZ2DqDt7h31hpXcI1OuQF5ufVW8oN9SxF1Y7u1x7FRVZ4qeRYCY4yy92
jyLSE1ph2u2EZi1xpi/PcSAU2xhMUtIStUrRxsZZXjumfoTQlhDBREg8IQr81mE/
cucVy9nNwL+7dBu6j8N9Q2RW6JcpQlqnmT8iBLqSwTJBZfvLmi0Xhe0KExwWApwt
n3PiaZfTWww1/IIbXk6g+7RjQLxIqq5GM5trhVsat50XkmhPpDuWifGfUKrpMmDp
Oi99jY5/fhlDfXBtuF/aKjB72WCGx2gho/TLF6aNSiioAfedsYmJwv6HnEyUnT/Y
uJffLhmAGRKeJzF+ma3H1vS1R6bgDp1+VvDIA//uibPqm+oXaJREWET0ttGuDJfT
1WNHJElemcjrxXB/IynkmaIj9+g6QJ5aiSTD2t8JDXFVQOYpxqqMDQGom3yNbzaa
QEIx6fZchWFltVWzeuiy5ZW5MRUA1R2KBenw+TEbiVKiY6LKYVB1+V79Qt3sukpo
lMrsB61SYtfoZEZpjG/ctjJXAQBWM/P2zpX3XBtEAFirLSCwp+fFfw0WDwnnk5hy
/tf/kTTRTx+m2JzHe9wNtnVwpSsnxmcrREpXA7rfrsOpAdLo0Hp1e8yorxy+lvlz
ipFPVTh1Jc3xBE+FA/EHChP4+pCaWjKAeemje+DGgigSc/bIzvOhtfllajPtxHr2
v7ICs+oaJorPBw7F1MQJoX6CsC1b2RLdgrHnZxastWXtj3YFu56bjO0dfPerIqDo
YVrtGiOC6n9c7Z9e9W95OgyveOChRBoNorUE/Sm3FzZN3G/xX35PTSUArvyQvc//
ix3ffdPafu1O9SNTdfEUPrtMBaSkfHsJZpxuOZqvCeKyGEdKOHtdmis53+PpJsrP
Y2k4BLwBb3bBQDR+lv5wifuGycVK5yOP6Q6MOMo4hnt0nOaFRJhQddUapPClin8A
ZJR1T/c3CxUBgGa1j2i8XA7lvMQNYjUhvYMY47GUhzdZN8Q2s3EsKsmQtBCdH78U
dNUXx/LsIMohvmfL0AEP/ecLRL1b0C6ZUXfbv+DVnr3+zUflU8lM3B4mU4QKrfjc
cxFHbWBQZ6gCt7fKxP8alPuprmldempkmOkVRWLQh7OhlMdp7+bXzILpEnF3mgTU
nnJSefOyJO13AW4C1bGMEcZYz8MjT4LCFOeRmPXCbYApGsKwNCk+zW4Q3IikojGl
QyApHgG86doPtV4uWsDh2ZTOC2SPvGdctYRkwMPkPpXL8SxK426+/cBH6i3oi8HJ
Ay6yU74WCsi99gIsIN6xx+9MRcbdq5x1WxVTbzxpHb8VJpRU+P0RIo6KO1CD12uH
tY6YmIU78j+73sJqsAkfTjbRdpkh3xo9q+NFWuBPA/I1YeQ5GPcjEPdAw6/7anY8
eSbWpJHzX18DkuL1zoh683OqFSZ5gw487Ctc6bWcUHez5+1OE6je98jc9LDMaHA4
BBxT54Rga5GyryhC4spS9Or9cEtf9rfXvp8R8OlFk9/+daIpY6nZVou2k+/uUJCG
BijmW49oVKAFarSSxvVLDFrbgiuXeyqRoCA9xGhcKtbJcB170BEUF3DFZPXCXM4f
kXvk+qn1I0m0SdgY2GlF6Laf55SQkwzH1oO+9twzHttcHr4cOteq9O19qJg8EoFt
kfdeACGhstlFWKXO1HmmDeTgtRXvR4GXbZ2a3oM1VlMExJJJ0AKQN6vj9hEKzYtt
7W+1+8wp8bHWhd+yFSwEUDi7HHDVGfmYgLsz+0Zh5AZBCU6jljJpE7pbmB/tIW+R
woP8lBsRLkbQDTz0mLaIjsS3gyUZnniIyXNUuaFi9rslODyCtSJyiUbgmCNrA4Sg
DawhvRyXU7sWrPfnLlarBoXFftg+Vlrn72u9CiFkvjHCgFSrHuFtgWacfefubxUK
ebbUyphv2T12tVwWUeGFnqB04azSTM9eS8JL/f+TGWa1kYqv9AuBWkI49sA9gpCw
/MVtirzIPpGsVrO+AzSMuXWUW6GDajxBUZQ73482JUjdp2ZH4RzTAqfs8AVjrdvw
9UBjUTD4Ouj/K1TMTia8xCzuy10t2oamtA20k6N6cI6XEmIxf441+0vz9giQpGuh
2esb4UvzFW2OzrSqJuNmvftu7GvUx03EFprE2maX8iaHVXrWHgX817py2rxi0edW
ok/D9xA4rxkWYauscO2R46seCi3kCEEfZreYTTAChtcfreszV4/KRhauZ31qtlec
aMlkamKSOOXcpBwPXaD/44m8dLAx3rMm97OaNqthZ/4PDfGFu7KTGqgzyVmeiFi9
rToFaH5RMCQQCuyV2ytFhfdK+bhBl8aTSi0f8cfuVzzA/jz9oQupOrey+84dqJNY
xexPM6L6Uhr1DTDnqgsRKsRwLxffQNtrYTn4jXWd1eFx1RjXU03xZrNFIHZp2K1X
qdpPRPpQn3hThFQhj/Gu6c4WxaSvA9xF34zKWX4MCgx4A1vC5vJmcDqSWJGpRClm
SoeiP+XEM3j488BaQbC9nKqknmpOo5y4va8zIIZGgZytCyI6xLe/07ZmXsyZleTK
04oYx1rzgXrqNFMfnEWYM2HRZYiBt6Sxv4uVQvEZXy2SqPhBVE1rORWnWNrrCBGK
s6EynR6leQQJvfumiEgdZGNpJMW/VpfJVSilpX2w0dLL6FRX9Q2R7RMy0GiXmGC6
shIytTuwpSbOzNDiS8ds/moeKj5WOvSJQIzvfoz4ADVOVXT+gPTKu4tuY/T9wdPM
gEhQ1RLgtFu2GFPT4gnAIA5bdFrOjAzuDQSPLBsNtQpXSTfENACVp/jFIVifIv8c
L+cEKKNZCdnJd8bJTZu9Ow9/TQbT6VH7BWYApE5vTvdvZwWXoHNo3lPJEM7m4oFF
0OGk6cHkj9eRmUvbxfDUhACt1HmmcVlRJEEWtEHGSq475PZQQsia5Y7NMxqeMJOr
yoBF3DnHbSZKpeRqESWc6Uovuqphd/Q51fhqobsagrmi1wSNPBxspACmYwXymuM8
em7LpU/avCBbtCahu9le4qYcAKVTJzsTxu985ut1pnFUBBqIaUHWIbq5h9gb9AHj
H7Eo58FMl988eUXjcfMxci+suKM/QyGhALp1ilGJwDeQUWJxxmV5N1VlXgL2wgXW
6EuAY59AH1LRV4QWNo0WOddLkg0n0id+wSY/HZUl0xGGVEGkBdKuK/1Czb7oZBrQ
kSNdkhw9I8CJLyPM9UC8XuSKCiDL36ybc0WESosB9n6yknzqntZhRn8qrkTtXR0t
kIJdxlfSnmlhgcgGl9U3RqiXo8JnznmMs3CoMOlFK+H8Zl/X8nS78A3ovPLObIz5
vwaHy0YRPMCPji7pkimnZV62vLz0IuwHacbhucVABqxUv6679dzJaxSGnamujEJK
O552E9vhSqL1dJaJPubDRqm1xgGLqISLgJwLztg90Xp8AVSxBncJhzwQlz4ZEN95
alF008pJ111y0odGFh63ItnJCG8mDmuTAYT+exV4B76KhS2qwIv3NgxV/I75YEC5
5hf2jeJwdEBO7RuO0xM8VJoJpdUfKxWL9kMwyBpI/0Jk1ibFt/u+9QDkdGGPbYWF
gClkdMBFVEVpHibMG7OQsXXQDXT/93XiH+5nLWI6GrECOG3T86y39eZefQCvKdoJ
kedyi5vhFysW9eoet0bBh+uX1i1u6FBp5dz56nj1XMVkRyXP6eZiUgB/SLjVrAn4
x+scCNFOyKsz5ZDhQYJ5YNYTImDNuYMDkzjXjC+0gS90Q1NceUtsWFDHZ8C/xQoD
AjObiMX4ubHy/imqtn1UGdJ4kbiypL+fXIeL2MkKX+vwfsXjf8kZViVoXwBSLv7b
Rjh7s7DEt28pXgdt5z6+lC50cwaoojPTwS5xra8PkUZ25EcXqFbKUAjxBCt8G1PU
4u59uR8HsMnEQqqaK6nd1On4lxKh+FI0/TlkbPCO7q3qO/9O92/7ThmSH2Sji3G1
oqyewQPXpxS2r0ZhWZzIa13gkq6QdoA4d4qu+ONNYlJbUKvCX7Cxa14Ll3NJJxzu
pEJ6JdRMlTmUefCzg3waTdQg3wHo93pHOTdUstPWl32wiQDrQnPTX5c87BZESdaV
UT5zzSNi4/Rq4Un43O1guskDdPneDZwyx+RakOmE9FzXlqgsQyNEDFFvAXArZwB9
wUb3bGpw/MbybVwBJwxnPFfPrQmDPkUbcnoQC70/vK56sterw4PwheJtedbi5dRS
RWl25i1wlFQjVK0YugQv4aNCowtL6fbVzj46e5/Wd1VCshyYbBH//lA8GRPjs+Hj
LwAwYj1mjkAgAxAJyPEEBXoZ4YF5POhzB9pUkG2r2G4+Xw+RM5SWEJQId1Fk4bpd
e0vvuv/oFVz481t7/0jESZm/0zs14MUBqTsvxX+OqV46pVXpwbj/PxD6gd3Oi1jm
zYtUtE3XCHNLfNgENHaYKLNZZPLEolfywwgImuzwGcGtlxLibyMpLbsKRp9QPJUX
0Y1xIuquvZ8Go4PlpiKNPUhXes29wVsj1ET2rX3kFf4BfKyTv2jxsbtrZorO2hT0
WeNyYD10m+JNaeF1p8Kafj3lToldGbCU10L46oyGNFNuDPbBv53rD8B1sb4bUQnt
SoIzxN2RbnfrqHx8jlnwPtkIP/NU1vV9wPIAUwzxzsfNX4/tTOETEVvgZbNOXhOW
xoIrL1uDafEP7pBDyBiLwKCIk/ko8rcPu93N01Gfz6c3TJ+plQ/sVoJrj+km7c88
Zg02hqjuoPRHnUjMyf3Dc0eiIcJ1pqCJ4xHv6QtvrhIVGDCkoPHni1jbNKtshmQB
OPTS+TTcUCXstnMVi0VHvZ4shJd6u3uuoFkxV7XHs2II7cAlh6YzHPuR/RYUzZNo
0fFATpH1itFPliYcNbZYErQhxrWUuqoIeOdW2T5qrmMl2s6ffstO4bkkGHZVVGWA
0AIoc5a0ErRFhpp6r+JOKVVTqb+C9YCKwSNSC+8grlyhDQeXB+iUF+2ts3Sbz/8b
cTYAC9dVOV9bIGYWenz4HUXa6pcmQtDafverUHzRwLlHBBeQ3Wh1jMMhlF2x2IFT
HofBc72IaxgXlCIS6nYOGTwXrhglP3HsvSxnmUay4cZq0gnil47XUztXL/R/h8gn
VaZT+MBLs7rtdabskQ7Wgar8MyOMT2KKxbGJJePW6/Jf6AOt9AwqJNwXXLbGd5xS
orSHxku8C0Hwd8RSl2OSd9c2N0SVK0MDhcREunRrVsL3e+b5kxYoeD0c7J+sSo8v
qpw7c7BK2JKUKC4Riu5MSdUCOVwoA5Bh07rSpOi0B15TdaiYnkvUaPdXN82oEbLA
klB6IiFF5SWjFJSqIvjEt6fPCb2emJQh+wqHc9BLyRKNRTZHtxFJ5kkRzdhoLkQa
/gGE44JgJB2UthGgsfJjYqb12qyNzJ1CqxXxNsY2D0MuID2izEjdHXuUaP0jcIIz
bzxBE4oa16ANk9W+tSfFgAfjbe8pccZYGDDutaFVxZnGkJuj2Kr72OSe3YuLUM+c
EOApAD2Pd+2cJH5PVRdWfBPKbcKE+FkbvarienpLAD81QockjD/j9YYb0Js0PiK1
FCeSdYPJoJpNMRlAmVH2fMLpSPKC6AmBlXKTM56qotEw1t7ECjAV1SVRo/q0fU37
qsv+9QGiVzMV56OMBA6g20rqsvnnzgd4cDS8/+9qJD1o24/n2LrfLCvdcYSF2Hwm
mbbRMXPK33/uOQ8zDChvrUc+Ph57vS+YCQEQC+Q8/ZiyS6KMrfEkQBm6Ny7De3Rd
PH/x8MJcM3DvKO0qctCPcRO8bOqq1xmnkdfa0bwq+bj5PDZQDwOyw54R/ebu8Vrf
afMq/2mWPEmCAP6QmLRPcbeXp7TXIaD3esC0R7W75jQ/3liXyHwonV2OiL8DIc4H
b/KlT+ZN+N5XhXFJjDYtg7y4pYonx+ty/FOwrDYZnaPZt3WI1lfvFHO5oISuLOvL
Ca5GI/K7+O79pfp9MjWtnfSeqzOcBiLtXJ2XJxLzm76dX/5pbH4GSckJA3BYPlgq
E+TGTFlFKN7j7ZqLcxyK5e5sqzU9X1wiV7fUpfTGnFSlaj2XZzCulLQraE8o7Ae+
icfdP41ie+oEbU9U3GraVS4BWHKD98uxYaJPo7m0ym3tSo1ks/b6APvQnGVWEin6
x8DQaysZ3ygNPc50Oka4oByLovi9E5bR5FrFWhJsTskhd9Lm4q8r3N6eXTNz+xt6
JtSRgHLqS+h8lJpErUVbQLaSTTKBMWxOdWzS6kYEGwNWp+HluQO80Jwd8rYxYpxD
zjhrBwLuaNk9I2ID1IifOS00Ux3r4uKsZdf3xL+zlaIZQSnXnaKbjP7zTGsE6ayI
MDLWSG7x+6wsa8scXaTlrI0tjRRa0iKlaG42lqky38ibd4hQdugbJmHD942C5Dtl
XkSvH7HZvIVP8uNSBO8I0nELr5MkH2XLo3VftIYwdcd7ZMuCcqNNwOxOq9S9JJKP
zaxiSCMA/snx/k5ghzNKrpS3F6QDejMDPkhQy6SS5LSzefWxPU6c9RTQjXfYEai/
gw0GTDs77pcF9ETWVxpNsUL8eAn2p9b1EYnFvwDRGmG8wbYCvU218XsB9H3PAsXo
tbftOFqDu+jKy0NPyyTr6PZpHgaylyDoACVssk53p83gwhTPAum7Y1JYezA5JsJL
y8aZzOgn3fCPzC+Dmup9iLq2UtnW3+/qyF8pwH9x7MP9HE02/R8PVRHDBgsyoFny
ixBxzIap2UhJGsxGgIfaN0tlN3xt9f2EKA96/KhxeoNfvAjjv4rKTHRZgZP2ojoD
8A0GkTWiIJ4XCXp2HaNI6D9vSPUY99KS3AKta7WJiX1cQ4bX2geTXFzskCmmbmHx
22SG50S44uQ5yzS8mxPIPZ/jzcP1uJAQRwnxwsyEZg9Db6j5YOQjLfpfaFtw/czQ
M0SpbF01hgfhmzfqyn9PKGU6Y4alKJ2Aft5CKC9j1+sdN/D04Fy0vhD2xMQqs1q4
4lTNk2qNbFJoIdaVNK0pdjs2KxyQz2EUaFQer5ZCfUIty2QP0XzqPixJso4pD49b
WntZ1N0L7gbuy9g9MYGEphTrxWzEg+71Xj0u4KfXGolKBP4PG5ukiwWpdbXS9mjU
HRXeRmWMa2zhK515R++AsESVJ5N0Xs8INf7wqM+EKujRmB7ITWaKqm1oUDwgJVdk
UtVpvcj1ZjR87DRYM5Xvi5GIsMAc1z8ysOMNpXLpT9D0jjA5tgpuzZYZFSCrPIry
5Y4M4P3U3mSY50wVydI24BBtgspkKKGFgFZgyDlZQ1nFFyoqmnvaOBxx0N3WPiL/
GBntfDNGmDWy92Mfh1Ypab4KR1phLJ+spZn34CGeqmPuTpVFaasd3yskziqomFyn
NMb+gzqiZmFvI+tbvxjN9XvPlAsr0l2q8MdyDlk8xOyQhs+wt4XUT/BlbMEVF2L8
vlWy0qSrX6SWDXEZe6vuCwtaO6KQSWrOqd6czXwkU7CCH8cslqJN9tFOtfyfM0ar
Nid6r5goC8tfrLDg7alwDC5TCYPsVfLo5szBIlbsZIT545ioUsrNujJjRr8Bm9+f
YeNiNTKIhWWl67dI2czxrM30QYfvi/bZ92ar2vblqNGRrvquUDSl4a0zJ6KVX+9q
P0TgjgFKuc0zcoMvKgjummZTQZ8nCPQqSPPMc0Dnbev330e+JA0B8QYfiuuAm5/C
tFhhd+F64X8XVU3M9f5tA1qXeTy8tf1E2RPKh2UNK5oOtArXvDbyTFx5AJ94GdSR
+C2SBvGfmJXzksv4u3TJmWCf2bRVpFBz71CzV+7+IRTu5CWf8wbYjAfLKauY1oFi
0oingUHFBMN/MZz75pAJ+Y18MtHUBpwTpDdBuMb1ImCe0u83RiNURA19iXVdeNh6
S1unsHeIccFOOO4EstBRXsoXP2doTtKC3zBZisFO/pV0Aamtr7SrKoLc9tvMGzMb
AjZeK8wbxUwQRV0UAyaPRg6kPfwHFA57Vi61+NDcSilmFuBQb0FOKT/MdKaciSAK
Zoy4kEXBPx6YJFQCBFevWTMhtfz6jA8q7pi0RkcjxL6FAHEchUarblSjmYwE6zid
y3TfgVO1aSOscdZJ1vDdPl/KIVGl/p6TqQAjJwMBFojQbFmIYoT7nLHT9+wJlyE6
iT7j+Sdq5fgNY570rB3KDW3KMMWYKlx7a69Oz75gDBDRFmkaQV5qeX+ZyUHtRTi7
oRZ4Yrm2+i7WhDRvYAueOmQnXxY6VnTLQfKrxHOStH75KC3Fg/bXfaKXXinQ+bPu
OMg4buxngdqRwl7aLFPFx+Q5s5gIuZ4SWXF/fsf7GHOy+mmNvGC94aw0ZW9qVZcm
ZYTgsB9X7AdeHvzN+LUSYbksA3Iv/s1WHJV6fFOMzv7D8Qy05NRmZOp2wXNda/YI
+Hwt6Q/b6J3fdC6aZt7h9iyjqlZ85AwoG3oWPFlqYV8VkHHTgkLf56se2aSNy3e7
ZgiC3p8juLJpP5BYIoi0Edz/+oqf/ZTN0n86ZJia/ZN4hh5+rwzzUYB+taiIgEme
o8csDLDwpjoA05AaHVsFsrcU5gv57VyoDg5KJPj+ntDJzpI9BA4NNxXtiqyugZuB
CmyQrYYFV1oa6eBgabDw1RqIqIxzy350rH7QqKcNRB+SkrAbj484qK+YmUkh3QMm
UsHv/92nAnkA6lWUGX0W1h/nzQfJ4VstOlPbw41A2Wcs5Zvl+6A5v05kKdajBa9F
K+PTQDh+vi2BmFknbuK1/MBhf4qvwE5p/nIM3bHw5bwO/cxTK3C455iGz1YNSgSP
+RSNEhgRTq3syhSqv68wUZxkSkQIHHRqBYcahEHsUZI7a/O+1TskbyXmLj3OnuzI
7177OcTVXal6ELKwB3+WLx/moJncCUpKOEA4LvzOK5fpyDdEkDFP4hEBcBrlgxy/
IEcUiSX5s8AVkk0UcBHWE9XA2yMdLdqLzXfecb3+atAYxMesiuKF9B6fnTF4/H/b
pgCsEdVBsY1rkoQqqeTNx2pKhJw7tIFn8TIi/+JV2V/lLj1L4TAR2NgCW8ngkxud
FPC15F3TNszTif+M4XrsJJSYUQqhmR/R78Fur61RSMqiYo8ixcvLAC63hVmWZrPC
S5RwOxsFP/k5A8vQI0f1VgaGDdJEldwq1KFBj9z7cQp12o07RiRV0j5tq0zp645Q
nCxEQGq/QmgqSVMvB4zOKcRqUavpNL+duEx7d7tuD/tuUTbF6ScXu5ilsXbvUO2W
RHLWOaJ7nCcbvALK/n/JsbKruAuFcQAi7ZyJPgj7pP6/tqslYFiK0zrsQSWAeVBH
ogNND0oN95H6hozCyLJwQBR4hmdecG5BBICQcDyXlfPLylTBSGXiBLTwwqzUfNbE
wiMDlcdK/c4s0kRXjHsoTQ1sDvUwNv2Crjs1suW4iWBym6udO8V1Rn8Fk7+Vyr9A
povRZl4y5WT0O1tukEwRsJHKl9azwXOrGpMmmZgKTFZJUHOA+FxiM++I7esTTy1o
O2FVkwSOYWWNt38jSCMSDozYm7YgVBX48jcYcgBicqpQ8TGmpBtidFFrqASOl7pB
sJ/AbYz4m/1x+MvM1uXiDqu4W8mHWZRv6nM2Q7xJYR8GJ1w49BeZ/FBz3mJwWQWj
40C9OscivETQCoBPKBc+zuciPYB/3xrqms3t31Om3b1seRv4ujIJ4fDMZLIIcZKd
PyVX+yWmvh3AVinciBfoNIdQOdih8R7Gjuyu7zf/VjKAh28eqnqk9lRiZgoY+2FV
eJVZN+SlYjmiSnrH2mgC+yN2c7aLiCy+Dy2io3WlMQHAzoM3VFdsqbE/v0hNW83+
Z7+iQfDksA6vh4a0yB22Ghhbr5W3W5HIYUiLEBxRAXGUps7Ntk5bGMNFvfqM9iRP
WBRdBs5BmA0HQDgrpxJ4mW+2/4OhzRoLjRgQPVxsiaSmxsgnFLWMUjFvMNn4+dLA
cOOc2kyrpmpGb+hBQM3OIHtjoEJsTPMMZnkm861tU1AUY2n5fjnA0lyh88tCdUiD
6V+pOO6Xmy7rrUrxgG+B8q9lDA3Zhlc4E42O1t58Q55JpdtBOz0tZHp3NHBhWABQ
VMAi8yC9of84pClQp9GcK7rmwWQC4xCdMOpmQks/xM75Ujo4dqFnAHwfzHwwO7np
nc0sxyJzXjmCC/0eWysxWqtiAKPtPu2bF5bC5bvy0yi1Ef+vtK0KzLASsPFEqbMK
cIlqyQOxIc4KzRVBBPP4q+pAZZYdJzz9FPlhX3aI1SamFa3BeR7pE4IffE7ImS+o
SWgn7MhbzT7SRcnkCQiIawGsuzPHRLyFBW+bbQGMpbeJkxwcKWQ/h9B0qSbPQl/r
uodsHuppjQPszqTaPkX1o0lWfmO0j5FztJN703EuDthmN/zuaQuUhR6Nz0mx1efO
pt5Nk7+sZaxWtb7miNKVNbpnJ6m5nfSQBiOw6wNh0aXrrpba0pr/fzoQjrg9NCTz
Y+xh58ZpubtVyuH7ZP7ZXkTaL3Rie/C8ZDpxThBfhxI9whgwruBQi1OFkwGQrZ8d
3gANZYkdVBLt44YhJFBzp5SFFfKgg03ULxyjKK7mmlsE5SViIO5Ni5fmSzZjA4bT
Sq/HSB4eqrsqXaQtJVvz6mhvgUxLceZplOexSoOLJvLVlYGf55beYb7DIXu9sp8I
KP9LAgkd6sUDvu40hK8krfCdAqR1U/jBsaeXnt3Us6wuy8fnDu3Fna/UC3QpZa6Q
PLb2SEHmW+007J0C4STJ8H+b8KiuBZPQRqdRoyDfi98OsEcEqgfOVt2Ab2ET5Rx+
kdajlab4eg58wdI+zI6AJavDIA66WtUt9mkU4tNZCuYZl7bET7qHqf7MKO0L9BVs
irMkjoQrWhbqhs9lWpf1rRu6612Pa0RtV3b7VPu3+0ZqvFvbciop/eAMM4yI0VxI
RDAHtB/J8vo7y4g18nXLf/yryg7mM/qpk8apb6JH/61T9tV64VS34No3V8YACXq9
v5hRzR5xcBN9MEJ7PQcQhYCxXpOB74wWj3Rnv9qSa0ctkFNEOGivpScooWqcW2Ak
VIFsEooNeE5EgnwUf6oIrsVGXmzVN0RnjJagO8OLqUfTOqcBY//69aeWQIqbZjlT
Ru3dYPQDdAXSaaKE4UJ1Zg8RfFakwXehV86Dp5fWq5DhSz+ikKriti6Kt0LNEJQ1
HWnwGoQSdsyHZ+aKkA7LIkY+Dbjb8P0SpAMzxqEX7lZTiNwMddo4Puvteycs1aO4
JJwnWtiMoqFg+fR6epXzFgQUeMDGWf2osoJ+nZRgO9nMLqDYKy8i57oaTjLWR66v
k0y0Ac4IIe0uQSgYzSc2sKVLYp13citQ6LMvoOoymSR0GQggHCNmM/VIZ2tbL24J
b8kdLMwNCaYnJmd2tXMxNaL1jsVOWGLQKCXDIEI7pUt9NPrZMwNnndINzU6ah91D
J+2u7As6b1QOR1T1mXRcBTS14cv+CxLhoNZs7lcSVbHUXj+etj5dq5cN1mWmoVB/
rS9uNYZLb8jbNxDjpu2KClzYMbxwy3uM6NURnvmtVXJR/ZRXg2Wu8QNUAPTZ72hc
T7R2UKncBuPi7Q/QIXr5b1slBYIQNRSVj3dT53O7Oxc1NcAZjb1cP1xlXj+crT5g
rORBRtcHPognJymwGQUu0SBTWhMvHVX6THdDlnBz/g1RjhnQYeY8+WneomGb2xjo
52GVqeDABA1jtyp520IL9HgEe0HLiOyBuOshLmxc/5MXuE+CDm7KdKLbKTFL//+s
yFa4AO8pP8rE8IR9K7HVOaQ5WlnLJ5TgmjYAKMwxDu5pDvE2NprhjQYobRvBlRqH
t4aZat32eppX7RV4OCnWEiiDzKrm8w5MmJ2lBLOIACpdujY3UPkpUdERALAE8wyv
G9YTD+I8KDU6rxTVSRIJEVCE7W8lTddPi4sC6T8RLRi4htEfxRB0+ACoULvZajsn
v7p18zwZcyFPUTmww5pgyn6fahO9NwaoV8lCJBA/9mTmvXNtLDGEE+inYUPMOevj
0tvRJfbAZMyPHZsdNd/lwgHY0vRUxe52chLiP+0T8DoIBPbP4kL+cKX5eJGZKCIw
90F+Rg7qOCgp8lKi4tPrnQhOHpbEaLFkWqbUzRnnTsB3MQiSCu9Q0YUOJIDf3Wr8
cCvI+XEvU7YdjZ4Uc+91enHAdbpF4SdL/QlB0bjl1SU8LZ3hb7sk0hUeqDObVVik
nT7kItOF9j9aCrGLHAmUqAeH4frDEEZwrigjOeY+mmq+rlcmYw0nWqvatC0bhyi1
bj8pIDVVepBHjvOR7arIRNY7aPa740iSo7dSaae/kWazQpTGt4TRug102Vl4j7/y
dz3QFkZCnmy36XoTCSKBp9ZybwVOiIijXOFosiI3eE+TERptddRdJBTOrp5pYmdR
gyYSjnl6mjvkb+tSIqO9H+iK3xXNGuuc8nZcxhzzREDDDmQYNFN7gLWabUFEMN58
7TA2z20QJlPK4GpkEHA/lHBzjG2Bn7Nj2pEktGEuBXIqhvUO/uBb64K4cLc5vGqP
qZSRkmtc5L8/uc5bDok5thduH86RAy6UIEecjdGfm77pdyHHt1iDF50nYO0zRp3l
vgx+YORNpyRGEbwQixx42U9QfmuLhTr3y/9m02lRPw4G4fBe3PBB8G/9cJrcHyhb
FnXQwvlEUBBol2QrKfZlVsp+XS20REWvZMSLXwFhgqykwzECU7krcqqT+ezCUVpt
oJkp9lskBRrjMO0lEtF44o4XiUpyElGLi568oFoF4uZBMUGHK5WcxgN4wo51b+dp
wdZ7wOPjAYoRyLSQRRZWp4vI4WTvKj3S2KDWYq0pCJZFQjRdb2gBTaE62MMd99HB
jq+pfLV1GLhwnzsWJPtOe6az7te5lyKDpIlR8qNmEbPKjR5CjphcGkzVVAMVPczo
9R6bclXYp50Lp0bjF5CL3HANMaGZ0ooRqbtFtB/M3g7342eevZ4XTt4ljRt5S6FN
9xJuntNkzr0BTlw5HFbMpjxK62csh4qsenVQ9lrcMPoc3N4j+NiteRYCizGbBKJq
wZOIJrTIM2ud5Nqo7D5dupWEhjwT2PVYoZg7ec/VdXNBKcu/srNbyQ3d/xHSuhoQ
hgvSBV27/JZMEsJR4k/CUi6g/Js3boB939MXX0tSMlXlJiK2pn8m5qPpRy0nas0c
7+i+eMU2tbhfIpiIo2W+jd0oqzDJ93i77U4fh5hz1+l9rktunc06jJmfO0MAkD0c
Z1ZUGEgP4gVk87s4OTyRRrvY7T1LS1O0P33RBppVYAkvsSkCTVnf0yIrYgGUErr6
Qwrj9/JqzxIhHXBxImfZPT91CSoKQL0gL3jSgKUoXhxRSN41DwcnqlGFrTanyueR
sabrbT+C2EQJuTwtQuaXG7hQFtlQDQuja77XNpzQfhPhQuqEgH69a+foSZcovx6I
XLv7SH5zPC0mZPkoo7ImLX5eORhjYtf2Lg/RHh0Nakr8e7dwvQzMSMiO96RpArE+
AP42Zvvn8iBMGw9dEgjm1KlRDQ5Nc7O5QdfC3x4myk6crwwrTBwiwsTO+CDfKtkl
j/s+hltWkKOHhfOz1y/hvtQMHecwXRlJdoWD0i72salG4AjcHj+usvhkZM+L41Ib
H1ENB+omJ4Eqm8QJfF1G2CmI5Hm0an3R3qc3MyiAx7z6VKPzEkKBpWm0CUPUryd+
HptBgJPJ8dmGExPVHfDAWpqx215TkPkUZ91pweO+GNq7Ht55+VdSQL08NBUIi9QU
10/8iCdrk9ZcgvLueh+cw5myzmi5pkDMu3uaGDUhDm1PU/2aYo7AE+DpoRbmYddB
CcdUPyMSDgryaAAwbImue714ZMiCOYlk/dKE4pIbp+5txBKCX1TBDFhxAsz42KDj
bHbSZOTQQxK/c7g5NYkGEc5pbxoNKkdBr7LrGGA7k7uJ1N05ovIumBB4y+DZWdvB
/SVQjsa8UHnw5HXUQCg85mblPGWZfsPABizvDAVwXiYljnA77XOlgco8qokVI6vu
KnVx0BDrUxFEvvkibn/kZBXQHQXd6RZV8KbAVPXl1+I0hOr/02S5MqsdIFvyqI+1
mMOPlsm0l85vJo5cX18Vrk635jZ1pfwAyaxYt3EKmE9b/EdADrP5PeQ4mCN5Tuqe
lAYy+Paqc1ENXrvI4r3igkC4T4SoYINK7wTVNbNUsV+Q8diFd4RcJwDzToMYn5HE
hMDILuHZjXfNqtmM/IH94gXvs4sD69g56dKwNxuTnJAC8mqqrLQQiY0tMbcxHXqu
7G1c37iINBwdDNDh6oh2QXnFZ0GiFSvOVJ9C6mLaDXWMiaFl0qc77vwlzMzmKdnX
HEKGp/m2TFDOsXaa4emsrfg76L/2QfToBAQiYwvI/kU9PpV4gMQS1OLLodxcAFRC
R2TFsUISE+dLBWwjp9wlNnXZzP/70HwClqkAGprRFa7WPpMCOCR+PrXBomjXc/tn
rlovLgBKWftHM20oGuO7R13V7x1/gUtExd/xKUpZu3cqVJJLmbeycK/3X5vPhDin
Ne87Fx1zWcRYxxc6aer15gAGuIqWRA8Gy0iLuUVgEyzzMlBcWtlBmk6rqE4bd6Bu
ULM5j3rSE9+e+xIPdB5d10D+iWwh56+68Ua5FexXpdc/BgZ5IhgM3QxncwBfd2ka
wsrpOLnd6ig5/lhEq5v/IPv7ofAbGadfzsN49Oiyn2YkX9+1EZjP4xot7HoqPql3
F2+sFsSh/6EDB1ItiYET2Q6wHamqt9o5IPA4bvWNHMhz2vSN3QdJPG1DIzjKYKMZ
OLdOgpxslLVC0DQk9eAAavfMEn8Vnk3pWC4243TRNFkCfdqt57N5CFBqiVsfYZw7
g6v8Ie3k3l2A+p5XDS4j3dTwLS9kVj06YA/fX8/eaMy8buvoBhzYqkecG7qZJ/cJ
kkUijKQCHEn5gojDnQdw4ZldD+n+c5EEaZN3jo9EZkt0TiR0oy7LkdKrG09qFyB6
ls6itCO2h5fEHjr3C1scdL9788qXZ1KX0R1H0WLZM+v1QW5jhz0Gcao4TyvPkDsr
/IW8T+1H5363P3iY3kZKAWJYgJCX3tdMu9Xe+TzOygavYGHJePqh0QILbJOD/YIF
uev/dF6ZrYA5yjvH4SzesfCjvW6109f7iEFrAQKQAJ0y/gl6XizsweVTvH4N3YbN
Xn/BZKRdJGOylvdMYgXLHUUdTDGpDwcdL/om/sZg9cJs4YTozp23GOVtJCjKSF3x
CpOCv9g3i1GUNMtXdReK67gUhHDPmMrwRponxiByugFuW1PewvDMS75Dh/uObeTF
rLj3oQYUeG0c9JY36BFfemXS/zcx/t+YIgiP/AracSXYy3ef0cbAVKg4EMyCTuIk
IdgIdKPxx8pYpp6lZlatNkHhi8M4gkW1T5+20TYJsK5+8ChHplHauiO0dvBqqHY+
GIt6MkjZypGNMuUPjJi0rlDJfjSQuQTdRslIIpj89sssM0jboyDKSyTG34jBUScj
oJnMJL1u7Ee9cGnQcRz3PwbOjHIfKuJQr8RJ6b/QcsNY9JFFNhUJlwBPMq+VsMTG
RMepbeAVQwstB2qmp2kvkGFIGW/v29uMBJTeZG4M9+EndMwUr6vkKfO9mtbmmOjK
towkcA8nSdcbImCdYxV4djORIruev6bLGhj9ByKU9bZH9pLIGY9oof2Vd0prixKF
dqrWys8nNW8RmoJdfITHy1cUXKv8jrwI0Zgc529G6YurTgtFp7cHc0J9qD08fJN8
DrvXttRiS1QmKcVZT3J0IEtWiPJmacJBTecYnkPsm06MYXXBLzeuG7wqps6f/JjM
WmnrbQC1XZm7Z91eRZGSs08LDeQxZYoOSKMxdGdYKP0v1olDdYnMRnK2yz4JpZ+n
rG0MYSfu3gdJyWuChUV1QByDizciMC9DCHoXHLdeM/LZcGjuhL15S8q80Xnmg2rI
3PLi+HZo2bARoE4EcRjt0a+BGsa1AbOUes8t5wc6ACOoIc2M4+T0uzBRRe/+06GY
xNBceC/JGky5LkVmlNod6vCO5QDeL4f7JBqnDOjyuLlGCMI5RGuGkvWo1hlfVum6
TnHbcBzfIemaa5XPVOvILROEYQNf1RtLILHfwHHBn5KyrlrsUGFE84s7uGfZj9jy
a/wihMRluQ2ObhoCrdpqmgjLfG9yPrfFlz/AdLNyyIKF2OpxapyEJwBAjWaq7xsM
UgjWwLern8t9Ks0T2skzUlWDdzqTCFFH4L5mX9CFyfbqIM3hLfX9Vp6UZjMkLN1f
KvWfi2+4EpWmwhAoXKSbo2SxkIgL6BAGX/9KA54y7R8Qcyo9UGDU7ZXWNWLQ0MPb
stdhiNa9YjczCtpi2SH/do9Rbzcg9Qz0PGb4oJLe/mP3dYUZ7vCsqST/32Ic4tr+
cyB9NAdpAtiochJ/y5LNlZRki7CLEJdmPL3MQXNZWBK+EHtSwS+kyoaxD+GPWdWJ
bhChyDqlH8tzftWVg6hKAcjVzy3uB9a8Qu1VEUtqmIJBmNX/wCTKyiCaBiZPHoJS
3sEZkUagL4eGtH+QypWO35Isy7JO3SeSra4vITUCHcV/k11ULbVwsk/Wf1Eg3cn0
FT4I65ON1T+xYw0XYebKeSuz9RF86A0MeC4VfGiulT4vQoFX2ItWBTC2YAvISqK8
PqcBed5d41NAemqVbSCN5fQDEUKW+E33M3u5dJHwvtIYAL34axs7WogS3yyiLfah
szV6sQzlM5QZ+WPy1UAxy5bzcwAjiuZdqgvXdVFfnXcu4LSPO0l8PYGsEdplgGWB
+bMZfvI+1vT8L+Msr6UnwTgOQjurFy/WW4pLCv0rTeIEG2RoHNxn3vk4AK2lXWZ6
gwP8tGW8zttCzuLtHP0Sir696/EcymLWIiBPY3MjbO8R6JF1mTvbghhm1ea9V6pY
3mywoIH8oVJdBnmNRhw1Xxnny7hiaKhVOxd5dGDxPXvnjeepKT3EIIoITr6jwXLN
J86sTuB4vp/0ok7OjExKcfkGd1Fhd71PYnUJSs6DbcbNXJxZVwmp6BD7TbEGMcq9
dRO0JNodGJZFvPCj5/oO+q0UnkxBg7IklOzYi1qE08T/IwdAW9Zd1pHXsQ/V4Ff6
NhyPYSWukfv0RJ1Ou1uaHPKcyg3iOLvolI3TsCJ57w63q4onvtR4Yxs97X2Cvwtl
Jdmem2oQKA+HZ5BcRA3YT7vzhl+ncC6xtYo16eHJ/BArE6I+FqoKQ/XUk8ljdXU3
Qhzw8fLFJIvF3ex1JkCBdv5jM0asGefKJQK8TNjqMwPtoq74v0w8rbUFYI0NfU9e
ZDG63xwEYbcdOi8wYQNG8M3+jHMP2L3xhvrTnkUh85bIlV32NbctJZTCqQqO0bSm
xh4O94WBHA91FrWU2vK2Zy/r8GigEJQKvwGw68rAkBUccu3NsILqOTEGR9BekQbE
Dn5tRi6hnSKhqXGEuZMEzOXR2+/ceILySeDfA6kPeW4xSnkzqW4he2NyqJ1x2Dva
W5dYi4BT6bLt+TBMicKD24YqRjOxbv0RF4YzjwB5FkMsnfITL77ZVW8MKDCjGOQ4
PFmviexpfroLnHPR0wh6qKjntRhLea1sF7F3HbWSHbJckW39uVsjEE+efxJFuZx0
XsA4Pch9p1j5RszMSyKQG3i1mrxIQTtH830OoS1I+egbs1faobP/fRPfHehKML0h
GaCIFAAGCv62XF0ihzc6QKj3N1FqkFvOnjb24Ah+hL3AlHiOQTlwA72hqnn5gCPZ
ALukkcjZdqh/Mz55FmYXUS+oKK6dNPKr7luYNaR5oSynZYWZ866Azu3g+fDERjhC
6avd3J1DsP+hIm1Znk1HGsi/tVEAfEBcpkGV0NxVYwLQCLZt1TXCveo+QUNLkOSB
ne5uzkL2BsGadjCyOsLZMw28PvVA/GE+Bq01o0Rb6UqHutyxFP26Yptp0iAKO8ou
ZoIGBmZ7bm9XRjBzSp33LrKMZrpdH9fGEJrV5KdHrOF+zv2IZZ8Vnyt1ylrwjGNx
DTxYmeIuQA9ln0G6FOu8UO7zErl63rJ2yXwRyAAILvCC1VlmfLPMO3sSUjPgGNoW
77AKHLFxbhxYIwKpfD1tzNmOgxJURrXLQ5RYrU/URlbxde2yJqAKIqxsjXsxpxYC
AzsZYYVl693SgxXl35NQp92y07HuwXuv1fgk4cJ8kIr4fWhoPPvFDQZfypqVA/fR
aXcTPGtwVctSdfQw79VT0Cvo7Z1bI8FayfFdowvwJvQTCqw4mt3Ml5+xmMprhY8F
OBfDihOSkuSVTJczMA4ZqXLxHxwhyzp9KCa++FPtUCbSH0GwMIch1OiEVQSuRxks
PP7Z4lJhRHLswPli/Lw8kVG+IOyld0Qf6Mxf73d/pXxbOMmD16cb5LNbBMvobnbM
u2v5u99vC9ICtuHL48my7Fca5qLSzNU+iX69QNPgoHFus7Xxnlc8UEYsPe9fBvfi
kulP1gQ450S8Zfr8VGT7rlGHpyY7tvlBJJp6czVWhwb8InIEWf/niCa/txuP6iGh
KxdIvqj3vSh8CrcXvchpi1v52Gt0/AEvym+CynOdLKxeFX6W4Bs+carAjPXSiCTm
DClLlJE8oTq1Ttx1jgVtkm4OTpAazrlUIXmxSz7wO4RGtamza9xLrp+fy7ZByWo7
Snc0wZHekA0obl/jqAQ8W4N0W3DOp2yqMiID1QMJWtRK9r+E/I1pvP7zyC6VsC7z
woY+RCZrAHJHFKQhPwVYjSwJ66eE0kGW4BcqBhliaHFBVg5m/6XlV5uvbdi0Fomf
0eimGgFGV7SoO3OGpNt6YlRbFYUelAPjKOwqoKT6QPVM/zkbA04outKryiP4LlPJ
JYXUjT+xpdDE9jPWTuDi9LC07pmfncJ0DE/KI7RypHCZtkC57zHPDdSHygtjpEhU
iqd1YTTQ6WLEFSQ8Ecc3PR3UwGLp/zZfIHTkHEZ836983IIFGSn/7bLe/ccS0Zd/
q14To5BIi0jsmWwOHkDhjeaSV7DllIZ+oVVEsegMiPTuyrmIKSC4o/fu8q/gQ+q/
LWSF3XGPQhw5Io3ngikebc3lW4tibm+jc9ZAYHnRPcpaVoocHYnnHUKNz/7N2WNN
MC4xCtSek2XW0opjah3Wj7ewTSAMs3g/3qwettgTY3jgILgUrV88j/ASnZv42iZ0
YugjczzkhVkyA2eoApYBCnobTrrGGjgreA//93g6efCmoKGIENxfmF6w9TIAgUnd
ydMREyg4Wsmzkwn4jInmb5MDIzES9B0TRs3m1Oy3zZDYNWIfIqY0UHISHt7JU5aS
1IYZZV3mKLub4EW6vGE+slOREN5pGsL14YKskGMqxiQJnPh67FpbEZMc/knOTBHP
B+xJSChvLR4q/8Zbn34EQmc6gK196DtWY48whYNkHM6vCfG1qjAScPnXFveepRBg
bmvvquyraq0E8TSspchD4WQCru/7JiGFdxID4gLstaNGEU1X9zNfToD6jN3aRlnU
UT+Ykq+2sZ1yzE/MD7ciwQjxEBrcjsKqzqs7cZ94vEoRpiTWLyMyjDnx27olmlvT
OGOXhfqqrRvL8F11GuIdkvwChAS1+KwSz0JQNMrfw6WUAss6K+YicqLW85GztuGV
ea7lnYEs3LLGWAK2242AW8eOQJi/Pu438+RdAf99sVvXiDCL3UZ2GIfquXp3RsBv
X0PcSgg3vL7vohwSw8eRdLEHb+gKsYE3gsYXPrFg+0GBvcCTO3mtqWx8jhLZD7M2
TGmuV7aT4eQIHcG0U0ADJKCzjNAqb3/xR0hHaOzJuQqLxe6y8eO6mhlkDsumWpwQ
F3iRGRJR7n8VJi2fOJ4IsIczYWCBtdhg0LQL3XEiGj5NlEyPLiuz2JLCwlGXV3+e
Qm0cjYxxvhuUIJA0VOyY5evP1+5Z2REtjN+o/WVkwAfW52u3WVjo5s/WLY+heoif
vxkssddpK9jwK2KJ3ocYi8nAUCHk/ZWdLjhjwmgdhoGfPjYMfMATVPbiNwzzabjT
dB36UW6wHDKBB92j0mWMTuLJtLOZg9YbxK7dMObc4GnRB1gZFB/FpNSDJYN3hruS
YinazCRG5H6AR+LsztEmx/1z4WEoYRYBQKxlT3XADpjM3TITq5K2tY8ADMUpyVBe
98XrtNu4Y1O1a+6ESLR5FKQartMSZ6p+PTs/Sv7/fsWcL5Ju/NMlGhZylbK+rrtS
Me2wL2kgFrR+RjBL1KVOtGWo+5peCQvJOdKDWe1F7bcYQe39y2YcQ5TEBIw0guUr
0e0dsGlDuWIAo2qz0z2+05zG3l/6shxLiP3dgAj8gB+DES+3HoQW2fgn5Kf03SoX
cHcc2zkUL6SGZwtVtK/I7b+I9bOwnOYOLpF1Hzvw2sY0oycGKQ7NMRRyezw397e9
SuLW+zkQzl56QtT4K503gWcYRK+cEDAJgf1y1P94rYk5fDsKz4OMF6WirikWmUwg
VTjyPrnW94fM/rZUwzjaku4n+b6sureSMVGdPT6r8l7jI5fpdSpMOdcZKjQq6zn7
SCT+86vqzDmbjJrL4JtoOt1Zmoxl2IbE3wVrS+xbnrevqm5zqFm3Z1hcIWtqlW+E
48KPwNd8Mo+w8Sp9KjKYpz22vV+bMEb7GMK+DG6790+Qo5z2+4I21r9rdPVGHspj
cpb7tXnLIXasoTzz7/LknnIBnS9i7Ta7B0pHnPxQJJG6b/F4najDzvY3l9tg/+uZ
trtTL7vGwhnHVCWUcJMWVbuJy2gNkFSJ41SqxmUs1NAlwdh901gPD9SfDO7ct8iG
iSYXkPiiXxgDmk1phME3BNj0leVSlnihKeSi04karvkGu9anEYBJvb+kZvtwUmnr
ifeFUHXurVqm+afhAsF6vyQDcoibrud670SY3oiRLlWdHGdvoyrxw3wxH8oCi7xh
EoVGFZdBaayzpSNdN1d0ZaLG/BBLnCp9KVF/7gj8C43umIexrnqcZwsJWc90PicE
f9gfF0f0nq3xWP3hiD69S4mZy6z3H1a1o+JIRGIb8WYi1p/mxuj6qzLjbtgG4/e8
k+AbzQ6wzaJ1eoFtBzATyBSFvgEzrUwcZafrcNmz0CGJQp0r0wctxGjrFjsD14rd
WFhuWiHSyderd4+Lnq9cnp37I/5dsJcjYTyjPQsCDsbVWfY2dRiFlrU5iGA7VUUP
/SMeeGnGGaD5VYu6Q/Z2wOK1jISUu4QEP5hmUkVyvkh/F3CNb4pSdeFU4eSG6F9Z
T4LHselb+eLCA2mKA/7NrAr04Z50BsJphSO37ROl7kNuhs5DlckOBgE2igH3mf1i
3aSf0zhlioa3Eh4J+kG4jNIYI/2geE4sAu9EfVO1JUqLPY1i5MG2HuEXl9i7cOgd
hUnXuOQmNoLz2cP+X9ykADvg0s2DsZXkoj7zftW7Cn+zZlve5XSaer49W/g+Ga+H
aH/Y+v3LxhhcIbhRITbv6CC9QExKT30lreT7VbnQNg6IiRpPLa/Vv4lYmvKjFI9+
E8vU3/uPsIfvqS4Qn25w5/gPl2xkxYgmi7cyl2eFS86ZMa5AE2y+ouVWhY2vhTTl
82OttUpH0Idmw6T/5FoUCF2O1JdiIpDyCnT0ebYHvmWy0+F4hrBPDdhbcOfZoVYy
uVE3xHTjCBXBBsD7HpFWs1s3shTkI9I/i4Wgmj6LlrjexObBs+cWVq9mQxcG/rkw
vVJO/ZNgpRWWBkMf92m7XyhYTDKWOVLPemMOcjS8oM3IiF7b1RCnM/KhufNe75mA
MRuCxHj/gG7uwk43DF5A9fs31eU1kJx9oRM5+0INUeXJoKvaHtC3RPO46t9zZPWC
Ze8a7UzT/c0C+9QYRwXonE7GHZcqk0Bc8FKQvMpmraKxM3htAsGN3YMq11tEVi6D
NHKkUamzMm1QlGGsd1zDvgNEjx/q4S7LreWmt7yCv7wqPXmPrkvSTQD8OgqgO9lQ
XdmpZT2QG9AD0ABsLiayXbbkxTzRsuNmxfp8LngvLHljeKPd9agXZ1AhkO+y8ORa
3JsalONkbez5oWnZFB/z8fLmkKagVt3XMpIeNQsVKX6c5Do9Zrwdl+SyM1t5dT1i
3BuDxRzJCWp7XP4TrdrkfENIvcAeuFvykPYfk9GGemJAL0NHsXXeW9Lj+/Lc/hD3
dkNijJg4yn7NZN5PcA+jX+1lzVeSsVBNwKtOsbCxYzHbRV9iZf6e/Eou1wpxzx/6
VozTf1ue1cP7kjStcfkNfKce9DBJkfvQI71DVBGtn6zESKk9otWLt5a72JjgwSh+
3X4QtnpKOWjoTkaIiTh8X4HQpoQdOoKsyV+l0Aat3Dq79CZEd8h2eLti+un2jkug
ymETyz91koedgRUOORBj/XgPVKv+4PkkrcOtyX5UtyIjKsTZ9j8MxofWljCX4UvH
qr/kWHZzx+xURITgi8LB7P3FA+TNalo9P80WvmI1NAsupoMFwU7e+pUcNXLgxrcV
rQXsWFeQ3kAH6unZzogwNoUHBt9KuGuh2s+WmF8T0N/3aJnFYdFau6DwQVBUF0oB
6bPhZGZOyloCoh5SR1aMs/Fu9bHra9+mftA5CT09V24GCdpEFxApOjmE7Zdf/RIB
0USiK2GaY7/Q3ToiVQNJkyRCGoQIENvLc1HhZZXrXjI7O03gaCHx++WiIHVXdFhh
k6hsvue5nLj3ydMwViYUl1GaSf5cVGt0c3cspxYJzbbAjNz/2Rgh6cyX3caw9rZG
BDDsKZDCal16RVOpKJOfT+Mrkh8cRZ/x7Fbdc5CBDqdHGw8OQ88mdblMqEY35cVu
IOIq0GSry7ix4C3nlTwfsi9DwdtZ9EdYzCb3WY/BuYJu6YMXHfj9fI7hr+kpppnl
I+fmTbbSia+uE4fr2hWvaTGJ2Pz3/aVbTyjz01jSgJPyGD2FmxyIQ4om/z79aX3e
+Ty0X52+VxFjCOM3QuzZKt3nMcFEtmy9EpSpI1ORBcNevWYr7987YKm9W4+w1odd
7hcPRK0KW0ISAoRTyqDQdVM4P3wAvyJlPmLonAwy3Z34UEzv7uaL6yVKI5csb7k9
qfr7kGhlpZPkwETyVHfZYXc9soCGE/R3SxGcn6qnMMDT5FmQqCHCw3aUD5ejOFYi
VlICCjIVALj0Ejh13yRQU6mtcJmR4Iqd+tgepSdF80esDtyvrK0vBED4xUkuV1em
Fqmdxk9MFy5H3FJ6b6KpVeDu0pSKZBbNEl32husLkJI9leXcbM0NBT1L8E5NSqvZ
1HltgUci68J/ch2X8/TGxa3h2Cyju4HzfSJTQayGpQ6ujewtfCfhdn4R+wqReiat
2UgodUXmc5CI7iB39ZHls+7lMY45nvyr/10ZBO85nXL9GF9UP2ScUXQw8oF8Bzhs
bfsQDzJyUeyA8gi48VJISEtmMpkPqpwxXkkJ5N+TR8UXl+tV7sWI9G+NkK2CGpqg
QjmM/MIba1vpY3WEdVgccON/O2WzGeK95Ey1rX4706rytPmQyHQ1Lml02Kyg0PrL
R8OS1Ftlk/S5ryMRbZ1O6Oec0kn1vznaJjMdgcxU+jIV5ApPSr6Ims5B053mqis9
TGZUshHL31jlZArZDILg9EizkwcLDOcmkKpOcWfCe/7SzVPcWbg5ypSjc0rty2rw
IBEdCODSHj0SIWP+ObZBbtmE29fUAM316hR7UKHoz2cXOGXDvSD7DupL1764eDGW
vQf8dYcJIkPx9f/n01M6XNi1jG63q7aZXrXmbALqMTuDaBkakdl0dWPYsAU6Bq4E
cPPyVbuGI2GZHOeQyZGwZixbkVQegfq+hnwP/0BfW1TBTz4NkNG97Chxh2GqIV4g
StvMP4stNntIt/6DO1FNdtdfRmMNxDeVD+LWPGGHDMUh2GoigVyvKDM5KlU1+5FP
8MiF8eL+TLietGwIO7vuw+skWUNsmXmWZqfPryNb9YMWng7mVHTKWQ6BT0nbGWlf
HhNUesfeBH5P9WoyCA3Dljd6PkkHOr224/0WPqtAAsOIpSyXH8doscrcpXrAGmPM
EYBNYVPMFSRGxj7b9rbG2MksbVbONuxa00MYl9elQrix/jp0wAw/ThWFKM/mA5Fu
9JubdqxHBdYPRIFfXpS5n9y8KZTQqZ5QQAg9lMMdeYoTsdImT+Ffn0NNI0Kko2eP
3yL6Go0RGeyLEhACaj0g+MTNfx2Waq+5qNNasz0uP+LKbj+PgrXZDTt9D2CgNXxo
5p5n3fTMTEMm/Ti+2Y6JY8Bi6Zd7nJflXZAYc0ihaQTKIoHbEzqQeL6VWI5WtRIW
P+KVdaLY+o43Z5IDg3CcmvG9D0PVjg3spgRA0rNilGEiHGyFr/g8lM/5zAKQIxq/
fykiZ0cHYxrRGKVIRb3ZI6R/qyhWy4RaAZEiBUsB70u78gddg0FKEl7LmZHQPi1+
bp6oqV3Dahv6fWvx02LSMjEktNUqY5FGgNjOOme4AqV/JDgl4IHfJDMtkhFJaBpr
oC99n463e8qRAriZ/zbZTu32ejSaEvEJlaewIbRrlRADAk80nbjyUKLDu9Z/HwS+
SN50twRJr+OQ0QrMfvTA82iL1iHEumvnaAwYlkyBnhLSZaCXoeslwbLhxEeLcrwk
SG+j7lW8zKxcdY+Y2JVOLHujoyXTIOebSNJgfhotYlTE0URKB2k5yMjCLZECvDpA
Zgd/Nuql+IaLYn2MlDcWzEFhS4EaYqjFaEgpMCUVgGb8aUIzCIUDelF5T1jUJa3R
28L3OJ9RA//GLVlIB5/aP4AsmbAoh4bMdSR9S/y6tO8GyaIRZpW/qOuNeXWjegua
45NDNZO8sKkwtIO3pQ9JRfttO4ncX/HnaRCKg/OqvWStBamd0PBV0odQHru5H637
MM4SP84cjGfDHufVOkwTvr0jkSe5lwoK4tZt+NxjU7LNwU5Muja4Ha6AUOZ2WdXJ
dw83DWrnMURlvFNLkl4yWjyQ3j3jIdY2CtfAjJEuoyQUNTJEDndmyZbZf0YSlh2x
W9/57In8BMwMJik3VBM0beTwXhnI48JJzF611qb3oP7kBNlwYCXINsTtwip6wP67
CgF0paWYGkjRzZq41q6EnWjiphRVf2y6b3v8s4W8SX0zitqtKgazHqNiNn/dKVLP
OJaTDfP1DyJbTwCHwjtBtW81wwPpWKwZUHZm1wFc375J0gPe7tcqL1ReLDTqIzBD
XOSf3WtZeJUiNqUC53fvNOuvdSldMMd6b4avDhEwJbK4OBfkrz0kKxCOhiJsSaUC
pld9TMXIYCevWjSs20MjCCQ0pU687OjujX/1D3l/lOq96WC60d7uuSnxiAyJMdV9
3oA97gBFeqRNRb45+lIhhuWF6qdX51h0CPBSAPD6MCNXs62Q+TC5qxE2ANOXkrr/
2Rh7w++tBUNkKd9/0ZeRFQT/y1cpzHMYlhKP9epH+4J60m3PQsDaqTpl4uLtffW3
0jDS4xvKqxM5JLKXXWldjQO8ENpa5QTuAzRDllYJgJg3j2dqO7Sq3DnZXIycYdVZ
fz1gksztqVLd75XnIxhuhSS8okpuDeOus/Z7XMs9cKcPkppK9OY7mAPNg0Ti6E2x
UFP32sfvKqusyL10F70DyUCQ1ENRJwQU3BGKYB6bAavsszYetHPsz7hehM+lVVe2
sldWN4k+7ruXze3pK0sW/6xhbShlwg0la5wKJzQy6L+8AGf/1cuKogOrHE4hDIMB
OjmdgxI4tK+qTqBnpkwQZUy0hS63GdGUolRXPA9duUCUESlq0MJko70fbUyVZcqf
8qxpD/blbL3nSI6HE826hNopij3UUzCFJijKCy+Ehsv40nP1GXub/gim//j+ddi2
jxXdrl1DO3XIYGpxrzxTH/KqUfVE7SaA30DcpH0HddyAVCZgE/mmwQolDKEer43G
G4xlIx0d5eaqAQMuuFfcaGQFLz6QHhpPQP5zeH+HTuquNqo5pwuGg4lYgbW8jIh1
xuco6nR23VQ1mBtOngGGsD87F2FgFI2SQYqeSyjG1YDlkXPVSacgsw+metBa94Qr
WtAEzDj0HQYp89aMtHdye9Nr6pO+xiT+JPzzra3ZoECbWD+E7XAfz8dbxuy0ZmoB
Ki+y6V1wuOtdMvMPysHcnbINsWRSOaTk3/fX4+Yk1XEeYbK1FGW+pLRuY9QBN9nh
9s7Xzcl6ACTaaMLGReerF/FANyQ3u/UoZn7pwSvig3MMVKXKOi3bs1y1JdyJXaJK
CYidK+rkLlgN2t2R8mUMSrOwBfiyQsQcfCxUpADPyz6DK2oP2+4j74fT5xiMlYFk
hxXjwVVRQK4bFzax12RnucGmTYw8Bm3vyfk5E8JdcQerBzEbM0OqWo898FZTmdR/
QOKLO+ysFrEc6AsHPhHZcozgBKsRvAq/jlWvuQqKAjj5G8uMh6+RF7g4R7MG/rWC
c/pQr3Y0eoTvjVNfx/jh3yiXPFyYX5rPZPd6eXQi9JJxtAouMzCyAWhmshsCFuHK
dclRfbKik6QlLxTnqtwTF3qBAyGoAOhkOCkzQP0AMKQDSiv44gmZBwE5LXscn80u
gJ0U7aHNPnBD83V6UzpsNKD1+X0fYWsttjmolcolc6NlnQhm2GMcvE2AopH4nVHG
hfmJAbseV6hT9r8O6pBco8OPv79XRCbhxEkoGn/vLKDXd4NId3tg9xCf+G2P3k0b
kNdxmMSMT+Z/vxiwBJnzE9iic7VRH/w2D0nRLNSHYkl/BbX4aDDI5VIfOItSpwsV
VQxOSC39syVgZHnx/6bgIIEFWg/QYyi5oWc3zytDispqYy7Ft6zHjHt2AVV6R034
G8ntMo4qMtyTu4sS7KSzjUQUWsCDX1cgnbm3UaVCNFFK9CywmgdM1UE4+lEoLLHm
9XlINI1fDsaGE8FXwvpclQ5XOpSBsoK2/OYKQpDQloEl8C8MUzMpFvnmzm3uhjQ6
RgV2KM9zpqN6nvMZ6MyGqKIRJPd1nZI0vyTbbMb8QcC/yK0L7z9faDiEe57uPMDv
x027kZfxr4ugbrF1Q2Oej05cEz1G6ctcJQmfGFBNfN96ECX6ajgPP67DEwJT97+4
C1/aK3rhH+qtR1mNi5j/5vlGSRhKkGcgeb9tLbEWSZ3xyVzMSwqm9LloZiDEvUZ5
PUtRBjUDtilE/G4+H1UvfJl7vEDymX3waviCxnJcMLo58oOoD3Et5w+3UUnBS6JL
tyOQoX1HMgOKU4k+S1wmyIxIqm7+vX4aZt9dlgqWKUHdpvmEdTSK8Wj6zba18f02
iSEK87FGs3OhuLUXKMMbv7qMuEJHDIkQBUhqu/jLyViCbrp4Yf4DwSyuCd1MT1JO
hJSx77nv7dhxaKsJ9unyfUntAweK812WEu982cYk+EhPx70hkPgVEZoGQZIrECYs
SZB1qF6MUVNFBksRYNlhh/ttKN2xk8ABHPowPSIXtfgr7hFl0Zbv/9diNVUS7FAr
lxwP1lC7kd+1HJXvqq6PaAKG0+wF2md6TVQHDk+iz7r8j8u+3Bis1vOBEkvCYy7P
QjnJm+ThhW6FAtNo35XOUQmEQ34MT/wkL2dpBAqxTkN6iHl7a/3NUCOT0Kk5Ebii
nh0FbW5D1jSXaX4/x1cQBYsXvKM1m9ZyJlcedE2NflBN49l/zfmP9wXI2KxGV5Yn
lKHfoAkXZsPcTv49YPiW/55VSAU3i/BpXsFXXnSKpfwuYx/cWRdqrS2u1rGlf/Hp
Xx59gjmu6Wa+JY4gFeNM6d6iFb66JcxQ4wWPJJw32txSC7iJ2IKHeGQDnrNLoRs6
VnjO0BskBc1zlSb6EF8t4SMVRflTBGMCP7VkEs8qexoEJZOuBA/2IRcc1pMZa/qN
EyQOGZijaHlQOBFG9ZoWCFeF4RqSbtCbOId1BjIp+pKSBV3lRnbx6i6aIyWb5JV3
L52GwZA5nrbvEYiC4RikJejjEKXW96DR5oG3BNZlacsMkNnYGn/zNHiPXqOsOzKf
a5jKvnzb6TKs6nDhiUkFFYkOg3zhhzcVA6nuyFZqVeusSz2KNetxWb4REWw55FLw
qPGzuT53VeKGB/aUPG/NZWI2Bf7xxK7oEAxjuOqUqX5pk2HZu30hJCx7gQcsb1dW
o7OoDnxFTbdHurnl0f1AmoHejktjMSaRe43n3tfd2rOr7UARDMcSbhk0r53ffip1
XuzRNfyntCt23ZYfD/XuZl0d2H5kz6t4OU9HwrFU41gzQEFpo8GxWKrCE9MstWea
MQzEwcRwjSDMGEhqARG0CEmJw8tZ4k5ke39ulnoJK9air0sKeO5z6B7StMdaXXZM
Zq2ghWVv6wRSiP5VwSNKZTXogltTez22eyVh7Im6Yzk6sC8zbQfqkOgvs0ZHKd3M
CG14jGhE2bFUzNn487fvg+3kgPxMY90xEJIrkGiW8ZrcpMH3kfvT1CCkDN8aAYSu
JT7U5PUX4h7FVfhVQAmowpPyUcgKQyVRCT2F2vu617tUevoFbkxjeaFq573sgCZk
NrFg5RdkSN+NMlbKTSkbJij81ixAj6YxU6dbNgISQ7fBdq0SrEy37n8wtx3Ai71P
9jaY2m2Z4AuiQ0w/eeFksa9yAyHkJvY4yOVi6vaxOe9Tkb4Vc45GaM8nwn8tLxHi
VgZTvPQNwJpK9WlOjdYq6AzVHnJEVrUqmBXEqU2f2wwp9+7Y+LqqELcY56aa7h1t
kgFCCuVN7H/X043HDTJNJQrLKwnBiuGtE8XpGF6bAWwXRpnV04V+ZekxHuvA2teH
QtWvplZnUdEq4FaOsDl/JXKJcaygC+cnCFBttaE70HGzf0QaDr6wi73b9fLIQ0s4
se3kOQcRpCzoHu/75UbGfKP99+bdbOcCousycholHagjXJJp/fIa1ta1LTINZwYx
c8D7pAYq2uiJGFQqjzB7i23h/T1UUQ2Cd+pKKmVnGiX0tOeADXpNnKdBk4PPR8EZ
8pHdrAsJK+KNiFTUhR/RU9Ja5Ej1fki6m6wc9vc5u52ws4tpvT4tyo4sNxOZgKyQ
QNLkD8ZhHE8K1XriVqJouD9pEd51jqkYZeRBetkRV8qQTVfxYp1Rcv2+AnGh/iOc
lnTk/72AstPFnagkDIbODGv1VqmBoW0/2yfcvb07wJm4EI9m/yJovG9kTVfQKn1I
552C2S4FlckXQltdltqRhgGDP1A3B9+9jUiUvDYGinAznLQceALe9NxgwS9D8OYF
AEcHjX+V1T/mS1DPuB/EGbq8KiQrAjQUKAiJ4uXZrmmt3YhYpZT6cVlZ9N3+4NyE
UtJIKxwGU7qlNK+ZgFHfeTQAjDacOKZdS9LNdG9XpgTM9zaeAOBhBSpIktNrlPP/
6r30q/yG4c6X+FDq2buggi550PySVEhpKg+/woQ8Txtrlz01Wjq9BR26qWwQMfEc
HmOAfXqXxmT09TzhAb9PSuVW472fnB7MQtYJiddXy5QvGT/SlkWXEf2+wlBrLYg4
BTidvOhpDba9dS3ooUYKHRuRj1fJq//Jzh6VdFdZBB31vSXcdGlys5ObSIaMQHHm
seIbY3XsZDDDd4v1Ju+7tBBlbpax/Vl9L8LDRl8B9Nael8ScSiXjXZXcXBvxJQBN
f1Un7mkPnDKG/nLqNp8yMvKB4GodGa7oTmj7/UYD0QM2APqQU5/+Fx1IDsGdglbe
WJZLCh5PBnn9RdJmPkzo87GI1ElxOYGa2tAhjO3KoSHdrpemWjjk+6gqOHFxj+jq
dgT5jnqkAvFCUmy35K14ACnTuqrqdV/KsoFuDfVWsXKTKQGgaaMDhvASP8dcdp8j
qFyXOtAMuANJ5K80r+jiA36oDAdBK9+jbPH4RzX+8VwX/BB5mPxc7MxMzQgplyyp
hIvsjnbFGryiF/e5L00Bf+EA4EoDDHBsFiLN5k1Ztqqy8f9Gf0Nm5ITlBYaOodnl
lwvXeR+TLph9Z0ZHzNvVv6azyAoI1wN8pko2E9yP7qPFTe8LQiJHv+ZP0hMxZTVW
YxdHv63aMiNQP9clSdORbA6VsWmVLlgXesKepRX3KzLfJ0ay0yyKdusgJboY6eED
nzdBjPeVZ360crmSFTODxHrQ0dqSSV6qCbRaBfYf9jBdp4G4+7D0elt324W8wjVK
RaXWWbquLfxD/NJWTrWFqppfM4eLpa4ydXuiRsi30gmNIk9OSzpfeHRDq2OBox8t
vd/s4K1dpBCRsET8hvoa5694gQS/BfEIbbjBTQmR7r8gCVEvMxNsAhJfZuHvW0pf
1/Mj7fXCkoCx9Mrd6aNOg4QX1ySA6tkcLYulgFDe9vM3tEK9MWnU0LTaEjDBQ1EB
J+7zvx/bQ1ih/BIG8qYVYl+rsa1p0Z9cMommdtDNpbY9+nZpgMtiB55Qj3NFI/9Z
iO/J+nOnN3TovUXRtslUp6HkpreNlLk/2SIMbxmnCJeHRKTHvhtL0mIhylruCywJ
soZEeu+hBDdnTCGG81r5mZhpMQyRXxNJemWiHqkZX4boykkJ5D8EpEU9OC9z1wLA
YJ4Scca+3ljA6kGqfKrU1pkRiKFMsJWB5sjc//L0DorMIamQ2iwdL1oJtX4zCGJc
5sTRShNAv7BmlkGaTlDmCgekmgYVsMEtV3Be+q2Hp1vo84ebKoi6Gal3WRTDyviJ
SR790QFXlRflnX0ydmrJ7PSf1R80QGI6wqwRb//pdWldUZqAzh5mOuncb1FWkgEV
wuMkGVzBqGl0RnBxqrg6ckp62aNzCg9Um9SNU8syxHyGKuPdS4V7/ZdZLSt59ZEg
QllPbEYkKJsIyUrq68RdYtlLOrwu1S1BU2v1LwNH0N2Hep7iVuW6Tq5aiF8gj2YG
tD3yBkIUO6jdNsdr9Ak2HiUf42b4DaEONHUwVIs4T76GghAxNtGrQ9rK9up8CMRn
J00I9KZ8C59/DH6M0ld3x0bRKX8OLv5RXRzjThQ9XD7HpGqzChXifoxsiW3wwYNK
foe9nX3lvWIm0OotGMwHmYxP2t+qwh1YHDEKr8HulziYdxKkjm6PT7b2/e/KYDxr
2b6cTIq/Q/8DvxI59Lr1IafN9jbsLjlmLLG+le/Myv0jyL/WjvXTy9brUHK90UEO
uKhRTbejXyDFTuhf93LAik3LBdhsss7LzGZbqgvuzJ/2+RK1wZfmcoct6IV5I8Lh
j75GVqh92+4wuDLlcOdxCqErxXFTTKl7t8/SEyTWxR0jjAcY8+fX0S8NWQ/DuHbf
9ORqai2UCNSe8s4o2HSgPfmsOrMYnwnMnkSfk6yOUkPocnFF/2JPm0TxW5hYS55f
OMqGPxe9coyMSTF9RFEHhsxmOrP12QrJVSXAXqbuDnqJ/joKcIGToRWbEfGSh+16
YhJ47m2aPsw/y3rJd0k/D34z4VljwW36KqL0QVgJYLPrVokHjRGeKJd8NifCCh+e
oSFEqFP01w4eZ+1W+0wlSw+UM+9bViwzTUlFW7B2CdS/ioOlyTwaHS25b2TFDucb
VPvMo8iMb0bnw5SLwDUzkgrr0OqeomJYmJbIbFPvC2mPGEhDOBTT7J0rD6AIBeTH
oDgyWA1qU58aQ27TlsMvOjaoSjHL3ePFG12PBXO6gMnE7pI9QNAReE6s+TbmSDL2
DEYd0oomqAyVy1qEZZwA2McAbPnJy/kschiTdefpqWfIo+qGDZNTbNVLFnVPFDNZ
BeJv1nfSHWpAWjZ3r3XVN9XKpXfSOEE7IuYNycJopPdSGHekeldcXUO4pL9uHwlr
P8Ez6MFmQuqZVe9tYc18nPmtIKWNi9gj4VNuXmCgAkP2Y26Kt32ehZiT6VHAiSjd
774CASjxySSlGuwMX7fGhFCfZ7A2wRXpwx0tGK5ew8ZR2cnEEEw3Asc0j6E0TToQ
0/QA3WpcDx8OiARyHhlEb9qEBF74xPR7o1u4JyErNXf3T/GkJPqQ2nx1xt+xtThl
k65Cc0ZHXcSu+M+hmaXyS60QRz/m1xIxeU9Rtk3CHCX+18gMnxFU6BDhy/BKjlY6
3epBtQ5z5y01xbiD6qWeAqJloqnr5qFEQRiCc+/Poy7upAzKoHedS/NGpS52HqH3
q8TOZ6UCIqtvpDABmliMGrKPPAR5NL4jM9i2wpWuRFDY/x/l3y8gIzepjlEkHwU2
MynzSU4RzE5npneXi6l9LhQw2rlY1fg5/603Rh0UDk33u7IG/PgeS3laQhD50u/2
s6QljsnsgdZ41A8QzVRtnXGa1V6N8T6p53isnYWBStq+Bk8nHiovARuHSMFoJecE
QBOd6SFdh7VM+J83R1P/xy5r8b8GEZJTWQbLEeD9i9kE/61oxNUx+pB0L40WY+oS
TOqzkoW0MhvhUkwyDOX1702R4E+ZJGCvbwLJKq/rcpPagwP8R2FaoMKcTD2pvqvd
8XCBY1ssou6qB0vVzKa6vWtZoAnve8JTEf/d8UNeYS5YiJS/4Ws0RM5uXparlV7d
az1noHRAhiXndc5lfca2xW+IssY3q9gTwmPzjUzw6ZSLPhyqsgRxZVVhASe1puE/
J69tnG7HRmuIA+/6F56VsDzB77cqzmORdtoAiJLjifnRM3S245iGJ57had6zu8U3
fGbCaciH8l8dOKiC4GsB/22BM8We/faqQ36YM7sw5aeGYrtfkNg+KiVvKCalPSFt
m6vRlGoYI78jGc7KpHvfTv524eunidUqM1HhGDAcFs9rmXGC6Kxb31TO3s1Oa1+X
CGgpi0o2WLOe/Z2eyOYvm57JZHfNGyGAUm0x3Y3/HGqD1Sr0LJS36WXAr8zCUszy
kJsdQaS+FkCnlTLKkLjYCrTP6fmB9PGMLvp16Vb3SsFauyDC50z1KapyYYSgzC4P
TWOiNY9z3m8de1nbwQWiVuIASIkzpd3+GiSaLRcBjk5YP06A75IEzJW7mF764yhG
J/h7Ajv27El2DP27H/X5bMSro8PD/lKqcwxqTB/KT3zWtDQDXXhK4GQwoxQjHsfd
wwyfAf0Le7UTET6oJfGmy+YEseEP+VTWwI2A+pjPpmd37jtz7PWEycAXmcdHPjD2
rQpUnIw1JvtfwepfH1vuKFiECnLu+INCAJC1ABIBA//no9fMwX+zyoTUmAFeRTdQ
3bhaYpTDcs/a5K99rpsIM1ZeCvkOxw5pV41KECJuCjBHzu5CDghht818lQlo5XWF
OgbZ2oaTJRzSvr4vo0kaQt4iayNyA1TKPx3HKjhdmvZeZxvRikvj6D8R05yDt+KF
j1vauH8P47M6Lmb+X0T3uRKfYgNNWVmu3XxZjmQ+LP7zLcnxGx6jgdHREpnH76HP
qBfT6XmmnNTji5Hu0ScawSya10otFc9vemsANPn8Uzujtf04rmpY/7EM5ZmIvqUe
tHccNIHKHKszQVPrZislf0mMb3DDmHQJjcGyOChfv/g8LBGj3eHehE7cKoDJhY6z
Iy4EqWauNH45Hfmx8nJHm0p6O6P+G30KKF3ca8BlhJC7INOLR9ODEXfwNOSb85xg
TRSyypAeR3wGDinypfjUvUX3qwpLpmKFG/yu55odld1NEXkneRcbE81b0357JuBN
kf2sJHDZE4cwhY6cfBwn0FK8uQrFu8X7UGMVjpnzz0uncG5DqCZz6FESElHUNAwz
gkuKfB6zUl6lLHdV/V5aZmQsNhRE2q7f4CZSYBHfMQBSTQPPGHJDdBeVO7YerAfW
EjtLMxfkI4newvwPxxhxbC+5RDKj9zpKGjbvwoayAEDgiZT2RZAnqNqVPvWn9ONr
ehZIKmHW4LO5aE468m8fbB+yfywMpzJtu5RQA6AAB3DFGb6zCFMcrJPZ5NeOGvbL
i/fi+HvDD6QwHp/FkYUFNnYqNk6ugialc/ElXQdhrxL+fLHPbuxVvt+9GeE8RWgq
hTLGjZdciggMRQSa2QfLvP9OEKheVCPM0523VbGzU783qrOIe93FyoOD3v7KSFi/
yvinGQkcCZAsRENUoEf8DDv3bqzoY5pEwm99Saf5YVNIiOOccF2LhOL6pLE6Akfo
jqRfHnPK6BzVonL9QUA/uMMHBsoTD3j2xWcnnr70vTzB39xjn0ypFddmVu5t9ejG
zWZjWhl1ziXZvsyff4YuPiLvOHJo/I6RAu77gP5H4/SkmX6R61VRZ6f6jtQ8QLuo
uAV1pRsGjJ147U3/p8Np3FZXAHKTnFYG7iwtb6u+t7eOtezCzJegfpNkyt8qSQ5e
pWt3R6YKP1p0NX3EbPZtZ2EKo3+ftEw6fsh8yMa/Ul+xuqOoNvIJB/YMKDja+zlo
qC3LXGdJIsWBaGEJVuiq73u7s3qFkVGhbxy9f3D+AbU4Y3LMY51w3rw7If7X7+j6
J5kBMqD73WZi3StTCJ4A5vechwVTIMCYSt7P4WAH2SeSITGtv+DeyAb4GaYZ6QiV
XkDZrPcgxvDAO2aQBiTAC7SrO+BYiAKzTxusyu55QJry7Rz4BfdOXVOZWVXsTvCS
ALhurqiDGXnDcTq0R2e3wU3u0jxQEwctEyofkvYlJl1DEqS1xc7ab8KdWRffhYr+
ivuokxnptsx4HLmjqM9ezwRfipG82J8NdmBe3syQQmRF+uVfmvXHpuqmKo/wYYLB
0erIUeqr/68+qiJHkvz3uss/cr9tLLXVEI874BlCI1hxRL8VMolrlKQuatZxCLvO
26jjnDaAy7giLHsVxA2Bj4Fu+nYTB7amcGkrWogcAn17mBjqYhrTEN4srXLbECxE
6irXauUZU0Fo12DTfjtNoHQ7o1nlR2Zn8RaJYqiqM8kirq9tkSlEYAu6KV0HI7z/
2ipwAB+R2aN9ecopOh8EcSEardABfysHxYL6TYuCo8Nhk1hjyXnsneC8TvndsN+D
GEbY5ZnbJALQQwlx02zaV3m731tPN7J+srvddJ0kW+iYM2mFVffFJraNRSFAPwXu
pmnzxTG+ihw5hCBKYPhtdIbbgowQEeCNmQRXbRKkzHJIvQsbvOFuWW2H2hVnqSub
gLKdf/d07Y2uZ6JdhX5qgkM3NL/TCe7kNZLWACPFPg6lCaFg/mg7KHbeTdCnTvBV
VdfQ6ult26c4hKJ4oNaZYdqSp8UeuWNz3LjWpft5LoZJ3EW2hnHyEeuGEseKTeLW
svuxSnOVtFi7yvPTscw0qrEmDipbUNcDZ96OpAdw6724F4rhDwQ8Ut4KDX/dFUvK
foqWBeyTmwqRvAvKfSlAx91T3qZZNe1Y9nDX4qKxrgPMZa5gbf4+8JdYNLUeajnx
ejzNsu2xwN02rNdvVo1j150MPi49l4fC/CCgeQA0+ZbDjK+MMaSl8vczWNtmBCXF
Nwk0Wkqq4I4FpxzRFIuScR2TH1NyVePtt3TWYit1lAHrS+586JK2E6tzXbcKfwjG
UtRGYbpevjWYVoP9x5XrHqutMKoru2A7LocP583gb103qpGhTwrJRTsFMAOtmZEE
i68aggIQ1bkyJhTm/um6hppx3yg8dI7TuAqkkpbSlSAoOMMDF4+Sx7B74x4Bvw08
5vDNIxdIH50gQsPzjlrdoedcZQ8sjKm0ywFzfDM/qLkgLFOoIjl/hh2AmN7RlwLo
so6qaoWKAOMglPsd8v71J8ppPFZ2X4+mSchvarNpsjNEBWv8o77Jm/WtwAT2gCuU
beGnPB2wOhCOlzfCJA9+fMRvrd+BtKWoW3UmEohY/UdYx09vDK4qzamtzWbD+zNf
Q0LtTlH1LPFJXJ4iRsjgJDgkeN/+vMetrqoBjDfjsj/jrQqWazF8nddsaGNud9zs
nX/J4+OFsrVI87hBeTplt1xiPv4SjU9+NlrzHtIEUDL4ISsXfjLvzUgBgk/BCBaU
XnhnXPL0mYpTaJ0zJPBVEPZb2xITH/u+UfRRp31XeWVO46rcQHTMdqNWmXq09sER
p5eO3Vu29HZrwl4jNhkhrD3soTzCVDQ0JUpHEjMhJgasvmtlboqcKwzQ9IeocEar
8abjir61JYspxthggYWSEncrVVf1OldkPa+nIJtRBJKv5eZXuCGM/+cFfpBUnuMW
AHoyv42h1Q7DVKIzfAvgR/io5dcTcFvWwdrAkewUQySBVE1q/tPwmLYoek86msl2
SbhX/s/16N/I+9qCE3mwCIL4/aFYOWdgLDM80sbxMXboVhfGR4qzUqhFLAAOB8rO
GYbM6SR2jH4q75BJw6gHcmq0Knyks98GmVs5WMW03sCP6C6enSSDOxGc7xxV6ZdD
CXcg/HLyyINKo9W7pC9l7yikk1zmF+l3MZ4befZBdQ1I8s2O6eG3FUZwn01IllKM
D7qH1DrAcf7IdhIBTuJrqxjqHsbkFJcOXHGcpv9n3RLeyODFWyCUcMFVcTbSLXHH
iAX5gNVgRHB0KoetLDHrbaQoyzlc5o8Ddjq2f/NClvQMW5GRbCDm4j8+fxPN6zBx
cbcErVdBvCMjvjrP8u5F8JXwBqLXuVnFkVLBwCTmInfeYbZETQ7HavvRJHR833tn
2iSd3a8ARx/CSSyDbDAdRxEqvjs1p2i2LTxnmtKweKPssRvZ2NUnbVfbSrrIaBEQ
WfdruRhzM7TiYfK+8/yEdAi15nr6fMEX6j7c15KRXX59Sus6Y+VBw1VtO4jHxryQ
zjFxJk78tYx9A8MNCNcNK0RvihZ7hTtlncbJIfC/7rTDGPuIj6+gsWSPleCIIlgC
eSLBZc4uDq8+ppySLvf3hUfGs2fRW+V/pfIvbMKebZEa0OpUAZB7njMjWoBQB6y5
r82XkcHBH74oclLAtTaEC+dX9oIYHNuQ0cb3V7GGqK9Y47L5GZ9VqAAQ0kqgOPQi
uZL5cmXd4zHvjVsOybMl46zIigLfvqBkyjXwx67clV9Il4Pzv1iyCu5/SG3LkYd5
tzsJrNFsjrmkrPd71kggw2CtVDkDGDhZMPlBMbAEn5Sxp/zL5PAfYozyzGBRAemd
knPFiNmtLRKxWxPYGDlzObssr3cufXRN7pcrWunSN7wj54bdY+qAGVetT2umV88v
p/XITgO6pYkdUr0gZNFctWGuqOIMcXev7fNSIkJdHknBoD5bcjFZjrKbNxACfnSh
eIYOuFjGP8RxHX1lDJbYKp3zoDMcMB2ix2mXxq/t9dGxguK9XE49cFV7AZ2I4T8A
KOudf/re8UKw4xYGDL44Jw7qldxF1/7X6tlO7/a5qE0vOuUXXumZBDZZawPgEYhV
l40oznJQ+TzxLKG0Bs7ul3drIkKBoUpt0/N1Iqs94vENgtEBTqimfGC30Ym/+u6P
GQe1Y4VXmJerIevO/W39l1BzXuszgTplvc1bkMcHnNAvdHtp0y+D4vofbVrqYP+z
JEbHdl17WV2Z8e4U9yS7HREuhR9fvWIGLNa/TUgMnUbuzkhtgE0xftWTTtCrUDnm
sCN/Jx7dexr0ar+/EqhFaGnZ9I2hu+jbnvO+s1X6JBDZqRfRVadz5fATd5tpZjKG
VPBqO7aRsf9g7AoqbbrrTt3ene7nFqDOQLQOYpnVXt3qDZvFmuc1OTJ/92vbXTip
XhhFye1hNH8AfBgWPsEfZk/OltnKM+70actnZXsRWND1WePqzKVKmeyZyY2gmP8o
6gXjPzlP2bTwnWnRwPL9xXEpPb7zAsItDCcf/VTqwa/fIvUMhb3AEncfCG7zjMHb
Pd75+1mH1czkArCP8mDB9onNmnWEdcT8Wd82jeb/2AoYNN7wMP8foFDNPe8tYq/e
VDBMNNDuOfoyHwj0YZeNgR5/KM95w+7BpqW1NAv0ieILhQmsEbtbSn1TUx43j4DO
ZioRJZHvL57/qtxj5+ueqxcHW/dke7rbGbK3SllX/WK/5FZKISAKrbhnOJVGtSKa
tk2qZzmjcsNicVnrJLhlfmTzZeUV3DZh5g5bMDuoxZdi2EZNotXONzJVYvUI27IU
Heqg+N7ePjTgmzwtBk7TdJPpLtHy7ngCG0ee9fOUegDP/UfEa0neqBn4uJ1ti8wr
kLQNFUKLeIx2JXpvWOzkZn5/W7OJVVNB13CALnwTmU4fel8/9/A4H8gfhEWM6Xnw
HoQfHcbgeBjPn+Hqu1t4hyegEeleBWgUXY3iYiIxXByQqcpuK2AlOyPeX6UZLo6r
uvoCpXCf7dFK9Ms5QQewcEuBJqFMBqLMRlpwGX5agN34thVPedkP757kij0b6THZ
c5TI8B3I+DolcCF3Qw0ligwvEOVLZKnJUAgNxe7JTZ71FY6jsvDedW1boVuV/6kL
aID4kQgYuVKsFQinhhz04QwGgKk7cByAzH8lukB5e4Q4VGkPgXPgvd2gNsQb6vvh
9b+eijPKQ4BQHpCgIKr28RNRvPsI7ciAWX3FP31UP0Qbta0+WtmfvyUfgFiGC47/
01EAmD1tBW4sFa7scB+vRixlZKqgEFAIZ2nfEdE0lzuqvosHNQoKQncSmnB6INd3
81r1NxUzxa9TRQ0YoHKeznmkUIWW9e/zE1V7ZRhn2730PfNeWLmDJorckp22Gx8U
EmAKqgMVqxp6qV2HbpJUEyWkPBepRL9eHT7WHIvbVvRimO0v/54BOACdjBVrHsUH
19pDLrPqOVvut+e3D46LgFfUJPc2yQHlZxXsA2bB0UmTUNBDs/Ad508/wSRs3FhM
Z+d7bqQMjJ28Mxh4qJ6YGcv/vLte2c31aQZddt0BUUaB0t8F+L21CkrgrkRpTC4C
DCx65Be/3ZR2cRWRxpzksuGa8/Ydg3eFvAYYTpWVA4uz4ZTgdAVc5KEaPBd6cKBT
DqH+1lVBL/17vxHX9c57xdej9+y2G4+AoJOHp7g3+DxP9pb+Vadn3qjJGJL636Ld
JpzrkO4xlT0rNoxYpwro4eUwroyVsaMWf9If5i5Stz0rlaBfstApApkAYFTMETlq
z3qE557u8sPLG5ldVFboavpOP5kFMnGj7nw/4qmiZ+uwMO+PoAN3PziBKo23OfUb
EF1uISWQWtzin/T+0/eyDWoe0AGx/KLmdI6Eg5IbZOMaPQf3lVMQbSKo9qgF7OTh
pCp6WCG+3yV4Qheyc+lCayuw1LKWF7Ab1GPFcK4iZ3mJq4yB/fUUVwfM25e5I0q4
gwyvTAESt3g0T4ubSYYVjvauMbT4qkBihAtawcNs5RFcQFQv3Q3mZPMNwa6FBgAI
iJhU2fokQ3zhjZpIq87StQrPzqrMvQmw/yyjaaaCZMIKPj7z8cAlJuppcmCRAQQJ
3vY9WyMPtcCBpIC9JR5zicl7UBmJD0t2Ms16Um1SNUbkI6E5GjTSFtfUjlGq772d
ZFSdDSBFZEhGrjJXKF03f1+3OeZqp5ex6jgJ1vpo1pBtOWvkcelbBwUMDssgR4U5
jWpuQpV2Q3GgrNjNlW4tNX9nK9DbktViQrjfYWUjhyWl8gJPEgUWoHVxPbObEnHn
ugHPO04SSZnfPJ+z9oDz3gSSycobEjpscAeECkFpKVWfMvU1Tig0dtgd/YUO86Gj
tTAOXVUr+w/w0D8d+2pGONmqLkG4Q3IDR4UjHeGj5mgbxxsKA65NtXs8qK6p0zXu
qnjS4tMYYcr77lY3Z/f3GtZBbvJxHpP53G2qqTex/9hZphIk1sey/lvcDAp1Z5o7
BlZV+lzpJo1MIfH/sIUnerkwo3R777d9A2yFJJ0tPz72s20Y2Yl7LvO4XkkIkXA8
SiIxKOd/pXs69Mjt0EN58o7Kfk8lAfEp/XgG/alW4zK9Y/aBnqcwxPy5IejsGfzl
lCm/5DHE5wDkdGUPcdzrM8RUvtOIPF4wlEPzoz9UPSqZSImw0bzUiEIwh6Itjqn4
Oa7M621Lqh1KP+ys0+VJijA8hVppioHuljPZnlwdGi1rBtvxySgX4efQo2khVvSi
AC00Rsj7CFCnH3zW/wgLBfUZ+ln+2MEjrXr61uHzT8e72hadsQHqF5ZhUppeLujl
n3XpY7cX34qzxBkjyz2k94zAgq4A+FD/tIUhuGOI4gO4glZaqCFIE1Jzi+LyT2tx
3IbH9qneAYZFmJuVgKXeXBr00Pf/bpdUeYc7R2gMS9TV9f83FGasnEvbAHPxQban
OrG+G/z/SEU3r6TIT4athopjIsgGmQp8sGN26gNlonnsZYP2GDUxNS3su12V4IR1
FJARqD8WMfccTJ8M+DgN/IEUATbDNoIPhFRDzemN9uS5/iHpqvWN47IuO7FV2X0W
c6TLaV50TqV6WlaJbrR7CKXapKHvzsV8T0EGfWBJoEte4GTKKqYgf8LH7AcbE9lf
ZII1FRlsb9mcib42BJcrxMKOzAiAH5q+YEpsxmnZaN802gIELQG/0rXLUKVBHFTA
ZizKzswjgmqPSSRL55rV90SQv5UMO3eRZ5VpiaI8jkCqgSiQ6AFVK9CpTMjcYYbE
9HCcVlfHX1TgX9ZEltE/Ozupa/xl4Qios2OSSPoq+9r7TDeUdXad92MUA+Vs/ZaA
KeYfS0nvnrw6NBctZCnN71p6vK5GjGtAKz/1GPhiNdz0acw+zcla2gK5vUfnj0KZ
i53ztSzT1DLSDOV18yIfPayxLSXCLmgo2OfDm7ULfEGgkuFcQB3j5Vcbre1mzVxY
RjjQ6WIwUc7KxJVqitB8ldXJhLCeKFYDSadDyeNyDbAHL3EMTc7RpMV3Kh2ATpkO
RwqhdIFcjuu0Qwra6z6xwghsWHS1OCxeGBDDKk2ASueDa7+dyj+hqpQ2En9zUnkA
RP5YWkC568X4WqPH/UNtc9kZCZmi7FbpXMADIEZdp2HQgmq2EruibWu5nqtP07CW
xVSyre/fbGNXI9e4xoA3RoHELenKzieB2x4z7/YMBUmzJkRXAgEvYMb7jAZH0XdU
FvT9FjNEZ3+Pl9IV2zqfxvd57KZ9chYQAygWlpaeDdkjVRYCHHBOgFQyrwsRG7v9
mQIRpSPD7E30x3rBnq/wYjeyh/BndQknN+ZdW/4v8rEi6lbFnq4GBxJ27qPd6BDH
eJMAXOXysEkv246b5nEMyIB3s7WS7QBWrEDuuDlAzNSlmKYy1eHVUabnWJytWouj
q2ZNo3mqjDbIOK1twufBhdU8e7B7OmCK1YtRoqFTbGp6eEWSXztZKXijVdIG9nmM
eMVSEgR0G0KmIiOWFPrsv/HRl9zD179SkNBQzGz7fYa4UHb0Ot/Up8dZlOcVS7W6
6rJGroDaU84RyrKmYtsoNfT9qdQ+ufiD8TFtwMQPu/W3TSmz101aUuaPeyUg6Vah
6ow1MaENnNZ2ZCH2vMVx1wswspFksv+FDKKUx4TEmAXTrsHeRTHe9qdgTFKGPPj0
LIBeJ1AeymuP4Lm52+s5JpaJGyD3WJ6Ny6CSXt1Z302xWZDfgrugg3KWDGIWaSOi
svwZWW59nVpvwtChSsFe0NBJQZXcGDxifmAedAo0D7eCxveDnmGrBYBLf05o9BQ9
SrJN5Sh1iaN1UH15kM65yqavbSPa+SHZRHE5xgjZyEEG5LvLpsOn0piZ6wfMY7+5
tYzRKeco8yQ3jDpy2d9OynZ2+wJ7zDc5vg+uarSB1GAZ88uBLr2111MK2+SlWcPt
w6iovrnmHoROmSrPg7BsZJ5wzbOd1yvdEiSRsWRXs9AXo/p8cCuOw5Q9nSGAtg1N
zUnnZtWORMJl/5lyWA2C7ZrY5EM6z6WTGcT9+MyZbs1j7u+qFtUVqZbpiyBzbtKS
GmiERSCJO4aMeA40+LFsCdzcLU20o/IKRvuuRp70m0H/Pj3+LQrkiaTQxsYvBaXT
9lwJ/jKqD4aoQHTkAidI91igwV03sVMRRm5RbmwMN2p3rfrdtMdls0FRzxD+xAvW
VoUFqIssydPW2WR92EjpywTFooTqufoDJh4NHo3Ocqclkqw3fb5dkEQSUJZhYVBe
SLlvBZcLX4tfuPoI9fGW3x2EPFOejMhiOgT2loxN5xCp+gLHvRBW5TSqYhHqnpRy
phkQ2kmzi4fxWGsslKQfFZy/cNyLCw9NQO63XgR86NZ4acKdWj6XYvy96qwYnMtn
4Sq/hqMoireNQC/K3qzilhEOARdKM+tFgLL4ZqQW0FJrQAXjbXQEv+APlgK98m4U
1E+BPfIiv3mXpIuMyMNvktHJ/H+BMqs34SHKH/t0QECxPt/MH5hNWuVm9jts9986
pO1ixk3VzCBtOhgBDJ5mFnNLQXnw7vojWyTX0nkugylEJyVeKkGgsfeVfttsHHlu
XGjXPjIsJBcsYCFoZNfqjXIhTN3j/rI+cv6bUmeDZc4by/2N7bLulwdV11RDtwoz
Wm9l0t1mM2xoPwzQOSNsVDuIG2SJqcQYZJRyjK/7WFfi88BJhfOlHg5Tba8pZhpC
2xH3I0HaKIIobwblvQiwEwefa+8JM8ThDISiLsvBVE4+SEVSjyKKOFjvjCEXuBPb
LKCt2lu848l1LBLkJ/kOzGtC5gzl46M0mvn+gO+fm55Fyghjl1VsJRuL9Wbnb8CI
uIU8JH2ZbpFat0840mPcr0I4mS80P/s1JbBnydpL7C0tgQYxleqibthVf4LhtCmQ
F6S5sWR9mTMCWv7ed0K7j2blpsZpd9q7Pxelqs6gdt3lFGSRPPDinpQ0EUU5E7lL
9wL3svpYme9hNAULYHpUH2/9epCjR6YuwlFo/PrwLjikeHbZPoyQwtfpCirMfZih
tfYbkjT+byrC8SvaUm2uDkF0idjdHDZIeee8CwwWmEqS/nL4o44w88Fpn5Iu1Rin
+CELGGEWZ3tU8HN7jEia/B7XDwNdackNEfRdXy7PzL1yo9hvRSzcVGbFBoy3R0XS
neCRiz3qk071hMycq57GJvQEnLZrpEV5zH5h7DtqBM23Pj+uo3UckRJWieXDOxY/
+AC8cqAmux6cuu3IrlzHlfMF9WNah8qkn8i+WNrR34UFJhri1FSmBdtsg7WocWQp
rA2gfcQpclyw4uHoKC7lqVrBQ1z45HaKn4ypn8+jybohRQwF7YN4m+O+Fy2oWozW
KsaUHJaFb1vy3DjedB1v6Ua+MZSqHDo8x+nquuPELnWJlmnpp0xPum9mbTovIgGJ
AG/aZ37INAS0kx+lcDbPUJmTrwUTDmJZ1fA4iWxXFLrVZDEAcNdxkcPHxT2600qN
RFxuA9qlpq4PFNoX9Cr9VfpuJ2FGhLUF+JPtfQb+MRp4p7MctO7cl+eW1t0l1iIY
XKcwcCb3KQDVE6ZmL1GLEXrQuG+wtsJUdKbm0WuBLaRzN1ziMp0Si9IZ/ugB++Oa
dEyKAfv0EV3gGMDrhx5s2XZfW35zYArnRgfiGqxZnArHr/UW04H9O7IQ/oYnNJKM
wXEPTnWc/GizFXrL2ykmpVE8QThph+murzNOgRHJU4Vwh7aJwCBngb71VJnu+6u1
Cmx78fMyg+4KC6Dv/S1WL2fXqBYwibH/2oTgfPLGGsNO9cOMuSnOrnvz/sPsfKT9
K8osccPBBpu/Mf0d8nUkIe3Z6ORxIWpeyDearY8sEUgi9ZMmwjzWdw5PTbkIyjQi
ZIuzV0VI7A7Ti3Jf6d5izUgyZre+pjN9eZ/Slqn4lZiB0BEcHpPIYwrnbL1Odvcj
XWe3IplyOd91yZUOQrZuK+01IGBwZtT9fvNZ4q8nnREhWSP6i+KJGDdELSjyQnTb
zMZ4PLibFKpMXl/W6ZKer1irlUpPx3IitFw2lIJ+MZ2+VJpk5eRncPv8X+V74CiY
iYZbaTwPQXEbhhu0FW13LczmNTL46PonNZdWMjlK9D0AciDao3ELzFPrfYCO4BfG
1DKOEk7A5gokO89P+nT0AvScYCklsN08LJ0RDqYcF379jzR7DePrIgww3u662/DV
CW7I5StAzxTlFS4Opxcab4l9K/b0EDE8ipRZCDqhzMwwHBq2aVDXg80XsNEVUJaS
+MexVQ4eZ3kYhb5kgkbwLEocVdkgVQEBrpp5RIX3z4mH9qA8VYqcpXYj6oU6VDH1
6AsNQQRZKcsbaVcA8GxN9akL2YTuSA6qaNHUMBMjeODmjT4SD2+mgVgry1sH5ERv
SR8Cq3C7ztY0CnKgsngNEpV0NZD/fH40RWoOECPCkt1fFvOkt63bhlLRRHIoZ246
fTtwFlr2WWM6qpbHN6IylGdEkvFAbogfjcPfw8kwEsdrRnOEA16JUaeGXbrBX3rN
43c0zFlTu09tVJwD1mcrfQoydkoTHqNKvZBjFoT+HL8YErMkqhwvPLv3J3UB8i0b
rYR8vhVrKxLyYFyNzZpSjU4W4R6UG4udJ0d+qIzNHexG2IYeUQC69tQNbjyCJtra
Zh7l6x1G7NmA4aRGHDEvXhkasJ1g1j0hBgrRBXgJuV+2bPinkb5ywi2iTymnordh
2lIe+g///16HLjo10XQlQWSmRoxi5oN7FXvh8RljKPfBC8Axsw1NEkTyKEN7YvwM
Ebtipum5kekCB20pNAoId/H9VWAOdRcAdiS8L2SbcwZY6y4ism2isyDe3gDeTZlH
cE+34gJxWkA7eVM02oXh67W0F8fc7d1Hq2PwALs4dF8UsJZfbjzRAV2AQJTG1QXq
NXlDfKh7Wuw1n99ieyhMpuvHh5AZdSR3tsNMWVQkJ4Mb1OnKUFD2teLAMXMgnJ3F
/Kj8Y+e/liWu2uNilTzbkzVZjafqdNvtOTcO8L+LM1lOI4tldVyLPSzjDdVMLOWs
RUGqk/mO1Gv2TogIqnpXnBGp+6Gt3oP4s+gYcluuxMAffT7NLvPxcqejRQdTixAi
y/+t/MD2g6Iw1u2Bp3nYBjRsKODiyBTrJkcY96F3/Jls7hWIlCTghVcgbk6ujXZ9
2C0RKaOVl3Q4Zd6WFw4FkshaZbIFd21AC/uSmNwy6jCR+PWKNihQoL5MqpS+JI8V
u8PtK5psbv1JvvEqg+fkWYsT55FrKdSDITiCIs0NBAt4CUv17G5WZgYzAsDj20TA
8ireLtLCwGl6WfmKMixUJ9ntC4pFKjPXW1L4ZGSb5UGcTXO9aNjfAbs4gmHXmbs4
nm6AS8USEcC1TJ7jg+PjyGRvx64mIFqIRws8zmkHTN97OWFdfaOHbINAENVAtMuJ
xW8voIw7xOtYZkFd7yzR1ANBdX1wu5mc+Xla9t9brkoSE9u9khiZ1mKdt80TDulf
HK6CnOMrlypMa37QLaVMP3v6/KvyFL/SS43jtRGfosV188R39FiAmeCvc7Hb0kMQ
WBvo83oBALNxlf9mf9M82wON8HxSfRrJlEUDE5LSU4/YpYKX4hGm5wPhGpZdnlhw
kRqeN1XWpUnqDLwy8njfp5CsgRmbv6v2u915PH8hlYuj79mF+DsUzSD6p0z1Xoh8
BGapCHgXFWsfsnCbcP68wYoV1NtApg3CX64+T1R/3wkBZdQnjd5EaL2iJW12Jc0g
nEBHZfKCJ34gmaeMwI6F2/+9H67LYjKq7orbytGV6aqnHbymXzISBokCNmVRbCUz
cgfrb5IGBHuiJk4MQ458XQ7MJxE2GmYF0eZU0taDC3dTmX7R9Lcx2u9POlUNF2DN
d1UMHZO5aqRUg67Um3L+KBpvVKG3dDf5pgPcQfRriHKfdkSl0FhWju8ViwQJlegJ
jGL7o/+1Xifo1HJGNculRrTxDU7mj7hV9fM1awK25GBm8GjW8uFrbCc6g39Bcp5m
qgrgkS3GngVJ4AJX3UPY7QutjRhblDHrHEkarXRfjxwbPBlywOJow2gjd/HhqfKr
+0goqtYBP1LDb2OZ9GzryThS0+yPvpwqIOTlD4A4yCQHXiwTIZvA6eR78aJac7kW
Gc3AubYRmd5dwmxzkIcTq9b6YoSeOZzNBrmPxQLBFtRcJ4ksbILF06CHLw/1GU13
Y1Xj5I8gPtHAX/sgw7ml9S1mXFSBvnqcvXp31uD1med5X2qJf2USQcONI+CS7Pu8
br3c+lxYrQOTd8AxWOWJHd9S9hBCW+ZYeUDL/rqNJaFNscg0OJfwzuDIeSvQI/7E
onhCkp61FL79vvl7kZKbhJYbrDMj1LopAWrTjE0dZXzkFq7A/vSlyf3rO7kmc/UH
GPdXAVwpDqtCZhXgr9YgZ6ZKmi4re9EtyljIVcw3bt8N2gSTSU9LQ2RcL6CBDhdF
nM3G6EEwUSJN5QLNWiJwXCfVT6bkOL7Mv5GK2hbWmtrqgNWCz7od4/eEH+URYhdT
m0QB/+Bwn2aQUjjDhhOANO9p4uQogTNSCRas4YiF5ZmHh7F8J1VusSswcf4ejKJP
dsnXbzoK/5OWh3KW3WAuIiZjE8reLtsFkRo2QF+fxU8yyexXGkci3fPCAjOPeWeZ
PjUh2xUGRVYmByYNtnmwDxuAGj5pptUkzw1UEwCVUXBZXFhu8I4qiyWdSu0IPuop
KJK/ixvB70y+gzwXz4dvSlg51uwcDQCjBwYyxJHxPHuS+6qMc+yR0VtpmPO7wkwA
XzOB0gEvGoOxEJXGJo3hqMNekvi4vB/2E9pELaKomAmiNjb4tyQGeduwLchyViPe
v/7Qa+VOLCLPVe5oHCgGTOPI7cnxqrNYgZxQNuD/Ziww97j6Ex99M0R2kH100QB1
qJk1nLjr3V0YAluLcQlMh1I/Ghj2Msma4As4IpDDdoAgVO1YtvyXA9jPBd0XOU9a
V6G4WKdo0kX83RPE+VDgekDaNlJd2sD6xcsU/DUPmJha1Bbd44DvRXasWfS1INiv
eigaODs3C1SKLbKP/9qXIC/lz+4PVq8g1yQzmjeXdbZDjrFTp9KLQT7kD13F68M5
XFNl0ugO+PrwVEz5Nrois016Va1T5CN/2o+9Ft2ykjTN1UKobHGSf8muzNTadymA
XexieOZ4jjzUxMdsl/0/1GmAXp6fI4R7YucbAVViJkIwlRrCGfmLnAbZ50UCjhIO
1XRKVyjUFFSct9LelvwXo4s2c/IdeNBwl0vv0Qm9D1RKwlGq/0x/u+porOKiSXX/
14h80wOqitJ3wZ4NOOQqeoP0k+jGHV04aDd0K/B6Vtp1jQN3IC6crKAiagNvNQfV
ez2VSR6ps1NEKgdR/DR4z6sgDETmIX/+Vs9Vq/6IdsR/5iDqWC5hbgZStsvXwVTa
JUuK8Ieb1Cbu5u2XFt+6+jPJhkCAftgrTk9n3T4conXARuZvVDdXUTq6nOASReej
5PmJ4aQhDgpSHoJZn2bdVD3hCfBl4J8NjsTgb1xBZ39vH7NmsGjUu7tgklwMPKBl
jqKABcv6y/CUTUYHWgdE/eAv27rItjSnYCLw3sosytUMmB67+1tfuRBJPhpyRmF1
DTvPvCniHXDt9Vr8RcgCKUGF6vA1sD6FyBIW3sH8Ze/jY47HR2PLOljp2fYc/hUy
tL5UbfTtwWAKFA4PR7lDsm5q89+3bkFOWCXw8cTTU3t90pHwbLHE6bl2zNm0NPIY
GXNRkEFsaaU62XhnTey1Uisg2upq9xplgJViUoDvc4qwzuEY9HMQGXs98GIyR8Vk
QoYTTtcVMnM53EwQHsAaO7P/Ro5g2o2zlXwnaAl5EQvo9xucTLRmjZOMn/7MCETV
Ce1prG/9FSTZADRr0q7oS9/jvmAaVVm3NIde/Hrul9/BkXz68cUGYONdIUBefAK+
DXBCGYS48MVrQVoMECERbvQwCAy4rf9gOmLhbzkHnfok2OtaVzyrWG9oWgoyPQ7l
yomy65r9oTYBaUMmQ/hszIWeuA5dS8VffE3TgFPBIcTdfyOviE8Tm9lJ1llrL8px
8QuyrVyZQwRtmBg1nFi5oe0D6jbqQ8t2XG+gFJHHOLrpn7jbmS3FXdH/s1Gv1Wur
l9G2lF9BjTeWcSRO9O9u8imizCaf04NKPxYACLFT9WN+et38q45f/NRz7xEOc2y5
g3DEp+XBhPC/tHBfpvth+vbmp3BFzopm5eV8sTnzSPlBs1SAcKdCdITlBh6ccZrp
FCxoUWy12WeS+vKMuvbx74/7CzsUl+ITF48EyQaQoKO3xhO7AdHEXQkiN8OiIEy3
Gzn4IL2u2EhPoCPSrgqVHSzPVnFh9fsNKEsotkW+F2xWkGrag4qd4o4X6IYfSSZ3
Qy0B0lol/GzNW2WLHIVtYnFTghDz/CW/rSnN8h5z0ZBlR29/wHMF3Hn7xYpM0RAZ
owfKmSMgohyD1wXENyIvpp5OUm5Q8H63vLQ5TUc8CuOoFvh5XMWC39cuE0G4F1Pb
4OSCdVN6cF8gl8Zxxhzsbe1HOVWsdagFtE2b2/+d22vbEl1DcAGiW+UpVcb6fLhj
UQGv9KmcwmgXDHZra1p4zOCJPu8j0SG1ru/gjmyknEfRuWJvSgAAoUIrzNBc4fyl
7wInowLFlCZCEAmodFI8hkJPEK5LKEBUslONyJcQ1i2vOX6tYAfyyIxVNJ0WJgZ6
5dpo1nRz02u+KSwpHDNMTTSMhpBzPoucuvrEAUpUPHW7jZkn8h0heb116IR4xGJ6
w1gWGjuHk5Lh9kipt2OVeFXPYGWYMZO5VrCaW1ymsPdF8GRm2KjoNArct2vCY7pT
dQbg9DKlDYEBRvvHKS9idCLNvTmyw3ataV+LojROiFNCf+lJk4lC2ch0LebPGcBF
lfQhsfUkmZQ2ndziqXTU5b5OEM79OUMtZjYrQ5ecXSwNy8pTMhKWTA/Wgrf41+tV
0KVKalWwT6Akaz6rYv2qTwOkNVFygVC6XoN76vzlhiexhLxDUoxcAuJ18K5iZC8p
63r1HCy9judbzGJY93NTDf08iXCOiEHugEzaKXt+Z9JKL1+Iew/H6EgCA5IbeFaY
husCidweuKb/iIcCGAPzYFIqpoIUzYI5aDfSw0DEZVaTfVX6SROibklkuZF/3YeW
Lst9v3Ibsy5S2fj4NHmsUeo7mwWox2+z6qsu57Fvpe6dsfp/nyrHxHwYkaA1dAzV
drKeFNPiXJsgm1l9veUgDcE1Hlnryhg+cOXJ4kPHHXuUFcY3/bv+hqtQw8rCDJ0t
boTaQLH/mE27Yk0wPlmrhyMf3SPy3CQgcKEZN68WKrFw3o6U3c6MHVTNLAMrbZu0
ggnA6umDrB6AYCfZmcKq+eAsFZOiJZzAvZ/fUrLc0wGy9ohoJVJfYIuEagPO3ne1
DA9Ml9BGmQthr67xsxswI2+6o/khCklOi/PsbNF44a6V4FDJ8jcwUFYjDz1WWMO5
jzAu15CH1C0xd1yHCS0ldCChlYVsbyrxbqp/qKkmUY/R8g7xa1IM3NRdl32wMf8h
/sIlFkEuIwcd8aWy4DZ07bEOj1eItvypaRy4N7ZnpmrgWdunBztAe/jqwLygcN3W
vzbNh6gnCr6kRJ/h34ELjmRyRToiQVgnDvwFY/4sfc6PWofCHWf5/JNPX813giIE
Gettei0qyvPgK4gYyF2xa/FbJdxi2xVkwvDnf8ruCiEJ1NoCWLQ9PHCxishXEy91
sfS4038+aRwlm4mzCr+3BGDO4WSeSopUuNcaESYiM2W6zoEZhOH+EuZTI3YefbVs
Qm5jeItZmhYjcS8LyyYPJBCkqIKTycCWuvWsVMvNflm98eC0EtFBw41q7qBB9r/D
3pvTHRhR8o+OUyfrK3tkOd5GlSuqF68bkP0DlpEcowdCjx3PP64sPxMRg4LGs8oX
tqkAF2wEsO9dJG2+cznQoCXXDehPvW/lUskn43YsO3e+eBpkhov/pp1Z35B2n+T0
lH+dyWfv1Ra2Sq6y3AybW6k4uEk83VWWU27uiDCsgTzXrWwJU618Be/BYhdhz31W
6ZwXv25qDWFnQ0FCAuFddv9HwyFAIryhYNhWS1LPMMupS1S6n2ql+WzaWe9nt23U
WN9/tBnyAKfHYc7gnZuwIh1r7I62Ad3DLa98ALJdE78IfGMoXo6rE6OYwgQDgNBC
RHBrWeKtuVJpWoG113PzWlhsNYSCExH94HxrUK3CLOSJxZmiuYUS8+tIKcQV3mM7
nQkDj9e2IPSJ2hbwo6oVvTvgf+B5BJXRi+s5uEmSnGWLzvSiKFgNUaWuieZkt6gC
JGHtSFMpSwx2skd3yDmfKNDZObxAUs1O51zOuEcr3OaPn/aY57E0BCPD/Xwm21AP
8IkluF7cKJb5SDV7W7SpbLYiksJ2Cm/FMMvNyGK2cOYG0WbzAx/nVD5dTcZVAUu/
Hn5rRsiTFQ9n+OtMG8d4WML4s6EC4EIeoRH/dJMWbf4bhe+ggp+xwkE+BxsnV3Ah
U58Ex/yyP8IV+5gsg36e54iVZmeV8pNR0IDegbu2PLDfXAasATKBzbWCWSgt84Mc
VrD0Zmzr3xoydh8lKCIdIE0RlTwc4l8BIjiXyE2mnChrgKLu7+14pPzA86AifniS
QUw7I8Qu7u1eZj6xqDKnmtAwHrKMQiCTl3smDbVm+K5GsyyNBD+aBAh+lSeVvoaw
dFp2ajjpI3rufCICmU/qcXDiUig1TngiJA0qqzfI6RKUzqzw0RUVg3jL06HyTxuT
mmLOG42WP9WGf6x2Nb4uwT7eCpmsdUqPmsF1WyNNNpscDTHYQZ2813UEiGGckz/v
NuXIK2twJ8oHHap9/dNgBW7I6il3MDmWqEVxgUB0eiW2VspzukSluM/pY9d6gK/B
q72UOFF6LktXUng9ldfmnW+8jIT2L+6eU3aaG4iuaPCuivWd6pa9crFZGchA1Syd
zRz/JghzQE0vQdiTaX7XzLLiYuwrJ2hsnB9uunSu4bOlquwKvenxhpEs3Dr4LFBq
fKphMMqJYgLxnBwCksrR3DIXyPfjTg2xJfvwbLPHPNMNgyexCUa5+6v89pzvERZU
RXiY+pYSpe/uFe+Ql3n5CmHD7JjEnjlFRMD1bThbnVOC1lBz8mjlNMrRR9QHYFMp
KwBqt+9mOTCIX8sxpvzwAq7ZS9THenEQBoLX22HZOirmpioodcxG4zGsRxD36J2O
XSLN9/Dwqe4l3AelxP67XxJ6Wo53bS/GwieWV+q+uYwEc2mdH2e4KS+KTwIMkfbj
V13CZkZSwu85Yyf88Z8jmmErGiOuLDBnHEBfoiGr79vHiCzRp17Hjd77ob3AhGxg
9/dIMZh7A5B7kGy/cHUVVZ+ijr/Po/J5zLcdFW5NwKld1ZeRGnl0tvN7z8TASovU
2Yln+S1zQZEmqPA5koX0ELuJr9mQ4Au0z+PXkM60R1dhacchQHRaCidaV6wzSfwY
20IapRKZAgVy1mJl3+OCHxe+m1pfFPrn8krV0s2aKFDm/XR2yMMmhn5SV2lgbYT5
6qZIGRJw709krs8SUgy0CYQQqExlduyOfew/gnHTx5sqsxLyKn1+GZ/bX11M+ThY
qQ3pHdVbUd4UzfE+DVFcjkvuZxh1cM6sv+cMLL57UbwemLR/sUfiCV4W1LqKrFT9
y0SWn2puEj/hH1kbJco7Ar0s06f9VrH2seXB6UonF3N97Fb+Ueo7gCXVSUmSX/9E
jszcRp8T2+jbOogSEBrSLNzszduxRX14Vz2oPE+n0g9T60k8u67lhJdT8s9s7LuC
mfMgeKAx2HPWTXddx4lRFWA8ULGaM35cKeP5lcNe/w+Nwv8MXKARyqaPGEzBH7wf
oo0Ii8Mi/ElcYzkHq87k8KmN15IXmOilhrhtKPDi6vLB92h7Hpe0oV9T/BLAHrZI
p5OK2SVcHPQsRgC2v5GdxYYXGs4T4G6tni2CB/570IbRnActsyVyKxCiNunIn/zk
qkp6RkPaAK+t/SDOonQIw2p0XChzdaVoF5axVJ/UEuYXgM5DglxSqOA2Q4azQaP/
g7DU2ORWVzkL1y4eRYKmvnWCxMRsGek42g1a56Pz20Djn81ej65sE4z1av0zyiIU
Y5BHnj7X3v7lqdFGI1disKoCXYZFl4ILCGkr1tOMGhprLC/JTuVvlPf4duo2nG8M
GIKX5XZYEpehPfQ45llcjKKhTHddiDj5lb+/QTu6kjNAYerk0F1yNhDr0ol+nQI+
3xg8I1R+wKS0hZsZ88fS+gzsmravdFWn5LbksSXlDQWe2xO3Qwc+7QnzJui5JxR4
393BNKJu4GCo0RuNEIC7B676ayJ5RQ/aS8Y9UxWMo62RhaP+oB23rWVsPpPJHLoi
L/DfUtFV4doNIkgZJwaEM7BvjgTxy1liUzvW6iAZi2hV7feL0Ajmij7DxUUucDyJ
FlRLMj6ueOkxJwKGErc468udUmhRX57rdWU+n0CssbAXeWapsd4Xq35sNcEfG1nZ
OrzI2sBXKkdEZeRvXtF3YajiL3mQII7dY7sRc8O+XRuhKhqHzf6TFap3WPanZtXk
Dsz6HtmwS38EI5KyIp9mubswE7cAuH68zM9qVJZvttZnhTuyz4EqS6FfXNZlrGWV
/8zExF0HqN8TiLhqO3AM+1s4VpFrR+xWBKPNi8WYj+PmU0VE9k9jfJoC/kF89axe
sawVIQ86ThA9zRTA9+9lBMP8NuGkkFHFJTKD/vvnMbSZlXCnTQtvcd3pbPOJf0W+
5HICdlDQe8kMd9wnP65B2vWK22oueYQQm462WbgQj8axFr/KLopsfRAeXkCv2qzK
i/Mphgt/FGtCURnlRtxsCMER55vpuj0mOgp0jc7kVejjy7C430tfQGvF/xR/g6I/
uOdXQjsAPBvXAuWkJ5crKMz6fjJxrQnluByHJBI2tTHNJnQlF5VPKyn1Exc3/hMN
bSs99sn5nJDX5YEehUQ6mxGpnSMDnykFd9uaFpwk9ur+6K4DUnpkhr56CYGS2TBL
MOWDNAsJ5mlfR/8ydbLqGVtbo08SiiU5uAgHKN5MtumE8z1gfUVuit8Fzr0vpKjn
jbPbcHvJ3Qa0JJ5jVVRk2gEH/bGPplHmtad09dVofcXrElrrixUGEPtqoBMfzXKB
8xkbiiXXOPm1exZ+igoAEusoOntbd59STOAQRqEsM+sVzWKxq/QfxnzyGZU5k5KB
7erewv4xAkKfnE2KNcgQyBFTEI5Q3J/PNTW3vs2vY0HoOgyyrEvJ89jUugHY49Yw
kTBmMo57MPdapWOk0ftdiHl8yOT8veqMkVldT0WocDwOT1sM/i4umXCfQjPtw0mJ
u8qxmL/nwNAZe1MP5UrsYUEw3RF6otUnsxPNrm2EthpjyjhGr/c4hClHz4nBRU6F
Tp8I/VDovIhQk+2AWFPlQCGlul3gTAes0uXXHEV8uBGJhavL73r8GpaHO07TY69M
a0TzL+hPT1YFtHkSW8rmbJ8k3S33xu2dmj8T+Jz0Q0rNTjuTB2Ogx+C//4xRxEaD
O47xHWVujyc+unbdBLId3a5pZja/eyJOGlbWE4OUG38hR3x2ZW8IQKDNyDf6bcvC
wSU0AhypJyg5CW8zU1e4wvy91TNPQrKxVcj5gPhAYU7mv68N/8h4qc55YsoPZFUY
B//tdHdjdtqjhxYelsLiXNypDaxIlc+fugwq3/pNKfFCnq/MZUGkYpHj/uC3elUg
QddWGyQ103UgmomZdk+ZE5W9tjmYSoPuL5ey73LKf0L0XZLV6M6H+68Q+7GBrPCV
HZQeRV07hK5ul/uAXzhDx3gXU26S9gcGUbQBPLCP4eV1SaZ3UStKOmf7AKK04Ix1
QDJzyDzfzmuUrHRjbhZ2n9UbVaBBQhVbSE8ejy/5AODRRfVAlx5/Sj0qTY1QyDTl
HVkfqiNeIy1SWfjHn9AYF2GNCvS+BpzMtDKPzAFPUFsrVqxHadu6ZnjPM12/jeqh
xuB62+k7ju0LljagiIVeMLj5TG8BoMjwcuQJkqoS0/SoZPKNVW4tquAnLYYSVOGv
wv7HAb+3lqkSrjqKUEJh6u9W3EpcdsiU4aV5oLEAlMBm17bm9xI77VoTH2WOALzf
yCbgYbPHVaRejx2mh9d+KV2qGjw2GJizbS+1QgD9b+SB305yatF9ZHNfBkGJyAwf
se4akiImGai2UbW9+JOWNCmL9OmWeiPiijsiVle5809enfTfIwUw4RRTvPHCrQCs
EMYf93SkMYolLJ7WjSUnOCzuf65CJID7oqKRUzcg2KrEkIL55YH/lsShs68LDtim
qryVYPgfftde/8e2jwLfQZNMaVoWXHIWZhW+jYKxyOWcRyawBPDm3yX7YPL7NyV2
crhQxibBu6ppccMiObS/ZuiADwJnYfgcDK/GYuTAVA/bIlEPXcuelqjOWmyFZt5q
DniCUdR7lrslGW1sSGWin/OujaGmTsBQYQxwPNiNeNaNRArQq7u/Kty0NdxzST9e
Y0UHC/+1bm01g72p1x0VVJqu9AWS880+x2t3qGYLrBCNfcSNnKcZlUHFvIpsgka7
/W6s90eI+CqypbdBQlE71GE/wJI1hU54GzrCEa4881ATnuY6fPZZekTDrIGrMOA9
IzAWmX5FCqiQ27xZRBxubowsRK/H+eg3aL6lAMRZnIKR5akP8zf0d0bSPFvMTUNY
TN7UBip5pivXLwz1EjWxFAT/zJaI1bKGbFrR+i10BfGRpyDTtprQvenyQHpZevoQ
PG/wWjLTTgpZxdmsdbVgv4Ucp+HQd0oV9iDhrh64OjQMJ8dbQgE8VEtYO5eOmiur
kK0RL2qXEJD0njb7/ur+QnsXRFXPot5D9H/ftrHbHKtJ9Ubc8C4W1z6fH7TRSsrb
FiinhoZKuyif4HmG3/qsJ5cs7DcehmKC6RVKhPMyOSJIDNO7M9i2pdklAixzoJsj
Er/wpaETE7yI0yHo+JGOVeVKyasdp+Rh23ncQUg6GVe3QNGHMD8dcBsLIhTlccdT
MWKqaeMTSO87pturObMFt3/N1tkYZhGcqsU2MZt5YsKJrqZgH5uFbr1EUzPRkeal
R0tte2rzpllEUVf8VSpt2AgkXp/FWa6ENBpyycf607AB2G5IYU4ek4kh88UUlnfC
y/1tYRwjqVzX62gYdasJ/l4gMQBYpmfDns/hWMVJDCmiGNPXcHfFZpjFqwYewXPX
Io6ceAs+HlMyRhnuQ7SqricyeoE8Kdt++U2AO5kkj4kbbMaijBeDtaJI4Qe5wilg
udXnzlyJYYVt8SP6ZCQ19haRO/9pB5eRKCg0/mYNN3F7r2CqMRqxMFKY/SMhcjIL
25beLXEwkWqJ72+pcdxTeHsomgQ+04jXzK7QEkBRdU/FS9vu7yIate3bmOOYfdYK
JBTYVB0jHM8PGQn9Gv0PjhlGNwdmJWtGqC0QFD9gzvdknANV2wAdWroiRYkhdlQu
r7TaCU61VDsSkoHm5ffL5SsZlFNUEnwzanZmoMdeHmhCkEMCsKYJ6jtf+/lYmcYR
ZAGXG8oj6+R8uPFB/tmkHAuofV+VVUIk4aS+DQ3AswxyWhtSQ2PXf8RKtsmUJuKK
bq8ZIKZjItZ5Lg0i+aa0lj/vwVMjjmA06hfujJ06266/IU73HRBu4kdMvMsYM6UO
ySDc725BitoUtfjcZrg9IqGg8DYhauzL0pifFR74w6AjUxhxKyYRJgV5liX1nbEx
hO96efbJdaIgL0OiBAAcKmy/dN+0U/p9t66g5WCYuFNimfaElN6g1XcG7wy9+wcO
jPQfYuTJ07hEXz1RKTdvynSBxLRToNks7skYUamw49wYq52LEA69yoIz1P0La6VI
rB8h8gWi/WNcSxMjfBZa1bJQIzir6q2kB6J9bR7QegvT/AJtNtoMUkGr3M7GDY/a
P/Xu9wtiH9uTOWaiP6JNenKOC9Suq0KlkeY76vhzQb3/eakDTW/F82Mug/5sOmjh
MeiJ5E4BTJuP1p0pALYlRE394M7voAcmqW5T8mn+X+SKY03LiRsBBfNp/qYjwpbo
o8RUjD0ij4viwIfw9vlIcyn3l1DXAQuvixsbRy4MTt1oNSivVX3E/9DwJxSqiYiV
bhV7XuK6X8RbKniodh5wu9gIa9QvPJKU+FBTX7xrd64TSZjvCnqqFuU+Nv0463Uq
zK3qLePXU0CA5jTtr20AtoZHT27VWoqWc02D1bnAW3DSo1nf71Mr1Eaxpu112t6b
huHA2Vi5Ue5+r5n1z2ckjDPB9ZL/O/42Y/F9UGChPQX8xQFZnRC1E0QCZXZrb5et
2PsTeQrr87QpFlJwjXmMwy3mhlbLo9nWqeW2AU8TpF/3hnsEi1gClNoWlEa4242D
GifYzAtKMXaWcv4J/oyaWy2EDGqm1PKkHm2i3UHPaUWk4D5y4Qm2zdSyDUb8wt8/
4OE+r/wmxuK0v+QIs4AdZjNwwYuwRviUqNODOs9aAtZmNk7NUU2UY+RK7s8SaQVW
gqzH4TgbTOCJgMTPeHGiQ5mnQ/sBVfrQ1TituK036MmdMzs8BlI+R2v5ogvs/paN
hT9sLO9xLAsiQpgeaw6iUKDQw6utfef6JAja48eRetDjP2QyyJ5O3QckX3iwy53H
9gZomJj/3XnciUWqHynZw7A0r7sO3lgBZoYjBrOtYzOpPQphiL349mvQr9le1xNl
C2V/lzxXjRkfcg2Z2RvPvF4NjEKjIR7KmAuPQt6QUUaZyTaENIb4Iq3U9jL92TO0
0MMAIM3C0yFE0wF7ygWBoRA0X+ja3CpAKGHFSPbZ9Iq2uo8SlA+xw6DvL6nDbjC2
LBf5FCehWuKDXt+BicZropORgxLhUqAOGq6okChjEo3bQuSNnnwRELl7Hk6CWMbk
zf+MC1KrIgQAWf9lavXGh9bofy5mXHJaNGjNMDKkAcCif5dCPMe6lMHuIpiof9+N
QiVUeDoRdDGaXPyWPIPf4+ymKowo3yFifAgqKsQ6pvWZJsRScj0Bokcu/JwjVZ7D
VqJRYgquQF/1mZaN8MrX7IYsZxXnohxEwXyvGCERu5Z/m8aHbbqOKlPWmS659zcw
QxFjmgtbdaL41/zaTWf2GiT57+KaIVmCsBlLH3ajtObqEO9BrtEtCuzwOKQeB03O
76gR7qj1ewM5Yjt7mvmv/MxOvcsrgKi/DGmpyS8lOGpESiPowA2jODXL47c/Hp7q
YTdCEYoJB/wlDsYxpocTtGp3q/I54o/Shca90uRBhWBVlTaQQed/Gqp8eCHF1l6V
++mqiQbDCstbHvi/JcgvswlkmbvVSamJ06As7Z8oS7J8Jevw8QYoxft7bzKo3083
YFcnIUbpgQuaJBOkAgGg3PGyYqrmLsr0tvJk8xntPwCtrO5wgEg04kbkOPno0vJX
R1WduXImeBEn49s4yegRl60cKfvgf3T5NbeQHMr1U/upSvgneg9aLIoxTsDaIx22
ln+vbtjI8LNqUuv3vUpGNpbMJrDADXW3gv2zDRhxzVLkY5od3UVHnqoXh0OzbSZ1
yCqul4viLzSj+43CjfDbuklpiWDP6MLT0fWi1H/vpV1N9cfVn+RiWkh2xdK4jlfq
q1zhD0UhYmHffDmj/nuNp+YDnwmNVouCyZUWXcb7MwmaAAw+J+0gUOVRicsk2vBz
G+IiSTma7u+9frl68/Hxj2cbUzkIJJbdNTsT44tZ88KbQtcNZ0JsONRqUMIzKoAq
k3DccKEWnmxsDoG4MR42nHFbCP4ZMD0B4KWuhD39OUjqsSxFwYLviqCof2LiEL8Z
3s5O4+MOqVNZUqm2nSxA3tWvm5DmRn3XZ3whbbAlzSVp0ufZhOlHaOL+tMb7i3Xp
DHotULPxxDzQX8SHDCkxjG53zxJtcfaGgW702/13RafovVmBteD9AYhLiZiIoIG0
OE+zkfboreAj+vGkFVQbTJSdL2tUR5aBW04jj9vMcrA6/eASO6+kom5bPVHVbjq1
kZSJeKEHhV4mbxz8pDvslHsyck5c8Dqrfk0KLQRa4wPDBNa9dkT1mYDb7XDYpsKd
ekmklOcZe4MLznodzWSTxyquIpF2kc3yX9Mu77lllfXHSa3o5KE5YJzT2iPteJFI
Ho7A53lHchHPUvTJia906B8IXzK2Iz8hEKVZ891AbROsFDAGqZlUIwymY5DMnlIM
UzjFz4ht3JiSctWuGGZxo8rQ3im73X7f7q+ehkKO6lxZHNiw2Q9GUkIjyObfHUKB
C3PVCF2YWRrxpkUXFv7ZwWLRJDOz3CAOSMmyhQLAb+qyLof5Wjy1J5k5VM7klhoy
5k+OIXY8UxT+gS4XWsBZH0lgUeheZvCHkgGLzjsGqKJ/z+wzSfJMoFtufyvoow+O
zgKxO66rx6yOrRnjTpbYU0B3yzTbqSGqv3HIcbyqZmklPcUHs2g2hrLO7X2QJOFG
fKpSNto0nZQQ0XfgypSo3iyg9g71YbR4ZNaq7HPxy7ZTVP2Eas30g2byM5TmPz3g
z0f/89nPEyuzovP/0lS2YAy4R+pw0/jhvWpoZZzB19p2Dz9E1orilkX3Yv5Zlzva
2C0BkvRS5hN9istyIVdOd02mt9GG3TEmzIAW2VVUL0kMEO/d/Q3ucCeq1dU71bd2
5Nffg4G9txc4peRER+seVFY76lKbA69ruvUmIz9ienLclNG6mnlKM/UFuL+Ab1Vi
+GP3h0WcrfkkbPmmsAmqjQaNPohxPFpWsOc5KILbMT1Ik8mOOrOb1REjrhmK/SYr
fK2rWiLbZlOYepOvVbw+90pTjN2oV5mxHW11Kp38T6CrE7WSqXezoeQDcw+7m9Sd
K7wgqwd1alJEUKghmiPI+oabArA1y3YJsjQ/UPVCJUsBk9XeoMyIbdoUCQ7S8bs4
CF/5lY77Tbago/CSR18xjxh5ErJ2f/jYikwnmXuHjvB5mSsj2NO6AYAxztCIzSti
zQNflRqVsJoSPYA28kqerKtvVCIvHMonI0naO+DgVM4YiLKe7kUZESbjEPSIw+bg
ZivzhRGQhCqM0q6p336Pbyu8ggFDYPaiz2fxSlb/ilUJd4TtPKr6zGkjW/m6+ErF
GCjrt2iHneEZcgBGUJPHl0LdoOfUKC7qEqjriBTIfp1w8WVqSK622o5HEEQpKL9O
XO1A324eyGu5oQw6s4HBWESLgXMNy1S8Qex9ZZDOZzEixJZDStQLnwE6+ajtzG8Q
5SyvOlrfMPEQNrSta5PaW/mSdgW8pNWnYCiQ3Yv7xf1Kekfj74MywiQhAU9t97sQ
Zgec0KLQ8su5QKKNpVqPVeyiztJN6cYdUIMmjehaKMc5ba2XYNx0wsEc79fbUoxL
gG8gXKbvAoamiUpDjsouz7HnB02bt9gAWY5WU+iqzjYmWTx7P/Cu178PktHRzz0g
Sbo2rl+ZtNjXfZhZCPVsPj3UprKYLNk99GDHfkIFPftBu/+4eV42rYXOo8Sz1n6e
uYa7dEl7QmQ5wj+mjeu1hDxaXcuzNgRWuS3ypuRMnpfYifp6bovP7RIU/kn6uGZy
Mcg3mu7gCtFnmRG4+FjFS9iAWZGmfMZNj6racjQ1hGzlorIjeuvvIdw4vKbipWof
zhdLNZhC6xLBHeW/Wqi3t+mHt7R5QyzQuP7XxkT2O2BF5TF3lAom/+DzpXn4nkMy
7Jeq6J0LDnCZaxuwZpRe+07ZgYjNN/U7NPqribeVZeEKl5/BGU05xYfMeQ4UZIkD
QYDIOGuDtzc0Z4iCBzUFBOu4nnZ3zy9b5A/pjVPbF7YWl9B2EfVA/qofkLo794ml
p5dXtDR9W3pFZUaUxhy9weNxektNi1nulUyq0P1TaaFlFD0e8R90S+D399lmfin/
ltlVinO/RtwINldZg5+u2T7KrMNayfKAwdVnXTd2UDFKA6L2xqpknTzKln7oSkgl
3LR4MI4yj26HtVAwB1LwTv49gq85Qb8e8ITDXJYLdaKmcq6mw8u6f4pGQapuhR6e
`protect END_PROTECTED
