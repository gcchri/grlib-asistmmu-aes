`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fDfw++A5SNVEs5NtACWPlTRIRpDesxHrprmyNLyBQCvNigVNf5dGqHw8zPISntN+
m6S4R6KTA8G3RZ5OpktE/u//yM4FDEyAU4F4882w434/wTjES6ZWb+BbRilL2f8Q
IHWo45QZad9hEDT2FCv8ueV9Gsdi2yN2NZc1UQw1QgE36nKbb0c7wE8lCch/Hohp
9XcM3vqZoYLYzzbL08zeEF6nfE8C2fCD4sEsE/5sbgt9IwlsFhVxFJQZ05xdwNcD
7bZl7gO6cxiUZp4V1bfpMO641N88aMd75m8xghdyiG1dhc7jCDhQukoPjCvktsRD
2UXPPPAS7gWVBoiw5j5u3Te+pxT0+WiLp+1tGIKuR+sa/uQVnrVe3gPa3SEmMydr
WICx4fcftCX8W+NEC/8vNIxhBWjIEagawYe1YpaCH4AlzVijqqQFWsXXjAZe3+wb
hJzLaXNAkZJMk/IaJ4aOznd3Gg85DnRAb/Akzd4vAqzRQ8oo3CSixUpnl2LvKTQG
tazV1uhHnDKS/iUn6YPmOhneos892x/F4cBRLZlpHitcjVd4RqdayfIAbsBQO42P
arfgQeedME3jcqUezAuJt5IxMXs2WeLQeEb2A5xgbDEOo+siC1uNevow7I5/1G0M
XwU1OUDf8zA3vrOJH8hvuWX+vY4ysVqnClRVx9kmNyVnej1QZgHGXAJ6PxFE6vM3
x0XIkZmU0xOX2++Cvmfa5g==
`protect END_PROTECTED
