`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z0sa08VX4AzcwIrrzxTrwQy6SMxOEDYReUmXC2Pmfd4dergx2thMACKl4h/xeUkq
F1P0Euijs/FsQHr2zQ43kPkI4939BIg8j5JbJNSzQFXbvOKJACyYnaqqIgMvGgQJ
Dk/MJ8OFkG97m0T8ocwNJXCfoLXSWNyZvmN8JJShs5VKV+aE75KALkv87r6xw//S
AyEyx2nQysWjsHOZrbwZ8fz+UrhFT49w6SkHIcJYwp0brxBMW3jke6lErxEKED/e
j8XjccYNToif83b+1Vfz1h8TIUZM0Nq8mX7y1UwV6lbJdsszD/TuO+d5c5xT9o0T
2ycpkf5rUkDRZu5Ihs9eqGOqu8texpZLQBv13PJOGsXeTHj4Lx4guNKRDvmapc5M
`protect END_PROTECTED
