`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AbkEuQLSvuJD/5x2vmDVgmyCPuR31h00dOo8TVF0hrLBtCk8AIlFYfdu7568gJmz
xdOKuitFFF0/40Qnj4iwrWHHqpqbLHN4h0Ub3FRpvsC84ZQWzagxwTkjbW7qkS4a
Oxlc8Fii/DMA0s1nOINBQlUkAYrD0sfxRGyba/rqEVSZA6FQI16cHb+ChT/lCpMH
3Mqw9hyhPUx0awrsbdL5SZq1vGb6S+ni3s7JvOBv8fSyQKdHZdr++HE/c9Z/a93r
ivXSvpzK83OYuA/tnGebXO4pVkYfR2Bup87LceZpUREfCyisjHL96iACidm0pbg6
uxVl4TwIu8z0WlAa9hwf7+QZ9xawss5MY5BJa3sPXRQsWBaLm2wYwmqL0spry9vN
ZiGepzjsqoI7URsrdpS1MgR2pV0QXJkQgNNArlHbMySt6sFhS26Ig/Xo2u7VJU0Y
yZs/UbbAAKze3ctyYXKG+33t7E2nCOBFdJiA/+sSH646bsoy28jku9TTMNhots0R
e58Io0AGDmfJrY2rWzki0h6rXKHdRi4ozFsTbVSXw9XbgmVTGtAlw+UjmhN0kok8
7Q4GlnaXB+EKl5CJ2Pqss6HdJXdrH/nN4N8x1r8xxYbb0i8TZqpL0NIvrfsHcvVr
eQKBRIJjD2Sh6CGzNJ3T/5EF3OD5+dWJeCW6iaMtFYl7HBbIL78Ocn4yxvQo/xzg
7ZS2kk6tairq8aNgSeqCJ+nL1Ur7rgYpSzW96U5aPHjudZamfISZQxK/k27U6XwL
ARCPLQcVScQoXNZL8zVcltsRGGijBggHrNDit0k7fj10iiaqlvjrxW9Xaw3WpZSf
VLtzIFbSWTt4cd3PncbdcSzbQCpbwoGSQ0J8nry3empOQgfsCJXYvvwGTrPFVNlG
8hMSd++9Uy2sce65MjY9p1jWSoFhY7c5PerYsvyvtzISdoGfot15LJc1RiQ2vjDs
Qq9AouQ5HDAHqfdrEEAu1LHezrgelj0qkhHWUReg+z9Mh0Re4NW5ca3emb9QqjKI
uHz0HmDM/wjUJFe+YqSVniT1IiZhB3k7tlMH05pdySLLYlKaQPOdaVJSkYoZWzF2
1x3iGSbSVYSWYtk7kYU9B+8HbkV7mu3CttZmwA6a0KxV1U9QM6Pcf1V8MVcTtYPq
XIxYcvzj8ob8BRTNindP1PGQjpKw1UtTKz1QRI31b5tMEU6I5+X2Iy3klQ2GW6ID
RgyhYR51unu0SGvfadp2aYCbKqMZk2vZWccbFhbB4AlbYRZbJpW3pESB56jB16hS
ZQqAhG1Tn0Y9493xtJdeB/lAbzTGWMbpODnu7mkaAB/AyItR9BTIjFtHh8/mk8Gk
zApFOvaGRJi8KN1Oifdwnhg1MY2+8pBWjrRmbTcfuspu+QYH9cg3MSm/LBqq7EGG
`protect END_PROTECTED
