`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+GSI/IJSHOslSAdditzsiXUruI+ztSKPwU1+zWA9qTxlrhdaGfWNaaO5viGaiLuM
yD5qvHh3SoGaGVrBqYVZTKCaq/2ygTH51PRlgSk0ArvyO3Ys+eQsOJtGeazlXtDl
XU+wrHsDYjprFAY2Y/fQW7CPpBZZhLyE1YVuLa5GmdZsF2Ht15Pfrfn1hiSc3yOd
zQMcTYyIvHegoNnt1P5S8XVUOj9JShCy8Q4ohFTpq61/jJJslwHUV3loYHvhYpXs
1flCVme2aaOw3oSpPxKGWg==
`protect END_PROTECTED
