`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fTA3VeCOWu1+Bba0zU8uL9lJyWSEJhZJ9rrsay1L3iUk2Yoxtr/S4XQAJT50je/S
RCo09c/SV+F3r7Sr1CrlCvQ8PE1XZcUg0RSgcE9FyDyqENTHusjjIIsHGdqWaOsO
VsYu/paNiOds3LtFSlxJAAHPFLizfQl4GokgCTlG+MCIBVCsY210xJpqHdx7Q/Fh
0xrYTNojHhYLdTYOA6s7yF9/Hwgdb+DI27Y36nz9ZeamWteVv+fKclrFCm49CapX
p4QtUglMRxeHhdd6Ft7oGswnMCd9qN7Njv8b1UOnpFOxwrZ0B7LdbosvESMJ2OJl
ZSu1WyTwUQz+8m/SaH1iYB8HHxusQI5TBHHxn0C6ubcoZc6uv/HqKK3eiKP6nEmy
OQ4NZD9nGh4PB5W342k/Pqy68y1LR6uWcS55n7VwdvdXlK8zw4PBqS2g+6SCEHx8
LoCPPqdmKZPdl+VI7JUkN+dalQyZYCNPJf5UgB07RfyCaCQ3G2Q/fEbwkzsjP6Rb
ZrRgvU3zhL0vdPheJf7Q1rU1GQKtOU/HQzMlTp3x5W7s7dWSpCHftk/ajaA7Ekia
e57FYdH6UVEcqnI7rPEm6TUbBW0hzAcQlJvfKo4NrkRxfeNcFapsFwOdZaJUoNB4
FyXQK3tESHa3ketiwMh4SZEr4HdMZATqSy78vNCgmCdtzAOd/Nvlii9kATItexsP
RG3yu93bkB0PDjscV7lekYcXm5KVF/ijwpjHSD9EScSsto/tStpSbo2nxBhbqWyp
L2UBvicKiLEniyR5xHIysqkpkKXkk3/vVArxO+UbkJf+MJDcASl2nQakQIMp8tKL
nFNQWYdRmp9M7uvaHgOTtEmX5vyPib7tA3ol4CaB2REWSGwm4Vc6eMPHJfToCFFX
2asvhFAZGYjJwwj8LkmAxAGZI9C3y6VRwq0VHEhnXLXS7LoJQsmQnseR7CGXBkX1
U2yjoAKot04DVYHswG7nOoD2RCGHTdNhLkcm0DZJ4r9w9aMHAEVij7J/2o+4JwWP
J0n0QwQyCL5TARS2X8lIuLoMpC2rVpZouBcwjTJONqEMaO+MIfX3QtnetPqXyVD7
30U6UlA/GHuB+/W7LpCMvnJLaam69fqx4YqI4UlwXYYNbiiVY5PVmY4fkacJnY0X
DniSAzvL/I4DG1LMcGNISodDfvZFEoRk/2gj3GOOx4++i76FZmT+XO4A75YjUYJE
YpLeo1Elf7DuFwEbrnEF/t1B/rf57PNT2wbjNLLcHEWnlr3W5juDCkqNf3d42qzO
PEERCj/3BtQ7nrrRfI469DeB1ST8aBdvU8gE0urxH5SSE2OZqrzuYtNzleX/fVts
QI+tDwPSqmcIgsVlriQ1ApKFYrNiSilmsoOwTNMtjySkdXnxiK4509SeMO34NLGf
yMibHt1hRTonnsTGdFsAqXBsJF5AstZqneEMPkwVbAd+SVmYu3O7cT2FHXwqjTUf
AjcBWEc5NY659qrq5g5FDOuIQX8R3xmaijLC3NVBbJC7LMQGgNC9YDWLY/JbOd0I
H7VEGuG6U9mxteHtIZ2X/w==
`protect END_PROTECTED
