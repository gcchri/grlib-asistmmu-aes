`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WzN14zFC1ejvf3X3SCE0GORSNafQXIi3QusEoVgfIMz/6nIiNTM0d/jOobA63nYt
N4D0RQhuuGx5hQsKpNI6Z7Vae8XnEESwtKCn4Au+gN8JpmWeQiRVytfnNcKeDCjj
gmneqUxrfECsF/Vqx55Gbd14irIHj5sARa9H9MlpwlWfCKJgJmlhTBtfxnxE8kM/
dai2qFJfc05ZPijnc5W1Gj/5Ukedp4t/BhD1JxU58RJo4CNns39rooQVjn9jKKTI
rcmLjzJuwmVZphMD10NnjQfQRkge9/FKWluTilSDwgZT1pREQM1tSWQ84g2frbMZ
E8EhHtAPxz/ype1lhLyLPGIVY6Fw53wp37gTahVADxoiUbVGt2w1WoQDYjAS6ibg
Dw02VmDh2IBzJvQ5zXN0qZ7VxO8HhVCQK2NgLBIEBlHzsnT0YE6SPNq8JtuwMFY+
`protect END_PROTECTED
