`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3DCBfwnszG/SVwtRUl1oEAMd4bCC6bOqNqtALGdP0/GVIL/urF8eRrwyZTIqWWBt
yTm35CGI/2bc4nTd1etdeRSxDOXSldbaPHEnBKaNiEz5+j7g8lvnEywJRVk3S+aQ
QKSlaHjtQo0AvWJ8cG8sb6zaastF1cO0zyNeM4t6ch/eB2v2yODWb118ldaIbICk
f26o9aB6BUHG1pOkmpUJm6bf0Z/nHrRQELnsRubBK62QCiEhDH+EAPuIzdXFZE7i
sC25Fl4i/LRODNUE1sQhlMqLz4VznyLP5KM+lD0+hWfXVmv7sJ4sGYhKpylz5rTS
mlBlfP8FgcVhgFZUs+E2pS4SGj0NNnFtBagRbhbFWXNaLWgUA5V4GHJjiec17vNe
WwetWeIEnTemJQXTQgbU+SNB1527urBPUf1rrQsJ/mxyezW2tdmgs7Mh1AwsX6RB
Ka7/RVcCzhEku3X9STr1uhbedwk923ceZpIEx8wDBrBLg69NVNSURRhBxb1TeSIv
jIx+KvHXBBoNPsmyzXzgclKz2gs5iAPXKtzphktdoNR/q+eDSvOUUpdmU09Y4L8d
ZNceYOob56Kx0j7MsoPN9bouu9SqY37y5LTN1mPRyOyqvvkivBvjSIOMhR4zOzFq
siAm0T4F6VAuNicNClMGfl4Pfx/u6jKZWDUdSiNmeAnUwDTwb2d8aFSVaK0Un8de
ppKAiTVIj4uWRndzTL0Ty8PYieYhzT0p8bQGHQQsNFbT8nHXQnDVCOBgYGzYpPTJ
8Wym/I3LqSeKvUoVWiT9zFFSn3a4lyuC2mYNy6LighJPu7kMpLPCnkYxTJPNq3IH
A6I8Zz3HWc0702AxuEpakf2D3C2pLvOQPdn9yhg4y3vEa/jDh9EPgek0bx3m6hCp
`protect END_PROTECTED
