`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JlWTXbi57JsDb6oBlX3zNptl3KLz0R8JiNFrRirHmbry+rCKfEXtLZQViq3dAlbD
iLrhI7bs0hM0ijxGU4/dxomfJQK0P4tuiww5z6nMx+0vS8Ggyu/Xi2vN2++hq9e4
+gXyvjCduzhJ2/xCE9NagOAl6dUJDihe+PT4qy2TlsvbApmJUt3Kj/JL7Ock5SWQ
zquMIjPmdwAzWeg0481Q76OwsxVmooSX+0x7S0ZRhVaKyVNuVj4ulMTsXtR6ibk0
rc0RAfwM0gcKirpsIe0PtA==
`protect END_PROTECTED
