`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9n3/76j8g5TfLgDoxbJkjTmYvhlqiWMfvB3rYBY+DJiMdhsf0WtDwpB3L+K0X0Kz
oBGWqkBpo9UK/fGqMEaZoWZTJzKjGRcWEePV8g66Zt4P31Uq/kqj3zLCSU8Bzx8J
iwb/62f/Hc4NBzWKzVqIWHGvuo76lLSbR56OQyhxWGpT9m8YT5td3JEnVdxBkFG9
z+FY0KACEyk0rcdI3LaRRCZkHYEyherLMJuE72JdOE0CebZ+ZWvverok0oO3MS+s
uscceIR8kVWnsPsizZueLTEgnn1eK/eM8QQ75Y68FEkJMMkQBPn8faOpHxISvZpS
cS2ll9aGjapCdWvzuIsN3w==
`protect END_PROTECTED
