`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
POFXZ88mMRX93jBFXCklpLBOaBaF9opXHfeUfz2KxjH7ho+ZtrbzIK8YRyUGIWVY
1UOLLSjsSX89zb0o7MoJIFODUCVoTqGCY2hunCKSqYD0peuEJi9y6DR1bbM6zNSx
YLZw5LfaaNYl1ywVR7wtssnIJCpae2/WJnz8PHmHZuyzdly2LUAFbGjVukN5tWxk
J2J1NTGF1bZqDVllE/6e81nzicD8v0tODEsh9WwsflUQccmLIUxjRNMyI1a4Qaj6
psGixtW7Ll3ZsFz/Mo7kaRJ9SoL4ISEztUsxfJYx6IK4ExkFy4MWA6KE5wchdtjS
uSRIdvpuMcYvNosNFARj31g1fqP0Sxrdr8/QnB4EdP9I2uEhAre9UxvC+HWyeQU7
FEOjGppyHIrOZ/GuSLRWl4fkyC+fG8xw9A2+0j3ZFL2PdybxCd5OmAkuKi1jB0Z7
O6Q38UFXJRWmkYVoRV3E3Rw00f0ZFyaBH3GTm9jgQykJNU3dy1eHzgBJLAsirKFO
xzymOXJrV+8gEOFrOR60F6CAaAaJ6x80LQMBxCZLwbEgh3GMbZPETbVHMq4avpko
AxNXgQpKPVZPEtN7UCuzmpsBuALRsC6TtoA+gpg/1AIQmn1V6iLkTI/82TOeX48w
cGhoZogYNafu8zRYaM8tt0NDEuM9XlMLGDAu17fN9pWWpBvlunARqWK9a+uDIFlX
kWrNLqKEFrCneNf1x9HWmWeNf6umdzox1Xrq9+jLMIG8XkOOtTF1HDxo80oCayRj
cEunmT9+7wcYMlktF3jR81m1j3EsXsrgFFUTCCFX52DqLRKWnlpvDlpaPdFKIb2l
d2V0P+b/chZuO6BHkEHpZt4fy/0R7MlQSfqzHg6HIxL0nEaWE1VqSAmMy5JlNJRw
jdCxCkgtggwio3kKAHSkMJUEmjmGx9ZPoZuCEZSPomumVcP6xWw95v4mZXhQO38y
epTQ6yoNPyikzEWM7pzNdP9khpcHWNZ5idjD8y95jKxD98AdzI07dDrlviYNwHNt
3rfvz4skMpOyXkjyYDWgPhfh1iqwA3/jF1Xd2bMhVpd6JknTLQW6bNJN6LxcJh/4
ZyJ0fNJ9/B6YEOjZ9NYbl34qc3Vc/9QoOXUMR+U0n4FU5FAOnsVlSSrQlhGFhXk/
+05ReggWzxN/H/D/x9wm4sLRJpRW8zcHBDsjK5tfQug4XPDA9t8bjkwHvWmtlEDp
FWUPQsirX+aueaYVhuPI3icVB8nnhC5AjLrlibvVZ7ZeNr4S6WJYcyOsjatSSXu5
TlZJ/RPtPfaw+k3UhY7C1S+CWc1vQtauWwQ+yT33pPJb9TIS/cbFaemt0v+3bIZK
aOTymYkzrkIUB7WtOtVe4N6jtP4rheSsYS335cPrmruqGVObXfSao6OPfdBqIqus
kHS+8ieUayR7dWxF+FwAKa75HghzXdwHqvNBZRjWlEACr00CTDki5/lTaAexxVfb
IuGMWZBemylUg2CJS52wMjnvMQ56rp5dLXD/u7QZBcOpuq1hS9edmUPWDisI3aeM
AwHvCy483wF4tad5iztG1pS0waKDDBMMwQDduQ9D2CQGbyjAT9pKTgAI0tFhUb/+
e+FBw7eu2wsOIJAPILRc+crYrcuB1LjMW2U5Jd3xBAIdiZY2lnayXMxIvIg+6Xmi
dyo8FgAxtcP+/JM/vw/PYPZT7V6SO0szNazujQeuTdbdmMhFPg7oC6yVzMk7pZXU
falrQk13VEQqW5BIfhwr90jqtANwS5GkyreLcnboilI=
`protect END_PROTECTED
