`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KmpDX3O9tUwN76S4Lkn7guNC4jPSK9fmr098VxuONRJNbK8ztj3+OZCHe/hphGMM
nE+Xk2fYyiJuGopEFq32pWa4HowcmGIHUh4BRJStWS3Ri1hRoJrCdvJVMBTAAXbL
4Drx3Mvrm1OISbJ2wj6xTrRR6eijHLNUNjyhyAiUaqEImtmvte1jmH0u1tujdpHm
Xqn0Oul6450NPYnO+yGbaXemXMFTgpG2iFEFi+P1xR6sLVzSLKNvyha8axv2Rpx6
zIaO1Kz+V2bEqtowhrm5kzh8m3C9JCJSTXMKzXJgAREI5icuuQeXH+z+++c3tvBp
`protect END_PROTECTED
