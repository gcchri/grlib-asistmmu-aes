`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bvFj3z/fO1YHSqIMYqioSz9OoL7kCM5iR6MSLisEMIkIA3ger6C+pmMKVcSR65Jl
3roCVfagD9BcukxzDg3SogeXCCCtr3X4phaHo6qXDnF6RN9ty1F4QNGf8KgWIldb
7XMttwxWvtoJAGdooSrDLuoiMZFhG2+Tt0wALIwo54AkFKuXHrJiEUYXrGtV9w+J
AYcI2NeD3+SIsMu22yt4OdtJOrWCGwUdu1gwTC8EwpIy/p/fpBaRz1JzH/jHMt7f
W4/sTZUUUv4KraUH6BZEuMnXS4p0zC4Xq/AJpMzrhUZ0YYubBazujTZZ5InU2wMB
sTSxRiMndvumfWg16vpqrTz/PrgYPuE0DDDhYdkg4zFXUncrNpT9R+dwlouov12O
o+G+9GIQ4DZku+nWMmZF4q2qYuqfADmVLEju1FpKvXG6LfOdK85IPXMqu1XACWk4
ElRqkiMizGNMy/lm4QGKqyUgvp+7oeWw4HsyrGwbFhKrXCfbkFXkdnWEY6E4ghXT
IGxVEI9Hdjyyo4QHZJe+n531jSPi2dU5egccBkfnK61Nm1Sj/ch2DkZ8NeEwAm/Y
tUev16toSwgGz1mLa+jZNr4kRSmxYO9OEgkjfzyo0aAygZLkIPce4GmpGhRb6TwZ
An0LYU0/cGLA76RR4FBvKuFVmG0FQZeAtZhggHmxtnw=
`protect END_PROTECTED
