`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
siAdIqc51OH7kH4BVLzfEyyuJbw8w7kdis0fM0lWzkRShsf4UowJPYD2tajzqiVx
6c9ZerE+tjWLCE+B3Ym2QwhwUNuIPvAGHNQLWa30Rm1Ea3U8Y9A9336pMtOflfq/
afmax21pCGtdOfFpI0eS1ri/jleeL6B/ks/l4OsCJ0mcypR//EfPh6F2H1sg9ZS5
dTfO5XLYV3epar9GYPUKqOBhwEAM3bFJ/PB+abxorCqHOlb9672Ql3nq5sebkayO
SZbMPYIpV2/2sjv2fKokg/88shQGWs8vEoGQdOypSuBXNAVeBLx7IaDvp2at4KD3
ofvNDgEPBxvROuaifhs2l0GMaWPbp/RvWbHVjQL3deKjz4jTC0sERrJAEfN3WWdo
axJ9e3BWm6qezc6v82eQPQ==
`protect END_PROTECTED
