`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aNqbOrpyIvNQIqKrYl45f0APqxWai/QlOvbwO30iLFIrYUzoGPYyJqlotrk/UhM1
Pv3EpqFO1Er6QzXkB+NwQUFvxmr+mXzAWKczy42dqmTx+pmgkHUThZndqRHKopgf
LuExdUyBeoeOawP5XlGFNg==
`protect END_PROTECTED
