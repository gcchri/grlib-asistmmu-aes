`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+dMgC4CleR8WxjDbSDwIYpieqhx3IjyHrqvjgHG2SlFU/a7m6wS8F7mr5O3bigi2
bpY50vZKgx+4ILfr0tb6DBuK565I+uOJfKi40lzz+hMK8ASDtcd/jMTcZejVSxOg
VFlNm2pzZ20r1NYQ6VowonZSbJ4oa4kJFM1OdYkg7E8zRG0HN4cHKIaAaMFLELNU
RGU9TkZRHlETXTTDau+ZYh5XyVSJqOv9dyGpVjy1OOWD3wnUpE1FtpxPIEMSDLwm
OPQPCfGGwBEC/5zTv5cYGYXkkHXg/2cJfjvyRvzv8zjyiXTvTKg0y9q394zdfvft
I8NlXGneAAYaBa8/Z4BpKDzqxxyi46IX5Bk48Am7EjqfVTFXEnBfGSE5mzxtlDbX
`protect END_PROTECTED
