`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ka66KbTSF9Svbyo1NkjLu7ELF7ZofbAVHdwaii7keuVqul6gsRDpnBWH8d/d02/R
Dq4fiQIlKteYPPHj5nHbsQj3SkN1h7rdoUwonpwzUwNvMf7YsWhPqeLQmO2+mgh/
oNcQC9S4+aecnsUfiQsuaExmC9SIDPtkpkJMrYcpvlsVpXH8ORTtsO7sV1CwFb/e
milahAaFVFlG9OcDjDymC9sY7ves82SL81DNQVJcJp90ZRwswMwJRkDLWlRqcwYb
1/PpoveBQ8loPs1UCxrdAMe9uEaLkuIKYizcribIMsPepP7o1JhBPu0DHrDhq/3j
iQriRzVLV6fZOe6n9jgF5KCrIRaaGHReWTruVUuNrdyULk/2lnaVepb3eztB64Qi
FeTzyo879elDvRxbRe+2OGN2D/PNB5Cwxe6/vS9Hw/BWrUoNY1sFVr8PtGNM57hD
d8bHlCc6a61BAs3Y3AlFvxDg9Dl+DUSIV1TUJhk5gAMrVqlt3RhHQp7gTq59TUZ+
ww+4+j4Oq7EB6VLwzs+tow9mW/raCafeMlWZpSfXyqEdIZeJqiMniSJrElQrRBx5
SdjW/LP9vKs7YldAClTQlvhUoySSTnwDiu0nObPD3BsBDIBBsvDFjF1TgKFud9pc
xZiGAbp9nxic16L+VCOcoKOwhCqdCJkobPjzz2SvdGSli1Sya7muKxIwgYmQQv9Q
PVH7QII9oQG4i3PvSS/E9HC01RokX7PJc+RtggXmls9ZEl82QYaeLIrXT2PCpqrC
dxRfKT3ZTDNjrugzER4iYhlUmXoMCAHoy1DyP6Pz4qvii4D5LdX1xcLUDnrYr3rY
97yF7YCWbPBmGLKqxmcTrA7fu4P6cnf8l8hRW6ADVFa5x4cjRLchLw/zW1HPOk6H
fzjqTwe5WF1i2kHsRxFWmSyF8f3D7hN6fKNt94INk8gxg9HGr6iyfJlVWO/n/hjb
3gMjL9KNTj2+kLtI6xEgrFDthNL5BHxxvudBaJa/AMePfkOif9CVE6LUg/0PXvZJ
JRot8XJzb3IdqaJx6qR3tiKK6AEmIe10KwGlTQm9hUGd91zQhtdE42fdp9nXflii
Chkbj40fd4S9ylNLuPg7XQ==
`protect END_PROTECTED
