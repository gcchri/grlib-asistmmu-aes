`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zd0OykrNTY9A/33upDfrLkgMM8IQx+xQrNUpVUWWeDui0YB2hcJI14zly6uFZWRu
DqeOOZYjDF0+7huHytJ7MhEmhe1fpQMcQ8FP/jq9Ach7x4NX0ZcwKEx44SIUN0Bi
cj4koU7hcmREd8GIv65sHD0Naa2b5XQCiFN3WgwtbvLwki32ws7FrqKOf/Q6mWn3
+oUNMnznLgsVdeZVnWpnCx7s4z2Gh0Q5MCB/1yjKbbKkr4fiy8+5vYSmNrK8RTYi
B03hpS/OlMhgM/89Eta96Y4XBREhcNFl4ZcUlYb4v1o=
`protect END_PROTECTED
