`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0M+qevd3nHDHGyGmT0S53wMYg9n+6BALVSXbN017+UCnZ+/04v292KdYBwV+ns7e
y775j7HB3bifQpJ8qmUTm81kvX24PQuGGbJ9SDZDTGGJd41OnuRODi84aa+twsj9
cM1tvE2suMcJ85eKSAgrZ3rLvJPyVJLaWiXFMf1kRORzbjxPwtUuttusd3aBgVTu
VhkZ6C23OWmj1ZWFMl6gWAC66D+PBeh4Y7yj2m04gbyDF7UsirRevEZTmSYlM6+n
LqTmKrIDMLQJX9htS8SU8xm3kaJfmSnVZrTP0nqvmKRfiAhmtf84NKvZpCIIumMg
sTRUAGKKh/N90qYfogjeB/fN2tNhsJNzjH0SGBddSRA20WcKNUPQSKo64q48uXxu
ciDV1N5I3lv/jUmZY34UphPz5HBptjXG8CQHuiXBOlKweIhlwv3RtIq2Q4LyRm29
8LV3Su4od24bEdpUn+Qoi0Iwn4/Cy4r+0NGSbky2RSV8BuXMEA+JcSAUW0C+GvFe
5wCpNl1G0mM4kgHw2fPu+QnvWshR6rJP91PkuzfTV9EC66X1j8534jlVe9KMYz9B
1WHEUitqAVsmJ0P4jypWOzR8mC5VD5/fLwno5lOAA+LCHgPUvwNTVrnIKMnuI/tK
lEHOmp3i/sdlVbF+87ncaQ==
`protect END_PROTECTED
