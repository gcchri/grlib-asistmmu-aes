`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SXKW1r3kbxH3Cx9K0nKaJB/BvHF82F1EtmSQTnae7YiRL8J2PAmP0s70u528f+lZ
skc4ehexOmS1/pQQKr4rZMib32hvNwH9PmvcVXuOXezh3MxPv3i2uxlykt73h3dN
oL/3Ducgfw3Y8HKWOOkjaadYoZP8Aq/FVcm7xDvwutyOlamP2L5DdUc1rPuflWjp
68gthrvHVtA6TxZJOO7KxwaEYsEZg4WjdWpspJS2fII3aS8IdBVgG4B+vmdUuPxM
LVDMuSR5vdcZEMdH1WTrfkBLcYWj9/8uILWD7pjQ9xE7dfa1d2DEPcZLJpbYBc41
rI7LgS/+e/I0JL+CdeQKosHG5mc5yoEkxgwtH71pWDvYehvshvY8PYrE7zshOR+h
EFCe4XiNW3hfxaptP3a6n44jWxUr66CeiOc21CTCLUw=
`protect END_PROTECTED
