`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bMqhJNC0ihQoBsG4L0Fbc442IYBHnYPUXftypEwJ/xvp/L/MfTyO3+MycuG1Nd4M
VlJPRmgWzBRU+kcDDh6XQM8Tlg5x/OOhF54beSnaDUyxvSp3SVBitgE80aRg+emu
3NZ5+YtRtyF91i2z0np/V4HpHUy9x6k2Hdb5T8EdJMynt82vktNpzz224MNyNv5s
jR1fXmI2VRRZdo0s1fHxCWS6rG09I0r5QKdWmkWhmGKIeb1RJUIBgJJ20luHiKqA
wkAC8TLDFZXHabOjcO1tTwXU7S015UwOlRok5bIWwyAvv6DJxJLcBq/ROls0csuw
Hcuuazl1XX11O2UdIpVw1aJcdHiH0BGn5c/u4QRjPboLLNOz6NjmY9DIQxsiU70m
ru412NWOoLdrX/kiRdGoQMWvkuJn4eukp40aqAfn66KVSea7p67Kz81rZAE7Ry0S
HuNEDiFnMfxOElJI3jzehb5NUXmqsPFb/4BN7KqVtwyHQl56uSpcoFiYXZyxftBK
`protect END_PROTECTED
