`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tQUIhyDDC+NjllllWT6oStlvD5wo61JVOVVNOjVtbN9MMf3BLob9A7rWpKjWChjF
h7ww2J/J7O22g9ZllV9+GLKC2ygqUCRGQxAI/XzlSLwMVf9lobrYzn7sPm/bLQhV
pAoCRWe/ZAfbiVHyEjqgLQqA8aqy72IFDECbIT/TupCDWllr2MT8wvx7VKAyDepF
0RoyayjGAP+6EAeVAJjwCiiPKaHP0XgOizdXa8iEWciOFlKofbyGM1Eytp532gBv
BB8PlzlMnwGFtJI2p0zW1lwXMZP7CuPBeXMz/JexjpNQWWlq6Eu2mg/LFazHQPO+
yaSTGbgPTe7mDwH9FsDh1YaNnFXoCZO5Ma7dnsYOtu8QToikqDwIEuTAqFC2voZ/
bDuKAYQNRfgyMIZPggbrabW09mpYIXUZRPdVLI9pIDyoo2c1HmT3WpqZvDFLa5K5
JvcI0SCAIyByyybo7cpg0LRR1BuXQWsq0Rt0ffeLm5UrPwb1VOkzHzDBNYrd0lCx
Fk1A3MGuC9+6sDTtztcoNQ487NxGLi3W5maUinHyyaHWnzVMu7spTf2cWr8UryqJ
zNk/rDceAa6Ph8LoFE7xW6R7XXc4tYewJny0u15/BVGbgIykU4lKkXMu21eAYi+A
PTek2dYLx/anDexOzxe4kzQ9zSaQDom6m+FbO52VKUoEAzfpU4dg6QW3FHIPnRE8
SiF7Y0LWQ9XUbDn7k8n+YKMUK7GslaRrU6xRI9FaaOVZG4DifA9ESw8SPxt7pNBr
Vt1y7LgGsDF4piyqFLK08R6kPBxs0O3e0FWsk+ndP2jhYNYV/lMjsVhoRzOZKsl5
W9Tc1koMjFcrWmGgwYQHH8IJOWMbqiCbosXLZLWad6T/QjyxIGlPBo9QL6xGZqsA
ao/kiOlgg01DJ1Up/stxnB3iYm7ulEYy02H2/SJL3CBrc4xK3/vLZ7C/elsdG/la
MbA1noI7Msfj0405jeKPUf7oG1LmUmmec5jIDnpA2Ihhcz0k7UREpeo2LjAfHbGD
6JDzffRFdfi7cGQGxhG4HzgdKCxKl/kOci6fACNR+6jEf6qD63WcW5fQrUpA/57u
aTBhWJcNMi4LPU52u6+i+I8WVfL+OzfjZf6/CGPR8jCZKwauo0deYhTw4+pjPGZm
IFYZ6e7+q9u8PlFhX30upcBsB0ePiqfQIX0GY6UCYQKsayHpto+XAGbi7u6FVdhU
A5g+Nv26VYICMQJYibHRa3ExS/BA7FgwO5Z43so6jEhT7BI+Rgy5VmxobcBRWi79
emq+25/v+6lw9rq5c50i3e5rASE8NFC5eY6Cj1eEumndcNYXcvpkYJN9eOeEk+hv
RHiwdUyC01U4idIzAlPtwaNWtvQKhu/2ugYTsIPpB7xwUf5t/VhDhyBNFESOSd2Z
waoA5oEk8A7fRejqrEl3QxpYNaD1ETiJyQtudbCJQCYqrl3ebB0gp9E3RPF3S+mp
NHb1GI632ovKR/uhKNZNiiIt7MOgHt364mr+boxhWjdEMc9/v8hitT6T3S+Nr+q8
pLjL1U/+IwZ/tnrNHOlCXYsRJ1+8Mun+6ZkSflFFXvG7/x3sMokyKj9pNnsH8+EZ
sNIQ8EQ3X7Dmz1w5kMXBlVMNAvKGqOvb2nV3rzEYIjbq6pl6sQV/ajM+GcUEizd/
XKD5ntxMiGOq6F8YPtkGDXgaFRcTHRM/xCQ1/EUCFVpIWl3jXFvZlK1XC8DTw1LL
TSnTNgy4T5Ls8ldtw7dXCyyDk1tah0Bw1ttl4SEtI7oUA+FaOVmHzHHR5flP3N30
Zo2KnYUAvL4fQUN+OYRQdYqfvWXz8x5NRbA0gA8XtznaNnrECwMCjyT9B5/tlYCr
LwAh3ezYrgM2oHMN5MDKv7UuSoXjIkhNnXi7KGrTrzZGz1dnbEyg2wKm6SR3A12d
40X9OoM8xobti1FGZgUhhTCQ7Z5bd4jqETkJg6HbSpdSX9P5imHq6Eq8n65TuY22
iGp1oF/shcfD6CBWQxV+LhDWsqaNnmp4NRj+Bn994JlRAuJcsf8Xmh/Gmr6SOUqj
kubhBurwztCqYd3+1QpNqT7LmSwGwyoJBVYscLSjokLa/wsW+nNNYS+YZFpu/t70
GK003h0UuE+4yHH8Q70bxb1C+CTZ1rSHWj0Pn1Xj9rB6Kd6pw1w1fI/oCEY7bAwZ
9XPpUvoeu9fJ3LJq5petLGAHS9Yd0NmQK5OIGh58gRkvHqTBY++9i6U/7Tcg9gBk
D3xAtTpPZi/c0AV/d613R3+Vwtgw4DuL4/i8CHcAaneOvAFAmbaiQestHvQ52RUZ
PjexuCOXGLWQgKHe+XqDbRn7TwgSc4J0TqO5K/F0GTxLDcHYvVq9k2VQVlyOuxqZ
jh+S+BgjhR5lFBcpiowgNxaHcx9qlO9OQIcQWVu6+5qXRp43C+u5VeFPj6PFYXZ6
ipwK9VaNh6bD4epl/saaRO87d142UzDUxhjrrWbAjEJWe2PrryaMk2iPiJetr5Mq
VBchPqC2SYlgafX05xSU1xYvvQf9iZt3oR0HMoIRE+UYqonEpdJjoUSHMGkgydbh
5KNrjyPgNBxk23bT+tWcbt1MFfV7zgYgsbKLctq3s0kQ1o0HOoBG7LuCGcIxELCI
mZ6oxOKj8jSxJTkA/tyo4Ej5fhBHDJBHm0gw2tgHS7vhM2N3M3Twj3JifXP0UWL4
ELfFDVcZvLuSzA+N16E5r+ii3+mf/3kdeZuuhmNFI9iJ4y+dLrWMDY9zCdfOjAzk
FH3ew21l7e04DueSMdexn3q1abmWWDd2tqM0rVNh3tTx8KhzNxjn+dx00XrhbTxO
i3JYAUfM5raMFSCzDbMWNVxAyQfofy0zl6Qce+XkZJJBAFuhzZqAroW9OsEEWnnp
jOR+k1Ik7jnpcAGyO8Mq17TkTMJcwAVAgkbu8gHVU2ONqxerkwtNkNSFZ7Bx5dPZ
/rLmRAPRaE0fWGKJZaVGk6Rvhjq/0tk2qdYvytklzl3suSnERz0qytqbc92YrmZC
hX6SDaFERG+k+DC01ORXvLd7FohLTc9r1OKmYujVjFW/qBrZd5ElM52SOvjTaxkK
KV+bBfQEhLxLWgeGJcMNR9EWol9tyc6KSgVzwU+XJegrgOgaBLdOdvC/JKLihAa3
JyH7b2AK28B7R1+pJu96oMPtqHOJAxk6y/lV7FYLbDJdfBCsN1pzAVnW9gTfMB4A
flP5leCY6fsFnFQx8itXEPIzSuLcUe+0V0I4l6uxes/E+6j2ft/jOiAGinMUx20A
v4xVY5b5ROt/pxmCsQbw6zTHvFw9yqW8OwZtYY3P/ZnlX/yWqXmsUOje1A+WM4ro
SZyxEIOrJrl0iCq4Maw71fLACo0CnPnLSBgMyNdXDFxwqf4kjOkbLYc5czPMK5nW
3uB7mE/Q6Hr2DSbVZJ0Cjw99E7fQ6WIEeQuoZseKHUconuLOwu0UpZ7TAOknf+ok
iLTz6KcwETAHvZNIX/jwZ6tbgcOLJmGj5L3aqWbX7DLHGkbpVv0Hufwsn5MKQSZ5
DQPOe4MuwsKTKl6jfSdehcyivBF0XWKVoR9Wv+DzIcog7izCm847iqxnNcH0LOf1
9dlbL8E63i+3LNTbvNqzqWMdjBE0id86pDvrpPuDlBHOtcv96X8yWF+LEg1O51Dp
i11Chq8+UaJModndKmQd2aHwsCHBPvqOlkZLp8MzAYaxkOaBKe+wTffryFOPCjY3
mnmNb9OBEDPIE/v5mEBq1J8ut3hY+g4zRZF6ymeb1FDPJXnZprWjGk/4dycGsKvG
hvRtCyFQwLTE+BAcbKIEqLAh2OHCD6kPk8lvlBZpn8sN9Kz/eZU0HcNvtX+nWpBp
NprZp/0SjsfKfs3HJi33BaZZ4vHrwT10bP2i8skYp9sG4UAVRFgQSO78IZ9XQeZR
LuDHhSFajMpMX5u2a/n3Y4NuQ5DlI0ZRlrbIwaSMnBnqjlK1XmG6ffp8LV8V/tN9
VnaprDH0X496ykFZIaHsRP6LZbRD37fV5++Z0Cl9U7Gw8tgkFkCK644X2JJH0w10
eswPrZddHMLuhEmU9Npkd3S6BG1fNMDmMiYcYFNQHhwmSZb7Xf/L52RDoHx/YA/M
s+XyplU81kOUBXlkpuvnQ6fuXxeSFGua3oWIdqHko9mEHzShl7QToU/Edt+PAh8j
czazz7RPDFBtmzYMS1TnKuTXAeCtOD4NN8dlGFIRaqhDZ6mC/jT1TdN0ftVmG2Oh
NHrV2UW0moCb2yKNV6lOV/YIoD4f3hCG1z9j0fhKQPkF8RzSRbMM88WcSq14SxvG
hB8KpBOsIvfwpHWH0cBst8ryuC4TeIiPcpd6MBGUmFw3QugTdsLKpmi1pNDxjOV/
NTJuDTa1E5RF5rK+pLYcvYoW+ES2MnD+7d1vitYxpx4gyTypzVT8uvRlXBH5ClZw
uJJURNNvTsgY3eSi9TEx43dN/LgEdc2Znv4fNrID4rmhbP+K6DUjFfZ+3YyQgFOS
PqpaJ12NRWjooQCkEeGmfW8WtaHOFP69KBm2iVB4pxzvzKyHb3D+CxiNnrYItecK
9IVPi4UNh7M9A7a7u/XJuZKqCpA7g+PDeSnaLQUPAeinqzg82uZF8XamybkMfFRn
qSymsM2Whwj5uN80KgW0JgKN17k5m/G49B1wRDemfw8JsOlWXdjEbePqk0aElGUP
I8b7mZeLRwkU2osaDagSqejgGrHujHR29FPNquzU0Dm1Lcz565hQ9uqZjIzN2P0Q
tLsci0ww1BWmi3gPBlB9yjgIwPD/0uhMuwwMw5fLABgXEwWt0VOUEr0V1ZX9J7Pc
3UsOBvgFwAjqqh4QQzV0v1hmMlmxaVjTJXNrpZRS7QNUg6dA2/eynYSJYqZZ8i83
x+PSEoPuI8UDfM6QQ4kt7sMn1wVFL3Iekgki0l5VbvwAnTVZjgYCAxSpFlsG3vfx
X8fTTOVS/42q0DD/Hbtn3WrzTmp3FH8xg4ZsSjl19Nd4CWyB5WDg+okbn0dXPY1M
t4JMK+PwyzTbhHF8b0PoqNcPm8Vt3z3hyaOijfvlWjaAAPwrzlhWD1yZyom5lAO0
yp8fgGN3c+proM8f4wZdP6ki0z7YDnU6+n/U5UO4o4n4FPnuHpGFuJlsSDtMSZM/
P/lq9pWt1PBg2ZWzCbbWU42S8V4pcoN2oysS8QkPs+e3+ekwSoTCz6HdulCLEzUo
74c9mPvGtgIAx7UQeMVvqZuj2tYapGvDO+6vCFht/EZ3ozDhvqXbhlCxXFnfxmCV
lpkJjOktyIlFMv0Mfiv8Z69TKo1OoC+WWIwFuVgCSMjra4jKabNX7ReOrAeWbFD2
CainDf5jFr/xOhAQ2USEPt+oh0A/euEr1Upx9xg+0BFiZMr0mxxUxnnP+0iqICsA
z5z5SR4+pGmdjDFBf85hTHWziYyo8LYmBE3x1L0EZxk0wl12jopFVfPoW6DtO2kM
wUnS5HEIZoyTHZpjZtwahU0NzC4EjX+jys4RrxMADAw3IZM0OwTXu0zcx1eOn9Wn
UXPdq2cQCt1dU4jjaSMMuNII8wsxD7V0icoNjBklvwgMDe7I0X+8q1xn+g2QqSMb
ycXaBjbTnU8w4DXK5DVUZQOGzHQ9oQQzIclGLxfuZGxumZs4xEOien+GUqBPg4Dq
5rK3PeZhoc6fpggEHS3GVO7eY5+SHzwcwZRUp9oEbMAB0RoA/QC7GYSNoNLJQVvu
E5doyYVk7QI4wwW/k6uAbILHcof1iv3QxxBkz1IkbLv1KomtIXUveOGQXmwIh8dn
Y9ZoCbNlr4sG1nTpfLvPOmMLQZ589Dxg/cTAR+sbwchGVOp7zXgQjhpmzxcJaQN2
2bDbyrasNHXynxzFLltZOGG5Kjn5ftUOtj7tu0tu3SzrsDGzgwpD+mqovbiq//ES
XvwWwEm4eKbDLCbFcULPCU+4Ts0YbqxYr9bCPHs/sVzTC4yxXhVrfvPPO5I/TbYz
2NgoBDhZiMOS1n8F9lb9mAlBgRJ2f+Ex5Ji3bfmItH1G0OZ9wolClKEvA9rUmiEG
RegefY6SwvlrJbrm8Hwr/Mpdf+eanxb547jfKiJJWcAY1VbisBGviUN9UOwQU2lc
xIfYLZUXycOcbIjKYz17ller6XKbG+vRq51cqufazzUUADgn38n3XH7pTgHoYi+S
wHdC+RfYvl9AG8dLzYEr0yZeieoNkApuymoSfYzi98U7mYeJPisbuaxQH9UU55kl
koSGHVLMLlZtFvhrf8LieGsIlnJJCgbao3u3icu5xN5ZmyDWpX1sCrIUYRYEcwmM
i4S5BByJja623mztfPOp+r/ciIz+PjHlr/fP9Lejt+WnYUZ8LLQ1LumgBeVtVwPQ
fD9r7xthJQRn2MxRZA/O+QgF/Cv23e9oXTrMy2A7pcVjyOwpwmLhx0iQIJxmzZQr
wVce8dg/SZNujSQfgRbPfddCS2OkRkMtti9xndNNKlb8RGp+sP0IOujgJkm3GkDZ
DE6YKmMvVvRZTCm8zuo7Kq7+XsmqzDSTQW0Sy7nQDdG2DBwid5RaHAaTlkic42y/
jt3Y7Vvm0O0M2ZyyY6zVeQFFhC042KMPJBgJLVKUCsuy5TKbEikh5j4VCRq0cTBe
hc93jdMsftzwYvh3RfAJkpF6sjH/IGYewQDVHYx0HOZkGTzbJ/ekXzdF6G7i3uTz
P+iJT0nZRgBEbX0mJnKLKUoehZLHxiRC9VNjqIqeY/OgaFPi9W1E6L8qcOw3t74X
FhiAJldK9Ke5Y2xMOxA270REzJLi32+grdP9x9I/GjP3bHqqTK2hqdXKVKIOlEWO
vIZSZQQGlT14uvxuPEmWzpGJ3BvADoVymMWuO7K4k4+6YRy1Oios201TTaVfXyd5
JGlDzU2FdRWkUKx67R9ARAiFcRUvme31LWIlPblij5agN3E/XVh4abzBm+QU+i4e
UiVQFsyTfzNlp/cF9Meiz1SarkznhOOwUGUUSZebQkgd86lEC+GyE2E84EefZPzU
9QM2NlH3ywF+IFDWF9cpVrUU5FeIKXSD3ybmQLRKy2svV4h47uwuZal8pTaQA7lV
4Dhhk4XjyNYluis85BuqPl91mHUDixj6RnoJIH2TZFryAQZ8i46BQa0HnW6WPvLw
ws+vzUxkbcLeSl360eJ88LSNFiS9CkDvNqc04veg93rYLpk2/LhutlHjLIDo/M6/
82dEZ764X9npFyo2Cz2moQH2rpU7ME2mSUxV+dwzJ8MEEpR7qg0sKakMbiVjY1d2
fjxhLzqwzdF66zEGKlic6815r1kow/1dSB5QrunX7QQ1UXBKI31dh7hKcZv/R8H/
gvnFvQyE28jEM4ApSLZdDEECTBKiPj2fL9Jmp1HjgZh9QuTLcDVDtR3qDybliFCS
SZCThP32uNSDESY8OaECMQhJEtGkmBYfykzv9nohTI8fVNPuF/w4bHDupUSwuqw5
8nhfkf9qRAYksyAcFlIgQCWzWnyXeHeiNO8ztobGYT2K17w9Vyp5+mvfqP93obXO
1wB9nbyqRBw7kAMZYt7bSox86joEF0AMM49F6Jh/DLTaWuGNjL8YsoKxr7YUpDCS
9OgDMmzz7+gp/GHrjaUnZu6gZc0BHhw60D1fLn+mwYNE/DdslOmU+ghDq/HIWE7X
jV8U9EXlRz6azrpnrjqlT4Igc5/6BNfkjsQQSM/Kb0y8mzDT4WhmVxLW9UJuKVIM
2vSSUwQWyEk0DoEsdLq8AI45I5dlJ/ZZdMrn1ZdYzfcVVennlOFcgwjevpoivXzN
YxDTGS9EwMNDNvHZG45MT9gcSsZJ7XvTOBP6LgDYZiqx7SU2TSWMddQDrEGbc2qP
gqrJGagoyYpOFkkIzxCotnYGwuYeB/tK1B1FExX0t/zJ6QPcmT+FeFmQ9yrwUtuu
RpRc01praanT62eQCeQrSYLwbz/9jUtqlhnfaBMv56mHF3Oi/o3wWVLDnE3pFP9n
n2+iKqtY1pgpqpY12F27sM4ydDk8RrWkWCg9Uz8DQV6QxrSP+LiTNmt0XV3pPKNB
p34N6YhdITlmEzshwNkHNJJAR4zW/Co0LuGavhuennIlOWcPEWICY/+yQlnwajlm
F/yKtsFN5FS6b+go7GOc416GAryfcJ5rjItB3O/t3QxqxzsN5nM/ZZ7jA/AXW16R
oY70TVtdIUGWZIyq/O4XhCmVP6t4Bvks9WO1VI9kO9lKbqmEdcIHBla7mbrQXIs0
H0onZeeP+rfR7u+jHy2jbH2mYeEI2qy+v6sV5risBHQHtPsXbkVdTSEbj1fI6TJh
KDV+fRr1GoqEsU//JS67AFDGLfe014XwXdN1TJealTrTHEEkUyj9df3kA/TOa2nQ
P62nrTeRbpTXPkSPsQ8LvsNIjq2VTuS0unp7v10B9k1vWJfZKUjIIXZ9GbUwveMW
kiyX3VaLndG6rTGE+m8CDg230ivZ1FTL5R6ju12ptLDXlBHgiCrBJKl3Yb7cI90j
8hWK0e3eTH9wrQ07PxaddXEqknkNmJ9nPNNlfCJMJc5zqiEcWLee61f8a8Nx/HfR
Cr7SMPtPLmwJedF7ERgTOojdOIKoCRpAjNJFm/St3xGF5JrjlBVlFhESnCrn6Ce4
Inr1MVhhjuChofich6BxXh819UcLNLkK4GrbD3D0g588Sb66YGweNYsOdmQ9EV1S
s5hTRcNghIS9uY7ulWG/F3zc/Dt1w1z9+IFt9L38gQyLrD4p9yA/mz2BovjtdeaG
UcSC5YACv1YXsPpBT+TwEINzlP0Uf8MyRcYyc0OisvkvjLJVuPmwtrUkBBIYh8j8
6pMUNhTkp5ezoigsettdzqHLTjkYJ/EwBSwRB2D7++rmDRLM7R/dzY4xWL2Xz999
FalmYc6ionu+EWt8opg/oY1aoyN3zJ56O76a89xlwTvA4qSceB21rf9puwcBV4jz
uWCxYPHXwdvS8vVnqT5KjqU3N2Zs/5cItgk+5KJ/VDncBmxbrxKH6D1wPYuAbQOU
hDbMXPXcO+SBWE+jqiiMmYHWHK/yynxJYdMI6mbIcFerVW+Wyg2Vgm9m9MlbI+gn
64V1fZwM3PZGt4RwU1ruNn3PkkdtCrqspRw6M7uU/1IRyZlbfkuky2sWQf9nfG6G
3adCiTRxchTngLV6YB+yIcumOVSJ5dTtMOdm38Xt/reosJgvzy6kGuVLDqBoHlro
D9ADk4fudUx34MOVpvLLTsFsGLkKAjwPvQZY+khxBOvtvqZRpBoHlZS4c+xq8zk3
ROu6BsQbjUyrLbr19eR3XmLm+MJ1x8SW5ZXk6Kmz/vSWHthezlJHo9nnAGfnD7Qr
2LdidBUH63Sv1dThVWx53faMCuQky95ymBiCKRfgx3+F57Pt+bSHFLjHd0bbmv1t
iKBoyLoTDqozQK1mOsPaRxUChHHWusT4oHUtET++VpO2/iAnnyJHiAZ2Aak6vBCe
PvkXQmzGg2yxerTCAgQhtwrFlBHBzQeRxqs2r161AbYY1Qpn4LzGLU5MaSJdiDxJ
SJZY+txt93y1jwfg0IawSXprDlNNNryMDiS+Nr5fResB8C4+oKPKPib9vgwDDFbQ
/xkWdoXstJjbNZLwL8GxDpksri0fBKTymbPZCqQrzMvaR/T0tArdToHgO4P9js8V
dlK/miV/0lxI0qJ5oQtZyKdneSUgZFNepO6ZgdovDuypEOYZOvMyxnmF+vB6zt2a
nXU1KUQijZcXsJGtu2We4KIrZzdlGVqYs18CVFxDZJp9LiJP6nr8WTDdWOXSaym4
v/O1G+Q2m9dkio6FP21WtxjYSF33T1PY75iD8jdkoba0qPFl+uCNX2dFLHkk+pSE
DczJZGqUGI5QxHtbNksOEvbxdah9PVDGxWqBy9/L7ZwJn21/5lm/SYsXyxd1mCPt
nrFPoWDWgQ8PrJnl6LnBNjRITILBdy2ggTWuOVWLR3aXtamq4QcxQ76MkID5ghLy
WmJp2CP8Lw2Q4KIQaBavy4wpVe3V3AKdjkcL7QXDCkQAglnKabKplBgz1cSQZBdD
BfvpiMc8W5TPgAdX6qJ3uh0PZka806dn0VtE+2Krb2BN37ovq8CSnvd4aaNSlvvZ
5AZdc1yqW03LHn8kybJht9pfNEMa6WmWfOt0ui3OMGF7MS6DbWGwou4nwGhKdeLP
wCiSMLnLtCNK5vPlQ9lnhRLpWMXhfem48S0wm9t1O9HR3obYU69DzhCPtJhZpGwm
/9ZoGMDI7GYokIfXQxESqf6I6DMw7Y6MNVqJG7pMPRYi4in6/kdSrVkc5UbLkUw8
5u9d2R3k80sAs/SedKVVuXegqapGRC7HAlj3EC1HFowAIY0IX3Hdvoqd0kYuTEnc
cjUsTOwFGrY37yAkRFexLwDQDl688poQqABbNCvNTGxhKOLJmg/s0+OxHAEM+CM8
N7j9E4fHkEJXfmw8YlevSG7YJosASzMzG26qKgxV9BUAYCFkE0XnB8iqf+mc5Dbg
Z2FIyIag8k9BVBEjvfPIOoNNPQFW0iQS0BNUundpcVD4MQ6uVOMMDtg8SN4xh28P
wOoBS4vQPq5VCoFYj027vK0bxljU1VWvxIOtlcUiu84tvjkqBDEqm6D2vOEiqrSh
K2CuQA8uisZ5+VBraXQzgmq4U+UhoXDVsdkQwCe/lwjrXeKooIVI1MYFeecGIADY
NOBnBumXMy1aTlazVlYt0LlLNX+89wze/kZoDkbVOP+3fScHTu1Y+gfApL1jZZ18
ll4soGDsstazl9a+CPvF70lowdzSEuZuB+igkRg1OclRzGSjA6cwnxdPq+ef9mV1
YgVN53yHNjlyWAKAngulX6EhLCKvGDCB0XsWEofJmL21yUfUmqHgCVTBZibYCGUY
c3XMPx/tUWX6dFIa2eCg8Mj1rIGi3WUtXBK0nl7k4viPxidSSaGUGpX4eo69+8KV
anyps12f577XhPRzgkBQitK1RE/8o7fJaaZEhDMnr4E7YUME0H6SeNKW9fhh3GjO
Evqj6aWS1bhSwm6GB0FqTURYxP/TKaQpHvX3fgfQ24ovz/uzkQhTq0iaQNWEYIsK
kK/H1+ixuek0K+8XCMGkTh7as0DMJ4zmj+g0QmTlqkc24hw3a+s1VaiQFPBo97d8
fU203R/nmV7rmfhtwYG5efTWjW9ML723Wkp2AbzfJTSQgUa5ImylM7aP4m6a6QEt
oxW6IIfqJk3w5Y/x8qQKN/chn10GCzrZ2S4EarsYzEOepLLH0lOl3ZqCTuPnUXnO
YevY/JsimfZ7HVjtpGtI04/dTUhUGpnN83sWtMltFngZLUefFK2oePEdZ2p/0e90
4TgDksya5e7C+eAdg2tkvP/gdnmFMwoiJsLs0hcUlUul4br+J6DysRb7SDWSuMih
cvV1Ta0oe/ue42dYE8bAargXLBM4yyQj4/mtVPgQrq7ALo+Z4eBIStf+ZkK3kZh5
oM7St9a7T9pcVm4f117QwksLRWuHSOlsyu9E01QT7lU/fw6x6W1n6ZeTS35Z2GjE
JZXf+VofAiucv52CnGED89YgA7G1X34E79G1Yb37cRBr2o0QtbrQDriHNOdG/Mtg
jTTz1unfULzcB7gY5tAYF6i5pF2Ed/UKqX4GIQbpDwfudZu6ziEcGr8LAQh3EOUi
dE/8LEyY3V5X7Lww1Z3IerqCNUeYw6XzL8AAxLcBfHxboxAi8MqZXzxo0DnfxWjL
JLpMWR/GQB6ZmBbWw2LKhVMIqF8ybZmCJa2zRvR7hW6HAfmthpJ+LNxrXwOOx8s/
yspEosYsTecg+DCH6bHwHL3bFV/KIn8fi+3oNpdwuXW8Vf6mfTim03KlyI0waANX
cEm1+q1Eyi6EfkOLy3/mQVWNbJ7guJRoD90tB+WRLoBdfICOCNvihj8o5p2448Az
ndapG2Z/3YxjBYT4A7M1j7MQtmnoql43tERW5kmTmj6TrfXcTg/LMFN5Ac6gugMS
QaGu/eJan0R5Gg+Uy+TgFilpzanHTXiOofAoPWdhqL9EOvVlP398bEE3Z0lRPfo7
5HzTkBzC8qO1Y0nszbsBRMeuVR+F4xflSc7HBFf7sluFAU0xcCxkC+EZ4fPm0gGB
uImr4JLaCegIA2TsHCs1WRX5W/zgTjNoOf0IbbD/OBiTvtGaXodSLtCWahg2RhlZ
oGb4qwN6+ffSC0PjdPRisUKposUBkC4Ekl66vmcoTJxD/pcDC3yYUXNgQ4I+dWIP
lYZhYcEJDJH9g41EQqHqZw+Rqw/X76FKXPn2f/yJtzJfLiDReAYopwfzER7QkKXa
nzFq+j6839AH4zpTtIHmmLlGQAYIOnOzp/bhKAL+HCmWGHmnQ/mTUwh+Tepw0jdw
E1hWmskH2S1w57+ZtH+kxV2DjCNgq6Sphk84WhT+7UHBWY/1qRZVcA+OnzPMCyo0
uTf+CLWSG8CHdwjScVdJwF0hlEmAZWq6nsEw58nmz/A1KaGrvr3VIQMT/CbzjsRj
2J7hn4barr2R2utCX1G9Zq9aK3KkjUluJZ5j74pmc490oq0xprknCGSZSw36iU+r
ZVM4H0331CkWRsGz786iwDCqa3q3kKh65V6zYuOiXh057zAi56AR4H7swuVffTMc
zhCScrgR2M9UE9r/2nYbprtoU/GQgCjsVOiN5ZvSlNFfRKd8Ikse9gofdvQ4P+3h
sKOkdKtVlnY0LzcghY21zFUNWiyz3GPPwlJ3HZmExoQjprP+mFttNzvb6rdYsAYT
J277WrY5mSEtSl7OPYIJSuAEQEKxPESJl90tPS15njPd6DMgrcv7HD4LA3+y806m
2ccRTBDJHyVWrFAcM1CfXXSV6LxZ71DSo1gIGADdgm1J0P4f6N0Xu8ChSs86h9RY
c1WtVlDKt6ai7OOKSx1GBlSPpPDoBwfoXOda9gmwFu1gdK+j4lFemIm01FiN+ZAB
3YyVH10q+gvUL/pH9K57mc0ph/MEJK4MccLebDXal7HCqtPMdJY7+VCU54u1/oum
XXML2MX7AdmKT8tAlYGwma5mrNHXTVYBs5D5ttblCUTCm4l4t+K3hne5/khzB4td
rX1wzHTnpWrbs/JaX2su6nFsgNEolb/lq6GAcT7MI67OgqeHbgLRK4XnczM+7DbI
PKOgn0xPZfysQb9ODOUtVA/S8pRz5ahBz5dJAGf7hKlcU+md9F2WBBFRqtyahe4L
J0xMwtT5mArG58M2v9AfEBGIsAkVpGJ38I8GEDjPi6VQdG3uZXOQkqj7BxF5J011
f19gypgZRFQXMx06KNTW0itCQlls7SlKqZlYjPPIXgNNYwUKt0KLPiVs6PdW2pLq
ZZ5pzgtg3/Fp1zK/ceGV9d4PYF1hb18oK4t/csW3f2DybDlAycX/Uol9Ev/Ii9T2
vXkRRXeLxy2p/PZd99gROeDlQWfcPT3Jc1SrId0UbkOc7YzzYfDx51GKbLLokkh3
wu4rn2ay0bxf7702A0bF1Ylbzu6QHtmes3igAvJxjQJNpiUNWYdlmuPvMC53i/um
5aGn4HkYTl2I9RjVO088R7FeZl1FTgrGANvaxCdBuOv8kyy2DmYWOocH+nDw4Uws
MTPmXUnlq8gIivEFVsOAAE1EBt5ZvByK0jzV8ZSozi2X+W6KNHwUiudj31HC+/Gj
itsUAjXVJS7Or0TIyNSfx5alkHFShRQGqGfCJJicPbCJbwfOkMhZyO3l/QKCoMQi
iD85cKVlmScdd0sA8Z7iM7uY3mminL9+EbpZMDuofVLrmlw7YleNmx2GnN4tX0C4
cuCU++0VP9XzxYHy1XSsoPd+RRUfWnPhWDTbSY3077HvL25nlRwiU0b/bBDM4Pb1
epzJ1UdGGQQd34RiQi4ktoliNf0DalxNITH2tGCqE23/jYTTZPY9yQEB+HTI0iAE
swLHKGvL/Qd2mVPTlGOWq0/pduBNjyyJ1l7CRhXwZ/iTUkXPBqRJLMlvXzOBiIzZ
aKlrO673YDRNtaMogjvwWSVZ5cgqC9TFTJFW2GXPGGPt+LuzwvklDe69qAUcxIXd
2B1XqCYg6DxjMoO8dSCYfwyYdLb/E0103np+fEMY4eOAa62A9k7qed1geTLeQBh/
KK5JewdG+nhQminqdITdwvI5im4YOzZw9JJGztxJC6bd9JcnK+7cjeYr3Tcp21SP
7h2d2niwy7kZi8YNeuIZkC6MUhIWJnYKiFbnWDHVPo/SkGfWonxEpYSQ6ITMPxtK
02zuTeF7UN7ybDZwx+Sa+VTjOqEBfXxuYTKuau5dnYUq/t1hTBPw8o24av+fCjpu
jCd1BDhCm4r6dWzLVn3PuKlJvKZbvTybc9DWja0sdzLvH2nkAqisadbIYLImL5vA
6QxowjsMu12R92y9mIa063RRBJtP917JXiwgUbhWaXe+bMLk5oVF6Jp96iJ4J0z2
iTGajllHDzPAyc3reaqChqAdqtqJqUxH42RXpnLWG/bdTei2x3UiVl0FzSVj1Pw5
mXJuhPizdkZOgZHRhvDThCjmfYleD2H/5yySr52eWWHYLMi7Jw8H1eulopxgV/Oi
MPidy/zNETZO6l76i3ayJCHl/oww6+/xOvhjGfZZB7jKSqR0abLW+hC1HIrGBsqV
FCn89W4lRLtejd7L+Gz1a5S/sL2RXdjMBwgRVzr6JL5zMxHRq1tSkEdwePYrnhTK
lq6ja7no6/rNTR7jG9npzj1C01fvcWyJwmZ80gC6ZX9maGGydGwUyfBU5C8FtFjU
eQBa6MgnQHzwHHVQTsYVrpkcaCf0KSTemIqnR2o7qQmOHL8eNBFjwunwKG5BI1DR
rsU4amqKsjSm/5NBU/V/GVIjc/9GPOVrQIFd7oD53MUf64FS+fLzY0AYGOku1FWd
peeFk5i8newuo0w6Vt1sapHynL3MXg+uYLbULLrSR+iKySHzLe4QpLipSPG/i7jk
OUmGIE16MyKeHwx2dx+/8DM7c2oEqKavE6VUBySJ/JP2bRFg42sShM8YTQK0pIgp
05rfQbdVv4TtYsGVvleUCms46ktlZzISJqN/dTFeqcFztBnX+jonmFhhzTFp1dOw
XELWX6McSskSn26/r9X+jWRrsEJJ0fG5noE1/vf8vlKxOsjZPmqs+7p7JzItL74v
KFTjvhxLd1pz4X0M15HeoOfdXtH5LWq3vAEDEc2foX4r6jiCANdlKhYQXfvc044y
zkFiBUIhzj7lchap05y/TLR2I8EzyyGG62J66JoOJKfAVKU5VDz7sbRtqPnhqp1P
8H/j4UyEr5SZQHN7Y7ili4byQHa9Zbe6fo3e9Xlsf3/tPxaP3bBanOqFPaKusuXT
YNzrDF2YTqm1gH7LihJwb3bB0CxolneeNzgAbKKcsbPwQ71og3wUY6qxdkuopmr+
wZXGzVneclZp6Q+Z3AGOq5ni5qQIfaTfB8C98uOmSKIqv/6GNJfLpDWmEOKbloHc
+4PdZlEOsOqlpkQQV0O2MWl2sDOvedj9rNV4F0dn8RjlEZgnHeMhIaumoxs/t/W7
Kb9k8LxAMVr3Hxhzm2soyY4WSSGRkE02sfpuRg5EhJsyW6oFJIUk6T5EX/rIhu+u
ezl+xFEQyIzaaYEyz3UT9broCVMfY0Em6mDtjVGsf6c=
`protect END_PROTECTED
