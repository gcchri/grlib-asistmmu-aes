`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i7nwVgSVDs9a0i0ffSnblbbeAoDWE+FIs8B2ZxSTJKaHYtId8l/utZdcjk9SVbU6
Lk6LYjpXA+rkdid/Bn20WPb+5sataeQl9szpf5RaHSR3YMZB0u+3SGnOOB2eitQV
SoUWpAYq6AE0Ynguni7JtbtIwI1b2v6d++ICK1Z5APeuky92biJcOh++LzxwxNvw
zyX5iFaroe1uoOnmIpBYNPYbrc3ehV312hB4hHPzq1hKu3WNldanfETl1RiUCqCq
8sRLStL2g02o24PgiCOKZikHRhivna2Q7igPnymEamQZFU/nWtmHLuHFT92FvuD1
rGQiqUl2BEWzAXqrZORCmNxv5/U4SO4E+nNEE20VK7p5j6lGb+Cdr3fmyBAUcxer
yKjcL7mHGjPvkpSx887fcr6ASsZ5XIhLMc3OCq1BkH+IsPmyXSDo9inYdJqOywsp
YcwI4FP2ZVz6peUosDkh64JdeOEQ1DzRFIZcaV8So/fXX5duLyP0GrtEHouLJAWI
jZ+/rHIzNveH9kg42YUfx/FJ2b7wTpVEvAXjGAjVIyHWQGKnJ6aXu38sabjMp15N
MTN9vOAXM0WxIRW7NY+bmm4kHQ68IfSi7Fsl43fnwzr4/PqpO/GvhbOdSjFn6LJ9
hidJIZEXGDX7tpebbWtnllRiU5ZRtGxR5NfYw2msVlgHzqTnR3Q5Qst0vEn2z5vP
UNeSvkBjClBdojOtR2qv9HcLu00VdkxbG2axIzzo5ndd9r8Ho6njbHorfTR3j6OI
VMpHPJKaaCfB4wrDw9zzT5iXIiBI2z2gz+cfaclZ0n9/n0Fs4BaQEGGLRBYmL2cy
/PAjstl+ZJy3PC8Xl6ElBolJ3Ngke2dedKZXQEhIG5SoLI6SfS3Tlon/IpZe2BJQ
36wYEbdbdpksFzRrm093DPWXu8/G1L0DCDDckfQsSfCt44FNmlLLLwwXGsg5kETP
zVBX3xODy7ynsUwW22HljqXWxVosiTN7n8mN2K7veHRVVJnlAinR0Y3kxkX+7JOZ
nEUUc2FK80W8Fd5f16mzGyuQJiWwSJE3VddiIDaW80N2/GmC/RCXHfQrYksfe2uh
NZa7Eio/ltt7Dyv4IBAnjBcdpR+tGgAVRs8jCxgmNQDkTpCjlP5/85D0m/LPZnXD
+FR+zpPIeVFIOl6ROZRfEVUppOc83+GwyCwcurEJEFaq4efA6pA+OOOnW1BO3jEk
8/L5ywCIm+vd+SQbDs0O3t7QORFRPtYEXuDxersAE1GheWmj5/Ylz/y2/5NWa7Ih
A1rBKvZ6t90DQb9k6EqaEW1+QUUhwhgEbyxggiX4BUzfbW9quZmiG7KrOvIf/VPl
v+6oWuu8xCoVw3eL5TbmUCIBJ0yU6pnCT2QPawJTLSQKU9ppWEua7sOUSo+2aWOC
3zOQle6g/2O3+IJSTnSsb7Wop30/r0k+VxMFiopVr8iMXERxsOY+mT3JaaF6exI0
UMRe4PfbuYq0WPKRzfjPsL/UQdWD8ZO89omvX91RZyJ+Qko+4zdZKvxYyR6IIPzE
Vo4Y7XrjC7wblKh+nlx025sktYSg6uTzQwBmmQBdxt8YV/ccetC2qBTm/pZXcOur
AiUL7IQC2sHJc9K6dwm282UwhDsxH3Hf0eIFwFys46/BXloMoD/tyTlVjfS8udDA
ItfXeLniGS9NNKXoBA1mt1iX6LiAjL3hReci7HokPQMetcktocNtjcVinshLoI6P
LnhZV8nYlRU4Nm2wiF91fXDuBo8X3S5V81kfGpriYeXMdDkvQKLe87daTmYB9AlB
nsYcX+aBRe57+u7WBTO/0GNWEh7sD8WQAgZGWZv0YkahVarqxnq4CTFEi7f88e6s
wCKmTQ+Vlf19yq9d6x1FqEMloV8EULxl9dCYAg03Vbxk3FSc0v3fN9lAMMpZdlys
OhEvxWrCUpCrR9OlH778FY8oT0s14P72Ze1sv5AXrEgJXmKIn9KdYdaWAMpq5wHs
PG7hCCZRvNjs+fhFCp9jwc7n+dXHZgXIWDNq/OWz14c8WYMywWy1dL8obTevWvBP
T8rCxm/2V1IE5QVLjeIVYMKj0MtIJihHktQf9sr8/LsQQAnJ3gzuNcCLL1/t8fg0
nkcXPhiHXgHU88n4BDxdbviDp+mNqwapa8cnXRQgsJDzCzdk2rOyFG0noKg4WoJ8
Qt4iALCfa7NuNzXFi1N7+H1Q1X/r5hsjk5Eo3yyqAxg=
`protect END_PROTECTED
