`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TfWRsJzYRiOQTP5OzCqBGK1Fyn3OS6g3NGXxGK8xzmq/bHaKih8Uxd3NfvzcY5px
GfTAxq+QRcZC0NXysn96D+yhQeif8p84VSCjdFBqQ1DBPZZtZ13pkuGcWUJtG4k6
UWQKKXo0lH/vglbUJccgGR1fJIpA5eCDiyLZRpjoE6KeZ7vq0RvQBN+hR/znGqtD
SchQxpkjSXAmVnIlXUKAGLRuWtgJMlAAOgz1De1r3z53gmhkn7dxfnPkd0OiSSO6
fsDMYDhJ30Z+Q3oW/XO7UK0yeaiA/9k74A7pq4Qm+hQTwZgJGlEpwLESH7uzOend
psXSiKsmNzzYBqTZ8WgQjeGfcsmTCQk5w/Z7BX4+EZurRMegjl0ISuM5DQU/+2wY
sbEEHUGqXlst0EG1kDSQPJu7GxeM2Xm+9ajospjwejCARtxILlbItGtudHbKlEz8
AjYIwIbmrYevEp9nKcFJLxNfC/Tk3A3onsa87VPHYl8BhKGESCnxcbhk2U70WMdi
fW9VqPWlMyDHlWHJUK2aWKVviEAWG8bBjguS1EtKJbpVTUj07xDVNijdLNfqq6/t
xbBbbzgURrWRD3IxbuLdUJrJPBfH6e0s7X95d0w/5CnpyHDrneoJVNP4NyRuvm/z
6mwTe5njtcLs/70NQusR5te71te5jrYrHEWQdSuJMwp6N6FYnhb71SGIvdz2Ms3V
xWCSLf2bTnRfpu1tiN7PzZMuj1tZSZkjDIAGqkRWteLHEmslfsNdoOe3Wx67PuyP
JET5r/VnranVYjus4wUiWNeiyV2JPgPziskfL8fR7IGCu7a4aDSxo825tyryIDMS
h9yGyqCIVGBsSj1+/PaIKMKBVTQGIEIjXyaWzqpaaXF9s4SaH1I6THg1yhdhYVn+
HBMYV+RC4VZzvhr814sk3fAs68aj36Jn960HeO1QsMtFOPJAVDtrPSItEUFKKyhK
h4xCtmBoxhkTdHIG25WcSYMSUT1YumUcAza+F9L3UBV8rtNsnD1vzx0PD45DF4JR
xSw5usHQZ0KBFXQlTHsX/FcMon9mzEy2sdLQ77hQLLG4KdJ8lRFSwYndLe5FM9z4
dfQfRMdo8dmjatM4Db+DHM+TqfIsda8G8poGqqPI0SEjzG0XwrAXlYBNPETzrB8Y
a2AbKxn4vGiUOmc5J80zzR4edaY5OQmj3G6cUqUpG4sWpKnenY2kPxVf9dhcyNJG
9GDi/zF+F+dYjqEfJ2tyDYC0h/AgmSPdG+rVymE4607UJdtzQzpxEhw0CubenrmB
8+TsQmoAvW95QnUzEhSgeUYWoCU/ozCsYPsv2yZWaDRlFivt4kFFpqxpQrDFnPQI
daPNZuPfH/Yaan9Ih/H5NZSll/UcnFUUPFklRglJDxp3SHornbdMjm5GbjxJs72g
bFrID3tUcjxSoV1mm5/B2CRCvGmj4iTn9JvGMaMzaEFYwNSzAETZ5g/NksQQTeTm
qhhQuHOvJ6ZdBiZdWQtXErRMD0ygVostUPeU+fxnl9Q/2ZLHovQUkqlY13M5w36z
d3zkSJmhGSNHj9LHw3oKU9XsUyDOulo3EPx6llc0pEJlri5s5NtZ9E2r5tuuE0o8
LuJF3S4DIwBCoNECa2HLl2XDupjwM/ag7fQUkKpjP6WDMbwpe4pc0RW+l4MQdLEE
Ma7Wult4RoRFMUO8qrojJVKWNTWVYkDXjf+dNTdx+ble4xf1NBGP/7XaNIMvG63h
H/C9DPGlBxgijBfmnQqzOb1BdWAQogUAf96NLObgZRhgfHVmSvgNqRbNNNuD7lXK
JrRNo7Wj1ndyilhzbD1rMSKAYmKAQAS/Ayr6WL4XzGyk8DpXgPWYqYHMHNz5/7sA
1J4HbAwjKlIQQGrLVSSS2U0esg90gd9Vodedu1DKKZ/lu+jwk1mwHgK7tnrWAhBk
OPz868a7153ffoXunyhWbfNdPsgNg0ijf0OX8PasWfU+SLrSk8h1m6WVhTq0sI7X
uBPfZRZvyQK6s/YbclV8nGKZyDoBILfnUulMglmouN10tgopeXT9nHaIt86X6dg+
0f4D+XgRSDHiKIG/C1B8R5es+UOkGmU/KRZKE/B6RxtJ7fz9MGCQRN/B3BPc3zhk
ha465WIrOLcDdnLN7cuHQTOKwBX8xdjEk1cKdU4KdAj514PrQo1c/5ajGxys9A+x
QFs2cCYCMLx5JFWNOuxP13meKPU7R7gCk9P7q69TTl2Cojpw2VzTOyfwtb1W/8DC
DM+p7aFki1qutA9MNFNOEp3NA4AiJvtYSOhQmbAcbCCKhaeiefiAE8GSvm/sKSp7
5N6Y9aIuSYkVHDRaCKUx82bz48x2/Zxkmrbq61ygDMPDEIYn5IbccYgXKt/wIwm1
F2+M2VMG0nb0Wl7iNyC44Pf03egDqnd50HXjn+Eldxjbd7cni9Mt3OQlwkmPIblT
EETRiG4FWNSk7Akwe1AxHITHcs6Y3GNodi5ajzf57SiCQwMPhLIOU8VSWQO1xMA2
U4FLuj4q6NRNHd3D1huZL/btQ4gJWcsKVYibyuB+AFfcFTR8n112BkNNGVmM3xJU
Q359iZMVk5GZySohy/GhyyYBQ7YWm733Ys7WoZU71A3SOH6owVpYO20XSsWQF6b2
C4cI+o4VIXYWETNyK9IAkdowF+96uKbMxtRPpA42A5Cg8iY4eGt76IcjizMUg2Uh
ixujk6Cc/7yi0likhy2Hd7eIQtNg8u8LnnnDMxYI3nvjTMubICXrxaRtox7hMQE/
9vImgNNCGNgd1+S7UI2ZvtakmwtHmSNkuamWWPu9dRZ1UvAWQK2vY6xaZpYjNN2a
PElBdJDwE2/kfAsslp02SNzEwcT5SbYPbiNrZX9owL5ci62iSRE2u4U+yc1nPzz0
UiI2/QobyQXqJd8/GIX8wwjU61HSqNVwTy7Jr4cLYqIL6b5il1KzEjOh48Jw676K
w5VVyJvW2rK1WktaqVl6hCtMctHdyTnDDroJHNYxCVkBW6xHfT+slVMmF5ZcBTsP
gvpB1mArfOPSKUZ5Y5BiiTZ11u3xGgLSdIK4PnGYYEiPp48ciw8UZ0vYTdp/fxR1
+xOs899JblM+5bSngNoF5nXgZFeriHs0Y1zbp8WX/7vifE5yDDsZzI0vSOlBsJrQ
99QzZePu71oatsR3UEDm2xeSTzhMIXxUjmCR+BoNO77+UnTj9+uBmvNsb4uwLgt6
HUZmxaG0SpNZb8VRLaGo3oTQZowsidESyR07Css6oP8ak7iL/VvesZE48g2mW8k+
NmDV0ju435LLS81pFrgYbdm4dTyiVIM6+Gc9j0bm0fzkyD9DOIKTCXBbfl8xCQ/C
s1Jpy6Uf6lSZg2N+Z+wCwQTMC/eJtANVMCogQtvvqPHaV7WclrSMymLrM1KJApI9
eqNUq5IixqFUq1SL1Ke1NZEJJZ+LiFMzIAD42bHwCoNrYXSGZ4byptZUp/8bDFdl
3fzpECQb8OIsa+5FTdY+JH3iol1mZU1xRcgkzOO358f69tI9ZFp4wLSG/bR7ahYg
eAUJbZ2nLv3AjVmlnCLpvihsITQQv5ZBCYzJ1dfAQ1QXb4vR4xHeJ6pUExw4gZUr
1tdSem1MPB6nm2/hS0esvPtZ3dk5Fnr60sxkqDOL23h8zLpZnzpRvPZKUxElI8Gp
wTIygE9OMPLN4VNW21pmrHGbUinBsBk+dvxwfmevKGhiGH4Sw08DsGnk4KzTrNNC
RNPMAgXJ+ARVlzfxrszU0VXGzYH2VWCeBDFM+Mfy7xO2xo+OPe8d7EZZZKXXo5Nl
d8z6mjh6KNTp4Vmk6z4kxJ0kgjKigyVYR862tuV+nGj6/gcP0e5lwQ8+oagatwaT
7yZg58RkUB1cp0RPp5yC90c2DE78WuFb2BHHdi/l+xJwbWK9QSmWvPCEtHXZj93e
qV+gIrQ5NuZdgwvozccom9TJSXZnbcZmyydrjkFgAXI186MnOLcYCDAnit8PyXWC
Foq+RaxvGhTrF0kjOAprQNUKY6yQN9jhBVRcBNSq5PRCCfIEB04b+VMBF8wJfDAA
JSi9iEbbBo+6d/P7C3b05ZES6bWMF2bUXE+NWpuvkHW6HYPnMkZFc1JdCtznEwPa
u2L7luAoozIScjfaa7hq9b9TWokx6l5qHUkHD5YSXNj+bqqdYd5NLg478AsGkF4K
o5F3MPLtmASNhdmMufVGl1xcFlhJrejtEFrf8fvqDg8b8kezISJslmxeajMn1X2P
zlCor40HDByyUPgLAXHeIxwdehWSU/t+Q64g9ZzoWck3hNRD5dNsTV206xcAZtQq
TK/lA8yJRvp8120bprP2dTAaXL/Z4NTcnInsqnJo4MSlSOVa6C1zixrJcD12Hk6i
HSGC8yfLz7hguSS7jQFcOCiW5wcaFLIzXO6oFFmt1MIXkzCPGwCo0cykeREkPBn6
0i4tCprbgLVDL3qVLmeoq0gBoBk+kq2b0PdJN0uUMs0/GXQnlz7vWQBk9RI8ILp0
6H1Sj0uiLUDj8yuyFLEGyNlywezAOHKXcmqpPn+1zkXcCImd47ILTfcrVM34KGsW
lSaFtY3theAntxeLNNKGSGsXah75VG32hm/WnNTgbsO8wACRYMytjy4/422UJiH/
LZbLkS51kQLSRA0s6s+SyeRVXfi3/c1rfy2K8ljTAmCGO71lf4U8dXZXPwnQ70I4
Ju4YiP5JPA4ANg0t3qAv0aAnW1oR4XUzgQ6QVWIN2XEynMBb/HumJn4hZeo7NGaM
VI2Fnz27ONRt/Fd9HFB7QqH6geoVjBe49RIXBqpzqCQmeYrVfsqB3A+QuaYOVjKp
R1qE3uMAv2oPXEt7SPWHMESbSSb6afZ7GoYa64VxeUErb9nNWyzsDqM7B9FfQTK1
pw84DL30j9fIvVnOb2ypI/eUEOC5wIicQhHGexZm1gBGYGeMPqDtfUYspCkoqWSk
vBhiGKIFKJ3LUQBw9tqt7A1J7NLiJH+B8SaUeI0tzytpHM4h9aLdt/+1A1E1WiUG
5GxdUQ6dj4yKHx8M78g2S4hNSf2RCOMAKJDxxa2zkrcC8134VK0XQB0glJmg80I/
UdhS+564NK0CYhcmh5F2DH2gBg19D8mTiIrLyDO/LlIcRV6b5U2GJndqMLrxlYy9
e+F6DlNdaE18EDTj9QWDyxBe/poU7YxvfvQSwHIwwABO4l0vqU17GJrCdKWZzH5e
kNAdoGwVq0774uVBc4P3asPup21rUNzgcpuj3uutJIUfLdgtOGBTLBIjtdehvQX8
aUnGG3L89JnlsgWT/9l/+CQfn7plD2wpYCX4mJdI8Ymni8NHY3iKUHYq3IK50gGr
w7tIIyzHoGXCL30N1fwCXniAii9nK9RsxaGDbenHgDm0peyng7yrducXQxKC/gKe
cJ2wfbSP+0OM3+Q3vgGR2FZtkHKFstM4Y56H4dSHhMa4O2+U8WFnvKRU/q0o2ABV
/HZjMIesrTZEhhdXOCGDwdzA0ZNHuWcuUPLHahyoN9mAUdUWaYTJB1A+FY5UnXGL
E2ZijLHv4x67MEIODJfx+fKDr0Aeu9RTF4gKKv9ZWYrhV6fSEJG8JClFR0l39Esz
8y3squW7BAWkDIY2fmfUdeYILtiN6ZmiKpIV4jFdJTTmh2i+hzVOeKm5GRol5ss5
7FVTRycqOB8mDB2OxmWacvoNuX8tuuomOi/37EiyeydXevZh+vp+L2STsVnclYpX
RB5jGYiJ1o29FLzC74vkLcFg3Sy8Y+uCuX3nQh2vNAtO0He3ckjfn+EgsQCwiVOJ
arThZq7vsFzTImMFAJDaulXfka71Wnm6fqpEW2/tr0BETZMUjfIoqMydl2sk1h2M
NYx4uOF0E3KTLOOD56uAF89JXROQLd0GHensfLXxipEmt1GINnJg+1wdYJ6mpaqA
cXguiakxiToNXvEWmlT+LfI838FJYVS0wYFtZiibOr7ObXrJ/R7TQ1NfBlt5n/J/
ho+J4nciOrpv+fErxcot5jFgoz3lbVx2lDF4YhaDfNGB4FUNX1+UQcYCr4RCVkz7
9s7TVwdxQb9wU3IOGd1Gz+gbAYPozcA/dJ1EXEAPpEt6jXDiVTLWbTdYjhyAbLcb
7VgQJH+YRQTqtbJYeN1n/1otreKs/dqoVcfMeh708yqvu+QT2Vr6tNl9A+q29n3F
ELNTiuajnfnDjUR/AMzOPtJzS0zJdWKzET/rePZ6ManjCrMgJ1ZLl0WwNfln7Xhn
nrHd/YQLoCNys4rT4OG1wd1uQQRom4uG+d28/CmftsunRxUiJCVbvFR8xoU4Dmoc
Sy/TclwhQHlqBii0VRsAD+y0Fwk9lUkZDN19ZHgdrQoBxKUi9bFyxX2x6Ue+a26b
Bf1DaQstW1JXM036RqE6U5D3cRgyaNTLGn/LuxCORmmwCvjE297HCpq5UkVy0bM8
5xrls5d5ze1m8zFuypUUVzWIbgQaFpAmIxAAYiMNO6DZgpeuwAdcY8OZJbc89272
Euo65p+2kyJjwnqysA9OMEeC2qx/XeuWJC1yEWgzX6fTMyUrHAHdx6Mx+N1JwUXd
ax0P/5fBLF1BsHORxTHT1sGQj89TEXgDaOi/giU+tXNdug/MhpLZ8DedAnoUt/gV
mAml3PjC1Wv0fiQy+eyPHqYoJS+rddbIzHnrsTSOcQW30f1VYwxbndjEN+bZujb6
A8Mj1e6NBxJPL/yGmskSGEBgxqo4xxfoL593kcXVUfddFK9LG9/KeTuPBTstpv6O
mt/IpWedBP5Lrr78IrGjDcc8NwJqYRQRb1ht/SP7tGCpX49elka/zs5zxz8QSm+F
arBiPZYr93x9vCbIWHUF+rVVbqT/3usPLHQfmP1YheMgHagYHoVryo8FWgMsvQka
vVuu501MsI01ZwjxzjN7DMBfZhZOnVsyfWl2xZDXck8U6nTYshqoD494MkJ40jN4
DAu4ueO8HrJC6RR9tHrzJ2CfQ6qH0xB4zoli4RpeehgPDFKX1Np0In4LFP0ILcoD
eHqBdrfQ0VlBvyOcFDzgVIMqDZVnzw2cYnIscCG5j/QRxhE5pfDJOX4jOPD/x8Ca
k2rsaz4Em8RT/hgmFx+sISxMgrrld8nkTEOGrclwynViZeDaLt9iSHNUEo3QLIPx
7B/t/U5T2YEHwI8Je1dZZl0+VO9vWXfeLw0GpE4kZdJriSlNYfFGdGmHFOfFnHrc
6fzf8DZpwjx+wSj6h33IYmnUjFyLjv/r35BJgi3nMqmxeqB0OKybWJGFlB3VL9T/
pLVfmlBB1/VB93ZyT2OeSM3ss6KKDqETJyWNbjXbYoc1xP3fNL+7+la8JGeHNb44
eQBiFusAaOaflExOF1IxS5PrR3oMe/Mk9qcCjlErKddG/hHCRcAilBfjCk922YUo
sWuvQVV8+mTHSgv076ymqzriPXrVVheyQQx9MFJu4dfrtNLfXA+aSH0904VwMb/H
TOL7mgBjRgi/1wiTHkQy7nNNBcH4m62riTpTD4kzmpb0eFTveMhDt8Dgv6DtPZLE
T+8jufukMro0PbqtgX5c70a0XXX7IAcLauznEyESiq8ffokVcAhhfuEIZNc06GE1
dZE9xXyJvC2z/2i4eEEEeAJmuGO2zg6jh/Clv7Ek3EPoOUS5eI1g1bZlDKxSK7ZE
KLC2xE/ZjLmacTEI6u0Y3QaRz6cv4DMf3iwjPt0j29JTjL9w3Mf8GA0BLjqRnUrg
o5sf9lCM5faqqMTqHkORzYre1RFz6O5OzPiBu8w1mCs098aEg4xcFeX3AHgfN3KE
fYA2CeEUDN05516jq5R853ry0ohKBeIzhnpC+joewC4iYeThuuNtzhB7HZrhkZvl
auHhaMWQ5iqtqp+ZSWRItd3WlXlFlrl7ow7mIUNsraZ9OLK84t4DVst8qbNHRXrL
f4EJf4OSa/5l9DPJWJmQI5dEy7uIDAiYqbQZhNiqksz7+Nsyf7XG4JPCXsMw8H2y
UsrnlY+7O3i9sX06aKIIOq7lBQib3D0IOtZa8H9Ls/ozWmv7ir71lFJizZWQbiwb
h6o2XmKZaDr2IECim6inZJThf9okb4tdLtvpYGjCDA0y+yXlcd4upIONh/ZBOPqR
Q0Huq+7RH5+UIBXMbrLcgfgIJrOypT7YeEIq02nHasQ6p7WNaElTjzCcTvtQamiQ
Hklp3Wg7WRbZVIQuW7E6S7OT17HP/BfIsKU1V+qLekoNH4EhrTc0s+4xfJJybH0A
BEqL6pYTsbeSARsqC0uHTAwOlCo9RZMBNIv49k9jQvzWK4qXP3hh+vsd6QX9Bf4E
cL6Ojp4JcsT8oytSE9d7u2VwU9hnTE3xF8KF7mI4fcRu3y3KaZjrJeEiYsRwMbIu
yEmSehCXTi4PmfY4HsIJ6EQESbAQzsTBUOSMT8vZ5SeX9WMGlHAnafnfrHisn+wl
tpersTLy3TEqcT1wu/B6YF33K7+JBYC54Rvcn+w/IczTFvw9u0SecE2yIoSUeRbH
qne3A8fxmz/Iol8T1X/MoUHC+Xx5j4DZU+VUF14oVkS8pyz6oEi++hNyKKxA7ECE
bxXvlxa4QKXcNjWTqd24oFQLUyOY+qjGsV9/IRufC1HMiHhq4LAtMusz6t0cc7ET
O00GYPqkd6MvomndqFFnxN8LZdqfoMP2egJY00+k+LvdQ8vPe4IJWx7cWAiAOlHr
MCpxtH/buetG0et2R+SLdwChmva6j86SSYxCsH3uRlxm1JXBFulDfPhUzGuTL3+L
uUhqjCluUSD1KvOxWv4MABM6cfi97Uq4MhsUfvWd6m+8A1pxwqrw9SqVJSwkm0Pr
25fxQYjgi3X8UHkR1g5aFgDMTwEfgi53rb9mkB5b7JGVvm+PKFaQiv3FIK0y265X
+GO0Jm7hyNKCulx+wtCEUk2DY1ELnWhvCwQ/2/RsNXFbKyQwZiQzQHZS9V3nSXbZ
F72zzK4h8K+tawOUjxOnPFPZ31xRStOoIIxXiexK2qz0jgbhoMX/14Qh/T9rvMh9
Ivn+RJXRKhpKhC2LUiy4ALlTkqYkhUk8eMir+Q38tiVNMT+P5yM+JLaJYKEo6LCG
85Yy0ibBIFaBAg19PBb50aF8QdIDyqxZVKGc4DsVytK4RLKY2rjqaE9v8mJ3gNYk
1UbENprVkshA02pW0N8Gqyym27/J8uF1rnlM4/7qFGg8bCXeinplXNi4LRHqnAqb
lZ9x216EhQ5U+V0fEKoe+ekbhRoIBuYfobyz8N7vn+mG6vrhQDYwrQJrYrQh6Gpu
6FWrNslB8YCSsf01+UyBPsQGycY0CEmBBICLO2gymulmkq29ixFmoUEJvVuAincI
dLKDCDoxvkd618vC1e2K9SNGeWcJUM70UkDdf+YCWTaxbwUqNJ68qIv0ThgUbZ2j
vp+4ZkceTHiiIYO0mTRDvqN5x4InW0U+sGjwvD4zPRUIEoi/c47ehULmpiscWhRK
e8TYm8B7LS9rYxB5vdecpf3ibNupwum85jPJeInPb2TFAztqknEC/uM85oP6EVHM
GHxlaZffy8V5qChQSgX6/Z0/GYzE7oVGZcBfwSwue/GKtPhnhfXdEwWaKE2cB4KZ
BD+uh60f+98ouunawjllMd7kZm4UH8/oW8hNBfK0RsqOjCTEdRG+W+Oi6oWGzs3o
oImThplx94ShgoVJqKQkBr/e5QsjTFpsTfs0YxIgJTTVOejglQvceCZk3fuirp3H
hhBSzCY00EYiYOOMXJ1zHZROUe51Gd9xOzlQYXY6ZkHUuNRQN//0zlc9WsFUZxdZ
s2SkCgWS9fyPb35NSZXJwwU4m2V/VnBjRYs4Bd36K2GMbPdedQ8iwa+WedJ6hd6j
Yxgl7fVmO2bHqUXW+MiQH4kvly6RGGsd3FTvISbsWD1PYz1GNlw7bZVlDuJYNwLN
25Fok0qu3kO+E2EjK2XGN8yjrMJHNb8Sgze+ksgFv7zQmjAE1CjcXXsYkgPL6Zs5
DIpfE5H8DZQDmCIF20NA8/JCMHvKN+gwCD246Um+KN6e1iqIYJZrE+jqBzZqY5Hl
ai0HzN6ywF2WCMj1TkVre5jcrFoGXQNEa5JLQ4DeazjWlx9CVPWgAfCjFtpqrEKh
Z4tLwCXh1urxXDmDGzZyB/TB+sziOTkAoSS30Fvl6YMiiC1QiqUfgDoHraEs6UwF
4FPgnzqiqW6vGgpMAopvd4leM7UmtL9PL/rP08D2QqGqMj4pEQ+e6ac/AQEhAGEA
QeiA2dQguIQmXKk6aoOcDcHYnAi8U0fiOXrvnfCYtkG82oTvuBs9MEHwOuriQ1Ue
cYM4zYJOx2zRaGX5Xxg0hrh2LWirQEUOFKlxKrOzGOEBc7ocZ759K8tqX+soNJJK
/EC1wrDFERuV01T17z+eYALzKk3xInaNMED6kX/Dh/nAuffR0UClSQky2q2/F+5p
kl82cybhtRIwUV9FmIjFk9GpKzXLcPpynZYVuCyPaBipEgyQ3ADg5mJCqdR0QY7K
3UCrStWg/U3b2OICiRrqKYl9Y0Gvpi2dgz2QDEcEi0bGXaSXMXH4ZVxDitPCq77V
2I3MzWcmIWNbLGjCuMy7oJkZG0IIrmRNx/H/r5e+BqtbwpRaxJ1tYk+2dBaeCTaa
+7xkOWuJfXf6Rl/jEmDzp6L2pnxfSsDT5svgsNn6MhQvF4nrdw7n7D+MDK0s/EzL
1kvHGAyC9LzkebWatai71EzjGy7trFrcTCtrscV9EzqOO9lgjvrqhoh4hCwgZ+1L
Xj6rGfBOttl4nATK+0bdsFs4q/D98KQWlwFnJB9mk7UDZgznJTZfiNffOTJk9w1H
KfcYwPXPDd4NSMCXG9gA5bUQFMmXpnlynu0vcSsMcHO4kHbrYYW92rq5rdcxkOh+
eJRstLuTwnJXa5A53JTV8o72npiSbunG/S4AQGSx4M8z1QcOqIV9zCQ8t0haOG2E
7Et9hw4JJ+kCDoTgcckBaWkA808t545r8mJpnEpLSSBWVbLE0uBxE6szeUT9i56c
bhds1+kXnEzYOSekC/UZzjCDEEadkIVNe5KZTMlSb3qhNridlHvrxdwkKh/0efEv
uh0gwMQHMFf+FSlSdIXxWeV+8y2UhwuiC6gMOe33fTCFEce6pFo4Ew7v4c1TlydF
awTx8XGF14eE+Ah1zH83ipZjICPqqUZnLwm9RPN3HULSdsatrMcsGBzQQsRbY2W0
tOB+ip0jks9DSIhUTsi0vKgVIYz6l3nzp+kczmhD0Se/Ve8V+13cadlwRmj5vUkU
vVineyh9TuD/8Ks7LUtlqq3WVkNPZQBEmCd/4L9yj4lcs0OK4aPz1oxM5yt6mfMf
RfwmrJo2S0pXhZG6dycn1TA/RTK0oPUdqSpwkvYTQtswF7fVMLBx7Vi9GRbU6BIg
4iGSKqqEbjqkRHFKWRg7dwzYYrhcA/2aEdkFvY2Ad4oyZaBdbpZ7KyVHpzeS0U0q
ycGM1QivIt9iZ571UOY+4uQcMJUMFnOmiQinJP761NqHfpJYKkDVqiC51vR08z3G
Dtuf9kA9icxax4xCJ9pqQP3UOETG3I58aMHl1w1+D99EfBFBoHcEGAn0ZB2coAh9
/z5MypkJifA0p73dxjccqGki20WRmbpo9S0LPcqf9c8ixv5tflRpz3puQJLfL95N
8f1t6MpVBszorEf9nMm60vcS2aiEwgbvdjkHry4ZuiOmajh7LpMZ7mL9uX9YznRo
d0cf/yyCA0wmHS6kz/rRKJoqiS0ZXpi5AhwgAD6fR/QML8xAzo044rHhYYAplzW+
V128sIbVIRmpZVgnNcxYRvsaqdQDvImmcP2LMdjv/jYlMRNQUZCEYOxyagpJ1+UK
W0+JmuiId1EB6CV4SjWXesyzYzmClTeCEJxDnmtbY4gLSyw/xNNNmpnDRGkdwS5H
Mtlfa0lhrV9uz13g6fnQ3rvd4HetjBciOXz2JBVljrAU4Rvur9Q+KQUxeIIfkJRg
MThyEAmnJV5mZQ5F3FyUmz5W3g85KGrVft3Ay59EPpT3RXipxs9ckJHRiZ3ECmu1
5G6hdGlPTFxlyFsXtHHt/r1+HMmqGwrSWL2FaS0ALiRZJtM0Ry6IVH9kqEdMCAfW
t806Pg5V1j+5aJATFyf1QX2n14MMMO5hsC6JM9HHxUXwhqGGW9i98SlmKbfcjyKX
nS+ldh1BiYfKenmzFZfnKzeAWyTKkRqW0x288AOWUAH1oLPisV0Oy5wowtMgDRJ3
DcQiat43kmJ8KRMAaJlcz5oBswNAj8V5siJuNB1y5i9QBxkeHtEFKNf1NdP1qQmy
uLjgpNFmm669lQ3gZkvMRPnFkhrd1XdF1oAD9BTrOMs7Y6v32M2ie9Zduthj758o
Fkdpcc6pU4qZROmWjZ6Gkot8fWlrZa5eo6tzCi8LNQ13Y5owbM33XnrYGe4tU3za
cgqmBNpS2Ir3f74hY35qpioyCJcTolYZhExP3mTOj9ljjzb72QHmWm9J+BpxEWbj
dIawikZQCul73LiiBK7+lUqHT+xhQQRSP+oBgsQfcFu4YhGtdWN/SDvrgD24OAHG
BzcV/Fl7NvigcybuLJBvmTFlpnB5JZUZRlBOehe5r/npUUbVEHXpPLXmWCpGrv7U
e1VtR/IkDJCxn6cks6qvjrTcuGo+7AOl5uJ7NfbTzRiPZri477ziRyTXYwwKmk7f
/KL5jlKvndeln/7KDY9NkXGbcWd3pL80x/WXQdSrpbHydLBxSNeUrQlkcr5VeBQi
lhhDzYmdjtDcacVLAyX6C5gcFOn0B87E1PVbnM0WHt6Roiy83NEk/9O6D9TzBMd9
4u1RwS4MHdI9/2EozzAWjZzTEFJy5z8wI6pfZjcGjefuQYBiyGUxceimALmMYPRl
h3dQlpAZyQ9dDmR4y/XiJIigZJiom1mQ/Tbv+OKwcdIdcahHtCVL2AN1pI+P54NM
ofepAlbEbIknTaOxLiVx+gjo63cQ4PrKTEmzhBZWOwE5admrQVSMoLmANyC29kD/
tPY59uit2EDZvqm32b5Yz1MhL0771vwOpAnMcDecGmXveAfAlTBQDm2QTzAkr6jH
nAmxNKtxtUtEKrazCK0EBNbpmE58top+WTKAEHnBJwvlrHs9cIY0CzfxKxhNxLBZ
shKw56rI8T6vyN+l6RX+BhPo7KmR8YsCrVD3tFQ614ZbGXYITquEHilhRPNilWGV
FG3Dz3vD774xV8Jl1wPos6cp0w2W3/vvjxjQsWCNews/kqkH/xQLk8dCvYXueC+G
owm5qJxiQ/1qIrRAEDBSiS3HmYpn6Ab8wEG2+GO6y7yJJZFts6zKX6PdN2YBRI38
L/+fhgAsjhzrKbJFjcGELDHymWsSelw0fAUIKKp+6jvWV9DbfbfbMyfUjM6d/3Jq
j3Yayf3sL2ro9HpL/c+hVfYITSqHew69Sp4kClvIw6MxmEP0MmYDTEUDJa4N88KO
qsJsCNtYcKLbwFGRe3KwQXlq+CpDcoHofjWC8xo3U5iErWLhOkC/9KEl1r1y9xGK
q3dArCllIC5fgbk/4x1TLFKUWbFkSVUGMwsIsC4EU2kvQAziS/9Y9cB800LIILlE
QhlhB1pMPdgg5Gbnfdgasxw1t5zQWQYWQN9ouvue4vq1t7uAqBfEkMSg5979q3TV
IltN3l0UPsmGBOpvpK+j0PZGQbgl/Ov01TY9K2UURbQ58Zs3Bya+sjuL7f8C0PF3
SlQ2fovn9DtkKjnJ9ZxuKs9IflE2+aWYdD4E1fL6IUKmu81NpA4aGVMSgAvzJdem
Bxaq52ciEY0gtO6JfPa15md+i+2rQl2JPd1l8VEVjjF37MAh6am/IqiDVQduqOUF
UR9bjiBLQSp9gvZehgVTcTyrjFxWdW0Hg+Jtthn0Ds6KNvbdiaemm/J6aONZaj1P
xa4iZBk2frsbVV93nwDYHW3we58YRNHFVunv5Jc/0Ud3S8UuPJP9E5dVLoO0iHdb
t5O/+OJSV/r/EeEqDrDzO3sgZVKsNy7dOFfeZEfqsOLGDIFsUblqMq0lm2ziUUyw
Sr6HM0O8CXV95mtOHYPbwv/fz5NQbdMduvC1cxbmePniHIY7rWBcf/BQMdcrppA9
ZqfMEqAJXQCxLBu63w4NeBs8kVbhEsyjTjIRxsTj4ILUZs00kC8y3EaliEeT3j6b
NNMsuqs1nvyRIOwYKBKuc0wBWA9r/BeCIjWVIWzn6wRT7CwuGjbOUMu9Y6DRBzV+
6hAkDwz5GDuhD1hAwruEACKxfX1EQkSL/OnJGFy/A+ci61GvP8ejrye0D7bnag71
m3L8Z/tCkStkI0kFWsHsKeP1Tpw0g/JDxLN4EQiTiFsAZ+EqdnU/hOnsi1axlBp2
Skx38mnbmydGsd1HpbEJ9tcVo7jQw52wINaqmlVCucCFegE9D2+SnpoVyAFu5Vjr
YpRfaxig+AZuZ0rFqmnf0c/Kmiuj0iY0ccT6LD1njod7Ew2VV/8+XzUCApCWlZXx
DE3GBMvIO4eqrZlJQtWy51bJAlaLTaDSPyoR/sm4vDlbjSlcP1AVtVjc1t8L+228
efOiMI/BqOXHYkgUhvPccUiOrgsQ9y0TojKXbITuwu/uD0xdIcs3FT/lxrpJL2w/
P4Rje3MJLjXIutCmNgWaxahNg2zEFxbEmYDMAWQq4ZYHWNPJ2VBgtoMuzBFVQrBY
jbUIH3xcV9URph2WfDwa9OP+1N5tZ9DNyAeSg276o1L1YWeffO4DzQTYfZWZfo++
b1Jhn8arAez3fS3mob2/Lf9eYF4DRzyYcW+g0yZkrGmYBRAEcphnqNqVRd7X7hYQ
fPUwJ4G9hy+I1pBooDeEk1zr+0yiQquU1SxUwZd2aiikCEoC8nsitUMKKDO5/hOM
baNbo8HBJPHIeJXiXoYW+kJvmmUgcDga2kbLxHY8DuxUQjx59magpxNkzv0rYC0+
tptOkj1P7wqi5vOqyKn1+T4WqPJg+0ZK4V4EJY+ocuH0eNs5GlDy8kZb9XzqtK+K
FHFjLNEBKKPY/QbZeVumDNCK5OJymT7SS7n/IZMKLpSVsE/qdIN+KZGnH91Lo0px
bFHyCEnr9eMbnOt9NstZpPH11+yMJ/b3LIe9zlXvMt1jDsgGg+QQkIo+7/dLMZ1E
e9UsTvI6vU6ZxxJTpPNvedX4iZS03XjTJGnLlAAcqR2T3tIV1f8v0yaQn4rfibjj
Tji/EQLh2VJZ8Xm7rggr1GnkkPTspYdm5QxOuyypssNUy4A+D6RES9YBSZpNzSMM
kChDXunrQ9J8tpF0ro+cTwKSzCs33Oobwdkh2AbhNimN7wwVRaad1iob1q1sUurg
+vBKTXgW+/jppvE7xdS6h/QjzEGPuwlqOZn+VDwf1mCV8rGchljnl++uZSLOxhR5
ZnftFqkEfDBR41SDx1eBwnFEn//bmoNoaAn2z7W4FA4JdhZGukCE42WTywv4/D6y
rVm8/k8s9Bu/9T/YVTnSGGBZcbPZl/DCae17pPpCGJ/v/82lc8GYNNNobX8GWXlo
O9M1lHV+hWzduxSJTlJN0FdgB+r59cp3pR++4AqXYz1W3Xt5iEPzisOV9CEyMxkD
2or2i0gQJkgWro5ld5ETTnjA78li2togEF/qJFAUMo4cBpkdw8wLswhPBJ/X8fvd
TQQiUakQhjrfDyvD41nnBzWiAorCDRycvrTzm3XiQAFDDcSE8ulXV/TtCGRtm7BG
tVnBM0o9AK0Thcpq69MsZJ9Wxl1ZiRVNNDQ7wFST6ssSGGcKhB9d8yo61EHRPVIp
YqcgQOXJn/4b+CEC8Mi46pdJcJGD4hCKP9xGk6wJ+5fx/qbyWyehX63s8MYk1xn8
dOzbbp0t3//GphroDwp0GmxD/yLBGNm9M1Ds0g2yLGQRJQtIiLhr3d0yMlGZoqao
9X4SRQqNWPeBwJs5Jb9VHiGRe9i9x5yQouZFYE0r1OhuyuhTXOCmRb1W1+dvB/ug
BY6U85ULCZ1jD61kyb/R0FwbjsxPyYWMPXAlUgj6gKzLmHad92YJrCwhg61W6qZq
9bfGXchdbFio4ox+Bb745CW2xKPkk+yTXMGmlnkf+2+0FMq208jrPEacdsKEzzVS
02L6FRSgsU9yH2Py3S/YyXoMPLMC4oHOIhej0EErNLZnZ2w/tRa5WrMvOKTh/03K
3Wy1JSIVMjak1pDq9CajNoepd0u5sGKExUl154B9aRR66FQYLS/+m9sIiGOfg7pN
j8qsjYGhpS4tH/rKHyKAvhQ+7DpN7JqUi0Oyg9ZVKUVeqhrogOIoZ2tMwk6Y2ku9
y+M12mi53WIB+AMn6jGTRYchv1IuNSZ1TmalMgmMHlza44Wmziuo8C/7IGzOmKMO
D8K0l5Iuk8yA3/Sk0GmqJpl6a9YkjpwbQhlBaU7rQO5Y+16qDb/6v86OPGP4UnfV
8US/dlumSI8SitdXVRlV5aKeUMf5dFWYwNxVRvbdrYOhh9+QJJYCuUIhb2uBeU7U
s/5OAxeJzMti9SZvSyLBNrkA7pYc1X2dIVxgqBgA/NF83E7Xxzh5gwbedRBbiikm
bBwS1hSA+W5w6KKcSaiOPjVv+vd0otbN9/NTEg54h/pBYjc8j9vVgWSo0jdhb8bR
jRtKDF6bfSLK7L4QNQZRpVIcScjOWce3/PVmfhRJmbRQXI7Aw4Ir84PzgljHUVTX
uskvxF+HGTAl0jzLYj/5ofldd12nKbxKW9UuApjFCi5zuudHNY7rh3syCPyHuRfO
ttzYNVkwxHQRiQa8JWf5JcT2qDhDApSoWIZDOiP3szZHMlDqRULWSTr4uGFr7YXy
jlpOm7ZfpPjbJ+FKKCPllCKhzRkVXJ/opWld2HIVKS47ELI5HzN66boyGPf9+rrs
8pkC+OOoLgwV+A+GuW3/8BKk6TVAoF3Wdh4J+fL1TJ1fJRSiFZwtVlQZifgaAebs
hz0RSE92Nxq8vFVdyCV8FPxtKhMxUVWSEyuMEC9baUrT5+mLiDePLITG4/fzyZcF
37ihW5xfR88NbobLbBc4zonjYDrCE103WZZ+FtrIfazSqynsD7+CfjJ+QPEyeiGw
xF6qv9IpUHIrQoqp3/XilbCj/6WrnhRYds0Op2A3JYcR0efAf5f3V93AcsrxpDW0
cdBrPohZPQWDAkQIn1XmMlY+tHuWY3bTx0s+w1/bcQkwsAw6CaxwjBgY/gD/Oa0a
dB+q9DBvDYCyJeyaRnDTY2yih8p2c+cw9+A56obkXkg+SB+XZg//8g26ih8ccLao
B+mk9Za5qcYzHLGWjyS8LzzcVN9C4od+TBRLiBrD+huw68RZ11L5hz/nk3twumZs
ZojWNmBO+yIY5nL+zLH1upC/jUZOdlKkSEeJnQXeiHk00t9+Jqt0q64t3AbzrODe
Myg6L46J+ZiSpRTEBQhb2P7WzQL0PNAuBtX2OtKbew5axuF3yw8jn8k5VzZsXVlR
Tsprdw1Qfd53B8HiRqOd/sCmBOhOI6zFDq/gC7nanOuTftRuNDg25l5Y87NVoJ3c
mfn85GYDuIbHbroN/+wf7t/VmIJKxxV9WNiyUMM377zM3f1avyVnRyRAXu0VOD+P
mBqKHSfGvSoyn8MmlIJAIlzQ4zpbQCk4nEmaA0T+K5aPHYlASOOFJ4m98zWFxirw
F0lHQOTZAIyNVasxQ4M2tFlctUx0mNaPV0jhyLA3CNVELiHpxOg4LD6Q+twp8Iqa
lfp8ZG4mxMm8KUw3/dgLNcx1kMKjlBOHxYZ89AFEOr+FpHP3QZ3a5jzr8ydraz5H
N8QCUERCn3e0hRN5MGvdV1hmD+Ps6RW2WkfzpEfLyNc6DgrMWPKAOYj0IXfv+AaY
NbO98mGZsr4nHjpHQrAO1PY7Hot1CZnxiUTmeDcUNRtlvTPrFk/dN1faR83YXamZ
aluXFXatGfw1LCFk9p/C1/S/9nVsRlHFsAHngB2q7/M56P/rhtbsp3nhpRI91dvY
jPaFN1GJNtSa33AONMX0rDMNZSSU1LWoJ0vx8eMSt0nR8d+xKt1d4alMoe8SeH0W
9sb5avQ9uNLj/ExoCfuYQYp1HO/r/Aosy4W/ADYLDeflYPSheu8uCBehzaoJOVhe
QHG5lwLVS3TA1ssN2Fgy6v5YJkekVh08rD7QvYu0TEUnlHKGAPZAzROxKppseaui
QUWrt6UupgNfeyvLHrUgGazKG1lMbuUqvrbi6wqhiBG0fzM/Fx+L/OYu7Z1hKyM7
/mSOuNyZHj9NYufqt+P0NPM/G7f1trMLgAedOhJKbz2vc7H6Yr2hjbhb+OSHo9Dz
ufcd0RMRNxStsfitFk85YpVONCW1ePy8Q0cOd2CRu0W1L8zEUG02wRy9RK6VDmQm
FBgScRzUy9NRqzBlaqMq2S8F/+4GBqMUNVzxk55il1RIAegjltAnIyFhqKiXN1K2
lFi+ORGN0SoSi2AK/hRhS/0PFk5njZzbuQ/bZOa3ntRVVqfJlSTkgIY6rkD8KZTQ
vwcuHY8mhnsGxWekzs/0+LFZ5yTyDCgzhNyoP2DMqYWoTy2ON84jJzOcbL787SSK
V2qQWeGTxyJZaXG3miRwOLV3AR6Eqq7AgndASBL1EFK+SFtidQ2lQsKYJnSLwcA/
P27Pbx0NwNDNc/cnWqloirAWnwYt1RXPrFkNsdwfUImulbk/pqRXRPxjUhl4bb8j
zzDtcby9heYZ7p1ok8M7AuBAVUIaslyXCjORGE6k0ILVqC3ttwybxyhMh6rQDM6W
5W1sNUK3iPjTpdo2XMm3mRc5M3NnWtmRpEtnuVvWBXcilyrxATUi/YJlPASDmhRH
IYhp99yb3vJ6mFGX9fY/s762+nufpo9zDm2pFCwmAjvISuNovpPWk+sxVGVzYdz7
dyvqiHPCz6wdOEQi0EcIzB7IaES+A9bpTuaJqVlK5w6GzH3tNcG4bpZPVTyAQe9t
B1PFD0cX8OZE3SXX/Jxhbnhue7tXX4lL8DTRUBlM6BKJAOYLk4/+Yfu0EmXe+28W
E4hPRC5dh32wxG6b8fZRsKDa/+2SlQc/51W+cVGQlxXWel1kcPnSDi7DsI5P4Hk8
lGUOuV3Gl3VncKZod3Ltequi0oAFMFfpaCoW+4jxWoMjHBWaRz/XrN2xO6lRWQx5
T20XiLUeCi44MzmkPGS29NQnXdGOtIOpyoW8YXg8q1AOWGTacGn5qV/XuDB/aYRl
O9fISd/M0KpzM8R7hrmQb39CypA67+DeWnIPXEFzufClmPiw6F+iJbJKCL9cPwcM
3DQjdVyTPCT2cUKrHUlMrx91YovfmxFWOevpH8A3Hc3eoTSf+FN6MSrI5bn/+u20
6tIGBmhRUkxHJdQP77b2aAToHQiwmhtQrB/5i8Iil2OJz91ZvYCiVFFu91ftKi2z
GYZNuUUk1X3LdXG/Glk2MBA4RuRY8zw4EYJY1v3ymSJNSedYGc2+uF49PLkiba2e
a9aMC0TJXF4uxIHdZ05l00l9nvHhCR9NB/RVoTwYP63JqdYwnhmwOUGenUgGNH/D
CZef6W7RDb2p0fsu4DjnDqSg2/RZQIkPhszb+HE627s0bNLMONgO4Bw2NAjkd+AX
2ybdcbweA6gAQ3hiGx2NzS/vkbSGJ0+WLPr83tjj8ffcaBJkucJxC+SQPQ2Ex7HL
Mb/pQI0IBQZSQz41GA2RqI/fMIM4oE5V92dKqLBla+U9o95QgJxX+insUUUdQ4Ga
v17i9QI168vcwHDB2McRb1cwHbtjiZffLLYL8+zpXZv2vDAFVwtXIieQ+V6SRVJx
nknDoiEaFlZziPftEQI7llqkA5wszRGDtbNm+3KKf/rb3CSVfdDhBHuxxTneCXGk
7tmCGoA7w6LVKo09S3hlDSZzcy4WnMQwxZNalvG4/WBEuFNT8Q+RR94UrvwJ5w2A
ff6uSB9Y1u7W40C0mb2vEtA/9EcFytdZXH2geqNPwP59CG6spdhGpIqP3Tk8mDHt
V59eJwxyJSs6vk1vUsQAjwlcLIYgFuMM+JN6GlweoKVSmkLgntT6MgfcU1ln07Y0
RwJle+r3zHTLhan/jt+6oNC5Ub2skFVGUA1DzwRX8E8XDXlxvIcDDidmaFDHsPJo
gA+yWLwrAID38feLOKjMDY0lcwo5pQG2yg9qjSGKPjtRQvzadn0pnce8x9SdpQfp
60YLju9JgjDPG72tmdqwx1MWjcaGbNF5AcuTNCrbbH2P9/rWwIH4A/MDFVbu1LjN
bclfbpNpBUUV5Gbb6tywGuYTEOzi/wi/EaQPI3vUGIA2MCcODSji5m9OzcAOP8jm
RXvCNhk7GuQSJYkI6NgsqqMLYLCPHaTkLpCiyxU+814x4Q5j6UdIcgbFk3dL4Q8G
wpdCT0EyJ3RdP1e8YScLQ5dMMTVCG5oujKTqHmtMZELPAPYObxATAhblT4N31DjH
wkMhyi1ugfv9aJ5Rmi1/yC1k9+D82g5fOES2lv+1aVPt2WwmuyX+w9WQTl/3J5dX
bPQzk87/DM0qVXjpUctejcdCNMDnJ+BRhyc4kKtLSLE/bVlx/Zn9aaIbNVKFSpbl
QZ143r8g24BlXjKnpJnwzgJknk2RVXlq9p3S29mGd6Jd3rU1sDrCI3bYDauRkOe/
0/deww67DYelR3tBnb1e7qfTCLjHJuhn1HXN4nUIJuJoSgYVh3II3WMbWY0XtlHB
YoHXNa5eG/bnZUcKzRVFAvjuic9PkMjwEvM2Rga/vWEmaZ6Wim4SM2yf4J1rRPjw
7IRNrf0PLCp4JepEegxawKbRVbuClPDuOj8UjvSBtKPurJBQ9zs21hKAP1/9Rxlo
b1uCAb9nIkpISx4M24RbMoTUaXcwUJXf3aLQOezBeCEddtfDx5orpEsqHRKfam/4
NomCZ6QfI8Z90C7tT8WV9HOD0MP2tZLIpB4ut7AZrheKKvMxrfepJzxskRiY8T9h
KWgRs52vuk88r+YJVylK3kQ6n/WsV7lRZ/u2fIM1iHKrv5HS6dOaTPDE90A/7i0P
p1pRnt8i5POjreA2P6r/LMxD3ZYuvLZ5p+QtL6QAmUJMv2jIMJbgWPBb4l9fGL1l
TBCnSEBiWpIO1rYHuavYOW8M7pP20Ex+Mn35O5z6PeYgJhnBC9U1TPGmUh5sR2BI
WaMN/wkLcIv+Y+QEZO3plXeyQ4/vyaOaqEbpXi96f74Zjd32F2g1cm7ICCifrsIi
oGABSdaTOe1To9wAJYDxYA+P5ExTE3EKAudUkB1IJHzYtVhjwMOIiouaJ4t60fqB
1kUeFptu7QpK/F3ohw5OtyeFQs5qxKhgvNq5QFA0rMRgXsLsO04UjZE3kaZldDLk
wpcFdX1V4OhcTcnGxmN8fdxk9thm8HQtHyxwTKZZFuPbGadZPvlvQ70XvFWKROXZ
oAiFSUxKmQ9RP4GlLXzyng4VFEa88IBWoSWxm71kpF0to/MsqJZmyaiNZNmIsR07
nC4Xp3qgDmaOzFlO/EO52Hv53F5yMO2BWPApRnA1WrEzu52T5xON+bPWWlE1IiVB
8QNuzvFINgVJDhtm2tKdFaogjxXvbQcVI/RFLkmbyWw04QDyiYz0CgrZgpT6aDtr
kuW3LhzZ0i74D8/o0vwIlUyNuTiLZKe6jWczVqk6MBBKI7zi6/L5Vuol4Xgjnp/t
K7GQTt5+X6tL0gYrmlnUfmnrWPPL4hpn7tzg6hCbLFoX1HLTpfiOx0f0zuWf6WCw
IFHhulgzvkRmW722HkKPWnQwsFlY1hfZ6R/8d+lBVTrfa2tdaW/plx/INJFjpubp
eX4OCr20vUFQVVD/0jp4zG3d0NHdQ+0F6DUfrcIWWFA6Gj+GbUlndM1e1+JbnDlS
/+JaLjqy0+CTLtl/BbH//1PmI3ws7NzK5EhDAmd16UXWosYnZN4dPZ9M6Wob8IHK
ixAWGqrvu5wLEgD8HfAliUJuiQv8nLpWlFrhilS1mI+ixo9daiFOopI1JSiVwmYo
M5fJiNt7yTt5egqtOmiOFHmEu3rouc1bXk5+UYryqfc8b+LEMDsGpea6bk5GxqUT
LC+XBqxLrWxRKpJDiMT/uAH5MFCkze1nOApWbXLippEJCSwUKVm2Nnv4gcYHrkbM
ADfciekvhZF5+6LhLRnK2thMWRfgIh5OWA+JOSe+DtKFMjJf73DK0d97qDhtfimM
ljkLdzgNrgiKzfJqu4+B6QMdnifPJbowkD8xwa81TA0zMmkWr7Jw9mXdorsn8Vt6
EFH2qzcu8FgvUnr+n+FnDuAO7zidVqFoqnmVXBb4AHe+UOIAMgEFPDCAuU9vBBVW
fcbeL/uCHuWHE0g4ElIxbSFh5FAxdyyoY+Nyd5dG84k2i3YU4lmLbgSw9jsgKz7o
su55gKLQlIyf8gNlcoh1Nvx1EdoXwCod2SkX53lCn8HvqUUWV2E29VWvFcP1CO+b
mdkDJ9PkRKYQzZ4XNaIsKdUGZBf1g4AdlauG47nuce3PlCa/tvfvib5t0P3QdWL7
qVLjTgmVYZfYAIDojCY4Aw+L+83vElVjp9r9AFoHiHlC1p6pYHz3LylK9abLXCAQ
PcKKFalzJfwmPX4Z4Z/IC7hfSh0YhZvVjiBvqa+e9arqFb4nPTD+Z4B3tT+wyYTN
14Z/8JLUi5HED8PHhDEVKx/zo8+EhUTRhxYHTpnasOlRBGEz+0GJDw+TewG3lp/J
2JOHBsDFB36LhvxCwbciviUWFjHiIYEH5ZIPg7V0qxsE7kqRQUXkkXqoAXxgLhGr
1XwneSlO5up0IJM1m3VlEFMfrkh8Rj9K0t1zcV2lfftj3l9rs+y433e6DBKIWif3
YMkDadQVXziSYZTUz2zFQwDSxxvqFCKbDIPQDWTAKqhR5YMz09lVHGBROUuMBNuX
YpFHABDDkNVY+tI4Z0EMO3cWCM5r9Ek/NaTAljh9HYhXibTlf3BIOI5v8F7lEO7E
E8cs8OgkYxjeWTeNFwncKIynHVNkgv3926lqVVgaS3eXTcIWYnl8ZTRMHdw67h0I
EjvQBXJMsb29BABo/XJbH9oRaf+PzwuH2WX6pG3unG/yju37W6oEtv8ubfA3mYNt
pWSrUEvfk1c7hUfgxsnErhLW447/wdKLXTKEVqJR+SE9ImrW82DDZiWSjvKRZGYv
hvgkBsTETgQh/Mooh5zJLP0OPAHUrc8nsRBXUjtf3D0mnPsARCSoRgcoB59bSaQj
phgbbopMcxh39uQfUVYldmxSOqoOa2KUJCmAgWRJYf2FOxxD3ZXiBufFcDZJBPdA
46errVe2TrftRHc9Lf2li4U2bhS2vbC+5ghLHw9pjQ6crlWkFfqwM29YYj4soZVl
YORrrTE4bfyI7DzZrC5TAuYNUDIFKYJ82zOgqGt+o/TFbFTen9fu3DGhxs1pTPCG
y6fgjpn2GDPh5EbGU0U0gA7/x0sUAEnMo13l3VumdNocKenGl1UiSNrQOk8mBFZL
hDIV9+QklYCWab4SM8rOis1mse2rEygqWuZBnCSSAc3fFB+fl6QI8OZCDbzB1PY6
7Ch2QWA4jKDfDkf7jNmiyqgV8whIo4Z0cksb10kj8gvTrORQsiRRAMnWP73da7aJ
EDZsF7iSFskn9Rk7pK4RmPFkMWhvdKjAjue7+EbpSn28JgzZ8UUqSLK2pUts2dDq
QNnT9CYliLqoMaLLQabOWA7a3Mce4PD9b4p4T9GaMwU7iuEvgREcvD4k9xJydSPn
Mp8p3LviDdwLlbyi0btzn0yckbmBqHNuYMiZfzbVtEgkI76vNZQzOWt3JUwLxD9c
Xl+igE8FBtjSnlU8pYfT57tt1Xehb+O8+QJhatvxq5/d1TNOyK19SXPvUomag8Hi
5FdtEpdPO3vhMgASPva8zZC0X5cZ+qPVCTXNoDHRXgL5Lnt6rZpeVvHutVU3hA1N
cAbd6LnqZseL0C1k91k3Rkctmdh2qfezXGxlX+oI18enVlZ6P6NwUGvLca/RdOxf
iXXM56fS50cd3R205Y3Zu5OKDtNyYPxYAjo+gSv7FzRmEJAjdvbYdvojhPxTHi25
+nq+itHYlpDDYduOWLfgnXNLi13ZB2eP4EWiee2EofBq7gQn1/wNOeCJpgtcoHmS
seIv3/Rd/8x4KMMVv/1g3S71pYQPR6hnQIaCAgWu4SWJZ40Ccfz6pToWBDDxjiKq
6R25yYqQvN1qDAzmPELiM2oncgtkxfXLY/MHnXK5vk6XRGg68er67XO+WFSkoZs9
zul09pBQPN1ip8VNy4k2dsO+1DC0ObhHQQhousuWzcgsxPm4LJLFWe0cNFDv4NBa
PgKBcgRn1qkXEzEQ06DgB+NFLrBk+QBNt6cKhLCBm8KNtneIKRv12d7iUgiy9IoS
gEYbOGG5QUJHl+QQ2V+aGqGip2lZyjfrvdkrjb4jQpyzKoFDqsD3a4osobbV4VF7
Pg2WxEPYoeYoQDtoq+om07iBthyA1MHXgJNDezZmebQpDLOWIC4U2cOn8Lke9f09
WSUOLoXZFBD5v4/YxKAB72a9RQOE2czHxO4D04PCC+hgS4dmYr5DujCWKrJOSSyP
+rvo/mSCLL1gKdrMFa2WyefVAHyeL4LM/Vk4sm9yXtFOWtutLZ+nTfsMeBRNFVSi
mrN7yiI6rqbJfofDqrT+g9BIN6wx93f42OC4LrPcj7muaPkTvUKHiLpVgPbVYcGG
zjF5HZCgmfszZNVT5nGaDtvy/raw25EeVDr8pjsp7bacVUg9y4wHJIXA1K2foEQj
J0Ap0rDDBwZWZgcPQX+RbBr2okO28SoFFvzGUfOVXifpBJeyJb6QHjw4aFWIyVLU
/3BDTdlegX4Oc2rT4ez78qk5XIAwBKgqR3u7xqcWwEVW8F/1aq0lSkX/O7+RJpGT
ySDxIUiTYx+WB2zaiqmkFPYakYNCrZbcHsTquilHItPvRY2Ab1wDfC1jZC5yipFd
SQH15O+m78pLPTDT+nqGYLuhifKMnR41pg+kJxrF6qYhRzcBWo1VVllPJeMYZHI6
2q0NGFjSpAS0yrN8Vx9CmJvIAZcmnmFPis1uSQNdk72Rp6QtvktyGyCa/0f68bZO
uXU4O0S259p9suFuh3aLsLX/eq2nFPIfd0JnWOocMB6zx0CjVTE6Sh9GNNdGKv8r
JbPRQ7udP5YpH3iMop7d5uvoITBV0vuvsrkYhHOmZ+H7C7CnkHIuoHJ8DVWU97HD
ANE/gP/txXBmhgVI6w4HgaSb0TEID7bMG1kKKblOUUQK4q67sD1VdJ0iRZ/I6esk
9QbQUDJwDHhaGHIaYvrx4jHBQdEy1VTncvV3rwXIazWeFHJgJQyS0sP4f9AFouWp
nEy4ENrE1O761HM40UCvsdBs2xZ36EJbbjOoKiRosGRB8BUaEFKFxVHEIgc6/Bdx
DRNC27s5j6gBJmv+qViOBiHeR/8cO3NX/nX6G2mBaliOltlLznpx2DQ1DsJXtZji
e0ZwaopL/M1vA9NsPjsombYd4NKePuxFj6uZVOm18JRd706e0i3cJxSEw02p6Z0L
aIcP0ulkd7sH8c1XE+c7qzX56Wh6C+KqeGjVFQl3fwGT1XjdaNiFJfny9QoPf2K/
A4n8onAfFx5h/WlCE9uVKZ8YLKuXuKXJb1+q2Ixir53lgWQpSq7tQX88aQmg833j
VIvQHGVL77gu7m+E8ZPxWsz6+K0qLytuHAR8GUNhjSYaHDa47XaLuD18it31TkvD
wnFWQwONmgM2eRoiTqPKYiTk+eceGQ/gfFD/9JiW0Ds1Xp+g2cyaNNvtbnjO/x5f
ZLTD1CQLtg5FpDpszVq+mNKeD/coYRrsPAYWd9A1DSQvtCGi4myJ+3HsSBib5IWL
vITWuDypKBTOG7dsxXV++JP0NI81Tnqxhgrs/pFExjwg2xRLtx6i8R+YHdRDsniL
w4S1fMhKZZuUmj3oTcpWYcoyg7EdbC3nkHMUhsjQ5QTkiyqRJBUYGHD88uefW/hZ
8aHl4ACIsy84wmN1tfCZP4oA1wcVMrO/JSxYJDb7G37dX5fZrsNi6dpwCUJP3heZ
BYT4ptWESs5cZwd2YkNOuEiVb536SniJfaeWk/y9p7HA7oPWLh3w8EprHojYxA+w
pSzVblXBOJ0fecta5jI3uZ/PdrTBlYbwt9ueAInhQQ139xURkhtHIYRuMJkuRKZD
Tahafh69KDwV4GNyHhtTsvT8zMLGboIc5bctu/Wn4OnvWV9tkJMlYc538113XbQN
QEUESFUxdi1i+GbskARr50aF3UJHI2kN2D13m6kTvR8cAsOI26a4UBZv2tpg7oGH
PWSIrodHUfcEhkIqZyLcEfd6p1T6U2ysAicd/URffbQxKDd5pdMzj1tUXcbBZ0uP
EsfMOxXfGi2y+ciurqpZAdDPVZs2SfRfmybAeVO72xPPGdMN1SXAFUKyunWeFHvZ
1i0mqwh/8iRuOwYE8Uf5h+uKEJtfrCRFXMbH7WmwIdmQeg/vW0m6f8Pi5Kc/R5Ap
pe/QzG+HTcGYv9HYyik9V1+xxPrzHAzFvEJq4rDnE7z5mhYlnEBft3tej0cbgdUE
lwp+jYq56qrjXlBIexzKjjYkvWllRo5TBHoazkzYBtvLAFzZxXNLMXaKZEa+yp2E
+DwsHJ8RINcS38j/PuNHPHTFfoiPcfHZ38UEnu402nEmG759kusz+rmYtMU8k2nj
omefy96fdnmFPbtwTB5JKy21wqdUsXa0a7CogSCePoS9booIeMKZyOuaP642wjui
cL8JDUBaa8ccAPknxKLc915TaHcgWrmPY/6mZcLeHIMY9LLJi7aCdJdcq4i+yWkT
uTcfXk/63sjEK4533ZMWx9bF3JsyIf4W9w1D5iAu32Xs3vNHbxCKnfSEY9yFMH+w
9At0rLlw+iEK4/mKcS0jIZmXeXM3k93xeb1+87ssZb1vo4PeexA6cYufvE/oMmrG
Kt+EvNwsnkJocFfsWH8eAxl+e1SBsefPgZ23ZOPnlQpXaOBKrL8qe/4XHen1J4IW
3xzR2ihkGMvYoAKUkMH6CWLIDbPG+HvPSzfdlrPfbAZj6m3MPnhPyB0BxeJyVzy+
FCyTgmISFiAVQZSVa34K3v+bu8EZHRdhKX9AqACIZlMVG25ET691iYGXlyoVgeU+
FvH1h/VWId6/Dcht+k+W1pfwFdOAcbCjT6aBW8u0YdnQMKx5KjrXZ8uj4H+R/IkA
tl1IiqkzI08e8CmkuRXhfHfzvkzFqvi515CDWoFVSbyWfJ5J8p7PuWlwD8CYJiP5
4l5TgYNufU3TgohY5DoTIB/8URMZphBeXxnjruzljHajD6fe8UyC8isBNITU7xaQ
Fvbc0aYfYA9y4n2rwTO5tgkn8A0Ma/Y1Y1uPvnVU82m3BV8ZtzJcECcM0F5bdHIJ
bqFxrnfy0aTzoJ6EmVwm/0Yeo3+VttoR26UKGMKnXEdSaLj3mbTtuiGtmerNjuGO
fqpQZ7FVcKneFFmPOrYiL0ZFauV1bviHONvZQonqUFcIyvj3EVr/0v80B5LM0ma/
G8TjSHS7FWJj3L7K1neys5gr5C51GrmRR+qdyJIwkD7iVLkJsCfS7O6pSswAbNr7
tbFA3l+tl1l+WvDdeUFU7k33/UuC2B4ZyOezB6qlPHqyA27U9dF8b94hjqYi9rgB
O4W1BGf4NsDftD/39PMw+kLGpxUGFyTmzSkuSB/wJytXXtiAGEMnuw5pnATUNlvl
eCjk6h9EYa/j1BxgMrMHEovOyQQkNBJzI3njmqZKBdPBApvlkBxvAXizH38sCQcC
oD1Rmqq5tU1EPv2Zw0DFYpWP2J7qlG7+0Cbua2PDaClgbsSPz6PNUDbolACrxUNv
9Vk8fTRE+5JL9v/ReLDYt2s1gnP5RIcb/BfZlZ43hluL3rhroWj8T1F1W8XOOias
O46qlz5K12f/o08o4a0ryDrbbCiSuTLlI45+fV7lQn+SeaiVUu6mtWnBrGV0f6LI
+o53oqBEK6rGpVPRjUGM2HMLObfeUsDaUVCqBMKBrVyDbflC9WuTfYP7KMluNsBF
V7IR1NDyyruVKLo4kd64cZFy7uf8VRxL0BN2nH+6Chi4aPK2fJqvXSuq7m0J7qOD
WBPcAiQVQubuBde0L4Mbze5bXKGFEQXKQJvauRiTbLMNqdmNvmbHeigub3Bw4YLD
i63D50PYoh3+rvef8UawjV+VvEynLXT+2M4y5ExjKaCucyNDncsuI8xBCB/EXZo6
z6uP5Giw22N3iZetTYF/otW/A1p3F0kMdiy5ykp6TkBqbxnuWgHXpkSyQZat+iv8
qcgX+CwAUKJN0Ap6LAXYy7VqsbqxjNnmxXTdj02gZnRYwAkmD4lG0r4ROJZKxLw0
X2OhZ2p9g4lJnnWtzWm6PFnq9G1fk+8ZZ05e8kvgNkpLS9YB8DttkQCjCKm4wA8E
gBxgt3HssONEoU4cu+RsJo9SL3Tb4yb4rfo/1iFrS68WxLH8RwLcJASsE8kbPEZS
FhmelIrtHUD9wfqFoMlg8Rx7PnTz4vFuIBsQfpzIZSp2DFqfRMYFzujW3qvhDm6/
lwm7QOw9JKBcjEsxYbREh7v9G+0t4jelFbBfQFFCKgAUp1wqyGH5CNVJ5cgattZt
K4S2t3Eqh2ByKlFpOQgGpT9agtFpEThCx1Fb5d6JGepyHSn87hB9IlYz6mB+UaCo
E6dJMx9/n5MXhxlYprz2+dHyUByTb1aE4FYz1Xa06S2cRerVlsyDxNbU4+H8ba3Q
ZDh4NLFFATtYCMYaycjZRDEFjSLzwb8288lCyrSpDAVOvjlTasa6PKS62BoS1NDT
33vbC2bn9QqC4BQYiXY2cRWUGLjnkkgM+FCMKbQfBh6AUjSFxNhFEIA5f8481AJW
xT2ZaNnew/0I4bW2HAmaDag2414lx54+z49p4wna2N1ImeCgAuiAmQSaXrBVe3FE
jRLWQkKBEeAp7jvweBtu5gftLZ9HgUMMRm6qIMv4GLdlY6zxPJY5jwS6RW9RRsog
oCz29FkzQUNR/dOtF4ECHk3k05P+B4wuYsW+inizZVe//t7TX7nccIhIv8yVRwn5
Die04dysSLf72wyWH8lFUJLh3n15aSkfQb1LyEhdUGzuwkDMmQDCF86KM+XXQwVA
pX5iJYtpuLNihBeQN5RYhxULfUWPh3RAz5Br59GNBTsc9GOf2sM3D7Af3/VJKkyN
rX0AxwyiZB+MrwX3pox+kw7xcBKhVwf4WRAOKwtGtTQwKRrPHsZMi6jI7yZ/8zGC
+uYbEoCF87iZFl5YR70VUjyZ8VdNuT8m8KOq20l7xkIf6bhEaVmFm5ZvV1ThKRlb
nwaUVbVjijDJdN2/1RzwX+uZkEIEcF0toZsq6/1vtnh4F7Vlg8ZCSoJNkdgvt242
SWJ1p5fpW79OSnt9Yx5rGTx5kpD7h4R/Jh1wZ5trzq6DxcIH8MSO1/bDiTFDsHEa
KJYsNaZQhI1oDWPybnKJFeKNlh9xKBt0TewypUrF1T8lZ/1SGSg4zwZQ+gdCPEF+
ZX+Vxora3+eVBSgpUks4efYhwuax8wzW6oNYwX+eyz8vkQ6jW4HTjQ/iwxyvSp4L
76gCJ24yNgTax5ZFNksSPVyaWqUWcQRr3BjOVmTwA9Y9tFdEP3F3NoYKKZhP+02B
ungEkmo24dHs9HFEqfJ2JpxCF6UIAup+FFyqmsRniS07+HE/eGtlapCLibfRN0bo
9E4DNjLlzICYPBljWwXt0IRKPajuinqZkyUHCB9YPaHNsYKmhMzxbAbTLE8L3zqb
dc447zFWZd/zi4wesMS+kpLMPImSaQR24UT4O4pjH0zv/QAtD8m54UBSZY5mdPb7
JJhMN37Ga0fBNhHSuPwlhasRgnpOibk1HdOLePp5LFdf8/BshFnva21Z7FI23xEr
ArGQGzFfyelA3FN5INuf0UOGw3yo48EEtCUx4Fdai/n6Db9SUOuX75Plcm/u7eSc
xMDslOVcU9aXJriLY/wYe53qdKCM5mjWXeIk12TICKLc+DIirmJtiGTdLdau5pB6
houImBonSIXB6NXJ3zgcBTa3nF0I0M6aFC2Gxc9q3tlBMfNKoUVsbNM7hqlFOe8A
sIrpRh46UPIUmlWT9A7i/8bTjJcTt1OThTfchwaBofs6gIQCXNKK+bCT8t8Ae1LI
7RQ1lcEWj1rsKXRIM/hi8CrBFng5SNQqTT6sXUu8pu2N57HUtWJFCQLfesAuKpsE
8Gtfal7aSlf39+BT46KrcBDuUXf1G1MOiqGAkGk6l4ynvIPfXqUhhDP3XVkAE6i8
93ihIN3N/g+Dmie+a1CyDaFB5YROsNbheO2IMKA7+18vDUPIvfIQldo+syrGv9T4
fF9v+5zX5W3bFk8Lpx6tnmLG4kh0iAtGLe9qtKr7Kf/pXhH79nkmGV8/pBfoOttu
3Mk2R8cH0kkYJt66jD+3OwPzT8MboOpgJn1w4be6v1TOo5W+CO33EExer5YsLYpt
ZKhSxg8pyRQeJvnkrUu4QBGtzzr70zlF5ByIoWx5Dc1DUDgWQe3rX40HaUdEdOtj
FrEkuIR8BKm8diMjVtXpgGH43vZOYz7wI3AT9sk+MiyhlD8uUBj+HoVl/d0nrJsq
CtvJpSXqNvdbUAcNRrWjH+zZaxy2fX7jdeHjRYbBlmnCuXvFU07G2grVuGtRO8xT
T1NTbkOwY9BCip/HVRB22kPKxVeBg73s6jUssHaIwHWbvf4Q12o9p2zp5ccUOfVf
nezB3KFhrO7n+JqgDdcLmc18mEWFAgyKftIbqRG9HIFyaMIMTG75xzOqOs0bcZrA
8+0AymJyLSpcB60e8BnWDapefyhLDbZS8d68yovm3M6+ggWB/xnXQ0GKgCmYUTUd
6vO0PTjSZXE5ChVVYV5nEWxTvEiGL2cA3FhxhzNhYlKOXqDCbvBodN6z7HqXOkBI
MNDDo9FV1wN585IAz8gHhcbHL+/SgjfZiTAybYp6wQKQlhQsKkIHim+c7nrgYCgf
jilx5NbD92rrrtJc8QzDC4YzW0id6OPgT2mStMy6aP3YjuSriBDW2aqEutkuDlBw
7XxpQuC4ZrbJAmo3WJe8RUngD1J7kDaFI4TFojKf+gnF48/2THzlMD1tTMZa3UdM
UkEehUTWimjRV4ZsPAI4f7ISNS+/Oxj9+0cQnKTk/hW7BaYiaZzSDwGNJ5Or78fm
6weEK6Tv2Jw6eLH3uWw4MObv+GAYL2Kjt81VRetc8MHDE4ydzJ0g5e/kkCYle5en
9M/ei7uSenC6XFO51/sRG068Tt7UDVI4CR9+0sibzXUoPfzDZ+MsVROjOkjC4VEf
uv6k1/KRm+RLanq6PuD9JOJ20Ub5BOdxDEL50+joTzSdTlJHYSylxQ+6cz0vb4zF
b28LXJhSJ2PmQyyWQ5Fwzrx/jqtQrZ/VTNeZDFBFh3yJS1IebS5sm6uRkk2Bqh8q
QFD+p3JRkNgZZzx0LmyUqdiSGIJLnAFNmZ/I+5J1VPXpFthuFJUUoriRzEf+xBzH
nBPe+7dkyq/kTJ122kmjKZxOXYb2OYgUy5xnNDpKLUBqfESe2rphASvGlkTBioaq
bB4vsM3GtdwufHOZZjtxpr4Aw/wkoNg3TBWgPBX5YMFcWa+TTPnXRA2LLbzgU2DF
fCEd4pvknC4SIlcIjpiiunsNmfIPCAtBGdOvSZ7ya85YL35OSXq4dghuf3cV/TaQ
KvOMO3OEO1rI1LxIgyIqUrzLEoIElXV0kKBuo2AvMNk5KisKw9E6BvSMPnrYLcuK
1qQ+MB+JJYKtyT/aQN9gqsnnVk92Xw98I+UcgF1Bl7oMEsO9KsfptPXyWKxpOTqD
VxerUPcLg1RgHGtNQ0k83fPvhyGE8WF1PrJxCUqo1BxjKbYUKVmUh0KL1JJd0UD/
gc7pAySyQx7tzgslnjb3YzteJ1eyNIdZ88q2znJtgqYyDln7TOBdSWbVAzDHnaLl
2I/ivki4nqiYjL/sqDDjpyDQpUvTwB/OTzEDZeCo1kyWnERBqp6bcdL6r0giHCEe
VW+35fZ59qnOyyS5m5nzbPoSFNAUISM9o93+tkoL6l+6zAPNH7RECbWeaJRj+ljC
ZuGoAT+1YrjeaYpK8mffeDEas4FQ9ZP+fr6YWAaffZXFDIkH1+jjZKbJUNfe7nzd
J0ekI8/NQJ18fRuFr5dmqHwmNAL7EKufvhZwpgEcwyBpcJlhlSS9FhNWf0XAM+HN
K5j4A6BxdGq44oEfI86g3mCFWJS3T6e8K4QVQs3W5OxA1+ewahczHhfQt85KnxM9
rpHRqWlQGZi4+cqASi7rbHEqxHXQe+eEQNKzscPds0tHuwBQlYTJ32NkSsEWsuoK
lxkA8s/LtC6oNgnccpgxtnTvsA7ZgYO3KMGqm5a7c68rNrWrC9+N8rLRka3+7KXt
QLTQXzSY2yfbyw299prVacP54kGIkExCK/MMQIYI9lqq+dEdAy3qTdzgUirSDasi
oG/afMkV4VpQAev48XZXNZWOd2BcfBOEVdVbKHQukN+9E/BEBKydSzPK2BxY5LrF
LxkNEvOYN8Z0mgDrzbZKt6un/OXsi8Yd+lPMH6Y3KnBtdl38DdvsZTJGQBaohyzm
EEPOylv+zpSpL5N/2nJsP/lHce/Pd5/5r5l5IhxFWAuwqJ+Gnpi4QxFCn6MSnAj8
jZYFNNpYpWCe75ld4yYW58nRSD1C06n7gdMiFwMl9BJqjvOAkSc35+dAibAmAsVk
oa6DFfS2zngR6q1/2oJrwu85YTPYLYU/CDERjfaBUl/7vEbEqYCmff+bB5R277hI
1tUpn7YRRxchAOKPdViJ7Rgf8cbR8JmifnaDs65M5wL+fj5Ki9yvWVkSEMyLw8iM
UGCbVUq9dkyyxXwl14g6adZCMuTtxGSdvODLZt+gWXenjAU5Cg3LbRHNSKCJwsY/
FwiCOh0u2WkhwTtAuqZGErsw46XpOFZq6tYwhscZ+MVJcevNQt8W2QbyyxQXm7p8
0qhEXr0feFuudCFGJv06E0mBU3xZLnAXI/ofLhIPDr+KyLhzIcYX2Hjn6AyVbxPh
oDUo/Xs3o4fQvCByx+BAqdyf3KHfWMA1Qc+73BMOGOaGXVunwvCSOK1lGerahHof
JAcvaO1iLkGKIq/k2cqxA+L1svkBfIBPrjWObEnbKmhyvoOGUSAh4fWyHo2OhZWd
Pkay0pA0mFXDdlnN70g+TCOGYGlWzUsMKSC01I5+zpy8moyzeD3/B5xEGF2408J7
bJn7Xec+5CYN1V46QXVIV2OjRhIiCPG4A/kjSOW819mYZgzo+jr+/7xRmz7wBYDn
B5S9NkTxYo612N1/k6sIQWAB1IFoxCVEmTOgl15xJjrWrax0tGjMvUnHYu0PDRdV
hTBzpzQqvKAOFam+Uvu2RE191hE15o3MDouuMKsntad6OZ9WldJ+Mg/yNK5TJmoM
drUS0wIbqxs9TWvCLc5cqDPDJClFDODpshuvAfXLmDiEoqqFbHycXwFpIFh6+SQe
jkhs/IdtfAbl3TjgxxgE8JGIwMxbiG0O/xOKjDLJN6LpOx0TTVb7bFenKi6h48Q4
tOxeOTh2OdpKjSsB7m4beWOF91APj/GlMGSecilqPwdpN8Ngy03bLrGpw96AT6/e
L4JK8C5Jp6XPC80VjLDJg0qMCWhSLqomI/MtDVACTBPqYMimJDfS0S3hQ6RDXDk0
I7O1FtEaslRlAiXsScIarjCNsR/9nsw6pk3ivxRDr8FjjpTf3Nfa/FIBY2hNcJmu
FSiXYfuaGJUal79NC5VrFMqzvC4Dj9FYJAbldJvzKsAx5FUuVOtU/VWCngJM4fBI
U/uO6gZqjgKE7yiqHv9SmsZXDm1rpM+RVT7UpRcpfTtGJP6I5BYYulQ4lth4qyL8
KKQRZM74GBvUkYz+25FhCUJ/+zmCpCiOXoScLzhKt+49aiffjrHXliIGvxQipo52
C/ytVZh51qJow5ltTax5CWHnXT5TvuXPpYnpf9h5z4OJHYO75eXJmMqWuao5JKVX
C7e3HmJzQWwMmOAMa6T8v4BzyVc4UDwAhGS4yVD5u/sjLAg7xDxEuHa7fGnqbdgp
dQ1+xwEvRq8Q8XKuxcjOTqN6hWqkOuX7/ARqk5ZJO3tyGpn4hsgXlaTrUD0EF8r6
+pFsffnDJGss8bZ6rTbBT1WX+Mmft54MxO+tTACylmteu98RlbB67voArRCpYzbV
Xr4X7eAkBAaX7eHjBVK/bnmeNjSvFeOaIAoCyiCs0tyWkw7sv77kwmAZtMFmlbNI
7wtm6wPwRheM+Uah6a7wzWPCwns0S9JAVDlMtRUoinMZC7o2IFBlxYdDajXh+2gR
AxYvgJg9ai4z15rp4Tdkp7dUaH9uaWNFG8fDm8jITszjx/wA2OYyF5gZhGhR1cRW
PEH3v460dt8JE7lMyu1nhadkdrPuA68tNNe7Irt0ZdG9T4PjreGOMl1LhU21N+fA
pi0X5Ryxe2hmMRukvJGbTFbz8h3a53SJsfNPerb+1M8vmQWk/QAgY473Q8mcgwo4
R6abp2p+mbsehtBD8gPTpFAVDBEn8I2tI1XmrEjcOh3c4ocCU8ROicU4LFbvPb9k
Ppm0kUUG53ymEk67A3Jm3inLnuaoZ3UHsKWwrTNh+oBP/FpEBPIXj03bsvS9SIiC
0xsuD7fTOFCqEC/d8Ab1X/hfao5q1DxdcMyT4jOzxFDfXc0TD7f341rCJK/8gKHZ
XlGS8cx16cZA0KO/gx+M+rbOSYXIsQcMGWFR3iv/1uRugNF6dtXul2j3HfNoY6lm
dNigzndfqdTEO0sTpYlivYp8zctGhmErgP6ZZLVl3hRv0jXwGnNt7f+adxZnNUfQ
ZBH4iIRqKqz3YBeW23e1Zu01ytZBi1faAP+Zp8hGlo3QcxvnN8dbQmhNQfZYjsCQ
fd5s4QS0C7j7Xl/uTiZdwM0QLIQizmtDBVemzrhdoTn/45PVuq69GNvuiY0v58TK
hCAo3cDEm20Fg5ci169NL7FIYKpSqsQW/gnpIx6ZG3WdpsP5h5GubzGSqB15yOqZ
K3Xjlb8nzPhQKSHLPBylspZwzVHZmUkeJZPyUTecpWG+t5FpRPz6mJC+O4hg0cus
jiklDr3gpjNgY3s0ej6WUyt8uTGRGeyhR1DandHtPIwwybCQAA4UIFgSruh02TTB
bqJHkcKZoy0jACElILSzXCBhMapH2Quwaw6nYe7RgXRJYuJpkP1k9GdVcDq5Sdvn
LNMbrDT1LJbMmrkVfVXbHPnbZBRGedp7ObOnKTenhnkcOGR1p8Qg/foxM7g9EDGa
7SiIChUzX2lJv9ANaYa+dAIY6RGkASTqExtcSF3y799ddInm3i8Iewdex29kakUm
Zgx+8feNdCGhJh0soX0INOEW+0DOwqdeLrRKx4EE047Y6FN0LHYlSUJDhfYzMSDE
g3hzjg+fq86Rtlt5NXHXCsUXzRY01bKnOY2hf+vId5x4szoSThzFtg5g074oLgPf
M6B/O2t0U5ZZbN6V9V/pXPXvTdCno62llW4jxfuJr34m2vxC/9WnklVL054dvqV2
yxQXS5956T5YioRks6A3qUJwmXmJ/RO6gXgiTY9kR1E5p/466a3GKWBCc865dk3g
CkEo+74J4lahGmmv+3Ln5EJ6vgWwuoU+RYCen7V6wmKGN8L8oSOLcwz9Y3msDfHV
zovUaDEMp8+Bjysd0y5I2L34neXyC5BnI4V1SV2NMTEzrs8taYMN4ZAPljQGxLNh
/i+WqQL32LADPYNhF5Ah9iIpb2aRZira+GTVyF+nkIMq+N4zc3K9+qJC1geSUBNh
Q3HDu1KcVBwCT8VWB1n6S1nVszjAI+y39c7sfjJRJKQvnhxC254jfWa7rKhQfKoR
pP6bM0osiO8OlHmiJapy7iGEhReM5360o9v03IsxDfDW70yvwwcnOTaUzGP8g5CT
GTDu9cJJqYt6fZAe5RvSToJ7HbX66SjngwdLFUqfYUdo/EU6TWYdV3cGbXwvBs6j
17mQb5BoAg8KLWCcL84mQSHSY3Hjglxl6ZrJl/OPrNtOJnUCJsmt7H/DsSpOTww1
s1HvFzokkI460AgppPdM1TlJ1Rqit+1UC6YzarUqxHfZBBp4Y+FIJESOEYlZOEsx
rTG3yiqDvcuETLE3t9L1AE51G7ozF1nY8U319bq8vkOVCZB+FCr37qmJGBkHhhKQ
nuR++qVBU3ek9hRBR/eEikShpjAe5W3a9ps7R6S9jOiM6y+tTSxSvsOVdMz4Zu9W
YUws7iQDRnpJl6DOUtZI3bRVNKD6njDJDbnMOTU7uZe6oyO0hVf1M+nRdhZ14Wxd
mc+hjmIBWi1DKHZseAFS7xrDelQwWXe4swkQWDyvwjw3C1l8GLz07qXRUGavjglu
0vLVwlmfqVAlh3VNLZ+IWr4WzrULIZDCqGCcH+pzO4d/IWxpoFq6u+o0Tc+TNIfY
6Pfp4H81fQWYN9Rcl5WmGRNuN1i7nDvwCgjrtrvwgGm9876B1Cv1fMfFLmH7LUXP
L6e7YpW5RUz7i9Q5kz+cwhbKzRyibJm8tWcAgFbyw5gUsRCxz4YYpMkfYI9W+xp0
NItKXaS18hWXx9n4mfBVYs47fOVW2JJVny4sbp/6C9fb+AGivJlk6toLIfNgkbJ1
GD8B+1VflLHEMXA63VI8SkDpPEaL2QJNidVNMmZfBDa241l0cPZsTM3mDPYz/K+k
HFMZDdTJ81KhdecIWR+9yx8amsvY9yV38icXHumdAxoPbnbRB/ZyWG4USLd3yZAM
jkb2P4dxp30ZnwQKGBKGxR+5Agli56zD5ZHM1/jITo1HQY5BW2uud70YHVJiD9cl
QkJS0X6z7EWJHDgETfwZBYLaxZNB85eN4O2sxD4ZvhxL1bRbhhXjRnX7GF5jume2
grnqHj5iQaexy2teSxCvjgMXk1R5MzurgNhYRC2UXjt0pHPFmJj33Su9XTLUmR/3
A5Uux0MrMG5WxhMWggZuAa3FSUWfHTSRF52Bng3j11YKMZkwi653FvN8KoZq4lkp
iJB2DmivvIgM/8OC3YrWCl7veSh/o3sPXmvyz5u5X3Fx1TofSl+6/G8Y+UB4blld
e2Xbd8369jIWnCXJ/uOresRAu/OSXd5RtSQwphmwPh8PugXfQ4NAVZxNC9Ps3qeZ
GHj+4WagQJyBhdGKv6rusxm4KdYLfCwA1IUiDG30ukgKycJDsQNOd6RwjDnejmxS
/VoaFsX1ZibOcJdw1yiQjfnlAg8HCZl8Nb+bQjCiuzXAIZLL5uvawWOIUYx6YbYe
MmCAVsbGKCaPKUZpU6GE1zwxq7+gEIBJ5lTA1+bQ0lQv+aTRB7gJqGGTV4WPUuxJ
gEd7x2RhC6p/dxmf51xnzwuo4Dk9C8NJIHqCbR61sLKUBNIac7DfUN8Ah/rg//KN
5m7Ok0BYSZuwG5aYx9fWr3yhd+dzSwKkLLWMSCQoHu7MV8xAm8iZ2CnHKIu3Lqfd
5mENBJhPjgRwn+PPGxvuXi6H1XiS52J9/mwqrlzJd+8+0EqRZOwIenvmzRXBwI4E
GvSq+khB+cyMZCYFVchy0ImtDdY419a8Kca51IG7X7yv90dE8gUa09FyRCEhuATa
0cyTOlbzHufkPcxrIb5bh6ID/qoswCsNJZ9dOsvg5ZacFcKVExDwA+YvGrEY5wBu
WsDOJ2PEsGfi/X+ksUFhpMzg2RC2pv5FV6y0QEjgUlp3GnUXmVUwb88AQkdhZ4tT
sj2yBoFCPWWCRvF079MEB9J1oninDE4ujRKrkomxfjLAsyLP9XBbpkyIEtQkS6nX
o10/OWkfLmqRzkMkjwtVYx/mq24oP794mag6KETtTZeTqDnH6pt9IptDBtWPzP8G
dmAsC2DjKZfnluS3g3Iw+ZvMGW2m2ns7iCWxCq6jikkoch8wuUqiaP9tuXrv1Ra5
7EZn+uTSplEPx9baS3cqJzaruHM3PNMaiiuhVXje2zQdjg8N3SXXWsjVLwPAvDr4
OFgU+YXzZkSA8lHFz/NARy0O755hRshWq8Rq4xl3+a1MGTV1Te4KY+Nl/7kuO9me
6DyIZkCDGjuAyGvK8DbsFwQQTmJr9KnKWrvEowH0ufBRLhpwn5TBHrwxZUu4PRva
RrYUzw7u1Uw+XheKcdJw9Vy3KjlOASn8g0AHuF+nIqJePLkuQ//oMXS6aAPNO0ZY
LMZCWtRvI5xOXrg+IzKycFN5mfAdwL4NH1xBuL9A98fRUQsPhRD/pr3uMJVnz+Fc
VD1xmaMog8Vl8YsL6YP9CWKxZ6B+ajoI2kRq31lkaVvV8nlzgSQqHsn54KHxPcnN
C3bBDNLcFmb+DNoDQ9oq1pzyqHB7hP+Cit30XJCGiZX4sFPy5wwYPuVTvzqnQn0W
FctxV3MtIl10lu1z1Aq0q9dWGcOJd07Xyj1hOCx05PDF4LUAlQ3zxQFvw8SNXFW7
kL6QNgP/avI7uRnD+6yDjl6f9fr0nQKpqHDBqD7rLTHI9wEKUOLwacG3M9vsgrmr
6qW68AoQaBQdmzoYcldBFb+fumh2o7HtUU+LHSOI15th9Cq7xCaeNMwfb6T/KekO
XmEVRCiWQ9x4H1PnjJ+Elor1tR9ltIz2lq/lxRahv1zpw+7E2I8X2zSTfCJFBPQT
8JHCrJu2IWqC0qIF1gJAG55h32dqipg3gcMh2936AItqL7WvgodOu8KTLvdcGBZ3
c1w8qaUsEuNcvtaMxQLBP2tFlJrrrrmW3mXFDSitVYzVm0ULD+BhK50ICnRn+US9
0HxpcLjSqI83K8RtwbG+fjimfGvms7E556f7XhUKUzou9ZJCZjkbXSmPmnyaGjFI
4jriZZhU0RllLgVy0ZFt9zLErJIwVqu6tOXyhYki38qLetmV/d0sC5TrG8e60NAC
B9go1VBFpoIZ+SqzjgCMAKVk6dyds7SWzpgtF9y7eYU/0c268ibjIX2NdihDXPQ6
xnUlhAqs53VkxzpzSyGdbEyt6oSupcIp6AyaIQ+d4XNE901ZJ/vjx3pDn9CBnI3Z
/dDcGerZWHonXn0FKQagxoHW7YIN5tQAs8ZBPTche+lp9NQUH2ex+dh4gJnaXlRk
8NIQQK2UUWeh/U2wpTZ5JguklfYZ4ntHnCFyS2bjFLKm0opNN4ptwuQo2wrNxxhX
EfPVcsz3YLi9Nj8pXy7oO7RcdXREs/TO/r4FXS5nwNwX0TRARtA5InKbs0gOjHBf
FGdGcR2BsAH7P14v8F6558fQCUiOmWmw+UjMLjpD3W2VXvPQuELJcV/NkgwcjS58
jPiZ/MZGHJHap+IUMXVJfNFKGwak1lXaptQxuVHg54jVd2rXTKqvQMHOD/mWHOnZ
JYoaD/3ghwSLylK3kDPY9dnk2pkbkTIxLUpI+ntihU/J11mrvJJ8vOGxyyakVLlE
XCc2mOnMSJytwTRujI7Kv6m4zsV2FiVoU0XsBxxUklrm6aArzCtJR2UtP9zS6rfL
PITVdaYXO8+5uHhXunELqhg0vk4En/R4uZfvkt9cfGr7ksUrk9iW7MllbPw+tTeG
g4ksNvE+hO7Ty3hK8eXIts4HmqqB5DQanjl++hJSk86uptCBMeJCR2vbjpQKlpR1
bS6z0Aqgd+QZbiDX7xuYKHPZRasRwbpyPDR46Gpd/77RoAWMQ2y+/tMoDHTbvyBZ
MDkgXXIhq9DR0ZM21n7lmRKDhz18qvgSZ0u0AH+eaq8KAikMqdGi1f0AWNBwFBMK
zOfvi7UCAnYQ4mBtqNymrhZ5mIC6+5NyPjI5CPezbfGSfzNFWPdwnMVBOsS1D6Uq
Vr3NrB+/6ZHi/+H3h4GmrffSE7avOaIZgec5Htd9oWq0bafrT8fecZgVC/lB91Lj
7o414i8G/t86OkSO1Wmzpf/9rJbeZ+mowJ7/RrGz6xm1FLssJ6JSUx1VUta6HD28
seNL+JQmTjrrVJH3zMUx9aR+apHGFyNsgpHoqBiMsME+s/dbq96tje7IHfMjM7nL
4p1ysgcgC5PZdQmiAqjS+8CVEg5Qx7Zxdnc3jlA1/7WwhZxlbL6r3KtYR2T8KGSr
MoxjQEmGhF+nmF8rxRxFPS1GTGdMqqPTelwLMaWPHqXLwM++qChe1GIWqm0f6ErS
GPkG7m1aT+7Hyf9yIKoCbM6/p0NYHNG1ek0VA8euaLbZfZRVJA8MwcU/3bpK7x/2
iDXpFz3REzcgPCaVMpx0bEhoEvjHd8aXY88AMB24rg3lK3h+l+ixe5GZ1Pf5JfEB
M6yQ04UR44N49uEyH8W5UzARvavRXBYwUrS14WgeWXIIw/wDUCZuUSrUwc56INGO
8lggLtwEFPSvfTReaED5SJVctiYr+08xoQ9eSLGNuIb97EuxFXDy1bKZpq5Mkbq7
soc7RnGxFlsl+M65/69vCVB2CrX24LjVqnbRNKLgrvnIXUQDEpdU4AoyxpfIRo4P
blGGhOc0Ix8XfVc4Y+bL8SPKNDGsz4xCWKLQ7YG2MWm/5BgHhDHM2Ox9qyTpTVt7
wqK8dYcw6hg3Lfvo2whq2qAGM3KiVTEXnfxF4G3BmIZhNLjP+WB64J6za/7h67x4
2XgjxgcNFh4TiMhDsJqon7lTJVGEaYX1xVZVLxdqhxCUr9w2lE9rE/iMcDEFoMls
qudGWb2i31hSlNQhsziEAdL1ycOkO8Ia61lLSPSMcDo79TIJUGmoxYzXx7VxCycf
rb4+FsOYglyNAev4s0ThAT5RzQAkWzvTBWDg4tNxknTDv+d/v4pVFRreNFvVKqHj
WQy7PcXve8pcUV4AZnyZTsybf9HgnzKwavOpnXQdZTBOcI6D5zeCNDXmvRXp2rgX
52Xp4XlkpMQnUXVxcBABjmoehyfCjX1OI+a2JJCuSv0376pP2F8774kMhA+LlvbA
I5hAsuBuFFRtf47S5JzO+5gTInh0XiXWGRgtiAzW682mdBU3LSbgW3/VSKEk/tiI
pNXWn1+PT2Pt0Um8ewrHkYf8M5mNnaQfFs6NID7gZxDuP+FUNLWkdlZFY38JpS5k
TFJC1xSAgBwkCw/6jW8X8wSWAMLVMqEPhcbrykHKFmC06UxXsqik7PPPadyHpAGZ
S31EKbDx1Ad08hd9wCi0rMq3juDg+FoZluI99jowVXr02fkE5vjTKWyWQTFVR6xp
LxmluGg83+pcU8v3md+jkq2LHwnAX2CgSnWqp2xwDRJvDLdvNBH6UMTcYQ9kGLr/
oOzJGTvnswiY9aC+UKybMzClRaUcmOnGxJLyU1o+108L/+DXIKHyzMI1+LMaRihB
fvqdpxGrFnTi3AV3pnmz3w==
`protect END_PROTECTED
