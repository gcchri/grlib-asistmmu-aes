`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
khjFXSZIPapBDyk6Tb0YadGWD86gn7O3j3NX2qLksl/KX4i0U7Gf2P7iLAYIqO8q
4K20djmtsO33SDpYOTuUfe5AtRgv0BTbLJWEnWcR2SYi4aWVllvtmzB6TMObCM7F
pgldRwum15WJHw57Y344XdWqVcO1x83W3DaBEduxbaxMhnkX2V4zM6WXE5ZqTKRX
kEDifvtXbkwrY8dbudYVdHXaaVkge5QM0x3AAjocmLy5XmzJnNClHtT5ly8VB7UO
bFdaKlHY+eKuNmjYCkPqa9gxbEry2vOc4WyPOyonF0pegAvlaBKg7nTgPtd0zYS/
s6XO+8VtwMmQr2VvHDxZfk//RQDFnltMal6K33oF0IV3fwrqfKR1kDZdlwJOq4rK
`protect END_PROTECTED
