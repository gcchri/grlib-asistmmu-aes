`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zxnA/YPbqMH+rhaXiVxM8v/YjEJlaO8xt2/daL65pkfwqsYkeBlSJBlDL/bAKr50
F6A8RIC+rfn5nwsPNI/zzISCtmP7MosgwcsJd0LMBi3vLo3gvMZA8X5LqSkaVodZ
IAC386gcdq1OlKuY9PLxE1wWmtPCzFLdf1ZZW1lxs9yhzymdR8IIVng34hqnBFej
Wr2Nb/pcuL7AdsbN4ZKH8yLnil4yoIjd4DoZ4hWARWmqKew7o8f+uppxoqhb+ouM
f0cT8MUAMsVTbJWuicOu2McYQWL/fO5VO0cRnF3ohztHkqa46FdBFWJk59V1fS2o
vUQR2qaqzTRa9+nkW7XlAlOf+TLfspWFVfRuyfo+k4XR+KK+oXMYKvwMwtLnQMe4
jEDoDmN6BCEb5qQKPu/qdz5yZRuBEV3a5tJnTSj5cB12sv1iHe3+oUkdL+/l5aIn
nZ5Q/o6IH/4jMtIfY6OCqu802vVWywl1FDrMJcxcpveIfqnjJux2FbEC9UfftLbx
`protect END_PROTECTED
