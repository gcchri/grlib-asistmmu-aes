`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VFsaxXTxC2dzpOy9sTtHl9pebcdMrRHKYfNWSwMOgUa6fTM+rB/EMih5YElHY2CR
Vet+9jfXxPb0SMGqp7tOfhXS483ZkkJkFsbALCdTtPnTcQqYU++gqTndNLvyCrXb
1d177fZRVTcX1P5aD712xo5wzkG64WqQMgXg/HDLaMnE/Z8LsHp5cUdMy29OmXHZ
E5jyrJPK3jUSJW1p655gz46Up74zTkHrp9aLlAQKPKNmlakl/UAheOiv/gLlfKit
NdQtlv9rVNfbSR9/zSRZi7cllt/9f2zf2pCAL6Ah6UOswlYzYtklh+k9gjCt1RCB
GY3NjIG+DQV5RzTH0LzHQo1OX6V49W/xkR43H4XfhKs8/yFJndGOkemsy81+HeB+
GZ/Z1icRsqQP9GTwAXx6d1SGHylGPatk/Ie3tWQoJ85NHe+OGDoQkBTwNHuqgsr2
`protect END_PROTECTED
