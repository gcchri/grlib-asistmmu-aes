`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fD1X0bDb/MqrpykPCsOUHeCL5MSTUWV7mCP1Do6yIMT4SxnfWC6oKnVwkOZNqXXV
7LO2FeKOqhsXLDWxnyVZz1PVHLGvozvCdOIe9Yodze+N4dtICEoRCbhQdB8t8U76
2hLc+F6fpMetpTPHrMjgjIifrowxBMeichjIJd1oPtzYzaQp3NSrR+Q2Y5+oUHHy
M1+bWMJTK8mV7fLFj1H2nLEMh2eY/LcMlOEW2rmK1dBvtp0Uk63B6vRklk7Nucug
idUgBlB16FtgNtZFo+fhhDMWmAEZUiN03bqStAIeTEnbNHHSriJ92cZi7OyhDKq/
+1jicqETp9C7kM5We9GjEjr+X+8rs0Yaafrxpfi6JoUiBJio+TEd9ox7bSHDz8GM
B5MTqczgPTld1pEOPjqR7/VXSO1X24U5/C2458/yMbBOmgQ2yL7+06bO2RT31kzJ
APXVDoI0q6PvWYIR+t41WuDklV08kw6C7NPsmpYDPEngMQcQIf6sREvKnSWFixZ8
gVJLTAAa/FIB2Cko6lGTSEEne5fd2iE7Ge8o9T2Ps1j2epWzuNWu/carnj/YMxHa
`protect END_PROTECTED
