`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TLuPw0fououfr1JEGiSxmip4HJge8tr2R4I7p14iUEM5h2LJnu6lKM/jbDxunSSV
JWwrir2VOQz3PtPj6bF+J6k8qkprwObATtg+VpoKVHonFYKx1a0s0fzokKQbbmn+
2t7vUGOH2Rgn7EejH+LUpelF6mqO3DV8zB3D2TY4PAHCC9eeq1kQ8Pv/zwLDSIDi
2WVmu9NsXlKwf44NEg7ghFtN3dorcIYTnk9io8kOxZMpEvLrk3zPkKNztvL2MxUL
ti9u+kaCwSqniJNviX57i7JaPpFsLVCjvqXtb2CE/GAVXU/wPAz14RjOXFHvB2ho
`protect END_PROTECTED
