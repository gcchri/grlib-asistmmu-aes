`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wrSgDMo/ZUONN9JOQxnRaoc/OmUhW5O/hiax2gl0z0X7egc2F6vTnb9/SMxmSYVR
dhvkl4nS3FhOIV03oOdo+HYa8nHGehB2MaamzRa6ubmonBVa0TWEFcr+TbC7qNto
3G6k493zylLLJDRghIm5d1pLh+0BP0hGHbhraJX3/xpJNC7TLbJi8HGb2+TFHy9B
lQauMkJzh4FZ5XM+BiN0XjP4eN9bTBfoU+Vx+mBTLQ13t8XGXO8oS1Pyn1xWjgRP
hA3uxznFg8U8LNDGlCQLFjthP2vyd+LyRlSzF5tWttlriU6DIkLbgcw9GZMMX4eN
gj3C4Gt3YTHmPGQGW911JfcqIhPsYKJDIAgdZAvgLPw64NcJpXvLHBl86AMr4E+L
GCwbsH2o6B03rgV5lR5SCp/Xn/Q4tZHrEzZxZ+SN2YWvwGMEtMcxYmWSiJzeb9yl
NbO7GIheOmxxycvsI5RK7dV08vLDHaMSl3FiNdv/aTIaNfJNc0ZagG8IZ8lY8HXe
3TF5XFRJKhAwyEU5zqJlCmgRla/JbjPni504zoGacYSoEXT93xQIMOCH4k9kQiw2
RJmkHOtSQfI+LgwJdXvlTKmkXd/z4RTVRqgUYUMrDfPjVwkmvsoZ1h747OjTuNDu
nE91KQ0zp0XuoBTnYD5SP9S7MMFkP0QrKgE646VKF08jPZg7Pa5ZyBrJepFdtLee
AC2qbsI/sROvnaULlcEmb7BJbRkQCnLgU0c25anxOH8J4y72h+Fo/0q66WVOZvdw
E5qJChxfkQEJuae06+4deX7WL9Ubqbn+GYJoKjrGECvFZosgo2mmwFt2n7hIE1TP
DRy13r6fX4KSYY7Fta+S1f1hTKowfn7yiQ0UdtHhcp2psdS7KyNVMxPrztLXx1PP
gOs1EzEpLHTH2qEvjCIbvm+JxtfLZAWvh5dilRKbGoDxvgWsGzbLBM6qgmU4cTGF
2/pJ9tGWWhpYuo5uM0SSAPWIFli9UpFzLx7qgkQ59a1O/uR3dM0dSuVfjsdKs9gy
+mouO4AJbwq1IkJWxel4Qz2GmT0XdVZyynbMyyxA9EFtYWwFnsSjL+9ob3Z4yhNE
ZiQ8Q8QpHXlWGjskqmQp1XLkVTGXEFwSv4Js/uH87CMz2iI4oq6QifPwS4b5vX7t
1h91LqgF9ZJ/LZRE9Qi9bBn/ZpnUSYx0vEa1xTNXyB+p5xfEQblwo7U4giDbMnI5
ioEsbQcEfwgNu1aMrQc3oaNOZZTEpdvbhhkU1sG/5iAVv1KvHiWb5cSMZPX6Tz69
qTCPYWlT/BJ+1kXhZ9kwVp1sDEaKrhkqY30b9NE5g57R/ZWoXUoE8psBV1Wben8i
fgnkijWx3wZNIahQ/h0N1U/FzeNoqcHmSYJrXapV0QMhxIgdGJhSWbrfiAFJ8+2y
EYzhMf+2akSvSau+LSXVE5AgV5Dj+VaYW5ToSnlGqotKKVnqAaglK23Xl9nIzSMw
FCMVt70zCV3R83Z09a012W6kyokA9U2K07esZkInxRRpyL9XRQSvSvVlNOcqsCYb
BugYV/Ku/VYJ2fLHEV1wicVeU2r12jjPKtl1U2z3AQUBy3FZYCCxcScIJ+cXi8HD
gdFPoYfixQeNSlvPgLKtUyal9Do/f8ISI5/x48znD1NFy2lw11acpH1Bhw0DeM7w
0Eou/o+B97R5sfpSl4Np9q5cSJGbCyA3RRHuljGVOOlSzlBC30OWk4ZCdSp/o7EZ
DLpux0tGqkrM6gKH1fpvA899+FDrhdb+SXnGE6ZVISNiFnEn+IJ4wvKZcD9Y5f0R
vv9LO+/lBF2DBleHRdZ1Nx7DtAqib1Z1/43S/1sZZLqDrCEEzvoS+d2OIo4MUhts
KNN8E+zFtW1vRDkbUCMCZo7sceszJ7ar08sfZfSSkyy5sjUTw5i+i0FQ+EkHaMtk
T9yItd7waFeB5r3Ch8uaJnUq6qqAbGNQkIFTDlf9xLYNQPHWMFZfhJhbwLv5YJUB
xzHETKqVGr470PN+IiGimyPJuvBNHW5lojJt86SAqX1Wwhty76K/HfSKjuPXZnGB
HO3WJpCiFb/M77jnpnZRS8Y7vE+GagC5SBTdOzYZdXBUceVMPx8KlI69YcQuWPWE
G/bfM0XG2BEgmdAgzMY+5SbERKomtcjkEKjmoq3T17zt5mHxh6dM0wAL8iskIcyM
yw73EvYU15CNgvE2aaBCxqgxzQbwcpha9S7bvnI32tJ7NGSO+dDcr8ncw/B9u9wH
uEhEx9AoloFaA93OPFNekW9imSMm4EUe2LzDqiNX8ClobR6jQPH+s5iLAQ5jBzVL
T7+7pE4s0ic6NSuLrP+SGfWWFjcXhl8Fn7sCA4Bx+rgNFE+IVr5QrD5VZb3G7Zj8
7T9P4MUNF6to7e9AFqR29FodQOpzQfzyXuJznqt2E/QJj2lqiaS1ZK26iHEF7JGO
8crK9zK3VU9z5KmNm7ZaH/z4ERMT1FTzhr49VBVsXodlQZupbJV29igcbTYcoQ9u
8UqFCWWprSqoi+G6dbX5iC1WY890wZlgnptFgLYrO3rjOR4D/8CKGQWcMa905Dtl
9/elHyM10rKOHBi/duQpZ/oPPiiiyg0BGtaB+8VHni4J5BEzc0F14Lkksi9PEXt+
EXItqYzMnOZoncDOEOM582MlhJmkhCzNd/a7brfVzEz7vYcy/+O7y5KrG+qOTwgJ
4QrJ5XRRA0MaBII++zAxPFOz4MJcpxsHXUWoIYyoAYFtXYlMozJb4JGMQjJuinLF
Xerv3dNqWfpf3Rcvz5zQpo7kPPHeibfiFJl5wNiFjn7bDnTsC7lMHKs88fOSmjcj
rWl7a48wfsyg0SOnFUmFk9iT2HAjG+SUGnJ85+oM3c22VD6CYm+p2fHcUYp8MwdW
oxvy/9jtx3NvbPzv2L7MXmcrrnmG/Yy85g8W2oEWw9hznpW+PEvwCNppkx1+aHH+
sBSL0s2xaCeTuBaicDTpIeuayJWdQuWaUzHw0nnVRJbK8ob/0EDlN58+s09+HhRR
wncQMXk8Sr0YmIS7Y86lVbNJAxFjiHG752NLrrXTEt4rxmgOEFCGNg6RCpSpMrfy
l3NGQ/HGfIyhWQWoi52/wI55Vmf0wK5lB2qmOSrcKVLSFVaGASeYkWpzDi0VUWtH
ovwaeGorKCGYhKl/IKgTSRoSkJTxRCAzjdBIgC3jTkiyVWEdiX8htLkdypxifbH8
KYBnIHk9VPVPFpX0aFJcOziSTD0DEatiUhyVRgm1gbvH/wwZOIvKNjs02T52z0Lp
MzEL7vECAxOrBMnY8WJgCNqzw9FRMH4zOt9e7FtVv2HYEgJbUnzyNjFuyOee6iRc
dPhTpmvhAwAk7+bkHjeu/l/kaADOTXG/aI0KU7NQOooVuVb7lyywi88sntuTleAC
sg3ULQN0SeoNOUD5lT8GV2r7bq71Nxj6PjiiocJWje4oVJvlr1FcXPe7Kg/m3hbh
h6PwzITFR572vDUiC2iDv8fW3SvclVIQyE4uEef5hMU=
`protect END_PROTECTED
