`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
seOWD13ROL5/VkUbhBbvShhAJEwOlY9hEjerkJ3V+vcvWaDcuXrXEvu+oXg4DaAR
J5W1wXo/7fuGBOz3uhhhFxt/8aXmlyqIEXOHlf0R24mM7YRXIKscfFxEbZ3z93p5
KcOiLHtFTqEi41DB+STX4bh7suF63BWsqHWUqfg3e8grpCwK7OvFtSER8HQy4uEx
kzRl5WUgne1r80tHMfndSXyr1npVOZDnG9n+mLPbwlQ4KWnZcVWPK/ylPpj0+NaA
swbIco6KrDdaBgng+n4/pGLGWI65/ItYa5C+x0m0LySbuyH0y0StqBlIyfUz4Vrw
uhKBpoYV227lW5Q4JIwroHbWBArNYQ3TrXCoCJ2N3OIO/z118JduoVlw+GsFhGEM
mrLE6LslnRvAqGk5JzOCBBYYeuO/Rf94k8mDiDZWbSjMjh1vhRofFRqFzhoGvjgZ
lrm6MdTt5++hn8flmMYyQfqJsgde8NrzmHAqmo+lDZ59pEQieSkvaDP1mLmgT23u
s6BHrybH+1rM2yb2VDgGAT/ISVsoSk9hF4b1WHuHn/Do9pj+fZSfbQaA5vnDhZUG
ztXMFOw6xMgQskE5uWQeqHBQllasCHftlNj7wG0W5HiSU9v1rFVM+y+UVZnJ8a3T
xxVTvgTajDNI3PKop6Zc7u0lj/TFSN2Llt6klbjSM3nuWv56jxmvy6uzttNw8Yx+
YBrz9Mt9CKQvHQL184sJj2WvZhNvKqHSrcI6/hKbrxC60+8ufIIAL2X3jE2AA2EB
`protect END_PROTECTED
