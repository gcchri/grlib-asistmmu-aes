`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
isA3Zu51o7P4FikdTFAmvDLd/Jk2kWG3rIolR9oDnHhEHXEo2E+8ENPvfDa80lSd
Rndg+v7ozLayj3nA89xSHqY+2QZXAGP7qtdC6KDj6feZ5735S3zyS0vVDElvEjTX
lR+I8SK1gKf46JhzcvIZHVKkiDNnPoCiZdO/9c4rTjs7+IDSt2iQs+qYuNCh6mAc
ELmc13poj2Sa7PkWiJDgnniWM8KzgTzOsBP5nMVv9gJ1J2YdGfRqWUOMWGSmBxR/
Hkv4qLlqm437yo7k+8lVEue5U7wQwEfhmUXrmWBKz0y1ySz/CwktNijma2QdXmr6
Aaf+DDhd+s1+zwGtTHb+gg==
`protect END_PROTECTED
