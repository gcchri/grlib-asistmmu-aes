`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WCDg0RZ92R+uW22bqFw7ISA/9ZqzNPi0HZPNaSPSoDT4lcGfDms5DjZBdkJnY+vw
jbqAvStifuITKQWKxRm1eZyzx4ZQHnc728tFs3ZvqiwGFpCnVEsJ1kk+7LcnH8O7
B1f6qNiFlsHNyCCH1iAY1FC+d00TnzmvgPBpxrngOphOYu6WVf0j4tH9FEybdizn
NhCInymaEGq7R3CNoCzzY1AdyKXrhB24UMSo5AsmyCaC6Z2Qc8wwgu7RVpirIm/z
VBqxBE8tX7TLngBArAsR3BvXPY6AgHZWwyfled/O0YLFIlJoGKHt5BvZG6lyIvTY
w/xTw6NseQL574gdltDdmA==
`protect END_PROTECTED
