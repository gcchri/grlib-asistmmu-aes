`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RgQrkOsg1nqCmAb5bNcz9wBebrIasKS87XHSbgpis/LArJlwif5gAE/TXnxZOpt8
zjYLeCYjwd5mPaRkVX1Yj6rNzu66VZ+6JVloL9kqOK5b2BMBZ+E4d5abqj1Ryi2a
fPAWtoxoUfuM+z4hr7mKc8AlaVC36IooqPJfuLD1ac+hAtmDsFe1Bdf9EeroNjGf
PGK5QpqDwBRahvycvNCC9lv/0QqC4qdy8ZUWzd6vnUY1x8nW6YmI9Bk+yoINhfRb
+os2H5ixR8I7gk6V0J1TKxnSbVb+v8dINg88XAcqqf0hp8js62gS0XbYq+lx4Mwk
QbYBG1pFsefPeJTzvzUapsNg1bFjdRWqzJjsSitKXALahoD5VduMxBKl7sYGirxu
/HMNj5ofZDX3KRc7zFGb0mD2mEyicuYNBN16g29TAFtDMDqwBcq7ODp7E+gg1ftV
n0bKPaOyrD9mNr42qR+fLjcow1dyvvTqHiRqXAedx/uaAEONmtO3VVUdyKAIhMZX
8kORHpSKl63F0zhm/0N11Q19qQ0XVugmhIahzeAFVV8PSBZko2bkXA53o9Feiogj
CPiNKxmwxVrDpXqBYe551A==
`protect END_PROTECTED
