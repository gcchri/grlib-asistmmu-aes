`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kliQidYzWMNl41wxw3ShbkclylG2iTjP1S4Ald1Q5ex7GxHQ1gntZa0P8bpoFVFH
dLE6d4T0mj8vDvaF4dFik1Lik8iVJjlEc/8l5VUjkuDUwWnZPLVwB03pD/Kf20vE
65PkF5jt7xcqN6aviWb5hTygLnqa4TIrhG0gN8VCMwSLVvzfRV7AMmkKl7pP/AaY
TawOeKT6vYxGQlJWVBRpbMuRmgGzSyYxV2rxPL4fg4wN7uvhd0tc2uLAxstuTW32
wnVBmBqRhHgHXmsTY7a9JbUNGRQeZ/7C/VcwL0cMLThQeUtPPVlqYlCS0Z4shfyp
C4qzc+Je/yHPKWHMssr6dZlnwTCpEd5GMCsn2OnRLSSjLSZRfcvA9VmTwZTgxutv
JEv0uckVT+sqMOv38q0aZ271XX7Vdy3LteiszHOFVa/jAf57S71BkX66lyLSa2CJ
jq1tvTEA6hLQhzXyvyWIrwhDBibJC5WJWPVEvGt1KRcwCcecWsqNnRebB1LT7CiR
gvsu7hte3weQx6iiu2sB7qjoaRAQXJWrXuWMWyC89M/gTBxGvMxkERTX9zGmffzP
7n29lXmNha06z4b8HgV+s3nW+rUrfxAYR9Qe8ZBAdsOwN3zo95fHXrBBSwK7dBlF
xFlw2snYZH80Ki0z3qKJ/KOmgu1IC0itSP4gJIYugprzj8OFLdd6dUYBvsi4SrTi
lCBE8nt6o4sUaI3Vlp+uMc7xJHd740vA1R1tfkZVotCOebpM6XaX5zXvi9S8T/5w
QlbQF5kJzcipTgMKmR+JJNCLWhDaIWuoTF5gIdApbSgL6v0XuOf0hbM1BCgLUAF8
qIky1hrc9uIIBoeeCOedjj3kXHFc33CxfqOA3yK6W+O12HvBoV4a3DwyFCm1/19F
0AwWhUFqsa4AjaBQuBmRN1POE/iSASKuA/1mrayl/lnhn+nd131qIAdAF+vbAb9E
K16f/1/5IM3KBfw9WuCESm0UtT7t3o8bDsNG/ziloWtBjHEl1inDXCgDQSbTz0sS
XHPc0cUeKfswYYFnBBBXz96mRyffeFgTkO723AdUD8yhXe2GTr1QdNCmyX3U+Bop
V7jAZeFFew1VI3mRt47gLREVJCtwbyrxt91FJN/FVDHC/VKa87IJABMSs/2kIw0p
QnxwhnYCxjQa7FkMbY1DoejZoXY9l824FK0CbYIePKHokVWgIhe35BfmnXbbJGqO
lZb3QeeSqSIuL5DEi0XukS2hVbMPz4VdvVeE44T2EYRg3CdpwTdpeeadqJK7dQWK
UcbSHG8Azq0pV1323RE0aIhJmpPOYA4bYN9x9Qdm3rBrX+IvOh3fl0MA58l3RTrM
f/K7dtSTXKkdiuRujr5cv2gLSoKST9RTTmBo5L6sqXV2A/bvl/RMw2sjUfTmUHKZ
e4FIPfid901MkWbMaHTPXyujAc71dpvc5O8glaN8UFjlHvbicZ15aSaXYKl3CUFG
H5lf+clp1A5lR8LR7dpOmQQfzqdGnKh+pnaLQukjnhCR9o3yBd5crJnOkmeoeg2S
/F17km2911EdrqPNhmvnDpfwVdT7vkHbHUZuVCQxri4bkEXbFOoSDW16gi/mmaHU
fhQl23Pjki1RfDsqfhg4mfY+km5XMI8mHZ5YLORKytOhYVOl98i3EoyfTBr48+2P
ALKmD4ALtM0VhM+/y0inBcUyzWw8Ro+OSISjUTaT6mShEwiCKauzlviNo00xXxBz
BxkxX1rLj6VMVgPE82kUVJROo8P3xi404dOR1YL8GR9NJsxQa8NrEiMP0Y7zhjy7
dE0bvnLF5sC2uzPoQc3skiCQxQehTx8jp1gHeCfOoXJoZu3OT/S1Osdsm7TPExiC
9bNMGWGO9tPUsKU2QnlYIqUq1oUJpZ37Jz0Z7t622kLqosNEMrMj3WSERpvn5X8B
udC70S+6ZI6lrR+YC1aP+fb+uUT3VQ3i1sZgwETO1lNGxwpDBiKvyygXYlxXr/uV
POx13Zgt/kGThxwqR/9edn93j8BttCE5VqHtuinv/E5iP6X0RJDtFNguePFiMHfJ
0y6YjQNSLr8Lt4rqFJcX6MWQdMunO2zi6QYOVY1NbO1zNxVzwg2kFawKB04JDAs4
AMnM7BMso+eqCpJkZHpYVS0BSlrUrrsxT75wel7hTS/FeWPeBtqLH2AtLjqx5ZWf
MK3hEkS1+z7nMmql00fL5UwKLy0npLi0V+ZCgWlBViA2sgztoYuyNgRRc7oEhIhD
kTO1Y3QDSbGVUrB7ANA8qmfjypm51umMxN63y3XE9cXjZI9kcsNZzgXWfu7I0Oo0
FCVgPiMOwPUO1cYj85OfNXL+m9b2juuJ8YOqHTSvCDKetp7xu0P5ypknAczNzMg6
WIPrvCd4KN351W+VD9+hWdnUeiGfGi14ixucY2zWXBFoFnlCsnzvahvsMb+YLpjp
jP3V3+MVYej368VGv2kJ5zoIdP+enJA6GA1higGS/X0OfMGk/4H0pHQ/rYwoHfhV
BBt0YOp2LB5wkTZN39W+4HA7pbByAOvvgtd/rvjrIOmLkWNyiENGTLbaX4eobv4T
TdkRziH/BQp3pbABhfyLDbj1Otj7albXwS7YP9FMHIuXkuF8mtzgRB5s2yHXUjLp
UakTd65bwPUmXE5WxbSz9RUgWE78eadmudPjFL7Q7hIgkx/UcRvfH/ba+rQO/GUP
85qpvrENyEp9Lnt3SA5HoIYTH12C5jfzXZ7UYJl0pwKe7hdfavk3n2rBJGVZ2INk
kGOOa3v1vWO6+OCxO300adEXqPjSDmec10K+CcMm/dH+e6KtMDtTbGSZX62v1eub
qeGuuyRUEvDoBUpm8funku5Tza1Ls57AAQlrzOsXWlOXPF8WiHUunmUHKq9dieJ4
T4QQf/b3BnLry9fCO82O3qL5iJqyLU/bf61OQTi4g6ipHjXx2rB4fXjaj9I2yET5
q9H31jDpUmO/Qkf5yuvQEF+lMBayFYMrGCvThR4mlRXGo1Fm+7yFvbnz52NTkSKb
MzhVhDzKTCFGsrxcEBBQajNJ5Gbl8CFS9lpMDQTmvv79Yg6j9jppvkVw0tEP1Nr+
dK5FgY7hkp9uk0i/nhUADor/4drTQVIkD2SD1yj0IvDPOnyVgXs6nkZYtsDKwLlE
NnbaO1NMsEdz4uM+BSn/Iu4H5jD/punOFws8GpEVU2spmCWO7a6ylyA12GRb7UgL
1maDf8Nn7XuTvXx1wmrmqR+4o7DM5iY4wFJboQUxbDAiuIF00DLGVMTNnyKcBu+W
XNcv5KY0Z6Y9TYTia+Hkzm/nWWEbrhk7HPcbMjBhQ7TaxHGZUdxSolckkkqAu+ZD
PLeHS8kbmerSrYACpiBvIQY9ZqBEiyMKJ8rWLgm3kXDpMjqfhb8IT7ri4+rbURus
m9DFXWPk65JwQnt4OBf9hinddUDay3QjAEXFA7WITdtGrB32h6l/5d1SELS5bF3J
xEBdokXRUgPbi/PZjgvsdm6yLPI7bTJj6uWNUoFf+FXWe6Hwu1D3SvpqcCuYH1r0
6xlDMEXYlFvcYry1HlrARDe1gLKM4CJiNW/1KWkcDP0hqOnucHZLOhQlYKi9WkUN
dsEW/o787Ph4nhf472jXkbY87rEoLpVQVi1Xs8jGtCtTxDoyzkOf1UCLPsJIxQBn
0htnhWJRzDTsa2VTxzqoelJOWMhnK6JHGtW0JLoJmJ/7YaAvyk+gipcRiamx3Ghl
w9Dbi8yYEgpqDpRA3dY1pED9VQZvf7POfa7ub2evJWujaQ2D+MCCILzCv5cWYC7b
JlSBi1OyHmPGvy853LobQqc4KNe1EEWsqmxY0Lu/QD1fuxTbEdXvhfRLbgY7RrUX
8D6l7nReLh3WZoZd5S7WWSCPkfj7aAn6/UxeutmTRYcN5Jm1PFGJtkBbsBxJOiYx
lF7qHWoNdIOSNUz4DumZIgzUzpsngvIX+RTUgQUdYQfx0iRi/1F4LEkKQ1KV5AJB
0K/X4uLzaIFZsa9l87lzKcSo7qEppPrG2b1kI7xPSdXTN655g/NaN+IL4+pNQ/pM
lasJHzMm4sAHFNLNb+t8YJTIg9H+j6+Rj5yVnZKIRx0A3oKX8Woz2P/97g+hsfa0
id4pWtIJDBQX9y/i4M7kg3anAy4FElgIdmRNtwj9X/vQrqhjOq1z5HmlCrq15gYq
xLl2Nl9CZLrhkHVaP7t7EBoFYwiLb6Cw0miFHk6PmrCHT2qvkgYABeOOzW02QdHy
qfVA3rh7FvWMk07z+3hme0c3iCg4W6hOt2LxduclEN5VViKa5nuzBUqSGsNZX+Qp
EmM8m8a9mlt703hTZfynh0g5DaDSv7NRKxGa727YhbkK17aCoUTo7c6e0J3sO13k
DY57jLuQgjTiFZ4KGLy96yDM2G2QNq6cwT1S7tm883vZMtPmYAC4DDuU74X5S+cN
Up34o6CxUZ8Mz49s8+MMI5coomYXI7uffndCSor8vgXZZ6lYkGRk8Ne/iBHWMu6x
3CL55BenTIoXLcDt199hjrpyAm6RKR/GOtU1Chca4tl5NvwLZHC1iGObxuIVnbVA
bpjCmdfGT1WelKVXPrCUJksuaVfnSSmjK+ffjyq67WqNlQDYI7SvdiiHmLOt/tfL
NVQcndvFuzsqaKfb83DSB6L8lepxIs1VyVCLxwdEGfy5q+RYJR/tGwKhMJC13mZa
bEGmddyEBtQbkexDAycMTTzHnB3xlrwcYxxJG6V6+WGIIVceUOtFvxCwKY29515W
VbZKzRTDaYB32/i7i/5tpfPPRdvd0M3ThXkNSRH+zcZPmfPlHefKHdpGoq5WlYdM
Y0xpJr8hM3KtUh2xZvkzA2e61sNwjEI7eNO+ZvX6DlkZjo2n7wIhfzelF6H+aanH
vaZWQLNmtzdnkxhMRyff1qTXGB89Ztxt4ObDXd270Gpp+yJQeh1GYBMDrGiPIOo9
wTAfkyeoEHAaNBTIXEimzPuxtfelGzgT/ckkYQW77DA0p4bKL5U7OUezwAigSV4T
dyVoYI3VxwQqd9KzfgC/3Ys/13CJ88EICWmu+fJX2xymZj5befYj87s0DNbbqfUq
djfamtFfD3E/5nrHZqcVMA24bIaBjjf+ESDl3aeFKTCxRiy1DhfI1HPH22ZAhC14
WJOm8qidt1iIuhwpK4OQwkMDEWIDhWBDbyoEAEgITRCuSp4glmNTTY6HFrV7kt8M
Kr0qZbft8DY2H1UGaDpOnGE3aDRRf2wATJXFj31vpxsdqIJP26c2Z2OGL2xsae5U
Y6xfhSPhig/MsGhRyodVcnAW8DccyTRMEDNeVb5xe77pFdCCZZLWnt0jAwcJM+N0
YYgT8xK7NW/EwA5EJK+GKfbfLJDoNawyPHjusRa+gsRMZ0bPPRkNGhTVxveXDt+e
NeTMaTC+GCUWtRhWuM8X1Skowc/gv21QyIkHzCmAdORGtBdEdA/nGtk60XiVmv/a
rJavVY/N/zX3UBoWdAU617Vew6ZEt4eyodSsqqRBKeByozzInuQleqQ9NWO5/N3F
Nah5EJlpHl7MWo8xuqQXo9dRhWJ3sm//dHNsgmKYP1Wg7VUGw2J5ZyuE79mdc/CC
k7oxZ5EufF7fZjJpTaKTWlDchSVx1S2NEQBuBuVNefrlBlXbzaSwXY9pdLk9kNA6
VkU2czNdAg41pCTxRb266WxONFFkr8eWIoAbzxszNxjxZyl6DRGFM43MMSyz1jUJ
cGJt/GMgVRHeJRTB4//o4HpN9Z1ikT1gKZqDbIUqfZUb/hvDKHyIEkOINVeEQvAj
7vj28XoDkRCFEaX4WhtqY7iP4E/+ApOp18X9cqfJTZEte4buwniACKOXtHdHIqbn
jCjkDNkdzBs//IUDNKs5qniW1VHJYK0eQKOzS970nNo2NJiLwkaU6/mxEev8QrFp
6h3fJgLA7nP/m3a116n1eNT2HgzGPi/85BDZHk7zxXvVQqh6m/8Pxu1z8WmidbqT
bpaJOXGdvROdJ8ILBQLk4TK0ucNKlQjm5LGu2H7n5oqOdEUjBFW2UOCUqdz6gDws
HjLTxTdX9mRdvl6DvBpV6dwB5zTtWL/T23Xcqd89cBjRE+TsJfbaSIZbRtEfzb3G
1tnGKqTwuJ9HzPOu78M//zC9aaBGcS457i7+5mbuY3g1C2IPdOyI1+Oi/ops2Wym
+PJ8kHSUmp7PETVvI4pCCnYuUnOquLr2GrTRtzdZNgVCqKQU2Co22X/wbXTi7kQj
NIvGW5sI65UsJYL0psCLi1iWROxi/dUyjMkTOJDtl1f6EOf5xuGmi48+sB/bKY1d
oWdFt1cizNMunNoShqaA56V1uUyepKZsaJ+c63PnrgVUiEVvWBRTwab25g57D3Yi
L4KB6LqzbCRfb8sh6Jy1g3uEVIKkjeOaliVy7x+83m+Ax9fA7MMVwSbnspSk3K/P
nlKKiGM6htTpsEpuQC1hQ2W240RTZCGRPczhrQjCwEUCi0+a6ES82c4u2oNP4J52
IrWy/l5YXlLOvkIta9ptHNsBu8Bh5IBaCVbff+5Rtrunha2GBYXpEJWwe/gZR+Zm
qdekImSqBUe0DcxA03kt37MbRtKxOy2+oHIr6JdyJ3CRusnysVUZpJIJ+oDfeu+Y
N5q9QMj8ePoAkjldZDxLlvkb+81SkCoTzFk8diaKL6Z7Lg7X1/hLewloDU3iH0Fu
i2pjLmmXIdsCv25+sfSnjc8cKANxS0UTlINbu108FtoPNO3MUCj6Mp0P/Uxf4kPs
4OCPnNbicpGJYh0ASyDYAO1UBvmOAZ8jDvMFqCICVtpT0Li+KQ6DngfmzhALGPOJ
AzNTujBeABVbeq/nCQWFuNeL93L2YSqbHRkItrxXkJBrs3I4QyZ+ojq2tg8ZG7Q6
N09ND/Vv5nyiaCz0nMaRKH8ff6+foYesvzkkujTUVKSRyMEuaIsUV8ejyWvTA5+u
w2fhc//BFK9RJFVdNXmnzn02BRWDghZCfTgiyUWqLLrN4KULDUH5lwGp19Ox0xnc
4IVOlvcDa+cJpxcHr5Yw+ONOHoIWXTz8WCFPRMZ6x9W8FW1d2fUYwvcgu/2z41Yv
9Hjt2UHlWTB+laJ9KV1XCKVNmyKXbLzvy/baoLLG7XPnnT9wHG6Qt3u4tM885Zxi
tBiRt/FyHKWU6rcN6P2ZeacCYKQYYCgTExmabIX4S0Bda4mSNK8Pj8Rn+PnOY6dp
JVAEWJAWxjizgil5dd2uZyqZ/qv522UNdH38U82uCQ6qXCVQ5Xms/ySN9XQMpAst
r9QK1PY+hPvN7gz+N1pNBsZryq0mPfMHvywMNkGvXwUJS6IRvT1G5jey0CA5kDPM
BeXom7Z2U9Y2/yF75AwTATwl5tLzdD37cwTMIYNKnlXcgRbR+iSKmfM8v85w41Fk
JFRGgRV+5m9PkRPBhrxRyguLQ62J+U/l1ECxwmaZp9l2DJzRPswOz8F5RwmhVDIn
1CbKMAs19tNI5tkOmAV415l/mSsyjSoyCj4r3zUwNnR690uW1Ky+w0KfxMXpIhkR
fgyN2xPCI7ETcV0Grtin9c4MWDqMkkLfwtJ+d/ATN56nCjRAsmk2uio5hwN1mov1
0eoRxGujq8Z6Jt5f8pYRCauxs8OB1CI69ApW5HtAX47Vy3BJoEmRPdpwinnvMYqI
JNSD3Wjh8+OsMADP62wjw2tsgFdi2DeRJX2icMKtzGxz8isE9Z7MTwRXhQkp1FeT
iHXU/TPiPwxvzANaLD2atnEnhzIsWi9G5vbqDm8m4cP5VpFOzZJIpmGqQjEmeS/F
hGfHanycv8EywQMIWZ3CHztTv/tnIM6moO1HxsSxZNtbOf+/WE0lmJ6CJahQr2dZ
1letUOpiCxiXhIhaumVu8qIJqFve9Xc6IP1YZlkWUqIYztgtJCOftYKCW6qG2MnY
JhEp5uDNaYMcz+1oKUkSjLaHzdRu3MBayErsGn0C4ycVPFRXy+5ZA4pSz/PxzWU4
C23JAyAp/eyi45aE94NFAK8P9VqEMGR4yP1WLWFe+G2xT/iwdQxUc0OzlcZ4sOCK
HNK094EOm7enlvuDkmiWbvcQwbAr9c6ZBfRKyKEQiLgfY76IFxALj2A+7s31/3X7
Fz7kLdCeolYy81teqtb8dbeuDnNHUbxuRl8CgiQzmS6i3N3bNRJVP3s4iY7JwEkf
wIztBgWZmMdEHihIELR58nySFkAX1ZFB17W/wm9aOjbURsgiLba8khln6hHh3dD2
ZiHstGyIS7WynGkX5HlIQk54E5Flg/y87jjD/u3MsmHUFmrwTLug21tlWr/d5fZ+
nR6prKMcn7uCgxjW9baQSQqL6VuZDi8FLB6dNC4UkaobDLjrYcmFmnjZ4O0hufBu
Jc4VLm6RvrQnFl5Aspbk+7Dkemc9X1ys+gCZ9lN4RSnYVA25804KiMd5RB1hY1Uy
rytNYkVwZveiIbGVTv4i3CRlSiuB8NnozFv/8a3vop3i85ftzWfGF7ZmwbYClMks
VwFAvr5n1PrhYutGWUFsHyQ5n0PlANe3jKiq53OVj1K2iTLkNun2JFV+M5GR4HRC
RwC3WF4ZZLImG6LFVRhGh8j2TByk5Izw92xI8b+7UQ+MfS61hVDLynXs4DLL0M3U
iLYuQSq1Rt8rHSXO9rZONmXdqvf5ElZ9KnMqPvlsUuvUct9zxSE4g5sm7225GtC/
lJvSW3OyVQUTySrUTPYAVXKUBQwr6NwYNJxH7bMYWL5gq6JUpcyz/lW8BZM58ZgP
qFgOkv8fpuyhIqEUQbab0lfiOB9QFGf3anCKqlS0Zxx7+0qSiWW9lATNgbJPAbkp
qZnHt7zxXUKuA1KmADQ5ynHwdgwILyrblxVNficFgfyFQNVDheBBCNxI8bgYli18
wb1IczCPwVDq+bMnk9/BQJz/v5WJyRnNC2wxutI0dQXsA5hKWPzaomydA1aJSAG+
x60UVmoDBL5n7KF6Oj6vV2Wqa22F9KnH4sdCNsWOOk+mNQB9vmpS7yqgPt4wSXDh
bHb9S7BQRgQKySrcFUULXez1WrAc0sivCaC0gUeoMvVDkmECFjBUhgICNHsG1/iB
bcaW8u1DhnZ1TT1p2HqL+zJSnxd1PqWxmqVpnxUFov17kv6HEAJtaba1UFxX1/Ko
meZHpG+bM2X9PeQtHrguV7so1GPN81/nh2b2+xRwX2tC3dhBaMJB4gU2dK9Uy6/I
92M7g+4ZQ1FDAucNc4bhxJgwbEIHXN2SFIMPvd7CMbcq6UPsG3GhJ5/zPYuBGAn6
ntjA4eKLMplJi8VQKfGzRV3fX6de9kIxlWgnEObB/DhU1Sr9eojieKYGG+zsUa8q
QcGtD2+0SGna8gGv9NxGfDP9VSyWnDW3vs2ne8k/jQItIS7UAEInKQxbqEhbjvVn
O9iG/YqbXXywp1S/+toMuGL6ExEkRSG4cmcYZJYw7GVqzeqwnCvQrhu0zNQZFA+o
ylgW2zdxwvmvrjW2UX+qmGCNU5FWRw3L1lzKMdr4KrebkxYc6AMPe4O43tRtVoB0
gsHvaemZYQG8LUc7czKvwkYs0A79PNfibpA+v6NMg4KXzEECEG4Uev/c/q7RIhDX
9IHru32BQKN8HP7QCP9g2Et4vEKwXDVxcL8jUtwRXvkPyEImTOEab9X6GzXmLYr3
fCWyFSCajmM6jwCzcnLkM6y7B+2JLoyrSx2rczB8+6Xn43SM35qUUeFHaJWr/WvO
7OUXEcVavXxr9V3jK0rYsfZx/zlzA8uRaDjrdXSnM1L2xY4/6LDTbdhOs/JynGff
+RP7XJhfCn8ItMc6i3ECk1v0ydrFy9ZBLUePsIS97PhOCJU9mdBTqUH9x11DgrNv
R+91UmR4KdHE/ZHQS2TAU+HgnS6vcwIyXVDeIt2iGNpUnsPoqEs6qv7i5l4qJrs9
TLupWMfIqWAfrazBXSasjmDPMHT4OB3HRaiGHunf04IvZdzD0D+2W8Jxv8V4b+2i
oMXTgMPoJG/AKpfjgUGije5QeAriNSuOGv5WGeHFfsjd/hWvqnQbD+LdxiT75hvA
vJmEYKsPiRUAR4mG2fgwViEq0qJ5mRtJPVKdVpWPGrtaig5T+7eGgu3GWuaR5mkt
`protect END_PROTECTED
