`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H7TmtYf379w+SCdTFwcQXvN36/0q9v/sYKlq1iXvsze2vcwXCsKrLmxxq5k0Riy9
rbKRlolflmEl+I9HnqquKylV1UL3aXrjBlWkTDFQs9KUAiRnwf1qB8gMFpDGMdfg
nus1HOKSTkvOB7OP4+1SWWB+E/zZ/lmlchkOtxJFPW2RAi4zP11MUaOMi6PLurKX
qqUjpQKTzudIF9AjD5i+ucUhwFlHHgcGV1MYl10YRfi4qsnU65TIpbpmC4V3YTbW
AnjRI8+F2IfxPR4ZQqJPHYpvA22QqmPi5mzW6nQQevdJ5tHorFf9EAKsz9q9m/SQ
AXRioxRgjVMDLIBHDzeeXNRasi0M7RBZf+nY3madyfvCu1aC7IqWo5UzLmCQq0QJ
`protect END_PROTECTED
