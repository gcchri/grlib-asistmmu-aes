`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XjGQRv/SOM/bk+hTZ1Kv1W2I8u3wdyhWka9ul4Vq1OuRYXtxfRLO9fJkBN2kNWsX
0nAHxWUWjNLGdc/s1YJ5omOc6x9zZUHlNGTT73GGGy7Hr08Xib/3p3+1a/sSspZs
BBd7jw6np6Izet+orI1NySyNE3aloVvGO/8LsX/uSRiqRe+IIfIyZABUiyOsEmkN
rGMc/B/dSYx6evsDHI+y0FW/mYbTrZObCnapouGFq9qjb3dWHOcBTFDO4tVUXjqL
Wa7jFDjGTTKTVNqyJz2gvFzDrT6VfkiGlAYc0UPvjXzI4EFgR0tQFwJd3jvU4YTc
SYp4BMa4oJd1okXL2QXcCc8KM6vcaqUNRue8KSzQlmm+nO1DEVBNvUPQvt7iHHy9
+DVnyxlsXztdG1lpoqIHp6UMxDwfsiorMyyDaGOLq1vlFbZuhDcEwMzKWWO10MkN
bU08TOOKfGVA1wIIJrOvBTPTZ4j1cxD730yqFWNApP3nENRv8wb4WRonQzjaWnl4
ycYu2gX59DttOI/TkmqCUsXkIcUNutBCu4SuJUbOgyr//F5IsBdMvP7Y9iX1dMg3
`protect END_PROTECTED
