`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gl5xTtL52qFbPRmQU/CMC2yboAUTeB9NhZe6wFj/Il9L7jINl9LL04Bf2BXs1UT+
VCv3PHZM0rRGSY7yDCPdzVI2bSwZfKbpEgxtQWXelKBfpDLcbQde3Slk9osQCzMI
imUzY2LhfNvJxQdN+YE93/OOAbN2fLLTP5MWI18UvgFebQDxQ6Bd/Xjs/M2Wiscg
IHb3gmATEBBFhbP+Kbs6VYPPii3RP02w3WyRntkVu2+JaaoMb527QLkDhWhTkb5e
XbKBSRkFWXkK2CVkKhvz9r84D8rzlJvjSvqLc2oFNbCABz5wewEJ7BmhFuE3H/0I
Mq56pUMO10YlCtBJJwWabiEXlESeFS9WwIqAOkvhPJYvzIGLUFuNPG9xNYmE6vXZ
FTAbSd6o8BgIXOgpILbAX44p5BLkabB7JaSxMTlakjgsmqnSAOkA2EDoYXX7nYGF
pB8lB0RgSerqnRJ59ZASwDeJ2xMRaWus0bA1pc+K1cABQrTtieAT2guD5pNkEI0F
rsMcGeKto1aq3UOPhfT4d1Zeh1flcSOHbhZk+s/X4Zt/Wj/SLMfx5AR1GUWMDqj0
Wzp5AtLslpqH/mXV5frTMfbFZNL439Io95Z3ApXSoiZUkeVcYrVfFAeabNhvjHgR
m6yBj6kdIVJ81XyjKIXUqRuvEnqXoyttMXN6ZJK/R+YF5ZN83/TZMmIYX2jn6jD+
NkH/uxJXb2mnMzqSwnuwmBIoe1D2XS1jWILZCwlXFjnEViLRHZhxPsmdfCvnWU2G
A7H/llg4+a+LpqfOA4anMQH/JFP1XgglzGe+AoZV3NO9r0Q3iY7WU9SbqUVdlalo
U1dXD/J44V+O3DHg6OSFZkjLZodEZBjSvHYoz/iBV+KUC+BKBnUujuS8VtHusOOC
OSoEA1yxMm8QVpD4knMrGg==
`protect END_PROTECTED
