`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
unVSeqBPxbpt9nbhEdo8vT/JqknxOlx/s4sl2OSifxmCoAq4hCn5N6umtqXuaiwu
BXeUniVEzDsOi+6l1/FIKpXyZEuA1dDIlLHC2z+qx00FEKVRLMPf0Np27yjcCf0O
oc2Q5mZPwSiBF9LiUtz9QPN/hUpw6yyOCkecZpiislqNOAzvseYAzkVJh10SYNhI
zBPIWBQ3w3ejfXxm81eEuE/1cQLobZ1IlnZf3/OUAIpo0vhOpTnBA0uY8iGVCGi6
ircsTL1wzx1pTaUDJ16hr5yedXFjKZc6Fsi22ELLrPEOjtb2FqNDKLacmPByLe4w
aFlkg9lU+jrIPArle8OJ/C6V8HR++AGyrlpab51vreVDJF3OmkgxYFLyM/9vZgf1
9J6NfuqcsiMUJPR9vsY0D+SzGnj08kydw2K6DtS1sH4aBdStswwDxyu5c4uwMppP
GUWlocbGbrXxz6Awf1Zj6NXsBf8o7uvLaiLdLkt5t7wzOhDggRmwRwh1R5tTGLO6
FGkmnjDYdO3mtzhIeAuNBMbm7DRZxn1ASSr6PYOD6a5u0vtwtZSsLYzjxzbLGeye
aeRhJLAJbkH8EvPXFFb64A==
`protect END_PROTECTED
