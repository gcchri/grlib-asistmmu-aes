`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jQRJ1rGLiE/ImBVDMJUuM7daDn+jb36NRFiHoRvE/CW66p4qyet60qV+Y5ANxusv
iHVTD6FlyEdImBFNZnEGoJc7SjwXlj6UWc6CQh8sqw3GOGE/yJJRB4Ns2JvAF7Xn
B+ja935O05lincSBraz48CxC91qycUXPUyibL8ZiucEsJcZFiP/aepe1NDXUJBeq
3eva01DM74klfj7xLefTtVxDJ6LojOO+fuFy999pYDoQEacfCDJZQqdB+xLAJCOC
PpgLqeF/pWyAZlXsz74VIafoV9W1upeinf03ucTmQgs7FkI2E1n/0J7t5kFR8Ox+
G7diUPomOxZI2MoRC3bz8zGSX/+HhDjo/u7zeF/R1ee0cUi2i4yBuoQghE9seYUU
dOmegmneknbrcl9pzJb7vnRRSr9BQ7DEIzqso0f+/4Dz+zPr/qPW+w/Knz9+wi2D
JKugGYz1OPkB2Feoul1tkVxYo1E7t5X5qtkrKBazfDrghzCtkn5QauGjBOwGkY5m
Nh2CjogrLGTK92CLXA5dUu0Fvu7SN7x/0OKdj+xjViMHt5dN70Muny+SDFMslnKB
0OSXuKm9ycLcLeWXDAQdDnpNZntGlFhzCNW3jLe/3T+mtYRwOYCslfWX+S/Wvpqc
Wtbj6v6zBpXs7meeoBNYtNnJlBr2YHde1i4lW9Q4FYqTY+E44qF4AsaXU4xHfTuE
H5lvqV22nLs74ZiBza3H3V3WF48KV8AXo9R2ayq0uswwLR+YL4CB03HCKU9NQ9YW
2CLge8G1qwWMmg+oazTYvQwPay317cJLV/ughv1yVPzqznGtqZ01pHqULT1CV4jj
uus+QY8ycpauWWVY4KJuvD7nsYdhEYkwYmqc4LnzOOIR696JgozBkN4Ja8vX5Hs/
HfZqn+Fdrr4k+odl7ubI/KWDhwfrkpLPbo2dzkc8Pub7yWWry3d2hYUMkGHZ7Oj7
CFX4+oCx5DsO+mrQ1YV9fJ1tzpRL/NeBJtW8r5f9+fA6WlFZr1vSqLJC/LDZokvy
NL/QqhdFF+jenQMhyTFHiniNffXFeIVHZHYMRby2CUiJFvNYTQnUOlQ0a6hQkYrm
1zLEAK4q+dyO7sTeuz3shl895ykzd62aaaON9egm8HOToL9BLHzCM/0VZyV5QHm1
Jy8jX5exqgVEWFglilP7NXibZeVPAiMFwnBEJihVbM0+sDZnC9Om5s1lcsCRiUnC
UP2O1NvvWYv8Eu2PYgkqxpbmBLTwhXZOFuJ7ej1iOD3FOQtbwJgY9AUNBBRf/Oq1
vXfGFtQ0V9bLRlyDdODzkSpS5PZRax44L50BjeTOXaINl9AMxUrwrl2hO9SEB9Jf
iIeA4tmWOQSN0o6z6hnGt71MlDWTzCICICyZLKxm0jx2U8k/M6fYMaQ/kTLcIfOs
bmfYcupUAaq/vpMR1Bg/AA+ZsB3Xa82pt20t87QVWzdUpEwvc+LbqNKUZGq3bvIM
anA9msrSWa0RWmfCfo5XpnxFr0GUw9OUsZX3r0aWpWNW3nnrMmmwQrNgLKHNxS0R
QOe13qGLyUZcnZr87cKVby/JJc8MX3ddfVXkVhRq5WaNfB9EdZeGzp6E9JGaCDv1
5rLS0qlo/hVAkHsmWrF50Tp6B5qWLGCJD2Pk9QGtIF5ZORmzlsvBf9/HNtHtB4Ur
M6DARn2NkiiRhNxD1n5awDY5FNA9cuEt0DCyJS3Eeu9yLEg/OU8GWWpm1kCwuJDT
tgJHeXMb7b1qacca/zT5tGu1t79BNScx60BzP/IV2smCBUUInJDBNMBBinQGOSm1
Zq05Cxe5sUU0y93AOAwCeE456m2ZlEx1Rc/Wsz8oa3ErzCSiw4Dix6aoBPVPVJBl
6Tbp63DVCN1MqXBbWr19V100DtEEWjrCiI/0vOh9C4IsKt7QwXzgg5GTSSiyg0gV
XDDB4zF0Exm3DBlKwXIVZ1/N2Dpr9a7UgxCz72ehrDUqbZHzgscassrnQP/hP+Nq
Nhu4/eGX+G8bgi77ZTRUMsjyYrp1ccsIZsj7NWDDLE9G1HQMSMVXeoRYGFhOeZ/U
z3QsOHTvXGkmLujlpUOpCS+TXKn442Kxxb3ZSGBLAhrM0t7VRxiCHHBvTssIQaZ8
EmxsfL4qNEK2jnux0xmhrTel1evirAfAlgXz60jwABIIFbk/dBL5yTrzh+Bqprnx
N5d1YKVUVbxwc6l2vLSvm0z7jLz/YzSnwISngZFyQQT22bRLY57YrvGB6fOgvRJl
j5bs+ED0Y1PKRi775ZulKUDlTzo4R3YA6CTHQQ4mm6XglCoWVNYSP52D2+Q8UxDb
MQ38wQ2xUjsmwDuU1P7tXiO2f0guMVjXPYTegJ+vi284h1pQHj4JvVHOb7yrkNWA
DAX2CpPTJr814uQCOTopbZrPILszJ3TQ/BXTfUk5+rqNmiaDtAmR3d2iIynWBqxX
+7vH/u/lpb71srUtVUqzmbVxNWWcTh+JhDS5FEx0C1r8wKeOBLgIYOm5jjRxxCgk
TtdB3CvAunhw7VbHzfAPIpV/6HfnjP8rU6kedB7QMVVRy0jT9MUkU0th74rhcarf
jO2GScN2FVYY7wEUcH0K4UhBnqyp5i75kS0bqUyXM3W8KXZlfEB43Y3P8TUPHYoN
nNKCEaJSTc/dNTVmoLpzYbtNUvBz7f9pP2FcBM9MsIZSjC0xirSKxKcjKBgV9Rit
W3qYXc/Yy+FQXhc3+vo9hiMS19ZLkbXmgjUP6Zr6zR8TIKPB1u7W3Pfv52v3LbNt
JoobUxwJwnGWpkl+ESChJmMv88P7n94M71hmNYGnttmmrmBub+dA0v77vp9/GEAf
j6I5gLMqal3aZ0chsP+Zuf6kQXnKaDfAmNjCPivz1nIXRg+inrWuW8mcqwuZMMij
wZclCagNVvQUFgMmmnFoSX29ZRK45VH9OYxDO39PQLX650xmjSsHMTQTPhdF9Ywf
P+/zkcg8CNWmBJAOX1QSaJTAyFGBPwpavplL99RV6soefbl6LmE3c9rA3QhspX/j
14Sh4JV/Z8R7mAqqUjSVWmCdj/Pjin9apC+jJXSzNbesRnd1ePQuOL5FShlFo6kD
wSbtPk8M1U2Wk43Z8sxdAIaJLhi74bitzLEVAq9iVl+qTTRwE3pkDwfsUbXHksRs
whGrii/YWgNfHegQlS7ehJzNiFy59TfNuMFvNuDV73tb/Q5Oy3ZDmHiEDJFOc7w7
pRaaeXB7hRcQwFcnagd2XB607SP4vg1tamnTXp3WC5gnu8vBjW+p6zryESqH7MtK
hEoVyzs3yCAVFm4IECROJNMILLm+8uJZ/aiG5arnmUeA+rAFiy2acHwQV3Vy0Ka2
I5CPgQyzStMVtL/uC6EwOdJfjQJhsvn14jmwCfuSJBLs4envWNWpppL68G7Tz5G5
tbg4W3+c2r4XHg4aPmQ3LWO7dS5bkxQyyGzIpfFrYPN/FNVb4WvdI2wuafegheQd
91SKkZHat+tkil2BixmUPeJbTAzHvLrjjyp4w79+NLyCedkYU+jkr+kowu8FoSGG
tcKY0+S72UO+0MNflLGG68IVHKx2moYirkOnvmT3cq7FAKFYu2qNxoxkcLTX8s2m
Y1vIKk/Ux1c3YyPS6BjHKnsnJ2JnNEDOeolLGuc5fpyhwcK0i8KkGfKPVhW+pvTg
4Rc5BPe2yIhzXA+xsm+jPfxP8MdxYzWOWhSdjF4NrGTV+VIKNX3uu1a7ud5E6kUE
GQAKGP4YlBlrfNojARf6ExmDpZEBzpfo0d4zD+652mjbDwLQQMbicAComTu99cLV
lVZYAqpwTiwfgsvM5UAnjA5Lvd4h35XQLQuJn4LnoOjy4cRguYQ0FXLNeiGFiLm4
WXV1OTwNyBH4V1W5vRUU+XwbV4oCDYALu+Qr2NyQ4v52DycgIkx9wCEHVm0JdvE2
NCXbaY6pOb4rgrBS6MNPhS/p7WECaVhtcKmiLkp/fkuS9h46/UVxmwt8CYN0IQRb
WL+v8nL62QsqpmvF4KphIe0rd/Bt08p8dhWPB52+RuW1Wo6Azs1j/T1eNnZMSeJ4
7q5vmChz5LALWEGmaKTgbbnKFUQN+lhOe4jRCFQPt2w0wK5buXpIoXsQAsp9EfnW
zOAv8A2+eAwaLAbnWab0cXfvxJnCZsa9kZSQPNWr3OHd2cqmX8c/0DYo7o3tW4K6
`protect END_PROTECTED
