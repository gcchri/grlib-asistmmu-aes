`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3P1vdWqV7t6EHkjhfGKrMb+GGiFyjUnoatAM5YGaqZcRVY73XzZ6C4EvNGAhghaV
uZ3OXH6FOdnpgUWJHTBbz+6DjsEVaUWvIh0jYl7lo5RDnz/TOi4zaz06CT0VoT88
jN+RJsEuBtYMG+dSaM0N2/xVD3JFAvOAvRDb5cjjwNtxNwIk2XkGgYtmg2KqcJH8
9xPBKZiDTWuzYTsNX3oEKf6xgHOOYEpGENZR5Q8+zk17DEbPgok/Rl1ITn1liofk
euI5eSC8T96GEdm+sUUDwBMjBk4vALvLO6Zjpl8VjBga/EoJYRpfFyo2R3X4xLmj
MtK+F4Z+IqPs7DHCZ0NkKoNwJjrd8/xMIWDQJFFxFmHoZ6oDTTUWpriUsrVnpkHD
nSeCKqt9TiAKXPDMH/gnT0zVU7PVj86dd6mkn9aKrwuFxsM2gPTpQWomXKc3rnBr
i3EyRowdGcdRFRBCGXydp0G5MpPuJG8hSu7xE2Qt3vAWbvRoXgNIhxLxbKWOdrBt
xODcm96+w7XtBklTT+wrGuhbsrpGY2N5GXOS8iMiyImTFt76lGI9Ncj4lMQPGnpM
H1fel9DPnp3juXBTKGmJyZPm9Vb8HCgJBsKcmg7+Mfew+e2lHV1G3MT9JK+8xZDr
uok6DUA2Iv8Z3kUNmecX+jSNRh3TiBBCqY3RW69wHvIcUv+87LbMKteiDkqXN7/b
ox1pS6Krb2iYrsWGz1NDBq9XCsQkL7gIaoYCx79ExE4Sh1NcIHTYv9x7oJGhvezL
/HyyRiZnpu4d7McVX4Tsa0May7q7CTou0x2cgHjVch0X6pKtjjQP62F2ptsDEZhT
K4wF/J9ggemr+ljf9r97n/vKxKYOmhxJHYgbWr3UXA0=
`protect END_PROTECTED
