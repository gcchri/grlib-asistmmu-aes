`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HG3nme3uXQ8yAulGj4B8rpQE/Xg7OBOvq1XtSUJ+doRlyAB/dxgr/CYjGHO0E/Rm
rbHECmyr7CrFukXnI32ZXDJ01h/HTjRY3pgaft4q6lYLBuCRvOhxKJkcLaHyZ6KG
Cjd+GvOdksY6v0zaVyQUQVAP1Zj0zbMtV5PilWt3Hp7HPJ6WQ+i9rV8SATH0nnu5
jMgLkhmCWy/TmWPxTMTD07DWGGHaG0WD2Bih4xd+B5CoO0yAh1vSU/pBuf2KNjwa
Procaj0Rt4y9WEGGZ6jwA1y5IzbKogt4If2Lty6ZBpSqONC4wIi+GNTU19JzZXWh
`protect END_PROTECTED
