`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P+O25kWSsEx5cDu4TC6XmU8gaFEsFuCgnzzOcdM5xRh+j0mrXhq0OLh1gF9WEc/E
f0CuSiH9F4LQVdInlYgXs2IzS2HQflK/3Zoog4y7pCFUzPDgGjKKmeCjNqze4F64
ZK6SD2Ud9ul57fY3wWUi4LCI8MqBnhFoPZFfaEYU6e5fgZlsxOUub+0pUY/7mS5F
hy7j4zkUTQFUzL+/kKIHdWN4gra+yI0mrlJ4Iy9uw3MJAemwiHSEbcCY+Yippq5l
+pJUf/zrApslxBXRj9h0JkIL1M+tY/vBcI+AYS0kCFLNhtqeviUwYfQZdixEXjQ2
rH7wW4/KSUDAN3lpXiIvZ6M8QDz10o1ETP7+vT7NFqgz6X2O8zLvea2rahhl4JTe
DT6hbmYMaRbV6BZn7by/EA==
`protect END_PROTECTED
