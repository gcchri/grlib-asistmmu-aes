`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7QsYVb6w50Rf014nZAfcNQJjHeCzVKmztrGYJnI9CkgrR37zLwwLstnY+au0PVHZ
TpVVLfE37ky4N3I8/mMUbahgduVjbIjgl/jR6KzcSL9ugHd3/VXCt0Srotkh5z3P
SlpmVoaOgKuPagqmvn6OJ4qz15lzPDvQTzWrryDkIqlRb4jUwFAMatCY0/KcIbBV
/BmYBQNVpb+R8KWTH0MfHTCfkuoS4+SBH2jA4mTJ73IOb9321WF7Sd2BxH/Q/lyD
3z9Yyq8a7+J17DMQ0YU7g8bub/jNjSr2MOFhTSLIE4X3LmHnS51FbDtj4gtgwrv4
M/p4EyfQ3mxTPqKF1JoD5doteg/dwioCltKbdKM3z1/j/goPspBAOy/BWiPDN+KT
kPUWO6uHzxEVYTD7i3inbErO3z61Txnhm+Ic8zId67S2jeqinUJl7pgNrA8ghzhB
QGt5uAIHa1OobXawF/ytQDPHXxb3vuQupHNsrm6mwYMgxe0Cpd34YPUNrYZLEG6w
KSSn93kMnU3etAAEzF8KDK4FJroCyACXBQiqWxZbiTlR7kR0ig3yNp1EITvUIGh0
hKMfRCu2H8GTVACPDGmtEAxjlAhLknB6A2+83rkhZHBDRlHtcMRZZpo+StOt7myC
OVH8pTR56b8Osy7u0Zrp372+h2BBZ4skpRaD78SCnI7msbvuqaYOgXlQcVOIvO84
MCNXvy/ZLijc8QEphDpCFhkDDoYO5W7D/3kIJmpAQnA2TAblRIZ8TB5B/yyW/7VC
77wFUVOlrnapFuXUjGU7yw5+q9uNJdKN+7ZDlgX98utLRygRv5fVjsVTcneKtTWS
ktAAD+B7IrqlTukPQbWV683EIh+U4v3W154Qc5NZl4TDewy8mm0U5Go7xUvzqBEP
/FrbzVZayrkNLut8v/a26QpayaUfMXoNTOV0b2HDFi7dF5QIFNDWqJVsYYuouXlb
oYuKx48lUM01wI6m0kNlF17MtYCyc42V6ZqdgYnZIMtJ3DnB6ccr/qCG3TRAhSR0
4yjWQdRR01SUb19HdoqVjpua4yl5/Q/BlUieZXsfBVU7sMfgaDM1BYnwa1htiIDt
Yg8jp9DgBYmxJq5t6NZOpZBY50ySKC1eRdquKFEICEpzmoAWc3v/sE/iW/uxGGtQ
KpZ3BaH6VdVdjukBIt42cxrPc0BL2Eg5lC/opujCFJ8KpEHy3W1z8oS0FJYfXkzx
gcnlWmzAOabKMwTfIQywgA==
`protect END_PROTECTED
