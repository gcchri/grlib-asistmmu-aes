`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cn0n7up1ZLvqh5lTwrkWKxLGLG79n6w0N/HaQ+zlaJ7N3ck5B5DoKZ0r6ciWaqUT
xkhYNkBofB+ROYwz8nfw7d0bFLFOR4YquMjcK5d6KNkb9LBXMU9JHAV2p5ZcB84P
ylH/DLL7jvPTYLWi4FFRMNAEtDyX5FAlWF1O0/g/PjkVw3APyBBcb3Bgt0067YWh
/4PEwk+pgjpWk6lJt08Hc7GOEYzamfbe2pEJ58+V1vSUESCzykEj5WbpR5phZvlU
DBhuZab1Yo1213tXSTx8+GcZhgwfW9cFTPPx6RzTfzh0+OLSxz7QpkNGb/ioU90f
zMCI8CaKSKaYhjDbTGPOYhzGLFQJ9NLbEKiz5x9j4P5u9zOsAUq3p96+zx8o0/RK
C2U6PAxVFeJEiWB052cKy17eQXSp0mJit4e7jQSpaOaxGB9o1p4yp3cbxEPoGqDt
Q7bWIeORWR+Bhp9b9+aeuSCxzNi3FhfbIZog2DPOfJrxV3SET1n7ttIkqG0N/xTp
diRH8wgSXIzNFQsRFDc243SfwhsPa68+12kcLCe2iA//uSTv4TEiI53+t+nVAbs4
fA2itsFnsyIQ+2ptGMh/pymN7CDUXuQa4fxFsRwV5slWTCwKDi0uIakt6qamTR0G
nU5W90LiI1AWfAwX0lg7WAVfQR7Q6AusUCXOEEbCN1AmxQGaufmtsrWZ+1+m1tNy
NARyOQJYu9IIK+trILZNdH2FYx1cdi887T4OMAY9dMKuM2k2mFk9n/m59qN9QZ+f
3roP0ldwA15Q5phEeL2mLHk37+GjlOiNOSVBqo0UC8zbdMSt4M3gmCHMIEmxDXMr
vijYkpKoVu75lgCUlyM/ryBpojEiqAI9agmr4MgRe4e//IFKfRkpOjF3jLmSsVHA
pCGGgTUtiJgvBiBLObZngg==
`protect END_PROTECTED
