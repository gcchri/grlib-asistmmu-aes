`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gOg+L4bNuPdhu9XTcIwYvAR+Apmkua3X7sFRDFOZHAfw0ugbe5XMoYK3vNOkKSVs
j47gV4ETY6XT/m+frZdMSIy4M8OhKyslxm5ks1v13lFT5yQebUq2RFk2ovfup4Ou
WuFoIW4NhN7hqmqWillDfAS/JmrX2Bj97/7EVN4Yp1T9x8QLBsrTysN7p1+sWYoh
u1ZCIbaCzM/sKblxfBwvmKOyCTsljaN3mGAng2Xr0d+y/R+WxFHfD66qfcKoz7Jo
Mi06GAItnDj/wjTCTHzUiOnJ749DjIAfLBkyajK9EObo2+CHjQLlZwNbHoY096qk
eLr8F9zLlU1J+VA7QgDxZwBUdAEscq7YoAn6R9d9Crd2QlweiaWU16Kgbce3xzaF
urtLO/Ba1uGy/1XYQMhBLlKoqIUjU3tHD7KovEIO3qFNRHxBYVAul5zrxuo3+g2F
`protect END_PROTECTED
