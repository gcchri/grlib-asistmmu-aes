`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uiLmjp8gPF20yr12w5MCgyqTpEGRwwlCUMgxwpJcYdjcxLSwti5JE4tXVtYQJp1z
LFih68Td3VYPcdYner7mO6phO6KY7AktqxA1hcmBN6xxkC2qpEzRtpxGsmvp+fD9
BiLydCWiyC9kDf52vTMQdTx6aNaQcgaK0HbPAFT0g1rvlCaPV/8WikYO1ZJPkR4K
SKbmYQEZ7+0X1yVobD+CNHb/ddRTDjSK4aHABSfuedtJZFrBA3AWFX6txcNh0WLS
KPts2y1opHt7bW+/9a7BiVBbT69BtyNEWQCiFsxBnfI6UHqygZNmyiEOX7gsoGk9
oXVQm0sHSBcP4JUeR2Gp8lba3PW4YU4nKE3DvjXWtJHgq3x8ccumGGSKGItUNlSG
fj2GHKKdNRd+SdGmbPlTB5yBNlbf++YdRqWbwLpxIrRkJQ191hSTUVBc8G9g64VR
Wv6W6O8WZgCLNwpgH/8JIPK6ut8F9y4XkDt0xK9AGVTDq5qy9pCCJHi4YPn7Ij12
Q2XjXynOQxJou3BaGUwox7cHNR7iH11DJ2Iz1SUfYGkoxPZ+pyQmYnqUrffL9HwM
FMWw+IMUQAlNRy97TtPLaW6K9qZM7ueaa5W6sSWPsUE7MIrqt/ES+tUeGaULUj5E
37J0APYMf3+JjI68UeLe95NcwahYwfbGGpnYMNvGpkz+ExBlkirNXLe/yqcnscsw
RtKpKQZqyLnx6OMsIJu10r25BEkQTDmjikVKrQY9RRHDij8UGe1KVNnXH/VvuDG0
ixm6bvv6T6YlGgBd47q4vCx4y8uEUIo0Raz9m9rXxXEl5apWCNQAd0wzAs8H1tJA
LVw+OpZDXj+GsxqCKgL//R4kqMsHwxMY/7Ng2gKgT3Exy2CINHLW/Fan+gD/+vWJ
dYxuBfVn9QCLeoY1v8EV0gEPga/q5TCm/fO8RUoSJWqolyOi4HXNXI/+CjDN3yqs
4nrG7NaWSSaJF8hZVN32G8YVmYu7GJvZWmNPSWIx0K+PqThD6ORmsdks45Goh7p4
psvitjr4fdN4ahuzzAPnBXqcBc7DVB+1ICbwuVwDedxR3TnwZPPDGMRmR4Y8SJa9
FBe4lAEeXDYw+X45X/UntOUbz+cAcYg3rxY+nRAKaQ8=
`protect END_PROTECTED
