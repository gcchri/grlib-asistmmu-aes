`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6oZHXzF8BXT1EtT0ttQE9u2zPgBCBwxfuew0Xtfbjzh0ppJscvuenIM3Pd4HMH/b
NYIBNNLTmj6a0TX+rVpaYuWxBkk+lv0SifSYvHXZmJ09prIeQ5sA/qAVRkxIW6UP
FsRATOMMGYNrRZ5I0G6sbbTi/zyuz2uVc/5jbaf63pPLd966sqdOCBcYOpzqUp0H
bKfzBbEbtaJm8ckzyTIJO0TuO9ISHmFBnf92oM7QJDfYCsFUstQw5AOzvPg44CuS
lq3QnwqCOn7KDXCtTUgdpUNyWMs0Wt+ewbu2HTyLu7S+yiuys3N7YmkuxxsW9mok
hNmz7nIj9/KMr43IoY4fog==
`protect END_PROTECTED
