`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TsKpnAcFlcRRj60YerG5KHQoAsFum+qnsIWILyhGwA9VrabRBAYzedo874TdNCoG
SnFwkR/98CSDk3oqp6iSoBsaQYWW/eW/MK0JwHbBCllZV1J/JHuPcqY9WO5QJ1JM
fpjpxYAdqIHkGvU83LxYCH05KhmNwdwvlqTKIk5+BgY11CZ00vV3/pqnsZ/vTpj1
IEJw/K88WMsh+7BAGAVUFGBn9ga+yVEr2zxU6cGuKSz+GiuSyas6IWL6fsi+TL6e
6EUvjhFOH9C7V+tF734xb1HZKxlZd6DJKrCooQgN1ojGzFiiQdZIGlMtLuVlojEg
KUQ2swb4xIKHiySxxY7t7p22jZQmU0AejzOMiAnUL9D2QWjfWhmzlD9DLkuhae9E
O3lJ53GNUF8BvyxHq2y/83wCEzLQ3faUnkFVTb7pW6Xm6HfMLfrK3+4AbcXhBR5E
`protect END_PROTECTED
