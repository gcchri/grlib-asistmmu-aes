`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YjRkXUZsiWwPx9nVNLPryzT+DgEAzCkmHg13uLbSZBbxQOdrEbV4AIIKFKh5Qwl7
C7CiiF01X/63rTXmT5YAOrVieOWz9rqAboGiKvJj7v7HF47KhilQXyx96/HsAcU6
5jvI4GbtXcnjJwn9VHHfmJEQIAwpI25m3i12FHad/XSHOLernO4Ej50jAM1tyJ3R
hU1ITfvJNz64PqOgo1RedPt0/LMmgtOtVYuyOeYBZ3ol4hPbC4+SfnHNYNY+Pk5k
kB8wSCkSrjusc2W1guYxgPSl9IBFSvMuw1NgodqqtETWoH2lD/gRsKPXmUVbV4Et
qUJpAWOfg2+0/GbB4n1JY/i9qtounIlH4eakvV+eaF4LhSZKrZmjvltqh6qDjWBi
6NoZQ9JdQ6roq7xWthfERcbmhRtsYJdpdHFyeyKUP9nWcVTNsB0Qj5y+c9iQoA/e
h4KLEuxxmeGlAEzL8ZdIIWwTtd7FMHr1ugHrjxQJqpCQUAMVPfZ7I/T8U1pIrOo4
OOpRefIFJXKqSMK2QSn4TfvNh9hdhuy+py/V2ee07zP23/XcYoFr1K+eS2I3qqV8
nCt1Bkits9d6DBpnX43DZtOYq8ZTxEAg4DoWU+RKnT0MsdVlgupSXzfhYrbklwjB
Mn6jhZ0wI7BCshyv38irn3mopcDA1v8FNbisM48XX0jpLtKbru9hxPMokWttuxgf
VmDhCufW9P5Gs3od8DHUu8htxPRHKJl61Wt0cixipKtlT+8rasnPRreDwuF69o2U
sS5qNFR6UIwNtDpjHu1OLMUz5nMp30StVTzVNKmXRviL2ygagwDD0Cm84PpHBjV+
PN8kJSO7mOsb37c5Z4zuhg+zsUwcvYT59Faf1u2I/iORLwdiyZG9SFW3uV8c8SXQ
x3fXpHPJrfXlxKoMQFtuTdE/t3UaU+rsMMMh+rCjSeuWtlMXf99CWx5a2z3wBaMR
hwOS2BiWZYCohkYaawsgGGCzpJ09sgFYu6aojK4vZRzwTdAA/9y1lpKt/I9clTCB
E9Vth1FJ5voW1M9NO2SHET1fnT2wsrXBUe6DA+Gwo8cuMrb2gBoaZz6Yxk53UQFn
aI4KWkz0ROvBJZvBYnyJj8cJlJHJXNW88SwxlsjnEppRP6hPdWsVZIOQVqHNr0Nz
dt66gTQvCuN1FdywuqDr2S8p5YJTU5w9+JYrQvwD51R9y7bkUWwSWhbA6QENUFs+
b05XDhK1rZYmNPYxW7tTrN9LWF33Bmi4dLzxGbT6ENSP+DxMCPunhDPv/hCs6f2b
DU2v0W0t+5e1TZp/9Z/unUVDEN/aHR6Tt/8ySmA3BZXVAWXjr0QHYhbsDcp/jOin
ilF+6cJvcdEAgU2u4TyND20cbX/SXvo489YJDU7V3K75Yw1VDAhnaW0/QpqXLtl/
PxcsOgDHRRf/raT6s0ZYJhEJ6zH28rdvFe75X893Ryw1Uvsy89Zl8tutdD9aMv27
1ZIQkdIjBHiT5iH3mrhx0w==
`protect END_PROTECTED
