`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xtzJprMcFjaQQO9ktaIW5bQtp7ojp8HoqcRGp3IlZE9pIM9VOLkKlJhJUG4m/MdJ
lDWipCcQIWUzoeV4s7eFdEKIuyhpy440vPNPkXxVYi+kJi06n0wsz043Dc/womqe
5Ht/AKd3hQ1w6QGkQG3ZIdEfqfk6eEHBAutFiYXFwiz0KR08IlVG86afGFySGuhG
qeoRhysdn5JDglUyXDUGnbIRngBS/flGJtypa5EtxapmYZnY660xJNAxhIXqIroT
EmFDJE+Stpr3nxw5IauYs3t9wD7V11qSY/n6DQVGt+1RwbR56c2uWAok8HbYOiia
stiGWqwAZc+g1101qf+eVG4KA4iRT2PzQpJGBvAIySsg1SQLaK55Cm68TNRPFP0k
WMm44gICFbXao5o1b8LOSk9zEDXYFDmxcQsfU4EIQaFTDMZILwpY5K+bZs7HARPP
Ob9QCj/4x8RvPE/77SCwyfQbkRER1C6OryTa7r+KoLA=
`protect END_PROTECTED
