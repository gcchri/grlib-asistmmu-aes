`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jM9rQ/ZqzrlCWZfp21XbOSsXhEljCUmvrmQDOJ1FuQUXB1ezEWcS/cILIkEa2ZDZ
HCTs6EQxGKwmAs8+VHPseS3oiiqmLvH11sISkydLeCiv8EdJRE8nZCDNSXiiuIb2
y5qeg2AQmWSIRjK2ZMiUzw0xdcUMzgHuqgQoXg2JPrSGYK/spYsGJgpvDeUJTt3r
4EXRIne0bAo8M1O+7zCHyfrjSxnzaLfpk2Swo7SuqRNkUPRBQgiB2X0yPyoNwlxF
Cdyza/dDXUFotydFw/6od77X1iRPkxAvaZofMNDhIgmJNXEm0M7QYt9IgIz1MEX9
tYr64EJKXf9W6FMAEOxG17HLxouSs1pJdHcxgGylizQDOsK7DxXmw/fi2zWZgq+M
1rBfF5AyhAC9FkcrUdRYDDj3dMifrjuPFzFn0H+Z69uJ465iubUOamp4ymlO4Dau
/5k06ChhU36OF/bcioSje0JRhCub3AhtvS/W5I8m/LaZ9LPII4JEemCmSDXFghtQ
WEXAMlMr7lRT3pDjTTp8DDwfZRNS2vFH3R5B+Gse0N1aWXjbYjCxd7v8cWdenwHJ
BlNFvEu/IS7XKBWDc9jytmUZLI6tGCMaex8+hFpUlnFnMeG+bUabR+fkjsn/OM/e
tvZZ1Hlk2tr2qgIesyBV3TPdIo8NshGaOMwcC6DmHSHadSBfOsiOTNZbc0jKgx5R
/sG5g0KWE6dWBDGWih+iUpXO1rq28N98rtWiHvfBIsX9kMGaixps4qcsF6KAJYjE
py/0xueZFJUQpxyqQkrWgtP1Yzegqq86ND5lKDLN106v49o7f/KMvoa4dGp//3kH
n+hUHj8MS7J2TpjjiSv43QdsWMDu/LzWK7lUA7eb+8flm7unvwZfkLT6UCzQFCvm
Hb/rn29UhhKWiLks6v4aH1RYKMmNCTzaIl4yMfhop44ITTFSuz0U5YZZxa7wU9yY
iBFXCPFrJ1O1Bz9YbaxEcZhYajWac6Ti7pMjpeL686TwHFKz4YKaVF4JWPhZFonQ
eJZ06JQz0R8mf/AyuqMHbPHQyWjyssCkrA5DV/+5auEXYwJw07IHItkKE2unnwCn
+GQylRQLJkLAiB3xM52kZ5pHFBcOsZrxIgbE8qhr/5HYiKj+F5yCJyohAGOOOJqd
5cyDIP6lLmSKBjpH9GvQ0GCQ0BrG2ljH8wgcMt8lReYzgO/2RE+dEFIMxYdQcEfH
bJGMBX0Y49qc70wRl0ifRsWBLlli1APd9K9bIinHXSEtdf0osHjh5wWqO8XFog5v
uJTLUXEPAT+igjoU4T0Q7kTXARFFcM2936bGgk2y45w=
`protect END_PROTECTED
