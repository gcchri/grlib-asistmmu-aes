`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HbENCS/oea1dgUIajY9oqbqgrgBRuZeVg084Da8Z4zf6p30UbIeRbjgwnJklfM79
T3c/t/lzxeO1EH7TnRW1M0q1o44IXdJDLbTWr0DrIsXwR+WxEcb119poe8Yn5rMd
2BjAnDjUzS3Peqfj+PYi10Q/Ct0uzPQn3s+yeeFQS3XV4kcb1PjCdol84o3sv8Rv
5SL96jRmN9lWrM8SXpCa+RYaaLTlqV8YXvtLkb96L3f+LPzpmsjHNzBfDW9Lo4A7
PmQ8NUFBHGJ00J7EyzHB+a/FH5g3hgyK5FneKRU5My+81F+0gsux55885Km1bl7u
EgxMtrl2c9yqstUrPaGwMf7QE89g3rv3WcP79e/0S24KdZTkp1qr/E0KT9eJm3Mt
7b9XmN4sRMbCRc+aBJPihbO4dPRV/12V47fJYcRqUKiB38Rp+2+XJwRb/y6mOzyF
`protect END_PROTECTED
