`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BV0AoHieZcBTJtCd+ZmSpI2vIQXdQwMr1CGNTCcq775kn/x5TT6k4IRsqquQz7w6
oNFNt2D/j6Nk6XK3vrn8DCvGCkhPYyE4GQey7f8P0WQOg7JH5ALG111cMPwWkDRn
8BJavP2FC0G0NUAD/4Lt//+/5HKPRVogRTp5SVNenxjudjBlHzStvqPe+gvCEY8C
2Jw3IIxzBQlxJI0W0jMR3d7HrIp/g4uhvuCGlzW+p+XRBpiXf72Q++XtT94TThqf
cIhClegD6MLY+oOnd0bj2jvVZ0yO1tw00p2SGXm/SfTBEXlfEwSszEr5Dub4JzVL
Ohey69xQAPvbw0Ps6eeE8CoZHiyBwIYK9o9+k0Ql2jYXqusa5KvAedhfDyk39LcC
`protect END_PROTECTED
