`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YaJVXaoiHgRyMuOoYcY/xpgKqpsRLiTM2YeksDJlZhuCXD1XqtLQgJ9QBVBswzJ+
zdhV8JiYaqlYXwpCYSJaJOcGESqGCt8xcIrzpxH2fzDIdp3SB5dZzrhI0GmRG+W5
xgogaqIMgyye0zw3O04t+8CwlgxMGUKEp5sllWf63q/Fb73sE46o3tbmH02wbMFa
sYJfgE9TE9+osbBtRQ6TGuX1tvgSeqYddj+hPBpa2paZoPZOC5/pCNhemuxAxUGv
0UyKGUYNaeHWgrGywRRGU4DZV3K9DxF5S1KEBXYsnfRgN9YqdiEXWLXPRuWEqkbL
w0TKsfDHLg7dpD477Cg8upOeXBxwS/9vwRC7VZcQHy+q96ryLidDrDMCALNkStYA
HO8ssdRlNaG6HVrNwx+gcleNq/+VOXPFN8z7cXtidbauzS8KhYhz/SYGfJFmse7j
4oBB0d+qXma9OVndjZU7Ur/UDpCZCy1rccZ/0qhezJtWV2NKlECdnJxsvJVC9USu
`protect END_PROTECTED
