`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W9qpBSnKSdenXPTySdPfXZT+UllLCINDfGFe68Br1QOFCbiZLS34ZEO6SaOGiRJ+
BMtA3eIl+HXNXvUZMGfm/x47AC5X6d5P6MkoxyS/VlQq50d1XOBRFPKYr9dLVcMC
glmNpSGPjjIo5XPxXE45bus07O55Q32oB0J1cLsIPhXBl717LXrxJKttIbneCy9M
bZg8IHMPRwyKJxLd+xR6D6aPsn49hjZOJnngfndJNYtsy8P3VC2Q9UIJfuwddUXu
saUSJMlZhYeT/ObAcmYd8w==
`protect END_PROTECTED
