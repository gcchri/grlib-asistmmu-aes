`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sHNUfRsqg1klDDMP5H5mi1gPIqAFbM9UO8mlK54k6qWGDW8yzMtFLzUPrH9lqlWl
VpI7rhYYuYOm4qmBQXdkFqrOCvJcfmlcbBudpImO+tcJyjNAW7QrrUnqJrq9IICv
VO0KHQwzz6dVJWg/HrDuak1+3zaHzZy6UBzAGQ1IOuvkW2fV5c1D7hCYpXjUlMEe
nbk+ciDyUVVyevPy2ERagrpVO1wCCchBJbcd7FpVpOqDKit21N6v/M7dzoQ9faYb
ze7S+WSERyQQtyrpDxvzOEZBdUJoKSR9IAYsSusi4IhqDFiu++xq5e1Rkae8O4Ap
KQq0yU3Jppsa5RlcTrniR6qYNQ1Bym3XxBPTwtDaJUbn8+ZdqXsAsFOj/sg5T2MT
+xDknH3axUZMqIp4CBUv6+LrCY5dHF5Ac4fuT5nT3NcWrvjalXhGs2mGGlN6gEO8
`protect END_PROTECTED
