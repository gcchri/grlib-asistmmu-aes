`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BxQwbE18f1LLcqYa9V7MPvrzaWae6RFpBrnzn/GrJy2Lya+EkUom9yR3SaA6yvCZ
O6GI8uTK36rYU30sxeOggTrYsRPkLJmx5oSPiSsdM183dwR03DQgP2Io7De4juvj
hVmEVPRON9l2m6IsqXnSg8mvAwh/0om5jgepyRrsT3o9EJQqIrLevVmHuquS/O84
bfMkkeQnE65J1Uarp2GvYqXpQEw5o/PhhZj9SY06rZd2vduEzVwq8HM19nrOmw/o
W60/4vq0swaiS+5crsZ2JrHGlvTa0r9R4sYcaG1cjyAoKfqOzgMnyhVgLmIQ7n8W
1VN6lqiJ8AikAXyT3G/PaDU1h4KLgexSu7R4V/C59JMhV5eWlkehvtd5Z/XCwioa
yIBciVspDXm3JcXpPV6Tmoum+lg6vJCAQ5u5CSd6q+A=
`protect END_PROTECTED
