`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DuMODejjk5sROk/rbSnCkwKTi7l2OO/cWACO09b5F7SEvETc1XkG+K0AXqPn9Qm4
ht42z7V9stQmkk14mrhrzCw/wDLBUVYktwLJyry562vv2nGFBznMn6141KnWiA7a
yiW7ljpAKN+NUhiNNqIa4OcpdX5pAjwJa7sIqPIE4f1X5hASs92ZjcA42DdvOBfj
GHPCMLQ5MqmghULIZz/kv90VMkilfXUbRbIpbUPuf1MBFM2JWzQp1GDiRZ5iXy6k
eRs2U0j8SVAguBpFALAPBYh5uulrJvWgGDA5hNif+MfgIl+LnXjlV2/uyYhq+DeL
8T8uHcMW0SjT94ET+mXID5DhO4kuYEOtazwYjVK81kTGBONVzmOj3k7AAJfFaxQD
L+y2ck+IWy1HrZ6OWzG+xmc9TOGaEKICu17pB75cKtJtNdHpx7kfHIUk1zHYvkXQ
yUmfs+Gzc1ZGh8oPcnNtk290WT5k0lFg1Slj3L1ZZ9PzLgtTpplJ3Q1fB6OaOy6l
za45eD3E9z/zafa/aVI0gM4ibaPIrxuPsuwiRBUTWuuYef1eE3NyEYJKNIo+V2Kt
QEEIwYhawSSRkwPnj5qkJkvQoJ5Wq7W4Zsg69u6Q/NZL2cnKlP9cjAGwxK2B8NPY
KeN1x5oQmTkbuwK4OrY0u+dkCNY5LgNvk7IWHYLdQef6LhjNSS5CyS8RIylL+0nF
4ka0yzxAopt0QQWez7N5RSI4PNzG4nc+8YdvMioU/h6v0f5TGLJ84lH1hwcDDh4c
`protect END_PROTECTED
