`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o/Z1eNoFlINrJ6Xm9f8GiBzmdJNQE2lIh716JsA+aAW1kWvvx/0SydRVlrCC1fpq
KR/3ujyR1MiWZazDwGKrrVRMaHacyLU0fcLM+YMyLSysWPJ9fIXGzz0z7IsR9DlO
WAxP/eWreBKLhVkUrM0UXJSXDdglSxFyeX94S9ACrQkSbQdPGL7/e4am6KNvC5RF
6WAiCbPEsQkDHcGWmicC922Jm0etbW9eVdHGhq6B8rZekKpd+VFGQuT3ciNuVQWT
8RzA/cA2YhionkNgZY711IEnGU9poU0gJ7Us8LGjpAYPEzfXlPhuM5XS5ejpAL9O
z2hGF9jdByQCmmP29eS/pirH9KfbLi5O+87g4I69HmXT6NJOI91BpjQRZeB0lXOG
dbFWMmTOtheS7qQxLF3P/omOdfO135rYzMZd5a7jIYABCD+cvY8FUESxuRXzqbmT
Q+aLm6UFrruZ4I/V8P94x8NGSPMErnTlZmKdYEP/MXs1p7W23xQR/3u5r7lZo/v1
WtMFTVjpo/ZKuW7rR5y/TSE2lMSEYX7HCoCuumLz/XbcN/aucW5Xp115SQHEpW3M
C1IWJU+f1nHLJA33Bqgly7mzYIJniei7hbeRALKSXQoMa+EZibyv/FwKRxLUZAlF
H0uBxRUitgArRc4Y6pFwwjNAC69y7qQklbegZG9w8AKNAHZhQJLWbQRLL3/fRkAW
hNGSBG3zoXczwM+CRi7W6WZ2qif57b+BHKXwFdXPYa2+naLVS2yK27ySwjgBoS8k
eCZTTvZMM1k2RrAbtGS2ZMK0mObhDWRNzugJQTARQmwlPS5jD1fGb7UPrqvR9Ozw
zql4uhbcQg9cdNn8e+se2YTtd3m0avEerhAxQRnJx6kf7JVYKGauEFMZtxrrGv5n
uUFpuzkRJrWmMDqhJUdTMWdBFXCEHXogQUSgpH2PuQt6CbcO97FjZJygMxOYIMnF
+HGgKeBRO8zrnbQvTVtYhg5XVVXYSkChOm8Hn282x1frXnmVDH5XvNrAZfJqKvK0
VK8RyeffsI7tlO9TP3yfjr/ZLsk40QjRrie6CAvnKU7eds1Rgne4Rzepmaiv+In7
kNFF8VkBLO1AiIv/mSfqYAgYKldKqF8JhHOMAin5SjGIufdcs1dFqW/uA227oxSj
+KXywUew0EeP8RAy3dYRV7UDSu8Apv881W6JllGJs2w+2FeM9X1s8LShOzPND0i9
Xz2t46i02rt9Fz9xNlX6wj6mKde+rH9dATrfRBXRx5/Lcj0jvYshC4jX8TtytZu5
/vcX2VhXav77k1sluaPKVYuPfD+3ETa6y3Asbmx5NfNb9ew1morX/FqhbhzH2sw4
VLhGH1HGyoJQmHEANWsbbiIta7jlPY6+SxXzCjCWwdHTE3xzeRyWrIezrbW3Ad+E
Rx+UP7lAgiGYj8dJE+JyhaW17u/OrI6TqWvkvjpDdVF5gzb7PQFQaqzpjFqzz9D2
GqN8Lz982/mzyCnYDdwTFUzq46a7NWnkyiR8EkMekQWlszhbKOiq98eggHhFqelO
zoehHIgg0e2ymPGBd+2vS9stMbNvYV1kFPXK7PpIkzQHbFVEN853dP/q3K7Tn3b7
2cQKzuNXZ+I2BRbcwRBfIjbw1VMGL87P6dNYLYqsi62hk9mdKXdDqKr+jJcwU/Ih
tGGb03fzwO7wJ/orMi8jDcohPUfGZejCZ0BRP8ha+v1rfVJyObCZ27K2/1NE83eg
mlwfI/IbgeeaZ0nnQDsZFT7pPqnLqLrFTJvBpYJYsoQcerDYAXNyrhW9oQlow0e3
`protect END_PROTECTED
