`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KX9yfzP+qOa3P1qEmN5cBifHwGjk4Ahtoa57OTzW5UBLmR4/xW0qi/wkf4BgQKIx
xmCKHykayMjZAnc/q0wnuOKAmL7wpui2juSkQXnE1CaJvR9/DyDuy9LX7Ko0osaT
I36prTOqILhVSgU3hXqytEkszqEFwq40L7aIqL0IJ9USJ83trLZLPno6+0bOfQ/o
WT9L7Pr46TOdjlgJZHsYw4VFcdaNUYYM71M+TLR8oM8Vb3nB9prP1b14Cqw7XBAO
2migKhOeT/rkQRHN5JifurAHxaFHcLtFGnMBZHd89g6shBpQgftXy43jT0BAwNHU
tw/LPvkh13PTaIrl9bZn083/SoPWRcEq8YoPpC9RcjpG/S0EOPau37i2idY8xu1T
AkpthmuzTRyVXCGeRdUOwO4vRX6fnJ16zruj7ICIYO1QyHD/3/A0Ww3c1skTsm5x
8LO6rIklyStNQ0hh9Yqs28sRp74tNqSHS1yd3eMiagM=
`protect END_PROTECTED
