`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jduF1Q6fOSRXgYP5cbXgWDvw9R5zUvuP79m/7Chm6/uy3827HB2c8uKaP8yNnmPe
tshc+djyYBgd1bV8XA7nUo/be4RIGcBYDmw6GZDynjld9OWxU+2txauqPgyB2WfG
Wp/e2SQAmePyKIOcWWa02zppkuld+k+DeULM+4AlDwg3SfBujVkrhf8GiYvCstHj
S1do+mPROZyi07+adZkaHf9jcSm79A/SE6L2LtaVHJDmdHwHZwkxXZHAwZ11d+Er
DmnHo05gAs25KlB9TC/6Q50c9paorVJWh7YE/76OQItI4YCy7E7SJ2634h6a0his
yr9pQvFrpyKWFj4a+59DcKx/Wt11c8qjrWr36INRvOYgb5QkeA6Tkcl5rewsj/Cw
1OJceeigpMMlbRWiDaR7ngsEVsUVnKXfw97kJWdHBN6TGHD8131Yn8tln2RUYA8P
0HWQv/4DAGyX6t72ftkKbHNiWcK77Zv9/dSnKozNIIZYes5uNU1wFzJdZwONzeCS
WkW9GbrLEgEb4tOQSfsxs6THFxcs+QmC/Yv/GtcQpeM=
`protect END_PROTECTED
