`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5EuqLilcKS7+GReLcUGcU1eiuVJ900ADZP1xJpxmq2BKM/vIqDWZGsxSj4eF3huK
ryAyWPuhCIUG73loBiULOf5h9XIYaPSxMzWCLtyL9TaXfDL1WDHwWcoseJnEytEh
O+2wVUUaYld3Pz5vPOCAiXVf4EF+ImU+YOFLNGYjLJ6JbGakPmB2aCwu6Tzwb0GN
Kvvs6oHyeyrXwpkpD0eb3rVd6Mh3jUVpunxvkMQoY+6x5Hzj2IHh9TEIGtk98+Sb
IWDEfpUUsbljs+y/YvdudvUZg+ZYYf+cHf5LaHZXtW66BB1hQy6dCE/A0D0VU92m
RXD7zCy2nPOIYi5CyfjuZvB9+XUbtJueXLA1WexRyR3K8wS5NCILpAH8amUjGY9l
IbzpCQJbP2WkDTNrSYSsdaEhodXY8usQzJ0FNxO8AG2Lk/t5l1aHztAYb/erKiw3
8GfU3fBGINgLS55I+LzW2dde/5te/MMzHXp/kdRIdOU4dsMdSRj2flbCPnfvJnUO
BU3tQnjyG3JVshbl1QDwp1gSaONegvwAzQ0dwU5Z56IbotE2uwdpg4J3HaHetW5D
MgpqyNpoNnaRbtD3vx5iP5Yj28BqxffjUybazsSZXDJCKGMOC/muqJKve8Ivz+CW
1xfkH7UgM65QRGnOb41v6ambP4BLxWO8kJ6pIKdarOB+EJsZdpafJe6aHTQqfhtQ
SagJq3BeLXAE9ulvMMXGN1lhlcUohvrELinpYzcGptsI3lNB0YygW6yBbI+x0VWU
HOLVCXva+Ec/PPZRNK32ueuU4n96+cUbLq6phTtkp+25fglIZ2Iz3cmF2tUtaJmB
yviytATriFSCF2KkR2JTSezeuvLCajvm9R+a30ej8Sm+UmPKEl9KpTBRr8K9PQku
QNB8K1R2fqi2gTKGY73xla08k0UmxCte6cOVNCOt12+CP4Vc58IIVTy/3QCsE4M/
6WQgq0r8qwLWqglUlUxlHTGoBt/by+cwGa5ArsOWloronQJHCGaQWcPl42oAXjEe
/YnIXqBJ3qj0NCIyUhN6GAuiWCJG2NJcgiJTjcQfFpjpkP/ANM5tzvWAmku8IuRs
GOo/yB9TMH7gwIhZHBj1PXc3sB3nscspWGxfz4w7LE6ILsbSmMBvQwiV9jO18SDy
7jragrapRHvo4k3qUw5A0cHxIEVdvhwLvv/G/0fZf9DQDjqoVd8C02V8ILGhkFe/
WRgGv4VZoHegys3hbDZ24uqMTAhmrIYuU8T/STPO09NbN3M42cdgK1a3EUgkJXca
nxPw3IDiWBVzxK5INTXvwntBKQ2YmEsmdLKSlUeYOo0J8mPciXyqXHcIeC6lim+S
+swLOLUoacGQ9wGhaVkgu8caPpUEvgOL9leSdDVSL/vBeI+mJB6K0Y8XTKeKABXh
l4YmrJ1tjtHyelCgw79hm5Oibrf3TNCfIfMYTlApMWQS1TcjJxY2R9e+HRL7M1EF
YrA1sY7wrxTEuIDtbZd8IjfgOzv5jTf2kB2uFXXK1YJ7q2A2GwMgPPYNuT7d1/zn
90lH9B0XCFWvfINKeoNP6axYBAbL8nqdd+SsKySboHKgfyOwDNx/lWJHFvfDSwrm
RFZjsh0fLWokR1+e7qf4oefBS5TPCpnk5/07PAMO34/M+wwJBeu4E+VECCu+7war
2t1xtwtAmtQPIlNfTClxdwixtGIlcs5zV/Pie6i5oSUHxU7uf+bK9odT7tqNchKi
FOYtkrwOUU1tmcaydv3/IYs4iaJva36PVkMGwtj1m2il0M8FTuqDII5ABqLLsEfj
sCpPzUXzIIm9BeKzUUvDMCX5Cw8aGBBZz8JFeJg1fthxj47rvlTIily+SRZc7eMQ
DK7X13i1ctTJEARZehFr+D+zaI/CEuc13BT5lmK8LbiPyhjfyztmVNMYw1RnKyts
wORGoIrWJwEOuJmxmoq0pTR5BAVbVaVz6Rr22UmJY+K17PBQ1x9jCso3R4WW1kBW
WexE85eyd0tceP3xnRCZ5uefONBBh2SLKOaIxkSPqcUgo4FIh2cSszlN29NBPQl3
/BtUcb5AnREKN86hl//Oqo+TnaYBQQ6pho6L4xHolv2ZNHyEDoJnrSHZsqfWaMI+
WK0GwELWuj7hZw/5pXTnWzjXy6HSN7l+S6sweUxGNxKPlH7o7z3FrTaonKgRAbJi
DfGuloLrKAJ6JBkxoIRhyoD9eO529i+ABEx8Ts0dKVUQG6iAbNRg2G6umnZBTnkB
Gv1Jyg4MvGDBbv9pQMWR3vuwF64jbRO/oc+IOM0DHSMv0/GiXpIZzI/EAjUyfj0/
dFF9oJwy0UbwcV6O6/QIJCy+W/9ZbOHS95v3v4qUjpfTjMWarMwBFqKUf5+hkbpx
s9qEeAAfvAfT7EEi1a2peIt0T9Mqk3hCugybQjl+bC32+6AdtP/tDwmmXPYfa5sy
Twbx3+8O2tVhu3mZhlqcZHevXiOPdQZRZDUfV30ke/N2cQSMnmg2liSuU0g2YIks
vT/nbvPGWQMMTJBoCKGPyBIGsYZjKJb/MQhJSDJ7UTTAl/g+BNBzD0uBIoKBjaue
nnGONhhm+vFcEl+hzf+T8ef60Y3iilwQqXszyZRaMtRoXBy5RKUu6Y1TSfXMGm4V
sDWhZu8vYs6AQVAL5/DwurTwKRYAOYNa3iMcahL+R2HUfsU1pwuchGAuVI4Rqlf1
BZU4y/roHvKXzSBsxlzPjPYa3Ytnk0izBdRo13lywFsiWRK/zPnTFFEG0BiWJ74E
bDA8Jb09dlp13hCCE4lC2pxKAD21eUuX3TkUNk1HaGN13T7G4DXDfa9a53HYV20Z
ndPjgYidinPlqF8NV1Pj2VnqyRgpNZJgPC8V0c3xyGXt9wI36Pq4SQLZPC/7Q62D
VZWE28gMjQm9SJhCrHPEJlkEnjLJKurzl31YA/wcTcLCvDqerSHiHDQG8ueuWRHd
yD5x0Fd/KsNHSpYZyu6Nx8VdlcEktzRtVSZ6sHl3WwRC5UN2CJIoW4hzhPSpJXl0
iOswEzE3WrTc1HHhZcO1sDYJ5mGEsvvDrYVel7XbXL65fjxCxti0E4zd+cAGcOep
ZyzDnxONxQtcxVduqDuBmzn6KZu+b6dkPOVNzIMLnL2o8CwfNBCgVHCGxIm/tJ56
HMncl9FeHuYhpSdKds/Vqn84CGnkTqeEckDFjKLTgOI3VtP67t+MtEJB7LktKmD0
7mJdFVPTC08KXpmb2x4ikBxQ9dcr4HcPeCdNqmth3JJlI0r1uXw/dhJ7CfJ004t6
y0cUlflPO3JXQer55v711+S4Mpoys0+b4rjjWK1QCJ8Xd6Y08PWB2cQi2B4yhR/S
WVxTZShbQwBO9MVdSNIJpobsQbc65JQvuXXawtE3SkvYywYh7pbPv3ER2Tudy9s4
wxXaK/bOSkzRhVv5Vmm1rNMxdywefKRLMkTseG72kHzPrFucLBnm4jc8PC7B6DU5
vTmrVeLCZr/bfce9WLfnWSADMQDJQsbpNhQW0QSmmODMamX1ZNyjjBCUKgv8SZYA
WmQPkeWD4kXINUPhZ9h/BjkHvXp7orhnVNEPmLY6USJEenCZHqfSZ2xikwGDFgJE
f00SOzWJSz+bWB5dk7qXb0GaYjQkqzIsKSQNCEz/rPnuN/bCrnHIjthBm5mXlTU6
BnHviS8bUtfCdSIzAw8VvZb+XHT5dDoXQi+3hNxxDSi4/pNKYhLlzUns073mVvE6
S1PIY8Hyyy7U3xipCTyxV1m47UldL6REq/2KFwcmKZKadZ7VM803L3JKMo3CY+Qs
trEXbs4dW1dKZJzZH98vwEWam5oXhwoX6xChTaws0+Pm+60IUVpczYjLZGB8dAEC
FEwidsQ6iycoIGjgG84sCswMDP5ZENNH04bvTRR3KG+vIOnZd/iSH0hVw86+SgaL
tFt0BKRiriH2zWcHAiBK7P+ykNPJ28ernNVvmdgUaQpRBnxcvb+BQubJgbj0wxcu
ziGpoJFXcOjJWpMf+rERk1ZXX8skTJW/H0pzl4ixbPLjE671e3dHxWVP3MSTIFeE
Vg4aNk9bdkzLYXbU2Y48ZZipXuwszxB17gQk4VHAVpzIdwDNHXr+2rygWD5qn6y8
KYedTmQ/771dc/etv+NbWMwxMQnQ2QOUUT0xy59IDe6qN+S97Q/umzYZMFrELgP5
yAe2bvaT48+AFizBhZdDHhtJm2ZlYWD86dRRiaiFav9FSc6KmeuktEWRJ06b3kos
bCkVY2JFh35pQUebodwKROpTPd0QrZh84QnQCye/vYfZLeGKwMBKxQ4evwThge1H
UD0Hif8Z+pPQtxR79chvCJ6skt51TZArTk4XXA7dkVCHe05xmFcJ3QtqaKwnlP9d
cDyaGCGWSloCSJvox6yalLLXlzPY1Pt6sT1993SUJBPkHje5xkqM90+gkN2pCsgU
mVgqb0adk3Oj0UXV1QsyQY9+sI/NIMC4BLSdDfDRyDPA90Xv4E2BHKU//oyh6pWU
mVDXlIBzFfl3xgNgwkBy5VAXwaluYyOdQR+2zv1f6U5ktt5E9rj3iauY80lcsdRU
mmgV8NmdzoRNbYmH9S5VzjSAWYsWvVC6Pw2AvW4j7qpHzvR2FpNCnZjJZfyG+sni
A7JfwIAboczyjPVotekD/wWDxzA1eyfNZdhz0Db8f0+q6dXTAvpkqtPICNirHYX/
OXcKUgOrdI6wbVpGdB/UjyJ1by7670WJOlVt4oUhr9ycynXTmjhj2jimSi8Vx2bn
iJsvkXO2ieIXVxAUq0dE2ojv4HuxndzeJGMMYh6V91Bn/MgDGG/Du8AJxR8aeyOO
csHeUvv3h8CYzUOvtahdiP2mBmSs4E1I6Y9JFI0guxhZCho1DYWOLW9kXj5UechU
eHNI7f77fqIfco0diIL0pYQ1Zbib1c1sxZUH604iNBnaNqkm6EUleSROzYJKREXf
aMTTm56fhFKsZ3Jmq6QDlu3rne57mBRdcGNWADY7DOvL9zB8zcbTSp/ewEwyafpj
Q8l1hoyHbK7OEgJbPdAZBAYeNgDkRyxA3zFDPgr42gmBG9qgW01ezMMbBam0Hy4d
ThcR3owmS281QwKSfmfIc7nZA4JNl743Yg3zcWJX+dTAQyeEwV0T2nTkc7/BtftA
wt06+EMg+mvgHN6DY9cpi5p9Nch3/MvdXC9Pv/S72Lv6bEt/mQa52WT2pCsh6W6V
q7uTMmszu3/IGyVcrMQSYi9bMCu5n/4hSra3ELoZty04ekWqZnS+omyx7gM1kBxb
DjFz5uhma2INbMpKRpFon0fSfZKSCOT3NKvlWFv5CxxcKv4m1Q8qK8mHLy0MoRTu
GTlYcC3XNWjWbKM/KigOxMOLby6MKDN32BlBu8/Vp+vO/6i1V5Q1nfxt60kemMK2
0FNoKWgqrs0Oo2firoTX6Oyd9l9oEYDru8pnpiXM19lOjG0wouCUT3g2TbP6zc0Z
PehvH23ylv9e5EhtcasPQ3fH6D+u6a7V9d9qcB4746TD8U+ENXJZgCr8BvOQq4yk
M3x0iR5pB0nFNAiOmglxyyR03qlDh5y59D2mBR/2Tq0GpXocIYG1SHzKYxb+MwTm
EWrpfLSlUpFlQEJu8JKZtC+TFlCaUHs2yukLN2dvwKpbSiMJlTbX87wg9P4fgjGc
6csd86TocA/UuyVV/KRHfb9voydtTFM4C+ys78RrHO1HRrBKceyHFkCTjdiYlI6Y
zUHBc5cxTRBA/OZvdf22F7XaUZ73A5C/0zzLMpIcRXZzF5ayB7QnQjuNHOr+oI8r
IVnpzvOw6fFfFIArEgWzrah7hsoOwyCAwKmd3b/IAsiAtb5tlyUt80RKRvXOD4YS
rbEh8o3jvwXdlnWn7iixB/R3pO2lvAm/Szwpdqg7MzpQaxAD3hOkPcMUpDmq/n+u
B9mKA+gDJzs6aiSoyAueCYEtivGh8HUC6GZAkTkQtcUmusrtI9TBkrNRwGM5jqfT
0ma9yI150o+7Zwfa8NgtDnh69J5mRzTNgwDbXqA4At2B7r+LqBv+e1WhkAp1KWC+
88NvhsvyW8jU5xYzy3u3VR9IoP8tzECzTRHnujxEsjjMM5MtVCaXea13YJWnQIZD
dECvCshE8uwmHmnjB/WW3GNilndGKGtMv/KvIDxgyG4twjqaFzsHi58O8KrDQCGL
H9n5CNPYBsdt5hAX6NwSjrbBCgONV8c4LE6Z5xvID/82OllbTuOm2U8Han2ZWK9A
czz6/ss0xna5r1eEt5oT1W6BUp3fQyMuJkvaX6X0gzsDcUOb8OT1M+SCbO6ocS7o
TA3TSbdqoroa5zVnH3g4Byoipdzn4G5W/kMS4rnC1aMXghf0JjukZMyh0Uuo/ovv
bNqq+RBobApXxcMa5dxb6MgLWjFu/CjYZciRX5UdR8aXp3lOJf0PCfqhoCVW8LPx
yP5XbpzyQvyF6gm9QQU6S4kQzHzZg+rTMbcAg7tcNMfs/GtYp+Hif3eUYXKDPm0J
6wj6qX/+qJZ4mtDPO7jPdpWo/HPHr7pJRfxDU4YwmDqH9k/wso2UkIRQdrp0ajDz
fEOCJEEA2+p1ZUpwK9QfbYIT1z4yqEarhgiL4BERORTLXRgNA5Cquf+aRs7H5Bft
DI9/T1fEw/YZuV+IOvM9y8qHIKBoEl6Wm2qB5EOq7+zPoHHcSscU4Slpti2k3W1o
ZG/rOBvYVwU6pqvqcnGNnUl3amjiVOpRrw++MfR0CTlPhEM8o4RuGcn1EIXhSs0Q
xcUcrUP2FVOGfchV9AFD4ltqLNxQELTOHUMoKWI9gdEqqXqnwM4A+XBldF10dFDr
zjgKdpRJLbD/FFpBLo6auDJ/OHhq+EUwxo95pdodiIddveIjuX99toTSwQUaz0h0
NHO0XlwVDK59EbJbnX7E9mYhGoSjP7xHdmjWmveHLuamBNCA7J7UK23qDF+TJgWp
BYXfgnY3FiAqmDsgNo/9puENoQ/H1fHeaIyWrxjj92pGGphuG5GJ4y75+ZSsyfGx
2M3lel0CFg8l7l10hScV5IVpMsDtlgGF/maAQ7cmfz1jJwLsDKLVaVtcK5E4XWmU
nJ+jB5DaNGA5KE89GNo+R5SjzKxB/SSD3Kqsc8+4BKD4jMye5z2zJ5aVGDKdjxg4
BAooZ50r9hOnz3dZ4x4D8msX34R0IIswf40vfAyH9KEroRvlFfZ6D4r67LpPIOso
NJdKvt8vvvtFw8lMCR86l4TntvORflWDtnUKOy4fkujw+OHQj2TEg3opU96C73Jj
qiUxmxy0oApLXCcZKMltzdbwfzHmZCQ0gHIJvEKUkQlfmPHH0UjQFLWM+7IQdObg
LEyC58N04vzQSpXoI23G32M3fVDQTlDS6oqufi8A42ojxJwJQ3fwG2i85z7t86cz
l4fpQtlvd1Yk9gsnZXGHC/gI2uDHQ8GQ3dajSTrl6qFMznY1nsHVIVoLgvBece+R
Hvwv1WZJH7mAov67IC4Fo9JV7QOx/U0kmzd6NTKa1/4LtxU71SD/DzWcGeWSoSMx
o6YKt4SxUbzys4DZrtRRhoRRSq9GsyXtCGwxUmmqAtljg4DxDGPcIy9UVB90MbMT
0ifqSxOcgKc6yvAq1NiH3UZndOAuw48aGiu/sLH5QrJf19ojHOlFFEk0uLHlMkjA
bvoBLaG1jMjPVWBQ6+jhTwfd2auih425GA/Krj8Aa2qTU9RuISmnImimHgCivo1J
rmqShCIvzm2qNUS4JDNJlbXMHsJMnyWi5Lo4BtJkfFkR/5677kRX4jA7fb1qgU8k
sodqXlwoQdTvRJwMA+ct/BLMO5ibSPjeq2ckcTChjCrRqj46IORpQMFRJEp2OFsi
/EDJdDDd4s+WWQdwHuazPZoHnKx1SFGMvlHiciTNKhZ7zk2e91SyQ0kHvyZTmnvA
FT7gWa1JJ2aczlDYtAhRxQ2EQdDTwBdxuBloARQbF9RUQ3ZGfssYmrYsqRNRZmV7
pjwjAh5GDPlE2Q2mrw+7VwrvxFddrgKpIPkwPBwOZqMpXrGA6Y9VBbbFbk89tC7M
E0m3i/9+GXR8vBB07HrnvDv4UBvU17Gj18x7gNM5GNyR9QBsITYat6QHuCj85Oo+
+NlLNFPJUClJ3J95AId2S+f2tfP7y48+EoEmcXyRqCbncxo0S9zdnbEG4iyV83vO
ihRVLsEh/+rI1rPm2CEhQTygwcdwt1oglks8RtpAKLwxU4hoFA1IUjzmtnhQEkJD
8vM1D2BhB+7FoGTfNRl5SP+ZK5XkOG4RcTZ5IEVKX5nnUDsqJkMygjmKE1OhZQim
p63+GqMr3vN6mmoSUVDZR6HwPl16iyq7lwRFoRXXIdG/3xqDzH3CCJOBrY6sxvbF
YXuIfeE6yv1Y9WuM1ENij16Mc71W7zvVCjWROUfXK4J/lJbJmargpLfNfmyudPmu
XlQbVqhzyt3vW5B1ijiRDzng5GpR29/43huKNjv4MhZ73yH3CGQsiiuwFLOEjTpC
HXV82rUEUUQyweYQo3+ZyZF60q1WxXSGxGMOX8tSRQALNMW3iMeQc7VRs8HXshtZ
1WaDbmENrI+s+oK1+8KlPZVlL6wbl57pudDAmeGJv3Pi5uIrFg7WUKE4qW0KIp/t
B4JiHghBWXsRm8D/gUQkasWoTKaKN36uqWPd0ycxOLXB+hLV0+WWLLcMQ7C/Qmtw
m+e7JMqIH4Kl9DXYPIZ07W7yrFCX3BGi/WV37K0Qfbl4kFB497g8jESTprXBtFm9
N+gE9y7iA+2/ir/+eChQd18ZUerUDw+W5+NdBZ/z6pOO/yRQq0Vul8u4FEGAgoyC
zWmLdRNN7nsChgo/lJrmm65+2gUKijCuY+eXHuNmAyYIhHE/CCl6yXESQVJGpXc+
KP/+kQLwSo3M/yVhL8o9CQ2iEX3QxgPbGK06jTZGdPyjIG0n9xBWnVCkT/1Aa99Y
K5QhKrwSCK6o92HqsxwXpN4rd0N4Nr3OpfGMjvYUty62u9Gco48m+xzeO1++6s/4
nOkrI/1qMxW4NSqmKcrYuszj4pURJAuPlknGnDFeC/mTa22FLbMd6ZfOtbA52QLD
HTlSOd7buVd3LOE3I8zB9u0gnZTgvDYdjwfX8qjZ0Tkv2JMAfg4cm1R0sk5mesbU
UzNC4xr03kMCrWHuVRSoVa91El5ob+W8JT7jd3zNlm9uUG6TxJAoTRF9OFbmim1N
9ugQ5wovzZeoCDqLiSywMI+M891xGbxBWd1gPPAWJcPwxqAmkt7fSlPWWglVEJ1I
j2FjgG8+22R5DkCLJ51EVTc6ahW9q5Sq7hVYytbjfaOMLUbS4YbfXzpQRTYmwaCx
9MKECxxHGwbtirSbP4W+20XYs7pTqT2Rl2V4aH3tn0ySfj6IY0TIKHaN3SZ7QIi3
LgJuK3CoNoowR9nCbfcdSZwcWN1l+vwm+8sEvS3WTfC6zUrYbFYZUs5gaEEe+btx
4I+eVKVd5x3kYxM2EjNzPxqmsHq98M8rImy4Aa3+wudvtLbiTy2SFoNaUT3ez6TF
kcr4yHHU22rXNSB/cr0p+nAi787wGs4Xkn+9ZffiC8GoiKxz0rlMMyoRfOvgIlP8
zfOS5c2mCjvZ4bBVSTy4bTOaMu3s4SESftu2DDZY+Ly0LogkOpY0Q9lIpt6dBhdJ
kGAcCy2/JDv4f8nuhatrtmvakXQETIiAXCVAkeGRyksgML5jFVK9J2VidkqxWG82
ov+FmvMw3VHbiUX6TBquR/+3z52gdd7n6ceKfWSJsIX2v3qQAmTPRB0LI5aq6Rtr
3rDjNRuM+7H29RVys4Aj+Sb2hfqm76TtjwY7zH/8ukM/vUrF3qwYY7Qk2TqTvGdk
gQbXdi6vvAbkBeGrSRDDzuaCKmmfl7h5WF5QDSBDgXPxUThU9c1zs4jv4s18EMFS
4i4YwxZeJrJVe9oWwM0RI09BmVHps14dahsCJMb/BcXPyD65KIcZ5Dfg6dvFJ2Aw
vi/cBqkGzMQ5qFhAEp8h1eVIrxvlGTmxOxX+WNSo1Jm5Og9/NOJb87b+m8X2ifmK
YuANB+ws16CeNcxRjfb/A7s1KP/3PphCvoS1b3rjc1Mnk1XvjONTr8m9y6ZJwrT+
ZKRllZRMNUW9ocGl48fi9XM+//PxQtLXpjdEYHgO5I1MNdOyIkLL82jVkzYbOiio
f3j8Pq7vjd3nR3YNh7jR5tkKCmaCYN2k6kqNCDLOCpfYWh5N6HshZk7ey/BuAGIC
UCfxAO9068HfIojiMQs5LozTPf2j+bBgNC3JO3jmLexGXrKaJeueQLtj4fEkypos
iGmQdqm2mzp7KLhm/18ix0Uqzm83jdgl3i/n55dkyPs04StixIElKu5tsYqfCwRj
2ls8aUQHpdtNo1baujtaEnDyjyfhnKmG9iG373vCKDn6PV1v2zwt7FMma/fpQ2sV
+h7z0H8ruoaODd7FVD1/S5U3WBaPwBKg2ulugbD5MwI8VDC+7V4fQizTIYOb8crb
AgtF/8/JXay1YPVgPQLhk15qJ/P9MlwBFNKlhLsdiHFbix7ujZK9LDA8lOL7ZPpx
k0Jp2QNcGYrUzZNrOv5BCdiX69ZaK1MaVmuFURxwDxKskHOkyhZboAkPQ8yr33sj
lGJHRIDgd8H/wi1dQQpvJ20VpRxO+B2RYl+kFZY7RisH+J4yd8p92AocX3JWqlf/
CtwJuJnrQkOGuX6Zk6ZhvRKHm2VdtwhDa3holLKQTIo8QXdaZJ5XG8QGs1W3dU93
W1cNX+qm0hSrGp8AYppmaUx2TZBEE83gVW3cFphsOZIyWE+cOnMORpms6SD5cw1L
oJskfJ4NrUP8tiqhXYIQ6/fZ5G35osyl6HQnx3yKTyLkPrL22TtnwviQBdDEnJH8
xD64PzVmRIQsUZ/EBLA+p759Asf3WU9BiZIatSfF5gp+veTcAEDHNCIOnIBMxdnS
FJRRA1k9VLe3596ZeZyaHzPu10UxIlGD1PGV/L1c9JOK1Aqfku1IOjYXFhjwszf5
DucN/VYyT0Rp/WFUSxDxcip0y3Hd+RAEN5YDzr/eLUzJXDBiLzfYxkDZnPcI87SG
kWjO73mNGi0h6ROjrVED/tG3Zzps18HLhSeVbDcIsH4nH1ePohKdNYzGWKnLiD1I
XEJdznMZBp51kac5lx9vs/3jAm9ZNIartarV7OjR3LycRHg1mXnlltyvfQTAtv9H
Iomd/DKR22casCukHYE98Oo5eJve7nSFAJBEAkHoywPLKZnhSqX/13+u9+ixDwDk
TOX6oVhZH3kfXUjxFbrB9oqBtVvt3NcsZCO4x2tBzVwATWWrOd7JIk6kwsDDF364
edjwjrXUZNG4eTkMOaJxIi1ScOrH++7wPX/zjGwMn60bW0WPtfkGwC8r45C0RS6X
1FFTGivusPf+cNgVB2rvVV5FDvA2oyBpk/vo9J9ypeheLmbTirTEVvvjWgY+aJaG
gQuieVe7rwVv+kyniTrOjJ/YggZHxH7EvcrxChiFefCLWAu/0wDAm1JwMVQd9O2i
jdmVNJx3G0J0hDPpA9h/JyhwAWzwsOpY6cOEd15JVdC1t+EL1tFic33b/ZbBq5K7
tXJo7vURV3rcqe98v5dsLAXDUc0EeBXE88fkPtKNUYNcB24qdNwuzh9zsbt7aLHR
fyJl+gidY7HNigdPsMOifaYLUH1qKLzfWiW1ASMOicbskbEOfGeIetyYL5f7cKKd
ZyTjB2jCBZ9YwaIujioBSKgq8LVxnijnKqckmpjmNtePQLTctMMFXsrKEOwjJvDF
sI6nap3Fu1Z8o7IQ2faNodD0WROqtmiKSRo4ie2QAc5eYh6selVtt8Zq3S+cFkB3
quUBSRGEsFlN3169wWe5XrGSP/3aDaPyteGYzLBfxx1VRddTGFM6CF4xtigzSYJq
TEZizqyhwsSRJHSrqGfU5q6LGrhBrqufe+R6J6c+Xy3T//tjrQa87OcB7vu0uPDd
HLE+A0LAl2SvhEjgqwuZtraypsQ/CO9/vO0rbkSWgHjU4gsH2ogqjRCtYmSIQZFR
VlPNjkHE8RYf4I0sebIU77S5UIULp7k2XAfqbusP9/BmICVXC1oVoOlbjEV4NGC+
SutBSvgFo9436hxpoO7qmXR9lAXQ0fUC2CTslAKcTvqKuU/XGeQKE5ZJgUcpqQH1
TH2/m3x1ZbpZCJYfUBHrZftIXWYiUUBKVZBiKvIbm4sf30gHo/TFDCIMrs+ncLAT
eZIXna2I4I2qHHeiPvGlAhTXuCnhehpfYpjzXnd8F5p/UbFeZsLiqf0X+uJ/rNRI
2dgppe3YTYQmg6Hp1UliYOwY9QNRZ9ezk81Hvzw/Q3xz33sKp36T9UF4aloMm2DI
lECKr8D2Ge9SPWMCmuhUw+kl0lYw6hY9eRHsDo7Jz4+Yy6IjMOg0hmn6b7D2dUbJ
gcUKt0T1yIFGqmayLmJhiRKCAH3C2YmmmHj49oaQ9InM8lgm/l27PzVeZl5e+3jZ
wfOuKoumE8lyJtRHsDxf3Q9M8gbPYBPRYFZE2dMACL2zop8NCv01nE/48KF80Qgk
lJ+AwXSQkMTJOOaTRJQcno5nld+ZuxPG2Wf98B+DKx4djAhLr1oV4it+NIxZSCj5
R0JcjQcKICJyKpJwHeVXDeA5Ajs7+fmLRE88TKKUYMwH1k5iBHHkDnM7YRqLm+jp
vvajRQMg3UX255YmPN2QW6QJ8LzRdCpn+jQdvtU6qKqE4untM6RGCpbwLTndVJK6
GRtn+TNN4jGQeCjsSr+Xi8tsbEbncePGKxzmLwQ7OfvJZ+/uV+cG+ltce6yFD82m
JlUdKVF0IU2cubHx601KAWrXBECakQtjM0iYY5a5zju9xkkgPGS3QOyh4kIcHyum
ecIdFhkvhljeBuxoNTcm8ffmkPcaoF2UViyoAeLQTVy6a0PrxZ7SgvQDnrMrOmya
U9Nnpg8GLFWhQqZmp4PYxMPR+J/zm6Y6dUQfHSNklKdNIHmicVjBOsRx6z16S+m8
8SteDrREaRp5lOhE3qrLHNyjW94HZo+iycjfdL84dS0Z6LPwJnbNnGXtPzq5ENCT
JXSbWxdQgQ5xmjyMz9PbERPQt9f/SpL2FET0QOKoPFvwM30lucMIM2P1L4zWjSYz
IPrnMyEG1r7A6+uhD7m/xkA1Dfc90w7JnJvcZHM83+vR2dw/3eVx+bZ/PYxInIp0
5BDM/Et+IkEZbR71BzFQGOcyhboVHF8dcWhEDiVChj9CuG1wQURom4jXCrh2XYI9
TdNSzB5a2KDdeYCbxrB7ogvo2JVWv4cn9EU5RzbNlADnpYpHY+kk/wtakM6xkfXh
vCjtIXOu2ib1LOta+RWapqglMmFZBU7slLM47Op8tcjtC0JqXfnz049B/JXAkHJ0
QY5yeMVDsBHzDzTMJ/TjymKhwBs9JiCz0GW1sZOffQi2KVTivuWnW5860ovJbYId
Q6+ibBS891xniwsEQzg6Qvo+uzi4TrlupCW1S40lKu145ftNHK2RO6fm1DIq/9KP
q0GbtRMp+AT9S8UEQPKkuLqKsGnMAvjuv3yQzb23k8m6/IYiwi2It+V6CB2uHyEi
ybJoKB2QgGw2CP7s59NcbCW4J1Un/yJtle0rd5rcBUg2v5Ll1w92B18iTFXnJAlQ
KxZJYDy+LYYLXH+FmR+hya1Mnpfac7+iwB5LwukuU2P636t/vNSjqXM0sF+X7uDK
A1etfo+sMxfJ7ac/h/oXbhrDjuCkUY5aXlE8s3pKWihBjtXJsOOdIqMaULuG9af+
9+iYBXvUE4dcHq99c+l985zKc3Szi9yO48GbINFIWXwRtzVjlA1UUWzYvzlBGT81
0hxAAh6tNb+4FDEcrs5r2+1p0UldJwC15ErHW3B5Ita/2zacvReb0wDuoTsByzNR
h7kRMIyVJtWG/FqKA6N7KZQwNJlXr83DJ5pSJsWxJasjcI6F7hLo+XikxkvpKZ+d
oYten6yZo2bl+XorU0tK9J++p4FLmNvRZndaeXyrq/h5uHxq06J4EpKUH9w1mESQ
s8f8NxxZGH2yWUXS4IW7R1GaZIq7Fe5SoyVeANSYcT1WvhEu9wTfJyL676CLhLBF
c/6Es6RqC//AF4oMm7+i5ZtyYXJJ66cILDHPHkFeYo1Cn9XiAfMds/bMsUPM8/yr
ZCWQ+7op/BcHdhGTggybUqmTKdIQWWE6Sq2pPCFCd1C2pbdH9pfFUcK0SIkBcncw
pY/+yNhPpl/5cj93obHl8vdJDCfiVFPwhVymge6xsLG2MH9JHk8jV13DHkaYYDWw
AvEOAfqstqjfsHLApAJ2dBbWNwPZzRNnNOu3L3ItfyJsWcYow0DVZBsx5cTejn1V
xcsNDLhNh5Q8ughaBj3jHr3VtRIVIabzk6i3b+tYV7ywSYTlcPWcsMNWUvJJYz9Z
uvm6IXP1VbviWrmUfxLlO8LIlwhbuKkAtV0R1wlK/1VN62LRZq7mS+xFzdrE9eWt
qV731px/EpoplDq3KQeWY07WlliGAaqvydqPbxbL7T4kkV3k7SCJIkX09MMcVgOq
4Zb8n1LUnjBsyLYLIFejaAzA5naweh6wA+aydUmm9oaw0/Cgq6tYWYo9leV3xu4M
lHuJC0aFLCe1+yKy4rbt4B/c2AflBTuK5Z85vTA9pd0zk5u4+H1nUPw400CPONti
AyzsY79LWgjQEfyyKo3WqqYqdA/CRfboORl1pbCABZuM9+8THRflKXZzfVrzqX1N
k1C+l9Hau/D3Rr7i4rB6cbQBBmRn28aJzxLC++Kd2RkmQUabufmDY2156go0FyiF
MHS+Vs8gN/oSmK6OBi4cFNoi03LRIchcZUWOGq1TyfofqtMlZO38nzRXzayHjsj+
Mnya735YDQ7QS64MUZHzlHHVwQ5sCZI/PKDYIxFIeJFT8nKBuVpn+y+ibXXKTthj
c4PK8qf5wr12o0va7N6C0ggORNBuL6WP9t9nrTDxicqreehFiISWTSeBlwSYCMUQ
JmC62v09USTPSoZcOHegXr0ep1OYdtgOuYKfiFcr2fQlC06sJgFclRSYKzdJTrkM
m30Lqe3rZfWE4ekoS8X9PFRgYBMS23xMtvVXMti/f1Y3kNTvYykzwbd3rvVCJBRk
0zWihSpBaB8BLmsLu9RvIc/HE2CH9K3FOR3glP2KOUcr8of0+XtTrzLwue/oXxHK
vovTYgTkkji9/wJglqg28mLdh4kU4e/LegGC0ym752Kbotvlln9aVoxNMw2AtOkm
qADLtxMlphlHVfBdmHTXY/eI8Ist9eTXAkW79Bi4dKuPBRJAHApodh4nRSBGToo5
5t4/7ZPngez6dpBxyMg2Igy7eV6VkB6vTNUBPXdWkja81iSFsC5O0F9NxMT0n2bn
gzQac8wLoboQlYbFEYVGqp0TUdzVMRVtvgMUPEhKcQDS+YjFh/wBg+wjW1yA/u3l
49m/WDLTj7Lx8VrxqUak35EhmnqiD6NcklRAoy63koPUP7uYhB3cOlohVfEEt0Ih
LQL185PwwP/0sz02hvH7RipgrR5ZoFR4UplCs1ctjBIHzjWSDMpUlZX/WyKQgSA5
3/CgESpp+aIiWoe19zYoilUVR+TnGCu8LHgudRlP2Gpbhx2SpO5wWqhoByHcO0+2
x/r1tBe5xte3nYsIIuA1XecrCXqF3rv0wBfmyua1jbKY3ddpv2dMbQMQUQI9ptBF
Bh19aZ7YX0r+hHngXAPEp8g3r2z9PIrHmpEjyyXJBoJ7Z7cOigX4vkv5ahtgqSts
CXlegVxkvT/5mlOK2H9ejYDrV/ZQi87mt/z7A0jX99rQDAlDz7C3A1N6Sm24OT+U
KnkC8kct+ZklodKiN4mAj/l9Lz06bGJZfXaXrbJhixtfthKUW0GenhwfXUAasyvx
A+z/jBG+tT87PDsTbx+g5CKAAZYDEU1HHqOjZj//ZT/HDUgz+RaGv/qjco5G8ios
z7MtsIlPv01M9NhawweUbbP+xta7xMMn7MG8Zbf+Y4xW1t1WLcgQXQOr+EFVhcR0
xkn6DMV7LW7fBD0ikh7gUHmSvTeG2TjLm5zX/L75MmPJVS3YD126yI4+gr28XFCp
uajF/HKu9TeupEbJpl7e1Lcaon8OAOqOpFs3JQ9xaL4gmQmJ6D3yx71KmaYoKPLp
duRqGvYShxi7BN9Ohzrse5DEaQe13FChFtJyMWNuxM0bVcAlU2DAZqVVGOIh6kxQ
MfyANhkl+cyx+mzCQeboNzIJ7bsX5bWn63YG1eqctqHwHx0rqw+uEavgb3ERob1U
DdCrjXZmCgUGqEEXzP4qsfiyqVGOhSY6GRlwawuOV4NXRh0TWwM9dTxshBSwgYMw
utpzxdmu1u3jcCmYUtkcWfnTeBOdmcJV8Xsjh3GqbX9bdd81YifhvEuhsOGZ1l3J
Aj/UZCEE8m7nxGoNnIVZFG+PhyvMBzeDdj301m99tlD5OFmIs2OnWYAeAFqwNdgL
G5YAqz1nfzERDiiGmpIJBkqnPBj7lROdsYSQicSWgPBVDi+43ghto5bqso8XMNHH
UDyZd5AlSUjTHscElPapvfrdHCp9UEXbz4U47IDMrvlXhnHsQC1RV3srGlQ5rA5l
W3Ml90uRNAxaz6ERJ/6ClIAKAM8AsgXNk2xcLz87NJ5204st32E2tPwg+bsbKiJY
9mWAtGH+7sTx6XBjgKif/l0EVs8kaXLKrZhvBPuvLJjpUOQDSXFWK/9C7JVSCRxY
6joudpcU+aktUV8PUkMSziSD5ErwvBButfoWi3w0r9woTpuHpF2Rxhub/if90Y5O
AP0e2NaJqhZQj+IMdZPJdlmWk33gwO2xY3sqEhIZlhXoHtjgaLXiLc5+DPdENHEp
EWSmnV4U859v1uLnwcU9HlsxYYMDTdnOUVAYhFKfP2XveVT6kSYjdibEJxnK75xr
IY7YEdUoM1VEaUQQQe+tr41jk82YFXZQACR4Dtjdz3qaGxs7GpPx4RiO8XI+hkEf
pB7/P3xQmGhkkr+8JF2W3VCQ+vMKkGiLR5BWchPQZ4LlKr4xEBhzRxMn0lG/U3kV
VDpPVXZ4l4elfknPek/WPrsdzIaqTuhlNOpPhtWZqTJovw2pq3zIyHLOatgPVWqC
w5qYy6cp37o+B4oK/PISbWxFZczCk/k7mdQKRlYqwV0XbjJvCxEwilUH2UnyiRH8
oO7ziMhhJ5rX8ewRPyMwibNrSlTZRrk5s2Zbbv25gFiDfhj0OlfoXzLXp5KWawLg
O5kA70mpayjYyvL8VWjFPpmx4k1ikeyIFTAwWzv6gb6vO/en8HtvFbCwP9t1zqYn
/KHoK0M5V5hX2eXf2YTG4hWGk8wmnaMv7t+IOUTlaAGAEfDPEBx/kIMvjLtVOBec
cw25CuwXuMnuOO6gA4KkGShH4A2+dTDwV0rXyPfANUerKYKhfPpv5vub/Sr6Vrb4
9BfJAtsHi1rpkTZSdkcai6+xQTlxqjVU8YtDoLnrj1qBrZ4B0MUiHVir+e/AZvwz
IqITxeWfCyozH6NYLmODYMaABwjRE1NcuXbjKq1o53w3PxNPg6YKKIOECfhM1Nxc
3SNEbz9r24j1hHW+fN2IOQ7JPSBtCodqqWRGi8oi5m6fVHcwQ/vH8GY/PvDIWw0N
jjoJ7AB0ATl3pjaTZc/7z3Au6ey0zlb9GZGih4KYx4hr5i8pXwY+nJQNmtyV5nXI
Xg7ugcDLKoIRlyboBbKsQKUSEuAf4eGIYYTs+cPIh3SWGTxXLwHQT1bYtQXWKWoE
mlwDscQY1cHLw37VcdOT6DXUwE/px/JdpAJX2Eos2CDwklmH+5byY7fdQIYaa6c8
bxpAy8QtcLX89fFgaQUzlaGiAzGuLj9YayUdVCcjzzKthvG+8gqEEo7gSe5EYWVd
APsCZV4jC4hgkroo6oiX4/VMTc0NUy0fE5QLUfcYO3xrlKmkP0dM8o1hgf7rC0tl
/QqFCkyh3KXHZ53qrbzumqmZyZLCyB4RSSu7CmU8dDgH1Uk9UoXFHoxZlAG4rgfG
cHmWKh/cCWt9ywYvIc0b3Lk7jLZ+CC/GjOsPFAgev1zpbPx6DybQWA6EP/HOZkGk
92YgYpLN6RJELw36l3TZryY+qLbvClf//f+pOTSE6F0Y3XQsPGWF2HHimmnMR4Ox
3zZJ/88V/gzro5LuLD/iOB84hb+YaQmkfU6T9xFDtn0fV5pXqkqDvgFY75EJ1Pg6
sSSag0BHFCVYAyBpMiy2CKAof/WzNJhs7V2XvB/LcHql8C0AGms1A5D98jwP0lIa
R88nNLReQEsB1uGfKfk5WnQ79mU0y0xeHiHU1hSuW3lz5XY6Ggv4YV3ghvadgJ9M
7NtVpXYBGUatakg4oY+eWmQJHjGMujlY0FYfAiyJXNPfjr9VaxLtrsgmYvgcoOck
UoreYVsXmsMWA/VdgPxeLiogimfrioLUK5xW6MsK/nS+abBoDcE9a4r8Cs7ZYMcq
dvbepY4Pzj1a9ywCPvN6x1ATbghHW8V7TY+eCsHKAPF+xyqhN/q7FNaONPPtFzmn
dQqxyr7bz6H1qqYZ4iX1IwzJ5P9X+7n9uDbZcwGeQFHFoMuZ1Zkzob3N4NXvUaaK
XmgHYLjHV110KB1o/Ir40WOjZF/ZSGYdJR8wVoa227JFbkaWOQ+1ITBhCthbeBWi
Vqf6Uygq6yXYZPrf/lDATSIWylgxJ2WxyiZ5DF3Nlf2lq+f0a7EQ126RFKZW4NPu
HkXLmB4IGGhn12nd0GT5dT9wErFuzxSESHNQJnOVqxUAUCjatBk+TFknaEFN5ufp
V9uGToUu4EOKZ0NVLJ2i39QxECctby/wL2Z97/vaXo/GwtCwrSt0cxxjA+KR4qmU
xF/JRw7AUT11YboBm9t2DZUW4bQvM/vyKICpPI369h34lVqNYMe9C61DtFicUnMV
kSbAeG4FsI96BRZR6gTm2N6PVLW55CToLWFQ+roggxRrk0ObDXCLk0lB/fQ2nCsq
qVu2gdRI4I5EYkbQebP4PM7Aw63pe4vlqqdjsHF7pve6Z9HNtroDvx+zYynNaM0x
cgjBAgaeLbPW9NJiSQm7bpxT6/fyCFMiGNp09dlKt9VrR1KXLVKARCYvfNuj4Jic
00EFX8h9Tnzl2JWBZIwwH4c/umhmZ1CejYCL+AdP7L0N1W0hNNytUX/G555m2hX2
lRsPocf1nZz9pyf8LR/kFWGkk885fGpxvBW6T2h/gATkdLrhCcajwSVRc0VztUrw
+seCPVgSB8SPf7TJA5YtzI5F4FvlzKdeda/2yeeftSf8s/eatjvaPQIQs+mG+G0/
DAXkYx27jQkGleZABKxeyg==
`protect END_PROTECTED
