`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sIe3umJNzMQclHTTuojbj50DXSXlgEEn8nB+yIrmwiUwzYVobYW+//TK1X2Num0a
u2yuUykz6XUUHQh2c2FUTY72RIwH+OmrnBSmkX+l7EViaSXjWJ/oAALSNMoglfu8
4gNoFp/m51sdT68WYMp+Vx4hflrGZD1b1PQASNIqyjmeDpPSlOhM3K0WX1dp6Joy
Jk618KBR25ccrrgkkcRDlrhKOerIFIfg+ovNw6b4/SNG7w+3cnUz43mgYrjrYDOo
bUICxSOLtlC12LsoqGcmghTzy91CZpLnBUcjlMdYb2Y=
`protect END_PROTECTED
