`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JgnxDLzLg+hnqyEdnt13kq3culwZ4jVPuit8bn00ss68adxrDXJpgtmOE+OIfpl8
E15041yjCERAJ9Z02MuAng+CCRlDR7O/ajawdhkzzwoNzTZEYhbj3S6DP8k2nEmX
uCttfeDK4w4eZtl19sDR0HAzQeNOtnA5g+iqyZ9SPQe2GfvX7mOAarxD2r25n7QE
PagK/h/QJG9gV2mthxgj3mwQPGavIzABIYpgCRE8UXHNYAHHbtBPGvQXx30x7Xwj
rHkzokUpwKNUX70Etas3Lc/jPriQ709GeSQxgGdiikZz5XjzwwmWWcaVcLNAAKe7
q+LBL88nQHNHlgU14cvTVphaqPbi7PU15BUFyv7HRvp7iPcJ5OqYr1EwtKoMa4lV
j+NTd6+v5gHYDtC6qwXyZN/8LQTkZgNzJQf40DhW3AnPknhLHtcbK+l+eLpja/wu
RJZVM2rh353usmbEnz2+NGi7eJcpMv4KVX0whPWT3Wq6I/c8ilFYc9SMYTpg7rmB
C6x2KQza7oukLWhWkV/YLeoUr0WoGCRV6fD7Rthd22FNdB8qd84x4dDluartz+NC
yB9z7BaUbPjKIPJPna24Fwzp6GJ3CmgO+byj7cnq/34/D4VpjIHNw2SoJjekXxHk
uOpUUb1hy7Sfy7xK3R+kJfZ8zTbhPMb77S+9mhoLJFcoK9qsYvj5ZNG8wZI+7UXP
ebPXmyb3fJBC41BUt1Kkk04xJaLNgKiGHmj+mcRgbCZR68o7My3WtXTeOB1o6Fzx
WsXK4AxhR+rYpz7o6Vds3kZmLNpApD4HqZzTr43Sl0UPh+RgqEJIsYYCl7i1s4Br
hTv4px04UwpwCWYAJjCCuUpIWIT5psVxdu9rRVXTPVIyHSjnCNwyRG5zqzzf3rkr
tF7sZrkjWa9ee11WEvKIdSbiOeI6Cs/eq1KZ/8npBTbvyFyq0+VzZM1C+EqVhTFs
1f/8BBwnoWWUJE01Rrkrg3cLLu5IHUMMk5gRCldv266N+XjTjOyw+lqiJpnE525f
`protect END_PROTECTED
