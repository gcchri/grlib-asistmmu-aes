`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wsnp7Kfk9elHTrZuPT6gI3SH2F073Pf2Z/7gUtADMgrzjJme51FR4E6qYBDhFwDe
nyQydYfDnvlRf1+dDjjobPrbzWG3Yi/6v45HLVpfB3I6gdzp12CXUg+Wj524wlg/
JFFJugOB9tZgeZheH2Y/I7FHhJbbTKzjACukY8le0YITSGHtMgVYTYg3C7UlBTkT
DKrJdGvvZUErTeCJ0h3pE8l5eSpmWv3qhY+LmmUe40AZmR/snPWrsDrjMlqVIqfY
Vu8DbLgkrVv4k4KO38wqcmqhVRRChffFLAKwxel9W+G27SU6hPQAGOFkkow3F/2p
JcL2h3niTM6LWijA1qqc1sHYokd6C+oWp0kaypARHhnpetlyeThI3l0bJLY3H2Tb
o1yvHWcXpEpH+icDV4X8+ajTC2TS0/yK+Zw4qNYFptRQPZ0rZLZeHoej0pbntRsc
`protect END_PROTECTED
