`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vBDWjg/OF23372NIMC4RIdyzfkiTTRuvhEgtiJlBhG2ht6IQATfONeOe9X9jowWF
vuggiBAcNDlwsgCw2q/G7E216G5uGuboQs/PW1fh9X5OnYCH0sGW2RFybj+XaVOv
nTXkGu7Bzur3stesFITIDSbG8vmLkVB6Vm0TiH7Xe3jbKCVF0O0tA4LoATZYQeEX
btugQd0CEXJSJiVg6clA5juQmfJowvh/ohCcXEYBBVT2NmZCHxvEwhHi0AAopjHe
2EdsikuvXAdMt9aJId5e0vzf6EI/6MlUxaxySYkg/xe5k2hkmcim/5ah8i3rvjG2
MQ0j/vD9tTh61p2uu1Her+zlcd+cEvDFaFi1tefvVKGuV4z/As0K00V/rRD9gWVC
af+tmoO4fvvoWVZ27JiaabsbiUZRAFns4B6hRwLEER0Ku0VhfIgOhSi3bETfk5qe
HQMlxeyolFhc3FaJ5wcEWFnew9nnrKA7z2pcRdsk3WS9eHBikOlsqhZfJ+E4GiW+
jw/QFYwVo1hR03+vRreUOkEKwRJLkZH+pfeLmCaX719P+1vVlfcypR9aiQkurLba
QdZE5RTYq3j2OKAgvNmhz//ja/bHltMxlnE2D0wbMOo=
`protect END_PROTECTED
