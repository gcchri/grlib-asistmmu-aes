`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hKYIIl9fg95i7Coaz7TqyaXox61AR0UYsXyzFEplqbPRk3wpY955Ehdk68DaHWb9
Yp6vAxEPEEsOVtofguZyG0jgFQtYdyYhkSOwjQ6y0uKbrcyHlsgZe5DNEasEOyno
PMjkqAc+CeMRAQuT1woOk8mwOmf4HmZ/mMVpLG4MILpg+bPjsGiIVj7Q1xT3KLEd
4dra3zDuzz5pCkkgTYjKOq+qeN3h8fiWaKnp97JmEBrJGJk4hSsNHjvfIyL2XmfQ
O/UbejEc5HvlqrFH2tnjoCLCsdU9zCJMhgqBW/oh3NnJwIRrfphcY78SJNn9TPah
M5ABZNIgvbzmyNIS8MAh1rKVZHamKfaSMpr7JLclm1NNPWgYT4K8kgE3PtIwljdd
MvW0AFQ0wdtLBBDMgUf/vOjuZES36pK3RqqmquvZJcwduEbGnxeAubN2sjLkMyPJ
vA+4IVcaoSgjL9zTr4wsOqLQWYbsu7Yam5XL1ADmWch7gd49OcsUfT66ed0NG+kl
rek7nDCRIcc0kQtBrG6fiQeUPQjGLjqvJDmJD16OWHlsZdsH45McWkJ/YaI1U2IO
0dpp1WxVTidoPLxQsSPSKJVkhMRNZC5sOGL0x7nwYHe7Jm8syMguF7Y4tPDK9AUJ
FgPxA4Y9Hl6iDL574vke81/1Ke6kkmCrhGeQM0BSDqhDEqsQyr0hXdaP26Btqjn1
4t/5p9HnnmY2dJaNyMUIf6wQMcb+Ct4iOxsnUVLo7b4W7pdkzNpwqSyTlCq0lbQ0
tEEpAzZQqSRnrrP2lG9d+NLOVg2TZrKzhsleps8TTZWHwhQNrdWlgd0XjUfGnPYe
SIfmSmsVkcSbj78bE/EjGAcnuoOrmPSLoe9TxFGQNqmbDnNfC42BwiJpc83NWYzt
NERyqKZpJTkrzXS8ldZybcQL1dSR35HKYkztWCzdRmkE5rZj5OG3CuqrmLHKguUu
kbzHISeVCTwevKmGxxzigpkVkpoKMnB062bHAIFPsoLAWAcRJmQCocGVx/ykSKvV
lgFxR1YIu74KiIIVh8GivCu3O8xY5Djh6UAX6qdbkC3cqfNU7on7QOYmZvvJyuXU
7QmNjGOQKFxKrJkastNwsjfT3RbWEAOIzUd607zauPFLl08b+27R6/fJJSWf4tU3
X8iYkvPr2ZlmLJzohikTxGdND501NHWt9cO4b1t/MMXSjsvNxkhJPOzOLqFaTvSV
AkkZevSrHd7XfHicVsrOTQTyL+eLgt6lmYWKppyEX+2IrNbHh8GMqI6qnIR+3/Zm
wxgZhKUcYOEwFbM4XwhyBRLhXviV/ZYJ4OyvdR7GrYtDKs0Pr1szEDjE2uproW7d
K+DLqGL2PifsWBX2M2GDv9HrRpP7g+8TjNuqH75zx7XFn35VRgxGIld3ekZTBpjS
IzLrW/lKOywF4XmdEp3pMK3F/RY+GT9iiSHT5ceV8htV5sGjAykf6w0FgHaaqFYF
AvwmKz+OrRMuPx6BQLADstC9LjD6rUFrS4A31ERLvfRcqoS8CyVEGS0Ic8KJpor4
PV5LAJw8ArSoNMbxHbKpM5qt0q3lHRUDzSPcF8KNn1XDUGDb6jf6h5XGgqH/I97s
Tfdv7MDM05P84ZbgKH2JJEiaA7a02/GFPIcpvYaCH2A2epVHU7tGSTiyW+g9MyjC
L6VL33fKHPDGF9iLx1iyK83rf65/7Ndb4/aOjVlTw7JQEXmK/BsldVIocvVgPITR
uf187nYttBGcC0Wwz49Q5PDVWR3A1TTkbVW5jE42ZlsFsOKAx5OD6JK3a0X5JMUV
hiL0LqHRNOm2WqAAZwYOUqvBZHxxy2VCPDmIAbxbxZAT1t/KLFL1Gs5c/fNCt+tE
Z43hhP3UeVVfy4naSRYAnxRnwhESO/SYZ+fjnVa9FbTFpU7g7QMz/xS7gMzIpUk0
1kxzzddP2hzEbOan3IY7q6dIOCKYJe2HnKxacsipLu8uAGOfvZWl7kFMX5DUE6FV
zBc7on3vK3d6cljqg64zQOIJwJII3NPRyTsAQuW26pNoV5ooF5pBrBZ9qKjzBM2A
WRN//9rpKLf3GTIN8JvndvRwEFh2imKUUDbam4KlMMeJXVzFgNtucpPx9HFIDCXk
csGCwd3su+Jm533696EFTDqfqBrU1qb0gr8cised3bWLSjo16BZbYNtCDJ39TVoY
8IzydW3dGYdOf4WC8NKq1TTWni0npqFLzH/41kocCOMqErcBjl9tFlFiMLSw+Xc5
/G+n1VUmdKSw9z47XzM5boBHATexKab9AOdpZaYQu7E+wFWRlGOomv1SLjLSzaeG
q9e7IgZWIK/fX8bhb3ycq8Z5wqXNTgFc965C/iMp92jj+oS3wsgvahsyNbRAEjvi
BX/P1vZGTCdK420CU6jlyCywyhM4tGv6KbfQvBdgHhBYQaXU2/eUwnDF+lWTLq2I
KFUiSwmXWDd3JS5Xp8J9IzRVvlAUG7+BVrr4CwYChpo24jK0tmg2UO6F2aREEL6m
dlUUxbfPRDz+KawSbI5Ic5kQ4XFrWcLNupsTRt51Fb2x//VEuhk44cFnPl0+J8zy
/tQVQ5k1Mktf75LSC4x82UQUvW4xO/m/nVmq5XEfQ2E/L0yTBFAK9+hzAHcja1DR
K11a94iE3vSIcJgONpS+/9sVPfz2nhn8ab9Ac0Q+uHxDD6Jg1yS6nzH2bOaWOO2u
k0YIZEvf84kivKi6NABVB1U6GQE8uqMZ5BxrVo67ybQUidAfuOgeTxYOQ91WTykc
VQSsuW/YdVqWmC79yvdMJ7FNfF9vhDCKaxQe9m39eNWfrwbUVuZ4KZOJA8B7ZcjE
LodNNA07At3jI4iddQCKivthPAarJGnlb64EwYntftqa9LHzkpxFFBGcW5q8beRW
C/gvj/B0XwefEwoV7f1d2RSptyAdrsl15DKIfoZV4yIocUooPGfu/VIGQipWlHkx
9CPhxT088aqYu6QRbk9yg3+meqEnMLrtTWU4FVzFdgzwW9xVUKFb7jL+jEjLd2id
EZWihMWmonKlaF+KmGs7736HbkU3wkCaSusWpzQuqoss4E/nY2dLI2pzGBnWofwo
84Lde7kMi/8LhUUOw8gVh+t5jDs/WklS0AtC/jNrMh3VVLkXITFm1KFUd9RfPVzq
omQe7uE0MsQlyaMNFkK143gxGNS+fNUiipqUd9GXN5pyRk71OqNH/x7cMlyVEdqE
0yWuDdGI3CUkh62PO8u77fPKRI9JdJHenHCzrEI0738lpcG0Alt/fBV0vAyKV4l8
e8OpBqr4a+gstJT9lV+5xrQscT42WgvcB2KqmnLKh/08JVApm7MHqu72tSlTjVdr
ttQbqTAoA/dmUwzPSj2aAu0uGfZSnMSNnqtEgYm8knX02i8ggTVvy8VeDNny8s/B
6NMFj495LGXKgjbieneQ94pTm4YtoGKKSSJZKz/xGp2sW66elIL1iOamhNwnykLi
29K5GjQcLhWc6M8V182k9VklNyrt9258hN1Ol8iUu2eQGsLlG0JrjfSHFoUQkMgX
PeBEG2fH+upEicWHcmOba7+N0Q8Lt+Bts/JNqsAZuHqCbEYwjydAqtFBV6fMHpEw
s51fGZVK3vIBPhCY23nRa0GJKrIDkB0TQ7xUVmytm/cZzwM3/frQExM7BUc0rzy2
DKAjANU43kYpfHR3wWWWLQ==
`protect END_PROTECTED
