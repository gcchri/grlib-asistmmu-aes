`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bwAqNZAHiRJYQ7tpZbZ7VRPPc5OrYo2Yto+UbJtkNKqUpakHmuBU7g6IoV+8WN2M
vre0R9s9/W4RkDpS01o+a8aYogmFwsWHErjeF+8c3VEsxpVRVr2DzcC9UIjgqMW7
IpRZOr0eMmhJh8/NhI3m++INQqfts5UjkBOybksdwGY7gLaqFg17niWGdIJU/aFo
axxMWW/hqh59pt0HrQOh6BtfKGNp7CwXWalEOtD8+tCJ/nbTKWWMty1L4NHWGB0+
51EZkaP+3exEMmhTvkM41TBp/8a64Jg1kzCjTU+VdD5jxAEXfd1lTvfbtJAGfS9E
dCQeavAeTqzQxzzC8TzK2WmJlJe72ZG1P+I62s7pYuaPqQBGspj9FVqqjyrkryVM
Tm2JjIUe7tJ2eLeNkGW9ztEbl9wmHb/Wj93M0RgG20kvpFrCtZX+2v04tq1wjmRf
NQBfjtf7I6bckKSEGzLMkQ==
`protect END_PROTECTED
