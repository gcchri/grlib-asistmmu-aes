`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dUrV5UKwUBOxNq2rsxarinfRmrWP0rACy2bKr8Y7TEDooY/vm+DpG9EBaEw+lE3f
lEo1qsup2HMfyX6UHhDuwiiYhKvCLloIy5jvIPO8Hp+QcmDlIOoTl9mns5aHt1gp
Ll116Pa36osRg91CuDgo4mmx//ETIO255DW5fmXNSvH/7rDcRCSFmuys0rIvuDP8
K1oT0Rok/TFENHejUu8AKUgu9wEoT0YFpEgQ4VukZiMFtiWJQ3l0a/HPCbb5n5N1
CNtcWL5oe6cM9w9DMrEswkRhMbKw46LntMCTYkZqIG4N7/2NeqceLvlvetYU5PFO
Z9VMLBxpkjb9a1agX8BFsSxkcoXCHlNq6HdTm0QjlR52YoOHOI4CyFus3+8xCTda
DaGXY0oporkSamtXESNjIe32cAtYwaid4170PhUqFFc=
`protect END_PROTECTED
