`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tSa2qu/lpwGG4FS+0YjUWGaKF3DxxIPFNdW7ID3SuFExrDNMR7n+wdorwU7eBZeW
nhmTY/1xJ9PqiJXXsTE7VxKzNMBdpaThJmHxqaCn6Yh5Arc1cSEZnJWrH1PQcmQu
NdewPTWFPlHxcXBKpQSpU3YpVDXp+l10tY3FfrcyEWoI9BNBgZBth5hAUxadzbM7
tYIXQyYoxuBgKc51YZFSXo6seapFsgN9jtMW12W4dgCIg32dqLbE1njt92I+o417
HOD9ZAIqth6m4Yv5eMajB6xBmNImmKeqT21FANKY6t4b/7sZYfLZltNFiV4yU4di
yXIvlbjiLLbyC5kLlIEWxCzpHxiYGqFhHJfBg2CRPwCx9DUIW01RBo2sjYG2ckqd
BAIzj05hcDwU1tJouVAyoWbTQME6mrHiP7rb99AhLr6VuNG988S+lg4p2n8l2MJ7
`protect END_PROTECTED
