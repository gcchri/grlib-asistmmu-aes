`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5gpPgi4hFgsj9xr1kjYoJR3WNv8Yy9+lUE6pwsSsA0eP/kB6SafTfDmOGW4q8nV1
EkcAmpPX3/iSz502nFeLPw/YoVtrPL9FMfPF4uUkYn04mFkQ9D+yMbGl5Ip3Jgv7
HOBepHhVui7Kfn4dfY7bjVuK1VHbaq5uZYy6jFo5e1BFeNO2yiBMHN1V40HSeFjM
9Dv1yBoFCkaLKnfNItL/AmQqaIaSxyzHJ1wzAkkBdW7h1lQj0hzbjIgQmcvNfHvz
zOUuCPPBOrhnCXFz2QNhAoipOdF81RTKh1dPKyJJ+7KBA4jSySsw3Kzd5Ln5A4Lz
bZU8f0or4GzX0n41PiftXBcVoMHHxRYmjM/p/mFRSe/Or88ekWq41+FoZpZcVGeG
4AFnTd3Gu3TQoFbPQqzEv9n0qOd4JObcHTH+cCMKoBXTa7sKlqX9NajPmjnau24n
2agKDnVk8ZDkM+NbrHMguv8j4/akb4zfHdAgonP3jkvdK5LvZoPSGsrfHzpTyfFT
HsfGXkZpjB3/OHQKSAPMyfBzZZafI+uSpwNjWSOeLtzw+NFVPo8E3vOT1iKFz1WO
28tkZw1yQ2TiercY88+94x7aX8aOPpnPh9Rwe2+5Mb7be4fY6cB8irbNSq5UT9cq
Hap0YFXswyQkI15cB5xYoA==
`protect END_PROTECTED
