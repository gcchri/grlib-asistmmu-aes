`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dihGUbNMYpkm5X7CTgLTd5PprjHAnWeo6dYpCMMStAqFTEVm3bwAOuhPAqr2grKo
HmbJF5ga7Dx1YXd5OzteWTjr0AiIzqyBmwSNZGt0Xw5rS+u4hBplQI5nkqc6AUkf
a+x4FNxCsUYX9O0+ivpXDGP3vOkm2E95GJXHHlErtQlwH+Mwi7v7jPvl19uecAnj
/vUyt/RzitHQL8dgveMVU8lLXomC69HKYBhxBZsnBbTPMIXwqEHmKdZ4b/ax+pCi
m9k4TELMFW4P/ZkgIzKbGmWapRJ2pwIdzOREeVio6vM=
`protect END_PROTECTED
