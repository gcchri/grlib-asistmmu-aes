`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OcFronzo2VFLQU5YTzYIRfazdnJnLkM7oiM/q/q5NF9zdpwMS6lWgsi23MAgwAi1
vNe24FIkgLNhPIkE/s7uNasfiWrkbbgcWhWhptaq3z12dL1QqhgznuzZe/6Rs7mr
ELUib582XBx2Kk2H+YGF9VIkudzgAWWbPbvZRd9Hv/jKf51DtpZx/kRRw9Yqy2A+
cbWeL0Sy8zIJGvHgByoAocFLV1Zv+BNOudrcxgVM/9u8uYzhJqDa2mel/XH5j8c6
IuVmxGoZ93nafvh1KRmH5Dmi2LHXmzAGk7NumQaoL70MgDfEhMUa3QILlausasA/
PPFcrcQKI607HHm62xlZ+A==
`protect END_PROTECTED
