`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r2Z0aY2JZjtoGeM7RvfNVdQot7KvjxJ8TEYIEEkm8VCNw9qcy1zTtAtK5vAHj7+L
2nQCUTvdhp/T607/Rkivw9instY1tG3oXOCkHunywWZsTal8KVt5wIzJGkSrYUtS
SC8f/c6OppiM9d20lKVmr0K01j1pDlDVSELTVGUQBVEX1+/oCOtBvXz2/ZWpkAkM
89QwkugKzvGhKXvBK68ei8xSL+WmVKlVTG/Ofo99Y7CrKJibe0szQz/VEHDhXenf
qxJKXbNtue5LatIvA4Nu/WFeDFuOQavAY11XHwH94fwPsnHg18aadxyG38KPZums
akLqwgGg0YmoIOKPVJwn0+ZJuyHZbJJ0QSCnjy1LDml12Rv0NcH8fy+7fLeQuMD4
IzcjV8OmaEhYajDHOF8GFvO9rsL6mHCahvsuzUNnWYkQBu/cE+2Sj3MNIh310xVr
ioqsulpDeyFgGiTCopFTufVGzHdFpQE3dCXfXU/bJo8LBtj1I+hINYiFQsde9hf3
0QO81J4AObXa/00XMYeb0V7RWkPmnCcGRdRPgWF0mGQmjnb7XXNHIQo6EkHcQHZx
aw+Yku+YyJdDgBhnv1liQhCf+GcBz+PgIAZUFaVkiWY=
`protect END_PROTECTED
