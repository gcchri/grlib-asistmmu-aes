`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5aUqR8DKCPZlrpIT4GsTBPbBTxn9fn886n01AwsXFn2cYPJWNGkWbMQAIIpxjzVc
ayJOFLsDkSn5L9Gr3F9PBgd2/xkzZ+elhx4QyFpP2v5d7Vme8EkBrEvjs1Lru3vu
SmVXuwAZFYeeh1AvhJo+NSDJZAZWtlHYCEZIe1dOWJpAHmfxWjX8kKUaIiYItMyx
YiOI7kpZH25sq6SeKdWH2IkTGdfFwdEz5iMPKziygz8a73qdz8W1aio35+nvEwDf
tfxSkhCSyiuXWpwZVZj/M99UtAMoH2Vw3qFshmtU8+IDXwR/1x/7xsgZ0KZsN+Uy
HzEfMtvJJiYiIaWUyfvGZQJ4zpla54Wp4J4jWroXlKrOvBOqkSOXZV9ik7tgJA/x
NH0N4YyUPueyXcUQloBn9DiVq8zZOrjx26I+J1cVnbQd0EZ2MVOMHGyfdOfe9IsB
lwtm/7ihsGX8LdlNeRjJjLISZpezUADZvT8Hmj0D8cxVYRrzC5QEUZBXTgX+c+CN
PEfa5isiZ7MVYpRNtpMIvC14WEkgV1/jvjw/2i8rkzPOCcAs3qtsgoZBaM/b9LC+
muo1b+9o+PbZzal/h4zbu0qzR07i2Xg+qSn8GeSKyzP7StmHSYUB5CmHrADMPbqT
z4aYMwAtQGz1+8v8HIC6TMGXnykDnYIgRCrhYi9gLna1y1W9fC6dGC1FYHpHPBdZ
UWI9683nBaaOU94MaBurfxBHKlQ00u1bLa/MG+QtOEJkGBuBPqcrhN/arqItzM4k
pFzVjEIA8DHSsbPbIc5I+NREnoBAIs7YlhaUjWtmKN2xuxWJHSybw0bk1l+NDu2B
/MrnySdEoxNTPLUAh6t4QaisQIsl8V3/UwA9Kumj9BDNnoeghQk0BLXa7Ja5LSRj
3seNxdzX9XawHLigiCO5BebQwOyiOglPnCdZmp8WFPSHUYvp0ntqCcih4A7nNEdf
cl6qeM66vcSYMuZOjdjV5eHv8MCzKc4nid307WJ8/oCiQuCAbea2bk73rLp6kGID
qQEDUy+WLDeILToXb1EzjQya9EZoBf5EIujDYk7B0ULzw3/NRjIzrat0yORSIQUb
dweoQ/ZIPAIUciLLxw164ILEgJC0lJwosBk6TNoLGX+wVF+ULxZDQfEuHhoCz81w
BWEN80HmGVpT1RmqOwcQ6RQz6jXS46eVrEQZKwq4rwCkHmgU1advCgDH/WHGc9dA
JxKILVL1Ao0jTLmrpLeBG7qcLvEPZNUeQ8oiHB3UjPZEQ+M0nQbj1pInKha/7H9l
IWnoQm1IwAidtlonfJOwgjMvw9MK8iqdQ9Xkz+bfrzCb8mfkmILkl84GMhoLZHXO
QsE9reolQXXvcmCCdvryNXmLiP8fugAudUTFkKdzu0368Dnyu/eRQru9AM8bCwFZ
h9AtTmT1Ldqc5VfRgT1LKiLOjyFeHZWpNaxNz1ytCIW7ewx0xypfgqArU15mC1xa
uXx2lxs2K012UBcW2rehxyCqjK8Huht/ay7siqmOaUOqY6t3ZxjosTOnzECgSjQz
LYdRqI+rP03sptCCErY0qpeflfFkld6M6CIa3MtjdT7WUqHWA7FzGlQy78oLPNgq
k/Xzq5BuPG6JT/H3mBj6WFR8bNPE1QusTEDzD6iGLBKZtU0QaTYV2o/j1DOR3Qjx
dFDokQrTm9nqJu0iq6U6H+WbSrfgTAxuqqz93cPc5bzaELnpxPhQ8q+Hs61cdP0U
6S0oOZxtxl1qAQ5RIuqb7EysIsOid//Xsr8etBGnmTlPMjZe/n6ImBa4n9Ggkx5+
vdjNzu/hhu6v7wpWTfsj52xG9UK91u8ZuucdxHeBYvwzO1TtSoSp724q8oOZMA3P
ueXMwJdA4atzDkmmn4cRX2n2nR2UWQnXod8JyJiX4cuFVNKfic7cREwVnJuV1qkA
fOVm6UPdD7RbBX/YZudKoLh/JkQDhhJ5wkdn/qQjqKg/btVAEg5d+mnF4MJxXgDZ
/mGMWPHwch27KmQbiJbtZ0YJmHg9Fx/pM8YEytBH8ybMCUZWeuIDIWx12V+z9sCu
TWeHicuRwSQfA+ZRcCthl3rx5NRMZIiiyyjJ23nqod1xdqnEMokflxSJfMg0YGTI
inkaiwtynUkWjOuMLDpqv/4wleJu8xADRSmKPWjMYifNIlcfKfWfq1YhE5wVXlP7
WTAjxHZKnEiG6+up96Wb2PSC8rxHzDAHdJJ2Q6zReOFsX4lygauulEX+xOc1j6/5
5mT5Sc7XtReXca6rW1muhWhpJbh1lRx+aw6IJxcXn7T8G6DvqsozJ3VIghX8T/ET
PQHmpkaFJBVfjr1iQHhU79+dwYGJEFxFcvRkYBBDyv4K3HoXg5NcuzwuxzlInk8H
7VmCNZLpC0noNLFqynQ6ujxtoLwFeheomtThm9VqCJTNI++IxDw7O6zAiWTlUg8k
Lt34iGQ1Dam8sgKZza5uMp+gvT3y+szrMaWFJyqNSLvh7XnnHUxa07NGfVR/V3+u
34++cv7YYwGNhzOd6pq2vT/xDmxuJf0ip7cNblY6Ckn+SVqbJ3hSv9JJNWV5b16t
PKbB8qGCLb1K9scQHCYdNIifc2eXKcfKfQ8ShIi/34ZR2Ico5JrZmRIBvcDMYuJW
Qt+lq5CYlgm3K3stJAq+p8tr3Oe92vna5vc+q156jaOosqMjVsSr+b3S67ByVxA+
Q8uFLXbLA9yjetiMS3mWCNasKy/0LyLPGkh61Lr94OCdnh7IE4Z+myugAp00+li6
cEs6TclodaG2BDZndxHQf59qH/BTeZSbPvHSHsRMSpRIgaiEnblbKUl+QEl7wPUv
a1udbfieDXUGWyl4pChTtzPbbaIubRs15qt1Q4ZzUIKOrHbb4ek8K/Xjj2rB6w29
mqoRr/Aun8iBlMPZx+Qgq/yaoQ3P3NcOSTy68kEhXjTZsCb/qo3xMVcTEYnDaiLj
qgCQlA/50nbPkwKakHRjbWDRwX9PMsUXpXf2lF6Lz8BSxP+lsgi6b9S3UEW6aXwu
2Hc20LHMaWpsJG//FM1HZmMSWAAlgJUJllxe1AKKA08m9+shapkDy8l8p8sc7fL+
Tt+UxbwoxFRyMA8f1z9k5dH4jJad8kb0ZL005Z6Uc8Np8w/CYvdjz1xycrDefhjx
Fh7C3Pbvz/ci+LDvsqPRuiwYVgadFaLFjQAf7n2LJsoYnco+9soX22mbBtMjcHbA
PHq+qLk2Utp3B6omqs7ryW8Bdn3jmQNiPyWuhiG8kUmwrU2CxAKIB5NOTdfEf67N
rQsyRZlZM2sjXFIwXRJZpiHaaNzmPO96lnJ4NVEXwK7ubR0jqMzF6RzwJbOXaaFM
+YbvZy+rPUb9sDgiRNu/W7qSDD9tgAgN7NOaccBIBIKOV/hvYv9HfjD8Berqtw6t
IEtwOYH+EqbvdGLaIMBtITpmsdzWv6jJya7gCdro4419us+Ca5fgYiuhX5gfqM37
nknm38PT5PIia2sHvUWxiNrV2X+TXbTLp8Vmk+QYRlPzKvJYA09RCfo6zhRan8Zv
7rQVRNTFYnCWDGsldXkdhOpI6jaz7HeLSonhT7RR7femH5tJiiobroCOXeEk2SZs
pWfSfTUVVof83/5tp7NSEub5HkVVgVgDlbFMNr3PD4rv7JXSfMRLarm0yZ41vBqL
5JxD8EG6b6HpwFZHSZX7txl6/YA/VpeRrS4JmZ7TV/WzOenHhd25FUhtOynI6vFk
DWUKTXcFauU7/+w+8y1xKUo6Caf67nXcJfJOqdzCy0jM3U/8z8KsrYaGIRG5Q0Hv
IyR/CGGKitmGz6MBflNngFpne/A7vA5HeogA5YUuUnTygR1QSGAPScY41UR8o4gE
qo9cuHTRFeku/a+Q9AyQzRCTbpMCrvPSa3wTc040wlZLBW2wYFmzsc+MW30RQvzC
inPJis2WKubaBSlZNMYtTTbPGJv2g5sa0aT0s2zaYeOa3pmlpQtEc80/40tDIIK9
CO3GkLITRKLprP+Yfo0qw4OJsIKWTgdgS1KUuPFESB/Drv+afcZU+34MzqhHvUqU
tJGHhD9Y6dAgMmVemcaiBYgaSblvH0EKFCFVTlCI4x2akBYRHZf/nHh428Z4PLIW
jQg0lPcYhX5/aNAE5LdIGO/5pTxyngDGl66HJk2VTEp19BepCt6YYOi0jrogGjrW
9iloZYnLoi5wB9g4V9WrZ4v2etQCeZuiOcnwvFOq7u/fxy6IaZscwmctBX3xrLsb
Cozs7PKMu1/JG3AgVD+s+TJKkz248p2lSVn3GUVr/1Or4Q6UPgjjQsN62SMu7ZUJ
HKhhdeKl8QyqEBVVF3dTtsA9kDBxvHz4+IM5Xf7094M9Ke+fnadSy5pVlGUOCPMI
yKYdNDywrxJvAgGAaHNMkJLpOCd/7PhbfBOqDnJy3YsQ2gTsy/27GT0gbDHw0OYR
8oom2BmKAEeDpseTw6ZVCN0ndyD6HzmqcNe5sNN6E/2tqdnFZcV0HmGpDJ4VSYDZ
ZLc7qVlO7E4EnC3bPy+so7dYtOdsDleRD41BwN0te/QqcOsepAGLs1qwDC341pMZ
HwD/zGwegL4L+e9zSPlxTDyzwQv5hSsc//hvJnJk0EDURKmHhFwmprZff3+N8Kdm
gJMl940LOI0uMy1jtMYGvxM1PDQEoEfB98tKRupufaTAqkHJ1/GApC5zWPKsWvWf
yq1Sbec8h2g1Y3LcCQ/+TV2c0B+CH4/MlcOs/asmFgcg0/xM+O1mz4VyZjeIF1/B
hg76l8GMUuYNj9gl57aZ6Ulg2PbpiSXW8h4Ge9VLxfhShfQFjF2hnrRz2UquxqZQ
02N//8o6M7MGG9SrsTdgmIX96DjiO4Zf/2rCBk6lqgJTTiZLk2k4UuXyJ6ETh8zH
dLH5uzRPgCXGDhIb4GmkJWRHZ9NcNKCGLkl1ku8KbvHEqYn61IUvuxM10W00uy4E
c30laJAGNQ8o7e9O91F42QsZEEYxLBw8epzteleLDUSGTuYoE+WIjNbn7P9X0ysM
tjufyWeCtVHWuwtgacZtKwYwyrr97K5K5nxit6vfmXIVcw2wVoEEeldxzAkkLpjT
RL2DDyobWgsjzHRZUojlJZbmxCrcM2yp2wckpd0TNpTmWm3vfu0GH58CeEgjeFLe
UnEidJ6fEc50wBjDmRE2jWe0bC2uK46DgMLHgt0sCtU1jq8HYg3zjRrDiyb56+Uq
BqQOymDIx/x30bEppsUeiNE6upmwtPPrXZyKHDytgFlywMic6YUNqqd7FRUnCblg
XoBysR8RQUQZRa1nxr4nCOw4GORLlvqu4SC7y0HFGD2FMJygSumSzvqFnR+dbRtz
2zG0ogXaMNHLbXQ8klOWiFVs04NQ2DiOvXzWxlEHBGDlFiLHK7wooNQ5EGAjLcQO
A7iV9Uuh/CWeNJSNpBDuEWX5mPpmQ+pFMeCuhI8DRaJb5pd9rR9bWffIuwYCjz/G
dFedMOGtNCY1bYlfkNHDrrlT8klFkYkzOLiByqZqrAUBqsVQE6i+lrijWlh/XCtS
ymdeuzjC09+5ISOhHWHdLMDuJrxV4eqPjZlTFIJ0wWlb0kM7ESKiweSOeKPllBkG
1LwUur5YrY2+8Ccw41QC66wn4SPdKKcRi5zsJbBSK5K6E/2/zPchuHLvGsZY2EvJ
XIEXjG+IuDlZP4gWTGdMHPgTqhn4t7VElvZPanMQyjeru6FGXKBY1LYU3fQwoNHG
Mym+SbRZpAcTOvzRv38GZZbkekBSHv+kXlgLg+qS4nAaRO6+wsn5kVEKHNzr3nEP
rI1spYYn+g7MSwWX4QQlqHTa2DDdREyZ6a0mxdWP1K8NPSgYfx+WKWWovyzUTr13
ziNxzIVSSLQgaKaTvIpK9oJRIR5ENWNkKcrJU4UOR+bBuIj09DZauQByhiY1uj/H
PastrWOjs1UBz06ldXkzrNM4513tGSlJSD86sTV6eM1jN09MOIfPry3VsVE5w9gb
gWOq68HiQ5J/0x0zczvPBYkTl5dpg76iseCHQRNpIlwak3aqXu7K6IktP81VuJ8v
5TLN2AJihypR1QMffXslztQ9+u7NbBlvoejnEcQ4FjKH8VTkJm1oSg3nNVCXmhEW
5ZkfXnNjGPjQz1BxY7o2N7ykOt6Zms0mi5AVimnYzJYDjzTP/TQMZcNWXistD/uh
ldQ5Q4+nFu+mYitf3E2ZXSC64rE/vv9x6IoC2ZYaCrphMPXTTLoRVdwX/bZ+hPQr
U9RDNVB2sl9Y1tAknx2DA90P/U3BXkM3qQQb4OORrCKbIo3CrjgUZI0brTkEqK9C
5HqilAtoAJ9MN0MeY0xYHX3SMqhIv0TRz3J54gpUvzflLSD/9n7IkRDOOovfwlCY
8tqAeE9IiVAZDF5l+o6A4ZCSLPAeHsERx+76OmQmDqNd3W5akTxS/R27FOZWorFU
VuD9lvvL//3De1jyL4PL/1LhBU0aN6S3/V2xilD+T6ATQgH2qgHmmZukc5WxcXMA
PIPFMUIwSzJyQBSLIG85HipTh6+U+SR7JTRU4OaUduaTTXuNrXszzrlVuvS9y0OY
NEAhvCKlNWsO3gzHizN0aZN/xWMASNJRZ7F32+3BKq66UtjYNn9PA67tonpg7AaY
6A9YFThlQFT2gQxHPzec9hrf/lE71Mj0SOLhKU1OomHNjlrIUQq5GtRCxzYT6ovg
KAkEpZxYgPoS1yQRLDi5O3dI16c7AKbj1BHpHw3nhoQL9O9h5m0ijvr7vRb2ZvFn
rZzu0Yi7mF0u7x9917kkLqobBem+hht6SlQ4WQn3zQ8rJzssND3TeMfldzSN6WmP
Wds4D16VlUi/L4CnGSwlqb4Rwkc2MYMrDL3aABaVsiOCh0S6FR8PLFbroUs3TZiE
QrNb/DYWECOOVMQdak0QRAde2M+SRVncOqU6DaNvkuOH8n5C1gpEua3ZRP2jmjfT
r5RWJvU50fX+u2ZpnxyuywlMCrUma6BszjqwMGiYh+Jic3ee9IvGLWckuKndCk5f
9KIzLVmtaxqunX7TkvuK4FJ/9w+x9G0Wj56ckJNCoIyF1sXlkJYmC1UgOo7sovQi
EGhshJKXrbJaz2Wo5NJkAWMlnAFGQH6XYS7jTiUFd61GH6EFSocG3DAL7m7m+mbg
byCwhT3DD1e7eTXLDavEfCyMGdFxk/y2VQJT61pdd/46HuOR1KfCM8tTwShwSyqv
XEv1r30b3Lr6TbgMi/yCr4ZNZ5+KtudpJ9d2qlvVia08NZqc3Y+LEolJSjipPZGk
sLcoNN1l5GA7QSK8UYNaGFVsZrK3opsJhHaOoG1Ypb8uhGn4Y+vdlBwKXtnSADWV
DvLOFIG4UprFwnxOgBMaiNfHolRL19SclvF8jIkw+Rxxy/ibYHtR0O2UF9NfVfqj
JU5pG1sPy8RSeTm7IeD8fRbtOapjr6AgOVplDAURtvSMfUNhi+WVawkQX5pr8fcQ
0TfnSLiwkYFbQqMuvH3/Hz69gc0TTgddeqxKPw/DW8U2pTfOT7oBHQw1m5pHAuOq
FJo67y4Rl7oDgo1K/G8C/R3ZN/Lo+eoEgaLhW4El3mhpF/Z1OGgojoairjMQOM62
MDViX6tpBmxQuyty5jTDuD/iLnE5kF4vVpSzRwCTClGPHrV9OqpQufPBnDEN/AFS
KFwPv0ArPqthkd1SZsRIbqqlhM5ryGNQ4120XOtmsV5Frz96gQXXQEmqiUrTK5Z7
6+MA6g8S1SSZs1kztJC296O2QdEhLZ1Nw8cptlE3L1BDTAIe5wjPtJQzxPQOA8Qa
XJ+cbr6FFwNTht21kAZv8cq4PDSjp2opfnh9++2m3a9K2SulzEF0xbbsJqzBzC31
1fRD7SWI8EuejIDmoNzBk8mqXgdrv8LEczvgHBksdJQiCxnwC2OJapnSjLZ4aDH5
96/1/C68y9OPJcgbXNxM9Sp66Z0GaZqyy2L4lEXJkaKHH+0nUxPqhW9s7WgbHvzc
/mXhehZqdeOMp17Skeu5YKGtCtM/iO3fCCDVh00accdbyFKLrGlKkSpGQObG83Xz
GtA8ybOqiCLDLvVE7Ao3mdGxmBbtHzLls9qRpq7y+l93joNtKhrDcGcDSnmP1lb6
P6WFCqYdLQs0sdgpGrC7dABz2HHaVx0EIEQkuCVP6GhIdpmDfFsiQKf05vL/xIej
lWdGkA35rZRV7f1WJ/UnRzTFPmmBbWsEjR9SpYNwi7gSD/pnlJ7NhMaKCk5Y4Gf3
+vCkx91xvFc4gYeeaSrgL9JUqekptiiOIYvlC9zxmkr5UljZ6r/EQ6grb/3+Kzqk
BrUSeQq7fJ+qLyDgGKP4QDJaxrvg2bJw8MRhm0q26aBh/V3m1M97D/RKosmDo468
umJVRyL7zmDkHggpnpCwrZEK9m1x1tJbdFfrduwQjq0rum88GfOIJkqSLhTkmvq2
hNj16euGFzxgc1f3S85+bIS3c6iJYplRXv1NBLQTV+rcqzwpUTB/On/gI4Iv4v2h
eLXUkYSLFjYS5pkmVCrsHHeuB2InvnsfPlubVb3a0rXKG03m7fqfjf+zbo/AMMI1
mJo89Zzwo6YUMUR7lJ+xGij2WU6DmHkATpEG+aThNODvgAilE8Bz8ZmOCxS4s+zd
vBYh0ksP125yF4dCRHyoOdPPxrOrJ/umUn+n3ldmxbghDmCPRJMP0k6gDBMmGEEp
oK48VeWvmAD8J+9Ao7Wy+aItL2dKusCo8DXsEO+3drdDkkRmKKpDkxqCEcyBBRqr
Uj+cRI9xQs0eNAZr0esRKG8ncBYED+fF0Tawyt7Rt3xJBBS0tsbMIW4W814jXqCR
omJefHm2UBTNbbbTxNd2fMXqfSEPH+o7I3ZR+QR+HzVteNf3alFtoDNLExmRCyZE
wb0NZwcp3T/8ZUon776y1TYXLRAeknmkrvXuzS32v5PFDgrCcqVmF/8EkQH8wDfO
HqLOSaoBYlQXbIFSP93fyc2JZVgOu5TUnOQ/5KVBm3wzWFtus5D1VaKXSW2hxo11
5N3PIJTq23STUSnfJL4G2gqPKuRe0GeSpfRELGMc7Ng1+von9MdNZvEYhqidgJL3
9mZM8ShOjyURUIfCwEl9CBUjIEMNrVzl+Wg2yPRL3LsgV5WDmorfnDopQXAAJoXl
ApiqI3HqLrBXpggbY909L1CdcbOOTE/FVf1hAvT7dGBOeL5TtvIytZisyQAOQSJx
aJdvGbA/RjZC7rVSRmHUaTiBQIfV1SZtlfNj3lFLLWlhYSwMaerB1E3Nz0xRPlcM
zkhwap2YKFFC8nQa8iBrAyJ1HpIA4mUY0t3EKZDzpwi5txJBgzgw/97GlvZIhEnF
ZBpkZ6Do3AoJjqYAseJycuYKTwnXFJlzaYpG880zc+jm4SqyHWZ+674483hEuIOU
4VuorKYqBgOHVznmijPgCX8ugnf/DI52ReV51qZZrQpq2aXFiTscx42+QuN6C7En
khJBMvUoy5IwK6GVrkgOvPG0/I3+CMghtM3ssxpKdZSM5bQr+nlAWh8s6fnUJTWc
30AF9sfGVgiCxXoUXjEWc6givkpWF3v3Kdng7eXMbK8TcapjKdb9B27QsSptMQPE
B7zjMAltjzVJoz+90x+hQwJHNTEnSSo6s84FtiGA5dXgeMBDgjhD7Du32jjqpj04
VdRz0WGwI5a9WarsXb7kbDajRFPwdzObyXiOopqReSd8b3ge/njxacKIOEkphgIB
SwD4jOWzRsBVkuHqk6HNfmjQq3JhRNHRg0gxD5/nnSl1SnMex9FPEmpcAzgJaws2
okRtJWWAaOUscvli1wo/xJESxEUwX52E5y+UbX7hLluahLLaBOyfxtBzLx+0v/Gs
uIwBGMW0uwn1E2XdcZbH0//hCMprG0FzHX76QSnoCqS6qN/C7X2YyTWtRhHqjLcK
LF/BUIcrmZRRixyg3v0TIP8R8dZqg9P8mq0i2muKCwn7dmHDp9OpLcNexAYqaRvn
YudooR0hcELE+8tykjmyhSKEXw/mPnZvA9MAgA8mF0nR0eyQyscDP+XBNfUBUEam
eCOUsmj622tlUprRQ4sLpsCNpHzi8OLX2oNNflvyBpSHhpEPdp244JWBC0NzE1ts
YJH/vY+uLRq6OnG+CiapsZdZyDDq3HnUGN4qH/cmvYYRVj9Z5rrHtmHsJAezlnfB
KCdXMyaJNx9TwuUMOD1M4oyWnB1j5HxJvLMuMJowv+8AOUYbQxUnKqaiU+lwJOwc
HeSkF9lSL5Cq23e9HIb9nTTvBbZb7KZY2SgjAzVZGYGYA+udw7SnokFk8fg01/5T
RGvmimlQbsLWSWRyYDgHmj8JFIHCE/uasY1V8Gi1wf8GqpRVlNl25TczyuFR+P3z
Ugx63Ieyhk9r1PQCW5Y824Py2jt563hAmzsbPg9F2LyhxJhudSJ6NYVqhbexITAw
JjfTay2PxNxHVOpSdjtaHo/o5ao7lDicgpy6mZrP2ywDO1qlqeHW5KeVeGNAGmu4
BuLwhGkiBwQmhLFLF1vTxNloyi25rRiN2KV3ypTZs4dvqlIQ2sOpwPRsgg+HCMWG
tnZIEkz67PLpbmc05rINOOZl11bw0H0d0BazqdfqAezPithNXWQyxRXtznkA2kIp
pfXM7ZKbFWQqiEaTHAVnL962bSiXPxUdCwdxAV65dauHG6j9a1J/g46FPAY9jrjX
UZwNfXREllVDpAIXKys//JRwQJ2KV4B/qwo8yf9ENzmoQU3BzVRkRmdte5aEeta1
LeTuoeTWeLb9kiQsr9wUhYSXe3lvpAlwJuPSzB+7VtYFmDKxfENfgVaNb54jKxs2
sjX7YHrBbEL2iWTB4vwcE4VN5eksldGpIACsqJSSfJ/S4USe7a5IF1IRpPpsrAhI
w7WyGQR3b1iG8z2eNrtS/Zi0JExncQgjfRME7ndTf+u0ctFnoWRmJ5zHzbdfKKjh
iv9szCMVXA4GN2klnOv3ocRvadLVh9kS8oHFws7FnofKWxw0eIqRzlCalmpYwJa2
3NqWBaIf/F5/f8AbVxIoWCqw0eC/RjoLiHLLe1U6ChVnPEGdqK+RUm2e7rbJKyXM
OpinqHJGGlOxXxocnsJzQiI/Vg3N9yh2tH3yJ5iiY1Szqgq26aglMCsvaNxE9enP
neRR/up9ds31bWHXanrsWrDEuaFhfJKpk8MlECs3pH+uBkLzWMO34uC3qyBrrE4u
BLp3dklZLK5a9eH+NbCiPi7ewVKtjOHn9RmvSzO3sNOWkoLuQEM+E/YDoUu6GRGs
BazvXZjXmNhQUM0U6Y47tg+HxyUcH4a8yrYH+yaT14vG4pjffDZanwoW26ryLjG9
txq3/DkkmA9KDNwoSFmPJzKV1JNFWHV/4p1mH8pbpW4rbDowEklWmxrukjvlImjY
GmQ/91y7k/Dmo+jyC2WFvbxft+n/lYLO515Izfov1ZYeN6OTskXdGApveBsmfH11
MmZMWy/ZsHx1+eSoHzX8F6fI5/K68HlTJ9i9uq7uPs/10HYhAXXF7bE+S2cpA4nJ
GAI8FcqDNHs9IkCR1cnLehxMM7oMC+TBI+1k+R8Fwd4UWPNtqznc/HtF+n5z949w
Ckn6ekxWTJD/CF+ffMOA+P/RjPHUXNNSFv888zgwO3KSdOGuU/lZVrnDhlMKaa3c
Rtw467+fxP0U0adw2igtugHABHHw1VHJD5nJJfzL5kRcnchPrKjiipsYKIQDyBig
hJOVh/RXG+pI9ZwDIy1TFAlyiPF+64fALdfcEDI2NYtSmoZD+BY9VDYewVrUZR3s
RDKj8Ubi7zHbiQhMuZTmPWfskr+mW7SKb+BpdbcBxGehI06DpRAYRAqHw695rZD3
TRq/D7COf0EnPJmbFpV2Z8DaUB82FGPA+njDIYcKVqzpK5+QqKn6bG3qwKv2RqPb
Da6UAPEUWKkmiTGEbaaSNK8FmX/OEGlrQZ0gmFkghyT/3TWRsk4KVWxqmghE0E+f
q/UyfMzUENQlAWWrouMDlrIyeG0OUYAl6y8e3PRflmyYqb0+Vaf/yg4AfNy1qNIB
ZLb2hT+C5nqfNpEq9/TYw0eiUdpsWZ/f8pTR67tu/bekYQtNFkT03uIpDKf+RjvD
U4wEZJKvFUNIKypZgTJER9bv9vhSmT+JrkzpQnL0Rf/paff3LUg0eOTjHqIfjp2w
g8JBkYl+jTnx9tHjfz25/lS09Lxy7oAsogxprrY+ddawu9riC3MQPZbiXrTgsgyk
PbVmIY93ofW6+bQAl9Tumw0LQ75V9bFn0aAVHeVBSDJWVSqBnb5ehIEIvGr61PbO
noDTn3hFOciyroy1aqXAG1ADodFQRv2oiqnoEsijNXTbtbKIosZcuWeM6hA9gtXK
89rQIEcVoP/zsChrC3y70wC7ebhM+hYC67X5LL2K1RXILF0VjEcKD4Jy+k4Bmupl
9kau/HNVh1ykFwxxG6x3kc3fBe+QM8JRg2U2yn7L9xtoL2l63Mf5kh7eIBlFRV+Z
VWh7MO7/tpGYgAOP6VjY1RUf1eSVTD8CMFdGwJ7IlWOqnyfLwsk0lLYapTqpXJiP
9b+yX7R1AfiA1dYFy1WTt1G8x84sdDvNXPcoXtWGW48au33TSWaQ2Dpz559Aj/rv
ZMTr7rS3bSMQtcrBF0UikYjRX6fwYCClWm3l6E8zfv6XCbxggIX4v5z6A/+bmfu1
HNCpW1sSUpzjfXi5LXCkhDKJF1Us+ETwpjdEIzqp0ua8kMH0GzEBjbrmTGW3Hp/v
lTpUHyj5KHkrg8fkzAbyXpS39Cy7zuCiAl6IoPwYfNlkc/oGQVJ3CXDhtGALSNDy
yH4SMrjuLLB5guKH1lF3r/5tuy1DMfAmXi3eM8/BPmuu52eYAUz2jTdI4KF94La0
WzynRaZux2/bgHmZyJijdzf/5Kau3iHRo6h+Zxy2j8xW/9JaxTbSmaDUPVazDpRb
3+rmktaKhvgnfokbgaJQjh5MgsgsuhDrM/IbhlzCfVIT4QvfGYZdCd1RwnwWwkyq
AAi/Doy+Acjq7Wf+NgjOW3yvoXbG1FdrDVjiAEtEmNO84Ey7yZ838cAoZwYRou+S
KAPZWKA70epAdB9akGEJhAnWF7R98+/tr4Ojo9N1U1BLvR6UpXpk2pu7CUbl2PUK
veIQl7LkKL6HJIPUDyMlxu9KvEryPReF47owx+s0Bjra1j/OJLap8JC6TgVLX5Lw
qdGKaN+ZOCWRA03v5piZ73nhuroCK0rzIpq08dlmU0mXxebQ8cjIGm/q7ft05Bum
/N90L2g1PVBw4XoZH0GVN9PzBoSdG4e8lhoUCLa3pukVHBasxSd2LGKHHkeIpzJj
SY14jGJEYtRFc5foOPFs2IprqvMc/0xSPGPNMKpv+zxDJqB6Clj5DDL+pIKCiLQu
M4lAqPZaaa/4ClOrzH1ef7uICs3h3ozhNmnf+R9lYonBWJghQ4JZxmejSapBmUAb
OSV4847Frw+wpVS2PEE0BQVOqh9V5Flywi1MIFH8Smmmeq2BKZzfwnQ7Ho5+VNXv
r1k7yUY9I83FOJYNq9RbmISSTv5VngAM5mJaZOUXU/jRfVHfxujBrV9/UNNTfiVQ
0KeD0UTvK5UjXSBn966wVUPoNACa0hyg37pHPbkpn5W22RP1jdR38t2zmTU0E1vK
0lJ1np1r2US9/0S9duAXoeezYBARVyiuMj49SAr7dy0TNU2375Ifa7ZiU1tJ5Zyy
jVy1Lhk8bijJyGUBUXVbRKObbGR4uYVH8nHSFP0Zl+ivlCKlbkhXcA9ztPXVccVi
LQ+YAKFlzXiJbhMmAhoDB1ASv63i9LmRevjJARgE5kFfaKpFsgLceu1zJv6wQuq4
bhc7aZ3H93CGdHSC1tYmd1qtyYbK13KmxpPjr+Z3nwJUKc5fNhUpV03nhE+R9kNn
+RTuQ/47rRzQVY0p4Bkpq+2JvlufNJKz6IMLtq4ub9cOEe3mTPoKRbTklKKAU+lp
+mCbRXqhd8XlMnLIKxM9HXxHLY4jEtgIJJKvjSMYcxqj3coUzybK2Ktb+a7MfdeS
3kYREZhY6yF10Eocanx1L7+Gct/Fli2e7ac/ad+JqDaq3obN1K58jLG5pNSci1GX
NP5UBekhnJOH43bNbI7T4zpQ1rQYCf6gSj7sze/07LYPfVzFwU1azbjogtAOV+TO
K33upuCa3PKA+6mmtiYuQ/oCKbCFwg5H5K1ozgez2DNd+z67NqqRMAhLB4aa7GYA
fNMwkmg8TuYQs8fR5zINbVS5hN9c0BMN4OiWNq90soNTHnM2xvyy1IvmiauFELYf
mZpaId7ig8Geu5qjN5iX5P3WTovQ5+O/QsNsTnR3E/NeAJCBIE7WrET0iSBdpE2g
ucGnAtmAE3RXNFVm1jBsumvRsLbDY1iX8zY9nfTMd7Q0EPu99l2AHcaIYaSN7AuX
fG2Brw+okzOxqswNckqPyxzYpIlnJzidn8lVcS+zzxP1c8w8QXhmS7aJHfVpQ8lV
sXZ47ZXN+MdTZMBapwtm+f5soyfOFW/i3lQfbCHVhgkisFdz3wdYrcRwhvBevEmx
b7ZRgDCaqP76sMuhr7saTtVvgg0IUQH+8Or7QyB8h7i1/4QdwGc34iWRMQ/kZQff
Q+bsK3gzfuzD15H9Pw7HvAf76Hxn3tnX1zAGeBvbkzygfBG3XAQkWFZpjXrNc/ZY
+HxNqt9hwnHnhGdg0r15aWf/Rc4+7TL7e6ztbGzmGUhMXUUeY5OEPTVL8OV/4gqh
HMwapGQ3ijgCWbCvIoBDW0Ju0SNeRKNYF3PYhBhUzcmsZPkMWVworocXtnJzI3fO
/AKWvEs0f67na5iMua9YvJM3gGad+VbCcWb148hNbhAGVgvMpdyVE8+Ur2jDKfqA
2+8gr7N0qLDj0CJcbGViP60+pBoPF/KccPvDtA4GVf3QRSAx8qYRr3Q/OnokUUew
diQxWwsK4h+etNkVxYxL7VJMK+7HEHtfa2z4hfZO52J3UPAQMvKZOsCAgDfZ7EVD
CuwPvOnFv6+kO5NmyOr2IaK7I8YxQxeSiVX34dKplZPlc2cqIrIIQe9CiHGaPpYa
GeWc5hjy7RpweZJ4VZ1J1vJzcX61EDphmjT5AieN6a+uZ0mjjtSD/yW+8k3MUtao
HjxJpgpLeYMe+d4Cfh1iUZelJ4DsvFkK6/Ai6yN7z0zlvJSOVvGWDCFbRUYx7fl7
mx9p8C1k4KonM8a1RVbCYW5VKq2JKciHSozt0qFO9P6Hvxqc6P/biFSrR0O+aau9
sikP0zhF2wIjcbSOGrlOHOvY3cwunRUHsINgyy6N+ja9TXsYJaZamCiXKzcvXY2x
sqDWVHhRu3YjRWdy7o2/ER/m7EYz9RLaxkAS9IhA+7aC8qetxv/SS34uyUyxRuPa
EprfluyGPiqSOslrTXvFo3cXBJ9Wy4HzFqWlv3Su/icEElu/9McaoEECHGehMuBw
SV4lKTDtjgfk3KSfXP9H6Eiw6u3AAzrP5fWJEHGAC3vSTK2r9cBLaHRrSHqTklx9
+34AQNqmSBkZ5alH1PdCIVIKiUKngHyYJC/IcCj9KGd67QVK7mD+OjtbXlXWycUz
LoCA9NuL0ZMBdSEp84gQS/joXRhzQ7gTmAIdKrI38dCIDYiXyeNUwJSR/U2+Ybvw
ter3v0wPjz1P+7E2Fd1/Jt/ZK4juGQhkcyFHReElZzP1Pk1DniDO6JOspoCv8MYo
2k5m0bHZBMvOH1t7tcMOguYy43QmF0/Qf3Y2hhraSd9xq10dJ2X3q0FLh0cKofH5
3VoWkirGEAFXdBRZn4bPODPDaBQSnq5g6qDdjaHXtPiClEWYRt4au2B8wSUMJC81
Nf4b8unA9NtWNsFIE89igNTOt5Yqil7vJTiosL/RwloD56ygsyWxBpkWyEAq5aPa
aFYgs6s5eWM8hIRjx+2ITFFvseu5nUv7xrb4R/rKnWrfEtFNNmXrpdR/nSsZfRQF
1DaA87Rjlz3mUAO98gqrbwK4LQve7bU5PTXP0pyYEg+5WgKF8LqPsP8EPhvOz8Rb
prnyaJoK+EN9BQqb+5OQ2o4YcR8fC5xcGFDZ4dOBU2wV19dx7WEaYeYetNvclKl/
OqBek3MQ+obPcgJzAAqmjS3FuxBuJPOMDdiqF1oOyLznM9bplvvPVpYLa5Uw+VOm
ELb6aoh6pTgXZPvCqf/DZeOQtDyPJFkgQiB5dPNdhKqZtndJuWA42NQ4Cz7D23W/
cC8XPtJ2KDbDvyi6SY8Ind4iQXoKdsdI+E5sP1DU5jmJKNmUfPQ88s3eAkSjFG97
Slj1JoQPfunG7fe5NVsmJ4pLvLyfWh5Pr/URAThxNeMOPU84pwkKsU+alIlQ4qgF
8HE5F/WZIMSvEQF65lMzJCJuvOvJd+D/K42gcFs0fRQNwfLazo+K03KjiCObuU2X
nJIwDd6sP8p5fRHMDhhxenqibZZTf3UZmH70fB48JNQDXAMTV64o/fGiFN0zq8tE
L02IsJkJFsAeovDoQELqH26bk2Q5Gqk8e9HM6/RlkwTnsd80d1Q9lLAlwakOQnv5
MsjO56ZiX2B5D7T0tzkQJkQr9kugiwCAeCDEsSkB2NkV32WlyWgN+yDax+oktDoa
ceOirStdOrK/LZ6PNwy9cputHM1JB095yo90EttGor9g26kgad913/ibrhCm16gZ
Cu1P0+79JAjQknSzZSUCWBJKva26pTQuPOSAY+gJeaFSrGvY3O6CtH9FEImagC0u
o4GiFAJ3NUkOmA6gU27+YQV2KjbcaCXzWE79uKLXXpS7JeMUpYy+tgjQbETpzfq0
tMsxJdcCAxNuDoYRwDiO69+s6oobDfQfEhkGIYqGwkNSS7IvUj2uPMMjMjvHGuJJ
ONn+pLzbwnHOitQkmK9ECzokLASKBwexwctxLi5MVOZP7+MTMatnhA0aS1h5lzQF
QbQUUweSnz3vuRmoI2vOesGQEEzss4RMYLZTrl7EASF7fhgtvtlhAMqaYCVvS2qK
p3T9XwGrr0dMbJtROfsG4cwSsStLtw5P9sVs1DJzWJG0AyitC31iLCd8dPkOOUPs
c4w4WQcZz4/HW7M4qo89RcRETcVZjFSAUQK3MK4ezs4tM3wIUivXeAqgJLVxfMxE
nUWamTWD+1R+IIYcsICZzyzh3BSMp7oxRndqglDxv/i3ESL1GJPgf/q45scJgJ3v
CU/GqtfptWvdoAINvZ/1wAvo3VSUrshV+7fPuGjAVAAI8wvKRO2rrB/hbCl67BA8
gV7LK/ePKHzUC53uxBr4WrggCRCIxmERVaFnYcpkoRKKcU0W9OdHgPcuPMgQMDZd
bHxQUZcbLnbeeRye+yxxNRrXqijthuNf5x5GgTFxwgMp8FCl2Yo19Kes1MKN/RZ+
TsD2KT6VLY5JGJ/A29y75zC9nyj3WpuqzDJNRu4GJVrnlBindjTeBAYgz3iWfsk1
Pbd0iDL6r91tbZ3k9rL7aM8l614QK/JPOzBOKDxMlNqhGgmvF0vVuMJkGyV+niqm
AZYYQqbeT6lsqGzngdDpqXt2ddgumKvpH94fT2Z4Lu0ibjguER7biizsBHxT9VfA
Nv4romSKRqhqxcYeCKr3KF/fjp9yCmzlurrYBGYUQjbPf6dM7qCFFUryJLZZF1Iz
kBgvQwcuAamiON0tfwbNsnFOaNt7zH4wrHSxxCdRBTrxYGTFJVZ24raSOYLlVKsS
cDR7343Bz8aCR0Do7gQxCY9ybvIxxvVENuJ9htmrIby6vHW4HWpV3gQEDgNChsy8
qs6/j9FxtbCQ1d3+Zg/Vw1ifcoR+gEbAf8C62C7iXiufjW/td04gO6T1xEaSNIv2
baba6wPBhtj4ydgczyj74346dc8womlK8ioZCVsgHWw7jhfccSaaGNPMJO5X9zTZ
JQBOWf8ReAgI5CMWhV9ZyWyokftauI5wu7VIUOvpqQTwKYTDuVkuAZ8gJruH6hNg
G8cEujO8n3BW1/n5tLY1vaqCFUshb45E8knhYibuPLplMsB4zxCVIjDmuLGLNEEK
goprt8gfvqdY9e3Hom0W1ysoBzZ8F5nuMKjOKkdQt3UH779h7ixYmxGIh2sY+/Rq
pldQaIsow36+kls1wH/XSlPLjY0iGHojTkwhB6ce8e44g+f5WAbJzZE6S4kPnm6f
TgqO+nX5n/YVmoJztv3ZaSDR50i18f2VnUcAIA3j0qyFaz8KwQiYRH0BXpfa1Hdm
ujQsoUsx6j1UqiAqGeeDVvEw4hROyzq9a2pTCI3Pzw9pgsMw7WAK/UfhGcjQmS3d
ctSs4Z2AfAO2kAQvzQD2uehHalqs5sssoPp8vnJFo5eo2/wanQS6fIRG+6STbxcG
5PD2pBqAKYnsMFymzjrtV55VkGc1BOCWr4iNjlzs6vghCo0ai25kJHcnQ2aqYApd
D0c7Omczjh2f6IW7TsMeAOmrcuta7WHxF2AOTCVtMBnA9CEfgkEjkoi9r45QbltV
7y8p/WFcBGeeXHO+MMAtUkEoexeRzDnBvxZ6pCMjww/BrzIIBxulxYZDwJ03Ivtf
GSvdmolnXPEI8S0R5CJsKKmmpxpk1YSsQWkFkz6FmIRDjqb3EKLG++DkeDz5cA2n
yorpCr76yVompRkKRhpJtsU43A04ySHEhYZMg9iPZ1aBv9Euw6lbPl3YBdd41qPx
Tfnjsx7cGOmWfqz42hi2yh35OEpP8zyne62jTNwKtpDkoL8zPDpce81uMyDKtvDP
KMBgX5iBlzcyreN3FWviW4srZqe31ljvYaXdHgkePdXgqx7z369aG/V5pVK2gODk
Yqo+FKoOI92mA/d98bfKuhfcPYXuD+Xv3jTPGOvtwJjjMCDR+pm1AxDxGRnr966B
jeHGih1lxcNz2os1l/9U1p8MW1SwzyA9y2jv6F4tOXnWn/l9SUTic/G7QhUTil7z
zVxZbWAl0/UHf671ZDtILFMzpovuujQTcQtAuxwGrX/IAKeiBnZXIxz1rTP2F7cT
+83x/JXFoZGavbqQql1rRc5ZeCJz0xzs8CTepxDaMgQW/hSYOm/VhP5IbelHOFks
hax9RDG4zUNu+5W/PS9ANz7O8g5b4/uKQyFO2ImuhnIXTO+KeQW5keVcaB68jLG2
N2cGdk1wEzSLjAhsus9zjXlup/w9i6jUHFfWRh6/Ko4ufBqxnJoAC9Jlhe7St1Sr
NqHZfMWiwpYpec64qN1Q/QtPTwo4zb10M9IlgCtIw8gbpt6ZiYzQoDD8YsIltHBw
Yh+zohkihLLfzumL9K3ycb9oSwNYZFX1QO2JrCp1qKVDtX/3LPEOL7Y8hFnt0/0m
bsNAgZADKc+baScJPzGt0Z63wbnrsDX1BzTn2Cm9W6q7vqe9R+iSet3tTkeht1OO
M6MMnTFfhHnNlLlkDN0FQspHCdlEnClueLCJfBiCHjL5Mtm/9YqqSrOSGrHJlp5f
LF5tH/NGHKBXdq1VNQhBIxwjx62QFcCIF+xxt9Zey2jvBJQfFlA0tF9BIHl7/7xt
l02h6mWeu/8gBXt03vLNvKnKZ07IuADBvOX+HELJK6wwcholrJ5lLWuHvgwAQpzO
BUVBWyAAfVm5/7ujUxHoCcmKJgcFFj0jhyJQ3/A8yEShj4gId7KYh1BLd0kwBW7H
tlEfsNo/WCh/MXHfA533FzEljRmSE6Uzg8EEmo+dRzydsMhKRxtSPUsR/jgq9ZCc
uAPFctOQJnbLyz7KjuwujDxFNFHpbiklLMmCXfu3Th+Fa28Hl6akOWOP/znFWp71
9wZx+XcD1KLw06G/DZfYKIMRvO7n28CXDxZ5oC+qBE+HwK5Tetl9beYHTrTMXRx3
BToKeO/BUbAlKEsbSR8W/gMtLJbgscV7lsJEMm9kr/VZiuDkt4gRitCc/+7Ue6TL
E45WRD98gp2I+4gbtascyqhjJQTE0Qp9FWj76ws0qNzJtcRFQBQZYUWrK3mgR7Kz
xptcx4cXW8dniOvFFXM4WBKMeHuQufxDGKZUN0f/5TQuSFTAxqyfnCHr33TMpuMR
yir3NiCRsqE+CQWTjM2iU4/2D5pSyFKvhCr49TPmHDt6rQve7JhUr2mVnsasZAjA
KDv3kRa7DKlyzSMADbWGU73A/HJmP2vsz3hXV2cIbWdovIR0dN6SdEAICpe8c/Ee
wKnCF3aP5hI85A7a/sNS4KXEdyjA3TGFYvqBuy4qNmzNXRJ/RaS/f2RDPMSdpKB4
s8BzSFfD8fEeZqY41ZE2J8LPelZlPzi8SJWT6saJ0+wwiiSnHVxtPDg3LdiBbhDI
7K2klnTBMbEpE/L+e6ly3tKEFwQJQVxpO4Rq6mZRj8zsWocPWLu1QRCGTs8wfiM7
oVjJmgZ+cjT7pSHagB6fvISEQoNft0rMnpWPvCUht0xw4eB77ZKktdW3QbVBy9/9
RoZ1hS+LNx0KgKFOENlrxerJLYy6U1EunX3BLuOWMeORxflgYCn3Q9ImldW+jmPf
tP85vT1kNrKe2YMNcwYYyoWyqyYDHYL9NCh8J8286pvKFPxKZF40FjbdsA1gdWXX
aWDSa3M2IJUYGUIi5jqEUp4O9GXPhK6++ZUCJpD7E2tTCnjmYSMNha6Nrc5yXswL
dbqRxliDhI2/0I/LzBLehxfUVvPQv6offXJpe5/8alt5P1NjuNI7teGeOh0CUFQE
nukLDkFqguKCfrqOAWP5ScCtDJCuXeoswl1Y/nNfskdJqpXa0hLZRIg9ogGMiPOm
hJw5phKnlUgfUSxIvbxIih/DOmhbiTQy6BMEZsSybSc/N6ck5bXpI+vnAMQe4pQG
uUXKwDvHj0h+6LOnvKpTbFPCIIrxs12bh3oebDy3+dU2W7kIuWsO/xgi//h3zVVA
OWCmb2csV4mScAmwHml78I41LGiWsCVnw9whEGHDEgIwh7m7s8E/sTLuXl/Quuuj
7vrpnS6FKsli9HJjSj+3UvNaSy2s/OGgRYUHpfr0QK4u7Ni4gPYY+rHZ/VeHxXjv
31BGp3LTKAN+ZimeLevDY3hoDVWz+lZ0CH8RL9mm9CbrkIB4oiSi3SCrqxjgw1fF
Fk+KE99Rp8tbW1kVP7vpiJtuOrWvKjzF/TDLKidwKXyDZmDzaD+MjaDl4/uysAEa
x4dgO1NnjdDpo/pOCgF1hhaWvmuUHOIOwJlmfSZLStBKqpyU3xrTZ/hGmPzO0/U1
+7zIYqvFMYmq7SEXJdUKgotpvlI5H7UGY1fPIJ2/2tv6nPCdRn2Jv7O2y9KUXzUl
Jb/HOyt8W+twjmC21TI5GRGUkdP1ibwtjN9ygUqcmc0FsrBE9chf86Jh6R8i6bhM
FyMpwNwAjnFaf42l4QAVoNh5QMFmqNaVQ4J93EgNmV3fcqYLJ9N9Jc0j/shlMeDe
qM11hutn41ZnDqmxdgHTCU2O3qPbMs3bEbtl4Y11LF01jvPR0k1lml9PUnjseYaO
HXsVpQqBdfeOgscFhNErg/1SX7doQ96RFo0lF1fn5iO4fYSq4fzUe3Vu4cVyI0HN
FF0Zqcjmq2Ppln7lYt2VKptom/btFNQZ4Mfn1hmFPzgJrbjpIPPu2Py343jiu6M8
4pirRbR8Kn/F2ta5gp/ewKmv678lT0Xjeh29+ypifmzXeXWMFAiHfLuSbdGdNigS
NaJAPEXrWafmUhRuaK1XM7gIUjwcXiwGm0QL9KzdkzA18Xo0Ro5zk4U3rLFF62WC
rY+EHu3LNndeQo12zpFZG2/+wt5ISEyPY2qFu385KOA8QRNLBWfLQJOejIEv2oQU
6c99aOhHxcwfSxymkIsRxv60AV6s7RiElDJN/bt+RIGyE0Cg07/zgjLNpkK4CBRU
VhuOFVA7qDCUtE2zjfDz4TJiKqHCG4Vd351OI4WJ046l8EkyNfqYB0UMNUNdiwM9
wdpzerNVF3QkaAqh4RqQ/tr3PVomG/33YlEvhE/pvalrHQ2oNS16y2tDAmiiXFpt
OPpDRkjj1rtN9jyq4jc0li0GonXhP/7C54IJZ9lI7MZZq6H1My3XrID8BCyLraXk
xMkMx2xQlqnnC9ZVIE6hv6ToDbhcqmfBZ645ALEMjX3OsJKECMQKcQu0e1zrs58a
KIXqZq9T7BBcni8cucfuUN2/Fn2YLO1xTuvSF/+aIVLQmMqQKdhK2cqYScU4wuw6
SEtZe8CNBM9uwYDIo5ognOhBUNu8vjN1DapWEw7agRXHdRHqAEge+mr32RuySiNN
kUfJDxSbmctUdgzQRkPCjEouPMWOXDCKsBj2U5+zHEsvN06qnS3sbjUhfp5I5XFI
+DM8Av2DMGL3momw9k3lyfyOdg+jwFdiRWREnI1rkESKfKd4qLziw0G9lfAH6INj
vYUc6RxoPhnmDGUdHYlJn8/jVfUk1+qibOVRwE2qYrU6eBTxXvdMPppGitaHFgtN
qY7t3T+P1yFa/6tmmLEOqBw5w5BK+j/wUQQcvBc4/MLakwK5KM5sm+H5LUuR+nZg
lpYCCH361KKyhr+c8rYJXT8AAs79rsR4zBjtim/F/I7mVOrKLAhnq02okNCZIcId
uoYgGhEUaT/o7T5HEBx4L1yfIvcJ0c6kILUuxLu4SrQjK6TRJ6I6rK7VjyHH0OdQ
nrEv//NgnVH4YSwU1Dt926E5L0MTkcDJSo8ii/InrIGPebQZ2bFT8KY65t8Mnacs
+1Ec/9MGGBSuZ1gwUOkqS4gjNIZ1oO7d7fjA5WRgqQhkeoDDnjkaei3NbG8VLwRZ
TcNnGv893XnZyz6dq6TrznAJJCgIPdv8KE/z/MLCxKUsQ9w9oyJb0SCTEsXVz0Ls
Rq4nAPAWVsvhXs0em0P/ydWL6VQrSDSdgAW9LZQqaL4iBRUxTQ+kx0SRHkvbhzvL
vRudxGXYMBQlRvBpao9asZ9QNy+JcTTio/cHTDtoH89TPCLHSN6SxieUtry9NQFQ
VeKgsluE6ZEHnK+Vtz4oW5tMsuGdeO7ZgQQeyksHIUAZUx+uoKwdS2c0bSavE5NY
b8am+tFJjU8ulSh82XqyIMEAnm7Dsj/ZZUQwetmTXa1iABrJ81w5Ei/GECxLeeIQ
6yEB7jWfTKoGmX2oZsW7T3cMlgIJKLPdodi+QEvJmBA1FFt9PPMXy5u2dmT9SAXk
b1YtD74RBgP4yRGkUqVl+xXySMkd8pU5nGzhMS70WauZnyONDBb0uMpSKTnVqPa9
faH5gpu/HA/pU2nLzEVAPAMZaOoRuOJ9TLyOUdzs3TFMzR3wgHkl5YK3ze401No7
4RCJT38ox9sjd7HUinyehRF3GWn5iY1YWvbGmSqxQ0t6gQdt61GVC8svTwXe5HUS
LcSxhbW1zK6pYVzPfNjuBwfGJKzeichOXZw7Aern8GEjkTe18u3MORiusR3juS7z
17gwSbY8I95q4QqUHmwHsBuwl52p/JLnRCeQ4dm592/E4k0lY+axB6lj7ie02DeF
6i4hRQcLFc4BS9qdPoqZO4l3acE3Vygh3reXGK/5fhZVuZN3XRA5tCjuuJOH10cM
uu7R91BcwaomhL7NK8N3ymo/QokWxAd7FzONZEmFLJDfEkZSTB2qKVWy3PNy7uYg
r230Lw4dYaK2sWdRKwWsPwnh8v5XIWmFCqh7Sq4vmKJgE96t857TxAQfUEKeG8mK
y+Dm7k2370bLqB8ZSBeiU0JNQJYsCegGUnPHbb0kqBCjseQLC4cA1Ch+rPS3XNPO
oC/K8TmQKeIirwbCR7OdUsf7UWZNhGjfSDrcIwcO0zafd1FpF9F/1gWyqDs5tecE
EVEANr54K1zz6iw3DGvaXKkHnOVFQK7gvVaU1reJ18hz2Dc4wfOPeS4oPginxnSG
/XQ+AS06uGz+wL4pJH4lSgvOUpk9rAZJQg/HYr6ucNXb+c3vq89OLI0ZOjwodTmp
3d8D68KVY4Z0PF4R/RPZfiZWNldlLrLOMYpTCICVXtqXDMcZWNw3ZX0Z8w1AD0eW
yRNtZZwsvmDl7Yp8Sled+AQKAvv8XYF1w1o8SyJ+UvyMppP+Srh4rKMnMZfE5WQ1
NsSltVQx26v1zftxTKJD/T2mTHjA+7L1422mV+B+bYhwyTEOw8sDXre3qzRI61Dv
lX2Fv5AkYnsGymNDN3iyXkelfb720MkdhkEXu8L+gpZ+qVb3ojZCtb0RPpBCsLgV
ffqixnv2f6M6YoYhz30mTcjbipnCZrAIf0yvflmIgO+n5GA2A0uqXO2cue9EdwG8
bfxdGGWcju5/b4CEG92xPdm6Y0HAS5g+hMKXlTHyIixhKfA8x9dTUEWq2kLamEQG
wKKaVhI/KsiVVTrWNKrUUOROmEOxwyWBASMmKIJVaZQApEm2AjDfk5LWgKplVHY/
RALqDijpDWxwpBBAVQm5LiN38MHfNGBCbMg1+5Me3mvfhWqWQO4am3xI9WZLbPOb
4o+BAJNNwMDnQUxa8DvmzpLdUeMXRnVdmOuvVjsXamXzC4h/uubyb2CiXa5nVkRA
NIC+cdubGJ8C6JOdDaszpdIQwrN+i3BdvNIvzPqvtpK5cIWzRjg2I2U4GUVltWs1
30G9y4mi57L6a+4nnfIXGTxAGYrbq7ZdjwMHoiHYXRK+5iOfImqLZjAPfcc87eDC
zNLNsOADb9iLE349GdVylIP436B+fruLLJus0YW1fmKwGTFjyaOPoIb8NTbwNO9K
7eU4/nxF3LoVZyFinzwH7N1TjckGkB13UxfkJFeHalA7AXv+tUy9oXBNqS6TbM3F
dJK1X4SZP9y7t3J19x3HTbJ4xZd3MyYGdeK0Nc9xktdEh0sdaUAY6xUK8za5Bht8
Hug5ULAbylyc19jpcDRTE6eB0YppJIxA21NOa7F3DU3E7qxCZ2n6fdrntBPs4rs2
AWakOOHfyIfWGwU4GcprwzXXJBiny9Oy8HmgGe9LBgNXQULoyThHn2n1qqHlvOzW
fIBQ0rKk4REt8TnAy7UNC1Mzo7vgjJUksijpY2TBObqr2PCWzJKBwColORl6hD3M
ASgaUnjBGzYjnrj3So11KmjaLefr4gIrCFejexxvQs2G7M2mf2qfvW2dxe04Z7ue
/Mnr7DYc68km48QN4U9S073zzqEhldB0sk5hw8DZvffL33UnDCXXW/b+Nlfvq6sl
YApXRvFyUxQzQ7OkfP4yIofyk4GqysQjq/kdd3ieVqZIe9CDO59QclF2z36sGYil
mWdYncGGv2kBUffAJicnPiKiY75ewRtlX/6oQ6UARFI7kZL/NZ8A5IygoPDHe7F3
15b2c5nIvOjhzTO3GmWqxpk6UQKKXRqEVXocsnHfQoDgGPFdnqq+jMEvhyuXWZFi
Wa4jrhn92NMbcEGzJjZ/WkBzae/EId8sLly9AbDSORglqrOPmhMcA7NiVc3LjrwC
FhqY2DRgE8leEz4CtAl3jYS1xPk/Jo8AVk7PL+JNWclvxKLufYBrazeNjZMvALIG
9EBlaYGpDvKWPib84rLqh258rBYEDKJLfKs+g6L8NYIF6lOqijotFsy4MIjKdPeK
QCsU5V2vHtk8W4W/n2oxb/uBeA3t1SiJEBrmd/fs4HUW0O8lj3XdTeF+fx3Hrtgf
7ZGfFB3H6fDg688otd8A0vsAcTscG+/HRTscejP2nwZ1FUgHLNiHoSEyh1fl+mSr
6VuxJpPtKgAht1RfaJq/xmTIqNy2DnMKn3qW2EyDuCogj5R9BngwIlvOxprroyBM
D/OBtrLslk2PTA42ovWttBk02cgXkhqY44L1BvicNh6gpjcx1UPwU+8o0VIEaCz4
bA240AvU3iRnO5DkZPb2b8TrjxWQeP+2ANX2WXZiZMvTmgQKe6w6RTm7xnCbhmNl
165Db+NRDLjod1B2aWZ0EbLYBbnRd9zDAu9Up0k5xXr5r6qf2Odrqu7KmAMM1blu
B4hRukUE1P5G9mPQ0OZdr4Nb0dG5b1zMzbLVihe3BhUqFEbdiB4yqFNublrqhpMr
u9+dcjT7qZLQtM+0YgbkqhUN+imjLjtFD7AKfL9rBAZpSzXdMBrAp4ReCQtEzVI3
MpmZOKET+TSdBLcBshrkbsRsUZv/e/QUbkzfzaC3O9IY4ERGfYxI+TUPA0pxAO5v
Pz1EMglWSz98an6CX/mQXOa7/D5cG7hS3x42V2qoba+VYpvOUP1AWqn3CHvI9xEJ
Vz5Ke7bsmP7DiQdysIttO1Vt8vNLy8iZ014bUwIZKpbh6tiRnw5YXE1AtPUHfJbh
mT4du/m2qTLUesI85ugRuEwZacMGyYl+ok7PVgeJw1TfMexvDvi4azt0XgttwhuD
dpuq4ara+Upp1CeFupdzSoje+rs7YPEH3T4j7ZhGzlPO8pSnU/Y0v4ohi2LA5Fzz
PO7f9gc768XaVFe+TjqVu6ypemAv5iYN7GOR+mfrRmwENwWPbFK7cQw/8Il/RSAE
7FTobp3x4kOy6UYlz7tCo2uPtOL6G2RHsgz1jeOuPXk3pYs+ZCSx9AcIZKK5A14E
VunCRxSlYVDT3ci5JfxZd2i3HYzj5HLaS0XLLJSFa1mO4GEJJg2EnQVFnNshXBtP
DvJKMcsBNCCQMOPV/rccAlPGjXevxTZhq0Fnm2nJTnxCNBwdjUz0g6zh3DdF6a40
ZieXDQ4UUNvvjJdU1Qri3V1zss4QRGvrxi8/SB4ghE95cBPMQO1aiGpnlOCK0dTY
8XNAPVn/Y50v4LI8KHk0CZ0/ydHWGY1j6N1XgO84hMiia5KqPDFMgapuphOxuDtv
Kea1buI7edBzhSq4MUb30MxVEp25xq8QRRMgQe7pUR/fcCtT6KkOb6tfZubW5xNk
ZygRHamIkc/emSfozNGas+65Vf4Vn7it8v6AFXO+apEs6q9s5XCpmKNFBxPj06jy
7mqj1DAOwwffmMSzH/pRKohCVOZu2ZClhsrcPaO9QSzvB89vTKipp9BH1vv4MJr+
YlhzDbwmuiQsisBabVn2z2Z4MRcfWQiuW288viT1m4+slZsAsUG9QvyNOHzwqw5W
p8np/T3v+rqi8lYjFP5tyF+2lBQtky1xqOwJMPvy718kmXKxvAB7Lr6Po3EYhpjk
T/WV2LVXXcI0+vAERpNt2jMgYKUccdi+gCooiQXrIzgkdat/Hz5Jy+u9a0WQJz56
L4JjX15Rc5etiH+1bJbGdg8jiVy6zJMBI4pf8qLgPk7RNgVM0KjuE2mtYBh82X4n
SF256Bhc/+LA4TjqU+rHwCBCYISyohj5G4Ks13PbgrmJQtiahKte5AT3Pi8/SEoi
seaqu5UI5LrViRZQmPhSEvK6nNRVa//kgTKPfR9lUA+bEn1TD27QsYNmN2kZZIxm
G/iB6XdCiryDXACCPg+L4ThXxMHzzNrGprCiuYTtqu8/fQDD7n0qM8NVfMUo6pCm
4QJ9EmdC/ev05DF7E3qY5G6vF5rLIc4l4uFVz99/FjTysWZfMTe4HXSP4MpUmbSK
hmzO2fhexGXz58qXBRAa2JlnZNYeMnqBO0f6o6WiWPThcuNAnqf1MB2sK8owX/ER
AI+P7HADOxp6BjenkHU+zWW6ct8cPysvGk3Av/L66jF4aTdpsj+eGEF8vHQV7mwq
krlH+XCrK7VZtns7/eO57eC1LmQ64/9iYtM+dGPGMdVikvuM1DkADgCIWtzEYoHr
DkJ/aQ0TLcjR78yPHP7rExNGjSQG6JRjtBgTdT/REllG768a6l08FRII0ZfvQwDO
uQ8Tbxfj3Gv/r8gAVJVarBcXjZd6reUPoRyuV4G/gJNDXr5tjpSStHgcqbVGq+rX
3XuwUXPaJzId2IL+4QO8tiCrw6fknvn3i0lQs/x4YO7nUcNVegtO+v2HoYGK/U6k
XlKwRx9G4osRkUedIBkaIPbRJ/+gWcPn7Z8tACXPtLi8iJeiYWE42ejcnFkzOt6r
/koRrphk21U++xkkFcKP2NsFQx81GtiW2QdDXaA7GBmogiahTnrec5pzrsINvZY1
uMZmPfHJS37FSwQT6RU8Aejv38ObDjP6RDLPb5qsfM659xnL7ijVt8TBinUnJxFW
p5K2tcBCn2djoiQfZk9fBSZ/MFOERuf+MJVZPUHglcEBZxfsFXmwPy4p8FRNW3FF
KWx72gPu6aKVHOHfMnACIw0Z24XeEIpxS8FpAT1mrpAUENjRj/p7Yi3k5bKcU7xO
PvDB3mCX71cXDZtzYycl8H6mGGx2BcF8jDECAdBU4KL3WoKZq3NlfhjqKFOCKcoS
7d9RgxvnoQ8tl4XHSWDj9PLru7E8y1K+ig01WAen2+7bBmH5+cYBCJjOLkHdld8+
JGnBfTPkgLHmNNv5EjgmnzY1pZbc1yS8TNBtL/52Z85iMYrT+ikn2SIWnXkfDMYt
xGn8KR3jn1tn/5+XnT3BsQtswpUK9BQw6+Vr7yMaRsUi/udPbJDD6AB42QbKjyqL
J9rujLEkBs2K9ZZXsiW6I6plESOW1BdDfTAMmZGlEEr75/J2BObouY5Ihhoxbu97
D877+GPzeV4jbL5VHpcfMzwhXs2i2XYIGy3xOOKJaOOgH/vPmJXomenFWrZKv1Pr
iQi0I+R1cOtbxphw7Z5zSCOpG5aM3jnX7rv9MQvoGDfDw0eet1+3rr1RCYzhWSpM
J4yih/ILiq02iKcebnw6Xz1o1iUm+iWhR6rsD9PiF/yrGK6zbxs1mTVCMTDUL/NG
VS8pKFtvkRwnzaN2KH0nv/xoGJqRWpjWAwC7LfUeH7/wZRZl92Rn2e3th/WoaLXy
9Qqr0eGejatVY1OEBSPAoUCnEjy7SWhyQJ83TX+Op1zZCxXENBeZ4hiPUthhavQz
8pF99f4jr1Qmvtb02j+SJwa9iSSAR9j+cKxelBubLpi2BH5Xy5hfKE4/TQeXbBtq
ii3eOl6r5ovJnGE4Q6NB9t6EunQYwKiWN4wbtgjWI+oJxybXDMBgHgKnW2EVaXRv
FZWG32Wk2hFZdsC44pPx6eieFJPpDAn5UPo9GiPNYwXa7UuSmPNoW/D2EGt04hJ1
b1MMUvn276lMIdiWxLBi2zILPym6nsKw4D0eB7sp4KFnT/6GGKgQ2IT9r6HBcnPU
iIQXWp9he8tQpHPQjx9UNkXmsfBXJJmkCOh5ijByHLvRN2ETnfk4Sw701eRO7wHb
K9OZ5bWiVGzTaw2jL4e2P6caz4UpOFvrakSVO0+WlGRcJir1lqGMdyNXnPQrUurk
15vranyb0DECn0EOttt47pzs4l00WBgGq2AtMEj/aSEBwy/ROojjobCpXCuZqNRt
UndSXa+zV+5fBwlbXcwqff9cAS9/510oL9nLwINTVzc/YdnC8yI6xYVpB0i7UWGL
XgkUUXCz9blyrmFj9P6+uvcA7dW5yH+gQBPIk6ebjZ0PVxlorx+qLBoG6yQ1yZHy
SmpS0N4mYYm5hftZ28eGjUZoDdHxKQzq7g4JGf6Srr6Z5lUodfeQ8ED9DncpGydu
3NaynBJtaDPrD8ncNnLscV3eQm74BiamkETBCDSbaevesoNouhfVD9E7oj6T//q0
gheEvdS3kB+jlauZNkHnJ1vSWiOxW+jeWwkfmHH/f/bwwUJkIG5IuXRdMccvmy5s
Qi/rvQF518l98EQPIadWyE6FMxvbZ3Rw63NYquISuiO9Jk590MZOp606YaMHHnWL
6wlomLEQZPeEEank9uSwVhvGv7xCbiNcCqM92OszZLUdFOIT4Nn/zG5bpxGAkwyt
7sobHLBQgiw++vgN4C6NEvxjYUwQlqlKohwEyRouFEjHl4Ua+jKdRUufwOibJw4e
fj26BSp+NaaltK0WSeX42Csz41/df+6YKzcOY3bIe5guQSTlOIw9X8i8HXqUnK07
tYQQJWn2Hj34hA6LAw+LzR6XMcuQ8lVy9LuMnwnP7NTjmlgGVZWps2lq/yDZ884y
iyXSSIS1aMaNcjkPumkUmFYJqvQzMqr2p56Kv//TtuGrY6/pcSkrbTqBclfqv9Hi
hDr4fFRotE7wZUsjIi8OQc2tqZKU7j1bxJO5vEj5MOkW3+TwMMooRTF5GFqojcBD
aOdz/FNHH7o7wTAHDfFkeqzrNqbwb8PVfUQgvM3YjIfXhXePAJ0Rhtg819LcgmLE
dhyNbpIZrXaBgoI0D2Sa8UAEZa6jJnyB9hEfyZreA+9bQfurxiyxvdxKm1X1/nFi
aAmR1b3R1rW6U9Mo0AZVurHictgTUOHpmkTdZJi12ea4wERPMGe/SI0LteNE1ah5
DAhkaW3EI+7YrVxepxIYVqVkclp3oRHBulUj+5hW0cGVdcvRHbcZ2gfhE/O9OIgv
ny8Ph6TEevxzh07D7AXnKnwsJ4HvP7D0yH1ncG4Gbc0+zNykZYYyqJOxXyElvHob
EFjgucfzhKCRFlZeCHEpKgwEEPjbqaAM9hbDqyqOITb2BAQ2FquRa8lmd5l1F0vX
kDfDck9+6+xdeK9GDjeWGjILcB4UO/RaviUDF5aHHTMg8Kml/U4CvLv8K+GKUUH9
5ZmLzHQZRcRGv47SofbkAbOJzoGDD6otAEmmAjBAew3KyZQcbO20kxtXyLBAf1gq
XecC+XBRBPpSAPSwi6OjjGY833C4s8h9ttbKTLKTtHERQhcgBWHRJV6IcuGJD1pX
F9l7AvEircZlJdhuLmPXmydWStfIl0RAsyCHbBUI2QHvddDQwSZ8mGMqXYGYZlk4
5usM4xvmKcmCcVe83UKSpQNECt5qsYIwO2MylCYxGYcxkcAxLqOxMNTPfwq2IpOf
L55RXxqg1Fgg5dzVbepuJFEYcDPA8DGgCtDsSfxs2pF6CopPZ2qIqUpqKCxd/1jg
OMWfZfM7lNjMNQzGDzaABp2Zk7KQXe4c+uqm90uXG1ge6YHYskrdtgiVhSGXbOrf
+8b8xkHXXqzhDWxRnX4tLqtk9r1g63363N/u2Xt3z+5PBSFyPXH/hTVQH7wJj9Om
VfmgfRl5He6Gs/mmqlyQWT6e8i9deu+hpsQGxRBKiKXYkr9hH1lqdYy2DprZh7Qv
im7gVnSK/4JuSDxuvhchZISNQnnsaKv5w4FIBSkBP3tsc+oWNJCD0rdboEqmzvCL
aGjOmZn2wEqOR6vPx9JjoAhdlIh+WgxglMCqHah/Wzt4GIKO+oQGyaX3k+Z78WEr
26MbxdD62SJA27yjnQUjMFZbB/mcR2yruZO40DRcJehCf6l+0xGnpU0QO6pu1+rW
gVRS48BrpcgEo/X/D1CI0juAEn6yeMN6CD4Z8LOXccZLnO+/72xT/gKC/2t000Q0
CVpzwzSKVbGfSQ+9VRLjAQVQtTiNXdIf7jX0OcHrt4LpoRCv6K6EAP5f5JQ9ETAj
/8o9LD8nxmYGzCthnIl4smmKrn03GZ3kBKWIhSiCnx6aCcJjpgSe/CVckkr/U7Xh
EItW2BsCdJb5rD/zKbmS+gordt/cuc54RLNpScvYEv57O2RVPBwMGQHwH6nEEDYE
DxgGMgh4LXCsRs5/D8w0/feJJhXQdh/RYVx9ERLCnufBREI2EPMj/kNh8TjD/K6u
nQMFBEjjaHypPSNlDh1V1wUUCa2a131NsF3EQznAVrKZ/MOReGRvW3k0V1WS2IpP
QPOLFXM86I75q/l1+MwloG1V6USpmRKtk82f345AzJIQ1RBQlBnwVszi+yIZ3Ylc
kl/JY3TeQW7iZe346v3yWHVdFF4+tH5rTl5GXaQl7ST4bNt3TO346YJLkbg6ape+
2VJWYyrCMWfGnae3ztYCSjGCrrHVw/7kOMil6jLgPCKF9j9QkZyFmHoPxJX/RXwg
hk8HohKHwnPW6oT7m8Q8XTgHtPHTj6MWlfbZ31pDPi3I7AHwwgYi/+wN6Ek2Jli9
Imacj32ZSRVxze3klHQscoyGQTvA0GJ4v1rJQX2cCFQQGC2Acl23hG7Z7ShQM6H5
xj96nrG6GIKjF1clmo4Xr31UV3bli5NO3GmRnZ0i65zocTQDyCX/WFCBFeBcHhjx
2gZltKYe2XVYlIHbmfp1UE8fn1gIR5lvR8nQ5n8ERoZJD6Wcf4keeuU3LFS0w6ci
ic6ndjNT2ikK6gKFJTu7BKplExcIyZBJjVi58tkFzPTbm0azjcl6rBHaJoKgf9gU
qCO7MCS/jqL7D3bEjfpbnFr8su7sXr7znhsEq+UK+PgeaECq4cqFhxI17mExAjLT
3u5Bvyzxl26/znpTINFV3Mm7nWXera/fd36YAbGY8xwGHUHKpCYvGkpdx/TUUVDj
JVXNN4/O+lk8+anw/dEXV8Ia7v5SjF/3baXZox+N9eZlIfFHo1hnZZ6l32UTD7kY
rGjeWc1+OcTcwxihJ5MIqiAGtftOzl9FSV56wYrBdiJdOlZ34OoXABxlzBaBzHn9
vwUXjuSJ8Rhci9G3P92jrvS0rioNwE5CU2VfpYyGsaGQnvBlsY/rWFReWb1AB+jR
sbGNAyb4FgF2VL/s4GqFYo2UVS+lb3w8Ie2nTrKLcFKTLuzudAT3ki71zmnhnpEf
UUUNE4OP+egZz61woITXVdwWaQwS8tAsdmxCtpoK+Z+fE1v58p+EOJU+em35wd7r
ZBzezsjKWhU94CMDFM1C6rXr47mmkJc1AFMDNIUeRC+4px+b273KVcSwaU0+y4d9
h11e5phj4Ti9fgweuBIYm13dNeRCijWPCIrJ8sdZqo1CchoQeszQ3hiGn7kOvUbG
2sCuAXLibi4Xr/OBaUkZtC5E6yonBzg1tXapjQVmS3CsOVra+3wqY2W4xG7vIIi+
3j5MuECSb4aDJjYWZ5tSZHYVkDdEYy8k6DmBAQ2XDb/Qh0nfKTE2wkaX8qo4Dpf2
mqR4pjUel7KTcUIzLksGgizqsiIvFrsd4hYXL7DE8yEQxQsN2n78TjlwYjUuJR5d
0ifb5XcAzcYuljngX4eW7pyf/83d0MztuPj5BopmsJOnYNJ2XR85jFU1EpPTABWR
o9M+8Ik9BbXWWeLb8L0eSXY8RwOgvTCpqiMBE6sPG1JeOXh2rY74Ru8tbsmn8h7s
ECXAF//gaTr/0FawCq1Va02Q0atsg+LL5xdk5EF9HiXjCmhxQX+mCtiJoiN77Obc
dM8L++UnuIcvHhgBENhWobngFgpjZwC/8a9PTylnL/OCFRxBxBUAURXTxJ+HsSxl
tq5TS7ywVbPUtTVwhvi4Fw5LlXwMmj/0PQpK2lWVjrmagEQpEo/WSkrndopaTvaj
J/SFE+JqvuqdE0Kh03UzolK9e+yvlH8vLiKYIHvC+psDb4TtPytWLb0wpUZ2Kvpm
0R4vMy50J0Y/bNGCL3JB+wr4Bt0todT/aeo2aqLgA5AHCpzLIqXcvEvRypbtq3ix
0bWV9/V+51Dx4sGdEj1IgsAbEHiA2oQZAILcSIiLpRMc4WuaEknXSko5RvU7mKjl
YPSr/pq+9TbsJIUF/NfFJ/6cjF2M+3Wx5yQooWnzoG46UR4sgbNGXogSKYs/i7os
Zcj5PZI72Q7DQx2LFetajzTF9Wq3Bpc2L9xfLJSYkgJ9akGVY25PORIVwJn2ZlvF
DFmvdSpI4EdkqSElUxw4gLJMjk7vbvfnwWbZoez4E+nj2YdkWjnvOPdYS/ZnxLbo
RDPM4kgzEnrLVxe5aRz6+2XIw5s5mUVVZPHkbm8Kf+WsbV5ZeEfcm0MEFeTBeN7Q
DSM6CE6G7lhTO5HGb85GBuH61cWxbTViq7R753YQ5ju0G3uSy1XHQIJgHUVUNDC9
Jxg3ae4nYv5XWbqWLszKQ8vtxu4Rrz9Se+cfD1P8+Wkfgda1AKBRPCwaqwWYVpPQ
jKraQ1qF8CZcPX5fh4Na/9VdRcLetQdkYYZ5NnCqC7SiTqc4VPLc8BBgNP6OJa4y
b/z4y2FfSJZeX3q9GzoFWbJHNfSdh1jTSKrMpPfRs6bAloMSmdouoKnGtl+CM0UA
kbOrAuDKuYb4BHOT7dugqBQkA71sE6h1YHHmR+SDzMUu6cQbCg6cly7sMoGxGN9R
JYJEfYJ1Na+jq3wkTDnHgOACN5XjuefvxDXmPawC/nmqy1Xpx5+0NqzgJxfz+lsX
wAbc02jzneSDVZnImtnaW51ZX/N3GSwSgErzTJmYSvrCnQ0lFe1MVPVFDizy/UN3
ZqvzxOa/kH2PEvkoz3b4saDf1/EtQfjIAPtyGmu7McOb5rIrWst9YICJoeJ6g8R+
DA5tY1l/vucyCsF773s/zv8nj8xQfjvsMqrC0BiJ6q2KCehiovxE1G72CcOudXbk
hJhwd/y4CrYz+pBut9jg/WTSCu8aCFrHvLZqxDBNzfSQ7B25+FJj+tpPGIRIPINl
zcOkQ1CGPeli/qnLbR2iJ5U/p67VIWFnR2QGwCezXO4ZMD/PyZp/3f6xigQTI0Ia
bdOe2PWI+J9kE2jkJbdPxB3RhvH34RTgE+36zTwmaYJUl4c3uErCZVFCFTYlELRF
1LWnR7g8icMvoWcAqe/TkfIEKLhRqYqKA0vT7QU+QRtdAhY+IFOF4FjKVN/t68Eb
iDf3km4Cb0ZQMk+xAJZOBbwP27o+LKHutHO7YrzAvqiCOVEqngyF3Ur0NRQNxf7M
F9WsZNo50vst4PgVwjFOp5bM2rUL/7bm5ZYevpHsV+zOi51TXQPDbQuYm9C8kZvz
FoXI5AdoKzXqXAOVSt46QZnsp9SD6yfQoOwPqdXYezMtIYq6scDT7v75u4rtG4R5
t9gBMlkou+Hwu3VshfV8Tjnuy6TmjlPOKPyqGguX3uuFXmnLJMX8j0MbaF7eEhTM
bQJXerLxuFKBzAL4iJs+kHAFBO4Y817//VIchl9zyHuXPU39ITAhXmI5+xDwy3lL
24NzUIFFIVThuyR0Ebr/rlO5lV5VUYwrShdSnGzet5F3SxnbANdc5IRum86rhcE5
x4cQtXDOYh2L2nA3lw55224uXw/hX2mWDK0Bd6jb4x6GzRfX3MZpQfJfGOBTEpS9
+tLFSVmzLiz+245GcI0IfXDXTnaIKhCEKXm2+JsA4YDSI/xtg/DSVAfv2cfOWNfm
4cVrVibQsmNrR1yjKoNFknXPbi82oJoJbXsYN3rgMaa5SJCZi1XR3ViAAoDsj8wP
LuF1Vq8eZ8XV67EXr1o+rI5RTYC4kVLvJW5nwCAzn9U8ZOxrrgGXgrHEgz/v93L5
AuL3DB+qcvB+VJofb7m2KAi8+scD75ialrVHwuT7gP1zIYwhxXvhaIWgqnsA8ndm
l9fOA53v3t/dfQ3LkyERj5pIqYR7ujsWjo2qhiC6KuOMr95VIHhQCrF7l24oz1g0
mjGdwZUShH8Z1v/mNq4hKZCzk6x5TeaPLKBZaezeuIX6G0+IP4QU6nLQrIAyHPXU
o+pIUpnTyvl69YJcvTulAjkFXTa/A5fYus48tSxq/aeM+favgHwU1vutgnONmjBT
O8Kg87SKx8SkDAORxhY68Bl5ooLjgAD+GPJ29ZL9j6k=
`protect END_PROTECTED
