`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FNa1GkiCJ1D6UJ5jQRJRFzQpHolZz//+voULgsuR5A6A7TBkY81kIFFsSUSWeN2b
IBJnEoJ6Js6opUijnBGm7ECjwIHUB8rfpnzY4gYXoRlW6ilt/HAyOQO0XIatYmW6
l3BLuZwnGVJ1Fj6CVeIpNgGrRHBCAWmH1kp8mtB/BSER8eh3j/NSCPh9Huornd2+
MwuW71530O48drFIlfBvViabwBBOTWrnrwYOza5Zfd5saucJkBwNhgnCLG8G0ZeS
dJZFW8Wec27x7hrEPbqRLILv4CDi3FBIcusQdqg8+k2BAVQsrY/avuflHDM5BVEX
xQISTA0U42uLD2hb9UCvevbIqe+BkZza35EoNFP/Hgb11p1B5dlsf+PJmKTLaNca
6wYUuju2ucO3NzvKUnRCilQg8ALMzH6c5dzcedCNmVY/TyuwYc0+oQMq3K1CPa1/
rWurHPstrstzAyPDaHg2HQiXEw7Y5g2ejy3PSX5PYl3UD6hg57ZmOtXnV+a/TDHA
3jZrPsAA4UmPDCU29OSRf0xGSn+k8sJzl+rnx7SGMQlH601AsbxA3hwd0e/e1RQA
ryBXLV03QnrGk1v4P3gI3ikzfF6zD25mI/0D3piq8do=
`protect END_PROTECTED
