`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KlB2nZmJHFd9O3aUXZuePmIk8bmv9JzedRb9w3IQuWPrdBSvZgxVXuhkMTaDl3Or
Ey5pVqePMSuTG3VKTG+zb/N49CdvTIrZFtez5bmn66ja4zjW2cJlnNipV5+cUlbS
Rpx9b8u8vdAok7O2/+Smf/8QUyF+BbYVH+qwqA1fsP1bMbZcLTzqYSXziDlN9Oi5
DG6gQJN7791x4MtTaRuhogQ68Yv/VUfazBadD5DGCYmkAakilEGTL3Owf9iYkFTt
k5dwqb3T6R+n6MQ+4aq45/mXdbVsxU0LtX5IpkM/LkFhV/KTUG3JFiTl+F1CXaFz
fnOTu1komm4NMiMfD6sXdduHECX1d/ptW2dS7MwrjCetVlMxIU66YTjM5MtDEX8M
9gwU2r5I2P6fH/T7/EYy9l1nC/6IFBTBq1oZc0SswoUq6Ne/j38kWegRhD5p61TK
1wmViRQOFcm/tZIy3f74MHhfmWZ4lfw2KUF/LhxYRJlaH37I89UvZqvCTGPC5GxT
BK66Ldw4ytbd4VHzW/lYrXeJSLdI869/Jz5auV3kwRCIm/TUL+xe9dUDkJyZJiTY
nWY6LsKnX5Sa7sNK2OT9aCKn0F2zUUUaElnxQXZWVmAl99JNvWCk5KzCbyZyvuIc
pu8zwEOKWldDeeIctV937qq8LwdfH+n5osfgjKdVgF1wllASof/BXEQnbGxKe/bR
6DWoJo5q1drH6VAYZFmBaXyHqiZYqeO9gGuOLYGi3iwDA5APhJMtgvO/xCnCF1FP
o3iEAP9YVKFuF8cKs6ngf4YSbJFSjQY4i0+jIQjYPcp7GdZYqT2vwSh3BIRRwjns
dsATKjyttl5jbvRNjeUPCKIE8iPMJwfQsNMs93KMYEh4fyxYRFNCu1wNPhZirm+H
3c0gy4YrootwP70IgEd2bv975KMTlyzowi2MlC0lx+lbgSkHxPJHXTc2NAQx7Wyv
yNwOP7s9mrNbfR6h54yFHNsiaLv5kSbIxVdWyw22w8zlKFMD8HjPjMjPGMnZjPqj
unbHap6BMrTxajL7qgwAVoaA97YPrC1hPfdfla7KDafRXhiWD0Mh0xHo0mg0iK2k
JVlCvc1QsjuFOWjKSk4OSqeznvl7Mm6tt/w7VhYfboKrjagjLBwkMQNXePmP0eud
ZitMbAkDwLjxv3NtvQmFN28vn2hgkdveu6fkcgFUA+qAQ/wJuhFnsFu1ipDTj0Px
PaWFt6X6dOp4UHQvuXmD8j4hwgD9K4EJZdJ6Z28/Tt+b7HvtH6KiqBQxCt65jrJC
1mkZRQifhoLCsGEbYht1PdbR0DwHpoMnumhnHTmwUaHhLcS5gV81YmHKDYERTsNE
HOGPdZRFH14DRKtSMFW/W4MDpZXFsjgWvMjllqgVHtIYCiNH8Ua8QvbNiPnkxJdF
Y6BOn03oaI+9GaGPVA65moO8tEqjgemY6TcwnjE5sBSAszflidaz/LrTknNVWhs+
rvCrEnxx+a41wUQeg3b5QiPMRl5X+an8EAYqtdUigVUc7cRIa4+NnvtT26vupMpr
GlDUI8rPSe+qFPtwFQcDOmcVPYX3X6rDXZX2i/OEnLlVp55clPeuBfy8QXgl4dWK
2EXsC9eTtDc00laa9BsjD9Syu8QT+6h9j4/XK0JoyfvzfFplwe+HxMfYEWsXLFd0
lrq15ScRWcGLvriwrAhJVZbLI+68Ls/9v1sEEFn/AkEZ9+N0GD3ULtRnSQ8uT5Qn
LP0S5k4uhRwmr3pMINnrBg5/QAFgJpaX+SpwkFDxYCgxdTC5T1HY2XE6Jw4D6RYF
0A3Pnm4VuIKM4ggEv8s/dMN1CuExqMLF1eTvw9v/rXIRlh2afx4SGHOgePzr6l+Y
glOfB10pdrTRvu9gS1mazKDdwircoqex5MfYEbRp3ZWJV/+JKWCGeUHv0JNbwygS
UbSsE0EEZSMPK45dEJWTFlU5t4B3pIRnv2V70CW9vmZqNJum12uGbrgZjvRKZrjk
cgrk9ePMt07tomg3yjkM+sUZsRT0OqlpH1Et31dzu3eMZy2z2TyWk+kVi0PDcyB6
yAGBNsqrpQl++4ac40QuwlcwXNGvksMDJ/X6k3xhaE96RhbM8Qcc0Zkv8qwgnJLR
ulvy05KLZhYl+DkhpQH+WLR/DSz+CC52VRH77IndPuHG6TChjv5Pk4gSkQNYDPjb
Q9v0djmx39iy61VvoejEp8VNXfPe0Z9hV4o7cjVjNb06DyLtGFXnFy9v/75oH4FO
qf1w+YlSGPqsENV5z2jbvRD4birGRcOhlOq1WOMZNdrZXE/JvKL3S7asb7xZMajX
I0Xr5hIZfbPXefH0HBZe50O6Jxj1xPEoB+n1F5mbtkbT/gi9V89bUYKWPNaTlS88
oPhymDY5wR3p6H2QtrvuhHHDIzn6xZ+WNVVxNmdpvlhwIZqHCZJ8RgXL/CrOvxj8
HxuoTZsd91IcfE+5jVC38+1zxt5VepXErsd0nt378whQbbxjtacHH816bd7xk8Tj
0dCIH2PGZtYs+tY2H3Jpsi/2GmFXX7uFWIs/b6qDHkChvDfT0ouOsL9u/QTUiIcC
UT+QgNS+KG/oTCBwdkGjRHVXYTtv/cKhLW6Zf/qAjTxFvKdOuZ9G2pN+eUWCGRff
t22amzzwPjJVj87/he1bsQIBi2xyINkIzwGGNjdpJPzrfbSZKMPA4DwONZSGv3Ul
AWQPZ+fM3kjwPzO7x/OavDF9BwlbXe0lnyK2KwxvU4RtgKtca0wybvzIRpNU6YWH
gZz6zam2aO6nO1sh5C8130Phijjb0BgYJSD+tc4BLD63UVUkehDtyfaZj23RS7uU
SmUPc+M/cpkhbybfgWDk5Qfw6SoSvb3dy2xcruNk/B84Sz2PyZc0YHXyBBIYSWND
A24GFMaZShFz8BKDL0/k2YUZynpFvPzkVIjbdCHa1HiVSVGsVpi9e4jfXrZ9fMj8
hl1k7+uybHDUgoPL6W1gro52ma8oVEv/RZAqc6+UfjCpSmUq80WsydJy7TabPCHG
5pDqwdUEuI0h048lWy9HGmKb5Yf/Xd1lBvJygeDk63h+5GR/E61K1NTzLiuCYe52
lnQ4ZIdvMHidEWWArdYidNuYWnnRBGtCElOetritIucy1bzqjoy9CJ2ujYRmnGjy
G65GjOb0UTFOXJDcPh4Lfep2ITaaIWoy/9wlSK4BfKxg5FObba/Lqm6j7X7n/Up/
PnCcCak/JbVjnVoQUtTOxftnQgT05/L4s9ihsKL13A14zHBlCKQY02RUFVFYVlDn
bVj4LGZdQ2l59ppXz9W3/sZjhCHgzoLuwPblWHKUNakueseypgZRY67SrLboGtaq
8dCY5uQOcrmsaWnV+9EkBwQWiUPIYSp0e0XHS7CnVJfaiDOXOskSpRmVbTf/12Yo
MncGkY88N0BhIbR2XwnFB9pfStmfCiPVpTZ0gj6fEITFrua664NAs7Ip0iRVHcZf
Fk/YxTkpGG3dS3ipvQ96zhjeD39naCSmlHEddT8pxLL9HdgkcriUMF/cpr7xWYSW
0kPtjWWNXOin9e8CvkBv6ZHHixBzMIyVFZw6MlbLtPrn+qY7WHKzx/XGZYHyjGa5
5yWW3HdH4HowTzyoFnT+WPlPn5ls8TR/i9JpuyZB/7T7S/gca1p4yCG/p0kPV92d
p8qaB3eK0iGG+KIjlLDL28Jh4/w8rMlaIkKo4R8nnOt546Vv/UrRgQosZsAVkKOi
HtK+5k6XXigB3232VRT0wXtfmgESj/XB1oVyBcYVf5VCbARFLCSDou7wAVrD4Wkv
a/ic0zwkRPNHScw9j2aOxPUVzGYi8KU7EtCxA3e0gAk7/E0CoJYBvFF/+4nIuq/g
4UYisx8CrodMyAINg1t0OADHsWhX18MhTckxwmbhz8U6piFGUW1C1smyb3Oy8Xq9
MzVCSLHTI60Xgg+dDRLl3m5BdQu0BVODNoFifptilGQ8ZZTuCgf/MuX4xsBSLLa3
eGsygjx+IQ3k8lHjwbnqj5DU+5aVAgl5A8yuJ9poweDsjkmnS9hmpH1TCaIThf7O
iVzgNBLWX8D9r0oTwRGkvyY54g4BElB7uThNXn4roBFp716/PSG+PawY9D8OHIYE
dqJCwIWKuPHs8sbFy3QMELo7htsFFYs6tzFDzW225dNlznyQogZ+Zt1VYSSNlhIf
olj7yoUi4INb38vdNhGzfGZnI3dKH2UYThWjNYYXzXiMr4ydJnU/gr5EoZPIBoR8
V8nbkaiciEBNEZQ9zEE6Bz+ZfJa21eD3wD3pKO9crNaNZv5JhytFXhOvnNeHf01y
+Ou7RJEig6MK7mqn9P3T13k+AQZTe3KImMkOrKLn/9r46WJivBD6KYVIOE+2Nuno
VZ1GDzs27jhpkEtSPmFciW8wddYG/9xDoemaqDQYuXQVM5pwqiPfLqEEoT/Ve1ra
DLa8M8luhyJx1NLxQEs0Lf6yJ9bRzVHXsQABI35dFlDoj+DvISlmNWJxxTJYw34m
NdZFIE72VEDMcGP4xBDoxHyDSfptDSNIyAXtWF4DNnPjbzF3RiRIbssWToaUjiHZ
UFoFmrlTtiwAl8woS+iIIUsM9XG/D6eQ7pNfWoEXtBsPjPty2Q56V+kT2f/lievC
KjvPDnCjP8Pn9HxJzeWD77p13oxydnq1rCnFkZg8o2AqKA5PfV0OJ8n2hvxJ2ZG9
S9yS9tL1XFziaU8Ko2kJQomVuoVB32zhZ6MP9ip5aGoYi9k8EVtJLVRo7PkExVYE
2txzDiWxugKjkMKfozCflJuKMSeuyNhHKA2yPnXwPefnO3hZVv276ibAEQLLjyJ2
638yWLOJKjRBzx2GfbduS4ud0P+T93yXONbUTvUjVZXQE3WqeFdz1XV4Vr7Num+r
t98svWfZ2RnkaWfBuTSW3J13GnH4lfbhvvyTNqAqTyuG/HkX4BddESrKV+gWjK1E
SrCsSZVIP1eou6osdxYBoiv/4utHlmgOMwyNYOqf4wCJ08MpXqIVkzE3F4S4LN0N
TKPHE4G52ZrmMCWzTZ0xISAgs6jHh5rFzSdMlWZSHfydKpxC421Txqhd8zb8LFVd
6HPYbJjiNwRI7au/ba3R5XGWqcJvLdR7vlkFhA3O06I3KhIxvIeQmlx0nJO9yciZ
FyJcFYxhL0f/MZjbJ+5mdFw4Xk2+Q4QBrA/6lx/WXi68eKBtSxBGaMk84/TxWadZ
xaVrkjkKEr2rMpExhjkK6dsQsE1+KTaO9P/Pw7Gwyts4GULlXxAXdwjgHG46cd2r
tmh+yExPwalwNbwrm5UcGkghMt/SKK5sMiGN6W9NDgFkRPDRpdEi6Lc1CtIgFaYp
GF05LEMeovTSGumkW9wXA+VYwK2Vjd0elA4Jx9SUuTpCkgxEAvffhtuu8CnN44Nv
o3gTN+aczvkQ5sUm5YyU6q/a6kqNiu/KZcVwBFMlu2T6OqHW5rxavMi0UL25ivIu
YVrECrCwT6B0aaGILoSuGh1Keyjd3jDx8OHflkLDK5//DRItNk4XDIw4kh7KkZBr
mZzIGRZWrJSHHJ0WTZ5fygonUjcS6VDPQ16I5p5oNUUMKjr14/grSz5yysScf0la
jvAiAZSkKQ/AlV5pMi/oLnlHoP4JnnVkeWYmGSd2Y4syTWzeofL5+tObWwFLXEh9
cAPSyNTKc3Xso8JegamibdOFNIhsuYyFGaL8NqNOzE1VnMFZsdDIlK+W3+G+2MJd
O35aZbvWAJg1WU/1Yt4vppdRPw2hDSe7BVZju0BCaQPDsUbkf2OKYE7sjJ5UvPp/
syKLQ7HVW3lFtjcjB6BIKe+w88JvfhgQLU9e12/NDATBE3gn0MH+PhMLEOWrXl/0
ySlFi+/8lRqnuF7FLUvALpP2ym0eOKS/moCxRpf/s8bXqohXjm68GWScEWo8pdqf
0/uPtLAk5rAAzJW7kUINsebQJ+Bbm8PRIJRxT6v7WB2OZYyoUVnsrSG2H0SCkL9M
NihLIjr0UVm1lCmk+tSwciWSN+B9eP8/ZazwVeV8RwHlQ7VWAxH8TKPE+AcZXACy
uH1Dg1uO4cE8FQa2+cWa7Unu5cr3FSFrbTwu56+Rz0yhHLj0+SKwWdlOKig9hque
U5wNp2EVbIOyDK76RCUX1s6OKBvf83rmkySjF88PV4kb08VC+EIDfRIQXrZYa52N
IRC0g5Xv5KsuVL5FRafvk5Rp5VqKu8HW8IYXFBeV5mMfOQgrfOhR1DTjn/IRmgV8
6vM0TUdgOonhQNGyRSIdIjx3dl0Qu5pXJzRgkCbQBr9L1Nh1umZAF/ypGrTMD9Gd
V0HdcZZ6xu9S1P/u7yse+gB/flUtU3fjhLU3KrmD3v/JJ19mWO1Kt52c002LLXdl
1iYIq9OLVXvvK+QMlzIxSlPcvMKp0EG3GvYcTXul6ktSWCTG3wR5M7XUdb2iOZQi
3O5sKMtjKWkebdvjqiCoNX42HtDThPS+8EL0RN3O5L/cRA1YKhOeBZun7YoR0lVr
ZWKN6KUz86PUFYVHZmwiOtbeRu4a0vxl2Ogh0vCop60/zV8noNiwwcHYKuEfGHmv
TO6AeXxX0Kgc5UWdrLzXa3PeYb/j66mn0YI63X7MIJQtgFIadRErLVIGDYum0/9i
nICq3WjasMEGyX7gq55kgODzwK9HZrClE7X/i68etdwai3Q4TW2OlnopKksrDXoj
7R9WODdnQBfaC6VTYSdLuDV/fXDekri9ZewnwqSfBzjfgke+T1RboIYbdQ+YaiRS
ykrYd+WJzn/A7Syg2+ftab5Lrnx0nktvcYavF+XWkuCdEbvqVd8o3hzUrA9INk1X
jwgmyifLN+fSCDsdJe1HKblsCL249piqs2Mvm7KtUMDnT7Uxt2frrBmx76vl8RzE
5qw+dsEiVL/E/h+668oRzkBl9VV5VdscZc1yAtwNKNzVOPtuey0AIFDFk6JfyIuB
jnEUN/qAZOI44MGNNpW3K9ywN35tafM2LmVLggn4LzOoT/Zj/xvgdhrazw0thziE
zhH/Wlqp4fU4yI82dXNZfHdx1bAWplb37fxTMaU5Y8198+On55M/mgEj/ispxjQx
vRi8oDr0S4CXopsNy1obYU7nKX0oeZlK65JI/S8NqfqfnxpdSL0RfQRNoP9dSgIV
zv/A575lJ1wYanbOxjmGyiCjQojBwL3vCHlEqw6LgpvvRtWLC1xrWAED5o0clEnT
GwofCMyEiS/6bGC7AZUvitkJ5MQG4VUkoooFaxPVMvVM+UUmRpuEHx1jFBSXvlh4
Lhr/dZCIkPpa6Kr4V+/UDWGLx1WEe6Ahwm/LSpQWe0hZLq+9OqCsYn3wP2mxAxCh
C8FSkDDPwzlktwE90MHbG4wPGI7JeUkDDXVDYRGzUazZ6RNF6FiL8dX+TELIxM69
NWa2Qn4GGNu/gk08w21yqOkUWfrUEehVMbIAsG0B3YMKPGNGOHwRtg1CGOoUP8hC
R36XetoPwt/5MVzcc1ylAn+c6gghpK6pFemOpQsusfCiDse2TxyA1dTFVyW0ZJL7
yFYsArhv6/nbYSZPAekEfLwPzhk3fhLf0FG0U2tHnc+nh2MVnO6Xb0mmXLnR7qms
aeBvPSmpAgfG/ynVRbAPA/WAWoAMSuZoGfC8LnHdQvbMVnYL3kgJ5ZaXEPkMH1X8
zcV5yvqfcy9gaFRld4CjmXoWywA04PSAp5bRl9k0QbwlzV2ofHcPe/EnYyvuTDWU
UXQL3kfU0KBVR+T1iuDrdhvYrFAWRGRPvYRzdp+nWQXPVGD/cOxLzwXMjI8RttJp
8SEEVg40Rj1fw2xUmqLloOwYgwYiUefWTmTKnjWJLwmHlAMEfB9hpHU5XiP3CQe5
veZNJBS55lqW97cyr6gnksFkNbcpl2pJwEndEsAY8jeYv++WChFZ/bFzb3gk8wCR
9QJgLhl0KrARRdCVmhNVCtVQezq6e1wWP6LEmx8AyRBwsPe+OInlnM2A7d/2eBMk
Fw13ShiUMXeDk0QHLUJ6BNAZ4FMcj56eBosAlu+jREp+5WLO3qsxcv+U4WCp3zu+
URnEjbWIUrN5eKNqHlNJ59WlRtvjhCQzIN5rm1G+NZHF7gf4j8+SgB6oG23SoKfk
ACaohd0RJdxFfI3DSZArfI4h1jzBLh+EZxPuVJ2vKJhsbprZ6YQ6tuE2oVpnnDaX
DmY8M4dXTxFyprp2kDM/v71erLaxZogC8SaiY3gLnf9tM5sSKqyZvd+3tuOBRsuq
XpEEAJdWlOLmLDH98I+Oabs1G4rdwTXiqGM4IXPaWZiab9Q/mcTbpvw89stQD2Pp
uwu7rWia67Ujv0H7C7MAFr/RjVsMQF4En/eCSiVYUxRb40UbyoYzfNu3QE4kH3GH
bJtUWV6dPXy5f898t12CrreCFLTSGM1zylsg+XZsJBBlSk1zrZ0uQB27ixWRgVBi
HIrJGYY+WndbfIZt3nWJ3rwTGu0VabpDcEllmfQg6tZK3jLHGzbPJHU5s0UPWdXX
2p/m1MEk/M+flZU5J86yyQwfI/b2EfVnEdTpSX1bXHcN0XQP/c47UxtEquyCxmP8
e6d1i/i47Vh5EBJ/KiP7wE5qqu8Elq0d6Cr2B3HZb8TCzACSe2v7fIHWnX+B+SJ8
AxL/6cw5HrNgGF4QS8DNZCPs+rOZUrsp6L29yDNE7sFvI+rZo0jwQZatZ4zL0WXP
Fzmc6b3ipa3wNwnROQce7v5bzSbkFIJurCDy0pLaDYaBcnMeJxKL77XNfW8SC8VB
uUSCkxb56v44irQUosGsvYlclXcX4WKhiKO8dm7mdFsskXelmY0fkCvv1pgclpKW
aZ5o7iAS4SeVuhJHFCGL1AgpHOglQhh88/C1CmTT3rmb51waOJ15Ra/SA0fvFS2X
SIPaPbItHQqWBl1EgOvqGkMePxEHHTywrkhco2x0rDYMbsy0ZeTy8eRUua3JeZok
a6yOgJdlu/0/scX+6ABKi6BuMlwHnLYoMRnVgK5jX312SFa6/R6+nlgUaaFDg1Li
3i8mmce2H+uP+GJ0E+/rVc8MopOD0OHexcSxdwLnqNtuKra6UneSCv2YRCMQkoJt
5J/T6cZ9UeDFNQ+KwtpHzVL10qFaL70DC5pvdIIbIlfRgHt6L7UA0Zgwqn7KcDRV
jIXcEnByG9JjW9aLkQcgevX+XLWFek4szCKZAlf1MUs/4iqYzjG4GaufUW62MI3i
Hcq1zy8uoDD1wzLDd7eTnu0/EMhLK6fyPzfIdeelGC7CIxWbax3fY1Q7Wg05cl2/
lf0vh0YJwpNBGCLMEz5P3aSsUp3miM1MpBDVoYYdkDz117+W625WMXt3q+MSeVp3
pTkZEPVlTshw1ExAEcy3qMec3C77WFCeL2H1ABT77THckU8HcQ0U3TUCGfnMJjF6
n7raiclszDb+IkqmrmTrAGfpxdkawTMk8+HZWKw9AgXbXbclhN092NvBWFNbI9AI
nHQVChOe0FPqv7zZzxkCvztMG/T1zfVTRLfhIe3Xmh0URembo24Ehe9HHrQgVEbj
M89CxFNGa+xcrTxkQgm/E6qtVSuGTjbL676q8d8tYCmhNKVq1Af5wtbignuUbkV0
GByGF/MkIF1pvlYMHSnfRoTd1bQchckdx4u4PGXZmvdjJWnQMGRPgL+j1X7Bd0u1
j4BylgDGvHd1BdRsg0FTq8woAD4Yy0eXAAkZoDmNFrfcZBOgyk3Jc3hXNlEff06D
DK+HTyaQF4KnKez22MlyH5xpjGVYwVV0Fwhker7qbHuxUCOiAsMTeG15Eg0wHf+z
9xVLokXsCzx7nv0YoB7kPbmTA4P4tVqQYDoEYmbaYYicExDB5NX333RWAWe2Dp0O
K7Q1cSi6EQP2C8ZGt3FkjHDDGao8YhGYVawFjboSqdnyKbHGz/0sxXrt4SFjkCIC
gDMQJN+zyWpUQ7do7awqSj91c7l10E+PLecV3+gdGC5AGLkvFTH8dEFOMRIR0t+1
jb7RWkv1WLdtmhpWOyS6J9vbelSJi+Kq4aK7uwXoslywaGT+0+MEuBs7XEmT+ErL
0hVy9/Cq2zdc34lY361BiJQvD+i5bXSeV++yiJ6hWjKs0bs41WUrQvIRkrkToHdp
TVA4GHrGHKnTnO5N9UshgZOkQDtM1KL6WtSTvrvytZNg2pTGqx1DnWYknWrl17qK
/Hfug+SnrXK9R5+smles2d78hiS1Ny6mL+O57NEPExkzel9t+dXS5ezSd/778uto
kZapC1Ls0kT6z5+OAzlRxWkRIGxTWOGO+MotpmfRzL6Giojh2yF8BmHzDOm0pGlw
RJE7JnSQnGoXgqinK7u3wezfm1nEFfbeYZj7tDt/xN18yAhXPbxNTxWQJcZuyyTg
M1G+nB7QIA7OTN0LBSVW+pKGAKWDZQ0VliaEx3JUu7ECA0Bkr9FDFyFy6H3RRfuS
ytDJYC9LhLOxHBcyFo0ZC8XZJHjMz1dHX0wEBEh20ZNuGxoCuUH+odlFdJOaZBna
ymnq6gMym/bQdBsLefiwkjcMBZ5pcH4IcVeBdnlgALYL/jZwalb826cLnLbuOUTD
9rgkDQ6UI65U5eGL58YuGvxLRc32TorWpHlXGZXQ19Mg4kxVdbYFIimUNSzLrMa6
F0I4yQir+gPkhlOXRrXnSfSpERfcAdbEEI/44S+f1K5lJ/lfWZTvKVVzwpNJVNhS
IQJ/fWKoRK6EsdQcP1xkjK2S8NLDdKxs+F8P6KV9z/BftIQOxpBXO8L0RcFuIfar
eqLTtXd6xvvKEHFosTRwJsdw53FLs8XTQwB/Sb93PaxpHGQuMR+nAxW82BufbzNk
/rk7Hx2FCvcwEr3v+gmnr7BMNpTaiiiQv/url+p9UNetd+eN4mM2RGWJoDsdPWE0
kfrHE8PtGYAydbpeYdfUf7uNSDpi7uY++9dofmlZpbCiL4pjxEe9+hQGrKV7KjDT
Z6PQZMItY9QcVNNPkDBl22BIfF/RkuTXgP8J7NT8ji38s6eKgPqeqG4RX6Yt41Kw
0RXU+MPsaf4JcIR8nC1CvFUti+sW+64uMJX47iFxglTCK7iSq3XFycvroxW9Zuqf
Oikskz7vXlqGUfjW5QcAD4olF6Ch2LL4nZPmR8QhaLfqHLQqfH1EzpTSmY9jVgCv
+ZvanJpUHrCovsGFivpcMXOzR1iqdWXXq63nQR30CUTCn8XcHsvuLvSqj2XG0DG/
Rh2z/zZwhc9rsGBg/j0DgmSlVe+ht/QwPKgdoaVtuySSVp9thTv0LPXFIF5i8TJJ
HxaDbXh6/297ViWLcVJCo25S0LlqBBp9ygYDUyTad8wkfQ0X2NILDh4jB7aRSzip
qo7gaUcaRZTU3mzfyb/RV3sBs5I1mBkj6WVN3WgkdUcMSMK+Y8QzYtrnAqbhuFYh
Dq/0WXi8Q6mIl+mRSL4MiTe7Q1nQssBRZNo47DMaVpHjZCc0JC3Fk+ZWqUfDubzH
O8/G/r5/TNY/+dpvPwKMs4Zn6z9nbkeH1VOiUKP368esH/AlR9TYlR5sK32DcQwF
Me8vOCSfnwDvS2m/ShMMjCiHmWhdBF5EdoHVpCwXPu25Q762oKn2SN7jgI4QMGSL
o5gQgPm7z2s+yPh6by8x32MKNrY9svOk6l3j6Eu4k3QsTOYYDDPQzf7g5IZb40Cz
n3e6VzI/EACN8AzGWBX6brSFVVh1+UpyMuQ+nCViDIsFzrm5bZzdSnTA6r6MW42G
wggNHPDRJuFjgsro3DkCFuPrO4Q+FXTo1ArEA6712A51QbULAsloX1sl742k8tEv
3be0p01bEpFoTr/bYJwUEe/f6OsNvzothF92uLXulKijmCGOn5IllcF/JwmMnUVf
LsnfqX8yR5sHWAQ6bh0Gj8VaNA+46HpAJrv2KjQdMj06SO+S+PzGIKF4RQ/av8Wn
ThybZIUxL8TMmMARBnpeJcKAofFrU/L5n0bh5YsbRgoPnEZP0S2oV8L5kKDCeUup
RbNshaJa6+myy+IOcXwFZ42Ue5B+/IHxk+fJhM+YZ7NSyJgVzopxyDDRUFYq5Fe2
Tcy9CtBHAtsL0l2FNLcapnjtiqk5qUOZQevZWuMmxycsMbvFMA1mLlEWEklCyGgF
LudLMPuV6eAN+avVPxutwPYTbs7I2yMOPQSA7qFI6v0Xo7xJqDQWMuHIa9GDNFwL
onD5xaFScETFczu7fL9wa541aLgYkwZgUbuxvJYTmlTFYnCilG3tHexr0KxwQUSQ
9a1IjnOiwmFx9o6gMOBDnao3b9e4dblxVbo7c/qAzY7ZDPLXMJiEyziNeqTkiJ8b
iuql8OzkX8qiUfq94uqSQMBVBTo15jOKMIe0HmAnVZqdvy1ye3MUfByRqVMD2eAz
FlY5RCDYhTV8dA9yXjLFtr4MV4QFC80Gj91TBX83fNQTKH3IBtYz3r6TIFMah1Ex
V6zumrjpwM3zacJGLPrZdnLK+V+EJkMjSZP59SISnCmg4acSCLLJq5FXF+HPX4wL
daots11MARlc/nt1LgckDEFDS4RB9+9bOPuwxnKq5MNQf8ZmdAFVyBiyCz9mgnFg
EXJNBchdwViFsIp7Nhoc5zyuvYNedIUBjIecr2d67WDJy80KE+r2dMHUiIm1G8t4
xskKIW+gj7kgQTm7qAS6OGzRusH0xkpsK9lGL1gbZMxbr87V9Raggfied935DXvx
byJK0ASje+ZivSqaZbO+i11Zj1Pij4xi5zkH1924uYlgFYDaeyqJF5fG807B/PEN
TohKFMSqgJ7mJ4fGHGrRb1izJMFYIfVolXNJK2FfMrctcWQG99l0M+5VAs2Uh8LV
DtgyDiPMUNyx+1ZDk7i2u6YNWvfrtXUydFdfox1kvxFv2WZFLnXxCjfOpRVqBTwB
PmTMR2CtLbVsVWYRAtR9nQkG9elGMSp6p127bHFrZjgZJ5xsdm8gKJz1uKvsYNSU
FHiHLHdF0PX9v/UBnv5SXhaK8ro7wN7VM31otdXG0SCIj2/tbJOA4fDp3PdTvcrQ
10UX9MiVPdN+lv5Gi9DOxVxE7WqnUamH96laFYMNZEZzz3QCYphmkqzZVMhasnR7
4tM0bagHktZpkm/Ho9YRe8PKaU/GQXjaUNXnlXpYWs/+37EvEvcuDBRp9sVkqMKt
UWccmGPohorGRs38y2zuabf/+EW3ituNV2L98x6XTYHK8sSOzLBnEa3bvO4+dbPz
9w+T8QVLMFXEzWnOyZCO7Hir7DtN37bT9+uTOA+rkdZMimtWK6Yl7wKEQWrqOBjZ
zhLMD9yFM+oWDTHVUxUF0FB2ETxqf7Mbo+iEXXlI0OBVtTAu2BP6kUBQM12Oz+CJ
ckjg96zzIpiTMXwQin+p2CLjhZ8RaUFn9Jmkp66boeIbqXALECzkPk9Iss/5Jkd8
AgeSYe1pr41Az3VjOEWqbeu9TrL6uyz5pc/QEUzN5B/WwGnQJa5+OMyfqGKhc7k3
/IBKxpvFqEOXOxDll2K3QmGit4/t1deviWcxR+43yFzAOEtctH1tmt+E7m9xN3xy
pMn68BIPbQ27VwQyXPZhBq1s6SjARuwOoJR/TX+ppgEODdhPSKHdEDHc91PXJsHZ
6VNc5cSiKr27iAYIKOISR+rP2WVqw4AxHbsQiJ4/W7Rzh77glF5Ug81+4HreQu6m
bgMB+oLCZcFhL2EXgHpS8z8E9QeenndprA2Lu4bajLwb988vIIF/Fvtf0X7hLBc8
N73cFO4s4WeQuDryQcJ9SzLSVb7VZptEnHabXKTI0k2KOU4bHfoPbKbUBc+s+fgR
u+Ukbf0NIXpDnjCP0Tk+jkta/7FUCxhjvZowXE6ju3nXgzpo14do3yy9t0sJsxHM
9ukeuouXM8BgJOXUD1UmTPkWBmVqvRqEAQaazJT4FOcd+vxw7PR4H5D74PTmX+hX
1MOGqUNxsB546H+i3p8b5UCcogp92K5fajeJS0UGzEg1szqA60tTX0+e+6bNRE25
BtCzVyklinipr7SOhj/d1foJ6uzHfJL25h76LTqOWtYYV63enkD/zKNA9++5HrYO
ScyjNG7gTUqN6r9W2jfximb+YJqgPKUcY4lqvbg8UH+eyCoUcipa/9KQNvUNqxdh
72FIcNuMpMAygULNJYIx6jY+t+1sKB0BYhqTbNmOgUmsVZXQWef1lFlum8uO1Uix
Dt3fuQiaJ1vTevWI9PLiHpE2MSQDkqf7LI9ul1qFvPQsHXiOjCegPC9sAeJku4iV
p80LVvkF2sJ4JuhFwMD/GEOhp9XmQWnZWCdiaQg46Lddf6oDIKseBXSqAk8WsoLf
CcolV6JBpAqPODEHYCVz/X506DbE+p7ITYnxAIN5US0yIhkDDc7Rmyv8u2wiK64b
nSU7jDQW2OgE4KMYFbqgLWz26T29ZoQ1ddP8sY06+Lpe9qswZBccq2GpISf5NSQP
6sNq9hvCycfq8qwlnFasAhTDthlLteLeRi5w2yYvkwM1kYZww8JPeGRjvSbpeghZ
zgYihSwTRPi9Z2MDpLcF/U3cnS5t1sjd75PKm6Dq1MyWyoZdMWtpphuhDMa2PM7c
cnBsIrSQj4DzSeKKGLAl4lwqZFwkhNWuQ9RmF1q0hMIV31nyUeEHywmWketTG10M
gQOw0yxkF9DiX6if6asfvlBdRZ6Q7EHVb1CHuu+kPHVd5wuoQkpj9uUXfgWXsLN2
aXepqyHAkRPrL9mWplYbp4v4Ehi8c2rwTawHWnACLuGImRDbkRVYgz0Ucf5rb17L
wkVW3wkVJDIU9ieHR4U96XC+xZ9+Cv7tTuzv7lD/twceXAIW5TRvvgB7dv45+AqS
FiQxlM4rkbLZKj+C1bMLC+cIFTaxJ+e9Zam+lHA6zVcFGWVthqcECtzgHeuoF5zN
cXdr+gnCk1cLNejEOn8pkg+qs15T8KSDJ2k98A4OlcmZIjMcrZtH+h7sO/KNLk4D
duelzU7n/rZWHvUwcZSjDYYYRippygoRk80gltt2/xGRCdrgw24kLWSEu7bZ5jMk
ioo72nVR0g+H5HI3XYi61jCBegIqF63i2mN5I+LbB2MBPuutfACx3/6f9fh584GM
uJm2rCwheeXxzOwXcM17ZmztMssc9dMdB/lK7ezi4j4BSzrogmI2MsZq0Qj4wa1K
W3/KyphrlnH8iS2ciGA8FizZzRuvBBMiU5ExYc/SlepXajkDV4nWQf0IJEfCMWsQ
zzl/azX3hKD/IbL1drLEo7idyk9Q8J/Il4tL2xqM0FUYM7e/7QZKEBA64KHGDRSN
uF9vx1J8PBUFfIgX0Kku7qoVCiSdY24JFrwhIdAc1ttmcEIetvydNa53rrAzkz7V
ZlWg5RnsjfBS6y3HvEpYEa1+3q3tydvboXcBRyOVNI2XsRIbYVkrsYNsZkxEIhcx
Y3JRD4BrOAnld3BVukuOfPLkbC9tr8k0zGZzvpc7H1KKEib6VhRPruwrxdAWgfFe
9cmkJpGDgIGHgnTotyIRycZuCPJgQfARMpSHuOy3W7gWvzd/KF31nwRR1sF4KLIX
2jKhnE54eKmkaZocm9LRHGIvYSEOKfseVPMQJgyYxE4NP1pSoubEdCcT7deNVRY3
gzSB4MfUkn+BnK8qSHJFDEbo2IlK7qUKobVm6ZtThMxZIblGWxOA/j4l2eyGa2P9
zwiGZo6nme7wcrNwDkvh147MW/ajNekspeQuCMOfx8HdJ+4RQ0qfTl8wxWZuKtR6
DKGrY37IC3bv6RtAcafiUoG7kgmU+6QzYEDq4K47FJSs1BhRIDmuDgpzfQ7u1K7v
5yyOSpt3+9oycw3jxHuR041G0OtNGubeZJ5ehBM7VBMoqXvpPyvD7xgjjt9BC2YQ
Q9B9t87aZPq+njGTclB/lugjGNbzAHsqrpcJ60w3tXCi9HOr5oFd7bH2lXFxcJ06
50DaKMeF8JCljHn7bxVvWHIAAq1j7bMDK0cjMMjC1kvFTnwsJGGCO4y3l0a/gOLW
Jo27iXYVg0US5l7G3pO5s/v3VTbIP1aqOs5GjHbQt5Pot61s05rVKzlICBCWbztr
I2cnvQ0ao7d7Mu+IsaqCcoFvEnFrcIpT7kZbQaPe2A01nhiKDRNsXfEtMVPMHwOn
Lgy7FpE/As0NbP6zANdECjzYXWIm64ZCWDkO375QoqccAPkfKoT03YA3FZrYeSqm
+v4zmz+PTgxiDBJpn8XR0ySZTqgvdwU9jiHHbxCCj9nW4b+bnOk4IwMGZiI1/Vzu
0Ua5LxTxKJgf01zGdjfmji7aZe1yvk26nRn1opLQ/LUno5202EIeBgKbQrCIVss0
v2kDkoi1u4j9bYo6KRqgudsyrfdgKCZ8QABQLXUw6cdoCy7fbkkL0frv4qP218hC
tWZRkTZMTVQIrOXNjtkmtGXnwSzxlrrRQUbCkbcSQUYtckkbjZHOFcKEvrz9t+wE
1Hkk13/FkEfIHsfxO04a2HIHPD5Zfy4X5VtGacJYmMDhM6w6H0I7DAbU/sV1XD0w
eK9czaKtTZuCZuWHKJFW1CpDgMrwhSlX1lr395R0mDrzSRnaSl5/GmDJZx/vqEKN
Xr6pYVGgWi86NG07nCLaaGS2fNAyDsvjSrKihXaVoikmUHp1Oq4frCK9OLYBGGQN
PE6VDV2+mmBEZb4HZlI5el+c72+6M48FLHb3IoUdQD/HTUPYrDRje8qTHsVRgK+n
ewgz9fD799LAm5Hk1jOEjyNykXWErvLtQzDbnJ0gG+yx85CvY4oAAjd524QZJyNM
dsbaTucfNTHEuD5YPJl8Gz7aaQ+Hvm8zv48V47yMECkhqL4ZbOGu9VtLMH55rGEf
oaBU4ybe+bE+sK167f5CdgnCxgBygEXWL/kZMMp2ccXluTgdcw+GZEyKKb+/V0Vx
70yK9Ffa3GmxUzciqL1ZTgasuBm+kY7J/ZNdinJswtX0IUcClcTMHUuDYEBwzPec
2ix/ANlHxvLUYzDCQBsE0huYuIMbtsOAptO0qID9PJ/LxLekvCyr93SR7lInwfqQ
BR/+Obwg8AvMd2tWiqaUJeqvYUlz1V2Z32bKhRcpCw7Y2PiG5T2yGQDdm65eZ1rk
Jz2uxfxTSTL45InX9/i97Iqof6J5B8Hwyq8nPLpftZKtvYw/ywx2VFaFX6Xschco
ZSQD9x/vRHlP31QvFEGsBTgNFq9zyKoB1SiOKBPpGHwLpWOWkMoYENO0cDnhnRF4
VlV/qFGgud2PIlNF34qNzfxLWAHrhXkHGQq+JjpCH2HjsHMGVk3F75Yw2PkdIC0I
Z5VqKq9OM8agX49PVsMbKgCCzttBV5uPLEpzj+x5fUjF7L0DT2yMGtnVMQA6G2hY
QljRWkMhUEJ9Z2yx4MwhqX3F0g5imzLTQc8U54oCvRrBzaOcmV5rk0rufsjI6Fj/
6csfFXebyn+Z3gz5sje7xHfx/L/3Py+rlZi0NzeByJRwSIOaHo2Mu1Lrb+AjVPZM
38gdiMKXhMy7SlRnqc6ecZQwIz6tca3nS7ryumQNOl7YCYU33curVfi0xgST9vZu
ttuVrjLESjSvdZcN+Yhs6oGluAmNly7UaE8o02Ib6sSrXIMFvuZzumDdx2t3uVi3
BYFRXXlAhzPTJV1VZ0+oZL9jqV9Szy6FV4wTi3xV6IixSUOdm0GcjI1SWWSgAff7
g+UrGyWMzjp6+9rAQi4CEP8Gc0N8SpXyseueY2veo9WEaOUgzMq57s0Kf4Syb0Sm
Kn7Denap4OQtvLQbobOmLPVFeEsmOQmX8W/tTwuY2S61OvfuL1RNo7QvB4LppP+m
AEkUMYKS3X0FIxNzWoab/nZJ28Xn5/cdDSQSvumhdbFQ9YQ4BBlS7Uw2oU0mReDI
nQyRM1yxGK7hyKesnVyYx9pkTDQIJXV9mVGBe+aL8s/SFRSxROb90uNI00ufBSQM
ioVd7QG/NfSEenpM8FK54RONHC+Ae7JHGRoe+sA44hcueQ/uELfX8AiV1Y00AYPs
2nXj+ciLYK92uRnX4EpBn2yLAZ02Bh5I3UciDv5Vt6O3WwhH0hBWLwjXO3DOMhKS
59IRzsixQaTb7J6oYRt020y78KTqJHZQbZDkbGyZbLYJtur0BFYUiTrNC6DInh69
fG6nB/o5/U4tqaErUFodGcpCpeEBe89yMItl8uLnZ29+7NknssyNnCav6CCPvIAM
fAbs2hD80nVAIqkaSg8MoQrtaG1cmll0zcQUQ6PmgJsngoWwB/Hqf67b5z1JRejv
JSl5CmxzMwmKHhRpv9WquebWt4Br8l2+mV2BLWSWQA0U3cgHh49VyRSK+M6YC+Gh
IUvGZC3pJxE+hb7lsDxLeLvK8VA5BHRfGYg2JSsmruTeGHf4G7lPbu/xU09IldIB
kut5MfvFI/9e8T6yWXH0sAPHJw5OqGhv+3mB+l8dt4LfyMcUpJIPzfCVzedKyDpk
a4dQiHPLiQWjPWAYq8TXZ9/w+PW4+wdStLKdNHohPcMMuy8K9ih0Zj/SPwfvJn9I
H229xJ6ym1RVTTxBQuvgBeWB0iowfxAXiHtVyGobDLsxDTRlJA7wsM8Bgu1dABnt
SBQI8eLne4KW3ZjdndZ88f1AA90ZrhtTmp3GgxyPIKr7gIvIWaCxdysTg3ic6vqY
qzuhYKX04eILdMqYr3kw9Pdw/QPbJnebovXAgsHucQZ2Vm2ZwXNtNeJhm3SdK/w4
y+jJ0PBcr7uuk9aGV3l3ee4NyzG1p4YsXjGDNL5d/4+H9VvEbVDLESUYw0pz7unN
ekBviN9tkQWz80ntn8NRFYF5jFL0vWH0MFD77h2h5WzfhEkmWIQNos43EC3ZQuNR
GCUvkh/Jv5TjvNqa3fq1jjCUVDdhcLJNxdGAVXLSkL3/aXmm57sVG/zuL6D+UOpE
8fmw1ETRxqoz2CyqdaYd+6zL8s7O4TSqVlLzipOfkErIsv+RqLpY870StSbDRsaX
9K9Q5Rav+BwW/CJNyROwBgvEZ4QxLOerSQqDd9sT/QYEw56E6Iyw/co3Fo+e6XRz
i43EfofwozKDloKHK7Ub3wkSxHJqx12rc1VbIaPnITdTqV9Vaxl6JSvdLR28/MGG
sDZGqFMfJ635RBhRTURywV46cYM6Utu2LWCnLVDVgLYU5O9vyAJ2l+mOIsWkglRR
8CHJ2icNqukdu5kPHRtqWwM17IxdiGYRn53CCd3Z4OI3X8ytjsQZ1Uq/N8kKy+U0
UV2H/LSnsxMrv5XmPcKNJTaJhgB25dMUD3oIH7ge+jP6qQVTPyZGiXLmt46CaMc/
EmADqpEhujHq87FztL1WETrrc5nD0Qs3cl7I62ypDd+VpNbUT7bYN9dzuByVYIl2
U9LUA214mgI3R9MGi0TOlHosSsXtbLlrqNPHzRI2iq6YdmNFisRGGIEm/ZiabsnX
/xgyTxTa/kRzE13aZQkAK4XzUvskG08B7sjo+82RlkihfZiFSx4yJeBkkFA/OzAY
4dz/SpVUs0ttBwTqI0cja3atuH6pHYf9jpaiI0OgOSK6CfL9qhyCxJy2yxFjLY5Q
mQ5kg6pZOe94fnoh0rybHfXPSMar+TNAHCFZL8E/xjy9FxPiXwvcumjRIcFL4YLF
2DwhEGj9j3/OrEq75WDn9U5Up2PNF7fI5loVJoAobPDtpcTep0AIJYgHrAErERI0
Y2LPUjnzqSYZjI1byg99IOFefek2HXDV1RbDTxSs7LpRYw7nxVDxgc5QGVegnu1x
DLl+H61s8nA+MG2HeERyXfTnC2EBuWEzfecx6JR4hHAGo0PYR7sO88TDuOiUKIdr
8vI9vmLu2uVmuwL1haUDE+ALsafz5qoeutzF06Ie/K9U3MienNjAd6TxGLGl4CXd
X2bpSMmgo6oox/QfEVZIdW1zsL/LPXQoz3YJB1+DDozTG03LHEhxo9pb4F8XyrXI
ghACmhPvK0feh7YCl81f+dTHhx/IaQHxlb9TvIIBN0IiWSP29r82GvPgsPhvy0Mu
O2kkbCAUyL1EAw4SFRJ3LoibCW47PRyaJVhPZWjj66HTRJo+7Ag/z79MqVcT0zwx
hO9CBkH31+Iuog1Y1X2DPqkWx10gneGkGeIe+nLPtPRmWTn7d9kD7tLq5kCromqE
4V6tW4Db2IVaxV+W3VloKQGxsI1dm7ZQr1BZHgmMbOzeVpAdDp4TaFn8Nh9QPHVK
kqNVfuUMclJ+7xJvJFZhY8KyHU1OwQzl0b6mR0yZMNNXa0Ou8lEVLZgUNLRbh0xh
WSxqPRqrzHm2kyOvTAWQ3j3Q9GwUgw43vyLtv9aPb4Qb0N/s7WZLs22lRv9IZ6SL
yfm210fn4ZF0xyt2H5vJNbL//5L7JUjsz3BAdmxZ7B33OZZuwbyiW1mfZsKzvocc
3raUL4JWvHPvzAKFcnUorpm0E9o03IDM7sec+w5lJoscb4ds3w91Aa295v8rJS6K
WuwGFpezaMTb6EZRt5IcAYDFJaG4umpcXTCWfePhkdb0VzGThGrjt6EDoO+On5Q7
rfmTeE/Tzo+nT5PqsYhVncO2OaepFFF6wDmMi5q5nML8WTHYjO3qMEy7K+bwsBWN
LjVK/kAMs/TSSnSgRajFlSWPUBdNSeAYysp80iqezGf6yMnEttFrPohsHXWnBqZf
fY1t4i6pDP00DcAVHyiFfUtrX+avBv63HajroQADeaQSN/ubbiOeCUZ9LAvy0kzD
jXme3inZznjARvq8iyUjCBI1hxNzy4OzblnGoFrpMr4uMvYRIOa5rWz3ahr0wdfO
0zIkL/VvbULrhZfx/yfEygQx3vtQCPqkOtJulRARZuDowF1aTIZAt4TNVJMXumFa
++rHZ/Fywqa2hilW54FWFtnvcA4xphll4FOaAJELFSQvU9VdSyPDz8ZWDVYisYy+
NQohT0xrBtVBSM6j/RriJVpIn+nPqOI8Im2TYrYTCTPdJE+xnHPOJYckH/KTx62I
u7lFrajDtKDnF3Py8IMRq3ehGVDV/Q2otxuylR/gHUe4K9XGivKwFITNraCBHCwH
HLbAEpFXGPj0QtMgrwirdk3IGrBGEX2Is5oDn7SkI94UYCfLaJybu5jqbIMXqqU4
3VM8PnnZi7FLVHbjWxZ6lqvFtKB2uqEDRe/bHQZmFFXWjJwEX4RbgZvwARFt5fjc
/5sNQRBg5+VYPNqve9K1Ygf3RisV2fgnr7Pw8SzEI2xprs8TkdaYx5P4tBWT3jOP
AK41wss9cC8L/U7S10GeZVgL+ubYDHk0vKsDjY5FILTEwjsIfRsPs5PsZ7yUf7+1
bNHqjQVxwt+/K6BtVI0HdwJkBG5KM/WgUnESx7mwL2jMaHuXpYjLl7q2tASPZAyS
qF96TJuWdv+44CAwiIkMotB4+pbzNHW0dWc342s2jkuFTiV7VtzbmfKdaVQBW81o
cUhDS4Wazz2x/E2iyV3EPMRzKo8kClYVeHtddY6xpGMe24ctbziIQ2+9Clsxsx/Q
/bTW8/Nmuo707DeIQTy3ncT9lKTh/FouBhmZpM/52/MEwo1CDPx4gBBXCAYE8LbS
cabmcDahvxI+TjXF5VqwcHNfFAZvFR2qCTS/70GM+mjmu+mDfcwm9Mmsd12N3R1r
qDuPjSiQDzyCgqe5kxMWv8UNlVgoY4Ofwy9Cpc0ritzMoRDLVs8DpgpubbIld0uR
l4IV2ZeiMccvbRCB7SC4JGzt0vxc6jEbc3mJfFge7GngAfQBLPUZbpVfL0o0vTjZ
rodgZzQ43p8o8l6DDkPcQmUko/tFZeRpq65UI0WjW61/ePiz7UMKWdPwtj57GUk2
QqLfDoMTRQU4DCSE7tvJh/XwRYG6lNo1OfmK9P3T15+bvGFts5c/9CkTpqt9t8cQ
2JrkHEPaRQIkc2bpm06QL6TVST8pzKVrD5tFZKntZW5PmIuEpIAFRmwS6aj5pBFm
g3SsmFy8oUQFFoihvO5s6FmpzEdkrfRWQ+dIyzor+GyGJT9vtCmZKOcvQFDc3+mp
sMP52lxvz2uniBnkJ/bPUXCjibryKngxt32Bap2voUY1W/0BjGymgSLnf8QWJcKT
G90pse4JAl/QR66Lbi9nepINe9n0+gU6VzkwKhMryuvMeKrKOJeWvs6sm8fpakS/
JPIPnGhTB30AsVJ+i0cedqQtLEkK4W1wofB8YyYHSRIj9zgzrjhRFC4BcJidHrvN
IXkWXoHV3O4uj4v8IDMsUU0zGeyvrnVchDIBD74CZ5Qd8iEWCGrY1rxtGuFYL/Kq
qCrln6aWejgHS3pFr4oC/xluYSgB19zFEIRf3fUu6XKlICd2RvPZ1iBayxIOJHOE
HOJukOmrYtb0cKbSveOpobrA7Lxous2wEdYnMtJH6/WKYWFpz0TTrzSUTeotA/7L
k46+t5Dmnb3nFZKnVYgdGUrZzI4P17K2OVPdYm1mq2Q+qLU/NA6kUT2BnebJ0EaZ
jFnUH7kIzlr/OaxOXGF3A/4cY9B8YLCGMqEBVIBhEA+x4682/RmZ9hbcRdSZpjAg
gpNPSD1aQrOxcOj5Nn2ZBmcEi03zr/oHUJUlJte5VLS+CZCueq8L2wL8bmgqr4AU
HZu1MdKsSZQpe4ONzCYgz2xFGNF/NvqQwOUYnKlHQzSoBaNajd5Jogl7RTRbK3Jl
Vtq2bYZXsfVWujOz0IsQHL4P1nyKS5ah5py89Pm9DJbQ7EJlyWx/3hBslpW25ig3
wha/Mf4QSdgMoXGpIgpIX5ZzJCwRbvx0G2tgzU+oe9it8KV36H0Kvfx90BFrJG+A
TW3Sx1W/G7EGpMferSWFIMBYgvdcBrdlL+ICOYQJCHJWVBO9ESx12XbRKoAvhqXb
DbJGo7mPe+pm5Z7MENpEVbybd+wnIYpRNHOTA23+4sHNUY0EAFOdeH4IPEtnHS0b
ysKrO+ZvVwm8WbR+X8LzGpW5ExPzNLmuC3tNtW2OJmEEOZ/+ZlpCh5WXkuvsHxgM
RL5WTcu1Rqfm/rIKDTzIIMM82Kd4QIZMEaPzBJldcz697rZ0Ub6WBWB9aNtaAIhS
wB2gwe5bNXyd4nSNas2LHOZjTLCOE52B743FNwmmKqVZOJ29Vx5lhgQs104PDsra
XgZkFpsVQZXKQhEA+QuX8hcQT99RonGffARxpFrIK9SdEvBzUG9qeFBkh6kPRtC0
UvOuVMECOB84ijYAeHPTFx/YYRiQTmbKcNf9w+19METjPxzTJivELA0+KxolnA+n
Co9H5WU1LJNKXHpXzLrWy73Omdu1kRh+4M1qCSzLfxZn6+i1l/ku0yaNZYFXGawj
YhgKA1kAfxkNupSjwTyuAgeWHZX7J4uJru9iBejS6DaBjOsLAVtrA/ecxGe0r1ZV
geGKx5iEQ160DrWb/xGBmgRsVe1Uk1VpCgF278geWJo0NtFG6aePaVksvSYP72Ou
OJcKpoTOOC1sWmkLNnXx4C4z1JqjQvumfw0aOhSd8RZDrIE2NIjlD20zNzp94Vtr
nuGZZpdwytwio7/ibOt2XayzLFGnQZg2PBommZIkYhfWwfcXjanJznNXJEcynwN/
9DklujplUMkxz8YP/uX+ZQsDJAMFNrfJRTv9D3dbWEu4Kt3/4YCepANiIIekuOvO
5qzMGcCOHv5sUbZRBmeaOypI20ZRvjNuqgdrltkc1lKHKWd/RtluuYytBNjp2iPJ
WTlWeQd62nRAm67PA4xLfCTJIXc5k+7LE6OqQpGOYFAwN0BmnKHC8nOdEmqZdqKO
d4JXuhM2QDMQPADz6ifUpQhWfMIxPSJjXZ1CPVZGUpbZRf1biRMsIAQX2y/4dSnD
420hiWyerVIPbRrY5lZsqf5WzpUxz+xkbxdsiBhKUg5qa2hpxZhZJuw8+bYQgE8R
46tKv7T6mRIJZ927717RE7v9bRSu7IyPNjDAB/j4c3sIrJXH0IVFsWqBeUmdaFzR
GdzQcPMVm5ji+Utg98OWzuWzorcVvwlndo3ZWSPIvdacxvUD+RhwPYrspTNOMxk0
aezkFvUlcagsR/2uK9EhzM0tdkV+yv9CAbckKZy8yS/4QDWqfFD+nWAXr+ll4Euf
9I5JYIMjuY7mSK9ZThD2G4eboJS8w3zLMl+rYnNOoJe8ZWoe+1akNiLBZdVew1wz
k42Yd4Jq2r+J2GGZ72yNTIkYWoisB3X25PM8TGxrQGnt5WNaQqGaoXbbs0orZ6R8
i2EW9PKeuTeH3x/NBf2Xf5CgI3Ihh/8j03DIa9oypPCTZNaG0YRTu1P+TkhmG1M2
YmSlaJH2QBqMQxUNPsHdM4uzjLfIFotTLFp8wa5XMitQCSYP89qn3RgdPiyfzSLj
YCUWyRqYqOyrqsrrvWdxe6iFtKIy1FasfBlnaJ1LZyCZGUAIyuE3V/JZRc4Xsxk7
ZZnNn1F2m6pIuvq1dfOYPmr/3PGIHiKJKwFHQ/x4xedp2ZMhD5SjnjKHGxgbO9Vz
O4YdY4P4Rqgl9iZtVO5n5HdO1n20taTDSAbXfaJM7KWGPiCqhZgOv4jnmYTo8TGc
TAsHIca+ZNGeHtBPDPxgF7JtBdMogqM4GQbCmfu7qviTgsf13kF8F9kyLJYRhv5e
6zFpLc+Es87LdlsqPQIh9aCqLgGwIpCDn69+FchcelcoGpljXRurAL9gO1RO5Nl4
u+XWFccdBuj9m+drHrCTFzJpu1zzH9wkLWBa0rKghojAu1Fj7f3RWF15cDnBZIP9
4fpjn7YcY633c9f2zx2o1tl+3Moh9oMWlNQZVh43dV4VfizYmiM5EHP3uu8OBEJ9
obxFuk1+fRfonpDOvnAyeV3K29d9oiWbutO8D5j7R7c7beI9uoOwkzHEdH5kws//
tYStskpFbjrRo12FUmsSUnUx3g0Ep0i9N4Ci+44FtZSh2v2eHwwPwsYIGZD+8XIN
QZzxxZa5b9InVu0ebmMgapPV92KZee033yP1Yrhh93OcLXD4swjwJHNPk3EEf1aS
8teqVYvjO5ZKS3Jif/i+IT996l7v51+qWpEYvw1yGe8lLEEqFb93Mjqdume/r4NV
tusC2TUg6CYUlv3n1HFZb9GKffvtBJT2FupNjCkwZMes3iXwxYQUFm+ljwuieTpt
/kVLD8iH0TP6D0eckpQADzlaWXj0WTf5rSXTq+4RU09+WACqumsWTf23Ax193wFQ
NbYw92s35cXlUnRomCJLR2PKVIwZa+v41bo09eA91JcYnrRVzs7Vg5CO63EHV8mO
uY3S3lnbJxhWqCBXnwON1z7cQ9YRrad0rsI0ziDH1DXF3Fpfd2+rwWXwRhEpRL+d
Ts4v3OWMiBHUkHLW0budRbW10aLDvWroduQbqv9jAw16uhEpawiCiD7liBqaCsmD
vpK2iKBY1J6LduGSTTVitjcilYA7tSURIPvr+n4a87MJpqdYnD9AOH/VGzkkVRpJ
lhOAgs7U3Z0I3wLKAPaBu+97FFJFkwzq64RA1XrNPYxg/5cSlmyaEI+sxXhU7fpq
eXIn+in69KhhgXigCmfLNF7g2uBHKvemSb+LMVMq5sEk2qFOcIyohdAJAjvsKmsw
vaYXEGPUl1nor+p1BY4tam37pOhWTy9taTsdsN5urxW/n18OopkPgO3Hexs8shVA
CO9QsgPQzlxRNgJqS2V/rTV5UwfnCNm/AyCGMFCnIDgJM8OeDveqsdw9ofBjkBBz
+kFdVPq2ym7rxYO3ML5oBLh3riK97A4U1Jdv9uw3LSToZhET/7wSQhbSVx+B5j98
9pFn1rLrcr8AezFgxC5+30wpLxBy77HhrvgyrvJvPeZ50LmbooZ/KQdgeWWJZRku
z/0uH4sCMhcrGZv9kEcOliKLmxgcimKAvIJwedecaPFs7Zjfw1RGAWr4eNfAHPqx
sw5KKLY1WUe3lNRXWtOdD0gxHqrHnmE/8khYCMNWIWmVC30TFpSPkfLJ6sM3GthM
TruaKFrckdcDGhykRHdKy/95NUPhXlZApBwxXcZJoD3PKLSCDxzvzifmqpfYBs5g
PudAwC5trBojk6gDGLjGVCoIT3V95Ar5T3RgcLgi5IkS0FDYZfYXxNJmeB3Qve3M
/VQn6ZMp5RRXV5dS7ibAvrzevemuvoa7lvjNnyHPAfoYiqGbQJF/uhtb+amK5eut
4Oqaovflb16jw7YAAuThKLeVUm5y8ry0V+uq1Gb004w9CbJ/4//1u+dOxPQJ85aE
E3jtcX9mcbrzV5yi2Lb25+0cgk0Cy9cq6dQ1+cHRGXM//3qJcWrhviJlxtjqDx6m
aRWR8MDlXxcZBB+Im8FwQYXAlCl2HkrnESD1w9pGjl3OjwVNFoHaCE8hTowH25DY
ChwonE0sfAj8yM60w71PQnhnkhQ7GKwaxbV1FtT0ZjzhyYTL+IZThl+e8u+7Nmnt
g1LHSAQDD3Jic3TFhDcD/8dQKBDLhsVmb5YZ0saR3VHBh4X22d6cFP++WUq4CDgA
zuqwxoE7S3L+2L1cZXFO/6CdEo+fhXgVzdnUtegBwPHVJc/SF/aBqxx99ayNTp+k
uQbcCMp0Svrors8eVrDIx+5A3mA4NQ63cwqRPU0dfZZjke+FHTwWWpG2RReNwWdp
kLtXfpurPDUnd6GtG38VkA74QFcbSuQokao8kDe+/EL7iusBUZx3YpHbQVUuulIn
J+ZOODula/4j9VDYdXKK+xXOe4USiTyk1VsnSEYKYpcFTE9tJzx5swDdHPfesYSX
2gJDxoVbtXkHgXmcqek4g8sCQR3PU/H0Dkmr28aj63hmZDojWEvV3et7xrvjxZ8m
XldzN9u+XxgEAUN4c/ALu3HCjFoLq32m3gy0fJx0XRCb1w036yBgEkCM+Ps272/Y
nJC39y9dLkFEDSE6s8obefVD962mNhpq1xEtsmKbRLd8zT6Sy+z100A2oj4hdS0b
CaLymMQ6zgePukXo7wg4q7V78hoBYcJxhURUcu+WgvEQkUFDhTzfcIhX9Plp+P3C
NeBTB1akrsr8G8ku5bFyMjRvOBCXM5GGclv1ghnnj8DSxXSLleVQX4O6IlOK/v1Y
zX/TLzsCRRFJCwOVC/HOblm/6pSCZbazFf+DOAoV2+6uxMnnNizu/JuVqJwp+3V5
8urgV8VpY6q/i2GMto1CMrFHLjceaPhtfl3jk04F0zD9rVHNfOLkUmn7MuBSjK5M
Q40Y7kSmzu2wd4jiONRU1N2isa4KYpffGRzWF7ZLXkjsWCYhx5t9m0StQQhCh5UA
zgsdppJJyANCdhabVOjf7ST64A/E3KyZpNZgFWGtHG3u5+FNMYFGmZzHsooWgIMK
B3P3JmJDkgHpv9e9T3vKoQv1xHb7ndvbXPqBjl7AU351Jo0ihK+dTvGFUitBSPKC
CSjbBLVEvC7xiWwI/2zpwPGrxS2EZmqOhnyIgMdhS8u8aFyI6GF4N89p6AhHILpy
EeA52jfWMM5V6GekHkiFWF6YA4QuzBGnQTaoAfs/P7s3JWj54VH5oQHwEOmLaMoh
qCH87AvfsEg2igB3kpm24oRgb9jjEgFeo14pPufUE+ovljLXXSUXgBklvaT78j+e
fMeGXsV88gd1HTEZ6o94OVnSBvdxWz7MxHx5RprFZYHKj2HFMgufGYYblS/DJB6P
8juAodfSQKd+LLKVbCAWUBTjI2abDaJhF0GJhmWCzhbYzET2loekSK6dyOKYdC+S
qyW1HEDlxDQ0qFDq4FarB/+sa5MpbvgTkUDLk6yO54zz8SsrdXXpkggfsEzcMbSP
VZbfcCPsi0OvEnVKNhEMXU2kBigurFm07ERXHa8noF8AZGD+EWnNuIcfmYY6fTb1
1ZCLDVuPwSIf9r9pPBmhRxWQK8jw1mErzoXWW6BH7Ki4kSOJa4Apm4mzKA97HlQJ
YiPdOIIqzWaRJ3atnLrguCZ5ZL4KnI5vK6plmmwWtHOZrHW/S5tf0ogOo6tfazaW
U4Bbny/TLQjpiWVsCawiF3eMeK3Mvo5Xexa1GITWmXe7cvWKIYxsGjbGVjKFptV2
B164AfL5egDToXUaL2ZTOGw9NAyfMHaoTJaQH4TDcbPQqqFuQq0jePZG1hP4EqM8
N8xJZI8lpwjh1eAjf0+XBQO34ysiG+KtpC1GxdIAMPwwhg5LKHjn1h6dLyUY2lac
VicwAYyWrBFW6uYm3mEcG+GV+RiS+W/RGtSiPgz52fXXDIsohrstvPz6MfRcvIv0
rYVjPN7HOM2hChSK+evrV5ucNYtCw8fcp8O5/DGHZ1WrJdHDHt4PO+OIAMn0M+6B
Nx0fVbrhub7MIN/mxo3LaYf96lApYf4I08M8RGDZ/7WHW4EBF3LcF6Lngbm6DEoq
Xl+q5TeHDOY7FvkhzNWa9NQE5fkDRvjE3WG6HmoA8u2Pw0jmfLa0JH5I4XGvB1fb
OLAH9P1LXQTyrb9ggLYKRu7hYqvzWuZFMlxbg/EZHU/4CHN+hHnywpRico5CS4Vk
sa2lXIXzi0CH65rluvCAogBF8ppK0V+oXRZ4T0BC4D6Evf7arqQEyHdWcmNbJIbe
eBGea5/YdHG1fej1UFX+pvhfYJUti7V0hbKWE0W28FYNvl5e95J2R2tG9TdOg10Y
6C5Xk2y+VKYav3ONhUsfjJpSL+4XcdNGrRbwYumSdtFlvjVIZjbK6xaQWWX4q05j
YhJbKuKoOvKUkcXekyg2t5PBM40W0ozSgDOQ/doVwoxa172+akcg7BCQb+Rv9eR2
wzjEOv2tQ0wzvAWqNmLpBRKIuQgUQv2e93u1CQMuJHSVDQ+38/816hZhVuMauZX2
nBUqesi2FhgiHe+anZNHDjUHR/D7HtKUsRZiLSM/0lskur2sGZOYdp3TwD5p679I
6Kj+DnyQawffpvwN3l6z0JXY8S2dpboo8h7TM27mLGY+GF79NMZfuq1yw6dO8TNu
d0MvK2I9zeuy/H0xd/GvOsox6jYcZsjGqI/IXM4iniof1hLU98ceZGXefVN83cCr
rix3AARQn+LXKoJsjeSs/aDyj73laHijM7K9kG6RRDLzdzdmVeTTmfGqOY1Y6UOk
z/8RKRWmV1edTMF95cMJdZoEIDSvTXVIW+CVAAiHn1u0lyieng66S5OWfUpot8ow
CThGv30aMFFBn2/MikKzJnPsiz+g00Tp98GSvTJP8fM22QO1jbT48Gbj0LW+MosR
e2jUypm6SKTteP/xTAHk4prjDMPLASkAyO2tozYy+wlx03vTkzacUKx0T/XkQIO5
r+h3e2RisKZEy2W2VRtwQ1uWkO430tLToV7MCTTzVsrOcm4vbpaUtWEPaEhapV5J
f5HAcq6G14760yf332w4agOwKcjhJzJAW/bCbnSMa86tw9bjynO0+ZyXVciaD1GP
/1TWKDQ0bjgbCqgodoJCUjBy2qy7laUiu7uFQqOOYrS53h+A1cFqE2GqIOeDctwz
/2e12krCSZpGwoj1g6ZGm2C5Z9lSc69Uxoo+SDkB7/G+JVeIkOdYJKSTrF92HAHm
/PcxFd271KCxispgBjr7KRyMU9UStSXV9S6ygr36D1gUmoPi28LlXQ192Lw22YNq
z442vieCy3Tg4kOYJ8V6cpisx56kC0F3ig0oarlYf1+Ljp2/1eOcMQnbasDsYdn4
h7LRKLhIorC2QVUMJQ4oOIH7RJbne13fWdpkpNPk9vdTbWazF+nVIsQAoA1Otcby
fJsMx4/q5KIsxaJ/98afiLO879pbnYRYZ/pFluozpMhEG2kRsWachjDzbaJ5tcy+
GTbaQUz2EopSwWd0ieoXY0yfSD82Qo68TMxteOmFTSiAXURGPLt3+Ys75p+C6m8K
zLy9hV760uFXTB+gxQQnl/cvYR+J70D1n28mdzq47A3nZfy6BwAAYoJFWCV7pwXv
3KYntfGfmxvaQrw+0FOyXTzcnRjhjLHFU3n9OKQi+u1reY7wJT3YjIxzQ0gRJI6o
DrnbJKeboXaRcpbdn01py1CriTyoGknVcuLK0Bml4Cp8DB555bDYOGLbZifswxGL
06sRPXzTO2uOjJReG8GWczr2B3bW8ech4LWuM6bRZBHGNTErCiHCfe74hN8X0Yme
rlq01dMNVr9mc8IWp16prTZDUUPgLAqUfTCf2arfjADGk24+6XOZ4qNd9f2DhOJT
3AyeR+iarNKgtAs82KdQ7Xdtz3atN6bnSSfqp+jN05d80Qc0cauUrf7uRFp+JK2B
IdeqSHWUN6UWdA3i5fRevMVlZo3IopOWBDmvXZ4wxXoe7KiV8p1gkxmi387X10Yh
ITrN4aeI7g+wwyfpKoRKzljXcCkBIhCjd4SE3AuiIk1pwlYdSPdc0KGNkIG5W7+p
AqrpLZM8lR30qDC1ogNWynKmMVHyWRRUAW/XQRmarEH3bek4VMvRIb+dYaw93bAm
PDmCbFwFA/KeBOfc/19WDPiUxyukQJguu37ZANUoawRSbiN6Y3WvbwkehSkmyZXe
dgrEG4gnqYQssFomhDfNhaNB99uK3d2vDhIHkNN0qpF+Xdv4rP9rl0VqahSbFgRa
SRtgHFV99nzrWYDaxSFOQH1HFVoWdjVIgA0cA6DfZ6VsRJ7jh/5vnWcuJAACYQ7q
SLHoeiaRh0eBV3It3Qic/zPrly7XiL3eDE2Oo1zad4WF+6sAQRRUBitB/SJNNP1O
hvZVmh2nssAFav49VUPjDF8ltS4t1vjH0GjO+rQOZQmlXNIaAXBRIUZNtqJWvBda
QjaRbtcTvs2wZUeyydvcgsLPh0oY9N3I1+80m28rwTOWOLHOH2KBl3W7GqRv7f0/
uUxQeFD962lzow1QI5aZlZMsmBVQweT3IkKPHrEOHTUQbhyV23qS3rjEoK/dmSeZ
SSboNWsgmPjYr/nIPOs0ZQ==
`protect END_PROTECTED
