`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SgcIcsGnAMff1Ln9qdg2cvRsHaeTujB7tQjTkhRVWVSIQpIX1e2Ea6x+Zc3rIp9r
q7xBImWhmEwgFWems+1BciXbqNI6varXSkXuwv+EvuT522IUSB50Uvr3XOQEGvUh
o4sAtbwLWwSOc7KnYrzd3Pj9k/JIeRZe1CkP1vdUIdm5CvRn68QzuNaNcbfQkDr7
k7EXICxnSMLNjCa+adlcfRz0kVK0DMchx6Pfz1lczu8E3Z97YHf8MFENk+GcWDQl
dexJAhX189V6dsdEdpMpKxo711GynWk6zMT5iYnb4rsfse0aI/MS+3h/pltI5Nmi
daTlySZ3unZxkcH8y0VdCgx9zr+yArjZoCTrDGRydSV/tfEl0i1Bmeu7XCk/Qu+g
2PMUeSvopKaHW5AoXoa2PzAM4oy363PhVpKsjhk/7AXvQclNrez4ltPPt3KTqeoY
RUz0U7RvI7ZDbzIJsNlO35IflddMNb4GrtNeopYPtsXzUlFIPNOCdtyRiPXz4IJo
`protect END_PROTECTED
