`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MojGUX4XlAJjVL2VQXF3jgs+8Z5gJjc+Lwdb90pxC/lY49ypXifGlwsTy481tjOj
yB71WTMMuoDORjJqr61VZeg0YE3oD6Nl9JcLtJYXrUengXlwWwESB78tYUYQIckT
HOVAcvTXlmF7eteUz+rIWYNZt1w5DLEzFihVLKppmOAZ31cbC8jacyvnf56A/vfu
NqwiJpqWPzYHQlYcEDsRreR/AKf3iJ+DQ18FKJDvQtpEK0RZzuPylwx7YAcHOeDs
HFlagZDNY8TtihbUWtqzcmQQC1s4SRedUS+HD3qlAt1f0cj8cPrZfRVxxnt6VbHv
cUoRJsFLyzEoCjbx7aFBif8N+6op5QXkle+4L9EMiWofwvCsMecbLSCwDI8zK4dN
AJAFmoIVZaTO2PMwssoJyX965c7Us+ZtOWf2fCeaiYU=
`protect END_PROTECTED
