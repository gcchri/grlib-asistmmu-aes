`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XK/+YZBqg77uQZu78yIt/l6dENsLSbh7K4pcUwNDTHVE5UBbkubRYSE7YPQXI8jr
w4GFoyBYLXnu9dFk5A6UWY7ghN5xDKiLTDOmK6fxD1Q2hoUkcd2GzH+PcZueUj3F
PnMJCXHb6XMJL/+gJvz1mLFSMXqXWrMQvkQlW4KP1vMWxZHnob6xD197Wm9/WCxH
AnwdYKdDtKMRSU3BnjAioJmlkaZBaDosniWZWqgtMtNifzgHKsLmxKgMNOr29gAz
SZuYJlXuAZ3ia/WYAeguIiEwBWuCFAFYGKz/u0NxgJ3ykbupXvs5M5wOnyZPcqa/
THbzfe+OrKoz1Nx11IHo3+EXzrDCJbBf1TmphzTmakpvvi5wwSaW4GczIsTBZUv2
6EHjJ2EkUpKK3vgLAivRWkk3/8qOzoKGfqPlqvx+Gj/fzhQ+MSi72i+fWYXf5FN6
X/4PjGuwTwJqMMxWRgD2kB0alC0Tn4oLtX3LmpW5wC4mcezazcSJerwO8+xCVqsj
eBuzL2NfjHQVS9jJJCopPxgFwXsOcGZ634HWrxYjATL0dJdlAELwHgb+Yrla1ypf
JI9pcHGPTPvN60o3qXct+C7Mw7xTBeD1vX3rP2MoTE4=
`protect END_PROTECTED
