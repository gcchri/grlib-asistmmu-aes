`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hFL7Y9X0JEXHkvxebhdK7oqj7nHrEM3iApyPh0dIU5rOjKE3PX4TDfjDKxU1HtUB
DnyzlRv8bQPsurPKTJ9wyn/KPTaOhxi6db5ms8nm/0X2sVD5Kv8i7eHKU05H7cN2
vevdu81cXxF0wZlaTMcl7ao5JTK+rBvtuYXaWIlr4cUBTL90Lv/RaHo4ltm1PC3v
OH8m4+00/l9AmeeCW2HZ5wp7QNfimit+cNJX0xBYX481mDoEnOQ5edNYj7OycgWh
f4bDymJoUrWXocNfZAyhpcRO+D57rCpVPslRCx1FVNl9zosMRm7POFWIe8a8cs1a
R0Gt4tu/xWkzFz7IV8XO0aS/mk/tBYdn/C+2svujV/AAxJ64BwjQjOBpfm7PbNr4
/N1QejQ488mIPOzP7f/KHbJHDdFCx7+QXN5jRvDp8ZeZukapvG3pUcjGmUGGOXtA
ag+U+FACH+/vbF/mX8PYLd2USug0Th5ct3gpv7wdsfHh2MfTk2AjmNIEP/tk8oxQ
`protect END_PROTECTED
