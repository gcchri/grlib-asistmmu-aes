`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hpKEAdk8rZvVp93pPE4TCoowKA7YPW4n+UsfrV1zDw6SJLKcoiv+eqADXpIUTpic
Qif14al5K1uOjgWnVAgW4ihQvaP7jJIA74HQvNwMmPKkkQHdQh7Me10Vfg/skWj5
uLmHhm1XSKZ0klmgfgcx3peaOGLSggdLMYfZWcJW2KfmCN7q19BzLeW8oPEa1BjG
pFcwoOLJQbH1BPDYV3U+b2lCeev66R3Oz9qKllVNRkQeR1+0kb6SOnRKQHcHYVpa
6RGK6GuKjHqp9PiPDduFUIxRL45yUwXveYmfcxXe6vDHWRy5CR5+WX5cHFhPQmiU
Y0tK9ETu6tt6wrgqyFuGgQpNncc/S0GWBlF5d7ZQYu+mLkL+mHYEd+MO5S3dTPUQ
zgR+ghIuX6441IGbGCsQn6h/+UMaDwbY0Obq3v57Qf/XFL4GwVU4bTJO+QQ+Ynts
LejMAs63vN5GQKR3nOxCbeUS3qxnrSdr6JOqt4PVlkcRLi4cNFHQGoopZX9T4Ogg
PgvNJcaYf5cIt+3t52Vaavm4wa2q38ocgzklcAvSHNOQ10pe/pDDmwbW9ps9C2Lg
jpxP7nmMCTi/vZkvJXHdpdRkUG0c6ZzEK0HepyQthtjg1EApHVvB9EPX+1L0Ky1S
k/XSXKKQQXUPpwhf4YX9v/VV2SiwJlO3RCsNAIFfYFZOjutCLJc5iRQby5uzu2Uv
5muwIXTxVBfy49Xh+iQUus5CkizPcCr2QE32ulwiv/G9PyIr6Mvo/+MIS5aRFX8V
HFtwutn5+6gb62Z+EiZRe32xQDoC74/C9nR++c3IQtfEuKLUiFpGiMTVqezE3d4I
e28SOxbS0ImCc1Nye+zajiHU56Pv34AB0Lq4/lUeRDC9dFs/CtzftU6za3kmB+dn
UjGAcjG5C/lISe7mlUUh1YtHz4uAvhlAhrj3eJXGRVJBsO/xQA7FE7X+Ybzsq3dc
3o3MJfm+2gI6Rru5yRYwChz6R4X6dXbJOGmXcMHZzc/MRO+RUe6xR+WtX7TKP+8n
KXe1n1d6qM/c6UMZjUzeaPITjEbp2wI+NIx+n0KXZCSEZ4218l+Lj42hHVHJao+9
QOKNbtyjBoN1mBOd108odw==
`protect END_PROTECTED
