`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fd1PC7fmbnwTwlwhp4/jTYzMGnLmktewv+uZ2Bd+SLQusn2V1LxyUfkDXNMe0GkC
nz48fHzXTMMaHU+N++Tf7D/MQHVz36l7Qj28JfJHeBD6jsKrgT53ZcDGEDYwFpnp
5glRCFdcQiv+Wsio1VtGzPhZUqwjK/6Pa2rrQ1p/ytWLTUO1pSeIuq3wq6Vyz6hI
uVpq5vqG2rt9U+FCNRC4h/UNcGlPq0sgrGybdgCOgr4XCK5bUQm15bqcTK9oRKYW
9MmRhhwuHI+/XHJpmAnWuGvB5c6Ha9Mmq9AbaQJixSISIBp+zTROOl4g6H+MVHUc
OM7d7lKugXavEzK7S5teuRQZfuij5rkMXHNZ5mX3y+gaNNglVuNHKvTJcYRBkGrr
wEebVUdezPewSdrQf85HfhytCgaQEU8kKfa7qqM6xeG6IiWSW7YP9b9U9d2Lb/tc
XpJR/ns1w9NIrePd2GgqLHOT+8vile6uleKYnciVW9pWiHFSXnlleR0qWTTw4m1j
CfDH65F50IVVSrz0mCG+EdYAw8shHABeMDdXApxFcJoA/zGPgfz5gtoXGnKPjx6h
M/CNgZZu/Y+Ap6WyLeM9M9nbJsM91/kzisFQQBOsidswyiW4fxqgNsKh7TmER8N8
9w11uccSzK6zjXZyxNXiUcEbIIt07WoLXACSJqUYKITwbu1IE49Fx/OPKgZ8b6sB
jhv6fH4j1PW4M6KkW0QVYAbg1Gh0C3xNwNz6DZK3UectGpxYw7rMnMNspRDivJ4j
MXAu8hO4jbTvLXXtgAsilp1W4Pz4kGjWgW5yYdx4H4YgvHMrW9dhHSukcwcTBa1p
T2fNb6+sDav7yTo+1XPhvMyZqW4z9j+j2YZFIa2Q2aZRtLTEWJyydaN6m6so1XGe
uBYVL2LREjGjuaOSArFmcQ==
`protect END_PROTECTED
