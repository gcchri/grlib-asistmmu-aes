`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e/8KGyOooH/tUjizJBaLBY5VH36iS1haD7MH/2t2QjTWOKq+jpamBKZM3ji6EyKH
zcmg+krZ/QPGHMq0MXpwE6mBnb3lajrxbLXb9yxP+36O0kC1M4SsABVAhdkQsJFs
2TbWtGActVloxWODMp4E5jdb0zxpmDyYkMjjCDGAPjx7CaNwLC9VHL4+gP21f8gC
geWNmS4d2u0A7bvv6c72fdOCPcIfIfvA0SQUycdOWqhcB0m83G4V2jCg03jWyUoH
wh/9XVKtB7kfgy68DKm0Qf/eGHXKCotrpT8SjQKDDTXs3OXBN7iHp5IW0B5lJ59i
FTfO/0ZXiHhOqkC0GoQXXYWuUidhnp603uplfiAR+E8QHqNgp/R9gS5DRpRjF5Tm
QZqvb7z4pzPEdubwSEGrrS68w+0s7+7Ou1FxdCARDoPQzcu0DopQ35es4rRTw0Jh
DG5vEg5hgQfd67MjyPlNRPdn37vwwVX0xi+/2mkSylilPm75ljRIoQqTkETMA267
XVNictbvv5gkWqCeHphgOOvi+A52kagemlv9d4BTt1JU84Q8XgMVpLTDB4xAUqjq
NqHO1v9WAdT5PqqedlSyn88S3CSYhyPYU1Eg9QdMt2x8lUTau4b3cZpsEjvhVIcY
MdqelKdALzYZQX3LVdhMloIb325UF98px/qrg205lAkMx0+jB/ZbEH9W5Cg2aiBe
okgmXFepsAmy+WRNcsZpmTPp41FSPwQGLEsR3WWTbnoAt8fMusVkewH00e4s1aYU
ztj6G1vZMKDvlUXGmFuhra9AspjP0omEq9qsPoo2bphFKrmPsfAlqIaFMZWuxxyu
9rjX3vj5xu+x32B5FKMOODbTocZ/sEFl4f1moZwEZF4eI/AqOuNWaSwAdHI218pk
yMTE7HD/oWg4dH4/hCDDFN8UolZqrzYo5XHJJPagIcGCr8Gu7IRm/B/s0JBwsRPU
9IlT2JzIV5BuZ/Hdq/YpjxdD/A9QOqfdoDs2V6SfnBMaUIk04DCiqELtPFbMwBGE
Nesxf+umPaJ+VXAlWrMETr1XUwZ9duvAL1A1TbpabOLEgulZBZrpprfgLo5xMiwJ
1PHfvLBNxvq5R2cfplqQPFASxRseO1bj64KKxf9DESTtjLHDWOVPKnsNYjMqrCkO
3TwVo/8852JKSXqhSeAFPO52gI46cbowtJtF9U8AimLSkmX+XAwnA6utwQgd1dYM
VPgnlbRGPg2GkVevKaurP41AYSizo5VopgrIj5G5yP3rek8sVXougX1Lx5MfV8lJ
Lb6h1wiKi7YxstkoN6Jtc60/UCeFYGSnf57P9obxJQS8kafqGfPuhKgm1KFbzqNX
wvVtHJCL0eG+NUz/q4iICv84nunPEBqSHCBO/5PkNC5cxIfFZWWdipSJyq1gbljn
MwHrfV5RFfLB1ZPHwj9rh8QYSnVbMtrU97sVOB3ybaShcil8pGt6ofTggD+A7RYe
G0c9qx/QhctSktLyBQqAww==
`protect END_PROTECTED
