`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RaiB00QwZUB331BAfAUXPT+Rh7Adeo984v6GzUHmiYeUbLcpGjmFKBx418Vtb1ps
Rmdqkx6TSXx1uPMmq4JcsO9/wF/FjjlD2LACayrKWW6RP2GehyQy4mG+SvubXvSI
79vA2vJ00YhubGGQgZD2YeVsbpWvvAXX0dmMIdnzylH7o9v2nCB/3qloBsxdlIUZ
uFvF4rO1G0sdjL/FJ3WoZz+i1BzrWzVxxJKkInWvZ231Utro4eNdLN77yh5Rp4ZU
UTWHuYtqnadcGjfBZWKS1BLW3py9faTiPSKQzfUMw56gdHlX0AQWFYW7IgDlXcMR
vBRl7Nzv+oONlpR6cnKvKQ39rE+QJI94PkOOaR8Uf5jnXACL62RnFY6sAcauGuC8
1g7kfNErrwCnUGlDRWhm7tVKHfwbCWEvK/oZHjaPo0rPvtpKWk4PS52Msy+BIu1O
hLXEQd9pRwLMf0lN2xbd7gaV8GGvcegvz5kYsOkdlIYWm/G6bOEAZrTdrqGDpbVz
GsU2GMaGJp+5n28LLKF9P6GskIpLONaHrIoalFO/GWmtvIpoS2YAHzwT0U18E1Vd
qIrv/R1r4mhwKcsQaNSbe9pEz//7pXyZY+ME7Ho/HUvc602ooPNshgxAWCDguyTD
4lTmcDKujaimmLGAHPBMhqkin77DsHkPnoWmrpGt1YNlg73pi8yEGRvukrW3RyT7
PwYaGNyD3lOEX/5bXypNl9eInhdOaYGd77h7d0njZzz+E/2/zc842RQT4yCxUdhZ
lsYAO12Zf/DDhRgaHUWV1nw02B3Ria7oB1RErwd5mFv7l48VXzXYYbxu5MdZylbZ
apsCf/JkWEWfHCCSvE8X4lY9OpNOLGWOuI6TwyXE5jcn0glww0YpA2Xj9tIZanR1
pGkwgZ2VWFaht0TohrOZ3PhVXcFM5zfAIZpq6XBHw1hqz0u46puKKTXCjWNxqGwa
FRVsvkDBQWq14usT6MeIXpFjoLy0skyiggN7C1IXWcrxEu84XftpB7fbs6yV+k08
USUgWC8ospzdQ/gwYUMXuIJZKlNLHwY+kwG+DlrZ+aUdQdLBIG2CKgGxFGzEUm17
YfIs5hBHY/dRClvT8E9OI5C2eCUfY90KbUg3Grj87RnPSMGTqpDqJhUKt8XLu+kg
gxv1RMBrxvUYYvDFlPJVmmMnhNgsvrdGRMJ68Se/R2WjnAhizoD61p4y3emtHJzS
`protect END_PROTECTED
