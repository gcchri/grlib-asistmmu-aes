`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VPkMMFTqsvtzbbw2pTxniBN70Ylt9++hxZDmtU2JLSem3iawNA4kEQbUPxpSMoWK
rV+SNxODv6gL2RnA2igaErTWq66AKHX4cPdh0FdoGm87EmuAx//LnEXXbBlMZDTg
seENrwao4Z8fv/q+j5b8oc2JSTwuB99a7HF7Xt6iSjBNqK4bAk2k6sPqJ5E1Ribd
I3ZW9UG/Xc+i0KMf/+Moe5NNNHRP7BeSSrQYQ0IWt8V3AtlxJWxcPbed40D6l2dn
PsQgSeBGNpS+wskXEctDtyOKtQEbc9a308VSPDUjuprvCmi44Eojwx5jCd3FsuDL
mru/VOo1HA2N7fYBC9hTwsQDAF6yK6xPqMhar7Tho1kd0btypizWDgwn6wxcDP4v
1FsRjzeKCyjfHqZeQqs2PL3wvp9BcpY/vaTbUEPqMxA=
`protect END_PROTECTED
