`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BuhYSUkQF5SHs/BeQBczF1EoVIgV/eJheYbvcm/7rKEo4G20BeptMWDQFrZNyoZs
m8pESi4XK23+ybfhF9NwoskzmMNi7IbQuaHS3XRjd7Fv3aXFscvhjoXkkHE+QIij
AnYhY/Rt6T3oPL+KQNZigxbOgIVIGRmoGUoZtTAiRPfetj1hTZHbJlefKu3BOpIt
i3i0eBZ4UvAKelomf4/Q2obniI8JpCHi2vcmPZOMnhWihJo4ttzw9RE+Supn0jtn
kc9NBdpDeU2Tj8rlkdZaroiqXyMd97MxO0zaCqPqGFN2WwUMCQNkhSiC5W2y1R/V
+58lIy+SbDCEnjXxUy4ZVNbVBLQLITo9+x2JGcmGq1V6JryrjVing7suSexJ8A/x
5UWwpRzU2xHC+UMsInH8r/MtqcMBSiZ6xoOOT8DRkVV+T+O/zJo6pMtokCeEeT/5
Plj0zk+BaDqLOYkEIYbbmPx/y9ijZ+LowxZFbP99yHGpS3xNXuXWeyzr6CpQONZj
3YSS1nixQTK/iIcRD+Fuvli8XprwR7wbk39cAZ+alcLgNyPoYc/5FhbLolZEFCGa
MHo49/WHnO8GrJegcVwR54BBR1RweIvuafaZYLX+5uyrPpIN/qf4ehO8sYIBpebU
isjf1B9DKfSeGQXEZ/L3UF1rSIJI4v6W+87rNT8b0HOF+5U+dcNgxb3n4CD6/3Gq
eIBexKTgS8mjlYSMuFS6ku76QSQIOOY6G1IbPopL9dA/T6WY1UFojh0ikJBFXOuf
JuS+/tSoAVTUgZsmt9hLaJrV9zKd66suqVBnWWvTsMhytWrzLncMTqHZ8w2Ao8AW
efXphYf0Q817xKzxGipq8tAcfxe1p0/VqZE2c1vTWin2p4sqWlc9ZM2tlxQNzkdr
iMflOfq+Dk0nd3KPPifaChR1NjZSHYW7S5gyKklnfB1gKxv5B4Jmrh/Kws79kWce
0JpibSYz9wwFEIcwUe9eEZL/OCOg9b1aNSbWUaQQUVD9HGg6DbYyTZUXUOwOfPga
fhjU6+wo4DR4YAB8DJziJlOTu+uGL1HCioqHT7evPTKGG+vQmSIYHv4+fWekBUXz
AgzEMWN68EdWUpc+dUhlhdXQfv+VYmAYqfaLL8jD07e00LjbpUszfOiKl1P0Mku5
Ot0a/pYUIx2EU06ubMY9gEKIh2OjLPwEmJrBpD298VpCIBvHanMK9Kkdkl6FCh9E
yNCWoJa78nOsn2ddFLQD5i1XdKn9bw22O/jyCC9OOlSi7wuyQl934ltLjphtKYDi
1nUqlGbcm40vD5TaNf7mZ66FSdtbncoMOKbhxN79xFJnY6VzuEFdxNjak9AfTiL1
mAyBOmHMZJDxAwwso2YH76KGoT6AaecBKuAS9o4kG742k+7k8E3tb+G/k6vNDh4k
swfpS3U1rVZMo01b8ZXVsa/0QRIXSTcRhTcx+ZXJyvG5ASjdJshn0af0NAjRTRfZ
bX5leLUpJn0mPNChwyoFbhahKLfho1NQF+dOOLfHZD0QpiOgdMdnGDUqmUKvQt2b
lHGTSHbnoV3PG+bkps3ClCdzM0F11aLSiRpvhGRpJkUNi/RefrwEah7am6SW7KZr
TmcZ8C2CaZzMKj+kASAtgdrDKubHpG75MV2utPM9rAozC9ZEJaX9eJphTRC9cwbD
qK1sndG5nGeww93g305wZISoELvDy3t6yHzo1Q/m8NR05mOI06pQkDCG96nHGkVm
ZuVrnJPuB1TvtLATYNULHalrSzogOcOXE1qhhW+2Ro77mTdT7I4hRNsXJ0YKpXlJ
YiwBdYu3AZ7rW4eD8ycwLTguWXh+rnRw/vtDtHajjM+N8Mk0i13/eoFJXn+Iq/dT
gQ6eCqfFnD7op44fb6m9G94W+uzvXHKcIKzE3ntkgbrR17H8JR0cRPUfViUL6PF0
E1YmpFRpzYlBs5sNHaKYXlsA74/JLRClgBn7IY8pcctqk3d1QYrYlIhGrxkjFTtc
lwqbT69uBGDFMpEnHeW6seWPbo5PmhVBPwJXMihdnhABULH5HPsGVpTeRbbfuhAM
meeJ+Rrmp9B7+pLaKgSMqpdh+/K4At182K9WzZoDJ42EqM3Eg5qI64a5tBFQLFrP
73TAk7T6SXeEnyFipB6BiJGri5F1VN5OAcuD/0O/bKFHk8T558T/FXhRs3JWyaUK
G/Yd21PC73B5U4OD/dCHShzs4dcRTRoYVWWIjzFdoBXgt7ynA6DgidcGuYJHkW9M
ZBkuJpnY2+Tu+d88sdSWO6M+XiqYs0mw5DkFYvT5DmbTT0fmHa/1i6B+QNB62/bE
zPd/gEW8rG/jH2m3UJH78ApI1/Jc8J/xjMTS6r/IgddPObm554k8U0dxVZbJesJB
1sdDba+u3s3YqH7+DXDcbWyuQlGlLVgb6w/XlC5FR9oe+4oSyiT+eC6VnQ8zJ8BF
XDFZtL+QMWKsqv6DPXw/CkY6CeQ0eXVXxDdfkdnxj2s/lznWb3FMGy7ibZrEKi5E
rAw+EFmi9yiTpQpC7UbRZEPAIVv1cOPBRQD3+lEtLKKpbGhJLkkV5p+xOGOgXTSw
PJ1VOZWmjUz+FIBudyjFx5wDLUf4JlJe/0dqgxTWe8sV96gk8UffLhty7Na8AMka
QLoSrzuhKt41BZdeZA28WstH97KADrm5NczagyEoR0QPykaTJqi1JBNTqriRttWm
wOJSbX2lZex8b1M6LA+/Rqjmsde0QQCGVdeRnlAQjD3wJ9l2PLKTo0R4NrM8Haq5
xJodl5Dvb2BKLLTlAvn6AsUkTlHyAbYct60WPOd4g6yUMx0H8HsZW1gjdtl+ePV/
rxVgUw5wjeya523+9qE+rhP3NvVFDV6QVn/HS5xm2SQ7QYQ7DU+OZ5DfZmqt8/SU
fWpaVROhDTiQ+i+vatoMaxZspm2HZUKacyO08LtoFt9jqX+OJek5l67JgtiYnJV9
LANrgKG8q9c0lKHIOY8w1uStBaVRNGzeU34S5hkXCwSb/pcRHA16usBybB1mSY5R
SQtsYIB5Tg9cLoUNxp0sVDY+5xxVFr1q0SmcZtC/Xdb+9G2Pas+IaA14FnIvmSle
I3S7j2XcMlihqYsAFcZCn6U+YgmELicNfgM2jWdSy9Y=
`protect END_PROTECTED
