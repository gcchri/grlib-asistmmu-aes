`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
veOW0U0n3xI6G5ZrBlVD1UItaT8NYjc2302hGjQw4ikoZnOtNoSu/ykOJVm9vwyj
Z/5j8E9UKhSCIS+nAjxGlelopiq1qClnNsFRAmmdSgwWnMaPiLpCb7XlIkdqcpXf
1YJy4x+nuPtehE6SrsfUwWR/H8EgLkQqrAbwGTLL6vTDIuBrrvM0axpDz7HqsQv9
093PaAI4IZq86GzhsWKuQ5nF70rB+VQa/iAhKX1B8k0BzCxoQHrk1UfVMtW1VkD5
EmycrM7/Oars1fCj4w4yGVAxe74/OHMqCwRIlD4OeWbs964BTtu7/BcAFkR+edJw
izXYNHLUSQ+M+GZxHyePh8v1wdwYF6KNhgWDTJnO+bVZ0yT+MGY49cxlpdanXQFQ
kZ745E4L7IZ2AKaLdcgnFofdB3BnNeXoeMhAYbcW0mHHJJVY154k/Bp+tWM794B4
N6OQqB8ku/Xl6MMT9rziz7zUkbQRJqtADTk8PCrCW5MP+SWYsufdbBIwIuGCEUlH
yderT4WHz9kecoUr92+tE6zKnT9AvzdZqBUCIE8Z6MFOJXbGNk71suLf5SBC+St3
NIvsaFP/4LX480nlohh/aeqpNlzYwVhSVfiTbZA9dRPH/fJaDtwCZA6A/xkUPIn/
6L9wlDuen7OgkqLCoezWSDwWetbY2WJRiK3gmntwz1FGbJ8wnEYwlPdRae1TwbJv
LBC7RalwkovpEUdyIMfFfTPEB0x167k3NoqENR+S1nsRS7pSvAlgpgl3bb5k5URS
msl2E1P9+ir1qZuit2piUFCOxco8t4Fj3eO0yKUCdvzrxOEi0aWxRagif/SLlIv7
DUluiqby0g9Yk/J7pSGwpWCqH4I5A8p1ChkdvN2xjljXAdGnuARHYoRqt+nCcFtl
rssezMHEticOct51YeY78A==
`protect END_PROTECTED
