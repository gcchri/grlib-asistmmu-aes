`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aG7UjfFp7NilXrizLl58jB/2gMkqAIhO4NL3qbLvbgkNPkIdDdlkVKKHXRpMGzIo
jXwl44nWgSmCliKCuC9S6tAZRvMAyeGsLAWDKj9iv27yfdlXrnqZxEnmNkCyEUfz
+mASN2ZXF8tC4W1+99EFkha9vRucHETQbDrtRhWz4j2hHby+gtAAEpjvb/Ujz38e
PbVeyeEk3t99nYlxVCyScSQohMtmjtyvIPJJTD/TmmmnWZRG4c1u6N7jO0nBhzbd
EEAy1qw4iZhYBRuKW+8FC0gnTgbU74cg6wfU1vHPWUDef+SWC1AWeYkct1uRHJND
`protect END_PROTECTED
