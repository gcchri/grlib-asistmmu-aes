`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4vJW5qwvJTQfLqrePZYLdyG0RKt1Q0RfbRgwrykZkElm9+xEY5mUy+9bYRYgEvY0
uDSt2sCThqDP5R4LDhwVQHLArca/51RRiwSL2s1Ll44sgmjQx6adgYOQUq0N1/zy
LOaY/XLjTJJGzK3qz9rgmC/cAQkH9yepHKQ8IHiBThrfbPVSX83NkdazBW3VvwWR
+Yao5mrU/LYRlclU+l7i7yMjHztoRiWjP/eFK4hamcERPFGe3+zQSTP2xuFIvdJF
geP1gLOcO1QXaANTaRbGBbeY05tmbzfIGHjpmodlQnDSEAgn0pF/lTrqBv8/pJS2
xbIHfJ6yFRNBGCBj/XCJOfP0uqg+MmIjxKdRvXWznvfNM06kbPe3XubqoHbvzGta
XnvvYIWahkFWH4yd6Kh0/h+S1C8V13ApevG0Irnwl5aDwnbEWzrzds7fd2PwdBQv
NWbPIqEhy2Lieg8+W/NKIWdhYwpKnnGJssd9Tg42k2KD++5P+czuxajOX2db6xm5
/WqWx8Hxzt+IKXvkKcSl50+9cE+AvxipZ2lDy5Rpg9Kh9J8fuK2fKo8k3WGrl+a0
ThvLZJU5gKaYGUJMlLBOe60pytoNFEfLsQuQU3k/5NM=
`protect END_PROTECTED
