`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
97Z1sWPJs38HDi0qQWqrvBCWxUQmC8cpwMd0EpcSsxzW7Ui2QqcBl5yqOMgtTcvx
Sb0gD/zaBnzRjW+oyaylChzcQtD3q+cAov0sFkMObmcDKoArzVIaxsgTSC3i+33s
ha6eLE2gpOFscdnVizJpVa/YH2DcQecKcuhBV/6HEOi+9OSG6KK3zVbd3XVarfBw
vN/eVqQBVRAqdKWpIivNx7CCtzC3VSJy6hPkeGfOEyC8uilENRx40MWxuUnYJtS0
Vl74L7YiHPWXKsDL4u/+SYhv0k293mJ0/6xyqNM1M+CpZgcP2xOCYXZ2mg7uo9mK
k1TupVRi0Bytbkyfs28unWqi2h74PU7UIX7N8GOqFl3aCS2U9AV2fBtXQDMITDsa
sjNHO4P8wfT2Fq/WdACLmt3Ff7+pUYLraMBt3jNwCoDwjnYk+iLnYCwb0NF+2FOr
u1CIEeyTcSVRy99NZ2p23HsyAryALUe7U2xdlEhCNvDhxhaJlnrkPnHYteb2apOC
s9WJWRZneqs3s9HFr0MDMRaayr0SoOrbSCtHVD5cAHFXPANVWeWzcNGNJ/eLsr1X
D+kktMOovnd5EbnwDZ3fig==
`protect END_PROTECTED
