`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ehrKVly+kiBK0VCboEGnERW4YxepU8HTPXXvbYopL3yzktH4LKrQinHzsYT3MrNT
BfN9o8o7WUsqQJ9syIC1lMZTbE/sPO/uIKo/jelT8bWG0Z7jWNEZrY46r0sDHVx9
8hrU4PoNQHkC52ZH8ptn/RFGVmEMKOyjbDESJc1kccNPNPqprTeDtwxb3buAMNeW
XNrbkWw6MfsQyW068Pv6Re0G/V0KCqMmGVGBrlVrCw0UF8gzjIKdNjz0ewz75eES
5RCQPdznNjAsxxvs+3yY/uVUrunwyXQK1Mx3Ewje62t60zX4wvCQFGv/SDZXjnmu
wdiUlhRIRuzwmQYPxF54dKkdeSxdzwdOR98ZxtCPoGPRW1rUWlEZKTZBraJX9s+/
hbLpSHli9NOSI+2kVB0TSH/STdSjaQ7x7nZaP9k0JzmQ106exlz6MNIJ7H0PfHPu
1EBvK7acTWh57uEsatG5gk9/nZXgKJlFoxe8jH4n2N9U6U5/IiUTwLQYZKi9i4Bh
VwOoAuZIKfNL50L8IgBR/P7Zr5YFM/qBNLw4Oci3WL2G26pY9tmXphoKWkxzXey1
UDfXI8MuyB/4xOsKM/mGYg==
`protect END_PROTECTED
