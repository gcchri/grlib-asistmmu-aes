`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RT1I/lCuYeB3axWXas1gjOJkjJKL6nZr/SXNMFhiMcQZ6kwLA8G3Yti2IEwcR1Q4
mT5ec6271g+B/dmM1H/8mt8KI+w/kdCx3Bjy8LjmASFo322ngspv02CpwGvwWFx8
7ttECtZOn6ez1QBiapk5BWUGiTSMJjbCXZl5XG1Ah1qxXQ8jsRPIbLJVdZYK8aeQ
tmhwEknsnpPZBgP+zDXyj3tWZyQZc3lD9/DK2Gt70CGtvJS1bk6JGgon/Q0dPVa4
rx+AB24DUFh++zyEwX/+Mxy1d5DGW6gxIMjUvUh9oz3TQuqV9SC8YRWPaxWwe12i
hwgOPbY1qTo1AiUjPuG7dvsW/y5I89xkMH8WfoWUk9geFWPnAWD4Xyneny7sGYbY
XBkVKQ/BHtF3dkYiEEObj2f7N4CDSsP4zzG3FqXKavBzlNy7OnTSLH9JxNzr1TWo
vioT3DuV51GVn7AanZ0+uyfb3xeuGfCwczGt0qFp3j9IBj1QduWiis1E+lg7Zl4a
MZ8A7fSYm57UuW+f5XnMJX16dfnKHiL4P0b7KkhNebCL17HITGrhnJInHiryfVSp
VtSitc0G2gA1fU2okOzlDu2rQ64dSOly5hpHPucBjAp7nwHM8U8YveiFBm7GpJxD
O1SNjsS9fOjWDGweBMwx8NTNE9qoYFp0whBXj6jK2QFXyobZ1iJxbExnVFAKxMXC
6TbRyIVgBu2Z895vdJ2h5hdNRIdQML2VHdfy+sMdD6dWfAnDIUpb+seyX1VHurwu
Lw6t3X4cny+Rt3YSk94vWEeOw7H4rSiZFSAtonFl1/GvRRt8dQzU6QmtabgTZkHC
u5plIkW8srN3yZp+5HwJXaNQtoNiICC57LYwOSqlcLsVrxICMacNsICkKU8Ss7z3
i4DHSO7wQSyIQPd6x/Zy5BfqBxu9ODicVpOEWGesIin/Op4Tv14SxnGn5PJSbbDw
Vl7I+LPjTjSSxrfsezI5MbFB0zs7syN8fivf+WuMnLVnSUTAwebrVVnjhNPL7dvC
wR3jbbAgTKFh6vNlsJlOAO5r/OuReAYqBM2TnT7R1eKS4pzTgq2KVoAvqslcVrmW
5F7t/dQacohafjc34GGtcmrpCQZ/LnkgLJsENV+Bcs2019x+TmI0bIwX8GzMVPFT
CgFtvwSnxAQnAmbVQ1NVU1BngkGoWw3eDoElmZ4MPF43CH8j7ifZy1xiJxl4azkY
qiWtDlbFtrIMBmJlQe6xZmZXpWKCGCDME4K4tgeFB8jYcDffhI/uTlNWVxw1mgAK
qj2LZwh2Mwbb8FaNKe5uzPL7r49dCdxTZ30FOPjYN9FQI9ncWQZuPgK3sWUPXrO3
nSjVvvZb1cexOfcBxqPDIgUQ3KjlIpaax9uhJrQ87smd8hR3V8PB8TQzWhvO7+GH
yk2l1ZenUx6VsTWETm1UViV8JwbuB4g7JRuleOIot6ACRKVdo+DocaYgVDCuIYiW
LDkQReFx3d0S8P7RapYnTMvF/jJaBHmedjUJ+mqhfaXSPaiJ3xSDtqFLibIeLugR
skGT0oJqH6z6vrKkrLO8yQ==
`protect END_PROTECTED
