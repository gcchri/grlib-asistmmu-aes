`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/w0yOTPigDCQl1o/R3sYBYzg4COHJTiHiuUucFt7sfdUOcbtIXAXeTdkDsVTF7Yj
fGXw8ZZoeOzmSIlLRF2t+Vv92wqOpviKfKIs9Mhn5kppTWpe8tIMRt9SxQDdYcOh
RgmVNJvduLbcgzyDEONGkyNF9pecVIohDVFfwhPMl1wNbn3qDwIAAI8yj0zgWE61
N6fA3m5U8NJs/6d5rvshlz0tNd+XEa8sszJNupQInLTRqCgNSgfKIrWv1bh09W9T
cra60QkZaE2VArllAXEbCFqkQGuHqj0ldmhGlg+SEygjFcRDkRaLbsYmpniSJfHY
Ky8hK1wJK+5SUAwEqza2Cw7HfWx7CtxIa2SvCvzdOn5e49/TtGF7R7L6SN5a2eYz
LksGbXvPdPkAXY0cBRHFofSSY++wY+vRMANxe3BkLkA=
`protect END_PROTECTED
