`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0qPe80INoNJ10/O8HAqM21z+l9kWr5IsJZZhMYDUtIKse12cewz9lq5L2aXUbsjF
gpt/1v7tB82/JzpL7Nd/9sHrUp/krHxHrublsS7p2n2fbDOjOfcsG00aubgEde6R
42oZi8KYQWxj8R3mVcu/dR6IIFUfddPoYMufhdcbkrfV8emhnYSWfFdv5hSe/t+u
d+RIAaCIwyaHHA9Bkm83DTeF/m3gguqNAfmE3DKwn5SoH6QoH15YRR2r91rn7ksc
G9F+A/S5xuVCUgu36TDe+Tz6i7DaSPfv9m+8fTxY2L00XxsYDTFTkNv5MyTLM5ZH
akr4Fdh56BDGMMU2Y71AI0E+VuiK1oMDqEQoeW8qoYUn1r3+IXjJo9dCYSyQoAQh
VuZ2MWBHxp3YtA5ntl0/vNlHjhygCoBqKJkUcgCWShbVqJoPpAsW0I8IgkLtMzyS
sMJj7DddfgveEssCvsih7J5YGfLchc2NSOOoTq0/lpsKELnhONrw0tmrvtahX9V5
zZJT68D9qKKtqJQslzm0UJToRTLUqlDrfOokNZ7Ei8hbMigx4phPBTu0WtfdMvOU
GD5rlsBou2evOpOZXmvRToIu2k4YOzePmiFi0WqmRV5b3i1KZSwKSrRYud971oCL
B6HHE8j3JwEPL4v+ESMjoqv1Mlpw88qWe2O0W+KT1baoVETSARCP3Qon4KQsk2oN
EthLVW0wqjI0J+Ff6FgFYVMO1UEn6EqA4D6JGoauFlLBxtlBE8GVUTYgT4r+r6/F
skmTULbOaR78Q7urJ0XXBq3oK8SV0tjz6ZE7zed6OACX+BTO4Z3HO7Y+XaM1kubn
zX7Mr1Tm3QqQS2lWGXQYkxJVpony46LVCOkseYY7Cb14uIiipYzyd23OMf9cfTVn
7n7E8j725d+MutoVgx97dV3d0S7miry8nNYyPnWXGqZ3wh9/wr/jRHYc+9VFJLwj
mCbbfou/QMq/TF2ZdsUuNWM/JjAxe859jM+8CRWgZOlEaJLw+jrxLz17LfaS3PJg
6HxjLH5mHV/izXyrMeWlIl+v5Da3Kr2XtX9uUeXgWIOVOALQH3CtNwbKbkp1KdNM
A6bdM1Kaa0YOqCEuYRVslGw6/+Gw7kTq+hwSU3VgM40jaEX/WePRuM45xDI7GBS5
y6DzTwZY4ephpARq6v5OvGOdG7h7GcP3k/Zj7nPTdKge5zAJIGb+g/nPKrIu3KnL
V4dizcSrohZmjpMCddbbphgmkzecCSvesrNYFFzAb1PSN6v8QR1G8BcYiikrh05A
9yInvziH3jM6JYtHHsedT8H86W4fVoo4Jcd5S1MyRS5rrstSU+rjG9BWvQcpaawW
pRaEf8zmunpwV1x4AuCShI03JMA7ggeEKCorjbKZUgK9v62NQi5eQFxohBfK9K6K
G0/6VriYYem+/8ARmxEj/QTYW1xRR2iLZUCiw9on1R1z9EHg6FC91V6ji4a+lkNV
QeU5Nx1cu/femfC58v0iucfXoSv9dpYT2bArXJTmfiyHGVvwd+aK6eCvkoJo/jYs
ii9zSF7u421308NCFumjPcciVSOn9MpxnTWMvJgG+3NBgxvyvvhS3w5PqzmF323O
r9iSw1r3R/G/pOmLEGlVT/plOn53BwD3jnrU7RMl+s21aqZ7U2s3uaCqDb8EAYIf
vym/qUiS1E6Eh9G8pbDyiRATHrjNaUIinkrymrQ3h7H5upmSGngntGWNiCE4QKYT
KZ+owTkKh2hu5lvjAUSIdBfnk/LClR1rxal2lkorb5BrskApSdtEoW/gLIGu7r6L
dlYoa5rCbf5B9iV7DmHavCR+jV+mk78Pf6vAHrhxybWW9TRjFxINYVckWJXpWRCW
o96zT/kU8Zr44GDdLilppwJUFiSD2maz3kyNCGvjzWXo9qivjeq8TGoAoI3OUbdZ
vfOiouDYLBlSPXFLBUh6r2QLYhOn2LyT2fZ786PwflYaTLXxw0+cekmxwyiBsl8v
mRYq4/ewDyt/8fSrHZjsTzlMlCJn4hSn+pnXS/mo/ReGxLatUJL+of6UJ855tu2N
8kHc9N5t2ZMvMs9ELVxdVxvd9hjexdw2ZzKqOwNo5i7BUULikj0ceIXmxnvPNCL5
`protect END_PROTECTED
