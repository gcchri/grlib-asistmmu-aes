`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qOgHcWBbVA15k7oTyLHygiPZqAAQJxJN9tpyOzZiGcNN3H1pu9+1k+/oZsyHbVJ/
a0wkAdCsWMFxTy9mGKK6qMfmIMACcc5HYJHGtEHIEZz9rhuvGGrH/l9CMsxVyYBr
9zqwmSOZxk8x54gryvMgliLxE1Fjub9Nkdxw7yuYth43CynOhm6OfcDO9DAQpT0s
6GXPwHVNnbR1E1oGAmufITly+zSZlW9ZsRRC07yRTGyDT+lG8SW1ywwiBy7uX0eM
/ruh4koHyY45hKLmtKPEIh9dy1abCSCeuX1wxLUji4nCfZQDQn1/fPdrjAtcprDq
5i7ETaSGcrHOqng59SsJ/fBkh4PpoTQ8k2YL8tMhYnFTmOmi0PaAVF+eSoDSnrjL
oHaxGIQ9QXT1lfMJbw4zNQ==
`protect END_PROTECTED
