`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Eml8xpTZHSLil5ABGZwP5dpT9ohDLKR5/WYQlDtUgUpntjSK6T1pBY6KFMIwyryg
pQMPsuD55agaIrnma+j2nanepcy/poHYbiz3eDEaZ9CNoGQRb/SnDFjK6uj75jJq
hRBDzt1QbE+Nb5TkzhtWOjKeIzlZB7Yr2kwphr4zHFjQmhsLBr+RBaKNxbAuRoQZ
LPywvvqBqzsuCxyBKSusCFcpxiLM3intCylIY1CnBWnzVuz/ypW6HSSXwWdoIdtg
DQUwqogFS3T8uTdAZ4h6/g==
`protect END_PROTECTED
