`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4fk2X/dH9zMKHYlGu2Lob6+tjnOiBXKht6SRYBFpxxzUyoL5vYOnS54CXjkl0hTV
2aAyeoeypOrNF5TyC7z+OcHKoAtMyYeRg9vHeIhy0T4YZTpgsseS6cR3hEPTRqj/
SdujEErOuDPZmQ3AByTgDRFQUIXNuTGzkbkZD06ZFazN2wXQIJ0IWGBlJzua/mfV
G3IYmeycPXLL8YjYKp6eLSxOW0ZDUSZgeJviZZWZPkmx6nP8boQbXgwSNpvgVd9K
R/JZ4Rhe/ocQnnFlZorT//6FuykGQ8wotuJDg4T5yRRGg3uwpPefCqamIKRo7TIn
Zs1Cg6n+H0zFWwBjeRXFmj/6DpVmd9Uan6SZW7l7h2loMi/wKcwr3IiImXYcg0sD
PUEU+Fda7Jl/n1lqum4nXH2Ldwl7Xw9/WP1awusdJJHBAhN40KHbGKyKBXAmOFi3
6sjHaSlrrJhq7JuD8AMyU0DqKtLXSqgKdjq+/v1Fo3v38GCDcgDZf5jjWS9NccAo
GrrNAZVFjmi7+tyl1ZavU5Jh9/s8/27MkGnDLqKESdirmtUzV96B4WmaFGdM/YJH
bm/C3TMUm3wIY/wg8ETBaj7nOFtfb8S+ScoxNVMrWf5rFwmvP2BjExTYLn00D/Pc
19aS/pVRNG0sGNwEQvvZRW71MOeNjNnZCgs8zMfB/kTjGpnW7V5TcqiyCmOa2sjE
RfGkyIZtRVmyMZyQjPGGoaSfrVO4R8X5desXvTG4FHCn5HpWj3KnBtOFniKV3Ia2
agxktF98eGPiRp2Cal4D2QyX5Hut5N6+79cztQWr+eSTtRukPBF4o91mwKNDIbwe
Jr3j+FPGYXy8nhoYoBb0c6UJC73As3HB4cX7r9pGlexUFtRBvLfNewLYZAwQfL3F
WZHoOFsMYnLOrfQBhCadmoMLa80Oel0QxXOD1HuuA2JTlfa3LtxOmY/OH8npyYN2
5/7cWCEwwzkzYULqK4GqTH+7IDoonaFAN3SOeq2OqqvY+6C/LeqsKFzuTy/TKshf
enjPI4R7KmN37UTfbtSBpOKv1nnOgkqsZbUM2iFk8kTKLTMt6NGg/4E1m3ySLqdS
mhChyNVLyrrhmTmKEaH0x/3bbR9Au11SAqJCDX5UrtzTxR67VBSXRegWZ/8VzPCE
4S/4Idl+yBmlj7xsAKJLTqBNvyQnD/DZW5jbiwLpJLD+9X8AxDZh/LS3h2qs1tWz
0zxReyfkCDwLrzW+WD23N/TVsYDKeahj+eThaYv7mNg/HxnzhVtD+HlRF5DTFsOb
xmMsEm7nIas1zBxCrO4yDI4Em1HpOVFSw4ZFsdgS2pbFCAIXAVgsRZi08dJQnprz
gdrpQSNrFFKHsf6IUwAvwcMwtNBQ/YZqv8XApyHt+NS039pPCiJOMD552fzu3VWS
hNqbqCICNumFNa1TcD+HGe+cNJHYDBAYugW+gB0AWz4PEGEZGSBfl+N9X9KPPjRe
9J6M80UDyAWrkRQJRwS2VBiqLB6ixvI3PSuR7V4ztfg=
`protect END_PROTECTED
