`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+5UfekFve/W2WOLus6c2c1WxOD3HUsxfD6LCg3U7Xh5DCP2gYK+glRyr4ODEzIUA
ZlIbfZWYHw5/7Kxlq4pZ48q4DjyJALsKGZa7P/hpzMSFzes1fj+JqN5T5o94Jxk9
lT6VFZkwB5xAkIaDf3nnX/r2ZnUGLYvmfl19a1TGHSEFFkPrWoGwFtBKKKLYkW+P
hbYqXoR/I0G3Ah77KAip8uM/DiaqbaTHPN1Gmk0YCIK9eWbXQRmY+uiSt/pjKF4b
0b7jPJ21rZEPWYq+XxxmK6lPLEw/xzh3a0zfDYMr2QqsUdrats1FscK6CdQFw46h
mme0WgXTQitDShg9vKSSBE/hMQy5H7Ycl7Sr6wqRmurMYB12SZ27VXLCT4X2WePz
bQ0DeZNQ/bhNUpgW3rAhiCdLZ75uX5eORm9s3e52F1GHByU+OaHiAgFTk36N2FRR
1E2tsOmENPgtq6RplQI3nR8fAQy0806V5HwSTeytAhPttHfHeLe13saXp752MB+6
aua/+Yboxwn2zGP6wUuNRvl+wEdJAvhx7Hk1JhieiV8PVkDPXukJahfc/0y8NQeM
`protect END_PROTECTED
