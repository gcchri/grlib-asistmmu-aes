`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hQ8HFFNO5CdywYiVqoTzS2xZ8pPA5AKfjVkaKykzAza8K+2uFO4bKkfqz8XL6YvP
y0AqY9Ih6YyuXPDK2YzCpxd6B06zbUELpdSpKV9yagvmHjc+CSaQXRodYB6b11Bd
BA7lxsQ9/Lm4JLqJvhWpWLd+sMnXwT7SzB2HjKx6c702FA1UHTbsw0IwQF+GdD16
2I+f0n0gNcMlGOZfdpjLlEX6r1gwPsyR2iRZkZBCnqclMIpaqb0oDlY3Nch0qsfj
aT3mvd6jEKQam/HcNP5xK7AcKjJvl7NV+O4xmuDVCaqfODFY9JrJyVLARCS+fw4r
b/buAyDHCb35nYGFfnOJSA==
`protect END_PROTECTED
