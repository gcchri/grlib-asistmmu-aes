`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G6/P2p84QmFsSQ3w66T7IgNjlROL7hdYsI0ntqquU5NZvKonWgaAbD9EhCJGHIDg
gqXKX+bQwHNqiu+YfS4aNKEefNfa3xnJKKhSxM8IWTknBUGM4/a50Na1Z8FCxtPb
0fPA7hBEJz1YiviDYcunZMG8wYuvt82opf/kYRfy+VKuJWYfdePsMr4B3NRLYQsy
IHLePMgo/a/AEu5X5g2p5VW5O6ff3isUzK541hUO3T+OAjGI+jmGGUqdjogMbW12
rQEtuxxK/835k+LoZlyka6L64j1MhdWEYiuLf4D/A/bzq+gSy2i5UFlLwHuQyAs2
BUfbpjmWPEPf/3VVuOTjZG4qvkx4flyBfh95+KOcKnha9/QLwTLUUMfpDcQrjEuD
rvEzHJATV+aQMbX1hJwS4ifJiWdQC+e7ZIzTNoYaLLpmRKSqUwRb626s4rfblUdn
TQoDqJaLrWc1ITieI5ZTN3i34rbtm5rbO30kCRyoL/Po88oLQB/yqIIZGz/yvanN
bTzLBEnJ9dxU/bNefM+/cLdd4ST1dOKhVcjhPteXZ72xxjl7+ZDMe5Zj8tB7evNd
0AZC2c/d7sSCy12f8rBraXyBaWPbnmXf0oDXcGkWr+/iCeVSssGGjXuhmbYpdvEi
uX/wPKigNlOAcSFx9KoYdSkZWE6eGjfDPbAA3WVd8EXxiRIt1/TBm0rQ5iCz8D9j
4Q/Yo6S6rpdZ05Ph5e+1S7mhpk9lT4RPuqQoCwclZc8y6ZC4fL9qn9CvPbUeDRE+
xDgIsQzIZ/L/OandC4E3xh4VxO3YG/PGBRorNHWbZKdh/3ybAfFECXOS8p8a69Rz
nI+vTjt72UCagqaxwzCXRpOVVPnVtGg2Dba7pwpY8p1my2y6Q0O2uZY4Qc6etcS/
lTbFOSUzi1YbU4tROWIRnRqkV18dQvV1C8jDkcWWbh5SxnqmdNGsfu6nXi21xA6o
S2cVKGm/aoN8a31WyE6ZUcEM2ePMUDPQWSX1AKT9R4fiV1sRtHSQGCTVb0IHbm2s
zMu0nOI9gNPZ0PxIumXcm0U0Jrg0ntUAdTkngHQMPTs6Tv1v7ROGelE4NJy+jBZ+
+dNZ3GqJF9GNPSXrc9wCXS0XkkacIkG82MNWrVG61c6F5TVny1UaCQbG8MjFy1ra
`protect END_PROTECTED
