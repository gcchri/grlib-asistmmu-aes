`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wGfOIkI8KBZJbUiMbQO39g/qLKF40QEFCzH+FZ76o94Mmu4YsXa20OtFqUg4YaPL
BkShrpY1E2D8n9carLibuAGs78ReopnABmGjVdsUUCAV14+/KPAdT2uyLE5JUtLw
q2k0Zr6AZJyWNEhOroXHDRi/Go1C4ZX+5VYbuC1SepfudTf34TY5ugygvFxnuKjR
jCsll8xff5XX5QiEmF4iwCKlVBd0g0NngXXDq4IvUOKk6fwy7LFB2U3hxolRe9BW
I9UUX0T+QXqIh8ALEeBCjpeJ+UHlhPGA4IyY+1/6usLWCjzjZ/rA6zXLv/9/wEai
xEjN8vAht8GyEfZ8x9IDBkiKAIFq2oN8uClhLcTM09x32QBFfSk1mCGNaysUhN9t
qUr1e/KulYGVUW8rCeSJ788VD03FX6rXj6TaDlcnNL+ixwJr3m0VWiGCfzHlpALG
RYwUe4RNYTQ0r7y+1+y4cf72q3Nl5FQfvMm+K+wecRc=
`protect END_PROTECTED
