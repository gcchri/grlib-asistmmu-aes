`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D0rJNQj+OPW6TxXD6Qy1fgnnGi7WpIeeGpDGNkK8b2qOo3byNkXbdmc7DI52R5ly
IRvK8YY8IjqhHKUKNrvdvusYRKSZPaOoNiGVdCTO0oeJ0o4jas4OPC4vT+UTai2t
MfGSlIKaa9enUlTIbiI5kFwEyLpexK3+BlRam7rtoBnihIIYFSbNbZQM8GpPHRk0
zaPON5R1cJ3gt2r9ZJtPOS6ufeT924O+LAtjPSP4y+0LyYFJS6/rYsUBfE6AS3Kh
YUFNtCsXN0wz3+WX9xrHP4oN+7gqTxS6gKzNBLPex46AJDOn+l0nHR0jglF7tIbb
pFCHaIiuFxVPEN3ShLXhIs+Y7TpUMQDWBTCddRSGPJOX0LwAem0I3ppRrAxs9o9J
3YRduaeS1HTy2mfgJDNW7wkcOHXDKnMUjznzpwAL0IWuR5FFGdzi0RDdOZl3+P0j
gVlSzUZqSwsZQjJBAI/OYwcCGu09LFhaS8S4rDkdFHsUeta26/aKiTVsI7OoZdeR
p4YapGS73opYzMQoOqWfdQ==
`protect END_PROTECTED
