`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WErtq+mxQRUlniqX6Q/U1BdjFkUfJFZoEIkhQWYCs0goiEpcjCNoqA//Yov1Cf9f
S67EeCrbT5IrC70IWBOsepucapqacZeRtcV0vz4MnwgCNMfqEsG3qhRrxQOL6hwF
IO963nk045A2Q3q4soR27ubwpm6Y4WsFPpDwWVVsERtFSb1s9PxsWbR/J1EVAMkB
psC090LRQCYyRtGC8TJWiYFjtr4VaI5R4+6Z0i77Y4JSwIDcN5xeffMkbfQnv+P8
DmNSfJmB8bGdeRfSghUwEmEavpI/pD0VB3Mqgn1Ye+/Ro/Dh7O64jeocSlfLXEFN
UEzj/cZK2oU5EMU6V9horRnQx/b8OXF171ERYUtsYjvsmcOQ4XFoO2l1XGcCsBXw
22A6mbm97jNourHMnNFhVso6prH5QRj77oZmW8ZSeBQUFOCmtlSTDiTVHqvERKwQ
`protect END_PROTECTED
