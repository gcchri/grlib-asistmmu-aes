`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r8iulfQNbjDUYi/tl9jKH85o+i/aXu0aXReZav3ERwJ0TZJPRHW+RFcPYkXli7aD
bHUhSv0fvCkPlGIyqXr6naoueBSP3rVxHF3LiMqcUE/NYlfvvJmMVG9lRVun5Cl7
Gtg1dkB8lJImhfBK9/VdkenjbNnJh4bePB7gWWAHX9L+DN5BqzZRquMDh3pM/dcl
VjuDp0yrAO/LeF5XnY0l8FrFhQ3xmFOF8gIlPL8wTsLmWsyVtQT/Nz86R9Gjvfyw
xYghRPHl/4+hJemCD++B1waQIIFDqcrK3MEVUIWMCpxEklLqCSRfo2yAJu9VFQth
+xE2sAjJhxYcJwlcIBPh7cwv7xvYiYLGe/ICNETkrfAgAWqSAFoNM8b9flLJ4ehY
W67Vtk35jws2X9ZIcrB4tA==
`protect END_PROTECTED
