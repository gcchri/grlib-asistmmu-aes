`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HDqvMlSNSInMe8M2YZ6ecIcb3bd4amxKo2N8efvPyH/5uVUigrjfJAdGZCxI9sc8
bhCGd8jYodbbt6DVTb7YCOpNVKd4JnCMGB7dV/MwdaBNOW1PH48939vYOxHVhCHh
z0UjoRZtXkxd7elp3eaqAjeSr963Lo5KJ++TOYrUUoeh6na1XoSze0YaEeCcFlZf
WPsnBrDufYJ5eYeU5XdU/Rq/hvll+BShcCAWEXljVk86GOQ1gdNAdCZ5XwNjGBJM
sgo+Z11bxNoViuqyx/hjnnzSgIb8SiKON39/201rRsdxA3H/QV3XwzXW+VLVGF+m
Tw8OMTb7oGtZO/26zUZad2MbgPf9ShTDyaoWOfWjjjlPaSWBIFP6XTLWst170iis
2CAjoMG8O4OThy1ruwo0GjBij4kHs/Sf9ckSpqZMP04=
`protect END_PROTECTED
