`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u9TrR7FMSRUjzs6T9u6DsZ9KrzOi2gXTTwrzQ55A9TmfMlJ4+3aX7+xjs0ZUfN9j
X8blstRhSWfsptC57TpsGhE3mPUK4Q9Cl2IbZgThtPit4QzwXx5bVyy1hAqUP8pd
bUC9F0XAbmUPOQQdBqsbPaTgPK8CCPkiWChB3XQeJi2tvr+lwnCKs2kjuyvHEpZ0
wRUvuyho7u6GgEFbo2VQdtAYWrL3xKL7Qdrda8KXKCwEUg2p+oWMcbIFZanQg+Gg
3notQx6aVxXfjCD5aagv8w7NGoZZE+VSwF3lga9n+NV6wzhTMzBbJD8o1KAEYxrU
QUy1HozzGxxAk0zYGKbBhoEnQHR4pQYEesDOInrg+g/4zUMP0fpnX8J7qD8tvb5U
ThEix+G+yTanX6ciCwonzqD0+Ia86Bz7OQmuRh31Hxhyc80KtFRL4y+lq9pPNROs
gingoR2bGXl/aQM2E74E+sWrIVjwHSnFCU6Mp4fnrC909u/36sM5wFXPT3koYr7B
T2YCXdWjnUYt8jkrCJAo39jqvZB3k2ZJiMkl5U+qLX/Fayf1NMdfAuf1t04Kp2kV
lKiFWNie2ltWbN8CmHIwrKBUDpVXZqFucbBdrulQHRByoGC/rvHadbHIC3vgUF3G
U52hW6yz50dH1WZNgv5/ZJucunl1c7atO/gEAP2W7wE=
`protect END_PROTECTED
