`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
280QDvsddJe6yuEs1phhJQ9VqtWjKHOmacltqj2+YOnWVYBfgcNUBd8vtVykH6Un
eCUhxAUtcpKqSc+kHBPr/FHF+J1sQgfT3jlQ29LLuJZdsxZELGsjlVES1zON6t5a
EjlMzmJFRSlGW3j3mDdTIwQC6njnj/fXHJnbTdR3XGMRvsmAf+XsGFzdilRCC5Ol
NRyJ3LGntPa6Jyc60PW0fdyUjuycsf+MMgwXRrKooPrqNRkFfoguQhFm4s2Xgmic
e2ucNAxk+wf4Hp8JTPUqmHan/VkwD9C/qSudLzwcWweQkeeG/GY33Rc+mUSZp4gs
2QBwYmR0yxVMQvHgU33q2atyObsKMeL1e4A2u+UF09wXNc/1hAkh/BQ9zl0tQFqL
N4GR9eyYEd3B1jexVNGGcfzv4Ucq4DAilM4iuynI7a6XvISWnf4aElwRPPIr78d7
eEtExRbHQzqgXtLWUGNjc6xO+KB6f3lPA91dfuTRip7g+XGqaFBotTTxsSvfiYjf
en+X74JCicARqZgpKMRB29DKbctGR2np1FW3qZJOsLBkjwxCgCGGIf0QLTrpzn6e
xecRkQWk7fKY3yGuvnUdU15YxqfZbATNlhet5ESwhGopKRq8Dibh56fUww/i6pKQ
nwrbAWL0iGjuuT/EVzdyRhcUvSKu62EoPzjLmx83SNR1i/AE7f6ahcHomNqZJUmW
r82CIEbQPidTYZdtIyK0iKoCQc1u1et4E/nOtV9q1r5LTR3unNIv7uk0G87tgtib
vd/B2RDq1qKTQvf+h2XJMQ==
`protect END_PROTECTED
