`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IBI2W4fUclUwlpxNcjjc85nfTcpMrbVy1y6xGwt92EqzcmFs6Oi7qPn+8E/AtKdv
LVXIJUPS599qsK4Hx7S8BgcTvAJtuKvYz/wzYnxyz/MW+nGZlIQ0saYnOcgsziHC
3PTEJilTxNN1ZFCDRfscMr29YzU6IAtWbMIYHaXzx7utDmbLgGNt/Q5sQv+ssqzJ
VYHz+6O7jGUKA567DP/rJ1Ob+UsbxHEjShMNQuDmpvehAtEE8qEtdp7o5wzJW2Re
N84oWY95Zzc8nDEkILRmWfzZ/hx7A7qkYANTwGryV1oAe8kwJ+8UfAZDIAeHTJbu
QLesEjR3LsM4MIz4xsEfXUGBy69Bjn2uuP0Nxm29QTOErZNeCa9aT1/9LXoHG9bf
sTxYpvCrTCs3ZRXFrtx9iuqM9nEw5K4RaDP8QfYdl9c=
`protect END_PROTECTED
