`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xIOlBPCVBxa+Mz98fLzHolbGIgw8n06sccpsPrmYrHXowd41L3Bcqve7Jfc6SIQE
tx9zodq4JekAycc+FXNv6XtanB1VcMjEQZp4zW6YYLvtG6HFUTTtZ46faDpK+bbP
D+PmEUwVQS01tFo6hNl+CPaxOoVESAt+f4jtX+l3Rr4jHG+CyFHpARWEc+LhRTrv
d9AwCxziWDoIKYqhxDWiWMeY5VijSu4sYaN792oIrWt8cA+gDFZGD33VDYRHOI27
dbBjStfQ/n4PqOne0roGty7dNhu4mrNiyn3XFYR785QDJIlimzK1FdgL4HPh4Pbh
`protect END_PROTECTED
