`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QEJLHIDiOgfU3hTIAVhKPvgbR6MVJIdUZY/0n+9HHQMsuKFWyNvjrwNIgP8u7Qp8
u6GL7qVqyFlQNXjyTKhJCjAUDfdjgTfK/TjrV09psNAJPVPE41IQMv6o728qfQw6
Dfm9EkbFqE7YxYqjp3q8AEmVgly+i80P5O8tDP9hJcsOe+1VrUgqbj97f02gSuSF
3ew7B70M4F8ybuXT9WfjzvR0ioKtnG5dt/LAzhz/YYIBWK4pAUc3+0ZvP/I5kBhq
by5R4NNAnymGN5SjBLmb4HLbmNgV1Ka8xfjJUZRXtQ5PjcmmwqEYZpl+WMzoyWB7
GvRDazrfM1RMx0RZ+MrgzrsCq2p6Bv6Fvjzfm949dRV8nGzKuu3sY0Nr2B9Qym5H
hKp7l1YVwjGXbZrZizX1zgMNIr0u+HvXo52be06fBnZld4/iCC/iu72zMXGf8R4Z
nDfz7vsOHUlelOMR1D/ao3sV/t5EQjUVN0qasxTFUUtG2qvEy/pA2GGlSPJ/8jVZ
bKfZkttm1i4OuwlcbxuxGKi9eRAfDPEji+69VfCDZTt58XOJih8KtsWMUqpPL3Pw
kcOSOyTug8cr698YUkamkgDc5hgxOQuhcNs01wo0yWNqC0hbvQbjK5w+xAdIU6xo
cuFDI8BW/jMfmEjiEwiJqw==
`protect END_PROTECTED
