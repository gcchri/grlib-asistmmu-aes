`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ZDtM5iYV3vC4SFbdQhs9k8iQiwqzc34a9Hl0M1QHPk+j5BlLxawHnwUf4eS8PpL
zeKF79yyj36rn572Jrgsj11hf4xFcQc7YqXUFPprV26nzTHP9nJIPOvgNwSDhnMo
qo3qHKGHcjXFB7EZgb8DaddaeLmv1hpVkEkHryp/ne2OcP68dSwYHHxON4YgRadL
dkhsNBLD2SDs5mhMRihwk21pQ8rJiVaYJMsMtm0abXEcEDW46OffEqJLUfpOfSGP
mA0xxlMtaxXm+sjf56kbEBfAaHolHDcjVrkHPBgVB5kKOC9SuNHPaqBHY7S7ijXC
kIJOISV7kGPfxDqyixyVSaFOi3ij9AwtuLRxU0hFwlfUQcCBFEFVJwSQ21JaflGX
ymD54UQQxtW0OpUlA2FRCfl5vjRHFpEe++iIEkvYUw6AjBTgMghCWxlADZEyNYOr
`protect END_PROTECTED
