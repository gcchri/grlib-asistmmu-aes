`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CeZvrS2zYJnSafisb+uliP5O9gGNx/5Y5wVMKVdze1s4OObwDQiJmoVbbNcv4HuR
W7OPswojxIbVzMQpkxOw2+TH0GksysIp/GzLibb4lxpyoaHXuRvSL9qnmBsJzjbX
Ir7K7Ec5MkoCJTdNoYakJbSouj1NBj6/I877qpJ4SQUFXoAXS/PtYotp35lUsnOL
5kgMtojsQJRIHGmp8Di55qv/Dx3KSza6MJwa82ckkeMXO2wsATXamj/zub3bpgF9
zFfrExbFLIyzbQXZA6vWIA3h5EgzeOh/iqMKQXgOIedVkR02SO28pdHJvDWjW9B7
QFoNlN36pmcdIQ78LnwSObniwca3oE6Wgs0IFCUb6kyFBja0LHL7IqN8Y0ni+j6m
JdR6q1zReJv0HQkSOwrdMRnS+jpHHIW3E0EGzSlhWNlQZhnTZ5RID8N1vsIU2tZG
kPS3DPgrLib0pQEXihVBZ4r0YdkuT/WESB6GNcfaVhLmowTJWRDAnza5WHVdOCtB
b0baEv4HdYrTMdTG0j27SQ==
`protect END_PROTECTED
