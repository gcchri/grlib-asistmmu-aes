`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SYbIsNLW/122RUaI2Mhys+lCs2EPArnk0tCQXkhmWycyJIedezQe3yQQ+SCq2+jY
wjcGpB1W4xIsBYFSbINycQFVguWNYlmevAgbzJ6cXo7qtzpLuWO5mDipT7kgTGZX
jQUVvINU6ZErivS/M9j7CMm6NlFr9/1GbcVyHVwhnqIIgFWezG7+uXmiaMoH+gPP
ykz9tJbU6PZJQ3HAKJuKKx+kKdANBGTwIxHHp6l+T2VieyFbyW7plrdU4RHzwZTA
bvpsOfL6nXD9hb+zNLxy01XHqHDwYma6B8RqHj+0mCfYplpBk0gmcFywxfvET1z/
lAC5Eu2TAgXu/bwk93E/y6Eyrel1NjF/xPXi509DTqRjSmemVDe2mGnLONCiMTU2
5g03OqQ1NjJNko+mSgY9xiHoQDrNT1E8fZvKvDUZTP2VwXXFFQsU+qXsNsvOvYhc
UBjBH+S02lD41omZw4yRwSkwGnsZqcvN1ixPA3MkIgjzgx/bEbl4gsx888cURySR
3g2g+Gikut9bUjz5SFcD3zjeSF1O6q9HBuXELQP4MfHHxFYJIYuobT/xE4OjgOoS
B+PvhgqlgDQje0hlZ6+sGQMKrkVm7fZ0vS53Vh7nfznvhee77j0ESJC4GzpODdW9
Eel4qBVQWJCopDHpjlL6OuvTtHWY6erCGlPw8C0oGyiln45BL0HrCQ1VlYH5LPMW
LJ9NrA3jZzgAzplJy6mqm1G31HA2DcfCyQuccWBFBAEjjOohd0E/wgl95RG/F/84
KtI/gb0JMwGucIJzwXbWlwVBd3TrtBgKTE8JQbrPWW7DEXTgFEpUEo+r5WEQUrk9
oFn6zTurnKozFcNj6RnHybT3nHQYrrQmRH3RCFQdYYa9BcCX8ADdKOUEJ4sFj423
BDUKUw7QMleA5UbYc+3AxzXn1zCwZnNFjzTBmiyw1SjoyPehXIdHHLkTdPz+0T7u
vgpvY4aM+36YMh7uyv8f8gswc3bdGdMMqJEJk8h6Fb6piB9Jd7B4w7pdab2K/586
hOi1nMsrwCHpb45wz2L7RlU9fVY/ReOZ1ONpupRFZCh/IEs03e14DyYOhTblQlPe
k+rZ1Le4OXnsIhpR03zAsNCC8KbM3DJ7VmNCiyYidV+sL6I4av0EyKgtRb78WWug
X88kHiCjHPXGLcjQWiQGwiVjDYLIfRhLHWVTlCjR5+c=
`protect END_PROTECTED
