`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D6TuM1GKCGbQSNvB1NIGO1rQYJdNV+Snb8IK9MJQoC9b70oOfJV2XgaW0Je13F44
4200bDm3Hp/aggYRkNi7UP8R3xBPHjwmYAVOKbb8MCASpK072fdhyL5ya+q0Io5C
tL6M2tB4lER6Xo9w5i7gAprAka+4WlfMLQ95rsuWGVXz1gpExMLcCTZ89G2XL5gt
ycK726Ko4HeTKlxMRFWeaur5wIdHN8+dibHeUbdCKpBpsmlA3WAwhpzTpPaOInqr
s9e9DvJErgHmBGBa9XL4FDLwLiS1reuTytQstOFKZqDjIOFFr17qn85CGHKJFBm6
zY9QbFCJ5gK+/zyo2l+gVHgTj39j05hCOJT66LEy/rDqCXOvbZGJuVkVc1R5BoMm
0AKCGeeVkVIdZBkuYbcNLmtpAmIm3L5HymXk/6dhflyrK7r8I6xmZIiLymxdpKuL
QmWfVVDVeqPy/sUIYDA4pTkz3aQcxeIYwLPzmuWHEUIYSAU2A1FAH52N3tNmRVPu
Nk6GDCnMKPhjG4oWfXDJNGouJL3Ib4LDUN3BXzePPY14LDWUfB+bKxZy3LirsSK4
yXVpO1o9nFvRZ58DyBAEDWyKkCL3FgvVSF8IBuNy7UjTTDzHi6s7LSTJyBSqDTOJ
3ww69FPJ685uG7RSiBvIBPjTKmmM8JmtOWCsLwoOd10lKYp3DZWxfqHAb0L3HrHQ
5agb7du40B7p4FBOVUPsqER5depnM9d6SukfqvzAnPtqZCV3HkOYH0o+DD4F64yy
fLsfQm0oLdIqTaRxbl926kcep4l64uJX7hjYKw+JpwQCRME5vOrOlIIAL9ubvEvM
Qqg5PbYpEnjKCgR8O28m97Dt3hMhC9pnCXNDuGSU5FQ1vZxufqsbzJWswrfTZa7x
4nmzMUfLNUkjy3UfQhh7Izysp+iN3tUzptzu93S7V6kzAET6ogKay9wbmNhp7KQY
`protect END_PROTECTED
