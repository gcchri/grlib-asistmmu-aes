`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BE7NePR12xtRXERyNwzV7I+fKgHYiyC4NZ7emA7x7iW/1xsbxEjYW8+AoCS4mwPh
biGe7HEGfwa+BlSPyrb2XpGJ1XaX4J9w1cwQZjnz7o9KmoQ5p3l/P1lEkTus2p8p
fQ/mNPl3JQo8eChO8naBDaVSh00gwol96FW3IKNo2nB3swenHQZegnHoE1rQo9dg
fJpdEYXMUVPC3jpBOXWND4bCLXsOSkmav0hnzBC8A37paRmn1ahXj89TcZSAvHBZ
oDlEcNwxyv0Ekbi/8F8BbT319CbRmtHqT+1pepiilx26RGxHh6YBx1Pu3J3E9nDK
8xBGudjEXT4YfQVcao/e88TVrkM/Hnp3BEUKx1mvc3eniFdTkTA6r2g7eHdX/sKP
dHQbiQGZm/eEgdv0SHdQi0cAuoqnMMPak2Zn/xDppui7OuQjbKe1waQAPUu2Axp6
8G9B85v0YddPq7j7RYEt7q2eqH3TeBVB46PY87rLg4T3jOyFULMv7dN0AxN3ETnI
grTf9jV65BU4IO84T3vBg1BdG8a8x50L2VvXt3UvZDJl26KrIfWp47woCPG1DXli
7Tw+8EgVd5tMLPwPbGfijklPjsJsroGBtjLCZprO/3Bmgd1PV/juyzcs1bzLJk54
FVT5ySbPNG4nIYUbr/4qJA==
`protect END_PROTECTED
