`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8lOMP/6FGpcemcTkcn7PRfoSQx+6qxFSMe4goC//tYsQDWKirjYBst4Yx/FgYUR1
90YEtRVZABo7bGyOQJtkXE2VNIdYPtgNM4dXTsdT5AZsklPnjKgwmafDpCTISbDL
ZhzYgcVXP9Y9K5DSd9BeqEmNmjd2ihqVYXOMt34MR9W6tKOpgFvX8RURCvRCq0kd
RZRtGCZZUWqMGJWsqJILG8qcoT2EOiXfl2Xk0K5Z6Aq5Vndi5vFa8alzcrLAIp+8
2zGmqYVi3p+iFieg9zlaKiTgdVT62/QjWG/pzmaI6ZU4XhZso3VMndo2Qoq/DFYN
jw+qAz2OUHWmh7RHJIm8iQ5L0Fz2+tz0/pnvquJ8oIE=
`protect END_PROTECTED
