`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+adl11Ocyb6DEycrum07PGnmsecPeCn3ls5QtrcZBwvjpFcLYbzViKplkK2ukh+N
6SvqU6+SurVHYdJgtDR3J/cEml6ojngT9+mHD5cgkc/OEi8uNzw0nHCOAa5PYXMl
Y3EGwhA8RFgLSIYbIdFHVhhXr3BhZAZTznNMyWTmCXhDNa8RhEFK1KM7723WE0MA
Up+7ONUzyiC2y7YZuDL29rzBJ0RZJuA0cuW6BlVrdnJZ6kjjLXI/eCwJRQUw1+2K
GrLYk5v43anQv90yrq5MDPfm7hT2r4CG3C5+17AJg+PP0bCxRiu0OsJJOlIqLtCU
3No8zS6K8RTOZdfrJPwEzAtDoZ1+NQrdChMKoDbcXn/2AtqW8+iqkLaPhvvEdLiI
lkg0To6wuqSizBQJO2equg/mUG9QKObB99K2dWpuCcbzbC45K+M1qCbKz+Fp3x2z
ht3YZJgnxOMltAgfoSaWGwCJ1kTtrPIQJLtZgvkFTiGzsWrpr4aFt5+Yo7BSOL9X
3NeIwDLsHFHbr2YzTU8NykTzcAq9R9RtSpP/Q9abFc/ukIxP/nTiE5/H6Ux9k51Y
yYCksoyruJT32ohqRS4nfJZnvdg9scQ9JGlEatlDvH5cv5X3kQZyTWv6DCUGdXSX
2Zs/Wb4j/jBEaVVeiBdsXQ==
`protect END_PROTECTED
