`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rafKLlEJreMLlsQDbnReLoFLog51rpVxywNVtEzfB1myMO9nZsXM299rV0g6rP/q
8ql/gHOxeUJoLSVWCFfi4TLW3XO1GOmM6NnCSquN5aPfpm7XoWTjfzwoF/OuGmBE
a44ge8huUrmKFij01/OK1cPxTqvwH9rob77cuay/Yo8kSykn5bLcNCm8ZnZqesUF
zER839/jlaB7hxeSNKBwvpUrsSTnF//BK2flblxIalph8VyQ5ax+z0Yn00aCTq6X
TNigIqOFOJWnvHrPkR8gbcx9hnI5rWqdupYfTPkEBwcK4nuKwrhWanCdQX/35rAr
`protect END_PROTECTED
