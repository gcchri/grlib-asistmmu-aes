`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E9DngPvhW3+xjZv5s9Bv+P5WAYD/gIC/tcDShAW2Jwm7t6RTuHXODqvhRLmjlqg6
5udUVoevE9rLnqaaQ/ANSvP+annvq0oe6ptdRsTBtdnU0EqpKu8NoWUVVyqUwxgM
TtBgIMrVykHuvymmRe03uD2tbehVxh1T2DHGZJdz4OfYq/DYfJTegq8tuk5NuJFN
g4mULaG0FkROvy7OG1bDUv4isehuMgNg1ewekBeTa4cxGNnUWqo57Yko7Pcr1DIU
qjMD3CVQQWRku7+BjW68JnTgmoQME405kkG/MBpgdd6ilrA6VagihyFx+y2yqKnt
EZQlIATqA6hKVA8HodO52Nn37mg6G1t+whneg5o8DgEXnXo51YPL8V/byfP/TjuK
`protect END_PROTECTED
