`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1CxVnsy1UCf7y9J35MsQr0d8QTctP+/8RH3Zn8ZkJG6oRKR9TtzaTMrjNpqWoXqL
UzUHRujtCxnYJ4Di59T2Me4uo0sOpShPsUlVGDdoYDDrVLbcGOJStKqNTNs4YIDy
FIJD39Ybr9zVDbRL+XD4+kDBty5k0iNN7jHtzZKo2yYLr0Kt55ngHrw4UMObH9IP
dZIXZ2B6nuexJRslUr8iEnruksMEXRRy8vrhHBEPa9Vp45xJo7X6I+liiK2lie10
gVW2x/TAu6R6yNL8Fziczew+dXhmTaZpPLH9P+6NrdpeqSc/MJ6JbXVZhDYOl7c3
bc0TK7eNcUthzWUlUBfvTN+zvtTBFkZ/y3pptcwVG7EUZxW4dR1Xo5d5Bdl84034
f7wxNMy0EKi2mgrJkX/SQuKJJXa9VrH9CnUjGtD5NlchyUVLV9DDKHSCgl8ZLoP1
He/Nts53xtnWS6Nv+VB29CX2G6Vmf/zh+y/KVKS1WXPKAz0QyzhNSiDS9g9Icl91
19TGGNUspQNRJmkO603jhlqvx9MlkMpAGIXdBeEUwkJc4A66psWblPNgBglrsAEp
jmd0RZbiI1soYsbvJjmf+8JUq2OWf4LoMA2oRPBYKe69ThHxQo1WC4kDIOa4HJIj
K9Hj+LoQqUbjTbIwIxLogwumeMlzb3yZMgMRWgZLKYWF5fZoeWY9dtwBjT15BFPh
mSADC5R+NPSSSqbHtHT/t1jThgdHvdBcLpDwi0Myxds0H0bego2FvlAbOiTp2Wsj
QqobLcWp741h/aSdj4HbXRy89a5YOeHK708xyPjJzpJDQX520be/f77cBIEebFFb
LVJtdT2PDIIgHMFlq0GxUNGfHTDxyyPWWz7E2eSMIwioeidC1wQVSN2d7xI9x5Wm
NV86/uRAwxd04kABMzDLbDpGjZOEAUj2JIw4/kO0G9FjIog+E0zv66NfEGUWbvMb
p/1qBme3iglzA1GGu+TJNwXruNQ+nBPKQk/37V3JxNc=
`protect END_PROTECTED
