`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tpv6ttWD0I5mou3ynCqkRX71LmtYdS//Y04MwUBSX/C0JKIWRdU6/EK6StWGdT4Q
5GhMZHbJr/bU+SYr7xLf+17+qa4+8fF0bhj8MWnhGJvKIGTr+EnR2+nzVmZn+dBP
f4aqiofHfwk2Bf+gi8RvtUBPNWNxHuRB0gHrKRh4K7jQW53xK2EH/hqPgoajrVfZ
L5R+6q5hyH6BLykD6S9/vYw82ynmlfx6T8O3QPRlUw6yVPfMpeWIYAFZ9Cb7sb5d
JUCQXBeCRoo6AVJTqww87nlDkKX8NPCg4rCufw7JOp6rxH9ktuM/m/WX+7g/FGBS
lMrrk4NsYVmwR8dAv6sdG11rnKJ8+7t+p/he804onhM=
`protect END_PROTECTED
