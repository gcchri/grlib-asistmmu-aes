`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Riu12ptMCT8BrFXwQBOUD2cLn1iWBE3Bk1thHoYC6fPIFw1dt3oRbD+I7H6/qO0z
oSdDdevNi4jqkR0u8JhVzGx80fJZl004Gh5TqxGRo0ptcJdi28U8Wzf+jLmlskNA
OM1LSccIxxSXRfIIYwZsR1EBHIY1zXRg9yg6dwTaB5D8Xsm4h3ESNzHXeZVCtkX+
ZTW1o7n9NUTmR/nzTsSrYlfTiEBmC/c/qu0v8OpvcpoWP/Jx1VjWJaUK5KWcdcX3
4XgIxMqk3O4O0oLUW+f+z7XdIODjHhfSz7ZHhML//2A=
`protect END_PROTECTED
