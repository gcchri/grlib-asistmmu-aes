`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hwiVMABGYT2sFtxni2IfxcC0lGIIipF3Jg6eRwI0utHVe85puUbHP7Fmy/NNIw5y
91ZZ0Pm9mOm+Qp5gWwliUSAkXBDhzV7z3236zO2qZTwbdrre9gSZX4LNVKzsYjHr
Yqo6iGeaVoye38rp3ItEYYb48HVes+hysPD7fyMUc93ZGpd8XKPHFL6q+ET7VBBn
4BfipBq1SQKhGr/G5yiifJSQIqOrNuzynHvqNcN04pxXogSiGJkZxufSNSh6BzSx
heYtmHrUlTy1Kxcu5xTYzqyADk+bPjyyi7blwI+A8bUUSQ4K5BDEGPeg0oioekGH
o19wz51jwVeeDrzE/+AM+DEhHxx5i/LHKsJcT1/KXu/CwMogOWadkqAnFDjTV7Rf
0wllmWawksLHzkYG2jyA3+O66w4lrzgcxGmuZ8BeqK/AGLW34NxGQKngH1HIgCYn
guV90f3dlS8FtMl+36BbwS6hMsR2lxTqOz6ZvwZZPRI=
`protect END_PROTECTED
