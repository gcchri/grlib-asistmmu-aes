`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3zejRfAdyWMDCz5mQLOU9jx7PWo0sfDNDtb/tS9WBBVOxD4vNwIr4Ws7ZbS+wQdf
wFxznDxLQ80QgSEC24yYQkCE0dObgKrRys4b3alGaU6BO4r/f36oe5Xam3RauG7y
lpl1oeVOBuFUlp0c3Xf9CyqktLoaJQ9GKPewdNwvBcfJY3drMTehewXJO2xcAgCF
7TbqZOcMvnIJ3XMHLBf/wOiqp2p6PHyWl0bLdyKtZi3wvW0a0jbRozD5Jag6q+iP
EAFzYDBAeOJnYyivv/aXFDweqE2qcrAI+AWwFIkutZh+OTNn9ANyJ/Qc/pTQJP+V
KPjq2z1UnXfY1mNxejnoQx18C12qr0jU5VgBcRk27eVznSdb5jTMRQXpEVHTokLR
5DkZbqQghZreGtRlTBITOW/Ugv3Q1uUqnG8FlQKcBT2bQtZrft9y/IQ5aAQ79x6R
+CmlEImf4rtu5bNxKHItxGGiGrCakIBWE/9Mt5Pqie2v9JAJV+QsTnYJGFqbPDl7
EFTK4p3t37HyjJ3LZX/y1444zFwYVV6hK60mu4pM/un5EvL8g9BWrdkkWhnTs3NO
UmOnlvUKcIYeIQH2JtwPOuAnGKEi0MpMtUAa0etmtjivwNgkGE0jp4/d7G0ZtY4Q
2YsEcL9uOiE6jWv1lU9loev7Y7IXWyo/aHlVZnyzE9zmIMeLSez8cZYtNolnsSZw
wZBk0e/bVSgzetpGrmAY9nTgZnd/sxAqW0Wlf9SPwyy9FzAsZ0RCbZiHmesIH1Yu
U/GfGalRU59P5uepeOJKNT0gfkp97mIyG0W7AZVZdZVFq5vgi3wn0jX763xxN2lP
skIkyYu9RANlRMFp3VM4MJefpusW+kMRQbLH4JYuI8ws9d5d4c9hAVHF3JHaFJPn
p5DlgMWnekA1YLbR+RB+EQ==
`protect END_PROTECTED
