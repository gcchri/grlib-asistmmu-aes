`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k4s1ZSajDuKzahzv3H2s0LbgQxh9rQ6Fumq20DSeea09cjmcyik6cfwULiMThbcX
iw8GccQl7YQdFnrk81P1j0PscnaAcWyf4crh79XvhV6Lc1YhwkUHee6HCNypDoEp
ikDIXJIdYK2+FWTlG65eTiY+489AzSF0z4cB3ft8J54OmLecUVRLlFMhAq8YVPvy
3TBgVYSq2jhUcq8+GSWG7ijSFEO1FJNiT8QTGoBSeyXr7H1+Hbi0dzx8FY5I3Djt
Kvz23Uqj7jDHaS+sLut3/XaJfuuX2dJCPe76+2UdrX2hjdmcjOxpUugCx7+hKhK7
oJhpwtIH2O7htp8dCPZda9ETXDBusdkbfZz7cnxTXOwrUNWuZ8FeacN/K5h8G91C
6Qmx2pDEmwpU17usSmNb6LNM+txIg8byQBYKlHNxWaxWYLz6K/WFDPw0KQDds+6g
`protect END_PROTECTED
