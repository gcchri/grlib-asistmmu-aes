`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tNfihaaLxVz4/UMYDe9bsViiRacJB8xvSwgqsfLfInTJE2i8zI9I8ny7hU45g3cj
lk+Xqa1Mw36yiHNo6poNxO7jFFwCmV8srubNugN7cMr3sJmT7AVjPcDBHkPRdSlY
N6N1e+b0D7ZFBEqJjhrjxW5Me+GswuFG9qizy38QzC2JhT1FGGvfOvcAAoeZ6AK3
3OtGAaDhV7XMekZv1vAcKKQ+j1c4cz4rGa3Uh5Ca8dHQimcTu1f6ylGi2kA4W9D+
aYdeip6ho4YJpyP+6YGyhfA4eAYXCU0lHAiQ5uyq+eeCf2SjY+LFAf1l1RThdAh0
+HuniqfGUpw7HT7JgEzdjwXTVGHylRlwIvUr2+tvDDdj9bKstk3qHsxjSD04iB3H
0IDlOWeRJCPjtocx6G9yXABhZJpoLMiJDOzhANV/AhgIO5zAdMywCsOoD9tn9YEH
3EqVMizkithptTBDG+oJHawJBlaoTzxVnUJ74s4qnaM=
`protect END_PROTECTED
