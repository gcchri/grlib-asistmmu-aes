`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yHBVlLfflIB+apFi2qZreVmEb37GPzEHldpmsfgr8T7IttawBOJM/TDC26mZN8lW
rMczNwZOZUzuvD4gDWEJj+d9iY9SM/8jf4vJLee1HZxJN4VGvBXIYt6CFUvovVCl
aCsKJLMkCkCFdqvMc8YINNJnDteKSfIRq4UQZOGSs2UvoNQeFzqFK4Kt4+DSSHBT
IDVgxUBGRQMh9AicLj+k2fcHb+KJD4ZogVKEaB/fXUVSL8Td/gqcdX3TaZ6vonQl
GQGzOv011TdklSnHGcVIg5iOvalBHuLW0alAfmajc/TnTyDq1Hy7ThbI0ahaNa0p
wD+WQ+7YW1gC8NMH1GIZDg+npNs5EIcxkTeXemrgoXrymdwIJhR6pwxcqbe+bwxg
qtj976iqEdRLV7zurikYk8lpC6rnL4XlShPOtN+uy9HAq9uBR5F4v6pafI1+LgI1
`protect END_PROTECTED
