`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jmv4QlolvSlVasOWJkqLzfqptJ6klGJlJ7XHFmfDwiUoAsBQziZg1g8jhVekC1Ah
VmGt/QNOA+0qQsiJ00Cy2o7KrAF19Zhifxlf3Wlb9vmtMPEoRlj0QX3tJxpv0UEp
ny6Lw4XqS8hOBcyyutbs1p7jFMu1QufKI3/Vl0qy8m9iKRUbENI6IQQfD7gbtT+s
WAPYh6ZJncO282pjBRRx+X9UzZK93YCq4nw0e9l+CGeAApVeq24Uu3MY53FH7cO/
Po9Uz3uJN9mpV65D54DmXA==
`protect END_PROTECTED
