`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AJiIc0L+5fweGkmOjNqNFbX5lcG+7GMamfvB7LZXszGK8IHFNwCba+H5yDqh2qwb
fCE0rcJPd5AzocyL4dmY+ErIiDr4OPA7v1/5s1QXODPa1ryD4cUoW/OXwfzmVEAa
OV/h0s4EPkJrW64XZrhFUoLOxsOvTDl5PqiTqU8ivY+C4xexnYOkb8JQcz+kzyf8
JTLQC3o33AJHARuctkGK2LHN3qeOxI9BB4Fro1EHaHpUpP2hryNH3HL0ks+yf4GL
KBQcrN2T/D7eLaLt6CIW7bWUK7E1wieD5mlBsoObwlQDXnE2aM8tDQl4V6ErBo1g
CAdHQcAycL2JLOy2UXR4yokEdctR5Ch6WoaAN+NuUOb56eA1YCgIE2QAPFYHEXmt
Vh0RmgG2yfq2nkEwQo14DrwI19cCOGuid0C8mTxudH9q2xKs2vcQB0LvCGme0KqE
z2W4iMQ4fG7JRSXq5+Upu35D/YSb3qSeBH9g591uZQ9XevqdDQbui+pUnXhLjLZP
`protect END_PROTECTED
