`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
efpX+0jyXQTuI87Xr1roo1ZAMAFL4uDNnpm/x8hTAyRsPtKIzX/6wrVu+PWQLIz/
Dk7FsoOeclr6QJNjfloHzl3nu+haguPRJ0Xc6B3SPlHAhq6JYlaaNc82A6BymKHz
AnAGMmVNR0npJOv3rf2uln+1YmNqmcU7KqHkMbRa+ME33wm52DVPhTnXLRZ2rZMf
Ed5Xlzy7z2DCvodvHBgMBshnhC128mqBSdHGQndhyeSFjdxcNeVDNfyZuiVP3dcq
ZAoBIkosf2Q8YyiAbmifLxib364WoaKasR+vQ3jAJcE5x9uUr+3XqO+jPmCAa6jl
okNb+VUFAV84uOZBrWXEbRhlhl2DrspN6KkcbE1dd1fbx+foLFHu/824+meFBM+w
/wlAKGK6pZqhkhVepW/8uDSD2RV4WLd/qZtp/PPpkBVqEWW2WNKVyif7bYZd+5lQ
KrJqgdZcq94/I9NfIeT+BIq1agXdw18Ih3rcIXCyzcdwo6WUUbbef1c1DdApUlS0
0FSNzOIXDttBEMCQFkOkR3C3h7dYRre6W1TKw126CbA=
`protect END_PROTECTED
