`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
opdcZ0wZggb4o87JY+rCKQAQb/+hqm99qwSNnncu6WCdH8uPCteyu08zJxixP7Zf
8k/GUH4nDM0vrqgXuhs+kgrbnFHypT0JxPpkpWws4xFlRrsY+gfFHa9a2PH8Deun
53Tkw5eELAAUInPFfGhlsYuL8uuI0p2qfwhA/qse6Cf0KhGuiz4983svZtCmZblg
5ZMUZGeqBAK0sd6zzIs/91ZozdVpVK7z6FlIkjlQon1QPE0JTioSGnqn08YHVf78
4j1VvEvV8XJDfi5DgW48ZP2gBa1OTAvTk3vFojH8r/qH/TFjPWuikkEb1/nX9bkO
TbH9Zt2rTYSasggiK84daA==
`protect END_PROTECTED
