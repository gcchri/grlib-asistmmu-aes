`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hzmmu5hU2/eXXDtF7hKj/nydY5/s7F9KK/44hA2XKRCEBPMMCp2Xlam6wYybd1/5
pR4atjmYCXbdbFSAqlTxOJzwvSAAUqaQi8JfUvovs+BLzvKKXW0Zei2hQTpTshNg
GY6wV9ezJCWnjdIjzcWIza4ApQeBjTGnWWT0xjuOKWjzZ2tA1gRMGMS+tTlVyZR4
C/j5l7hAY+5ZlMVITCq+R0Yqwzjd7tPnpEVaf+FRx/aMKtQwssvGSA95Pf2KhY6D
/QxkSAdk4Oc/xtyXP1d0r/uVFHzyUGmzvZVqfYltOs6BkeZwcdjcYyGjyMQq4JQF
5DkcR2pE98cTqd/xmEMdMUYdVV1vCRHMho53xx/soJ2q9OC39tJV8Sg7sriwTXrX
JIX96xqR2klX5HXnmdtr8TC9D+QN8J3wBlddVjRNrThOmOH/FM14KbVyiW5e9O1J
pYLqCAvYDa7hAgXSJyAjv/LlWKU/JVmMN5TdaE5rQkZJvI6tqI368D5pW7K0EJ8k
ZryWrCIpJ5SNW/TjonGz/OzPcGmKIaLs35MLHNsEZHD5yvIV+tfKieUwtAtKFCP/
hnEYDUKhsM7jW1pE8Yofbkbk4Oj8amQEGCJQfW0qRb9WcwRMb+WjsOwXw0qU1WhF
DytVds1UvxI0F09KvqEZZKJVJikJec3Kar9RxzRvBTR3UpKQFj4U/a6GaNCnUt0v
0kDUas8pldJQmTOw7Kp3hJMOmmKkpFz+K6bXmOt8PhWg2h6omhuJDPtntOI/xuae
Kl3frBQ/H7LQQZvrA0LTGOPt480uogc13HwutNHRuelGnYbCBxrMZXQgiyPiNhFG
lQ1h/GcGU+vTbrdjCQRaLRxS35TXD+mhm4/EkcEUN3Giexx6OyER3kz9a+kHj7gU
5zlBaWL8dk0bV7+YLUdOk8Pm5ixTOmcnJoCLRSaW3AmJQaNgl744YurCtJp157t+
fqpgsom6txMPhpV7teGy6coNcuL5P7deb346NV9eOu6x3nXFoPAp/LkU3prjTglP
DhutiuZjeU1fDczA+v4bCQp8OWyNLzYwbb163bo1Rg9ipaxo02KQofQz89628g9z
IlhH4T3tPiAfitJtsG6HPBB+1uIDDW+JzDeUY7gF3Hk=
`protect END_PROTECTED
