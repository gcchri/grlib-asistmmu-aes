`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+5wkLVh+mGcGg5/0gHU/CESgQtllUznxrRyHKZOGH68XQyt9Po+YbdBnJvxi+Kct
2yuWz5mYUniybl85tx47qvV3JrJO6KTxLaGGAS4nl/SWDO2f3+HwfKESC01gpfvb
F74ytoMBgMxN7XHeUxXFnaasmND2YdqkwdyvodUh1dSghpQ09ImfKK2yJBmilOpR
twiei7j36Vq+0x0f/siQgaPtOQKUFwK5KcnucG122Mzd9d8M6Q3Rt07I0Fu3FAYe
yRvchM0l3elaWfmJ+JfrF5XotY2PMWf7riCGRElfZ4wp/+8lB1t/ccFDTlnBGiod
1Ic3Hb2D5lswAEmwrVolYCjA3xdebb/2xfqwuLSUOL0UCDtRMucNvp7/020CtZLG
m0y5WKkrAfk3RXATF6/ZFp4XVnWn4mnH3u6yLMcjMI7KWIPNyV3tTW0HbS/i5ea2
mSVGX1mIu8KyNaKWO6YMCBgirmaGPMOGzOPDB/+Ov1/YugKVLGgvuT6cFSYBI3S0
5tw1Ki/vlQ8BUpeY83rOXB2t+1x86agSPHJe3c6krthLaJoA1SQDJQ4IjcFh1Aix
XP8C5FEFqfhTU3Kv+cJg8LNA+Lgt+T6S0ChnvicD+2qMxNeoMZxwHHIaA0h0gaus
9NIsE6jOWPLf3QgRmNtzTIpfeZNU4GG5u1sPuedjGKRqKNFTKx/EDUTOqxBK5D0f
JAASYw8HlUzy1BW5qghs0trCiI4MFM2oCn1NvOSSW+6/48HpFwGK0JK3FtHvTlDG
JH5Wa/lLd8uUPKLAVzUzUQ==
`protect END_PROTECTED
