`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RvRoWvFqhF22X6MRGfkSm+H437+1W/+k0PB1fxLoNcRH9Bh/bp0xwbMoLHoaU1jh
29itUk7TYWYko01wtygbnX5771PBU9U/tqXz6mVaXqbYTytWSh8hFk6IETXlCvM6
oLDzrCxG4HYJ21zCThvZEBa9FE+X/gJW3CToU/2ezbfshOZEqidJm+DlBLxECmsv
3/RFydsFvFsan2S30pAvH5ql6a0QKrSpxLdP8tOyxrs3kABCVffq2w2U1lAUPDVC
0dKJBlJA1iRZS9NZWVoYVmRXr/EOSGycmrXfvY2eiCc3udn8U4cBVbE8m6iQIStJ
7qARcoN9dy6lYmJXyO7aUvvqemHwgYgRh3UC+4LmXgxNP7ClyFokKz87KzGkO6do
1nnyKGeHOl6pkrV5vxNyGIkPty6S8PERsEB6n4ab2DCR224gGLkmIEcnKFGZbhGQ
`protect END_PROTECTED
