`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cZOb1y1emcrQATRVQj63ICHdZCPY1OXMjR0UZfF0Rji3unPonYBzYD2vnWrbktta
eKHVUjbiqHWj1R4dQ8W+gqw89SzV1jYVrHSItrmgF+qdH0uwntQ3uceiLNBT0VtN
0qU4N7VcicMCrVX62/nF/jwv2JsyP3e525GJAmoEUZwON7yZKYlrM4qxIhUpqTwB
AH1kaLPrmgs567zPtIQgM0RbxUyg8lJPNuLe5ReEZdugb1oglLjfhGRjyjOkPoPN
auC7YZVS4x6UQNWOxMOmbXPE7ngCSKbbHCKv7cP7E41wuQSasVOGNvNYAzv77BO2
csJkLAd7s7Y50dTbiemN9fzHRKtI8iVvvF4Svz2z9Ht5iAxHqVYHHM7zkIduo+Se
ZJA1ZJrqmze/0u9dSzdc/g==
`protect END_PROTECTED
