`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CMw6kNNWxpcRtYyQxp0yLf2bGhGDRwaMPgyDSE+2QVFT1BUMZyuyH0Fd7+KaA/zD
2eFRbadVyeDt7kefJGU+9sLtCYfO0fsRkQ/L6Kh9oMYm1IBzLsAguSfizukfvup0
N1lNsotE8FMp8axUmGEf1MdTrSYAbV4JImNyTKTyPgyHinlo+WGdtjFXyw34nTeY
eGbQ14oc1ky9L/RqwOBJI/n+m+JYNyLBkf1a3Hg6TzQhQHfJSxGaSNFz3gqcizKc
0hZJ/JmYhEfP4+UVBVQKziV9KQPuxI6OfDvqdz0jfLEdqFOb0dCAvZKvRsiUJOrN
fkgBnMS51498/LJJLKP12FICL4LrT0tk2aIdaUl3bdjt6vI2NQJO36LMYxFeKEX+
LOky+cBsX0Iqae3WpoXET/6MNxQjblm/5fTX8PhcIvkp9kqTgZXExOSq9creH+Jv
MIuf0hT5agBI5yNK9IsBDmhUX64NJTvQRVnU94oWTM9EbXWPPK8fHNIPFRJNdkhg
aeMaEh1uh6wBhc6BvnPtTemg+luSxPMRYrJhxP+A3mlRW4dy4HCDH41aUi35ScP0
zBshq9QMi2JWGcS2fYXmnbd2FO4b1pEMPK13BAUrU2fiqAcSu98S3r5iNyMUXGeD
`protect END_PROTECTED
