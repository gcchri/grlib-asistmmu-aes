`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
19xGsiHXgd5TlZiSqiYqJvB9oA1vvObL69c97FdMgQFDGGM/Z5d3doPQA25ptB95
hZSt/KkDAvSF+VcsER7uIDBAH0JvW1JcA6jYtBhL8ExqVtauzNAL+pHA46OtAqfS
n7c2WaNO6YsQxRP1VF/3homFmJHdgPUM8c5Ajw8rYBKtqR7LRgC6fPEYayC+57eg
NqoQp4efm9eoE55LPZryGl4Fldentwyt8O7VRf8boNeo36hGqhnH4UnWGv3TxJNL
Kvqd4GqwvS1SRE7HKpcvW6YK2/UfmVKlzFXpE7bFr79K8MwsJ6xb61IKrVjKhnAC
LTM/3Ob9tMhdV2DpWemooR8JgMgaGTksvcAXHrv+eZ6aGirjCLIxhV0AwGDnd6h7
MQ7XWb5Qr97MXIoVp/MCX7t4U28gnzYvBTJLuY5JryZZHLD/boZK6wGuW9Gm0GEK
Gz6NF/MT8FUb1hZ1obwSRjHWRYARvREbdutgDirJMcJSqIQkbTrIk1NGS1XFV18c
5+xQ4tBLRnCqqfI4wMs0G6NrUDLIFyiexnRPY/WY6G8PxiGcO9LYjLsTKJ2FodnQ
AjhI1pzlqxor0dl1ZSCNCHjZngDOW9+L9tqa9NIvDHnWtdhjrq6f5KiaV8jUXesQ
q59D0S92TqKbYTOWFOiC+ZvdBWGHOweoQBr0v8DuLAM15dYZT9jS+FSy7+8cl+A0
/b8fbE4cQtfx/Jhfja4hWz4yYhiVfCRaXa9/nU7so6LvWVTpD4Si52w6ofVc21se
nbt4LuHWL+fKetAfekEOeZ5OeXCK6Z8qx3EPYlgZ3vTMfs6pNPovXUq8abK3wuTt
b0lbvylj3f04jdq7EPCy7bDEy5cEbbKaKKR5/5DnOJzhN6f5mtAlkBrDdVBOI+Pl
KrWG2Y3YaocYu01QlITYIkqvWI9+hLbEBrvR+OifTpKQqLQat0ntS3wIpVjAqzzh
ilK+BUJh/Ng2OkhQl9aVONiPYj4tLSld9Mm7YbHFpLrCcIXIaK/98T8UbTJQzyMA
xD/HUNTxdltyj1RCO57A+39KtrAbJUDS+vT+baJxCLjl7aJgXHlys94UQQhJypEP
0TLNzVPWCCw4hHQJNpPsbugkBvCywco9ize3SyJ5zmLp7Pt5hiNMcba715Z5P/Wd
00X7t2qxxyzpqnY2Bbw1FauPFXMTsg6hfK/WFBUwGNI=
`protect END_PROTECTED
