`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yJ3cTyDiOuoRAFlOsEjb3wNhyLi0+u3AApbfYpGEqWvjvEi5lR8oNvzTt+JRWmsi
CrcmdIt+4foaPdTrAiNT2ym2Z75KysvQS/3g8Q08CmRPLF5GBh5NO5263ioRIQka
bRTFZ4/4mNQerREIcqqQ25JsNiNjjsGZawQYziCzu3ktWttaJ71tDXm89ErGXqLO
h0inRdrqoeejzE+NXSzAQDiEuK+f0Qchy3wONP3Sbzzd5usyyc5Sv/FMrpp9VF8P
OmO8aj1etlK5nCaFu+XOY+CW/yN3j+2tOvKXI2LZwtBTQy4wgmyTxncVU1EeYJy5
8odG5G4gCqt/jI55/3EytdXl8KU9PNFCMiZx6YXe/H5exfGFIgF7OMzOuIrtk2kj
3zZsbUoHTYXQrpgW/7nD6GgANXMTySzTksIcZF7GoHjaFDDHHXeMioXA2LCXzFVk
TA1UutgfTpwRAYEjxxPnLoSawr2Vbv/+YpZXBXLF936zQ2/TTDqBhX9zkqs+/q2f
9HMFdpECYivXMDY5DssZ434hPA3qN32mok9Fv0N76Ck1ug2sQFyLezR+bn0uio8z
ImAmgTaMSHQ0nt+GDcdpIg==
`protect END_PROTECTED
