`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
54LRM+gqanEUbhSgLanGzKWnpm4Gv1saaGbl/RrGp5w7Pb3ntESvwxNG2cRCiD1i
lYtFi3EIa53Efs3ntwy0yJ2RH3WAdch6SgPfkV2R63XDgHr/wbEwcMau4OfbYA79
I5FqV0sj50Jrx48zSAl8xSWamh4iWnUks3omaweBhUeciDFUKM/RbyWxfgND8j5H
h6oz/H7NjaMvO97Amin+AnUl7/ProLaAycGRb72+pZ8+ECqvF9eWDYuGOfk/YoCU
TK67ofBdJ8H2l9GPGWSPh7esm29PZjfH5v174QGEed4fZPBPBnSCPfXF064bIMe/
dHnNQm4PVyzDGmqkpQtM+Ll9J8ce4VHhqoGYWGq/q7vE82NrSTG7bBBvHjLcOGC/
1ROYAKU2pXa1jXB6897hijWoQbv4GxcdiQNdilDXyBEdKmCm8it492enrbtSOULx
N1l8Qz1CFczDSkLhFm/cPnwWHWBwW3a1dTS4Yt3bwfQ1yWXXzqq2wsGFxnl18+sw
`protect END_PROTECTED
