`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TC1wG9AViIykZbanOtY+AOi2Nu+y5HZ3subeZuB91Q4genMu4yPPRFI+FLBF++3S
+G+PKbhgyGQPTlUh5Gcu+vwzNi1OfXk6jI67ULYaNXztHy8SArsjBFmtiiUYNr4T
7DcItlMhiy6qlAXQDoz61AHXQ+/dl7grKjkR3cCpQtdY7dtjsuU+xs7eHaSsDAhQ
A5UwVW9rx7iGDr+tmnIODzwyG4qAXqGxwINmmHpHHaXb0wkLCWJm3ADPzg01oJQC
i1Jk97NjfOFA+ENWG/PAboAvpJgabX51PBNRM4/L+TJuc0u9F/oy/b3geEAlkJYo
TdMjYBNRZAyvc/eYkrna+X9T4lxPckoQSuwQbGz8/1vgKXb/NQrzJywxqyy4qpVd
KTrd5gzdQGdYoBcDnT1Ukl3mJwPX5u0ivzwziVaC4Ta779CeVvDCpxZw7Q6FdHb/
Q7O1oFwAjPWgr/fEs3phMHDc/agZPTbl/K6MVBgl3PdKvv9sn7p4u3jCDOvSESfk
4S/ddxVCbshwpe1G9tPbgBZgsSlCYqnbaZu6BJiw7Ao4Y06+0j21t2jpnb0V+i/C
krRRpkmxTVDhLV11ZstjdiqZAl1Y8BCJkpbQGGgHJHpKvmP8zMP4AAlcBUzAHFLm
8NdDcKLO/IX6BZdDLwYJZRbwfh4RBKo+j5SlUJjI/s77XuxVW4UwMxvajtgraSBH
dwwmPt3nD456+Lsk/qhiS7cwIyqRzGrIjyCkJeRhgByHJCo4HJ/dKPxWAcJraSaH
7Zbt7tqJXuFjT2AsOpXp5lHp4JilyjIG0Nd/uzeuwUCvu0wp85PkYCtuEahSxpVV
Gk3OWoqBs7owjwT9i1iYl5WQzeKQUi3YORLIvMZIZOK+LTx74bN8sOg9D+4k1Gqo
UNWK4BMNtaPl1Ld0O+toQsBYlvmgWpiDEXWv3AXzr2nVEPK1+eGooh96fstLVS8j
CMImXfEKc7xoTC0fXDADurAZJ7uShH/r8pFkm+xNa926DICT0qEkxyGkj12DDiqy
QeTAH8AFbDYaCGH1QE7oA8DztcRum+RsWxIWca4aAUcyxaDqzdAITatFGOs1Qfrk
0s8hgboVRUle1Qnh1s4NErcqFnRufpBQbImZIGlXV6TWmzPIUdhdPXT9CKdRHnaO
EVixVIznrUgeBC9Bw5SqXVJdK95ExBDsAy7ueWwrKm22rPw9rZSz7/Gg5AMhCn0F
IUOOUHDdkQOn4WqH1FoNn+ZLzkTC9aSJh9SL+JKkeiRnT612/EKy7y6aeK9tuaK7
/iBuqgsnn+yhEEyrm+vR9aP5n57BnzNtetUfJHuSvhbJaPS92yjhvmIAKy2Ym1Hx
EbrZbInz2+XkG5u8ufDgodgYGmlwQXhO7AhtxEzmcq+WE6BNZuRuIYoAQ/2jH4yV
`protect END_PROTECTED
