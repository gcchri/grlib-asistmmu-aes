`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/AeTmAkxLLiJUAeGQnmju2eWfoK4xEO8YRncJSLcWc3ba/2rFcGzrqt0mUwuKSyx
VCfGcdZfvghO/TUs9YyJTx2oE6a4jg29FqoCpobUHAgLIMODMl0FVrSY3BGBaxPN
tlJMcx1Fl09T2LgsOPm3A0bDWvTyYrh479lwn5QUtATI0UWyk2SbQSO952SzecmB
kYMmjlDRDtKeo3TXiunLi2Jx7XSHevXGGdlCWeYBFYh3xPLHa1A9Vpn9JTLidIqc
lkcDOmW3sw/YqK56fiijJbVUQFp2gc1irMkvsytISVxs7JayaI5evyBvgYA6Dkge
y2WBbjPJQk7afYA3NlGHGSS+xW68/Fh0W8stHGoOp0obPKA2u8WqwN1LMr0tVYBy
An8n9ySJSu33zexRj7mqS7/nly5E8SaNO2RUS03vQc8kYhIiPc3Zx9korhhtN2dc
+ehgncAMU7rnmE3LhOxRWWtIwZ3+sE6CR3/GFz5//by1dHLyHaiey6AG1RvJ/On9
j2ULvHhPheMU1VaaU5KLW5nmaUOc6GMwI/3bRGkLOjEFMd46BNmLZ1WGiv+EUXLX
d5VHi2i0WkenUc0ClPheKVWPsdr6MgHBuGA1MSdQ1FRULrJYji3DHQhH5yy75qhc
2FNvPuw8w6Ii4Fb9pqAkKFQ16DD2cj+IyDcZGIp2xtD/93YcKdv5VeYGPF9+hKRa
GbpVfmdLBtvOSvIEC5j9oLnvV54/1CIt5Xb3204jtE8mx4r49C/KzQh0EwLpgL2r
fX+BM3M+wudsl5l0yZaXsagXW6fS8oOoJ+LY780/Nte67B9eOT5gdJkz+FaKG4eM
/YTvJcPYNlHwWa+ttnSFpdyvDG9U7lkTaT82tIIDdP65ZbdHypcfqWz6QiB6apSy
bfmIb4vxO9fYi8gL5JvJinh5rJtsu6AzjE2XNSf/FLbxLykSXZsDqcADxSsagMu6
fHzZ3EMSL1kFPmn2f3CIlipkrAZ/8pbo+IvA35RJpwRfCa87skMU7CEg3e+6LCk+
FGW4bTPIP2rhzbET12ivxQ==
`protect END_PROTECTED
