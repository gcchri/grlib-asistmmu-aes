`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VAZjbee/8nROwBrZrnxLxRDh1npRmuckIhNfSW1S2bhcWs1HhdZd1dQQM77Pnyza
m27c6A2Y0VlEEhlGHgstvdybsE1TLQUzGyE77eAKPxYJ4Ev34ZQyDUYgAzGIQy2D
mbp88kndh2SbW0FP6G7ZgoMeOiQw5ZiBtXzdnr0pk8bdPRfXBdiaF51Z4gujsiRM
YsNmrvagFv8VPt+5dEPoHnMvS4baqy5kD+ljM2snbTVDavi+X5dMIFTzTGx9WyZz
UhxWLNr2NKxwoIgOWTJ+MnXqZgnKDzJz70kodjT6bkFv8Frjat6OBlp9NPK/YXDK
O8U2mBNoGT5sHRg0hAE2WzGkehcELnCXj1ACMuAebmyf4VwpMPj5f6NgwpH0Zr3X
AuOU2ARYlNqAQ99ENX5mGRIuUV0H7v+kJYcEPDCEOvfoH3hEyEuh57wFbTWB10gA
OpX1q3RbRz508xNK0b/9rJEA2X0IMq0LLtMfJmcYmywUDaf6vEq7Gzf4zl/+Zh1Q
NRY1J98HRaYdWj2A1nrBvVwYjoWyPlchjaAUxA7o+cMjn3vaqDtYZmpTdHFCd3V+
UToDxOV6isZtGuWHIEEuBGRaXc3jDJKpzhk/1f59umSZ7gPozmnFfyWUjejEyEwe
NLAUIC/GvI9Isbdg05MtoEuFFY//8NvQvN8L78ocrEm7xv5E7OxMghu/k73/mBZi
FzYadYIfcnWN8CjoV9NrBINS2t3rxdsmc5BNc5uL9WCvRT47fiCbPnRhsWIJYRhA
`protect END_PROTECTED
