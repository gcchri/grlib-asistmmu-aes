`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VPl5wSTGDQdQ//KVkQK84gVhkcaZNTwtfQrVXDg5Chm7g4vgyalCNOGyxbb4ZPWN
0gjStxh/xvvjvoY01fo1Ter//08OQ8HpbhFYbLMHktxPgxfIXjTM60Zuf8mS8B1v
NX/YZJGM9b50KHRrKcSWCeDzw0nNF8iSMkWpcAf3LDwUKVL46i0ajmVuWz2zHrKn
iEINNo4+K/U235V01vMs8encUmGew7XzBxYTO/cGPjG3fO6DsNrcd43BwqcvIEPZ
fsuZ0lQ3b/s3V2U13WIP5+hZKeWJYGGsgWos1cKr88l3hLKzxhhA2Q10+U5/pEZA
S/AN5NfaxHH/SvdS4b24wYtn/fMNaSUgUcUFmLZ2MonG0MjSBJwSSsBMDq2yUUM3
gUTzy/E89rWfR+yIrJ26wiAQ+VKp2OJpEhxkrOUB33piHiqAWAufEdBbtg0ggvH5
i3iFLRUNpegWF6bQMjDIwVB/o/7Fx5YBTjSF1wNp8q0ZfkzM/T619CeLZOZYcAEH
76qIVmLgauT72vfJBglUsV06BgMdQOh31pYZTSAuHWFgLShpbsJNiqGy+NuyMObn
gPyIkZHYAMxQ95u7XtE1MDw4GIDvHLVc00fHGbH53hJz+Iqk6LgjgoZKGjLnm9fX
rbwvPElvZdNCTUaNByXQwWJSSQsRW9V/b7OaMBORHr9TNbKgzA3qofUWwlQYWBQD
pUICHMMwpKWyyGoikF8hndfSV7xUG3/1ed6NEWC09HtUyE32MNi9VE64cC4z/UHQ
VbTg3+gUnVt5IaSmn3p8ajVm+n9+LnAA0lZZMxzapv+iRjLoE2AW9PiiToLwxcMN
1Oq2rrcC/M77os5aRq3Paui2nPEO9Rs+87Jm1w2cP6EgzojpWeO5nd4UQbn4pq7k
jUiTlhKHc0XDwnSMJ1xiHPuMojAMsdEoQLn26s0DKVP8Q12vWBfMiG21Qc7UDjQg
WULxJ1h4PABGKsXav5PX489Zwake4lp0qMhODUJYbJ7XFM6+xbrsjqvePZeL8mGy
fuYso4uwOEkImw/sR0iNuPBxnkVoz2McRSiK/CMOLFWRwTvbMf4sKPIkRVwU2du+
xsWqBYgxwsnKaXpS4Uw3xHS3fp+Cr8OkuBU6CjIFz26yS3b9g7LwNzoct5pmp1Mt
cEA34O4n/Cx72ZVfQMALfxNPNDChBPkPkajxLV0e+WdlZrkGVlZYfSuofstEfGTC
5yticL7rhqMYT1q9ShUCwME1Mqed0i3PWnZAasSBM5/1vmlaHWpjeJZX2rpDwcuH
M4burMGBFkvygz8O9V2+FDA1NlFivCLhOJF4vzZiAOwWnSqqLnpoAwF7ok7Iw5vW
0WeczjDT5K5tg8ORsDxeL3Ij+ZU7oa3kHbChHHu6ItX0v2W1MgM4BC7xY3WCZqLY
eDoTyBgqF67Xzrk7rBz9C7qKJzrEEAeHeXz87bA9kWTjkIck/IuTWgvYDf0sjU6b
2Txu1JEli3fu18v6fcNhhShKS8d8/J1j6CPbykxnkphEeqD6G7Qu0QJFJOqtwcr+
kmK9Va9LTtbE9oF8+2vySmqCEnnPCtqPar8MDyqRJ3gSCusfnsomah+UZJVzkivE
0jUcSlMACsRgYjOvpnpgy5lzzc5WVm5XfSzzl1E8DPuF8JtPZarR92f40unEJSX1
ZWJVoE98qsATtgrHXOFbhf7HjrAnHCF8bGOrpJkyIyGaiIT8sfEa89/82LTCf413
oL6bMBKzON8gnRr7sdCZMKIKXEThfv2ZJlRGwtNg0QLFKm93Uc98rzoKajpfLqeQ
4HHu12aRnRtfsVFvaSuYYztEQtrLLCQHTrOYWmTdnWzCRs+brj4jPWG4FVUWr2Mv
2dbFKV1lQaWpTxK4yfKSLD+Gf4gzjk9YUH3Kv4O1eWo0FR+aUv8mW94/RhjltxXj
mIViVgTJ2hC9j6cDWPWjkwG5AR2ZLRKMZ7offA3BmIYeI+5KFOYNN97iQ1c3zDXd
0PsnE91ZP6dVD3K1RPAMVcyk+qrRywrG0zu8sdNlAWQ6SKEZQrxiBVMPhrK5MdZQ
lYQ+wLOLtsdlfWMk4RgNA/XUsQb8HwAaAVeu+N989q5qmCfV5KsfA1QQOIHhO5Kr
9mMOfBBNSM7pp5ywcRu/ER1XMRLsmDiJrIn40Md3oBCK4G/o0RyDKA2H2pbhp5gO
kCtgIFUxLqqw8rRVLVfBumXvNgAUI1lzOHte3qq9QhTK8JI7353aA44DXu6cPrQg
1ivo2ntplkZrt2CCD0Kyt/hqZdILJcKES5rVYvQykoRUI7K/hiitkgI5wEyg71rL
OfVRDzTz2Bye5zRdCy7Pjjvh6dVEc146wa+CGBzbef9FvmMQmAWTGSxk1SvQh/i2
s+l4bSNTrgYePEa6/lZbndRXWIdvxz5tLmSkncjit+3g4oZT8QKMMiqrIfEbKiek
JIA4CYzKN+PX40zMnN2dTBqmjGUu3EV2U+qiLvl+nOEINJk5YI/GeMrpyJGI/ubf
C5xMoSwIbuqrJ82NLWv1FMzavESpDV6LWnpWbDcbMcvzjUeu3Pc5NPkjzQM1HS9p
MiJyN6BO2hpAsoCrtn1aVLZXzb7HNqdSM4Fm4YzrZZuhGcETxjQ1RCSwFyEylQVB
Q6JCNjwOFCvg6jR3l31lUzQ8hWdV/ndr4BAe/hh8KKhn7unBngA4zt3vsFr8CyDw
db5jgean4AaPrJJjr4OFOZC/v8jExClbQrIM64evRZP4DO498iacH68oNO1UFGZq
wngNAOS4uPglg1uzJDgtgBgXYn93PMqGCy4a2AaWQz73IfHQg/plyguEbaHJozrI
t8x1VELJvs8GaH/atTsMsxqs7scEVWOo+iO4M1bldHHnPgeAQJagcUtsDjJVXwAz
V8Tu2e/Slgk4KOTrBZRya9od2kBG1oBwYSUVt2r+7GXWGukqiS70cHtUJOYKi+yn
+8l/IQhEHE6GaQqJrfSD7dZ99IBBCsAVGJDyLRI5OddXSCY2YsTIIIDH5E44d0wt
a6g0+h7BCHFpoD/czL8MPjCPg9+Wgb8lZ08MbU/k2z8MNimT0dCCKC+hsCMvNe4B
lZ1W4pH314G5tRaWKcwNExUeMxwTpDMNUCbUN+VyI6yNGRjo2tjdKi+n2zL9zFiP
119P/puuF8g+dxCiHGwit5uE/OE855TDppL/5hpaCc/L7tZAjJxyiL09eg1hy0pW
EYOX0W//LZFb8CnWWkOIFC/kGbJW85Jps5kBNRjQzByysgH0FdoM1FXZG/p6QB+u
v4ginTiNEYQNxJcPUuUyJmL+RMD3YSiidV7AIBecqoikalpm+KL0HJfFM7aLi8by
NWTRsM3wNb0AbnrvWhpGEeatK3GQCeBkYfaLhtSHxnpLCRjF4aQSpNECMvwF0Xf4
YyJlwKRVM+ddmfOXjwdZ2iRUJbgbxk8TvhzjmRTIah7vOGhg7echgHC0rCFFzvSd
F6+IEJuqLnqISIvJAgpeN5W8QRWtI0H8fyTSoVmwM+QlziW1PMoUhqRs9rQ3iV3y
7iEpuRhMX/LKGr5mu9hUtQvNN35Pu5hcyK+pyc8VEYe7vddG+VOdrIqIqA820g1p
/U5nb7PP5U1h9AeyPZfp3Yc/Im58zzvOwVwiPfkGzaKGSOB5igaQnYjhCSOBsVYg
xvc/VYu1s4IHyp/HIa2LudkGPyKn1LqtRhjNa4rigc2uqBVN6yo8mNmz/imey6XZ
Ps/dKdVGrXZouVzlO3IxQ3mlxfH38c2sr9ycHilu9z94bn82PEZX9lRKZDd9FSZ2
r0T8Cv7ITb3DKd6SUAU5ePENT0Y9n6pxtezzJplKvG0xcmPV6swiFe49yIC57HXW
HGVDfCGAAg6/bJ8m7CnDTSlP0qYIAcsiQptxzpgSRq/e/EfTy0S5BmWty6V0t5MX
GKYZiZPoYh0j9QfMNjdw0BCARRg87xoYjP2VOifmYUoAG/qg6ULvySMOcj/qV2Wr
NkeeWw+tEOR7HHmnZixCUfn/qYyL2m+pmodHE4zHFjXvk6S2PqwLM75NGcYJTKZO
Mmfg1Wf+rxFqVszlSJsdcUpOOtytxFzxYq7AoTp+304iaxIUbwEJFGH5B+nio50X
IF+CKTnfzaJ1nuyf2+olcZHtspsHJEya20kOs/KIEckIv/w4mRX63D7zfaVZGafU
uE8NqySL9cVaPVnuOoWuhaEiHJKNz/GpmrZYDhYFLQM3o9NPPKmzuhHG2rbPwt3O
f+FzgUMxfmtFOX3fgLf/rhcrWFHFsat47I9h87Yz2VsvfJyERqorFrU3nq4jtPur
VHOLofFhOh9HCQXpVbKRw/SJIRn7tPeUHMgTYrc7BCJQGypRVwuKd7Xi2GpJWVtA
H2BKM53QvSBfgEvq1N6pB3Wt2nXnaMLVJHu35E2p7KwYJ+6JFNLYzVWsPoEr/uAw
v6Ne9I/d1Fx8z6o17a/DY0pOgOIML8sEKUhoTvTTGaOw2bOn8nbGdHydhC8eklvT
j2+uQ/l5nj3V82GoIqjn8ofnDKAz21jeYBOArapCV2PUzfv/nl1JbpTkKm18051H
29RbUFUyOBNTCpoHc8GFv5Vl2uP3aRXWwfM1yFPu6HCFs8Ztqphx82W0BmWeXw5R
MItdgVtdtIKzM64LuO+bmqK2Md4H0DVo/cgeZNy9uCPjKIxg7XuCwByKrgorSRMn
vP6+3XUm+uprmFYnA6NvIyxZbx/mYU1qO08g0xnDEABvA9TkbZlqb/jwqi+adTGf
Pqh+WBtH2n6BYx98d81g07H259NOAsVmviefStRyFud3xFOj5H8AqM5zcMLWWG71
RqOq25yYuz0ToEghyxIh4+U8nir5pWjhmkflYx19XrEYRhVQfcWSmClzELTJJVHP
23drPE8Aq8r6HNPkvs6wieXnkj9nGXUZw0beyPrBaEB3uJchVTQnhNUQe+2hOasf
v6sKkOi07NL9q6nQrB/qWIHlgIbRf7Y02ESRLpx1cKusv1Dqz5JngTS1psbQbT1L
W972XTNofrFl1m7DG6ksGgZj/2T4BptMx8amgRzqHiSNdzPpW28WpLjTZ3ENR6ZP
gFwbWBjOGs5V8HE/xT5i7Y1xMXeGw0OwACwfzfG7piC6Csa5StziF5mMmMgh8ssZ
m0MTxwYEEAxU2Woho71ujgXp7TVbyRNY3QoFNR7Ly3qqorNdocwh6Rua2qstLfFv
b4dJQOnIrjzWuWsjW4BqnGJSbUtS52Puo6a7zlpUxVpe9xImfm1dqweq5GR/RQEm
Qcdslo8f+QyWlbnFKre7wyebyb/wQdV1TFbKFmNnO28wpVekrpK2aDG4b2UgdGGF
vT63ZAAZAcaQZjjjhh6Zk+Vcz0ZYNquRK4RroYo9C/1Oemblp+Dqa/aPeOr/w5Hx
czlLx8e/zqj42mXzOKpbw5bpAikKXv82mTPz98p8316+yCPGDaQBvqH55lza8dTW
V7qOEE71EG6FuRxxda3+ngachd1IJ2iqOl2fBiJCqXQkvhIUlh7k61CVSFqoK6HY
/Nd5ruCk4fUJP+eXUYYxpYIVP53C4WwCkeMTrjDf8wT7qa+9ieWQUPUr/tYGYJwW
qd5j56wCov5RN0aPgz4LVfAGk4PPSPZftNhGoFPKHJEOk8Dw9e9vU2WQs6JRKHPm
XKPe/LJ9yf43oukTAVpU8XkrmHDkDbHsC5i0i54cn2n411Tq4XIh/ZmmoyPba2Zb
bXrlwp85RoI2RH1hKTQVNxgfLYdTMEQpGjl+5vpyfocGpniZKZe+lgGRzYUy7NMr
hvodhx4OsQ68arHcwtWahxNsY+8rZp3glIrcs0ZqRqmogCegZtWIDAyH3ov0u1Xv
Jpt96EgR1quhbU8Tr+wsKRLhE9FF09HqsqIO2vKrRMjh/zK2IrMctSnNErO7u9lu
CxaOmMIpqIQHrP2aTGxB+McYSAGas0tOUk/A950PesHTPZhaCKvi9xXeh7ow79JX
tY4wxHaa/B3gUHGgmDGRaJBgHtgOmCN2FpfDZISVRuygBaqyujrFv8v9Z2VqoHGn
8H/7pyiubALcNVXIZMCUiWMWxwKetJjhKQc795t+R767hYsJKq2Bosh36FY4cD47
JftLDNfdzyRG76FIvg3dWHHKMmiormXXi228rd4gDsKo2/SvS20QoigU9nCkC7ja
zh93DUivyzXP777ndJ+mAp+ZtZP9VFYZC/0asIhhdN2RI3E5VV+qzhAfzSbwLTFy
K1HGEVD7HRoe3I/60+JDDPCTnDON81GWKDR0tvHv4mKLKzi6SvYErsR8HePORXpe
VdqFiB6tvUqQPKd16aNN+dGBNgbrnCkiPLiqVYbzedeGoMOBtHkwpT7oX+jnbZ8O
0OOxmEwxtc2lu8q6LySuY0soL/+76NK5Wo5wXrY9rWWI4/p0UN/W8tNsgvkI5+0W
7yEckbME7GgR9w9N9BNfw654GYdrvbHOw06DjW11PbKjo/ko9r9o+rWQqAr+kpKf
qtk5kia1bSOUcoxxRQJAM7aLJ24KJwtJwwD57h02dRxX5bsHFbiRdqtM4spXOuzH
STeKOneAwzuJSE7jsTEJ2E76IRMEjRaShsAkYd06zErf1nzP8BTGWGWpTPx6LFGS
T/SMhh91hXJYYXekqr9rlivL3EzOOCPuoHz1DfYaXMyYvlTTET6ETh8RCwQgHnwB
0Z4SDhOHNb9UldZXgw1aMIMaGTantofZju9g50fXhaEEaEIsAzvDTcspj7pIRyiw
r+4GClXYi3I+r9/Bzyc/r72Nxu24AfKSvdT1nvMPEq8t1u3P6rNm5+Ss6bzauqRy
INY+dvScgLdNw7u2SsegpHSC56gcxMM+cDOrvB/ixIWVJVTiPPRKwhgIm7RPDPHh
YtxPp4F3qfVeGVmXrBLndenuxGlu1NV/XPXU7uVHkL+W2XFgoCiGZj3DHK3f22w8
sepEe9efye2BcC9svgJ1jrF0H1/+DF4RP7VHY81QwE9y21gNSYVlRes16K0pznVn
QQWjsXxAPvl4AJkSosomXwhJURyK8KNEDkAnpFyQvvSpmLAXGi2m9BIDPWzTQrgW
70I4QFNatDarta2k6CrmXyyu+7kGMO1sNBIRmYMPHTjN9MGsMkyPCCEFjN/QC92b
ejq3LcW/EFqO38PJyls7chy7Y8KM8XsTLRQI9UZVdGeiyDJP9j5AeblZMchHH3OD
LVZYd0NldjoS3rE1aQ79b5/WRI8IhhBgB4zGU59shXj47QrVq8YMUfsN6fdQkh2q
iwWR+pUrW7TDwzRxUipNL8f+XtazTRAD0AcZMZ+OFW3DSXkR/RXUPcOy2mwATxCW
nHaqIjDoYgs2nXjBf0scTv2yqbKlbv+qm6qwey+ujnZ50LuQtuBD8Im65qRYAqq8
0e8QPwhn3IliciP5IZXD8nDT0qQ1qqxBuzQ4Z7AB/WD62h4Ef+HFtyv1kJkQZVMu
V2gup7E1KpZcRE9gPCDSiKyWHPxIjEflUtzCfvrEdZ5ikBDYq2/VJfSGuXlWHX4U
N4b0C/+hDoXz+UJswiSGIIdwuKmwB1qFJGi8UaRA6sNVo478Mok46wzZaGWIPYMf
ag86RN2yTjVVlCKk+4hJRJCioOBVjZts7xIIwk+3uD0eRXrbN/XZq54+A+VRxqiY
/kuT/rU+jDaH4hNuiYX1So+WZFbAwEfJthWN7F/Zp576u8o+lTI4lk9iiEZ44RZt
51rmDxc5csu3WqaEt+TFvuql8UDkTZYMSUWmV2tDXdQ4SvsQCrAUKJmgNW9gPwmQ
blJ4FMtXVze1Vjjlwl/crcbPb0GcwVPhRDi8VB/Bh0TILLdZg8yK9wYiqqk2Xgb4
uGP057NEQKirhwLtnWKu5UAJnnyd/55HbIJJBbvVVDHt/uY4pD+/r09D8w24U4Br
4+43AXNkiqxlUJr6q8qS5jiNskoCHcKGKDyDtPG9s6fU+2s8SXd/Lm79oRj0GTP8
cqGxpoxINo3T+I3tvfoHskPv1TrCi9FJDhmeRHNOHKxneQBCg2ftakvefLO7+F+x
V0RAJ+h0WaP22EGE9XRt8ohIeVEHqY19bOrzUXzlA1YQq8erGgI1aVf3epw4AKaS
GfDLSQGwADK5KKJe3m2RBv2Q3UUeBkEU/3oMUirVe4YFwbnEo+hbJVbozskHsQAj
p7lNs4yGVYWLxmogkUmcEAsuXay1UKDQlztwe/861emssNfqRTfpnfFWqcVzHwKC
vxQkhH60eptJka4BBU/45aACtN4uVbko8nQ8rPs35RYtqlXRITBIb3LL0lEGos8H
Gr8s/1bx1wYxocoqgRydq5+I2EZ+tlu0N675haanBswOkAAyqxAYeSAK1IKi2u0q
kKgA4yhz4yW8WVGEj50faCyaS34aHUHnAXwD1eBUr9u7ztxmCh+w8IKQavWF5uA0
L7xSRrA7bXEU7vGvT4M808PanuOGuXTPE3kkYTBhxhBck7bR+MOg1UzXvFq3eLGv
t97u3e2JXAmz0MP7uzkA5m+op4MSKi4OdO69duJ3kLmJshv4uQJcXbpYfAtN00MO
i2qy2KyPA1rpqt+Hcl+VrCzRfWHGGKWaQgsgXVhZKyUYkG/viyFtoElgmNhG7n/1
U2HpIl/uFtA4ue9LgN5laesgtc8tfMYuYkNexamrtMaIpRJPW7Bsv59Xc77Sn8ez
ZFtzq3WsF3PJdqSsTy8/Js3Q0xqjYbVVGmP3EFKnVZGC76uv1M/flx/q0VfzGnpK
m4tWS0gSwnLLXOBNhZtPIxL+8xVQqDuCymXnjAVRqtCuLpO1etAg7fGQLIc+1Ruh
pElaxKYo6kqIsTDahM3IrfjrxBzWGHCiN2f5xlHxOwM7oiuRs7Vwrt9+Ncaqbxri
3Zsx8beAEIT+2gD83O1nwiLSp6UqY8dUR9EA4HFO8W88qZQBS/TA9zNDJ//bycAT
gP3NbfJrkS5PR9/UUu2z5CUdn3MeWHEaBuZfY1JQ+22aiOCPXYSPGKoEc8bxr7zc
+FjDfCKk4LEFyH5lYZnvFfyeWn90V9CWRZrFoe9WHZcz45FZusNr0Uonf29T/DVP
F7hXrAydSMu4bFg/cuDDoFiwQNGjTeNTzanIK3+VEztf/wP7nkeD2Ksfc1NDibOZ
7ND33udNVkxIg44kbpVh+zS0QA/FrE48mIwm7Ge/4nvnXypLWljY5cX19UcGH/9n
TXYIP9A0PfpSXRB+0ROv/G903ehFLDHS/kk031RzkchJg1htDJRhFiNFQIR3g1sY
kiNGuLmqPxdbr+Zx2mheQCDZB0WBuhkLnkvrq4MGVZ2RwQ76ko/B47qfz5GvIDf1
EjgWKEUHkDpLTizKeCct4V6WhcKBfY+aV4hedPI7LdmEFlBvOD1PXECt0lqjQ50E
9KRgXQIYnJCOD+U43A3HJwR5C2fqvMqv+qSsXu7Ya+UinIf0sp/y6Fq0nHe7QtrY
cbexWvlijjJUsb7ZmHV6MaUv5/rgfSKdNi0cbj5DFZKpeWviNKXjJO6Mb/+gQeTx
MB4Y8vbhCmiWAsXfWorg2zN0WRUTRCgnTUy3twtFz/m6FeRXFiHPYlXm/UBxJBeh
oEkMK4mCn9WyrR1wLgOUnB6OUfcO17RKJn1xnKEr9pu8WETs+Adl0oy298tzPY7P
IxYioQmqD6YYyfHqZXycoYoKGK8XCk1967flFhtbP38MsqiR7iKzpFdzSZSOhgzn
DyVl1ERogLQyyOpL+ZABVxtslwOFWDA/+088A70EveUHyihegQrHoCOKpTX4PW+2
Yw2uF//nx68/79JPInpYZPnElqS6y8qyKqRLAEI4T6vfBFDGD5lpWXyEMY0Gdjgs
5FEUglVr6H7RUMoBSt3GiHU3B+fg7oGFofRKP5i1JORVun99UlhssdDQa7yydvLk
EKJHHTHibGfW6IKkHQBzvLM18vs1LUHXTsaIgjVBYEonLkIs5cy2RcvUG5nfaYXR
QqDfBKE2BQHzx0AhTmoUY8xQfF+/gkADH0K2P0acQHuZ4+HvJc3Q9M302MMYaQg8
n8GTDh9/YJ5sX/Nh6bAaRhIjk4vdg/Tyvzs4dQNXw3/gCPcQULj5zim/FlBFU86X
XDS+wLWOY8WIMn3O5l+FUePQ0cNDjCOZ06rWyPoGJOfQIVTQd+YRk5nlb3PGfzJb
z+Xq7yhDMCfDeVTXFGD8SQCXPEK+KJ+TVAwknvpROQPunO5SS7vERuHsRBq9GDCl
eJHpH4bMBYJB1YY8QuQdabUU3g3vKweyEUYrDCsk9NeIfc7lw3pU38DZJv2wyMTw
IW+5G533boFzmw+JikDgBHAaYGSIeW18pOHHSfOaHKgmBLK9zyjwrCHHWguW/uak
8LxxGC4VOct33D2ICGQpcynhYm7CpQbeu2QFbNdLy7Egzxlj29PexrjRST/z1MT/
JrQqvkR9Ji5/8G8BjTEJIu+6AZOmkkJxrevmt+aABfShrCdYWfZ7EZenrSJ2mR+L
ZE23x8XyvuwvTSlDw/+aENh4/xE4Fa9CYUM4N+P1BjfN9Csjw9eRLPwmsxn/nlHt
iKCLWmUCqj1fu76iNJLg1YeNUX2W4kmucb3v6ZmlPOncxquIxYvdCPz45JFo4UNd
SBXzROXsau4NlFi+Mm99UvPRdGjDR68laC4KSeU01PoixXsEiDjrNnbrREk+41Vu
LXrNyaXmJvjN2r1TB0qZjZBddMB30/5bxS1zQAUXUUzlN39QWnfBVxxXEvvGb9NC
j5zMJF5VrRyg9H9AuNlkY8Oc/n8dgHhzkPyJvoN7XbpSApXq7tGpcskLWUkPuy7I
G4C9fbL9KcPVO3TJCf+Q+hzDqDY25gbEd5lx4D+elxviDonIxkoM72FSt02W5oau
2LUeaSs+VTf8sX9nLHMUQJ0PNe4WQvu3Osmw9vNF6HHcJ6mDiuFOopT44X6SklKJ
2fFthN+UqjhKlHd10NHE3+9wlK0r4GqWupexsG7+CNQDXn5FSUP3ulew3E0Xy0ur
bWKF7lSzdlJzduBszAJkhbbicdUTzg30pJWn1UXB4mLuW1TiGKV7LqkBb8woT2dq
L4PBTlFcgCeEn5fLW4GtEoKOzyK2t2sfSfyMpbsElG1V6F90zHKJacqmIzg7GlD1
Tppi8TqPffHmPCIF+0zAL4WtliPGHeYU3wu+RoiR7S1/YNn8/gQ9DSR8WSwfgj6Y
3/VaKfWiuVcLXbo9e82q4AuTm0sdrwHOds5a1n8v0yTqpLMVNxQD8oCcZFCkBnS9
EIGY7zMuKfLNgVcp1u+McAvxRDKrPPdwtCUI8yqKABVzhav/3Fs9ZSpfQP+pvE5f
nq+FCTCK+6Zn/O4yfXF9XTtYXh1fGCk5xvhJxzzA+V42DTXxKBz+eAf5EEb+8Lhe
bTsbPbGV1pMEt1MuzfQ7OhwXBioy8ALMs2N9iI5rYlEe4WNfkGCthxwAjl4TrEzp
0sSy4VSC64AlzpFVtHviVY/ARLCubNSY8vqVwYDZkLVmeqRwt0euAGT7gBS03DH/
yUia/9lDuK6wxL9rGYj6ZjDeWnHwPuaf+HR0w/PscLwdCS3zx3UZNzfTMPuLRpv0
`protect END_PROTECTED
