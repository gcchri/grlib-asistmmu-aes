`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JMsA5V48h+FqWb273v8AsSIBiIz+V/2rRHFQuGNOF0mM9wMDXJ4rKMez58iUP8ua
5lnSTcBQ+SS8ptXwDiQp/tHSTDWt1FizK1S1CzbuTdankH7JnY3dY0E8yuw34Leo
twTUEWSnO2JHGn830iBE91K8hLFNA/lQUKNmOQgmhbzryGe56CjgD6/DdKZJhSfZ
oaYIJKxoK/o0IbHXMbca1A8Ot4XrMOuoI5Nt0X+eAhx05CL1aTuRzRlBQ5BhTrsl
85dPEZzzhv+1Fz0YtLU+pybV11ZXBd8OnmyXRfTcgg7tsmuAmGDw/w6IUCXniHD1
RR7qWVaTAL91WvyKf7ynordczw1OSIFayGrNA1LV3e2x97gTxYivHNDiTQa77Zh/
`protect END_PROTECTED
