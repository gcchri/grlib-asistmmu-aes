`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WL3W9ltZz1MEdR6T+YeDNcF/eu+kaLEDm130ztI7Cqvkd8OiMRdQFJuXqYWFmo1k
MKiX2C5Lck+r0EF4asjGPtV0sFYMk2FL6bx9Jm0EqAE25BPR0fG+IiVlMh/sRZIa
bdBO1y6R0fPJDvHnZ0ODOKji91KFo5ydUZiHOdYJhfOKwajncSkT6tKa8O6y+E52
PsaE+IA1V1I+hyqScBML2rdg7D+JcM0z26B9jhAvRQMcsjzrd3n2fIEgOmC1MSVK
/Pf0n+44W8Vj8r6kV+O1RTwirmHWE02WyHu3+WvHR43rFxKXAOGnRzKLwcrMgBpG
jZqFh1utS40k6/yy347/lvY4yZeL1m+sdFcK823qfSElE4B9Blbk2sRJqOzoCzk2
c0dvSn8CEWML6ppVs5P2P2tfZSGGi/CekjIrTKHQYLc=
`protect END_PROTECTED
