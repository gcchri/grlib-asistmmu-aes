`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HKWqxqe9PCmIpEgIFWskSCaocSjmc57LeGrZbs74k/QmE0qBU6K9N1G6d/IUVUsn
oJrUxbM3UScRslPEHC8qEuYywd0SDvjYSJHZL6KhedkJQtVg9AvPZjMNw7umt52r
gcnhBbegXB/SzonsFbxygyuCEs9sWzqUUtloHyoosXeaR6Jhfk6AxweVJDxaddwB
8XHK++T4wos7kBffAgtt/1w3/Wpq0TuxhPWdctGdIkHpEQupeSitI4/TiiklwPFt
9caNR5PVkaIZgWRH0QXBfiSkk5DxdL01qeVbYRLUi65lUePrnamyjMXrWF8Kmkyj
X5MOuFKHF7Rw1liR08nd/JHfky0/DLPMLtWrmvloNVr29lrDAzE9dVa2vjPE4MIS
/E3Pc/xeOjSZ8nKuEKV3b8yjs+0v2q33I5hgzlRhFa7DvBLD7T/i8Ebw7ZOOVBZn
OoWCe2mygl4bELU0ZrlMmW3FIowPWYNKqVckTVE+EKQ=
`protect END_PROTECTED
