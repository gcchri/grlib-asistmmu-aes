`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mS2Zz7NXpFE3MtuH7oaJKAnp5yL1a958uOHnxjpefsjKpC211jyxuKH/LedfYxjB
qb3JhVLKNNXc5M3GpLp9vX37LZLR+Wnt/4eeCdDKwHnm6vGi0WnoJT+rgZ1bXdQe
v51FExVQ5GtnVxCptPfMic8L1ZokF6c9UwYQ5flUSguVCIy21w/eZ2oWUQWDj4y9
knGCTJHJFE4ZipGBebHQraGnH6b1nF+p8KupcagtxY1HboJDJ4mTGP0jLlidA1vS
hjneQElMr5n2OYfXScVCsIYg1OI8PuRp67rPE+JVm8MHMWPNH/M5gci9cwGOIwnN
hWQ1MVLsHraBQdxyh5FilUUaDveowlZg2iHZ+x7MjpryYgPUceMriEw5v6V3v70Z
ZY+MHGMZ6yWfhTbjHINU24T0y5CfFc551Xe42dL1VjDrhH8AremHZbjO5DsSUS1x
`protect END_PROTECTED
