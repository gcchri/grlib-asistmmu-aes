`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uOW0gEdFvgpwDb2qrxUmHo3piVdwD+p31qDHvqvLLvgr+ePF+UEaYKCQALFmryEg
K5hfNl3Oa062lKq66z+rhBno1kb7do8zpkC4+MZZkh96o/2362hXz7sxNfcBS3uI
QAJHG7CReDWttAyB49Ktafq2oWui6Lg8YupXHNVFbo6EDDhXAKbTX0ZWzzkIG1sd
PTB7W8bpBXYwCjDQmMU6Qe274mgYukcYTJAlZrf4Oq/2cX7rLB+1UjAttd6j7Wpn
EqAu1Am/Bh7QVo7ZBdlzJnk9Q26pEhBQf3AOjFoX0HdCdBBAkPrOeOKCasJMQVuA
DM+x2QX0osGKtJ7nA81hKA==
`protect END_PROTECTED
