`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FD2LJri6U5fIRziHSsOyVYiFryc6n6Aqze9h2x8DoQLcsNfQnAJrvaQL4TPZCWI4
VKTVkP5OgMxl8KVE11g1PkvW4gSk7H4mA9lA3Z9shnGAi8/LHFpN58NOYW/OGwaH
uVnVK19l1mF9g6/Ms8Ti2WkZesz99jI8XMwECzpoXiTMTtZiiOX5PBAnw3BpoYns
Pu5xbEJRb0REQpmE8CjPLYvrmgTBAF1OZfPzID084dJ5zWb/KEX7/jXSDBhk9G/T
dU8eT5IT4O1S7Xc2sF/GZCdzUl+1p1N0HxCaBUBLecy3ed83x/lAR/bQS0CYwrbv
`protect END_PROTECTED
