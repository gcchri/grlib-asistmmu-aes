`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6T/wsJ4XozC8ywBQv7DhqTmU0zqe5DcEdq0/5ap1j/tSZsak4mYd8I0r3T1tQmPq
87TgoQUdFy5CQ6pzo7aNT2LUMQtqylIKuPfDAzgkSCcJgwFI7+YMIjKUuY9+VRoc
ynhfGE0B3TUleoyubQQWETKvg3eCi6NrCqZJUrdbYjwyhtqKQV3y/6NLQhD40YL2
VT9ojPoTuVf+BStDSQTMUuxu5pgEX56XkZ8RIdHrgctNgmO+2QSxBAo17dafZKde
1UE/T/dGznCTlAE0mgoZsWkUOu9Et31+aR8YvDsxuCdAktSsBc6cviOo05kpbrMG
AqeB+VsFV71VUhiuQ9UefwJaaWetbTEpG+1bJ6ct49H01HeDfRc/mS3qigv5mnaH
FsMjgoVjoKvWz1n/tpGgNtv/CWoFWml0z1GFNEmr+qnHO4/mrkX6pIiLjgqZbukm
07j9AQ8PJtL7q8QLEysHx1SxurPpvEBd0JeLy2f+0ktIKqOIYPewWjEd//wIqZby
/cLbR1QtLBAjeg7zzguUVgGvsb51tB1QIRQX8ub2nnhsRW9pfIdhLkhk8ONzdouL
MUfq3gt60Dnvh7xVASLS3w==
`protect END_PROTECTED
