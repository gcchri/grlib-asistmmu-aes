`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ktOdOeviznLuCYU9rnyQRd0rK5B0FLxjHuvStS39SBTpGqNgFpjLKGMugTa4oIp9
RpTmbJgLtwqWvTTGhITSLT7gogjxnVrp7I/i/eXhRJydxXogcR33nCk2fUp1svnX
pIeL2pk7sYisgiDX2wX748iOv+9+LTisPo4BkulsTvGNcF2AL3zkw5vcPlux4Nwx
iv9op9Mjaes9y+9rL0LJUz5tUL1JJD4Z84p/AsmHaaTfnjXydNPmI7ZZ2aaknc4L
SOU5W6hSqK+9T7zu+5aJw33pxi71ZAU1hqv47KdpvuiB3jC4fY4KO5oVT0WmHL27
MaEsU4EKRV3tJtZfqfLOOH1LA762umYH3EolF7fJrPPHIRR5sdlI9X0YQ/thZzyS
BYaMijtfEGmAMFug2GhjwycaTX5kichOhd9fOKnPiNw92xuVmOvIc9VDr1RcYBmg
Eg0MuIbG/Ao4GsYOO2yreYbKv0eMASHJyczuTudj8j7krp0fMeyR3Ti12KHsHRhp
N+mJhZmiCQpCUINpxEdU7/oN5/Ey+HcobNoeEouyGyzKWSL0Sgu32okBgbtmApAw
XOAP2TDfCO6LsYsSO87/eIPATlXqhAEr7eVU+zdlkGVqmV0+HAZ8L4P9vGbsbMBG
ThQ5geTgOhP2NyQPKQvNxLa2SABHX09yRWo7dRI9V1samMNbs1R+LUOKbwsE4c/x
7jPGTpxv2ONJq1jWy1y3heBbFa2hnNiAGRRv5CWQoNU=
`protect END_PROTECTED
