`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/zRYCCVWRShhNFp6bDi4/UbOeEEdCdsBHMJTAuA+7/eP3C6R8WVO4fEh38/mRi2+
TGq4EKC3CZfj7v/691Fcev5gB2eGDPTTmLtVOHRTt6kpvPx68tcdyAo4tCw6g/uk
DjXRtRy0gNCUlM0JTbo8s7fbA4qrl5S1YstN+X+qp8mKDyIJWYUK+Mrm44nPkK0q
RDzgZXSmfLJDEqJ2ZaiyRjdldnngCa5PAqQVOkTirAhAnYNrH+Ogae6Q0h0KrJ8m
SGkZ8pQPfy5URpIHVuKDeg==
`protect END_PROTECTED
