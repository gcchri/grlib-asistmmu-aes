`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
btSZ7tggKk1ZNQnT9JsvJzX2e1yP98Lm7+n2f1JlFtrZ0nIoghINjHSaBJyPRYle
53qxmezZeG6VgD7hN3urPJFaqUXkXpoIKLAMlpqQKxTj5rql23x1erZmRTxNgK3m
czD+6oEpU+I+IdgxT1fw3R0NX/Pap+lQ0oPZgPLWGgM/PFHcoFe9eRjYgRormFZd
6Qetmxx8Bled4c3s91b3xltpTwqi7hRqysRErraJeWeU88GQUYFHWYapJ3S7OkM8
dzZ+AP1Uwag+fG6kN+IFJBIB/V4NJygA47fZjg0+BUBwt4lV9Oid9rnbyQU/mJ8Q
j7Yi6z7G1vgPzYCh0LG5ag==
`protect END_PROTECTED
