`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1vxnI2Qf9hb9Gt7hOMi/pI6F0bWlpSX00TjCUwSn3PPzKDhvJHsHaucVYrwga8j/
I8pMb2at4HSbvZYqjKMrTPIWg9ve4FaUe1zcP5k2xvnTjyiAs/jyii3oZ7kPFpbf
2VgmOxjeS2IIe1MkCPh30BoqgzyROGqXDGEup2dpCVMZ90WWQMPgHZEzH2lGlEZ2
tKM9seYLh1c+JYhplJdoo19bSXeZzq4sbGPWQGmoMhvFP47pQPPgMQ1rPlImBD2j
6PtBqt+SPCaMNyCPyIGqkL4xV6Io8MXaSntqSnaZAXjaH0OElyF/YC1f1NvFo0Ie
UzzAyMzGskXjKbosfX05K4HVPQSW8zKoyL4Dier3JBWXQTX1ms/CdZY8lWrI9xaF
MKMT4uteYELoB0Mmb7jsYvSdbPGepjEIfarjXTuESX/9xiHR6kYEINMEDpbI43fh
vx812/Udd6lGZ+i18HNiuxkajZ70XXcbVVsrwYR9z0H8VBz6b4fv/1CZ3piXBD1h
1oykN+/ME3Vke9VgWTBkmWKtQ5d02Nkg+BWJjyD6FOaVOhNhkYamkNI1mGoWB3f/
hQWTkH898gPILzFmLCU15PClK8urCRCGc50SZBGzITdbBVLZZKsdJT6gP8lLBZ7p
3eIVJUQq992AfE9YNnc+YQRCcnTzc6k1fZILmWwmFcVat1o+ODiA97SwFWnxCUF9
1OPj9zbldG25bDD/NYv2IJH/CgK5gw5h7GW+FTHWs30InjWb2v4Unk2LEGr9aYwD
7ueRwxzEC+Y0W9xhyrGdQbuSdT89ijAeC7k2W5c0Xk/sZdP6RantUWIpcqRYkjnt
ZYaVHlJKI1ECVqt3VUFvmI8tjv4U8Pse0WznX7azlhps03qlZ78jFulkN1tS/UK/
NUBiXaSLN9WUuwC5+TH+jwWpVXgi1Z30saS4hqHNQMTA62HZj5T+121/rvZgaLqE
ghQnx4Kbbdadn+33DJKCrdF8WDdtdmASVCrMcY+mnIofpgAPiJ79wKD+BEPEcGTo
5u1qVx65ABBpd1NiiX5m71x5igZWVRubhpVH1s1Pmm043OXqOCecz6we1SMbugkD
4IKARaSXblm5AhxBeAfn98MfA4Zfzkvf9eXlcPdofoRfGl7w688ktXR8YkV51OVM
va3rBQhyYere94yLAi/G80Y/t/ZkxsfY++/Q5THkb4zc6TzBorD2Jy5VZGVF/iIv
1ABwcVO62Nk+q5SxlvHubmFuoD7eNzhAh69hdDiIxd4QLt9yNau9qu+qXzKLmB1p
JNZRBhEF06AQFxKpujcbCTIlxqBET28B8hFob2ZpBVEGyWPm+iRiHXC218HgkJPa
hKGw4RPvuS4loeRTXtWRWZCjqsUwavg7+nfAufWLE2kVEIk6BgJwha8mRmdlDdyD
d9b6WfNBIQFS4DGJtSDgQEM4noXSBiMQthehj0cfDXPhZHekQJgKzZWOCGdhFsdm
l54kgEAUAlqzGPqBVqujLkZqdBAEW4X9WpN5cCgCO4ux/3CMh/6k2VKOuqheO7uf
VpJqZKtiN/z6Bj5X3kEp3i/F02BbFCRQPSSSUciJU2dGQu702bXRRIHi1hmvTNoT
oxwUsFfLy7rHkWS+xHHevQ==
`protect END_PROTECTED
