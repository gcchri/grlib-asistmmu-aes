`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FfQby9sTMFW+PlHXxEOmkoAIcwGr+YzTA34WUYk1C3GLAza1MEuCaI6LFzYbXKT8
MoFuhU1K5HnLM3VOsOrk2hhEbpamzEA79aLEdxEw5R7VXWwQh9jSR1R8/erqrB63
Nrw+/bLXKc6hDBf5yLRjmffZCX+9cMIdIAFzaVemECONxik0uBAw+tvNlBmTx6jD
EUfnxOYd3pshqaGQWyQVzHlZ5VVA0O/9ciTffRIWeIaPMdsiW9ENnrdrP60h9oej
ido5JD5SkCZ8zBuhr8N/GLZAPeo5UsFqUt00BkA2X9TuFvsp/2kEU3h1KFMC+EKJ
75d7mSl2t7DqyK/hqcHeTGsJ1+B/5Tk/TUi3FCXvQpRjKL58mHRX+OxU/Ryz7nfp
JCy3vmXxGJDE3VmQ0Z6PcYCLX4/2GpV69h7zHUngFk92ml0PGAvo0pWsdYt+QwV4
vjANVudyNcCDeC2oeEb2zGdSB+MKnMjS0c16R3UkNls9efOsrloEhWQ9/YEGI36O
sXkBWqOcbLRj591REGb3Es+T60QSuO4pqEgQj21T13rC0OEd3xXKNYNLRt06Mpi2
dM4lHy0RrYJRNxlQlSxJmCVqlRprwdSCDOHJL9hHta0zxg4Qv3pF7mm3iR1BVtRc
3LpKEPaIZr/muhYELrWOSqIiGZmFq++rRifc5EGEkNDgXrdi3jmwbnFt0tEj9O5I
WZ85k99YU+KSXbA0es6D8X6DaySIO/O5bODyUKBSVMMn40aFtgwtZGgJGemlF3p6
rB8ZEFFUZL0D7MdAa8AePyrEN6G2JQm5eJq3u6dILmuDTXN+IyzQgaChkw15ZppQ
oLbWghifL6suwwiXy3JvT/68USOXXL8/5sxPcdU8UoJcfiQET1FtO6nH6PglbBbD
4VIVWZrhx+1JWdgjYHGJoVa1OUN6vVdsbRBpjFIYyWBZgT9rIZa+g87fW6e2aHl8
W+0VCGA5Nxvswy+PGi7wBzVaLg19tW8ninapURNtCJQWrq5wbxvQf8sVopVurIeQ
eC7pUQboOTAbR8onZrfTWkt9ryt4nlNJbrX57fy/+juLBf+4WhWKB+D/y0YNtFwD
ySBDgE5fxZXsDZcRmO9HSKF/nFuUSkfC0JGhDQrgDcVTVA02MgdXa49ckzYhkJ2P
LJXXL1Fx8dAUuQHlHHEHLSeaEDJGPlGkqo0nMZbdqdFDmHpD9gYT57RYZgIQEIYI
5i47Alzol8pNFHsbXoYshDjJAN+fwqDm7ZH0cp1RIcjiFwpYZ+ddNwV7tVBB76SS
ovI+U2QIXRWO87agjII44gPtxTfqzY9yiMgHNTbNGv/X6lTh8Kj+g0VLhd9Snt9J
j2bxrLdPtXK4N0pvKAJuvkRdOdtgrKpw9wKOHxuUXL5xBJd3I6/wXvgKFseDVsQa
T1+tgkslOvtj1GrtidjNOs59yokpZT828J+0Omo/zqGoRyyK2C/BZXbDwWvQENe7
J8Xt1zKhfOrkWGWSCMZO7JhPKgMPWMlrMRz7CbGP+Mk=
`protect END_PROTECTED
