`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lbBjy1q2VImETX1BJNlwjtlGlF9G+9cgcWQC/uxuDN4lCJfpOMIitO3M7P5mc1J+
awTPbm/QdNUG7bFQLRnqw2bviTpkvejgZXYrKIimaMNeVzoSkhCr3Ow3FTY7WQkL
F+U8sEJsWFIGdF/He7oL1V5Xv7FkZi9SpO7QIMJ/Fnx/iT6KmBIYzy+7J3Hw/c6w
AEXmgflo8JZnKbyV5mHiv6ttYyIPhHcmRpMN+y10n3UG233FNizKJc8mrG9q9dbf
F9s6WB+ZslF6vwbroXrCRZK0JQf3jqQ14qLlseQLBYKosKjxqPguRyHWG6JTTNoN
LY7MG5Uk1TwFDLSwax034ZeUCG4iydJcA2V9l60BZf7Hs7rKsqOgMcXkMiR9vGxc
faGZj7HntpXyXwOnzxvI5QV66zNaNBJM0LTr/75ihr7PUU70JppijIdTuWSwfqMO
iu9bClMh4SJFLZdsLJmKztXT/Aty9ftVJBEI/Ah20JRDcsSL7L6Xh3R3gR8/Jwu6
`protect END_PROTECTED
