`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BzNWRP9XD63dLH/XSGspGNzKyJiRLuh0QLvvBOy40Zv/ndvU91maKCppA+M5x7Tp
1Wzb7KVVGOI8sv7T442MIYQPD9/jF+9ZE/dBJif54Ny7gRr2avtLc0zhQsbK58KB
CuosgcrbShUlb83TE4fWTb2VRn1bEMVAWP6aE2XzYiZQHPRWYHQbqr+TGJAyPrps
7vZlU6O8tysNbmBW5tHGrOSc62gZm31Ap/FW20winO89CMCRxGnJKTUSR9tURQTL
z1jawYYBNdtq0rBp+Hry8PQD055mCCFlC/Yaiv+IOHh1jXY3FwkrgMg2KWPekPa8
PbFLDPdPOxvzhxtDnxq63yQItcSaSUIFTpRBE6Jsa7omjYmmvzzcf3B2LRrFVS0u
Wqy6sUJMvQ49ecRxZNaT6Fl6dqS/0R2DKhyt1GXkJ7OEPasyWqjr/kSBiRSwW2tR
ga64qSDjKIOUrMacMG41bN3EgPXpX0FkHFfkpFQtT/wHUZRJDf3WFZceLqIG5V7F
YJJ/lY76TcVirkgLuVMm1V7XSlMxb43/BM8Zp4Cf2PeCmm5eicwhTwTthJ+9s5Xj
nxuSkgobDcEhimAZ0KNsMbPJjIkoXms1WVl2Ht1dBxIP9TGwpj1G6RUYl3TZs1T7
3GgFTnfCBf+H8wThPHhe+GT8A04zINaxFioXl124ccoNfltVVRhHDhwNsUfX9Y0J
mi4R++h6aClwXqF9LxLVx2W77xYCC+LpsSjdzxhF40Yk2L3pMdI9dYWZ6IuVZwK8
Zo25xLOTczR5pcsxG0eoqpdx4oD4GKWie8KtMKGeIVoKaXVyIrdWh+CWenFZseBn
19j7d1MkogfA7Av/HQ0ruEb1fOBG3rAOASTZ3aBS7dqso54bTWmUihJ2v6FcLW0T
+M1yaLr3a7+M0ysl+D70S8gdkPemmqQD7JelCrUVHd+tUzpFWKhaREjvABr42PEY
tFqCEm1sRsUYt6+HDg/rn8uD+D7Vp3Mw5wYIKSUQu/vFVhFDMcX6rQlquVSOYC3H
5amST/I9cxkmLtPS9H155QqKQLd6QNlhnXR4m1TcnI0qc1mUg5o8vvHOhGcbmGZx
gLEOWHeFsceICACb8sYWqMn4nad0dmNPUhT6NX5B9Cb/b/+0ReUQw6IvASBRHDF1
5IT6pbwIWttpeGHBLRVAiaWj8J9EZjhWDm/he8DYbxB/VIlif4sr7WWvambf0xWi
Ll+tOvA342fK3HW4evDnGXm8DjAOuAwns0h7iC/zRBXaOFZoxOGII3+Ac/BgzS/C
JTx+56pzi8pfO8zNp05jS4LCVuS5Skx15rgE2b018flMDTPHaQYBXQe5ODDAe5OA
FbzvQuaJ6tURPdgIzsPkKOsdSYZ6iLAptmjUPZ3KkAy5aHhLXhThxc8dgM8e5wC5
sQc1k9zVTa293kbz0b1kpjB6nNI3WL1UEyxfb/t6+7LlFqtdVEFAHypdEjnKoZaC
vaqmecEEb72ItArHx+cIBNmJ2j6aKlYAh0+Dv1OH7htYHBVq0Is4HkphG6DYnaro
k7gEiJp89B9oZKmGh3FvQNddOO0NW6lIQH5ThaKiSgqDLAbOluNLK2YPH7lwA65V
fxm7PuxgRukdOZM2Hcp2ZoYI2OsS8g0ia4F3tx/uToZHXPWOfqDnrOxQbNz9at2R
I8ROLzZjxERAHKb2/tkk/HWSP2z+VDg9xrc12xYj/nQuIuChytYmN2MbztKnYoLf
H4iPJJHZzrLZEIt+bGQueZZ/KNL+vzWn38ZdsZX97+Xc22Ri4wiDXJ+1CNZ3b+QO
BveeiIE/ufcbORq88510ultO0tOrknGwodNzRpvVUFzUkAi6uJDeavc/7pMVbeiP
gqUzYra5S5WxVX5ePFU4qSIWt6jaJa0EwNBU9dmp2dUg40MegKMEBIkbnNC9ZXEM
yN8J9ZcDCG/lQ3aO5YdjiASyMvAfFfBREINdgdhBcT0/JG1mcm/nQT5DbhewiJTz
gU2qrQ87YUxzAthX1OvJ7By/3V+OeDkZjod5lh45nh/B744ZUZhdE7xNqw91awAr
3ub6pBjkmOrDVMhmGZ5AXgmk1khWcZ+L8I52doGGI9nPQskZX8nmy80JFiGMDjKh
xgKHT5V/e4oRjZRhB1W8lEhQshryVFo8VxJ2N49JP09qNs5Pyn2nhVPVgSFPi+2W
MKPVG3QuH/VSTRTfXrSIrEWZ0534FgyKNC8kKfCOfpb6b0KzUYh0J3r2VPsZ+Dwz
yejd5IXaIU5IKmhhcJ0E222T5r8L1t7UNyFl8MqrWSKCD8mOKI8nL+FVsMaIwRdT
7zoLKlRtVChjK3VofRORlcby5r11QcBNB12VTS1l6T6KMpEoe/chTB1/7hOKN8Me
PN6YDMUtYTzY6PPQ5AZYUFi7WGGqf56nbhNlWLO+n/g36XkqFOT6bUKhsbngb5h7
ybYYYQb7koOFb/xugEaLGaRLdVD1RmqkvKeCEZkAEkyEXoKnG3LRGhGNLZt+OlZT
YvNlP+6WXljIgOh885JYzj3aZIyKEzeYFLAeObb+Dsr5h/LFoajr10L3zZuEsoPv
0JZqUbLYEoA3DidiPGT0XJQ1BsqFs3JrQDIU1Hebc+JD3QT2c7oWvD+o4h2FWFVV
`protect END_PROTECTED
