`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bXpE8ntC4zqoi+vrNjq9aaRDkcwV5c5Ty4T4H3J7Aj2wSxBulRJ6vA8FqmKhUs2x
XPtfytvxTcac0D1RRwBnirXjioAcsWGGBlHITq6WYpi63SS2GU9z2pXO43dJnDFD
ctJoN1N/CkZFUgBKBp0wnVq/kr3uSQ4eFwx5XLSrgH1JJFQzc4G+hKkNDx2NLqfJ
aSi0LOLgC1C5B3W+qhmt+Ig6U8WhtQqZ+ABW2OHL7gsIvv4lJEZsvyiPHIB6ReOx
0V5xxK8idavsCREu5amJsu7emW9mt2XNo/UDGRNsIPVtP33PBMtGIFpSEZ0LgRT6
6c8ksIZcouarZyOJC2yHLA0MdOSk+06TAec8q6JY6cQQ9pb2DvTK2qis+uZQ50KQ
yNcNGI52RWlYXlr9uvJCr8bxYr3g+9St4GxAw01VuIYQEQZZ84OWuZvHRZVVxXrX
cNOtgVQE5N7O/o8qfIgTw9GKvxim488xFeFcdtji0Hge0ySCpsjg2anqt54w3snG
96pftLrAHUUtVnBtnyNKsPzBXkKUU0t2sBGuRGbiTKH8mZ4mVp49asxub6BBXNYD
AWrKqlK0QvgeQ5XdvGiPUYwZjqEeaB1KW8tayhJJjsRJlrCkQVJWvOeiDs6ZDdrE
tUC0JbqR1AT0ojgPfO4w50TJR1eJ3muwrhe309aMoWY=
`protect END_PROTECTED
