`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s+3zVvtsg3sPlZXuvAJqu+BfFh9RbR3nOcg35G6a6N5NUsWf5WoI91xsbG0baFid
aFEAtBTkTSsP9G/5fIeHU6ENyriP/+Ijjwqr+1g+slQHiaQGJ+31jxBH6zo4fKhi
MUog6euAIXL9pxIcw+epGZm/bMQG0X2fnCIszUDFCQK+wu7IZ2xd5+tKf9wJn94Q
nhGThNG33R/zZMcrNrWFE7KCRy6zTD4/fJK6b25l49WoQyO7cDNDxqW07NeOxZRv
46Lyo1v+1KoRshBHc0zRLOSU6bvTR6NvCwFOCjcxTYhOp5W7L5ZVp76jEF5+jRPc
TJhgN3i17wbkW2COaq5ZKg==
`protect END_PROTECTED
