`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Firgu6b9LbObO7sC/Ed8pTu/u97pPonhQce1K4hLMfq6tsiyNSGLNYRgIU7dJo/3
oAWJKHCUFevVRwXKIUa12H0xm528kJRtKLYC/cHEBH4rZBYKt7EQFdFfY9vXfQDG
+n99Cgew7ib05ELgYO2zXzosiJzquKHLwW/zLlNCE3zq7Bvg5E3EgPaxD4VdRw+t
aljNwCVZg9zW51WpAf7aJmQKyD2BO6RxgVM6y3/hyCLehjRaF6mMJXm9c+jL8U3O
tbPDw/Lqbfd/W6wAYz1vfmAqaB71qZXQMXkh7kGBR711yJZnCdvlUZdGJ0ckcX/x
d4QCjlKJtmoiaLDzR6xeDD90j6O8ubuC/Ek5mb32tmDr2tQbnzCDwG/6cvLZLnah
9/RZHPyD5YE0tjF3JRULix0O6cQQaHmq4xnh8KlT0vRfZPkQTKhqnGmXqN+3hnsO
tl3BbA95rD63eeegBUAK/IqoDgasFgbkSCD1ZhOELCC2jxYiJ6fuyqjG6OD7l0WP
iPznFGbdSxsEkDJPmdP3EIdhU/9D3HU6pD6zl/OvCoX5bzst94mlH5SCLTP+rV7b
`protect END_PROTECTED
