`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gMGe5PeO7bWsPtSl0V88oWPfKoiam5TahfkiPZEfdYCQKROa0oxPlLf6361ZG68L
6W9BGzys4CiaiEp6utwP23jPU/Njzi2vD9+YO4jPyIEc6UWWWpBPbXYRzf7ji4Co
k1UGiQlnwLBssRFTjjsSHvoKIGOL6RgpeAzdY4gPtwRRqJttJ/cwG8IIpyJF9+uA
QX36UNzet4bhU7gErSKI0buqSxT2t2FwKQBgvGMoSVGIxBgCi0zmYpeWnAulvu0y
7mi8jo5vp4GhInAHaj7N4rKpHDmJ6t3nOj/aUJy++5lFYQS8xKxHpJ7MSL2A3kFz
P0JTa829sPWaXJOyRS6pQWkGmvWt61oFZ4A3VSk8iJeSlu2gluUA7vZOwJsKrTmq
o6h+gNVxiJxFyRoqtBCYJAH+VWqff65LDU22PhMPuJwnTBLtUevapKTXI4g6eWVE
Gdoa38gk0s3F94ePxTntlIUacLOXt1O30Dx/fx2rFSJE+JIQRTwVTjSOvcxIgoSd
txdOYniCYzc1Jgy0AZTZxTVp/ujFPorKxbraeCER/5bsLnUHdk6k3KUwfKhw4GSk
1SEiTFh37XNgKQZgEYv2grR0zEer+dWJo9cL3pc5IxH7r9MekWyTS3pUWGIuOFAZ
Mkm97/gxPt0omX1zr0rlj10z7auhkpNqmdGpSk1BQ066k96X5xxq/Rl9bmvwPUiE
WfDH8QcWsBWK0aZCvHdKUCEpucndsHF5HB/YJjrTsKpG+HpJkoe/6eGELlp/t8R1
ecyE2hb9D4eY687CUcKa+7o7Pq6Ldqj63fYQ5xvmHlykLPRGlnQxA/ERVp7/RmrP
HlidMXy2fnS8UJuyAkcOsJlaXFKvf4POMI3mJKC3Nzq03JrWmi2Zws7mq7iKD+L8
sDwFk2JtbFg1GQf71j57MhpqzNRmwGreAsUEqCdysk44XUYuywwg3jJz29JydMRG
qmUdMkomMzL78PDxtpL/eGI6b29+Y1HFjoG7r9hxE/uKbgYrr4UEHgs/Alm/oONk
LNxXMq38swqeakAnt+MuVyCy31FmJDYUA6SrYY3Xox0bfBqv++omJY921A3Lbma0
CC3OGS4yP9yd2gXO59lOKYCS7CEHYgDn7CUReehNYJc6jKQ3m8UtQhbUAXuJxt0r
zBEZVoMqEdcUTyma7y9d6tE/4B4OsP9+TkEPkLUe2OSvzlcRvpAllbCx5H1ZMLG4
emcIFnh+e6D5N1gqmK37Mrp/4m1HtN/zbiORBzsCsN302VhfV0L0mam60VAkalLX
vlaV4kZUgdTe156vTzAYp1BpvhCLW5RP+Xwhn59NvyC8Kd9dXVMh6hNeDlMKf+ml
7oyTZ2aBtTYacZW+duBEDEJb4wc2Un1GPVarj00x5uFocegCoJJPrNg9wFy+GD+G
0Dp3hSkpqyT0M1cyAabQrCHNzrNTsnx4sXGm1sXTix6GIPANWN1ktu+YrMrw4Mki
OW3mjpux/O2XPoLg1SytkBdolI2JREYOdT9OI8EsqCZq6KoxHwcS4agCgMSgndg3
2suc4JN6AVH7AjD5FMUBy0sWIlAXNo0nQTAaF4f5M8qrw85j0EY/jD1lJWlSz27Y
JigHGnqmw2HJN2LeCKcfz5k+EEuHu5pUOD/DYZAKx1zsAbizP3t2AoR4Q63Xd2R5
9aCwiqqYV16dotOSXzxYlDe4I5cvrS0MTxSgg6faRjCvoAQmnTyuVixYVkZSoblV
blcjslepEO7kGzJt6q7Sx+Qcc+D18UIGUXguHz63oRgNWZD7avrWGocdqX8nEXpZ
XeqTbpd9o5rFGuNn7RIvJpR0oNdEWtN/qMpie2svrZVO8P3eD/z+Ew+p8QiN+AQx
iyqT2rc8VgQYu5iSSI6L5OntpOCpB1kjiV1tIQ+hbEi2ku4adVRqQ8ykMhbn7pMs
4uLW+EHNDdGoFz1gcFtbcu7F/QpEyC43LQYzv86zkGfVF57kCPovROnmqWSq/yfJ
dpWmkBaDbkG69Vvi/Jk6XKsW5xA59LKVz/b2RSh7Wyru5zdsctH8GzGDmtDb/vEo
96170uPkbxwmue4lKsj/VyrvMKnkmU2IJgwOsHFXjDe89kXzVCHc9Gel1Te8nzRq
nThVPL+QHOApnNxQPfo0xA0ybUOMTTtQarcWK0zZTHrf6riWghHyBV2plmcuHusb
+Hys0id87vT4YtyecGU2hHui8D205cMRGGkBwhuqJTA5hdbldD5cPoZ2y/BuKp0t
ZISWxuMiEZ98UxE3jsgDIZ2lL6+RzSjoSRA1cP7nFbFl4LYui4G9VAoq5yxSfCeJ
PSAPvJSbeoZYdMrkpaXNiJ0Csag+L18gZuuGAfgK2Y4B/HjvUBFSVMfZ4rO4heF/
ZNC2jN3PI9Rzj6PSBJLndvQjxGJMJ8RS71/p6IQjk2lbzu7Gd0rTmmP4j6NHkB6+
baLYzBSRmVy9imFCaR+tDwwAg0hE4H5snlY1BrAd0QjsGlU0E0WadNLoK7F7KLtx
h4XcJFu7tLll8EwwAX8XzlqwE9zPczEqI716xK6+gRq8pQwKFmo5+S/lr4/Qg7Dp
LBLNTqeBmImC6emO1EVTv3Z9GA2PM0TKZozIFffzjL4ynp9+12FgngNzNXmcPo6J
YatgIM6pwMqKsNxnTnu9T1GCuwGI8Dqz6DZC5Q12XpnvdOHsdeI/tcAeH0vdagIN
9M27J1BQVagcZBegV38yex8JkwqQT5Kuv0Bq3FkmkGph5gtWRenwXKfvIy6eelSF
jz1lyH/JFU7rjCDtepQnWgNLuGbAd/QlRnWxVNbsKS6CQQjmGSf3XqCNo1ivm+JB
Z7SzAcAgwHWNTqtGH2yEd12DLFEnIvivPO5qcIc1my7tD4h0CZZEKVxLtYUakHld
`protect END_PROTECTED
