`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xQdquwZA+KuxAIEVRB7YENZtUCQH18iSELkXvpoMakXSEofYTkcdUf5BE4SsKyHx
9fy0kAf2TzeCxTjLW4pVtfNp23pi8ez4F50qXjmixF/cfbBeOue997sHuPu040bX
tXucgPmbSFOY+9nUY2yUnBS32sZCALyqET/eX4aTwlbjf7SEEa3skh/8oFmwwp+g
gPfaMeK4IuLsn6Rvdms27NJ8RFRt89J3iGYEvHkblxFOX9gWdl3FVz9JdcLSOV7m
VoGDh1z4lUZm7E4+PdL/OhndPNXhCfF0BG4b/ziCnbDi/ggo/kLRjXUdRM1q2M7r
IYv1iPSSFpl3jp7u7+MtpRNDhtxyH/+BJ1gz/oH2hK8zs8GqWo686BCbpsNVmENO
`protect END_PROTECTED
