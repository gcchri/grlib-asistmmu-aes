`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WL3t5K5KIC16thO+cudzbbzzkBcsV8GpMe6b8LwrY3ZGewTS4fV6bwKwD3zG37h/
6NFDsEgpOmceaqC3kwFAZATvT6gFcgfGIr6vqpp4HA7xI9K9W/EAihNbshs5ZDl9
Hwwqu01MRuVidxohcTBTBc5EcQSogxInqHtXzwVEziEbElEGrexElFYmv+IL2M+H
wJOIf/aiDY/pgbA+iQaHPiNdR90/WncEEpKeCId2KyKBjdkqPBRiNQyI8tlyrcZp
yO38hMDm4PCRd1RvWs/UD94b7Bx18I+nMmvwak4YzOMatXFPVs9fcvl1OGFuV+Y9
V5SXcFhmxk42NpkiLCjXxWN9j1mAQJ08Ec5Ga8Zwpw6o5u5amyemNxwEqVu7YQyM
UCpDWQzRFGPXdu1I2P10Uhra3ba84pe4zMYER8Cbmpw59i1DtcHGrRX4Y95GqcoD
Cyxs3/FMXRhvIFd1QX+9+ASPMXsyDn/x1He+2gkkxCnpfkT8j5BFLZpai0pCCjtp
+mOUxuyts9r8aUVjFsMvjyLZD80aF6006/t04L8NZrIep9rF5JOI+5/EyhkqYsME
NNOjxVElh1g0yXZ3wuQtpSlut9IDQhy0Fkb/k6azcphd8U+q6tauJ6ljrOBhPb8U
aewm0ySfh0DwQjow0wL3fiqhWK59D6If4BO+JWMQNI7mP5T4r8SGtYmVp0zetQtK
ZYdl9K4DGW/gWaJy6KbX48LYeyJcFYdhonsctQxjkf4cQrSbdY+qnvPdG4NRoM4r
+PKik1FgT6uzJhvAfYy1+WgrCbKJV55/w7nXkr9wsQIQF1WxbEmTy763KD7oGipA
nLH1GfESY0RdgadHreDoaldQIP9w0L7ku4GA5/JgytjPVkyX2CKpnAA8mlaacHxf
1B+eM/VVYMqytIKIW/cecDQhqEG22tN4mPsEO/9aW30nFDT1dyawJ+qyzcCfLGal
4Rzc7AhMaFZJHjZ80XKrpq6zRbDdVIQw/rLi4kG8PN4b/cLjpx32tnj/kYFY5j51
YyQV8B7AJRPcc5XCh7Kml6WHlrj6TGRFA0apwy5ffOQ6z+WA2rRgQwxNK+Uk0pIc
P8jzW5v9DjDjAdpwsKwVkVf1L7HSNLlG/xHCHsa4wayEN0uCAaxlPcJ6wHvLkv+r
6nmCO8BfxORIqkUpAm0Xoi8Wzr4EpZM6xtwoN5JLL6TjQ6mOEVXZZERCqNA/rVw6
MhaEb/xD+30o+0ASx0cdghnAWIj79hmtYt1j26JlAJm7FFi7dbveKZfu4N4wUjdP
MTxvx9pmzCk/X8Si/GLe01SW1XZBgrXwkxPySpVGWzjA/kTbBbJzP0rrYmxU7tz+
vD3kDY+Jxvii90Tgz60EqukzW4sB1pnyR6LKZQGgXMQ72pCD91blfIZ0QKWp9u6L
DxMrcn8YLq5d8l9aovoK2IekLXrdE1oDc3JrREBcs0KUoj91aU1mS5LDYmVxGKrM
q9u5OinD56z5AsZTm6sLA48+SAo2/1lChzz+XJRLAl3ks3hqSWDJHc5Sptw1FWsq
TlK9nVfol+7CHByarswTd+TMdX3CySlUF4BkRyvODeqwaV+I3kQCCgFLAsK2lZrW
tFynnttEWfD7Mx14k3H3caLDNvNIPemoFZ8v5Iqx+zYz+tyYVsi0UgwcvCDocTPK
3Lu3UXgYXdwMOBG2l9p0fRiRkYTLZ88r+N6feD8xc4Kwla+LtRw2vpKLHVO3+C7A
PAHrCOapRpc0BXkEd1Te78jpcr3YnVYkQjUTjFBUOJrk8fNNZ7ukS3JZZCO1TaY7
5SE2RV3ryQwbaYv4d/n8MJelSYOuajJdnPlPw8Hfr8rsZkwoGgpB4RlxTqwifPVZ
c+Gva6LZ/p5aTY1uIUaCkFJjwsIwWCMSsdowAmBThti5mJoYfwXy7PhgVhq37LB8
CZ+5IZioSBQSa/yHLmN1gVyHGBB3Qwh6zznFpvQXFzHioHa7YjOYwYw5tw5M06zd
m119ql4UUGe/R8li2SYf7Z/MoFA654etiN3Dsihus+PkwCQRpcNjyfFl6PHSm39w
yBed9Ua6VeZ6XbWf9/SA4KFPzEjXBGk0LshnmXdxBPl0pdDTLPEmfolME+Tf0HlN
aEUDoZAbU81juYugPbabZpK26g1wiceBUB82CQsnszp3kYzqT+k6x9G5icNakt9/
YGox6cf+90l8BqfhMxT+udvOPOLZ+iikUG3UKoY30k9VemmZMPlSmCN46/qgH5FL
IBEFy7QGHSNnXZWXyGL2oGZcQdGJ1kwNIZzvL4/jojLfxgA7vQgkZE9CcvLCb6hG
OYBRxs84H1rhOlyuSnMbGnXoRraRAJjfK2Td3u7llOqVv+AaGpU0gVSUhkdi2qW0
8vVMVP7fQerC9prsmYX4zp/+bO3Vli/2tchySkAC6p04Hf7Nn/dh20Rf7f85MBdv
T9T4s8i696Y3ZlUN8nG5IRkBillPDjlRJ6FwJgCmDQRC/djjR/GHV7ya825D35sB
i3zUYBUW6UhrUjicMvCIggdlwi3xrcSg2qU2iqJcz990mvzjhZjdgXL5gBG8CJTR
qMFGn2GQWhs8igMHHJjgpRUzTZtD54PVqNAb3Rihq2f5ZX1kA2qa+ZPvhlTSNxzq
YK1fMwSMBWv5dX/oqcskdw3jhWnNalYgoMj8P2vTBdH7kAVc2EDzPGRqVW7lzUrg
VvnvPfxu+yE9h9Myk3gxb9WLmfEkvVLUBIf14cEajkhfOz+93ntyE70wl3B4hyIo
kiH+auKBIGGmB2ylacs3TjOrR2O2hxcFlfDIwt8taa5t+B51hsGJOVap0ofaeEG9
d1LH0vCxY2im6ABQkFROfgtFjFjgzt+ymxsLG9Kvgo6SPfAxhUzD0Pq/oRdYfbDF
3aat0TgyToEu0IQXskfwORmwM4Z//arKBfQIqWlb2p8/XmmWRcfgVKUq7mYgu1G+
UuqTA/LOuzbits5TcIzuoq2t1NZ7g9B+6NJzirjlAi8lpG+NZlKy/3Th9vftc4eC
yTQhHOY8juRbXUgchuGfDcRnVBbhCujZWb8lkHXUmmY93BqIvgPdSelOZjXwWk0o
7tWPnhcq4KJfUXHxBoKjGlKF//H/dPBvQJAbRYsgw7Zs90Cz2hbp+EXboHgSv6K4
jiDiquwZS3+1qoYrVSyvaACdavOENuTziLvLYIaL5ybthNR6TgW94YvthwTNLZ36
tt86r+5FDx5evxWkuVVpQ6D1X2sP7zQ/TQXD7DCv7LjGLi+sMl82QzJhuQJH1MHT
vVxUfgUL3xRmKLhkNw5MT8jNJWlaV+VRPasWd7ayc3t2takP+cNeq0DC27WPXgW9
zlvr3iSOaLQBba9+ACx5dLSCX7e5Rvw12f7VYs9gmMsGp3EP/DPrldSV3Jpa9O25
jWfzFxYIEvaGWMl4yQ1+gdI4V6JN8NFes9gRIzkl8IFmMoY8AF+oSjUxvLyRfry4
P9oQj7NXl6RPyqgEmTQlcHGyg32I1QSmiCphIsMFZeRxhdxueX5r0vvMwv+1fHZn
6EGPEF2PoI2kFiCVenXpo0LSGNrZX65aE0xNmQE5dB4R9SAAyCr0O55w4bl7x9J3
`protect END_PROTECTED
