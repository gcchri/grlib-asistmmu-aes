`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IF43nYSdHqRGXBUITRE+BwKlh8Ycg0wLY8qGYVmzIO9+P4DlvHLI3ySM5Wg0/Zsp
QMjcmbrPbr6iZFNXCvyxZtM7CY/r/EAOsiuIEHcKV1e9mv5DT/beKFnjjKYeWrKG
WVYEo1ZYbuPc/CM3ekc9Bs3UJnO0bHOtzHvnS5mEIsqwE3lxcG9UHU6yHYoMa3JO
UuLN+7AoIG8iLoJtut35qFdWd51inCoq8fHIFv4TryDnad97JPg3JKh1hlMnxobv
ZFtywLpCw3r+J3an6h5XMA==
`protect END_PROTECTED
