`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+JYhcsWiAmaMQJdqMu8W9d2IAwqkB3EjNnqGozJqIqkh32+kqfPwHW5RKql9Bw2H
+i/vHx5QwRXSL7fuLGQoos0W/lYpcPHAjQ4u/dmEXKBlDoFzv8Drxb3d+ZhAj4vu
HRzfm6L+FeZPGtBfUA5rNIurBE5jOpAX1KzRBWshRe6hdlGZ6Y7FSDuok4YHAlsw
Env5tPlJIexQgKzwgGbQpCLEDRFNy1WKIB9tKe5gEMjCxXCIwuFO/PHhDbSOFRXF
w0O+ewuZPB+e6Nl4TN6kPdDPj0EVFijfIaoyZQ1n1PDC7fhVa2M+NsGU5UQfU1r3
BZZ7j+nYrY816l7eWaowx4fuUZ9XSyt0RmZvuJ36iGngWOIXr6FITwpHrJmAGfty
boqRBq5yCI+aAds/l4AGWqKIldPmJ6rVZJO13pjvHCI=
`protect END_PROTECTED
