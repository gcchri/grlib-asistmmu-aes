`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fCB0EcWMHVHPvwb9HmyI9XpBgCjpghXQbuCScfDpMMIOZF7/2eE+Sk24yhn7j4zs
faYPiTe00soDCVZ61ln+ZXR/fyyhk/i5XYCaoScbrHCsZXGmMDYe8Nvb+OXRD5bs
Hw6G+XbiGpHfaBq7TOTMl3rIh2yJImEM52u9nMWecLIFlLC9Iep/NB0l6WQB+oGW
ib61n7ejZOjI2s9yfC6gAnseeG0uXme9Qtq7AwfuvV4gMWQ2b2gym3xviTqHTy9k
ocjfgqyIdTjoGFTfuLciOhn/cVHmn8wVUe3LBctgmseHzLbHIWbCDEqnmk3ZUwM5
7erRXoe4Rsi5eu1pg4dF4gnrkFMgfrIZ4E5dUcu4uCIOEqvXXNGYxNvJ7ZtXN0AI
r5eqJ1O5Jdm9dps90rWdw+MTP8ejCxSB3BMlXd7FJnQlqndms8VPFSRbkj7JFpRj
0ku79drbyxJp1BKOCrK39ON0alGbcUax0oA12WiJT8bbQbmtnr1751GXMM3tKBoQ
WjHBFrtDB4odyxK0QLE+bgEG3XCSthO7RHUe7KGEJ5lxjuujdcI6JSXq1wjUClhw
WGtqJFrxE5Fy9WDlQvUm1wVDPi+RhlBK/Vm9yG0AWohgHCWDEJUntVUEzc1bKbkQ
sOIoSZATVlkX0G6qbO1GZXgFRKmZkCZ6hSVWWb2QkehriLUktAjbUkw9fX1Fsn6I
egUNmOiZIrUJSOXs32NcuyAKlVnqw7jVAbUOisFlbpa3PUAc0a2VQEYwI2ZhR5mR
iVm6FTCR56xut1dR6IGoMbcweHlLfwDbEEjyIqBmlEsK5uiVIbky7c245eH4VxVj
dQG5n8DVZwlbhBRAvl2UHfD5ZoFqmPFDSWVQ402c2WCF5cnN3kZsyBjkxXkENSWj
qWH+bCW/35jCGwoknU0XaOAqsanFn2ByhMHNKgCPMpD37F/9AluvZjq1IseM31kH
VimJtKO0P0NMD0hN2F92//oo9uUGutiQ1t9Yc1OlzGBHYidi/aKAKhBVKlwH2YJX
54T54rmHjWwH6Mc167s3IMw61q4WM5zyn9XV1MhLIAIFQKhDcEYLTwPkVT5WCZGi
l0+2k2DvSwbhu32wGHg5kcJ4fjetJxkFVt7qg4iRA73saCCFskXUjV5lFuPeKPI0
xE2ISpFHmofMfHTtIHxt2QSIoeUYnHp3Q2Oy5hwaXUuZreqCm8eq9eLy4VbFVUcT
hXMAUXoT/oGMfR5Fap56y4kNbwrogOPI67ODcfKWr8uy2jyz/XXTfWk3HzAraUcD
ZLjkIpG++6iqvi9F78YoMIcRBBvcl206RgRn5vLX/mFYm6P51d3F98bM172T77Sy
cyJprZs65EwLR53d+dcXZO6Y97lmNH+auc1+ekqM3ot/apiQW26NP/Hr5v68jhyJ
McWGjTOznZ9ub8QfNiG4Xa+G2zaktJWXkkEs9ImKaiKVIv4/ORoGu3TQi1bGxRHV
lNTNL4pH1TTie+Fsm+JTOAvqq/tPjXEf4z4Qjl7y4InBuQ5PYHNdM3FUdh3k4Q7a
FkbJKHRqFcjXysRVoSFmd/lR1itj0CJM07yAwhWK3bv9wZmJbzhW6uDxraO9FeRX
zrbAI6URVTWprLNquny7pTlHJZetDP8abfmaAQfNVkY5E50yLZmbOUEeZhw43tXB
flwM0cEkT3fw3f8yJeRcrRZe/8xyTo8ga6yVva1y5pSFFYRUqQ6D5GTDO/WxZwJA
wEaTUuNPcmRDnxzd9pF7wtgJKdRL/vj2s+fUHVx5zm8H7JS0qy6f4mZowykofxMp
qMxEYw1ZbjrxtSh1FRXvMIDO+lmm4D8sRdWY+LwfI0mwPuZtSbHkWP5TWFVQ3Iy2
0sUD1ZcW973lS7SmEOugbA==
`protect END_PROTECTED
