`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9iwrBvROGBynxZ2uc3OJpBHtAS0ouAVwEEbbmlj2BKlMsAjYlZWnNuU5QgOP+Y5K
Kr3D0+dSB4s1B1gWMp2Qci+F6xn0nifXEZxlRYvbk/QFWcc6JmPqDdCIe1A0e0rl
774mZ41GDQjiMLn06XcqQMDGpjLI9UNC1Oo6ZlPfN9dN9rD+KEVhaybdBRsMNQvC
tGz3YMuiMSzrHLsMZmy1OoBCS69hBRBsrX4Hgw8Rvk3dtJsJMf1ZdqcDcQvuczum
x3bcuD4jgZaXnh/aIHp17q8JgxjIqt9hAtf8oCHqpJy6k8YTuCYunWaVpgJH7HJd
IDuIURwy8QPzIqBzUp2z62WJPFpnjjyNpSLXc4NBcElEAP85UP38F9rca+cSbHA3
fxahs9FbRnrZOgzmD6GlNfY484clv4TbD4x1YSimwwtlcEYT18TqwElAwJEliGF3
V04CvpTUPqjCeS+qWuOFjLvn3CIqFzYYoMAv6TjtmGTTWjlTnLbJz71KRj3fy1f8
ApwcBG5i+pJnX8lxiD3b+KZ1TUpLRSmkW9Phr8UQekXKFBM7BGA6LYTljZ5YegNj
ZlPtnK4RoHAmIxfHnWl/eRYOMghEMIt3chEDoB5qPaxBNAxKiqHn8TWPRZkgKQL3
DJtSvmhNxOrq6Scuf3PE3k6AL2nWykXjbJ+h0i3FSoEl4UiihEQzMrLERBEoWPCM
VwveRsdltmjkMOhYI4cKgXYk+Z7EusuGffPTJjzHSy6P2OHOgvO1ZuW/5NMsYkmN
gDrT7zW830o2YuSHrIDXF5KT+DJM1rAo4XyaUkFYbGGd7YPCqXmdj/3UsXqFf1Wu
+m5FPBC9ZuRZd+nuVaoA+HMkIUO/AM+Ji4MFFNeI9isGX+WdC6CdZj9nm9+xzjW4
0sDEWKEm6KFM4D7hzvNI1CMC6w+/TdmXp7sMAPge/OhsuHXdGkBX47H2YWfUB4K0
tU0gi1dcJ1BwrXb1Aie8ecq8ga0y/uF0Lx+2WAj6r8JddyN+6sVGQ8m/zdzIjIMr
`protect END_PROTECTED
