`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7uJAFh8B+hAZIei4fgRs3epaXQYnGrwCyKyJqbqI0eF7v5zr91jOu6hiuTUJ61F4
mRXPifnoUtd8cgJmANRZny/e/jsD+JTP+WOX8oyBuQ8tLjfdvefREM4uAj5PWrrP
ucJk+PxrA8U6f7s5wZJUgtASk+E8hgHisZT5awOJx3msW+F/jWSP3Ux7O4fWFDdj
hIQ3TLk062f5YWSGIcqRxPgpxg52hWQI7JuQMTTHFZ2pO34oooYbHHnRm4g5y/hi
CFXpuF59Ef8OtHh2V0RP6O7p+QhK7aaeFm90cXGqFvdCT3iUOuMaHt4/m9scfchp
5qfzGq3f8F6N3CeqRg1mL7miEIqmAgz3v1SaJ5PaTTOVOSH3cNJrtZBmNIuljnwF
q7Wq97gAGpGNT+Z8R8EA6+y88v1XbRVwW1VU83T2Lz9/VeuH+aPbNIYjF6v25GqG
YBFlqEuBZgC0yfScLvX+71fwo2Z5BHakPpCHvGmdFCdeAk+xcYQyLjFZ1lk+rSYk
v4BMStVYAtdzjgUPuAXGfucm7fDXDVSbzek9kVFZ3rtloZEATQZk8nc9JU010Wa4
kxvC6yscuitwmmCXdLih7uNPvHR+ALej5RQ2CY2w/RsQvNRvVkwlN7zKPBTHYAt9
FlkSn+NdUkl+arBvKMH4Pt2sIw3MBmy9Hzdk6flaNglRyjKdw6HHybJTPL2qkw5+
kEeCdNsqP5DRsazJTxv52/4EdvKVD7rp/TvcAROOTxcIQD2MMrbQn4UHrHNSfB6F
Ph4ngWgdT2sTmLC3YM+1Yo8atXz5vTHkytHkdLus8fTY9SLs0f3pNrGj3uMEgks9
LrqqQROwLcvviITcUOxvCatuclpkPHSY2hrxkBLMygmpby7+tZv9EUEN/8s80/wL
8/g4p5tYgVIFNEHrFYXVfjZgQCnQcWcxXJxbcP4D1lhHSBzZ0eaBpj+d3o/9/pa/
FOCgwT75Byyx6qSzOJW/ZYaGCz73X0bzAoezXVLYPAsmJN/btIjzCy+zOnHfvqfc
VnxcDkheOqq1EPajMM8drQVAY0iHl5ADBUaIIYZhWEpPV98mY5TCs6nbDv0e/2uY
cXZ/755nmfUnw4W+vDAv1uKAt90G6fTJtQPne5dJn4iuQtoJw4mUZ8wXrxP+hDhp
6CM1JBOSDU7zebQasf1YET+w3+6uryKcXc2wTdbwgksnOV4iwH8NiwrA4Fqv6QNl
A2rCaajk/KvV1TKMddC5Kgy3gHVx9T6O58d9bInfAWlOa/8Y63i9ropuIpcjdGAH
`protect END_PROTECTED
