`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U3udhpDrImCkwZ/w/s3UxDmf/UEqN1HtTkpHqwlViyrU6ocVRpLqYwMIYmmgw3NG
ZEAYSjOotraxrO+hcrAcIu/bIx4+UoGPXUGHCTQz65fO95u2mRDpZYAQyKCSGkmz
IBO37xsbD1OdSKhux12wQ/4cSbJsOs5GeHe6IH7h4ptqt9tpPn41l3k5HYV5a5Tj
zVNu3HH66r1usyZuBzUFtu0L8X7YmOehpRwrYoOCP2UabWTp+cR54YL8+3slsyhi
/bY+NH+MGd0Ww2JQ2WEZVdjAYbzQpu2aU3GrD2GR3KG/9ZJyJ8rPVhKY+XBDWvWy
3di/Xjw+SfQIMXEUfBlit+nogb/N3EDDBd821LP4SFW7tkk/8hfRiYFzfda45amA
O2AwpoBPjCroMdPL+T3pWUBhz0zu0v8PlGRa/i1VptTqCPP5/TGI/K0HWu64GMUl
WzVbzDpx+GGjl3ImnRqp6GEJrRhGjiKBpJ7Tmk1gcD3XkK+BZVVre2UVAOc5vs1Y
4lXALCAgCyamoD1LN21ZjU5XCEN/3xcLG44FRZ71XerrrK2TwUHj9qoGSwOkGAGp
d+EkUTO8tIJapKAtAuIiiO4IIc+EhhhY87lctob+6NEAORNRUb9YtBELjPQFubYC
AuWoLuKgRz0ZaE/ZlveqVQ==
`protect END_PROTECTED
