`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OC++AQkzyezlZVZMaRvOTZFw8zaymy/DTbNfwmZvgyAIsoV063DyJ4s8gK+/ZsH3
1DpJgKqLtXcK2huUc88svkSbBuPZKjqNg6pTt6x0CQYCTeOYiRbMZde1yNJ/1tK2
qkQh3X5RTOL2d/cuxuluiWz8O263tkeVZ5wvT3j8/7bBV/ZOiHDFGHlpJAhh1ebo
0bLIzYJH5JNALBgM35SFF9v2T1il9i6LhIJ3T2iHQPG8lOGwZ+Vs20i8tuzBQ1Io
ERd4sFtGthxLT5QiFOPs9IXq03A2ykSIHdSvp2c6LIqstklHDWaJy+AGseNuS5a1
oQAzS7911naNl3tIDnmlUw3qW1+ZADQgjFMUwn/50uGfrCY7TfYHMgP/E8BIkA/L
2MkbNJqI6qul31yg/cBNBzZUEjJFMMUIFrw5XCigb4P6XpfIrTyNeStybLqkdxiV
wL9FAWZUvhx9IDuVbKc5m3XLvX/YqOvx8rfoYQolvbvLB4bixy6t8lUUVwHxn4Hz
RLE+T/HzzFHzVi8WY5CTz0cV3lZXyxklKvmsP2it9KjdWHf9Uib+bEA3KRc9fgHL
jowm+nuLwC2IEBl2x9+hP9AarmLk1coUyP/moSdfUAACXqKaozTaDrEYzd5DjeiD
lHg9t2VJ5sUyLjviRo2hPh94vB0ZHOMzoxAfZu/Wzj4bOQ+mwy/M7hCg/QcEoLTU
ZqNQARz5rLKZYMAOoIOIWmJfOC/vQecVIvugvD4knhm0nlAUQ5fUVqEWMfEegQoD
8MlllII0CQPlGv1bTo5L6nrMbKjkz387I2lM5XhPkfoUtqg5ukrwutgSusLnsneh
Elff7X6FSiZiEETPIqlR2eZ2AhHO5YxIAWEON158JfvvrBQI2JCft93q/ymZ0S3D
WReD1eQMS3Gw+AVt44S3ZKkcbjCOQoFBfCA+N2WHwG4fJ3VBfdA/Hr4h1/EX+U9X
1EUBrBjzRiDwTc3G56FFF22LexXyErUh2nOYITwGXE0dk7H5ZkSl0YIteljTF8qN
2xUU3vUQPre24BKuWMjh94xO/2YYn3Z4Dl3Pk+naZFS7MCqM5Yycq0I7HXtsbQZj
KSp7HDGiba0wJt+uwm8TAdbagTkSMP5zxUD1yT0uPfoULGDjYl6JZ+m/CUHQpVWK
`protect END_PROTECTED
