`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hNsyeeBH73h4LFCsd4p8Ijy51RLWGhJuRcZKdQXmI0Ar6rRZ6MrFJUMJg990wx2H
2UOsllhJXkPJnPFnkfRWF0NAINVgDrTiSfuDzD9zRRlzRwwZ/ekV5wT9j32y9x3S
bDlRWBmP6lPgwXHfkRY64AaDGKZIyUcfVtJhtyDa9o8HuTuEmu21OrF0OEz1xHMK
/KKmrtzLk6vzJW9lzrhEGStrJ+9JH8eF6ybNv6T4YmLKtHTGA+B8UiABWxoGuFlg
AKycTC+eVqV4jpyQ4bnJRpEuvnk50zD2k603tDtvu7f/5KrSh2O8oabp+BvIJ+Pd
nV17ubmIcepRQS7wgIRMkHtgXq40EIkgLtNf9nP6UB2sGR4c6vlU4iXlWQcl/sQ6
qgK0mlqQC267xuoiGwq3nzI47iy1NbK7/oDEIVnyXlv/e4ZOB8TftUitURfhqowG
w1Vu7fT4CeKX3w09tgEn0qX7L5OWnJa8VLUC2VXOLw2Ol5Bdvf9gWAqQm74RFVvJ
qDQVfL1i537DVIjoorIGrW+Lr59nl9eubAYYNhUWEqSwJPFQjxTySP8cgm3wvI1c
khHAYuPPclgv7tufhrexBLoRsTSiz6Juqmo4RY5cTVlzMTPmJ7qGwMoIjVmnjY3H
px8ogsXnqAd0fLrOIUpwAA==
`protect END_PROTECTED
