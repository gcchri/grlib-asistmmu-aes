`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NdnkTgo280tPityjdLctLepvRLtsNWgWnggNB2d4LvYbkER6cmMCkFI6+v6RwcRX
J1HdyK2dxWFLEP0usZn2lQb4vl4zZgX8SsG+6PcpBZIPEH/T1LywOI7nSAK9GlAL
ufBaHLYMNRPn4+HafZHTtJXICNaOvo+jeM80PDq7D+VSr6CxMhwZWekIsfa71jse
xvfDKDp7vpHhHARZlCt55q3Io9XBI7BdRDklFqX3RZUfTt+04nCSG/rUFQypAN/0
YQ4d5+9foSXoSafru9c5jg1n5auLpQuy6TSfExHIFJGHiDADJ8x4jwUg6T2bWcLQ
G1md2TL9kb/FE+yFv0XFCr66EJscZSe2fwm2oL9zbTXQ2FEEf+EoG0n0ZwXAuxYa
r/D58yrcKKWnYFqxj810y68WEzngVZ5UTWUJXaAz5BIQldNnfXJLGdx72uxC4ggb
jzX2MZwUBuXmRJyqRza+/Guvz/jQlHVMwL6a35Aw3hQc6OmYwPTydmGTt3WuiBSv
deCYmQwRfkpwxYmQcNHi6c6mlPej5kaE6PBlCeTKUdmxTDzbdgNFW/Keq2scdoyh
UGoqWMyZ+sPgoWTFXsqeSuXwMxNAwW8MqXh7GZNSB3dnp7NcsrMTlD6y2mZgWCQT
IisXN6WxafYCTHECAax20NaOpYjgRLCsrU7yRNrGJIqjQwsW/PNtAESG1E3eLhH3
8QE5zkzkOx6GH99dI4QskEl/c7pC6zhoLqBX84ku0BiLrg1xn/GRqNE2+yJTcPNB
6yFUsAXcRXuAcD9mLgJfBuzpP2srGVDFC/Cypcz8AnRh0aImtLVQpB/HWbItYIrC
YWWFqZoF2/0QcS/4J2JQak8hFNxSzNX09yn2Yg1BIfikDELyCfsD4SLZ1uPBQhFl
IARK3CKrona4buT97Q086T/J9P6B8DXn2463sfLDyWETFHWorWV+0jmsz5NEYizd
DB70+ad3zL5s2OybMJIOO2f5kFhdDzMsImZC7jeiQa6gnVtsvf2f5ryW4KDpfcwq
2GuJ9B4GxcluDxXLyaFtpLK01ljfxcG/DYfpN4FssLQpdq6v47uznALX8k57B9M0
X0ZhoufRos2/sCkBtdGprePt84brRl3YcO1QgepgTPc5Zwta0lW1oT8K89ckBuup
TYNh0jeyvxRJN1u5cPfCSM53WQAnz3YXEgvaVoKO9SeDR4+SIzemsJJF+dHTKOr7
JrXkIDhhRGlO2SVDgCw3dGnn0zO6cyF0Z8mYDfAZFxuLSyXKhZYuHCnmmielMUDf
KPFk1sN9JcxRXHscABOkYA4AqzkYUElnxR2wsiZ8lbMrqPkV4Qvc5v6h4UcEj7uD
qlkmk+6wd15hjbxNe63nuEYr8ZshfcRVjinXiryoVBgeOUvo/AoDfFJtu/eR7t2N
SsQ+VK5/6a7MTO1e11gKUHkyW77j8FywTBu0o3uOGJ8CR4ISpE/WKxDvtB2ucqru
7dar69jQY3ZskgEVKFbfH+Ll7OIIi3eQji4ZtBC7hoF0rMZJnWH76oqwH/MxKRmW
POdtqj0trdJEZT//7ZnQ1fnhELQUcmZZhb7lmdhqK3953BqMgL4XoiBsCUm3ZQcp
GZeiMjEMs55/MUJ/lgo+ik2jwMZdkUa4EDJ38PExNRh+COBgaXamv164gwXll+3B
R07LrH5TxCMqukwQxVJr24B28Xo1eyyCX/9tM4mglRqyVuEZaT0VhITjvwbl/dzP
XxEYPb2MZXEHB866U6Mg6G0oUvOfbHMYS/2rCru42S60qb0XmbTgaraPb4Bwsb4j
dixzb1pLe1PevApus6nE9P+T4QTZC24V4bHQrHDvAuF60B+7iFxgkMIj8VlPEaUr
Br9WW/Aj365vqc99pHMS6KdRc+ViI1E3bHWV7kVtWLdJm+kBIOddPPCPwDb4mp/l
W27ygrTcRHPS1NMIZgKh4JpJ7ZRncopVz3k9s++nD/Av8Vhj4zbFUzVXQNOu705w
P8quV6mO+YfRGGVLxMzOVARqR/Bj+nYyi7YgPPKMRQORqBF5U/EIlSNLwYpPReij
xHEXl3KlPQOhGjmKGjRJW8LUyb1WUrfrlM4CyobdtvH5c5cyxvTdWFR3GVP61RJO
+rTPJClfR+7Idqk+dw44xVH2zcGhGBHM4YrpHneL+j7LsBII9+CAgOb0jNOftZ4G
LwqLvM/TzV9x6ibuFN5AsmgVayt16COi8ZRwChfd29fIz2DeKEwNGTJ2c0AlQHxp
uq1kv+vXwD37yl2C9DSBHdh/K3arfQabXYYq4RX+MCCzSlqydiFLD03EkAv9zBhg
lwhrMv/bhr0epHyJ2zErCs4tahPEgV245x3w0Zc3qwOypcoNhmMmxTpNQiNUPn7b
9/QaK67ifRwPeMzgmBdkQwwQpJXZzo9OH0rXRff5cU/djKeFARUBE2bpVY2NFblA
PkhQop4ojPrj2RwiFeMeCWLQtfoZo+YLRettqyvzUfA2VBtMp4A/f+aCc4SffQIt
osxUDiEcXLzdbnuX1y1U/g+Ezo6BjDG5kl0qcN0DhidfRuCNzkW9jiCAuEG20aAC
i1ZnVrALg4+9IZdZHSMnmbQsu2Giin6AxLDx+q9Zdo4Xd7khEhZyJ9ijdZLbLCdh
KQiEX8JXxLIG+eLGUfx9wzBtqTwO4jYcSN5e4Q0bKWsB13IaE3UKLbSXeF1qMdSJ
9GWROfkbjv8XRmIH1gRHOyvw8H8HF2nn7zEit/l8m45IATdClF9SS/AcXgZj0dsA
DF1US6kpCStIEJfqszPo17x2B1Vc6v1M8uH6+kQazVpBqrU8SeoFQ4in8QhsE48s
H3WOPEI0t+VQWUEAgYduihMOgcTBgYr5Ga6Z/7+DBV9LCoY87/3IQaxfd7kjRZgf
FzWBrw2x/BbkR7d+shNtKeyKOx8ipb+hFF92NcANGleNYJSHe5UbTb9FqIczM5UE
EGO6MX7xYurVt7aoYWkfYnnjq6duiVPQhmu5xqznZ5EUJUAuwYBi6HY2nZn1D3MU
A/2sOPEB6Z5F/KL6e1GpiJXg5RfR5dZYDUGY59m5HfbAN2ZrVzerFC40Vk+mJukk
6D9rGv1uCDhbCTVmj9QSO73MuChU/ZDvKceaHrK6tI1f+wQoHJ+nWfzfOKMfTDrh
`protect END_PROTECTED
