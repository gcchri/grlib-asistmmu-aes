`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dag0s2GwPVSNxu+ji42B1NF/SaOu0OVeHEfhAxO/uTWfPVL4uPmS6mk/YPJFaG6P
C30DGnUWwcuSrVmJ9C1v5Td2jrnVwpuOqM9CtFOB2XaFua7c3tXP0AJVjMltNz6y
jL67hDuNATR2VU0fEaGNmDmpOANQsvzcKUL8Xrhs12XKIdXNRo/xxA2EoYQLJq/6
BhiIRgC1PoNgqq/aufezjjtZ5RRi2Ny5qGkCaLKgxmuN/IyhXq0hTmhiZ4cl8U4R
YZTlgiiL69U29Jw30uJNsgZCG3IRYbdXG6wct6TSZBPYgxjZ1kQP3RS8JwgLEXH3
zhwTYPpfRCdudBdHE9q9ZH45Ety6DZ1jtuI9BlJGW1sJtYzPIITmyuXHICt/hQgY
kNX+KKc6OE2Vm6fHQ47J4Ci2IkEAAqIKosyDmNRz1OP4HIIOiuLkx6gq6ltNp4D+
p22GcPYs/AsExdRRRj1RdoMMyze/VddywVyf+fCjmfxB/CFqTGyMhrSoZT5WNA+b
u8Dq1e8Y1GyeKUQrd0CawEoCAKMIrNielruZbWjRYzgLJnLAIZWN31YRNXgyp5lG
oxSpXGBOHMzw9r6x/aEtbU6k0Zjxf6fe7kB5hzIsZvRjpuAc01L4Jz8OoUcBrnuM
6wFtPa+v8p9zdBTF2mX+vlpAYZzDqAnMaOgEQ5NJRyU=
`protect END_PROTECTED
