`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gk7Ad/1DJh7gr97gVhNLeUqDcGUPLs4AZwKq1Ih0saq8ZB9s2szcegZtWUj/l9iC
07ZS4ay7MnD5EPVvvvJoXtdFqCr2pOx0hpcZxjd0yVta5DQVbnWmfaxF8BU2Cvjc
1/OSIh2diD7FNY9IBfB4IyCGKHRqhLdPhkm6U2Syk0ZOv7+RoMR6LUc6CaAi6xQV
/oKQLVrDSRbZ6HPXI5RqEsrXkzspJBclg945M+8JfG9A1brs84qNhFUa0xyPwy3C
6issxhpsSkaueFG2fVe3/OlYBjM+m8GvLYjwU6G+lcXI9QF7QUpJdMBOrRqaOkDy
qO6Pwm9ADnjzEYYfMzNcc5Nh7ys/xQCUUImmMaoBPLFgVsW7u75gNxCEOXnWYjuL
7Yya6SR7TSciUEBSBIQpAYD0/g7TpW9lIW5QG7cC7Q/yQKKZQIorxG4rmX0K/SFw
O/xzlFuiC0TtuErT8XIHrPrY+/zzp3Vrh+bJxHHLOZ46J2FYjZmK4rdm68RSGnxl
oBE+Q6ZSi5K5lv1MmvuaFqOA7kRXjj2NwQ2NxzXjfBbbpJ3R24ie3KzOD7FyzKX6
mrUTfaSikdILq7YNjYAxShxfNqGFiUFW3wyMkqUGdURlUa9MtHo/kMJrzD1bCm2c
0gFvsT++jcL7+z4Cqpp+Fo3czWnppWi1EkdFk/luJ2uiK0MiIQNxWISGtLr3X+BP
Y3Lk1kooPpeBEKSdW4dZDX0e3GSTFwbsiRoWdh4TLjFUPz5US2da7c0XFdimmXcY
VCuhMiFgWX+yib9itjbDmhPu5syXXwTUr+M3Euo3VaJ9c/r/0fUD/qKB/5IUkxEK
V/cgLf7+PZbcMpt9OIzhNNUiUJD0Wx5s7aAJmsxrXYvBmlUP/qOioGLpELXNrzBU
pOHZYgjXY/vrdO4NI3uJSEZg8NVQM2l+TuebeJb5FVqV8YLEpRsQII5bNMrDDFHV
Xy6X0FAFGh7aBFdQS/0zx9LZnfvdb7EJgqJ23t7ZhiyuhZ/nIvw+k8BpAB5edsin
6Gbc7VGgQ0opDK//YChJEJmDS5pwl03OeLh2JWYmA1vT71nXEyH5q4ga+OvpmhEM
ZVPhxZNAqube4zCTYojgfCR4We/viYalU+1SHoXcdLNQee6HQEsJ6J9R/VjMk8Ys
tQs2IGaUhOZE3ITT9w3f8X0Y7IK/cRcTE3NjBdhUZ8oCE3KiqvMgEq8AvC0yEx2s
M+kOQ8sjAEuVuFMD5lGjwnxRkT9rMVkYnLWCjxtdzG4gqU+k24tOS/GBrR5+2q3z
`protect END_PROTECTED
