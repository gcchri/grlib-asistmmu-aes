`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yx7qXhOyEAcguJKcNoOEsfOjbHjytvnW4ov4lyNUBJK+VeDwJXxsgt/JZ+La7Mar
6YCXEKuMIV+oOaeCAlcjxg28Q/KxnhnGmiTZxupaLRmGCbEU9vYKcF9y+uVZqrBE
J/mAOwnK/+Wvjot8pxD3gR9JQdZIc1gMAvB6+2GPZzsfYmKAexg86Sz3fGj7Vdl3
ubUcyk0XndimJsqvIIzTDrB5LPSMhH86wN84cRS8mBhG4sKx5gQVKm4MvG0vrZdy
9NP7MY1RKm0m+qd6J/ZSNL/cdPILr9Sr6exTnOMmXpLdxPVFP3V2pFBUbKG4ewBG
nkDVcwa+zJa8FiiL7yA6sL5P5QeQsJ4vWL7OVfvXJrdfC+IsVp665ISyvXBu7M4k
QPKEafXWcj7Dngun0wbp0iBLGvKeoJDDoatfz2nDqiYnQph442uZWlwsj3zY91dP
P70lE/CDIQ/h35ONZ90hzx+AP3MI93agedXEh0qNYy/beRfO2eA+NXSobBcs6K24
tv9+J/4hiU3Cn0zh32ElDs5+CGehBHJG7QBIvYQiPzCoDQkusSc4mRCmD6Qw+qbo
A2lG9/L78uFIIVOv0YcRfvw19hLuor00/Onu2oKjbTJIA+KMIa/WiMiKulzl29ms
Iml5LkePrDT/7F4F7HEnhfRRKqRgql66eltkE4GJ2hYrthDdN1iNWC4n3yBH+bZ3
i3H7jHUJj3dVDarXLqszWBAExmNXi8VkremSLQZe2rsBOXSLPiVlOofRa9nmg7ij
ByUlxdlOvZdmkzBQjiamVWQp9KIYKTFuA+NZet7+naMEVcxefa5hENjdwSdr3zIa
7i6fRH8OANshL/GT6Jw8mWc35EvjU5tkZPy5MUE08+qDlIHV3sUff4aUbYkVkj7o
1cETcjYO2t6CsWMcfsAaaHLf8PcJo0NXnlxUqM+I9bFp8FSd0Pewg4mLjWPXOR+3
3mHYMvB2Yz6MIqZBRhgM9g==
`protect END_PROTECTED
