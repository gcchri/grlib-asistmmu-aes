`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Fcx9EIj3rDqhS1XJaLme6M1sajfb6ztFIZ4IeGHWWb1eSaK4kvihEkuJRYt60xi
v6zwqBLFZl5Q+0bVzLX4S2pAL94IsFrt4z2Z6RDllw4BX1IrLR3jtGxKBLlZgYWG
pHTn+Nq/gICiqWaCTs+xdvBizfwbVd6f88CFthwgOvudd+qaiJOaMfnTTLBpHreW
tHkGbtQkW7BWwcI53m/S7BzhKlHCTKKcSZMgAT5r4SB5Dy/G+jbMfZbWeLbMLIEt
ajB8kbi5JK3Zs/X/bmZVuwQBqwwT/BVJJPfTe057rkqVldIi5xTDRK0WWYj7Gjeu
BhScI7MdX+sAmGD8Y5hFiqZulUFu0NtV3wPv1r7sXydtlgvZ/LVhmgpwu7mLVYY6
W8j9Xx9ik3c5PpneKpDPVQcs9xsCE/BAsF3oYakUVfj5Z9eDM8iSZWpVpvkd08KR
po68P5lZayvD/mHj1GG8bJVDMIn4ijVJ/ntzdr0MWbRllnNuMOd3ZqGSR9lF4MY4
+WgL+GLu6nuLHdjZP06AsuDsQ7zr3SJp3qi2HIk7WppkfojwhpAwLv9Cxa7OaJEn
Q9F5XkHqKc3hdVxn1RemRuGdye+R9DdrGBYzEOvp96/fl1xpaOuQPG56MWid78UR
PxoKWQV3P/TLIjLVFUBH4Ij19I88QPCOi5/E63HtYMPMBl706F7MZEP0Q7NVhuOb
p8Yrj7G4l/36FsjUcl4mdj3rkp4luznp9lMMEkCGanesvAjLc7+lKMoYy0aS9Drs
hD9b0qBDSAMuvIZUhGSwV2RJSlggfqDZlsdNNDYmwZhP31tJrBtz6d9k7oqpOasL
P2pxhIBVEzoVM+eQNJl6RfEdPtA+fBr1r1Fcasgn8ObNQTdgybS/vwJe4pEk1Ott
6wOpqQ/KL0g2e+FTgSpEEw==
`protect END_PROTECTED
