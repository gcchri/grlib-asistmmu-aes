`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gqUAum0r6HnvchIKLGA6wRqIOkaLm9GzXv3LVPZ1udax5Op3Gm0SIS1ZsWxLSd9H
bU+7h8+cRYmoWpCu+tT3V22x/cjbSYe6+bDFSSOqnfGTcRUDK6L5tpkIPoNTvr/j
mHI7BWGVCcd/I4J93HBHQyX47j5Fjs63gkp6VPPTaHVzwJku0QmhnM47AHD9Lkma
D5CqGjqYX36SMrQ+AxPjvB126HbcO9NwbQyAHb5bYPHaM2SiXIxujdb8ti+F63Gf
dxEunpoqzN80Rc7h234C0Gq97HdVzqBmaRJ7TzqN3KpFBsU4gLYj09IMF9QeZis5
r0VIwxjKOBivHg+M7RaskLj+Uw3I34PHdJ25pAbp6Sw9zn5eQszTnwkqRI+ZWG23
RwOt3QgYAMO9MpmEAecksKN1R1CTJWuijTcHu8vcxLvH7iFTt4Dki9cCPHNCGcDe
`protect END_PROTECTED
