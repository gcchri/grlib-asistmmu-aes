`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Q+7BjCjo9LGeSvEKeTf4fP+CNOXdLRd0XwuxvKqAIB0OOLskmb5Wa//7sMZijF1
KYRECCON1StAortELBCc/03HVSfHghMcrTCEbco0X8ZfJUmMKYoRX6c56W49Sgo3
Z2O5FJVqLR5E3fnpaRq+JnLYMfMYNBezt7WehSwXz9mmRT5BClRPtd4UfLbTZvFx
AvvclQBxRpA3Pra8Pv67nVBetanEswy08Ax7MRLP0FDNKLh97Crnmjx37HX0YyET
e6yp4x0W2bu/puwU6EG12vud8gx+9v6pOTQtwvYAjVfqhvqvhofT4F0H82W4sNdB
p9F9GngtOGXbosE40yRVGw==
`protect END_PROTECTED
