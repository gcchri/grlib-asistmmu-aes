`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DosRVzIu6w7mf9CT8MHAVVd+ID48diPR/EoG/D2RuiJ6lnQmnv8Tg1ONPEi3UXTE
2lLcwnE758LTqOYO7XBda1ldn4M3eMF8Fn9iepxI/yTkHu06Osvf6QN/813xHfWG
GsWNxI8A6pnrEIozYS/+EUbUfoao7UebKO5EwMRDww/opHtodDTaOKeSjQBFDcJx
y7EdlDi2n5LjcSxQkwnQl+fu7qbr93yF22WamI+/Ms1I8sRV2vfIGQSm6maqjE9N
54FpDbvLLyHsgrqfT5V10FCScPNYv83NLZ2LxpM1uXvcMaQ+MZqyAV9wQ58tXpZg
p2slfjtaCwSKxbx7kN0Qtp+s9Fq/LsTlgifkFcxoMGkW7ADk+Wzrnn5/+Dm18Oa9
tEHEGPHQcn0fO7OKr5RB/HTA5icKcCFggYapb0zaMFYvObOG7SAAiZJF/YLJaPkh
8MyJuZ9JkzVsjwHVBQnSmY/jB1USuQuY17OsitqOOk/qXQmQ+dGc56TtrrtyCBKD
M5EgFxqVd1ZTnLdViK3ng/PjAJm9ojRGN+YMaByYJRkhRW8p11HS6IS55suyvNkk
DzBTfF6HT9+0o5pDlY6/UnbtJyWyDFbFO2E4O2E9eOo=
`protect END_PROTECTED
