`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C2Ln0zowUeQ9mo66TbaCETodjp0/0MJJ96ZyEALnVoS+sXHLlHMOaLZek0tFyWO/
12ADv9VPZZ6X1Lx1vAhgGNYkQv+5fRDTiGs01DHMlvZ2Gn0CM8gfcv0zY9VBiI3w
ZQtxdo8Tr1RGyL04on+JXQfY86F4XD9hbBsxomalogAutLdhIO7vHNbw9xchjUXR
F3o/jv2DfyIF8eaFetlFRGyk0BvUlGkLrqyx2W7RdQ0A9dPkxPmVsnRvE5jEqQ/o
0daoDl8esJVTYZ7nllb7ZA==
`protect END_PROTECTED
