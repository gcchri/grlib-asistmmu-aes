`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ZzmJLY/1qGAfMAGxzTg26xjoHViR5TyKWn91jpw0rdi2K7NmNJvQSlIYaEkugOk
xdk2+SbDaa6XKrClxK1ak1HPyzoIcdrgS8vrJzlwZWCCN9xojeIl4KIERolF1UcT
1RNZuq5J9H+Gqrd3wj0GHza75KScpw1lsl9nnX8cWp91i4VGfxZTRerLC7fUTTSq
6188oiBDtn0mvcKYHadr8Fs/vy4GgKwH1JS2+JO5U2WycEt3nSy/Unvyq92HXfAM
vTtIAwt4y4SUHNFjneLJqL/l6gCrrJnQbRy/jFLL1v5U4MzMwMwHyyrti6B9f++x
Fjh4L8PQez2/1FIA+2zMmKSwYjocGT+B2TA+vI3ol2S/snBa1UYq+S8cJdbl5tEY
GS2eBzGBnt3A+jxTOx3s9iE20j2A/ZNkgDP/Krt/94DOTA8rIy/MNQ4fJpE5AQmg
j8oRHzUhKyEAW7HTidx+PqVfhkRSilYHyqshpb8amD4DbrHZET26AMoj/DXZC0Yv
b/FLtoZai2jTwIYUjt3RyX+YZlObzCgcUUpN9/DHwSTNnTfNHHBRUqbVYNrYeCNV
LJ6AGLy8llSj48vxeYNTYV+NG2Dl5BaV6YvZoutXrKb9m6ZmGJ6Rw5yHGErqrQPm
wa+UVaXuvcEryj+K0JKbGg==
`protect END_PROTECTED
