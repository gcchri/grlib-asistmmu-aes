`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OuP4ocjp4tMTynm4kOKC9INH582Ge9VGWKoQ+HQQfK0iEOerz8xPGHd/Ia5urSUo
tUNb81LX8BoLZBS4QRMrQsceWlb/9/TdSGYWzCXoIKlq/5Ph9xTfeOjXjTplTm7T
rwtwnw8nnMV/Vc/kD+FyMv8sM8hgUII5Q1lu73NM7aT/Wu9XTk5UME0aR2l+6psX
I7kh6XfGRiPxNtsnT6pXtdlbJovEb0o7qPVbvqcTA8GiQsZTGFED1lFq3S3xnj1u
3EJqfcxKHkKM+xLnwiqcn6IJSjdA7+RybbhkUvF0FSMPJGaAkwTDtk9u6IDD65pu
9aHIIpkGzW0HNPvDhk0WcKMo2yHwy9R+pIW6mAcYn9AB3mqe1MAjLcBX4a3d2cNs
+1Y8FDWyRq/ON6Q+byDbSN3SFV08cjqyIhfbxXB5uXWziAOnfNzxhmnVr9EkzC4v
/oUhxQAKJ1pQRz/O5sdyFJRnzUyCO+lufWyLT7uUfMbOjsb8xzj3FzGTbLj0Zptm
oqmGHcvqNexYcRrb1kOqnTqhnnynQptJQzx38inRyb1VhdcIDQUwdKIHMS9zD2t/
aB9SAQXEhWQ1nVVerMAmQAQqyOKpq+JwSlQyE0PdlfMDxd/sVpM24rzYvmZuOZ2A
voUN0Zjw05vB+UgaPWZ8aIqLwn6XA8YXstf12HkfgcXm4mpxEUG4eEyMbA/lPBr0
cHSukOIDrnYLiAbH91UeD6xybx8vKPg1xzhNzAQsQ3NXgky9bzp36GDt3SuJVoiz
UHiTwtE+zhxI/53XrF9MOn+MQavf6EzvlWHdEiXOakvHCKszesrRLOgK5nUp4Pks
NoCv0j2dVDYaHK9IPz6bqklnfGOy9lXDFuqZG8d/HMA8YOMTddS89N3ORxZhMUN6
DYHHeN5WZZQEKE6/DRpamVN0h5U08vNymwq8vvu5noQzSuAnOpnjfcel5VPLKhZ7
R7BXGzbyXswhh71xXxvRiAmvFYmafrOJ4K93vC6x1OkmN/SjzlDnTM6rWc6rxySd
8XfcomMkPx9Fpl486yX3SQxWqdhINZzYnZ0GurZCs8mOU3hZ0TuD0wGERPb+cGyc
ZY2T0kPVzQ146eQTEGDnQwxDZu6ZdRA2mVV8UOIv4xJ3rUuJ5wOlPZmdJpduFyjk
nK84W2nNG02lIWMNk2UdkDTq5BeOW0fq9kWn7N/efY+B1m7Xm3BsjJFDFIsggXnJ
tcI0ldPtInpXyBbzTdKnBnrF1umJZhJSnLqQ+M7jeBUYYfmsihHcB6tJHkQssqnS
KHRvIhy2eCL15E+bl71z+WhWt2Bv0yUFvTKTDTfU88GfbV1XlKN31bUAXptdvDkV
nw7UdEWUwy0GFNuNxQluA/MZhJI516EXJanleSi0juljrzxUb1ykhsvm7JxjwWvP
`protect END_PROTECTED
