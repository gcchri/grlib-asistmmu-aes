`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YW6B/ww+dQ8vbwuumgQPS6VpD5Kw5VcvCUApr3deYX0h0nk1EnEogfv5nme8ejL4
NS3WrqiTcimy8jbGsYC0SwIadQlHQqSShbpKutX2sK3wT38LMjCRojZsfTLqHnDY
N+/hxaChzDx3z6zjagjRf962tNa0vERf6K30I803ZnLqIPxi9PbHvO88STg0gtza
jB/GEs7qDsrWQyVROPqhTK7lJxhkZ+qNDpJF3n67JI6UKt9XB0eVjZx5dIU/Ekvr
Lq+6BiGC7E4eMr74ggMBFlMLDjYcJVNG2meOYvmlYNfodl0eBzBaFEHC4N3pAaA9
s0pCcNLIP/j9rY1+/2iUEmwtB5pyYj2WAVsMut+Z76kojLNRd/j5ou8hYL5vls9A
LTHA4yTyar3J3eDYdAnXW/08j7ng/ehg94qnZQspy9rFDQOAwVPPgG4UWlkLlhP9
xsv4fE1QJQqtYiQh9X/Ejp7Omq2FVKrzXPG7Ye5w6qAkiDc/Ri0dz2kLjUGsDSqA
7MT3sRRMisQ3WqomY9JqhDXQaEaMawRRskOnuP/4emuVqc3Z1hM9ohcOjdwK72YN
sG4AiGfLLvUv1aXDSqvdPEaNtvmo2nWnHMUg9TjT38fGNpVdqyrQZEc5wguXOTPO
2Ksnmc8ymAe3D6fR9TOPjrzBC1r+b7xFypqWwkONO5f0ct64mfZbBojCmLDv75tK
1oU8fgsXvefuA4FsJeOLmQVjZ8PnLKwzzO93pSk3k9I=
`protect END_PROTECTED
