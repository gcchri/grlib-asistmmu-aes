`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+px1n8ZgkiOGtVC76aILjZFuu5dS7AUUKdbxJ0FQ5PgS5PQoFWZU0GEVVqPPZ59/
aC6gm0Z7x79yQVj8P+xd4jJBM/XdFgSD5EJbqoVYV7ApoIl4jg8BmYWfGCYh8zhF
9tw+xMpxD/VUEOlF7DYLSDDvCB2GtduBntlRM/k65ZbZ+xm9NmNQBPieewUR/e3d
GOw1YlaPc/Fx0xXATYEj/fcZE0MQ2BHI/TWWQ7Nw7RQoD1KcDGggFM0rXQQSH1VT
GUnhb06Ok5ORN25yOUdE1BdmOlG01DatfCZKjGV3NjOC85YXHwL3DHJvh+jEr50C
TwuUMXUWeSbQkqqz+e6ZjpV1Nrb/yJIQwTSEW2KXvUsPoyiR0lJwYIak7Ul6AbuJ
3m2wp1ROMyE/r+QhuCMPSQ==
`protect END_PROTECTED
