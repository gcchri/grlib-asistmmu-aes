`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DxGTtcverdMKYvmqNkJG0sDapTyWbPdBnIQP7n0AVuMGQlNVtEb6f+5FhXdq5Hxs
n16CgKw7jfC4YngvPI1GD11r+UXPJhKzc/3wgM5/9G38EiKqD0pszjzlKcGIneOZ
C+BCAXFl1zHFjat9kbGwQuYdfrT96lZZvDlSf3kM7y1HsdJAMMGQKIkJPNzG3iSV
OeIU0u8rrGuzgfOHFpPNRjJxrhTe8jS+6B28hqRvd2kQhrxyJmrN4ufeWnCS3oQE
zY/DWTwzhGev1HmfU/kBsVH+2VBJIq/A4rtM4bVRw7gUOg7kHGAj+CarKPN2HTcu
57mI3RZxZY0m9IKHJyl5vd7GYN7JqIxmFWkS9vXnXbl7BUYbpbgSPUF7EfwhA7UE
2cATWCgfeKkU7hA1c0UO0tokBZdvQ2nllFE89mTNLwIVeUQ7o34wJYOTErvRLPFl
BbGB4nnUrVx5y33dGZlzorVkZDw7SNzel2cRj9kjznS7g6/9oASQLY45SFw4PuTA
r4+nivUBIZRdpQo9RWQ/La2jVKG1JpEJudKDI7faKzARmH8DCiD+REQo1KIGpM2U
M6sXR/mUyropYZqA/e8L35d0dJD03HXwX5XSLB6BvgPiE4J7Hbf2mSocLYKPR8mI
ZDxNxL5+CLx2w/YrD8/+YuZnDdyuHWYeWmgaUpAzNk07uWA/mcoMYagbbNh0X2GV
8XaMvMN1R5+ExJLFJ0W6/jsUH+tsdr15RCNRVUC7BiN2h+3CZr22fXNt+k+UlPYQ
WHfLB/yKUKKai1Dh8k8ZIQsew8gpfxSGDpVuytn1xIGz5z5JeccXjAsSEawQKX48
Ab83XrUXFRTZmPDTRbbdqX1TYpsdAx9j+JahpRENXBEUwKxNWr8rGEhiC5zqeO2g
mC5XfiD5RheoLwffWGbBrHpmO0Q0BNA7nyucaDgKVilxYRYpxFrQc1DqHH68E0fO
fUkb5QSud/wuWA+U2N5VCWDEh1XytCLbXwv/frPLNIFkU1DxKOP/ikKiHAhxQXoc
kJMmATXLon/kr81zhjerVSeHW9SHm19veTPdz9nRqWip5/4ffhLqVpwMf7QnMj2k
dPZi3WSNbY1/ThmQvKeiEYG+V0whM72Mm8IhGXNLtHqRWHkrR9XRo0ACOZs7TUIN
HUv9iBLnE0ZFjHT34H+H6u7Z9ZULd0YW9P0mC8IINCbVBRRYxK9+ADvmUeEzzmlU
cvQ92vjOv+Jb3ldxuTIMZwki0CPrPmtWgTY3wZRCuLyu5589NMZUEereM4Olya2b
leLslY3LUoK+lZcMiTxVGlLzDs1BMIzraFivSu4Xs2GuxUfsRC6cNwkd/QxvwUQW
Nsz8kA7iK7TUNzCbkvAoGsiG4v7S7ZVgDAqfCtlFRliQ3Gv+d6eRN44XiQ8A2Yy8
3cx/W4EcomAAEoQAZCKu3xKcr33KbeFfcpexl65bDFIkjUpbS2EkDFOwX/NVE1tE
EsnygyWSxLk16KKFxqVlFfbILVV8ccwMhU6hQYWovETv0Lz7NA5sac/uK7QwMqan
aGPnhVb+mRIFCJmxhhWiIMLxC8zic/4G0FJ/ZA1Og2kBxbtHIP4kLplkdNdYllIq
lgXewdXjel/W2bKpDs+8F3GJBVlfO3FHzzM3PjJxqmG/FQbmhdWOX8lOUinhYYcw
F8mTqdMah3yjeb2JrEJ3Dl3TieqZj90EYrpnIi0p+LrT0vCE2SKmYXIu9T1wTLdq
0Ec+HHT/+UmlwMeVlpnkG3PjJ3IVReCzCqg1lSNGPZJCNO45Kyz0EgXa9iee/Xz2
UIxsdG34565ehRHF5LsmQ9bdeeSwjxlSb8PE1GEO1d3vczdqU7EU0c029eSUZQZA
SeliGBHLvz7O+VmLDHgqwru1KmhNXTcR2hNDAT6x0ooZj9dki9oVrpIg0kDuRGI+
KcPLv3ZzM7mYIYS1tB1o1DGD1MZeKUfY5Pz+6DH0phVX22KTW+3zy2tM70SRubmW
mY9+1zBhYR2WMrQfKdaO9w==
`protect END_PROTECTED
