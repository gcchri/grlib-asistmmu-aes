`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qu2V91BBoV+hO31QJPB++DpY1d+vYbryyhQFlBIZLWonvS/5AEeaoH78U618XN+P
n+faMwW/CIJ2kroPpMmVTjjkAzzVcmrLNjt/r2MAhN0vah3x9+a/A9Kwe3pKCn3f
AYUGAMUSE4iHwOiGXBmsiw==
`protect END_PROTECTED
