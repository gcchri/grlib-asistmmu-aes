`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m7U3oZ+Lc4pvO7nDU6C7QG3RYEKCktvNyTRpinh8dFtFaiLH2d/OpVMtcjSZoCO/
2vXSnt499mgQd49inLcIAh2wWFU5Wccei/jFbBnxMFZ639E178plKjg0qu6Eflgt
A7+2pq4BPaqvP8RdI5W1ohxhA3M8UkqDLJsLwEGgOWoNsIASjk9rIfYLtrUR32kD
VwiB5bv3OZrEC0B3bAhoafPZdcWwmP4J+GzK9oWagYKVPESMnHicMIuUUD4REfNa
8Nllovwn8cgsQJrPa6d+f1sEmy/ryl++fh8zOtMhQB3vum66L8jZJy5wxuutedfw
jBHm3Bq3SeFujrF7ZjsegM7wZp6ThXYGQiIUJ/AEEAVxSTWnPw1ziC8SVl/hcyok
z6Uf0tnlrtEU84DSowd0duZcd2UkPGe2L1p5U/TX/p6aj8IrQfIY+TMXBS+YYFio
`protect END_PROTECTED
