`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6N8dut6Whz2SdklNf3QIY30YdI3DM99hESm0MnJRyHAcCkze0N27K+10TVBUpX81
wfs+eRv6G4X2RO/CtQUuICKTID+v2aeyKsuRhz0P5L+iZDjoYSNuzJVkhVi2SwBq
vrHr4BTNWmUidKgrU1s5pIEFq3L2huTNwYZRvAnhDCHbdxpQtT9/Ql1QvZ3TovKZ
ojUDv9LjzqFrVXw4llbG4BchGND3q7evKHb8jvZw/llcGxaZE7VpL1N81S6tQtjz
WQqoXB0BUD4k94xIvhj+gfVvpGARE4eZQMw9WD0KOuMTqfiipbvv5HL3kcsNDM4S
xbJbVbqHj95g4+sNSgAOwA73zvEGIR3lEFZVmBMgE1dpQLy5VFbjOjvmfPEASuGd
nkPDE/61sO4CGiowVu3ANXCFtLxHEA22nMBrvJNxgqQzsAIFgTynRMSEy7nti06E
1yAN5ixUGlffC1oa1TPFUcAsLvVX8FCf45BYpnH7UbwJf/XXL+nWcblD6VAAMnpb
g015HBxtOnpWLTPswmd2NOIro+SxrI9xsZTJjjmnbgu2SgjD/hJcGwbvQvWqCDiP
lkf605ZPfexq5rctADGa+4Nw7MXGSvv5l65EemunqZke6XXGiDrJcnMEOYvZNC6D
XDToZ/Sr1Tyg0FAipPOW9c53fmt88zGH/gAIpliwh9e/6ZuvGnHnSsNK1dyT2BBS
0lz/FRMdB9hWZktH3x9nlT8Blg3B/N21KH0OD8i0k5u0u84zLdoHWB9W1Gc7bcxa
84qO263r4/0umS3qId6/hu2k58dewHySb9ksEXQf0XmTOrNnbpmfuMiQapFD3RYS
3BknvQW67tI6bsrxXWs6hY4rxw9Y7Jh1f4L6ieXBNFf1nb/Ga4V54rpQI4+ATjWS
nG0ozhyucHM8l1ciMPc1hynat18cRM6PcR2msg7331Nfg/+GFoI8Ix2gh0DzJRKK
XXlTm223/dk+ghSmgBmZhgRCmg7fIEzbvvt/oWaStQOhbJzliT+dJqeHe45x0WsS
8/MbX/wEyQnq8p1rlX6XdgehhdqAMWGjWtrOL7F60my8wR8gHu4B+2UMjilhXg5e
fPysFSBW+VTNDySgQk24MhMjj2cQzK5AO3n3Q90DqDSfvOXwn6hFE2M4y+0QdoRc
TOnE61SmAtq/pinfG920f6J/0X1Cg+E1e62M3IHc8RSQs0M6o8KhzP/2aGlDxNk6
jPpuRVQPMy/yuBSCe5GYkEVoKvFgeQ4h5XBWS8D2BLnvkPbiPUsvecGc+uYHjsth
s0K2e3mDt/mRrNqz31+MjnlSj5SsgN23ojzbJWXbRaO9xEEqmZPqLp2WhXCuyqA8
`protect END_PROTECTED
