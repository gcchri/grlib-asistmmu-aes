`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1pdD5b9AGwcNFYII34baNR7IoQ0MzawKAfIgKcNIpviSHfRfTTUPgbMv5yo//3LG
/499IrIjJ9vi0Kdt8E4zZC9O/RVOrUoOfQVEerDwN/lqjaUgX5Or8ole99YSWnLp
+GITJJK/aB5LGJo2vMhtdtEEB3+am4aQvC3Vh0yL8v0LVSFbZz5xdaKoKl4fCkX0
0SJfRZwJaXkXesVju9TrgKW96ZFPrT+UNZFBXP7OVrnMaHpZL79mE8GuwN2r02ok
QeO6ZE4dfLlgHiw0be0ulZZ+K4tuFKv5kwhmbssey4Y=
`protect END_PROTECTED
