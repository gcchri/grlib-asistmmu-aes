`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1G9QhoIa8J4YNApMHWKdEYC4+LvuVQOl/imQITtXJNyTujIvDT0SFYGVDArR/usZ
05QLZMEhEaUzXPR5jGVwP7cKZTuGYQgpACSKcPlS8v+Y4IB3Jb4pAFZkeiWwVqNu
CRHMJBbhlFw2myCjibbD4IqffAYZVZ7e5ALHxGumDMfweqiVj6QB3VMUNT+4cj1i
BVtTHM1YZZqyBotp8/a/d6n9tE59KPAvBYonxirGDDO/AqCRblI5lrKL7n/qXcRk
u7+KYKN9DhkXEMVVu5nUT10JBGQokzkFAeEW3hQqOAfi9hN3rxxpwoiuK8nf67EE
u5cb5jdPYe5bBAlUF0U4BDMIrsWQnP0mQrNfD1us0BWZTTtEVGCNRdxmRCyFNIW3
+FNScSNS/Do3wCq9DzArbAtQf065yvViaq4EgNG90aIgifrJHpogpA2x0xeupbv8
LVqV8KDLtiRhq41VJdGWu7h18pqxb66ZbXM6jF4E2gUgGpMNE9UI8K9FQfcTRRZh
TiHTzonuVsM/gJ/nKIWkZvYjXi5y9E72yPv0DaWoXtCRa7/7z1VVxPpnGXMgx+H5
YtS0oNQuEVjYI7MS+iDKMMXhwOOeolS7OiQIBOeIaZopa+Npq32tTqbQyGB+Mtjt
ZhdtweCkemN9g6ymxEF/pzzIR1khxIN7HIbvJdKv3ZQ6Qna2hLhuIwSdqkXmsKR4
HvMcV4iTH/AVqd2XDIHWtPhW6C9Qc5+H5rByxWKCI6T+2sZ5QdMofIcxT4dBtvIy
p+vq1ZPjzlHC11mjz5rijNvln43RUBMWy7NapVMhC/FsGaJXoX2R0pQjHUh8vYet
wTWaL1KerYG9oe83XkhncQkj4n/NEQDomj6ql+qL9/Rg0i2mXq7ZNzKA/C5km0U6
6PCaMlWDgt9Pf9lAoInKVpzmDmrD9LPxi7XJvZYvlfG3zRSCSY8Ft3Kjkl41mK2g
g4qZ915GD0nisdMcD3pSFCh5s7ud/3zWYQtITsQBeZi6RNLx1GUllFrhAyryTQQd
b9eZFg+NrZoXDGMKWI5hE8WU5IysYmHJ3G9osmKmCZukGpbMbLWgJwUnke2MwFaw
0zQTaA873yQp09Bhoip3hiIZEe239vWLLdD8YtkN5UX+tixSmknwvOH33GdPeS0W
I5JdsNPJ0AYpucTznvo0cPXI3LyxpFDMfpLpgk3H3yai3hNiD1JP5bIHWJ2LcNoM
jG9ZuO0gc/oLShQMYzB2U9xQp17poCQR6kPvaDaVLX/KJwWptWaXovdE+q5Es0+a
29acM0nzp9kYPaTZ2d0j8sGeAqtW+y0mlUu659AxWGC21TWcoRjtk5Q2WwsQBlr0
6JAAxTkWwJY51a1Z+oRLqMnpUfVOBn0wWF4iSvntELCWWPJmJVQmN3r45VP0S3Lr
aZIDn3DkXglS2kCktHM3/RcqIkoP24laYSOO57mu7YRdUHSU0XKkgTg8TjFixsie
NntmVu+SqvB3j11pllP8jeKQXqzUM+sRDJLaRkQb9iKJ9vyDqVETFJBiGrKutBb2
Pqh+5bqAYKbAZD7eVjpniAkhglUpn+mA+EuyFWiStdbUxHBa1G8cNqUyFXuznigo
ajsFvV9plT4w5ZWfd/6XJRtsKkTItYMQEO4tYCen4B0/9gSuqPC1Ct8Dd2gecXcm
WjxCunGOjziviImWe+0nrPfnCZ5HFC4tXTOVa5cLFd8/owa6yypS1j3u+9RXLXfY
1pzTkvFL2UWwunJwtN9ggrcUVJvDoSocP6ZRCgSx4cZVXk2FuIfV+3QCeXdcShLX
iOYs28UKUdQ8EtfVFqOyQ53iQeu3IG1Qp7ZNF8QJlEz/d4DDUv4mJW9X/D8BdptW
OBMsqFZCxwbAs3Lbep/gt2F8XdedhUWOGmxyDmniuZYDzBuVQb3CPKnc7QKrNxCB
6Ox/aDIIa3kwFC537VW3gYs3O0Cuu6oZPWfWOEaRhMWlNko6dy6AGegrNMOlBbuW
c6xqg2tBmYV65bnppfjcGlRTprOBv+Av3iYb/yqBYLzfxgaBFZ+DDqEkJ+J63A8s
Mn9h1KvOaD2Y6XGIFTACffmWsE4LA5kYfx3FmRIz4btUGhkI0peH208GYwnBumzd
vcbw3bMD5td5DTXx1yIDNIySUU7kS5kbZ+MNOa7y5LEjy7JDGqTcTmsLmGD6gMyM
Yf3/gFtZmllwxVwDds1YGJfsA4P/MwWJFNQW3J4REFHaoTiPOIuTQe25jCPx0J+J
KAq+2GOZxWWSeTkiPL+tI8u0XC4iU+ZKo8Q5TJnNfoYv47FqT3glw+yqTzL6CWIr
wojdUDhnUzJi2zJ0JY8UrEjiy6PQp6ZwIC+pnF1iGzohfChU8G2zKihkgU5abg3Q
+E3keXa7KDP0suQo42tnE81XqGvVtjYTVjZcKDGjMGPvbz3UA9HNY24npxNxk8rF
v1PmEIHt5lsyNVkjyP/ZXLd2QFXyOyLQ+OkW8IX+6BxG7zR5WYAelWl4k3eAq2JE
nTgiu1W59HtOeGNeklXoFUdvb7nkmUjnp6oLpdBqcgBm3LOsiFTrb3RBfMWBWKGg
y1LbQMJGdvpRKQEMiTBy91WzsGWfZqP4zK0SagRGHYheKRac6c8IHgFFTb+X/DJo
GS2slAqxKIMVZRMekZ5gkXLUF1GiCyvWOIihmukXuXs=
`protect END_PROTECTED
