`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VMduRtHJNlVrswjUI1q7M10Fzic/GqxL7tX3wAqnmaq/3T8LvjCTOeorD+3enN96
Sb3yHb/wGRbittehWena5v+7g4LHiJY98g3OhuFLZd6exj1m+bFxnskPb45Qo0tZ
wUAMmZihOiaEDl8zZtShWjpVPH/ZxRNzOWG52i5FczVeoROPo4BXBgniZXkydc97
LyMlnK9RvhVxLmQ1ZxUbbG7aAezoELq13o/ks8VDjDxfLwF/9Mo3qkF2oQCJsaRM
h+sTQJkj6K2EehoA0xayJcYMsXsvRc800BaBQT0vEVZA/omecqWSrGjT1fQj2JQL
kXlqLlOHoFPTBNGv2eWQm3dnFgCwsRG8chxQ/FaNwKMYDmrGlFX4XRsCLxuf/2x2
WULVJ2Ron0TQ7/aFThF9S5trrFDSsQELUFB4cceRW/YHsvX7szWnLbdB/1XxVjp8
LS6fBsmVOAjZwQHpvHTRfmzxy+dnEQnZHqQbqCD/8ibjs8r/lSMhyiIihlc0Tsln
I7BO3Zu84JX8WPwiTz0W5I0xkBEWdBjLSwtY4aneNvrBccRfMtikBAmTEwdsv9vM
PVLA0+aFwGIGTgxhDFOKbBmEJSHQXJHGjcpTuH/DmTKuH5QJ/Wkzs/Ls8+HlNIl4
VAp4Fqi3rLTX3WAaVQRJEtIjBrQfEo1kxDPd3tZhSbp7Jf0I6DeNqPYPMF5cM3Jt
ISPG2TUhGztJuuC1UmUNZbV8ZgmEhnTIZBCGkAHI6wY=
`protect END_PROTECTED
