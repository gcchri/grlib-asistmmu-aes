`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9tIcmoNireMSYXKg6Z8n2ubgEvrFtQ+GfNYn5jX3d/GEZdfJblVGdhaRR2lh0/KV
DNB4Clbn+QCMRay+Pg95FZ1eUuCfqGqsY4Kx+rUJwKpplUf4BrSfxQhoZm2g2utT
hHHJGfNBeERLlGjG6lhAy+3/ka9eK9R5wMPGS/gUAXoEhbFkDqfVCy7S/hUw3h6R
RQ9O0a+DARUpsnkcA4tZK+4nUVYoFe16b0HyPWgV+wHMD9T1lmg36f6xNxJ/BSRJ
bzpgJqNKCvPcKWRv9Hn1CQ==
`protect END_PROTECTED
