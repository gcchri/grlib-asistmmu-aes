`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9FY8DO5/r9WnD9XOkPyU5gBKdne5JNNx6gEd5zlYXuKwyK+iwQ2tVXnzkZlsMmaP
39Ufwj3fHRz4SYaddU6xF14PKElSilLWxsnA9Uvk7nC9eogsX0sYufM0918kVM21
1DM3HCsOhz2KelZkmicBT2VDw2KbBKofY/3EZhsYpNkZGTNNAzVV6FhOp14wojd+
oND1UiXP4dM59XwKgvrmsVeqYqWEjeyrJuO3sDtC6M+rt3i/bztM5+v1l5tn2Iy/
1SaXjknbWqQobZgVXXbpX8yyoJX12bL/3nMACq1w6RBzoFanceZyJS7HRlEYquoE
ptDhtzgEQVbmdYCajjYaxNSq7Te9Pcl1lS+5FKhaG1tkSJQF1WituAQAIAWuvhOK
`protect END_PROTECTED
