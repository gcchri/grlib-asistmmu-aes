`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HodfHpCX2yxUCbM0wCCFRRw0mPFKuGx9SfkQfuyln58AHISLTqWQITP6z4zavCu+
y7oq8lbY4DrlTi7n4AsuurleYxHEnQcyEDKEQPSmqGsS2c2m8BAMnTNiOuvZh2i5
jj7Qy0A5N8Mvc62MxYXdFs/jKSfSJYQQ8WgKCKTSaT6thkyTL5JqtfZ6vQzTjO8Z
eENnzCSbgh7ZX/OSvBya9uw3GnA2JryZvzSeYb5tGCXuNhyiWgF1WETke0GUNQgY
MTyQLBQzF9dziSZGgsS+b4H0J4L/B4A3/rT5/ZnMwoMrq6ERQ4eaZ9jsV2EgFLCM
F0rZhkNXlLmzvPJ/ECoPxdrY9AEKhj2zaOR57wnPrYUzbnoNleVYXtAviVuFlhss
GCRjF+kf9jIPhAb23xZ2AvKkfDkvUzRqO9hhCfD31+08423HVfFvigOIUJsJSljv
rqitam0qZlf1BoG0+MH20QsIDOz4hSPNNisIT0RNCR+e8/g6SQ3NBZ6o8e9hPYms
v0oP3z+PuXeoY+S9+h1CkoyzQ/+G8Pxfuz6WXb09ne9ZSqrnK/BspU/jv6FcnTvg
Qbzc6hxPzZyVcINlwMDGAqr3bsFaEIytwifjbe90p+vbAl6wwDq2NR5rnSIzZbEg
y8+i+BzGhyPJopiilXGYMxdj9WhvUim32oY7EMUii2X8qonqZCsQjc1h6pUbtkQX
r1u8ANef0ofGgV8DuLwz/4mEfRMGiZZXiniEmE8V+qaf9J2vIz9gqrrRhP3rWj3h
K1TYjngxTytHqdoJ4uCH5Hm/FUQFBoeV7nA5rLwaLebhjMSOffz05rLVa/lnJrUo
Q7ZSW83FFqjg9iGT70iiGYzjY+fTy+ZlvqT7T06GvumgCgELLPCX/X83Y/rJzSIL
3kTqmUBP6pSnPhbIskk5N3zacqYUjssE1np5UGdzsPQ=
`protect END_PROTECTED
