`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4gjaQzgPx89mJdoBFyFT7beyCV3Wbh+Qjww80E3kFzAYbwCPkw0jlL3NwbeM2uBk
+89aqCVIJO87bfLlNHaekn3/5x+9gEt+QFVRrw+t3AaQt+yckWbSP6sOdUqjAggM
WljLWEXdRCz0+aKj8yoLU4uwZVlbgkJOHb6e1mpt8/KSz/2VUY0j+zbIhY7GNssZ
Lqd+BuVvKdpRPmePuivXGlrq1w4sByxPs3PY8/iC7witAtNkmInNcxBnae97jZIz
ugRderCtStf1HWMxJvmVPG3hVxLNXk+hRg07HEJuVKpqGbYvyE+MgFYttUY62FWP
`protect END_PROTECTED
