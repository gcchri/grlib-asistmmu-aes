`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DLMqA/qmoy+nWJUaQD6UJoHsrrEOEmZIdhSEyA8XEU6fWadOUwzjoygILNvBEiF8
BpDvNRBvoFgkg9yzH9dku40sw7HpqK5aBxIqCkz/SAiZNLzk3BJS/okwgRMtSdDO
5rE5vaHaqg1mbtbXHx5smb48M/HTk7z9OOnLG/gMCMV8gZjgg9OO5gZdi6hoi8HO
c6EDSgv/vm2sB90ip2T49vqJVVjEWLfcLEeNNZDki8Esw3YlZBd2lazwgjk4/UdB
Ks4knxTIfb+MmrdJgktboV3d2Ph684Y4mLc4NjAAsZSF7KD9jNyAqyo4kQnDhno5
De9bj9/NF4+NT2ltRTIDNV7rHcDMRdq7oVq5IrEKXy0XoCj7MttCiGl9+7iUSpk5
ClpTHhYyoXbEzSwQR3PHy0rrG6F7r89/Mg0mEItBpb4HKRzjtJQSMDbhtmL1Vkzm
vjoDhczxR8mZdevPQXFLCnGvITTKR2O61ikyAL8Ta0n/aTK0n7XcbjZk/gXhfMX1
ufb4u/spIyuA8ULVa9Vr3V99PsBbviaHDSk2tuKvFwqWLvBI4TK4pWIYHIHuKKvo
mK4udHaZHSLVl3soRftz0tFt9e2MM8x4+g/PTGF3iW26nBVuRYJP6tzq+lZvWlQd
osJngPbwrIPwcgWb5m5vqqywqkroRALjF9nSvuOAFUTS6UyHnnDgeuKRNYWMbapE
dfWYu978gh8bQw4l8E0zklvypjvFjZKhuaOmi2xpRN9gkfl5EntOZk9wX2gVaCeT
qrayDHjt8dBHupLqWnAQXiX7/bCl8csA91PJ+GGt0zhkoVKkOhMbCt8izIY1L4Ij
szCgGVsOnBlMZ3AJwMDBB/T+kz0HOAgBtj9uy/shiK8gvXzDDbAUp8wDQd3AHmi4
MUCiHCVchTyLtmxpMSJbnz8vm5AIclkFmH0gJxWLZ3tUdv/qu1ugT3msKnr56G5m
gv5VLB3DxSh2D/sF1+i87PhgE69MwyFkDfY9ere8T0nfTkoJr/bwIoaEO39c5ViG
+c053YS6FhEZq3h8rAitg9ulB5T3l6RSrDwGDaTETE1jtvCnL04DcNOF7/dZGYO6
+zh3/ItwObaANhL+NfKzCAAc8VUI5oNPwXB/mAL1z+qfD6qeZWTvCjjX5DZLw1pM
6Hf7thNwLTtZniALBiY1+ChvoVqkpd+85xEHCp+dDXKTj5HDuYPke2yMPn/ar2Q2
j692ZPlIaJniLf6iQGJqDygERV5+Z7hof+nTldo5Hx32FPxsNYuZthSLFgQM3M90
EP6jd4Wzt4LX+CtxAXFoIje6EmKJG9nNvL7g4xvC8hI7pdcVqEdAlSa+1HL4qH/X
o3+VrSzAD3S9WeEtpj2cs/eGlw+mXcPdfjXESZo1IvLaP0+M1NI5B8XBegcYOeET
TIYYzTyniolwPKQO32/fa0fUePiWb+EYG6H4opUDnXnk7o0+P1/EJea4UdejNFXv
rQJkqqy7snaxc4DgejPUnmVxuJC1rAkn9XZLQIXu1X/aqWQu8iKtPRMBCf9kGEZN
U2PErBewx8ea7CpMjNJrSH4nBVQHU/mjpLwbX5NtfQ/+TN+xlTBsueNY3k1jWef0
cWKQUYC8PrXkwPpiwybajl3yP7IsbVgv8gTOIHMzSPVg3X89H1vJja0c5mRauYqI
NR3aTvETAEMs/MZWSooadER0PJ34lVANsbEm8k99RanCjtSak/jY3JUU7xyu9ac7
fX97X7GSQ0OzYLBNWxvy+quSH39gbnv2vwuzECJw0D94CJGWNcY0La0TWt91AnAL
OGJZf6iK53YEI1ffpdm+GCXUgpOHAn8k6GsKVAeM3ltivaBy+4j0QxYzxIBlpgzO
Z3Frphg7j94jlIsVgGYWcA68PNCnCP2k5ocaB2OmmwI=
`protect END_PROTECTED
