`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rqNDQG/8UTfahw/HywQ0mXEFP0XW4a/B+FjP8YMb0C1QHPSXIMuzWP1T6GvepOLJ
2i0BL3Y/sniuqiR+VMBDlf9CCc3QtivFQw0G8bv9Wn7VmWBkpaT4N1SIZivkCOg1
DtvuxwAS4XD7azQbHCnvhKNuN9FhkxycdHl3kdY6EcQ+rsNSsK5MS1f1mbb4leP+
iWGcyVGe1LMHMXj33LZ++EbdVSHewyHG8XnQNuSDwzhlm6gl4QjSO1ZsUEhRnmjq
uRYR9BBDxWjC88II1dWmYuD3GzjvRcTM9mit5cAf67aclwJsrLjd2QR5A1Uvkn46
+m36jDrxHk62yAaqLAfSjf8+YMysa1NgGHJrA7to3LSHjuajJXOic1Tr1Nyjbq5x
MrCHLvBd6B1lM5La4NgEjRMUmyXfxwWKnakq2guOy3ubBw/hf8+kuR7fCQeZG7X4
cBkKF3SeFqyq/V2+SvyrEhgjl6bmc3aiZYl3R7Wh0f/4CgXMum7ul+Y74TNNvOW7
H2jH09WoP7JxZwRx6VGmyCnA5t49btSziTt42JVJteOLC/fIsyVNJpxOazmfsfpD
gPZQDDgpzPTR9PAd1y2Lsg==
`protect END_PROTECTED
