`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DG9R7gH3Sea4cxzcG8+ZiPAHeDJNUhn6LNvwWNV2WU0aJwX9nJkELe4QpLbRYvM4
KZPczGDEV7IKDg9hfQ5YNF4bhJ1O+h1VQxv0JBS2ALUrw8pRREk0g98o+83LGZ63
wgp4fzcTXtzduKrnKU2PNNYk275gtbQj5lsqxVG6kdHSiiXpWhjawOK+wLRIsAGr
cdYED55pVh6vdCQ/6AVG1TRz3kJ7HaldSZftFNDpwILN6h1dm29jBMUZbmgSKM9W
UBEVT9QhvGzqQbiV9P3wjvEIi6rXAshqS63EY7b83vuM7bGLbMhGDUzcK3Y7ZnJp
vWV7YMca/qUJ9sE9zrGvANexjgQz5xKI9235Bf1z/tsPUUz2h45Sab4YHoUMOhuv
fy2OfmEndDQy8MgFy0w9ioh0YpHKR7jpePBgJAVf9qUbfoTlrdCjEuQuYxp0zaUx
rReCsfmcpXbsVgnOu18u1UINO4e9ktvy2ax3ha5ibgzNE/QGXQt3MEiZcdX+Iz/a
ojVdtiSPLu55H6WWDRIeXuIstFTmWQ9LxAguwKaKmYgFdFwGQGS8nGPgiAyinePs
LDD4ckC1kqVmTsz49KH7B1i6HYaRXXO7l/mhaokPRsYCxiRMEyxJFGASbLQMXRF/
ahdFkuAE9MTvQouSIjtBH+/ISf+4FKlrLGsUpW6KXBYD0q0vpz4bNIRtBOkiYZjM
JS7e1CQ2OyFRqT31U3q5lfJNbCcQ98kKG5ZFib//KROeVTSBOurast6Eoa/5H82k
e87TO2L0WGQRKkl27BT/8RZwnm3YeVFKUgcyTi5j7E2PKEN+hw45qK2PPHiw0QDI
KnJS7PwJv+ztbzYfYfVzF/Dml5cNb2nxPMwsxpucNjUk3vpqXClwy5ckReQVRvvI
F/WcCXApZyMKf8G0fWt+ZrS4zsbzmthoIsdzUmltqiCf9iMF8VRODyiwP1qlwpX9
+fmQ8pG7Su8bH9VRZFTN1w==
`protect END_PROTECTED
