`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YwUHwJeI2WBVHmsjCTsbcpzeAAP4PmCJUKPbboaVkmLDVDH0muzSRqWxQ8Jov30M
m6LRFvDZgm+aWshlIWaSVJL3gQGrpVQij2Znys+shBEWgG6acqZa3wb23amag5Wl
QtPvJfIYkgkLxT+ansDk/vY57EpPe9BG6d3CzNffaor87eQFtHAxTz7KSpMptLcX
RGU6I6euExHgmUPNUlEno/eAeT5KrAKCGvNO9AyJAfPsLj3lhgC5aBPZqC5tePRl
awmerPsay/tzVxSVX/UhDex02v1H4m0adPdUS+u3S1ZPCcZZMywnK4A8mpHvsosi
ew9pMRlWbmFb3VIx8ZWpKzRRzgfZWCvaTkHvUcIh4xfLKXJOb7cZXajbrP+Q1T76
+Z9NTBUh3wvoQ6Jg4iyeRjg88qct6fr+eNUwv6sMR9eGjMp38qRW7GYm3DIKp6pp
`protect END_PROTECTED
