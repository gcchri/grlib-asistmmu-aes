`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pcrJEwjWRjTWY/GOY/zyiSiL5LOYXCnoVTD83Rb+FXHUinh5gkbweIC5Eav+tfdY
K0gK7Xg4t6WWBk5xjCgvhRjK9HkBW27IJ/LPulb6uh0psT3ln+d9KTKv8eNgtjNl
BA66BUHZrp03ibfngW5eo7lFagZI1G3cSAchGdasvQ0VYu6pmmbZs4UYKk9ghIr8
5UrrUO2DwLLtdvuPgEn6a80LW9QxvOugY5/nOCN/dZann/zH2GmpbP+PJa2HImzH
zkoQsNJDuialp5zJV0l+vINQ7l7e1aogkdcsxfYWeAtOzMxpQ+koWupuau0YyMKM
2h+l7JxRsrtQNTS6J/3W6TmJ2PGFgzeIJbcanOPyIEYjq22VFQ+V+Pf8+b1U1dMJ
uct/AU/v/NcMwrXuQrwBuSLwju9j+oVks9dJqWRSVarde5O+MXZ9u0enIVNFYm3+
y7dyE9OhBf1BiaA0aOmo1J/R3ujFsXkdTWEW9KQteWpIzl+sNOXWRaG3OgoLTk/P
v0I3WonAnVmiqC3RhCvkPlf6+QplaJzE9nzv0jgJ/b5Bdq3T+i22Hf25WAlunRD1
CVfJYa7/RtRetd2RQaXdxkA8XQenfCRBO48MMPjJuNMPp7hszE7HbuPSq65mkwHM
fsjZ1oRob/5CE+EXkCPwMUSKVZnc3cEK26Zra6MDokHv7sW5UVetbt4O58ctSBTp
cISalsklrQKIJBKRjqzFWYFPOSV0kC9LKtm349DuWG3t5y/KEf8mBk89EtkzUe8v
gEcgq/XYlQfTYhOtZxR+Z3whGjrUO1LfSJ7fq9ggL0wXavAKN1tlD27Hv/U0pRkR
LG3rsWbITD5dgb4tEJYOTqdeRDJ9dvznBLYzS7OacjSOZ41gRMFz6YFI5j9sQm3B
WtXfghYX10IQsXW4mcVlLIcscV+k3+oYXlPAv76V5Lt+VovDeVgqXPjKOHhQ0nYb
b3uiNGEKT9pBH75N1uz9HVbn5LzIvoCzfwXRbILEwWViCeRI5OY9ghvuKJNsFNL3
6WtmmDrW1p/QocGxNDbNrv5hxlg0KFRGJcuxAb2lb55G1YPlhPIz51BKXSflFjiP
V+CjP3sjaztdYszTDHicbj9r4+/wsZ1leLOfEkql87Q5zYkbEUeeIA8JgEMIikSs
IktlAGEpIOVnvWLRcBnqhazsySASQb+PT38Rvgljk1FFHC0WiFeh+SHtzA7+f4CD
BXp2hJM152Krl8zfnbOtmds+pzGKbDekeQO79+ovv05eyz+RwkqFx0SX/+NlYOqf
nm3cbsDxjpu/l9Mu3vWozr4Q0CrnlypSm/27u9Ue+XryRvpTwaveON6WV8t1woUF
NY4NhsmLaQrGocjoyL5COCldL8+O5XMdrNuERVjEZlJdgIDvDhb+IPnKxYD7jxDz
iQQCZjUGHX41UJPxJwc+PhvmCdfVUcJ6N+u6myj76Kp7kk6J4WzzMODAHyJNNyPT
Hz+C8IA0by3gwDdv55oNJ02xEdXEpulixSzRN8rhsaAAA+On28vS7HxQp/fwhoud
+9qUcUU1UJlUfCmBGY+MPlnV8IhSq6G1q1b/oT2xp/tyOSOAva7TIvyp+jv6fH6z
NTaAGWlLhi+qAUMWlIuDbFFCcbobXhr87M+ydmtZLRbR+fBSFONcxu3Z41TulXcl
QeWUR7QyBJaFAKpqHFGHrowT1IXDA4ZhReLb30hgCLv5JZpW55Sz8AL15iqkvidJ
MPrOZUeFqOoJUcIoERcRSLMl+W7E2xwQo+iCGm7sDZYc1SPiX7GWlxx2l5t76s2v
pn3ZvUMV6iRfdj+tecJF/31oBEppo+je05ctVyn+9+MVoQvrbrWKcWMVbKjr7LGX
YT3ln3FqgGpykAYo/LVlGeNWBubW+3zMQPk+h3p9HhRnQAYN25L30TOWIrmr7Opv
61idSkIc5gq68mP4cV+x3R8OM7K0wfU/GwrrUyKdPpDb9rbJGniWqcp0W/78hjmx
+fk9HWr5llQ25Xh0i2pxpRnvKJk3uHe8sHcJNK4W2Nd9Ad+S8/01E6nwcg1XADSc
nsupgiUfKZHEZfcK/pTrx9wEcn3RTUWzi6KzuA/AcfHEJIfISLacGyZGgVwbbw0l
UBEFJiNpOd/hXlU9d9iwUlYyt8woQk8bJh4F9dzOLpjko7ETt20jXXEdxb2QGJIr
EpfVwsBBHwJ4euO8Uy6/4jA2/ubqgdgs6btSZHggE6wv+XhvdxuIKqA//YXQZSVG
7K9uDxNKqb7+ggxBzxK4p5KJhxOgXhBvzer4gELoKlsUcnTef34xK8uW0QzX/JSO
759c7oe/lph2xZe+sp1SNUHEIE1gPcFkU4CPUhwzOk9lKri4dOJZDqYj9nv5m1bg
NkkNQz+O4L08i4BphPU71fs/RxO4DrrvP/lS60eQxAVoDi08HysP7wQ8UUvBe/94
F3nJ7a62KPbSgWhnBJHAIp7DlpCdsnw8ulAMvCm72slJHUWyVLuGGxwWZFmNXFNR
cZqcjwJWRXOH17rqrShJJ6GigSJbSw6l9V1zbOZOW1z1YkjcXDp+I+wB3RvA5vdn
ynT+J1mi+V3GW0oQH20odo6ns7fDcKNXQolNXCUX0HPvZtfB/nX3mZG3UT/WAWMB
JkKpLoE3W2xS+m/V5sznGmRm5JDadCUAv7/zpYjQ5JfVF1Ne3ebzg2nZI++RGTJa
mVDfPxBJtPslFmmsmcXyEhyHFIYZXFsHKTPAy8cOYatbzSOfOk7hfjfMYgNqHoLh
JGpI2PLAJx2Cv1nREXCHJOaogx+6TJGS48RnjHtnEvN0oIpaLDaEqJfh1q8/WmxL
lJO+vLnQ3g+4qsXln1XzPlh/P5+BH+A61MZ4/13yPXRyi5hHhigs6J6U4D1USDnf
xc2QMggKP8UH3lY/UFglaYaCmeoPHGvPfzpymHxUh/pyWACp9YOtSG+zwXGSWtm3
sXMLq+E5Qje0pS2w91GGz4sQ3/YJPQQF0kCU5sXv/r3EoCD+YywixW3T2/zS4F9c
l6YCpdVzm7Bx+8j4XXOSrIyWdpwc8EBHtKp80vcBVIYhI2xYbvEAy31of8NIYC4v
RxUiKJ54s237YXHjk6rxW94M6ErSK4QI9pbKLU/dvLAhSQnv4adS1VvIgdzw6wP6
a3zIM7sj/prJr1AZBLJ6y8DWk9+p09KWd/ATmHP+FCwG/73KpnNYaV+6ypQqIkTA
hFNoVNkAq8dRL01Ejgai9drlFY9lq4KXnJQBRlUohcbLiBvirdJj9wTRUixezFfG
ss/KG3+SEDCJTE/QvHa3VoNnMqygEsuMd3My1S0aoIUU5z9Y2eegUY9pHJArYVkG
1BYRfrQmAcVCxsXBREEePZ0SWfriQRgSxiOdLJ2++oOtU4iaYc9v0SQHbW8/E5H+
eCoan1d8jqL+/c1lpo0/VwGvbkvV3pc2x8jMIqVst6JWaI/MyjTAVxFu01IfV1Fs
gmz0x4t6MZPHTWxEVf3nQnl/pGMbzKr5D+V/+SsU7LfX8IZOqDkIk96WbJAlLA7K
ER2YoRcECUTALaPGms+g+ItD6myvbAWYfs2LJiv0ftaIkOEGRVWR5H6ncqMkjtqf
+PC8FoDzX2a/N7GojUko7WDoJiywQFxilOljqflpsyumlXCrXr4saVkd50+CRgDC
9HuYCbQjNYFKudQ82lTd7/bqkDDYPEztGVx7STZswU9PnW6wGWxCEOvd3kFb3vx/
G0p542vBhz/ODYdzPW2Jdr3npgeAN7Nc//I4X9TmFv5acvGwDUur5DnfbC4rZPHj
VTN7Z/t1X83I+SPkAVYQ9pVheOvD51BW4yeFbEqJTn10zxAZbLYQcoQ8kSvLrAzw
N3VWmnPWrDm/bB4dNwcxIQWinfe0H3eDEXeBYi2SzDSBmnHFCykx4y9QyNnSYXrq
ZFWoHbFnmuhroknxGYRU/9pRSZEZWbUM02BfV3Ui7/MUicVzr6bQgXrginWymFFa
n0eIMuBy6mwNBV/xknG12opiD60c7Xn12gJ+laIATTOK98iXEp6vBj9icVrdA8/g
KqmmDcaMC7WzIKj1fsfdUBjJQ9yyq/mMJa3GFS+AaGiRVGyXmGqo1m9emoUulD3J
wfIz25dGaOE5dl9mE7xQcAU1cHMCRTFoJhGP87IFgrbziYeEj9exlhJVEK4439Xr
fAhvokTLMX+iuyQRpFzdAMfYmYY9lRWMq8Mf/7UuQgNNod9aHJd4zFSssGklxV0a
QkR2f01iC5o223ggU3EN7rMepOMekrAUJx1CVJhoV7syfAedrecGwyUsyhu4Alzg
Ri7Ib4TgkUouBu25rbhLN0IAplUOOctTbSKt8bXXXQI82KWAQQfpfO5wU2DeNybc
FI2rgyrCjkjdKCJG+iOL4+jYxuJbMvpjSVOepoJvqlJ4Cf6AiRnmr/zwJd4Z4HJ1
0USKM3ddRMIWyyAk4X2lrHuKU+gEXoMMJ1t0MhAOQDwksp4mPag6bx8j09L3Z6Wt
PWSTG4GJNaxbj6x7Qk9SCVgbDv28Qfjt3MNTNX5riXDCES6hKeWaHaNlR4t4nVfn
Am53yJU8FqS1bp3H4Fl7eV+Rjq5LHYPugiDe/IramX+/DnjJ08zzByZlzXd0fD8K
CQdIOXoHHEJqVsKz2OSozlat1VXi8v3Wm5sc4cVJZf7n5Wq0xOxsMUyva8tgBVeg
AEs5NveE0VLtyJGdST9hUcPmt8tX5AM4n0CjwbRmHQnkzsOO0UHUrdug5GNrWJGK
oT/h81bEXyJ+8WP8dswB3i7eXNnL2tIRMvv8hMZAXbkx0vhhRA2wzyRILMxk83z4
gXJ7pYk92GJ/qWItTtcMmLC7AGMAjVNdqJYRbh/LYSVSJb8b3Iylrr+xa0CK6T5u
hVXMYdPnOhvrJdv/lbhAz/YjqzDXSIoWozhOmVOoWoZBy2n78KVcMpllphAb2iEi
2tBq3ahrYUlQWyHKFx3hOCK4we1rGBw2xmB6B8G2Fjyq5nOqewV3XkvR08sMCTEE
y31TE1/85Q41tuNjXk0R5SKvjyB5c70zjq9pwe5zC1UoNMWwhQSPmP5fENHCiO8B
BJNv3kYaM1ZlT9VDgsS5/CFuZFuE1VHP2iScsL4SJPO+siIATYXvcXJsPMB7vISl
uf77Fm7B8TRIi90VUzG/OPNF4QRQoypKo9ToBC5OjntS5XrY6VH/XJDvfKsfCRi2
+HCyCFoiLZOvAh5++SVdpbeag64cyxI4o/dC6DgB3vTxClXjiY7LNtRJ2uqPyRrE
W3AYOpPbGJFAGnh+H3MFSA4vgKli1f/n6du8l+vGK845h11FDHxgO7h0Hc58QWdM
KSnWZrQZ2aliVPrWP2ivSGPYHwZtL0Ox5GWb6lbGoFYkQXtvYmTqNO1shp+jZxqr
W9SZyQD/BFf1qdIuL7+QZQISRnfXLBO1oGnk29D8sW46SHsV+10+WpKnuGdm7cK5
cUMSxjNtFvMqiVxqAS/QpPwptfojSSnhi2NRr4J3XnRF5s5/HF/v6Y7PbZeA22ej
LU9BsCfDvPu6O8YutPzYd6IwQMGco6GUMYrmut+pLIeq8rD7Jmk/+/TK9o93pS5I
wBFa0jmPtNZj1hDE5MN2K219XY6k9GiFSGvEvhP7l2FiZEaujAYbVxCIJOo8ira3
ZFtPDBdifa0OnKLsxwPEVIUZ3IVvZuM2hyV02Uy7JiZKU7qa/57mDWlLV0rNeGIw
bmdq+N69Ewh4W/yYBUTq1cJOwL5T3vor9P2LZYgnVaPnzIqz0WjTMRwhj+juTWHX
wgkpw/z9a3Qq0D/kkAQ3zeijpJ8lZjiCLpEHfzTtkqWf41dJUJ9CGBLNlrTv4TUZ
DEUEnbgccwE/0z7T1ESi6DR3Gz+txYKR4HFgrh7nqCldjww3w2NUweKbU4yMV9Jd
cVjeWw7qVie9D4NsiKuyWIgX/sLTOmZoN/FxJXik1DNKZ4ZpxAqdSHQK05IqqFv1
VVoaBOs60sjFlyfEP88RZzzKL8sSaIbZTuzyjHykgCo0vLf7WVpsc86SVxcS6rX1
AuWVZaB2COqMoJpzdUDs53soMqYBwiSNqcP2xZy4ko32bDP0IHPhYkaNKx0sveQX
gbN86U3UqCTM8IyYRFoaHgvhmcSk2a5NLn03hFfj477R6fkD0/DvLc0KVcMUshV8
j8CxmO/2kuutiD/A2LHnU1F+nTZelGclHSMgByTlOlPXLfOtUoQPN0GnI1e9nn3q
jYUl9HRxlMsLj1lXdG8aQ7xwP1rGdfkvR30oe0tw+P72m4s0LwHlbhKb0tdYcHKx
2Xh4pp555+V+C5yAixBGsgNy6QFitr0/YnZpY76JeYkQZbX501hBagUNiQ2E91FX
pzQr82didUlP8NaYMPzJV+9gI7ItX5y99NQ+XzBYfpSyiQtcAfMfTSa6QBy2S+5l
XxUtaBYvklpI8zZET/aEkI3n1UZmH12Pa/lY4Vqkbxcx6z0XQ/blayOCggirN4ZR
cWDc6SeHhvCUFU8LBGIHxWdPU2B7aVk+ZhtBtUzA8A5rwa2/OaeFXLlg2eX0k34D
TsndvuZKYvf6bNJFU/Om37GASE5oAoM/0Dx8L0LutloJIRZ0FHePydXS2zxifJgU
+AKWl9S3qqtH8x/wL1jgBpU3ZIw/EEH3bzygVi/FM9NlHw2cT4ZdwCqdOM1nb4cz
Pk8onK6BMG0PhTpIh5FFVrkQtxaBu4TCroMno7Zd0NOhu2qIWVjnHY0oxi3g4Bar
NTq0Xfz7Ii3TR5vCtOXXCl7y0gz8TpdQXuJcj1iSGxAfR0SrGx3rszhHOFGZQfYq
1qGAuulq2sdtnbEjd7VIEaOuDPwVqx6G8JOlPCRLNhyD46WQ9wHLZ4RF4Y1ZdrXg
oVaDbotMp2u0ME2pgghq9k9nFWtGffk9g526N82JP5gquEM1VDKV33RNscvHmxCv
CG9kUfRgTmBCggTQ3lgH2WUYNxAtmmLW0clD2FhgmnhI8Sx3sT8NQWI6D7AjtDW4
QC6i9HwlbExhfaZL+6C5uZuenlsmklEQ+u0NX8JvsNK49qvATf00yidBRME0QzKg
J3id9/DuBrRfslrTvQeVDJckA241XdLQ/6e8li222CFslEWaOM1vnrv1K/2Ofbcj
PA4aAq1Urz5ndUnMj2Tk6ZcMq+QxnbBrGYMyEjbvB9NzSrC3duDpuHpNBnFzeacd
KS1xQzGiH3eakswxKhymDPDhW0KZMtjYGa2yClZX0C8HuVHCnFrJljzr9ZFDo9Ap
dXIERjEkajGIABzY/L4a5ayG34zxQdBP2BFTuxvfAdXqjmdHIKCh+ua/cxZBb78X
iDFWkrD5HGfOTaKoP1mL8AQEAQILk7qr0xHSVZiZ5rnOVztHf2KMkbiBj0Y/eLnO
BLYKL6h7p6ZlKX3rbQmjQiavYhNHbDPFnn8rdzWQ3RrEl1qeQvigvbMSwTEXiNRK
hNMez6nZEfwD8hMbxYwO+s4wotDHLvgNjEb77BG2PZZzdAark1vPbSaWWel3eJw7
9BAvvjxMM1nfffaZFcXkTWam8XhpA1ceB8LqwIjSixitCZ9wMcS/+ujIRCf14QiC
texSJMXUQzjSubZ+G45HPLuWhey94S+Njkgowh93MDVBLhgbjpshG/Ae00zuy2PH
XCYItCAM+4qJgqVnjpLdVGGT92JFpmDxdSnRuYA1uMNfBW4dhpnl437QhSfQVsgQ
y73ysxa1O9tP6OGzyylQbP4ncgKV5m7B1r0B0CXcZGFwgmb4gv92TQvgB7j2dmrP
LsxY47a7reeCmdor15DPGB4ZNfFAm4WbcAcNiphte2HJEWVTSzZGXHQhqQgJKhdi
ik4Ayu+f8GuD5RKJT3hxZNF5W765CLxYzavAF5skwxzpCdcBG5MWUcYLSZczd9Wh
Nw9GIvMFjzBriAmy8vcl5ByYR3Q/HCrKO3L24iFch9WovSfjVelnwaiDICVRKdHI
ecvsoEt3ysa9VMHTtLsjFb0UxDOSjhqT7pj9eMnbFP7rhQ7eGBp0H6fPCNpp1blg
zB3+d13md4bszo3d7ulgsT605TK5cd7p67JgECU9ilwkoGPc8dUO4h+xWbn6BwjZ
52g7tFWxCVlAgLGNt16tKxLQ7eDLf+2Y5sVipqevBVHJwLC/cTeov2hD8EscAGt9
qlFqxRgi/wPuMxsl9+WhZOVE7MbI4ix6ouMG6XvnAmMQDVNs4vMvZw12HUqT4s2D
HMBZr8QmBhUWOL96rapHHYNOFx50pIgqZ5ejuJL06Lft5DVfZ1ZAnh0aVIWEBntv
X5XkEO8wlAOo32T5M9BcsOZ+VouEAMbegCZk1zAHaLeobasuRGJWIwl6Gp8q4G3B
tDRHzcL4AA5ygr113E0QgqvKxiTuM35Br+2lMYC33iuf0j8e/kOWaLUTdylPbpQw
IDoqxsJ0iSf5M/pETQReBKjFN7TTfCErXkKfdxlHnLVJ2MhHYMf5t3ZyRFn1dzqW
vPYAaQ1B6RLdA9oYtJsU22xPEtIsWnQR27cnCzh38yajPlO9M/I6YCJViHXQIJjv
Q1fMUIS1DHDhHH9m9MnEJgRQAzPGMxXW95V1pb6546PegRqRWDaC9cl9TQjGgihW
LjDxBXxMjl6hiYHV1ukMr2knPyk7PB/Zlw9M60boTr5qzQPxVwslPwWf/F99ZZDh
Xk2XVhcDZXLacniQBXgNOpb2RN5LZUZnk47puRVPrbIiadnU/4TAsS6bbJAN1vbp
xnlvJ4lvf4oecRUtpx2vNxb1TMi2QUJiUhMPKBmxO5sE5MkuU1/U4isHH6KOxFcZ
tg/FQ4xVo/S4TadpFB/HGKwlKmYerAvYN5hAcluhY9z82G+/PbcCOb3IKHei/LTO
nf3/CTm4G8+64UyusKkeSZbJjuN6ByjdrLKXMkpROfyewqQ0AvbU6piqGOaM4KfP
RqLidJuDRe8elIvOJcYd2T/jf5GXYrjg+8PIW1mLkaHPty3g5HmjEteQI9wWrESG
R5HCcFkyypHOnIwHH8V3yiSsdAJoMVJTNXrH2ihB9Vo7M1c1BshkqVbcpFes3Hkb
t28Y7HWmr0TsEtYfxNGflbv40GK+pdqSQ8awYLKWzqEXN/R3XfplSnRbGcu9jyLX
wGpWX29QT8CLDSL8QiywdwhCX5nSG+0o1pTHkKHFmqvWwn/1nCPKY3mYuJi/A84H
qTTezU+qwIxDslHedYyae5FkpN/Xuh3Km6oZJVgvBaXRDXGSkKjAqp04l/mydtpA
Z/ULrgGhmpJ2pcmx5N0ZeXVRluCRhElYk7pw06do0ToUlrsW4B4QinqlT0YuYyCb
34iLkNUY24r7eF+52yC59d+XO1aPa+p/oGTVGJ7b/Iot2dFai4Rn8iVulrxsepne
uW595huo0ax8kF3/gcjs+a2Ez2zHfh2OlQ9pzFRyLbBp6ighe6MKwCFL/H9ksQdK
+ZSnKnAhABW0OiFStj0il3XMay1pofuyjRjIrz0xFYMfxK+gFlFYJ5DHhPPXtBIT
YUqkLti9K+kTZEy/uus9U9O+64IxSav4J8NGz0zHZT70icthKZVNlyRvc4JE+AJ4
IlzlaOUv2SFdnx9gNv7puscUGOX2PvlyY5/K9BuWZSk=
`protect END_PROTECTED
