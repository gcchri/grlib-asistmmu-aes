`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DINyIFHc/Vf4HkPZJlyg3kgIXho1oshPle2IU1cHBuMmGFQ8N0KMpjQHXZb44tTG
HjEPwiFzge5C27+I9iZ3Awq+piH1co9+0LYYoSai3aqiEtYAbrwATxrzFip71Io6
+aQWdh2PHr7bfWaBI7DyUsGsf1T/B6tUKJJ4X/srvGAyGomMB7W9vp2CJKQvWxlM
nSPAbfJaHTpu52R7nlV+d740Aa5AQiFOm7a5fbDaKu6v4R+ItB8ivuVgzlAvSoWn
oCwCgcF2g+Kdr5AMPjwqXOOg3T82Y6O4dvjex0gpU41bTEPPtBMOJx7rE9t4Qbmd
XGuJ+bR5zdisul7PcdYkx3P/kIoVS3mPETWt0jZymx1TpdGXvf/m6bGyHgxtxXS9
mulE8pzljan4EFwbQO8Ym4V1txrJ1cMa0mR+BmjfHzq5Awy3+1DSPmD9eBhwb+pz
zZgBSIH529eb2c8Fl40+qHjKUmPVobzw0sJOvHVnlM6Bl0sZ4M9X0K5CRuBuEvpq
`protect END_PROTECTED
