`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DfPzsbycJjTVpkIW9F5D3pqdkx07ybEZTk6M3HkJPaNp/dkLP1BuDYvd38iBFYUi
K8KV+bEyQTqgcazo4BxCGxdhVQS2si7Ze8BUcGZ14BMxFiDIuzFZ2YG9VnUGmIgw
Ec13nTO540izhVGUcVj6azXT4dJHP3azjgyk/g0XqX8ruWYiTu/y6QPL7Bi/LFsX
yrnSbtwFCEImTHvbOUOxGQovOOE2FUDHa6ZgyIRpF++P+UY4ulLjMtxEXrKilLg8
LCWs6rF5Kqr7JrO7byPkzEE5ES4xzozXaawD1TkRtB0lV0HcrjLd8HQ1HQ6yqel/
dsODUXYC8Vo7CBE2+22bIncvQSO9APS7yW8svGFo2oa/yAq2Ov2SDVhVgTbeRYiS
sk1S4Up6W5zsCFnCyTWYQQ==
`protect END_PROTECTED
