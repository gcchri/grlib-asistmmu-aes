`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WqKjLYpxKC72YLyr0xJn++Gh2xWjZYEp422seOI+fOgA9X6g/b2zP00QW6V2ADAM
76Y3vjOaz2n3zfNLHgkxXmbcLrYpAeb0Ukfi/xtxjo66PH5yr/DUdSVrelKrkZtQ
RX8SQMIjTCrYlyDQEi89GsrmCVTv1TJJr9la2nd8F5zoGeuHqSAFjtqq5uj1ZKtR
Cp7H2sl8f6nmMjQL/of+5WFaLpkm0YbCY9JWymEdBc50dfh1NA6n1K4qSs6Yr//4
mjtkQsmvWo6VuXkhdkO8lW9JsT6Gwyhkbcrkhf62WXZHj7cq6cFgw1wHKQ/0tC3w
iXoOKaHPbKd7+AgqFUNvY0Wlx3d0UGTLgsD8Onx/YFwZTainIgsrhm0tS/RybS59
FUoL/n2PpSExPF6n5KBPOOG+imNh/Sep6gqAj2/P31bGRAAxAwlwNUH68TxGHs0d
k6VqYJHWe80OoQeGBMs/0JRN2phiOOq+DKjpJCXclm0M2JoaEl0OjrHkqefqJW8+
6G/ROsndHwl9lmFFc9T3Rre4Nn1Tz+4hoZpms6+UwXxZCkKk3YI8uzLXUTsdhIqz
O4KiOojyAfYS1a5lEEVIkbdqtDDZVVDMFNV9r02SwLShvezDbYUb0+hqX3/2ZZYR
Mc3bPM9U8juiAmCAgjhGsrLulN6sjrxHGV1+/a4CcXUutrxslgM8i+8dtTOYYeAG
WVpfahkValErus8upcLMCftw9YwpE9o64tBKBKOSBFM96nAoU/GT9D1MSwmjyd0G
MgWWu1otaKktL8pUhALolVHdJ4sjgmzWMNO2ZmvZuwnSzwjLeh7b/w5vm0xx3Pu9
YM+sPNT78FhuLmzb8JGr1jqAhd/0anHDNVrbVjqAEHt3A1V0NlsdBsGloY7ZhNik
RT8TgCzsExn5PLamQ3EyRlweqbPyPv/xNvoF3y5kGE3RYs2ggiWxPv7Z8gRk6CNd
6trXECZEsmprwZRSs2qMZWEjlIUUFBkZMG6KHgGJU51jhTfdAtsFyFFgBGMM1Uat
yGK7dKW+LPDr4/+UGJ94R/10wFU7w7znh96ryNyi5gETAtY2i4Ye2IZhY3E5pwcN
qG6XUSiHIrh46ztKY+pFuAnYcrzNmGJLVd+UdneIkQ/F21B/Mt2w6zxSxqHJMGFl
`protect END_PROTECTED
