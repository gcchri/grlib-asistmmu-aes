`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o1WRQ9ORuJe3XBYsHTKwflkEVD8LGlQlh3Dv8eGY3MTkdH06SYVTAj5UCeXo3d6/
c2KwZONFOrOAs9EFgcloA3fmlfQ9WYQOJNsRBzQyyMMYf1SXa5RzlDxklRzH5Tci
W0/uaZr8q2Fo5lFDcX5WSlrerQkui1/UadirHrAxmzKHQRiOuJKPFIfrFdmQR+MY
DZvVJ+DhOW/5KpIdxrw+KWjq+b2z0dLTvK2dxWHNZV7EI26JDR/lHr/3xFJrmVuX
ltmq6yVgJCMTtXpozg7Hx7xwPJ/7L6RTDiM1bTXlI+VIyFPIk0+Rx7JDDzIIvSr9
bvR3TDVAec9TT6HR7zfKDCNra+IBM3nLOA6vqQaqTapdL/zl7z7w7W8OcNIkrLsN
zu8UEp+6Ric7FX5DdexjcVGh8pZmBGeI9gvhGauRBShYEq6HpM8f7RzBCpFHSE4P
DiocVufm0hrwc71OlcVi8iJQrANh9aQPiCoExVtJrNAekzeqfPWqdF/XIZruoiz5
8bx7ENJf7K04n+FvfNoWeNNbwB+giRJ/TFp+96wBTJcBYAiU2mlQBLQzOkpn+j1w
U7JFtR6VDDbOUU7u5bR/KixwPOXAqsKXm/WRm4G3Ig/iXsTbyTz0fwEc6U2J0z93
LUoBuLDRuwo69GNwfkin0Z14DVAnhEK4J5bLwBvdH5xnnmGp6dBCxOMbUahcIP4x
+/EOmVyZ4sp/HzEz4Dm6lMD0mabIsb7soCsKuUuWXRzUPZBBRE71K0mO4mO6sGBJ
/EdxhmSfGWakPJKpxonLDCg9KzjV5LSjzo7cVbEhesN+wkVFgIxHG4z5tm7xbO95
H7C/QGqDxf+kiiU4qC/FDi8Xjq9f9GNkjlyf/g04hmnsBqsThXrVxxE5jcl1ui4n
BE8bFoHd2jbTej8MuB88JevbzWvWSsNFn6ddyjsoTC387lqEMFLF3M1aVmQ6OX3e
x+vqfXXil4j0NeH9xx+ZH0pTpomEPtZwCi0kSRZnscc7gw7yB82Wmc9IZ/jqHrWW
7pSF72zAq+1YMGLAWedSlIf2OzH8tGljzF/pB/1XWkWyvISfeyz+O9MO3asSnzGr
+36elarPkktWatHk5aQiCOBNPvxyp22w+0QkhSHKdPCHZWuqaeM29dpfcVFJ6IY6
n26fYZGii/RJoQ/TQj6T6hXT4A9MxF+WPGaWpkfACl8/JEQDUltSwmpPOeY8dBqT
QLg6IOWuQWiJQU1uF8INqdufijTxtpA32IrkOzj1jn1Xsc96krKSRXckQHG6fE1I
XmyUgepk7gOWwaQtzjgVgaWu9A4+oRQApDkm4W4OHCRv4H5i9l7Vqasmk7glxfa7
kheTr9qpJMq/mNgHEhj58b1S9OBlDiKqYDK1QEtVXpKdam2wUUNxbmfyslx5JvXU
NPtHYfW6jc2mO+5jdBKoumZY1CFKVRIX1hoQd8qPTvxwpcOd2BoPbNebjS8o4xpM
BRLTr2y97ZAKpnND+WqPgC3AzC8gd1PN07tJeNLkznCZaXmtGdJnHdzH4wF6qPyZ
HOWwxpgGUUOIZDVyWSOMxmJ28GwxVdQCYptT6qfW0yomObG412j2c56JAd5jeTO/
wvEN/OprNt3xX2Ny9nD2LfnLBQVT2TKhhY9v+4ckCmrpe7A5wEgXBPkcKtTGUgsd
DeW4zbgbOOLjp0rZIMx9PYKB7LkizC7FIzkYCB5sZYHM78K3NkxDVNxR1U5jG1Pn
JrY9VmIA2qJ1KpXgC+6KmunNthrr0pxiPkIrRnvz3T6ZcOeLLAnVaCekOODfYUkE
xrTMMDbpcU4AAlwKP98Cq1/89joZE6m9CNPXRyKi+oWhDVXxmxojP8n7uo2plPDM
kLKuY0frVo3zeWxt6qOJmKvEokizluwFILw7XyHSni9P+Or8ZSqjfdyr2+uL7NgI
2AyM+318tdMN6BxMXwReBQ/jb1Z37sKpi77parXwY9yINqyixeyI+/LGkXG/2IlX
fqU7ULJUuLL15l7bCUo6pLaKWRQp5GcWz73eA+SWAVBqvy04bCKD+E5GFFu/sAbx
8ZgGfj/EBrdOHH3RScn7cN4VIfVi+zf0kQj7ieaj0/+LqLjP410Gxez3GtvgzoTN
fjB60uUXdU3riWvUr3X2WET/dDlssscPbw68B/pq8iueiZ2R3tRFQIbH7HE2Mmpl
wFE7ToHll8EYqDeyQNkA/pFZsJ+XGak3DnG1a7oCnZqOQwPX5qc+YzB6SY6kQRXe
DmYAUDjEptVCdP9/eHnWjLlzUXExNLKRXRTP2XknEz0PJ9SmZPv7DtzTH1zrk5nS
BGoUNnm8No/2by5i+81VR4JmBv6NlRvlm6b8BzVpSNWRCpoaO9uiT4bqUXpvOVfs
nMNMt0v9HGEDvAAfy6PYR3Q7QzPz3yBX55nmSbzgZ0Qcrb2BFGdJBqK5tw+3F863
mtADe+AQUYdzfmP3WmbXtGkUhaPxZtFQh8SOnKgbHfI1u6xpVVCCk8PpN9TnMs84
fgvQrMaYzs3Awi/cTqaAGyeWgtaHZAkY4V3S4KOcYSORaJ4gtwXN5nMNIz/RD1bv
3zl8fPjCIK0c1OnOul9iaoombZunskGynfmdAFW64wMSzuEBph2/hHPH+lA7g29G
KwUG1qfenYWTwgm6ST50BXR5thB1soXOZcCTFxC9ZGnalk38AE5QqhoeKMRoAfvO
YvwnIpKrOsHR3PmSCWlpvUXtrRWyhZhBEr4vqiGlr+X9/T7+pOOcrk4mvpVFTAxE
+H+ZOGhQxwT59vfOnuZfUYSdWjfSeiBgy8VdjfH8VXGBCQDTk19O6AwKVB4OjdE5
yomDxrBcxwIP8oPvyuorjf5hmByWI6vbLsqch7ewUQ8daQ075RROc9q2kHCUv+bO
A0NoeePMm4Xs0VCZsGIDDZPQ4dtTh+xuoDhBGc40y30yViFaKvfm6FiVp5MDlXzC
4sWL/FInCIKQ2OQjrFw8g2+YsdcnSIiCNI3QlUe6ah5kJLbu/4f1sfwGXA9L0Cxj
mX9p1EwQ8Bxp8XbShSyOKCjomhpmrtj3XlQofdyZR9T9N3QD2VpttjC1v7u1Ff+P
AkXrSPwqXzAMNbhXzMFduUCZzLliJY4xlrzymlKYFWUhlQRlurhEx+qkY6uNjhGh
An+saduerqMoiLUJcwhpYhuOD5mJnPVY+f14fM6nca14f+wbIbHiRSVqfQFi4NxF
tsvVQb5t0fFM8BoAtkR6TeM+4ibh0Cff+7NWndgsqo/VrZ+b7Fbb9gWudbOiMbQX
Qp/kzDZ4eoflU1LRfXhKjCzstfM1zBbOTD8i5e72dyugJem3GSLsT28KgCoMtijC
MQZfPJZsak1FfFg1ngcTDCnPE1bd+CKi1yihX+IXwi1msmrEXQAvJ7ybDKe9uLRO
uJ2p2DDTggXH/L/ytblVRw==
`protect END_PROTECTED
