`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9veJGUY0yRlbvJSM5kc4qu8Sbt2vftZvnrdG8ORj/yQ2zwrRDXPIDymuf1AixSp8
om9/vq3HXKmI2tIb4afq89U3Exili8pqebcpz90UloN7/+83XNEN4jKcNiDVBvq5
KExRMJbp3mkY9DFsT9HmfiH1HzUWo6IwDPPepv/lEXPB328tRdUIqpbM8pxDdNyb
9dxpQ6ELh6nUivXT7tFJJgYLd0TkGnVL6a+FSMbGiXCpOSS2jJV65UaT0iBDrUeR
PISHAZm8q4lz88zBTC6xTc0UJdfeinuGSr/JJUaMKopEJXrFpf6W0Ptw8AeHQpMQ
9A2lCa9EBaC/Mco6uLXxVPveUQiYXIO3ivVrVaNoFkFUsLBd/i1WuXDEZevQIF4l
TrJ03Oqwd8louz6U0JA7p9988DVSYozH0xCGhAlyHML7QrqQy9/HWYQmSilC6KfR
791YNRsTrYYhNWt5IcgOBW3D5T5pNTMQOMSeRyYlJCE=
`protect END_PROTECTED
