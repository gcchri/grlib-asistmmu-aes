`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3PaoMjyY8AasrDbBB9enk6iEKEN87h/r8TV7xCu6Yb7+r4WnvKGeVv36qwlZoGMC
UT2cQsVIPfGzUPj8CXDZv/dMp4LtQBLh0SyU+zO83pmCjFlGoOxdID8lm1lNjpUu
yJIMkXcn6sdYQcYV3bEhHUMQQkpMRKeK9pLRImsq5QmL1xMhw7dPrT7qkHSt/5U3
RpP7CMFLaQesopjns94+FWF1/RVt0P5ay+2zzw7sUosloDBNojXvSudxAJBEZsTD
IMmSi7u0kAFUkoUEz15hNtqZHw9bC9gmQfrttGPgDLMhdAnjj1HSRlmb8LF0Ah+g
uES1gHhxrKdd4Blw41KM5GouzxxXB9SVijZ9duM1/7c=
`protect END_PROTECTED
