`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WTGJ7940AjChwZCvp7F5GjMykuzlWgHMk5gMEOvMh44gC7JAcpxZyCWfheZ4IP8Y
smuUejhKXbzTm+uqh0a0xsPtZdWs5IQf/Ll1PCcPu7PRASE3NCOINQpTS87OsHv+
gbhuDU1xHDEZ7tvP736G7VhPw2SYk9z9OE6goPZN03tD+VtzpZw4X0akbpDxy1xg
oCuG4cslhSHa91DjPKeurgZL8nrhHwvLX4rZX7kOtRjpXr9DlyRSxrIYlFDJOOjZ
cP1Bq0THZePVpaSSt98VjDvNJuQDGrjgfzaT4G7fxgezzQakx1Wxb6zghuE1WeaE
tXrPAg6SiH2HpbP4SLfnU69C74Tnmh7CJ/tKuBQ7VVlgpjAgm7+K99OZw1fNz7Lf
ovUJhUsJkYhp9D0pm+nCJXav9V1bOrq+/kREMN4Un4p/I+IEkKftiU1nCWdJ+3BD
zdQI0+ie3nrHcCFgugcrqJCI0LTWzocK3flKgpwggDlOLRmCU7TKjKlKgELhbJ1Y
A1V2l4XQ1SyVMkyPYwaEIBh8hVD6D0mbV5Am1YDR40qKJf/Srth5/u6SgzlZ1fxb
4j8aeM92La1us2oAa0cNAQWhaRHOjdz5Nr5hmYsF6M5iR934K//x2tGpw/u2j2J+
jaJf8ANfKWdv4sY2hJMNL1axzAkvvewqjfYKa29FfkFt4AOHrau0hPzMn90S1Xy0
a0x0cYsoNXpGiYboM5DfyVnFiu+WDJxTzuGKHwy//RT1V+JWpACKAV2VNdVafpMs
O0C/eB4ZzpSf8+6AmiiWsg==
`protect END_PROTECTED
