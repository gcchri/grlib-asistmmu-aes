`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K/l210gGQhp7nKCt7Bt/iEUUYHbcEF4XkEoEaxGVjmm+L2oYcYwbWRRKi7coeTmr
99NGodqm+vn8E+852L9GwdAXR5esDOLAfBeNXyxkV/dQM+kY9x7SvkHyprJFbv24
6egb42jPA9ePeiNl26LMXvYdo4u1tY96Fo/xjTY8NgZd5x0djG5shqqBeDRN0Oip
Iwy2v36uHTeqhhJ7OKC2FqaOXO+IQ0BBZe7APUUwdF+fgjFnzV5UnCi7Pi+sLJ1r
spwUbrS/0z2pdcNQWPuk2lmfZfpDFR79ExxjBWH1hMWNGm+KHtOWhj7jj0l2G+A+
EEyCWzs2XSl/y55GADhY/HlqK1NA5SOgT6drFUDxIlpHhNZ0ZkzhAC4GvFGX0MZv
cHroqdg02CIDJcxBQ+1h4OW3TmRGbi3Ep3k9wfh7DogKgGZa9d64HMVQnWRmDDOr
xIMsxpILmKeRC2C+4pyznXGBV1GcGw2oiz/ippsUaYv1iJDEkWRR6T34FM16GsBt
yfkT5M4FljmGxG6zD4lKB6uq6ooekwZ5NZdQe/z4hKLYXd5CQtt1wbpl9d7UiMp6
RgYZIeW6R9W9Vam00inWV9njw6cVqvWR9LwMhxvw2sp1F80bU+j9R1jIlBGBnTcO
Qj4OuUa0J7Jh4Jo0t+D3gWmb4cR3h8BM1VFpzGR2I5DpyduI99Usp6heoWqKVpPM
8aacgpFqzL2DFxtT1wnha98yCQo5kcg3s0ArzFinHhrfNGn75yecgD+zhnz9Otrh
RtTsin84f+eMfTaC9wQ31raTL7LKnF+u96x5LQxuPv0q/e/wrt3EwK6tuBf8fXIA
TBRdF/AZ5Dcpjlpdf2oEsegJrkqSxtl+gNw6PBn7WXlAIJ3hJjm/QSG1V0BU/uNy
+sHbF7waPHTlUTj8vxKVHqCQa3lppBXZ9WH2xR5/63dNvVg3MoyA5OLbJzMBtMn5
DPJis1pBboG77F2cxQm/T6dInlfPp8O9w9vzTAkKG0CRULVoIXMXybpPtlM0zFjP
7YdlMMwY88+EyRHZlU7R1usjvmD3gLqOCwXtybrqWOcot2URwT0rN15MrGZKbM63
Cn4BY4P5PBVeG67d5V6eyL6Z2txUXD0zdmtgOBXPnSkZtvCoeStvAO87F8chyN/t
`protect END_PROTECTED
