`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DfcUwt16wl1AlLY8USOD9x7PJ/3TvzjYrnqzJZJr+6fBiQd/wY5q5PepstyPVLKR
arOAn/r0Gq5seP/WP60qK00TB5xeE1B+1xklmVHXyh+R4ndiuynXyNMOoCC057JB
IvCO7omQe3wJM8cxHlNap6tsEAHXbt4FDpwCaISRl2gPe9BjKLy13gKXVuNjmppB
NDjyB2lEMwCEk4iTw5j+O9yTLYFzMoP0zGlWqjWtKYj1QSlFXjneiPDJgLH+xv7R
IzkCy9ZUyd0zGE4kASVVj4hAt9rPI7eVeJzVTvFRLYce1QQ/ccn8CXz14nsgK3Vu
JJjmDyxGES558Xk/oQ4mUA==
`protect END_PROTECTED
