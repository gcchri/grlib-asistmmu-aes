`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cVGmM+FWPWwCpJD0lKrrGcPOTid0AWCIozD1nwhCb/MZxDMht3aXw+CHXYUGIUbl
wAU0nYH8ntZlDAQ+4VQ9bWa9gTfpRj/sVhR5V6j9DQWmn06nrN8q8R7lVRxwjscU
hXlZLjAFq3mTvv8jmzwqAcdesUdpKSpabn/i9qO31+l+DaPUI/NXtUwpl1EYo4x4
rUOWIDZDRV+IukQRIrKY95q3qDg8/GtgJMA2NhKlWfkuml1UMFBg1FyCulN7HQOV
jIkS2P0brM7Tw5gSfzdpz9zdmAEWesxtESiAxBCd1tWZDCfokUJKV4jMGqyaGkqO
wknJcP1VlkyaifXqN9ijHel6QW0+c/gqd/4lT6LRL9B//r0TG7R1VDbblSMt+xf8
/zLWbRN45M7M3B9XsqFUgKYI0d+iX7M8biFyDEW9SElTUCvYarscRf5gYDWPBCdE
48cdGiIozh4IEIxeO6te1UcmhizzLreanc43xoKT4eVtpWYUMAdp7Bc92eMyt8uV
7jPUjikpv6qkYQEv9kQxubiYERol8j+T+5Vx5LIlNs8R+TVt7SZtFYUvODiR9qjN
vVngwTBVhOsADKAY8GTJ4ZfO8YjIxnehiu7HD7onygAgTDljT5BG6I47e1Mi9EiP
NcSwPYs7xAAJ+02EM+oqOYs48go99RvBeTSzatKw8ffPB+x+6TuHUdtT9j3aHycW
H+nMk3QUq84vL9AIYYeJrZvIoE9gH2nUlKX0ybYcHPgnkjn76A+BtRbvIZ4qHmws
N1ni/l1p/11tfC0x0ZE7AacBuMfbtBcalLBLos8pRugnj2F8mGNfzoRy5esJNfeB
jpBRQ91C2oAoMG7fvjGRRw==
`protect END_PROTECTED
