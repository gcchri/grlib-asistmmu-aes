`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bd8lvmYUmZZvAUxI7BVBY3ykmd4J3vtHyehvB3IYiwdxS4S2FMQr2rQ20PriNStg
3sWzUFSh6SgVen0isoBxRWuoxtsD/mMUYUwRKrXhOqtovnOj/Fy3pqsAdAM4H6gK
TOvM9Lci83ux3mDQjXqeEdoAT2B9S5Ruw7zKluWbG4GgywZLMyfui7Uu7G3R0H49
ZrL+l5QHlILQahZM6Z2kUOUYT4tFKrSRkbzmL+VVpUiInH1EI32RYrSlM4ZKl3eM
wjIWq/IQu5lIaSJkEaCjtQLQPny0eKl0io4+o2taPgEfYlpuVZMLIbp8Di9+1uSI
PW8a/V3hdgRykYOrmLjDuiYoF5XwPNlKwiBoOEqq8U/RP9oX7eHiR6BKZs1MZfLt
m2B2G/RrPqtq49R0uMyx2WlN8rpdzvL1GzX4eqE2in375OU2O2OPGsULAP3jSqhz
XlZNSU3kIIXVhcNPmnPxZHLs7K/n62IqYeVG42WrvJDYgMR2EUi4ug0vpM3Y+3Vs
kbYEMNcdlLV204JsSbaH7lUEljilS/B7PoY41xqr1NTp3YPu1YnFh8eYo1kIkv8n
C7liu+aHZkTQQiVGGj+pSMDh003puqkE3l+zQ4iLb2IDGk/OvGqMYxg2YMFF4qZO
RGOZUhYkudnnBMdy3hPWnQ==
`protect END_PROTECTED
