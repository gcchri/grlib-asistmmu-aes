`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KsfYCmh+lqxvUDlFQuMt1yg9lqDbpD3u9ZfnVU4dAQCSUCNh9PqCVAWSwAsl3ne1
x+aWauoaDg5wWpwvlNRieqJ4uRxQ0cp8dw2C/dhu9hNXxi3ScXh63chzEHsMT0E2
MaFjXM/Pm7wWrxxXZOTJWaM3gjr9oViLPC/2TCTqSeWg4kHNeRQGPokidGAJ6vlQ
dYXS/3+hL2ycDr5YvOUQMBhDYR44ZzDT8y6mT4CheYPhGudnYEvb9MKHo0RS5k1M
txUvS8BswoCA9Gi1x81x5cRi2o1qyOdRvH+4pF/sgu0kYAahLzXTcRXv+3YY9xsI
X9Q4P2FUqZVKxytgggt4BYVmmHBzr+SCX5F0mloh80o517G6J3qD3u7h9tu6fSRO
iffkJG5+XhKHKAkhhbBGBmm2R7G6BjhS2CXMpEEV0uqeO/tF7bvw4ziuY4Zu3rNs
kvMnHNFRzv6hKRg6KHieUQ6wC/LG9fulxpjZ5+PL8HSufORRANfLis4Uv/kPWnMI
xBdC18Jq34OCS24kF9Qom1PGalQhTIYIz037HE/LlbnP+fUd5q74Wv/Q9AQEVLAe
76nMfBVBGWNPaqQuGFBnX/bCOqlGe3PJbpL9+cBFoyNe/3j6VaGo645Bch+s0H2S
OnR9Sh91KtQBUqR16NYfbOeABXKthXSOy7Y0QYxY2mxM18nCVvVB6bqNkQ7TTzpa
mHrb3q3K1thapIsz6Wqk94anS9iyXNgYoXD65Y7NKbzPDtXdbwwG7NpxO9+EnY5R
voYr792iCJYIIkTvLP/yleDWV9E8KS5Nt26Ktu3DAfb/o4jGmOD6D4N8Jn4Z6yOj
cnHNXdmWIRdOx4x4pxMxgBo0/dFgkurIh7MCagmUBTE0UxQnL0p22Ri+sE++MNsw
jrS5EAPsJD/Fnn2isnZuN6Cx4fMgR4QSERReRwQQj2ZbDqCdGHnyGa9Wba9aiOQu
+VzZh6mZC6WiZpzgT9sqKCeHg6AnI4lzTd9Wb211Sjyk44jxdOmp9kYPyTa4LnwH
Tb3a/BMkxIdi3buO2eoMXOZdjhM4PRW03jViXKLebCRI8c0tmVsGs9zXDGKfohXW
XCjJejFcifD88lZm0urQtTI0+wq+aPB2TEAeepWHDklDEFBiUHrQ4rxCMdJZf9nB
3LNWv5b3wodH1V8AZukLwG1yWqri91cBYv6723hf8cc5Dc3FEZijQi1WUJtxixWW
3lsB9eIVJoj4DMZlSSMTnwa95kC75Lz2jHUbj7zspoROWaX8PDTcgaznavJHN8LQ
rQ+peXUCbo338So63rL0K9HWhWddHy+Qfz3WJAOu/Ol0gLF23lC7lmt3wyCwDWep
PEhZV9qTlthx1Te1DNUEj0wRGcIpimvxr09EY3r8sHOj/BpdwRRIm4DcevnTVvR8
hSHvpdWdUcG5Jwj43PEZsEqErynY/7DuSxffznKRc4cqk0fwXMXZzDNRIAn1v58I
6YT4eEqAOUmjy+T2MfVmZSRGiBBddwjpmK9qnRoNsdw1im7NOk9hBdjHCty7qtWQ
/I/Djws/laf6bpqZYZ4v0PUbPbXZguoiW8Bp4CYopfINdi3F1jmDaodYDunuZofu
G6mwsXj+jKcw4KACM9h+s8PywZv59gKS+LRY60Qilj/CRJBGeUmoAs6FwmPix0KJ
hTmM/WmfmdFoEHJRB2xs/KOhGOH6d/9Kd38qMTh29AZn0uG8GGZYmv/eXMuzQ8+o
Ch/0skG9O72N6+FvHlyr+M2THFtr4e61SZITY2HT9unc/fozoMFB2NI0xlUU1saL
4w5uzSnFmVVmy4VcfQ8xTBTcHkbP3huAiMpsJqOMBgvwVyehJIwCvNFdDboU6IpP
1Y8gvIH8QpzM9rwAy3wBmHWy2t6CpMYZPPsL+nuXKipEzbZhqfoJrwB5Ou31WL9o
A+sznat4eNOT2ShKt8TJjd2hAuKRWyZO4fFpcesh2X0nY8NbLzoAQaTzwUJefQY4
xTVImBIdK69iLPxroAEETsjqs0WNutqK7wc/dDwjMRvqak839IQQQFvoo30Lqk+K
NrzU1OQhPl0f+QlzYjmvPjy7tx6ZAt3XPvGhsYTELQ0P6dYb0+b4TXjDoCGa6xd0
4Pjmw4RT6oKcLB2huujcmdBtLM21nh+1r4svpWnvqzmhv8MZRBCg5YbGdQZ3mBom
wKuB8KLkCochWzSRGEDhIbnk20L3uU5GuA2gNDrYq3NeGKRQ9i91aTn80LHYZ7l2
gLHacLmVbk/ePfz3zGRZbxytK1DgW5K0qYtm9HFi6JuaXGEw4LkTMiUUIXMziFiY
p5tuZ3604mnsOxdwKz5BiBERRsVCftxLFEm6WIxgmBLt0DssTqkpSHEkiszUKHx1
eOGrSGYlB5ovgOoWQwZdFF7qvJG92tBlsyBZg0II7ErxkCYBfhuqIlm+FkIohw3B
PYSEsgEHNNNpBfjIkcmeqUU7oe8irq5KGkI8/m2KZ+hA8jzxYM0fiSPr2OxCBp0S
NoEBBletqyWn2RxObQnIhwSC2nOrdhvnZU5/okMXzvShuYrR+XwMhXRx7yQOvOMX
Gb3NaHE//nBdujPCZ2IYZaRwaDrRGjuc5jpnYfgBHinmhb3gy5o4sb778A+uK6c4
MDHnd/gvhSn3iGiu1mCNmc+VZJrRCQalchW7XZQEtXA1UCppDVMpYTpaUK26snpP
q2u3tqZCrOWSleJGiuPpz9Nksir5DLgrDwbZdsxb3KdlAU4ITDBvw33TT2ctsUDv
Z5IFlSXZeXpVOMHiFg5uoXFSdxmE3Pcyr5ONPgueAtMYfeDAoXthlcaBrbhowsHv
EKXMD7tt+7SewCkrigyrGyqF7TYEfjRU5cky2rE9c86d/iul7s/MCrzhGdPE2ihO
2GWOYaawrSP+Uey9eognfEzrZipQpp79P2JIBiWlz4LRFVwqazWXXHit562Y5xM1
SKzebQdKmpDHLG3AKT9mLPXK2tk4MkVAROUDkeXAhP82YRYsPjWpfxfG7NaseuOw
vT87B2k7o8uOepixjtKMs8bX6+pDOZsY8SZfecRdhCzNWM0Hpwkl+XD5xjVDe0Rz
7gE7hu5S0T/97x2JEYWi9ybeREbJNRQS+2NbD6yWcj4dA4bYYtzPB1BzOKpyAdE2
acQhUdRLKqCQ9VeT/bnAu1MkTrchbCaZVF8o3U3D5vWblZRV5h51YVBmcgKMgeli
YWTcv4EWB+Os40QJx4JWkc8SJ7xuBRHUHRl33hwwNYg57qX8ujkvfg7RGn0aNqke
t8bCjMIgYodPF3+jdZD+tZmKfGthT1LMojA2VQuRRcU9MCriR8eOUeAmRMrPsIhn
RYAu6yVa0WtpdwUjWOBV/Yf7TqumVbtkH3PXYILETI2WpGfN4mZNyfEeVVbpkHNo
VqSBNmogsiIk6FcQLmdxzkk/bAB455n1ozTD7z/RQHOkhDQrIXfctxMuAVuz2tBr
9/uz8JN0TDBeUOTDYj4j4qErMmi1dicH5veTW5FgvkflScbjwzL0eeBrfVOoBB/j
Y+iiv5ZBmssWtJqE1mu10A1vxMw08oxmQtXGgM7n+hfLAVhIKm96qnBRlq9lKtey
rvr0iHrSDIBSSMsmgXR990q31PDlP5G1cw+UNre3ur8bWKy0dnq7UgCWCsI/QnVy
T8SSNvTTsglhUEccZLZidnMTaTfWWHOwQJHlFukG3Muq5rr90mvhF8mKkpyXv2vd
8ZTZG/zUsw/bO9AMRwX3dun5G6FYiE5Ho7O9hvP8Srw8e4ANUH8OncOSKAffJ/pf
MrSDYsc2EVkPaSDpchRvaDbSUpcI5kskGudO42NHxiroWjAgFIvL5xsVPlsLz8sp
QNWUYLHKd/TgnVPizguajVtImJk2ggj4ToVKFvb0jxdTQsygpK+wbtq4pI+YDNUp
h+8+zU9Cm2l8VzGPy4CUEuBmpzRNzfZLABNVOTflioVDKgnBwpGxACDbS98zMRqd
qX4KkqQfmAjkdS6Vh/76xxRxl2T7d0rvTQZeI/dlIAZiV913lTTQmOLLp/DvjH1J
1sMWhSsxPETIgR4mt1KqfIytQyH1HCmRXbLbvssYDhk8Sg+CHh6W+T2wKiPS0jDx
61oKQnl4luIkQKpfo5eN4LSmLzXAWBARJcy/M7XcmpGRwN0Xu/kOwwpf4yNiSbkx
wTqyG1/q3dFaO7+pvNIH/wXTs7dtJHvAaXg++mUZleCdykDcidQ5Y68qXuzqaJg8
yqByyYCyERMC1vtwuIJGGxeGaDBDJ3BrqDOljwfDy/oxNEvmsqh4QGLShVU/Ww4D
MFsZPyqyb+P9VwlHO7VaqfCvB9OjZQPH7QlSDGEYsApnu4H09bdusHa8N1tEahW3
/tG+bMqpBjmCUW38xgtSCB939c83xDzqhuwmk4+/5hb50qKc0oPJkiQU2xBd8wUi
E3iZ7KE7k+nRJ6tz2gLPHVETL/qsOD/p8uJy9Xbo249+vZYZUWHRady/SuneU2M3
BDIgeksiXwbcg6oHYNlT3lWR7JA2XdgIYIvaLuTMS1NkWaxGw0TqbaFJ7YYI67+y
c0scpSGTIkxmrTK452T/gym/HozhewahndGk2dWGPgMFCV33ROSq38HQfWBGQklt
Qsab+ya1e6NnzbEjMK3n29dKXi0LKjmBkVmswl4ZNzVS7L2E3KiMZosu2ShpvYPb
Wx0fTlBYvamGM7hF/4dTP9xBl1d0/FqpqqBdRbSvilwRYEYQA1xpWH22KCxLlJq9
sFXm++b0JubtB8po9PlEjDkSj+rxOti7kmzT+7NSvDkN6oi98kAx4Guf40WpOrwz
RlRhvQRWTI1ZrVQb0txLVd6IHJHDIVmiTbpLTosKQojsv7nlvB2z/G8s0sr2NtJM
b7mzEofTJTqK2Bl5ZZfTXwhhHV46hFUZpDeSJinZ2yN0Yj6dZk/6qL4h0cEqlIE+
baNlL+V7CbDViYhj2Dg6f6vWeauZaU/43+N6xpQy5/bwDpLMKMu5VoxkNlCtdJL9
eJADr4UjMDIp+wHBoOIHN3KtDyCDBS5Ka6hwfqdguWUukU+2Xv25rRduIWV6wUXm
y2YLaW0URSalJc+tZInQpCJPDCG0u1Q2tZZnMx95UYh9527jeOMlhvAeFqRZFrom
herc+odKtFfYkZ1Cu2u+k8BdB9R3X6sfTkgqqgKXthxVcm4Pz3kYyZ57ntt3OmzF
ZA9ppRh91BGaxpleuwAf0TgaCcVUbbwLXKdlse6GuxL0o6VZgGJFIflfVx/fTdNy
cUqytcsI1fio9yzZ44y6KxfnTjd0PQIhwWP65iG6PD51WkZDCIo8+sHULtbBZMAV
4pG/nuhBI8TNmoUaL06x00BFSeMJT+rID9AOmQCatc4EZqGTojbrB4cFMrsgjvhW
Ktxusy+sS+VI0QNkxHRlHuOAkOmqf5WLxGp09uuOeUyoEMeiAcu4GwHmRg/g6wDr
JCW6Ni2EMw6/WAwq/jlSdWEJCv9fnSM4gXvqGM7zRnNAAREmc6dQAtC3nOFwxW2g
TUTSbxgtIuZRgCVHQz2OX2U1KXi7EtJp1qnEYh+TJ9e9O+I7uMf1X/e7BfnP+pzk
ptmKkVRoDg2v9dSDI4mFA7Zs+LhLIt9fJuTtpf/bIJW2nlROjOuz3QspZzoLtX77
5uSy3/lLMMwivQjHtpD3rZ0KFqfhWJVDAfVQTSVgROZJ2NiZM0lmNj6V/UH6D2VD
C0UrV5pTNhiBeCpPPzAAt/LUJERpHM/QkaYt11B7EWAzjXvDie9mXibLp99q2jjr
I0mUTAmeBlJtncDPNwc1FDmSh4Gq00E5n/E0gtkVciijEisJkU6IvDzOo+a9EvNt
ke1eXcv77eDjs4pgj1hfCCfDIvBOqUOM7o+LxQTVVQloVYGscvrc6zoMvnWM9Lhd
q3u/YDrOatFUa7bhDfvwM3gdenjIaaBpO+3KZlJtP1q5AEufirZ98P9+NtqWVYTy
KaqIihO+Aqs915deT2YJqWNVQWFeI3UqCGAoCUpwJM7V7Pw34/lPCVg7ifeXc+hu
kPu8cQXYj2Y45NK50suGDXbEtoomfy2vw5nH9WyzYxDuJiSfJwozT+MgLMKBmyt5
vodQcIrDPdH1/AFYp8ITcjtFqSJ4tGeLzSwL9UG+2kYSKAvJUsSbJ+UrjPpuJ50z
INIs3EyhlhgnivzHwOg+mkOTCvIMAvUBToTHHtbIMMZDfC83iyTzHkJfDovhH3N2
M7bP3M4+X5KQ/fmX5Z50MDKT1I9RvVmaFrFe72kdujW04iD7CzeSZVcG3AC1a14n
mL0+BgwRrAyhUvnTbKR4IKtFcnXwy/G0MC20ssrNPxLIvxUfKwHBq2qkgpqxvk8c
s3blmU9dn+rszi529SIsHvsjRoEh17bjm16r+jk1bJuTXSaOtOxz+x45fAE6YZvH
rMwsF0y6za+GaTQ0yg7dYZ0d5qU2X2ndTz6ysxxwZvQzoC8U8vjDaxyi95XlPyX4
MXveGNSfpGGytaWFxFHBlPWJHF9gYzMP4lSEjYFkCTb5B2IaRsxr/Fj9p9hWw0H8
UPqbAhPMJwBAQyoFcLRR/kGpwb8haS4ciwk7BSyIWQvIpZRJAdetnnqRz73pkSsz
jaEjU6Gte2CbPQocF8wRDy2CK6WfezqSkKpmSo23NV6cFMQiVFzaeqqi/TlVahvv
QIM/QYA5M3wtFZJiVvj0p9zgDC9YkjlnBpMhvzLcYNRxXA//8qo0v29s4FPAqadK
2h/ay3tZjhpwfSC6HglhellpXdL5L2lFW+gBxclSko8PHiZLnb4majqf1anzlx18
YoKHWG/5j1D9nbteSAfM26Ekf6DC+RHHXkEtKHKcaTKYlygGGpUGDzS9zDokiWWg
vXFi7Yu/VCuKxX0HocLGlGLTDdrHbJ04TSeuQRkSWFIGnX3n7BjTRN3z7M1f8LFG
lCVMN6YSKUpgGNIxCBmDCpHDd956COZDT+SRyVL7MxOxsvyXfKd2OTygt2l6IZqq
nJEYcurZNLzg2LIaKmdYQLuZ9j4L7mndOYr6rH085pmAG33xw+lsWx763kEx1mdQ
VyQVbVP4PguvFrt1VZYN7qvPufkO9PEuMihzVBnLr5GveYK05+/XORO7pP4jdmrR
/OuaKs7QFCJDd7Yl8viDfGJzbGFYV/ocF2FWyZ7MfuiYTWXYqP3KC+tpC6IhC+uS
LiiKlX913t8Prlpektext1b2FDwkjcEpmFRrMbpHAVcb9VkbfVxfMDDGUfm2uadb
X6z+YVBWhmjjsg8MRhzS+JM/DaF6AG0Xowj0bCro1UyB0+OKmbiNto9s6TCe88pF
eZQ9blL0XsEZIpZKmpgzbrLc+AavfpSK1+kUxBtOupFF6QweaURk2V8NNcJ6o3L7
pmHpTKVdrY9edot1uOXOK0oVK0AwcEnFwrFZzFAVmoCSx4sisij1n4OqJBHLDmxL
O7gXedLxVeo+moDBruHsq5dz3kdOAt2tbuXGX9nS0BT3lsAsDQYr+6C2xJW2+2OS
1fyHrvnyPx/jYGlVWz5keO1Sc8CG+Vma2l0vEWAtscueupI8iFk9AnVUgfTC+yH/
A8qmLegfsIp3mJmoM4nDT9ZnVPnEw9v2qviBsQPnzGHfVncMOSqsWbxtxcGKIC86
q0mX1OkeWDMOGJCw3zd6EkOjWsvD1n2yI5Fteok8p9j6eYMZZNKcC5up6Piaa/iN
TbhYhFe60pSJvOaWoYQ7p1EiSxDu7wDWJDohR1gfGngGJEjuDXll1CLcBHt8atdl
C9mTleKWI9CDkH2NJ8U+sOWVA8+TJkeAl1g8HkgQeA0/MsZ1CwUyOOZnfvbcveQR
q3KYpVtPa+zVC/TK1qOOKvbIBxrMArpY9+0sqV1pGPy2ko7KC+XAcJ7OGDxGzuqH
ildTflLVGwsE+p0MdwenyT+DpVfuPV0QLjDGSxCPaZoMcquNWCVsFdrJXOytx/Gs
jf8DJSwYJlDXWzKrS3BGDZIF+ZXdFU73Upm8s7xAoFFXSkq1yHdL8dO3te0fuZ9A
2QAnt5pXQUVGBYN3sBPMhhOVLYPEEvPKgZEDiCrL5vPOhgl43IeJ/zV3bRE8jWGL
C2JLgRrglUPa8yKtx+xTuCAqdED9kekb9SjmfI9z6k6SK8Aol8s2VryZ2cTMrfl7
/ToFQ88CZSArzMf9QUsP9imRfIslmRyI/XCLIo50u5IzgkJvp9IUmXNFnfyd4vUe
3DDz989v1+uoFDhiKJhp+Wad1rUYZ/IKYNpw6f3e7U3EaijY9Xk+0sBpCx28Tgqv
vfc2/Jw50LmNypQiNE5D4/I8i/xE55cOZKv5x4HFMPWfgSxlSqgB9jNyIM6WYRms
UxLKOGIFx48k/ago4+SfTaWdxm4r4svygTfvajPeNRmRFamhfdiiNSdQvcP6DPoR
SdKYW7hz73bTDcreBhJSqRWbj9sifbAyzxdiVqQJsNQJc/fMn0A2LbwW9Vo46mp4
4yYMajv0JOIj/iHp57Zh+FQ2Ml1ngI9N0bRnlEe2l6Ci5kAkHob2kl0tZNTS0Ocr
s+svKiYo/um6QcQGjWGOO2whGqZEzSJrGOFtphI2mig2Icm9I2eTD9GN2r0UK4qD
pYseSb+fT+ITkylJG0kXD5cGwTpwkoUKDqUJ0eClYOmKAYZRkCc0dsWGhconaAiI
jFAOoVA0bNy3/dK/4+ob56QriqcpgWU0Dfi0/gHX6Pv+kynfVefn5RPSsVBut6qW
qz1jAwMAvgHGoJ1j9XbAdXw7BS6f5XT7LfAlPvPPDEjjnvJl8OUNOWFZPQHvSYIi
FFW9OXV2u31NEcA0JG/piBu6M6k6SmOhNFNbp7MI20zpf7xOZDWS7E9XNO/te6wD
vp++hY9iwe3Oc8g2dFshKWqgNHKQprfqUy/f2S/P+CNxniGg9oWnSsl3rNK70MUR
2G/hg4EUwTFt8dlM84nyjA==
`protect END_PROTECTED
