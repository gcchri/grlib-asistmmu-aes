`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Az0oonW5FWpGdlC1Wl5tmn97K1OPj85xFx9Aa9gNj8K2Mu+rEuDdovZ0NQarRk08
xq5BpwMI/PlGEwlRDtVzXCaG2juZOAJGX5DFwZhYyRBXCrC+y1NWgaSplJdftvfc
YEpcTz7iLzO5VKlzovQEKrfQXRVzZoBOqF5rXGV+hL/oE6Vl5aLA3vZtaaWcKoEv
TTILSqvQJO7k6NNmVDjmztmo9Ac1Z/N7wYjJ4O3w6IgT2ZMh/U+wOqBpB9z4nsBy
md8ACbidN1VRp6OhVZvgzR6t5FvFbQ4AGIIWKmfcdd0Z6RXUHt69/ZmTeAGyVbhe
xCcXwHIJHa9I/WFPrdAeuAitt/pFzAHAjVrzlZrAuVvKKbnujsLFnr1+OBe7DFV4
dXlejNR57Wq+HhnGkT+qtzJ6Y6zK8SAIpakqJ728KjgnyYZYNpTy+2SzwcPweAar
DhgBHvbMt1z4wJrVS79YEsYUEvbDXqR9rQT1Jmj4b0xVraUGJwfHpbrR6vY/7Bi3
ZqWuL7d5R6hAi/JMhClI1NXCDuM8gwC+unkgS6f/yzDkJ4tPLepIVIBc+w4p9hG5
uXOdJvRz5NZW+3O6gboG71t1exOE+AP0aJETPMD9CRFXsMKkUj8jJ2p7PQp78fG6
ZBYC53tyE7CUa8uXYCJK+FGHxgjBU3OpszSmSvI/fceYQQ6V9ZLntvw6Z53LyyGJ
PziuoZzrfZvzZAkGGkxZwAFuKgkO3DwKT2lYfAvy72B3RyPd6A9/PejCDI3gpC5u
KQO+KXEfFuEBOlbjuoJkTQwwy8JNf0ndfazGc3y0aS5P10+k7eNG/ZbhfKqMkRfT
p96OD4wP7eHr7oKCvS2uSG0NFxHOau1ey3puOsbWhWOg9FEP0potso16tYvbowij
hcTq72ZONL6cx+vQksvX1O41Acw6mIDn++/Ij7UhDTWRjiMSMSPvc1P4Eyy9UpIz
6YIoaueDAasrX3/94YVBb9e0wVvX13Wu3Tac0EYXjcLv+JzhVCZ9VzQphhXE4uBU
ljwlqUO+G8prhrRErXdPxCsNYTTsvXdcoobZWJk7W5j7tdKrxPrtsI7qef/9+X4v
ZprK17IjLuxCjEx5caOJAF5LQZQ/Gh7TWvoFTu8WGoDrcwoVxGTvSbdUxpDZE/0f
pHsOlAd1cZlZerj4oU2IF+ykWSjcXV5rLBndNy0qaldgVA1QhuYKCpEY/626GPHB
+yJ5F5xUbcjORDk0H54UHPtpySYlBAGCraJoiqXXFUiQdO/EWjSCnrYnQO4Rz6oP
qtLtJSBXWfZbve0pDWIosyAyZgaY1Mt196JhAtQiipvnmaserQd1qwo6MZPj4puN
Bh2iesYt6o5KHaMw04x/8wqy0hAJmyE86aGkJ/8QWenyCqLTb2n2P4ILUY2ere8W
Hi97dcYezCLZTIIhNam2HpLYQPa1RCWJ4M93TMFq8hiRrFE5gIp95uYabftTvpfd
p4DTosqj9Hn/0WBk9tXt7cs0YIYtV3jCVWPr0Z4QRDQhr5o0NgSJaW4Po7/O/oeQ
8TpC+LRTG51VywmMBZHpK8uVcqiQxsHi0kXKrD0VVs3iDYlsSiA77t30PKEdTBc+
duXjyai2Fa1uOlrbIWVEkvzyuxXLZPnExn7ZH0Rk6jFSos5MYfFGDiz79jSk2Qjh
3ccSqIHFMQcxe7yMTl45KDg14QnjZ/4a9rCZin9VKmloH6vBfbmKv/RSctZhofOt
hDiDvi/OsbI51ZLd0get65PjFCRsag9yBLSh+/cgFviEK2ecUSFdiUJWCeybkxr+
VDsXrDsln8N8RggMfQq9DMYvPS/36iXyKePyqMerWvEfVF7xmxr1vHwuKQeKpvEY
85q2wQSIHomnvybmxkpU/od0fHI1abhR+PhTxnfzIF+TwtgEUEXnkzFwPEfbUA7H
zlDTIyZAnsaBGJ9w4szATSh72y7ig8pEzCiUSKeEccb/7xDC6mLfSUZz/DirA4A9
IHz387TX3DEoSVhyxT3ueD+3HXCGo+ZRi1CSNSKk/rAhS041NbP7y77WCu47X1h6
v4+HKUiVFSFQNbcIPemU7FcEfC0tSaiSBhPb3GL9FMNnYI1NF6oic2+AEKSz9m3B
NXczey/tAIVrxpGSKxFQLyb2Xsdk7amnYWsZzuI0kKn+rzekXjoMGB1eatdHaG0w
9H4+AxI/eEZLtQliY18ZoKvQNd/OXBr3jY7+C0pS5/OLhIu/MWGuY2HUWtKr2hJo
Idbc7NmAny53iSZthSDKAe4Lmsr4oOYrQlX6I36W2dYkeGxp9LmB/O0xrMfUI73r
oIcrFTXVPnDgsbQdScZIvVEF+Wm0YLaAzxVCon3oE0eocBFvua6AWcjCtO5WrvBt
eDB68tc9Fpz92YeEOTAWDD/TiXGgZ9/IwUUUPH/YecVPq3vVKuqXiGsmON699RY5
7mzCn44VPvrnPFdwf9uzHzK5j00wnsAZ27V41iUt5BHK5wfaTyfdppj/YqM9EFpp
fJ3UUYeqSDfZr5L+Dq7d1rOoO8oTSz4Q3x6DcfHqWhez0YZQSPdk4vJmjZjJr3Kf
ezHvK/FUaVSem2sJd6R5BKcdbe/1Ar1qQfqOCjPqcnqFbnxe98ERyFICDeiKSbh6
mEluISBBOjCZRObGF+SJYF6rphmEYydxdknDr+TRLvx2K+RjaIc0mfgeUfuU9eba
6VJMR4QMdW0JxvxDRohhBrWWtG6jiRYg2Gy24hoRj6fDqZWaFSL2AtsQHCQPs3ab
A1LY4/euMGON3BwTjAUqjLTXIh/3W1tsydqN096dqPr8Kl0hc6Fdqz4dvhwZb/7r
u0eJrCpDFvFTjJxxjIlg3cRWS2uRccsl/kyByz6r0y2FXzFdGeGfpAtrmOrps/yL
L/+B9qR8EEfGAW6SyzSSoxfkWqlbleVHhw/buSheVDx2raB/bEZs79Fh1XAuCJMe
XmZBy7vko8+DjtERGnmjjdrqdOxwAwcpOQx6cz5B8EF++wL/Uti65PC0Jy1oCdlm
Suk6cxox43LU7aSj2iYSf0lgID5xDDJswoOFDtfH3bBtVGkV2dr5Ysi5RWRrNzOu
yKbtQ0bCZkvPbFT7U96SA9vmqzf+Ahvp71xacLSObG76/0M5itpqQGUhVIdHVL0g
cL2n9VbqjPIRMKqESmXlbWtdOm0GvqyS2g8aKh51CRS6K+/QNd7MADDHKP0flsL3
hykUc8sYW+jwjyDJg+HccCcEulJkDV456jG0LDp74eWgSP/shithjPJkItsRS04F
UGqg8dkdbPsfhly5grW6tZ4R9zf9wpFFVg494R1Rik+B2ROSM+LxDt2HRFFVmGJh
V7HvsxZLA82+aeIXDlYeULqfXrBgWXiz5sdfaS61tSwUTFmX2vsxTSdzGC1/sJUl
90ztUFdYv7TL+sNbuBcS3A22+VYjfvSPYHvkDXzKbHYhxrb3SAhnwk5+kDcNWUIu
hOjZ+OHl1QiA5SQmUq37cpEwC9U4YKHJd9s/LkthGietuFzosffCG0FSgYkXjyP9
pV4Tf65t4vDQ81rlxL8JM2ODoLy3j4vdZvS88RcnmOjwvLvSYEG0DDpFxzXw5nRo
bFpj061l3sAnhe8KGzizv353HH9S5ZlyaZLwniKzzmrBKnRNn9XC5aPV/yF++Ao2
vtjrUcq/q5ei5/EB5Sol/ZB5tQKTGTAZebKbeTeKojvhHZGEi69OrUavRfha/uMT
Lk3wd76XjxlCNXPrxkiJl5lWEu1TROO4clNA2dFmaOytLQXPOCgumUHzB450a3G9
R1uGUeWBivgjmR8n3PWtYuxQ9kIUa8nYptJXA08cl/VtK4BF0fzWgvu9LQmWL5fe
7PwlXai+SxyRtEuMWxYOSzY6kjuPaO059bcOf83Zbb9FM0MVQ8SC5HxOjhFEkeey
Y/GKtjrKGey7NLL2CGaKF65YgMaYKmNaWFT47wnu280IwM3HdRJlbSRNXgn2edtN
9PMR3hoPi10jaa7Y6DV7gcADbLDrT192wVLqDumOOV2OjZkbDODckpi0AYPJuI7q
xPfvd3pD8xSrGnzu1dsD/UOa+bk9ecSREok6ZcwCkHp2bNRP6kv97nCJsATOVDgk
HQXemLAjD4RWS0pQMRlonBqgXeeWLYObegOOjMeLn0ZSfPqlTdZjqrtS263cvCN6
ETnQ0S8uBjm1dDlGbchKNtskzL9kUCdOa7Cy65W8eCI8KwH2MssxAgxxX16VlxP9
BX/64eRKMfVFjPnJFcjACYqIqmrFwmWMjjv68Oo6BE+5h3jf0QZ+KPr7dfIXp2wT
i6f8VwRRWBhcb14PFaa1AJDYJLY+Zju9aY4/fbVN3Vs=
`protect END_PROTECTED
