`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4p0wp5DU5Cqn6PxKj+ApDS3An9dBvw8hvCYVLbcdu32kzJMZEmOZUgtlABkQSOA8
ikr8FzBOJqtrxuMmbm/8iBylFBJaE4Skhbp80QylSyeZmz/B9W5dUVTrFWYBAHHe
vqi8mP5zyQEDdosapdN9/aBMAPQOasPtCPE017KO9kYwgydcLZ36rh2tNSwp20ue
9Uei8JFIDsW3kEogb3tdktQxtQQm10MbASHdLMcvz5gW1tOnIB3Z06gY9OC109iZ
+rgYvd13gjIuMJaZAg/cRTZNwaMnlYci8lT6G+O45RUPSg+yqv/STtlFK6YXX5cP
Ylg2s/LUqpiK0O8UfH0ZB7VfR5JCrKeQ8W63m4ixW2jCokSMS33HIfCdGZNgPOVu
isOv/s23jneTyF1wBT7B0Eianc9tLghCKXWi2zbPteG1nA/lhB19/+i66XoBZVYl
K9eCp2HjLA3b4nQtKbVXquKqVYWHwWPrz72aojxnsfiVl5cUhfq85jSckLCkWGc1
7nucjdumFYwKrbGlIHU/Fc8h6E/R/3BbGVu2rlyoz9mtLRdecfv9cYioLaMhOJKD
8CAgwUGX8UckAxd3JzXiWnDNx6tysIk9MBLUyG2LbqM5m8cjzYE7Qp5EzCaHDEJ0
tr9/BHB+4pGlG8EawnpnQsaRdujlZ6k5jKM86GZBn8IoUbmahuKGkM5BWOXO1Qs5
UmaD4j6iOD1nB/2C9aeKondMzcTPaONojNEdc3WtIFsLrwQLrcWPhI9y7wawnnvs
VUQquXWXhl4myC8d77cncQrqKM1O3ccOlYZYe6hac5bbCCEyu5DgnplvIJ/h+y3g
8Jsgac43Ve01hVfe+YqbZ5hZq1ugPa/qsbDS98gKfkXWThY32QXxa1jfi8dNyDF0
QvP8IhV4z6TgbItzcEHt2G6sAPy5IamUZPyAS8HcB4tsycPqufXiBh4BXoOvMdME
M1OV/Jj4SIHsTNf2x/g4YCpjvgv5lzFDAhYnYFymUSJglvY/eN5czRdO282SNr9G
5JvuxAS1Fy3jbAvt6ho771le4CpEvFm5FGOfgfSCtFU6uRDsw9M43++QGJ0ths6W
HyKAuAwTwYZb8S4XjV1DOGkiM9QPHBf5T7rnmwUM4xYX5za5MIBrnR2JDNOvKzA7
XuRGWBpjf5NgRVGJknKcxGMw78icA51nLLLGbHO7yUQEACzY5weRQF5iY7Nx54yw
oPMVM7jZ/O3/1BnwootnWeZYyeS6ZwBhudacsLlk84diXGtY9p1qFj9x0H9XCTJP
ctfzLh0+P+X9VrTr4X6X15e2dKcL4F0O49qT95VVi2K4ZHpavVPsGUd8H7Rnvj5x
T8rcIlCeqrF36k83cWwVoku7bDVRFa8Jgvua+o6H3VDkt4RF8ZFdpKqMo4FuMATW
faMVcaVtxjmqi6ds+/D57L1TLh3OQwcTtVBLy1puC4Eb1wMw/Ljy8yqd4m+HIlPX
2GUiYQqqzz7VC7erAXJBUlRVqpQrrcN6UIMrTmxtyV8Atj87KDcraEOrx8lz6jeE
+22mBAcvBrpjP3AvWVYgjHmDDF8qjuAbVP80J/3p/H8yOnpGFceW6MPJWJsRQn63
ZDZosqWI/vXD3XNv7EB/0NO7tjP1WkzfoekyfJwKP0ubu9fhs0EZKvZgAft/Or01
dmgRSyufNL9sHiAVVAHXQTAG7MtaSXOOyYmLxIScokZ5xiBedYoWGeWHAlLd3zm9
XLW9STZKT8azvO9X9khkG2zoGHbLdRHo+oiKvBfzGi68TUAniqNmRw2d1GJeH8Zy
WzJvy9/7mPE2VRSShRKxrWryy2PKDdQl0Tpa7XNwpiW/9jZ77ngPIqS/3zzJNmob
gUurYNLW/b405Rprg/wSaQSkSgIZN1HqqhRC05vfGRELzaz+DWvprpL0DoVhoEN7
2HT19OHIRtEhiR6AcbMoJaz08ODWeL5t+eXBO2g7l1lrvGquXhgSo0/tojz22Lpb
bBXiBJF8bk3XMg9DNZFz6hZ0wkvQ4UdrkiOnKVwzySMPmueOljRFMRYNNSVIuWl5
45EBFHEZP/GEd1l1Ue6get3+QByhbiPAM+PzCqrj22G+9zJ3b8DgUUkRGBkTSeRw
0Nit5KCdF/jASFjTgVys83I4UGffoe2u6tjFtaqWiMQMZOCiYgXffzq0IrYhQcMz
`protect END_PROTECTED
