`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rCTfXB1NhDY7hekAiYaMu2zbjBAfOzVlcHSfzuTeVzruxYzNdpauADZgBim155S6
A11wYovZzi3paI3c0asw8GiWuBOqm9bReVpEf2jnLNszkybIxUuf5LXanuLrseAD
sv/NcL1ioh1jIgvl00Gcw1AQEmGKmiszJFtE2EvvsxzVzyjmW687RTMGgg0bgtnq
Dreaygeg6DtTe/gsMt+H3fnXtnx2tkd4Joell/yF70dIDiUqh/Pbeys9WjyAR/4S
sL++kFe4Yrzlxa4XywnN7/l4WSjTfGYZzWrpDLEqQKwVKFre/IyU0wBrD01bpJHZ
F8C8CD4Q6l1n2Tfdz3X9fSx9EMQBMDkgedvfhVz9L3P8J18lOQA2DuaGDWXodZdo
Tsq6xRXl1thEN2F8RntR9fNKTUFbpcrOgavu/tTaYcRLnPoTjHBWlVY55j0f2Xxj
Yl21c7LphOY/2x7zw2aw3x3KrecPYu1P0jsXbgMGNjGLx/uKG1aeTzCzMLdHvBzL
eeWsmC/FrwRZbnCLjAH2QFGEbP/dr77PWOwWHnnD9kHTS1CnrBvR5U2LQzg+oOa/
H+PkTW7sNrrzf5vxU/bycJ3W0MBJ9YfwvvKNIbYeDDc=
`protect END_PROTECTED
