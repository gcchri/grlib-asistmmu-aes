`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ARgePNN9y5uUYfgAfOm9rCy7oyqae2fiA31HYOIsFYOWORTSDLxTHcoLG9SD05m
7/6AVIVgXAekNdbadAQ8B7+BJbRumuLzzTSnL4NO8IC5nxBYJo/Cv5bdcTTNoQLw
5PQLGLnmPfycFzmolihx6SqYh+3NYd2HkjRkdkXCWImR4wTv3k2hVR7Id0A4NHMo
6M8zcxlw2Uqv0HooxV9MnBY7PtnKEuR2MUhW9ZeFQ+VI04N1kL1E0BmNjf+h4bj1
W6Uh10Ak8nlMn/k/OQvHWANx1jB8wgxZR3B5aXL7K94+MC1C5KXgUmqHBid5FMcR
UE5w71ADnegZA60FnlhN/8ezRleI2SmSu0SOFdCGkz7/nzQ53TVWegQi0fa5T24q
gqV0ufLA7rkEllQRTs1thXA+2GTW23xmxH14HUXCMoSpBj1ndpOTZpIObAkTiVHw
aH5BhDHyBNYtr/wheveRrhQdgGwh8rwUdLgrv0ObaL2ILWoysNSE8kU3vQPsZkoL
dQYrfShHJKVZVFvcB/jAM4qq8Obxw5r9UZCu8kZ6bQmye8yPt1LbIPzFbNRDevHs
5R8Q/x3PyIaZg/1JuCLHOSqH/tUnxsiz+GEhctav8iZ+ndAwrKyZOkOPyl54ZWwh
if/hYjx53FxEFWyjGs6jDcsFgnRsuIR6cihNJVDF/22S65q6AcpsKf49zOj9cK1o
0hANr35gtA3gzHHsZJFGXk3vf5PpQWkHLObQ2abu+REMy4bt/25b0DwnKcx/aZ6W
zM2TnYvdFD9M+Y5HgMVfc7ZsA5HGgJ+ogMZm0ZkZgjUFpAKrzGfnKfM0zBXtlZBO
QZY5uviaQHebk4xMuIqSWdQQWFyXvrtfwFyI/wJ/xWUajuL8KSN1rRL1IgmGdoz4
R8XInH6xiarXRMC7qcCoDzmzdUkk7GPnkE5VrBcNK8siWPW3sNYYLYMDMrbVOI4x
Qe5aURgHgOmRGPYpUXI5lG5Q4I08bWRQjXY8fj7hNf6C70Iui5rLflX8pUjpUgKB
zkhESWa3EIowAcpMgiE7QC1SSXH5hp/62N2M/IPbVcGHGOzeFCsjHMs1M7LDzLxj
0mxfces2fIxu0fKBYGsZo3XGsTHEVxGhmv9bw5j7sW1Ycv76KR+cA852bxKg6y61
`protect END_PROTECTED
