`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c1J6hTqj7vh5YwggDfldKvf9VeLLQ74rGhbUyj87+CzCpozK0++rxjiCDYDOwNf2
c11UDU2d0xD7Q7i3HRqMSczLZyDRFdQt+ASS6mC6q2/o4tmbhTWUdkgpDL3Or/hX
it0Z8TvXUiSvdiLhNuGyua44JC4Hug7iXRywJm0H6FCqwp/I1LMWgGBQ21Fsc8jX
5TKaWN6wjOawzPBXJc1/CXZ0s0RXC2ZjxVyef+Ywc6CqsfGC+m4uAjnCIqoYO0Mn
Y8sOpAi2YgMnpmzpaCTVuMqIPR1wj/5uyjAiU7lyma+zuA81Z7Y+OEecl/I1ZXH9
aNbIaPo9qDle8Pim2RzyTG09HyAeav7gsZIXOtK2QuIJzBbNuGjFu6dNGRq3gRdq
I54xXyS63SCSAY/1BILUuHzohTFmHS1JO0/Ih3pwsx0=
`protect END_PROTECTED
