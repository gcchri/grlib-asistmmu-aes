`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
21bVWEfugrJGQnHak5vGpDPgv6DqDWz+xoBkGckhndXaiVGKl2Q8TxokP1+d88Oe
UimUzhSaCm+6g9vj02xyDPuFrtUGYd79MSnDvYMrf0hn75jpNur0UBWTT06hcOLF
TDiKgQ+T1q+14mQAjVpEnKQpImWp6a1XZnR8r87X/bRR7zy6FRzE8eJbTBu5yhlP
H0+akUAfDN4qJ+suYmmIo32e4c0Wctc+/+1gfGSg2jfw08fTR7v1EQcdas0Ys1y7
hnxaviTFrcR3LyzANcOiOOmKxytttDP96H+5l6/Nro9beblUONqiFgtu5VWGVJLl
cAjtUwn8rCKyEqkwrw48jxIF3EW2r4p6M4NW2WNgbyE2Qs4LSV8YaJ7x3Kpl9Mli
e1Siw+bdxh0oGo2Dizsd19gp1S/gImA1r5lpu3CUzrI=
`protect END_PROTECTED
