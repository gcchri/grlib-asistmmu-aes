`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UubTtA5Pws4asEKv+UUY+IDKOXziHgdkjqBlyVl6VTZPWhzKLy6nITegasLYDPOp
tBNvMgPjYmVspxWWOtzM8j6U98t6jyM6fVqD59hq3G38bGOjZI/9LAQOF78JOQmV
AwTI4CzCQOKlxYcqRQ/7XUl7EbrPfeldqqUKQkhwi5F5rfG9RYTn7+VJVqgmwGvQ
xIEnEyYVlkxri8vRKDxcm40l0ASKKdhKBsuKSMsHMNyMUrBR8MQtNbb60M0+iIYp
Y26UFolBugTxa+8W/JAwwKI9LuirYOqlTtAb8JNGvslJBvHTbuiKCB4IEY2OPtu1
+BXWYGW/lsYIcUfVjfCLr6r3KcDO22CBN6LZ8tnCr7DslcbBlHyHplv3Y5fcj9K7
jgAP+nTvhLI+2H369bKE+u2zdNm64z8CgP90AZbD+5zBgMRff4YRwyQYRe8hvRY7
lW+i4BtZyzBB/lRruvPtFzAczkeLQ758ucrIlfTIUO0=
`protect END_PROTECTED
