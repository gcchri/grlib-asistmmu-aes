`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fhtedu6nf7iPyJ6xwsi0gkc+QJumjh+M/pFTHxR8A7ctCeunSnoGlWnyctIe9DWQ
bXfltUccYvL5dj1swjucVpXzpZwb74daT9DKrxBilghcINE8R5bg+bZwuNhMDtjx
RWyiXJ8j0zfVaHKTpx0lLSsP9PGHr5V/LZ5oT2Zcz6+q1W91HfUY3tP63RDBttRb
GIyb/B7fkiZE5CUrbjTjwIMCUYnsIy4k4bZHTa3RjAFzYYb5bZkTCC6Cm8HDuQon
JVL1m1r+r1K9MC1/3HUOugCprJN5uEfPdy/GEVYSYZoEJk0hG2sUxPdylpdZMW3p
tIxhbjoUWsZfQfLm86VnvR7sAqFdkTEtLNdE6FTE1PwxReHLPjkeDCKqT+QnjFQq
3NA8nt4j/3S5yVsSok2sDSOcHwufV86WO4wTodGd6r8=
`protect END_PROTECTED
