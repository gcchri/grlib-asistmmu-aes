`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C25rzjVXaCuuJRDf77LWw61809uMKzaYmkcvEX19TDxzUYZ74YIlnTfyEDx66+/R
le58AZ0jmOU6VCCAEIY6z4cZt39cWl+dwh6mDmZCHoVPYZlWcyzjIZt6jWDccPnR
d4h+LaYLfg/oszCQYgT28gQHalMcEup5UzljG3MUvIpvhzXvYlOS9RV+WALTxbeh
p6Cg2zHLBhgM1Uh658zf6gvqhN6UFb8d5buU+SO57m/UZkitGRkbCqEsuL8i7IB3
x3/tSaYKgM5+ffal4hon3Z9X5CQWRsw/ccwGc9BthvHXrVQ2BnHqaEUb2izFLAYE
ltTAdSFjC85DCGYUCN8Omg==
`protect END_PROTECTED
