`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rqnc6ZKBvpxjo8IpAB49Jj/ixSZyOYtveWnwytgspz7vtHY3BModE9dRHnxecO8g
PdBXx9V+C8+cM8XFStQW7O3I3I3Ithqpav5alQb5riObkCxh/FxcoyM5elnct7GS
0BXj9DC5qqLH5BsEgfZQeDFCFfDJ7teTz5Yxdfa43/Csprgp4p+s4Egb/vun6LWe
g7WTOAlaMNuOZbyclfwGAnm1qgXapmjytRU1h8lcE0Byh6EF0Np0rwFkezNeUFqq
qWwR1U6FjSfbBqMoOpE9rjB/ShGsKkZ8q/NEF/25Fch/EvqswN7ERkDuU6U4+Mv6
XwAwqDG1Bl9zvlJRT2W98Q==
`protect END_PROTECTED
