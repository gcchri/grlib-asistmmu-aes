`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N7ay9BOajrxhAFIps8rzoDbRxCf2ibVtqKeSAZyZsm4YLA1ViEDeyxeoq7n4T6Po
zAY+mAVFXbyyUdAjLGMGQXhNb7oqyyH8qykel1jbbehaHjybf3JZk9beJuONdN5o
MrtdC1y0flpYwxKlLqylmEDc6t/ejO/8gO1aY/hZSZ0dy5yLOn6hSO2wz4rzMzHM
8ySDI2tgSwYP345sAPx56wufLPSflYvy5bLUuXbAhOjkAOOJyTQgihCj9RiNOgaK
NwmP7GbdqvKbwwBA+kPcCJvaBDk2uwbTFHy0X7PKMXdCDwdPdcqzuHkCmIfHDvlm
oYxvbG5YHrjkNvUJOBkZk9VPLuRuR/JnY6bVXYN3fxesTYLT9LKaIT/2RUN5eaEG
YBiwoi8tYVI9sgK5h7Ryi1WFC+3MllckzgAhMMWobsZcnW05ukVukWzG4P7PpCMA
vkiNl4pw0mIkrBQboVfvYCDJuJzsT8IXTVM5GQ4E3Ci/a9hbGbdD8NOeff5cJV41
kRMoh1ekCR5QBtsvrt5rbf5IOM0bN81gVq2a6W0N3esbS1w+xq+Mbw6RAUuKAXWN
MEb0QjcaH8Bl6nlI+zs9xbxye2ewlagPANZIQi0mUsuEge2oj6Jrli1hdYamPQPL
/q4C0uCW6Y1Y5Os951lQf7r03pUrRY3kKdpST+HKyc4gspEx8UOG2txeVGKqeptr
Grjhw/ssL+XqhdYd5AdCYVd/iGN6MOo9kBIX5RcQAwJE57l1Km2DZVNRKumwwJRq
l8UYPdotlR5+g5atLoD7H9O2PkPC06Lq48M3i4Ct3zeQhWrzuRhzfSNB5V4SIzBz
k73Lal2aAXrosUoC66+GSmCUB6dQoxKnBP0FldlqchVwLVXeER1ZlkZIpKL6XwH0
NuAMwZrQ+3mpn77+ytekpGi9LNvLofx6ZteVamcNQLP6d6wK8Ie/dW1ddoLRrMzc
rgFR2pl/sQ0EkWS8tQu55cIiggeCqCVP5wOEPOpkv2PIG6qlS0cq3Hs8QqByu4/9
iY/hSfg+5lDes1OwYho6NqJoxtVVCFOfrm2Bf6c7BGRXMqfAqQsPs/VpogWi2BRw
HWUlDWnrQeI16yD+hAu+f1F7xOU/OFdDO3QvdOxA+efT9YMSoZ3mAt8loEw+8K2I
9xZU66asNNFNZffNJkKu+JU46KOZvL4OrcKBi7lbiIV7XZE26pj14PwahZdUdqtl
LQw+bpnaIFZ35j/9D10D1eE7ODT0Ry4be3hJI4TFXAuCvqUprTbVHw0I5uzgbJo6
uYWSf9WA8DVgu+2QPHU0IG+P+lDaP2eb+H6i2gpnuYjSKkh92aVZiUxKlvHfOWyT
CTyTYmh4OUoRosfWbO1nvA==
`protect END_PROTECTED
