`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
noDlXTPrVAy0p65eVzzeAYZOMhvxjRkbeAX3iro4amA9xJ3W5aR/X40KuuygCiLm
dMf0f3HRsxWVSjYs+p5Ac1M3zgbCqrIegQwm+NWoAaq2s4Xy3KQE5R1cQikhtPdn
W0cB15VdfvDeoGuuWfN3lByYSSiDfklWw7PeZSMiMgdWHZIPGjqrItC0AvQFy4FR
iLBX3INm+UDa2wf3uQeTLH2z0DPOs8a6Af9W13ZtaQHNER890/6CV0qvWvIv8lcl
UluUjv/YSDj3hAWaXaVjNVzWxYMHnJ6XPlFkUEDkMzMqq1QUpsLOb8oxElhsdaGT
n3g4tHILh5287PyrNjGjyfDRO8GtqLTqIPSQertX0Og7GEfBxBWViuJnoCyYsPdT
Udzn2/IgdTL2gbdbf/iDF7ax9nxpc5p91LqP/+2fXKy5qEpntIoskGpDgRk5U/lM
/CfaMAr8BbX3hUM9sI5cQr/nf5oUl+YHcCQtgLEQBUINo/TluBBoNztbmZs8JjTT
`protect END_PROTECTED
