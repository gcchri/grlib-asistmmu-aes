`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pnq4Q/MTw11t5v6F4mwDad11aJTdDgB4NIvjzvTA8SroSwDpZnqw7R2fzM2uDn2w
CbGAtSUsuBQiqq+Zd29jeJIXz9MztOdgIfTz1K41lFf6oA3CGd5wnnrGWJ8Vm98j
ADLV+QL+OPfVh6ORiaatiEbYPC2fWWxVZ6ssHp/ycpNCh3rCk4L7owRvD86hIrE9
wHw8mwBK2f0tPlItUwS8xIyJc9/mMe2lb70Sz2Da08U2GXlC7SFyDmW+ZjEEsSdF
+b+EqOE47IsGMjzNHG7TGJQppMmKandjEnSrdcseQo9+vIVr2mgU1UqZCPTS9uqf
zb8yTIUsQOkfIUtecd16TfbtwtUyumkWmXvnTt/oMrrauI4ajkMNt3u1LJGTiA1/
hC6MmpRIo7zoNY9n1n6GgxP8Hsho7JnwGFsey4N56shixyqGXSKJVlRZfa///5p3
bVnj/6pJ2cGazlRpA4YqNWWo5j6WJ9cha8kr1RhgxWQ=
`protect END_PROTECTED
