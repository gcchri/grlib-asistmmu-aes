`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nSoYbDFodPHMfSepWVn66qjwifrD0b9Lgs5wQ+1/sfYa6U+2dlnYUogGXuwzdB4h
on/n2+je8XgOoqQ7e3Z2KL6zAGHE1MyRoag7ipirwIalVT91ac64WSotYLeXUC5y
072pzcM++UEUySEExabBbH0iF06xlvyDhLwxybuFw+ZOYfoHD3M/usoX11ujXCtr
qTeS0rEeAbT51WIugWBd8xBk6LwBPhSvnFmRtWm/Kg59MEEY2yIS4NJQfAKwny6f
5eCYJ41St3NmwJ9r9an+xGgXK29ik+staKGZu1d0QbLjzmNE5/WKx+Uqs6q+RsgF
`protect END_PROTECTED
