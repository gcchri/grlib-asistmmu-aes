`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5yoQUQI3uUXJdUW9Mcdq5C+JP774gicyTEiSPEpQmjiBJEax4qWz0zugkLRcCD6C
+r75Yl2ZGAlijXOfuwx6tgrziLF/cxq1roY7OP/ybWKZWxBKtDGWsXJeB+OQbP65
VwBCRNijotD1IM5m/FNVU3G4pGpUneStsGVHCTGdfffF6MWIlGUgg1XL8wFYM/nr
z5lGqtCBS+d9gjormSFiqIlsmse8t+b0z1Ye3wsQ6W5qsXmZDq+gv8Y9MT695Mk/
UnIo/gUwpNn0At13RjgwngGjKOlAXr9dT7Wg/gzAQuPOLSTGCQROI9xcV7yS2zn2
i0afu9uyXdvl12LP/qMpPeGWqbOYGiVb4Pd7PrTy/Qyr4f3Hzy4WFGxckGKXpK25
sK5sR04txqtYmwJ9CRg0qyTi7Tz1+ssY2Rnk2lzmdVEsVTUMj/1DVatl66uMIzL5
H8rd7sK3/Sq8LjtimM/s5lVvAdEJqkKN6a9J4aIXNdVOrzlcwvy0eZ4KoH8i0PIu
`protect END_PROTECTED
