`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sYBnR8qmGyBLaC4GGthwysp9vqB3FzkLkCcStIN+CB+slPijCyJgmyShzOuKLo6E
Gze0JlafJcJJhe93geP+X6e4X+mrAqHdgzhEGOPh4tNP5qgSm/Hf88OpVUeBOF1I
kZXxD58hFQrDXBeSvEj9ML3esMoNuHV1NLOaOLTUUTbxYxWZUfdYQknx6Ma5eG4d
AkQ9Riq0QjyN6gA4hba3XNwPUyADC5+V4gHEasvfnrDggMjnhmxxkIdEBXPPXNUy
h/HpSOhekMdWTEZy4oQzvFGWEEhJPhJWgx/bdFcLS8EhJw1BdlGY0T0t2U5w9zct
yw8gzyaLiwjRipGLFc0/gvOZof5Jw5pYyDYfOFGkWR3uzEd4dOFt+NhrIZWMKekD
fEMROKDNrH7y6l1++/Bq5iMPzDVAle0kqc4CmjxkNR/DkWTclVPW0ieqyEziYLQK
0GmPXRL3U3i+WUJvzWF/h45o9pdLM7UQa2NQAQoJ+P4=
`protect END_PROTECTED
