`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RaOAQGw348ZCcCxe66OtwsCIuFfbKUsn9GFAMFN+4EX4LJQULjRHWU5GvU23HiDY
TG8vBBdR+CME6w5cCttvFz/INTUnVlavHNz0wz0+wq7m3K4/IVs+omHEcrhinO1f
jN2JGzHpT+7x4jHlCdylYfFr40rTRpds5rwCjJe2ObGi4KNT8h6LFXQdB6ayasEg
fQs7zAnvIg3UogBXgHA1Bk/UQzEezPyWXsrG0HoRYyo6WdiReCdyuBiCuAlJn95u
ng+9yT5pDYdO3eQGHY4wuDyhnt9pvWjuxpX7H01xkJsiaOh+GpcHcqfvCEhSi+bX
A/R0k9hBgjE8L0Lc1cAijtCz3lInV3ry/YEqQW0yNQo81tuW9qporX+neHSeA+qz
bdBtzGJAuln3+rkCc4t6mD8ayJyWQmGq+pEA2jhJOOc=
`protect END_PROTECTED
