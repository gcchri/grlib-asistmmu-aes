`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ykElKiKBWQmkI6mmLGsmxy5TPoATs7pRHoERZHLs+oejQEA7lo8jgoWQAWU6E9ma
Brz2QGBpocmFLhj42fLH3JfgFHrYZSKLt9u+NnXXLNHkHEHiSSliUOhoVecQz/Ep
opR2l3gBf79g5C9j/ZBUpZItaQRltc5cqEFPdJeI8xxF8ZwA1N+uN3IK5sBWTpnU
pSppSo1SvGPn1ifZEzzzs1QUlJTeFLAelULAYiQ+Bx8GF9RdJV+ucF6GTTaJ1xUI
HKDyRYVzzfGt08SqPnXFWeXQ840lhK33xQtETY25IL6+92PnnhR7AFPLvx/Psdoq
Mue1MkDl3foNh0fHc505tim8zq8rAh0z9nCkLOFPdq5wqNWEpycBrTZyW/6jgzXe
ZKmVg4fOzos950iuAYMCDQr95hF6np2v+WrgF5j/SAwDRHFkTS+kbRJhakMXwMkF
e/re8nJbAV65gZo3/4e9HHobWQZdwOCavsXvAiB9nn0CRhnqIEoS1sCiGqtRz8Pn
g0GJZHhqoM6tpiXvbyocAw==
`protect END_PROTECTED
