`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K1SEK2/Yk1KRWfZWO6gWFw3lX9TGvm93Bpl9761W3Cv3a7kgTZi0E5f3qGXw+ul1
/AquA3odGxpOsVVMDTDoxHKpIvKFFnQwmY0Hy7crnQnDxZG6UayLznYgKnM1X3Pn
d2ZiL01qXEYK0avdZrkurkXR87XtH9LmhvAmrhqk2bHxpNrJccuoF010v640ku8n
5/7Oy8/HhorljWs9vCX4qegHdKRfE7WDK+3VKaR2iYsaYB3LfKhxUTmdLT69tcHE
7t7CL+FMt08HvKQAfQA2rUFGrkMgdErUbfiONW9SckjIbhqzoFUIBcpicKuTtBHA
0KEibCfeVB7JcZxUnclsH6c2MCTIqOKwshM2HuY22AoesBoTgV+ZNLyOkCTREd7n
Sh+Y7I20GLGwhkKPOc0QiJQrg60BkGz5RN5OHV2au6w=
`protect END_PROTECTED
