`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lMPlGt1U/3zpzQOnhjMH/XGQGm+GtlzXKGsIfA/UiUDylw423YjI+EB2etCfFLTr
aZoXxDSEq//SuFuZVo/trHquruX4ab3/XEs/hcmHR9N/AyYb/zvfWdhQUdZ0crNE
cWGGDWiPNWvXdshDasrn9wyBucAL+lL4qDax2RpO7zIrUB9uK6IB/2/pkM6aGinX
6Pwc42RfKjkI4bPsWO/buRRUbMR9jusMNRkO9E8mrRIXBFpO6cqaXluaFZgX0QB8
U9xZUqinqcoCXUPbC6HLNU1dJxB9vmHFt8B0ScxW0Gi8Dh4dxmtEQcjHtDGI92aq
8EssXMeDlwe/tZj7bK8sVUPgz3N7CY88nLhzms2qaYAOe8glFbeVRD0h4jUWE4Z+
nkbQcteEKB5Zft2PrXi5izlQ0LFUPxpn8TByTYTbmKY=
`protect END_PROTECTED
