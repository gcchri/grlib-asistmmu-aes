`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YmFUMnzTvMkCHZ78OPZ8HFJEUIpVUUBV/xSp2z+EAG2Q/UrncdFIWJCCW0uR0ylr
x8ap3yb7MGcD1wjs4gmm0scnDS8JwoUi4aQWLy442Yfwj36Q7B8sT5fyybhOMcG3
x1ig9Z+D3eNw/AHznTRDnzITo1uX+bpuDixm3aEDttSJVLydGHBZr+hj1/SOY6Iw
j5YwOSBoCkDRzKrcQ62/sDLF5ON55pHlpeTQU31kQgH4/KxUqwDK2LlS/lm4uEwe
y0tp6KuFuUxfvMxXH7dFtVcM+s7USc8Zmh0kAo0iFySO0JrCkpvkT8iq7R4n0644
tMxP55XE3FTM7peF8tDM8AMCt61WyaZ8dJr7bEWuavpElKyZyZBa76TcTVdm3IwX
uZvdCcBaCNNdmUHvGjkTA86svl69Cp1mGAd1NCwAjdfYDQFSkzqq3uwMgL9k6oh1
qrv9iy01A3oeMX487X7wl/AeOoBJn1a4KPvwwg9PnlnrV6jr+YZhXa/TVjbL5INf
78rAoBG4r9dTCu6g0Q36A/82oBTcfBSIn7Fl89Spjcn3JwqcWPZQxU5kJ16w7Sod
NRLbxUV61umXLYUfz3a5Pp2BWBn1kAI3JqxqLT+EjJoox36A/ndyzjeQuGjsIvlI
FsOlCnyJxm7Nub7d4yFQG8GMu9uj2YrqDg6fh6vVwOL4tN5OJRYM3FfVUl9dt6Ic
7JMbMxggjpczmQllPJRCV5e5aUmzCo6eX0oDRF5s1XTdpZKTYZznfQSNxjklhYZX
XeWjHQEczDd5/S0Cru3MUGI8GG2csrsdBLQwduOcpN/J+NrlMhQfYHpnsT6JteSM
kYSRjUumaS5FISpemzbnIzJHWCOmlOQoMT56ScutvLj6P+egtfDm6NIXLXs1yG1J
GB6Z1LQSsjhYMknAW35XDG7xhKa9Q6U9WgqKoe4ayiKkiHWJMrXfrpoZ/7Vw2dV+
3erM51W5ClZVlqHLqDgClBomRqlp/JLSpes79VOCG13gahCuuznFi9VV+ZhstwHK
ZIhglRLbGwBYsyLblhWslL8ZDyzoAJgHsMiYdtV1OKOpUkqJ6JzyBKqMeDLYCAz+
yKY4m+odGnPU1BE1LK0x9DbfWXVg6x1O9CsURNjA3KYAkYCTcjvKF4cBh+efKcp+
0kMRykYhYGoCsKTdisDWEQ5kaveKff9BivbXZgQHDOa1ZnD3qsKTOM+Bwc31l4h7
fO5u/I1k/Bns9mSKVV6EHDI8HHj3D7TlgNqqOtIq8RZQULLd+lLD1GOBEpF7GChO
k9V6RL8j29SDbdSzlp+PfoSUuQWAzPyQrLmQ5O0olChzfC/br4PXkk4m4ZvRRQAb
P79FM5y0pRupY2gMTN2ReTEsViRRWmgbqc8gYsaRjyGRG0Fn3beJ2xz1JF4rSfVS
Vtyce+dazh8BpHcdhuT0bqxCDC7RYdCNWk1nwumPmSQPg2XWQLjg0+yCcXBQAdT9
kL+w62KpiFFOQyTxjx7QdO8kl6xDUb/52hGGXxsRD/3XxJyeDxQsRUmavdhQTV2T
mcd3oJnStqDhk9Q9/OcCev4FIEKrK5ZUIJLmbeJeKvhA8PE//8DBIz7AGSu9mnrO
pbGlyPleTiajFvcmefh8RGXo3NK8434anPTKc3VlyLPuIUK1ijmp1aO76UkQjeeX
MKrYNHwnkhltWQlu8ioRf3HjBBDvDJi3vinubtVxyw6YiAvo7svdr/u8WRtMCAds
aethzVDZsmYa94CHGDz3NK6kY4T5DEKZnafHLEvZJb4hquTKElWqRuxx6YANeTlX
6I7afbdmDxTIzYPK9PL3XZ9TqTkdpY6xrMqrNa2+54lxtpS+ayPpkohu+Rv0jEIj
Pm/5nX2GLENUMl4TGN20YeSo6PLnIEgNIkcfBTdJRZXzpJax8wpVeVeeOGzCbORk
yF80dDPCLEl+Q5POUDNAWbDWtl285fPULxBtVGeksQ25nOrqZk2zUgJFrs5AYOle
s13ODRIKbwFbOSFfpqaT0Ib7ZFCuHSVfxxfWlZ3Wg1eNQfK7TRn8UhxqSuTFb/0v
IJzaBMXGBQYPOFwHHnUJiKmDRylSGp0jPrk7qocaQzNzGnaDx4pFV5P86UAThfu8
vOOvKmv3o15tQ9vgPemEwiJnSFOBHSQaCARk6N+MvtG3vMuU7M5LLfpb/fj7GUdH
7Iw3M0s6zEeasts2Q0aqJKasGMw56DGI69Ph5ZL5tzQ5zgFe5qckiaczi295Qw++
Qks2n5E068Zz07FLfGTe7TkMfP4YsHd8Rl2AgM9KlMLTYHp0dMZWAeyweAFSZ4JI
7bb+xdyhNB4C4ARlhh43Ef0feplHo/i0uNUh2J11egHzDFm11PqbIX5/ncdlJtr1
qvevfXso9Bl1a1rXN/nnhaZ9oe3d85ajcN65qDFRnmaPUj6ypABFFsn8TApce+5F
rZqjdrXk6UqAzDFxWOMBe/gZ53T7jxJyUGWvbc9g0AyBt6XLg6tyq2XrMq21X/jD
QmGiERWG4KeMvLbyP2hsWQs/2KxYLJtL4we95c2O8874itP/GOJtIz/fFrTMPVOr
ls9ff/rM4tWGdB1TzKVuFs+ZVuc7tGi6Qy61VZ3z/5Rqj2InHTTDltG/1FVMYIx9
cBtW0NWW0GgNfUcOaFogTNWIN1pRWxGQ2/2poghciQAUPzWxDywIr8XwfUgt81CG
2ydTD/MrmjJaOVnlWBWwTFkHCP+g/vYwmLkrsoCyMcH4y4Wglxm0yGtY2ImrDUrH
hAefPf8QmFB1Pc2srPDfztXkErUNcoSCjZE8fohiy/HU7hW5L2ptsj4ZtEP+2oo8
t7ng/DruSKqumBgDABqdDbh2BNXEjNOoZ5LFIb/JRenFj26AH+u5MvHQ3GISa7t1
a5WOqBxdlqxYQBuhJfP98OjLiX/gCC7DE7jKBuBvO+TICzTgWVIFwRVgpTaS5Yg1
vpVpwkqhmM/Io0rrOTxwDr+VidfcfM1Xd9lU2MJ0Q3GDYcVvl5KeHD7+LYeRe95k
n2vVLuDiYXb9Au0d6CZoT4TFGJfN8PfnMolsZM1dBNqVw82gBtFW27qWg5HFs8DM
YUjyIHZvHuNvTdgAx6HfW8suD+QvdkGHZgTuCU18ApdR+6usRpJezkNJ7ac3Rznf
core2SKqh63Z1r5ZEpCkGvty6VSw5lU6iPhlWPQn23WgqUKxAYqpGj59bwYc9LPS
KAzUqWTycSxgeX/ScfOLA2BA6cTYxGVIfUQcH01W/P/opfzErA0gi2EVyGel/Yhc
xW3BQmLgBBmSWTOdqIEyIecurxmh/8NGw7RyHazebe4Urrd5w87I22D0WJk90rc6
QvY47mzlKQ0q2AVDBj3wgFXx9fdZAKR7zlVXALqsa+imwkyyivZNCK3aYnys5Jbv
cYKMuKxLDIQXbkA68V6LgvzyqcGj5KiVsiTGJwVSMwP+0qkzarMygYSibCP09dfc
OXa8PoI4TJitQlVWSScbUBm3supHCCk8kgqba8Hh2tXGFBTJIlbjUh9zTMd0UGDv
gyyeVpnM/JEh8Z2T2GRHv+w8KLtpLRBkXjQ8aCCNsiaFLPTgT3F2dFMs7mTgZKtH
PtuOUVGQMcHbgrk83QAqqwO7B0gjzkxd4Mrl+ERV+IMS6cC5G8n2Z10exgcbT5xp
MqBg7eVq+fqQb1/eFKjoqzVtZosVo9S9DwB4Qw7/7d1+OvepubNIpTx9pdD4dELY
LJgBdRd1JuI7H6pflit9G0vMT2qpxkhwYZwouA3dOOcT18YrN/goieNHZ9ROFc+y
4SLpwQvp0hLxsHoWqQtaBi9QtHtWvmVxZ2mhUqZLcZn0wuV/5jjvZackV9smiDDy
ncQrACV3HD6OFsEEn5yODRzN25ahdQLEc1suW3DmIQ7/f7HueCkLXaaY60A3O+Ev
NIOAc8JT2IZ81csyIahCWl1pkOeHhoiLqdiY9EE5NbaZKCdNvZ0ajUAE9ySgI2kB
L540llgCm78nwdf4LahSCUAOyXR6Cb0zk9wjgriCrPjR2mjbWSOYAvSp8cIwkgal
gGMiwb+4J2sPJvgi6Uvm+ng+1Fg2KaDGYj5PhVu/M0Xg6Pil5c3mXDqs0/Y5HQwV
WC99BLX6ePOEPNY5bgU88Z5pUnY6ocKSKGkVLj303O7QJpmtYs+CKzCKrKGh6Dx1
v2dJ2RzTS35JDk760rYsKOUlnUY+j3lXmsM35lU4hcAG9YLGX9Y82aQ7SmXdBZFZ
g0JlTPyAF73unH8zIBen9aLWbaJaAnCUoZkpEmCBe30NUC7p5Rf6jp2EywXCUVuH
g7KtHeR1O7kiMvpyRtLDWrz7NBPbBZug58JY+AjEFjUPTpnDd8aatpbL7ZWaBKaM
gKr/DCk1TujQL78o5QFDCpwbitWnA8KDVM7rVdhhLS778BMXC1x8BBKaHaidW5QU
MoUjqlrDF0PQsXK9gwePpdKyId5YhLZCZ0LjYxBdbyQJBPt2M54jKY4IhaFxqxw/
oI2jjafz0LAj1rsVUMdgSDepuKrReVs1iB9xVpXPSEiACbZ7Thp1+JSBA/JHNyfz
rusOQlygM8qTVWkeBHUEU2yoOKqVBweUUsN1Ch8cAeHYAbMc3lNrB/1n6IW3/U8e
9PhKp1xGAUcFYwyduoeU/S7c8aYmX1jNCAkdbgO1QRl6ddRhLlHDQayTo6Z8FIgo
ul/e9BKhJeygL7gef9Wm6i+Hd+gNoXylCbrI/zL2vqqD+XkA3gaD6F/2P3FgrFuo
N5kAkpQqeo6Q6PBoOlIcH7JwQXtJukV6G+CbseqdcDEVvoe9p23C2TKjtDkzavLN
DElHvlRG6k7S6IP8rWu/j6Bv/LeJTDFiOPmRAymp8qZZBHW3Q6TGXBeDGfUniIos
yW8Yrp91p/33BMWMFmVvT9AiQIeiKMeIl9yf1Hvc+FuUy+jUiIi+0JL3ca3oBtJM
2bbtYbcp0+DCBO36WxcKKZ9lGLeJXjL5X/Za+z/egys1CHU3PBlT8cZMvpckM678
uOpYkeyvoLVdzu3DgZtSrjQ8JTAzq5yznNzFLcRUsdIQZhKzXkZkBVnkSmaDpgUZ
GpFCYjRdi5HztcZS+A3UC9jNJNLsWg4pp9fbtZ4jm3Y7MU1W//lvSYv724e7LBV7
mtmJ3mTW3wEJyT19VIRC9XGexH9srjxoi1y9kuR7tumcNPq6AH52Vtsx+DhJl/AS
nJl+mDEoXt5X5s/Mcl3E5fQ6ZhesHCQnev/e9srCzeVnjfzpj3erBUT1x8IQift0
Ae97VFokqQjVCozG77+39/2KXZzI8q9xxf0V+yNyg0lgRg4upO8t8g2L8FrpskoC
MN8OBh6d+x94ZIstNUjor4nESHRPZAT9gKfSergfgVepkoDmMk6nnS2uORf5BLO3
3Xi1582OtmaWrRJpJPh1U09t4hu0IioXh3D8VC2YFytVAG0XWyQvJMcYV3p2B2zi
dKAUEPCbHJB03VbrHATBivA37IGloqK9uh1GwH3ZXsxBAwTPaaiwOXDcY5TzIb1r
q8yQh12q7gzpM0+KIU9EIFx4TRiDJQYcy0QXAxj2kr9tCWct3RWwGKSQLqczdTI9
pA96yGcfCr1ys7YLfetPN5kJpAQCEkT+GyqRgIQ+MdTlpL8H6QvkJKUJiUXpzAT8
abRnDmv5CingqN0N/Fa9XRLQshiyp0NShivLnhBUPJDwzgmUuTmroErB0OyyD1Cf
z7qLNmB+2EXzpNmSxglaVdvFhkfp0Yc2NwlFHoRFtdMMg7GFTnPuKRa8B4oytU3Q
fJoRYfJ6fZFWjPqCNm8DBQSkIpXagcnmInhY2z5U9ulQLlYh5sdMIJe68QCyKx5P
xiZb+ZqOlq8Q/mTqBZvCUUAKrmwryTEIbhQF0jlkWGSmjvs16yMncmqlJ1W4QUK+
XCZrRXVJyL33lTZwQMKae3Cwzx5mFFbf8/ta+3Pnm3JNhH0I4BNdjjADNZv67C7n
FyU93TdfzupG/V+6Nq3sQadD+lD6ru/QKmXoFEjlaHmybM+d9RXC2HKm4JRe69yw
vS5zaLOhthShfanAWPe1D/4Cql3y8V/YrjXD55rMC45ugzVAM00KAjtW9vFTNR8N
uGfq2on8z74ggsrs0KVCufqsCxIBQQ0lVF3HYCdiXaml5TayU5r9yi/IXG8hUoL9
ofhTaJeiYs/sjNOT6DAXN1Zre2syTcrEfWeFPnvCAfwYnT03zjJsm589WgV36yyZ
NQQdOGSHKzz7JCbKmTglG/odDCNir23cDCyo1dj83ea7ypwSC+eDngmyLxQ8rA89
B4q26DVZOctLLluu4hc1iNKob3ud4gFxBOaXF+0336YkW6rcpUzTpXty/smrJmlb
+MvNPmwa4j/aUgUllkDKzPI4gwVJkrGCHoIK9eCxaIyXKjcQXgHEyiDJP0nmpWQL
HPT2+xjtqo+siBNaVsi8+fzeUqOq7uI77cqYvpns4GsxA9XdseT3o98u+ziAuq7o
Cc7DgOWkP5/pV0bBb3OkHetI95yprF6WkLH7vz9cquGNOCD1UpWlUwYk1XIoZmck
e117LdMsvFy/LnwaaJWxuK2OZuT+BzaSwPn8Nm9B+idyqj/TlYbm4/I3c8tjic0k
RkI9/T31BFZwZJiavSoAViZC/0o/+mo2spSL77jpZCnr7Ws75fdzrTlGLHvRxTRy
SXGtAS5Kb6Gwlj10lSw2Mw1vPxw49VRSc6luz90swbnd6dPTRZN1qagMYeJD5Y6V
3IjQ+EpKbwijpLWkFRKSMYLJtEgZRdMdAsALAuoxBuAs3wyoBbV1tP/j3C9t10i1
TbeUmuEwjjEbpTIkQFNaf89+Dre5xvB8UGdqh+ytc/6TyW5B4p19sIonxkgzfInK
bJ9l9/A55z/i1KL7QGdcN6IyIcqrtZFjvBtUfQCAMQq+UCuRLSJXBlHHvjbpsHE3
rBgHgnZL0s6ChdRGozUm6djR+OsHKqn+b2fuINsXbbnf64NRCTYAbWpm7otM6Pmd
spnhG8x/X7zN9GX2S+0VYCaS56m4CqBN17a+vjOBJy2SHok/Wr68urefd9oYLkXK
5InyLk4l3JQDp/gYTBJ/5+NL/DscUPwB1NdfTY0RHivWgYUFUeDzg2/9/ywplN+W
SCLvfwuWYG5CwZ2fmKdazr8V84oA3IUA3KbKIERTS99w48K6dAWqVkaDQwjMYdCq
gT0T+ORPLYOIBMHRfHn1S4RevrQJ0ryoz+Axr8a/uajuk4bLuPkZ6Lp8MqB/mdBJ
L8ZTmUOgdLw/IT1GQTGfef8AY0OFALXM+gEDBCtq2ZMc5Y1g1C0t/jUGTHWWCqLd
6GNVCMx6drWFYfu4yCIpRBO2/4ulE8/XxiUIPAzey5tgYd+ZmRf5eFKo6ZngnE9v
gf/1awSY9wWKG6N8syYNY5ga+wdNU0we9MEn8fQbUt0jaV62vSgsUZacdSKM+M/i
KBY3CiHOAPdTWLChdCdlmpzg2wlNVRkA5qcLrnEKKikUxn9k4PMUCdTuLJqWkGAa
JI8vdUIhJNTZtEtq/gCeYWdWzy6GgWvlZeJyNqCsZQcyyVRH0sHxbtiADrYNq/QW
hm57EEKyIPNA/OhaSnKs8eIu8hUnjXZBvNHGbA31lNvQWFG1S9Yc8pFgCCSsIVEx
4OAckfBb8HuLxqOmmP9gy1n8YVfYrQ4VnowIAZubDUySRg1N/Va1ME8OgigwlyHZ
c97eHhZ+CeC3Ren6eiYuaoH5MdgoKmvv0agD6lWFbvEKZiKIM80hPJ8SY16bdLTz
E/xgLShui3t5N+E2gs6pusVWCKe9wnV/6j5TE8ouXDJr9Cy8KPLAIioLZ2bh2Brc
qeNwMwgvsKTROFBiNpOIk38MdX1Ecsg3fjn7JjlmeWd2mECgyi0Ly2iCYs0YkEqn
+afTcsdnNkQO8zRW+39Ia6Vs99SnSe6S9kSEa7MFiJ3GtDt88LiAW9fp/gkdxK2A
S0O40ytZR54MYsurwA9zUNkskOD66GF5aebCpxydWnP7O+3JK4PtZ+D6w87Z6tH1
FQAHrkfbexk95G9E+A2wMzxgIUgdFl7azOELVyHG6UdZHu5Hb82FP3b1rAYdHJDt
OxaXqjuwLCf1X8sB12ZlQHQbQzAUgIUbTXV7Pv8fdwB4c6KoBtzFmJFXYoeORZ0e
AUYoJ0eCYcCawHTDAsEceEI/wjZm4RMM5cyoM+w5Wt53TcVE3Bu8riX70bMV8grK
T2OPx84PzOkFmGe5eOlv02txJbJrZx6NDTv6YFlzTJB3h3H8vt+6ltm0z76S8FZK
SPQQ3kOVeGzEy8MwPNQEryedtlcZBmRsyaidq7EhXj8muDGv2jXGoQGTVqB7Okes
fniHJKVfWM8W7byC/ORQhvhei7MMQtmbsjFWcETdYnw5rvukeNLhLzFUSsUuQ1Ss
meFOhdhOSZ6Bf3VTws7FoINjSTUbJXY7mX+d+gZzPQn1NFrcZHVzyd8QP7G3TxWU
+IvCySuuVFLXdVS8y534f+4Jyff/ouVwALKNUTnzwpLededB2ct1L32U5mZqaiAo
ik7YBFuGo8MsK20S8UZxu2q5FFNd1g1G1jcDXj6G5iB4Veb/iLYhSpMdcDS6ZDYc
hzxNXl6VOv8RoSzzLS/5IfHVtZ4YoW8BFgszuBUXt/mQmdgjYhkMAdzw8j90aUSJ
gCWN7WU5ZMHIbH5yBCgDhPe0Z5RvvxafbiYxZilwJNH/e2zRjN1hStZAMgDTBi8b
VSSPIcNlLiP6EwIlDUAbDlctFycNwW8aZWmMTMMx2NC1gx9ieNMMM4Y/jd5bWl9d
hVGW460X5WVmtw/lAiQJfGTs4NdI2m0nvS4D7WWTm7+Qao9LLpCwwW0tiz8mUciO
i+gbnToUY2EAKEqyh9y7F4oCkgLV9GVZO4AqwtugBcvgxipj3jtEgu5UUfr3QfJs
/Ijq4VZkHZ11/dazVHaYvpo+MU8IigAMUs4J/G5O9f2SR1b6As1r+DfkSCmgXHe3
7sBU23NgtSGffrl6R4+AEbIGAqpSQ3oWiJWbBXgn0HyyNZHaTPwdpF67+WKe0bbt
B0DYRqRb00vOTbUJA4N0vvcK4s/OJ8cOa8xuxd6N6zj2FbtDFI0UULeI+nHcu0Pi
jbqNnFCvL7t4NNZcI3ed5E7jxG1/GPEUf2sJn5zkp2AWBmGjds1dXmH+ut9YMDrk
Ws/5VTVFxgvxTm8QrjxTSK7ZMf3syBxVpJQxHiuxgFHXNx+GTVIYWHFuB/io5o+i
20tAvX8/uK/CBVNd1QWYQDG//yiMa346lsGMtCmamklxprbaCw4ONrX313K188mX
NcSzK4Iy5sLJRPh3fn4HxmaF8rOrr8dUauzFJBNZvvSmgJ1du2usnxI08h7GdA9m
2bI6flQ+kiH2u6e7mgYrAbLtohbIVORK7PUTGSdFwnYU/gea3N9Fc1PZ7fyxNBIN
UkdVx1w60nCLzJKFaxdO2KIOdSWYhV8cJQsxIBes3+ZsdMcZSiaCcXSS5WeOR1KP
OVTFKOq4ZxLeAmW/cOLgb0aA6ppjKPWTOIp/fwCJxHruTw1CnWSua4Oabmp2tksH
U53ZOfrW6QsIARRt8pXikdoZ2WFy3ayAZqZhTsNYNs+P17OkA244nHxWxUVF2WO+
LNmX7W0Qy4tz8AmsXR9ylwU54iijnvigGdvrC8I95Q4H/oHwNtTC4Xy1OCHNMCER
ztEPio4G0byPc1VrkdDW0zQicbb6h3ahUoiI41nIVnU8I4+oirM7HeeSGmxsdDMo
oPv7566acBmEmjPl3/G7Yi57oyuyih7iDJVxcdAcfDHsGRlS3WHiYx1bCT9qtEPS
TcgUQSMSlqeaiDPYirWO1T1FSbWgHZ2OHbXt4LPwuVNPbUiPLHHilfIh7b8eYqLD
/JRWVFVThE4qK1DGiKJ8OlI91caeQKL1iD95w4HaVVGKMJdBme5ZY3OQuJj9q7Eq
aGmIShZ3FK3OsVTHiEPH38gqUvF9Am+CfP+5V6sdw+y4jVo0b4JzJA/QplxhjW29
7zzRdMtfGBHdnjdc4N4a4beJIYUqPWecjYULqTN3MDk7rvsFcu/RijhIiJ8NNEwY
pGr5nbEsC8nQB/p7hV/j+yH/cY5cNkEO7D7CKSNzy5wtYBKlWaES3SCXGnTqGg2B
8pnCVftQp+fGbdjoVcleOM8Zm/6TjRchwLr5BCG4RpaavYtrP7VhK75ZEWhTAKbm
3ynD6tgYhCsbeqsZklLJvHbcA8gi3+/lb0YTpu4i7bUsH2gl2mYTQGnzWHnTwR0p
LAFkcn9GnnPr69T5bo/TcO/SoQYD1/tEpo22O5zIavQA6WHVzAGzFbRULE2ewG+x
vFuFxiRpNWRRWgxuwMtqW4S3W7r7P+lXdyeIJ5htegB2ddlJ8rbXNHml/Hdq1cR2
KBKOdKGm/qxHDxuLVi9IpfGIzHa+3MLDsGYrvISCuasPF7xpuBDEFR03vM2GKpFt
8siCoyX8BB1d8eC9+aVc0Z2gvSnJcWZ/kQEkjIOkefshX+ADz5G46j5fG3RplHkA
2W8UcDxAIzgqwhaM5LvSKB3/6/PJxstziFVOtV4XYeJrpzxgP8yKabBedYlbhcgY
gY77jXIJ6EzWRJS+R78wKaUXq2OgQxJ/efo7mX47RMYqXBPEgT5HxBQNAGUfqMB5
dkbxLdba2f0TixCrBexl/EeB4+QZixtN8IGqJVn9AlU/gR6eMpcXT/n3U3F1RqLO
UzlhmJjDwi6z7q2Lx/+hVBqZFUD29j7RgyT26vRY5axv5vVlDp9LA/nVv3EK9UiW
4WY+eneu7OX8PoEQVfSRBsj8VmTyscyBCEOTZWcILT1vOGUUuhlhO4fb4Xe5A1KB
4rntj5F2vKNMdFRgpKbO7pfN4sM+WdlFITxr2qLJ7A/DlfzrPvtXERj3g/n18nnG
M5ep0bkQKrvEPM5KslxWlLpKY6bgPaonOMru9dBq7F94yr/uOlbeLlB/ovwEGnqn
OMMI3fMHMJzY/HViFRkFp/XuHoVuof/YygEn1McfFPUX2bqPElO5UpGv+pNvfL/H
+uLE04oynwO1mQXlqn5LLNBv1bAaeVjhJbax7AxTbHNFs6n+5UU0HzwtLJ3LhMaE
sKqgLqQwa3MW6AwWqLUohMUY/t6vYSIhbTRM7x7fLVKcDRR9CFv/ZeAgAMyUZxQ6
w3z6h7/8muPjq4xe+U5XQst4vujiAuQ8OKmIAmgTD8adVpiW3skTuqcUfedoXxBN
nvtFRd8XOUE6rB8ODO6zdXe+N/rGOBgnQK6Pc2yusDbH1jYstPJU+CqSHszHPMJ/
QhUEoUk86rF5hU16ZKIJL1a/+eN2q94wT95XHamWTZr0sPFLfUBlnGjKPrpDQR+R
3mrKtPo4iapjDwHvEKUkW+faxR9LUIsntEkGrDEvkD5plrSYLGt4AXmLsHetWG47
TG44Y71B0Di74CmeB5KCrbokqYYAEqEBxpVL0wV8mWfZUzM7z5fZ1nsOKCFBcod0
SqXBusUD5AoBtwbGDALBB4Sy5JPV/uamXgw+fFYPsSwYOiofUubJNl0iPDMJUJLF
cyDQ1ohuegh7BETkkANrO3iYQ2rKVL+vjlFeUE6IHUqtPhbMnDKmjvxzuv/awn1x
5XkexWqNJZphyY2ZvB3S0OJlWypodC16c2gzi2/jRNzZmPLO7Taa97Ye0odbcW+W
+zhD+eb3sSjN+TjmbRFTkhxe2RQ4tTn6KuoHZlKDPptMM87VtmCk4wKDGBtM2uW0
Bukg0A0WcNza1CKq1ctT5IKBD8rrG70adDFVu4PC0WKWnbQ1Q364/gc/e6fCIhI4
zppk+gJ+g9WsjxEFmCJWvgDnVkiV7V1vibPnKiGJvEa8GLzEJ1kub9IHLlRQ093C
sQXH8XV7ixQ772LxdWcsB6GTsiIv6EhTGoJf3P7SB+jgWn6rk+TibB7yID0V8+XN
4AI3058E4Op795PtFsiEKeRAN5t+YbzDSyGCkY5SedtW7IqaRaRWMrpVyWSzg1yb
lDZ5/5ElIQqRQY+svtWK97Ipz5FEKMU7jTcVXLcEnCxQA/cRZP7fk5VY4LlpRg84
Q1hBGPzFLsnlzftffcROG0oitGIlgf8ITwBVlfCH6gPfqMegLncYkyYMw2aFp1mS
O36442xl/Ld81m3Th+5gaBwq4wOp5hNY+oCqfmaXHLvmttbilrIrAgPaeF76WD/5
1uVjP5a49XF8l/1m8ZIA+7D70XZ1HhEqUKXgLRdIjdlfwN6SbQq5U2a1Y2ZQciEw
45ySn+WHBnuXlUdNuS7QHjsr1ynUwqP6MC92bOT7qIiXu0/7mkFG2thk2zifFWe1
eh6XBd535KxRHbqHQaUjGyzd33ZvgSTFx7WTQyW/xyqgkCl8wm/Jnaq0/Q74iT+5
Qk/1EWixxoPav6I+UywECi03NlU8CKgE6W9YNHnP6+VNdv/322mDFTx0GzCBcuOF
vE/2dDiqRht0Q+plMu0nUywnwt+kRgOH60JXSpnveSuK0S/oJip1Ay/6yT+7WNo9
9eTIgBpYs9wikkcVQ+oDRinEDTYNk23qeMn9pMBFE3XWWNAkYoM+xsq/yR9ex34h
jUIwHifXbpjdOgJc+GJf2hpP8Pa1T4sevdHE4JWjS0GjCyBY5p6R1kTpTEHOWPZC
HfnMvJp0Q4HW3KRntB5aZ+2qNdivhTNK5TETdFm4hoWBqJxd49kGbpPB3OBLMWoa
0UTSBfITEkeA91D/JIqnmjbHbn037ZRHrHFHsG9neltSmk6Y48+RFWcyMd8WV1We
5wrZq1hYbY5b4PpSU3n+nV6/iJnR8COsFuDGdVtzrN9IgcFC0ZoYuKPNsDBDFP8M
eHtVVG6TDfHd4UNShdm7JYuZAY0ug8kl7/CsAdXOZtFCHJLXqRFts00aWXqZK6ho
ifLnL0EkuY/p38Ch6pOhAxcpfPkJwxcEhtcdElC2LqPt4Fh/Qe2qdw3A9DXNnhqh
a9GVd+dOSpxlr/JB3yDUuqG7y9KY8pbypNX0cN5KTcMse872Uxl6Shx+UEkWE8UM
jIT+CO4vBG5wrdgj6YYTNnzWIkIzHGmbbWeRSSoNKXozEEJDYrKXOFNGPVbV78Bm
Ib26VwiM49mCIRNFJVpc5mt8elOmR60itEY9AxiT25P48FdTPq29z7FQkU3guloh
LwB5PgiYJIZzVIeWi2lvwoFjcmqNnVu/OPVhEskmoFR1lq61jXlYp9Ohh4ZF0fkA
SNW2/aGRnn4dF7vqsVpyZJIehZ5rkPaEXq3/BzyjCUz8ziy3BI+ocNPl/ZxdILvk
YW2fj9RVHoUZFH29PcPUbAICAvOl3oJdcPINS5oTWTae3AxCGbqHS8X/J3Ds0VjZ
ghOy87narvJop5j2cEsdBjso4VAQE9sghn7THWjWMDviFv3xLGnIw0Eaeblwkuf4
l9g3dF0Z1PxURXTVDBDCBi2C/62Zdmd6FyLl6pil0fHq5U/PvL1yhwSaLbhRsSwi
96m1DAXjodriFuNJrNZE1uF7sRG4CepUdctNG7XQKHITuWNIz4fAQeJ3enO3MKQA
sT+fSMRClxLdZ0Jna/U6uFxkgTjkDs9enYML1HB0NLBSmEwsXo8Nl1rSFNK1RQ+I
wP0akm/BCZpdVRMut5JfhbZ1JjLS8X4+la7FciDE9MBbR97ZBSRLspY3U2JB7tnx
4hHD/KmKLVjuOJoU1Wrg9mh7fwC8CWAVAxfR3wBAA/J0jVkIKrqIQaC5mFdg5HJH
tbAUt2BxjfFVNQI71N2vqdxAdS+6mXTf+aXcITOk5DCEIc2632rQA00J4CH7k2OK
GlTlFonnqhymTWwzxydfH+XteuVQrJVETutCpn53ZpaBhxZJGKBeKQCJ7YttuQzu
4HWRdm8A9WZxIV4WXGnIG7nmRATMukmgjLHno2zX0L8K75+9wtnyUnNxvJPL/Ikl
JQivbRzhfq7lnBsgFrZsC1GxkqZeNe+dM6W/QtMCWSKhWfJy3zMeMzo9fc44RfiQ
WRJnq3ewWsccJ/Ba3SoVk9ZVLDIMIOeEbpa9sdH0GYJxZpgzTPSOk55JxwXugzta
Uvuf4yTFjNo00mM3FQ5+DlbeVUU5+u7ctB0w4luJDXfUmjQlrIGcVlHg9znjNqnu
fv8gvEDotMSxJW2lFXUCRlilEiY83FILesjo464udBFTxL/0imZL9wvWv5VNRulA
sDiWlbFVZAmFtyIsgbJKZaPwotA3yDqzZqF5+mhj2rWx7lfpGN0csFYJYvmXcruA
WOjYCgMCTjieWYXKz+/PFESB1B8pkZF7Q63m30hSK0ifYsFIZAMWTctJ3Idc0MR8
koBoz0zMvMq3lQTeG8F5NL2guZycGuMkl4xM2O2SAwQx2RqG53tOyP/okSlCUyGq
5dqvEvpqcZGavLy6g4l5oeh9nnx7lyHFRHrYmCdcLESomJxFys1H68t2fsECiglI
rL0Cjt3tR1Upz62ZoGdfQ59Rre6IpJXllfEtKiLiMM0DKJoqSvjt4h10lOuvF9Nk
FOj3eGdvD+H7Zl/VY+rPwDwyc2fO7QxjrnGRerSB0RXhkWQRq48VjDQhOOsgzH0w
sOY5iq/E4UTsfV2GpHDM8fxHoLOlZCsfpVV0Dk8REK2IyTPONXwGNPupJ/XveP6R
MLV+LvwpqXwxD5EiSHNhK021QO3MC7bhpMKKMeaPiYd7eyFFeS9CpHp3ByY/gggv
hd2URjcQbMEXcAGic1VKYpT/bJPuvjzpDchWu21xmeM=
`protect END_PROTECTED
