`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M96VUOdqpuXc+A7q/i8966VShwlnWPsUQjTYvYhuXHi+TTG4mpQ0egs0Ligukh9h
AnYeWJuzNUsUFB1Vwvwwt2xaufxq9ViIk8Rzyy0flQ20LyVsWHRxXbg0fbUplSZv
oFA3rIqtffhdJelluGwNkbmJbqebPOw+DCn3kvxaYZtcjvtZi0zx1/pDp3BUBQ9o
FffkZ+DVdWjl8wtPdCdB4iqOoEoMdYIIm9rY6buRHQBITim0gKwwSiHU1CeKZvLD
bc6Gp0fBPKFIHAniHBITbsWhmGklNzu78F75j8Ik9psZy/BmO2gHZMl81yqwCoe8
tiSqL9jWSVb32S2agC9Lab8d6BX4vdV+rvMC9ypY3eSeM7QTh/CLchykb55F/Daa
0Yh9CxV2iT9SWY+BkYHHOvGqscBxDyAAyTZbsAQxqEEP+fZifnVTcf5ljMvjcdu+
9W4F8kUe6Yy6d0qp/TftDgSltmLI6Bggs2LTgIAlSX8=
`protect END_PROTECTED
