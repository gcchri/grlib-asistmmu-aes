`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hv+J9MqiOc75HFnTkiNFFvECnZyWWhxbBFUtt44giuaEpBZU6fW9kZe+dksqVorq
w+H6tP1HR6rW+sWDeEWttjkamAlXeUGHeqfdt+jpn1w+ph6iYyFfjzRqvBWovUYZ
8bPN0+XKvVaM1Mfh2ttHzuZCgOlOrHvypq9oG936i2SIzV/TpwUeSu0yTBHmMNjq
gze17CEcJXK83IFG3IKi0P5d6YYhr0bu1yeUHLAWSWJrHpXCSXSJehE7qbAK8YEM
qG2+wZWAijqG71WPHJVVA4aAjBnBxk280yt47vjAtQoRV6SMgssbQbR6i1R3Fdsq
efpjB8e1hm4cC4+hMuHrXXPZAR3ItTAOJgvIIIlJ8SMoNqJXjb2aAyR2EpvsIvlP
G1wWzMdxQ0Uo7cuXeJC5FZgkzviJYK/zSkczHcnOT+Q80/uL/KkHsXOG50qpOekB
rgb2cCQQbxKP1ikfAHsvyeds8qI7JJNtRTeA6nIzynaWaRmjZB8Tnv70CiKMUJBL
`protect END_PROTECTED
