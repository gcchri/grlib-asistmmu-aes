`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4GIMai3WgvD9Edhv7kxc4E6JKcAXhyMZerbaTwKvXDOmfHSq09vlIJaRx+38J0b7
MT65VjigS9ctyqjxxJbyOBkJQTtZSd84jYs/48ShKUVbF2Lnlb0RVicJRK+pmNDy
3+QV/FQ/mSsIRmXI3k/Pa0KqqvMm1rqmb0u9NIDfedyf+M5g32vBl02trz2qHZhs
/9cgM+Cnc630iFGIefWfuDIg21c2FQxaxA1SZ4POeZfr2dnlsj1YwDpdpoGoX7/l
dAADWPHLKduzR4V7i55+aCy9j853+oFVfGvLB6is1RbW2HEB5j7QUJJnbetG33mh
yoYd0EbKj1bA4obBKnkwsMzzQ1o8rL1F59ISB86wMgIH+nXMcbLgERPD+poNT2gV
tzK0vGAMslSnFADdtuHirF8JAsZzjbElHnqH5KCCTC9AzB9dvNoBp/jUCWj9ZvKE
rIQn4TnwClZtnkNNeF09Iru1SxUGPPhlsUhFJhbO2cFbzTXw+BSy+cMrTS4gddHO
GnGrsXzd85JParD5juQWH+YhosszRBw4LS3LmXxD2yQrcX9CUOwV3m+KQZqIYbed
rYSvieNQfucpPiU7d8uTd5d4UpkBw+7xUawM9nRMxvAmu3sl+2SqyTKQ2WaIE9qH
wfyZZLgt1Wg2/Gte3DxqtOqXwAp5pkR/vLVvxWlyMPLMK8jLAZX0ToYIOWNnP1KD
oFAOgj9pQKah3HkSlUgCdmR9yyCIQdvo258t6QhcfEMVXhyBJFLLvLB8AaRTsE3Y
m8fjRHM5wymM/xuN+CDFTihPR9U7orQJQFeCWbQHhObQS8KgqZ9s6gxf8SjJPWxG
VSrgkU1uR4hhe5XhvGztWg3j6LV1wumZJjDDyrKWjeKFEnAAt+14RyRrkkCeSy73
SkrwjyXYn/nDPmVU2/Qbyt7bFbYknTj0t/Bixy+vcIDCl3U0kGXfelCg3B12GbvC
V0oVO0Vcr4XbXXUff7th/g==
`protect END_PROTECTED
