`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
intoD3wS8cGCPu7UtZEGz6tY4UFgOpzla8BmdIUkKc9smnL7eWUFIkaOqAorwngj
aW+X2I2w4rptcIgil6FUiVVKwfCjUEWJOazp8Xi7gJi0UjPhRb/wFY3/iR+PCgMs
MrA+1vrWmVzAZ6SUEgwpmUNR/QlpeIe5VS+p+/9x1QVAumPN8nP6HHkJzkhWq0W2
OdXNVPg90bjz0SvbOFWcPLuEagLBDNgVpNzYIoKAieaLNo/S0ZJGYctJ8OAl1DqC
Yw1+xCWhc0TclpuGJfJG1+4ogLQVh955TT2aHwtJ2E6zlrfWs1GDa6B2pRpFUmSb
7OKxHo9OwU7u1RlxBb7NM3ECq86T7tuVD9T9UjZfVgcdLahfZaFp/MHM6JF3bE9K
QnpAXDytpnCMAw4sJyFmSPtRsg5tH/KX5Fzsw8fbBGB1lOqPf7HH4iCzW47jijuq
Iq/3LYIIUAlz2PNL+OJb61TyqLVwMH5I/MTiMA7wKZY=
`protect END_PROTECTED
