`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OPQuyrIoXelkieaf1Rxjm5Mik2xTHNSKK0OY2aDH+YcJmMw5eoLHYa0xF3SiAa7y
MR9cqtsb1vlztOpsJGMiXPZY4YzuViGKi2fBvchj1ZsXN/DUHVq+vuzYL1o4hUNj
hVyc4vSwwllW0zPl7+YQH1CNREn+cu1Nb/4S/LD93xuAwZUV7KNuoK1h0xXRb6af
giccsnRtvfOA9H4xpfWaUG2xMtmF3+4IrlSdKruSeJTpljJivkLl/9K10lQDP3P0
9E/xEOzFgPIACHMnVSp0UkY/0OJd7e+OcglWGGKsgdZvQb1pWVTFV5Np1wkH3YqY
ypesVrFBWisBiP4QHtk53lJ1+ICh7AK8oDxITuaFFFAIeKRNCYvFnLl2fTp1el4Y
4ts4Zl5If4iBVVFDDxcH4kU0nvs9hcAqt/SL+U2wRlufHyYBiE+qYFd7VEye/LtR
vNm8gtMJtNlNtZECHPcyFgO/9FmQa+Zhmq2fqp/UKplklqh1qugfrIgjFdNBuAuU
bpgimnf5XxV8a8eyrnb00x/J9Khv024EcxxVGvf5oikTea96LcSELhThJSMQmLmj
N5RehbI8QoLT6gxGipFrbM8JUK2liAAmiu4pzhES29Y7KWWC3PbgQvHsJmQQDO/l
Blwil2afEh6kM4LBrBUHXAusxH4QTU2hh2g/KQp6JxivJfHCZkM3nvurBB7SkjM4
gxjk1GapwSTxioRzBJXRScTyAYDL7Bw9f/7EbEKOn/SUFurc+WtDvs2GGOznroAe
w+Uo1YKkSAHfVtuYaea6wX8DOvg3ZSXDCSDLCr4FDTPXEZlAA1aHiZ5OxaNdqGxP
80cCc0lvxSv7LUGA6JPdLUDVwn6DKfCE9thFRw+zJwoOcP3xOZ8gv1Xix5etFy1F
igY1Jy5RaoHvt6MFR73LYmua0IZjgCCWuCb0BPOWxIJRlPF/nFXyksqzdT5GefD7
9sFWHRc+9W4Dvy3eHPVtAfABHsJQzzgIDLdMfOPfq8cVeCFk7bdXBtclo0xk3fhc
zBgdCRVrc0HDr2oXgL05evhhAo/+oi2uPBeV+RH77cUup1xb/yRmR5fSsmaPdBj7
LTdPwPWRSFH5qWm7rAKPBFmMOB0Bmv85QjV3uLJLcn6cALayCIkZIgHdAcdSJLwc
`protect END_PROTECTED
