`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+LPDwbgzL1o+DWry8gYQmLyHuxlOFURLHQbpbP7aPIbgMLOO707k7YyM/yMelZNY
RJQbH1KEq0uijudTPSOxnqR2ka0l4EmsGBf5PVZK4lMkqa1VHjSIAB1UScJfKtgn
Whm9p7dGXCl01GE27F8agBuww/4NYEESI7+hmd6A5XnQ67ljVjnIQkHayUcZ4HL3
FTFic+bNa9RRfzno9+iulstfE1hnqpFZkHHIJV4QJGIxBXYL4CEkH53osjJ2JfgO
qEDtqDkuTFGgBOUgSD9wBIUW3Zbw+4TrpJCKpE1Olo4C6EP0MjDa8x9AvbTfuhcz
dtiWOSwTDZD2t7gL74TLxA==
`protect END_PROTECTED
