`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QYb0UKbkzvKCYyoYyQh3u+/LJvb2aGeqEaK3XHuHhHiIGEupujkIosXWTRwTnohB
9o9NHIHMBB42foSgE16MMv/L1Kt1h69/K/H67JNFbGElh6tXIGDsgdVCPec4BweO
7PMDXQR5zwnPJIWlBnNlI/3Nuq85itUnBrTUZio54I8b/IbIR3NQRuWF5nmMUOl0
OAXljgEvLaEaeySFvRljRjrjGr7CWaoJRAVykxWgOBFe6MOgs+PlCRjCpAmZ/Srq
fm3hMCL6WbWbrF68QwLtv7O9Ty4jYfkOWoNyZQhpFOJdJNFCQGbuTIf0zwKcthmw
NShPMIxPDmDBZqyYVpmIZjUsfiIMRMVGN/PxzqyZCglIm+SEdY1kCi+dHJs/STAe
cZTo2fcjD5+q0wwA8OLolawZRB732422iDXP7pgErztfJ86HG2VjwcJBNsxeJT7d
QtZ2Q7hXFQRUQoWAbEIBXWB7giiUgp2qYLG5RdC8pVuycSxZ0xb0bVF+9kh774Sj
FecMUGC6nEBtEJWakZoqhBbakNBlp71g/yuDKWP/Tk6xVIsEWHJ5jl7gFpRN/ruD
PvSbKJrBjxutygkgVNTQeJP3KSmh5tuK8OnoRzSrw28BUudqLrzPijZBt1wS9eVk
i+/Q5xeHmGXv0yrVJ1Qz152bcjRlRkF+hnS58MKkWEuPUPMp//blfljG9rFueGka
Ck0+sbQAxY7OiQG5HpJP+ro3pLKmohZK7y1WBp+8hf3YFrJZzbDRLu0mneZqHWeR
v/M8AikZinLUJ4fxuZqWdTGo62tFkYcRFRJc1afzZr1Cqgvnd0As3+Ni2lg4rFy8
lkCdqQ/kgmX/Nc/i7lasRlA8uuMNQCBq1MB5PwyFLU09fsL1FCZ6MdzsQOhUfgMi
P70fdYcwy8pgk81nBobQHCB8PWNFiYH8YkxUqs4g9A38ERT4tE8SjD0Nq8wCHWzC
9NKF/DruxD4UlZmcY+tKXnVbf3e/5NwwMm7I6oXK4q5X0y8fue8AgiOeSz74e1SF
rhgDFx544SKKYiHDbrR3/DTTQ8faotobyRDfxZUQ+nLIGERN61yK3SMfDydLlYrX
tm80WNEhT4MpicsmQNbMeIZiD0q09WuYlBK6XcPmnbQYGtuv0zUwc0Exrr0kHsF2
ExGPRF8c+K15bU4GGlSAZkPqkh9MQjpJ8BEouhLiGY1MujEvl/sIBYSxpr2Y0tId
PLiYmErgy4OhJRzEErBddzYuUtTcUJPkTdtj5htksdJ7JdKSmskuHNA2/cM8tgbO
EMXri5UuKjAL2qTU6JEAbEY9wDywGxmFwEYhJX2rwyfbZ4PzcR6sTYHxx3LA5h6S
6NS1wHDVLW2RvL4kjsyRE+VMctDfuJf8PAfR9TawqT9TbjhRGBBKV4hPkjdBTQbQ
ggWPP9AgdlwEEPjwlwja9e6UicbngTKF15h2OTkVO96bDVJ1sTyC2Ki2MHp3Gbyv
UK6xrp418wxBakYF3kw5p2ecNODwyIKlYOZyaW4Z0zY84tNGQfKntOjomRHBGfFe
hJy0ftniYKPftAQlhrBXQ31Gs2W7AAtvrHtiArgutk/qtBer8EFwl1wIdXcbyJ+x
wjQFeUcg9PgFd1+bfdyNzCPMbHmkjowQYiLttXTDFIFEvaKg1Uv97Yfec0P4ihT2
YKYXsaZ/E77qsSAvFnWUqgGXZpAu4HRwlnRUeL2GU+z0hY/8NVUFTrNSlNYxQI1T
+7VioguuGCj0nXiJkW+Eg6xMTaKVSrUeeHfAotlXN0oFhT9oa7QSterKrmJPnnQe
4e7Ye8HxViszDk0laKTLjIsQi/SRblngfGlKVc30qcZwHKI+ttLmWVMPuVR0xNZa
mZTLWMYgpGGtbJq1/apArGCmDTwd2pvRP/ohF63lLJpyKzPZsARp34suyGz/KKO5
xdq9cc+XiGjf+rWM2uZCwsV1Z5FHuvlyU4vIUbOngkY=
`protect END_PROTECTED
