`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GvgttGUr2ZSpZw+zAaTRSTut1iC5FrE+os8oRLC9rb49ol4ZZhktN0Czh0+pEOeK
+Blg3CRB5NJV4oRqajWzvuoMavL4oxw2x3QE5Wx208AsA5nfDnZDHtiRUK3gItMY
agP5VqjuvS14449qzyqgWKGW5yL1waprO44bL+lPrmwLRc9r5DvP2lDkrhE7MmQQ
FpePp8rheFd8kca9gLipKH0P+IKhi/9nRwLKxTqddY7eZV/Nrz9gSk9Yx/wn4+RA
HUzLBqZiBWM0/QKQZmHlVrMVoOoWuOKfrtQUjknzxjISXesGsLI8gm1ahSBKxGDR
EtLP5eaKYlKsXNHQMNsIXeklgWGbienrKedxBn55tbE=
`protect END_PROTECTED
