`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FgR9H4ap4BvDFBq+eftzgN7khku9kNih1nvEEjVt5OeNbeCb9ADZOcAyL8dW8I/J
SGPS6SCdrGaSbDo9+C1BQ8DnZZ6T2XK4KU+HprImJBxEMju0/9NEbLLk2lbMaBPx
OaOSg2LhMdTBA5V2NmdRLJTQvy0qwZKusJ8rXqJDyaAUkygnMY8R+i+5NBgebvzk
K+IixcRZtm6YcnLwjJ5GVAtH2ZqJvyWppPC1e6BlQxvd7e/bOWP792X00wFB/Oex
BFgdv7G/ei0AHIgWlXDnM83veED0tuaGCcUM+2EKi2qIizrQPwHIAOnm8fqsZJi9
W9Zdu7kb9k7aiBkK0cvFdspnXYWwX4keTFt1i//9QkB+sO7pjH5IscHLnSlGFbqd
JhhqlmHpG1BtU2GymCxnSdFEtoQyxTA04beeJdI4d+peuhvGZiIkjZ8xIkiZYDy7
6J1a54tAcFJWV4OihWXGKn6lowuYpjYrT7Ad8KsKgBe7mQVMmbSSCrzhWvMHLa5A
`protect END_PROTECTED
