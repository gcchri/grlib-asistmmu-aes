`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ROwVI/WjkFi5poGZGU1wS45zNwye8v9DX0Gko9PQTHmf/9ZZq3l5/YCKZDG+wXIF
LLOnaSln+55gb6DWRn2q2cS96lw1Qo9uKRk4254/Z46YxX2Suvx65qVH+2YaBLDy
eciZwWW+V6wOYUHfw8UNeSjHq53+L9IdO5PTS8bAZn4Mm4mdNAchNsKPsl7sPI8K
Dz7WylZoS5U8H0q6UA/ByNx0vqigJ0veSYULj+o7wNuEa5esAVuF+2JHtozpP59W
/16BXLvlmkzRF/0A6vm6k8eBrvQvLQHdBLhVnLKALa8=
`protect END_PROTECTED
