`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TRqiqCdUyp7s7hSZw2JxovoSNPzU1GAEhXpPt2RfnDUjNzCorBX3ZlZh7jidLddB
8QzGf8oyqtlYBKmYf0CXwRZxXz15O6/j8DC9XOfpRym9ijSgeiCcEsjmrNdX4jhm
TWyIo/IMXI3dDcE+DLcw/1ISszz/c5DdVCOlaWCeR6uPaFX1p2O016h/mWRqItwk
fK4QIFn14fqbIg2bQFMhzPiNwsU2wsxgjlapeTJYZTA4jyYWR3wsBWj+XIrT66xg
rTJ8hXG8X2ygAVf8CwEZscVllFrXmUXIJ3d/EkXc5iz8VUCLg9rm984dhp5jx4jF
FFAXd8E+2vFmpl7XC2F8y3WudzxPZrmbYNNsDypFgSuI51kSU48dKycQWD3JQjvW
OQOw9IdgFY/fsf4RxV2XLVx2XPZxcDVOqFQwrMg5s/fglc+tHbR932DCIHFm9ZQ0
3ntGy5ORDK3gqrBr6M94Jn+p86kRiLYTVhWkUywVGgZiG0ZXLzuoYhtwDMrItJsz
qI/qS4omh1sNwFC0lssxYH+0JWkO3AUdVPI6mLPKZ27iRI1YrRZRBymLOyWwABnt
g+FnTwYcGPET3mYSDKFHRWcre9zcrFcnjioYgO4hPccFfczySnN9t5feG0PeJVIa
Mx0X9PPQa4OR2szr7GKMOYidI70UzIalMVQlTP+GlLhpA8cNEJL7qQxFhVJqoWHp
+eZyDE72UVfui5tmxeoMvcGJXRIS+MiX0dNhZh0Ep+IAZs/bC0b6A1wiC0gBf9gP
8rfoQXf/1Ks/PQJp6dg6oqriljjPFzX+lQQwxByKTPwixw0cv6VYjlIZkUqiI1XH
wFAB8tJJ9ma2kKNI3L5jeg==
`protect END_PROTECTED
