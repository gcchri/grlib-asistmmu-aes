`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QBJSiy1yKd1o6sXCIX9Yx7G9TYxIqxlG399mY1yZgi7fBRzXK6sGt03rpnbeC2Nd
BoXvR6TI+VhWYUd7pipoIS27sEawmUyn4K8qWFyQsZamEsYy/5TLe3+MoBrfKCx2
8lw8Q/3Jc1An2llD2kjwYONwgzvD/zTOXdLUa225a+zrx7Psg30MnKP3oUKpNeJJ
t5c/OjlMKg0bDAEpb8VpPKV9rn6tWuA0MU0/cZ9BMGdMKEgLqZssUULl+xKslQIi
UKaU9OXuSvRv378r3kVdTEaP8Z5vtxJ02AXR6QHOv7ViKTtArqJOcCSTqJvKGDj0
Ju2CKJzBQh8eC5BaPiLCU3jVgupCO0w+420q1X+f7EaZUwwVsOrKsZzbC+Z2ghNo
3ycPW89s/hQ96vBt/ag4C/DVEvbMI6E7O0/tr/VQgMA=
`protect END_PROTECTED
