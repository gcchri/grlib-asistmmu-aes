`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TBpop/q81SQW3UzxOOjHQosrzS2K44C3RXTO9uEb+RPEODlPfd21KC8oPij5TY+B
E29mnPeV10k8KKJQg+nLD7XexxNORnL6Alpe60QYJS2d2JHQC6xwNdwXA+yAMhj1
1P8oQ32Tbz+jvGbbRyIszTzOjMA7WsY9Ovp0+eXeldFxy5zfKYiyMBGS0OvJrqdT
+KmBiZCt9wwJHG5EX2wRH1HgR7xKB4n0T7PqcU5C4Nap8Kn0LDesrkkZeOqe0ah0
gr7QkboMfo200oGeu/XhpB5s23iiyq/q2kw/YnaiL0KnG40gzXvdUsLKFbqMJE4D
RYF4AF5RQH0NFwNl3AFagQxRnfgaq5d0843CzTu5DyjXCx0Wcgtw8RThZ3Uv5P2Y
rvqTlRCMxi0RQhN2M+8HM8KNHFqA4rwlm9K1D2u7rwASDgcRCPbmh0TCpVlCWSjA
GyjFKXYJuLIqXahEGX50XbExtb7pR53MqNijS9bzLlu65Toi/Sb7WBREUiSP+7l6
M6YlwKlrnsIKeUzVayWFCCXnhF0SYEPd9DhbUHFdm9plooqQ1J2tryesQSkGXBbT
IsPinqNVRQETXyzMXcUuYjeNiRW/VqnvlGIq2bGAEcFIGoyKX0lv/tAOrvtUISG+
RtbuE9IEMqcxhRHBka3Ng5d/jvYHV95wZyNwKQqEzayyWrWByJi6XaGFOTSOqVSX
r6eSNNGHwDsoz4haN/i1Zm8ieYmzrkK4lZnop9EjbeltN0C7pQ3qttGlm9ySxHVl
6cW0bB/lmqWMGTy5BbZNeevDQcN5Y24J/csRAXAPXc8SyFdjf36S6IM8GQnBHf8Y
gcVkw7GZok9nflnBurBbXFusU7fxDgqyhz4zSL36bR9UV14SzV+KoUqU5ynqMoJx
tniB/fKOHmHtw+oSQiFuPnfMAIJb+qOh1Iy+uxuCBB5WQrmC3ZWjMKpkGHK+AIX2
TOYbAw0M4IwjfdtqZFV7s8NbNqOCQM4DfNNp4pDr7e4eqzykDdDutDuiIPditQSu
r9JUGUUtNo/CeN4HZbuscjpA54OJuxFTA2fQheaTyTnKNku7tIO+m9UkornvkUrT
P0yuo2shEQHy5RifDBx5yYU1+2sRUiTDSNGDK/LMhort2C6BWbv/Ci2k9RsVMXsv
ua5SCAORYCzi5gl2NZ8Xaoq35VRvUoHb4STafucsnNsnyJ3taMv2l4sNZ2I5gAzT
ydS7F2zzEhyXbF7inx3jWAe1Edgwa7B3C+klAw4+9Swm1m4lZ9oow+4bNFh5tnSe
+T//FsSl/pcWVoQOvqTAnN4+Okon44DeaJXy+jBJtTxZF43YXeltS7eAbAY0K4uW
H9QF6AId/VgLOiMyHH4UQyz4XIQZjXffSPU+u9wwV2RJ6J7+m5uTj+1T21Ajz3rN
yEwicHBwmfSESs6EBLaaImdnmSpAtKDXbNwEApKWbJak5N1EZ9KMxE3nsa8N2FWY
IuMlBUAmO+6wcZWACJXkZeuS7RfjYYBWj0SaDynMkOOeJiL1z5TB/63aWDSO4wuA
xaPgfgfArH/CBAFkzaJOML5nf+h71i3Mv1QDtzp+a8YXhRHYLRkjfgLCrit2Tjhz
heRDRx5tKND+FmmzWe2LDIwAKUaHbO+i+y5apT64vHYt2hJ5kfWlLr6DtQlo1Ja3
LGEhKjPSfzfiYTTiEUgfYHtvQMSoi4AVQJ5Sx6vNAHYQGwems9tYDlIXZDtOwUvo
RjK4krpQAW3FAbtiTDKLL7xsWop1T5jVmSM8lMtKvdg9ZLU8G1Jqv4dMU7dBePAw
r0gni0SrTdaqylET/gH7HNABhf/gZf6Bs7esAvjRTiPpL70YvU8gIwDMy13RsJi8
TJQcgBUgteNJFdcqxkBpC3ZpUhVPtZKL4kmy9L9+UwiYxxE3+xVujptGyreonTzf
ylfQrZp9fym/+n/ypksX3kbsHBGbyh0VRElui1zxoP28mW9zJLMxVk++aGEK2Jss
u0dlAghuxW9nlftgvnfRcjJ1bh0cLQLN0K/OXHGY9ZIr/9wFJRhdXglpIO4lku/L
/pgKZHLeIxwUcNjc6qrG9bzXzGn5sYdIfEiZ/Tqvu9UgRNhV1H+OIShP/3+pADSv
9c6maJfm23WVxurXo8tSKsKidOtO3+mOtQqqPve1xurh4JQiqJvrjg2o+3yOzMB8
eVRN563XXS7RYrTiBz8A47tOSF+bUldYc6lxPOSMx4WDeSKkT56KwPs9JQhVoBEM
EEqMc9OPXHLYHMr5aoW8PhK77yQBVKN5YBraqTv4eYI16tbrH43H2EnR5jiUOYlh
XQZMR/GTtVc6fglOhSnNkXJJ/g7ITZbtHrVVZ/3JQG0=
`protect END_PROTECTED
