`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m6HZd7Sj2LXcqwHqxdbrl2x76ySWmc0/R8MnUnept0zNV+iuwy/ugo2TXT82Us5q
DuE5ZMCG4vaau3oO+s4YrBYdIW+VnH9Lz1jMi2d2EEQDDy5z6wmayqoiIrPtF9pe
GGtp8fax74WPNvBc3whiydnOvQs+puqWhbwrEKWA3J8Moatqw7UXDafNOgeJGyMj
B6Kg0LazK6wVpgGJ7fF2B5KaZUhXN5HB43qk2fKObuELv6sGH6U1Hme8ki7aIsEA
5smPnsN0UdnqTaCS1sv1f0+KFcjcKP/cY3RbVzvD+Z3BOeZcBSYAoYiBGhmSF3Eh
lHwX7Xu3ljTf+a/9SQIsPNGPfiQM+LLhyyisa9nIQZguTjGyvjUjKqawYu0uNxVB
YWCB9PeX1Xn4W2uxkUv2Mg==
`protect END_PROTECTED
