`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rkqc1mAO9dZxgXi+vmuaoHY0U+zBC8YHR4q1ZV5Eegz3NGHpRelzNRA/uN64dg/J
G86dA13yYCw0QjWcMFMCzC2z/cn/Cw9nOJfQHOfGeyFw6qTyazjwdUfge7bpqZ8r
mfVEN9sOfdvhdWZmN86oxd7St59SCD7kNAz9pG2GDNoCDag9OF0sF7SgObrPWkQo
Ht2IwprvY8gBAgRZ09oxuoh5oZQuheMdMqctcc4U0/lPUVd/rC2VZixATaPB4Dha
gRsv27o23jJ6v3yg3NIjHjtmIRDf8EWM8ixTqXQzRfCnnudxMxiwq3erHyrkxYlK
jR7OihxZVlaZLuxxQCLO0wkftp2lDqcxTnGzfXbrBFuMuKpVHMw8ebZcDiU/Yhnz
ASBTmUWWbW4X4RqRspUH8WECpzKfBIvnENs0m/GwnqDA+1dge3r0U5pe/eXQed9o
lWHJQODX10tlfmPHA8kw/ddLYdlQXfx8S4aoIKATQa9R1EsKPEBJsTgTcHf6WpSR
X6vfsRHDzHXq/qKKpOKejPcoUeuDmRRb8ljmbpoG6XDxUAQ8ssLnc1GwOHgSfdfO
4JrQD8KSVpg7w1ZkJLBNHJl2mfO8TJCpexlM88NuJbBjJTv40Mi3z2fzCEAp/Lkk
+/QVGxYZ7+jyw0FKTqq7jGWj07DTviAPyWcD1poEKuSCIrCG4lyT1G5KrB4PQgQ+
PPpgSTJ72ti9bDiOuoj61BJs1NOKAMmMYQ3zHSclywwRKPsMjPZ/xzEumt68Q4uD
YtXjt3ZfeprYob2eWv0PJeiRLCK4Azty6y1Zn76mYJMiC3GLx7ctimlVYdUFwpBU
JXW/DEdkCTF6PYTijT9CGRhNg0tdOOsElqCqptTtyhztm/AY7efkXllejxiTr66g
FPAbPqg42ED5Ol9Pyp5uFcYnh9REM9H8XStx6QVGkZecWJnmKDg9i79kaEg5kPJI
2kRdr1SSH5o4SsQQX6daw4zK3kMADMJsPBX8e7dx7KONgmx5iWJtKOdeFJpBvh/C
O9l7u8h/jNbxXPN7Hdqlhy1AAmAc8pt9K+wcAcoivZnzt4VUu5DeiNNBrehpzlDf
U6oZLOxgNL9J1Ro19tz2JBMUpZunTVozBo4G3DL1ApC6LCmAei4S6GZhMVJdF4c0
epQeIPLqKYf/YV9Gj0DaSKltB4HNBPrutdENexLEmu5Rf6tcHZ0IP38b1ZtCyY5c
w0Abw4uTcUyhqOzXJJZWx/jNVdb/Zf+VkTQvBQVD551Tf4VJfx39v4RgP79UAvEO
ln8L6lb8RiTFZ1moEi+2sK/YV4F05coBCEBTZm+uhG60j0DYuMQfmUshGElDXOMo
heuLQ2F3YV+/a5trDRI2WylzfWqUVc1Fjz0Se0Jx+pHIAfM+vCNrx3/niMh1BLs+
CuA8OfslIWUze+A2H9H1DYBzFHedSW4LyPQiKiw8XovtCnHPclH2dOHbhPWq0Tbl
N+NdbBkPCuKXVX5ssxhC7W/kD6/LOQTyr9Zs4zz+a6mHi2986OVa+Smu8fbaLDb7
uL5FE9HdEcifRP2cjwyGH85Qc42cBBEa/M83kzZBGHhpeyRNMDRvGzV4LRh7/P80
rT8aZQcR0/EplbFrJjpvOqYV771kuhob2KZQP+MDvT2V73QtbOuFoYo+6kdOPD7d
UCFFomWWFAE/jXOiw57keXG/TT5OTgnra2dMNbhc0CmrvgdipId7XhHCv9fFfbVu
A6hupelKnWBhTXZandI1iHK/3BObkplX/34oImj1Z9roIn4UubY/gonsPZQHAtJG
CXYaOXY932fxd8NfC4dTsOamXuyHt1cjHk1MN50TgYW6VZHTgBuN5UTbxmBZexnJ
dS+MVuTebbyZvGJzT8zx31x4oMI2eKUUqGvyfkcRbX6ykrgh78etlpU29VYqwvZS
ngOEgv/ZapPWfx9mFhnYQvk2C14wSn83xz9pGrMhiIWQg8hzUG4Ve/igF7cwyFlG
f5D7Sl1te7xJlB4w7M7/N6l7UgzFZYGO8tQWwMxHJULDaqfkEY9+uM39FCmUeGiu
utcVV+b6GOBOMjzlqZAszNgbWon7NENuZhprar2oy2IpETMgCtgCR9uytxCjd9SI
zZQFr8DMxD3XoZ+MN+EAUyfgRXAS1YcHnKY8bcQ1IIaRX9GVScRE5QggixnAljJx
nmu3z+nVp2RjOyhTfq0bXAR7vfDBsada18Y2rxISKMyN3/ssFB1X8P47LkeW6J5f
0Jl2608ss9tjqvaqqA/uR/lGSPE9zioDLaIOm4MA8dQRjfaMuXccnPuU97sPP9vt
kKOiX6xCKChbVUMQ2KnSwdEYgkp9ueX/ZqqxGwZ53KMKlv8kpbcxKrbHNJneoFUY
soE2D2p1u811cczP7TVZLUH/jOPX633FMg97/zHuFvjdh+7ZKVZnKOk3ZS8Kw8g7
GLOPfi0xWuMWRCB1RqP99KRvSniIB3zI563QPGr1elM8uD1Jlcga3wlVtpdXYV/I
D7H2hkC0Z9Nvz+07lpqNEHAtvSVPovOuJiGBjJst0FFdXeo7IMofUFKiOLXhF6F+
lLxroiTQGTp/ARhyZfwtaDpLOd+IfNviUev/D+dj/Qj9AOtlwKlFxZDRY5qlftfK
Rg1isYe+qKsJZUA0fSjM/qqS9Z8TOyUDKNXgNpMDBiglCVRMOBW8q2XepYk5FkdN
bbuSvqirSN5uJsBEq6NzBVy5gT1TD6T0gboytLNqu1dyQxhblCthvjWr2vMI0nNA
TBoJHngdnmWO2+61GH/jGMbjBra5fI7JS/9rUEWuy/C0oyvWPT804UX6FyTEaMTV
4vmMzVMD5G2Bzcr+3pFFsxJ5ae676z4cOzI3K67j5jJqgqMlp6voKEKw1yfGbFGd
q8zas9HD9EMyhHdP3KXM56VtilptqPr8TNuGL8FsB3mA/V1grwELPzrCVqCP3Txn
CG8lOBMMXx02FrY6/wCdsaoo/7vOssu9F1K3+NDhRikvgPy2hH6Ny+dg3HTiUzgu
wvqdYI7yuj0vtiRcqisVR9ulzubC0htuclzCjzkzsXx+VKr8wgu0wWBCEYk2D+Rm
a+hanP2uJ1fmvXZbg5PiQleoFIs5HD0x4pNUHsnhwvk9mc0ySciq7Q27g3PWcHTm
Jf6NysL1Rx6acvYtvRxcAYvpyXWcVVSIjvvrTJubOIsUhlsuK2TNIo5d0VJpChIm
hgcPwBUr1lX1jXqmR6hOnprxzFhclmM4YypIsRTX0fM5AmMUV/bU9h5/3xvrMl4j
FrUmpoLsM6VgIHZSmEYIpwtAjSTMT7Q0ydwTAvLB8drggr1qi28rGneoBhsyzIqT
XfefEhbDnOqoRNSKWREy1MA2m35z0kGrFD0VyMcCrkOm1kKUfobEKUu/3EypcOvT
cE02Vb4k+FDI8MlPoHKZ+JwCCLCIcLMkInsdQ7+f8bDYEa5lSpAOJ/qTh6w+Xga/
UJkEtOCdloZ/Jcd4GOJumWSR0N/mrH3o7NOhhoB+6fb+TQnTbzenA9b9uIKwazMv
m3IWYV4+9wWxXdmhgQu3ALG5ZbihrJbHVrOq8xl2YP9ftWAHkFnC7w0A07a8zDeE
fZC9/5Nl/kWubSfWOIiglv8y0DW/kwU409ML/z+Qd9gtOrS8zJVEKj5Zy237vGfy
bRWj+FIbZTdjUmt7jTl5Ik1DkkoH2uVpfVyq5qUOcfE8M/hMVnfRo5K8ZXNGA3qx
a0d7j6sHzE0+Cp+fF6f6+1/3Vagpet9/dcq4igQNpRKNIdP6aTJbgyiOQ+dA+CuK
sni8IWocem+g3idHGReOaC+c7fnJxFR6cdkOfzKB+RUREg6oHvBkzYisPWfzprUR
3yzUU3nNg7R0g8+ZlYVCJhUEJJKJojBvo0itcIEII+1+FXA8gru1ZFMEJaHag5XZ
ME1QrQwH5UNdyCgWj30pnj4LFswchRrc76Cwh9AtKTagt53V2uDAhvlg8hCvi7ku
/0OC72dMzmvEfXPLDycoXVlYzKCDwWmxG34AB2Ihca1eLyn8UuK2PSN4+iqIIF+w
VmNq+/envsmUbphmU/sV7H9jmpcc9RAi2IyUsU+2N2h2jgTpxanc1klwFtiuVN7Y
ettQpEt3+2zBkAnlSPOvnvunpRzDZgfdtq8gv2e9VhMFYLOvY5XEoCpWx2oTLBJm
xplkR7Bh6NuOxY/vo4TFucp/pBGIMnDwhf7dNklLr96K7XD4UJJpuOubIoPVh7la
4BZXreP0kgXJrI52agN+Cvcr59Q3eQ6RoLtb7i7y2EewVCx+4yQQS/t0nuA87REB
scfDYT03YqGUtRmQYl6zBhOQET1W3bqvFAVSaLNMwPITF4iZcd6vWKyahI3LRAqt
rwJLIPHYdcI7N4lMqutjdOw4DJ35H010WVX3Ar430tEk62L0Qb0cvFV1IaR993hN
bQIgS/rdEZ5B1xAM2v9fyBH1GB7+i7Yz53rKWftmuy2fJZ0F60JVdTjwsV3cz+On
nrqozkF56fv5k94YrwKtRgBoSHLotK1kX4xQGKUWzw+v40R42VXpEl/8iaMc9ug5
HNrglRA2i0nzjattOzDj+R821K5Nbgiv6aLVeWpvPJZ1xRIND2T3FcTJjAaLJvqS
8ldjYigbr0xn0USc2NI0nZsjOQcweJ0gjYc0Y01N44k6kHKt2S6KIN/Nt+IhHtfq
jhRMe18ilF1P9aN0m+w0Zxy5m7eDEXrAREY83A+p5kMBVJryFOUdNawfnDvpWvSU
hEJA626TL2BiwTSUQTgjECBsHLxlzejxtWdCalKMKRL/NTYD7H/iRZQMqwPeWq1b
blLMqL0iAN+cSjsy8Ld7ldhYs5ErC+QIhzmiLG7XJQISd9qnVRgOREuRDWX5XTnk
d1Ewm3bCiS+Jjj52F13jMhpG3NxjizclNYp607F3mvuY/bZpsMDWTbact+pbfsD4
UKE0hSyp2qS+C9DXg2luK0LwsvhCAnwaQ8BUhDYzEjq7yei7tzw7fK6y9UGhytQ0
ds6N9JHgfK2dU8MRBHB+hYpk88rhtf4Sr+u0pjLdo1Gt+ksCeHrJqY/X9MT9cNpf
spsE6zKH2i1CmpZ45ErDtSC/xy8dXKgBt2Ku+vGrXG5yARTB68tQBdNzbvvuUeCw
3sM1eoMFPFuyTGHMmw6gcOyEAyW/Qvx30UsjDu7OPRDA4Z1/6lapkYHMjaPeVxYZ
FnVHWYfa70SUGjTinOHZQu+vRx6m0JevMF+wdHjNOciduzfy86DxMWVsjbCQ/LB5
vGZmaT2lXYXHtncdpvF2lbIRf1adraP/JHnsylsJPixo23mELK2jQqsr9THAuFAR
iD6pciW8lUmbaUCRUtQcLbhpKfIF73glG6AQksDgm+o0GbjiVmLVB5McJHSjZkMr
MKtXCo58/TRV9iyMag6e22OMTtMrFoeL7eD8QlUTiPvy0i8yPSMg4cvdglMBC48h
Y7V140g8yjNM2BNt4pVqPP7s/gIkvsuDvbBdCH0QND9pHHM1/wKyaHg0Kvlu72A+
GTH+GCiozS+HMnjJHd4o0AkfzCZDBvrmcW6xpbBhHKIjhOHtb2EuAH916N5yGxgT
bYVnP3a2lxRe9ePfORiUldRBXnpv3J2JM0ONWj+rIFfMQVWOVJRbBiNZGP+oI4eG
G2lJ6RANY86lNq83yrKmQ6HNrRQhFpspmDiRZ5rwY9Z77SfG73sdTDzzzoW2plTm
paHBJ43vplMSL+obhy5Mfn6Qq+6/YkW2ebDqt0aCPLtZnwiYpaH2u96kOBkBYAOV
aE0+WEeTCP6rWqsl+223nX71LhYDtGmQOygxYZfJNciV9krW+nVcV9XDM7bHWHcl
9+5k1yOEvxIHNH0UDSiHzQ66FsaxMLVXb8/GWWShHbLP39ui+ZuVFOG3FDVMnhfi
CgurojxK/ZD0v1nbCjB/impNydmrhWW1uksA0IZ1Y0LgrJno0iobUhr487Q8hNBo
B5LD4e0/GmEiGO+D0cYiODicP/h/+cMjQu1VBX8uU1P+ymQgrE6JtbXt3UplJ9pc
w7i4zglxm6Wp8yDyzK1eWFslUw9uZFDp+YG+0zAkRg5V3acc6re4pMMRNqILHumA
sxdKfmnfDFM3sPiCn8VT4z/hrjzKwuAbjXfJLbUj/BWkM+Ud9eNBLlxzzZy+HHLh
RQtEOC9G4iMYTqUmmNLvnqtMoMWI95oytJbP3MeTBtBOgE+NMYzU0/Ej0VX0eOnU
3WJsIlAWTpIWgNSPd8gkGGn/fqMiVsSSvcviiWO/jKjqTMkYz7az+/bgwpHyg5tT
ZSQJZZaqeJsq16XBsPyygzuhtyoYrlvflUBrtB4Mxedxe0yYzIwMXZK+pHAzBVpA
hSq4Ccyb8iPOJQm1zt0/OAmCi2rWNDAb8O8f7wcpLwBWPcqApe6T64HvqJUl1g1M
sSKFxwNbG6hmjFzpAzTX5MteG/HPzcSrhfsXkewJaSopFQ4ymFnTeh2osCSHTnFN
bDVJPQoPQM5O/5jpa2YKeQl9/2owQevu1flVOsb6vnBH9x/O1JJ444Ejg2JLACO1
AJSs2l6aoFMM1IHnAVTcLOBRwzMAenQwnuiyC+i5JedcKQLp3qOtJxiBNCC4iRjh
3EBTkIZTIxMIFfK0ZWXngCNdlaZPgslrWImFYQDRmMqrSFk69m6sQX5Mo6+oWX0Z
79oZPOil6XdCH8+VSlCkG7AwjbZT+dPVt/bsgCpEay8o50dTOUTAh8OMUMcSu/+b
zRyY7uHLc7AZBFWpRsYroKSBpXbwPQA+vThsmWE08Y38G4oIf+/2HeQos88vsbf8
3nwM/kB3Ax6hisbHBsmfuqw/BlAF3+13U4tCW64QiGlyeLSaGsRdcph66sN0tNz/
AhYufv6WMB3BM0Uy3bP6aXB9I6XVyje8b3DXhvnxvariv3Fj48gcjFycPm8bTEW7
ElGsMXW6d6isk0Tnbc3BX5tjo69lus10966cX2RN0Nf7owuPBcbl4KNA47kAuGwo
uBHjhqidA5SZuzL3seh1IG3Q40oHRVk6TTUYRhbAXEQUftJS7RPgkVsXyJLQmvCi
0K08GPbsmoJ6BbkxAnJuzGYfr+sAKgXLFMXzKv19k6gnMQ5UJVCAQIPyK8avo5bX
b5KDSuLFGnlmxA3JL3qlKHd/tDE4vZO5oGIEhMjHgRzyU7n9jBZFoq4V/7YYtPAK
S2zIkFm6v6o+/023Qxl5AlvozxnQzCTo8lzn+xnykpVXRGBigT/XtaqVrbz6WjqQ
9Kz9iJCNDCkWir4d5NU2YYwX7AgW7de4qY14c7XDoPv+3+W5VkIykT/jQ/jXjVI/
EU98+Aw5Yj4HHeHfHol1nQiaHUlAf0JbKz7ryDWabfStqFZYLCLQnl4zvZ5XoWaz
KKjhCfQY4ReToCTv+PXoywm3sulWWQKLH5T3v/znfNprlafqfhSsAW1889Rh8zMl
6meQTZ8xIXNmjHBTroigRUhS3SoZ7GLCbN/LzL/pHVQJnM58sBbGe32mVfOUloxL
GpZb5OGXhdjd8impqxgrGwIbMTLmWV1MIzimDMQaktLowovMhRxjFe/LwELU1QtT
GmA680rnbwtxdG+QzYAs5wSlMg6HjZiHxKOISMuW3tw8SMtPfxqBcTc9+tMoGBGQ
Q+rlIyv/QLUaypHJPijWWGJHN+IpdVXc00hhQqZ2bb53+utSMHK2O4sm22OejLkl
Eu/qAPsIMSNLtz1e/6zfFXhVLzXa0/uBiQJ+lNuOM5mNV2zGig1wh+19xNkJ2GvB
kWJIl22NNG3v6ZNXuMrTWHtpz4vYDe+IyLxvKrsu9gDp7g23aGyKOVUjpv6dbnGr
NN6ufW8YBDtdYVkjQaaE+HAMlxryE8YhN9TQpgzxnHuwzVRM5/1I57VqEeOFgMm1
V76gcp6YM5mAdSNi+7twsE8EtXaQd3bporARzawEHoUDgI5Mdk83uPNJvG81ft9B
25sRuHK/mIHaf5ih99RMie7i+b6HbM7K9mmZe9FRVHMetjPK88C3Lb7kN/MD7RhF
H2UxbCs8V6mGkL5JADXGbUpTjrKAMwLJ5bsXvjcIF5lo2jknK8BDC5dBonqHjQzP
vKHgopxrBbAdfkyO/iu4KLk8mG/6anpfDHMDmDJ8TqghI7Otp/btLVw13yp+bHw/
7YNsWCZ5J6Btv+m3LXVO/gIMZBv//zASG1S/5lxpsCWNTT419UqiIsAQIomC5U/A
Cd79mZiP3RDuX/jN3RwOn3+qKNlKET1E86QoUZ2YiP78rtKRVpX+sJGmv7N+iAXM
tdlL6PEDfi5fcxB3Yy51NpvCmdgJIJG7v4rl71CuVvHoxByZCYlQxC1oGsB5SaVC
lsk2i+St82ic8avARHlGvqjc6/6v07cedi8RTnj9MFFCqRQf/lfvBJkiChjdmPe8
kYiVOIWJHwI+IFxKApl39ZYCnOeVUQIHXdswhP50p26+AKLzICryKz2yHG6g2t6k
mbhZ+R8/0tsPJpGSy+mx+xOfRZhhRc1W8DlAkVYsm5ajZ9cJacqA5LwQeJyUf9P4
GnBgj9N4O6panvBknFvmIFDH7ZwcPbar7mnEIQgAOqAD1raoXKf0zoAbkuC/DRGS
lLX2xsB1bTSTjFxA5dnyardSLcur79alRKPWhevypsr8SsCVD+HLs2lAG35zWfXh
0jYEgdhadMby/wXcFhJhq0GNqZH25jUYL/rzJHUVdIdptE3TiG2rUr9H3b31UW88
EkUsUbtS54ArzxVhI+Yr1S5gf1KDDlAr/XEBOIrvhLoIspAbNG6LOBEVp4UZRDYM
q2wMzjQrFjOhftMUYJTlQ5ZCzn6zAfZD1dkUFf3iZievWV8/tsFtkykytbm7yAVa
azwXsmPfI10W4bqNFWNcq0IZu4y7FJuTCa9RjeYBU6cwUgkzvPy7iOnIkyh4r/bv
tdBWqHkcao05OtBnUUtm77vneLZnpOUXbuqx3jw3xNq8w6VPXFgtmlGQa5TD6wZp
BMTXAL37ctABWW4GGpNdG16LqwnWlmoLD5BmLhP1WUUu6W180q4GP3VfHBbzYKX5
flg/XzfJKWw7vXFBdASgwxWRx1poo3Dct+nYDUhrzONGyztBprA1G30Okn2YKlJB
ivDXZF83bklVO1qCbRkK7a/+9EUJuSwoPDAF6p2F4MMQUZY1KssxRaGGO51cHKF2
9aMpntxm40Ilhy92vgQn6l8Z22BDyEsN4QPoGuJOpCPEB88yOPYqTefw/78/BSMn
sgo3Dq5EBmX5JTdJ49cmcCygfOj/hhyY9XTH5jQ2IkyDYvolzXkVv3WPnO9Tsuyf
W4NP4RS3vNcf4h1TyJ905K6iFcRlXU8Tnnj+1QIvBCxuJbjiHAGhd7/uI/21GFa9
moAoSo7SmWxMvXrkcTh50pHJIvyWcwAM6hjimeq/MVpK5JEapZO5bUH0Nf4JXv8J
3C68R9TJVt7jeI6sJzxCYh9t7J15Mb0dxqWF4yqdlCVg7+X9BGX0erAKhtquz2RB
+YfHsZ1tf/keyUFqw3QsUF/D8i0l3FIWPVik7XoHisZ8Fk0RfekQ7Q1bTfL9xZVg
YRvFbfYc5KAGx6c5apmvHJ2U8dnYYzUTEe34o5y2X7fnEokJ0TV2VhDRZCYqys7T
CdpmPWw5AQQ9vBuPGYabXgKLYwTe0CXGBHR6V13KFxGbL8fRl69pNbzb4urb7ogF
smB+gvTdqnMkA2fERDurHyEZ6jb0CLsHwNSA2LEX4SX/q+9ouPexV0uWaj/thJek
yh8swlbbLkpxYvvEMOJYdIomnePFfE8pm+3v4fk2WMgyl1dh6XiP6TA5cD7NjcJi
HKvprPLcZmnSvUGj2yJIDmZhSSvLe1usYZvXbUUTQdKyLbLDEX85J05SUXnEdvnB
Dfb/QF9gsF0PsDkbSLUOoeMG17bCbIAb2SmmErSAMkpDM3ZUmgZUhtxF6vKQBtVm
/EUDOBAZPGGZG87+ZNrcUYDHlKGzpi3GiX6SC/NrkxNE8XlryPu/erHVAG77iiji
STUbv8XgvMj7MSYRqMXz3nNv0M/snwCo/+M0UW6AeZPboWoPWPyDrFoCpWpchRHf
oV8Tk1O3YMJhP16TvtWpFVhO83IZ7zxfw/gOqeFw56ZJ3pS8U1+6wHpBMazhRx9P
U4tQm2g3kztmBrnCDQCmEcjTOPd52DVtxc+X5e4amOrFUNHzeIQoE1pw8GYWKnE2
asG/pG2lFw7mM5OUwHSdYxEH6CY62IoiplpMjRkzahAkre+pjWVxz+WM4jWo4jWG
eMLT5BubRr2iaRW/dJ2ZwVRMB432yuWHOEFoSPzbUYgYK0HJuLtY65prkU21jpwu
EjFBKcoiwe+LaXLZDh9fwy376IWsy2kWjgaNNTCwoeSehkPnkH0BRuc7824lrj7y
phXp2df2dDQQNLCf8ZgwZHHbn8WR4Sb1G+d+St6k4yKsdRKxn2z4+b1XYR6tovxf
yx/wHrKXNdOIxDRTUaoDiJGx7QbqYSp4RPiDY2TcTjVHCCsnTjPjXk17peCvzBUL
o1tjeGoqUVdWaIcJbWWjAFu3jCKFxR+VNgyzv99yzJq1CwIz1MZJBbXSXc6m75KR
SxaBf24Z41jdK70duCZQPkCXOJweGExgJRtsiCx5RePhZ3JRTouZ5+cdPzdZMu3r
BcHXIFCpDn1haH/9L0uIiWMes+fITYeY9sGPGLNBvGrI/13tTHCygu4/QlbXH3A/
Uq48RwIeTnkDZsFw/B31ldsGM7SaGxGp0+mj4crWEvAzfhdyLJvn24TYUpOdjTo6
lnIQaLL4uRdk2zSgGUB1BW3LjHdjubyrl0CvuM3qCA3HklHmdW86efeRt1oWi0cL
gA49Wx82HYvx5CucFtxij3hXuy+4pRZ9GDOLYeiPsDRYqXMC8VT89gVsDK1+Rc26
07puMrw66jUxV78PQ1z3Aw7/Cl0y7bOGjW22jPMxeQWgMjxAE07nLqXHBT9kDkGn
2qEG5nvu4VouCG/hqC1jpCmlOKO0pZ5EJRDiZ6Z4yCAN58Af9RvCJbdHE6lYmxUt
s9dbLlS9+0KJxnq5YiJfc4MqvMTV8bCcD7A9+TQjUZvCStl9CCb9l1JT2NIoHzqV
d6Tx27fQ7nFWvbsHBAUVSDn93XH1fZv9/L9IwJdLNf8lLBSY/DAOShvlrLyy07u9
m31GgIdjlIMVyBkUYC0sB5+x+8ATOg3HddITd4pKRpd/iuoIh+xB6ffW00vBz2vp
7FmziXK2vf5+7gx+clJqVbEOWRHxEotXioT1P01MCNmoWjaK4e66jLMRjZVEUuG4
`protect END_PROTECTED
