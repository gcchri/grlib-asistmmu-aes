`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PYqRTuIkOvX6jp9iOPIEuy3FQ9h+enwClAQ7k3HUbKAEVh7cqzuoaLAxo6DAggXS
+h2wS7AZWc0KkI0Al6Nbq2NlEPSgtl3gE1glwhl9ix1hg3TzgeU5n3EDJm4JeuQ8
brNj+/ld2RYVt7iYWXv0jDKKlTBFZ5XaCZj3yEgvvpGW461GMA5nCaI5QgjEI6WO
IwQxYOH6ZByHstsVhsainO7whJmnthAR/UkKaOdtLYGe/A9K3lh5wB2+gljWYhqs
8Rm6rKOfbDKiyH0vmz5cabvv8h1QlOJ3me9Q4BBTkmJowbluFJrWdOMuNGTXBgA0
V/E9wJuCQT6mq9ecn/8tya9IDsv/KxJ9yAfHF82iijUIZNxX3+7+exVMj8IcImGL
9QJ/HqyByvQusi1kjJkghSxT9ArHrQ+QoH+he6Q4d3MMKJ+vO2Y0RglQKgmQoRKp
`protect END_PROTECTED
