`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+EecgELAY36ziMtlUDRyuxVfHZj28/xmxvZI1WMyrSlQ9KRizQtW6ZfsA9O+uV8p
YY3QFK72Bal8o+Hdtrm9LubL4YtgJ1B7j3AkVZtlvK6raP6BHA//L80HOZgjvPip
dYyex9uD9lfOzo3eQQH+jzBzBo0vg7AX16kqDr+bLSNbLb6pxqkpR/RhSphmVYhS
4Fwj8VfTnzcKTYuer3OJ3B0MYPD71fIhZvufCvQREz+DB0sFjrAoAbaFoFcFlBNh
5dXN4ULbN+1DPBxjS9EPtvSLLbpbKlBpj607Pf7VpC7dLMUn+3GqQXaPpelbAJB0
enNWhBnI9aoJqlFz+XESdL22jUhzDezmh1FoFhbZqIBW0NZxPlLwEUv2IpVXlxSt
QsjZpnepKCq5w0i9tDE++DxaEAwybLFXIcjuOACVW9amsq8KPTXw1VNPW/b6eqlE
dqFmqigtpG1yPHtaD3PHtisOS0pkDGqhyxDLSJpDofvPHtMHre78YCtj09ShIOUs
XoR2YH/rZCpw5Tv0848q5TTCqZhzB12wl6IC6rdFkk4EtLTUxeFRHSybiOMxxNNz
y1kwHyuQcDl29kA6P0QDEA2RoE4oE34vhGN+FAN8t5JkuKVGRhigRKFyvSrUp5Wv
EA4mK2GdU7eC0nuXm7LSFVfYlSiY499kTt3MI5zYPmMYbqNgXxlq9XrInb08Gn3T
MT4tHV8co2poUYuz7RZZIgikp0NsRvlN0hzKVeQghP4nLpEYlO+sCLnliJfbvZN7
/MGKbdkKWlqfBdRnp19WcD8ezHQg2hDhngBJOjS5q+fxN915C9ykW3O8dg2dKqyJ
r1vx4ppzqlQlLggJCrrxMAbcx8p0AbsgfEH3YX6pPGs6QXMzvuNkrmE4RsFa2rSB
gPYMW/W5GpGiUvwHehOwxDW9CKKQKCvPUjriVjjr+uGWG636tDnKHFD7ssmW8B0S
T80FljvC1hBdxMdBy4pe2/56OisSyII7bNonrUEQN5Hwbeul8rMcIm6P+z9ifk6O
SQLDw3Vz8ZigGpFPiPZ46+a4bM9iMPCk2nLtlc2575UBKZbEog5vr+YqbriOUvEX
kF6nMlcK2Mwfx/xsmIHJxHq4sPLA97JnVsfJ6TAUjxuQjD3HwmKYLj1FdmSF/4Th
DE/VAfhMMNZTzVpxkMePL/1on7lhxnn5QY6ZRhd9qXi4WDf8whWBKSn5P1l/wPBU
RWmIw1R1sqa3yDOjYl0G0JQ10r0nu6m7S2HrY4Hr32+mo6Z2Qy7HxGkFK8Yjt37m
3wfkE9Z/ED3XnD8cLpcgWWvqM0vu1Dz2vJzPjO7kaIFatGW/6nlGHfeW2+8ufiYu
0BXPKvZcB4w7mnCJfA/eiQ==
`protect END_PROTECTED
