`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cVo2MpV4WgP7gjpnG7FJHDLjH6SLCYWRzrzMpnb0kb1SLlocR+jSFOh6jQz3lpxC
SdJ/DJxy6yR1wec3gbkGvMBKqzghsjuDS3Uwz9LOGUDShDI34Kp87zHfcxtahyWA
cPYh12wHd+r6L71iZfKv9kNytKSDHUBWMU5dtCqiVrDajrjZs++bAxsiJtEG3C5/
O54D0eKeB8EiBiZQZGV9YpQS3MMVAdhbqkY99UYXVWruE/bnfsYNhDAB6qU8ELR2
0Ul7VXwCK+2K/aTUiIV8YpCHNkTk6KAvoYPmq5ixxUDGeZU1K+fFDfVTlZY3SYll
HcEIsA4+bAkoXF85DE1kuehI2oLvNvjKUnRNiKzfAiv1EY73/Ksxvh3e3KtMC8+x
jEPmWc+mDbJC7AVW8ul/gWpY2/vi6AvdOI7TsuSo9lo=
`protect END_PROTECTED
