`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Ne+35uNncS/V/6Ndt33CG6D/qIrwANWhjh7HSyRg34SveC3wt3vgpbdXDpooXxd
B0No5fRgcmHHvqSf/6t/i2AJaYyhfN9vR8Febbiqq+XZsDbc7q9d8o3KSR2lyGv7
hVWVpCuNp9E628avTjWPbrqNZ/tzfldOVH43UDcI1424GUEB+zy5NU5fY1+DuQ9s
Hy2AFTc3YD3o00z8undaE1Ax7nmaNMzT/TrPg/z2gBUuLT8eLFaVApy6/mZbjOql
hhOxCuql3qC01F92a08Ao40CGLs9B+auHtVU9T1lxJFqOgLgrMqLU7qfXj9FEvqM
UPku22B7ffDImYRTGbLAn126qfmBqAKpNOI5aId9q3z7YMwa7E3mOrfyfA8OM6H4
FzpC7Gz13BXd5x9CwLKNGw==
`protect END_PROTECTED
