`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oXq+6DJ+hMcoau3lm8j2CLwXQbwHGzfdt2weFt6mdcyGIh8BFKkdH3wh8SpaDPTf
iDJDPP0jD+X3wgWoQOvlIXneY+KG9IKEXopLeGg6A48jTsRFWB1Z1MbOGsFVJ3v8
5HfuE2/r8YXDUVSghMFXmtiwl6oPvwG53qmhzBOUgyWImYZ9QykBoFmrW9BzEU7V
OoXB6dcpC5dpVrO2kYWImb8Vb80gFBt7+8AOjCGUImhV3hvBoX+Mv8dJfYTNLMy0
TQvov5EU4ZDgl9EdUx+8ImbmwbFfGftN1Z2y6GwHwlKsw6XBnTeRFh6xw+cYwZox
j2Ke927XAjykqoG/UtERcAbrMKhd3W8mi5BGtpLbvFd1WsnYkp1ovngordW33F5Q
McmCnO1QMUzeOuC7tc/i5Q==
`protect END_PROTECTED
