`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qKwno7itTdyaobzuPhD38LRRbjcCmH1U22rJx/PrNaIAF2d0AkTydTEGHgzSeTZg
9NNAgoZIE2t8A5CVJyGezcZkvddEOCM0SHEk2vo/ycgIqfdLIROHtVi2uSJEJd/m
m41kMFGqTNQ38A8/spPFSDtYxENOcac3y8LKEBJZD35iJxFJbyetSeRmzj26yxqB
sEbEs/lcjQGFyBb+pZjVRyVGXFYuruvWykaSS7IArpOr0gKq5FWrefnsluiUkRVQ
OtOD+kza3WXM9wsHnq7iirQodboO+V8igUW5I+FF/UqzF0NmcAm2vLrJ5jN+z0aS
PeelTwMEb/eHuAdph9tubYdPoQ6AfHo6sArhqbSA4DbmH4BOYZtpgffZAZ3WmhNN
eVKx34kpv1Rpu9zmqJc+Y7F5t+M3lshYvwMEOB5m4CtZyPB9FGwdlXKQjTquAgWr
ZC/HWzWP01UT/muQrfUGUGLQk9DezqnxSlJc7NEBTqRE5wt5pj6vxq12z2DTL/C1
DvsEG70Y7F8GkrLqz0aCLWBMtON921iYr456MUsg0uzXNiuha2nVhFEkfjAu8IJu
ystbMavt2RA29a58QJLg1VzmSWJ0t5b1uehoJViLprUsUrIIysZjOzhfzZwHcKAg
ddCFe3P0Me9bUb9W/n+zX/ZAIANWeuSLKlErZtMVlwwD+SJ4yJkWuvshujTUHlsd
UGfQxBKHGURiY4Y+8ocHB2R4bS0XPD0NiuA6qTp2cJ+29C9Xg+ynUJYV0beDgFR/
+7D8JKDGp+2GCQgS8uzKSTM5qdOnlEb/8YWy/2uNjeDmT4zJ7vcNpNbs6QQP/0Yx
WcdIIXC96oD9Vb/GNjY9nO7c1XCPizgfEg2GKg5ZrME8scRtUjHKoOdBDupJm5ih
n5cXEgFwbbzCZs+nkH++lYKkzy3wnfK6GxlEIWhJ+GB+dc+zJbXfcB74TGiEzbjl
83lSjanavWn+KS/JG2dd5i94x0/KUdIdjR6KyuX+hZhxCtflbgoI8pFdvBMGADs4
XaruDi+lMRKntj2v0BA60HtFqbuHTS/TIGk5f1mZjMVuF80u0oi5I7ThFHJHkLWV
YruTUchtClX7jczaXPtG+kIsfrknRCPWz9Le/a/vqXgWISVAyW8PZ9WdQAT7apJS
IJmpir+kFK20GOC4AfymwzvLG+yYFQZPhooCxdF/i1q/AhVZrMCCKatfPftrLK8R
D8686pgidDszmIcHYyHmeEO0P9CahhBusLh9VoxzN+S85pWHfdRhFkY7U1xlVeTF
sY+VqaYabfDabXCtxb2gd4bcZPo1D0R2HZ4UeVwLsB+AHTanO1XWyFt97fYqMUT9
T3ovcVMmxOgOMNETSPzWi3hABI9UhkzS8HTRafup8RdiSOLpLtjG7zIi1c5fM0eu
WhV92ABeK2wc52Q14KhBa+TBXOlOjvj0Jx71Wfxyx9S6UFtO6ja6jQ4HVWyZtWHq
SqNYgapM1TWWuCPYdxPU724gq+C5tv1gLtCFbMkot8jg96t+/5QF+NhZPWPtbd+b
jj1oO5OuFWfZL5brKm27yiqJJSYlXqfWtYsCEj8ML0Aw7PRXrvYIRGhPkPMiAvf0
Vq/cnrrS0B1Gw3xqTBtj+B/f5j26xSsQEEuZbtvXqSZDRqs7VrZ8iTgXuMyeC0Bi
78lvUrgSYw7cM279+7zIsLpLTb5o9KmfQPCHMGau60ToL8JhBnEW5Eb9c4XUYtBK
n6j42T/52nkozuaMCysdkONHO5m84A7ACOZjcLyS3+0qHJunj5wTq6e5ALGgCSD9
5mx65VMASawFYsZWE8DZQ5CaNaISrDqA33LUWMQEUc0YX1zO1WtmV8zzsXaPXtWK
gVwNE+35EZs29tERpiVrOBe0MDz3HgOszQHbfTBDEpnX0uPE0FPfCzapqF99Ouv5
6e7fviYbc1REuFWdRYQRVDlN3Iq6WAwFu4DbByavMQlgVeT+zyGwGGyR4w3YrfwW
ttH0Hzh09Q1e3cWzSZFKr64M/CbcD89qvCy6PEXC0XdVcfxsRO2Me5NyB0LQ0dPs
K5ofVx+Gzq3EHAtSluKWtAeKQohJNMwCuMeZnsAHrnFSnGul3vmbdIXaf+nyVSEc
UCpxcXrUx91+JmHcVVF+8R8XvYaCrYW1Fe1ZAi3IEBSsID3GWIszuL7ZtiT/9kRi
W8JmmWi+RPnl/aUUHwRm3Q==
`protect END_PROTECTED
