`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UdFhe6xrFbsihdp32opfqeut7gLiav/IbpyO74T8u/ZwHfl1eK6b24m5HIkytrBi
6VArBy7Fqt0HWL1V4wciQyfgbFYAz1HjmjUJLX6Z+1P6kA2cec7UrNJHcFVBi8ny
W33bqqwKjGEFi9MfU4sSNhg0SgNTfUrd8Lhjsomho1eFEG4Br55ahrvhJ3U6sG5O
zlJSEbIbDmik21GAMpEfR+JXaZ5inOCZyCy0bJWx2iUVqoyFyio500bWc2I6egLh
9SdIblMn7wpbm56gz/lcV5Hf+B6PMT58PQecGMlV9JjNNASlz2E1q4DR7Kyiiji0
2BnA9fZihikaOh87r9NHgZFfTUWuAiRUtNZckkPYGchxryYveGna9/JkCw4sfYX5
ciompfX2zE9S1UIMkJqL3s/FYhb6rC+VhTYuRzZt6WXpLjejMXYuDzsM0KE8nbaG
tZ2/fZa+mkLCibZtmibJBdab5YQr6zMP81gtrEtBVQVqF/b6fObiFNkc7utdDi4T
xQ9M4iDHAlHJEn8+lZ6/nMYD3R8C1Aoxu4LyQAz2OWUY10yBpopB6x8Kh7i9Wz4t
k44GusycRUTsGoWZuYLe7ZOps5CjrzTYtjcah3yMd+2CHnKfvWlYyYFnvJFBKxZw
hEEWbePzXrA3Qnqc5ZT/G9HxNmu9/zKZbHt3mtiDRI3mDOf7Ls1ariOZfjK6RNZg
/4FUIxLKh4BtHjSZW+PcmS6QxJmktmiv/XB3SXWqYLOzSckW83kXkjD4pyJ3sIdF
y60JcwbAFzd9HDZUuR7Mu74Q91W9o0jXrKDqLYhfUmqZmHQ9C/ffhoHX7yeF1iNd
wvSkYhX9JbKs9dCuViXssxzrmIv5nU7RcwA5deYjvTqYu4AN/vMmxOxIMrtTCAIz
uZQFilmuTuXfmHLWVmoaQoEeHIkTULMUw4PPN9CT2t7WdPbOVJxUNZMd2soQrv/s
yZN34fek/bhgJQHWlJp0cA0nOj3K4rDUtkEsTH8tDO6yaMuvxtIHszM8Jg7xUo1e
HuWEExu43GtaGVOBS6MKi/hS3RGJ0wmUrLZSz1ih0l9cqxJvK3absaMWkgPcP7aD
D5B6jvytkM0wXYVDxTeIpGCWWPSNGV8pjaMAW6cqi2t66Y0tCUuzbKSv+ZbiXkpr
eM8sUmOnPYDTrfR8XAHgeXMWxRUAtxdV3FhO0LXJxJ/qPabQBZlNHZMzPgpMRRDP
z8HBHsbTBtgFMByw445Gkb7G0U3frcE98DlLwKsdQjWgA/2GPt/Pte65e2mcUQtk
8+/bNM1ZvEv1BqFv0mm3Bl73mjzmECTeYj0QJbpC5f9TlPH3DSABW0yA+LQZT9Ai
mEI+b8BRxbg7OSCXE5CNcOjlb1a+sdY36uqBWZIQKiw1zHparTzUyHbfeQNLa1d6
1i1DLPqGMdLeE71uCzOwuLSxudDo4QOOev64FMmDsrjUnFAoQmr6rrkduo08F5D1
jPQPLBT9YmZ/9xIi+VtN28tvhEkDOD+OFzj6cvm7+x027llbcCI1R/+2fvTNaZGg
HwS2YFkPbFbpYG0ntk/4iYX1psJTnW4upYk/0RjZI+tiYL0V+eDioYpJuf8WRfty
eeslvAu7ZjAMAAREjRhZXdquy7Apz3ALJOZfSkMlubjHQSsJ+4JZVv2WQH3S2TGw
GqtvVD2rqPG9k1IvHAjobo+S2i8Vzwm/AazCinouXPnshbPvNlp0GzA0FNyjZWvU
8NEEJ0HnQtMADd8I4M6/AD9WT0dT3nrkov74elrHrvlNbfG+uuP8puAoih30V21b
3sO20PrA6uHdB1Vx6x9kiS0wyGh3g36Whb/dCD5r61ikXaSjjZP07ZASR4BTHSTr
An/XYnpbvSbGJrRSq3jwehhWFL7YEam+T4clSwwGs7bmKEHuVag0HDJ6l1I2bqlg
euwyqYnPuNHK9kiIjzQs8LLXYM2RsAaXTelniTLgWj0D1W+MeFPHxM2qH+Vz4FlM
j6F85Y2YFpVDYqpk3xYAnT6Kbwtq2WGITXd/g9qcbUINdYIw18iZly+bT/WAmmUM
HwdS1bKffw6ZK+F1zbr+/0DmsBwi+yVPAcT4/Oucak7adr59GHgsnwGoGtMoPGTz
b+X1LuB6hxW4zL8BdmWYrAs78rYL4CSS6M+Bh1nzbylGe94FV1Q8Wcn+9X+Xxpx6
BSvRE5N1UVQVc16uv8CqvRDWMLkPgqiT2Cho2KgnW1USmfM45YdklN/ivpBghm57
GEumLzFLwMAx5AM/oMqMWV/LLzye4aPf7uTbmZTdPqbbLtj68ayiCsgdCUp1CanT
8KWmCJUxVFT577n95tzh0CmOQZbs1T5bHcJ4gnqEx9YZm3Rlmr+PpCIbpX+OiD+2
YpPY+lDW+x2Qt/iFH81K1e364hRNaVQ1+5Ws1RpRKME4n3aNw64CVnEOe8VG2WEA
mH95zMGzwUFwlkWjkoYeztet5A4HaMUbn6o0aRpOx8/PZ1MhGGopICxKn7eXWyEt
kOqvZfGqrr7wRMUHDO6+nGfjVysv44sc/hBH682Bs9OsiVxTyFfo5wHd+f5u63hw
KrEqjyeZthMzZu5FugVMSDdP5V6LdKjUXnUREjCBa092oklC0najuYS+5jrBZx9t
IHD5L/UPwfOkBHlaaEHKwEDKw95LLa85mqjd81djxEV2fKgjdgoDgZdhqPWCC+j6
EsMwvPFBdr4NvRdXmNFSC8ZTAR//9ZwotuvpEYgVAJGtJZymjM69VQQlYRw1fvb+
Pv0vMR5hhrav+c0DBB79rquGp7EBhBiraTXV58uwrj6sPBFtud/2Q56RS1UM5k2s
F1VoZ4/qViDZuxwWrdNeFhoLkzrJPYqZp4+GDQF5EE9Tbw4kRB7uwkH/DIcEtqd2
lU3F0LP/AHGBgjMc/HwC+zT2oUysTaPfm4IMX6xGtYS+a+rOIYcg5oP4rV2gSDXW
2lwM1skx5aKNv3Z95z3ME+OluTObRGKqTYECcME3yG6kzVOhCT5cnkfFrArdSJiJ
qeyKW5yCsrrdu+jcfPL8FOYc/vETWUVdS925lYPNJjRS1K5/wHcCAXHaJOLp6kRu
zonZBgNQ/5xpVu9iR4X6UdorENRyuRWMvkgrynSufv0C01o0i1FdNYEbYuK4WF05
dlkHg4SDcJRvBzQUiR2foRHlOYvat8I6v1TweIJVnaXFFc3K7zBCh1ITpoKeTJcC
1vGnVrfzzND5U1nPi4Mwoa/zLQc1llb/X1MlWcJwg+wOJQEhOkIe5fDI2Y8lJQRi
19jZ0M+wfrYNRiDIHnmCP/TZkZT+jaFQiOAwVf4ZrTd8Rp0jP8myYOSM9IU8uT7t
0CA7tUfRT0IhmnsalHogINceX0Fxbp8osy2qzcl+yccTiVhqkSdRhZDtsG4dz6DW
BAXxzHbp7R48Y3BKT+01x4ru78qsSlqLdT+GcRigse2ISO/+0zGHGlrcqDaVM45O
pxWJd90gyhqHDJ0dFQ228bhd6Jas/15+rej8QDaaAtbG2eAueTee/KRls9Sg9iCG
04bOIIXkSZpIujnIHIrpfZ/qvYmG2/dhBiP09ISm87pcSpYjSOMUomXYAjSi/NEw
34ihx2B1OGTNZa4sLmEXVozpnfILB2hnwL7fegDWlVUbGx9jj4S1SUyxCfUSxy3e
pP4lBLJ561mPc10/tcUMNAb5VuqgH7IeqUhNkVm/GX43dmL9zDKcwwLudpCRxR71
BMuUIfROjII6zqxTh1XppT6lpVh4UjxUhMzVzQplzSAemlh9u9jMInDElbixb/82
02EbsvohYDwxIjqCraCNgcXeE32pmNGwB/M0x3WRKDkLMzl9v2eJOfctbj8xSa7T
24CAH/MFG+x97k4Jb6q0umbgfKSq1YTfQ5Z5m8/7g68ZlfFa7kvQnFW2TPTMFNBs
7oUDvRiQzIYrnC7m29Cq4oNoHA3B5XYsv9bR6vAMCCwsWZtjB2obML2ianvgVbwN
vzobVVgfUekSE70oF4Oi3BC479+z+vJKic4AcxFNL5Y0lKNgF1UBz1xAvepbm2hB
8GzDz4rDGBGAjNgQMDlW2qkjGpIxv9t975jnCaSyGZydZCZhFBMmeorIXMKWtEgB
/jbuY5tFnPjhsAwkWVQsgJZHslCWUnes/G+qfPZAX0NrXktJAhImysfKg5mE5ZAO
iYxayDCoKQ5ce5RWzfcMYxHQwWVzuS3iVrlvDyPLzCcFbR03ZEHs1ENOxbkfFpG+
nyWWy5SnJXB0scWU7Eu7DEd97PwhauhcoMGPDTL8VIOOgC52WO45qlZ9FD5Udpp5
UdOb7njXMy3gIG5W1ChclxJrDrm/veYBbxHP1sPlL6z5RAvicN/Ga3nC2cmBx5Cq
SFDB5UMXEflF4okh6oNYY8sh3ZC0aGmyZiXDvOdWK2KOSM8Gi5sTjd6byJuxxQ3r
/b1n55851iWa4WJG4EDtQnFqyMJ7MphZ1QvRhsF0FN6m12khkYXFkN+WKqWZUVZv
kiqoZeP3hxNfFyk2p+9+caqJzGF4DFfuAh4sjz32dGzB/WUvwWlFcv9vAfFQ3Tpy
yXpHxjFnTJUTPO8Lb5cUHAQohyRm+Ia1+RIp7KZR+ZQql9Mmclp/vw/Ob4DjPSlf
Sll7gWwO6Zbp8niNwUPUaLBE4bXFy9Pg7ulYVytitK4nig5U/WVmBSbdtXeo1zqu
RM2D5+kP7cwyZDTD3mOUYFXit1uqlqn31bNdY6uqK6vv9q3qPejswHCA8u49a6yb
aS+PD5wdhww8gp/IhETGdfp61pph8MuihtL79PhxWrQOiyqT9LMn9UgjBF5D9xof
fyYNfqCJeo1vPQtrS2KkvHoISWHxaRBKlu1gCckHv/UjkjCs+v07XAVd3cBX4Nr1
q35Mt+BrJG0/C0HCv7dyi+RkWtGXUGbD+zdH7/UOUN8gryQur04GTXHAMOCdVYPJ
GV2HDQszxswVw53K9nnIdOi83w5vs8Zhq8iBQ7O0BBHJKGQRnDRfl41iOOl45/3K
inDSybuH52hSMFDvz7yfHY9Vt8Q5vWcZM33nOltM/LvazTX0YZ/lqn8uf78yeyHU
/4GH9WlF4LAVW5nzpOYmS/gLuDjJ/o02rvJ/OrdWkyrL1vhWKftIb+8wNRMftgk7
N0Sn5MsEdoHUlzwtApBMxxsxf0XHh6WNF4S+mMyHyu7FBfcRcvPlgd+9wRjTb25R
D6tn6GEbkXMa9x5Hxx985RjgJUYt15p+dpm2JqI2PrRb3mG2PVUIRiIj2z9fmyFI
NNl1jey+7OydX0qClfTqc9xNQApFcI+xD4FTjI7ge7+OtpzM7/CwtO7qxuAxbWXg
bHJMSyiyoUqe25VMLct2Ujiv81fyEKpgMIheur6s6Fd6veVQw0nr18zBIvcFCnq5
F/nChMa5ur2GqBb62DcGCZ6Xi0rNNf95tAsmefloH01019oTVJnkHbhJDSt3Uzl+
ej2kSuPFIFdVxEntckj45l2ZdfTtPN9nuoV4W7DzePvDJe5B3mrFWSp/7DBytfMd
Y2YGaYwBrj2YfsVqQGJ03pV1GlQogcGcfm7iupd+uKV1SLpao6pwx5qqLDJ6CJC3
m0ZaiyUXwIIS/33qACA8uBux5zUXmgR1tqUo4jeL9ZYp0G0padEejnJriY8MsKwP
wG+vb7ZWFBmYN8bsRCg1gdxsY99896PT/sUPR/lKjQQkurMI37GD0nb7bQ0b+scU
wOPMDZnJdwh2UrxazEOiWfvejzAmLL9Ws9G+NuaHLogMjijo8l6z6k/vsNM7bUkH
+4ucoDXNbL/BqiyuZXe4ak5uMxUa9YRLRpeueciqE71hEuQ95isQGd7tYGRBueQm
Z7BULAz6mL36PyHWfS62STUOKURmGAIjIiR3jjPqY5RpzVpeDDxu1j37TSJ8QF7+
yYK+avTREnOqbNQ2tpDoP6Ngc2/s/hYDqjPbWmthboOxgGJwh2kvSHfXOcfyEojX
Al0nxL3ZVqKC+32UUfcefsJ/sRs0uEXjWJPh4fNx53KrMeSPdaCiVDSgcOsPWLqk
trD10JCA8NBLhnwic+BYmf1FgPb69F23h1DYgr5zYqhOJr3sXWvup+GZ2HJXT1SP
R8DycHtGZtM0kSVfq1YES2PJmHkXIzKcWCkfmeC6l1XZhh9s7g8ZUjpJ85wheQpF
b5txDYA6LJkY4T+E/5iH98FqpKY7GqqwooW/ZLKM9czBXzUagFjmkEF323fbYICV
HaRqvicaFfjM63tJWRF5Gv0jJDqWMomWy1MWSJvItuL5cyahx4caLip7ZW80+qRI
QlDn94pry2ouUJ0G2h6TC4uw87nhLIHLdF5t/LuJ9JtO4heUCm1QABslJjjKb2nt
RsVCt+whMUKsuEMz67eONbMMzS7xFqa5iOcW7uWTylq7tVONzWjOt22M9D2o+LKt
31V/DbCXPnQ41/29OQBnA2D4H/ZBmJpTp8Y77CS39QvXqfF/2ObMSkRtuvePg7ri
igHv+/O3zyrIPq/eninf+5XbCTt5S5zgTWXWYk8IE3aSxMDx+i/3WC2CEFkihnlL
w9fucS412twM0CybrcKA1b8s4HYfjWZMWYzwaFg4YjgV49lewoeY2peZTA5eyibx
icDvySW129jlQVakCilWhdTM3lwassRIyC5KMz6sc4jQKG3Ty60m3CVo34woEM4G
l1zqOmYyX6sw3yW9lNJHk7C3kPoRRhvfTRJBnPKiLEwzEoJaCR2NjCvK1G9pzOy2
f6VH0G6ZS2LdmW+Oj1CJdXOyAhk8ATqarEMvRfZBWnAWkkcnGdcHjgAw3mAX2N9u
dqRpBdYINKSuF+xabVMKaHhD7J6d0pivqGRXZ5R2KE7VcJlOSWI4jSHvEBV3LpgS
hw+lctjMCRldzwbQMtx0rad4SuNgSDZ6dK8U0AXdYGQ=
`protect END_PROTECTED
