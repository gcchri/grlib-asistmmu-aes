`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y6UL5GuYvLw7ZMEi1nlY9o6O2X669feAHZ64YakDfW1sG6RTQDWvg0LNd5XsPy9T
lndQjGhtSLkQhEGijl+GFN1ag79uBAdB59DorN3nhtBdBP8uC9d606VjYvphIlrm
ZevhTThdvhuXRzLymqQi2WNf1hUZMvqx07wE0TVF8eTorQUXI/v3sh4Ag0EQsxw7
7oUyKXAyPbqaXiwZ+Q/jVGna5S1DhLL4wb8CYcWeFN2m+ybHg2QKbZReEuC96RH4
Kg0yjS83gkzBhG5/hFVrGjLhLgd8qe/DHBe5iGAv2iAdM0pc3TvnhDCg0beMyD1r
F9DUkIgVf5QR7jqRQEtFuJPJX0vEnAA9mF54ncF8JS971M7J1j903iMcSOuDCvjd
2J4zCwwionWE0jtV0VQ481ZqJCcvChL5Rf8ZMoeb4Kqg1Z4i6cHe38TpHcD6COsz
`protect END_PROTECTED
