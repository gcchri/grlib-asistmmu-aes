`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SvHKL5/2T7mv014rHp1LZDGUK03kYaiHKcV6OLBVPEaUzqM3KzImK9VRml9znqJP
Af9/NEWBJKK5qkwgS35V3fksbG4csyhYsPDLRL70VyavllPMAKE4LcIpHeJLmI/I
n3DPjSJ6oiTt3ywfsjLsYdtxUs/c6TIOILgA7b5kfLmHAdzv7LIxhsLziJ43vwCI
jKcTEGLNuSRyzKAV08vKM6y2eoYsXSh5a1hZeNqPZb81QpsvkBMX0c/feUX3CP8W
AmVBNE/vJsr3pW50CfCXdFKdLvkJcsV552IJmDM3b6/jT1rBQkjQWKfd8jg4AsoU
uzxFpyl5pgIt3/OWakQ1mCLdSVQkQWMYAwLJpEbqStlF5k61BWtDuWICNc0+X1o5
IOSlp/UWWNJXiN95MwMFwL7MxdA3utqc1zaSjado8zqN5DK5GcRs9kWeKhjANL8z
EfBSkK8iQBlAQnbkrrS3mDvC3q8vID7doxFVUKn7lUNMGL3YX6uVnr/gqWqzisDa
db5ttEw/EizFuCzaNTmD+q3lX8vYQyTDzSOd0jFOB8FPqfpoAVBaWZIDlRs1pjCi
I6z4Mxly4HEZub4Oy7Kj7w==
`protect END_PROTECTED
