`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N+sQcE2mUEitrxgY/WO44n3rKuoAEZ9yo6p7MWrZFjgO0ivrRaMeS1PktuT4byU2
Mtm8JJRetQNKMzHQclnRoBtuOCVCVBQry3gJX25IwXqOnl3UmaRDlMrqjXtH5nRH
QGcVkuG4Egbq5iikKZDd9HbfskG48bN4cO6kkRPkPC06DmxvF+xNs9a6bZp/IxL6
K7eGwKMOJhmXOpOpkFn02MJh+A1vzWuax7FOy5CrbO9izGfW9z6I9UWOpqnFKW5I
svJS65yE7f1b6CVJnP1eDkaZ4yiLQcIJ9krkDm2hO5lBfw6fgEMY7wIBCkg9ILoa
w/SgWOprjKx5Ox2KXZmjGcviarmM9Lk/QOcj8dnk5+wWOtjq+kE/EcK1pr76tp8R
wwJR6rx9JEsf+KXYtOkxWTdKwYrUWrRt2Vh7wPngRcBNrxlBYQwQ+umu+pJoeLbk
VvWFqrel7dp4SryAU2OBedhZesV9WLw2teq38HbW0WdSfU8r0xCh6wBkTxCEqezO
xF9/OnN/6VsT5510ap8JKejOWlOynnRFwlqIOzFJhmeLBOvGqll3QEefgZ0nZFts
5HOMxZQxJt6Gq4X89XTXynMbCpzB9OPxA7E3fjcO6D54PUBmjYMpKeQ0du1vOrTd
19ItlhBK5V8SE1BdK+QYaqWHBQBINuziZEqTD1yJH+TNxp0aWnC1MhIhEnUAUpsg
f+p2J+Nz6EoPqB8pZ8y6ug8gVJ8Eup4kbxbqPR36jl6iBxwYLK6FlcUtC/Y8CdLm
iH2+i1nrAjkZKBm3TxUrgo+1cVvB+mRw//rdz/kwm1Ll4BKNSB3Qw4sG47bpoA+o
79EW0plaqKfAtB1dJSbg/ylhsyWuGOIdPkGL7OkWNBCJLxaH60GFWtg2fgHNL+d0
AQ+37LWMAzt1VV4gvpAuygyD2gdL3qi0EEcnrD60wxNlq+uWowAXFpND3cqUE4t9
pH7R/zZf46hcDmBoue7Jyqz84wgPsnVgMKmFpK8YqBPUXYq3E2Vo8b4qmC9McZ3C
XEXs3dL22GBCrIi7hexW5rojbe5W6/8Yi9AUOEZBajINRjMsXBg9SUyLFyPcb96h
FHLjPH7CUwToYVoyFerec5Of1BzG7ytWeTo+tG3+suqKPFPC/8K8oqMHAbs9fRHl
Icecj12HKztAui2Q+92a1ftdfZdtklaL+SyIMAU3vp2u7ai0OKzr5I+hV+EeQcqL
yEKpqc6V7ycLzMNXxokbstRVY5kG+NeNlT686u57zHmkg5BAX0dluxxZ+Yu2yRE0
o9sZ0B/67bsjmjpx1Z4rqoM1Go3msyXQFCpxSayhefw2UVx5UMX+OpaghLIcqYp/
UM4smeEmsdidrp+nArixHaJWvqnSkbgsks3ZNhWU4cOjgG6xfnFu8mqcrOPYM0bp
Eg1EukM+D5RCqqQ7xpYby5tC7NyYMCNTVJ/aq6wJaG2BOai46CGLCYwvMIXUt+dt
GxXevmp5iWZnohJ2nsEbTVIVV0Ir4gxhhIRIKGR+UZRZn4qFWOcQGwasvUIGuWLA
E/izpny3D6Wv8QcKEsEQ+FAhEjO9McDfdztLBM1pL8tNlx/ALNgyplk6IkLUrjhz
thzoXgZ6h2Le0VHASdXmiIIc4tCexpIDoqUt1rOxS+5AinjkSfpoR6R37wV6o2YP
OQGyzPo+70H0FzypQH+5EE0sTXzmlB+iwOVnKZOqy9Yo/5X9jNNtOaqafjoiiDuT
slgMpcXTKvTY9N4/llXDhk6Jf6AV4nZ9TEDzoBzWSKiEn+z9kRiV0KebaDFsYdXB
bxg//7g0YS0kSb7CtVmYT96n6G9WzNzM8AOeqGYEBKaZfyJzma6U5Af8oZiVPCiI
SFFCxgn75rSpTbMNXDVYd6JmaLoBO+8cVWdt2qj48JX1rce4E2DsnFryG+S6h1gu
DjXFE3/9J1nhHVKIl+6pPtxG/VtTrWSVUQGCZGJ5OB/hzEdQ+VCoEgLj+XVG8K1r
NkSI+1KNVM38oILPoiPbmKz5pj6xZ/3/+WxqsRbuGHkFcv5cuSpuwniJlAqr5b1/
9D20gDaSBmSRv4xv58GP7kkaYRAnhxGF2TUNpHmz8D0Yti04fX8Bf6893ry9udOh
ATyjDcDfVUh9MCHWPmC7YVgi2ngkQwYs9rrw7xsSgde3NWjsX1FBr7dpl4PQ9CgH
tTt95QmtMtu/2ygVTibm+q9XhyCNZ7nzM60AgdW0nbjet65DuzrGO9WcXVj/tXyg
zVymx7JiYn9bYs12yqhitpqqTq3pYxKotfSTZdIRfjzqrcRoRHOLNNbGb0qsb4Ql
XY2qLOuxPyI/tSrOrk1aDpXkniuCPHe48+Odx+aWkK5GXaYUUtx2VoGUZfdyELYw
YXvS70Y10nAXUO1MHTDexbaBNu71YnrVWcl74ItnmbkyYLNRfmA9nuU6NZHC+nDU
ZJmQrTPSsRgO+ZG8MhiA4W6aSeYB+RpMkI0t1cPnKuIenKHCujicTE/nCd2ucN6n
lwKgkfkOgRHo4RuScXCAYN9wVacZhPC/QpgPvBCUC4SRjQDrJMQZUQ5lPK7FUKCO
EZP8o1ayv+M8Pyz3VtqjOz2h8tSSOyKGkm4WB0l+2k3WT2+UJmZb0IEo/AJ6Jbbn
OwwBBaJ9gieBRRmoybtlwgblPRie9ygw1DNe6kaIbPIhwPd6ymDdLb/LIOnVkZlQ
XimfVMpJqM8LxEsuU+WbvCDVG5s3InoykRfSguvnkZ4YNJ+uuDZG97C4EtTcQCQV
hr8AxM4d/xlAIw2mYApWWSWZL/a3bUlNgiO7W0/AL3EUnzCJFO2VSzr+wsvugsJ3
UM5/a5YpQb+i4AQF+gN2+sL+ftAaQJiXffbXWfD/XEyOrYj5MhC8OKQYLQ7txdZB
0v5ATBI+/A3ziVxr5Z8RISQ1MEKdymckPEYo18PHfop2EBr4dpQkwItyV+7o5aSm
iEgvdqE5/TlOFKbXF9DJGQzFWzlKsqwdHdQckvhIjorBAJb+aFYrfcx4LAUs/cm5
HUqA8RNvByBWugkolBw3wTJMDcQ5dPe+y8Z2gllGZy9TcWBJ5MAbAAXy48P51E7J
wEsuKVZosj16schwNddqW7BNbYwhFPicDqIbOWqDz3sV8/XC3FaxCUe6rh4PzwuZ
27HdCMdfDJCXGN7af0rNxWDEMOa7r1ZmeRAVvsxzPB4NSuXmDzuLtz97b5wfQMzb
fjNZFZSXhcEWszSv3o+6DRefGlfM0WvzPTEuxIdddc+kadBe6ftm1IJTan2SYtm6
1uygg6zHP6aYk3FmmoOYkTEyypb1gT8Ek+EWwBJwEVmuDdf99irvI3F9ywIYNDkU
SXDw2wce4wZ/nbhBQM7KmPZvFv6wqWFsbBxK59MQvgl2qDT6bKN2RIaSsHJosgFR
gJhJolzV1GzyPJUzEdndJku3zNnIFTmTgceUc603coE0AqxGN8IgstMYdGpzwS88
g+KAjjHz1jvYMdAfpbTCCETMmXNpvetBKn3B4hVRqWAMuovl2xrN+mY526cVgNl1
iktGAb8TVRM0rW/ZQRLLLPbGMLXWhqAX3UPZnMhKtPRiVb7Xh6c3Fy108j2fg/xr
j8LY6pngfv2VpeCmuwTo0w4E+njMRPN8mgpH7XvPfJChiySEPspGHBNUXNhHYYWF
//ZBcK+2XlInHPaXb7vXnhGLQpWzHAiiZqVBnXvI5vMZrltVnHZRz+HYGi+u4Bbj
`protect END_PROTECTED
