`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MSu4/re0xh3APB52H8ucUAtfHu/ipKRGGPoNCpnXzzXCmOOZknAVBiRljD1Zbggd
LXHYXi8KGj6mlh565WF+4FLo+fKt/05Ieo99RI+g73JujY209ziwGeV87VsLyi0H
HcR3dRlby6WNIbAwhzULOEwYGKs6yL2j1uekq1lOHLgSnwuSpqz5ybpSqO82n/YH
qyUjUeH3FRwm/x9rW5iLQb4JY2Ppfk5i56YEWrUj8QAvKdMIovThH5VhtLOtfdZb
mkqrJPGJUZ+iFppeRtED+DHibZLgbKWzAxo8xAPcj42fKbuxl8D0KKC8/VE88Y5i
m0uWlvtM95ihqtVcMjqBanB/XT6ZdKb0qoHu5VHxwrMeks/kvSDTAUsJn1XJurIo
slZX36hSCq5m9n782tJK9gveHU49/jctkkU6bacmYlU=
`protect END_PROTECTED
