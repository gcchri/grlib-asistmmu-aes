`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
91GCNNsPlMsX1tWrW5NCNoPrWDFfJD2gAhTXvnlTIg/LIAHDnfPaPllXYZ3veJm1
x6ZCSQQFNfTxGGhtUiTvsfowUHELQoDoN8B6qCkA5JWkwDmkELhw1gTEVotMif2c
1CqULjTCTPURnDligykUfxKNTHoMua+h/jwCBQ2uWFYxTPqtTVGtBX6zDsCAzWsf
YvZXuQF3Ty1fqIaivjE7Wrxc2g+t2Z/dh9eLlOH0CQ0ckRd1hCMED9L33iOdIKSb
+2aaRfw9tA67QCtR5redwg==
`protect END_PROTECTED
