`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PqYqFuuza2sATlsacIrMsO6vTFWGbP8+axND7VznFrtB/MCXKkg92l61SfOJKwHI
w72vWGSnbA13IEZUICN1C1dBUR/Wqc0L6lQSSsjIxl3GsRsdomPheGcFelwY+xgj
+f76EhebBf7n6RAaep2K00q7HpxghJP5DE+DsHUrPUQCDWeuh8XlLLrZCAvvAYPM
FkKXsyaUA+CJ6b2041xkTdRrh7YCCrnMjQn8PASewF4/e+xbeGSRf0+CS0UqoZqb
E8eqnJELALjoz7LFCAX7CPjaJONoBCxp3E6gJHdg0qmCHjlw/rRAPjkKIi7nXVSt
ZblxwzxJpCrgXQDdiMSFkx4ikY+9lXD+Iapzt0sqcOTTs23h5Qs0iaoSKJUCoYcX
B6aR6w0NfVGjGlLf16szRHWbWBlHDHMluhBJ5/KvTOA=
`protect END_PROTECTED
