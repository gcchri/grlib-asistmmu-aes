`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rtf/ezFOjmi8Dm5jaMg7F/Oo74atrv/o/hDwZDlMl7uSkoRjREW4dVmgTL7Qsv2b
GZTiXU4SD+pOoyBPEnhEGBjrwOEDBP4euZKi/kJ6vUHIzMfiUVw2vQ3nGgdnp5Ib
68KYuLfkRq7RqD8y4QMkkYcX9C7Z5kKSMVTTsW0AC9mkAXcFh4mQahCvRHGK95JR
qA3OmmiE5SXZD0wq3PTYZQ3xbotRL3c/h9ve544Q5h+RLShspsSlYEWhtYWCTKgZ
zxo8yw8FaUW3CsmGM5OC2gFtyyfMlqsAmDfzoWsh1uCtZ7QONnajxK9+SouqwdHr
5Q/tX+tC6Mf11jwT+n0P+eWvjMdAHnHaOKDnufRDPJvgPVe9RiARrdV3I25lJ2Mi
`protect END_PROTECTED
