`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uNRmXL5qEPh7x77G8raR5+mRaru6xoBT2h9goP89CBTJG/OKydQ9EDCohqo7Ep6z
D/IaaalRufLrTp/uCdKLMztS2eaKHvLG/Tb69heYSSkTreR9LPp/lBC1KUTG12uq
wKYAFABUqDQ10gVI835MUqwvOAouBHAloiqbhHbdjeTUznZsYG4iCFLE54T0XpIp
dYIywI3IIBwaLEZIeB6hb3Ggkb7+D7pKjvVbq9jov5+j224NsXzHN2GDj6pPP2P3
fbXuQBasQV68l9uLHzsTViJXissf78T0OngYMaCYLsrHPjwQngEX/B8eY46EqToh
myRGpkITYn/nD05e8B20f5cuK6QBFlNr02E00XT4f0p3bvPiCqsXZgHJvL11eVpv
TAyRZ4iVfjM5q7oGRXI/kTsUzr/WSA0dUyDeIvXO2LxVJwRRjQl1Ox4pH5zR6Ku0
2mv+1jzun/1Xoi0oozuArQgmiSx8bo7Vj9IXNZI0aTNouklB2VWdoToJaZ4n//SX
d0VqDZ++rI3qmYIox/kbUd9oAKDWrvl6mn0WGgHJ+x3FWTLMQWCRMdSM6fwbMF57
opVt5p/GLaOpOtNqTnMrtBIaet9SAgIG3yo9UBXlaSRGiipyFy0KVOwZojPWLZa9
guRVJCPKHP3IfxGkszbG0rfPfAPQte+WYkPC4nQRlNVusy1CvO2wh86HOhKEoOeQ
cQBAPXozdPHBn3u9//4W7/sFCu4U9PlLC9SXzUh6eNCJSaGGy1f3b9GoTcdly06X
Zgedu9IsPyZu5QpMfqeVcrC5UsUtOLfPQ3GvHxwHtR7MXgtWzp0RkkV9jCRXRurw
cN+ZblT67RQu7YRDFs0E1ILn//6mX3IBF2vlCS7pmivQ61/xElo8y5kLV0Y0ka6g
PWr1mB+7EeaksguPh8neYA1G2zwyruQBoRTA7r3TkBYOmKovv+UX3KM5Od7GetbV
tkoWTC6G4Oa7U0RIgkk0l7w+tKUHZx6SNPwNUlwOw3kZ8Eyfe+h7ejF9PIaJiBKL
lmoVfUQUQhDFlUQPz3gR1ub/+B3ek7hSmAa1WN2X2see7sPt8N4f027X5eZuWBkg
BkjzekrIsKTj10UhIOip7H887l/SAbkiESx0orWbB868GwfCffChZrS1R/4vUKyW
qleoU4GC+tHdEuNSZGayDim0mBXSX1/XOrhC4hU2nopmzd3o2slVnCmJq72Zp9+e
vzH3sMdfTGwySJU0AbNNXuyF1mqYtvRc8pNrYt9KhJGqhtxJjNg2Agr/Fg7doDUr
MqH/bfOph0JTrqPihgic8+lV7SgJUSVXWe8i6t8e1gW8jbNIxOqfYYgkLJGVhoKR
S8ydEakZPfUDn9YyCMRbIARfk5x3oG/klMQw/YAtlRtdwMEBshve5nEghJV3TTgN
61i9euPgmcQeur5Mwl6y3g==
`protect END_PROTECTED
