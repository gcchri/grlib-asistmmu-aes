`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
++/AobySZPPI7uapZWOkiR+CDbNagtJoTPJkwb9tpMFXfIK/lCPqT/b9rHCGJ48c
2wuTRKPIgZ3GhZyOp68b56StgqsIEsOGhC6fgrsp7oH5S89wXu2BQntHTNB2bRn/
Mo+pVB3BgriZ/wlddtJE4NmwW5AAFtKpxhbqOZ5DRu/v02qNoUVBGMo3Yx1s1ti5
2e198Lyszp3czSEEiLqP66nyEd1BSRMKZflp6f9Xc9Bh3d7IfLwHERIs56Eaf9br
mVMOlPFPBhhC8xkY+afADFkqfFDlBWP61WMOM1Hg2MmDB3xGr4P3wPkR56AqxMuw
sUkkJH+jR7LmsMrUuDFUoTc9QdNHcDIGMKXg7tQ3VS15crPPuhO7KMBjkbrH27/v
La0+UP+E48NVW5+QnWBIRhz6JsGd3p51JkC2C60zKkw/8dFD4p5DyZJKagiie4P8
8SJOU9A0+QxAsRdLfMTqUOHw7Via2vcFb4ormeepIwi7BOvYisY2F0l7MR7On3G5
`protect END_PROTECTED
