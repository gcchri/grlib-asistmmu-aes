`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5G0+alk9ej85Hep8yi+4H7Z412xfj4RP0vCh5axtJL3QXJ4fQO3ssRHJRIxA/v9G
yxmxoN8Drm7byjlUe2d6TZdzYNFqqA8CYChO7bc5eef/ZRFBqdGsFp/8yyxBFDB5
CImWU73ut1DMIHxU6a/2CNi+V8qHF5JR8UANjOqhYYX7LXEokPghIml0f78dyljH
w8Opi64Nq2sIgnE4Qj8LPH9/TBwhj9nyDYKcn2aftl8V5fhtDT5vY6x3t+wyTl1q
E6Fd0qJm5bDYHeSvupkUWP3CnHWBsL9NFjUHv+BeQ64=
`protect END_PROTECTED
