`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
clC/3YniIwVPdkTOdL7QyB+NkuaucfkG/84fxNKNTdMk0lkMX84Wbx+EkWIpaE3I
6FL0f4i/YTFvR/0fxEdh6OpgwnHCntRBRDQtXu4/jkKFVHnkbGz7O7OCU/N+wq/0
98zcPiSCtxfkv2a52Sjj9bXqmLnTF/prSj0aQ03rIAHTSe9Z0CJg66zkTT0NigXj
51mImzXemgYf7KNME67n4dc6z24HDmFvhkoeOYIuL4u+xkaaBSObYtepn1iqgHsl
sCO6APtRAV+ivJXfQMDk5QPqW3L5yIO1KFZsXWIjzAIBXx0A/vHzyaTq7Hag8evA
vDJeMwpm1gsNgITg1BQ9zy2+3lw6ehT9keugKoZpJzo=
`protect END_PROTECTED
