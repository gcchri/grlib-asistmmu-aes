`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8u0iHV5q81pbZ08uWi8n+LCfPq0unJ3TAbqx6U3wWhrsx2g2lc6h8+qxAKbPi05W
m5rVPnBcMhax5OInv02zoxcA4HQuIZ6l42RWDSpzfFlpc/nfPf1fAmVW0b36kb21
V0IIHNLO0wiZtA3/Mos+VFfcPTXfaGWO1SAhLiAu6KfX69VcGibmcwpwLOPYOMgC
UNBBogTU9CdTlIs5IQ2WwnSwkbZ7mrs8UoSKv24vIkc4UPEYZvZGdFpbMtlWNuQj
eLCQoO+sdmFzLurOZYE+jSzSKmIn18YpoNpcRD70vYsTGATClyziHxKBRCGQEYIL
weMXaMVoEl5KLcbEfrWKdKcaMzqcfVdwq1bE13DRZqIE/Dc1jDOigcBiIPLoMb2m
6Aade5+j0tob9vawdFeqdVnYa6KhBnWUBWmZ+XkeInBR0r+8ZGxnmVm6SjMNvKEY
+NEg8HO9/18aiNVRgSujMmKzMKFCenhnRFpMfs38L9P0GuGTS6cAbRwSeZtMRnz+
TsesKXnbFq7W/PL0YPyo1Th+OmgnCKWpJK8HUotGsiAE0zEFe1d2MIEv/vxto3N8
s1gSs3si2DpUVIhbCgBEa0qFNDcBk0MdKBZ353xbRDUU55MsHIaaT8ObuzRdKTBk
yMpR8h6Y6kxgBJSoyfY7uA00qUPinuwv58+GoziM58qbksz3l4fcXzvCexqwuWxe
20/Q0NHobPvTpw2gtVMhnP4SriZc1c6jJ7oD2wDwqydNgRaSXhRxT2ZkUJtA41ef
meSZAbJ+pikP62MogaTo+tvJBwKSjhwlGhdgVRSCIJxKnIu3YH7KXiDDZwfX6pGv
1SKUsCm8xVMVQyG842v3WLDkVduwvbK62hdHPaRcc9wCeIo7ZkV8fydsDCb+zkoh
s9gBirwlKx7yd5k+f3wBkCo0C5ZbssTwuCr8rkqW9U1tUGDmXaplpB14tLjiuV8z
`protect END_PROTECTED
