`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wsry7oc5GcH5tsHLGDUCwsY7jUzrhZXa9nozyPcueIIjrUdb4yNLzwiz4gm/ABcC
XsHDP6mwNHc5dNGtnfEplnZn3iHtnvsGPLUZ6F5OTAl0JvJVJZd4vBDNLK250MP/
P2z4pUL0mevQ9lua5sAFiQukwwRGSQV9EY7DexYCvk8CROQieqN9yq6xloIYZUEl
qFZupW7NX646qZsCwoj+Xenl6dgO0zqGSunL1xFnY2A+tigv9HwHQxvC2EsLCLcT
uD6MVePSzqXBZHLdbNtUaKJvX1v119nj5jxPAy7GIFOWitlfowf5+lQJ1nznTm4+
LJ0OiwFDYXYXHBEIazJaYkctcgECWSZ7LZRt06qr1thIi4un8SkngVuJmw18/GuJ
XVDZ4ulcgU2KzKHza8aa4NxBkzI2mc0hL8RzZjpSnQSAmoWQvKCU7o8x2SoA4aC+
8P1+GwhXiGJ/hTbVeHBHDeQix3EEQaQfpRDObFEOaKSlzOVkanYnBNxTyeFC3cLM
ZfHPKKnkipT9EJ0KDRIK7KEgCwDxr8g9zNVcai4LrVkC7sm89LGz17Dw2czzxqxI
vtQph8RQij7ZnaFw5/6pK1oYFP1xdEs5GVAta3iNNF2i8OUv+aReR44TTcrhRwXT
+i7TxsEDaSQ6LjmGO9ObnWtgJF7qGTaV0yPzSMP36wCTIH5qk6KvfAhsTtdhHyks
TED43dRXViV4IdMk7cdPU7jsXfUrtBGajI+GyInnBiz2yNSZhWAe0SwHUWiT2xwT
zjv3G42HeGjOxW+P0TKxL1u4OhIHJhkbuhbOugOJQfuqEz26sHZBVwJwNccjiIjI
ddpTfe/3DaAcWc5Td/Iml+IjljW6wSwjRzLfOVal64Yi3YbBqfZ2blV4IUvzAEj1
xCKPvpXNA+2TmpHGIYfaniCX04kwpJPIIli0dHvUyrybPZjwhMxRDmXl49LvO16J
uO5DvK5rK7mDgvF+o5Rr9XWLE6dDCqdMxLHHDJLEXdaoyfAewcCl49YiisN1g5cB
cIfa/86hjTgoJuoSpgIT31G3eCG5V1OWeQdaLp/plM728MCkP6ZpPy0mqLPE8PlU
1599z4bRpq0o9BOTV0d35gRgIJvEYqfO5kNEKIh2HcGjrA9gK9x3YC3ILFnWjtba
WRkk44hB0+RG3q0tX0rB8LVx5jnUnLSNLY24zFVqJ33A29zI9m/XKCQeyMQcVNOG
OQU1VrSvDfcZIMJNpEAvpIs3RrhM8mj0mq0KN9HYg7bt+fTD7NFl8ZaeUv17zadK
1c580Z2JfRAiqOWZWnQce67Wm6IWAsGNNPJ8yMCvOJoJRID/5LyLUlKaC52zBQWF
k76Bs0dRbGWmDbvKZvP14f2ZfMGOfSFyZljqE64C+qJjWi9InzCFQaIF2H9qNwyR
+rKMi/sn2I7/n/tuT6n+cu+ccRde8iYaK3UdVyyb9MmkPQpKztYXJEkQ8EuqYwij
q+F1gDyC8iJMti52gIDNBBUZZ/JM6/r6eCiLIa2HWQ7ilHn1fqJp5U0WbhYxIMdJ
kB/hYQdLR1LlmH5/U5n0W+oN/7dzGiwOZloi2brz8nvcOKbqteSz4NuwFL5o6avK
GCz+TIAA5QR1l85Bma6kttdGqyvl/q1devy5l169ehBbyHdEy8lD8eWMJkroeX2F
K8fB4j52A9tYF2UcsnpUL9MYWklIy4P/PAjpdPmeENxlq03IdHVtqwWyetq29wrE
GJfVYvBC3ye1aMndvv5Sewyvm9qWG6+As2eRnLUBaDX4rEC0kCqjFGZexhnLKq7s
P6NkkYCQrFHEkcBFtYTtMx3AimEaFjgzVdwxUhYPFouZhLlb//U3MnrxVl3wm32k
CP7sMJJ+tcgxVGvABE5lzHewzieTowDny9ij6+HtOM3Gz+GCOrQHtiA8JuLpItDG
oXG9BZuWB1QNXsFGRo+lERWdKJZcjX30kC55NFJjedeYzxisTsZv8a8LzuTBQjKv
MkYLQcdvgoic8LFj5UJOsiS5j1b+BJsm4O1i1CEtVzI/H4rd3xgH4tD9gj11rCF7
Sm1wWxYUdBN94F6in05u0VqGi9iCPAV/WzRSHc3Nuk26s4oMd0Yg0oHKSelE8At5
4+9Xx7kxGlNka5icpJ9MLUsJrAzSbgCjbBndsCrEOtQdGKNDuPL7RZp3Yg/STAX2
7PNWOuZSMXE8horFvNiz7d8jNyzmDhTXOLqV3KlBON7/fXNiRGbrmMDrCAfPZrSc
DEelDE/YDsv4kj3VSEPj/1K5PtwvIdZs1pV475+8hzKsOWsOGotx3OwYF1+mZfYw
soe3NoxMeP8/8JVOBE1YXvp7lcL+2A8HweVawDvsJw8vnQXSJ6cnL6NSMTJdu+wU
KyT3Spv7+DJwRtH7RtJT7dyrguHFNedTxSLhUYJwvpNVD0cE5ygZf2hzNZZMI0FW
PKCxI6cDQY4EdDC5GocilalmSSC8eDQprBw0BsZNm/29vAGq3uvrPKmUPLFTck5p
d/FUq3d9Mp8pckVBLafa4uwzxcqKWGAcC/2433vqk+8UmMMeb2Z1cMG1B+m+nKDa
ZIgMhiFPgENIoKr3LEhN2IB2pFIRflCVo/xIkNghEJ7xxTjany+NE+BBxZkFZvFH
`protect END_PROTECTED
