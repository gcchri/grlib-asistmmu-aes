`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UFG+8LJduX5bBAT5wt7Q7M/kAgopfayJihvsvyG/t6PBnEJTUYjuC6SyY8svuc6R
/TsyHen18qSVan/ePNEPyD1Up1RQPKLMPhLalgnbsJd29udefp4icVN+V+nueBEK
MJ3G9cuI9ibzGFrXANIoi3HNuSHX+BdPKhuYXn6vR9nunYVjna/HVtigU4JwI9n/
wV8FOQdGP7LlThiasnYefaTSBbWsBpPJwCGRkVi/2EF9xy8djFjjAX1Am4zlzqiV
LH2SSRwxgR7TJAsQ4VaHgk7m5Q4I82TENMCiAnCcNNud1E4M3xeK9LN+LTU2z9sW
9WLVk2gsWZuSnBXfBFn2XvhJ6sckGaTlfWoXyrIpTaBarrvjnSwWvQiESuLUDixZ
w/irOASn1J6gqDBg1FJJPea2H3bkya/rJdpZV83ZkRYbXSnp7vgTXYuz+/eBFCQp
/bImzyknjTjFye8MKLTFc1yc/2awUvD4aHps9+wxYizSmyYya4jeaf6JOgWsC1au
LsaLhHtX7+y8sySw0oVt4AA/ju1RJG5S2lFXfJ5DlWj14/MbXM9lR/FlH2cANIFt
4vAEVYSTVFfJE1M0IuuYP9S0wfUGQo+FzE39b7J4Stnd24IMzMZixFyfVudkS6lD
wX66jEF+mhoNZRKxCYbX0tm90ALfjkUTyj6O97UdK1G+3aa+UaYLo7T2DzIF3XTv
Tuw7k8WjhLAGBBqKtGIVRsIEp4Tg4Dz4RqMEecnspzsrzDjD3gWW5D/KUo8L0nkQ
J8qAATnZDbjfCunZw+q+gGRRuUsZGCsSosypTriEByvszpcevoVR4U+oOoJ77wSl
0GUT33lyGSqeVdxnkS27EzweMUcRHioL4IlorkVdWIN9WDv21LW6664yjMsZk5cu
u+tosxkBqmMccNyHqOzvyPZmvIA/EkkvUyktnnTF9MzejFw2rV94j1zSdxd47AHL
YccysQC2fq+viC3a35I1Yv9YmG4kOnxv11KignWdyG6KvLORUR9TmoIqARSfnma4
EhjxnNpEftqobDg/P/6HyypBFSLCkk1ko+QS+/CRX6QBKNPSHbj8WJgM4g2m0YaG
YNgE0+MIbEJVvx1BrtuVEPxMjs+St+ML1dH7jFl2l5nj19dUw0QXn6hrKUFtYcJj
9uc878bQ9yW//bJhcIDV74ag6zYrhMld+X2u6qJ3FKlvxYtd8UTVkig2EUvmldsM
cylFXMOUB0YSq8TAejjTzIz5jEBT2A3petUKzfptSESkVkAYSzSYR5XEoxOh5zyU
C+hjbF+Sb/8Co9kEDgL5ZRKeioeDKrBLLkEtLDZhVJL1PyrW76wA33un7gmLqVN8
t+xu2WtWLce/2VWY8QJdn/+O8bSo0S2HoF1kAXUlUCSyiPyu9vkyWv72tDgrjAha
wdto7nkiFuX/Es97bChCrBvAOwQ8cBDlWzZzQr19rs90bWHSXYbF1d1msgrSz1KF
Q9SOT0+AiRI227U3E0DbDsNYjIha1yHxC2fg6EGW+6eL52s8lHP79MyJiwkYBPcP
OALy1O4FZ/OYaToZnQ/VKuFE6MxzDQJBxSxeZ7zaSHHo4ZAQUTole5fFuHJob1sz
aYpEfl2CdfiheOXyk4XcVfj+zOMuoHCPebCFEkEQ0naHHV9B5h+nY0COhtFKeBp9
dgkS1OEo913/l7SyP06jJRW2janskX8pcdChApM3kBNbcb4jArup6vN7Szj1Krqw
HmQK73rVO36fnVMU79F8U1/66sws3gsknSW5KrI95Z6+9qWafL5Z8SYeZaY94P+8
H/+nZAgIlaeYAOH3tfndKDrcLGSoys/qBZb8ECooM6bve3X1TYWl1KqRanflXu5Y
XUgEfGsFHQeKEymFK+n2tMlpB+fhquStvS5sll07jDyRxAFzmV0G4jRaKrzWcdHb
Jk4XEs2bUsRHYix/jr7/MILpv35UMdrW2XwAOCpTCFqd6yCQ75mi+bR7lCu3tKRh
0GQF7SHWr22Ycy3yEyeDMePFE9nXkK3ds0ncWWM1D5uyvZ+TzgWZOtA/ooC4tV1R
`protect END_PROTECTED
