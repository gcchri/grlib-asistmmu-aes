`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tkY8yCFq981FT4oAenFcJDkT6jcsyZH6gThKK9uiXIqafJCKHaZYR87rOQRSpMqe
mDMsbkx+q1ADQe4eT5ipNwbJ23iCD9Iy8QYVaSGuyVFsU8oZ0xUr2pbd69aV16ai
EEZiSmcJMfpuTWo+7O0wo1kIIkfpi0m31ERfizmZWDUcOA2AT19koFGFpDXmCZii
L8hXEDjrc0rdA5A1G/OmFa4RJgL13rH1XvZ4Jo0YFB5108XiCIMUM0GGRTQ5urVS
ZTKJA7qS+LiHLCNo9dy4pnu8ICiJM02mWawjdA9k4d0fkpv9Mrp7ZHGnVux0Bfcz
Dkgpwvwvmrl33FVJNtGOcWwYUHY/+jreO+Pq4vKPVwj8tkkHY4gj36MD9qTBonJk
BsCbRrFNPvZ7GF/F7r4mOWbY/67C3svmsLp9FrSZbwX1yax7S/AuxYkTWrNVZ7ZS
BFCsFeIHBsYbNcdcgjGvXrwT/mlGH41DdNVYfonqBWTqwIFTEK9BD+uUHkJ+y7Lo
`protect END_PROTECTED
