`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yBWLNIOdUU9hraho3EXX/JJZYlpR8UhfERmX1n0Lq7NOPJQkEPNHuHS0e68phWDo
Q5ixbBACRZc/sqhaT5kNu3V5NaY1wZnhtQbeVJzbuek9T20dZVap76m8/lDvsUIt
ox1D37f7yp8J55zKqJ9rqLfrOonmPKLB3u1TzPuRzXCfsr+26bDjxXom8Sfba4vf
kWppsO7bAKa9qItoVfxMAGQ1iMl8XQnNBEVsb1hKGZbJJCRsHn1EgLURLIB7Ep9g
tvieIZxWoqwbIQM9W3Z2Bg==
`protect END_PROTECTED
