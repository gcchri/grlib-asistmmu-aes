`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oDPV0a9qGyPmCK82+muvruqfd+j1uFkDd4WdVcmoWT5kHT1oR7aI14ygVYx8pB9f
18g1WpknYBVPhouaybNY94gaJlBS2rBiLfr2J3phCmt818xJMFJQwHUskMwQhzKf
OlzrD/vVBFpazmAlbAm4qDcTASCtUKiG+w88lwPvSfae+WF3mdBZYU2ZSBTENXZV
Tukd0ce5Jp6xYPCR78/nrrlRJw1AKswNCbYqWDhYDc+JXYsKHdrI6CPSBX2N5hyE
FAP/Q2PBzYPrp2IGKJi7ibAy1fHcPqjaaGLyOsYVBLKYB4ei3b7Skxgt0a+8omjd
Zy657+HZW8M5SsYnDIUu6bedQ3Y/tpdifKthKq6rsu+befYqNtxPb6MaDh8PFJRi
bMQdePBVijsPaxbOUbItkIpB2PDNO8kEwxMzghiYo9f8p10aMMw4BYCGbdWjANWy
putLv1PTElN76eFGpNWFcQ4lRAX6j2aXQUaFHwEM5hIkET1ni9jMvA7ydv874QLc
f7gKLzcsgWzM2iMdaVxz3XfAsp0Y/j51BFfI4XP1yntY2UmcXXlItMaWl9QEHoJx
pCQn+l6/5I3SVANYD5pG5cBh+02lqdxoJOdH3wPs3LFH9NQSAQnIcmiQji5V7MVw
TOC60dOV/idxZIoDx/QGtXjvJFH8+z31xV2YYrqya7ublT6zla1xGJpy1i2QsaKw
FDfgU14bH50NRydwOW8LszPjWzGXjFTCIi8H0Fc1tXmtdjldZnPc3DMYyJ24/eSu
usbNrXcttMdwGLnvYLpFhXxd+EkXNRatXTjJs4NB3kCu3+nSnKryaI1p8XTtqgPr
Kzie4dkDo3sb2/AVHyvlj1Qj6bOgt5ELbD9mnnaULZJn37refgQk7cS+10nTdUd1
cNlZyvfS7f+FUWDxFj0WHZfHAGevq3FPaG3oAGhRA5qsKXa5fusitJ8bG3wFtBRh
yVhh7w8H2TIa0ToCxMvFoafmk8V9b6Z5acianL19ebbB/HUJ0ofOfZEhw+ZIUV9f
Ocdt8Yw8nqZZ90Iw7F/aRUFlW5fnA98+8zqK6EznpPPacap0PSf7pDwkI9drz+7t
Vh9mOCBkufcHNlTD6w7Qucxybv8HQcq8d6k84w+v4kwjVBu8Hoqv4vzabKaNNHSS
+7hbyT9+9ThEtf44t80KmiwCDj2TK/qnAVHop45rVjpU7C4wvKrkIZgB7Rg/mmb/
deJDulYICVbs2VmnTpvxJiW5W93puBpCGFSQsHTArD6rQJim/SR7esQ/RQkGwZ1+
k+471xwS/0VrTxIwGaoFr5Xtm0NPUohoGSPWGHrj9p4PMOKTPTydGYc5dEaq/eDj
J4fESBStferfafkjOJ3zJ0PQeVtll4bGPNm9RbfSjZqdlUqEoC9+LyWbcok5sCu3
ZqkPBIvHsCXCD/ngvedaiB+ZTVPRGudgapHxfOT5lGSLWp75j05oCLb2+9k3V0gL
alVaVxC+BBpQxG2oPA1GN8r/916Zec4F0DGvZDHtg30AjbN+iXouGp+V7w/C9NRN
Q6njoqtFuP0+sv8yG1d0clLEIie+8YJpDoMimtp5US7547PKlHJpY5JtEut6XZlA
Vr7DdwLs1HlMcQz5ZiA8hh+bGmLkeh3EyIT4ZK7dGzCfHxxsfAZgab9U6jylWC4k
bQBSJGKRg9PI6h5wdJ6ceh3VeZwx0B8zDClUp6UN5evAw/qbDrjDZxL9/9ai9RBi
Jmxgyon5IlD0X8ngfXYKZFw4Fcf6CyZmrmmAoEs9Mc6ztu/GTImzn/inFPIC0HLV
wrJBqvppJlm2mpNI+YMvHCcKUpPyPETOAF9i5H52zYgJYR0VvGpOYSVCf2M9olLQ
6yTwF48czSh0FMXNbs90TTnd3zMrOeWh21KUupvuJxu4kZKXmj7E3QtWpHS2Sj21
MlvsoSy0hSD8GuhVAAl+9klIVrWgGJF6vKPH5DM9kkm6deV4+tL4+fSvbZPlFDDc
UH/t8a5aYrF9tgo0nPCh0epN6BJYYHdl8YlSZwgLhG44Rl/pOp1qumaIfnnT9VIG
v0qaBigcXXvFDS+bVDPPvlMqHzJNPj4y+ODOUit1263XyI7VJL+5rE2mtVdjItpx
gxXsSXf5oP+x/l3h+IjyYlHIAhG1uMAbvWsfPOI+zaN0A49KnAvyPJIa0UQ/dHL5
T4P43axNOgwKXQbEDbReYkf8NjzSF+g4coVoDPFAj30VaukQhbibdZkJHzGIq+/u
WgxxqMQRVtPV/SU+H3o4AQ2+nJoScZoHnc7KUfjEpaUP/bGXJUgAsgHN0BQhjFQr
/tZe/Oa/oh+8ZINyWYBgkdrphBDuugA/rNUfgEKFhaido20Ld0LNxLUN6Ne0Ksi3
5H0a327X9fRNeTNGmfNrA4QMHSxdyNZgsvjcVgzokSWaEuueXPK6KMnX8w2+YhU6
F3Eyd1wKA38GcOEqINT+ZuChY2+Ag4m+VBUleWHw9Hks3LMVCY3kUxNJpdtIl9EQ
z6jAgKsmJtsWSCGCsGNQPlkmh8zyV9Mm1sBjv34+lGvkLqiRgVL+Chkq+J4o+syu
p3RnJBQV2afPqLUC26OBHpPFaWOHqDvADUJU25dwoqnxF5GULtky1rO7ja9KlXZX
KzGnyX+oimo3mOo5M9d5NY0h8A0ai769Zf19IaNgf65skZeBP79fDS+tAOvJiUlZ
d64VR2nUpj04vAa1CdqcjfwUF0WlWrFgBW6U3vuAk/KtPX2LvP9TL4LW2FY0R9VQ
gKi5d7ZJgcr7qYHduPPMkiKKZuJDGnRVyFg+IIqyHfWbJ2r3UJhkhOfAy6iiEsfo
g+R/1r9ijVsnHgpDpwP7yTuesHD6Gcn3afquTWVfW7tI5T7tesiggTBujhg6hTRV
HbihCmfK77k70uH5epI8Z82dRKdAj0yL/gmPwgnyFfE2SHunT0/x1N1GCqBSBPrW
5zBCc2mESRxNU2ZHzOZ54Pgq/ZTX9HwNjfHalBFEYEp6GqInuSRokekBJGWp9uNW
+Epyfr6H4RLJQczq2n41O9JsGzW14RYaDzglriph/zXaA+G3i4Ch28UwH/Mmcdq5
JxuyETCO96HczvNlYZtsTFVeBBWhjkZpHaamRjqSZmPL6+jfeHPcUh+qYUw2+8aN
UoeNfaHPeoS4QTsrufu+1YAJLjV8VR0aqcF3rU8oCAT/+irjNuvAzDfnLAnC2zeE
QBmef2fi5wyoUvVwSgg0g5IYBXOGTnl2IdJqsW/w5Hw282MDoPdclu/FefGFcWh+
GowdjTBDpTUqtFaDeV9pGNItoYKkINjNTYn9YxL/xkte+ZAA24wJo+l+IKkXchUr
DxW+7NEu4C+YFXYDVMbDZIWS5mIJwkXGXsWpdiMs33xGP73VaHbX30Rf4z5XFX7l
AKTUnEB/blBdD0/a+GeuvD6ltDWPFHRJCiVCWsmW1cnD+u/MGWLEjWxwTZAuN5Y6
PJ+KwLcj5XHVesImvtqYK2QeCYHvI3fxTYhQGV1zc9lXgwCxwv6wLtDacCR4QdML
pV05oVtT3nYm7iGJoB3pVuFqPAOxEsN6Zng834F7DlpyvUsAJw46zc0UT3PwQoPk
2CRascXmTOgLzPURZMGrd+7/DtKP0gg8oLGAWLWnSA0qRpe8HZeCpc82KrDDTZBn
GejcpmDlUssHHKjYuWIBDYJ2iOKlI1HB3uy2GM/gRYv2uFZjAmOhaqy9roww/909
2oRuV0+xRJAGhcF7Q9pyg+PHqavDaAGLlnaTZGb+R8PUx5eXJwyzTFZmDVAAVdFn
0qynvDE+H5xvHPtKVEwda4FV/GZt1wVeJCF0UN87ZMu3Qij26g+Whx6d5s1N6sGC
oc81DaTJYsYW0TF8lkTrqkzlrI7i2/gaC4vdhrtFWnQsN/dGMoO5EX2GN2wq8kgh
xS110rqhdyeUJ/x2rIgk6wPEdWinys9WM2xcCppdMmfRTmYXGO06/n3Q3B86ukw/
ZMBcOEg5Cdhwuv6NMwI11J72WvBsDf0DTJSQTCmZRMbMnHo+6yNLA21e5yn2sn4K
qM728rsbwXYKqcuxGAUWbnma1/LlV0/9TfK5Spx8vt+B1I5lZbHZhNiA/CiovQ65
1986rG/vpu+0+7T7HWJTnoFaQNfCvbCvhXdjgx5/hL7MqdmMz9oCeCOJerb1tJb4
szRpmZC7csiUnCMJqIZAsou7OLR0O78KuzSlgt26KrAjTgHUj0k+qFUdom3oIs9J
3lXMRv7GyimkfnbLU3vpoAfB1hNtMNLbhha+crs/eLMq6hYEvH9BWwQWoVZ9mzDa
wwBEPeneSlRBeprsRWPyUkPfXVaqUSsnqQIa1oQqnliYRGv2JH4WPKH9z4QinZzc
nZhORLHbwXy3EwvI5Ti6341Tl1frm9usEmWb6vZEeQzinqTRwKvmfvuvXx3K+2DZ
sV/KKnIHuEnmARHc4vpSuykVnGf0WMi14ekSAGO9Yc085aocYGgkdARPIZDARCVH
CZZtYvpauz1Dg4C4/74GlsFx1PJrqAnEzb+x0CJuf36EnNe28zzQv5AkwS17/QkO
H5o+6BhfN213mIp8rnr/qAuK0VIN3HBmv7MbYJ1om7m50tXK01dpBDrL8dN/Iq0z
CiycosL6CRnI6UMGww4a/3x0nazKp2kEe2ufOKz5NLkvrA1R1jiha1XfKcA0nRaz
xsRLIHV2yYaEe8FOpSIlb/TSpb9exhypVpTuquE5KYi0B+89XkUyhVM7bvgRSXnk
6NzhvRmWCobuhJFbaMtvra4eCTIRtCw3l5Lvy10uF6RCwKQbdOVUxo2qGDvsSTlX
5/aFDA6etZgkS8BUnh1NUARKHnbXif0zbHQYClu05Oo7a5NcJD0lbNn1bghtGDLh
2MgoGEcBtk/Oy+hSuli3wujwm+R5gU3KRtYQeAWgqjUgmSJFE54Y4R/wrX16TL3F
ysphF3FlZJ2wuN5ufKCI+m/p3+z5gWF4eeQyfw4l0J5vcKcPlXJlxLiu3FLqLnmp
f5v1sYw5OsViQyZsvkeJqvqDevWPWLjlMif07K9qxekjRO7mXUR8fMz2r7BFgoxd
D6YtOPOV0pMtkh9tK3sPZtQ6hc2tdSRHSKwtdQhauYsvNyFLCvLb9ZAIdmo0f4nW
NCNnE87XcsRt8suXTfrCix64MGWQjxFq0AKCxWumvEacueUviSnJb9HpXcIX+kHO
29IIdjBcn6oKIbNGCplipciip9dGG2VwgUTstHrLhL8f566zX7adoW7/Rza7Q6kO
6RpaA1d5jlWNSFFaxVDkhA==
`protect END_PROTECTED
