`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iq4EjmHZaZt/tGCu1Km8YQLVybpIh35zlz86WNPcl0XeMBAo+ZNBHdMyjhd5g1OZ
eTLmDbxj02hupZDrOEuoZxzkNE7NDbDeGgzhNBnYsoGi4661uGBQ0NT2aHgvD0QG
EkYnMJocKgaUvF6iVfnRU1ZaTbcbCRYPasLFcvCjq9uW/axlyzmgImdpgQYSVSg0
e/Kh18ocwd+6IGvrzpKl/dE8iUvPw7bD86csXyqFMLolFlcvY+FRIHgxewDPDJsm
LBZUUlnsFZZjUBWZQTu8L+3mStIbR6BYNcX2v0oJEyVFDvLO7coCkGtdoC9+tfic
Hytva0P0NkFpnWglhIhYC/ZoIwwQzZG6c6E6xKjpi6CqfNWkFPjcicnvx002lFZG
0xQkqUw5tWg5RynN/7LKVS/URqh13cEgW2QPZTpKfjvYeFcWw60l/cZ/mQb34Uzy
Xp7g37WxtYIx5tXz9HNp/H26fS9kuAHsJLBAWb8VlGBTQCEv55rRxjJ1RDmMaFTA
`protect END_PROTECTED
