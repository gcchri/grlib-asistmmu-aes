`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GZe4SQI7chrO0ad/0RGpBu5YjjcW/5evZQEzeF4hDY1Vo6IFpROULHige5uL3kx3
nq6YcEA5TjveCmZjQP+Z6iXs5SUw/RpdSlj/PO0gecX941yAceAbxn7kUGeBaw5t
eclceXbO+BMdOfojLt7pmrFJQEB4Oo2Mzfnx8g22V7gOhlShkO6SPWDvCVTRP8i6
QHsG52kBzX7w6byaU/NzAg==
`protect END_PROTECTED
