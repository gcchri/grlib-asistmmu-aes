`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yTnvvm/XmnUBeqvvTEvxpqUeoVQnzCM0YXWeaBqAIeu1Ih0/vJpIIC6xMS60J05b
iwgffznLvot15R5tSDf3QiAye81lnddLCJgam3Atm4GxPeDiRNjD3NObyXSUIyT+
J2NH8yseOgjuOKcpXKxZ/dE360mMICh0shqnBw4WBTT6IumbPRP1tJTJUMOolWr9
XwK4QbLAoamgzb8cErXDC5lZga1D8qw9PsCph6r84bK5D5Yrted7IqPZWNv/Ot7s
3T0207kEHAv7wURP+0kZW4sQczTo/TC4bKdI2ssW4vuuVkVX/H+JWgPWqrT9HZKv
zm1uen05r/V4YPG3FqjAfxHkFgViNeInBEQsPB12O+cm3gN8SHtzVMiMcASSYIL1
MS+XFbZlrYpWRnwxo9VZppFHs8CNb/nctuw9sO8AJeXs8U2IqfpOqFZGFr465xZa
`protect END_PROTECTED
