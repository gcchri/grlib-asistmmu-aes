`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cw574BxzQBsARzywawhTsL18TjGdxpJJIijBx3FSxLw9kCQZetXe0OWQiuPxz5b+
9vujxvvrFejPDPHG3UANOFVVEGZDwGuvwe2ML2trTtvfXLVJ4l/aLjg5vgORDcJi
djkhuwz9A5k6Go3GwVl0uoal+MQHJ5qQ03TObJTp15jseMtDkQBItDEGqUc4WR/E
NAaNAyq4db6EyoSoYWY5mQ2XvAresFIyvO414r1ag5F1M5znkUybPv0jbPLqekdD
ZJUK/Gq/K3jew04Y/K2lBDc11J++BWmHN/FbTEN8sLzAnbD5rAcG1zUnAhvWmWK+
QQXicMP1C0+atsZC1QTGNr4TKZ856RSMVz/8tV0yiLkWP5y3IJnGymlFz2xcXqKN
REXFPHlUgm38+b/h0mkWdbEl/nsV8ROMeLqfUJ9gBnMtOfwFZLJtFB2u/c0sFdZk
4MFbXjU8Je+mazk6iGERxl3BLJSS1slu/CHbzyaAPa8MdMffaMEsB40G2+Tyg4HI
9jM2Fc525o/usPkV3IJSAwl6LuBMk3+nXbjyjxKG0x724VzZUHJH4sfIJ8PCPB6E
1/TbMhDqhRyyJ/HJN5bdS1NPOtc5fb6IKGS3Qr0wgRwV2boQzg6m9Dxa1kb6SwpT
CBac5S5lZh1s4el4fTTTQMp9g953V1P6HYbGr4G4FUxwvRYaOcshHH5szbyTT61L
wtbQhfZS5vKW3qBMaGI6tLccliKhx25An07xub8T3s1bfvq1hwTQGPbmfsiRk9Ze
uhss/JWi8C3iBaWSCnoQHlQq9ru32Ov3c1ZzAySvXA5Ayj0bfbQJVjyhhi5aSQiE
ShC29AhKP97uzxUE0hbN1W+rqSpkeaREJp8BUp0A+V5RLQIGh06Q5gPJoldWNTtw
CCJHmQ0M6h5qXDGhScCl7JWsvOMcvINVjt+zC23TGUYPPdqArrfdwikeDnrB9HYv
Id6Ngj7+mpPdCccygfyjuPjRrYW+qmi2yeitra1nKp/K8n3Duk3MLLyzKOmDLvMU
sNBNnKD86HWg6WreNnbORIaLoMxNxH44LmfLpE6rkPGlk+HVR3ElfjhZDSv0vKnu
lUMWUbaRsMELliJUFmqqlLNbXam0aDlO1vKJmcQkj3SZ6K7oBA/N5WpZ2msx4IZN
ghDJ8/3fl73sHVoblTMrC7T6FRt2crvMP56B6A5P33G+PfpEvoNIL0cPL+rEk3Nn
A9KIL55UcfbICbkii92Eeg==
`protect END_PROTECTED
