`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EFp2eZQv8HtpNNSmO3hoG2YDRWlE7Aasa6VvuPEbQzIWViVhd8MLjwkxX7AuxTVG
bKNPfrbQopsNi68BYPqc+DjkN1Wfv7TwWbKWZ2m/ho/hDcx+FgC8vOie46FzcqBi
bnCsLShUH002k8wNgSTYb2Kp/PCCU7oM1zGSBtPdcqiQI2ypwXZnexmyageS6+1M
cijTe7hZ8OkG8Jd/Oy0+szHe81fbXQZWSvi2JIfORbeVALLrko06DhVyvs/CsiQI
jlv5mql99FuZYVTIMPXUaFS4suw7+zIjTIEtlHmKfVmib8fwJtUCU1LiIRJ5LV8g
2biit4weFwv1ZWVWEJGpzvW1i7Guy7JbijfbMsfbYEHgWCTCNNrpVaqpOEj/XZX3
yOVxLLPbCl1Kzz9SdBET+GRB23bnf5jrF3dg5niwK7YR2Nk3jxDZLG+2uUbtzZ+Q
qdL6B32CcJKomvGZLwODzrntpqKcwSKDe/5+ozBwTp454gfvN33B2XAEUU6VLpPh
WviHd3B7T0arUk/1sIqdSB9Zasr0ieB78LIl7n9xjYx7l+GseI1XwxKk+QGsKBNq
10XVrMSQddkmaoBkXnIZMRVqxyKxqcqvfHvQT6jNNpsA8ZAY7oGM46t85PCcTidD
rScWy3rHLCcSgua81LYdBrpYlq3vR2Jm4U7e9FSIHkU12ZQtFRkC1ehU0mRW7MAF
2HhXnuyxAMnRdQhc6u+PzX/dBIkrpnuXsh34LVvJBV0pNymYhy0I6JvgTmYbYCNF
UP6KQVSJ8MzxewLDlm4LaYMWxhjbGiCqUQdkEhCvBW1XDRfuFGya6m9bYAZvhdtk
0P0mMDSrv2ozsAALSOMrmjALhiI/SLG2BInLN836Zgs+8WHL6LRfF7iLpUnL4X6R
s9nhJJgN1ncbjjMA3Cw/b5X8Z3VK4vPkIdkCGThPZnT5X0I1zOblKV5iqPpPbD85
`protect END_PROTECTED
