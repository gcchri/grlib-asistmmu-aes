`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gkj2onh/tOcRWTAdC0ebeAirYf5Yy8aJIMeHwr6c+akHQHiQczHyztedgV4/3UaR
4IW77/8q7oHGDOQ74la0zvlLBB3VlnRcBeYDNLuCEki/TICpUxSJSuHtb+Xj8DBE
kbtexz9h83/LRaJuZysPIGCORRxhRkzNz8TQ7aPG83B/pfMwD7Qh+jbct0HB8iT3
CKMDWYf19xVPNRHXO4iBfNLBwk4FbJKDS/k9j94sU/lrg2X9VMjOUnKqd0ky31eN
TK6MEqcchgOPnxURFIo4ueep4gv9L7Whx+rDwTBf+96R1CPG2MQQJADKhZfXmKtc
dppCfQca/byZ2MuTkpiNNWSQRhDfn3SG/tTmOmvUyZEN+e8EzRCom8ByWKv0V8T2
f2pmTBLFAnlFhxeA87Q99muRR4KnMGFnt/U03AliYhab7Pe7q/LeTBoyLyxFBdqR
EnPrWnMfDlSyK9/pi2UC1KJPl/Uynj1IE7W2zfNdI/dbq5EK5OD0AJvwEGQdbjU9
CcW1I7+5O+e9zpCeIOaWI0Hj7wSU/7wu6WrMdIdZN7cU45effzBCInadjBn1f0+V
DfFCo3eKgQS62FDoRelVJZUtqbJ2npIoxpf46L8q7gafcG13It1O8WrntVQTUqPY
35XUKNxE4FC+i/C7zKPNXcXJGdZAY0udo5syBDSAhIS8GE3XmoCXMorSVEUMvOQz
cOiiW6bx+VkM4zB4vWSHGzleLEszJ/3hrmj4vniH753KVQC8XNdnOsixsMlvoBws
xB2QbRJ2fZQ/MZg7QFwYvYrJu7ABc5+mXLzSJvozjmo=
`protect END_PROTECTED
