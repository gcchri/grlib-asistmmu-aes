`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YTToTS8WOIPO+tPPittuqhg/yn5chFGc5Cj9EUMVsI1kp73Tmt6k+pZbePz3FGuk
Iz/fNQoopagRXdV9QUlhkyRGHzreduNcdbAcsXy0id7YxeqOG7QpU5VFhTe1mRAV
fzvl7Etr0cb5fm7VONGtTcgGXBGwJuQRBEJAS4q7ucs9CD6Zq40Bu2xo6dSOMftl
FfVbV9qbbqd3ScUrOE2wch16swkeO3vqFoTekTWGoaYFYmpkvpOnZ8gC2zc7lWUA
hiWf+GtiTJc5OyE/IB/wpt2f3rSxJX1V7pKpvG95SyZ83ykEwnnN3geqRfHOZTpX
E0BTMe9KyNfKxsEryPZRe+DmegsczZ05EbKZ2IG4gAViMNKYfzyL0pDe8Dg3OLSw
hUki0goyp1kOabwebzNzLE/9Iik1kcdM4d5zTllTdrwqwmkHCjHEZdAHSGpUw2j1
3NChDHOB8bqGholgjtPiuLw/cNr9vBm+wUQQEzz50b6h7jKl2CUIcUwRhjn2hvPK
V/fO72dVWXTakqj5ys0md/UGOoTtFvLCyEp+WgRuRMBfyGS4F0rWw/Tg6qwxJQQW
zSlyjU41YXzvKJfanksAJw==
`protect END_PROTECTED
