`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nco2IaZRzMuXFzfBephy46uejE27Ge639EPYOXR0BgxbQIC6ZCQBIo0Xz5Ovkcg+
7xt1j6ifItpB+fdyNRf6lCOHrZQCeIFIHP8PjEGvpvUIlfoQ61EShybhfA3NoEZ+
dSSyhisf0NDD8lZ1PguTkWtd4m31hqFt706C7METrNw25JIbMWTawZNUBZwH8zcV
w9Gb+aLeXgu1p5jP2sWOar3h+MuJmivWzYGrA5f7CudpIT89oRBAaHh2uzMwac6r
8MLE8Du9WYUiM478pBE+EimyGX+M1p1lSjw4uZdimnx9Q8DVjlzgbkVbozVfBktj
Uxh8kn9+LB+JgzYv+7r2J2W6ZNYETaGYp3FR7zsU3lrWvBjgUdg9dHkVJkCAW7vE
ZqV5yuW2bWIue6ZdQ1gTnU5yO91AE5QRHCMrq6EMzELwDRIDwWCkGZ5/3uQA4rTj
CJx+VLW2SZGkrRf4ASqNa0/AY74A4ezaSes7K0Y9joO2ao2gdL+VYEgN2kVT9JmW
n+j9NxdObkSlqewBrG245mmSdoea0xa1OEREuguNAdV9HKGSyRd4TW9aQsljXn/U
mN3K/COHTNHlBCxdkgQYNNyiQieb7LT2rRNQIanBHIA=
`protect END_PROTECTED
