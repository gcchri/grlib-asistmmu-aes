`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FKYTKwueq1bBGcT7iIR+wn2Wk3nrQO6eUPmULjz7vEErHYfnKt9MOHnbV5xxC8Or
w4VWayjlc8yG1HF3dJcpARQe2qkwqVvbQMj+g49vSnZ2vH28o0LdAYKttjPvKjbB
yNO6cWWS9nTylWhrBfgieDX1HJUDmHuvqJh39h+J/Rul3yGvUS5BZ94JfKkkkQNl
9jCXnyod1uICSoncwnwnDPPvi5+T2xvaRRDn1WuAz0WbxOJwksPh8nHp4MzHBVr4
EmJWqJCPJYXPRlbHopWcpUys6MaXJ6cck4QdfPxH3yjmFk7EntkzZbfpQRPwhr52
WXpxcnu/MWG5zIFzjcqLIFwdaoOvYudplryhwusdaSWwkWPxvhSXRAZtf2h9c54J
EE057ZbNzNmfjWiTx0MXTMnQz7DG/0OoVLJGaw/Knd/AOEcKkEr32MvvWu8xf2rf
`protect END_PROTECTED
