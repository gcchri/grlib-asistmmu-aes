`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hTRlhsZ4NKB34pB0WvAzMLF64/YdupxOcrcE4x+xgNBPM4If9ZafAIQV3z4VFl3E
yhUj8m/bz/Kq9UzAPb9K1gE65YLKEAqVep6+te0bnnZ21Aelis6/PaczuhgvUlGT
CjOF7g4fGaM98nRl0I8qFuNQjyyQ4DjJWPDwcIwBVAMbd7mrvGPr/Y/8PZRCEiIM
hA/7ifZLTPY3gHjBCttVc9b8u2KOlLlLgI2NThLDHuXxSEoFkKhN0COKunB6jmR3
7an12053tfZEg5fFIGQxRQ==
`protect END_PROTECTED
