`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x8bRHnb1mOMBNk4HQurypv9CGqNI7Z0Qxw0SPw1r3thdA12Ky7fzYCi+d3yCnEKX
696fF6ZeXbAmgydBGCtukCCf3oX1yQ/2kEtXiVJEv7gSeIRckZZEGb2PYCNDY9tt
n85S/h5zhWfWLXg4y57F/ecFxFp7JuzHJdckX4Ybe/Lb9bFwBuzrpJFkGiHmbNzY
agEOydDXR/Usrm2tev9BshLzUXnE3ZRsmI9RtIVqa1nd9fXAE+GE55z30Ayp+Ooy
6/QYehfIr3BTVumN/edjS29bAO8YxkuxFLwnnJbipbw7NLMqURkfv2KP2yucjfP+
TrRZdofrAnuznnHKeNfibqfsCfxlkgcmzm8i79KRdNkWdZSKZpWyp0VBEcTv2A4U
4oBnlBfxfFwK/B76t9W/1000YebqJj48dghHqMgOiZ5TsFQ65blE/WpID5lnilJ7
AXysbhy/YgrBFxkxx7uojspZ3iLAd28u5mNERzAImfDbx6FjExxh1fWPG6xgsAQj
mwHw5688HN8BQ5qBjXZXtU63pCpYi7+f0kquDmPlWiOiwM9i6+y3kYOCcpg0XBz9
W45CtbH+51IEc/I+Td1fD9h0bX0oeh5zsDX0Zwy+qPgMfiDmQd6bYoSL1cu6LDbY
3yP1sb1QRUr9bix8a3mzM1hCg0ll1vs/1Qm7RdCYhNW7U+9lmyfMrP0Nu15W8EhK
zUimfsKmSeVA459UMYkDYKlPqpkLnsa6b3SBTEvF5b5fs8MGpNlNaEd+VGIAbey7
dTo3ufrywhCseGkUqVEyBCw1Oq7BGFK2Fz7GFjdyPcWpOm14bXtyd9XPlO3k0R6E
cR7DNclXBGk6fcjtiIQayr6V58xykVeIAA49cW+m41hxYMes7T+009ZjwQhNsixV
dEq/irtC0OqmBfrF5j+7d2hPtoEg9vb3WN0lGY+fBwHrkkr3+Y/R5ZoWZik+hISy
1yStTP5qQkzkUHZhM9BPAr5yTy67RjGGGKLfUkaI2lhhUH+PvO6CexLakdKBfOIM
+8v1LMNR/gYnxfGvqTpLhiWhSya061SWn72WOHSTWHaw2+qBNzlFlT0+d2ESgU2s
26xccmK6k4rkVpsOKNjgpQ/x8tKTOllw9BW4TlucidyZzc2zfuGwy1CvUWa9GlJo
imnFG6re5ZaF65UzFz0+zFjY8pL2ysfHl9RjElipwdH3X15jEj3n8kU1hw/0Pu96
vmy/Fr56FVaMqIXEZytepfiBbjRjXiLwC4JPsYnpEAZkKYmR7nGJcN4TVyCJmcIC
ddelG9ETVXTJAWC61B3NYnrbaZcKAmBrI4BzYA+bc9ToQYf7AkKhIiYmfUVGnGYX
2snUbAQJeK0zX0ryrxIcS6m5k23oTkigShOCC6m1wNRbnp7gpmOWl7idV/9AOV1K
Oz3vzr3+MkgUmhH2jrrMz76uwhQK1w0K4EduOWrnH5H03/8QYBKVp6WkfqIpmUok
qkXi4G0bVmh2iyuQccZFbE0iqSdjD3k6PG/wy8rDtybwOsa8+M0gWFdcNmXRr5TM
oW2wYz/GCQm7x8DDWby/wiuTDQEKT5iGbBcEKhSjhz4VmRPWjbgjx4+EXvhXeuLX
+Cuuzgts13hTaWGytv5nMQVTKSqRu+InXrH5m/ezX1v49AdEJYhAZebxg8+chudj
KkrcMNEtpzCENHMEiuCz9LxklnDk67b8oAmx1Xect9ry43vAl46/pJzwJOlfr723
wXh7B3DvXBiVCsLoux1KFDd6fIysDjUO5K1UoRfd6Y/sXwQlziqrZ/Pf1pJ9Mz1n
zf1w9r4Pqh1rJ3G4l/XSIjuw4k4JZjnzbyVpwjbpSL9xlht8cdgQgS6GKkLW/9iL
AcLpgD5vLqhIz9Rhxy0pveYQhUq/ms06/GzjQcfidJOIoCe157s579vqSNvYcfXL
gmZWCAeNo5kCyveZ4Tbjlw==
`protect END_PROTECTED
