`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BOK53qdQAv9jEPSCNO7Cx7Qp0Su/fwAI4Bh+XPV4D03LujEzr+I4UHxBCj2ZL2vq
6SyryG8ooDanhZpdJ5bPOvme3DFChS68DIq53OMYHpbO3hdkcr8H270NVT4O97CU
+CHTVKi7u4OyTlV5u4cBIG385D9MF4cesLDesolOgRwzdw5RnREai/bSFVpedRDe
US43anH85JvxKZWDTnRj4T5ObZ9vESoEQ8ES2rdNGLTboraNq+0VMjj4zwq5F/RX
gD3STR8mBUuGGdnb8Y2sPpbxKVgTzH3iUnS1IodUPiwnGvoft/1jEBoNN0AGj3+i
P3OaPG3en6zT58gCspqKXhgP56jHrcwLC+Pyix5ZcpetI0NJtwi424uHK2pJJWDr
VGK9UCd4Wv0VENhgbqKELuiu3mNfYgg1czjTWK8gLQ9rofku0A0Sgn+MnXh1dlM8
vhwd0ozgXoRknHVugnHbdD3ABLhsgVEGaUp2uPebU7gK/WMH1x8kRUSMX0nG+kjP
F0uom4I3YrxQVjK/X7Igrmm+P8W5YXxTkQWcfgbm5mWLLg+TvCWpKqkeU3W2WAV7
bA9ZGbKlDHSVl9SiqdNxFZFEjlYmu3oeBN0NlvMFJsqbDjhnS2HJhH5C+eI+tZwy
ltdxczOvJtJcVrVJPZKffUtnmwDlqk8+f6B54eoBNTKZJCYY6jwkzzaUv3EFLFsU
SKJ8Hng5cLYFGUMAYZGUGYRCYVW5qzK5FsgZzlmuIy55fTFHjjHc9vF8YM+As3hh
XJYm2WKR5OBaOoqaa5cGQmTsgnvW95UjU7NqJwKgUui/Itw7qLKSs5Ug/2z9KL7z
lQVetb7fQJPvBy7EWshGTKrU4t8vleORJSXHUPV2+Y1e+2CDXjUuV00oDEQuGO0h
K73VHb3/1V7HhXxbi243Cw==
`protect END_PROTECTED
