`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
79odnm1iHhIBcpgKxpqfhGYVwqqKB6Es5aADyyVXpN3ZJW89Dt9L6CpIYgN7Gqvr
mYPEck4d/GNw9NnUmu3/OaL+Z5zJcPzfKrajkZ4oFET90YcpLeRM3IM6mfKdD1Ic
qP43z0lkCo86Sf1g7GfTTb0OgEKtcB93uFtnMqEMxnWvFLyK+TRic5y39PjOir1y
vJW3re52LGWezLP+f+xRYIMmlxEV1bTX2VkCbDW+rEBDyZR8hNdCOx5uz80hUxCM
U8PBbw9VqWjmQXXlZ68E5rAZTwnitvnDi+Pjt+EiyLKao7dJ48acfayz3bC4exao
q7k1emuEc2SUzRLu97GDvpoPT9C13/bBiike/c0QyCpyUC31jbB+BFNDuj3zfJgZ
baOhv8jtFqnlYJ8Y6PlpLZUfa2ZptUTSsqG23961VXEKvvqqi9LqmB2egR+sxKsy
Xl4LH42sk67pIyTqQ4G5wcrEIPwLa3tNUfw9PlO+K1PkKTVaznj1L4oiHfzBbmWY
uQ9fXcZH/Wsx6X20+8ct0Ii7z6QLyFtV/e8DEXToePL8aP+W/3cIxomXltM3g/ty
moR98h2OYwfgIjXENCMt2Sa4YztdHDS5CshhHkWq+j4cs3k64SVtjukbRIc7CFVT
5B/O8ZStVVvuEJX3pS/N8tWE8ETVvUklSZ/W9egxONn3MHIAlEJFTmDV+CBH7wzB
i4pEPLKWAikrnNNwhmbeD/OEAeCAXNkedb/4R67mJv1S8haYI73dP/c5LdsB+Zmv
oS5lT4XcQjGY5W1CuQHvvImN49L4Mbv5Ax5AYmuxkSBuVtXOZ3IUDGVQW0TeL/GU
ndxjUzASGCg1Q78xiCvkmMgAxV/GLjn/fVN+G2tNByY04SOuo9fCGA3s+htdZlJ+
LVRTxPCE2h3E4qynny0Xct3Ye6Y8vxl4xVW2RcMplSX7XByPoVtVsowAPob5Dnpe
qcOrd+NXfftQ9+T3oWJIYKkvYm6wtM/spyaeIFukai3r4A+2ZaO0VVfK12D7jGLv
fClzUkoR+/ZbMkBecR9mywbOrUWf2W3J/oPgRI73X1qZypyf268NuXT89OFD8k6f
mjFQCGBgLsdnv5skz1UzdeEGvD6c48WsY36WgJ0w2/PtAsssLl095QKR0i1GBvQp
9KHYwLJAeaIF1fWy0byOT1jZw8xwaVRGRVU4XIfTYtbIlvFr6f0uWOqXtMomM6le
V7yyp3JzDqBeoZmfky68XZIi8Q5kW6yIZaYf8c7wL6hutWCYJ3KcI7Ct6ZozGp7F
2v/77BI/PCOEpZ26AOSjq2jGxpgsERVIhBV13KoJXiWAdKy8maz8jxOpKC4vWOTo
Mfqogb3yPbqo3Q/9mepAvGx/L2P+uEJogxKQyohtGosv7bteAQ43K4495294uUg3
SxK5gaWpJyYe1A0cK93W+M07GK02oz+385e1ZmuB9OlyIauDjKsn4vtzpFGvQ9ji
NQMuanMrOfB0E30IyG8OVvJfWll6U3OHvgFgnjpMmYfVmeveEewBPet5BKG/MQQo
+fcmtq2bVoyGzN/UI7M2Y3UiGbikFi+hACTqWgtbOD35r5/M9SVm6yW6EP1r/PRu
RzuQU02hP5JaopI3JKDr72gdlA6bvPW1uVwaZoJi5fWvx9CSQtsyG0sVMhcfGNNX
fGrTtAeTeKgVrRTDijrHgE6VGGUc+vQKG2iM+JMaPSZgtMHWq0YW4Lil31BfPYGn
Xf7Ahhz14HodYAFz746BtjZSiTjjwhcoYG3GdYX5lccV1aNWxCqH4pis1znexmM3
VuGeLbdpk1bNGmyhRYHv33tsZB2+v6wExLmVvdxI2EQiE41Xjj3uvXwlsHDHOCpv
og9UzhAfglpFssncXKzy6+6LDgwlcEYKJyEEGYd5jJmlzskplqb2aeKZdRphVLRz
UYD1hR9rxEsu3CftFiSPOayRWElOEYQwdwlxLUSJv5hTAc3rciSMXjYT6/eedQPA
5Z8ZBwlnbb3lW4a+YsZwIjl1YN++VsGNGyAC+Ng7tz20xxN/S+3XG7bqcq1S7w1F
6sOU6h2hMJdl+JzKNyb+F7+eIj8xnB9BTdpUQUg0ZQOb7CwrLwK/eOwyLbjOBhfg
MdUpeFkpLSQMjdTAx/OVp1J043q/5ij8laFGJd9z4g9TaV30aMN57omgJF1zMTE4
P8sDs0yCnTwS2xZSZru8fdLa67HbhA32CkP5VijCPak1b0GN7LygrV3FETIIA9oG
zqujJuUSa/cots/F7+fnGwWaWRcdBq3YoHOj0O9c23zDXUFGFh+TmtDqK+zcURYn
Mgj65zpalPQ43e5gt57dJGKofUD9bHSM8ph+YxcvrmDa02va49V2kpXLuM+g/kY2
3v5wyYI+AyW8jgr3kfxG0lCl5XVL3XS+12EDUE1rzUjKRXkPnbnmS1FAAy4ag4hZ
hbO7LtNwf4fGXRxtIkVd28HgZfLqQ1K/IvfbNNecrWG9HqWeu9bhCu2Co+JnaVL6
FO/Ks3vjAz5ga3JI4PQo8EDk30FiFzz2nuDXgfskBT8F+F6wm2wiaJGQOdLwm7+U
JmA+i70ouX4LncY521agIbnNZ43Kg1GYxpYqbf5wc29HDlfimkgOpxxdT8rWKTm9
Z9OgPjFWszAjiPTguInP3a7gwQNIF/TkGkT5Hls+AqV3SEmW+PvyBlZc4KEA10hc
2tdvgtqeaH6JXrH60KS3g2RFdiQ7GARJTlHNJOjV3FSs3yTHkY/tWGCcb6Vswl3j
agUMBxQzRqYOeQlkh6qfk09dW9sRH3ssydBhz8NeVb8JB/C3HAdRfQlW7Ka6XLaA
L4LWILhjl5p7nq6RJfQ+vMV8flYLL/HQw2gU1HQwIyWskASGm6KyYcmKcJ+x7hMM
TAVBEgV+wHlzQ+bY+zu+ATrJdyPVu6vaiGH7j5O0ZI0OV+LNGiBwHQtSizcbD1c4
9tO/t+jCNcs84k5UDsuIbiJ9kRqbijvsKLLa3CIYabiVgL2PyHGLAy8MZ4q/SD+W
YVztbCrc9cgbbLEiXrihsK2ZHgeITuEx09kFyeRHdPUoxrVGTaisRz1RVN9SBOib
/7lv6jvcUCn/jDcyj40mvNDbmWqMuckqFQbOqkVp2LtrUqq50Etmku8M4d6DCIIv
ZGNk9SgNC4WTaqc91ruZYeGEpthkTE9vkNG5DlQ8fYn+KmZHbeCkUieHs2nalFHj
goteb7ar2WRiMyDY8+xBqOQwgsUa/7S8mAPy+BxisrKOVjg021Yg9IwjZBdDyLK1
xuSq+gw4+hYh3nK7t27Aq54gFPUAOdWjUArczipTESpAg6H1+ada89YR0tGn6yxm
ceH9JOnBDGzRw91Cl1Dfh0zK/oKPQ/hd2S/i0bq1YFvE/o/OKNLBO6oLe3dCDSZt
qVq+yANS4gk2TC8xfblrsY12xcvksdJ0aYwyBDTgzsDBy0K23/CT37X3VVUbs1S2
m6F6YsccRw+tmN35AAxKIW+cAAcjCfLjllPPB/gFUQEckWMHJ/2dNsLu1VRV2Axw
hlw76JZtUQDvZKRZWbl5QsIQezUJGInwi2/3cSUFtUDr50m4J4qvZ5GpW6f3xrhB
28GHGvy6G0rn9z0180uHpNn4vdAf94+W8SUaNitjJa64FWxlB8sVsloopYbTKheT
4HppBUj+zjYTRYhjSoe77/LlCL5kTc++TXOjJViaQo/nKvtFYN3X2V9Ihe3kCJiv
phJJbRjUQO0wkM0PezfAURYBoEEmmeT6LGTE3f9skULbin5jnKu4zvDKbDxLLX9m
02WPDMlzHNQF5pQ91j+x6PFP/DNmx8XWfB1LeBCcWU7u3DF4u+hrxapKeQIwViK+
7ykWxw/GYO1v4MKh0JgB9eWmXzX9YsBw095p9l5gymD2MmwSUUtf0ye2/W+VJOfN
9Zap7wV7nbUSbWSK2TX67H3fRU9GH24iQ5N8IROJlQFfIWcqrhmDuWkKOOWAAFAP
OQLM2MxcnpxKReVhnp/Z9qj6CI9lqdethJOntPhqpeavDwr5UcE/0guwzR31hZt8
i2GpizJ934u0CwRSkUddACpg8n4IzT+2eKHVdc3pa/N+FA9Cog55ddI+d4pR/+C/
1U+i02YH1pNLzFPzBcxgiXPRaiMYlTCo3UiFh46tvrG5d3U7Yd6KJeqp/puTacp5
SqLALnP5NOAMlx5h5sa4ZeG5t2nZdIv5+FKBjuznRBef1/6hdihf+k4+zFJr2sju
06mvuQpZMHuhzW8igFrUx4y8mqqz73RWh4nT48SXeGxhFQAHXn4/yumnV1g/1D0N
gQ6HgOIbgjsUmZfJIk/DViurElMMM5o5ZpMg10Ne9A51CthXMqAQ4qnAgbBLENL6
c2jkfTMzF1+6Qvg40Q1KeqbdHsjtPwcFlbLF5VRpoxwnFMWueS//oDpT3W8vZ6Ae
sz9jPrPPZn0zshzEZNTKJP4z8w22G1iCLG2VypmykYkESPa39Qo/QPC2UKm7mynq
fdD4KF1zUy9pfl0nmRz3wftYByCYXH/qbqypqJgUX36CPlBWm+B2k2HYF+afXmHO
wcncOQjRwqjMBq8CLcIo3NHQ55SirdryRnJIFk5JdY10p55r9EvmMYSIMPMiIMxq
O6h7pGbNYDX6rbcJHqd3GYqLBAEBREAe5GQUW1jOGay89d4pvcINwmOmasdMdG19
WN07zOAfUQzW4/GXWWMwTm53wbaus3tn+PJC/LPK0BwUUrOANvLbRSGt34r5k+5k
RtA09WacAmHoHa1vGmVn7uO5fzh5zNADrqEbv7hL76Q1sAcZv6XT4m77CGuycX6I
Ys5yJVG5O0DL8EpHfUpu8zPk+Pq/IEg7F87dhB1KziAKmUVFpg5hEkLf+VWS2Oe3
gSb036cVYT8SF5IAkVLLXZYAG4C/ZTNjU6lDaufFCLTC9OI7xjzP73lcAYyM1TSl
Y2pzTbXiUyomG2STW/GALnv1cs0CXfRSJeScOJv1xWTQ+EhINoa46qkdoIUtYxXI
Aa0jlp68ej/lQTlQujxzLX9jnlPTnK1f5a2DZdJTRf6h5Gj8w3fLyBcAFDoIyjY5
+R6WwY6E4hkNc9MdtZrMt/3BZYRgRrDNOMKvzvqd6HsSktZgvmmIqLyQtEJsT1/z
e9BcD9eJ/HgHT1AgTsTq9fONx8iwU2ORR577TX4X1lmaZ5fOfwL4KVilvc9n1Q5G
e9tRs3K7zJeS3qxmbxgfbq6aKUXpBlN12EUewEqBIty1WN0p1a4a7oPYpOA+3t7t
UWih4t/L2vprKIdaXuPhQfm8ufgdXo+Hix7hu8gHJ7zZdukCOdCn6mSxGtsXtY7t
u87sYp+QdTFha387f9IRA1f0bHszgOCJy/8yzBuUQz7k1wXuRXBy+3tZ5LM1zxyF
VqQXQWY0mHCUsbzqLKcj4fEvgX9WaDKbqjbDPQ9/bVNZrzLkcidcvA8BmnwL/ok/
ZEG7hu3GhRsaWdpUei48X3Jsb6Dl5Mg3CoZwzcJlw5/yT4TpemflfAcoZpTSq+3w
ddBXechkx37/SFAj14mf5b15o88J+MTq2pobDtN5uP25Kclz172PBr/1/bmeolKW
HguFMSrg2+omrvOZAgVI6aIUsRdtK78d/Nal8bbcp33gu7n4Nfrlub+UXJ0/k0KF
PZs7n5L9ujueouSIn6TZhpjnM6YzrFDjVBaylI1ds00Jl0jUqiE4oRlPvbFQXj8Z
qeuDo9pM6XycVIR6iUFxwGtOyXQI+L2p8Mnh40VBi3rCxemFrezugmuClawUjep3
JI02vcKQ09Otjt/q1RQ8U7VDUJdR5ZJ4+jiRXycaFFumxQ/7R+W9fW4ijtRPeTz4
MlLYzihtMrF0FvBn70i/WDqbNbnF0ppzfHOeu3bau/SRN2aYwuilReo6gJ6xAqIb
+anzq/BXVW0zjvxom6Y8TNCR+fMTIJI5Neoon6YLW2gq4mSn2pw1BZ42zv8fenR2
z7yY/u2I1CF3xg62LrG1fFsxLotxAZ3QvjJSnFq20D6Ucy3i01gXGIfovC07Qzw0
Rhn4pf0hK1aHRCxVK70ce8Sq5QWhxXwLsgBGIJT58XOXFXoajYZo8KmrylkxISm3
z0Ze4v6QQ+VimVaZlgd6E1lhH7VJapK4F4887gdOvJDcmyYFIivytqmCWHK2RrwM
OuJ/o5J5ZjgC13Ykw5IqITswa4oaLz1aGM6b5VCSJgyQ9Y1nO050gpevN3IGsUXE
6gjK1pXotZx2JVNPxJxGO7/19HmYzOOJFoAHzLmCq6ON/nF5nA9fANL3tx11hKYG
1Fw7Uu7+nrn1srJSxyd4yTZiamMb3U9iMMGKQl5ZUPfyXn6Dyk1mFFvQt8HDT8An
B5/G8Ak+qL8QzCFCSImDqK9ETz7J+5ZLAJvrWSvOrnk6wBMUaevz6TSTD1D+hqnj
PNCmrvKtAgvvhUfx4CM0VFRQdFPkjHNu8Aq2ymH4bhDrzNk6kUl0zo/Fzmjn1OQR
Tj5Rep/1vJpMK0ynUTFi5v99+BZz22UTMcjk7Cpr4dkdR8F8fcvfozk6TICTe3l5
7y4XEAXjm/Fy1sw582IDrqM/XIad4gnz/U78fjRmtm9fYFQBpPOg+RbpYc+XS730
B4HEQRdrpz0zBGOiMKYFqQ7fN6vknzlkCrfkHe/VyY+R9E/2wvcbU7xS4oODPMCM
ywqAW55lMZq7PeACiw9nmztYHFm2zWgwH5iVSEh2q6yRTAZGEA8+AmZawFDo6/gc
uq9i0/dpg1C5zrlUHF1X/Vm+J1gAqO0u1OhMbUCYDS2M0kEN1cWNn4NFx4EOe2PD
7N1awXmy37w4UHWyaoj2qNWnfoLoMmI85GlCLHQFWigt2A/IlpeHgWSecBBVrgmQ
yF/GFzoFkTavhaCsaS00f+nOMyNfKhGP/Jawsg2Exsv+aF0rc60p4ACq/3i/9GP0
ZLmYtCK6LKskVVA2sOsyylgKU+31nnA264IjgesoaWj3F/sEi3Hm3LlyZls1zogD
tRq9XcJ1tjn+1cQ8Ii/bKrUQ6J15dtK9+EfIAVFd3+UQh5u7UkLH+qEXJ0qp9HCq
gNL3prOPIpjQl89nbhjSgQTKechtJbxwzlevwM9e2Quv/hc6BApPdSOHD18A5i8V
SWbmnSCKkU4WT0ZxQ9gDklqtQhRLlO6lNRlq/Gz6/b9Dkpe1c+GfbF/pZxeHENDy
HptZ3WmzsUt3LEBwhGg5y6/FNaOU1Nl6n+BJESIZYfhG7Go5lwxn/Mz8IMVJKXo6
JDR2G6io8jA/WxCqcusEm899iu6+SOEiqunNQ/VdSQia7W7c9a8a/m24TiAQiuFX
eVR+zpsIiZ6NHQa8DvyVms+587NgiXwSkUKDoe3RHzZ5UrKql+X8lzEfEPV4YB25
tW40HnGKRO1rhzrkyIH00X3wGjNTpxqBYMP9STrjPTyTa7YHXdrjac7rX87ozE30
MZx2nywrXoIDal1BBoEzsoy4WuwFShQmofqA801Re8ky5JhsRuv+EsQuN7D3+OLN
nbVDvKG/6/ObWv+zKONNm67LAw7ifDQXBmEY+B/kyIiCwnkS2rIp6FB/mbT7Et/i
ThHWvQ2ICEggQa3TpsQx76nYrf82tUGIKEVJt21hSi5ED7WelccuDR+vvxe0Ul7b
+72C2pAPxzPV12Emg9FD5BR+bDRTN4eMIF3p89BN4ow+Glcvooq7uDcDposmqpBJ
uOdx3j/X6pCnuSY2D4GqPGOSeVGLaFwO7j6Hjwtf2VNfd7LCxOP1LXVzGZmWKMJ4
MEeNuMklciqmFXp6AitM2SoSwMROdtat/EhjRfeDZ1IvPauFc7a80emX2bPo7lOY
MzfLLYk7krqqNMmv9Y4jXFVLHdNRGDweh/vQOgIEFWirYTn2QyB3GRqNKMHAqBF5
yPHSlDmepZHntpWMPX0NkdAssP6hXQegHrANnlDLESkNhZL4hcQvVWqMYaFoMgnO
kSNQj0A3kbLOdtpG0OcC6r6NvQgH97qkjtc8H2wREHDD2qr8+jf4uE2YuTbV64vx
XZcZjhB1wjABIGEztOLCSeTNqpQ2jUSgfqL2qmDY6RD9VYWDQFUg+hFFc4XsFTsT
ntRh+HthMTuvU029pSSmypKHIhKXDKgsKgKXGJiJhG71H3331CTkprrb0zwwiBKw
E1sxlUg/zcQytcJ6ksdrDAfD6h2UgTrqgM2NKL0xndFR7zb4BpdLnwDANRIvx+qH
apdKKHYxQXJvErHVK3jruHO47LR95JY75cMDi4ER/2VYXmfAoDhro8bBVPsbyuUl
kgDnVoMd/3piPVtP0CURQWDntE/a9+CcawFS8x7eaLD475c3C79lKUinE/Sq1//a
9KKVoBo2GYgyFAXzkRg+ieIF0MiCDxc2VwNgxr6VIqoaJ+f7eBRFXaq+zIXYQ8BS
O+fgeww1mBTP35yBEwjPAs61bkHtcFPzswP041v/HyH3iHbrNtTUpRyVEzdjoXUw
lZcCEgP57856FDj8XP9ov3yFJqX6Lw0DMRnS9BLa2cM4v7MG9c15GA02mTlNVzkR
6+huxxnJXYAlcELgH+C0DqedbrK8GBCEJoM8FhiBciQUp4RgoXbl0h6gQZ3jR7fo
JSSalAm/Yf+Q9RTFEGhuRHjEHsw1ha6UCQlg1oEXkqY6KjQ/FhcPWzh+rBFp1C0G
B2SFvga/UNQAAT9LQWyKW87gTMiBWtBLJ6Hux0S6GlgM4fNtMTK2uE55PscBnPBV
7XAk95VIogt591AkyRybniUk6MPvSkamoplWcOETrkm9sYiV1c29iHmG5gbnfT8n
p7QcIo7fQdz6/LVaL8GTrgSjd/S1h/c/gs4evMRDgYnkR8dfr3fnmM1Kidn4JZL4
XzUE91xF6eWGzBzGb6ip5zapuE8CSoDU8Qz4H+QYIdmsrRFqwWyM42TN9dPobXhp
qaVcNDGgKsDbj3w+QPBEqK6vMU3fe3qSK60szUT+aMlv9dHKDTHwDpqyCZCDAxFY
jAsG0HK8N9XkbSLEmfC+SBHXGK1CwWZgpJdtjONmY5MMi7H+8LFmbBv548h+O78W
J5y5ZzECu00C/YI193b8eJn4UoWe7n35c+6QB15U9xwwHcIZVWbL2sfx1u8v1cNA
mTRoHwtNmcBW5h0GfamVLU7zk4eOy+mGr6y2cj/qzPcIF39ic3HuyEzzFPQpqY8h
GHfevYnfaGRtor1QZO4MkweftYO92KjJezPsHOsPHPoMnyjtlXWO3pm7WU19byO+
FBrm4yE0VoJOALXUWSl/6kGM1ohyT7s6QMDXhG038lcEhJXDypJ2f1UWoCjq0Kti
8Bc2mJxhAplTsUy/XakH6yRsv3TWG6vMypq6hV8WN/O9aLPUnMsJ+yQOVAK9oG1b
8OSdM1XiLku5xJ1cGs3NNurdcS/9rfpF3oYNmD+2emzO2WDAg9V0KmVmY++rFnHP
uB23/+cINf4yFauCQeUyI2Or/uiaeKV9lm5Isp4JSnlzJVTdCrA9+EdWZESoci3s
7oKb26v5VuZjCKDB00l+1i6DmQ5Rf/BQn+h3Ysiibf/hoc349sZZar2ivMZtcPOI
NCEHhN2P9lQG3XjYGBuIpadye49+p+OqPoePKDzhydYZm/GVb9B0/Z2TNuyYH+7+
wC75tsEVU3PHQM/ZDmojJU5ljpWYzqi3ZaVeWf3Rr/CBTCEVHRtNhEssWPsDtfsK
C+lZx3WC/ksgOosfOG9Dil9yxkVjywRcFfTKU7TKLvLxzxoQIM/EDO0Y4AgRyvKB
/9qU7xTIB5ko8PoENCsX8qsS4cC8i0M3+ZjkD2jApITp76hXz5Zgpj0v2yLPA6S9
GQLMBtGj+JjBJATqaqn12Qlg9+FoEq5xSwz9rPTfmLvOc7XZaAiTkLf/dlP0LBO7
pyD0SYp2EcwOZy4UyFD0RmLSh+t/iISe6E4kpqYUe8TiezZxpLNBz144RDKbBGjV
FHttq7WVG0oG8UkQgFVxYjwS7QVmMWJhzlFNiB9NfWdrH6YsKhMEQ49ExmBRoEc7
xZJbdEjJ5h6OT5XzJ3rik5SOTUjQjhD3ivtRkxPxDeR/OD30ZPQ8iZv3xSZn85D6
agWt2PY5E5eqI/pUUkD/D47dyMDr5D3PL2b/CtC36iVXwARcjbgtHW9VP22v/YWL
3O4Pdgt9HDXXiUumoshzeaohJXgRQz8jeqM0gVwLm9w//5pySVLRU0QAXXPI44Os
82AiGdIuI54r5KePeqkOueolA0amXCHu38toink6YlE/QcDnIMN3fPnxhADLMVKP
SZ682fTp0rU1Nyl0prUvPIdXlR6FB48cWit3larKzwrFmE+LCWz8lwaWOelgA7QH
ILVTzwhCbOt16rjHfrSdshlO/suPI2f5w8F/edZpP5RoCAWpgaXibFMMRVCTAJq7
yzOlR6IuHieNTPuvl3ycpS3CSfyA6DeVNu9D6F88riNKUSBW2Ydoi2QIPxAWfRB+
kqxODuF4XnEYx17RYeOjHu3tQZR+N1y9+X0HiTlJZJM0YlHGIGq3m/sUlvc56FGi
2FvXgUFeb6BpMFlUDYGDgDtZvcSLu1KneVshn/yieyqB7l+0XNhX92Taup2CSVM7
fs9fqfOLIbYBJQO9kecz6vbCvMBvs4v2eHb5U/gNcxMW5oc2i7BeUaiMQg0RxXKi
nVmPBkfi0NTzMFa3kBwuOt4vHPB+U0XlH6+Ow7WsCanqzdyvtrrx1ex+vd+hHnXu
T8EIHWwBdPoxMt5xHrjhxP+ANvF+uJXNcjhFbJEn0zuxWuQAohq0TNEnkpkD7zpG
nW+RCwUzyF1KeUCaLEo8s9cRKDonOUrchmxUHSmc1r4aXgbGseAhs2KU3KnMNnWZ
btjOceOdQbwQc0LhLxXqKOovLYWp+fcjYuK1DdZEjamBE4Gt8+n9b8a7SFsYCdxU
bENOiOKBHOMTYTPiIEOKBe1djw7w8bv977YWnZCvxv/WCg2FpdXrPCQYjFIoJnqH
INdcc8uN8Zd29GC2S11v2WXR0FbIkXsRFAumXccjDLVu4ixPbY4lG6H9PeaQS0Nu
Wrhrej1wnKTkpaKtMJ1WtP5Aa2qGlMBaNM7aGbL1JlpR3q7a44DlGfiddrYSlToA
WiIh/ISVU1gCg1DhyYiQfsyys0aF6SMWwWLe3j+bZdF5LGPhalZJ0zREn3RIF5Lt
jVzN90c+9TnP0pZYiZbc/3hBUTt6UaQCeHjrMXFrenSHSXKdd8VL0hwtsOJZodB3
tM96UyBMohUIYdSy5uc67JBS4l0ISojJBdItp4d/BTEtKG4ePzirBzEpptkJLeuD
mNyABgkTYNGKwNk5QfDDw67dgaaA6sv+XREclN7r2GR86t4pvvDjbfi6pkUTnVAf
T1TZ+R2I02SiPMXz6L7shCIn2oJ8e+mL30BPoUyV5i9zzqStf1WEjtrlzAbCE5Nm
k760EYQ48F+2vX7GOBJ8bO5qxDPFPyzeLmzPUOfJzsk0JcsifYgws5sjsgjg4Pkx
4Jq9QAHQs5EWaHvHcVGk7OUxfY4RFLnE4lnnFCJRBrg5T7T5qtss8s+roKcxWQxk
4y1YQNkhqN0WushjRJdLxQ0+gjX1kUFB6rFCJdLjhcR9GvAANxSsMKvrTaiQqGuE
u939CvQh0EKBSBxyKU6yXKZlwyybADWcXhDUBzgd6mgYQCRytFsG4i3/AES0YwF9
5Quxh+pF/+Zq9c1P/6+C0PPrRUud4pzvmQYcwznkk2SigsBK9QFQYGxjVeMDwMBx
2ggX4r7IXzf784SiD/GWNgvQltxA1Wu9MFul02gUA9dbSXNV+1cnUG5mVpJxaYZb
08VynXkJGFzvsFiUCtqWAYhFuy2VdktmTXZ3U8pj7QON/trBrZdndE/wWLFEoE4U
c9+eY34q0J8UmPOxjlpUEXonRJa1Lnjyo9it2yY8WigtH2P1GfOZcHv56TxqJPBg
ZE/GwjZgCO0Aww4H5iG2mqaDNm8F4aPiHhvb4KU8HYO/HC9PSgLc819jFLDaP6Bx
PCfo/cyJQaoghhsnWS3tD92oWb0CxddbZZYHrekmE+PYL6gEJ5BEp2xiYp5hpI1Q
C1xwMZaOPfijrmv8/eUYzPBQPrkb10pi3ZgMsYihzhrxBnzzq+xz7bnL9rtbfVRv
CgKrY5m1ChJ3L5fYeedBDKTMtPdnxsEdtI5mSzFJ+TR1vCWavP54GCqrwzdw9Pub
HEy4Eptbj+tB2/fzbDqS1DMObH6oGfzzjoP1MCzEg8Tmvzw71JmM1KQPdEJLunxq
yQMZMwbDctHh7S9kg8totQIffjA5ioTVw3WhIL0iFLpWj1IaBjrYYi9ppEXoi81P
+ndCnUOoSLaB2somLJaslWlnrfkuo9wKphg77W52p2P3rfkyLSSy712y2aS//3E8
p/irlYD83qpaauPwh26vZal0R6uHaRqJUfxHQKxLVUkSOYAQvbl1GrcSkvLUMCbz
aV6os3ZcKpXdp4IfSj5gHpXvXuOfA4Ln5icUnsETdNL8M1TqdlDM7gcGCxE0TEIq
7ON08xiOBvIthHHpthmRryjZ8n6DPYXI8rA8ZU7EUhBBIVW3uFgpcyrUUOlKUlJS
vFr8yPsZc6Wqa78HPyQ6Xi0eOgsH8cA/q9NEAaIwuuCmZbziRmQiJPqPCL+oFsSE
B50HQkT/AXgLg1Of0oQqyM50hFKPcZRGOIVkIf4bj3d25dekaCp0p50p7jlS2lwW
3sVawHQ3M4yKLjBGOSvhA6plXvmVj2ttTq/y4TntVFxwnOb/wCTzAyXdQlYMDN4d
RCet16ntW1/NwhseOdpzHIWIYWwgzvn5EMsKuPy/n30pBCZDTFGdkR9Y/qbbdkQi
ZHO2myrnJral5bArYgZEa8kwu8VtWLJyTpKC8/rwAq++abFtrzvLgzTtgXvob1Gu
0OVxq6V4AwVzKTtyyQ67+GV0eZu+045fEo2yKqAUZBa9hDaO1EzGKE7EhsIVRfsk
n20c/pkeiQPTB8mlenyXsXGQNKzyjPuJQm8FeCHi8PSn0msNdcAUQsCslUHQBFXr
+l0BKe9a8LX9gjoRU9Bf8InF/XaQEBdIz/K3hGHK51Vj6+yTxpwfNw+LS4KyPkAE
vb/mkoVMieB8aXHZn52uMcjLN7i+r6LGcJrdm1KfJtXL4bQRXvFOpR4BLMSaduko
7VnU6bXnXpuCtuyObMgIi9gE/sD789otBrOqZJZXVzz25mfihbdJQAZvj8Y1qaYs
ZEsYvUpUu88tH/IUHHXDmIN+/oZvaR8CEOZj7ruXTMpT9JKnLQSAWPrGaM75Qsj/
A8Mnv2XHHPmidOPKoxZ8bva5WgSPAtZaM0luzg87J09K5W8MdAM6ugcYVs1IVled
pggepptJvzs4HcQNwVT3QTthaylxeLXOPBEHWiQ1mGV5dm8H9SzSnZSu63XSd1Wg
/p2fIHnFMKEkcu6cHy17B69h6Vdnt9iVaFWBiIJoatroCu4LB3Q/wlg8C+/fhvRs
jJmLZbWMXEVp/81EOLkaAFeU51gNIHl7bgFWzGAziQKUU/NQjFmaJVvnDDs2oECd
h2gPr3/Ih8d1u52cyC7FEqJwurk2nnOdOYbN4sStdhN7rMILSS5/40NM7NSuZNg6
ds2WXHt/vls7MNGkOOjZ99H9+jfKNFUG72cz/bYtSg1QR1LsetHtPL1yf7XSAWKj
rGd0u5B7M77MuCFPBT1Rbpw0CsSQz38cyPsFtbDUgL2zElbG+AWu3EET0JMZnz5L
yHSo/l44BZPItwNlfGzR4yWNg/HRc4Lf76Zl7xQ2mi6TNmsz/HhdR99Ylzet+1UD
65b/krox4qCKczWQE7h45c8Hho0PUcy0a0yvAoIXKEjDyT+BtrJ7m0nxxhhWXKYy
+QhlbvhcdbmaOAX3xpAoVzMo7rcArdzzrCHxsD+WzUy0MuSNJvn4lXLRiRGAY/0l
G4AvJDleDuN2W8ZM4xl4aIoAUgSwTR5AAI1ePJtKnEDejoOaY+kgsjOKMWJgWjHc
vWPNYDPi663QjUzkDEhNk3+PvvOvfvQnipEZAESYTvz5pBJ9i7IJdMCOI0f7sgMx
g6pOJPilhkydW07esMd+qRfVa93pLd9is5Eg3CdK2ZxWzTREzaE/QxaIz+QeMiNi
P/h4Rr21s60Na+wTZ6CkLcp6XxtwuVqKDZpeKOxvhr4xG36w8ZRq5ZSsJbYyJ0O4
MfQt5M0mx+artKUwqp0LHhuq2acUxDxqI/mS/oAILueUZC4jTCodRtOlQ1kROhHs
BjT9NLi6cJE5+GY8QJPBjDE0Jgdu1Fq6mHimwOTB7CfezCy4RKByH+nFP9XbLpQD
A9ITUWDP/x/wlqHU3fik9wwwtr5xmgxu2PKytAU8oL2ffGagkU7L65VgZ1/LKquk
7+dIuKF32LNjpQ1B53pkOJQhlJwZxTk5SM1o0J0f0JsIA0JOiFvI+gSWnUMaJJE/
/3NB2lvWrhKpdcf93FTAtcA2KWEaSkpcHw+ot16o/OspkMQ9D07zyvNp+d3aLiks
GvlNMK45QC7s9UUhOMqafBOilv5Ypdx72XV2LOKmW6xwdJDoeapdbnrtZjRc5x8l
W7S+oH6zgnXWztaijmCDLmd6QUUCegbJPAjnUrc98N97XQekiERGrX6xpFs9BpHj
uJcNtWT1fhiJ1DTpo3QTaUGBxYXotoha1YYlYZqv07ui5COEUCl/Ma4ldvfv6uV7
uEUN0NChnHRQe1HZzuoibtk9dF/AaGsoruR76ufoy4nJxGxzTFjzqY/D3uBdiYMf
kNkUQs+u5owh4KjWwU8IH/YH0psM/vaXvwM5y2MPDPt/yhZXouUKK5m40IxBTYu4
M/oyaE7lkOSvhyuCYvkKGwd3esWdZIPuZ+ndNXXNX9GcscfneLndm+Kt7C6t7uN7
BT85XG8fKX3hcrP6IdVs6ArScagZCMUrdYtwGjoU0Eph7SH3xx3Uw9F0fOWGdx+u
jTbTRA/uf8QBB51oRa0PbAd6rEEsfjXKBaVlu7CbtIgAMOEs3loYZEa4eY1n6/83
cg/5/9P/sInijp3UbVek4Te8PTjDBFZJc2D8CZryJnWcfv5yvcgAqgNQaiLHQnlc
wWizxNp9YMziYfXpG2eLGe1iQWBbr0v6PMjUQ5veX6236DjOttIFQ7MN0AJ35tC7
qXHZ11rJ+hjJ5qCXKn25AeY2J5hCeq0JEydDXsgXzEP9eIv5iO+FNlRBHYwHwKZt
Gj679s0XYOHn2vu62HKmaUU+mmnrP4ymF2qW6DudRfguPqo3XMSA8lPuOXAUetBk
YvHBCZ17yIdYtTGLWKQ5Cfv6AJRvnj5xO8tJSvtzHAmXPKWLjpxEOQCkSNofk7F7
ujXzl7QAxEZSu1hu/Mv0DvdwPiXT3HTJ259lj6si7lRPzvAGK70ltA0YXb84Kyqc
ztAYkfxuikIWDq4K9t0B+ULHuotLvYkICdE4vo4ix/qHmbPIOtXkd0vtsEk6XwoX
QSz3/24TkgtsyHCVJ68KSGRzEAhsPzvTS9/KzsxaekgMizgSlf2RdeAI9qdkhmp5
75H3NDn2KD0bjPozox4Vnn6Q95SjLCEdM4zgzI8+9atyw56U7Z9dQCpB7hJq07Uu
wDppiZ2QspeFDMvcrydBgfZ0kX598USdRSshYOPAfvxfTmYvC4lGc04nmDYqrrB5
B6qLxjmgYxz24YHwCo/kep2T30hOOWnLqB7+Q18C/5hWvyOohJ1vou1yW46qOzbv
vlQ56fG1+OizgvHOFnNxwpyyocueKVutWKFWnW3zGVrzdxA+WLIc9I2+NkfgXILg
MOi+YalmF123XjO4KQ9xoIq3TL3AdfWm1pVtdIBmEOtI/35Uw4KcC8PJ80hngO9J
ZJbsp2p7GS/OFocOfIs2mz2CA5cfIyR4N7E5Q34QnPyNlaikgHAcFj7d8B9TQ2FW
j8S8Y8Dk949hBV9nhI60cUlyGRe1vaIb5Z/kUjNEwFvXpNTViUJ4ryA0xM1+GccW
yTvQNe5BW4fh9n2vdt2Osi/3OzX6ewH95ms99ooyUs+DGfq4d8BTVC4T2GCIj1+U
8SUQTsWi+oIJEwXu/ajqbiy1bmdveEYrzSgeeuN19SQDbNlDj+MlAD04dr65pWcy
coGPNBt+ioSTvVQFn6iUbjGyIlftSnAzSp7Ib3XRDS8tILhQat1kv7P2S+1f6z9C
5LNI3UiXeVuCXprjdEjsJfIzHAA+n0l+M+ej6bnuS1+HKzeK4Sfp66qswLGW1EJa
LRtaRlCAoo0HSpHcyG7KPyKMoXAZlUnow4nVpgZBL6GSeGBEL/r/aLGAKyWgqRyF
Wocwe1X7z2aTnbxoCxeODT+k9ZTNxRtjNhy8Iw6yvcLb4XgAS9epBOXsvbVK1XI4
u4jzeQ05A4J4tgzz/+O5WMyC3mAAngPQi83PRfXErh3+BZAs8CGeSSAWir0BwFp2
S445BRbqAJucq4udHJknimhbOGD7bqOi+BI3hzxHpYnYj0rGENL3nts+knNGlY+E
5qLVsoeNDiSkHgithqHLwdgYj5sPCIPEDssIytE2IY4cyoix6HaIZQ/SgLWJT+sT
btJx4JWo3mDkbisFzXFnAdQbwQAR7XZO6WVgaZV6me/ocDfk3sA7I2X3GXnH3R4U
pS/3UCuBVFmgFTI+X1BEyzezDtBTspsPurge1DQ0RoRFdalQ8ffLDVC1vwbTOda9
7d/E5zHaIa3bBoZMFWbyWACpWrqbFj0OqvtMmAdaGoqPtH19RgVI5BcA2PHIwCNf
WQ9ukK6Fk6Bmy9xVMfDBUlOLk8kzTK4xNk53dPR04FDTPmmDn6aYMEb3z79Rs5eH
UHYpC3qzMHXQq8LOcHCDCDnGWRoCdLWL4qNVuoOnEQW10IEZejq0eq0iEsQ6hFsr
QVV6y2pXY00rgTI/Tiw7sNrKn7Sf9yLhr6nsCBlD66gSNCAQfryEQODICam+fIpF
VWObtJSJpeO6spGij8hsXU3jQXDm+exMOsvv7HFvEgFKSJqY+QbeHbB8ZgkMzAoW
0Ye9MNrAQiIs1yRE+wcnUvlYLqbNU1JrgU/wnpeFKX2myZWiglkwWL0lqm3N1WLh
gaRlHkxOeeIFs2/QFgLQt6mzQ6Phd6n80oAS77NWyYLxESvLHLUHgfExbdRb1Akj
DHrLKLYNNzNNbYg3DM+xxKGvdj7jDCcg83O0l69H2Y+tnYQH/W9kQ6bPRpG64I74
aCOSN6ETkwJ7bj71JtxYjtio/8Mc6ZKjG9TGwnxCx3aT1SKiCUPk+koZn+1YHByh
2JVV7Pch21rnJbhxkWmJ6BYYNXD7OTt2TVPNgNzM84eqw86fRKKiwVs+PJpXQJcG
IAujxQexBsC5BG1i/lhjW+g778eGPa6JKx2KcCj/dYigdJxjX8PcPY+SHY6TToqZ
69eqqLR8cR06dKDX9i+F4bJK2J2pPMMhLPddaF0co8BoNe7SEIsvaB6bwa5PnpXV
+wyTlJiRlh08QZOFx6kRA3/m9B4r+0X5QLXj2YENqNLo/A9lpdL98gzdSoTiQhm0
lQRaNTgT9FzVSmzJ8VWnjTrjNlTxR+fnySBnARht8q7pc1F1YJQzSgM/9XyR1ZJA
RTIYdbdRAGmzdErf04WRQqMipo1KV1XwukgZtkxwk+luUUNw1r3zCAWKmBIhBu02
p5A2oXsWAmJqSODEY0FtajojA7wsVFhvJiANciGPn2IjcA8hi/zaYjWuFZQeWJv2
nYBUIme62IpTmGZYWFmkZybryJIcFf91yXxRCpuqpJg6ZtBgYw0+EnQGAUThW1fv
s9Ihy0ge9HFGKfjSZpn1YY3Mw5bI5VuPjmtk/uJ3+dpYLmanm+dZgQFa4bGXX96A
5nDaf+8IZCUBUeFObb/tphr/cVhSaT8dJBw5nqnh0hIWACPs7nFxT3ixIUmEZfwl
mnLrHwbKJ8TUayBqBB8wH0WYc6ktrGyUYk+OZH8DXM6u/zJjIFWzcfM0jLsRIKtB
6yRFZhDjcBf+bMliGqlpQHFOtGs935ykZ5jH2pCgs4wVo/dZgMM7frOt2PfzNPtX
FzJaKZX8czhmUz1b7ARI06Sib4BQ/ATsPcm0W2iNPPDVoyGH/WVzxOIIL21QWBV0
PXHtmYtk/f6SPlzId6xxbd2bFtDgc2bU8DrT6vdmWWnSBX2Kt8uSljO3GWm9NzR3
qd3+oHp6MIMKhPesrXpWKPxJtmBEjlm3di3RB8pbHR2HCrnIJSuP5y1pbTlsmFfE
CuG/f3wAVOm3PKNAa1ORhD6sbLGol0w//cBAIwqyMEFtZ6q6QyUkStRrJu6mx34d
xljE8jhcZht6wESw+b3mWtRbxtrigVEzST8pCkubY5ORXRJdpqyOjFBthdFI+qHW
dLkgYCF62h41A/MH3R0i1q74B57euM9D32l0hkJBGuJzz51js9dkfIpQZhysQNAv
ocynasWFdaaw0SWgvAcFGx0N/hQMi+SFMvq/ogGM+87ROCXNg6knVaIf7zO9Vthh
9iLYFJnyA3cWk0M0MRfRmt+7VKqnCQCLltNXla4jU6pQ2ohJQVqPR3dMd2TlQsA6
3IYn4s0+MZaebiQusmUdtf8Vgdy1YoDZYxSMFoCYSeXW0vlcdSabCDquoBjZ464s
5eoj2eVZqfkDyFLvLnLe5o2lTmh8HKG+Pn9OKgUcDbYn5ZTT7NKb6fivFiiGWiU6
Y70F1IL6qEdT/wgOEI/wcNq1bxfRv3ZgX2bDoHDXekMGNeNeMeSvvfaAwmHJHkWr
YBu54Rw8qFHKdM54KFos7jDsiCpU1oYy/5DYZuG1D4YrlErDCxdNRDKtViGnNMyE
Vibwrxm9agVLwcta5Tz0s8dnOKW21VE8liKFTk2iFsb+9sE1l2AxOPxcDIvQoR0M
0pfMJExFkE/ZapasS+TtFRVigx5N5A4YSh/XqSz6mcxH+0G2X6MOSNuUaf1qnEzt
gk6VnmCS8qGV4kxzohkIh9f6mmRzcDHGt5FpnU608dqGeRbnwUzMa5OkkdJsx/ib
Jy1EMA0p4Ba70fsqpX3JVRoyj3OuLohBoPRfHTgUBR2sObO+So/897o40MKM4jOH
mCa9AOEvhX2Y+O03dtTetJAFZxSH++UJLbVicnrQYYe9bMHfz8A3cl8jW0Gizep0
Uj0c1vU/7GsXEXBUJaMO1DJeN0VyPEgLeHikJGlLyEKafDmAxmD+e/bsHSYQB9yo
+v8LuaNNKZbpOkUvWsaM4X+0KCH5JOOU0EMGvfCz/Ipf3r9cUTQahzBzNeYJ/b0h
auQAYPhX62V39XcyxYkyU4pWbzmY9HPLJcidinjHleADmIoPQiCsg3aVl3uB/MSo
1y4KE9i5OgED23WtNGtDDr8t96bGvTHS36/3GP5UKKbfNpFloReYaJoh3vfwQrIy
Of2jD3+1HKzroo7EvIpMNGFDRnxA8EZVoRc79VL4954Ym0vOJ9DHUgO6rmTXIRvi
oOypcGhI+bpfj2LXcl+L6mfSM6R+OGtdd5vQVREuD2iYnoJMd4inhOqv62/yI54X
Rd5QZsrTRmyqrovePx333oKRERFOpepg/Ok+TcXGWiMD56LIC9CSFEWyMIOXQgXc
wfGxduVhjaY/xp1cC7sBEhaQPqH8/hd1urtNBZaiIbrphemgk/UdpoFd3ZIpGG5N
9L0uabNPTpzhg2fPL/A3e0ZSRVy1TM+TmOJlHKyYifgKu1gMB4PmmO6ChBFMmyRn
N0eguT2cv7FZVbiP4VNxpodxMK/hjkSzwj2ABsS/5+1u9KvcO/pSM53kM+1lPSDg
I2r1bpsw9EUgQ4j/GmYuhwIka17DpUBC8bokIIMI/YvQD2yHsYGNw0gzrge2kWzr
3iDr9jW/RHMVwj/v/DSxF0KgAVbAQJs/FjMrXgTmGAM8Lh4euSObf+vVfWnjUMVH
2Zn5nV466np6+Gx+N7AkDVdkeQCUm9YwwQRrOImiOhKizRDZiBI5sx4AE6576fGH
1eG6KABhxn1UJdUXt3quH//4lF4vzI3zupXk8qhmlnPfaQd5rrFIY7/75BnPVW4r
WXOON83AQxdI9yC1sJ3w/uyKYIkGFIIMs5RLAeRQ4jtF/k7D9YUbkgdB6PjCoCT7
T0HpKaQ5Xv45MzOFA3kFlF0TvM/Q0ZEdoukC/w4creymb7lQS/9CFAQxdhud68J9
Xng6PwQ9elGtoy/KnKlNKrMCPd7RXep6P9vzQS5VDSRIZwdX70BaFoA1QGVUwfJe
eG4WBZJ/H51NNMcKke5b3zUuQlmRi7rnBu6mh/mSiGgbBFdr6kMN6kCwBMITXLYI
QODOtuhrmFpGkYO6yV2IQSVq4MogOp28Bz89Lvj/N3fcMsE4uu6vmtH076C69Wf8
s1gZQvHdH0TLzlYNn8/XqWbwgvR8VhPs6DchyES+p7E+O+RqR3d0wvpp1hf0z3xE
OONzIWbQpMHTi7k+BhXfaTyk9L0Vrsb47IQ2BRWIP8kbRLyWhSxG6lTazFPmkenY
IGHZrMk4T562bN8885/ou7NVkJ5gmJwR1VVughjyghWU3BYSN9ERF+WJXFxBp2Ca
e12sMmjQ5OtfALhUjOSQJ65HxbxGlCSxBzWko95duXqQubGasMWlcV0H1BCrgnyx
vCBvac2alSnx2OSv32SOLLYXL2mxFJxORFa0K/lv7Lz2QCK5xBFQFFrIRt6KHJRX
cSIkiQziHaCosbJjrMI4yWP7OBf9Zw6VaAC9DX0HdedCkaenBmyTMJSBTlfl4NQ2
1c8mbPB4QJ/HTPN+DPiy9G/lhBrVBfqYTrRjtIvecXGe51rouME7JL34ePnUvArH
ftb+hiw2stcjEwybh/mIb0PvGjmAfe9GwEXNyXoZvlHUWQNrmqS7R+NAFiUuZlNS
fS/FYQhf3U/EADEhNX8abQ1on8DZnEkvvHNQLHv4Q0zHeT4sgqcz5WhprZxQGuCa
G0vVmWIaN2GMT1KRWb2erxDHHGPlqcJb5DjRl8w8dM/nUP74JuhT6imD6L8pq1ur
oC/8wgDygBRyeE2AeCNxqaQ7CVi324p8n5kCecZaq8MOq6XqjG76Y7SMjgu14+jh
90sNzV59h/ozCqkw7x4F10Idm8lcF863dAeASg+okGzlwGs4Gq2GW0Q9G5zCslDE
YGtEmHshyVMlTzEGZoeEIIKorUzoe0dLB5myhgwzHQaqG/RkexJZtiNwJD3sgN34
/MgZblfihasWFo4SwzlQV2R+IhS/hUIHDNEPrlQK8VEu6hxb8jBKmgvrYeeok4cA
PhrYYryVnYfdQFcMwiXfV2SZZx0E7BFcU2Fdgk7DQvdMv1OXI5JeYhQwoYvPCI4k
Gg9RA1eYpPJa5gtv8fsSHAf0UNJJb8eiVDIBCzleIoS3O9o03RaeviOII0tOVfup
btNlffntkqkOMeD96Tee/PN66wYYCsLlPhQGQ6n/qBSEBqMmRddMnngR/ERUa2nO
IulL245mufFhjbtSN+3Zv8KT7xtOSlEvcfPQv5MXVs+sIq2w/zyr2P5TYpTq2Ack
TvfAymkRN2liVlRunpbE2J71pFg8nAhF6uPo5MuqFvV8g8STETAUDEj88avBa3Ul
dLdZHPV5ff97yyGTsUiMnLarh/GqSY3wSsNJIrGgNSUJjjgzjFJGcKdMJ/DIzV3q
PBNS46ZnjDf36HpaQEdzSqR25GkmCYsvflyRMDhppadgwE/mO/qH1LN+OmMhbGb/
uaRhureuwrQ7zoC7ZB3txn6dWWBrMysRRSH3d2/HQ/40w6/tDxZzDsBgk3e5765/
MgChORb+5+nV8di8qM8OjEWZ8Q8bB/UokSXy+20VbxC9Df+cJ+B4WMZ0h9PbY1SX
iEPVVOlOd1ESk1f2kIC0mB6HLsDptl8vkh/2/V81adTUWmzGtnrwV8a0RMOsVwIr
UN0vQcqvZ5ZSBUSBS29GPpEIG6lUiuluNKbpAYhY+VknULPs1kqJXQU6laoZuHBe
CSNTCjA26k+Ual7NQV+Izld1DXTcS9Urg/6iDsTc9dQmarKouior/IEzQ/gbUWQR
8L+VomjGUR0IVhwBxAs0qQP06RTnBX09/G1v4qgRYWFb+3My0eyhINT3XIqy08K0
iyngftLAfQ8Q3a+WxyKJ7QpIksBx5G+TKZM/hV60ZWZAHbKKxq9skCKoQBTnLk7v
L7n4el26MQAs2hcSyKhmkS20d/DpDGlZIkP1sR+vcgn2LGgy0IJyJhGP3DcwLFoz
aFkm4TMh3kqYJGie7iGDpdQAQEesxYNSjRNAaUXrf9Heh/qsGQemHdUL7C40IldA
RVjWkPmQYxcN3QPDdT9bJ5bTJ0CfxTNfSFMtalWPVIagHJneh37qrsWfY5vzJ5sh
N3RM1BWOHmCgzc1wUNvM7qujcj28TmrbYwOr7fQtH0gk4Pv/Dm+DCEQh0UdzzB9b
p22wyCKoqJBlbQL9Y3jKnwSa1fR6hWlUcX1eS7L+GYWlt+sg9a1Nr7Hm2v3u20Ur
B0NTQCzGUWRxQYKEr6tSs+GFGb6RcWE7dIJmvP3jxuMWIaQ4/zPQNPHyfJ0WRYvL
reKZO2iTW2rzFW+2FXXhyr9xK6tVsDbBJr5ydMuTgQUF1nCtgtU3oy744M5blC4Z
MNMymXgkQ47psyySZWFOm60M7rxMmVLbfpxZanCrXYJd/dxJ1HPxAHQgR/Un43EP
Mvk1yRWOQnY4VGhbafvIfSZbZrCZQDdmU+YcnC9FhoVxAfr0xrU4FXZwjbsiLYh2
gl2jdTCBhR42F3wOFP4Dk94fCMwbHGHKdG8FXgGKod70jnsp3Kqm7wy4MHVd7QXs
A736XiZ1ELWL4MXdGvgfRObDYFp475J1J3QYPA8Z/W7U1i7nF0RF8f9tbozKJB2F
LS8c3HiPrGw5+qywYinpE/MU1orYU0Z3vOLqJqQ4/0tF55EOQoIPEyT26JTSMNpq
GSmDKyP1iHsOKT/rwovd0pij+I2mr4XH7kz6S7mW+jjm7O/yOlSBGDFilRD8dojz
x0XhDD/qTu6b2MNNi4l71+lT0eKzS4oMwb/Cp6guHDJaDTiPOdsv7xzfUrk3Tj4g
7XrbNIebKVlXl8ctkeVlUeKQALYgP8Lnf1ZoX1x8sbRWFfmzVJY+Zu/wf44W+QKV
YNQIdSv4c8TtKhEKd7NARnxtpTIMngOioKaO5fjCNzbgPp6RkoTHMZFCWzd/Girn
g/YMVTdpoNqtcqBLqLiBsfmo7ddWlqgVXChwy4N6aWibpcTd2R6q90+JccFXgwZ2
YWnJR04RdPnwE+WcKjBgCjDdd0K0/HSof1mNENeQNXJUqyvbLvlYccswkH5tYtpu
/5Hi5+kDHR8uL4Snn87AMyJM0YFI9yB8KPYDBLqDpYih/S7nm50xhRYXQs4NG1ss
bu+82ON9HMTJwtQfho9cKMBmxz1x28dxOmkJGrt0RuTUH2edmvyCmLUhxT4zxnZQ
ewnu46/S7O60Wvbk6d85F/NkRjKeHeQIQUdD/w2ZTkFAemuuAI0aWMHfX3+8B4iC
VDiXDaAMPDql0xPZ+tJkcTf4HjqcvV4THziN8vZykduCtf5KjqOlQTkmilV6OYO0
Wbdn20HR10uxRDCdkNY6+YGrPaMbdM72TgTqLgqnqQYQ1DWr8fUZbQeuDHwBi8F/
p9dq86VVuFxnz4Osw0LAWmiEYYF5S+yWcNBf9Uz+1W5RHufpmdVgEdj6Dv/WURlk
ok0XqCG+m+mWSGy6NjPUmOpmIB6RQcFr+IQR+T5sQ9tFRi//wKdti1ZPZIsKAQ7+
VdtbViVDJUL9eTWjWpHcxFEKg2pr0HLTl8JAxEVQPg9nIUq8KEkfKDF05RXqGmZY
1Wmqlpe2CrTR2hLZAujgAs5yYff2PF0pfYCRCNuYpKKFOkeHU0b+Qt0T/X3yKojX
e8xE1O2VAG7s1oOedwocB0wE8CPcfizxaSkJPwUTfQFARbr6An8BjVTX6dYGNcTN
G8CYD+fLcB5Ck5bvE1q85drEmfpOqA6o6R3y37IFyX0LORSG6RnIYGDkzmoN910g
GZLdMpJUODQ7IBFSLCPmWD4v1/93QE8oz/izhwrwbxRjZzDGFEXEyIMtHuMn39p+
pgZpAsIYjJJlnkmor0muJ9vkTuFc5Sp9Fn2Ni51zvkJLk05DHwpC9mX7aSarihY7
NSNo12F8NfP+wHvvpg0AX40FSETak0jzgDPb4hvdOvnvyvSdGdtJOtkfspwiDl4r
L7KpZ4lxCUiQT+w5vd8DI1k8AYyoEKqJLhBrDcrgfKeetjmv6BtLcGsldIrRcyon
7dpApgVkjuuOxj6IngJeIac9x7pJNgkieVOePHErd9LkpcF9O0jLsGjC+/SaQZhd
czORuuC4q94EBJystKz2E00ZGGr77TmLWeNx2zSjuUdzp9IqKA/lDDeIIROG2O8k
xU7oHxlPsUuVimLkgwvw1aIWQgldORWQD2s0a1th7RFiqZSmUIvFMJvWo0R/KUet
TVntSSivf+LMI1cYvHZuAq9XvRQJH4jI4r037AeTxgjMf0XE2HNmWoE2GWJ5660J
rbuN0C1is+LZaPlIUCG6BFuBQriMZqiv4Yp2TH7lhyxbbkhOU36Z/hCQyXHt/rcF
H1BbgPQ5HBgQdpduZKNoZMxQePQgdIDPHOluqsZBenniVnzPeQ1Qjz0RFbMAZeuJ
UomjVDN9cE8F28/YqMRjtHMwxEmoTxy0VWIdr3oGqMgy3jpmmGBqAPI6rNLGSgm9
RtD3VJsOvm22dLchhT8gl//lVg8K+lZ1H+VRZCq4zUMz8EObqnpKhAEo94jxqJ2O
D4GmBkKqJwESjltrNZfE6QqXkE/Sai3GMaN23msaJZYuQFDqIsNbJ3P0yvCOYK+D
qocnVZgyfGGT72CRm/yHDzEeDu3yVdCXidd4eHdmaF+0ZssbarJrJn9ONcj1FzQT
JQdAj2qbGPq6776dAvGiU7DeoRTinTSwatiFK8qh6fWPXndmhWQI1dlx/LkgNdJ3
a5kCwJDdUeIU7VBbBhlicUPFr9MowkYAUjUtyaOsuJzPsDLfJYaU2r9uIBjgwO2Q
wrZEpnT4cllEJq4EdwS9FVHLjFnVm2QuqdEGvmKCj0dUOorDZ+g0cl4ilzKX6Err
7yhZcQyYoFf73eTTZq+DrBAMw6x5ajfh86Hw7USkfUJmH9YhheeY7am3LlD6xFkQ
AInu3EIKk/8EHGDBWseJv76U6j0R49xW/UiXGq3S6tzQT9vJPTbjqAhRANBTM+2o
jUd2EWsurcC/6xL/2pPfkvafzudiauT2njzofW3NcW1hARk0o8k905/3wEoqE75g
jL85xPwALmsryyDR4ZRRGIOONSy5WaQ2sOKy7tBYZ8iCHCu0WAnvWUDl+Lyi2A9X
Vi2j1b6mwSCYO4bgTlEY722ee3RLf+Ebf4Of/2yUAUjQc9gJMGiuQrKA+ATeQlSz
5WQby4ys5amjpmewhp8DCey7DwaSe9VFfcX9rEOnwdi1Mjm0XY3KDJ+6xNAX0tn6
Sij0LlUasHjltE6Gs07BYXfb/8jIWGisX3gSA07Fz3J/+J9d63cuBT/m1YMlaRjY
c/Yv6qT7FQtS3UMX19nHiTukZY0wqDG1PCfke1gl2TZdqDP79lKvMM5IKYxPDF4F
UMCFFdOfgEMDABCj8Qu1QPFG5gO8Et8bHRNZkDkXVRj60/og976q2DO4cVqib73M
bhJsFOSyMEgh/FrK83S6eYRETXPWBrgVp6zTj8uhm4DHN34dZsZ8hfuEjyz+VD9R
Oyp18VqJuVSX/Rh1/3gFzovVw1NLgrGN/DdqpOn1aVY+EqoneLsELPPg/PyE9/SP
YvAPTkK/Pa3R8smy8U2fBCeiQQFIkbftYlpFlJecl8uTUIESXHOl41JZBL85uoj8
osMgZOeTYf2Z24Or37hlw35mnYFp1sdTcVD3xW4UHVDh/YKEcv8IZVi0+qfdu92I
/Al7N3HACUSyGtA43SKLuYy/mSKHoBf44p7BjCPO3t0r8wGedqcgdw8+jaH4HQ53
AktWdvM17m6a3mh0gOtR75Aymr4/U6lcqs9tG+3uYKXcIgvzafIPCKhEdEwJBCnF
xerwL9XltyZcqmtmWogRfpDSuAxBWBqLsgPBdeMXipezqZCM2AB2oGrwXg8yupo6
/ARJNhW/F1B10wUay/ui5KwMGA39H+7b1PGZzbHdQEMZ/Y8xXXoYNlsdDP5XbL1T
NbJNxxwQkZhV7JG4Wsp7qccWkZQUz+13zXUxgobEgDn9FLniKPHp0Bin3W2pEAW8
NbZ8CAMElV4V0vlNTOy221OChebtKQD/jupUNpeSL1vq/bTKJS5mm/eIrFo5urCA
dJ6EETiW+piWkczkR6t2KxmnQNdOKlcPhBtaCHOmkm7aSytxFkCqHRFSWyQ1FCgO
Zks2MfTjVZaff/MlybJ8/Rm+M7iuLNntmzdmGyoaRJ6t04k6GaVc/aXHqiMMduBC
KoWEiOFHUreGYNWXrELOyFl3p+6JEGMCp/S5PhoJmGkDWvSco0LZG2TALU3lCIIS
k4kZfig93tX8rpgsiNVxy875yz//ki6Njbkdtp/wE0HjmWqpYQbkbZKphcGCjUXB
qBPmP854/fjdrrOJ/a4LGLUBxdlZlGNnyYx03nbNQxxBwWKT9zbecCzXS9JeZ2CP
YuH1ywZaTuvd3CZyKyL9R8xI7u0mxpTjBbANrJpUsgFcVs3HpcZpaOXKq8f5zOXg
ZpMhr7+hA4yoNdfxCTR/U4/T1Tbtp5EUN6wFDO0fqbLqnE2LWQQesxRm6klxQLn6
bIHSctVx2ijCjsWtA/YHfFQs7EebrzRrLQhiRpa2b+mRDTLhC2OMZp5E5e1VqOjo
gG+WH02CAmqDr4Uc7ZQJ71F2sUu9MutMf3oFLdO/F4BabjTFUj9wYQG5PXURPVGx
h4Xu1/UqJBQNIdQ9gGH7J4zhTGS8kdzRF+2iwFvGP28WnWsOl8lZsA6AG/48U/ar
e++ibUA3qK8lN6xGYDkjONFLmkLQxoR0DKSQuSPSZcj+Mj8APAPnjodxDsH1qobs
FXSuu8pTJnVF8v87mx6nfU+vAK/iRqKvAgqT3Y9eGsdGXdkkQ1XlvWDsI0pV0Vzi
HHxFdlmJlNhNV7eaXamnMIgOg8zK6xyG+aCbgl4IIkjNP0F9/rvRDvv3sqB0Q8tg
FwsCtTJncJwqUCTUm77CkOogMp3upbbxmYNgu38AEG9mwfbZIfJU8bbVAufgs099
EwjsfbGN3fCMtMpgErE15Myw4QaD5ocFt+hY0T5e7yy8l+yW8yqqXkFfirdsMKBu
y463+69pwzwrPp0zTQ+yUcM+RNLFFB0XQRuvN22XvLKfOVuBKJLicdiCu5gP5JDL
Wtkf7enkj9dr9tOtWKTVaDDHpUrZ5WOAG4mcPP9WZvfzN+2t3D0tSC3zw/Oy0nox
fWD8Cg/mwKyTHk2Adz6QYoXmqwSNoo3TrZPzYAgdLx311qoPntYj277C7O3u6S2x
QvPj9dmMjX1j3P8+/GZdXMxoq9DFtvDSRq8D/POhZw30cMerIKn/p3MUqrsfSXS9
5N4AqGlRxDa8/23FQS2+2aq0PlznSd/YRk7y8Nji1TbinsYWuuAMUpmnMkPecAWA
0IEIj8IbL3aFiRSvEOtCfTFXIvmPJCIpOJQWzxWCqz5oR4l8y4wTE+Ue8lkIFmVo
Kaua5Tp7sHo7G+z6HoQ7W7dVhBM7cBNftruN9k+Di9Q+KFr0AAnfM6OOCBsUVrTe
75i/6o7I+LfoSJULy8YE+xI2BxFxpTXL4SW8GUuZapgbSNshcyaThkqqSG5DKUrh
JNnToDgE8g5fhNC5vRu3rwlQklEufEUKr5mW9Rw9xWyvFFA0XAIPgJVTfdLzcnUY
6ETamXMbhwlGJPB7MDp82ef8bywI1RRUbodOHAAT082cssCQuPkwSPUKhMHspGJp
Yhg2s2yDqZM7LqQJaVaVhEuQdBGgo6AH2UTUSHY4/lIU4XtPhGh95gVDechMYhk6
emHNVLf9myPR6UoVVpIbZbyRLtoEFjt+kq/Gsu/a6FdOBtyxKm3mQj3ztBCRRPeX
h2WtaoNquepstQPNnN5vmzcGdFNHhJdt6IJw53O6d945Md3wX8nI/GG2JqCzOHul
XajDCJKSJnTjTVEl0p+e5tCVDnfT0UJIe2YKtU3adSTP5roT2CL+PnY3U10N3BP4
rI0sUvOXyvlOafBZsSLJahIKHDy00ZW1mnotT7MoRUDZ+YOm6hbND2dweTw4YOFu
AAzwO3C0hRgSlaPjSJkb220CGSl16sNJUAcxI1I1aIIevqhLypFWw+cOCPOyz5IY
9t7f5Spf1GPA3ecqUEuVXBWH2cbplDlteWJpsGczQb0qHgUeb229qI6aNs1lEEtK
/KgwYxFCd7H1oGQp0Cd8DkZApyzsj+8p13dMuTJ1f9Uhxyzw4AGPNzs0dv1SJLLv
Xrs3Es4YVbe64eTjSaGcFhqnSiwiNfAN24EM4Wf3bl9Jbxi2QbulSW4iUaFtYDfx
Y0GGQwYIi1hZ5W6ZYeFsfE8b3TOq7Db1BWLVRTZ7hZEE32yDgK5iPSq87ctRVZ8D
8g7vDERqcWmO3ERuCmx7iO85keNiat0QGmtAZBjjDnVFvUW31JP2Ox1dEEr4YqBb
`protect END_PROTECTED
