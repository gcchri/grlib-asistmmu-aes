`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PY9fpMJ6B/2l6gVVfgHdHckM0LxAg8tlU1tZ4Uk4Fr99EphfmHAX+X6W4EjYyTHk
4inc14K2W6heQZyivWYefQdbBEDurPp6edU6n8wdhuyYBDQFaSPkClHXmAFLHu7W
ELJ+s3PzExxdxlPL8+fvKaxrMDpn+HL6zJRW6gPKrd6M7/4Pat0oHF3MDNCwYwss
/5/prdLmiPRgAXYrb5n9RFnjbkXBCWiFhUidWk2giF3mOx1De5rb9x22lefNz0FO
3Y9ZHvpDygN8FL73uc/iDmG1w01sNe2jX5k4lidXCPM=
`protect END_PROTECTED
