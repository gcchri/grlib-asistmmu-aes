`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fxFvdfc6p9PGKzL96lhN7qYjNQyGdZqdpHuLGaJ5GX3e3TIzcf/2muZvt262QGon
CaDKyxIqoDerxJhS/osI/RcIuJh09lXuadailCKVnburfk51rxbdECMsYuv8WBoZ
Dco1w2H4iKyE1H1FIHBagKgVVNt7eG4LCQCXgJDLyUHUETTpMxA9h2Jpo67YpyGn
ls/q860moT3v5Ji30+uZ5mBkRzsj3+2bL7lxNfS0odTfbb8/dOfrMSkesVUjce6X
2CWCApMC9TOV/ybTPmIUhFS7HWB8mYG8tWG9AS7kRLn6z+NQ1dDncztBloqDh/mI
wn0NY1d0t/Sxd5oQ2n9zbQIZAaPnoEqLXQsU9NT5dSS8m44A7/WLv2oJCajyRZPe
U+mRg+ENPRg6nloRhnMnFWLF4XJXplmxtNHexE+F28UZ8hLppuOuEGylPnqTvyoJ
818M+7fp1zUcBRBSr/446J0M8KAV62KfMMmL/nLdzeoiivIe838dcV8yoVlAgTR+
lM5BW3Y3/xE4sJng0HA15Cr/pYmZflK3Vt+yxTNkvBNXTNT5fkxJ2AsMOEEw2f+G
NJFnGapLIjnxqMzrgt7jGzpS5mXhIg2Y7bdDOF8nsKG+7vH4z6VeciYDkry22oYp
XlgZdST7t0Y5zjr7pY29AYdS8ej+37rJT803/zAFHnAAIZTjcnpgDDMadd1PHkra
RaNSoZyVylZVS5FwTZTMH/Ov9szNaSyLSJsEc85QpIH1zv7Nrs7SCwRh21OAY+8u
l1/Gda3ISY/mlp7Y9XvU77XD8NTFTt9Mxo98pwiRU0Jed4+FuKBjFMNoV4DD1u6l
OwEWDwjBCJ1/+9p7kouvXshKShUYG9t/7MiUZyb8ZNf/6AkSGE3+rFZ+TIaicbnA
L29qWj/9qtjV7Wbt7e2cXUx7R2TJMpVKOeisKa7STYezZRmRScIfZgFjq+hIn6yW
fOK7UUR8N4ac9KSCZ31rogsxHrJTLeAMqgT27NZ6/iM0Umxbk1Ij7a33OIY9nSk+
OdD2eZJEG+Jro2oxKadHD0JS1m9f3N18H6ZbwK4sigJ73brka614eWpwDPQPca2z
HyS5+hLo/nLRmjArOZ36/+95Tw3wrQUvqUYYSLOLyDhHpCHlhrm9S6csclNm7brb
N2KpE4a7rIEEuakZ4TOd9Pr0JDexCSpPeHfl0gLmSFVrXZnKkzTo1tJtq3PC8989
apaEsbSriudY9at3bVcCF6G6JRu588FwrTbBTctJeC+PCYCtJZJVHMR/McWoPd1b
Ox20CO1RswQL3t9x/x6/z+anmOQTsI1FKdanVTAgqezotvqWBj5igADhUL+88Ofm
UZ2slaYMHiwNr0Fa3bQnLSsSlHGEaYWYYH574rSccCbfBUhapJz/xG77xwVFbLCA
rpTC4B8c9P7ieHmk3J5vMvKRueATjjdTFyA41eGqA8+fzjlj25zaH3HVi+V2fizp
pGovyhLugFdkQ3OP3sms1FgvVErrh7rwdZ4/aCUibCjwOnI4Q/AKDCtNsKMnwSwI
EZmHoq215c+YX6n/5MLbU1WwYf9cR6/sYPMArmskLoBCNAauvS2A3aSN8Z96RK/V
ens7hGmZY3GzXdkBjA3G5Ridmti+ZFxVPHAPMASkdUTDdZ3wqlJ7lElopZ4A1OhZ
nnCmp1Dv/Qc4AsE40uD+khfa9kz0MtWl+LwSr51NlNY02UOxXxkvq52bnwFmXd1+
i5QYRMZUAhZszW5LqMNKk+9S6vqd/ofw00N16k/eBL8VilEhLz7L/qdqWo1dz9VO
CYrEt5zyGRTZllioU7cxoFO5ljOdOcEt6MJ480Y6vmT4OOtxsxiyH1iaTxImMz0c
wf81yoQFSidHdxgxqZeg13iA4QHDBp87JBfBAdrwyiuYZ2CXzq6lpY04Ne0X/1FY
M2+KtvQuJic0IHd4H16OMrzoVaQmESL8t9RuY6ou6Y38Qi+idtRDgRpJJFcwRL61
p9JEV9njktYvqNJTWr85CmrWRmD1XKaMcp9+mvUDAjZ/G6vmFTnpx+OsysdjM/fF
0C0jnFsxr/SOpGTLoutB0Q==
`protect END_PROTECTED
