`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7pqWgYdHF0NM+yBUHKqxiqaq28YGwpkCkguKyayoyMOPIrl2pWry0nc76+xoK/++
nBczUQSQ5MPvqhkldlPQj6TGhYEz0KYNI8HqYqawr9Uh3zqa1e81VtuQT/V3hDTM
wuCADj5lfkKGOaf+Ne1qWoetyNvhtKAR3GF1StBhYtJVS+kIjE/UuU8LeXbxHdFF
rkj1cHjJNiPaUmPe/t9sVoqO+04U4PSsZqNaNXRzntsBi8yxyJRf7/P0v/ppenf9
FXF59mxuxlDC3o+zwU2g1LKQJKJqjUy0hxOb3vfs4sWvi/h+M3HEo3jVDg8AjEIo
ED+81OUwFyb0AqWi6wreqoi4G1I/7SPwOXda6PiD0QgjSRtzhpYT703UAOmF28fW
S2Qoj7vZLJz/JgNT4y+WySTjZfbvZJkYo7iJG1QV95wpyhGpa0L0838MPwT3/giz
icXMLlMFenQuv7NwA8j4GnqKepUhii9WDm+/jpWv2zmhVoEm2v1GSl4xZ1Jw9Kyd
HaTEmq0D8EfkIPjRs7/o/kk3uH1sCE61vFW3N+hfLt/UujFbjFcX8cg4iTBhSdrn
T1uZcZa4DoE+GUWQAFvMTKNTWP9P1TZVdq7tuvS/fkI=
`protect END_PROTECTED
