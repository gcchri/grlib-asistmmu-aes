`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nz+EttNTP9JYxSqFX6NDww8zL9m/6AuqpE65QYis5MIEz83ilweFcDCbMhildOXY
YVZ8I6aA44djvJgyY7RRzbAdSUCPfma940dkm0Uyw+vBTAB64MU2TgAiXvaPF1qC
46zrY5d/1rkexeEh3K5dsyesBkAbouBD/aQFDKjY5YYNvAlGAit10Q988P3ClvmY
awERGTvJuwZzUh7D9XLn4Q9SqyjgeXXkVoGM2hO5EzyNOA8W5hgn2arqdKPlShmW
k0NrJKD0mGKfpkwrf8KURw==
`protect END_PROTECTED
