`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jQxU6DtK2zGGxaNkfjHehkKVOVbrVtNcSx5Sw7WyR1vS9HNltmN/XapZWu41nCN5
j2y4koJzriNK2g9XAVzMmgC+fq+yWxxIqDDRquDsUn18Yi2FHBWsnAG4ZGMLOuEo
jr47nvpAl+lwHfHFkkVERC8moVDeCKO3FcDyVYdf8MHkDtr8INMSFfw2BgXFNR+l
D5ZPEctRBfmPd5YgD/MJaw/e271yAbfm+3wjJGzdeR/xSk12d9oMbTZA2ncFNHpH
+8Z9jEhRMxENrfSvmH3GcmNWrMGLyVS1E+GlIfXWYGHXW/jP9X8njReaXVNAWspd
TP9r69UaCzP6HGsWeinto0Cpox5QngsIm4EQDGRQMCnP2r0HuBDl1eOqdiS6jtoc
CG9T3eRSOSZNlWBZDV2xbzEPELEbYc5Rle12US3Qr+I=
`protect END_PROTECTED
