`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WNAoiUV+7AqXNytrZDtPZ6cIkJsDCY7wIbyel6mZdtpjCWMAtaJ0R7vHA/PtcMyV
Ycevrm/eQmkkzvqovp4zIhzRcs777dScnGl52xdMexsi+ljXyWY+LfldH6DHV1fb
uTd5KRQ4K/M2cKfmlq9kTqc/XCus2/4Vr4m5zizB6ji6n6/ovjm5RKHbzCJIUUyH
v31Un9IWNZ8n0PS5fvc7y4iGFnO/IGXX7IJI4Tx/wetP2rLwseZTjSzpR05B4wgR
`protect END_PROTECTED
