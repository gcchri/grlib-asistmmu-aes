`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PZ0GQC0b+rmhuos1O3qsUtV9Kq+/O71KGm2LZGz0wJFFYW88LJGwblb6hfKYk2yB
AoN6L5FOml7UhGVI+CFUnB4JEtypDOqUyBtbdRChsUvDS3TWbH26wsSzSqpS/pgE
5PZXAagM8fRyrhRXFAjV78krxFVuZJQBVRqPhF+dPXjjiTQxvCxQd26hYxcItzLZ
KBcVQQQTfWyIPwnS9MsuqMnzBxxNZ8zLAth15yv/uyiLnn/W9MKh0tRI6clzpMK0
QuWwiDOI8AMkIWDb9QTzRYZ9m/KKWLxsokGgHTle72HRwOVdwZr6y6XwucdTIFP8
Ojw5NXQJrXAtW98RHstvDMUVjLrZe8JowMInXCv06J8q8RL0WoMb543Lzg52WuVq
lI/pnI01j/8NUQCINcft2ZtGyY7zztAPIs40pHyHVP7DsvAkcybrKpo/Q12EKw9g
fKBnlVyrlhUPyxH7i3oZ/RyIR5OxlQRpM/oCFLVp7FiUQodQo8Ib3q11CjF4ydAR
NtxpOi6MXAr+bDAA/8SKifWPcPHZdUyMOlGSsiztdpZVCv7ouBn+1SvKxZ2ERga1
wnaTjytTRwKRCNt42RGHPAGKgn0UkqPme9LjQ/z+OexfP7ezKA62/Zy9j97WcZPd
3JuATBjGeonEsAWxZrjEHQ==
`protect END_PROTECTED
