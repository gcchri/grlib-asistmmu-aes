`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o72wVyofHFLw4NKVcmjfINzzOrplkTOWYWHNhTUdIDYGDkebZXr5KoEMDv5zMD+r
gspngiygw0N4UGO+JmiIjteIiiIoxb9aF1he4gWoNol/h5xBNy0lkSPhNvxOYK3f
21zMgOhwEuDA2lCrnPS7kLu/ZRf7Lo8VqMAVoUaFOvTXDKYuT++9DGV40Q6wJRev
gpQbNgV3IdiowgdClEjdR8a8DfpQy5iyK6AzZcsnXivsn5mmkxdvfmkcHBgd6A5U
5PyOVPA9hnXHMes7R3C7WxRd1pSE2pacECNmhyKTPzdyeNVWcuVsZjqgKhF8y0Lb
z8uGRD+ko1MAaIf5jhNigqhLyUkWPAdAweKi5ASNVcaizWByVg5XP1ybo/ro6LUr
taga03cTIpyTnefHKnW7q4e/cMwd4pJgSsD6AhjA5ChsRCRzuIqj4/4+xbBjAIc8
UO9B4JStFWr0yEfphH4+mgsp7Q+48/K+M8ARgfVzRmIGkjgDdmviR1pf2z36uSYQ
XHyX74lHxdUUNz2W11PAj2WgeertMHuZhxEK2/o8UdxN8PxmAGIgtCYHQVkYrvTo
sa5e3yt9DYwbL0VlJR4kByfw/jfZvnl/QkEcUgffzPVfjyKpMIm+GNCRJje12Sua
X1aOneqbmoSw426eA4ABvxfpWB7CVbDoNpFnV85zC+Mu/1rxlrE5WRyNRBRx7O7w
EEP2y8V7dByWuOdR100fwVfK2mRWyJYkcULqptfTsJbeGx/uxjzDsOPQc5nVqJLe
wyE13+lO1XjXYlGiZluFbE+PNYduundmQVlT07alvxon9/DLz7FvGhueF8elmcSo
IPgX/BmPaRabUOkMxW0nKRbKdfJXEJ26F+2+azYqSgLy4vTofLyLqnJATAQj5tZK
BcSC/7MEBy9BxYGaePZqwg==
`protect END_PROTECTED
