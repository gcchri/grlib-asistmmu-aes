`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PCApxzgKn5+wfGl8VGL2pStfHziLMsTB7mTQ24rU5zMdN4aA9t4acFmgYY7qerLM
mmBQVP6t3zoUZSclzYo9z5hEITtOuQpc8VDPid0AcpLyWs6eEPTU7HxlcvflbXjV
u8TlpJ3JFe0qeFnCWrwkMSKuK788WhM/JJMbQlDVhAbRhzJBZVfCqRRc4y0ff/mH
Ji96D9m402YmzC6/ofpXqsVA9F/X2ven9Pfdk2mdtqpEHkTM7FEst6rbKBRWYZGy
o7zIQFy0g3C+abAx9MDDSh8c1V1KclkvC9Icp4v3P9QuNW+dLKGOYUB5ZIqBnQ5P
9U70DqbGxzgPn02Uthfhxeil2d11NZKmAE+nJY5HWlLathAcX38nVhWvPq74etTM
VRVGHeIm0Nz+6rmkQnF0axjaCzfiFtBaCEzGV4PbgRWa4ITIp4ojtIcZlUGVwi8P
82WPLMBjP9bXWZubpX31xllyiIgLECLvwSF7Kh30U9FWJrfdfUayNODfOiyeu34V
`protect END_PROTECTED
