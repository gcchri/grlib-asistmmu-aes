`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZgY95fXbK1e0rE9J2ntXNPS/+QqRtB+zd4EnOFJ4hZeR8w83HcB6yRCioMa7r3L1
KipSZmlB4QjFHfszOaKQWUMPdfPVolxD0f74eI5tObHHmGAXCeAWHodYI5fTL6LH
KDItr/7/nopwp8XBDwU/Z93sfgq6Xfj0i6yfqB1WeRxZQ3u7VJO4hxA6RjHjxeCZ
zVqUvG/jFoZz1ZIbHESP7cwojZ3Kt2jA+KMobEu7Eur8t+AeUWMvYfK9/S5Savv2
aqzU1NcYLDosioOmAMUlq5rCgrPnIdOjbR5CEpeNwH5Ck9XQkJpkLCAE2lsaqUgb
Vf6Mc3fpj+Ddnz+E1DxwRPDNwv/N6eDz9bcP/otRZMSRcfGhKnGbAfqVgxNBO+2Y
z4dBsdBbLTrhv+Pe4NxUVTOiahW/yGDDsMzFcGAsjW0vPE+wSjDFtlm45MT6PvAI
x9IsKOlPUqf0gxgHUzrmpRSI9AxBfWf0oVtL7SW7anYUXMvcB2KzkFxbbMPL24kB
ewe5dgf97INgIaKSDaiicBPRkrMFgGaLaYCmSPgY3zDj69/3iVUI3xzvcO1JYXro
c1mAfJyIvKGVjZVQeTqwO2RQfmlNU881P3lLZMeyjtCSIruP/dckQOUmeupHOHQP
yPecOab8yTO2GeBf9KQtoNuk66LDia7a1uHeB+KVCV1i0Irq/F625iEjCFq9lovO
8qkw5v/iBcoImsIOUOlBQr/Or3x27l2mrecT2YApUL6gwjm8OYTEOrThq0ii3LYN
UtC+HLiTELPTh0TwYvdy/mA4EmnQiHcgE5hG4ehfx6EaQGjUxqYtETNxzfTI36KT
TpVoYRlvEtXFiELZgu22g3RwZ6sfSpqca1CmcYyClVgg2/jrc/ZbU+jMuIVcEsH7
BL1bBNcHKIPgGsIj6VaUvJpAkuwhrHTG7CxOyBVNRsmEohj98iipG0rPc3D6kjir
D4hzd2Iny0DeSDPe/oIhz6Za8Xm/ZaVdQQGf0JvRE+BhdajP/gQM1dZaMPl/1y/P
reaLT+b9iPfFxBio0BreJw==
`protect END_PROTECTED
