`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sNwhLdQhT6n/dEaZySCS/bMNzFlKeYYwWwm2R9DQdB2RumSY9FfoPGV7NPPHY9Us
CUsdEaYEmtPh+FpyuxlknKClwqqpFoyqtWNaCopvj43Ta5cG4EVvVzs2IZ822DoV
3TRciB4kcLxUvPfI2OG/uwCRZ4ZeFQhLvRImPs9jLYm3PQ95mDw18RIdbmn4F1UR
/2MLj9KLc33zloBzxANjRRRxEAOfYubirilfViKL8vgayaMYjuKnCeZBdcBW8ezc
0lJKsQfh3LGBMTT/QoMNQ5iL0mfUtasAPBGV2IaYePM1MrpRo4ib7pOSKE8ltbmB
JrU4maCez6YpOXmNSgSqOkQcop9MFsVWcGjMH4b7xXtN9+tE62aNvBje3tmuBLxi
cBtXYhCE8deIgyOVprWy+DqwsnCyu1sSPq0RwvzU0ePyyqpM5Ja86n38uC57pBHk
DQ7HPOfrVBsQca9FiVjLSAX2HhYUFpsP61aV77fN9ZogV9mYlj55uYHsfIayikM0
zBJBMDnOBo7vratPERxh1ALGjlIcFQhsRfvcOjIF5f+A3XDqH1uXS0Mv4vSMm4JE
9IT1yXUETRZVnHOdFyBF6ElmzbJF5mAIgC3aX06Bnec6dv3Uu40ealSJ7ak1wJW9
TOKvfCsYPbebN85XaRqX9g==
`protect END_PROTECTED
