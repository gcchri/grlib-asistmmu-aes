`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vvYjF2qzB05bcGRsHxOyxqr6v/62J1QZNXHW3fFXIZBAsZ+B/JguIBCvtTs1xn4o
v6Fc9aD9BMIToMEQAzbMOt5b9DkwZSKtRVu1kXkWOt7J23fk3ta2iLr6rS7q+VoE
JDvB5A9KFE2Es0lpZJ0qpPMgqZoyiF1INd0PikUxFV7pdBm2mtDu26xLJD8awK15
liwj7/U16N5iBS603fDemao6U9U3vI3Afk91hJGaXvGiSrcpL3RUfvBkHZWQyoki
fQ91I6q2BgrNNClx7UstUHDjZVshTYfdAavqLHOkAZfvgyWxyni9TgELhXmJNrb7
Cuupf3JPoV/m2bZsjZg8UWEGHqyeR94+1RqSrnCl+lrYG2Zc4obSBZxDNWLKVhQL
LLxGogsEoIZqx7OPoQSYj/B7rGbvTHttGVRlqOUvR6Nfze6HNlWI9DnHVeXq/YVU
jnuZiORWOrM7Y0r7CJ/EG04I/jHAiaHnoVvFc2PBqqt+snCXhIACp9AvWG5Zabzw
W4M/kdq0kHna/tQEienmdRY2WH6JH52kwPrW7IZPLOGwBqHGd6w1IkR9/NDpj+GW
4v1QRoHisnfF0tS4wTLdbSxHnVWjz7Yy4Sel8IooEYLOWmuV9Te+En8uEbWrr40w
E0baVgB3nwIEMqhpGwckIiC/eLCAEArWbWLyXxGLfvvwWyvi70BnRTyLLXZQk8Mi
5y++pEBENkX6lqui6X5V6cUgTezIfVFQcnQAwoiD3YJ5+5i/CcWrU/sgC5meITsz
c6KW83Pqr2IcxPX0CWrmghTIiBEHx8S7vX9WSsMeU6N1yOOAwrbVc0sinBDpHoCB
rykbGzdiT3JZMJUeA8DeISW8QBqCV4D4FpxVF0WMnnR+jPLv/JoaQDijRy36b68g
pifWuqI7GRrxxRJ65PMXR5If9/myxEjsDfwFzXe+qoCkK7K7eJ1xZERdGMnzjFmw
PPzjl+OMXbA3TxL+Gq67U+1hEw7QbhLn8U6sV22Jo43p7kt6qSbluF7S19lgB2RS
X+D+u1merLNAfhtCJth8lmRIChk8HFogfL2F7WhzVj4sGJ37UX8pZ7jHt8XIiiHi
Q8p2K68W3t/4g533Rv9fmtb/j2/bmG30JD9AbdxWuqiROcxPzxU3v7hYZ63jzsqH
2SLM3voPxcaHwMB8Jwv9YDumx3z+2zvmjoBGh8xCoDmw6XQyb11995Bv0UFEOux8
Di8AraC9LbpOJ3cBSkxiSJIMkwoYyrMvmY+jRJAt0/yXJQ2PCPv/B3NLZGmH5BiR
c/u30gr7NQ9WX5xFDWgX6K5hnXv5kSLUgw8bnPkffYrK2XiplxBDiMyi1Nz/uRGb
Mh3hRZmRlY0rvRTjJ4n63FUjJfu2kG/joNtrUt9KX5p2pxpTCiHNv3CO91jAHSUu
GzHQMk2bgEIzLSqDIODh6xDRm5nTN3Q3/nybcRtDfPSGHzEKYKE0t6LdUIlb5zz/
LdUt+RqdAyofJWLtuYvwMRBfzHG5bbtx/UF0IrPkNNfMKZAMpZAC1JRKQrj3zvQs
T+vLtxRYk6Skcm5f8LF+aH/dqTEDq8N3z8D2ENvYPrX9e3o1uTTrx8XGnORyweAh
rOo1Mzq2xctyHQN9cBuJn5Ev1jQuhln4OIccVCVh40q9ioS8IpOTGqY6vMs5IN7y
v4t9PyovuMa1cHTA3TJaDTBVvD0mtRCx5vNizAUOqBgonjR8EVjjkqhnfZhyaQ3s
VZK68Cfj3O0J+84PR3nL+nQfkyNjCS4NluDOaIBBB8nYeGBvt6fEX3MAX6G06sns
NkLLlNzQtjB8wo8uX838qEFYCtNduU/DsFOGxJJGPa1oi67Wn4QPJBs7FT4w+Gcm
aRraJNke/NN6NCynVvYIE3HA0pTnj5KMdyOQhfP86M1XTq+GCwUTNABmGOVjcj0M
`protect END_PROTECTED
