`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mbpAMdefiPlZN7RLoYCQGHyrWg7+E5uhZGNCpXqhajBWtVZAIgDMR3z7OKGM/LY9
5Z6/EBE37DZfipmN96FhT+xJ2dwUQTbG6U4ML9heMzSlOM6cqBRyyt5H6a4TuTi9
LAlpKmVZO5uIhQUaWeyGCEIHP48NkAdAgTIOSDgVKWOxH9A1xSz8fMB2SElz0+fU
PLbDACj+qIHW40odZzfkuYR5FbyDY8ESQ9NsMKo74rz1qWwCjv7x8EhPEuwSmclZ
h3Bh9gUMnGIazAQDJb7P8pDY23xXvVzz4SkfatqI4jcN+Al8FpBsArjMzfds628m
RdzGm0dOu/4F8K509zasT7ETnxNkB2oo5gXz+IzdRiPfj+YuB+mny1fpADTEMQUf
`protect END_PROTECTED
