`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mpHIM7VWvEBgwIMZks0ujHvktMCEAEJLeG3TMcS30IYFcNr7GdrGL7bj1eJ7WUmr
UTgI3HM57+hrPK9Q2/5NLABWSJSjsLhr9EWpjWc4RmiXJqac2lspsSgQoqjFn04T
MODMTvPU38Z6dyejjr5A6kHzcXTYX+m4bl5i9HWnzg9PXVz2Kq4pDtY7qJFP4N32
/KWpu6wvGsIndXmspmubRAsfi8ISZFyzs4qcdZq/agly2Qa2s03XgjFkfayJXF6E
2BlSdLFOkRUmuo8t5td7OQ==
`protect END_PROTECTED
