`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JyvaidK5keTj9QHBvq/k2Q85CqR79AGLr+Cxs/NE/su6XIurMovcjAZ1KHgW56ab
6XlCEDiS/t97oMtzBcMFa4MwB8FntzWmjclb8Qs1Am6OK3r6eITJtNBhOK0Z3QJX
Wb/6BZH/pmVt8D7H1vxqNacnPnWKyMeCRyDNuESp/C1EQaOztW8PS6II4SG7YfQ0
wxyk+jmJ7k53gEa5upVgzeJVU22PXGaKPEayiP5miaNuynWhOPTNisd0nuQvf4Qn
pRXyAHDbnvyyzvsSQlxaq/BJofAV0KNDr4NuT0pkiXhe6LQ4Lv4ICmor3edghF3V
LYGF0i+oHJycE43VQDHlUPY7IdQ+8DZYOYvcZQi0OuHyZIXcqwxue8jL9aivL8Pl
76Ooth4iyMFi5vmBCWnciHQ/b5F/tmAGj7lnvoHOjrvKrO6A8T1OgigsAhaRAh8P
QLHiA0IcaWokJucNljvytdIj3g4Yx38lxer4SD9/oHO0Of/4+OxvGBqcwReLzgT5
no1UDqLP++9G4YF0eDEwQUE5D/+s2EuIgE1V2cjtgxYj/KZMVI27jKQjuHiTBxsa
SrOCHzdo2MofJgLWLhu1SzhcFejnb2TyDZqhQEwkHsYiJvnso76N09JvkXsfi3Tp
ttU4ecHpEfkzMSos3ykerWTKtlFJWVlplaljfodz1Tov7C2bHuyskOxjPxXzvMPm
UKrCy9FqlFRbplTBMofNYQ==
`protect END_PROTECTED
