`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
929I+CipeBlSz8j/WL+yNHMtXJZXdRo05EA+fP23g2QJOqYyVGII3vIXgyNyj5iC
fTCTBAlWrUzp9Yh8C2Jf7J5UfxMubltVoauH5pl6frLFFZ73OJkAOWyreW58mWp0
7H6kEEgNild/+bOIi5ASAjsM5sk6X+CFdSE5scXIWYsv8ywgnBSZVs8JfKOhzyzC
w0AncZ0qs6UDx6T1FOOP0i6Ug+qitcgVounv32Hs/tU4gaPfvLCgEaNMjJi+jN4s
JGR5ISa+P7koPP90e5y6CKWZ6u2LmaUjjRs+uGguJoF5pQKfQvOUBqtoQPFTK7FM
Gdx1cZn4gemnL9qCz5xsKJJWGOQJmoOBpRTSMPjoRUvMQkroErFz/jib7SO2E6Kx
txtU1QaNyjN0tTWue66vifVAuCrmYG+ttmpsaRjMqSjLrJmIb6iu1DnR/yK84l9I
oGcPGI+r5ErzGMdgprDZ5XavwoChrPDOG1BMu8XtsiXqHRg0Z7yyCt2suU+sUFGx
cyxTGNoAITufZ8hJfjbTY6cnof4vm1Tw0eNkYhAZ5qdrRMqcegzxAl+vRWIs8vzM
eQgGmWG6VC9ojWc1Ej2j9dxzTi+n2njGf5mL/rTsJO7xOMCi6676yYHKE1c91U/9
sYVhUScqORELfkmVQ/TzmF2ThHuoi/pED3kRPtaIp2vtPVvkzmyqrfdsY30a5U51
0DR/KrWLMUc1qiapltT/eoRGCGeROr6b8PMyhzDEdbN8V3QB/xs8DNWx6x+Dpuyn
+t0ZdOJIu+a8KnWgC3bk8XovChBmjk8ZTjOKs59zW+vOhY25sho28Ex4NNA1LL1S
TsgV+hFlYVZclSEgAtO5yiHQeOegqxgd6ozebwB73wsZA/lPmbtjnGAq6nb0ZvBR
O5DN6jI2q5lXS9yfClXdU/FIu28szc3txoqLEid83lnxOPMlkDgb4klDWvQOGAnq
af6VsFh/XIZv0quqeDbY23DcdI7MlDd4ndjOe71GTbqC2MOiNJHHHIOLgnSsipJt
3gd6Ambrkx721X0S5+F+trXO8sVDa/MP2BgGrBwGSYovFGA3PBqV3i9SvEstHWFr
EhkhSQTwTvcwL8c8eG4S0JUE56BVxXLm9yYTsQI96qXSYlmsDSpntCtOnS8Q7cYc
CntT5AI3zT4GsuWBLWdX3gkZajoSDf3vuZZPlI1RbUX2a6H2613mpo/qPbDd6VSi
LHoFGQ1r9V+nlkYZk5zMbGRIb+mJkr/QUsY4+KI6MCqVCCgAXmYTMi72IGTZl0Ev
Bp83009R6+U/VBDsrF/TtVd1Btlty/4HyUVsd30Hx6yH9AYUHgFdxyYkxTTzSHs0
nBGAa0UJHKoDedFgpjaPjvu+0tTi3dqBjqCWJ6MxMnCyZNlPDyg4939WPyqK5xwQ
tt221nfz3HYIXHkQ9Yr7wz1Vdz8NjJpg5N1VhvzABJ2a1wMU7a9yQ7qPlpNnH6Os
tfx4424O+osPDELgSudViBRAIpEiQEwa/30OeApCJz+d4qNpGFOB7jBsZUVUCaLp
mSZumf0RHiZNlEC569VCWqWMX8S1rahDbV/DsDPWXavRLbXk2QARMw90AAhHNs0K
EymA5kj8d5F23DpuN0/HJeMgSVO6Zp2nNmvUZod3S/iWtJydgKPzUujpHPtKiAvN
NDUU8G0oa7X6hhZrI4lczQ==
`protect END_PROTECTED
