`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dpsqgGi0Hi16bnZUGxcZGZYFG9hP313U9qAZjUOIoynpg0yt9NcQyIgeAfFg1b9K
spcMP96+I9+1x5B/m2RaIFTrO+kC0BHro7oer2ZiyAhC1Ox+C+SAs+5ct9iQytyS
0aHds12+17oidgZXCc0eg6N4h6PGIVF/hIEQb6INC7ssNGVdPGMbzYSWHZFmcC+o
VkBt4v+ARsmP93rRIVJcdpFPfuqsEtKyAYJEO6r27/UYUwvMJ/YhE/jn/VkS2Jp6
iKaXGdOJVHYsKNEVY6V9Q9V8fhgkM0H4qxlPoCu/a9t/Aydfi/EEm9EcalZdSJov
H40lO0S8AvanwzcKIj8TmHXE7da1Tzz8/L7tJ+YVMFsludJLlJAPcmdkxDZnjCo9
XJfFo2lzMyCVxLQBas3hcbCY6ChxAF0yd4LpcqemNRApwv5sH5KPMBKmLU7CCQav
VBlD43q9EmZc+yCvoXzTuvwAnCJXerhxyqs3vCHdrK0Dc5YKTq6W3XTotGIU8tM0
nuGC3VABCPDyMiTSqCMHM1D6GOtQDJi7t8DY5+V2svdr3Reh9W4k+nG4X7bnYSMp
+aRsCgr1sEadpI0emuI6aUFCUAXNXkicYQe1Wm1wpSPoUUMa9bvauCUq3I/sNVZS
9tg+PAzSFomjoYe1+YIi+IaERWPjhPhRLHh8SP9zqFzGB8V4/iraSt277wtOCQmQ
zYURpJsreiXl7+lzzRXZVbwx8IouvFORifVumeY0ABa7PQvlrANwXqCMvBOhMa9q
4LMkYu0LHi1GgFpNZNgU2TPtuDQAQeLa88dBgdUqqEGyV+I7eGs08f9WpZ7c5nW2
QW5ShhRq+r+xTc8sm7GiDNWn4tAvM54SWVYuc90tbpX/Xil78zDfARDEujqwxEPv
Xc9MmMxAmcAcCZ2LoesgAwatufJ1YnRP2wtAIKu/BYXV260cj+q3WgxMy/oKvmMS
H/8Jas/9t8y7E5gS35HKXe8PlzzsoylUgg8TAJItr7YbPe7T8paKKD78MLE3BnJu
8XdH46HvL/Hbg+MWHJuh7ghU8vjIBzMrGSBDKfMuOWtUB+UskDlJddAg2nyq4NJA
9hwqEv2Hf3gvvygthyJ6WSd+ahq4JrMROo2nLTKZC1GR4esbd1hJxRxeYW2H9q37
ACf/Crydm8beAfX0Ov2Mz4c/4uXAZVqwgAmFdAn11x0/v4aiDBSHtW8OYURpzcu1
CZcK9STpfuXbd6B/uyZRvUW9MISBgXaMoFNvtXNrICdnHD7j+/opoX1ZcDb6rv1A
NHYoSyWFd2LlryAjxD/WtVKuUxOCYgnLTEQ+OZgv9GALd/YNcrooXDXV59HoBBbR
o/0zTiQ0wwn2lhWTd0yoQpqegnkMyicyHjmjWJ00hB2ZI8GvU3vKC7Q9gberTA+D
j19SLvTchK4uPB+HRsPCBxc6ZmlrjWZp/qp4koVEK93U3YqyWEczDRCvnArC3Y0x
CDG54PCxXw8wGnkDRdCTygpuzb/C5ak46ph4/iePT0/UvLIvBikpccuv9ahJkpk1
+zy49bWW/v0LoP1PuDwFANl53diwLqhcFUTk9VYWbHTU5m2sQBI6GFIugTiMl8Z6
MW8JMCklgL6p8mkGYsOpsA5nD1i4pPkfw08ZGAydcIoKuHUTqFeZEDxUa6edoJUk
QpMOyjPiF0TApQU/SKVA7Viqa5LYKvbMvJO/MWPr6EXw06eUxi5qMc/auiDRscpx
TAFHbOIWyMU+sBkxVOGfy8mBgiDHc0bbuxgXYy762ad/4eFysi2OsWSWwAPzP6xK
K/T5/EMF4vwgRowWQng9QzrhVXmqhv+qa960zIj4QNWKwkwlOHQt/QJ0m8TV5QOq
d1WqbUfvqeZ63ggN2idwwdNEQbled3LVc9q1lvLXFSRey+P1mEe0mHh9jAmq5ogc
4m1WOiZC7OxeOfiEbGnPGrO8Jg5Ru4ZhKJzun83TpfFBpktpdSwkCziBc0wAtRNO
oI9yXbnwDHSCqpHtsb9TvdY/ii3cgdPDoVO01pmB/OI+VD+tQBN0+ihxDTS6mOQo
UO5ELZcRICevs3QQn4O8z2JwS7y/RIEpvu8bzekLz8o8uOjbfytRGXTMSD9eAsRx
73pdLpSOJZdo04wwtN8a2DQNV2SglaTjYMySHa9tmEAj5czEgWemMh10haSHhfMj
J04c6jErK5jOluY8RUxMqg==
`protect END_PROTECTED
