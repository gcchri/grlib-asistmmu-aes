`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZjhkenoD6nxF78Kdovr8JChXjuEVIZxvgKDXvnMV4p0YYBf8Lvj1eg8WjCZhzAnX
WlUv+/s/meGjkl0k0bBCexhHTh71WPD3OsANOMeqRVAYUwXDKyPf9QoXWUbP7Bim
ZayXvqf8tgqBMozxk/jPBoZkhjvG0Vzo60Vjz1oDKsaYir8lGW8KY12gwxSqxxBl
qt6kRtZatCGXwgcgL1ZDmJsSz624yCnmGjqFqB2nJgz3w1ykpZiO5Dip5OWt0h/c
sWxAX1H/3aKno61qcD6YWqmer9Q10xVWBdXb5EWB8Nk=
`protect END_PROTECTED
