`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sV8GCcZetTAYIPrAC2qjvqLjH3T5YtHI6JXd5i6Js//XdjIJIpOVffEqjJ9Kmde2
GDt0ZX4bBDmWZmLLIXDl6JWoWKAMshtQNYdcbhg9GohJUv5ltrV6aSlSNfKWzS6U
WtlUbJPBArxHaoLFW+3XTM0G2SiZNZET8QOWgzLzZX2BshNkOVYluLQRRbVcgpN0
1JlexPb3pVGEqHd3SWGpOnt/O7Qkaxw4+/5qBYnbPY6V0p8Of8kjd+QPxco7jrmO
cBvfLcW+qZ8trlEvLZUgIRXpM/CN3FU/yb5DZ33Y0uA4MpmCP4a+CbAo1BKknkla
i3vEQnIt4Y/NqAh/OpjsWpcT9F2wnOT/igQ/uuL+6WKSLItYTMMAEYNnfL3eDFnd
WPOX5gTG8qMuiJXXimNIvOvByQVSmF+aSpsL/huiaLEfl3gYrDWRNEVSAsKnnN7B
kC8Ogg5WVOMn1NMIWdhOaI4NlFTwSGq4yCRSPD3XBOUfaCuFK0YQbLOZthbYIRQ9
NGvl4D75U5k7K354u84XOQL+qX2h3R5vGE25Md6bEs+UwRJeEC9VHVN8b6YypCie
hc/9tJ0YDQRO8f7TL25yRIBp39fZTIwCQmG/Bt31pAjeMSUnfmQkECo50V1Mec/o
RRrIcjkaefqsofM4CAqlTkPpg9XZrD2DncaBIcgTutB3pVb/YX2+aKxyhwuQcko9
Oe2G4QcWeo3CHFbVm6kCXn8UdCwaapQ5T3pVpjR9SbirszWyygJk7ZbgRtAvFp8X
4sgPJ3ta2aXmeL2Bfl/yaOL0KSM/cOxw3eoFTxRJu2zGgwQ/DI3yvKz1s+EapsJi
0A0k4aPBx3/w5TezirDrN2fA2dl2Tpizq0gFqOhYFoFsC7kvP/qfzDEUHP6we9WT
Ajatui1ciRO1u+PGEw7RMrG0bGHvqSwi5OdNoGq/YRoe/I8lgRFrn1rv1HSC16LH
uqWrbxz2uV4jmp4r97olh1sYD7zghsz/T0LWdCJyGG5PLDLFBM2Intj9F3uNFfyh
tc/bUvvH69LDXcEN186eTUaSD12tj+WD+9BCb2aADIYyBuafpxFQeEYCUDczsXWu
EEj9bG3LfaAnLetB32IZ3+VdWbmxGZ9Rz8FLM81Hws82SW0jFV+zQVaBWX3vWYhd
19evICy9CrAHEokbOGuebCGpI01EOjRXTuG9fnZGQ+oFLfU6VbBvafHGWbPMWC07
H5xFTOhOL9fRypABLQwUHpMCcbWxq6yqnBpKpWZSl5pwWfvIfa1QtlbfjoMEvCZz
/xC9mKJDVrCfSr+ltMHLvlQsBJm7Px1o7El2iG0mwZ1K7jEmT8bXhW3MkGDik7j5
eFjlVQvnzhTKRPE/xXyjrlZW6ZjRIKgr3uZOLkzQCyzcuIoOWWEbs5hWcm5BHHyT
rPgkILqFNg4LquGj33I5VWCkmHHXGbV5XHDO1ZOwzH61NCFRPy5NYZyMJtxa0g53
VXadu5qhBbRNCp6xdA85MTfQ0AJvrfuyJ4RMBz+21PVB8GZQJWVa/BAni3Mr3/qc
1b7N7BKUB9edHvYYg2ce5ZPtCkR4+XrwPbxj2WRAW6NjhUZlwKi5xONyElPfJyHY
U8SY04eLrZr58IjWl+bD05F+7ijZlJILr4Xx/DgL7nlNPh0aFbBQ2jTbeBB+yNxV
muYOaX1JMu7jqwoxOEAP5tCKETDOQflHiRPrGGLY8+AkGoe2FOG19Hld7/N6I7Nz
/40iw0IX+m/hs8x5Fbe9WjTJpHDUL+/L0w8S/APIVa3D2sT/1Am+Bi5TLnY+Vx2L
hfhkeSHPNZ3cVv+0UrsLCswHG/IV2aM0+YXxfwEYJX4ADNOybcFDtUJjWXs++tVb
1WeSllmTwjO7XAmS2p9F9rhEA5VLmFjC5buKe3LjtWBDEOIh77DWwNvdQ+TBqK1y
+uUk/x4J138bn0AoJ+zMLFIM6+ijQHc/d99wifGfUbTHUvI27mjAAO7hQQStmLwK
AljLdRXFh4RSmC5gf1i4gMKTYM/ma0qx5PuqKXy25iPJbHdlsUFJsQomkbaqVDix
MbEPmnNGuU9RF7HlHlNzRnvLgXHCCk0EaSAYuvu7CdOUpGOtl1iuItpU/fHpvPJL
ie8bN/YPrWUcR3G+Jo78h1k7pzWeTUCmWCAluDsiuthB+qoqRDz7A2FpNrajoWKf
WAavoV13+r19sj0Zno7U7Rr/dR3UgugHufLWyrqnUgjVy4Mazg40BNURUV6lPgV5
yHKRlfqVcfz20xMcGAQUTGKA9fUFbYWUNG6xmtsqSElFixFQlfY4dM0eWplW76OD
sd2G4Y+iI4g+L7hzSMMXMh+ymaS7mae6AfhHS7wtkUWR7RLtkcsvZ7uKSVmya4Tb
Wpo92fNzt+DIKvsYrB/7Td4vt4t4vgX4qyw5empZVvIXZUM/38YQa4OEbIiQb7pV
nZEvW8dyDtXX4ba3T4t3y/PNlHpu7R96q+PjXVWc48eMEuofAMUpoMBx6HyQ7frg
t7JsyWvruMSQ6i3WZBxCNZQxLGtudP59FiI8XB75+C2S/+yrwX+Voi1VbOhwWN8A
uoQ4d7MzMIpIFp1F12C8RWeUVdcdLlfLWiWlX6Muf4JqBOwpD+KMLmzEhg0eOvyB
K74x6DtciMVu+a61fY8xy++ilwl/HsHIFqd/QLnQ+56dMB8KEedJsm4WxKeSLGA6
Sb3z4F6SsCbN3WfGk6YNEeuzw90JsQJyer/vv/KY3mehBOfdwfx0AFPBGlXj5YDA
A+plHQ/MNCm1uIVsv5QjxckjfeKhI/ZA4foO6gpCwe/UvJbsJKN7mkAFctUXjStX
n5IzBCcRSOT9khBNug8ZFN1ZP/migUK2+9uKMGFSJNfelWJ5Ll/h3ljR3zWaflCq
Mvnp1NbP5FPVj9TXCAszwoTw1Yez9tZVVAfZI5Q/WXOYWgh7DkoZAps5u7Z7qSDt
Tl7CBLymVu1ZBdPw1F95QWvLPz1TPINMiFzynxRawe3adzyRetaZiqj8Pl0lc6pT
48IovztdbaErqhEGpMXM71rjQ8RmNT/iup7S/ehkE+gpgrPxRqyt4/U/DD3rafDt
chs04wy/obhJr41pQAKFkvrmkBhczKSCfPyBrFQCK/r7oybGiYQjAd8cRkduhVPV
IDvYKRvBVblfmXtx4Cv4qiHokn8BlgN3ILdqX7lhxPhMkmu8Ki749zZQUPzZxW9v
ZbzRE1PjESAV6Mr6Oyibaml6uonfn7PrJj78an703YYX6k2hqSIHtE3GGjg5ROGn
XyI2rWD4/hkAO/DTSqyrh/a19iQDuQWmZVfiwYkg5Y4P2O4CoKVx7bcYDJjvnK2o
3yxxvMHl9mReVfNf8vX7RasB+eJm+QjK5vAa/aBN2jR5W6H29dkwScpif2WO+/9i
9ML33cOg9SUVJHqDXkVgvKMh6pdNl+EuizKLIP4hpNE+VD5HHrLeER1ejkTiQ5X1
evDlRd3vOh777qrh5eKQjxTaU2eXXXthXITS9yXbsr3c/U8JRuXThBTXf9i8C/Tw
Fvmtht6Aj2BwXVUq3Lj6ziEb+YulCCS9BdkhSWQehk6J77l1tqcqkhbOdkbT7+xv
FQxnK4vFzbQR3LDWtn+znNx1TlVEHmRrMPrOc3c9rVcdtV/7GEKN2ckjBlOSPluH
+rBnWU9avK/o5Fo2d5o1aYVmD/6HaLsMIvwga/H35HMgxzwjWjQ5d1cqHNZpKjx6
sKtdBLK60yHPHyzipo79M5SQwYPbH0Cr8u+ZjaE1oi3UPULyYF0qvbORDVJ2ybnX
CzB9uzBwWWx11a3NBR0qyTgvtHToj9VVHZptHGL52eEFU732g++fI526PVbl9B/P
GgxJj+kavtqMbY8UW5R8Tyzgnrpr7SfsIiGxdYYbm7JVsucKUKk+xuJSytEje69z
54wG7JlDpz/gxw87NvcCjhbQZXyzpM4uK235Z04ocsEV9wwFi6JQP1xbENyCCIHr
cLsfHiRInir+n726/RnOLzPzzqiWUS6qED3eULiUVvNImaOUcOc6MSQ1ORxqMMMU
D80uBLp7499Pnr3vPG4hqAsOBrXGDummTGW6qAlMEmq9VZdLWYgvvtjrVcE1mLB5
f1HTviTHMuYsvIOf6yU04c+kfLZJoQAWR8lS+PYjJ+bV2pkbUIK8+Q5iCWBSokJM
ygWJEu3Ea8LPiXAcY0P9+bJGTxBTchLTu2pNkIDT4WfBknScWcyhD6BV1+jmDXes
lD5fQfYIvZ4lzj9WEDnuW0Yftbcb/WWT1YF3qds8GzDELf4vtCeDATtcPFBJnvC7
VziDQjLlmH0n3SZ0t7ITWAhJdpduLPONEduIhD7viOVYqRzxXUuK1CNKsGRSotsk
t/2tnBB9rhWTGUUNR+4dqscpEGI2nap8GIxoXGKeVsP2/Mg9cgiWB3H89XofsiNe
vkp0D/ID+0eZzGAhE1BBoRbxGpNNwkdAkUyIMHyC66q+UumcF9DB9UKb6vj+7K+K
yKgRLXAq8Gc/IJQaarGW1kai4BRbN3SEzhvu/aXhZYge9h/hGJySziCxA6eQHxBS
j+tYek7FGuZdx6K8CO9SbXo7Wx7Glucqo73caRN3rQzg7nqcXmusz4Q6okcJV2u+
lSgdToGhmVkLSwerNpNNzNwN30e61eECb9a1/+W3GrvRecOJqFmheAAfvLQ7kWV1
V1hGBMIqsxaNvBEObKO6sZrvJ1F7QDBu0WBeLRgokBZW99dpcEIdJhNx71rcyZLl
pnDzbT44IFZXMtl21VRKZ95ZtvpyZbn7P0CTYHUS60XF39Bf20m//jxJNnKa6Xre
8cDO9DuztluWeaGwMnjwM/pd9P2OuKE86oWHS1/jMj43myHCYSh6sODAeFLDFLN9
0M0r+4MeStVhlKtfg0+rW1meqhX4bTmr2mH1dhT5kfVI1J6OYausNWJWzKf+iGtB
nzQQBoh3AVS74tITP5DgAuo6ujXZm0SSY12+7EysbzwXHnIQ5ff8ANOb4e1FY3LE
waYZj+VG5VvvgWd1d9Q84NkXehBX79/aBoqeqB9SC7zntLwJ8SntGRcXxUyJT6hF
52iMzx5FlGvlHxm0Du5AelQ43fKABc9o4/M85Mb2CXq6FyX7TUdw6AfTXoKJk2rk
tNETuaeFW12PhTsJ7IZSY2bn4b8NLBZh0XkLSHHvBiCu8Tcy7mTNO0Vs0nwp/fQE
+I+PYUA831AeK/07bhklGQ7rOD4DOwRbgM9E+WewaXqfyjOX+EM+h3T5Whnoyq/p
Qia8hjEuTKp9IzNFcVJK36FrkR73RRX6+TSCh9XiAb4q6qDufNWuEX2ycV1Y0kb5
dZZOM+ap6IoHAoAc3VjI8Z2nCDzHf79bhuXXdbzWcuxatheNgJjwxj4V+/v7OcA6
A93L/2yGs3QkjCA5laSUohJzVAwV5PurO4LjNzPRnTWoYAtfmH1MwyywWf2z4DFf
8EGFtv0ULw+eO4bd5KA3pGqN0MO5Bzx7tDfh0mSAY3l57dGuj68qudZxkak2gm85
T7/QOoTMR9eeeVfuyuJsV3U0ulOehAXbV2T/1zR9q8aL2t0t7ho6c7JRYWFHhMz8
eluiyJDPH4BPLFMvYkZlYGVeRWIsvWPbfiM03eRAVj6MMroNmrOGncNlAuzB5knK
OApo6hWpSm+4vZaYRTUtJrSXzU3w95qarYHJI7onFZk6e8E17nOF8UvUQVQOZ2p1
9kyAatFIulxGXyzhFS3E2tpDfjZMMQen0Gtxx56cjrX+r9qIa0B57bGTyiqB07hN
y3BdDxaVRsHlyeWnof//skouHBEE6PtMvQcqjaEpMaCTNQN2JDaKwMJyfzM8zMfv
2rO8oiSmmK8L3kAV70KYED7UAOJWiscZ1iXTEGxZ6C86ulYafNDt7nGmX1MlrG3Z
98yutv9OXNuKD+sfcHFzZjZj+9Y8Pvyh6lL9Ui3+vFhsT6hAxB9zob3r7/xMDlHm
M5q3iPqE+xtOxM02RKg0HqRpVAwVq2a3fjbuanuSo9MTUkKa2rg1NKIMD8r4invs
6HayRszzs6Lf8EmfdwcwczX7KGRBV0xcCnvJ3CnnGSYPkVRftmnNHY8yESZfzhFb
426abiEQlrNBs73erxxRXvHUqIT0+zxZ9TRKlr9RvS5LndwnrR9nnN9jvO1eL2H/
o5kWahNuYGbm+wtfjq9WDi67bC4tY7CVu54ZyfsCdhRaxH+/LfoRHCWi2C/3MTBO
Nt+5B+gNfK4dYVZurKYRyYnSvPWEqXmUAy7/UwC7Sz4vapvQzTMDXGFP61LLz17b
Sg/+1sxDC++bWniAy3Xw17/yXotSHMwntloFx5oKN+01hMcxbrBWAvCbIGvTxLjR
MhurjLT9fXA4teNzxvwjYI7JdNDYz4RBps2sya6hnwek5cRDFW923LPBBaxIb4jy
BE3OcUgOjhFbsUtD7eePEamcqepYdPfe7kxZmFQBhXT1oO9+T40Hmo31+shj0xzP
RQfVqtTTBDFE9o191EeWd5iQRudmdvACBuQksOIWdnFQ3e2v4jAzaWBFN2s4g5cx
9gRhxyVCKXkZSNV7w5jFAXB8/YMVYosTglbveGpj3/ZnPZF0nvvWPJegXOyjQdg4
OXBm4h8xhtZh3dUyjArvdOadubCiGuUSmvgSIJAowQC+FYgiDr7ZRhDPmvOmLWj4
ByNIGtRTj2oQ1ofwaih8e7Hz55I08PSYoxzKms+MQy5MQYdqkduqZ17W3xcL4S5g
pE9EadtRCG8npS+RCsL+LdkecpDcRtRxGftcQNv9MS7VwGwDFijGQ1OyLvQX+5Fr
hFtiZzJOrvkCC2SRx0u1n6T4tzJjqd+d/Kvjk5BXoywRKSLP9leevtT1r5vtxL2Z
t/cHfuZQ/WNVXsulHe9MIOny6nlUQbmvwG+x4UdCHmfTvNnolwEXeDxwE1rsMwLX
0KTO1K3ErISlpDdUVM0GeFtJe2+NoAQv3feHXtTTmSYRhKuH10mrOQUtQNFgjOQD
sdm6imc8kItva1Iiq7vULWn93AlbIb2wWgxr/BXmBfvmRqNax33mJUaV+ek+OqLr
2cC8UAuA7wKW8jxpbQTjh0Ok7lreZAKBdWEgPgBfwcP8qwoLlCWG9jFz4wvJGn9F
9uklMxZjyBHP0EDarlGjZOxsnsIl4nCV1rfCUPgUmCECNRm7QnXUNrqE1yvRWlHM
E6Su9jvvYhxmLnaMPq4u3Dlr89ezNV3ZIFmJur26khKkzYkBiSbR/10978AryPUI
8zDkeeqYVCBjmpk0FExr0du59s6Oboh3MWZuZnNoUPp2qRcHDZpw1/MpBo/0uY6A
DgSYS9ZrogdjFnV+Olm2mhrBmnCtOHJYEoYkaor4qOB6sSgpn9PazaCUQ6wMan/f
9WDLdx3QgUDjTa1Or+r0GiPuEHGZrdlLT7UDWw5RRgiIo267jwIzvLcIAbjH4yqf
mwg9NkGGLymCXoA+xgCWhKMLoFf1l3soxlywRJb9a0+GLFi3jxXWMjAiIAOH1dj1
SbVENHiJ1giiVn4Ue2GMF5Wt5Zk+VRYJJljz9Dv4305hQ6yKLxs0jUnSFpy2zxBU
J5d7ilWGgd9eF4WzznM+Lxoii6F010dlQ6zGzEOFQ8ap6+itRP23M4HZg9/C04Zk
U7bzP2TQd1Hqj8he2Zx+nInBhE0FzMeGyvWK0oSyVtuYL+zyagP6uBwnumiSTIZz
bK5bSVKEij7pnSK2z5onzZ3FCMvZz6raCqQi7GtQMYbld2wGnED/xZdLr1v52dHL
OWlpFabn00aPyu40sOuSBtnQ7PyRxN5FD5VdkLSF3ghGf4tV+vV43StxvCoyf7L5
fSbyNPLU8geOCYz+/YEpipJBQ3NJB505x4gQfb2q6gCNvTWeE3IXZGdx0PH0GiV/
I0Ak639vIEaZd8t9zUwG+O7swRjzIhUpu3dL8t4ao3A+MZd9evdt+0nSf4xEejCb
F3vxVJ+Sgc3kRyD+ySDydyoBJO6RIWajoAVOXJqO8o2rm2PbhuGqeOTWtLqjfAdB
DeKrfHUtl4ZUc98iK7p00RDD0UdVg7IDHnOUZG84yyIamhO3QPdVj9WGOvh9J6SN
CKXinMXqtbWhazURY2CDmslMJ20v74+87tVzW/pqJ8sKpQCClHlWIsx03x1L1W9x
RQwR1jyALrHy4LRn51fcfNJLGLfc4WN6JxZL2RdnpKxTy4OfBkVO9t193gHPvTz+
z1OI5ruy3l3wDGds9IINbHQ424fVCNF8+HFN5eQFESqst5eGfGcmFLg92DBn/VZO
kWYBCnxqh68+tBw2o0FxFzOvPZFVxm1FtwNN5ApBs9cPWUGNX8qAl1meHv5y5Y7G
kctZxAZMDu8TP3DwMkX4YdvxT4SBhrJAreyc9yfmSzTLArHAjshZqW2UOvlA0+dA
/JzXVeWBPNxgqg7gR5SLPfXjXLKqo29Yx/qvX+EqoauCHELbATVxsQWoyF8a27qa
5fYmVmCXvfc7hn8gzliBkYqfqyJMsTEKTe5AMmCt379vV28unVKHoKPjv0jTl+7H
`protect END_PROTECTED
