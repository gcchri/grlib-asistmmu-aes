`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OBeLnOeeg99/YohbKUxsO0P7cYRN8gHOWuATr0bD1wJ2je90wGRkO8+6jOnlNYDy
9pVIwWWCzrMkBdlZF2xhUUr5LaxRBK/FwashU3htcOrxkym5EiWVMIWXhnCNHyQr
TaFH1HHcyfeDNBED7HD8Xs/D99eeICBCQZo5RP7bsN3O4s9n39BLqW6ZAkWmxT6L
/tEekfPYZOds9auX6gytlNreiSCrMf5OcR4qo4C/b20+Vx3aY+QhOrXe8WyGp68a
dSDnwFGwLcfgvnPUqMUiqUZ9oRlaHmtI9iMsMmVln2n18jl4TscEVGqfkhqqFRBz
1e51T4jdLv+Bcb9txzD+S3jC/d0tBwRna/Py/0h6IEw=
`protect END_PROTECTED
