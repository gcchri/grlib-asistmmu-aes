`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nHGEvvVIqFd4hO3O1LGr+ROger5aGagvqo62oWsIMvppSxhIWHTGZIZdrFBXyb5u
Xxp6LEgaomVV0d4OOy/EldUvIQP1s806WjMn0k0+8atOv7StCH90+jmZOk9QCnHy
7GcZF61lMJc65j4O2xznFTDyPkXhv+md1hCSv8RGYhBimS+f9YmQYt6uQ+GhbCmy
hgfCbKOwD9Pg2x47tenMyBGzZNIyQRlsHoMGMxwxL86BZCzlCWEyFbOa/Kr3ywC1
LIW0DrKNlisM0jpMXatgKjB4q/gkVIHOhVZj5Qtv6WufGtRJ9QSaHQkln0e6SfDa
ti8ht3V9Kenp6Xtkz2cPd7qN9bxtXlwsspwDUQqNCW5fX8DDkG7psZsYCpyMoLcJ
lsNAneplIFFCLSB9x0jwnnO8dKJy6ana4bCfe1Lc6/L4K7+sriOcJREaVuAPCXTL
3PLKReUhVPoDjEgH1k7qv8LDZECwHCsgmMqK9nfD+c84dOwQoj/4S9BajZQokzjZ
xLk27vtDDOetqcIR6LpOAIM4MoDhFAWPqOp4aQQE34mwd+CXcOXtZtND0zonqE1v
GRDWeLa8O1dLkOy4gDfQkOtcEo0jMZjfEQgwAbx+mRQ=
`protect END_PROTECTED
