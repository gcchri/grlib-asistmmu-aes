`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xwwDaSyDsY4vuoObMDgvdKkWaIOWADon9FrtcVEhcQa64JecNIvvfPRR0TkXJLmp
YtyfZZjMawCKefFEFyU7kUZz+Xs+SBdjtpmEU84PSFH/ZM0poKlxtLy/nnYNRgpr
Of1hF4ANApvcGwizXhSoZHfyVo5qwwaUQwB/VaSCCs2cdNM8kyPF1OLvJRtgPtNy
Dm2lZDd4xMsZB0FeRh9MNEfWWOO8kE1j4b3yJwar8ZCR0IR7GRZatfu8SEePuPjy
DChqeWSSizG9Az+vXNlvRAvr4uXceeB0RnP8L1jLy9JFQjeBuIAAZwA4Mj4hRMsT
PqLwDu2YgIY4hXyvoUvagSANUrue6YcCjuPMeSI+S7+6dDzFYraXJgLgI3GFztRT
4n9QKXmBPw4ukQi5PKZMWbEerh05PCZskkEf1LiExGqyLAJ486N4Cbq7dRAUMZOs
yAQRvEMlFc/pOl4Mhb0OYNRZbfzUs2zj5oSGVKEBvE/zDOLE3QRNZ0gdkAq9PUqQ
t0EKCw/eV7kttYozzv2wSiHmqQQ5IoivMbD29jUIextzOsYqnAmYB/XzaEjLQxhK
Ax651THaQrn3kuminXiAcBnspLhACnJVLQCE9bPgJNW5OeXplXDBYtQ1UMBu45n8
75mK61puWO6Uuude/3A7f45kOnBeYoZLEYpWm4/Jtk8=
`protect END_PROTECTED
