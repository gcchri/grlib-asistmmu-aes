`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uj3qORVV78yJBwkF9tpFniefOrQgAgOTx0Nr7I8zGKwIJMxxeeV+3fGwBGXuC1JK
T2d5VPoDuOMM9VgU7GsrUSvaQJijMFUKnrjik1DGIdh1JA2QKgTX5Oli94zl/07r
+yDbyMF1ThE0Woibo4JY/DEOXQ/xkLFUokIrLl/bW3eOZR/C5JOBPWYhulAe/brf
eCrnmGw/oaNL8OUpfAySx3/c5Wo8tlPfl/Ez4uyA8xCgdhyJWs9NJFtKLPrzC7C9
m0vF1BibOZCygYLQSPq0tg==
`protect END_PROTECTED
