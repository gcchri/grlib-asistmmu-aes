`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M0NighnTTZe5IYSbUc6KmfI64/8V2wLPGllDQvYWAxvwiOKLGR08T6FJYlCZuLPQ
PuEZkaCtSav81iE9ZPEzdliCXmMdTl1mwNtVNvkOP485rEPnUs7jCUsUdTGVW3kC
dnEu+MPWEX1us0NCDuvqYriZzmJVdcEzdR+lbor35rqJzgSCrJab/m7X3XZ+YmB/
bPo2jTJpRcczhTFnO07Fz4HJJD9orwDwT3L12Fsa6rPTwffOiOw8XnQt5JrFe9DG
hoy2NY3JR6uQarSO+QxIx2MakL1hWFdNUh1WcqMepKZSyQz2VarmjxkCdFfeaVka
CiwmdsdJDHkve2+nCr9onk4joWlknBE0gb5PMR2xZLOnVBXtoRtjdJ/13Ap2CMIZ
nfdCl9HOdjwyvdvEpb4ueO9UO/hvHMGo5CqLXYsMTwItBaKJoHoj6V70xvcpVAuC
HG3geWPmmQMf1lyAHMOb46y6BM6yEZFQLLjsY6c4CrKLZx5rGspw26K2DNYDb7uQ
/iyY6F7iiYFp3gIIBeHISb6Gg4Q/A8/UUx6vZ7pkRDyN/LB18zM0+YkendZALB8K
edyvoOXt7neAaSHqKSVTYArY1XBxG1IG8aLzOxbqp0aI2t/HKosEWJyO5Ws/NBRh
zbhUruW0Yto/B8buYq7qoSCOi7CWNZdpfubuyoOGLPOTxYBdD6PzIUEWcWtIOE41
o3v5tKr0w/8agDod/OeXSlaYC4ydLFvVILQjaudoYc5EjFhAkxHtSnPxFDT20aoh
ctVauJgOihRuk2nHpDH9FyFAIWxQ6+19z5yO2U228gcBNEcJKpkMhNqdH6nsabxV
pY4NISNYfZnaduiNHC/pWRoYPEH9/nWa3W3ZfbQLaH/E0nYE5m05y5+pb7VaYdBk
YIJbJpfnm90ajiPCmC8SVRNAWuULbf/US9ceFJFjmDaMDuZ+hEpzAyRaiDpDH+tp
1PheEUhg9UQp3vrYXGc+iHUMAkcLYIpNuZmcvDDiX2qw7OpbIBAAHqAnRcAD6BEl
q0Yikr1zGj5t4RbSjU2T1haeAP3+cbgAtFGEtjhtC2vLvpaDVEmIW9ZBvChImbvj
P7uy/wjsqZzRMpe6tu0WKJibjn4jgbBrkAveByKQi9TQS41VKBGBpbAek7rOImJI
gZY80F7LAqgskvEv4jo4Bn7x8eJpPB5uV+pEzOIH5pEHefIu+YTO2Yb+05q1alIN
TaUIYCOyzYh/AuXzI4Cx4h/mWWhw7r24N8/OceXDq27VKdL5tnoy8BP0YNgccIaH
u8fqzigBL5yL3pEZx5ASs5PqD+CZk5HdyAoNo7dwsQlHFOTGEUza0jshWqyItbj/
AQffQqfvTV8gFBLpfjfdI1HJPcWd70ixt8xl+uG/ZtyQ3PfdA3qDwyFWkx1qTq/S
q15aXhpl7pXxUJqTM416fKxS226wzNJQZE4vpEsaBQJLBz/cBlZyAukVn4Gz6PO2
/5us0DLsT1g8ScFHhh7A8vB4SdUWyioDoCfnqbhQTyTIwFSiDvVQCTZQoxOCTO6y
0kaIVVxav+1lcVjO29IPFevM0ZVegERe5IcD59dxWCo1w2ByNIODkiL54GeM2RGc
4ZN98Q/e1BdkafSVvbusZPckC8du4QGmPs+uEW5k+yV57CT43irF4gzBElQsHzeK
6Dm0yloks2c7AzefJEFh1e2ZUSDLLubK8uxSAp0ZzOIiPsuJak6Z6VVhBaCdNnba
MMeN5LzWGq3bQIagSadMLBIMmkO+Mp3qcyk2JZPT9z/s5PiXexFIieUXkwomjEC9
qXfgvLOyFxQNhxtpIPbkLHlQJDMIaTgMOirLuT4hGJRma8wkW0DvjeFMDGoDGzKg
dicOkbT3Ds+sB73Ok+oQWxrGMV7afcCQfvfLQNH1DRac3k+qCmY8WDEnsP/f61HT
lYWFj6bvry11xZp3yY4TqE6QApfuYXIFjU+5cbMzWWCIhU1RA8ChEWne0vE6JVS0
3gBgpsvRyA3fJ+ZvSPNOiGWTQi7DoUvhLB0bn5VxII0ILIeLUDoUOru7yNJ3C7J6
awGDqKiKO1tUHFtZlHL7jgEe6VVzKdJB541/89o77L3Yh2erAAtR8kQeJRwWhxok
OwsGUWSf9JDmG95AIWmslGp+yKve4A8lwEEF98x7KKmuaeyv+jLyCo5mLGDDHMeS
EtVCdEgaZ8HeE2XwsLRC7ri9wV536jHUEvFyk2CF+k/CS1rpA7PUEF53uH4XKSU4
zhQEZb1Gt/BMLkxhXYCNSlQ0vdvRprXUrjNzMigtPo0gWXcoJNjCqgGM2vru1aGs
Dt+rIKwGhiqgYm8Kqfj6CqeYympLkMdHnkRJ54wHUhiIOMVEDtpu8pqL5Q/S6J5f
DACoEbn/hZf/kjwkXvMsXl9pp6+5LTZk3lpm67GTD1FmiNRv+byvg8iE2Auj+gvl
jH4Q9IuiiO/PkpWo0qi+oqnvCfAjgL06QM5m2telbtDdmyP6Q9ircvz7p3G/qCl1
4aNXVJovjipET4jv7fSBzK/YF5Gl6c9cTTI/g5ZWUZxlldNi7MMnYpGNaCuevyaf
k37KEbhhyLSPaN+e+kRr/iz3+JWLg2Gv0XHpxoQ44EL1iLZtBNt4GnvGFniIqamy
uth5B6QR1wm3ZdKw+TP+ilHaJaMGf2J/ccQxDGnAIYcsbWVWHvWHcTIw2Ww4sgH3
OIpuuG7N6vOxxsihdkBrolA5GilE7plvqV5nG8EHJ8yCfDOzhVezCO8bECA1eARj
OY5UwipbPQ7wDXD94RpiJLx9qutptRpacQnklLIV/1dScPynweCJ+zThOUS4mKLl
wPk8qvFRfcUllBdT1uK6/FGlDUDxVa4LaEaO7Xkku8o9dTdAxR4nw3Pp4Py2tsha
Ny46IejTGvNp8/ZIXp3ILfwt0mqL+QyAI+0zBKY6gEJ5Vet79fNE6ghUSP+bMGja
tUn+iEWQuqpr90GwtZWu6sr0DJDqFEHG0Xj0DglqQp8RyWLmJPbbOtK0SmC8g/f8
A07sxAuNlKAM3ZnxT9VjL2ZzWzWrtOUqPaSnGAEf3i1JJeuB5p8+w/jvuUEwJmrl
k83A4FiCR2zsZi4RqSI0jlkA8KJbIlK5+G+eg3hICInfPVfZprio1gxx6huKGwGP
MED8eRcpioBHrZyDUwXMO7G0moR7quTxpP3JKk4HKIGO/ec2vBRalIKV1UhrvhOS
SqzMsrlVhUm7cOW52UeWqytlcPV0h0rvjyDwAzNPHOKNQnFrMmg5uGFBpBEdQfpk
oz+C/2eyRaIFjyPEKGv+Ok/VbvjHXoXfvsIr9zuAk2O/ok/FjrjyqQVFeLAObfDH
Il9Im2aEP7q3ARhWrp92jocTZ35psgIhRalIcvoQ10Ukn9G1k6plbosWUIhxnPSn
aHB8MZl0Upsa34jTdlX6ewuWUFoRBbpw8hHNcp4Wja7MTY9xOdNWxozY7ieuyVtj
+KnuJJqEbkply8r2c/pjU+2lBH/fLsHeAm16LPYUjUWaAWV1FLjEPEY9as4vFFv+
DSvBL2848X1UqAyRKRyTbqhLHUTtKAxwGQ4/eIBCL9IggnpxiQBJht2lqiH4c/Y7
uAV5y4kza3owJEw7AoFFDTEIqC6sT40SA5m3efpjFAovbtYDQO3THHO8YJEgGFhv
zvV23aE0ZIjFPkwPaZ8F/I3n9STr09MJPX+dCjErNkyU36pw+hsSgz9CCsioDFF3
yGNLq5SY7xO/tYH3am5+BrrJfKl5shI0mxMoFDCLg63pvZrz3pPOaTOzq5gaAIuS
VWlZ2wvWJtZrZbX0xpXuuB6O7niz6ixQ8lRmbGo3q6dxwxuSOqZCToAfhOItfZlg
Ql8Rk7NPBIiL5ADuJmOOdiSleRx6yVkmDydbE85UfqDpSUWGvNfzxuiNu0jZE5S7
9qv2FXddSSK7yNrB4EeEUoCl9Il4bp+P2391mC0o6G+BkoGr1BTPQ8mTuuYmupQi
sq+x2dr6YXZhB9Girb0IgXA9RFwqNS9N0O3n5PytQ+gtLsC10Z9vwGNpNUPBEFKe
pQMDrHkZb1djznZ7GvNUGc6KhFbrfzfIi5oNzNn0DfrKBIwROIIpXq0IMgbhEEAX
BdyvFpkwwV6QSt++fLwb0klZXVMIZrnkN78Mpc2PmjvfCqxJtXjhsXBjLaaIdpg0
KAoUGtHsUvzQt4AQ8HNM8un0sTqHuyUPSttmOhCsH7fHyEzSdwgx8L5Smw5UXL2z
zzEA895taqGf6qXPDBbrsIN9i2ijyL5+l08u/Ody2P0TojAfXMEU5utE2/9xbEEl
xzHHAcDLDf2qVwP2MAdtI+NXuLJJgMFK7PR5ABntm3OqXzZWiHKp3IV7Zi6ZMcec
XdVHpi638h1XWAGgTUKDU/xezF9jGCMy0/GITThHArRLRAfhgNVu/nl+lmXA04o2
0NqQ7J6uG0vHPZKPKD8x/5uVIAIO0mrzL7dfg4ahpDYrcQYTgFzT0EvR0LzdoRqe
432WZ4Xg8QzsJYIm2E7bb+q9Y5t+lGuOy5PyHMJddFGFXQXP1XB6VKIZAug0Zbu8
v0IZct1tOzg5e4SY56tXTvODCUW7G8GL2gnA5h5UH3Im7tqeTjEj538AySPYFlAb
8lOpr5PB030XjAXQbbGmVrA3C1kyjASMYZlIarQwHU8H1Uch/zL48NJKtZedluZQ
l7em2dxoABSwJ3pkt3M4D+NQOpFtXc+MlQMXPxdV9/6xp2ITBFK4xqywf2Uqr9cS
Xwu+9kaLs8GayBxVFibHveyS6pLj9BgVsBjLU5NT/2MDSoDm0hmQ0feNssdl3bCq
YfXGBXAXR49tnvbUhVK7haQuizESRjnq/wxyRJl+PNSrG0uqsqD9VH9H6WnsX3Rk
64ssibBlieSZPeLK0IXfNvuGhf/Cq+ezVLWWJVg3yhMGplChAoU/bXsO4LuOxtA9
nw7MA468End5Xx3Hchl33NF0hmwP4uxnq+k4pnjkXmwAdw7c9yGLHM9tDQr9W8+X
HDocYM9zMo0NlKbjmi91PCdf+az2hSI2hvmeCALQgXEoK8iP6Xm1ibzcbIjH8iMp
6bHkvgvdzlzXRckfH+p284ne2jncQQMJGgQfMJvpIac9H3WzYzB/76gdGtwydbpt
S2l3B4tL6Z9AQKwvaOCFxQ4l+3Swrwtm7YzbMbDYTPu+cKkOpTl8m7r5dIdtfVSu
Y46BwhNhIWNGJnolzWbHhc2lbXnDcCY9J1ExDENT9WlRKDX+3KFGEpH9G+JHlvEQ
ofqp4OHoq6DBj306VJWR0NvOpj5kuVFtf/i3+lqcoN4EBonwV47uTPzkPbhtX2S6
SnAkH11Bmxo8uLbybWiq6tubU2Wc0ioESueXYzxxtaRG7Z0XGvz5zol9jzYJur/M
S1JUcTjE4jlLJVz9zJ+W1Lz9WwssUSkYuGWDdHusquiz7Tx7hH8pWzCmjp0k0cvf
42LNObC20jrEi9Aw0kOtVtlNSkKC93VCndD3MhUVkztLh7C76TsnOAG/qqLYwIlX
zuE5E5Tla54p4QMQKDQZG516+F965oc2IZ8Ms0w3ORcbk+NNYFo/AXpgq5D7yVBV
yzZuUIf8l2nFLR3r8fItj4XytkKUuWuFkv768H+5+y10TqofURwoBplWgeLLOnKT
27dinEYqcm4hkqR5n82TQO5JUS6qDEuWxAh03Xq2qsjBYEQ6sTBUajq9T9eEmVYi
jsNLBWwhNqzrUAcsoPDXfMbMv0RSZpIWmyR0Yzqamx6yPAqyX29WOuWQVsoJn5wS
`protect END_PROTECTED
