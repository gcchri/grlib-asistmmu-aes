`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QOYDv6ev7vSay7dlfPcck4jd6qFq9+38qy/PQPGrbjqsUefFJNhahcBPnyB6ppic
RVxKEH25sE1wRjQ3k8itR3E6vAtsztRWB/m/Zu3s/3qxdsK9VpCZK5wolfnaiBAj
N5sUyCdbV5zgqie+Y/oBoXWm9cPgHPoasBVNxioFXTqsDQp1ojA/EICdM3GVWuTr
oPn38VpLbMZhqNLtaOfN708VUuaYazs8x+5TQEgnYLHNTsXGhO4Gys72vO/mveqV
ClPRQK0fcDCiWly1W1EKFQudjOtstrSr67Q/9q/I7TEfpzVzoXvgYqJhPNb70B/6
aVRUOABb11XPagS47FB1iQ==
`protect END_PROTECTED
