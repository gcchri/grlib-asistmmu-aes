`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8jtiCPtLc2UHbNoYOZ9v1pXKJCsNfEwf9cYoJ2DJR2ht3kw1A2pLLK+E5dk2s9YK
sJ9gpnD9pyn07CqMP2yEhSV21CKCYpmCkVa718InRdouOZ/cQPvEuyD7aMFh8g42
3cESp/PYa8KvkPmC0D/1S8PxeT8yZFDBiYFv+amTqU7x69d7lF821iSD2wa0QNrL
S4uo8D2IH/5Nj5Re+wxXg2QaMXgxpKl6IdBhbbckUyt6q03DtOzGOhZgykwjXUbb
5c1U/Bbu4rMj4LdMfh22Y3dNqbGwCbmF2Q67CmiiN526wa6FjyzMKdJVt4RwoM/j
gL69ShvhOc9RbmJsqltJf1npTPvf1KjE4hO36f0viS1qt5VfGDGjvo+BoQXUHXxs
UwlFhfnbKqQD/ZtGVS/XJknnpECVlVYNLbyBZgiDDJT4vNmsG/ZNf3Fyaf36ZIbU
uEr/Bm9VUFk1XoBfe02Kk4vWMx2ZJK2iq+FGAgbZDXnT/Vp5Zvd/H0dTzGmgiYnx
VgTb49/4QLcMyyDX8x3WbnWlyFbH9GGnTmrNp8GhK/Bwjz2JU2NT0eWPyoRUyKxr
OoqTeVNBKsoMmaGeJRJcRDJnVXFhltBoInx4xeEG8wTPL2ZEQIstBzSpC/Y/KWmS
Lb60lsP8JdaTjPqAdaRHhE8ydfEbyZKQxEyYbw3uPTSRhZxlRWQBe6P02BH7znS8
NNuLdX/UgBKJ/5SSAJr/dA0JMFdPPVti2JUS5LdNf8RpC29JPEKdDW5P0cH6bgVs
VN13r2KqgLqpxHi2/vnPhgc7pVcPRm+yvJIyluTNvRcQWMtsIPugYlPbhJogaiBa
fAvYURYmFUf1RDebhYsBpOk+UJLKhRMYDBz18OFHM9yVHu3fq/xSasUCLYiuY2y7
kLR4oEqZKdGLjQBTwcvPnuUncOIuvl2Oy81C7h5zOlLBaWUfzkzOOUjmSn9SAUPV
u+LFlvjwM9H0GO8df+I4RAIWppnW4QsuIclLa8wQdW1Ul9heJ2u59vx9irakv94+
ESwy2vMy05MvZjJhLKzjk0cnNKSgV6WaYwhccQyBnlPnTUHz/vd85Bi4FncBTnpO
NkfVrDQ8J9eS8rwlOL7Ceb0Zqn6TCSy2PHybhn32iaPF3eFIKqt7EwrNeImA7Jvy
PmQvISPCJbqyKoA6ULQJ14pTp3OegwOEpdE7dezzjFSq7bG/1l0rsgiA56B13AgX
/p8GVwnxHWtSf2EuMa27pCO4Yt4QvWxJQ5Vj5ODOfi8vICnUSovMereE/5DzTT3Q
7K0hheRnRSdtVZkez6VwzA9bQybRlJWyrE0bCZMiP1sJaSu34AQbP1UtyjGr/RLH
wlTPqdT2aCxki2uuw8s8b2LxoTgF4f1UOarKleom5UIm7sPAQUUPFLM2Kdr8DCFC
RKOZRr2TdtkYSqVvS3bZCW5NnELnUox059p56VuIHh+m81tKv2hCOpd7TN4XHIQW
PSlzCnGgHhdU2SfADFL+nbMHDu4HT9E4/1d1Ds+IS/dGD2ubbWq0v3lxmPJ/ke86
FMxPu/2anXhe0wKXurBCcmCT5WFQC+ZIo2OJ2Wh889l133EyWSZQKvFuOn12ebWq
G1xc+4QuJtXo3tpUYJXcjbv0ZFnpFyfyveUkxTbDIObJVIS6Yjdblx/O3YxPTNum
nSjIXFt4yyiSKa9OqT1wK0Aqfw376xQ9DexYWNSxg6o3ZPaGyXjEhqyQK0MQuys+
nl+BKoO2d4hNGnAh9ODyEQwzvY3jmbSH6dP9FLEIITqb5KRgSpa4IiwrmeSkmdTc
jAaRZEd91vt46oa+gEVlmxv3BTv8K4/l7ZCkHf2fnpTN3Ci/21nwhW8anMs5Nun5
U+B04JTXN/okUH+iHDXQpO5PYZw+foGlFikzMuDBxEcdnjw7Xx2jvyOYdDmm7qMY
Q969kEMVe5+pYfeeZvOh7ioAVqfwT5qY4f42A0isYDQXsw/7FpregM8TDy5599oO
+M7rzNGjDRVGrjbwu/L5HuFRFDJPchRvb8X941xnxMSsYl1soJfD+rWeV5M2c9+a
iehaLybMVSaR8hNW01783KlZQ6mEle9u7IKKFeaCSErzAe/diKLtbaB6xIYS7iuk
nSbWSaUyXGdQ0+uglnxCdC1DZ4rScG6opKPIh+G7OsKb3poWN3E+iHVodD25vA9y
m6lcrr4dipNJfkvJ+nJxq2FsAbIBxjo635kC+wKNCs3x4Q64oBqz20/mJyCHlUhn
yFgSe4QZXWEOxcuz6+ObAoyqC+rhcpjiSgBThXeeqKKUaoVjEXtXqyxFJuYtAyvh
WJv8zf3Vy8kvZHeG/+LETIeK96H9pmmC8esk3QP/FLfASGXMQ0/yKbJCujlZ75T0
DwCMbNadfGkCdq2d+IxN8qaNNElWRH5QEkOwdotvK5DtGZ2FqkmF4g848P6ja46j
GCtWXfTJxg+S6TMZ303iBjgdSqeBmpRJtA7rNqQlY3DI4u4dCZ57/GVPqymK4xuM
QENByXEFF69t/vP+DReTv3BgfD9cEu2uDf02tw13w1RrENzV5+7A+LktbnX1KWhY
CJvcT5iwDOSmLh+Ns/0wCC27VSa4HfJ/Mt1OIGP9LrcB/upclZ2ZXvDJ/w/KyISc
iSV0QcgIDGl5uIpSV+ZEu+E0stceFv7s8APrc39HyM5ORWJfxL2XRNfukqRgsDr3
Rt0SgkHLNUmKIB7QG7c/eEks1qaTC7wtiDmZW+441DvCXGG+xDqVF6vw0tstbh9w
RTN1+ohvm95Zerpo6PuVfFcR+RPgo4kunabt3ov0uTLwTrJb1pisC//SItdN/Alb
7LlVWAeo9Q2+yRipmK5QZ98DHGr/Xi7EpcrvhC6R1X1joqqFDJmBuOFl3CWDvpaB
XoE7qL+e55Xh6S2VTmPQKXWR7QacIW57wPT1BW22l1fEcCnrReZZ/uZBSU61NEfX
`protect END_PROTECTED
