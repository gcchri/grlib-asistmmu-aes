`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e5z1zYXiiweetCZE+Yq89d8+txP4+YOnHCoFP1Hh44vtAWUq0pSEnbI58sX/a7tQ
UvZQXvwS5buzZW3ixjx59ztpXbA6KNNZ4WFkpc9n/1Sm3/nHuMdsdN7G2xGS1jw6
BSiWIEAdZcetfPv39ZIa9YzdAwaQzF5XQ+3XIQnTC2VvYMEoZmR22Nz9Wj/sQxvI
XO10HRr7mnNebNi/IXixNVyH1yDwW5i1x9AQWFfTaUYJuvmEZTFLGDF3Z8wem3Zr
NgNsf+UQYhfFHp+dAgQ5JiMD4p+CH8uliyITR18LtuI=
`protect END_PROTECTED
