`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GFMISUUmzwJusnPdGr5WnXegJk/vePj9VSYxuSwCOCRo1UAFxQlcgkIheLQhwGR/
adDVO5zA3CLb+uhgBwC6My3aKVUTrfUY1v9AExkgEdSxKjp1lpsz2jSQpi2qM3uq
j+8kw9ybwE33jCnYHC1Ql+izVsMkaXX3IyAXlvPcQ275wZtH3a8doGKZlJSQ+2bT
7T6vKaMAr+ogdk7VFh2ALoljCjQlpbHVgSkFOyhcwOgCMu6TRR0dWH9v1bqW7vw3
IX8ZANuqsEpUMwzfRRnf2QMNJGJmUAIvTOa3oBtpKx+gutG40+3TUM014TJFBQUt
PIMYZLm1aVOc4YY/68awajWRG7q6/2wXxQfgzjaEgceg3WgpKueafAgApKL/i9nY
shCO16Kt/1Uuv5pU4Rf2L+XT0M5BUOLDifJrLzKmslyVD0ZhJ3IJaLuUwcPoFvdS
gku3XCYlc/bFwbtdEnzXq92B3GJlYRpMdCvC5PzqtYT2mqycX77LVE2CyjeqvEPu
t3soK1cxWA52GqDRrgWI9S/0cL3VS+1QVuIajTEupAahZIISMb6vxKe+Iw24KQzZ
GojpFtflCg2AQaIH5PyyTIcp5U8gCxwLuzOQ8smfWSg=
`protect END_PROTECTED
