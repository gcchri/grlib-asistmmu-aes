`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3rp6ErQiERdTClOis8uBsUFmbxUKUn6PKiNATWYiqdkrBxYtWTzaCzR8AL+/o315
+j/Qq+Z7XF2FLTPqM81xccOZkjj4wz+CVa11aAE3gHR7C5iWPQcqL0gnbIs0gfQ/
TUvceE8uMiYYL+Vg2cZ988dEJWBQFzO/d7VWFN8e33cBJ7A5m4+/a3L2zWQbVHqp
TkU1kkYP2k7Dwbx/vPnXdvQkrRR1Z+YFKPBZxQpxklo4DDPRKITHbOA2goXnjq0x
QBjjCaJ3i1ngVhwDlPI/4fjeGOdHB0Rp2SsX6nq6XyuL4N5EiQ1YAq06T4V1AQoe
MdFGrLpSgvW8bYxySE87Ho52JgLVHHEjDkq3s9DMY+PLSF39MPPE3mTRSTfhR7he
Y9IW3seER8H9e29cAJ3fqssSyUfTSGs8kICT5iIcVHTEt4HkV8RRvDHBQ0DDfCAs
8QJ7wlhIWrfDJtZ4Pv3fSQ5Wh9UU2P6PXUxZNwW5LNoociLEszbNTGN8FAZfEssL
6DyrGyLEINIaCKkqr3CMteczA4YzGIk0l4GsgAnoZVDx32bj3lKy7SwZeDzjMnII
fQ+lf+D2f+rx+WfFShPSbaScl4/zMJzJ4JqPfYetc9GX4CsTJ4U1TXV0+a54A+LN
wIBU6UXkQ/jQ1i7fHizJqA==
`protect END_PROTECTED
