`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6pC3D9ChK9mlctkCW8kIGJVlSdwNOQMGJMXC2B/0JgIaLaA7s7BnfObaxlgfQkeA
ICqA6136LdU3ZLoSb9KJ7jH5IMloezCypPcElQcg8mDsKCRdWrjXsdk/3XTMNGoM
6s+kxK8Ej0vcghsFYs9cCAdakVh+4tXjqR2pPfSaXs/b2HergeQnDm/vJcWU/YmJ
HV539OgI43BQ3HbRRDCb5y7of8+oEtI60HwdTY6N/l/8OtpX9cQNk4FZ4vLvVWI5
SlIrS+NbFS26xQm1nuq3oV0VxZSy3pcWWj+57oqVuACrz8LpH/Vin+XoU3vmMKek
l2UWjOzWn4ZGM2ZlTX8f1xnxhgKKXImRV/d+2BkpdKL7Dl6c0mg51zKBKyENnrvh
6D0dtnelmJMKkFLGAqa4NGrgDt0eqxv1JieKrHC0O1ZVDEML/3KBopVwzib4DUok
mSOkqP63yAxiB2ag7lyT7ROcqQy93/jXubHfA8+Iqouh6M+irOYUwZiuFcpiU0rN
9RKykGBez68+e6u0AUSBsowIh62ZBVrQlAxeuGpAVmbOItL+sjMZk956PDfj7Lo+
asXjrw+Mvxc+Y8nxUmvTsJplufcjcD/dPUY7UHILbcZLR0dIhsmQw/SoqHRgaOCl
VZ7iObqXGDJgWJ2EhnlkjLZ5q2jsx1b2LXqrcfhKcSReL01xcscVZ4jeGT1wLaDq
W1RUA6++eFfVIJVJCXEId8YZRVfZ7smujPSbI6wSkDG64Qu57LcyFjKvv1Q8MAe5
yyXtBrre8rs158V+f7YBV1GQOOhqH94KJ4CHvOEr9FziWCGk3HHuumpTBIeXAMKq
cS+/K0n36SmJTdTZ3QV6OK1U08WZUZ+nu6gUxmup8cW3Vb/GD/AcG4fjtxsXJ+vJ
CdhbB6+bM7yQb5LTMlbnyFWREDB15DJVb6YTX8tvN2zgGgBm/cjLX3GXerVRMN9A
MJLkVCSvcIKpYDxH9rid0O2Cui4fT4xkJ8shenxdM3uYC4IA8G9/YcnWCPegyxU8
U7z1+0Hi4jSUkzikVXeL+/GXbONYe9iywuuZy7usBspy9hrv6hvNJ7az5Ddrj/UE
HShgW1fRl1XEnKTBBhwz5S8dHwv+TJ6KI/z2aGzaD3aINDDElOlRzRh3yPu9oI/h
qS04RpMMSyI6NaBEpztbACkGyHAHoWqN23tkt7ND6hR6Zt0D5DK9ptcNYyya134h
H42E5qKYzvCRvITkafUr60Xg7NrADeS2gLvIO6QchzSaqjRiqBsQtiGEb5APeY69
yMuFNfchIUbG22UYbSwU5A==
`protect END_PROTECTED
