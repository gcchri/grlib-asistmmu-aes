`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vrZoRit+CrTv8B/1kdzg/d3z70BROb0ek1Su8sZHc5BHPtUHXiv6u0iEkre21co3
VxctV1mVVNhd9nd2323l92agRtOU2f/F7cAExPXcj1SwWdF6Bb3Sn9RhYq36Gc+3
5fVeYpBUeF9UCFT4UXc0QFsMEvASVQjYYauHFBfoQadWStr/UgzG4x38dl8aqTMt
wxcJoFHIe239nG/2AC0F3OjrAt5S6fk7hfGeKZ/JBvD271SConsrIIrarCUARmXq
E7VotTLp8zkK3Ua/yjFoPrl0yB5VCAT1aq7XsTXXX2GdDy/wzS/eTadP/St0LdpU
z/nEQeB1l4K1mZ1+bWszc2QIaZsZ3O6jeAosyLxS+DTajFW2E+DvUlgNSenKTyDy
`protect END_PROTECTED
