`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ScoFRFnTP3FzeW2D1nosL2A/g5MwgW3CPo8YUkfQ5JIq14miiC09rm0dz1y00Ia
owme0KwKL9dSb7TkMHyXdqQ0DNAQvXlv0MmZhK0H3leSd7l4QpZeAisAsijRA/tv
puNqRBymUqMUMR9phy1bC0CBhfznjWIZV0YzcsjpqLa9//A3kwL/Zgmo0gauO/ja
I3JGpIiHX3yOI3Vbz0hGcJakqp2y9KTs36tIx/JAL1FvEyWQCUmDdSPflgm/PibY
pOtYW7G7CY4XHf35V0APyW2qY64PEMbYR3/JhlJ4EyGGzGZFgz5zodMqbp4C8c7K
qkeYbnAd/6+csFV1FaGSbKopiTFsKz7A4ZEbvvUSIAXT83BhKhGvCiGsQIw+/Zzt
Gz8qDWlgccVDPsZyHbt8SSoKGNeJk2nttPlxSYDsW+SLl4iw8QoJSTatdgvfAxAj
y+f8GDIOlFCm+P5xWTzMm9N0jq988pxDI7hodtDHi2NMrAyqmquwX3qZDkk2Y5HL
y7dtlBeH5l3uJ9w925hYma1250GCy+/kV5dBX1V+Ey61RCOH73yKBMQLjpbSOw/c
CrKe7tdBhgEJ1YgxtSvFkaOrejBFKkzI2+c/hYkeXxwPEQlOTz5iq3JL2MUBmPW1
DlEFaPBoOaeUpb9vsoAxkUOQ9L110tnzsCE/4RO3+zYbsrkm6KgJvI3BbuljAMSt
Rjyq0LMF5+25p7CU4g10JTHf8bARiA+QCFq2yBPRmDTkNXWbspQrHjifkgl9neFw
91gUQDlJjZM1n1KBi9+2Rx/kYAlR+Wo1tgznpwFrmya+tPNlivr/lswUWGmN7ld6
9et/048v/6a7lvB8sdBRmlzRCtiqwg1n+BZlBCFd5UUPRCNsHbqRR8JW+nkpjiA6
WkjaUcuFbbg6PoKtU6LK1A==
`protect END_PROTECTED
