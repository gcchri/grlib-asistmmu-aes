`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vg0rqk1djfcIwYoY1V5NpVFqyZKoBgC8le8vv8XuOR4ww8kDEv2S1Ds/igP/4KGL
Q+vrsKNGvlAQXQ6p4Ld3EOmi9hcyxsheKTGrdla5BpgCOC2f1o2v4Noahqm3CoCP
sLc63cD4DdY22EpleYg9kiMx0mBXui+/awgMClYldGlUp6KOxYepKSeTyPxXtvIr
0yXxOr2R3uyZo5rVe32U6MO8y1HDnRa1p8XlfvInjvK4UV2GT4FXZFUqNe8pGGmk
QT7qqqvSalbL+Oqoi/1F5bHLPy34XBNYlx/HLrU2gQITiXxiRVkK8MhgeN1XflEl
BpO2+TF/1pkksZuqhlOcU9jggNXjkAH1u+2hF93hWgBDYM0LsiEFk/Ehj90wbp8V
kYdLhlD/pLHmCn7ihMgNCA==
`protect END_PROTECTED
