`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZonF5El+B2h0+Sn/zPbVCRIuaFNAZSx+XwqrbzNDWjoKoW7FcgqDxrArCRHHKJM+
lZ2nSTpP7AdVYlZ2vonF8vOKNwun9ZpRizZKKy/RNr2FE+SjFbKQjDdOTxbH8K7J
iTCKdy1dS2IbWXzKfTTRO7/6Ee5MLLNUDN02707B6Xt3V9PtGxi84ixitpWuyRQD
pfjukGCXZoDO+ltHf8HrKNi7y20CmaXaWcNpUKhuFMIB/jRMzCj0hx9iNrZiOmi7
Z7SfzqFOAs5RXnz/On4o1DPVHOgjYm4+owQmzXAB6Zqg+xl3Stt5WS74oZvZ+lU7
RXTYxZpj9pjLdQZFZMlU1fpopR5+Ys31hJMAdTyKOlQkb6W9ybzLKrFvxQuXWsIA
KUxMATF1Ry+YKPYIGV6roJq26xSH0Wi3GqijuFLcibmIS2PPZ+p8clM/aaEkowUy
vgrUJRTWshZP8JQfg3yn7tS7Vu64d4k71vHRyvnJXsNl5M5HYwEAPptL+pq4boGT
e0wlHR3KdNn0s1XcEIm2B7QnarMCgF2857307ThcQajK07vJ8icDC2Zy7hpyZwYo
JSapTmimERVZsH+AFOMjv5AQVrr7o1FctQ1cK0yxaxsljgtm8BsVFIdw8gYZ1SfX
j0R7ID9GCWrvtH3INf2ULrtXOgqmtnqzAjQ80+ua5clbsmjVpG1S0SAvJ4/vUm/l
CikDwHxIvKTnf/mpELyN7Z8QbLQan+jziboigPOD3d0wdjaPfeLH484ALpaXh/VP
qp+FcrjnDdGiBLyLzlRYJIeDHFd69POW6RvQFjqgyZiFgAEA9sdHPvn45yH0qyIX
6tEXFMnIKZ9wVbwErUkoc8FIYQdnaUPaEDPeIKnYz41iLmG2j1/0AiClASb05Gec
N2chgwuRqRuReAcEZZTIGB4RAzBGIiPtjDSML+7suYsDUzfKyvzo4hh6m1ffrChu
rthBtHb6EsLKqcms1JmkUL2SJWeRmAIXFzHg4ijadqT+euDliQF1JWWR331F8o+R
FBcKZGvapT2GiAxxx8miuOSH8ZL8BEEKlgD0IzzHt78m0g8c0bLHQXTBV1/MGKbG
uYFERbEKleUttJzwY/LKrvRr982X5176AMdg72jlw8WC2xYIpSiHM1qG/f79Ho18
pzwz6Ra9HIW8cDFNzNsq8F3N4eePdWeK5mq0yY95dRbEbeMdRBKM2o8YrkTvLrCa
m8g17m8HoNwVLxAJM9ZuhlY1aiBbgbJDnnys1N8RtAm3dqcNZ/XBFRcZNPH8Bo9N
Lm+hIUNF0HaqbeagiQQY3wU809OzgDP6fz+BhtTsFgCK6BK7f3AV88K49kVzslmT
+WDklWmGaTBcDkHYw2sqjqD0WxjGvo3td09wz5X2G0WMy5rM+S7JPf7up3CdQ8vY
o+kljBP55mIanoghIjcbtBcr72CWZ2TOz45kvUUNpirCFbxNYXesg4EsBTAi0Byn
gS0zyRmOe+KKg0e3A6RfIRP/b6pKbfWOzdiFYafUqTTwm2QYLVu5CZXw4WN5mEZQ
BE5WpyUX5eFYFHD+uIEcrs29Io/NZQD63aW8lNeUuiZgUU2xrYGBxjyj2yPzVSL1
AoZF1/jyIAuj1i42JxXZ2kbwP2XnGLVsYGjvcKY7ABLssxRn3pjP6MuVoZwV5ii2
fmdhgHTAT9uzE/jec5BHVfDZqQfONnm9/UWXKf1TFkpSRXJF5KbWYlhtNuGFkiB1
DFr+60hXOgcxC0mokrGQC6daWLsxTwCcDNc4k9lXUGPInMuXhFQVJQWe1PM24j3m
N4GGMpBh0F22NB6g+JyCOBjkKWUmMFbhbKUMOfa6Q0/CAzS9PEkbE6uS9ZqXPBEA
steJ+LtR7+FR3USO1FN2+nxVLKQHZ5VGfqK2QlhB7g2CPKKlZmEA4C5WB6TBuwQH
cyiEJTLuSR8vE25r75v91+z66z5HMVBos7btItysB3DKl/YQmBkqgQHow9Cl8KJQ
lst28O9Ptonael+upr2GSj6mubvSq+/KNSwxcGaSiUUPt4NKKnqidn1063d8LygB
cSUgHvJxYEVCjq0Jl6GbPm2SV5fochdALgqcO4C80HOpNBCDSzEEFqGjkAUVG62q
KnzuPg0gp/9H4J5S4FEACbZblDe8BTUTqz+9Kzkpvhh0MKpbTqbqF8g0Nw4f8XkN
oQI3zGH0Yqh13vKOU3FSZvZvUxhptsmJjFEEE01wz6zlD/dnhuCULyqOvVmHLLQO
eVuH8MyGvaC3KM2NuVJm0riKA6ZYGZLMqX3UOOWhwpbD36ZRq9EzPdlx91cmGgzb
CfalSq7L1Ix0DNGo2JOd2Td0Qah2DQFMs7KrzoO3g/pWA79ONtuHErEeT8hwKTrD
+OstRmSwRMnCWKpkoa4krfGENUX22GciOMZk8G/3T3S2Je6R0zMOASqMK+iAs4OK
4ciaDTGSeaDj++eJfG3nEslkqNNcxuGPrSpNKU7Zl/Kes2mY8iXxWjBqvUpakLem
ZPy1S9vagAkNklndmFeIKJqM3jwsU6qxDfSYRVO2xOGQ2tUmm99hdPxLlt6TJFya
WRdJRykmWS6V8+rfUVygdZaOy3+U3Al8kFTdmhmWHcQCC+UtLGigpY+2sJzbdEGY
EgYDAbU1gHpjZoXD6QqGRjhM+LWQYio278yqlvqc4hUdaNl6m6GRNJ3TXM7mJjCK
S8r/tgs4/6gsjoJpf3SzaYfK96QwsMKOZHld4z0VjPEGBtIuvNu8bhd8yB84y+K6
jCGJCwCUynCXFKzRxo6HSjzweyTM9XJVtkW/p9Zp1xMacjQ6M8NLV3yM7USJqqJe
sb0IOspx9A17Onz2sqGtH6zpzFKljekCEliZa28pRU/0+KxnSWWaGMbIhMa+ZDuh
lRbICpvbJx2mC5wqsPu5BR8GpGi1S6COBA1vDgZDqiTLPBg3+FIIct9PxrWxTjC4
2GnJBxgZQU6oetYRTaFcQmteeT5971PtXWI/ydRx8lqYWAYnhJ8wdCO5gvOOtXUL
FFUw9VnajQ6jpZE+IcNp7l0cDgHju6c2Lgx3bgTgU7zv0DHce+HpGKuy0e2mLLPc
BVCuw/sawyxITPFWGHG2Iay7UdBTO3CkU7eoYNbmygvRuQbugtsUHU//T/kQ1GBD
EEvvrcZuRgHNuHGFHppxFkKwmDu8yWaw9PXVrnDR+v6rXI1/PxklX/FQEzH9kxoG
TFjNdjPgxH28sP0SKd+BDnnt0+N/1FCKw4ZSiMWKTt8wANbPMW/sOESz1MR5/+0q
E+86y3fvBtWy9a95MLDyosJ941Dp1AmlVkHRyIR41FgeRVcDDk+9OOSqBf2Ul/OX
XRHEfwEWNf1cSUCZUiRYjQYjPNuJt63BEDon8VYnwFl7hASvCO7KgeT9b6bGrhLH
rbE+tB51/UKb3BBmsNrUGuQvSPhF7O0KLSwKvQgeR8uaUVkkhBqOQ53CUvAlzji8
aGXeYSi7gAjo8Esve4tZIucO3AuLp2IDbbYX0UyiroOnmy92jysK0JwPDW8hjRyz
C2FrQ4UBNFTeoapeCaP9ucQYNgalWQoX9jTmW+Vdgl04GjC64owcHZILUpsYSYur
t6gQz8p44Sprzh1w6BWkYmrxCoeCZ4SuLP4v6mj2tFbW0cJQPULzHloYNcYGOFSd
B+uSYWYL/CWmYP4Vtg1FWYejEPSZNE5yb1x9hTD08L1PHbcIR0961MevQITcWseg
u+KVOCna6SOpiT7OVeJsXCZ3FIlatHDEuPibNvPcOGalLWuGRumWMCPngiyOVvGC
MUNDisUm8zCI1S/asNgXMawzTJn3UMgIAGPJv/ANezQE/htBQ70E+4AUYDSqOdyw
OLpn8gRWHo8xU9nX4wCywQmoN7ZqNIVo9bjfD5Tu6+U=
`protect END_PROTECTED
