`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fnDluNbdgWH8y1WSelJZy3SNkCMkYQvF9fbf1rZLPnGsI93G3E/YmHaYtq/8f51K
iw5rapdN2g6WmZl5fW/0yYWfqsDavFu7Q8pOANnxxzQdF2LIQU8maYbMiDGfdPsT
mrS9+mQ9WmF7AqB9kBY2MXxp2RQvLwtOVrQec3A2XndCvj8/Nz4CSXbKz6HuvSHD
Mo6MRL7OZieEzmanm6jknXsE7BkAqyXzYKh+5g2EmqziX0lR9bdGAvTPh+xTqdW6
XHv2KZ93H5sX7DogS2yWceJ4KH7YkJpXgV2XW9QbmdSy9SupQzJHcp6uuoUXDWYg
Hj60XrIEt1Tr1YT2E35H530NR8z7SpdxUYlgMAGCPHd8ywvPlTDdjETesYnj9uQw
/Md498x6KDXZi2yVtsmRpacLtlp6CF9XVal9pmcRY0SVRV9UbHLP6WZecPC7WN4o
JNFyqNas5f22Prv4JH3xMXHfSxd7Z9ldFIJMbJ0s/iy0gYICAhu3KKboiAOJokWM
jUbzAufkJ2OLYYvjTd2bQ77sci14Z4BLHnlpof+mMVg=
`protect END_PROTECTED
