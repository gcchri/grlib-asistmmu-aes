`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zzyj/Jb08ELJoceGDgki1Nz/OofIV3AnPR27F/e1u6kLqBc/uMk/8TnaE7Iic8pr
2ScrzEDEmfMYkTpVzYyf7fogG8TQ8TnhVDp+BIZA8QEjnA3vt9ZJq9jVWrT8fdH2
O6+vgemdy5kywNqNqeLAh1VmboaJbv/5aWfQdc5Ong3JhXN98C8eEYpzk3FJ/beK
aK2LovAMCObCE/K7onDJmtvFqz67OC7RntfNVD5eJizp4ymyTE8b/vSF4QhgdjcL
0O2T+OLVAU3phT6F0EmNep6g+n+kX1t97+0yIsw7LvYdzOZq5462oHxlne9kDh3f
5CQFhcqWXM0keDp1NtNLEEpIu6U6E/vP6zpW2HIor8B9fFqEJJozJvBvWjb7yj4p
OuPsc8lgudisC0ax7I5GFosdXOTwdD1bBskneEF15WZ8MQYknKEm9l2/tFd1op64
5lo+yR9Td5VACD9vgE5OUvVAkGRu/GPFWWg9aMH4ihC7b4X1ur+eT5/RuwvQ+Axh
BJnUe3HXi0g9FLuh3s7EY/H6eyk3ia1b8Iw76/8PBn9LD490Gv+zlBotq9ZCTs3d
b5wiOy7Tz23nx1FaJa58RkVWXVgzVuCQy0d4FIfpHG427EFNddvxUJBgPRC24w9Q
hTgxgwTXUu0rgjy+DnPh+e23t4wbJWsJfBk5PxfowT+tKEIPHguUjryTawRYP60f
64hYahzMmWwS1NPPde2IUOrqW+M7x5dvAZvY8wBlvqMPRpW6PA7YnKIIy8qYoWF0
QnWX5yj8aWJs7GrQD84B32HB5WTHpg8siU6y6En2beHeKhEmurDf+BkRef3aX/k5
s2c5bUfLIMaUsFkRGTCApPJnyhx7rzlf/rZ5vIjupsdMkHnakW9yZWCZsKbBUPxB
nDAPozrfTv7V8pc5RFgpwyAhIx4iRHwLGgbsxdl8qACUfF+CrjnIgoLoK1pOIW/g
F8g3dsVHr2Ce1UF2Cib9j3gL/4eqw8cpmH8yJbuoy452aVEVzmoL3FS+HwWG0mqq
dATATKej96XKQ/WAHdYZM1nzn3o/91ANL54Xl3zlYZX/djQaszi1NM+FO6oYofpP
CsF/m39PrmOHacU2Vyf3nCcvY2Prj7rds4XUVBMB4aItvFw10txbql0I2hD2t5NH
h/qnbsNZVCM5rzjh38kx1JfPmP/CQyfIhLa3EkW7vtP4dmDIIqIyjKaiSxdjR66x
9f/Mk7jciCj0QSJz34+cuQ35kztTbSjxSvqgjkUc04SpnN5q0Rr1wHFt98yMjMZp
CJxMd0Wni76b8Q3RhmE/EI6tckHZRWI1OoEvKNvg3vbfGq9dTUfW2SjMhFZIAuKQ
eRX1KCc9trBGow8mgIUWdtOxAmhaNPRpGA5QL/w2czUmgKEShepLq01w7Qw4S3nV
ehVj6v0GnmbNfZBrrfIKkhwEOiRh5H9yQg9zBaifZBZ719POac3Chw9PYNkLSdIA
KHfTBp/SDO0Q8giDj/3ZEU742oJYxrj3oL6Dlpu7ceXQpDaVgdezBstmCMSogJ3V
2HTYnq0iLHN/hULjWD/IK11CrCXBrAINIXWQPowFlKC8+G+++ER4zjoC/5tf34Z5
91L/zjZxrWxvmKnssSdb1idH3ChlGiE1Z1CZ+tLULzhLnT5sPaLpfgLqfsX06oWk
HpG1yjA6eKMxKGm83dgNflQ/9RAFmfQLSp8i6lZgIN8twNewO9bKvsXiSAD0zZpK
FAafAbmx+Tk2zwShMN7FG4ITXP009t32novRtV1lJmNAx+r2x0/Bclfpnf/cUfOB
AfqcigHs2DirFCQzGRZmeMAbJ1fFwcagwqV6fwuZThXD0QzIWRHJrJvBGHzGweKW
I6dNyT+5XcMWRL9fPSwnTFH5wKF5KRSjP62JvKyJ7K7KtHutvRm4+iqJvAm7uVvr
KAXZ4o/ONRpB8ul1wWLBUVYsOPiz1Q28oKixtwJfN6owVn/5+uxYWnP1meyjrOFx
5BhP1Tiup/VKd/G6VljU703KkbKrhMD2iMp9cGc3c2nqPf9nLKHpa7qsAVVqGMP0
XstuDWPulwp9+pw5G+yApoBSrnsLETyJONnL8zwu+okUQ3ZT+CW1qePD4XfCtHNP
CNBF6yv1gBBLnQm3tn7uIC3bFUJYLl7Ehs6TUtG9s1geHzbuAm48N6p3ZbbnRFxE
1TKy/tY32QC82IWqizdXHZhWTwjyB3CXZPr0QNPB5MZXXsgMnwVuTPCRlm7I8bD2
F/wRG04l0Ynb72gJXNzJWgtypZ6Osmup3QlQgv3y6q1Z0irMQ561z+S6D9fraenq
yQLNsEPQ8ICBtHdQsRMIUUlmeOirK84HirKvaPZjOqo3I//wRwN8RiRkEVi3JiCx
g4k4o//QyelD0UXbxmlwpjbY4qo7HyzH7xNyQcNIzCQZ1Uyp+iPVnGk9laz5D4TR
6Cyf0nmg/rMkZgBSBP987vMf7pdeuxCAS/87twnQdbUcKVt+CKZEhtZNrQG4XM8z
vUyUaoPxd7Ds/IYM/czPmZnzRcneV5jdSlx6IoKRUB6P/t9BEbb8HPmQa8uI/c5o
8GAXG1dNagBHBs7miF4WE9VGPdt1fwLBtGExHwTU57StNCsFZ1/HgjqaBfgkUeY0
MYeMwp1BHpldwWE5Zwes/49BKB89Rj9LKyFXpsCaPhNV2EW5xkkbO1gCWjGrQ7oO
bAXsOThY9+G5QOvGaQolWpe4AWlB3+qlXq/BOBn2oQGcAmidPIymtbuIlvQ4LviK
mYUKNlMgj94KVQXTaU/RRQ5au6fJ9KX25UuB4fVjgRa3tE4W8/S0/H09HUSbMDt5
n8/abGTncDuhH+/LpiqvFLiMG537WSjAZXS3UyJqEadhNKZ8nF8m/o3Sp+S8caAg
UK+0K9845CnwFPfL5SSRIQVXn28whlDyG9zkHYwCzPjbiFIFrnX5/vW9Caf+MdXb
VPKLI9DYFLajWTPfhjinCmZUdhJvBMEZq7QAetayw21JgOWHNq0J/q9ZV1/v2VRg
VSjPPXhUEYWz+uEBCGFi6ayv19vuujxvei6SU9JSOjFKfjAO2/mnORu5kmzfQjda
2j8+4SlooVoEJuwGOk2zamvhJWzz71eDhGlyGRQiNgZVBm7CZiZDMWW0pASw7kK8
iRR+omNZ/ndPQMbZxTqOffq8f8WcgfZWAcBwnvrtOxgpbkJVo8ZLBRxSLSoZfS4O
yjrN3QLTbu/aKpvmZlUeTu29UlPTlvpCjrbm+MsoyI7F4EyvD9Aru/RJfX6kyTpg
N3tMktTXHdfL3We3OGlWoPDWt9JBPP0nsLzzBW0ekoPgl00YeOnGEDuSPxdhi0a1
7wAnKOkKcd91elFl6IB5ejjDQjmOkpjysntwZochX643zEebrnGpZCrb5HCXfzJO
zkVSTgD9i9Yee35zhJ2HPPUBRxT41G+rD9pofsFLJQiqHl1gpRmkrBQvpkCMToLr
lSX/aZSuHIUpJKivDq1zwtEXN6o0mMVeGkXkhtlVydZIMPisZYo3691KgCwl7G5c
UDazWOplvyeeBDjSt94OAFVeNRqNyysIBMx01/tdUWj+w00FXo3sdoVVtvIhgpxv
uRFhdi6xJKKurCGt04lvURYpONyqXh3YsSCVMh3+U51p0rQYgkW9/LC4ND9Suk5q
6sgOAy7mtvKyGQQrgvO+pqo37icIUg9jDchzCCSs2jqjbA9ecOxHVIA3Gyo46gvj
t1O6vNduHJmk+ignKe1YWkOBFzg/LAtFKGskhbnWQ8J44ZaUnybmVx9e/w8jcLl0
kZNApLsbMTjNkjPI0sYRJ79lwYv22JebRPa0+dHs47Y/GA2bxY0Oyum+PNhwTh+l
R12dm8cNvVohmBTXjLvwX4auu1KZrK4a6FIbuUunPZ5HWSBPV4hnkKda3/vRzXN5
a0Zwp45B5xrEcSjcxRy0JSMRS5mICcaBCItJ+kggnQFY/FPQPYDz/z2wJblUBYjL
ChMddDI+EshMRW+sQITlTnHUhDTCF7QCDHeFhCXWSU6IJu1GnHMrJeWm1lqWRixa
XV16fcP+MMif6jk/0toBDwI9X6cMp2AU2vcQTxxt/hyNpjV4Iby+DNPPiXoqNSI2
+9YBZcQh+Jz+RxQyBnTuFbHsiTb+iaZ0UjmwnoqgHO84sJErQvj5fjNMJBrklaaj
iVrgeJOiHHfzWRR35DKHo4RGFnvArdTE9h9BgpJ5zsx0gyjnbKgEbLYkZloMwIAd
8AQ0FltSHm1/4id+pPFZP4DJCTDBYXwbFc66jeNxDFepNq2NziMUVuB8njLVg+4H
aHP+oB5qic1Anfvb+CluEatYBpimrGlUJBx49cwynXSzB2SXmj2UlmbZZYuob9kH
wDdGuRvG/dEoDlV1EAaaK29xNXxS3/6XFcZpQKbylDBWhZzACCsw5vFrfNZSHuBf
GnlSw9JsWE/dquobCpsBynKwrhxHBVwAi6dWTO++PrgBtcNUUnnqvHJePGQLUHCZ
WeEs8wAZCe7SxtyeE+nKnQKgDUVh/nytP6lI8waSiFvwWI1lsJD9iepEFxi0NvqU
5bgTZ3NK2+pyOFXfH91OLM1sHpYEL0QK0eHRU/v7GclHrsQx6ZgdBLke6faE0UFx
s5HGhPXJHTFtF6gUS8jNdlHl/Ae5CVlj/QLspQ4MNg142KdOdkaErfUbi4Vik6xC
3jJRx13NRDYmLeLjGHxmnnCYWzYKTuxKS7QeKNzD4O8YJTCl4Z3BsEyqUGU6eE+w
T/a6uj+oQF4rXOQpgIhiHlbBAOR2ozqmkFuC0wyguqNdoORRhiJ0Zx7hdsV4OSSU
LaR1jfo9kfy1DmGo8/IvsQ==
`protect END_PROTECTED
