`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JkQw3j4QBidVhYafn4TENjQ4Sd4O42Be0j4OeRXA0hbqMXH++3/g/Bwc0cmMtJpO
R3zxTh0X0E6gCcy/TShb4Q3FtIwsvXWbKKYIainJCaoWobNSqJqgy4gw4x9SsZ1/
/j4L3G4V9pYRnO/FTeA29e4qWZlwgtEeX58NCTblNTee89zVDOVgx16AD/cN9XXQ
bkLgBg3busEV9XSsJBPlRljOyZ9dHiW9Tfh4JL4bgq4p8qxR94w6l1WCpR8M15us
UHZKacYOORh8FudZiBiiAlXqjtFhaftGLXPKX1NOcdA/dksS1tZGJzfa2bJ6niCX
z9OSOlI0uiEngtDeRa0gX5fhuFzHydGhJEewE0aABi/Z6501BLCFRasI1NRRf9j3
UKCN+xvwbGS/52bCKjqOz54VWlY+FY3jD47/vYDXB+uAxdo/pKsPYjZZ+iJ/xa+x
Rzki9v0riSNtlvk3ssPfjqwG41uBXpok9lfFaeGgb5YI6nmYqZe3m1yQKrwwo0F5
`protect END_PROTECTED
