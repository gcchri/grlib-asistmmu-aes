`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X7+2JyHMA90cXa4Civv17QjDY1HWJYErI72IRbDAAtavNsg/wAS50pRBSC+FT05O
WuC0G4xrU9mkgN+pWW0IuJ6VtdACkP6pUurCzsjoGRhSEcXAUrkL8kR+0v9y33om
4JU10X6TJ2oxi0S4PpPbJuAMiy4+FsmOWJVEshEHsdS3nxYmWyK/APrthIOXyxh1
VlEaKGuK684Qmo9XYbm9k3YMwwDnI51DKISS554EFJnydv3ojkIaKL8PpG9342E0
SufffiQXpGso+PP9MUqCqdVDkEGH2HzfDHnlzd166NvESCXsA9q7AZa6KtT7ZC8S
YqC01Isan0mOebpll1kJZsHoLTfDDuo7f/3lTrnFa4uGJcm8e+3JuiJjTOo+2jDZ
wGvN9RDi4URVWKZo2z5ty9nJA5qMSvZ0VX7PNna3Bn+YYi1YnzeL86ZcSFBSEkVv
49mvpre/WdubG8yW2kyebw==
`protect END_PROTECTED
