`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MbZhw5qM7h2fbEJFg3YjjhVzQlwV8Hl2bQuPVMfGJFguylV827FizReiIQSQwGvV
Y13oyyI662TJaLo/jxwnUHPzzLjsZXrrKvK/u+TYrz0i8Yzj0CcxPPxHlQW2Aw8S
tp/XEzdNPWcyIDQhgG6Qh6pqlxYaRym0OwVmjwRaVH5tU29n7dSbhSxJJ4FX9HZj
ZsTKKThPltKW3KLrjP5a4Wz/OEBUAVdKSUvALnoHGCdZpc3Sdy6IH3GmqqahB4RS
x486uQ5uaWaCfnLgq8ozJWBs4zC5lMIIHhDPtlrFH8Xh3Ol1sZsUeFxjJURV5FpN
JvNOFi7C1zHXXZpiTTcC/w==
`protect END_PROTECTED
