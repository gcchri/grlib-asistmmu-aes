`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ovPZ+2tV9uaiwVAxvGKUKFlkUU1uOPdYLz1gSJbAFK/LDQfIg/buLfxPNXmKwi1t
z0u9EOznTQmYacIxHU2x8sQ/J57wdk4F0kZ0J77/xKJXiQJh5L/kPVyiHyRRPXre
adQCr0ntzz6nSFjQLPV7a4m0Rm61jUy8ofHszrk9em2HpHWA4MqjMCuo4XUInXAl
nXeHWOog8h+5LrtNVrup0kKw4RbFHLNacWlo5yIhDBuvbFZzgjRNVMrIk2c/mRSt
I8z3MFhtEx50GZcfssxsNq2ZNgNRqULxlPsEknWUwecxJXzfMEvnYQ+K1l87zTK7
K5fLug3w38FlOjPHiEsjXz6W/5zofnFWQLWM+7Bw3xITcbzBY0kXgwdCdPtKv+8l
ZoDmocoXHX7STXkK3BoqqTZY64m91PNgnu+A4YqgLI684lsWz1w0xDnbXatpvlnP
pgMw09sja0YfwbhqaOTr/trwsyDjAPcuUBEPUM2rKul8PEX5qNcujGhq6RLfqk4m
vUnGknZ7qOTPR+qfVt3Hj6IxuxzcOwF+m8wJlADZf0AJGGiVfPXecREpP9TRtZLS
XuI7Cp1nWsy+p5PKgQmoAi2bhavk4V25/UjaOHm+nXrJLB35sGlCUpDWFEYvI3xY
zqlXZyiLQMD+41zb9g+DcyhOQ4E5f7Evy4WS9BdzsWB9mISCZ2MIOyLxka+KfZjW
hJdsPYU+b0DADwjkFa8PUFav7Gw3jNQf+fbqpRYH+E6nyS1Vf7XLOxTrC7XeDQQW
K1DdlNaoGrq4sf8h9ToHczMHezEg2cRg/PBSIRvZ2UX/an21TVr5OhpZRXGNU0pD
+qGSGl/WZKhTdHGKIgymtGkBxa0bIIdn7SQA/ykWcohEEixuPY+wx7toGLHiN04x
`protect END_PROTECTED
