`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kFY7hAcnS9yG99bDW57EIQP3DUgW0DpzOOYtRV1o/7PtGiKM7ofH/8IUoDD2+QFZ
wJVcRKXz8hLl5aqbGlUV8B4rTz5FHccZ9wIQc3Yp1M9vzeYs0CgBy67fCk+dwwg3
Bze8WQ0sMdJLWIHV4iQSb86zsYWgihVrTB2L8JK2aHZ4NLjb3+8Ah5vYUWMlzvtJ
TmFbP4aHt7UsILGBHNMx2ynB2nYb1/Dexk07CFsvlTxv3b8J9vNT3UUQjBspWb+2
ZlWvAcRC+sSwsSL1EtThhsS5RFoji1jBDpux+r1Bl73/20C02i2dK7Wg/vXRGsPj
goCHXVc1M5wNibwsiHn/1Y8fURUSWeyNXxb0YXGuHiyIkFHw/zLixHxfL/Uop/9v
QjqP+VrcL1+eMWRgirilFGvDCw8c9Pixbl/MHVuCOzeHB1/nTegTTPXAZXTXISf0
kCbGBp4IfvLvY493gFs6Jw==
`protect END_PROTECTED
