`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UDd4vcurG0y3UYXvQbVaV3IL6flvP/aka7+2cXu0e7eqHvZG/urmMTrzTxG+7yP8
j/Eh+BfjZBpVGbbLjdMY3Xh2hR7LXukvye1rhIytKGfN00v3bsbbavVUYtSPay4Y
rLPixORKI5Df8RISgHHUk9cEo2/2mYWLzqYE6p1Q+9QgcHpvlpj5Mpc+ELZEPZnR
F/EeTVW48GWDNwGEuabCIOmKPFVE9D/RW1Dle5IUvUw+pI9JfWDeqZuLqelQkoJg
8Wu6KdrEsAf489AgkW/09rRjxnAL6kaRPNpFBRi3HkrkWT5Hds8yq4ktLoPj4s3H
3QanlDl5rYpdjWCQh1qc27ZX3MNF2GaS/BXBum0fliLT6GeoFc35yPgZpJ2wHnG7
3Nhm3nEASyZ1bj38dV1oRq9a1ODpgGLdbfN7E4Mf4WOwKnattaLSXDG5wZ+4HnKY
js990LlL8i0TSH3HioXGPXmotpv8LFzBKOABAurUswgK9bIdthewcy+Jnmlt6XUq
fgYAVVpk3sCVEwk3ZnJX81KiS98yOjF0uk1JGnu2RWn/XZacs2B0RQuTHU55A0wK
w+AVKrzea3vjX7PqmL3Pa8uImKEif4w87t+MUskmxn/5F2rOSUXmN6XbNQTwekAd
wyCAg4wTCPmPwxviriB7lYCqlQTlKfaUf8wSXhcVcdO8IR8FVO349nggzKf/3Rjh
TFd+TrxTuq2nNPenNCjwuAZOAfCg+MzwvQYNlHUlbPheS+5Ry0A4zmyGgZGQiKG9
LBLnxcDUMLUfo38HzP79WjyAxRLA7chAYpAS6vlZ+KP7sJPr8LNIkJJsxt9MLILb
zr+HA7GN0l6u9usBmQg4fOw4z+wtyxXpkefjspB3oos1gEzoM2BmNRUI6FVMRqdy
hWx3s7Swv8ixF1TXE8PI5nVaydF02uObuiB7743pfiVgQ7zPRn8h0mwEClnblHiI
XO/0d8S3IOFbm8VysduHZw8NiB3TLHIc2P3HCov0XpvLMhAQZfY2Yr7eHTbcdLTR
aJj4eBwaWgZRJhdnIoiw5hqz7gvqYdkRW/xCTC1lZZAMfddiXMkgCMUCalba+66I
xNHSYPxxa2uQjenaUu02IQCs8G0Byl6LGGMEQpj5VXcppXIKz8hNS5KZIyYFasvu
sa5/pR33X1+8VBHZpfDNcsj9eh3+xHmDvWXAhe0/J1Yi0qXCRjBFvrZUbs2FVkBa
q9OmjASqwcuw3QwJpFGUnnbwEGpaimLNKuopfqg+oCYlgA9wmaxug1/AEk423xZG
rp9wTpEZVIWBDhuyCOgtAoo5lLAVGMVkqDrL1slc3OWjit81r/bNUqzbh67vIxLq
mnz09NpxU4gcxShBLnIt5MMEdksaQ6MUwuj0uE+N/5nduUBd7V8K81CMQ1NiPRvp
wt4OfUxxCrVfso8o0qr5ZnYRLdkNvtz+N77QpR5OM2fHep2yZV2IMrYHn5h+WtzR
vi3De1mcZ/m0S3a1ki5tdD9hi06NYOjygL3wiT5T5+CSF7PHZcyKphBDfJmsYif6
VMVnsM/wdZLZ5xL4yi8HUsJfZdOVWzN5DE2RGIsyIldhbZHp5xC/V6Tl1CVgOstF
KR85PoSaIuwRpz2iSd8EFFL+HlCVJDPNDdg0tmeRZvbR2oCgj5ZV4YcEcJpS8378
M/uuDqod+rnanlSrtEH64JF36wrdeUtloHcmOiuiwqYN8VNyfzOEEpBfa4btysbX
NcpsoZL6ZQ6Abm4WGWl2QAY9qYdCXsj4ko7qIazwlLqpAHh8RtVU0f1JEiDfW0cs
aDWfTFszS1a3sH8PugJXjvCZGf8jGObwl6UUF89M5j35BT+6vonu7/GLtvK+HnH5
MR6+FHQhwhYsYpJTO6AbmCPXQa91SbPEtAtnuZ7aZXnG5+bFECVOye6VIr5bZ9kx
qLbnnEPKruMKQx8iqWEnBgVB4tg0nbMi+jjFCvG9AjSxuG5cbX2yrFefxy7VR9WP
V9CPPm4yC69NXS8mC0YiUTO/LHCETsuW2WRoiKQEkS4VeMlCsKIIjlhW6Lqj+EGJ
yqnnMIMbMnXJe6YVy1aW/bmRNJuTtj9S8NgP4UoQM3choRZsQ3LY/u4T0Y/mj6Gd
v5j362pU4VV61cAWF607P3l0ArrLGKvXEYxB079kI1IsWqF7BJHhZ3MuwWb1zfLv
pADMttbgC/P2B9dZZ5CCrSqlCodxGt2dQ7Asf0uEm492GLO4UizYz+MXVpvSWN40
47RL3A3bUFsAQ3cgX66thJUnMBv9fr9yQmaM8wMcc1jw7Lbq4hjmuIZluq4bZBXb
FSoe7NCBMHjk4AbbHrTilVQbIBY2K8tmeKS10n2onoTh0G05nQXOb8fwtusZsOfC
Sb88yKtd5lMMbhQoNvajPeMZZJYWAH/9kyxHveSp7aCPPRCD2Ci5jB1+1R71XrJ6
ZjuTpDf5EnS1X83ftsd8X41r07fk4f+BNkbJchlJf08qQlycrNwchlH1uDvGqrou
NP1qqnH848P1bDT1+3GMBrxAiANq10XthzJcKv4J9vk66IASkQqxRdNtqSOhszKp
n2snonHYY2AGkdXjltpzP9SbhGNgaXT4h5p8KCvkIkMw+SR0ZyuhkH2MD0osHptb
tfcaB1VCubqTsHp7S720RL1kfDZ9jvKrpyxVYVHBHk3jeUjKwMzF3aMo6kvA+nCc
04BvOXuaYROWifMrcDrT84inYsBqM3feU2lbn6KR7OV2f4E7PjRQhCmP7JKc7N40
s4AuncqtfY5fSzrf6VywxtMMUvLQN3j7XdUktvtvYC2P+LdJoSqg+XIyPBpCVr0a
J/TO2dR1PMjW075wxXW57qcBTRFzAocjhEQYHnOzx0QAMqvDknfjmtlRB8Kf8uVB
j//t3x3FYmJmy5L/Hd+YZlpqxbqcX9aReyHmmrx+If25iItkVnsOBV+B/cOLRR5g
DbEHplOBE8wbnjz4cGvV24i0OkB9fH1hDz9NOzMJh5RKFm7T7s2D6C36FE5MKM+m
L1IwXP1x0vmigLVLSpGxnJ8r/FBIUUR5FgjVVYHdb6o4SyN9sPc7KlvRa26VW7dF
r32kBBtKxK3E4GoEcOI+V8oyPxB/9FnXOEVZDnFyqOobDnTUFQXZHaQ2iq9DC94u
Rls4LNFMMHs62A/VGfDnyKvh+jq2SzlCAiwjx0QNnujKT7qPHMzmaxnV5DIrjMpF
aifVIEF8o6dBkK60VxCsWohfQOcs1ElOFflLSx7Z9W0ilFl2YKzql9bOEoQ+9psF
SCF7w+1N6YDNWBjZ4ScQFXxD1BDdnDBXpz4XG+TTBOLPy2xHiqXHX7U8FHRwU11S
KPUQAV9btgmb5lHhQl/HBAk0eyUbk/uQjR/iRQMS3WsWhoNJShjSXRtNlNbYQk5r
mTBzkQgv4JDCVHhN88BiLRBN3O39G14oi4Ca5cVDGPesW8pUPH/0kGAw7KvtRtbO
fnkjByqDoMlQcZcNvSaalQnpAFNn/ZFHCVCdHuDbVSZfyfaQYiSjGxnGmi+me+Jq
dlCVuoPRdWs+zoXCEvnc2rLZDcoyPrdCkmcbBibGCP4=
`protect END_PROTECTED
