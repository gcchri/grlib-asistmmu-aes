`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9sHHG31KmGbXXLhV2yBMqKciQliwBn+31FJvEyBqCU2QVNO1fnQ9gziu/sYZ95Fr
vBJTZUqdzsksswJhONa1V2Vg5OzqPMnGiHlgbE8IBq41W8zMZEiMiQxH06l/TxTz
k59lNgqTVvPF3yxDiIguRGxkGhJA7cpvymTkLv2CnyY7X9QeSl5n2kGt3zcXkhEn
6P6P1z9TKuL8VLlpYlYze7G5cRc6CAQbWQQd5bxkDI2x9fKXc3Xqcfr5muB0oI+n
Gcb2HWXyb/pOkVNi6pwHtg==
`protect END_PROTECTED
