`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sL62L9UMmzB1+sPw0oMtsvcHXFCTMmL7udtcRKmiizgTtPOUTqdq+6EpvEINgBjn
A661pxF6z54/QStLiOEHD/bcNJqoZM9JC1pSDaP1DJ1C20TCAw7NKWAdhkLU5L3C
WrgHIx/qYcN0UAGGXw+nlImcw88ZkfrKa5yNsjM8D1NvqUjcp2uMscgWrRyd+Kun
0cPTprEi4wfHYomDKyUKIDwo0Pe2gwIomEhMDmBrqX3dxx4K6tbCuQhoULjJzw8n
5K0ZoNj+8/0JKU01BIqUkEIXOtc982kKryaqIM+EevrWCAqV6d9Gme/EbLZDNfLq
z8rMyvks5H0dM+Q27SS1RR3Rj7HSakaYQE03uoYM1uOc8um4oEt91EG1S8RpaNH2
IjRkC4M71/3EZ8OKPJe0M/TCPrDBE4JlAx8vHqo37/LrqRbokc12hHRkVYJmiaZy
`protect END_PROTECTED
