`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+hElH2goRB5N3xuPEzZ9UFtWCIEvKKy9JhEyisAzprqrBa1+L0iRhagoHZd4lD+o
3aLlposPZNQM5q1EEFhvd+oI1ggNGJf1dS28w3nN+NMq7N0KKM3r5qxcCBRLVMRa
Hlxady+N3iDhSasQuYId6Jw3yL11TxCD0T2TQyboa5IJPex/+Qhe9uH0vvuyBWR0
Bl4fK1HU4Dy/GR5lTZDD7pN9pu+/oQQHC6WOwYJUXAUkH+Gt1IyHIjc3V0RwoOWK
iwvuvnRkGUCHJDfqPa0/E9QFPCA/2xqA19+MxOjQiogCeZXuEliZ4mEenHEW++u5
WLpbsveNNhBgtuhwlv3b8vKxmMg0hErtAdw5I8VroCCWge9dAPjZXGHExz2jz9jY
k96d5ItMj4/2sXl1VKTv5iwRTy0IlHlAp0SnM/a5IUpWRgomTrHC6Laxkm021VB4
CKzxAbustF97RAz8zrb4wWU6atxvTU9im+ow/t7bfZW1lqpP3aaEiTvK1JnibV3P
owcTZlD83IQnMXZ1xILWWDBCMGgBkwSKWOASU4yn/qr/FyWsjA45E7oCY3V94Kyk
h/IC06qVRNeow9nFnP1fi+K19FfAm7+9NX3Uz10UzgxaQjfATktV/RLIr6qYu0PX
XUptoq5tXgfgYWqBoMpVnQ==
`protect END_PROTECTED
