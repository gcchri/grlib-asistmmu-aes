`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bsEyGRTsKJOecyHdYDQalhZWqbx3FnESQh2xkONbwH1l+fYI2tgRuulFfk0C3UGw
6AN0pyc2oW8+TNZLQVPbn778LP3WLzwi5uLMOnOWo6eQ/Nf7lpaQopWT/uVAgCyk
uoSfUTSf6BsIbIbyISv5WJX67SfBF2e4xFqFy0POtG7yq5tD5aMNCVtLn/qLjAhC
Nhz/oazNXlmuH5uoWe3RGKHjIE0k2Cx7gTJaIVH+L5KW+15ZDBykazGU4HAth7y2
2OwT3Yg6qQvAbTXed0plmw==
`protect END_PROTECTED
