`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xSG8WRkNoWsLHFjdEgK8NgjqUx9N7BesJxInut+gNiItDFIyIAhkUgCGrlb1iiS8
wnuepH4aZGf9B1PYMs2MJGPKLiC7lxD/sVQrn92vu/cliQtvifju8U/6zIPj2pv6
umBkvYnC9F6E3JrY6TW30tNHqDEiwnhzq8052O1R5hy3LsPXtb0i7cIf+lIgjzUY
BDZj19W+KctWvimIiK6tcIpl2pnEgFFNCjwaKUbZUBB77Oez1uGsklDkSclom1pr
IApu/Ov6kzXJ/JhLFGoD7FxafXGPE9FqbDwXsmjkDRaMYtGoPZivrT5rdL+QVvlg
Hz70HYRa0sTjW39pfR2d0YqV2ElEwtc3/MZq3JMGkB5tt8i8HZTGm/6aDPDKzMBj
GS5sPJm4pkWQSGlTYSNXr1TvbrDFUjphS7BlQGZbAvM=
`protect END_PROTECTED
