`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7XOEIYZD1Ft3ZR65FjnL7ER5Esc4rhXAd9CeeZNVFfAECP07SBTV+a+ssNPBf74A
6l3XQn1kr2zalwJ8QjvvGp6i2i9dkml3giqAmWr7dqmIEXEruhwqwWr5OlC/m325
vp4cu2CV+H9z9CM3z38mtqrzuQ9bm5DcoynGM4yRdWBWeSu0ePjOvd1GOUwNJTol
k3VjFnR3PXOcW9EYRUGNwVCQDgrLdlzF+bUtJcxxKzf3yacTFoB/ApYjo7C1aG0C
Vs1nR7qoj5wZb3mWQtClMBNRZbetN9n6/v3ZcJTemS0=
`protect END_PROTECTED
