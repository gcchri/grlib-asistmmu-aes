`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hslfrx87lCYzbooDnuEspYz/LLFSp9Ye+SLovz+ktTsSm+jvPTZREdwbjoPvs9JP
08wo4VIDIx3TAWN2R1nDZQnWvAmMz+aRRJ2Aj8XsRD/pltncjtmOkSfF0srnRuxX
D7+NlAkUk/rZPxocOaGKEdpsglYKO93JumjGFxp4RjMO7FxqCVNtIONwXUGnqf7U
QvSFk7N3y32PcLTQ0YjFc2MgecldTBiBfh0E8b5EFZWWjUfh9AXeZh2HRcUQCTwN
WCLsdIA3tD2XJC0YdtqHej8q0iJq9gQqkSkM5xyt/89ohLT6shrfGXE3SN5S4LGt
Saw8ItCMqsEdyTHxSDvoNby7FQbL8y93hmf5uSSSpzRY7PyHRUGQWUIPS1jEwNh9
Ev6Y0wK5PTEIvAy50Ph0+Q==
`protect END_PROTECTED
