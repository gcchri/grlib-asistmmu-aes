`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Cn12z5F2jfSxUq7RV3TFfzmT8ZAdfIrwm4a+u7Zp5wYdkwJt6wp0X8XSTNLHFhX
mw89TPYhAJLXw7/vxUdz95mi599Tj/ZaZL2ogqp//hIcM/Ey1yudWjE0SBa2y0td
EiMNycO5luQ5or/zXum8DUCvQ7xFfvzWwabuVd0asxNmT1HCBbOKPkNg7FcTmSZa
pSoE1b87moVkx1qqPKac0o672kVzqlvNhIuWL2ebvIh1FsZg9yjFLIhS7hjaY9rl
pZL2S0ixB3aYFgVQv6GJX7AC0fB9rXwpGKex/+roiSvlMmZwGVjhUENwNNu5DCqJ
TTtgBgHZDiWJI95w7HVk8k80VHp2rq1WgcF22GaZg3UOqnqKi6QyfPoBpYCrRTI9
+7P3NsK7QDXqEhTavt+DN6rEb+tFeTtx+1cJMRwE2FOOsE8pZSA6HuCwwB+vXMmX
5rfbsMCfoaQ/ArD/sS0Hpw==
`protect END_PROTECTED
