`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ahiMJzdlnf7Wsni+sHMdQRoNNad3bhqscvIu7bH4pVubdnzQdKZvm5Eg66KOSnKv
1Klv2lJVVZ+b9QziQSceq8vbxJ7oYh7gK8v2kbnyW83QX9BK86018J+Xi9l8x2Db
gRzkWNL1dWlJwkwSUDmDok5E50g7NCd+EIYl2hq1show1avffXYYt7wRh/Y21nLp
LTofoEN6irt5wfRKO3G7LV/zqR6c9E6s8nTzMFR+8caGuHOZq7sRk2LMrnW3u27F
+eXXzH73+K9oe3mN9utFxD/QU+XcVyHyedswCingiHkZd/vxA1YlDvRTaNu3eWAg
kmOrkKKrW1SHaYLcyGckgA==
`protect END_PROTECTED
