`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6dvUeDJ52KttdVozZEwiV/jJoudKhnVDT/kH6Vsio9mrtJM6ui2vj001gqCuknfm
RIyBzLotvPyFt8xjS74CwY8ejYpQ4GfBVSyz+1aRg+bbK2w1jGKJa8DRZu6w3KLY
NTYlFeY4GbT82UAhjnKi8MLSEH0CkEl7tSK8srQGVfwHHu0SrbjHt61hks7h9h3f
efHwAUa0FEJEsmeFUXlg6B2ZovnKuwBvDzQGit/iSyXVLlpsUJFM8rQ2kB3STO+4
JjeA/ed1sRcBB/qdJh91rpvVaWw+8v93wySd/72RwWY6NRZz6SHHBVt1CNeCNa4p
xas3Aydn9KmLpNCgzmPgAmFULLtJPxqb2F//nj6LQAvJMu/AO5gmRZha8MVpnY+Y
A+3L/XG0Uylx62a4BkunTu3wrZnlB5z8+QkegJfwIqYNbBkqnzVMVByQa7PI370H
ws4XVbNYa3mbjIKYHa7g5Q1oUSd0WDLawaLirybMi37k6G3OYDNJVlcZ+9NcdX8y
E+OnF0YBzOi4HpiMzvcu6cUMGjmB4e0rptO3NAzY6jXgVdlm2FCd65A4tN4gPL5r
jA+rA6hqynQjEINHCecjx73viJ9Ysy/FtdrAXzqh8HcouWT3fLsWbssMlp4vwG/w
jXDb8UQKu51wPUwjgI+PJCgw7uCki/pYZn+QUpl97IfoD7gfDcCjUNPBWcAHi7vF
T/8E0+t3SV/RYd3ldHs9T6WceShqXrFQgLSvaf936z4CF34s4IiShkgMzX6mMXY/
Q8uKwDO7B6g3S7rpreMlgdhD/bc/Mf29v9C5VUQXLnRTzasxVd6aqq1Klh6v57jg
HJiuqXMjRQKTdhtf9JTJd+hfQrFpjNJN2VDmYzp5OPjfhpmS5/iKidjzwvvRROkv
n1YoZNq7GlsIJyWaUu6RBlBXCndcDhFov9DqNLlb3ShwBeIpQ8M896qu2NWm0L2y
`protect END_PROTECTED
