`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ozpzwaKWKhG9GhNz2D8tFel8uxWHd534Lk9bqX3p/3CjkrT7Zynv3JbiyTgSzLX7
fHDgTVxUs/8uNsMUDMzAYxO/pdrhOGL47ZKn9N+Vc8feSsDM1nIWbjfIs15DN9e8
DjaJmEIP+w/aBR7oQyOw0M/vrO/DdcdkVFqRQCjvzuxRRHK1MBTF0rCAXW3YcvrK
jDOqY1+GluBSUHlY3zzenNDEVvhUoAHrKE6eeyAJ/yN0C3VUQMP/IJBBB+RabUQ8
vu1TKSa2BOMPS4MPxdSwTBELdzUrCay2A2yOEr4zaPTm3wq+wKsHnNRZtfhd6XgD
XcTKzECYpX2o7N81s0qx4pwUAy8AsUjnZXAqaqe5hNRQok7gndY2pk9x6eNkOQmn
ZUJXXfQjj4ex3UEq9gzvIDcpgru9pNJW8Ruvpsi2Er95kcMait15YAC1TPxK6iZF
mC8oD6FWaudSZp/xBJG9p+h8MZnx/pAQSwCM10ix/xhEMbpACfg57Gxeah7se73s
eSzTMwV9b1/epKSB/ZkdpeoZGLw+JxJwsHIdxb1pX6QmD5sdD4dBabFlW3+1k7JH
O6zRHrk8J/XTbQXjL0Om6uGmy1VhjhkXBqE1nO9onhL0NbtBpRVuxfvHRAqOkAFO
BKzTMucCgAoMVMCZCqODAIW6AuDaDXBprC9MJSLA0pnUKZm8f/CI1GX4/o8idQJR
YAA9QfKY7kMFCx1h6If2ZojqtJ6fmOcbnOWD9gKH0uMrYBEYlncGGXfxva4DOolC
X3VtioSFh1BP98vgYjIQIfp2r1QetbHfJteFlOKWyfSx5M72YLqUsgClCUv86LOY
`protect END_PROTECTED
