`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yWPIm7k9+8f+j9OS3HSHHRqdOzkekZqBWPs2ed9IM4X3QYIP0Du0XrCeA27fpvOG
cSZRW5nrq8WU9+Fa+VIjk9UdW9m08x+ICdMUpURRjCRS4j66bdlQ+LJPtioZp8tQ
wiqBI4QdFSXp+y67VEVlr1EfmQINL1SWO+RNrE+ghZ98SngaKbYEdrW3UpsY6ADy
AHKnVfG4PPGtIVoLFJNidFtT+IBg9TnsaWsrWUu6H6xIdgntyXv8+T6ugjv1qbBj
Fb6qY3em3VFL6uleq6Nxy5arU4MCe4wNSHnwEMIfWnK9D8BKdYpECRPdq37BhDAQ
cxVUpYtDk50UpBHzgq+livAdppXSS3scoceSTJuml4NGnsJNeKZPQzVtf8pc1dq+
nLFQ7o0LqHtSVKHE/tF01wRbLPZ+rOgGM+uZjxiLTc31Rk9Xlr8wMYGc2svZSv4h
fPjNkGb4yIZR/jvRHRt7dFV6XtE50xFgPczuBZ5vaV4xFiqSzOcczZ3mp+nMtWtY
CEG0oymvhD16nTCdYu7qp1pIL5L77rtHO31aDLhd1OqyP4wlFktJjYaHiPrxlpQM
HBNwtnZww2c+piVeWU/RU3xZHi6HcMlKTgt2dbstjRGqFkJHYMUViXPtnpFUwGWd
WWTdvhCPViBaQ9odceDtuYCheD20mCeuB1CT/iuGyD481Oc7y1OTy6+iYeNNiszx
nrLekIpcF6b+ev28OTD7l9h9ciNKsTALWhqBVI8T7KC0Wqw7h74uMI8DfqPw6nqb
7SPWE/FdzbZyTr0pSVf8HqTbtbVfA3hC32x33Z0iaSC+R1KRX/0itnWw7DKgvB0l
tmzz36w3Bg0CWpp6njOj1DCPF566IM1GUOFxyJrHqZs=
`protect END_PROTECTED
