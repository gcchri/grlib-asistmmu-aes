`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iM1t1ddtfjLE+3Wau/4n2CMqtd26Rf9tcXI096vwEtlbw8PluIvZNN+Xn1OPGUVg
UvI2ABBP8WPkBQZX2doYgSX3KM9rMoFsWuuxABIOcMPfWH8/3WhUhCWBhGLnHT/b
sMUgGOX7hpekrHi32GQKntu7CBX633eC8Z0giJgOi7SqSbKEabrFlCPQyLkINKaW
XZiY7kDcABplyuL2VYTyLoKCS2ppDxXd8yr0D+PnHyrb93nNgOM6TYfWnH0S++Yd
OIoKh2A7asU6sn3QqLCSIZJQKMsLhDqIJsSroboH9wL+5AcTZiGBjMbQ7eX3ctCB
um0ze0ScqYVfLO7nnY2hKdTy/N+4H/HyyrPnd+ARLF2JdJeHSfpu5iQTd8sCvMDu
4JZ5suj9HAPV2SJ0yobmg5MmDv9ej6vdzQw+cEafgz38h8rPEf8VqyO+SVzQcQ3b
8FLn0oD5A16oy5btdkWW9MwbV9WmbNUFas7u+LnvNb8QktqnqqdfwQVmsFeAWo+k
CDnY15TfxZlgELInUq77y1jq/IjTY2T++jmGS+PlEK19cjVuJw70IwZU1B2hUM2w
pvgr767G71eQDbqbVdrMxQ==
`protect END_PROTECTED
