`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JSnfxKRSh2D07eDCfMFrgE6ruYFvoPO/8R5NrpMIztZPt//7pR5BFQNG+k7yOYB+
/dtUTGqQXXGdwEgovyVAoTpWY/IkKDSe+0wjpqTvntwZ4esiUVeVo7kfjeNB9d6B
u9M8H4aGKvzXxeduNLJNtZaq+VNMASimAZLvr3wxFcf0Mad8Lk5ALOsV/qiS33TC
8Zb8dEhrRuBBwrVWzOgAzWL7GWBUvtBcQ4WRfiHMPjfBWuGX7VAoJ8Fi14ffl0rG
39zCFNRESLQ0hmGKFRDFk1Q7PqLCsRfQdotG+V7x/s+b+F9aP4LGyrs+vmazxSsW
t5FV8s8q0Ki+ik6+N95rE41FfaD/V2G2e/nMnAknXcvLDKxyPuFWDzCNyXLtImGg
XtOvCFsvDZuntyQb+bR3/uClEZ3EaRSlpDXvohJfWXJvTxF6fRMjxRzWzfRz6jDA
/X7wtPXcw0XYVFCvJPozdnTN+N5qQw5b8hgr7w/YA8/nrF6O7o+cKCHm1XR+YAPI
7HE9hRhPN6i3B63eq1kr0Y354tRyOZR4FK/V/Oi6KyIV7MXVSYP+wxfi3fHWGMD9
hmw1CadPFyNh9/dGbQkIhi0iwVDPiZhEULFZTWBmymBe62wMOd2/LIllKLedLtJI
qcYrEhwBjN9y0jAAHT/NFXXTeJBfNn0hAwiDPbhdOmtdsxwbkrJWjCpC+oIBk/FN
wA6oMap/mDXO656l7RkWFPnbrYmw7njidbxKlTClCaAX5sI9ifiM57/2qt6RVvAe
24CAko7njpcKQgxO6Gato7TZjKvGMVHREFdATsCrGN4X5dCRvoAyM1QpxsjtJZzf
oJ0f1yljpTwS4IZOYZ7aUK12uSKOqVx5+K80uUO0n/7qM8ug5GixmlFqXtIbcUgy
8CYfRAJn8+StEzKCXgJT5UL9rQT+Iu/z99DpxedjNz+/UX1WfBesdj2/r0e5iyJr
cG5WBIDDgBL6N93iRsVEWDaokIzx265nKMQqwQoQ6IKQ6hqztCfEFAZV3bTeHKVZ
qy2KpCYWijDc4wLnrdvLPrZQt79Ps40t52tHlwjA5zxjO8WIv8SOYUOp9T6QSgv1
hBQFpFEKjRw8XkMaAqU0s4ayk+YyOQvRVywuVbZkvT8Vit6f2lqooLxhC5w7X0Bi
L4nyBQ2dzSoWf0iWNE4hPCiTb/qAOQIoJKKUGcWDM7AIHYB2cNzUvGalrCDi3vrb
IBl35l7zwnUhWmGic9GDThGJ/IGIAMsIFO/S3JiMFKLlFbAh48PCeh1bw95YGbC/
6Hl0rAENMhfmvEYQtWTUu+eOf37i95V7N7N0PMT2W9yN/dMVTQooOwKRFizrVzNJ
rXN/6QHp+nxUJWXfFqMmTgqsh9ymkIvJbvVZo32wDxFORsMtTmrWiN65Bh0HxfS2
wWpQh7pf5kVMCjRFes+gHoh5rbr3lvuROmolpxkY94lXbcEc25eXQXWsKGAlmDhw
tjj9dsVW6FYzMOOX54qXf9ozJov7KyiUJkqn8bpoWLTRxYz1KQ+4W+eH7GgfzvXW
zLNZg85xmqraETRUzeci8QcvAVNlU/qOHuwT/Jirk6cDagYnReVtRHmCH8UBp9Gc
4vf+1eHeaR4UtyG8dx8os0NG/p+5in7yRPPQCUcKkz8RzwwdapjGoQa2e6XikgJR
0atZ8Q9OjBos6BRLp59n5wWmfH4aMNZKuB/czT4su5gdmFELeZaZYjYNFC/CxlTE
HWS5Ii2f/JX5X1ftLjBUC5ndmwob26zf2y4QyjFj50vssxGeYQhds8e2udp916Zd
opkWRGrKf/4yLCVptxcDS5TNqq19FsG10ezx4F7Jxmb2o9HTJAJ7tfHx5o95dlue
uVk8zaUiFAbQhVFceKTdksbVy3DfIp1gbRkWvl7Q6rEzGLxHSOkCr1Nm8BsqVtUL
wt0Pxoh/UU4+tzN6CKxZ8kNSAXHMI7SMbMrV2SF8MTgEsfnUCUxRSwlLY6a+AWci
L4OtKJQZoA6NCYrHuIjxjmliq7foDv1XNHECwfv64aRPDURyIr0bQo4L7P12u2av
9wN276RBSQJLpgykjG1jcSzhbIMpAi93uZkYphXHZTpvpNhguu132CBGguFSabaU
9aRFu58QDXRgKQjixycgHQuay9NjFtpe6DNMRqBVCVE416cxwXFPuBacdrA/RATj
k0vdUYrgFfCxetql4Wjs1H6rULcQTMxRQD4c579B9UAXzqDOQym9Yyax3TKwAcBc
FFHvRJRp1j7xrLs6F70k5DEVRiLzVJ12VfzLCgJiUDdnMxmtNRGs7sUkCFmVVLCA
3/0fm+Ct//03VDB8GASPoiIAoGCwRthXV5qa29Izi9Ri6VazgrcfqqEVtnSMeyWG
6xFN8jAjZNvHfIp8mi11v5oo/oHx6o53BaUfG558i19iB/l8ffCe0wWGxIBYAypw
8v9sYGI/XSimMdd983hBGqZWaSXAuJ6MdbVO04HjdvJo9BkQ98HGkVGoOigEJy5s
k5ShFX1HlekxQr3n9vMN9atEHoJtuEfJMLStTL5iPQMnctOPP48Mj6FYaaB99OEc
uRytuij8LMNhosJrvzd/n/g62hL0aGVYxTflioJqzSbS1eKjP11Mbdgk6nkwkLvd
QUK6tfYv7bgGC4aETQIKwsoRkmxqPCxTpLZLkid6AoJJDeN1c3ZKusINBffYQHlk
zkVgz3SAXXUobTV1I1inQNUBUP8MNngNsYexFLMUC+nAIMpsWG2nOr61JVIBFJUz
uo6op2+1RFxPfD4JWUMetuITiGMWf4JXg5BfFHWTYtTXKEUIHpYpt2mXlelGej7j
whqy0lQbMKiN77Mvwwiisuhesg436TrvIoDBAD8FREN1YHDv8lWtu/VHvvm/eJpc
YjhdBnwcCANfLxl5tIGK9ZKP3aP+/cDitQjjX+pD4eqSD6Y/91wyBVvr+RDGYmyk
+jSVmiXfzAYaTjh+ir/5ziSM/OCm8VzUySGWREL5wFo4LEkUctqL8kwJUj7ijAn1
yzBJ7QMd13bDO/G9wWYuQOERbnhQQ+9k4Yq7hfUZPlLKaAaE8nf2ad1w9gqqFdsU
WuZwAJBIkPvt8XVfV5c6NOnDXqigxAsUM49FWTPRSLHWXnX7zoZCk6zWfb1wi8oC
07a3penbx4+6aGY01EmxApVsPOhZch17h9CIfpc50mnKmaPzE4an2fEXcI8sFCbM
8Mr4lMOiI3ROUZSFW0HDEyCNaczoaCFy2kU9s+EaMqh7c/3auHTjwUgHh53HHEr1
jCuvlVMgvPGsc2qJYKghzdI22+F8sHI7Mzppkckgni11kMCnh5PQ5tjaGbzzKBwA
98Yr2pbPHtI/UDWxo4KbKPtPapF5lumfg8hxQ+rq52GH4+1GPaFDliC7aajaS14E
6WIlnaCHGRxVioPJZ8PeMt2AUIAsaKRGO4z+S1zQxavwiW7H0PwNir1n/FXchOCy
RK2V2E0Z6p1d+X4cncWyyZzwcVf78JWYYjAAZLll1EkYGeMhCS9vrGN4eWnOVFCN
fqD4yvT9YrWzCVEbcMgLc7t68mQIFPFBRMybq0yCCQ7n6q/VcWnVvABoVFZdH4aj
vzSB9sBc75uQgaL8wAwe6ZRB8dGg8qUTrEPOBoANnVh9j7kZ4jKVvTfQslC4Vn+c
I7Lm+D+ZNXKYiOZrXvaMxic6HU3EDJ4xzqn5hDeeR9BtsodEsisQTwXInlW9Tya2
GSmdiS5GLrHSUHVNduZVEg8FgmYIdCIk41+Eh2joTkl6IuOgGzUlX+4HiHDcty87
BK5gvzhQD7DUpnZ5l00YBCCdTIF5iIENB2CSvHfZU38s/SCb1cEBlcA02sAy8ZrZ
hMEsgDw2btYZBH2VqSvVxG1dNe/jUVSMj0w+78fpOsD8DMzxfeo/iKAkcExjNKPf
+TwIdUiFCwKpiPmueHJY+89NnkK7UW1Bb1LDRZ0L9v7OIezxMipWYIdVoQsJaNa3
ZPwXdct4hEhZCQPGByBNteMAgnNVYMBGBL88iC6PqmCangg+aIQ8NEbyt8hKVIcr
oAb5KLiJ4AxRUGoDASBmS3bKQlFByFK5ra8H03+EU7/5f07CCHKRqvlWLiWv04ZD
OjhRPTR9kp94PjwCQNhfbiRdy/P6DrvKoW4CD0wQHQSs/IuBQisjylbix9sJbvqC
b8mC1paF6TGk9GX8ywR9d44G20PbIlfjX2oqItoS9dYwvskjgi3v+HN4dU16kKma
0idI4hBWRHz5Txi/jDsZEVFir2mRO2PoYVuhf2nMBEQ0RerfEhte2uuXKpmdD3Zg
SKEaeuY8FpSz5tkqxNMvmjjsksEdmeVQBuhBztnbDFCqO/T3rB89uNV8X3qwzS+d
r5GWICeO0fYioi3YEQzY7AkSjWgR6XKVkAdZRwNDnJZIwWlzCajrbp3Cgzowe8uR
13qE1Z6FHD+uQCL4SEy638p58h3oYXmhYwvNnUNOYbfmdOiE2txFcTHZZoRpJuOs
QYJAKFIeWf+Kn2n1YG1HduTo1rHY24YMt1WLQ2q5aUoG8RYnNrbi6nhBxIwIBWi0
DyqOYWiEzP4oXoH2P9KiO4MGwwYHflvLs3BlYaFh3lKeF0AKPShFaEYVeoeua+j9
NINFg5a0aLmGzuNMN0RipNVfW1sWZLGa1NMmV8m0nPAzMol5qoX4cOqdxDSFfKTq
z+jEQUtpQFU+pdgsqHRr2MGBcBpOwi48n4CRH0GlGCukbzZcKXTge4GVuWZih7KI
3zyZcuf+mJ3pOWAmlVwN5eUc17qPHjuK5lmffT4RunduYCB6FMVVg5sTyPpkOkOP
B4oCWwh2um0Oj6N0uPovyQPusgt5NQFILSmnHP7uDctkXCEqQNsLNbvJKGXBBfOW
dLh2iuMnYBKQ5NI2vZeDpDdnhrKT3qtcy16XSM9CwWwIv8UzS0qESKRkybQMbYcs
dU67TBs1Sr/YPbrSdGXGUiyUD2WyaIUJ3G+++onMwovgQioQgujw4G4nxeiF7t0u
mrfb8tWiGVZHwNZ9Kmi8N66WfAI3Dl1ONSp5c1sPuZYI7viuGpf3+xnHsq4yhSGg
PRdgw4mUOST9dKz5rW5a7d7UAnl9klHizHa+1bCnu3lBzKdIr17TS9txK4dqqOlj
TLNbjhNgtTkxKSbvI01Z0pp8Jj9agw40MuHwGfYZQHtdyTbnDciPiSwa8rjzDOMq
o6sqV7s5iinIzQuAUi5k76EFDFzmZyOQYsAdHarr1p7ljudz6x4jMmdDSHYPoA9m
KxODHifuajQ8faXdB6Q+euvXTfG3Mbebjv28xGu4rJ+axFNrLjRD6HR5PhMCewMN
CaxXP64/i21taxuu5BjqpmCpXnXceOcsHqa8GFK8UJKTX2kDmZXdajyufdAe7C//
NzB+sI60ryV1hxzCJz+OIx+BBmFBdU6300BFLVhXkaO+Pozn44d+DZUHH0EFn5uJ
pVZ1uH+zUmCLM6S6m8sAoKwUgp6orKi6BoMD53BB3WgDwfYmpL+4ABJ94KyRg9XE
FSG8SvEKEE2p7/aGw4OBjvQuFHRMILC/0DNk03e+zrXypWriJyTcWUf1940DSMod
FIcCl6JGe3aVWv1K8pis7kEPMuWl3Obbyc/K9mKgwkUjqB/T7X+cf81oCQwunhay
m4leqwiw4jUqOYDHiUzjCjyND8Ljok4PyIcPNzqtT3s/IyOqP2adnt/8bafPXkG9
gaxmuna1BQuLmo3ieDvjTEtfcD6N0mDzUB1/VNxN+eDBX+LMrDmZqcLBZ5DJKhDF
CteeHj/C9RlvrTXORI6rvYPa2dRkJBkyx7d8PyTYVmLWBDQRMt7oc+/qqqUe5Ahk
MMSkcYDQvd8VfZona/IKCGij/abCzY+cEFEvW3ei7ucPNEEeOe3BkG43MhxZXrS/
UOfg0EX+1+30etQSGiO4eyOM1WQklsSUAEh+uB0ttDeibSmyAGlsnoXGrPQmeAFI
4oJVIta6gGG/ohJalkfepIiGGWvFjZUjDe8YUADf7yeqF7MdOH0i8KuZ5aBAmq2g
HqlBhAGIX97Tn6HRGlHfUAHhHl4p0CCti5u0XNO0PfrJfmcal6r9ofpaGZFT2P0A
q3J7ID8mxj6mp+ZZ/rUU9x5ixggwVks9LslmnQMyndqW3UtqwnqtWeeYlBawnvCY
g8NyGTIv9kaZmJG+pIPY/rV9Mp87YK0b3X7ghbAJIUCeprv2unM5/lFVRZ4VreV3
/Whq5v0p+epV4n5v6AImk9hJWFlDbWYgv6qDu6fFFIeK46qAq1pmc3QvZHc/EzoW
UTGw31JaF6ikIEMX1rtKAS8e0OmGOySxCvnOAHSQ5364YmOYkwunNS6VmOeitBgP
r7ilv8JU/monOygXh+GpMUA4On48psMDdzj/7XwRJpua9r4hU+qqN+i2UGtsMxGt
ALLQgA0FkMIfiRbjqKC+VH6w7KR3oLSR76nt4I3ax9ESobzkzU/Hyq5yUPNYOt+M
8pSzzpXB61D0T38G6y43yeo5wnQ5/j7FyQySz42Ch2Z9hpMYlFmGj9SHlamGx1c2
vZTN9/BiTA7XSHAmEi0YG2wP2Yh2G/nJMgcBRm6uSvkgU0OjvCYJcOZQ8xLZxw4W
ftBCe6AZ5lZG6m9QzvGyT7nMaqtUeXFCQn7fqpSY0Vk33yiRxfyeYbYvCKoznmsB
RSKtFYd8JH6uLvGyjXGC72FswH0ZhaI7mxajVFfKN+1C1mosUWPb3/HYmn1FjISs
j395Bl95xJZ22V2x786UYLr/X8UCtY0E7a4xEE2wzkmULyQBn9M7VOb3n/193Xxf
/3YMmOGsqYiCQt0/vU6UGPJu3zVhMpRphNm28YdsW2BN9iPkEVAWnPi3OfspIes+
97qzG3g/1e1CqS1VWpzHyJQHFtRMJr0kyBLOp4u549LOhqrIoCNTwQHBHIlRXoVz
PVvEFol6PflCzgevlyv+D6erSfW+AIHYS0b6CZT/SoqxgtY15QqXmxH7w7yhq+4p
kvxVDQjSxZS+nOuf9G7T268HJN7S5HERH/0e6REqmTCsTL89uyc0VJx/5FH9D4CG
wc3C5OvfwZMQBU6Xm0evyUOH0Hn4SJ+7PSUB2Wu6qOiy3fMjM2xONaP/ZpyMJRdu
25K5sikdhBVGPXUICNb0OyWTiMiTX8GZ62LYRcgRVyvr7cxkRFjFznhFaH86c5Si
DMMN8yxKS4gORoDYbSOi5b79OXDqHCYTDCGzHeHspR5ENjclhjl6gaRRu7NvbKlh
fbp1F//AH4IEfzxYLEI/QGS2km+E37CKnzPwdC69STnMxrN+SYKjyz+rxHr3I1Rf
/l6M9JvkXKTzjE7JNRgVU7be0rkuksps7fAPHRqWxA05wYvOqCQ49xp0Y2EFptkP
ywkTafRapRsY5V54d/2vpTf6HcEFoy/a15ax/wScWmmSMklbxTQulfqnQXTCOGBG
ToHk6fs5+Ok4pCBEis3kR2hk8nZAT3b+OcEoyJDyRNrJCQJz6aj0zinMoKSu0sbT
J+vE8I/Y7PEaZCkxB6xVXhVP6hXxtQ6woqYbi+0/B08w/Nz9182S/bcC5YeRyPQd
O2FFooQeeNSgtaPw1cA/7pKNxkTrSaQXpnLNRP+ZSuXkhKu/5dvetQWWLXBlcXSY
GaAxPkmEEauYOww6LyIPxoM+BpVIqESjtdtavwlyjArhcgE4DGO8SkxWY87M0jwM
PSfUWc3otYWe/cb4RbdjAYu8ms1y7F5ky01cR9hgRjqmAvCua7FVhIA8GXPIHyrf
fProJEi9X/ObdTPvt6l80mVRcjpcatbXZHPIZeTcYJMejRSx7ikXBuwtFXlelHnY
ZsJGA6Z8rE75T8YPVBIyUq9QNXi9xU65fqPGPKo7wt8CcluxF8YKIGgOE+GqJC7W
txzGmx2LFYQ97r3gMziWwpRMXR7P6XsRNdG9CG+LBg+as/k9Z+BnS/ZGXshPFBy6
lBgJBLT0DEMV3zxfFZNgYAcXxV7MJXenF091ZUcBziTAMHDQ+iXCkIXoFibVuVIi
uDFZJTfPdSG4FFb8d6l1mhqwI06fBYMqEc7nTdFRUizzvOzDF5kotBtQ50zcM//Z
Sam5ydXjF7YVxJa6Q7xdmj8HyQMK2KgQRMNBpl5cQcB5UA4YvhVZK8TbocK1Nd/Y
c/5Bz0u2jaGYsy+NgEKS3P70lksDrEAQWf3gxF3HmF4++u7crmKKhFtvmRpzyWNd
pj82F6xO79MO8Ds42vig2mQLsUh3TMvSXK6NFUEFzstiPGKvG3HmW9w0Umw8F+oR
Oz9JBPSJjcj+fPrEO4icFbuqljEfJynZZGBdwD8M5mvM56c/MuwDf17xaOrg4XLq
2Rf6P7PgKhk8aSLSnvn7qRAGwSTs37lgNm8/bE0DcKPe5BP6y+CWJ2dB/ZkRJO6a
0EVnSq5HWXtX82ryayN4IjvgM0nxSaK61sbGiCkKu+WZdi5okuURwAtgQ8By8dqQ
AQpDlDYM+qL/D8OBJ4Y3tRtYiS5AcFvhaogZhkC6syT58y69tLPYsIgIfAdPY2Po
/5s1T6nU9WJuXbcG2xp/21ue9EearHh+UqrXc1pVG6YRENjkkI9WYDLOUUfiQjqY
fNyNsLRFOEmg42eYtTHPWhzvxZqvRPlxEcr4SuxESAIfEi+DfD2TQ6EnOeAxDFZV
sDFGD8N9xqi44E77ediNR2pBxB2FFM6FOUpc6+QKLD1fvaQAuT8gsnNq1s/S9Jz/
csV5iOTcdtPe4icEFbrXNprxKu7h05cYc3dpbCqGrzigE1hoH0jw0PoaemWP1Fs2
flxkTSrKnBt2zZVOmXBsuwcRMCXD/jnuI8dawp583kPqI8y7vOMEQfzrYiXQ3M6V
OL0YlN4RK7a0+ko//+xNDuxNPRM/jCp38RFNS/b9EZRH843F28Z/s8zUADr/gYQi
/hAol6MLa7o9+cxCDaJn00aL+ufBgiFwuDriin5PHN1Wew17aQRLJL5FvNBQ00K+
dQYt71gXLh94hNDfuDLemp3vQdLwARjqE+HCvlfhwgaJFaIoh7IAwv6Ue9aL3gYW
LYEQTJFoWkpX6joXo7PMhGGZe15GVmHHkTP1euMxFSRjPN0j44pRm794bfUTsbfx
QhXvTlENaR5aKb+xR8rDL6og606+BpKniorqQLVQb75gCcIA+tzhs1tvUrHGN1io
+A+DP0bsGHbM2VMYYJn23PiS42RSpCgZVXnFN6d5QxvQkrsPwBIk2F9+agJeruXg
+MgDX/izTda2amZy6MuIr7k+6djWteAdY1ppQPwnJIdw0osB7jrPfiALGwRnnHT/
36/uWCXFq2avu4L6smwb85/fWUfjwik/13fJBUEEGHJTqLXPU+d85QA51MiPuncS
H69+gH32X/7ssfohsjKXmAh+E9RKBcp9kNbgCSLw25x+P68Nk8MYUmaaAa9nBt7X
wAfzXc3tFeL46kBIDY1HW+HTK4EI9Kbexhfz6vh2so7sKeznPJ2kmOMdPvcDrPXw
+KUaYcXFn7nYiKK7/6l1OuMrcj13SW7XVTi/sGOUqSiAlOC3oo7Cw8gh8Ev9cduC
yhn9fjpBLdHh492PCOL5xA4QMcaMgcuSSrjdHqFXIILUdmFXjbo8iU6Ej0cqD4xO
G5UqXuZS3cL/Sgjkzm9LRLgsyV7KInHIhBbJbLKTDrIjw4J2MuaFaOslktj6Lg30
8TmmaJQ8f7tyriiyJXaOPY2AaRU0a3ee1w1vH46xsXBk7ju90VSQo08TMGejsXqp
xFbEJaEYrXKcgQ8BKoEZyrhCauYVUkPhzDG1LxZFltjSZr46FucyLEOq/xZKAHEp
zHf36NV+XllcaMNXMHBaIpFeqMob8FjSIGfIeJTweQ9YIw9Q3Tp7IslrBhfx00kK
JlrNlQZsP71D+aRhML3PQTYW/muDJLUdjBtlAHNrvhvR8ll9PxDnkyq46Km0NrKY
kYOGC0FlPES/S6w4W8GbHWaOGVcZ4XjUvMBWZVku7hkwmgDHfBwTL0/LPHseMW1s
wh1Px1MapYmS1ePaZdfqJJjFci6ibzLE6Zvua6w2pKkifJ4pMXv3RyKBd0m6mpU0
D+V4M0srdWtMw/cgtSRtSEAcaUMnT0B2DNjcHsd7wdeRZ6U+y08yTvSy83c5m/C9
If25ciPWyj0p2cvVe5eeb/1spcE/4/hijwNPr+7jUPnn/D4AOnq0/h8NYcV5J3VI
mLv7wl03uqylSfIsDEMVBRbUv0OA1unJ25K51oKh6m9hZkU0LwvzsjsvhOX7bnOw
qtbQEvCehVN2tEwW4/ATG9d6807GxmFWkXgHVL2pEqE6fJaL655v8N5Nrzjs4mfj
zvrS2BbPs6uCLwOSzDC4IK46oP1ih9u6VRPFLPw/I8IDz3kkV/ML1spIOhN0VDJR
A3I+UxgJH3bs5hQ1KfVmLHxQ5oVDfscVa5zQs11slInG8RVvkbp1Qdx7X4rHccYE
OmpK+DAH70vQQVejt5Y5ohiA5vPCjIriXeWlHtINbMDMc6+Xuj9nMovdNyc7MjSc
BccAdtqcvbT5zKT7uTq0GpnNyXNNDazyNIugCBMX5m345zn7o8MADEw0ClOTXeXx
O3qok8u7jn71ZOxD6oGKzMEMRmcuykJ594UYq8pbOKkRdiRIM8zEljDcqNUHD2H+
TJpQghz4WdGiEfRrAPXPfS8LLKeQ/2XNCBKZMhDIYaIMV8DHuichm0bL2r8hRSlB
e+zZZfsNjZpVyJCU3Nb1YeTQ4021u3FPpc/HUro+MFoBjqiziz/KT+W/5J7QQCKm
/ZH+HYuk5ZgldyaJoDZUUbjCj4Y3h2tBkw0ADn3BdDS2aLgHnn/spZ8g64Z7U7ES
wecpQDA2GXueFkkwOwzX2SAXrYPgI2K/tQLRCtOksgebO8hIjEr0r9xRX5O0hC6d
qqv3zwiVWd0ZwSL0Mqfwjq2+iSh/tiR9s6ESC3K9wxBnKQO+TLYD8WtxZmnqRsow
eV4mzbdakwgmZOxvh++Uvga3Q2tZoI3Lj9GJ3U9vD9rC9aqEUvSljr5abRMlOSXt
/A6W0lAd3vRGBVE5r6I7WvyJ3Cnjp7jfgTQNfXee8IRdQt9MxsXvpY/CGrm1mn5D
MuV+cp5mYJvPWA0HwOZG5QTkall8dmARlnntWJw3gMsipfU2Mf8qLA96FsBwTtwI
T8gPiI5fyO+Pe30uAiyV1oKVy9WnSCEGdJjrDoJnYldNu49StB/Td+YENpWZ1i3b
tLDtHSvkPNw1Gxo95Oow7h3FH78Y0633KZYuy3kPcQt8UQS7n+L+jsoieSChAtT+
aAHDn7sQfEg59zc8PPC+oR3x7syPLI3fYuwfwqyU676wBxPWUJCRb5mIgIK3koaU
qrg5OnC6tenceNfB85H593/wzZ3UvVAigOXykvWKsNxiQ22dMo8YjEIydSAb0RvW
mIRZhCUS3v+ojmpevGxOXLtxuwMah86/6Jw5rlWw3sBaX8f9Wb5IopdEXdHc/ZIx
mzZ/xVuUsFH5ryxlJM3Dx3oxCRGKFP46fydC94Iiwa9jrZuYG7WpDu7UYYqRkMM/
ZltxKT0Lu/iXktdMq86AKzz8A93fqml+huq9E9JGgwURib1Pj+h6miZJJo+cejsY
fOT0iItvDwqkb7ZhNivuGIEuIKxFYVFt+rWgnPn/MNv7Zq8H0M7+tnBn2oGUjEFq
mRMkm2lCNDJ6TzLtmMQnx4+8tbbFSZPzAlKFY4yz+OtJc4PEjHu9MpZQhW7FTSLV
SC3O1VuvRhQ5A1agp8ixy4rc7YlJLou1U/lzSDFDvRA18T7J/b2yCmMng1NZ/mAm
Cf1gT5oK9JtkkwnI8iRhVCjtfgvYFkVbqLCGOpG/psYD0lnvh8vGqeeg8iWuCY5J
DF8RPChqCYdZsfRZRJuDNu8e8cw6gdyMUKn3tIK4MY5D4sXPXpXSAL2BEsw14UT2
EHfzAFCa4fEZMm087mFRAmbZ8sdOwwUi5qJ4GHjo7ysL0V8tCVfghKQmbiTNvgWn
vUX9poaHUCyqzw2t7YcMmAEcpWgU6qMjcEcrcTfXxRWOTfosWB0kppZeXA4H8yLX
189U92VgG1UXJrmg7uob35vF3gNwWkoVjdNMIIIUjM8TxMy7KpzlQN0mTTyNNvnc
oDAW1wHiRcqBtA9f4IA0Ab/kknMWiowZQcfaOymU2JMqpbcmdREeAEo6y9nK+kVm
d/+TSu8zNRW2MRJ6QfSvLYvQUua4pQJvQBeYv4yCaXxsUFeI4W+udasyidgZniep
Aw0m3PfnjReRSO47IWD/IJ3VZEwlvC78piMCETG6MrVetilm8XOne4WJu19N57m+
tpVxytgo0uO4I0VVxYkMC6GKOb1cXaKxvqDPpB9lPo6DkhtL+xruvQqr2m7ihVdc
6w/4bxS0XSrYWr1ZysRr4s8f2lmD1/g8xLxuk3iJtxLb8Ih006PjqZoOlo5edTBb
91RrMOt8Hvpc092WZwFVHfo2IfAxxbiVB/k48p0X8tCFSAyqDuH9dqUZKbhtAsYC
bCmP6MuMmpBzEHPSNOvjXVhmKlH3zw2IxVTpxPyGmcxvZX4psTi0EMu5W5GWJuqk
gZZmqrPubYee23A2rQ4uGIt+/mhoHF5+SkEguqUcM0s6DlgApZE3zwzFv6mfO1C8
h9MrPnszOx0cOyIujOmE4bNN+eKeznf66KG3Zbhahm3bm7MWDjoE6YDCMqaDQdxk
cIQI9jz5d47QAYQRg95wIbF2uHLsvGreBa+5UeKMbkUawwN5DcuIp1GrcHmP75kG
Nx9Y2xLJuNn2zOAB8sIjCtHHPv/5W01GhYYJFNMd7MedvAxHkQXdV4p9xzmV2pU+
W9VBdI0QcJstaRMXtJWWGrGZCdiLTp1nkMwfsd92sAkFUG583TsmPB5ymuSbch9R
sdJKX8uh2tAeFvPNvrjNNh36DawrBzcM9DU1qAVpQ6C+x7JRJcQoC51MKRXL1wd/
FupuyBr4e1SEStwkcxeAsmn8u6XYg68kHGnOOj3NWTGERLoN0S3im0w6Dz5ZUKE3
DH61XP1cje0Tf4kqIJF5KVvn4xPi/IAsgVmVC/rxDCvIbgROVtZsHNobXcJG7QMj
tUahWCgHM/XKzKy0wKib+ayLpJ7cfB0Y+MYoOA1dLvV69/QhFx6KiktfBSV6UvXd
boYYFCgmmjPx8haBPj4OiWWFnRXn0JVfj1dY3tm7G40OBELyKHm+O2ZNzFMzk9ID
sEgKAvjU1zeN6FIBD8wUFhbY0ctm201gK0R1ldovZS07SO7DhvmE4pYEgw0FCNhw
ywaqtc1cNYF/Una3xbGWNYqdzijVvYHepZnmR0H+XRCyeyd8sLr+lrpTCJuLgNvq
ZG73DwfLwECa8a2nfBPhrb5EyVZSC384vZdjlPy9dPh92rWu2CDQToXeayc8Grkq
qbAtbwgbeW/zy4RUDUPjryTjRFdHw8Z21iE9pkVJCa7s0VodR/YMEdokscbhNUZx
gvjNqAueLi4/aZjdScP3yC+U7oScn8iqthweWm6ZvSHCHLIJK6UO6ncW3tGv4HDK
9OJ8MWqaBNc0+NyBHzCuQqZgxoL9eLsqE1eVNBmvTqbsj4MScmrsDipPEYnbVKM6
MSmwOTLLXrtN+YmmkAt75pKcZQ+SQbnDSa9oWf3IDsnBowqHfUIPTInc2S2nPKjK
qt8HxunrzPzcAamM68zOlJTYSN3Y5/97k0aKgSktgTVQFiGZPLaMqZoyWuhRmywF
TYzLEdMKQZflcgi45eQWBJm7bjGbrJbGBeObIP+Yf/GsRca7ySkPEZ5cSTw0UEEp
cWMysy1QJcLbp20SibDsUFqklqfZT/KIpz1vA9Bn0RcCRd6HmmwtcgWE8kE6VMml
UTDxgxQvr0fB1RtXDSwTzKp2YOlnSkpuZEd2oCdkbtWBBt9ISk44fexIBhRhliRQ
TBNDzUeUhIbm+vbfbSA8qsjQyFUgK264SvZKCSDw3Kqw2y/DD7+Hjao3NgcaO6JA
f/ssYeDJlzZvznXrFxqBhqMVgRTAeFrfzrlsWrxaBbpCNAy0XQajudsou/I3BrXu
LV/4B4qTs0TJqMuRB1ckjUg/wErPun6jXRh3ATplBg9k6ByMZl58G6POrUegl2Ic
ByE0nFo4RjklecSydb9rPfnV7hsz9ulTIsxa0HNVkD0s6PD2VbCh1nYkfVFWlySj
xw4fTmaPNw1qEOlokXmcNO/aP/3fzBtjURPfpG52v32fDNrWCZYmK1FXmjZhkcte
jnHW3JNP4lJW9rWLDcVlhjfZCKLZAFDHf3yBPvoPPfU0TZiqpeyCtveHMbTh95+U
BXRhj3ATqF3JC5BZcayf/3IR6kwsJKmuZLdXDkQfdt6V9FPrhy98B6/C488wP30E
a6nQZ5HAr7K532tsVB8DpwDZKSp2ECUqZiSTCN7da3nRWmNUfUWqlUr2sjFRIziQ
Bb0viN4/81zJ+Nd4KRbjduWmlu8AWzzaLYfH3goS5jlLqF8LDdtirNJOEhkKYM+2
d2XaL+UybIX/49Obta29HeW9J/ttAzKzof5AMfg/r7yQLvt0MoovDmrJ8MOfvS9O
ALQJ79wTLflJX+9YMrFhUowCmYhQ7UbwWdty7z9OQuD+QQVpjfCPnoMFCbC8vWg7
qrDLsk+DiglcQdWDAJRNrqe2koEywBqTYXdJvbZXh5jQkQRpV6ZCjU9iRSsu1Fhy
jQBhODUMEbZB0W5BxCRPTR/bgek+eiIvews1Mt5EfMQWoO8PVVHZPzHyhqVrcJx6
303iw7KiwMcaYV8Q3dEJIvbZ6O/sJJlnWOa8AC4wwMzJltARRc8DZDV02TNClpX2
Z3h0AxuOYRUiC2pEUNv3Q1VQ9N2M8ROOOj1yG8IavAUMiiUDOtRa15yjP50RCp6c
ZRwOk1gn3lY4zxII2Mtx/gcrPJomR64oMk9R0ji/ob0GowytJtiV++C8PFlbW2sB
YoqGjQHrFgPJXU0sRlgmU1m2cgwXrYDiyNu5VkK2wnHgBb1n7n5JPcf3TNrbjzau
Zo+egH9PvYzrUu83dw4/hFhPCtGCcYbTRY7ujQIe8CUoJ/QsmgV7bWf9qZ2s2Aac
L7itd2y0fDlpINS7eEmNdNqRm6dBUvvOXpw9BVy/5g8gQQ6I63dwhPjis/GLLMCI
prIL4x4QBHPkj+vmthzpyIhRUxHhK90AIs35rvPb6GCHAwosck/rhAw8O8TFy7HS
HssIW9oE5mu6ZglhhBlitOOpUCfcftD0MStBPFSHZQMC7NhAB1FEx1wsciHo/xDR
POMKea35yhn8nM8AFJ0rh4Y5l2SC46fLDqp3M7X0gZLkx0MP3hYUF7UA3AYgd1He
TlUXVPflnt0drsCEMBwk9v7izuU39PEyI01muzmXp7cVfI5NGO8OJYkoJ4FLsIqR
LI3O+WPIlvwQTboVoIHBuILm0UNADOlwfTf75kLvLp2yu8aRxOqJTMzSZ7ckCRxH
bmJuzuqdQFxM6FLMhIBU70eTk2nNdz3a0R395i8usNYLVRNaViPpoYbHHlkWb0Lh
x2GtfSTQQ6ggVRChkDURLXnqjTrcPOfTWVqxAFoGKZxtdfpOQr+G4d1BMICFBoPY
gqCTvz776P6M5fp8/rVME5/tvKJqeskHW9hw6390DRoGNWQ0+gXBfC4jiSe2jtPk
bwItysOY9UvJcpIzgVwiQhRhrqaKow2wufSi4UfXzkQkxtU/IFXF71yEE3tHNqGW
WddTF7EozIsANeoYpwJet0iO8AQRGbi41Sc5WSiVCl6yFWqqvMrtBQctieKX0skY
QssRrO/rNemXlNk3JQb1zW0AXV7SonwF5ANIOBvlQsvlsHwMEY9ufK9twt6q5ftZ
gFJi1KcrP9m3kGjs4HHbEIyU7eMBa4MDZS58J+2OWCNAf2KKA8jVAwxsTHIOHcWw
xVLC152kSJRH3ZeD3Nha7g==
`protect END_PROTECTED
