`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0N7WZ/ia+Os/h8xAc/o/Br2BcNySvjiqHm6XnYTTp7ypT7jdNPxIJhka6N84qzgV
+Ewe8EmxZOUqoiqrNyD/tZ1qbuiZ1Cs/c8B685oJQ8u/W2RNYzEoitx0EFzvVKXv
q2T1fYT8iaxkwkRTk846thyIwCZY+TQCApkdcbuTvQrdQJMfltzqnlveMGrQ1Ki/
+M9PPkHsnje+i9CMK+4vhnPukLwLOkNeRFxnc0TTxVURA3p4j/wcD0XyAqGINm0M
i+3R7qHeRBWl30kRiVRjWx5Oka25Lk1q/oHH0J45SjJEvsAAfI3mnQgb4zp6S8J8
2/y8hxsN7Yr6Q8UBLi/uoHlvUe0Kw3udVQUXXAzUiRxSPFjhJIf63qChfjCObiX5
97clIVBzMIp7hvyidNKKz1pShovGCC9leC9gem03mR179/zFg5XVPvm5PXJCMzaW
2rLdddPgI50pENtmKLw6nEFzsEV4WIL5Cr4p73KH//uUs7+CqWv9uSoHQXI9ANWG
t8svkEoUpibE1GcfrndNspw0tg2qJD9uKIoxTBs2jZVwTCSxEDIH+uggi9SCk4KW
978K7VcxzSJd5MJ9fQVT/N8fOWJEBXrbw71KW7MNnwzDvs5J1kA294bIWUUAANXa
stxbxoN2DaZN+SU9tNZGLN5/KMgs0zJv6rLwTIayLjo=
`protect END_PROTECTED
