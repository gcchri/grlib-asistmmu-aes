`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C1riJmeQ5lJV/9ejmyM+FazHKhUPJm7aYSWFu1sNKThx7m+Oc+JV/O/5ufSD3vyQ
UtfUR2zagh4x39qVykbxu1OvZhlgD6LNX45GO4VV0yp38Yo/cTh9G3RFO8fsAD2o
c8/8BPGt7MH3xM1v3xC45S38xVoyki2CX5dw1BNz117MvnLkC5hQ4H0uGEMmEvMJ
HKXCFVZMZhyE653wh6Unz5pUqfkXrXuIYW0eqTzwfqZY2nWUvBbCw8BuDWo+rb0S
6dd2SvOKDsYKiyxFwnIoHHeMsGJzLtgbnPr8jwS65fg5pGCqnRNGk0RivZPvwbuG
X19RyVjw0txs7Ld1qjehk47ngeoE8AskNsznrzLgCSAfuhZAqfFaYgan0P5kuDOl
9EhDN8JVB6HchplXEWozufurxKu5ar+oa389zgLvDggFRUaaSKYs9Aup6ilm/8c5
Jdo8mL6L/NV6xuDlnaHysIXIc5uRGnuFBgRNCcei8ZSZApOBlzSu14zNqeXH4NBq
bi1oAr+7ufoJoaSyzVL8+m7Z3R1pNu2aAJ3u/VWfoXjq6OSfN8sHAU2ko1acIP5Q
iBf5J0cWus1nTtIG0k+0/AS1UADgp33lEj/OdHDTGo1K4gAuIRXTzs+23S0+l4rB
FPN8Z4N7mnZoYZNSuM3Dd6caVeeUZM10IR83VNENSAQWWQZ5ahQKOzAZLHUNDoxm
CP3iNg2vdwdGo1sTniiat16C1wQmA9Gfa2cMj9NgqD1dWnbX+iwpLmiHOEfsqqk7
FYO1DEKPXIaWyHwEW9JyRxAfpSlWibJAWM8rcfv3c2qsQzkSyf8Suz+y0mU8GI30
7AlWrCeixDsgP9uyjmSX/42VG2Z/piAkUZOEAjrDyMDItKYMe0vUKzq4RJeLx+I0
zPIyj6i8FkJqO9apZzNGbQ==
`protect END_PROTECTED
