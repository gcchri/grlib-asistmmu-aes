`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8WuqI00XhpJJUZRtjZc2YPxybSiCyVZw3+IYi8nu2Tlbzfwh4qiwUaOztY1xVGGo
OA5pyblsYSTMblmB/UtlVae8IG3cXyQ4IfpMmyVe+Qm8GqaUpcO2MKtE2QRTyZZW
Pmk/DLix54xaIsSD38GI1Yh/Np4zfckxB0aVMCMjZoCh1GA6U8f/poMulMVvhA5m
XZQG2TTfQX8BosUDAfFFDcW/5o6GkdpW6y6JJElRYKB5JNRCmTS52y+z2YIOk/Wg
ng2s3g+/55+kd90/PBtHQdL3TfO5apCms7cXVH+DVgPJUxorVdKdXMu1LCOO23lF
4q79wf9qj+RT+6wyTUNvFA==
`protect END_PROTECTED
