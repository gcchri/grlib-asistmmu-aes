`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uPYeRIeIpbSkdcMnZ46YdYJNaC0h1X9pyRqpywqrOzFschKuZCNxqdXKcVsVcWxs
g5id1Ky1WPlNAgFYje+Ner2o//D4tJ1udjEZ7DAcRDfBE/sBd1Tp4J9FhoigGeV1
D3B8kunR5e2LtmnYJQkz0CEtA2phLeAL5Pk3vjzUTMBbrvXzHX/4sYAs7IzI/fwA
8aReG3/TUfXbfdiCvv3hfkar3UhdlARh08aiCCmg31TVCLR6QGuemk3MBwRAE//o
ym4BVDeTiaC2Bm+rYUPn82j4BY1NsUf0QurY7aFYrHXbGutB01jkVTt1MWea/4RL
8vQq54znbLjRlqrfsT69s9Aw4A/SA4bqFbRzDLC1PUAG4mFxozV0qaVp1rgnFwhl
IG0Sk8+ZhiPcZ9gpPlVtLMI4Pj14z3h/SGsoLQcaoPA=
`protect END_PROTECTED
