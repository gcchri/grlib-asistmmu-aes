`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QHC56Ivp/bHh+JRutiQVQe4XDQczBCVWstCqkZsPTRSf+U5hp2cOGDMBcMvqOx6l
q0ZrS1q0qe/NYmn45n4ew6DYznTh6AnAJM1eOrhtTWXAvAB78rgbE34lCtkMstAH
tJlWfwILB657dUO6aW1KAeZhbOOocCnqu6gVOB3Xb4se25V5t3HbEoIWAKjZakey
13+Xvv8dpCY1L7bkd9IAThQRY2Fhsa/u+dIx7SpWHtScGs7AjmXV9DDXZy+zmtCf
hHIfdd1c4Hcn7CLyn5TaiFQII8tjTTKzHOty85pws8k8VtvGA5Gb8d38XsIOlpMX
hqV4nsbUp3hClX30rbqTHVHrBb3+DTDkBjg9INS8xLOF1aR1EC7fwpJiDt9PcY5c
U8POjDubP6NB5oGNczrQxRX27QsqyhaXCA1CNfl375X69UCdJgFJ7vDUzoQlDxNy
kI76w82bp9jotz0QCKsoW0B61hXDodTH5eaLYDzBXZdGdcXk6UCwaiBdSz00sEF8
`protect END_PROTECTED
