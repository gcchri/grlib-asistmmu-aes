`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qcg2A7vXJzsj7X9I6xrksnui/C4OfS5o91++WBh1s3zvwBFw9JWXo3Fqq7J9uCHh
BnJeIqemRRnKbneQ2FeCUm7f98kT9gmnfG4eOaf1WmdYUL5s1L0mncIoLCV7BrEf
c41qBvcOevnoPV+fZmvSgX141gRNoBHeNnruf/7UKIc5l5U94txesN/h40FYCWQc
k79WiV2MZ/0Bvpl9lATG1TcGrI9fBvPbw2rTaqga5xO79gyBhCTBOCNbpxTRT+0F
b3IzNCeW3VMOXb/45Op3dBTO7mYXtaPJKqogn+6DRVUOJtsCnYAmMjJlLcZLi+VC
fQy+3JQPWIWpzqQpQMhAYoSEVqO10XyXPUWTbh59LlqNQZ2KGmc8YJ4l/37uTmMj
Ghi4X/b0x+I2aqJ5ZfXYiCBMQjKaxj9yc7Xq5+4yrpY6OvKoeNOEK6WTg0OlvN1B
XvP+IBlYGgl4adCRVaANrOZ2xa9+CsqnA6xKTKppgr/sqZNqebGrcFp+UTtwfmbM
9ca7Ki8xf3/FcyGLrIy4CROelmxNkdO/MDZXtoPnBX2qNZE1I/KIzd2ktDORPFaY
tyd90MGGqwGzDlgTfmVn7TGOoq1Xd1P0ESPOMppwV/Q2L85mAXcjdEH7+zjrfUsu
X4ZwTIpJAvEOLUHAIRKiBM8kDHLagMEDOjP3JMQx/A65E7R5wvt+ic/KEcndb584
9/A9PsukDJyDHFBDQWyakAC9/F3cVQQdRrNyzVhKZwVGJ5LliuFJrV9XPaDOujNx
GgiTB0M4Y3XA0tP4npasZ6OSWxO7IsN8+zKre895IaRLTsCcM1amW8LO7+d2seB5
NuRX6EQa+Wxg7N/ZQOEoa8QB/NkFKYB3XCnPfVLGtnFz66jeYe84AvsbKMZK9Byb
0S+K8WZh0JMoKrAeYwYlxa6MRsxH2lnFPfNV2jH+ayB/EuA5mrWyQRjOUBQjFpII
B6sTjKXqoj0qZBW3daHZuA==
`protect END_PROTECTED
