`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KAuFXIm0LkgDkGyuq7qRG/5km2sMFmYcl2SfZQZwF/ySfOxJbDByViXXcjdKnF5S
9AlOitL+AGFAh/pfKQvUowJnRYdjo2/bvmP++S7XzJGzoULVsri6nQYMcZJvrZTb
dbkyybjx7LgAzFqJw3ca/UUlh1My+h9jr329nOeOO7zDrcOEm0r6yaoDRoXBJh4+
7A6XMxiVj2NSpD4aTHVxP9G2rH1zqnwQfrkd/6CLpW0qYIGCy+xHbgjXBAjb5L06
ob67hr7uRhQeden+B/pNRIuHZc8/ED5Grix3KmOCGSC0WG4zY0pbd0SrEMDXGedG
cwt3GRZFQVdwTdgyZSDKVpkuuP0RZBnE4BJEdDfKxkc=
`protect END_PROTECTED
