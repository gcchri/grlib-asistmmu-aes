`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wAUjzBvxtMcLd6qpBjDJBayDjRxLxUSvQXIfi6TUZC6wDEeFXamkrv7JvrYv+Bvi
feWgr28rkVk1vna33WUlFEcmXW/NuVMR7uvkqFuQb8z8c4XSBol1Avf2Cly5o/Vn
zJBdrIYzPr+vxcvQH3nmtzXs6Q+TuNqGa6d4nJMvTV5vmyUrsok6lWU5NdOCsm2O
DwO9+cpKCgtyoTB/9nbhKPqnMPWCcQpLl60Nb1TkkmEl0YZWedQOXkQjjKQWAPQG
V3MaAO86OQRlVAc8XTV1Mpl2mGQYgRitZ/uE+fRh/ymKunGED/U0hhuOQeYdRpvp
WLCuAoUQt5aPn9tFpacJY7l3BF6K2X/gY+kSXU30C2qJCCDMMCrWYY3Lsv1izhTA
PsN0+Oa/8StVClk2QFV2su8PTmwBsf6A3hfQryOAa60EEBb1+0zqjW4lkA4Bugic
`protect END_PROTECTED
