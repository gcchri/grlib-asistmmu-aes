`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KP00pRab+HuaAMw7melvYkBkBHg2SH/6qHE8n0uLVC9ul3gD6P8ON2lPUn701Hr/
h/Rsg+zMbPm9seXPu0/E4DPNYk25NnwtK2Yy6RlmHXhgoWAwna6t8ITIqSP2XaS4
hMifgiS8+vMaWCnA2b5vIEM6ONExmNfw50sOkIPphqF0qhDEIEhhyEqeHBbsejpH
6HyVgxoxTkfGNb+mdy26ZW/DF+3XLPIm/SyTYO8NDc9Ri0G8ShuKwfNS+iXhtJbM
23EqaVfjqOXhnnfNx8YOXXX0OXMR5Tp9Ey601TgppHqiaXkvq1KgThQYj58sDH9I
tSKJzBrLDL7505W5hhamZKrPB6ZrP6GklA94vWfxPARK669kzpHJ6UsPoDNz5ozI
GoluNk8MyVBb8MfaeZjiBFG8iUGubNzWnPxVppgVz7ZAxgLILKGo22Izl6T+JuiN
cyaqSytKwV8QYXYqbyG4BoRhPMPc1A3RpeH7xfITN/pkN2TZ8sX7yL9sr1Czi1Ve
Nij+WWsfE2+5pEttl937/OboxAipuV+liRGyP7iWmZ75DHNnI+/2wYRqaZcCXdyc
fXOl/vOIZXEzNAdGKgZb/xSOHuuZFPlywvvK9jGjPw/Cnouw7mjuI225vA/X1HA0
LT4ie+oIERSJsAKe2zwdSVsouOym0A9ArS33bUAtxOIGHKoEMGjUdyp+Hz1cDnJr
EdsFioYilyyfsG4LiU+koEznaMttTAAMBKP5IGZKS5rcl8T1lFEY+wDjJG0KxKiz
Mjf6L5MloK2frjr5HCUTh2zfnzb4Q269AxKG0jBKzmvReSYXOrGOtERiHX6B8MSC
KVPfnbZXuDaiXWGiL9F83cmNZlaJToRNyWVfboFvLXGDQpkzbFuo9knie7cY5rOu
5QKh0XvRTWmEvwcaOofaZzU5NIQ3UkXPvu2to5idKjG51Uks+wFeR6Hb6yxQimLj
LWrXk/iTVja81kigaqc+Jd/4YW+vf8ik3ddKaNa2I7CYPBuYx+4hbXvaGDyOdgZX
mV3zfsFYq7rniDbk8a17schHEOspwBbW5hhsP13EIs9hjHtvzNEgnKtiwupYS3hP
XCEWHCM9wxLAdp1eNxMPvY+EXgWWnofbLdGPsXwDw5BrBSRV60d/NTKSfyfntce0
exX0D9W3hmEq2gTSpSD5Jk5Ui992vanLX2kOZibN7A34R4j1uWZlb1yKnIFd9Mf3
LOvN8sGBAuAQVrzZflxwwTZvp2cPWVfH+IjZpkm6BimILX954eG5u0k8VpWwE58w
dyoelwyKK6x+e95ntVxSXWPq4/KOGJO//T4y/jjQhPX6QRxJhRaDcLusxE8TCKqa
/M52pSH0qYy9Ya/Hm3wYy1nxnDTZZZ5DY3wj+CM8/md0jN2LMCos6fAtRwQmXLrK
OsrAWF0oHhNIwbPMKM2XtG4k+SzBoLodyD4DIw4Qn8XPE/n1DNKgmklMhI/f+6J/
q4+ctp2jC2euKmmruJhDigf5LF8T9AO05ULIBtYLxCh8cUJaOsqlXgORgDcOpd2W
zNxAa6EWoWorDcKGMnK4LXc/FlhRr5zWwGtID1WvVe6J9C2c/rXGKnQ90A5B/ofj
VUFbSM5ZHC8CgTLuDKp1+MuFpT/EX4YHO68GKBiMRXRA9AetfV03U2gGgYO/bAMu
yCvcTWqdEsj0nbzNNhFakZ8YxwM3jH2jp8sicAZfik9wmZgAFc/Jg25gQYAbhcTg
+q7mERb7z7SGXeDr9pvfWHLEVBwQgox0zwO8K1HR37E7RcD3bnuuPxHy7RuSBw7g
L0/CUHJPVvacertEYVQ1puapkGZ6QVKHVafyutW8mku0sxiX41XzsWkCkVx90SYn
Kdbr8BULetGOIVx5RXrf2Ctya3lzAHlObemuCGn45xyDCU+GD1PDxSmOOWQqkXjo
Chd0gx/bxz7p6riezm7IPhBrEsmYy/fmbqQeR0zQ157ElWJLn4KomJn1G7k2mCdU
Qi1Qh3gEDtcZ1Llch0QAgR04c3F2csEWGCJpUnbM5oiWtX3xY7+7r/hWHf5iwfE1
AC+MAGdBzn4tbDULbTchNuEJiO3zRVAODoTxZKUamJYNFTTS4KYi1ElZAWMb8Rtv
HqCe7fWZSC13tvANg/dwaIEYQH+lighX1ZmD/yES152OpJjpgqtMpcT0Rnw329uM
RYG1u+KZ8+9bPoRqR+NbiRTB4uelErWBPPPlAy9iqlnsbyM1KUP2LJTxQcH8oQMR
RDsGC5znBXKci6mloiC6NiRPAVrH8haIk+XY0TJLmRkFJO+/M3J5j6MxmN0e3bgw
5QlZ87PpPNGy2RYdebCLAcn4pYol7UUOfFUNZxPOJCvXIhaEP/vfapgYkSL0cie/
0ZnM0PXJtSfLIMD1zaxkXaUjQnPt39Woye3KEgUS5YiiowGbYm+hqvpnGhnFXElh
B0GH9C1UM98jrSmarkIQ9CPcZ/oMxXcEyj2WUoFB7xd95D7m/wuSAnhcG+SZwh0l
0oEyqHpP/DEd2wrYivszhbeGGhFzznnLJq3Ceeaviu4CWND4q/tiAEFB50eNnU4j
LJ0znkaa4524J4HwOTu0UjhPRq0kHh5SKVgaR9wx9oWKXYJH/ZwL0KXDHkbST58d
w1xPiGiARw1EqV+yq9+a0TjdhTk7x5Pxn3j9RyDVIHxCOuhCdZYFDAFQwleubo08
dE1PxFaDHm5+0r+DXRIK0lt9ZqnROf07sKLQM1NuB3uedU5rEOm2J/FyjpVlCA5w
f3swK0Z8vyjglrwusryUkrNjBZJ9R0uob7mt8z7002uxurFLsRaOddd0C08OXRf6
GAP+a24EZllarXPAglwGX+GIkmccZcrtHCVUEa2tmYDc4HQ5BnCOBFZUMYYfrPb+
ISL8N+MJyv2Bp7o+8/v/MUGB7DT2tnksBlKll0x9oi6EBaktyQEq7+S9JPshb/yB
Q56YYvh4jeMe+rcrivd5I0jiDXLFp2mIITXJWYs9FucCkqRJBjisrH0ruQOZEA9r
Yk/XE7TfGZToSkeHZrHWEEy44PFwGNAz9SfPLB69ZezZL5+b1Y5xA1wjM+LMjKkB
gIAGrCxhtZh3DJhv1E+xcii2WMm19yfX03srmv5rPqkQ2eEPo2EVDPUVDy3tR7u/
MQ3ip/CpfGR+zUfN9G6gtV5lxGM2HxtL9xHSFRf1uSKDnIqcWlO88g2bfHaWP0Fn
kOiiuzgT4K/Ffev9a2YDkqkLkLwvkEy45a6UNFWxR3pWecM7jFHMgEktUuaKiOKb
pTp7pA+VQHQCBkFuCz/hujEA3FrQpqHVGZv99WkD8Jr8LF7VOlhiTklDYkGYyv8G
Vdwq+foIRUmlv001Ivho9V/wE7rPR10TJvBueKrfYCRjmFuCsT0m6Zz/AbuGTcdo
Qdqxjv8LjKGkGH3U0wW85f5TEIomuX8clpjrbPrOQxfZaLjAWmo5E/urP2Nh9VZG
odgzDK7gEdfs14v73jWm//kJMvs9LdQEwjBZKtlgoWKD/3G9M44tMf2a4fHq9VgO
Za6sUsssZis1Cz3Gbhm71Xb07Lq3VmrwgIb2DaQUIyokjC8W5+bxlB0X7XU9jtCb
24wry/OMgw8Wpi+/fhtwJLKZXgQ8Inrrg6O1kKSHANnK2nh8D8D3RunueP3+NoaU
tuWyf16h9VTvFfsZPYcJrssQ0/u1SRvcS6saWTKd/WEtnJoo9QM9Oo4lNpRoeJYl
jvmjWZ9zJwrwE/gGMkO2Q9UV2z1MUYCDKNkrxwUSufO+The0iP20EJP/+4KAjnWT
zuRNgENsOKAGoPI6csjzXp0Zy8DmDQMx2Mm71EwgEwlvgxVLqtZ4DKNg1qhd8Ygh
26no3HV1BuM1QDlDuquYSw8bpguAtzF5+P/Jr8QYKG4vuRAH22rXN1RsyXatkJWN
mVGGScGmBcp6XkYmrI9Zq+o/2sFmbVktpxXqlYhi6S3sfuaLUv79KV1zm2mKJ2Hj
nCs8Ey1E8Mfh5DgsV5wWwLJZ28SpWG2xGYCSAi5ZcT+ro8SvMzUPd4RGUbg/oHgg
dAF9N8sXsKbW7gxkMloSzz40xR+N/ygAeM6DtfbYasuYpHwTN3F3rlkJqY6kqgdc
9M9kFsl5dtGQAExwGKe1pBs++Rquo5SX8js43UeaVprxCrfba6UKrSHcSeoSxjtF
tOIfVr2tEP2qIxxHgDRj6yb1aEgXphfhBBUR961G3D+ninmM55yMvjzbVokYNu3K
Xy46mrUsSwq4DGRBRw1gIh5zuTmoyBsDo4XFone024qLQMlQxEA+XJe9dLhp/RNd
wucaxIlcIBGvd+pgjTNvryoMnG6pNnNe67cLUBDcQ1X6kXWpuG2xEmnUfAMeMsaZ
HAXRfnLIHLIoUW4VRjOjfYeHixQzKrhQkMKEuGB3x3e2g0MgM2PPLcw8RsyzwA5I
NvtfmEHtxlN6UIVPf3bZw/QKylRs7yJXK65L+AxH/BPM3LS3QSEqABXCVqWLLcI+
pMuGAMTKzh881hkdzvvZ2kEzyltEyw0UtsEjMteUFzCukmPZhkMzwlri3f44UtII
YmYXd/esQSfzoNVGznFts2q0b5h39opJo62stu6DCm1LEIuOLcpim++rxR06dCjG
Y3UzfpAxhF64LPdBMpHu+x5RjfFezlAw5g9Mul7chZwZe9Ilf+qg9ffDsQmNB3gF
fIp6vupjrYzuJd4eO509J9sgjsuMnI+5LNTqsDXqopXmsU914mD0HRS0gUU3nVGH
NM/7NBPB1AO5DP7UCD6gQzkLt6BPZ3BkIvehm/spYx+V1Xr3oT4KWqVJvngE/ZNi
xWuSqmek6nDCJDVmPSdZGTiQH566xd9H1MlouA/2NmsclShKR07FMvh31o2KYzKa
c5Bbrt1IBnwiCyVMec44+sU3rqMvoVWrKv/0oAD0jgFgZayoi8A69cA+V1SCKUju
el6+pOj/cZzktK8PxPTGqMsU4RcFFcpVopa4Sq9i4gzLWVFLvW+lLAEIps6QitO7
lHQflgiIvyLjMJPBszDTUj3D7W9e4W/DwD1PRMWIBboLT0dsPCOAmJgMq4jtijrm
6EtFedR+sXhCNsj1knGQ8vTq4LED8GG4c80B/o73smr5OsDpjTOsnOnUX5ZK+V/8
i3/jWT3ysxSe4NavAeE1/YLElYIMuT33HDhaObvszeehsl4r6FZoG8TgyMk7w5wx
DCizLfzMUo4oiMMkqJcAU7eI5TMyYMgkg4RXD/ufbYCv/pNQ040KWBEhPknCfmxA
PPJoZ53xhbVCzpAsaOFjqJeJAlQc/mk/hy2FbgSa0BDl1yFg08qV1tYWcxHNaY+O
Rk/hWI0XXehas130H2IO3A==
`protect END_PROTECTED
