`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wllavkw5gLDf1n6cHs8cRJBImX6knbDyOAV1GLKEGZ1RRQoWdDr+yx/obXBriDvr
7Bq8uZ9IpWVNod+BOAXo9YFV1WJnl72wopNvhSi8e4HjoFLwg2QM/Tn6TWtxGztO
BMu35UaEVoPheLvEMr+VGdBCkimHSFbansGE2S8ey6GxAQ62+q7t0WbGvkBuSjpz
aschD25wIdxHQxoMXd212vF7i3F0N8BYsttgrG+Op1kcfwmPyAf419U3WiMdBrGi
PMlQd1QyJAdpAi4hyKjfIlwiNPyQ3BKpgU79IO7253lhUYzzi5N7vUnaZAlG3SB6
tXOnrStAXB2bDSiNknT76JGg+dcfdlQPLJInpuN7pu51ILKir+haRcJk3c6B0pQ8
JHlzS4MYZx8c53W0us+9nhPtIfYIwWmj7KIXSSHrxuI98lC88xQ3t+3xq2IhovXo
`protect END_PROTECTED
