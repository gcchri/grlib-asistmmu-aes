`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4rS91tOkIBD2NlmmtKe+xs1im0tL7qVQ3l+YqEf1FY81F9N47qSZlNySOMzM8h6Y
HczHOgbt9jO8VRqlxcUtTodhWh7YlOyMt9BUcQ7TmkdGm2JU2pyDSdtWMwFCOVwP
AUo4c5iOLJIdneOvc9HId7rl0s+Q3Na+0lJ2qokh1Taf67u6x1jAgDXxLN3zAhWU
ulZZgdDy3CzIPqlvrra5TkJ7DHfqjagVebQCC1/+KPi69fvE9V8a0EAt7eyGdndN
4XvSNszYNyqfGpnERuS5rFhkSpXxkGBB6h8antMCM+cfpsJ+YtpouuA8IhjkKsA5
1gSGNaLjiaAx5rYzfqWRUrbmS36HSoKgWHGmVIioK+mLNh3r91rbANEljEN6VV7y
GW0dOpeNsCO5oOzW65eBoqoKGeSviHw7ZObTYCq1eBRZBJ1NwszgtTdvvNd7y8dw
Ja3MDnu0/rTlVZdxLiynlRSyyrDNMqQZtz6cEQFC93zZvy0orcgRL6zRDl0LC1Y6
rvpen7dsH4/R7fSTLj6ZD4dzCPpSMS5mdlXJSoqWciu+TCgyoRZL/1DZQUAeaHHr
y3HdglCVf/PcbM/6vJSU8zp7FElClHclmEqD6SCZrXLMyUMQ8kHwyy1T4WHzXEbe
4yzldcpDp3vBR5XNjt8m3bhKpvXruJgZReRE+IZo3yhrzjdKPb3FlHAn4Tn6HMHK
EanA4aYdeoyWyjub7XSKxF0Gt/kB3whINl1ETILWM7lhnbmLKdg/nuHfZCBoj/jU
0Xm5ks+MhdMUjrZhD5Lxgg==
`protect END_PROTECTED
