`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B162YFRLXKMtGjyM7BILOTOniLGopXsIRv85hl52JhSfeaFC1/sEIxyHwQ6xK0O7
rbsENnDFuL4Ete3fi8R5a4oYbTWG/cBBccHPFayUqBgjqW9YCIcC32WQ4Su22Rsm
kjO87Uwt3vAxbKOnQJ+dh122wuIbKVCZemEwrisovW1pz4mlt+Dhtdta5LsquSXS
8bzp7JEcFHoHbZbQSMm3QjoCHjskPeVUNWkPArZlmCfNCFfXzswV8AZJbRuhRW4y
Iur0A46PNGMYQSZsrP4rdprRPrxAY+ufwirTEwG0cMG9pBUJOl/KbljCtGNMayW7
kgABtrj6bq928KSAd7abyta/G0o6B0W2GaPlto5p4WQ24JRx8sZw6HH/KTkjMZau
fbi5ZEZhzKhy8TY8JBoBbI/XdzZjgx0FNyGsjuUJmxRCkqqU08ySd9n4hw43WlNf
axCl7CVnoRT4VVr2fvemrUDiHLh0AbjC+AGw9Ce+MZBLRCUbLwgXwoHPmHfdQ82j
`protect END_PROTECTED
