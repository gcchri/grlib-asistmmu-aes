`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
37F0ubbGyLfQ5PjOaWYWe3CBQPVPPTiIjCICvI59pFBXvi8iCzvIs79H2IPVwVjy
TJsCOmcNLKNBdHz4Jq7G0DpwzWWQ/IBPCg/JxoHt/015i8+54eaiyenGcuONreyb
95xKUzm92FUq8U1Hb7OLRMW1DbVpnzyUj197Y2Ey0kuWHqP25rC/9o/dJ/UETesq
R0CRwkFB6fllb4K9E5ToBmx+Pp1B2BQdz3fo6Mmvuouu1IP5hj5t3AL5Q2RLERzR
j5Rz0XlZBklLaHjvtfo51A==
`protect END_PROTECTED
