`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AIc8bDeqkYT+VHN4SYDeUC2wf18F3dbDXP2H9XbsTvHmRV0/ropyF4Z6dG+Dz9xR
rSBWJKaEtzaaSXrFPMJbCYDJhr6peNCwy5cmtt8PqCvx3yuzOHqQ/SrEVQOQwo4y
BD3KxZLZANrRIBwbHEcAwewfRxrCWKxb1Y5Da4xPI7J6qDIy7ptzDQ6zHRC1GSbQ
V31C8D3OEMU+7zlNmC5ozXL3GS72bYN1NczScOJK7nj9IhRFTVyZDlkiaCEuBkw8
5aeSNrh3gPIrASx1d2iWHVziVv3VzPUNWyXSdDnRioSu/tDDU8OGg6nN/5i67Al4
eq2n1tuyUyjfCuYEMk/VHKfEFjmh8hsHws+TSM7P2YARkb5TIL6qyorGIlqLWwoj
Xjg/eR1j81jRkdYHwMhoiz24MqR4F9+wFiXFR55fQLvhD/Zg9lqOOC+yu/SxrlVz
WwHjFM4FNnIuc5wbfe1jNLqnDuGHgKcPu271T842e+HeARsoSOEG4F8vFFMhqLWA
4sXDeh3dRtTOUco7Qq2yTapx08iAHgyu06iKt4UBcJWQkJVu8gAyd2oXHswX8LHT
LBkjcPZ4pRq9WyKPcN4KvvBaynTX38tV5XeRmNS8V7Hc8T1tln4t5Al62lYd9yWa
xVKKD1MmUUiP/w8YRxbU6tZUK4mbZXAX4M3lW87qs71efbso/CenxnUy6QgTy8Sq
e05huJACdiopGRl1fsOS+IWNElICyXAExfXgV3Rj/Vqcr2sgbmP5p+4Uire7A0gt
jWyZfwNaZiYawLV0YqKCRAqdKupySQEdLDAsoAdyi5cFOQxE2O0WixWX7PrAyw+4
Wk41oIW7y6Q6QjspLTk/ROD3U4afxD1uvpcpUeEIK6vE7GGGgC95gfsSS4wyGji8
4x5MRaJks7t3nMzaq9OuU0MtFWnWeG0s7wUmd5zJSDhKhqP4lgED6eZ1fVv7bO0m
kH5XLqBzcu1Z5CYG7ERfQLyt1wU3wKTLnDYoccOflPmMt6vqb/4W52wVP/Gal5om
oO94FJCUiQi/ebsZ66DdNpYwk62rCM37+GnQDecRDdUGvJtJgB/YZ/DLU1ai19jJ
3zsT00jLK8/JgdDz1pA+dkHqEg+O9nDJ7v5H/ArYOAgXyR0G7C5VntXt+mcNeO0E
`protect END_PROTECTED
