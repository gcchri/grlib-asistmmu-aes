`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qb4orq5/PMliLfr5+PCWk/JFdr5zuH5yuUbF7oDxRK4zdKay0wcwOTR07wbwFQwX
t7wripoqnabPydLPjnTigJu7OhwzpsafXs6xmbs+GeqU9UCaKeEJf6UaFHGIs7x6
lDAVLwcmPg7iBGJRAYCVH1avJv5T0CaL6TRaILQFVcAtY2aIwKK6BC3CmeEh3Gu7
aWXEHZHvE8e0MRrFo+n/Bg8peMOCKAplQnIIt8cutEe++JSoByTbvh+N/rr+Lhq2
ds4cLSApCAPA1jC2fYHTGItpABcIVZBdHFEoDtUkBB47bwzVVDIfzLmbouUuoXi9
2FqGCBkNLkKHTdX99VeKiGnzCfqpahRYrbVGeH9VzSWN9K5u8CiAG6JlZWlhIHCa
wHRwSWFE5kz1pYSaWf6EhLNrNFBGOuUFdg3H/huZoZ5bW7IYkEOcQkjgUg9IjAiz
`protect END_PROTECTED
