`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uBhHxaF7LrNakQxfTdRFCNJXoXFKW2e6WhvzzZheDUg69N1ZR494by4tnNd6tQFL
hmX2qz/DCdk+hEQ4LN1YWVu9o3buvGxNODCPeJ0zgqo8HdYKHbEWskkPmOD1ODHw
3M2rq2HCNxT7vSDkj5779T+9Lnr96+x44cNz+eh0Jt8XGN8w2OC9LyswqpvQ4x1Q
/MkhoN/a24D5MajrpRWzVYfq5Y1Jt4psoVg5h1lPMKwZd1XdtN4Ir28e/Kei5t7o
DFpaBwBZDzZB/ZujtRUKRp2aGOxzpbz5LdKySi7kbDWSvkau0ZFJ5Eg8xINZbXtY
6ac7Wgd98NdBkLnldqT/cOENjbPYqRCoG5+NGczFyFoKNiGQ4m6ylmFi84Bkrudq
tCWxz5iz96FR/vVziNCARsQeNzDvI/Te2hvL5dLAhAWeQhjeRHWhEqaetxbQGCi3
+JsjX4QcUELO5K+TLS/7w96fCJT73mQTS/LDka7Q6edhHzcaK71beUO3+tRRU8du
LU5Px9JfHThOdFHajCLBwEB2GdxUhG2ZYAZCyzEZHudEjTRGZMUUDx0XPn6pUZ8v
aDLfUA3lX2xUGBgwyQNLMXpDUtd5+DSYJQJZ0xPmE/wYQjMDJE8cFvc9gB9YXYte
`protect END_PROTECTED
