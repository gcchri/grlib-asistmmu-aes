`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bUQUOXAURD4L2EOhob7skPro1mzSWWusZ0SRRNRdMXZt4FJALVEggfQJtEn4xvoH
Byf/wyASlxeOihgclrNN8Cs0OnbvYCHC0fYUxVAXD7rs+UGmePDyff3wTTyRnLT4
FBC5XOYwMWKzivFneRivP0hBsWxp4L8Y2n2sqIOqjSdnkN+f0jNg9MXCIKZwg2G7
GWPa1k6D7d4UOdjokWH2fBfAtzjdIG4xsCkT7ErCGVH35BbldWZBMpf7ah3o4b55
PtkxUdoII5C1Jg2+igOTLl8oSYjaF/MhrbYBMoK+yCYUAdew6cnAe6o1S4HTBBtz
tXrceycTJitUZ4tcGLjR+A==
`protect END_PROTECTED
