`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PJA/Jg86NYNFeBrbIy9bpHpbs+fpvofixUttN58mZ3pZKykEzcnY8KAtP+uFzmW2
D/GJSDqpJlT7bqkOqIw8qZFxktobMttUELJELLjqQKE+zHhKqWMkeP39nXCMmK4X
sq9EoroK+SnXhlRxdql7ken4DRkIw+y6ltzizb0+fHkZW7ZKPc+w6fAhTvmABdbk
EuUoNW3Md5J4omVUKfl2JhI7QnxZQ5q8Ap/K6eK6PKmjLoAoO+HhKxVODu2iapPh
WYCFL+Oaf5tstm2XY1YCYrazjsSL4Dgfb5c11HPGaU4INGTlRQEI0f+0Im+ZMCl2
wkT7ETm3qY+iMfy8MGAQdWTNvM38T/LPVRLVPOyRBmS9RqrxBolPAzvw1z02WRYM
bXzPW4drZ4DRgKdMzaXPf4nVfGdz/7poM6W5LZIhBaUT64zXhDA5xVByfpPPqTrE
`protect END_PROTECTED
