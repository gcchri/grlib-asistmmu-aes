`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JkpGEs08LTnG8m01eONY8q0kX2UTq4HS0UcCzD2yBSHCBSCKCIMLDykPFGsUDxit
dp44P2z5WO0/PlPaAquZLMMfL2mIBr2SPEpCi8puBUbBUWBtFxI+qaaBZ5rXfYv/
d2DUgeUEF1vdnvcg79ZJ5UQPxp8iFboI3pOP8th/WWiQBau5TYYoHZGDcWxgy3JN
EKOLRFdmmQxigNbA9LNpfpulEd2NY/5g5xf49Ixxts8zm6vbUcvaPK30gfQcLm61
Rffi7T8ZtQh7OCb19ggSINYHQ9CvBwbxL4urN6iiR5nfQjVArA65cwmNxB6LvYLo
koIBlEDZDKCszIL8z0h2DyS7ENrhPTMIgo8Rs14N6nyLGJ1Uh1Ad0Si6aPRwM0Uk
mQuRnmLyVNf+q9EVSUZRvzp/OqdelZ9lCCoQMVZ+487j65UBMEUFm3a+CZMhHo55
`protect END_PROTECTED
