`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OuawTZtp+IDjAqz7ITOU3+LccX3dkFgJRlhLfloz6mtjLQpmlJN74oAmuj4DlEeI
Yp5cRQi4c9McsCWvRqopKmif4KLqx3uh+KO4s6P+80Vci4JBe5MZYAheOOAmboeK
HNaSTtrT3/RrBs6q6HwVcZkAZhaW6RxZ3jXkWleOpZxG+C5lK1wy0osS0ineVnbG
fgy+YZ3jYvOShiDaOqpCz7BAXZXPq58a8deTOI+YoDnSlDWXgHXrjQdEd0rscz/A
AgZhCg46AN605v+xgjTQNoiCgniDqT8bofKS4lw1SREwjUWnojp0K0SOU++1fLDp
Vi0YSEApFwV2HiZortgyxJjmurlR2tSmOVBFBXNS0hnbDwkGGW1adzFqllelOs1I
ztQ87HNYBiUT+OF3lYC3R1mZxF8lebdVzRpzz5vP/wsL4K70jZoGZ4qJYj1aY1fR
pfYsZcklEWp2t/XRqZhQHcayZQmebE0iTfd1UQFkXhClI+7ZuOvxvltS9GEZ2lkG
C2vJjTia/Ftv5Qa4IcohnhwSs8IQD/hhAirCa/0f4Ml2yOGD+TRQG/T1/dR+QpwB
mLhT3wjkVq3k1Na8nTB+zcBh2Y4WYA5NcJ+rn6l03GJwHNbGL3fEL4GKVhztvK2W
622g01YL63soJKeiQcjYrg9QxhnDCXzT2WF2kK0dgjWXx2a2VEH7FhUe/mhMFzcV
kcLOkcV7q6MLSNGN/krNWUh14FMmHNOnLL+hsWMtAu3wFJPgLcouIsmJ53hNfU0/
8FOkog7k03Q+EsWCz0P5D15mrADFZx7cKKRm2DSLaOyNoyujKqVaMsN4BRZdMiTE
hXS2eIz7t4dtjeY33tgUWP/kwi6yGzeC0shRCiDjCfkrTbVfXa9IN+awRYqFYSgw
1zGi63uvk4xvUas067h+IwIuIDo+z74PK0RZk03+XI/MfmvPVmj4v8tYyf2ZQvLq
sLhFbX6ePzWvYGx82ygWcZmoGTAntQZVNXFRpjhm9rEcWlJ7OPH40yO6pS8VQ6/a
WSTHKAC5oOvjD8Khr11luIhmkWnQ+t3weqZHzAJuVUVY9IYYZrtJo9sw7gOAPrTW
`protect END_PROTECTED
