`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l6AEpHM+aGDEiU3vRRxKBjtHJ2KwmoJuXmKcstwZcC8Pqg/Hp+lF3TshEuHJCZqk
oNwfZOoKtoM3Hf2UTuOFIfvHqVFm+rAwZM9wm+ZEmm3fP1skHvGC9PWRMfakuFHK
hQMpS+OhkTCChWb4q6K2/MOsrAophBgaIuDPppii9oHafbWADsD3rls02d0El6Jc
Fik5WhMyTTmTeH1UXV8JqBYN6r+SASDBVSTsPZDB6aa3pSPkxvJYwy6GJPLw0Z+E
PBoqZEi/fmjpVV6GWbRQawVMrCbfE6qMMU9ztDBlloiHSQU5HbPJLLjITuuiF9ol
KqD51N26ivB/0RFk/zkekkSlL5BuvLC8WWpwG4LoXOawelw3bPTiM9qQrOAfD4up
BrQb2rY4KxhTZcy5y3iRPXbKRSWzdYdfI5uOSfZyqGFJHROYdCz2JufXk+vyQWJW
R5uvoHnV4XNPznw9rUCeKAEMzfZI/YkuZ7laRugQ2cmFuSSToViane2HgMtPdMDp
siTyKpLeu6cLwwYIJZktF7AiTO6fGK6/vBcRUyYwm5H43Xs5TYCiayN8ibYuxZpy
YhDuga+cLXyhU2m8ApTLinkM/k16mNCdViHVC6BptDaabqO3LOl/3Tq9NS0gmnM7
+DJOHLfBQ5Ol7DFwzkj869Phj1/OB5UqjwcAXvFhgj9B/k31DwX0JrHuoneILzdY
CaJKnz6zB0hXFYNCvehdDgZ2bUwpYx+VnFq/HI3vOFTXkuAagl8RjQJuEeANOUp1
8JkGmesBEvBQjZZe1OB9l9nJ9ReSZQ9TaS8DWbSOrVMc3ljapBrKFC1mWUoopUGv
KPwBxBiVGw9BwmCQ/+lNzBP2L33om/KChUD645xktU7qpcy3fo/B1SP2XjL507wG
A6G8gjDTH7RGiztMBA5hdZpIoYiDhXYj0xC5PjRJftHSFJ7Tic64l9N5LOkqXTHa
njYEcKi9w7es7sajhWwSDLBKB/tjDvihxW5BzIDzzwmVVNp2Cqpx0+KWXQzOJ5fQ
hqw9HDmGRlXMGFe2jhteaA+r1XiTR/6l9kvP+QMAbUoQ/1U905yKf3E3PR8T4Ehd
DQxNKK+avy//Tff2N7tWz7GZuxlEx4ONdYLvo25XS/5PSo3LpJ/9DwcnAdYOymNG
15EyVDAJ4N7dCdRsS6oKaKVtZ9TqVjONz33yBUbPB8Rxyjhg9N5lgXhfD/CsQ+BK
QVbYJ4rgCeTm8SR6nWX1Op6Fsz/9NoLJGzb+VR7cx0+DlElR/gT5B12dRfgLZFKz
BMQDbuYykSFVfkWyXjVxM+N3MooVRsh7Z8VuacvFdRCusyX1Q4D8WV3xA6yUbEPG
/ioxbnMJ6dEnYOkSBgw9vSLeqQQmGH3FZZXegkWFkY0BCFkCmiRa8VkC63blPJky
2+BTp5qx5LVkjWSbEgjskdQl/2rJXmpkrVBqEotu3QOc/qU4OUlJbRDrTaFXZ3Vx
kqwCcHGTZzww+E9w4cimfmkSahsxkE2cKUfWGjWXKnBBXRDy0kejY5vvTFHmoDO3
xlK1d90XXVFexcG86IFVljLh9voVZr67rgJ5qrrkIELsXDDDx7tyHRqVbtCO52U3
KEv0AhshCfF+wYZic6w8B1bONq23ib2x4X8i+csrfPV/Y/TiBEq8ur08tmeP8M7F
Y5oddFEhWXV965CgBj0yZvjxHhMsB1ALLgqX4HFUmwIppNRxUmCUzJHz3qFf0nc3
Y68FuMbd/A38Uu5sg849+HY8Ff+DnedbmvYVfmQy5g9AnoI6IqxH/ug4QFWpEam+
mvcyIyDRS6shHgcXl/dioifnXe4zizgtY+C+X7CXt5yUjLK8tCSZl/YQXl9sXcgw
acBxClMyol7iNOm1aFmhSRIIAQQInMZF/6ULD/mg+itZ5XjXorK7fyu4nOrm1JPG
6sBMG1oJGMa5mkCmvsyTlA1IxbRrAyKhG6zIFEUPFfC0HMyAqciaa03my4PLwPCS
ETEtZldeHHtrsHVJe0qmwZK4EAWZTmjNysIHpNKhKPRhLwK2MYAEEMvIcFK9Ng2J
3/DcWsUFKQi0/peSqugQIHhxvXxeoq0m0d/XqPVyQ3BINCZ3POg95eNsYvEA8sSZ
cZUp3r/Apa2r8R1SQRgfw4sRgvHDI+Lc6ySyUWdBnvgFO9htPeDe7Wg0K2N+VdAi
eUJsT9KXfmQh5kFbt7ydvft7T+lXwy80AXO9Q3eA/adG9XbWmK/IPYhuG9dqknlx
1QVwe9U8X1hsQaWmdroabt3FNgFmh7ASXc1PQsgD6La9VNgLy7pkfmTr+COMAinQ
rNJXhL5R0haSmWfSPVlK2mE0KmjSBw7vKuXBrtoq0/IYbg9tOnRkXvWjqrJe2Lzz
ZOahOH4CQWxmN70sz1JfR9rnILdDyGUe8QO8z/kpna+x/mxDMNtftnJ+Puj5nYIY
TMjlsyAd9RFuhXN5Sc0k5nD+4R85ZlrHw0QUwwyKk4264g4Mst7Jgz7dfNisi5aj
gq+Fmg0/zNUQ7eKlmjVjE2Be/m8Ha8OKmhrw0yZo3hn7aLRqsrEMpLfxCkbOjECE
2KWuDWPzEIj/mJciTmCyit9wxhGclqSdkWJuZsKTJhYZV42iisW4iS4o8pxP/yHx
veoKs771JbmhSnI6lbi5uNvSHdCQc3+P59/PPAJxUxJ3Iz8J21KHvOoWvU6ZbMre
eQ2sz/9X69zYH089/8xiLQHTS+wsOpeLVcQIB2UBchMjscJjnI18lR4Q5WWTKl+Q
VlNDbp+hUgs/caSkoIRMbSpiz62kj+K03MhAokU693kvzU3NJsyJX+163Icb22T4
+uMNExlkohCUHrsF4GB7PP/f1FI4HJ/jA7puoAssacI7k1HMHaD869xpCNFn23KL
8xqVelRYi+zHuiiYnT0yG+c4lWVS1dXh7q0+GyIQNZ706WDx3LDm+YtY5y6pM1wH
KpAAKPcrwxNjlMb602JAlGBHrTezzMPrnwDf3CDVwv0=
`protect END_PROTECTED
