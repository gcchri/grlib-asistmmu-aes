`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PIiUyTWge9CYodTww/bp+OoGdL52iwVSs5wkqvBHUF/5o7HAcfW36UB8pUmwHxr5
axEPm9zdWyWA3U1PCUD/M2WORGripm4YXl13LxHABi8zO4wr/kDFWNZ4k5Eb4wEM
znHA27PEd+1LjgiHHIlkiRE/wKXOuiNlgtOUSb1YPYOxJ5zWmAhfD0HY5F1XIkMF
CX5/aT75ppUuLYrZcdX3B7b0zz7CRhxjjmrHcRxDulnm6Psa+4GFyhDK7W43NkxS
FkvgJDYyInMn9MyT+N42DmJa5zLahhqLkPzFmUeCVNL4zcWm2hjmBDh750wg8JpK
ZcZy1PPI4K/l2WP5qxJmUYtb6YO+IkvPNIyBLC3qoswgATqxNmITrNwBP4ceWUi8
4gc8ow607518/rLUMGRd5FU+3XEeMlXru1G5q8t82FozGTL68nTkkQZ6uMQg/M6/
yiEJ5Jixsn5Vn26KYp3aK/1O81Ve+/o61jF1V8gLZu2Up8ojgQB+NVIAYp08p2H+
V0ZVIvaOjMXJTd5M7H8T22ZNJB048k7Vy/WBU87KHl8YoAL7WdcOR9tolnQ76Ami
TYkHmdLNUwrnvEmncb/LdSReV6wemYsz5ZORb/176mZEbRcGvClOTbFdxCvceLcr
7xpPJISXkVA3cPTvDqan39eN/QJv7jyEaqn924B56wPzvUQ8pRuJHXQmREprPBXq
Ujb/ZtI3QeIjCQjfRvqTPCN6aDhLnVWxv248uO/P+Q0Mjhq/XxfmmdgFYV+m3K7G
cC/qNud7q3tj0nuH34s5Ktfh13Q8oFDKJue6PrtlFPKBIKmi6lxVrIaWaiVLk/rK
Um0loiamtDnk7jY9Yfxrk4wfmYqJ6bM4IeG+0DIDYoLTS0vJvIY73kwm6uDGBrQV
1G6H1xuuwI6vDNig+HHLi9/gS3wO4FcZMQ7zQMbpnxye2CTxOfGPUBk/qySPiAYf
xdezivQnheZ2th7FlakIqMWIo2adKj7No1fks6SyMUMiyIbKF5Z/6mxy08EJ8Yjv
sATMtYbU1oO/Jbau/AoYmOtfVs025uM1zklNdQwoTDiO9fEF2qw/W4oHfgE9/aRu
ibARjOz/Iv3fmtr3djC3K3+gA2sHnQiY7+Qx89Q+64hMUHQ3chc+PRe2KMNr9lUR
cx9jvh7gV2hobuFOgFq/owmQ3Ip5CbnSc7WTczU6oTkHjkva68woPBzW4DoJg77O
pvBqqu9NBzdPk6MzVDJ+KWi4zg7m17I7efe2nzyJNrz6k0lqQb9d5Q498nUqgWAq
SXbqJYNGpZwWX5M4Vql68FDTnoQIeR6G9Dc5K7DOAXyfveYzvmVVjQVpuJGnT+eZ
DW/h+Qd/cp0X/sXPDk9rbKsjQAL4gJ7U7v1sbGvBNyUtKTNAlUio3NK1ZIxIhxjm
DO4pxboZ2jgH4amUzUAYhm4/xKy7Q3b5YR7OKkGa78g3mTL2F/ILdGrg3qIFblQz
9d5czSksvOqHHKJs8WSZxJ8nQtpRa5oh3aNuugNUEl5/NG5mEfflIEECJj2bdxvv
OKk8JdhCiH3GpJWppNRtCF4gvwyC998SjBDZsz9xLPM5B9DCN500aTF7zKBl9K49
EJnULqvc58ksuEbQJQr/ePgVWSEYb9FG8v4kJC1X4fu6oAxAOiiY0bZcoWePY0eJ
wrTaTpkXGwebkIByjESfyLSfygEM/WbVz3L/B0IFnzV+8n/q17aNeukajw3uLRt7
AjY3tck45JULzw+zngTJo+JjLvCptqHr4eMCFOStiRAPByQ06vhe0vb7qihP2XK/
JKx6/bs9SDXVjtR0icgdAvL/un+V32vH4obNMclgpEBpcWkCR9nrUmnrbi0Y27+s
y+3gHgqG1VwC1ETBbLhWdqpkppTEwrFIQF8aSVW2QcNptdmsRcaGy0+lo+qiCjm1
36XtoGWP4r/pj3uiye/uSLCRn9kw1EWBxxK9FIiojeB4M5IgKSHYwIpsQEZrM3LZ
WeucgO8K07vhPP3bxlRpJeZh2uzUro8n6MkuuvpctO3uHuhuFB+7xNcpSbuvKnr8
KEZ1Bw5jWa6ABEZoU2r8VdYvpKgQJgGNbwiYYutH4AvuuOoQmltlbCsj0QkusYFS
pgnCQ84JUuQjyXH00NpPE7Dqbh7cMbwiP3Q4XU46PvURiuvmOPsO1WIdfZmkBv/f
lbSe+ocJDC1CLNu6zmCvfCQSPiVPX+zZSijTvvGORDe4aqYp5qqN1SKHmS/vKlJu
CuKqnhofuVd4xoBNFb2FP+FKWNxubxpvNkuVyNHWh7qEIvlhZQj4TFrmVe5VdhAG
KepkkQDbKGB4yT5HixO3mHL20uu2NOGnFJIJEfPgXS2EYzMGc2ZoNKdTHai074pA
XarkRvhTamm6ZxJV/KjNsWgGkjWZ95WsCDEv1uRcY6WR1+Pw5Dxt7G8ahZ3TS542
B1T8SZYEGXG/qkcUMSzfFcPA68qqhlwVD8OhuKerQMt05OhjRlgrBTtQqgDqj/bZ
fFZ4BFW0TrSjZX04y9vHpyvXC7uv/SPR1DqxWCx0TibKdDGlpV+z4btphPGHD45p
jAYLfuek57ZoN/S1w2P6HxTMoGzn1oProoPq4ffliWWVtoqFlgWluIsK4wGgRErC
FbHxT01ZBBzDMUWP1MMdJdmJIBTb/wFhUaC0S+6NjYobH+8qMa4WXfTaKnnXSuBc
L18ixJZ0JWJWTJ3FERRJpfWH3jk1FQPNkk2KgEzbsLAZHBktQynOG9kbXwE+COWJ
vwNX6OPgcCMFbGmnO0XfA4TVwj8QiXUpTIH0rJxtllrUJu5v5xVJSls8q6ML4U3J
rWQwX4X6di1XEF3soFyglHzQFg0cPVuowlh9sUwg5ao3u1KUInpLvIZBtebzKnaw
SqyMeJIGHmm1qBJyxEGCVxLJaifE80Dr8XnyZ6pFz4EfkB/OdcA/WpnHjyCi160t
BJdM5pQcuQWIADiB6Aoa24ZIWrEAEUlS1SD7nazedWvpQgPQStBewQH+rRY4v9IP
F1nQ77Kdm23wF3xwnhr0gTDhOtxQVby0wSwJf1X+4zaqMp6lMEwLl/wHCNZppHJC
cVjP2pStyzykIFEFTPLvQiHwfT7hn1j7nXdMAO+L+hRFw0yhsA4rK1LHwwBFrXqP
jsACKa9hbo1yA55fUBw7wdYFBo2wlWHoe9TGuXe09A1y3ZE5b3raHS8t8Y6LZCJ4
j/SXKdtsCe3VKuQx3+f9tRgzsWPV000McDQ6fy/RTK4WhZ34rrc+HJNmmuK+9UGi
SadUYoTsXMv8zERZcrDbN1z5MGYJlsJRsiOo9/jTSVyRELJBawPGTDX/XG/SaRDS
kAYK26Y3a47TH+MjCrRkBbs7w/hq8c6dUXUF041XFwxLjDY3ltxShFtfblkb2ZNP
1CSUnBtwQCgvsvPg5zaXshQdcmGhdyzJ+nB7ahGiMKN3HtQ0g28DNRLucaz5ck9/
4wFhdvWjs4tUcRDqFeS/auhxGggAp4Yz/FwsEcboVLdkxwxAgEUibewPdRpPD8ib
ddH3spQ/j/h/n74JSmxFIhTxlbhjN5MFy/r7fYAZ/bxFZCe3jnZPCzrggrKWc8Bf
5JPI8lZeIDlFLYcEkKcT7eePH9pFSu3qw5q6tAVLsBs91Z04OcFY+0wqtBlOzdZ/
wFz9LSh6nTwsxy1aFDzK36OxgQGJy0Vo/URkckgQYuno4djZ/8rK70cB8OkVY34+
uHhWx0YlIdmN2HVSI15PgRhrT0OynLovNOaWOyLta0fk7R2u/r65xDb7n6FBz6gm
SUD/tGwl2gwKoFMvw7F4N5V91fCaMZ2HV+J1g5G7ddfYebbTis+nWm71N9GZ//9b
ShZ5n90nB8Ossh2OvNSjjW60N1+27XCOo0yyGE0AQVJG2BHhu8ko/CrpZm2ppG7M
39NwBdWfqgSsLlnjsuwJM3FkZuhBMsSwt4V+WGQOBN+dCxQrOjLf5kufgappnUvv
6Y74bqf2I5udq/PguYBWRskWdi0cD9xq8tN8QEnfllQo6noy7UuImqk98LVRvj19
8q0AuIIyW807p6t3vXUtqGjNz8+mchEu5TfSSLprQcJuw9MzgMRCR1N7bOWje4K6
viZwfPi2Rwt9xA98GUPFCHDsrdNHFPUxGsWhC9gL2hKYdWzMEtPbyosZAeANfOg8
yYR5ThCmmSlE/YTLmtCwu+RjBEiNk1gnf+aT5jRB+sSCbDuku5fvJ6kEBCiIM9z+
YIcZqH3gGrNu+fY/yB2jbsmOzzUsyi29zGC47+9nIzeSOFKlfjjLYcngYv7clm/S
2uCMNmyrz7Gy9Oex36mu03+RZzVWJffbylyjkhq4u+DCd1ArujE9Nfdq9lCws9YG
cUC/ADmbMDW4YesCCtrCJQxZmlFWIGRmGyEgayf5uoJPNPnB+1mTnQoq/g3b0ghU
1zn98YY0tK2MSxeb1dvgHXbZNRI2QgdMQVZheltzFAEOPj1R8K4XmHkm95L+xJko
2/i3uox2+vsGooZRUzQXGqaC4qzy0TmN+h/rz/zSA2yLgJ7g23Gha8nx17IjHj9H
r+85eXoP72bQRm/Aw9cmgc0scjDXOWiIJqS8zB513JLZVEyaQzxY9zidhRcQFzd3
oJvfXDxhq64qaL/osKS7I9M/KBYPJXVXQc09zACYpWNU+kpVsmq1fS7LcSUwVz2X
w6kpOR1P6VLXMfJaoFXNcjFo45Oe2WF3K7/O6+l/hGnCSYSDsCBiRky14HN/sXxM
jzBBRgv7S8txGVDJlfN7bw449zJ9+L8ZAwotgzIOzKxHOONrTJ2qQaPmkgE8V28P
l4K/PoGg8llq+kFC/dgUcR9canrjRWhlJppJpAQQ9Ykh4N6lZeMC4LIQ+FV50Vl3
397ybgcRpOP5UtzATzs4bb5sczvFxq//9TAz2yi9UlzRfr92au7XVLaXuLNOvAXN
FSw5POkhslavKH9jzQZNcQhfiwSnxdCi0csghGTELK/nB8VldZwdBZN28dQ/PxKL
3GLmtVhRPK4kbrI02NiY8h29zfnf9z1Cm9PjQMIFDMMhI3YOOF27Wih0kG+RbQqx
atn4dAZ3O372AQfvwyt9WQfSskyiFFem7aQ41IAv7Mhik4ASeqD6l0HmoN7ljTs7
h9OSpaTyKq7NmSbqWQD4aRxrEN4E+cui0qgT2gPEkIMaSqGO6gVdxjWmXeEJhe7g
ekQTRHmMC2FzfyzkRU4JvC2C+6ARXT+CbrDKKzIzvItr/LOjNvIlSGAlXoNjC66i
2344h56tkEDFLemIFqswBIxovyGaTDaR2ItWnaURDdmups+A9InbnbKD1fjkymWQ
sF5Qjzy7cNLZ0V1xIaT1shvbyNQobVBwXzxwc5c8Yen4/yjbPghFA5IIytgBR+sY
MFwbL7H3efFhu8ejHa9kUMU83AbD4Ovg7FNjL4nX3nRFZtR0SX+Qfrzg58PO1CGa
fzOT3ZS7LIa/o4ARphFG7Z89do10wEUBPogpgFFujfqJ/dse7P+RB9bIqyro5osE
KyLbBmTlx1DPD3Frqiqnlil3SMm12zYwelFQT8GlfhS/MAiM6SNr4hxZJLZPu8hu
dD0G3MDzZqhTx2AkZkURd4LkeeGmdPZEW7V/nJKCctflLNxHIZ7PiLOGPeRk4qTq
ebHlxWjPnoIkKa1iiAJzjdte305fBUTv11nrJJ3DNnnlZAXFEq1/YEEnip8SOaGA
INmfdqx2oiGc076uKutDmUnV2bEn/BS0PhOEAyJTffaNvlJf2OpaClighpvb6ivY
PgiPtPRM+3mLObMgqKU//pV2aw/mF8COCs0x5B7sNw6vN+jCW54QrKqPSUWbgLDD
kRz3vJ5KEbcEKJ/eAuLLe+ORp9yin32RaoQmBcgBCkJVRYUqbWHVLrTmlDlHM+6q
fcXHHnKrEQhMbVeC6N4k2OIP6XPFnrfA0t7IweMl7vrbWi84MegfcA2QyBmjQ7VC
1UZqdwESe93/AJm0D0WTHExgmkq7Ui61MMv3EWLocFfB1SawP2x+fF2zXIqqNjU3
FCXLS/aJUsm2qsNANkYs+sgRaO1yoTPJnSnpVKLFzXKzugPbQXm9dU4itvNCoBTv
Tqc72mmpVQqwD807ZDKGkxGLvxJ74vFqnrLou9J2MW6CZ9KMinKU2kCihycvqSGf
XSN2khxPumD9XdNWUiMHFbYy8caePKhlP8IjnaOQo7054mBmhWrtzsPFzVWdFnUk
UxTcc++wgRU9PJObYgAas382M1TmOynKTn0MjJ2S127t5kt+ddzsUwBnx1uQDZMu
BYX/4PLrlMAGYBueQaDDbpOf2bERE0ciHbAtDylejNgTn+xFyxVy29XZKROtGrj2
069RsvFCJnLu7SG/WjQlkfVMFZ+FSXxk9J1vI/wd+//7FYlwf0/+6uckww5cidCc
qsmDJcRXVgKuaJz1bTrOuUSayVnNR7OAQSnoUwKUV+UCEOEnbA1Se6B0H2B9RDwb
x9PqL2eeH9ty4HYwosLzuL+/1BSWX+oWBvKPeDd5hqooK/JpzbCM9gih1LvTQkmC
Sh0VXK+3ARXK4VIBNYuTFthKFGNiH3/nTCmnsG1svrDNB7t1DC3RLMq0jCmlMBNM
wJcGHtrAe5+PDG96gvn2YTKegKcg3Or49zcZO3LAGRQXbV2kvqO3EY+/kPCcDIPP
LugAoG2H9FXmORViS3AZE7cibzisxcMxJ7lYAl8iCDTotg4bIEjYMMMP7s5MjCly
BKLWsnNg4yj6kkM85L++njv8diEu34EVIDzh7Hj0SmnMtcVkHftV3/shEBc3QHIt
N8sKO2AB9KV9P3guSHz9HaY9aH+RDhOev08Oh8i0ydlSjfHEjV3V++sz99g0c1Dl
/WZ/UGKPcQHGRU8ccJXL4hb8sT1kfywcnk2ZYAFY5ELgU0rH5Fxs+gvKYwYwZi0m
T/NVqpfqBPJ4ejDm7MXvv3NXHKDmfV8yEtw1MAcXSI3IzbciqyWVo6/KndBPWNgX
ccIaeJnrAxODZfnIZdYBpmdZFljgi+kAAgWBwt+IMwYEVFloJqxF5Dly2UlrJjdC
CMYy0rbF1K8jTIR7dNOu69bUaQS47oSX3ZW9V88dXszouQnOtJa6Zuf97SKO2VZl
smSEiI6NvYyvzaSyvzRyQKzYepaJGMlSHZyG5CLG1FAkZN6Exl6kGuxb+Cek3PCq
DQuODe2ol6aLJ+4DruLtvF1QjVtQBRrz5JBeYx/sGu251XYLFoRALlH7R7Yz7jDZ
/E2aGoJmLYoqs1dXHKW5FCXwII7iyHdAXvsoYZu+bsAxRG3/WIZ+9JK4ftDcdldC
0ldETjZ9yrdcTimAUPYlkw==
`protect END_PROTECTED
