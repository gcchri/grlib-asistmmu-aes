`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aWR2wZ4nK+SSFjTfc2Hvrs24THO7k6e0gv7ndqoXy/BCx9HSCVHHUn8ATLQPHZId
8O+8619MiKw5UgV0/VJOz3YOtD2fBNNkyb71e4aMFYfGsq/0FePX/lOBCigI0hs/
FeZWiXazsw4soL/M3NU4MyiJ+QgStmws5EmbsXnPbBqaeX9hWn61yZPa9NNQekO0
rqVKrPHbwVssvwqg/tZ7OPdFk0K2EvnFc2R2yye9yMz4UJbvcJ3DU6MTR5Dt4THO
u6uhCVq3260yXznWGzEUOrWOaW/OfL08fd/OnxX1DqwNDhDw8aDL3ScXoozaLMeX
b5ZwAHyOiZjeRfCwugXb4rINXPEin+KZqWS5mVVPIYhjdqOtwxsWD+LgSf23UkGz
i2yCO/rczCX1bPcSbSo1FO71p3Z14zWWPy4le1ZoFqU=
`protect END_PROTECTED
