`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kKg+pw1mQYhBGDqfm1nREqpiMpH6etDFBS08kaxwur8Q93EmgTgh6cdRbq7grXpW
LCq4rYHwmpSRWr6IzXTZii990pnYmjCaM1Ri1/8EulWFs4HgX4fJOqdHarUzoW8u
lAW7fao+NY78QcwFcRGlSFQmESm11dr/MmIZM026abv45A8n7SjUPZPVrc3+Xb3L
qPcjnR2Rr+lZr2zAPsQBKNG4b+WQQKGDJUb6CC2DngG2rNkMSNqgRZdrLv949yxe
ywcETv+GtFLiQE/VwRoVKtN0y1clezGXkxGyAleo55XNAyjhENxtL0fa8X78aXvD
eurvkt3AvI494AaM9TyM4Tv1oyTIsVsl9lKqCo2e8yBn2FD1ILLG7zWWvbX4+4sG
`protect END_PROTECTED
