`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fNoOmi6c5XFZVqZasOnw5p/uetyXkKhOJbmE4YZpfMwiu+1OLrvnStJAZ51FMyPz
9dC+7bKBGSAxIINaw2up2kx2dRsArOY0D70W1XxetGm8+Q0qlu61tnQdzhZzauoC
2it/OiTHy5vZALgPtC2CZVDPAOD3rebCN/67939+nczNSdTSDMeIcsB4udLpznCX
aFoNLtE4PAr/VDiiP5m2x75wCTkFdXUYfuzfAu0a0I80zH+P0Ipgh/0eD6vhS43G
HpXWpCGMjiPEVTjFMPAC2ltgkD9lBhnwv2mA37w11K/gpy4KEhPmhrUGO4bMqI69
OgumIfdfLKc2q3+ihFovGOlyvPuyUfT/tw/0/7hlvZw5PnuG2a+7jMjH36edsxk3
ZczfoQd76UbvwYyIVCFOGthrOhXzPeNieYgOx91HY4i1KLNhQgfqcEbJq1OBAG4N
V1CfXliQnwwVJcX0dGZga9fAV682Dy446SGSppAu9RjIv1io5sonkYnXOAs7g3Fj
`protect END_PROTECTED
