`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pm+aS/cl+n7HOXgpSqx9lp5IiCkCS/yJHiIXTCPAaKqMof/Ukkey+9w8lVL13/zv
4Drp5UuCnb3pXR8vcn6SPHEexOvuyjEslZT6dDUxlbijh+7ftvA2FWeVUB7tjw9t
7QIYuIZGchnUrxG13B0zWngdJEgAh90TQr6144BawJ3CcDRLFZW07/lyfi9gZRDo
vLXflCOtEikei1Q749kdlKgQwbcHN+8bR8LEM/EfOvyd8lGbrsuskvjC0tli78Da
FnUA+EYS8qqHGP2z5u5v6va7ZjULaxP5eP+gf3zJywa1EKv9y/jNZsz1/Hte4MWu
VStUlj5nyk/noArpa//2I057dCBIcLNOraxUJdkpmGd1IWlxF5Hc1tFwITL4a7S2
ov+uazXJ6pf0YRLLGDY7yNTloyor4AuFrYiZPeAPEGE=
`protect END_PROTECTED
