`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KEvDe824b5Wr8uyDnEtxMKGbBVecMcm/xldTvdmdmTZlZhJAeZ7KsW9XN1mxuY5g
RNWknWOZjrSc6AdfADyyjucRVcvLSFoU+Oq/6SgRo3CGZr1VutTuiNps8zBy0uUd
AGq5N+YgVH0cvT3SbW3HLU6RMyRPdXbskX+Tt/qZ9Bicm9dEeYdq7sXhYQn4S7Oe
Eny0McLzEnxl/VL2DjbYCUnWhx/DRqdpUUAsJ6gQ8aHNZIeCOa0jfM+4K47LOe9U
Q1uRHk9JfUavAUyCT5pUuL3Kz2cq/4Lg926pj7fcUqNrSeXIumo1S81aLDswJj+P
oOb9upRB9bcCrol2A4WxdviaGt4YxUrF912G/yBvjiTynX1kFSBWs2/VRjzrfJGl
NHP48ykEbIcAttI0Q8FBSQ==
`protect END_PROTECTED
