`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w6quZ/uuXkAeqtiR3cSgJFLMnLppJccbygvwRQRcmWvE78wCFZJtBc7ZgZnlv5e9
FVhGjiQgXtHb0LdSd/XA4NZmHmDBj8rESnZfZjzNHqSAGWX0JgHW1hD/foULrN+k
yELL8MFkOZnpvOz84RSBdgPMfsxHWE3JzCJMMO0S6K4wQ9StXEiy9Qo1UnlBHrSD
PqVXIXtKPHEbVmQFs5st2ROcBdC0V5s10YF7oFkUtbiB61H2nh+D9T7xqpRbQnV+
ZLWO8AL6KC7ckjwpFu/rT5tuOLXaCh9YUkJh6W9judnBNGzkJvslfou9EMrPB+/4
WECfm80qMPaYg1KwMjXgPBh6Cuz0dxGjFMBUuADqf57jCcfb8wuMA0wnhCUP5vXs
FB7a3NSDxuizNiC7Qtga0MJoWbQgdrI/RQ+3J4pi3kWREUr2Z7256Z4Cg8gWKa1/
ESa6gXrq/H5twWLcPS20zlAO25BW5Cuar+vw20b5KK2BRAM0cV301s9vZA2b3MQH
ZXKnVc7V6ujJxXCrluePFCTk65f0pLko0yB3mTEROu5R7u9CH+0u/2mvD2L5PtB3
aP5mTrmOvoiLemROAdm5X03Fz8hZ/SmmaGARXDzphD40kE+LtI4cURIe5nOKNYgL
x1873sEs6DuPvUuwTFppIA==
`protect END_PROTECTED
