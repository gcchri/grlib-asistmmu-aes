`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MUiXQIlR33Y151X97++u35Bg72C2+TG+xvkG4XeSFXk7kwUIfA4Uw8PEu8UL02Qj
DAGFTkAT4YmQnQCLc1PDpUPpGTRGvDd6d8bjT71Y4RONJ7H7D1XVU5jYvXUUIWR3
VLXGeFstHYYbCsURE2nH1P8v5kb7i0zW67rAlt8xrM7hwNBZaKooApWoZnAuClu1
heWL3vM/EjfuxrbNLM9uxLF9AOtYSLGgyLUYeIaSR/maHQDhGqEADF/4mnMQfy9f
upT2OvWqLrCOCjjbB4HMgdFpXsC++l8+lle15G6fJfg3+ednZaTkRItpYF/Th2gv
ZkeZ4eDNdfoUCFa8fPWuE4y4e83ApHWVKK+JpUCC+IhtvGnpOG431P30B/vPVmo/
e7f3IQea4JMsTmPRN5YO8Q+NMK5Nwot3zfBnhSt/9/03rGJxxiKmUKdv3aU3Xkjv
+PdVUDckd7ebdEFniMVYPkREDzExlFqCheFMY+jyAtQ=
`protect END_PROTECTED
