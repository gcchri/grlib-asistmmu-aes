`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DNkrX0dma/jwrB99ePz1TDm2a2lhH+0OPQk4zZw3XsEfTR9g0arxLnHZbFwWQ0Lg
uGOp8div3AebE3eGp1QEBq6X08Ay5AF0b/QmFMMDTAjreAndLksigU0t0cuzDIHL
WpiCxVmbBBhaALzvN72BoeMEsxRh4JL9ay7H9xzyGQNKQ8hqrRYqRMYrESbQpKgB
UXmEbnSRo/d756bKOXJbvFb1pQ3CBGQofdCivNImA9maqtw56ObpB5IRdjpQk8Kv
BFuZEnfBmSunrTXEg/3LoKM0BhNDnxuDcJyRsNFVKbe6aRYIi5EF91nNn9CDADaa
zkY7xp6QLDu4O6ilzdRiqfEIej1lP9idZGeMEIsrdCMCOtzlzeb8GZLt/kIfXu4h
/M56wWKoJ92vmmercEAT7M8UMkkeFQTSk1bwxeAIm52Bez9tPwD3Gaa3mjP60C0m
6r96B99lvHHnalJFyn3A3kLwJ8oDZQ7rS3ec0F73XJXPuO7fi8Fs6G3/NrD7DKeT
P5GKxsy/9hrdhDwDXhpHLOtegslIzeOWZTnNs8YOoL+G32x84OsMlanI5fcvec9o
uDUpLxWYIrMqHmrZteUkew==
`protect END_PROTECTED
