`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U56+r5AWy2Nw8HeIK9XHDtWlSC6TFCFaYPPB1Ddb52ZUCKrS/gRxRGdpXdYUWR3M
CY3NroZ5NxV6zNCjd4OaMCSIejI2lvUPAtuRuztK6XoJZLDjYhY8sxl0NnMiFux0
lK55jrLG0dfF//+ob1rBg31ubYQ0cSUd6zhj8rWxeLvQARrNebyfS9qGj0Rdjix2
obc8URhl27lXq7dGa5uOJY0Wu68VT0eE9YrNPqa9IW2BCLjS2OezjbJ4VMUwZh8r
flOUaP9oEwCQD/oOUwrhsOUzQ3XTpwKX2XID1o200j3pNKuZT7deSNRzpl9xXspM
6ktH2owzC9Z5Sg8TzHjLodDQApHV0+HZmQkcRwfYljOiM/PcBlYMtZ6F+NyqxWOn
dTB8UW3cuUcHf+fOAqDTDj6gDuL+pbDdVuzRc5W1mZxwu4JS4jK0EgsYhNpbFEKu
2tfntYq+RRikCiQ9dPs+kQ==
`protect END_PROTECTED
