`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f2IERl1N387EMVFhvhCjyoCKkEpMWqd6C715qW49/Mckxb9+taLlMiTiAnttG7vu
6lr/K3uLm1nx64GdI3Po2wuHT8kE4zw605+3SuyXibD84+ZkneFSjnU82XJI53o0
tE7P8LcnQ7cNOlZy9VmQDmJwYgrgmN4ZflRH+X31BK6RnFHMsyfeVrmEXIfRYNJG
nlHt1R3UTfWNik/izkhL1T9636zdREysFTw+N/27RMNuQVgWW7EnabTqbDETcd8m
hPKEzpj7HO2NlHwpUU6LXRSix8V0uN8HXx97C+lS3lX6lCP5q7DIRUfncV7EsArE
RAAaS0ebbY62CTv4MFO/n/CpRX4pYrJFxLN7fwHcrZMPDHgQQjHGvkMUEnk7ZPx6
doMS3gCWdsdpolXnX7hBWBw2PJrxlGzBm1zVbc71NZc=
`protect END_PROTECTED
