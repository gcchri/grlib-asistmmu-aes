`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/faGYfDopmnaGO6oTiGrZmBfsTiOpaR8pdihcNMt50tVF28HMECsmhaooc3Hrdof
F988rRXgCkEKYa5EuY1OA7bGxJcrzUZ5fSx6qHmdgC+x1Y8Js9hVtkjiZe0qvVqo
NoM3tLZ2Bp0aCVGobWC5eF95SdjkAWyJ9XgEaKKCE9F6arcAUVZbl8rfNnaBqkVE
vK3O+AHRk1qOax2me7E7+xHGZJgfAMjeTyGtnMz3ynELaD2RSMm0yJqLt+VlBs5o
maET/C22RrcIghIgyU+GJuolh+6g+ZGiOfmsawLAIdLVZn119lpYI6kGFUjcDfmY
z9FTy18yrPNAxIB9hpuY7LiidsCGt3eNoWCwmV+lJMU=
`protect END_PROTECTED
