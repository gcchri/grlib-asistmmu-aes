`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
biSpCBvnllqlTYvh08PSv8/OCA2hFKCJGAV0iGBEgkhN3PYF7RqHTfPe6ntuLrzb
lzCqeuk/qA2fdCD6gNXvkIKlTPNlR0rQYW2T3Vy7M43MgP+xFy+fbGkAqk7p7e+Y
ERz/N0sdD1iV5Tg6/GFr54vIqa7OIeFH7I9/ZYe/Z7JudJofnQ4Jr2Az7CXN1nRG
9oWAO0Vq9iGFuQ/se/VuN67Vemltqj/C51JZt/XQ0yqa/QToGmNv08AXQQ6oNW+O
/YUifhvk1GW/1BnYVVHUaiej5euEQoSy+Me5NBOhDBMF5pVYmtX8CDQXbGwp+6FR
I2+xQgkiI1jrbDRN2D1ToKS9zCJvhEIE+0PDYBSPn5KEsPR/U+6fnLjpgeIgOGaC
txYyJ1tos7y3dJ+6M4YabugO9iwoEdPzIECn2bTyxBMjhzbT9Wg5OGyf28jYJUNF
pSiCeyWfKf66pgKWRxoxrrZQEgpxAAJ1YWpGbpBdN1pIkfyAIXOYAd4q6BFT8y+O
ieOPup625brntHwSQ0WJsoqkZNxh0bQeJWEnQ63w6AaqMEFPp1KB1mjcwYy++S2j
SnETts13Lz6Tr9KjKiCd0UFsQYZ0gTqcZ8qyQI5CsPags4bexldC354Tu6KIzsWL
qCN5OtqTZNdLVZ4khhUGT0yTzWbKShKHp3/SxAVaDcnZrX8M7hD/LsIgEr1hVoOC
a9X5FIks1NFEQF/41/3vNoP87HCIhzRo1sE+6Yy5ru4ruwDsHcCU0BKdtb2XaGFk
iTTHxjT2Kq+hSsyjm/ZW4OqQ2NcU7QR8sQuloibK0qfGYzMsCw6xXmHdmdq5+J1P
9OknwJslRHgHNY/qMscPhk1xgunZYrUYLtHf0OZzdCSTzT7WfUOyJ6N03B7hM3In
b7wilR2/R1vPwr9JCHjj07eiDNSRzkJJ30t3scTWcXWkx0HBY2MRg82sVdDhmuf9
byZVS3xQ+8b9P84fsHPbmh/sg8vyeuFYCqFHZNC44keJvxHs3+QIdaF2WyRdPBSS
oYfYg55RNwurIJ+Buy1V28plYc+d8TxlRKuJcFiG/2ZqfD6CTOfbVsNPPtHDqaKN
Xp6YL4o07jrUZpMGcRxKhzazhQUeEEppFYZ5J/NoYlv+r5twaAGZSqMzwGzQKr9y
/oaQcH73+CNoyvyldOCR7qouZ0CEJOOcdenI9T8MzMQAiCK0L+lvssmo4hPgn7+p
xwxZ1u7EjAeDwjEF0dtltsPe8kd9l0KP5Va4GC4lIk4fAMFaAx/Rp/qus+EdN4GV
lkSN36Ic3tUK41fEhVgtYbrXvQN6YuFYzIXTaTPtdV3GbQVw/ZOTbhZKohFYLpJM
zJ2HeGWSWzH9EhGOetq8N7bsMiTOZ/pBLkg0EJ4HPCaH0Il9A6jx3L9BKRdltYFS
ZTZjhc0Sv7l18ygXDYh6GBuTcB3QylVi+UaJE1NrpvYwDAJs4Ceb/BK0rMwGl4cA
kpq4pM03AsMLFMArBwdhEqGS6UMDF0zDw3R2y95LmH5VQ2fbUcKVaIi34VBBqpCE
pHqSSNCTx9FNW7L7j7u6EwS7UDmXcciquu54GYozLVuVmMraUQdljUdxaIXxenk/
rfNE3wex3QJvcQ8bZ9955RzsxV1Oz+GSJVfMkS6KjHhd+YHXM4dJNZsrpqsOSqDv
1/Vh7tMNZkNsYtCifzhuOtWt9iIEEw0Yidiw6GK8IW1kcRyb3FqQfZ6pzqYbm3Ve
LypBh/uWPCvPyA0zjUQa675WMujp5stsqnV/7FR0vtsi+P9Z6hx9I98C1gTX3DHF
KRpdh8Su3gBhQX82JFCG0VY1Drjc48sUF24RliPYY6nEjN/9QxIDTWsNnLFL5YAz
SrnZNhW3yaKuhSzsXpD4Zj+7Pg9PIPs13BpxdePtcXoBaVV6R8S4S3Q1avYzpE9t
Uj0lcazCZjGtYZmFplMbgjvT0AHUT3MV9V10nNtsZpibP4pSvtWpb9KRLs0in2t1
Ybucc6Qy796bZk9ryIMuYNNpJ7ibNhuOr1g3hQgAvKwucQ543xGhiBuyivsaAX7N
k3jdoqDCm5YYyMghunnWyoBZq44DiZwmGwL5nvqcDsFAVQpNT/cgwxi6xevFbfjW
PbdQYYCCVZdBXiYn3JP5HY5TB/L0hGDy1XHhxuxvSZu9Mz6bunArfXLkWJH8HxIj
WKciVjTYrbq4pGsFH1QmfAc5W4yCbEwpetOW0XLjUMGHPqZlOJqwXpDgT88Qf4l0
6scT+pQKgJyygbvJnoGjT0pwI1W4QUmx+ZlA9lC7LVBrYPeW9lItQlo5v//GyYf6
ppuRnNEZe9zt6cEdyW4o6NS93T6qdAGwlY0KEGVW6+S62LKT+cVuqXLMgWWgnM5y
IIIRP6V29DTaCorP6svqm10xS8pVhfAhQ61qa6FuUq+Gvfy8AbgcYKhEpUSljJ1V
ewZn0kjiQwGQ/P1D6XGAjf0s+dKIz3H255AZLyEnMm1PkKh1FaWkHr7eEPGXuZyO
XM/YhqMfEOZjRp3ibBFFQmXrN6XeeIk+5O6uVxQMPUnNgB5z7OkPynXsLDksV1K+
D5Sj3kuJCxV3U3/ZqSRaWMUucvkgx6rfbWkQ0wrDTy7gqTFyd/cBaw+4SmOkRzn+
Za/nm2D1Czui7j37rJbWcuzdF2KBDj28hhltKhYzXNrWEhyY+D2jDUY/zSmFqaXd
+afheNJfe5q4j091xm2V4egsCJARL34tB4a2I9HEvjdyrf+nwda0ps29vVTYLkKJ
KLERMFuMjD5SFGG3uKlom7riC70/QGqpxLvjm9d7glDnKmQm6fXG1GXYI1msWjvw
Wug5LUD1wjpH+vpu2TK4ZM1ICs9RYQss3IJmxNRtU/SwzKEoLsR79Oq28VylvstX
ERWd5UYezJ4sAkUa9h7W0/F4+phuw65zV+yq0sRVDdIRfLs9N214K336+KdYm5G2
3espOW9l+JrWD3R49O9jE+iMO2e7u6vk2KofvEvCQNvrUSLvf0NIobVv6soV9TUt
bL3J7A17k0pHZtqIGUPp2+I6Km5/TzSV9NBIISgL5NgFw7d0xymlTh2X8b8Oat9k
OPkjoRVHb7nur24mRpBYL9Y9yzK23bOJRvdgaG+4s2VN7zBaGrEqyCCN2ra+zQLK
IwD2vdshYZZ2Du5/ExsCFjL+6K7rdu8YHX+00SF02r93xxPJQZ81PLQlybH45giW
xWoHC7WEf8dcn/P1pul14tfNzIywdhBixOf1dklD4S/60TXfZ211lH4jO1B0wknX
Z0WJxowrVYITOHC2hKNZCypHIi4v6nBIPnn0Ap6TpmQLrghm09m8o1iz14XEwMYL
BMhCg1rx0nTcvCyuc1KxmY5u3ZGBIXQtNJflDOOGrznxrs0IBAOVWshhg/i3U4N4
YJsRERk/SsJlKuFZwQIGe3DCTBIDQw+GL7Jiq5Bf4kmHm6HXqmawYQov3wVTO/W1
R4EI3mcRh+nAQCpEa6O/iXL2Pi5/bCI1/CE4jGUZJLyHqXUVZ8LDh1FD7F8k6YIY
1bZ+d/LKSwJt8+0H2zm3KJ8CLGD+g8iRFx/86/ppalRn0ftPTck+Yf8l9RYmfqNX
6j4D+B385sr+//QsCNm+ZsCXgQAAA0GbjZT1pEAkt6+PqcypktUBBHQC7UmS6Lks
smaSBt4j+5qCmFW3OPS/MUpa38DIg6qvPNCKC97aCTtKmiBBXyuVPwqt/fy87LBI
zeEWyDYDH8kXQ5YmFE/pdyd0A2kpX43P0kerbP1KH7sOEU1+TvbY6of1u4SEFoxn
JTbHtdxWGxTIrJPwBVrJX/BQ4ry6tYQkqOll/hKP0Bx9kZNyr1tkePh8Kftr8jwW
RW64lYMooAMPbBKxPjPkH2vgLP85NTmrytMnQxczvrVrIBJyBokYTgaExmWGy0p6
xAb8cMu2P0VQz2J1n8WWWi16G5j4zOFaSgOqgoAKpOkGYkk5KYLma/W6RS1CPkL4
A4KSNXLfHuyjC522LfybMbtY8CYOSSP1wDO14cG265z9WUECUW9cE2KXrRfgjs8M
5jkHlyurNV8P8RgOetORqCcarPJ/teeRNzzlk1qj1YXNLIYct11pPDGNyM3GvX+q
ssBqx6x4JS63FCMHkREnKCqrqArRbXUi9rXIizXsSyOsizKb8eM0Hzl3IIupf2v4
+S5gSIIJksaS+963uWbQoDW7pdK02Gk29upibECNweVB4h7wYd0Pof2uGOq5/m4M
IlSeYrUlHmfkRbOC8iJuzDHPLeCXmf639mTejJmyY2XSsNdVFBEGM1U9dqhJemon
K89cJwW8TPHqk0kJByO8BADJJ2BoVwORu6ZP+2k7E8g0yLj39TMpLf7Ug8x5c+bH
zgxrnGDzRKeB89iVAfG35CrWh/naW5UeT3n97Zqp3Y3ZM0n9r77Blc5pil7niWjx
S/5m63YLfXAiQNGPhV+KnFryQWE8+XNpCibqxWN2hTaFDzVZSJ5+jnhPNq3Z0AAv
A+mAuFT/0KAMSOBGLEE9slZsa5uJbEfHSqjzDhd7UITQFl/pBM1TVOnx/niNSDqn
j95DLMRPwDYy07MgeLtOpOnq3lzerUWZJT4PGvDRrwU+0Mta//Duq+4dWUJpsR9Z
DOd3jLAb5ZFzZ/gUX3vB3w1f8COGcVcDtg1CxDmVaz/iDo05ft0KIQJ11XyfIVYu
yq1gXipfIxwXfigKNUhGSqDDFqQLyufZ6vmzwsXx3Sa0kalEBgkH2GkrOq6docoh
oLIEK/Qex+GmJDc8t0UrJv2YcIRTzXMpGG4bQ6VsQZ9ebeprm88us0YBZcv8CEmT
Jb/zXbyoXkXQCWcMm0eogcRpl5c/O83EFndS9kMpggo+AtApQiRh/bZF9MLHNfkF
5YzunJCpBIkQ9/ZCF5Yf4xKcb47fNidEKLs64ThAlWfxABpeZRnNk8k2PHYu9Bzx
n5qFYzVgq+TcD6mXozvuk8JrTPOQXivki+nGjlXkqEjEyJjvPq/jT2S03POG5f5d
XjPAyVEeCphY5yo2tOSOrARN8h74ttcVU1eedXtlz3Lg5lI/tIbKy91bOoEpOq8p
XMpASb1PBUnn6h+f3hCAFjjoAw0zETO5Ewj15EK7pKPMmxb7EeWLt72uWXilMJQK
IXvy+JZwwyt2BL3OlfLt6RYD0nsv8Dgt7k+T7A48OlCKv7zb8tOsUzt+4nGAZsMN
NVNjDkF2jITbUfeCBN/VIZSvTNJE/9GGjT1fXNlDkyzGI21TsuUHpvy245M3klJ2
u5i1wh+lIj+CTY33x7U9CK/5b/5ebpJp//moP05K4d+Kdx5g6hIFj/iSjpQGb/GU
InRN7MoXaTZHgLpQwsVlm4y9mofq1tC52meFcWIjPMSUFwaKLOxeg9BTBfU7NYWF
q6dwc1r7LvA6c85y8Hkb4+O+gf7GHnujLIxMpgBxVxJNgRkozx52AjgWFaMZVe58
yQyLj2GJqizgAmkQWEvS8Nayqh11485uST04jcy+viv2+l2Arhoj29iXyh/mM4i0
jbhMissb0YB7yaBfhVFSmJitd8Dh8aXqoO6bAwqA5yV1XZZSez20Ix/rgxR1TdI2
fQuSrcVK8pM9khbZmDk8Xdb8LuBi77gr6a3SJLcpEPB7tyQBWN2Jr32lRbFFjze2
vetWICXMNXZrh0lD63LmnVGmOGVXM9aKCVwnZy8f9WUJqN63iYgH2TgWlkEsKixr
KWlnE+IyDUEn81ZaNzkm0EYoyMbUykyW5dEUyQlOUjZ6SNw0ALXQqRC9uTXrorFQ
r33bqGermf2NXXxKqGxpcslZrBUZ5skhBdrIzH+SAh7QNJ6Zh6oWT28yJfbDegzE
LZ4WqK4p4ua88iTZWFipyxh2jkzs0XBGdsTomfVB9xBZKTTIj4tZ312REAdICSxH
1jHotcvNMLJhvmdJuy4oTHWCpiJbH1qhGH4LpCskXn4Q2rTq7t9cxvbgZTIqJKG2
lPDAZvID3U3WDOnudYByjPOCeJBQDU7GvBeYbdPqoQM0be5DjewkyZ5C/JA3rCB2
zKUSJx/Ile010aW6Gsfg5r7y7Be0gdBJSIvL1u8JLnvv4M0jxpMLjO6BbMDIc7AH
SmDDO/31PCHRCvzbaid7397DnP1U7sO604mq86ex+kq2GHglOXkbs2dUN4AFlHqE
wCSCfjfe9iWavOHvPZRJ41nmo2g2zGR+keh7V9CSIkuGjUeu22c3+yeMG/wPxE9L
mtIRI6+b0jMmdTONhcAEIuSz0yZLF8LodxIJWdZ2sKLhUTh9dvl3jyquET6y0GK3
EtqqYdFhfUgKe0/+H5RDYoOjTG2/aqB+5nh5FKK1NP/bCZdqXzUzAm0i4XD6svSJ
hnWW7v4gaGv9oYzCcMIVs2IcNTmSwMesGZcH9+N2MOBoESnjjnvuFSXNEVYu6hci
D5shz/l34p9THNq4YjGh4zM6HQoRAEyW4c9lZfz56uZEHxwn54itJUF+eD8GoIVP
1787nZobQBb2Y6Hwh7t66/a9dsnt7b+9ylI0FLZObxCiKXojLvwEAeIbZDt9RJDa
Imy01vOeYfDQmPrVF0R4SNTd51ypCmC1Nb2wpWteJWHUrTPhBemhiefUO5EA3DH1
bRr0VVBR/Orq4A3hZpbVh4fGyHuvet9Tz7RZwEXxdodJIK1ryOlscRUFJgNEadZ5
cxT7lKoI9Kem/ATUus924XXfnSfy+BLvrRVoPQ7IKr6i1SkLSnpgW87fGXbLSnog
YH5ZAZrAByI3irKZafnF21Hilc2oFqk52iYEG4oS32M6aGpcVUAqLsfyq6IZmeur
YWggHnfepfwlTO171u/W/s0Dw+DheoY8gUozfcckNctywfFO0UCpdp6BYXnjDRHS
q/rIGRU0x56q4j2NlsZC966umNvDJfmlxPe3FtLaB7xg7XVOH3R50aL8IjkFjJwl
MiL+ggmIZSE61qsnfQmA2DEme99tPzRm4c7VevwIXwzvjAkWRIYGXtwqC0OEcvTD
OVcaR9g3vd/F2rxu3tlsWS+aQ3bTvlcOfB7t3Qvkdz3A0QB3CHQplHveqhh4Gt90
TfOh6/i+Ea3LVucPyZoHcEY9NEfkOVhFJQmgkBLoz7wuAyZSXRk+5LwrqzmVMmTN
rz0F6IzzkTmFd491fLp3UVQM66olL0VEqrhIdnmTOfQzVW59O0hayGuL/mJiPq/F
FyRC8GB94rhfv91HQPmESZ94RRSXrp+EpaHMfljCL4deJQU+WreMrhu+GQbHzx63
SviOgl2nZ8TjNJxvIl6Ejk0AIJc/08qGAAhnKTZlNV3+glgO7wd9xoffzvYCWRO8
RlRakr9dWq0RG0Hyedw0TFEj4i4F55k2r6uc72njjxI6LneNu0XAVi7jqlayJXSe
lISlI5g+B2ZKR5C8jW1ekkmXnk3/l9gnKyeGCe8Yha0PYDAWLcVRGzDlrh8a0v7h
1Wqq9zaGACbL4PemSev8ZEOV0oJ+Za3sOa/Vld//wbrTBHGfbF9lBl/1QYYnJq7Q
kemiD1NU0DfC727c3D9bZiDQWaJL2244rfm/pTC62di+tJEOZnwyYtXkvAs0oWb1
YB6H8Xj+3eRJA+vQCmX6s9tHhKPBJSLHyfHdKS5bZYdCnJrniUbAIxEZYzExdf8c
0pXCr6lrkgSF5dCArZueA3Div0p1MMujW2HsWwGg4yOEQXBW/RN7LYYWOQT0Sf2Q
QAOL13KdN7UVbyKqSb2J29gnb0yp3qwDX5vH5/c+/m4omk4KpUM2rsoicgfyn0Og
P4GjU+9T3RKXXY6eBeWzMqX1v+/Gdr9hhsZjIxytJtLFE4beZzw2tkfmw07WI6Eb
d1J1JZ9dDVT5KoednfsI41+x3QL0i6y0ewKs/cQid63UV/TzEeDkGojkN6Kl50DQ
0DF6/dTY1JfrdInvbfU42BxIMMg1VFJpp/jNnFl8+DeeNej4oRCMxsmt/bXD5Rum
TGJmMQAd91B9fIs+HOFss/qcSh+ldVRskRJtBzbrJLFZsw1gJgOVefMqP1SOc+rk
BUm9AIQhLhTwcZAQU7LorIS1bHAuun6IQp9lOBJLODQJjTlTMb5HnU54CdGFJSBK
hFFp52mqPtRDZExjjYKnTIw9RJdhiRg9Yn1KO/8i0URKC6Jg/3jrXbNQX5XDJKgR
zb/C7jDS9b6U2IzvxgQV0xKkaYsvrTlUU1VYD5z0swBHCPViHxY21HliXGvQFtXg
ypOuBObOJnypivvgOZ2O0FTM4PKWx4b0rYvpzGx6e2EanQmqtKsQb+muNou5etJA
RZBBb/do4WXR2tHK3cZVQZxqLWMjMnWR99JOxlDxuzShzL6eL9MEI2yeXMpDzebi
bEIkQ2/dbbGmp3rJb4PKronjc2NResxi9Y4QvzhB5RtufNcwuRX/2URB1+PEdc3V
v9rlVUh2x7xdI9CZsHAI/1ut+G0RdfkYlP/G1RfPdLCSAKtvpEK4bbyyvgKt6t7d
VNB4UC7RrY5yGP0gXuzxRqHs/TUB6PkrDxlQ69AE0g5Sn1CzfHI8aEP9BqGC3X8o
6oaMU4w8gHUaBQMJmW/oqe56L3TWhnw8o9Z61xQKJj0+Kq1UOV7T7MV9UFqphv3H
nUKnLHdYguwiz/or4aNjrnaIE4JgqiG8CCvxXoWnluOkRYb8iSvorldg7BCJNgZJ
00PS6sPck/ragX9Z3PFMA/RUKH2QwrTZ5j6aHHAvTX9vyZZC8nscYl0USUFp/EOL
zhRXOvgSDd9N5P/aF+bMT56plWv2LzqLHrdL8xwg4KrQwZUby/purg+0QXgb4gNI
HAcaKBtCZX0v7uqQVYlQzFPLJyVuEETguTVqeq4T7G5PW47BoXWQ8hZtfRZjlC75
wr9kYtCuq8ujRFin+MOHR4NKF1XKGx0HRgVieN7f4iDpkrEPZKnpu8y9L5rQmm8U
vanP0s7SwEX4cLbornql2MZbde0olcAt7hpPBsAP4nkL7ZGT2YF8X9dr5hddfftL
oZ9an5iYJkTKXQUmoiXPnbRGL512AmN+4PE+mEVglfmlq3BAVFkQ8YlBeNwN12DJ
29f0Q2P6Z81IFD4gjbldepe7AUEhVDuESpG9mG8RxR+3h+kDwBQ7alRfbCIOkxn+
NpZ9qpz18EmyysKEjjet6GL0/PRy0olaSHmAkHXXaBf3vq7OKmLlyI24C96H+bb/
qJuecmv6rSRAXJAivXoHg6E5Lzi5sc5wpwkLyT6zxDQ/dYZnapBuUP2e3Xd2DSn/
CfJSgel46MtODpLItFnMoOStLaKDicScoAWWr/GhBDnqpVtAbNqRf4RpckEW7iUl
NSF2RUMAYtSoFGlwSdd1NaVozv/aaQLx/kgYFR+6YVh8YMCWp8L9YhuGHDoKq+yb
+2Bl0m6YIxyTWZT3nokoCxuNYhBNplKTnol604ODaIiug5htYe/31J+4YRHhK4k0
XyaltqdAtk0QRH1vCCUWuFotePgtrRNN9DiJGnz6ZmKs0+YSj26+eqN29J+4L/l6
sOYLgprYM4A4jQEcTNL7VEn7IyRALuTzznKJeH6cEE3VW8WPNe5Jgv5hTYUcK6/P
BURumuML34OZouYTNK7c1xojWamXZyjqsw4/GB0B9JZlFW9JS1UHZsadl92jzj+N
ReFa3tOl5n8CVQNqkK9I8PARKF8kDaPd38GXcKNEgWSAxtjibZ7L1i+RX8Md/5Nh
BZkJct1KP8OaDH76JdG2jTyQvIhDq5pHzWTrxVOSW9bg7kJp7smqYWxancRVJ5FY
jHZAjwVl/t+2JgahE4wXvZntQPb8wxdIMHH9wdkp8QNdhc3tjp11d/AlULdymtIO
DZgL7/6xqxwAWKiYB7n+z1roG5MR6VxPZeDyYIEMlgeGoqY/iRJTLu0f3cqK+88X
56/QbPVzrfyukUnxKx+GQpSPiuC8Ph/V3WhzEZyz5uWXk0HMNj0XVSY9Mtl3ybO3
Wg2tgQVAvmTizs1raTvT8+8xsZI+9aH7vRonmJZpozyStmVJoSZozUvePa6p3xTh
JR277+f7DL4NUYe5eWkXH6lJGV99BU1bJ4qJJBgPdzQgt3/pjTSeJvAWeH03pI/c
3KSYr4ISS2oZ3kLkso9bd+ni462fEK9KrvG72/niBV9NYQbOpFtHVGHe6IMRMNjS
g6iZWD8nQoGq6puQDQ/ql2Ph6Z7q+S/szyMxd0+unDtFYC5cqp1v97Nv8aJsEQMM
eqSa99oJ9k9QgOmb5b3Udd1NrryKIg3msKERDY07S3SdJTVWX2Rd5XMWAdIBno8F
dj+Zc46Fik/mr/WzLBdyD2z2gG3cqqQSSjFyqx+hvOcfTgKREUxEQIPjnfP2M8AQ
yRFQ6gNpTw36naciv27sPWPJnf/+Neh/X0iQ2frgPbAHbPk2DHsez/PHM4zyFQ/G
9BSCPn/0TFH87yNXYEcMzN/caqnlZPrwvZPQ4fIVIdS/0Vkh53hZ14dwQxCj2ZRh
11EJxOPVZzi4pmNhm0978sYJCk9QIr1yBr2pMXqoXWfY3ElpS+bOWF73JJVB+3rP
jQuZ0EhH5JHenV5feLtsNEk0SrAcwntYvoLaDuQ69FrfvX8Bh0ILBSVBBTVNUObu
5+D/sTIOKmz2K8dHyLiS8e23HWN+3O6rvCpszIQxocCe/qprBG8xeBQSIcrvKDSl
AIjz/3Y7ptGlCa/VDzLAwD/AAym1Wfs7VTqMgcMNKffPTAPonNI0QX7BqtAO8qDo
o22Odf0AgMIQQMB8MNTZ7oIn4ka0Ftj5mkpIFcib+5gkLuvqbiKThDjK1j9uNwjl
Bph/QUcXtanso4xUXEm4INnFSENRfbH0pzyO/VZWMGUPl+89tVa37W0ZwoI+BQwS
ttSQVZQbq7AdN53QGhsMb5pC+KIFOL2ufBHZzaj1o/PJpb6exRYCchn4ZXll0REu
MFvrInXQCdql4M7WJnM0T8x4T2gz1pW6Aa7wOl9I7D/+AN6nZHyFH48FLCy0r7dq
C4aw2nGxKNcYJ6wxpET5PQ9avvPYA48o+nEvsWUuV+0HZS7xFmVK5NX2XAa8c0V5
TaEOlEkI/NRyc7EiQyvFkpvNLVYFmXWxvUsjM9mFZkFBi1EgjNwZJFlaatyRCUgs
YY22T6EKWWF+K8FTolCd97pIJb/2UwoIkaIbimbKKP+LZoZly/510UKwoNewDshg
GHNXe5ZEoTug2zI6McFUxBGLmpCqPgcqY3R7SaFt8HuhvPgrCp6F4N0q0n3LZ1//
nUzwrKA0FUNxNwxY6MsoC63W2AltrtM9naHCz1JLfipCdrLjtu9WKWIL/O6VyE1u
6YCpSSrKaPSX99k+hxIII+wy1HY1cJyHPg75Gzyzq4WZVt6gtx/vwaSiZb2RIGV0
fD+rERYldGpCi0q7sPphYIqzmbDFLVQKZfSpWhMms2B9CMGDQcj3vWGyz7mdHOBY
eGMVGx5xFzTW6loFEiBnFKTBc5LfTXmP7QzCsZ/lApBLKTPgLT22inDlFeyb50O7
zcOLny/UxdwR/t9X8zsosZfKj/5NMOpJbdk2hj/b1SpV7xYdaWqZkft1s/djAzeO
X9SVbmwGgSUqkgaRhG1u5O7P9tEboiv4JoHbeMa4S2KTdY1S7MWtenkQ0bSFeWUK
IUysPVOHu3SV0Nsecn0a7VEFpbhsDTRnTcIHuIYUHCu/Vv+Stcc57IvlY67jaAxL
7IlB7KCNPY+bR1mgVStse/JtmytzS6PhzoMD4TdKnvF4MXInEN0Tl9PuwgSrxPvJ
ZqUSRJiTjG5oqPriEKlI3QW6KZWiF5zlIc8ST9Qr+CcMCJdMT8Am5NkEAvd0fNGG
T35B0sVXwcymxDL8Si2bjazL3zzlMNCSbhcC6w+vxolmy/bNLkNi9GlZd8uy3HDj
wyL5wM5jxjn5GGqwiXlGaPavUHG10VKPuaLLIpAm4ihsZlmt7HmW1aWkY0QNXcR/
ZS2nJPZObeOxANn/TDpxOHP0FeSGb7JzyaRrQ8UOPrl7JvJFxDjiafZJEI+8KrQz
PGRjF2RGRpn53FYZaI5Fn5z8M5A1t6Mp7EtOJHlqAsa+KehSJ86yrJb3xolkyQoU
ppM1jbvLCorhn+/bGEFXpiXuYPb+05H7whmSOuIHczCCZ1x3Yv86LqlulrDs4hmH
W5AtEhdFfeJUIbr3XiHgfIMBKdpCpb/U0WvoJiUl/ehx76BKhE4UDxy+XuX661Mi
jSB74hTSdV3sJCM0G15ncCcb2SzVHvgrEDFmY5+Q6mPt0A/JK2QggU6AVo6ha32c
vM06I6Db1ryi7NiuHUAb/X8yopSbEQHCeTdfeVhvS7MsLAGTlsZx8Oiz4Fwfg5OT
nSpCHHLPJXKnqHuLJM1VGZRYdONgH5qjh1zU8dI+IMWU8iKj4Vb9TDkz6ELQssNz
d4241NiwtInnvb9QKX1AM7CYTjKwUoVpGTob+B2dQPDew39JN7TkCleaH1/qOmuf
vKcNhY2QiLc5rFHJnoy3iyX4QBUS9yN5xeudeMTpBsdsOhrq/AR0YvaQMrQP+yKS
HA+SL4yC2tVxT2+6+yiPwwxFt+8Mxoag3pucEwrD4uszKIfdQ6wmzzuiCgSpfkPk
AU3wUTdMNv+yfDg5inZp3bV7STFSm7HQfFM85Nasrwet7kej8iYvpAudyek6mFLi
268Zxn3Po0X1YnT8CMZ1+K3VX5RoHlz8Au74k7JYWu8jAMtGLdHG9lUD43Q1D2aR
fjlwCvx9N3VlrhqOwT6mRHf3XB8cZOUVcRZuxl8FUM97Cf13SFsr48ZshpH5YrhP
txhSC5gy6jGrdpVzOqaWBMd7LhJz6MRJAfJ0bLD4bZvaXyvNrA4GUl3iu6mIfruN
+l2Tu9YDVP/1MmKiz6t+lAgA8RQzu6Fj0rMY0Vq8G3NBBPAzwnJUj+X1gZ7wT1s3
9MuytdaElb0asCGiKKJxy8HVgtUmBkFQersPmL/g+qAFyS/BPCo1W8uBs7k1IVQi
pL838DfLNKODe1B1VnmQwzF2Fp8ERkjDVZxQJrnWaHbOVpEvLNmdVZ0RKu+ZxDSG
tKGg9GMDUegsSUqDeWI5xwW5nhcRrZ5yxEwBApTAajh09xOifZpXGM29OuxGUm4n
5deTbJGFvuTunI027YP/w67ti1akurMSLu+OSfyLGHAUuzsDksTNdgd6tehRm3Is
03mgTTnAIwvJAs0IUdecGGFMnMtPHaj/AoYBKPHl7ys0kZyhtgxuFrv3EOlgtDwb
XVF1LTCAlyRaXMaeMUpQzl4eUs3JkhgRyFtLm4gwFEydwPzV2thqaVCDhrEvIMpG
SmExnioUhi2zZOa7HOS+9DxCaYuWx2xxQjzmTtkK52PEWRgWqhwYBPMcKmaoisB6
Y6GA9+wftR5ogXBrqx+GYVLuYa+bOIRvEJQ+eW+Ywt5vDu6uqfDTZx0oReDNXh9e
+AkYHegzr4sE/witw5geUAePCn+470U+7gP6wFikxnZlYF+Ud+RbSUrv9LGtzoMA
noczVAhlMixljlncwLSgi5LZ3eHt8DKIQqDW+MV04uA22ixC65uv/7seY6FpABzo
H22E2wIMN2fh8U7N3YF9zgDYetH6y4XCktSALm6wDOWRBEBbaq1bnoChOWUFkwtx
GqVg9VKUrB9EuqumoISYm2LsVnQ2My+s2icNe3xEktHjHp2V30H9abLF4z97XImf
NtlaKqzGqnN5jSTFNWRDxnC3uv3nNyxSDwT8GFGBPj74BsdWSQG/4lJ7ZOtIt33o
wWXZLV8RC2mmxK3WalATl2Nqe6xN+QqGix7b5uTifvwJ5p4VHYlPRYGIYTYF17JD
qagrPDKXx09qtkkoccTHOfSDmoHrYMjVWrO1gpX1II5wMynthkRH7XnqZMAwQL3D
EO9ppqOVC0D+vxBMuWkX21dxKyV4Js7fLCPdxeyKrizlTPQ8+Z3PGv9ZvHtFYGQX
1AxpEjQI/EYrkljNoNHmjYT9ewLOVz4AtOOs9W6BW6IzCAibk/wlty3GCerBa9G5
kOx/+SnoC1wsMMYLKEh0OFCt+iuHtqNwgcRr117jiD6i2yFZnXzQt6q5E6T2ikid
BQkM2+ElSHPCk4R9WhcQ+O8RRpCXpFJalUz9xc0VYC5AHY/yqMvvC07tAoLxZt0N
Zpau2oiW5MbzI5TebZOEckZGXJj1CP0OsaEsGKpMA6OD4gd0/+Zvu35xZcI5zX5Z
zaaS0rF9gBNLlunXYv7ANtcd2TTq71T5kElYSMFvNPjAJ5EiylneCiOKdEYp5m1F
fs22Pa5Er7PR2qTgpRylM6Qefc4VwRuc325YVeeH23AbS9mYnJWxHLKToULC59dN
xeueQUTy76M/xGcOis9ZPhUvsMoVKgz0o5x6X8zubBdm8KO7+0sr4ibQ5bJE7XX6
n5lAx+taUrPmMhamyAnjA/INUAnMor8lYlPC5+3uVMcaJDAYggh7vXsJZy89LIKh
wJ4NTPIYowMINXINgtQuLd2kk/KDMrUshBxJLZYyCYqITh1gLxRNnxAwt2aP/eNS
i6alCWmYj5Ys7Iu6PWJemfeq3qKjlbiRZzXmQyb5Nhh2nt4yXmDKjFVAypveIVEQ
8f/F15x5bW004wwSMdbTxEjUFH1RaWwsVZ5GTjGuH7HhlJU9d/E5F8NTuqCkayB2
Z5L7UwYiqKJ/8zoikzJ7G/Q/2Uloqm/0EsQ76r3kkzlaInugHy3NbcAZeEkchnh8
RRjG0H4gSS+zd49sK7VeYl4i93tJHnXF676BN09FDEgUJzn8XYONFEb9M+jrb472
feNOz1y+t0YRFHp4ex6/6KzrOlu+pNKc2V/H+Cz1wl0+J8AyQazua0KdTC16vTHb
rktw2eIEljbR9FKfMEBArjsdrpq7DnU/M7bhQcKeif06I26numdVQ+c1s4Ue3HqJ
dYLA7vmyhJuH1H1rolpxkB7yivaFueFXXpUaNnWJrWJYluJNQgH/45mHU0Ir7asy
grSMdiOeiQpRXHArGqkUZ15YXylux+WLO5FEFgjKDGQKS6j3KBOgzywswv1Lv/r4
E2Gckg72C+/xCNwBYEuFRrajPnE4723OfMQ/loD9KMiLCS5Azjnl6HHP6AP2unCU
nN0RlHL6tB3r2kfFEfioEJWG/VEBLYPyEEMMP5kWJWg8a7NhF7Iv/yfG7v1XjW7n
oTWsaqP9V3K/EsnOT/Wp4IFq7ylNjCb95WxQu0fLSuSZAr+SQ6X7tfUqdYx5RAa9
IqP/SN0vo4xHvoAm02iahEAKItvwqbgX0SgScAhtB1wk0A0Fi18qsGgGORYiDYka
Bmsw7GXzzlDAavPNz3KlFsmmnGxF7CMvHA6MDcSOivxldvvgbgomhXgGfQGJGBd6
r1ZS9nZBtq0+q52AtTUbA8BgYGnVBWGVL3PBTAzCatHXDgvueqOLrpNVq6yNokSK
uc3cSeLoPrP6RiE+F5rINvcf1XNBsvJGzbC3Hc4rIlx7Ea1grsAz44ywWag0mgPX
+eSTS2ergYGq208BWhlHYQKkLTZjvoKhW8Lx32/W243zivYFjZ0j8zHnv37P3zKv
nGhoFZPzBNY33VfI5h0IYsx81X8c7une8qWJxrA+1ZEpvl3jRlFNmQLsKHtJATyy
S9S1HHysrTDQwKktQX+BXJhUwodmdRfpwF2dQ/5HnHY+R6T2LP7O97ZhDEJlJtdU
FGiFArlHRLmFfkP4v+5ljIYvgfcKD8QyhU6V3cuwperf7zS9QNzRTezzSuZpYxXa
74fTEGw+rHNU8KI4CmZ1nfrj5Hi0zczJT39UhSuXEE/dMezwpX8O37CdwqB9o1Xr
Or+g2AXuF0/QEEggPDTtBD580QDRVOr5dqM11gcktdHai9Qo5OvLGRADEh2LChgL
qGEvMTeIj30djDlYVKywmexUUELqGw7Z0Adskte7tbXeiAkc+LdeZDAts3HVNUKE
Rka6ICFGGtfeXpAomdS80tvX0TJZ5SIZZumxC5sYtrR+LNCFDzHWuCXawoBSPpdv
TTL4X/+cAg0rKsfggVs2Xx+7TgiAk0P/3f0d8bok+86OFFI9HPOf/cn9pCFi6WCz
f+gXYatQbKfwSLmlAe6HjwWuOVegO+SIKWwepdrde+zQWU0isUS9Nu8IxToS+FyH
l53zK53XQruGc2G89cIHP3+2IKrYyM/4EQJ+AkmSJQrbx211RyAsmo9JfylWRYIt
YhaW5UkNBe1jdgGoTMZVfAUQZJITdgAO31DOcaRzJUfWp8LqcHYNAGTMQF5E/2Ee
U+rdweYirSFA9h2Hnk6W0xeEdIfvhBhf0OFQf01jFn8BQV8h0dC7gizA9M/K3wMu
8SS+G3xvgA385H0VTfIhITgPnTuTojkvkSPHchvLQsHLEaZtOrLDKb7z9lr4x/et
iv4/FUnlU7TgYzzRltqEd6xKDbQB/LdvPzc212L0qSVSQK2VtfVgQxA7fIFOez44
94FgiPUxwg135T9na5o6WG2QILoeyKTAS/l4EuIM/88fY2BNAsWro+lP8zEE4mjw
CKPgW9SsJz2aiuCYOzp80X/2IA0/jFFZpcHgdOyYL7kSlnxtETJ+IfoGT1NarmP2
NJiDtieEYsyBCpD8qrm3H5/PtBD9HU5BnVacHu0Yj+hs7TIeP3zpZCMmZ2DrZARs
MVJ3vcslsiH2nlMjLEEbCZruxuAY2f7qNK4uTms8QBsotcLRx98BjYy3e95Cv3J2
6C73kr8qBfoSwN5pMyAlfyt3lPwfZuZ3gzfcoKMwp2k4uymmoXeLdevIpv1kj0J/
+ZWZz9gR0b7pgUuGnYuCzRsXJQLHvldBqmO9HCFGczsiPSSMVox962glcycmZmm4
ewFrUCgULIz4TTHadKxrdWI6nNHj1uYUhq433DzecXpjTGu8ORyPVzFevaJ+Hrk/
KvXjWBkvI023xTWpeEA0T77qvp7z/ZGSqGs9LFfQDN/DS6Q4ReCriIsCcVc8KA7j
04BM8QGfi6tYYkS9UiUSoVVhtc/m8EGthe6+WgLeOC8HYG1u9Zb3by/LywMm1OXv
BM9n5UDon64cYyornso+7DwKctQ9QKCYbi2KWR99pNXbeS9JJFwkf9v8hWI8CrRt
c/WSE3+srBVUrUP6ExRc2sDA3EiMrV/Zpf/4wM5RBPHgLgfWP1qidgaR1sfe++S7
7nrQQQqUjc3Q1KDyyHhoYeYPZOfeptfizonhxpGvoIYuNXApx4RdahJgg4M37asR
AdRLmX6D0XAjU1uPm5FIO353EZH9UNm+aQh8GsyFRcdMEsM5BqO2zyQH6zv3Giev
jb4lt1k08iKkPP1bKqO8TYOM1cpi4AImfA88OD1JsFgCsyovsmUFDUIzCuDq/Fmj
O3+6AgS5pt4SIlZTWhBtO6sSnSxl2zNw9X2v5ea6bdf+gO5BtUL04S4o/zeEI6Xf
glW0cpi7k65xEw/h6g1+jVpS4EWYPOTIWwohfbjd1IGltfYHZ/nYZW8liMz2QJbT
uudBwTV4mWIVcxlsC1P0QaEd6x5fTBChVom202LWc2P3fEuosb5K86K07kmcsBwS
ViQI0wWy4ul08TQHO91jUuzcEdhuSAws1lmIc/EvkCYRJScIQcGyIBduFPDPMeD+
q+il7debMJ+zwbj1H2FCXNMEvdGG3baBMdTOHPuUT02zQN8exIPgmfkrdCh7w7PK
SSzjnRTim1SN8LBpDEIYFeVc1my5sPp5GJUFGC+zuA/Gfbrtro3u9fSmAPsRfXMC
YWpvoLR3bUnPhTfI2mw7ZpfBgnzeOhq7CrQVjD4cvuIHL9DZB74z+ODNWbU+MlE1
4hi80RX2NguyGMlXjf7cyGA+zXNYpaa7n0cvzKqebX7hNxRHJLrSYBHx+IxKnCga
WdCEZghKdu1cDPCeqjxVFw1lCYSHJUJLiFL6vnFbWcWkzFcy1BrKm76RT7eUP6SE
PZBieSEzFgx/vX/hkmwtq+2Z+sS5CsAttApg8njlW+g+1PYCZiSsCD5PZlFeykxC
xsrNLhEfSVaQgkemsC1HHtWwzpVtla/xM1kT7khsHELhBRAkz9Jt9uK7/SwMd6uB
r5c9EEIJMEz7ZnjlNJMl7zawEHLy7WZTDP1pIQKXLDhUJdxLEcTniDBb68LefurG
8iSHYN7LNR4hIChF2TT8PDbw/dt55n8QSyO9aNv1g1QItM96NrLJ7DJz/A2Seqzx
trFtPeWCL3mfqJZ8QQIpzC+zTqbEb64XO3vy9lDufYkaWHDkNCjQlMYU5B79h++Z
F/C5V18soTN6aM56cHhjW+/KFELxoTFyTlayq8jKj0wWBSrRKsjIPupkXXfUPGFb
jt32YIqCWS7exiQ/nwBLnSFeuzvo82xSeZ/0dwy8sPAsBWQpTORKSjB2OQdnyXox
rCE7EQ7m8rlY0Zu591iAXODtuE+rIe/nJgQL7nuSqOuXaUdcnru3wNwstphIZKvw
DorklpnFCBqUyVeFLx8eAQ1JeaQzFXs6avso5zqAH0nmmp53UlD6hMxPw2Ck7wU0
iEUSrOFnOSoM7VcoC30GtJEua7xUg01qfKX5fw9XJm8Oy8TchmMns00RSDbZHpsQ
oOrh2HcTku5hyCCxFwiVrQFGKlh0zHsmtF8ieBIcETtt2jU/MLz5o58YmHciuoki
mAZ7Ac6rRfV7pm18ZyREMLrnFlzxMQ+YcVO+yUTtNn0CAjBasB6XzkdTPuGnlX5O
wM6xdaY8IKsW4YvoZNJczjQ4BjaxquexFxmWf+oosVPAmcBWIN2CxjtfoCLl0NJj
H6u/GOEBeNO0tCnSNHuRTSf50z4YGM43cRV2n45LygDu9UlIMPTbPVGmITgZy9f9
vwaUGNwRREESXuzshIm8EOvDEu8Mkyt6pgHQuu7uOPaNizNpDFYIZn0uXvj0OQlP
lCJ+6N1XxhLpZCvdXx10sr9heoFB0kt3OEXvvMn51i2XQK7mF0FuLi/F+cr62TxC
Bw7Yy5eWvHtowc8iNQstAhzdTvSag94u7U2OguBiK8FUY8tHH+SPtHI/GoVcbIbs
ddhAfrLbXSNQwZS/Frq39gQ+/pE7IvOXAqeUKbs3LBS/kR2bhRzmo7Rj5bzoFsqf
jHRbKYIDNLLNoL98ZEnR1Qvm312gvzwxtqU2vTv7R+naPfsLUa7feajP5vrylFPp
D5wLslcsUFTdRBLXLx78a7KN8mU+WP24Lx6bpY4Ry23llyvAM0CQs+l7JmelSsxB
SO4pkTHhfR04OWdWows7Qim2uabOVXlx0QLk+x4ApVhN5xeECDk9R80gLV0IpC5F
WibxvQbJ5qnX7e7zMoQrKI4pRda95aVW43fofx0z5oCPFv1n7ZbZrY/0foHdTq/5
7eZGivjTIP5I471eA1cvpicnp/+caZMpOdFlFMbPRv6RDtiYaHBxprj651iQDO4n
H18135jZWu2PVCNOr6r67RFIzs9IckeFoVmUJUwEx6q4UlNPGAfcnCtzr4aneXXb
4nUno4rQfVnTWzGzHg+VXbiXYolS17EoiwB4OYM1g7ZUtWfY7Ih2gf9ri8PAPyJt
JYhsWuCeJLqPL77GwFFhgbiDoO2BGCL3FHxvgVoo8Bjb/wBklLSlqD3loyOktdWu
z8SzDF/nRfC0S6AZchTW6zCUclBgqALg97gKulJt+NSqfrGF8QpHoF76dcWACvrY
5hRL+DvcuUtKVO7KJkFfI4mt5Za60Hx5BmrW5MsYVf9qMhCF6syYGa7lueqcNiY0
SgXUtX209t9kUsqWel0Rh0Bs+JZAYeCbCmFO55VHukdzPeNocn2uQDB7oyF7fKz2
r9csWunejmmhetNnz1uEIfa7SvmnEF1LyLXqAkH7AAU0mayi+rW5CFpLP0anS1g+
NZwOfdMeNN9z6RxjcidwAWOgsAwH3+WyMvad5JIZIJ8yUA4H72y98m1yRAAhY1rx
BRJVu9uvnsdKX8W5lDpA6TJdY1nPZV3deaMQmLoFQ2NKcq4PMdVfQpIq8KET0Yp8
HIej3xYE47tIO7ZAAhN/CDn9SOixZTarL2+MXpQv45kAiQKKZOp4w8EXn8PxX1w9
JNlfUfxRDZ2jwD1k2U7CyNSmI2ksZO4MWTGx0guhDdkL4LPs0o1nKgHOxGORaVzU
ButQBGCnGXrW/Umi7o8xa0UkJxiZf6AInKCsMiMxfZO/Ik+GtgqvjMunzJy5us06
fW75Kw/ervUpuDhMEvY75eiKpk8c6Y31BsvReStfaCDZnL0t0AvCXFIBCfGVBoi6
rsLj0CCaFZ01RGXduyhIsNVZkoDiHT0tnIgYgmcgDSbTjgJzLv11AflL5lhEbqQt
SNdvIyycJuQJrhp0nP6UHPhDNwox4sasyW+hDkeFXjlHhLTmdAl18ZMgNAE41XHT
j1jNjcOEpzpPPOS/6Vjj3gLsU2EWdY/ygzfgGvUiupWpzCGFjo45RrDLIwMtcCxt
dQxF9Jq4JiSPZWjpijOku2O5YAa7OoxaeNVOO26in/APygzaEEpw0z2phcNxGeHr
FZBba40tiUKw2/VPHrC2XTivWjrYATHStcOj3zaf6m9eUCpO5eCt88WnpQgrl6j/
hRj5ZRkIPxnJ55yY+FxB+DgVT6u+ku/xbegcAauRUM/h8BanzdWcD6Flpjk/tNnw
4FztpAw/teBgCDxef5Qa0C/RE1bDzFXDyB5/eSnhLnFWwh2BEiQWWvqTwF9TXfQJ
C+KyiuhtdxMUuv+6IIFwBtbBaKpEP3IMqtfBqW0OWXiR6j4vlZzEA5HWxGaZuMLp
4hVA3OqIuU8UdsonQyNZZt8tWcNtP9t+aMcmd6tgaLZ+t20H0KD8Wo9Dsk+oLaWn
5k43izfwGD/AJwFPcLNsH8EXt9wJYluqmtgthw7bOy8hDMbgFI1kn+qsniGCnsY1
JO9E1L+Q8ZuEAciDty/UF83lOXitXent0H8q4zNeqtQJGLzXi6M8rymOadXt16vq
a+VwmLOEo4a3RPaT5j5OilbPnNWVpOl/a+HxKfcFgaNooYtkzOHSEsx/AfW5akHM
e6tDUoW9malxJbn+/aJr1Xvo5Nvbe8xpTB/kBVPRCIueyrd7xGMAE9rLVPhhGdPw
C3DyGREwZ2oOLgiK94Libzsxi6mK8saNKvxMzL85QfW5W0L8Ua2XkllKsmVGr2zm
6ziib6efgQyLDGqf7rEIo5JIPg7rTg0itFgPQviD9ME3BVIubnrTGS9IYFpbRbes
V2ym16N1hfbMX5kWwb2pSHluRsn7BQUoq7bRNYb1xAZWFTmUaKJ7G4T2kYLaq9BZ
AT2RErHRijvI8dS4obFcF/4KYxCCA2WTiIlaldMMHQ2kNjy3QLQs9RFP1I1iOv52
nK8Nv/tRZPBfQPOb3yFZE0ASSClyJPofM7L1X0ULrgzNm3ch3YLjpW9+EpSc1MhN
WFO/cSzzONFF5dkvv7/MKfYdjZlXveURb9ux5oZZFzSw0HdDpOGfmuXocGFmwI2I
3ZPidNJI9XzIDpnmM3rMRs73K7riXl9LeZfRMMaXEjzkuzjmE2ilT9iKCNQ8CAnK
XNLHDxB23OSh550opoxaRYlX6XWVpLZ3VMB5aJcOz+KXniBgaW7hLU9FSBE+YNfJ
mHOlUYjui4uxe1Bj4fL0XBagqn3354Y4sDQDFFWMKqRRcBKJR0gtXFvBFu1WVZfA
aUU7nk0o5Rv608DwzATsaJRL8xZiSg8PbSvlIeW2IXi9phimWhJVWlCJ4+OlteDs
ppMy+8ZcgzdbZaIHLBFhdUKUZ4je7MRRJVV56rWodP4dPS1AWusJZuQULK3urKEh
fO6RiGe9GTxz3RMjQRTCJ1lhunTX8+sJ6P95RZrTUWDbyiX6fymvkFLfksxzo1tV
5wIJqBSphdHZ5MgCKJauMJDwB/EkOTSqBrKHVqxpabxueKWLkbyv+Bp0NRPApPAx
Eiqaq8GKU50NZ4uZ+x5z4HfSe+3j73zyC9grDHKG+9n6oap+TiIrBbW0fSlwXGyN
5zxZzv57UQuta8IQ5VW46ftS6t5xlEHChVO5DIva8nUmYwhs5E/meGFFW8ipi1VV
+rIhtsDSHdW1LSx7jf0SsVkIg/M2HJ9CQSA/XnxrEq0e4MKNnU45kjY8LW7lyMl+
z+DCCQivkYEWyYN7p2DqjICX9Rtip6enKnetjAggQn8B5SPKDqVRF5BgjevXD838
U2zIp3HMkMR5JwZdeqlFtB5PQpYfCZSigo0oW8TnP2+rUVcjWiDGhuj563RaZjkr
a3XV4P4Ud+c9qmNmo6Bl8EBfCF9h131EUh1tq42GTVmYneCs9TjXl+gE5vGUIBto
lHVhDo7OBdrNDnFPrqeMZgoAq3ZkvSt+pCXykLJZcJJuQadSn58huxZfLijWdzoA
2ODrPt6kBDZvuO3OOtLJ1AtmwOMbnCnFcD/sEWeGz21FKzwY6idDE3CVFzwiwSu5
rm+0wvxOQfV8J3QaKFw+gCWollIXElQLBmyz9vsOkj3TvpY2TGMzotFJtJL4WWv7
DqNZUF4FEghiF2EbhDSj4dabUD9IDEsWSxzpX2r9dyGpgSGKw1X6iqQC7hHw8dcq
rphHipDmNGVPLuP/gUEEh+YR/rNdEZHiCmYg1JXQV/mt1PFxNeI9av2rlHbGePjR
bP5SnPLMhKhi/biRFb18b0D+Jy4l+tM6RA10SNu9FCSGG6Zyff8cCeUvyzrSTnon
8oR/zh59GAp2ZWAnF3o6VT+gp99oPJX4py6VA5jO2qZk4hOHb1hvPRfvrgH/6KyK
ui0yIot1UgXnDmnaTL12gR/8yw+F4IdpCVU00w3bWZbU2J/4PJWsTGVQLd+zzZ2i
0+eiTjplDw6qIVjwdxSl9pbvNHjy1B2yhW9Ux/7lGpfkdOCu+YgB4w+XQ5MCgOX/
9iE+e1RJ1Bj93oalsR/CtgYAaXl52bIJ9HwmChvugRWcGaPWelMS/6u7lsJyKFIq
gIJEoUgzzrUj/W/PShz6OTTjoU8syCyAtzd4TiGAaag5cicE+3ry8GjUqc1fz9st
3LCYBH4sMvrzZKhQjorbwzqMtCpAsQWctGhFMHfwlHWvmxZtScqeGB0PU/Y0ShO2
qEHyXRSKMqVhTVPIYOVxrmLiq6fakUT1hUB6EemJpbSwfmpo5P7RHKPqPzPX1amn
+ao9oudaZft407X5Q1mpwyXxAR3sJLY4nhPZ93DhHuaJZorqnIpv/bhga62vCYe7
uZUNr+t07IZNA0RKMJ6lbpvQVNyQCE5WXqg/j424LKMTqkDdX4USPkTtCrA9ojW+
kIe9moUICvKVp6YdjkZsulUTsFALCoBflzQY+XFy9fdji5ysTbF/rmrpoTYoiG7T
zGGGSarxMzixTThvL+38wexjvcRCr8u5pHd8HC2aY8HM8LUWEkYHMMePrm1ZLFJW
ndqmswYBHFAZPlrbcgs51UaoUrhN8o1NtSq7Q3aazRRUxxxwllMHtbEtzHpWkbZf
8lneTKEwBC/CkXs9t3PQ7pjXZjU2WtlKpEVvT+xxsmwyKYDFOyBO+Lda136bLoMV
jwqWRqugRx8zQoKk8LfXByTv0Nagblmw3LCmNgYpMM0yYADajblEyxdzEW8vps91
6SEGGeZXKmRCYOSBW249rxYg2+CQ1NT0o9hOQ/88/TmjzQBC1XbrT1tCnCGeoNGU
GYHv5RHLYB85KXILPmherTJDVvkm7PlUnOD7rgD0XmesuvQAf+uRghNuR8AMwIjR
Z6OpjN6uKOKJ21qd//6kxrPWj1OOKCq3gbk8krQvraUmXwpHNsN6qIVsxNW+zjk0
DTFSvIP+1rTIgHMizLdgtn8LRj5loGKNVsSjVuLgxmc749aIOoCruHpLlip9Eyfv
VIUZWGq0cQET8chi+22FSFSLw/LcHKbSvglHlc2dw5QSfZtytfZA9R8XRX2ndVHi
UHH9em81X7uIm9/Dy00HdCJrCtOVCp8Tr0Zu/a7iIRYi9X03NH+LVzgqCjyTi2zj
L6VAH4Z1PE5k0ik7GdtzcNl5EmXkUFTDvwelD0y7k1djqyPW2n7aZ2y61WH3XhaC
JzCgOWYPAeTQcbaApLRdiEotWcjMuFJT1KDQjYwWfu3ipW9pZmtK5V4KnCiPE5XF
IMPHUzEpO1oixHZMnw3i0Gi64YNOo0INFGnHOZfdAnGVOaNFh1zAQC/+3vF1Eqo+
KirK0nEDcxSHqrigzfY5YUqxIJv/LL7ODbGo1FA2lhcm0zjwEA6zG5cA5gELmxHw
nhSDfugPS5ZdrxFZ7IVGQSjEnxlisT8xh5e2Z4gIPcsVUpBDhZ2DxgxrFtKFYGuJ
20E7gHbJMrwi18UsAlZfXjlwOAZKbQApKZp0nNumELDqtrndfJVSuV39f6NNsQBn
lDLYyeKbcVKOrf3fEjxWkpcFuDU6DCM56PjqG76Zv0Y4ffn3MW0cxh2bgfcHNbZg
xHUkNFMLSw8fTBPURQ7yTGVzsBZaSwQRGxY7ADZEE/i5uJoGcSilabUiJIUrQp6x
EBpyiFIOUnq0P4JU7d4Czod90dLX6ukk6nnHriEgc/0U1PfIwaWHMr+bYwBWzHfk
QO9sdJfOKSHC+LAico2r3YH0dqSBulmciqyfFo6oVUEqYHCFRiiCyLT6opSMScwL
pfRwWtdXn9k7iOaTC/+WR2sjRLlTTk9x4NfUL9ve+WOdAt0hSGngtkPOqGYnVXct
vBN0sMplALqeM7Gptl+xL3VfD+eXskcogU990KPDbEoEV1Ecpt2n6qKStSjbd5Q+
m3+F1shZV6gUuwLQqcw/Ue7ilTJN31KsLsUV0Rhv5thof/ySMJpltNopDnUWfLLF
agv0v5iRbEN03zykVvYOhEgctCNkYg3LVN4VMMRgO2CLKH6neOktY5jNrfWoglz/
7KJ3UPHwk7Nx+2t5gNcNC5zLxabUZGvBg6kXR7A+nmoYmgvZdBUtJrLOLR/VPVYm
EqBwe5Waw2bcMNWQJYr9cORO9WdBGHZqOfWtNEC/8t0PHn7+HZ5LWJxAWfNKR7wE
1QqgUt+xYRcnZiQQggHz7K6iEcVfZbFy56fsbCqy6GG3CXMH9NG9basOCNVHrNVu
BsH9FFGrL62WU4qh+p1DEe4RcR11Xo6YCprdNf88P1B5e1AvDeY9LDkZAwU6FFkQ
o63QXHHY/zofifrDIHJ+xe+LgfbEOOT/KNB6v1hcThqNaItNxAyTF7HiukLF76du
0tLorMA0R4DqBdtYKS5gl07pL0lF8EqAFZKbbf2ynYbAaVgUfm2lz/wMN76MLNwI
o+pzhG/fDGROyzzl6mh6oVH/lctoXflRTMW+ThgVNWTWxKJmx/z1j6y6l0HIYAq9
zIh6Pzzw3oCjK5kET1PrupCFB8plsDGsFVX65fJ+IICP7zWJmfbNopfqrt/Re8/u
DndLj6BUHPySI1Meoev04lEH/4TpK8/f8pifROWz+/sZBV/EdlEHyYnK5DRJNyhM
QZSJq59akzbMXbLzU/n+OZioFjPXTRkq+JuNmm2S/Fj4d/UIoq/8KT6L903e0BPf
VxPbGgnrB8otGfUCSm0OdpaFnspO6D7TzKq5WVaMmnNKkqvyu5TUsAt21h92AyEW
q5W7LKOn4UV44MGEmX4DFq3XYbBwDUSAEGDHgzp+0cXM/SYSFKrP/hzcvW+dXDSO
wPKNGU5Ek0tF4NgtQhiPPBBUCput1it9d6bvyEGO39IUKuSIPvJTwOP+mjoaJSyl
7BgPrWikZE/YlRzGnG/9YDP+DVAFL7ybMh7U/W98+3UOMGmzVb7FemlxJjyGknRZ
OjQTToLgQa6exYBEAaSgU3ZVc1vWmTl3O8iTwgD1arL+Rbj1CeZs5KfkntP6xuDt
LKtNZ7/W2X0TTjQcom6CBV3RngCy7dXHis7scO+q/UuZABYOefh/XwVObwRHg13A
g2a+KQ6CGZPCI5rYfjOhc3ZozAh1Gak7XQuQd3NI4v4NXoL0D3Byxvgn5/igijCo
poXAtn4ieDsoLc29aPJUuHxrXtOQozQHTSbh0S7+4aF7H5UDhikP4Ov0CZ0yLD1t
apeNe5exiUyxS5nj3y6zEDCxdQK7qbNoYzZZoYGqQM86JgjL6OoTUsWWrxLJyh01
QNJWQdhlWFg15xtvn5awrwcD73HBN+X9u2jSTNb4klTOgkFwaay5sSp1d+TJP+nk
u51CQ0WOaq4dFFAaCcB7YuzaHGwl+caR7zTIpZu86zSizGCIK3Fq89dMoXRclS6W
6iJm4JvkgXM93HRbb45iiwzTo73X4LDauO7QaP8E6phZeUYjkfOqqVAEHCKr0keQ
9IBJuYptAWMKmgGXFzrQCPlTdamGvKWLxOEFdCoNXugw20hA2eXsjQCE7sbFpQhJ
pKbFciXCPzsBsjGs/I5FrSaD1MS8At9/nA/EFlU17VoPZ0Aj3fRtV0pWbLvgEWYU
SydtWPuF9UGkyY0WzIIMdqLFhlnGA8c3f1LEzW0TarPO2TestRXfRrhrN1N7ES+U
Gox87xMXOL0hHLsGriIUElH9v+GZ27ayVZzDzhHVNXBtHsJ3xUfb9s7gsW4RDH2k
MwKqJfpcjJZC038lT7ETGFfU81L/QdvICgSFzj+YDY9LBSNFZpq5lBwELm6faKSS
nCgux4giTu3k2pzndQ5d8o0We2idawfhsNG+SyuogxHojKcwa+NiuRmWi5Nkw2Ew
wBC4yOpKSYcePz6A3F2Jwf6zB1u/CZ/Egs+TBaDUUnWUfI5Nw+6srwWnVfyShwNv
TW9iev1VKQgtkQ71cESYyY7C8AY4nKKMTa1wLwY215uCwwO4AWKF6mc/VpMFEPZU
o+9luZz3W8ysESDN7IQhJn4AVYy9SZxWEAa5gEuDF9F5TdWsy1uIgfHbq3SPDmmX
FIIyUbg51NYOXyrZ1Sx6SasbKe84XUzMrUX5QKQaLzizvy71bWh1DqWB7NJgKYAr
UGZxduBMX9IXM4MYacsy8jum5a7CauPQfX2eRRI/dhaJSJp0ba4X0NIU9vYVoKKV
HxuOyFl60GGP8GuaF79aop4Ih06GAZWJZDcoQQ1S81KfkJbLho15SC2LC5gy3RUI
466bek+YDaZrMT608AwGvRPF94AEmwk1L9NA+/S3UPgz/gF3P0/OMQSBvH9F+L2r
jbmvPz7viJiBU/eHzTX+XCSnqea0JgBB8/bEVMyMoiVoIbXysOjpM4pllBFba6pO
qhjmEP4JciOk3enmv3DDwWiH53+yeIATMS+XxCkTHDIrVp7COUKjvShxphDDNPlD
jB8HsNU2DP9qB4ZuD3jC5vr4IDLLYLoFut98vXJyj5wL1DCD6MJ3m5+919iC7s88
JaqjWy4SqXpKd31Xf3JO7Vv+3xdjhT00ipFEQMTnTg+lTnyeTuP3enSe4JvQLomL
U+u6xHyidET7TKTPMMGuNJ9S6ypkzwoZoLsHd5QCpK7QL62tvY0G5o0uQoajI7a8
MbmWgCEB4l9i8uCJGH5rJ6b8nrlEzLiyRI6nk4SyY8oK749KbELh70k15vsF5eWP
jXXXzYuNPr9xmw3aykXbfO7zv4I9Y+diaXRisdkkldya/b+NE7qg3pWOpLY395oC
R0BUj186JVQv+6MJXBJ5vfy8QUPxkjsmz2eeZI9DAbKYszUe5K2e5fRarcOBdNJf
bqkWfNYtyYytaNdrXTsUci95aE8BNOI1eNyoUNS6nd8BQ9ChnoXkAdmxntgUJuIJ
X3lxgmZPP8PPcWYVzyOaNsCOhbRjrlaob3G3M3HInZIk1UQMFW+pMwpQeqVl4gEV
mP9vHZKSAit4084grq2Anwl1ovmiEkPwy0/7Z4xH0AtqR0FUn5caxoZmX9auCQJE
76HD3LPThE51WAK5khpPll1hBWdMIjMjKEY11cGVxJGBFe/r2M8AaNPeb42Exsrx
QrYajp9UWxgch0LxqGXDGg6qg257UejcYKc1wGt75L2uxF5mJAFXU0gRscfadKIV
w+PnKyHtGJQZXk2nTgsCvI6UIlXfaFM37iiYbWT4BMNfwpypO5ghGn44k3U2vn/j
jlsRfLMRvcI0NPB4EngTiiUWZvFQgigZwsIo4PexgJSMVQIxPdzDYCHhKpYM9XuG
MV6hgQEEbbDG7G8Dr1zCifoeq5+YHYLqbRayLqL2ZGMU9f7yVR6v0ALVtyPyKD8v
BftwrLoh4dDaJQ6Ov/W/DTfA4S57o7V1mD9uIwgYMIpnPL1DrL1hcRA/oMn8R2Os
yKNY7FG18X/UI3WrgKQEiKf3uvjrQfEbx44FIIBSlgfGaxPVMfap0A4szZpi9vFs
yICe+++tBhHkT5aQLlUbEfKSUUYJmo9cmK4+nsp7VG0EhYjnfHSDEs/WzVHNIBV3
zz6UjfCo8MrBsORwlZZl5Sy+Jop5wfJPXM+QQManXIAulY+DYOSTK331drNEUS9n
rH5y/YVPPZE79HY6ZmwP1GIem4hV6Ka75HRmxNvu5wym2ymVMZqfT1XddvQjOeob
cDLdqGegf57LVIKDUZuCd/KHkObFLtl6G/pIjodYYccmkB71q8d/YlxNOq+0RSgH
eIOIGvW8rsaphsh10nG34rIw6dVwBfGOM3l/aUop1jXl/tDk+3YbXPcBGh9S4jf0
vz7djM+1KNDvKzhNhIoYkBKdoLU7kuwdcEw3cJqxtDJU36Y+3Vs90KgYSAy1vkHz
pwihr6mftzIRVvkOToDqwTAIt+98h8aaIS5LZtFcUGMRkcNSejfTurYH7QizIN8Y
I185sABFKUspZLnF6Q7p/VDRn19+658/olw4adcuTo339Hio9rJyb2pv6MvTW1nu
rjB3ykCZRDxfojmWWkFbaHZqBn1GURCw2iduy4jZ5MVSGliqLu/oakM915YhSZhW
KrEk+KWo6miGq55tqtugSkvozRdeC2VhgTa3hgnu1wxk7z0JwUjA4BaXyL2uIUJM
Qn7IvipG3CTH6u+Ux4sjBC68zsA6ppUozqLQwOka5BdhXW8RL/TnlHjF4WZ+zgzW
Wt1A2bJqfwRqiKu1D1+oIsMOS21RFHNFPS3QGjgaOkTVupPmqquEqhMpuwJLkEFl
/vq8YsgqMbC2PdBR13scO5H1hqtl+IFYDSaROes0Xq30B/VfVHB2E7bKKdGTtp0R
jjQpTG/2yiWYb1nWTK7oYDb8l0McxP38XPBdfllVPv+H1afc1DmDXugHtVnFZ+vY
Ne9kWHlbUKPE5TuZjXWhYWk/hrKrPRg6rLYRHHrjMVvd8U0ICopVjKxu3FlmgGTV
DA8V3eZsCXRkMGQ6wedAgi7gofxToEkktnkI9YkWh9IVeqDqm1xatv8egyoKIdzY
L0HHgEUrEEnWgPZf1o/yqf8f0xbmbHc4t5CV/FrwL8OOsaD6iNWqHUQmzs3j+U2Z
x8o+7xAyTQFpBiy2junbtOzHq9xKYZ0KeYvmcyQBXE/hBQeNb4ypBDqgoymIY4cL
QZ20eo33IjsVZJuwBjLOoiicCvz6rPoh/bhrMftoHAar3JI8lJ/btleWQqbYdBy2
UG3IXOhufh0DLXcroAx28azyXPiagE6MtJDYeJVQbplUM550U8ciQXPzdAWwnevV
W9O4iktbb8IzlFmdgz1ZsPVNOfBxmTZWbFo3io9ec4c0cha7HwvPhYqBreRICQXx
Pxyhj7G3NTuKhRYPjJdyVVL2hS/cVthqQ1QoyygN4OG0WVnhBcEmZT+2yBZXdIuB
nXX4wBI558/WMUbODs/6xfWx1A11a7DmUkwiBU7okWop+WESrOzXE6R7Wi8u9Jx6
+N9g81WRSQBfnObPu9/sNnNrayDtmk63bAo2QbtcVmphEmh1HCDxf2zcggJ+F06e
/IH3urQwfeVHu6l7Vjtjcsziw0MESD5fLTQkKQkIMOsyrhtbEqtRagtKp93e1st6
TM6R9D+G9W6lw0USjjiwl0N1Hw9/ShUUH3Y+xa1Ia8S0Lwdd1qE2ZaO32B9nPrh2
xAWNWZsZuy5j8oS3Mp7pBrBPqkmC8aHfn0YTpL3psRH59AWYOKXNVZsAH4GpThRR
JhoUmKVP4sLr3Ae/6aYlVUMuZbhzDmClXDlo0RXuZ8tISpL1Inq6cj70cBU7NrWr
vJOgfBd44Pu7byc5olWyUW3KU5YiofNSZnq3dLpE60k1uYUzABmuMa4PpsV4m24S
VYWG4lnmMvxp6PZhc2NR4IBFuI+DUs3YF4718JuW7eibW/NlB8b7VXJGuQtZG9GT
VIIoy4JCf8iwSb5BStVJ6NwZz6Oz7wHhdA4wirrrflIWI/WOJ91iGD4p5SS+k1mg
hze1/R5Tp+zWqyDBJ006fSgDWughSBeJllCkHKgXsUtyekAfmTzIbQk82x8WyMpp
vMu6TPbYubDJvrr1lZ26HSd2OWyqcYsR5smlCh4UliXLlyICBdyCX0fkN4OceCTl
CcbwgBsR+C2IP6Bx6DRyvCNZ6CmyyU17sIEnSHMGGDhNya3lit1f/hyujSG8/b5z
KYzOhgsDpxbi4bPeEuKrUaVB2OsngcAFYU+YTl1V2llTmTAQqd+rHMwa3y9IN2Wj
Vf3NIT/QThCbIb29yhiFKYUhAykVjwmCH6M3bxSIC0p2hEQT6fVqC6hqL1IVp2Ew
3KhFlwCl4wSj3MCgUnbuplj+QmtrGU9UqS+THMJ5PRM2nCnzoofW3QHcn2Th/ef5
9x0LngSQQVI2gb1+GeVGVBtHcxP9PsKxr6MQjVeiGY2LoJiAOLnqD9YorOcqtBlZ
DKkueiMkDocA2pgSfCifcNdrG2GYZyZSkeiydBcIjBNr4QkRyhgyEHDtF+b/7Crv
iIt6qKfmjdFC8ZQ2gHUmfOdSbzw9A0VJECmif5ksuBYbu/tcX3tMpOu5ZVbATV2h
CJWoYD1auZLwKWxT6AC2ZKdEDJ/kFG/8Coukrz+NssXK3DhajyoDgL0UvmHp2hNC
mbVtZTAlGlSF9YQSTZlalbI0/O7HaR249TvZMjl3rfJUENnz6sexfGp5K4Jrjhuk
CvDXXyF462kZ9TwmB50fTTeGkgk8jP9FckUTUXZdqiqw1u4L0qZPL+ihsOAYIkGg
7Gbiu5ZYAuo6NS+1FIUiHHYFSeG9iIaR+rKdhd2V68FN9fKbf1WIYsRaHJQZZb5V
p9bMO+Xr7nDnCnN0apdOq7mfvvzGTraoYPeMEprTlTq4xigIOBxLCFVxr4trEVBR
5w1iuxVyMZXXHa/0bUrp5Ct/VXeOYpq0/GgOzOCQ8ncgWxVNVSadufhxTcgF2cRk
27TJMU3Db6lm+7fHdDWtRVYnFQBpo7/WelDNuohoH9nJsme4hSnPwEBiaDPLyOgi
rT9Wb3UkVAGdwXgBB31XqcgN0hGwdGCXJM+Yueb5imzQwTzPyBfFIWA311l+d4po
SMeJCTBxQXwrG4mdTYN/Vv5INN/sEnGKINk5pXY3/HZuNEWGWVR/6/oSoxDjlURK
fQdS3njWbgZtC+VIRHlqs0i0IBfUxODJt5rejMRXHjazwWfDiFDrwPTdCPBjaM+1
dCzr86iPSUCHRwaHMGmZA2Ro8vJgpyez5by5zhGHctE45tiUTpcKltmFVwRFNBUb
7FUzRAkhabwomabVcT2gAqHcidUYB/ymPvjdC3DgbDXlFeUzzDMOx8S/U3V9Ee/X
8dUletcH8FzkZme3YJZuUptAtZIc9vjWiMvcyazFtvTG371gdjFyAj2KaFKx+eE9
Pb7mNvJExgV+DrzGweiAMAiShNIfK24tX5no9v5EV9O2D/x9caGU/I3rKKZI5jLo
eu0rELx/zQ/OuS5QEcYsch1vxjfy6dEOJHH4JcFKYRC30iOSVy2gzJFm7DHQP8J6
BnEHjxofM5HXfxGJHRkKpc4vj4VhWDmZhezKufXViYkiRhDT7gS5VPqI0ttKqiBH
uyXUfVDSd4Y+AEmyCB+3bDuL5Oc31PfSTL8niavc+D53uEsaC7Rqnvfs3jhDph7l
qgzBoUIEcmyP2Zg4mTsJVSbGeXfLQrVS2Dm/04eFAaBu9osScyVDKZU4JCPOmucT
0vlK+1pnEs/l19PLPflpsGhGZpKiELFip5locH0wCLXtzhFynAxUKUnnQ5Go8YKm
6JxtdvKRrWABmwLXn/U/4wkuhgUWk3FS5OWlwzsGfQbQbt+cVcbja/hhR6qx/bFh
WdFEDtClL7gYHr9kskUmTUUFsxodCwHUyTPy0A6QEsytK3h/ouze+dn1qAwia+R/
aAZ2x+cHv+poobT+g6AzjcY13M+ork5t6PccrnMMwTUupLawv74bNsjrU1OEn/2F
sPoOh6WF70G0QecwX2lA2eGpenmvXFtgP3aNtWq8AJjl2Qfk5AGuHo059H10XtiL
ygX3DCkJPAW7stpg/wc8tcYElYX6vYU5cBatBFECQ6M58GgojJXk8bHNpeeGaZxq
y+Q/9LhPwaAvBaJsb9e0FdFcWOokiduNk766b+jYLQ8kJBuHPx9HoIA8F+B1M3Jz
Bkm3NoerUoFxaZs8u5OoLZ5P+hQB+W/idjVcuwzypGzsUbWcVG3sRiDen6B7r2Tk
KmkBb8K2ySJt/zP33jETk8cMM3NePvlJGzwfbtjFQKoymTxN5KShvnrNCKtLVn29
VKczJQAgvStTQwcB2JkfhFtbuslucyrLzwimq5fgvLdOuW3TBPhv2q9+PAYqNaLb
OM7nly0f+dueXDTKGcB4YGA3PPQuHeo0G2nbqHrvDhkJ0fWSNUyRF4BEqjdbXgcb
c6Tgl6L+aHow0fLckd1StOZq/UwaBZYTAwPp3EYRmImUC6NLODBRfVDnHD/9P56O
IhrrO7BnNnP4KvOR/leAaeF1XPl4wVAL0qtsRTq+PkF3+4AhQykQIafli2/e9iv0
Hu1+aEvz4bAPiFfAcolNQQmSNq0+Of5uahYiW0nzr2P942mg9i4Nut01sQWe75Ba
vCooOHbO1uM/s4Gh5/Ui4YBH8VTp1O7AfnVmLlCAgc4ctr0aD2hCoy+JIpVNKGC4
AsQEEsiIKSBP74Ydipkop+0iadC9dRiMHpvLOo4u1pVn4TvZhLUiWtTokxJCbDgE
bwLELVVc54Zr8DBStpXl6e7ZSwHCeUyK5B54lJVLklZSN5ncMBq51a/aHaZn8xyK
MOSw/Ph3jlbDq0QdOpIYZASPllISPoO4FZv4biuw0nZqjdAtqbwofhYPYm2XPxRt
SgbnylMU4L06Akgf6yND7Zr3102/X0LaP5vPUYwvNkJcIQf4y3b3GgLjrwaRX3Nr
yBV+RYo+VdGPpHzmvb1qK91rLnvSjOYhrgyDxEAL70RTzBzs5EhUhePJacxinE3k
Jr21Al9Qw/EOtp31is32+mb19vh4pEEQOnZ0C0OLDME4nvsFyYQ56p9DWPVPqnio
biI8c79CAg+scc84mrIFjWV++0Q6fVSli0pF0SzjNm4A+Xqu9aYyhcgrihIExmfP
7bbiSxTAcynEQAYkaA2WztFuBQW5h4Mm+DNDGNhfN7cQnNyyJ0jfcH1G/1vqFnNU
RSPWEAgeO9QkGF0CpW5NqXCmy9yGpcaBNvCEIq+2/ysKTIqNBPsj+3toWGqYLDJ+
dH3uIOYjBfgyVUdDZDMdS4pNGVflhnI1VfShljqHViVVM4idrLQNvsMLeB3FY2/o
TZ9SRWo2g0dxDJcECFJMj6VYL0LyS30m9ab+Bgu4HStHPnHHmkpp8LJFQEuB+u1T
6iKMrlD3NyC3x5diSaBhfWxF6Ls/nueR331vNU35bFLb+d7wmWyER6tSDKIutPYn
inxUDYxIQ6F/RU8A0MXqBz41oBe90/nPJt/M4AwMw+M+1+J/h7RSLD3sit8crE1z
pzSUq8Gvk0fhA6pBNtol3EtdVU0ODUCuXoWxX0KDTvzx8Pp3qCyLCnVwzu6NinjL
0w28BK7A7zxsnStLdXbALyOV/Sw1HjhUfnaaC2QLb1HrYa1j6jkY3zzj3r4DMDLC
VUPp0caalS+pB0ch6d/alynUT+cfwCexsXaZlAtPebg6rwjPB4E7kj0B92yUo6aE
Qvab+/DRfveW6HRtkPAL+uao/COPoMwg7SCHpKx7+0ZcrDykgFPnvvXAz/UacKbt
DKGRdp3D0htPsT1a3jVepl+OtImex0p1hyza0WVBVPnPWg3qrPS66BosNX7bnnas
GyzsFoYBw+nOKcxAbzxr1CHCGd+Y1absG9849njXjL0G0+Moj3mfQHlClLKCaLAX
r6IOVJCJQVFANqFcZpnJmbtDG/novh+IWsNmCuKfO49F8uURTgq3nSkQrG6pQHCm
r4GQkbbLD/fidnv/e8XkglpHrak6FXho2u19Gv5R637EfRKf+M4D6Zj0Bywymz9q
zZnZcuFSwtY8M30gKb2wxpqBulPt4ADbMhILPdio2c/CqQLuxIGYgXIK2AcaLs3N
Lt02qDmD5q63jHzTCQlPNBjzuB0HTAwS7usRQ0phBT159Xc1BPkBtJsOEiAjwOu/
FDVCez3pZErKUO6J6/o4Kxy7JQb5RKFZJpkvJmYGHzDKuZx5T0Z8hcgpoWs3z1Qr
O0RRxeGMwqqb3VR8sIHdQWRqfetodZ4SxJBO0m2KWH3zJ9PorW0embRftWyr5cO1
GzcWiJxV2xkS5As52b+CyW64Zg1BX0XKUFzLGO2LiF6QFE/S9dv0YqP21OX1CMAs
vnHuDYLvTsOXsqysd5I2dm38dHQiZKhfyfpenyedwOiWgyLcj9w0VAKxMc/H8MTQ
IWuLpUrDWLwX40IHAN+TdqIIaRZAkCjnoW9D3xjNC44CAlqfdukNF5wqxNZXA8BI
963w0u8EllRJ3ks4GCcgZwEG2gYUTHXgxMdHps4dSfxWGkFXXzcUUsbF1saa/a7n
N80oI2UuGs818+Y2eeaBloYhlbC7DPHNj4tLOQjbIYOE6AkvV4hNpq33kxaHwecN
4QT0sVuEQLFmUih/MVQ353BdBcGiF6cvkOijnlUzBw8GuAVSEwujV3j4ZEYeDZx6
TLViVO4qdmiKQS/LXiaBkAmCLIYAgLC01yz7APMJkzNxDI95xPQD54IpvugN3Sey
dz+P3CPcPDfbxwxGZGBcSblFUQEPv7aT44gE8BrLBMf7vRhVqvCUIrg5wo6XtOGW
1uh/T0EtZFJGDydQ5/7AlMgeD2yalGtAwAGF6Pi1bTaTe5f99wTR4+60QTVC7mRZ
Y4BXYMcRLXf0uB8EJfijtJxGLqQxF+Vo3Z+UW+vgI+sY4AF0pJvhgkMSMLlbA7DB
+rs/6V78Ifi/p2GWG2N2bsBEJazLXQLLd58Pa3PCXVgb2ElWNFqAFw2+LFPW4aqz
YZMWIZz0+Np2eMi2P6tsrHG10P77T0oCaNHc/KseytcB/dqRCG8dNfcOknAORhdt
by1X7MxZbIg6W2F0BTX9VS4GqkV99nNksDQTmXaQADtbSzTeXLwQWHFymj4JwVfT
oH6BZHZ+Wni/MDRiUwl3YmZOfeo7ApJqwNK6aFGri5KG4zQJ7zlquyRpMm0FFSVN
qi7am4z82XIY1Sj9W5uKrOY7I9PRvn+z7FQiD/mqz+Jephk8oqdPoxqwK+38Muj5
78iLd0DJ+o92Gp5k7TM64CPnHrVen8UUCuJVqhrfjciLrKaSkFnWSKuDyJtzV0mw
85C6YjZ+wwNIFnRMJt8sCUdMgN4TI/QQ6ftwCwzRTpDj7XHGh1w0AHCvxeNcUjlS
tO5sGhyR9FbybZkwD0cf8Sbp/2FgTgoH3/8wLIsh1Y+AlOICeMk5tHc33LPSVbp+
sJEZbmZWE6u/hh8wqhW7nNjpPjSMfzXvvaf3uauTk8eO4tgmYFCSytYM14M/87f+
Xigg/+UjDIoHn5yEKC+7qGzQxhgUTw8Ba3GUHC2cV34T4jtD5KFVCCzn0kc2Pjc6
Eb3MuzA+a3fbaZ0SLSZk4kFr+QyIO/P91bnlLf3ruKZBc2LKcxIr/PLXGg+Qanxc
8Lk4WgtsQiyV+5SVw+yWTO+l3WlD0G/1fCmmy4t87v8U6/ZWDqGTAln2Kh/irHdh
YxG24eAI8wwK70FUZeN6M/gr25VLjDCbNdDPQI4q+tcF9Db/BibyrxOYhKGDD4Ci
vsk3Mh2m6oC+uqRRXiw7STxqx8593Ddvaz7A8/z9YCWzotbZQdKWj1Fly9Srh47T
ek0UDDkk8fbbtwWnGAgqrCostZNVWNK/w4PGUaeNoQVNHB9Qq3znreqS6rTaAewc
crpgB3dDk5qa6MQCcrcHzVDI8c/knzjbEs4lPQtp0wj2D4p0Mng96dqHY9/FN7Ut
xTnU334DL0tbGM6ymdy01sSjIlkXEJ9R4hzurO3iOTDjIC6s0PyjUk9iUN9td1t/
0fB19rmOP7n0+Fi+vWRHFAgEodnRJXVAFukmhS6ArbXSTwAGZopp76WDrBPAqXAe
s2Qp4WGrGhIaSiklq7C0rPFbPjPPEvtU+TvRUXs9Nn8ZgF5VKlq6l8XBU9vfyOV6
R48R8p3Ndgx28vjpFwH46b+hGSY5i96ZNnMK5rPNY09Py8SluxclGI+scjdWuruk
MMQ+YqDW8Tr7xzKbAczXIFFAvenbB6gmbg02MCaEx9dv78KPBwNybzjXS55OKAlJ
NhmZzx3eBvY1E4Gk/QNnPo+t+VGLNWFV+U/YPd4RDuBYBJ2WmVdlcKbwwE/YovIu
gkLv4gxn+CO7f4zBhchggn4mRHq+Rhg2az+xte9+r5UVbksc5HF6ta1MGFbDO8rR
0BS6nLA8wpI4VlE/IULHWFe5uaXplHC/ZTklTyPBGM0KB4bQzvksZs/ENk6l4zGN
lxE/Z17DaYnwd7nPFZQUdTOVDuZ0oGXi0XJCKrQlkSHXtptjWiv9jD3/7Sxp8Znu
eB3GvCDrrY/o0MifWxAYCknizPKXApyZa5krdqIAzgmCy7sRIS8fLWvI8wxp67oB
ZKVRU/vqEgsc5qYGUnW49kdRMlvjw/Xj395O4+VfpPKvdH863Mp9AW+GtCStxhEd
jhykOiTzvqyqncXjnoHb0T0RAg1vvL5TLyg8XJfRW7Ptr9da1FJlAhyJtC9uF/Ms
Du4mDglNaIEydoKdnugU0Vfxyu14uetGltb2iMhYCScWdImLqhxY/3F6W1bENGZh
FeXVRzrUCz6B7J588oINxDdSAXeKnu+UZwPX/j/CZSxK+W2MpyckkiQmMZ1bC7LU
fRLy4Y0wcXDLbBjNkx7q14u6KF2HRPKMeK3em53XUpF3SzKygnxfcoBhvKMRl26A
KRKs8+CXT6r1jDW0ck/a492XMPso4MaAeTrDr8NB212ktRXxDqtmso6t2xXcXVyL
Y06hFSfePcwDSxC7Vzug6FyhEz5i62KLa9zBESB1wE4F33U9Xoht0dbEXVwyCJjT
Uz4fFYdBUBYt4EfUANM7/xxYVt7Txh38wyM919SkMz1xd4pmIXnmbithsnSVAItU
thjCMJQPOpoThbmikWijLl9R1LermQI5hv/46D/ORVBeAcYG64XMkCzfvcX9F8vj
/Ev7l+b6qlyrO1Ku629Kx6SUHl8gB7K01cCUMwijpInYABdHl5RB4+PP2CoSEOGd
rv3w9Yo94vjaVMkLdN8H34A8XTpBrp8WD1TTRMyS37RXf8cH8SZWrgA5RgAC9eI3
eLPULWsNV+eTlN2I9t1CXR61LLFrh0rK7wkK6gKtUkKRP8gDCgax6IA5H1POmAad
Dz7I9tTbJaLvtDdZ4JwZ8j88VNlFoo0YWzwkqbkblqsPog8DXWIVKPdBVtpzx/TC
4fiV66jJdu8DwDz1BWVYtfH0Bx3XSIxI2cH1/9BH1pK6jE5ewcJa7AW0I2l/BVPu
3gYVko5iWs7BWJI9gxqVzB8OhbDqzbu1HYASA2Qew1HHULOUzU3K9m6+7K2JdPHb
D2Oa9foO9mTPi3lf6V0yJRD29LgmX8SgMWRqyJeXRnkltPpRX98VOSOb7YZao4yw
iPSd8th7KSDJvkBkqY2WKk4T4neNO9TnyFH2iZwSBGUNW8SAzfMYcn25xhMactWi
dA/A2IpJqbuTE8+a3Re4LUMyujp+XSCjSnD9QiPAX04kmxmc0Y6+6GQAK9D7ydy1
PDz/YgRpDl9qZdj3ddwXxCiF/cLbTupLUk/Du5nspRuO+zuRiwRS5RziR5HBukkv
ZksMzeAG6y1+n6jTf2EHWxgFpHbY5ia0Ztz6fIfrTXWmBwWCiAQWViApPIMZa7II
42Rxd/JIsSdDvfPnaAJMWFQjg99zdbQdiUz1HWQR0iderVyNK9WTfC19Bf+x/bfz
vVsEVd3rDN5KOpekkg6IBnGxlJT5CDMjASHBVKfWV8MfEOBtwvdbgh1+wjWy/3l+
J0xSqrxVEvxNeaawzfWxkdt+4B4fUhJs5dHiNJ2TfflJu51u+S5u68w6+6N7n6oH
AmSUkpQ7B+GZYMEwtoQPYzOWVAAFwL8Y/GfpOuiPE3w5js8blBlL/mg7txvlEJSg
jfHL6jQGEYgldO8+BC5UYIyoG4iLubVpKn51LdtryzlIc7ctrYqp9N7EmuzsTIBb
lZKY1izMRsKMxp2FG4auSikz/MK6klk3T9aqLA3LqcRtpZrTr+B1SvxbwEH8mL+9
PGwGKjWmjojVGgh7En1IzJWWbvqNJoW1yF51lrP2aQyeEAQRELgKPfdzPQSd0Hi0
2xJZFlwUndgCDlNl5E/WPV9jFyEs+yJj+rQNeiMd1RRFdEfGy+9fzx/Q8N1fCqz4
GXaCcy2N3/sLU88od+jVwFIqAF1gyzMqQq6Lh5ClTRoDY8TdeGLpzl6Jbf2M4VoY
xPm2Y8L+cpQRWkKbPKkK4iwgXb46zOEPB7Lvk1VjU84OinPwcL4YJwbokR7aZIiU
SeIMvMp+W146FwunEEg2gkEkFzHBjBTSkC+TS0HiiqUP3q8y4K48pfIcYqMSmC31
OJnKWFvKIIjExlrPLLFhVUl+e6rE9+uoFLs1OEHNMQRyyZanpm5unjPDj3xy+i1L
49fedPJCkLeVV5Tj0NBjfGUqILoapUxyTmI1hCPSvq4hH7TNokmCE9IQcbcLrEX4
+TMJCZppCRpEoDyPcNhGlmOr08ZnR3C3SDfBYThq732MxAHcmvEzhuGAJTkB9yge
v52QaJZq2lNhwGcEmYe4g0thXETc7Aueto9Mm7eSOOcjh6SHtK5FoptSQYu36OTs
9VcGaGrQV/2xKt96XoijbAJsL2YBoe/eGXcphwlYGuPrwU5Dy3pwlT0IA02oc9vB
QKrYd/4cNe9RPwcOchlAWPT8kID6QHuBjwUVfRisUVfFSnht9SSx9kRKBEBC4LVo
HUq8vTt1HFOzS3wJdKTjrxUvXE7dc1oqoV/tSiXmEE7ipR9OcU9fWXu2CYCDn8CA
yM5EkA140yO3ukUXqOeSMm6WBQNyqTKq/P5Hxw8x7WttmXdY/wMzX+dWubSs4HRt
B+v3oTeTSJYMWCRnVFrErolQgC+M4AD5v7Jd17/zF/IcGI+peXMDHNE+cFhZB8xV
2no+QNHCc2b/C73CvnSFGelzHBJP5NbqySYZCWMsocvjX/sa9np5P+dvdvTTQrj0
rHpouZO7Wi+HqqtpirtHGCItWZZq0A8RbUhM2jeiWnZN+dE/SyMpgzZg7fjqYeXC
6wnut0VCx+pPd1LYGoz389KINLuDbXbjawQn9vz11aOp3Pih6DB06w+8y85f5wM2
fQr5YRv/BYsvbefcYj1ifiqy8SkNFtjgDI19z1cYsWiBdy7tfRtT/autjThfcXX2
bPByzVH6KRUqAJjfBWHb+q9VUZ3lhKsFy+jwvrS3i0mWG3ulH8ZYXvkT5VZcGHCM
UzsABa8aqmkd3jXmVk4jHJLXhKCRQoKFL2of9pnsJ8OSqa9E7qPf/lJP44UWgbzr
DjeUIL1qB65zrt7hLxizrHZWJPZ22R1Ul9c7xT/8bdD9bYTdw5UDqtB6ciT4rA5f
FQDjKjEpx+595BvuPXC5/4dJtO1Ik/5FLQpZQUfx7ovD3v5JRlxrk6AJAovyxYfo
QOWML3FWdSCuwCfoxSWW8yPvotALZHPEmmKxyyUJGG+jj2zCI6rP/jZDY8voY+eC
Rzhp5p4Ra+zk2c1C3/H3btaFgLF/CjMjoNg+ZLvcr3MVY3dSB2dPbnf2QOVTObdb
9xp0qAzz0yTy4Cr9W+spia3mVDmOkFuNnW+wGh9jBdg0HRbqJcK56lJ0ReKjz4Op
k02u7wkFBisaz9pSAmsxKUAKfSzV7ulL0X5locy524jPZ1wKcTnS74UbCFs2VLpy
I+m/vaNZeljLu+NNmbFWRrnwoEaaQcZjF+SWwDynegwIPwr+V/KUxvREJDqc34Er
0Jcu5pPpm8sJ3DjYPVRHT6qquqNkoHFPFuLz7gU9fkAEego9mo4WQmMH1TIjO17Y
mpS3Oq38At0yjgmLA65FB24NtbSv4jKOnfY6DJkohsNbFW1vfgQbotN6DZXkOzRv
tUDJtP2g4O6pENUpWWLJGzD2siauPLHOpHgDgMS/7go9xJhwBy1iHSMiRQtcLBPs
ckHJwVjuO7KWx2Hd3prvz0CXyfJPRos/sa30B29WAy4/MNJJVaCR7i4gbL0Lh/IE
fD/QDMUHu0ZxgWqhKQ4m8DCOZYR9SIvxKNQnAXhr2LpmhIEaoDhywZwKbGU/Nq/+
tWElLBqGG0XL/cFvpmPQXsK3Kg3q7P7OInmVzzC1plHsa3LHO6jle5QSil2giuyO
doNzfjn2evfqR3qXeajy4LFIhNTNWAJpxXeVY61wwMwq4hO7dPqcUNFyneAyr0aR
ScVCiXlVZ9VYVjFATUd80UkLo3M7Cxyhg8eu8MZcn2Rs/Z8rMMgz7YDvU43PhTlk
GNn+ncl+et0RxzvT2KwRFsL2JbdFbkLjyZ98jx3axYSI24ckkaPrUtDB8b1uyQUB
SZI5u8xHd5UTZC6rFzf7ryu38mznSMatinl21zZ+DnACqdPCFnpDyx/rajZZOsIj
axGfKz/sKqhApqjONWOedSVb4kELDFUAQulTGa0t5kRKDaFlbpwPPJGifjMEQt1X
yqVFNkoUUWWALxhuQ7F7FDrEzyxI7k025CVWQo9socxinMDiyLehUyD/xy870DTS
YhZLdCAHLfaUVi+TdqRNYumq5WnlaGVKdAUA25lnohuszNb3m2WxCy3YiFRwq10f
nYSZ/q8Ip98o9q3XF6HrI428BRp/39/8uvdMgqr9HEaK/CEDac4SE1A5jJDZUfJ7
ChvcfGLQpv1cC81xgtZtWRIginPsZEEp+S+7thTHTyyp0R2Oxe2ZrM+Rban5djSD
+cNbhMi9TdcLVLpBon9NPdvukQFs54FyBbLfkVNniSrob6hj433FOmEke2jox+kj
XOf1ggIerq8nC3XLI09Ru6w+mNe+DXPFViID1E15hYWEDm1gXcWZWCFMnm2nl5+h
afaiV1Sc1844sflN+satBPez7nk5bTE/KASGJU3gesO9kZ9AXEyqmYZ+G5tezHL9
jXMAUpY6LUgHlauJq+7sXEY2NbtuAz08Q4V9Yq7NOMnMojpgiUOUbdkvS1RgeJV+
o5LSh6C7G3R0xaNrMc/+cT8kbo/aEzgk0thIdkwyGGPCdc/PYtvpAu5TdHwrsrmj
v+zKlbfL8pa6/ZOn52VKUHa17+ROJFhgSaZSxDmDdyQhc/KdqiHWNWLUxtB9E/el
BDdO8RtLdHtqN3QNUB5BYTDxtXkiLs/18EyrkLyoOFWUpEwz+a7P3slNyzcs3fD0
YmUeQosau30WCe+JH4HCoZDR95maBtoFyFw1l6khcNtZIbejo2MqqhcdZONvciXL
U8HfxjzPpce6I9DzAezUpbohPu2T70zafJ95CfbRuXqLXHhk+LNgGHigLGbTyJXu
RmT5cAaF+3a9cfCp6LdP/hGeUtN5z6hutT8nyOu5Tr/VhqIVP0nIhRerpLDYMACX
5NRqOOOT8EJj1+Og3T74CHRUmZpzzyHLQnTVdNvhqr+hXIlgoG1MWTvSI+KEdYab
SMXyCNnvrKGude5OHPQxNeS26+u3hpruPoJh8AIiDJsykZNgzVHHqlQVtzQS84tx
qY4JJmEqPoWON338k3oTE8V/Ige26xq1pUR5arrjuPS5uYZcsrnVK5T1WJ1NOx/h
FgnidsiTxNa8WRgZg+tzmrFhuuHNHcHNtX0OHnwp6VLefe7hHb55QkjQV8nap9Km
P3WsYHfzgpZlhriiwxU1LoRMgS1oMo6Xm17EC9FlQHXrmXTEWSFgOFAS8jtlBPqt
/ocBYm7CbCNeBxwZXM0Sd/HuOFeYx8uMACqQQ7bVcZGq3lYgo2pU91uxPM6XeMV4
+sFTdRH0s5JBnBViGS1rnQiur2IhdAD/uuuZYiL5LSx3XkcRz02ly2OaiMcyW8kH
4hN4XQ1iEEQ0s14UzaUTjQXGE2yjkLO6R9SdV2VDVuLzbrR4XeuA5+qWvJ+LrGvU
UHvMlKPJQ7CpqurUgVIJurL8dbuAsXjrQcrHhQtfesfWq1nN+h84Svdaj06k8Se8
E0X4EghxZtk9HZ5kogkMDgha00KzRMQcPL2srJ4H7AheF+mDOE87b3Z+yAsr5HEQ
QMAZ/z2yPtLXhm2dEeZfgAWEIRZVKeyieb15VTPjr9JJ/dHU71ZE+kAnV00puhLt
n6oIyTTPkKfGtQl0C/UMFXljKVC+SVdPnJgC+aGMPSvCddmcyhBPEuGKjcQ/Nn/w
SbnIELwbnhK3A8bOrTZaJM87Hgm+pqjKIpTePwHb66y3qXT14akXkVjgDDFnyNoT
FdUpnQDOx6VlkyFvjXanuZYY+oZdBLv6bJcW1eYsxfbXRCYdykScPaol2h9ToeN9
jjuN1URp81XH1LXi9tGUqyjjurK/31FGaF2xbFXdu24++zhVRZPE12RHiD9YxI3V
KEmmXv0lwlzl35q26JUv2v3rXVAclTQUa437afXPiJ6zOJz9K5/PJuBTd39NjSHZ
7fqxJsMYcR3vY68timVGC4QaWtkZDN4lux9ILx44j9qiIY2ilPLF38IzUGO7fVYL
phbOtOIEGWlwOAh9gLsBozU+fi92WJQ1AJ2rl5B5bAAao3hrM4fWcKevSR4wFWjg
eVk7/U0Heb40Y9PpKPvo5aYGJ1D5IfY+ajSHlbJIcIG2R8OozgvYRtZ1wrmAapD2
Hf70peYNoDDymiV87I45Tyg8Z/OLF2yPXCbBeLvt/qK60Mb5z4XH93lYj6DHiE5W
b/H7QiSWrQ8Mg2s+NFR8wzl2TGIqFvI5en7zZI4bm0SWMehT4x2BmuuKEztcVUe+
bNa0gmvMXtnUaQXfK2B0C1LcLLlfyPNG3mfj3vT0Z0Jc01YE3NRpIyuh81TY1aBP
VpQv/bJKIjwRwRzVc3D1fKLbXMbCHHiFjZIT48Z1X5j4KTWbtyjhVXD+5dwjOsTi
D5Yql82QAfKVOqKXDqjphqj6GcybjHgpsiniASYaGrKBCaP+00sf40h15EsKF/Wc
YrUB9y6HxGwf7Ji9Jk4I16AUEsa3Ei4e4HwahWRr/och++V0i7IGTJWtQRUESLo+
xM0XP0fOpOShm4PssrBswBmo7V9LGvwonlIjjUwRrX5PbAajnYSqN9Wlh7iV5jeH
En7H9+fRV26xF/Bs4qFtv6jJPE7UZgdvlltX5REYIa1Mv5UqD0LizrppJsvbr3U9
0TiovSPpG4ZBJmSpplTOTo3+Apxg0rzNPcpDNgWTBsWqdyklz3P/KShc7kkZ2ZRo
rQFF1sDI7CgyIhgS3JDRYKy5KpfuSiWnXu8/b6EowcyhVefrMHrsv9Nv8iMBDeZl
hl6h6fT/evvmFzEQ5rqJpVL8CdA4/Z2BMWOYanw9UGzDCwYyu4UZI5goXOscfdoC
CKtswmGVjApfWDS+RJGeITGxf8kwTQ3r8tigr/JAFizo5XniFtJgpuwrQNlxU0qm
EwKDo+w4XSp3tP2U4+bc/diR9qqd75yp3IBx4trybNVxj2ccnOnXFad+znzdW4OY
WHcZizi6UnfPxWJt2gmIby9yD/VLZbOBZOpIlZwpOXhchxrR1pm1cLSH3x/Mb0N5
fX9PKiMwZ7+KAvgE7Jg/qF5130C/D28EaZUw/QpXqGRQTBlKUUyFZ4jhML3ccvEN
cz/Scj5vKK1Wz92J4cmqUZQMP6p71I97aYBKBbFbK2LKPA9E/jAmbjbqzUVT7hPx
sMUqlI2Q99A7DFZrpmWkIU3fTKspGgIuaJ4P85WJtO+Z5GHmn9BwLntQfl+6p6q1
vnp9XHYqDK8CwkBsScEAlPy9pLnG4woO1F47+axqKjEV6zPBrAQmR+DpKE+GhCrs
aEBvQaRJR0p8V4mTJeIYMFw252M0tZ9m+mHc8jPyAPJzQubdTj4vbR5S0Zn+idpv
X8y1hNj2jFxupbTiTnZ26dkd5k3zmMwEkin5WS+8gAn7VCKQOYT3XJRqrmQG/WHW
EQTuLubXRrD88aipup547Gr/K8UX4mv7OFvdHk28SvB3xt7irXWRiooTgvt63XO1
pSlctZ7IqjIBXelluNEjmK0C/qpBBQawlxJqcT16cL/3qicAwJuQJ6MLuls9TdzH
9TArDogxJLUMLAE8ZUNW2a1S3C7sGCQZANBArj0z6lxA3mJurAnwL4FzF19NYfc/
XiQ/ocHUIzO/y0mKYYEyV40gfuUPiq45btGlEarRymX70VxqQyiH9jwykzazyaoJ
EYfZRzLp6rDraTBu8c2S8M4deOjEpdvhIzinDClFuFgdKMXIQlQbZXjxDtaJJJur
3Ultka1437N4uBSPKGQv5JnQ6a6nLMoPrS9EwYy89Z98QahKt6iip/2ZQlKAAsuQ
vb7abFimhtYFp/V2ol8oLwAmhHcvLXsbz/f4pppqPEVL47G/o6lNJt71qn/9e/Cu
eWL13Ec53AFwAcNRQnlXSRQspFIXkn1qYZhgTbcHyY7s+xavlyv/UsqJlCdyEww0
Pz3kk3S9P2dG1CEfG5ebmZ+cBrdDds4ujo5KFtOvg8zdqqMxgNwC8bwgRCz3uSWz
8qmcP5EyCCWOJkncCgM09s95z417y5F/SYtjFZVSOpOZOaS0iokTnt6bJXZuLn8v
I+5TEDaqf//X7blT1ZNsdIMZZ2cy+ugCnP1B0srnBqPN4yYYqRoIDagFgnCwabtT
NGCy3h9IVIegEN8N5LxnIOiyV89fKVVSoCY+MZ0REqXKqOqAmVKDjkh/mB7UAkko
xSMUOv4ik8bRjkMd9t18tbvfUyJhuu1eL6g0yhDEJJJM2+YBTmJd/RBRg9E/p7oV
i81HBovEjw/Qdlfehox14Eq4Pgvc/sB7G/sA3ejqZmXBxVJUKiif2IsB++6ymrj5
mydrAuwFYnPWf6i2Ynj7mDp8azHHHzEdaKF0NRoY2m87YkuO+9JyQq3NECY4t+NW
A/prg2y/A34rig6p66YIbYdP8i56LgRiAf7L/GQT3aAG4Es6uqdKqBAAAzANjyhc
qu+9EcWncuL3RCbcz3eArV0M46lxBTUOvrh5bbe103lxd5mH9BChINibnVCZFslu
unlm5CTJJPQN6141uvm2alnCcvIwXQw8nG4T9g7EQrlS7BteqxwtiGCRXYKtaDu/
CiqBpVcawPHm3KjudGbejtXIty1fgPhNt0axKnNw1p7/5NSkbCkg+xzGM7Ji0RH2
4dVuHJK5VyH1dzQ37fd/q2203SGC1acOqO52+TMbyjVms/43lAxWTouHLaSo0e+3
kiOk/Pur+IzRp13q3W/SjuQQyj3iFF+CaR9K7l+72MBQXmTXKmKa2csg7WSwOAuv
IlGybDSLSaf/uK61vSTszUDhFAhvPDXjgDnEVPhyohw+u+h1iHOXjFoA+uxPPMsT
OQv/RrnHd7VgJWJQc+kVwGp/7u3P5pJG9nKvar6zNze7iIv0NW1xoxIBxuT41znq
4IjGneD/GERre4/eR5W6pSEWwh0SiUNLomE3pEkdhqDh+fj3oIE59ahtoU61M72C
pcEYqmzqXUaRYros70ys0sfIOeKJTYBj8BsV7WiWm0HmgTroMCI/DWI2RRva7lTg
urdWov2QvMgtO0StRX2fkxVecHTNBYTDor5eaNsFTZ41+aLieGkYBTuT7VYBWxbU
DIF0i5hdNJfVT8vYCrApdQ18SBw3x50a3NxhuNEPszjzDMu8Mk6NPLRMNsx7VAxt
7GMot0OCfyun7lM1E6AXOs8RYxRtoCR1rjsDDDWIsqYXAx15KL/oglTSTczViHGR
w/cr0J8J2x+u12nxmTawnIiwjeFi9Xoy1FJcTmliwvTFytz5cL/bn039Q+k4XQuE
DzY9rOWYn9X7i8YOqxXCamqXyKyIvdnaMvJNh5Qpd3odq2xbLXFV8reUSqWfN67s
4OWU5UQAKoRXMU469Rj98dPFLkwV9m9L0CqMv49m51xn9Y7gMhxhGxHi4acpYEcg
di6ypARq4fVxr6I5nbZPjoU7yg0QQUrxWQhgb8/Sce9G7jCV4S7rc0XBKf132HAe
gztVf9n3kGTWDqijygw03uVa9JQYLAmjWhgJPnLWZmU7N6Osp3+ltkC1+9omiuSz
HiVdU6mX8UmvyYokzVJV59Z4UWEC+dHAss5nFPDXADRL9R3q31r7qQgBblEqPP6m
Nh/YnJvUewqTxecXSoOzB5QhIUYT4DuyAfEzcOKK+9sAiMWuczxsAbOY1vzC2dTH
TY5/6UtoK5vf8wQf6yfkoJyenyBgIgdt0KzOwfwnaykxaMpeXNjZyd3J3AXqclvm
TbXHlFM5XtsFIfukety4QvVr7X6GBd9cjevssJeUr2iBmO8KeNjGEod2hAJc1ZsX
ggoBRBPLAMvk0MuBMNonJsXCOSb47hzUwqVZuRGpTMq1upUSUWWecuC8n9aVnwr2
BaQVjjk0jnTjHbcsaMJ7g6fTHU5BfzocPn23LbC3zYftKpzxyQc8AgNwhSW0+ILS
Irw5YEvdemKi67HiMFhtPIuRuMUCezhukMJJVklHS8QSaVwIw1EcjZa5kf1fxnoW
XpH8Qy7iYwazZjzabCJJpOaZiY76WPJvuBMS5lxABSNBrIh4SDAiCgnOoBCMabCp
P0iZbdjQP37+Axu6d5kheCxKBjw+dpiRSAVzrMf1RENBvstx23CQvwlO6x2b/I3L
RGZdu/zluwyuqK5puRss+I3V54kBuhQMPeAK3IJsbPdP1cvaWtyRYfInpXY8eXmw
0nUgiTBT3webBmnp3lWlf/t0Il8d/PHNSaN3QkJkcwbR/ZlIuiaO/s+yMVCyGhVy
DteMIhFRrlz9a+1v7ew2p3e3TMNvePx5GSC7ANOXC0NaAV7kMrRqFrOcrAsfhsIJ
DTmOpusqBdJNtYk9AwRDh5Z0KumQFW0EpX1ur5lqF0JCO2sYQif2QvvvbDrBsnPK
oB6baAzwg6lkjj8eFOXsCv3UBnsnd19MGCMRpEYJYWuiP37i6RvNvTdC8NSULVBa
t5Jj3fIFz0kIiQnwmc1sXI+E/XdaOkEADQTjloOGoZFCHF0Pw91B/PwHD9yCQVfr
2nwewSvej4Jh3m4lT7LsJiepBLHy/GFIpsVy2OKybBBsjLRmj4b5ollkSaplnR6l
VRHhauin8i4/U6EtocKGgvdrX373ttm7QCYHI8AD1zBa+4D75Sa/1mRdnewsn4vk
WF7AmmsoRo9XD1tnSOkvEAQ5BT6rFy2RNQnNEDPIlYe3/a+Ef30MVA9m37joNPXR
IDj49UXeerie70ughklV5Lk8336HJndqRSL876OorioM8qhMhqfg02403+3qE3nq
F2Gsb9QZqUrfamcJMltE12OnUI3+j5dkM3lPAYTSgs4GC9wmEPLe7qfKSX39o+a+
eBp9DQAP9UX6WKidglgkbunAx3wVZKmcnSnmmuzmBcUqDm/5XQqQCD8cjxVRhs94
v/iTif6kP7nLVfiYKFy68wIXfUsgBSA6+aqwdSfIO4iZZgKsmT+T5vkBY/3A161R
ZeCEqLCNSVnYhiNzG/g03YpkqOi/0ZQ8zdOir6w5jXb/Ih7c6WOdzfVI6JewZxPQ
dufWvrBCa7XO8BXx5lA/w4lnbzGheoOP8v6T856mC1dEGMfcHotdiseIhfy6Xy4G
zHHU2oGr8VByBlT9fuZrgMKOj72DbKqR1DKCIrPuZSbCdQ1Cb4DtdAbYQsHcN3VN
v+pZjf/Wc11RH7R3VUCnwhU8+O/i2r2v/83cEB1y10vNtrtFPRY3zPGpa/pYvHha
mfLDybJSYfKm0CENV039FkgdZs7WtnT6BSpqggM96T+oPhZdyMeHzvznyJT1rSi7
HVDbqb65VqLThW4OwWxVngKeBsTrWg7O8PbSOtmxaLoJ5u/Xddn7ynbv2JJCzW72
iyIglMhQY/zyFF/BhZ1odFsttumorFiHsZRpYIcUTRrr4Dg7/iuDI2LkfT7S4Yr5
Gl+fzgmF33oTr/6TPfGcLmQEr8fQiGcfW3Id7BxrmuIntpDPGRI/BuRvYNsFitPL
FJlPocMqS2n99kxL41vojk1AkgaKDXMAEN0CtPRqoazDUyZ+7D5n56VbUmk6yGYd
YIfDrXEYnaQr3w06wezlRwHSMzFZy/jbP2O9YypOnRmohzefDnQHhzGOFoySIWjV
HWG7n1CwFjEYNRQuThVnt2qRmPoLgNAOxhNAmwvu/GEBzDgDNIuYC1NuYhikUGAZ
Q9wkvhJa9eJ4JWZ1f11OtoG1aE8Cvwu8q5fTHkGqADWdLASjltlwcGvCx5jE0bXc
Jh3uPTa9QUgpmDq1jKM512mJnEY8Ebs3DEfo8BKG13Za3dWNzZ8fEpAddpYZq6oa
HU3EVd4fngqUqGWk7GVS6J2a4S+UBWB3bsdIOVCeSSC8Roi/l8d8DwnqwU/NDhIC
zfyXIBVleM6U51y5B/z3y+TRdmfdGlnGa2Emt7L2P9kRXrFFdg0JtWeMTQColHKj
Xnjz91T9C03V2W6ciKXXuNEhqZ71wbDhwZAwk4MF3GxIPxaup4O7C6XBU7NtNE+b
AER/TKGxQ8WS8MvEvgKOy0VAqx+10uzgNrbenCRdKqieeM/Qn3oX9dPdegq86gcE
6n2EdL+Ihj3ONb/I+Dncq4J+UZAYKE7mvQ7fiksZWTfz5dVnhoG8iNsZacJJ3XTh
9ZzRkwVnYjFXw71ejQE4RC0hrlFvAjzYYZZlNbj3aLAg/DkNOmqaCy8b8y0t3r6t
A0uktkbiJMrUOmIUE/tB0P2H2+1ZOVeS3YUs4v+joBBrEVHVVIjRALNbuPSWfwgS
qClCWWYgRXhxbWY8fBK9wkKsYJVAY5Y8zFmzs0zUsQyZpdN73zdcHHa12i83aslu
9ktSLIDFlFZZyye9+qFu2tHbTXT7gzauvF8z0vl5Wt8hV7YGoWDlzs3+GmDd7SGa
vVOqkzUxjQ8Mxy4tOxzl3XCrfpY1MJK/1zNWK7RTOPUYhB5NPt/OJg0BsmBTNIxp
vUYKnCPmKu0vBdtSGwNmmout18EEPwxId/q9qpxQcyrHmMrPxYOwIhsaqrOSy8lV
jSD91VUOhHWcOeGg2aJHHxVtu51zIWUkx6IFYDnWd2jv9gZOQFCh6BJOzlwYFqz6
Jz5FwHdpeU94NWkMQNdByZA4ZbvO+3oL98oFdkrboMyePe8aSxfXTMU5CadHAew3
GonpcKvcvWkuUIN1rUMVDgsWW5ypusBydLxN9ylvMmEHBq7ISf7aHUIFr0kQpw54
rtGbNzcVn6Cva80b8Xny2aR0LXkECyiSViU5xByDWGLohpweKzVRzlvct+FQ6bo4
Kc2fvtM3fVvCtMqZTtFexbowBhj5almhtYPUECl+b6EQJF6mtg40o+YCB8XioAs0
M3xFAzdL/n3By/Di1PUVmnfdqzXXRCl5PgfDUbFcR0kJ/GFOxSwf80NP+SZNJjQ7
2IU+CWW+S6KXFIwivd1alAZwUIXODLnYrv+fxR9ah8vYqiJRco6+E9NxJrmw7eaX
hr2dOBwc5hG01wmNXkEtzURL0PH4nWn0BPW22qiOLcfd1ZtYoElYVbNW478QnThE
/CtXaEW2jruTJ8LFft3b4xkjRwpzeH1hjf/G2IAcbMUsW3Ns6++eeakGH73Vhwu5
rWDGXjcJYNEw21O6iPCStSW0/MBqLi4C1FnHUlgQvysC1SajUJaC+QZN2vU2NRUu
uSlaKtgKTFvjSZxypHzXXAYuusLIeL0Nd3+qD1WNEZClPRlnDu1b5UPuTGPJO2oM
PeK53Csvq3Mqui0yPbBOuxpuJvSJ5CSTA8tfYONhhXZ/B4meDpvzyKuHCI6FNYFw
WrYi8jW6yoKVmNvaezG4UUKnU13QdAllg/UglqnAzj0AleZxQjCmv1Fb/VYN/IH6
varzh8NN39fsdENbXqFhVW5pKYDLCgZx2O7jRbQqEg3hF/niCdunUQ6Yronid/hN
wmjtfdalwTUsf3Ci+Mm54faZFEePs0cnnh7+Sz1jLzL94YVAnLgmRpz9+zllIC6j
HjA0w0VX3X+Jej26iRtF1CEdRvv00QMsGXzKYKcXJDXKpBF9K0FU6MyUhF5veh19
rxZiwlUXLR3lGLlOQWP57HNjpdeBH2H31EAf0mqPeEK13h7ejBNLM0P53Z3bAqrQ
txMuzL9O+VZSjrDZMnTAt4gZMEDTILjIkAaWDIfMWgf8klxFzsRz5VqHKilUrKed
TfCyoaQy3hfAcD0tyaBCUqyKtDbAeMpjXZUt3DQ7XxoVH04GlyXwfsiUC15zBZF/
3ZaG3OjnjcOs0UwZWBbfSkg8f982rJ9plh1JnPBURN8NPVEFeNfL9H3gUtn7OCTl
LRV6T6TMdADD8SyCAPr1Fa+7hurW9Yc4syAc0vdaM4mVCEw5NCdBOhGX43lBOEl7
jy/1XqmwKW7PV24VzKNiEbeSdZSsEm3VIpuUI95ebmfaIee/zwqkoz2vvJNTIo3j
Kdju1AvFS20oB0nM9K0JGT/R5+M8BN8ewsBiWDNAuPVTYdA5bvevxUr+W8Sju3Q9
JXoVIutstzVaLYWo54nQDFGhe4IytWa3//d5qjK4co6zEgd0ZnvTEkYTmfuCqAtX
gk2J3K5TfJL3LQYQFOiujkpqDNGrG9LDUlCZErRATjhJM1qFaFHrj0D67LiGJ5Ip
Q4mTBQoCP9s7v3yk7lZRGJbqgRPh6LnIspX3woGfbigfrLJ0/HzlPcLWUt/ZY+Uv
4yLHsfPbHMpne6MlRInCZ+5RfJndVe57FR4mAOTfufY07nhQ4tS4QdfjUS++ozp2
HLnyXUjnfsxNBpfM1yexG43PAyU779Dm8DvLGzZjYeOIQBzGkB/Xoq5EpgAEyhvm
e371azUyLPXkNN/fvS4eTr6pQwLshG6jEJdHqcQYq3LibdNQHeqAnA+TO/JZ73mD
faK3vn5DEpZRroyQu9Q3aWFuK2aKTW832ShCaJN/7728CzvzMU+JfYGet9kInG3V
FWAUQ7ZfFgD/CLND5UhYouKXzpIf+f+wxnZvw8W5nay/l1U9wG1AFPPpzcaQdbmv
VRE5jNRx8FgSrd07I0l4IFN7WINHodi0Il+0QUatsS9KCICS5CE7NPDhGYGRRRDa
++tOnSoCYWuEfrf4cZUFnQkoko/54WgCX8ol6QvgrLRvK82qhFlMfNakU9GQpAXO
ZgAhHBIutfbk1JzIRFKlfkv5p85ukDX5wPjlndxD+l5DWVMwUuBaOdZZOQAPZfl/
3qe5UrE9uU6DAUU94wKAqKo5KJnflZdz5P/LlPGAjqW7udrfujKZ6PkSAaOHNKqt
xyDnV0wXxJfSLQB8OhdAklKiopEd7i/8NfenKOmG6eFknMWTALJejZObNp+No2hV
mFlA2Cg3XcufyxvzQMNJyspR47qBy3htpSUxcnAcfxgLCyA/q5gt1msA0SJU3MqI
jTImeioBYDujFp9cdZCibhCxB/j6Lk+fWGaXUMMqxtoySxVPBZxxTZhjRz0ySWel
RLJaDSXJAlbOdplIb448gTpYaQ7Tw4VX3aDWmJLaH/Eg+/2Zj/Mh1s/5663m4qAh
ctozt0NP3dnFnCFIE4oLw/9g2OzV8N9sLHUHaZ0cj7lzZQFIMvhoi+H/ig7dpq7k
Bl/8Suyc/Q8568kAoUTm47+dHtBKP4Y5gUTmQCa1oJw/9ZBU2UhMmHhmXeRtdKfI
SGZ/PBMIsQTFN7J6UHK+rq3PAfnC6dDPb5CSe20vEBLJCbjJ7h1X5Xuapm8sHPbd
l4RbsLtckwocqyQFYRtpDO6Yob3HZrnKsgu7nFMOnlbMhB6z8Pc9YcsDzkIPn1wv
uJYbeP7qeB7uHTxGpfxS2qZ4XXYRWe/SPZ8+wz3WZouRgDZ3JMH56QytDNmzckoa
H6BibKrjsOJdLUzwTS8/goANwc92QWYhUGAf1RdQu9bET8aneS+Br3ccg+gv70kM
eA+ZECw218gBiQQzXq/1Vh8aTPkOpHAlsQqD9L5fIKjiEiGZ4yit8JZNZoYB9wGJ
P3H5v945L6+tQu62ECm9P6w8RxirB0XqS38NVIX63vkG25KsxMkpyqrpwgt9/Bhj
sh7CqDBJVZgqf9IC+fDdyuMCEBLaxmDi6xlUWLp9yeLl7QgTAPlZJlb2k8Q+j+1g
2cHqGaqNrp3rIgGmdaJDTxd6zFz9Vr8tmVQKiQKNVCNJaYayQirnYxIF2+TYl7mf
BHSWyZs7ywrrCd/jUmLXonPInum1yOjOYht56LZbJONs+MauBzDqzhQ+rAIfTVyA
wG/0Uwqj0k1KBpFWde7nbOX8xiKqWHBm0EIDL1frVz8wm2iRJIyvP0JRjSYCjsfL
OOdN7UKbQ4h6mXk8yXqP8wfUsHxq+qgvohz2W99tRZR5PhbAHtBQwvshQhh3C5Oz
k/KyNeg+XrVvfkvwQhwAM56rGO/KrK6U/SkusgWD165eL7FdKmdVXAYKGy3t8sgb
IvPhcF4cEYehERFkiz5o95t8JZM+fYEDVRS0TKNPHkTBdfWK5XYg0/L/bkCMkDFo
USPFIkWNpcprSASeUFSiDJWm/48FYS37QlwewtEFZ+0wXkFD/jIRAFpMl1dROdzt
915vYsM70kMENkRAU0zWlWTAviBXcljyfqbN7NSiCy/yDt/H3K37EdZBLTSDWD7R
G9blJD3YuZXnxtHumAKEwigK2SMFMU0mWCKOtlyQET+IFvNGbx6GOUkAvjWaUJwK
wzw1xzJeKl69wSAY8Jwlskddz2BDN3pSVg8V8id7mSoDLuUxIPubxRBwMoakmE+8
4Sdsz50iRws+D7BEHkzCxBW7fdS6uT3RgMB3CNOyaDYMYPcwMtwjqi2D8qW/QBra
ueMsCGItRKSGcJnTr8aeXgYj1hwIb8OdU2uAwSov57oVqtR3pQzbZqyqXHJoVFMh
AmHPkRFRMmlD4Ue2GrLhA2RYprnFz8MYLL3WGKyxOqI7Vi7KjQHLWBg56DMpYgOr
Q+nCfjFBJk8krZLVBkwLMDc/wydF9x5+beqAt3yCd+N+syfMgPRV3sG7hxzSEJZf
vg+jkZURlCuOLOr8TZXeCovpXcOTIADqo5GZu3+rgdbhTyqoSWeIczlSfshIbFiI
bIVH136SXtfhYSSFmlOOGNEjV1ZIEbAuVqCP6radSc22PhqUtXJFfNqYTOUhemF9
wP+z3c74v24G8DTI0AXLDsa32lmY/Ftoq6AtMk8DLSjlcZbAa8YkOjcNYwQZzIf3
tx0QifOczqiFXA2fxAJ40Opd6AV3CTNAcAojBfxZhJ1+siYwpN08abQgt9z+Mawb
EdPgOaYfzPi2M5lp2dHojr5TCD2csrKovJ/cPYeOyfXucZNLNFNPvm5UIn+rrwYr
zA76Qa/cyyQf+rrldskW8HrXYxHzLXGqynHnl8EBQ6WmJkoHYkiPetV9yaoQPsYk
dwZqZujKKTuZHeQLFDngrMqRoVMokvyN5KebbRdErJQ50L0KFDBVjmrB8CYxYHiO
iec4sStxjIeAWiAbhjiCPWnCOtp0ND1L8gl/DyfUQY7g+bSQ+Rk3D/8pbEAww9C0
ysl3/FgAMux/YRhMO8cvNsrIocrao2GPtjkCR3GjyfpGt6l19JJg+AhGh5TbdPAb
Bp7BMdyu4BSEfqNJ6fIhhld+pW8rj+TZdojVJvvweotU5bbjbagOqHdu+cE1dDqS
yKGUbNhcLwUJfQ7iyiSen2M1QBJ5kQA6tH9y6fKbNfllXi/TNLKa0NKs01G2/e/u
pL3sPf/ixbj8eRlm1TAD+BsYZxKtVZe8FhaPAfLFq3ou5MnOIpqWGFiAr00/isgc
xlYaqXQiFWwMSUyYuxgSuf+eub0spP9/HMger8sza5ocpvbuWJFG/8cRgAaj4ilH
WpD2B/zR14lJDKL52awfharTq2fWUGHKluxI49ns4Oe1LnBWgjjDl/kTZhcZ14QE
a/OdwAMW8H1RxKtEl5l4xLNaqF2OuDKOO/utfbp3sg/Yz95tMsV6FgrtIvR+MU9L
TodXpxV2whDuz8N+t/+T51MyxTcNfzonioKnQBlXwwpok5w7VdHATCKZSNCvBft9
WoGLIw9jf5bIZJ0+T6+3RLPdkbHB1hNUZsTWWGS5vjJeX0rvs3ldors8I5NtupwY
PfKjKsOEbFAMoJC6eR3NO0oIGHWLjuTleQMRiNab/YscGTj+IV9Gx0sZsUf0ubxc
mOVozX39rItBMvmd9NP2r5RBm6/kLyPamH874BtHiofFwM/RiXtYvpyXb96R/VR1
s8meE2kwkTuG4lw/94PeiupY3/sQOJFFAYImVMHjRSDl2nWtYGP1VJyQhHU80s9L
Lk+UeCUopD2jjWFmKtHHNW2r3bJrVWxT18X/3nBUx1s4GYWI/QPGqrGLGGLc07Tb
oa+y7N9kbJIvIU6Kk9MWdPDhGhblM6NecRf3t8xsanJHMJ1xIqefI074EUr4iE5o
Ef/6pBXDNsXTThVz1BWFg2OvvlPYtBtOprDfmpiTIRAzLGc+ylXvS7PFj6IYv+i1
iY59kB/k3eJg4z8QBY7KG4Q57FkDXI7qJYw2zmnaRUIkQ5LziM2HQsuzuaS2qNCY
G3dhKV9EEkhvD6KGyQQ/v6GdsLlFoC1MPIlQbGaDJapKxfUozNQZ2uChzyk9I/96
i/WMMTAqy7jNNA57Plom6zQmvgiZqQn+Q9vKZaTdERIZaNghpfK5DKHi12uAAndA
5a3kEBm8M2X1RmafE9seLNqYUXvObvRVSDnDDOKkCr0qNRRVBvVvqLsTFhAyRXVr
ASBGP2Mjz+CCRfNJrgMEukSRkzMLpzYsV8XEdy1u6fDbhFNEh/MGVSYg52wDbapF
9k9W74osoeKb067NLpBgzeIiPzap/USyuM8JjBmzrAg7hEdXRl2ZO6QxmztEGTYi
ZI8+6QA38liLv9EH8hqQMmUP+hW00UKN8yqN1HCPW05LDtqCBn0Ni/5+VhnGYxXo
ULPU6wK9SAGaiBVVVq8rVb9OHhvF4H3THHhdPLy3oVwrSkiQp5rvE1kgouDScLHE
`protect END_PROTECTED
