`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oj6yHHuqYlcm89yhrzFume8Cn0bfQ2HIyau8w5/WfH9deeScEM4Ytx0b0TTtKCa9
kZER5sPomYh20LQbWN10HnbeyHeIyv9DJbGKh/lX8axbUFfOqOs8nGhm1NEtQNRd
wb1PZjdevFEISqfPWCwdfX430HfVxC6F22T7KGqdChnc7nXVfqD6padvwSPrSVuU
J5p2vNdooYBTg6YEr/U7EImsIzVf3Ws02z/i/7zf2kZH/m8khf/WkOTeunpvpXsN
yXgL0X693geLTeUdaqWeiLCNZg+9OoKV1A5mZ2XcnnBAOO8ZQkYczdQa2LqQTC3Q
N6wcXYmxfXi8ZJk36l88+tTHpRVZQADAlkfmgfXgKd+5JITNhHSX/tt6pLIxTdWw
+4DkucH3Ni03QnS6OYyN1eFw7sxefhod7PzpqScugoWe4upBXhl2eWLyCNVdcDH3
xl+Um7g8ZrrczNleBQOUcRXUqLWD7vL10enhIRmcv+JFPJ8JErRUtdJWEFmh3F6t
wt8hQ9w1XOFDE7/YF9x2yLcV7FttT1OJimCAOABb+87uZV0YgeSCWQ2WkMj11QYV
SWli1KFJDob19LWmMYbCgF1WdkSP2CK+wx06OhkMgRa5TdgDgfc9y5XjHG7KGo3A
IKd0Yr5P/2A8ereH9/LqEz8J3422TBROgCca4ZvbaFLmsQQx/BjZZcg9Xs0E515i
SPDaFK/JgEqQwt9MHJEt6HyoF07e3pgPj5/viFt/mqgYGpWNo5K9vMXT0FdgEE+S
UzXzt4AkBacZ3OPYgFLmJ/UHibnqGnlbn+ntw8LBhY3uwdSJmap9P+z8u5w4GgbS
AzghSW4ZMZT+M0A97V+UWg==
`protect END_PROTECTED
