`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fd6VsWt/D7NRync79biLMCFdnERJKJDZCkMMdOgy1fgPdJZj+9HVhUc2H5hTCK07
fVy5ZSjsZT0usqjxj3kQblV/+j4C7Vj8Mw24a91r+0vBXuKaVZgoQmywmdJQQ1Yh
yAeT1rr8xMA1xW4HprfVs5Fe3juQZOxxWohpIZvgFFwui7PKjIdIYEIOfYlby4bS
SJf2O9DB+08y9i3RttYRYZohwMEzdqrVM1nrJ5Ko+kE=
`protect END_PROTECTED
