`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
az0/XgbkluFT0G0xre8ILQ27tdk9Dm5lMKEV2Vg0yhddqixXBH+qxOku3TEtOK38
s9e/toZ9sdgk0MBpp33dVEEAg2EGjaEcLxr5D9o3faj/6ISn0av99OH88BE4zR25
Qzs3Ke9sMKhm5y5LnANC+KoHXeNTzGdzkFKX+UeWW+O82FoFu61RDJp3BzqBQAwz
ikJUl0fIyXdDn0JnGdnp8YhSlMapqUWriyLhfVipiKnowZCLl0IdlGjL3Mdnz7QQ
Lobh1WBvwthCoQ09cgWQt3TZTJzzbLEhZWI2lTFeUsBdFyoBqTj4SH46tRVWW3T3
R5TdKJJvx8iQWOcCQQsaWsdU3t05TZW8pTJ1xv7am5WMig+BnLjbI4ae9WBzBwWz
0hAzorynDG4OxS+oBGbWdzjxo12JuZyE6hfR0Q8tvJ6rRW+zbS5GZokkVRY7hc3e
Ygg2664FPGFSyQ3g+y/LKd3dD9Kxqvujef+MlYIsdkcMgMbEkoXph9bYdOnv2P/S
+5H28uZX91oMDWDOwrxis1Anz5jmMLz6WRn6pMG0fzELwCIVDdS+DJJGNdb+jaz7
69D0WgvosfhXThpS34pdVg==
`protect END_PROTECTED
