`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MVo3KBKF5mDdCaj/bvXHOfYjJ887vM7Nb48h8Lqxk6rZbjQR2gX68Mjb0ZzTNpmh
714W1Gf22ktSAedSSHhPJ5+wqjjFplrWk4JAbEVv+qM+372V4SL1Zlz66a5j7GLM
np6Cl7sdlZ53b2OD/vrzQNW+MseHs0xTrFCuIPyOV0B9A9AWhZ0qfWogoz6hF0R6
2Tt1xgpHI2UZ1GjIcei2kCN/tfphLiK6OrcoOdLIWCKNW2aUhCihPA1XXsQaG1uG
qp+RgYBEtHHSxh2rsBTBBAuzJuH5McK/Dim8FQZT5UsDfndP5vCYRPKmcUkHJGLR
ZPLASSBJCR5s9awZTOxeACOqsZpEKuELHn1cYhssaDPtum1h3e0HzC1UE+fKt6l9
`protect END_PROTECTED
