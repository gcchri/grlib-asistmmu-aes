`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
725wPBqgJZAfK7ESzq9QLrutDwxHjQtCuQRRojh7qOqoMVeGVCAVTg2hVoFgesml
W31q+QxFN61o98IAoDyByMgY12eh+UN8SKaUicvj9p3P3Kv94DDISCBtJmT+gWGC
9Xl9t/ItPX3AJY/b5eOO5mefhDn9nawivPSB7/yyVKC3k3Jg2n1gk/8PMwUdChg0
pkWIm0k9KuXQ+y7oklvsWP4IoTWdHKEim4vHtcFHT6HCgJsHFyvJT//HQ4Q4FT7B
2PddW5eK3tKc9CSCNtQBOXVJinEQD1IHqaP99VU8AwO7Wvpjx29hNQdyqHVfg++R
iJSEeLGUCDMvXLyfvGvUgnIFBX87KlbH+tNrz3tu34W01hAsD/4gDatx4BrM5Eqo
55bW9YhgClOCJ+y+Cw6el8LejE/gsNth2W5T+muuGgqIjmOA8rBM1NTQmPu+/qAR
N1d+rqfPWVzdAUi39yUeDnKVhSKmqe84k8NTNQgMZQ2s7JDpBegBq15MavAAd4Oc
GjCggGo8oxarov6cMVfnVrgLH9sVj1b6mk9nApY0yL/mYH/G73kV45pn1eNZZ1Wk
9ANoh0JGbn2IcfDFUf0Odl+PkzDjp1EEUbul26dSYKvr0wIhxsVwo7mJyEPqZ1ZX
6iE7n3Qpn1SAxsBkPh4LWXS4Axlo5tAxo6b9ITaB3eHIR32+j8X+QaLGNOtxP+yF
LpUX4tuIKAIagU6MWalkYwLmSX3PrGc2s3dpzdLQ2OFBH4wxYNbHLSy6bomx/h86
XIZKq/RpZoRFCp+dazyqYIYq68/ajg6g8jAwnoWhEkDsKCJNniDCFQKi+/kg8g+l
nuWDK5O7wnsJysFlznB6BgV2mWszbnYQ5Z0/y5+X9NLCEKLaK93oPNyFUdyfT1yx
ZrHHFACEOs+sNzXvy5D0ZD1I7pO6SdOb6Ne/gOac5PtYSM16exgrmM1W8604Cc3E
ID3zjfPnDONIIfgoei+ND7X0CYhFkCrIy8iq92zyDur7PjzxoYL43ULukz+UHrh7
wvp7hknrTyMy0THCU9zVxKaRZgNZw+FKEbdoyBw3FSPzoA6LYw9sV3SlGE66Nc0f
QsVUqcu7Shd2Bho36VjJSeH0zv5ZFV9b0xoFdXAxEpgnUftUF6rXw/sC+S4FbEHX
ePumBvQ58dhI9/o+Jaxjq2mXtNLdT/9mA2mYMMD8NP5IfKNiqI/pHWyLZKkhZcUW
skRFQkrTih3LUZ3wAHKVspWCeS33GCTWVc11CnHltNI798z8j9HcmtYAfhZSFjjp
O4t83mAaMK7adY7jGBh/3eLZIBFgXPuERHKUeX99wYrm/PqVGZQ9M8SZPW8CMiX2
d8p4Gn6kWYY93LyPvhgsUBJI79ZlBuV+zci9JysvOaqaXb6dHeBgjyiukfHZbXOv
2b38WbGHt5NyyBmj1AVjo9u9hjmPcRL7kskG46SMv8x8wQnEwYn8I8ng0oAtsJCO
NKU45PoZS29ajkwUJaR7wJtSTKlbhCqPXqaVZPv7T+P4q9yLGUYpPQ5M6HjzGqBV
LlK6VFmiXbRWLmYhzdrsga/iFsxEq4Y3BEym5MNVQ0sWKnDfaLYVno6s7qYJB9uj
VN/sheC4z7TJSctjaby9OSiLzL04Hsrno+djBVCFJe8O2wNnH73CioOfy2Y1JTGt
Keyn9mS9Kn2Ps4adFAiz9KBQliFLiQd0k2aHtcMa3ktahnYgEm7xytg+WqnDgNrl
3R8pUqlo1xDhDdTFueNcsBAJ1DeusnZYnu38PGc5TwJWseFkYtSimP8V/3IHdrp1
fWmbDs07Q6zQQrUAMp0FuAjOOX6EZzjuzRk2rXEE5SzNjXAY7GTQn5+Hmvkn8aRo
zlWZGCq8mhKv/Tnq0Po0+SOuU05ZmfcxUcEpRmGtmNoxlO6a6cn8ytThqxcUvgWP
n9T3DL+P9VAEi7RSa55ujYmGL2cgCtNn/1FmrgxYAZ7CjbTXolWaxTm5SKEUpRPy
7SEBbj01BvUHbhgQYxT1XvB/FkzOmh+FU10yMmD1BLXq9qIKEM7vqBAfBNEkrb73
OzfWf4u49Az4M66RHsJJv7puqfqisSgi0hH5TNS8kxY4q/JpoWnASBfQXDaf62Of
/6dwK2ke7VmaLGIoI58PirK0JORFGDvxan9GghRJSsd3jAOpuhaK5PcoSUCRyymq
xn5L01nyymPZvmuT5LBYAcAn+kXQHvZIWtZ2aZxlkzBzREz3LA3ehxCJ6Yix/bp2
ytBFXYPq48uGWaxw0DSrAfHrYWLUG7RhGI69XGUA9WozbnlDLVCCFn+jcXrZchf/
HURjEZo46180+ULnVTpBS6zJeNrDJGxP8DkypoLfNaNNMNUpTLYxwSnQxzZkL+o9
1wOO7+ZciF6XUHqMULgk4SlD0I8b7xlxZC96v5XuoQjFMZJ1/raUrCyeHPgQQDWP
3RZV3foQu78GW86dI0vxCEo9TID1mNnakgI7Ng7MmccXJloh+MZ7V2lgfzRqyqau
ImmIQnzjK6C8cGViKvhmCX/mRdjHAo/UGUaehh3FBvu0tv+OLHB0LYg0DizcZXp6
JJCpkWme+RGxEllFwioyu+Hc9JN3M9YW5GbTzI6tlND/P9eWt57vqtXenVdhLmZ0
Kzpef/IBUvy/CWThfHdjZE2iGhP0gKQIX2hnXqiUTEFnhzTnZ9CIdAm5KsnmRNFy
BVdWZW1t3dd/C6PejfI/fir8IOuJeflHyiCyBntOSUvdJHikg0uoqViBDYy6/VrU
i9CTeySaS8SJUESNZkf4z7mrmAEhIhnSe61AIGHfSU/eBV7tE1zDUH9dVd2Fhb0L
nFuglefgbVWeVRIhfYTsKVeAtNrakxhzkDksdPlXnFLbNvsFq0JPfm/hKH//ZZyD
Nz/APxM4iJba4XfRI0lY8KqyZuPaNCXHL5Y1Cryvo9xp9P4Ew2uIFmLY4M32GtIU
DjBcHOLaEOHHlTDItw3V00EDw0jwrhvPwrEtFlJkdH0=
`protect END_PROTECTED
