`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+g2/Z/sV4pK3kgjAEyjNGcZdmBvwn9bWUNZR2BIR9SBHzuC3A3aNf3JKn9Y3D3Qs
44OKXsDCWMYJZBgEvlYP1EcXG6DPR1j9TahHC0ZueLu96Op7sfAKiFqQwk8CElZ9
MS7v8Ee3P9HRlsvONzjjrUt7t2EdJmLGzRef6h/U2w3gNTGPC6tdGNAkgEExRRbL
AtfeoLSiXI0MIu8Npvjh40baRG00/7wTP1IZu10F0cIUprp8/C4uEWkwJeOs4rTt
ScQFwqqAmpVnKiHwcJQ8fZGxawm1ycg4IEanvMXmf95329T7J4dh7bgdrZrsvEop
MP9t0bP0k9plLbAPus+9CHR2O9US6UDcXDLduJ62zu9xyaNc8i/flULBoTwMeAXr
TyFfI/m6jCoHAH92JxIv7ERNm+J2Ydwf6S1RTJrbpDn6z3ovKiT81ljw8oCAOE75
MC0PD/s31nU6Nq+mAJk4lF5L7GBC8/uwlRqJ2HrX0NVr9J7dd+2xVGqmihGNnrFu
+lGy9kRnOpLhr6xdaOTzZPNXjpRHM4izRgVIqrtcjLiT/nFPnoK74LrANvBpMnzs
kTGTGLlzKKQcEs08DHTFVAgCi0Vvp9PDVFfAzOxR/2e104qr/o5PwRett8Ue3Eli
3jz+lFFbP8kDfQw3eLtX71a4eCdkYf22t7J6sCEW3sGTGAWY8PnZ1j8z1aX5SOO1
JKObnhrRkaENZXZ7dBl0MdIShkGVOlhx7oip2I74jgwBSM9Ls8THaWI1Po6J2qxn
7Wp5e3w7XlfAeb43diOuLQ/X5Mml3rHzASYsaEVgZbEAIh83Cqe/v9BJPyrEWAbF
6n1Foen28jzmVlNPIsXWJV1W7yMvfGEUiyc8UNSDBYq5DqTewsUVa5NF0zX0JRmN
Vqzo7koIZMz2T8RFADaJEAo7CUSu2NLoHBFynq+p3YrVVoywIpkgoJFTbECJpRPk
DoWVqIX6Cotth/wSkgFqFjOc1xySCrfUI7EXhu3SRSYPjG9k0FGoYEN4EQWtHXVR
biVSFqd4f6ACNSYPgNoQBes1L5YntmTBV1H1genvzRYUQr5xZIIOlQ331Gw79+4I
Ca2s/CVb9pues8v3oPfgccLlEPWSLjW1XO1NLa4acyOrU7i59FPuRJhV5CddMvcC
vfSiqFOxx9+XKGwyuKz4Tfmlu48jNP66/lujHcvc7unodVolm5qHslqxHjRT9fQV
kbPeiPSIgnfi3JH9P/eGJvOSo2nNeEIx+EUcjRw8zMkoKK6vKhbGt0qVQT7bOExG
1sQJRaM95opNoCzF2Y/K/1qE3BZHn8mDVyyT4J9umv7v/vcDHb/tKPhg9EL8mCNU
rZfToLQVeHUwRuebyMH+KfaQKzgaEbGeWDC25b2u4QX5mBlTNpgydAGRu4g8u8rc
E5fRYLUV2obegSfRGBDE+pMQVMLQLxRtnc9oBHDutuL8P5BVev4X6KIeJhT0YM/z
VEh6LzU0Z6HZHt+McbLdnbKKO9vmhZ4rhpCHtMyqVSDrOSp4Q8MNdlFJlosTE7E3
DSocyIt6nNXaTLf8xnCnIO/vGuotYA6X0LS052sR8YlGTw5s/YP/bvPDNr6qrqRa
7KoqKzgjnBa/vSshlAnht42Jq0wB1lTg3/KYmHSiyg2j3njoo34GbK0J9vDdpWm2
TL4RTWN2fGAs59mUdHXVeomsKtekqmwqtXnA35ZrGFerj51sIVHNkp825jiIwSR0
JGR2850XBD8je3DlE+IxnYNBYFT6NWIRDtD0TWaOG5JlNQkx5UbiOsQ9DoouYGMV
aKkR1NMBLhB/SG6xSGCEQQYDOynuc6MG+DJueizk43vp3mqhVuvDo6xEQE3+Rc3h
w2bSxU5NWqlobIPdgVB4PgZhKuXF3JAQFNX6ikm9roBQrCqx7ERPnN7jryrEx4y/
BAibcSMeke8IfyM89KoQ/KtXEiFT+1xRGZvadxcG8FA766j7a0cBSOWZl9Tfiyk0
qoIkNT/ZlatyNGXeZCbHizS9Yxe+wPR/zpfyVxp0cQa4buFpa5kJl4KUOFU1Gax5
X7xmYrbY0eb5vA2f1i1mny0sLS5F9pdF9M1Pe//vgmRzyZ7HOPadHw9skYIRF7JQ
O+Rx0VEaG5Eig3cDO0gNyoqKjOaHoRz8wZZHEjQoeJW8T51jXwhDUBWkyvGOKqdL
LzohLSTiXuqUNa5pJ1rzAkBOASdL5bpIA6ez/Xeku/U6rM5Kse1VxhTzgrVrtw5b
F8fcstlDUGte9lQ0lXEUqXbfihMCmZcZAgAQUgYYivLJbdK8YIE8ASyBooJxvr2+
kdEtHrKThbpFX7F4i88XHrqDFUWqIHeWKmpamOO8+CeiBDMiwMLkjCdeovtHJ+rH
MSZRsyfsN+LkssXsWbD3kxiIb+cYnlRlg3VqZOC/ip0mYk4r6X5P6tnhuNcgtc2l
3l0ok1L1GH/ISvQdr8XW7CEBMNC5dte/azdjgTC2Xe8J9CrhiBl0YowzfRzEdCX4
e/KRx+Eqd0h4o/YIBoH6J5ZDAYvk5UEjhRcbaLehXYJNeCEz35+pV2rYaXtBncV6
WZkNiZ4dhUJGjJmvkbd/1wdMLsk7u8IAr/+xgutcie/omT8YXVfmFThF9eqnIFOh
LlGVp946bg6L4fRLhN9xbiQGJfnJ2NeUAmFjOBT2rjGNxvrHhTmZuNTJmLoEYyqx
a5IgA5I5ucLnkJ1spxybtKE8YoQSk6jS1YACl2coC1D47aStJ+Dazk1KGufpiBrk
B/BuOEomxX6GdihQbWnSixTzHa160pL9yGBspfxX4mE/LjyFUZYsoMn1tFdMHlxn
GH6NmFQv/HgrRxy4kUb/RNqCKXkpS+uAH8d/el32VNVXcWFA3tW+hDbmKnAOWXRK
63iUkmN0ZW1UTfjBN4aHU3eLTVtOT3y4LocuPekwFcTA7VnRuCNDTlmLWKYfS7gx
cwXbMiN0g8iMnj5yW6UXWgckmb3TseVja7tysWXvOroBF5PGP13KOg0XPi0lCMZj
d8lj44H0TDgK2lnMlG53O1LKSLc1YXac0IYPZuvnZn2kVWabKxzjhEsLB9DQc8XD
odPOLxmAo35fGwr1MmzS+tz9OItXi5TO/dw+w132GDo3adlJav2H8hfEC3E2xlhj
b8flPDSldY8H3+wFBKfUDkT8+WUFQJodu5Cg6AL8YrwBNZGtZZZaIRHkpHvC6mHW
qbAL6weZqcpiTSke3vThQdDklViadR5XAvjC9776G57l5XP/wF5GbVgXNJEHLui+
fmJm+MmnjWsQ29gdm8VOOn6QjNpVH4vqdrpYy7QKZQgtv6RAMY3m40q/arCxAlFu
KgcwcxKZQCM6pq89R7XLx2z6PavSwde3M9TwcAlyKTIVbw+zzEPyMEIoAA8H/tme
DKUwUgUXbCPyGeQFrGpRNgXO8kL7MKLsyQ+ViUqJSgEq+iN2sPbW12TjWuVj1vDd
SHtIU0bF2s/D14yGO05/icwWHWZ8PiSNthBa3lQyq7WVVQBluYJnRJKamqJXPH6s
1CTfkV2GeGJH7EIVq6mSGVB4CBkTrx+EsgSHQL/0WkzD0aRdyioI+KT70ydAd1jf
7c15oL8RlAM1CUwVzPgBMcadZ/gH5BTNEr/1dDZK5SHepJxinJt8FrR63OIC6gl1
gjjsZoRP8jlLbffcvla/7JYzXe1/mfcIvUkfB/rI7dABl61+GSVacBdR+miVudxo
FfxflO6e2yrNMwY79CWP4+Jv3kr2xZkMkhJNq+o/W02Bduk3whlsBcIiXHUbv5U6
ZHs1L0bJkMnKu8LuWfTiW1IO8DM6aIzR/s3k/vJyDNCOjgqtvTsQnTlkDAyCkrgu
9GjjU+FAR1SbsmsvQNJdPtv+EOMX7j7YcvIRdyI1lmHSRqpS2mBaCCQHfX2NYFOe
TgOaBWn3HvYFFFnrS+0qMqOFtdy9jO6KkILL8OlEtmJmcgf7bgdX5ntvg6z1EI9A
akLkvYoxMHQOg0W+qOjpmBztkdwE5H5P8O3aZfGy3E0Azl67OJPQLCvlGMYSh+jM
l9oCFfh3mkXGL3s0rgXv03W6Az8uLdp1VzbybWOkW3TG1KPLDihVj8nTyynutVr7
uEJUhANXYztMjwFis2dCT20/jLwMxNqQwcl/EyGUJl5KkJdpcppsY71Qz8LRs89E
Lvw2bjKbh4SiJfSEkfP0rcoZIjAaq8/tnm0Ow8Fp4KI4EU3iDPRikaq/UHx8AFkc
PiJJekr/bjrl9jPyiXueenyUEjc+qNv5DjH9BGm7/QWUfe59XTBpLPKZwDWpqCcq
kLTXhR3hRtQSzKIT5dm5Zuda9QiUrsqhj5PXxcMTtcA4dEuGTn6Uirj3Dk3AHRUu
hHRdOGvpHW5ZwLkbGK6rNv94mDZf1kKQX9uFNxDGBbn2NQGAO29hAiR+IYUAUi02
kpryxPgbiBklu4NBCU3ougO4Bqt1gNXmBsMv5z0ZHs2XDREbjfUSd5In6byC0E36
GN5arHDy6yUUHiGQEVn6qdcDBqLqg8UqiXQU05mIWNbKwDRKBm37aDidIC+opPzs
XjnMYY+1MOMjjWCOlWUfa/lkRp3TMwlBDrNONftrcmw/JyHbCOwzEBH4CF4w/afq
p5e6XTqaQlyR5zg4G9+6m2IGR7KIoFx7iyQu7eXxVLobGxFlkk7ti5Cu3N5d2RMU
0zLoP57hSVavpCp2Z3MmanaarMCL4KMGzEed/EUNclouV22oj6zquCCPTYhi1/pD
S7Tnmr2L5cT4BJu22vwnrlWkCpc3B39wm8vjM/rOcZM6QRooCkHAOORcxfl+bXqq
zVOO2mbMg6JGIAbDc933Fx8nukeYXTmTggTqtWIiB+r9yVnQ2KSRpWs1dCT9/HMV
W02UX2XT/cgrEOooOnoN6pY0wy3N3DHZgxayx+yvmhcAWGPVq16BKfwKC2HkjMZT
KLDTl5dPCoG176Y2kZ1zkYlc5dcgE/52617vA6B56gVdsKh6qVKwOCtEhk4xgfh7
ITQ9Dh+jwcLj6K0+QZ+m3E6QT5XDOOtS44vtgcDet6KJWjvjpkg/wo8BDr7RBCOS
O24Ktrshq/0B20ADZ1vEFveAHMTU6wiMjcSqxUdClTof9qRHhHv77oycF/sW4o9W
WX3SDIlrNGyPGfjJEiB53kpgcrr5O3DzMpypWeUYbjn1fC+C2k+JvhqpdA16PGkX
1LfH49PVFw9zbX4PBQUhAXXorT/qJ+hmIQ6O6CadTtbosjH0V7XhXoEsNFghTnOH
+dRujDw90In5sPBsffvTjC2kJJXZtqZ8AdDdCSZrcdGpfio2o1/yAGwY2nPAlx9X
N8U0amQdaswARJfFvO88JKoQIoJJ9U6W5hUrwL/+23sWp1rtiVP0WB1FTmTDSPvV
/iOvnpr97oHyIGwgV0S9JDwCVRBsuj+q6J15MuNgtmcgrReqVq7CdzoXHsr283E7
Fg1MaqRziZsTzuL68f2aIR7sUM7hg22YcUbMbgD4s8E2sZQ5cjmahY5UHEAn8Pg7
CVWu3SyeWsT6siJyM1aw9yTZNPF9BC/M+Bfg7+URvvX2ZRcy2uh+HOSQHobiExIs
IF+Xj1uwQ54mXwlphAi3yYQI3KSprGMonmwuGZKd74zbHbr0oSrC+Q/t4hQK5LM/
AJTkOqxESoGlxzieeZZyaT8xVX4qmtw69YiaaiEhQP4ihBZ373H09C0zWpK4cfXk
24ON5MPOVu5gP+0yhtzZLhoVrWqhPKtL36YMF/uX2+q7EgzwDKCKnEJtP2cLtHgR
6CqROOwDbVTzmdW1V9VQUjtG4R5Z1eV1JA0YaDLvaZ3NJ5jyo+wzIiEySUMYO0X4
I2y3DYt5HqGolGoBolTlXQwqm1pCexpUL6u5N13nNw9hkUXXIzMbs+2o0ED90y7f
RFAg6xTAe326ZlApT9WbhFAHYAKrgujUXGNzOAoZEM16K8L+QC5yh/c9pgRaCjUu
UeclAryrWQgdJXPX6bePfy7eulj1y0rk3553BGaGQqnXdvhbXW1WKB3rYd8Q8c6g
cRkC+7Vg8+Ct9tn2YqR+abF+bcG8ZWwWrLCbjB2V61Xv0jiuN8F+bXQJn0MtzjGn
IVCXr88YY8gqTCHi4nPTYuhweexsgqbWc9Nb40U2GGx9VNIpRY2aDvzFY2+t/1BR
pDdtwYTpxGYPwV7i8Ym89ba/M/IVIA0U1TvzwHnfyDkp3ISHE5HQOMSaTCMPRpJd
yMk1iIvm7s9wR4dtLX6cB2ecBatmylWcg2wdSns1X9oldD0g2yDFRt3oQzOKUkly
JNmTqKHNIpdEXjvv/s87Inwhq7NVmUWwWIMB3rnSHQz3ihR3J82Y50tthRZP00pS
k5F6Iq2kgTOkeY4y44bfb5L+fffzDt2PezgNjDMo7PY5OksVHvAyunZ7W4EQTaoE
KWd7ZNy9yADcY8m7zenKQZT0CVa6MYA0FZXBui+PbULqG+yZThov32weciMVbUe8
2JhW/dr1b6lag4OHcXrYJFPdC67WfRLGA02p560QnH7MsLg9JV8SiUjcfTOuOQQX
K3ABaBiilaGHkfoxdbdKINHEF1thGCGg6p0LEgxOm7K3hDBKmF7Y8Pmc2twTmv3I
fgUXqw5YQlXY94jhgWPFOPDq38K2cwpO5ujjAlon7bmZsV9K9vHMO91WIaR/+sc/
zQsUfbeDyDnAwUM5fEz06+70lPFpQ8wgjPU29lk68oAzZniPRtEBmnfcp+QzSTa0
at5BR07ZOlUVIYHFVHAdRG5RLpK4sG+22A1Sl18bQQzkNFY364CVvg4alMd3OrTI
SKGSeFn7uAtjOvNlylKpBW2kF1vtNLcl5pcgC7AUhsMGBKYb+Zuw9Eft+wtz+XCQ
xQTgpnvAUgVMYurc8J5bujUewtrU791VmWDk6LwuAr9CHBvazDpo0HHp39NuOjdq
H7DuZFqAsOy8WU3Vfw52osREQElvVZUfH/uW7WqZyILCAZIy4vkZXQNAGNSBHTrq
8O+NZHV62+WiO200Q91peTfSzws2tBDxtTaU6rA7togmpqnGqLkSsBkOMVKBzpqs
y0ET7kiOUMRjoam/Nxi3Iy8GvsuyJwGXvswAogfGv+v+67FXTzWg/TX26p/VhlzV
UKXWxOuFgcZ79+ZHEEgxtOyPODBqNq3N/kt+nssnUSNljN2f2pBPpyQUEHEiHAAc
bM5tt0y96+3z1bdh5pI7poPUOvNBYR7FrzRu8ZhvvEd8sArVwM6AIsKLeNCAQFv2
zeq9vEV/cMZDORyMXKR4UjmAe5n4mfoqaCoymOAmWavwSlteOjl3iLOND1PflNde
DEPaDJMoqRoICktUd9QZTG5rwsQadNmi9cfj11lKnUEezGNXf0xEuHgbzobsT/4I
SjiAeuqBowQxVF0j3MXvL6hqLdrRQgtWTHBhIfsr/H08rSijAMnEOVpUHXo8qvm3
dXzfkCgfzupMItv87IOCjDd0NSDLGnpzEsr/5WZ5WhGBInq8IPk50N0ATOkB4is3
Rl76h/4sLTf6JlCPVtrb/ZsF3SLkZM2DiIaHqqRD5+lUZvsNk+wX2sRE6rz2daiM
WFh6WrLMOkk7WzfeGO1GZbkvEqt+CfhztJGWjVKjXl3qB2Hcj6d364U5ECcLRu58
YhVS0Ht3uVxj63Yl9b/bCZXac3Sl7Udc+Ws4ZrslECCXK5p0W85087dDXqCcRohc
FrPz6kG1RmEvQ0Cq0KnSZCRPbixj11r9pEEfe/GUJLL6EcrsriAc1f2IkrWVjYML
N/VnU2BxA7WIloNCi6YZVAcJ4CO9njoF99mkNgiesCLjdNGWdWhSnbqatmWvIzIm
AvX5BBMmLA4dPVQuDo08N0y6+44t4bwcVJaoZ5U9KSh6WXsy1PMZ/nREP/Lsg+Vn
KhwL3pZN3mUrpXRVvPg5/psOVdWZUFhCaO9k4p7J+ajOXmf2Ujia7eexCwmERl/C
byU9/J9/AFgPSveujxwdifn4X7s5D61fM9ikS2wWSEdSbBF/CGBXVaWG7dzwzGuO
2uTtSU1J+lLsUl2ikWHX0J1Cs5j7475axflOtQW0G6o8x7Tr2SbLkrJYquPbpOcX
E42D4WwndNwjB++xMqkvIJbZrv3GgvyntMgjLQdRGzdEkghi6QWEklss69tsgEmu
ZYzcU8ZgV5llzDPAUnK4wc1CClKac/+M1noV/ZYC4VxgXqzjI0q3+mzGBuTzQnul
YHSbSBYkP+TNy3/JDS24Ts28nPEsagdfk+huDs0gf/Z9yweVNSLVFrp2RIIwFMZS
bRx9q57SvNEN4c/95PHgdOu8HYZQ2ZQ7wo7e52WCyMYnewZnpmV3kjUJaNxocHOI
KZsYWoVTsQ0/L6qkQ1m1typCgplLJg1fQgRaw6ijt40oNJZ8GVn+FSRaUVJLqvL2
PHhqdalleHj49oMox3NrVm7PDLKKAVlX6gtgLQ7CLL6sUV+2BbytIFiDPcxm6OXr
mt2/3PA9C0KnHj5AA0cl4Ao/NAbTNIMk9abKEEC7imP/jiF3A9hRVMJl5iE0WAKk
eQtNRtoq+GwQRWMb01/2cHlDc7Iooy5vSx0VNYiRLKju+h+uAr07CxDN1fwxSSsw
NNPdbFCZby9pCFG1k/qdJR0j0xh1XjsmnwdMt4dFe1UbYde3/OZvGw+RC4sKUYaX
1juns7Z9+dKtOvmc7zQQdBM4smqFvC/EiQZBc9UEEej5Eehw/yxTWwzFXhUuDnAa
GF5/MCULlukrMeEpEb0ex79NjcSF75E50J2+C28QCBozdRCUm5EEeKdWMETikFhB
V409t/fcEDXvZ4GsdH09aRwwgf8H7diB281lm/RBZeNwgQhBv6VcWFcMBA7eVxKs
4PfAEVTr1bCdOSklG60MW0shUC6mzLMtpIEeg8V/KqOPQlR2pek9qcy37Xwaf26V
hvAgSo7rfOTOGt6oXF5rYyx4s0eUmozcxBYaVHIHgAMjUbcjQBmDfYsJD8Hgn7SR
BF3w8IgdN6yQm4IMmXEizbzQm2QVMw6S6vVehkKuzVXXy13ESOxWkZrD565bB9PQ
CeCykMiENwaWEMKN7poS6VLAXrt/O8LCu5jfRZ8vhUIm2U3pKOXS1TMtevm/oy7o
MVBI0V+MNOwaogOrjyj8o4AaUij59EwEn4wdcL4QE1eR607ye0v3Hx6NJqTyQYUH
DXm8Vv4PSI5l/HP2sGdRUqJkWpN5m0G8Q+q7l36ZWLkbD/ChUKe9U8AlRCBqnhbY
GdtPEWPEMTBFTneCjLApqDnaBKn+il4Y2exYgy2eMyA3IKC1YJKxezD/B7+Q+YIa
k8dAChP0yDFKTUpynuuMpwR5lSQjkp+8o9iR711ipwY=
`protect END_PROTECTED
