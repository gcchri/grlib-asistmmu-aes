`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IVHT/LQkqO4/Hy2Y3YSv8UpYZ4xrIYtF66Znh3y2ycd36AGWRtU5aOOdqPn4xQte
BfAy2jfm2Fers+eguFRfFObQGdOtB3jbNmSq8KqKOknrcGagrTJXPbzwvDsjqWPZ
iPzb3Xog7574wtBXPe8m1j6xUa0Tvb1jGNVGAnMRqip31qFLxkQI3njAKbdmGSfX
IxuB7Vk2uqhm+0tw3P427rm2UwQ+xZExN9O42G4w58QqlMFKL9OxAebJ1ExdogTc
xs/dwRYA4LPATIV51W0+lkfYfTfzj7ffEEPBSqxCdUq3b4PQ++/GYphfcD/9QYAb
ejZ3IdmogydydeNlf8tfzd9o4eW814BaWplvQNibT6pY/hOnk11p/+OIwJKOq8aN
97NupA9R4MryepsJEhYapQ==
`protect END_PROTECTED
