`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jUib+qKF97pT2We9Zy4K9Wj1+4zTpol+KPO1MDGq85os7SzRODROABRET/g4Sb98
faO67hWZa0/veeFReAU4T3ih226wHq7giYmjUPMCe6w/ag+SeOJbRvBjI9Bn/ZUn
HxfQVxsAkC/9JQZMqPpDiVJyoWLWnvkyUs2+zXzJoCj0ytLxD/90bIsM4uq2469S
HRVSRdxxNBUi4fAR7fgqcH9RfeiLtMe4siSnfIXKI/ye/938Pjldd/QrzS6FGo+w
+je5Jp1iuvoXpXmxZ1T8prVUExbBLJOM75YNsMIvCWGRbFnd6gs4CP84ONGW214V
sfkrZky0i2kabrI3YbEqlRI05oenka0iFUk3CQEyqNvnMWNTP9eTndxq/kXkSLB1
ACimg8aQYzL6ydxgOu4bIkrseUYh71K4CFOeeNFEznSk7++N6+klJMVWc8hU9CIY
5r299VCkuZQmqrDhXJdziw==
`protect END_PROTECTED
