`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O5d4FxPjUfa/tpP3Ahbd9hTwFEdNkmeEydp2rtb2Sof2w8gdW31E3TnxcC8XafAg
xivUIlFCbk+0YlZlfdl3Am6zwDjKNhzLBmngnBU0JYQgu0tXL+P9aJEpHTTvuaFR
M+yT/Nt+h+o6WPGB2u4nPHzXxqrmvHDQ15s3Mszxw0OD2GdqzBqBPyKZLZDA5RfY
4ArbKhl+XcPhaF4ElrVlkbUcjSJmWY6wb2wMBv3tbtRnQ1G8Wb4esRR3ej/GN5/B
YIVyQQAFJ3YnR5xGsx4vDyhDE5o+w+lHUch5QhxWdOE8fBdOb3lbTzNl7FVXxC7o
LKzbw/L0ytacZF2Nd9KNyQ==
`protect END_PROTECTED
