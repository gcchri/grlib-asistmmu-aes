`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
35F02ddBpeTbh2Cofx/KFUfNyNC1H2z9RcsXGrOYUCNLMDbiqvDIFMrKo0JD0wAW
nVyXDyk+FzC4Dc0mhuDGQbhOBbf96RHouAxqZag0YJP1BvD2bKFH3nusXsn3pDHJ
kOBRsp92xFEwbTtyLuxglSAsDW2wHI9WKQKdj1z20Q0JVchbxOKO3n4f+1GFzqRL
JOKC+ITUA4NMRQQWRV2MbqyPd/tpwlm0f4jLMS6isJ51kRmx/Xfrqg/jH5sptH3U
kNlj4lpHKiBo6BdtLtMEryh8BtfQkNITm1o1+x1uFUqhFHtun2LGdOQDZl4t0hq1
u/3OusSIvZ5TxPimM58oSVyZvDMhcF1PRTjOpak8r3x7gh5QYhtVIe5/HNOBIuUs
fw0q076WFnbXe9DVA6fFvJDVqi6fXJf9NoMqHEY6ebpbU3lrdqBxPCLD30PgVR3L
z1M/QjfIzMknZqnxIwf306fgHbiC/Ne2xau8TaOg/ByzsVrpP4g/HF0WKUTnt8U/
sSaqd4Plptm2XbC4ZzCPIEMOiTr3jr72oPJIkHecIBfTE/W3tsXrh15kPfhHhB9N
a926NXnX82dcBxxFULEXUXMmlBeRyjTRRW9sdv7ssFA83gg+8VDtwPZ+5XYTrmi2
9ANTiKXFYvlx9ldpDVMJSLsEzjjG5qA0S8C+QHISXPdZ6AIhokwLpKlYyIBnUZPt
K7Op0jRzNgDxA71yzLPAquOpUVZPaKxX0XhgdhIMjyDPvyXGxAAZBXLyursPaSaX
2kI+/aNGwHoq1CLg7YzzY8cvEaYmSAfqnJkPMuJHNWrj3vxMgptkViKAbTgI8h/S
oFMZgzz4PQRwxVWVnlhzZpskoOZaiWogUCObQ+g+qPGg4gW4MuwN+p6oxfgWdEBx
7xCP6QLZsoyK/ml/xRnADlTuhz+pfaCzwmEbaNDoss8O09b5npAC/CkLkHiY/K3o
ESEMX4y5lDSpnD22NwpfoA==
`protect END_PROTECTED
