`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3wRXsFORptOfdHuwYhoUFCZwiWzJoeCaRu9RYk0W+WNGIBbw7Rn0tNWOPWB+gOwp
I0wJ3CNsFrYa/JbONspmhqYR8/snbfTy7vibX18V7de0cs2lHLrFe05ZTRFDVFj0
U8WdfhZmic5PthdOUa4770baxZmjB/wFtmdzRgrHGArylEP3uv6Bd3qTN3EoQ0n9
8Ltc4ai5CKVxFvQcEs8pUelo+Oy360/3r1M4NO6apRVn0/01aeBr664vBxKypfzf
8Mb0UnYfOT2SKxSYQUoX3UaH52JeMsVDKhPgjc9IZWyvIMw9SrLVp9aWDfNDw+bi
7AS5CNU+kw3KOLGv+BEO/p8/zm/KiYcpE1t5lAAHueHdmIzzKvlCTgtFa0ldDH5N
ZdBBUUsw6abo36Q3euBG14jv49hNDHM1oPt/BLchZHupMlQyxNrmVRQQJz+HZZHu
g8PtqAXV73AfMDZPvYbbwqnYhWzP/2Xwf6s2Ujw75XlQxRZcr4YyVnYbsFlrsI/o
Comwuuv3dW/DNNVLsXcn4ldjKVVJIHQo7t+SSTSS/mVsS8/i6JTkLBShI7ItMfo6
`protect END_PROTECTED
