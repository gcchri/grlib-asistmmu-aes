`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S3CpV40BXbtDDX36Tlp8aNsRyDMOaJYmfzPvS2cZ1pw4AV70WF17WjxRRi8KTEaC
kYTz4AlaV7kSpr1XAldL1puwQvI79pVCNxtCFTWeueku+3W86BxotyIHcn2BfZS0
N+k7GpkQv0pALFHNAup1fBRpvRMNlFyicU5iTVgtTwiQFU7kNwtApVMzGlOIa17S
Oq1rT8ICQYk9q0z9H2wHAoHAzT2MvVgNYONUUVbEYHTy/tK94P8GrsiwCkfRtvSG
hKcaKb99X5O4iQ3D9b9bHd0ww8dzUQAUz/vfK7L1MmFsvihSHAT8sTc88QbaCE0b
DITUbY1ayLvfXcJaIP7xwyXOFqA0pR2eTXPQNUC85Dd3cmM86u9eIzfrnyIzv2nd
oMOJBPWnFsmPkadOHoiO4TcvZrBGYTXfKUAXkEqVkVc=
`protect END_PROTECTED
