`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UKrvu3ek7q/qWK07bGBu+c9+qEZltLx+OByOr+vUsPV/usGvVXySeTdXkErpY77Y
05FyzmwZDU550CA/s5c9f0tWXFIS7T9xke5iGT+opRU8EwodmHdjpeKqN6lXaWv/
HRsPZNj/f6Y+XJWWW5v38Idzha8/LnRuQecPAfTcRQjgc+ZlA2RfPlsmBc8NYvTx
G6bDp+ZpsO1okJ12F60An+5ezafboLqsdpXlTtm01zWBhT3DCYOxSpyupx7fBWvc
JIxxNt08EnFg5kfu0u3yLTifiTip/6g8+Kwk5ZywDryLNKVPFQaG7xFOMLu+G7KZ
5wzqtg66ggP6Q+J9TTwVbn45WWM6xDTXEdHA3mtmU0f3S3+4L5MFB6VcS5Fi6Iit
t6+TuhovzmsZ+Bjk0FhQrjh88PXxJsb+BOqC6jMAOrxO36mNDdOxw7VUICzs68jV
ZLYPaBPByNeGaQ4TiM/egjB0Jzvvj+6fB1ACbuHVcmE=
`protect END_PROTECTED
