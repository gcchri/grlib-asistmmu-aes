`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o0h9OW6dVw5r99XgoanlMurENYMZGKLY/GZO+ELLRLRaoEQ/UdhmRv/4i3RZ6R/W
Y1eprcMHAfHyf5jS7NQA2s38Kd+WNJnp0HkbZrtcRLFuflkSpwoZDN7Tzj4AHBXg
3AFu59oG2e/FA0wRdXRR1C2w9fV/xeU5qTaxVFzbfJmeBhhY1JXZIgFY4gbbULlR
AW8aBPvDdLKIVlFO2oizD84m8s7vkmTUkDPZIW7xCfK/WYFkxDwVaKPcwImOUk6a
3wKHbjqwzFM6Ae/Lv6RxGDwlCMebg65zUgMYnrnD7HfmerBjbsGSn0q4aPQmdqvm
hF6tHs/elG2AMBRiAIJValYUeZ99zhHDWyUpq53EJFu6nlRBjoq+FhkrtumIydLQ
TmjqrakYZCG3M5Ccu8HIRDYgAnFf0tnuZbWI58uEyEFxUObdb20gOm/II0ejDrqi
7yPw9oBsG75TWU8F+34kE/JR9hsZ6Y+70tyt9hoVk3q6iYppJLY9uMzwghSiCNXM
K15oWEpP1lSE5NpC6JJVfLV2XPLKeaaA6WHrtx6fu+zovbCFHWPfsx9+C+tkETKf
Advgr588JF+FdINAXam3r4v7bGgXKvNENKvpOiSnyCrCNFCKYVcn71mq6WPj6i+n
kAC/yZU8Pa8ndR4AFvh8ar4FgTKD+TyNNCs7PESCliu8ttOm2sNw9ia1MJI0HgUU
hsdT/AvTgOepO8WHIzUw6/oe3+bAddlHaIwTAVRUs5DbZV28mI9zUSQXSJMUa0M4
Ru/1MF0OSl+LuTCOUyArDqQTKOHRmaNuWH10Lwnz2NywOyhMWZiell7cfrFSxe1k
i/Mf2+LftFeoX+wo3++npkCNMKXDVw/SM+0nNVZ6UVFIVeNn7vQN53YMQRXLExjN
6fP3kOnezfDnm9EqgfvbMXjmKcIceP4fiaJ1FW6KThxu1xWfeEtsMcmed08+mHeF
+S+9lhafRRUXPFefDK6/n8vS7uuQJ8mK5qkOxO72jfw0LxifSfSGDqV8/v3ZKgyU
BPKiu22vjlQc2Ti4SYKrOfI3gOOCNc8kzx1NXK2CThx1AVlIFqhxUSzCxxz1Li6H
PZlcWWPTaB3pMtO5R1W/LyIr+QNCPQui19oRh3J+u7+qFdAJvUC7rsFzU4aEq0zd
5Sw1BLAZB8FjdeGg6eJFaYs4upjgwb/VaXlnqU0PRHvSXAjYDo55w2Q1+qUSyyOv
L3HZBtV/aRnFCb+ViHfFTlj/TXXiem29J+frgQekrwgEBslfNyFy5yNarD2WvNze
yvL1/qFZ2Vr19k3/f+ucmFUuR7w0zyBFrlbnuBZ8IisyutrcDaewk0KoLZyMoYEc
tWaHpEU64u+N3zah1IeMv1xRrUD3NlVNoeCyBpjUM4zjvYqMUSRxrwtiyl/W1jEV
fl7RD6+z4U6q3QWwwZaeK9jE03z+HtPndJrUMN9VX40W9XXOQuWIE5u0md99eBjU
V+j6NLhbIQde7oCTdwgZi3umApv9eJcT4dW7TDkruoSNz2J0u3e7E/Ojke3mgF1l
ufDCqyt6lT5HFKcB4CZUxuzhUoYHo5MIrBX4h8DY+sVPzDrpzTsZikRtK93fWA7H
BorCsh67cakL+VFluxV41OToYrBi/XVf2KxG+kiFhwnNHIlQXJG6vLkQD+AZBt/D
0ljUIuBkvvyaCCJyXBylfK/rPdkqiuhVBqb7RLPmXtJbVCp2sJ9feR0DT56x4Jlu
P3VBQhxtOkY0X1XPYHtlkQ==
`protect END_PROTECTED
