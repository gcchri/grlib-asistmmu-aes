`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EtMTR9R6DCRHY2Qe4GCV9cIJJQKiTtXxpBiKj0PT0wwvjCKHqNFbgcNpXAZNsOZe
EXA6PKn+IgD+IK4owsIqzkM31j5xx3nR9zDX+nS3uFbjJYtUkAgFSNJeI8O/vgLT
9IWDXKsqaV2O+j+kzLYz1g4+E8/TIg3Ayy/lD2uI6ZBk1q3QwbZnJLt2LwiOyxaP
Um0+oIKFKMMAIzLQL0whfTUwzDq5swFUu4bJQHAcSVhxiRsCierG1MW0P9SF7JUI
/MlrlLPlNoKNJzuXn+kjqOHYTqS9LcW1s1uY681F3LH/jWp+5ynjTgOTph/fl/lC
9KjijonHd8n0rBhOCNZgDQ5fODNDu1E3QtUtlv+BI/36qhmsCU4m7pv+nLHhv0Lr
cftNZ1y/txj8DhP9sBYGK4SfDHn4i8vyQx/7bwm859qiGoZGToTUTyijmC5uXtb9
chYTweJKL+TLGY6ZLkjkiI1n31CimW/Q4gmlQxTovgw=
`protect END_PROTECTED
