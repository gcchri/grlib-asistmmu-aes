`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1rNmhrDV3ppOS83KNrPogPqpIDTTlJJSqgLct7ffPp4KP1oZHPJeQt7RZkknrAoO
V6EMrSxphogI3+nYCX65sLIy4Mktkfh6Kf4WmuvLyPSC+qu03kNKHZjnzbyPPC+H
jET0I8UTP3LtB2PcizLstZ3pimtJiKYfOoF/y9Y6t32LZK2XjNr0zLOjHH9BI8Q8
7YWLm8hK7FxD2obxhQkvyOjDeDY8AveRGGMpdJF0ml7NlHO2XoPQ2Q/zoljV0zYl
6NjRsvJzECcPEFomaPO1UwblBP9VevZEoUutdW8+BmhMcMpdKu97k33MoPa5EEQj
MPUx3g7pY0Nhnxq6NpK2IWuchYnFfSrEKxy+C9gQsVQE7IepPzf6Df0WHfMP8Evm
b7H5myyEH1bTrqbKoOdEwRQRIbsLKQO/AQ25TvYfLONzSvX+zixZBTGv4ltQstbf
J501f3b4Z6S9jnfQymPzA6QRu6LyACc4+8ECeQkLDlZgqVW98Lgccfnpe06cdvtw
X7HI8AGWNHYLlv+xzI5ZhZiGq5s4sxaAfGaSYxOb2s8lu11d89JJHftfJuPwHKOA
XdT5NiPj2x9vZDE8LQgR6eTLY7tei2TZSChHjv33p+DzvizF1iGpOCjXQw5xz871
k1dSUMMybj43wLy4SzBriv3f8oZPIm2J/uIpiUCHZCA=
`protect END_PROTECTED
