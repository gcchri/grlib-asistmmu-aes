`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o1qVJRF93JVCCcSyv1zaJMOcroH12l2d8PCCm+Gk1sMAIxRnlWOK0YeO9mr2Mhnu
zCHaEHNIsAyStkWuxGaqJ1C9ZfykWQ0GE/y3Do6EZvuD5T8+I6BLysYm4iXlRsJK
hgzQ88hCZmvVqEg2O1DZNwFnrLgGmCUYvOcW3vKDqTlOM8WNc4oTS60AyHRdrgZQ
7oVCWcjZQQy9Y4CoClNfBuTiuufK0+pG0Ypc+nqJ1nMJswjaeHHrXfqxD5VdjzPN
OJmoYg9oRchPPjwH86ZqhxuBYoa6obUQkfdiXatNiYq2ljRFrYNPGxC3QllcQbiQ
sAD0G+60WviCRk/KlqVpWU9GmVDR1Pzwz3ULtAMnoyk=
`protect END_PROTECTED
