`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2g+94NRAqMxRBkCh6SK7HEb/0G/v83tSj30rR9IN/iYDKIxBxCF+wPc+mSbdXju0
Cmb16vKHrd6FuMFfgttQUkpUKKTFNNdnzCX9enh6A43lO4/uUPIbBcxS4sPtxNn8
0ZcAeEIwlmM6HRfjRfr8hZhOmne0XMVSxnc1cX1UBmkHKNlXv2VqYMoyfnn1yDNw
lUmATKLzXmQ2aiO0PdDFzrijXoxHMrbWWCxVi09ypOArSoCRX+ee1BhYTeckjab9
NEtkHvW9Yo9iQijZ1lGXq1FugE+1dMEFQxdqOvrBDpR0t9KDxdl7ILzJNt4MPksI
WWi08HgVmIf4lQA0TmMwmnCnrVwn0zuwOfPAWEC5YuUQbeI7cOQqQRc/YwDyE648
g6y47nkSMiusLBFOwNIYDZvxl/Ev6o4nVEAg+dkvbzMgY8dc1EdN8SYGhBFgscvh
i8g11F+7/EFU5uwa60ZgltLfBHvDrQi+8PmulB3dvQI=
`protect END_PROTECTED
