`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U2s/9OYu00ekCVi14yljIWgTwEVKnVzXZQTNGMDqsdH8ErnaKVhkSr6/8DEktCnB
tN1SIlF53SGXO22E4q10wyqTGqTW+56z2dC0loQ/cpkI9iH0Eym8wEuPIn/9HYN7
wxvfkjvh8OxYdi0hhU2dig4KlncBODwSipcCfciFM4fmT3FM2F23T4quO61OW8vi
H93rn/AWIToHNRDO/CSCxGFEo2ejA56JzUMfHMV1IFFYIwTKW0oWLdud+E9Gy4IJ
AIqxTUB21jdFAkxNZtY2b480+fldQ+PsGYpH5lCsHnw=
`protect END_PROTECTED
