`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rVcUrKv/4ftvy9yizYg0iTEYTr01QHp25CnsuUQ9tsF33tsLNGS8qlAI+0opZcB4
m6jGY8ItJl/4IsMXanM4G510OMuw1pbzPLNODOSBgEnc8+yJBzqUTebE2HzZt0ni
olVlYaEz/2Dp1wDt2PeT0Zj6XgB7goDU+DT5ZCqqaXv03axWXdrR84TH+fUhi6YA
t5NtnAjAecEG+RJ2IuQgYVmT1LK/lcqLpwPAPx8vLTNJwo6mXy4W7w8HljW73YUv
AQe8OM3nQbDZydndX6w7RVUD+E1S5R4ynEj18HFsqdhKQPMWMd7rNMYZHU7fGLUn
kdFzOYl6915/0dCOq68kdmxvGKXXxaOXyvN5lvCGDYJuNOHqiG+seDYag2fmyjzz
QXaZmwE+y/JZFYuVRekPGHhRyfy0lheUrQFBJUQYeulwQNraJD1GRRVzj0miaKq9
g3JXL4De6r2qcbhOkBIU38Rmiz8E8Qmb3tU/LKByh4geuvgpwAznHdOvYFm9tF9E
Y54XmtdMwF2MTcLES3tiDVz110oEF7ZHjn/7rHFwWpoKZC//w0Iv5RkmRxozM1hm
MH+qCIXkvugZcdrGsAekZWHCtkNOAXaYjOdPymgR4gwgdDXd+hft9cqKS+35nrJZ
820enfbcD2O6nrtTH7gNrcO4+E69p14I0m05s9w84OSLImt/jMYyWtL5L+yTnHMc
1zH7VJ7w2nRKTogFWFt0up9H+QtAtG39F1/TK79tJevQ0+Wsk4jK26RqdqzV7/yH
f+/cUOhPwPtqnIa7SsVO8pZ2taxBC5Vz7JwHCUXlSXiO2uhPdU3K2lZ5dgQApjAF
g5o3uuuUfeZaqrVRVyozLBun/lUu1R02nXfiE35iCeJ9Mo/aFtdMma9Wwlh2Mfh3
L+g1eYVdaQ3baUiCDCLY2HO6RmzaH80gKjR4nVUwRWcGSjaOy888afXaNvOtz6tY
QimfHYhXogN73C6GUx2urn96E67aL+ytX0aw5VqU7Ajy+6tKVrVFdwcngE76/+UB
mk206v46c4Umalg/hM84nDY9trSfOznZZ53gFZcETxinblvtIk7cAgLkd5xhnM98
j29tf9XcVnLjcsxb0nR76dzLSE3b67nO8BqVYZpMvljLZVHWyUQ3ohAfsnSfAFqu
RaH7M9JMY3i17j2Exnn06HyORDdJG2PGDLVcj2kYaBaGn4hUOP3jAaFBYPI2ad4S
mU5HmfciSgm/TKZ1GLZUGWvCJQBeLAnN6rwKR7UA55ficiRm4X7UuArBodLBAG4e
nlNLV15q5XTRVP/7eMZ42+toOd74l21oFX2V5mu4jm6V+erbZU8ONAUaZfhX+NR8
Ru5btcQy54HIhgrX/1WyUEjOV/t1+YAZcBwZvtCZQGEW/v/S1XxX+l1IyZXf4wyr
kgGKfnFaqA9HixdakVqEbeYYq612uh7Ab9WswMWUewkuXzDz006WAoOlNqWtpAkU
Z/N3mVL1meUufldmRxeAMQT3hoRmNqYXiwXnUOigikUoIKp/vPokuuwr74AYX5MX
mn2SMqjSkjFsXjOaU52YltcvkY/JcbY9DOLtBUWCSiWqXqcCq8/bYjUumSRx6MEp
4svb5U7LUkcfuXzyNxvgYyGRcHHbbCHlE8SKVyHgJazVJl2x21e41tpacLDfamlH
/BHnmCqPjYNWn4gwxQleYJOcAftW7wpHXn6FLaYDHpwuql2mP+g+oL4gWOzEMz9C
fGBmzdRv9tlCHoYohKlpuyW78ySXB7kG+G4G23CSw7Sid6E5lky7OF6B94XIaL+L
8q6ddWfoEJjgdhMwgz11HD3kcBwYqaA7GnFXwMDYas/Ybi9buWL9b5A8ugaogg9u
NmozeR3oop3IF7hfsBJky6yFgYJXToNh41I5qBxQFaI64QRJDVpvlAt1h4vdb+VC
M3kbdosKFVtDQtbgO0IWU3WqAaKGgfzas+YpOeD4fBtkNYUD0dGYJLi6ECE2p/s6
lSe+/i6d3h3jtE01kTfz7q1nLQ80NnP0sYC4qENrkkhg79+zYlpmJbNym+u0P197
3EqTlb8BG4tiqxHjn1jYO4AGXlukb/Ce3uts7opvccr1J9n8hhud4/9cNBsOZQN0
TZw7FHEp+Excpv8HcJEgPjN/mmTYXhptTuvznvelwJZwkQIFhJx7LznMn4yuJ7Ju
vi4SZk5sL/wvx0v+no/CbwpFBXoRHUJStmXJBVvHjjI+mMpbcAFiLItF/jB+wKa6
gGtbVTL5m8F5HsYJfedLAUevdKtviEN0iyH2kKtSY6llehRyvsuuXKy8JS4Xl45v
uDtoXjQhpzy6GDzBaqMiGgQg82iIygB6Csf5S4cfTcIuQfoWg/qeGCfgyKN9ijvE
F3s1OJmdJsKqi8vhs5Uk/FS9PiuD4xY+2JpzRzNGHkmPsUmfgOkHDsjOXK390ZUh
o55i4gPhhPmIukD6VYE3CbBOqllM/ExUK5jF663o1Ji8p30FFJ1pyi/DXbm2ap3s
CUENgOe/QupHYfoxx5psasVRacfyNcFrY1MSDiJnuWHa7iYcRlp1y5L39dMOSZHs
cOw9uVUYFCxxy/mG+2ePgNTmgOuysb5rRt1oZfRNfZX4EAnruYo9Ou0RKX1TyOiw
wzzWx3T1c/FF7+KBiL+e7Q==
`protect END_PROTECTED
