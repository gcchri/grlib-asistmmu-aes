`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nG9CRdoKn8s3T0ORc3K0f5/l3mCP//ENFvlkgWQCLtPv53tbALbxEIMlCxjUqWbk
J9BmRP1S14cK+tx1hqORyCYktgJEBjs/lFEkdScvJxbiZM+nkh4xuoKSz02uSN7t
KRt7sH8yXC28fW6imEwTLnl5N1VQwZCTyd7TLVhRtwEwwZ9sS1ANDxNmMvORYYgW
hvxhLZcJjBg3Zx+OsNNlpTl6NcH1sfszJsVgffjzgwQDyLosWm34rasC3g0D+Wnj
sMS//Pfrkf1HG343Ly/gWx5HTO6YkAnQfduDV/0/ZuO203ZVj/0vCqFbTuwg9Smm
hktzxPP3cmiNZfKOIO96UnG73I/MLQeqVcJiVSPR60RUt+tI7AG7uqr7DNul6bDi
891LnEFOgV+GA+eZRZyFRn7Wepy0GMph4ofW6HzeZntnP+RHHiMU3qLSiuSNLU9B
`protect END_PROTECTED
