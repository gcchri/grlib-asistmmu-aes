`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JAO+vF2r0A34eBda8Y+w09jCV4a0pHE1nrRR+qF493zN/0JpltLGNL1NDpCsO0PV
BR5pYgMhcAQAsRQNxZm81FZ/fa40k4JpLC/ItvxVWMUq9E/w65wMhp2Bsb7CQRLm
qXVZlnTGfrNM+bx/OrbROYAnYGmZIJ6vrLIMXZdE20F9OaOLPFr31HUuMDXksvIx
AW23t+yZ1UhG5IAFqRFXJuK0quaoGPbYjMi/B6QNceFqbRg3STSNukq9UJtlNNIA
7MUm0OeiXRxhZkhqWfNHaZbmkLTM51e14JIoHvNnGfHqs8o4FFgEBwbYNqduLXf9
bxbFqffJUeMCTmqcsNQKhiqs+peX6iyw7jKeOq9NEPdmew+4xvVCRwG75SOWqOgz
2uThmBCmSK5y6LnPkmBZjhkqpynSOj18FaK02BfMYJdBKnXoHbZP18Cm8xzhTBXQ
GNKESzM7FvuBx5Rh//Elf3Pk+j3yVBdIvzSQOrRjnimC9Aa6SpLR10Mt70Jk7Jup
JcBnIHBe14B2SBsnTKoRP/3IOXyroILjmrYcF+7jpQqr6XfHBsyHgs/fv6++d9Fl
n+Ups5YzICgsGCYFJa4rew79NflCxOIhpPAZNaPQM5iToJD+a1A8cNQdxP5q4P1z
qfMfYYXKjLZXu+IPAOzQtu563Chmx9+7YarJCDf3daziOwXlaNPPSezwhfmm2KFn
PVHvdMBcs4U2//9wVhDqIiXd/pvqsec7SP7lJsbUqqO5NDKGyvo6hk5AcmX/0kmQ
q9p+CwTLYF6VABxAOhGgAlz4VdR990UeMmxMw3tkAQmM+mEoIPRjT2rw59RIR7+U
RZK2iJpgscoLMI1ec6jME3m9vlFj1TBkNpvrQHZ0CD4YuRwlnJIJZOyaob6xqk4z
DzrVqP3xuNKZDQfCXmHksm79gDegz3zRqfoGpbRS/jr+O+Lb35teadyNGmCfdhAz
RV6Q+qV4WAok+7C0wtLrXTEmjRWNzO9nr1/F/7kgNfGXnyE8F7gdVq2BCKET5hqj
sOHb8a9G88Ng42inDkvFlXcgMlHbSUFDIuJU1O0csyk/c32QCk+NO9wQwnArwi72
40+siT0dr1kml7PqH93ROQ==
`protect END_PROTECTED
