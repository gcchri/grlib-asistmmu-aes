`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ev5dB1rUwx1s9IGGfVNp9HgwTVk17xctoUiwTPVpIRZjABjPpnEz5+a03zzR+7gv
BNR3fOpdJtwr3EpxUWB5WSyMl9x3GeoiQy4025zXE+d33N/BLDEUQhtlAwcIVs2J
OPxVDXdcxqPVuZd5Az2gwU2LXochg6sA4A/vNkI4ZZdeYnfEpah0VVIHuc6UgZSD
krhm7halyV0xy5Z0tzR4KwFtBmOqW5OI/9rFhR3FvHey6mSX6xWMXMepYl/7s0nd
F9bdYXDoZzDgevnAPkF+dPUG+ZKdHMCkC30d5I7E631Ev/801/rtt3s5vv7KYh3m
GXvJfpaJblWVq0eTm6+8wof0PC2Lm5iI6CAGBXtbFlqUUDdnJ1HjzXSDODnLDj2P
vtv3GHSkmyjuKR5X4AslJtFW610Kqbbrxlc/T1dFr7GfPQBiomQrh1R8bO6Q+/aR
5J6vxrf0v/yu7t8SLkPsiowbKb1Xh59UmwIUsnzHJ1r3RIMwsfSkvJAADM8OcqAU
3DHcUuHKXD71hqT5zyhgbfiOA3g0ZgPsMVClMitMUZHoMyly6LzUtxTvCjY8/ZGr
`protect END_PROTECTED
