`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xbEl72GEc0sQ3sHuAugrmtkADnxe8AslnVTote/CeDbDvxSzk9ZQ/S5OFVd1jKFG
7gmpuY8E5TudUhxYNRpDwkUAM0Mww1tG4k7RFj5gPoumWdxXuaIl+sxmQOblN21X
sKxtyhOaScIHRhcNdDYMECkNgemJGsQhuosFNY7qNt5VG2FwFz3ONfiJs1jH5985
c7m010GAJlvsHrpO/UMLkgstTMSOPjkXawMll9y4oePrwc2NGVQCNnltJXrBV6P+
6nnN/asjY0E4Aqcu79mX+VxRqMZ9MfAA064UthXJ9v8uScp8MFcsSnenZ1SWvkKx
ZaTDqdOuIXV0WBT0XrmV4HdG/5s1w33PUd0hvfQYXaoFajdJ0wGiDX9nIpTBy/Qz
r4ArKtY0JuwWvlgDNdxZIg==
`protect END_PROTECTED
