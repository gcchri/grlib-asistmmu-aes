`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cVzIy4+5Tu8utSh3fDelvyAgCa699lE6lFljD0UIkdgS5JrBrhRfVvkZKb2QGNCb
sZzG9p74KCj1eJzQKEsKbnDX27cxI6l4Mb4JQK246hcwEuMrE5FXuaQ4KrEj95Ji
Uwqj7/a0N1fdinF52FFbdgXEoiOBT5Tu2vLHWgzxLK9HN4r9XEcaczIwWwaZ+iQ4
l93WGMymyQ/9oFx3Rh59zlNiP5Jh6mkRObmWQTIiYO/seaupi5cyQR/CuLLMYyl8
Nuw6UMkscDw4uBSsXuiAM/JR5/KdDMhN16SK/XH6lfaS7XnDYCLKSuv3Dkqki8I2
AOX6jc//lN5Pbg7AnmJPCZdkkfFBhTIRolshfgRQ8rk6KJPLpTjRGMg8NZuZU8hq
Wyv+ev7I+D6q19eWN+nOZCvPz+Ln5ix4m8lz5rkpGszaPeABz4WEJaAxadImEThE
QuRWvJq8RCcHMetkptuULk3bLsPk8aZhXiW6H1NtUb/eOCkJepD3TXXFdGYZ10sm
Jrcf5SOdO+WFWtNkR3FDVO0/LQUzcxEkVcZlmYFCb5Zp2fNEaSc8DtxE6TGEzbsV
DL2GiPE1EydVYeGqWwA8HQ==
`protect END_PROTECTED
