`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pUk5eqd0s0EyHhOzSrFcrpGaPi23ubNYkO19WMZ2IVkPROKGMkputSOZGUDI7Air
7qlK+jBPgdgiy7Sz5qoA7xZWtdnnnEt1V9SIoFOhxdZGc6ef2eu86mZdfPbtXuNp
Y8+wxRgn/wAoZqT8LXXyLxd7bSceJOy4D25CWeArcuUNetqu/pBwvg+l4cAlWlfT
ah0kkLA4gUlQn+tw77i3zU97JtJxIBL5TiZyIiRQPYfip5+IJVC6nu/wAv4H5cts
O8S0iHtAANyh7/HrHcGbATSbp21ybnC+idvLLJnZm4nF6r21j4NHzFqsfTZwEXOp
fNYQsjRrJoC82Gi3LpqpVJG4spiUxk3C032oPPjrRAIHhwQs0kkeIdRNrNN4BsZX
uKBT3RCIpgte1Z6Dk/0D9Bp/vWngWiCh9ui2aESrEXdJcU+gLhTu1QBlI6SiqQFQ
hXuOCu6/5lKMkBgg9pPty8KD0LErcofqH65BPzz0EE1eUxr7d14rqBjnjknX4/bS
d8udrA83X4G17xHl7pi3AKIIWNAVgTkdC7ARe28Qt2M31gIrQ74Ts79lKx1LQyh5
j+N56eAuzTfbx44NlOR/o4SLltacJub+BCDVgjg3AuT3Eyoj620zzVcsCNiksaSf
Val4jlT1KKVI1QCtYfYaVlcaR6+nX9jmFOCHNgtvjtVWEBDsSkFCVsezee90yP+B
`protect END_PROTECTED
