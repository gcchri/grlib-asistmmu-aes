`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8b0nrU3NT9l3HWeTdEDH3CFQGyT3DsZ/CSNigmMXKYo63H9QiPuWRPUQlt1wpG6Q
CR4PWK1qV70DGXfycIhmJJpIRUGtGKxiXlGcp1wYuFNTRAGSyyamN7HW7puQEKG1
iW69ZIWi5iMVyyMxmFGqjLwMlUqkOlXBTcTe8R1aKby0yiWqmXjog0lO4sMI69vh
XZnKJbhmia/pM8dpzdLgGBI87g0xoxDPeeh/1renROhOrSEic5fz0OB5w8JeyjdE
0LNFUh5NIhnAHFECEjEtcF0j1mSvewzjkfZRI+RCsrIyY2QtUZDdY7qBtbVgesyg
i+ZN3BEUOOSrVbFoeRkI9Zr9/ZWRQ8ac1N1nO32ew8uy2m6RlS8+vu+T4pQlbEv3
gqxzsrogYPhYXllocOOQn9UeTFtIu9XK09jzMWIt+gLrtP4ZcdJj/9AnCbjVozse
7DY3aLu/BC/RVevCqgDUcdaxEK64l7w8Mb+h0zQ42kgZIlgDEms2i4zXHoh6fYhq
0aD6uARJFeQ9Mk4HxQxQaHE3mqnImogsxTyfU7mhBJaDkwuQGhXLCbcHnkd/bZ54
IQ3OBsEvvIkQ4snwKrUSe28FN/IOnm2sTclqIZSy1tIx/RdQPRb9NrapeLEnOldy
vh+n9eFGVXx9t77MtknLIDo0B0tgr088BKkdtB9XXhkVgjY6cvXf5BdFcZ8qqkA/
bbaKkpWVyCnzi89Wje9sxg3zdTXxo+fZ4W4tfk8O1k0qDtZadP5upe9jYC9CkGVJ
KydHWc5lL4k+YuDd21+ZuTbd7PS6cG+Aji/GnumYsTdsPYoPCxrhX3yQGLSK4hXO
hH3ghbBlAVhrOQlBMRw0Jw==
`protect END_PROTECTED
