`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MNih6uLmsZmB+yxpxIJtvYKSyue3bNpjKVlYhFk6VJ2RMcToy4aysoL7SehvYWHh
XFz2B5q0mDwfMKPOwN5O/zqPFhoz5v4tmq3FtQqwBtc3evZqemVwHf9MyaRhJyPY
kMHsr0gUWBzwNGH2B0naa3KOOOTgBDqW7SepWc7M+c4SACP3DKgnkKalUBkVzqec
+SN5FUrTblI8gigUXzwA+PdWVfo0dMZuopO7BwUkzVa83EKt/Qu5PgZIAgJAQvem
CzSbKY5sJSAQVNRZOwdSJ4I7BeCB7UiuhjwsepkqNxoKtMCjpeys6GDJrT6IJ23l
9pET+vkVWdT/LjONwc1E2A==
`protect END_PROTECTED
