`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SAvXkLvpSNUJahFJzMhlzVEl5/wyGCc4Kv6GJFxrh+ElIvgxPlbhnsrib3BjJVx7
FLsmXmTaeP2xCUlTSYsQ4+Io240+jEshsIV5b8qejM8hJRot/Yc55tfzQgZur4Mr
g7uUZ8p0oH7f5SDAHYkap+c/O4ojT9Aix3TkfbPHgaeTkN6A6b/dcsh2x3AF9HO/
p8r6Ioyz7QJisduowgBQKd2yAbPqLQlnq5svRUellIZZ9K9uloi6laok2e9SawPr
YjLqsmfSaCtCoxV+ag4soS8Wk4w6A9xVWXONJuZawwUBfCBkgLcPsozPALHb4VNC
YriYoLsyJsMwEZwlKx81ypoTaGQKl6KztzrRd7gp5KFYcZl992dxfI+GsSeuaM85
pl/Hii7cJ1DXL/yPZn2HV7kc6VLgj8T+3hvEozRaVVIyCRBE6ACvHWpiJVZFiPiJ
UuS9MwgLqPYqfoHbNiKWDAnZZtGmphBsYmWpRLXvJ/ftUtykltFDd//nlevX9dzF
KGHBrEV12nV0qrNw0C9055TqTuqJB5FevDOvSN6YGP/gP93aY82Cpwkjr6J+A0wU
4t64to6RCcM7h29gdHwgsGV827mSQy1BJYYn52FLTq8AVNZivNo414PLDa07Yrjb
xc9Ohym0FzMO+DXxQHtmMA==
`protect END_PROTECTED
