`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pSqADAn6Z6O3yR6/mefdHH+2P2vIScpZQg0rSFCpMrwCK51TPk4DzyT2sHTBuz4k
K8BoFKoyctCK8wijrBclB0p////QJPlcr8dfXX5YBA0moiXOZ0fCIHM1wC55aa1T
afYlqdUZrGrdjVBl9Z5I6fPwFGMn2C6yflCrm4ojDydEVF1mpdof9BWAqk2IMT0n
dKfnUTxaG0VdZwwAjfb2t0jrjCu7vnor2tU6JNMZxEAiVyFU3TdNlzB+7zrqx/fk
A9QofUj+88Nu6+8iaK1Y7iaR55ZO+wikwTuNIi9KcUgdsekzDf3nHKf8cG+okObD
ogThC+M9YW8YF2SAVVbpUdrJqdSJhKDuJF5yGc9nsDe3lRlSx0GlWZOH93vq54D5
ao3w+4cPM2qu5AEv1UL4bOogkHE4mf0z1ODwjeK3C0uyFtm0DzFGRNOiItZ7AkFH
SEmkPb1764BDVGn0Z/5FDSxQBQS1diQDG/JZrEpL7w4xmtvLOkv6LMXIQK8B8ylq
FcVKXz6mxQhICeIjKDRpIkza6vIuMlrz7AFnXAufYJOu0Wn/pVxme68XKuNkZAJw
XRl9GgO0AojS+RCyQzGA0/Za4pZyFRwdUNjfahS8eW8dEJG/YNwSJEopcexRB7Gj
g0H0GPt23pUAH7DTR4GuxtYwfEmDgPtssDj7a5JI4CKl2oCzb0WElVU1FCc78/xD
wOeFvzt5zWgl/QQ7zfdt7tz2BfwhkPqu/zsf/L8lxutxS2TJ22YNb+CFBJeODk+T
3pqAkrbRzQw+ec3lIH4ptB03KpuzAd54C5RjZjQIvrJ4iQdOKeq8zQdxQTFmW3tC
6Xy8vS2AxslOefflxRbcuOoUIZrdvjCugUBgXhDLbxkR4whF8XF8jjKg6Us8l+OS
MuWFRFPljD5jN0U7kEBeIX3IepT+Vca4BOLdNaL2q5tErN72AYDVlu1Nkbx5grBv
TCQ77D8u7PU/TttjlRhxSwfBUSDoSbYRXTkF0hEx1HA=
`protect END_PROTECTED
