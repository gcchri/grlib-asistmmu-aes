`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zz+Zp3l1MfhyfLN05C0v3ei92Kt/4bqwmbkxj2WYkpt4bw2rzFCxOy+2lg8U2yG/
Ov8u5om+goTG+hxuaBlxDr9oEARCUysyQQFkL2SxUG75OKSOroKX9CGeIlrPQkgi
dSrp+QkRj3R3s6czIQ3zny3IptlYhGNR+DWyoEh/1lLvTDnHahmQGPLDaFBHWh4I
9RSXtOmPyg8Zhngwvcpd/5FzXI66Lg1gsBxf2fwlWmQeN35J5S3GSpNO/DI5j7UO
2qWFdlaVkVoPiOjn9xa08vc9LliVb31xWaROgQsx68hutzIWDbmwh/GuPz0D/joq
GQ4MS7UEs+5sjSnjWgaeOYEGFftcc2hlNGXXZEKgFrAxVyKv8KcMjxQS5iH8zqI3
lVUZPesT8SxhbqnxvOUqiN7ubWRECzudJA2kVZHHxVfGdRUUZqbx5/SPLUIqp9I5
RxAF9+pCEFwTjTEV4ak9JSlCuc50TeYQq6YcYDnUlidRRKADHoBy2yvxht9PneZr
o/xmKsUqqVirhdCAFF043wNNubvdvxYwqfIISWi9MBSTh7VjY8qb1sBfu21ruM3Y
3WSL/D7qieZ9w1l+S0r0xc08QzPsrN0Yl9wtk8Z84QYujhkrGE0bySd0cL+g1/ul
4QcVXWG93IROw/0F4U4RICz27uhnjUGFVztDwNv0TOViPA3hnj/OWfYQmCENd/EZ
/sIiCDqqFMi/njay0Fz2i1jU6liq5sVtCN8VE6ALJJ0qmZHixBtG+mo7bYReHabo
VrU4zHOOkAxWKjVB5m7934EJtK8Blqshcsaoje/MIEPaXiQMYlC6XWqpUHdo2zhY
Ibe0S7HTNLEmW7gDd+jBCSU9LqjoklB3ECd5AIz45vqhO2rIp/fwjLOinGzGVc3J
8x4xFvxiU33TxfW6PEfme6i/f8Sf30Ez6BB+qeWF5w8mimK3fNOzqaeAmbj0CWXJ
zw3MiiNXSIVyroB/gYba+kRVnKNhaWw6lALDfAaT62I6usf1AP1LJqqj/RpQNDVB
JOQPAF4V0mNM//6X2o8keb+bCk+dPJUF3smHvdyR6cb7nxwoCWb1l/G+ZegE9hVB
SFP+Dhej8VfR1p6Am/NDtV+vcJ42G8L53XqlejFXr/GM+/wYry52t4jj8T8l5jKE
Nx8h8v8jghSyA6lIG/ozrxuMjL9OafxS45Yp6gAVt9ZZxoDT4X/OqBkw7nDK4zcA
Yg9fwlch3s1qieRRPMJ62we/vVz78b2zOC91Dzkf+iqCJ/bjrj8i0S8oVOkQyhej
ShySYRZveUm9QNwLPWCklhU/7TWXnW2jM1VtZg8XyEO6iASQ/N2ANdzFYAv/MvYy
wRRe28riyliS2BK69Zi4yKYKpfNcMhwS2ll1QNfd35zoXomLIWUBVeDieREDKEo1
HbXj4977R0HIZhmTbak+Pn25CwFG+/1LSXQvRjH3sYMMxWkVI+tGsNDe/PBepyHq
h+RiJNwZvhIj3v4kXlthJ9GtE8Huifm+GCNwaAnWE+NUH9WGTCpHMYgTCL+EF/b7
mwfRqzbAsPTgqqoNNq/+dMM1s2Lw7KpjrzUtoxa6q5kMlIVuQliT0nFzVc0fI0Tu
jbakF3pu2VJJFAOo0O6rHk20VTDN7JzLqgSpPgkQbbuoGWy7Lt1AkspTr/FILjWy
FPrZkNjiSKjeU1KECMSugUerHPv0QwdYERXCcpNo6S+BIHps5C1yaI5zjoCpBqkF
0f0HBXeVL8DcHSDo9EthvSOpvHJTPWzCWdczGxg0MzeedEtYkTDgdaF1GDU3K6+I
iwoWyKW/c2v27uXdb8tjiQicUt0Eh8B507wOQszTKh6s14Gm3HqnQTkwYP9jNPeQ
Nr/Of/ZAEORruLYGDhpp4ZNAS/rYEQ/X1Mn30r8/N/s=
`protect END_PROTECTED
