`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5emZK9H0o+pNjUsC8oGsU6TlRqs54/jTMfUzdSwCb1BMMWD0QMTeUfDnuOd4prfW
ZJRUFLClRX4XwBX5I4GR/euAHHLdUuYwoqX3tKJd2uAfN4zxBqcmwy1kmuNLa3cK
dRwCj3hE/xpxeLyt8LgTh3QxUiR+eiZhPhnxzeW5iGfYevWM6Q+BmbYhhdI+jAdb
nsxzkGkGooCpQi1OJitO0IbhDXoEut+VBPMlAqx6BV2eHR1llu8d8xyZ9HsM2Nf8
pa3Ip6okvMK6d9ObZWNmNHWBb0tkBMbhxz4PZsykVjyW08y0IDMgUgru9vUWLPy3
ENf1NkOBQKCpHaEy786lG26/+9ENTSCLYiJjK7uNEEI/R2JS0ExRrex/1mTZ7RfX
PFKSf0m+aFv5hSBOh3A6Rx1UQMnf2EQdThyavXSSXYVjvUzA+8oizIDHB5nXhEqg
Wvhx/pp6rbp7BJivtK2bO8zVz3L+2R9pvWZSxMQS2KwEba4mgmutWeLh8LtmBbJ+
87e3Z+tWF6+AUE0SgdYPwq4yYcsLzk8qGZzRfyw/NN9oKvlI8nCHv64el55T52KW
7kkdv3gWoXHnrxYFa5jiafO/ng8EXu0MCStOWx8KaEyhFY7e9DqxWuN4piqTqMSj
cOPZnHalxQLZ2xUvuOZcOtMn+4qzkIO7hLlK5mjzMAhfqjZU2LPTeOIEtvX/gvxZ
aZf7h1hfzeli7yeiB8E+GqsOquiwBS1BIGNmcDeSzCu6Rre5WDShtP+uhVUb2s4m
1C2uuf+aWMCfQpZrftG2EPW1Ar1iHc1FECxFpzDH30D7A5VcGWw96HnOtJ0zkDMc
ywCioSwF32+BC761t/KNA7k7C/SBgCTwMJhSzPn1o6CFu9fKCvZvG9XK0BBD1w6K
TR4VXK8BJi4pnN2OKtKfXCtaFK4C8TSP6hkW88/FOV0nG+ccA/R7DPFIpQmR5UVF
rUf4N69pYTjgqKdEsD0YWQu86juEaYFtM7clFHemIP/xpfaq/zmzSo+2Q/4Uo2eG
6gD84wKfE5tQrJ7Vs8bGV3cFFBM1P0KzZY7P0jSbLr4b5s92nzkY1H97Rar+8NwU
2E1FgyG5lwZzs8S5GNepvFrbppeAijQ9U2T/1FtBQlC/UlG4asKfOXZot4hNWaEH
uCzyoa1CUee8wmhNeaY2yXLjj0m9dBxihEY8o3bJa8K+9l4bOryh0jC130fUhLiu
zM/aL1iWcBNwpp4CfOPI/pTpFy+ivbHFk41Kem+gwFwiAondrj7Pp3BHxRX+FU4W
MuIoPa4X57kYEqWUpAoE7RQshyek800RBtftPmQ4xswG9IwXBL1+zwxpUYNFcKtp
pVVMB2t71uXTavB+OUHihH28SDOr6vAekZBaeWKhjppgoqvoWH1vUAAv1YUCYjJH
RJ5Er23079LkIIGoiJZfCjKVpy8G8LjXFG/0N/WH9evmq4kvYoU/qgDCy3NjB/ib
JY2AO2FvIIkYdoh/c6CcevLEmRGV76y1iC8cnzRpLZp4eHO6ttw93wk19ei5jtOb
BWAKURqEApFRapSlSnpuCD9kSXIQ8qYywPuekdQpxgti0nA1KSe3YlB1aK/FJf7q
WeLYN1umIKmMJC0yZH1NpeJCmR0ldOjIgWBq8rTZx9w0pSvPz6L5jVTzCueEBA1i
UX1rda+gFIuEFTqaB2qmOJS2xyFZAXYYKldgmc/MMgoKFnyRYM/fE7WEZaiJiQxa
94Z22uO+ZJ2H/P6l4oZWNL5feNKnhtGecPqORfQE0lgpvgFveQZCgRIndXjLGDz4
sUGI9dktHHHL0ESt0qSSlYDDW8Ben8z2FXMirPyew0/7gnkd0ciI0QjKBLkaUNVW
LSy6cTb2sDH3w1bTgtDwWt3+ef4783p4BgVH1PSn1CcJJ1MKf71E6f3aIy2ve3om
ShtXsGujNnPgry8Svnpa6bOYyA6H/gPWDSaTE2KH7gqMtExEeb2ZyFjWeHGDC/01
7EUWmhETwRqt+XdWi3EA6VFmp8kENND5dQjtQ/hariTcm7B6LDxFfgdUYom8j4VD
BeNPlIICPNdeMSKlS3PnOpgGd7hlMLnt4IeW7VfEbb6w2QX4jyFKy/WycZoHmsyg
1OdCH0FjdR7MmdZhGHpnwOtylNxIHZoo5QJFFO/0lhJLHnIo99UYP7JvG3B5X++U
H9ctZG2xLx2SLOqIn2OnQzxc1Sup/zNMsw/5YXb8TKprCIrcsWLH0ncc3vblUBxQ
jIh+UrjAFxyvt+HaaqMgM1y3PsYrXIwL7M3A+eo4bTPjzNnfQzGxn9XhGrcB7kHb
2OyKGDeI47qgWbnfN4JpxKD3ywg9jQYPJFMkfTR5Z51HgmBUrCkd2k4rF/xb23c0
9H4KPAZKIiJlRj5ly/eIkNXEsR3ylbs+b71cBXRxM38bgItVolNLq3lAndt9FbWk
TeSPjh1tVsTVSmqT3EaO7jmwhVE6MChCgzoWu2Aa6b7vZS8HcV3RmA+UMQYAjZWI
2ANKnzi768BZQWHxoMWBBunqLrW05KCI4Zr0tk6Ao10=
`protect END_PROTECTED
