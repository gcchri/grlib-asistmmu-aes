`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+BjW3dohzFtiKI5zvq1o0KDzL9SdqshCOJrbf2zT42NEh2vp1LsxkZwqYWBXEKsj
w0ITbwAZgASREX+G1pIB0W9GH9rAnYzDpH49WG/azOgugloFbbFvnaSI3GHQbfEs
+SmJDhQ1aRZtQ2eyrvxGGQRMUa2OOPCg49UtTsNr7qB8vvpa7Ywz9NOXYjNNQLZu
rYmLnXGYIfl4G19rrks2lUXwhrXI9/3ZnsOruc1FN3Ds3EPgkkIeqkRV9fm0cEFt
1EKvGKM2KXoeWt2yVmq1o9WP8q9CbVooInuCoFlFPYh52vglIq84L7QmzdJX9h8C
wx9cfAJ0jY5VkAs8aZ4t6w==
`protect END_PROTECTED
