`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4EKFWhdP498JNY/Kss7m3TJ8RLY1taHbDXye230jkr9glLzts3ok9qz/nMNsgGvL
d2Y6g1SnHtyLXV06Mu0s0ua+uts9mieUrJBIPw5pZ9phoJszBvCWAIKfYhM2rY8l
mGFFt96gZW9uSDXW680Vs0FMNt96Y8Qy/9kdYg2ZhJPrBA0mTwOkx8LzutLtbFWu
phsskQ5CA7nMp/iXbs5B+udchanck0gTpDWarZevDWmwNasF8sAWuVYgzcvMaaeg
71/SoXk2jXqbXXh0wM/W+JVkAUsisdbyA8MhJyNku0vFAyR7dc17mKRFlAWeaulG
asaVt9D0l7SjzJLL/WfAl2KyK29ZLRfn/EoeEWOxoHN5xsP2gmqtxSyDLEghWzAP
4U/bzVLNd4wOAsESL7CPtKOTlswP/aI+C4r/rSS1VtcyepPd5j6uL9BjNb/ykKHI
XZgQMePEGfXZ930aKXBoC4b9hw9QVD/lGk/VaSXGNwGWNmW37oRz9ZRWvTb2TdlB
zhJTzRe0fn+dEEfLqVWvbTv7nPqgNFuH2BxGGOx0mh7yz3nvwjG9qmGmyfTqOhqv
kwHjM2LDzqEmqHcMP/aCbUuKm12mufDTkYEZ27l1N7WabRGLGelk6lyLebVJsNej
Z85SGqQCFo8HQ43waPRnUu6Cm7nbLDkOq6Rscxobsg07kxBlewjeIIS0EEbsEHRW
bKj2LX4cdmtgAhDq4ikgahf5J71H+11WC4NtdFGAHlwbNPEmK1ZsgsCJrEDltsjB
LxJ14PmvyVsPn0UK6zZM60vGmVp7vTRKE8zuJXel2WJnnnb4bYZEl5n4pxYBw2aO
EUmI3oMeli5uczv/+xMajgqMUGEzbP1eGt7tkf4KzYNMRbcDRT5aGkUzmJNBXKZj
soSoobVno1nBoe3cC5xqRg6xbB//nHLsQXWlK+GqpN/Cb58mSRrV4KszEEtME4Rr
mXCnuPxyKFnzkzIBJU3JIdunvytIkNidScZ1RAtJwz24dyIpdamNl55/I6qUHbJa
FBURkVF2qSSWKAEohC5k0J3DKW6QKfAlxQaJDtD95ipaPbg/f/N9rrVCLsbSJWUy
dMEJRaY8kTS0s7z7qUKp4wftmiW92GNi+jcVlxQNQi1wtsWQ6ZcnKVG9FLHcGhxW
QlRB9A9J+iutVD+xzJBprA/ss2g8EpDSGV8dyJAIbCs=
`protect END_PROTECTED
