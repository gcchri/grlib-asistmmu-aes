`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rFGVaqkAcMdBTMFYUiaqtXYAx4gTe2yo2bW/z5TmhfwbLFVHDRRwB5BWj37IDF7a
R6of5fMpyGUZBgjKEmpjTZrHDP0HWreR5q0gy29jbUYcWgk1Hwvz/85gjbqjGSSq
mYEa10O1v3l8Zk6IDNZEYIdPRJrB0s9hFdssOgDFzwY/w/XESkquMAGbAguxbwf9
ZdWNl6B0ckjEvIctidcViN208I26TiuvsVog++JERghpp0o+GukhVaukSCk184z5
u7gJYiRD5bEDtYl1oV5tHtaQ7lTpN3Xs6Tn2QZUQ7b+giwbgJcaRrnMirOMEMVwn
orawQDcV2qVl1q4TOL237A==
`protect END_PROTECTED
