`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G6LGavZP18N0Lb/m+BDVgtYM7vaaAdDp0zQdHZLEXRXXt47sfFHtdJ+YybeoXyZp
lOwqUHI8C93CqF8oIbKetrfPykwI76nqf/PTZc3koGFN0+fwfmzMo59iFosYBFvl
xNheK/POco8PzFtm3cRI0LNHLLTK7Hgd6qZWfDNOF64yaVYAIRUjjrtV2qwpc5lK
G8RXNaoi1cZXyEEEsZBg1aMEbjjvcMBVVETmxSPyeg1XEz7FkdJHVSURyFH4T4s4
WllY6/kc0XtbQW7NthLP0zIYb1BPV1HzZNcxxCFs44sCYoMt4UUqMhDpN/6leU1M
NP4GzjanKMfN9z2rXhZim26KBoU93j49SMeFiwikPj9a8Us4Pbkg6Ld6Z/m4SN/z
5hLSSQJeyd8Pr8PV6UhaXw8esDRWSYhMCxRVGlWqq5qNbzRTd9rf9Nhvt7Ja6vKj
P+GOqy9VbxYi7cwWcjpQ4vcqO4anIFknsBvVhk5vNtqp0/hV42suOkQ6K1Rybo3F
mNkqp8kNJt1WFuCjpZx8dabKIR7wbgSBQfn1JU9kw7Edo7xJCqZlMWoRS173WpvB
qZK41XGX1swptNvSrcnKlB1l/SKpJ3cb7cFIe/5ypW61xAM0fKU0XvjTNNYhfPqj
DJVZuFUHUmLrjbVcQr8PJJLvw5KaiEH/WzLHsjuxWNUVQ3kOkBExzbzoYKFzxW5g
bk7Ikj0jheJELSB3Vb6Hudkfu0QyI84LmNkL10hCn6k7gpmbN1svTh9MDCbRrNh2
h4FbLRkGmGyU/4bPYsYvO7ntpYcR5F1Hgdwb6AvQPPL+/8pqrdNCTth7xQFVBzoq
Xe0KgpptfZGGjXb3VwUgEipuW7TwsBKdfKJAQziYZHH3JHIRXYuyQEkkynH0CfFP
+wzJg2I117PbVObM1IimGjgWk9KexHfNY1WsbcXVvP25CXbcWpmFh/00Nzep031r
13HvMVZHrXcKpyHpfQyZomXRDiRb2DzhP9zMVn4kIFOpKj7KMOXLQEBTRZj+nSUC
AWvLdToAGGk2O5R4T1452elsAAfTO72gkKnfk11qxBX4Q/6HpeOmjxLG37zwAEfR
`protect END_PROTECTED
