`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jkWZi8CpMpIQVQnKlg53WIyciYM7etw5Vaz02ooTWPnOTm/bf9Jymm7rGfQf26hu
9E29wmNcSR2uk+o/h+ww7cY5Ap7Mdd8lDSkFSOSDn4pO/ttNODy8bIHVI2tWWag+
ggn8/y16A5qY7DQ/8QYwGavba79nkCaCkBE5NRZphku/WUQXnb8yIAKzyaS5/iyr
DsGnGEujAaln+9wUMJm37dmLQlK9dffZHCu6rSdWiFlLXL6zJN6sg59eYb2Qshap
09kiAPe/HAJJUoVSQEkE1Q==
`protect END_PROTECTED
