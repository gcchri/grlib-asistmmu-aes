`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bbsix8AmD8RPpTXelE8atraEcQG/yYWqZKq6Pq9cv4qTanwiDkNWIP2Qzp3HoIXd
VA/jilown9nY8+JtqGIuT8AN9tm+r1ll0NZOg+rdXQrJfopWA1Uw4sxcvLm40Jfd
n8E8h+lBZBjhX5u1/go7YBBXm5NjlOKKthyF/16R2uC4lYSGPjoi45gm8O3JyaB+
+cDWmg/nbx2UJ6RK7haNuH5nRd5Q7Vb0u4LXjOtWYtNWYiBHNhvdWkKvbqSTMwAv
+rkiZkOPdxu5TZZGCgJgpKaWGbkxQ/+kQBzOnba29Es=
`protect END_PROTECTED
