`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J8ioIQKylHXVPwiZQA3hg4YWBrpVV8fRuVNR+TZ/XCHfjhsOd5MroJ9YgUkwOKuG
PQgQVV51z94BqBU0urxeLqESvGOuOkALtfl8V/OeTPf2sk2/0vWGPoxJKtZYr4Ak
OMVnI9yai+Xj0i1nKFf5lrVzz+THTchkY9xZNkZrE0LOZeEBvBkT7XLEYbswes59
YizMnJ1eLpTOoKc3QFcsd2BFXEQ9+sD0eGEQIXRcqj/m84cViNI5ivVoqGIsqR+3
vd7xh1uls9IvNBwm8oXoAm7CrBVGasT+Iqj/m6jYnv3PD/24rh+U/r3hFZvWZn7b
0lwYxZxWzFvWJ2mVYOdnQy9rs6RmN+VqAfjW4LZ9VjavkRNWE4MPD/tIcb6uIwzj
H3wdZi9zDHPf3NUB3HSlEKe+hmyC4SBQlEuP17qmMBGb2l05P9EqZXvSph9kZdf4
2/optd20q1MkRpIP53VA/YCBTJWygC0EYsvvzgdz5R0p0IdFEFCnZKdKStCA0Xso
uWQJlbCHLubkaz/fr2EKhRzqclfAuEcirGiYTAoJ0R9Fo/xQce1u6ZYO0HKKYJZc
tg3SAsHV0aPiTmlmpxxjbMNjRJYpVLNfvSVmvvdkkbuCCkbbR124K5073YEPnAce
wU1EraTkbTaqwVeywYgKhkSTsJKAGz33rw8yYwRV+JAukfjoCFcrHRSSw8mgfWcI
v7lWynPCdwibRNt2wn1zamhjelfu0bUSsfpwrvaRP3+oTKcesOVLh/OBksPtQyhk
H5883Serk3bk/UUYvh2JbuTaiAoY31y7iVCkh5VA6lpj+zrbDwDW7eq3i2OkgpRi
KArlQ3zhRae1pmOXNh3UmrkcMT+Jc8f7yymQWLLrjSHORwhQcCEuZu7phQ8G/xG1
srwiS86twOxeesCuRu6ZWlOxXXoDcusgB/jF+A5RK6Yu1uZfhkHt4/AyJmUVl8vu
A4lsrUyTYKDsbuXhGhpM5Dhvu4SbF1Ac7rH4LWrSBeSuZfME3DP4jzT0tJz1FmLO
WBXVCPfS94ma03DJwRWml934JRgFE12vT1rE546qAHhvPO67NbRO1m+3eMlzy9BG
bOrx6k3xe6Hvn4GO6hpg+8tfqhJKvxAjLAV/faI/Ll/CJ/bLf1nLeMcunSB0ytgO
P4vs2h+4vvRs4CgkCCY9pX4IbJaNxZdI60eEvlxxGSDByXedNNY/i5kH+++yTTIP
XHHxwwVKdTARhfzVzEy6n5PBSVI4CafSVXjhF/ZMED7Wz883peYFA42a18wGUHhP
qZHi8jj0pGrpRkSt7+zb9EIXAvnnukvN7fiydjVgAISWFCr8Yo+fK5vUd+fES0Nm
6+ks8znbiY6IUpI3L/a2+lGwhNJPCWsuna9Mne+nZA3XtAgl5myMdSfQ6RiV3PoK
/5UXo5KL9J9bOcXuAtKLnHnd/KLMVAyx9pVAjU4STAlmBPIr0gannYmp4Vpn2YHo
bPvg6bhxsyvObLQtEHIIUzeZDae+uvy7I3W6OKxHxQSF9leGVK36uswcfhGl51PK
wHXs3aQ46RQW++GRDIiZcOu1jFOc6YcSOwI3w2wPw39QMK1PvhrfdIfEdd97eLAB
4AagGeUuK/fJlEI8QroI+5rOrOPxIcvMZ7xCyEk8HdtuQt+T04qlMjFrooXiX4CX
WUxIOFGLoI975nbxC38ealr2KLT6zddrF045UFxFB0o/PZr7Mf9aOzUQqcsJHkGo
faZ1pL5iXERn+JjkyuHwaYdYg6tpkgSkmnMrJVqyB5NRVphv7aQb1kduAwbAGbWX
VMy58wyj17oW1vx5k9D9+9ExKwSlVpZCyZM1kRmxiaGnWxV9Ya99aIrGik3rJGQI
CYRitJ8R6xLHOBgIZF1sSDL/KJrALGjw30QQZmzMXwILqpJn1NU/ER/Pz8qWmpkY
NCOgP4EgsBW7MVofZEQv0xSApVSf4IHFzuIrgvXg/At52xoxnK/zZgKB6L9TmTEY
kYwKLdZ2uNR7/Myb8EagJ8syS7YA+z4goA/Gblsien6Lc1e44Tdl3WqYlP8mHKfG
OY66Oc7qnB9r7KSvjceopBheRlOT5HSww93tOAcSWrtSGKgLSIGrx8QUkTrxe+zL
jhk2ieVfKwSj57rO1n0A+WX7pwyBc3cpEh73yOapONs7ZrFazsd9PteJuaoDrker
UWoJwq0xact80L9jeXqAO5nEshu5yTt2yA63/IZw2MJJ6j+fkEUqdvotTSkH9xhX
SfhUCKtIkr5ZoOP+K4YKSkHyc6F0rImqWYO1aScNTNBVTocNMM4Y1ShulRgVW1RD
GwEDLXbEugWeG1ALrzUqWDsQ40utrB9XcrqcSzFmv1uTthNm808I4JOdeaKT1v6N
/POsoGnLBf4E5GHMjbiO9hBwSsC9mU7TslqQSEMUXdSaguLhhfunt2jUP8EOwFLc
mble2oaYX3Vw4VLR74/iP/5CAChdWg3kZXe86pPv5FdYM+M0bFwYnROz49mWzsQh
Y4XW6I6SlpQGkBlbR2JfJjygmGc6JPKkx/SE/rEyvpahvBlSfxqNNNVk3SQ3gxtU
WpMumOGsNEHPQeDRj+aLnmHmosZobEL1bZC8imuYY3HTzeS3eQHqDicMjr7RGJF9
gSWHIMPtd3galsALo8NtcCJl4P0T0uaaGB8jBo0uPU4BXcwXcrruqDTQUnGZIKOs
GCCGxWAVL2yb5/uS9zEmRRm7MVixFtHw+pR186cio+iB0s0aYKNijXg2lYPjddI/
zwJ+9MD90j2lgbeLuTv1Zhrch0qFMcwyMoB2R7Z2RyeYzaCJA+rkcMQYBmLc3bnF
S2mSkwWN4RLqCOUtMcH1wmmGEkdb3WBxbH11csVv0MD+vsVr4oY7NLiIpm4UUA/m
I53VT13XSGUUCEXwx4l+sYJihEDKfD3EF4XC2kTWDqrrIlscXQaxQF7L2pwwbVYd
otDRQbY+cXgRfhq1l1Ga9l5+QrLFw6kWi+vt2nNWO9p7uxM0UVXwaFRkait7Rj4h
PQhblHNGyJU89adc/9lQvkbEHlToSvZ8RuAJpVE+2NM6WlOTPHTfYMKVdHXhFTwT
FodBOZmGDqoBxJuzpwRCz/DWQiQvFJ5PQ1zNkeyuEcSdn7qJtv/XsXUwzWKH120x
ux1XyDHQYwR3/cqghhsS5KB89ArA5hmk/9Njv+tYyTtFPYwZnu9sGHnwsNoZcrb6
zFFQRE4CV47lO4EO/NtkzJQCJ2uAs5Oqhgi9/cWD/6AXW8A1+y93lQtvhPCGe/uD
jpAkDsCGxRUueoSRhmQn59u6EVQim4QnioukAMKVAoJ5XapgzWIxkH420kCT4gUE
4A+9g9OkkBm8y58lfjkEzVhXPnA3KfnvPTu4BZ4WEOSmIcdXQzfRKBbl10n9QXcY
uiUQbMP32eZAnRjQYVKHGI3hY2F0c0QjXE0ZYJpPHVm2Xlqu+aaQK2BqCs6rhRKc
cE0IKTmi3uhYaP/fJ+AKgN9tgLWR6Q6lvzlfgRcMTnMeke2AAN+EK5uF9xAw+kAC
qRYjdez+TVexF5gOduDaHd4fwsxO47uSRSLZZd7ZZfSETq1Z1rF1r2Z8C6aR5P9S
zRL7dFn2lFqeD5PSe5w85iusRRZK9dROC6dJPlYl4XpfYWBK8N0RoTKBYdivdE5H
h/t08dG/3Onw3lL66X6w9WN9OrJhV9XInOGJucQz9Y1eHQrNm4SQO/y+eVcFekiB
6oFV3XEiAo96S15JukoIglYuX2aFy1iKf/8+RWsPJBIaK3WrAivLw0ovbrK3lbnc
aCVypFyvhvXCJSDabskMzSmwr3NhvyAaabBXvQum8jp3i2AtyXREZLX44cqivmLF
wGg0a5VjC8n7tEF5Lgb7pIjxwFAeOqGlnf0SnH4kJtE25so4zUt5d1sCCv/GmXW/
Zi/70Jt+4VyBtchDaSOAs/pS/uYaeGlIwo2+PMNnC9w+Tvyv+RXcbAAhM+D+JuDn
cL58rHrFfJSeF80T54TAYUwUUN9L6vtd/t64todF21XddKaOOuo/pFlJRKBJq9k+
w9gfBYrJIPkids0AlvueUXIaW+qWzqcoiOKdlLSmu9Qc4HMZ8GrKEhRau0zegslA
zl3Rc5B5VZfOkJpaxvj7ZoQ5nuSopWI+m4OlEoJ+eJ+UzoDebrXu93zQzWWgWJoC
jBuyh9l92U96PHpsJqrK32Ob0hhIO/Em9rNqOF6xsflZOFZUbcOkdSUnKRklSzcV
K7Q17TUV3FzRpsdaVKQRpRCtzsQQ/cjZ3CVrf11YCfiJZobOGBJWYrYyuEMnGMUx
VV64TVLh9ezZqyu0nR6K/Zw0Ie0u6+ifO6qY6iipm9Kb7yE2xuci25l0mE71LyNE
/ISDUWlGkt6RulTXz0LKIKIx14QoK9Mk2v6rPb5k59qLqclzM38EW7cfnI0s+RjM
aCQ8uVGdDZPuVJoFG6F6PEbudS5LoQjCJ9v8lPNdzEPgMu6+TJXxlzF8ONvkEAri
am4HNunPh4OuZWVjXzh7LY5WkLIeLfoMUUsCRd5bFBrjpZ77/rjU/lPGuoMC0ir1
cs2XBKqCv541BRNW4xA5RmHseDaNncoh5DQgBOXYyOeakdaqmFykEXRnpgaVCYdI
U1ERJodakJ3OSMegJPx00TBm9qtGCbnEBh1ed6qsKOvMXGHxVcSDjop0d98CZo1h
QWdMqlrhtQyEDaS0Xo3tQVDzo4mXF5WpX9E+rB0OnhK2HiWtEuh0Q+SK54+sD644
yO3+FZpoyWFXbmOITbUid9izoevv1nERvbPsziiTWIIuvRk7Ye7inYGeSd17Uglj
8YFsqRPlJr2EcTzMcQsWtVMRqVZ68j4tqkWWpVG4P7yDCtzH8bddOzXCft5IZLne
YU4mw+UgNWmhy5vtZEboQTrMnivp4EquvRQYQ6CcdSrdnL7xP3o6Q9xeHZ4zc+ll
geTTUhx+7jiT1hsgNCrYJdgpUDeBzQpk9/b3eS3Bxbp3/sVAPffv2Y2gmQmwXocd
JXS8zZLLF1Fv71w7Rb3VkKyKPWxKz9ZMmz11gMasKRkV0BCpr6lQscMaOMNSqJH/
dB/Jf1giwNl5YD21RLDPCaYXkHSztmOQOnE64Rbft/5HtmKyh7WiGAB/psM4VK0A
xOAIzgl1bA3LsBQUZ+HhFvJlBfrmJ3kLyv6JYEX62LC9Bq4n3l6riotl81gPkwd/
dgCm29snd5AdNjliZmxijq8nBbw+VDtYPg9UEt9FzCd1Y4LX62nsWQpcTHwr+ChU
uTXcCzmup59yIGYZLW3l0iwOZBRZNbBuOyaNuLHbJW6NCDkWy1UUqauGjcWHkMIg
M8s5U7SGOg4i+jOxOp3Ew0av7xTqH8H0pGUMc008+NfhRqQGNyipN3aCsFc/oQR6
2xaSXqymX5brLjN0P9rdpCzHtRsa3ubajac1cf/GbJVa6ceUv2cmhYQDDBR+8Be5
vDr6DvifSGqZkHuZVH1OGgNRFSg5kxVr8qKIbYMTDE0y9EMJd4f6iAB52PsUYY/q
Nul4A1dVlXIBVkqrLoyVwA==
`protect END_PROTECTED
