`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J3BxUQZTt42GDEMtURWxhUACg11l5YSsqBxS3lr6ctpwIXlB2rA7+j+aTXChQyeU
FbF+QYijfjWQENch3N3gkifUld+3QZYI1VytVoBXmARgdAPiCBKSJRKvwgo3FVEw
f1MaDaeUe6PXWzoh5OiIKijNOxIpDDmUUCCqCVdTv8NyoQmCO+B++v13NtxTu505
lS7Tvt0BRhvKdz8FjKv6TWcJPvOh5zbXRK/TJRGGf1LBFYox4KI4MYr0oC4x904g
AeaaFv/fxRr6SbIEN2StyaPF6AgJDx5yYMsBBpO5D+QISVZE7oOt71+SzmWExzNL
+UmFzxd8w8KKQSWljyfMLtClUy2ERTWs5GPKfps8WtdcccmpD7LsIQ7RFje0s2CW
`protect END_PROTECTED
