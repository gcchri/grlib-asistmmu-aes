`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s5IZobxsNKeRFfDY547ZLtbj/E+pqRuUXWYaPqoVUHJRwBoYLLrj8w+5AQw+/0jB
JhPP1rAdb036VbPFpKiGVqFOgp1sM+CKwfy+7WAIrUBViOAv0LGhP8HxhcymNEW4
lnyZVKhHJaKSwU4SOPomu+d4G2dil5BLFRbaBCJG1zj6QuY0vGya6x4XYXihEkN3
wINh7pxXz0XwNpBur5JAnE3jDDcWtVa+7YcuUH9vjPsQ87BJK8QTCbtoJBSRqfJm
IFrsGqgdCMjVCnWc7fX+ab7fZsYzxtU+tjqX9ZUsT9zPLj/dNElY1Dju+9wi5Vin
NsHoZhdRu78VJvSxDA0Fo9bs5W+uRQ/fr4vWEQJT0wGXtQRy5VboVApNwlvEryr5
SbBa/ScntP+b7l9S1KgIqHRsGf4H25jyX9c4uiTRqHWJFoGJ+jWYpqZ2SgB9cVe0
R93KbkgB55o2bIC1oHCRpsA8hcQL/9cF9yiUM8yw+rP+B8pAdQBPwTFgp6kPisiE
b2/lfB7cfA5i0dnwCEX9XolX/p1ewCIM3loQROmH/v5LV7n5EFtqqJoRB0Xhuvvk
lu4nwGZB2bLm0bHEo2zT+NNEUIZmAqtCWzIknGn3zKK53/MvXmOMG/tC1RuRh18/
H3fRK3fvsKS2QvTfyl1Fhg==
`protect END_PROTECTED
