`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kT2ANg07qkvAWXVUU3ac027U81EjfyY/a12SvWd7/MrMKlq6B4V6846U9LCM6tDC
qBVFDh7B5trA372fN9y9tMr2Glo7TfroOB2njpix9g1YKO4lxlyV7WMTKyp4+O4q
E4RF4YJ0B+jnQ65VI1W1IpLRqqjEb0U4zq/rNYlr2pwFIpvf5TBaKsC2fRo+TZOS
aaCMjobux+OqhTBURFEJKIR9sqGOgoB5y57v3qt/MGQ3XpvTclrFrhXFLdiTLj2w
pj53aQmPI5E5W/NZWDCg5qo6nuetwJDb8GtPdBE40B9sJMyzhszp7vN+CPazh2//
w0Y2k2BsUKI2DFrwhzmW01f/qbTEI6yq4ggUgBZjEOo1yfjWOS37zW0XYVzzMRs8
`protect END_PROTECTED
