`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OpKHdtpd/w85CGkvrIV4DpZRhNGlicslbPcH7xuWG51sx5YiYCmWGFqknCjHWnan
QIHv0D81iXy2E0Au6d8Zpix4HRtzcVVsovlQhEQOmaO86qwUoeMIPI4pvDyfXbTR
FS9HKTdygmfHBUkqXoD883g6Hs5/XHZSQnEINDOi6kAgKMemfKh2X/cmn5YWw/uE
a7ETgb2bp95h27MNLvX1KO56RDlweohZlFAzZRDdGdIxUJThRmYlTURFzCsfMIr5
DRlNoVrbxYHRnYE8kwYNIqMLo4T5eTI9HTVA9IKJMTkA9PZT6jA8hs0Q/wr2FUjF
hGgXOFqpJiLLcNMmxISxhiJdOOrC8I5dcMMfLcdzDhKBm6TptFrUL8zI0ZeLVQdQ
Ws/dxpHYuNyW/62/iQT2EQYqohCV6f8+cYkTIs+iVe0txWvRxxxTNL9E3j9nnDH3
hVdjTosniriJ6tRzUK4ir0ptE5ffprB2bPzx4N4kAJP1SRiCHZty52sRRtYuVouw
j99SC3RwHRunu0URS5Rbg3FHR/pNAjY5B7d5hsi/0oIlXjHxiEZKw7weN0orQg5a
ufPyXIxa7sSmEjdIIi2ou/T3QYw6+/KlrWXvlfjsk4SavRQwMNUsnYnNxUIAW8hF
aSmWWPu0lSchqNIQVN2XFRdWVoLv7YX534l7jBKXOFgLVxiF3/OR2vcWaaoj0A1H
dsbmTEJYNo8acFdNtI1zXsUbVOzCS+wzF0A3rhiQX+xuAIUA/BnossKSfG9ZpTVB
NfmjsmD7NUy10Tk5w9s+l9Ko5uLurWIqH0aQPHTq93By2YsWYif6LspYr0f/Gg8r
527M2HhT8HJui96nLYuTXr2QUOkXDC6RC9jcaUqZcTO+dUMrbWBIV8NvwRq7rEHX
`protect END_PROTECTED
