`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5j65V9+exQGjL15mTMlop+YD4lRUnOtahZ/HBRBMUPExgqjFJONHQmjgZEI0hs+L
MAFiVpDgz4cP+9jObKtBCM+nX6rcKr8nnTAGSdn1xFacCXl+KYb/x9S/lLAJkRzw
uwgmzmFVkiA/JAtv4yjH49DGasrKMP3kgzhLPMrjF2qts5mS02GE7qPB5IsAo1ZU
3klZzfaYi+dTPHT2ZDxiMXEqaQvZRAA6GE0GL7KNaKNDEz8n2s/sjUOQGiOIZUoh
OYsFHFYZkQgmYDQMgNaOVghX8xXwrpqefpahqbYXAp+zMp9O2BnUlxPL8eY43xyL
s2IhqxpjpnEcFZ0y1qu74YC62IhLix+4fPRoUj9ghBI=
`protect END_PROTECTED
