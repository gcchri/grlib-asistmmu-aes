`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lpelN6xHFeBva3kZfs5WyBrqe03ZcqZXRJvytq1GzbJHcUbHJdLmRmjfKzBt/Vw9
MaiQufvrOLS+J12QjtqmQoSUPHD4RK+hA0vvPHRf95poc/jphQF5SwvDptM5f+A/
rXtFdJJwHnP7gM3cK6dCT8OOog8bmFb97EWASjSLedHU0BadIVCPnF+f/qSSQ5Ya
9mh5o8WcjUUWSrRmtyU87B6RhE9wi+OCNl2w+nbij85hi+ZxUDZH+c0p3Ychei+1
iBD5o/WAc/sAEwoPUZJkPXg56m2YFE/NX5um+n1pT4sD1FHStTErKRcMgaMGxqY/
xo7X+aCNXa7Tii1EqhXBIyGCz4FL7mWW77GOZ79Dbx6KGCjZOjeHGA1m83+bx70C
L9weez8aF6CRgvwiRXh3vCxTChY4goGZVyCb3P4ossTSG9EQBkrEDky7NNrlgGQn
ggffNCJ0w8qkOqJiRZFIJoQGdmGjuwUf1w+ix3Lj+2yc7Z+INvOwXA2CWwRxw/PV
6CdxU4rxYhF5SKR0tY6ik7WKqZR4SJF0gc4OzFQcvxeLnur6DXJICvzPWOemqOs2
B9xcm0SFt4PpGL1fCPS1jEIz6pL8BPvo+bK6ByxPhERVp+/l8IEuPDcl87P+CspC
AqSFTM5h6wZX1P4GXEGOuHGBjaSjHyp03kmK7LVV0X98LljIWk121kDwhyxbh8KR
kcGOldTxFmxaq686Fz0MM6oH3NhJ7HSY/QVkB1a2LNdSvOJ6mu4EJVhtBFHs33Lj
ne7kuquXiyZcyqoNxgRWTA4yJXChH2tyjPaz1+hbVmJLIXDhoAttASsxzuaP56Ek
SqhuaX+injxrNtKL3CnKR1vVBSwV/MpqL9dVWesbLmWIc1/oF3QWypZvYtLSeL4H
FLHDoXcx+zHWO8nZCJubKce/EIsuRLkLI4wGiEHKDL+VuLVEMmrkYVlWhRnQEzFR
UUEwtthTCcpXOV+ANn5FczPLh5bcemEC0JELo2oKVrfr8ZgX2irvOmvXMCIm369J
WUZmDws6OpGYptUrGqPnkekDtgfDzWPX938GD5jWnGwp4EyaYSlDUWTw063NzVZm
RYrJEgVHQVkBfePJUUx47R4QieIzqtZGxYtElh9hmI2bqs1WrcrD9hDWVbHMF5uA
v2UohB8ntg76vcA5WjKI2WZPSNAynJ7gXtyrl0JCpesRy/MJjGEiVnB2DuJBQCN1
6hk3t2b35EW0rb7Jd0UvAfU/TSFStBaWqTS7nLE98jjnzRQYOTkTwqXzBMsLwt1e
qNcFLH42dSX1sxeHAH4F6cGVG1SKCUx4EuSdH15Tef4=
`protect END_PROTECTED
