`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ccfU8b/A1EDDqR9FDK8lOkqzSvF7JPtTliyu7y4ZhHL8meOugeXsdhRwjwENzHR/
85T452FR2bLNnejVDuY2pYqhAxkFf1buly4/C2Qowao8xHn+melRX5oP/3ThV5kD
aJJRkk1Du2A6RwM18SKqOY6gNqXBG/hsSlIvb1uLr9kKPAP2z4Iv8OLVEWiAfSYF
QHc8GuPjThrgvFiS1GG1EWvTYxY4BpSK26io960zmPPuNyO29qfgdzd9uGIUYk/5
Kypmk5h4JRbNJvd/ern8gA==
`protect END_PROTECTED
