`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xWdJ9LBOyqyq59HndH3LWVahwC2WK+Qre25UeJMHaRJbO4l1ayUJIVKZP4JqKKSW
f5Se5LMwtYxO3G+rLv+siCg24AOIBnQAB7oiDKP8t8226f/v/F8ycfOJjxZJvvn5
56JgWqdpKQRBm9kLuM4dQz9MaF/5IG2sKET7vUR5pMgNlvgIBXOyX/sD9Jo13qhD
sk2LHdy0+siNFC+DY0QT0wYyQf1IEabYQTw6grCgiAQYxNp1N0KIlycmby0HXho1
tv/SkqeKKjfx3alT4C1YQ/i+LmLHdRFsMFIEDT8q0dzMvW1fq0KiH4OZ/gri7TjU
kzemXAz7fs81/J1WWPsJzGAp2Mh6Qi8b6e5Ys88MmT+0irnfDgPW0SvNka0jAdoT
CuwXPjoWs49JbQNqEBIrJ7W4nf/ptBz+qa7LGYZG38j9YVVoo4svJWE7LCHrC58+
ggY+OFpg4IHuI6DMSgbUji3XaSIIlY8iQLK9q8hhKgx+v6iSAMIJa+rV44qxHBKJ
SVsSqoTDvmzVsVSJHSLHl6/I1CUbjRmsxg8Tw4E9vVskUu+k2zJ0HNA2L+owVoYL
hCYsG+0Z8YK6tGw8OiAFbt19e16QrDLwQW1hMpVNvUnMiGTfSgevuFsSQt6u9Lyt
E64kotnxKSUasKHeQx7hsQuIcEIKc0XVOj3/aZlF9CVMydgDA1FGEV8fgrj+RTHB
vG0s1ep7/Sns4vifkb1m0VcsvgXU8cqb7YK+WaYSs1Vu67a/vomsPp2atEtMNzn3
+my072he+wM4o13x9tmwYI+DCZqu/LcH0drAZniKRF7/DyPkZtvzHBVNacAHaNfm
dXQea6BGvFDlAd2CEHXAO44gly5YthjM+A7LPltotVzW51/Av+qW0SZv6OlMBsbK
4QMva/+VoxX/g9WqLgxKqlzJwOarBm7fbmiS9zMJ7J4djVmNnBnEZovnVyWtXoZH
kLEWpmV7LDXEpK16owlBmRhXN0LRbMkh6hUyJICT+q17H7t1PbVTjK1QJki23j3p
tIIrD5Cz98bscfimCx5W4mAPH5Rd3Mcv96j/LK0hhyx++Z5lwRSxz7RZoZwzodlG
dkT+pPoKru9IimV+vwitKe7pNgl4DwT88PxZBE48qTigcBHaZftdzU8ei7RsdUgP
940i3Q/U7RafiROOtWcAocT5VJePBxn9S6WZVym5DXD58hsB3mWGAsCduSTsOGLL
bIEcFwvSpyB78VzhIeLrj863TP+cAMBZQ61Dmqvcefx8TN9EPHDbQjhQrCP466wT
T7FKFVqyLWwkkbI8nhyL1DPhxrcr0+L1sLa3FKLosQtRwZNoEEcZ5YVHXx9EVLf3
pC8FD8Z1fsrNsx/AlzNSWQ==
`protect END_PROTECTED
