`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
64Sh0tQKE0+I3BiOSLDapcPR0eZIdbpNm4V66wWuLIH8nFaCcAgJOdCmwIrFCQYs
aNCjVGNQKDI4BS9HGvL8bGtnrwhFx9hrxSRYBfaKsbBO1kKE2y26m8SFqfpZLx8z
ZFGCBpyUaZM/RORs+fYRGJrkdc3AIn45lAAk9wqUcQwGk3OykLJXN+LOL/A3la3H
1uKx1q79SpcA8aRqeSTCr7XrNT6/apJh2OSekLrZB7tXCQu3X6AWCeQ4Bw349tkC
418XpWffZp5k2H6FUFU5NAQZFbuxj04qBwaqUexdEVLGTUhnaGC/41RupmQaKnpe
ADlLTIN0V2uiSezvZeSH3A==
`protect END_PROTECTED
