`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RlEu4OkZ8OjZY60s18Oz8hCajav4bF9TALnoFA5vqFA7cnCc+Q8MLu9z50Sfkg6R
p8+1zwCcDevyFNXzUjCUfO7DBbel23MfhVNN4e+6Ch1SPmFKNlQ7IfWqeEDSs52l
v9be4CCt0GOya1oQjC8mrL4n5cPxfTikbIqUd+YRxSZUhZjqhyiV0M2/i+mRAbtH
Ni3+AHz98EkyiuANTytTx3iyWWBu5e2b8aGpWyWrhIkFNHFX4PJyPGuR2REGfBOO
HUFL2yPi0Jk9RqkMJLfVLQQQ5kK/jAk42vcJBwOvmehEP8bREcRm2MNJHLkF7+MB
rWQlLiCqjt07CETYsaY4IaFPLUS7NazMh0hNmj9ElZkRNm9ECm31mX5IdezAX5JB
1dZ6smFKnIilET4oer1Pq6y8KWZJ+EQAFq1DMiZUJVc=
`protect END_PROTECTED
