`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
21SMwmyNh+AzPHAl1UePzhhh5IohRfFLdVwLIJS2sq2xappCrJ8zeODXrbOGbCA8
NhkAjVWGn26HEwwYdbwDRlVgskmfwNV1oKDAKSEj8+ktfXh8vzD2ezfmIwWL68vJ
1Af3PxEl+rlxUhYNo2YJG4TDGA4GGTqrdVM0tgAFdi0zJmXPmlBeTEcB+WuTzy6d
HUKYcMoZ2lSiABzyLuwaLTNzDV4ov6gyok6DqxAK+ZI8Bz/EMxY5Vb9HcSHd1eWY
ZrjHNQ/ADB3DUlRz+6UKKZVcGCfn9IWFCnMS0YiXF7ow1Ghk37vY4MQJwoMCWoSH
El5oIXbFDmsWw3Eu1cxyqk/lLdNkxmTVcvi5bgbnkhQ=
`protect END_PROTECTED
