`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zNg2SYtd6s2zoa9OKAzQQpMQw17dg2hffyWY/+7hHUITFG3w2ARVPGqzF8gZG5Jc
Cs9wAdMUJkvT0hJV6uUXiSgfkIqW0yDEUlh8bxzpn2RO0mMNFQSdkzuYQBF2ThmL
ckPub6nElWGHqicw5k9xyMynOGjJbCIuJuP50gotsBp/tuwQQbX1Xl4lxpP/5FfO
5uAoWgOIVP1VQPon/QDhIoLkx8/obvRYtFf7SWopXvVeK15CZjTha8aEwwSwZe2N
saJIlWUB36LNGI6ssZwshKvZ6kkFw1uR+49OaZcLwyI8hDJCLOtCsEw5oB2zve+c
/o83G/3+olymqXq86YssolhyEh82aHvX7vaZNBHzeQ7C0bSIIqv8fT7LVkOjTmAK
`protect END_PROTECTED
