`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NjtrpEgleS/8Dm85KfOKpMXzYW4jZrPcFw2e/SmJCHWlA6cq3XAn0vtfI+zxja+K
JlZjVGedfkCaF1ttWl5QvMApfseF4EyWjK06+VuJu+0vfPlxpyfbSOml9l3Gj0kj
1OovkvabErKEdU1vtUfC5ZQd8xWhNcZtZr98+fcMPJXu1H1NPbAOdIH0oIKRQ9rI
0rV6W0oruMehB45oTzaXosGOx2UW/8c/DxpkuFi+jwpl5P2gkS3b40Gr12nYdslK
bAE//M1XQGGnqIsFd3sSXQvGTAmhr5bu+CJtz6uUZzZuHqOwi5oUPu0gvNqq6ZLQ
ZBr+vXuz7rnOJzT8+4ZClQ==
`protect END_PROTECTED
