`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I83PxV5vgs8XO87X+bnj/PKlHIrZdhLOpcAtfXqIzv/UGt5Jc0QPpIoY8Pz1gavJ
pie301uREiQV2edRw6VL1DPU1o/6f5NXk/o3jX/PC8inPF+z6VHCUhh8+bqIna/Z
0jsenKGL9BliSRh1LO2ZQL3A+EbAuYDeAZcBgcv/LJD7+JlPZ/qkKSVcjdbYnOxQ
tMaqKTJHwqpnqcfRpRhHKmX8MXzzBHdXsQ+MGRkXI1A9n8zNJC1v6QehPbUg9Cuz
h/Qbf3IoQRGP3/S0YsTbvLUinJxKfcVJtB5Xwl5w+oOMhutBVc+XAURPnhou/R/9
2zhADLZdRIjauiaAtfsisXUZM+KZEvyXRQUvE5WFU0oSW5KkZosbhGBhWHcfLmLK
UpXBMUNk/36s7H/c5sEA6vdX0/f//+AMcGugxZ44UBoUZzKNiii6SwLCjx0ffwbO
`protect END_PROTECTED
