`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FwxZ9fe2hN+7+0nqaQP7RTHY4Rk5xT6gbBznfwjD1LN8jjcU9gEHuewJ7d/l39pn
LuW7iQlzsoEVVvA+iyXyvrkCCeftafdU7umIKiYX0+1Ru8kzIPV2L5jtaelmOymt
MDJ1pJa1rNOIoXmZAv8h3UZ6/rtcXNZ5DuSmG+a/mmXVmZ/zVaNDq7BfUBiMJqkw
4g7+ORTA9vQzLYD0JaaSUC55jfz6KDCqWlDxOJjMz9rFoS7FakoCa0KUz+fZ7ywl
ZbJ/p4tZEIQvDxkOXat/+EgQTbxI99rMaZyk8xMMhipNPOIxDktDo/B5p48NFpnw
j4SylNjtEUGkeJfDf+x92VBY70h5TU3dNo7VioK5vQLdNg0+aYLPUqaIvO75iEmr
CefkIfGu1r/NZhnf/2noZgoB7mTUg6WbHUcvMrXpUxQqVyI9Ll8Yz/MtgwClEC3T
pqzcaeUJDtTLvn7cDjE1uwRL2a9VBE1jGfyJBkLiXwAnGcpc3CrdklfLi6o8zmrU
I0NK8s/p+0U2PUsXelMSl33XkVMRK1juSQoHLefD3vq8j/kLiyl1mq4BXz36uPKJ
MWSBBDbemKZQuxkII6y+2I1RaucotEsBJLzJ+Bl3UcsYmmsjccxvIBNBDMkeeUl2
HvlhkNLJ1r7icPUOn/I11lVGQ2KKuA0FzE6ZIZwuz6M0wnm5/UBNenjRAbNnYtDN
0R/LlQleQn3AmdfIYYYPVt4733MeesMQ6Dj97p/yVvPdglPucEx+pCjht3WTcGqY
FscSIlwIEkc/yocS7NMx2L0DHjkuA3XGkHc2G2G4rVuSnqMFaE1+PRA8Oqfe3xDU
zON5eY8JgsKXwWsNxSjyhh2oFgHfsMnwAEuMSuRkyjXBgTcID0SDJrhrJbd7ttgV
P6GYG6HiH2QIKjbCt9niVAQpQxQBoitjY9fd9Rt8bueMZO367fZRbFXK07U3UmNc
vQMNz9KWOgFEGkO/sXdEhhwH9YmCeHDPwt3RPRqtbMsWdZbQgZxKP6YXvZy1ipEW
`protect END_PROTECTED
