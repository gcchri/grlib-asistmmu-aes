`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ggP6yhab7GydBY0a8qeQxoRYVgPqpQlJHmI9+uNtNlar93qv4n6NHQtjQCT2agrF
Acxk1+cT8Z31D7Z4BQOlZdcx9hH/hKvWzMQXSqMy9W3Ix0R0SDMC+WSh2/ULcMmW
8DhUg1yfhfKd4MmsjbCpcVM8LVnZsS//uBvSaeCkoDiYf099/KIeblLuMYtoPbM5
B/jC5Ay4IE9rL/cThAxW8fSfIv5kVdb46BjPckwbATKIT2KSBBn8EICB5LVGOaQl
+ySvd7cYQ2TIoOSAkCjfnmvRSww7rRzZ+xikHkRWhLcDuxA2my3fIqzqqj0rQYtC
Ar4nmM8M+Dcck/ucDxSdH8V4zrqupERySXdDDAD1oPOjYSpXdKVCnVa+o+r4Nr6g
OTgIfat9SkiVDhQJqFNIFHsdUcf84x48lAQwuRuOYM66o8AJSYEQjerRJ1d+4j6s
+lCDGQCQYH/v3+ChBbzdPtXgmDf+WOHZc7E15xgZbar6vdxi6/TIspQZqcRrzf6w
l7qwffhym6AtpJHJPXpdt5H3i/6Fr2+pq2VTEJh/aXsMZtKo4gmDAHV7UBj1dunz
`protect END_PROTECTED
