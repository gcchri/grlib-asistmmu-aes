`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B9JHT2lmPPzQ8XMLzUsBZCJYEre8c1OfRPxHMcu/r6qpym2ZGZAwTb4CLrwUnRXH
FYD6m4UcAaUT9ttt5eSEYw+XpdUBnMTH9ryZzK54JJnGQy9d9qHta41uYjAlmuXx
gED4rHb5qEokx4qWTB4bY3lOQeu7q+pYmfikFDC1ecIsw+7SdSNYeFEhbVCNYr5a
M0g/E30OMvPeD2JJOKclF5ieFn5onnqvwFPBrGDDzkKO4HlhCoS7waj8mGYUcw6b
TB7DiPkASPmfKnbddSuTPnM+G/+FcTwDwru+LHE41RSdTz20CLnQE1gWamoBaolJ
LIy2OOFoh81CUgzF8mokZRGg4370lBqsL5a01VpEJEmGHRA4rGkb0X7hi8GX3xW1
znj0hZw3xtTd2OG5i106dLpTpLiOOOrnRGbaUDf10+gQg3UdWl8NNHSut8RM9q6M
hvWkVsPi2Dpj6u6CM2XA+2n0NMutXWQgicovPEeSU9oWKc3vvD781RFVXnfDhF3A
Nxw4S5zXiO5AvLB9Uy9P9inTbGVzDyFoSHd01i+nELvc3ZMoJFKOoWbltaIvf4sh
ceRs/RhHrNyxbWciaehWneyxj9pa8WzF35+WE+tFgadSw3uMGntaaiixBYklUjaC
8FfYzNcvw/26+1U+qrz0Z8i8lTp88bs1Gh4LXRSd+IBiMZklPhc0+1mZNL599SKS
ZrQQb7H8Op8dIlVQX0qIh1M9Du6+a+MxuQhHnuvTz8RhmPKuio+k1LZWJsIDWKP7
DDjXWdJ6AAa3XF2h66OfWY3ZXY4ZcxRNHNrSRY4/As/FuCwMJilhuYHX+2Os1aXn
p33GymABhhlsSPeQcE7QNAGElkm/BKCYW3BvqqK1HIOd8JzEOfFfIvUD4/OUlW7U
3tJg0hGBRbSKXn7kAVeI6biGLkOOLCYRxzkNPCF8L/SWpEovKQvKvYbH+IxxJt3S
AMSZCe77eEZ5dU22cLy8JfMBaESKG2h4JuAvIPTGb7P87q7tdUUuTs2YX/8U31pn
VJfm6/e3Zf/H2PsQQ384ws3SsjA3Yan3T6UssxRJo5x50ex0vcugF+Q73+95J8y5
ehpGnsp9Tecrdv2cCppjZ6Z73xAMH09Qwqrkbg0MD4t9yMPthmzW7ZKuV7+zrHLD
aSiIrV9ZZ0eWq8ygYtmUX6N4NbVl/Y95SI5cXocMZS+sCMRcMN/6Fmeex4lKzn59
5eX9vKbl/wRV3srykK5WGTqJVgg0ipsIkQC4ql9Q2OHGX1Xx1wo6HMeEgDDL5lvL
KjCHuFjYTSG7L/HizykMA5fC8lqCpSEtoK4aGbytyPwploMZUYwzFNXe3lX/yhL3
YeeEz1yMjh0lI3m/YB+rEHfBM3sT/tOGqSg9KauTdyoLhF+4/qnEM1QjLenxr0na
xqNjR0UnDlFDAwteDC1xr47nbRD3AN+c3rKdveLHGz+6oF0qWBL3IA7LZT9xkGEE
Ei/fVrmPo6MechsVrNLrewDU+SaDQMNV0X2cSJNdYMdzuyH23ICeLHvj7gS/sg2I
oRUMg0SrDgsWgqFZa9XIXfo9lvTFLDMa6CX+7WAJu6ZqWA1OJvfjnf60qknbCjnT
B4INbwr53JLuYJqm3ibzPESDy+5uLo5XQe4P65Sltovc2HlglQ2htdd8aD1A9rQe
mbOQaf/6X1B6ZsqC2gx3a2xtj9u4KFy14q9d2N5ur7rouYddhtlz2rymFwMRBaeR
/Gd9sAh+3glRE1bHm9+mSaP8evDzkfdMJrEpJh1s+Gz/W6d6ef4sB8Yy2Uxr/ik2
D4ZtL1FQjYSDZb0c8N3CJWbPvbOT4bGGljG5o5mQqqzRYqzqvr97iq7odKpj7d6R
babkIynIf5bOYgMXzNP74tLg8YmG7aIe/zVtPCa6oJ07TaEOrBGv5eObnNkh8c6J
S9qR9ZhWu8cs3D2YI2sYYEyWAG/MnK1nEu4avBFvPzQOPS+YtWF4t2T06Maj1Xag
HHM+QRMbwYbvRkuigY+XZ8ArfYjtvF2Ou5q0p8JbRao2+VlDV7Bwz/97ZAVS/Wyw
Cjxjife3WoExbERx767Kmr7n2zkPkeH3t8qNxJlf7+7TbHv54cCy5BuCR8S6r2RN
mh7VQdHfioTUyOat3Y+u6fx/0pb/aI7wQEHLBLHiZFPdMCyr1w0Z/KRC5ufPDduK
FKPlflNYCLpYrfWAcrM2EbOTs633l0Rluwn8qVLg0AibVJXbE0aCfNmSqRY6r7vR
IWzJWqClC6trsZwHHyM//uQe3inHtr8FiK+kBEaLrABGUmm6qtXnEUPNUC+W2XNt
ZRxqVB1Xwj/IPbYYJ0wT1uSj+8Yxie2NBsYuqr3/OEd+MRUI0H8GVMMkl0zya7XN
RShS8y2JwpxzgCy1IKqqR4kVayryoe9Ueg3sSiISgGC7REqpbr5Ew3LlBkHrniRd
Alp4fqdmKUFqsQGOPQafNM/8UrQ6ePw/qiHJRHmsVuf48C4P1v265aLnR0JvU8K5
estzBGtGCMrTcXLpipAQcakP8/1TxlbmfonfSMl5vkEsfdfFPLfLzel2UUIIl1b7
GBjfo9A1+weR8bs0grvAXeEyJk9ImB1cVpSW+wLmh9I6haDtQhZ/9sFev+d6A0g4
y5070TsOt3UlVGa/uGPmojzJT/ApS+bNMlB5N2JbyeQqQmzwx1T5rdRGmongqlyd
ZTiJ3FtejQQEMCiSi+Jkykfz8bJ7RDBwG22bfvxmrB6Uvt8o/KEhceK+lu8mGanF
eOTZLkOZt37zp+114dn+ihvjwQP/z24oVT4MhQd0pgwjYUais3sy+42w0sDrE2Ns
xt3uK8cZgmG/svtcbQgel/V+Id5pVEQRtIknQmxzhC6uXt2XLlDlFUb5zx2pvsFR
MYs5KIiNM4Bj5e3Xi11smUhUosm3sIpnoXkQJVskflIuYR17yzeutveE93ZGP1xF
HWvyI1SIsd7BnL3IwftWX/8NfVhg4FQ1XITIH5vzNgzFd6V6t/nAqOxAco4PMm0W
EoR757DlJVpL/2pLL4T2EVf9TvAkrZ1Jtm84EiyMkzRbVMlLZ2E+cjPCIOCY6fna
TMI9GYIVysVUFRXesRDWMcZbDhX+TBThX4c7sgN3KwJ0EwfhM9msPhjSDUPkoio8
tp9tR4xH+PY7WKaYj6yKKZj5O9UZuveKFPcqyXqqcV8wXNurpb1L/MAKlIb4RRnf
M89PGdrXETI6BCYjwBCDXs5oMHcdm/En2f4a8hdQuhFYYcufZDKYbLw4OJf0nWQY
xRuNPl81uTVztDT7vLXT06vQZ+R32FeMbYcaVIuwOS+F2YwNXObspbrc/UohHQYU
r2GWuPfOLsQ3095rYXArMgcb18pUmCDLxNHt/CQ5PCdgUJbI9y3e7xhfKwWzH0e4
O0VxUa1fWGL4iKsBqjCEO7B+Xa2y0jVz6EjPyPzWJ4lmHQGLo1YyKDmnW4zxuYN0
LYvUofy0ewftVJUgFK3OTTD0xR9aWMJcSChgJ68gI6HOlWckqQItcmunBBaiaLZg
bbBqgyYTa0lWgkri4BVNppJOxoc5Fd1di9Qc39Y09Ny0CHT08kIeCn6ypgkEEbcQ
Xq/JfItMPvi703LCXCY6I3QdhfyqTux6Sz+PHRIwF78IMkAgTXffedcZZ4xEepX3
6Uz3XxIVD26v6XQNkO9+Q6/Wci7fih+WRowKawL+2aMbriB27ZLWtVU27N11AgTy
qUvUaMtvy8T7h3S9/3luTiYiPMpX+iF0paYf4ghH2SWAMcywvntWyouWC32fvemC
kbsv6vuR6ymiuSIigNwLHvwXXBFwWt7TmHTYIn7K0Prk4CmjP0wE8TVFoJyPfkXU
sHxMu87JV9HgsBFv0rgkWVeswPWEp/M2Tnhy4TBZ0S2itn7/FWas8XltkU/VtG2G
/rmaAb1Zcz9GTpN0HGN5mcg4XEGkHxgGJXkecostx3Pnkbxz3q2EkRKkJkAx0/D8
KoikHzdAYQiN8nkNs/t90FJNrUSTX2B6NbuCVpJqMfbf41sX4Lmrbsw2iM+CYm3S
Sm4bRPfzYFoAoqj0GrNOMhaW67JVTb0tkp6dwOE87Pk2AF6PD+oU5VcBt19hdVoT
cygdSFpe+6qrGlSNxFjpxCWl9CZal50ACDGxjwlo/cbSmvIXxDvoh96cDGOj4F8U
iP8MwLxGOvnfCSL8SkawzPgP4xbgcMhb9Q3HWFtUXs2ZYdjtIarySUK5DgY/ICYp
NQhuZeWNfknoIHmbSuxutjdAgCiNCgJ7feP+Zm6M9gh0Fxl4FesqMmbYQX8PIgo2
GbXXKD3IuxxiNB5y/Zmbat/m1LHhfRa8ipq/07a7/fPosgGBOuiUqpMno4zdyAFQ
i+d+O5E5+i2Vx4fHHAIByXb44KXGFS46b1yJ5XWG6iu03yyaTyQQ2vgapS3WviHy
CMFk/uBnSmVhEwDC9s2ha3IJJEMfP6yzQyg5JtDLNrCm7FRmRmGpGJAHncXUcrz+
9MaRWeMZg0I4PdXm36GRfdBfCKJ4weqpQU7Atkn10jCme5uUS3V+jgxfz1QURghk
wVNIhcmTPuMopJSelHoq67N5ktOPwj/8rLlbJWDL4Z+jFIjHPtabBqjZImr+xtsB
thUA/9V1sZ8R/Te8B0mtVUyMZS6mbJMmgXLiT4C95rd8kYBLQ5fXdZHoj0CtT0Ga
TKcjMXWIWjZDhIgLXzTqSV9O733OF9J5j++8Gb5n0PLyFKUy/TEwgffbRW3SAp2h
cMgBeWOkldwO6s4HQVIo7s/Il0NHbFbziEothnsTCDeUsnJkVyNUH3BhV2T2MqCT
5qLr579oGCxrynsg4qZ+SzFguTO4V6g2a0n6qY1lXzpv53Jf11lwxQeL7HL/0krY
Nlu58tgd6qh6YkYXKptknpYFsPwtu4h5sh3FnHvPb4FVpf7eevPMp7I96mQW6K4/
9cVR+U8YbT/xrtSuebC8auAL037Gnzd8hqsX1yY1guvDTmMH9hlf0iWpglHZq597
QpcnZjgjx1GcAa+vKfZHz61TPFe4HXGg8bgcCtuOmJs4+GFrVW5+LST687zbl5Kb
8u/pOnUnraGJqKIsncqFqdoWFSGSLxRNf1y3FcgniYI958zJOMgQ5QgTZOPBNFmB
8ynxRSKAbTvQOQujMLUhAxMHPm0Vv3avtUwdQX3gRAY5I6oZH7KPo73mE4Yepef3
FWmjP74Zg5REszDLdjodekVN5ba4G/UvbBSSxbK+m7pLsyMuqUAcZZoN5w7G4F2J
aoTXuxHR5zoQD6Bm6hifqn0P13+QYxQB1J6IaTOIgwwzlD526qmOVfU4mte/xJnT
Ikh5jWUg2ISay5elkYUsmXFNgjZiSrP3ay0EtCj2YKfZdxyQtrOSuTz43fOAKSIv
6XD/Mz28JGEFPYYQyHQOyP4rzaFCj/DMgagpGOM6MDH7lv7GmBrES8znZ88cSrpq
seLEHqqwEtUlXYyfvHWXlrmNmAqsbmVrYUZdjCdGkFJQx1x0ViJ3BE0gn3SNtYD4
Qj+RAZrPUdNy02QvSokJVt0XbEFFrQT5p1RnoDz8+3Bv/tjdEX09u8c2j9/UN6di
uKEk2E446lcsEGndVGZJkO+026vNYPUMI2TTvJDCipuFmUBWncI/xU3upwwXPoXb
WVcCKMcCr66X4TDQnktZfL5zAB1wu8hyNwBSXgMnKFXB763IeU3kyRRfoOk5JbHt
YC1cBOR2jRaLE4BDVmVDKkRb+oJBOiAGf2hP3Vl7EcoLCndSpRoEy8QWY6iTK3Qk
zuwEK+stsikokf15yo43M36PkHZibVogfb9gxTvGEwpMkcLl3bAjGIIGn/4KIxeH
auXv1re/uFAvA86dn7EMqr4DCum1zenJk/djmkJjI/jDaJ5D9v6Ap4PlPvSlEN3s
Gv/I0t2F10p9goTet+iY4mmpyRhGKD2g+0q+F0URYs0BNTlxWaowIzJuO5Ef8A06
3NtUuaK1Mh3Hu5Oqulg5ff0OUJ1xek/YjzdaxGP2PQALIUbgpxs+cSgowVIgLoCL
cFjUlAV2SA6B6MY7E+ABPOZ+76Swo2+Nzha0uE8DCbGpxqK1bH8iVxhS2KamUQHj
j3a8ezGkH7GxQbGJ3MCELG0Hcptl+wf+EjKtngzH4bwbfpD9Mb0LYPezJ8Qcu0vW
dZy9hsU4nhgGeQC0Og+GWIKIu0b1F/sfCqdMP6lxS0wLEmh4BP9YoaHauoQbJwi+
03mtwRXl3J94udeBYQg3o7l/dGpnkS86TwhTTfOUy3mjJvoC05jP3/IRhuT6Eh9q
EHXNHgkw3oHdw/HTSR6qdwExhi26G375GLvAiULDxZux6J7XfU0lq1Y2HBbcBX79
k6cl9Czv3gIJrSKTZ/c994ZQ9Ti3dwSuLUSumuobuIA9s+Oeh7Q/eZ2wXKdYZsii
1sbleU1m4w8YGhHByvSE6Er+TToKFWCe+2ODTgpzJqh2iR+mcIcnGA4vBxpdbm1e
mJwZDlYXlPstvj0xq46UXMOGoPpQFqQmCJ0ai0i7auvL1mUWI16RulWMBABdnFXS
k0x1/IlfNzCwmTcKEg9DY0Taqe6QTV9+O2LKAE+z0DF554WGznRIUyh7Xmmii91b
UojMda/58R8FPNVYWVN2L2TgO7JQ/dB0N+GweVWPg1w1p2Mlxq5OoAZE4PxgOJBv
M0UBhJQlUTjTP9IHFUYPXV0G1X9dKok7rW9vY48ulhHHlvsCuQyihzFIZ3MBLnls
11Lp9MNIyjBLGHYrqxB4mdDmUhUOvgA7XuvmzAJ9cQAOp0gRM2N8A3OD6Qhgv5r/
0BvP5d9RnhIbee6LiGRnpDANTtf56j6M+GSdsIMCjMSvoukp8DflooN4sqjzOSEQ
ZUZ0289h6BY2xKTX5O5BiEDCWHb3abPVQKNUw7feDoAMD3CMZS/7rLcOMZXvS20S
Zls3qD0dHMD1mZWdd0hHnIJjEzRy9GDb+Yny+Ct9+KLrZnG9v9ueL5HMZECGUBdd
K0WyN0xfpWhBYRDme/+6P6n0n8jrgopNBmMNf2p/trARbd+Hmh1UXeedY9sdCceh
riLrfEFvEnfQJJ2abti6swDj6nJxKMgyTwp3/pnwzxMdPIA5RIcRB8RCxpfnqlSo
Q0BIAjI5do+jaAvmyQvY7PicT2Zn5/t8uxR4NJwHIJt3RntHRIdxFpejN9MXmE44
rp4tSRzCEc2GH5tGnY0+TEuv5hBm9NUPytRrH6WJdTPu4L36PJ1cR2bDcL9X19JN
c60i7uKN66yiVXQVlZQsqIwPxnwnMHDOUAw3zy750b1gy811tyeofqwuTqwvAnHV
E8Dvyg/u1og7fANkUhTfwT3escyLIivl1lUYmfOhBN28HPva3vHSPOnKTQhZ3s6u
+HWrrIlV22VKTy5XPkkOuEJAbZKvA5F7HATQUPtubKWKQcWMksGwhLp6gBkpG3R3
yS9gn5EIswkUr8j86HbCYV9FJwJkAx3kzZu3g4FDynALizxyIBDQubQmuvJDajws
G6d4tgTbC9Nij7S2pq9BJeG960mE9COvmkiMN1t/V9HnLORVgBPmLmhk4Ujne3JK
9bOEcxYYthoJU5mGDRmrpp03f8+QFAz0Y2mnZeIY4TwFPAHs1adp1+ZMzx/CijgZ
xgwPem+4bV/BkvzTXf9ZftiQrAnB2KFcwsMMdy70RnvxjbbvfNrLiQAPsZfIRKdt
Od2Rfk2dapgyQM/sEZ2fA2Uf2yaiaqd1Vw+OUtjg7VJp7E+sKn+KCj8aGnlSWcAl
fqlF0mD9WSlH56twCV1TYRmZ6ugTAsBn/edpxKC3gtVI2M+j4Hz23FZ7jgeILcis
OHGSQtOirqmlS43rb8LV8eQ41Xy6JXVGLthJ5K/Gk/hqzgmGq9lpYh39AHJJlAh/
98jpDyFZgH1bns1tJmGm6YdGJpeAuMKDtPG+XHXGQ9cfxbKfgfj+oj7JV3bgwOJH
j4Iopb3WDtADpRj1PwoTSi9HUOE/rY1tsOcCay2q9LnJdKj/Qw4S4uLoJvAo/aGH
cBiZ8KlO5fvonQaBROmOVGLVPz6f+qnVwnLtpk2q38cNju+xE7NCWlfVMarxlsrh
tfNq5ZHCwbFKxTdh0eGobHXdpSxGWzDKw5BVU7vGel7o5RHTMVP68DsPULGRT1K0
uw/7LXUJ+7Uno7WOMTNh6dJc2hah20CO8VQvUN8KmT39r8E9Yln5liwfUUNZm6ut
QDtVFwUmxQkMluEgexGrcg56dzLdiwHplFzvFRVSCrCDKMtHALdQvp3Vc9w+ggR8
sYxqWW6iaPHdHQnMBx7gnui2Isx0n23BquomwojCvYDtkfL7Oy47KJbdqClmtkXq
qH7xRdwBBbYujBPucUGF5DRhiDYU1tG6bSL1eO6O8FjVmfraOYaIKZsjPM1N2gIs
KOWD2Diz7UWk0xddhoy6DqMfQmCBkGSlhMZNSJ6V0jdvJWQRV3an4pQnlAakfNxF
yd3ozzVoCPJwb5cuM551X11Uyl8ZOCThW9voWuTBEWjBqyaH4WWYPaiULtyw0as5
J2T7604aAVw1PCaYAcc7t9ovYGINQDHxABdINC1WKYDkAuls3DkN1oAX7ur6+5kb
CI517AByFnu0eyZV4swIH6eG7Qw1TJuadMB0UAGePaGNqFckcQgtihcIx49Jbt5s
TTau7RJxN04knPVHTfNJRiyOOxb9aqPMS8fVV1IOUkt8Ya6RwvaeZfml570NGa7t
2M/DjOLRWQVVB8Ut6SVzLRo/fqqibbxX9c/fkBvn9++IC5TcExvXD9VprS52fIhZ
Ra9qbuOLVtOJ8/zDyHhvL42ekMKKPpD81TiKF2IMtzgNuhQH8236r3nItaOZKcg4
YyJcS+SRGytE4Xsov4bH+n6VwKBs5Akjkm2KwtLdAwmklVgJvhDkbWJcMMfelsuQ
Y51fUUDfXKbPTv7dP6uUQhhCKQsy70i5yk0I+2XvPSCUdCF2yWZTrKp/UKmjRx57
aYMxC0jv6U9Yyb3zaFvRO4PhPevegaT3jmUu88PWZLZ0FquE+ZNVd5X7DCuVeiWl
Cq2kFHHJen466jsjtN9a18sGVIQDWBVhbWyCCXmw8G50fMgCR9KrEUT5pu2U/+F4
Ak4FUa1rVRlZLHNuw7oXrFmHFlU06yFgJ+eMrcK86j5CA24M9BaGjwPnNieZxB6A
fSgzVLif6YWGQ+FQhKdeyWUYSfZtim2eVgLNahP3BXQFA1t8n//3rWbA71KZd11L
J/rUVXwz1nWDtkwtm7HVWFVXFCDmkCXLuUtXtSbavWatKrpisLApzQRlFeD6YWyQ
3ZX1ZM9h8Jo+fN+fRd9YjTt8++QRUhKrVDubCNjifX+jpu5v4daua1EYPg/4V0BF
oj8twt6J7X42p7B0VoFRnIJq1YsRnqjHFSTNxMoPDy1+awrY18qYsqweyEFbAoGk
vvLvvt4rYhy+P2PJ5kSTzrzB+SnXGXAt+WE4ojKnynG16kwn75RC9B3CtLg7af0b
x+W60pKq2UUYaRaB1qQfXodD+HpzCzVpyR6xLGGsuev9KYsO41UNugaUIYSSjFA8
Ol4y2KfGSkCjHdQPgxg/OKKAMMpzf5cZtB0DElymYAXL6pZAtdguTEJeC9TzUl/E
nMRiYMHWgOsIQh89982d5v8LUYhxS4Xi7rHUoRnFDcLAK4zM4x+ltNrwX7WYyAdG
cP3C5LyuEqE2T4X6e2Koal1DhTAjJL+Xx7EjfEFuVJJbwm4FMKxf5818muW6u9uu
8t5yUgz21gK2yqwpaRD+18iPlkTdL0y2/bDfRWdve09aUmnT1iyETw9upkuJjGwI
563OqQUHIYpQX8WWkc8KSv3pH1GTuNdYAUPpseotA0KOqLh8l6vEFF8abPZQ0gMB
9mcjI6Ygu3DrC6KMA6QZm5L7Pe+gHvh16dofdkHiaDI/XGU9SWg7lHzhAew2+czq
MB0VfqmBQ4/VSW0VXhnnAsmeMGnBzawV9ppKbC3g6cFv9YCLHplMs9FdM0aCTjs7
oDor1lrn6qqcCMabRtul5iTqPSn5Jr6jTRP4nPYt9PJVdMGbJbvQTDGSGT+P7Fx0
iU/iPqiqYG8wGLA1a+bT2CyxdErR7YSdY+ZVmrM4tfvxmfAtgAdEm2pdnDkkl0iM
TjyZBvOnrbq6Hv591bARNHzqYXbafcuUx5pAUiGW7AOuTkxxQx+CDI/4ta9GsDZm
B0SmcjmKZx2Nv/GFAqI0PER0MoLwQFe4PqjgptJ9viGCULLIOvRAI3N3PV9FEPcR
3xTdH0iWU4bjeMFiZrQGl3e2BgBYBkk51N4c7S7QQeDmpYuCGrLLzVifuthzOs7b
KX3KPdpeSkESrmR/JB+wDYs3od9XhJFyqqXtlgjvcpP1ZsssWcKdBBWxHGPILn43
lE0Opdskj3caEpjDewbOtQ01nN1tXDQLUoy+S5+yIpbMK1PVA1VJmzsqCwqt+Wda
zKIBsQWLwHZzkLbM1RjwL8GiKArG/FHyvXUXgmXf2S1gKCNqxBCqtWdgeBP14Skk
nxeDpWrfQ9UQLnSYSCVB5b6GoSUAP96VHM1lcr7r+6puq+QVmfUzBOrD95XPfI5K
YeWhLw0VJsthGS8Rj5kGytxsIU8RjKt9HGlfxbynZnP0Oq1OnfbVUYoB5e7YbUXn
Fu/LSXlzzh1HaxRF5mUDP8fCZYQ9skm+FRWukArfMLDTQbVCpo8fQFEmWeycxXCH
iWFBs1PlDFzDJErGmjkAumnxoZDxMpCzGJeeXRL3z35gyuKVc4rrIGyCBlgMBF6w
ganjcvNB3NpErH+XstS/IX3ilKEpyI7lBFbvypfjxscDrspHkNyrS+WYPNaHSiyX
xNSM1fukwYsbtUBFAvGktRV/p8JlYSEleWpmv9j+4ySsIqUYZQzK9CMs4pYKqe9V
+F1kdk6qs2r8gRcqvmN3ZJOs3FbXtz1wuw+eetMoKhooG3FZijz2f3SihruueYn3
ZX1i2BpsAEhXtEIDhmo4eOwcmSYCnJ2uk+aO1yBB2xYarsT3Odi9IX36UqFB8MjG
/KS4lJLGEtWA1p8+YU002nQRWu8EnGfteNv+aAm6ikQ3VkuB6I5iU9obU1Jy47dE
2P9Dk7Ye96HLFpF9hbCLURT7Z/3jcx/gI3+b6kmp9Wj6jHWaDQkdNm+UQ8gqpfdK
Ila21W5YvIs6YyafB3qwCt9AFa7f0wtKiWiQDypXw2cnk/p0U1NnSw5ngM7YG1pt
fTKDvrQfkG4Fnzkq/6V9K60kUT5Uvi0inuEdKHI6kHS95w81z8KD0Vghei+vgsBz
ZoGq5P4ag6jmf8K9QkJeCq4yWSABPnjVgfovwKIxkTPzFtf5z6dYv9ddL/3ZT+9L
BPHxdaFiK+uu3mcKL6macJJSTIFnB4X9KE0XTb1Juzz1fkV3j4FPIHhfCVawfpdv
0b4LDMIoKx3MV5PRT6JbF+6H7L/bzKtBVAvgwf2cQVyfH7+d2N9inaPbbE4pHMpw
4gHuArsFWyAdCk/4jnKb87V3QyYiQnXlbIf6wUy55URQaN14nM9GuejGNGetghgq
1xWDuMzgZNR5LZl+G3NH3mxPTd9zpoC/wpSfKT6OkUu4284Ie2TgSYJ5Qe/tlIjo
mJ4A1bW+KWhfsOEiEwidZUBCiyPyKZSnCKkTpGTho7I40EwHkPNkpcYILxRP10WN
cBt1Pql3c/6WfYC9OdKtBS6HmK1H5VqJU79P1Yj+P+F4lpGAiEN2C+eHcre8a5mt
YXy5Okol5LWCBN1u2GqrTtbQF0Lq/jkzvzFv+nrcNUnYamYOUJkOW2XjTaxGW2xO
WMchpon6KVNvXzc4pL+iyJm+/jLUONsvbfLGcDcd1GLqNomJEO1zdwRXwSAP54ww
lcFTstD2zqvEysh1sGdvMa3akMp3hiLQBSb90OifuZ6LiLtb5nOAszFnhKpyp/yh
sYQbAcGv7VdSzRM9i3uGJABda9Vi/eYxieXnzlVaDAjILK+iqjVXsmqV7oG1Gy1V
7t8DbI91eYXByGnddGB4F8huLr59A3zMqDgVvASlzS23fz9hGDlanjnzTXPHSr+D
DNRHFDsKodCYy9uedbTEMZP0TcUQSIKR6fcQMJ45UgZI4bGFiM0dZL/YzzTxjbsm
NqDsd3PEEQZGjpRSL69xvZ8YOgiS4EHhIU+vFvmOQWZgWSNn7/pbBmzRsfhSOjlM
CrHWsTYClP5O9pbyqDuOeYOmJFDSiq5tFx9YGmCJxAMcXngBzAc9u8whlKYYbHkp
guUJX96S6m6QZrTqmy6MeDjHohbP35J6DbOA2nHuqDRwk3l+O0PnzWsd13iP+9Y2
LxWl7fUjBwqXt1tXh79w/k+VR88IFQNjBPvopKOujm9JfdK9ljjvogV1gLoxSyeL
NNfoNRo76GdjkxZgOcodXTZAdJZDgI1wE0p997T7R3XVbcicjy09JqJOvXAiKaFs
99VkKMz9MQf7R6bPBAqEBNt10SZQuVHbedJH6Qao87fd6K8g28EKVisEccONNQO7
G8oJqC/p7DF2KTbmoiW9KWLA8k6WbGY8AeZPyM89FcITXc1yhU7VEDt9baqGrJNV
8t05invSw0BvjUJPwayCIt8JBBQCg15FbKoa2EzkRKp3bofxX+algjFTIAQ3qGxm
XDLWutNvPRvXvgi0BF4CjJr2/FB9CM/epJTp/zhC1CwikTOHVHGMkWCfn624a9vM
7GyQ7wuoQaqs+e7FF6gMWo8XTyVKHwXSaa/ct3DLbqpqncsTNIMGcPSi76OndrUo
B15CittfiNCDTKEgI7wiDJY1U6GuO8Q4NF2gMLe79DQ53Umf0f4/FPBP7tJA95Ny
1nF6GqNJeODwT1YnIJIOFkavLdw4ubyon/ipP/aq07hN/A+Tumt1pllU9pS3ZvH3
qZu3l1dfsIWR6xMYBZIpLzt81/eTAlQUi8VZlwSvXd13Ev9656zKCSbYwiH4dbKh
sYDuZPif2XnIeE62SyasW4ji4XuZHaDuKFSavB0LxWty0Pr6LK/WJLBPdPzZqsfO
kzgGy/Wne0ZJVT9rfu6Pnn8Failp4OtE3wntb67d3GiT+jPBj1Z/O9kR/dGa6lfD
UPsomf3g3k/0dt8SV76xWzMgHTQ7hb6df8iogoJXrnQGOxr4epML5SiRHeDdSzaS
n7mxRRGawleUVokmI2gowMGVLAsOANIqC/HBrn+wEQvNM2WCZNTWLj8jgN63+5bl
289NMQObJrQlJURGzqutM8Mw+xSAWKy6YHiPqq2DW8T9Ba2BTNTyteC25nhTJPBF
q1qturHSdxbyQd1SNSwAq2UI9OgSs8BZ/yYUYzIqBvw68oSQpzaW2NrXCa73MQnD
4kDuhfpeqMPK5oneuQ5T/XyT8gkzaSEOjQB5qxKrH342Hk6WgoOBc4WBJfOF9GPX
Phs2N9sSIwAzmlyKYBRtF3+KaX8rPlwQTJMZL8F6dikDB49vfHcMx6qgxBt6gCe3
OWGkIHFQ5MP0hXtFEIRfB0SG3pnO6HwPh2LwI81NrYmGIEIzXh0gFBNesEOMHzt+
82LzRsczuxncV2L746PmnF7Z+T6B9G2bHAOsc6+dJcCZmfeAiU1Szh/a+g7iFG/9
w5RgZLOPvXewbml2j3b5BAY4Q92u3ysVV5O36+uZcCJ4ZoU3erGjOiRoDs2Qja7f
86GrH3qColvxExVUeNuvnDZUJAlpAhJxjeiXXc8xb1m3GmC9DNQSnKqimpc5/PUG
p2UFS/lOAyWxB7NUFMZofmMLlGs8Rtr1E59Yg1xv3T4hZW+aSgbbIWYZ9Lq9lhiX
WeCjujo67or4MG7hBl+6+vF3rxYQSipGeid4bWS3m7r8qX44FrkPiRpNYMeYeI6T
WAzC+SjfOi3wVOd3K305aQDpCi1d47vFxRJ+JRNEcv36Q1rtw8ZCwn4CezB0UUBE
T6mYd6xr2XTRnAt26/8d3raJ+q5vOHjTTp8AulRwZnnNbkokvDFc+e5PjA+GPapS
kUFJ3oBRwU1LhnUFHxhLRKXUhj3VYJd+C2tfH+U0gMt9je7HPfjS4XpNvpSepXmR
CgQLXcRKkd83vVn8lWOALBwYVsjbfERBl0lxEtzvXEhsxRmMHiFZXa7wFmWa8Tis
tcVRVtHPesCRaxb8v/iO/ocZtSHgE1JQII5i8bNRiHpjUbg9GaGiPmUcd+r/SO1r
BqT8JMpK+llz+MEandLXgBUSvCM/CVnuQuNuTdAFn+UlSlfV74UBPnHhZPTlaQlm
McDsAxV3D1WyBhfPb4HED3EPaam63rW4nmstsN+jojuJ1CjvpBzjOtHSs4CQZGMq
75hQDhkAj/Sbe7GD5MS5F5qtzUOUlwlUFNt9ayLFbpi8aetX0cbrXDj0i8B02Qr4
hRRp+83GpE1H/M3vpK/ugv/HIoREh9p9Li+sR1rulhhdyyzryzCkrTRhXpT3yMby
jWKuNr49r/P0dY2VHmXA/jjWmJWkZfezT5BD7Ss1MR0tC+7+oVnZLmH9vu0RKSUc
7gmrJuu9nchBBCOjhJkF31ldH+3xaR4/mJAuZEFetFqCJSikKd4YUaD8XVkkKau1
HAShts3RStt2vei5V+eUpGPSLUh3OnosQUfN/6jcJTB5s4Fae9TaZzPvClwAWD0M
xJHbvot53xbhjmHT/Pwlzi/YGD7/7GtsfvZzz3vZyyBwSnUvEGR4vQ8Vkrgu+toB
`protect END_PROTECTED
