`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f59FZGInfzETJUjqAmrZD7KMgMafg+fE4aVEhGZiftdL1FppDB1W7irBmH2ZBqy2
Io1YNSMBigTNpRR4+BXfkesv065sOXyVI1zf2NgjgBNEdH/wNfQpfLG4o1LWHqxf
dQiV9u2ad0v4nJALhAzs/c2e1miMnNMOtMki2YdbUl/MG/1ua4zPFKu5hA8n0nEO
e2KUTktjf1uDIu4iLS2BW8Lmu62cEsWIkU7RupwLAYkrTNXs5TYmYDlT3sj2l1mf
EdHXVXmHT1zkhxPADQx2ln2OUiubeC1byerfc2BS4lVehPenaSxqKH4y9sR6Up0c
cw+wCylZP6g81mTBLGxArT/HidstPhC7OvC3tugZKB4yVjaISXeZJICEVjFICuyo
DPD2zWZtjam/uE6TTSieRu1mGkjOon6VzffuxEb0FDvT3DJtmJmIe33FdyxGQbM2
iWI60OXcM8tpQgC8iwsIL/mxQk9Bs2Yg5EL6dY2kyJvng8jsZ0srb+PyjSbBpy7T
07cHB3zQJlJ+rxzXfzExixYtQBQp4veH5dmUR6MQjF9rr8mqeGAGBQRTxVALH/DX
/sz/ftEsrAZbta/qFVODczLDD3qLpHXQefCE8VX8h6QcnsElvoQpIugTAo+BAn35
DEkgyej6o1MDVpC+Pl0M2a500HEhlBZho37ABo6FQnD8Ve8U4F/wLkQWFPRDZjZj
LCwaXNtKsPzIZRdPIKsmYWCe1ZMGlNZEzF2Hf2gNCNw6ZvPV2CV5afq/WgRIFnvK
Nap4Ew2/Fwtt+Jl2WfDK9+OrTUiuLvpLXxrgYe0vllyBwBmpHiaumR2/mLb/5Mx+
cEQ8AMTkDyFyfGdh2GEr6Q==
`protect END_PROTECTED
