`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NoqoYWY3Su9JDWJ2IZBMITdfJZIjexqFsAeJBMcZIn7VnrZJYtbB2kytCqZ7vh9u
3Yr+NncmRhrXr7IWajs6ab1pe98rFD5zs1oP7qH+TpdscjE6o8wEETsxnENc5kXd
e270mtVwW+78mkSuCGbytbay0SSMIdjZQUwPDG/pDn6H8LKJN29p8AQlQmVh55Ft
Yo7lKJChRDI8ccdOQ6XFiQkcqp/XxcJCdP1/j+ZmcQ2t/LTz/WUaK1N0heP8/zOm
rwT77opeYUpqIbEOTJ8wkpmYOpo37Wcvr3LmKFmUwBUJxh2fr+xvceTYlxPd0s/Z
iQQweuALFdbvqzKx8QhBfPSwGu2Yu6ZKU2d3sYta3vNg3IjvuwS4U5aHNnGYVX54
qi9Z5iBKL1UVnNMxCvf2d/KU5/iQa8u6bHmtM8FqaKbffV9aG5EtgJ9isbowpfkX
khbbAjdztSwygHAVNXoRXJKtkuvzAQ9JWyEPWY3sejwTBsRBZUj2avZ4s625JGVu
JF1TL62CqY6/9tzL5RDguggyDBChvRPRpxTJ+2XIlvMYSqXVv0z3a40TCzHT42Oa
45MjecJthVawAIidzGIn5t8nypA9WBy8jUKGxe8V4DQRGc3WCY96HSCHV7K/Mwbz
HRfMP6Klx26ssnbWOtyiJd1EAXWuv2vpDApCzDHtRtc=
`protect END_PROTECTED
