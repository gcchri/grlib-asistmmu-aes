`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7CJWHgL4KMhvsk4Ya8iIEyKicjZhVP2Z81WdK1Ce5J0OQxT9xUgbjjjxkjBBVXyK
DOOYLYkFW5KFhDX5xVJgerCDB+v/7IzROOKDcjJ97virYNLJlW/yic3cBRWlTPIK
BZSdu60nrsQRPCJr57PeOvRb8h0rNdKV8ytLxj7XDtrs2mDkPRmcvG0LGIJqT/64
bcrmJmn1WKvSd3/tYshUfZ4orpx5mRkQLOX3hYLga7GtXsLp7SFWeI9d/SFu+U3k
IlV5hgqGuxprhoCdnL1FeWAWNRktOk2GxR+uuJXrLO5Egk8q0UNWWRsGVHBYd/sD
aljmldUMUQnWPrV4+VNdVlDRiBg1UGVyXPPAipxIk36/29GgOhV1Q53QcN1PFZsx
ZDMImxmTmCQKYIazpAKDuFKaj1oquEgvvo69ewylgfo=
`protect END_PROTECTED
