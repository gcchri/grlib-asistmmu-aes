`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FHIQy7GSOORFwKgiSFUnWlFEbzUoJ/01CaAyjrS8QhjzDDwGBtcwp4izNjDtyOR2
U9DDHe9DjLIRwPmzDsAHYBpvoxKx9qrQCkRAloBOPQXZQw0lPT9joBh0S0jMdNHv
A+MdazjD88V4gyCILJjCOiFmaIhT4bdCzFpNCRhAzkweGsah062k3kk+qTWEDYdT
ZEB120ixJAoMdbdieWHNyOkMVSAO0cj31XN3BOJGSGtY5dWyCXx0GS7AsvWXElMs
vX7qKuQhmCTfwlTAflrccKl2jIKFCxgDCf85v/Q/daQ6HqoCp9E8ppXlZu/HbMQ+
Mq1erExZiwCy/8qhnC2wNIswWAuBPDTyrRbMYPXEUzz2NxmOi6cY7+kysly5K0rl
B+Xl64tH0nzIHGHndFGPyTj40fdY3J+GMIeo+yxbeG/EAjQ95azb5cTxSTZHIwjG
`protect END_PROTECTED
