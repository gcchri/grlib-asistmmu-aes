`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8K3myV9Blhrsd00XdwsggIESO6osymBoA3q7tR3WR4OoQiMM0s/J5flmLZYJQh2j
OF1Zlq+moGXsX6qSaV9/oWWu2L21HbLosi9p5haVg7BAgTA9p9CT1KnMibxWO+0K
NJw2R4y9F6P3e2fL8JBMG7Osn7x06xoG2+wlt7/rDJ9B0mhpVVbc19JIKMRQvdEn
+HNkQePwvx66fFtp5sDqoNiFVSIX8RSREPUDVULk7JoLFHXwOU47PwMTR/Ra+d9T
laa+KmY9zY/sI3h9o/xsjA==
`protect END_PROTECTED
