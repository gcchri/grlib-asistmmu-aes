`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AvrA2t4n/MmHd0Y74yB5BlqOinuqGi09pmkkd2GP0hVp/r30gP73ihktplCn7mS0
ImoYPruvNIviHz98GL+QoGudd6Ox6icNfanI+UPBYxlMt4yHK+GMjLRzie6jtIUv
xpwM6RPIRSlc8PGGmYzFCW4rQXw/lCowCiHRyGZA6Iya7VDFhQ9U1evIzO4eYrZ6
0OOpb6DjPRXFuqJsVr9RasAQuEdRi8V4MfC4qfD5kNBYo/5qKorCl2rRGNLVFPf7
CtEff1gDVu0QjKqUk8P7L8NXvu/C7aaKluJstMcXZ+uZNMVM9YxvpowuGzqdGK/h
pXQqtHIUXxW31U9z/6b9OSOEZ94aZHXAJ06EYyAdqQkzDlJ1gpO+NhkvyKTv52gh
cqrlpseOCKIl4fardBbJUndNY9YHXkc6U+WUyLMMVO3WMrsw4YcJcsbqzMfFO3gG
vNP9vpxTRT7FqA+qCTWYYwtZIczludeJhoE601PyhwG3VSK8U4s/dUQoxH+UzJZt
fqxl4sbWndkjU+DJ5twiMeUYJEMau7zkSqBd4o1KR5sxWt7moImyfUPPIceAktCZ
+dk0eBzUrlWTqXNHME+4NE+qzCFs6aDEKHHk07AEeJQE94gadn5tLMbkiqQPtS2H
f8r+iM6FRMrpNaG7EMRhCxFk+iHx8KoMaffAX/5r3zKvgeHUMOzujYIT4JkwXE4m
5t/nNHq2oet1jw3WMsD/K0kF6KmY5K0H11DLubTUOkmtKPcJ0rsrDLuTp/QSWrFp
vOs3R+JQAAkSo40PBueodNEKMrk+0JtgFn9x4Z/lHr3Depm4pSiPAKgP2/bTG8QH
yUaJLfOkszH8KMMl6jFWSR+1P3OvRhWDwHQPsXfKYITwkA60KjTih7bYlbAQrYBK
qW+FMsIOOyQ1keHACOIQtMXkeHo0RStHOnlfBMT3fqjKfaW4GOT12pYIqtuGd+5j
A4IROGs+ElNtORiv1+aJSvs0XX0HYoHnfyNEoiWn7YC/HAtaDxdq/GIPZNn2PlA8
sdTXBxcifr2KslLVgo/vR0d6miz3t2Dv4AnoQy9MEMMOEh79EMtPgLI8dy6oGuNW
gzV8UmLJHqVxMGLmMGAWFGtTeP9QLKbSlB2fuf6mIkAUyKMW19ie+kZWYNsfSDNz
Ts7M1XqaJWU+WrDGPKy5m1wxctRY0x3kFKuNa5ymDWgLbNntmHSEjhivPjejS4lW
97FcvFeVI61U5xZMf0LMlq2ExQ4BFR47kMMB0PDe7DdlvDGycu8uk17yCkvqlQ0Z
wznE6PQOf/k/v0tA4Z0IXbTDuZUQbS3QMdFy6p6uKJEJN8f2uS6Z63Tr+cuDu4TD
lDevI/rtsH9lD6x47FLdJOX7O+sEhT4usNlIVGhsbTBKwNp4ZE+hwRIKxrd87IH1
mOxdabFRjxI3PqAbsdXvcr9v2gPea1PBvO+NJnfCt0afR5azrETyXhTyvYcP0Kx3
mii/IZdfFVnqmSR7gwyu4J0GvKxUp7vEQgQ/SwXbamCoHx7Ly/gk1RBEg8opmTZf
WCogpKi0EvVlAl18NnrinVDl/zspFksNbHT7afbfeYNRlUY4hsbm2oQp9QYQ6NZZ
VT4fh3ffMfsz/SsrZJeCqEtWpU9Jvtq9hGIAo5vu3L7HkZ4SPnUST1L/s9U94XXj
bhgELlW7y1e1N9OK0thk479+NDsygCdUvPj4qWZEXR4FdSHkHTZeX4yCyLmPI3eK
Ypy9mgMANN7M/EPGp3SeRMO40sY+tVfz//LlHmsNij08cf/WGRbdu/SmzfxQD7d1
604CHIxVKommYJRLvZyD1YIgNh7pwWLx7L9yxme8a1bBWDy90uUWDMUZl6YWmKH2
IHFoGTAJJTf/D3ai+0nweVYAqGEBPZ6mrxK1SuC7Ao1+4ooMEMUTVq/4G4lYKNBR
N4wWzI9SZG6DkitbAGvLU9TpLCmTJboElIrbP51Vn9BOAhVBnu+zk9cEpE+SMAFj
n8pmcjfQKNlppdm9jsMYSGRnVCUmRwutANEPZiOb2ZfNI6ZBJrUNCURrTS3P4PN+
PGjAjzzuzIpySwqcqjaz3lhJQTdJuuMU+184dRJak4VhL6RjNfoWAbdePI1pJIBT
p+YEKRdqfkOe0d7e+TeKCMrhe9aWEespHmH0IBkBw9DGQ0dAMPQTPNep11UGvYNS
StJ0QD8+2+aXxk/8ODWQCFD9Jf9cAT0uiqm3CZhfEl3HPzeg6gA5KArf8DVTYC5L
Cj7MgCyeMbNzZ+NtuPpqLAQlrtkaeI0t/2e9tlWNZcQoLaUDXG+1CY4iCivNsRn3
DmNnk7/hoCSoq/stbYkmAOTqgUuThAuc/LtxvxyhstE=
`protect END_PROTECTED
