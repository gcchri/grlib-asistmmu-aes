`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l1nLPZ+hTKG5DX8xCba37F2W0eIKrA0cVIsH6SqdwF9LyAz7J83rwLSq/tbM9Zew
EFsdMsQfzbG6XXymE4LX8JKvbDSJ2WYUhUcbfk4hci8azcaremhvaMr6XGy4ogct
lHJF7Bmnrc845iXXp/77tHvriCzZrR9wHOFHvSB2yYXaeRvlqXSq9gEUhvkPpSk0
nDcGaHLxqYmYfeNvqMkvg21g8e2yJfMhxfCVZMEzUfcPrjlCUsh0bVtu7XgGcbY1
ZSSBvwqZjyqk7d3NlmlRnrkThNtKObXCrBtiaECZf+X+WZcOJ7d8wQ/3V4vtCpiH
K2S9P8yKLk6AnOvwrhgaaHwNapnOj4n1iAJx8Fmp2caSTTS5A5dE1MpkkX3ehoap
UBcJ+RwNLyBHSrhkwtoFIpl4swYbj9+krrcph2t1j8NV06S/062G0UfLiKpmmz5x
XF9tUUoWnlrjKeSOecC4KFLwhFKwRttXtALXd76BDRWE859DiBLLV0dQXm3GmkGN
lD9JrjcPoGJYyWxpH0OxzjI8rmmsOLTB9bT87MpesCxdGE/VaGSQ9hGhDAvIXej6
pu4BhBxE4RNqNMIt8nPQ+EiavrXuUvV812Ce6gZRerMzTrL9rQskQHKtkKPXkZcI
UtZAvhUe0rMlBL7z4kWsIpiTqKbwSNQm4KmWK9FM/+wZ2TgmIBZpq5oqI+CxWyKQ
y9uWMvE9lUdWCYElc/yoh8DxmHq/MWcI3700FUJuoH6yzlc8hNnkqiaLqubCe/cz
+6WIQJpaAw3AzrhlYdP7VV7/ztda19bOYgyfrsJnhkX9db0LvB1+gCeSjolFjagM
uOQC0Uo+yursEdN5M39tyv3UheuXu1TYARSgQvLaROrDQ2yIvPqXL7mih+iSYIPn
2BKEoj28lz2S1qHL4RVKIPXiCzoBTd0nSIo3d2D9dltE7cfq7q6zgPn8GK6QgHj4
9bE4ZSOJJ8+zM/+LUOTcE+fnBVsQ+iDjpRv1/G8dfi4lVbAtcsFf2xkp8UZCI8ut
U49tqlDFbtNybnz49pNHvRC6wsLPZ4OnZueFUQ5wJRa1qDllPjdXja8SdYA+V0s/
13gcjLN1+HR4s3o04VPWCJ+uS5wrQ7qYfXcapwefcCj7isWLVU9Sw79LUY4pxT5O
to43wXM1+1VMaZQ1QEvbUd9um/Gnna76DDN8xgXwPa/JsBkb1mkVmkA1YIA6r2u2
7NUGZ34tow0TH2iDGHHRDRGu1aytAaKQNFj/BxSFxb/F6aTLxe3A/9R2rY+hHOqW
pEfcovAHurAtnfR/HDQMF06s81W4EvVDMj21mR1Gs1R4YHh84fEO/udnmfpo+k+m
6bGCigYrpvkdp6epaQ+JULBGYnFEQXlJ6zDqp15FH1q5MOWypnrC8jHO2MlWXdV4
E74yCHZXCmRmrte1MuEAab/gyOxjvPSKIgNN1NZY+poJWnwDcKDHVJEjnHzctLeH
K5z1L4yPvggX9w3defLsicCjWwZjY+TWEENG8bZefVwMZqs6xRKlroJuwRLJYRmN
yvMBKilDT4GBbh/olybJ3OgFu2GxJxptEuSiPJyRFTKB/VevIfXYKINI4LdXClBg
0rtFpWyTTrQZUOMkMIittTwVAsZzOPzCObO/NNdzQovjDrFPUT5hx8dIl2fRJVuS
jHOfdUBNpPRzNhHUhA2VSpTkv9pYvMaWykwD+5qfrD5WkrhYHepfqngmdsPdTsYw
IOOwmbIfq1hu70/IgPIHwGRZ07NTXTogEmyjeGcFIboQZSNpYkH3sN1PnawykQMm
tgpzYM7aPlx6dsi3utgdE6REbRu6eBGJ/x+MhQXmcJDc3/v/SHk1dpCP9ZecqJTs
7re9l/vghHMyTzd3PMmBGRD3367zPTvTYHX88dTDslZB8/C0L1q7g85w8cdU2g4D
T2y6YIqEZHT1Qz1HXVv/D66k3Jmas/5hrE+PHjYJarP5kZtEgvioIqeMXTCbpBeT
ttTPzoc9BRkAI8kpClcmoap0DNPOiP3oOns889YPEFuFwKa0B/vWaY0ScPvOaKcK
p4BoG7NGWfTf/7ftGoxUcUOwvAcJ0CY5zViwVWeOeIx62LT36lZA15izi72D4PZz
/eNugCHjo1MAzezedLix+g9KryCPBSyqlAOs0Qk8oWpA8LXZt52+xfm/N8241U0K
z0vwCYYF06Fb28bjS90pV1mxsdX6gSEAL//BlxXHI3EwctWNty+yBaD6PJyUwug/
vtj75DxDEIXa5hLDKAUjKaAyd9WMF6XQ3vOgBe0r6VJ3zoTzzM4tf4B6xiH8TVqy
AlQxD2CDFBB50VmP+K+fMRCf8sF0qJQ9+o4jlXUdsHGhtlAHgoequEhMk3/sDMdW
XByIefDQ0H9vKV6iK3+IEKF0wqs0s7b+AuOVeQ2OuYE5tmsPGyCcgsdS9FZ/iv6B
jvLNSrSzInXOszkFYBUGWD9gflhdiXs0kdOfy7KaweFObkCQ7H0dY389y9K/Kbx7
1hO3FakN9hYs0kDU5h2GVzJ3zapoZa4iP0tSWvU68zi4/EAxRH9VuU7+cf06LErp
n1QvABrwU4LePAip8521yCVyzdBZOP5CcPE31uCW95duxRIjeRRj4tfmJQAw9j/r
ew2QBpD30I8CF6w6v4tjbi257a3SEkDNppAkYX+ZSlNTmBRYGESdh0Nh+7hgEJxb
Tkh8ECct/q9bTEXQhQvYEDHRud8tX4+8wFkgcfYeFQazqTObJTRqg9+5Yd53fn5Y
eAP4vSiUrRsZ+pE2EGU1A7hl/GmooilK+vo2bGrWNXryS1q3MeyJyUoXeuCDs/tH
oPXyhqCzZfM35I9fLiqt/hoXbSveQ1ZkmaA6YKOwr3/l/9osVjfuDJXaPBalquVL
oSUuR+hnMg/dOEQPc4TOCB1zWfuPseJPhc4Y0p8fr8hp3aiCjQHw1LhtJBC2rJJT
1iwvp1leyWxnbOhnRXHCxlAAPVHAucisjtfRkP0/xPSsfUK8yqXI3DJgvpNPkpu7
vWGm82jC8+uOUi3Ksmfbx42g8LmhPGUnhFPIUm4ljHPrfON082vsh3nor94BWbMr
ch8pJ1T1c21noUDtD/JdhomxzOEtJJSeekqBrbASPRBUGvM31Y0qOUkHaeN/4YAO
MOG0ohXHcemCfZo1sD4lhUkDIT+dbI6UaLExyeSBT3TwZk1ulrXWlcI7MgW/89+T
s5t85V8GvikJBTnCLhc5O40d+ljTW2Tel9ure2IARmmD1Gzxd6Nn78ro9bsDlti+
LrOcVxDTY6ZSBhLQmja5sk2VlGUqpweYOIIH7AFEStdE7PfRo3Oghfk4u9aAXquT
bnRhzr4rMYFjCEyfsz1KHEvF9v0DCnMevwbjERUDv1qFzHS17h9fE8dVejLzPcX1
vD18YRQUTYVCNhX1pQTnpq1Lye5t5VP7SOkccdbECnd/z7QV/RJ9UNrOtv3k5ayR
EuFGRzwLANL0OqPF5ZdFtrkjKbimf4oAT42BLDkM888DkHziUJVWEYXLC/Q452oF
dyBONef2aoeKSqFFejQpGhhC8ZRbtOhu4+QusmhOgdI2pr8fDAP0++1XD3vtv6zE
WvPVYAMZpQsVozvMjRfMwtlHSteGHAUUGovLJkKzuZ1Vf4f0kr3Oo4tA/3GNGcUL
WpCE+BoVV6nLTRn2dcVQjUiVXps/meX4pzgPx+5TrU3LP8ukbYtfVpXNbzwEEpYd
MbFV1QvKtjJRZxn58Q11ILQt+IkeNTZ7f4CHcjPrD1z2sVSk5oSmsZ3E0fNhZftI
eJV21XRpZPt54Tk6TFyCdh+TLCThd6ktIghObmt9K/MsM8FBG+xo6oOPZePPBa8L
U4DinXu1+cesuntOkCDzz9bubWrvygGg3To/5DF7hgLSB/5c9WiT73KH/HnPtJGE
rxMPdYpotmyZL/QRsQ/9Pq4KlSAJQ7gT3PUkA3zbUfqSFyO6vUsUVwpDFQIWrkto
fJMCCjZtOzR7VPtu7JZ+pWkAK9XAi8c0ymgfA+irdPbzS+7sWgvch1VnzDglo9tD
cgPccf2J/5r/YztCtKVR+LJdfjaP1ax5r8usx42HoxxBrjV1k9tUYM93+ia2g0S3
9x0IHc6t6ewHYzQe3/xd6zTk7NsW784KPq+O1kcnAcXO5YTDvMToz7b2JoCr+bf9
lvSuZIq3jYVyZg80sXZYNFu7JG/TGorvHEkhGQEX9hEZUtaB8yxUmMHUso+MNmRy
VckW47M7zVhkpWCzBuJr22rEUWZIwdmrmtGFkNzEaRsE/FsQITqYxX1fbgpVcEMi
JK4QsestalgCR+QYHViwLIhkGVfZr1cpXh1QWc2hND9F3sBDu1DlqZH0N5mumIyH
zxXiU//pBElGSRUd1SLb0QCrA0K93jKvGLUp83l0XqygCpEr5KSLhHR5MLyGBX2p
ZlOgrWWVQj0zN4cMcYX4/6JuD1u9bZJ+haRWwrZteNR2zI1Xo5QB0oYqKeFxs01b
wYH3c6JnH6Sn1tTrWMY5WdMlJzoOYIe2x66ww9Ny1Y5lGY+9c99ufUq6IftcAOBG
Kgx1APbriUpoTwA81Hhk34jdTM5WxBmxXR9q6FQz0WVDYAmIqJZ3GEAuc9mikgR2
D2vub3RoM2vXkwsvgIU/56E0qaeuyDRA0iP9XiomW5BhU3lel3dUEaW25ums/V+y
TQTTHT5NevzBeCpXUUCVfpPjabDP9G4zBGrXtnvyBDCOfGQU9XTtUj/Vl7Ma+UQK
Z6aal++ZJUoh4nd6CKBNol9/w/H7odtCx6BHdp6r0M1qdA5ZFE1UBfxqRx6tiVRL
aDR3y7l3jXMPrv9bd3vF9uitgUYVluuiwuUGrygjiV2LriRvoCQkruIP5dl5VOId
NqT9gWmr9ECeQgFRUKFP0z1SKoc5qFNXARpoH40XSz2Eocwo/hEhJfT6cgoS3k2a
lKyLXRN3GNDsOQ7F/nO1L1La/D0WOBRSZVzmRIt6EvTN3DW0kZOC1PT1LicL+NHZ
9TPdcYFqcJDpPYPkFwDKbYQFsU9BG0gh00jC4yHt2OkF3+8wLmidi2oorQLjN4fi
4kbJbn5/vpVz/k6nQVHuLPiAWTP3CRADc89K3AMqdwAt5d/D8A0PcGJubyXV6V1Q
hDF5D5q6gulDEyrA0KpmfAalq2zAZPfhUgAxTxtwRqAHgQNYkGMuAz1cuYNxhGop
Sj7P5OyLdFTk0MDqnYHJnf15PYfT+yUR9IQlorztqb0WVCPKG8Phbq/qIiRyyTBZ
RX8pclOoj2WGIxE0Q7agh4bRmXkTyWYBUCExG+FD7dbBPxw3Hpi8w6YkHa3r74uc
WtZqii1lkXL/kbR7Okwogm+n09k55ms0jBRRMMBpUnSa5SsiRWZ4NZ4o6lmOaKfY
oPBCrf2y9MKCuGvkvHwcw+56JvSSWC9fPEZxeUd2qc8Kxd/Xf2aMMcM10B72qm5R
qasUGMmUEol3rgqhw1Y9Ww+jzmxn4DVpiqhYq37a3T6cOAmO5gF/1OXMLjTb8cjP
BVwh3T6MhVANAedA4ilmG0xyu3g6dh/Adhm2WNLCB0QMC1jYWMxmuHPldrSstBLV
wNqUduqXGO/1+g63BV1WbCKVADQpZui4oqLFCSM56LVEdiyuwvSLp6mZ1OLeNQ85
ry8bzmc+Ray7vLh0Q4S2zCRc6f72utELHbdm6cZvrrP+CRn5zZps7u7kOm88oRJK
sW7fzH6EO/eRSZpGWtUsqI56C45a0x2Ed53LcPADCZvdeZIGCnnKDJEziEIC5bsv
ksx3c44qNu8TM6V9O8gp6lgonmKYwvToRlYlBox1YutDWv44rZKPGhw5sQKDNrLn
E3fRta2UYIO4QGAU8LnoRvzkUkRkC4wrB9cCwYSH00a5idqrRhwp5BhUIt7ilx6m
TvEfI/VQvaCp8/6g7bHdXCj+E30OGkkS39FP8aTcqevphk7GK1WV7woM+4Svqty8
w0Zyqv1/a7enLCWGoPWL6IzCpkqhGlC9k4rZzL6oiF/8Q63LN6Yy4KDh73mu1a8p
3f3LS5eiEK/MAW8BoXIXAGr3DNYsgoDz6BGSGBKnMyccErygt6dgD9EaVogJHqhG
P2p1HEakzI5Lj31NjsMmB7cr5Rz6jbXBhoBY25Y1crA2y03xXuGvH56LwpwLMI8C
Ss3fhuB0IVolta/p4ATSFi9GnSYzxuTVlVwaUSoiI41xdPUEimPtquy6xlRDKgfi
0ccQ/IWyp0PTTFh+agar0gyFiDAnB4tjDRqKW8qXu2MOKaj9A0m35V4tKirXlgEB
T6VyiHlilvrgvrl3n1bdZ040qfAd8myDUt1AyMtE136YqZxvhglJl9JVZsU0brKW
28bIEkYbjt1DZB9Qw6DYgIMcOvhpIDJyb8rTsGJwgC97H3wFs2HUCSLg+sEwCc4R
ttYcL2enJ5gUR5iq8u/6K8+3hrkAIHT942f2IiamORn5uSN85Y47e4pc4QGvdcNS
1mzT6K5AyUA9oqOMReYxz7neIOi2Io5EM0wZAe9jkJrvOeOo7FCOR5Ugg2cN0XZW
gPxE6gNaDiqQ7MDoqnlrc+JTt6InrKr2mfGxBUuiinf2J1vbLu9jxw0BG7XDLq30
0t8i29k/DavpfJm2akAQZIZodLaqSrdTRxyww0+3uIN9X0kXxKn01ZEYDBI58OXx
/u4K6Oc6a/RNZJ2VpFUHoX6BtdPk813nRidOcMkv2UyEN3/Q70iK4C117mVMsAFe
caUvv0aZapJMXR4T2VJqcaVbVi67WShwPRbGw+WDqClB2bvdN6LJKeEN0TQib2wS
xZPDbnYF8yOsx4Bqn+ckOP7p7IauwiTbfQnLxBnAx8y7bLe3KjpiKzNTEpyXJQMN
uogWSG5rEMRPI0YW5WC1hxvZG/yg3cSfvKYELnPlBsRkA/0HhurfUwFq+nNQftMd
SZqGdui61JDoGNuC1ULTJAA/3RH0/H4kOq7DG0ztIshAN1fw6Y0RD/kUgY0laRbc
bBL4AQKVY2CT3cIXTgGs7hiXrBfTu/BQwdVIArc7N4f+XKURvgokXrEL3Ph/eIya
H8kFs/dGH6wDM672sAK4rPPjTdlEv6PQCBZsNq5byMmp6JB6FLZWt98BF86xqk5W
8saE1GmYtFz2utDySzSVyx6sFd3VxK8GK5g/yX12H8Vs/bB/j75CB8rhQkqHH/UV
j6C7jx69F/TEb5pL/3B5V2a8VrO9RJvR271wScS2M1F0LN1CblOIbLhfH83VkPU0
m05TnOjrB6UKigmE5QvK3E1ufLnBcgJRwvHrPnGufWki/vBpH170EGB67Xzz6pXE
Ny9wqtido62vJPgnrfOGycnx8IQmhAEsnPJ0pxDgTc5B2G5yHSA6/VHMcLOK9+WO
TijLw+S73C9Yjwt/CHgX5qn9/Aa/+8gW+zsiVR4et7K+pBxVD0m9SKfHymuV5dKD
gcc2d2YrcH3FmczU90KXJQYuwnjVyWbAqSAGM37S7AhVegDIMAbn5ydKzWf7I5ZT
DVIx9Iv858536H3txq19UU19x3p6S4Lcq5Qj+3WbooRfhEqS20A2qkQC5D8A7qZU
U6B+2+Q8gbge5i3UEoAqyHRIcCADRtMgr4CZnIKdqh7kwoP1MHJV/SfLdNsksjBH
fQTNIlXFcfUdjmc1x3d3q3QTZZIsPHzjwIfmgELIuoiVf+Q01Kd3YtUuy1OOssX4
x92DNGmvDOFxLTVTLpP8u+cFElIq2sIX9jiyex1U4Hljw9zWvpK4+1UPZbwQo4dV
eSpeb82EcautA7Wu992bi+nvVhV0imzwdeQbzqHi8hisVH47t4J+i/xkfzvEjnvl
aShj4uiQm+VccJNUeOAUQBm+CdpT/GAWLAHMKcVHMqdIJKG2q9IRxu+FNn6d2AN0
uQLrZz1GngpvSpfk/ipHqN7jqCewqqY7mbkUHgGq7XeVDX/jNwceUtjW3dTG88e7
2Qz/SHvrvvXKteXWGPPoM/+KKcV1GoEUQ/7pm6Z9W6ETQjVo1m3rwg4SFCw2kEPC
yzCPoVRkDdmLCDU40lvLoHsdo33Re/c6riavQsTfQuDQrZCp+oBhaKow5W5L3Rhm
jz+btHlAISAtefa7psoE3uO7cYMM8wQadT6gJS3oNgUG0nJOyKYu55YZ+Ul5/DkQ
PKWfiniXSixMmzGuPNKme2UFWx/yotWotCD/ymoWPC1o6A2suJ1OrWoCE82aY0LD
OshPbspK8ZHiwhHx5XvbD8cpOpv0yD6R2eB0X4WGxhtDnXchrI8zLs2OcQw3Buu9
b/loxsWxR5LWjeuMaIV6fXKmKWXAfTUUwwnbLQwERp+aB1DojLqHPVtAHo2FokbW
i/uFbPEX5v23hjd3yPGj24eWufHuXMdidhzZ0QusXJEZFkEZsqhS1SBoYHB3ld6o
VEmn2bFz3FaX27DUVrpDJMIr+h4PJpwiwtE7DZaDOZMB1ueVdC0/J3mn/2dtLoqL
CzP4tWtlUPL8ZFXF8GGiZDkNn2MMPIa/nC6mg2qe3gFVJsogdUbtu9K1L2/H4aH9
`protect END_PROTECTED
