`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1V+yRnUXDH7D3yC8CgVcydZFLZNZU1eP7QELfWJcrTGNlsFc3wJ6cSvVsVUe2EO6
3tfPE2zE7cOetvTcHsrm26xiAfQqSp0rJkUHsKBFHejUwn/ex6N14//CHB4mstyE
SL9wNPYcfdJwyzv/hruPxmtrU9jMUik2Tp4x8NJ8bMMOXDwHfiRqUbRrneuhzFYa
mhai49KYSHMWWvoX4SY6tqR8aia5tJhIlJMzr75r4A3TNjSsoqbkMQn+gjqowynC
p8fayplU5vGTCDh0rA8Yj3Ra/uHD0JGJA/9S/WSGmDoikRVdDC9giw+Z8eQWEtpc
61UuCbywoK/ktueHl8GnfgKeqQZA+EagS0IjurvY24cEDwHbWQjShXqZd5zDYeOB
G6AfPIAztIa6+Euwy3ymgCaI2YlCS81sFuFzAc/Azg9uawm+/UVm4+sNSIwomGnf
GgNmtSfYS9M1KTcCjWUlg4jFBXuvfWQj04v4BjeQWxn1I/U7hfCJUGdV4Xcue8LA
cAw70VMEcKPyGWPlxLjWJX5fHqGOlvANSVw3DlsidDg0h3yZc3Ko6SFyE9kySCwQ
jP+VYf0gXrASmJiIhp69/XRHNOX04Izi/tgYLgbdslwDDEPp5IZbQSc4v/pxaJXy
6ZluXIznuUVNR57rnQtkpie++fpHtjd2DQZwKfi0fWoCckfP5Qo8cAiQ8URR4Vwo
Jn7Sh2jOmsgT+xBKkUbnGe9+upuvvAobgOL/yff9A+d0sEsJpYKhjELSw5cxo+//
t+Ma0g1HSQ81ezf39+dRurkKyae1b2wPvEM//HB7dR6bGpcOVG5cKPofYNv/Ft5k
VD9mwWV/Iay5pNhwIAskiliiDpqr4kDQu/wmb5c4bXMqXn42lOXrNbS8PrqJZvBf
tEN1a4GqFs5972ljXehB4wSATBsWRgS1IcOJdtXAV9FD8aoKIyL+qzd9nSV+SzUx
AxgoX2YXTshW4ZSlOv7fULiTdWt2Cayt214JlZs1iPJaK3H9foEh4hbH57DvHmVO
Jr6Bn2ujSMlZas+Rz90g5OvLeSH4/h4YwGbqvDhvxqpzQzkXs76/dO5TtV0e5lEJ
CHQPJklVE+tvq/JmwdYCcD989O8qPKlLueP4GdPB0TeoA4Qi8dtAt1MoXAhV44nJ
27TzQxvYqbQ1UgdcOUlLUJqQ/ttnSuQ8jSgnYXoMY1Or4TueiGut5cQ7A/oys1nw
5Ul2N0tIG3f1J31fd9U7aDvbOWBXvFRG7R4v2j/yUcpDK4QTBrBp05nF9seR4FyW
1cmkLCic/yoD2gOrO9A5KNyx3Em5LRGYh2ukkfdtl9Jss9fFQFYJ37eezsDlN+A4
bz/MrROq0gsoU3+wnmFqiI5VJ22HUJ7VCTPCJOXYIhjMuKSQzd4y/YxzN2hH4/on
PN5Waj/5YYXiiRJrpyjPq+PKr4RKSt9I8I4FD+qaIA7rWywm2s9yw0QeDe0VpuyU
e/rL8pftyMoJBwbAAWauV2OeGDanoABI6go7QY7AFQI/ms87+GQ72t27AGYjDBZF
rRvso82fuWaIs+AcdZ7c/DaIb49tH03Gl4oDYiCkrOWJtjJpBluEwM93q2FmxEzb
nZZ9BuZvTkGjyX02+JUzdA3ofLj3FkSdRnnnHg8TIZygElNvUf0BJso40lTUzhmn
2IOhBFZiV0UHmqX+dPIDpgRb0WiD+BDokPY5D+nQH+JPDQX5TbUbgzUkqZKS2YYh
cGdkTj2YjmcKJwIsg5+UmrUl3n7m4qfODoxDCyimlQftubrWXLyWaUVFggYqq0Nv
VHlA9hC8CRYRcr5NZQ+YxTRhQA3hriq4Alq1S9jEOqe9BH2z2DWb0KjLkKp35obI
1qiTkdHKMtuZKQvEDaJ4h5A1vnTud8pwGFbflQpsqGXJLtCuwQavEcV3wYCyvcli
Yu2Oot15uGGW8n1YnZGjICu5DpQqtWO5Vfo4DMHTmbQhNUHzFG5HftIYQJROCFSv
ssGf0qVh7T5dj6qChM+gGIexzaAigQljLGBDff+5etqb0pEYe8agd9SCNSWLjfKs
LRIM6M4Xn4wlexLF8vlvBhA8zBalr10rSOLpSDFwHBWxkHN4cCJnMC/j9roO2kd4
CZVw/6nTfRvCVDBmcPPW9sI/NTxYhHB1m6bpWMpxwCOveTla7i4G7ZDAvllNJuD9
IFZKddTRP/GDc1+JjqeKgjyZWM9MTE5A19qCDLlZW7GLBh7rDEBhfOEhi/4Ux3Sc
jl/D/ZgoiphBRrtct2OMHiSVg7FDyKamNmcBP+fpx681cpl6SlNTtYGfsdE9y9yl
yXWGu3BgyCU2OGLqeeedMdCZxOfJQgmbZO+2ogLc/KCiXJBHocWpKbzM9tzzwrQV
`protect END_PROTECTED
