`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HjgBgNhlUVg4KdQtzNDSk9JPKSECs7207TxRFY3yK4LO2xb+FMfnjynCW7/Axx29
4+shmWlA0r85/x/7WLby0qjm1NiTOEWI3+wrfWqNPevSAjcjbjSDnDPBk67bXDUQ
+k8rLLQ0UgFSFEFkC9nB9aS6QJhBY4M9fwFT3KgvZ3OhDOQiGQKYTqZLzgDSnlqR
ZW+tjQYWiPwbDjmCprOv7DSxYQDOzZ8+HvNitu/8PYgbLWNTi5tANLpoJQTvpV4I
xkC9PTVQ1/hNAqbkPk4z4Y1i+r+LyK2IhIzakyN41yA8WFIj+jLiOo/dxf5QdmVX
ahoLpn4ULb22k/B6SSNAbGhPsATNXSVwBw/5OFUu5WRJqEPZa95BnhTeTFduthnD
sU/Pdy5T77iVz1QgYYpWo6cey7xrskpwvOVTcmhAl3eXkMmDILG9AC3LmQ4OVdTu
x5bdCRSk8lx1lsKd5Np+tA==
`protect END_PROTECTED
