`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QIZnPpJ34J/bTv4ofxsYSRHrzu5joEJj5dMloUICXpsYbc9G64HeW6DmJyPGC/Qw
Ln6W/OBO+49roPczfPrOIrGXwhmD48aWMmMJDSioxb5MH5L4BBrOSZsHH52522hh
3jRXwqctH5/adjW2KCJUQ8NRe7EfVajo8Ga8aMBNpVgE/pX3qQHsbsqr6cNu1rFb
J1PhHvQzGapEDbQyRljrNVOza1WMrsZjEzBogd+NdF7KFcCbLouUfotVaRf91c+X
f/ZARhX34BzXjGrgfnK8hDFF85QClKOaKFPGyLvUv/j3IEjgTMPI5vUcOHWEmWDl
CHZ5E1hkrpZ4K0wxPfIT2xoZc02K0lG4xKdX/QfAKgEvL7FoA6tIL1yZrWBldBW+
fudIgpyDfGnG9RJqL7EXwbVjiTe170y2Rh3bPIB46ymMfk3NU38p0LZ7K7dLOEdG
qVF9+UAhRviqCWAJHpWildubLZnZi/J2d0AsxGXsgZ7o3KZJGfhLQ8O5C4X+2AX5
DDZ1xAmKU9Cl2Ti1SeFwRejrImZ+WXDHntj8O2/36erlxLY95e5ARcp9ylxiQHJR
ywkaGDw37weYUItVQCn3kmY0MhBeGVoV++BGEZVAZFdhgIJiUbH2TwmWvRKVojrq
fvr4CEtwSfnbG5F1ZKB+EA==
`protect END_PROTECTED
