`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W6Bku77V8fKmAVFg2GmIApUCq0l2SiVVkQsHd9PO4L7Q6JtX7cEGBmeTzhD1DJRN
w34y4BWfmjhGEutkZgYcuHYoQfvqKa9WKsFGmKKhwi3IYVwQFyfx+dloPNvI8t7F
BgZHLOqQWJZLyh55McobpipAFXXwJFGjsu4UwwJzuTzUKNSk1/0Q/0kk/RjQWo19
t4Nfnb5471tBk5k8q156oLI9yZmjVnBv4jN5Pfcq9M8uzLMt99eLjsPAVq66tz+3
59afKaxKbQsBXWaosZ0aQJkMRPEsYtCs1Q3O2PxzR4bAF0Db0oUXBc3mkyOsyXrK
v2TuNcrY6N22NPdVUU3vSSZsnG15WLXA1/puO/2GwHFhA3TM+1bbHo3naoDgOiUm
5sThiDMk6HJTNiKUyJRBlYP3rxb6EFPETp1Pu57tqUtdi++ULzn4nBZ+zRP8IO1l
QovOCvmjfXymY8wMcZQnLoQs9ZNZv8IVEhju6YqUATikpwDf+PO8tWZvQ+XztoRh
CmffiXxm2YZ6Hex8S/Dz5BpynH+5k535+0IClVs8DNE=
`protect END_PROTECTED
