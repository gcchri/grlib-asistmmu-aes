`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SPliBLfdmY9Ek+C+8fUmeu+dNZ0i2DPDVB6sBEab4dG2m3ska6LtBoEfSK8Yw7v/
9A+ahmMA0BEYeWDhFVm6zx7542iuuUZSUWurlf0a8EH/Ov9k3CQlAZQrFGlBWKoh
SHmczELBLAZ1v3mfcjuQVCz3KMAe2IldhfidawXL/KFqjlS/V3CQgPmQT0iAJfT8
cxyiorcO2P+obAQvJqg896uUVc8aQz8Ipyxiaud6kaoU4EPwzGMVsbkvg8H2jnkv
KRMCUjq/Ndtgg43Fmz0AXvmE55fJyBswDclHaftPorAlREOPW42d4C1V5TfWz3nX
OaO15/DPVckSvRGVzpN+xwgSmyKOwdAa7FaMmoNKf7lN9V5XyA1tX34gcrEg5Agp
fTF5DsArzrnQOuEX3puHD4VE86ilbVSiTibJ6fhkGghCqest27Dm/F2S/JKvW4Ms
OH54uLjY/IXv3coMwUSCO+dnBBHo3MPekRhj4gpUtTJojNDI9f4ZzEbrCehLk4r/
ZhyU6NPKP67+o2B3FRG55ZUrsdJUi3pHDc76d9CEsBJGLSq6yw0LdaYPlAIPgo8F
SBRk+jKO3u7pFb28AtDeK7NPYzC8H7dzGK3lPUf9Uh/TZ6N8VdN6GSq1bA2fgcIP
vIHYVEuE08GUTCb22pelgqZAY5a0L5n4iGmvn/AVHwGtlbOd/vFgmiNyOAuI1iNa
7KCMEnLyWHLFn2ytThggrvLr9zGJIEWeb+Fp/7aCrHs5HkX/OvMQB6YBHglZxvVF
Dr7hqzJesm1zuRVXSl7QUGQLU730jOlswrp0nM6PyXXYaw3J45XPtWHH3KEuoG6T
MPO/gpd/R3gRJyBeW3F6O4UD0OcbkF9IEzCtJYsiuFOKyWFz5dG/WmNwsn1Tj1XV
HckMcjQVgPLqVlWI90HHEOxVAXtVaXBbh8ym296DtK/MJEZ0RfA/osIcceRoQWtu
AMAC1WBL/qxVWxApgM4Mvb27gkI6CcZD6jzbGz1w/MtdMzepSftK0ak4d6uK3dDB
uCqibCH50ThmivP+4yKnuLRHukoPj5c6V9qpDYnDLtqKjSnfRXCG6hEVW2Haqr53
2gh/ca+uyzwpeuo4cYrA6cNMM9nN/56feKen4VIYO7Rq8zNheGxv9SrVy6tLVUK9
Czm/IBCqRZiysBPacqskyNrKk+HTFDKRgI3hxg8m/DQZsZaR93cWhKlrF0Z5jZ3r
1z258qzL7LDQvizsigaaF0MhpsTVuU9XmqL8MfvnEszGk68vxWaieN6ih3NXme6v
ERRhrVjtca4thEgPZdXU7Bnl8BN9EkrvGaoQIDDb8aJEhqBeEiIXDxBzdM6fhZZs
hVd5S/O+NTyVMDx5kXuqax79tpsjNPbLUEN03zSnsLw8zeOFEStMwyaN6FpL0QcQ
llgtCGtKZEhyJfYtc8CMW6o9rPxaITJnwpwavhgAEYD8tCNmVrqhslzlbxp7nkuc
Es+8YnwEs+EFL+VYEMlY4ivRT5z/WLYjx/mr0C2qkpH9NTPNXoeWxsXtqpEDxpdu
uN/ITFD3TdRxoCSpanXVs6u23w3MCq2c4z1LSig7tbzt9kgimEDa5cSgTzYh/GPE
JVMB8hbRvC2JCiubPl9sKFBtUJmwXR15U2VGToHV5fYgTbIQHSzhiQdpoo/cl0+G
mLGJLUKESxA2kLW5BUsNJnYZRssi78nqvSxqDtQV9JAbCHRc9IAudhSx6BPGgbs3
bzhiMBjoDwsqN7wO53QY/TKdJwQHtbBv4mVKd9YKZV5Y71eliUVALrBEzIviLaVl
Jj3660mw3Q4yvkSIZIC6NBkulze6ynuIri2pBPvS376o7gdBLsgjkewscBRJdi9u
J6k5Ijt32qlJi/KZmbHwbJIPlD4NSME5e+IxuOzGbQwJRip+6Oj743W+82r30+o3
XjNbjwCBpXFAZNi+H6VRlmRbhtmBWhmLDAO2ME9EL1BBx91mPdpJKJP+0QcjCgHn
aEeTZl3XXTDpQ8bd/go2IcNn8evD/nq2WFetnIW1Cqh1TDRJkRRiNr91+sjooX8Z
F9W6vw3nk1bDeHf6OSHglPp129sGQ7SVE/hjG8jYJratRwg1s2S+EUcDHpd/uPXE
W8gm/WJDF9iFkhOS3s2YjR/ae+egdJNaHkLEMHzGTQ8bGQ5DLs/17Ub8ZWO7XYyB
Ne0dbpmJlcTfFnrKkOeKN+8gTN9x4g2UGvQ+ItjzNdMZ0YEbxW70qiY2NiJtGny9
uzZENTPJkzt4EBYBDhPcSZFCVSklfafvCwCMstDBtnJe3acDtRMd2ha59Po4Sqgf
px9R4lVJPKcQ8ZMKLPDLow==
`protect END_PROTECTED
