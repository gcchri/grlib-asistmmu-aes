`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bp7Bxy/WwPLogFt40Q3unaE+ay00AbcbGU0ILGpbKdElp8/fI2t9i/GLseI82Vri
Wh9WvGz2L/QRcOe9F8brflMj1rbsv1Hrh6YsBsIHDM+cpkN2PBmgpMN8BuMk5Lt7
dFe+kn56BhLJrMAvcQys83VPWWjEJggOFUQssAMXtaEkqJ0yOB7BNIECjmTmr6UR
dvrhkSvI8KoWr/dYMYhk+B+Gxiv3KM8f83ELbyvxW3dTnHRV5TSKsLcSCmTkmeg1
UtQwxl9MxC9DIG40aKPDtgIiGJHDIKcbq62NBmnAYwz0GkrKrBQSjcFJIt7Jb1s3
hhq5YJM8++e2O3BFKMqiBB/CB7vYo3W5RnucesyeyyZmEtiy0ZtC6AFe6Su+6rNh
dT9Sd3vwlWgIhROZVVgkJP/jkI25H6OavY+/ORWKRXw0gU33cOfu13vT7S9WbCOL
/XPNsvmQnjVJRlRurosRUZHfDxpFOleeBCkL8PFfZpoLcLTXGB8ce0AaNJzIL5S7
AKpg9WoHAUQ0NqgstyG6Obvfh6RHPRgIFAaxYMH+Fd2kidhWTq+GbkIk+qL8v+Gn
EqtI3jMzc6oNJRQ9W7jQ9WlGXavC7hhbSZmjvxl0TR0=
`protect END_PROTECTED
