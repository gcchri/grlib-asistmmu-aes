`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gzl3ZRO7R/QL1lglPOOwYGhpW4fpoE0z+y0tz8ak80NPzwihL6qRq+sXUmMrSVsm
ndICMpTOTxtwRFeI2n77DXsgRoeTJQaZKm1g+hqcKWQ0WaRZWjJU+kd4G1SGso3+
vaCMmHKJ1s2iLCxHfUY4P24YYQgLqIFWpZdNQe++GmavPsxwF8gx+5NEAK/9M2QW
kw0n5ObCPunVwnKLHZrTmYfHPu3pSWhnTSxv3/9L/xHcmolx04Iva8QBXniAO6TG
6rOlUCdZtdXT91PQGC4BoOjvvtVPeW3T7DH+gg+zUOmnDuszum6LSR0ua9WoI77q
MEQ/CftH++wAYdH9RDOD2gsYgg+KmHX/WxzoMB1iDRaXfIrgDbo0BXsHr6iN6BKO
9tSDDE5CEEHGlNsQcEMWqmCF4QCsP+SKJX47bwJb0H1YKQpLGHhZHPPMBKm6uamd
5XhWM1qpp6y4cal2MSW4FywVUVIOIMupdvz1b1VxsPy+fl7XBjYIJudmcfk66f5N
MXB0wMPu4NvNwcRjjmq55n0IFY0LffNKArX0ncQnnJxVahKM+Wy+SbkLBMQuejX2
dlh+ePBieQzYwGejunmIKjBcN7fdwpcMErXCXHcqt7YVQGZeasEJ4Vn+XORe6hWP
0BonaUrj3vzrn1Cwe/EvSFukGcqupwllwsL/uwEsj2c=
`protect END_PROTECTED
