`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KwkWQAKVg15Oh8ZpxLJhGjlKQnmK9A57+whPyFlppj4mXa6D1ZpToIH4lqNd7jDP
td5/XCN9MDAP2i8NW1G0igqe/YUhIEAH3vLidcj3kmi/vibMizOTRXEBcQGoUPG1
Wpm+FXnrfA1kAw/n4z72CzUj4Lm7+Zl2deE/+BhB+2sq4dQxfgbakxR3pN6u7ZTQ
Izj0c5KVZORmxgySj0R7/DpRFN3jZoOr1t90JEhcJjeTxaCm6GbWqgUlsC7DED1Z
4Fw44VIw1S8pMF32KK25Ptcg+z04dtdCGIYVk+7evDyHYxN8q7ppU8gWBuocKLOZ
/UjU23R9Melh5Yi6FG3BkQOEr0Ahjq7URD8He9/pMK7ngsORJXfVBQb1VqeQ7jW3
UxEjSGfp72V4CWXiy+JI4Zop7sxW3STGI8nXGhxD6c8KIWXp4DDs3w6JxveCWQij
`protect END_PROTECTED
