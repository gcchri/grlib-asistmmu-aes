`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4BeTt+HCV3xac70YiDh8hHANNi93abvDTunOApx38ec6+iwYXzVriH8tictgv8gL
uo2Jdr0WPHl+F4WWdJOb8BPazjqVddcquP/nGBzYU9z6obEp9PkTFS6d0z3c+Ltf
89quQEMNwqAqEqebx8j15Dm+Bn7UWCPeSUdOpUojKEe7RW70bX1niSDt7qndtBh3
UfOhFYEecJV64juLpGkh9wjc60ssn7wvqiS5X81teFbUuNzd+W19dtCAxhTnLcnL
kbqbhnYL967stckh2tv9MtVG5vNoo5qmq11yaA5t6zcCM590BNVgdVtS86076Fbk
YinTjJMrmysVDmfAkGQ3ob/MOBkRcGGFvP8tZa49we5F+OYvN1LNei0dm5f4spKN
dMVFcAa3/lZdy43H2yZnTrklP9QsDRMr0Ftb2t6cpb0vFg2kuwDy+xXMB4d2dndE
YH54PUPDm2tekAUEH9AprCSW+FaBXcScjRu3fU0H0wzAAL32t/XhcLxd+vSu/LaU
2lq5h4X2q5RfG/+/mHTb0gtPiZDSj6SJ9PB2/kUzjVoPiZFkr0T24r9ifnv9iwsJ
YQzpXxcleR6Eg9U7SDbZg60HifgN6QgMXwGhYQ/ttfKMZ2cc/YLM7jQSo+XTSHUj
1t9ds5ibhrl2whseA/wiiu2O8WppcxuX1FsHgaejulZIW/a6kRUdSBilepwxkail
`protect END_PROTECTED
