`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vfNW/2zRquBYKN4fxC/RfIUjk95NZfxQ+/L0lsqbn4cB9u78Ll7NHfuG5xdWsYWC
6IlwzbPnpVzdXv/IfoDu9U3d5kBla95/5hln3Srwxj3p1h0/5vl6pyenUQfE0nYU
b2zUluX1JzF2xtjX8jAhIBlCyZyevvcbkZl+Td+qYCV24RuVprWXHd6mdwgXrdVu
/g7iaQ2lXgMK++SapoYj6ByzKXWJF58vI9WueHjtUi3zlcMn6UU4s1EVzdNkMZX0
KWtBfGpBm+c08WdkfX2BhCkRSEF5NBORH+3GLViEp5BidJok1fpl2MeNtD8Mcmig
9Lu0jI/K3a3EOfen0VHrguaUqYLZQaQ36QIZZEobldAKBF/F9rqm1yzw5A2LYXH2
QgSX5T7D9qwALoUDF3A5I1rYM6v8f6AUquPBFqw3sdJ5fi7ZocQ28kCQon+zXajt
mSRoZQpQYw7CrlCn4BBYSKAZUILcYmZJODEIvhK1AiAIKYVcOJjDUfWYjwcH4tR2
RXsE7EJWWYY5LvACNrY6D3rMnB4DycnaBwxCSc74Sf6wWlickLeYFqvbTdghJ72D
LnKYzYYfdOx8TLtaxKASbUtVCT4dkCoFO2Jiz3Alsf206ao0uo1sD3KCpH+ASYWg
QOpRE8EVz27sXRUMVpzizlLsQUDoIhojr4QnPL4w68edV/40I5/u9R8AtYXbGYvm
HnChu9wIfvOWaip8dXcyxSxCiaiX+uggp/A9hRrOzgQ=
`protect END_PROTECTED
