`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U0Vi9g6vl/JDVspSYRs3pplKpBlPSIhZYZEZp62HdFANV/75SfSUtEClVfWdoUYv
tMlrs6HjKVBWC2sk8EXMVtFmj0FThW4GYxrfNEEDHaexD50J/X3eVdY4HTwmsnmY
m5wKCD3tV7BmdzaYIc24kXvCccutaOGJwag6qc/9Z1+Fdgi7O5TxkkfRmPNrz7dE
2bsS44Oit+zCJdZ01IxwN712JsmpW7IS3ZTehFuz0+uYsGR98zdsNiHh49vcE0AI
NfvG0JxdtNd3krYkydVF1+TOIznr/dt7Nbp+xPFEqs95v0zOC2h2soxXCL7jNDi2
UorFIao/UFbLvRcBECN8yK334JJZ2c9DqXi4UuzNV9EERE7Y3YVAEFd/vhPnXPXK
mII2eMlOZStCeOlAVYYQqSLKXlJ/lRzIhzS9Mf11aIyGU0AbcZXk6slU2j0zgYPR
w+fnJ2QmGeezhVHXbvob49V2UfGSEGcD3sZn2O5QOKFxjSNBqQoMs3jplGYzvPl/
CQxk5yCcneE61Sg+jv57W+iTOWO4TmQ0YaOha+HtSxTsg0b3KnDxAyS8lhHk6nmT
IT9YrmC8ZWEirOun25F0ZTAmhlzkl8BTnsJNl2TRamYSbkXvlBAznaBOPQxUOAwL
hYsf5b3SuF7BvnWkSc4pYCsWB3U8Nb0nQLiZN3B5Q+nzd3LIwBKOwENzXlSJ+iSB
yhQeq9scd6NJogHb+dqXXudL1t5m91nW8RGIdtk+OlBTRKlHiWnSHkeDV6cODYof
xcIaU092sdAV/OwZG0lA3h0O0Y8Jo+xFOfGhcYS9uXI7zQ22C2O67x7L9qCxoV7J
ICDLgX7wZjaJ28O2JlIrSLEZbudwV/ebycpVl5NBd9w=
`protect END_PROTECTED
