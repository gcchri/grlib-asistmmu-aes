`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y5Xp1fzZ8VTG2VZl/08IgFeBCcsqLxytnJXkl6oa19X28nkjw0XIBQt2FFQTa5iM
524cpaoMDVEIm3Gg0AMP0BvzvMvEPOB3Ox7NwLQpWfCSyxubejGaOrOgHZUdyRyF
ghRH3wt54Py6jTjAewye4ygPJnVB+UDtvmtRxtnR6ZYszT/9LIWvSSX1iMBukG2o
y0bim1RtNTYCg5Q1CoaTHpxG20qjm2gf5U3Db3r2Ka3gQwDeNkyyK2rZ4d7ign9w
Frn4XaHmSP6W9mkgQvEbhuLpe15B7/imOQ8SsK4Tlo1XPWGVlDnwSCea3QMQxoub
/Pf+c7l6mUPm2RfCO2JsCZPOm46bYvxhHE/tRJyarIUo43IAq+aPVfmHfaoIbrNj
OmCuKyDM6rziOIh61fn5mjRTMU/lDiJ4LMD646KESF9wfRDbUy9UYxTgwlLz0XIE
QmDBcwmk1Gj7qdX5L9RodEKanf5i43mY4afiMPrEWNj0T8S2G/iXXDwtE6IMNVEK
rXPJUijt8VNRTLtObkc012+Td5ixHaDeM2RqGYpKjle5YIIv9ICnKVVzCYT5SEC4
vdVMkEDC36KGnOh5VwWJJEQ/C7YvPxOSJeuLUbR+n2qz1CO79qr34GTCg9SrQmHa
+A/00M5VuthKllsbp3L09uTOTXRXmXfgn7ceIfIvkdkhSrILrkhND9PiZ85o90xd
MXUmP8hcc+Az3E7VyVsTS3DzEkPHYSdPfu0MosZ3UKsWgmqxwYWG1bQ3RbqtjATe
hvlLuEfrfQFU5T5aIFPPUK/G8hGDdxS/g1olQmb7py7tRsSYcy1hVERI3x8AG9V/
QNYGdsRCYIzyN5YI1bN7l5/LwHohiWSGiTo+YdLKGjE2j+DjLT9XyprIej5ufwQT
VpsNfMfdU3N8Aye6zQyqKw==
`protect END_PROTECTED
