`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YBePo5fGETHK+jSetb6EmbTFwUhQa1zJ5VX1hMUyE5OdUtJ13wvlhcbd9xNalgFZ
vSsIUu/4pAeQJO/8/FoMa+NpqPCTpN70ofsEpguvsKrmccqwKeLHCvWqO9ku0afs
3nooQ4Ew14/RKmmbkE0RYhTban13uiIbcWBAAf+hny2h6BDmquOO8cqkxItXpfbq
GQuTP/FL8817TFghvqeWCkZxi/LNDMeIIrJxO5LUeK1Tka4DTAlBcTY7lZd7eskX
rhbewO75Il5VIQGdOndvFYXrV/fXniDBtn2FNheetOvwg07vsXohybC5xDuQMUfx
Z/AGme5+q/pEw9QkWq+fv/YXK9r4m8v0/yb48M/BlrDoUEi10BBhYjxHxrZ+Zb2J
cXCFEbhjFuyQUmUN50SYROvlJXqsHcORhVMqEY7Nt7Sf1LTp5URldMvIpAjuJTil
HeyCES2U7YOR7BrYiwHMsqYjtV8ljLA0lhO6rIU58bVMN/B8NuD4s7g7iuu0xr9U
BOMx4LGP3lRjzjLINyvCcDSUWAYPsFZTr+AQhVJ/0cgT3L2SS541gevkYK3VpTaV
dGc/sOeIWYv3lMNKzYN7xq5oxPTvra0892BVZZtHmJU=
`protect END_PROTECTED
