`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aA0LxmOSNnCkCtJ4NC/mAkkHngywRr+4/ETISf+KiHK+jH202QNK50fMd6TpStbd
8VmiIMdrBVo07T1Psj8/b19Ni8Rh1m2m7y9vpyVkYAvM4/SU4vvyd3isgaGMtG47
mMA/2h/iBnlMEzJp883xyWgGLTDz3ag7wDSk8BufHaM5Hn2L3eK9LAhlxGGxe7nP
6C/L7A+KO01+R4wRc4+2WKPrByCzLJEuBuL54Jm9Rek11EVmvi25O/1LkVnNsFtH
3rO5bZRRHRR4vhBZ8AGCrqrjwGiGMKYhObgjg+spK/39indsP503ax1QxC3cKN+m
moJU8KoKD6RKFxyqBFrSgZWaK+5LGGDuj8kQtH1fcqg/9GiTeRXh84ZWZY/Tq/3p
y3qRaqsDFAtvlO4hDTCtuty61ut/YkjouaA0VsRhGwAApVRiXx0pbJCV+RvMi/WV
1nmtVlMVsAdgXStoZbxctSTMgbA0Fo5f1T8nSnx3jXc=
`protect END_PROTECTED
