`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7jmXOY0FXHWk5ykW6wZotYtH283i3fzKfOJCi0JSdobPgTWJqQZ7w2NP82cBaN9x
7tGEBRl3s7oLb4SZ1B8CD6wCmfUzH/eCQ6tQETjhEgCOGnUYwgs8Ve3pA4pPbDD0
rvOuqRzVnQ31H1h+zyPvTFbzUtNZlEP2OM/e4Vgh5xi6pIlfv3Il5qmsUVKmcsEb
XKiK6uMwUAGWBuDCPxkVlWHzaXtuW8falOou5yzC73sO0BQJVGcMqJSf6TKN750n
tj0yb12Vfhh3P8ZL/R5lKDXmGluyr+IBcb4IhqfWW8IPsApkaCcRHaYCDkekpMFw
2QuVwpbmpW9xYdHRhrTUSJXfOa15lGjgvlJWQQnblvOKmo6w+BBorK7XSj0Tcv6S
`protect END_PROTECTED
