`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x9WZvjX+AgWyjIZnSsOqMqXB4X1yb0Xmy4fq+boLAZo13cizFx/hzuCLYLSx2tru
L5CMQ0mSfoa7nDlPjH6qFFk/6bLI+C0MasbIf+4A5qEROvQINsEEiYkTs9h7JfZq
JQVDMcnx9dJsUTjSUV66jDk3zo9hrRYncNLenGQn/+6f+vtJQhlIBNaE9DVZogXv
JhTHanPlKyP4rQDJxgpOLR8LWHI0gkIRCYULV2Z+uGkjVh3NwTFtcSu+tAE+iQQT
Z284zq+fkSehaFJHGiy4FlS5lA+sXoLmzbw+5MqHuU5x5Fh01/Vkr5k7V8xtNSpE
KTWTjFuMq5onOxlbcuHrPFOes/mO0xgENk2ckEJFy//4YeKFYGmXHfetIZox4jTN
pd+bqbdS2OJYiCF0TKGIFWH5j5EjyZiwdGMwV4vRbbOvPBlUtbNQvKbxxU3yaX05
`protect END_PROTECTED
