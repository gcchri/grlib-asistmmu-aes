`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eZyvdMJlcHCHzCCn0Qcd/aeTu9MgtJTIUiNekcBMahgPcMuzbt49OOapO3Jzcw4D
rYQxvTJqC1kXR6YhbCHiiL0qN2L0OY0c8x1VOuRvbik9yU1l8sNITCVst2EKsITq
/Vf5CLG5SgdSLr1ihfwibxDeMu3gZa3I4LjFx/oEePJDyI5S66p6XOIwzq/QfKzr
dAMEyQobDPhuWvzOYsZl8UZjdKBdIOUqaoqfazRXnM2pLM92xwqrmYfi/vC6I+dW
0hyqwUvP1SnPIzMrqpw+7uSLLYls17nt0ZOMjcn0ZfUETCg1keUN6Pory29N6G5P
1Q+gEbgCMAgiWvYYl+W8IURZrO2wIIJii5zYU4oAFIW0OFa4h7AFX+5E0Atpu2hY
h+klUcquFXxSXLfq98Qx0F6Uw5uoNmV5A7X9IXd4zU0zEYcs/cbvLgdOU0pBAZRL
s+FTtYaWnsPMni2+yTBoh8JfjIgMQ8Uhxf0ozwXUUF8GctLUq3zprHw8/VGPs/ia
aKKbDcLTFqXxNTuDYHYjmp9L2pWuRpOrT+T50mLIut0q3owiQdTGDMVCzQevmDMN
dn7+APxsOefhXSmN5mMXHf4azLqOCaUHM3rQWRcQ5Q4QClWlmQ8DCuuHSnDR0g7R
whWtp/Co0VJyYsF2lfEBHg==
`protect END_PROTECTED
