`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lQ4PItgUzJsBWJLHAkK8YvRhhWspk/zqIeEf8GmsU0m5NHI/FbefCxeLtf3C3co+
fWlfDj/kmxiWiTKWGOTA+ID2BLyA5Q6vOq/ySgMJfPOZbPJQhPwOBE42mUQ4UUK6
qIgXl69SyQSfv0LBG7vxv4hUw7XdE9zleF9H6f5Kwr0VSMAANXDq2K4gy85PFcnZ
E+0if6tkjikA2vnxMxozYkIIukaUwzxAS0yinYffg3jQfaNf0vegRZCsmdgZZJ4Y
WsddNUTKXpAboO7UWua7Y4o1wdhivYg5qLAR22PKfd8PrKiZoYiNDm0UGTwEouu5
cymSfXIqziNCOenfphd4f1C6bLqw5m+dRwTwXtct3x+Oo4ROs7HHnUzTwZTpaMrG
`protect END_PROTECTED
