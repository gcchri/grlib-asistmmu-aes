`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GEgfniYf7x1AIRjTv2PtPb4dZffr6JJKqnc/O7m4o+liCdyLzlV2akl1Qsxdm2TH
VF3J8JeHBJQEV3aySuo72v5BBmBlTrLXQWazJq0tjAZJOdFY2x2b0YyMVoRxsonS
37ezc7o4e8tiL3+id5Ylmk/i8MS0wJKaYoLd7F0uDJCbwZ7VP8Zm9M/xG0brgaWx
7ebgtHPhUV0JkGRQErv1nlsfihGjvqN1gmI2QNW4OcGEfqoRydej6cep+7Ed8NUj
/66OcNBkEh/h2iYbRFeWhBdD34v2TQ44MfUpfCw8QEV/W3wQQ+RxB9on7Gg2Npov
EnvM41eFREozlP5GIFddRagbylq3iGxesRaE4Q3YWAu05kXgHpgGaHXLtnFLhz7P
w5r4KHbfF5evYdv8Qv0SU+hBhTboPMsLt+I3PXFOHVsynCkBMPd+Z+2qaK/9Bd0p
SclKbUPsGfgr1uPPq2r27oDQcMskIIqptvK3Sl+SpJ1vLOnlojY77D+z06tjP5vw
`protect END_PROTECTED
