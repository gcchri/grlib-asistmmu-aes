`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M3UWsKjYaTBJpALZL+B7xrcYfxHr7+1br7N42n6J+rVLgSYD0vlEbY9txBHIh1QJ
+EMzwf8zN8Ls/X84l0Pq5tsUwDDqqbPBYlqpebfsAgOZkhl1zbJVaj3o8QQDhGgl
5mmrCl+J4DpzNMfofWKvZfG11dzY70QMBKX25ghPE47rDlHr7oNh9MhgetsTp/dX
ibYc2meDY1q1p2Tyf6xngPm+g9EChQZAXmjAErteqkE6krLnLyFXeCQGaxAS3rcB
1YmFcHe3ZC/zB74tIXJ06cSiwzVb/H1ww3Fw+PCNxq5ET78HrueetLJWSF8rFC+T
`protect END_PROTECTED
