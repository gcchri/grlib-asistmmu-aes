`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
68Xzn8Wjm4J9+lwYuY4/UrviDQZdIMfwrzaLZqZ6ZcYcQyBcSby8XG68sYTyGUx0
VjAMNQCIHjRTdC4SBYCiK0KPiobB27ZOo2YGqQMtxUJiW6dqLHAqjwwPvDdDKmaT
R5qU7Xk/P8XIw3P5PGzlPlXZm4dJFil2QQ3askaHdHNRdB8luhWBUl/0w5OH/MGz
YY9R6lr3nxOpl34d3QKOmd+TWlxu9Aa8NQbgTjt7lAO4tiBjdynEzYrrDbqqPZpE
yfxRP3RjC2+JJO2wb9BMlO1DrZty8CUNZWsHJHWL9mw6aAa6tRSat6i1MP06Fcyc
7yDXlTuxySpfns8RvWRbfur6tJRHOX+kKTSSxltPI2lL633GGCIvnPpl4Cb2mNK7
5xxtJc2+0r4M+YxiortXTQj/rob3zoJKBJzohoQ4V0GQbykLXeFeuZKGmNT6flNr
66Ll7XTTHHSrma7naX1+/VBE0dbQzhdzPwNr1sq2nE4=
`protect END_PROTECTED
