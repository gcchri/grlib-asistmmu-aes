`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
udORIhgZxVySU5hlm6SsiTHWcmn9SMUq2/EpHwcJPS5quCDgh91fc+PmBzozRld6
0nb40/LjYAWkHL9aS2Nq1dCZIycnXNf642go8IOxis3zu/YAefe4tnIc3dnOi99p
82fl8t9UIpde/ATHtM4rIyIJqAeH9ADPikMnNaFocFxkDWjP63B3GBohvXIv6UgF
/639sVazL1CzGLUR+mPShPqYT3h0QjmHRaVZvJ2+nUN/j7pLzgzED1ah1atyf/FC
QvTe5Tng5/2xO7tg8EAXe9qE+CSZlrZd57ezuOKAaRe8Q/A5MZKXjMrow+AviTKO
6pVD2Np/hWqeUdzwm6HV6Cfa0ahdL0xyxViH0KbVJFxWNV+97Ad3YeLM9CThEbG7
I12NDzaPMcHVOmnasB5/6kIozvq7ftuOzSxoSi8i4S9BIY0W6Lzf+oGFAuB4HbqO
`protect END_PROTECTED
