`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eUO539g/fap3z4DSH2SQhUi+wf2PadrsQj48jWC8Z9PjPcDeHWQ+ynL/mqLx3TeD
ryWCaifgXWXORwNeMDgwimtdqm5NwsJhnc8j4NPI23CwOY9YK/JmTxR09VuRF48l
DUEJ1CORtZQA9m7q/gMjQjCOXbVDKWEQWZpkje3Kn5ZaQDquPzO3VLvvG72F0LRT
rAknlKbWX/B/nWJMU2sbHhD3Lw+7E3AR1FfJiBkMJKb3YBv+UcBoe9rE6AGmVPdH
B6tLxV3wHxsj3CijbP7qNV33q7ipiQft16/lymbbvytoECQNBTtEWiiunmqIP7eE
xPJiaw7VqlT3ypA7jqp00st0ZyVLskeNkbpkGtFH2mL6wvTD72CJoVsX8CoGguDz
hRIeYBcLimrjbCXD0B4ZGC2H0cIAB4FJ9f4mHBmHTOn4GfGt+xopKIyo+toUrf8N
cvJrzZapX+Egrj6noczJ/A==
`protect END_PROTECTED
