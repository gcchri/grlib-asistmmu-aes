`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WtsaYvVYYI7QiME6BPJfMniCosKxTMne9mbE6rlwMMdJ3F8vsKWZDUDs2AmYJXLZ
++1Fy8X777AyjZI1cxGgCxYg9klUYm9x0Phu3mcYTdD+dtL1FKO0ExN5/BoxwXVP
0XqipOPo61sVMBcozj+/4f2ACLQBvNAtwvSjeV6aY3qAHGu8AS6RvHRlzIyMy7b2
ZbK2Uh8ANMpe0GtEVrlVwVrusBi7ajimaYVwHJu/MGxjoHhRheUTBjbdin2NTwii
l70Ku1W6TZLrem5QJhEgir84605kyRRVhB1QiRrEgKwAAO2135+LN8UijlYtkr9G
jehO9zp0aiaJEqY4Hzz8iqK0iFgH2lPgL9ES1lXdhLLWGjv6gYLWC4n6NND7hbey
jivepUb/jo8zUdubn6nSxGaUIAwrbOW8Uxul97j11hOcQ84rAs17EGLZ/ZF+w2iO
`protect END_PROTECTED
