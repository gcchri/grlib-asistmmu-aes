`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iN3YeoYzC81NHcAcLEVgXxwT5ik84D801bhkCVEBm519AJ5sj5Cdnum8x7J4deCu
JU142/M+qh4u6tfUOwyf61tiAQe10yRMU6h8sCISUEE3+ATdXzPpufDPTbOvUP0r
GkMc6vhGxfL7lhCy7ADJwkAKzUz12nDujghEdIKnZpHbrz0561+GZ47C9hW1CcNE
Iec6HsyNyPVzMN7aP8H/M2gZP3p2bZkzUKEPE1szilVhkCzuPIRJc4lvduvQHtQz
0aT11fLP8sv9XvoxjYTwOUaqwdqrayLfUZPidv5Ed7uNOH4rOex7UDDTWm9hgVC1
jLOaFLJWo4g7cFra17YEEXJBczcvzzmTWszu9JbTuj3mO3sx1i3RXy6bHcenK+Mc
fPglTDLbAJ3rcqT/eFMFpeRLjeR9bpczqwzDbNHvWTC8VAu8OD5/d46+fEc3EXPK
F06TVnlpL2jNR1Kn1x+fxL6Vbv0GOIjzIDCBBGGYBgAPJ2vnuqQvuDWn8uO5lH6O
QUDzSXB65bYkHoB4rCXeOcOW3RjeernCmg3hS3g2QEvO5DFapk00HCyafDT/0597
P/NYaXo8uOJY0hT5JrwxHiHgfXHRFB7Kzspmb/TrsJH9w86+hShRay6WEh8TMtBs
bUuLtS54/bHz7eIKaUu2kWF6IdRV2zvQGqAZnJO/ZTPDN/hUk/yfKSqA01xd7aps
hVjqkU57O6xRKezv5in9tvp7gkFjZGp0R3+VVCImVgE4IJ8shVia55bXY3TyYo4P
XTen9mt7lF38aK9aF8/rvA==
`protect END_PROTECTED
