`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cXKubm4+1N3AafNY65Ws1pGPqD3JpBXr6xeqj8MbtglqP0qnu88lNbTl0hG1JZyg
bkCRvu69QsoGKytauj+VtUZgdH5A2oiG7n1SnKX/7NkneJ7cldhdvnSofW/UTQ/p
dUbgNuAvlAwA8uUfuuRqSE79pf9W1+KrjPX+iPRw5fDzE+yctDz+DYM5kPVFmWmg
Y5m0atQ7TFPQ2ZnfXA2c/p3324yLjAMLcGLZD/ysoPz2t8iPX7HoSI4VKhZkH1d4
xwrSKeaeCw3EHu72IH4xoX9DZHma9zcd8J1w0EHOCdSxzyXSH7jYaJKNg0/GqQL3
8nl7KSuVKUtj2sGexWI868Ap6DZlXzw5ZZVvjZL9m9W91cZh87xVHlpItndfn8Cc
WoPlCrwBgsh5bZVq/dvfcL076BWYeRYVqTyYXXMuyYb2u2/N6QuY5FZJzz2GMHD1
Ky3NeWtrI2wO360FUnDz4BjFp0S1o8Rq/gHduXsncHWYngkrlZmIr+MCer9qnKav
`protect END_PROTECTED
