`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+T5XAbecMpLdwJMgwVkpoR4IoiTzFccYC/fiAXGLeYCfIpmDhWjjWWf63zst1L/L
ZSTXOuUXC6hUnZRhX837BFmhp03n5q8Bp++ehCya3O3pEgLrBLal7DNnfX5V1uXd
Kb1zCfUHUcx6ATHxKNqNCH+80a1qmavwl8L/VDyoTherfUkkoxHfpFxRvPKY+ZRv
LOq76O+DQKWfTUDwurqmCFLlSGrkY/4bVfceDLlBoehq1wQJ8H2EwpwF07dHK23W
oA/XEfs2ht2FRTQUpA4f5r+3bVaeYQ6NTNs2Su1VZEse9pSzsXhqSaYiREg7RnHv
iqw3yUfJeXP4tRW0+pYSv1WPVKZCQw3QIUufRP5fXEAWtCOrP0bMqgQB1m8OS3Ib
nB2ehY+avISsKYi47irMRA==
`protect END_PROTECTED
