`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jg47Fe+4qFZecq0UbJae48c0uiq20nL+zwE6WDMrmP7JYqt49Fge3j25DAnFjzin
tZ0mMlTUFqE6PzPd6AqV6btKX/hYXTzxSiwkEg+SG4JjC8TYt39joMFOcitXPsMT
knw5PIJLKaZKen9bdOQgZy71bDDFuWs7g+A/QrTuKb6qmygS0FjpwnRj1vXCtfYH
/5f2lV8oMdcGiUkkKvoZ+lWwchQOIQewAyow2dEn/G4kDQQTZ2CSJ9NJ8Ctzatvj
dv69igai2Sq0Is/g3VzGgbdPt+UsiibdTDJ9ciCmd5GeF0kFmbQkLz52iQEh0AKr
qMh0hmcA6OJtmJgJOrGEvP5H6RJ54oC7Fwh5Pg1oezchZDXfuB0mRJInIX3/QzHe
jpLmWJjNOMax0SqkF2Yb1s+DYFR9SEdnVnLSedLsjo4=
`protect END_PROTECTED
