`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UZqUPGPg/SiJ9zEU3uEASCi9rrMnzR2U9CI+U0kr9opnNja01DN9L22Z+9q9csTG
p8/7qIjWsL8/BM+YxIdFrDrSfrcxq/xzGhcWuJGKX89PJ9BOiaiIFvnKSJd5Eqh2
CusNrvd/1uXJQpQR0SHRYaAPa87ALVjphaFuF8ZAlcjGZrxtr4mtHCTYKA23n4pL
nIZ3Nybry+X8V3m4x8+xCCMynGDtBndBqCYd/KhelxOCu/eASXt2j8KmWO7BZNQ3
7OUjXHKRm5OcurOoOZtqeR6BTFzmaE4/yy34fckBbq/1OZ+O7AMSEusmdKLpWNl7
U2lNBIQi20M5ZsI5ucj5Kaso4ZIsb+09daVib0BXmPCXF3Df3LpCOG440pu9lMPd
2SN6pRuaSwlWPSQq1YOsuhjpNk5jaW57soC5+3ojjTNchJspTtgVHnnDWqEw0pOZ
gee41sXwdzg7Lm4ghAEOJJ7esgnxIkBP79lQtA9Rm5syFubZfzGJlNudBBCPc0Sn
MYNPmOWp8Mv/Rj7Q+mPsJ82HC3VUZvkZflQLFUTD4N2QgzjCj/9XzvMJQI+xxIsG
5SSuXH8BNCwuuIl62VOrFAg6t2q6TUZaxswZaKYdwKph5hoZ+hhgAWk6N3HDJswP
TQfXhtXQTd9qlp0ZLr+BVgGLZRVt5uVj/6yoLcCelLTYSRXToItOX935U+L54cR+
HFtfX/IZqQW8oYqJqE49xzA3mxfPnrkZewDWSUO4ojRSQ3UGt+0uHCxF3LmORm36
plTHG615734iADc+VfaO8phT/OsNs20tVstMWKB6wQanU8sIJCugk7P7ydLDJoUc
Oot/EzFIqRSPKx2CxI1otS/OitLAH8mvzfD1Rcotqt6+1ItiOiUhb1Hto/RA2tbK
jP7TXk6AFkSgO90Ti0LLAgzKw0tbmxzJe+8RBMPMQy2Mwtw2DIRFHnTCtclVoC2J
q28h3TOQPG/sFBd+jnJDX8YGVn7cZsaYKSoAEJWZSRFfDIHwzlQpzwV34IoCkVj4
+8jaarzyE3VHNd/K865nLdytBEm5aqY8uxCi/lM8dSxgLoAI+NbNsbrHmEE8/xtb
LjyOgrHD3TMT3JIaay7QdkXlwgqUeArGApWWIU2UXK27iqwadRwui/wuB8vmovj1
nEhV1TL2sdiXndsKkaIkrREN09bFxrg2HVH4lbGU1DheNp6NGQrRW4CjZCW8DczP
r3Wbj47fywF1SdgSfRDnUZiY/dfxcVQV/h+nsUtMGliXEHGevTO9DUDlcBk/tUsc
dtff3OsEQ2Q2jx1myE+UjO4annCwQfPYKtnlmQPTVP3ayCXg9feNUH+IMHG6wGuw
bx3QGMLO1Am9AqKqTWUQOmdJ+fZSC+7OrEPlA6/htlZsx2BKt2g9YQqdJ26N4sGB
LmA1OJPEHSsA42nJagh5V+VQ8t4PDirlOw3O6doudkCzOKlTWI8Nrshf1Rspc7c8
`protect END_PROTECTED
