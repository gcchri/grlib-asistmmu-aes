`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OgyGUediFWihdb+IqV2ZiT0JOwvx4xRuIcMhs0xO4r0594F1zZLdKPHp56wgTpS6
KEitpE19zqKEIeg9LnACszOpdG2VW7YxY0LBbDASskDWymvSYXXyz5cOFQj2r/fe
LllLlZtkp4xc653ewQ71Esr13kvHo5iVPV91e7sOOJQxRCftFBz07m+vattgfiIC
06neq4lTz69romyJ/A74hPOd8rEVEwxTb574UJ525D+UDT/M2Q+ynG0JER8T+oCN
BBUHN90lYXH8SeZv69/OTY+aZPsW7JUEMD7G3Lv+5vVkysO/4V4Y5DN6R0gnGO48
E0zDWdNOuiCEa5F0SFiyNzMsPh30+m29hLKExveh3OczI8JGrAJJz3a4S/7mybml
OX2fcxfr6ZWmE2yE8H7n1ZKDxhzEYvCYUALMVlgyHnk+ASeEjFoZENVF3p8SqXsS
dD81hUjlvXTZwB5nNafM2/OrXLI/rlC4J03PAeeUF2D6r2LY7/hfZyZ/DwQi6w60
8bP873gHpUukJ+hH18FmMZo6Yjo/On4NiUyCQ3nIgEm3+qsXZR/uQ+wBGIJbmviC
JhQ95ep5UAax8qkUzJ0pD5qwQ9AzmDIYYb/5xHmWhqx1Tj4cEdP6aBCf7JSQd+Iv
P0HHA3hqy8giWlH80KtZRH+WmqP33/1g7uLZvJGkQWA=
`protect END_PROTECTED
