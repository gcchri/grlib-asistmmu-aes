`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nsNMCe0Q5Tb1ximo6Lc+njFWMEqpR7dmCIXq2lOhF3M5tO8QtLxebkf20pXbyQlT
+6QIhl6qDjAS8uND3jJelUxceFef0l1qM8Z2Zmeb0nKu6Ean6Etk8Ni6X2B3rKSY
7U37zoUSJVu4T5BIZ9BbBg2pjJx537OOWf9T+KgoQq1ijNjRmDMW1Dox143pEAN8
rmtGQHRdGDijgscRwKUqhcK0PxMus0KMrr6L2bzq3GFCEF+Tgj/o/N9EIdCy4nIw
uxL1IzgR3xzjRgJtvH+vckwSpuci6EjIsxtC5+hsds0khN5mYEnjtqoGZhQ6AvjL
u5rKLs80yhHg5OMMWVLmsp7ScRGAEiHSseJ+L0I72K+2m1wQe3EnXVJXXR25+vQz
QhP35Cy46zNK+2BcKozMIwVskyfPGzMwaT2hY009plXBPgrdknQeiJWM/qHeevAS
FXI6Eiyr38yv71uTt+SbhK7d19eDxhXPuf1xZKnsNYeuHA9Kf4LTyziET0qwfuoy
YqWmu6gCHrdR3FlCS+0vO0CnQ/aXLFIbzG2ORrxU8W4OEddSwMESZ7PlCnPJoi21
s3Q5EzJsUDMPvyd+5EWmHS8MqATKsjlX8Lojafd9vlvJJH3204Ijz9jC4sBP+gRE
S2cigP3HOsqoR/OaqV6PWdtMW3Pb7Gr6EV6tmVh80wkhgYcetyd7dEs96+q0CnSj
qDnZayC2msKmNVK7zW5iSd5272B32zmcEzelan/kSm+74PBnqSLqbUOOrEsO6VdB
l91styy8rz3KIoepq79SpXiyee3xvwtOqiXCiSgYTlX9oqmuxPotmYS9DGSze1YX
tcJafe1bHxZmc2gMmD1ryvwgaFqvSsn7vaSTaJIiuA6nCswpF/HF8v5nt4YPHHqk
1fzwLJfhRmgGWzpzZ0wAHE+sE3G+jGZMHDKbkFNvECXDKe/Dv3IGGAoU3ItaUwKN
3h7JOplNh78TZHqq+EUUmiY0HgWmqmEdqjR5TvexlIfd99tv1RqcnUHbUHkdIESw
S3t3mAjb4AauqbwCPWlGAOfLcnJOZnt5Spkb1sny24CD3RTpYEu2YUnche5OnHbT
Oi30DWBzD7AeRiumoiz6z5rTE/7MEyhqnl1qmuKX/kzICDN8fSlncQbRPBjRHu9z
a6YAG+VFITO0mfUvMYN8JimPqgcYzzMvp3o1saG9ukpl9Ks2O34BDpy0MA+F7ybF
sjsp4vL6Q9hblgGgCGDk8RgsFxkruXUMCjo4SmshNRVIrUBpDDi29NSLoCPi+VEv
AuwH064sqjMinnT21mFYpVHQo7yp9/AiMIhdfaRVF3S7J6Ov52gwBAl+LKQ1luqb
Z12NM5xjj+8GweWMMZmOvsBliQF7/JdXndsQqmtPJaH9VUubu5TvAyogtHj0P4q9
DtDa1znGR3zMUm+BKgEWcqa1I+KnVbyooSJUBxik/0KLtAOHIwgFOgA8/Ajyh7YU
rPAlItMQt7TgG0d8U1Nr0Plo3McXjoTCahVpWHz5MOf/9hgD3UCfn7dhkKJr2ozo
hPdCQDTXhHE48TcSGkBrQeKDcDrUiakVPkuPw17Sbyu+vu1pYaI3rBIdW7mQNpTk
9fK/5sxqvVxa0EGa/cCVUhwGDemnXGIpD9oyE2KLd02YQC91YmkD4xTcuUqLY2S2
cbyjlugNQ9IC/onun6T2b9UWup8Qv5DJsiQlOE43zr2y2L6o+sK1vNp3EZD/Jo5j
FidejTNAvFI8l+ICo9MK7Lgd9TgHt9LXB5+Cp06eTi1ngl5mXB9MvJsvBpdc3Nnk
tSntneWCWazYdwSmaxJvFhylOl5P+c6go6b/iejQ5bsx+m+qqVnbOlPobOmbNaw9
XArbEqObHOKiyeWLaw/5xK8vnUa4G/d3LorIl5JYhmohDFsWK1GMZOHKifImTTE7
OT8pXBtglwEyGwsAOAHLCyz8iqF5ZOJb5gJtbxnY7hyzh0fN86Y1o3+PCFcMElah
9lgZKQBX3KGxbBe7cmT3tsW1KL9F+f+yJQNCGh9ynjPnwdZf1GeO32DzPlSQP634
W2JKtUaDoMi3nGjaxz1nJZF+Hu7p7ctIqpPvtibaS9LsqKuyNXfhm3cgC6NpVpNP
sP76k/t/VBkOmkF68Do2ZZ5zfoDoM/ds3N/+maJ4Ppl+WQiKGu4SiZzA8FmLLKio
BVnkHMtbIjk9/KkwCxqeLST2OOHlvcHNzJGyFsqMLRTzbmHl0Ad4MBqG0G/9drpi
G+uaKtfIP0Sp4tXqv6FUAwLsj/PX6meDZl4shryB/K1BzzflD0Na9uk8p6Lofb5P
OLumziporrIp7vXI5Yoaa+G13Y+GyPf4YUtmnRC2QoOJ0J14FWZ7DToPSXsPmL8i
UG3J+G+F3csLXFE9d7U34NoD/rsF0ZR8zFEp2ApuW0Y2wdqzjZbIvbpYJjDSdDmw
LN7CmfohIWBl/fbw3FlLQaOwKWbqv+VUzL1IrCQ3hILraXuXhLQbAVFKzVbOyPrp
JDmne8YkOEXUoV8J+RCqZLVq8RLRrtZxlX/A9w5JlZVSuo5CLqst0KtOS/b5r5gb
I3WSQ3k6OGFlUUWWQUB5y+zzuK450iDfxlw65XvqZoB+lCw+y+W43WzERlBGKX8u
SfSclNfcsXxb23I7SAIGsXPuKLVGjGK99KM8/H7x7aFSML7YftogjF0+QIGcwsR1
t2noUksvT/JfsYnOH8KbHZE1Q5+jDPBOHfOkQqF7dSKp1pdZwuroS9CzEl6HODvt
88US/7PSbvhFfmxMkuR6+kKDk+ZNL3E6VsRMvBEGfl72o75eOtaYZ7qICSuVM/yS
+byQGCKdydOLkaOd/kp1U5t3o3N4ayxqchs7umwr4QWqp1vVXCm+Q5Qs7+7GTXQ/
mOLgljQMuKqs6s15KrdswMmfk25loLmW5lDYQWObaOyOwQq42oP9AzvmJP0sRy8N
o8OPUk6o3h4gTE3JVfQY/sGE3PSPeuh3qKIux2GWIY7pfr0Ics8go1Q4+Eaz01wy
1yhRSKrER7217ufRn6w2yeN9kGYLqpnKKUmVe/7J8ZlGfFjeajnJ0OZSp9+MeOTh
endp3hFCzA6v0C1GeCPj8nFZ2PKojAbOozDeHZw6H9sDm46fWXLu1GXwDAoPmTev
JtSqpxhbY1y0bTBROvn+sSS9l2Ey+BNHb0oNanrrmmMjO8vnHMOXqPw8r92IDIOW
BZP6EzKlUD37CEcpzMA49OungKv0CXs5DU5AMpfdC/O4JHuCrfHSHL1Hv4ICkRy/
i9Sxf7rmKW0oZpR9ppPNPwGTjwdUlhZVm9CdNo+P8gZ4x/T/KA00vHkvSIzSIgTg
qcNZyYLfAZ/iX985gqdcXwiMHgoGE8e1Na4ZB7Mzf6643DWzvs/MsY1LeJIO9y8S
/i4ssGEAAOatAdCoyMVoIrg1O+6U415fXDj7zbuCP2btJagflfUV1X7pzPaMU/uq
+z6mzF9kmO21PiN5Dk8oGSiGLEsyO0oL3KfOCM6S2Yf6hwqClsN+oq8KM8BKJ/Rl
P+fZYePUVjPEcky3t4+im8Qy+zgxpRdq8Mjc5B3svITg1hLpUgfrmlqljChWLR6a
cO/xXEuJGWv4YAi56jCDhZukL7FgUFdwoqBOYQkmGDRmZw3wN4BR2clRrgA4vO/u
yQuVOYCLXc7Tu1VT2EOV7pNWD8upcmBDVW+LI1SaJBaKCna5yZF3tVVFVZ1qGy+X
bTcCslLg3ZLBqwi3M6zWWs1rV8zvwjU9OcZHZkKgxiZ7ny7oj0QANkXiJG6ov0LM
nRcyj3ixzMsQ0zITEiACEp9dKC7suYumlP1fQqszc1beAvD4iUMfvodPx2qjOslo
0/xhA+N/CaAbBANyxkN909aDwi6Rhu2xieMH+vBVqDGLY+eUsnAs5QFoRF8tOuoa
DbCuJCDjY+sU9gmOF/J+RQNH1+rwmh/R+q4BXg07wizOqPv834qvZGIDXJ+fxAzR
pNV2mFUtgYfI1ApM+KTmQfFYfjTkl0Rj4B/SK3uZYf1CBLBPVdkBmMGKuYsF/eVa
3Bl1Jt1Oa9xC9f436uPsrsTx7xM4RChUQzY3GYFI7lb4C8F3eEJQ0IfA7DwHCqPm
8EQ7YpEnVy7rCopLJaXJzb9RXNmWznd7mY3GCrYh0+lcsKLwdAdK+tfRvyEkQXrX
4Y/HekRn8T8OAxtT0GQyBNpf6SKJRuYvXTL+yhgFNu4EB93r3VWPlZ9Y6kMTOLy3
NGbXGU62I47+4xTg1ZDJuLlzmG2Opkp6ojFr28Y4FYkaw1fNV5zQKBHWHZ4QPAuf
0r56FvN2CKxSAqzSKIEdMh6EGnvqOVN6VO/SgtjJXv1KwXHOeT3p53SjmeRquKBU
IFM2XXxm9GfXdLVRZbpmzS6ddiHYnUKijWb3APtSUv1quymFXuX4pNbH8a5jf6gX
yTmBkfYmX7xzPVfyun/VaJyrvdMMn94U0TsZuMTTnntK9AMa9zJs0U0zHJR906Wk
mqDg+DwZAXCeLbhYmyy06WbwHmKMAQRR7Egn3Za8a4+F3cq2/2/YUoyaWZ3UCELZ
X9mJDXUEoSl4ltz1VKN7Yhgkev57SdTQXPu83IrCZR82YIyXaUP/OHt2H6COUZ9j
eVUFNNOSafpmhnQ7Rql13YGG1tRKBnwfjvd0CKAAEnO9qR3ChPE+jG1DqO/DVHN9
Z7rM+GifV8dr5VEKwpjR4zBTJ/Ke3i15zZKPuN6ZpIFDp70HT0/TRJmY4rGJZjX4
nioNR/9TeFG/KHSMR4j6PvALOM4CDdiU1pa6tBWtAfUdQcAolc2VJRHIHkLa8vlN
EPwdfx+UHRGmXfXLTz4O7bkZyv+NErHOWDDYAXvFPo/P2beElEzR+JT4DTge0Fym
GVr+ZfyzBMEGAkIpuW/KMUbvZmj9FnoOVZrjkFaCTH+77izXwqfkPfT04Q8DLlmi
ws0dwXKoENj51WAH5XncohrSFpjC2g4saFm/bSNfzILNPmPpbSiWq+f7vcE2w+Ov
5V3pJM4G9qYyEqo6ofssKeNMpn8jbtE9HLoJcCc5ey6WO5BlGEC/tuIFSTEr1QtL
7J9RDCw90q6liWp/VXh0wqfchvyU8Pmorc23/Splcem6pf9w/AC9+oP8izHYuJpY
D85I8LJ/bCwStqE4OFcn0nWrlBUFVs925kKH4M75aKfy4wTfkXDwLZXLYChvuqaN
DniBGbWDrnEFIBimhlhCiutRqRXLRbMASe3h1P9iDyQQuLFN9A7NEUI7AuvlkQwE
OJiyE+aSk+yRtg2xrjrf8hz+CYOO2Jq88qU/XrmgrvfRguuPHPe1H55O34cKuh3O
MKbGD5+ZtJ+BQuG3DTge6kxiHJ70ZMDKmnuqyb4zD4yel43hDfvvwu/F2hFNyZr+
9xuuyIaKuva6UqjH0lfBTPlpG/8jR8wqwASIQG35qNxXJgySdxSg/8xSmEBio4U1
RIb8LcfQo1tGeBZtE3L/aGhcP5tkLC5Nm79Cq30zCHIFKBUwNcTfdkrKSnLGaVV+
lDSL7hX+b1nu9M8rDhbAILWIoWQqZZpARkqopl6pGIJV60NDnWG9os1aCe48Hj2j
9jWme22bncuqQ/jDU240cLeWmUfTVT27lt8tGcKohWiEtAWBxkfuxFysd7Rltk54
iNjeYDeLm2J+CL9vPIjvbHkf8GjQB1dEoH0gAmI6Zu5+eW0D1cBx3Qg+AfrKoZZb
PQz+p7ve4w2c2oE7Dwjl47MNbTO2KjBTdToPozHxIL00oPDz5cAndtTDcOo1O1x4
fJzc12TYYDiP/NBhLbcniBMzRGUwIJHo5rym2qP4E5x8f953LXoYI3F7CdsJoZqc
gGkN7Bn4L9nI+aK+4JL2ZXEIURDBdVGkDFED1moauwjhTZW1Kjy1WUbiAIIGHwMO
T9+1rjw3W8tOYaNRwJzv2SFbPVhVoo9fir+2pk/r4Gl8f+bIdpNszoUqielG8fHC
xrvZ3hbIDEg4LWLaS96gM9mj/Gr8amtyBnwar6VjtbcaHslImt17jyBYlcQukmTE
ecZn6cPQ42goIEObMJc78NrItyMAmjQjpiL+F2CXQSaa7Lhs/CpV65q+ulfR7DGR
+8hsjRrPkD3vQE8BJyIW1T5+LB2T9qQnYaOgN7hOzTKH9zgfGlHiYHZwC7iJyJIQ
v2YUAf9FpIoqNv0F7Xu3+EcfWleZXELpfAOUkwnakLL5B1AsjIIJdke4o3JrgSqc
3VlcBaBpiqGHnBh0jo8XWv/A2PBOc6uDF382MRM+WvRijY9IipIwhDZnSWvOghYS
G03rrxIKGe/00PPvoMTbwXdMhxSxy01nzzEXc2sQ+agE5QQ1uVI2kaga7F+1kauf
upFHKACPmwI80A2yXG9JDdzvJ3VlsB+AHIP0czst5YbOlrYvA7hu+Ha24OEp3YGQ
1Z2EsnoYLYGgcfZ0GBSiKrA5+dHIA7h73iUqhTJHYmLUMLc7R7Mu2e1y1x6aNXeR
fNUrlcx+v+COjk+Qvx7IzNylwZgs+1HQzhekJutlznQ1Oq/2pxyeu0aUDlTnOiNI
oJz9pTKlRRQ/9OK7NZRrEfhm5xWEQZ0ddJ4G7BD2Vv2mJji4S7RPf/yipQFhWHx0
UyEoEjaDkV96NEDwfgBGIPSxSLEtgP0dNuFpm/ldEZHD6SU2yiFC9afebqYl6ePQ
IzNuN4SNWgT7Zf4K6zQIJsy/bLpT2ektkNTxsUsphG5Da8/oG+9TsE6k03mwUuZp
MzH8JPNs25F0KYgQKz9hgfBDr0diLRS9t4/axLIK+8blU1aOkzw5HsAqPFJiPgx2
mUUFy9by8qN062WUQ87XPr4sH1zRAH+9jbhDMzWUn8YapTPNdmygleK3dmY7MIy8
7pxZqZU7EjdSFmJJaYJE4i+UH2NUwhWqdpaHbvKDHNcLpHgPKFTisL0vNwM1WDgq
eUSJQvn34C6upNUmhr6Pnnz6emOBXEaiZl7/tR2/8OPtzusvDGS8t9Olab66Xn10
7W2KFDX1h6rfZJGi0uoXnSDeKs3V3ryvslET4O7bQ4SUWKTWnkdmZn+PMF7dYW/7
S6hyaoeMHR/6PGA3gGzEyX0z32Svr+r1bQwu3t4lI3hdVI9uqKvfxN76D8Wijpr2
YLlySk53gm9KEdK9rWb9bHUBuHqvNU9l55cjh/MdZOZ8orH/sX5Ox1C4hKwpKEK2
U+/1xbKsXNXTiMxIOJCuBLEqVqKtzyZDmKStJjG7EYhuUaJCfJuIpOMEKHjPie2P
H1tdtr2jHevP+Oy7ClOlIYsy0zK5NcsEbbVltRf2JLgVa4RHyJwGYYJq2dBGGXjd
iDqO9pE7lneC0RdNAl06r2VKktzD3BrP4HYHP+oPF3in0Sds6dgUJRoiZ7yEtrrm
jNIYji5XKW4OxfihVqjsyr+erY6asYSd1xXo5ss+lW4iilnb56goLWy2CZn+frss
e33y+nS5dHqekWENH9c2FB9VuGWYLA8RicJ66L6+K9r/cyad5OOHlDvGcp5q+jyS
fXwcCsN6KXasjF4sgifr2A2kFeEbzJ7P+BvIS5//8vNtljIOz7WztevfwMzj+DNf
5MyHFEhBPwYgPKZhywFc3wlq7TIopJye0dAezYEah6Td/8hguCen9ZEy5AstKilO
47xOvojOkNTE/6HIaY9wMsPDO2fAmQYForhJeWnjG3KLi24dml0D4QL2Mn779B/u
5a7jk7+gKcsYQyv7lz68HkSUJPpljKnYML8w6vkMoM0SUERllDtiDZsTWzm3JQ+R
hj+C6Fv0vxxhILuPH7mdZ1vE+E28wM/q99BRDbSDOCgWVaWsgdvkutm4+0fenba5
J0UoJryFZGiGgqyHgI7D1e2Al4oHZZOct/nEqn1wMpqhGX1o8EwoveIgK0DG/Vuo
MIp5Sv518NPcCzE8Dt8gIVGx1eAZ4hKNSI04AfliA13yD5vtlq0FNRQFKxXBkrO6
hkrMZwkU6ZGU4SzeOBNU2aOws52Q1C56/SM7y4ZV1wIscMDZjIW8t6KAeQHKcMeS
zPt97xfBhmBc1TzHKgh+8YEDZ37i7o+KEM74KR0P9J9NnyrvKFckQaSc92eRccbn
csx4m8m0aP/xFy86hSUjstMhBWbaUopAiY5LWpoKu87UQq77+Cd2RvegWkjNe4Qp
y2OlNUk8zciNu08ch2lBB1cfF+GRjOhRP7ezufbIacmS2QHE5Y95OJu8My5kfA0M
Ij7/v8WK6Z9Rem9GTaXNe2IX28Pg1SMRmnYzJiaug4kcp+CZCd7owmkli1wGdz7+
PRW7BOCqX/8CxXs3toU+2YVkkNqeMrQsirjyedmh8cafHdGjEJWxi+434JIzBJoI
ofh325ugVQB5UBUvWABSXLjPv+oiKpB74RbpPeLg+oAOIiPcmZqRJHTVfUEJqmPk
GkoIOvri8YvjkQj3aDJUi1gFF0EP/uQCMaVUsYuF7xDp7JnCtshgsblLGvAdPK+I
eYMPPYHAtQO/W96zKqRa8oTsOIdIzfXhgIKZh28uy3HCv7Ib4evil3CLHpq2pfgZ
JWFeuuvXORCWVLnEVXOrWYqlXUTh+jfIh9573Qa3Cd9NRAb45J+4a1IL7gUCJWTF
FDiD6NP65NM0hm/jcCFmzPxkt6wEHLZIv7eAOToiQUg6ho49F3CoSz27a8dmM9Bm
H4RXB3oAg9CsHPxogIQe/TFmoUp9mLVc62E7T4d2zEkbbhfV6a9mJ4BBDJKu2qW/
YxHYbSKk6VCzPi6TaEeAtWtSaICyQgpk0pcDeAK0JcMhW73HshOUy/YhSWqv32KL
XHwd/gFfRaC4tv5UDG6YNYq1LrQaVXp8dBBlGUIPuc36KdbiT4AYl2nG3E2/GDA3
HUnkBDMFb7w3U2J41cwLCSvYXOZ3LQ2kS9o7HQ9wBYhs7VKifIa6MJyJtxECpIKT
+9Y1R8iNB8mYXMcjdfqO85RbUZEvr2OOZ7Lu58SQilcuM44i7TxnLHB0AHCEpSE6
yOVkilFK/4KrmVT5z9dWotPSRVKmpgDtYfWaLXp1Z7eN94yI+3S1ol44sx1UxYBm
lhGv/BQ1ImEy8ukn9nFVtk5bzwHo4YrN5cwV04y1+o20kUBZzuOdHQUtCQ9tJZhL
eRrgiE9hXixxam8qpK4JyIaCddzb7q0DhYRoqFwkKhZ9xd49rk5KWrrLZNYF13p5
KtqvCgKOt85Wviml3ZdRgQ/o4McUN+MXR1UgR+pJQ5dEeNI2X3TEHh4HaljS5TV3
s838xiD8IknhpCYo15fHru9y2nU4vPU89j2vUEvAeI3efBYTJ5gqo3jcuyeQnfkU
eUfgF6SQTETtZ5cG2oMMxu0py30OHUpPAn/d+642jlNk1DaNWlLTTu0gp7FEMRdp
yx/QLqFdmwseBw72rR+FJ87JZtberlmsbzBvTJDRBhy/dS868DtKleMRF6mTtSrs
s3uUAd83Y9S3QX4EynKsy3NCy8Ty08Y/3Gx42eLPxhmYyok0SIGkhYRagigV1fcS
cvuG584sH82X1yU53vIEtefd8j+34P4crFZz9x5hK/Ndi/WZ4xmbbNXRma1vAkMs
V0fZrZV8YGlf0dsLWG619U3IdbJ+rXmWVCyXJeCo0lKzmzurxMOQG70uFxizH4g8
Ji1tQfzhNNMHrYZTTGeFownYLsWtTk8FUQ6s4/yBYwzMAVsA4Sb+d0mTTfLa1dne
uKh4hAYYMV9SRxxp/zQqOxNYxFxp/iv3KkAoJweiVohgbx3a12HXj0xu2j/WDRcd
mXGuHvfBA3WtHz7N3y37P96Jpi1zgxDoMGsMZq/a19cb9ba+n3yc2nswC2LhXZIY
Ed/9rn897SRHCZyLby82nwYWlEm2vrA/lS+RDdIXAsHxfK87cvr/PnE4UivAkpyx
ZqeVpp/4/qUYjo0Z+RiTsTwBVKAwkt8hRbstdxvjHqePs16miptWyBDD/hefRCHf
bhhBGx3Ts9fNBtnI4JL7Egv08Tidgfwfo9cUzTDMoBUL4treYvuTEG/5YsBypS/c
me73nlDhlDP0UObNrjOWBgbX3s0TfbILX5IdGRBGnpGU3PlghjxUz6YwuqIDSNoi
/VYnV0STAu2Qhg4O50oLN3K2x2ai4L13zzEgwLE++DkmvHlUadVnfLR4TDjLi9zG
HrVYTEiAn8gaQNwrADzk4iot1kPIUFw6CnGP7SeBbH3VuKcROp+SWAGpCWjgYtIP
C6erxeUHlw9iCRg7F8r6j/r9HrBdD1cLLuViW9DR2kIpEHvd0Afz0fQonyeOuPpc
vYF/SQcU48bGLUCyZOnYbPnMvSDhxqn56e/59tUuyBvIbcD3FsxfJwP7N2y7sepA
/blbIF2yu1vajju+4R0XOkkS0zvB7D3qh3SVRCAoXtt9XQvVk69Wg4d4S5Cws0Ep
AXfh5ciukATQa53HJo4X0TE+zq3IktG8QPsWLMxQsrkQAcN2CW6Xa+gAKWpezGoI
gH5hUYzCnXkeiZrtkM6EYEcqtH/Bt4q42CEcKiNy3oi9WtsmWEFza7ut9Fhg9bv7
dDjvxxF9K0Wk25iSx7HFGR18GBk3hU7gBcoP+YMTD9NjjgDJo2kmkDA1HYNgjEPI
clP0c58y+BBB3RpcLHy8+IdqM7ZjhuLuWdXt/is+xkjBFhG3KaMN/qZQAdiE/9LP
O8Hc6JB1y3jiQl4dGmkq1lGXKExtALxx7Toz7zT5dKySXtT9pBj3OlKJc5dLYFbS
OAKVVzbfxrHW9XUDGO3AOC57zyT3MmRBhw4aQXxP4oaaKtf0NBjq+WB7vOKcQcRv
q2o4tmb3RWR7JM8b28XRgoFfxsg/J/Acbtzbr9JDhgkUkbTeahfiIMlvtbY8kz0S
MxU9Pwkcf1wfGZg7sWL2LKr8BHaA/wcjzXNwRpEnILbV38clQaZPxPswJQuwVewY
NV10x5kVETd2XIvcbkQt9RNlb1fyg8Gmqbyf9Bv7i9IIWLcAJNUQPcG8QObN/vgU
qQR5b69EFiSw4EE64PXWzDmKUtENnfRGk5RbTiTH4qxyyBx2kKbkX60IRQg43OVm
q8vUZgCVlCaGlD7o/ANhUcb9fW4w8MocxHwOYUt7bEWzF9Jv48fpYQI+69vMrEnh
BBLodqXs7v60R6ZZqjVeIzRf9AYHv8/veXqxZ1yR76EqpeX/OKvzjyIxD/7Ol28f
IMb1ftFbKsPOqb/GYJVjgmAdP+wcKdBEHBO+9/sQZYkVBQ/MPpvpdUeHYqXaRuiz
ZqeAPT4BCQqqF4iE9rHjFpXwwSYryrXSRfHmKH4BemyedsS5ugDTi4iHNfqyMhfe
KPtfVySLKsrUj7NTCWjFRS+++F2EahdhwqvRywT9Q8fUPuhMgd4WsOBpnNdCJH2e
tk+Lmb21YQE2HI3WXdmO4lqmUqiAIFeSddYuTKgMVrLZ2+ZmPtAwos38Se+Zc5sZ
rJIeVNFXN6YVjEX3e+LcHNOCB/jEfal/FmaSxbTC5S/VytoFwgOwzKfO41/QOPN7
WVErppxJjr/bspnYZnBbGQ2zylPXbqj/UxJVApaZCrb4s/o4uA4Y59V7DXBFQkD6
sfwWbO/CSv27HoKU7br06u7j6lOsrEU0kP7lHSd4RKMi48jHfiB/Xy/WNjuvwctc
Bb6BYCwHsP1LxAx8Rl310IGa7GTrOUduyTfgytmB1Av13WzHa/atMOh2cgcfQSF1
PnV00k6254VFIRgwwkKIe40vnhOM+1NcHmEpywdTsPW5wImsKYnsS46fLXt+CQ0r
DCy1mW1L8/MivpwdQD2SI0Go2Ifp0CuC7bGXhyj8yAvvfe9qvW3lz3A2nHpN18HD
csU+VeMbhJkgMm9ZJlH3rzf9/IN3d6XXLXyxUa9aw5ewfTi8bwwFSoRUJYygYKr+
DJPRx3Qiid6qrNes0R10hLjfWlPLlzSBX/dzpHQHtzfi4Kumrvxcszzy6njtqZ+Q
D8VUNq4V71f6/IxRMFlntpgR28UMRO5Pr8K/JDnM4PadvnujEzhtOoiHi9OFQzGU
qNs0jql/cz54sS7KF65PcgsH4j0n4VJ8pA4fE1/SA+K0sbVbQDO5QuHpCJ8kadkE
XJKJ84vs0KrMPgiRxGreVIN8BCEtm5gBk6OLJY6Wm80SQxn21GbNuY5HtCG2UcYp
pg+7A2Lw2RHQOFXxWbZ631Mlovymg3esdE8wf57jCjWQCDlAZzoe1izwF8G/b3Z3
PMX/D3GwScUVH0iypDk79EuMQKoCzOZvkUkrbbuNdi0jR6dd70z5fmsEX3ldk6Sg
ji1y5flzUmNGF3JormDwoq8uOKBMdY9+480jZHaZ57GGa+7mQgEFnYHHO0o++s35
Mq8uBPF9x/ZvesQ4VzLK9aSEAbA+6FVgl5ye8gGGYhz1o0Vcy9XdRjv18zqZT4zZ
stoG/iX7xJiqXLxgUWlHNPM0yGSoo/Sa113u70YVj/HT5Ryegzb8iOYMtylf7/yg
GnZX9K0bS25PO3fR1crkSuMButuvPm0cdJUTV7JRBeMYFEKuEt++Oev2Xee0sW5n
JqBcYnLaDWVHKL6xmzGBN4TDqbsIN0WHldbqFkRbVdUEYO8F43zJBr+y9QmpylGB
H4EEbyFsE8WvyvmQeRnh88UFa9PeZThhNztQLlUwNxhpT0N/MQJbaXT+uWtm9sXA
jm3O6uNuxg8veoAhFbIFfrDPaDxEPm/V1m8lzZc/9qRE0c25kN2nVmJN3evymUXX
1JEtSapACj9LX+ho9jDmrpqnv3/Qr9iBU+1auPcoqpwHEl1TfQeircFRf3CtxGq/
70vXYwaasjeBrtIxtEGf6/+7WPasR+n4EJ/gLjELVUIMgGN+pXlGWb1/kF3njHRt
xEuVDArfCFFQTtefnvPIDiT2unqo0woGq7zwBmrMn2p+g4/kU+Vgta7ziuydVFyq
iXBeyRpwnR1UDs2xvWhJuegYa4NE2bHHJsnf/AbrJZPdNS0S/ttZ6NHXBKw2blgi
l6zUPxoDCFBADBvGDq9zPo5MXh8VY7Wxh7GhmQlgrJK9rem4mP48TZXyEAiySR3J
YqwSP5l4xoo5uffpKGRqopUX3JNXMUvZcOsSMGGSmOnBD7Z9TU4AHnBBqOpp8flI
xllvRjTLeuh8rDGvJcE9qYkQpUHpq0Y1SBKVVyxzaUtYA0Ge3wEmPM2DpDDxx3Av
xk/ldafQX7EfTlhEi8VVQPkoNjTeeGeRDjTCu0ngM9/ZIfk4HS+jgGzxpqO2mPlw
3cts4JmEa2xSK9i6ZJDPwrf4FOyPB3DPaCHJTIHCtBsdFXnPtEpXtQH+njfxzdg4
7z72zZa0xaX9Z6+kMTuzeQGTMDGrnUtJYcQDK+aeYonERR1ZFTUwmIc5hPBqM87x
zywbeTO4AI5r2yaL8l4/SIjhc/4wEIWEn6ZwsUSqRwudiF641hcD5HVfsLuS0tbm
AjdEU5a9rJbC8Mc/UdmPTBToXCwrABt2r8e1jXjzWMItFtfKRlDPaTceUQYgzSlB
fHjEMloJ42opfPup1bu46npqsZnbDopgBsw80eN+F+Z9BkvZA9v9wIb2LKfgymMN
1ZLcLtu8/LG1MW+Hz0XZnmYtOy60/4xZJKgSvTeIH0/PzVLwEyTrmJiPWGtofJTM
lx2sqJelrTP0vXQLbQ3mpcT6GiASTkjG+xnQaST+BBaDTZ8cFKc5pIV0vXjBMYpx
iFtD/yf3ai+W/r+qSURhsueCcUuveq2sej7yv3nCUi9gwn+9xjKrhNm6dwwi16z/
gMfMd/DB2JW4WGDXxcSYALAb+fAHa1FVTKtghrCZ114k4L39gClLJCiBfD4mV3pI
wzNBuU+SY/G99h6UFCJv4QMJUmLqG3xtkSSPimLVtELIxiK0T62YS5MjbmUfAnYv
kdlboW4TkhM4ER/+O7PydFnsgIESYF39ymmCgYCSGuIXVe0y+E8cg8W/3yEXqR6w
633JkI3o/MjbMcWamW+3AwC+aLpWv5r5uYsHjfs9rRDvekec5lilGpL1EPSnhkZh
TlLxnGyJiMaGLyW7JL/MUlbzQobT202GxBN421IPxPRFkUjAYL5CGNxZEf5KPMeO
oRHpp6QWjWcQ1j07qIqwIwE9PPQKv/CqIE3R8mVYZh+CbSOgWupd+9HoqWl7Y3lF
SctfQy8qXzeCSQAceevr43q0mHGsMfgGwAMsWICyGOKOnmAH4Wz7MFtXKWqiHyBp
teClA1p1QJYENLvTyC1b7t0+AuWH1aeOwctyJ9FggA9UVRoYDVuH3cIzFeNlu8xO
kuwea8BbqPV9NUWPzJUhKQBfK9WbOT+o64w12GJUxGTuhMtr95Phz/3EkNXaaK0P
mHiOlYapbqtAyqONMXSSkn59eLrhht/Ss1tcQ2mVW5nQ32SoKwr2iGJsq16PJ96X
tUfuSzVf3otr+j19pIbCAejfXeXrYylBwuICBFw7Iwv2SYVUgfIWmPTKADTq35a8
Si3LDOOTDuJoMLlZLEqpfeZkBq4vzpDXngTRUeej4UTb5ZlfS4KEXPzH4Ydm3aiQ
S2OAmrIYQq3NVa8+sEXJZkM7JR6/pmqifK5JQ1iV6ttZiwWRq8V65Xnj3TUlWVgo
dIBk6jUfr/HiPRteTDNL3NmIqlAJLTApuZGEQVdsFZaP+fXLNmD+JO0YPE/NRfVH
7V4GXw1RDgZ5q8n1N813ZIs1F+vAkebGGS1OimAANJzuAZpkJQ2TggQLEBiYpS0o
paAexzASfJjykWlSNNYc1AkfjrvaO7s0h8XG27EgdCC7Nk4xxNHu6FvR/xShnI2u
rLKjqs2vtffDCsPRXf55z7qlfgdwhD4j2ZQWvea24APnbnY/XRtogawrbM/iqAXM
oksMhFgBgfXF1yARdY91dT633iEkZVQpfUve0OVy0u73cYfbNNToYQWZ0COCD5ho
gkEjj37sUoNbdExo+xt6vJ/tFgEI8zS4T/H/XWQIkXiul8ESwpM3H2GiaHqIFlBn
3yo2QI+vyeaCTkL3CLiuEnVdbDwPnrRDlP2oHsj7c4oCnbU9kFvYst7KJTh6wD/5
kegY36NynHCY3N2s7ILBv0VvfesAP4R8nwXUXM3BlRmgAXuwO8gVRpcanFUuFsuJ
cU5pgDxXq8V8C3565PZ6JPgPpdxlt0hKLip9eqDoeRP7RnDhABYSAKHx8fOxGCHz
cxBqP7mU/JNuQFzbkmC1lNKk7V63qeXsJ4wHDIBi0u+lsynJgFlUzN/qqgsfXBIf
RQzhp9NxTLh0MNMPv8X8JlgiiS8/PbvcooodhSxbg+OCaWDFtHlf3jOsxo5Bzuj4
lGR+Z1pGK+tMW7hqp3uZ+fe9JrMagZK/Y7xr+zOuHyj/XlNHeS7w6U5usf7g8wKe
ru7zDeO+P4eSZRJHRZWc42UT3i1QivElWWELCg3GosXjx2jbQcPh2RDxlNchDebT
RhoHOyRekllZpROpS32+f3HqpylAAPNOiaRGbdz/n8vgAP+GAbn7+rXy2iRbS4d2
jDNXoseFqoFtuQPiz3bcClxOLeYzShM1HF5FtIS+u0uczCQ5lY7RUEeO0Pxdjywc
8SpCIzkRvNd1CE0flaI3XqCD/mYOihmb0r+A3XxMQXPyTapYCNpxrg0X+Am00p7t
plI2OTj0vclHK+Pr/IUA6eNCO/tDnRmQ+ERxvnJXoYf3KjanpV6M7K5MZgJmsQ8c
neT4pTkj4pJyy7nEDy0MvK7B8EIQEXRMgZRTozlzjJYqNx8y56Cu2c4WEAmB2yyx
HjCz0QkmVtlqc5iibq2rhdSzUtvh9g1WefXjU60kDK3RSXReiY7rT8KTS/wGc1aS
e6ZKPovVRCr9FNkkQmxoueVmqANJshvrbYNSFS0OHMM1NJgj7pZxqbtyDSVi/g2W
hUbai9kX09dCWB2ZvcvxSXjxYenYPTJZe0+t04wqY584qgZZ8p2WhgEyvVFA8L/b
DJSEL6nbnQbS6B1wxzx7Upr0YC21bEaK9uHmeuDUjewd7d0T3CX+Z1jhjLSnZ650
4EyKsO0WQSMQ1P2cPfRXqbMVjQK6ZX5ikejXBo5TqyvVjeXFxa4AAqJvdoiUIW8Q
UQgzTBVmXiPdl8kEEp4RDCweWjKaEcDOMMNJ1ipadfQJ/7WSi/TLdFGMXwtC4p03
PEFr/c70SQqU2szi+oD5oIimidzV3uQbKdh/4RjeUcVCJE9NMwXH6CuE3vPir9Dg
tIHJewBC1zVfx4HxflaayBYyJP0r3+6IVrpQiwUCjDUHVNDjHwtMtgpsqWnSBer5
Uk8BPyHu+arbf8b/dLMzqdrFSJA1fCjgZYovqpVBCoUNuwufrGA/UO7hpqUOZUCz
TUZdENkhFIgBzWHPWsv+y/fAufs2BnyIK7F6OT/MxZzlBIA+RWqCMaH6XtFD809h
NlksV2yz+BkOFhzQaoPAMWUqWWYOV6T93irk0iLTsSs+PpYuJ8RFEb+nje2DlBqn
RErAWeRo9Fl/NiHEQzIUCEEhBfTLh7bBEPtRsC69igDvpIW7N8N5i3RnUcVQsDUb
gy0fqEw0pf+94IoyWbQhVHip5qx2FGqpD7nsiEm8ENOzbMInhtsP+SgYuQ4Il7BK
J0aMY0Qgd/5BOxCBS8PqTiHdkm6TnXeyhqWnbc7v6qL0gw55YsZKZn+8NRc6gbyP
czyS+Lf2j0RgMKTPxtwVJbp4G2KOkMXX1mw102W5PpJT3ruWduISD80cjjFMBLaP
L84hTIpE275oQJlfura9SdP+I+GFC+dDHe+8CJVy+OtjYPrXSTMkUgqqmyjHpB6a
izna+1n3rxE9WxBzNrV9rhcCt2rQVn4ZEfetBNei2TQUIR8Sl9u3lcPTPxFyuzgq
Td/UPn3UOf4CL2bwpWTH29j2mLoFSYKAqmaBv+vTuyDrD8qjKQMxyLI36E0Aju0x
ioj/PGjz49aNbk9MUTQSQ6Pp7mZUJay/1cqnEQdyRWCfzNpdnapzN7fj1cnFC+2g
O5VK+wFkgyC7T5Q3bH2eT/MhSGkomEHg8wis4uKMs/GUVDuyUzM/9e5gVVXOKhKz
YugTEV+erYimOAEZTnEMsGK0eGHJ+fwofao5G6Jk25fuYVdk5hJEY2D/CBguBQoB
8e21q+LnogzvDN2JxcaWmcRERPGeSuxB7pP/R4obxTxMkBKek3+SihwYN6JdR4tD
9sBJSzJrx5PR6KtNioPQrmAFIbgYpUGEhJ9Ow3+8mJmzqsKu6c3PEJ6hvqRlk/7/
IRvKLmvNMMnPY1efCWW7tiPzEj7K9H+IskL0+jSMzDPF1rXdCYb+OLKJNXogEQDf
ycBJPhLeORWfkm8Kp5ka+vFTOFVWod8bnESBMGYeN/3nzESk2UbUGQqk1nU20o2s
KmOfgFChkmuvAFjpaZcgmFVka7s1I4mlL6wqvZazzCkiFogX3BcxCMVwyoNMxvZG
kr62IrhFdjT7mN6VekTnGiw1cvS3+bWf/+mv0D9mqWT3VMqdLkPTjLxGU52PXVyp
mlSsKZoe1FNdngxmkoxUSq8UtLtQCA3IEDg+pftKe656gxVMYLWLRFRhk02UBDdS
/SMAdkZsj0XV9Ul5kS7MHQ4xshNKft/LVvtG+UiW/ImpqOzXp1Wpvutpds3ldWho
9sbS0Am4gr24AQ5FDz70TuhLBG+clVs7LesTk6nTneGWT0sVku54KcX5pfK5U88v
DwfepR/eOEhB+PHsiu5WGmdigUzWZKn18w4ldzHdjJ2TnI+DxFnumUYySLxLnZAW
dDVJ5QLgqrrVlbW1JpSjoKmbA0/wz3+2EDOiRGLltxKQFt5dMd+TggFthDicRF31
JivgLqptZEHmW5Z6B5wMWe104XMPbuKP0L6qh8SDMMMPaU8kLbVk2Yd6iriz5ktc
ygkUYGkqLKA0hmgw8cyJb4e4nMOTl06JdIeiyP0Wm9PQqBH5QGDZPALw2ypsEFtE
KU0pcGFfWTXwfgU0aOTaCBuuM/cAo2nNHsCcWqrdk6T2SHxFSpsONUETOnrZwdJw
DS2+oHjU0L3SvtLfq2nXWJVdH946O3dF7aVYDy5QtHIzu9c/2+Jp7EzR0Wesx8in
SM3m2eROx36wNodnrG16+nE48sdFIR45IQP+q63LnxizYOaymYeSRjLjgqy6OUvQ
SEYu8td62T3ga3xZBqIO4f4Lexq6vaVHgW0CymHK4ZjWgt97m+85J/XOuMAfbxc0
Pe/bsNEwGaxCZvohIwtx7bnNBzB7NhlUcW8UJbygYzbDn48OiUQltlJVZiNWCr8l
EtUkrvgGLiq+IP2XtEZxh9zxvWS5GloCnrhs/TOhNB/+rSDXXbHd1kGZh+9Og6xK
NH+skZebN7lYsWHPVuboiRiJfC00GjDZA0jz4u3xXC3Nhd8s0JOfu6lOH67laFLk
ArASPOVE0+vpiXQIkgSERRDzkK/MBMg0D1lJboWPZhmLHlyok9FNg99gsJZyEOBo
yEQPXlZfgdRsGVqO45gEt9jBngQrXA+dJy1E07sZmrWf0eEtEmzGd82CflI/Hw2q
2jseStowZnFqfAuwkeAtFsHVbpTjE9NDkehSTVnKLZwPnqjLep33qVDz/YmEjkYy
tRqfNpkZTIZXjkTQj7cRKWnezIKNbfiGiFFTsZQXhlAyM86uVr3ou2MRNmAVGUAW
1/+BVV90LqSTSWaIHAReY9EYFa2ZNH/UBx9sv25tMuYGX2UFGW3iBkYEBHSU8IMo
bNO96+VA76VNWWZ/DyPgeDqbQkjgBKSBLOJVL+6eNOHbo+W3e0u2LlVYUlk8CfAH
nOqmVYYU2BZXC1YRCj0gEkRvsPmraBDQVSEjEqWqqntT2ULC8jBqkcKnvHdA/QJm
/ahyvFjqff37ZMTQvJOYBceed3K2ANmE+THmdyY1HD8QaEDkVJJbU5UE9w5KGPq0
8cAjmg5rmkZP1BCz0C8hPwSF43/QTs+ryx1wdOQu6wWFX0xJlQgaafrDkXyrtOAF
EgQzFukGQenfBxSY35qBifS9/zDPferdBrpGbS5KqfS1dGiNYYF14BZPbw/wQ9u+
mP+EqSIRzWJY95kuwIOBge9ivt6lOxxas2ty/LeWwtaIsILKJGJ5URzcJAZiK9Sg
4R/hitrDYCAlA1LCrP0LXh5RGpzcQcUgA2VxCcFP9LqYCoRpgvT1PjKryXWwphsZ
surrgfYRhb49kCT01BE3AgUahmLJy8+wH4ykx38GBfV1akjJY8qxpZnBdrzNHomo
UPuWsL+kewqi87l555DUO/XoSDdSTHVeiwHNDQvaGBZ/BxjJRfIn9F/YrYDW4e91
2AiYElkuTU23u+GH5B2VYbbVUFPn+YXK2LMJdXpmcFgBXmsE3Jb9VfqeRPdTNTJQ
jfUeGhbf7T7yQCXNlPYwe/3LxZ8CvguTms3VGMcra9JncKTzMxwclvhHKaq2U1eX
eAECdiZFYa0+YRW08Xv5NVjzlsYGP+4zGslIWm9pw3709Lp5D2o2Ia71Falg7GGK
Ot1eEgRci4lGs03BGyDXQNpFURZj37QBnLCUddmP5H2G4T6FKbvrY3SLg4p5Pd1e
oaLviv2/ZxEN1khuvdjcbzmlwQvLKbykBwOd/rH1fQ1FkqOx4kRvx+Y2Md4dNAXz
oZIElZeuyYIeC1+N+T06lzMDj1IfavwrG93tOOp0B6Me3roVfCW57NNfaaLw8x21
wBS8KwdOqvltmjAD6iToGqET8TCaYF11MzsMacZtmVGpaSjM2JZqukH87vD62GT6
s2luGHbFXbt+wcrcNRNcN4mV5MJuEpSl9uFDWVi1hd8kCNOXbpx3js8CpP8e1fdE
qBa8ZSGfI0Qze1ed/YsAJiBmUHlkigtrXoCoSzUx36vH3KtQFRk52bR1D0f7U9TA
NG3IjEwR983R+9FSH99yOJd1BSO5zJDm91T/kn369EMPj1ydtlX0Aea+qob4yoXq
mLEjV0aZAYltCjvBUkH2fAXaiMwrrap5EhtHoDn71o51OMXg9QtgeV09pGVvbGtE
kdeRLx/yxeAzwTpXzVywMTyvAQcWhaGRnyUEUG9NnYm7Cq919D/OCohdlXIR98O9
+FJSZNpSbyx+leeU/lePaNFYSD4JOLwbwDLxK2gL14Vgu9BkkgioUBf+hgwT8DME
wLhxpBnarl2YU1Q443exUA==
`protect END_PROTECTED
