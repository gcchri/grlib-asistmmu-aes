`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tS6hmKJt/wB24K1V3+In26Ec+rEhehHqL83mbzXvmytlNt+iogmnCiAk7W7KHYNJ
347F/RZ02a+dQQQxACZi3CrcheqPOlyUJ7jEKyFYN7Rp7q+pzXAnhxgi3gW0pXtn
+kToR2F6EfcuTnAW2l50zM7qV+PKYLgjpZ7mxys0k3hdbTf1Ug/YgHZCIch1QbC4
akoU5xN6yG54SO2BGxU2+/WqkW91Dz4oVjFnT/o6CY+3E0OEy6mWcgxy3zwV2my2
5ASA9BGfYM2SfFizU1rmNa0rMV7NJOXWchtaKxvn+QQFEwQ9BerCeDHS83Z1pgei
afMiViXvSQs0QUR6rmS4ghdeZWmtwIkC5ZhNZew+gyPM7B0vAyy3a8tGmp2K5Gye
BXuW5fe4jLY1wVGz18RBPEcAFB7dzqlc6kaPobQWHQhABrG8XFmFxsX2wVOrnvMq
1mDOuYCMltn3Idp103P9+EwBt1HoEQBDGrUcu+QE9HRdemFRgQgA3qJef6y9e+Xn
DnQxnbeoJRo2a5ly64HMRGdaczQhUomfCBoI1ujVZQtT16DHoXxJffvLastn87xV
iMHsbLlSYfPgOdCILpuUwZirEOilvTKrWktPkVrvuIpMVDTJe8p4Z0A00OlO2vZw
nBZFmWq7ckMtXD1l9S8veMwDihJ2QxF1m/70pYF5Icpt8jz2/qcS2cbTsDAiXaaB
cIWRHISmQU/N89wHlcEOqnaXCAV6MsYaSTCoTqdx9sGZvjcLKHl496QhD0VhHzfr
9XQv5aJpobNtAoPYJwIVpA==
`protect END_PROTECTED
