`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K2YZXopGxxywsYKRiRqSIQ3ADBz3+bGIddb2AJShF9eKQQDkXD2Und13FKL6L3rx
n5JIM5Xmj7YU913LnrbV7W/JWAeCkFbpIYk1R3g13rT8A7c7a/wLBx4L05VhvAgh
8xz7y+9d30Qu5WZR5C1s59H/fn72CkPxxOSxQZsEyPLlnJx3L11ZdolqrdxeZv24
yzZyUFPriP83EeHMlDFWT/2s5a6f9rj0bdMucd3F+RQt2PQvbvHnsm5D7y3yjCyy
P4OghMdzC8GyGD1HFb6m/cJ87osMGDzr6ck+AdhySls0qg0xnsaTz8DR+dx6QVUh
YE/OUKwWuWVHucITlgAzUQ==
`protect END_PROTECTED
