`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iPCBBfd8wTdU1Wmqse0kEJ8Ahq/ueJFIDkc8Rqp3r/zmJdXP7T630VtPFJ64xMWB
EgRt57G4xZtztEcBTCqWLHZOC3q0AmYFrHLcQvKLpXt10lyPlvDGmVQOHOYxJ9ng
KmPpFy94Ae1ttNDPJuP1T33vYEgPxK/FA5Dzij+GxZJq0SJIa03nljTKCHx8L8pQ
u3uapYCglV+rMAbvHEVdEkMeFhzvBvMbY+DwXnihLYZimWZAG7C+J1+Jn+sRogPg
SxRwZB0LgCMIT/T4aC+ZsAQekOd9KXYmD0cfnSqX3MXFP1+3ZQbOFVQcCM4AYelL
qNEGCGijc2IIZlWjjugbB1IlbKnbM9eYXL4o07c4EwwkmnNPTpAlduWlnvbUeKZb
KD8VyQGgR9Itl1Klj2olBI7gLBD2uLyraq76Sl3X12xIfFLWaJjS+Bd8Ma5G00qF
wzxNwoM2uxlJH5pptN65US1TecRDKltF6RbI4SqaybB5yWY/IUzbmCw/YhGLKoNl
a0zS7Z0NnUPeMZGsB1fUBtC9nKtbNXUqpQq1FGqGvTAc4lRn2uTJFcsYcQZV7Swl
Yu5Rn2liD8Ic9FbwOO5t54cSBuCOO1sy/FBYXPg1DG4=
`protect END_PROTECTED
