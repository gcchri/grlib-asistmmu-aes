`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TtDuHyYbQ9QFtrDloq18xCprTJVg5s+8ahy1LBZJbwzdmwtooAqGUBF+CxJ6fNFz
7Uv2ayJUywBhyL99qlQO3GZpQrnYAv97qkNNA7/sDCAVxNUZ2ZV44zDYGYScSqvZ
JBaU1Jyq1TVmKUNnwIE8nTHLQAmoI6wNNpgx2HnknuXs1zxTKJMhI2ErX0j4uUjr
WGDo+C2zqdsrmF5jf4UoWV2ccwQK5D8Sgs/q1MEbFoB1l0c9PACojM/Nlfq74FAE
CqgAmKWdW54fktHajbvmn3WJ6XQ6GJg1WnrOTTG0Oxr2wHOFkLJZK4jJ5Kl48ghw
1EgF767U45BvqyRQaTSbYUfvj8fYlsBw3U2TSfEe3pdqFHQilyS2Moce9QSC5cx2
C4IKxB5g6fGIt6X7WA5CPmS9/V+pzm3U7NFAhdGO2Lx+mt0+mZBd4s+BTlzV+Lly
TW8hGgsRdDI8wOeBKfjqXChwszAuBvz2jkzgN3yt/F8=
`protect END_PROTECTED
