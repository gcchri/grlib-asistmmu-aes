`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nRD5vz9bAr95VvOpS2TjD8/c0VhBLscZlDWRg0DyYMH8XUHXHx6SMfKCmnrEJr4V
9wjQMp8VP5rC0tUZk2050zISytgTu/WJ0CGUSby46WUOYXNpnKlBhyPWcmJBSF0v
DmQR475csaIsPOZHGanu0qJ62PQPVs8cEXOD81ehwIBmlRexeywjpqlobxFFGZme
Y5/JzOjRZZtQFzHoeWqqpMnkd8w9ldiCqf3GKAWMzGrqqSKgoF1X9OpbACDVgTXV
s22iRdz7Xto9eRD7zBHyYA==
`protect END_PROTECTED
