`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cLaZ8o6y9NimPM4j43Oq6fdrAoDh4uot51MAXNbZIOEqPWB/svZMJNMWG8d+tLA7
Fd1lNGHf0wV3SkuCue/wgm8TrYYmif7eOL9TEeVVuqSPke99/ITRKZjuq8DYJSZj
CXM8rqkxWAydswqrNwFYjspWxSBj7G85VnolZ8Bnxc8IHzZONAiBHbpGh+C9bmuV
KNobA3nR94SzO0rsok9zhUqnI2M3v931gKVyBU9s0Dx3qPTPtaqYb55oMnFWaS5K
bCXds++7TaYJvgVW0Z/9V1TI57eNQyfPXaNTyP/9RAEliyd4Ophctz2UfriLojan
8VO93KuajP62BjPU4P5fdpjpNOq1uNFrHeqJ7nxj/V5p/Emkb7bE6B/wE9QYO9QN
EK8ixFrrEKI5/f19tXJT5fH9WQWdri4Sey0/xKCm+y01ikEAKDQoXTVWq0hzVyLb
MTf9R2rpydQGCxgyFRtB1Ql0JlE2z70a608n8vKx9el2XRvE/QbWNMS0Zm568J8q
TEjOwXVP9hGN89bPvliFvYNIyOiUrjf5tAwTI3TLQiD/0+ez0u8CfynQKK3HbfvA
j4C/cb/NIUg/oLqh70IszB2lu71KIaCBlJv/a3IZtlieJHJ797bqQ7x0Tkt5uxTo
xVjuNMHiOMz+aCATTiU2+I1XJsV8moYOmgR6yGnBUov/HLX94Be7H4vYSYvBAFw2
`protect END_PROTECTED
