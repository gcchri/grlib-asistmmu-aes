`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xCh/7FKAPrHoSdqQSxyResoQX+Kvwm5k3O8w3e7VPe9RF0leJ4O9VW8MpeURpi3j
LEztCrCPmXAO5SZlCTidYfEidJOhsF2xwUwRx3WfduBqcgwXyGjm0ilToJMaPIIw
fq8w9AWlH/Tt029MsI8EE2WlHbc2BnQB0//vhYGzXsXYCEUtXs1U1jXLyuffN2fZ
leaTO4bOQZ6F2GRfPRBR/QLHOHY8BFrObagVZM/DTmbCcN8mu61whuoF3HqVvyZp
/Zv1aSdVtaZLGLp18fNjY1S9pMTaH6GTH/Gt3+Xf6Q/dXO1QvImlS+toqVtVoYWK
ox4J8w0MZ/0N3WrXn+b5ZAifcyexKG29uW7lvnRMjJugCyd4qSe2e/KOyhJqcrSd
Rm1ZUqeGUD0mRysssfS3k7hWkKzuEZRBWjE4eqOs15p+OE2ZDo9RNuY58I9eLyiM
60UPwTZBI0Y7Dl4RAvR8bw2R8vVZPUNgSycsJiQNZ16iBR2/ynJuxk49+AIFkpva
NxmuYcQ48eBPa7b6RbasWppMbuWk73sY0Vx2haITHOO8uvY0DyyNGbPumzv4NsGk
QGFQgNPwUpUmwZkp5Q6/A2n+XRroPzT0gCJXawgh+lScZY0gy+iEAGtfBeKvIowM
TEXoeXF289gU3h7sa9f0e7o8hQeyWIzINpXTa6H71r8EuZFsdY8GT+TVNPY9bd+w
UlJlZ5eWaYeGInzcmRFlmJ74/DTWQKYduoEqjYU/Rq07lSowvITu38m+Cj52Hx4t
Ik22+C4s9G19fCo9JijRWxaOv9ThYi3M1WK9CdPhuBiIhCe7dvSU4oCULCxS0n4R
uRgAXwFacS0h2AvATT9Dl3ze0mBkLPU7eH1FLqdQZEoup7SbL6w5w0944jLsW9CC
zv1HAKV68GmlswSpFRv2+GryDWAlTYzlIrgpFJfpE0u1NaHa4QosYkFWOLxyrp6y
iXxanEdbxOCWKFLtzZPkxMmug5E8gYYBqlQbwoyDyp+8MBqXoTv8TJBmNKtseoxO
JX3GghGbp7nhGvASmnyFmXmazBFBuYUxcWwhtU/biKOTXuCjf1B6FgCIJ+RDKT3K
humjU7ub5wBoJGGFvuM70yEceM+xrP02VgGiKjvUcOkiIH93A+ph5b6p8JFfM4PZ
0D5dE2brad+4yrQFcOjMoGbdwxcmLtc8xKC9xd6OjvhsmkuuJITno6xcBc4MENLV
yLcEFibWgcOLO35R9eJzmos1erl46Sz56APgpO5RD9JwjktGXLVQOtJIq74DLLlA
`protect END_PROTECTED
