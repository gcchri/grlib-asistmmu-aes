`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OUAcTiXD4MB10mnRSRGpyeGIJ9vvRoq6ZkeRZUYsvR+7KrlUxRHX90gYRI5aYyEf
Z+2vtaEcnElo3adYjkmryf8juLW6mLewB0444/fPKFQ4kzXwJwn4zlzlBR2z6Y0G
f9tlP1NOh4RYWVuSieV+BZ1tSyZ5SwLGUWJ9/yg/jgZoP60qAATlN8Wbzy3UpM+k
cSFpEKoEEmfundUisIRS65UG5H/QVmNVaSmEGsls0h+kRD/0glHeIfOrBklisvqc
dG0KsnhZmq/U1YIELYKf48ifm55X6fc7Lz2r6uHU/aGIsjT7I6aJ79wXL/hH0MQS
6jHzF2mJY3g+eheuJlAMjXjWRizn8FHzNiqkWc3Dd2OP2CNK+1d+dEybl0xt6b9E
gfcMCHHhZC29i2M5sTjkw7wzDAAWfWleWthlGjKsaFDZlXaUo6L2s4zYebkea3BW
4GN6//Z8k9bNaXVSBQc43SngTFrKbeOkDW5AHppfbCPplFb4NL/bsGpVj4e0nDgB
Ob+RHsuz1iU6Dmn9BT9iMfGY2ftsdOylUMO4l6LyhSM=
`protect END_PROTECTED
