`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n0i4W1yEpL6uKcKvGg2AYrQ1T9+ESmwf6tBFR7evZPpnyG0EL5jMvnP/EONm0B9A
IEqmNbKlLLh62aEYlbtvAzmjzJ5n23GSj5NeZw1VoUYFmI/ULjd8HGjSiLo4CYcj
NZC39zBpF9VAVT2hm6/mYorSZceqmfCBS2srxJNrIPHxCyN5VOwX0/qc1NPRws+p
9OshTwWKC6rBXGW1pNNSQe6tSv+vbNF3PT11sJkenbsNe2zk9m0DtnjiZYEsvNKc
8Ri04wM3avul5L212mQOG4o4GQAPLe0v+BAA4+pxpgS2JbUFErPlKD9vi9RHYvnP
xNNi0/VIvJDQ1w8QP9B0sLac7HLNuZlUusLALDi3FUAI4Wd4IyesQYmXWQbZHCs0
MhFpICn9XaWTsEay9p0Yw+6Y5dENR1BZ816zRf32BvYW8iDbZWNzznlAf4ubvRVB
A9NP7bjYZbE0dQ+EHp1QK3oDWZn5LaoXt58VrNDgbJWJJVaz2/AEB5eKXsiSwZff
43dJgQPvMfu5f8o5Ns4uf2G5osOJuF8RzizoYvD0uig78q99P7Wr5X5iJmGpvXXk
gtmkvrPlRLL11/Cd0wXyTdwOuDfJq1j2FJhRJ8xWj0l1O1+qWBfNMZQNdEfTORIa
l+drVFPoEvUFM/Ys+8OC+zPI64KxS02v2TJS/ujADjkG8u/2E5zyfZgdnq680Kia
zbgk1bOBAqHyzWlUhxqrDTKkVDlK4yywIp57QGEQG9VRmNIzAeeu0vJoWHu7XR1+
bzSc2C5UR0DDBiWjM9tQn2uhDI1lcqdhM7qIiYxWwo2hsQjawCwaJnqOn0SwRHhM
ul693fF2sVq3szzdRPX2vxUAQAdiZslWVWZsCqjeOXldMgltU8IntxR/zn+PkKV3
yfxkGYtbzYIVTaruYy+DGPoyf6cNi2pTiXrmbXC+TOU4q0I3ijfNM96i4bhwvBom
xQWyZWfEBT7sr4DdUzedKdPOSs9YU7M3bgG+KXsruOumoNbDgSoArf3VDsr8HewT
+/3wOVAr+yKnUAwQECWseQheRqecoVghXNr1QkXKOrptPHvziU8eiA20a8+vKh0z
XXodiK2fD4SFK7oOoWw7NjBqB1/OPRxUvaJJoQIMIT8Vpgqgq81+/W09plFpJWNa
OIHaz0MP1qQaNLmFXfQzhFi0HxjiKLJ4Th+hjBxirfeYy0KT0/cSPypJ6vJ8ZVm4
1TNf/8deVIgnZL2JpPtWdMxwrdwJGwNuvWShMePTumdZQZpfPLOUXt56x5QFgg1F
xtBL5SRqtwxhHk41Gs+iGEf/QJu3B2vPLQlbLzRzwkkjlbx47byYY66qZcVMgQuX
vq0rk8O+jEpkYKVGkFxYD2nARu2qeLwyqBcROsH06ODEwhVAnqCDcBmCdjtNjwWN
nfg6/CvmYplka5/rbEuOYW0KC4B+BQs7F7P7ypUZWBtBsJpyOykyUaMOPun8EId6
IpfFBFlX+GATcek8svKLLxrr/cKZAdRgwSw0WhyH37mvaStbYn4Vf5+jj6pt/Hs1
U/qGvNEr6krhfJaP24bXufVkfONMSKiTe/o4Nf04k6jowK1oCEQ0SF+VwJXpdPO1
9jpUf8+EBuLO5gXwiG9nDNr/+dl91dKiR/PPuLEav/q7lbbsq4cgMo6fub13Q22d
8dTGp5MedEYy8329VkyXyQirKVr2OXf1jaWJ5FKqITl2ctsmCJLBVzUg0iCIPkY3
fpIIhA2MmXCB5zbOWbOMY5BeiSVyKfS2RE5OGrdNNjbZPeMxqLkp9pGW18a1W/vq
KpiOvA5BE0PLF+M9E5XIMhaExs//4YI0RBgG0DhNVuWW6thuWS7iSOAKeUdl8UIn
QxoG52R80w7FRDjeKlxbIVwNaFo26f4wOHkYfDpv1/+d8pvV6SOy7rJub76DmdqX
bnL690v33wCFbPQkMznh7rFvCUUFrexl4RGHjYgt2kMpoV9nPUL8gt35EBJ2xTLG
9PsmT0d11UIXRlSPvS+kFAYdAbPQLdGlmz+EUQWO7vaO2iiiPa1HcPCz55OS+SU1
/JzlzEhs1i3oybCaXsmD9/3uJPanrXAwAgl7agAwl98=
`protect END_PROTECTED
