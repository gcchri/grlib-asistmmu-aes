`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cg53jZgDgvX8zyV309toAub2ESACwa9n3pbK13DZUWB5X46RIbd9joCFiMtpAGSe
bh2zPjgJB/W2Kv7kAj5ptrOhIni6aYslLkfrBEkCJ8E5gjmTABFweIXZKJphBU+o
bHWban+QzcHCoWxlBdv0zB9MDFU5e/aLF3iqs20ZyTPR8juW1YQ9E0EmYb5mf0lZ
Lf8cBUWBIVRVlRDme2n20S6VDM3cy+C/ivOZdGHS/lR55rFUGRMF79Vq6qB+RPS8
uAviyaWAS3aMO7ZWaMtjFpt2VUW+BY3BWRazc9xp92S73Hf4MkVRn04p7XTPyR92
9s5Waqd3jtQXAKc9FfMy//V5GKxKIXCFpyvjwMXQBAtQ3hz07dm7wi90wCGvjPMp
xQpIFaEPBaZzZ2EWQM1T16cFxsOgENVc5FEWYzdevLHGPOtEhYBRO3IT8/5ezFBA
Qt3Rtmt05GJyOQfKThyYxUzfSJhnD9QXwLl28aaRztv1R4o0mGxm8hUfqcN41pM8
XroMG4yFCkuC40SLS7+ZVBLJMmLNAIjsyzwBcKx+pSIQ2NYBD+///gYswLnYGMT0
h4eCv027beMULl7w3UjS7ITPS4j9Owt1elr/lyzw++OKZ+p/Xy6AKXFUTsstTfjB
Gjyk7oThAFvunDK8zXxp4rI+y2yhhb2HruuLUspTlhMQevLDscfVcO72ZCSJRZsN
GGuUBre+s9abO4LyecwXnzSErlc/ARt52qaafz3xQxPZyLNXDwI0N2o6WbFwoWrh
lDS7Tyq3684FWM7/wmSD9ukFC2XR1X5YilmxIH+xEKGOa03ulzmqHDBwRBHwMzuH
Ut3BFAV1DxaVqKO88RCtUdEDjUcJEOxq9l/9YLOGHMW7XEGKA8/HRtYxu699gMh3
sVkulDh6bJO5J0olyHnvwP6MWy148Rbr6aZXy3kSqUok/C7Pi1A8UWtHpZjpc0wg
2jFUYW2e2V8kw13YQ4jHgxaI3BwL97oKas3zMgkQDRTEtTY5xvthfnjTsL6UbeqD
fgP54LO3xchhuRGLv6aR1LBDrwh0eDAeKVtn5d/v2smvd8sWd50ch/Tan1xPzP9h
m0mCRf4eqwpie9mAZJVU00ErU9djbbY9a3jexeke4Wza7nNVex25QvUrewkqBvGu
zC3JbuOf7zwK2MOZQ0IzuD8eMUBZDuHG/NeVDuU9SJFAl+5sVsFpbXYR9FzeTsmn
pKHfvg3ximd1ULyVxDbsOUqOO+nLxVe4/5joPlzFsBn3cwiaegPVJqLY/p8EA5d+
5H7PeBlNyN7BFGqT5JV0H6z2yE/FRFUZl7wwZV/E468FxV6GeMG/M83g8+wgznaF
LYYGRhef6v9pPhVyK2oc+VsqhyjiIDAj2OyNCToiuTZ4T12RCKvvtI+quFOwpmRQ
rr3LQDcfKk82vPZEhNqhEe1AEfa+cetQXov4PyBbomzYn4mot2idthzgsG2k8GoN
EoYJDSvRnG64Q8pdo/llmDt60VSo5obUXu8yppNVXoR47mCRd+ebS8zWMDZG0C2N
tUdb1RU8oB+7gV8vOaZD7hteIZn81KiYrOYTeJWyAslictJMfc7JorQ1r/Jyp58P
RIELdunAjwGMIr5PkIkz1g+htjX7QWzFCCSK1jTnkYC9bUbnimgw/NqRAzkNFRvJ
VylIpEioDkHnUGSPtEZNRztmb9RDfKKfrmpWL7TB7WbemDVJw/qChzm4VZKE7sCC
oszKhBirEIBBrxZH3fitR7EoPVa+QdnGLDUfPJ0zwWZR8NaWKu094qQPasQxV5/D
QptTp5n5NWYM6Ju8gt8f2pacQ0cKsxtEu660QKR59K7wsNxeftZfk641XC9Hc1n6
hef39QlIx6BupP+0rEti+QkjnFamacaiBFjAwbEKFA4cKEZqbWQ75VDtTBO4JzoJ
xpOxcKu3dBrk2bQO5NzLTE1hVPW6aJlsZTEV49UeMVAx31P8h28E2B5Vu3YrHfpT
YSZzQOYj1+EFgDGT59F0BC8k6U3/guwk5ud83wMpd2Lz+NBSpISgG9mjxl0AX0Yf
A3MshvETluRVwSGZyfA1QTwbRtzmidyeO9U1HHxVwgq0tsBfgCB7jzakEzE45VPV
/p16fELZBcQe9bhWJ2/CCOjg5FbQu/caNHXJHjSUFoZJAKnCRxAN5tbxYsO7aSPv
AAiH8aE6soTonRJMu+m7l0PiL/G5NhKtmslvBNFDDsbhqQ0fBgcmnJsa8n9XC70o
uO+zhRBD/MQSbZDol4iRLs+qdqgboDoyi0GbcqeWVW3NrntMnif6a9SvSi3BjqR2
9AfbpmItB0vWfrxMh83jO7oE6jPeBNKHk30unPp9qZ0BUmbcy5UxN4LGjNxKx1ox
hy5b1uIilVJ+T1Z0n0GuTHxLPKLYd5bfryTtlca80oPFr0Qbxt8f2Ml7yrpWtSw+
HcqIiQufEmki4M7MQgrzhWfqRSJXy9W1O8L7EFfuacHFKaYWT9DdhNEMiAEhK+6D
iYRNLrI9RuXM2EOqwpUdz7fC674AKFofRgJGXZci3xaS+5lsxkaFgy03xxYlXbQ+
HxrDXu8KysBAudCcMNZc4cuoztAnj49Ady/77+ZeIxH/4Tbs6o8dQz3cUYuy9gaV
J1H+9BTgRlIdIW0KBoV6GPdfHk2bAIrTAN+lpntgpd1zDGITizQnzzmH2uB2QQxl
/myQUgWT/Qc3kXzfUUueRz4MvKCbz80w6Th6m3ebAWZpAJHYRXUwJ4XCwtbY8BUP
30LZch2ab9AjEvYLAoe5rcfNAIjzpFhOfjpS+/EAz+WNY6dkk3TXTzRCCP+V2vcr
OFJp/gk1bu8EfE6wnYzTUzxUwSU7jZf6zariwXKeVQk3oMyW/MvG9GaMZXOY/9bp
0wux9GgYGFlDDrHbnz9eHKH5xzOdA1q5IjDkLjp7ICbWSo1lVHxfjeZwbGoNZdWo
hRDR0WrZDTL+wjpKAz7hTNUWUMz02sCqtqFueTBevYQp6cwNhi2OIOgsQdszH0Cv
IUra56JpZzQ0Mgz3EZfQYeM3a340/hj63AZ+mR+8Q1nlKVPjQZZfLT7LKGMmfxDv
2wg9UJN87FibYiAz+cESfekUT5YYWd1G21ydEMn48O5qx59g1xjLTtRzYkW+ajUS
Gyk+91/l33GXZoBX5qPgxuH1F8yeHj1jMGPDXYwh8JC1sgS5X4OCM3Mr6i8M4rkh
nx4Cn9M9nf9QCTcKJvEbjlFb2qeaDW3hkDGiHL4PqvpQ4bis23V/jKMw3wq4iUCk
WnYJaU3JISCW43qnAx+Mo9StYOYoXeag0yymZ3eXK3kB32aZITon6P8lqGPhdzDI
rCvEyk9KD2lVIDtZhPdo24BezAY0596nJc1Do7fobD8yDtVHHlCWPCJ3bRrt0kOO
+yKgJSMiMlBYGCEdVflxUx6lgxO1eZgg3IFlL9+ELj1wl2bsvu6V8IA2Hgxc+5tj
YJsA6ywSKWAjwtC/OMpKGSB3hiW3+RQTzw8tbp7kABAVDE6GEQNoeaWUcAJb6soP
9ox4BQehE5DGDwoEM28ikn4u0nUVTOP8f8hGCIanf/ZP3MOmps00LeBi4yJi6ZuZ
F5CBRBNsJ1xhV9sBL8RYGpVpD4YgcomTTFKyH8B7JQ5of09O2e6wrqd2QvBmam5Y
ZDoLhcYl299/lwcCcWSHOygJgB99A/UyvuTlr0n0f0Gro1rfaPxYk0ctaPwzhsOe
0kpAi+h5aSWdJdMFTmS65zJ5MU8k4VWEzpI9Df+M6f08fBiRd73JBMjrcT98FM1+
hg1Jpg3s+GQcte6x/FoeFT3QBNOhCOdSyUE+IZhene/o7DPPqdFEfC9dR3d4uJzz
WluZlvzHBVOzS+72yR0CJztY5uM304qpqppZoNn25u5qHQF8023u7rBt+08lQFIz
MM60ea3Tqpifa8uQGhDJqw3YUDjX3AlHubaasWiBq8/oBD/MQ+pmOPZavLHLHpZ0
JtmIGVX4CUupVn1Z1+Csric+i9e9tKFp4Yk4ATA/h+0vOSTYQnsfTJMWYXYbHMNr
VAiNPINL8FcfY9DyHOuDhAuMfD1v2Qy44irCJO7BhoIczW+Mv2IHo40ja8JNUEkb
dyhd8N3gI43kBpv4jrs7ADngQ2as2S6FiKM1TpIakQFJir3JoG3iiKqCVNok72D2
gpKvXvp6Kak/Znwj/88gdvtry11H+zkHW/RGEOwGF3jbOFb+eJ+SQY0tZ9WVrZyE
Iop7uXCGVelO1BcAsJWIb24J9o6wmYCLVQ7igUDyQkY3n9/JfBDpek2k3LJz6iNH
5UBNWkwJYTFNC48jR612UbLLrGY5YM0DWu+ipHpThQfPsP7MAMlCoJ1wnTB9gbB2
QzF+rkay7lkR3UvQn3CZxpn4HuogubIlxe4Oe0sfloCmgH3lGunhyevHEmBp6rAP
ssbSlnvAaI/UxUm5zL4oouc2A7zi0Xz7EuF8ejBzjjONpH8/ShyIs5Q/2NlG0LZo
yQsltahUn5bmRcQfffliMMXH+s1pym/EzLjzEWzlgsKzQovIooYpNPq8ezaJs5GI
GN08OhkZHIo/L55TBRJEBa6z6iW8kKMO+JhG0RZHohp1fF0f+7aom6isa8vLYi4B
DlFwrI9jpyN9lur2UJGcQ834wEl8ca7I52swUssMD3LTbsdoqJquRuA7s8TBkJHF
T/SUjw8BsmPQ0ivyiWVyGmKpR7ycG/5bQPWq0vIQlWquPqMQ6mrgEhcd9ffaF5bN
d4wwJM1Pw8lWiaZXOjKGpi/5NOID2ACWVNArIb9VQ2Rp8LLbSjR6ZZJQguvu/paI
QiY0VlesEarY45ulnlRM/V/c7cxDFnm8jIbpCcm5pdm3vEoLkDSNeJ10L9YQhdum
5vYwHbrSTQ67gROXfTmgOo0BDj6QhA06bbpjCAIN5durJWV18R7jSQsHMGadDHYH
jdaUbnAXCQITMHTBj8+Kuyr4ElPrbdAZUOTfFJ7D47csKJMvUGdKUcWQ68vrVvL4
W5RDpQQcUgN6pvRtKDdvO76c3QHV4tjtd17724aUCfo8ix/n3mJXHPeJNIBigr87
xbUSCs9VSiE1p4diygRrUU3N3r3laZuYVoBP/SZh1ao39b+XBgq3SktIaAdG6a4J
aAIIl/VrbjNz7Rt/BR222WU27RIeywtYJGZtyIdCSnv6pWbX7xzvY+XfW+qdkajh
tYLlUEoWX8H6CdNbY2UucVALuJRQf6TpsJ1Wv8RHmhfUjLJzODPfySeEtVz1wOqA
0o2tWqVeDSRgvbHrGwf0YRmdC+PwjVBsnRIc0jaRPxMv/9e9gELSAD5tJK0p9upV
CvD2X2FMV60TnGcaHsZ4KBGzWAnBCNj8KvRyGBnkOp+lAzodjvH8WqVIQdZ2CRac
dx+y0L1CXCvj1xYZkDKbMn3rN/4KjfwDJmmGGmvVZKpEmelU8LhT0kNFZuVrTa6O
jSld9iSwDeVPcfM+L5VUf0Ku6L4s0MpXOr4ia6MPWnQE4kAgKuByrztwn2ME/ex+
zNZKMyN8dwYjMsXOSw3Jy7rC8hL8nJSS7+ww489Mp6TSgRlBmEDcAK0U+xlgZFZa
FhXIfiB0W+Eg8I4J0Xa82PDc+7wn1FPCXK66+UxtGxzkhbLnBz8OtgCr9pMtplZF
kYAuWoIFB18qI1S8j6gEy/QjNKGobFp6rwilCqJ3Ou7QOGNc3InW9QaNQgQAhfyg
PR/UWeJiOJau5Xzs/vqv6hO/mfsLD3iKgjLjG2c5hH/lUX3RB3RMHW3Rg74UranS
/n3TFVRXNlb9OynnlhFnynNiT4UE5AnzlY/a8Oaatsy8/vL069JHWYRYNDRX7MuR
eCE02YNIr/E638teuI01trS234W3apYrmGC9yy3CxAahRy1QakVskyZ0Oy0OIASC
8+vrHZHSNEWf1ggT5mf4+zbXSPTJSFtiBOW804TsQqtt52F12vdpuHDoPeTYdpwA
Zf74+Bq4SySIprmNyLN39Q/qyFm+xo9ln1YAreuPIQ4RWkDlddxE9tt7iTBUP9mA
VqrIIGa0V0/ZG9yWFYaEWNYXp8jL2qe+KId+9aYY2h0RT1fq5k9xM9EArAbCIDsg
qDE5rH99ThRByOiPEr1tiSujZetPYpIcXzsOJElL6UWcXMfZ8YqZ8YBFqxGiDXFm
ri8MmCEy3OO8l4226OEv0Wdp/ctBMMDiU2F5UGHdjqdJYDPDsHXU0c5+0tCbvo1b
nFUPR3ZayERFKIE5XWaLuEu8GTTnBrRcj13aDjw4o+N1rZtEdDTlbF+3xYQUPgYc
QAdrBH1jAUJerx6P0QSwtUBaefQCuIp8dF9SKaP60ojj/6P15N1xsJBv790hjbU5
3x3FSsMvIsad2MZ4y9gx4cc1on6tMnGIouPSSWl9I41sh+w9B7Ao9BOn7/2n+BP9
/hFkn4uEW2f5y/HeSl+fqQ==
`protect END_PROTECTED
