`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cy9M9A8BxgnGgdI7/wQdUIQxJUpPkbEk8xgjp6uyDBSkZC1Gc++wFEZUl7I5XoXF
gB03wcW8bGQrQvrvFRLuDP7tQ2FaW3zSbExH5nuB+bjZvw4FKuDIq7yJXEN91VOn
5RI+A1RNx23MapsSQta/xZ3hb952nvWQwKF215rJukAoEmj2Y8X7etsleg0NYW9V
FWX0BijkCvo0QcoiMxGZsbhhOm2GgIKyfJcPUAIcDXOMi+et3mOV5ipk2SUL+aOX
D7YD437QSnMQjfGP9vLDLFiSmZyfi9/FWWV5bAzup9S5kwu4Z8Lpu7J5A86eRPAn
wqWotmBfQp7xwNZbBFfXX+HhEfJwxTu5kTn1FG7mai02IzHYA0lX1+va/yoDYGFF
JUmGcTxoJATrxnp5v2McpjgtY89K+YpBrTV2DHUygDXs+uptzzfYGAuGx3bHkU/2
RPvsd2l9IlQ0CTfxtRCCvhb4zUhHVDGkg6KTrWI3Pgsb2xmsYKxQnBFO9fJDiped
HScqfEw7gfYU9GbynkpQ5Emo7aK5yCCf7ZpcfY4iExhxQn0yep+uhrXhCt7oZ58M
jKnwrlt14E93CvNKXn+dpmuPDOoUoqLzHb8Wnu2e9h9DjbGGqFKPOw3wfaK9KntY
8vBI3XTj2nqtcc1HIf0nX2V+5BR79MmQ86oXEeAeY3yUm9VKbZM45mP4lS8AhWiX
frDJsY3/WYpq1EFtq2xRfI8rD6iy6N2tr5MOiEf2kS/3lk6tvkyf+IpK4K55Ul7/
igIB+dGLDtHksUu62wRxgml5Mvwl8q9EmMaVEkX2tsaltDRKU+88ZIKAe7uOSgmp
3kyVn/hBzRAptHgiJR/qAykv4BGajh9/hWtW8WXmdsXezTPEVOkxs2i6FlvG0viz
RS/VTZz6SUulpYBnsqDKi++Zb4A3pkWQ5Bc6wAAvnGaVA3OQDRUBYdLTZMmJkxWr
nrVCodrpJcOHig4W54n5rwY9Xh7DnhXdcIwUIU5ZWorXDwcsf2XBfYxbVK66FBoM
9JssDv8qgbNOS3rSYAvKDK4txS0oztrJwW228NN/GiQtY5/C8nsUd8/hklCXMyvL
comxudrbmIoC/UwBRADU0k2hPFCxsnzAqAGRWRVEVp9/jXRot76dYftHqrWOybuQ
MgEa0xSObbu3WIFkU9D1KGxEdlQWh3IU5BN94YBbTCMPOyJTCQh32PURzvAs4eLg
n+qVYZUeK8bf2eLI7AAueKipjaGiS3g7u4bkDjtXhv5CcX0wdQpE2XzH1MCzel1y
DqEpvAtVV9QWiLeU0zheqlLFGkBIzHQv1grh74CmzMkxi+OZdUyHtWv3QPnx0jQK
zqLzhBEj5xYr1GpYqdjk3y7j+1OeHWJGEQB4OX7qSDGDB4QlDo6vx3MhB7nBMxtJ
k9keHNPjn1V9Ek/jVQnDcxICU4TLqy6PPCu2Gv0MjjsjZ5eiAR9tClwkHt4joDJq
aoKAwdanPiFeGTD3tPlg1FUHH4RkxkvTR2LSOd51DAKwUH2ss44fAMXaUhZ9pRRj
GSEYQF6x1ibcxj9lakOmC8Bt/K2FDFlUYfa3pXG0qHT9hpbF6jH7ZwwBqaexhzVr
huRBn4zNaqWaRvgRKqjsuUQ3F9W0gCEumUOIsVdN+2d66WU4t+DiCaD2NYo9U2k3
OOJnVJcJz0OM1iU0BBNro/RgAyhaLpqgsNuoLcXLlIyHY/qRq/nEJk4Y7cZCDxQp
+mP7lEDm0ccsEFQNU4w69MWwUMiNiXVYYEcHa8hUT/2Mpy07N82Hoar0+ifxL4eN
eOVj7g9YwBhLPKm4c7bLIVVBCrbff85e8yfDUWDbv1UWA82Yd6iaYi7YPZV6gsF3
NsSaSJE0aP3qSV6jVvcrz5IUd4sZk/5+9rk14IILIDAX1yqc0E9BFmSX91hXjxrj
9qGjeecLF6LnYUtDoW3k4WDdno+GVzAt+JgZ9Vu13BjiuZKQWq7+Rg31zp6shmuf
EgTr7oYbVSnGkTYd4IB2CIjoBe0/f1RfaTfEWQmdqDaF3oQARwyEaEwBzgs2QCMN
`protect END_PROTECTED
