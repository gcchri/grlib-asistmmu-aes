`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jTjSOJI4xNvud9xiaQKq3hNXQmxQTA00u6i+cjVgh3MxrX8lUZBcVHkH3VbIocAf
Ck8qa0LiR2Jj0pIOohRHcX0SAodXLxv4HL1aTfcHJkF5LJZ/7B769qoRyET1BQA0
VpPj1SBu4o4vRYfKWjM9dOY8IMZFF8KrXFyuCTKRUqQLYHTCUS/4UYp0ucVeOdoS
a7+lCEmDy1QSd7DXgiMHg5HXS+hkgDCUYgF+nzdtiI4Hk0hZ8zPviJ5Md5bHgO7E
fRB8u8JQ3XzaQflCHQAeqxvYdm4/CsinJ4nEikGufm3pb33uP3EFKCaWGedJRme5
3/L/BPUGBMiNiSiRJHe4X44u516kG8tIvcfoHWKuqjO5c0aCWPUc2oASfAPpiVl9
7k2Ie/UpppPgirPDuhEobXvIx3RGDZLV83rY//HcXqHUU6HFEffaRYCPcDtbJbQG
LLGsk6XLlhFTJqhZM1GQVzhdzolOzhO9NirgFOp296Y4Rrjo2tcleQQB14Mr6liu
OMrnMhwMUzMtj9cuTAIgNSm9sfcrmbcRUkQ3pdgPZqCQtilqxAhA8UkgnHw2yBiF
/E2yr+i4CebJEwonREAmcdzpDm06WanvS6//aZ6JodTV7/XufOMuA5IXpTjpyDpj
QTp0P5MCWZ+4yyYXn7juxDhi6+7m47OyVygwoS5hFEyjxZbmW9aWa95OEQtf3oTV
hAjPb7C/5Dl8VKrvmQK4OcsNpalnl/ECzo1Wfzz3sl/haK4DajNbMKtFwNu0HFX4
zILgUS2fFrmkiMsX9Vgy8k5HjKAeYNhwe5kDvEMS+jmW2fgKaWTpj5Bm3gwXqoP/
sn/9aCyum0uSgtgA+XwpqtKd0ixm8zNugiNdQ5Tl8bJhx9n1RedrM7Be0911LgIX
zf8AjQguuZsrsZz3TU9KH6IsE/6FCNmVVamA/O2b/CioiTn9YZDdMHgHGtd03uMM
XGNEL/KPHJENfiOzWScKybmxFTFZ3bWdv7EExX+NavdQqmzOIpKVVBPeitLiCU2x
W1tXkd0BeZ5VdSbt/04ES91hh6BjVBa7rX0NMfmavd/enLFxiwFJ1x1qL6bohl2M
aXaoed7IFTwGLV5/LZ69uTPE8/pWqM0pDQxw+RWLItEORFdL63lzggjctyBO/5sN
xbJJ08yIbg9+d6dgS+rYp/TDPRmO5M8Y/z+s/ohTH1O9ybh/WLJxLTsNkLsjED/3
x61YI0pb+4cEN5DfMK5Ypvm2OrnJUa6w1TkSSg0DJpXryaYASogkaYTh9cOFhovE
kr02q0B55SyNBa8/85gyVDdif5mvmC5ibL0dAB/FfEU8TwQ90Dj2+Za+/d2kGOWK
o4JMzFDxVQ+XJmsrxNfUtD5U/wFC320RaEwTlS6K0rzzm8RcihuwFMa04odxM5GG
1n4FDVkcN2IG33T0dkXbXV09ZCvNyepO7PGmvuckKmftP6I10wm5jMj/Sw7TZ0eF
2O4gC5XNFUdAmagGXblc+xEwIF4y7m6uUy47gsgc0YxEuP/9Oy2rUYV3E17Momc6
ZhMRjnS+n3GIAPRy4iIlLS3v9Xf+25ab5pO6ZXKJ1BMB/0n5tpZeh1S6hRbx74bv
w8v1XuqzCv/92RSlCZ3WQrS/CiOns/BfQvw4YC0b7ksD0CsjbYf9bdFfC+13oW4b
1HLEVpi3UPdhBbmWeG0Bd6dxH5BRlMXCk/NmPD3juM6ddSZFjs0uMi7rse0Vkeqm
ZJvJuVLTYFY31JfInpVTfskfnSq5vMarErXDACYqWTnDNI6c1iNjSpR3E4Kti+Js
tRcYonNngtXxay6xK/q0/LTFgnR+wMRKIRjoIayQ2EFR3cVyS0RdkOYHPpHr00Oj
NLNgM1qpbDk4p4qDd6K/iJ5/2wiq2xSRSJBJkwu/+nGyfxb9lKMovKSo54S+Fwq0
8rqqxG2uvyOcUFZ+c1Fg4Hc5b+gCe8uolcUx0TYgNpMPlmfwcDl3O6PCOljY3Yzc
wZSS5NiJ28pTQV6GRpl2jS/i8V+DVSIlmwUrRbDBPMt872osHtwLPLyCzJYVV6IK
c7s4sdG+ohRJeBAL8xr968ghLzi5mIc/Ag270/QMmhDJfrYQLXwAEqLCHHt4+CuD
tW1UsfXb8/zd0/YyZ3LnGwZCwv2cCO5gA4keuPrjcNYZU9pxkqTVy2ncRNG5CQiL
EisSL+5HO3OFJeK8wr47WVXxSGT3RDlIETXJMg2bEownhFw9cYkD1nLl8eMbNmeG
`protect END_PROTECTED
