`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cyaYXTgYTRfy17/c63qH7NcSZmTqFRTt5GEPTMPWY38QRrChhuHDJO5zynkpy/45
Gz1iBtBkJ3rT8q+n+Eo6KsGjSicO2mvmFIH0OpKK2L2gw6Ie/MnPLuuXPsFK6bv0
RgM+M00JCbbG0HlkxKoaIQi5MoQVC77lev/KSzfnBYMf/j1/ma/6fQbTKHIAm8og
l0r0Wi28W+ma6iqlGdfaLt02Gcp+ur1IZXS+IUkRCoAUKZ+/AJWOTb8kNAbmcKDv
T0jGIhvm9xi/JO6AyCYeR0TFB8tBk/Zd/CCJe6aHszZ+JMQC4FLFPnNtQHlXLZPq
YN69GJhLKvLA5vsTOgVt6FWxnkVe86VkHzbGxBVsGcvHmgFV5JRpn4CBV1SfMLg7
EIQuTDCqBNeR9j4sYW35di3tcOx2lD5TRMJWbAt5tW38nE2RQDwu4/dE0YPD85TL
cHvtipTR6kOBt9y6gCTpWBTvtQlYkrWCtPWBIUBz11kagetoUmQaJbZm2qZttX+0
W4DHxs2JlX6W958Zk2HbUqGPcvMO60L7c9+RXaZwz658mg33bl5JWMNJflaFlQU0
zwWMa7oZ0f7HWjwQ428/cO+aBoXt6FXRcAk03SxQDuYYhqsAwSXkNutL45swsLvg
igo7NJ5Kf1JYpcQut5Hq3tOvR6hSx5XJ5fg7g3mj93KRpLM8N8GDwmq528c1rQ6f
gYP+2pi+crFJQMy/EvLSG8bIFHPCIxQGXMoKMH1of+NL4RrygDN1x8CKGE1rHzSz
ERWNcxxg0ysJGxIzjwMm9Vs3L2IOquHUcScUwHV1y+CDdKYqB17SJM3dRnk4Bt5d
b8D7XmuRdx5k/SR9iB5/8F14MF/CTPTWwvqZk06/wzbtGHBsmJNMjCabjnYztL67
PF/B9IQxcHGviqJNJ7jngjnJoXOyj/0LXwKPtRtc5tMjWT1aNWfHWMO2YvCnBWwG
kQy2B7ZkjsBEdcST5CerGz3WdYMwj8njg568xlyy1tVH4FgM9WpTw1RIlpCBwjAQ
QbLpEk4anCqVUe8pyfvBUrCPW3J4JbAKVkrUeOx6h/FLo3ExHxnfucH5U1cAteah
bM8QZR3fWm3Bbss2n838XvtwfBCOajcl781E9fl5eOn/M0fI41Z50DojpqIiyXDe
ZDlaac5v+Q1v8HOslzQE+BmwHbo6bg2HRZgG018YGjOWY9kF7pbus8G2k1Z0WIIw
uke/dn+z5uPdy9i4zm5oDvoYGsa9apjpB2xs4fArLF521IbuYzx8EfuxdVwl4ijF
TSrZqXCTLnuPRagQCRITYX8NrYKnK6sUdUavDga2DLcjT5zdcoYfGnOGQCfzdWzx
r2dfkqZQMj7ClTKePlEgfVnkE9CC6WY8FCAAhOFkYt3x9IC/ziaT5TnKXIBmp6Bx
AUTmWmVQtbYHxXJARqXOojF+cgUnNkKuK7sER7V6XzC+FlVHndK/j4NaL78/m0cc
F1nX0D0XZGOzmXiGnGY06SI9cHARK538xpVQYRSAjSy8XBHGKIjWh0K8jvhZgyAv
h9F2Oz1wI5GBw2dZOBibQF+uM5jy7BZZKjoynMrcMlofsjA02KaCU1VDBVqUXWcq
vLwPR/tmZYBKWWclfEJ5x0MoNojMOcvjhYoym1QUIQm4M+q21Zn668KEZJewiJlP
tylmrbUS3BU/F8pj0m00nLCTw65RDLjBl3wx4axZEbo8kJ9fC5BxmrzxvnoydIhv
LvvHm7+iQdIOlVJJ3WBj7PixNwnVhFxWWWF2O0K9xiAiSIBZNxoEc5aQGIk3B6Ll
l0lzR+90qN02OiBLoOIs3JMCHtLQnlgmuUWDY7LXIC+pKOg3YcFi21xoZ2Tf9j6v
6V1Pidu06QwIhTGmjM4R6OpVsXlecrRziunkFNikfMF+8+YdjF5UJq60cyq+646V
6i+hLNGxQGvjTrytdUIDADI+HU4F2t1eW0ju0IfE7LDs7Go6RmN++AfRsOXhLGut
6q3TVqMx2UTm+qIqql769knIXSHvRGco2m0M0DOVqr8cfOnu2A7MUaWuNd/Rdnwi
/4x+9eTmDFx9HJMvK6se9+IHLk0yC8utSA0q1bbaDltZAPYOuJEF6tfpeqDkJ+x9
5OTongAIIU0ukoz8NUtO0ftKKf4lc+ISFLngXl0TabxR7M5t2h6w+SL5IFqNjXBx
AdVIjuIdjpcBhHDCXt6XwXfEgAzolTXy40i069D3ZzCrPN5Lu1JNYB6TNhqglj7J
ydPAZOHPONvu60YyouqnOmLCdtasAAPCzkuA1vwAPVp2w5VzqE0KegsNPFrVrJx3
nv7vrivu3drdHQcVZLDrNRgYUWHGpuMFrqQnAgvR9mV9JreQXqTlj0HChMiexnBH
edcwitslZ8mk82yYO+IvT7NHVDDzu2hXdbwNyc6FLCRNyHS/POGJlm60JjrV6EYG
R8RtEZ4kaHzaL+TRNVb/ccsAjD7v3HPpay+CrdTR4KDvZyg8OfO1+aSHBVd/psTJ
ima0nK0VX2u1Po+2e6MyAyIKv6JkXrL1vAmndgZWp4B9kL29gwBLk0RUOXS7qY/+
MxP1lDG+iBvPJfUwCcTZ+AofaR58YIbXCTVS6CQTL9Q2m5JX++574u1kuzT3wuPj
2AW7cwJ3mT+lglbzTtEoLCPlIv9ouN9FPxgGOQTPQIDeMTfLpgXJYUAGnHvjC+iN
VJjK0ZdFhFEy4jvstHrwtsAfgJ7gnxB9UcDgmpX03nt8jfWqTSMWye5wzlTeCRQK
N8OdkpOB8g0LKNx15hNW/Mg5xsDx0WXvFBO2n0wae3pAvLmyWWXIpVezfVSxpeq4
E7Ot+WUJl2/lMoxfSVG1W38PO49JPjCVrSF7Z4kUzK/ADwP7g2g8aTwDDwZ/GuzP
N6ivnpX1N3hkzYpUjly9tV+tblnGnRHotZYWF5sRQdlFsIs8kfmrufj3aigpKdIH
rXrsdphYB96Syv7P9N96w/ACbUgATcxFtyl427WlS/hzi5QzLBrI8tVBtTXHcOLt
XaCKy9AjcR2JSEsW4U4MhY5SUPyN/JvysulXwY6weoafH3u2KAfa75E2vn8gl5tc
+U7IpRTqtelIsasy8r0EF4cc6i/DkEdSwWsq4v2RJLNm56Bmh1oHV+oWrSpkRsm4
54TnhKJ2SafTu1XCR9rVJblQtTbM1X5p8fCrfX5PBp/fhO67vVoDvoTOvIW1n6YU
V+8QSGQJLEkpThhZKIwntGhFIdgFUL2lRIBl5uTvN4WZnnMmt1rfspvQKx5Rm5Hg
T/jEndup8OF0D72XUsZx9E6oadY5nK7Fkg8GSwGZJa4dCoDEHidVc6mDl90zYxB6
q5miT1keDMs6Qo5+LFjw84O7tvamL06eZs2Oj2HGuW/VZiblLJhMFKUTEUcuJE6d
O04wYY9FF2/C1dz9UYRrhdnAijEzY0OlRPxkofDVBDfsDjPFmWwL0Xkb+OI38lRg
/KtqTQDr2eOgSCA48SLQjP/yR2f7cRcm+Mk68aOo5VztDaAS6Cz4FijJfWIa9tSA
YXpZX3hQgYlwMq0faHmJEaGB2KDQfF+5vvx/kSEYxOydKwcjQfM1KlX7AqZM3A+U
awLKzmv/ImJQeonwVH3vX6ACzpSFnh4mfWQ9njBMlewP09G1VAye59K9g7opWl6v
PzJqxQc5cmZnXsJe1X1cu3kNkfcHEi8RdPurtv/Rrp4UT8xYacWaB2fH9WWrE0AP
ia5QkGBSGpVnccXbSemLx4vGZqWJoWgX1S9dWiworHdGGdjPkIm6rDgqFJl7JKF9
3fgrmEDLlyepT0WSGBmaiHxjB8ZurzNokjIPfjXf+dXYRxNCF0tcl/Jem1qNMfIZ
xMDEFwr8s/vwYuq0uJ7A2Q20VHGRMVmH66gjXLof2rjO28ZeoAcGjXRlGUPuKDyR
9hTz+dKUIIEv3tQ7a39qUd65hiixKk+/wK+iwlZHL5owr/exmya+HMHhQfVfMsRz
eYUpnHzwBnmKtf0vKCvHwSWEkAdfUlLy3rlwI+P3LA3HBm7g4iD8ODBz3BOLEHy6
6ymsp8iaEABoXHfX4XrrxexkRob6x1r1XfpqzZNM7ONhi7eoQ6YdddtZ50e5Vbb+
9iTyOvOz8KYmxHSVFQKgyrIDZPmeWJNqVz6ZgjaG2qW8NV8X13ShoZlTp2TQkdJv
y34FRxssxvCWQv8Tf1qlGfhXbCYLXFe2QjL7+iiRce4Ls0Hln/DG20o6CA6DhLHK
j/7qPmZM2Sw4ahK2TJU5FvbNauNXs9I1vQiOZ3ChXrBiWjJztmJzrFp4jOMbotiK
IcdQiCETcFyewFVRWPe9ot3n3aa6qz+JS2GEMUPhPuNkOh1SMt3Y+Oe2tIbeQwKn
1GuKL3ZSyb66kamy6n1rQ7Y3ex4wwjTKL0xEKya3WspaRm+gUKBrRy6HkcbepK7g
crj18mend4Nfa44WdcI2hgJnDpuCb25irQ1+/7PdzQKEHrvZah/KS/WNNiUWcv4v
WEPGgNZNAGqMhqbHjuZazEwj2alYxfLCz0joxNVUPfWHQjnXkinvokuX+1fBSZ08
vj85vczqUxakAiPUi85cRdaSZzi9tmxB/adm35tQ3+5qdaNKPYS+cl9uuBQ4+rcq
8cgV4D7ttkOyCgZg1Mlh+Aq8TjbKubm9d11YHeiM/kTSvpHnJqN7f1k3CFi7x2DQ
dAsmROIzzyOBMpAhi7IcVvdudFTa1nff0sVSkN5VmOHCGYuadOCxpfLaGyb8MTwG
NOF7PDnaID46aMdgCVbEtKYtzkzzIE/ug60o2MqEZQVeyXS4KKjY2e2G2zXR/4M8
BA97qK0u/auH3OAT+pmpHGaL7fyLpSFs+an5LCqdzRZIa0VyquO6Om9iOhdf6Fel
i12ptmwLeC43Nx9ROA3ZGLMYRfsRhtfL8ko3P4Y91UckqKGamhWDcZLIR1/YJrZA
QClsUnevasJTlpFe5C7co5wZxXUU5uvZ46FzW/QNvx7Zp87vYdsG+XWfmyDc9Lte
owkeGfN3VqEOvDkQ6cDmMUA/+G4HHKJ7NMMCyImoMYYiyX2hUlbnkohvQsSJMvOP
pz1NaYz/3fEGZ6m9Ezpb3bPbvb9nyAEqeKAl9nRRh7ASttinGX6dMx4lnMuzEdgw
5Q8vqDttIc0paGwblXuXJNkeussQ39ZhHfFf2zt3l522hMBoJ1no/bTj01O+okcr
JCZ5F4OahlyLjAIZm5amhW9tgFAE+He9F9Euum4tTFPO5x76MOopVQyyJpKbl5BC
eeZR5VhXPHOj5THIonshPr+jIyv5yX3QBb6w0p8dN+7AUPAOqTKsKjUYgfQDMFc8
e9fcygv3Sbsvj5cZxu3DuW3s6BYVmxV1+/UXDKM1/UYM5Q+wKGixr0EO4JI60D04
h9IaOY5ojyYtOhXLJP4bm0VbzMGq1L4lM5BK5LJ38nQCpaygWYL6L30l2RgxHNQk
nEpQy4/jndyeNAc+7LA91qxOua6KyAqYGWiNvlX6o/QTiRnvRhkhyAAFLsIaMy0i
xdygOiPGCP/0cmkWZ2dEKo0/czVt4RVyPOzDqjz9w9ftCz494KfbuoLNL7oIjRaV
ntQkiF+mjAVmUtLB7veszCsOyYW6+D1uhQ8UlFXPXgNnZ7kYbhhmxqFKEe22xGIG
JO9U3V1vDV7AkyxkhN7f12YzaZdwVWsgI4pGy0+IrdPpXDXC9G2tSdgYlU7ygHi/
HL7I7DbH1UqjH9sv02MllS/5RYf0pOrX1/2Qa2EgzAIWlnZcSis1odDENXd9+Nbg
6P1D4BPb43P+4ewrATUxPNsFHhV52CKOwdLheT4hIJyo4W3xQUpodAXaw0JqCHeW
fu5EC60o9nGggGbGHLTluwzuNQcTQEZgcjxkn4yanjLf9r4ig4bhhwyFjuv8+z4N
jIhQB7ccnsY85O1BCTvJnQXJDGbMSoeDGbhB9eOUL61eCCzd9w7HV4Yh5+3JqvGx
pu04QtA9Vkggbf6VSF2bDpWXL8Ewc8bnx04DSGPI1lltNUYlwIRxrm/NVyKH87a1
hkeFAqr3QJGaTlLI5aJ9UftWpXg2ug59yQKROoyiVP/2MBa3FNMDxNKiTqyKH/v1
ctuq4bt4K1hxN70qfpsKF4bMrqOAapgndRujiuPv3I4iECYFqbkphZHh8t4+HIaC
bzWBLi4DRdx1jKn3b1sAYVW7BsQrmcj3Xvar2r/fV33WhZ+cbVVcCtY04xB2zjRn
zJZ7oqtTQyIkydUPhV5hpYA7WhYgQnijiqJQfSBD+cVVh3d2jhPqj/3eGhEFgVSc
Ra2yMm618YRC93MTrVq1u5slCEbiTJK4SZbvRSLVOCM0nvSFSzVCmbMNndlCA7yQ
c3BwPiRCo+XYpblkcDcnRFGWZuoZsAfaQpl7J4zlQlBuP/NITzOKzuLZkhnyUTJ9
hVOFt/zGfa0/cnkU0JRejsAKnvFHT+BAaWRJ2IGKbsy2q3jBV5Bf6jnuhpU6BkhG
Ecgrw57XkODtvbgcqYVClE6GHcD/NAMJdwbsKi0zQZfFLJPWPxOGpGpgjJSpnI2F
faOhMywDaUvsOHYVsK+NGHI+htv4l4x3SZAskjz8osIDDz59COV7+u6v20Z3kl24
LH71xBAJ1SbkD0iNwq3ARR3g+EPTehmm9d3PJCNdEfhSEIZbp0L8pBdS+2yG4Ih7
Hti8lkKESfvzdaqKBaoGa+HzARwpgST/UclNBKvXJf4IO6w5jrL9C2HxP84r16LD
PpUVv46B5qywx6pzOLBpJRwe75j3pAdDuWD4qYve/JKKqNf5F5DAp7eGgN1SKLwC
glcsMB0P+u9ZUfqMdIl3MCZCRInOod9FU1TgIS2MueLsWmaW7ih26SRtw7si4wGL
kgc8pK2A+m9XIxcUGfnqUOZ7B9ch7qy9iqhT0K3x2g12FDeEG0jYQttPzOykTaJe
tj5PGyGKyc5gW70rrWGHZOqQzjA3ePpOILbxPfzaSh8nsigi0qoyff4JVWy9+pUz
ujGVuMUqiOiupmgcptl9SSjm9n6YGlHaUjRmXSG4Kh5Ga40EbXzahvhBUvLhHION
QUb8PpJhjpFrCL3OgfgRAu6oFLAtkWa8vGrVz1B1oRhdFUwtMAcpJIQgXYKxBDq0
Fel9DuFk0fiX6OVOjG9MISKVTtIx2PM6WqRj3jAMzhKlk8FzhB7u/jKSI9u/ZCU+
nkULV3BFdeOyf7/SDe7dwYNo5kvd3vfY8YzdRFCilscxs62UapXF+ZRip3OrWN+4
Ep1tCzY6XiO3bbFV8e1BvxqKAzS50eCybbMP9GXasZNmlr2nCnCsI794yEtUVhoL
UHwJhvXtDFeLuvEbGDth7AuJX3s/ViEZcKTKiPQeoMjQoZw/mRA2dIEPOl+Ulo3a
faF634QrbZupQGkygmeWVTXPSpJUmDBFI+/R4/5IjkxPPelvptr6IViFj4SaryD9
/lLrMSztaXgd6JBsF0qgsBskzwwsbQ+KO56tSJn84LcvQoB2ocyxzWKoOM0uqi0S
68pDuYoPCxFae/9YbQ7964iPmfAcF2ngcMUEZSgpAuasma7uRlyJqMEXN6VDFAUw
xKoJVO3vB9Hiqr+hTcFPQFyU/EHO7lIa8CMiU4WlKHT3ANlkM3S9HSK+FQXZLPAp
dmP/7Ie9ixTvSveY8ARCpA5/g9wN3FsRFdwFv7eBiMfraMd+uBvFdu4a3j3rzj9E
E3FXI4KVnb8H/FHzVHGMiULJ8GuOZ0NYZ5sQChbNJOwYTROErAOEMAcw7/zfO1Lo
67RbHThORR/zhl7ih5tpaXBmQgeP8QGuYzYA3YG/06OghAq/Zh+Hc/WOe6SUv5bv
nf5KlKIqbmUVXzlwY4EGMSU0DNJlCCYIS4lw6BmX70QTICkJuFN5vy95j6NDpafs
3FxGBNc1YTDlZWt/S1whkURGq1coOGl3H+M98rqRpG9LHPBxp+q+M1ukbrBkiDDH
e/BSbmVXecENV5lbif6lBi8MthH9zzoiKSFhwDfEFdbIan5LU1Ym+He6O5RF8BSB
Jj1/lIca60bKhFebHSgYQcmZ/ssWVtGdlZhxHXZd0Uf5WmgB98oJVFdh7WGkIDoj
ggsDolp2SiqcQF3lXQl1FujPcg9iteoCy+mYcpQSbLUGYgGRVOoz4Guxu7p3b5+n
zkWImA5+EDakgCEIp+Fw9k9ak1ir4f4KzKOccYihC7P3YWqmSXkkJllTxz60TPGT
A9u35asX5eL/0Lws83S+/gSFYBHyEdCz8vOcfy9P7z2zzzvjH7CKtEVQAk0RUrgc
VzRuqzeGMkhuhXn5j5mzbT7OrRza+AJpHxG/CiIDPyPb8hncVF6/nEJpEk9P1jnH
v1OlqIKSpdt9Q4HrYgP/MBj9OG52MdaokC8P0/10E+K8IqRPCuIwwvkBf/6QGvz4
wSwGgWoEAf/uXN5fmeG1yGwPqHjF/p7u/X6K3OJTbG9sWcuayFGeNhAFTor622MD
bXhC2SDd1BdpbACWA0Tqr1tbkh8xEqiqkrHgVTT6Sp989x1wLfX5GzADdbPkCtjj
pDPT1L5IYg0p40ywfEwnoTumngQzu+wOkUgRI0WZmQLlDGZzWCPVfIUKhwa4vUD3
KaY99t6SmHIcAMD3ylydYL/CVJWdIX75mOarIh0WdTnDJNSJ/jCvYkPxNHvBD8KH
xL1onra3fDx1507OYc+uG2bCWR0lUMfMto3xEySuutPVau1r912SJb19/7ZX1mZh
wjO15SFStoM6OwktCG73pBY87oxuohlxlU5j3nNWMy1R63TZ7L8iFWSO8nvlgXLd
Wc+M/BxTYFsmGQH7TPVgpNt5SZkMT5rPAZvw5YkWFvMvcSRJ/XqEWNTX22rinz/R
6+W/TcLTw2OAPOBgRo8i2nFcjpbDgIgw9hhEuqGY9nKYe3eL2L/+DH5LEJ3/41Nr
90Y3Hq1Wf4dJhNYB93QY8icguWj6I3PFatYSd3AJ5plE6cAaQhdil/P0N4bLMVKl
9X8Gljr6o7dIGsRvCB7lNw8ysM1Az89kIB/w1e287C5RfIESaj4fEYwtl7ANVk1E
vctQdGViRSZehD0uQbS9MJ8zQtmfsYia7mBJ9htnT8St+jR2nVytikkoDkxH3OI3
CK12c4Pbxcr2Pqqf5yROXs7NA0xlYN950c7Im1gkqWYhfbGnj6lZlLq+EQUtso90
+vV6ANh7gqJ7VNRiB1QDRrk9lixUmhs9JY/eUg+f6g8EHuCdKikz8VIwPx72UQSz
NYEE8rDhuCjcDxNHLWsoeJ/wjglgGmrCaFW/PCkDzoYVp1P5Vh44/mt9lTpPxcwp
tP6rmFwBIADwDrWv+44gX5V+LXlTScN99Yxe6iDDj9oWPSWb/itALlaFopE7GArS
x2W4JaN2Zk5cIz+bf577Sgpfho7U53jU4FY4PP70iPywKzRAFIPlHIul/szpf8Bb
nxD0qkel4At8Bhr+WOB0Arq5I8b5CK2F63GLk/ZlTD3jaM2fcQMr8Yq+bS1t42Rj
OotXD3CIzzOsqia0Drb+npe/Fv5hFHt6G0yXyVvzp8PyN+kG8JOoWc+6Twa5CJDg
h80mXTjH2pcKeiBPlMVp5znm54boGEKhQK4cJuST7p3HlfU16mM22rkFvNGkFSJg
BhT+eTH+rg1q7LmZl7H3a1rdXhKYdtifPDxe8QSjQk5nY4Cne4gQalDw0dEj4FJs
uuTsECBzE34jmJMDw65jXc5EYHdfmYUnVo1eIe1rdaHdxhMggy6HkHmk/PAYz5r2
xX/BY1sCk1vB08vkJd3vpxyiEfli7hizM1rumLnmZUyWU6GltaXU/yadwqZkMMhW
8by50V2Hng73ubw7pttbWlvMOm/UGqqiU/f5OJUU4HIwhuxKnhL0rLLeelIBm9Pz
ul+SOOvK4Q+EazMzq18S6a+S5AbzGdaf2byjN6iQ7rR9Tw50djzOZXtqUy0ZdZ23
VtIE+K/LRfTQ14jvk710vArRBLS1v+QUxxWobs5SNMLffpCS53X675UtsSFeU4Ay
RvEzkcp/JxLP/9csNSz69syzNY1WRYcrRaVnE+6Zb/inmeVNc02dTENWgfq+JTpl
yCG9jreJpmmZrQUhgicHCVR5YD4hqCajXrnBcQbg6zqs5YoFWAr0lcsWJ9Xq4i5i
tOXIICxJpwu4ZNYTUCq8knNEnR1aGCvRH9tRUvNdM9AxWDC2FQP5u0VaZBGJ7Qqm
ozH1vH/4zq5hIolFnqSQrRmV8PzKHxZm7e77B/du4HlMwOTnPBdRmlxH3Hzn9YzW
0OPvL0qtQGnTC5Oyc4OWkgzg1bU84YhlvXcjk7XX7L1hgzxmbfUAWcFoKVig3jcb
sVgTiVD7/f/hWBi4FkPB798yA+LRIjLxFWmVE/zuTzIX8EGumS6KGJUSlQ/jt/Xx
zcGfhHHH/9bzu4X+pMME5IMg1JWUHcvMatwWknahriCjgURNuGWNYe1d9WZvuWGc
sd8d4xCV0YxgvJfwgOI99roMCsZ9efQsFQVaPMjMzFMyi8DbIDacI9eGSm7RbOT7
SZXKl+wKF/uJP175YVxKWQPRm0fABBDOB2xCpx4IGmT/3fXhalYmI3NpgIsGr5hP
H+WrzN4zltG83JlLV3OIvzufRKZ2F+gBFJ2hCFc7eOw/xt41+bfvsRGhdhUYkuuP
IrpOVhYb6+knLW4rRXo2NX1aBZFchwZgJro/+MaZ4DPplWZiMaxSv+2WFz0U3gsX
qzddUnS+BHEmDAeJIZYIajW59+P4o5jZ3XFPYRuXC4RSLcQSiSVhzY+IFu5lpl7i
iig+WaonXMVJjzi98k8CuyHcBVJPhbsWV/ehhiXHZNFW3F8RF5egoth60aqz8gL/
GniHTuQyrl6MXMOXeWc9fF66DxBnsrBsOZ+WyUg6uvNdLJ0+XH16YguyZlAKx4n5
cbkn/HxkjxyrTU5XWSqzHzs5EwSbB+8Ous6dia21CsJUTXXT8iJ2O/rZ2sTCckuL
FpBX2cRHsVeySwqfZEcJXGGs1F++vzJuHU4Vp/nWlQ+NkS+RHhA2a8V0/IiPpG5W
8utekiAReLQL7ki1WbElOzFt2WI8nVwBrPpIjuvNG1dy+vNPjd9Opy8HiPW3AoXd
AvH3jFSh6GifxQUTgWNos4WL28p4iRG4XFwD23OXeTzy4nka7559kD7sJcWiR7qW
6j42bMfNY3AUp2Lf512OM5szLCZ6AdnaYJgp/ghqAUGdzFe5HDQPiaf1rxoc018D
ShAUTnuCpoXj/7ehQOwRVtjOKEKImjPfSbeknMxJie6Nl3t5QxB64HaXPQmqFxOk
kgwNcvYwub5KUHGUTzl7uoi6RlU4EvL1kNaPuG7uO4u/tM/C4OhErfMVEPLNU39I
nlK57Tr+JfQRjWafJsb9t44AmJSCj8sxkUjio2sN65+eQHX88I4+hWXHubMqXiEI
AyneVuM46a14SiWbv03IFnO6ONmXpzGosCzL6x1WeX0AuvlhNpOkfisnWm5qBRmk
9gBSmK17r1jVsIduTPhc91JFzx/3XZ6GMTQjJT81e2fhLX28H/WgsSCPlc2zv4UN
qjyukKWVzP8CklTFHYZUIQYkfyrtA9+5uWWIlnUKxEF/AulE+tvJo6oKFw0KkZia
sodnPsPSfMpqlp5PJIVK+agknbxnzvNlXg302X/Zf/vUS9vYeC4tFVcrFSu8GcDc
jK5A2Mt3wbIXxCTrmqNiVlPsaXikZra6AC8P8XSZiPwtfnU63sib/6k2Sluybfb+
ymphZAH3zsE6gz0W5U5FLLT+XpUjhdjzgXomCNBxymklqJHXOPflMtbErPH/hBPY
Hc54jIiBYL6A15aUbU1IQEKFhnwp2s7XNsFQvHd3H59Rh3ctgN6gQDniMsg/sMub
ujgOYTNpJcS5Y2D2rBi9rH51rx3k0gfv4ZLMoLU7LN3eL7W+sTvDBtMEWePLF3Uf
1PTtyVeomjqi2h0jZsbswgBAnjpo1B9D8OJKdjfOnrBwuRjz49hLKfpjKNuSDBGJ
RJPHQuKupIp+nL8rLUqq1bYXkH6JUuZJcB+FoIqVQ8nT4u+7L7Ehzvpt07gb11fs
f04p4iB9kFLDInc2ztWmKQ1Bu1y6YK0cMWJulVmQuv2cIz9NXDwlbwAyiduW4oMl
nD+YKC7ZqwtkoPEiYrzeE8CVzqkg1IpiRbCtszZSiswGJJyIol1WLciONw30UwJQ
Gty8KGeFzm+x9TAbZEKeF1NBDehZ4p4nL/CaGx3kSi9lNofegyFIx9JHGRMIqz91
zxkvF7hywXWBmTjDFbsXnS7aL0ImxseFK1xD7CFM8AhklArzAzZwzbbjgv+YQuL0
0pv1kK6Wy8uhVmEi1ir1mcoK3AX7FuoYbhkxUWC0lCGBetUlxQugr5LPQF96rqLU
Jf049JmgqHAKFjR6gAhwC7GOd3aI4ua8e4oAF4xAkW2LlGoeKnMYCIdGcC7OfgUL
jlAVDcyFZ+PSQxoJu1ZEvNVU7lOWWZNLqAVltPMaBzy7P+Saohj44slTs4XtmfBG
k+0e8UPyyPkNw7CnaTbwrS5DQfBlTJFD9duFzmh9uX+FX3rf/CDxmTWEY70B0ixL
5B1BNkiR11Qxqq8dZCuMsoPmkZ5lcLwvUpQVkYApkSgzmwoXYwSayfvLUMSetARz
KUkZAcfMNOlRmKsU4gZZAKVZStQhMqvWPctZ6vY32yE=
`protect END_PROTECTED
