`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xN9GByICCfvb9EHLH2RTzphmkjigkY5BbB1GrwGajWhrI9+jWlYMVucqcnCd0caK
q7J2zeZ1yRxfCcUK5KFlUEWiKsVFv95qga9Xvxvvu8mGSoB7bSKigmh0ClqXkk8u
7YCHmm73lA2bK2xZ0IQZR0jrcOqeqjBfiyLZAAewfbXH/5fmA/R2fBGPd8+2SERP
+2z2zI6KR4J0uLk3GVnXeKassEHsiidgkoEoRWJIR8++dw8IXPgsYgKkXxqeae41
3OQa+wf+uAyyZ8aP6j6B0FwmG2HDMxdBOXWPz26y5xgv617wDA8v3MHVpFEeHT3Y
GU1jRnoHz9DixHF/sMoIIFQsgfvmEj2Q4eN6oNkRp3kxWZkhgWcB+31uHyIKN/jy
StO6iTdPSBEPS/FJV8Gx2A==
`protect END_PROTECTED
