`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
czHdXxBSrDOEiL7dX/+2H+O2WskSATfRkqBqMhEF+ZS76QX15wzuPopJ59Yp8XaZ
DtFUHYl55M6jgvQQKAu0ExFbHsu0TM54tJUTEb1vCF1EGI/LjBTin/Zb+ur3Lfc0
nUWJNzYOfVGN/tWBJaZ6JD562v7hXFBWbgkKBeat8gt8rU4sIuIaObO9MVBG6y6t
VkIXJe2NUvbZAU9u1RNLXLyGzZt55Buz7kmzapuCq5puk2mFhag7xY7mRjOWy9ye
8Uc8VYlU+X7VIqq8Azcmy2xZKDSiUOwVc2FWwHQGfYUBfkHje+c83JHqwzasK4Rj
GKX50nIyFgmGkRljelKvlJEQ5yyG+Q+fmHJQ8A0aseTJjJOyPxGWtWAwENDQZq0U
csf6+hr0DYp8galbT0ppyqAj15KVlQqO3+UtT1Y8gKHAQafzWF+vpu5aUxnbfNQH
ibZp0dYcR2vn78jCejFShmYR1FVWS85pi9QsgqWBtbQUySfFlqBxne2sH4aZnPAZ
6gARXKNZq7HefRDkS2DGImGhWVy2/BSPnmvUirJWSrXmFKx+LVMBo5dd0t8c5sbV
8fMEiD/AJ48yfBeYRcQlVho+UK4gxXxkZWVhfWoRkAYr/26EIMYBH4VD2sDRMKsq
WdISZQMJtwTfDRIKTekTp+I0cMDeK17rg5uIt5pCOutqyiRDOnFo80Yq/dXuH6eb
SuzMiAWVoPMo/JzLFfwvaBQ5jztvr8ZsyaHKp4DUpsQcs5pTgzWiZO3ybzEfI1NU
u0wGkySQSDw7toF8CewG553bL6Zcvl/tWJIvK9ExK7reCU9xQkgRg4Oq9Xi0vIEO
8Z0H5kEdB/S5WXTSJwkw2SaHwqWiTnb02l55u6hERTUt7eko3IiKkNSF4bkvlxh5
3P31d4vMWWdHwACjfqOJuA==
`protect END_PROTECTED
