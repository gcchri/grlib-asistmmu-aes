`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G0hA5crBlxPdMAhHmL2WKuEdfJtuXvOwvg1L3V/3SEPskt6g54NZWPS7AjrfCM74
FMr9LWxjhx8+0IdASmEqPHMVL6ovM+J8dEmP6yOKUenHQPS+LgnBdQwmqMpH9qTC
p2xy9tMM9HsVzfuZMHqDVNVJBLwgenbinYElr9jswqd9buU59HsyDE7cLn5Cax5r
VfOCeMYytc46ewuC6mGhSDqV7dQiwCDD2dcNnMIfyB0V0pSic8JEDGImGFQYx5gU
X1VN9AiNA++Nr9E36AqqKK/DhgJhxqEhm8WKLTDy9xkWuA9SdKePnZmleW8/fOEY
2h1TmhZbfoDEyatbS51GnI0LCCgs09ZUxkf7z9CWC9RoNj4Mr/Qw68ErCoxF8Ewh
3UlFgp5chOuOKN4+4bDObEeMD8xUSCWkClKxcFrERFVFp3IvPgcBU0sKQWfKCINZ
yjsKwgZa+qAbxTzggSok0D91kg1h4mTHG7hxv+c4JtVagf4/kB65CCm7mFtRbQSX
2ygyG7a57vqUIQcnK/T+qPuOn2evwfhUt+I9QVhGu4EwX7lAUkn2iEXy7t7iuzcD
SknmdXPD+GfpQz1dVXKHpvL3jKvSr4KDh9Tkn6zSRZmi6eqcklUxq94TTjiCPLL7
vu3u51Whs8nnHpP1kRGw2f5etQEXo2fuGKsgeqsswg4JzaYO954OCoLDos5DVPcf
I1iTquE4+JsVZM+geBxXtqpdB9Wth5ogSSpCHBa83KXiuQ0UUiBcV2VWjmATXzuU
5kOHtDgiAHEEV3b+zoUODWxekrfAZsfaB3GKVhQsl3L+P6xpH/L9l6na1oSzB71q
Y538FMCTql0TECDRghaQyK6uFN/iPBTOpr2W/ef3rZ1qm1fpMVzhoRG1rTIfbeBl
y9DVOoM3HM/E6FrCmtv4ItBPpAedPCP0zWaCNRj0cxAy4JeW/6lwGvLheEZg95/V
KBP47xB5gPzPk7fmVRZrdg==
`protect END_PROTECTED
