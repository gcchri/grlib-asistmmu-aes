`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SB387rysr35cdaj7TJ1uTdFX6ImVirK+GjQQTZx5jcvtADEeqwf5CLWmWqii1wTx
JicnqIA1FHdmhRzpKOT7FDIinBcqAhp1NjTKq057MYCXUXa/Zn8oAf+mmPeELM3g
Fj5uj9ZOZ8Ra7Ux6HwbuBYL+Yn49klQr8Ievu+hciHWxhiiB2qTOqFbEi117dzRb
4XDd1l6ShQjm1nO+gfIWqbH8v0EYIxTdAaxUdWGHjv95hvEk7/IDbul6wfRCrzKl
txvDKqKEH2qGjr/KTPdW4rNQaExFYYWtRvcZtQWDm3xIZSwerrWA8Kqmia7dAOMm
wtmNspzt2EA5zdjDGP8uTo8C1zRH7W9QGg/tZ9AUzBa9cdPkWtJvXNj1DHnt3TzR
R6OgngY8q9occLkiK7bMoB9r0QIVYmiY5Qxb6nKtfC7LnCwha/lXXafQXou3Rk8u
7Lwh/MSr1B7tLCx634BPkBATIcYDgeRANyB1oB6QzWP2xgi+KLaDL01UkGR3fFKD
74Pr9M2tXcKxrpL6QpwjEXCiGVj+gngcH75AUpQzLjAnhehU+bKVwAWjH+WGAkNZ
hX8yKz25CVkLQBWO4RfXu35ykRROJA4HSQB1qf949nNu6nw+sYs1WI4qFr75v7d6
mkdNkXVLfXJihFnkkp6wlFCXtRLXjlrHIkaltZCl8aCiUHSbmzNunxaaHq4UDmqI
D77EqUXr8arNHKNa2u8LjYzsLnwv1f3QIVAatu14M/4TNa1mN8aNKdpFzci6g2K4
/BmEKB+AYf00dpHt1EH77pL7U2Gr1Yu321rPPHaX6I4CZpsxYES+RG82v2O45DVk
6kqpnhrFfJpSg2TClDNAx35L/72dLh9FdGWpE9udZf9T+pujjL11/c/d9iiQVdHi
XfOjvmnmC/nSNodxFUuyDVev2DrdOkDEzdZzCIVM48pNT1G1Qi41WYikqWDDWyvm
KvIsmJKYjnZj1C71ZXtNk4C4iTMY2+d9yhWqPhMP/E9J4lIzMQagoRdYqvmiY7/l
D2KnY9bbarCnkIpFljQqae1/K6a6WNDcnglzJ8K/QjES9tg/Rl8wqSoNdeAQ0jWB
ZdRGfMDGZH9WsAyafQwaOQ32sSQdWMpUZjS8Rdrd3jG0RPrZ/juU5ha/JS53Lskd
VqWYHV6YnDWsizU6nV1mSeabrCJKG/CusGW4wJQH8ZiJ0Np60x3/1nqeX+phgXsp
+Z9gQADZezKs4g6MN0BrUDk3nMiKiW9pvDSFy6HGEhX1Y84BPLcbaDwUD77c4YjY
90Jg0e6FgU9e2EHpdxZIg3r7aAT8yVywbpNPfh9ox8BJDzIsWRlApvWNl78nfmpv
PYWtKxVk4NzyPQSqU/jmeikHrhskM1lt6gqmdRwNePxEtqViPY9cPgoe7r4j6Ezb
drfB6EyvNrmUoWaG3n6tUtY2YdA31qmrTSFt1D36v5i9PNHbSMz/OvbR4Fjg51zD
3kSM5Y8nspLQuBqh7Yosy162shoeRk/yruABxU7IjJvnLLxfmfRMwOdax+/p+oNg
GBCc6FCGO71fhjn0kQ0xIOQ47QVC/448aqHftWNia1KneePZVZXKjEPRPRjOTfNz
E36Y8XLaL07k6xSnW/oDt7Wr/DKiFUDIrNeWuyR0ScEny5k/QJTe0aoIi7XkAbCV
N2HQ6oNv5SrfNKCW/bAgIuBQzEZOpg5SjpqoXsaJXa8Fe3Waklqj4Xa6c1h69Lfh
UrYL+ixbOv060W7eeHa+3wE0mqrBuphn+X8QWxhMCAm/bu3n6VFbDDatzOz6Kg0B
dcHEkWe7K1uRnscsKpAqH5A44bXMIfix+8ZjzfHGoVncJLzNsshgwIBE9D9Vt+mG
WwMhEKPFHCMJlriJbDsWtC44cvXQVpcFXzlug5tKDrizfUrQjPpcsGZWqCAgl5MK
HDCzPoAy5SOXuXuFcYaQxJj6gLgUx1IR6XHBF+87+mixuSzcSgln9vEEusnB5yaw
0NLXIMG+SvqexTr/rd1gp7PbqO06L8Zd3AD4fpR2yptAWU85jE8WVi4b6wqZcDvL
/z2zE+x1ZacvomqZ77ysX+K4qrGBVXIAhYq160UJLIrUw/DYm3g8W0a/F3aiJRx0
o3UH9k+EzGosooVGAiYtORPeZBHKQK1OsdMdrcjgzuaeJ4d1pynt1JWAUqUjyAfm
dgqsHR0ft0sJcYts5kD4ULXNEMe1icy3J85unK39eU0Yb1Y2ZyAoQo9nOXYBTxrq
kLL51xGoB/CUOH+6f/4iCfqr2uSmjHCv1gCR2s8hx6ERrtPWwGXQG4/ZDe/WNErd
F2Dlqb237ER2R3r1x8NX1FNXGZ6D+OeYRjS+50yowsFAkKxRR/dZOb8wcB4cc7Fx
/+GXl4QNtPs/2j3Wm3ULky127SWMDMokRnkvgCFHaLFEbVFHyKCtbmC8PDh08hPE
ozI3Q1I6/FvSN5WC+PiPuRI7Qo4zeLV3ZZkqUH0QS9mLf6DkEEoJG3gkNXI5o6aU
89Fb1SCI5jLyzwc18IE011DzpiZj0PmJhHkZiQmE3V2+MXiOS6EoQiFE0AHeQWLZ
U9FFqYkhzVY45du6zKhe0+VSkoGeHb/IKkk9RGs2YYb6Wyz8M9LMByqWcKckkEGz
gU2bUQrlHTFzw1LFzL/Iexg/xYTwoeKo2JxcW5j0MDvmYxl0qk6wgQNj8ORKuGTJ
BXn+0ZlWSdjHuGZ6XPfaXhgC1+cnEt8kCdGXr06p00uWn1X4siWxZpB0WNOAJ/pN
BjZnyHgNqF5OQ9abp4xzIBxyyZROb2WaNq/VefXSvpzvqh9Wr1CHehkbh3mVzyak
cIWpPWDrQ+lgUdkQDPGHHXfJkbmQKblHHTmbvXg7pk8QKGDA082TUjcZNnrb2sVi
Du3s2OQFmXyO7iAHy2LICequqCRYEJpO9T9p76DzpShijvK+bhVRj/kEqN8VNvBi
gDQtBQfPw2OzzTXwjI58/8g2Bmrs2G+UZIe+ZFk2IkaRc63oRIWCRWBb1pgKuNbu
nm2yy1oTIeH176kehX+jK4okYl3DzYnXWHzqj5N+F6qYVt1lUa/m8e5Omdd+bZAO
5REU4Oej/1C7H/fyxIZ3QWS/+jy0rjK1WpiSY4m8h4z2GApH0n9z4up8BWW7d4Ht
/BMm7XSimyPardOXZCcJuwuGy2DMZ6cAlGbRQsQneE6jKNRvH1aKl0mnKRP5Q9vW
yFPRu5ryBL6YhkdL+N29B7RQKgHwk08dv1ro9Qou4OAO+Sqz80x6obQnOxSTLq/u
ezXUfFsIk7wAXMB8UA4epvd9srTBVsVSxKn4IF79Nz6gGk0wAePzBwCxqcmpNV4J
jvNDMDFxZsSdLBQXRK8oFkTDa7mpQFb4pGz37jr/EbPAim4CpJhvHeltwX42Tlyf
RC3w3mUsgNFoZ1sNGEdXhk6uNb3yh6yb4gCt1uwDCSaSvrZo7eo1XGjsjKQXLYEJ
h/z2QtHVhH2eJ1PWJYQxls6419IkYXImUm6T4liNT1GGD49nfYXyDvweNGhHTRgP
q/zAskzjEyd1kaIKpw9jSiR+abFdlZstN7kCGWZqJbzvZS+FtLBlrhuYDhoaXEln
tToOANg57GDZlsRWhrcFX9bBpwjgQwGoIb0T8qQeNV7cF8Ej3sa5rR3AUXZEBWvn
ptbL/jx03hdnH1wo6FD4f9TYc2pjq79R9+b5lObtsEet5KPlDl5XJcD7HNAgMkV4
X5dAWSd4StNOlQPsyUjS3MRZ7XdB9EUUhHv2QV7HgpccfJab7QF5UVisLgtSsfaX
iSOSA5DZtRy+r3eB9/CCZjtK27i8MwmustJ5XneldwCeIj0N+C38fFoZh1poVp30
+NrUn0MQyMafSiDd1DlzIvDdge180GweKPraw3Annt/I7oWRJPR6/Ky/7cF8vSfX
ee7humFcgeDy6hmNCRgxi2Q923Kpbcw82GW3uS3OdjjH9dyhown7CasGXgrUWlCs
3irporvocAyylAuy2+NQ/v1Mf45vKfuoRyTYQvoJ1Z/KXiYgPsHA6nXOvJRU4Wzq
Ulv+gED7lrmRShr6XPVCZbEvFkWGlKwNm5iS+mQWI16oEAfhdEnx6YzqHKS+Lwq/
PT/aLZwWSbMcSgEcbtnV9e4NioExzwctWQ+dJsDCbyRaw1IMNwJ3v39RFAzdofrY
ms2H6OoQCB4aA/WoFeFnzUJN6ydFzwTbkV4ZxaZx+YTMbJJ3QnPOtj84mtXI6rBj
N48LmLN3fmq5ejLu35iYhyBZQv2N50M3Id4Z3Dtsf2AYc4lNMoPvm8uDYouxiMTB
kWFVfjdcpVQ/UV4tzKYjs/mkONaOF/2Z42wfVUmZstJtxJyQmQenXUiYHnUJxZK2
ozAwx5gOX48/qxwmqPA2YLGyW4YUNnKRMY1eQMRAWl04QVDzeTUf9tU83/MsMCNt
2qjyXrRhNs4Wb6N6jCekd5lcVZLAeKTO5SO4IjDcTZm9ID2z8kZdh1d8+i0HXxSg
RzK/qvPjeWBwF8FfXZ5YxgdImbPaBOyjnLBcCGAyfAsUdstmwmfc0YYfWD48f6oE
eTtRui/4uEIRPEjRcrKMOo3r0ssnJoCRuYML63uKPo+QYXPldw1StnAzugChI6t1
jUx62oyPWJofdC/ffxiQ8QVYGeB4GcdTIkcrAVMbZS0N50qnvpWBrvnDaE3F5oP9
r8f83HjPAYX3fp3rQZ3iH09S8k48pQMXlt46as/2cTX/XGbCX/swxVbUJUDWbdM1
tCBeW0jJ5eUGqpRpGphfvPCc1kidB9Sb4Jokojt6NAECOye4qHhIrH58i7Djituf
TqL0gLTpA/u1zgorOsh4qLC6ZKNPJruJCqgFPErFn4bJ0n+EIZew8JjUGziBibHT
ZRlwBkdVjPa0rkLViY+O6qtO4P1ysCLtYXKhrM8BerlqzyXILkY3PnZ5F87WlwO8
VL3B8RJulwFejHze4n4Af99yvkZ3Q0GCZPvxvD3Ew5cfTBkC4UDwC/7nQIu90Vv8
tp604gO/sfwVzkVjeemUrzFF3AJnIT2o2Z9odzm50fLyUKSUXlAXsuT8Taveh3tX
sPc9sVDJ/xjEt2IARxVIv/4ZPGppwEe42IN0MhRwDlkud7QppPY/lbQPqdRmZhMe
04AJraxBsa7w0xRjbbkX1neyQazbffMnIBgQu6Rn5HstosDzoJ8XoszVooHQVSKB
r0e8BSWRVwH69LSULuOHjY3+2Va5hIrnKIcWC0wVin5e96IcxIo8mS4a77A/80p3
yndZewCAPtAMZ/TxxiMc9nyEkSHbI21ja77m5BQ5WDmq64AZHPzV8fYuZO6s68PP
5rp06ETSo4nJawGHQGPKN2GPzGS8CcyLD42WLgK/SyIbk+dCRoj2GXVX5bu6oRex
UL5igQwfZXCo3L1UlWS9OkfGvxJaWWCvjoUPqh21Ioc6UE7amf1pwfwvBJFMHW2F
jV1/l5F7agvbLqNZNd9VAHDKwNd6kFeS5uJuB3uCBorz66ULdrztbIZlqX8FPlG7
82sw1T6kcEyFpi+69MfvguAa+hfDH1pqzT21AaRZ+RqURMN93HfknZr6I4EhqfYC
qOjadHsVhnQeu0520aUSuP2MRWALcCZggTuTMsB2aC0iCUJ+uZuRu5wJFWJ811A/
wBxhgQGgBSxHNaaYDeg8t/VyAYvsfL7PgjpQWcynFjrKi7oVXthVehAbbHYeoTSC
wWOQhk5mMoes/gBfDB3RY2AS6ockPdO88SmgqEdKlyk1MzE7hDi6pDP0P6ugLZcj
QA6YxlHYbqpZUlm3C+dM12EL7dKJmaTUIB2CBzoAhEKr+GEqwIRVU8ecnli+y+ic
/2AB+w9ZmGkuY1xrzx9y1EMs3N9dxLxsaRdZVwYk8fnchs8+V5xq55JpRbqLLJLk
7EwRIkuqslRDNRgjqAZPRvVAtZtIziNVicossiKFmYyJkW0qPgWo32HAewwv1OCi
OM+X3FZYFJHUG/xi4gG8aIPFlL0u09y2B9crqP529pGRdSYmFRowFoWoDjfkyj0U
79TB0t3zYV1cQor6a1jcMkdUrxRPt79KBiIYB4xX2hgMPKzMjpCnN5RFKp/cQ7Da
gapmyN93uB1TAcMUgDKNiQsISpAAWH3YDdYOA8sUKUKGN9ZAxYdjsJ5OUd1pPE8c
wfWhnXGRnwSG6tWiA+4ITw2AwxHs2blWn3ZHmYK8sJ3drhP2NZKRRur9rWERFCCh
KkqZLXPLXKtZ7QF4TD6rQLGP6MunHrxeDDL4BpMKDNbhPeexgiZn07113RAfniQe
z5kJw11f0Ke+521nzjmYI+Bb43GhVqpsiOl+1IDFN3CyH+UwRkYNLsKSiJpVPjno
p2Y8paiwlzqLORWxVbtlWYoxoWhzRJvSfK1NyF8PV5O9fzPjcgh6epNVeSBU+A0X
Jf9S4ibaa9pP6wlWkhE1vaqPolfpRK6aVk4LESI/fXrlr7K5Xnnfgh2Sk4oso6yA
NHYSuqLfHrrBgLfGL9hsAfp/zeaVEHxTM2V+MZ+FynWi3jTyyfUe5moqIerpUI6l
lJi/euCrM0ZF76yJ94VVNnFuwzCG5igT0E67JuBPzvdhixDErodeZ4EZkPJw+xcL
2j97Sg38i+tn9bXaAbcyp9cK/nUWis1iDq/IJdNJmqgTfmwjCv2KEdj/lI6oUXoX
9A/fGmIc44qYDkGxFegcAjQXac5/8BmmV5itEMdHk+J+Phim9PzLAQYhlKYxgrdq
bpJy2fQUQMCdCagamrxH8+V+jI+IhozCqFpMXnS3MgFdzO8LY2Mt5BVjblaEldqf
z11JP9i3gMZ5LH4pU0/rB5VgJxdPun8EB/YRAXMEIZq2cBBISpF7nJZGHP3dSgLT
Xlpgtjuo0oCrMImPdEbIDky2V4UYxjRfPhfvIeuEhAznoxYrDEeRmm6ujC9nisDT
z3WAK255hSTIALTfTJiYKwn7UefsotYw5CBO+r5W1+vXTFKr/EPyVn5betnrO6Ik
KEWLpkfFNvmdG9SlZdjy0VKeeuMhaygAAMt6PMlQ2vOYSXNtkQJgrQNvmqMEJbqF
0twwRLxcql1YoOwiUBCrQ3ADq6Ivvet+BB7rqvww+n95Brgrluu9jUAAtQvtvxTd
Q11clM/oc9x+uspMWWdj9s3S5hCRa8dPHvcdNna5YDufK4sNLzedwCz9q/I8ATEf
TpLYAV8x+r5w4V2JSf7j9Bt3IAAq7SAbfFtoVYd2i3y051kC8O9sNIk6FYUZD4QP
o/UH0VdJ/jrb+tE7a4qwOvWmU/8FdKE5co75BOaZybBSN+n/0MjrdEHcGE8tcFLy
SlWGTIO7ifAOSnNzWusiAkHfHg/i4RLH5cND5HXCb3DI4DXazWQOTsiEmP6dgN4M
6BW2zJu7zB3mMZuU8zjAMnHaEO9kj3joH7snNB/D9976uTix5uD7Kg3dTNy87+Hf
J+LQ8Pr5C32BdLi0jNvMFMzOwnJ1DNk2h5sqGzE3cyMxD0Vtuevumjjnpwz0QpN5
jLOniwpyWTwx5Z/geTKgt8uziJLM4xJkoI8UpT0BPjg5omh88ZKuxvt+2pUmimCD
vBPJZGX3Z19AmdiViAart8IpWMd4bV0VhAIjYLUXLmdvI1yPzpwpRS/Xoo8TE21g
YXAiWupbKOATwqTC7jc5rNO0fj91Xh9w+pZ9NE+WRxYPkJpGks+KJEYkiKkGfFPR
TJ3O5RYNYBzystYfZeJKtSjiFe+3ehVQwj/4g56aAduTdskl745BIvYhaOpYXCe3
p5pv3tQ+Kkc4sJk5/rlrYbZ4+LCqSarjnOgV5yPU8xGtup2ft6iz3tgThCtGEeA0
PGOxTj18gFs2mKY1TVojCXpfFDVnvE9kSYxaMuvQiEZgAQC3lpv1apAD11ANwQkO
eAg24q6UzLwFPlhT/U3ym4dvhQop2TQu+iRlaJ6Dy4Z9U1+ffMbUj+OxZAvv+oEi
ZQY5YQct3EjVumrO3WHB+tYPTTqaQ0zkF5Z46ktITB2P7MCG4HdWj78XiyCffm+m
K7jKbVlsMOTljo/K6Q2+Cd/F0ZkeL9oac5GV3vQ/rpzNJNzhIDGZuIMIBLyXIZvO
Pu0tSYLthn6yFLIo0wNSveff8TUUNKEbi2KRLBz95wJMhEJ/HbQYpbbiPPEjNgAx
B1brQ/KEHpxn6gBjWTO5Uvz2P/5D/uCe3p6cFrz7Lh5wFgJJdpLxOaxxOWLDgyxS
sYDE43LBH6WOqU4kKkusAKmIJTBlVAzhz6/FWZqKD0z43H5Nk0uimv9+bpeUxckp
ILjxtrLWQt2QvIg03gOOzTL/4UTuT6or7Lm3c0vjafbXIxP4uubijrdcXhKuxoMh
mhwOfSJtYi68v39ghXACMELnM5YRuiPFurJfDwuKc9WwczSbNDVVr3ILC1zgkJ++
/GAtO8arbLdyCbZ4kP4MmFX0B86ocSZmcycmR3jgGJUcVvNj88vt96hCTm83vgx7
T+piYZYVUwppaShqk4Y4FTogxMy5DnpArPmu4FdBqBCWeoaxcjXEPo5LNiZSxTm+
FTg121SLWjg9oL+UEErqcQ6FKgFxBPuhQ34kOsRB9MU8Lq+c5EfASr+/vvIdmWmH
7PddTYRZ05JqDN3H0dmvDG3eGQmxZ/oWu2XVe7+JRIhoBM6ARbfEOgEoBws83d/y
lobjc/eDeIXD7Qa3jum2njRtL+Glgc1i3pPUIJ5fF0ys4ylx+4GZk5wE8igdyUAx
Io+F2WPHwNN6M0WmrJCOURcCsmVVGoNn7AtC+7w5gYFZUB6i2drUbCiitAvY3zTd
hn/YjNjQo+krW/uQaSklkrOflPfNGORuaAITVZlqmY+8kQT/hs9NCRvYTTzunGx/
Iermt5Wobqjrf6c7DUUY/gZdaD48l/a8CLVURai2l16GrErcRu8z/YqDsXjyZhMZ
CRcM8CR+1//KNnX4SbevIfgVYimPsxDapfjV4jIXzzvMxAvk5hfjCUXr0Q9Karwm
v2Pv2V48UtV0VUpCPprFpl5OstwiXH5XtBLpMLpykP0oEtNYWbw/UW89/GGfu9qx
Jv8/Lk2V+kWLQOcE/QPGEueusUylw1B7FcH9O/xjOcsnKcoxfhgDsF/ZVmPvOQR9
VcX+CArr3Fzx+I++45EOAiyZHGfQAw9FrPxDbb2WAQ3/v4OKUF7QWH0Xic8X+ApK
79Sv2MkSHesNoUR6i7wPYofWP07remiIf6OkZPuZ3IkGIGzIXC8EFDJ4OMorDplE
vJwBY6AO7kaOAY1TK+K/kx1YoyFoKn4FZU++m9i+il7l7/YdH83PX/5C4sBnX2zL
oEAZcBqKgyyk7OWvNKM3S237IVS+3RHkmCdQLsunLLfGL+Cm4KUgHDKzCpGbCrOc
ae1ilJQoAZJOP6mL747uicKT28hmwCfLU3P4lDKdDq84kJUoz0lVa0ik6l1nQYug
ru9QrF8Hjf35IWRb6v80GPQO4NaUyxTUHrZ4ju80RU3wtbQbGDqEStEdney2UAby
/hrOI/7DN6WgA2uZ3pVEqG1tIcACvmF7zOwLvN4/FZWMFtbKXOylE0ij8AwkZ5RF
bJZvULb0FzsGrbrvZKgQ3zNt+kk93Cb1IooZfQ+VD0b0REoUYyCmkBEM5cliAoJL
BxWU0CXb9GuTyNp1mpCkVnzXGhVldv2XT6wp9UMOVPZfdq03l/9x8fRyIxZZmGj4
WqIpcupGW3JcWwPbxb52TAH6Cfl3pLsleX/26iNHljhxD10TAwYKuJ4VV6l/GMbL
E0aAThJfobaAt/5/s0UCAGh3fnItgDfNH0dPxamFTYC+aDMSqLOcN28OlpfrIm6q
0uXTAaKCP65OFjuHe+ENDdBPwaTxi9IkrMByvME3tR7TGtnV0ycMBZF+qMrahrT7
1hHOxRlcUH+f6IPmglvLJo5/7qwRcrm1/4cHTZsi//nIkqTUAUWDMMdWexBNpkyw
3lJyEGEbjPlrPhmOsJ1BMKZeZ43Gl7dKIfY6wR88W5ENThbwdteBGXpF1ERTEVPG
+sxx1cmi8fXKC1o1ZA7kssNY/1WoWdkOY6J4EV9h4hDV0CdVhGBGhBOoGPx/XD5z
sq6tDCd3W7j4M35XZWzCFCgHmEh+zJfVtnEj5Luuu/qLpa8fv/f7S43KC/Sfv7lj
FIW5yaz8kFoZQFd1EigQwbq9HrjsgfBf7G5vnc2gQgTIRGgq9vrTCWPBz8HHC7Jn
BJRAr+1YeY7nz42GJTmBuZixxvEa+HQMFxxolSh5AZuVnIzVgjZUmSL4c4CaMjEp
I+8f3fvwaGbjUlgotVNx3B+OVBl1rRQs8Wkd1iys00nSxu5DK3MWIHQ2WZZYtXNy
QoFsNIWe+hMaiLTNpMgyUIKZpVDuY6cRZ/ea5P0zc8NczMavn74Kt01v0oC3kZS7
eAu6IDb2Z95Pcr19yQdpESY7tGaUALDKzCh/Cuh6A6JjaKXdHbsD06qjtK8TrKZL
IFgzeHOoLWaH/+U8tn3gHt904OLciD9G/F2wiugcNWVb5AKoFinqZB2l6lsI+KA3
J6rseo/u2wu72eMKYsdmYsmMFXJJvabzzZVo65vnU7PGuMsUGkoF2W9Jv7af0eTM
8lL/7n/xyx5kICRoPReRJOPScAId2ShjFm4vOLqevtSquIPpnqEN47e0KOPZbX1S
DrDILnUONkURiYnToX7koZbvw2WefimIizaz635rTbqOlXz8hajSetvlKW1iCTgi
SiWHwED2EeOb4DLXW6lP5Hndht5m5GhYhP9eOLIsb1fWYsgoelB8944OfYpkxlc3
yvP/EdAkBX8t4oX2mRvUNBnIeEo0Km5yW60JLZEe2uWn2ls3boXsGpiz+i2VFbNS
bc6SfVdsKGo4rqOilqnJ5viK9hNhAXOOIyV2Hzy0Z3PfkfD5iP/zb4G9brLGy2Bs
LAG8xtA3u05MX8m7SQ+kcsSgbyRy+48JUoKiIUhZRho69v+Cqq/l0cA+y3m4iyQW
kNwl8+90fv+0shfV07wtu8gMtPmO9oNP2COBxjlh8ov0C7eMD0gcZkT/3NAyU/ng
QrbINmRnptNSEBAj9GPMLSeAnG14dyrakDjOGzRLV7IszFeb6H+B8eO71mHHldpQ
QSUXYziKWS80rF0cULiIGKbHr0rAL0P7nDjj71bmCAvN84TmWbRrRljmOYSioEXH
/E2Md8mEH/m23yXORTgJJcnpBBPfgJ31uoggtjcfq7nz80/PbM/HaJYgieIaamw6
BWjMD/cTXdkcoKWANIyDnvH4JuYP6r71BDBk8lLrVHh6+NOotH3HJ5j0sBdjaZvT
9+vaHogkqcv8cWD49bje+YlYmBguC3tebAVbJe6wfSEBSiaYPsrlGP0pVKrJac3S
0cQfZTuxNMQ5IZ5tz8dEUNJXb1aTcEWroPyz7VyojoQZsbCrDVllUtnQVyeLtxNo
tRKEwgOMwMlIbrjMWfP46wEVdAHjRqM9QZDeW0iAo5sXSn6dZ6jHQR705ZNrQrZI
Hjn0OaxpzBmjUAXZPkmKAadxKoQUnMLQOaYD9+r09aHrlBMrHxbrpLxG1H1WLCeV
t2L6j8xW/wekVFVdqSa4fnmEhfngPkOk3iqGzi8l77/PnrXayQNHrNvAaNs1O/WM
dRLFR8IhxBBviK80CjDmcRbdZqF5h5GRL7IiuMAI53IN8c+WHA46L4NBY8Kmc4sf
o/B/sPLekipd5hrgRyhGsp982xqLvK8tDDAU/eX9CXSlu8Zcp7wERoO3fZ8iXzoC
Ma4uVtu+aLLN8E6uL4frgHE8XpQ4DfXAy6luc4A4Nv9d0ZiOtG7JX83LqXcTDzuo
mIj0tIkT79yeqHlfktMGMn0c2xZtiIlC6oJp5mkYp1IVL57UW/Fwao8ygR5zC/MV
oKbidmQ3k/GArCTIARqqp9w1qU3H5YAwL1Ovly6z/JPBDuUxClBEgkqh4ndv4zml
AxkqnjLqX1FV+NgVAAEp359T3Qb7AapGn5VmC4MzoEQVnhzE5L9MQcd8qiLS5raj
ohSdDzLjF7E3BQGhorveC0eD2Q2cPsIjEMu/tRatrgRx0q5nm0dw0vdu9xbReqK8
bcw7HWMkz1Fw7MXRyy7PefdMlikjrCJ2eNCw65i70a0DQaCAGqn2mq4xEUlqzxdB
tUqUp3ltEdm3GnPMQbr9kHmABXrr6FkzwpwK8YyaT3MQqWc22Se4GPo5NkWKQStY
ApO8Vr3ZDFFMFt3x4w8S9kmhp1o8L3U76B/pLvjBbi4K+vvjIWJK3q6YvZ7/KaBb
fKPnThL/ZNGVfC6C2lC6LTbJ0l05a6NqA8KCgb8VT7IberdzHzu9q7aKDO7N13Xs
JcuMV8QQKCRWoJrjF7WDEsPHMy6OkReotMjMUfW/+A+/BG89rrJbGdDPolZ0gDxS
nuTPgKb8bWBoUgi72oj8v3aoE2/a5Y3OGvcAJVC6jmHeUBeFRfcfe02bqBpq2y5L
AXnept/Fw85RshtftDidb34nuCQNAW/nXT7H/YPATZE+g9wkVwqme3B3SMHbDj1c
H+jgNn6j0rl+S4DcU4vnhQqo5ptmEpZc7JNhMY3g8+ZnKtae4VxXjc7mwCb1m/P2
0ZOIsuVEDP3ghZaoKnioJdJYYngkC45kbL8mApl5C/Xs96rHJN36ehzpDAh9wu7j
NxNsZCa55K2oFxwiVw+ok/xr0y7lPUG3zqnQIwQdKKMcHNXirHidGqkEYklVNh9M
Awq1nOTFs4VAEUBjlppIKRSQGIXWh5ChxP/93x1+6Fj/l2LUAY+Gl1WW020ci2o8
qkmSF3LDP+s3/uyNn5U1mtdGMTuDBOtFLfIZFIrV1SeRRgtjQEJp9wQ1kHctKHXG
fB6XTLm6Y7nVIPh12HFOwc/1VkZI6d4Ghzqk73zXmVJoh9+3nnxaUATC/K4ghTgY
WEDYJ61vcEBBh/+0nJAhR5JJKx5rNq7ZZufAvilvUt+ehJNQ8XZk32p8SGuTYtam
2KAmD307tX7arch97j+QaoU0samcBgJQnGQ4XFWOS9aSWIug7pVBVJ+oytOVkffi
PtuIGIA5boCP8knVnvj82wwzphs5E6/3PT7ZNbAZ1sjOgwKA3uWn3IhxDNMX71HU
FrrXs50SM8Ys2YmcuqzjWVLVOXRWVuTZvzM9J28czgB67dLEIa1CDi7NzlWHu1tQ
exMY0FA4pcEDlVEaP1PnqfJHmmkMKedmdeDFTGgYfQin5c36vrBVy5iRC/IvZLSK
upr1hgHzBOcab5a4y8uSZzi5EgYt05knlkIbxoAZZ8udxDbx39O19bzlTLyWiB7W
UC5FJ2luUNPUL4IEHip1jzlYwPh5xkEpPMwIyb0lVIQi3AGj/CoDY2qvAxJApTQq
nCdNIbv0AWqudi2CjktbOVOr0JlIhv+pCWsT1wdM84kE7rKZqj+RVSwjyem+sI7x
5NBzZFwPFrS3SmWdRU2BCiY25ljCvhtSvzHJowitGLOfOBMNECxTJ5c1xi/cAX0K
QWWP8DJKT+dg4RYqm0ino6jRRwMu12z4L+124EGDKvzeZBfM4uf3BchxwmQWgk4e
mDHunhu3Qyqp5aGoIfDti1PCW8zT2pN/mUn7R81+J6cWmn0/Z/XG2XNtHsY82KyM
TcQBcZdmxnHDPKWaKcWpJ0AASPNs6Mzd9bim8yICVtaEYoryqZHgqvhhamNYrKsk
+eUOfGoKjuu2wcKaOTM/LzhtwT1TRGERzTC5vpjaP+9Bex0uDDvoCTVs/eqMenY/
goXXs57zlibljEmg/wsLHclne/Y2lWf62asG0W9uaXnIHPvy3ajhsCmJZ8Z1Pp/5
hEkElzz0S1MLlaVkBSKvRIZ1eYhxSfUlZbf/QHk5nuqTI+vO0Mba3o3lKYZAOY/O
iq45B6734CEy3iTrRZpIR3Agl0Ypzq4LFHh/0dl/Zrp2Kv+hbgQMKGEoj8Y2BLcY
Ipd5jfvhcPlUJ2jSZGsk857auegztEyEQlUAM/CAHlzElaiX9td3WpcDEcZEeSh3
wmd65kfF6EtnA/7onImPbcTTtjV/JV+zVerwuz7isgh1TnuCcZ3y00UtForFfPMb
aAFuX52FP16XMJWRv0wRCHSzDa5e6ov9yt+UbrFWSAQvHJcsYSCet0Cfm8w3PA6U
qSz5nlZW6EpSHOTWIFnrbhHgcs511CIxg2c776tWjQJuex2Fk3dsPjuqDB6vAF8s
nsEBEnj/2/kFNqadyuve9KAK1aDcWDWHGagJUjnkJ84GnDesDSCudY13nCpcCWJv
eh/XphEgqhftL5CjnaL2tms2TLZUaD/CdlL9ZrtnE2mf8puYMGr0x8lUlJLwh2sk
Kv8LjMJOemXXl3npdjzN4hrVBADlebA64n+0JvoCLvmMCw6WCkjMHLv85jHXlTJA
mwXPFLi3ujQ90a95O5a7DtWM+OVYuSWF9HevI8TNwsQLPzY5FC5Pp/x+6Zo8OQsw
TMRYeBMbUORJwCHE7BWjKvn+S76q4UczpLd/moBrFlHRJo1rga+SmbrwNehmzPwx
tHzx8vFbVtFWQu5CazMUi9d82ke1zBx4xZX7vbhWR5j9HDQJMJwpfD0aP7TDfC6M
2/bUUesliEiqdUVdmgQXAFf3g0HZmQlDtRky9wm02Sxgx28a9HlEI6l3kMKjLa6p
Ehc2E+XFcOmRk+G18w2kgbHeDQupnKThJg5PRLciYfafojGrjyLm3r/mj9Np1S9y
RNbvPxP6+FhPxCm1NG4X5s8sfZkUx6hNx752djAMXtYK81qBEhlFx+zzqqGRa/ll
LHiYePnTV+pCTf9oiQV3j6FSbfWfjwoEOlNKO/6WK624TEe/HuQ6eZO25OuSGBfg
+YW8+QJN6oVfvqSbgApLfi/1ib6KWwOiyx/REuiUYGWnuWKvo11HmJxzDz94mnu4
xsgl7U9QuA62mcT2LH81+/d7e6U19FrNd1xWpmRLneL8a/emMTgaF0KLUU0B3j98
YQiFVpX0PXRCrONig1xms8lr+HBCdX/izn1VTsZjK+6umtnxQ/LRDo/cY3x84ZyV
J2ERNEUlfRNbFfjjqvFA8L+TrIc8VM1wDmKmSf4ZxeZanF1mMeAeCo3r8K98oDMP
J4jXaKxonoKm6kjCKqJwJnK2iJumdpKDJLi4cuD9rCgeLR84XMFYx3lcG9gIXW20
MCBYAvn+Jsw1l4W5QOoUcRhRg4+XAHj6q+fhl9G3Z/rDXiZ14d+QAMkCDhrEHWuq
1Vg3F2kSY5u0/bdxCZZRDX4dzdfqFCL+eBXfrc4FkFbg115Sd7Y3yXJE8FwaCG3s
Vfk13WI2mkTrAKumU0kc8SBW/E5a/l3wWP0K3+lRfo9etcyxeg44Msb4vNp0aHxN
lNc7SsGxAnFGRfOnMuuwVJfbDE3WqVGCqhfOZqsNdm3orNszR0BefkGzHu7dKxRh
n3/lKLc2xrZ5vpuP7LHkZbMmLL1TkBmSgno7N/mHxM4XTdM6UoUbHnzgVDtOm7Dl
b6YFA6dLZwh2nhyM3yGL+pCcEQk5CyxT/wmvhYj9R8UHgKKojDL86LEzFehBbBCb
5rqe7HBZjtA/hyuoM1/cmH5+oVrp5W9wr26HqICC45clgxAhftqjwaMz+kIrPJBO
orpd/9WFvZ9E0yFQ6zHBy+k654v/8Th3H3vzpUWvPnk=
`protect END_PROTECTED
