`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VK75LwEKWYIFYHgZHJqMCmNraHq26jeu0f1/CS+hI1BkfuFapZiLvF/QnFsnTKBD
uASM/IEoMr0nuFHcDz472sWEDp1HUHmUySG/bXf2w1ylWZLQoSqlYRDtp4k6tIfd
cN8n3UfEWeYxUI8rPVHouCpuw9CUibVnyASkyDfjdhwU4EBVQJN4ah010Bmdq6Gh
OTkhVZTl2qzgDpnLY0+Wsn+ouO83NxAClf47rr3JqgcimoV5P0CxyjcoQfDRYaFS
gsZjMgaFr3UuYlxeiMTbquaPCwbmO6UU/Kn7ChR79UbXaKqkf/dAGV+88+X32q1m
MtebKmyKY5exYMwV0WlNKPBWoTJIC+a+B06NPu1ZhubimLmJ9x9qmdahGsZAKQaM
MV4pOdUqFGnJ7k0/GAheD1ITRpWaX9DGuDobIW8so3lVZHYjsoE46fO1s5WleZH9
OlPGJYKjwbMqh66iTBssDrXxmxGSxBJQWgtb8IqZEa3rVcKbdaKD4xR+TpsMsFZG
nvIasBGtqbgIYoXA80a85qOpPZ0WUWL0FVVBXNEd0LJ2cMS2ZGvItegZSFJJuTtY
mVsLzb0y9A0To/YBUD7gOzl7KVrLtHjoPSoz3yElQHyFUHwGlZ4KpLLTlNM3DhO3
T7gjojLf39Blkls6U2Nrf7s9jEcqEV7//QD2idzL4A+a1rnEtY8n4Fi4grTi3uIi
xxF7UeSs0VupDCqciBHb3jNZVSSDtYqwDk4SCSjBuo1OziE9TjG2gTBOKE8KhewG
qAHUadV4lOludruSol6V3vd5dXrEigdNcg9bkGTPlqX2BqJ2uk/pdeC7tDCIX512
Gd7w5hnEzYn3Uw0QoO30gUA/dPrUSMXtJTbBtfNiu77mIEJBju93nQTRmF2yBqVy
4Jyv+oRTstQ4dDGSEEFwRM3gyZBJeA49Yj7OJ/EL+DUUPIrtYNRRM4Di9IHrRhB0
JJkohEtxi1hSKh1G5GO+K+vtsk4wkXEXQG/+tbShxz5KH8rm9I6CwChWC09Kq5o7
yYv59C37sUVpaP2DQEmodpnXFyq6txBjAYWUASPJp2TnH3Gg8tv3VlCJDhHZVJHh
67+WsSDKUhonwg/BLkmC5oPy8a/stmt7PTbSF96pPaC2r2EnTteGi9Ji7FiXrkce
Du1/814AOOzytjVMNOptfbGn5Ci68i6uJGxIS/4OulJ0VrAjXJByd92dVXM+JM5B
n/frYmiTPPY/RseaCj50qgQnXqFrUxvI3gvFwYAIYb3fiE0sfF2ZgvcosWmfS5Lr
vb2dNfeI4RUb8tIm2cKdczqOvjU/mYGFSQlFwFWcttc0P2VNlUtmAh6YCc05Kf0R
ckA+lDk1NzfPmBhurTeAolYaO1Fg/cCuFf5N7C1Q8H2WKTa8vG9hao+M59skOsun
aLJxQUtig+9B+x685QAiaDUunipL9Lbem48wrst1y+QIBSrtzgjRIXS3oa2NCKf+
Zz6wvnCoOdaSSx8B93/cxm6yo5PERgN2IkYW+yIB5NUjEC3b5MtzvSRo3xCUerEC
3RrXUCYijBidBrnPgjUQkEKlomFs1e7KOgnIm7tn2NrPw2i3f9VFrPMlAncjXRRa
i783Wq1jStV2NjHqa9e7MRTO5695sXcUXjjQYU+y+m0zkWXlXcR110T+WuPXOSwv
D34VSR33/yzaYfPFaOlcUfxCNLciJF4GUE1a66vphlw8Y3XWGXYWrs+Iv8aj4lx8
DhL7p4x1rPbfLUDyWDN17zjGW0UBJuxqhp7zuPzDdO2IfdN+tHI23MEfDH+bqS/6
GfY1VKnPFrEO+kfQIH4jfVnyLfstFI2BGOtC7u/E090JgPNBmy5tuEnFEao8ZYN6
BmEbbpis8QT/3H3a26mTkcZD3y8v3U/h9bafE9jm7xvojxMRtcvdCtniCvtmhKsb
VrLCtiYsBfwOknopDjbCyHlkcl8b1X6VtXnLofdmJIK1DMAi4R+K0oxNfiZrqvQs
8c3XOyPylL5SI8TVWdntJcDsa573VByq3zeEBBRXdVCDPaIpvBFY/MGmUZ/2U6Du
viJJrULeSV4TnI4WWOSaiDAmGFqN0P/qeIFeMcphPJfNYlhvbvXZCu7UcjEkzyFr
LELPfA8RtRY2kWriQ+sQrFZzNQ8+uleaSq3tX/beh0FfAZSL79wiaBpMMKLjjvNL
gY/+Z0xnlddCnC3neHOaT3qzXkov1smrjoiCkwg6lECYQLnihUXfcZcgAv0v/+iy
KruJWMD8x6gIdmdzMNNcfj+Zo7VgAGP1s5fh+DDvOyYjT9GMHfTHVfRxpqXaPbAD
CMZF/Lwm6hx5qvUU0Xf49IGUZCny2Jukid3jxhv006ZdBILG9G0NNx9gAduledQW
HSbsspRj3JQ04zT0OenkU3Y1ZhCP++s+8NfBSF3QFmBtIEkYh0qblKi0HMs6ZKgn
0WTeXnJPNCgcpgS5yJyTMSEjXIMaYTbLq2cYB8pKGmDLeAWBEJrHz8pXY4KAivmV
x4sWVLyLWX9uc1vs5R9M9ybiW2ESavXibJsj9DgyAgDaF4HLP75fO2DXJJPBV7mk
AfXBAVKC9FhS2GFRXwFCdAvcCm4sgggoKjaeZr8QugPuebIsRMVan+/5EcpFr8+v
JBzPElvCIQleDSDOIMkjrQiVaiPKBBDsfF6/gBNnfkI=
`protect END_PROTECTED
