`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/X0/bSjLBfL9Kt+RaotDk2XDVBRk8+PpnO0Kz6+X2gYbn+MLZDkPbRP1ZPgqtJpG
A+YvRW4c4KJeeedgWnrPcwb8+VRaspre9lw9sl16GFHVOdAe1V1j0s5wW8YoWwF+
U4c1dqwlIEjZ5Vle6nFghpBlllT1oAP0q0ldZbPwxljFzbxIgEDPTQR5evCAvBn4
RoY+z7OMUu3oLDdlovZ3bzZb+fscuAo7Z23iZ5/mTaLcgDvSq1KU+d0wLW4gXgQz
7vwp8KXcjjnIPvGb50nlSPfWB/5jzWtgmNE0hVKhJqXHoJB9NJcyZ6eR/cS7qVOe
vE06MsSYBlb/L6ckGMOQWd+cH7ASIBJrfx11YrToLY5UTwNe1eT+J8wrcU0t1W+s
azBJ+FzFLXwXZof+/5o4ez7mMTe025EKrzCVqLAtb2DTZbad3lmMClRvKnZYj/Sa
BrEp8yBVGcEa+E/nYQPC8JMYlZJCIc5qbkhSrp70b+DPkF2LTrNS/8iJbFZdpj24
05+FCdfpkL6KWeldgMQjXztpZX5Am3bzUdLK4uPie71UoBnMuaAB3wQUdmFR5GOX
Bq6D8sns6H2N+tSS/BPH8E1detpmGAd/EHkuTSjplgGQlmXGdwkTClF9HHCL2vq/
knuUlUcsEZwOCALcoS/csZzmupdyZmX9qY4a7r7iXXeGFzrG92NX7nYzHjpIy5+K
YQl/ZCofX7m3ovt2If0af3rDysMHLZ64dsBwMWEAauRvaEjuXx4+75fikLMcxs3l
vnDvooOI5z1d4qZJqnUxlRtvRwP3p6ERiGcln34H89Lv7x4qU3P5YdXP2tqVN+JW
JgpYSdq3yGzhFkr6pAd3tyqLRbDTe8sE+FdRdtvPPyiu0vrl9zGOfAth+JMZWzZD
QEuRqCkQet2cS+y+re4b7msniFHsFXQFYT5jVolgEoeI635rMYhCM2dNDozNwVaV
KpZPrwittgaLIDOobIFA5/uGWt96ZCD65LLm1SU9Lfrc2kF42MMmV60SdvrZqqSI
sipLP17uJKvJBQ4L/VOJwr22nNY2BP8ahQ3VP2v9Nna+p2fB4W5ZgzC7AltfvKD1
igXk238AhLBc8sfk/0JF9kcdLnmLXSmiQm7fcafAY5YKQwY6HDj3yf4h4KVKhCPX
IqKPHp+vbaYo+WxFQB9UlDgkD7I/dELidodc/tT+u2K6Cr/iw/GLZz69VFtUqUkg
oj5tKBHy13+3Oo3mxRqEXlnEYMuda4i/1wlNvQii2HzSUQG5vWvK/l2Zcrk+zUAH
siXvn9llRhNFXpRmCHbgnSmGQBBkVc4Okd5zbAjY0E9BRutikVhHsXWERBNiuA0l
iiGLXXhWzFYFknkPMTmta3Myd1a6Ujhj0nTnnSA1OKEzZzap3sZPB/042ae048wx
0sGnBqP7vNMz2FywdeyguHEV9Cbh8fjKVhWJjY2xq75PZ+nii7cnh4Jj7Nv+D0zV
ptOYDwf3yqyQ+OWQV5PY7fUOIUsK4FECc/eQMklltHt0PGPXV/NVtyzKrbVEOEZh
eImPMA1hRwELterXTcIEZZgO68H3dnmppVKyUMjC/Istkfsu1l9AOfk9IeIPYCkh
XA1x+EyBuUfZw+J97wjAk9lQTZxCKx0+itpRJ/fXNqgYIhZwSLkCySkCQBWsQPO3
ysgQi8WF4S7uBIawkPEFCpGDk++tbDsFvQDKpU+AxBFSjqrhn/xK5/Z5qN38zxT4
p6lW4EwmgqTXdQvI/PsdJeAqPVBs447iiscXO12BPZc=
`protect END_PROTECTED
