`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q0Jl0bOcVj6vPH8bRAjLHXegqS4Mj/JbGPIQ4yqNL8obTcW00LbzBCLAHBOdXgiP
J8+kwZI2rR6n/U7Lkd4G8+I3An+2rySbIwk0yobEJOW5l4yWW0gvs7maelJQO8cg
l7ggIVtQbDH2bBK8bmZOzrf/H46VpdNzLeO8g4jWzD96YUxqXjqOqAknfnMRIV6i
piGx5AgJgBOD0p+Va/XUDAuUkt/lh+25LswlM+EVgWnB7UU2pgmzpHsABkZCy8Hr
JyceI/tEJe7PH2D8zkT/gQ==
`protect END_PROTECTED
