`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0baGhs0ERNNIM2JpP2XEMNm1Yzq/mMfXkhoXQj3HQ+Qw3oLPkDbiZNkHvJlhNE7G
QBfP3zb7faPst9WHgTwN9dE8uQ6QgzEW+9gHkVHsnJ6lX6ZfUIf9geP2rfNn6J6p
KM1KNKkzUvYtTtmgEyy5cauA6fqpJN/hW5JLHgocieA8uleVj1YM6+5ijLeekQYO
h0yrRi5kHSrRJb0qeWQ1PxHgRsuPsUiUhkO5oSz4byTtKTHnZjUqEHSRTd0GXwzK
vJ0pqXho0WN63nBILRRWcGFyq7LZI1RZ/NuTt7hanSRUt9UqP5zJNVj+tmgi9151
20wNAYYZHyXNG01dtQgysqbeOtM9FOQYh/0XefUpqnQt2r+w7ZBxBHWnAUxqHu5e
yvU+jlBiHsO/lJu159EfLSQXdvEnBkNXAPSSMY7CO+nkO6dObkU+QeJM0Jk1M0U9
Xy+CfcIL4aUag55scYRaun4IOm3DLVedEuv8ZtbrGbm5Cu7yDxaqby4ng96tM9vN
BwoLJjnxTqLgMKpXDYM3yQzeGs+sqPtBsOkMgqM5ynGnyI9TJpbjfccITKLucvPz
5mrrJT9F2Gcm+4WMP2Cper9dOpO5a8ZOjBmnIki+LC10WQP93kyuQUaVoBcfRacr
yj+iQtBqQoNDsjSHm4Q+pA==
`protect END_PROTECTED
