`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RCwpAznMu8H8awVfVTpoiI+lc8xkSlSRdeY4TyhOxSEybJoAGxvf69I1RLEoU45Y
wa/D/YxkD4UshHD4taKhk4pcFrXa7toHutCWdakCCDUni8pd1HbzUZ/EoRJe76Vt
y6La59u0ZjP+kOPpApt/gq/QEaAVnkti4hvq8Ap7iF2rYnYXHriWlDFDiKFasolV
ElIMgN1iycjkif7rhIZ+8y2LCBj98OW0ZqBz2YAbLxrq3uzCBp4377BA7KIY0izK
5WIPC+dA047YiwWhYFZTew==
`protect END_PROTECTED
