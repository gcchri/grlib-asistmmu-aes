`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wtkNbtwCP3UB54NoP8XX2QQzdD0lm42g8lPlaervPmW0bF+mrH7jKAdHAVFQX3ob
Qu78ojbQsawyqUkiTfnyA8ChLDB8512ItuzOIa5RmtypU1DVN0T5Pd2IDUZYk7Mx
BkXZpVDnyU/QVvFh4llaKKoPxYXffZFroiiRb5/fpyHvG/4+2hFDte2FmWZCxQ81
skY1z6dBcV547TI7nKI4WdeUaGedafaMPWVGHa8qzfRKyjCSNDqQz/uK6zi0dyH5
F7N+wQvbpIKzE67lPuqOIkdtFzgr8yB1zyN4nQUxRBsgFEjyaaeMKC7CTYCKCABp
UBuFTKJt0Ux6HNq8vogWdOXqN4nAUSnIsoFaYd0tlmrUdIcMRqVKsOSrdAe3cedx
hsZe8BL4K+vWAWcq1wdhkpTq0RhVcvT6Iz9ocuQMQ30zG919hGOnjLsVsLhF8v6A
zLobJN8FjKD/mqObqaoB0IsZdxIO5dvKJ+hkr0rShvSIC6ZL4qnOvUhQ+ukobXed
pHXB7RnJ8+JrSkyLFR2EHjMsF2n/iqPIQ8sZC5ge+vJXns8Ub3iFWIptm3Lx1ang
rzTn2VQ8PYgjnWDrAqqjjJs1FFeChqIrZwlAbjSoUVi+/llPJUFHRxGIlc9rsP+c
fA+XBl4oQ7xpXt/1Xh8XtZzZ3iDK6p20c9AO8Ro84mafbcACHhQdaUHHJAQvyp+o
xUhFL/mnIk2Ek6iNQ7LmVFi/tVOMLVfBuLeA1759R3S9e18NBSVjBiNK1BZCp1OO
K7v4Cf1FNqFM/skMbyL62wldLApNcbtvMZZW0n9DqnhHYrUGUtD4uccu41fftJdP
JuEqCW+Kg955rOSA1IE1fNOiyNhyN0l5h+NUmWl9STE9cc3s1yPAsyCEczfffXla
zCVkAelPlDbOEv5lZYp05TBcUuLqfmgMfq9MmtSD0pl6Nn7eA6t9ysYc/QvH3tLO
fV6UUxLPIU02HJaKcrSKjrHMiBzCKFkj6qvFGzsf46hYV20VEJkvwsDWVB86VIl2
hgn3tnG7BKteG6tC2GXv0760Fdgyfty06YlnIRINkxTdeWObYf1JvdJUHoJXsnaG
FmmxSUWVo8toOgWRO/UQVst5N9qnzA697RKm3PXioAQVJUkmQHl+GoONmL/846+B
xPUlJFHndH5tNjHg4NPplG50SmnektjN87juAMxUAbg4Zp42iClxjdxpjJ2xPzcM
/qMEtgoTWBYa1+vLCAqoguj+/StUrKQ6Q502VJQvDVOXcT/dEgLslGFceXJvOIQB
MBDKPgti3Cz9qFoSY/0aaN8dU9UxhRjrcFvNpuvE4OyjUlko1r55kONy6dbfu8NF
fi+V0Ve55x1ZLIonEDfwr0gVQ9LOlOfkR8vH5mu2YQFZtQ0tIQtpAOhKcam10vZg
mawpoP9scbkNxXWTZ0NcU6wafvDlkA68byvTOp5y2JCrRqyuEIlLowazewQEtkig
G6BcWNoTmI7oB5nDwVga6H5M7G4LwOlIAzCB88I8zIWosODRQJGHiLUhiIjYUtiK
n7T/fIxv1ZoBw1CKWtUpavmR4oY+Q9tlXygfdE9MGuDUFWjfAju9DKpp+gbhesbm
MAx6aMjQpVF1kmAIAKPxk0TYybAEq6nnf07cVKIM0Kla6gJiBRckR2/ULcacWwIE
PR7KbNmfsYqK0UIbr9JL8zwQK/mo+EiOC+of5pUjjh/4DjhyhuQePzOHaO8pF3m5
xKM6UxbQCJy+LfNlav0oXZ/pt9jrTYFDJ+Zm1FaybsroODvgletaMY/4pygegUxM
t7lwRrLjEtQz+k99RcNboIbshTrbbt3gCNzt6Y4/t3A=
`protect END_PROTECTED
