`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q/GSt2gMm1a9iHc3L/P3rCgGcoxeeTY546OnPPrY8cpIM4nTUKlZl2N5MnXDqxb2
j23bkC+p/yyE94GvEFcCa24BB/Ydzpi+rPqKsw4jtTeOTQLkefAftDi2RSw3z2zA
yrNjralA+2rpONE0K1T8yriT5QzWfCllJnB0TUnx7VBE8lB2P2hyJqQRC7Eg0xG5
DfdWKVaBHRZdIFxHRa4VlAcvsjzB5h9fi/POHoudC16EX6pBDJCiH7VYLFR5wGh7
trPSbCSEJscoRLpagm+9iZ9zsVOdM5BG+YZ4pMBwzCOuxwEVwl2F8hJaepk5h+gf
pNz1ju9eLLjdTiiG2dA5xXz1cvFbvJ1SLDgQwlNs8wTQky9N4eM5RTCcXdG67lZC
eN8giwNYeQEzd6oAiBxzgk2R4+dKYoHdwdGBNSrq2+22/japbyh7nxD4zRRUdlBr
TxqCfJNTuTCoMH2mWiMBOqq7xpZ351uBU/a+UZRS45s=
`protect END_PROTECTED
