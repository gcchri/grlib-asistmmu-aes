`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bOD8R012DPx0vwddJtPIwqAnOyoH5uTq6jtCBS6zIn+ShJR0RGq7UJOmc3gJnWkB
GQAjnTRKYTij8Zmmv6AOUioIOZFYyD+v/xvRY2RiBo0wB/5UQp9g/1duK6zRHAKW
gbdh0uXScS5uRH9m7RxfefhBzK8151u80xqzhq8hLfmAiEf6GpCu1AqvYoHo3TMD
zl3kLzAIQlJE9YyvCqspGC7zXGywVTQtwkq0XuMItsWS/b4xn5uZeARxgBz89vl6
QV50/MyuwqU9vrYKysO2zZw7+frVx6rgBCV3+e/onp7CIxRcN1I06gmoYCInMvAm
qn5iFeQ3R6X+uDa5Iw2diPzCYFQCvUBnkUukkqbpZrytgFri4duRGyWz0Pw0605A
MCdXztRv41Yw7ImQITg6ag==
`protect END_PROTECTED
