`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bu0X8OFgLggIUMWiJd7o2UEtJXbkrAX72W9ynRONC6MP5ETZaI9yAsIwgh3vd5bj
uaW0ZZjZcZ1C4AQs/vLzNIEAKuhtnkMFbUTCEpOBf+2wjjvKw+UpjaiuiDQMefiQ
qQihzFtVZzet4VbaeRmXUfzOvWPho20XxGG3vxmaWdA6URGTfeeDPYNbTbKRJKXr
mob9N06f180Cwk08bCCF9Qlhk2BddXdd4mQQXOzkV3hEKOL/H1WhbepSeIqT1/yr
hQCfcr0tqZes6OeJpGhd1HVdYvWFIKIJ+pLfUY0BQ+Cbz6yW9dYybkHrigLbbczV
MsPNrvIdNn7foXajlDQYmiPeSVWQt+tI3On6453fSfpwjTc3HQ9iADQLtyHF144Y
vx4STEe9MjZnyTS6y3gyOwk041zk9A0iCFUXt9fBq4JEvK6yCFiajo/m1JghwlFK
UE+20B5N7BrC9kb8F4DTBKHWd5Ctt5FZDeBxoDA4UeUGBt4+TDU/5YAOCWJAoVky
`protect END_PROTECTED
