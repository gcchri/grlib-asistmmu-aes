`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
760bO6YYdpYMip0yhatrMfoLEuhfPY5aGxNJtWqculQ7jmePEYhxzbqx7qpS2r/e
1d2tPfqTbgmN954ggkwaK+DQD4PsebnzYqxlth5K7ZSgPh8UB/OXQwtNG1SVYSXE
roAaZY5SKq0i0Y56U3caw1WN4R457HVAVttKSUhfXOla0ox1dTd2HBkQkxQYveLk
J6uqX9XwaY1AA8YszsI3eQaYIOOUbW6RcxWsB2bIDIpaEdrVV+LhtZ6WPH8mWmQP
Y/nwHDGSE3KOCVayD6xChZTsYwfTXqY5kRkilBXMvpR55+CbIdf2bW+XwbHUeeUV
rv9cLyBGy10QlWENNmT4ONyCmwf9VpOaUMOVHd8ulXTQoUv3/cX4yo0ARfqokIPo
KEkheykkvXEpLzcAoiTM5L7F1LQGiIloLurXcqaGJ+psm1M8sKCyvnAnZVa648M2
puQBzeq8VFcORAWEbOfSxxRBjCfd+AJ6Pp/MdALK3cEAeXJXSBTD39I3CSx38Lmg
1BRWTJAbRFuivWRoWMZt79e7iPMCXrkhMYbtbK6DCs4c+sQARrGWro8JfwO1fmm5
`protect END_PROTECTED
