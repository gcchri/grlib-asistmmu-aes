`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RloVbbxmkwXwWUD/nnOGG8/wz2iv+YzsjFV0DybJ1Gfx+VP81W5+YPm8KI3c3YS9
W0x7QKuKy0T2/VV+VZ8P1oIVCWLaNwMmLKnGAL/JXtl4uii6L2SzZmu5H9mJ3jqs
2ozOqp23yH957bV9yo4ins3nGvZgJr0KhjTpL5PJ8R5II2pJQ+8hkCwKC5S/HMFB
GBegkAqqkhFffVvjEwb4TAGBa9tnS7A6fjNBeTPy6NXYblUI0RYP//R0hoPnls3l
nFgUKEZSpyZaiUDcJL8Qiwzixc2GmlxtgZ4LHgiQ/m1Ua+hB4b9A18HtmyuCEudw
2tNDdjSGPscq22xDtLB2mQ==
`protect END_PROTECTED
