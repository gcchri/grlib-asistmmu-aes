`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y3aXTN7/5taUwnGgSxPr8SiaZ+v3xdRknc5bZJ83WMk4wq2cuETRH3L2lRPktcsB
0kktTXTUcCd9hBwmDADMil948EqXT5Hbg/ogExsghEu2ulU1BjgTWB6orJXnEquk
vRB5fxn1I/YGSewLihZP6sDm1LaLDgW4xfyC9jTengXOzD/8047+xSLKJXtRtjoc
dKPgk91C28vDXNOhQjMLbDJkY8TLDX4nG56DJzy+bCc1qvDyWqB6HBqxW8sdLWy0
F3DIgMSaGdwIssYyEhboO5mn1e2TTeFYK6UZGN7Q2YVMFRqj6+1wSr7vVVtde9lj
9KeH3FsQGmyh1WZrmG3MSRVGq8Z/KcYjIumZr3R4zcTU8pncEC2oHIfJybJWROXV
pJJ1kyi0dWjnL5cG2Cj3XQ4HkA4EVE2Nzrxc1e08hg+DTiZQC3UXI/TYaPRo40+z
EwLOoB7n/pQ+SGfYCUZoglZEPUeQeP4IzxIWKwurtKIIPiQBZEuwKnwPBD9V2TwY
`protect END_PROTECTED
