`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bohSr3xgewDp/AyGsr0lXJSByxFr7Qzjx84b2Wzwf81eSnhyyoS1grHiXLa8OoJH
hlvQ7Xtm3JI18hw5w83rhl+Xjn8HUJ3yB596Af9iKS9UapFnYaCnk+ritihYia5R
8DqOcn/CcRQVYc0SHw+SU0/XhdmbGx+AFgLUWBrhz3+N6NDwN1EPLvqokswfxyCe
v7/yhrcTJ+nS+mlpul7kdzefSBJqi0mQXXT7CeeMu91JtzP19ZwSpyYZx1PQAhVN
fGE6LGkxW/4TgULdsBu3PLv2bPXeXzvCdfCwUbgU6AmMTZO/g4TD8ANtnuG7LgGK
VQPR7VM7HN8dpD9G8SUHRRzLk6sJo6eirm33nKeCOrJMfAAHikCqozg1AijZQovQ
AE2YR34517FlYhvxjxNkrtQa+Y5FgFEEihskJOy8FZPPd4AsxNclDAyueRGSTOaD
BxJqz7s7YImMoJusGMUtfgHXoEKdJVQgRSkseINgXO2DF13V+sRmJXeBriHhHK3a
gQSGoUcOnBmqOAUpSswacVwCihdWq/09EE0LDmu4yCFJiERBQw4xR+5YwiLL5Yy3
bXnI7uFJpZc4JrsDMuf0IzwGbGkTnfOVbVFmTu+B4CQ2ipivyT1/yWusdgVvtgrX
dNacRjxVBORg8WQ/jMmtvj5AC3GN3AqT6LDB21nuSTzPoh6Cw6XR3MKc8wK7Of2s
qglCTrD0Sv8Qwus0Whmi9VJecyRUpYG6sWYa8Ur4mw+WLsiurqUWjJ0a+q6zRxuG
EUIu3DMNBMp3nbSnMaaV+kBAsf65KXMH0NUDgMsREvpgAHhxPi7HdtwCri0FOlrx
OjbA+IVPwahBgDUXsXr72th0zG3aXI1TZOVUvS2H31FTwowykIXyYo4YzAo+AoJb
Hgjuh+nKuS5gUiYNsGWffcW1SDPxk7ljpB5ocD8nXv3/DLk0rYJZBK/wV4N4al1D
R7FkU6/gyu1KCZrFtgi9UF+diIZy0qElGjt6xPWNBe8Xgrp43QUqqkDMC7TggyZr
QRZJMjQrkDaZTseYs5lZcSvBwwKMDCYNK5AXBHwKLGIOoQfWO6Gs1L6HoWqcoqaz
dj32nX8Cwo0RK4civJrO53tw0nhSp0zcLOmavL1hxPUJd6fOy40iArLFrw7QHpz6
g7ajqFfHCdNNYVrs9sA3u8yrYxz+50Ia2aNQ8/pMFC23AhJGvIo7KZl3ejNPMnoP
+Dy14qWRnvdhn5wyp0zFSM8tsiw14ijWpBz8cpYkdF447wfgcy0FOOT21twOedgZ
/iHauItPEFrpFP/6Xor0DVo/oxjgXhRv4ce0ExPVYGzDjRO+z5LO9XkaWNO4bvML
mDhZf6DTcFp2Wz0dtDgmabBroWUyTnM4ndyM7yMQFTx5HDA3zHqKVsknF3UruT7d
lnSyy+TdH3Uz137va5dRcesqVUP0G51GclgJ8JGKFhBmqJ2eyXq7XbRyM072oCBC
/+jQE8K1GqLBodcCIPcPlCffFMrQfl8jioi3j5p54ZIV9WP5Ei9tQ/56Kex6a8AK
RD0XCfyn/+eu31xMJ4hzjG5CV9o1K5fVY1Q6zS/hXkTR9JVoB9yVUoPspztBEHwF
UY6+d+F8tg04UTDrrWGYcjRqPXSheYfmwekfRq2EJaQ5U6pc1okGZ0dkm8uFJaqP
bLk52O8NFzCrLr24QVU0zw==
`protect END_PROTECTED
