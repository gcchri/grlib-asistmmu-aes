`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NHyGOsCRho4Z481HDZWvVZHkhNyi+FJNXTk/7rH+dKP0rUQqMi4JrNH2TzQtQStJ
Wl/4phlyzFFf5g3h39oc2v62rmWl0kcw+cQvqmLIcGEpvd0TP7V3pDnezAvY7/MO
YOyG/drXmYV0FfoUXn5JWVqJ9Le1sK6YFDVP1Iyv4ORzcjgsurs72m7o5Mw9ll3X
8+pCson/H0T/us04CZw6uq3nXbeOC6jP3mECrjd61dBuge82mHEpGaxTFCEZ1epi
tFczaIF2kLpjsCscRo4kWtt6YZPyB1FKRvJJ8BJ6b8NjXlnWtz1Y87pCeD/Y90u4
23++x5jNX4xjaNXlP9Quyv4it/Skq38DfD264WpuuSgBFphybXhbP6064MpaA8lM
I/8EzP5ql3arbZKfYvHmwlo1T2fmgD+wQLu6oZTK2kyGc+Pep2v7dDDv/UIYVLAl
HYa99FY5n1rYdqLG6pAP7mFh6NldQDbr2riUVfeiTg3GsUmtxBEDrBEk2HV8U6tn
O0NnMpYXfsgkAT0/dDyj5gEOrtqRm52mmkjB1L1yRd0=
`protect END_PROTECTED
