`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SDiJ2UtRXoruhCVO3vXQrRvLclUQtZoe+dD1qgZX0/rtWzHXhmdEv7sxRW7fKai/
CqSYnA5dOF2A+Tr015hTT91OnYL+KE179kX0lkD9T4LkY5H4Mv/++vFADKDVtIn3
7Eshs+zsE938R0ZaiamMEz1S4VMuYMGe7cdlgnn3b+mZNejxnB7fliptS9s+raC0
2o2QimR+oYsw1K/EwqaquFpvXsfRKHzMhh/wkBDdFbyXh4LIo8xEhhftrecVczoE
JyYXpb7pGXSd50I39VyNyaB2RTNJDeftgxzuUYJO/fVYXYXa9g8IqmpQAiyNkgJL
ySmr/hRoUqdFRn3Clco6Pv5YYQ7NxzAfu9drGvRwPY72ZNXBufiCASDDuXuEKVzy
p9Ls+y65d284xB1O2+cj5YytD/enGcuTBw1LmDXqGX5CT8WzUIp27x2Gqsh/yk+b
ZuK5bWkeLU1cyhH1e3jF3y7zJjSE4mK15R+GspKYPtXRZRxCKjKt5zFvKL2LBZ1U
9+XPNmES0e3VdsSZllh1IF4yn7kxJR4LhsmDfVmGTxz1/jbRxfA6CmpLtPXKfxk0
2c6xIryCxQyTjQU/d5iiqFoN/f9DBhJOGOmFtrBbUe+yuPAWKQY2gsFrDbAKm/cE
xF03URIr7vEw5+9sRikYGCM9CxF8i4wCSVT5o6CCqvH03LCNcWMJfh+jaURTHOhi
QJaS5onHZ/J18sIZdhG/B0eGLY969LAEDDyfyUHwmfwaU9R1CWj/U35FaJEJFnef
EJXpfbxdG5+LJDHAvBgiEhyBrbOV9f4fKXrNKeooAZqDJygw849RbHGmpkvwHvmX
FCfbrt5Uj4oQ/tEnt96wN7s9r3YSUTNn2nJ/7M8rWpz+NCeaGani7iiOSgclpmNG
F3ZQLmY8gYrHlLoRmAbgEzp2SKm/acmaAAAL5v5+THTeXCgF8h4GxQ2jTb1cl9dw
coGt6PYcWTBBYuN5lOdwPYa/wDcUssM9MAwxMDppkJ0Q0kVLA8eZMH4jR1r+3ZEC
e2ar4bJ2M7DawV1RigWGRoqimfcFIRQfWVfzjEVaHv7jbRu9t8e44uZ61AF0ebDn
um5w9JcmEA4FZA/vSwzuYFAqd7BxAopLWVxa3DwMzouvoDgIbgR19EM4W+fjsn74
5PNEeaIJjupn6qL+zRhrop0qoEhQ2yrt98x1cFkAf+DGlT2iZqQQy7/KoXVbI7RX
jq6hJmZUaUdq31kMuca65DUXpBzn7uc2KL4eFlFfXOsBfUOw1zhowpxi1Aszt2NO
vSXTJFbaneAk6F4S1gFtxQVSQlrGeUIoS+KJGcPVGKhbneJuHQIv6qJvvw7smNTX
04IiFhJ/CQf1rI0P1tcGtNRP4iR+81geTeJBpSu0hbrYqWkRh5YWHZIyQEwV8Vpz
/Fq9SMgydhxVVz8fU1W1cOrS1wmCScZdwW2pPR2L9ocy5bT11WC5iQMam2QnJlNs
MjMl3n4u8jx2HroRLb9JqnrFBk+v8JpCHUsCcLNHzSrnkPwKSxhrNVBV6Eoqfvbd
oTA+F7QU/oe0chtwCF+KCjQmnwva0u2MkSMB0akHYw2yKqzUAfPhCgbNsBtH0uTV
0MhHcTqimFVSTYBxcnBDSZAjsdxpHc+yPasBOsTejIzDcBKCch9Sb2vxELVB59Jq
OOqw6xScleEkF867mysHyu4IaVe/TisSpgB8qbdiYLAwHkfewAvmmlMwBArEhdVQ
7CpK/Xq0R3UDbTCqvmYyeqhmMhiV44Sy/wAq81WWJzB+9NyOujinvoO3LUqlbniF
yUdRVSgthr8wOlzaFFaliLzd/nh4T2pXJwvQO3EvpQkw/QlaY5oL9suXXeC6dwMM
qlDFmtrRLy8WOGWQN6DEaqXu9t+43xQpLiPY4NSDybx7LjxTg78cde0NcWcsRTua
9M+uh1ZE0oZwHkhzb6cnNWWMWcCTvkIOCGCdBmM7KVrKOPN29ugLaw0TYStbwXuW
WxGmav3TNu2gYO2XTg26KWhMs3JYZCJxpj8DqsEIgNGHN0fGyCWhxTg3f66lx0Du
QDncaDZVi8mUKoK8jd3vIDTyfPFinMQbOQs5TaQ3+3OLHk8Wcu6s1Vli+AUnwELt
ayCjwVLvrpbcDHZoPrIJmwJCOJSC+PxoCqfI5aPRrRryqZ+akNPW+qdwu9iM+ge1
Dxs16IMm7mb7dCD2dsBx1lymIlr00DWjF7SMRRqQ3J9Sa08d19QWOqDI4g4zv0Tb
AJBaA1rFogV7/8cuo6vsxjGjlOJkNG6rOnxBMcT+wa6TSvTF9xQCYzvs2LiDfBAc
RXfAqPSDh8HirzmqSxCCSzI6+HUP7Q8GpcICTmistIVTKDw/x3fKhAPyIRGjnpjV
n7Ljuwnu39vnx6j9DSD/MkKrGWc8p92sq6LDO6P/ZiNlkKWlg8UsQLKy7X0+Ca1p
oXtGvUIz80tVLJAiQ0v4nIBL8DzUhTZ9UrNjG1NvsCuCv3lJnFg12KDAvnX3pVwL
W+iy1VLQY+t3rNwHXizhEfKxTsGAiMtcueZOMtu2sjmJg2oVppl2c4/gPscuIbrD
iK2XJ75V7G/9aCdoh04y5g==
`protect END_PROTECTED
