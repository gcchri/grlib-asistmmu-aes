`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M4hlvdl9TC/rFRYVF/PsxkFn8UNZ68B9AkkepB9p6hTcGgG9f/oLzUU68icPcxuD
aFHqW+bUaF2EtEXXJq1UmWzfroR4C+t+74U754QCsjhocDg9fNzcICnFsn89e2yq
5JAXr/1+kbuzkGT0vqb1jVt34Oir90bnvF28LiVsOe6Orcso0Fp19UWWAgkchJJR
NuyQgvShYkckdwYmqKEvTbCdPe6FaRF/PBIU0ALuO9z8ulP8XF4JP6mzUNe4u4h/
43jBYQ8CqsxVvnim2CpD6pGjdtr5fYdNuFTisANqSdcKV2S7y/frg6vsH3b0pumC
Wfm5Tet2NTCL/9049G8O7XZ8NRKMJx6tQLoeIYgYohkt1v0hcNKiTq6F2FnfSPVu
b6zdeGXXpl0zjTHOkx0nEGmPpyC32nkdzk2WPseegewjaaMxXMwAZN0IOosmGIUh
S5Npiy5OhtDjyTnW/FGfwbkkg0DFRZOGUvGTHSIH46Q/NcquoaQI88EZxoofuR3k
RhnJMOBNvwYKzgR/TMnpWA==
`protect END_PROTECTED
