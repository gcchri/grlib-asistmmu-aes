`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UMxYHo+9F2VlN7kZ2g+sFjYnfCUSmNVYfDi4YTgGktUomrC2lAQzj7E1CXIKVD7y
P9xjsX45zr7VybsafGE5/Ra9rCEDCe5q8GeoXXqLbsF4GVtffR8KR4lu6HwRvls4
Pq6rRdbXRUhslJoCTkKGqZGebIw5hkagq+L7rXDk4YeKr8Tp/wzH7GlgXZLeObE9
QY8YhTbAdljvwU4P80cTm7zI4iS0MD5PUsDS9wG1ByuRwq9Ta27MKb48flsCG3Mo
Vdt4Oj4zHSRvwnuqHAD3DM1ah+LoCtc3bwkJfCSLqtCHEaSyEwyEOjPGRvtSubBV
fcHI8VENZJ7e7PPhCKcYW4+yCNNybRKd3wOXSFAyOGCAORN7JDJZCNxeipRiA5jl
4dsfP2BgRIvTBc6MJVCoie0MSaSXc7wG8bx7cQN2QgPx1ndyyZUSm4y3Pel7rIIN
3acI7gVwuJqdQhw74L919bp5sVlcIv5bwLCtXELMcvGdUoYoCku66WvN31x0clu9
z7u8+2ELE5kRp336e3l6TaQRL3DyPt457VzhTPRXFeIzTBjfFfVIwaM3cFG5LZ5+
cJcXx5fY8+PqpJMpIOR1h1t/SpbZZdyxCUVB5vQMP8H3sjQG1d89joQE0nRK/D6Z
TkD6c8r0aRl7Le2Y8oXub3DxHdUhedlT6z1gy3rv6RLc6GytAMpBn7tOQnik+j+G
zr7cpwmpPfaNOL/0x5kZxaHUM/LbsmcbTdVBgVvmuUK6qIw8K0Pi3fJano5gRWAC
9VjIik+vatC74SrOCWvjm+0ead/sit8JdlFwYXVbK/GwM4watKS2q3XR9bNPkvZF
RLNhrhH/zCTcOPAJOsMO01reIpFvjc+s6WgLDEf0Jvy39uus1lkwRHnU1LiwTCm5
IchAMwefOtYutgEwQZH3OouvN0UHm7FEHuyOYeca9pf7+K4A5wg9Tt3sAYuKuSA0
s1XKUo4tUVkX2xrxhKJaFW4O5qH5BvswERj7PAK9EtM+1TXt7r0BhcqyMe6HchFN
abviHg04T80RuqdhYkc2rQ==
`protect END_PROTECTED
