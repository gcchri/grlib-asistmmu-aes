`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rMjxnuLbvEsqzWKZeTf5am2XQYIPjN0EnxA95CWZ657zynf4PCh0nNYmcdnxjKVq
r42Y1wHSvbOYqTHQkGuA7uXwA5eOyPqx93LrzIF8xUbCNx7W8S0eDM69JfTrBDuN
KyOwhLAIvyNotwR1wnQGt6r6yBveReIdPs1h7pvD/n9u7i4vlO2Cmw2ZXmcFh+L7
CnyvosuDrYu5DLa+kliYc1Ep71gLfsHq3OjirywFjaLW7tOMzvUYnVjQV8yfhxz6
mMN8+w65pO9CBqv0mQ4cs6q4d1QUyJbEfwcQlMb9o8fNn9AMQvzed1wX2oHmQTxY
yd4q8YKNsDwj8NbzGcSp5r8a/T4sfB8oCK8HFPZMZ+016SlwChYaSAQodxq+X+aJ
Cr7DXFssbxn6+JzEyj6NPkOSpMMVQZTNnOPnjtNuwFfP/91E5UawfVDZgCacUSgb
PSEQuIet31ix3pDU0zrD4uSHqvicfGUry6jdyDsvZt3Q5pfiNbwBLw07YIuPBYDD
fnuSzpN06J+s4A1CM0oGkO81kAoCwPMVopq8fvW7cKSnfwB8bMIOAYrCNXmWNYzL
yW19XSspwGPLmucmelJqtzyHIXNUSCVJq7+y+4oYQzpbtot5SYQ10F177dn7Vofi
XgeAFN5PmhmCFM09z0+69kB3N9RKqspJBzbNCRYIuKq94qfKbwVjPyX/FeNXax+7
rcjusRqQpl18iqn2TP522sGbI42o5Tp4XcniEhMIEbsCTxybCdm5ykJntwTyA5qO
`protect END_PROTECTED
