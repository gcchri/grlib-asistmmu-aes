`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wHmjP0CbtRl83gpX0NXfG702sa+lbPQBpNilHmCCb9Zruv744WiOi6I9ikV/bb1d
8gPHIONVMqe9Sxg75i3oKyzHLB1S95k/d0W0gGR9ofPp8hAZ9P2k9Z4ifpy5OSiA
cRM1+gR2fHDBK9TZYTO/Ydbnw1eFedoVo7rft5h7urbEPjppcT6Yj9ooZQq6lXOo
ZJEKatrDHhmn+bm2n/vwPI8IGP61JAEwNkQ+tba8znrGKs3r2GGOUh0AGMTwlpG9
PB3ltYf0El9P4aFNWhYS7ie13hjaPP1FsylmIwjPpYjYRc/iqkhCHU+4d/uOh9M/
TBIHugQ58Y8Xf+XQ3JjENjwv5/R1kg2/Td2cVf0x/Qvz9zD0yTQ5w6b8QKmx+OWH
JCsAdAarV0o10HprzHfmyS9UazJIhyM2xNZEk/zlY1vR2AekC+fp9mfqFe4aesux
eFgkrfg6tfxVx0yCWV1FWTYrq21A9CyJdsoxV7dN7K+PV5hgNaq0tVAqCysI6AqM
`protect END_PROTECTED
