`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6pBgPTIuHRvF0Gx5BGPk3aIJNkAx6zOZDzWVk56PNyAEYRmwSopZdCoRzKPA8dEU
aCpb5j/7zkwf3Uf9TrwuqAH9kSXDCpOKliDS12eWZcQPL3JO4EAIb/CMu25VykxW
uR735M2xY/WGNmwq/kGn3CNj4T4YE5jVVuNoW0LkP4j1UYybadgmt6F0LcJzLMMC
dcjBckmchOasc4ArKN9Uk4jrJvppPyGBMcjVVgopXxU0Nh4H1ZbsdUlpk/Dw/AmJ
HLOp8bqD9BqOWes63bKj+5CYGHUSl2x8xf0cIj8RR6C+6jIr0O4jLGUvtqPv+30V
kqfzeKcTQqQmS9BsettZt3zh6ufML8uGyyc8lLrTbGJsN53pYYi7MIN2pHvFqgps
xqExOuPqmtmYZhOcxMVIPrwm+Q5nXZfuKCx3sBXAdT/mQzwKaBmdA86KwNdh9WC+
e1LfWmPyJJKhEXRJwWKLWBZLuCyhu2uEBjn195U9LSY=
`protect END_PROTECTED
