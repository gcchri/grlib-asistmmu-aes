`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UfsvRxbTmOL/YJZumo0SBCElRPqT/hEV0fMB8xGMJaB39rzbQDl+Tg+u7jl+BG+j
BTG+NX16kF5aRdiREcg2u9EtBcPRhx9aQoievIZGsSci2IdKGrHxfxhXeUdYYtWu
VCJmM2QnafrroL+k69o2XSOT7S9VMcDpa05gSvIy/R5yW6NErtifHeSwAMveskZW
57tvrCr/+LKLFJj3q8ShZY4qn2KT80Rrp/kZLXK2AGlZp8qOtC6co4RY7XCY/UHD
VAkqjD7F4T4YtwRE9x6KH+1jjyYFhW2pUVK48II3tCPpJcr4C6BQr12tvaFXU5Lk
`protect END_PROTECTED
