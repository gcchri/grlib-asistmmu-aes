`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gyn7h+dRm5KrZTJBxS/GtMVLBxQT41DcOKFepRRpsVZW/h9HCC9x8YAoGoFB9Hb+
BtR7chnPRNPjC2o5nS16x1PVRkpLV9aTevsBgrDvjkEPY74intXkGcsI2HgpxHiY
TQKJ4z8mVnMvb/n6UMFxzzJ+76G/+Dihyh2Tk3f45zuRJaz4lt5Bm6mDFmpfaT3S
VqDj8Id7u47fnsXQVe4oh7r3Bq2OdfvOsDsaHXHeao6mimtc2+FInHv0JUoDEFI6
jCZLjqv78Gb1VeqqezoNs5O3ENGdN8tcchu1MHXp7vJSXJ5kebjngZn2qcHS2Hih
EJg9wAK65GGl+a6mNlGkoC3x6TyseyrkFLfChdMvHkbeY58oDL6myu4H+zgVBePb
UtOStj5zOWkLnWvcigq+YsNKcOCIpoyX3bKIrPdpoz6Jt9bkKO8vSU5wdJTaJhe0
JAwR+knN9gKB+uXZPmycAwNRtLVmdZuUQiGE4C+Y3Xpd3nfKc0KX5tNauR6cY6OV
Klx8XzNwJt12b7sVURx2xb6/f7qsaOjgEIFbE9+anUxJXDyPoUbLRQ91Nz0lCMG6
uOYoRJGkd+LoIkHrr8C6NuM+fiWCSggkmHe40J4uNgqD3fJ15SH2s61VuimyU9p2
CCQ+nx7yQM8NgpYB76+MlQ==
`protect END_PROTECTED
