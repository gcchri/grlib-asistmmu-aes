`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wFKJ6jfGt7k7rj02NJ9kimY9QNY82vcjk6QWmFKGWZSp3a1C6o/PSTG/LF7c9rza
iopNKI4FkpSoz8/xRj9rsQRi5nyD4fi3AUdgiNp2CnT6gtgwCExUE4aOaZmxELKx
Z4lgiFZlDLDB9/NRMqTBemDNLykke6uGiuOcnK8LWGsxS0Z8+teIxS7zj7slHkXk
Ba7WCfojiwkMHxMarzk97vX3rePWxURk/AAa0a9RKP0=
`protect END_PROTECTED
