`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o8SCjTn4Xj8i7PybIeIMX3VJvISrzF0OApeAScTiS+6ezFpBI81f3Vun9ve7tKCV
S3PTRYD5iMioQQl0xKgvBlhHe2NXaFwGtwwhJJRy5wJwn25EOuqVjQzlwG2VwHC5
aTD5mqLSJlr4Bhtm/buwNPBZcLIdw/Ymm0QmHKccIjfnHApPozCUIIn0C/LfvkNT
QQzW3zFguuLebEVfSRfGHXuG3+rUb4gB0/8JuEL0AYawUALddQ2l82G0LmZzDBup
VGKNBTY3BEBsE/JAIsR1345yCJxurziSPJRahE/pmfjpuOw37NwA7fU98Wq6jQZc
cQtSFXuIQCF0rbKvW+dWHSLiHyGuqIkT4frtA77ApRTgBQ437S5TSX4JolzzEv9D
cU3QLwhx+OSFYDh2dhTY0DpnON98lBb33Ql5dWFtasM=
`protect END_PROTECTED
