`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w0wR5KlqSW3Njn38Y07yJyDWzTfemfadN/xReFxay5tRx3jW9JO08MmgcDf7crqO
ZmWXg8kUGrfwTAgKL29G1W3UxiiLFbGMh5xeXyMqJkpyHq8XgDYsjypBEY6ML3KY
WxGZpG1ykFKUFmV1+mbxQrKA1+FMsaPRXkvySQJZ5DVaOmE224W0/NL+LzmO1p4m
UkSTfiTNN0m9a+LrO7ydbrftidDALEY8xUcE7Egz9nPH8h9E06YZPkv/x5/vD7Rr
Ndx0UCzwShQZK4qFyKCph07tB+cZkDTpuQgVZMgRVaJdCuS3bczZMw2yId0hRISH
LW/BZeHR9/SpmrYs5nDm9B2gHNUbdIoNG1C8Nl5w10pFsnMshdTS7g24e853+CzH
vXH2AabYYNHgK9UgmEF/pDdrmLblx4z0ZXhiRHi9GmcoII+AW1BtrvlzVnHlCylc
jVnfnz/JIUB4mppT+q4BPh/bgl+l2hKQ+r7wBwluZknaKhnzcjGp2yh4uphX3UoA
GEtNPSxQrIGLIOwwJZFx23Ch9NFYs5GaSPbbtAEfpwRnvBLFhNZvdAaq582obqqU
RAYZGKJxN+BU4Cwv357IzlQSxDppKIHgmCBCgZ/2bIzmK4iSyj9bOpjVSOM4g+Vh
8q7+WOisx2AnMRdLjV1nZoQcY0CcmC9tldx9nKApa0hnXE8CQTtQ6w7r9q0UMS3w
4J789kSJ0+A//N4qnFPVhXuFXHytefGDtrx1m6/q0BBN33JxmWRNcL/vwrsaAl5U
9sgX2vBzM5WNRRiFUvz+yZm+dkgl28O2tsvDa0NOTSVtaGnudDv4iovVV0RGzErG
5Ftqj36G/Fkv3yqfdc8fgX82uAoI+HeJekvZWbzp47348ZEqLeChj7GK67MpCpjT
QJZUsY/AYYGHuX5S91qcU28JshfpHUddnc457t4DBrk9l6gqilgeV5RFBo/mxqxz
uOqNZVO0C9SHpAf/yNCWo5ftU6BYTuiirhvqycSp+Dd/GlYXeiwaGzQR1XRdzZLu
4W35G7cyAuizUlwblcX0yNKV463fTG3edCCTAskWNOlCw9YPbv6UvbJ2O5TfEiTZ
zV5bzASHoiWbCCgUVzcrNBKf1ftFW0heRjS04d1ttrYuj1rr7ZuGckvzYbvBjLL6
m2o6MuZu0EgEUx59wzI+AcmBHc5rz/i0lnr4Lptkt7V4jaxMWSvs0NBSVb0ULOVb
UT+aPFCMSFAR0Xw9NAw1B6yEVQg3CsIBT4/FRE+yCluBma/m3pkRHNVoEeFaK9yO
rqANWE4LCbTx/+yy4kO+p3t5SevA6gVwWj69uFr/vIh152QlRJRjMlk5F+RoPmea
DvSVUf5KGeY00mLYXpdDHTNTZmeinvKi8AGdvev8xF6MqolmeRYXOYDMG4U/Sd08
`protect END_PROTECTED
