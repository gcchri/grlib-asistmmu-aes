`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HA1BbXjmJ4ylzn0nLu6ywZ8EgMBJQg62UcWAcBPYKfLdfhob7OTLZTFf/Z1GefZB
nXj39sPXBDBozH8FLPB2r8tF3DWkAQmvWD98aGLy6VokEEAZTQsi99hns+nMI2j+
Qab83iV8PfAKDIX6/Yu79GZGlcmOzTOeOdjAjDK2o5Pk+f3DRO4Vqd5gQ3J+1lUS
obmL0EyL+UZqyQV+il4y2ZTIB/M94CM4iPKCBDpwkk15PUlw4i9LjIO72nJU9gvj
lueuGMReAlEhQ+efeNyJLzzaf4tvcd5s4QXtWVoedUxjfZOnoRCDqzQil8ip69vH
i1U0VdbUYBh6bph62OrVSfGjnXVZojxwl4ZiE12wACS9bLNcQwmssS9umVGv4rWM
47Uu0EOMTnw/fa3cIY3QY9MZ/FBtLFpZ7I5zzQ+UJViwUjLY4cyP/Cnwz0/gQl5z
NlwNIbNyMJF5l73g8Hth9/3s66yCq7dvWMz0U0ZwegKHN7dgA/WcECohAD136I0d
8wIxfTN5vd1P023x9Je14jVxnnm9ubRWenvoGInIbwYCJWxHbxe7EoB6cs206aFU
VoB1mC3qHifvtJNqKXYgg4oXca0k/MCOfBRukjh6gAzRSnqC/RbQyCio26UYzho2
Xn28Yd37MozSc86SnkLVZKIflLnGrRp7R64N95KohmAyp8757CWk3aq6xZyfcC/3
agj9UsFgeaqmt5eGrlCULiG5Q3OJlDcelQB3uNEAHnYETBKqdp8mwmvbsFsLUP5T
uSoq+PoYKxYpCdBP7B6y2losZ7kMj1Nf4xFWUwNVl5HncrfsbICCj1R2xDEsKwNn
ZyU4T18xJInYS9Ct3y4qMNZ00ild78F12DpIARoYFyjY2Gt9re+T8FWhQW1R2jFL
Bd1mXf62hBnWdTPJN7rNfsPMdqqRclfjvvMH9OGff6V3lPIr73e5xXWIx/XA+s5F
vBA1JYGQ108Xy6jaTIRMUHjNQnhMSyjB4Fzee6WyfCJWXs0qpDR+7165uAyFgJHu
h5x4ADvDu3Zb4iEGahsbTUqJNPPr/LZohKg7G9H+B3cme57/55VPyBZzGI8Dq8tC
RfVH9k6kQD7q4WH8/Nz8RAHltYzkNIDEfvmLpKl4uDfcnjiYQ+VmaamYeXbjIO6L
tzxbiEQHZVEIMu9DjU/x8/51J0ITFOGlx+DNvVXLtoOs4rbvUQ+mndAWpoQjLN2p
gb0Cb2Ufi8c2AZja2FT3DeEw9WuJYHRIFvhsxGxUg5hfDr+dVwOYMkkpZK6BbiC6
d5AUqnpfInnG6l1GA1uu/JV2fkaZt0xP5fcGfMm85UHWtBig4JQrAwEUd59Fprro
EcJ9WW+au1h7zTFp62cThb9hxclww8wwYlpzxMnBP7h+sP+FTFGMWUFENiBDq/gu
acKK6PHFuCdM4utLd0iGiR4zMOuVbxwT72yJ6BAhj4qX8KvQHN4u5fw+wa/jfEuB
cRUGej6xOnfupdbZMnIXmpYEL1t1pU5FQaYj9OToc54ot1cBA1WHR48PSCBB61dj
d2RX4TRRfE1EW1+AvSRBRaxnbMKV3oGNWKT/Np/ZSeH6MQ0QfZfMQBSDBXietobp
X2sjIS0S1X4aEomuJFo3nl24Xsbf81WT3CLx2m0nEZYCw2cNTBYESE4trVPMdsZ6
POWjNZVgM3CIofd4Sr5luFmOAzuM2MZjfnkbg/VROKz6uw7asJHUftL/BKp6NJob
ivIgRfhdthTPd8Ykksd9sAkbqbfQxDq1BPbbqeYpubennzy/GJ6oqOs+B0ODq8IP
hYJQI48T7pwshWsyQHZLfM+iDT11Iq24dHdna6SqQQGTJFJ7sNV9S7mxtjw6Xy/d
CSjZXnu/Q8dHmgK+dxJcIaulmnujpDLQR4wTOV28RNBC+e7xsktI3Re1SUH2VScl
3BtGagZj57ypIJJbt6fjpFBZqJppBRcZGwOBitk8TW5pGO9f2NyqCLQ+DvDA/zmv
sCe7mP2uXjqxKLMhfw2AInZvMCrPEfS3mMnaoQ1Cff+Es1a02ZxqWkV76DK6BO5z
XHoF7aSlC1Qf5r4tpwDCyEfPy4n7mj/qdg4D2J/WK56rt0xWiPuZR5qGbBvAeGtr
H7ZBuU3rGFYhiOhiVBtqfzg3YhPd77JGPwvw+ZHoPqBOoGcGU+ILDRKmQzhAZIP3
6tEWSPDo+QvVoLqf/bybn1GQ8dX1iH0/uvxJEYY6qbfTMAUONXrtLKMeTbW85lS8
7tXiy80yoK7rg1w1sGifMonxcgxj51ivhEDw/ptbwps92EupJ/E2Rv70B3NdnIqX
o6kWe3N6P7GGstaeuCu5xxhTQp3xZYYDxtrWQ+RNWhbwIR/auv0DTFwNIwTC3WsA
2IJrac4mA6J86mbc8E/kEpCVRuA//1Gzqx+H/q3vUeHMDVtXzCBC4S38Hv1BEVJa
+puiesxfsE8nGhdXE+EDy+uQUl1fecqWJtUlX6JtpxD2yeNu//jzwDlpzRL24MeY
nnIKYUSN+ZfiaQYfXrOXjkPvaawugcT/T1GYekVoKhZBWi5Zim6YPrMDhKwwDnWn
ssguwJC2jQtBt6CSEwNem79y7XgEMihCpDcJPPVVUc6PAmVkbepMJdCdzPvBDw1F
0lYf2n58IhDhvglScb2m2KrjK24bKaaEi3aiNc142pduxxyhJGUa3xGEmNet/fU7
tiu0KHKGYdKeYKnJ3j/YY9p7D8LsziIHcWYkkAnN7+gAJthAuY/Hc7dYf6YiaSwg
cailSvGNSWtl+TMLdRSFiqoc7LnMog/whxdSkLpufRYW5yc5reHUPamKREHW3HST
140ioX832ISEHoSBdzG9WgPrgEr+BRLT9J3BOc5VRtinOP5mrZiXjaJxQ3XkyieQ
nTNhEDAq9sC2QCU+ov/zJizHeFRCCD2+8KvsE6V2rBfhksG/pgxcC4xKUr85T7RK
C51dPPfB9X1YxFuN6CpsKWcaIho0Lbi6HOXiLfAV7XZcbU9VyW0BZ3hz0rHtU0mu
GRerVUEvuxW9p+3FrWfna6+NFS2G29MMWSFcJWMQF00SHxZ5JGGcSjJbFunOwUJl
zILF76mTHEF7xCAaiy+ZF9dz/+lLgTZ0iqOHXCg0pfrcWq1u1QyZ0zxVmeTNdwC2
Vd1PyXJKBFQ8S5Vwty5U8rYy5dq2Widah71NUgl2L2jP5wudAdt7BguDaeDQSnMD
RyVhyxN8o3jrV1MmJPyxyyW65/NE1GXBm1FDL8ryWv3vuxTFykDUaIw+RxVHAKiu
tPZkeho/zsq6jhEWKAEYsEsvLqP6OqI1Il2lbZRyX5k5/F5SJVQKrROxXN4jBC8J
C0nI9K6T/QSt2y2uVkCI5QEBtpfYvfnJGSMTguPXVXw5M40dOrzEXDtyZw2SbDHE
0Ct2iQCY87cWFmDKMYG9UfE48XVNMLkfiuJBHMwp64spMbT8cIjTAuWWhSaDwnQ4
+CVmUk5ratLAfphgx79a4M2aUTily3QAyIagiCNN2SioqbVlxnmmUVMV0NtdFeaY
BUZwLFmCOHYMD/jQkd3U9QhJYVqDWVIK6D2Il+B+jMbfYrSBy+pyYcSL4mgIK22W
DxzNG6KQpH7xpiEBqCD+Aj89EzqTMWh9U1lgiZtq3oE1bTz63dqzgp8WPrgxeTh1
eOIwnkaGUyJzer+kFCbuwVFbwRb6KIDlPGXTrCtRdfGNEvlZ7/mSXeGsAzaVYa2d
wO3m8//ilFMT2D6zmqWI3fJaxEcWlR2Q2LoYZdnsk1NH7fk/IDHXrd5RxAIIpldN
hPCVdcKxD8d5iRDXvmJ/rj2de0lEEvus9Je1De6AGdeUW2BObMUak+dH2xtTJjc6
sHMhd6dE8HR0pBcbtSb3uzhp13Xf783+k1AF0tpH6eya99FtvyASqFzNmUGs1shq
lG8/27ijRYfCVecOn/m/hxEGjoSd7i0pTNy+ktOUhlMeaMmPnK4PlX6y4xg/4cTX
Cj77y81WGmOnsyvrMXT7nni+0/60D4Pw4Ql1xDbzNIFS0bhhzh5iNCXtj4Tg8bTW
eoqEPJfVkUqjk9dj0Dx5r+Di0wPlhnOXmPSRd9G137B0kHSJ55gulhbnvyv6JzEW
NKZF4jlvLy8EYQXWhm1Iiol1YSaJzdDRGgVpQscEALZT3mkAVdZ8W1ycDauwbi9p
kCpoRXbR1P0JMDWfhEUFzIcVTH4HaiCULOkHHoe9RHMesmCFHddQgvObAaPJ+PKX
s9Orc4xWuWaBS/KVYqQ/CJJNBKI4W+fCtTW5rTWRW4RSUc95SfdTPQ/Sv/Cka85z
k9UzhTbtnl4eFGM3Z78pbwmAvOanmWzT+f6iUl+DkXmPY5biBuVvPFJeBdsS0rPl
4YP7eFwL4s84RgP+BSCC9dnh+5bQlEC3OZhKyM3jghab+wtE/be0eNQtz3VtYnY6
j4fAZXZC5dwF3rZ0cL71IoDtd9lDetfC4v1YszXqAduynUysIzZ3j4QWs2Hga1Qk
AAEne+o2GRaKI2kzn0zsBW1wT9sI9Yd7wLZgODUmoDY0zvGMbQtR+Vy43iVPj/lT
mRR11Z4NLptWFQ/Wmsco169VSjLpsD+h+3JCgUKWIyZcY9GLvGopBaHmliTjAV5T
yC4DjAuI5vL/IDQeonABqVJqKgieY1INI+g7AnO5q0W+q1UutKm3XKa0vXBMm9Dw
rrZa0lNA527jYrlPUI5XoFQZXMJH5TydBu4MYz9swnBBRDqnzNOQVyNe2EKmzKXi
zwgP6PJFKOvj0vzgrWS9M3HmYp+th7r3zbF/iSAURprD0tOq75p18PCpZlJesCui
oI5s7/amcJaPkUuDAjoxjM3WtDX4kRt/gUUCg97RCi+pTBipMiQDwKaZ09CZCwSC
Y2a9snyZfPO28OGYyqCSzoi5+mtmB9dOnjPkCl/25RYkFDwjJjJCQf2uWxWpZJHJ
hNVNAtb4mCLXkOvbNxPp7z6+kePsNPjSAmFRIHmYP4JPauoVzLuALcknaUJkac1f
DxkuSJnk04zkMb9k8vIVVBx/Zzp4o6JioCvafFJt3mSfuWn1XleA77Eu69j1b7nh
anc6qNrHqzIehhB2TEb+NIn4EfHc7m/gzFygOXmt2RH27n+eEb755cSJa8AZZNTf
Vm7A+xINtXT7yf7ulOz2gHC0eZWE312k8RRODYx7/J5EgzQ53LBfmz131WHWfF2U
1G75EE9SbSk97RSZ6VL7P0q6FjfI6tY7FIn/du3TJv1V7jz8DXRvv1nMmGqXO44n
UORnkvxP4jRLIUDDzQZUwQY0fusV4NCfy8Kpgh4SIv66xosN5f38yDlygtcgpfoI
5XYvjvHCto1J6SVPN6rJY9OQFPSt2C0nPft64QZ9Ds9EMSDGH5ma/JR68WOQxKJF
fmBRnK1SWIvmxCiqSwPnMoGVJNiPapcltYVMy0nBgEN+o8OTIErq/7z2Dd8nzoqS
UQGC3AYLSJZ+Lgpp9SPC4vnmum7oYxHTpNdjTwQsQkQ0jRSFsdPLqtUas7m+o+xm
Hcwvty0JANYWz7qvZdJBZj1JZR+4EFSP0xaiAhEx9W63NBwIHezTmL52b7wrnbkE
9bkFSxLqU1l2ev3SFlvs6qybwnPG98zNA3/BkMP1/BtIGuhumPHrluepxBNS1ew6
1ja3qRF8tLNSKnUYNI+cIUmn48lK4ottCV8Z5MV+btAwJz8yyleAkz3BfYmiG+HY
IB+drmJzbdR4h7+8nzAeIo8BYhkVYLT6f7TaVYKgOm+L06aWtwq32nrKdXV1szXt
804DQImMP4gaRT0KuIlEvgB1Ak/RrQR+Dym+m5Pw2F345j7t/GABI/gPIFzQ5JkV
T9EOq9KmanaUn/MUdDzi0XKbXwtB1Jw4Gr319EW/FUgPk8Gae/BMVy5m5CAYhPfs
+PM+WreS54pdQtFXNi9pMTU6KXzSg/i8m491TOsxruh+uYLD6Ob5C8xfgtzqjMPt
sZTbTL2zyY8iCwCbIMYfNmMHDlTRpIEmHtYlHgAwtrtaG8aWhCizTrvcb8oXVJX4
GjjkrI7CHvYJgnKV9UtK19N6EbtLUH7EyDVuMe74/4MgnvXYgiObN68AfgmcR/29
1C8YE+ZGn/M1lhF61fCxUwq7h4YXtQmhUSIRoLwvR/QHouoBRSDtjn5jNZ8FPogm
fZRAgPXngjbuuzKAyDF7pnvscs2RhSJS4d77aqkcPMbd31k/tnv8947THkWfzcQE
NsoyA+4FBRpXq9rzVTMS4/xpGknNSIJVDMvO+eEWdY9j7l5VEzXAMPxN10PCO+GB
xwv868Zk6XE9FVdxq1Y36r6VIXemJ+YNX/tMyx45kt6rN7I0pak4A3CXYBvpLoVV
mSvwzLhnOMMeuwsAE0fZw6fLvOcXa0qc6IrJsEIvBHXLVQpnitlrub3HCjcdSfpX
JX873HUYAbf+xoCXbSSL6hmPVKrtvJi+K+6bjTHKK2aJMtFvwNDPklSlPstcwM0V
Wxo1j4ZFg3nFvcMrEU7ruvU5lcgAWzH0y9doxePSpdH7O2OSSq1DW8HRxEGyMs2P
DJAwmhyLIpptzQb9k+sqLHSHYW5tKpB9GH7Lrh7gJD1EkvdQqv9XFJiz/rB63/6S
azoKalSJ+NqSkGr3J9Rmp6+sNC89ciSRNy5obOKicB+a6eeK5762V4iLc+qY53pF
7TsC12qVbhUOwcDksBM72GHoy7K8qYR+Qe0pw6/DAkFL7X6ZP/y4yA7r3NRwxVuq
A+RjP67t/QJDhoL8vKXSJoVQDmJJJOvqnFLQuLAuPkEivwI0uRGKFXHu/xCnh5Ud
Cts36yfGbIwFyCXmkNyjq8gMMXevAK0RWSNkiJ0DunBkMBlwReUl1AHwguTJ68Nq
38alrEcB+wQl/DGWeutDSGHOw+0YpJy6zsvxf0ScCyGGtiuPcjoMvlxgnWHdK+y9
WJqknHooMHCIbFCZMV+2+KrnGlusb8a8DZwQVKvWZDuIVBJm5ufnqZ+EZqoc/xKT
XWdKEyayb5axVpj0qWtwkafoG+MM+4Nsc1lR65yYXk+1CpUIU0wOZLKltPz3Xwju
3z+tTJdJR/vEO5Y3tSocFwX7GSE5AI0yikSVAEXwVpXbzs64crrD8b/P1cjB5HDC
KlHahc9OfZu5F3eS7z2ubqt+s/9b8o74r3AhsNdWvxX8Kmrgbta2ZuMCE0Qy4n+X
Nycknyw7uaJGxBtQu2qGISI46SpI4FYmjN99XeK5VGU+waFRjOVbcqrNpjDQeWFk
x0pJTU71UICoMipLA+ZSK9Dq3iFXF0BGJlr3IfVaPOGQu+xWt6Cwk9C/QryrdjHw
IXGCL40xafxYEWvzkYJzMcvzIiDp8l1tQ1QF9NUxey/Tl39qqpro49TzoR1b8Gr3
WGAr2F/yr/iQDuZmDbkas4qwxzrdHhOPa4su3EbPJjonIJimFc/Ot6GKErDXfQRq
hT9uQCux0H1LatKpHZbV330r8GG6Tm4Obsv7EJB4JqnV8gfvhILCS7SvbCF0UtGH
VJ/WVMZIFIzVO3uKMYSCPrjZEGCq1+26OLCIZibWXFuZ0U3s3qWbQsFs85NjXRJ9
x6i3h762ihFo1EOvHLIM7twRpeudrnp0PDv5FwsLv8NB+tYSHAphLeikR6wGaoY7
E94wnWTxHZjaY6FOqt18diYhbEddqYv5Mk6/aDRyyTgoeoUpoeimIcWF0A1ek/gb
e7r03mRnXwL6KR1TCC569+EIeTVsqKlWY2//7plHA365EShTqAKPh/F01wG5u36X
gva0eqa8JwKLIDushO6YPDmJYCG9M2OAfeuOUH5KmZxO0BBSXDj1pg95A2/ld9U+
tHQmP2RCXMHYd1mBgRKRnZ7skkEwsx6NQZDQo0pC20wDNAMv3oOxxM5Z7+ObFj4L
f+259wwbQs3lA9DsJ9+U6OZETwuK0uZ6vNkt0ROXrLHl2TYWLWroabSarggN99D4
hox0c4BGRaO6cgY2V6qVZeqpL81mSelRh4ee9f9zUGBPSrmrodJ6ZY+4ow8aweiu
ZaWzoca6/uWMAjuFGJ/RJPkOLxWmv51ITPjoT5qfcevCWBTxcgU0/TFST91WB62K
ovUR/zYiIwXNCZTQKvYu94pxbO9cWu0Nnz2fP/ZvCDqgIyxOURM6K1w+CE8eDaef
EsbtQ4nRTbvPm6Q79VPie3265eN2ZfPCyCjRGXO0UNqyFkhH4k99be+9zz2l9/HC
tWKznWf9b0nTMkdw8GV4OH1zEYIi/KBJi2tbTxszsrToZX76Eo1EP+DA/D5pdb4n
tziewrRZ97bNro5tXec7tFGnJunHSZnrLOjCTLVWVFeHCDPAgI5346WFj4vCEkM5
hONF1I78qEYOeLwUthTDoz2WmIXC/+eHsppICWIR4pZnxRoN29TQMqd6kAOPH9rb
61QZf6LDqaOUlEMtFLDBehVZhFLJuirIQqkrKs6xSLriy3FBYFR5k5J7dHWGr84l
IAIk5j3OfcqGINsNNd9mZpv3q37QHB4lLzJ/6Ai6tEZP1pTvyMeEjVo7q0cxJ0h9
jDzLN5tNKA0s4A0ocJNMwvBnG/G6ajWkXwFAUew/7F7mEhiO4nz1ObVvdp7ECJS4
d0NF7RIK5lygjI4Gb7G93D+AWjImjmfM1bHtLnXrdjtb9puayAiA5oq5zwLocefh
9S1Lzaw8voZVfc77/MUHOwGc6Yzc7KxeL5E+u8ZMyNozcl7dlegI0UIQ2qlDo+zo
JCkvIOtt8oxJrt+vdHSQ+glTveY7rJSEWIQv9lzsy9qzzPqe7O+d5zBkynrp00eN
VB2NeYp8BQA1xZvV8ke07bkLi2mLRNkMdHvF0BkPS0HOsszn9DZBtBn7+TBif1Ze
SIZEMLAOXvi1iduFu5ZoCzotvERajGq/4okYPP3SLvytVgcSRNk7zDS+hfZNpWny
51NYmDOD3ryZubDZzz+MihY6FITIAlQMPzY79+Qk76Lw0rLcmgRYc1TGQKuUR+nA
m4Is+vEotLH9lSUkoxi9l0c+Jc5Iu/Vn1yGum32kLRsuHWhZ0IDRIJbx3x5KsUh7
1dz2q8m0mVCYJacXGueZwKmkrJV3+vTqR1knTh5Jh/kRYb+GROtfLqwfc5StzVdQ
Ws6fxFDrDXJHIFPJ3F8fZUfOhzhdSBes6ppYpoHeEqBQ3O6YyQNqFvQEHozcU9U9
LgJIAUHUtvY/6XKQVLV/cuExIgOM1uOXPB1KKAa3eFcf44TBb7AceLaYvZgaA+7O
zusoCGmKp8o5rm+NqU8ZYRo8gd86fdwd2sA8XXAVw0wJEMTAJeoPSEbTL6f6njSM
Bi/KnyR8wfNpbhCmsFvG9BPkeZAG2vjGzM7rnwE1QKkI5HDmXC8RS4U+djKuD25W
+JleIpq9TWNP7OGukxKILxMW84HPwi/01eB5mRr4wieTL6CQNbwUSMlmCRLL5Nfl
g8ZXgWpi0fvsDy9BgM/so5wWLg6GMDuuCPP1STu3fpJCLCjFq5iinaQESNwrdbxb
M3Zoejbo0wO7dmgOUTN1nm7uLpriGsrwL8TWy5XV1rTTevvOFJwloCwFohAn7tKI
qQ2+8xnnepeSqVLJ30eNmpXDhq9BM+HqrWSK8dF/x0XpWc39VfotDUItYewoy/It
1aYxkl4523D5FnlsoYJlVAjYZBx4Ry8cHpVez0v+HWNtmpuFhU/mr5ewrjVglpkh
Hja95THuQNM3JC51ye7Cn5Fqvz+y40pEvzw6/9gv86zQQ0BYKS00xEHSdmH6GvQH
rOjAA+wCd1EDGpbIIcuqKNEJ2uJX1xjZ/w5t5bdBo8GkZwmvTVRCqGUaMev2YOiA
C8p+yN9TSKbw+SEGm4xkdiETbXZAjozKEZehy/dA+sJA0+k3NSAZFAlgpvbu2ltH
iIPkHPvHGdSxPzcOod3MhYJ7TSdS6vPcDbi5Ey/7sqc2hGvan67pQoSqrTZzixSr
TFiETdl7qY/TNBj1l+w0jmN/8l8AvXrsZJEbdnVcmhy6xkkKBieDJDMKbhzR/rJm
yNiITHQ+kOaw2HSZ4sinxiqlruUuoj1xePymvEXqcVRywBCf3wtHmra0BmcK+FAX
pIZdSEZg0bZF42/a6v0r1edMIAjhfwuvKSbvPSt9bRKuICTD7D1kDd50OJ9fS52a
CjPRRQz9nq7etQwIJMU2fcwhTtwU6q16NLsYMHnEIZwj7SoO8WHVd7a+FOuN9mjt
MzcZZDvTG63giAaVOwCCVmA252Fbx0V6iDDDdvQ+hrb+quNIpNFy9FDjwV2I32Z4
fJg/fQY4/u74ml7C8140txvb5rVEbwvgKz0VBj/XcoiVCm4HYktSXVPCaMx0w9e1
BM8fkjV+8XG6Y8lMp9I+GjTmpDVajPgR2nBpfk0A3BUTKy+4Z40enAKkUok8+yaz
hmy7jY9c2rdNAG7H0OM/e/YqzJzFoPeDOse78g+Im71bj3SeS/c2VmLbDc8/6QAw
GYeRCDViWW7qFhkZUBWsfLGFHeqHYYvAafADwg5CU4BHzZFW77nEhNHfyMotP7+4
WAtzVqfxK4Wx0BYEiPh1jKhHguE76qQZ62GB5/Q2r+93z0TAs/YIuYrJ/RDdqvPC
owWa17uN3s/iP8GbVpsv2Q2dyQoYOluI0wt9EHdov4l8MEReKC4IbbisqoyQjHWG
HLt7ggXxMKhrRJIEDOUqocgiSSgLIU5xEuniIm7p7dEMg4ELwb4YqOQp4gr9mVFL
h+o8/SZvhTj8FGHB+gXtkKlJB2K+w4Q1iV3Dwt8DPGgqK/laHyYAznTmkubqRj8W
jzdAusjBNIkV/i1oU0bEiqjbaLW1LGcK26g3NofqdCreEXiRUQ1iJUz23O+pjTyN
acm/o17XoMU0+WOA7qL6kOLPqQtnPWaKeHHRgPK8BEscbEFzs3VgVq405pyoOKEf
NVH1bNxK3OE4CrryKOj3XSGvBPz84dkYa/BYotT1/rHPtnSEN9ukp94j+p5a/TzA
hyC4nmEVMW4dKWQW6Ktm9Lciv43eMDaiPnL/fq+1KUvMJCGy5zLGC8mvZs1zpKEU
WdSAUROt99ht35hGETZrV064N7x6eO7tsxnAcGeNYxffEF47CMBqjZEadNi5Ex/Q
0yuUrgpKGOyD0M6gOJkZGHcTeSc3KYFb9WfyYPzqRtTx9fpmTaKlZs3vH8Fs/fKz
ZtS9t4f6jh0tI0VZVtvUBi0+tq2nNfOfCGeL4r6oTBdXxbx8mUbxC9/sZhxIR+lp
zx9nxi5aBpaBjBnJs4if1wjmSQgz2wRpT2iDcsmj2ez9oqRkHPhtljW4nGZSw7QK
KknBtNrXD9Yy95nnX4mqR0e4XGmlloOJsAVzKaJappG3Cal8xtpUWiy2jZmfh9Ba
0YdNQPsOfVbjVEvkyx1u3zqgIpsvyGtyzaODTYgAC70o4zHmt/R7n35U3BE5l6uj
svaCYWY3bz2oK9PpJTtj5vP2tlIhvIAvIqIXAymJlqASHj0W0Y2VWOapwv5XPfTK
48sZPq4/DEqeYk7WaPeEYIwqi/iUfHxVyOeBJDod3a3SA7hbnh1usf4RBWB3EL1H
Iw+/84O3l3reNYhi8ZUGcem84ARQcggF+WAlzjiJJEofYrUu+pSjyzj5eeEzg7Vk
x2Rz8z16srKIBKVzl2PI/JF2jSmec4on9bC8f6uZV+rE/FhSxSCrGarCkBMIIjCs
QLB7ibFMIt3tFOy5CH54VqMQCFalGrGPLFqvZMgPkTOLAkO3ZtiLrpFYhi6u/yOK
v2Z9KUWNvQysZrDr/531iaN7TfNENiFzUXU9zF7eoBt9ea/OeCaEZFKvPzoWa2tZ
VzlIhzGLrCLp42Xj+UVCDqOOjSFPpbxDfxcwC+I9WzH+86CkO8SQYBUnefa0TK+W
xcH0wikIimJjPVtX54O6Pi6nnyz9ArZnzamh00yQqS8VBBUSltls/jpF2S/87j0B
5tvdQkoCsjEICyHq42q1DvLAahqNCzyV7osX66aARHBEzNond0ECSrd0W48I8Jwe
qbiwMlyzu0BH+AefK9y2WDs7kvnnTx/VOTJsndsHDQTTMD2EJTc3sIGCaxgTC0ij
cU/p7F1YK344b+yWQNGH0Pr9tTcQBxb+7qF3lWCITwu8etsorH3fQI5RWSCvzFs3
/AetWV/qiW9Ms2x2ZJ9VmBXFbNm8NQi+P6txQZXZLpLxk55QAvzwfwCYViUVMH9O
LODNcJFiDK/ViAdapAgJ0HUFkmHzyf2lLEQTdl0y8otP1oGDPgbkyNaNK5ysxqOm
gmaDIUjBtxON6g0sU7wrGbEqbky9x/0AsNhpPesVkB5YB0fMchCYhIhz5/giWVpJ
77j6DdO1FCd7/L5l2pikEAEL4NFffWwiNR4G5+S1GArKTgV8TNhlquZSURUbq7zo
Z7eGuhM1wdbIG4IKh6AXgubrfkHUcTm9eltco6IeWe2dqPOzJbQa+GQAu0MrFZ6g
600HBOvJBtyYnkR5C5ngFO0Qrnn3hMdE4Ttwm6XpVtqP40k+0M4RfsvJjlrzeitI
fZd3/XKrzi+X0k+DzI1SWY/AVl6TcCY59f4iSilDmBBh4VPMA29SVRjXFBDyp3G+
jmrAvB77eAuL2GtGEXY6gS81oaecYPpKUbmk/UBQpiHhdaow0nSHrZIHyE+XRyMK
1fDyOLgAGkcnCoXwtUu6WeYSq/nEEoXTfIjdSMK8K2aKm42fD+/jkGwJayVCFPVd
Lh7i9NrWMPCMifxutYG7nkzh+IGxjoNRqplC+huyqApoWxyRKIUQDtX48MviChGy
4/GPXWy1OATkhURFzyY+ukNieyNeOtZZxEmVc4uE7FNbT9IIos7sfYCRRRlUGxom
4Xjk9ASzpViFR9qcpB5FVrk1ZZ5pvUIdXw9xsvF0YO2tQEwdSQEP3xcT7KIzU2pc
8ptdgKqZZIZKxjyy+YUGXVBGPTxrtCI/AeJ9dHqsS/HPLBOg3erbSc8+Nyk+SUrt
igpJm+kP6cVO2aqJQu8+On/818o1zvVIh9g3DXNc0GNlcd+LYB990nPv2e25EZX+
FmYRAKXRR8Xo9HK3N0bBK7QLuPtbQpNNpOWzNvluzt34oVfEOZIB+h/kurkGyxgK
HwZgpWXtHzIJGD23lgFqroDWqvaJtnbadPxSTJCULQglUfj4f7f8KVENoUI/hKYe
5mDTnCpWP4eM+UOslZ2EtYDOetdTCuYRWcBv15DgS1pwZvvTLY7V/4zORAbbUQEC
/Arx+lhIzyn0w9TUkTyvuCzpnevb8t/K6EdLRlZtuU7w8Oew5+Q+fH8RbPPEtPrh
QIQdltSsD535EOZ8XEwxC8GZ9CQIDIEu8a5zJYzGBJLn+K6bLXwv5IDgKfmtmXka
35EDHmE8lgwtoHPCxSG5PdOZox1KDngBgAEoKgbyfUgZVHTc++kBGTWdcp/b4DQo
T5Mt39frGUBj4Mr4FDJTmFxzghalztH8L3SIZo1WuVxfyUu0uAoNT8ua4d/JLaBY
wlMRMKNiZUk5gPdbMNOmXNUH4N4CrAHgcyCl669ZFqa9Y7zfxLTqci1/tPORbzE0
iTEKpbtZajQRkI5lYT5ztm5l+4OM4RBzMr/DNDaSYSrNpI6Fh5TPHo6eMYWyuhZX
DeHYe3zV5xbbdI5+puFXK/dZEOKSFDjiAB88J62yrUNgbQeq91VVGNM/TS1Nz1HZ
DF/5jhK96yAHonwprmWJ5n03zBWLnXt+UKW2W8tO7Xo=
`protect END_PROTECTED
