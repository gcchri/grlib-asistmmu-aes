`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KWhKmQZFtoxWtlP9p323fqh9sYBNNHHTi8ByyrUoGctTolfW7pzc0+DQzpNh8K0P
mrr9c3y9bik0vCs/sWBD6OGk9Xp8YaSXtJ1YEitQZkTH5vpXFY6umtHKqqot6woI
xFDPm98qH8klOn1M1UuyC/Lk1QS0QGgctyKdpepDZrKPSkBfL5rBAIt+nlwIFu4/
Ix9MOEvdEWvGuVsZcVutPGfT68ENous1jNwHAueI7oCcP3e1PyVSqmLawER/lwyF
OIhUOhszaxNWDayijd82mHHtyWvVGG7E2Ekau0eORUuFfyFDhJTEIpLGAxIE90Bn
o7dn9n8vxyuUhmk8DKJYp/TeovrS280F6FusuPiNciGlgSotYaNc7ynDM0gYP0yI
XaYseY0qTRs+rFKqUMOOct7IX5y81FcZFlJLWBbWqUipGZwE/VyEcK4GcKI8VUZ+
`protect END_PROTECTED
