`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9NQZD7mdHSchUL3kG/QOg0BqYCj2bAkfzLKtkzygL0iOkf9nyp5Z+iEkwoqRa9Q+
Gmqhw165wI0y1EUSZkHp6LOvmFZhdWLSQ4Cd9e5ibfRzyDcfemA759OwWsS3gdqV
nIYzUJacg8KT5RN7Z9u2iCwZbHJLgbNHFCPXgQCpJVMI77fNMfmZ8m5btTah9E4A
UWDTDcU/bRdK+S6eZ1Lr7SzTA1ACvxx01NRjZdSA7yFLETcSjIOwLXfS+3+flDzc
04FylTnSZyR74sFdYsQ81w==
`protect END_PROTECTED
