`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f76UpcDbSGlZBarPYQWWI7W5nuqHEFpOYqExMkA4jW2l18gb9onbOMQUYswqqwk9
EAKcfWTCSCP2wtsWqL72rGsZ9vyxsoQCKrkiqmId31rXbYhXKWFy6jOZKPBvkL5c
KLudpdSI5YyPdEipHLBCZBBgCPgWRoydfkU8OkMfHg4N9tgaMmvcX5ACETfkwl2K
sUQgl3YJ3fjW/YlgTAqQ/daa/wwsJeEXlFgvzQ/IWClTELJoU0e7fVXpGnHy2Ihz
Nmb2jrizBzUm5IPPq587GFmaJE9v2p/6XGvjPpffsXL+xds8Yg4GFEq9NXPBK9Dk
vWZm+EISfiqQfpPuQ5IZ4joD1rIbuxOsxkGrOwfGu5V56KXNHBtfEMUyN/E0knkJ
E4Djs97sFTfYl6ICQsLFVaRbbzuNIAM2l86GP0uIUh/W4aY1D/v3jcUoyWAZlUzd
OTVFlNunhDQ4NBac3qS5as42lvbQ9UcpL0NGLVDsQ1Nbknc5T3pMuFQIU0Xyonn0
QYCb2zuCWOZnOSEWwSXooujOmC8T7/EJpZZmpqtmvtE=
`protect END_PROTECTED
