`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F9lGhiEdGDy5uiJjAd0an5AlJ+gpau+qRTw5l00eageOPAoIC3eQLmCKVtPaD/R/
+e73E8cAb8/oU84heWBH1HYVFcoZDtk5gcEw5R2BFZAoCy1WvnKvtN8BjIP5uuRl
JNx6yNKMQg+Y3RDKTMbBYyd3LktcJhIMyKM0lGrM/iMxTSFrTt2haPBshX3filsH
N0krIgOXkltUHX07Sw1v/B4p9gyFsEx3KB9Kc2atak5lHNkXCQEKyTdk1YmM7ov2
BuKn4x9njqhYR7BmErj+NjLsrH4poggcOv54RObwzeYRnwBVw/B2zyZFtWl9O6tV
IK0gAAtqCn9WZFcLQsOAqyjZETBPgKYu/8dfzuDORgPmwd5lUsTddN1uPeujb0EW
kEorTq0xlWfQKiLbs1rxRg==
`protect END_PROTECTED
