`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A26ImeGC8BQ8ix/UkAMDumjOs4P/Up6gtyiGLErgzWiCvU471xsZlDpWXEXpi8H9
F9VuNaD/1hUXeRT0GDxVWAgDnm/q5DM4UwvM0wRemoLHP1oPN1RX60aFNwIL9Nu6
bDC1nlxNPWAMSFTg5soMEmyA7FtBghvxbV0ld4q92rmvsjYcLX0efZm7P3js/zrW
/MbF4DjSw8WH2owbIllhqzcsbW7yz0Zxom5pYYTq03aEF5iEh8PnFR+zB0sMNNbA
/jzDCuXEFe4EOu3vX0ZZKFUeN9OtfC2w1m56Zwmv/aND92hJVFRXCkipcm4pZhAy
79tfEyhWQnkdT3FzM2CKjvSiknVKsgQrg9UxU/IlsMtGLBlG8iSHsE2lEdJab8mT
Gq5GK8FD9Fs7csRfqVG8laa3GAX9iNleULMe4a+yMiwDkj7A/h1tIrHluXt//dy4
Z61QhPR52OkGafzLWlWu376opqeQuMI7V/xdYAA0mOUJgu6uvJ4gnJaZw6bLAMFf
1Pzg3jH0qa5QFyJPRtfOvfwDbBo9srik/Dl8iRYHc+QaYA9f6FctcfPO3mEax36W
IXn9MzSheusl6Bt2wQoRvg==
`protect END_PROTECTED
