`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+HPg/npRmFyyvzA1l+umQgDUUH3Mj79n8HN2pRfnuf8Gffp3s2DbKPG1jH9vzfMv
dFKCi9qw6JA1eXVmOXR1P4b3fU5I8QD0xBiBSErHFs/ccmUJhiyYHvhY/TK+QO8m
AUxbMGmj7XYUG7+58HkeLk3x6cxIjhXQxAVk7ig3FiUpmailRBXjZmzhSpgxMzOx
+VkZXEbbOOztTXnGxYsQPzoVMRLnjSg9z5pUuqMxup19HkPsxyfjQG2pJp8KCu64
+q9NfaIz/VZTpjy/yoT4tsxiAKl4LEDxZ++dlAuBIrnjI0fHPs7JLK5oEfyM6DTF
aejwfUNdS31ldd41vHqtJooVZgmRt85LfAA7rrHsS2BKWAotGVwpzjepFaiCRtnI
JBfEh64k55Au5d5svQ69GJZL0YZRtOt3ZrIgNo48tg12DH79rVH2I7ZL9MkxPRF8
SVc+1JJd4vGPuR+sdwThB/O2pvbaesFXfBwauuWz69MuEj7nZ6ksFDK7egMHhv2K
vp8bVveWaYfEIt4av1oLY5RHL2VofgmDRmlfS11/ehpRrnHbdhHedoPQoFCtk2Gj
fkys+f0yjsI3yUCDEpa4OD4YPn9aPwtCR+LoAXCkBWb11G5jOmzhxF1/E382/2LN
TrYzBnYm4/D9WljmotJ4N+G670tV5q9P7yTRqsk53WCKbNWihKhRyPj6g56tHTOu
cU9XVtEP7r0D/vIeUDyVP7M0oisxcqi8qRlPL552bObwLPYr978OcUY9Ajx8vk0W
p9QlOERfSouUX2EK24CIp4sOmNGNsSIPfmh2PVbzE6cngwM13cpqOQ2O8dOU32um
mT7H6hyJ6rpMn9n5GjpkzvY4E9gMcvf8ZAGOlo3tQzXovH4XOE8/q6x5n1z9ZMq3
cdoFxt9wlCSwBh+HmLZL93EJmfxWqUqMxOdQkIMLaGk2j8Un00BVB3vomCmuh1H9
dtjG16g+mngc11D5G/+1goyBDgQbRyvD4q1NV/xDJtdu/iJapB++F1wpRRzDGV7n
LtbMD6qIfLn9KEJTTcYKxf5Uq4Rv2/rdAKDqMHhmCSzizc9a9OwkMnAd9KEy4wwY
RdB1sEWFW8qpsLr4sgWFjPLXy6HGKrCCPcJN5F33mgDqvyiq/MDU5GOkuL/TK27A
WmDtIAl+rD9XqMTiYf5aDKBt/QaKdEYoop0VPTzrgjtQ1jLKrnMiZvmVPDGevK3O
2cs+ElgFHmkHuubA+XfisZSkp8/2CRU6SIMkf+PB1w/4PifNJPoZRiC/M0Iy7S9b
BlYcHogJlZyt3FRvgDfvyTV7pxiQR2FrZKFQr1xSYE/6xj6FP1e8H58ef9BBD955
WW6/ZKEB16WmHx/E4fjOo7xKMLzucuG76l3zIkaXXqYSQDJOxL7uaGgy+n42kjDp
F11Gi0E2ADKYvIGXUueqEk5O+9lABK+6d0w/5h5DR3svXBv3gDXNmvgvbOm6qGQF
nw67D00e8pynA9InGP3W7AAY2qvWZ7Kzolnd0QQTVYQVYD/jsbkql19Bj/KRQCV/
c2TqY7/+ZZ4X6jUzi+xEdlcXaCGCJy7VSkp3iVyhu1E9mRS1LX96ZIwuny0Oc1iY
DQkwi60d85wsUtzPC0lzIdMxoGuFtPsPisH0DDGtXoQo7Vs6lMCG1DJ7kxDK/A5T
PpJTZRl+7iE16MDPu1PKon0CVnUJcQT6dM6vg14R/GNx7d/+CQ7YGnA61Zc9kCwl
ayxQ4z0T7Fk/kL2J2Z79ptOA9htya9KpPfSqWQ1YqIV3BLoy97PonTk/bbPbmEQu
B9rXDfkrvLeehm3zoV2ahzKHbc4Coeeic/FAjzgJxBH1pYmitGKO6W1fccNTYve4
J82otO9C8MD0DhVp4cBTDxG1DGUWGXxYkAydR6WYkbbtQW59Wk5PRdgPT6o4i4mX
JyYDVp4hrtqk23Z5VLWiqZaQtgSIVEHbMV/nNiAz/jCCHAALX/+3hlfxOSveCaJk
XpVm67n4MO4mUiAzrD89K/IMoWQkWx3IPU7t27pzTRj07YbPynsakMP5MxVQOsDs
bITv4GH4uRMLL+w+818xoJrU5A95voMTQcAG49E+xo2DidK57YTmqB/KOQZAKYnr
htnvYX9M7cimjNzsR9DfsmH+HTvDjQbzwNlrJ6leJFYcgwEQhKNektRIew0iDcyz
mCm+FemZrZRx9L0lLm1pXp4SnFmJ5OXU/YTIcilWQBAA8D9DKNijVF5iQK4uJO3R
p8OxveJtUShKHA3dUFNV1UfCrhE7Lq/2lXsuEbtyFb9Z9d1L5RBuNsmpinft3Jk6
vcJDRWFSfwq1/yDZydyhKr5GBXhyMSoMEkOVRAjpEx73ifO55IvZ6XwWT6i3FAKo
vY1EnkszIaNdvIKfTBpEv5gjTIYSKoMSlj9Qx6nWjoCakg3Zo8HVWlBHwAZB27LK
iHYb+D5iQES3nVSvQ5vm5Yl+haIMetafpkp37EWlLh1Kylh5I0Srs2oOsbHayu85
RbHUw+hMEml8TQqgLbweb5ug9oU9ZAiKj6TrkqZ5BDuEX31ZfElzqXPJ+lzfAZmD
hiKvdtRXRpA3fUpcEjgfv3yTSYcGKRpyxRVFuqk88fR4pej1leWjMkCOttDct0mn
Ipz2ELHJEdff4TafLcDRV8WoB4J0G69IzroRE7oKVNMAuG3EzAI0xyPlZ1OLNTG4
ofJgCl4SyOQBxHqLUUniZV7EDADGeT9Y+mwB6o7Y9jWaU7UTuqbpKv9c8JITC2PS
S7BYHE38lEMb+V2+2ABG3zqPMDg9nk2smZFjil0sjs93//SeIcEO0ijhxAZmSmZ0
xy1OmVT+ghMbirpwSAFc0u+7pPA4IPwmRTteUtVInQuDZeX8VY6hecrar49gGOhp
JXcjajvNOpVmfBGX6W1GmQ==
`protect END_PROTECTED
