`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RW93xFOogy6Qvg6AbwglmGE7SFosI3ASjw7e2XZm8hdVSEtTy1tNhFOD59ldWVHQ
uIHpbmouVAyRltPOVHlpNOyrM0zfGINsiApQipC91Exe1wR8xwKbXSV641yJiu9F
/UZwxovH23LdhobchcFhCbwGu2+p3VYn5xHDWn9psFyJJFY76tybPLCqW9gDhxh3
x11SNZ4kD+hGSZIJY98fyuA6HW2hHjkq0OnBkfCVhMjFVLj7AOQfUDM8PbD6+mcw
pWeNl9uOXSNXirVmwXD0iifkTRq7xq+Wbuak0MrR/8VA+bRuqfChGFAVuWtzkeEf
CVXugzuqM8GCKbGDE2AqAvPfNDgEPlunqy0dFigO56qtLolsyybJsxmCsbNgEOHr
YJQ3dtvEMrjnUCAGuS/UnUTVLyNsdt7MwC3xPJ4zLIul+JUiPNOBVjEtvT3PGG7A
eGoOoZY1rHz76TU70l2QelIvo7WjjEn1AfXR/YBt8K0=
`protect END_PROTECTED
