`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2zY3NLGStiFDPBbUMKEGshDqgNwvT2BFOH6ZHDkhNy3LLcwObNptjOK6Pv4g1sPN
HnTnxVwRiFqyvv72mStq18PSc6jLyELYL999SgDIAxAZjInlpzlqlhWR2IJMabi4
hk4baQcExBMmIrSs1tK+6nM8LoeGS5CZ+T2c/lF1xtPsLqETs+IxVpvDjjzQ3jHK
+DnRuySNbSOBYLzs+lQt6uMhhfCO0uJnMnhPtvUL2rHKj419ACxHijgJjoGoxNnl
b30G0CP+GechoG7iCADFwA==
`protect END_PROTECTED
