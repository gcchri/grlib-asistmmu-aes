`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hXnbBWp2+W7prumrNqSGkhzMXSCqj12O7TSUMw9Ftvqgd0pN0OX7IoveXYMvHC/I
MuoC29H3fgj6zpmbBC6JhEK+x2KeZggOgHa/v5I7n01J4Lzd50uT7Chqq9x9AJM3
3QBf25LeWhJ1rVay0JZclHsO0mvnA9MS4JU5ctfq12xPWjxV6+pc+faTDGIj3DUF
kKXoq6E+2Whvp5vYpu1mK3JLcyZHYmBsoUkKjAwKPjCoBiEBRt1fMaElVsqIidRt
WVms7l6tzP4SgF+aJmN4C8P1Xj8UVVDOqu5bvn/JItvGnnlKh0uXsiS11Ulwdawz
amOYcI6BwqAqQeHfhup8Fq2WwyyaNWnPNuoap5/RZILW5LwBBFulUWjLbM10ORB+
v87cwyJKYSHRBxM9xbrxDWfD9fmEVyTVFuxlMYPhbCA=
`protect END_PROTECTED
