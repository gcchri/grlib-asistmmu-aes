`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0HLv7c56YOCtSXkRXdz9CjScQjygl86nztJlRAEaEQTjW+L6o+dEUCdO3UoNgJQy
xs15j7pqwtj5npJHIzv7BajfHdfS0s9HF73zbwM6dqmigQmLwm23MTN4Aw3UdDbg
bN5inAsGxZnmldY4IuxnaCj0kxsd4rfq2jg8CaffUAYLENgQBozKLEE5+3ft+4Sd
n/SI9YYMtNW6a+MrCYBYQKbAwy5tbbDuFBcPw0ABwL1/j28vW5+99X6MhO4CAZjv
3gMQhlT/qfQYfG8SVDyylugZTYBgbdXiKtcdxBc9reXQnz+MmB2hnKwP3dDXa2yK
8Ap5kIO7rksa0mGgmhk8hzd86Gcr4FOW4l/0UA+s7fiiu1Ef3gNVDmuDks2oLnJP
sln9236CELk1SFTRz9lAspCfxu1ZfGw+HWl4jbc2p/00xBHRzMM6Nrcd788E3AQ9
NZlAd/dk5Sr4rAWXLkdRkXBAohrjOeq3jUtQYb2w8VSl92e23at1PG+CblHrFTr5
IZaToy4dP3bpVUPk2fZlHw==
`protect END_PROTECTED
