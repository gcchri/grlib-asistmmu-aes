`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pDXf1Vcx5z8VvPQEdqgb3PnjNrE+0MR7b3HNbzdQB4KmklgwYKFpffPU7bziWpVE
UGbvOXdUdgKFsg+nbvPTnJXU5mLCbFt3DF/ASoCC7Wcl1+XDa8g7FkkyQ2jk8Z14
e54+a+gZWESmISUH+x0WIt8cs25WdQJniC4z5JoMQeIk0If5ME7x7IE0Pg7Rioxr
5XDZYHoJNq2/MhIBEwHZC5D6dOjP5JqwoR1M4b1UTQ8pJSh3BrSLpMCqSD5yg52+
Ozy1rmLx7iQnDfVK+G4EfSEhqKdnaYqCUDtub4OLExwOmwKfL52hluaSflByHo6B
CN87pwieXxFRzaIYxFe61ILla674q64XMq7ItQzpXEUxH+OwSXOMY5KwEFriHU8X
M1leZGl2ZMSoj0iwIZbSQjZBQ3NUQXW6CToiqmHoKKEwO7MqmbVRciFGK21UQz+4
5ExmSj+oMJakJY2+Hsheem8RnlDDaDisRcpf68KLzYPtiSCJbcwioL2YVQ2qCENN
Grkjkht6TvveEC/y5H3xPjO7b2plEnpoyBwEC+D1nwdM+TkmlqRXqv0jFoYkgk88
RHjjlQ42GOQUVkuhyrdFi0lLS7CiF/ay+I4qD2y4VfOrNuB1TpbbuymzAOdYOcVQ
tn1H7i8NU3TOncCiXqFit6FqOxP5YBIg5eNH5eEMElf9hneYPdNSn6504HDC2gac
lOeEOj6hTqipdU1ZzhnqqQuW2VXSpZkIsa4eqaD3cvZoG1arLLgkBVPq9aztuGUh
tittdlJ21fdAOGZMTD2LTOXtMc4L0EGovID0oqh1wTVlbdzsNCEvqSbHMcJB4C0T
b3MLgpDyQGDG+/gyUtcL9Ip9KzX2bzYm+kJVRpJOSRUWznnj7caZTBY65Ka8wCZp
eiKbAGOWgO2rjdpL5RwywLUNYMQjunYgZQxJBHfExTKDzj7ZfUn7Y6OW8yP1xluI
YBMofUXmh5MXIaQP8cP3CjlFo+oZ8c010Ov1kY7P8ZYSKE+oSo24vR6p6HNtCrp2
qndyZsEx6FCyTzG2Xz/MbfHe4odB2xUtCCdtXSAgopIt40i3qJkXbO1Os9qaUuyG
B6rgfBiiltHRwoYhHmpWyKgrypENH1VyDUHDQRUZ/TjDCxCIwbZrRdnAXNpvyFeL
6styexDby2iFXdpeXxYO90oYty9y5KUVMrzFxXIZJObbFUSHXj2fMYx18PUxNn4R
65kyifr213gUHJ3jcg0BsLXZ96D7ElQAVuZIw66hTZmYt4xMTlstk4eOLWaKYNSQ
f3uL6IFSvV7sAGVZqKG6z1PvgiKVfDE/iiT8flc1I3kOK3Qn/XHruSPVgoDOmKYM
85a6AzXw7lkQ7XDoaiLJlJ5zf41GVBYyWwI86y+/48NltzsngF/kZ0PN0nQoJVOz
`protect END_PROTECTED
