`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rhr9/EGggMB0dtgd2uwZ9SBXl4S4O13YFuza/sAgFap2wK4Pflvm/RCgh9cseLcA
k9AmbfPjg8FTtdHb03Es4xTa/5Fta5GEgE/1MwASjthpl/2XD3H89+Kv282wVQvk
97bqUpJLnxg1IHLyKHWGzwirBa1skfpfs7AFZRsNpgXk5x3a1VdkKoocsqvCy16v
oLOcGpGeT30hUGLyST+1z1SLDXG7Wb9epQzW6MDaNiomPS2BkywgY9jLX3StDd9b
md5oux56rBTnL9PnVV5kARtja3Hb4GmZOPDla93HppPm2VmR21rzzVMTKwtrJFcZ
7mStD3dj6tDxoX141vAiXRUyQ+LhpBYwZ+9vrHZUHR6mxFWfWVG0llx6l0+5S99b
KTv25R59O7TBMm796iC4C5GB+8Pb1nDbvMKHKqRCO68V/BLIrPpm4I27EC3l7nDL
TlnuFAC3R0i19mSnnqsi+lXwDR008R6ZbOFEGgwiPs+cf30b8HQRLUeqe6TEYO1L
ZcPD7aD0dpPlt+tGTkJMLPArVSoXp97I6S32COgD6tMaE0ZSOkybsnkOLeDz0F82
dUGsWxh5/cRDpZPKPYJmGaVzXchaLttS+zPFOB6g8orZ4cP31cMa18ZuTgzZPNND
vtP74w5Me+o/TGswAAlm9l5OKzPJVb6nNXw0bIS0F2wGpX1abR58owgM5ydVeYNm
XRfxFMT36j+FRV4LgCFQL5xDN6RgCX+UgLE/BQiOOnaBiai6FnbTWgkoRPfSdz/1
S2+wMi/y290JrwvKdaGmcQixNFMI9gF21Xr0QLUrB4bLWvS7RjGesLK5AC9N586D
CIfz/JKJdWvjNCBnJiJYuv7uOY91n9MPGwWZuLRJ4tsaFwb808Os0rstiFIgnMjF
M+6ISFKEPZ4Cht4Q3CXbJD+MlP5g4uUzfprI1LDSzpg=
`protect END_PROTECTED
