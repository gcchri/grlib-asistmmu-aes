`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bvUG7Sa3HYMmQIXhqnU4syBEX4ImiYVvGWvOrlMmYjeXjGYWdeqL/4x4eDxh4a0T
CfGK7DA+8lrrPfNtT0XjPoiACteQoGIYtvKT7oixPX4++y1L0QGuhXGjA/BELN3C
ZcdizYmwOiZjXB7oz/oF7B1AnhMqXnL07olxr5TRYqNitabFwqu09u67nQNYcVyp
d214qcpN89nRtupSeg8PY2v4Bd1F5nQL4HExu8UTm1h1PBs66ZxkRp+pBjh9rnoI
TfXEo8xrQB4SbY6NBBZkkTJAN5NBInahUK7Ovj0lGEJFSKFrIvQzvkb3C0EoJL3x
pU5AcmYg7fLKzxOavgXc3Q==
`protect END_PROTECTED
