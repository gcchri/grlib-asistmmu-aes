`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WWa5yug3Dlz79CncJRJSUitG+forGRBXVwL4exdenyvYmj0ar92I3vPqyup0y1eK
THK7++NyQx/xMBGpoerFFTFhSDTRM/bTFOc5TBBtCAUreUjVudm9FuIuyMSvkKol
hpZ9WMSN8e509Yw3AmafNfjs/BuvwxQsdiitcn7TgdphcWqf2Y/BQOgHrjxUrCnu
Jeb/nALvdQvy2aY0ldvcxi6iYziDQM7hQM8CFCB/wZLaZwbqcDwVuCM6aQOQXMpU
5blSOvTtSQmKp8BSB4rNZVdK56eEVBzQ/5OMt79j731F4HWu00/f2ZvbcLEavLXq
O/yzFFJrYUIpWaKkvaC4kZ/S1wWoAw6u6/aAi5cng5dbksWTjx5yCKBbyVhEmBu8
Z2M8n5qmF5+C2U6JpURTnDBAA01SdqnRO+Rxx6u2Scbjj/z/pPbnG1pIrc6Roxq2
UPEaAmrc3GjxNPb5ZTWzpxzdK/ioWP/GpdADscxkkh8h9wHoaY0THI/3RhV4++rj
xOQe1O34VfY7hZkYE7dqXiNHOlS/2YeGdFyFGIizXCwHbqGif8dSASYLCs6EPZWe
ErYyA+A54AbnayQ8BZywu4r6NVbYX1Zxmw1IcbVxWYyXAy+80BDbM0zZsJMrdu2L
Al4M9cZVgbItnDuE9U6DM+xx8cXL1ukhGh1ytfPPfibfJ1waT2vghnd2LCkVzOLs
LqpMkCRyZmizU1aEkvuTX9M/QIrItO2l+kgpjBZO5Mvw8eIDNSb3sBe8ZwisyN6l
0qK7MaMRfi8Pj/4xRCh3eUA/GjRYCn8bNzTQZAhcUsdXLiIG22UD5x9JxSY09vKl
i4HLspPIb5rR0NnnM4O+F9OO71Dmeag6Yzx3oMUwjkR2caVSVQqqbEWLMbNSkYBa
4K5SI9Agmdo99saG12GE2DbLx1feaZXme4jMIZ6UH37pFtoOJAVIAjf7ghbwQFF8
X1yPJ2YHsdaTTd6c+eDtuRLy1jIyAZhI/Sj1NGkurO4RDA/POFFfc61to1Ipnheh
lS8Umm6UTosLyh9nQYT5MHYd09ojkPAkhU8MiVMi0s7U7/6oMTZgFV75SG8gSQ2T
KN+FivNkElE6q/6fUaQaTpmGnX5lYkyhoNQWW6Bk6d8nlzgO2fbQsRcKbwvkAUBE
5Lzhd0YG1RdEe0ZpG6s0FHRSM7dT/AcJbio+kpM8S3QPv01GY/fJNbTVbFOub7er
gAcvH4DTyExv3ofsJL+u07v5GwtXWNCWZyi1O6sd3moQ9sw3Aa7sWU73JeaUDmQu
SlWZ/Mjz3JkwLAI71SFKHBALOEksEf0Pu3BqYi9uz3HFJ2+tH3GYgI3aiyIClaPW
TpmxxEdLmh7kPV0B3UnNsktD0Gt0tGi2QzF9vg5pVBepE5j6I0UWnTzHNBdBarXi
6lirS6eypFEH9+7rKJz2omhOZBlkr9pmmH/PrUsMGTd2QvsgKVGusgZRo1gGp4OF
YvmCZdRfbYSL0YIpGi1eQj0dkWQ0ZXsdqatR3J6xgJv3uRHH2nsK7vOhg7NTJom2
LlIsRZ4NgSwEnel2Owua+sFkrmDgtat8/pndEr1cjYxTKx28sI0FnX8sl5/P6DAp
53z7RPQzMkFjIqu172UVdvvhQaUVIF9uY0W+/HEt5AvvzEwh77fVcrL4WK3X573l
7Sew5/+iSec3gymfJG88kq4FPW2TzXlSbKNlRoGMJUodoxlR3J324vbmZViNiYro
Q2+ZfRRZTjgQbXkNQJAhDy2fF4/8qqqVlDKyhcNxZWU7FKunhl4nxbMWkHuRd7Ix
mj/42AM09/TE9fjyiPKRvQogQKMeWawkVhy2xOe6cluNxH471U+rtmrfhfLf28+N
bRe2Nm99zayioGshEIsK+9TyUhvqpBatHq3NP2PzjwpId2X5XoQ4p2Pxy0Tjw9yi
GYYKJOBM8KZaWdYnjk1L1xG+hZOMtUKqWLuFYWTTlwi/5HRL+KdbAxlBAPW5nK/y
josYZP584Sg6KFrJgrxjs07Wuggwb8BGdSIOSnd92VKE4XyEy7RPoe8sj5uNDYDN
owJcAnh14Z+p4K/huz8XVbNd5U/Z228Sw8+pyQfkFBeSKM5Ecjwk7wYs1t2ya6LB
1Ypba7IvluS3eLHr6ZfVkWAyC9Eu7GJzjUeCwIhBMPQTXC2b1syzk85KyU6WpYe6
DVebrJthieQ0vNAXhZBPK7MovDyXaUfKjewZfxvUCHUxHT0wBaqKzI9oIqflsccL
/tPif/MtsCigm+/OCwQMf2JTG/T81Ycu57Lv/Snnk1Pi4+2ROOjcnY+pkCTw7X5q
utnDzRQ2sd8Dxwt28VfgfQNizTouxwvHerATwAWHjqDi5kN38ydhp2n2oNjHYMmr
yvihkVG8NFJS4947xKhsci7hI3WH3zV7GvVmaSxd8n6Ice2oDsVaBDNa/0d/0pAh
GGPoY5N/OH95GvfQ43gnK8I+2bISlQaKeISjOywvE15NcSLRNBt2IHP1ZmaLV1ZH
1zIFG6cpnm4/W663LlPUWZ1dSYfzdm61cUO72MS4PoRdIoBtN3tZjOPojXbtuill
mAam+t5Pp3mQrgVmjz7lJbGZjv3yCljtWS2WPS87V0yUOXxfxtp6XV6kTD0z+lnJ
abk9zvP0uDeamY0fszpoRlvyd+2FqWLVUEXpLDDv+yEGbrT8PFd8bpZykKvn3w5U
5r5LkKOXirav81sual3H2bZ7vCxeMejaPA3vf+x/W/fHV9EuyUrEqkliGiC97YCc
6vSfpReGnhhWQvBXyYp5GS2mi+kZEgD0nj0+f7Z/3x13X9YDs4SX29pHyCKCECyf
65zwasYOCY6BxYyFlvLAPyN70FP3qk5l4rYKGdqIUJ3SCebjJfiezQpB4tm7j7HX
woQTjcfi77AoNLihi64GRkLSiXUScidj2ZPktPIzXNGhOwV/ecAY+kXNz0NCOBac
5dg/JDb+djK1tBwPRD+QL9Q8Y7zICl8Y17yf9sIlCd72DfKmLr7cJ/U3Lg/I/3ct
1oBnrQtWzS6JGLjtt0pjYdNVRfnTmQ40bEYcddbudnwMQ3e7DttD/8Ev8iAPGWoc
mmvU0aDff20eYdZP6BHe/Qi7brC7hw5set13/SIgMlfPnwfYM0VtQtjuGAZqCf10
pvB8bxJFx64SYP8qT39qMYRavLGnygu22Nn/W5z77Eet1ZMUZn3uoQl+xQvm6EaZ
hJvhgT+crZB2YoD4kFzkDgWKmjBXwtIFeNld8Vzgc+WSfkYizVZcVCt8EeDV+4s+
442lANaIZ6qENULlBczl3QQ4w3HrzI8tJ2w4oGxUVzhHv6DsNXyePYscrkXUk+Bt
+VPrUiD8PaIw5YRqmA1Fw2HJai7uHbwu72vZha/VuFn3GW2omwGlHIJnQjFkm3AF
FpGRlqnA31L2ZrDZqtr75f/dPcYJgVMpe7v2LSKt8WR54ZWLZDkoZog9Z+39Mp2G
AYtYFLN8nDHA/0bAq2yrMyxnKXm+BpVFb5DvPAC0VH164IDI6WZSB+fUuglI9jp8
TnzexaCk9K1ifSop+r2K6Q==
`protect END_PROTECTED
