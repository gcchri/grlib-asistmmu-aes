`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tJn69iVMQrz7k833CiPvvvlv04NnZ57kUCweWvvldJFW0yWctMBAzN1zNPjOVie8
JLtAbDF29ivlY/PXmU8DllADUqTCigkdNg7jUCLRpFblplPQpACHC29MfyOJsGWB
mFKGc0zDydEwvoRpEd/Ew/qALC4sCLsFS8HKVK+uh3RIKLMYDAOnf9vWruymAjyq
P9wUyczOEYMSDpx3Yzg/P4u4opnlwwynSUGO+ZujabrjZZ42oQJGM7xA2uIqt25W
Sb5HN+85Et1VLmMSPWokfaVw00KotA/wPPdvNlGrdUcgon1qSwlgpBFi0d+FlKqo
PCaStDe9GyMD/PRoLvbcxQIlbk6dg4OXqQmDdo1GFBPI9JdU3wryCoKvwekdMsAU
AcPKsME3Q6LIfNG6Vu1pwzcVFtjDuCs/o4hNwkMnv3Z7/RRzuEQDAbekcb4zDKGo
V03h+asFUhLvTe/ra5r3Gzz6PViNBDwMuPbiG4FePqBo0w+yiOsyNByqPcNo1dPd
qVMzJz9f12BiM94t9MK9IA==
`protect END_PROTECTED
