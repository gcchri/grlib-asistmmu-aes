`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R0k5C8xon0YkLxVHaYdl9ZGxF3kV/kflkF0UbHy6aUmo9TdAO9XaUk3AIO4MGY68
f1UEnlkLzFYUkEewFS0ar8CGm3+B65u4GydSkNvVjbXiUlwg4T3BYZtQxGPyScDP
LbOSPtf6brGluZpkZT1NU81gdLORV6UCHLtabk2M4YfqJ5w8tQjx7fNbIn5Ihee/
+SLQLJRl3xfx6zILa2KMjBf4ZqZdoLfvp+WRUUyshkhfsSqeYo5YiWXcozmDfPYK
g9su5PVNsvs5WV2yG1pN//Obt1l5IVSazVEiLe42gp5VKfDmzi6fbYH3Ii7yOto7
IufoIh8ZLIN03lSclzXbUNABhuQX0GszD0v0sUxzqqBQIMC/eNr368D05iPr7ysE
RY8o6svJNEx+IKEGxvWwDf5oHxPkbgjx4cuq2+qvPFE=
`protect END_PROTECTED
