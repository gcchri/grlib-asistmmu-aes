`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K+QZB/3CPVo0fNgY6iuqIywGvxgoW1fqAjEegGY+4UqSHVkEKwMLtk4cYPuYzU3K
IekTLVjh0yne90NPtvQgVWDEXRFD5irsV469TuTKw9Igc3p+EllI0Vz+4cXvZH0l
X5hktM0NexhWBEO4f9+A5+SdYbxOZ4TvQ4V5jv55FrF5Hzjcc/cUhrWcwn5BWMOW
VCYjp+SAvEUrhgpqFzsQL3bU/TAlFU2h3QUmFhxNbF/PpBOoq0X3ZMcy/cnPbxQP
3iGLjjn3ftJpb+s5cqGl59P/U9GEuufT0eeWS+pYVYcUxF3ajbVDKYMJ87I9miQw
yQhhWDFOmHZf8gaA3+KVf0zJRpiAQbUBcPNptvjwCBimlkf7j2zwix6fNn95X0Nk
CuMeM9BM8ZxmuH+8X38aL9Lrrl8eiy0D5bxIW0llX0EeI5/+qfKsnyiVl5yZ/3C4
UULnjKHkSl7U3qOUJ6Dt23vygyTMEqzUONH2QoTDp+YH87fO8SQ52xBqEninKhrp
C3exxai5nK1Hy8daL03Odot6YZ82xhb6ofYL5LgnoIYv9YK1IrMnuPgEK1qPqojN
OInRtp+mrchlJsHeMrm0Sq4YLRqipNkz/8uUbqZb7QC/7N4x/J4clePnss84Sqej
UKrczqRbiTi+oCA4qAwnJg==
`protect END_PROTECTED
