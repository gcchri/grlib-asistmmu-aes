`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O+MiuSnzA1OGQRxsKZyZElVjHYvwq2Y+g1fttkRij7QN1YKgVKjxyu2Mj1EloD8z
ce/EQqpE28U6AYUNBhW88B6WDZ5NpJnwDzCIbF+SyKoHEKLKLs5o28KnPN3RljH5
KJkCwx+YV0k8QdG5NCi2G0V8u0NygenGIj70S+3i0fQFmQ/HOAFjn7jqOxPjBvlF
9hz6Xs9V3C8WxbL0udLzYqADaxMJmybmTuciAPIX7Z4RBvcqg7fKkuQ8vZgU34xF
wnUyazU8GxsvOOmSFDn7quH5eiwfFDjYKnz7AqS3gs4TtD2fGRLQ0EMjAJRPisyf
QTuow+fOFVTno1RpfrpoSBfTRr9KtRk9NBglc5eWpMBeoqUmhTHZWRzOV/p7Vju4
nZC2xwxukZTDlDWPfaz+FJnftloWfoZXO4HOGXjeWrs84ZW75+Vzkw0C12Nf3Cyj
WZ6Bc612mDX9R7v9zT9SylxK/YTKVJtkLtUI574ISjbGjxpIt99TwcudxGEfe1k0
2dItbdg6JOtmu8Uko+HHoZqnLOkkFVsHq5hVbavca4saohfreWUsK0+sVN5rcaPI
TCLa9AYTciL+R8TjpuGj+TSmyrMd2jPDva1tISbO3sqLs6dlxJGZIT+xJkPiy7Gl
ihihEw/1fIklvtn2XY+1jEuR43GP2zyYCy4ripaDAP4RYivBr2UBNEYd2b+vyAoE
XZ+/P8Zs4p8r0R+CFEVWhuW2A3uoezmviq9uz8QrXIH9CnUjukwk/EqYYXAFGbkk
cLmlPSFVPs+Ol1meguYOhr59pz/zuXoEJTkwId3r2hD2PJ+uKB57vcGorCQr7Vh6
HjVqzNYdSOrbSKF9P0e0wG8GQL+gPtBfN53lQPBOyBENG/gvvdERMA6Ymrujx+5R
+wR7gsq+9OOXstfGxceGsiutPCZHXPm3pyry/F8GyTKkiJWZQVIuxx902WFg6vu0
eFiaklDa1e0U0VpZvX3O3+1mAuIr4FFCoJK3CeDHvik2tFu0skm8LEOGhVra7ozX
bhI2onJHBhN+2dm4CutDGIZPmQBtKwKDCN8kvhYqNLgzmb14pdI33ZCTSpLinMCA
trieaJbvRf3Fjx1pwBW2iWC1VMwjNwlTvchuODTC9BLzKnwEBibl/Pr8nEN+VpTE
/HpohqOzkNvcNUpA3PBz4EOqVG5CSHomnrs9yiugBRJXKb8HfpolvnBPLt+ENcAs
suqJugCPAGXBGgpKMNjdeR2As9vCSBmheBUegy/DE8zsrBuZVgrfpWMk8a59nSB8
GAulTKtJtKw68nWZwB/S24WXTq2saniAAnslmLPoLshFMtX5/dMWal76bMQrPJGs
VdmvmMzsBj4SFb/hOpThbPNFdQvgj+u1YFkBLOFDq53tkIUp7TyC9Mj7Nt8BHWha
YbMcgXE4S6ziIpbDlTKobxqC0IqBqVJnAciyfImvrMwTzbs+ZOTV2c5kwp+RnYgZ
DkdDK0C8/N7ZkZQPTtj54TpN8VyPb1PuzVQd4AtRMd4BZYfsNOlU72hX975ppCs4
IyNt4G6KoEDn2TP5eto4pXrofXZXFXZ34jnFaV0mvhSthmSDoo/AbnGe8nuurTNy
ntF00Z5weqEy1E5ptJSLp17OWyy2e4HQWCKpTwseIiE2oBuLZukaWhzeSHZQIvt3
80OXEoIRA9KCxw/s+NnN3tqR9BiontmMa+7jHAukGUkapCvgzFeBOXx8rs5LLUse
2HIjZVgpL63ecoKmTNzJJ/pJAqmBbeWq/H+yBJN8bSOrlO2bnZ3OOmNGxcpbEohj
vEbT1mfaJouGmpmP3Yinjtr61A1BYQik/MzeWYPXVlLhkN/lZFZYoJ+1/b6iSavN
imed8mu8sMhjV6eQxHrreMcz6pbQnSue+Wjpo8HgJGnM9OR/t4xlO1gtAoT5ZP7M
ASeA8UcqcFoAKRDfnrbMfZdIk2imXt3lPsria/vuakbKvA5dTtR/h7lMaLIApHKi
+J2CMf4xFjmQxLu4VQB3Bb52o9JtQtUStCv9CDmbTWLnD+OocsVZ0Ywp2QwevEEn
IbFzaAUFRqVO4AzgpNCZ0u8yU+VrJVRg3YAVUZrevBILX0koChXa0YiWBafGnhqH
ameKVsme+3NEUHB84rBnbbSWgSY5eatMh0TKwCurvICKGokLE8ScEGwWm75fH+/w
RkMpc33LdpYMoM0JRj9gyJlXu6mxZtkzbvUDb6qwSsS8jjDAk5O9Nm/DrfWWqqYL
G/21Nh7YWiYvkeIRT+Ot72uZ567EqZdD20c6oRF3Imj3nBAQBTGqU6sdXPnKT+m1
s8FlriHOv8A8lDqMymRBqkggjVSZmUKEa3UsoNrCG8c4ZBrTULZgfMVjaksvZwnv
omMBpbeAoLxuUT0U3+pRwFaJ6MvZXg9h0y4QK/ClA2rsEegQ5DbEZoX4TJbjUEjX
JW8BE1At8swz4KLoCQXp4+k4LyOHiPux65u3VgmUHML9UaUpA3wuGciFidjnKzWX
tFLuiXAGEDfAzD7p3CndWbINA9O69n6mSV4fYrFERm3pLVqLbSBrg8+9GuweQ22z
5VGiM/pOI84BkcsiKxbBO9rVSD0NcTjQUKUMVrM9iXtSWO84tQuQQbe/cRlDp9Pl
GzsokANvqcxIH1l0tfoeHEvRYLh9boWXlDh4xgJLiyhb0YCgeHmI9OOhM9Hcnkop
0Q1l0POfv9qooSX4ueYCa9/akcc4yGYtXW5WN8S2kxMlpRLiJD/dEVFBHkOPdfHr
EnPXYA/jOyKCFdsW0EVu5wU9iF/GFb3LkXXgRU2fQJv6WyttZAM7dIGbZMZBrMSp
HuW0CfRFH37wIyax0xunVR6WTXQZyqpC2Bb87YtxdE6H+Cwb5hkCti0dtZ+0OsSo
Uualcgbmcg3ENHwRXHS4dAlaZZZKP01WkS0Gil4zZmFxUfIcAgVGo/THuMun4nlB
NlAi9UL02Gseg5xvvUHgWowLAW6J+8qqVsrz/S0ZwoGv4GMfqVZZOMJTwv3R4l2O
FJaoBIXqBqkylmHRYqsNbI/Jbzss5AwjURPB72oIYy8x7JIi5ZhPaTwbRhn1Qxcn
RYT21B4DIum/+kv8qIhaePS+7DdTSTlVvUUikMOPj5O0wMcx3v4abb2HU3xqzmZj
54ja1kQJnlVH0kXfq06rs1ZMpecMSVhXielzddV+4/GAz2ZYUfrSE5aPvaL7G5QQ
7frJulvJy5VDATRurI8y+0O0yr/lSqqfXHebaJmRBiTaIWcJoy1qZ7ZATu+19C+O
2Y44jL27EAACnsJNcJ6We6PDW6zucGIf794pv1mmXi2JnojqPeRuKC4b0JIbsX5V
lDvUpUNI78I2uWpo7eV9z0ZEZ5/hYiPZUoB8+UgPDi+K3YZMf2fK4+C8gBxxD0Ly
UHBVB/8EDldNducNoxT6iKd8eDmLRFEboDfFtc+rRCFhkUyAbPgt3jtQ+A8rGsNT
sP1pMzWmt7Pa3EBeR8tLKZtbB3R8oSPNxy68YONWX97djU9fpVV09+owJttq1gdU
Q8UxDVCjKJpQ1R0w29syHmcTE8FJRCUURS2EGTkShka62MN6o3jlO2KK3N6mL5ab
Qcsrg+G9QSM3kVBUBKf3NLfB2b7miPp6KfJ8DuDA687noBnPqxD1zF2lt+6p0WzO
zMd3fAxlWoYI+BE5vFQKlMfC42QfiG+GGGUKCD1hNoJA6nU3lVAvQ4ZoAhQuFbF1
2jCgpdn2SVamjOv9+S9hjtS6MIpmOfbcc/HYUYxhA77Lnmxibq7PBhr02p4BmCA1
X5ra9w2Ql5VhNGzjdqjnr4sO/xMdKX4JcY2ynnT/kGlfzDXZuAf3VUpIu7REfqL3
sL957wxLmtGWUFCV8bGUN8tpOP06Dd22e1GUwo1td0nqRxOXSnlCerbqyxjqCsMj
rjsnkHFEOZhM2FHjcqaMp0oycMJUd4YaPHrfw8g51rpB5lGkh8h3WHhddEoEA5Vh
PgTpKFGDBjJLUS0tHm7KEm4Bzqw783t/g96yni+zdijV38U3rA63Wbwv47tgkoA/
9hOHt+vYEZj8+opw7pUj0gJ+OliCjGWWZfjz9TClvCYp/P2NwWSOtGyDK4mRvCpl
T8MaNSJXa/imNDtk81UnG0zHw809G1r5B4/cG5JqYco7KwFoH7ss9DNxJckYB1vK
jXz46CIwBdp0kYm686dloPzTciwy9si+QkfcO7cEU12jON7WFJzItFVgEFtN5mz5
Kk+ZY8WLVdk8fA0c+3IEPQmLcE7AW1b7uIgRbefJCmcIWMTcbNfOkX5q0tmCwjUU
jzP89fAfqiqMsIliyNzKEXn5Liv+D+mBXiSEzmn7nF4lPFZQCMFxyr2SNbJiqhs+
PbWjxrkfuDUKzaYR8WJjXy0cjHIuWNPxD3nsoKVMdOR2zqANNR0RAo4aRufOGZw6
twc3PsFowSv0z43bPKiEQ/nPJea2aQB7bs9RYjBBXOs1kBuFZtNn04NAzGE0RT4E
vLLEzjgQTsrQ7ZpnlnYXXDuZeimljNfge8KOkqm3eyauiuD98cFkh86b9olHRpB7
/FhXzKIjxAn6U5ocWMo0gnwiJAyZargC+2z+WjLWvm4kjaIXUEbNBNB4nwiJDoDB
kxmUa5fphQLN8cvzlJjnUOCfK7121/H2olpatu9Ij3BPNyI8Qbp483xY1Dlk+RIA
us08f5RTZeZmq5ALEFR45RiNydJVFlQgCRbyUTx8NBDr+Ku2PoCqgv7Om9kkifJg
KOwdPQTfqiGXWm0Oh8UB6TF/OAVGrVzRazyAceUTyF3epvzzRv0igZj/7JYFv5Ng
osY5GgaOseymGE4rXV4+YiyQTH9fo88W8z5uKEtNGaOYfmekA0srCOOlbtKJH9QC
US3R61AA5S0KVRpOlV2Nu1nOZr92dlolG8Q/dF4skD3/xNTk/5Fr+0MrgrwDWs5V
ISjH6YvldrC+/moOE0xu+dYaImM2DQHeDKOVR8TQe2XRC6bzxKzETSHWFMZOGxFG
6DoAERuJG1OjaZAhpmDPDtVlhzVEggmxq9FBcFRYtRli/nrqZ+VrID1JJtQyS28Y
jHhS4+mKib1Olg7e5l9Xjw==
`protect END_PROTECTED
