`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tPuaAbY/z6xcrKY015U3s/tAXoc6CXjNH7fIQh4sGl0oprh66hNeu0PuuAcfs9dJ
GB+/gOjYxDVnlIwpYxHAcaQWWQqKHcwd3TyNnutZrutmvZlRd/CdWVrH1dojuiJ3
lJuk4i9XXLbltrOHF29Av5YvVNRTOMQ3Y2FSUrKEeZN7KMyp6w2av+WKNyIriOWI
0YG8+RXjQkd376znAcRlkC+Uo9DJhZWogZkIXWDsO+a5dZ0QycGKHJ6bUBW6J+Nm
hiFfIFI4ibmyW1sSglri/rK/pnVTouBNQ8P0VX39m5AAeJM1lUmRbu2b0Tscz2mB
P6Tb04q7cf4R53C5T1T2VQb6hvdbbPIWpu0dVdFNpEhLF/y8g4ujF1BTaP6vujXK
6SDIRGV9g/4YHT6/wiw52eZlsGlnX6VfyqkcmPrCSp0RFs4M5krBZGhKAekDn2wR
vsMmnk3iUehgt8pBHLVNORXyJO7SQS9dh4DAPBeBpFGS97mf9E3TjhytMB+fKOM0
rjmWRFq+b5LrQADblx6T7IyVpUNYTnkWz55Gwr+5EteFK1rY1HR3bVfEuZbn1nvt
R3umAZ03rtaAKlo4eamEQg==
`protect END_PROTECTED
