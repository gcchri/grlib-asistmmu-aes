`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gT8HK3btHnprZtLzR9Lzh94SH0XWaAxLffjsy2tAgFwkOtVkJx5Y/3pApLuW35KE
F+LD1BcK+qsM4k/X2igilu2owbj7Ylo4Otkewzl2taI4SPtnhxVAV/HnUtt+dAUp
mlVMJ7NKWfovV4p2ZvEZrPGIKpS9ztRmkqK9c7xxmcoWa+v9oNPZrVZUD06keYW2
D0n3WSUXb5T/LtCS/ohc3jxzOIMZrYInuZylRnVtFj3qZibl9PgdCWOQsHi5af3o
w2IEImDxlQ1S4GqO7R5uH6oH2nZLMMSv4cYHQSUSGz9wYSogkblucDF59mgq8Uog
hfffEboQTBLp9DzdfOjhnmfq21z6GB5TZsXfGoI+qRk+Fspg/mhgbexnnvtXgFrm
BogLmggIEu2Pd2Fo2MXSZr0vqj2pOu86C4PaThTaUlscQ6KLVhHeSO2gn8twH81F
VRY+nJGkbRmuNFNuUoUaJ3NbTaJzdWIcpC1DlcYU5bxT0miYrIX6FLMtUq8p17wy
WVNj4z8pHi8Xs+u7DX53ENSWnPxQ7/7ElGsxKDKMFwtacfPZ/TchVfAiXc8g9gBQ
w2DB5YOFWC0zjVvUOh6MY6ulgMHfylylxd+OPlGEugjbGJiXk7xV+53nc/1qCp/p
AYmRu/fzxKjANrFeTjxHa4UoDxmQOXTDjlI7GzxlueNGDuKguc0ztZrGKd+vfbUR
IaDx4PGRMEleeV4j216UhU5AOzS7oY5gAvbJo/8J2wEOw+S3Ru3Ue9nUyv6lt6uR
T1xrWosZa03fTE5p312VIEaNd4dxiJYnFTyqkrTDZUOGRQzAhJfxTea6ycJ/V2T+
vvrc2hQ9uA5b4osICBy2EA==
`protect END_PROTECTED
