`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CsGLFQByVHHEBSwU0CSohRr0tgUDYL5XsYflms0DAaaFmLiU6jUsb+DhwpSTHPsw
NaxnqXeo7j2cjpdnIj9gYtzq3ep4CcUWP7gGpLBa6pDADj3N36OI5pJ297/yjf+q
Ld79hb9L3O4SqjVp5jFOZUWwxg8EnNJ0ERmXDiKyrlNmPKz/Qv5R9g2hMC37TZw7
+KvxGL+da2lqjJl7cmGgBeySd/U+oFb3giSA5iREIlHr3HdCe1Xi1f+ri870goa6
qHbaEND5/RzlYA/XZ877/5AnanAJL3bqCQVb8IjSplxYrlCVmQjnvI11ZyniN/60
fQVtIx9nGtce7wL0FPN6V3up5pVLAUPXTqeguqD2yTyCyHNbLyBW/W0Am4SiS81q
Xqsnsxwb+lUDyh+UW7v8JnGGo0Pb62H2f8v6M1TdSCrYvcROoJz8ybxgsOvJYkM6
`protect END_PROTECTED
