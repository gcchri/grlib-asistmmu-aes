`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pTdbtgoaKI9EGDEvAyiyGTiwHg9AvNbvHnSxQchVaro2PFcguGY6jCggHdDqAphD
t28RlHQ0kVOfD09R9H5sYUClZp4nEHp9V7usRhb14/MDOfK8zBv9qxrGyVVowvHv
jed8BSD8uV09yEgZVkepNw+/46TThvaA3+kkpDm68QgGl6ILkMVCMdye5R4YXTZH
zfQcFkJkeg/h/hRoiNEYPeAgFaOjzPGPe93wLzuZgO809x9jHKyjft3qDMEIIj88
ewTNt3ggSEswKLDZlTE2cw/KgvcXUMltQf3DnUntIOGMSgxl5dBFYsd/VLoyWg16
qRgh9uE21eZm7JiDgPS7JCcsrUK/uhbjDpZEe1AAa7SdObJQH2X965W3/NgFda1z
hrtBUWKwm5htnQgQo3TYxpKRyx+Q1Esbx3SRA6rd/N/0mU0X/9jB8gOKSQ4QZQP0
z14Q6jXMsnvwuzA0MM+qE93fv/JHRCmvC8oTOgxpd4Bc0OoiF+PoJeR5vDzjvs+N
8eTkLCt2GagVStwKqJXDASDPwkr3zXCCDv7RNuSGoMg=
`protect END_PROTECTED
