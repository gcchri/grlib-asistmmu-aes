`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZwN6WVJqLxMrCa75favqU8yqJR6XxzGyiQ+c4m837BiIWBdc2llUD5CrTRtDuCSq
Y7TDeUqu0636dOxtWgyU8zzZcBX+os4qMNdR9slEzEkKxyNQCIR1njIMeqI9XmuE
A9nDWn4UFxE4ebHoKOHbwv6vsPLxIVdy4fs61PSM3r7Wq1wU5tllMg6Ttp3/47oO
RT3aiAtN4HB4VXYCUpk/oXqKgT3koMlSan5Y/540I2K89Nin9HfjSVmp6S7j/tHM
gcE9VVtwHa9wqKNJLmaK8gi6qHxU/ZL1k3Upwmgg5spS5Dnf+AyqWFxm3cSn5O64
6s+NTEzghtuOreaqtW0foFDQlIqCwOAkEzukweHiHhpr1aoKsMOcn2kspTWxvb8T
53S+LQjuWM4dqUJTg81bVSiQJ6siQxnPaDHY4MTc3nkinQmEk0LWo2+sWXhRg3CX
C0Ug0LgdipNMiclA53cRc1GWtA3cH6qgmtoKiy2qsdD9n2qUqE40rP6v5uLYQ1eH
VwkpbyE5h8l9fiamBKQyUo4TRV2ViI3eyTZny45v7z5Zxfl39+gfsLdAQQ2Aw4JE
U4VmbiHAsgqrEOUq2NwnLfWxDYdzNXOnjsbqE10BGaLLBxa5FhmCLWOZXcy6enSi
++u0Wvp66GchqLVotj8kNrAaf9DbEEc8EeDbfND2RyH/d/KXOZOV3onlJKcf0/M6
N6Rwd4oz5NMKq7Y1mgTH50ibz3/hTP/6HifgX8umsnSOOzeZ1OWI/O3EbtXlCMW8
4oiakIpNKlQpitcq+AXvNqOcDh3PTG4Bg4+twQNALStC9aPYJRi7MKuvrsLLWJdp
EOtpDeGSGLay0mzhD2c9mYOv3f5gKQ0IWwmrgLyL6eT33gY+8QucayOoN36TnfX1
YjY/AvpJgyKRiIXSbZgTgXX4uEqKGggVUv+ZY803c96UhjmcvlxbllOJhH1PTqYZ
`protect END_PROTECTED
