`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tGo3NdCt1GoNoaacTsm5x1JEwUCEjb7BtenpQN4cBM5aY9cYLHrGxRaoGewnLXWO
oE8U4wELKSKiQSFut5+OiezlhwVQqOp1zXC2xqId/yWIza54pcVSlvTbvcPh6fIj
qxKjv9q2Z93P31HJPeuu90i1Jpe6M1MLnQViKLgCLJuCTeJhOJrD7zsWxQF0It2+
mYOr92DwwKjyYXt3+SSnpsdh2EpGLe/2sKZGVeN3SZWHhSdutM4f5gQjiCV3u2E4
nqt+U+GrQaN3vWvBkDTpvo/5loREAl/Yi2pQY7nd1w12pybLrwzQ6ZFb3TBYA8Tv
eB9kvgLOxgJwIDwwPRKWUlNE+TQjFhJUNHivRRD8clA+uhmEtVd4F2MwJNBKir1W
HCvLAnf87i0RsNF8Yw+qdz72Rp1KFi230E/3hdguEzEh/0s523Slt2VXJHDs2Dud
oMWVNRADgBaX03drXUmg/OzynfbFI2+W6KiLM+OJudI=
`protect END_PROTECTED
