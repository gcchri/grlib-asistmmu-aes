`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A58dg16raBUzzROcJApqzKmPQPrqii5pc1imFHJy9mbx0nssghRXtVQk53o5GfJe
mOlY6EGI2xd76yRZOW3tH7lPTa0hi9Pl2JZfnYRmkhXS5X4gu3ZcuOIYYOh7XN26
MD+nBfkXUZ4ZJn98sbxKzu3tOPjcdcTmkaiMihEjZeZeR0DiIsbzeN2BiiJmKNqa
Paon9zdFVMfG5J4bnja3Vty+Oo2VPoq8Ut4bLzh+7Y8xYF0e1+M3tfheB7DIquOm
tbVdOFZWPUXkR85hSRm0LkQ1WXaOINJfY+t/SXdtRr93A6j3lULWwZZhwUOx9oPl
Io6WGt70tjLNe6Rweybj+nNQQuqFuWx+FMN8uXQU5GmcT0r/WPNHMFRDM2sgdbtF
6t/tDWWlfsqlttdoBLf9eftdtUY5Yi9y+A2z9xibN3fov51hVtNLCpod4o8Gu8Lw
0lSb50wkTrDV0biiwxzY7Cm0A0P4ws79KDilluW1b2gv/VCHrbSL/j2VR4tya12L
7iH8/XGhxFdhe/F5C9xyMAN0D+YLwnl7/mhVxUaXz5eZ+qSc6hjGWBN9KSZg1xhl
LvFT+c9CFvtwpchrE97JwaM21oVyMgZ6vnwFS7a4dwsXjGxIiomY8HYHd/CJ6yFU
uegJEauMmFtTlbS7a/Meeznv5wCtEvkcmIf/AAEQUOHcw2MmZIcLr2ytf2kYxnbB
L4cwN8r1MytazPbcYGbUmJQPoRkNqnuFxNHyEkdvD3plGZeDcSDlY3/cRPqqUFWB
LR8fUracl8XSgTQBMc2dmA==
`protect END_PROTECTED
