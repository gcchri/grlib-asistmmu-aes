`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D/ARGQd0NVHxhN7gv8lLwoJ9TXl1GR3vS67ESLqzJTiGWjgA9EvZJKDgVNaE1xGv
Q5Z9G38xGVnoYyXj251f2wfc0dOzkchfMHIR/jOwoPR/K1d3TXySdnAYfV+jUpwl
6AL4bGm3k+llasLMNdFJdcYvBrbvMIjUj0rGnvo7+we3vPq/EhngiB6x6MTfxbV4
me+wh8BoNx+viaBUyF02U/tMlX8Ykw8V+Lc9VgCZCSvYbCob4YP58uqKRsc1SJ0f
FE2kPc21g7+/5kQsV2CUU/xAiQNM48LBb8ochy/jKx1eev496LugikdoIeNEjzyr
lXUYU4G64ibPnYdPI3+6LZhQ1WbAixzDMYb0rFdCUOYyGnsSqbHQMRy0qM1fxwHs
+ukXlGOrTjmB1bV2y01ImtKO7S5jAWjw2YdI3pG3PGw=
`protect END_PROTECTED
