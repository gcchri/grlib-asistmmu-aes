`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zQJcbALA/t/VmrWlDyKVMbCDnJpewELtkE+2NF3genXglZ0E3B0dOQNyEioMPrFV
BIbODa/AJ666W7h/Tcz475ye/AAEK3hT/8veYwMlDTaEV5SLox/nafCgs2A2FQtn
9RQju8b7gJMvv5gh3kEWbDV6IwaQC2XhYTrx9jQF2yEbobs6JICn8hPmMOcXrkDp
ocEiZfaLkI79RnsvIgqZj38P7LcjuBPlAFc0A3r6wKo0T8cVr65BdsBtGdq+iouJ
upEoZXTYJg99zLRcUo0o5I1PqKUCjvOknkWA/8R9IOb+8iimhkNTYn3AJpL5uSu4
g/JUQfgc5WhHHRT7oO5eVyRBTXAHxQ5kPUpma1oLtr8GS3B39NmOEL53u3D6f5+x
ZILYvZTMh0OhEY6p4GpZBlwuTImVHr7uvfOYWcvA3PPQwtW8twPPoNHDM5RXIsFb
7clrCNkogAoo3CKzssWQ4uSMi3mU0RY3pF9IuBlVUF933ERIzpwIyngJJeufte0J
wSkMzQhn97f55XGc0iJSeaGMyTHKaL+1RZmXz10nljRew8kPD39sLKoHU8Ivk1HC
YZmYbkHRGItk1XNO9voUUg==
`protect END_PROTECTED
