`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YznLg5mzo9/OuApMiB9Rwjn9Ihh5qTaeE0ztlc0V+UyEoO27s2UCdhKRoMiGmB2I
XSyNnoy+Qw7yoaV3yg44QwbxAKAbi76CD/fvH8Aqm9khlwCGI+XERp+vbiH4G1oD
kc6ImNCY3yVMcjDTXr963PVWbfDGQriR+rLj4uUkNVqEPRdgQ8aUagFTsDKhVRAQ
dLk3R5o4Ir4InQ+y/FhsswPAXBHyd59PyG+2hmKGdv5F9bEP3J/iwG6vhgEFnLiQ
6s98WLD0CYdxROimNB1iLm6J5OQ3ewa5x0SQCqqJZ/YpB2/6KMuLHIgYg6118pSn
8TPKckY4m9fFLv8QcrjVrStbRmXu/fhtL3gb8WUfoQS+Qg1c3PrujxVPNgF271ft
roCwaEKygKjTh6Ar1fo3grH8BCA2+HsW1gZv6h86qE4sQ/DnBZXM0La1JIH3i+/3
Z9oTMm+rsE3GP4NQIi1QmUcB+bPrWzWEScLiUrc3QQqdeTQmnSR4bp3o8uqJCQfX
GKuGmDVmkIbKuk+R2vWxOL6AexWmrjWwEkfeb+Pbte/xBDXY0oEpm8aXFoSktcp6
ieaI4ATX63ZCtko5TcmNuJqyHx7TtscJQ3fJOOTaM7o=
`protect END_PROTECTED
