`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F2xsBR4wJdy6J2aA5S3HOlUaR7m3ORTl8eA1lrJJCk9irl8Ze3qYMif8qs6X6mhD
s7V9NaJK0hjC8WiWBcqhXQykAmktV2R116K3FFygAfVhlLFKscsvT0Huronj+eR7
uh3OYJuJJUMRFfWOYdGpTn+5iqs5rEYdaCqQa6DyOnz3zW7pWguF2+Ds03Y0LjkK
FMb6C67rcBHbcIygI2NI72SxmFshcmKlnRXySZ0vs9J/mJkpl1BRPlObOqWBZSu7
gy8mlO6OEY9AchgWScmL4UPfH1WYxBcQ//xwMF7u9SLwY1xi0TsyWjnE867QdU6B
UrlrDGCjiYEEyncNdceGW7Z68C2Nr+RXgPP+jJekEDmN3R0W16Qe0fHD1m3sn3Hz
m83rWkfzAseVl2eoNcuLeQ==
`protect END_PROTECTED
