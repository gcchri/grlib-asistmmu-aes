`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xbP9w9Y7VhlOfIXn/eR03onUL5WBXhM9E1DZkHjEPDPTI62g7a/1rYGcNXgCfGxG
/1JEnb8wA8PqLo+nebUm2ikKBGkIhHhuNAVpD2IpQrNqMdSrQ694czUtiFBKSwmO
+gf88OljFkoZwMr0LeDCCr7tK5i2CfDvhhOJjqkUk+vbeoTz5VQj7iAt2WpB3Acl
AjDRi0QKILXBYhiYTnbm71BeFCRTV5CjdPZjSJitPW+1HlDVFESOVAjPKQ8LyCdd
XeOIzwgg7nagIRaqb29mtPcKGB33McsURhzhroLjqIpcM4AGsBJlSZ3wxuzv8c4o
D/F1DiOeG131EOhs/91sTxSrPd21vo/XFRLlz8a/Cpra+z6NFIHJU/tMfbEVX8ZA
4xjPrVXzgIcq3vT1b+zyYgSwW2EwUa1qLvdtzw4ttBGCGp7bqC9dhymoHe4Z7gSo
W3VpW7gzHexqNMTwzBVSxM+uUrx8U6Jh/AexBzaUsQS5V3WSdiBIPL768OIF3l+E
pnaPcvfkSIT1RFpAAmozMfGx3YgA4LFlgxm+Spz/4QUUJz71Wfg2rYyQBQExpptW
aR96y/OSTXZbllCYobXnn1JEiSNqKEE6MSEqQT6Qs+T2oN/bWeaxsarZ5nKr7jGd
RRRFOBwEQJsE4qKc6bFRfPREk37KRQTi6tsDnex1rKjP/d7s2g8uJjPKGTutqGab
WxAvEoKQbmszpgHF534dTVBBDZ2RJCtHVNo4YoJUGlc9HcrKtQoPYQBJ6x4Vmhu3
ANDjY/12AeqfTkoysYw6PSEYeKEQntlAJm+umKVEbfPxDAIc0w9P4jDS2rycDZCW
9dsYXIVZs065zOYZqkanIjKnNujfEuDPbI9LGXYqGm5AQhPHH7TJcBKE28I1gUIy
WVvBbIKUIK7z7EVJyz8WAagpgHJXQQck3DIovt23P+Ss/8IcI2XiGKerWynf2f0j
XZkGi0y8/vrghVNjAbBTV41hvrDUzJKf4sKCsYlbRkgaP3Fn65LMkyCCF3Z7m2uB
sj66W2PuLIIqHBSktjZ4XJ39yigSiSu3ILi/mYBcMHTjSHtvh3OrucGfd1Anp7Ew
CgLUd7+jWLoLnswhVhMZoi5BiXugWh/jMbNeo1RY/Lp3kqAtdaX3BLmidEdw2Gl+
uNvysSdkgV4gJ1k+dAZOzK3Z2Mlp4JOlmF2sROpZutZY3ck+tQ4j87V+9RFmJJXc
AS7DKlP+0dXbv9cIJRTPB2rfoW1N4nA9+MBrHUOu3pBIsIlhSr/6j63oMPl9dDaO
EvDPfdOnPth4cHxSpfbYmODZwp+G3FUPYRCniK3HQ2K2N73nOOcW+I9E+GHjh/kI
dITQizGGEl94svmGPb71BV78a1GTNNmm3PVkRvl9jBx+cxbiwa5iZgEK8NblXLBF
Vh1hXThH/YFnyfyYIC3HZ5SGutX3Yg6nDqx2E5IYFVdKvHI/GoZBpySRB59em+mR
BoyL7yl95NXwOHL3UsxirwhA1XLlh0dUlbGqGtJQehCRscNRTXWJzHdcjs8XgqTE
JXgxHNdoVLLCiStRNUwR0hZeqgn4nKbtJ+IJUKV8bCtNygQtoO3r6VjUCxxtVFoz
Hm8CKFWMPw313J1+j7iefCb+PnWeozfrK0ZfrD9MZ1/GFuT5HUfi+2geONLgGYsX
0cKX3I+GdpwfVBlGZwbKchROyF/XntNXtiFr+2HzSJupx8csi/rEtDgYfZZOwVyP
EKmO01evos4hIroaBNFJNWsWo93RfoxfqYohVpja0s2N1O6CIMSImI+w88bHg2yS
T971cCyKX+y09K03nisTFJ6uB/3d1o2iCmLraOt3TD4u+RIUZs2hlWmdJDftg9pP
mUpr54uw+VJwQGiqpCtR8crxNQ/SaF3hqSrOWvuK2ewwmoT13pmPlkky6dXd8DMM
2VJ58H1g93qhCbU4JU90gJF1fRtUEQ43d5j3TqY5FhiPT7KO2v+d1dvyQN2YPQ3d
BfEp3sEnWIPLeYYTuXENE3VhKyqMZhiabz8Wqpmx9XkXPodiP7qgM7XpPRF59nTX
woapSbnbmzd7cRSGhg+XeFqpjeXvKVzJipFMERVq/sE=
`protect END_PROTECTED
