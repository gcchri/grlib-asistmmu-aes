`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bByZgi4tIgIkbCDiLxN6J1alaQK+CdZTVInx2v2cWMnk05Mvrd/cz4Xf6j8bRJui
XgfOB2BH1QZ882ukV9YKg8FCnkRq/zjAMWyttRUjDjFXtKum2zdmN8fTjyxW/YHl
WLHXHUQem2MaPHz10Ha/Fj/clJxMZFW+eLWuvSbpS6xZa9i+PtmNYB8Iydr8a75Q
F8p/ok/Qb3SzdiXUa5i9EatPw4uDodHBZ4ZHYP71NxFnqu8mJhLj156Jb0LQYstK
fg7FVXFHVEeRO32p/0v5qpbQvmjbh3jQVhHwVZjOADePh7g92QgFihgM2UKwCIc3
u4+yrRyRBFDlTtLp0jFJpakLOG8XuXq2crTvX63Fjb7iwxcasueLei3fElkMfwrS
pqChiU+M/hs8cjWfy9LXyyv2w0F8bHNSVuD4KyXuZo5pYE/Se3FOVYF2mE6tlLKb
2tIFmQfYtmBFQcxgcoU3RZwLMPTMt0LiLgrA+JZWfFT27EimHkCiiBKQSTRsCp+0
ef6qzQfH2QDhJYdKK7Cq6/UFPEjhN8Mse0AeTVR6GQ0wESWdaQ5eqSWpThSkLFPZ
u8bR+c+/higSWPvUKm46MaFx/uyZWFbgqHH7hOjRVdU=
`protect END_PROTECTED
