`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8JMOi/hp1COUFpMfjmT47TtRRw+AR4PrJIqEbX+0vx0bbLAGuRleEaT+pJUZI6k6
eY9K0q/yHyXaJtDS1ig/Ij4v9aLDFuxB8RsVOYchBataO9B6zL2TBLIU8zGkyWny
HTj8d/p9eQWlBxjpA2Y7Hw3Xb5GEtDNwU96cmuNiZaum98shQJKloPJVxfbZNRVX
JL4mEbg/GWFN59IdvoIh3CLejReiCeQ4IKRVal/1r+rFU3f+4H32D9BqcWvEXK+v
nOoMWQsum8btg58okrjkD5ih7D2kbLi6ID06jSq6SeHkQIiwhPhOnfQ3t3ZHyEUT
KMdVsE50lxJ0GYQeR9R52yyY1lwSOKFiAsRfLRn7dNGOBZXnjcg24genT63JierN
BUiJy3E1vkHgO3qMkR6EK90IbWuzc8dc/6cuAqA2gUPvWpNT2CuN7TmaTMv67otS
LsNySxFTKx5q+yYdrMTveBHroOjxq4FAAXtMa6Z1qywQJYqLlXWYbZmkfhkx2Iln
oXZdJxkDumBp+Y9vRh7mx+w+VVEH/ljAmAjTP4GJo3TxLscjwaALwEePRY58uUnV
cOmXosXZF7793JE0YmxJTpM3V1R+bCX7PiZtK7Y2m4fNLIWYEuEWCi1LQ4ue7+PV
lx5OoEPqBhvHO9iSprpL8J0TquNc2ZEIlNDerJ6sz2FoMp7X7wiL/5TUstgF5B2s
PFCfHMbq1+dtZ/nK07sx4UiJNgeCFixoGMGiVI7umhPfSaubxSDfbSMTPhCPlrw9
vyVyA9V6n1qWSqG3QOpYByAk3H9zYr2ACkY46ptApkO1iZbWSAz1+iINTZXqjW7d
/hbg+MqS6XxS9DfQ92HnotKg6rYhOHETKDEiVVN1ADq1fDkNlZr0UbK7SbA0PxmO
xvikkaIWraJzDjRA6bxVX4X2UecjGc65u+CWizZxBAN22tQ9Kd9cCprWD4SXi5FB
BG1XoIp9amWR5DmOWpBldd7VQM2tfjadwqpDCA/OlLWujMlPXCJORqXZpw3xvxLa
KjO+UMn1OPJ4fef0GecDxWSsbHnvRr4LLURXqflQtceveCsxKWoQbM1zk+nRHNLo
dBo9O4cYk4jhzB7bgJdn0QlilxF3nP45lXcz2tgOf/BMLG1sQC6d8+whipuXZcbh
YBF3834gFkoDatHyRLOOOKDUnHUoMrx+o2RQYU2F35vYWIiH5mm0ayGUVxUPQDNJ
2v+tYVpranhC+VcinlcWtGpFvJ32Xhqb27HqOhGeb2JtvGGaYPfo/kcwstEk+IM1
EhvEOeR5b6TP9qQUGyVlspbNLEiuVqYXMRhuVBQxNLIlrbRKRFd6Z+xU7AF+Wee4
RQGJFyjFBggicABu8esrN+UIt/KPFeWgKwb7jyTLRNBM+JhlexVoV8+7+gfRsD0q
12kKXYRvc7S2Amp5+jqHGlnMVTAgghphHsd3lPiJIYsFQF7XUG11smJF/Tk50wAa
fgvtRRoXI361atst33mqEUu6cgh4/igRHelLGADxGlgnEUfj1mVr9+DLH0TJ0QEa
+7WOaSHtXqoLRnSKY1WRvnSBUhXefmkmy4+U4vhVPnw=
`protect END_PROTECTED
