`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rgAtgNrkePNYd1s2QOLomym5lBQNyMya3/Iq8666dS56WxNKMtGAHe2woS0wd9OH
lYP0QxG3QuM0QBe9cFNME5lop4pGwSXQuwPSdRr/f0pFnsGAqfByFKWLlbwQYC/q
QDgKWdRAbjHy4icErOta7sp0rmHHlVtjUC4LCHw4grFzfx1MFfm4TqIo6uX/mx0/
Cv//hN1zy1uIjefD3uFDkrpRzcRWS1YDIIm+rfSRXLBJ1tmHYkA6K9+VHWIV5+Re
kQjeNbLOGN6VQzVfbj3ln5hwUJh29h7QXim1POOr+grMv9bS51q530ppHY/uC/Sb
`protect END_PROTECTED
