`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JE2RHNje+mKOsJeDe2eVCoZwjwoTVp3qvzji7KlaOjDuft1sXHs7qpVi69ZzNQSl
QZCg89ywcF37Tl+OxWSbaXoSzNcQoNOspRLP+kvEenmOjX9TJOb46tyJn12lRcf5
0p22abdGNRwVc1+kpOBIsuMDqmdtw8p/RJACjSkTAmNBpMthUyuGRBUFCZ4pKyS8
wlUfdDmkdq5Ouw6qEtFoPOspIla3zAFZKK8L+FpeAyfqlwzrNRDEx/TP2E2/oM7M
hgDz+dlABeIJGamNM+sF/hjNUu554qVQd4s1FrD8hj8=
`protect END_PROTECTED
