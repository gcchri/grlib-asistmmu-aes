`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zTqULHbg/fHmGQ7okCvjEZhTDvsFFg6XXKjSzW7vrEhc1JOsYC0qNGyTXDXQ8+7a
wNkw7LLko1hiCIg1QPByDhn5BekmU+FD1YXSlWYruQxCw8jrD+J9WHuQfWPqDuYK
tl3R1Ewkjoj2KBylB++M/U2U1h9j3vVCfT3Ip0NnjB2WWwZUE5bQouIUisK8Bw4W
0PEvxw06iTeTwYYOgdMXN4kcKWuyg/o3UoiUC8W3omIuRNEdSso31u9i6IHUq/W1
V4cCo4FCTm6uD2bomPcADzcHXJSrdMl4I4/IwVEtmvLlVvZZbQnMFSMRp2RvhKMI
M1j+1nDUCQaqxb0IUn2sR+xEkoS4v8EA6nKnX3Rqv3mn+HTUpI1kaBRxJELTQn6c
ah969ccs4ZYCzdU9/Y74tXS5PNeMWZ3be8VxxSWy1NbPGK7XLIPWkHqxqP6ssTxQ
RYIgCOEjARIFPSNVf/pVotykkfDc7dCjsErGvXgLfzA+sW7tg4WfGV8Hnr9FrZtw
SeCyisXu8hWdql0T/w9ZcZPy0vp6yQI5XKgwZcnxP9A=
`protect END_PROTECTED
