`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m3ha286jLXjixbZih5PScPinfiCnBk49zeYbHjHS8mPIexuh+RNVGpgTasyEPZAE
/lLnrePRsN85NqRY0Qm9VKrw+ZBmkLN8aGOQCcQMm/Ywsh2KVfUBxQukky9hFl7R
7M3gehITH4qq4m796VfrXiMtzOa2rVBlLQXne+0AYqiu99Sdi6quc/R2hnyyl0Dz
bM6vEIJmQ9XOmdr315F3Z557yU1tbkam1yo3xzGcUUvLPBhbCbtz0CdaetAn1lN1
gUZAeksNqjD/sLhFu4DY8SXmi8ZHgrW76JFe5Gvi1MdPgPnlM8mx8/0vLiH92244
vwowmtZKWGbSHj4SrWXpk5suXT0pfH5Jyg3vZlOgmScKVnSODunG1Q/dDqKxV2sJ
l6lHQEJreSfklumakDY+fXH1gL/as5CCgdDUxAa3D50e2dh72K2fnDLcdFZSpFkI
0bE4HM5/YMEk91ohuXKmuxG0FhchU3VewwTWg/VjiE0dONY2ocorgL1Cdkb+RiIH
8LEHdRMyjCLpQeK0rajWs5gMwsHLEkkGPl05bJx3I6irHljaybSVq6P5rUKpv7LL
RpW+6lVGs5Z15Yi8K4I8o4OlkcxWw0gkueNRC6u/NYeMzAkz1yOMeSxi71O64UP+
B4xjXkTAEtTRPSGrdasCOVIciWXP4sVp6EDEGnXND6xq0pP7YMwbq/jH+G49LVLm
HruULUqXXxeLSpOxxBrUpVPtOrFZmWdKOzLNrV/MDwVOSl9zQn0CIY2jKVVzfCEA
P42DW5DcPLxRPWUv2dkubA/Z4nrm/Pn3BXcf3xyhJ3Seoei0fmARA4ap0344NtAW
BuDMzJpbZLWgotzReC05Q88Yrg7/Lh6fbxc+O0ZZZs/AaXJZoHlcynMJ6HFKKaiJ
VfVoo4VjKR/4eiJOG0yPh1MSsTdkSz42CThUz7tf5IlLV277Verrw8xceHm2xrTy
`protect END_PROTECTED
