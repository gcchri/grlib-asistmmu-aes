`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k7Wy8dRD9GKLkOf27aPLI56pUxH2HM5f+1zrAfIs6o6ZKkadj2gL0wbIhWAsFNSU
RilYT8BKb1mM+Tpp5gYxSfbNM/QDWAj5u6hqbhNyofL+g6UdmAxqgohvmW3nWBPy
d/l0vidKYrt3FpFqzrCtEDPpuGik5L7+1wmkmYigsaUUA2fXnV4TrBdPXpzNrWZz
8Suk3zGmPkZHweqcu9o/cwQPtXc7TmOjB58f/uz/5OClgNHxgRFrphQDBBZ2ky+x
L+TM3xR1JOJHbI1HKuR4VsD2SLbsV9HMGGqGHkXJY/EKxVDToLgD0bxreOMQjL3E
riXoVVLa+T2/jYbu6oKqZykdg+y5+LgiqE5f0RxSmcTmU0+OLEoApftRCwiXS6Ji
VoxD+iGpQYkg6lZ04Ez1twoq4xh8Hi6TT7uXPS5rLgM5Jzl32xQiEad0HClT7CFB
iNfS6W3WsRBcZayylTI7t5xwl2wtfaV8seswFVZPoCeNsS7VACxSZqaC8EH42Av1
XjB/lAffqwwnkIRWL4/gxWkgLdWvoa4stlL9hV4mvDvtdbPyjHOVXScVd2MRMAZ1
v1qU4CJlurcWA+Sv2KXHLRVzETGnGuTRSMypOaJC0Vk=
`protect END_PROTECTED
