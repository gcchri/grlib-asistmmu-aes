`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M5M7iU2myEikNYX5ew/DIY+1vMni5px0Q1FtaGO443tmdUitFL8GpkAO/Pvk4dst
En2uybVuicLnxQL7H3ktBzYJtolCFyj9v9SF/Sni/iFbgzS5EVpbOyn8/Xh0s2kt
yugBsOfPpC5Bsnyk9UK0o0jYBzJjmhfFcAoaZ+1Y2xsfXssOAw159ja4Kww1X/WX
II67LwFT5e1V/FQsd4w/4pX01tlEQ6PHSeotXi4aIt3KcfsHpZ7QqW17uSNYGtXh
Hs/WBsKwOKsX5S3tNeE54Sduu3/XJg6JAfIMZVFXtgATie98P1EAm6dUZ6RQ8xq6
MJqREYIhs8/TuMrGk/ILvmh0V9zWqZz+pf3RDQHnYXeawViOkfNZoKa4C1VUtlGM
VjXpYBrGCIcs2/uyazYKNfNyt/3wvNx0K+WVLRG8fm0DekXiywddLERIMDj0mZAB
NAVxGMy/Q3MkGMq+6Lo28zDcm6rdJezUney0FF/2OuwlubAzRRkyBsw8ZhkZ02Xr
NtPJ0OWR42a7T7UQKTjiVo+rn7WmXaUCIEOk6Ik9HyKuMMik8RnfqWNbQsfBlAhD
N7LS9TdBeZAeW9s/FK2yrV7aw4lW54yzlHYSqFfzTxtMIm6IP9z4drpceYZaeWBc
AV1WfdYThyUMud0zvOu+O9k5Lf08/8odL/FQ1dpdgZubSpH5h9+3hMoClYQV/xxq
BNjbdeXDt6gTqY/zyd69eisU9VXcRDg1sOPSxGfKYkTUF7MV64ypGyPLCSJf9VRi
RBV/0JJlXbnBPYQmuqdnLvQ3kRBrTHGJ7KRcHyLc9rJbAzISXYHSAtQFDwX53zme
Y6u7DGjsyZs50BSwrmBiyWLpkdszZgr/26/VEYevIAOKgF7ZDpFw5zzTVxobpBnm
rsQ+7XapLSTO6ot3WGXstw==
`protect END_PROTECTED
