`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RdeGbqZdcp6ReduSwzqzDuhP74p0gPyap4f1AviDtF4ox+qt2cTBR69n250GtC92
sez+6KZJQVtlmEwXNr0aJkmtfOczNPHOa4MkXYKVnat8muah+L1AslDsKtYeMX/+
k1W5+e/Ys3i88TXBkWz2zSETsPf4AZvJdu0qT13+qOlo/EHBCIsa+QCWt6SlYeYY
1gVp0nhz4pSN4ljdIF/zrw==
`protect END_PROTECTED
