`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BadKfzZrNvhP/Lj1zFN/lmlPwEIkSSZ3cX0LHg+HN53oL2hdsw25n1XnvtATvw0I
AJHWIcwlJNMMIZnwNEKYPpQnhjTkDARJVm+am5aSf8gdInP6XSCpyMGDfbe20l6j
tmyxmXACxp5EW9a+ctjVUtX8tA5SzoVlIL0AarqMJCQHNthL0RGq3Awvur3bzX/U
kI2/cERyTh9BJVan/cRr4TLIt74PNfU18jPaGk5eFxXeGlBjJ4LXB3I2vTSllVt5
WQxra3P9xU532FlV+c90mx0AuD5OiGhxy6SzAnSUYZCET1oDUQm2SLIPdvddAoy9
jdLLEHNxSPd+ehqGqNGouA==
`protect END_PROTECTED
