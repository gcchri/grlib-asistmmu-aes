`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u7lzck3v3/xxK2MGY4a0CLhgwMXadCNqnO3aucaoXfyxJKSo2NDoGWoecUJDrhBD
NlJVJviTP7S02YWNMc3KxhImh9fneFaI/xd6Y2mqIXfh3SbjJksM+Q3uLVH9xr3l
5XWGWtVIBdi2lGYQSHgMizNruukD00aT9vsziTMz/aXfjvKUvF6dJesQWtQO9IK4
1gf/kBTRhA0uB53c1fZPUB3Q7vGeDVwECd+hTMbNQxT8TQqAdGfx0k9+bXLBZ4vi
6qMtSfgay0/07MQjgTRIqZJo7SoknHhvtKBuZDAzzvTfRPv0Jrbd+R7S1r6cV7Zd
17ZozxRGwu4Ixn25FGPX7OCYi2tcsx49s8unPiHJ+3Qz4i6t1AiaEcAuEzUNxpci
2XAETbNQJS4Cgh1sOnfiR+vX8tn9eVxbDDj820/4wg0MSV0tng6LeOZU88TPM8N2
npDQiQiwxeM0yj5DzcxK8kWIWHd45rmT8cosyGxeCtyztPny4SMiQsuZxYIYS9Ad
sO6lyWdZU+OMG3f8rvjhhmQy+7vGYiOJDdIOQ3IbT5+1rhFv1ccdRGIaLUHKIAn/
IvJgTRb1mS6wz2hD0hwyF5+sADpIacBLEjRtIY81VnoegEXkrN6i17Yk2LzG+mOU
UNSdXsx8bFDzptJfsqs3CBCM7K4i0h0D3aoN9Wm28IW0q/3bDPqDP8QLQlV9DFpj
Ff+s6HsM9/OO1j/3plTO/8jRiwYk73qTVeJpcJ/lZM+c8MAIVvtL1IemQ30F8MoB
bhRLA8MYHYAWBgPf2gg5ECjlyTFZ+s8UFI99nCb2v0kfVziwkGecfXoftghbwgzt
8DdcdWfAnm4txWn+PwNBGg==
`protect END_PROTECTED
