`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FyzhOHSDEy1/qoqHcIsE9S7CSWL9PVTgSzHjrTNCv+5hZQPX4iTen93dN6C+BinU
hSZwS2BRNQROIepGvujn74t0Rgy3LAu40+3sxSjhqTmgIEUI8n+ibGLawyNUKFuD
V2FsF4Z9pugXhat50eRJNoVz+neDFZbpFAAbsVniUcHXGb+Vf51svA0YVd2RQKEF
G86YLzR2hqOE0UdCHjctnxgeFZLMYPS7dprZ2yB/fdBxd2tOY+ohoKMVZT/Uf199
XeiaeStk1wTZLtkYLKPVbA==
`protect END_PROTECTED
