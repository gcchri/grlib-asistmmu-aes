`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F0bAViXfRjV9YYO6xXvu0IIVYNr6lpq5Sw2eHEUuFiekCn4CxXTV0PHqpnOxRr7o
jxjHY7A+Zi6DaWFXlcsREtCNgGiPAIur8zxkR1OlN9KCHgOBUul9XgEOLAJ3jQ4C
roGLtFn1fFtm97BjnblidIzOWKfsACeQTgNsb3i+TGKX/TAUiXSjkJmx3Bav4wxT
xDNNM1ved0vsOEoc+n3kk9JwlGg27tEIOftKDUS05+jpgvUImN1OmykRQHOSr1R9
aSGN8bk1Yk1VOEwwfQSnUPu1wP/5Y6ytyU4nk5cote58sYbmEOvm9ZSuFZlCBBR6
kVInisTc0EInB9jMFIg9fgKJ0hSLzfJBJogpYxlpx595eljFP5QzBCVeb0iITcEP
h+Sp1s8xuAL2rhdnWP2tspx+Apw8NR/4ntOk7CHzVgXPoN8MC1OvXGQsLroqPTLg
LPBIJIgnA/iUE+EbdtPAlcCbHE2aAgRzF1mvIffuvvvSHf5j2nDwVtBe8eb7DIkX
9U9pRb6ib/5dFbDygTblIoKMgAzGKmlXQgQ40e+nCdCRF/P0gPVqqWxtuKsFHkGg
ikdq43pZ7t6ZcwrkzxAWkxAipG81LiPdRlYXPlg+9+gE/OJ2qa7/553YPcArNPor
s5IjN451DuVsIzJz9EMdvFEPhOTqPLknlSqgffnGrlqxAJ/0OsI6D73lap1WVazs
iqUMNrBRKzOLwa7eZ8CIe4r4VauM3u2Ffq/oUlIrk827KXjUsD3vblNQihxoK1p7
NnGQF2DzpJCfHgO6VzPJDd0lmQaKPNG0fsUw2HN4j6ASpdk1JEUdGsTsHFXtlyCt
01rN+LLgwy4I+pkgkW4dws0ptPWzcEI3vURUkRKDeOkvXOsGtWNd4orgvTzxNPaN
LRIYmRpfEjbPiuoycODwlJL+jS6BJuJtuBGy0qQewxKVdcZXRcF93hyYtiEiS7q6
x/Vmxb0VqrX5FSz0id0D8X630iY0sIBgJHvE5glKJTs=
`protect END_PROTECTED
