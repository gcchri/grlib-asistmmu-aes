`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BEBEZRtNYRn4IFmxnb6cuBGL2r1/Lzuxout1fYdfWHWPJ1VmsCx8RqNsZ/QTooAL
PjEzcpg21CRLBLBdVeG+czuKOV4z98t3KuVAaLkr0H+SfuZuNPrQniiARrepm7p1
l4aDVyHifkkRFLiloYId02MOxDT9BMVN1fX8oh7zToJKP6Rp6A6LdcRhJUOWi8dI
GUXjVfo0STeN2DuY2OTQ5opT4tlmwXftjqDujCMb2/75QjzlhbN87MQA1DTpFot3
5dLsz3gOk0Yuv7+WrqDjVfXz2qMqBBfcaSHnl0HA51e17VvVSdK4OYj49gj1R8QA
Io//XqjawAgtx8963iqVZfiHCuxPF0/+4k4RaWy3xJ+eNYjvSkoExWAV5conTPXm
VV+ZAHy6gdFdVZfWLOeR4E4pyoVbuSEo0eYyJWvgCuSp/WScko5raDQtktVN/8q/
fe0Q9fp5NXjgsDKq4mYhjEqW1KFwTvAF2Et0rOEstEY=
`protect END_PROTECTED
