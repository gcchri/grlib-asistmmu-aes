`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GBe/2KJBG3KDso6uP2duwwasBa60FnL0b73ugJ8b5cTH2jg1n4HlYXstoO4GbMmC
IyyJOVLuDUg1wN6oW+hcD84NXQ9KF0mhO5VeTlr8bMPOpUDEvHoUPKlk3bynH5jm
8YyqxopDP1pcNX8W+VXwYS1CTvlruViBGznzlM44f+MYFhGVPPB1ZzVgAzVjJSFn
7zE4hEoFJJswHSFBhwFkjg5MYT7jxL4q+Iqt7eAz78yRYYs/bnx03ONSyDgRFtwG
rfzy5uUAJlky05he5/DWruoPw4wMLU/cH9daF/ARf3ia+UAVKRlFxA7PimzZ2urJ
EsQUr71tinUgCO7tIdg2oC3WV5AaIY4eUDWzGbkLn7ylR7sDhE4C90q2RTrJk3Yf
GwrvJTuSeqiKBzpC8eWPGmZAm1gmrT57BKxMnFf5jw3LxDcdoSNr84Fz1rIyo3rG
IqPpRCxA/5Y7E/UrlyRKR/Uw52Kaa1+/L0KcHxsdz3MSveM+P+NVtWJFo7xglzOe
eXSnPoj8nkS41MYAg1EjhHgctG3Ifj9RH4hZoPpOcJd84aNnuQlOHdUM3tEXJpYL
him63snixkRjnFFRBQ/lVzN71PcIdotxfonDcsIY+mFowqm9Ebon3KOprfHw4o4r
fxAD8dA9f+XQxDC+SvHOQ75QiOi9+uklRZZP0uHmMe/45NkkIUMyUwPdKe1C0I9B
KGX8SSRAx8uxLS+jp9OSrDkI4VyAnrxkRybb8AOffgnO6HWpIg3LtgrMuw23p64j
DAzsWmzX5+mlItDDapAkncpUw1DTobJrV/hZmc0+8rrSp343BSCZ/yfENALWwffl
8NYqDXID04itrhk31HJUQkRikK9e3tqIYQ3x/0Y+ErFIuKp8k6IrlVhNXh3e20KV
NcLPJ6LCo8U7j+h08MSlKsjzedP1APFE33mf4xfkXNbO89Y90LIHSp6KTeR68zGJ
ng3I+IvV90YaLy/R2IWqQT8av4yBNvESKs2BHn3FNyx3oVavyPitjPEo/pCY2HM3
prWT7iUMmWhfbAbopS4BToHuYFfZZ7dCWFjGH56oIaK5O5GZUcT0ge2WN5z6yFaU
pGixESZ+4NFM6SJ6gKlul2/1nz0qb0jh1oliQWirD9lqjT0aG10qAzlgKFbfk/3G
ldhOhbxyBAGxxIuiGyTjGoxpy7dOV0y8hyf04q+X0PkPjtEkEwQetf65jtq07wmr
5y8jqmS31C09JsRCZojGU80unxLG7zWA58rZ8ZkjuNP2Bcvq0aR42EAW/xv5DRRp
GAqWzpio3KRqnC67SAMfur2BKYwmCm7Tvk2/TZqiOv0xx5ATPxzGJoVjNuG+LPb4
PlDSDkwllr52YkreI6WaZslHI2yO4yNyRhOBNEj1JwXRTz+t8YXtmTbZg42hwm2P
YBZuRttEnAmqYaVLo5+e8KcgFa4/4udwYaZQPMCYPrd8ay09Fbvn2M2wooQK1n+2
bMpV5aQTrouMjAMjpHNZik4UdXZbW5qZr+suLrcN6k9G8o3jzP9wX6mR7OHaY+3h
N0DdzQo6zZyvjo/nfNxM2RBjPFmFfwYLR6yysVSJala0ruJh8nzCKIRh88s9/fZe
zLWblO+anHmY5kPS2XXa3g==
`protect END_PROTECTED
