`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lFxRyy/NGqqQeJq3BfMv5hBNIzdwQ27FTHCxhey32jMH2dUDaIHXBVH/nJ/3IQQP
F7R8MRRw4fvTBc/BVp7psqFO6ufPNyVSgj6MYKpighXEVVc4FURryDK41W8l7zBJ
WrlnZ4sKarIU7eIKVic+xA+sB/cC4CrWypTz/XRb5OlHCn/e+VeRha4CUWgXui9a
gkGRT43tP+2G6IXjoUd2dtl2Tw7Rt8t5/DfrKdbEmhPRw97K9quqgQUc7+7Fumgz
hUi3VQz7MAeZPfQEGcQlLjyCzI2iwMYVyYdAK+KmNZcIN7SDqS0S+huCVL98M7M1
c5Vlh/R9a9vMOIHZ6BvBX8Ay4g2VuXGHT5K2H9mTlwSp1Ubm4scXeI1x8dwu7aWG
8nxLnVmy+Zwn4riQV2rHcmclaoAWNDogdnuRHm+vqRKLFUIamhB2ZeRhs8D3+KNm
hY72SXEmQpLqhXrOo2u+CFztkMINMAXd0b2Au8oC+UOcwbJmHd7U5765UIePFKpR
OQ6lzKZhYZRGbViN0WkAtg==
`protect END_PROTECTED
