`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p8fawG+lGcSwOQ0m6mi0lU8evMn7fNl+ICwiBljwQST90Q7zyhBFMYelWu6uxNuZ
lhWQT//qWks9TeFjKe6c0JHBArAqEq11Fy+Jz4BYTSHaomCOdW4kvOQkp/p+Dk6z
BwAzjcK2mqMjG9ewDvnpsWJVFps2LL6dI5Ei1A4MTjBMjUT+qN2ZvZcRhGUnrwbt
/idwl67vR1wLMoVkfFvQiLx8hyLVyxiutN564wE6+RQ=
`protect END_PROTECTED
