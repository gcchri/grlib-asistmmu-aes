`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SoXv8aYU0B2LIyXNnDeUmkxdgW/Adop/Pb4poBt4gTpGmcm/KPBfakcOJbZA8tDx
fz9qKmANygVgFxeoSFOC41mR35vANdWl6lAyCYbwyMQD1SjDELelWV/mIYssLKSz
bOnnSAAn22m7wmdWteevpTiHRL0pEOOBL6jH/FZXnnesjtbB4Qg35PHLOXmANhu2
Sgkh1Rj+XXDmzHSshAUy5TfnQ9fjHk5Ry2Cyx6EOXp9zZpSLvPCWujoyNrf4ST6p
TBepXFHJYsjQM+f5dV2/Ar7hUkrs3GnDmLpo9iE/oFWCzi3otKcHAE9wdla3Lnqj
mch7f23ENMhjSprS9oHLrtqw0QweA4PgUrl+Bui8u5DKnyVWoR6da6wRiaVMDD31
KnFN7XFbRhhL6S+4Zoc/uTRib6UFtR/7ZrtfiZ67QM+ZSj31cB7u15HXYcUlAAdm
j7t0rMnbpp616CcrrYu0tgc8ny6ZmwWVArRLk5rdApHRTBhzbZ62ftaspn4plnTW
aVdGauiK+gGrxW8jUoFlkvaWTxQ+mg2IijvnSp+BQn/T6dawSgJlFxmn/7vVHIos
mca8YAPDoHULUc/6VIizIauxUtKe032mEwCQ9Fq67UQffqaLpfJXOa1rI6CmKSBu
gTeaxOAX0qfgmFb/t1Vk/JGcQxfcoFGw+Ir5ksT3AvvbkOeIIQusckA/j/tzpMFB
hjylaaFHdeOm5U6MAtbIRdz4f3aRwZOCClhtXqSpABlpfSo0c9ACgzV7dm0QPlGo
C3YFzZgHE/a0Dk3uMzozgBwy0UZRc4ORUGtXlD3eAmdd78vC80LETZMPGp/UqH9z
Ue5qf3+XQocPXVK3b08TnUxAu7dgqWj8na6rpNwHrDhmsoPd/owotahsyEqaZ4Uq
nSMZsffsAV72/DGQTfUUvGSce4tD3C1M0fAN1JmJiMb+0odby4vLOI1aQPEje7s1
szhREhVIOn4ErAI7QTl86tZqVuAFbdBr0I6WbalOZWj+SAPyOfAtqxtrhCY0W0+L
I2dQxgiamMMTr2lCWj5B7/+j2H+uHgBSVpbYCnJHVISTF6cXlULdm/KPRumEQ0UX
p/WPYWinAqkjMUx3qvbb3Tagqrz17mOHwrvzW4UmnZ5y4KJJDuEd3XYWB8btVHt7
R8+EcBWoQxlzC/S6bCHa/KyY9hEz1OLteP30ib23X0dk9YvFNv6SHkCf11UDMaod
8Xon2tbfl4T+2iTTuGUhOpXD0s3FLxdwROMZvGiILQ7oU9VOvl93THst/k6bY656
5vRWLip4cnGQpZpy9NlvqxbWYeZaFdmrOBfvEGEQ5eFSWTgD6ygm+y5p3hdCilYq
qRCarpKKQrewoZn7dCI/SBeen3kKRRX/csQMuPCX9SNH2WxoI2pNrh56r/QgLbYF
XYcKDOENdSS/CHRnTvDK+op0VfxWMomG3iTP+jbuqRuvHs3DBPyd7ZN2Pl/KBq0T
oJ1j1krKO7vmTdN1jFP3qeqFZv/WWWUbR86/pt8VDt/tVJDAbHUXjc2W+T1UPdiG
OGoCfqzAVhiufxRJ0WJqsdRasdUVegjGd5d8yrEk1bjFZcVTXEAqT9kaVqzwt49B
C9gLUnnTLEX27HCtZoI2tfDfdwQtNqAIU5uH5JXHgEHMxWzzCERuCeBnjAi2Ms70
lDIMl6DJnjw78lDsjjqLkLXKUcsVUo3xREWBYsSGI3o6pBedQvwIbbGRv4x91KuO
mIeeGLN6vCWyuxZKy+4QaTROctWGJzZxScAzpMZ9XrCruFwbTCY+SbND99IjqGqr
2kfNWfvqPb4+ZAMkRj5V9xrpdlhnkAFrUjd/Rd8csIAGB4QEheVy6gxIjpahqmQc
Sagstv31UYo84YibegxC7g==
`protect END_PROTECTED
