`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N4XQnldPpJTtC8Txtaaq1OjRyqncrD9lnAZr+vDtStxvmU1MB5jzTtgG7hpF3+al
1KeQK1ow3Ebwmz7LyoXVByYjIP05SPzY6az5aoU5sKh6zPfEBrEhaYnm+++p3o+A
gt1kMhZ7Tp8u7PoHsm9fJ+sdsokAN4afyiONNyMJRHkmyval3ZvXaXeWLcA/y74X
CyRNkWXrRJWo0cJUP70PSCgCWM5qXx1AoskDM2bZ4apU2NVHwa4DjqC/Yiml1hs2
UzlpMcK/VQchRq8fWuR112Pov1omlNr5LL6R4XMdqJRndBW2NeDwwfuuhnE13JIA
dbU0GAz9tZhumObYYkzKmdhHfvO0tyTJFbWx60AoDJcoLPkahuJ7HlpLgvVp6nNw
nuxWqxoHQWyKXVBUcUuNZFALDGatuQBiUe0iboho0mM9LmRG4EzjEWE8zO6tPsCD
EwDDozh+UVHn0op3+kePNrjR5tYJXA7o6hiDwHcjsqmsrutcu1dIYki4TcPPeYEP
YoCPjZW0E15EpNnckHWFJJ/Sd4PbIpBVX4O2FtrAyu2MlmHkCebhKM2xRTP6A5vQ
74VAyKBYbO3TtMCF7tmqWiPKlyoISqdPmTzd1tXyNr+iBa7kuMQmPr9ZWmAl6pGx
d1A/KENoTmxeKZfeCIOGEA==
`protect END_PROTECTED
