`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jJbEMcz7cA4qTftjWcH+O2RGrtN01//bHdMFpaaRguaIod3Q5UVHsMlxmiRe9E6n
H5k2VM5R67Is8CKxU2HARBR56iR1mnNSE7VpHi7QydsSI/+sn6Gi+Ej9+5wpZoie
TJ8kl60pR316ll85vRJU8Zf1DcGyX2SZMEEKJKggvNC/ZD302fFkBIhR3LhK2wXv
TayhBSfYthinPq7PX6IxUpQSnK8AH5N+ilxTfnbSE8mzADcFDLdZn58iiHq4Ef8j
b79x+Rb1rfIEfGj11AMiLl4xt8k8NI12UFJAsU8aJvWCTjWQGrE/jekaGirL8yC1
VetlLFA59KYfqY8qzlumo6uDuFHFJn4UVh3wpiZAQoWxS2YFI1XGqJK+csZmXKQr
wzgeIR3IxT7GkWJSbKuNyTU9Rw6Z/nhyCOzp5tWqW1UInUgJwjwGegLYRJ+UFXb6
nCQ5F0SV3bwru1FNDtYjL7P4UAN/SCb+2CegvNLSqteGoTswVDsLwOZ1ssXcbxvj
HDpEsbrR5+kRK8KSfsOupbMm0/8eULZthvBekOUvo31qcROugECPzLypSXbMIohc
TnmHdDhcegrU+C6fc1dzlO3P00gw5lrqgh3CXNRenrVhiHI0bX0FmN8bYvCQb0vA
vwN/gbKmqMQgYQpLiMJWBBljeZ504HzEUxUQliiyOIlGbslbIDOk+HLzBsXmN6m9
GLe0zoP0bgWgUqCu6nLm22gtDq1e4OxtXAJS24ATjEQNf94xMzIzsajwLar9x9ws
q7F0JNQZWfPJFaqNixqOoupLkxVnbwR870Ggtm9RksCSLa8J13LEOEu09rAX86XD
D6xyLLsbk9vmVaazlLoAESjiUFiJ+InvMkwmUeJIt1ilBadV1gCExF1uWLI+c/EW
kgHe+GyAjdoqF6RNGd8vELysfDWn5fb778hxzN2A5uPMNxYDi0DenUkKpiuQ5kSU
ktRgeZIodxX9RxPCVdBKunhTWHepIWBZKN+kLkH+PjDSgYBD00XIH07jwXxU1tNP
CSHL9yDxj8O8+M/M+p8kh+nsv7Jj/WC6Bh90egPRiDC1KmdKVUEpsfszAwhdRc2f
cHZ94iwWJPh6fYwPXwrOgJVJejloYt3SqIXeD41PeVLrTY/A2q2T1B3UKJqJpg98
V2lk32gn7EK7c1LDrTj9kszMqihht8kvTZ6nv+AZAIMcqM/Mc/NCn6WZuo2C//5c
9HB/gmRnX2b5St8oTMzHfA+QioTW6VNqLX/fE077CBE8CehT1EwxDeLvqbsJSjP1
FKZj2GKJ4/bbR5jSRNrJ2HvYLowbD+4qpu+SoBsMzsEaEonjMei7QOpPk5P9S49O
`protect END_PROTECTED
