`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0k0ZHeRWX/63/6KsaThkxLQqgC0siAFoyArnJchx/JYP2cLAU9kppk4dGVlTC+Xe
8LlYIRyQvToEnlxK2v6FoeaDIPGKbzZ68Pf/q9Ve5QU66J8emN1nNgai99tOYV0z
muoq3Uzdcx2BpXzTig4nBBWL/wvryl/qcpvm30CU+1pT0iTonR6CkGwQnAtcyXSf
76Fb0ZXWK0uhw1fA5bGMZ8Q+TLOrgMRtaVhiqKYk2yd6EWi7XgbYzPt6EKpHfT8m
xoBOIOgTm9oEYyvX7e8Ebw==
`protect END_PROTECTED
