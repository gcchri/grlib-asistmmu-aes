`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7BD6s4SBHS8yr+ergDpFdj1ApnGp78LJUWEyZFQ07gCUeSbsMiPqEYgv6WpMJ9Aw
lkcANDFmxgDBJrEc9i5La4LX0nHToTm6dNIP9YTKHisyoPJuMdyfv03z97uNUw1N
YCDg5lDKT+GEN5mcYs+LGfeTG6VmgVXuoo/1sPQoDMdCN2OnLgzQXIDPuHEj7pkQ
Rlbpdck/w1uyBZS2kV3sagky6WaBzkjbqZwTeJM3rnMioLGLAOhYCp3uAQPNMq+2
rWw5NiaNjNQzKx6mC/1OYxYaEY16o/VwkiKZbNIdN1iG6fevw4hD5dEOzJpuvwmp
cUPuXI/WPkUVyy/dxQX9HpaVJZCMwzwejZ3ylhTPBPLP8Xcuqzsev0UTT8W28ACl
QJPJSrQcQRpQ9WfFutZJwntB6aHocf0eKemQOcAC2YU=
`protect END_PROTECTED
