`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NJ5hu1YNaBBfDl6axe+2fFSikj+tlmsE8ACd8Sas2cFlUh3BtGfLqt2POtfcmifC
jsYadcj2N0lljXcc4BMXKy82yAbxZ9obPP1UjTT5iSJZoBsu9ywGqiwjlWBbWSut
h1ihKZHPtxp4NIqu+EGWCrDThkmsKmC8BaF1f5pTR2t2x11cZR5g4pbRAJbHZLMV
QH/LN/9UmHiRDCuFQK6tClfCMnPWt2ceg9+j2wBDSHs8+XGxkzHq1lVs8fqNs9zw
85/qFUq/NNF4YpoPkFBSF0Lk61vpJsJHS037567m9wuAdizWZPhTUz4YUyv6zVf0
W6kbHxn5XKQ8Dv5Eu1F22kcTDcJiIS8vBfTwpeu0o9ZrkKE3TiLH++/fNMpby3Xk
NfhNcCw4OFLPA3gXzE3CdvXW7/p5BN+YQ5iSBlFYLxQ=
`protect END_PROTECTED
