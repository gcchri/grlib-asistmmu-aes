`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6WZ8PCbpqPA0wibIRaU2XNpcFcf9SMfrw231V2S6t4X6SYYjg40k6F3Q+FHGrtVJ
0eezhKG34N+UEZVe8Qdm/RZJKCFTXkMdiPHLgigIMunJXguaYJ77H6y78nkKMJt2
LeBdlzTRn+ePx8H1YoCjhTN0ku5EiUaU8E+8X/xSM9XeVu+fdT85eukXpCP/jyVz
N+Fl+ExVail4aBVU7dO87SN+2jzwlni1Xr+HABd5J1K8UeSgU+JD08mRxliPAS+9
bgT2G90JcUekLqNG2tauf/HSuO+3x+qj7bgX7QU77Ye32svThd0fDeNpQ4pjljcE
xK0OCwWaE/MekoeFfmTZLrGs+gQF6ZgPMghmbN7lat+lliXgKXWLkimH0WWsDD34
LKbic8aCu94f+kGgMGlNA7A1+XvmagZup6UVsUgQWOMoAYHhobLWDCVxKdLTqBRp
rROAgU7BV/7x37JW0+oA8WF5hCBHhbQSMOOXQ7bt2EdvHpDOB9sI0Po5DFYB6cJ3
Y12k6eL6iw74D8udNFYfquJmzRy4EoLGIJquqlrhnjB2nCKIgjPABgsUG/izcoeB
e62kuFAjPSe3CNWZQW/xbNBi+ItlHYy8qCsLhYLAXuORLn8wjACwMWrvwhwprFDI
HDImzbliBZr4klS+poqLiUfn1arb97WzdDJYAMgah24frkiEwHvxr2I2j2eDNxLk
/XqP5/uBytCodIgMcf5Mwed2P2+q5ThF4E2sg+9mFCUq53M13XnGZ90TpXCAZAOD
zZ/35KHDzn1pphUJ5405hstQYhboFBl/LPfqz5Gj+q9VKUBfTpAcIWLVHRa7BR5f
c6ALhvKYpJzjVaInF0F8IW4oXxF8FDgHAjKa41Sb4XAJnbvgh2qjEdDjywvoyKS7
qw1PJ6GPy4ziw/WmtRpyW1YIiChmkXezrzR2feCllnyuZ0pLJGu8heZpXJDhS26d
0JMb8kNuiR9We6BesPgHDD/souuqtfGS73BrXGNweX21zNJ9l21WI50KNUaO4iUx
8whWFhnf6Ie//dNQHo/ao5elFRiZ9nQKFvU9nKeq5k/JeeA3jEPOVzSA7KTW1hll
pD+shanTl1OMb21ER3I4KfhL+GeAqcihOP/kbIweArOh65ooUzSV1+leGes2YwWB
mi6eLq/6yC+rN/DLlxwMj6AKPNbO2b3GakPQlYlj8TOWSQGnl3OJ2yT064DoCkIX
mb+sPeQg0wF8ax/eqVi7mD+Yaaw4bJSS9EXg4QigBKA5B3DxWTzv/lLB+m46XOzD
w7aJ4x01cey9DC6jU5x6i4y+fAdKv5Ze/sZicDinon6nOCDyod1P3XRdI7wJKR2C
GkAAnF+op+qYN70y4kLnvCMK/s2OIe7ee8UMZwBKvM+0uKWlUFhSx9PMq6Il9CxN
6v67ojSu+NOTuiKsE6NcalrwpxVxObl36cWMiRhPwivihy31WMjurEZbsBIuM1kU
5vjjF4gQZfjCfBGMrq7MH8O7oQBVRciTUCDXdjqvlQhAi/psmR4zHar+fYc7ZS+E
rOiwfJVWTNF6ZWITc0VIwllX1YGyAHsnzwNVEXM2Gpc7Vi9WosCeka9KCaP5WpdU
UikHzY29zNs4DyUV8TQiL7iXcDAwbGm+wQaI4Ji2/k4QrKRn52z3fzB9D1/PlJr6
JMgrmWGUCQ3c7h7xE27Qc5Sbp9aX6MNyqCRMKRLdjF/Hco74toz9mLPy7r7IgyAz
WVNEcyjhPYMSYxfVNEgkDp4Sp8sUf50xKjncM5uKvu+wivn28GKgxDZwViJbILb5
RoQsNbRwCIMv/Y8zq7QOinBeiwPRINitjajlKKO1uzN1CaCX4SLb6PihctoQUGoM
FIn1NGDkmlZ5xRBPhCUcsZCSQ/vkM6ke6f8odHTTT2jq7NjBOxVPY0taZWnRedxL
Rdr6AZB70+sT4ZVcKWTfYi+RHoC2zi4UVjeyVnZ8S5rTDhIL45ATvqY5uyIPZVJY
PX/AkCIvDFDJ10BycPnu0R0pM7oZ33ZzNZxeQKDuadJj/+7aPSDrZhIJGvBN/dVk
wIfQgSYktpH74Ab266Zn8ELUXK5CfZXdhP4YUook2cWecKKoVJ3LHkmZiflUNxt9
eNUkV+NQfPa9ChqNNS1+WkWzFPZGEUHONPCPndGhzRqQ7DXNQ0t4S/Anx/b3CSzB
WiyeXY6/DXPU+IFnqGvUtB3yTUFxw1W8est1Iqed3Dig7ufgcJSifBCDdqAWeLdX
DkGU/PX5XIGodnJhZ5/ZG4OHzqNANGSOI8WvkE5att4wQ9RlLJbD1kbxvXVnxOWC
JlhzLhFnYal0pQplRKO2awueGnFsdOLdKOmdbTP8ZdBxxw34tiBDRx0QX1r6kmgp
RaiK9zIch2CX9go4wlCPbX5R6lQIH3907aRATfv8rCxlWQLJfefkCCT9/miQpm4w
jXp+7v73cKUqv98sverFFxGdCzjTF36qRvCZS3aSqi3xa7FNs2Jzq+2IRgJ1s6No
6ZUZ/Y7ttQ4Un8jsTXRakZgVX5qkW/55EYYzUviOIbY=
`protect END_PROTECTED
