`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HOKQbKtxpmsLCrKH2edvcj6U7a2ucKq1ryNvm80IvtzrtZx3uTcIzQncm+Gm970w
2dov9orv3yoSP2M0LVRpUDpj8jJ1jscwT+eddaPIuPPAUpWiYapgF/p/OebdDBZw
DSv2VtsF9IO5geT7JHuO6bzW/pdJSBtmkX0HM7cvVNeZMYUvgaYrj2pqSOGZKzo4
lExR1v7xrLXU6hKzr+baGYTrNLfG2TBW0AZV/Zsf2afAcoPw1/frZQHQuX5GT1lw
hx/ROYf2Jf+hwcMRNF5ODQ==
`protect END_PROTECTED
