`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BtZNazbmf9rFaBnTJ3G5kCVnvcogEb8zcDpk/2L18aIXs02JJaash+WjNwK1qkNl
UkSsM4z3bc78hgqBFV/np7hEkp+MvJPjWWh6iSfcXe/L1HfDX74mf1/QGoEnoz8u
Y/XvxDpid6MGoNiUUHVpXP1AdzPvjaNhYSvXhwfFi6LM3efXoNixuGVxlUdwWvzJ
JpCwloNSgcrynBNDSE3Iaae7dSFi6DxnbBJVgHtP+ABoD90mc/zFTw3mvLhk4XtR
bxFD5HViKQURKSwbQ+osZo4oidQMdWv2z2Bmn+OErrNRKoPxAsB54YssK+2as/97
2w8yHUsbipby+u2Ry9/OdeX0/qCvtBYmBVTfCw9WTJz6ZzEYRGTUsxdqyQBP5rKF
kMcs1Mfzrmwi2ZhKKN8yUbFNCQ49Bs+Ivrp32et+TeEZGQTmvC3ZKXj4YtkXe4Ld
1JRYUff8W3HFjbWqqIqxE5p8hwLsokdZgXg9FQZky2BInE9ORV4ZooKIzRdXV/qI
EWsLih9xG+YdejgG6OOLabuO1rKDXdT/1fncF5OvH33L/mWOu6aKcmApddpyFdQx
eGt+N3t2UoHMjcA8aeYFdgi6CsE5zFxRBVYluGQOpmI6HEIQXoqwh3QwrKzD9Omi
1rPjJ2EeD1Hn8vK0DwdRbg+AiufkS2tox51A/syZgnl7hEd8v2IK8DXRGRzTkSVy
bSl7zWThpF+zmqT2M24lYS4jLEaCYY6J3ASOb2eMEbRwept++2J7nqBs8zzm5cFL
1M88Pp3E8QMkwYRiYFRHU8CVoYLLCYhULAtPggJHvk429LdS0KFE4s9DMjMiLoiK
aMp76y4Z8HuuSx14zvaxqjffjWDptxaYe0sTek+sZmyJ4B8KVQwzmC3qRJG+4TBP
+JR7YJ44O4l7gxyB8tB69mOOrYZFlrk6LLSBA9WlNa0taSs+BLU4GpxuZ0C2Kgza
dOh5fIzBVhk29FlFYKxuLs9dgueGtLYf52DjEI4wk3mf+JW4jO9F55bLctL0gm6f
/l17uaCo/bTcRQJeohvExMJaroG5ewtiFS9ca7BSyHrXrjb+/ukt8CZA9JatYdo5
hXFcxGB60fgbz2dt3qPodoBHN25ywVqhTLaHf5373GepiRLVzhamTpxjO8k7bAqx
798TKotX28XM8u+MM+xJNIQWaDWQSVI7XWAEluT6BxUp7AM12D3XyR2MAqTqncD9
GG0+mBjsGQQhh3nDGKy3HDvZtSGpCWBdVHUWJRw756K0csZTOV3xIJfYCscdszPW
8NjNenP6rZ0V+9XzrvIgxdlasEp9naLxBLBZQgdLFPGY7cPVH69//YNbkNjI8xH+
VlzZ7oI4fy8tZ9GOPlaKCljD7lGF4DmXV9DFTTkGas+Y4UvFcUY/xVOsEnZYLyAi
+6yU0SSxGF++fXhzujPn7TOA286W0ssF9cxt5/sLs7yWBG3u8wSdLE/SRNI9GUum
DVVOi4tZDPWuNiQoZZBMA7AjmSKTUIQ7lIzobvNw9kDXDoGaiVKr7PmH7fuUIN54
tkf5kcO9u+tFRw8e9cPU4G9pu46diywZCWqrjtlk7QERu0bXQBwAMcDgJtIDO/uE
XapnArf5G3UgGWQmwP+JUNqCpW1ypDUvsFUtO5wltXInaBYgAAYywhnzK5m6OAVv
N7nbR7nMtaVMzl5XDVmA6Kh1qMGTMu669cCq6BBS4Y8DBKa2WmXzBLnYpdKk2Iy/
h3hQGFAVwBeQhMHBj56nQj5bbyXo1eaoRks9aC0GOwo/ZHSJcDlYK/AJ0Q52Ju5w
MFAx+QhyMTgGT0q6B0Wkv/+TKsbKpDgTAurWWL66OslgG5VtETTKeJSPczYZe1db
d/BB7a7atqj62rdSVY5Uq4Q73g7oqnfWDu7MW4xhry51KranZ2HWdB3RWZIcMwB3
c8/3kRT0jT45BKF+NvSl6VbIhdvtTNlCKukvagX331/LDxdFhR8vT95YcX5X9iIA
vyaqSYRJQDiEyY+AqzYjU1xVeC4h9H+TMDpmnN84bSUnCuzI9FAM1geHx83kO+KP
ruviR2yJB7CKtH8zMbmJS+VdaGU51wqYIHVXraNHHH2niHaQqW7wfVSPUJpyqxmd
v8lH614OX/FLvFCv+dptsuHUPuY46rzNagm6VmaQmPZ6bPM9k+BwaGIZ63eU+pIq
k+gzdiWcUZ/b+/43tIdT77M37HiZJ30GhIfQIaNRL7QRffmNldvRAwk1aClI+SoO
gkkl92YP45xQYwo7tHOqAHthCfnWECw9OfhS9mCO6Ynng4Gi81tGLkZm1Evr/Vff
Hr1bekellWgJJz82DQH1RcxVvyn6L9qti305+EKsxyL+02g5rlIJFsIM+b19p8Yb
yNM9Z2Gke37uRsjarz+ahcdCw9RVQDMQR/xOlOveVCGGokkGLRJCfrNTY8ly76nJ
v3ucqHxKUpK7PP7Sfnpi6vnqTUl2RgTR0Z5xrFT9M/jmZ/+ugPB/baElPI9IN9bi
OIgY8/mbjstqJSSTeHVFV5MHGlrG/b30i3KcxtmdIiKTeDUS3BX/od6dtw1uH2WX
DPtg3jZbg2F8ae8d28smik//XKrvyq+jzoOrzQCY6MAxaWHD7sbe1+KDki32C8QI
403jFCWibIYWT8Q+7Aj0YK0UAFXDLH7xYIyZJje0UmtudBaptToe0nfqwO5A6KiC
PbXlGQBhrzCtmXItm2prUJyUhme/jHoGXP2ob/seqgGE0o9duThQygAYXkH0Pocr
XjEG2YwWksBuU5knsGUkn+LT43tIQYDyA46p1EEFccqneS1GrGSlVt68E92ZNuYo
z//CbEuUeaQ+k5SYl+CqgdDZ7heu99ojA1ptnxXx6g9ze4VzYo0zLk0qmgO1gX0T
M9FI7gUDFUB784B7T9jtWPV7Mri5goRmz989MrsZRyyrKiZHkA1haaq5/EGF38Af
R2t+EG11ILrdc/47zHyZNLj7cb8cHff8giXNm8XI9vBwa8agtuI9A0tE03tFS6Wm
TfrHe7C0+xHPJ2RMgG/cdyvbaRUk+XZv+C6sthaHMf1mo79It5KQszdUsHHMdzyX
Xrv95N+Yt18ZwY0/MjrRz/jZLcazOXye/q9xj7jYh/Kma/zYKHXpntvVtX4UxXEN
YqMGhieT5/5bxkh3Z152LXTX5tnQNTHmq02yy8LWzWkzIbUSUXa7YEYTa/NSDGxX
UgqUJsZBs5s7L0vpMCBFMcde0NrggHapWfpbwsAATrSS5123EXofv4lnE8pUxeAV
`protect END_PROTECTED
