`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EhO+NLPMTzL2MvKggD7mALz362s1Y22uFRyxLmP9T+x7z76xOFRUzzCKMo60/1+k
YdMfZ971fu6SE9dlgTtyXSaG9WnQOhHvngZ/X37al2XzN4Uzu9lhA6IfOkJmDkgX
+XYsQuOuckvJWYZd3EMpB8mg3w6cSjIk3PdudNo6848dyStT7pRjiuV8g7f71rXv
5fn9ERZst4lXP/McVhUjQHf6RYyJ3030dijLJf+DR++LSpi6c8venrV2pVKyy3FJ
UfhurCZc+MhB1ZuOUau4YIqqYby4fpGRfzdERQ3TSX12uKDfRSK0rEe5+7vvxCPa
BJSlJgw3dY97W9Edz9GostHErKmGgXaQsx3UCugsIPlG9to/2ksW4aqC+eBUNiyx
yhK+Af5zsbynvlvGkcXMASGxgd41AmGKhRORFNorKsR+tBiE+sCZ7oYGxFtrCtyW
8kxSj1OZBwjVB2Z0mkOAVnqEeGppwVJkXuxDcGwE/vm87TpdSe8pSSuEL4iV12T+
KsR7CXX7atyLBgyJosRWwz3WnyUqmtBxO8D8Ges+B68Cx+LcAjueUWakx0iGORCE
99sN+4gnN4PZG7myTS7CCCFgOKgdN9orYvMhrSSZgBm02GvCwlDwkej9UczhMFRy
i3Kon4tk3VYoFHVeVBLALA==
`protect END_PROTECTED
