`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4ZPYodvzV2dBFxa8g3FaXRDUBthp8091bj8aZZVqnQ44jx4UUr/j79QNfTEUlAc/
kph1hgSskd0Wh6P6nEi8BpoiQyw03caxszEOsiSYM0c0p6rFWQ9UmUpgkTuKWOzT
BSQuWq80KpOPCXLeoJXxaxv/B6QgIq47Q3kz/20wi8mJPm30kslqQxA7rj1dqSLr
ydgWNrOBhMeODhEhbviZ0kdQLWJqUh9Xpcj7FEIqILZT1V5Az4TDI4VMfvqMTR2b
DoKWVVciHAjTKVcd7I9KSsuRt8qxd+dvbqzYu5xNCS/6rvIALOx8OCx6Tg7ruZTg
ow4vNkWsKxHL5jsoGkyuF9cRcLSVU0SKGfwP7f1ZTrbVKUuU2H6e0dgYNFjer60y
+p8LAHjPc+hRc8dtrZAEkFEQZCIpLSVwsGHlzvnKBIqjov3MyoD2dmwCe/004+y3
WRA5x8e8lWv4JjNWdjuLWwZLkHoNBuuTgVpA8GDgckKldSuji2X3xvn1wsgQ54ff
Qh6vTchDCSxX4BFNa0vWjlUOutoFU7ESWl7jtXaH5ZbglgCWHO4vAP3YM9dn3No8
DglfZe1ugfZ+H502m7qXBobWFEcI1iL8jjeRDszrBNNAcKU2Gatt+JIdA5kgHBtE
wtToaXWE9FkNGShWjZYAOjPlo0usVg/ErcvVRCryf76nzoa1cgeNIl0b4E/CH+y2
cTZq5VyYAmpADb47zGzl5JGxjHqG10vDDtA3RJndz8NTKRJB2JUP3vEhn/d5vh7c
Y5Mrmme3bGH+yF+KXeSwCg==
`protect END_PROTECTED
