`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mBKVn9iPKslp5I0uzx8Vfm5UptH003jz5LVvzeSdQUGctL8JBYCV1vY9D8dVPtOa
6kfgweWdNsMLq28PBZCekzT19xS3nCoY1QMsk1xhleJSHg463rr4PxyJNdZyvFXv
ozSoBgx9RNKerAQIQv27OVmuLoflnnpe9krb9jKfTNcQGjI0y/0HPHOvCvKmXxZ4
3osDPmhaDr4C2gxFXMB0WhogQ6VMvUu0aWQQ3r2ioJ5xL5qKlafkJ2z41aubThes
3p9GVLlM0aR1hlG8JWf67dZnkCeLbzP5MEzrbAmpUmOIFNXJHs4NHd64dchKlHiY
qy4jElOmpG6DFdv3GNycepChHWPXrIz9E6xDD5KKURP1ORZ+67y8xLUZcEIzEn9O
ieU2/NzG15MWbsh+8mJnQFpLy3//lb0M6he5Zcwl16g=
`protect END_PROTECTED
