`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o/VNK2RiwuGgFTdxCX4HUm+Z9O8ROXaM86F+6i/onPjoPMihqzPjnVgxTWka4j7G
oNepFEArftq0KQ8xCkNwC0+aVi8VQWUzksHx6bJyT/oelmUdf1g6UXeA5t4hcgtt
BA2Jm1ILuj9U95nTma9tfcdjQlev2VissgS7DhanOzWt+pvOFx4wc2MXZR3rQVEf
cWNNyHZ/JRqRvWrwrgcsmtM/jYUbl7c6uNkGkxqU/3fygxFYcIFP7ejIjrd9PIhn
ZDE6j1aTiEKt0woMU6cBXR+ClnI8+0rYje47Nhe/R72XRG/rGxhAYPgj/bo9ewD8
eDYI84sVOG6B1vP9SSHNiASfrwQnY90SiachbuCwjfjRPodda89F0GhwznTK54Va
NegvzmbEwd9q8KzK3DEhn6lQBQIwkTdDkKC0Px0/sM3RggMOf6ATWHGd++aizvQo
`protect END_PROTECTED
