`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iDj75QZncANboRjMeqxKKvoOTqPq/Ar1mw/fuLGocNHdha8Elb0OZhDOqG5TWe74
9DqZi3ezLKFrBqHnkeONMqPZnWRRnT1bsORHDCU/G3cyzHPog/C1OwrfX7UbEfQw
As+YtBfeEdWmhn24pYXEgZei5OgWwK4y9rUXwETfbrNEQTesEzOHRuSXJbhg3Uqs
z1LLJL1VeyqGHaWZEoyeovZwl9mB9u/kZXUb4eSTdO6Ks2+otc0fZUY0L2Rm9Gvb
8oCnyv/P+xYPUJPcH3t73OnyB6b/3gZBaJrqJx+LHKE58Mc/1ADE8yzlvrcb9sqQ
s8S2paZ78lqxmCT02dReI2gj4y/LuY5IyZ+GF+lnHPEtgS/xnbSCBxynkiU14N4g
/Jzfgnb+ygbefCt4ZY3oljl336UuvlxDxvHfJL+NWUMsKpTUUYHI3UQ67+hMtStj
WJ7kKYaFJlIY80FSiRAS6lhFlR3exhj/yReer/ZgbS7nMpYiVZ/S4C3Va+8nXhrW
yfDL21G+kR9h8+8kOPAm/jnJAvPny18o9nBrkP7FZs7Uf0iebhFxkq5sE8k/OlrK
TllAJOLjIa1/AugVxYrfZOxlhxZoCx+iCizJ8CXlYYjx2Q3Do3WvofAz/YxJbplG
7FGe3YG7HZRqtYpZcYCW8bD+FZNB0gejqRNMEe1XXebGe1UWqq0lx/OuyX3+5imA
nT9zghbpgBpswTOfqrccNBYVsxA375xHCglLqV+NyAgkjeHMQ3TK6npzs7ERB6k2
UGJ/CoUC49xKgOyaq6uo5e/c+vrMSLCD+6DZyNUGBQUHU8yjFVn/KquK7oVI4SGX
5benlBCAhk3N2qGUHKfI4Q==
`protect END_PROTECTED
