`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L05QpzQiez+m7nb4n9pPyAsGXnxyGaNcfdmfAmb2awD5yyRP9HR8hflQscPAM53m
v5XPqd4T8sPQ2/DxXDDYL7eSSoSdg4LPrJ1gpAtXduuBzZF92G9ExlHLrpWrfcUq
tAoCFxu9fhYYw0KCFCHmt66tVJ4+lTD038UuoVv4KfrEBsnoxFi7TdvA0AETZHK8
xBDcOvvMJCqe/Uf/sjWVQPZd77iPAfljLULjjbD538q6np8ojZy6QGQNgzSEEPRV
6dE9mG6kh0R2KM2RTam35DU8vtGHYqacn6zXo5KYmqCbpKq4J/X8xWv4Oa9/2/pz
yrLCLA+HDoNDZo71Mf92ga+Kf1rIR6bwZc9jtmlmyFzN2185m0XThOR9mgzJngt4
JhoXljqigY9LHTZB8/u9MrNsJXjW3xhAF7s+gwQrjJUsA+hfNkb8NdHgJVfEX0y4
`protect END_PROTECTED
