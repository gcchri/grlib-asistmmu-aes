`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
16DrXvl6eOidTsacHWzaVMmRKpSQan/gCziF4UfJFcvtBhz9Vg/l+Xco9zL9qwN6
pbqYObbb6GqgsofDRg0EkUZKELTaQiktFscrFxePxXQMKsLAmzzKfqSSqKGktly0
vQw9KIhsofcM3r3TLgaPz9CJEbOc7YZlBqDoZ7JgdKVgEkNIAQhJQ39Lr8oFfwnL
5yB7HJxa/GDKPG5E9yFJqSdErH+TbYiqpdf+tZyEZcTsjpmUyGNAfXba0GGy2sSh
OnMWXPydQO2p1rbXn21WRK98seklbNspjMjdrXQqr6SyW6yY6H+wOhDFm7IukZxO
2a1eoHovETOARVeKoGMRCDaj7Jg1ba2Gpj35O0ec8h9TI9VHa2Z7mgqayWcgA77y
6d7XxwHl6w95NRRTH0HH86DZdLVvDTKE0G08ivVQ9DbNMSNlIdF7SkPxKIubkqzz
AyZEVQalsa756vsaTqajJ33zvcErmuEuOmaPGbAWIWhkbgsxXMs5TlkVb+AV0JbS
LSuhcHi5KDr4csQ3YJcRmwsFz1Oup84Bes3ZalH98LO+YUgOZ7GWDZX76mmjFzD0
cyllbWPLFxr67MJmnBToAVO6fC/28NkXNSjruXA/KLIiW1ucs1e/m1B0KIdtTOPc
LFCFyAmgj+mCwjnxyitgJEW1HHmWsAzTUz7TNLZnYbk2PpQXPhns4XHh3kb/MMQw
Jw29bx4DC2yf5nFZcvqmAVAsWGA7yBirO2Yctp17qKGuqTp8Uo6p2TnPWTpp96iH
s8kTdZGX+tK/spfTfkpPkKNQzEpnd8SdLZrnCelFMVunDf/aNW/IgqaDqW/UrTHX
ZB1rdNLPE6/fQ/7Ks7bPv62qyu4V0QDoXju3D6oqHHeExZZ5EU6/bRaVP0JwByuL
HniV1ZJs+CDOXT7F6fx+Y9I7adW9bSpdrvcrjst3mqg0KlUr6PIVR9su6ZB7Fim7
myuLo89Z6XY1B+c7TYDN292chIKui2Yc0km2ONsWOvOwwavuJ1OjlOfKKcVEtpxM
RqfkOMb0SNKP/dE91nS3/CVZyDE8AE2GT+gmfJO6Mr56BZbD+BiHaHn6gFyfi4/9
Jf9/i/jDShve5fBnVuyZJYFpqerMNExlu2/iUIjp0lrQ0juuxx7YxOhc4lkxT/Yi
gZ88GL7wbpFFK4byPvI/nm+mAeySp18Md2xCU/0lJvtYVJcrOsdmZl7eEffSnVVa
TP25heK95Ag6LwEOq403c7Ld7ms42tcrzQELjM6F+uRqBS5DC4fucXKiR9lKRuSn
cNkYnyE4cwyuak0tAoJ5SMaYRuiXugJIB3fmvUPBXBotVvZ2igckbAmSK46lX9rK
amYNgXknw5dJy2FgbHjtYzRp/yp33bQPBjqCw6Erf6Yaj4qPoenuvci6KznM67Yv
kjmJEjvqbcV1lhjwWnVu4g==
`protect END_PROTECTED
