`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oh5dn7jJ0GqYkTRrYyaicSPtcL9tOGXitwaiNDpienENoPtZ0THih6B1yr0cK27Y
SXmh188KcxaVtQ3eUJaZmYfZZcAzcpJbFgXih3c3UkYuB8rGxgEIrmBpqcUtEcLe
O3FIK2TOzEMh3HMQXY2gxAoHD+0wE3Sj8jKuiON8p8scj/3jZH10BO2OroDXvuZ0
a8DBp0DQeVKpGYI4ekm6w3X2JjeWSW2OfSNjiKd7j3hlvFbunMp/nU1zxFAD0T/4
PqmqsvhNGCdsfCEzMCSFvxVbfYFywFCJMJGglrS8MpzKRsuPgwnxBiaMiTgoZY6P
/5ESmpih3wKvJ2ekeuz6G+qL499k9VRL1pkS1t9X6zKaj9WobNSYofazMTPZk2ff
ahplJ3SutnoZaHjIt5gsJY3/nwR2qF4RbHY+2QoOEbC5WTjJThyFd04u5l/w3eU6
EpKu7pdbuELqLkKsJItFn6VkALcZw4gfTyLO03kiDBgvuj7ZhUFrC7LXlVDzBcIv
iaf4pYu6fEl48N4Hy24OMxk6tMSU9iToKueB/idb0du1ECGB2AoZJFDzPkWQaBo1
MLOL0T/KPXXxEOmPKiqOlpK3QQ2EBS8N98f5rAZ7oG+x8FQQzzcbYl1TYn+ZKEIb
PWfuSzKdgv14a4WRXeFwV7228lutiC5DmEsnC3xy0WpzKKmhAciRNu3kYOIAGcre
CB7k/10rirXDfaXiOC6qWlHo+C381yl1jKYzRde1RED78CCFj+VOAy/uLS2grfRk
FZKfjj/z2lqYJoQmBXDNJfPywjoIJaWuiW2u1bVZD6wK/tgyDSvLOP8Qk/38gA0P
fwpmTRGj7YfKkyJDI3NQX2x12nKqyPSEIxHMK8ItSDbgbizGAhPG/A7k30FZVbkE
EwlhSeNKuYqWrb8HRcz5suJGusx7fapmmWU6U4a+gA0=
`protect END_PROTECTED
