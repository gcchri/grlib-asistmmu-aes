`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kF8fwSJIL1oq6C37WizlICXMlKZ7AQD8jqYOq3AHwjU0D4+2rmFJVUrzOPI9gt7l
rh6b5vaZR62t+1GSB0WRVfiTkaV50JfgNxoPMYu9gwdGe41sLilInXW7g09yPWU7
Zlsspqrh3R3qGbrZheARKBRmXaFFD/b1hNB1d73PdjbxGhATvKkZcnu8FnjzeZlZ
bTlx6ReJiCkYr5ca00MDRULWCIuEiNR5PkM9bbT+af3Fft1UkHsRfwFUZ5C0AN9A
k+a6NqQZpi/i/GSmIFxozwJQzfNwtRs0KCT0AXv70bvxsFFGU71gRddbjX2y8qoo
OiNX2GNJNB6Qfn16qXW8OQ==
`protect END_PROTECTED
