`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+gEtU6Y675R7s4P992zux5n9mDe5ADgB9302LRuR59N1JgGfXHO8g7w01U+Hsit8
/VAXJcMBsT+dY3I+4E98a7etvQe5GFS4QBEJA0vmgjgCf19ejw2QqcHtadHucqiY
MnmNNS4hAxjaBMBqLjK0Xc6QrnoE02+RXI/5S2r9++DUlVfWXPHjxc0bOrsdjz90
kNnbTfL2sf0QUaco9gKeu/yoVoIk1D/TPsqU2NENHj6V9ApKdgrw42IrjIQMUc35
ChE21Qp25Do5jnZ5z5nUEW42jehD78dcD9IZtgR4r0lHuXEXYiIgR3R0y3sVUREr
aJZU2g4wGiT0J5YNDoG98O+/YU4y2T5Dg+Oe+xhph+zKsLxsBwv9wkqnsXL6kvAX
wMcruHCdw8OemOsBJezTEc3LbjPpkOVxSf+KWNRFMdGFnNFfn+RriSSzSsRQ/BBd
cBlxpcrFc7EI162ibLiShwclGYzWZNkXL6aQiXzCoyNblll3R0iO6veiQAO0C4PE
iidRhcj3mAxWPJQNnFBtGYpRaNE/phYn2wXp597QXmQpPXVbgvxu3GA8/cZfM2Q2
TIizgQSuN96/Ra/n1p7mSDWWDsJIh2ap14wzkkS05x7ABWoC+9foVMfx072acMa3
IpS4GUxHM8rg96PxwOK/7g==
`protect END_PROTECTED
