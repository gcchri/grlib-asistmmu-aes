`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gkpjsVLCa960+MCyCqSJMNkZwgdQYo5jrQtEqK27GPjhMTkrZtUXXsoCUP0RYTUJ
2acwoJWcuHJSgLyD5t9KUmjHjymPbj/eq2xeVfSiFo1h+nmxF7/ZhbL5hJ5a02jh
oPrVF9IeUnSDh5NwVMCx5e2w2ZmUMd7jHepi4KBIVPneNWHuYKeNXbL8WC4vRG34
bCb7dU7B//ITkm3xQa2BsbU+52GrOF8RqJTf1Oh8Chz+WqmgjGbn5lEiNBuD5okq
UplPXIHicpqnt8alx6BSAEOuA3k0VxJ8DYTxF2+dVrSGvvzQKutVhCwsepRwae7h
ZdFFyHVvEs8DH8vg/CsF79kPZCcNqIh+M91I7TF280l3MkeaeP3FoU//OXVTRKG+
yQIw0cjg8frRtmzfgSEmJjWDKy5r3ccprU/fRriCgzr9G43Y+yfXA7m0E4qbc4v/
+NUhQ7dRvbvzcnvAo9Oi1+EeadBOatYenFd/sV+PXy7gPbJUZyB/92+ITQPlL/23
`protect END_PROTECTED
