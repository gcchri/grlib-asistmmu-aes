`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SgKwUKT1SGbX7J0BZ+qYwSYrzFySMrieatnvuvWQYo4+9d1N/kRauhLZYgE2Rrjs
UnxPx1MwWLFtAE1yNSsXdqNK4zjUbpEwOgf1at7QeW6nxaabATA78O1m10LucSOz
KVaXXPvJTHxJy3fpNuxXsYPYJV5Q1CIqPVFjQPUGkQUnOgGFp5D1bWUjFUApkheO
idx2AqEg7IN8vvSAKJGqxUCmYZr2kX9vCM2ShTxfOCrqLbiCG2LFVRLDxT7OcS+x
J5+Tyy7YIjn4TCcCmy9pFuGOO692bZ/5yHXbJBPIFFq+4NRdENn3I3lNbFn1519A
azNDvvlfuNmnxCZ63ZjmogYYhhSDZj9B2lBFYBdbyfGp3j3tcgM03ipIL9QQVJDl
TRWHrEK5OIjJw1z4+4gi7cNhDyUs6vD/ZMqpqpgavpYLYpJ64wYIk/llUU+stRkO
BWziu+SyuFC1gVWQb0Po0yYz68F/8iUanskuOj9kN9jns3LzdWk74DMQeE4LXTSD
vx3BOp5A5JzTfQ8fev3aphmO5ZtrBHMh1dgniqafjQOWW8+9xTCdErUlzFCzkucW
hHSp2GLJyb16EqGnZmR6THo6C5owjXhDJErzWzQL50RtbWZlslu59e0y2tfyC7Jm
QtAdQfk16771gTEhOan4hWljYEpjeLDuEJwR8e8XVw3b1o+0FBDQ/vYhjOnJJZIa
x6KZBKzFli2TKMShqPoD4myxsJkXu9lJ+i5P9ObJUt19iUHNZiuCQJL7uIbk89qd
SqzAcIEXy0dkJfl+V9m5FA==
`protect END_PROTECTED
