`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0f2mXPQ3IYvnr8bI3ILYXIVpxYEvqR7P9CoEshtLd2e+znrlyc4yN14bvN/oPjRd
JjQG8p6OBtDKQbiqYkXsiDxicpDeVOV9aK8+jM6dvojabreNtsFyyg7/zhIzag46
lBkMMJeRGwHZd8WopMMS9I/kjpf8tFAnjb42oBrwGfkBanfDWqFkIfJXK6x/LFil
FJJ/ULSOT7pN+aRKsbT8TdTVO/T+0oKwVEh8AsOE/oEdaC5oDZMgVtHN/EqUUQtd
N5q4yqZoSwFhTKm/QaIkiuyn+FzlPQc+HuaRYnw97rnm5Si8HGkYgnGwl/ElCbih
kqIcXZiTjxIOuMiyTVaInW5Ilshjkmf9UIUULSQjVnoEgrNZNgso5S0KialDXCCy
FFhQpMIl8mahCS8MTCwBS0/pTSWgsqUV1vxoDKbLUMRMHqXrsT9v1ut75bV4vU/5
lWYNQ7eXoQfSrAQ+O8aKAZSaBVLTy4C92GTHYWse1oGe/TG+Lsf0sW1Dco1VgnlD
gBjkGWn7mXt+lDk6VZy+m+AJnkOXhPJ+0WLuVK/BzyOvZg4Adu3IGopNResPdqn5
x6Ro/oCaG1uGRLIiXusLLnIEq4jjYPu9rMnEFB9qaz+SuFsiq4NC9Tr6nqmHeT6Z
Oc1tOzfXYHcYmrCtsm8Mwyv0Fzyr1zFKF5PNB08x1pSJwByozwcVlQQZlr+oFTQ3
n3sj1Wbd+GopQBBiABBbnCvqPlRxs2HYe5f+f5/1EQY8vEWNt5YFfcQXmoD0/jOB
4FmaJMa6YDTTG5ZZCq9bjeRJU5G0pBdk29NayW/WPAP/j1vyjFltCSRrHLYK6O9U
UYsTFXjd6nAu0sxzR03M+zXRfycd59wSRoufDrBoYgXGsadUnsknTAxwK6acWtAT
kSd6IhSPXYhdFd5ktQ75S7LTF1hO9VuWdgIdClWxFDB5cslS21eSlHOGK/Vis2q5
rw63HSONYB4Ml4/bDDE/84+Vwo63GiDNfl22pEF8hSQEAo+IG0NbkIgy7Or4Wftg
jvCE1JI5z94qAHg8ImaG9mH8PZSBL/tSevXwW6ujgh/bGUK5IB3BCM5GWg5CEnOb
s+GS/xUYviS3zHwtgLkgYZ/KH3mPZ25/tqbjIncbW/OAC70qduQ7AgGK1lncdt5F
4XF17gZKQvfCOqPEJPO5UConCMBX0LRyTnDD3hb2+qJZ+AhVPkE7QRCMHTKsCzTA
kOaAAMuu4oiWgfUtkAj0fTIm/tqOutNqkCsTmKLb/GXwCQBDlulZgWHyTA9VoX+F
ILii4Y4JSb8vqh3/EweHhFZJ3PTPhU2Y2KYT+mX6Zvkt+rul3H1xJuCjuR9DjxNt
2cKe1uMLzyIP/U7JsmHOZ6A2H70AkEykSZAUvOiYxtPcBnz3Iflit8XufLCoqB1d
0v52x5HJemUFKVxOdgo4kuis5D1QD0JuHJXktwU4rts3Y3hcCHU0Mj5BbLbH4rou
iSXmjWVi5Tg09vxvrxEUhj65G1/oF7kPv5nPav6ImmUs+Tys7y2wq5FcyHSyNaxo
rIwOxwPWHVE1aa/pL0Z0qgGlN6sJQdF6+PcyLiT80f+nB5DUQqYOq9EPqkvrtW21
J9vmARnEEgZdQjsveRfulCb3ZPulZa1l0hQlYG/HYNqZQZKb/pCojyEbMXZ3rnF4
gXfGa5M3BEhF2w7ulCDexDcPzqfIjv+JDfTYNWYXOLxxYP6OwQKlfrtS7K6CSq/a
cK0oUqPZn8YnMYDWQ/XKxOI8xxfbbmt+84l9JcW4ybRYTogEZpyM48vZV0esLhgG
et/cuHPa2R3TRDxD8kmZqodSlbJz22xXUE5Df/tFQ6B51L31tTRfOAwOf0nRWYcU
z6/Y+JWFOVYjFn7GRwFrw2gWZQOyfF8Qbd2yLmYuqlybhCOa5P3Z1HkZ63FIwp38
JYDe6PU133nXz81EKSdJjA==
`protect END_PROTECTED
