`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iQGK1xN7ooqO2II3xeQMrym5MvmyDgsbZo4j3Ac/TnMuv8D5qjKncfKRRLxwpntR
HlV0H0Ms/mxYUagxoJqgg4NGaAS8hRvbG/nkssIqzgJ9PJsFbLcp/8FFee6jtmck
k0FRr8APvCQ/R3iyzjnuXDOu1909qMkDnPkZ7I7+057Abl0X5I/K3tQ+ecflXUqf
+h3NbaJpPyRNv1MuGIrJGSKMoCm5rYl1xWpI/vZ/xG+VYKczvjnWdGP5QWv+ZYP8
PHpXkzG+q9+w1fECljtbvTcLYH8bdAjnnm4QAD3kZmmk2fU/0LAFobGqC+KJQlCa
JBY0tqVXTYQuiemnobJlKpDpNfTpAFK4HK15dlZsnYEeHxCpYvpGQhsHbE/GmOpW
ISuGZKE1RbK7eJXbFtAAv2AnL9Pwb+2CgGHY8vwE+TzvNGaN5QqVaaGt4VuL6ot2
GOY8g54vM+WQ2UjlE5x7ZZ1c32aMaJ6Sh/6gFu89Q5X5FFPsWzUuxPOoO5n6ILpu
u+YyaIGlldiWvHAYOL+uUiYHjcu9gN/E269w4QxQvMz2dQRy3v0x/swhhVFQbYJ/
YB+wdW5D1q8HeU3aDWXgmbG99SpnO73R+ons47suI1QdMJvRsvBZ0dneex2qqUBL
yhqdTzbAAt8NJz1p4b2P8MVwx3gEcA1nKwiTfu6mIo62pFk1rWYBxB/9k5NS5Sbk
uqOOfSqpenkf3UAbiaQvm7sZJF/PQY2m84la69jpXyOe2aWDiKFY8FU37sH0i0em
1EbcmRp1aL2JGaS1aVF801n9c6Z2+eZPO5ztqh/QHkXOW0xW+zWPw8Nr1BtlL1AU
8g4S9feTHvLfD8roIN9aMw==
`protect END_PROTECTED
