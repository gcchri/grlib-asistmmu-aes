`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BRdUI8lCKKC32Kx6eY+2jg767lF09uptn1NxXE4N0x1lSrmxpytj+8CVvice35Uk
VQ3VI4jMc58cycpY2bH8JROvlkDD87CwXFKU1M8U4AqrtsDCsroORmvyznQklI/0
JbiGKW5Sy4V9HoZ9iTTO8X9KlEvUZH3/mnQsd9CrK7nMSmS5k7uZVSxjrdYAFoM3
Efi9r56F2IwZXIMS9QTACwH0K+9tjZDs1CtI4GaJ1eL4/TLPYKTVWsbxF2F11P03
VRLrirBSeJ7Zdsz9YQn+cY2P/LhyKI+i8Zptrtv4UyDRrCcy/WpSakBfRVw/ypEZ
llZ2d0O4dlafnGQAwyGAeaUTjyIHnUDqpbfsvGvvEdbV5H8orgt2AkIzbLTG0MKO
qukVknOhsTr49HlJzTUjEJsirUfP7AwvRRXQ9TrXdEFeNioAfdw+gFlsRsMGi5Cj
iPB+b1FWkFFEvuy5EV1XH22lY8yNtmQiUMhBU6byDCsA1KleczDle0jrtpwn4cAy
yAtryAvETHkdViOzz26/ADdnL+nFP76wqdz02EZFjksvY8F3iwu4shLqeZHVY88O
sNC/JfnY2t/BTjaQ78az7oKmAjDpCYA0nX8G8Ru6/L4Xg4n5ESljwiGREeWpYdbS
Bbv5Xv/ril2ouAfcddrKenGXQcC9qRvTj5c0jg0QMg6geslZU8kYkOEi6R4nmoNK
`protect END_PROTECTED
