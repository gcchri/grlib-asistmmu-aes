`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e/xuV4Apxq8uE1+fGfS/TWJ9TVllHzaFok8xrzl4WyCey0Z3ZFbkjPRpm1xdyOY7
JtahR+Bi6B4tEWl5qJWh+lLUG14yUx8QYbbUQSH/Tb+JsVo6aGCQ8N6f9XFr3Gou
/lHfDjzqyR0tuNS8lq7cfDdZHPnWFwKNWKYykhCpugGlpstePLKJZgr6aYyUQD4Z
+nKzijUMYQdBLEBb6mN8zaSO0CXAlFNH09CEnq/d1yTRRqjgkZ3mcHnuOL3sWY2e
/HFAm/HGPij8ryd0SxX+1CglyhCtEEFKgWSBT8I/S81FpGwzuAnwM+zR2e3ol3Fj
0wSWfYtfLgsoPp3C1xezf4ZTmyQLM1nxRPCr8Q10rm6MsEaXFa2BoF251m+h5UXz
wp1lta5FS4LQIKij2lwJO5BpPagG+k7E+AGqjPk3yI6kVYaKuearCadR+CcrH65Z
4/ZI5zxqfz0ZHLUobINRh9DWTZ2vTf2FXX6Z9aoJphBifrdNVIzey90hpI4sNIto
67rpZOd3NSgNsf+0KHuzNpdXhdMIfkr80Ir0fdc5cRSkxydK/Ch+CmDpdPiWwMvI
EbQXL7qGkOI8KertoBq8KtY0QNMxYjwrKaFP311HET+0bFxuqtYrd4Y0kYXRFvqR
rh6BUGwoqqs9+uGvOjzWvAOAs/pPBgyo4m4yBD0J6AQk5U5aM7LGPm8d5qX/iACL
xHn+mvbmcXoK9JB8nFf/WD8N4J4HAOLY7UAm1lVs6PY3P90hT+ua90duYEfaBNuY
ri76vAplFj16WwFStDKHMLJ3eWlzxyfo1Yzue/xngG7r7CLTV/ytGE9UNYKJYrrb
k58mSSDX6mT1d9Ha5JHF5ymFn9PPG4YPUTKfxWtgae4QiR2XrEUjteSrMYxmO0rc
IhzyObczEoSwe5Iz7ROtpV7nc+xGyTheOye/MpFt/IQPS+HM4rifeCrNjeoahVHR
ps6CfK+JFhCATrt4yUjXu3ldcup2eZ626zc6npFkL7Anym6fBoB7XZKVkGAidwQh
hNv5kCXLJiBv8W0Bma1PKtwiHpgOAobj9b3S0+RwKQvBWNlxsZ0trYTk7htG2xXu
mmuZZUrzrXcyNc7pQZvzlDdaLM/BNUl3qOO1FKCPR38tGWc0M6IaN6roThaAv10T
oz5pdMG1mBH3T1I+USoUI1T4P/l5NUJMfD1SVkVm6yclHfXgKSzbJueSJdupPbqo
nUzN1OwJwO0T60JKHy7qGRaeng5bI/UG64YRZ1RkwH/HprHy6KAFn5LMMkW0ozvk
2JLhn/gxAT5wVGsd0RY6cc9r9pE3sTbogq5ov2OGcOTy0e0maOdXsQGObIXOv1Di
2HAed90ARzL2nyu85WI4Ox0jiRdbl1mWV1C89up68B7VUmxlfj7XWUuVYIyB4PZ7
8WMn4WlsGl/ivjU+/dDaC8i/SrPSUlU7YIe6onKEw/c=
`protect END_PROTECTED
