`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UWVTEp6Rxcf/QNyQbdcLeKECPqlICzaRV7wYNVfJ5+rZSjZQDY63KgT6nZvSTYn0
9tv9oSpwRKoq98STrtyu9KNGOqLI7pxKivBZSQ4iPRY7D0XQOaLYS5qGK36D+e8V
+6I+47o9HLN57aRyxUx90ukcTiJ9N3Gx3xlJT9k0wGqTtw5KRpFwUMoqiob5rnWE
y9gOUiGNsYjlWHbFWFSbwBLcgGLylqDox7Vp1+1fHvt6wLiKRmqYB7eabcOkN2Sl
XNFcUFn1apBcm2f4A1wG21KzEiRrWv3X4Ch29aECOjFpc+r/fiWSGnCordMXdYs3
9XAOm/9JGJdI1iLi03MiwQX8kUy5uZHyKJw8OE5Gc8uTN0QVDciP/ZkjNJVOtTGG
tLDp2jiD5X3X597Yr7dEUQ==
`protect END_PROTECTED
