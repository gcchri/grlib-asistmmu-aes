`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8kTz2OTF2iR+zZ5gUFtObvZSWsVtFr1bHeEROcWCgLMmruJSN4k1t5Sfc6CBr0LF
LUZ9cO2+7gCW2hvlp3AyU5yTdjfXsgvEsEPr/egrZHrPsVd2etQvtWaHsHzPDuaK
peYMgNLtmawMY5pvNzGdxiAfOIMf4hbgCeniXwyZkLzZ1feYEgOC5MsuHU6ax9Jp
OXNKaiddPjGwMjRDanfWr2E8ShbtV1OuwLNjHL6S5epv0h6e4Bt9CPyLFP46yXS1
JRkwMQH09LJORL4KcWnym3B+Ww96zVf6J30uT6ot+NxGu0Rhv8pNu5O3NmKVOiwE
KtlsHsy54sG6aY2j/IMzWze5PYfbWqaT8HJgbqGurEDqfkfZ052I0LE7tvp4fPmi
VeUbGY0AEmenpEtlw8eGxpseoYWKmMs0DkNNmQ5sFeqfJyhpOI1z/+J6YL339qXV
2afPSLZ/bOGurKfrSvuGXh6pBf0x+VJx/M+kmNXibbt7Ain18H6PvSJ30PwhlL7I
`protect END_PROTECTED
