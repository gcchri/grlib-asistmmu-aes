`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IZmkQJL36zEkBAVGapgMZ7ktjiQ4puI/qnLojsMnhrzbsXE0H9d+zh7rYBuXjKjH
oZ5+BqJSYZVQZKL6vitCPs7yeVVMLdVrhMABr7b5fHJbCVCzUObP5bVEHuWUZfW9
yBxT7GYGjJBEvV6S066Lv2dbT2dTwk4lKQSIRdRoh3aUNRw7FWvl9tdpg3cL1Po5
ljkCjQj4aO6ET0uiZJX1Q1zds+vhTvSjUnOlOIQSa382qTwF+wG1FCzoJjlYngjq
m/w+ggvkeQlLRui930K9n3r7phnDR9uOf7I7HpmpaKBtbBanwBMQQur5H45ZiJNR
Bt94WPH4INpXW2p0fgmC7A==
`protect END_PROTECTED
