`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KimmtoJxH48eFs5VU8uBQDRzXYUlsgXA3dhRIWCa4QfhXXMWoYg3ZZSiC/XedOPo
3TNMfOMTJL/G9OwaMO26/2u9IQsWfVNn0hcui37HUBkIyKEnpr07mu3xiSIRXwQ9
TnpQtdlJIUAvYmuZ1I3vP35AJ6bXhU43YvNyelgNrrFes50HcLlfQDbPJvbPViTs
zdJIL9UtnRE8KLD5TtjIt4aabG8IXvLgQGN5upM08hcuFIkRg0t+ZkWvSKj0GOUS
0ZMQFriaS9xNXHGc+Wl/1JE4JryFVyLUOqLyO1gkL/jrKGAbyn4UTvrZg8debcWI
CDXQXE3D5iOwylMqLCv0MZ08wRCMk1Vy/LNGe0vjrwzDuHAV/0vUojBcZg9qG8Ip
IWse+6fIZ5/vP7QGKRLWtInB5lZO+sZCdfuAVCATZ6g0QMT+x3XYblRpJJu+HZ7i
b3NwmY8tDdGtWzw7kYCt2mKj9Y7xqPPnHiKznB5MRDs=
`protect END_PROTECTED
