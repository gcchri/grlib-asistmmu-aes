`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MmeTV0b+4AOP1F2cXP/McyJCtyy1JGNLYXkY2eW9ezOyEETEHS4lAoQwPa9xxdGn
0EMXSzuIj/m+AYYdk/1YS5WVLWRC483Pb9CT0flk3o1bigdsqtMG2l0jyia1RHfx
kbxcIkxUu3YUPIT/6GqHtJmnTePz6GnPwzYUAcDHiV1baKV7xNXK+QWN0sU5pac+
o5+f7bL24sGij+5AAk6/TiYCRaHHO/w1Y3clZMjN2touPBiUe2wdjLSrTU2HyTaM
j312pVxryktfkV7t35TxOInGmapovLJ5Wx1fpdiSi+m2EfMDlrLHvBSJW5pCVwlu
lf3wh+AUCk+i8Y9EbecGx7hgYOXYS3vQs+dAf3w46eFPJrM2KiYZAKjZ52EHcWPm
mmIxVk5JU++zOg77CHFHIcSBLK2teI9SpOWK/vTegtxmeKDidWhPa88degFSe4LR
sDEsTHfmQ+52F4PI70qr/lTMDAc0h8K+rFAtzZyVqVU4JiKYV3EuzHPArkPR9OiR
caDCV/aa0DrHWQpFPN9SxEYXZmzPmznVBswjQdyPIbioYqPJi66cuFjZMv3+iCQK
qfowzWvg8ulQN3AqcKKtgQOT4BeaGGUDgBJprW3nFpM=
`protect END_PROTECTED
