`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gdXukDdMCStSzd2AW6LDEXGSICfWRtxLbe5IKD/6/ucklWjxJSwDFNvJJWyWL62T
iGME+sZImBwtkstG5K2ar4x3rZ2FBZG3gy4QmQ8GSvaxECKAaoFVlIh1d6PY/7tN
aP73TlUrlnso74j9HSdp4ZpIb59DOx3uYnFyTJMvebbeujubzxESq7BBQArPy/qv
3RX1GYundcDevkqCLomp1JARrTa48+zTPCMPv9a3fHZkzQ6/S26X7pDUgA9hnAYA
NyK8tuoGwzHuDDJQRxnGJWcHHGfQgf/cl9NZsi8XIINoYRDe0mtEwZmJjJx3aUv4
uNsMBfKn1EmnExbMLOirIw==
`protect END_PROTECTED
