`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GdGOqORWIrhq4YvW/020DbtNz4CiJChRjYX26bFbZY8yglcYy8cwKXscqycdjvy9
uk/X2voqnRww+NWiMe44LKnxmDR3+sjKI564acMogJwzLtEju5KN1qtNw1tqtqmm
gBra7A3yJcDqaoL4v857ceUfQfkXR3oIbnQtzh1UOcrQ/Kpt67WMKkd3MbtGb3lO
7E8jrzCCLgig5aHY5fLLMwYXtxM0KykNvtMmvksUqfnASe9wTXhKp8stNGrYTZpI
Z3h1E+lgQ4qSlJRiCl3RFZiSidX1aO9tBi1rSVwLv7DXlUtX+DUvPvhGJpX5moui
BK+u+w2osTv/7y3HzHLseYEokI1/owZWpQdIsreUED7SLh11dAzNOqFsyAaxDiHx
VRNSbLStHupibZ7cA00LH4BsUJ9rVkSGDeV5SyYZyKFyXXMNp12ZxejV88XMuOUg
`protect END_PROTECTED
