`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A5ymsYQxqBEX7OBEWpR7Dq+kZ+eZVQgL0I3+XY1WmJY9ifTx7DZwAtkTX2i+YJ9M
eI7PoLgkwpDSWZ5qqgoUj0+38A25ihHbZGSdP4hZxMysG1L85TKMqZ6z+MQvvZMy
93JRdizQcu5kONKzqXhDaKGgVNdewz3Dn3LVF7aZfO5yp80EbSlHQr6MBQoOWUO/
wQo7cDUeoXg+OF9rQ5GCERbxT2gQmmsd5cwUPn+I/+VvHnguVfG4eTrbgWvvBI+a
E18Tks+y+WMtARZLUPGG5K585W+7l/WA1pjshknjtzykt6LeYjKzk4V3ekyTyQSD
dwm5ahMPV72GNAtEtOfus5TlVgxX5B92skGzbjw9dBS3daejqdoe1ZL8hNobOMRd
y+UiyYN2djZuppOEviKIGIsBMqfRnx9mlNT6P5qmpiVW2IidVZ4id7yV5FJptZHm
VSGC3aZ62bEBpl3X26O3blSpjwfWrenj3K+G9a+U86QTMxpsYf7XPiBrP6FQEl4e
4IEeAWQYPg9jubArFixZLS2kD89bEu1M9NEhpFsR5S7YnTPBpqXjUw1WBXgkQFiE
VKwdCuviLIFo8d8wbdEpCvVfLAnpXXRxePgiyhxmf1CevPoCoGxyNFk8Uvr1IrIX
en0t/8+xAD7XIUYzRr+T9Y+uOh9fwb6+LMKfcceDdigF+P8fk+nxLSpuASHVv+bS
QD8qApy7MJ4/Gj/7vhHiiQRuNHqMuFmDPDtVq6tA7wjiPnmyBG39iAiefAxYSJy6
XWdH5Pl2XzkGp0lwvAiSva89m3pgjDIiNJ/4uxCaE6wUaQQ79JeYFDQ5K3cdZ45C
KDN3E2OnepdMeoHYTYsHp1w29zGmv17f7rhIw9R2V1Kfa39+lBwF7NMVSgf8uuNX
RyUqSSHV8n5gCgpN+9zwtdD2eVbgot1CanGLgW6VQTj3E+Ld7DwYXpv1TvH9VwGN
Dq9aVmsy/6z+kgGWvZdQiMzqxsinl8Z4c4c5h5hIe7BH9g6gmI9MK+V+Rf2PCRmU
cFvH2sJCsQcbEzumHTAXC1q+jZf+YhKhOj0Y1bheP9MYH3I7uwluXR3TtbSt3nM5
Fm9aLgpt1hGffx/G7ZWJ2LkdbVoJvLYuPgL69+7RtbAg+7lJibqaQ0vizyXNCkTL
HFe7BgXC+pas85oFSUfNZhmnD1K6c1knfkD93rVS0J47VzM4fCY1b0AD6wI1U2+s
MKOEASvJsl5mIiPCntnKzeN9w9MFMxgzCFbZ9BMtkYRTtLIrtJFQ5mM8rDl6sVOu
KQxUizPOPe6/SYk/5bfVdWpN33TdrXprTNTPddNMz+KOtOnGGekdWR+tPxC/OAYt
jkryXRXM7oby4tjknN0/RYC8OynSZBACe2lWbTdjRAdIAwpo10IqFcDkoqaG1I89
iB+70vA72duCfuZ9Ss339d2wiiv78FHY64M2OTwyqxbof4cMVzBVEqbmjv3eWQyQ
CjlVUB1kMfs+yff2BbpoHz8lebEORy+xcsXJxS5AOlCh3NnFR3R60IwUR/AjpDxc
sBfbWWtg7OFqAi/WHDrP0Ee2JdIYvupOP5A4HDtdO8A=
`protect END_PROTECTED
