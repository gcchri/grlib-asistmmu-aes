`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O3byame+UEYyYWcBBp8Zzze6vHvVgd/xG8gBvamFmxgDPQ2XlG/aedyW4Kt21y+T
CeKtRbSBBlhi0erBuiUH2rORvOVQwWf85P8w4Kn2c+c6bBwg1uR8lTkzWYyj7KSz
mhmbSky4H5FKxW8MGH/pyeRAre+t686rV/tbqRpMiuFS80/Jzw8kIoJrxDIAd0O+
+AjFecKo7/kAXJD9IQGLvSs1TZUw9nThMEMwnqXAxDJ3KbzAqW7D56fg/ycHUiOU
ZEbwjWN6YaeFxL+9qZ/V9ujR9vgZesx+WSlAdQeU19Zd/F4SQhMUxFOSMNcsZWoQ
cQfGtzRcvBpepckWVj8ErJbkvjWEewlb2s4T108oV/WQFofUOdvMAdjxp3xSXB4H
zOr9ah4keHBSxAxN1nGeK69Iw6SDwW1yigaZsgdpcddCmVRkJxl/FjolA8Xl02Wl
tvLztKvUii51Tycu5gwXC7IOt3K5o7l3vHNFuEkomN3OFc34DdyKycDbTqzbtprW
W05iZMvJpbQprLnhnEf/USUM9ekZRZ17yi599/IuyPk=
`protect END_PROTECTED
