`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Zqsxj8SQ69Y6W/HJGlF8wqLeDDAExe0NuKPtODUuNAi9bwdRcy9w3c66L61E1j2
Vsbe0EALZJkdVxdO9XNiYV0xEZ5QD5npX8qXV1MU9xz2dSDvWRMogIXslaoRWU71
gL01Zpq7/I7r+QlFhNZDDw/Vsa2rny1Trkf4FMQDZcEpSQqxZNonbmRWnQfDWoSO
Yz/djxbPh9yjwa8pUiAKJQ5utjQC1x9hTWv+nD7bZrMxfVQlr0yJ2dFgHcThWHwk
taPeHjiUZAmIQ7Oj4Lh4yePq6h1Ws4FGIxS3SlTN9T9queQopW3DMUEmJJySHJg1
7wAT75ckyyFNvzfWGToeMZdkvnn5H3u4W3IlGQxARVvngbgnTXt6lssANuulGWra
4CbgO93Km0sABqRdylJCU4P3OjfwP2cciXL9CEkqjDLufldd/2tE79HqHFXkOPj8
eH5WcYYbyIOpU1qf++biDx2GmkFSWy05wxXRCU/+T8E29XR9rDLqTzuSuvg4eXkB
Q3edYG7uoPp/GYCzScBZuiy4wm43ByoeDDJ8JTKJON1NOG+n3FpULC51ucF7Es+j
tAGmxwaG1Cw6Uj4oWTQP75C0vrWqrlTDoybvLJDR72AbNq9GwCPScXYUOAaVecop
FidiqxjTiCNSHTzPS1Vlsw==
`protect END_PROTECTED
