`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2zRt6CBKSDfx1+Qmc4momVg2CmVyqKOWEQhdUsOG9Ch428bsdnZwXLSjEZ9uEvbN
FQJMRxDjb4RofGFkUTKfaHhQoWULcOUl9STo9sgx2Xb2k8/PiIqSkOxa5aRATZUP
nLjRvpDYoEu0BQlaHEiLIPSib0n+l5KqyUCaL7YdjX8ptmD1ZzjsPYqPaEPV+FJM
xwbZkVRjcmpZ2mvgykZkVNm3B/zyzG+oFgGnzJmbPHxhrMOadupnK58C1tdG56Gk
yw8RL37A1yLAfe+GLhAB6jKl6Awaq3im6FqELTKrNEjCIQArg4ceKDwQtfLCXEA4
2Gt2B3prbOo2OOe2NmHVQljKswkTCAlW4j++0ptv+czeTU+3OjOsBCuMKlRtetaT
lO1mAio7vKwNBssKLKcpslc+59mH9wupyV4S5791ciciW3HGR1bCVkYginkvr3CF
CBI4RvY2RZYaysSpEuLF+9zXn1MeTEz2JrNx7pw8ze9RHi6zwfQOaRgp23cS1sJ3
Hw7xGFHqMS3YxU3H1C7jJZWAQwPXsC1kjyApvrqbsFCL4LV88vebvf0E6oGTj1JQ
/BjRcqvlDP5wMRLKkXxpfh43GLTovgfEVFF3NqOkK4GjLMuyXiz/6tBUC+HwUHKx
x/fpqg/9gj+1S1cyUtPu8rNH3NTJrE8TP1KjaL4a2MPiP8JH1rEoUm+nd59MZ4Bh
m23S7he82EEGBk3un0Jdi9GAgx9JBnJd/LecOY5C5/ndxayXXW3GSLahyxRaDKqI
jj/srnSOb9nvXq35k6A5cQYul/R1cr7qoxgWWZdX1jF2uIGaVo01Ew5WlXbcmPsJ
0FKC+Kdj8DIvH46netdEIa+FG0dNum/0wEFW9PdqYGB0MpsAQ8lJiWiHX6M3l1dj
6i9amTJ3COVhkkRMb/mn+A==
`protect END_PROTECTED
