`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0uYYp33BKu/+BSWAN83/yn9mogQKOF5oJcj99d34nMzJVOerj1rR38vPRzB2GCBp
mg/z7PoCicDapJd+yRF2YfErSNkdUBAFI91tuTIeLJMjw6htSh1q/48fCfYpGAu3
ivzEYru+YY3JK+NZh7h0PctOa9ma1v3+mjUMFiUTXX3scjme6EEZ8SoWWeAqZY5t
BPFJkPc3z3MqFARFe9tei5XkteI+N8S0yhJBzVn8Mq0lwbdOvFWYhUJQ6YRry3k6
tMk7VTe/pf9DjQQlZU/I5sfyZ5biOAbpImTcOOppAaJHosmOGlUzxjBtquUnPygc
GUQeE7SV1r9QUe6XXlCE6m0f7Nh/PkpCmkOq10nEuv1hZz0zA7ZdIWGMSp/5iIBG
oZ5vbSZxcIFnh8Vbc9fXtA==
`protect END_PROTECTED
