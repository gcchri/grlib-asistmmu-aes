`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A/efKg8te54clvY7d8yyzE6txLfzB7ktwzMkyJ0O1rXgd4sBfoNAs5isSklYwQm+
Mvfk4WDDXLrbzJxgYr7pZJ+NNvZyFVvve0DXEaHKCPrM6Fi7Q48KhBMDBQ1lfnd4
94SVc+cUSv3IdTN02gejDQ2QTr88Ce61RzvTl8AuXa9wyEEKBQmTb5GvibqFbC0F
VnKjmtdF5kgLDW72cFNrUtZdeTT3rFGmMMzgHhooAsYR/TQIWHcFGG0XrvVp0m30
t7V5w3TYjdOzx9GqSvAfikFW14xiVUASZL69LT3hnhZIv841Ri6oDBUql9G9HGg+
aI0g7iEhkLE2zOFCCWUlIugs9GKR2z6Ia3Z6uw5924l2OEGtbkRoTNxEYsxLs4/k
Cqho3/TV8/k/lRhKbsIlxQHOga+oSUzTS2KLftTJJAObgsdwOuBCXzWey4Hmi/Vw
ku0gp8cdWB6ql9Tc8MBLZMpG+3RLKu7UmbaToznhPgAhCzU34aD0jFMMtO0etbFm
43JTMCEUr3d8rdsze/+Xa/nIUCy9ehUSf6Vb4wl9A1xF4LLX7Rc7vsT68Cbv6EX2
OgjjX/PnApRO/sh5JKcPFcn9YYHxtmvUUNkjISN8fPkPsmWN0K4izD0/DyC0CCQe
Xg/nBusSjUafAZ4+T1Qy9adfh7ClCo289WDblGL92ogQFkg7iabx3ZakLIXlrJkD
CLE1kLBglZZnROCnIymp4VFVMkfONN+IyVbPADJZiK59AzWaZ1h6ytXKnpt4svpf
EJvEsw8QrqEMdIUqKUueJKvEGVopCtxxhiYJ3oif2o8FbMzG7DY/nrdiQ6ISwNW6
akhlGzijht0n0y1MdTAS/0sBnhtDg0IrP4/ZXY+IOyFlNcjSnbwxP5veSYkos3RH
dHW1S+B6mcK0kkDcNiSq6PlshFtlhV0/R6XPBvP0VY7JLfnXRrl4DaeKL4jBh2jg
`protect END_PROTECTED
