`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Mlb5+av1MVsZWWC7/d4h0nAEYAa6+xJk40kBy9JEH8u/VeSIAVGVdUccIZxKXuv
IS+JgPuRCw0Nq6RFYf/knWO/O2lLrGL0Td49EAfD0BhtNPlKprn4y8lVMnnO1R33
3qDyhkqohXulAF8vMxIMiLxOYSJfmwxaOSxlgZpTwAH0ddALo9UN6gZ5cZ/aYL/e
JRx7h0A902zyG1ibhGf2ghDSt2E/9EK5s6aSqKyWq8XG4ru0yvLxg6xUGurWDa0h
cH2Lx39dTR5B4I2+4c87cSN3kjgS/Q8VXU5V2xkXZ7/thGq7fKrTVxyx80xV3pL+
NYLZ4zOtOKmNXsYZcLi1C6OSZM3v3MbkOluRxSaLLtel0+7CYjLLUGGJR0UCo3mL
4vsF4iYZ456ytRdOCzFxBByayYQ/tbLLOL65kguvr5+VTkv/H77aoU4+X1khjUQC
`protect END_PROTECTED
