`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ph45epVifBC+QU/KTRSfjD1DjFSHbZ5Fp9IZ4iEY2qEUvg9xEprMU0wQllNYTU4m
67oaClsRiXDHyH1GWeaEUXG5P4XvBA6KYfXwoYfP6QG3Aar93hsqdqg4ejeXyEHu
BgVrH1fWxoocpCoWO7/j/cFKW9H5k2QI+AOglZMrMHKVDtY+04Vu6veBUEZz/1RC
fPG/OE//sZ0ea5+OUIWGDJWGjU1GlYKaDIap2OmWJvDEzISqBfp4V7iAbY24W48P
icsCwsAvM4qeA/TKrRLusY9ZSdnI5uiyXUvZ4FHdRb1LmHkM82dhksZgWJtLATEu
Vv3Nldno981Grq8Iq17JaBQLhXOYC2lX7Ze1LLQkJGKl9cTtzNOZxDfLyCFhOjtx
igSESFwsSUwPn/KCxNUtiAG6OWFbtZREAeHIizcWr/wFOSU4Y79ZTxdeSkv02I4r
He3Ikvg6V7cuTzTwCmTrmAHuNd4YctXjM/9YM4uqr76W/nfVBPHU2ZsdEdzxnfUR
0zLpBQseL9j86Vnh9a8KkuwMvGBu7Bf92sjNw3LrkTGPDubSESj8i1Pxe9omCxGZ
30evkaVaka3KSFIVFnjncepnQ8KkP98eQZ6eqdJqeoWsyJo6HmZEK0GyB6jUlMz5
LvVFLiYcazPHb5NJni/Gz3LLQ3NR4S6eJ0xQN6VX+fAYXDoC9LnSY3u7UqewzoOJ
3ibnuA7defATX3fmtU2TkhEWz8TR2iSGAJ7Q3nRM2o8+r5/EIfatZGQ+/AdJOifS
VPWuILW/kmkcc/4j38GcjQw7gecy5jVwgE/ONWrP+E3gLlcI7gFUTdfvN9UCNR5q
BnQ+nvBW68cnfU9nXQ70J3IV4byVoeLYbIvqpMnWuRW/pG04yK6njm8Gi/LgjB3T
Y88jwcHH8bicuwIoxroZoQ6qPakH5R96ze7SL0jeC1lr32Q8jX9KrHH2LtTMu+zh
69+M06vgqkYVlrZDT9Bop+KEgev7f7VDyY7dSmOJ3grPiLRARIRaIIKMPfgp631R
9VSo9Z+pN2/CIqwTp95HF4aba5qPzDnl22F/5yO5lXeywUINKB13mlWS1JlbLGHq
4d2mqc7OW/8fTPDaJ9vY7gMBxZVjlKqcjhBVulldBO3VUkQwDhHGyZqDgq4CgLQl
n3HM5EF0k/xKE/SrP+b5W7Owga11Jjf8HZECkvrCiRYb/8m0Hcjwpg7U4zpIJlZV
CMjntP45hH3gqB6WLLACJnOjvmI6iT8/TwKou/D5M6/cPMKZ4o3+v8sr/wbWop25
DK1ixRHYQcjsI15dFcvRbri2ffoqAPIexPlZ97h5MZC5xC83EPpGFnSH171LVGTB
3af1KMLYg509Jh38bvO0OUbTUipgMcA3A4cXcyLMQwHQsQtzG+VrjU7wG8Op2c2u
93UXFUnkKzk8SHszcujf5AqDsN1yH8B4wVQXoimeJHp2USpVC54u03GRfj2XK9Cb
50pw25w/d/5MYDT2ndZMjoF7Y+7q8+sS4pmwP6nQ8qdkJ5oAxy1w2iA9UitJSUTO
`protect END_PROTECTED
