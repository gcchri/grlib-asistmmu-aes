`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gi3+Wne3hf2M/GikDaMIcq/bQyjBOAXgAJ871F1CXe4bBh1A2AnotJIgCV/2A1UB
tKvlqfFfuTjc1HcU7QCazrWgV5qMpXvSu0R7ZiVS389YcBlNldDaVLH56BhQuKCW
LSsKNVY3eSiQZHno2tizIEexzIxYa7TB2CLxwMvYbufX1F/wPgXgCnvHdHHp6yVm
QYtVLqCfTKVyYsJiKhvWSyJSzZ3OVADOF7dGsfIsEL5IeQ7HskRoT6OlvRucGBXJ
/JmBzd4hVRwHHthSog8IFU36rrXadfXNl50E68l5y6an3mjx6jqzIJ/xGZ2T+04x
K4jyke8MfrCv65CNt8P+JvuMVu+dTq0UznN4MwsbmyNDP9r9LZA4cr1/oeDMYJT0
/DmCYsK39DsDqPa4Ins2RAIi29/KywxwxdEGPbbMBuYkpn0f47qG+1LvdxKV/fvg
45hbEFbOPSl4JZFvvKnV+Exwmqt0niVXMDW1I0gajM0g+4hfKZ1xuR21zHMycyKU
`protect END_PROTECTED
