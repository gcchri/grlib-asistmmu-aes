`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dKjw5tnq42rah4hiNhkhna9WkGFgcmIEVLWLzLIGZSeVMz4ET3UtWSlocUl5XyR2
yANbi2+9vlXmZ4TgXU/c0TTK2uDytu+P3WfLr/v3i5LS5fSVgE+FcIQFxX3LxwNW
GmawKGo3KhfI8G+8x0qPP3TlGbdNi7N9L6ObRgByn2ev+c5xyj1T19XI4AFlbwEP
GykGti5zWFdq0dBJv+tOo5sDhatj5Ioty+sPkeOkJZ3SACh7rnTBV4eiC7U4CGoa
+UQB9X3TcNs1HswWM0ah0ATs0War5LZCmLheegAhlq0A/+BzYfco2JRvlcu9RHEs
/HloDvh5s3rxHGPyQvQA+UdePIeCQJqpnBChtX6cMR00CdNplI/GQFYEWEbihs8X
TTw3TMXMBGEzu8kJSnZ5cchfEm1aJk2wLt2D+DiF0kW9/EGjYaMO8jD4rYywc94L
+5y9ixYY+OToR1FhltSM/BnooB+g5TbKRLE2PSWMTcQIgU5EWzmi5lZG8xBztwHm
ywbIY/KZpU6Es5cUG1MMVA/+pXOQNBnqLSLdO33u0E+sNn1qHwJtUrf2zEXsy6SO
IgPoC2pCZHcZWZZdoLSGGQ==
`protect END_PROTECTED
