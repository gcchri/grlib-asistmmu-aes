`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9cxC7RchlucGv62kiFq5h2D0e0gbDwpLVdR3gDNmvgwLL4u9qb6Yf/+9UQhLXf9q
XFxZnOd2UTs8iWNRod7ksQVSBj1MWDdXv0T66L4a4inkV0erUImFnLb+e+SfAKOy
XVxc56TL/6KEyeVHA6AntO8P5jQhRnwY8vD5mkYdVrYkAxnpAib9yAm026lilhF5
0pZrcBk4a1sHyasQ9s7VInA0s+lCSTf9udwWzCpRxzDex1o6HIi72vGBWLqWWlRU
UsAjusFsnoponSe+JTXQ8dK/yjkjlvRPySy7s9kwoEawZxQm/K1ZUc0HUQwZD6l0
HkJ/Q/IbO0hsub8vDaMReEgAmmEFg9LH7UCTvp3ihEfOy8h42OzjmgQnvOqCzvIN
`protect END_PROTECTED
