`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TxzMbRy+VLQ1mR0o8FimcswlgKbjuSJQnm960caL11Cv1hHkaGyhfWWJNcCQWmf4
2dw+gdiaNf7tD9mCmoq8YkrdTyeAqS9D6zrxcSV5Cqmlqstkykr3Z+DRDXddg8/S
16IqNC1XyRe/cZlNJebHumveLek+ajqG5rtKM8sXnRMx2y1ekDQONCLJrTYoFkbU
kne2kiCYHaWymaAV34qaXTFySbmehnnwEDua6yypaNcj11EUQwL/jAY9XzHT8mx9
pBvkVTMPW5PrCMGWnuFmJ7d+m/b/NqpSAz6i2dL7lciweyeNY2OSBvnW5STVjY2H
p389kcV+U5Cjtt+uJSQ+vQQg6cE/Pjqm88i7eUCxB2jVNe/cqk+kwtpqODwsrOuj
SEWQWltLxkeShi/Fei1X9rGL6qtznEAfU4A3T+1+IpraXKdbiS2EW3ntakNi1lcP
iX/bICVZ1F8ANnnUA2sV23e7it+HAWW0UP9FIV9L7944ndYOT5AJjYZObQpo76kY
gcEpQhSViFS4yRAvlQSerivzirk2D46mkiSoZJ+FP6B4Xbj/raq9VpLBcAfMYPul
f86lPl7QeLF9gITOL4cau3qncy4DhRYYT4vKIy2AMpOCQV6OZVOCNGEJfvPA2VBO
6WV6ZH1Qb8d2JNwhY9u5Yy23ejSVvriBLymKkrWHx1oZr5eBFIWAX0lv/9ZEW6/d
fqmSRayCxTL2r0MRy7TcNvUC1SIizrQC0qCqfKQYPZYxnkuYVh6384J8VtJYJmW0
EYuIJ8R1iq46Hf7jD8XlgL01VzYLGpWEzOmisP0+V+toFajjYBWB0tOYScCzPDdB
o+fUaMdK/xs074c0bcYnBknPq8nrb4nukOD+bc21QN7CuaotfUMwmNue+X66FCY7
7drlAO+kEDiAVFhaiz/MfeR3qtSdqjd5vb1DXWDaOOMqXlF3lJHjDAsddPbcEgD/
bUEYG7/UpGUAjCaQgtK0+39eOlBTRkvXpRVN+71fqawJmHrVXlj9TDmy7xubegCK
nr5vUpa40iFqwNH1rn9F2FHyy0I3MRRTxuNQ7dbJgxi2QMpUVPa/2lnh53nn9Fwy
wp80Ij2QrwMJ/LD5QEOwdOS7FgJeoaCGKeIdlnlfp2HemEcz/8AwkGlKCg+Q4WQ2
cJrnQ8PtFDzV1aJwZG5b+QTZ9jCp9qGUFbkk8BIUwQmryL7bhtgBNqsWEnDmKwsQ
iq+bDlDq/rOtJxcGQ/Il651n9HFy3uM5Izc3+inGEd/vlkF84OfMM5d0bnyhF7DB
sa+qkRD3+UyIRuWn4ZVIo6ZN8PutnkJoMuZBBQ326pa6lk3H9g6adOo12n+NMIRO
Q8o9m3pbXc5eztu4fAj5qO4Y3QyON8keERbs40QeBW1Qf6L164zCCPZtnGm8Ci2f
zOJdRi9fYhEU0taFLe6fEU4LaOyj4NV92ez0bRONnv/F8RbmlJP+QxaG9htGDr81
ltf0LvSGgF8yE94sYYL4p4heMw01FWrwaQf0/M2pci0+ucQX2GfENQbZlh3YBDnD
3OUs3fKeyG5BhEzGEmXhqXh0vEXU2Ii2+V90rF+QRJSX/Yb6SH8J7oEMyoDpABFy
/Ihz0aOC/YU+BvbWFLTl8CdCZALvsmksUrQd6wlHcuJ1LOU08BaifUG/1kzitZxd
hJt8Q53JUjEkvNInoHHVTO2YCCbbNZ2nHVIJFeFIy1VnoJV3wHN7IAOyeVLEuZJo
ons3zW2/ZvGucdcdDWLixtKZB8J5XaWvR395lrJ3UP40x89pirkVhKP6lbZan3jF
LAFLVprN0q74Q+UJ2FGbK+jOJEveruHuqTTdDCOGANo1u18Ie5D1NteBL+twa1ma
KI7FxBdZMbWMWcSAWmWi8bCvcfN81M8vjN9P/BiAihS9gUHbH+35z+WN4f3fVtwa
sy45wKfcRcXEEsXWueSHR0E+GArL0g3BF2CyJsOU2oPDOndD07i97Zo09ViFcdYr
YqAnWa3b+0zgpRvIICJmq0Phu8yg7moXGEncHlYgeD5QLG3hMJKSp65wUlUCvpOT
Fn8b0p5iv8p35TNsUufmAciPmLwq7lHMFGEbYMe+qq2NbfDI1V8vJ5JZz+N1oLum
UYm0oxYt1xOlJ830sHzmdbA42ROPxY9ZPRs3q7fY1KVog8Vc8JYP/hEl7cv4cFbe
y4XMxZ+u4sTAMigyykJX62Ohn+4PTo93NC+Gm3h8xOhTOjnwOnMTWwnRlHrZfSj+
Bg5mHJbQ2wLpw11TAW1iw4JelrvTXvZHbt4jmih8/HthTsq0ZDsUKruYrvR+n3Qa
dIMWX7hwp6JMlkSXim8sLAYhMCFNfGGhWeVtq4Kdys232FiaONddi/+kKtfYKg3M
BnD8RCJjsDWdrWVbNHRUqjmcsAJcDmFFIrqW2bXzsGcVxy7QEQpD1RwPDjJGb3Q1
pYEJ7nN2KOZFvJSKcR1oWkgH3iKZsyIBxrfeFT36xRHwPLDTm826QjkyLJX6FkCN
bvAq/ZRYmx0e/AouZMmPzho3aKhqZDU5WoyRtpaIe9yHSaZirdoWwdAnnNq3mnzr
FIBSmH002g3/WeiucJOBI1nGfqOuOZ2BjjZ+7+4j4iJgY7NP88VUCl+qtr6ki20m
OaYAYz21pM9AzWrGZdIkLlYaQnSnH+mjtTV07vP+hlAQ/u7uaLxKWFrWZ8hMme6B
ui26KHZDBsQ3THnc81rgAfowJQ7oGrg+cxgsw4P3i+RtiGfxoKBbkIDeV4j8iWBz
i2opqu1zjN/v89zKHRRlKgB7QXxxieyEL9xphe7fvu3v+1TUTRLUaAgxfTh0z01B
RKioxWIt6a/4ZB0AaurAYoeNfe4iwdE9HNeUd2ugXzGKmNKU7y107G+nMJIiT2Ee
7yq0nn9wzNoDxGQVfwsnK+Md9jL5d3suEkkDaW9S8kyfdOKByCuZkBjuJac5DUbY
U/G/p4WRc2mZgMJOYjwLt0I0eaklK2lt7E3LnXAfI5YAQJWd3Rcd0qko/FIND1h5
JzJ67GoNRysKuhJAsBFvXDeTCG6ME+e9owmuGRSv3FKMHw2e5Q9fWsA97mkElp88
2rSkkIPKji3NQJUShReHzvFYMBeNjuUI6UWPcmhoh0/mLlkRT+OVWEmqkGNV3Zzk
ioIHtFBX0OjiodotuNPHEFWTofUTx1uDM1PkHYxRkpTzD2Xp0PnH4eRNMR9LNPZj
yhAw/3ZadgBp9skvyemBRqsiSUJBSs8X9SJktQpeL1GBt3WSbV3lXzi9aiELhNjW
tUBIQKGomGAataoST/DCLz1pqnDJ+DeKxMpVIas0lEUqC04F7FaZrGuS6yznUnpO
oXfYmV+UIFrf28PPDv4q9CgxlRDEv7K7i2WsMVZ57QulbpmXKzbPPGHviQckSpLd
ZTVJzRlZZQSMVFo+AQPfDk+1G+QPnCSBkG6/fwOmr4kxEtxuV7XsW4/k/CBlsIlX
mMm+MkMlvy80aB/pl5ii1HglV2BdMoxcQXgk5iKspPQG6PMKOz6cvEFJ+b13Xutc
o6UPBH/byi2vYU1L4tewV0Gd5lJy/UaHQSUborUQcWojOjAT3WvN207fi61onDV5
t9xB2sJ6+3AdAbwappW2beFRLpEpO9QGfMrpPUrZf6mmnUSWiwVtEyLJ3Fr0scaI
7vSo2RnMntQ8PfkgfeFtc83HSIuf8gDnYh1MXuc310N+b4g1upye9cdV3uO92eTL
wJc+Ei8YjM9S5hl2tQfJTQt5+CEItrREr2502I1HP7LBzMgykB2tNF8gMdSvAh6I
NZdWDjFA0NM2kl3Tlu4oVUbTFYCmjSbruDxMUd3huu1L99/5x9MqAsBVmsX0zjtF
rRRnp22N3diOyGEVxygzX8frZ1ZfrIG2LwGaInVbAygLeCU2fc5tKQSSyZD8+b+y
eUBbpW8XHk15lEHDeTByhVNQs2t8//MntV4POQlsw6mLO0l29jnIQMdINFZd5Ucf
nzxS3IgS+clpPKB6OdGDdyzqKLQ3MWzBjv5256YYBSLNz0aKnLPgvkU8trytmJgK
WE/1SygtilHqSI3Ie3PBOcRvYCAGhvfuvuhASx3lM87M74Uj38Z6qGsr5SOopPDS
gUYi2vWmYVgu6uL+37rHXRTTmQ2CijFdAxedCrgEJ+Z3CkRDVbthQDjJrMOsU/ZE
rTPSS/4Nk6xGBa/niS9VdWWy29lIoZnq9yAwHhqrtyqRxogVpyOhKqWhzMNj0kNu
vvT4/Y/FbYrLOcH2xd7H4sC89IUmA2kwnrOowtYhfO/Ljzsiwqoc/uVdT6T4OVOH
LkbO2ElvhAh9AG0ZovfO9DKoLH8NPGnl2JjnuW0RHMgaQqnYE3T6Gs+rUxa7BTci
g3mOhZQkC6IzPPqwfZDoCMB9Wb0x24Ecxpd7vgJac7wOLFb+69Q4Tx2TNMx1zDa2
S3LNqwflmIEYpVkAujfiapmYmjVunjU9kYGtWc7ikEB+3tcqfBEwvkwLoGaMLWko
I0jEbnIfrdKw+c8xH08u9N5/So22VvpVLQiuxcxGfwr/7BhbbqQw7pX53lU4EVj8
ORJp11T4c4k2CwTIBO2PvgvDZlMeP7edprkKAydZUIe5UxBjTJvHA6ObPaId17gU
WDTtVsm5KE+XEFS3GPAql3WezP0hgCcODOihK8nCw7hePpTzdXZ+QE9CmnPOl6OG
EuYDbxs5uRB1qsZMO6n1G0hCfRfDwvl8KT3CWNjAYzoosW4XqbI+kIFy60q2x51s
/8Kgy/oMMX669iaLxUcT7i5BAkEZSj3E16ByUk2Cg9DOD1opGeAQQJLBiy8lnXQD
oaKZT+MaiorRQ+vuz1v9PtrxdebEv+9tvklkXWL4087Np5fMxSCxA/+L0a6legdQ
RWINjESSeeys6RxoJZgvonArTFVKjTEXz6xHdwp8Oy1tuK+sKcOjoX4Op3F/EoqI
/vpp3woVkAApOug/iofbJUtZ52h8Aq+XbmZn85P/gOc8CkyBZNCBa+U1MhwQiW3x
pdcjJ0nwvWm2w6ND8Z9Q8rUr3kgED4IsBqpUJfFclSLkVzy9WjJH+G1TfsHUGzfe
Xs3NERMBxfRLZvwJZwKoSNoY6JTh7OqL6RKsoNw+TDaUgEwcPI1MEWikOsPGawAq
eBei4tCF9ithQx3ZyejYuDvxIWJkNCM+PACFE39tsgnqzz+CKc+4r8eWiZWYF4rh
kQtMbColFqtnv6/kVl0iWW2yjqsUvleHXR9uJWnNNwgA5tqKI8upfQw8ajvhU9yr
4Ggathd3GOgRvhNXYFnZlyYfITDau6YMi0LQoewyWZclMeDQ+41pXY9wqPAE8eTJ
xx9PvOmfSUB6SHz7+Gu49g3ampNuoL0wK6f/ZuSp4GcFz/4iDiehWK3YSUIVgmAp
tiVgLFZIjThRtVn29gANn4kNe8QbPcHaJy+tA1h/kZEhOVM/3bIe9iK4syJ8Btx3
17E6Kwdp7lEgE2KB3dXmjwEyhOG2PuJggPRhtKuU/MK1eUViWG0ekjXK56PBcOm+
iqgtPfuZgxOdnICzCxnYmCAPREV4gcv5x+W6dTwI0+emraU6dhcsvIIQTghq06Mc
Zc2FU2X495Mz1XP8JpwZnvJCoNQaY18mp03YEp93RSUWU2VZ9LPIbLyA03Htlg9X
VgUIEj27Z3qHvaaRNMA+3fVdr7gjqy87xuOklgUFTovkW/wCEXQfynVWVN/CyumJ
uWattxLaut4fkvpmckDCf165AEl+OcQhGOuE6UuseaTMziAUkr1Ns9dlbbdYEam+
58hgWa5ydZbygWM6YpLEeQ8t87p7HLrbO0io6qaL6S84RW6kiYzus/EWnk3NFyX7
yN/I8o5TpNFL9l0n51QUEfGo5BtoNG+nNJdhjK4l6cc507vFZz/DtM/mz8bZNZUk
3Z2gOV1ZYlUnutyha/FBH89M/+oFlSBSObhxPP25IrEZGWD3ZieYX7rLb1i06z1c
VfVl8ANHwGz++WijJRc7HgWgzeIQnVc5xKMhxb6cG/sTUbdM0yngnEMjIPq4YHsI
l2pKt7r7Xdk96zYKKJ09nUMBUjlES/Dq9iCmDVtSEEcvzkocGIN9VuvsfupAI2hR
kVVBkqV9UYu3wSeWvQ2+nmB8U5xbZ/6zAUaKIcIGT/cleCYaftUnSDX6dUmoGjrU
gftJdEJRpuVgwlTbejH+ZyMbabO7I9DKHQNBufOVYUfYXiL5lXVI+S0eYg418nzu
P/z+8jHxQ5ge9LYl70X7lOwKP/VOs87MKuNw4k59vajdIdz2Wo1WxoEVLXnh67d3
WtAFye8iH2HPw8tOXEUnrYOoLkO2qXA8wIBXLEeXkzIumqrqQYDiu09URE4yeYO7
QnwQjGsUOIXin3cmzT8YQDjo5AXx3sKliaS8TUwySjNHycyZWMapCt2TUoQec5A1
g+Nik9ILvtrxyqR/5Bb/fo/T3Do26/kKIFSRv4URdvSRHfmGDn22Sad45Ry+5HxS
+u9Quq9tTxVW97Tt+gbVLC9fHW/j4tp5lPhpberfPeu9QzSxo3y3pPif6Kd4YIsg
DXIYTxg8qv8PC67NE+iQlGHWjl5H5g50sqqy98Zpxq32y12ndCHjGVacQDIIUc1t
xuKXRJXcvrLmjHIu5WhLx+OlveIinTgJo+AP3GjymMiRwp1IW2ExRXkKxd7NbQH7
KMgtJE4mIzRhK50SCioy3roWtmJ5aFy7MJEUE/+UwTrSzN77koa5kxF5sEXk/NbZ
SuKOwX7bjWXYh/PPMIbK7FUTr+OWIh6XUT6I0OxLi+T8whFVXdRKRugEvwA2YzUJ
P7AuUWRE0T7yuYc+T5McYFJWWG9/BwKP1rI9D2jtk5v9W/UEtuVzAdh6IpEyOPxX
qzSBEF5cx6gm4WQar9GEiKIlKduGhHAtq2eIovdA+nX3LP+0OiGn2193U6UjFhj/
QwZPHhXSKgND7mvimD234pjDtMdZTXAphQd3RiF4BAqSYkNp3tYMv9Jai8RDQ0ir
alKGWgXywUM73d70lNEzC69K202IxT7ZKMmZrIhCFfqtVJ9Rbuy6Ov8flkfnTVr0
rDNDRcM+X/TpX9uPNcEzmZ8MMJVNhoPvNgfeoj57ird7RwPnfmXZSLJcmCcIm7aP
0Tu+iqGWPNzhHLqSqW06d42AhgNYS6sb9RmuONOoimP87cY/Jol/aZhpKMY5lbRa
PbGw2/PZ53GFT934PsrH+tj8c+z3lxj7zZZgLtwsGBEVNCPDXFJ78Gw0t9HnQAMh
FISG/ui6FuXTz6P/XtbG2DKnRjirRj70KjoyBREk4pKj9ruaJfGUFFn8BDbQpNHh
qZ18AeQsEn6pG8wbPXPzwsuM51luxDCeX/QkC94zPQjLIFRJrVjHK+oYyIhsoiN0
bbLIcG9dQzWem6dg4NFsW3ZORqA3E5CjFyf8y5H50T2+x3LAPX0mZ9iNDX26JDi/
sfh7erziUa3ViaGMZooPzNsxc0nBhHweyb/l1M3gpBpWF7W/7K2u2al/rfAm6tM/
ux1Uul3TdL+CphqQFPZotPFRLOicLwyzErieW/VW8ZgpxtPmDm+gSPiT53zzJzDh
S/sMDyE13GNkc/Mn8fJ2x4LEKTjhf0wxwht4Rk2Ni0tCJ7rJxPkK4ZmCMbjryv+g
GwrzBQV9DUYURYM3DvtqSTlvLf5mawafk39QgV6WsPnwYRYthw4L7iOOgd11Xxlk
24oNkveObQST6c2K1vZkR0ibMffDlCUa06codcTWETiM7vqWczG+xoo8XyvNKUfk
Zf4rggBIsrT8I764Y6S2YaXqTWyoTqm/ZZ3kBE+csi+cHJ42nCH56NNrDeppjTDD
lEkFIWM8OThs/9wO5T5dNMO64ljG5nqRuV/AfG0PL0ZvgrKTzLMlfjTum8v8nNuJ
CU3QGrovf7+VNgU0AOnr7C20sLs3HY3YdvhGKFkt4RsCRRc8Hw2iaGi/ZiM89oBb
L/PjLYt4vB23IhkMfHOeJoQNA9BZvufzadGHEDCCINPORS8eQ6oXfMPfLiKdEg5z
/EIXduDn9oSmxykc0QMlSBniezklbincWeRLmuC5aOHuAXw19yWma7wncJLwtNXA
XnKdT08eIDvt1di+3t60nYf23AtzqlZ8pVzkOlL7YxZoESIKLQuXVCii7iimN9u6
/mHhochnzRV8Uom7g7VdHVHroo3CZOQxOiQH5eWw63WtNFGoToaxkZzsG6VMjqkf
ASPZj/P2k2OqaH/BfYwra3wsvumcqb71lti+kcMBs0lDVT/Xutlb1pabWkbk6HLL
vyj24Ph1s3KOaJFMS20/mf2SQpT6jVLy68EDXNHPnAbn/P6WYUV/wrDfhiC+JqdF
kWnrqokQe+0oi3wg0BY4cOpq8s3ZCthtKENWx91Xu6kd7mykl1qlFqhDw7NK9VeE
UF1W14/4w3QXnW8b8nxHI6P76grzdJLwT4ezuoZ5EoEZAGMvE4K2kjgCqg00jKP4
ydQBD1Tzo64ZEAt4len5f/c7NJXZghmsC1Je/muVuUJKu9Kpl4YDBxYCOXZl93Lh
P38X/CYJfmtRTlTnlAYzLqouH94YUBReTJ9AFaA9DeEMhc5QPLPT2etuoJb4hS1p
LzIU9IGPbl5QGHDjWKmgC1xZ5JTIMXGiOO9uU/T6QuMfaIbhQgifw+kdZwVb1Bm2
U+kWApYovjooFFJvURGzerHD1AI2QmeSFto7hdZ09vNYx10INP3dH92PAzXwUWam
sJ2FC9GbOLbDNFMVRFHeE007Sk/cCZEC8Z/NADIPrrnH12xGkVkWfrz8sOoWStcV
XoriNU7UDVgXhC2vNK7/MQdclOF/CICHLGZTIgtuP0+6jhgmcwz++ehzBdrzJw7g
s0cjSbOcjPAKrDYbSEjRm0dmegtQTD/kBl16wa5rAvIpPDs/GotcCoroaS8v/+pt
Nz5va6oL4WvushTaVXMXBV4CbiJnJV4WC2TRX4PZElqPWc1tX/MAPTtdJmRIislv
y0UGpJOlaMlLODO2jPsHU0725lX5m3ihZCrKTOuRDczNnU+b7u//ZjtIZBLApogM
EXu4VCNrkwLLVPDZerNo3r5faiO/TSKuIwt5DalH8trzDXk3ZOoOOzVINFnMb03V
r0QA6f0W74vnGOVBAL7a62i7EqpDuO1zZZA+xKnp4HXm7/ugLLcbGuDFQcL3lRCk
TyT91UbwXZgXSF6xKKWt77GtL/yYQr2rTZ3hVz8w88n22SAAHeLoO8kDCcfU0sHO
IulQNhM/CDcdeOEh6mIB865BbCepj4WzcZmj11Fs7+nRrPrTusOJJ6ArQcxdMuRO
Eti66DQMUtQRTVKZ32W2jlMep1MkqPbQR0nCBQl417KI7c4ihvRlIw4s1GU/fuol
ST6Em5c26TvjvQbtIJlq6hnHIJTrIkyaoqYAOlzzhpHmNc1A0CdppAB4J9nBMscS
r0n+VMS6uSc7um1EfwD8YudOD4TmCHy2phXlTcIYOwzAGiQ940DggrphJzzF2/pu
IqYz2MnIK+yZxG+eTgeRJb4pF9T+3oiTWb0zngTkCtUfw5en8IvG3vLIT709BwhI
VDTUifqDQNkdotymxPqjzoDOKBzw7vjn6sawiatFdD4QWZ6TgcBU3hz9MLVPWW3/
ssW5W109xinh2jbVCGMppmbT3TbPzXAu1Qxh2iOn6XXYSSPul9Ew8u5cxdXNH7xf
q5HleUVi3lTdCx3NQLSO3g2iFsHEpfxnB1a03jsLjyp6TgKUgreeBGettimxXB0+
mD7dXeAor23QKc0KLXN/TJmq+9i4LZ6mbtOXqfPFkWApUg7J3/BE91uPuN509wLN
3t1DhtI1QKrV7NQpQ9OFhc5OqfmXgqEGrXZNF8aTP6Aj/8azl+BdeY53DKqhMhxt
OMPVbfUC5ylrCTNOuVca9t2TyE2HmXs7gfVJQyRYJhIwrYX8vqNZOP1oMnG8aP6B
J1jjeQk6r19JgSwM0gHnQnMLXoISjsoiP07NQprMBsxXal9fdjIPzV2E62Bvdagf
VJx3ReC+ra5K4tPmRSG6kPWaEuHZ39fQYyiutP103hPcXSN332T+VHyZlsULOXiW
tkUzW2/QqnoDKGlKXnYS+XI87QKqSUCUjp+e8iuK95bXhAZWL0nPWEAxHtlG+sGX
/5cQNQfb2aAmm+BLHmbbQEDnbdFv6evE8Uid8oNFMT0s1W6KRk0UXRgPzNkqJPTS
Ef4Nu35KUuUaDoftPzsFRTJgaIBEGB8nJihlVSfPdM/AlvKQVGRzlN9p7RhfqT5C
yUYBShgPU7UAVRNd0hUnEw3thg4IAQGVyrAv+PzWr2/Es8mPC7faWXFGCgSAWqe+
JbQt/msPzlNN5L9d7Of96UhkDzfuJX1B2BIG9p8Fn87PCP6z7l/iTJ2WuZc4Lrbj
U/lVZ/jwZZLdhT5BZEg4+16D4F+qiMYGQLfN7SSfraoxfwjFB5DmLAdpKAz5qPKG
Elh7UGgUuPikza+ge8sa/z6f/a6pEMEgDuyebpx1B2/qYaNOarrrugNCC4hxzPw7
7K6d/gaWHBWstowjwtYkhUxLQe63k4xsXHYLnIO7OQSydTi719skJQ1yUvYxY0+q
fC5r7x6FaTBkQSgBHEZC1g4IJkTN2IZeDMu0SiT9D7Ubyx1ofu/yrceYNvvbuLyC
kzsMjuK2M2VlFp3d61OvzA+wJiT2e7PBNBq669rS4RX1QGeJ9oDos0Odkz4kCWEb
S6ADTaZYONaaEzfPbgcJehFb1TYy4DplkvvdsJ6xx7MhFOugmN7x+lWGixO7OaLW
1fSIPbNm/9PTUT08FZX6U/dFz+x53tKmqpe1TJuKa8alxJYcblzr+JekTXr01fjU
q9bHOIjmuhawGl/Uy80W3yXCjAbnx35QFf/eO+B606LrgKzwkohpnmw2qloAnpk2
gKrMARYjpeEY+0XAPpsRs65W+WNbP1ffCDST0SeqH2b5U3Rs4ivr+QQsN8N5dZOO
Ds5STLyP290VMgMU5sHRpkXBmHF+yRA+CBrxCV5DnKmm9RM5LHWpXmTkvLF9MLPC
nrrnA410sP9gw3dLSBjt9qLoGKQXvY3ZPZlCkzGXTfGWdzbxKLzDoYue2/Pcq2w6
x3zAd3sxxi22YLsBIjJL0Ta9kKoeCTwl2D02jCQNOdN0gK5oZZhJBCW52GYBodzk
yDuuNLLTGi/VkIiiBF0iOw36Ma7fQvB1ryqxeYCTH/HjO1qNTVSNTUAKDKhM3LLR
ZEjok/H7fSy+kvJDUDagMye92y3rHEsCNb+wc7+Oe8TejGmOwg/JzmG2JS59NVoe
KkbSR62IRm08zH/A24HyJIbEcUoCcK3anu4pWQaQ3vNs+ysduthxc08IadFU7LSY
QG07hL9RAsIiGECeB9sQS8KN8mmq2CSE1kA4eiGLSbTM0T4SVO1QYpwVW5DiHqIH
0JKQa9xp9SUc3hMNYrZ9+P5T1qiQjo12Qw8weerVcNzf91F91vi/MYfa9eJq8pgv
Eqqsda9SerQAHfZV0DEh6c8fQ93pE3CZxvSmqZhWJs46/57iVmwXDzDIzbjh6/Go
4N09IjbEVzndAevV00WUiHmXp+rPt8WdPCynLId751YY81Dm2A8DVPP4mcfcTFG5
z1cmDRhnioqnsGYdLr6gNKi/6FCF/z0A8/i7tBx8OL0+nAhjggdIWnLWy6PL0qNx
CHmRhTUZ5tBxkRHOulXKL4Su2nRfF/ElvBJ+jQzZeqz5wbI+l6gcOEEsWemdEL40
0pJ3mOzhxPLYQCD/ebqKbALDnuksOGSCv1OI8lTsfbwmNkB5kC2Ad/WU8NGFuzxY
5hkJcveCj22mnMWrA68MfDLXEYCDxprWSeEFE7dwvGNMgNN0bMp07Zx4G1LXSMKV
CVLq1YfMsYmydmu4zgvhr4U4eRfRN8siBYRSrUuuMU9dxu2MLoI5OmURR507oYL6
erClIMCNROWuXg44YXbZoq57QGfc30HxZcik3ObYv9grEKj/hARBDM9GJqipW5Pc
FM1MY9HmD+GicQboYZIHuCWtHv1dZvFjmKg3m34gCRvHHbD6tFes6uVA9ukmyknI
6+IgsEHwIChbfcSrSvAEoBZBIRzhMNvmW0PY+RV2e5A/AraTnP3fXckcYQVavqKD
nW+D27llI3DFazHCYndWRC0sXYyZK4d0oRWYWYmZ7wt2F28GcU2hilj1v/Dw/FSO
cxSo163pCULG1av5HTum4kO4ECpArw/rqyvJoiZ5aRcbWajuudFpOdHZ2NJFVYDn
ClhoboeWlHHZpyP8+pdU07HUiMlOouuKk909ejkgDsOEGjrtn7WjkOMqbWBNQ3eS
2iI02wn/g99FiNVKDCbSMlD/MWq4uG0EepSwP3RqgEvBV1waVCMUigjCn5vncyD5
kq9oEPkqW51TqqMcMX6ZKXhEaD3VenhM5iM/GJVPo1FnBUt1Hr6inlE1dZLcgHm/
IxjwgsmpnWTvy9L3zB1CQ092hdovUdQq5aF+ILtKqX5iDy/ijaidYpuio3TEX/Wc
PTBYl6n8fKk0Y5jSDqfUfXk/LlgQeRh/3eVaG9XIyBXIstn9U4uRuaKRPo2KX9BB
J1c0elB1tnIvGmAQmJOCr82aR7fLXreNnMj8zjREUJaHUNDm7bYFTWkprO7G9mhB
T7LUjYkORgCjJwQgja02p6sa5qAmjsIOXjotn5NH6cU5AYF/m/THNsO6khtrnq7/
9tdL+DN2jTjqTA4z5FRa/iepBdjxK1t3uVDaC/J1U/Ial1sDtiDyBGmuhb/YpQBK
EPiO5BVoZneaswJ73k/2SRA6MDhwjxo5p+1gxmUBc4vwu7DEL/CDLZIRsJiRfuqx
lL4VQJYPk5Cdg9myQlHNtdIo54dCIarJ//N4RuFd6SW6l8bY4GkyxIKSI6NwE1zG
hmLr/KMFUyct1IPejjp4kt5x0O1t5mSuoT8vwnkBTWSLhcs5wT0gu8kWeibzXyY0
IHT0JzAUSIr5iV4eP/R/19rua0F65MQvCFN9RXnBHSxYIdZGLrAuSYlN5LZ8MaIm
xuns5cC/IUNEUOEtXxv04yMqgS8W9mynOmtCWMSaHUBYud2sKTvNIeRgfeoXuG/l
ezeardmvPuwXnK0dPyrky+C2HPE80GKNQ9F0K/RGAxGDTAVj5mmb/0wwyvY72/s2
aB5cIQiGHU+EmSHWH/vBHCFL0sX+jUWFmSEvq6pdd+WNXTa+OZpdjRZiKxMnJMgl
4RdrMSXrFYA+nKhHUNyFrYm9WgC+lvret0Sv+mF6X249jfEwh3IdpF2cYzvsA6Vm
FM25iVBewAV0VSZxRJgroYLGRleddn3JRKjYg8eNMmtPQ3N3cavtNKD8w/eVqbSS
jibY5Y7JzX679A/dYKbiZIxPftGAj/a9O08Fyw9dA0M4HQT6G/d8HQ6X3vR8un6t
Lk/J8AUBKuI7dOumPEAiZDKfg8RNjFcx988LDqURimy/HSAr8cSyVlUx88qTLS1C
WQjEHQwhQGcbruJx5n7cnPe/XOkeZyw+9QHYAeaA4v6864iFVph8wOPjmSbTDWe9
A4ckcGyL0kT5ZyHycgEwsZsn/pAv2hEJgpAlfotH/OZvZzvHQA2BZ1M3o3hwMMRh
g58QkJn8Twm0D5YYT9cZT+P5SYyjENWAiSZ4x2OoKbQqZOhHagj0MtVbyfyKhqEm
1ho5c+pVeJNOAYcwQs0RVVwO+wAsoGE+mIgZ5OJIREjGK8Qqt/mion7qfj2wHMd+
j2UgIsSwKdm2nWsZyY8VUIk7O/7TpYuYtiHxw40OxBj5u/ck5ZUnrmmQlh/K2uGk
ae5NMcPFWMREZGF+NI41JdUJmOCjmMg1cRvadvnbtdqaEvNDNcye8s3W1g1sx/hb
X0kERlEQb2YEtwgMStqs28W54SY9dU6+k7fAHjJk/uUwXtNEIh4hKXDNz5+mJ8UQ
5c2X0r3u5ZBOeM6SNK4m2YFSEdqQ0HiengeGCIl9iEQGl5EN6e1MuIWhR6FZz9Vp
0zmpqUkjCxXe9PNkgHI7qJ+1UtNvUfJi7SseDHLBDoA9IQ9B37Zx4jTCV2ja2q1p
FW6YqWf/epq7QP1yQn1jCK/Y3LglqvLbSZY7Ub/2SMZZhQLTe5YoYNM3UmXkljLv
f9N5OPH4zd6XL/UcAmqWDb4+DPyenTnPTa46qyiu9KymS4LcpuyRXdTnn58QeZol
ETgBAtwz+HjHK2k02CY5Mrm5ZPy2Gz8lbdaHVQGmQlGeLZIXVzuMghIT7xdXO7Je
mc4aErTTSlXTqW9ROnotzaWKYvz1sDMJ+ucTBpkEkPU2FL6PsQODuh6jnbdyRVcS
/5IXl66klb7VF1fAO9r/kHP1FbTE39vXYNsvCabB/6qukl2DOQvGUtwS03GaGRPF
PVgTAiL9fwucSlT5c3G4UyhBeB7gzHDy/mb1y8AiyyAp5OS26oAIQUzJI34pArzd
TUCVntHq/qhUpjEsmui2aJKvvFJSyh/e7724zca+h7MikNOU5y0yptbdOcWW7BSr
+a9FIWeZIj8Xtm8WD78PaAqx8FGVRNNbxmr9XkAvWvbWYOnzoxSMes5LPTIy1fZ2
9E3/1K8XyujUAYrcg1EycdsM95w2IpiIVIMZNUxTOPT1vK2mqMdGjkMkaftteAqw
u9zbS9ziR7sRuCJQYFg5cFWTVrIa8/CSmKcUDA38BQeqLxAUXSxwgOIh8ZWs/5/y
hJyGj4hCWUQACXO1WfsU1BSK1x7upDk0gHKplEf8nKa3il/3brIws/Zvix9hvu7k
ox6MI+BHFd0FFEcY4PS8muDMg8EtGOmDSj88vzFcDeVkfHwcVioHUqnSHT4/Y2rV
KSX31y9ts7oHpOFHJIuoaUXKnqSMLkf/JbwnHYUTdtMkUXohfHnNZJS5YVsdiqy5
iamflo6QktLTjgMoAL3oJQKHK5yrrXvx3Yr9p7IWMbyHH+yqqHawqPEw/dcQ8pKy
vTW8JxT3HFXs2txLu+ChIzMNxTs/52oTTS9XTYaonoYE45GB82rNz7LV97gckqRF
t7qFKfOO/RcmwIJ0tBRpqElpGxHo1Z/EecvcAsoOAInzfMkdpOMmNsgZfTmvqTlg
zRpeNaTzyCJuZxTHeCxoej6S/atLGy/EXz/j2gOpr/CVYjXtINPKmiHig4uPCcHi
ExFAMPQlskyXlgFfn5ZTvRvCRJecExrqP9Y52zY6KnRrKghBKCtK3GzJrG85xKIn
MDO4SSHPO7hufmE3Odle0jgM5RUV4T9fyLkcCbpWKhbihkHwz/qP/3B7A35/yR3h
8BpUij6vFdVHPTamicTilkYLCgveVhujSZ0sx0r8mcAMFsjBRCK/58OLV0m22PMu
nn3O6QK6DIt3pT8PRTrxmKoEOWRFO2Kp8faEVcueCYcF9h0nA+3VexiQlr6yyMmJ
ZRQIg5GpdUY+EdnUwV2qMavHabEqd/4IGEScTj/FBXCRH6txoSAwVSbnmnYSpRz6
26U5ze68yIzdNTiMEwumfMWEUMTCCPzxmZe2MEFkQhit6nvlLElJM7NCgwziZWbb
hTSeZNFmT0iraQGm+nRmKZxwXqy1aTW69HWaW2GcqddxObZ7OeNkfRFuSvPPCBWL
jfUowtCa/iGpUezU1cvynA+q6ANgD4A2Y5Uu/p8CABBy4jhMFJrBKgmh8cpSrgnq
AMxiEGP37RkHFwbk1NIpCfgwlmlkkACehj2ZeJ7uC/oJiKu44ITjN/qHQLEv2i8B
/PykxcApOb5m+DFzOLWU7FiC2PDWcU/zTJ6SK3zA0go6WYVbXQ/ZsdSl1ZySL+X6
b34fl5flWmDX9jiHpNjVtINM9xR6oVcVLftaoVBFZxYvMdqbggtxnCyO7oA1rRP6
6pcg+q2YXHT1dytlpptjXAIEcBX+oyVYi6bYROWwKGLJkdoIsS71LZhXk+mXCSgt
H96Rg1jfbjIjw4rZdPxF7jAAvKSUGVj0SdPlcKLFExhDhjRkgSpsRsz0ZSw2CTIZ
wD7w68+geiRM+INo0+AY5jKzSgUbUmlvO7dHHz8c2GUntoOC/8uEnoKKcyQ/TqJ7
SE2bbLbTAju94Xzwwbtdqe9tASL5RBb0IPu00PI2dxZHMLwT15Tm4KVYXDH0y8PQ
xKS45ZgTmII66pQWThOlzD2HD92pzqeoeg9ESNDDf+SDtDdD/vYEAMLu2+LPg/tw
i6XfB1rB7KreqRBDZzjB282DXcblCO8vNE7RH/Tl4mWh7hcZjs68NkMeTlqIHZTH
MmFE4fywZB91rBTSlteGud2qrKtjQbLR8havO6qCU0tGV0zs5sV5XFxqKGdXBlyh
pc6+gDlUH6zXOu3bRxcp77F9kFMa+LA44n16kolYUWU3oRdlLdzbmDbq573LfcGT
fWdR4Z/LUqevNM7Y+zDH9O4me4UJ04XPvjArBa9FbBM9e30vrhwLFl3wBT3ZNzdy
FwOxqEW1bDxrUZRcpON1KZ/3FHpxx0nc4ie3tsmBm4cVIHtR88NtYB8gtreZ+cmg
njy0imsjRpWj9A07twmAiDzYMHoH+/oS++8XhSUG+kEUt3ZNL5i1R1PcPL0bRjH8
ZvDrClOEVUHPDvSYmEbOh4eiVz0by+xVodi47nV2Lq4Ur5rDFI3hJC823/EjPqUx
nz0lo33X8PQTfmx+X21KMhPK8oLNADMGm9DgBRdmWjhSb/lWB9nla+rYCb4K4a1d
VnHklquKtLAyOZ2jvw3+iaJDBB7+7wSFFAlUmHlUseWlVWVpF7q8z3yMO1j+BBwz
i2FFRHOQ3dUk67eCZmA6roT6RZk8xb/2cQ/b6PQazHEp3pySkv1r7cqSgUqdQISb
cjJ+wneYnFua+uTpZz0YbLJgeyFEMchi/fOdU8LB4s7HrjkRIomiu9qD8SThKYr4
DNyMZMu6OJU9xhZv8jOJD+cPqu+HWWoJb49SW4MpI3l0wk4HXFUVJCR/+MswtPg+
4vKz5RJ3WeNDuY2WpsusK+f+8AXBX8ReSwnftXd4npLDL/9W0Ja4qIRhh+LO7QCp
1kdlPUi6Wg+9OP9fi19hzz9/gl1DGX+yij5Rb80/kIo3QF3ySOrqEDFlw6OZ47hd
BIyaoq2LljSR4AYbVF5FWcr1KlRaG6P2rI3CW0CKcVRQ3EJJKKJQ3RyrsRpQgOgU
YZAzt6RBe9SU8mPVvehbeDHKLrW+zydqTVRYarSnsxUQRB99k3Lb18oZO8kpjjWY
7fVwXZJIZhcVatKslm5vYXDT2pUviLzh6nF/kUaQ8n67x38Ce0+D/5LujaFydQ2d
DR5NPDF48W3UvL2qjluMcaY+Duq8Egf3dc9kxkI/xVL1TzNjsk2QjZpLiXJTC12n
xFSjcxkK1hfumc2OhUlmGZNAYn4k1jwgnsXczhMyl3do20tF7SK9k5elU68Ko2Dk
udH2tc2gJCnkKYZLCq8XFXb06yuSnI8hMSLFg2gX9oYWRjfyMCnHMGQW2SJ9erbg
SdOrXoXljZ4x8AHeQQcbFbAXiktKXjhhq8muf4m4EX6QCYP9/CFY5yuhyrKfJYyB
SJUozT/M4bWO027q1mvCMeSm1G9MC5dU1zwX0iLxi3LNsHUx+N9ocg/z4fDrqXR4
vxgvYypd+8TwOwS4NFwwHOlKGs06UfUj6YuYJ78ySbFcWezOQneDiHgHXhX0XEii
6TvjaSivFUXR+Ju6QOFxMNJI2bpRg3e3KEDR6Rrkn9lCO7PXvqwcXqDn5mdVNgti
IxH7B5w0Jppt+uTC5fv2jaqMMZ3o3H2jalHrHThIhtGj2sHcH3iTB2So8uTHxLu6
aqKl5CHWvStwga6ZTNo3KTn0m8SLxG3VUSzNHZaa3GnU5v7DP/xFpKcK3FA8aq+V
udiSLvavgrcEqi2vcqJ+hhpROhM6H08D1Rkc0DcwkjXOdpivd9wzMR9JTv8N7Fgy
TbkDL0MemAOSP5GRvo0trp3QbTzW0Ieb/DoAxwkKDzMCK5sOgvU5iRF5DA1qoKao
HbHjUVFUDu0H6GOld6GYGuIz+MKXHzHCITWiA+YO2QcQXWFYUOcqEN4a3XoAHdu6
cDREYkW4E14BKQNryNc/ISdndpYc2y2LvcZQHMLGi7T/TmxNPOwbzU1pOqBJVt3R
RIAcJCp3APhL1a9MORxgm5KMRtcb/TVd2Ws+H+NDjrYUIYTszHlPPsixW8jaQrPl
+mAHRwffITTlet+80IjLdu6ssbaVUr/5lhTgxtjUhtnn5vGcaezc5zhCBQaAoLwd
7tJ623fbBJT4nks5Ttd6pqmoS3wLan/b4uwflGM2mPy3WK8VIlDSc+LJehRW3bMu
dIFb/PcvoRRvIOLblQArCnFlO3yZlzMJQ3GSAMyuTZYGiIkHB4J8pHdMAcmsPReb
OQA0ATG/qqHX3GxHtXD2dAEMKmzV9xH5DEKnUE230LPQ+sCXhwdOCsT1RAYfoTMn
tZvOJFy8JGaJgfqyKIYaDh4DR/8yeKdnEgS45UJZ/bjwGmptEzyNqsEjV/JyuXAk
G2cEo3TYrRQxcNd84iUTrlYmczttitPeswInkevR4RpLiqiXPLYmdX9Fz5eKrb7b
4WWRahubYQgQYNCRcDJ1etpnfO5RqqmBbx64D2C0b+SQcu4G1qtXMBJzsB7Un3Oe
VtS96Z37qs2sdWIWsvhWKw/ZaINZ6wyQdhfz48BKpil+1S15vsKSqgW8b1UL48YI
TgQoSQeyagykdPFJEBomhD/gXxPeMJDZGRrOEWOdc3f5BHnNCBBIT5rOtWKMhhu7
IQu2xgsHNW/tXQoRleUUOIGPq082Pp1/SM+VPIhkmDLAI/GoGZNXiyopGi/3+u6Q
MRhq8/n/r8dWtirZqtaIihhaqneG2VL7sex/YI/hpHnN+Axkk/80ilWKmIoFkRyI
h0PHqx8rEPOWTKS6bcBOA2bI1vSYysGA+Xbofp8Buxua+zzDlxFFlvl5Xo7DkmHC
PAzzi5mBnRmGCPwuIg7c7m7Bh9g1NKYkneb3lO1+Wx3WqpQFd1uQSErYBzmzJX7L
cqRUCePyLLSr+4VCrTolRDEXRSvckd4s6GT61BTOd7mh5uKYrwojIGdSooe70mwM
ODwogNQauGiiISzp3bDGNv5QydDWnVcPnuiTFs84SGvIJtWv0hxp4n/gELQ/ESkH
Gm8kyweqKuIVUq/YT/2JVuxqSaCInJnZzWoTdggXiZ1vsmjPHrxURVXZ7J+JyEMH
EvZvNoqT0MbB25jAQMMDPxWR8iX9/3kf+rqxoOzWXE8egZpm96R7AjRVbskmYvp0
4n6z5lpPeAaIAGvn8/t64SknJ5OqrVpga3TVQFuZ4QKDLSHOw9B2LEbKHwGSJdbI
ghB3O4e3fKbwOmsXlMJj/vXUcsqbYQYLptkgJOwSpQf/mETDTDqtNcHaLTF+Y1QO
ktfiLFWLOfR0BKigFTgS6VjKmuLxWgkUNIZLk64RiqA8ffq1Ixk0VYNK/IEeiwN3
b7SorhKoAppMvjWzRF2W9eY3dzOK71nFLzv602oqH3dMxJo5vVzDBIEGiaaP6fcw
Hes+m5FKrKzRdlBOXdH//PcTL7POeqsD1v/PJbUG/AowdXOTcma4ebu/zUipIo0h
cRamdJ2aTppMccOjWNSQHUWxpQAVFb76Fb7cDU2g94eSBWnxMnOrqMIyUvnYFGuj
KIwhs6kvLTFYN+NpT4Y15wKhjTn+6YuWOTD3ArBbIM77wDn3XCQ5ffsOZSzHUijk
o+ssnu6NFglf8NUjDOkezxsefNSTulU4VpCrv2Vv65gWXoXgaaYaGY61HUHHzmZZ
JYHBDjQcoc93ifgK2FxzHh6ZrqNDgeFH68oQL/Ysa+jicJgemeEc4NrlFI/gX+re
Tv9pD7lB10HecFXs5H+YBdeWCdz2R+aUC8HT7OehUy42+2kHNoL15Aqk9UraMXNT
ElupkDjV6T9u0pux2GRapPT/niIAsn+voeBgzIq1y1RIBotuzi9bt1FTfvMskEUn
ZsFXdhUdP1VeuvQP4SV0rpetZnHzX4th6nSTtOx0+We188BEv129kSYEqOHW7Jly
WrTKQtjx9QpowSKzqy1vvNweBQJk7FPq2nVMil2yJliKyGJJS2iy4J4f/txGIDx3
rNfjjiN2IwG68jaJ5ogrw4oN7yUZXQdAEMRUmrjfZtNTM8rcqYN4CiFjvVvZRNtZ
ayS5wPnoRBcMu/3/hXzLSNSl5b8mt10TwzSCDMoRhqfWBjcQG6ZChzPLJBTHbitm
OoK3nO1mM5m+L3KeoO8oud4K9sUz6HI7HD+qjg4rd44klTjqp7eETU44kqXN90zt
4OOkK6cm/vk6LLQu8fgDPljMFxR2J8Tpd8AHy06WR1Ihr4nYb4TfH50vLAe5QjjJ
MbYXt6OPsrQWat6/HJphWUUycPSnunst5dtUC5sQ6v/T0wMa9U7X768tGsF7sI8C
MCIgEXExmIaW08cwiIWmR9Bfm4TFSK+QezcUy7s+WF40InqrZQvbS/fI513Vqa2U
OT0KgwJpYWS/PFNCFJSq/Cwh1fNiCC+NwykY+34d2/PfBQVp0o0IPUQvJi47bR++
6OXQLsHGEUrz+6RY5XKmwDRIkmbBWAW6FJR1g5kuDw9hA4I9m4UBj1QnqQOuTICf
PSkmCQ9bow0xgFDGX0RlaPIWGRC6oT+daZVwmzVMHwYkURQR4WD0xJ/8ht5OndVU
L+zKCD7Bw/IXDl6n0kLdzzB38d/xv/yK8uiBgcTZHfADW5vNS/syEkji+sIaNvjv
hybHsxlbUQCyvyQF5kngNdZwS31tslJlhsU9jpUqrxeBiYYWJBvIrWmGy2h2KnNS
wI0nHk5Kj7ws/34+8D502IRDt2SzxWi7HLDwHtUH6G0UZy/bIoN5WCZSUiSA4f1i
dMuqtEyCwSqD6ZyFRwXXdD15XxDiT2/gwarVtsMJ/mbSWEzcsip3uijSdFFuIRfI
xd8LwqoUZ9d6KEFu8BwmRW7t9mA91wUx7VdHyR0SBp3DPLxYdr2BzEhJUnXN4lxM
TqHLnJsutoaMhG5Nd2hHXDIS79AciYi/UjND28EmW7HLTIUZzL4iq1dGwmQTdR0t
YPIQfNXZ4Lq4b3f4H8Q9YdBy3MUFyhxB5tbCVYbpTMFkfeSrvsyRtrkSB01cjwAf
tRLdVBwp+onzaqTURdJQeBQBcDy5/VS3/dSK4pb2rYUVQlEtzHvHweJeCwfd4x2y
D7Q+C5liZqZ85rdlqeyOLEIYfEYlE+Pz9KLrT4RXSOav886+ldCEkPc2jpRr79dw
IBfWzGTdNN4onclvT/vAomaQJisZP1FIbG+vOTG+kd3O1lVGMqwud9uB7N2zrI99
B84xWks0dVbCXZi3QtR8JeWtqvBRX/D6bUxANT5QrbDSMuCHaj7M4czIcd/nTS8d
qeE/CfYo9yvKVsAlXKbJAf/jgx9GVy3floADkURdj3/97koTKKZqkn5b828H6pnx
gAQ3wgDWYOs2ZpHLSVuBIS6EW5RtWiUcHX6u4htUFNbvbfPKgGmzTBl/wRQWkKqJ
SCLV1Y/QZbnXusWTp/mWNiAeZDjYRuZYMUcTl1UsMpT3qDMQ8RzYU2BpM2FDh9VH
c37f+rA2FdGuLEWCUUHEelpgRJamNZa7nDrGt0IX1GCjPRB5G0XdFdvZKTVlwx/p
5q24pRf0nXYrIqOnfTUephcMa2+EtlniUWdSS7ZSYMCCj3Etano/lfGCEicABVv+
h5KEsy0QLouxcJ7NzH9VT55Kd7CRvyejHSmy/qTn1Bvvo9JzNjfkgPrfMlB7iyWh
MhuAXR055qkUBPdZnm6dTMF3+jBPpU05ITsFrmHNmcKzur8XquGFf9IxoENuqB9Y
Cs71hgipppnM2o2++EQXyH60XYX9xzf6jXsIXv/BTWYUFpaU3mGA5Ofojf2nQGXg
YSrrUhXl5ZBav8E3k9VlhtUxrGhC2N+AsgutH/LLh+mU+42YN+4jc0BCJHaF5zyU
lrW7iVHGCv3VFFd8uxCzTYUDKWAE0VC0Mdd8nEgVTFcPkCZOx9odI7lnN1Zbvz/O
3enbqoc6bFdUe665owWfYtveVqwUNjDb1whu4RtL3T3HJ9NeJwm/J4p8Py5BgZy+
i7TZGBCmPmrXYhgcQxHSz7AXlp540+HDcrqoi+jbPub7HCbrcQP8tr/jEdyp6IaL
zQZabkGIuJUHuSIzgRspooIu197qLdnFumc4PMzhziCvL1O11fWMvWNDVsM3bUtw
FhWt9fNfUtwhUXr0b46Mb5Zbh71z8XQtsJig4T/DjIEqZfQSGRYuaC8WeToXxHor
zwKBRW29zMJ+qKqMQMmblwNc5hbOb3sHJIojI0gN27KyHp2W8LBP7gfxOIEChweu
nHP0bhtKcjsbKh8KTwelRB9r7rwbTyzvMy+y6AykB7MK6JfcZKmap74EiwABhfAa
EjVR+X7un1Oe+k398blTwQpDElMtfhdCmFL/lVb6bleIzJOGTQW9fei0sbKZEH0T
Lhf9tBBbHFudF+O5D75jhCHsxS27mln5+WILKroGB8pIauDUaSgJlS/J9K6j6REN
ne7LntC+k8n1RXVJC3ven3H+avJsteB/vspYufpZijgWq4pkRJBTWRuPct9dPk6b
r/4RJItmTbzTGeZyQEqKKcKJ3KBPDy9r3C5v70LrkXgZf+EndfhmOpQq4qcrE119
HYfn8JoKLAL5IFbMN4mO2F5LPTPnoW/kGC5r67vh840DJOAbY9Ls8QFr8l/biXMh
kRMeaX4hHfTU6dxx2s/wh5SMahPggHHQujChfoa+uxmZNm4wDlnzb5usuCzFsg5V
RL+b1dOGefaa8PWvUQ7rhAKdwy52kyR071CFZr/QnF/o3dU+8pB4bxYaGNrOhg0S
+GQX3hp9WH6hArhvd8MgPHI5s8g22q9Vt+LDLCdBGU26/KsGm9IebWQblt3idmlk
tuP2p5X85JkidJ01L/pcTWW1HM90pOF8RTh/a33Npcyhm0LKlQC31o/4A0MPJIOQ
/qlv0EpBshFuTSwM35TTP0sP3ZHO3Iy/Ll3UVbfuhedFPbb4Y/iIUSgoPCE7XqrN
DWdpCf8zoY+mP/62JZ74nQo3luD/MSZnOgujQeoDZhgo5G4ajBdVPzIkMF8ueR4+
2aRg26dpV6UEBMxyTRoJdThjraUTUAUnlN1luUhrk6HWO6lQAUJPwZD8Hgwv9IkR
b7G+SbzH48MNy1Icsn7ugOVoHZYlfPd49upAmWVi/f5I8no4B+AdQbFnm00Imom6
WwrKQ0FcbVoGFEMgwPkcgbXbFNh+XY3xkfCTcxHnTTetrTOUHR4XBAinafPZ6pfJ
e72hjOYi37JdzS5sM6sD91YQn3pdO5BIGNP51khmLC+AjBbqaraeyxVm8pyPmQS0
xYQrP9KvvqCif4Sk707CrSZMOA9g6Va0fxrTmL9gM3ybZ2LJ1D0e6c43vXZc9gDj
vmrKpM2YQ47FFFex/bfdel/M8Dm3au8IVlvmxDqc8iC0bHZeqizKBm8Rz2yVSQHa
viw4UPO5CJAplFyaUY7DLiP7Un3WR6aa5LFe6d+pmd57r4UmpLtyCS74mg9cTg3j
b5i0eLE2iD/nRc7dUu3Qhiu8psPMWNKePJbSFsD4KOQZLKcBGw5yg9SVV+jdylOi
St2PUAFVN1qhuRjHYxSovMrU53Rcv3BRIGv8iLqI5vcKUhtsl1WRwJm0dSpIFAoA
thJFVYRfcQzvkjQSamO0EzN9r3OxSN+4e8bfnc4y7SQ8CZrp6CGFB7e95QfBVj/9
23/VXb6eesn19K+KCelc2yIceZ1P/QSYKH710xlexvcQpnsGtQ990dCVMAWVqqdn
+p93XkGwn/HG3kAKb14h2kBUpK9f/vhL+1uRGIIbq5sPCuAv4Om8vucbfb9c2iLf
6Rg/54hFKoGiW0iiJMZQ7EzF3CyJP4/xNlWqK1O7tiDQRuRAo6MK6idXSXPNswWA
mV9p6+EJpWsm1yv+Jw2sFwhyijnde01rG39sjdCGcVWJMsNpNrUHG8n5Br8WijlW
pJNj57YSID3oLBRiIyQBJRtUheybpsxDEPh4ii10JsMrceI+sems73YlsY4DxT7u
49R0UF/WVuj2ZSoyUBs2ckUvz4d5MJS9LPE4KkKYadINWgbMqFPAJSx3H59+iGiZ
Dm/e927U21Y8XMcD2xAm3GNQGRqd0P2UH7gnZAZJlw4DSMPIFxp9xBEafon8/zJs
hKAY+f3L4jw2UmxGIjez1by4p1xqRzks0M96db3NTSsvsrLDOE7r9LUDcSzqGJ3C
RhV5bMcsdsiFUxEgi4mKDxApYewI0LQjI/Ogf/LWvZ+fvGVvxlAvZ3zYIKGWdMnk
1+UspynrV2FvipUFjU9XzfnlP1lUJMCvm5wLRhfZU+shU4QfDBz0VeTFj8kJZ/NE
I8YjbtIqCxm09jGgvIGFIQhAAhOiXumsDP33+PEcl9ehyH5dgBMypLYOUIMfslhw
w/w26kEC2uU5SV/LYlIeYIV1eoUUvMIRIPNII+lLpunlxSMrcRQiUmbop+didJ5R
O/s3jgBwMYdY614tneO81nOHB+N+3Ud0/C1SVzGvIYLv4dv1crm/499CR3A5fIGD
g/xvY4spV2IJ0H5fFghcqrQWFUZATcKT62mC0LGPb9OlTW5CgNHFb8uYbQDXTa1L
l0vJVlgfKm50lP0Vl2tCqp9hlaRBtZp37P3w3LUi58v1tfqWSJFtmNTvlZShLZhH
tjsLNz3itbiypKCF1QKWxXhsPzzNMwY1rf+gYKOzbYwfDG9Y956UNDxO36ivcFEm
b5LtZFZLe/HkiMBGE1B1ekwJEokV8DNqxpQpJQziA+fnwZvSvAfJs07wfD6TyJ6m
+Y1KTNqSqfKcTa3apFHSSInPX1AYM0y6p94KfgFYGsIqjxn9QXJpTcPLsGBH9/PJ
tYg90LyXVRY40i5CHJut/0XNrKSXMmNlIO1luv8Ixqz1A6/XtKIQiVAjlZRvGi5m
uzcP4PVL+j3ckjaPGl056ePQQ/oFvSI1usdWZk4LT+YFSGj6fqc/smb5hw4oM6nu
BQxU7MEVBxKOC/690tmnsE1f8cmqvc13d7q+tEnxJJxN1yMXo9PJaDJrM2/vgvJZ
xfW9bnpz3x10xh54kGHKux3hYkyaMkHl5G0hFtag3biKcEbv5wWNN3X6vO6nDkKF
uO6XtNANRDTkxktsgWwRd1SrHIOlh6tMQu65/hqcalhogYj/ORVyrZs8yeNVTrAu
vVXI1EorRQJ8WxFVcuJjv54uyU6/gUbgQ6ZpoWjEYyz7G2AgXboBhYptaLLpyq4P
8OTOUmgfkZsmpsedcwx28/I+KloskJoyQs93VYQGEmRNtNpcV/vkhRYI3G57/9ZQ
26ZEIlAeaI45hWkOVdBiI+XkmODIpAySzXMrU36IfRAtdtRpEBVTwzsD+Wd+z685
PhrwyOku4flvh4+L060AJ2ytTmB1zXv5g1gyqgVzvbEvn1gG6fa9GBpBa5LRZDSO
4g68qUFk/hRzROnQlu8n47hmlu1/6jC9rQ8ScecCLWDjmCNierHmLtJAiiBG3qwB
dkJP9p31DWsrwBKKvdje0cEFXtsGo04MooXam57x+//Um4sbKO0u7/g4syLifuc6
iXof9IoksVGMUPxHmRh2np8LBIVhCQq5xtwpfiGhwA4FCQSI/f6Um7Ind6S9WesD
q0wF8bfPY/cFGZ1y/0qeQsR3MRpnqGSjI8dqT4f+6s3W/zkC6cor+mieuf++VUQV
8z0KBWPRptY5TnqCYnuuYcDGtoSiOUKCfhb3buFA47gR7SeGsHrQpGKyLEzvi/fo
CBIgLfdUPAG3nKmHmaos4PXBPV+qwm5SbMO/G9RNrs/aqLWpASreXSDRPCkaBs15
KlvJs8Pqjc0CMfRtTOZ1R6YuIVdeFqRv7QkHvnTC6jzQ3km71xvc+fMz/0yzThn/
qdNIgd4Bk2W50LFcYaBVydJ+40cwEX/evEkP88gtIMNYIVA912wZpH4l+PTyXjZo
+NeODKhiqy0GvburjjQfgkvTwc9OygVLUWA6VKUyLJambOEjoT2qcYzmE0cU2mLs
xabXW/NqAG7wVvp6hHnobgVjYPVl0fi+ZvT4a5VF828NAOoPLmsFPyT5b8OI66vU
n+OZQ3Iq/So5ZJUFbldhbYdg1rshl+R5takn5U3Ekgqo150GGvqmcVLRwsXQbmge
0UrZ3Rh93MPoc2CmplXJ1AfW7N8bfUcCB+ViMILUEeITrMRLiXdHfpGOqYv1o6hz
wIistO6dH+Ri/HnZOoUsPP9Qaiyd//ugHboVd77KouAUHKcvPHVxxpYQuSgb82GK
MENbWy1I7XF+u06xlruN3NwK7fvygQGeUzpLRkIfFMmCma4pUE/ZKnIoDv6cZv+j
mJV8mIKtCadWp1mnWlacLC750btIYidFvBsg13B/7Wc4rTmIH8nAdZAwk2xFf0nb
P7YziFR0v7VpdpFmyilXDuJv5tYGFVgD9TjWdIsuAVuzcOkQfdRvUMM4KaOmFg9v
390nx6QDWVHkcCMwaNF8gTAqqpwn+WOihJk8Wl6dfrjt58PHlk9qB6XOyWF0+1XU
RzgadGJe0cEeEwLCljB0eW4AIlsmi1t+z7ujPE1Qq389HvP23agzPRtgX7uJVxNH
xSnb3wstu2s8qr8oXEK4DXF+tB7I1rDOq7Ke4/Y2blz4Uxig2LdN0yj1hN3sF+zR
AUu0M+HqWK+J13dq4XUBj3ddjWEginsqkYc26hh5iSmkF3zpGAbRb9Diq5vcskGs
97G/NB0mOnsNbFfqobdJox2o/MAezU9nuyyEeEpjEq7ZbwIfNivEp32FJ4Dt9eL7
NKQdFxdwmVLc8ryYejqAAgz7WqZatZZt7XS60d4GwUbQc5XAXPr7rzUudSgl14Nk
uTT3QFaDU5yRd952G01+MaP1+od0L/fk+Dygkj4H+qB4NBrqYpMoIWAxtlspNzqx
5NFTFvI3fYaYFGnSx0OTf7AjB9x8anKqOUdQ6+dtaFZVXHBm+E11tadaLEKv9Fqm
h3VCxoiUQSNRFIjSUAkJbnvKUcf+edRsj0j/N3GrzWIxlAdzzJIz4Cd9M92Q/INu
WbDQChH119oVNZ1JnjCUiLxMA6r8G4izdP7NmXcHuMmEd8+oMVpmSGATwUx4z4Xo
VbArB/Zi8R9WY/ZFgF0Kz8arTCrxNMTlfg/rc3IBeSZJObd8+F/zAr7Gkm32z4Nt
jYaueR8usO/iOS6O4k3QDgekMa0hAcZy0GShR5HwTW4w6SNM5rVl/ZYGgY/zACpf
5ADVHjMch6HCeNIov1MJlTuehIgUxPuO7a+6YPCHFuyTu+LRWs0lOao4WdDNgYLl
wkpICmsGxW0yrQcaX06pnP0VO58YVpiKU6eRAAVaTSZ0JPfoc2xIudrUF+FV3L44
1pAlorwx3031HvrIOWiFXfrf80ykHIDmrbe0k24CZS4kSFGFq5R1neuUBsfP/dRu
OQO8R3YrvmVGlBQ1ClTxRxQxeHCj0s+8D/pXYv+slsUYJ3KUc4hxq3o6whkTekDO
vLe3CI2p1JJEdMJ8JfoUoUV5wl0yYxvkfMTtjnS9Z32i7YSPT00FrYIHpOhr3cjZ
vMwGFNqT7NEX1R7r3Wc3E5ibiiGRDh55nUgbANMTmL14jJybSaanixYWYKtC2ULl
ir/Fo+bw0Geaur7XCfKFDU6UUIqaXIOPzGTi8ndYKmDIHWEpknqakCDrqllZReKG
poXp8sbSFZCG0oKI7S6CfZktImJHR3l4+OG96iUECAEzo5uhuQGYyexv/EySs8Gj
S/fypqWZ6X1ew9jOT/Yz6T2qKVx/IK4Hx/sAJXyXRMlq7Cq1dI1UGEuMDfhskm0x
CthBS94ls2uYnprcor1pYnGDqnkZECDUZazrhOy5XXvsXAO0OVCXAWgY6y36AKZH
lTwGpw4Id6YRJFYJleUZY6F1fmE2ac4GAQD1P8iUZjKBmYGkI1vsdMYt+Jbn6siU
TEJdac7jXBy3szlGXoyxR/d2VUJOkOGml2MkjkzZbBVxAr/Px4jP7NVBjg36Z9eU
0vE3N3QEACPenuFdYFkmzQbgm/+3uC+0+DHyjdBFXFAKmcd8KOmO2yx5EV+MxUtU
CB66T8W3d4l8FGpWxtg3TAbpiyuIdyNzmHcLbYZkSbxqnuE8pR5qPHjAzZTf9iMt
d9lFeWTtvrGIsYacz4AqB5mhDvnsRgw8UCEW7IYq/lurvzL1YE8VSg+twaiiIAjB
sNmu2TLFk2WWuJM1q3W30H9awgGZ28WabiqqHvUbnxDWITg5y6FOkREBClHEPVxz
Vp7aMtRHtz6A14c8ySwERDsmCYfRxc4aKXzooi5bvIz/DBmpyc4lXKCNFV579Fte
ccRRULWqBhqKVUM69zY6chyl4BX50yEwrGio5TafrDi38KBdrFiP75QWxc95/6EP
FmGFnPV/CMCEKf/QYLPYzmCcjKDNBYO4rP/0exLO10KUAZg1nEXH8UJNBPAYCfKn
fUgYTNoScP3GeV12WN+WSfv3B8TZ2MRGmDuF0uKqp4QOc1TjRH27BVqEf1u052VL
2fdRjf69EqI/I/D2ZXPSTsFJX6TGF/heqQ9O/XlRJDRfnqlx2Iu/c60X4l1TLvJW
S3eJqwWKGu/2oQAN784wDNMwefHx4U2WJ67Jm2fDilLyH3VHlWeX0s3X7mJjnx5m
vKW0++EZOdkXWxtYu8eKr+l89Zuqo4kGzB2/4sbuL0Qsjj/sDqrK57N5pgNQCuGi
+cRO06jeRHiT4Fn47PQNK+tFpcmbO9S/mVnOJTem5Cst5ot3/V3k7wGfCY70GahE
14NBESw7jQqYDXWQsai+/NZjYqU5q50LkEhofQfUilvvr7wDFrwJ6SSFKNE21Ivt
mDTVmEMSKvd7zetYH62Ta6Y3RWWCfjPA6kImioXS6a3XctGiYMSwiuF2bFLiCVrq
S1OEhkkl00VV9rdlagS9ivwpfxcaKGnlnRPmtAcJSeytSKJ+NNVflyeoWcDlQKBB
33vwCD0FTsD4jcQcy0txqIOEhzHkM7/h3/qhGmRmnC2nPlARATGraM+WEnH95Oya
F/7EUwMoiLX48EifXIklh41XweLxSVdLCUNmVHvDxnriyALBpd007XbNLgCaTScc
rYibQDFvwg9LU/MRnkKI0sjzNOXP5lNgA/QCbKduP6D7+coiafcTbkpixxnTcdSP
9bu8Ork/JTha8nvHEPN6nsUs9uaNO0OGhL8FSoTIRomf4vVTbSaI0Rn2dY0vwbLZ
+2zZiWMTRO7NBEQDLMjXsR1R7g7Vm8oP37OkfHkknM02OcXBzA8wlTdodgtzAb+5
M0nU41kulajmMq501cKixONQlZsf2PjtFevpFf+XNhwKgkk5Vg74PgECaHxGCD67
ObpTIySZcrwNFt/OilTFMz3mdljN87f76jx/8M0YvLzEFuY5SwklhTACtbLk3nsg
SJEtNsTL5GvrFI8HNpNN+FKbfODNHEik7VdwciuxpmL1Bgu2vh54kGdHVwQ8ISxV
g83j7OufmB1c8fkaAj92b1dSrNoR5svkbbaCamNRRXg3PpEs5jb5i3Q92ASR9rb7
OgFOKQdkM35Cyc0OE4EBvYsSgCFvjUD9+5Q/uHLcmcUY3bvpap6ZMgYOndE+/pNb
kqAZxNR0gxV6zi1Tz6yfMcfdlJqjVIvs4Dl1X0T8pW7FkrqX+G55a7sENBMv8GNn
khwwDviJS55aZNlanxM79GkjcuyGJC6EFoocHKxDdicZMPg0SyvFdgU1OZVIPLqX
+sfK/B5l1ogUxq//WVm2Z2tb0XT2qUZBpwzZS0e8U23qL+cNfW0meeE++Kp8mgBD
t+8JbQA3BVFcv9aYXUkK6AZaGfVKJ6toWnFCMby1rhnoQHa2txrBkdzNaiGugMzb
IxEmGoLN7Kv8qD/DuX4qXWlbJNdsPtgkKH2jAjjJlojPwk5azGcAumIxsslUSGlh
xi6WG5z6HXnhPA60DN2WLrj5/N6U0akcoEXsv3j4hQ010mO2o6aYVldCzHR0nWHt
fJtFwFgC5xXQdi1q/SKA2/GV3yMRnxDhQWCAVRjdjOqhk1eG3l7C1w5XYgo0OfkM
WaCziC/QbR/cTfe3CN+0hXfhFjngsUOGLZYtfSUrjI4S9h781MgnB+9F76S11+t6
sD/7Ee5bP86cJKUFCNwh2Pn3LB4Oqu4RV78NNY92QstuwDo55HREzkw6+8MDbbFG
ZNW7qc/jfsPQA67PvZmzC2fcqThbNxePFP20CL5PXUyCtmkCnzW/rQlzk4JeBaao
tGYFkBgJD2wxCMm9ik8AAfWsfIrmOPFwBSXOKs+YM6lVa3Q9czNpeIe1Rfj+GWWU
HxT9qay/Nwba4SgldWwg5HMdYq3IZt/5jztsVzrT3U4+ekPzSp0vXk51J82pRfLD
Rm9VCoW1YAwNLCE9Jb8mT5EYLbAVXovbFDM+K1FKp91phw7FCaFqt9k8riju6ynR
7n2RCX2zA+vxielg2up2/oDybymS7Dkg0WxYNHglGiZn96wo+yLJXKbXrSgxWhpZ
Uy6gUx+PlKrRrEh3cS8qAdecscRC+5SZ/6f28E7xq6T4Gfhfb/7p7P76TMYmIVSH
mqhw7klhJPk52XBDY/6CEQ1hE21t57aIgU71Ibtf8bxTBWTyTCbmjUckWKcAbADD
syP+NMZ7+yApeDb4szU/Gcv5GSqrBYdY8uPeg2A6Ija1srAhl3V9x49tXP+aVoz1
TS+vWflKsI4QciipPG+K5sq6OnKoasQksjidOognL294xlowiF//DuruR7NkyQn4
UbtvCKgtKy/EwLVZFvEA0EusaerOqBzPdGbJQaLXy4htNKgpPICJfTDSpGrrOiUY
vmEO89cSQ7phT04Zfy0DwsGvazex07hBptG6VS7CHQiu+wtt/neLnlBMGtag7ulU
/GufdVRP2HeLyeUPQSuldYk8OSLOrn57IjPK/xobsW2haqy3ijNP2cY9WgmTpdfA
0NP6zXZuCFQ7fVe8yBkevG8suxkbASoBPbtWmNJ9g1A0azTNx0a+St1PgnzqjWEF
+ejT/xP1Yjw/ykkhmYfeNiZlpRpiX4csOpnqqlyUPkRYlcuBt64bukvviLoiWzum
yS8osO9Acf4dhhbfK4Ig2ESUE2AAJAyKvTsvkmL9VGINUhoG6PH0TQveKZWkwqjD
v1rTD3THsCU5oiJMHyX8uVWmEbJ8fSLE9+5j/ODZxbdybbBRJ/6bQjUE4uFXPgUo
jjUSIHKzWzLC1zHfGE+ELXzsDVHZFc3qRj5nTwPYx7VaJoMRfA5UUudA/yu9w8Su
54XdrRd2HqpcR+oGdjrix6+TM5VfUfvXThm3AK5EPCT+0ruludU5q9bXvzDkFssZ
xC7nzCCjS6JiU1c24qc1FTVIpridLStO1TZWJwd+QDPs7ZtEoJxN3BL3KXpOMqfi
JnuPJwIZdxy8DrAyQTdFkcYCk/LZc2UGuVYnw37zS8DsuNXZ2nor7vRcA5yYEVgH
UkN9n3GoXeHEHkgihVeZZajFWDJB3xsUIRtfXAATySzeRlrten397aBBWmtRMLxj
n3sbhnRC2nPPiBF5ibemhVpnoYEWgcUJFBla4EW1oMaZUj4Zu8HP468lSmMyVvgA
GFoe+ncYyoBBd93Ks2ntkZ4aAGd2wBg1KBOOkNqo40SNmp1ZfJF9/YHqAKkyDZOf
egnihJ9spH5jx5ztDpIp+rr3VYzax1Jn8RBBaSfXTGb9KkYFq+W6Q69Caf+OvAIM
6kjbA6L4tacgCUk4jxl4/d5u9RILiEfwMajA0Hl7b83eDoNJBtpjG6BrymGQ7jkl
21ejrAbvdcJ6vCLlMtujDQYsbShfVgIhBuOuCsUDkH5XMrYsvT+By1pqxtaCohHg
gJwH9E6fQ0A9KHgPINfFPsOWboWcWRhVyIKKdZ3jeNeOsGvptrs3IEJifXemvT8u
dqPjWnSIaJseUSlU7Iz9MY+2YbusN7jAtcZJ+aTfXlDpRHnNTpsira+bVp4OZUgw
UBzf4hVC6ophSWIGZLICupXlK8dvC7r5TNEq0LTTB48XiwA5RNIBdC1Ab/6wLLPR
qPv/H7OSaxi3g68k+T6Vcb9QF+iqUUWH4I0Sgmwl+jpHjcznTK19ygUYvB6ISJ9Y
ldqY3QmPsaIIkOl0TCxKo9dKzgcFh1foJ7PeXMPkrUJBa92P1YDkWI9jUPolOykC
MNq2KO1lp+YfuSN3i+mmwae8cvm7LPg0g2KBwOG/wv1sbix9b8fWsdQ6pCmfM8fX
TWOq3t1QDHjIfT/PNCxR0/qxAKUco/o719xfBDrzeo8SxvpDAMnIkle4pWtq7rD+
biTP83ky+8OVaC+hAaMYwNP2cBgAGy+DLDaJtSdPYUF0RRarE2CYgBDtykonwtby
A3AqQyBtYQ7SglUEXhTBbrtG0caVePo9VnGK32okyL058GiExTtINlqnhuF+kM8+
PKqL76bQtoiZvtYfMoCu8FsDmSG/1ZdRRs3dg8p+SPmlajRf7eTI4/Es35rcAyrp
xJHdr/N0xT4bci++ERL2qfXrxCvuEu+PiefsZs44BfDmh2uMszANUdkxAZVznT7m
taynufgNP9tlae9HdfIGv/xNDBL/aaTsUJ3Z6UCBcrgFGLZj5os8pQcvTwWzZaZr
pibx3hZCwR1WxheyOn5ycmYrs2AxJ1y82y0xnqU4IJMqQr53o6nneLsnDyip3xJd
ffy6oSoX19v2qdocM7F98IAGw21QYTOf7fMuIEzpSPf++htXWTshb5eNsWYg/g14
fJRV4Lc5DGLq3qGxvNfejCAIKB+zcNZMlQa9K85y5WxfIei6i30ev0S/K8r3/F9+
jydEtdEvXuLa4pVNVCRGB4Dj0g+pNMEVfALF2FJDFtMgahqw76EBd6nCtgIQR5QT
fpFLeFSdGg4MweTYF+YXeovhWyinEWIvW8dsDEzAA4gM0HaArUwMrIa4z6167nog
OlvLMNT1lnLOhqELgAJ1J+TeohEvy1ItyfNthRFuYcwMnEyJlE4/ZI8ntzL8lbjr
jqtZtq6UeVdyw4HrKpkSTh0wgi6cwPgkDpNPA64+FMa21WdYwxlT8cvGzfbOl4dF
4uS0fNxZYCMTFmYvkCf6P4GpEa7j0atxja67LIDDJgNK/umDnlEa0WJfKoo55zNm
mvR8rQJNga7KqA6/Q8JVaPNgkOanCqwt0vZjwKotihvrhccpEwHUN4ZJWonCDsQ7
mKtG3iv+qc1N6bnUEz8nv8nxgVMwSbZB56OferSRxEr6xbCWLDDVCe53YUPUo6Ss
AbUNWl0XSZk7LSmm8xIQ3NhgpHH4vvcEoO19kOUzc+acT3liAvzpXFfmBsL5O9lL
Y6+QzS0Iff7x29i7+QQYOxelAbJfTOzD73A3SE7ZfKv1wG/utTXg/APlvqWcypK3
dh4yaKgwTrG1YpRR/18wFEpIHwZSO1kdmIkED2H5A0Z81CIvxHa0YAQBv0rw9P+W
W59260EctL7TOy4F8GPDK2Xr/ybyLNXsE/ILCX788sG+T5Elb7yJDUmdTEBVpf6t
oM8PFgFUcVmEN7zXQ/8JxM+z+EcyYi/YxL2cms2oI5dWMrCGi4YMAPWlAkypTqNC
Q0J4WZhgDyjK63imetqxZJe9hNh4u7c2vHpW4SldLKyOOq847tJdZY3CTdBKG/Jb
hsFZLYFnvXU/koC7NyjccAlaWJzHQmtFh8lDj6QFFmRZzioUB8IAGpOuCCiCAQbH
FdOiCHAdFSDmChvV3/2PcTquSOxbTEDQ67XJZ2K0uoPwryZnQqLvwToRsONBv8qU
p09BwXv8nHEKZguKmz45dHivMGkp75qj36KULo0esr4Q95bM6SBfjd4/uDhYviDm
f0Mdq1HanQqsnXgraP1FtJtyWMNfl631ne+rH7e1HSb1F8HKR62t//oK0xYLLl5i
PpBN2yPR5Bl0P67rHxKdK8bI5j6hOIF2x/ICqCRocqE0YHH2cPRnoU0xh1n9/TfQ
kJOCje3jC8YPvhuzOKbn3TZoPFCP4WDE+0CKTPOpT8hjbll4qLKxbpSSGCSbQgqv
siSHqIntmLRtQQylJmcKK5LSSxXM6bmE1h+NfoaadW9uzOa+pE8y2sq/ot1ZoBkg
55Y1VYU32WDsfPLjSVIkz3eLKqJrHYmixhBrU8Oq+PiccvRdgmUIfyIO1UtSk+tb
LrX/toq5G6ri5G8mKybi8TiegYnd748FK/1HzYR79VJshsbfoij+8muxeA9gBqhV
JzI+1vARzcccHMCBScLIzVqVfUW92zEQ5HV55vWI6VcNXYOiYRizD9XA2bPe9FHs
hOhO+zTS/yEbx86/6rrv1vPFvgSfuxwsyV31KbFhdIwcjkUsBZoUFoTRCssVbkvO
HKYbwLsTicYFlIIiAofJxfPn1S7TNbFkuoPhc8S7mrL3dR/b2ASwt7DvEl7+C5Z6
swEf4Yib8hg9yg0hpUL7okXMrWy5ke8iVx5Z1p5+jXPjIuPcfVzdiarz8x78cycH
ug6+eZOKICq/XsJbuN8zkVkvH3yXsuCm8giWwfX4ErWf1sUsuRepo9vx+TtVSBM5
lIE+zdsCVfsDqmgW+i3Z8GPrQZQWMYNJEzgnXv0hCKkN/LsNj+rrjU66l2LqKxZu
kclY6QFpbp4qIjHjyqf+K5Rn6SzIOxW44BvVNX3Tbr7CGlanJ6ENzRKdckG05qz4
Ry2GhxNDiCzHu+SvLV3CJFdsPbP2P4G6LB5u/ErkGQkO0gVVtYG6aqlaeA0bpwXR
frg9l4CB6/WGGr2ph3PKFxZ9s5xoReeC9F9UVVggovgrY6ASwkXf35HjlKOsk1XY
tnjJqOo2o+nqG72phr1pdpBugXSciHpHIl83tzyCiPDtpmUGRIXFg2TCTb3PlFUN
RGsVR1aL4NlcwvTu7lCltP5ClhEGT5bGEPtzLbmHP2vPi2nZagObuLrfZLXw4g9d
T0DF5w8cwcuHQkuNdH8V6O/yHpQbXAxoG+/0Gyj3Gl9Kn8BCJKLd/Y6YZMryPjkj
xdAiXAVw0y+U5+qdNCQH4uN0OwgPtuH0f3r5Vk3gTDbLSiub1v2ockr2WrXBzCLp
0ROsC3+SRmGmXx2/xhxcgul68P3+VPtAsV6MLtsnF+Q+4C5RWv8nYZIr1WVqn30J
PWJR5aT9gFNvxjyl+UmxEC8iqQ0px/uUNhwPCdmLi+CsXWu5RYWL7Pbc0JZmFHJP
hseCVSxgM9cDGBlfZrQdsIt/tTf3YbO38dpmk801uq3YScZBLZoAkOa6HmWk2ak7
dSfyw9HrYtdkBuYL0GxKk/9blvHcvvFsY3P3n9AWr4VChUUrCHcWEqDD/v1DQQiZ
c+z5y5fTB8ltAqCmFWrhSkZROgXZTvFaCdNl5/Cyle+DkJssqBFLac/tfYifAhEu
agkr8I2kdPgQXhX8dcvFCdFs1WzyXfp4yF6iPm/XwGD2/ZiOEGgmmpc+l5i4MXfj
PxBuRcrsi+KeVPl/z9LsqAwHvHzhT1Xothwfwo8uhb5WHxub1p3jWQZgSUIPf7JE
sv8hGIVDg2dnUqUo9Vn/RXO3FHvBJhrgvVsj5c393hu9Pggq9NVAcBcGS4379Vp9
gFdw0mW9zn8iuN9rF0Pj8C8XhsJAHNWRAvKIVcoFKzh9gQx+8mVhMh6NCsljQg3W
wFKC5uvnuo9m23nzcZ0xRv95hVJ4KijN3xUvOoW2cAsw4EdbTTUT2g92A/W2EVfG
IWOSqoSzdRKVNIA6GU5ezEcaB/lrsIcapbj3cRTON5iBd0TpI6S9wepfdbXriPuv
9RXlbFvaWxgvP8/1kGpWYpwmEu0+WsROECxtklPk0lTyPEjfAELwXf0TJFBvocaY
6lGEsnA4bnGRyKz9DViu7O0Q+JjWoa/y0oxjunmC5/guzq/sB0sfrH3mcY4J5jhK
Zhggg4d67JCNMOPFxeIj12lOXO8J9J4K7UpZ3Wm6vafC34FH4vz9xTH+Zyvb7vxx
62+3f84B26WcNXRHb++nLx22zdioq/i/yVWrdKM71VZNBHuRt7lmXz1LxQ7svtYs
hv+lq1uGucL0Rrcw1E4DjNF+e5aicfuK6AGaSZ2YiHppxCvfgzxs7fvxpRzR8vwF
nkHECDeQfTFks28hV01qLDXJAjhb7lpi2MsT6nDlAb2u3F8w7URKq9FfBsruaTZg
vgSUy/ARbMqQTxAeDfKI9ch7OGf8feVoSGc6TMlNfhiZOnUqgC90TCJ81UdhTH9R
/FYA3UMooMgYqkYSb6ogg9y9D8M7Q3vInEoRNE8Ttcah3YCOGFBqIXM2VXgfmBQs
S0uKHeWuZDjUt6LC+PCG+zDaBBROyFAEBuadLah7Rta0Y7A6UNb6xK80trhna5TT
49jLrMMMGl97LgnEOqAurqq+Vq/j+TO1GScM32U84UJQk15/5DQkxGiF838J7989
A6W/8ou4By2QFj3VGigzt2hqPIawc/a65DN2yPw+auuGvNgstOU1TYyu25piIwh9
VPctpvXypjcPyausKgP6w8W4vvnrOEqfiZnNtVs/NkrtgVbQ6NK5sz1YW6pahug+
7CZLhNOcsTiggfZA7DaXm/Bk2L9mmRhkNdubjofIru500vZNIyMfVqywNG1oicvT
cNiTw+5Eb1/WbusPDAPOluqUYUbR8grGIem8jDfkdtYp+fQe2/BnSwsVPFB1Ji+0
AinNyMDZ58EHWcdZXP3qVna+kuhMpYYk7UTv8H80PMxxV7eNf+ejfE78HWkXjK2q
MXOLomSeHx2UuPRdCBSciwHbvid3+jiEgOEmTBaR9pB3Yjywv7moRKQn3PcPRH9H
TqxPpvrdOqY+VWlc0N7fV6z142UHh9chezaJtGcP4WYF9StDiwEtMcFO89rEdhgK
DzqUiPVINxVIunsWgqsNfdLSbVWKjo5xMqjjoJKhEmAjpA4dtvMtJB+Rj487Sn6i
f1FFD5MuDgNTlcs0WXtfQwsCwYyw+3TsgdV0hfo0s/QLjytt5elV2f62FTuxWGqe
n+24QNr8O8dSWRzbspLozdkKyN2upZUUdxUxD/WBQ8Sq07SYg+VsRC161ek/Oa7+
niRFV3Mr6IwBNEa4nF8tdM1UjfLTlo54kY72tx0BCT0hh7R37PXZV1xsPBrHq64T
NZ4i9SkVsDXRMk0WSyeYehd/LPLayl1KmUyhxnNBimxz6JhZmmTNvJxQadx8VSq7
9Bpb3BWWEdmEFhaEeGCP53tAaWlu+0lxh4Ld/dVDy09BBICWn1JP3rzQiw67A58V
aY4xg+JnrOyYmyIt8ZcwhFL9zZNbTVpL5PX4dq+IkXFMnWd1VlHRv4AjjjxSO0H9
iNaduo+NnXRE0/MDbUeX815Rt+C9Cu3NHUYddAvOjY+XXHrqSdwBNfLPTK2BVEtn
wzPsMbmvrbAk8n7ZlO8mphZn0BQJENxWq++/d3tLW9FfMO3avXEju+b8zyHhvRZT
v5Hb1b/B+21lQzN8MLv1MxY+CxqvEGeH9Nymxng3F7ijfhd5JvC3pCwLFA1GZAL+
xfDMi6+e0rE6LDNKGg4mCso0lqmrnUk6zmZIOr+UlOQtgiHIBl278X/6npSzItku
nnG43aV8Yam7hm3A3VbGlYJvg4r0uFUGjC8xSe7S89UHCsPae4Btdvpsx+sOMBBm
H2aOkO52l3wxIYZwCMMutVjzUpWJoti0DtnQwq98DntaGQaqAfaIFvRdzywjdnP9
JeAXAeT+rSYzK2GdJ8VF7FzDJkzRPwZCj2YXNaZTcEEI/tON1WBPJqNy8gN7xMxO
GiIX2YPlTrpCAbhAfrsa8oeVVNxHjPgeeeszr/Cc8rPi3tlsFsToQshO3mrf01Ir
gGYw34zkfnh6pb3sWmQxhJ1rj8NoYuMtvUEZXOHa+Zkzd0UhwpA8vOe4fAv+Tq2o
ZRB3GFhxwILedKjb8PdqB9pw2ZMAxAO+lt/K5ULX/ZYaQYN9xZxHwEJkYjwiHv3t
jEgo9qEG5kxfQTpFIDS8QqGNYgeeNrBSocDJU3CA2W2Q2WhXAr+d2zsNWa077yfL
z2L6vDEjEzDVNFN6nbZ2oKP1d+3TIqh60fNNOg8pztASnhpZgVjEQwB/ohmjGyit
HPofsSn95wZYBtYptPq6jchcjUrFUHyGvrtXI4Onzc1i8oSxNjzEeExjvpTooASo
eGsjc0oAxF+g4LhS6Ah9nXdWrrdq4043dZspOC8lAIRrJNDlrPh7OBxqLgDcV3Oj
tJFATmQvSgCXpL+WVMRGTMjAk+pW7HIW7gJCgUiUKtmM3TlD+DtOsTZGOLFmmcTy
4TY5wpVXVhzg2xY/ixYUPW+aI1KBjl34/fvD/X7Zn1c/GThv8S2qDE3m4lH6DybY
Z4bJZJDsIc1Ai0K14NuwJE33H5v5Tew7WduMyJO3QF6AFuVB5lAdBxlv95jiwSFP
Ts3/eY/+dDXt0AcUjwoHZ/grfAVHv/BSEccUoXnDPQ3vlJQe/Yv7kLjVUu3sq+XH
miwt96Ee4jBVu3PVdvQmS+zlfhq0UQTg3a2aRqFh58jPfaaX1Z9Zessjix1f2m5f
rqVBx9t+B8nNqUNV9cyY2/SPD6fXAvYxKbVRIQ5a/PZKFBNLgEHPfS3pcvY7BjTc
1PYbTLIGrgvYE5QZ5u2mrvVefX+0qp8nS/iaw2vfUJII3Xzq39vemgfg4fkl1CRD
JMM05r3AT7lsYgE+R/4XEDbOIk2Se8EkR7P9rmuEKk5JjXKqMjFOHRJ33MtdLYkT
LlQyP56NVsN2pT4aQ7bp0eLkUuvcNfytUHRI6QfPmkeImvaOSWG/CW5KKevj/5KR
+YYd847pcXA+ywixc7jiRuxOjo5lhUyx9tywYlWZFDfT+nm1y8plcegj3hX4U4zb
OK3uXrTE+NNwRrUPbouyvv8+YR0co8//EOCpVZD0O7U4tIgOUJLEkKt6VIWf8Lnk
J5BvicZ0+WY++lZo8EUZ3l7eyHbvw6Hy6OYp+dJ5aEVg8iqVCxXsV6oWknH463Se
K76rSxaFv5f/JtZtUeKlKJSGr5cTgslypoaSaTkLn0cyvYjwM2JErLxb+LC2FE3Q
Hv5R5W87ZJJbM1t6Y2/DVztqfWud4h1bOg+gqrCWeIZCtPr7ZeffnUvohxodgAjt
WxENQNeGuwhb9aToA9nDuhsEhDM+oBgdiKBwR8sD0BaNoH3z6L2hoqEZ46XlC1Cd
QWOdGg5/7sx2vocTJQh4nXke3sNaC8zEbib+YQ5qV0KDcgTFWmpUlkaI4ImOGFyH
Bu5dYGN4FwTGvOaXgK1d+nHFDovi3udCmIqJqRUHZFLh7VQgVkCJWl/jSvb+lGDI
lVtRRU+grLXuwrAaih4h3V00VpwS6JH3bbZtAv2pW8APHFa5DxgxB0GlBkVZI5Eh
BmWSDlu9997gtay8IO8wWj7aeBdNTPOV2Z9FauBvhLs3HgXEfIAN61cXg4GZSXmL
Bxvj/PFBtjh5ovCK1eod0YthFVDgWQ00tMrl3RzxMAGhlbd/cJCiYgiLkGKsndwR
Lucq0/oKDHAe882gds3UXbZUV8eIA7tGP477AA/BVRauTcZ3j1M0pkzKdsKxviaS
f+IYEiVamRYobhlmcNAxuxZgV77y3RX16hCrvYpQZwwvLAc2aC6KiVx8A2BEaxy0
YsoClZXWvvqvypJOq84GqXlz8xUI4zcUAvXN74cxr8/0asOgPJN86D4AdD+nvo4F
De39A2mysoCbydvJhmFHPFxgwzoRSanPLmwabdUfUn/K4knbbW/dGxKlTQVACbQM
SJh/U8aBORBilOG95mh84wTkv6MKvlE+u3tHj5cuIf78wGEQ2zA1TLUkSXveXa+U
yonPKlj2bzNZADjJ3uEpo48LIz0Bd5BhH0eSG9mTQVVCX0GUwDlaTa8bc2NMeo7G
C7bGyfn22jXCuphCx9qZCYYnUNO8oSnTsHhM7bAj/7a//SN6yF1xbHKK817ZeFOi
Bf+IK2/2/NmwCheCdXItdR2hJqvZftEMkpSw7b/MDq3hWo9QGGJIprxo55zEetrz
GCqz/0LKyEBgXrbjhb1XjBOv8aMFq/1rcPvTvBt7BHiQZX6qroY6mFHXMfnGcYQb
8U64SVeV/TqGhF9VbATx7KA7d60pAsfpvPsdVDUIk5+GKb6P53UxA3hpREGlutLP
KoxURbAwlNuBXwiI2wxeQTAaVGY9Lad+g+KEb9VS6pkWQVp5YupfYljioS4K0zm4
z0npK7XFelvklhwua/OAkP9KH6VOeqtUadxxQnklW8T2v1ItQcunWFbInkgYI3Ce
Q/2Y7on5z/54PMaN16HRl+7QbHHADRVNgTT4HR21SU8aPtZebOY7rE7h5bJLF/Q9
1cJnqfSZdxm83mPJ/yf+H+Q/Xlv2OkOBuxI8tBNaDfzp6/e/nK9PT1KEWlHLoQ+1
9/GJSiYpMVAaREJSb+N/iiKTQcGMR2LfPAN+adiBdPJCNFOqalFNPycnNeMfSgJK
xHtIX3bSgWPMxMQlbLuqCHAnY8pmmh1Nmpr1PdKZYE8ptJWjvBVzZaFIk4Vax3Oh
Cr0Djm2cWvt0zudPy8N4O1GSJcimRPzy3d9o8FKq14MoXqkVhT9dU1oMhfuEKqAY
HM0SQZSs7GHQ3KE0801AWMe1rO3nq2wTfhSNnRM1qqPae6aHZnzUMlatTKRXGm67
SGvJrRY41aYQykx/4UBjZ3WQhIkBGdm/17Y04csYfnsUmszHB01AM4HsK9wMfgbS
jQBVlml8dODTEoUc3PNEp/ipywRlicY+CxSh2WEAls3VJF55BBFtil5qRx2xgVy2
EmUnFGNKdJecBUJbCywRr/ip/cCabgalgNjOtym0DEDmDAuKUtaz8ZDpeXTiKP+T
mHHyuAylLAODopaIgD1TMB4A/nE6ItzhB/U3XQgik+QC/8c7lkSsXcg27MgcUezo
wtaigdmX2yN96zr/3OMY27j8JDiZtVIKrE2Jc6lhs7P7vQ7Lx4aTgZQxtDsxmRxT
fq+rbpOCLNuBI/I7YRmb+CKQfJHlfPAtzVih+fzcF4cq6JbXjyDrzFsfk/ktNqwA
73KCYfNtHD80UalPXlbEEjM8cQSeihLbn0ccMXrtoPD3uCWHP4cSWJteT5weftpf
MnYeZd+oQqBTxAiUrDbLlEkhWekC7AyYCFQ9zbqZIpSYjtKjpw8JCBP1HEKaY65J
C6iX0XcZxo8aXTAcM3pExYhfc0HBSRLdk42lhAHjOse0tZZWxskQLrT9deKeDfqQ
fY07DqQtNelBi2dUkKlR+f8KeuffhEYRmSLMD5v6y9e95YbsLIMyO+SSn14mk8HI
GyfYep2/sPO3VuHFQd12QFpj7mWFsh3sDzZjCBdVKK621ZxdrpO9ZItVCXNOg8h3
oUWaq69/mRrzRlfRempmOjBazLATfCi9NrqBx6IkAzJHOifxbpY6riTGeyJlqoKH
Vvyp71scdfsOARweiwB7adUow4vXfYfEL/cf+DPavWbaUWC2Z4HBB9AXN4HUbVlX
T2cfYPkkSDbNDBpxAMo6H2Hk9so4KfK3WIPcMhGaAApZapfXEDIHqwtlm6Z9818f
AqKDRxMll6uaoTeyP6RfDxfl4/rQVJBXCsnTvvR9tFwm2I4cjzm/RKhl/fO/30e7
pixv42odoW3UKhxQ3QNXalS6hSv0SwcTrvS6d/bQY9lazg7pflU0Rf9kWMUEV2OM
Z959hNMPunY9FXJ3IA5ZxciiM4utwcu32/OwTz+cz1ntlHAcqTjWIn5mEdO/IaW3
h8u/aXri7EsvO6kmVTEObTBOk7+MwqLOJI+sdl2YeMrwXEKF23WB4VP1gfLENYEw
EN3gRZ75Tw8kRhFriEvphKGNLeBsEwe0offaUwJ0YEMz08MboK/BTEB3gFqpQ2Ka
LxkZ3JfTG1975dFM34n46oLTjML/szZoWaVQqeIqhWgQcraO/w5jn9IM9MHzEG/j
kmRR+57IgF5x1gKdX9GAgsvwSvEG/oGpC6tZ7A+zwCwKTTkxE6jh9LE/Ll5DcIBU
Hq69388ydM/OH13OwkhhVhsAc0ymh+gnz7m4o2gAdtqQ0WdOpmBIlPwvULMfQEIL
nUYKLOfmx37aaXlIgc/aKcrNw++rhV5wNIvde7cf9CqhJ3Ai3vXxSUSHDr2fDSjE
5/Ji+FTMR5ZJIva82sQ9zlp65vfFWRZqFsibmgGTKJJkZfKE42vO/yuZqDcFs2UL
F2d8WbZi091EcvibgDVl8zmMOgqUOSaGS2DGf+duHr+11CqF89DZwo5FWhSt3eIW
MQjM6f2xSA8IQTihgdZnBwkrK6az58gwBaL8pE+1w23CPo9tWZ+cMSZRZnEyZJez
JpSql/xybcIbWDSRKiQL2pmSCzu+GcSwRWIPFzWkt/thBFqZVHzbmUUdUdnvO1d/
WwXgcoBk76RfYSUgwNgUAiCd0RS+jrqVhdXSVbBiKmbzNEfU6aWV35GY8uWTq0NU
Gn4rgBXu8BZcrCEjSWGfGwj4l1LoGqwSJFMWjLcpEjFnKEbcVOPiM7+xSSZVDQ9c
Bn/rUgWuPI+lSHMSfm7q7L3XfUe2qf7BXgPeJQKOsiWESgH3WEixtPrOCae6YKX2
57iypfmqEr1MB4MhIKmTfJt6F9AaMhKaonv1WO7Gv7fj89RsT2UrZJOUdRnch4wX
vTfAGGaDpWMI2A1NsvFxFhS6V8QTbIsUmFoXUR2smIOGPaWz+CgYOt1TMsaAdRQ3
4xmNv2oYWi5VyXaQupv33r4Bb0gEC/iyoGchvARgW239XaxnTyDqqvZeUAenfHK0
kbIBtJuR2vnGFuHvV0euts46pvv4LpIBzIBgYFBB3Iv4YBdK1AtcmWW9Vp3kjiMF
aKsJOxeS4yxuJUQ7DmX67hsWkPLT4UoDOM44fOkFND6DQ1xiIenDJXve8ZwvpSqa
qFzqLwu0AVjGKAx99oUtfkdUVH70YRhIZcY82nNTiHESkiTOWFQ/EW2XenC2Bahk
/KWyxHXtbTbRRukUsxLXZKShz9dLgPkloLbEURRepVQKvuo2UUbczoA4rUATRUeA
7XJ0qQV+IQpc692w5iO0QEOnBrns7HwkZbi6Dk34qhb6p2XyJrlwfSm7r/w+6oaH
NpiNzOf5VyYK6+LmdjZOJWN3YgLoyvI2jL9pjy5zHhZWlkfP9wwyYtHcToQS55ht
Xg3ohNo2oisbpopWxekO2bUB6NJRnLDf1Eqk45XzZUBAGXITgiKGnB7+p89yxoC9
ZUlr/u+UPZKLfFQZhFl65Ijs4xnqqiD0ypU6UakKh36gkSKFUgXSH7xJYtoTd8J9
hFmDloO1oVs5ncAzZcizWVnDT6GEbZreAtTl6uaKkYw8IGoF9/cdSMyc7jZ9eaVJ
TwzrXfmy+KNK+9PTqg1qUP03B9PSn0MDQG/vALOOwbu7gsjeawDlmRd3/pNBHpL8
`protect END_PROTECTED
