`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TVh5aaJXQnRW3yYqheQ31C7cQfxlAdHJ8cyMLIxoOXVwkXyFKLZ5k150fomurg2D
LEPLVkABCpl0OK5FddV8UfmBH+DMzEO19ceFuvYZIoAi2HXeKjlxaZtZn+7rzLX4
1G3qQHuJfCF4D0Ct7Qq4DjDyCLW/IBVNxE4OXnYlGeD+MdnRZZvbDOjae8XS0SY/
HffUZXqFAVWVslnl/n6OJmy1K3LNWCwti4wY2anu0So+qBnKSIxPJXY9nF8Lba/b
nIQuDAVBD2MT60wGQj8qyl5jqXsWihWWrXVTJq7d6NWcAvKlHuBN+JKSPEvfHyOZ
7G+oFqVb6b/b0FbJ5HpHimynH6qQY5Toz69+v0imyuDdile3Q8nqLgKOSZmcwvdj
aNnSiIYmrsx5g7c3IFAsnA==
`protect END_PROTECTED
