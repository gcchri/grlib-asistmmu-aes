`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X2SjGCBDUhtNoPWEFy6tZ8xNezU0vNz3wGH+uwRGg2QIS7SB6wkx1vJ+4cefmmNe
BLsCmnsWDZnBYK/aefpcYxo/wby1BUcMypxHrWrQdbj++aFD62Ty0fpMO/WfMmwE
7sy37OS00QHi+dh0duOq+nHh8AscDNznhmH9hMKKgAYBs2DiK667LYZqa8899yrH
MdczID/ZaofJfT/wXWz4C1kPOs0PX0OpnH8IJ1cAp6ufT9VlV4y363CpVr1v77qK
XUl+fwxtBswNXWPR78dduZ/AXU2saqy/L8wZ7eQw6tqA9b1878a4+w4QTWjLFarZ
h0ofk7o9U6EnbCoxfjFa2MvFHnlFnFjzp0W21Kl17K/2Vu+Xe+Pvm3y9RzrCLsx2
4ml65xUO9gYJ/xGgwgB/d9t//pTHIW4WwxotwEA4HOI7fuCbfIaGdu0yHXA4Ac/E
LGQOqoO22Wl3zdbNCLEsVhQOaxn6GATo0CZm2J/v/QLgEQwYB9I29JPwNuOzIt0d
UeUQLt3YOlNo2TFyYcZ2K8SLdD8ZSIReuKOW+aAwFlntLemuaCqxe/1qY7mEY138
e9UGuJJHS7HwLDvMZgpQ7Gesmf3YJIYTKxkR0XofZ6RH2nPjnBb8QdBiLnzgv+pZ
daG6DpKljiLuGCe+tV6w+8cQONobuc3gU7ik88q/eu4TJrCKckGFf3D6nRqtLPFo
buJtO8na6PknMA1/TDv/oW6/cEPIAJ5aSYL3qYau7xToXgHIA8zG9xbPtnFAmpNG
Pj8PXU3dqCfnetbEhIh7cg59I0aeZeEanPjWvYrjbzNFEF75jAilvP+fC56QAs5a
mgTArXaAt07NlnGkDA0AVvE+RPysGmDX6NsrC0rIvIPAfXzv/sPiClyEkG0dcNes
nmeBwmqAA60nEZuxSezCffdIVA2MxFZckzN5lr4Rw8J7IEdQs6OCZTWjjc7Z5VrO
SaJbX5ba6QROnGh8FcyOAzCcJvjOazetdodcFQcRwBarlZtLVNWSy2j6eN76jENE
SRGCvWbJ8pjGn/biAH9w5ub3NeAtT83Iui62IHdDQFhv9IGjkoAaHC9QbL53kD1Z
UTWWK7XFBJ6i8PK2azHZF++tI3Qhx9rYFHAssh6UiIUdvy3SysUkpQVUJti4xapV
8XI6KCjZ6QvcP1JOJ4Xet/R6HILSMqVNCRNDdWLnW2uJrgZw4wNQRnyH4ioIAZ8a
cdLddnUFrRAQMVxo2AOCdvvxs5PX/jcqr17UnXw2ngzwhdjlUNl8IiwJd48xRrVH
J2qAJgnV3YpfsodJFStNWA9SPdyE68RQm4yR5qpCoL58zN8pZR9NaD2CzOPAfHoJ
MMVdqRgB4q86/Wp+Kxc3zwVZ7K40Odl5UTAD75s8SW6ObL/MqtSXk2gGANishW1c
SGkXwSZPZEsekW2bkAEGTQ==
`protect END_PROTECTED
