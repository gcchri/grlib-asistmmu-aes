`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
62NyKCNU8UnpdunKHXmHaNoCzZ/a/kJmnuobuDkYpKiTC6L8SsxQj9rBF6s09O7U
5qiZvmpszv10jIvwRYTjgQuVTE0NFEmbKYjT035Jnsgr3QyUgcblX/NAPjRoYROo
CnbrFIZE02FOGjG9tO/xFTVxvlRZgSuTdlcXUerpDqcz9grkFN413H+mvv4DRpgA
yNEJvkgtEY+aCkRNXZ7KwJB2t/wEXYEl+OsPpdnsSMjzz59q0DnkirJyDjGo2vap
Y3O2cAyRVFTW3udS3+L0dtmk+8tCmNIihQR+++vW9My3vk4HLZLTz39okGhNEi+R
AyljLvJMT2QOvOahabkGvwCPe8r7eNcUilpO094yVb4=
`protect END_PROTECTED
