`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oU6BbwMR4L0BWxKRKO1R9jbRnleq2EhyGmPou8ii7bh+gC3jZZI12p8RyKegoeBo
uqKaz6cniG25yee3Z1HW1ZW24ztn+xJy9wUq5fuajps7Wuf+O2drYxwsTxkHSaKO
NqPmJphgiQP6PhjyLa52bq3s+0Iqs0VxuYQu76BbXKdK6YBcfnujdzy8n2Kcfa4H
Y9vGZG397QNnIEPZw1cw4gw7TCg8DsjBsZun1JNsgXhYVfKZu9p2EFGL/GIDyWrE
B/quMr/eugK3xm1ZuChj4CVcn6loNf+Zex7gFUvoRzekrVGRRg90aswbIjJZdbwa
wJ/3t1ryx0Tpjrm04RmjFcjs1xc2z1eE3Fw3QcXIGgkZEtRTzpeFqRZX2jcnad/9
9fLDzup4oN948FMncF5KwrjEKniKfK1xeu/dWYK2N5lvOOziAgzwkVnXuqH0xTEe
KpVyxFHDbncZ1xK+S8pbY2+nDAFd1/uD1CzNm0rzBDpPAmiJ+OoUQs48lCGwPFa9
GvXnV30vFL40mm9p8I8LfKkbvmUw91vqJbbdMHTUNSiFN3nQt00D5p5GtBsa/cc3
ea8L0AhFW3dtZ5t/Tsvj2Mt1DX1thqWdj6R92pLTodqirlG95G0NpdafHa3wdWNv
bvtwqzmgZVsnZbiTqZkrZWa9VY/VQzfIrPiZLaNTzVriRFuj2tVTCHKquroQWtOS
34sqFl5gEnkR1P4Yp9vN8mIkXYlbIDE8XiNBiHIK7Cdg6W2E5g2r4KwNMTMInYh7
9FaBEqovi/WdHFyij4fxv2dYM6v0VLMVOaxdKNG6HxD/3FNNvTGoXn4kHn4YZndZ
2SQISoV5mj74Dilt3VqKbnoRrJYDp0ZABrL0JPxuTwYNfL5aouDH9Yfj0jvztWNf
TJdCn56QsTAd/HGv/05xrvSKUe0YjIWybraNbHdYlVkBFgW0Vs46J45/zI/kLIkt
VmpwhOdB3Nw41nt+KQkIjZYudJkpQ/Gt8SFiXI+fdzhpaUDcLHRzL0MpQLm+lyjQ
hWeDAXc/Jntp1LaLpiRPKoz+ICfth7yYekJx0SDN+yCox6LPL67nP/gmkHaI/enu
tdxNXOddI+Xv8S9PPODcUHVwFZ2Er8+x0eRIcwM30qA9yqDUniHAmmlblHFdJrRS
KVzPBCn3vGVA9k8hNIvkDbw3XyDNwbZ0BcA+f/OvfGOp2rl8lLEJTMQ9b6SQMpeo
vd5IBEe9CXEU/RvUCIdfhXkWxroPJ6TiQ/qMYF3jviM80GJ6IXNv/PIbCEe7X/6I
LX2uiEF80Hn63SmMNN+f++WeK15IhJRIGQPsYlfYbmMuRno/tWJz8HMFGYt+/dql
BQYe6jMRpfq0whsAFCDjmZ7JycuHERqxXw3IUO1FLkdmvqpbZshO7hdlWW241C+c
7jsLkmntQY64EBM7taSYNk0wWc0hFrvtr6yZvFM/ujfntOSv54Y/JttQy2k1p3Iz
JtXsyIMoxQ/b895PKPBEvqY+baVT4Tead3WRBcwkEcVZDVQq0md5rL5KxaU+5vyc
rwt0Vpi7sQyLYceMJM1Ms3PTvlmumdm+Te/2L+VxhQYNY0Wm8R+rl3onTD/hoMKV
R3HBlK88OCEwaV/OHZ2LE+PUddRxLX5mlEa9frjrX0svkT88g1m5+Bvvjkvyx/YV
sJ2N75LmAJs8rBbK90BmcB5Cyo2Xp5txI3VrPtW0SFBYtnoOt4wa89oG/JffAJ8l
0ruxI6fiYtKg81YCY9ZmzLZnIHm3Agcjjdcb0jh6qOmlu424RLZrvk75Du591EXD
qnSmEU5xhHDaJRyCoFIy4RfrtpfwtDFbeWZGxpw67B1NE/E5ZFoHWONnuV0vYxd3
KIs1bC4j0k43HtyTmzPcf07T5KIrFZOIRm1FT8s6xPDkz/K9sUM+N2hP+bQpX+LN
ZPSiwx+NaEIHHJUGsiIudz7IvSEZqMF4UJH32btv1565aO21P1RN5lWA8umtjTn1
hSFcqw0FRezAw9FpuLkO1qDUgWKNowRdsk9ZOClDZCnFWAvJ/6G1DUZsN/lU/XzT
3mFS5HXjK3o5PSA15K2/8g+zzeeLP/S51q0zED/7S+dRoNJz+gKfmCjwoaFfFPyv
V2Yx2A5PNRplCHm4Hg88HrRbpTQ5UC4E8Ks0SNDuVqxsAKRFcmTAwpOacN5MHKUF
LKAFgWTAChToRqVPCmLQjvCzphc9WnojHWK4Iz49D6KO3imVNRK9D+1AAG0uaOrJ
e3jgCa0cVXeYUMfbGV4tw3SECReEjztMlcQoPiTM+dky2loyEG6sLvFTb4ky3Jzj
n+5D95Lm99OiYOpZBbVFUiHQ1X9BHYOHvokVkFgKIl/MdEgPGyjkscwBjvW+hIAc
Wx5QjX0Qui+4ZZV7AVdj0wd9AC6R3tusG+LSVJWKL7G2IrDehT8Gv5gTwW1PzuSJ
bXhrvCY4yT4JqIq8XkW/SlzX6gG1v2Bauz93i+8eolIsJnL4jqyHYvAXxcyyJCSz
N15g/9abj1lehGDjqe8JHlOZ8MwtzKSfk4hf96OOUNVyhyHywr7ma0RhWBQVWTaI
nStiLjYmAIyxamOzK1bJJjB0aPLuaN1FQvm159ACk4r8nDnk+Foh6zBDidM4Yg4G
++3GExX4r5BMLZUh/dq8jXWRk7mGhsz+zGp8m64QhnhOj3D6APXkGb/2b9ue3utL
dzYfPvBHPrOd28stc+ubK8EUwdzG/DfV+8UlYjMKR962c5QNe8z48eqXGfCNZ92R
47kXe9TV9DBBRde7kshyIyagZaXBcmRKDURqmxFhUI+nRqaKIF9bTP/bq2pMSq2u
aUKoSXqvGny26oYsdJZfKYKwVmaqKSznwmqtAhKydCJwCxeND1jlv1IuskuFKDSd
gw6hjdxA89XSDDt9pFHwZQxZQUhsnVsWEXhj1azC3VkcRdhkGZqxCyPUgN7ZRAeZ
jh0USR+iewyIY7x0HlmGDg==
`protect END_PROTECTED
