`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sjGZ9D5itxZnx3FvWuma6jXGmPFenrarCn/Q6LkRlqhvHpgNQgVOi+U6QDojEfQA
N7mbdA7yhRPhkTqWPEQ9jhecbcyyoifCjt0w8yGQ1MwU7QkzsH181oeLaP3pAGvt
Xnu7qHJ+A6RB/2ABo8qhwTgKvNjxYymcfsG+ZHvXkJcM4QS1dz4iyTjJimfn0krG
lhkytSUKocp66QMGVXwi68YgKWI/uBSyiok6jKQYdxqbFOVWZiffqrU/yGdR6t/h
7/Y2GTqMcxbc8D2ljo2G1WUr+WuWloiD7gveY9vWYaZLp4wQCifcBQDAUB4/KCQC
eX2YbyVpmpRt31zU5LPKG96t+00wlH6vBIZdEyQqSLCdf+FzYPZUUXON1K2jrDjC
d4pSbaBxzvNlexi0uZUkJY25Mh0+Z8803zNmmpH5RZwgP9YYOM1W09LqU225oBSF
gYebUS0cOK+LycL7oucGF6uf/jgKlk+tOdwG83cdP5z/jXUwZlPiF1knh3M7c/Rt
0X9ZhAzlCroM9VyuR7EZ/jrzrb00egIewUGR/QER/C/QC2zcr82REE6Do5WB1yAY
bo4fhbZp8TyYmAiY52H6ydQHSu6nThYeR8UlUMHuj9lPd5WVSoZLOSUrN37V+m18
6RcVexQWHSgP9T/06crNZDfqwuAlxbEFY+Wu72egCWPK4dgjoUgFCBilIb3ya69J
zcNwmRLQXAMqTY+UZPTfQ6oyy2Kxu0jbus9Ri4+fsKrg6VdHh5KUSF1kv6SMLVGh
EuHKPd9kJY+n1tLlkOtkzeGTRQSI7dITFPXUlhQKbnWp/YjBoOQi6l8LO+fBAC9b
8PGJGkmjOzDZBa22uQ4GkDUZRp4dkubiZWCSnV02770NJ+G0UPFEzXMIe9D6VnxP
IauhU6louwmgacUddnsy4fL28ArPfidMyRaoqllIOT0GJx4HMx6Zt3Tgc0+hKFiS
Nw2hpN3AwIxja27UGy5sQuXmIuY3QfTySFND9WvTIUR1baXp3dBbJcinhoS8wOUF
`protect END_PROTECTED
