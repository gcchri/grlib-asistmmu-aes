`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a1T0krwDbklhZizRS52L4CXW4tkZ4kvfafg+GvxAmKFlB8F4EuSFVbsfKrBLopq2
xqrlZ4ml0MltmHxI7WBBW0Zq++BO+b8dn2o8lw2SwJSICOfT6BYFHpBTCdF4rYmY
AW0qWD5PQenpjbhT1RcgVHr7G4T/EDIy+7yyELnxSof6Y0MJble3GFmTQdQiiFjr
jVApvJ8ovmSVdlj92oN7hRPzG/j4oS4kUfcLzij4efEGQHZoFsISylFyV6OrItbO
AfQmT24wllLf79JaTAzmt5eg+WASWLoEz7rI4bAY/MZzcORwppSpxrX3nM92Z09O
n5cGXTZRklz/GRpUcn/cDOn0aK0z9S0w6lewJ9NhaMAhKMoLi13e/EQW/WnjJkhL
ucf4IFykDJ9rqFbx+qP4V4lWk6zgO8GhECvPaqB6lm7lkMAVwcAW5D0AQG5kwAtE
SEsE65q3tVyYP2BszIjqiyZpP6Su5WXgD0b/xhh7ubynm7F8VIi6Qxg6UCxMTcoK
4d7acWj3NWzhOnsQcJhafg==
`protect END_PROTECTED
