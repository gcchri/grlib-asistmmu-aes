`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V8GOqnbXPuRtcUOu9H7QB/3srq/3Wsf9JuKzpibgTaLGXSwldx7feE5UCZqJA9Zz
M9j/ORTgvR7Dzkav/ObZfxG7R3vwf/TP6KDny7HmbfHqL39+DsL0UthSlawAFvcC
wDS1cJa4C7oh9jMQyb0c6F3k9CyQRTwrNYCNPT3pm2/qk+0vnxT3ber/nVDdEi+b
86rjltYmH8f8qj1T9BNWzaW1ubalKzZxraL7zN5fZNRbG9DEsl9aXh0NiEq8JdCU
AiDGAnrNA1ldzUM/ghWfMUFdjXns+OQAVTKBFaPlnXSx4k/DXo0evSCXTvSTTyXE
EIJrVfOm2vS2tFVeKdkUuukUD5gqKzCEs1lAAFt79naEoQNytHwKkTHFf+KYjNsI
rFw47FoQAQZx8mQkAZx+KFW5X9f6e76WPd+gVqXDhVzQ1KhnNxePnuTEcZGfBgjs
p13SQRryx9k3tC+GauRcBsis4m+EVvHEzz4gbCm4o+QKi9L0wfuCYY9fXga2DxjV
`protect END_PROTECTED
