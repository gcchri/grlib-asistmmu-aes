`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SOMtDxzTTiNak5DXLtx4IMkkvHc/OKmkTMTFeDA9YpaTh3gGaLjBJn7/10KXmdx9
UztAmxlJJkS39DGcDr502g0/1AOrDYV52opCehvqwc6FEn8UIoSTg/PDjWYZjuKA
td+EIG2u9/eZGKYItIafpKklYUs2qwthYQGA48UNCoRnQVtzKvm2iGUBO/rhjU1j
/7x4WGGPI7+q2FrTqP7xSv88gXaBWUVPtmT5t/dM+2x8oaf2jC+7Q84IvjJigb6Z
YCeK5Ds/1J0zwoqdV7DH9uX/Ta2JvGH03ammfCOw9k2FEV5DrZaHtSX5U1dHSqPT
snbLGDAkCYPmfgLre6KhNYBjXqluweSpPwNGSxcT8z2iZTYGvep7Gtw+iXDcOUpL
uN16qSgupHsfsS1kIV6euS1JYUcnDJJNPySaqKFVA0fVVUY3LovxqXvPv2+wXb7L
KFMpWCDM3rFmNx21i+mLtaCcJfEZIMui2CWyM+Za1vR5etizRRmK7J1WCD6R5Ro9
STyb5SG3utcj5/YnVr2Ru7PBhecp60qEZN0MBcJBAxi0BkNV4R+K7SVKaIp5bi0l
f6MatSoqy7v8vkL0Dnc4mRp2sYkPAGH9PRsmlvDDEVbVZH4oPrbUtQJFOqm/SEup
8l8u9IqO2Uxlk/lBHsSToUavopuvp6lRdScZ49h72+c=
`protect END_PROTECTED
