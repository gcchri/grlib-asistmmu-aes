`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iY0C6/tu7nNtYC8/brjlCgWz1ahTR51nrjGuE5DNc6BnGSaYHmgMfYu49VBI5fUN
6nvrXztG1tLW4PfEl9IONj+Ci7Qa30eKec6b+H1RqFShcSiU0ixY26NoyvV9n+gH
YMwdx5ErbateDJOB3D3jEFk+yyNC4Ggqf8U37K86h4q3+rNWtt+Ckj++mRbWsstv
Hlv8kUN++INhzeeDnwtqqOxloMD9eRUghtSy5Y0nE5utJ3LMRyDrvKFt4sToUq5j
Snc5Ed41HNGYoJ+iEaKNS6uLFQS70z4Nh6wOkrwZrDU+2QkQUwXqUt0f/vzCXv/r
Mk9Jy7gUqH1D0+BtS7eCDcEmUrNAKgcWmeposAxQcCPMKoD8cxb8ikcyD0PiSkRS
qsfXND1TZpXj3x6lRA87xF0CPOLZGUD51GzvCX70uuxshjzKYoLWVN4yD9tq++8c
Acu6TUoTzhHyNsWyRl6S+9D6EWGRlUyFEdWBUz+C4MmHMrjw1zEUFGklaPttOpgw
jOxSZOFz0EmkLHBGQ6fQjj3rQvtvXeCNaAwqt1qQfiI=
`protect END_PROTECTED
