`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZV6B6rQQK8zSk4L85D86Aoo7I8igb3k4CRcg0ErSCrvpT30uMZHFheooWb8c0/SJ
QeC8s5r/xSn/T809r7k5Mgiu30jT+/Ex2L0agAf7zUz/2bz5rFT4ED7isoNBA8u6
GV+VNHH5WVbo5vJJ31inUUStHcMIW2fubbu9NN6IWKYVmrV13QSjTrnuX1/xLWxQ
JgFAN9e9Bm9cqsJb1+0oiu2humv5neneqG9+H97rFweTBvEhM+1jjvY+tnIWR1Yp
j3kL5b5jFfKoB8LLA50yEkJa0wy1l155TYxVVOGYmhNRNPt04b1Bw/2P7jyWE+xT
mxxRwCwZs8UZpOlnnyihAUxNin3aHwRStUXlsjPTKSxwJbxVyeF3Zzqqa86jHMP9
+Qg725ElWm1QQCZ6NT8MV5yQ1cPfKLp53HU816ViCJedTWj0rqweWu3rQgORtmlJ
MG3VhphZczCQH1lH43+nP8EGuLIh71TbK0BjM3+Qt0VPLBfxb+rT5a5WjcCbcCBp
S2vHrKUhesp6IJliLrjcrR7P2W1I1W03yRjEb6S/Mr2EJCjet80nzSUH5938X1WG
+GR/KKqyRXo0RanA002FDElk3kFINtpb3N2CNHG3lb0IMIyu3cIrrXAXFxCnPwFs
vh+yO7ddDND2zHyNPleDwGhL/YfqhiLVjOAlg+tg84hYAT4tx2tUC29dgKE0rI9r
WKPC5msngE6PbDlbBWoFQg+QK6ogkUiuAm3VwV0Fcu4KH5zMTCKPDa1gAzWjWT9m
igDTRsGyUuRAi/JDMikcbozUrtYaGpV21+h3uIa1SjQx75n8YmBqQe81Ejeb3TIo
reU5lEP9beHHFrydM0Ju5cAbzc6iF69jjmwKx3Q+holx1MKx+Dc0SWczer0oA73Y
wyxyu9lekgU7HD2ZdbIW/J7CulSddraN2Kmmhlrvervv6CTVHgsDOqJiHLF2jSsj
j6cbFTESvl0itCJp4lnRN/N/rK/YFkWZc4zJW1DufqPlBH09jugR6ns2MtvgSCEc
Apj7JsfNaM/sAjxcXzFTdhsBQH9xSLDAJyilUEeTAyEvAlTtNNFFojNYgzqOJcmh
hBoc4+idrAWPNV57ywE5QqKjieLksMdG4JtI1otvzV8ICsXr8XzaULMiMnMAjmW0
Hqzh8M55nd7InsR8b/ZwqyZpXoszhbd7a2d5ksojBa5Ns1K+dc/WmWokZhVrQ2vI
68g+ThL/QiPe6NdjrZcv1Dof7dOgS0ObdQw4JXvRyc8mTrrs1PZN/ycuGJaqMdp1
DD2EN6yfc3EJnRIk5Mx7C+xZ8n5XDNJOIcnTmIw4XcKKZMMSszQAJk4PmVmp50zR
dvM+e56ADxCkNo4JCCdDP4B+4yVPrLbkTMDgCG3r9TQUvJxwb6fa7zNT+5sYZnfU
M06s4S2saxNCWMa6Zm9zM/j4XlOP4NbzXcSQnGGLzoldfzfQCLnY105D9iFrGQYB
HT4YLcdBEHogT4x4dG7I8NnnaohvTNo3BgDIFUxv7K/QuajP3yj2yEzJjspGBRiC
ZBXT+UNBOeFDktNEqR/YWc0LWxFIv1mbjhchy6Xfu4YJIargnr82S+4pxgzEoogZ
`protect END_PROTECTED
