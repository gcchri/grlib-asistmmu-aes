`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JLZt0JJflSTzlhR57fH75HTmOxNneUT7X+htm7bXhQXGkHqhawVzoPFeoZDc12vd
x9B6zGOUoCeIyzNZ1c0yJA3G4jIIxgg/DYIDoBOt9a57C3Yxzsq6MPjVckJROr2h
VBaphlzMaFXa0a5nE+ES3kONDXhgQ+xD1afLfoq5wZu+Cg/q9I7zzKk9QEONtPIF
74DlfsMCgPf/1obYfX68DhIJCVoei01u01RymLOLkyWyzESE2t09JzkjcFxYMb6C
mQOCRLjeBlXlWI1FpxvT9+d4lOI2oAhFQEq9iB6Hb1o=
`protect END_PROTECTED
