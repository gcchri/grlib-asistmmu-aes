`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lEyTOyNRx9zSiH2KBGOVfKfsVvt0uksKFkICcHFnTFwe1oGlLNMPSWepED/kRXeW
xUkg0YV3hoFtqXm1GT8L3N0gxcdVQArmw9/Uc++vp5NAQyM59/hfd8RgaXsFm72z
cPanF6zRF8dBK9TfRV9QDLJEAnsEE9xC8ZuqqA4ZuGd0/osbrckZ54SN985RwjkZ
R9bFGNxrl3huOTdqLX8wijtS7IxQFBU7ETG07dlKHwBT34r8pFcysw9FMTPxX1iq
x2EaB2jZ1h8pq1urG5rTFbTq5aO6vNTFRpLEhOqnt29IKZfpTMI+fnqcnIZGX6N2
WT5qCpjvNbeRvMfY7jhAUl+XLVi1t3osseEOBMVK1OKkwKLBwEv8e6/QOISa8YyB
MN1eCSpIMhcseNZnCmBUT3XatV0qjPdLLXg5iCFCdFXj8pjzDsmtx79QWmppuSkr
`protect END_PROTECTED
