`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GuJ4hWI1apCtunj8esp8yVMRyidwA8uMuXH9/Z/MX2ZMLNcIaPx7btenzEJZs84G
gTvVgfgrOXD3qpjwWz/DCTKvXb1YJj5lBtSsRGjlqGqBFzXnFJzq8mCdkdv0hUTv
E9raOlvY/gAn2JXoU2KxT7ApHahUyAsYzJXcOQHsbzbmK3R1EIEbs5ZnavJ3bbCK
DvOoXH0wIsUjb6D1asvcP9H5O8C91YALV4krSdRvXNyRVTQWHpruWaQkoMQWglIG
e0nRp49/Ux8wQePVow/b7g==
`protect END_PROTECTED
