`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
15LAfy8EJ6YVnhK0k0Xj+sxPiSf4Z9ZQNxKaAPiygBYzBh7j6ihNvhlkY61c/B77
FGpsYk0Gvi3IIvWr2D2sF6LwkruoYnTX5coYdvwrD1jNvMyJvxT6VxTFlnZ9OUEq
jbcr8L87CaMFZeqruTY/PKqn+8g262yEmagvWvWDElD4U9hzqkyLEh3kjZXhTmeC
IdBZbl788AtDVE5GUbw1DHmxYy75x91/q9xq+nNKULdGzhITKr+utnlhwAn4aWjN
V93EJVWFRsXQWX3jyoA73coZ+jO/OUGwVlyhVEMI/qYnCaiY6GhhA2nACS0n4zvu
CQEM3uT0Iq1cVphOaygph1/aqn/CvfkEtB63Bq0UL6GLyUbCTySzbvLahUSxBXTr
liui0orGGbL/kNQd1W7WhqYSu+3Pr7ok/FIAcbZBev+ArsAO88oT6up1UcWhbBxA
Y+K5W2g86iGmSB7cXM9nKMk5Z+wOfau7urgTAzzLjNmJ2SH0hp8HJ/pl3osit8AE
oWXKyIowQswmzKAlHFzUIzxOx90wWQo7i1Ru6xXkYLsczMSAxz4jRryAWHqr/tfK
jjrNee8EBKHdyu7fNCmJ8vYjzFFPBmJ3ckGQgpVULpG9mJNI+Nffe0Za924yW+Ji
K0R/2UhEf29OUvjP1rKZGKDO92lRpciuP2ZEy84s8GOhJ74r/hC8ZshW8mwc5wbk
+BdMa5TDpIS9rWq2uU2bBoYaw+wuxFeEkJX6QDit5wrdU/jtujg4++PCf/mkBkmk
sGPfFdikQOqVy9TS8pQljd9zMonSfc9Pn6sKE3A5YR3gGRykxxQOtBCiKpDZTcj6
G+IIuGvPrpONmrVss6t5GhepbE9FvC509K06PlFe5uxeLAzEXIEAP83r762a+Mgn
mX77sxNhu2QOmVjQFPzq3vDxtgjj1GLzugV1QcEAYvOO9QIBp08P08xuYNyGuZoU
0JO5m23vAdNMl1RvS0nwdUbxxUbBNS1I4DEY1sk+twK98KENiLJRULkfTs58Joyo
unPfDhmgyCDgp9nnBcEYFc3Bkr5fftEmb+IUZQVyJcXcWj25bBPpks0A3khtj/7f
OM7iDjnlg71lrtzk7mknoXYfdvG5UgEUpvq/GrMcWDP35joG029LJVjnXLrAY6Ai
IWFKm68n5n9ceEdsI1mGDAUJJnAsKfzgJT7Kx3M38jM98KH7Q/Jzpfb/eWr4/vT0
U6wjHFoV68DLbQNefdfzj3oAozWZQyLG/qjzWRWpaR+9ifVqLTEvvBB1R+DdZrQO
seoRDcfHYAX7LPsO5SSil7Y6YyLDA7/w6LbqQYjKQhVS2bEyYNdavLKuU4/Gbyj+
XoIfjntAhbcscp3EgtMZHnC1dJaS30xepsnFa5cmS6HU2t5hwx+R8NI6+C1qsYYe
gGa+K07HuNWhm2wbva8R/9cDOmafP/TmpwU+BkbONBetuUImGnDPwS3gLXGjchPM
gw9Jd/o/IPkVcc79pItcCLYD8fzemZAZnGOvN63jOY8i72+LWEsnDHQcANwkHCFA
YlsI6Qhx2DdzJ20mc2muPKa5Q9MO0X0GWsBgA8uolaQmBX2R+qUn4TEa32K9dxZn
0ApfPQmKa1beK3UTqMFGoCGHsjC+WezKvMJaATfDsTnJmBM8pWmYQ2GDA07H5zjj
4rcwkaA02AoE86dFhod5mBWYgkmSa0OZqh8ZvBO6QpJinM6I9tZh4TJY5/09CyEl
1lvdCTaorzhpvVZDPUaH8C9aN4f0nxgYbckKVtdJMay6k//eH/xFJRUAYqehCkuQ
YLWYTcuqU9/9+PdpZB1LA4QdJo+UQxVmIDTuL3Gtz+tQ6kIpCv4S4YAvKBtvA/Gq
3bXWHWt33K+bEiNy7CxV+sN50skbgh4e5iwSEeFb2gfvAg8dNz3FeGBgceodD1Uu
BK8zhgYYABr8/cU7ktW58J1AHtbarPHG9TVtT8U/PzNKetMXtHxmDSUTfiMgQsmq
oPtyqJ/x9izWJ0zC8fDk+R9DYjXAfFxXrs1hXsveoUpZ3MeWSCi63PM8KOqJGJu8
7HXGAVNhAcThdt1JOoaZ0O0znku98kXe8c9+m0sAx09XsXRNOB/UIvSfcZLCoMQU
fBA8DikWcw5qiynHrhFCeZ+Ev5qEuqqfJvXp9Bm4qPgD2lXeGChDXr4AqweDT5Cs
/QYFLRsbCJz/iQPwIsPxxOXNWc6f+9KIg+tVQypd4c94SH0Rw2bNXzt8x/kWugNT
P1UIsIABq6XeLpGWq2YCH14VpOkhaSRAI4pM9u8oAVWVf2t6FYrMoMcNesgKQPWO
+kssaHZrFDSfiOWGKLIwH/W8A6g7JN2HSA7uZ/QiXz7UTM/N6LTokQQ03WYJXAhC
b4ATWbwCzI01ZZYSvjGck/QBSmbEPHEx3ZGZtbzEg+uTbFa0eFmKGhZPRZxVhSkL
Fz8nqBxO2bSUQw9/JlgSuwoe6xn46Uv4Z1UwOJcMhD5PrnRQni0sLWleiLNXPg8+
6eHnkb7ber4bDlodDruO+NuY7lXJrm2Ov/0B3Vqh55I0TGykyGO1ku5zKnbbCjR3
lcmd7SIi3aowCN5roixY6vWablfT7ZW4V7HTc6EX5C69xm4rLFMHzQQ8+K/Uth+e
vP2OiEbVBybfvpL7FIjCPKex4PWstxO0SF85V/yj1aefz99KDhmVwAFQ28pKIn26
qbpZp1YySHBA509CFUdqNyCuCRD9su+VD/IpF49tHEPOjgGNSI0mvJ+Easm+UVeI
cz+AiuZH6xI9WSEkqH2v3dXWn4InJuzXteBt5Lk/tLBcuZcxoywNo4smnk7rOYMi
7iBShq3FufX+o8UgifSx8EGUzrw/h5tzP24WpwY+0fQv6mkHro/o/XlWfXi62KXo
/iU9wCExRTh5Zr4VgkFhyUoLEU19PBhpgV2Km45XXrq6pTt16b/8NjexwKpn9H8P
r+xWP9g6xmQFAGBxn0oVs6rITDilEnCXhTJGSfUCApl2HOkfKBUdMoW/ebRUuKgB
SFJsgKz0FXgeMzhEwGKea8E3bTJrZoAoGxlF0uk6CWjKYg8YgNYECRCHtEOFRN52
GxcvBVgPKoHnpxuk1WVcuX7fUEj8riw12nOsFoRbnUS2e5an5Klw0k0hZGz+tSVh
7/iZIjwRuuRoWDoo3lJ9Cg8IAaa5mnjUAP5W8GwWumWRXleL8zbsYY4BF7Zx9JQf
w9+vovjvTJw2D0mOCuIo49tJDS3dWFt6sJkp5uQT4/knJXqtsqVjI0eaGKAUwgFv
4d3DXy1sw68QCjcKhnnKNXAHNtkU3A1qZ8C07+FWufa4mdyI30zvOnQ4gztsSuc2
ChXnCROY3IKM52i/4eAxGHRQk3NSX4WCTOCqdnZnUx+lP6Z2rg7AzPPsylRd+O7x
jv2PyHLPPOyBRiMFe9EZaQwJuMwdgRoYXZE/LEsESZnDfmx3X7WYwp8FLpEEUdxu
+2oOnzYckJk5UWKcn+Q1Xh4LSpYYKm1oH2L8sXafKOacs+H/hcsAQPru9icSspKp
eeGm9OYv2HEKWM5nz7Rmnn8h/twKWkzW7Z5Gktv6oqK+w5E/z1ZeuZEUKNrMsxNT
UGZxo3TjInJFhfIF1fYxfUVdmscBduxqIF9qSqv6NHzhedfAuCe3eDDCr+nzC7Qx
jhi8dDl+pLY0U+5E7pVM5KZPxfovCbSZx5lkvjy+qLWqVJPqQOJPRVxT/nblJwxk
uZ+3S1URm6FxUxsLOTAxMx07wX04fsHMW/33KmVri9all0HVifShN8VWcD1yAdJk
QZEakge7XHyW6I7SHdwLlBfSksaRhWy/tQUyiaevaX7E0fjkV9oty+mFrbgdqplx
XBHZoTZmcCfMMmL0qV5hLo4aRsv1k6awj3TauNc9AdC836J46EeYesKa2tmuV9mr
jplEGnjKdrVnRGlnVjFgDQexda8nn/FlQfMkZGwW273GUWKxFPKtspF5BFPNM/xw
j+8YHBdg/uEPOttybqHYd0C+yXQEuIDV3aq65jLM8mIWxaUUNE5u9Q16+oZR8QS8
RWl2dlKGaOnhb0MM3z2Pmbp23HHO6bmYFAvxN08nF4LxjAr9PanVxaBS6InoMM0n
EOlMIn2Re1tVuLji9J0hR8rhvRxu8DuUP8Dh7NhmaTkn9ZslQJBlioEQbUz0XdQ8
9OrX2HNZyYwBWwd04a22PExmSNbgJe3iE32ottRJpNsWwJ27xdy7ITtl5wrVljlM
2QBwMkxHDRm471Hoa7bbcURukzgNMn8k6akZMivgf+bQ21tDyDLPJuZIYBvBSi7Y
hGw1SX0xuKi2k39zGoyco1a+e+wf/Y9Ka0DkkLOgJz4LGPoTR4u6LqgvtP+N+9uo
JMZhcEBNVapgwTyFFJRIc8Y1L47ZBC7nq4vtXtRM1iYg0IalO48s8LpUhnzyC0K9
zPf3pMrPBmG7AMkqGSgkuw9b9OUARngeAuiFL7Hw1Q6BrKohP/4xYCEVSWco7bzh
iAZnz3JswOTRaQCU3PIk+lgcqssPlNCisx0ZRdec6Y9aG+Ub53EgQI2Oocf8Fkdx
k6QhXbcGLrE5o5oXLoMMW2s5mf7OuHPKuIsdTgQoUhhQX6G/l+ZkXK7yJ/yWQWgo
uEt/PZddffeSR1lmqkX6d6+ZBfbNBesVEskcPKdFQvTGAk+fqh7jBnD48xlQoYwZ
rUmP3ZfQUOxfbBMHARcz6EpImwVmBIjtaocEXkoXgETEWPwqDawerzru2Ol+rFaK
3QgoU7zGV5xr9CKDLOvlyHYW0r+CnV5W8uGEc6J1za7ZVW9/GT3P74wZthUnTQ6c
rtxfPXr5TFlXpCmWgsLTLacXba9cPYBnRpc5HDj+Zsz8t2G2CjRCkvjrI2+OB0LO
pf88scGdFtNixM7JK5OuxaQB/k+otVD0BHZUJ7xLaDPhAAgUXoWX2Fwsh8VK5TRW
dQm+CSMRedZnIQmCQdpE+KtC9dyfr2bFPP7GSc3I4uovjj29Lg/W/ZzQwR4J7C3A
0EvRL8a8CVBLyd8NxuaFJiFtzEHhmrybQM4hVdNjiak+OVniq0evdWTgSDmNPxBL
dVaqgA3hTdstVP8no3IDo5uIkoeIp55Oe7v1g9GLBkyEHz6gBhWRQS4pDc4SjkId
zyp2c5mzlnIP3/b5X39CXIgI7lO9+NXwYi7wFNP5tk5dXAX5eKY2yLdLBw5u7XS8
pEJnII/iCBDpwqmPQ3LPj534Eqj5QFf8u+3hPZS3KzTDnPgMBZCjjUD34s/TNwEI
gND7N8H4DoI3GxQhLPvtluQbaoCGYEpMQCua+ybmpqVyc/oWrhk8nzCzoaFNkMH0
05tbY3vMhOEr1eGSjt4zsNJza/uVpH5T8YUUw1cDSNyLCY+EpGdpa0bkatMBLSAO
RQhIpUST0uRuZ62bkkpE7zWvD0wK9hhD1AK1Ps6/CTX+2gOp95CU4JcBsVcMDKSn
N1TcOVptOxoOPAQFxlXJ6gzqkv/GWvCoHVKier91r0l0wEqsoH1pf2bGO0x/wOWC
NXHOImZH0DqMrg4uV0+nasGMC5yrNZ2iLRF+YEcK8qEatROooGTgvJorJGVYalmD
AfHz6hGPHM4BZXaNd99obhko6eDlblMAoBw98TLQYJWKpnmjsGfOgYJeIkKCaFB7
beebtyF+ogVrJTkFv/9pqq4cjHx/Y1aSM9oVsxgjZ92+UviVkOTK8d5o7QzgkpB+
tDXmK1wtFz2gybecXFaQTP0puYlTnHXdBaMXmaVu/yc5FImeU6v6JySoMEiSmovI
rk4WtLwXVlFw9lJO234QkNryzgCiPpFvbq1ugMYfgwcA4qGfRZFhk5FT8qIcI0yl
xK6C8LV252AqyNZC1sICNH66y5SqppuG9hWr2nGlrIRM/5VOg7T8He1iG9SiyBfb
eqU5nUyrcJ/3ljVCPjmmRPX6BgVDYx/pmYjN3NVAKEGmQxNKGk37fAn5jmyfS8ou
6nQ++LQCOcGAiTHdFMf/eALOFe/pd4OF0lZ35dRtJC4NjDTPX/4RRNEHJ6MkZqyQ
ukl6Olp6tkVfZk2n+wVBBmt8x0u99+EwekMQaq3hr1TLcNrJgxqdvu2rBivTSdtW
buPzGmEzUKGB5szjkqhtN8Srmo8+SlgsmRvFZeTac4G/giORR4RcWhzi9087Pnkh
fk+8Ppn+r5pJfbikFblnKm4BqUiwB+fS9iyoKUsI4nj1aMy6I8xxfrIkuGcpqmIu
NB4yCk2z7E4ncOcoVopyZiaMrxuA3uoYxfGG0+CJBEEaTxw8oKmwFldoJcFr2oU/
tzdh2swKMtEwYWCEPr2IwYc6O6TQ06Eq63gZK7+SblRU3n99givY34VzqCVPQCf9
dfQ2iSJp3gfhZxVscgyqWBCCcJz2xLAGKo3H86LgXAH4mzDCLpyy1U9eNMNKLHfh
NfQGAqLpTSoSGbyr37mETFQctGOqM/yPrfXFII5r8NSIi435tpJeyaejA4KoT2Q7
rfHmAnqzS6wz9kpoD66zzjl+YjjFvErn6yUDlMIBMcby+yhUBdOvEhWWvLljgO4n
kqepVtPU1IBdOgi9+xaM+8CZN3abPzBW9lVK+vsQsL0ZKhPMvpizQF1yWog8AaMD
pumzYAnKjj8qNUAyFtaTSo8NkkyTi2GnfA6UwhOLeXhDGyGle53OaGCdQ+b2Puqk
Yc3l9H+mgJ/rsfVu4PrG4gz5uCeUpI/R3v7knrrZu21BB5bR2a7KsA2BV4lk7Tk1
H4FSsRUfAUo8y/OQhkMlaILHCGwNOsB96z8aQ+4pEFPCEWv28fNxZ42jyVC5Bha+
VkJyJTCGXg9Rwxhoi7Bnl7ahACsh5twitWd4SvrQpJUdmHmG5gyclGbpaxa/XTLF
6Ok6Pv7CzHqHr61mOB85MKGYTvvMxTSNCv/brKPlFCkNM+clCvGdzxX2X0Ct+/WV
I3CfQ7kYnNF3vACaQtzL8f84xvZ1ex9pq11g/tSUfDNuBKYZK8leOrtB5jPUvAej
+mAJWv/++P0wv8B7Ud9KwBZI5sQYz23LvitcLKaFz2XrulSiaKzCoFBOQ9SNadOy
mgYwh5SGN/VJ6qiSg6iMZwPA3VnMqzgGzX1LzFhU0ry+sUYPWmmEj1sImDEQA3NB
HspZEK143nZekwbEPcOc5w94QqbjVErCY7crDGQRdI+O9e9cH2aDv1zkcR+U1LsJ
6weKjO4/oX3YM5S3mCJ7OOcAjzVpr4VEBNOjjmGIlfGRfWus05aGJ6xeWoN1K0S2
NkD46xHf9HKWKmtD7FChHpDLmYJp8/dXOdwrxmlRneS+nDiC1vvoHTTfE83wWUhK
qGFC68NaKP0/Lpn7WDUMzfpFjsMpuwou60Wbk9zFIQs=
`protect END_PROTECTED
