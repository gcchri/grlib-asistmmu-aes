`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q/zMj0r8DDoM2Hkg//bNBb4RRmM/1C5tNklXsAodqc8Qs6DhOm5avTVVozg/dbu+
FLH9VJN/63m3Qtk/YDWemW6On2fbzpGoNBdOcf/RS6ymUFsxiZuh3ttcPoa2kjHj
C3WSHkGbJlQuNHbLW0Sj43fbo1GyLQex2AaF2ryHidmvP4k1A5mN03y1k2lcNUbG
afyI5wbf/tJp3itDmeQ8uKFZKF29qbnudcfyKZtwD0/QJx7L6xOLGO3zRwfeK4Zo
CwVUp756D/nQ8gM7AbdYw/m0Cj0f1fvKBar6ugukNIb/qUf/BH36tob/WylYsM4W
W0fgovd7stHz4IxbxUKWlzb2azen2P8vOPIqCLR7Dm5E2QdvG2QhsLArfo97HhmW
5uEtwiI+SyTIgZDDvU6AW7CtySuATnnCmSZoK1OGKDrJgFJVGW1vPFZiRoW0QXmG
`protect END_PROTECTED
