`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kH5DfFqHkZeeLZb32Ue3W0VlzAkzCA4iBLnaZ5BUfMg5tLE/iCT1cXf/KqTbfyqO
BSwHtcCrXY4irHxOPYF+b3YzfxrD9s9RU16MRAjWqaem703b6bxQShD3DLpsjYfS
C5MmE0yluZ/eqsGF5pnH42X8Yj3N0OrOsrxdr3vzSERMVWS74fmzk2vsFYFSyn0O
wux+ssYIxdY8WWbOuBkP9yafF4CLTAhnpzctWwDLAFIRcmA4CxraOJd3bQCwBsHc
tuvh6uckO/d4KpVBVg2xUaUcfld1pxFOPLYaakwHJa3/jtLCUj0+/B757vXFaUKV
Y2KRkfSwFMJ4O5lMaT5SWECnJaZeIIc6iwIDoQtnuWo6aMZV6pYVb/JlbZ8z+KrM
/ej45UQzQiL+uiQ4Xwdf2rGMZ2g9qp+8Z9Z+m1ytwnDzZpZQ4gk8AXegVlO1EySf
2E2VEd5UK5pe7roo/6BciYzcNHdTeAhBdLxf/Bpz5G2Gw4MihedSPhRdhLbMa7JA
1b9Zrx+1Bliw11Ankl7hBttGSABMwmkVrYm8hzJsNOrjh7tHv2MNiEfHpXQFnDMd
o3GiBnj5Rjs268QwNG/OG12NNtgr7hOQlhW7wPGPNGNJFHCJ3540y/xnWDWYeagV
rprpW/vqAF+VcxDgQeujF329L8L4+KktopORIpQetOfj+nVlQiIgEEUs20xvUOmd
+q4Wn0N4f1TA6lhJ2oU/gIrWAPVTfM90Jx50euI5/kbVpVJw9Kmu2MMlHLKPTApq
Z1quJGvNSmT/SThLvLMrTEGMgptYv6cLx8MHhlI8mKjJorU5GNEE7k6zGdn+I9d2
r/mbBQ8aFGZAxgZo3aFr8XNVJVhOa9OJCdwxItqG2Vr7Kwcfg2zMjqchzimpFfP8
99XD12VpASrWgTZ+y61vcMaC8Ri/VxP62QSx9RG0n3loinsYV/d8mCnEQq2qWS7T
`protect END_PROTECTED
