`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RNW7yJoYwdLOQZP3cFuYdzkk36TJEPmI/gzkFMd/sU1kLmtHgIEmBKN5+dEbOH2/
FU3fAHj4YtSABr7p+VnGQnNBymZ51RGrstYZs6CgZGvYSyURsaueCZOmB873W7Mr
Mq1VmQEnNJ7pzs25uOFfcV3UNqAkXfqfJb2JFCXK4WHcY/OZvaHFcmNraGfZWZtT
d1ZZGEv+1EGyG5QgdWNmC9NMB2Y4fs3TBsdEr4hAsCDISnHG/Ccy7cc3x+79whM+
JRyVrbqYf0Zg/amQRpNBEKA0jckQI29F7/K59Lw4gnc3WGBanM9a1ckik1ejBGuc
dYLgyeYqxWygcQtlR0kWMEtXQimsO9S3vwVS2fwWU5sCs9Ml+oBhb+uaXaymXZF1
hJJmwb//EZpX1O5eguaCUm6iuXnNf6GWrJkTjcfrNrq3ADkj8wr8JoGmUepttMyy
HTVTS7+Sgjw3KKEtLk0A5w==
`protect END_PROTECTED
