`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EFp92lgIrn02Y7I8x3dsrTZY1bYv5Q0RhFmD6C/x+rgYOPueWYLzoTBKffTp6WtZ
NJCHY9yY+omq1BKsESAOjMZooengU+/W7+65YO38W4lI2BlO0T3LwU/8W7SKkpKb
bgYgt3fTt0A5ylUmVoJ8MOde9etNpoXG2mJNicRPr2XJFbeXdGqnG2xe9twmMzX+
QKYweQ1/oEz/6yTfZRNFAPRUG0K8Bai03Tvmnqp4jcEgRb4CuhWwGRVa0Gl2FPE3
L5Bj/TwVaIPLRnm8jcXL0npRNuubC376W3XB5fbJBPoQ+5/ttNaFZ5RUzqtfyRQe
StkNQzFqc53WuexU6r8F8Q==
`protect END_PROTECTED
