`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K7zu6U20k5yNTKlAoaV1og3cUzLFRXaeh2vybt26n4l9BR/WYuhi84lK5mCYO5ji
89XedJuR+8mdn6Jz/RDHKqaNVKa3WjoMUzzuwTkgpvZhI0q4rSEhogrEblG7viSd
DYoZ6+yACzdlSG+jTgTewO6Pzdex/hxBrp2/0A61snuroCDU4d+PhQPZEObGYSk9
KYrW6ANti0pJ6Ms9vuyBVKRLcW7QYQ20WKR8GvYNg5tXpgKxEXwXYK9sr6One9Kn
pNp262LPZa713/S3w8p5fyXJFUXLi0Z8x7ZOaMqAMSVRfeS74ncL/0fTsrOicGZo
Mjp76NTqPPJpkbHSay6Kv9U3GW5G1PozmBe/ZXPn4BuTCN6W6fLeOFyOzMOxTEAy
`protect END_PROTECTED
