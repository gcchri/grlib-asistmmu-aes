`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i2JZHvkcbIfxezOwr9u/RiMI55Y9A4Y986rdtgmI0HK9uMqpFP0NU7MOkwscWlY5
6J4Q1bt86/GRmUCGfwXqEQzN8ZEkAOEG64yFxgki2C8t+YNm7fVgcoieKeGyW0gW
XchT/qJH9OGQGafMC7TgFpX0/gSRm7zd1b+sAUCZKaKSGnaJnsVSL9SS7M9M32tS
RQ/U0n3XrA1hCLhOKNxYZnhBuJXi7sIBQVG1IY135aV24HGwn1ZpT55p4lo7xp5p
AqsTsww/mQCOkIXc3wbRi6NtZTmoQMFPOCem1BdtCQrLMhQSVMpaGqZrol6YiDAx
P3jb2k84bKnEMezgVg5wMPfQZs2CJzeGmdDYBj4tCiz3/dyF8VIOi+DQWRcr/3xH
G/SBD/y7ydKO9Fb0SQa6jQmVMBaisvon7Fxiu2JWHo8=
`protect END_PROTECTED
