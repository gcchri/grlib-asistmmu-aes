`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sQiIpsODA3/WZXKEVzVgDwS0vhb2eaiAxh0YCDIuyD++4tPH7H9/7QnoMxL+SJsm
eBPwojHsVxM2uW55im1WS8gYeykVV7FAEu5mZ0CVgHAxs1wSP3iqX9wXIoNAUMX7
5aQNU6Y4LNGvHDZ2zoEVehM1gnVp4rOLTmTJgvMivmMwoCImdGZrE6tQ1I+V6+lk
BN7iVkilODQJzXWvBRnaCsCEoZOrEoUSOIw1ii0gyW7+zrqAwmGhwwiH0Qqlcxe0
8gbBlMFhbnAAT3XnyvfgcwvjQgW/vsjWOYBLnxhTbCuDYqfR1egNDwWMpdrVyzCS
VYOp9GIltkqUNxVLr2bB59hYBlZ72kI7W51yM1khcthva58rYrdJ9xjmXBsJQUmr
ZZLQ1aKH1m0jzqUTdO50qR1vSxmXbxdZHnc/Q1dvj5SS7hnD/kiNkuhsQ5iYHAok
G71Q3Cl37iWv4U9InqaFE4JG+/KUQbI8WQr+E/Emp8vzerrkSgq54SguZCIjICQX
CidgXbuXIpoh556QbmGpmNDJ1hI/Jb8/PODSwJu9ygGznSG2XLzuPqcXjrKiCpW9
JeLez40lCh3rbBrb/cZ3/rcTvRjQGb5cTPGB+R2SeUBHzhL0eENWlz676RJKidHp
QVE46OApyZc7eKlMdw47Bqhu6+fowhftZqB0rfKQto7CK02HUytVxPtlJiac0nd7
`protect END_PROTECTED
