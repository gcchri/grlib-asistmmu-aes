`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vdr/tZVQjA8J/ZD90YN4T/32PPWg6P6cMTgAojOsxaOa/b9TFwQj3HnimC86Ojl6
3tZ3nw9KVJ7TlU1gCGzrLBovSf8tMKSGs096vBCITFLdpqjKvc5SHqI82FDX3oge
6+D0vflXwgaJ3L8gVtBrwbIKblrGv0CKp5b/GXPrriNugRypT4bKdZfq+4ueLFra
XVGcGGRooCr/Wdjivz/6W9wYV7z/EByoaMsQe5B1wwH5o/YXjJo0FR7MVJMlJx1c
GiFn2m+zPstpJpfpePZzbm8BwXYWGeFIhW7ozhaSUaJf0Dxoa8JqnScegGXKudqH
eJiCIGEdQh023L63UeU/lrZW6mkid11H4r99vmH5YIAHd99JnIKf8LQdNzdm5fqc
E1ILPEn5VVDrdAbtDFt9jske+XqLeSgB8TyMkzT/vcUyfUz4A554nv1dj0haAQxd
`protect END_PROTECTED
