`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/25iz7hY1hX09OAlW82K+2l1xtWBEVOWJxpDCQ8Q1OrGKanmLpscWIczwa14jCGX
IWASyCoPXg2gWaDIWVhy41Av5INMGlYFJGKhUAZJCHGqb6tibUEllUFKybpiskIu
JPrJ1joh/YPLmPNavdQax+qy0sHgFYz2buV03zW7ef5DP2iX3nn1AizTBic1A5D2
N6ptgvXrZgeEUp96pZqwIJ7vEzkLaM+M0NYiNqmuCEtD3p59dK/VyUrFjM2YdVyM
1te9QbHitFzHN8sHRq8YLIxf1xI6r1EkudnzJqTAtaM=
`protect END_PROTECTED
