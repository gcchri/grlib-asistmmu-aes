`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nymWbspNCFxjP2X45mhkqad25WvtNymj93DuwIwPad+Ywp+aY4kQHqcsKgRbQXGy
ZnLGT1CjU8SbNaGUPvvnLM05wgh27735a98aQCsLZska9R2YzeMZGyATcXCSgWaY
RMjvxyb0shjrrejGidJf+1t0OHaPSjcaKgX2cptsREKPWRZ1LM3OfddFwmIkTLkT
DKyN4hqB2NhqTIqC/Kc5r7a0LpGzrHEtx2YAE1wI7y55h/YEsoLYR4U9y83zzejP
FPSC7oCHsWoGGgu9c7zgnRs3I5bzv1kv1RCzk/w7dJGDl/TDVhGg2ERGqOHdEXAv
`protect END_PROTECTED
