`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hR6p2eluQmYCxdawtvGMn2WJ2lbAYkeMgtAxuc4NWPjwMzZsEdTPmsyuLdqnjS5e
zJTs/jipVflOUevUKqu+Fc4dOb7ZFQjBLJNDCw/r6Zrcwg1BdXgAegyoU83s2aO5
sVS8V4XvUJF5m1dgE28jtQ5ET33QpRXkWlRPkKU2XdvrxTTQrGfK5jtluPmrL8TW
tyHoiqVy5p8AcW/yx6u//jL0C5wpSMvkG5lUEoicZtIXOUjqk+RiLbWOqVoeQzaz
p8qs79lEmJRJryRW0HMw7idbRPt2IQkb1YooE65D640r3CN1IR2Stn+8eb9sY10W
J5N1rrMMaIKVhBoHihC9gu2uHK0LOpHI3BBIFtgHlJ5Y2GAfPlpctzyYNiFskSz6
v99j6cEccLXAD3n91mdZuHDGpRK819e68RiUqxGqf+DgZoHdNWqK+R/6IaPbp+N+
VLORnx94dVBEF8Iu9ZukHzbAw7ZDz4OKXySeUIwi9Dd9bL3oia9vwnLaaYSQwVaH
2orwA3dTXtE+UrWvI47AOFiqwT5QvcD8ItxWgBQc9i9dC2oFMB4qhNIjf9wphbIX
GxNpW+/W04T6m7AR8YC+uUEzHWOGI/iMqk5eerhZVnvD6zcIJIb2IDV/A9vH3fCY
Z9R0OU+Y4R+wzKmd8UouzV0IJQgiznIO0hWz/8Y5TXdXlSZOCxoVSAdQZhUMfHDH
qEE6EBGCj03ugGl5KGVl1+VD86uaeEQYkpC2IEnnn5Ij+0/AeEi7u8BvKa4rb5wg
1RW3hhkPUcFDp1+XBBInzLcTjxxqVszv5uh6R2EPEJdiJH7KDRkSu30MFWsJVZny
rSepGTEo5sY4nv2n22HxOPVjxdeQK6z4y/sOMdy4MASV88LIzxZhauvEDxaNoPbl
Hoj6u4CsVEE0uKlR2fvWFXzqrbRSrs2PuVsc0Khf4ex+onF5O2e4YUndLRd+PDY5
u/EMyFO/RRIzclxyWGNSONZNVQOn1dOs9bFkFmh/n2t8BVkW2C8Mbgd8RScvYG3Z
zhyHVzTzV75vM7AiVtxBan9yWsWvbi7YI+Hs807vDNneS4lav2azv1cPQr6gPS3v
dlZxIGCMzaWaopp5h1yPzeNO7LyMi9yAFHHqDY/u5nVxJqnYAFl2R2PB18KVSGzF
h1YU7nuhV9TqdJ42xy/EtnDXzZeQvpok4LTErrZI5VLonlwS8RGoF9V1npGFwS77
TFDmx2Dk7rjp2HUECaSyILQ77UrdQlE1FgHctGUvXtyB1GMsv8lmF7VM+dryD06P
g30r4EdXdII5RaIP4V8OOh3XEcy3A9Vo0MvcSQ5PXG/HEzxH81AQwT167lO3Oyp4
o6AAf644YOtf+X8DmGTpnMcDkojS/7E0mdtsU8w6x3pnUKDBnX7tPh6LXkyUCci0
4mDfefFNSKpRQUor3LSDpd1MzbS8HvNc+pdJyxlPRYD9ugTT9CYLwiT0Q+KV2PV+
R8iMT6L2EA0xGgZBneA01fw7t4tmH1X6SiL7XLqX47C98Z1uKCEGpoyAQc9BT0I4
emAlL1f3yw3ANe2M2AZZIFlY3yMODQv+C/5gYiiFN6DbJPkIH81m9AfH6yPe5oms
2viUeTxNTxyM9wdvBUtGPKG8FlCwrQeOOHIn3JguW3y2ZtA+a5UQ5avTGqMCMC8h
M/CHpq07nbGt1kTtuxqixcIFf+Us1qPrthOASlM+ipqjvI+Fz0gixPnjR5GvpkMA
+M7N3d91+w8s1H+vA6IN37xZtoxrS5D4REoo2Yzutd1ta3FhbudIb58NqOnIzR3R
mVnuQS6ItTeN0ucV8YVMgGMc/5ixetNH42n+GuRPKwW+uQIjdUuaQFUdDnV8DD0Z
ji4/2ClZ778sSeRQm1Ox9aYTu45P+DN1hmYjujYi/LbUmflHXVpnKI1WwEmc3sbx
alKIYjPlUllczD0s79JkY9pBhT9N96MbL/flLrKMQiwvd1XdwNaNbwUSgIy62bD8
DIIVEaXYACEuwaDyGHZJlF/vsdfDsC2v9Sbb4CzKC35yGxSgkyp/Dgb1+UWhAvdj
uPBemsiUpd+MLY7xUm3HKbnxdqEtdqlDsBdOkJCYeVEDP7huAwGTZdfu2Px2bX4C
45fWGTUPqgg3zlBDL6PCoauyjwVUVBemoUWWx4mYmgg8JJipAuTM2KlJ04DpW3Sg
RH5pB1Tcj2Lz0VJQj5K0TxTNJoe97D65VB+JOvHVcUp73eniMT80rDfERM3re3xi
ZxKiBvEdFjsEk/RBa1oPIWTbGKuV/hOQ7FhTZW7Si3tFsCzgr2oIdUZArOreR6DN
dei+fennSRwodrixd/Eky1E3F61dF9gfICzfxwDln+kY4pRVtSS4hqrlRXHXLt8P
qLsTVOIf1eJKBsWfPEdhQ3GeTf9ha9NmrO7WlNXOQEydBpvKPkeKpd0B0CdUGWQZ
cKw1qI9cpYiS5I7eU7WUOjLuEhPfUV7+x6cO07xe2c7Hhqw2vsU7XXYGvYLfuA2f
pAuMLvkhjiCbLC2AKL3PPxRBvqlxqxDIVgjquWAoLmhKoOYm7TqbYoCWGQUMhPbV
GIJr7GSFxeKjuBdWXpj8N2lLbzaXhY1+eskyrkbfw281fhdeWjO7IBGcStuPe6cD
VAqkDiIbnl5JsDkySReeIFsOAQ0Qqva+/akKWyL/6ig5ygeg05qmCxdBqcttQ9yc
1lqcqtG0cT/XNLZKZWCB3k9c5pY+sT6eNCsSIryXw+5dmWYUIphr8BrpzVJLNGXj
enIWfj0b9wVzG/ew6fhvsmNFCqZMwJNDUljIE9O2SlgOypg43rYtmA2vtB3HIdZx
/K9bFLQPFtZ9Z9Ifu5TWGV1i050i2YLuer3jEea0brVZL2Tr5pNOtGeYeF5gsI/h
ivGN0qyYXBZ+B3Qe8ECteYhb5sjNpiAf4Xr3v6GT9Ds=
`protect END_PROTECTED
