`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cEEzC7C8/wgVSJ5UjqHfBEbdCHev3BXPANdjwA6H8bfvU95fl1odojU/UGvG0Guf
AiuswRTORU/nqJlhH8W5HTCA1OljfHwV74sNhihhyki8kkqmo54tUDFs4JMfDxhw
A8l0c8D3WecYceLq+qJi6wQDw1XdrhF8r0PKO23VmVcl8SknX+q1QjANqN6T6M1q
edX6ztOT7Y2lik6fsS2AZg==
`protect END_PROTECTED
