`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LB4YDTfUDFOz9eXU3zyH6ZRWaB+DohmxPmKHlkcOZXiP179CtAMAS+M5s3S7x8xK
ug3FKBv5nxWQroe5r6MSh7w5kKYa6iB23jwIGyQhMDeYLF1amytabrdpXiBlC4SX
F0qyQUi8tTzovXKP4edHLJ6SK9KI4QvwElp5Y36vZulrRJYI3HaAbha0DHO9ecKM
Ty3AfVFwnXVrllStSrlP2Vs8olEiG/elAtRDwX8K7t+Wdm3S//u59tHFmrXmdmaq
ITc+ZY9bV5H1JrzIfvb8wnwzaLhkqDbNP7YyiSpw+TD5B3UZOSs3ZXXfr9rDsRLs
EoqzMRLNUATRM8V/PSIQQWxImKLlOP9q3rp/prDi5ZJIY1biFf54HO3g66PcUI0M
4I64DHFQeo521md3nyeCjQKmAMOXTE1NKJVd/+XcOUrVdof4AEagNQUEJiVTQCp/
C7EMraKrUstdxX3rvR/V8LMgwcGIzSIrnsSYIWqUg8AsUePNEOu2xssAOofnbXD6
`protect END_PROTECTED
