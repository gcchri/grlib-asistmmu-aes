`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bkKr5s2JID4v+n29keHtxIQBSuicA5u/EhdS5QGAIKg4LvUBtShXDxajgBnmyySy
ozOc0qBiBfAYcSGnp+JL7FvVnEht1kTTXIi7da8So3gzR0cVroUKLGfeP/Zu1yTw
e5xtNogZz1CfI8UYd0NHq/FCgvFbWGxC4CTb1OsuTeYEY2dpPPRDkwDDGOS3Aufz
70DAOPtIGjwKcVKO5poBMedi5Ow/13XJEpU9urQ8QJNAnBMG7ljLa9dd3MexdeIe
DNoPjMYOMbf2k5ubUVBzS7/RSOc1Nk6adOSzFWLLqFjS0/hHZ4EUgFs6KwCzpATD
vXjqKdQ0DAfEC6bS8dBf6Q==
`protect END_PROTECTED
