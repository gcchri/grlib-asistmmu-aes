`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KyxJavfQuJ3nQLCzxBMElepxei71fqYYei+hiziRHH/CS7njvomxCxYlDFY4oTR2
80KZSlEA3bjAK4pfmGLm2hQJpdpS8P6+0iuAlfWQU9ctwTj/x2oy+fA//4uiNwUx
S+yRn4nvK7Xi9ZFcZC9aPj9DMy52evRApo3lkE2SBoRWjp40iXNu1xVSPM0Jmg/s
KmZ0Y+84DdRiku8bpJy4AA9JS6oq1rTaLTHz6JlUKYAxkNIahvEKD9mxTkx7fV6p
PIL0eev9MzSl6iRKKnBY6OMMM+8JwC03io/n/b/x/pFxO6AFTuQs5tHTVmgBRHW/
jk8PRkfZwVc5evMPLfHXoxyC9UQKnOvZBh0FHvdVAWflwGsJOmtOyE3SZ3jc5ojU
fkMagmGXPmzImVPiGrUAXOKvySxjVJVXCeCGMhJUm3gtaKHUz7EJVjnkMESSmrc0
gnQg5TvYlA51D3eEc37lwUd1N4COGe5XOOvUmshlxeWZyZRJFdNjjsW0aoVWKgmG
ooeCxnn2qcoYtU0k0n7jA7YWbCDNGDwatd4P4AtY8Z+IXFvFaugvc2BAsMDHBzLp
60/YpENYUVdlvj9Qcwt3vDbVnxGwYIljs6R1fw+rkiGbHYhNLgXrq5h/GVUSYaek
UnSj1/upp/aOL7AFxm/dcuiDzqp6fdtdGe3wLfYkO2589+acObC6vodHNyvR0rLA
dClUgEWvVDleBwnEXub8pDVd90yd7OGAU0IjdvR2qDFTUKUirAYVqIVds2+5nyDf
t0DZ9SpdgN+GPBnMnUZj8XzTy2bCe6lQwDL5UQQFrYAXhOXBjN9Ly0/Ku/fLKy5U
lR931jCMRr5cqnuH1wxlfV6rVVv0ZeJ7d2ZANvDJhMGgFgoo70CEd0d14zDolGCV
aB5DxANklz7KB+NzhrDykd2x7Ly4RNDXMfXWG0YH5QuE+M7ScBl+AYkR3QC571JR
KpMGkIJYRFl8tJv0chIWta+AIxTTzGUHhD9WnJr8zcal+zkAx5lkASx4CpBdEu/C
iXaIwbOKcrRPTcHk9vq/6qn0sn72FOtPcG3fLHr173zNqLAKTnqvOBflFSbZJEKT
DARSSBcsJ0FEs99l7nnsu9TWvg4c19+G5y0gylvbjh1MXNFUKZaMqSwLXTRUMgw9
89Mgo16ENHwgHXsG7jjg0PHQ8PKA2ajf5FdGBRluNnxv8zOEgJwyRLHY9qcm6cW5
3IUB7vcG3ggRK1wkVZEqVr2xwh82Tua172R2LTpZefLqMRqF1QGK61TqpkkqRtdz
mx6Y7HptxcKdVoqmxbvWBxn5xN0jts95rrJaZGSjcUWQiN8nQivjedqr217gVkiE
fP7yqtJVkmHbYkWWIs+n8bLWbzqTBuvQNAkC2OqIVpBXo9lGHcbIgFnBWU2xEq1T
LwNNJHpOhhNBN3z18BZG7u+S3GhAaJ/6moLWlHrax4Io5+ZgTCAeibrgkMaKCEQm
GhIQMid2clM6vPTWvsFR1B4qjtewzoU4w5fXc9UjXc2Fqra8B8Q1Xewo6mf6fuoW
Ehq6UJu6ew4WbENSMTDnA0MvV4rQgBm8ctyGaLbK5syc0MXg2Pci2tCFMbCjliz0
5kjESx11iyjO9cx449AWzHD7eZZiE4CLY4gumzLNBPHwsikNdNV8ltZU8Szqlow5
MMfsj2E3WoEt1lIe5CT5QxKlGblQW9E3N2qPvB5eHtNMt4ZXed4ZnkdtJrL+a0R5
rUZlw97DbVldZC8id77zMqq0nTphVu6lDVpR+5vqgaHGowB+8wPr5Qd1nzj6X7pt
E47WmScKAHWEnnqKJZstARxK5NABFTpnjf4Wq1g3GMPr26B8y6240otvg7iTQEvr
6fowKyPhFZLkZuwHEo1W7rxir5fjGX5csUIW3DiaRqzZGBMYbBmgnqkX6BWh7KN8
h/1MQeSKWd6LYjtN+RE31TZLfIiNPiG4mPGFEWqgefebF0Kjh9YlYa809iZSENhg
u/ixQMcRzC6AOQeybiklI9d+ViGpi8LE0QuNKBnAEfgndNsQ4MqlUSyrxLLou8Tp
nyuJ2+PbbyyhdKQiP6Xuo/Df/+Wi93M3armmHcn/FgDPy53GOREBTrX+iVOxy5Fl
iuUq6uC8DncLmv/9rmCGElcVA5y7jWBacC83K6PHBAA13E9flZwG7HeXLyfqayYv
HWIVwOAD/yiW4nf3VNm+11ZifCIErQvCQLxzoKYZ82J3ydB4WeRU84w08/5FUhA8
B7bZvmQdSsE1J4PWPByzSaeOAGwcURAt9oPZ58K0N9bkyzcjjEDzBisl1Eb3hqNw
9tb4bIcQMAmzQkP+8TtEYQMp91penNpA8aIS3SJLhG/2Pr5bOx1OAgcJgmgF5gpt
`protect END_PROTECTED
