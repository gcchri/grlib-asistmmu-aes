`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UDthnPmVRwmGGRsAPUEcJecjQyriZgcA5FcdNTXNtYmzBcCe9AmZDtp1EfSTi/Bg
+vtDo1e9FebWjKvT7qZ2Muf21bgcoGR4I1FTRlP3+qbGvi315Ftqpy1RjGi/57gd
DjlEDOhDDVDeknytYtNBK+Tjq0yHJnGgBm5HLfKoMR7kC1Zz71fc2xfEBseZbNH9
vwkHMRvR7C+sClOgoS3UHd8ywDn/31BYu7GB/Gs1Y35IDC/EPRrlNYN0pZcw3nJq
dyvXUkU0F4Fpjgme1d1VstmKGFGCcctbg3YLsfoh++NWUyV4F3DXoiXG2Uw9phwf
fwIpF7O55s/8CjBzm+5Feb4zje8Zxy1rRxKRdiDJz/p+w3TQzU6Dhzmp376pdWkQ
MOJkykpk5FkjWYlCdjwW5/rRWN1otT9RuoyE4OXYUhuu9lAy9apEDqmDXl8V1rw7
hJarsL6A4vNUFi8nMURx9qk3+zCFSyZccw3ZR3pQUIVLDFKUlRD9yGSa+1ujDQkR
meXp4OPFpptVyb2KDSShAKtJOk767R2vMzFa6dYM9fqjRFOEqssBT9TRkMHFnyj3
B0dkpRpawnID1WzrXvDoxTlrAJOtZPEgkPthioNnHyioI1g6iyHF/XvDMerpxKX3
ds5IIe8Dl5VG5YPj6KH1w96f+chveqGagXw5L8XfR6/zqXxSJ4SAvypZF3LH52H0
g4Wl7aqjKCGPdb+y62zR3NDuXOh4L4lClC4ethEhQbKRleYX+976cyU8cswyB4LE
rbqyE6T0KdHe4hP7uqi90LGvPZRBHFKJ8O/UmN8NQneFyu0g8D/ONt7C3sd2AIMA
IpmY0lX+SMZV9BUxqlm0DYUQW8EB6G+KflW/0s9J1l08LsjDjhsdsR4rPh0Ocx3e
/IpuzfWec9RqG9Dif5ODg2FPVkY5VOUOgpWAr1H7KvMhaay3iYg87zB4S85oE69X
HAXc6KIWbcOd32zYpkqzoFAj+Bb96Ogl7TSa/E5jYjszea5wNGsgfjI+raua4EuF
oauB7iBcLR2rt4a5VjYqXRevk1TV5ZcFjRDovcwe5bbjUrvEFSv6aFfO5RTE0SFF
deJVoFGomt0vcfUD3TQt1xVKf1tu7tfEZgBiO0MOyczmw/s0f5VGb2KgP9+ZOclX
zrkohWPxHvzhnLmxG3H+ZdCI/Y7njzZKj5QE7khJ4DKHq3bdSqwptz/GeWl6MqkJ
M56zBbf5gn54uWdMv6dJUJ3/h9brmv1y7FcjYpdMPCuU/oN+xmQMY9qDb6PPAL7M
g1EiTAjyEOOeb0lVAMBeKYWovANG/hAmlPwLPKAyeqxVO9a47lGDNR2Hm0CMYuxm
LJWiejEduHw64SzZ6i3g7Fo7lPV9WmknGySQuks+avKStqtAe0TrOJ2Ypvs8bz2F
jy7olV+0i2Ml4TgXxv4A89+af7JEEB1q/Gw+/4Sk+yV3U/U8hTkXObYUuKgNt5K6
+iVeIXTAwzgFmycq3S43/Mbx+hnfeb0Ls5Tes+cXqQ8IgQXkKIweU2UKh1lZpTml
yvd6V6B+ikcG+6dTWB8wCpzhDVhXIA+kyTBSQNhQGTUVWnbFoxhSWrkUqemQfimp
FJOLQswMCptOhQ3wx5T7SYLmCgZtRNGSFULLT89n8DZp+Y3cWKhnkArZkhCQaJkp
cXAj+KIWaK5q2/TuTnz/5/x3vMnqs0gdIsUZYBncurLPWxSmHSnV6+5F+FhdjPXP
pYGPUZ7BEtwTo/vRw4e4M1HHneKxq+jYiaxpXD8xn2oy1yEIDB0nZ4P8AGooYl0Y
hT4TfGvGIqrI/vNKjfNcPK389qyLgvcxeYfBfd/z3ypvRy0k+zBMiaIYr/QMAzTC
zbTiw8PW9T1EyB8rzCauoXPDt48A6yeZ0yak3dGfeUHyOITFhPFFlR1IfNDHoY83
omzCGypJjQMqE3h4yyjJu35Z2gDusHgk+NNifymeVDJKiNnNAd6g0hHKCQIfcyMs
xD2+57De0z90WXoV1jRwr3ptnhstRBjmfflLypaxnLlKy+LaDpUPAW6Njxeup6KF
EHk6vKDnR+7v/fdsk/HjuFO8OumTmlXdVH8SQbuKFC6wNLdM+JcFAjut+82N23FS
1Lgna3CFlo6zftLOdNIE/+maAoQTBcQIhFY0j6+rs/dCZA++EpLjwfXfPyxNrrwO
tHpAE03H1yc4YF5tPVztu40ajmSAHEcMAm5Ja1i63E/NM57CofQ34Vfsh8aKNlJQ
H16hfaXH9FBlMSE2a7ryGvqyZs/QX1pxB+4+LRVcxMN1rHdJ7yHIdMVzSh6ebaLw
r+50MhBi4BPzxOG2Ulw/dg==
`protect END_PROTECTED
