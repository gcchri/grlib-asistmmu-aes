`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
63lkqyqHhSyGSnxN9g7LIqtcJWl1FdQZG5fljESoxziyqYZ/9T/TR0tq+uM5ul9H
c80WhcJzaYn6OEGNSYPnXX7x2K17xEl5lCthkz/BsDnobM74WZes8mimsoDcT5lm
okYaVZ5h6ReeOmsDiUH94D06NFOfgpw+2RJa58UCMo3p+5+agMjRJ0SSJ1OB3g92
wqVDamlNa7/q5JqBcYkIwyYD2Zudf01m4m6gqrGYYRMIusziC3En7I91bxHBtRmE
C4punfkkVQY8kgN2pmleTH01CMQ6Ko2VTs/XSUwOovW5wZxL0pWvorWt4TmeaJ14
RX5fzK8Trr1HoeEvyPaqxnB63MH73BJ3Qgt89NaRmkpuOcZPSgMXl1iibTpfTF6d
nFxg2RKE7BhpBHy5UnIxClpeBScsNJThrZKVgErd8FfSdKO8UllUgU5PMEi7ZveE
xE17P5HGoyn7DqyPD//fIWuxCcsxgqlFQeuxQnyr3W5gRpAYzQ69CfgOZf/nqwl3
0gu8eIP8CIHkDIxBrdFhXxJoUGMbm9SZLk8J3p1SZdAZ8+7kFIkD24d6RAlioc3K
0xpSTbgSr9U8lR7Inmjz+WeZpEe9sRXsfZ2ScPx3qskT0W/J56+NRqFuG7VZhuqX
ayPhUxt1S31g7WKPtVqcEIQEs/IPc8KtMmsUhRmBmJdtcYpQshV06Yx3nKOeWbFA
4CaDAMDzf00qVgD19I0UrFstmh7FdSXAspeaClKZ/VDNCnOHv/XHSAM43B2wBHC+
YLeY5tDdhicaMucNuexTRZ72CyI5SYVsRLsjI7S7Z0smf3MIgXv9CpkiJHlKcWSa
aafSkC5dmRqnRO0oAosNfocGKMDotXT4ftuUwtjAX0w2X3+9+XdW00I88chTElqA
TokTuXgW9j9F5GN2ChSv+om4sh5Ikh7X6wqz3ZwtmuZ+btBz2ebpi+nzjyOLBuRJ
QeXrWJNlTdctGh0xAfG23ujXnxtCkDhSgTirDZDhBn7WTuude+vsldrfftQtZwXJ
FHunZZLeo8vnmfC+CkJlMz0KZZksAVbnzAdKakIWLX6oYjFeiPDOIS+9cwAZE/KY
Je15M/ecXofZPkrsYFGeTvnTkYKCjiH+vEPFN6QxrFSiL2YwF4rIM1uYK+lVWJ9T
wHg/N70S+++B22CMFsI4780sMK/0EI5vnovNH1xu8pnB8d1Yyxc4GnjlGLxlFmx4
vaDyezlwUQNZJ/O3Zo5dpwm/4bjnZw6sklVqqeHON+nVgqk3ASFWYgkryslSW8/7
`protect END_PROTECTED
