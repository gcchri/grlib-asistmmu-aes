`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HMgjYfH6eA73YslJJdcoU6nqyImb51EXndcMucedpHkudacI5stXRm+OZkSNBmsc
8UQofHfEwXDp7DdPfPXxDoimDVfFQj53kolKdfZd8ubDvq8GZ3C3zjrswlCbKeps
+u6wmcCZzXQ/CMcgALyW9XQmzI/28uhxStm82L/U1QWV9pbUF2OwQrpJuN/2Y66r
8igNhuoMOulf3XVrUkxrj9EHFGO+E8+McOuTDn9AUFjNOJUU7fmG2VYoIaZE6OZF
r07U/oO3BO6MN2JZhvNF455YSqXmWUqp6y+4B0YnG09+B4VgcBCgb/OHCjBEcodM
ioVzJ6l1XeEAygTxEw9bfCLqv3dBvMuUgATMntY2ipJKPVRE0bql7BQltZpRdvZk
Ewy/CBAvLathCPiAG3qtrvTIL0l7BmNdaMlFGi8huy5m8JzKEMXUBcO+frvKXewG
eTuiKJPo9yUEwd+mGWynAjJ79fWNezxvF+niIdJ3hSZjIWNl02OHe3oktIGP1kQU
YtmwRgPbbX9xxCY+ObTOCqAcnjy+i4Wc12E0o8h+hXtFOQW1po/Cbb5rLswLxK3H
wZFDiA1z8m0U3MDwiYqwjlixsVlEohmt07NqNCCFMl69bnWJx14bOVS5e8uhbTQN
WDbpDMNm5OQm1caQqVhoflhykd3JYJggGNX3WpqyIZjf5lj/SfJvp3R9eNWtH+AD
E/2/LuLWNxJIoL+OPaBnhXfKBYTIcguxDRJv2pPIxVAVTfG4p7MV2X0zJv0rAU+S
3cQfSdmefn40yG+wbDqjCHluSmNrsi3OgougINew5mcRqVu/qZWH2rOfOrktmZsV
0TRzer0WXvR2hg44nCyT7QPT5t5e34OaNEM9Z+cBNb+8VTelO5B37lYgDtxMaGnU
qWvvfFCBvXuzqRnaWwJ/aHA24HFT5vP43Z8X74us12Ng8HjY6Yqe+Fy2g1WKGHVo
z7Vc7up0ahmrtfP9KHmvPxUc7wUQszTkuWuJlkxPlZV4W0VqvazE6VwROw1z8YKa
fLWrumNtJrsPeuOWwbA3g9pmXXq/trMws++CwlTZ1elpAXS7ZLMtLhsT2PV+JFdk
0U97pJeN02UJlFvlaSGHAtDjq9jLDETCzxIhz31QcurRP4sAKFBZI31at5M8SdlL
PLsW5k8C8CbPUEH16XGON2sWBdvWzvT2VM7QMVAWzgpGu5Uf/T2PanzpkWY3rJnv
NnQQNnEADjtsv4wvQQ/J0mRba0DOl8HjGjOMiu2Od2obWXf8gD6qW42o63s6Nr+n
NAIOH1fb50fftngKt1apAyaWdvB3iVcolJ9DQAUoGhDDA6vdA5SF7aAIpMYB1k6V
GZkFUAduYRd6/qRH3sUi2UPRXtTCWTtemXh/44DyawOiIabsyZdwhe0Jh7y7fVwo
uHU6491iYHw5zI11W19tDqQQjWjFya8xjXoqQ0lOPF0+ovzD6LrZ7expCbD7bYzc
duoo1I2KMGPabSTWDbOcC8TLQFqs18UOE8+GP9N1Lx3ueUSSOkjSoAlA5Gx/7BLg
ZjmsGl+mE93t2IVRrSS+JmZFsETmvP3EvtRl1jTMvE7HanfUsPoWq9axwiYP51eZ
7iDe//WMacTSaYQt6xc4ihK380fZmHsBUqLug7/VVIXjzdCJwMYkAmAIcqaKo3u8
m+vZ0W39ETOVZmUevDdCGJtHvDu/hE/7oKdH1PSTgJg2C/lyBibOeB4FaCbbgNGg
pqaH7Vscf7hEUILXQFJaXu1UrS4NVZTaMNzTKVT5XuE+00FFygez6rzlCnla4loF
QHGrfqmSHne0YoHpvSB3J7PIoVborcLdd8ZT8bLrYhUsD2J6/ou/CWp0zj39uVsc
3iy+x8r58JbtO3C02OdP8uLEdbGHHEVmLDrvg+jF+2dLBanQy1Z1fLkAYsSa4L/o
rLTsfIS7FD71QOJM3D4xWRe57ElJ1FVhK8Ho19xMzaUVTLFV0ESzXY2cYOzQ00w7
2BPFJWlvpmfZmDkxA+KtPF9D6zRY5RqTtGfEvh7j8baZDBcX+cCJuGXk9qYV9nik
mBFOAX8s7zBDpQvnzv3lenWN/ckBrBymDPeHn7E7s2Y5p5+xIkGPiTPpvlkKqrYF
b7YvylQFUxeDS9mfjcDMJOzQPpmg7z01E7HPOdOR0eXly60j3k6yb2egCm1aAMXQ
QCsBwUR+rlZy+jL/okMgReZ3shGUsDPKJd98IDfQT5FJ46Pt21i4lnPo9YcJCjY3
qmvy7R7qN7b0e8kfC28/DqQpk5/4B8/rmJ7l+FHDDi3lj2ela7OCIiRp31oHk70w
t36W1yhc9bKm24FryUZz+VsBaXWWdvD88Gg4HbF4LaKMLw0QTssFjxmnw/Hp+dbA
UhtK83Tlhy+aADJyTYs8i4FiT2UogIIrg0gg3DkLHPrXtrzBdOnaM/a8YLtG+bkg
L4OBkfwGxE936O7rbVnMPT9qx5PPRZ7xZuSg6fWRo82eOXEXd/ggcYJvX6ZkA8U0
uHAqkeFpyYYWvQcubpjOOReB0gHdt1oaQWvLP7lCGdfFxrGYjIVSAtM2wr3JaO1U
+1ZcGh/WctanvDu8LIdmurDJVg9M5balZ26o/d9XS1FClSllfuRSph3xKifywep7
MLXO7M7Ub8TRO4DWE9ueLz5XXK0D+Wy+eTFgVI+D7MphEFHOADemO0vLW6l+nnBZ
vZsN7UW9cgYMG/4eNhT9dr0y2IqsZpp9I6TGHqp6njFxFLowwEYOvqmxRSUGhZQ8
syFgv8n/AovuPEPBAHK7rquCdXLY4rbGnWO3pz9ptO9eNMvAHX3wRipWbbc0PMWR
DohWn6QPVlhHk58d2OYGfXy7Atud7SKol0bnvbo5Ls7koD1Apkp2E2TgA0q3lKcA
G0cnaRrrafvwy3rdUPDso05z260W51qv72X9ZG9So9QstPK+x9O50gvatNXP0C5O
QMaHX4I6JM4TycUrdkj2lBG/ypEL1y76OJVgJ2SllDQWuouhfIbiCFcwYd/qhLXQ
59lIWFzCUuxDBUudAkFpfdvGmEToGXhoNRKD6xEFkP17UBCs9A1wjPeYWdjMMWfH
Ka3bvNM4qlDw8EHllw2ebpveke7ngrDBD2MIWYN+QUXgf6g5BHdCOR40tQl/S0Gy
528a3uuNHqPfu65CPJxzag==
`protect END_PROTECTED
