`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TJI20GTLxHsxPi9n0Ljobp6FmZzF/gHzVm6+VbLnKOl6gHgUKdBY1nMsxQ9Rq9WZ
/Lv1vpyH65+YPnCwkCV4V/6Ga0JR6Cve5RSQ60UR9llCC1JiJh3XsfLwqyAy9VbI
gzV/UIRCZy8c0Qb54NIpiJwpB2uHzHs6D4cmcTAAFkloY1vBPCqY2VWu3Y5pVk6z
gtimU98iG5LdBGYFMoKSBfBYBV+T9rH/KK2DQjsjVM/EORCijM/tN43GeqnI9ykf
4D7etvdPVojqMPbSznq2NWtJFZFZk7lu0JEH3R2eQAisbJrM/3wfsCIJFJqRKDsV
ZL3dhdzhkPBJuGIaBY1Ym5/UR2F9Nx8CI/VwWYrXmPCuUVcjhKES5I5rL+G6RToU
ZLpXBQjmPFbBDW3J07sAf86TIdv/3KxMcJXlc3oVcfu7x0CvZtxwxLUAWrNASR3p
wciN6scrc7zgPy4YeRy2zR6hIotIKW1q1SfUXFgHNsBmHWls/qbBIs57Br7h3Wwj
j89QGuJduuQTdsBffHDXTmxZfMJEGXMZSN5+Eh/Q+BWkilUVtQ+oehCmrBw0gJcY
y8DL0GQfxqIrwb9Pih44cw==
`protect END_PROTECTED
