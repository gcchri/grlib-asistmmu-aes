`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x1YV6sMKm3PjjwMzQxVxbkWAp2rK4I59N07uNcfjZ4LjwC1XKFZ3LuZu4vTvk5f9
SVhIlSyfUBFK2QTJG0hZFGIC8Z3bcGW/XjLOXBn0WBRmwHWRCEgna0MFhrNxJxxb
fp89mc57g90oeNNAbIfSwnFA/WNPRzZI3ogSsLST++Bm+Hjyv0CAK1QuzvN1RgRr
LFmx9weP3oGGDoav/Gtp9WQE4QbG23zBAUw9il1+VsPuhaPPIPvDcBOL1dY9UZen
Eb8h33eIHZAYIwXvsRkSuA==
`protect END_PROTECTED
