`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HqKUk6a00nprYlWNS2HmNAgz4lTnPi1LUjXitdYTmvzvDE39mU2HvtDBbVUbvNa5
r7iUtqVDh3RrGb8qq2ziqG7PL/PrxBBiZKX0lrNjc8ouH3jlyalcD6c9VSfD4A41
nvrBu9GU49c74PVTb5BjzNAUUXoccYIs/msvV6dTgzzZA45v6TofPMBRrLuqsBTX
M7he2JOVPR31thjPbkgXQA==
`protect END_PROTECTED
