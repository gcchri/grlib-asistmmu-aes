`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OvnKPSeyVpG9eaBvmO4G5UEKUIL0VAxPWgkYZGkAgZPH32p03xarqADoNGc6yMaR
DPk00o/jWRAB5Qq22U5oolD6JUtX3csz1zMjFjquxi5Itg6d/sarnr6V0/hyYYi4
4dsRTpV8daMXl0zyV8h0WUDNA5lqWzS/xUJjtPvNTghRQx6AIbSwyAkVddXR2h4t
uvpsZy2QS8kSzVY2GmAohnolnxhIf5CWa5EfT+W+23gnuJmf4LVZmWB6iaeCnLab
n+RxVj+aCMwuHYLxNuctHAcKmJzKex0e3M3GmK2Jqst85tK7xjsW7kgb177s7DKh
zeFGFsikoON2BIX6h6hkV8IV/8HRfnAQYBEyWzAOrwhgzlCxQTzaH1f2cNSWvZIg
kCtyU9vKnfAbWjHkEuCYf3+BpZVnxwHTqvQog22PWnXSOQcM9H2czT/VjZ7YnmEP
`protect END_PROTECTED
