`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x6leFLibdeAazTDDwGFGxkT18FGt7VsjK63xslHr0lAr+1YNmpeQtsE++xeisP6z
5Cul/07UHGpGRBrRM6tbQIFk8f9x7Q+HImG+W2yhilIHUHx1kdSPbLovinYy3J0t
aRXukxtPB4YKhaSmGOb+Z5Q4y7WNZKax0u2VmnaTu73CgouTlRtld53xQX6rmMRa
+nsG2DzGWYYPZFg9FE1UUCkLLw8yTls9A2gm+A70/J9T+Gu4pD9jRLGeSBOrL93T
nP7Ic3dPXD+B0UeEh4D5niZ1/d2YY7tZAVdqVWFqM09X3fpYFTAdOaoNQRqHIAxu
GPjQxbGPW2pXn5iAIBa2/cAjwzdFxsZMJb6WlJT7vm0t3iz6SfUUZpjV/tTT9LUb
z9k33T8Z2Ow9u0x4uZBq805nByMiMJ/KNBS/JCemzqs=
`protect END_PROTECTED
