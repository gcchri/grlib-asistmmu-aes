`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gxrsdfUyJpQsw0RIxrTQW8J0j29IcrGFGgKhPu3sqIFBQrh4mvTsZOYNe1pdz+RE
HaFcR5c4Xf/h2otpQENJQ9m6MLnvla1RgghTuzw9VJPLHj+/3jv9CnjAFWJ5RCMw
hlxn9DiG0TVAS6ldsXrayXJwaDoy/nkFnEKxCFRYnFu4B08lsE2Adjo9u/tm5Ziu
PY3VqOEq0yfQXlxQglbk1YkpBpMJAiP5pf22xz//Vk95e0MOMC9G0AQ1kC6gB5ud
uEY2uUeg1FlMWQClsyhf8JnwB96plt4pb6aZaUpxwkWesXc2qa+adcGIwVv4/Wmx
DwpnBifWPJ+hGqGJNzYc3rXS11m0ZA87C69H3RAcm9L5/BjXSaXARwWHJcJeK0Ib
v7H+uc/Aq5mR9hu4eON7oFAtMDAIkcko7V8BN2d/T1a5aTq/tgf71/Bu1TXF2cmc
ZRCWSt1CO7C969VlQkENCovyeUDEFidB71+ZDPcG7POhPgazSnj/iktpHIEOTkpc
5EJoN10Q+180WJ6eWSGeom9L7PhYkBC22gDAZ0ZaCZDK6vJJAYDprLnlaFBbrC62
AzxR6cXs5fzEMewml9IuIFBkbnLngLlZQYxRu/p4Z+/lzYeVON8mDGWyt1xi4you
atGouUcTJstK4QmzOS7BEoMRx27TQCXHsTZ4IFUBHc+jRQlWQrNyOdVNyyM+qvWp
J6CttRlcaJGbMz17Pbr0JavKbvLqsTxVp6KYM2kEmkgpdzTNZ8RMhh769E3kSMwR
T8ctdFzZbosRSEeWe6WDhHduxtswhiLj9rE5Oh+M9AYEVv7/m7FL5/RCnhTGhz2N
K8teE/pnxBGgks0NVZYT4ObpEwnQXyUOf3c30LwsKtT7aCL970aXP5AEQCdHbaqb
EPJFUZZGMCJO6FnSng71UjdXud38sP7AuCttL0XbxAzJaPNziZJlR3VrnCJvcfsv
j2VWdplhrcyS91+QMn/yuef1qw8PP6RMCse8ete2OFkqd2THF1fbBYpGOu1MyZV5
v+tBDZfVbmYyPJ+MLeRQjNjUHYBV2MbOiTWisOB+diVTgmS4qJserGgV6wy/uweE
xM++Nbal+Bz3E74YcUs4zk9VxOUxnKorLIgNUn0ktyFn6FrOiWIilPNkoGBAcjQD
FkuEO+lw4bi/+lI8QX/8OptOzjRqbX+i104tUurflT0iO5Glm5Sz5NzbrxXR2227
YMTh+/lhdlFLVL6XJBo9Bc/S60mI/8zV8d0H81IOUlCF1taa1oYHsqLkNDIe/wZt
ug/w45ddY+6tEwQoJfKkFeX+FkEF4jtu1t4DoXojQNAOkWHch1G+/ZRg+b+pYcfQ
gwhiWgsmzuhNHkPg8tWcxfMaYp5IkRFWyZtCM7BwDzTtpYclbe4YQpDBD4nM4S1/
FK7fFgWvGPxbmWEKH2gjVqQeDZ91SEuei++pVgyB5668f+LAYAY6eK7v1HZtHVEb
fwseNU2xKlSPpYjn29OWQsvpbdnRXItT/V6IJo0cWWR39fs88d6FjHHXst4FI1vA
7v6tXei9ZBr89jKT8nIOQaJ3PJXGlXgLxXZIxD50EE7UVlIdEbJoU7OyWyXwZWrz
oxt1aidasxIHbfd66tJDis3KkRNPI/9wcFkdQNAY7GKXQ02q3lDpoeDNkQ2uWNUR
7nLBwms39iJyEu1+UedrVb6HCgrCnS4AsD7kSlmhiIoAo+8aSk9dYQt12neCq+g1
iORZfJOrL4T2i31Yek/XAPcBvgrLFUI8EWt4lq7RppcU3T0lch7BtiN5lZGY/TIL
eAubPjnQIQvb1BlZ/qn/KmjDDH+pQTHDxzeHDnS8wk043kBpxiA+H+4NQMqMpoiY
3NrUzkA2Y6ei+craTNRlf1jrALWgkYCNPl+kfTApGCBr//s+q2tR/nomHbH0QAC+
cd76p9HrP2UppeI+qZ+mU16/pdV1uQAe07IYNP+y3ZUHt7VUbs3mHsG8AeHruNG6
NYes1j1HCL6A76cPgb8f17bFjxSmRS7OJy0iXtmtpEK26p50rnziWrMIsAsHHxHK
MHWuYz6vN5Osy4qiW/7/7TjeY8vILI/N0YqZ80LYu3lihQVpLpP92ml9Sc1Tx31j
EpDFLI7Lbh5WVeZvsyThXmqFNXwp5J+G6OK0oIvI6/3xsleVIqFBVdp+0pqQo+nz
CQi3XZOHeWPBVqzLIVo1Y6S4eAnpFSdNBA7qBip9QIbpfg9gBlwXkJkte8ybFeA0
cFjcPFmcvUKK+mNuycyNSkhNqnem1uTq4zIOEEGCZGB2hgoJ02nT3pyWvPdPzRp8
3WlwEGgc4wvUR2QscB+vqPZJLJFFHS6dh6JiBN5qSuZhhxHVHJHyxXucVE7q8X+R
44ksimbrtflxy6kzP7L+P5bwd2F4+0j++4oxjGOP3RlXUs7+AI6BlDGFXZypy0DN
KvCwvUKagk32gLIbHiO6OfhyeUldgT0/9M34RtPEs/skifJuwQ/aT6Zh2D8epVnd
/FWXUkY2OPVlciSQtKONHDhephP4b02TqvWZkm8rFn0FJ2iycewdZTmmJDuRJeBr
lSxgcE/A1aigxQaXbA5EgdTsl8E809hnr8mQ4e2IglTrel/ZhGtYVTkOlRO5MgfT
lD99ipomKpNH2rQFcwv9/SZLJOxygzrqGQe6dNIlPJCwBvGkutNSKlFocrzUvoA7
49FOOINVi7dR0f14I1rzm+kMQehtszvJuGLCYRbYNeJr65vdQgLS98XlIWzMjHJ+
bd0OzeOZ1Cms4FXIgOa3FLJqxSvsjindhWMUqmhQGuis0EIsR0Ahw7HTIV9OI56w
Ocw80S+b4Of7RjZ7dbapXuU12YdzRmiQKpUlE/wdOCE2cFzWwsHJRadKZaeBo5g7
kj1wZ+l2ejrci04cXbB3CeGHxTro9K8G0jlaoKtGsUcj77vOzO3aH/8gHcnEdXH2
gH018/Y0680myMaD7QFzcWvnRl5OegK0ofPLmS97dkfkXJewxnBc91RSUXPv7P2y
6ll+YlnE2cuTESzlKcSUQnXWF7joa2GCZy2136ssbc8VjJuWmox4bA5IwQHr3pFI
Zmc2ukIse0TDqSMPKGgc8dBHkqpJlb7vhc7aTv4bJ4SXyRv84RP5R7seuZ2Nh7ao
eyvXwXg+LkDzpeNjdWX5EnJNe6CTUCFsF8+DSLhj4fVP5J8TG3X0OwpfRq3mkUuk
m66q/2TlJTazuwmmDEH4sWUR7v6xGaHU5wFCTtldPZnQ3LkQ/t+snyKbb95Cz4bf
a4Tz0M/uDOscs0OAOMU9PpkehQrRHCAOZui9kClXeJxw5q++Ho9kmfKuO+0BveBI
vqkD4HX13ejDxADemF7+vJQRN9rFfK97hr5IBqrhLZ97eaqBFXOk8cFcFBFvKsJo
c1NjmAcoyTzWomK9MKQMe9Xj/va0j8Pa03OOlph7+7GIwmORD8sajTIGvOKfAS6A
EmJwZqDppt5d26Pli7T6ZbUKeysGByKkIboaR0OpSbhLwbcwL+qOtQ4M62S2Eqml
VjMeXcL5RVWjPrYZKp+k7YhP/K/TTNbH81fh0PvHjHnhmaJg8OXhVsR+OADP6idv
VzdsFF6l5VXWi29Ng5iOxLzu1XIlQvklF2mR3KMICJWnnY+32NWhBf2cuqmrDEc+
NoPG/TvNXk4BhwTqI5TOW5ojmlnlK1Z95K6nfRPWFDtcVbDCc7C9IYdNr20ulHUV
dt/RxLIqkrD/h9PBHkljM3QmONwysq0qSjoOrVJTemgZxvjJau/nCpWIt0hIUrA5
hO08XBDGtT2JlAw94WDbvLoh7k9w8jENlP/hZZ/LHSnXZr7CVXbTcebnDIjOsNoE
+5tC/6h9DFMNl97/3dwD2iZ+ALxploEHP7SGhAd7m6oEfZXDw3W5b29HmPBL5K+h
aIQmrPrfXTo3R8VmSHADNnJ6cO6kE+yRid2Et1uk+buDkkLbFGuE3RLEoV8BMOQb
aMUC47w4W6OIHMAuVZUpZyAEMbSMLpOX4iaDqCScfH+oTC4ltGPjh898RF5CypNs
TfK1un44qiyWsXgmb6WYZbKONMZwP56eHNxpLeo8Di2e/sZ/HpKFMHQ4wgEr9HdD
wZF5fZ2CPJbt7OPJVrv7WjSp/e5VWhdo120yejA8wH1FI9ZHBYwIl2Vll3ItzqNn
jVz5Mvee1dmygM4o2SpzvHXuMJ1Dm09H/z4pxAG6N1QWKYNCLi6IfZgjRhUfcRbJ
CXRFyHkdbheHp64kaI55upzeX9vEYyaHF+moYoW9B8mKfL/tSkGVtIjuxa3x3XYF
rxAFDZdLc4YWBtWneyPt47ZJV1DEEsb1XnrL7xO6Lq5t8R0BpVJ5rgK3PMMD36BQ
6xMbhQr0A/obrFpiJxcFHHtRi1iClKpAhaLXU8HksPka670ScDvp2D7sGw5zoCxQ
j7QosPVPmD4lG5J6NaUTDwx1uj5qBrgi+9lJ0Bx5KDRKiQkvF4avBE3yzvEQzrlN
tljKDhf/QjZO/aoADoLJ14xp0nmBNnfOGKP299RFAlAOTutpnW4judZJajBwghVS
9VC7w9RlC6xKbYlHIEkiqJakKuQi7Dc5zsqUOopaZTyUhppKrtX6X8cD1Z7KwAP7
2Amjg7j9/gsvEWjV61uv1bCWKE4l1g6oNZwnhyouPmFZdzAmMN7LBWth02otzKvD
LA13aYuudIK7/ZMz5GXWGp/1MJqkvNcZvgBnfsR9OTzld2EVjRVGv4fmKpwKLW/R
ZjQlxhMXHbYPik0h8kcToiiWKHGx/OTqTPhiAAh8T4UzghmXW4/eM5siFVOARx/h
CaYcJ1qwJbyHWi6zC7KUpe4A+J7fe6BQwZ7M6nSue9+rKcsE0dLOeSFdo3M+a+Bq
QhjuPDsyEJz0MG5J5BzWNeSw2bIPCxhtppM8y4rsWTybMwlpg7qHI9Jn7dDfkSgg
ZI7VPszNnB+49wafgNZMfIFHlwPY1eR8zzSKH+Pr90Ng3rHiFf7inf//FYlM3prA
u7Xv25iLWSHKAQpNu2sUXjD8mO6nBxuLnIHLLau+KvbMafXWOUdw1Mo3+2tgDB7H
WMtXgmOi7R5dElwV5qanezEReliJRYmYh94Ri++NcD/EgsxVusPvKYGaKMva6Srs
GP8gqRgwRBKP2Z7rPD00K6eBIXP0OQ9kvigQFRyvbgUFmboXqhfuFlq3as/qoKHF
mcUlvAA3j/RHHW/3nZ/0YJtsnTEKoWiSoDzLxEyO4O4PIA2qzx7rdRCq+plUsnAl
NIQciiHjcpibkU5W6OAJYXNAILLAAlCTXrZgVN+FaCyGwI5u6HPgbgH1odZpd7ql
sMWZHKTN1CfnHQ83d2dfttXnuoRH4oWgN/RtSoaZkItGWSDgIsh4AaiWc0Nsyil2
re6lGqrjeICv5zVm8uz5wuPI/7lHfis/+0kP92pYYs1CZKZLqGhr5Kwtkj0Gu5tQ
7uTTtPa+KIWRGkYYeTqy/kUVCEKP9gqzuqvwt0YaimoCKk1JMUx5WZUR6mh76Vca
ETS3H0at4VALulx8s0i2D4Z+kWcI6qFR+jgL36CyDb8Szj558p09gtZEG2ELkocC
/PjyVGSs+sLA4MY4c34gkLjSaHIkuEbZ266DfmfdcK4YCgxz2QsMnH55hbRYl8iZ
YYvY3ONrx6jm3916SN2rGqTf5VcbV37WbxTWl+KCKKbZV9bqEKAb8p2XzXTxjemp
Zih5fHFrIFVPRP5HDVLnQXbN2p+UiPKd92yBY3ubM0+3He0hVkkihAEKLYup8nbB
wRMt3uojb/mW0SdQNPmSfxKT10iK4Gg31EPEP1gBhNbMKM9rxDOTAIO0rzatp6lM
1bAOH32t6Vr7EO6DHLyNgGjAqnup4fd/P+6i9l8fgIWp3yShTnaYkKtVkxxNtXrj
dXRC1XbnGRYfY2flaRxhpdYgF22VYiWb3D9wYfUNLoX46JlIvT9S/r4RWKsNUW5j
rwI8/PbAasKxfyqJR/qan2QGW+0jzcdOXIXpSWERtMCbqA2I3uXGy096ufV8xLgW
DJehX1xbHaOnvhLONMC7J/HX2fYxcKd+5LJ2uVFLPoH7uLj10FkjKhLjWs3TfVgn
+17t71bzVMmm7O+k9NuaD90r0yzEoleRDValas5q2NvIDb9qdR0+cMprs6EdVGWS
N141KL8fC81bcsBWyMK7thllHkzACeelqux3oFQsMgdBWG1LbE4DL4SXQLPy5nnS
aiarANLW2VGXAoEYqR+GqRchVQ8O2ZFIKB1Jc7/ULM95X9B9AjocdSKJq2A0X4QZ
B0TmX6pl8r2f4hUwWguMI6v1MvXG3b5qSu7q+UD0vpfjDO5CGedt9bIUbF3w+O/j
ajwCSYNxi0mfULxu4uDptPRw3eeI75K18lo788OwzQneLqT6F3bparLFHIExaMtQ
hOSK6BOOpIRXMWoEz4hvFb5vu1S35QQU56tmlco+kcd8X5LfLvXZ8R1OHiqGQ0+F
taXQVsQ3j8iX9ES3ovuPAUm6pxf/NX/6/p6NYJGfvjepIVQFej6B2PfHTrSf5gMM
GijuJKPzsdl5MkfC/sxIVc9m7EusUp2M0fK7NFYWBaluLA7FW5FFXOpbiybcp1pK
6PPyELu8n7UdyTCBvzlqafLZiey2+rr3Fo2tjgPEPs1+rnLKb7GTQ8YEFWsqzwGa
cynRPVU0b3kWirtt2ORxCm4+CX0f8gUjV9ZcvfayoJQpidCkngDQtf+XFuUYo5cA
lZslu3VEpwuc0C0z5CvNckllhsi9pfJ7JNuGiZlaCQyrKK40cqOkztlpmgB/mF9x
P0ImpbtZjivBMAL/Dg9e2WD42HCjlmw7HqV9XyqGXnKdw5hUeBNCuAJ5tZGynMJB
8CEi/pY9DVN8FJ5co7UHy7DyDpJibdO9uQlCaBg351wC5Kvtpe5hOj+cV0rvcEEc
hZOsYk9dIf7eLDW+h/vTr1FTENciUEx/+3HeVn9iZv45GOIc58FGVGanPR3qcMya
QRSjTzv9l+fCMo2fvKMNGaIzFx+HkbNo1qqJwl6+1h3vNqZ9PlDklTHVnPHpun3Q
NW/iQQSlq9UsLMBb+6w56HkxevC3jpLaiyLZ4Xe29bVXnSaliuOrgrMQ8ha4689i
229DoaAdRyX6f/IayNVOPZFlQ7KPylWAEQ6hdSMgwH10q5ZCtb+OzNJ6pAnj+jLj
1fYC1r/ZbfVX3E7WBPU3Ch4dJ7jhC/h2C599awrVMOWmMs2LBJXZHIkjqKAqV+6C
BlmHuE/0Cn7VJ2Zcm06G/ybHf8qZEj/ZK0nVEf704uVIO0owI/9XmVWVxHHHM0rz
7lyuRNNzU7rpa1EKAk9Hrxl7WZstAwbOacvcD/Z8FqgcBJnofUE97U2BEo/MOoq0
vjRJQ1z0HodrCaVEG57Mtb57QASBkYHM1rUZlc8a4AdOEsxyl26b9IKuWGHAb9+A
gI+oYYA7Q654tQFdcgshPj0gZx08RrOkmDEyiKXmjcYaiuOrOzKn4NIV8hnHMs9h
CtUxghySvj0YQI5fdVP2teJr612DUR2w6bjnF95oo5Rzy9Bk7ja8J6MBw+SNYtWZ
SZ4bPe9OM+T3Av3NraDWjZHq396alvA0yfT22Brr+PcW+0aXa9U0SACQBfLqxITD
5dSDq0BL6A5MhX5Q9JPscsp5AEGXZjGCJrGg9IwreGbPT9ukpsI6X4rsQ13Zlo12
eejeol9g5yA6tHXqeLf7PA1MgBXYB3/q00QIG3u5NW6OENZmmU2AEu1iZjNfwq0J
S9SrS4I40kAZ/AmO890+xsptou+nH7AN2UtCsq52qhLlI8F7EqAv2gIhwGBdqDvT
8MYB9yGjNtB3vr3V1l62ck8Kle90VebeL2f+AXFnTpQQQ3cMFPmEKPzyN+uN1M+6
SIUjy4UMxHfVEtp+CUKyUnbg4PgYauXUl7EfnFrln9eHukICGyU/IkKy35fQb23E
/4uQBmVsPXiFqMo2XtzGVVI0N8uaGEi5IYYyb+415V6mTzhOvN0FvW7Eg8u5qoAV
cHEun5XRTVo/tQ5FATSHCvcpXAgs+U+78McgLNxJdDav3bl6YJx90e+TClUWTAoh
l5k+4s0yHpk29WzgRHfo8AodWrGk4Wuk3cO1ZAlFPmjRW3OVRfbYecbGCVmc5DN2
fLZqOahWON2+uDxnLsIV35IBSm9sVZptQ+Rkr32PRVweumfsqkkxjjdbHz5Bonhc
pecT9JkVasJcuSIesguWc8rJ9kTHRM1gzpLyyA7HuIG5Aweed45fAK3hWxqq/a7c
awgtPNAPFoxuamiLwayBBnjvoislRGzzfSQZsxvzLAKM1fwBt/k3zwJj4+EdAmP5
DQatiVcBmFQbouBRfqAwWYdiYSOBVmuvpyOX/iAbOo7wgI+DISs9c5xKuIBS9VI8
oZn9eeDMs1kOKK47bb3pwm2EqDvvjOkQu+tlbRdg77/NK3UNlirSxmxJAu6SA3d3
OsDiDUAo3QjW328kOvRHNZW448OkJ92Yg1KcB1xtVWynyeuWR/QpADVTZyuNq554
fNjq5HdvOrCq6d9sGYnzMyRfWQGgbquahM+ULvNAdbMZkIsC0E1L6bw595TEHj0e
PIoEv1/RVsKVtqYWReuaXKm/ug5S4qanr/CvyRxxjGYMHsAvt5PbpGOks1if5adD
AqPuA2/NfkCrwE9D/abWiEOwVdPT52hjFJOqu0ja85wWzHUpmq8JTeQjfnkjAFsa
hWpUBQaItpS7u1cZCps7D6vxtW6lA5t3zPvCjkx3xCtJ81E5adp0byA2muv8vDNW
VfV7ZEPRs93PUhyfuvUxdujBDqH+wzj+Bs1ERxgkiihFIHpgf+F9PTHdIzR1T4bw
uXHnIC+VLI8cnLGpA8vWUyto3pjhiOw8AGihDf9iw+jMEgOALrxPeOonaiEeNVc1
htg9TExcnWNxXbMeqI1BvD3Tr6V2f1nB5KEw/UGtcO53J+knLrwferQ/1aPLRSDX
nmJVdEaX0RQ1Kzc4MzN+EPNT68HdSM9vP+hqCb69v94hVlkxVblveTRZb3YmSkjp
s3AQKqqcgFY3io7cJgKabWQA7kgOyLiHNuG8oZCapUaCh+nDvYWbv8xozQUKvPfx
JjTfMiL6DCSJNQ26BqtIGWhMXDlEE5RabcGQzsBJDeRg+tnBL8eYogSRVT/9qomd
ZyUD8EZis7tnPNmlPtJpCWUYWhoRILU2yvZtIA/AEuZaMfWf7fzsvITHpQ9ZAtUZ
jJE2pWaozqTrXRaMzwrrxUKNL+qKJshZxYSlhTdrbgKVkgLUqWP0rUAHqsDjVtCt
RyDmnNYfSHIkzjEYJ5rrCvOdTR3sN2u950ED1HNsDDHOFeAbEkCVuYhz6CgFKlim
dozF6WAPR9Hh5C+78QgMxH4C3sTxBsjiPrL7FRRy6gGxdlv/FAmC27f8wplU9axF
SKkTqexWzwn0qobEcJtRyoYs4RoJp9tk2hdpJN5XU1RS88BLVqCVIulq1/82xigZ
80OZSZUlQyF7WtmzBf9jpuVOztPFkLa0hqbA/BaHEfMvXEyfZHBydB0TSF5fe2SK
LU0lFQnN0MyPEZDA+RVRKEp+0dHFbg1VCoQk1f3Y/a6d0HaYBohc8VT8cNdHmnO1
iEbqz6nbRXq6U161POMIoSuSw/tbm27WcNZiDn8eqfp+tKyElftJymrYMvvztSJq
hw+NpGJn993mWcsXiOMrlXFOz+NT5f89TbZvWcDlKmDeIdwEc/BalqO7pRH5wZJI
747wZegMGfaKdVK58ZI39JSpDiSCSpRKT3ftQXKQPf669YskSaWl6xfXgJ/lzgs3
Dstfyt7RbJ0YSgwPkTi9mdwEfvQzL/Ka6Iv3yKI5bOEjEPg0M/N8LA1EsUmqu0Hc
CtzIZFqbQlcN9a7VydkQMJQb1G5AZUTVC88LgRmrwZJ0TYe1pFbcnrF+fe5CAbI/
afxNrpYqv5+XjLbyvnRQ119DwcrSB3ZDLJxiXKpIlHfYah9tHBFFfg6nFokoaITu
HodU0+01PZWl/ZxBmqvgLYVCsNV3cWSD3Jx4W8xxbKIeoCZ/uYlWikdvDqqSG4Zb
0V3SrYi5Gl7ssBT+VpWGcDyp4JwRSXVNh1gaB4EhnoFvndOS3fPCVk7+ARiEI0BG
CUvoqZS7gqyeYgBYSR0R6Kj4eu2ArPB/WhdEWEuJ8g09WOMqFl351mJR9DtUCom/
HLC+8ujTL5UEs6KDra+TRabawHUu17sV6sSzTXVed7f/r5ePT9Q7uPz6CMmzI4d1
OdnbSoiHUTU4MCxNG54DDDmh1cX6Gvp7iWtntnRt6VH/Jlbw6CL69rQH+inhAXa4
NqM7BoJOSppDMKF9joddr++kFU8aKmlq5BzjNdiDwHR6SfCt7SPABGKl/Qk6gS3z
dqvBmKnLo2i/NJyJwGiazhXYA6jnPrYZ7pf3Vnlta6434G1qYR+blpQ5Bb6uY+zu
5D7ZSJpLzf0Dw8TU74TloesUnp84zmJ9rmBU0s7SweZweb4c6+qO08O4YzQUNy3q
hSZbtRYswH1pVc9YQ3iO7MUSK4S3m3uIGt7rfTSWCB+NXXIW8Qxmh0r//Kn2WIht
FR4hYIAoStZ9LCI4fmIi2jUOkMYs20fAtDhpsSweXXKoEdrz3Uy1pOOshRf1QH9I
IhEHuhnELumxw0gGUP3JhoIZ6yw4bGLpEMlGQXEUyIQgSfs61jr7Nl+nNxPOFvyq
tthU3STMynCI2kDeYynbms8enGsFyEQG/YOp4X3SeDZyN6zZF4PUZwjLjPCwg+gY
ADdJYOccL9wbqNO90A3dJ0X4NMXTnnRiwrYkFLG8i3N10ZFVMBbkg9cd9k5Nc91B
rNUi2U4JiKktRmnBizmL3OqIqeisUKr/78aG15DsARj5ZrDqt9p3SpWUPKuwujht
J13ouf0Z7eQGmaFHBZg5UehM2Op1X1ej5ka5bBVtvs56jyAvDTjxF2DyxMcfiaiY
uuMjSjaWvmBYQ7jjYDx1zz4LIPChHxBT4CYSmAQRHEtl7VdRKRVqP3hSUtxNXmNH
oEOb0TuHFnyWVm6TnPuraFfIVauFs4GtMScG1XrAkyiiA5YzTxVWavjU2IYg7SBC
vFi20k+K4Q1VOcgkSk6LtAXiYfAyCyNgOqHna8CEo1TnuLXbCDi96pmgYY1NPkgM
js1VNbVz/v83Q99mQbIaTTs3VL/7bgTfqm8hqklKuAmiTOFxDEbHFsH8uG8xgf5g
IABdpiqPYb+1RkhsCicB8R72paHWujJ09aUzGpTPR9a3WBUlt/h3g5xhpQvrcBst
bC0R8yjhgG9+FwPUIeE2ph3J6B1zKOgHTk3Zsb0ANGf2zxXGiCqdYWzDOL1q3xxW
rYkuu0Nu5qNX3n76M2P8NWtaAJa3SFsRxraHLyI4vCr7HlAR9LbOR8mu+IohWJsW
EokQ/biTu95zKGzWAL/w8/Co6I8e57rgrtqRrHDVZvv2pyDZFXtnBTwEYfiZowzA
cHoR8fQ7USISloNM2JmEH6dmhuah0xPGsfTFEE/nadKcdID3MswVnKDXbuCOydPW
1TmCHKjgWGceD6xfh2gJ9nDi5s+3/XB/s/Zb0J46evGPBdieXsPmYv1MMN9hxuKN
lamZ0Kb0TAYT8TO82VlfNOMtCmTpIEsc8SSF3Q9XLKzeHVJ12/nXLBqYx896DwGX
qHfo3wUZ0O4Wpc5/OxPNlbRZ7SPLdt1HHW/mKiKqM6lRxaehKXCMJMncbVW9HYdM
eTEgBrcRY3Esi/1sZRxDqtZAHAHbZMSDD7R6KKUf5iDa/fwaq0byahlg04U3id1z
Jq0Sn/qHrx5M05RIwAHDHEIJdNzy2oxDGQ27Ox/PvjL6Xfb6EjOuuLqboGewtMCQ
akt01z3idfkfvXcO3BNMJZo7ZYF1vWUN3ifS/NWYXPOjsBn5BJ2cDWB/9/rCzrcY
VlkHyIWbdBZec9YdCrgwfuIZWD3UhaW8Umg2xqIhHXVXcodwt/UXh8rMIKNnucUI
kWGwpsyuoGXuIm+kvzjSP9ICdnkuKYiWEA/MjFEb1bPTmeDvmKEwyEl30pbjLqO3
gJj12tWhbiIOGbVaugwsvqd84H6GfEOKZTzJEPsEcaK0uYM039Ijk+zg+70/GHIG
ue7Ce7MoacQIQneNnBbdGvE2AfQAZL002592HkBrX/IjUERmembdYioz/ycPDJQe
y+75cwfclzgMfKFerOw9QTtkqCoixP/gq3OA2JZaE8/1VylASn09rA44QhXcrSLf
mHZeYIzq5L/KkyN/JpLAqImjx1dW8bV9/chLnq576pEJw4CJkLejSoAUoKa3K+M5
PrfnVtVuDKxoBiMfofl/gdrHBiURBXlQGHU4dcILMdvuGr8nOydiDdIDr6hU3t+G
KtBMJe0TyCw3thZyYsdykHGrCYn9H7dgFEnE6BCbkqb+CCdH6UbsOSamWWE0rlfA
YIBhCJArmd61oGtH4gONU2PVmpZN5SSuPgD6sCs6s2Ql0vIM4oUT+BYt31CmGp28
6dgVsGYjFbX6H9EMRL952sRJ6sVAim7DWNdb4GKWEe0eEo97UYaFrqmfYwcZZvpu
oePn4cYgGQt3uT8n2T+cpwzP8HYYu4jfZTf1xzI9uZNp5ZkbvBIi+1H3EBXlk2Ij
`protect END_PROTECTED
