`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ob1a3M9gR828y0ZijxtGoEUiQ48JtfOOBkvFcGSqMP7PTH8nrxthdeOqe1oMVujl
lSaHhlyqX62EUSRwNXc366M7a7Tbp+bj231IndUj/8/ttyreBc/oEsIaOqcyqg4D
0J1u3z2Di0dIVPMJxxXXPyL+xga/4yAvpKJzERxCFNK4H804h5KcwzySPe8OA/TH
ziyoswTng48T+ssffswP6LN28PfmxFJfPpgZhuZ9lnff+PxDioztV3CvdNEvwhc8
5yhNk2GZzX0I6OGx1LjeI1tIXLPNj497wlvnzuo/fpOQ8jIe6n2PzY8mereTK5QZ
APf4/j4LPLLsj4vKc0HTgxBQdqFgL27DnwdrX+LyqYHNUrVkt/EILKXl+bYUjaIC
4EDpeT67nUpEW41QEFSF6YKqlhzMtzmOYsemW46MmCtgYpkUS6HsQvEKF19nYdBa
IgcYTStQLTboulE2uQcUVzbfdoLuSxykTSxG61Yr9Botr6OJXQe1/gS2LodpQ9pW
ZhAlDTATu4T+SwCvGx1W7rbyJFT086W8nqUA33c5aFvjcD9TSZaFI/A6FU3AfArY
FUpNogAvBgknEIMBlUKTKZWBgFRYkwfef4GSMzvlhKaffZadQNrYM9yXJzMG7NHe
fxgiLnOQ/dHRmubCtJ3yQ1Da8H6cZbTHZ2Kxh5arqi1pcMFRHFhGPgOyljG/Cjdm
rmExij564tlozg32amH+EJA42FA9LJiVPBvHqpxxtKH1CZ7mSVCB4yXasxt1b5hE
mzXVzjt5/luz2Q/nsMvYx4oJ5y6j9G4WdbaMJHVOYZ4FqPIn/FLWVSWJAJdcgUHc
2ZcF7UjQR1qlPIfUcdMMMaZyR3uL20hB8eGYHfWlJ39dgsG2BvbXm9/YGswct8oW
TdfKB9iGqxHy+r9x3Oe8weqd8+2D3hwN7vflvJv8YMrHLJx1YsDEpGIdNpmld68h
Vh2AMA1zDoxCTqo9f7s4Em+C61kITgUAosxEc5jkl/HZsVLwokF4GvK6beKBPBkW
sbm2a58wwVlI51LGLo6vgiMuVbVU4uTUOAreuEjSiHNs3tszEMWg2As00hh5fpe5
Cwmi3ZRruZDZJx7/kGdPPJZFvZLaE2K4sFzy+qiuLbrvbGUkRViOcU0slHi5UHip
RCZ539ae5dM1mQXDkN47rE2t61b9GAA5ZpyHNHOwSV9tlEnEqpiC0kpAjsp1gFB9
u+M3YQl95gqwDXvTMNy2jNs62ZNBu5T6dvKTAIFSpv2h8zu4gCQHzQ6RgzekGPM+
`protect END_PROTECTED
