`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2kBAMc3IAO8zVAP41aglGPK23P5ljJf8SvNdraCImqNl+meIVw2lTfelgGSs3f4t
8x1PtdyzBy+rfFfhzsczn5n2st7aqO/uZ3NiFVU9I90kAavJ4MyFD1bDEKvgmkYQ
FRQYmmUL4AxFqhI5iCfGQXIcFX7yqg7YCSk6ckE2f76vk7UXBo1jnhfM/kQhgOsH
EY5tj4CFccD+8ixK5Lnjc8eXd+5FAavx+Iu8eyQ+SQDHQZAFfab11IjaGOvGbwwP
x8MyutEqG6X49P6Unjc0sZrP3JB1vUlv87pwCaoddP09bl+Yrezb0IpZ36bqdzHi
U9zP1OQZG20O9HVf1ZTkRVOVwVCCMiEb+HB59QHXlBydqXGGjDXqXxbSuFVPuMed
6l4U5czV0dynIxPBuZu/EvMQI/BWYjGA6z4+QD1nJ9onAtYv45N7diihy2r7gz1z
XTOx0mCDEpDpU3T+c2QePquJk7LOktyZN2VOr4VfAyXo1JMpF7g6tFw+UKzngUX/
Y+PsUtj9WDuYQGxqQuLVfiJb3QE8FDTvwV9dSjwlaZqmlxsZ7FNySb1qEjM68Ukg
Fbh3G4iUctMmKJza6/zrvl4csZTnnhiYv3AE7WhRumSjElVHPzLLBa6I2Ec6OYal
sVEREGPwslAMy08q4UQIG1Y8EGmwsIIwr5Xs/jiiuoYIMz4dUmNXUIY5s1+JyrCU
PTR6yuukVZDfTsJFeB22hRgnoJN7956WiWUtLesbTrl0fICr53CoSvxq6uWqt9zO
FlPwj0OvWggtDprriWBxQrHC0aON4rcdnkkoH6gGdkuuun1XFFLOW3TitSg5Vb8f
LIn5B7CicAZZdE2q+zls0Q==
`protect END_PROTECTED
