`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+uKlc51xkEstflfrl2N13uJDyNb9JhXMJLix/pgUrMAERCinWaNsYQ7oz2Dd8kuI
srK/V3NHxUE0oAS4atqBaWhEw2NM9Qj7kkflnVVxzCImbQ5KVkBe6UMyfkJ5o7Mf
zZ9AIdTGXNHfoegJ195aH4q3cUbWTHj7KnRjGeSI4kOMXLUYyiaLZv+ZiPAjh0Qz
aCMcZrz1ltiXxgpgq6uiqoEki75azAFnBInPPRUaLSdCXwOfnHcGQzMjPCFMVSNa
OxiIaUN4HyEMj+0VsHfMvrqAW4XOzQiKc7cOxD3J67JesBcuAfuO93fTMDb2t6eO
wAfuSffzDYJwEk0hnn+XAZfcLJ+Vswe/GG5FfEG3V1n4GEvLkP52x1pObHZ90+jw
xuwH72lXBY2diLChmYv1u4Mr6zoNYlAeAa6gzYsd1B1SVKd90hwZVCPGKsbJI8SH
V5J3x1AIBcJbMHa/8SD247Q7OweAzKJpHjDOVF/k/Sv8uUcg7dn1HIizvDAHjczH
kxorRgYZJRhFgObVEzT0UrSBMezfPuQ1mpp9uBMjnWM=
`protect END_PROTECTED
