`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dUnvm6Qm+7vtszzbH4UtTs3nblDeECfQPPbsZcK2lAN0JJzd7lRDmdUXBk3GsU3q
p11a0PJ1xyNkGxDWLAdDQ03Bg7IhiFD2WPX7mfRxZl9SkeVuMKp++0p7WCAtPsTY
4RuaZGQT/NAZ0+1u9YBENL3TZxH8wQ0hYHvkqAwMKewR+2ZQ4fcNXzlbcWdDyGQO
Cf7Aop8x9Fq/VIj4i/Ji1r8Qvh7wTrMrPLDZ8C+QPWlg35tXGuDQhNrel5mM1Z4o
BdAxg1vIhcVNADBwmgMQ8gQEq08wRXzbC4bbnIjiafrQS6YhS3r7eEsVnJvE7lT5
v2jcfboeWNW8ZdmISitbw0FQ5FR+B8oGeSvBAD3f+lofm/PPdbknA9+Az+87zdn3
yyJmKQCre5T0CWQUCCz3o/x/HQRfpQv6jg5zPl224k+Nsyty3FIV7Y9tHttP4AE9
g7tAFcigbUCgqljEw+I1SCjlVz29sZglR64aJovsBf/EJU6vuAAgGAz4VUzqLqs+
5xQJId/WVGzs9CofpU8bcDQZrtvvTPTbpZFz9ghfZzS3EU5P32UmI5G09YSdBAWl
oSzcg4M406a/6HWEp6ggiBUm4A+rNfyOQnDlhgvZEQDbjNxOmleGP4dwzykioaSh
1RW9OtWRedeA+9u4nmwxCwq6VdVn6JdZ8hE2uvr60EeagBnjTWXPGHtr+zENXtyB
G+UqHePQe5DYQOZGE7FsEA==
`protect END_PROTECTED
