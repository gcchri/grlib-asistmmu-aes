`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mkfGgzsZJ4RgQ48yv/T0jwpuMBEdXTQ8Isgq+0UR9/uEGiL9Q+Isdd/rZesuHXMy
P5ZXa2OUXDjBHSoYYEiuWM43wursgGtx189fOtcNDrRNXmvz/O8hriRTFA5y/oix
xhcc1bQvTWbxIE0Q7fCbUWWnK08OV3NxMYJMTUHDtNpea7C8RsQUlRtA76QF4vEi
ArStbtPZnEHwMkbh7EsgFE2GXyvQbXS/f8+z1ouvgG1OWvALkV4BPzCXR0YvF1Ox
qePw6d06YvBnx/DF89n6HL136LswSewI0mRCmT17l5Oga/BJG//bV+0c/n7tXM5q
zKq2506UelcIGg7Fyt20YOyvTIxs7etnlaNjVZF8AHr2ucBGzAhaClI+SlwVpHgm
OJDzwYQMoZ33I8uBTkjJD/qQWD8HfEWxYrlx6uql9PVHajEsAvg1pS/OO3xFHccg
Ck+Yq5fWhl6CG1Wgyf/1Eivdz6dOEAA1Xtj+vYQhxf18g1dP7PzWhjdagw2YMKbL
ElKFJwe+ZkAHk6ndO+aR6NmBU8xOUgufZjiD3n5DmC7gJaZD2808+5wQHwCf8Qdk
NgriOkBP1Yal7GQ6wtQOH7J1dH6qVwCk1SjuTChcvgB1eq3CgjwjdrU+LR1vdQdo
JsRImTG3VPY53It/xHMszOO3Ej/qtVmMTKibCNz7CUrjqLtdgdnD1Tx1xRbCh9Jq
TdVApK1Ag96CcQqCOiQrartbWq+hGmHwx7BGkmUsQKxplpNareS+buR96c4cDd2Y
JzRszhdOMO7aMuJut6c2eRA8RhpBSREOv/NiGLEJ+oDBg6gVRnXg5BKJegKxsFYV
DLIjVIo/GqTajsNdlayPIPKQzCQKVxWa5YP2h6wZAY3Q7xvIr8gUmaimYzWzmtUg
Dd0YzSkkkMnZ+wsbI6rLE8d7yPRjKrDdZPByF4BwcURITRMLCpEqjEiFwNL2iPyh
jh6D8V1/O2SQRBbeNm0xXvJRVtnIFsF7whTJ7G0bpHm7GSkITU2GfyH/2j5b8Dqy
1zeaQP/Mf1V8enZsKgnW3akbjFr7vxewX3HZmeV/z+hZfB2hu10mR3JdgewvIpp4
J8IZ6ZcPRH1rtZrj+ko+yoyDnX6izM3+zom+N1PAhAiGm5aqWbibhYfKliMKqeGe
`protect END_PROTECTED
