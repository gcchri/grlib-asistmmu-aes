`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h6Dl5h39HkoFDab8ImU0LCkExXB5Lr3J+lojBBPX797AJD4UKQREHv6cwJaHWp3n
KsENLXZqrgnCVTN7WhHN58YkA+HG4wD4Qjzx5eLYzTbdH/7bDpo03Ils9cupkkgE
wO6MjiNQxiwz1tcIeH4shr6M5chDqGJjWUviGxcXYJPLBcrHDpD26PdWx+zibyEp
LCFetKGn7iGgFcqF0fLw0/ZowPUr8LpVbGut0OwH6jGnDAiEx4sCx03jRbk8HR1U
R6D0lVSQxUm7h55GD/NcYrQpbC6fowtUzmh7HthDDplEIV3eTEmvcwbOQAu0WsX8
a6NA/cUPPHS0ToyV3LSi8aCqKgQkrKAYpCQ5iY+zb72pW8mQXE5mol6qoZdQhJZ3
nfBaXmJSNfPGqLXY/mYeQadpD7aaihHzcTQjAFlErqjk0cZglNdsK/KWfM+xMyHk
X5FIwMuRYg3KIWmhal+hAw==
`protect END_PROTECTED
