`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lGPkcIBWCCajWfwpT3WQ6+8sKHR3Dp4B6/CmfUcYz+tCHrenu+NrsicnCgkSuzja
AYI4EHRwrhjL42QkpPEzDY9yRSo1fcGwnWY3I4jfURM2hlQUcvZ322fUWimexPWD
iwrGA1UyxKQ1Ljx/FvVsg5E56YepH6shWDs+obFG9bfcL7tmsZiBHqDAn5ZasMxu
5CShvHyvvY0ADFaI/TVVvo2ceJmo+lunDJO7I2AZb4m2LV2de+jaZYkAnPjzQ69B
LQMoSRnvL313ID8hnsi5lOdsobkcQu7rybkWZDnQsXzWqWsR666U/Kt4lYptcUIQ
7tEvNMp9foT/gWw/GiJxhWLbpYemS3bXkVd+BAl6Ch/8zVcIhj9cAskHrwCWys6u
j1END2kMGTalODh7eb4UD7Bcn0F/TFTcscXuhN6dwCuhpBEoLJAcyGSfXrSEN+/r
dbVMRYzFPGOlDEjWq3Nv8lmoI21kMwT6K6nks86TmyRD2AWo94wjW7cxTgK/IqRO
OM8wCgwtURNcAQa+ZdFfrvke13oH0D+eLYwDd+a16is/cB2E4HTWK1s7Jk560Q4E
fgbZ3/j2jFDkFx3aG1IUzt7FqABn6gCMpngNWFo2YOldkix03jhQjDKrw36RX7aw
CwPP0b7pc9xqtTSURn0cy53x7zmWVClzqNhxgTPSi33iMJile6chBXg7AtLwQRoV
z8CpwpkHjcey1+/588xGKuTRMxki8X2gofuis6t5XLhAwvBgvpGrP+JAiBvy/vPS
bqHNun8IwJwz+v25JINysAxe68VsDaO6G1tkMVdwWjYko203J/iHQlUsBhKRH2OK
f9AaZLLttHLP5kSlvrqUe6dpYNW5c5hbt2VXyoS9mqtKD1mBFDTHRbBEBvrGAns0
Mx2IoM7Ya632IGRi47/7qDLox7LgAOcC+1xi+XJbI2VWh77jlkB0iyuMlmS6pE+o
3LuUbSx8kz82sKT7W3+QGEd2FE55df59h60JJI/WAghFBWF91Oa01/J04X+MQCHq
MFFYYEKO5jrj1ZkWu1psZM2ij4AO4iglciqHTowk9fcAB+Ky9nDnqjAYHTiZgFzb
r/belJHioL2+GBJ53BY5ZxmpoyveBR5cChAhd+cmkauMGO9PiTXRtOhTTZGSv4Bd
o5+LyeaVGVHf8XDWR7ctYWQz0tM9wn0qIBv9LKCyOL+dMNguLj1x+ja0hzgtqros
L+Owrn+iaRbqNv+Ueo30mio3FTfzZfbK9I/f/rCSEAQUv525rYeLbRpFgjdIuTTS
`protect END_PROTECTED
