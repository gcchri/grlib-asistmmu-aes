`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8rk6dxZ8KVn8HDDwCdw1FzzleqITEGEKegbDTe6EyWdRRbBVx4zR91WG2y2w4Ml0
CWpo13XRzbPS63eByz045CXDabfQ8FQSUBwWtWeSIJSVwm8XfA7KDOg+jX8dqyBQ
UoTV5Z/IWbuW4W3zKL9DSHMAtnQmXCg25V1cvBoFM2NGWLNfhRS9h0wT6RO6QfpO
zv6D+9kLEnZDocM9AF2Mx3iOHWekSmzi69LN6rdCf+4ak8lf/pxqH1s3ZWWZfuY0
X6L2Sww2Hz7dN9/W2WI27g==
`protect END_PROTECTED
