`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qx2RiWxyH0MhoZyTioOMWOjbW9NMYu1ZOVRxMV168vXs8BQ5y5KGMuefgK/3p0rC
1slv+iqxg1z7FL709v1Sn1hqqY9EQqymkNAUQpTu991xuc6DlXLnNIDETnAUweIS
WOFS5etrk97W/5SLqtM07dWoWu2fGuXyirkmZo6IlXhfk8B5nK4TPJ5JgARL8sIq
iSWD+hX7MXd6heiK55gXfdj9PxLJvpCRTSj1N/s/4XqCAHbQ15MeEG96N0ZfdCuL
ENnfoL+Q9SDT9lVNeB2CK/3GNhxLXUicMV6Jwn3kBzLSSXeaAQ++KtQcmybtLN26
PUFeCVY3tX2i10SU9M/NQ2469Je7JtAnCK0pHb2aJw2mEk9TbrMeAksH39KT4CLb
kXyLP7AdYA1ze7o4dTR9r9vcpUTWdEQbS8hNFjC+Z9p2vsqF2IJzUnveUY/mq5ic
7smY30c7rb2/6y3wo3m4nmB390XqNa/JmneRbWVWiigVI3A5iY2b1oFxYuJ3iYz6
yBj0WPIcgtupSR7Oid0UyGMaFTNIEa623bO0sWGrmKq77K0XcVghyhpLl96s/dUq
ljJ6eE88XkeANEPZ02UVIro+uCygpF+nnNkFaPy9V1yqgh+hLGRb9lpa3Kd+i4vL
rH6MwHOapFEJhHP9tKeIeiVkLeHAYucwG9Axt0LoglJ3SfMW26eAihK05ccxpH3a
tiwdgwiPRXny281jz8dcwutb0GlfDu64kbgluUjfvR78cZ34CIBLslc7TUjkJ5OV
ATv2UEsd1RAMqvucpYOD/3j49Q7jgoboDCy6tg6gcqCHzrPG6a59GEQeTfpRPXxC
NfSaoZCos0jM09eJ1EOncmWkw/VP0KSFvA6YNVdmIujIaG83bv1aAZXBSMWdXXa5
5dFzJ5RXFPtuiVkG6aTLvmGl+WF8WiknkpPkEpzlPrGeg/ASkfA3hrQNbdP3CxpA
YDEgIKaQG55gYGCHeaSu2ye+5eLr6siCk1WdOL5XmxibSm4tfYcUoAeyfNYRXNwn
xW5SQOWdCO0swIeJKbuJeOcO1txHA14qblnbDPMLTYhr/8sN4oJRp5/7XlfKfGs6
CspSgZWw9gDfqhFm3tDOjfxrpYG52WVfiQHvEllLKcHcTMPUMtZ7p2qAKN2J+0rt
6qZDRnYkv0RyWki0sJ+THuMM4GL90MarO1b0u1+s0xELlq4TdtlVV+RHYQ8iCF9K
nv7095zMw8ubtHlgtT5iQSck7MJVcmLgT3tYK3SDNzdk/jSybGyCbg0CfcnE9VYx
3fiubpj0UtJeRKO8V5jfkKxMpCgW6ptHcgsPqoMzWEdZuJgF9tu4hewbW3ID7s3W
IPu0CjgE1YMR509/MdEWrf71DI8OwHuY6oKhCWzTFQSWvtEe98lYMb8zEL2HsRQ1
wxNY/fSfAKye9ZW8RwIQQ/+ceEZ19Rxdpj179k+a7EKXepdimwCBRFowjVYxiyu1
dgporJhf5mPclwUDU++wxTKSXcjvsgHM3f4yIgZYNVyQSOHLrVWEGn2oC6wJKMzE
ePl90AkLaAmUFF03HnpEDuLCz5OS8QO3dPg5niy21cmMx83KYMeiI1fswTkkNS5T
QesFhCDcWJ7388JmJejpt1+n3MPb4ebg5GotkLFjV/OHUVsLUdq6dNUbuWhmb8ub
KLG4aMJVdTiZml0ZFtutahFGfQ3xJmKgrEzw+pdvysfoxYI8/tH+UxKoUEGhYOf1
5l61zKYzS9BBY02xBPV6GI1PMFmyZM+cO3dh6whLMDbOg1MtkU/ymFI8cxO/bW6G
3Enljp8Lez/UeyiRUc2OljwSx/ZQQ33QaNGD4MPWdTwG9frziHYZh4LqnskQX0OY
x4GyS/JWr3Alzzfe+JzlApKB1kGM/Suh2EzjBvdt2tYnVmG5s/LnBLmpe/WU7VAY
Ov1/Qo1PYLHZCvw6VaO6RStDRfMePQK2GhTrgoh7hlW2u5FH8CoKFM7LRCwRiVTW
G6iuNcLPf0VjuNc9cEUYp/sZdOsYok3/L9XlMxga/x/d7IvXkX0VmUrocJNdTNi/
kSX+eXjf8892eyNwgVgn8wjkvaqCmYjY+6uiKsVwnbAhzwOf/NqrbT99kQrSiJNK
OEJg7qSby8bYdKVtI85nXiWTi7BG+FYyRtBMd9YSBhFJD0JgpSiY3Xu/sRDJpZ0b
`protect END_PROTECTED
