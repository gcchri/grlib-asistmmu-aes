`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VeIuuhKeol+sk4hQ9/hvI621Q02k7dya5o84QHivh6/23ccutkpekt3b6E32QYxD
fv9RN+V9QXMSwztuhcoQGc3mmPWPl89uaSIXYR3485uRBf4WauamEf3yQc+ADXHH
CV2GCiczRmvbbndiLrwB2G1tr0kXkuAz2pUE3/FxXQgfUEO+41Gh97e5CyT0Sh51
Te9yEpYDm5d4yflm8jsSGkO6t7iYL91j6h1ZxstucBS44taLeDV4RRAe7m1Okbs+
osC6WgdNj3CFHiOVt4oWw8+sc2nDNKfl3SMm4xMxBvx6/89JXQ6h2NzeYC2u1mKv
hrDNywTKyR76qosbq920AL60Yb1Cb68vODE3N9BDWdklSTzKEthIKtPo5pupZ1qx
x1EpPycxFhFUbSjwPyHrw4Ru8DUaLCwSgurOiZ3QaTOATwTKHlaM4MuS0evatrS4
hMCno2Ai0Dz3rgyYC8rN0K9qEWz4d5Jjt7zf0JvRp85OVDFqGj1t5zj8diJ09lC4
yhBRzGNEGzmSkDzN88yLdPyOY2UaWcTraHnNXk4ZyK/r3Zyr4JBN6tF9964OzL6q
fHW23iPD8y2XEiKN9x9xYErvxLJ5ZeBWy4xtDAOPHjuM81CKEWQQ3//mHmGTIeSp
tA+gxrZ4Zvw5q5+qHqUYQqYVpJhr0fYaXokIdRVgmxZIBZKo17CAjJZww+wbw3bv
qaanyIMOYDr8x2phgpkMTKjYu4v8IIgh+MYANlOLivUf1sGtziQcjM44qn9I2q6z
cY0CON+uXR4b09KYkXowI9av/CgYeR145TEF6+AnhtOiuJo/Zc8Rm334htzWZOhZ
D4OYHZAJ9SUjAZktNH/fjA==
`protect END_PROTECTED
