`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aV9Tsyya6fDxhtj8urVcj7TGAhTH+Ni8L0JAY16s4O+g12e0yKDWQDznhapIwbAZ
4+cHghgv0ddyvmOM/GTQpU08G7YZ4AE2GmxwS1WSDlP9jS2SqjrHzzjmg+Zv4WGb
nSNSrvcI+elLczLgAF9EAKRA7gA1LTAUEKQ6Y6jRfobiS5GcLGo+Y2y3YahwagCQ
Zd6mNFD5SE6iUx1k9owJiTwOyorUB2J8xMlN+7uU0FI47jKBq8jJh18F6AQOiad0
4SwNWhyCaFKux4FgHOb05ZsX+cWHViS2b0zH6MEzYZ90LvN4nP/JgdYTtEgg013u
OMxMSSskL2l5T/4Mpzukt0JlmMaPxqGsdBcpa/McNl6FWgPlhwsB1uDfPmXN/WOl
`protect END_PROTECTED
