`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4hoDUFC2yPeAaqVBfjOog9zPWKxSs/NHHcc96aIJbyU4JdBPkOaW3S2M1cPvJhw2
pJB0r3oMtbcH7/8byLohujCutCbkyWCQipfsdwJAmORJTB8B5blcG0/yDwcfKDSy
pXEn32oEl2DXkKOtEYSN2vIRDu4jazh2XsgLAI9Whi3g2O3oIx637XhywUKBYlxN
BKWLSvLbTeO+VGpO095XrnuDgb7DH0jEbw76OcZs+uob28c8KMk7auc8DJNHtABi
wuQqaLD6WPIJvC/ZL1zJnki4HihPSN3TTQM5u1q37ysa/0iikSwQ+K0qvsY/dMNg
zjoC4DiGqiOKVRozJVVQmnh0wKrTC64+M+RWc3QwsXoj0eQ38ADcW4xo4/ApdDZl
gUbOVHdhBGGVdDfttEbJQw==
`protect END_PROTECTED
