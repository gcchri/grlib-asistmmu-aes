`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MsiwXkzYhvUkiReqcqPbyEfuD8EBJo1+SceqW+WwwhXFHU9WUZfNtKncDM8gOlm2
7gMf+N/Yezo8oVc+czLedGH0brSgVKf/je9TY/rOPoOeFFTaLD4MscoSzj8Ql941
kEkaKTUIqx3dJ43FlCT/vmgPdp5f/tNfvkOrp7/fGQ5tbiVf55FjGgSjXXrOOeGf
zirBH8Jzp43yMZ9p8FR8piWB782AhMT23HF25pr8jVteeIK+NV23vl58rS7Uv8G5
8P2I++94Xq/ZwhfSlUxORu3uQPL4rlSJZA8Md1q09g9R0KEv9tGLPl6zpiwKbIp2
khVsR1jLuzqjCqGoLL98c1Gju2rGxIv85L8rdccRKe7Z9Sud1MWgnZsbkgsbJYA9
fMsF4s8eBcqnE2bX23ItwwrTSaHEiPr7Cf+0NnJxhDmIw7ZnkQo8fSpPL/jmQwJM
4nASRLqkKbGOlyVUABdDXbg5W7t633fLMz2Ncxt/oXwIaou6507XrZGEkY08DONA
30CEdow4+NforpxZRD7goMvbszP+hQiVNsckbS0AxDA/XARL4L9b7RZh9rcVJL1z
RogvkSx/WmEMkk8hyy8EGQ==
`protect END_PROTECTED
