`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tcA5iifn8ldu8jkSDCyJ8GF4XyO8BvWTq2XvJIDJIy29WF9fF7AwM0NfkngMpQDV
4pP7SK6fJf8rcqT7LIwPTxCmU3/JL6dePTXiF5D/3NXSpGlshb6BYkzZrDLKsZ8T
nbtWw4GuFoStQq+KGnjgSBr41QUByGTHu3sT1Jqy6YvPyx1Q1DAvHi9LGW/FNllh
fL5v1U0Oszki4wxZ8Dr9EnEC4PARS/6PP/LTbE6e1dhsnwKpVHA7vtobBXyrs4n5
/quo0PpI7FavFq1xE+rqsYBMz0YQxhCV8ghiOsRch/42WMuBlCUS0MY400NQvl+T
EqhYD42BR29u93PXWHt0QMSQ/PhQw19vBzAKsSJbHPOvMGfTpD+dbWBQ6uSeqSUs
`protect END_PROTECTED
