`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pPdqFEyZTdW29tXrhB9WYXxkc/sETAi8sOtRTYRc1Se0CbKivx7GU93slaTioMYN
daR3tiIEqVY/opSbPkaqU5i0hdW/QIS6QHIV1RiMUC1lATpPR/u71K9kG/SrUTRz
OEzHMCAzCOdZAFJh3avszE3GdmSBE4NBKm70MexDKFrr3hNw7/Eia0mrtSuRPbDC
SDrqQHi/7DLHmQvNsySbnSjCToqC4Jv3X/AvEGcYNLATEVniFC1S60SxmVsegqj1
jzgR1edlB49gy70MzRSVA9TyZTNhziiAUaBC9G1jKrd2e0ZTGnEtbHly9x2p6FyH
xREf3EtyVuY/gQSUOPH3tF+tcTB/+WFX6OiP5vKFY48SFajIY/tWWTKZhpVnT/KR
4ajJ/d7xAvlBTIyh5QPUPw==
`protect END_PROTECTED
