`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eUhYjonKedV+0whkE/yEhrQSRxnuyAAfEYQPQ8BdJY6dpTN64EBgtRbGyhnxp2A/
stn8wiIOpK8NNYJeoT3KwFwJ3pFIHtwU+kPR+Unhlk8s/ARqlIKmKDrRU21UAhF/
l5dsCLaxSdb6YzP+9V9my6RXiMkZ3/fMSlVYchSO5gMRzPWlZvcJ3ViRuRPxbM4R
+nD/VeEiqqp7YyDuAmF2Xg+aPsYS33sXD2jaefOv0o2TFE8gmhbQjuk+q2btvbHU
BevRa738pUQygWUSlWCPan99fY1q3G7H8Wz8Lh12vmxASezeRtxa7CsP5k9y82lh
Co/cyvxPe6lknb1CQCNPWO9umbDHKLw89o3+BIxTJmHPwVwioaZ9qUfVJ2G335K1
jemXXjFOmSV+6Evby08lJc4+MHJU0RHJxQjoCNwYuWYxiX94kcDt+tK6eJzbTFg3
jaM9ysWN217DmsiAOij/MWEOkAXysb6sH6BCRAUTbBY=
`protect END_PROTECTED
