`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+dHKuXKnKiiu6MTuld+ky6QXY3Cnb0xUHQCJFvd4YuYAwCJZTVPcLFthAe9XlNyL
5781c0uojit397FGR8O9u33yajPEcx01TLRn/CuFN4NaYE8pNljyHOycZ/6kp3Rd
jnkXoQ/jBF1sPKmf9aMbUKp+Ky5zbLp8skKAg4OH/3ALpjTZBca0bDPDphdxPQ5A
SOYetEcb9GkS+6Febe/S0aUcOtgLByaqcloPGR4bbCuEPGPeGrdTH401ruGBPY1c
KgJaI9vPTHTd+3sAAmFKmKvkgI1/E5VMLLXvEsAA+AE=
`protect END_PROTECTED
