`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ypprctEGYht9Ku0ae2/SslwFZb8bpIhpkMl8igoJADXxzMeSWOkoWo1WCWQ02A1e
+A6kVS7H5sPhDMCYD0x8Q1j7UXvgShQiJhAlO8w96Hda9Ak3UYv/Yu/zOAkzK04R
WcU1rn0Rqkx7zTA8EJNDNqDy1cG6VnDK+Ey2r3pNTbrsCbfg/0CJ8r7rGd5+PyI0
zsORHj6FcxtoYV2bfxaZp3nrY/ZRdqHyLKAZ340zXHg6J6NfcKdIttgrJYCwr2r3
OcoosM+8sO6NzIMblbB4YXIK+SQCeK10tAEvdcHyZhjLuMX63Tr6c7CF9LoMirYa
Tx+697iuCI6WoSIZoV3AXFKuzTePngGzoS4zQGrUeFDXcKgoZeoEIewBAutHJ7tv
Ag9Rr+7Rmnf3EnSxc6DxSk+jmXz0xqavUiW5RoWiG3g=
`protect END_PROTECTED
