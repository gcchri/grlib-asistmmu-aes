`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oqo2LVDoubpFqbk/DeF3QW3QgU6cWijsqGTkNW7tEuyGc/U9F55IQe7omaq/ckbN
TPe3jYdwsxs1XZjOi39/tTSuC0kH3H6l80BaacG4XFETkFCVzzmwYiT9yhGBSk8g
erpFupwl/F99QZVUVYGhYPKJxLcH8K20Dgej6Al7gRM9/n+DnqiKOnmhTOk4pGs/
qM6P4TGMWz6wiR9xMGjm5keyKbcDJVLH03tQGvOZ8+MmTV++ElMIPoSBaAsOzmkq
ykkn2TKBaA8pH9rKU7SR6zfX8sSrFADL532MQ9tVJzyvC2rYCfxPr1eh6sa7xhpl
6YlDoc6S3FKqlNG+x5jwseXEBq0ecZuH3WBdg2mQYXNU69k8bsrOdMfl3G8dMV4b
XW0/SLQjVsTXSHS2jxUGNjJwAkGUyQc8DybdARDsOBIwVbC2mvZTjj/Gk7L4hp6e
PeZb8pOUPnCddZo87ZJDkuAKlQ3lgeaDD5Jf5jjQusJPgb8Mse8fK8QVzvoa/AXc
/jN4/mFKo2XnDl7l7NaFU92mrSqqPX2EcpwXGeiWbIzqbL1nX5Fxh8KkiXca+bGv
uNzOx9EybSnXTK2g8IBh4JKFc9sAhdoV0IR1E5NjsEPvB5ZEV78katmPIKcJwyUo
qvsryglb7+Mg3Ijgne2o6g==
`protect END_PROTECTED
