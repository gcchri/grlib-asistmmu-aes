`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E/d1/vUUnN+MOzzgFWL8hckK60G/8pxncMdXbWAbrouY2TZtxcVKtpuGDuTeqaSz
e2iWeqAWeVkpUEYOe53KveZNIjmvdrOdRX0dMa+K/8Q7EcVfW0huKr1gTA5Whmxl
iQtqfIQN0JNCRLEpkpOPjYdZepLBil/7b911v4X+5gHvXiWvOiH2FscrVDsU6AWR
benoyBuNu3w4WFThE6CrrFm0vSgiAyPNBo9yRlx44bpduhEIJXsNvNIG/d6fSZgZ
HzgOA7HFVfCbJYDd3AQH0oq6+LXfjcvOOqtZeFV3W/rXpk4dk9TOchUGAaXkmY++
25Tgn233K6ALZIDaTcbtmTIg4PaGOjYp0ca3nb91RCuZ3844eoYIeV0aZ7L6iRea
ZaZYXOTCqewBOm2VB5kI39Hk8dPLkZ3aF3lWCuWu93ewyquM06BTvObAFSeBPC6i
qxP1jsd0LpeGtIQjmH4jNHrm6/LhHu+DbwqcsKW9zOs9G6BsOPaj/TQCQFLneueK
4/Blnngxjohu1X0590qXS8YA80IlX0OjKytnOdHqFSG+IleCkotTFd5VGKN++oPo
Bisoe0uQbH1RgKQ6BPZ2sRj59dlYvW0Lfn04HmI/+0MojnnWNPgXgz/PpA7bhBf+
rR9Q49iRO/g0GDvPECINLA==
`protect END_PROTECTED
