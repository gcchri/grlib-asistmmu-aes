`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WbwlJPG55FC/4Jbq1pnlJvQo+MmZtnPKT2o/oZMhKjMrOyYDMvCAbiZUnBPLgcPa
Uqb+dutRHC/RNQaM30cdQnqIrGwMjbK3EzuOYzKHi8+5GDx+TRIMmy+dwWSBDCtT
ELHChUDRXaZu+3KBWzVkKWFod86Bc+HVQfHvgxgKCakVVzflJR8gqmJ/ny836dGk
vZdcE+7i8Z1Qut2M2lnv0+YDMo/f4Gba/UsHHImeel1LKGX/PlGYKJ63upX0qaan
JzOhYhN3gCHSoOsHJaud/AIbL30PDfih5dmIi2/bFUd5D81vdoX7XqaecI76kCPg
ts3ZGnvB5KT1NbzpPuoKOdf/a5oYcdwfzhUYr26W6GdxJ+cVKIur1oViOXyEjtWG
HnynY/uF3dXsdGLq/Hxd4/EsjeUUkiHWVj9jPrpVAdXjHilJSXYV7CtsH6eOOldK
elLBRaDAdLgriErq8yF2FvOpQxw/JzT+ZcnGLeup/TdmFaZQVBjKxBONRJVz4zpe
hSdqmdTmtHKBLdVH7cPQ/RqzPcjF4VIzbJA2IKspu8RUHGFFONDLAXLre1kcvt1+
Qs2w2oeZe7WsY9aoHAcSl+5dcWgh6oNJeoM+RpJz/PD/xPCK/mYW8ryPYC/sK3L9
nzOI2UrsGQfQZPj4xAY4q2mOJHwdbhA4pvMP6s9SvO5xxC3vjZTQ0orHSWwRarxi
9ladv/98tyryUNmjSbi4cJHfyU9fju6Cd8SpAyhEWy4Kdmi9Phg4TURxd1LqPuHx
sg2qq1ywS6WQGk32JXKHjQ8eB3P+Rtk0EDzayyyNZ3vdcgtJoW8QIXzSbpE3+2nj
hQ6v5vYXAKDjdAsfD1bT2l+Kg/dmQkCfeEKXSMxkcB0DgKY9siMo+s4Sm8UoSD/z
Ob9uCv9ZfR+Whq2D6WM4eP7IDUtaAnbLQeJJUBnEVhx5rwF9b2tet6fQMH9sJ9BJ
Wzs33DE8j+LgZClJ3nLhNZM7kWgQrn3Pe1mhnP7xo8MlpFKwqYCVW/DUdNvDIpW8
TJ5QQDLIcnAmmkvZ6niRR9InU11CzOBgmaNWxIIgZW3VRpaHhJ/8ye86+kDtjocM
cLScazpOs514quMyg87xsZxKZRY+iThOXUhXlljz/AQ7h8yG4hkShYeHBhvCNAEq
BDGJE9StmRBQhZ0r2lE2cYGGq1tsEEPXEmZiHoBmAomkf4+OX4d90HW6Tqx4e6sr
JRU7i0mrT9oxyN7mxZcr8BM5sXf0UgpYqYv4EfLjKX3EoFplEnE65OxorLo/ZEoN
Tg8CKNjajA2CjEvK3Bf8VVmGElmFuntEDUWd0NxgFnWK0ss91DHi3DwAvWfnAmm9
zxcvtjVAXiRfhPStOTcfmPznaCWXhvvSnY02Bq/pSBEBQUJ8LlDZwAvXI6qEbMy+
8bCCJWQNaHRCZf+0oc2CCa9kDNHvv9wAViFwjbr7luX7+B2GnD8iSlIem4GBk4cN
o9F6hCwKCvp3RYAtuewX8VnBv4xlvLObbHDKotrmZKrmTu1hYjEG8Yi8e5w/BY3L
iBCAD0xqpqthUTL7/8Yn8CdWKQCZuOz42/BAdY8z609kBQURo/NZBhdSJ1Ovr4fu
`protect END_PROTECTED
