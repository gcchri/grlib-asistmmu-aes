`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DqTfraFyRvwxqISgyoVe0B4bkrk+d4z8eEt9YUUC4vsVDlvGuGe1xcPiNL1UJT2Z
VMy2Hgur7yIauxxURDz9Jb9RMPyas9fZjdDfUCaBZ3YXqxzFMEQ9xqUyoyiV7wnB
3qhsxfJRa5SAbE9dfwEp/qNwpolTglXHcf3xmdnoTfssIVLW5Ro9P9KvdKXyd9DZ
hKecLsPvKAf9RyqXiP+SXPa1YA/WeEb9JZgMIsoPVTQkIapt3VEokKkPMB38SNIN
w2SAXqvwwHSOVQnxDdrGFtPP6AIAThcGhdiqiFYNGpQ9jtJaGMfwGW/Eic3lCQjx
NAJrVfqpRRG98T81fO0cXuuBvK9pAEIrqdzM95qdgxGnIGK8BBgBU9yfGJjyxepK
5QqEXaYe6dTr05SFEU7uXoFExjilRV0HXyQoH0MvtLwmAE0O7Ma3dTGYy5gQeVC8
0qctQQ15GMNg2Z+p3n8wK7n3oKZrgU9JMnTO0Cr2RdrEQFrSsa8qRZ2zNU51r4zW
RkiSOssPz1P5OuxLcJvdZ9q9TihknI4eHqKr7fCCrLnAKmbhKDkAJU6n3xRisfas
`protect END_PROTECTED
