`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ey8zf2H5wyCJ+3E2i3gIBWncJvZblyibWmDiuenrUbmKA0O6sHRIUxYC//9FKikL
8jwngSmBSqEWGKa6yJkkUhAX2r97MAHfXWe7pAgJYJpdXl1X0WqBu/KcX+/YtY6i
v9IqqX6P9A/BeQ/jdtcGv6E0qZq9DByov2GrnXmzbaJy34llq4XxfpuhCRWnnw8G
O7n+xr3NhklPi5C8G5Cn3d20AHWSoZ15AillBa6dH6lHy5bVrw5TjKo+676WleLz
aZ2axbU+J7x3icrp6kpXI4c2TqI5fs9HS8g3EKrlIF4zNisZWda5hJoeBgixm+0u
SzY7ZoTmCiS+l+0ZfJ/35A4xr8HqssWT/gSMGBxJTfW16QixhrN1e3FARbB0F0tb
UxZpeAJWfz+BL8PPUYPa8qw+4hYg+vYzW+PFxoOAIsr86vbEycroN4t4K9jO+7zc
b3ly1xeaPw8HLyyccLZipw2GJqR5D2lbq+Q9NBqVVyw=
`protect END_PROTECTED
