`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KCmTDs53b/qTS7rlYF9b5dkT6WVe1VeblGVxBIFr77JmkEnxTtCYv7OCVGMhlit9
I//FPxiQLiEAGdBw9id9MsLk+g97UeR6dR0IigDW8pkfI+BpZd73zv+MdPrrd4A+
NfQRYBjPEB5giYlpfo4daiZheSgPk11lyNy/PQF/OjEge0x+66idjUMEKeZL/Tpt
rFEmytmR8Vtm3n/7BvmAI903gkVWXxja+CYidOLMTJKF5knkQnu4V2zjiBWc/h7x
FIq4eeFRoQUnhcI8pGyogA==
`protect END_PROTECTED
