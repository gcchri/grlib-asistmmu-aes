`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ty8qmgtDXfDGkqtO7kLSVMJkZo8WKTmKUagnl74YjMe+d3SpiuB3wDaRoAQQpQQ2
WIGClj3iX+RY7fuvk9Xdp+D1Ynds5+iH7ktUvAKLneKfwLyCTAuBj74ln6UlCUEG
Vsx2SXDbzl/j2oLzZrvOSbtMJaoxS1vSFNBOWWCXX4xCfTnGqQM+VXLqQOd4Ur9O
+ehZ9uemCSSXg+v/8Jj51x2nVIfFSMQ9VrsihatOEhnoegz6o7NnaDFVlJtui6ut
HlDiWlIfo04FHoXPLE0yTMMDf34uqtroKs9tkQtAX2QSoAa6s+JjDSYB5C78+yxH
p2oEeGyO9TGQzRSXb0PXdqGO+L8vxc4ZDW85fbRUytk70qRScq/ag0xkM+1bd4tv
v4vkRl+oYs2XcjOOKaGwsWqTVlg/6BNZOHmM48f+ZAY=
`protect END_PROTECTED
