`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+p1t5FBlVwaXPvzrq/RUC79rxXDkV+u0XUW2s1+bkmE2sHLFRuKrRgFz3lig56ZA
6UwSC4KLPMRAL8W9YRwt+ItL8nTD9YrauMgPDP0QDNL8+QeR8BU+OcEfxpLbYWjt
On/hu0MeNsvx6YPyc2FfPTFJXndq4sNSd6iNJMxTIPd4vBrn5UsUnSVGG6HhXPCN
Fc7pGL+fKxGB7nhfSk3Kzygko5A7MZpjlMcD4dIVf664/vp4Mzuf8UrwU0F2f6zw
QNnU/NTr4ndDI2/Qz8B9GOw3gxDqb94SxT2KTbFYBs9JWadLrp6jC0jMhEQm8vzf
92iukCarYkODqOQh7SbVVz0VDUw7Y1LZIYDANzUAj0CLOutyEf1eWrmDk+HiS+WB
RmgfpCDH14uaSBvYMCdJWHPO5mQXEiF33+qvS3viTW/B7wiNzc4SIrhgAEsMfUgh
i5LuppNl0+IGxU4x7VMyU/m0cLlKrdJqbkOb+his/yMHwN+vubgZJ0kpiM/vcCj7
zKCRYMDkEuKT5qJlQzva2GNtf5raC15yTDJKUS6RES7ikvqLpr5MZBuo+NbhEgAV
YM166ASS07ds4lO+BPOECyRJkYnlvbsLyxkeaFmWDtkosQasA5M6nNScy+YBhmSa
1AGjRsjkJA/nO5qNInp+fhxLE5erbo1Nxxz9lYgvf87cHiPWdQJOp826XijSQozV
KEpvd4JlHh4KPkYIQw6zeFKJrDEC1CgJnF4JKc6+VaQI2nm+rHPI1n1NDI7W/crh
`protect END_PROTECTED
