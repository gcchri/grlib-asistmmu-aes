`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NvBnDCh5C53XemSLuCY2Q8+qyXQpxi/+MsRmknjfVMme1P9fCMKMC1VEsx7ITmh8
kR8DTuH8Xn5BRtRalf2sKpzCh4mp6+kLuZ5qZ19DGI+vy8dsZRpOT5NZwBBRn2qK
IIu5Sk9T5B4trfNejF6gkiWIFpOLwdq7vVRdKnVrNFsdnJ42iBRnF9PhHvPnob8B
2x8AgCVtoo9dESVFwzjdlc8q+bvMtyd/uypJ7Dwz8Guv4OMBNGMxNBF45bcQhoCN
mWsnljHB4M6NMBcg/F1nqjeafw0rVyZqpxNiVeUftuNWCFHKkJ9v0QJzB2QumUuf
zj/ohv22AAFUIxPP39TTVjmkD6Lk58sJ5vENYivpsX6NOJp91urW3InfrylLLLdq
77bxv7lMCceAl5jGHKPWHu+oDsDASFNpYeUu0r2MbL7FrdT4F1PfZY3q2yX14vdG
0LyUYW5restpPdYdiRIJONLbY4ReQI3MT7jRcGzNzLsDZD24yJVPfdLxeh/E/37s
n2pRV1KNARlRB9eSvVUhe8F5va+lPiHiJHrRNHu2VjHHmStWkkkaIGLW8iK8zAmR
wMhbHiK+64p9vHQkwjtWpx5UayyTY7tt68+H1X5a51Y=
`protect END_PROTECTED
