`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
menZq+EGN0t7yDzMIWrqp184jbdugJG9Hi/M0LWLo2CJvYcV/tDTNi891zeuX8Lk
I8+Xsx0ChbKd6k6xjr6wdifZopocB7rXMj8SLL56LO39XEnSyZJ7exgQW6ZA7JSU
W/1TCIS2eVgmos2X4tTbWtDCZu6FnDfZIn2CLDodiBooHSVjklpWzw+WYcYT5wqS
kFw2SwIn4TrnjbVU09wGNAuuKgJqNP3V4JOd7aJZD3QogdJYDtdB/k3YZtMxoxbb
g+6Lz8hp6L4hhTv07PNj/6kLbIcE/8d5Vsd7BHzb/3hl6xRr/0mytpN1K81uE3KV
dW+f11ljnviDtAm38WVRKAPuV//MYLAkIB0FaNvRvyL644y9iT0rfLy2um8cSVM/
q30d4ra+fSHB1wlRN0ySlSrGbtcGBcLahxeiDcM1r2bkSv/mXz0QprEHP1pshe8F
u6Gz9pvjjmylxvD3FQIluL9/Y5aXN7hCIXPVp5loM3z9Ji2R5j0ohc7OURbsf3zW
VohgVNFSkVELNvG6LqSdVV3cEXZmd/uCANOBMrF0RkVmnNKfi6oQAVRvrkLb16ay
jaQFq/imhCO/3EljzhM3YVGQdNhveJZZI1vp05lab9WQP6xha1DRiATf1X8fhNT1
62Wcb+7eYXe0rrD8uA+w3HELnnPv6V/8qyZYMKl41dSn7oa+ah9wLr+QFcNKOg1n
J7sjd9h79MbYhd5zaP1WuMYDZZ+u9rnH6JGY5bshgqVSArzyPPBnVgsMdZhOReZp
g9OI54j8ldiVDbQM8hRTebssUawpMuZDAB8Ga4mra4xoTbUHBcWWXnTzdcoUT+uP
vLUNCbLvKfrYTzqz4bCKq6HyCS1V62w1R+owcsMh7hvZA1VZ7j3k0QnQ4W61iaUL
zHg6ANhsa7TwpEz4v7g7fQej5GMpdJ8/EgILrTTpev3/mqkQ/AcxjDOO+jvmIy0n
F/G05koqa4kh6nFuUNA/B2/GiXXJjw36n8g0/wF5YgOZ6twLXV/TjY3iDSqIGQD1
uceXwogpavgIE8B32mHXKf7jno5vKep8wht8XXO5yun+j6ht/Q2baSepYGKdCTY8
PiiKgkfPDmcwlJPvvDZTebewI6A22YLIpOYUePyAESEh/WRLICs8rns4U115utM4
BKSw5JMftczNtB+QRLpoJlo6g1vSRGE4C30Tj4N8o3GwqTMx0KHQUPZJAXhxW88/
L3FNw2cdT1tpv8G1dOSUTvHxPXR6JPv40zi+fru6NariwPEU7+YcvwMXlldGKuBe
CFv/C8GlrMD7FI7GR4leySaiftVsxMbxzlP3moL2kqvxU/YCE1a/iXVbzjcayHy/
32xor1KX5djegkZewH9pDO8TF4LBpK+zmbbhOrHwSdMsyXVtMqZo2ci8TkDxH93B
23tLRhXQ1LL4bFvNTGIjjk3O5RKQ5+gcDXmeIjtOq8WYznu3vYaSPxk1Uy/9fMlH
2ol438FztRLcQbmTAHA0AOogxbgSEwbUEKl5fSyjMt/WC2te7eKNCE1nPLBx/+V8
0dvb0S61VoBN1x5+65ll72bteaxdFd7xUhfcIo/E5XDqTnOe3+lu4RJg6VYB46ME
IFa0VxM5wuDgT2RJ1TzpqCSgrldt6uO0B0AuPl31oRybO9vtRI7zgoi4Xsltut7l
3NFvnVLsHCNvUOFhrk81HlsGVwRWXGKOadSg0clqDrpq3aaYrWe+67EK7yEOO/pF
J3mb/04sq3VjLCtuMN7XxhV5ZI4qzIFcM+k8vhQR3ZJ5b+VmvRHzJ/k8+etk57cn
dZbsfV2+xI2PwXGxAIlPJO90W4i4YffaHNMa96M+Szpmutam5hnDqIJby8MT4WXE
CLjSFmUO/AdxhwLdmUJ/G9TRXtXCWig1oj4lFL9nTW6E/zd+fsKmg4c0kopFR96Z
DAdD4A5GWXvcjDkti9V1+wgnnzqR8/OXxAJsTU82eLJP4Rsf9f3eSTwwOf6PAFnO
lANXuDGad2VwCBAP8mol05bY08lyzb4uV7CwiQOLeLPw3rir9vO45SoJwJoDycaT
XceACiyrCWrj8TBF/8jrQ9QJELLMWnk7KewfLTCmoIwN4GF2PT1qzZMZgucF3GnI
I6cFKnnlO9qCOJ29goQ1rHni3pGSjRqiK6/8p8Veo/iqaydAkOiUXE1SDjzyn1ul
KyjQVVjbl7a5Euou1I1UDP+ZYGs1NN+qGXWrHWLV5/q44Q1IDqKd4WpKD+O4pARI
PYLzSL89tb/f4HG02j0BrIgBVfzVROkWxibO0AcHT5+eK/hb3adUZEovk3xmxw+n
hVJfLqjPow+f2B+NkfIDrcy8oOzMZM1boxMIwHF9V2nu7tvi/YFkf5yAUlH7FvVP
adJpqBVYR+1ua4rI6bk7DS9+ULkXIkH+iTYvKAJcwKbOfBT4yRE+hFMnp3tkvpZR
HAbHQeGujwXMW/2LyfI23S8WqoUdvTkp3ZKArd6QAh9T0/5kl8z5JM5wbel19RSz
Wft1XiUSLJwIgDvxc8lmkocjyV33TsW8EcbQE6oJgZVasOa6oPEtD/0g1Uc2mP8j
2MIQLf4fHdJd2QMkpBeqAnlCtXXfnE37xizVbPx8JW9sJ2p0JjaOlaBiIrHMmjQE
u+KHRlz38T+4gKNi5gT0gPo565mwjnKcua5oPF+WEZyCNwn3CPpkx4NL1r5A9O6F
ffpOgVnjY3rP0qMkdx0p5QTvMrEGfDxHwLxYpUFlPo+dkNEvdgZbvkrUxtIy6knQ
tpLLCAhl1sisQpXMzmNPCnRM7mCoWOWKh4sXTGPxDdBz5OhxnnEUHgbNLXbd2U9L
fEp28sn9D44fvPgng6N1ckK6MOiozldSVhYZMQ7thGu0D6hry/a+lU9tjUjpvvBb
PFepy0H9jMH5lNhrWyPRiglKelrSXwKnfop6dKpmB3IG/7cKlz0Eel1REVD3rtVT
1/OJRhfEQj9akvb3ksN3t+fqFQ8fRWWn6DTEJJq93zRQiiymalRKwbN2du6syGON
Mtme6OTiJYjTOfrcUVcsAnXarp3luyleNMlTqrzR/YJjr7WZHJkVWfRJQy+qfp0h
NqinaUsx8vixkaroX9Fr6pkemiHLjOZovCVHYBpCrQdxfVv1IAezJ99pD4RFaFFQ
6pP1+fTH9Jvk8z4Aj2uQRGOHqIjMYs160sVaZoKFxLy57w0ZoJ9zSER5skZVTryg
sjVMybzBc8OTzLLEyoPcJms1g1ukRoyv8WU5fEeykUgC+HiTOQNyNspJnKCgEdL6
zYvXRiDvk9vVSDBKcJKg/VUG8UGxOmQbDoJqcuIejtwtAcYTU2aWSmh3F/UBP0fA
FZzn+6DEuQarPWlymF+Ljgi57DkjrWbjAYpxyNbj16COPxAwT0rwVsDU3dm2ID1h
FnzoUXVN1mJr6d/mq2Uxh/Z8gcsHhjLnGiuwB02bPsx9ky/PaaKWSL7S2B3AoRH/
sNLUYwB+kwj6mokUIYaEU/QoDjCp8wV7EgkGynT3iW/xijJhbMJKCjupQKgz+cTm
wgN7CYbnHZBFqqxrjNd/rktcC+DXV8gyZKHv/abyeSAUesZYav/HiS0L9cMVtfoH
qa0s04UBPabrzF09ajvzchsjUS8YoowFbLlYcaIZj15jOWkTflj7ZBWwuBNL7Jw8
8cHzbMWPbYT6teM7zsLoKgoKAvIJni2ivn4AuAEFRxVLbXWxNjROyjpj9LPj0ZIk
`protect END_PROTECTED
