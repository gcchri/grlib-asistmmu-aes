`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CUwpN39FxMyP5H8pTFhjlgKkweMlZLUGaPmSBnbeL1zQbYpqL3JaUSmY/EBmfIbf
hjs3sIiw8bWndiYRKFACsmxiBGa0m9imsLrJDWoVKx4ExlmZt0FVJ7JLUMu7o0iu
vRQEdljpBMX17npTvL3B8efs9ZS1rcECgMkQzg2837hITfVoWXnRlyUyIpBygRu/
KpiWPrX6BFt7M7fmg36Kw2/2DPGQ1phcXZsCNL/nPpT84u+HXkcNFVAhMmA57BUG
IKlD8Dik0OMp22Ujd5AGnYs3l6inys7GImDN4kvApl0HOktBSl9zbtWBptZPUcRY
AcBmYM9VSJwj7yaDek0b/MqwwbZr7V13R0wcdYCTRyMRqtDXYQZwEDQ+VCfZpyfw
h4LScmSggQUczcdAgPGPbR7+422LsMRBVKM1eWDKEnquFq6YwxcsR0goKh/l2ufC
abqN8ljT/sN/Wt02E3WvLZoTFoMAepsx1ZtE/CsH9yaNkJtP3p9GkFs+rLDsgANn
Q9+CasjJWaCLhhwGUCBUIS9kmp8WXjsdAc31NOmC1vRPraz/78Jgmq2DsvTchh6T
nPJ+u905W0yqX1B4HPtiW2w07zR8glXNyEeO88GMFBPFKgsqCODbK8TAkktBeg7g
REVafZzU46kYLgAckpWfbtprWFpAX+q8eJyjW3cwz3i2g3acZ3+tG/WV09RViVm6
lPRjx1fHx9ywmUGiweiQ4DGSXAaTlWlk872pyl5LIkhiFzTjFIyfBS/jWBFBZdSi
AvVukbcEM2HrrALD1YTRbHyqFqHxhk6JgjZEpG0zRgWjXNx923IH0A7oU31taqV7
bzAf/z9DEdgT9qBV3Y6VgimL2AWyGhNkBAeoYDiH7sG5/2JgD7dDwwwGjXeHHl/w
B9IGnDnmyIG+V48Y1vIG7LGRp5iV6n4wFrbRguEjYDZdolaPBT7wbrxFGoACbnjN
W0t7vxZfzj5eHxK+z0k7y2YQBbYPXSr5MeGMsswBUyOGvLgThtGRirSyQZSD8gKL
BKdc1VfwyvtlvNuOhfYf9RQVwvrn3+ePnJGn5AwFnnimqOvLvrhPdS4G8E+4qB9k
o2SxhfuSKxPhyxUOguH3KKZ1EJWKz/eAp3xesKdPglnSfsyGJMPhP/vU9/BQKNeM
GFv8FHrWBjpbBHHhOjYVSOvofqoErs6eE7YF2aDd3ArdNooF7VG/XO+sxttSVK9F
hllAvsproQtC0TCdqsKlZp0sJn73o9NWU9wpsPsnE8S8arLM9qn/iMHaoYvQMtTX
fQdlHwb6xx5UOmF14OAXgnFw2j95xSO6srTbUpkIg0eVrwpratECqb0miuVfwJaS
ES8S87MjwDrDhexN0Ix8pg8N+O2ymG5WqDhCngOroj7wlhOC6oeLZuEfExCzRkKj
1opZ66tWnXVeFC/AJemT52wbkSLd7qQlEgCD5kzjiVeAa6T2grs4l6eZhSxwMwer
IeY+FsSC+YCuA4npSL/bAhEWs1ZKEHGTmwmDoKCq400AIkDWOweHfX7Ho7GtCzsv
BeA5bmZ+j5exJXznhzKdDC76XPQ/vHz/4OeXpXL99GKEdzN9pZzQLljtdnrDJu6+
nHoM5Rdy5eNH6JSAXKWhsirwFFTNkzYaaYoFqnFXyQR5TL8wg/IXih6Sd3lEU0Bc
09QWzF1bRLsw0Dbl58NQCKbUvYsxq1Z23eYEW2etOwLPuNgO+h/HbnU0umVxs6CX
JTDZe/mI1hmBDSculQSKZwslPS4OjS1nA6elG74L8ULdlGneUemZvg6IVMxP7o3G
I2Clx42a1F2oVXKPi2O+eD9tYbSbt2Ctm5rMTp2PkLLxT+kr4TA5uZ0ZWg5j5fcq
aVTGJ5rx74KFv2X1+7UzU1b1HbiUBJ9OqmKinYK/h5oWhTPV4+RXU96K4oJmgBk4
Ie3OzVaF6GTr5f3KYYvykkgV/ZI7OnqK5Teur9vZLI6WC5d6jT7ikpaapAbks3NE
iICUH5bJ4np+LleY49PVecc7faWjCmESvkNpRU2HBTUURVZ3ngDJ0PhfNNj8ufSQ
+V9I1J+Dq5eAMSJw4Jim0Er3oXE/3cZ+meQq5RAkz3ngkcEUjpSJQ5WfFVUaE5ZA
X9zhXEVTajPTukJ4oHFwTzmF5EJ8tBE89Gl9SXBEScHKKQfz2AuVywDedqD3YgSS
kaT3QHuVz7aFy9U+Yf9hUY9Fr5UTNmzB/MGdMKRzMYVfuBzfRJaqZ4pqpZXU06h3
zsG/ymve0C9gH7gIzoXQF6hX7fi8CoeBvRcwOsCW8T8F4OYsnEEbapy2GlBHjj6B
G5lVlbUKKmshhA+V6zCYCaB/KdxjNNmqfOfMDSTOaECVFb0K2voz2k5xynvj2fz/
fs/UORy2CzrHlYKDyM0+r72RngFmbbGpLAEr+cVDbjzHEglnlcBdB/sIyMY6sAUp
IwEiL4wbIpTqQ/uoJAT+n1ysBBpn3/AzNf9tLBvTqmMYU0t0frfDqwEJ1CvxKxZc
8aFCMa4y6MaYq7tsT6gUUVzQMuP9iGPoqrwRTmgPGdzkVgnsq5av9tg5Tm3/uyYu
C/7PTuXjO5tXoQID03RJV6//6eVNYMe4wdgiwHTnfsxnzCaPay2qlaiTNrVMtWHO
6AZBUHzUG3ilx/VM6EwZfe3LMQGTHwa7Es3X4QUXRAOyFrHJxSjGFxn9VfLxqdSr
8qVRq62BAnRSnQFGTWUupf0L9KQpFB0OEYPircxsMI27xbW1D8v45DwxIULkJFwe
5RnVc2ocZQ4VJ5hgCzGU96ucyzhmhoQv1NMAlJ0zZLacZY9YDOYkrI1UgQsrX9Rx
mF++PL9A//uqHm/gW8QxILJ+Hy2rLfT7mWsln3W3MQIIXwPSB9iEQkQdVlfOtX0v
Ei2xpQafWx8n5Q+DwK3hWaZQ4pGgwgIVOMJiogqS6quj2ow/w6pQyuHGBvnpgEnE
K9NKGOIfBiJ1gDgHsBpktaQcjNsvQNaD5EMxsGWtnE73whYObAJ3clmcvYVn/CN5
G/DydQE2V4p9j+CGB89wUzhYg9YIRbRU58UuIBIvU6Kt5J3Q4wW8BVfsDWF/Mfwm
ekaVR5HLEM/XIrhk1C2GuQSO4SzOuNMtdxA/jnLX18Px02JxGC7bCkiOjX1GvVf5
tzg3Vqz1OWiNzE8oatTe34cgkjTOmEJSd1IJ2ayYoiiB2+hGUAsiHRsjAW4tSVQn
4O+y4jdWAxjy67Clu4ZWTTJ4UPPE+DN/Xti6xgHfAbNr12W5QuhrbMRWHkJiry5l
IEWgpRRwI9i958c5KtKnOW5O/eebMCRO0ZVkxarLoCftgJ3VSMTLqnEMpF9E9nif
2YPN74iKaEJqanH1Ko/SJim6b4dPGT1beE3NzMUMuvCS+6bzuJ8L86oGx5Osj4G9
gayfeE/0DXbTgftCcEUE5nbcU1oQUOxFQvz3EPpWj957DAt8Xhfjcx0zzPpYnFvY
Y2bfiC4d6tCCG3m6quZjFdiA/QiZ+7Q7fPIBDCLK9nIRNeYVewBzsXLDLzgFOk1v
F9syPZ2RPZr+8N4646Tbr7h1zQMjIdIlURJEzzzHxy1oO2n65j0kWu1VkdSw46md
RjKBR1XjD2ZrMAA2E6h/OArPmlVIQDi3UulDsLsr/EVlx4ZAqYFc9aA6qsei9pRf
wclehkVRtZxp7iXxdLrobgzLd8VUZR+3EYEknA26xot5reNfASy8Qg0Em2yftrOb
DIHmNDn2qHKKOtcg7I6c58mUtwNoHvMzrhJ+6ty4+AUAFZbRi+5fuo6n1wr2i3Kt
c3f1Kmg9gRaQoM1+jveJM2QPB+rXnSfIdoIgkg910hVh/1mrpLmTNaks5sv2izBk
xz3lgG3Z3PNc9hpfV3boPDpkGA8BZqvaWFPoCOR0ERcu/U9rWrQw+1zayVUBD/hG
ssyCz/H1jVRh4EcEeXK8ixizdtSxDXmJj5GKqNU/b9v35SXhz9nJxEGJjhQSijMf
6S2MXxko0GNBCwbTs/3AH/6XK+4dIGbY17i3RD8VwZx1iTem97l8u8CUCJ0ND6U6
T9W1mYl/ZB8LYWHXgT8307tbSbyfpV6m0BGiKSMdyw4Tdk4N7jRMKHEQQ589B/Kj
oXXzsvC2PHfEqcWNNFHcprZN7kwd0pnvezDw27zSP0Z4S4csMAF/XiNo2Uj5RGxV
1T7l/UWt3Ne04Eoq4T4FaCEGQghwcTpQ5CBq8Hg1HYZHA26GvpArevBTpZ022TbH
vio5c8kf1M3lRPsW78Fea2zXsaIeEuWmjGt6rBDonDLzFezP+94xnq654XdQmbbD
BN9M0kx6NAXDxOApGm5RQ4/WWF9evOF2Pp7WxBTRrhwuAeBnzOx9D3ovMnCz+F/0
ELpuDmOskl6bopMxOgBXIAnl9wWQN4nmviwmMmfABmbzRRhapCy+kkK5StZ1CBw4
jD5TsSbdhYaJgGy+Ti59mhK8JgWy7ZdCPgtqwUlGnEf0K0+q0oJXPYXrVVDsJ0TB
tlv2jMCZa4CmLIWmdBBEiWD9Lx5d8eI8y4k+Bbyx3Mj/ryN9ixZ5jiWnWNSaIePN
QIEeCM+F3gOMeKrWQKaeqoojXuRXRXbud98Zk197Th+6lMXIZa9uLZWl4RBVo0RC
/YGgMARyHu6K2DgOFtkEjlWv9+8N/QNqTAtC1Wi5HBcFxJpaMVzskJq9iucnyXUy
qQDR+QoVMWn0uKX+KsQF+tJaZidtyu8HxN5ipAzxq8BlY1Gv2Mdni/y+bkdujQbj
AvNVqfF4ltepEuJbyhUzjdmRV4/r+xpk/aZRHwqP2XG0QFoZGBYVWBb/czDeZOsa
mIJmnpRunpswIlEVj1BLewYgey59m6+2RAa/sTeujwrRgpjupn2y4OS23v56utsw
gFzLLHTjiApLMGqlGoK19ZHisB/dmBMI0iilbTLygRFiXJbBeBSsnw2+raTG5VxJ
mvWcKgPs7iZ10lzL9lDh9Pallz22+D8szyB3t56lDXPmkN4T/Kzwlqq5MPGToI4R
ZpfhtxgpzTBO2Epa4BGcpp2EFiglbRgIqVd7gB2aQRX5o/z+Ohs7loX7/7Doo+0t
iSO0GaMPY0THl5qirJsMepAGKonh3bguNMZM6EvPr7N86j2zT02fHi8HnxSrPJ0F
5lHzvPpcTvNmvmaUKSjNodUlgJ9tz6saO2kZa8QD5ImR7u5WD6Oa7mmu18Xf1rWm
jRjadJTxfPel+G658GmxiHh9uJkw7bWUD6SFE1rUR0V5GFfT+/72S8jIKE/egApZ
nd6pEwJBFjDStRZ9qxQcxowlA/ppReK9ZoWhI3f0sRbWpsfXdO430eVt/Ykdqxww
TiajgPrdLHWPOYM/JaFr/9g/DYOpCL/qHGW+UhD0nZQ4lzAK3JDpkvNpi6bArfxk
zn0+fFLwKyHr2kcJRYIoTlCPplQfibDpXR4f8aPtTKelzVp1MpsSJsoWmaWiLB1S
FWWk2Jba5SsLoiDyx9VE2gck04/aLRm2sVFuukC0qpR/BCwG/kus7uiKPP1gg9Tw
S6nrx6vtujeUqHyRkgQn2kyqyHgI29bzgy4hu43U/WpdtC8ybQFxU/4djO1XWzw3
0xCfTDNePUw29R5C913g5SNdKy90eqWKZnDgG2RbJ1vu48zXe8tGEcxSqiIzFCeZ
neb916cw5dv2cNNa3cr/+MmLXchfefQZ5c4I629cOBiH+QqR+1DEDUNoRYimNTHs
ZFTy8QvUbNiYobImift2D1rEGW4FDTVssHJ2qqrVTBWRXxOETjb/9Z0b4MLMJJO2
sUlmfE8Wrg/xghyvwUHx5ViXvjD3Y1tFgWcbZ8FfgftNORMYuZa1JXrRpYIzYGhM
5hCFzvEAE4mSfm0/Dd5zBJgjg1LRgu3Lihj5S22lsgOLWqaBCsGOIdSmR6/+K7Dw
KyvLLdVLwB3Uvyo6n8NKMZMVrFFPGTO/inr/z+ZCFX58DlNOFtIqhZBZhYzUkV2j
Qg+xwkU/ppseaxmNNERB2wf2vzzGmTRErpt6SkQKZlE3d+xoaUrGljHnZR/GhiXG
XqANSkgsC6U7pSGm3PVZ4Pba+nYPF+b4WUI7cy+aEhZ5n/7jXe5O5dSFBrSWHvcW
xcwloX8JhJKYKbvgbQN8tcg6ZS8YOJWgrNgumZCQQtekBiUZ0qMcAACZcdkYdTl3
97NONL+d+PJJhWUyq8fbJ1iMuRwmw8EnTOUTo4nrxTUlkLjqi4GE+9a5BJXcIrfr
xRCqgA9S7XSfq+YQ40D1QPZh4180h2KLm0hiknQhSyjanXTk9mdT7Vp5W+tb2aFC
9XIEwN8Riql9rvW852t+Z9h7UQYrbVLdzNOG1eRNGl0cpeIzkR+P+IZzCe+bPxqA
8vCfGmbaNGPhXNfL2gAkym5wRyAFUZI/RNyRR4qrErN61nPiQazABBcGlbfsexLs
rZovDaz4Cvjhsz/b2sJxDP72y1nRUXoyc+pZqouJ8QiZnTyMG41LHCAFcA18kXYC
eAA0X/VL1rpaGiEAGRFGU452cm3momLX7oJioqNj1Hln5TU8Db1vvtsrK0xjVq01
sK8bGIOzvI3OnBm1/tBJPjJ0pHvqfDdqSEJ8VoPxR3p4/TiqOp9umAzSt8tl07L/
wvpfKeex7irA17xaIm2WH2q47iw6/8tBdgElqD9gKJ6JZuu07Kx79qe97vSIcH8/
ITB8j8fUV/JaqFEtvrp5Sy3qTCXNLOv84K1vH0PgyN2RwZSk2/o4OSW8RfILRWug
N9SenRN6HkqNT1BatD1tGrX0EdRgV/1ieBspEExEZO5Oqio7GHxZ5nVP4mg5pz8v
MEzvfNWCFyvu/88S7BfpgneeG1gbKBqv0FZKLhS+8Vlk34aupBSRe6SqSnbWVfzu
c9JODQ/2Tx5E0JFeDc5H2CD71V5u3uL8heGdnpUQzjVUWQmx2UxggGInmVgIhY3/
W4EoKjeTSYs/gsjzMfvKCAvUqezidVNBinAzJs/m399OPkaVgFpjHTk+0xXBkelZ
6C6mi3JUqkgmA9+AhFShjfnpO9BnvNZWmp+G3lkDAzNfQ9GeqgJv8ZVqCUy2+RtG
hQ2umJOjbq/4hSyH3QVm/gNjj2KuH9eU8upKX55++r9XB/O5sqhhM0rRFM62j55j
QHrZcKkuYXt3ppGLzU7tCfSELlPruO2oaZ43S0pFTdsLycVGmRSudZXbRBd5NXYG
BBh33KgwR4bXHStx2VOex4WOJ845SsPSTg+rIta3umPJFwtz3YYkYPXU/pR2Qh3y
aXg01o1K5jivhCKsBIvDquqB3mLBcFQ74KkMmk6IKoKJYQwGHhCZPGFHZGNUU+RY
ZUZDv1BGoJv/Rh+v8zrK2OYPbG18DWeF20YprvsvZ/g=
`protect END_PROTECTED
