`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sGphcPsgYKNTbsPC6EK0d0J6+SAyTqH4HthtYNa/4mcdz2Ea7ew8F4DmMc1ZP9fM
d1xfCGbxO5FE5E4+PTPi5f2AyScFwQbylNJ0y+d6o94+v2YS1PbxCVRYE7S6bjVF
kaIa3H9PrKwxhlsxxQLoJUCiatetMFl1ixSQlD1Cq4MqVrUMkbLMJ4kY1tzJqUkG
L6X9tVkT6JCOlU9h0LejmNtMyDAyT6WHHkw4HVTngxXTJRDQXnk+zIYwfvPNqMX7
y6ijR8MUI/k6JuVayvK0sGb/mTEzmljuAZ3dhQQMDfcKJSAltisEhG47a+TbCOBx
lGSPFGFN8bGiQZpeXdC8YkpbD4gtaTaSrqMJbXUVZnBHFusR7e6OBm60W3S4Ps2y
VQ5pWvA4DyMQde6HC+zWsFTl5PFy9x8+MzcL6Zr5KQa9OJO2mBKB0vFY0Pj84pS5
TXwc3VOCx6Odl9Pc5fiRVGdpwjI33iBYgnLoO9YSoc/CyHKlop4WWMojLrLWSx4l
EsWZWjGk7eFp1MBndzwcXD/I4Q63/dNhG3/Nt57bwFJXXxGnClEue9ve8QglLDmK
KqlmcOpZ7udRTE2bzpMMCQ==
`protect END_PROTECTED
