set vhdlList {
