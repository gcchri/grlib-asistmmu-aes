`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QEKtLWswXaiP66lVPJdKVDXUgk19P1JuWNwUqw04jesTId3U1+I+ZjxODJEXurcI
PjVl/XWv7Cjsjkce2S/qtu9RgExHcKuFWEP6qI5nXNoQVflbp0+ZG8UvQ8hNFRjr
+y8ry+/WGdZ0u6VuG7AX9eTKY61L1q7LeJUUrE6+IFbqe/k/EJo1CF5Er+onfvag
xAlaYbyfJRtgKaOhcBJQy3jINJnI4my2edJTRTI1QuxGxwHcvtotpvrp5GW6RfhK
hEflFZnvBLp+HX9LFIVV++NbRUjv5sBE9A8G/u7vC79rT7u5Xn9OU39ecBzCvPa3
BgVa2vUhbP+H4xWmb4htArDViOkhJCoI0N5eCP4Q6RZ4zrQISkhqWTAVPWT/WqEC
GoJgGcy452QcX1OvrtQClCNYpK9g1pVG764P3ILstfUJ0baDgnZ/vK2jp9KfM5T/
ewGG8YWQkhBG5vg1LGIzTruhXlxQEHMhiFVWK56qEwo=
`protect END_PROTECTED
