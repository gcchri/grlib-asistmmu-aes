`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XB9ZayWRYq+KZjPKbIE/QIGvMi4saJYjPGkCKUpcE8T2ieLEUZt3c4T0iq0W/dfo
ViRmhgIpSjk7R0lM0Syi2Lq6BRJpEfKZi7XgPy3X1REFbsKTnWmG2SylfXnq4JdF
jB4oc0tdiTJaQDykkj6VpdAlyU6YqFMV+UlEN4/zCup6XJLvSYXFMlVq1JVQUlbx
yEpkICNFdJIIseQmnh8AonFkiv0VDGiKionSnoG9+vMGvIX9Z/c3jMHQsYA3h0A5
JCRNC2wXWCoTv3yB7auvXci04pja6Aa7pdmZT8u9U+68n7IHQpeHVeFqJhFVL4XX
2NhmbQYfmIHeQAq+w6nMJHJebmc4Mg4qrKYGRp9lzl1DkVUZk7ld1hJvEk0TgGKh
YYjc9Zy6tctrU218qAarZxcbz/1t53uw7jty72wAyeI0lZotBTz9AEuKSVMs7CVy
ZfhWNhNGE8siuLNINOkjADXkWuXqEnA15eGzCJZ8vG9RhzoFTWQ7spMENsJvKu3j
4iZCUY8/jKB2IMshkC2xswM+fD9Ktr04yw7fa1pqk0axV0NILnvOg8OcMsqJizAk
rc7SOjd33YQiM3FMT/L8n74NNZwA/ZtxtGgja5vyGO3u6he7xAETqq0JbpWYftjh
1SLXx/4M7xalZYQjQ84PP6ScNoFqQTe+/ykx2ZdCxE2DCgS030Ngg8Bzlo77WvWx
rwglISGQGEA/hwbq1edV/OEL2bCefNpyabp0UOLi2WV4wbmjOBAAu+ihLnHREvVl
49btasp6PF1+/bOLBQiTmMXNhOfXtgyPb/OtKCLQmU7LFRP2zMICwwCwv0cImTri
7E+edfDExhbCV5swJp+db2fT0u3KqXyMAkfEAPwWqfFfCcl7FWeOxup/bNlOIOqI
VlWb9aIHa05Az4/KP7LHgV8gDpYM87b5p2zqGWOTSk8WFeMqX2RktY9uPZv1/XL9
4ylwkq0oozQq5qqB9OfuIpE4Gi9ECztABsGvRcBpNyCtJwC+V06rxQ5sGU1yRd8K
Smorz+NhOqHKNvooJm0eb+GHzAt9gYYBlgvnykTGXLwbkat1k4i1TBgUQJ+BkkVj
486zNCye75OF1BYLJxtZBuElHqmUw6BLlVMUkl1JZcr6ZTrZBUDvKU9EzJoxxTYA
kMY1ejWURTt+mYhxbDpsPVIAh5J7lbyGMnXQrZXma2wjeVuvurSvG+aLfWxln2ZS
bEzzZpoqhdB0fYL071LDL2XZXvyflLjGuYEuxke8//8CR4KuFn6SHuQ7pOitIM6J
oYgLC1Jx11mwIUOCaTy3q/kGmC9iNxe/A7/SdneQbVz4Pn9A6nA2QBba57cWX9X5
EMA30UN6YBJzzCMILxJ20Q5TkvhmF6Nb1CwFint4qzdbxyRrcepnVi3ksNK/POC6
8d09f1kjzmcBlGJJ6PETvoTFXn/ewGcfZpNlFydJJ73xY/WYEL/+MutFDMIAgncv
HQFE+3UV0GpsunrVAi/JaiZuZOCNhTs+ccy2OMoxsZooTSax2hd2QrQj/OVTNG+N
e1oL9ey1UnonAUV2pMP1PUZsW0Uhoey/JG9y8ahOSO5rznGviVwgek50G8Zt1Uqy
nGeaCxtHmAjNYw0r6LXwDN0a4Pjcrx8ojYjRszAHMhP2GltKfhB1T7tMdYl/L1Xz
b/dLUClMrJZ+9zOMLa1GHpb8SDh4KtFGlKXW3TMkGvfyEpfeN2YuYLVZR6nQd6nu
yzvCiTX1aY+MkJenPiY2SPrcyt+8Fy9CdwA77KNw1jorGJKgiKrw7f+9p+wvWVjK
wgAdU1AO8FDHEb6iDnhqs2Gxo5XIfGnwj2V4QywQHKHtu61amWvVfSM6aKMbO/8z
10UTOgZThepTLZ9x1r3UVlHKjR4S9RpovhjA7/ykaI8cB4/+jc/dgGEJ3TYtA26f
R0H7e4PqFVsyZQi2YKLPUT8bOJAAKWYaWrZFLMML8kt8giY+ZlE6lYo3WzhsiNG7
2ja0ve4PlAy6RtYZs3KNl3ZHbv4I3Kp9annAAehmD/8qppe65SKvqv6GP+FKYwsm
LjPk6b3GqooXRrfPwGDfQWvGX0mEpzqNd8vAidQ/1gJsMyZ5izrkNgdV6VtLecE+
6iUA6SB+6zLJO15HrpOILo4zyI6Uk1Ps1nMqjE0LEFq2OPuoKWAdETyEtASq4SaR
Ajb7DYzXGelDKolZgxXcq3LJCSJtXiM+UypbN5CqRIg5ywDrWMZ/VUkJ+T+W/7PH
RSCXef6bwY01n9YfA9D2YUfb2DR6MJeImlnz7vnU7djuU0u+bK0sx4i2FYpnteWO
5YZraVY7cgZSZ9zZmh3cN5YRnWjNo5iicRw7U2d+NUHsuh48vfoGF3fSS6wGLKam
2YEWdHcqxcaepvr3lHQpXL98ZXjJL9x06v8OLBXKp2qty+G3dn/ZYTgI1pciXVYp
UcoPugmuHwGE+vRHKsf6XTlNvG7ndDO768cOPrDjWf5qBcgDG0Vd9VC+f/JsBc6y
zXDpXoMzRuvxLYaWyRVCVcQ0wcF9KWVWoamFgKFj6ce+neJUCU1D5NhFqMjl9EKe
JGLoxvDziwIuCH7vMVaRVNSXiSqDBiK9rx5HWBhD8iIID9zH2im34UmGMVk470xe
t6xOYKkoN214iEGqo1m/TxZd8zzABmAroIZgi5ErUR7R90F+Dhwx2YGIb76ytBLT
khsvYLDCRNi6q4Sy5KP9MJRwUzBUVhPTWcQ7501eQ91Cv44+pW5s2PDeQHd0D6r2
6pMpaGnpBz1LHv1pHnZuvQTGXzURBu2ekrFo33Pw1JLyFB2MIhMYrRmcSmJTsNNI
8Iv9al94RPPYsMEydzNRBFGMchkINX8N3cwPRmsa9pucn355FUEG6Q42bJ1jSVgz
ZOLHzq+C5p9ysb6qoyLv1ULDPQgYo/8rhvX2FElu8mjExDVR4zChBPQv4bAfiMGf
uGwYg1KPqix9HlYN2Df8k1Wt9Z7oNMWFzdOCove0LJk8Xsd0f+EJ5I83LItWk6Gu
LOxIsjgjvgLwNTc/rS/qw/WHPJgzMNB1fm6V+rt4ByDSjjALQoet0APA89KSNz3/
tMNnYt42lVjDq0yHVnwoxGVvecetEWGj4/t0QT2UTywGz0D6agWllYjDFIUWaQId
gtRQa6HP3a6h2dTYVUz7C2PfzSXBNQbhhRBzqF21DG+yBuAzVNwRwWgsysdF9VS1
1Vbuchrd6lHEs+HeL0s49y5EbANmWjHXQRYJqZbzVAkrAWIO34ovF0QMoeefYowi
CsRoA3oRTga8BrpLKH/b+frU/yKZ0H+Y+EpP+N1tI96HUxofAkRGj5mCeKZzb3PG
Ck+mUP632c830OaGU1ayFo+wjiYFnpjt7tEiKKSWpHgYuU/UdPWvExw3m4GU6hQT
LKDp2K2gigCEzRV4/x8UB2eReeiq1QgxTexl9obYCa46Ku0e+u33ywlnbOy40c/D
NdY2ybN4zYUqzOaVGZdpsqd759oJreR85CqNN0L1twCV3LptFf/7QmntkRoiEHwr
hSxuplqpM9yz6fQwfOu5qHMNzb2eFzEu4i0zxNxo49ee/YWN8vdFW1CAdX+s1FKk
v4LkPEcDqvhT1J3TEqujFOwXx+BLMuGjN3vi4vU3i4pGmZ6qMnd+4QNtZnNZtrgV
5Om33Sdiw/8jXYygttpnODRr38Sr2OjL/VQu2HpJHR77x5jQKqM6zQCZGAoZ2fXT
ge7wD8Cqc4OuIQMhH7XvfH+toDFznF/SYbR9vTIj+nREepdrUf4yPoOG8IpmMHL6
EYegultblYleqhrvi7YZRXg6eu9P0NXQlD/TUU8m0WgYBLPDdc2C5LjzjmhFaLBv
5tp33sj6LeUuqyisvVhO1kf6uhTBWK+xgKt5/xv64LWH0lpm5bSO63rxrusLvyUh
bChPIkioBpKaHpiqeiFBsdI+/XxmAAdyTFNLuWL3hLWb/AuWzUmqnMD+hPXTycao
LyS2CRNF+ZfAc1yXahE50sD4fGTihUSNSXTuYtu4yQxausEcysPUX2IiHeF5N1aA
zqlUko96UoG8k+5f4l3KbL8WB9fchsRIupV4IF8Oe8C/a3nWl+CkVeN4uIhOXRaF
z9wtW1FMWGFYv+E1rqvCSH5u+9V4QibiXa7m4/kObBrR2jcNZW2zhEVtV7bSGlUn
vhwvP5OdPcbXqOiplEJV2D64zoTBzsQ9Q0RLUHaHqvdveu5tBYjE8zMVjNSS57mL
7qH10BvPNmu9K+H6brGUIZ62x7ywRKrP98gDLvgZQCyTpYNSHiMDOy9cHESqRXi2
KmBKc4jim3EjE4TCcIDmTLOHX/KgTtwEwJBUJuOTJ2X17rVTpxXethekP/xx3MPi
v5axfS1X3o86L5hj8E/1cT7S/Z6uD5FRbHkfU9S2yQhkI3f+ogdbTxJK5MLMJXgD
431kr84vNI0WWHBvSFEF5wagThZpzlhuItbiQpE6vPWTKhrvpP2d/2YZjMMer3h5
fpmplCDB4RsHVGfmvrJ+ZWnzg8PKTuAVCIYPTeADKdUjhfC2EEKU39nAvnkN1jn2
n247z9qGmaYeeQhTvEfntpJF2/2EhTw1ZyvUPbFb0+j7ZNfwBU4jxFdPpKibBwUM
X7tUkgMxIrpw+oA+44obBMfAU6GmXsAo4a1EQonyfQHZAOIkQQfw4ftITZNcZy7P
rBnWj8QATJ/7Y37dOrxYQcSwkH1+2pvv1yVssBdvpgsaUJyGEGb6MX4NtPkkM7+n
PP3mZ7QBBp6Tx+IGqZn0bsPgCEsWHapJ0pykD9sqir9ZosG9wx1jILeY8sRwxPoI
S69JVmmhsZx8ICYkC6kyvanOUkolHvGOsYWD5Vtus/day4fV+6rxo8qjLamwZadY
lxUoJjwbRi0eVtZy6D539cR+9z9ouns2Puxg3OeCZGJZyp23Z2ztzuQDJPSJfUJx
6RNm79TdLNS76rGEwKtRZ6Ppos/kQuQokb1PiDQjojruugpLP75t1SNAwtuiOetv
5iDWbbO/qvvsH05L1hFOVHNoTwUgTUIilWHTe0bsLBh9zzHNSRtJwmd0dX+Xqcmq
xChQ911/vnNJWWtZkWnF3qtAIflpn4jKVz0kfmLw6hFu30xE9fUjC50pjhnfhByb
o1yQxrGk947/Zlorhw4JY+LG6kRhMR+FR8AUVEX/pUQPJQkHJJbjaJKhRh24sVB2
WsRgjMZg5RmeSwHUoVgLtKhjBIdP2rdIGqb5WBrJbIG3DLNPDi8ADzSLvo6mQRZB
JLygM4jk0y3/4wwL2s0OTKkdi/iVk4vZWK0n50yuEI4N/jxfnBUFYX2ytj9MEhD9
ZEljZoLeSHzXiFEdIdDU9oOqct+uToWqGkyqYxGRV2kv7KW90d1kjdQ9X4hmoKIk
Q6BdypZLoSDAVQZilRVDF0Sur9oobkCTEd/fS8hHRBXGwbJ4DJn3rljvdAT+6y+6
G1+Wd+hhPWy4W7H5+2E4E+7aBPoRyysipB+Ft7fCCypDzGFyLvT7fIJGWTj7s4qu
zZBSsC72cJf48zCQI48BJtl+UrlcCUqH65XW3iURQ4rPATUPcthu68fbJpvmeEh2
p3NK7eOh+NuXBlqtt1D+7xS9Rj6q8V/5TWnmLsoQue7egAofd2BUk1nXe0ivcoc0
oqyiGXvWrPC2xCIeloWyabiRRuMv7UEcXbrfipG7nWh2WEhCPBFtqFkK/8LHEv4H
HOGpAnIDqiBFOn0WDHWoJX4yNXO153glOAAAl5r1lJt7EHqPXG6Bi/3JTmT1kx/S
61QgoWm40qVVFugta9z7F91qPNRcHLbZtSCTjdJ1phHYy9Hu9/1nn7TCy2AifU/w
T+ysAFnyLdGUJo59oFp6c5JV/jCCmweyr0ypJDASfqlWnvCaR55HjdUKK4PuvcJ/
BKc4o9AmWB5ZYfJR6DogS83hLL8xumpq6K7XgtrcLNBOvE289OBHjlO4KcSpVSs2
y8vBbq5YAFYInWaNmHUCEPW9Pt7Iy05m1YtHvuOW0xcr2OXHWtKSURUXO54Bi56l
pRrmspRdDonYoIDm30QwEQToVSSBveAc4cY5xD3Pc/to3GzJebAet5pLNO5y0HiI
cSWbpTAdti5Snq9KIfCJEP8JU/9sTJQ4iQ37CA//PoovufKX987VrXUYCQPpMwML
ZIa8W+egr0FpNpJCuxXjEoLM5wmN7N1ip15ETvKuUseu1ELB9GR8lQZ43MYwqefW
/6LAZRoV7NlEeNr0qHlckNevoDMLGbTD/Ouk4zuJU4MFanjkg0xGMc/r9iWADxBX
PcYo1G2nLfoI2VlzXaa17qdqUrPI7cKERpH+ixGysoBWKs45Vd5+ck/DHWT0e2Gx
vNGWQL9lqaBmoH4N+vyS9x+4acFAsd/lYYZipoUl6m54yZrzhBqOSiqEla0V4t1f
DJbOrCc/o2RsjmPbVYw8d1+f1H5YUJrK0XbaqBJqCmvHRpwT4QkeWKuTDcH/2M5Y
Dm/4WJtkAaWrKAq5jCHg06VM9/sKtFdbGQIh2sapVvBZhSJGwttqkEiPuVxD0WoH
3bb/B3271jy7JWZsiUvuxfme6HjXRitvoPWB1LwHlCv9ShFWa2dKr6m2fFcTaLx9
IbcLYJ6qBVe93PGBjIRhEWP6px4hW6UQclMWhHzUF7iRt6BbG2wIkM657AoZgAL8
zgmcM51O02fri65x6uobUkB/O5/6hxY/1f90OttU0w0GsGR+dfURrDAHjEESAc6y
ehblIRtHOj48e3rd5N4DdA+M0opQS5iIbMoC66uKKEVAHdv16ja1/M9BTBLS6l1A
EFGIGngklV4B0O7i06s63yb2kUkhUkox33AKJ9m6ECtZ82V8lqOg7SrxVEHmDbQq
xLcg7uw58RZSxo80b8rjtWFYJx9lGchkcvy5Flmfnv4g6Mgr4YmXpJG00BPdbf9Z
ISO6kL2GlAWz4SyEB4koZTDpQ7wkeM9GUEa2IX3yZxkgcrY5/onXiMXvGkIt7dlq
BsRWK256TZCEa28DTuQMTcyPO8psE1ENROr0MxgiNZPnqqsKJs87vaFpuWSLVVJk
eWcAfifapD7zy+yrGWmvN9JB3xx+sPMcTD/p1l0vWASXq+C8Eum5H+NuUQ64TC5z
lQ/V2lTzI22N6JV9RRkqyn2DVJLbDEWINI1gohQa1RnshVmFygdhZrqzkZrpW0jR
8dwNGa6giWfl+LcjYcSPrxtLD+4MWTUBZcA6yrWYJbvrR3PWpmTRG2GEr/ZTj6Ep
P8Yg5M6eQ9UPkU8xIXTp9ffTCLkukaGL4gaV3b4KEosVpLDtgB2Ykdyj8hcBJyrc
Rp/oJoy7XKiCIscnJNr9RUbQvuuZHqjGFyUSAO9BndSHuh7dVHGD+duz8itEkGwh
uKyYD5h8BH4iu14m27Weu7FjHxQdaTpfNJYTGxSTroGxj+YgnWijpFtsOt4Nch7G
YN/irm7TIuJhNV3Cc81BsygpR9mZUi9YK24xYWADfQJOu7XvtvTaxc71vE9VKne+
AZfIxeT2t77aawywoJGPqbq7PKWjC/zlhPunKXlHTbJotr5Sk2ccuMIgI1X3Z14K
jHv2+17SgOj66Gn/bp8jbo+uZQ2EbD53vjvtvHd3RpJzcALpfagSOjOlkm1L2onw
yE/MhwAbUz4SEKiee6lznBXGYJnwf6TiAHjkIPgqnbVFUMEmjmDIn5unDWRel5ct
MoQe8UWsrWmrOFu5Vzs8lC6bRIYfBjieHjGDWcbxrAoVo5URqXlP4jrBPCwotxNu
rs79SpS3zRsGR9zF37/hlBvCv2irIcchqOJiUe09NA//ph5YzWkqJ3viUAM4CtEI
XCcjh8loqVYWk9dZTWFLKGyBb0H713T8knukcb+po4S9HASwNXm48cXyYdsyntq4
Rg3pI3+8qmah6iy52Q7UlfVZdiZVG3Fkk5TeX+L6gvMVDlI3XPNH8PLexon+7XpP
HIFmTk4U8w9vyqXqwG5X93+kdDYQxPK5VHK1Yhf4cFeIXFrqFC0qPKbLqRYhWGaw
Sh0Da83CvbkGb26YDhh747C5GuQvyQK1Mha3rhbDxW5kcdUDS/7d7akYj6yJnGlv
F/dirfo9Ilt9nUerTt0gywhm5WYRG/CD0Vtyos4upqRT0qAMz/i2nibQ0egKS47n
4uKCb7tE9HUM5nQ5LqTbDhiL5N+NQp97Abft1MSqBGkFvy3kU/vnrv0ux2/Xm76J
bhsW1hmibsaKTWBQsQgNDFnmxw5I8ub3aaNatS4+1UBkjWLl6+nIwvOL5ttPuiJt
oPlM8WlYcCw71VO6jugllPAuz0T6NthwTriTt7unWGB+TQP3A9P530vYC/Mv3oyP
Wpc7l7c+SO/9M7harR1IK0Oa6vAdqwkWc71oYu5e32yxEvBgWur86sOV/7HypGBD
aB8Ph8Urm+AVe9mFNm5GZzX11u49n9dib5mtjFH0uhsqwoF35td5YJCDG9Tk8Cdq
jxR+slhQJqBUnaIPsvUfcacRhtJDNyZ/vsZgC7qKaWeOQ38lBhSnwz9Ta/rLlHWt
6RhxZRro9kEDMOBXJx3Bx+wHoWdXgwqJkCUGVktGbBASo0fE/JmOfW0X0VJ/kNBK
vcaF6q1ep/Tq91KAZXEy2LcDv0jNNXsY3r3SsV8jGENSkIumqnNxhr9/GOTJqYm8
HxI7fOX2LncLg+mwBOuyjGz2C8RS4qVv2tspIOdeKVXuNlzI4Evpibi8PpqqVUbz
0Eb7cwLFhGO2SlThgeDmRHhzZMbpbNLL76TwBdCiG7obuhHIOHRg5aM7Kter0kmH
CpSGglbJJ8sefiLl5XN+rtkD3WyU+2F8vHPBqoviL4qXAUMOeiYsevKrkrwDVFfF
SfzERUZLTcv2tqYZS1IUwMsap/cNArNw65lK0bpGDib1QlJBXO0zD7gWeZBPQWCb
6PojfgFql7Lo7VH7Fs+KwtoQ1z3pzE6A+xRcSZOK0iCgwTPlIXUHolv2Ei+DYojE
H0MPRzlPQG2OUefNFi4Zb28m3LqsJkHKW/c330AFZJ7UXpF76iTpzMfWAmWcMZs1
sHi6uX2Pt9iVTpF0ZedpVFoHJt1twumhGxbkjlHu2t/l28AXMRFI5N84yE9OqWVr
b5iKBUL4uJ24UgmFl3ZHNGx5hNZ6Bd/tPhq/SWWhAEBG7hW6OSbhJaD37SX8wE/Y
cg9/7eMjvfms2WJGd6eOIQzSxbo9ygbX2k6kH8eKb3qSugiFrSaLN6JH6VxcHB8C
aclTTAkUTvmorpdCEaEmifX2cjheinN3uqAyDwRhXAusqDKpx3NDBwd0cosjx6em
w08Boxkb0eZpCZiRMBZ4bJD7McmSPLyvYmmECkfhJfPVkpTLOfcNEAcvM5l7rI8i
J/aTMuP1lUSvoAY91YUfQDbA8yfQ+ZjN9ZQbNkWWywDXKL8CFo4SpkW74VBgl6BP
VzvoD0vELUlWku6s5cUsv4AiiV5gH6BvciQbdSs3n7f6q2oihZbWQqq+LWVcalHr
W6D+1x941Vw2y+QZ8SbrUdfoDdYzw4vMOf5o3QHCw9hjfBcyW4kdpHWvnLKkMBIP
0R2XkkBbPJ5YxNyWMC7/F//hQh1n2iGKU9Mvy7AHJyqwNOhPpErObMZOAtLcz2jt
x5CA3so33Hz9BSW+ekHYI2ct/i0q5JQztB7sF/wgz3BHs/aebhFwU84Hl17v+q0m
08ij05vUEu94qz4A1oelFJW6jhWVO0d3HHoqBoqHplga069uTG2Br7MbhFGguaqP
HYlHd8lc+NOfSG/VlVd4EPZ+/WqkbolOcAFJh23VV6YHf80BW/axbo/l00JQCYgQ
ASPNeL9uGw9Hpbqyf5vhc1agYOMkpPM+huLSvGzOAsxhG0UFrIalwfT377Lvpxob
ouiOzBNCcPVNoRvqHGQ9MZSzAsdkdCLbnXj3+uuoDgdhHZ9S6Low5NI/0ARqnAXG
ABJoukvZ9Q5Uu+qXg7p75+sAvPRtotL3IuSNgpKdR4X1auz5YdBAmK0G/qDeOi3r
YtnH5O2PTdg/kQbuQDe5tD+S7pbZY/kR2mdUq/ai9GWgOVs7+3EIznniX02i3Ge8
Xps2BF07MxeVP/pj4sZJOzEbk+4cX0iZ6UaYuVC5axokk8HnOJWrI37BTS9eGREA
7qeH1jplJcvE1ri3lLIey+8+LxdNqBH5p4/q6tc3FMcpL8JHduBwFs0CwtAK0E9l
kGXcdnKjUBY6rlWM8hqRY2kgWAJ74tF7Ihc1c2hFHU9jZPaV8AdZf+DPaoxESXsz
`protect END_PROTECTED
