`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nVzaJb1OK+Wr546zYuIxVq8LqVuNitixNuKhl9w64+q+4ncX9pskQDTyHohnPG6A
sDKWCcmkyJUkFeIM7K1ucxk5eL84+Rdhrun+20zfHprFEt1lJNpRA5iG0ea+7bnH
7jtbLBOaNp7/z6YcQ9QfY7McDdiNs558iX5osvUJjbnqTCQ5gY90MiT2iKyMweqX
oFMSeq38St/kqGPAUz1tkybyHYCdE5T1ZPf4Y3wbhsl9y0FZhqs3ucWJ4eGnH6jL
cNfoK3V2DM6sX8UmV7ZwdK4Dc8JNrEezZWyggao0hz+wvB3KKaq7YaOy3LNsVnr9
ToGXKW1UNmwo6ae13Z6HxRhEbCRDTatYAbLWldGrXHZplCvp9zn5FiueuQzWhed7
zcCxN5/aPtHT+ke7asQIMSLFxh7Er6z75LekgNOIygWRyOba7MwE78gXwGVxAo/r
SKtciJPeWM6C26BV8cBv66jOKxSYI65W+Snbvr8Ev0gDRah9eUSfPzcn6+R6bv5Y
`protect END_PROTECTED
