`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HZr0LNNWgm1sxlxHgmLhYC5A2iq2yqYrGiZeAjru20Ln2Ti73mgcgkce39tgc1Dz
cOhqeXBnAZBaAhsqT5xIU1VrbUoWuvTim84wkg/u46FQJv4qkUgASPeJpeQSflwN
rcWFl4trIqAxqGrX9quxDI0cwVXNifBGmU9ONbRkbzz38KWTjqEaOKsdWVthDBHA
Mwj8jXqmAouEaO8U8gKkdhqi/HZUqWO1SxGK3i31vfYXxq6ZIa858xK+NqzMkCxC
YI39Q7lL7/jjScEV2lzJWm0g4PJYzeVEGXGgXdreF7Ts5xw9bpC835G/tn6KRyPi
BgMuljk86PXbRofA9zPiG7s0PYZEfwF7B0r6GZE7FxfPV0kLu+oF45M9J2k16UDZ
it95Jh47WkHQ82yiCYh1AETT+cXFGjDHCOiB4FucRqU=
`protect END_PROTECTED
