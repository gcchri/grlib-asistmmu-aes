`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v5OS3mynh44MiMKdcD4LPdufKRKh2iF6YA+tGfW44TnJC1UM2dnTCnqXy/VJDMIB
UlMkiwtIKZCBnpEoA+GPSXwTkIy969Gur3oBmouPjy0m7grjmdPJ5IewfEQIPVJr
i7IC/KRTEt/++0KjNZ9NbeCTW4iDdWttr5IePQrkHjD9h2VSivbGZ797MlOLXtp9
SyR6aVArxr2UaNF83Ru3r0x+ZwLIHM+YOIkTWhfKbRtfEIG+K4PTxWenXEauGCVc
DWt8YuipSUFlNpocF+1mhXcXRN6FDeDZwCeX6K3343DLT/Wr2MIcmDRkO4lKFLAg
llh7+75DhuV+1kRUCScnFCIIQwn8NhNptzFWWGiRNcwpSVXYKNVNre8bKOT9gGyZ
gdkdKFGuvrSK8KKgIMRdUu9nyb/b4EIYk1Imz6UoqwrX+ZpTk51GL4Trq6kznDSD
DZcOZIlIvf+Hz8iztx8dnGGabAtDJlZn/vV6LC+pPDJsyFPVhYHPkwmdvb55xoIZ
`protect END_PROTECTED
