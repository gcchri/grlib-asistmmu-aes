`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tQVkfocSLPgc+Q6Dmrdl76HYjLQxOd4+kmw4W7ePVzH8XoE0WpWDyq6fuOfW1Hw5
dOFKEzPe1syh/cpjXaYGF5lifdV8he6wXXugOdJKo+1gN4ha9AkAS63k6cj3BPdb
FBwsmnHjoootMVhRL3ih8Pd8CL34eoua5VTmc3fvgz8FXx/0ZrCh4JUCFEzteKd2
psOVOHAb9GAQvYNlYeZfG60H9aQDqu1yOfZwBqJJdqw8Kis9ZjC7/1mN4K843w2t
jv38akx1/CT+I8WO0gbhwWYoKBRPooTPd4ZougLmsRsirI+ZTmBzwuoHW58trmUL
/h8aTuuQQA23HpYAOMDVif9UJGGl/KETXElFeU6IRaAxMcWQ/BzuBfn8qtTjbgYb
AMtPgLk/1wUW0bCU/K522byiZYpcj/+XqARcxoMBc3xd2tn/QBAsUXBoSh1J90H1
Mjmhq7yWi/AQ6lLZv5l6/BFxG5oO8wXJa9CFLCOhfzYutiMfegK88L1Cw2Fhx9Zj
jH2muTw/Vj2dE6z8K4ef+GUHNUptPvei7Pj2TIwSrhnKgB2T7cVHBbw//e6hz0dQ
rma2urO198CVrZZDeqbR4eDT2+OCj5TYEoTPqw5//U4xKHuBz3QcBqorhrfzeUkW
Ce2RiVXodAH/y53YjhbH/qNSMicH980arBhjQxU/nUAE0LDN+3pmCM8c3ygqb6DD
lKkXKWkYwpW0cklu2VdD485MqRvW7PXfQZ1mE2I+u9B+1Z3c32Gc6l7gF0QEPX0t
YwAQHx3RvzyPISHPi/VB2Vg1HdI83KTaarKE3chfN+iD12u5WMzzKDNcKKMKyhVn
fNPiO7QXQjEjFldBOWpNprc5FNP4HiuYU41EkBPna5plNtFeJq2RAX+ulNrAXuBx
pTDH2yEv9Z4V2LzUlLbPY3IDnMH8ePKKEjtexznW83W1g71TyK8u6VyXqVylYEdx
niDmMqCdW32+gq7AL2D1N4YqdIqnmVpQJ2FN7ruWY8+nI1gmN6xwev2m4n/bo/M5
O/j3BOQeuF8qSHotcnIrzrSXBZ9Vx75PwMyfRiKfBjn5J3Pjde0nv1ljS8aXzuP4
w5nLPWBXZ0GfaeeEs/XDEJm8hvSKflTYmjQiwDSjiFWthB4Bb7HLGAoGKhJ59ePF
g8RT6LPbq6llK6hNZ7Dg+qLGUdYzHiVHDzJX8gBGttVu0RkkeHAaj8HaCORYjxwU
zQl9JTyHPI7WXbAfh42sThz1133ug+V0oFYNUO1Wq4+giwir3srTkL1JcydLRTQy
qxh6znjDqxgBEYUMzzFVEeWM+6jm2sTXoVqCKrWOyXBW2aWrEuyu8R0Wbxu1HsRV
RVIUC5k0fIBKtEGW2zpN7S8Z098HT1Bh4Ftnyf7z5U1ShM6tTmaZ7g8lIAvsnsYP
HcHGUrQ6zn/05PyVYYQv+m1f7w8GmEqFQHsd1o9zJe98QF37elk4KoQtqqtuEg6A
Hmo0qsKeU1yOB4kTDX2IOUM0oKezXTzKoiaWgZPbwmGfyKGbkEVXjpJ7zGQpJqx8
bjvyrg9a0w8lvd1y0sD0CCq5dEzm7blH/6vJrfJ90tdzUBRojjnvKf6ZFDP40LwX
YlABo+cy+p2vVdwiO6aCXET/FBT22KvPxEOb+0i/srZjdMTSdZySar11fdtRc6gZ
/vh+5YJRc2PQ5jWzXwS8qQqAPu1AL16YAxFuYwUpCNkxVjmi2ehRr/qVRQ3DUw0h
nM9NvCA8/MNdOOKn2ax+yy7H4+D7gm78Ej6bDIqNU45g2fwq1vu9IL93w/+jLHT0
QLIynZXhBXuvPNT+eIVUbKEog9NZs1pu2UYuzbTQUvDrGIuPWvUG7n28WB+TLFPh
46JdjemyPAwXlOMSw3IA750MhmR3rJKIrCSZddY42ccv+0qUsXLfW7y5RK18PsJp
xoN+0S9RUo3j+XFoVk+RXiXUEMTH8cEBK0IbZLINWcEmCYVQjHELo4NXHyptL5ov
3wsWOmkIloituGY1faj4V2Xcba5n4KNiXbczwYh0D6wSPpt2qpngZg4xYY4xI/gG
yDxr2PoGd2JqujIIpqX7XQzgPDRU35FVEq3YSgx8Uwbs5Fdxt93hARfbiBy6uEVz
H/z0bKt7L9h9cp7YquzlCZf5YkiegOHJTTjmYuMBRAU5v9k9wLd3SkMtPj52LtUD
G13GqmdF02DBiSijL0ibzgY96aM47s7ZgbdC8+1DVeBHLKHIKSk5/8MfRNNDHJFU
FL64LrYaqMvM6NWNsq9OzLunWoTsYwBHxmzns1O54mEeCT0XZU2XpHI2W9v6uUpV
uDZDnb2ZwbK09Fvetgnr1KA0UthDwZg6XyiWWWMoOzI2TrMwHaK1EGiXO3puX8Mp
R+Iimd/RwrfI+xV2UmtFSCCvn6mFENC5amcLChkTlI27CE1Uvjx+q63bRfOVH8LJ
/NJKmmpq/6bLc/CJEbB263qULHpiYvi7WguTzmlxzphPNAJNhoQ/8h0ml8u5aiwA
U9O/Nq0futl8lAkZyOr0/peJMXy8J7ie0WqafYFE1wPR7QT9fpoXn/9edvYNB7/M
gXcVNvxDhT4eecXZBAvFhx5ZnXPoDEn1r7qAo51EkqqlXM6XCq9qiB+Va5R7YgII
m+pgqWvKJg4Gokfnty5XnaGNyXxf2yDs7XT4Mpq7VHUZTD4ppRxlWLPvv9mYZyAW
PVx2d7JcLyTQ75T9ji4uk1VSvVCrZKJhY/x9Wcb+knqN803qrIyyrBx2pOZaqlg+
O16kfQIw01+Pz/1jhnP5N0mYC6YHdAcdf3/vbZETET0u2BvuXQbaKxkJyOh2TmFs
udWBO7o0T8PTHhSB6J4qeXANw5dL12LZqxiyCc4R9FY=
`protect END_PROTECTED
