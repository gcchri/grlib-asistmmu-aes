`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WwpbfpVZ2R+3n9K+f38BW3YcpfuC+dplnryhbeG79yIU/SBuUDlzUH/3E2yRn8u+
s32u6V5FUixFQHBGuvQ0QgxxLHhW4L4rLpUtIP/c+pbC8jHQb2Rm9ydas3Kv7IKw
14rmJUk3gm8yG2RUD+3z+WQN6ZNmT7Nml+9hnUba07vCCvBauBFebIO77JnbqUnn
MGVWIiJMgQj7uQjqq4FcXTuh0GTz4eNxjKUeu2VwDgwFdPYbVXf9G0nvb8fs8+Rs
/BWYurbUldTc92n3E3Hj6Ziwuuvfv9Q9vLOV296DjDqqXM1QKgW/b2lVWD2t95/9
X30jN2lXSDjbEl0Bl7uzpDgRiZPL7cyLwfF7YxwY18Ndwyxm1eOkxKDJ4OzXdlCu
laXufOBX+Sz/U+VywK5o95O0JEMGtrZddDIxudy2Jc6wDO14RPiEa4UIy8DJen4S
eo0QaZanlKaz7JMXZJxVMBA2a6khEwfCUs/pKlhVoIGzNc//iL+2nbkm+fHvuawG
T+sySreK+jSQrv9WwyVpqKy4dmDJeQ5KVABp1DEKQQNtnOW3ysJHfUbcjK/RZLsA
85sl4+Q1bHyTRR56sFpK4wyIIyLDgskgDR1zwKj8QSVWUVyggOB0yzSl8S8dJ6Ke
0QIzXJer9R3+nijTG55Zs+cPc9xL6SNsEC9RSHpQJvB8vcMtpQaGm7u7raCBCWyT
pLk8l3/JSikJoASC2Nbyemg3sJmIhw14BQ04JaSMGJo=
`protect END_PROTECTED
