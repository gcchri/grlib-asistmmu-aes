`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
19IAlG5J6PGxpvkik1nhR2VQoSeZT+deUGFumjY+Am7ziWOI9zvKkwY8VIgSBybD
Jo7hVw1G39Y+f7UQzHCJpWdc01WcxRDUDznm0mgNHwHHOFxbQFOW/qr0otq5Pb4F
JOBU2WbiGm2uMtFVodq7ESvVh54+rsLdYMP6dPZzjvtuxzic8s2FlmQhCTjR/LgX
Ju1GSeLQu3HsCIy87xKZRoQpnT1A8VZHHz+ZoifK0ljzZ/4PgMDg3p9YTyxC0XGF
jLXN8HyIJlFOHEJaXFoFFpra9aI92f6k3WHec6A+j2Uv3B/n3shMX/ZyjbTithC4
p3woQimXzPrFqKBWvIWI2PIU/7UBmn1/YmdK8U+gazlCQtgD6ij6K/SLKDxC+CnO
wqFhBwuDOR1lLqz+QZCPiPlhM86botwnaGTcc9r8E1gw97zG1IcJc1lyTCyrtq4e
ZbBug6G+OGMFS+o8H9z9W59zeCBznkSzki2f+O7Gon4j4t/PGXkvEVUSllAYp1Bv
xkZanIDjVwoO2ermbPiwCiYPOmnmRQPqS4VhXvpcFowBq5cgzGPKbgIDOB02yXgb
MPk7nreLFNRjExkMBQ2V58JoewlSGUK/6ocPr9ydv5s08X2/9EWqGRXjD9zFlRci
Uwyxal25H1BE4Yo8h7xN4q67xV69ya4tJInuRWlugEbGYuWOJ37dLiPs8IRXLZHs
xZQmM7Bmgosvy/u2Yj5aUFMkdpEtvUMGgKMcoorvXMiZyQkHHvK5/zzJ6K2ALuv+
bk9bWtXunu/9tSIIeQFDy38uHoWGRiglMUlwnszpIMzzvmJiFp9LzRMHV0gveKnU
bre8T9FVPYixx9iez3gpcnIjjLoCmYde73PB/yZ3PgmDjTNU4ukHUhT/Ey0IpsiN
xenzMDKG0OS/YxL49cF/QlXXF5oQk3ss4IKTV/xbaG2oE3x/mRh6fymZVaiWlI1X
p9avTXY57xv1lJpmNdwd0FGGIvojNZGcncIVq0ZsRPQkfJd0529ozFAC1+R9AyH0
YojoBFykNKJOgG1rG1alJQTyPNSnR8JQHQVYpasRoN4PsCh/wzyuVJR12olXKaKT
2afW5asUjL6oyGUmJ9xQToBsM+BMUMYmeYgIhwTBxq6Q2qd1P8D7b/IzK6vNAA1r
rvgAjUihhSxd0IkY8z5Xl4rakjccfBgdMauFhkUzilh1t6I9D/NUA53M7LmpNx2Y
rYjGyfraOIIXKQT+20yps7HMNMIx7ANeX3TETB3tP7zePyUEBe6z8z1ZFFMV4xsQ
+b8DY6WSo07iToNurkVyd6VOEzWeteUFSwaChQkaq5/djxmsgGqTyxgQSW5NF+gq
FryKL/ufhzUD7eCqn1UVp0GF3H5vMpyEQYmxfPCAy46/unzLMVfPvHQ1E8RiBsgD
sLmEg9igRjIGK/wmVnVR/1hsM/gkEI7Wg7WHcmzKVib23TtYh6VnGRO4yj/Bkd9h
IuVlDSQe9QJy/aR3ldfj4AZWEBqeMcq2TUfVGi1Bmjux05NSH8xQxbYzdEDpTJ2z
sDOPnYTNYMGQzJ/IT3lA6n7XCJHHIeDQI9VeVGBo2aEXNk57wf+yAW6WvRjUgItG
OH87B6NfF07ycgKrvkwisntEh4BPCz17cRD57oB3iM3pdRLrd6LUAc5EpyGfv2de
egTlp6ORYQ6WAwWNmH4l92xrKiEl9gmsg0YOjleOcL0fMxddsHng2nhkegno0YgY
FpZ1wI+M1zAA1PDzrMh3zSh8vGJWF5pDkaEM5PSxbQGLf7OxdN4c5f+QdxK//+GQ
hfezyc1EwLOH1t4JB8m9+9T92wxvjwu3E4W2z6k4WrvJtCY2CxF5+zXG9u4QrKT5
Sa26+dpnNozqcBeKsnvpfYomy9KeiOIKkhsx8y2X+1xfv5RVw9FBTvrDW+80RfmQ
daIhxiMgp5CDtxbJYJD1N1HSyFyDmnd8WfHi//biaMNW1VGOxxvKgcIA739X6ESJ
npFLbVMhYL2SkRnqGtK4fRCvohENvnFTW/n5Ke/EqaI0uQ4rzLCP8YwhDMBPTywA
Zryorm5goitw/4hNVDQFOY3ede48ODJbUNZ5bNgol6AGwYsHaqFHAMQHsa+XblN8
p5Ah/hA4Kt0igfZJ8WRUK2QWx8aiXN1zuJbX6AQ7i6+5AVecdn2QUbFZtVGJxEWL
/tZtNycXqZXhYfloaIGoP6sTOhC7247rsEfcZz4NE30mtgizlv3bK65cTpXGVynn
wba4OGInqNhaLgf6isVTaNpjMeUwcmPVSeTKYQHjJkLbWTyg+4txWU/dV/xsvsw4
QwyIYlaqBKyx8QTLcPDyOjQbKA+fzSNJ6oT0o+wLq6y1NKy8MvxzPO8SWn+tggPp
6hM+apFTwIUg0uKczkEP1W0RH579M7wlEP9dDFEDAev/GCob2OBMydqQwto5c8kj
2v1igXevxQRO5+g48YXjozrX4WlzhZTnzaQrUCHRF3L1K0qvzEtmGH8+5iCnnHMf
Ic+7aBm8KxMlWd5BcdcW2ilDbng8WOrFQ2W5m/hIy5G8QLUfLHWiI5Cvqo0+17WI
lj6V3TlWP+B4dVipd5ysbGTdWg19dvctyzmL6w4qHg7vbhfLoX9QPX5VPwRKf2oG
/mzXLXppkz4xmBFC3DBf09eDk85WwaYj+76gzR1N4EQBzatDa3g9IgUpfcQBiYHe
88l+6rGPyi1biHSb9wMWUt1Nj5sQQAvR+H4jEYByKfeo9ZUlO7w5Aiditax4jYbH
8m1/WGo+f/8KtT5FnVB58XEMa9VrdfxK7L+HnvC0/yAEx15JrBpNe6lDgPn5Qs8Q
FniqqejGA4/E86khDpqzpy5FSFQmw2BhhWLvGb+Pb2BUHNfMnQl1mR11n81b/d/F
4aEeNqG82zu5prnaITdWDL8jLy3Ffas8npUVH1tjs/jKdsjgKwbiYL66gvJTQxBA
ADf10qE3V5xzCPk4cS8Lv36athIyqMfqJbEKk9LBTdfE8wO0e+EDm/CPpwQd/hE+
at82vzkb1fGolFjI3Yy/d21LBSCpVEXS+TH9krCKmCuOHTtbAJDEHzyAt9MU5HSa
BODTWo6qPnLNrHjs7XUqemwfs4O13xv3oG/XfJ1MBGn6KnN3ihZT1RJOSAgdW1HC
bG2buSydu3h9QTunZ7HN0C8nGzy1unYR7Vgoj6K9CUWHYTZycouWW/uhawA51GKN
`protect END_PROTECTED
