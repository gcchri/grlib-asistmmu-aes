`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YMdwGqm6WnaiU/mUElNR2EhJp9SnM2z5AynlUZq2IvUxbKPjT4CQsNEu2YmIxv+6
g8XZLa5rpjBG0r44uDbbxKfdGwAsmnrB+NxLrL6hRhnYKQtyUnsKcZ1OZMz+PLz9
osXwylwUOW2MH13UewU881oJmMYR4NMVFpjj5dVrsJT61qsEaYwk9KvoxZjdE4im
KmOy4BRLg8Vi0SvifwpAaTtFdU/1sGz6Aw8J3UjldTTeVXwyXOeoI2Mz1a3PbWcp
f1Hlyg34pgfL/Vaf5fH3vC9mGqVEfF5VfvMwbim+daKxpx+Pk9saqZyJCcze7p1u
YFt7wJzWINhM/lqk9YwUPA==
`protect END_PROTECTED
