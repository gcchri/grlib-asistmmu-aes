`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xXq5JsUYYLVRNPrBNa4lRs+HDiJso00Ev2kyR2V3et6ZgN5hY3QJnASDGKgK0yRA
fcdQ5yQrMGGN8R9KMoiDl+XezIHZYVbK3yqswvnzudpHECMaIAd6bi5DuTdkY5XG
WhzjEwu/sJ8IPt4hmrwlCcihw40rDAToez42yKia3vxU94vJBTypCDKohttesxpt
ik5Bkr71S/mwv3kZ0M2GOmiqf3+eTmOa7+qyhGSBUdF8cA63dRff40V3Ik4JAsEo
oGFBf3kG0p7LAUlg/YhcrQ66tCLEAi4LcMhY1Y24zB0S+11zclTxq23XZVfHgc40
SLMuMW1Ck991VkItHF/v8l3uIExlO40pDEBxjnIQOF4ftJt71BwEl1ewUBrKX1ol
3xnqAe50E7oaJS7n8qWLnbaEYnGm6CGnCxiSdGffYCw=
`protect END_PROTECTED
