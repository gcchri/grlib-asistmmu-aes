`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AvGDQCtFmxgtq8Hl1mruOr7277f4CLQgLmslAAoIDf3mB0dgxyUFDtNT5n9Dgd7c
+itLa9UeT9y0vcgDQXuql6/EyYJlGCckrrkEg8LJxuX11UrRc4pv0GtQjyzAVPzP
yW2erxk7hG1o7iJnuXfyZy3E2kC2NDD84XO5dToFi1nhzEShUQKRkeRXQwCBVv0S
IDYo5hG/6loJ6S07I4Hl6yN+02B6ag3wN/LXlhASjkXXZhcZb4O2JGci7JLooAi/
YDgk+A5Qr0dfzDawsBUKpCHMWZeYmtdbyxymfMNCUi1GIiiuRpdpgMmFyLEcNz7s
O5I9SZtaebDzC+FWX39RE9CSQA1XHm1oMEJeG6f/vRcXbmEqTuId1UWojkRZhURJ
fgD/jLfQZ5ABxsCbl2ntJxOHGPmWudE4SHQxz97xfasUr0lHqdb/VrdCut0V1w3d
gX+SiU2vJzhAiHvLZJOIA5qJ93Q1zDjmlhcodAN2yMzL4ssIurReiFQ1QY2yIL+t
qjoU2655JXZ/Hl5hKw6Xo+AT466ycJQTYH/rd9z3d354YGM/6Y8x9LHkBhbNxNM5
+Lh3OPi/ILs299U8qzrufA==
`protect END_PROTECTED
