`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XdkxCjyLkt2FWpudi0IlHEuBsvZ0mC5YLLGFU4f/bWzo1fUbZv+RxbcWUyrVro4N
O7zMV3m5yyDj3BLgswpHQ4E6K2g47dqgRyZmINPr/DLBE0kLg+il1CRn9x/4bWeu
UiwHVzPEsSLT9J//gKOYIgo7mvbVuMti94XFbCVxId2pK9cx7nCF4bM4WVrtvZUS
/oyUhOoGumJQgosgHNYoRHjRfDvrPUTOeLTzhn3P9Eqn9VOZMA8lp45rPGoD6HvC
ExebOtMWrZ95NEwGuCIbANFqZRVgIvGv4wMU4EVTfhULtFOnAoR4pHDtT5eK0hCF
r/nHGy0HSyz/DzYgaZj8mCmGx2mku7vl7NPFWdv8NbBm2hDbspXMJDa+QDlZQ3YW
qMmec9SEoCSD1nEKQF8D76OkvBwaI5b81wj/QFNB4bwnQhsC6mQ4B4DPDj1FOwLS
gz+5ZS08P7/5m8yPifMGFt2eq8zBQom+LltABM2vG6bCVOENvywqgneMkiqKJNFA
mx4hVJjjN+V0zkoVKPJ4YErZP7HE3EHx9thwtuU/K826JJSxSdABmY8jcDRmq2RF
kX4i+rQM1pW4ZDmwac+apvJ/zLS3DAikt+zOL7KEWwWpuFzGzg89dlqO6bZr4ixP
GW6VMqwEOH+MGyL9JURwxWiKcT4oWYrbO/SIztGTAKTWgdNGa3FmlOnTR9sfVHPI
dfcqWEqEdzXn6yEXipvAUz1epInG6xNcUvewvDTTiPcPnwdr1LSaLl9vAQ3oi43C
59yDXQh/+obydCyZvBYnOzfmS7fp+luMSA2ywYwhwoygPXEOb0oycH699LQPiTCj
DsIDx1hD1DlTcObZzpmJ4zsaBtNX/mtFVNM+cThxXQsD1lg7trSfVCDBFCp20rYt
Cc/0DKg/Qe3zlr8HS6uB3aqcNMw+9Pr+14QgdeZSCye3UdPRh4jxjI4Fz8PrEKnJ
drBBgbYEqgv2ZjVVONWwy3pDZEDyDe68TPCyK5/pkUgxgX3YTjuB7D/2DZI3QgLi
Y7ADh80fn3Q9bovgcrqETqeElbYOjIiydEtqWSWg0FMmpSpRvkPwcxrgHzDjSYpJ
CeHS1zOJ3ux3dJtEKRoS3IHflydTCboVDTA2pbA+2ZsjhAJpUYM5d+DXoiPkngMm
BXiR+4+Eqonaq32qvYYtQ7kdrYrzazZffmgsBHaYKDzIstqlunGDCjYddnY1yQkT
yHJtXN/Htf+QYeRbo48T1E3rUjIAjdRFPUql5tPYhkaoN9ijgM3mVbYjmtnRa7CJ
2Lnm1hUOBtJbgAyxXKLJfx0Ga19Oc117lqjz0ZcDuVYHJp/fn3ZewaPM1M7xHyn2
vJ5OF64CKAL9MxdhiLMVD9HQk2EK6TqQhEWdpA4BHTs=
`protect END_PROTECTED
