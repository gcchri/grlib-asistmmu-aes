`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IrotxnY7tNK1mieOEJBYsHEkch1dsJHU9P8tn/Te6+mnUMZOm5jPRIOZPxfq1UcF
gUIUDgQbGh0JDvkctRJ4AVMSljNiHZtSIpLlIlCsWNNWx40yMaw6Ci6zTujlIgHU
GvRCzuyKavZ3mJ1YPxtPc4naYpOzAG7wm+xSaFTSWKlRYtUlH2U+La3/JJrMhT2j
aVODiRj4v9ZD4KY7frxfh4fXwPomBTsBppUYhXJdVrBSwFhFaQ0cIruqEAjQIAhn
tr7ugkBGhAWbsVCR31+UDq4rFw6RLGwFeiRSyVLxzvlrEVA0Uu387CfABDitWbR0
xqRoD9cAnFW5PvvQoVLMKB9LgaLVa7I0jxtJ6rCWuRTtHVaHJ0/sBjMi6vafV5hH
D5DeBMDI+4P8K2ZUosx/cRkS1qdHLFWIdsMMfhFUdEYoqO0jWG70vTPY9jYK1eui
rtsdcXHSSH8+oCPJpN2sBa2PeAW7c5U5M+RtXS62Ey34OVF4TdH7i9y0ZgNBEQy8
AKCNKtm8W1jl+rtC6yB/YjrNk8g+PWt9X57J5+nq46PVI1On7KAR9RfL1DUvpqUI
FuKbmM8KNe7L9h2EVmVxEqlCP3L0JV0acLPTMAGotIXVLxwEv1vjKoyyl+CjlbQd
OF0upPr+u82O+RCGENFKv5HIF+2VtkEUm+5Ygv3kPBYrYWCLWQt+8xWp9DnU+Dby
yJFce5uuzXtB6xCpRKxwF677OxRIBUu7wB2oIzkmA31Be8nb0S9kF7ElD8SHF8LW
q6rj8OANsls7P+3SvBvlFIXtIcdIOfyq7OpXZE+sJPyOHHe/lcIK/YumASLC+7uU
0puLcDiPsdi1LinmqFED8fgP7mfrG8BzA7E+xBvlDO8uquwlGh+jkJMm9ULvrKEv
MH6P+tTJXEswgrmpXmHyMx8+pjQcgyWXy13SBrrlpmxKgn5epRYbBtABe89N4PIR
`protect END_PROTECTED
