`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HADXG8tvbKT8vNLYlEuhkbfJi1l9q7pQ7poNtEtGyn3AU9hs72aQGFzRdI4bWYFI
xsrQJ4G+EHC/C0T06ZZ4S2pTBYZIhvog8aY1QZeE77GhzB46mlfLjn2BDAsdoaqg
x1K5ZUPuuKF8gXPDAxBfpgXODSZCJ/GZb5QLu44aBHoWvN5wswKYY/hnnGKcPm34
LOewdNJNUKIaVYCttkWGmMahPIZu8mzP4d0YbfDTRRGyBWjMYDNhqZ9lJ8XXjLW4
LHHaNvJfmTJ02uHkrSSD0zne/pW+GFhHEQFjfDsvD9Bg8oM4thtWOBz9+FKVfzgz
A9huCBHwKEnK9s6VmooaWFEEp+ZudgBZx/GS2Xnc/+xFrnWwiECrbga9a5ok6nrj
DFfL7IjxSAr4IN0AytusNQet16kEPousPFYpKiEuEGzUp+Jd9Fq6t6q6j5N+imzE
1utCa26x9INcBJI4IsichA==
`protect END_PROTECTED
