`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d7Uc+YkxU2R69zlQT8t/fw7OxWQ9jMvWdIZbd2RkKwszLD5+Kh+3Ui2Zw2iQjaJN
dPXhcknm8OJfIpeUjM1LmkOm4UdyxdYFE7OVkVSP9XC39bato/k1Q2qU3jIfHjhJ
tiEbcgAp3Y0UiHW/glFmJD+xUHE8dvtjsA0y/TjM2sjV8ejK9WLN4xr+6WwCfOsW
+X3SsGwo4onp60NVBSdCAiL1IpZc1wrgkuy1jUw3ENhkXGsSkuWXvyo+E5a00Qa4
ltQfSB3oVRbmvEAVKWPg3xipfPiiaZUJoBpVmXif2DOWSdHkeuuIgesHoa9IxrDj
KBVJmCMhYMsTUXr5zQUFKUqKsuxaAupkWic0KW7yxDzDZhY0fYskhdq0zCcq0IJJ
Lf7ZD5hnIZL9Bbs8x0mxjOSH8w4AFZYHPr4KoaPiZuHJ5ZhaNhTY5BYuZVgHwoUs
qI91gO2DDacZof+2HS5htKFbmjCu2fBt1xjdr9Q8Sbc8QcCMfRU1Xm+aZryfjNyY
DN/VEorW/hl24IPV+xqNWOmKqYz8E0d32tz229ROzNGW8XEBEpQHoI0Tjqz8IUBF
c5sjlVdkofwxHVzdyLvhu5yDFYLwyxCJL73gbHkBtrTGhm+L6ezNNKbSZK0qp+BX
F1RnnQpfPVKcUJ4nRjIzkRxh/UcSdwG5atOuDIB+iw78a2ehI5sRUaw8IJyyuixg
2jU30rfoas+2dHrc44w6Zg==
`protect END_PROTECTED
