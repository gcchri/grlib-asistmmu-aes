`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a4/EFISFsb7WuPm5H0EPinXaVBIr99IDLqfXIEp+hvr6fiTPpn1Ir6ca2PGK9KUq
LJaNWGriutr0AflYf+CvzV0NGgSu/XlfHD9pWY3neVt9GeyCVeEa7XMyWAC25z4y
DxHoK8ll/xQCbAUrQxpAl/NO9dEgOXMSP4dWmzsy45hdeR7qnyyR94hdL7/ThjQq
ac3/pSwmiNiIdCTb4PDgDnEm2wyR1lzMPKnOp1w6DEp0eCbT4qs75IKwwEJjWOmF
pv9I1UiNVY1teN2M1BLaGpIf50N7FqyZ9oYRQSPSO7Ys/0aCfqFws/rB/IMif5vx
ZkAXoTKuPjQh1NT/ksNPJvE9nw9cFlyLgSYLsccPMrxG9oe+RxnZ2mUP8mEFANEt
kuMAhfJf0Nqtmuwg5pNhEl1wmw1s1diIB0Z+CUJO8Vf6PuJ1NDR0aKddqZ7nAIyy
`protect END_PROTECTED
