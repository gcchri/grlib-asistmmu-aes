`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qaYJdJ53jJRskCE0Cl8UEj/7NfBK+qhXBDbmHiz7ARqd4tkVF+DXyqwM1fqBS/Bg
tlpxClksjj9gJKtKmK3iPSwnPWrUPWYGSsstMav3WW4oNc5YrvtMkleHZ9ipNV6c
ktuJX63npZwnUTDFtUbDDV9Vwn3+R621/a6czgd632Xjap91jllPaOojcFerZ40+
J3HEQoVK2CyZ6yMLqQM8Nc1hnELFlRiNK17X/vb3kYfKnxI0DrePca4SVX2tZ9sv
VpBmCnqa7q6U5nmyhgG0JVl+O12qYyPxAE6sGQ7VwpIopku4SwHFXMB1EuwCtLT7
SSBx9blIg79OfT8JRe7dGihevjQSoCZNsNwIIjH/DGAWAL4qOGuSUBmWcnfmIgNY
PQvMRrEkbQ+BsOsb1cuY81kRFPiAsZLcvVTRFoVDAgtPUxC8hN6/bjJWf0BCLb5T
BcEIZpL7c/RYyjue/wfuPG3ReF0QzqFwhda5fq8/wmY6HKOk3WGQ+CXNIsXTQgn0
ixnj016s+jyB2UbjFwjOjDAWfaRk0Sm1dyxBE5oiqENL52YdXz62PK74+w8xhqmV
SM5zRyThIe95yt35MMgOsbVbD9iCtGX/CTzG/kvT4fdYyZvRkeksA/asembZhuRf
Po3+B72yTeHk/dn8evXNCd6K34TPyohq5Va77veLrDt8vlfa8WAQmphhsDuR0A5L
GdCQ9nyR35T98JkwijnzFBOshJ1sdCereiCVLGymB+y8y5cP/maK0Oj9nF63ZlpE
fajBmRtleJU9yr8lakgYpIW9nbGe2iKZtur89ax0HVQCKso8V19Ux5sqO4p9ikp1
Cvwi/NiIGs82Zbb4XRboU8XVyFH8f8dGzOpJ/c6VbCUFbgzLMImMnm329z17bIHq
KgY9MaE450z0kPBMPNR4esgiHRsyPcwNYV5FDCtgbjRzfXzZivmtc3wGTgd7Ec4M
KdnJyAxESr3gqB/u85jOh2E/RInPHw0zC/Q0MW2SSiKyh5LQwq8L7pjNDw5K6c8m
kzX6lxQz5yZVTsGtu5tqBawiJLQybk0ln17l+e4Abg5Fw/Nx8m68Le/k9/rpl3aK
/Lzs1p3Uz6ovbv5e05dcrj9hrUIs4gFnj3ttMn5HegSFyi6bXH9bS4S5OeTkeU8Z
A8f4E0Z4dYD7+uZKCLJ2kJWs7OEgB6b9WRJ5jASmUVhIEO/DgvK23wI2geye5yn9
TFJ3Eml1eiHyVVA5lMDVWNbozZ8uy5ClYyqqQk/sJjmNNetj21VIPXpIiOrNs+zr
ddKY9DcvHbGaC33sdyWXzoIJb5oSZYGM6IlHlO4nT1FafviuRykayFAD36gMYjL+
B2TmyMucvT4CdMw/3FA9eXVuFgAMoMJtzV5zgmYkx8MPeRyCJls2vR5l81Afyq2l
lfJnfIW6elobYpO2IdcppNjOgz+w8CXTTD86ff+bin+thtQ0qXJWV9Mtg9wiB3xq
crs4boL9ep5B0Wf2sWsz9qhKYObax4zFuAkSCOeY6UbZtcU1G8uFB7naOHnKu6kK
w4cItZF3qo7qSaJ01NUAMWHf/1Dqqx5J2qL/ttsLwniwaREVBmksl2xUy+OclPVu
V2X0c6lqG9y8Z3a1GW/F2AZ8KGC9vIeR1YUDL+T2XRExvtQ7wwfH6Pkz9/HUOOV+
HzCmGVMNm0G7E1r2iDUKuovnnVV9hO9bEMc8lCtTdctlr9fmvzpjs3f5qUdX2yFV
ode79Zy5QoxjlJS0BdBsyuXz8j92JiE+TtdXSQ0D4Nw2zQ0RONRZ/sF5PDx6uL86
DOXEvAC9LGcq8sGWSs6PgZNpCBAeisAdsaT0CS2JB/gltZzKdzJ7TyaNhiKbQQJG
OUqLcX5LHeYKB17+iv/UJQs6D8rIO48WCi0htHlzQWl11V1eOQO3K4OFsQdDE/vP
T3qjLQGY7FpN8faqCIjADQ2XwC0iSJMvPNBga7zMDtKSN8y7+hX9/dUEpxCo2UTx
/yHoys67jACb0NFLoVIxVCo/3lBFFTO42DS4YzL5QramIg7aOVPzyE61zKutkPvc
kwt7H1cDodgT8bWv38VmfeWe9BAIlUnziSlzppbJV0cZwSseTNiR5ldX9oOBYNQi
8pmTwpmCRRrogY6tJg5qeo1trebZgkVC0+1qYOEU51sCkGde0HCcDxhYypyhjKze
x6dXLxLPLS2byqfI/ec7I9b1+bkwaefVEp8/2g9SfDeRPKjCOwKODU3KL2qaiuY/
zUXDCEZu0ARPKXSERjBDMjOVcup1khtoptiF13/n2vcgHlm57D2Dzev5nVomrrTl
6vNhAkWjZfAkvPkAigwP9xQlpg7C3saJoUHKxqoWf15scvk62+jK2urBTaT8dQlx
sCANud1bppgJGtXfRZ+WU9qpCfoL+5qKVbqG+QyFS8szpCCGYk0yVIgvmvUceW30
guqrtoSlvFtJPWnPNBHO3KBQWahk87ix9paezF2WZBTcbHEgvLhRWbmfEOdxnp8g
1+tvROHd8j4wMyOqlUXfbiFLQGdCYX34WJr7iE9uOHWs2VYwXJCpUuh7Cf/N0RBx
asBG4YO0IeOu4LScJcqYg7yJrqgYTyr7YZpjZNoaLcT+kSMisjqdTRNHPKFEPGOy
+/2VU/K4UH5aSHCMn9IotkhBQoDFd1KQE6cyXYt3sgI7JhOT3wuxPVwVngSmDqN8
YQ8vz7xr6offjd3XcZn1d/wtYuzctQOKtf4NBPi2k3z+gJraI4sVka9Z+fcKPDnY
p7mVXnX7a8Mfajvu6HD+/hVXlbenuYaaJubzUGPIOmm5WjcIk5Gr1E3UQSfToiXa
gxx/cDg8gU4EwC/wut9dIwiH5O8//SbB+tmuL+qheVZzQ8qn7kuXL2TVUBY10VvC
5Nf/QgLo2KqBaJ7iwvJaVbj0NiQgznTQdns4qB+RNCsnjMzHYdkIS9eNbn0lzZJ0
EzwkSZmVW/VgSv5RVlG3pVFAqgBM8nu2JXmgEpNysT0=
`protect END_PROTECTED
