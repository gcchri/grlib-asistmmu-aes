`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V0gkYKTIEjLLvTU+LAq9UWg9mf9fDbTwBUirJ7iLZS/tn7h3p1BCo1TbvPL6r83A
lDbcJKNNIDcGacUx6hHPhn3J2YgGfIwlGYnc1oUYZ9eUJucgRcLm/ay8DoPIIDsP
9NlPmGIESqjLGIToTSX+ad35bNtRamhzM5xlODL0ztaL3ehgg8KU5cTo6xMaj6K4
AGXgLdSBxlYKGdLgjZTJExjBlh3dkjVpiMX2tl5vEB/6xrwwd7gwaiJZFjgJg8aw
ZCuXBU3tNBdxni/V/D8x8s7GdJFy6RrP+otVZpuU9MxwhocaJFtho3XSl2TE4UEw
D9FvVc+pYk9fXDQ6K17pG8HUpknoNVZgutwgRKdg8AL1i4X0MWOKsM8wr4d5lEMi
RFLyEUTLUvo+INdH+nOqlZlIAzM5x+YVnDQwAelI04WX2hwqB2qlbS7xp+uW2oaS
eYvhZJfbgTdNf7hMY3ctPUaNWy/od7/T3nJmNc9xANk=
`protect END_PROTECTED
