`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EXRjtwAjySZqE0D7O2vV3qjtikZHjWTqeVutQ1UHkCg6DyFLDaOwaSb/PUGZYtj5
6wbceD8SEl0VqoCzgq+SADGj7kM3HnQnjjObmNmZuGWQBEUpevFUJgLNfQIlfYYX
fTGO+k8IEX497jgZhmxZ3A7Cg+RFx6lJO+oe180PCrpWfquAnBPezzWZSye28HUU
uIL7TFadWWq6F+Q4ptxdVIm7p7W70UCm5MhcvOcT7hnwZAoP4LVSS1rkkktYYQ1q
86VBkaWoQd+Ejh+ImKGLqe33//UUp6tLib6rvznD+B79q/8xhDhG8vjf1UiaqTOo
4csUWzrWyp3hkd1mdJbU5kYy/4FmVbuTDORsnV1cLJkIOogLMvE7ZiyVxRQLRCN3
zGlecXSxuzNhC5Gw0eTHm9qz6JF3GjiYJLLwCXIzJJXPH95ruUupG3wGcgf73yQf
`protect END_PROTECTED
