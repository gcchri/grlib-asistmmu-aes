`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OX4mlbuEE+hGF1/RVavq17BjD5n4c1TQe+x/TS8f8pOWJGIRE61ixc3+hRsNgfI6
Jl7n1uTlLqIynO5PxU5HIfGR3zbaGM+yNzxA7GeL34f/iXhsNbhkX7nmuxqndwSK
8B61EPezFf7wrBDbNcEEbkP2AODse6YbO50RKzg2W9WchFtWUFpPv+ETJJ6sR1SJ
Sygv60vdL5hpct+fWWug16VlswRJAEdyXX3p7oTwfZDyxVB0QWnv7CmRLily5hPq
3UF+4iMhAkIY/VXf+h9oiUOhxfcQvgAHBZqnZu9KvryLisEQ67DQ7p7IrRD6Pt8N
cm4qQ/5UhaBhLKVTqA9WEm9gLK/ZJl2+CRX6QDUeyQhUkvcGqnYcGeVc76fGPGbo
vNvgwpGxzE3EjR3ZAxk03YGvoc7iuEH7rPrveG3gCeq5iiMl3D5ilE0M2LA6D9Lo
+JR3W2jwrSXBAVLs98SWaB5xSEOBw7rw+vjzYLmJSRRGxVzMpLo4fsA8RQr1I9Kb
FBVTYQtk9PNus2SEY1FIgIgB/wmAIFhJIFNqqj2vpoFITZHTbAFGxNp3LvTjbuwT
nog4YFNqFhm8vpPTiSk61lKDzF0kHG6ZFUZUXYB2QnQPwT5hGVh3o9Nq4gPCK9P6
cL+Dbr+s/NBrnluU4JndZWGq0ZK0amlnSeDQOsPASSBDLawrDWP3dGMXHS1S/LaF
pOmkyW2foQQNmBW+SpImWR/ZisHZHgotMQ6oz6kO+wAmZnVizPVj6A3PeWn2K1ml
V7UUO5WT91pdW0y9Hr9x4ZLHb99iI6rRLCRMoJBQzKa2bfQT9AyXEQYlKwHzJzSV
cHHR/f1mGt6yjRhO7YB7nOQy5g4VWzjknEgwa4owNd3jZ86TI0GlRH6x1BNjI7tj
5idzuFJXkfGZd0I+bNL78qhVP6qlmmGP5sXvGObMqxpeaHJPjtjF66cKPjF1/ydG
mzzL1hnfdSv+XatWgoRkIQhiFLKaA3gSlrBFqcR9XUA76Zg+6HDf3j5hJ7LyRrIK
8VKkSca4fgX+uzgAsBQMUGtQ+TTC3XhiwMsyttGNMXOxbCnb1VVJgqkRBei8by4F
zFbNvXBUiLwGQh2aia1IKUXB0ZCvpMPwdNohMvZKSCGFw9vkfQXQ3bWnjAqn859Q
yHc+p7Giv22z8OaelW0pH5NpbONKLZve4dG5LxGGQgSVAd/9259rmWclLaC+H8OU
c/nhgNhDVC82lTeT06wpkQ==
`protect END_PROTECTED
