`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8WQkE2tGco+xKoZJb4CiHfSbE23FG1Nv1P3pb1RHfgsCztjWS9U1JrM3pS6fyq1x
o8FGsqH/tnP5ga4FL/g0uUhCZoRSytHa+649iOHUuD8jdYNucgfXeLclCm4But3m
EIaZ7tm1qGe5JajkkTBqw2E3AbQHtWne0FrbIBuF6WRdMLVtMrXGiLQt+U5jSdpk
VRX6Eofz6O3KK1Wi2NQ/1V4ZKFTN7uDA5O3VS15wyXy5P+MZrrAHqlFm8zxZWC5X
uUuMn52GC5G+Rkpksv0fWSL89vxCBIRW597ISm9N+lzfUvmtPYFKLj0yv2DdoKQ3
Gv4udNM2XEP8wdQYfH0WJxwqSxwER0CtQ7BqT0PP5rk23XX3BxNnv3OlQm1brsNh
0XsInKBm3L28EvnKZrMpwFUXUpglucBOG+S+S8zezhjt3mX+mJ0qJqauz/2Kc/wG
Xn0+9HqUSOsq9g95xbn+CKCb8LkWrS1jFqHYSEcXzZqzJ5kjPlFtIJntVFDBQ490
CQtfvYnUhSNMxSniUPvp/NgSs+wI+wl6QEphmNypD1dZnfPAt/GU56EVZbHkS17U
Zj5WjGuRweyF3rv9MU1OxRBGkHHHDazB3CRcZ19+hmTTnPcEJW/D33OUjmovY0CJ
VBWt9k2ee6uYNoqUjCqYsXFs4KGnUW6Gy6+Zip8SDuOAWTZwrl92Q74o/TmOPVUa
HmL/q3LWLMfu9aXz2QnEZq4eDfCCynOA2RjD4YOapgtg40Ril6GF2Flv1JcKiq8x
ye5AJr0WnH3BcUHzdqTmfrXsWiFJ1sdUZiOO4uVOjhY=
`protect END_PROTECTED
