`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w32o8AvG5Cu3YYv9QZzA325/LJBA+1DdlA82QkWVwpZUI3+nTkHpLNqDLc14c0V5
tLt08CzNKBVhAVEKnZ+CSA4y2jnYdMDwR9q+vIREfvaGUG0YBQHM7y0Ttnnxafa4
zQ3tUtGBTRUhzK/oHykybSC6TMuxR7Zyn8h0netTT8Jso9U3/FbnoHw4I/2NuiVl
yyM7shzCU67j3IBzGjiTFDV53/NEhNcvDUlIrd9ve5S7ba5o3mV2BNPUPc2IDPPR
o0SzJC1/cAT0YVIWejQ/4DrNys5Fq00l2kGU2TZQ0IxkU7YmV47TZDDmJSksvy5R
qscr1MaVXwMJ6MODSTPu72dQ0/SBv4IpgO9Gqq7FLXs=
`protect END_PROTECTED
