`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cyAcA0XqX9CLcjD6ncx2ozl+KTG3c7MG67k+zRqT/JfpGHT08/Wx8st9Mnj5eNWz
26LzwYgvb3XSUljG4dtin+nyRLEBvB4Yh5F3zjBLSwmWQ0KVzFdJ4xpNc1awFK3/
bPjXg5eHgY+A8SOET/HkUsY5YsTdvqxk+CcTHOvlkpmaDtEvKr+p5MQrJAzmuAng
gKf3QtnkihHPQ487rbFUCg662SwrFisGOCp+BtcAEKm4frRh4zGgquMolSTkyzvc
SGGX/mrbY1nwrwivy2PHGfWM0g1SPu+vAceMGkA/aUTdl6FWX/SE47CE72oNUctR
xkx67DOnnvjxroOghpmHZbHh3HlLFku/oHmUz3OcW9yfkDU2uetPrPUlgoyi3lwn
7vIjo8uvy2TZ1OzTdzvLhg==
`protect END_PROTECTED
