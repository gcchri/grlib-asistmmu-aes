`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/7YCp9Oc6iSw0rUE9KK2fqgkjOgkh1G0mss0WWpu/aEnv2+lyAQcanGHE96ZcuUV
ijnURp09zZzpF19DDm0xpQwIygfThEs3veDow3brUSW6hR46xo7TS0dNa09tJY79
FCgZADs8ihGXRYudbwO9/s2znAln70dDnSSMdndfRqa/jNb522YY7go1NA43ON6+
erepRz+6ALpOWEBembD2Kwk8aYZJnVaxV+6Q00ipD7vx3kWHn5qm0eEGoevufOVJ
E8FV4egdTHDNza15d9N8waye0kAd70bFNulGyodTpstVlgDYlAk0rbb9HR133BmM
4NpXmRqUzmb88+Ywi9YNm7UoDYBhaM1DULV1ao6VsMUDugGmpYCyOu9zWJ8Z2Rom
IDkAz/+5Q/c8YF61LchTQJkDMjIdZ7V4II8J4Eqyw+He8Fzx0n06PaWwtREeOfax
eu8W1OPmyBHj5yCQfiq7pw==
`protect END_PROTECTED
