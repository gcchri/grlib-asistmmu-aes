`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jwUiG2HCwuX/6bEKLkA1V0YjkMHHZVXpDS6780rXu54fC7qpk2wwP4lU/VvJM9sA
Ih8D4qmCqOnBJSjE4OiXS9rX/9pOYh7Pf4nz7I8HzKBbmjefhw7Wm2vuUQpowCaJ
C2TJZKCpOFXEnr6KIaKZjDYv+nDVUoGW1jGV4h5aIMFzq26ffTEHMYnrERwNc1pt
HIQSgGMDe2EfxRaVHOQEnuBQjEVTV0bMdLo/d3V5P0MDyHNCjp/xj3Y9pdi324Fe
hGEcOfMrevTlUwExASEAdg==
`protect END_PROTECTED
