`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FIyQ/sMp6e+Cy2Pk8yDpfd76uwNJwhVda2K1u+RyEXu3xnfhb2gDM24WLs5KcYzs
GXK3GEGGl5bKcb5TPvGyzpLt5yHcSVzDv754yexjiAEVOF1aIW8GoAXaypWib/OE
K0/7pQhcHJnHgLxIJRiClfKlx6lkPftzg/mstxhixW8qU41w3XYsLxBeUFCgq5sQ
JDHYn28nPV3Wh9jQurHk6Opc0lGFSkFC63Cu81zsxlmAtQ9+rfHoSBU9ZOErmFPf
BM9JYdQZQaD4tWxhE90ZfkZcUqILNJanwSI090Vfl6Bi8EUxuOTHER4hn+po/LPx
CJO7HRGPYMRxlpdKkLHmTA==
`protect END_PROTECTED
