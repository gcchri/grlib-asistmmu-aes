`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6lDyw3xED09MqzRLc78k3KcYpjEmwRN3BHDxeTytbpKf8+nS5NMi1rHBl/MIeVtM
QhN87+72q1pDHSN8IVOoctojAj8DlyWVVei6v1QZy5KY9zqG20cOUOAeIWfGQ2ea
KC1B/+e+jI5UCF+dxwLB9qZTQaO3wPwb6j64incgSH+wdT4UE1Opg3aeCy9/s9IR
6QAvV7DpnpzVNUI8AIt8hxOWMZ6DncWj/KTZk33V/D2wA167sxJddSvrS6Vant6f
GuLaAdBNsLSKFGiavIqK1kWLAbNCe+/83UMP4mwvn2hfgFDMn7Zc8yIfAly9P28l
UkUwpSK5mE+yelfr4SgLyf02qFyjBIzuZ9OXBRUtvoRSGnditTd+YYdz/9l4bwmO
mWutp500WHg3OxsBIt0a/YUas5bVcfJAxFZne2io17QOFzExjm55lzFGJKNF1H4z
OUf/wu/X2MwQ2wRP1mkqEw==
`protect END_PROTECTED
