`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hsCR/QztzF1y/2EBN8zbUaXVinSzTT4J5RUX207nNKmYPmenPkTD4fkMva4S/ihZ
QOkI5BSA1MIvFaALzD5PmgIsLzMOddtnaGOIgKOeYB/8iPvBLsBqmhwYj7ddl/TV
8Nm0OZdse+i6ztb/04T+AXlZljoHZeAahaAYopRESAiHxrAkGuXJzB2ccHJVSBOI
KNZ58ZrO3GVuneh69PWeSVPsIYi3QqAMT+L9/HxQm72pIdn5mSJUNAYBcTGSg3jf
u2Gx2xWHr6aBkdCyDzTkO4DgWVwqe1AU5voHTcZsygpOKOgjwDaKDrGZ0kmlJ2F6
4cjOuhwWjvHAelxpwUt46OBMC2RjjIk0s95NT++oNCvjpzFW6wXjNu10qUp+NgbI
d3o5E5kLrmfqYTdj5KMbwjahHw8wjbvoR2SgmHiEj4o=
`protect END_PROTECTED
