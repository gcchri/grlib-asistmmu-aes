`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y3C+KvN1m2OAK9iXNAfy3ZadvVS9WG60jL+kSdYaq7Tx0f892cDaXw/fWT+R1etB
nr0cXIhoTAY3e3IY/SVF5i9bWTcJvmI+qf7AbgFfnnybnXfi0lZfeJL2oUM0SaKX
ZEKh8wUzTqbbNz6Fuzr5VbbtGzOg20ddLqu0AM9jChph+zwUcKp6sJrk29pcIHFp
qX+H4fYHlXYQCCd2tjvl2G2XCDghq0tCfMEjTF2Gge5KrQdI07KbUgfgfwEzdhIz
M1RU2oBOMFdexob8RT0rVji7O0cu8WQeTvM4nAx9UZ6XYxm9UcUp5WyFkypWcduZ
rE/wbE639p1fVqxqZVNrhQ==
`protect END_PROTECTED
