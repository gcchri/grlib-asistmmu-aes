`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9ulhdx0PhQJgyha36/7n3sHoE2YIHgoQBOeP41hBXPQkIa9Wk/Z3suCtKJyxGTt7
TXh64V6140Jg/3b4dSQhrAdJ/TIAvGkRUxWaRSTgnQDt58HQcbjiIPd2CC1i42xW
4k3Wqdws5XtilFDvL3lpC0XaFe7q0vEn4CpBw/xmU650RrgleklX9PV4iSR0rCm6
ytCvxHBxpTU34VZ75A9AgUSG85mUewZX/lCsnip+72pjVGo+xQpyzBPUENWaobOk
L0VyNms9IBJBBA4XetJ/SVJAb6+92iVfX47+EBwsC0gqSYcZJHpiFLYHaq/HLwYs
psJMmxWu8PaZ5j9ud0aoeIQSMTXorI/QaXkjj66V6kYJi18NO3dDi5PZlHZIpjHP
yNf17sw405HCC1Sq1DKvmOlTZj5fBHsj+ogxv6+0AJUMYRJb0VHgfCwiUiE31SSF
Va3aQzKGzerxdvfVEU3dGA==
`protect END_PROTECTED
