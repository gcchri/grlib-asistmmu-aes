`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D9DMOFcq/K/CKCVsCpdnpCCKry1QDuvd4EQDO+yFQDvRzDN/ozCLsQqZdSJrPljb
8+7D81OYdAbxf0gyGxfVu96vqXkX1Ow0kZagO9zEMGWoXQrpfNiXB5phJOj6nRJf
9nTtK6dmOKFhZiibCFhSfZ/9BpjK29fSfdqTnAGd3pWH+GGmxIX4uJqtKfcNeCvJ
RwVsCAAF3kKdsTXdk2tGThh3cvXLHFoAaljZhaAWcIitUOvGdlMzgQpWEIsLu2oY
Zmt3FcwK1KEuDm8YT5IPv44xNTQhfg1q19hk945JtY1E1gJ8U9v+LWoaV79A4M8/
AiWSQzmoegC6k4tC3I8BbILji3DWOjNTTIMd8TyKAQjK79OyMGguYdJUALzY1gDS
QNAeXFsARbsjtmnVzPKPO7gBTpRcVRrriL2YfRBlQR+gwFqO+b76rJiQqzD+mv7o
Z7aqLt2UMFsJXFTWBcrSKS3m2JGw6lJ2T/svyGtUGKK9BXjJI1rs33iO0H2sHUJy
L418pUDwbXSmzAON5MJcKT347Pw6Uxj7ZJQRZR5kakUVAw+8OfS4d5aewbWgYUBU
u6S4X9k7pEITJGcKFf7uB6O1ABuOvqMZ1bxK7Rmc6QrqdKZ1HnjVqli2vfo2FipI
n2rk24Z8G+Ieqrr+7xQFslEtlbiqKI6a0zN5Qap4AqNXcxVNZaUDt9Ba0rCdEdBO
yxSjEJLs7c469aAuseN+kRcXn8SlWPWKNZWKjvvcD7rpsjGLH7+MBGL9gb5Ubnva
/bO6vzZffpC8fQQA9Lq9dlS77/jWKTDVjSyqdXQGiZl1BDjqzodxLrJ4+G7YicO3
cuXFMHux+3BRuw6H926jXV1KyTY6gkjU7cucG+ZkiP7OSyDXn5lTQbBpOUJsIBXq
icmD1HzodOSws09vF0BgG3ABB5oJaOXgA5N0ecEyBoN/Vy9KsvYCPa/TFD/ySlF+
fBQPw8eyaS3dKZ63SkQKcIyWzJ8skRlbKpyCq7sNHcxBUZotApqOhTJ4EJbVX7rq
XF5iyhZhC6CxMYMWF4PLzGOc/sYvt9YNZNx56XV4OmsBF1qlDHgJoWMkWPM7/4J2
Wk8qL0yUSOYUQ3oC7v+v+5LfmvKLOw4xJXxcKl2LrETd88s9HgJfSrvPYj77g702
hRX5z3c1QS3umZ/DULrrwighyNFDufRyXJqG0rqiuihMB5nyahhxtkMyqSwwWRRk
7M08HnB9my4KclpiUSDYCI57k2N8Q6JFELxFdhC+TDvOSR47AQDpSUvj9jZ2GKz0
CNdKB8DF/xXO1L4mO7S4Bmw21mytcp9bLYIa1OIfQU7z6fIl1nKP39mUT1lUCGYY
25TbLsuyY+k5ShPrwcjKVQq8zEbp156oFu9hOsTUWfMukxzdpGkbphob/WQnyUVR
6MJ7OFKSEnBJXmIj2eCcWLVSZN8Bv8eGEGfRpddp/RCoxT9HeP+K3IzEp3R8uDlX
eHiE2XWZuH86dtaMGwID06gUcKk5dWK86CiKQkX6xn3E3LfRgudtP5RVzgDVxKCS
65Wb5wpM+p+zGnmBArH9JTl7mIXsoCbvyRG3PkH0YlAotINKlqw7BXeil72KBH0U
bj+FKbq3N5WcHV06dv1Iqjc4fHR2gfo+hZcXgXmfpKwgNz/RsX8n6DKj3T8ixlbO
NaQviqPI97LPfKvDE+rbzWmTFL7jDsDP+6hJMGldnlbsusMbJ2QOsN0bKiQYT8A/
5Hzs/6gwK0hFcikrJvxEyYJZwyulI4Q7jKpH2JqWA5G44MmbjGKfvjnvsOvb0A2X
ToA40WL3DWZpN4ZmR9EvEv6v5qDpI8SJ2kktD2+YsMp+MPRfMYRQIYz++a2BWpqM
jrxNHIWfM58UxXnnn8vaqn1hvCz5L/Z6kugM/eDR/kVPWZsNdzvr/CEd5cx3cyTg
5N4BnoA8rehSqBLV7/7frA==
`protect END_PROTECTED
