`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u8aejX9TRIJ1trKa9djhvZinJO0EOFhHh+LWF/Jk421h4HJD8aWDm9xiPjuvF4wk
24s/i8ru41v+HmYFFBnj0mgjizNwLTFIXkS+aDhIOzuh+J9Nhwo0zRe5M8sXNhDS
mTxv31MyRhUKp7X4Z6XxpkMjzMcIbPUvzRiv6xTLy9qcksLeRzfkiqVHW0JA2aSD
MaKYSD06QaFVX2I/KLo5KCSf3RPh7Z4plZVa2Uqwpr6Xx2Nf72jQ6eQ5oVQ/jn69
5UMSC2kH/MkNPBBPH2NuUw==
`protect END_PROTECTED
