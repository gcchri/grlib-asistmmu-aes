`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1sqP5luOvU2HmmGvv4XfOjWmAQPe5FPgEllBWcL0VV0iSp+o676LuxY+krY+Sn1x
A5MrbPV+oNnGdl+Tplj7rjyArIRrRh9WgdTNmR9a6kymxccYxsd2q7minHzBX7rI
u+U8g2LMTpSkhP4iXYnWjV+012sDF1AwUn3JM9emrmU+INF4hJ5tejy5WHcTohZW
UL6uy4z+MxsicB/TscT6ZuLz0Lsjwm6ewQ1oWjM3B9jLULDNEk9mtTYsvaL2oX7Z
XhKuqVNjhzhudTK0ddh5STbVwoFYnk+OBq6d1pPR6lPq/EhHCxYw2GH/dYpt/n8a
dyho0tID3qarytvH/iBqCteItHRs7N+p7BdtmGC1flLJ/FcnqMlze32L4/HrHAez
Bhte/EPHp4hPL6zzMu1YNAg7cvG9U6bkADeYYjPSn4kcFuDAnVl+fVSwBMvchHUL
uOYAhCDuzja63efKcbCpY7S3Srl3Mv9FAZ3vYUozx+8sI/wThpPlS4xy7vgzSLZh
hiYG4pAxeVr4W5J9mRC/7/56Mvp+YDJSOS3aJCcUzM2RsUQkPC8fzvDLSDPRy0oD
FlvtDb+tBovyPma4joIKAyt3DDuC5OgfJNW07jpP2YwDcq95LWoVW6Rpngo5quid
vLCTOGAEqVDs/tz3JfjvQ/1ELv1u2Nv0SbJgxww1Y1BAeVBjxqh2IN3i408m+pX5
bmHgawUlC1pITChwtpwI226MZYdMcJiUSx11JLPO2Gta0RxebSuE81wtcaIxLQDI
qtjrn/IzEApe6ZleTud4+R7XlF4n7rpi1ovNchmlowUYvUfajihsOS8dfnUCM/bS
Pd0Yh6R/tPpeq8heV9JQ3/rb2/aDcKwWjQLiyRzujRlMTvMrgze5Os/oP/+Tm8In
RJ7pEr11wQltu+IJRK4iEP2w+c6JfZ8KH/BML8EwplNtkK370sN/7k4F0QXLQiAQ
`protect END_PROTECTED
