`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8U7ntAdr6m0bhNC5u1jwY9HMkOY24sjQaMfvrt/NL/MaIETO38QEk+AOWoXXfplB
kS/VCo8jTslnQgxsS2gyWNBkQEgVOE80VeJG8JqEFBbB7xkuLp++P7b9VxFM8om0
cHjANEwqgYQfeoO0Zu3Rb/FwI4UiobBPzp72wAC1gQmzvGGIJNUWeXNmD5PZ6uqc
tRVWQ7LxiANw9qpBP22IF6ZoAxRtzkqgpHk3bLqiB/3wLDEP8xqofA32YwjPN5YC
WwZIaAIoG5unD6ju+azve5aDIuySKrdpCDTUCWomIz3Qlsa4OPtrpqSRaNzsVbNg
6T/dR6Xlb0JBKTH+uKwZVPdn3HfsYSkdVC/HViFMUAQPJJxOcZTedk/RU2QKZcO9
O2sTInJiSFRxwIwGG16ljiZ69bZF1Dol1N5sQbGfLINq8gTx1wMmlJlMnRDesH3+
xCJqel3e7gv7tbdrLk81hcAaZBGg7P/J8fcH/3849Nt5XX39Ipg8xn3Ff0yZvEWG
x0l49Zbvxjl9EEjTCPpb+MlySnGBqyI9g8cCQqwr06MLQxAvJUmFX3mSKfMBqCjv
4uRUdlvwe0p2ojKYwSDbun1vTcO6Q4yb5uk6gDCkXJdPz/7thE9bWTjLC4hrIx1v
0THxTJ+uTmKxIlRbN1oAfjq7CaVpxZa2iJExDsnY3jrhepQhxx4Ybg4tBW45JV4d
iEd5elIqTfeDbAQCWYjJtQ==
`protect END_PROTECTED
