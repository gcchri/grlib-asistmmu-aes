`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E0/Hm+gjwun952PVtSJ3y8IXNcp6jBiL1jV9htcCdH0iKkfZF/l0YCyr41VHEBCX
jAm6LRKk2S8AaNsnzX74SfRoBMPjYguRuHvW+vvpxqtSaVWyitGYoRtOp5NTuX+v
UZoPH5tL4Q+bmSYvOJIlX0+shaZc8hSoEFHZENxsgbm0vumN8R/MnDohA+q8cmvr
F267wqDswN7fsx6S/OyUlbwe6vCWRPgc1F92ueo1ctM8g2eS+NqDJxYA1NCm4+Qm
3NE7HmRkzNodOWYX5qecMKfzFdO5UoUf03CW1okL2mOlWh9wA4RH8gekeShVHGY/
IUlXBLAPLzVlmraVTgG63UFfEe6TiRghW2XkADws04jpDD/DTH2j/NN0VeskBBfG
G8Q08e+LR+YwDcFOUiyMldZzbnoKHAhUwxZFVkYNWXd7B7bxiWJ4D0aAvpkcTyJr
zOTKMoNvnSTPSI+vHUVrmq5iZwCz1yNHCzJF3IPd3HZwZ0ScjVRQUhSsYlnJSI1Z
`protect END_PROTECTED
