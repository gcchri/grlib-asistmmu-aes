`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6RLTFGR0BN6YoqkmvUrL62OoGDJHn+yyom6KtDw6mK5egcUI7xFArG+a5qTZB777
Vy8TaUEYM8A2En/Sl5zXtiBv50JkpIKvY/Ves0XyKVbfFvkzN49v0EDhfDULuPn1
FcUS/27xoBLVDm3BYYTw1ABc1LZL1XA6xvMvQgqajSB9aWFCefEFr3bcAFh2C4Fh
rutWjpEb7lWl0ub/qXu/QYrAkT/RP7ortXyS+49qufIqd6+jjVRJX8Ff8cdz0G1f
PFu2wIxBqpLeB5qPdNcFvZKveAqlz16JKEP2YsoeZyrnBrrStFdX1mSDnBJmO7mI
use7OJ+WZKTt86b0c6Q68VlyUvZ77Rm8CNwPiZQkldubxQSIB6TVBSlOhYo0wpj2
FKyuiJTncQ/egZ7fnDFcpA==
`protect END_PROTECTED
