`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ya5QUpwlKXl+cadM8WUD4GR6npR30FPDtwITjcce2kI6ww1PAnbc/il8Oyk8y6Gv
URHKGeVCR7Pe1hj9A2rmtYVLnnRovYiN2zSrNdSLENU2iPZnnSzFWZzhm3MMVoX9
VFWjut36X+opqxa3jn4zJ2sxmzDYkqSxh7Hi49+QgjmAhv9fDm3mz6YyrnOya4WU
mOL1tW2bCP3IcW7YeUfifvxfyY+/T3Ipz4Og4spHQ7EkzGRb5/JfXa62dO0VFw/O
PBbW5W7MKfDZoz3hEVHSJSZtxlJiiUNT/7phyTNdR0C2FyKMDoZmOOGYF1pt6S+W
fgIx5qvbAXQYG4xtWhvTBdULmmVSNZDetxUzgrAOt1gKutH+P8O85+sXXpoN3rnD
olSlMFa0sYYPE4itetGRyQ7oph6MoabqZ6xZ+GCGN50Ks++rNrX+5LbX3na59Zes
4G5ohxYlRmB0kbh4MZr7sa/Iz1ZhXdX+BUvBH1B3ddh3i7ajMpfhYG1/AEpU8CV5
`protect END_PROTECTED
