`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QJ+V2ML3Y5R2t8v2lTtGsAfp6AoTSnE1x6Ee8A/2QCdkYCYYzd5z80+gkbZqUngU
a/L2ROMI/k6Tleu/GOafq6VjWqqhn3/I46/PyTmJ9ZSgeog2qj6/XKdXKTkNq5m3
IrOK1Cj7/5u6JobEmx/CegBWnzbtLMcJNdnXhYwjoZ6BsuiSGdQTPQvZTY9c62RT
8u2+mPS9cml+cYpBfsqTDo+w1b5qbjmp/4EgOwkfj2xRiigbEDYgikaCMzZLqjjt
TLHYiqJqMTBIPdFohCuad+eEIk47obfNMcgwqNzZ4zlK7amT47FI9+uXfxgmADTe
N4s96zzd4LpvEsf03uYk097zy3aPAtQbqb3v1DjgGHozO1PKIcDkd34XCDgLVj1f
VTBkF8jsIMJyru497AO2n0RzNreucWgxjQbDpcBvyD9wOXMwxid3cnk0O35ZYuJr
/OGlFPs7tvTmhmq8wv73oUTo4XbydFSQyjjXa5/jMeALkMDXyAIQAmCildTP9FG5
zn2mlhxyyT+yxldSy/39l7MuQc4dP6XzvoJLxa+8vMQ=
`protect END_PROTECTED
