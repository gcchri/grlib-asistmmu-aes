`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Q+nrwd7D6WWGCGOJJR2QZH2rUct2r3nS2ZxKHj2Pk6RQCFc8QTO632FazglgsqF
bvW9DOe5/+UpYyEW2jns51oevQzNxQGTX1ah9hvJENe/g30WDKlKY9KlruuGfT58
osIYNdmzO22w1YVdRgatR2o5SNOdR5DcTLdPNQFfi6ciug/MSELYduMLHJ694qtp
K8Q2adfEnpDvGAWxrGibwg5G5TwQXoQJuKqw5TTAPSZPhh4GTi7DEAkN3J+SLJUu
wJmFMOst33GfeaHk1ccezTfNxDwGQIl3vT8GQjyzC1W7VG6frA16IzudTHr7wWkj
Lvxbqh5YSWEeUuvCa9bSNg==
`protect END_PROTECTED
