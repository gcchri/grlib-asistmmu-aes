`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o+W6ErR5ZJwtiCWEwbCQ8ynlHFxrS2L01Iw8ANz+hjPtcgvOMbRvxHwZScwXPuHw
YqFT4r0cGYN3KVP1BCy5UMnbPIiOwsZQOb4OGUc8ilzlGTvaZWVMv7LLpDNQpanF
LASZQFWMUZ9rP4mbYj5EVKlU+jup97Em2ALd2lYT55Ea9Hcb/8RkUvXAPeQRlnlB
CqTSElIV7w2sKSPX6D2oUUEXfXJRcsYqfSw4CLJVXYhqgd2tnNya7/S4PzWnr0FQ
ywOeWhoRv9gjk+a5pP0d5x6mFppWOrAZDShtnW1OOHf/OtTyAtbLizO0cuIUObkM
9XcCcyOeoIiE5lqrH+QX4tvn/7KjjRolFCKaNaMsuOEIhcS3rODE+ES/Lk/sxjfD
WWWtBDGtbuFchiZiQaTRI1tan0FoMFOih5OjDArOLQRmClswuk4+ZVAJzfBdgAZ7
CAR0PmcNIZRd6YvW5oo4sMVUrpSJZom8j67vhbpFw2XHOCSmuxmOuOG0rckZ8d4x
sXJV879js2IVxvXyuPfDJtOAXfh9DWzVbt8nXJI9bKqUJ+82Qxh0R7jNW2DIZf6L
tBtVPROWuYB4Vfv7Q4og+0MtP0mSc7ooxhHXx4o+cg99G9LdXP2ImSQVU4/oK579
6LBFwfwMPR1IMMm4U2fhCHeaUd+2SDfaEbmR5DvcxJX1nggIIN8LyXRnhTSnMFMX
JoQf/y2xtYfzjatGjKZpOouQlUhfhTpU2JJEiqPZQiV+h+5yjd1KVz9HnTDXrmNf
Po3hRrhTfDY8Fs+WRiI8nBC9Uv+9HXHq38dIZUOR4FaEELDC5vhfRijIufLWFTu3
ZjvuIROAsKDBrvPKjNUxVQ==
`protect END_PROTECTED
