`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
daNDnEYZrGzkDx36IEMsHz/sHM+D5OnFqsyfZeX3uQXRcva/zTmCVcVsvhXPXZDa
Mvy7XGcA6gV/5VkcqpWP2OAiBtXvQqqW3td066lchbByh551qhnuRnPVt+etNyT9
3SscnNeWUdigTh8+cIE2Upi5dInzcUvIBrByXGPoRiThfpum+N2Kwb07Xyzrh5N0
9s14GsLGjEwrVAA+M+CMLZ65rnyUVK+4sz7iNr6LPNxMP8aQYn+mCsWuARq/ozGU
R9siqIrSPZSiw7MKcwde3GH0y87TsO5d0a8zZNtKqrs28DIIPAeUqmJ5tf49hUP8
EGvuWk5oCwiZS/RnX0lVrg==
`protect END_PROTECTED
