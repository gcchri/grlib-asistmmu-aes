`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/9Sig0KlRVeoydr9hLCgfKSPEPNx8SiPIgPz4gxcCXoitE6y4VByPzt1f3i2m8hY
nUF0YezP9SsiynHX00hknZ1tSCs2vCD/gZsSBbXXc4V50YU7fiijLDrxavV5SdpG
SEZWFRwE9fu12OZavPky4N0GwUdyytZiMx+E/oVQLUyQYvr+rvl1WrG8fPu/yrn2
XAfhYFVK+BbLk1KgUGRnKADX1qU0mBq3FCerJQbDYcMI7ZX0bJUvXb5v8/t8KwAc
ueP9KhV0F2GqzPgaSXA90hTK16j3nh660zpbSurLloSxmd29V31oorWbQz8BiDd/
nbvuJG5VXNFT0y456zqnL2yOgj8pFAnjcWgw/xJ2hGg=
`protect END_PROTECTED
