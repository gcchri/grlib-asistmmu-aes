`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/yQIj6eS6tbLKf8VYtO+LCNV0H5tbYTMSwO9O51zd4eCezTunM8UrmzEpeC2OrTD
lixYXv0Wlzc8eVnwKLCaoa/JajN6fei1dRgCYQdvYGiUXXNf0brCqdOww0TbNyUe
MNVmVozyepJOP2b40uYSg4XOB5lHDBXqsfbz7m5t8x7IK37+B9V55p5oZOj8vjIo
7kK1+4u+I9o4Txq3Wgx3FtHUfpvKK853eFR/XXqWiDZUQCr9bV9ZA+zgu25KSAX/
y66yAJuOwe7SkkoxMtrqLBhM+HMZTEcwx2Gu7lm/RVeId20GqFVf1TupyXHaXUb/
0IOGZPYuCKXwT95mq4HrQPonLGwOaaa7+W1KqvGkBhT7TnGupawC2H9o2ge8EldN
IRgRZ72tRQpvTx5qbp3wBuNgxPFIaHS04l5l6EFiRKtvbRoURLYMwImaCW31b1PI
i0HZfhzp3zv5eFMx3Te0k4oLQADI55SyRNKD0OCQ8X+IvEn6GIs0OOW+x0sRfUzs
`protect END_PROTECTED
