`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L+lEt+oCNl2ukMPQLxI3Vp3NLaHY7VjRu/iZepkjyL/ImRn35ikjUPFESyWUP+d8
iRBNfEM1OExAlnLxDeODyvcvS8Oc04xzlGAIcMjQYF17oQCnj7W3GQgq6bwI2/4z
8nUY+p4xMmIv+vpENL/EsJKxwWyCAA3pH2kaAfY5oeA2Es6+56swys7lAECMG4jp
5yWJBqbEqVU+I7AFncHjCyNb6YSMukKf9n+Ruw34BEYSuYquje7vAVknH+pbwUGx
vYCf1xGtshYKTcdHMI3sROf7Bh6ZENj4CbZN5oO58kEpmomrjb4fz2e9kY73oD4o
GEMOOoJmsRdO7FkMlRJOs/Ow2K5IP1+HZ6HMHxzs/AyLrVEJHv3m+tGrexH6FAaT
nPZLtKqKd4ZsGsK2j45Bg2Y5w5d9Kt1UAAwLRVW7/bA65zqoWNOa6dUwlkaZa0iQ
TrhFsVBWi9rBx+LZ4sDGVaWsMCx/4HCCcs7D9zhWsNJrNq2qCacUweUbQa183i1P
gJSZ+4h8a4iA32Q9lh8LYB2ULtXJATOeocUpS3r9bVZOhUHcPIP7j2Is4n98wZtq
px4zJfOTqP3gZibAKl004/015oYK73iFnRnR9QypRQNhVb4j8bBi3ahjW2aYh+FC
LxIcev78dXDbUQ8g9b1+jiXQ3vZhRksPHMs8AIc600X+YX8HHj7G1idiIvJFIvHf
nEsklyTOIrRT3WtYU9GNnHRZqasP4EmFhWXkp8CQuecAL6w/Ib8MqIVUnUS8ExHV
QDMwz1M2Hp1QN7r0nzZqvz6FoWL3CMmEKDT6WpgdKHvbdY7t0EG6tJqTt4bkUIEw
EymLWOcZb8c7F7Gj6BaaG7gBw2y9bnPdfaVrz6d6+ffX5Hy8vWUYjEQNpyhLTzom
zUk89pHiLA5bg5rXyd08JT3ujyvYmmwXEFZaUrvdZM9u4d1ZJ0yQrbMCJ0K1PoGq
K/wnqcmzF1Gnza9BkhiF5k1aOYFzR9wIPPf+lt1x7dYwxafQ5yDlxx99dC4HAOz4
T1BR1zvEMVXGvfRkrCQdtu5qQhvIwdGcIMsOLyWcUCls1MkZDi/4hlTU4b3RD7N0
B4Q01JPtI5FQxGOMAjZTWA==
`protect END_PROTECTED
