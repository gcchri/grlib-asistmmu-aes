`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K7mXhleSJ72TyNS1xgpa4+khGjSq2o+YTj7muF1H/FEiCdu9u5/4saQsCL9rdVNQ
2hp6F9j/6EC4LZEXWHwYPCidca6yLXY1l5EH763jvvPJWkfHU6ex1jWh5Cihey4U
zJ1eQ7mHLdTJt6dUrEpHrC5teJqU3yLGRTlvuB1xyOjjU0WpwzBYThMj3zEcJMRx
N9BJFyiLi0/u+/5CD6Q3GZYmFbPwH3YwC09hKxzzeVGxOPrJuq0B228qlCeZ3PBx
/6ynorurAFT5NrDJD7vFsDaPAyeSXzRNDXmbYt97pJWxsedWUpa2TFGB9H9DOpqS
7uKX1ciGEwiffAV33foy95EbeT8CVkZC2SzA1YvknLrsVAisyw5FfYPFWMqRj95Q
RtX1UP47hZE2ucYh6p66cOsGc9HVW3uY6pSo3f5CoymujugAewtXoSE5y4/z6KF8
mYdWMJZvLn3IX8djrCf69mwDyFwVkb0POF5ah6d+Mld3QCt3UgGrTw9vCjSh8nyv
4+6hhqxiWtPvV8OPkdZT7nji77Cd2mDW75MaXRNTWyFT+u7j1YQ+M3lnIomog+cT
Qu3LtPcXtjqeotjJFHA4+kc583Mu6ZtgW/NAe2eW16WF02/GeyBEaOfwb4cVbHqm
1yubBKbughGinzbn5byqQ9qFKC9gw52/1vY/xzjeILL+LgVHg2OGoeRQQ/tA40Ux
cR3nDs3qPLxrM+d6R5mhVRUlAFWvkMXIW3yXR+6Watq9C5LcWrCNhiJ8xmBgw3Hr
JO216BXfRHJS6wJ7YZYZvvukvOr2UvB3xnWpoDMaxnw3pqObOq/d7DXXgE2W0onc
FqWxgxDsKexQDXwnI7zXKeJO86Slxa0bVeQBWM+mP9PsiRYguLsNumqlSdDJA2An
o68wp+Ub7Qf8X+CvXEdEtw==
`protect END_PROTECTED
