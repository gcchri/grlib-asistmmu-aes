`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s4ixD8v2QbCma1Nqlyl+HLIEtAFC4WtrqZF23/HF+Muv+i62igpJmv8zePG+Uthh
blHBRvGpH39l4X9qf3YA+gLpvv9pV4A/ZzYMJXS9Qd2hJAhFZhiRInGgv4w2GrXY
L4JbYpXyyJWRiX69LnKLKkXKfppuxCkqIogGVrTSquSX8zq9KBKncFtgt4/rdDo2
fECY4jmzhlXVIpbY+8UOTFG5GLMQeqzLVmZ19Xh21AtAItW/1pFnuFT33zjnaS90
HSVGvukx92SqgSoslkx6N7PXtJsGaLPLZHcpbpougPmrqUsdsQKOpL2SvbXidY48
K63ID2hJBLGP4aigyBqOSdDlr14uoyFZ5msbQ7psjtDRTCETa9lmJBdJysu7opMb
5dRdTtkyLUAHzjDw2MZWKOv6ZaW8qoAnlZlP5ZxVfPOYRra3YOL0MpOnooKpd5Z1
sqAWMLVgz5Bj5aHANBHqL9uiDsLM0LxfVISefR3kvw7m//QQZEAxUzqVvCDEGcly
KwG6wZpTuH5mxOg8/+vVjVZq9YUh45Mm970T7XWGODxuVLz3l5llFvDm4qnXTvST
bK8JyGCERDkZ9OJLGyGmcSwSYNlTQLdMh3i343LJMPlHcwLn3gs4AQBTaWz+ASFu
Nie3cIqrxoBTWdyYsr3A316yvZPi84jWRAw5+Z7Tghav4i1bFmT7YS5Ydyw1Sq3K
yelG8nj6arnlWRwy8HNDUmljCQHrGj/ZFWjlMMXueV0wchSweC0R1CgDfnH1n0+C
KX4Kqggz8lXm3wckssVTrNPaQ9KPLA5Me9gk5RH1BNrVxNmmPDXoIpbJkQ/BHTEq
BXB2vrfIO3CwQPhlDZC37QvgciZoMj1PNkwtWd0cRccTjsRhoGa9j8jvBiWQZ72j
vOvU45nwsXwnNa5Wt84epqVeyRFvTs5DV494lPaRDi1XkKHE01p72qYNEDDsl1Pw
3epC77kzaLvM8EGn+R+bong8aFB9lXHa5007+Q63wGVs0FQmzuclLZ0BfAAG+2BQ
NlwIKY14Ej8sZPOti1fzhIMLDKpBTPNJtQfjH2qh5qqpAI2aCy53ggBfEJyTB+0x
rOk+hNYWHzB188RU8Ek6wB4y2yoKLdx/OTSZazDdvWwiKx44MZHsEMXkkkCTQHBO
eLQePLjLj0F53Yu0ECWENr6HT0II78Hj8VAL8vZGyEN4WqDX5TlQO3k1Ch0GTQqn
coI9xXVv0BLlDZwDpgL2qSQbk9D9LjKrQyXvGjgilvdgM4u89UsmeUuAVSt25Wek
3vfYNUiat4UMnpU7R391k6Gb8NKRv2r2HRJ/CILKXuFgbea7l9Brtb2ILSjyy3IU
D3YjdMu6cpML6Tg0mh2bXH1xtRvQoQKbwRmFXCzte/A25V8pzz4XNZImVg0q6NTL
eIYwB4IsZMNUj7npzkxKrgbpRwm0FGFUrPOC7BWCQtKcZ47kMx9g0FPBjMvpl3ev
Lut21aRlLv+ieYlJHSmfZSUoi1bQ3rbjCF6cuUzChbJNodEFloljibxi2bc+V36F
OgRmEIhKFrDVMppUkW0RhEL+DgMq+HuIFU0uXgOAfz/1YKLf9FI/M3jV2+uayanP
QScGnIwt7e2i1ki77/5cXgJq0ZBN74EPPjx5R9g4CFKsYR7axAjgD72qPQgXFayi
QsvP9iCEXsdMf9WJpXsekLGJS+nVw2inriFO7Y9Yex+cDx8DKI6jcZX8B5SM7O5r
+y1afKSqX8KFDe7hZY2uytyRJ6VJ5ueefTIC4+ijiiQq4ejdZP5CI+bcgTq23xMz
VUFrrkKGhsrQpSbUwxvEcA9R0VItZHZcirNMAPO7f9HJ5XTFxih4XCO197qU9aPr
l0NrRsaN6XEiQkpBUe+2seTK7EFHBEgW7KCE8S25OeXGVjJxMe4833wIen/qMONY
Y/ejrkAgf7Kk2+MlDhpMKqziHXY2GNCFG/+RVny/cPGwPyumVRyogL6/XD6DiRF/
WAIRcS1zP4bD1rq2tS4G7kxY1gXnLZhbwWIWByXFUU4=
`protect END_PROTECTED
