`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e4GKDxisC3ORWJN8bYgj3rIReQb643TrHFp9Kp0GqH/J5FTVk/rPtCgKoQ6X4btZ
ENSt8CobLlfqS17wfSrVP28dFdkdksDcNtprqaFNrSm1k1U3/CFMnJo7xtxti2j1
C6hynVouUp00fIYHPd8zEfp666dHSyHKVQVcP/2ORkH8VUQeoH98uz8TxDh/1hy2
K68uKuEYzOc/lG8l7/J6VyFIyZUrf/asMZymjMdrzhnhDq5X87WftsZ++jcJGxZ+
uwc1hxSWuWrU1n6uoGDYePoy4uI7do1dHeSTUzLwEnQSjyTV58cYXhW7BeD3zxvc
MD56fToFi4Z6/cITh7ba+ZIAwAsCSrY4pVXqhtzGa2Xj3kMK4eDMAJSn2p2MNesU
S0R9eS0XZXBoTmpaYawfbuGJyKajmgtiWAapU7biZpA=
`protect END_PROTECTED
