`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ffh5UkXg+80HZoRqLS0uPLJ7Zv3Cwjq7RLGqVBEfAFhEJtokmo2ba9ZEYKfNptP
eBjByIuICk8/1Mb93q/81P694RUMPwqPW4rDSkIf5rcOh61Cpt4ylJtmYDnMomRk
4IVBL498cQhTqEbNyba2rWGUYaRCA/iY9zZHa86M0+D0L3NeDcS6eH+CR9nnwf0p
DutzbieYQKDmT027K7Fb8eZ3pegKN3OXHYHTCFXnanSxWi8hlY3muXecIPTa7Eoy
jPhGaxLudRHI21ZWbSRXnOpOvLqwpkUZEwsmde3loqhVJWG+LNV47gaNMRE2eyUo
77BC3HDr1VrVD+sgkP3H0gTbcg6cBMoi9fz0wJUvDRkOe/5dVwTB/GC7ZLwpXYv1
NHXOXx8/j+t+6hAq9LVm9ZeYZ9ij8AYwp2ddSwAhYMo=
`protect END_PROTECTED
