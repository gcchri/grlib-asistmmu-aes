`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WICQ1O9HTqbMVVu2F6dTSfzzIl9B4TsGmMetzc7MbeAsmUJwXD7fcEQIywjqCWOx
XRvYNvc8qzudlzoNfNRwwUlt41/WKpMKG2tOefJh1Bc0abtPucnTUm7rWeLZQXUM
2kMYIh7XoyF39jhY7VMYUR7KgUUTL0n4b5sA32cK9zvriK8hsiJArKwe7Yzul5Cs
fHxHB/I3LhpiyjIc5efpR64Gdw2cSgC4AY3EymUR/xr3pMxMwmOtFR7IPIy6xvO6
YEzYhqRDzGjne51un8k8nSHQJAoQINWX1FKum2Lnn1h4eV1ricAzEhe2DSZPDWit
Kbe4ajprbm8Af+7ZBN57EwUQwkdS7FKv44n3UWGUwAwVOKVDKabjGxav7qCtralv
LXno7c4VylNXs688ScWPd/gltqfC74//LDPHaz5kJRHUacw33/jEK+LUMx22HIJf
4MRCpdDEpGR+SKu914dFTALkLTNaP662HPMXD6g8U7geSeLkgs1YAcrFOW0VMVhA
U2E/T6jiiL3SiC8XgEVJL6zi2oHYVoPhuVRomW775HSf3y6QoVloELL6HEJ8CaNw
I/OFHDtxVNvux+B+tDtJLHnIU7w98Wyeh2V9pe+tjGiU2m+eCO59GuOvmNr72E7P
R6SUkydpoWyylDmYnoyBPx1FYpkburJY3FmRuxZ4GjbTPYgvhAmp9LkIjSv5SYRo
+j7TLDt/tpsq0Ze9tXAB+s1V3Cx/GLlZNMuiB1fP9bezkbQlc9xI/BuWl/8nFM7Q
psM/t9z2vYqcYM67AiGg4OxbsQIlnHpFas0P8xZXVd4ZCE8x6FRYQcmge8kVkzAm
MzrnZdJHLtcSJdyzH36IjjNg0+iB2kHYNA33Lr8YxU0=
`protect END_PROTECTED
