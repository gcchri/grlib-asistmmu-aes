`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wtjZ/i3W+exPj+JOxLM7kv86o1mqxB/DoD7O2GGkh7zxVESIXu9R5ui0rH+7oNIo
5k1w6xDXW+lv8g1rlKSpgfT8XirGbm+MHOwaIfrS5Jp2mltB5IDqwDJhIVYYu0SO
WhPh7g29+ctBsAuezcNkilIrgCJdRLR1im9ONganFDgV7D3xowx/RL14jZkNlK77
VA/+k0OGyvCQ5As+CBbtn261RJLxJ+pkA3kJNNBqHMEt9xLwG/JcFDaUdMqdaVF5
96VYkANGAe19ZUkjSULgV4l2/Ufua7ODF+csOBLuhfbcSS88AoXChkl7fUp9tcNR
UNnuEGV4i5bZKXBI4LTQMlfcs5EIGrAVgmRYRxEjxZA6gxcSOM9RlB0ub9BoTEmU
nCUI/++Gqb42B0LO8T/1QaCAXTzp71Yhd77EtsnW92MtPSSFvKPuT3d2b6bC/Y9I
K+olELjzh0OgVuxm/py5FPq8LXSg+fsXRDoqwlxdCelohRKmQ3IeEnjlSSTGMXxO
rhmD5VeoR7rq7Bj7KN6ATtOrfMhy2b0sBXo646kAODf2xGFwhKfyRKVe/3vLaMGC
ESTp7SYeuNaHFs3n4jr8+9ubh6ILIeTGcpebzMqnpiC0LF5qpmEHjfRE7NVtnSOg
MeG2J9t3Ukz8vICXDyh98iZTzGx8MIUR7myXMWzPXAVPClNkk8O6hHOk9QzUOFqP
psmshqCuXg0coehI4kmSwZT4vGpXHK74cnf1EN4LpBHQ81MXxqb1Ys95+QFyCNtY
Vhq3SHf/2NC2Ta32L9zpqMO2lzYj2oecXy0szJpEFqMBo/9hL4r3T+AqE4nxXcYD
DI5jbNBvZ5D+bCu2pgPHMdmjtWTKbSeetQ+308zY5Y91Kog4UazNpgjt99b/ipzD
RGbojOhymdxfm8lFrxjJYqkBL5zx5kvCAikwMl4B3SkyNu+Fv/BTF/OhKq7nj3+9
vLR4wU4pXQ2UCYV23RDDbiF6tJwPMLpN4LLZ26rgfxI1gVrrmzPBym6hbtUGcDaR
5hqoV51TQptMfj+rCOyvCjNjtp1g3ErDG15jCHoKQrqLxZGDtk1WGzgzqHl3+m2Z
Ace/lBmD0QMgnD/ZMUIW7+4c8T+5QyBlY9wlyAhP0iJhTd4wjq+CaFGhSjIog38a
CVK2BcQ/OLCl2hasndp/Y7LWidLeuOlbV0HtiWWf6IiNL3RjaGC4brHeawry3OCJ
tKgOI2Ump3x5QnZuc7kB8VE1H2vp+1oxoMKd4jS48W9Idsw/32eIjh4V2x1bgpUR
`protect END_PROTECTED
