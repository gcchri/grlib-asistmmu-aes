`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
op9FiQIaetO5yp37cBaY88w6qvOaQRTcYG8eniK+htQM5UVCwTkSw/0L2bzs2uuw
cPgMADAXBqVibu7OAWHwR16jbg0wnL4Ohak+7eMfZifHFvNjjd1RDeT8I10j/J30
dEwUbD+0Hl/OERA94GewxlTh+h5NETsHiDVCNURL419ZgUxZ2lEYZbYfRu2Ghx1n
5BG+GVG8ZkevCbvMBD5nWDPLjWmGh3M8VSOyvI6IAFTB5RqedjXil10IMHJX/wxD
gWxJggUurSLITe4u/T2z8AhWiur/AVkQ5NfPc1Un2cCVmN6tjX2vBUZFAyB/otVr
3acn1NQ/ybhR6b/zE6ryVuUZqXM7JhItPwUlol5Ov1KB76skB7raUCQefbc3nfE9
38ZBe1mUMmJmlpqrPq/xQw==
`protect END_PROTECTED
