`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2aonyVYEjR6+UFcKLI+7oBQlIOs7HeNYvaABnXx1/VQY7BuSjon9ovvNHhP4uvRj
nn9x9rfA/gJUcAEpTI7BbHPjopJ5Y2lTv5mlbKyKKwqClwMLlp8MCuep3t6QW/A1
UV9U276u8KvRm3eoxZs2UYz7JERq4eIbWVAediI2/xGTrmA0En1apU312AyPajxM
D5AClxzjjP2CvlDNN4VlSaAwBXqVJYEnjDr5XdJ48BJaYCSqPQUO7xq0IPQBdod5
a3zRCsWXj+l3IKvgVxqR2vhW+XhDYVNoLnZDBMcu9gRtyAz6FWVprT/86NecNNQv
EYJcSO1iajyoNX2zy9q02/jCVggQgD6/1wjpPeXyR7+8pnKI5U1RCi3WHLRo0ARJ
/rWGvOoHojA2iiqtibSr7VmsCvmQz732AdkzuzuG2ciW5kPKJaGi0qLJktaqV5DP
ISxhZGjA8ola8TXYrnKbUFj3t+Qq1BO6pn1g7mW57MXpgJNCUCZucYEL6OYeYwC4
hsxjqsyC5M30Er5v9fHROj/X0/OEH+EcR5l08toBhgEyjcs1QyP3xpYyIg3yCO9t
hAA/eaZE2eY5aoM84RkkeLRlTUXSfo52TVHlwkNQHV5KzHGsgmYAf2T8OjPbWXkm
qfT9SQh7lfE1Q/dscgxKh1MnKxuq/IjQSuHIfmD9puullM+JUHk+bfWnIW4QqJ5T
bbWAZKre1e+d5uEcBDkxSUnSXqZjzErtkLAYQgVpErD6bhWAzqh+NUErFWMdPnYk
YNjKLfffAq1gZ6VBrj6FkcjnDl04t6/KvMSeHeai3y2wm4jqqbwrKNmyGFlBIC+G
33byEOKkIBpAzpP7z1CMfVEpjhOa1KlvaR0f0QcnutJG9Kbh1RBfITii/KENBNi4
NXygkc99uBgQkdxa9w/Iw+TEgbMyaigBx+EHnTy8LJib+mP7xgjozd0xvB4ZSEpY
a8k8uNoZXlaT+vyEA3gZjJNU+ciVL2WNu0LBKl0RiDClRaU68ccb/YPdmoERo55v
EJKwU+1o+Lsz7ghQOy+mvj1vs55GQqVqJ+ZWIRKbjADKfuOmPUHTqW974+hKYPE/
xlZMqlfHaXiOBZ8E4RuCwvHOcpwSJR0XuSozmy5pTa9QeJOYAECgOmTnxIe0kQxW
wDfR3zmQfIoiSQnAUuNgjZjW7zLOizV3tYOe0Shs8Lwzja9nX4lSSyQyYAMR1Q4g
9kumAfWrvBwaBDa7f1DTzXezQ+SO4DhHfJBwZ/h7mwOKwj3KAIsJl0zE7dh5z16+
HbnjeU7BP+R8X1macSF8bv/06V3OVBS+mM0t9Qb9tJCtJh65ZT5oL7s9uTgqb0FP
eujlCH4T0fKdpt/Wx5Cb786Qvgu7mqnlE4stAu8XWl6IpupMGTGtINXe+l6Dn5r4
PnjydSYj0SB+4/VFiyjsw+oZwzqc09xqk/iOAfqKPdzXj+2qDfsnKA+UKXZaXpkj
4lZKtnAaQRXRtWUHlKQzftfcGgTaQPnwXeeZOKSjzIRNxqAwDX+kKnUdHETxzcEu
JYyDGg3gs3CVhF/kfBtAZ2r4RzzVLtYu+CjVDNYbkvQds5EvEWIO5Tp0rgsRPMKw
ys2c/i01ZzXddIOGJ8/s/MjS7aGDcixNIGawBLg3b3Ene1mGFy0i7d9thv+fvSjz
zVoJPzPQ6+BO2batT5EifyKhzLLoaSgxao3BTFeR/W73gZwE27WVRqQ0TTFuX/JB
jf/oa6idnnCGdiaa1PzZ5Aug7gjERO9sER9rV9oCND6Q0I/Kn0m2U7UXhvIm0pwx
29OYWL/Ej9D+M3cROQtcMvr1pqFnjxcoP/WGsPzpQU7lry8Yj2SkdBHiAGTjCDNF
gvjdQgbtDHr7Y4B31VHL5Clnj7DJHf3l3fJ+cRtatweeOG/VfIX5avIjqtaOcK1m
2TbXuumV/wY3L7GssaIfhMQUUOy5wHH49EVwP/ELjLrtFaC0nR426D1mTarY88N1
bgJkIkDFicQ3WsTJI2+xYxwe4KahcbniGa8S2Jx/vSl1v8lfOqOL9NdQumCAL1lw
V4ImC1/Dh0v6qHUs0nzx16kYs85WWdUZaLSYkpi8f4nAXR/aDTSviHnVYIwx2d9t
I2kQPM0ElKsrBtF8fFev7VTQJPtnn+XIbui3wZwvP1U=
`protect END_PROTECTED
