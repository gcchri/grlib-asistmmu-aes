`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y5CryNkpG4UOXwJ7WIu5CHXxLGQTT8Fv8kGds4BVAmkevS8Xvy1TIdRpmhq8UdMa
dfkWsBl91kcoq5zUYVNlrZnLGxoJ9DVDYazPwGaRwfaIaCWkrDNa46cjBAF4BV7k
sMIsyCE3v0tzfub36Nn8p+HXe3spI36ovV2rYjilpRhZJJ3Va/2nSWvL/u1Awap+
hD9L9FWUFGydG/xnL6bkzVLtKVwBono2yasNyaHFXULU1dYbyaQebFPfaLB1i8Zp
xp8bkS8IzlJtjCxYYofNmZmckszWQP8xe96RiWy7dSc4T5x0ttlTsSLpEWUHbjw6
fCNzuebZPZvsxmicovmtj4BGaC8N3IjjDtfBAXo6PIgmWloodNktd2rH6WFNeCl6
kLVY/2XnfLebbhXZfH9hkGL1dXNkyZ4gOOscWt0vCwlQt0FyAFTZwRHaxw7noU2Y
`protect END_PROTECTED
