`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iLrIeMM57l63jzSQVf+lVJ8ggjVN1foGGrExdFYs+8fEeSi5PXwzJBM5inJ8QHUQ
raR6OHCMxtf6NJFZvAJFP9Uc4bWlfA56IIXev3hytpHN5qE7oiLfQfeBOpytse2+
uz1e2vkXIrW8pOyD/fpBF66goQvJsozNaqREhr5n5bHyfdneB2pj9FfX8ibPJEg8
KiDwMWHCk246ypcapfHWcIW9NgOFYHr+IK0E3K093rk5HSubOTSAvvSdG3m9LkVD
GIJtEJKkCLbYFyXWGQG9LcjMdibMHo284FsErJF4hpNDL19JCX9S3ONH3AUu+fxa
fAeC0FmiXDWs2jnRGWoQGdLDsN9K32ZEBQELaFrEsYi2yduECcClunL9Uy+U6J91
RZV7Exhm1gZMo/uSKMolqgwmlDma8T1AbG2ldAv6tpqsky7+ryt9PT4A+G3dyYOJ
2kEElP7vE4sbgvdzUzvoig2ZkjP3Mbvcrdw96U/7hiGMNj/JNU4se4bKpkt+N+ie
8q/CFrQj70zLBIt4R0nMg6jk8a1TGJ8nkLeTl++YLqFBsDiQxSlE85pn5FGFaF9e
a0GoH9RGvyn5w4sR/MMCCY+vxBX8fLJI2IfbUAba8DOnJR1d50a0ynfOIftEmq4O
CLJ2GgEH/UEOlpOv58jSoB0Jea5DsMbYE4LysMC+3QGg2t8HQ6jB66emskPEwGwy
PkN22vd+vrcjG7I1nSqKkWzPQDf9Ein1Z2bUNc2MqYLSfkDQ5s8Wj21BhuvbU/mQ
GSsU0iUwXu/jjVSVAgeMnK0fcJOM7r8kT+BhDCqtTSU8nX6+4Fytqn0Yheteoztu
eFanpkKFWKffBLJcBbyjSc9T7vvsl2VtkrPB3ZlOv6K21pHDXtiQkpqPsIG159SI
qO/A2h0oj2JR8HUi2xUTZ4MVncBpmaFPR1KyAQLyfUUvwXIoP5NKyYjnwRF8KnvQ
iEJ/ROqbLKuQVDt4wYJxw7jOqSnDoKGS43XTBThpCP+1Db8kQXSjOksMjeyhNIIZ
ONXrMWvUnFyV8iIgoLpRx7QYrHWTa2uwOstyIE4pqhMQeOK57PQw/pFpA7onxnkG
J0F827gfjPr6b58fZluHiTsVCpHBVCvDzhfNOI5EtSuPTa0usUF0sOCdCcl1qiQO
0dwpP76hNmj2EcaZfvg2TTwU+I3gPlxGejV+HHknqbs1FUmOkb4FsHQe15uEDVgB
WeBDTM/CUzP6oA53un+/GAyvWJVAgnPhx1jJsVe+6+vAOrhawZzC/I3uZD7pnIwi
1A3UCkVJfxIxDySQcA6xSGEintEUk4bYQOsxX/j6nbFIO+FcHBdWKiQx5OXEx1oC
vnzUtYKeDv3D1ng8OijZQj232v1EF1U/RuL+XxqV9lubnhWOef5mvyfwIxQgEWfP
L35zZ4jl+9n5ojj4bAYdir8H54daSQWYXPlgs8ZsFPfXbtZvVGJJj1wKOTsrtMww
vwNTRrLewjNsqtv51YKNrqqYupdMrfWhqLHff/8LkFt2bjiHR99dTh8wXW5itsZZ
7UETYqEleOHBJx1z9LBtutbjImtN2Jvr6Flpzn5BVHQ4gaJ9FuYt7hU00Yr/nWfn
9bMK7xDI/Eb8Vjk88NPr+uLuKy/fR1Hwqfzlozz8X0/4sL7QvOevvQrEzPPW20Ou
2h+t0iYOd0mrotoadpykAtRqgpWVHBY/ZmzIlnul9fi6kpPFb67/B+6c+VO4vmMb
FopfjZg7I3rkdKsrskJlx2mvLo+QALpl0+VBj9WGsp98NLfnxppaGzye7nz0xDvz
vBkqN/+V+y+mtqWxnJyQORPf2HvxF0KLdgexgflKZ7X34c2FiMxbXAr7TPCwjIx0
WS1eVNPfTqU7SD97IOx/Yc6qHLPPbfw1HRnQCCXzUKMi78pP2L1z+qyOGkgJM3Of
1QF/ig4gYDh3kQakXD3w9qfvWtqz+8liqZBcNfBmC3z3LKEeXhvJ1+1+Ia6hyFF5
ZHdOZFMhKmJpP23zR+iG8jAIjKUH78GVyjhJ3+XFmqp7w+JJRxN3mP/00GktMC5g
uNg5ThsX9bbhw8b/y/MT0lp2et79HdItrLKSv20P2ulKx0O/Y41FcVYFks6uM+t2
fDtxrgottknKLYDofBEMvKjlEIutSikZAIUlpZP3JNX7hI0FL7veehVIlafrwUNC
58Usy71yTP17vo20cmdrbCc+Jj4wyauGUUUTB/EeZyR7fojrMV3/unavwyKG9tZn
0zYyc3GfCIFHNCjvLn/YuafaoNZU5NbVW2MgZfgbF8OWNm+0xJhQ6zP39XZ7p9Fp
SIHb+DtEsBmEd15kWoJYxnM8rTqlsGNHWrcVB83U+VDmcJ9Dq39RlXmFfhzyThU7
yPCEjHOTjRWrpYlD/7AmqKTgCyBeMdzHQm4q5JQedYVoB86C53w+tQ8OglznFABb
bihyY7Gp5NoK12cWFaHJh949rzZogT6aenVzXYzgajJFHduROPDur9c9bpEb96RX
by7N28Zxi58igmv0FjxV4JhRV8U8CbRJpXtWdtH9Wb0IO0nNgYpwZj4ZNtLfMgdq
rv3ZVo+EDXI46CoSOuXzzT8yGLJXDtOVKsNZBOeaUJqrRvaoGJnPX/G9cEO4pk3q
gx/xU12Q9WrCFLVo7qlHoXJ4LuSB3VhnGo3AfZqOKteeDcRakGrnQQPfx36YU5Kq
r80+18TjEdLi8EoBlMz1LvYad1wuaB+Did7r1XpYudYLJ0jM/VZbdYMaZKKpt6VA
FCy3Uc7qP0X1HcT3sPfSz1lVAPlATX5bubkJ3SXqf6WovqJtu93aElQsV+T89WVZ
5G+TH317zJ9NeMke4Ushpxc0wxC8eJlXO8NrMzjdT089GgjDDRa6d4e+Cg6yXAPL
clUBxg8A3BY7VA2aGOjeZAPSvwwRkGLgRHK3ane9u0BWsJXc26KXAjNsnc7Fgq+k
aIbD8kRCZQw8mMEgLNtYhn+HCQW8knP2HnMQi9UDTme/H84IG5Da+RCFFrD+/40D
elw2Xbl7dhIe0ROiaKQRl6z0HOop04D3RZ9nReN3pJ+G6dfRtRyAJrhjJA843hXh
wncM6LA/MJydZxPfp12a5T+PU4l5ptj9NPf0W2k4aCQkDPFXiQgHEH32AYkvc9xk
qROlw9dqn05mo1f602gc+vHyx07SfTfzWGR+NYNPHMd9vVmQj0vkVnJLkgrL9jFx
X9vIhFTTR/7RSy5PGtKvvzf0acPPd3Hhs/NufHl8nU6aObzT1BhYpWeKOyL0TvK8
b0eZ9bkzFOsD2WNG2FD8Qd5wIZzL1l9o1VthnZ0v7z4nYrhE3bESOvB5fbCkYScQ
f/HLRC0Ar4hvS1CgICGBSA72xlGVk57dj35tEvbMQJ9cb9MVaRkKoQNhttt4F1v/
EejhGAkvHdR94E3HYOMvrlqsiFid8DxOPV9GVcH44Gvurd8dQ+/srmPZSAnez7fp
hpWWP/3if4j4H2BYoMfO8eREk1IRwyEucvyZj7mA6HQ8JR4f0/m4y3uRlNPxv4LG
C+iLmGrh94jfxFUqoTwut8rwltX8ISAqg8jGRP15UNlPYM9ZEL4zXXCtgh5tOe9W
SEwvBRzvbFlP7lO35KNjUu7Na+RPRNlBMnTQsYut7krgMcceDD+2kf6NRJM1unb9
AJ9Vrkz9fddG2vWk8zTNSGSXL02M+X+2Jgl1PK/5TKi7VM7RnQVm5rJb8i1L5vjZ
ULJgjGuuMpfcgpDqqa47/CI45zkT9t3aAlJkcnNtPro4w1Wszgxg35IrVlJzRC6b
2HmKyOZohMOy3skmNIWdbBf8lxengtCYZYr2MnbuQrP9ejzmaeGbTg46TenzZIF5
W+J2I3gQKAogDiT2KJGBEdIFpf8VkHlkDS74l3msZyBqm+SHckw92iKc8oaRGzKX
Pa6QgZMaGcF1FO7huZVszGJXvq7TM3+DmONusgDcRHOz1IMYIrlVgN/fTGkKlN9w
zg5m0czq+PhEt9nparElGOm7BBF8RyURKQBJpsdPUePSu9VxxcDSueL4+Mp/QO18
1wEGfkP+r0+Ye+ZcdENQFkdSBgK8H2MONxegBvy4nwsEf8iQLS6bx0eQ2oMnBn2q
Q3z+YzOa2cgAf7bbTk33MWGza2aFpaYRFcM1gEhkOByjCQ7WHUju6iOufMODLmZE
GQOMXc+hIHWcgZ+/sU5gGqZJ8rxwQ5kue+2pQWdEtJT5S6D/T1d4Ib01UPktPQwM
cbTh1JgmC2n6JleXSFn83EfYghFfFER8RPljR14q5nb6Q/IdSXdfvd00+HlizC1V
2pSIPiiyozFFGdznDP+7uXCB2PIS3lYPQ+Lx4Ny1z6DlPP21kvjWVPJLv6WWpgJm
6Ap+YAHgO4a5GIAXnxoYuh20BqXE06lXu9vwNkW/o3KcdGBFAJ4fwIF5mR9C17Ew
koaVQeCh4074D+ZKzMe81v+DRcQsnDMikPpPTOp2fJATdhAVtJfS0zfWUpIc3gsL
UWTiNjhCVyNSUpRfWm0oLwmCgpP+5figfD7TS7NpSi2sN8Kzy2NhSuoKF+MqtmR9
2hO3mJ6TlaWC+befzK0YLvj3KbVb0NwaqygbWsOuq5JgVJu1q3xrWrLXg6O7E7J2
q51bP9nGJg2GUQ+tNxkdc34ZIWL6NzGdX96i5E251y0=
`protect END_PROTECTED
