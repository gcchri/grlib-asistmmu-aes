`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dC3YAFMpovHWmusCsMEA/sKXcOyjYKlzI9SofKQMvtbvQMQBc4t8FYUdAQ58FrCs
eHJY96SDZtu7AuIpnQDxRxgGU9n79qirKhbRSvMDwCLW8JifnieBNj04UfJnNxaM
NmNLZg4kqzCpKL4cP22S6wjtEyoYNgb0FSGOoQ52xnkzMCnJWAsEdV/5M7XuSUWO
TzE6Gce/mfNGQbCR81uGYTKTwqqwMK8DXqft6WskRvV8moqx6gFscSgr1x5H/gGc
jA3ot4rsTCPzjTyZWuIbfXWi+GJy5+OKaxn9mnZKLHC5Vxi5mPKaLwpdUTLfQfXB
wXPYU9HDlth30OOtumOG/qeFu/sKFvXPxZjQM1U9sBXEO6iCYQE+mupMqTzz7d+V
0pjOfE3PtR8oJpajgVNqtBzz82c+T6wuAUBcjarkgUebsN9phr0sGnXVzsQLK6zc
bhvnkDYGjFOZck9q1es0bExc7/9MXJ5DUHOOw1dOaKJ6lDPIc3quxtICwjeaPWyh
zKho+FPVNFp/TtMQjyczHZM7FcmT71hWWf7mCMU7eJ7zJan4g0GTdaXJkdvOfMTs
yktLBQqXb4XzKBw5ak7s5Ulu07FdCdpQ+t5Dj7uY+99xkgmF99nzDQ8wKP4u/L4m
WCu5bAF02ZK2bD70tUmBxz0ngLiXG+cCvsJnn7+tAKAARjPcJGEnSCVVOgBpMsQm
uNqIaihXRP8W341di5maGnDQr8q8SnbIFOZkJ29dZUYJdHN8f9hlJ1F8wSWB4Yuc
pOamPXDXr8bGTFMVf7fkKMNXKK79YmFbqSo4HEm2xoY1XZIuIENn239tchiAl4qz
P68FrRYv44Vy2GN4XjtUEU5dO8WkrbVSAMsNF1JPSt6Nf70ai3ffcK8ueYQbCR/U
oRwv9k72TJtqtcma7cl/8JHqnmmG9WA64+/FwMOqNBsXWvpvYd7Dah56ouw+n3xG
smoJAwlTFYLJp8fpZr52duIHsdbQ86Se/G18bf9PAxExtzn5KWHKK+FpiNwvRwxo
YfhR3y0epSUdgBS0ri2hIkqVqTohQ1kUkONGb193/PwV4m6dAlHMkwFy7LUx9Uqj
FFTtMVU/xZ7MtmGRQswok9ltWFp5IQabhQNOZYKrGcucV+/tE8V1GFbtqxphT+Yb
mY/PsVI54p66bxatfVCBFnQUSrRgduIF3k9BGgmPPVHosNIeefYHI2yUmHFqUnf1
zm6HUjhZ6D1GFQnPLy6QOC0EA3jA2rentsF8QTpxu7IcqC83qGKl9UHZjsiqV3Z1
PjkSW/B4rkWuw3MJZMb76PkqlTau7zw9A6VU3Vc/jK9HftTBF79o+Vz+m9EBZJss
562X35qoW/PhMRocLekRmX/kV1RtBPksKCYU4gPSP4v8N/neqdDLIN5sQQmKyGvi
XGVVrsplRr51Co9/hjJRIgr0ppNF8E0Q/AVBzRRc3xc7rmS/6HFPRDPt9HGSo9ro
1T5Qu298gBLLhg52iHVEdqIaIFxYXv0U+3y/Q4DP/HcV9ZXb322S3uCpnt+CDJt9
Ty7VavF+bANeChQdh6MKvABPNpvfFYlWHNuJO637nVnHbWWp3bYvcQfPoWX78YvU
RGpLgNYlJV2TBCsmjQmIq0tCkybEjZh+S2W8oO4PprRahYDkpfAs2y6nQAAcuHkk
gdKYGVlyWlrLUVE3yZpdvd5xCNYnpli1IRqrii8MuOvJPHXfRjFaHAwf9HlaLQ03
VGVJx0yWNY0jpeeHehTJrFQwqvK/xCPzNdMtbz+h0kJVRUh6XoSFvnMZVb6+piMd
bh3a8VVNDfSAjxRDj6SLd81Xzd3EHpY0wr5FJj+3hY7iH/nhhRRV9/O3wfMbtwLb
HHjHTrfoOvsM7PNMeGnGxyKbsjDf8kln5acU3oaLKfaxP1Cga7Q7kx2svyF6MNnT
AuC8QxiOSsc6XhQnxnjPXmF3i9kx+PT+yDm8/Erd5+6ptq3W3IwS6PXhV1eq+gRO
qK0026vYacpju7Y5oYlguBx9KrB+q2+0psOGDKy0JI8Cjkb0z/eFsBlbhunSVEhW
83etMpHYxJqRL9xcwtFIAZmK+PjuRhlPoQbFFV6swRcBw3oYkhGTiM6Fv3JL2ULu
+zunXgy9UvXuszXnzNovY/c8FzH04I0OXINxetPk7CIP5DT06586euj3YmSP5GTO
vaoi4b95Z7VxdhjJFC0P6wjpT4aMxI/5MSOtyTyhKxh5uOD7UdFD09tS6s0L+3uf
9jHMqblDyr2PNxs/RY3x9uMy6yD/c3/AGpXL8DfsF5lFrlM/KUEClbZUSxryEgeW
mDwQAUuT45qbwYG6YvHGDieHN7oKagdTWMfpvOVU7SAtjFwsPvM82MhGNFQC19/w
+hGWwgYUIPhpd8ZWd23MsMKvjcTEfUjrgWZ9pLIBfkCOzFTyC9MvRY+PoLyiJRoJ
wJSFU3nq3ehVfZMfi6IlpNrcn/973SV6iMDIEP2L2aEAW8Qbwd6YwOEzfjGo3xHe
3CRy0wWIVe/BgJfHCzs9IOz7aLybMbV3aREb2nTYmDKKtFXJALr6JsEGbiUAHKEO
cjdxm3lzwQbXafT9kzJ6oQWnmRdS0+RjdE2eWbIYKJXco/xScemHQ2RbMOFv5cK+
gKYTrqIOseV2/WE4pslCw819Wlm5UZ6FJiGWD3sLIYm8Jm6OVtnl+Szji8MML614
2jBFeyPByzGB7Ak4cpQnxZiCBUzRS/zqiU25nBfkpoGSomwRJ+0zE8zQmfqxk+21
SdDYRKta1sw8/lZjBTikr6uxd2/2YPXaynW8j1MbS36KL7HTbiEh9piY3QfHtDef
YIvUmgK5/oSXecPcrDrEp7eG+y0ebz+fytnB9yTU9ZHQDih4+X1CtHn5GS36rbjG
BU34kcAsyM24IanL8GkrFX5MS1YiZK7OjT2hlqctTph4bYWxZ5pA3/sMXgXzm+sh
NfUKMyOAcK19nVG6bdb6y2SIRiNTDr8jNzC0KjSiQxssXzxNfBmLvGce89YwCw4F
GI22j+KOXS0KyTkoMc1wLaEkxPZJ/QNLoHbQkxDbqX6kdgMoCUWo+i151mLv7zco
pfBgk/LcpS2pEEJ+UItIlmUAO0TABJQahWz/xiOi5EncX/s3gm0+CkcTEEOMCCI6
EyFdhWTBUanMbtqD/aCfOOZUjph7RnUNOs//BcT5+egcvIAlIexrMz2eRfQtjZzf
MdltzUhADWIwE72kJehBQX8KZORIqT+ZEXGbM7zFDtr2JlzqgoMLd2wxECMVTO7S
SP9i5vKHjpxoRlQsJXOZuxm5btk4/vsCJxfGUBCDgCHPOl/BOVtDDgFJ57rRdgKe
HhOtTJEIjZ7aKzhWy8mJSsDRauys7sstRhVPDZ2V/t4fQ9jF0XzTd+5sCsS6VSwU
Uso4kh0ZJhtRNh2gFBeLEo/T2voWRkNw6lr+3rZQgCdIkZzSBm/TF2Rf+HFu7lDp
RaUWuISt+QplCpHnAs447bxs/ZBhWKbJBnA2y38lsrQF3Kn2bs5s4gxWsV+veoNT
bmfGv4EWmsLH0exMtclvsCYRAUo/IYtBRHKhqN70Xp9z7hY4VJ4LeL/0n5JbsATX
JaWn4ZrMfUe09FxoBHL+aFcBenDRJ37CHsVe5x/CGZVcOw4B16bKHt4SfH1ihN5K
YA/aOhQ2IcSJda/20bJdVYJyfiRZZzhkkZlybjnWGKPyVGVNroOp0pvZjXjpo97Q
IwiEP3n89Gc2Z/kekKTCHs3sPSQM0GWm37lXyLaDCwrrIE1UEpwZLEfOS9/k00Gn
8aCpQE84319aSR6V5HyLh0YiD2cSP3uEOLttQ+Kwx/l3xElCqPQKn2d+C/nQTaUq
Bp5aws1QeERoazR0s9el/OaTJ0SBx8g6t6SVqFrneVHf/X56ZFKdp3nbw7X8RL5d
dlAhDLqhhFMjaeCI/9xTwg==
`protect END_PROTECTED
