`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oSrucR7kvfQVy7B60YB1pER29z8DHGPkfI5dD1OXHxxq11mPoeyEtK2FVj7Q1VjU
kA+5FzAp6dFWrAbX1+LJn4V3ku0j0k9hez1jwYRCxczgBYp8acwBwKKWi9Yr0+kL
59oYC6cjnbwbs2+p1R1TH1QgDrvRluiSx7tZff4HSDFkX2kR2fU9sO2g2DeWFv4F
lC9VM23K3UehTbOA85EKi8PmBd7OfQLOVFnqL3jLZiSihpN6g7CC+qlLigGx3JQS
Pve8RlXVEh4FF04oXvhGLdio8ceeu6ZidOq2hIoIKwiucnBFGSy2sVRTZaPt5PnH
0RtV4kjvLCI67C9FarU10O8YwPGdel68PGKmfn8yI/qj5v6Vc30LlP2EHGPdIsqI
Qw5Ul1fow+Nf99BXpIpwklh+ZJrZJ/OjWgH1x0d8liTuCjzUVAI8wqO7doixLwwz
P/SUsl59noTgwHIiyglL52QgxXzkA9OwcN1/3PusyGj/olIxVvXtpQwwcNkxGqEx
wNxsHRGkW8+IVNPfzN4VQfd+GVyoyG22crYMbmoSByJuUws2OjAkz4sDBpU0tpmO
Git3jfTgqBDp69U0/arMhTXcMvsf67e/56NKEv/p5R/tJeQ7Qd2GYo0iZVGdU1wC
+4Uxk9BZm+4eMQvVfgIfNA==
`protect END_PROTECTED
