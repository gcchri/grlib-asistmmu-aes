`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l8k91oBKqkq2BsvMd/iW5zw+2Q18BOy2V07C589YsDsISeX1OB5cZojhqhEk+5K8
iNtsfuH6Lw+yBmEWK6eGQmjGNzLk4RVELcdbQWNLxnwOccNdTdxlC4t1usrvnfX2
NhzalosEt4BzUp/0Wsz+suoKqYjEM6RpA/cJaGxNSFvcNp1IUnWfNMh0MPbqI8t4
m0sdx60r48LPcf3FTlkpErp6lpmKQnb5nnbYGthpSvDiGz+UwdbdNV7ldGsqVZzI
wzcszuv79aOgTZg+0oQUlUQtGjfoLVpMvP+CHNwEXMDUL5jEiyX6b8M3vW/2wijU
DQcPd8Ws7jvzJbzsRUX0oNFP6snAsevPkvWdV018UOk=
`protect END_PROTECTED
