`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
irccvOCr8FQEM7RwwbYFijcCwMDo7qP3u3UkOkuDRcOu/WTZvG+5pOHKIItKUc+z
afw5d3GvUp/+HCWAbXTYGMEpZeTHlHJVMb+b1Ov3WNXsCogYUs5zF6x8+XyHEx49
TnOEHXSuUJcQkYfJRnzIGAgOsgg+r1+PHZpG9qySBLY7EOhvgiQ9fvXhQNBONyvO
gPw7zn7maFyWlfChltLoqX6p8EzIVRLgRfhwudWomB7ro9jHaBKaV/cdg8QJrCML
PrLg0sfZWyL9K8Wb7ffjshXke1WxE8AZZh19Z7i9mgJlv4t31oPtYSR4DeEr2YtV
jLIQwiW16DLnDbtOxPHebeaEoXAjHRPSnW2i6zl+g2vXLXq6nJsx33qPcDe2LYqc
`protect END_PROTECTED
