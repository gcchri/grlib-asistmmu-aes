`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ywgVoobHY6h4UQ9hky9E4nsAwtCC0bnLXiD4yg4ZcnTZOW4kzlGNT57cadtah9h/
NHGhNrrGy5sIQHmvnve2Atrm5tbUr8fw+uO60AWZSYHskXgTiowdyCiV+EHwnPrY
w/OnLAWYYkV1hI3xLbF/bwxvpsTqV0oz8C2XGuwnQ7YWSowN9Mp9NIoh59NGTswF
kdiVTwzN/QRhqaMyw8fMGPiLGWYaO1z85H0sMwGrV2uIvLg2lvK6svgIxnyo1JeT
Zek6nILQpgotMT7OEoOCUtYjxagxX0NABf1q5/pr21bR1fE6SDkOZZBE69VInYQ8
P9cwnykp5rI2oco7GugApVSOH2SUuWd1BySIK6aO/DzhHCOmOktBWjbVOsDPgVNv
eHXbBfUMng6zfks/xs8uyyXmdn6Bnekl/1GlMwldvGXf/GqFqovl+RCNfO0wKOYx
7eA/G6loWTK0b4hF0Vp+swWiqv8WjD/dYEyDKmG8Za0XvzxMCz9XNhieWWgyVwB4
VHqFWeNa+d9822sh/6PdZncMMdBrdKrb1SCCxurZpMA/y3bbeVX2/twdQ5pbdLlg
2O2L1nsdEyPz5gc8h+3chaGbLQ/0xPax4LN9SGL6WbHYhVoVNL9FKDcbgX4itgBK
/H8aiELMkvNCiVTCxFsRagkquQ5XUMlArKeT4KRJamha8Y9B956GXKZksB/bsodz
tKpYwa5NHnYY65xVSxoC5+QiYB7rSuhpOW9PfM2e77YTtqJ/B8OcAVa+D3ckBscn
wZM7vC6SxeSN1+KDQLbTot2vQY6A5SL853ugXkUTI6jm5q4CGmDU63Bw81iOaQRW
MLlrXolHKFqpKi3egsY93kipMLF/ox1IHOgljJ525/4+REoidI6qX2cGMf6UMBao
i+U2tokhH9cu8DwCeETEl3JIfhbKZEeKvUxzh1NISPvslA9Zs8VMSIh76S9i+f6I
XlS7hRPy6V3Au7EoG+Wk/aDudPBOK5KOgr2zrLdbN80quYScaxMhX9rIbNN8uC0/
TPSBUt+dyT6m6PIoawQJXVRC+JWaHtS6x8E/G5mrx61XBvdUJUOjQxNQxxbi0zCM
hNcacdOPbDS6+6rsGsQg3+ZYmyXc4k54G64wLXVwSxEeIonsNk9Emn8AOrd7BfMu
vtGOEKobsKT1d2eSFjuVwu5Kmw+3zL7kWjSav00gK0RZJ9vcBK/n9+RHAPyGz+vI
QODCGj9GUov3B8O6Hd3ZNJbWuv4+Js8nwlqyNxSSWfIsbe3ECqS43shOEDibLTtG
HktA2JyQxGNBmt+5ggFwgICl6QUApbj6W39yt1QYtRyC9gMMFERWK+oCqfDSOxh+
bJC7E0+Qq/g8N4ij6FEe0ikwYWuXwkRrC209ff/1GmCXFeYABp7H/PVDOzVTjIpd
v2deT3pibYjIqZpR86luiLMtHVyx3DlxoNC9ytW0JNt1YQwKuVBCf3A9W4vzN3f7
XjN1ySbzMsPC70ujSaO1/URlIRaEcY/S5bG4slxIzDY3w7QRlj5Rtq9BoFfQMN0g
IxOxzsDjsOYpSwwv7nQxslkNi5qJG+k1WLoJk7DYSoQrbehdb5LviFyJKl2mQ6UQ
2NGkGzTD7gACMW3836py3CH7rahipfe3nTJc1ukrgDK3iE9EOrA436v1bTY14pii
IUJNiLqDNhnY+SO54Sa8pk45u7JsEQyPOR28ggBNKfA8WxrhsuQ2O6jS/ITtpCFs
wtXWj0tfWxW8aBDZ5fVHkgbAHA+1CWEQqVSbrkjxA1HQkrFh7k3szurfc0uulcqr
jhH2JEmWYnbB1ptpzWDZu8uP1T5ttq/Z5VHBFexoMP7r+2VE8R5GG7r6dx7HsS+U
V8+nWSBZTKm91Jv81fD3PxZ62ku1zwtV6adFiiLrxtO7PjqGsbpJXtjmHEm/kzBT
3qkGmGc+t7QT5Pd5xqAh0Pnfn0jEVxa8k/2/Q4/iyPfMEaoM5/Xa6KcdJjZlb7iC
R2gWOxO3wHDQQodT7vjQhbyMQ15HiA4VpnXFjRod7uq3Hl5rXKdJ/SKeTrG094hd
2ISRp2ZgD5x9oaKiQiXWQuWxoo57IO0spS2kGlvQZ4EeDD9WiTRztDC0jz1a7Z6R
w/jQSKcZphwYldHsOf0l1FAG7H0wO9Khq3AEHlkyEEYwlpiuO395OFpiB36dOu6V
YShCCXgAqb8Xsa2PWbLYe7l6WI5jybUD7Bw7FHnEw7WJghcRV3JZSmR7ytCo0JdI
Wdwyng8jv866fbXSXzSOU8xLriPISXcfTz68fpthDLcLfWWr4F7FMMb4j/vqQe+I
j6WxrNhTmJVL6UCh6rjKwV/BXcspg4wgjOQRqTcK2CV/Zox0vrEW2s6cef29Wv6g
/3fFfgaRGTUzTVbKnBJcrDZu3Nu9HLxvaPuEOYTdoqs2Y7ZO0TeAY2mKKdrbQSI1
dg6K+EhATHyjb7d/V4BIW/yTVmUd5e+8J1GcHMz/WNjhPlx+Cj6oeNhElfGUVFuT
9oHLBMxUm98JtAvhsj8qOBicp5XuYBYO9ugj+EWOWIHbOKiS3/nk176qMWG7fTsx
QEvuP8hb19TscRJRFVkmPLejeXaIm6KAdu3SzPCOnSi1Q+DDI2h7MgAtGA06Yo4G
rfzvJiPY4F7SkM/c9EvI3RH5u0a9bAqT2Phoi3sEntZARZdqWJs7N2XnSUK6F/Qb
G6mAWbyCT/1FLqyqGNQgHpgoxJNgxWwJvIrpQt6/Tl8T/ZFXvpaJB/RRl6RWML6F
Hg/ZFWdajBmQeEGQ6ys9lumbWkTFiPZj15OTxGiwzDrjI0/O2FTZD162DCBx26py
to1wpBTgln1buLrqeKZ/B/P6OiIdygYpfTNDZz6UTqT5rbWUlAV/k6qsUiCbfhwd
c+mk0V8yllsUSdDkdb77n0RGxaXnK8mi/tjF/MQevYrJkVqJQZWpDD/ULPRUNPeg
QG5V+53qYkz/jmvYmlvHHH6UFU5uu9FX5DTpLTH2KPdkslRLtrsLrCrOa8mNR5D8
+yfXh6F10Z/xV6jZiweqLmePDFbeqdQeY4AIx0iwyMlzNz3fvP6TwrsKo0pc6LJJ
EzaB6bYsj3jAKXwRY89hX8QaKVjMte7LeFlKkPN3Je56IxHxqLlx64v76KfwK28m
VJRRHziVD4Qhm6qK/hdt18hgGmU145Q2ni9YT01l19iIV2kKOHteAwdPkEThA3O5
rxfmdGaaUmMLXj3JwMXRS9SUph55IetgFFZGzg/PqJlubHrVbmGUtoe2EwYA7/QK
cU3SHuKWdix9pyV7M+yUJe3JT6PUl8Bx6kPEg14s8/7PUrfsV7tb2hsqhmx0jkb1
Wt/kTi5d+qEaPrDIxE5sNtEFrFiYsmStRh3GX4Ut6jWkyIb/Y+MXpHanrnrnPb7K
2OkorDk2Buw2ec57NfmFGuEr3GJ0OvAxRjtACnxh/gNy6PVNgl1i6nqLDAApvUUx
EP1ZzmBckuHw7cWo2Y1ouNoY3ODR2MTV3cURMEmFXxqVVCqBU9AuTcMsoPlsaqAR
cHgI8rw/vzsfdDrMnN4f0DPfAx6BHkZXYOMAUWF3NrpwnXdZp16H+hRkGF5elypl
QHW0njWEwROXl1UJOAOckyuNfiDEHRwQD9TVeaJPpOlGv+/a+OX8su2C43f/mGSq
0TDEyu4VkXJ2dKG4VbouLuiVV1nsRYd3Vlap6LYQUQNkalG7nQRO7xgWQhwvVSTU
Dniqgsjj1CxxxCQOT5G4ecZr5LbX7X+dlumQNT/MEcS5Y7D/IQgY4fFnPiP8w8fG
kIp225oKezCRkzbO5D94s19D719pa/75IDW1z0Yiikp8LrkYnO5gRACg7zqZqt2Q
dVSK/VloQIvs1ULi5de5tJl/MRGw5Mqy4SSk2OR9pezsYsDVZAqugI+foAKfh18Q
cxiCZX/N3/X2gha1yww197Y/mh8BzEfRBIOYOma1kJ1rDqX1iTodat8YBbQegWUn
mVRRR+7bZyYpHL74RENLbIMZyrpuj6SpZ27zIHBSm5GPPVGMkB6jxMRGK31Wawdo
2T6l+srNmwlS+tgvvPvNY45f6RIf8s6UekCvnFBOkte3vT6AZqWcaAzha7u8jwfF
Yhj0Lkz1pSjlzHlYpx8PwuElZLEORF0cXNLbZ9fZyJ6bNgA7pstXkYGGgaT1IZnn
dnrK710cVxV1MHoYhi1g8pFJ2O/IfOt4nGZALhLSWFxY3OqR2Kdo2Th05uWD41+A
Ce5mi7TrOenzPdtPhrmUZErsYDgmR02XSQbML3c59zXGs5xU44STNA5+mQ9YqLyP
MKZj+CVVHtNbm+1ysl8KqqKPIScMaIkmqyRW5gr3Or4Jf3ljrYVYSEF+b4HbcFg5
x+NMt0p65NSz+cXFETkj5+6dq8vD+fs69Pkh9CSMuCPAj3KKdbx3xSnIXhX7v9Si
KYZ8QKHguPsSGfqH3mU33g==
`protect END_PROTECTED
