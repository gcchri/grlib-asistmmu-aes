`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G5BrevvwKu0iFGecn61ycFkFQaBnM/ocC41FGX7rDNSLUi2K6gJOxS6A/J5xC9O+
uQVC6jLpEkkV8m1l1RXn0IVZZbFUnuL6pstJP7NICOELV+TOxwXGmcDM3rLeUYY5
6BVm14920N7ebql3mUgaukjabBJ4xXL0GbJFuM26vpnpCc5LXFFF/27hyMlBXBoB
0+6PKOaJcbdFkn4Kj8aIyfkKUy6TFBtXAm6pOJx8gx7l66L7tUo8G70RvNwAoH3e
obmBRZQxJAw9YLlwPplI08Jqs1f7BusNA633bG8w13FTXMGdjzwfUS1JOG8r/IFk
U7/scSDKlB0PnWAL+Todr5tcFjzqJZ0is3czAcWg9Ose3Qjvl3OF4WHOnxf2HbXR
ohhBWkxanA9OVqwn//HO5K3zGvOiwlRH+bo82RzLxwmyV4g3v1iyfk5tpbfsA4H9
IzHS5EGizLxwoWnqN3CPLmVirpWm9R9HKkvEKCtHopU=
`protect END_PROTECTED
