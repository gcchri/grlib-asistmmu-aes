`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mrc2At2mZoz4X1NyyIO7QHHdijQM6YkC97Ld2JfEk/7PwwIjkWVv4E5KIzC2IIRi
yYsCBCTlzofJucCCB1qSM8GhezW3p+E/dN79AmoAoLenTKQhuzC5EAw7cv44lQFv
5JnOmJE0jA3fP1z3b0tR+OrothVXPAZ3H80U9y01uoAFi9mhbMG/7OAYP8RosctE
ZtGENGfa69Z60ylma9ZvAfsKG0CkqCcIkADQi8uYuYUmIrsqTMWt/Cdz9SPnQUMQ
UDRomK8Axz/MOzUStmav+V1snqX1XK2MxUCpa+tl2OBnv/e+Rsi3LVWyxvb9AkE0
BG5bgSyXlYIseUVtxkxjOpA5oRSlddNex19PUijntv/Ls4/onOANtI3UkJkoYrYG
K+3QqRGx9j7YYYj5cMwSaQ==
`protect END_PROTECTED
