`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hmD8FoBlWfxOPB5wO744v1zXjnhVGcsMJ7+hCB15cmgyIb8+Matx+Dn8Po/Vne3F
q2uhutZkX8X6Kd83foN8TlOju9AceGIj0vnj8IgHGbGQY1Tr669bEIFNAyJ8kWOM
OOQ60TrklFVb2UWkWoMX3VOxf8QhIlhLZ/CKCtx0cfPkGrU/m7xl2ClLj74gi9vX
NWTN273+Fqdly9Hfg3jLz9GQrhoYJL7bLVV9kjhVnc/bSpzi7GVZ6u6I9z1d9YHw
IV74VRozvpDcjrrukkgUQ6zWj7WkxWz78BzdQ0VXeYzECfo0YKkkw2MkYTXrYZFg
tyvlouNf9Xaw+v1C6ZFI3lojuUECTvufyqM03jh02fdFAziGRnEQ+P8rRxKRLgpF
gP2APJ8imHFDmpDyJOgbrk4rLKzu+bgyArT2OtjaIHQBXeio0YKk0+muuI9ZswVQ
66TRe9L5nRn/7l6fcUPe3I9E4RCF/l2AeXkdq6MRT6bY0QfY599VUvTBQ+uqJbkT
qR0JigjjaNxsIDX5zGgiI+SuZ6wd6mczrB3evjNSnpXQwSagtNd5+wEmmFYxpiC2
MeHmuHzqGjVQ0Olz5tZYypIQFQGqMf7dnTly3SHkApUvIcDgjxGkD7Jftg6llcMJ
nw9PmNRYVQlkitsGj76c+LslCoseHTPa+GRNFZKwGalN9SjMnrRJ9axqHavkahX0
37k/VUxSecTUukNbR3DQjkGBp6CLRKvuyrFzcByRmH0PldojSNDveNjIjOznS/Q+
/QM10jJTpFkR/jGNO1MO2bJb/BLL5CDYWMAdoaBKpKL6LdLvVPVNfUDN/U1KJ4PH
JRnuUJEVIMJMjw4UpVshQy5KTubVmQj2VW2ccDOi5I4V4iEFDPGumCALPRgq7qtn
iAaySchJZS+4nPU1Z7yi/eDacZS/yEZj4FVJaxtVCTned8l2oYsRQPXIV9WZr99T
rEZB3rqp9MCT3UXht6WWDr5azsv9V3NRduu11KxCOhpPHaBFIlhzqnYzEOSAlw+2
T6qN4XpjhqD4RTD1q08HK8EqlEozmZGQDGZLm4lCAXmFKm33s+sESe0ugsbWlS5r
E94VDkKT6/s7BlpiKspGNaTaLD9a0yyklIoyQrvzVVDj8A23j4DIf4g5+4sTeykk
D/ZpmdLn+B1wKTiiSTERF6ElZSUzWn0Jr6rw6Ibj4Od8h4Mgx1zq7TV89MiAoeF5
aHZDH76uuct/5GvsYOzThvZJk+PGERB0zked6QW3isga6DXeqBQ9azcj1bAdYMsG
R6GkJ2YvGf0WzszuG3DXLOfRofSxLga5zD8Ej5bzQTz64Zxet7dwxZzxONlQ5rzD
W8COfGU/L4gpd0pDyo6LLs7z+3B1wjJDWB51HybR3tRe5sYfUcEJxFvjdUpp43CP
S2xIwFFoaOyYEel03XsefkbYPRNc/rJUK5cLNlnFP1YsIWsK+CzaTFaDsUTYZVUg
Wd5V7h+0htLqsAvc4oWfrp8fL5wZM0G037iM0qfupmCsSsWw8vIJSK4eRnYi5Ykl
WTi7iBtX9rMG8dKDFfjNE8biEql5ZYXlRJtSfJtr1NeKlaNrYcJmtESUTvKeyNi0
3K0GxwwAvZsY9tFErHCXql4ICKnxJmL/vyVXRvCifwc4agjtFFOao6o8IM8h+vlJ
OV+wNgT2F0ioyI2XgnHNMwmDLztuy3c2cXQ/7TuimlBmq3DjwHksYGzP3jwzRp8V
CL1xpU55x9cVcFlIt6vE3sEJO8mHuVmXqpAvabrrEp2++VolBm1bj43zCXeruCvD
+14GpczidRp8ErYLlRcbsX8/gZvEur9PhPZ4IhF5MdEzCrFxy4TdVZ0B4RM1xOz2
IjPFcxnvV1mDFlXEjwux9c/K51m+dnQvRBap07turWICD4FdtSJAS6l4WSXsufXX
x0ESWJNH69JhVzmxGyMSv9NEAHnf1GoLTPU7YRULXRDqGQq9wKm3hNj6uEkHeVlS
ijO5qJ9m9f82zAWRNrr2aoHuCWWg6BWT6nzSkAjr+oEwo+DHJOACEFeLj293xA4g
jnMjjrYW1PgotC+V4C4mKxVByocA7yqQNiKSthdhlL4P4fDrlBGtYGpZNMcLHLhK
FXgMo0ryihHLUT/ENXgR8ysTuMF3D9BqjuSR+/RNgDm5lQ03XD/u3/OvmV2ILDMp
3C/Ldb9JZ+eAeU7ko8AsVm6x1URgWyQZ0zbH5UERYa9lZfkXoRnR2fq9u615RZj1
BfgdAbipC6pzIBj8miUto5hRbvh442ObEH3XVP0T/xuIZuiyiBgp2ObYh6u/KwCK
7rRKXagjAgXw2+DZtuy/LpBubjfgyHitzGF054l+S+G9e/Ge02tivG5GNgGCDGXc
mPZO1OYqCOhBPEhi1bGR2L/0u7Ayz8N7ctR5Mk5Mad79gQUtEW6ONAuVAD7+KFAf
Egv4POCh1pkyVDhhVYRImdIUj4D948Mp5EsdFBlfpH7xlE3zpm6ys0QaQlq+5Pmj
YNj98P7abe9zOpq6VVnj9LLGDAwq1gib1rFjOoJJ9eKY5dnEKzQ+SOiFYnr4VWAt
Ht6CWwKCYGv/sI73O1zRbjyPooq6SqotCMbnQ9ednwmIMYHudW5qOX9dWk7d0tYT
wRVDDO1+EBFtioc1jIgCi6u1/IbXekIVhZhzBlITh8EJj7mdxOmN7sfCy5iqcGc3
cwpf0aNv8XQFqZEAwbT4bYnqQw5mQ2uK2/20MF+uIUI0IACoerbGxek0ISQqAtuf
n/8QPpEZKT9M6Q/nfSP0nsSWM+MV0DZ8HEr+65USz/QfHAkgoMp/WUnoFCwJu0kI
jIbDDrGp6qNIZMxpJkNzRy+wc2op4Ztccq4z+bEK/74Ny3qrFyjrvDYGpuIqKeNo
H0jp65zqKpiisD52x2XVUj2rY2I57TG0a3K9kFrn614y7PmBv+gQu+odlFyUZL3A
krhRNqSZcNEvra35JdrOmF96JwSLHsfVZFhJH6RYTubcDVanEcGmLB3ew3Jssj0J
r5NwvrmccvqIuM6EHkfIVgO4DtNGAUORns3sHjo+zjn6ut0pvYMCOKTb28LVzGRs
6u9laV09YcUplVU3jfBTnhY2JMbawCdiy9NmR/Wgt2cGjzB1FUq57UeOs9cPoDch
MZWRkO+4ff6oLm9HasyjF/6LKFMB7rPtfQaqpnaMcRyfkQXrOdsjS89e5qPZt+Rf
n/Tv9LCul9f1wv4LaYfujquMzdVFwLXVxRT9sTc5lTzxlWlsa9RwCSuNYFgrimBW
wHdXnUFcHHBAdJ0zVg1InxYTOmLOH9qBk3m1c46Txnhal+hCnXHhneQIz9lk7OiT
qQT209KtkMRm26FipJbguXF0iHlJnnYOIWgpAtRA8VL0tkYQwuY+iidhGPwkPxBz
Ir2/nlCpFRfRCuAYxf1vgdsT8zmqIa29rqJe7JpPV/kT+mdcBlIAFzThGeY8CLqi
Eso0aXqIdCb/3ELjhpy/9QfqZPz1qPmYnDgYc6lwRppa3QM95xrg0rIY+/I5+Qal
0r03+p+qjCfQ307eaFI62hy+HWo/lKk2zq+Gp9Dqy+jxFZfGI5b8dDy1TEIxS6EX
aEafIxVjx6aSSpYAIhdnmZduXAHYcoRVvVvW4AcG3j2zNBrMl88CZeSyNzEbeAVB
p3lsnzchmcm856SX2gEMvNG1DeEJZsJU8e2nqPIio2RPXoFul6+qc/DCPOJbqL2P
M3V9wySbuAyJCrsE/8hVBFtpWYkOVLhHv8wape1+G6cIYgpE4o2hKkEwHb7Q6Xir
bh3UhSWytC3DKHFokoW1z1LOaWU4uAyKyNABfjg1YVCoj959dceiiXQ5R4UCMo11
fhwGADa8eoe0pXRCWZ84WHBew5D5X58LgTs+98b8xzObbvGj/8Vbo2PYS28bDibR
mEqOVt4WxSIfjmuy3bxaCqQu2E5coXtM9V19RUQFZKc+NPLyASulYco5Kt4zapGj
Dla4T5uosKfrKEPnsiMUtipmo/FOKcPlYF5JUetrxwXx87A98Cound6X+z9jLlGI
ZZ3fiSEAjVr4XP92vJf/qpatc04ewfw6hqcgLN/kREezb6n5UVJTh20YHm00A8JW
llMg+BvARoXtYLbGDIHZcJAm0/DrGOsb1+j/YMeJoO30ok0tNxYQD9r9+hAOKCg4
kCmj3tPqyiHFPJ6KECuCQ4a5zTsXti7pnVLw79hvl25RAxgqBjkEvarDmKePLkaD
mUwfDhQYWu2ge5EjCNenajiZOVhhDi41e2stHHB9Punx81IMVVgMJuIbOIc89/Jm
QKKlRevNlvJEJ6oOeIWeEwE+NuKeY8t3nI3Y1lHrEyOb52xM4jReEqd0Cw4ywu3P
1V3aWzn0AtSdhMQ/tFPnB4tSsS22dk45z/QUfBbTYKCK2fLCPLLFIoQyC2b2pUmN
t5zZO3sQynLZjk9/7oHdBkIHBnwlhHbyPBNQ99Rj2Z8Zw+1jZuwIrnYEzJdn16Ff
FvbD1nSqmpQChT9RruZb5XnLPM2s61F9FVPgcjr2moQSxH2sR9e7JEAVssJt5diQ
G6z4wYeZk8n6VAzplb8oae7vQzUp65RRbW2kMik0AZtOJj+i1ZtojcQ4Bu7a/9tG
1F9/B16VdJttX1eDVduot1gQvUTOSH777VuCA1bxAvc0LvJm3kMwH6F6mk4CnmvL
HM8xmtu87/oGBUGaqail5yCtgJu9kT0kPvrdg9jxpfOZtNF56FIfOskoPYmjI6Hf
n6mElZuQ4kbIxqIr17+z4FOVwjM4rhmEz8kK9AgxuoIKNgoLVBvwRUnr0Dc+BvSZ
lXFv9PvyKpIlGXkvlNu4vlqelZoTP2C2NfbvfZwmvSPixPyM+/fuFLq2knYwgLr0
Kt6MSGm1Ui3laE4GYL4de+dIvHzRU6YXScuZhiaSBEISkdlHBAU6zmO1F1v2Ss02
/17LZW3LlmGoC76K/VQk5KptQlGUcudAun9hadc1P/24mpg7aYgLlLsB6vANFSvq
7GNZwMwwlWn6dV546qW7ontO1EA6RfG2QUIx4MjKsb9wvgeUp4ilmL40lqDTZggS
d5FUoCvxKpj9amPVAXxHk9hun+QuWTsk8gKQeZAwexMbD7VaCk20XYykCk5+TXSs
hGqjX+ZtHXZVZRGH6PvhvoLH8gSzl1MPeyz4ez7pPGLUNNJI2eddhn5CTeCNRinv
OsYotj3aEtdQCHzxj+38iz+3cWNADc+vfhqfyktC9GoeoBaETnaaob+oxMbe+P3S
XbDFdmzwfr47bLv+0ogAiXnZeW4eWdbQg/tA2TuaBmkabfwCpt057t/K+N14gD46
kYbATcGAcSuFne6VPLEOaAcXhnQgYC6ihilNsTL+VdKbAjDy+JTbVlf5j6BQZRdf
n2SB5ienkzVY0A2vFmxTn3DVDTCnDXfvz/cG6S2VTBnLspalM7KbblNDVovFyNMM
AyieSF+jLuaoiueUL+Uf2tUhe83Lr9y6tfqrI+deoESQGm9GHn8kfaSLSgffOk2Y
Cz8qPEG3hzDJ1A3u1tkNAiNwJCMmN8k/Xw8izMURMpy9x7uBlaygKp251FRgNcbR
cFQowQ1nzZbH67y54fH+1xV/C2qXBNscnAAW85THvtb7edPQCIRrnlCq0omMtLk/
wsxzHxvENuLHvZ0u67QTRynGtGAnHviWnPC9RH5/Pjxfl7oDY9uHoNiV4Ya2ZSMu
aHDCM8+zhqD3amdukVLUQgba27BrZCeVtwVdfx8sC19X0iqc0nUkafIghTkCkKyv
FvUPnR8PyArlV+/kDNCrMZVKy/S9pqTEetDQCSeHevOr3ck8GPMFTgMZ9v0egqyQ
zHk9S8e2uQQoTEGipsTAvT2jL+an4y4duV8Aa197mMNcZuHPaFYCtOvPH/nIviDl
e5q+6unfHCXmkh92lXoOJrVTu0y2fgVE4Je6ldlzw3l+T1kHgmNwYVab00+qkKXk
8+/SfN7GCOTnQaIUsZedQc1ytA9rdRZgNuy7rPfaefxeMHA5H7h7aUQmnO3yV1v1
IsRryIt1vteyfqXk/TxOaMdAwylhR70K3aV5uJkWYDtCLKjTC1w2HMHusrhE2SGJ
5i/kTpMMAy4TotQOWS9JouD+KVtUCl1wD3LPgkZ+H15NkXfF81ZHHDDasB2YOBFS
F7GmW3QGSoUTHZhBuDipX+FCSG28CVLadxHuWjrWP3sqNhWsVhdk/KwYIC6XTSpD
M3Ruwgo9O/0AaALZX/zgGbvzHfdi1D/D1N9K20mvO9JaVbk7l5PdbGEsxtiYD5XQ
4O9jjn5p3McITgP1aZ5BNgGe0U9YlRYO94B2SBMCaDsATowE9yg9Z/gRgHw7Kx3x
28rztOuzOYOfRkmMTkepF3Qju2BDq7bUFbl5Ne405WhudqvhWtanen6oxOIOhNiz
5qEINh/vtCJpM/xipszNklCSXvgaJL/F32HSXT72fd3Qwk9JpRcw/9iPUP7hFv/3
n34XvfqB/VefzrbYINIUqd2tAgYyZi0Dy0TIWFxu4tQElyOXNWO2nE9QMJSpcgvs
HOqhvt8Ps0dapGN1zTbLwpxJHETXJc8UxId0BP1/JZhF/P1+hC+VBipKeNZ67EwU
fH9JtrH5hw5Wk1+/DlX9QqSnI3W2arXUQtcDEQUJWCuR/mPDsl2o+hMf6MkDaCtX
PvQg1zMzgQRqwNmijfA5HWhwLu+PYa3OTtopeCQY9W9ReQBT9ruJF6njVNORQnOW
mYR1GJI/pP3lwM5oS8g4jWPzmnrlkARZvOcnKm0Ced9EG1evDsRT49/4iUw9KKaP
NveWMsT7yi9zTyif/d2nwxuEbqlXI1o95EzHr8a/3DMRUxWihJTgSpPtJUtycYaM
4YUBh9efRTQzLzOeNOu0o773zvdVmoNCyE2kK+3oPV8xun/+BK1qW4wh83h5a3CD
ol0OIQ0NyPNrCLwVTtherH4oC+/b4QzOTkTC3mp+KBENxyUMQPFFdoMcpoE03b/r
vBsY5r17sD6grj876x9dvVzR9xlhXFzxP1sLyJ22cv5B0mzD0nmJA6a07Oj41/Xv
6J15QlY9jWnGMgAcxBRVpvHLY/EekrZ+y+jDbQchn7S8+7D1ulafRpTOmJXgHi7z
RtF1i5PL+ke46zSJYaNEposPMr7jzNv+JK4wOSbWUKtXNH+psrkLRWjLWn/P2S9a
RUIde/eHt8SSMybsjg0vzW0m38QEUgfJ/+zHwiWRE64AxhwMCAkTqQZFkR8ytWYK
Pm7EQRAeB9KgT7W5LfTDQCKtJBf0L5gSkSgImiod2Cn/ra5oPSN5FHmwd8axKIe1
qAoY/RsL5vKQaVxxVWdzA8XNM7Fcv1Dk0nHh/gkgNw3hm7lkZaZlRZYH0omdjzxv
v6zXK6FXZ9mqVyLBB4R7mBJVD+nd5sanK7wFwXI8QHjasSZJwJIbSC0gFxK3s4zR
XoNK7/Z4uxNn4btZ5kdcIX1G1WwwyvjAQ7xy/qCB0wBMVTB26TSn0B0QwOTSH9Dw
JSh/HzuJmeN6uuM61ysXQi3WJdZPcw49wLiXpvKUdJ6fzdQRIHqhaM6bVuQ7x7O5
Oh2XW6dXYj2K7ctMTM8N+H7gtKlNJaTFs5D0Su9agStZ4kyaDkKq8eUAZ5qqifgM
4MqklkH9SgOySZEsONjJ/xTLQitrGXot0MQ7L8WpT+3r3X3+7SyPjcYUb9W7qNQp
fPAHhQ5zK0Z2iT+tbberXXGJePkvbiatDPlGnAKyaOeHPUH2B1dEyYSqnWNzGVqZ
OPfHkWCAdXK6uYpkvNA3dkSM8/zuib+6N4lvXpT19KP3OGkKzx1PBpPcnYiC+SfZ
AuAhHlHfx/4uvF3auN42BloZEOIdnhcUxNUgfy7QfZVpTGPXI5Ags6ncqGeQjyyw
MvTeh7JoG3ogYuTDgsD8u6oM0oylFWvLcsVXGqEDqLxM2LCnjmNk9Xrbfei9LCP3
eTfa7ogt0R3BWXD7QliuY9sNSVxsm/+kmZI5/dm70LWlGKKm+NiuL04d2S03Pmw8
vHreabeAdHdLiV8u+04/vluyf6WyHGHTPL8CH/tbNseRGTJRwpsj/tU7kkLSjckt
Y1baegIeVmHWC+b3QRjS21q8GjAbXx1rtZSZ1mMmYh/uMtl0GChNfMy9WPTSVZjs
958PMZHIm1NnkLqAiUqlG2CECKTjvgaF1QDjJl+ThRIAbUz5XvTrtkmc95bgH3OK
2Pqb/be4/jmOnwvTchtJLYvCOuEG3HvOSWgik5ai+1ybEdrawZHEFRwiNAhoBtul
HBRUDxK7hemKZD79cholHz+KsEiSG5sXW57Kplehcdd1zxQHlGWh57fE3Sz8poDc
gyoHN7T+9C++K5nl+NnDO83/EaSJImp99VoRWDLgegUVvJ/BKCArw888wtn/4ukt
ljmOSWPdCOde7Z3GZIJWbO+eV54uxoN+2vmuGYi/NrSbOARsHZCNXLgCCpPt12be
hx89uOnZt7fCHntxIjV2ZI/WnDJ+GMaIqs+KOIrpIxj2mWLc+gPr2TKVPDHiXmXh
NGsXS/uzrXNFi0Ejo4lU/ppt3OydVvBhgKOdKlyESiYj98LPqRugn9TpIkyORojp
4k6d09LxCwygl4gQ5asJwMOJlLnLaqhhAsP4IYldNKcv6/duePREf4Tw2XJ8b3VU
bof3qZk52dkunMLMRmrHpfdZwsoiz0sBvlunUUejbHL9ABeKsqtygiHVe95n8jTD
aOSKoLCLI9/E+Bz9RfbEKEFa4DLJZw5mB2J9lXsExI/IvmmVWdjAaVBvKT11/gkJ
ew0+XyMj69z+eWsDAo41vbxr+AF3Ap9jbzZHnrVHg+YwOipXvkiEVVjaECOeJKda
fkLtv5Y0C1j3unrf5bqC/xidDKRPJX8jW44MVMc5NyNyOeVM5PcHBFwHQqa340xj
7x3QEWGLkGhucCLSN8F59ixOchYZGDYIy88gH4oHipXiJdEQ3CW2atEY2xWT3LNx
8LDKtPEOPQTJT9uq4i2ktSDQAHCfc1SewVre0sbIFcXOK9GnuBoXCNZmZsmlcnb6
Y+OFtfzoQqvyrVGCfhu/Za6fBXKhY/TIfzUsu6gI1hIuU8wEQ5sKxY++YUTXB+aX
BdDFHxqOmSHJj1gOqKj8gj3lvv0Wm4xrSX0Fz3kURl8VLAdHLTg8y2ryzsdhpSz0
X7Hes+3hCA1B6mfaYw1bylfqItUKbapnR9Vh/5crRE7cXtGfiyH6eeLCy9r0Z67d
yDXK9Exn9KBrTQyMqKBnB1d6AL+lp2qlhORfySNKCli2OuhDxRPSaR0W96qPJDlY
Qys9/EEXlUvidE0GQnK05V9p1+gy1YVKFsX88tP9j3hLVBgu/mSX1pwd0JjR7BYy
y+0lHEUsjGMeDGNQ8Zn72oLuhg6U1tSvMHxCJpL8yXVlNM604852XkuasjmWs8pg
3WIebqEKdpENNeh6MiAQLGQqWaa0mIhz9qnWSThKsd0m/OT1RBLX4ybXkI+BOGmg
ErZDkiki/phYxvxP62gFPbWNv+aMEVZjKS/6eeuYtOJ49XvLfDo+Z8YrJVfHtoRC
LNpcbl3zPLaRtH8rv8cyUqc0fyJ5ZAlvE0xjc+2SQtc8bIYVYC8uRl/UrrdpifEY
gzuZhoxe7NkU+wU5cmRiTk9DaH8CaDVVITwfpqVABpNpvYTylIFFOn4tibpAcW4V
/qklGUwt9gc1XfzWGrqBcugN60hUIm0bT6vS3C0qBmMT5AtxolpDJ0qnDT8VcmNL
oHVroFiTnZk6al3MkNjA2LGvyDXhjf8YWb4CRkvVRnXl80zW079wYjlkalxFko5r
abBKhoe5BIfGcHgpX/+kCt4+ug+BtShfJUxiUpcT5Heq/i7tCtrU/E5lzTuJT9Fl
AoEaYq566u/PCHbCQuNTenUphuIiPe9l/Ldkg9EmSyumYnJRev+Yxwq4jBqxZ4o1
ojwyayY8KrAvzdUgmjFhNMCrSQ3CWC8TY8O9KPptCYCYk1oRjrNDjp+Ktwjq0tn8
U2IKOBgqInLESe5DjwkKaedd8UM6//lkLGr495pJA4C4NjHfLHts0f5XUHYUB8ju
xsfyuXm9n5JkszdwsBrqJWidstNM5qkfu3o1jsWQ9cwEz/+Aor4MgG6HH21wIILg
rK0JX87ScSGctQHgje/psYBXHexaRcVO0CiF69zmo4hTQjiHDfa8FVob8X3YaRZ/
5Tc2Elau8hafJQhKudFpWK2E/c66CfHuws/N5iecaqx9X5C18QOT/P6FfYBc37rC
rRNkR7j80TQNQKmOgONrj/YRflJdrGFdWYXB173dXo/5G7TR3JJ/XQB0IZPQiiTT
xMxWY0+Z6gxCM62YrpaNyXHWovbMY0DO2XVPiwHcn4v3dnW7Qw2rj3iKyMtN+LFj
aqd+9Sp6o+Bt3FUTuMnP6XnQVF1VCxtD/jYVorBZWPGlG/1q4HbbmQbRT7w7qcDH
DB8/UGWYYg0FIOxbN7x7jzdxl9i1lRfjh/n41jibAeO7OhnQbSGOOXWQY006BCpH
DBI36bqx71TSCqcgvuKMjTXs1/FxVAkDB0nPNWM3f2KRiRcK5TLVZ4WtR+V8pYXP
VlG7pv82Boaxrf6lvCeGoiX0b7kuAI9NSOUOQ/RR/gJAOp7ZwcUaorVjytKLs0/N
SJFTf661v9WGW7WAkCPbDBthJD1EGjk1DPUsLQkQVMI+VLUyw0yNRfy7dcUaF31s
xhREs6EghwJxdfRosPNMm59hyruyaRlM/nmXkY4Ifk7aOwmOha7wa8wPYiOo+3i8
q0MAaCeIZ6wgOCJx2MsTvDaUqcX44pJDnUrtkOgIBpQkd2NrsgtsxbWp7msWFAC5
Dro2GWX7jztlgrrJPQ6QBRzh2E7y4toUJ9vctcAOqnxF1i1EytbSnDbQtSxPNMaR
8SCtjwrhOLppYC4zjtr8H7baocsk5EueYv2Gh7iXHjU41UZkIokdGAAayKztuJ4W
9+tHgCbBQpEf7rYtymeIJnTueSGOGzXlzECswUgWZ5n000wJqR8vQnZsMgCaHHIp
tfMgY8xNrYrNSGrq+RoFsMpdzsxO0Yx2A49eDpI4p+XNCQ87b+sRCC1/jIedHQ++
LJtWF/ThvnHifU4gSNeAT3YdomeHCIFtGqX8TRg0qz6ep8pU28DRQCc7q/xfEoh/
XVMoQNtNkNf5sEUB77vGtY/TPVgjCNHDxxrBIutpGdpM7X2PQgFjI2hxQ1l/d2GU
56tad9jSpIzBjLkgklqfcbxjF1EYWeWiyFCdatjL5DZrS3czBHeuOo4Wml6CAyVN
25S9TlC1SHRghS+NsSDLMIQCQ4YAX6kFmU6x1W+nPOwnUy37t1lfMlDOH8F19l5C
F3d8mwq6gEw+mij8EG47aiBGAWm3WbwUjG061EsVH/JHvvRXlOSe3K67NAqqdrpV
V4jR/yEvMwevabrRINd8QRA8ifFcn8rcZPXBRRiG2CSt1R2enjoBcVVLH5X56twn
n9FmhDr4ySrqi8ka6UQa+9vSPlqUljQ2EEy9GtC/PwFMFnee3IjIxTFnQVoxuei3
kmqCQrE7sWeFP7pe3Phkqe2GGsLWSHGTkAYDCudmbfdOiEA0Ene4Js3r75SWi4w/
PgDVzoIpGZVl8ira2F6JYKPds6LkLkS1dZaAUnN3jQLK2xjGD+q5UbdeL+ZzBXa+
IpErgS7NdUJMScmPjoqYyiDwu05l7W3i5GMGygqX9TPaIQDHQsFFej6vcMw2puK6
RD5+MuEhIT/hx66OsXfaShRWZaC0nMjqr9+Crkof1mndJiv9L5rjIiOGkrCJTg0G
YoN94p8KvGAn11S+2dJiz5yIRbwdDEIh+MVmQWtyWE66uYsrD9fOiX54hmypM1li
uFt+WpzkmRaJpSj0BwmE6/N8NkWBpDv3SdORVb8zH0sZ0Q7CgYloZu+h3Ynkfy/j
QnyJGS5L8DleajBmJy5oC/z9OHG9TvdxO6RkOst9D0QDiVx64pXEteJ26F1gXggn
6Lb1YxngJ2tK21lVQP0nUoNu6ZsPgHK1o52Q87H5Pc9UupYLMiYEsTZI7TIW+grv
jK2bjF5mOr3O8N7haXxpkyoa9DRcDPk2OTso5cxBMf3eEc4Hhcus5cIhJkzLFHvA
R8wYftZtnIwysb5IvM3ZBiIoQKrEtdCANm7jXBzNYJsc2jKaDQL7OMWjIjVUbLi4
6CZtBxQtyCVWsHbPGRtYp1KrR/LiyocW1hVaCpCcSeQ8vObWJnjOZWJySEFdQiox
B8SIgI86s7O08YddAnCz1mZ/IVrnn+ctvOKwCHXRf3cZT4eqv+VIgMNj3k1+GmyQ
K/EmyB9uNzIRJqJFTK8qpEZ+8SP3zOPykBtQN6BmDMAdnTiIBoemnpY35OsFjpL6
0McP15L5wCcCPPJ4Op82vz12hrp94CCMh7edNt0FbRArEEu2Al/c1MxW/N4IvsQi
yfg+foucXXH4eMUy/qJGmnQubLhm+O30CVMRSRDAQcyp8AMtxwozuVG04GvUKKaY
b0kGESOngFQVU5z2Tpb2NaXlusm/vbIoST/6n0eNHyhdiQ0QMZOwK2uuim5cho9q
7f2dkTSCY9HIjIIm6C5ECS12c+wWyKFMR35oVLxe+VGPxbcQm+RG5uW/rT8RfyVS
lp/4FkcPfpi4QvVLJyOrTfl+60YqjQ7XGsMWEUr0zfh04kYWFV4rge17LtIIhBNv
bmrY3Dyz+ewJWqX+khiauAv0kUR9ydlhSbQzUdsI9dGSnv6Bq5dcvgoBR6zxF+Z7
GNCeduGQ7XI9CZIpptHASZ1fpN+kKycKTNV3xNp0BuW4iRTGH8aXsHfgSdVUGA45
UjHIDs7VrC5pHazEFFwFMtTBTLGpNL5JaLYCGEFx3v8t3Ed3ZTXn8jp2CXkQTGgK
ztOxk/rAjXWF6XsDY//gDoxMlsxWnpdvoMmkZl1m/DSYUMbxOKAlEELVGnabJjZo
Xz3RZFXSqtceNZXZihxyA0KzfwUWx/n+FH93Qr9oVL+SG9eXYEWFaxflr7aR5lgQ
9rCY4jzw2mcmkps5OUk02KAZXDv72m45LnkVSLgpkRcXIR7nwVV4duFe3G8GKOKv
/xzScObBL1HFNQT61abaUCPBR8L3d2iE2y9jAXl+bwUhbUGRuPbV9HDHn0aK6AMW
yNP0+AH60cIaBFJDKwidmHXwlMbtRY0LbXEVBxvWqHBk5gG2J1gPPUBp5GApff1R
ZNIU9iSaDuh6NxN+xB60rP5BzmHtR95KMqNhE9Z72Hm9Py8oSbeb55QX2ZS+NXIp
LAfeRVJoRdyTcOug/xEr1dfDy++4F4LtTW9GzbwdMGhdVOUcRKBm3eT5CL6xAut/
19hPjMYupZXgS2o7YaGIpUTMml2YC3UHOyRdq37hsh35WmlCKf1HfZNdH8eyze4A
LO5jH3dLJ5BVrBhv/706Jfq3RHrJ0D+kZWQ3OY6PFCtLKg46ayuanDYBd3n96Rib
U551thzVVLXkvJY1T39aaid6QMO/AMy0PsaONxdLDnRXV5WcPxwkotkf34qf/sfg
oTlPZwOSjzFNII5F3KMBhR0SJhhCI8J/mBBRjoSQ+u1vmr1JvCjZ5nJT+EAVSJkn
ILBQT7i4lsT34Cg8THxEeVzoJ4Ak11b6GfxSp+GWFeZe1jBBhNKs5zM2tEtWGWZ+
obTJMGyY9iJf21efDsYPh4lGmY1D0uUtLOruoXxNTHS0yazHbVBF0m94Ay83+FVP
sJZZYnpYbTj1GBgyrLe1xJOjvNGb828TyDkW28oHovhEYmlwukf28y20KF55ieno
7Q4DRQaUN6z+8mkN5j0qAEHGyvC2mQU3PGDl04kz88sWXT8WZpP6D6NhTgba6Op6
9ojHcJcgU2oqESvN+PMzA/K/nkv7vIlyXE70n5ByVqxhmIeMVyQD2BcoMFYEw9UY
IA4+YZ4WOzzVQDQkyp7BL7Zwizk5bEORF0ZI8run16BiDvT1BudnPB3zu6vo7Oja
ESrGUa+4L+4sQC0MW2m/jiPc01ktkWHqTRfXZibZsGEMzbVIEkGMgtO6inpU8ps1
ZokT0O7Phgbc4jXX3OZSupOCnSvTbI5+w53bz65mwOA5rqqldnqkDQZmt9a6Rtou
aLoxktc6B8sAJHk1Jy+wp17Ms4vFn9GZPaRBnmTyufepKdWKRqMZH6WuNBdyCcv+
+q7T/STRQqgSNlwiy+w3moCTIm1WNN54xim6mbvD1BKl35p88+wdDNWhtDAMEzSz
wSz2KugrsvbTypL8mM8q7R/5oBzc+1yUNEsxDMoaitppQQbhTs+BiRgA9dUemp/4
8HYTFKIGTmRCu+ziX7whQThxXRk+MLU9Oa0bxVV8pHHEZ/ZWienQrUxicaIiAvOy
YOOiWiPNb4prtcL8pW9YxtLD4G3wyvrVm0wL1qXWfQZ4oyXIRH23xj+7GuhTeaMy
8Da4Mr9CvMBWVK+31awwyEhT53PmdFJGO1tH56Smrd7YgSPYRRv++kjpvndFC0Lr
2WxyWw48TR3iRu9WG8SUF6z/JFclrk4aXgYGpi8/gMkQbX4/vIClmNOEE5T/M3ua
VIvjc6XZuGpQsNHMQgUYiA2FGh1bJqUQr0KOCcsy9JDhT1ZQ+Hu1wosngDlD+Ih9
kWnMzEps9nOaj16WC/lM2K2v3iXHigEbaqUxPaSAjkizo3EC6nut+y+EdfoN8nSX
3fOzO6TjrvSXxTg+tfAyasvxRAhkGwnwr8mUKJ2pMsl+9b+sFrfETs0TJo7VOhnp
lrS3DsglFC3qJ4a2MkRsGyU9xpwZPzbg6ag82Gn3r5XfEH+7glqjoylkniqWHVFK
+jd7xwzUlu82Ul3F3dgS5nLhKvysXrJblnsqY1WztIiACcVea18dYYooGcEIt8H/
ofbh8QvwMCJvDKJvs5LttCJ0ozeKKyuI5PqB3jWYZ1S0tFmr8dBvqFpM3VERT6Xe
DViqaiDx66hO0yK/8J/2Kq05L+eDB94y4qLFAKbSyvZHTtvwQCFIvwdghUtYwpQZ
Z5Pl/0JJmQf3LFPlVuQQzk+4kAfOmJ/7eUwLsi8aV45Ho3Ez/XdYLN+jaKfk0tCz
6fZHKaDTA423o5ac42dkCA6O3vzg0YDq71qLDbD8njLw41/6zVv7Chh2HHmIGvrX
450l1SrUSscRuJ65vZ6LfQD67UzzX7Nv7XcUg7aZBpAsNDDBkHAPbNqtTgrCGv+1
MPnMoqfiRxsLm/Dv2jGhMw7AdWqaLfwIfqo4+0RrJ6RqqTrXwwRQUUKkhYPk3i0X
B6whp05wINQ1a8XY38WzDashoKH1KHEEvs96nA2SuI3atBpT7S+QOvRyPUA64eo2
CgkxKx3We4rAZzNk093KCDrT+qj7dfhFbtb85+R1edVhvQKA8cIXsc6KjhbX+tJS
w773hxy0rMHa8Ozgn065IxvvKfTkOTIG/RSZWwWWB18z14dB3UttFcFv6a3dRxsI
inuVZXZU9FtXSjtF+jGXdb6B21J5eSS2011cAKCgzv+PqRCi/YWsdIaY7LsEyyOC
/InfMBamckGsRJP0jAW1oLmuoGhUhj1BsH9j3o4P/xrgpP2gQmCah6oU9i+ApDl+
7BBqzJg5LGS+61Nmg5Zqb+AkrSv0Tm7tabvrKI784EnXDeEzXbYAsSzRbCxBfguD
Xi/yW+DjefkJF6SPVI2WTYJDLl/9V4eCPXIaInu1BEBY+RHeY5o/zjLES5UG8SIP
Jw/yR91rJZNFK1fT+IEGEvvQ4IIvDd+5ThxC++D6Z0wVZnwF+eACWYY32IpypnJJ
FPk6FPxYaRsVamMxLo6QYnwMnaDhe0ZoGQlqUU5ddieXqKiUZPZDMkMiwlBLarLF
BCHJqTn7l3lS97VXDLN0v1JWzmWlJajdJ6niiWGjAXMVKxfBD31lYpq1VBQu2CbB
Sof0xn7t7yKCiABYmF1HuQprfQhrwmeOg+E/T164Qr7ZVlvBAUDgS0UKD6sdpEXn
yWCNW1rMHtbxoZTEfxnJcG3yZ6xt0ELGLiYYsXRsfTVHqL9d4XXlDIxxZjAD95CX
Z3nWTIoA3yQogs6tS9xE/XnIM5aM4DaGmH4NAYXPt3mdghckGRp9VQOsUKCYR7Yy
nM5nsLSWfW7f6j0HziEmBu1qWEcoZEjRvUz4NHVhoQN76H2yHBikGzCwKreZB6Io
oXc+siI+rHi7jk2gyuwDgwGpdgdQ0RZ+fW3N5sqa8N5uwDaut9QTQc5PGE3k+Rru
pr4E+1vBqoATGTqBzyOvtHTAE5IG9ig64l8TcMleXKOnnqHk+kxD/5b8PNHCGOtV
Z/L1AMhlndHHWTpDpONipwdl73aQOZDkEdWBOU3LB4iQHXXFLL6fXGrNC5Up8FzA
70FwF0fmKAN02kWtxAhQ162JXxksa4258pfo7jEPbvw5iOClhCDBZ82ajatTyTk5
N65eYUOS/PELC+YxR8UDDgYAozHkvJRPmDo8P8WlScvwZdVTedAEXqwJI2AlXXlL
dlu8HnFhl4CxwMQ1Yra5rNPcy9yfUT54/nuP3jwNHkDY2fjeiBMYebS6EORkp3zY
S5hZpK76PSuZDnhxrYSrCKglybIpFgrFlYkjLAkUCCbmr8/nW5o6zbPkN0f2L3DS
dddhvl1pymQY18h2KCoM6wFpiLM6qnnmK41oDUtFd27VTvjN11da/5ViwY8+Uydr
oxZC39KDlsVZh3TC/TV5bewFesnWYg96USR2sWcnrMGx/ZqEit/7lLyaLHGNSdDz
LNuwkkatHK7mzh7x+SCvH5oiiJ7+fVc07Qr3n3qWKsUCjEr/0kfwYXiC1sGdO4ss
h3FnC4+Xm1mB+M2Qkvei/dsMjFUR8genANaYK1GgaKJdW4+ewUueSDaCgIR07mPQ
yutRw57SnfIM709NOpugSWqDJ8QIrqKvV/6rQ69cRIEzZW6No54wkuSDu8WRKrO3
6lZWKyekT3aL5tu9bPfw2mdcyNZ5gk6J0SpFDG4e+vi1E6x/NuAy6sy2cjiw5ffg
4GZIj3kZUgI6VKeL2xnN9A+KvaJ2ZLX4gqjyCXsOlCRx9X50xkBCi/ylRiJctBMg
rvGj2cH3zMmxU1R5YX/L51KRfByIZwkEiki9QYMja3RP7qtULQNxl5kOd8iq+qa4
UYAX4zE//pjLpbF2PahyOLxKygFRXL26SH6qVNGnhC42NEAOWJR5IkNHRfJWoAJj
YE6N5uUeJVgtGV1Y3BjQ9pc61CsITaj4r0V75DaHvig8kGN+uu2ku79WreGtJlCj
0lYr0D2xJIqJ2GzfvEUMegBDUOVBI79bhRffh5LPBZ5byXDQX/b+6LJeHqHybNC5
BMhNK3G3XdUZhkxsVMjGuyd3lNHCev6oQsE1ae0TFdZZN9wIpjh/8pHs31un48yv
hFdNo0oNjWICl41q0GpXfOfk6RUVm7ejXcOPdjXCaCdBXawnbRBSA6Cvgh0r696P
OeyFNoxGQa6FdxHcmU+yDyKlrzx6zS/VWlytcsDWWBeZcf9UZGg2BJhFqH7BwGPK
f7CYpmgRzaAxuqJqOBfP4r47cGu9TO/ZgSmOs7ivfWeFYJhw73ZZXiUe55P/ktcT
Vdc8Ly+r7uWViiY5l/xeRiCocusJWqRI0qACDoI5NeXQw8GLiAvSw/dDvzWqzxYz
P92+ENNN8j0tp9NhrEeT1faVeTMkZvRn1oglAz6Tt7bBLe5aFswY+aFhuFu3VCPn
PsVFLA1pN+gQuSZVTv/lJzRza9hnl3nnVAMpE3+BML87xotbRPsHdQ7tC3TjGUYW
5KQnltoA3Qsk9aiAbf2WRXoJgmEyULiHahRP7ZlwqZCFnw0MyoTi3GIKOdiFQ9No
Zd2h6xLZ9e+P2tidZ511/xRz4xCDxKcWl7lFWvf3lw4NG1ePC6lHjaF0vScVjvmS
ucUQSfJtqhIdUYNYrIhFVB1+jNiuVWNtl7Am1yA2sBYY7sK8Azab5Vb4m0BgINW1
FVgg+cxB3czN5P4AFx+nGucydm0Jp+KtrehpGzcCa9J6aGZnbYrQj7LjaL5TpCuz
ndsLHal+D2/h0NoPwonTUxLLVw0FsiMcNszCm7A+hAIgeV2oILpQ7UWm5qUzlGbu
nx6k9o72vC1jAXBp4Cep3WDzJXNsUpXzOnqUVB4unCKulHIaVvkBOzrwbpOaPzO6
6V71xiENYeS5hhghyDyxthlsfrMgLJyejp3w4GGSHJEW9tIeYC/vta3noNIoUYf/
SLK2qblBZ2aI7H9K9UZ9FLVB5t9qN/lsmRxs61RlWP9Tl7KN38Xz5DYNa70DGwd4
W5p2ST1IulQhLhe8etXWYa7ksJzFOnxxNfIIU6nedlMB2Q1kKyhQ/mfTHt2h2Xw3
eO5RQ/i1cnjQQTlLF8tZenHuN/rwU1TXVZz7uKy0sKzceMOcXHlG5Pu6fUjVweim
JaqjbxXr63Tdi9q4rkUgvqqG4B9Tov332oU43qXu9bfJUXzDvG+KU+S59TLpHYHG
0bUuQlAcAU/begwsSUT61d5yv9lmmHHF97MKboJWvqHwU77loQMQfxDwLYPkhAWo
8avg6Gm3aebcGOOprXPSQrAkPmaMAZXPpG/ohfB1fofjGbNucsWsQdoEWlO/c9l+
kBy3I/LlTPKRE4AVupJpllcZ3NsYxkAwMfAUAOM0v22OSfQYv1gzThyF4IG9Frz5
/XeMCeNTkFhg7/vjEtgw9IpoBM7p0HZ1U3ZADlfADBZOCPNAWRnY1mCcOFAlYdqx
5CWXC3XfNJRid1cvs4uqWMFziQFk52L/JJ/WxFu2sUH/VRcj2vXGYXGX4YYRJNSH
oHwTmTRazdc+xu4LHoMGK09Fejm+HZ+BfWuzgsvKNM4iETUIKn7xVwUO4Si4ywjG
7Dm6KYzdRsmUJIfZhz77x13uMYm4SIEjwKn1vxQclELTqiamiV5Lk2u/iplBchG3
ZXSwQ7SvrMqfgGm7WqWXuYGaAqy4UkQ3pH4WCwvWx2dgho1450yduwxOIDHJkRbO
u/sYoec1i31dXCaGybMOI8BpDOijAMJJu3szAEorlVCagcNKPWbkKkkIX5ym9vVs
2g+R7s+s8W73Uk2qB/IDuaOJwl7ZGNAXwLS/Kkgqj0pFPVTV6h/08thEoFoDmnYC
zFvIIFgSkUoz3wxOeGs8dQzD4Dh708DE3vgaQV8ookWzuR5iNlYek6Hwg+1rVvL0
fIcX8cwvZ84aWSdJpZYgDJfmaZQaSSxPaAirHeBC9t2iZOyNCp0BM08JnYV9VWIg
BydgNS4yUiolBQtpl2vdEch4Qlr6u4aZ3QiXulKxBRcFj1Ig9VMLV0Oru9BYaVm9
Nk0662UNsfSrHAlhyOaTav4ckRJLbyZcpTn/AT5zw6YNPaAAnu8jNur07kgW5JbT
6h/RW6S8KdVB54lbMjUlPHuNjcdFvJP3Yp33bzmSa8r02o4CZ1mCCTjt9duKok1V
VFMd9+ighLaLaLooRn6ep44L1n32RA+cJRvmL+tNMpWsKvdwfs7P+M5eU1gwh83Y
VB5X5oUw9linabmu9ryv2b25ynWZgEqD2NFmI5gKsItsIpEX8yBPaCJyfbjcW07Z
hgmjwrG7tgX6/hgMoyXaouiaCxrPb4BDm7ZkSMlErkijvfi70/YNZkpzusAVAzVS
qRJ6O5dDapvIrWvhzsH+/ovHutfzeZMa1LlOl5xhJaG8nd42qIM68/05mEwgTQHf
iLHlqpWQIFi5HFuOGOPyn/jEKhJsazydXmcWubdjD6+3J4SGlurYoLwXsxCWyVQC
lVcQq+ZlVY2CdDLPhiWaMt3i6SRC0jPhvzEEKeCdgXwjZk1qpii9dX+eyFAXapve
MnExw/LeQvvy5BwLo910v/fij3HkqHndzGPbQpqs6pDZ4esPpvlR+aA7DAruGy2M
62eUrvswuc2S6NFTfSizE+gTGn7nzDRyAj5Ji5RDSQfiEz7EsUbnjSfNcwANIqiJ
QRtqUsPbt/5J8DoCFq06KYi+/1BAEUMyC74WAmvXWqr4gnGEWLPIkC16c9rLL4pX
Dga3R6r/uwJF0edWaHaqRMXL7m3yDVwS72kBr9T37Wsb4U83GfeboVhz3JaJDjnP
Cuc0uVx6Cdql/E5Q2zuj6riNzYzCwFusNNhLVgQv/KhnJEHBHEwj3YTsbBtgQkQE
yYsuBgb7I+X8Ob41GgzGLHVxDJtCbswydJJ9o68a3iwV96lO+2kpVl+xnC5jl5lN
JH5kuhwCKvl0DxM7t8Vo3l6gVvZX0TvEiblEIRVhYIJK7oa9rMtkMGq+TEIjGlfp
tl15h4SU28C+1S4El8yMszoFlYKLk2Hbr7tLrxYkBRbHAc2Q8vCZ0iN8+5315V6N
QbeLO8fTlfhynUHuWcrEXOLW0HQXuM8k4jA+Pu3lCesBk4jnKFVX/a1XV3S8AWTv
3U7lx8cZFsZtTjmNE28O6BufgIAZmMYrkLd53NKfLtVrg3HRu2hFFkwY1ixhF0tI
ezy6XlfKjYHUO2I2M3oZnVeijRfmbkWdZy6MGgKexoCaktAOucZP5dIYUsPQ0NZY
9XDos60kvFS1cgGgloijjxxiiYkBFmV3ReXKhXDlw15S2VZdI2jP6NnhF4W2H1Ct
3FiJqgzkT0lVkKAH+tXEZ0UnaQSGp6cgqoCzEo3zKFgZAj6qRVkEy0jvVNxTttYR
7TVm60hn4nlsqJWXX2n/T2oFq0tAeYoOxz4WsnQogsV5ScxU2sdFBsQtlUFXfX9b
RHqrUcGFVB85DgujTXXJv6yLwN9jkSY0k3MWaNjx7SHrHj/U9fWnHZPjGpUbH2C1
B4RhW9ixc68pY/EUm1INRnvJaQHNE//zGc7W4dgwp4MXg3rrnWl4PcEdR+Mq1NN2
886ilb1Oo1GggHvyq/PK4SZvRahyNUCDQttnREGtP6vvkLQGEc4A7yqcBZxsoxJC
12s+0lPQFRdshhStxUM6uy2VJ9zP5YRnK4Q6HMkiQZBYxBkHThLXAYAn9uIxG2qL
9qkUiGsARvZGTse/F4wAN4d2P3R7nsVUz6litP4OD44WQiCzHigvurXMzhNSMxGD
JZl7J9JJtT3DfgKXFozFyWNCvh8MbJ4V918aehVRxOqyw1Juoz1UxL8ZPYqnONoQ
6wi0SP3+tx3ZN0kvAGWauihLkNI2T8YkncaRtWpusrs=
`protect END_PROTECTED
