`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
79Lz9cRe6Rig2oHhK+MUDrsBfP02OcJTP2wuAKL1lkwD07MOcJ6C5hQD5gDJ963B
qs0vk1sunigq77RniLyxxjAqOXrNIFfkFnQb98xZ46rfIF2irUK4cBUN/g2Hh80Z
8wyFgoA3gkaQS8CWxB7KWkJsVLYj+Ke4obPoxd9a2h0vYziMWrLHC75ty91UT60Y
OgdvFfPcVD/Yg0dHFZlMXbPEry4aAS2kW5bqfnP7XtJtj0j0AuloyqLMtwAsmiVh
sngZsdANA2wspv/jKqBlT0HF1mAVokMd8TVYOHLOYtRItRfA2gpYFgx2yibHmGdS
njh1iXmJz9h6yo2ShCf3Ox2O0z/xRNYJCF397PU3BURWYRxUMe/HA0A1SaJQP6Ar
HbKgjA9/I6pmGgCt9NIFUFR7F6XHgTho99F7Ln99wb5upIxryQXScqb2x3bH1Tyg
URxFuk9WWNsGkEKq1ViFESHk2AsE+6oh8l+c9bX+2wu2malZuoG8boSoEfJvin8z
lcBD0lpuk7FlfiQUYIv4Mq++zo4qnV8aYfVRiAVkoAqxVJSQG7jl5FoF2qZx2Ihl
weJHvQFNXqtSN43n16vwCVf1Fg1wHUQzyxgJzOWmWQXvtzOfO1vaI5Wemi0OULTE
yb+oxaf4YJzziBITYlt+7Z6bqfBSUHwYSiU2DUEfwi0P7X9Ue9H+oJsozmcNcnpY
OK47sLkTerZ9uigYrJQ6Wimbzdf8UeVB1KiGHKy+fmuY6fBtis8FEE4R5WQl59Yg
wPaad7NSzMSHf0SJZJmrF+3rCttIgxYE+ufv4qLJKlTzH3DVWL7N+9eb9LeerDqZ
gF2/qT8d8y2oDC82HNzWXRdhoShUrFz/RwERt1tUbLe/Yh1nWVZ6bJ1PyIJK5+4t
xKr4QowDZKTfnf/Xg7AFQ8Ou2qahdnR9TuG3z+CQu81Zf8PsGjUTCGSL+860RKiU
q1YX19lVC0ruPr5xtptc6FnbLbkFBCAwopbjKeWi0zY6iA+9bqCLbp68weXH+ryX
Mxkl5bMGVmIFKrDNyUmddBN7HiOaH2ytVXjpwVKUXg8fFd0OixLKYSVrG9xHS7dJ
/Vpeu+evXFy9ew+khS4bMxA8eJdBLoVYl/aZYeApZgaa4DMYorSGTFylXiS7Y0ua
GXNI2cThPrN1GEVPl9penHDwB1R1uqeJMTUOg02ZqHMH7mJoYZDei0gYvMMwD0Yt
Wf2s8KeY8fSaZmmDzc9Dz4LFnUHuAD5bwdjbb1CgQH3Y9CvaO3pDn5GDYJkiXUcD
xhijUuth3UFTI10crcM3Tv5WJ3gC8O6k+zEb1YsmMo5WS+V1L2fy6FMLYzCpt0Qb
p5J6tBoyGJw7D7xsovsCRLUqfPvSFhB0s25yQOTDUSvAAFLBzhTqzSO5WBMANsXs
lWqxUm3TB+SKKyBC6OZhPXiPk7k1jiGCcfEWTETN2uwfgcfOUXpqBqlAjLnKjuTJ
5jNdde0YVPO7bFABrTqm82cvuhG1WAhm6a1DGAdQJfv39sjqvvnO6AMwtSARURll
fHMt2oe7LrsRjdT1rcZ4Np3rmRh0I+3Rdn41HL+4szh26rF6PFJuq6Gv2wTeSFFT
rNIB27jPjmTRsM2qQQZv9cOQ4G+q3Ux7X3TeHj3VenDQU55qVibawlJtUMl2g6Wx
MCEpfWHULCaJpmy092VCLNSFO0rSClgiT1NKMqGiYQ49gG+y4n3ZtIzWBguk5f17
KaspAweXQJuXt3n+9Fs8RDV4arLS7QEw1uZcV9T8Y1STmDft7tQJtCyxsES6/j+K
G1Sfug2NQA3u9uctScrqegL6UNFCuomkmn4cHBRQAgJSWag/ZZwBfBIdDWCoJHrp
/eJ9vyrHPuNxJpahP8Ng0vf+wBtiAiam24gDKYKBD5o8cokGBozuYwYWEsowv+k/
idy0uzrXrXfBW90/jvI7wSdkwi7WCbHS4wtq66I2EdfbV9ZyBml2zFNVJT5CR3Ig
I9ah3gepehPzLzu8SLR3YG9N1YaUJ+c8fgNE+DeNfOSs4Z1mqxj3+Y24IAqyoMQF
+c77nwh1f+XZ3aNpDvrETHiokWIkPo/h13XM0ggLtdQuh92424KLFdkqouELu4m3
R422xDxdr6c//nvR4WuZx0nX9ic93422exlaUU36ycsxo+Jh/hb5vGKMTS0N9h/b
vXa7UJBAww+7HnhHhTbrp7j/0SI6MyvDB673l5E8wNqPT1RIwq9Zd0QFIyD/ETRE
CzeRCOS+X7L/jM4oX8hgkWikZth745Brqw19t/L0xLxeAIJ8zVRrBB8S+E6PiPXS
MqI3tey/U0v/FVfy7i1QYxhAVL1MT+BFDMz3otTd/bk1yQIzKek0/lePpJ9RLGj4
tB8Z8S5wI1yCw8pnisZu2kKamhRciFnxSeh7b8R58f4n6bSdpMkbjiBWAgFw7PZs
5iXqG5GxlSDHnu8daolUy4CdGiBAS+agV5CZ3kvVKsJ44S8q4MDdFQ/iPYgRR2qE
csLZC7yxDR4P4GzSWgKUiNkokOTqtIb929Hyeoxz8jR3PDh2avAuvsu+2MbBX01n
oM1kWbi1za81P4HrVRRPUN8gTU3Be0H8K/D4fMNzyzmyWNAvEw+ozKU9hgTIg9+V
+uxvWhZOO3waIMyyPvxiQLgIuK/ZGfxSLJ83ZpQry2dxIhagsmE2rY7soQyQZlhS
DXs/ulmQRIUEHQVHnwO/gh9aIyC/+6t99d4QhhcB0ykKwYVRb/XPLKMXtX70VKmk
VTPIadio1hdHtw7O0KX8U0dvmE0npUUjn4wcq6vB83j8RES+9bFUPOxNrM+i7TWy
4xKjWliUoBj/3wD3Bt7oQgxZJAKslhJYy5V+sy4jMdBcDyavNMNEzPqQEMVwqakT
TRSTaleFes1oV+xolQuNXbMSXXFWlUeluSyLIMIj1HQ9/dwpBMzJta0+AifwRI7z
EYFP4tKiU/7q4M9y9ZZ597/hAymXuKQB5INhbWAsHUbM+PO3NWBhwQ7ioe8Nx9aN
`protect END_PROTECTED
