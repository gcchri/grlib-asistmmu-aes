`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VZHpdNeUcZ9qHoTlbYDdMTMYFBgemfLaKmklU5nIUacDnRcTtM1VFTXCk6hl5Ti8
SMqqtac2naJhVSUJkc0DlKB+GuO3Hx4z0bOSQ5v3i0vd/+Vqy+54dX0FbKWT0bhL
lQHkykOigoQY8DhzonC2jqhN0g8szBwR5KcYUnZfMjUMw35PapxWC3MVEWCXLftY
xXzHmEiRsmtS5r4CdfHVoaIDCAdyVORYRE42oy2nnqH5O3pKwqwMqpMHuyqZMIgE
iYQuBI1s0cQpA11MADjrUNR1+OGRuY7unumeduUFi3G6WRtpRxPWFE1sNzIyJbqy
duMRBAlcKNH30dFuTR32btvQM9lnyA+FT6hvpRrIGSo8UNVzVPX5Vcjklab010K5
d2rb06SDPMP9L8UXO+6h9x/XFqGKfIvOVUiwy9KGIKMATECato1pubQdwn8hfU9y
K14VOzU76/xcyvuhp8sf9k/WREAZdAALGuxg5960iQf2hV/WHhGUU0A3sdNcbORQ
`protect END_PROTECTED
