`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x2GF+DiPHkmhbBJcTbE41gCiNbOXGDjvMHUeL781pAuDPzUoutBJr11G3RHgCB9K
xSNVb5MrlFjdu9AOauWuXmE+Rnd/YUm3UQaeRzkIFZnOUwC5X8oCCj46BYH87vVY
AF55zHQoxLSBpJ5H3XsxCCiQh+fxUG1qq3FU5rzoJlN6VqrS4GXrRuMtyxyKCWrV
dGHG6I/9g7YV77j7XT/xwJiB9hDbma5tnsGcPDmj+3Y2GDBVF8D6zfjMpcH5GJ+2
P8cYr8kA6wD8KUzghFji99auLI1gUEcJBJ8ky6Hp12hj6BKSSA1mWmh9Bp4HJy4Q
CsTptI1x/IrqPrYpQEb3UQmZiUrwE5cjV155CVgZc+jYcAnIEeRmVpXWCwBoG551
Rz8aKOO1mf8iGRO3g+iWFOCtvcN16KbFVfG0Jbh51tkPVmWByMf5FB52BwZr20r9
bxVYY6o5e0gueoiy/ONEtDXyNB+SNtx34NMw22Y441Hzq1rAEJc6bgu9Qgap78qL
SYi6C8litjP66BEH8aeLPKcC1+++sP9bZOy8Far/w9uBC9FZPRuU83mDdRCCR2kw
t1Ch/N9IMvwGrSOaC7iDJywW5aOqEDWT9JrIBo0NB1QV8UBZSPUxXV2rQAaiVY4T
TclzX/ry3iiTaU36R8XxSpe+OyArHFccOPt1XM41hxYE2aDh65rjtbJG3z7Arf+o
i8bbLQMzK+kskIjXF/kF/eymITv5dhxdm+uzOvajusO4jMO2jUD9Ly5a5W5eAe9I
bv2plBz2EhwjXLzW7RB8IF2YUlTNiZ5NYY+MgdQop7872495hanV1hrD9kv4LkBv
S46MD6dDl1KsjdCxHONg1qtoEZG7e9L/YFcp44ZcKGg8y9Li50kaDA4X2+ko+OJg
IdymeNBXr2/STdhp90/CwY2LLGp5gmPy+PIszxHfqx0h73eNsmYix8x4/I6mmEY3
yOZMhJBtyRoCG3aqGE7hr2yEFrtv98brQ1M5e+W4XzVFNkgm5MXahpMYtSDeJpZ9
KHUPSEwfmh5ccn29oeU44xBnnQP6yQZAvxDtQsGJTSlW5kZQXdO8+mF7VafLTh/T
jgjtyhDUIOXnmKB3sXVFDtZ8zZxN82/tmczTkDVQ2V7NKJfEsbfzIlnuZIuLwlWn
Uwz3dseqq5aRPYmmoAw86blGk6YxLVj33+acysn/GdvHhhzR4AIg+oLUdjScoDrj
8QubRmuLt3FKFobExPcy1qprQ+H7MWoZFMwWDDTr+e1VAxLMAft1FNHwExCfohMG
08BaRH9XvhVXEdlwGKbueWgNlYooIbTM5lcPxiaIaVa1MW0wlGXcmZsQUUcWpzS0
Seux3K9H+6JcCWqc8fZ0b+nePUL1BZiPnCKo6mWs9FOMXxOcIEtG8sLLsVCxb4lO
rtHBE+SIEpQ1CvohO8sNgwNcsR8ArHMMzn71dyo3a746f+Q31d1D2uq3oTRIEc0D
0ZYuUhNOc1010A/YWA5R9vKf+JA9pcWnZseAC4DMJ7XPBETa3aZ5bL2IwZSTiL3B
CpYaZY/ysSt4fI2fyMDNyXNuZJeWIFCtng0YopZUXiIrPEffxcL88kd7/G5+TGmv
xiqx4w7K2dTAeQx9mVEfuMwTiswXwMf4h3EpROhEfUw4o5s9gAt6qnNjzIHeqlfm
+s1Pi0MkcSSwopvVII156j1Gaxgngs1l2dyyCONGiHYVJB7SvZd+5OwsWbFoAt1e
RaOJbUnzE9qmACgS9uDfO88dnVEjOD0lYNGUfa+neHQ9hTiOlpHUFN8BWH6vAaAh
RO7e0cBLjpLCORFczixCD07tfCEZKx0w+W3aUeh5Cxs=
`protect END_PROTECTED
