`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G35FDQ1iCdkad6Goxx8RqlmoEOIYlu7N+sWeZfMMtHoUy9WORodyZeah6KDUyTy4
HZHqFvzaovK3f0iPLcIz4ZN+Dp1JPjUB+2sLuZiHJisco8sbHNAjigczhH6SYuNz
BkAlEd/2h2hhCZHzBlNIhpQHabxdcB45d3spsiymWATsW7g3kSPFvPKKaxl6G0kY
pBku9C4vh2YNiETJAf39TYb8YG7LouQP/GN/kCVK1Z2Ywy2bQXPcaojdaDRlY4mw
OBIgyf4kVAqMo8sLRT5qlhUonqY5GfElRhD4Ex6E/wzpzR2RgYir9ZN0Su6GwNma
CLIxFybBEiF5WpQvM/rcqztfP+sPrxDFIKDpKDgWfwNstLyqYir9Ao6lhsRMjsy+
/bhSD09J/MVvzCMieWbQVB2OeHueQZfCx8Cd/EB26+tSHvcrQvFXsr2Q9T/Z5k2y
r/2i2eUyEQ3bHoVN4gJuN6tfDqlCoDrw+UNdKnjqvDU+Eljm/BqtTX3YUfjvSk0r
C5F6llHLYZBwsEiF5gElHbSNHhi8sluTk8upswoBPQ+GG44aR0z8xKF2HVH6QmVN
p5jQItPC07rhQf9G4skcNQ2a7TGQpBzR6pO2bAzph8p3FGAN0pU70dbEpnfjQ4KZ
p3a7RGZ4cPMfvsGHnMqoYw6BGQwHQoLYfHAsoE0osf1SVxSRJj81Zxz7ZU6tUpbr
jmE0uvR0V66M/sd1CdmbzQ==
`protect END_PROTECTED
