`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4KPWx1yodej4LsP0pil0BRJ56J6KL/jNxF8oKhwwlp2/GhzqufZNOAOTfKb+3GK3
Kbg0iLlcdxs1pGj3q1WP81uXFNEiXDbOoi2VCa7zgD0PG4+Uh43yoXydj3I0bqMt
7Z4kCr4UGAVTkP/IRZFMCjU6q6jHFwDN+/PD509f11y7kosNbxlsnFYGXyRrsuqd
ThMHhsTu50OnW8x2tO60+CK7om+wBarkdNzj9IAHyuCgWAy72vcOkcvCujgfvHDZ
vl8fgX6UuY5ZUZhrNQxEd2D8X0DqwQjzSWpB0cqQ2+HIo1BdXQfq/Qpg+zQxdhGz
oqZVE1+pHaV5wRxyBwvHFbI5JyBaQUL6GfavNKO4TzZ2aAZ1nBexchKezGgbh2vX
ai0Y++13bV1tQYWcst/iCD1RH9+6YJaUJX4MaKlNuvESXf/jGroVHfElK3Ap2xXN
xK8x3BIK7M1AsD2ou5+pTRizAlQb6drLNWWkVprBz3t3zSWysJtSyj/OQkcij3a7
eHM7t1CDwMH6uYi4UMm2A6zznKxMwdu1WZ4yi+R1vD4E1aOyB8p6X/GQIaWfFPPD
4/rxu+PlerYpWkyOV5MQ8KJ7Tm5oY6T/0tSiWYGKE5CT/Yb4iyx91RBt9f3vYAOn
iQyYcjUMcCPdfoDsaX8qA/Ekw4qFo9ALrhDb/H9hTg6HWsVj5V6f6cvkyytzQCGW
1acNxGTfCIPMXFVmpsiO+ur7kITQs2bvNGde+rTi9O2ryTnF+2ufg5PKyJDT+fMQ
FzID1FruUT2pkhfMOHZD1Q==
`protect END_PROTECTED
