`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GD8nw1EVkIOQgi9VGtvfEjiGpsxLa0s1HLU0ogB3boaKzy0iq6UDk+KU3tq4FzA0
COcENPg9qJqjRVDVtAMw3f9YwqFaCTb3MzOnL+geiXU5Tl4nx2KiFmZhilAB/7bF
KQ7XzwAdb09LBDTpxqQ2mnMq0TGanHcLR4U5Ua7ZmPWLKjEJCIm3MTsVpxLv1Kut
GhfP1yMVoVPz91Mo1Md0Jk3sZtiRcGQ7EfqTv8y8Bh2ZPE5s3yb7mJeWaYU6hVAz
pNC02oVVUEEp9eHSawEwmBb5yYMksFJnODLJ2S+lUngbC31F/5jHXjWQS23ODzlv
3Q/lfxmB3lJS59e2eqvSz2X8XIVyCkI8+5OVXPhv/8E8dR1c40EsYbJm83hK84Lf
fRdKuUoKvej0zqdhH2fPh8yPiBUznJ15eJLA6Id7QDNlWwDosCrNzeFqrg4ufO+a
hAjpV1rS6O/KeEwUDTSwFa7FRqreLFxy3i3AhVPP6IK4o29Uh8B2wt6V5apxw8RZ
VHMnQCFMQ++wFYrrWE054O83hzTZNhpCQl5/Ev3ly+0c1cn7Vfaxbx/ZLb+N75F7
Ty5Aoxve7T4BhRW4Du3afw==
`protect END_PROTECTED
