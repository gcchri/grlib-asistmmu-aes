`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
33M6XiPJGqVZVoxtPAzEggyvJY0vRM5d7x/1NaUDnLJt1ROvX0BL/jCuIFzHVtWP
YPqt4KSc+qHsBptZsJIqiTnBM8Pyp3nSQoNbPHx5JVOLtfSnnTVAjmy9n4ka6iCx
5vV8V7e6+gVXtQaOV/zQRkJ20fgWT4nyuFAxAOJfNGuICEOrCUjIcuWMvPcWr07V
0k84LgjrxQJ+lKCVwlt0zew+NKkKjouoOGvy/MGmvpXpgSbd57NVODd1zxXtjlVU
kZHmNQQd9qPoiiG+8QB/y9cewoajG44b+UbYC0AEcW/5s+Bk2V+jrO983SOIZfV5
aqAW0Oa6M645OToK2CVELqtzUX7r8f+KBzyzGpYyLoPXu6tzHQA3JDchCFrCCjPV
MAyP62STiho/hM3+3+aPMo8EaDDRRIPXcsX+RhKuhqICKCrNnZ9XF6Vu172LyS4a
mkQLFLzVjAcJqv6wJBSK8pVmH+26sh7xLqzJhVxkwdWu4cgNPIN6Py22vISFgAbD
HG18jYMLzY3e/L/T0/F61zXRvvyDe4wPiPtF300BcNtK3oqBvSC/Fa2tO6WND5k+
A/+CXOZYGgpTJXAxdehHlTvbU2xQD/IqC/PTyHLgpNTe7buOPeNea3K6mWQX97zS
hvcm1Ed1732QtLRcdtXDCSxS1WkdEjkLqbYhEYQLNMZ0PPAFdpTmRocub7v1XEyc
l1+34FUZCoP/IG/SYOjebUl2gZ7Cki2BcUB/T1agsMiabE265leHnkIa8SgK7oKz
ttMAudog/lMUBHc26ajmyKAGBQrdOcGywkHQNwe+S7jh5Rtimucyk8oK/jz37IXs
htfq4KgZPl/7qZ8ntf9w2eorokj1gnOWtxXu5Sqi3GXXxrUmRDPDxiC7Ftx/gMDH
J/EsW+PJXXNtFdhMwNeZRhslhYQd4f9GTkUvRz0ro4JbP98nrKO9v5u5QR85EEeR
OKcVWQ7GdyGFNQro3DL4ldMZBijbfs6OEMzeEbD93WuHAx5jVDhxAW2OeLbuZgW6
ySaIwFfyv9Wr8o5h42AydOqwYeCCKHX0ul8VK4pGMajLIxd9X2AX2/5SfD/JwS+3
akv/X+DZ03Mc7P6HDkla1wkObBFwcmFHbo0fLqaGYy/4f6KrIwR82x0BN7zslNNL
mULpfxtku07YZkqUJd+f6uY3jFziOQtKl+9xVLMmZ96YfqxsQmKA9uhTccXQTs+W
wc3w/ioBDr+P4YifwsT0VvLiGqbCKwzpMlF+bZWc8AfOaClp/gpMa/4F9pt/yCWU
xSJzqgZuzJl7L5k+JC1QzFrYMaY5/C3O8zf+lqhY+vCVvK8b/Uf5GguWnjUaQsFV
h0V7lXvCu2VKv10sVi2HLmsoiugUwea82VgBYw0rmdPM5ZwxoenZC1BY+cj+4eG9
mGBrniEWk1AqlFXjw7H8KagMm0y3rRWZa9TPcGi8VcnY+rV5bSSuTzoRu+hB7u5b
5792Oe5FfAcvxjf6NtNxXt2RuIudojPbg+04GY3J8iqiuo/xxiTey3sbQPBWTUzC
1iAH3RV+RSjf7Rf9j60l6ca9oVGA6VAgEPPhhDAFPQhjVzdtPF2uYr1inRoUW19m
wuQf0Wv7Z5XHNODRU/auk3GLBYTZ5XicB5RtucjNXMb6RXKZxb2m1bT8a3CxURpN
2r/zj08MbzNgdQ4/sIFc4LwtY5TdiCVA0UhkRkJTVEOexo9AccLyRTdI8B3kazF2
npYlidcgkWXdym7E1NOuz9KbnLwQlpbIPVBvq7Fea86fgpSk6nKUAB/oc/hfbv/F
WevdViRJOtTk2WddouWx9aneIBDMyf7QY4CHHsRkrunE1WNUzVLSwbKNOuXtOX2A
mEJxKiQXwT9VZ4GXwfr6sfLKX7RvvE4nyJbImu0scqZv92ksj1wRdqodsLZ9nQuq
JHkv5LZU8wB7Z1DvTurkkVrjuUdaDS78rrd2sGNEAWqfJubspJscQ5R+AFEkpLGM
+MBEK9SNxcsgr/CQH3FqzOD704zk29JY/rcpMHR5rnUqTJnCQ9Cb+p/ZbQ5ojBdT
iK1KCTs/mE9bklwlBO0FET6fgBdf7HaYDoQCfayJZ1opD4KmwgNQ/ApfWaZ2Na5h
ndmOMF8cJSBw3d+Zbe09yz5+jqdJaiIVOG2wQC+iYRHY729tDwcOK/CGWu3We6C/
fUhgmMOym3maB9pqmHIYjoW1+ktusS1btWtVQuimbHTgGwVbFREKZHn+DgjaHlNj
c0T6kv6KN4auaP/S94pBgaeEs+xvNrI1varmAV42WkQd7W1BeVLe0mTRY9wCs8ih
l2y811juEk9T0J4Vas6KrTd/glYHFUWvixOYzvR9zWs/6Fnqes5aGhtIg/ysU6KV
X3bpDReHKbaB3lRNbVPBgme38IkeXXYwS7GRxnqx2phvcPmvZlHNDM5imnZ+pCg4
PS0VseMFnt4rHVdcFWtq62yN2vIqGsaK0LifAPBCmmNOtEKX9kUA9bxMe9muEBxe
BH2quOdJrW6m9frCG3dTEISWxk1R7A3vVo44KcRMprGBItQpqWB8HjeGCrI6TBf4
lndpyDh/UP8nGkO8p2JEo6SDdReZY6vaheCmCCQPls3JrHeq117Qjx+annz97GXF
jr/CJGslmtipKI0f4hA86uBRW1x1lLbNXEi+c6vStyapsriAyBkkMNwbHsLS0gMd
zrZoKM5JV0kKaD0wQM/3wVx0l0jJERV53uLcUZ3l0pMMh45w7+uaEDmMRBW1l37S
3bSTzQ1fTzhZsRVVEtBdR1N348C5OYQt5KMqoFnFVH73bfHm2PRLK6AmYSIFbGb4
3W05rnWNtC7Q+yk4VUIi0fFKzYbc1mIq352F0FJoEhYVINqzWPBfDCGlwvcjzXHz
+F7NtnLSKBWgV50iRDPaPYSOCEKv/p1tHa6rrJJLv1KmxeiYdTeuewNRDrUT3Ny+
kQR5n6ttIGiN1s+SZImNhB9ufgDaAq8OXHVF0x30Q8t1VwjHs/UX0+4ylQKKqsGA
HoU1AwlOpeMijcLALHpUoi5GYgCU1MCux7sKar5ndcjRVRBqul0Ovm2mPDjq4gV4
l0y35bqq5/vyQiDZs386ZW33Y07M7Fidjorx6zLzPMv08aKrAe+seMulwhkgJcVn
gD0YFvh8QPvoF6/QwlDcWBCGCNz8wLcJ+eVTJBCc/kCjdRGoFk/IGs94k5bsJISC
0ccIirx4PBEnAqcQVkpFiqXYzEaPZ5NvkQjwjA/jSR34L9PdpX/1JrnF+1oCUt1S
gwrqEzJq2KJz24yCdln7xph40eAVW9GSSN500JWrBYWT+xgDXLnE1kcR0OqMCB80
EeISXrbrb7VLZNreS0xgKwUr3Mb1SXolb5mZjx0aIlhBh67vu0d7Fcn+rtjKXer9
3/rl6Mw7K7PqCGkihQvxFJ+LJ/vjJ5bgE6t2yxydBLXraxNQCCZaWZfitNJ8byKe
abtZ/lW/c4ZqHW+l/y10UGhSohk5HzVADqLnqi9PUx/p9vufRR/vxcMCljPlInJq
Q2V2Jh2HM92fxoj1JF2QPTsd2QDkrMWnCMKIgTikKuiO03d+g47OZ2NtgNYjufSV
FERpx+Q0e/Dh2nTcytZ1UbBpdGHTnGo+WSDCmfCj7oHoYlCGT8xXM6cLiZu9dUu9
CqOiZUniwo9eSPOw6nOrEJ5wFNv3XctA7B3/SpBH2xg10plQDm6E6jindV0enyGn
DIL52W1NQAhtZ4fAEjcS7aga2rYrSVSaozjbq8hQgRSV7/8TlsMiXAL5hl1Ws8y1
XtklqcqvPDK/H965xD4Dyz8VqDLNTCafzJ/hBageKPdRjXYxd0bHnNuqgRF0iPBr
Ke/Lt203Se+KeT82RV3yT6BUxbpQ4dAtFSR5P40MjahRq8A3Cg4851JsEV4E6BQG
OkRhV/V0mUl5YNexC0bK1BNOfBwPLOjw4fxNJNjRdO1lOYyd5cKaDrE1zPuLXrxM
0A7tqjs6c2bNcQS39V+fkgty/cXpXlZA7RswU8BkGaMC5wCpoHfSXoUaO9vHpMdX
N6HSsElD180FNDuKQlWVO1Nv1C/x1HM0dtpx9r5nauwbsXzQ+CsMPbqCrTLX+pIo
+0ozngiKYxk2zJHDBjnwVUQAnKamjAooNYOk2BpRepUCTmqRXHWc/zKx4fALdgO/
cN5aRZ6ZDNklHhLBsdNtBauVyteMlWE5U7ObmFtDaCjmevEXSA6Y11VMDYFocG64
wWfav6HN0jR06XwXYBpriovnogCloz6u33ORovdfH7X6rLZXkLrhvPi8kaqdIPB3
Noir0GohqI85cSjsk2/8j5xRyiYIg51cQ2Hx5hLqYTNtF/roIAheitXrO23er+Ig
qkh+y7HRXeay66e4kAFd4JEDDzKNz6fFea+gACxGHOONakTWrmZToQStzlA6m/qD
x/tIclRiAE0bUQPwPkDJ8v6ZRNKgS5WwYVAR6thteUtfw0L2tAZRMVtyMiz4H+zy
0piwyD7s8dM6Rptvm9/H1TO+I/X4ez0CpsphlEIE0/VIA2JU+FPhXszZU/cQy4PR
uqD/N22ZxRjOGofm/bxjqCGN1qtXKG/j0m3dHegPrWVoVVJunYDQf0A121rA5iay
vL1pcJ5EARQZrNJUHjM0irAkRZza7Cc3/0ZLX83x7J0C8WY1FqDHKpLg17C+aK6E
wmyzCn8rd9NJFlIvS6xChP5QeVcN6YFL9+ZbEqU8Ug4HpOxUEd4oPVvVC6USX8GZ
qsn5IPalBhgi0Qo7Cj8nJg7GNfWRexO1ZCoQdMNnAkty2Ioxrw1/+wameqyZL6Vi
0okr0nGpLUvyo+niNS1m4OvFnYm/jPphLQ4vIJ9h9KMPPRw/QEht1RPseDxYBxby
9BkJ5jU0i+wPOLvSqoAS7o0NYM4/DCXTkKp/rN5mEkEbvJprtJNz9lx8seX3+xmU
tUE6iv52k6+T+r8RlQdBBhbnD4j65xD+tUUPsBs0rK+J/pR9UPGi3Y/yr9KZn9cO
p2pKOZnEnnF/CKKCOxEJ6reqgoxsnU+zx7B8gyg+i1MsaBi7O1CBdNQIaK0rfmLa
s7QchXQdwoyS0o9DS+uX5xNMqLouBc6uoyQXq5PTgrEWAJrqUekWRIzXqsR6Bkk4
//BMLfukfccMWahLNJTZTcoZtOppHBOJm1IpVMR3dis9x+6v2k3dWaF6XMQiaLnT
d1RDH5nLgwLkBrHw3x31NYboUkWl5pYJi82OChpi39AvAakrDFD5ndanuwUFQvJ8
jmYObOPUvWWetQDuudnNbnTWcHfJ6g4fnqEfhq9d+Vpa80MbpAXwKl6iwDIzRfzS
+QiT3JWg/d4Vg/Evp5W3+1uAnAzwIpunSLZIpiWXnMnW8HQcyKONqW0K1DrVBOOI
YLKUujFI590LJUwI2wcIklZma94ovYAhGa9KxSQ7qpLdlDHLVBulNQ3Uqn70J7vR
rcEr/Pb4HcCRe1aJet4ioZTBRnec41+33DSEO1722RP7GoLVnsNvqbg1DGk9l7yS
g/FGCOBx+3//NMCgZ4aJTJXoMkzOoQYfcWBuT4m9zXOK4MqOradI/JmeB/Uk96//
z6mloysgSbzJvf80cyPyLiUuWGMk7nnrCxZnU3iZnFjonpdTOpGKMeXpphvp3OQF
exEWr+IKWlpKXiG2fXNZrvkT6JvjIfmEtqH3rTxf2YamRx2IhpSXpX/Tn4qTSUxZ
3m7jvJXCDTKOo0sP2bOHQ4CYwBXVIYIimYHbejLl06WazVFw5lPspGRWCWfY3qPc
V3MEKoVFy/5GC5m+D8es0qJiwqApofI/cgEBSKxnMVfIwmbWnH9/bbHayYCnr1qt
AfvjZyuJzXWPfL+3kKA8aQ65p+/mKMP5aoI3UnNZ3ENY652NAci2COA+CXjaA+vr
ln5qUTCHRReGy206kGT1yoJzuBgctn129QAVVwP8YIdzBB26ExhSk5B6GEbx7jJ2
Elub3Cxe8s51iRCT3TGyFi4rYLR4n0QlMpBlxZmvmdnumvGZqdLwcqTnEQnvVuMc
vRfeWtq2UziGXKMxAbRCTtmLNvKFv5AutrdloLRIkjcZ8ZPEJgCYRdw7As8fVYUw
STVDyDpndUVRX/nTuplCVWVi6JgBtnrHkczlpXSGq0g8kUeHCRbmBRqD4jnyI4Fa
AdMzm71IeelS2C7b3Y40F2g7+uYFxgOhSHrnoHQlvLpFHaL6Jat0iPgvpgjBJHo5
NcsKeFj724IfTrp5roHsyHB+cEsmSqyL8tEcGApHhbHAcCkjLL6PVH/wXeKpahb9
5AfmdTKGAt9ZyRjiZa4DG76jxJ50kQWnrGFLZbt96lB4MzbajGnBT8hBx9TPz5qq
z/eylX0j+RFMER82HWAkE/BFV5ahJRbRiSXkYJ7oWfixcYiOwrlM4Pb90cjP8pox
DdZOQ8o7M5JOwRTyWPc9OREcJi35JyxAw9r+2E8EKesvV7nLl1marz7qLuiBJFFL
jvSKNKATQgiaQo4oRkw1SFXyh8BenimL+d3R98QLZmQfzaEJQuf67D5Nbil2annK
hrZhtQ6rgIEKu8wKeuXi/qv7Dmx1rjgfAW/9fo1/GDMRKrzzKL4uQDPZevO36GQd
RrplWw8UoghcOroKbs974IAtqT5EIFDziHV8JrQUpVaEgGCtJqjBXsb6vFxmRhpj
g5jPCsnJs/6IcUPScAWjrPPYkawDkHuwkFRLCnINfiN+KWSGssSRIgR/5dAJukii
8mTIxHqpHyXYq99oa1vN8bhY39S2QH/v48afVG3JmxqO0JLJgFAdrVO/HJQbolAS
qVO9I5LaZii5Nxl4cfd9IH2Zyj+3LbggReRef/I8LjGrUfEj0frSsXnqLY/Tnnat
TczomDEFkduzE7XoQhZ6wiQGo8Ry2wBffqyeavYaAlcGnGMBxUNhY91kpBHJQld8
o4oJDbjSXvTcMUu/KObXZnjI22YAEsrxmfAKa5LN2ks8uupw/7fMzXRJnBpkHdM8
4EwvtVGSKU4b30Fx7/sjMdwYlZ5t0+6XlJ5qHeo3f27flx7ihi/7GWQUMkDFXFaD
iwYU/lwRNr7nptUtSPfM6VWYA1y+XAzSnTpmLqrjxXpaox8Z7+se2TpOWXIKlbJk
3Rwr+dWUEPdH5y7zvrzcGzA45x7Q39KDob12ISotplYOWS1AlsVG+IeyzqFKAqEz
Te4gCYLGzuuu8Yo1uhmCIPZXrVyPIdyXf89dJWcGXMvNJw4y3yjHPit1v+2sRSbZ
ivzDgXJHiL1Eso69hBN6rbdwgHI6/HtDfKHBey/E7Vq95OsLgZQt5bJ/hsnP7RhX
9GhwvO46Brf1UD2KgWJAJ0+NNIyM+4hLOWNAa1QCB/cVBcMVPr+8SsK3C0bR3u3X
CEXFwVNzSw32JQTinBQu+n+HdStfma6oXwAG90lThVWrm/72DitMGF96M7EvS5Ix
NlIMvHnLq+WoTEJy4w9vvNksowdgtaRMhkJgUOMdQjAYxiLVSzPSNJ+lTA6rmIFF
WwItj0Lk1NfWpeA93o720OnYUxX1ZexE+upMrJ7UBss7gq4EEQae9gDvSGyCVRWm
5y6Q+EHw37Z3sajSJ2Su7J8CquB9Na7hBKoWzoX94RBFJmqRKA1BiyszbpTAW+at
XUwOxE/Mpwy+QomNbGXZltFE+onx5mTnEdp8LTbLMksgneTvi3s2a6SqJN8ru1e+
yxM/hwPHC1Gb857QW9SiZiXKwfoIpv9smzjXKd7wscOHfZAHNU/9+hpksI6POk7A
AjGcEUq1oSu+TUoE3mQ0Av94g0x5DX8Rrj91I/8cr8CcyScv/yRrGt6nL0V4V0Wb
xBSz8C/eHDZ0YVhM6OEzZz+9RZph/U3SkZXdBOHK3diJE/J8AK65OPMJPTDgG9ME
5+aFCsJOKpilX3PSQB9eYmD1PJWP0Gph0F8qumWEIem8157GVPqjjR0AV52FQGOV
UuholISHDWZ/XU41vSI9EAStUv8wWzEGAezJUZZ2E4Dn2n2CTUpnovvuB+tWO5NP
2E1n2iQgXyobLjN1ckgKsS+DlpoUvPSYG7Rhv4ZYIsZZ1zuemG4wB9B8h3PBB0jl
uVlbRV1+1/9JCGXwyKSPxIvVxHlPzB+pD+GJ9Sg3yQmEwzctnfW5UFxXN5/hoRIg
aySmCK07OJOF0cqEW8kNfNCkM48fyW29kkFRGr55DacBohNZzli9P5sXJQf9oDuc
E+2T1u9xPV65pbUvPyb99diF2z85hwValoH1Aige/06nlTMGU9oWikx0EORK62lv
tb60fgszhZKnbfeZBBXyGATc2lhIbKHPXdyYThkCHpC7lovX9q68JvAgLnEEAoTZ
NmQ5f0/3elvv4K097nNcBkoDAC1npwZPkNNolFtBgtiHnxla6mCQlyMWSTUyTtAl
Wm/FWMazIyR63wOheczhelk75pXwPpOkuL/rgJNpAiejBR6BDKxtGsof6kqDJaKU
Jd2kMm7BZaRnpo9Zq8J9yqlTWvgyACtHkRCAo+lsQNyY5hs/7j+fg4HpuBS3ptDZ
jGtBrgQGU6WVzH6+QZDyIC9q3ZWVyfwkyw3pSbhJ1p4pNTWcuHdk5ugAbqMV5G15
GveqriqeopxnPpgPRtO6wv2p3I6hPpKQLhpsHAFaISc3vA7u+ORMKWQHf9fUHu59
BuQpWZC3HZtBypraNpny7yQE6C9C0FQb2wMI5kZ7CtZ/82NrkHEQPZYJ0Mffi2w9
vkRUHlfaksjD6vGL2l+T63Vaffh1SAiFtJ1w04KfvoAADv6Z+K2tOM/RdSB/i4S7
lfVJ8rrGoOPqcfa7eNH5rOWJFiTn+q+uyqCMkaAT4pGFAz6z1XZqCgPlt2sPk+h0
4mMoXXghBA/+PrYnzfFR39Npdav2dzych49ANIdoWgwy1WDICELOScBoh0zcpZ+C
aNIaTHjTX72OO1tDY4m2EVDXpjnaQeCREKtFeiSEkBmSW9xIYMxJfaJKQAw+pxLA
cX4ukWTcdvtZ8In4KL4Nk+Kd6yeQYKVXVxv8YPR8+gA+YS/PkfJ+qWy9USKY+TQi
xf5DebXmUd7hRqkXxvHTituBQUNfsZ6wvRzQwSUE/66JCRTLfW7H9xxYa1aIV1fc
yGwqyf8ucvzlGBfsirvUgmCpyXkW4hNP8W2LMUd8zA57BkE/2TJjqYVNUGiLArz5
14yyLaH/u3H+1wI8/IO+Gz1PDlKVtcXkygYas+l1gz2WSit3B/hsLjNoxdRJIQ3+
FDRAs/RV6JLsyou1MJp7etiBH4/raXyfE15yo2HLiC5RRu3w6cwERnCF8UMiN5Xm
9RxWJviZBBnsf/vHqVS0k+lxtKOmumWcCf5vxNGYlETsSi17aGp9jVrnan6DlVSO
GVl/3LCae2vYgS2u9YJfSCURVGmxnNa+U920CTR2qvT8Uhcjfpn3rKlVC9f/zHmG
wsXctHY27E1gRCCLmkeF364h+8oRJCbtcKli3vVG5vibUc8Fc/VbTs5KOM7DXIVn
/0It9y54uh374b+JqEglTLY66+ZH4XSPp7EJTFYQ+62LbVHY2qSY09t10TFUa6rQ
kkSgInG3/KF/M0o87XP/Qv4HXhMu791Mfa/C0UvM9zN/SVYI9821Ub8duXaESjf0
GraCk+by8hNRSoxV2Wjt8yHyxLpB85F3WIs03d5za76JDM0KXbg0M66Iz+OsuGwD
ycFIc87p3AEiATvZcIKrACVmIN62AJYdCsQIdkAcLKZ0nx1cybkr3etfNO3LVkdz
y3dtezjt32Ud0hpDCO9vVEfmYdOM70b8BLQtdH/UTsp2jhpdspcS38B6M+V8nYgG
OIxiK3aSKkY8QsL8KGivF/31OKMm0utvgah6tW8BjqHsCDRA9tVOoVNgzJ3WxQZJ
N+VrspUIFaIwEQtupn54sTtr8uHQLszFeSiq/CHcq3DfSEy67Qve6TzoNlkYHtMi
KRVgtFgQ9iCZjPpG3OC06Mg7N25lQHyqHtusrY37RSMioCjsn3TcwXRL8oepjpHM
XcLLLcLCSRE+SqsO0V/IKMoXKQnmM9p0If09QfKZeb7PiIcsIAKigoGPfLQI2YtL
EnIWZuXOePKjJ8fzUn0c0zPbyAcyY2QGgfoSItLMAvGGM+H4Cum/8RT+AaWnd8+o
JKm4qoegfr4ounVksZ+BjOWc/LvTvll5AtBRUClbouPdb+668UJZ5DSioetOfQRF
UbYi3og4Sb/YnSV8X1UAmdDqPKrbpHKGxH5xCSTgkWRpDZGwRjVftIVicN1AhBtS
t1KBCt/UCNOInhjdGttEQT9LbwySmkT4/YZCDJ68m6nLHkWB6IUdxLhkKdX/43kM
UAdPRGqNez4Ektq7FjftrFdMaWd3FPYhvycOm2/bcgrtkOLERiIpjOGMpdTSVo2O
iq8Tevfqhhac7Up9+ANckl8MJ8f0SDdcLPDPMcZvwSvY05c0EEQLI30ew0L8D2yY
KOpufhyjxeceVtgfxMo05fiWQlZqusJQOYWrmcDs/xy0Y6v6tpdk27Isd1iYEwtU
xj8N77qv9gQ0wfNWCxEOt9fRRCkWATAAxLxEu+i2CSOlPxt6Ot2PXJJK4+C7L1P0
N49GVIatfvwJB/DBotEpbmeOA8bxt1kcpAKW1xGg8bAJmz1Oox1E3sgd3geUh+k9
FwuKNi7WZWSV3Pbq4q0LLCm7usbqM9Y7zh46eeWeC7J6IH+u+dXPjUc5rLyl1ARy
A0IMLsL2WYVXTqpn/acdtrYlD3M8irlby+EPsTTmqrLFyJkx+RaH4I9dnjB0jDih
fZuh/rdTj6I5izzzq1aFV6joGAu7V/g6UBpFNnuuiJsjs3Yzvu1WGKonmaE0H70b
AXG8eGgJ14J/qzChEJwYN1eyNYE7HrY9tFXBV0WvH20gmGuHz7lU42OjVyuwptkU
47YGcvb+LRuqB9wlNi+86wtRIp16MrF5SCQAcj7g14JdtoLVWDfy0EbpNJ2V/pcr
BNA2yVQqNcY5nlRBjv5VNQlivFt8mr7ZB2EnoiEKh6I5GWmKFx1efILmFwfVqdSd
rwNTv/U67OQ+HikgO3sLYcZ0L/T4+Krfane4mclM4tGceqTCldJNsX3xIf9ykeVY
dECYk0RpYB4+JniZxbIxcrekK+wobHuHmi5QfZ7Jq4EM1TbHEyxBQXWTgtepiQMN
u32OpQqJ4lWG1GMoBCbBq7/pmbDHFFfwVrPRuRKHr8wiisNSeR6Ph9hFxNFS5wbL
YQ4iak8LCFoTDU2/+lAm1D0qn5NuWoQAXLN6rcpTPZa3p6zXP3TDlEGItWt4hrSm
wEhSSUIaWK0tgjLXKftlDLADIZRk74FOyjnxEgk/8M9anlXwIgVP8eH9/8GafgO9
y9J9+bunY6+oOLYvSHzGxB+e2maHAcTmUmMN5TMM+pfNsntwmSiZq+Yd8yJkTFz6
KgrLNY4Z2Z36heCF0DIZqVdsSRzvW0BHUEa4ZywjzBtptltpQaHII65BvH5RaUal
O47e3kDb03Kl92oM5WRs+fVWYHkpVW3lYb/eM9rAK6ovsT89d74gnBz0h4Vlqw9O
f58ByGL4fYsnJV+He9CIF0IbPQ6IgMfu2zIR0jdwpBeI6+I+7ID1TcAH5mmvU30r
8nprhaBSB9yMHUyXdYpqcGxzBwIAYRVMqIrMol4Ze6EYGXtUzq7ANSuUF9cknjGq
93sztmn+TCRJHZelsbJe7ZmdV8BKGTC89prPtiJla9XnwcORgh0AobzcBN3Jtcfr
+MaTVYtCG2ZbkyssWxFwToCIHiBnqNN++Td7WspcblcS5eUta8otIGk5Eh5iZmeG
GB6dVX4VzoDht3/Xw4GOs0KzZO+FeBbIENQDOZZcP26PdCZJ5Loqg8woCHA0qbKF
YoL+FKebxib/+2PE3/sGakIsXRyxG4FyF2CfxtPO43R1p3hv/3yTp/7yLugf7pzj
gIqzK93W90wTrirx+Cmzg4r8gXONAaZw2j6UqkKuQhY6/a9TnnDtS6Eq16ur+boL
la63HQQZsR58T/fi/J1gAjw/ZkO00704PZbWuChYHdWxoT6b0KXPhmZkough+mqs
wfL747YqXpTBiNaX4U9tI5cjMgCLuT+vcnr8rW3VvKmD4L5UYDffgD0a5C3+Q/k0
V6suTYXCUkcaV0pUXRxFCEFXlynjTmtsvUfXYoNKqWGtkOxf3MqIqemgqiggaUy7
0vdeLJyxUU9FzYUw/8KI3f+XHgqOcGxxqPdq6TJndJz6mIm6fy7xxLqSVrjp5eMc
X8W3lS1kAY5geAA+rqI2/Z0cqvpuPsxwiMkPm/Mhi8fHYu2Awm9qDvHj2jtFsCyN
pGN3jQtGtk3gwyP9LR8rKbHnCyTz7Iajmp82Fo+uE1mQNDVNslLDVVmj2nVpg/2K
g0B15FW/+JTccE3YM65rVZAEWEOfWpF5AdsUhAKkFKg//LZvRpKweIgkUrGHhQyz
aYjzujrNajtPd5qptd5qco37ADztFOAPx9k+tsCKPHNlU+UDNYkFH7QU5pKeHbyp
53aVZ9JEEGe33SkfhTgZZrzpz9HIggLpbNs/xJX4r5gD+xh1MSElKZljhqYPB6z9
LoYzlMQXZhZkmN6cMbnkucb4sRX8Dge0Ccp3Ey5NQ/sEfiiYKHuWUGoqpK7MVoAz
puZRmtorXcLtErJ7k87IKCRcO3D0RK/LL4PNaHB1kmoOUeEdznh8WvxV0MCvb6m1
N6ou+wyD14naKQZbOUIKfU5mvVW7tvR6OB16RyhuWoLma/8D5LR5E3zInYUfK7nx
hXKP91enbz+US35suH7nxr0yJ6tUL6EPzEQz2ZryvWN2N+2VAyYbIX50ZHE9A8YX
PU+vFxixihK/pYSAYzdNI9VbdPT7g1fz2hz3uBMEJxdXC+2XyZE12lpWt94jJBdj
WNQR4tdIBAsdRvk/dMBQEKv9DHvuwSgDPKQ71/nO4CrgpuU03YGJnooPbHjmQoTG
3v9618gvFhz6DUupLEjWY+MgCksBG2srySqtnz1Ltn+jScDPxWSVOpvjjkvuPyMM
hIoyNLfuzaOzVpkfvMvEQBU+7pn9Y1ewEvZu/h5ztaQtRWw2jIbeYUERK+zlcjco
X3mzCf1LaFX0duBWAqB0NGEP7BsKpcQbtM1HWVv222LrEEwIleFLMpSv422/IBQg
5yvre1Nqmb8kSpQPe9ou/4aPo+RQ2xb55OZTA0AP/E+ayxzl2jDj7H7cs4OiPs3Q
cpZDzrlKU5HSIKQMhcwi1JZJ88NNviEi7pWLTZ8ropDqC5cmroB3Hjpl9oy93RBZ
VCMZ4+832FhbiK9UiRmP/cewWfTyWWI6Ny03ED+v8yQU/orFYHSiwkV/wyuN+jFl
dIKdNUAJRwZPiYTA93uIKtAuYARKK4KRS6qxjmmDMiqDLJncsVdHa+e8pbMsbYjQ
WUoRNiDiFOuOIOmZov+zH1HvyWpphu9ZEJK5LkVrxShGT6MvuwqRW6d8Y8u61clR
JFjFlhQspNa3S65IiOULuxj4VfOEDspoo4+7ickVHvR4p2oVJk2R2Dq9cTxUGhYt
8mtISNrHGjWJTicTynp90PABg/+Q8w7EbzEY/2aFKxPzzmBSgThPVVg5kIiPJ9xK
EDFky1zFrog0hZ+KKomfliQtbzp9e2oL4BlcgGzabd89tbpZmGsf8FhdVhDPgS84
24KWKz5zBLucltDE/VNOruZlQW7AVQwWHvPzG/hRSg+guL3jCPdpZ4mPGDXQ7Z7G
nhA2T1cp8UIlQG9lGT/MiuBEg0TwntXxlQstsxF16HtmG/OrN8eIO0steMTRtFgC
gsIF73OlmXjfWu1kwy6VJRwTw3rpVTps1FOfzalQglmVjFLPS9lNbAMnURjHl9WY
/Ml0Bk0Jm8UzduOKMKZjGZMgRuiKUK7X5K7J2JkA3dsAZPzp4RMyaZywvbG3KUy/
w6T/jbFgn8DrOLSULHm+EzTkkZLpgykRjdkNqyuDccjGXWkdTrXr4Y/9q+mgx7IY
7KOB+Xe9okIshZJAH3rxptR+19/4n7ADDSLU2q+x2yEc9mY064J+D32Ka+9jG1ES
CsbfsJWFOKa9BXMhLR2HGDiqCRNIAS1k8bbJH/c4ne77tsgUHUaMViJwzFp6cIOi
ZhM4BwKPFHxNh/Cbkv93DKO3Ot3GRO78d3alEfAvrk5axJ8PtRflzpkc4K+p4exs
K/QxlDe6QHdphZ5jOgefZ+B+/VztBvgRIxGnx1ZglhWc3o2plEC3RaDQoDcWPH4I
+x0lkRczuc/B+rBYYVz37OQEWtwEbtgIKlL9lRkTTTwdUhTA85h9hroTiOuUwIz7
zebrvksS5sVOs8CDwv/6u86/J8NGp1A4hV405SJxpX/w1QfKE8tvbiWZnjtQ2mMS
KglUxm2jJoiDCGtmySmaH1X+Ey6w3P+Ek6VUxibwJIfQExIvpEBp0jhlmUVb1778
qBwcn90b+pQt93JguTyMpufJ/MMKpxsFjsuVBceL2xAATiJ5FacdZDXRDtkUiku8
AKPwaLqkqKtqFkWUfYM9MtGsKD/C16rP2nLHG3NqNGQQZNTZBHn21uSiy1Z6UnUE
ElAIp69ja/6HzkBg/UqnxHG0mox51pfqJwJcB3VTdF1515xpwMZNxE6Dh9iqI1tg
3T2AXYieeWVpsoPob3AcZn7dK21KEQ/NA7FBKrrf8QPIkGn3ANxaNo+jRyplqoUw
Swps/smZ7oUs8HQq8RSisCEfdACr1IsfAEIJ30lq/1db6U7UvHhzBwp5MT5oZxo9
1bhbX5rR7t+2+QNItAAlFfFRSvxp5qqygBkVHzE8SLokCsjU4qaHsEBEvhgQnzsr
Q4w4Cd0l/Rxd76WWY8OG7OgUeGcqlhR35IulWTGRxlv+3YGxoHTYwhmzjy7UlQ2P
aYM+hipU/YPWx/jOBx5amZP77nTPeIZ6uPSj3ocL1yHQgoYfYK3JvuKYPnsx04/W
3qmMrLbTqScVXrt6t1XIxMfKkLYsOG5PeeXAKTZbSA8JsDbxxEfWay/NSCm2ulGn
RSRq4MZjV9O+ItCxin7Zr/z8WrXuAnskG38SxLFcn9ZcfW5JanNdUcLu2/aSOwPK
CL2bXrbovbQdgb9PDJzF0ImD6vRiXmmnecNqaYVc8CknQZ78pnw6VP5YWxFr126q
tCNLmckZa1gqnM3Vw+QRt9NtrYKX3HHZmGHe1Q4aZYfuMAhcbEv4yHmeYTin6tcS
TENeJVuEMTwSJWSnBckVTkhTTNXSwIPSak5aIE644GmKLmXPOkJFytzi9qJXKYuB
QGv8wVOGmIVLkaAFGTUG9m8oEQ4zcYVbX/MdHKaBN9EKW6nCsopGXHkGiuda1Oa9
5GHAhe6K2c8J/3eDvvphxjlYAElOlMiVhsaEXK7ZUxjePm0AB8we21yt43tV8OWB
5e+rsOY/MULjxbu8gnDIR8nKBw0nYBC+nkZ+J2ojuD8ZUCfTKoNgtceB2OJ2wpbv
M7+7z+Y5K2TFXBH0sIBX+9emw15cb6P1ljM4TWDDKLBqYptJjlr9SJJ0DlItkOCl
cfdr1LV8upgzrPNodu/klIs7nl6+ooRHtLVbfXQU5n7jrMyBPE1G8qmeO4P/B1xB
f94bTfn3NsRJ4Wk9MWa4LOk3XlwkP7iqRyJ9fZFVyJ9KlBTHl4J/o8hcTyHX4P3e
aA0uRbezs/bqkFd9EAGE14OM5mV2I+hIJPujvAv2EZKQPRCEnyevw8+gQQAQ3zU7
w+7AxcMmpKre8/rn4TplgBIxGVms6sy/yZIqjL7qCRfseeueNJa0Kc2naFSSnLX+
LegqED89fan8qkL1tGZHLLKbBkOZWouGSVNTl2L+ObB/A20b7i9RAww1bkhvKs9V
iBhCLlI/HliV6FxN3WZ2j6eCte6m6JL3emeuUmJAlqEyjKauquMe9J8pa7kWRkud
luOspGzU160pnIOU1GCigNQcVZAdX5uv07NM+CpLvNN4mWbSrroUwzY2Q2W3edKt
tGrmaCT+7NGM9+lmKEIDa5bZD8i5lBS766Uapb14LI987z9LT3jXX+UflD9ibnnj
9K98UEmqXeinMZl2MlwsVudC0LTKX/vYU/8Ri8GPHVNhrG8NbwXv9vadh4rGQDVJ
SHsiFvvw/ns7r+8YOMkEqLxj9HjHoAC60EFPtf/Esd+UxG+zPwJkQZxey0poQRFT
bZky+he6zDEyWZYE/xogzoYvqd0sCh5rCFn5kae/BRfezTf+vp3uEzawnBQIf1WU
w3KZrNnlSUCvO7YCdoKCaFxgdTHDJL1J00/yHuz4NKv+YKjnu8qUAbACv6Ww48jT
jh7NeF+mMfQXu3my6JqyZ/1oJZeIOqn8BL/a6SxLJszB/1VERxSkR6s4dPCwAfgh
czRJSDPDxm3GEk/r4x+jMT3I4bNDDR2GSzSwSMpllWqAJdfHCl8Q2f0hfRCRIE5s
0e1HyWUN9ukNBefo5ZAYgioEEloM0vMffsgoKNBYkyavkBcqSnkFC702NcZCmv2N
XMmWNCqpVqkbXEffe5Yo/Tx5ScPW4uSLc5CUcvKBMoisv+Xstm8WvKSjWZP3vXYg
sH/rL19cuO7K0QX374zUhwUZFU59WrUzrKVebq3F9N7PH9ykcP9R/QQ5YL4/kbHP
2/q1FJIO4zRxthxZCRHgCgNgH5cfYBaDDDMWGVHxYtbCrZl4jJnuu24c9wXEbFgp
jtEFr1oOTKnARea5iftHWOD9IOtsb3E50q2zvkQe9LjNz7waTBrKlJrzvR1XGorn
JL2mdKpY6Atfw3Neaorlk78D4JjzNhq+YMl/vExfBgE46VgzJZPZXjI+XLEaSSYo
joJU0p2X64sjO20UWdtwLijoUNod4qyFo+oD+jhEMB6eZMIBBg880dwvMzdtoLb+
05dk5jnhN0BPeUBDmOUbm08cLwy6J3X6rjHLwmJPHe9Tib/kig8si9Pr1gy5QDU1
Zfe5lFMEoM97UbG8UAIWjMIo96XKRJfukrWD0g/ZQIrORnXmVeyuq5XP50elUmOA
/JF1mDugDMREArzAZHUOeqAxiFamEwfYOhYdlXxx4/P6BKRKfh09K2g9IwSvyWyi
WIIjqVuKKH5HdowS3WKq5dm3NWZrrtTIlkvaHtQ3XzdoXjeAFsGkN3VNSvH1HzK9
pJ2HbhRprqzHm2QnZby4l7AgHW268QBWSDy6e24ofQDdaqkW2sbWkzvbP7XosfSD
1irj3pKEqdk2oT/V+fSyo4w04IgH/AHzutSfU14/5kZ8dqD6ViuUw2DqlrSmi8FK
ye2dNZKeMZUf1FRTh7sQ0uFPm8P1VGwBDujH6duqqQqd1pxFYxeyXnPeLqIzyjZ1
Pp0YJCUEFO3xkg5VEZfjVtRClIuoU6WNAA/jtN5LWvCuPAkBudNod444vhG6azu4
Cgs19leskmN91suLy1P8zxAZKx+lZPkK6AqBWDGyif4xX3qe35cVoh3hf52CO+hy
aDBFZm17JgEdufgeAMlC/qALc0EuI53Xmbl5SMnDqCIbjJ0D68a70eespr5QomPW
XuPuo+2AM7Y8tH6TVkQ1SzhhPMuYgz3fztojt7FedTRgkNAbdQ6YkM4YbHRY76SH
5JgWT5bZQv39BiXcH4cJQkR7Bd6xNpPOFQUBWNbPDIYbydCJ7UyLMP0F+QeVujED
RzPfvzljoXssAybnu1oZ0PXeb3XcXU2E98PlqIS2MWiLBNmTG4fo5gLlF07wMoEz
dLkSmTt37aHoQ51aCIMsiqSbp8RSIZ1w1fBeDNw20FiOz4xVQ9jxgD4IatmsuGlD
RpZSq4BhkMTf0+96dqbN6WmGOOHg+PYc+/Xf19MrnU9ixmLGzoFVl0ChzpEh/OIt
IqqEtesAwsrLymsP4sGTSKy7aD8GfLKGSyM8kmy8KDjYyVi0iX29tWWgNuDGIBYg
rhrfJTJu5aEmJxYWIST9egj66zMpwijzE5Rmh7TREUPr69jAdRG+XtU7DBkvhnz9
/9Wm4rLzf42SVLwtgP5XTUa3ptUqX0EGbjScq4TjPDEo9h2CZ9YPzv/6qt0SaRyL
6EbSvsBC2x7ZI6soRdKD+zgCPYZ1ppKoN3da8bK9G5w7liKk20mR6yD5p+H2/9qC
IHcCk3tZzBE6SlNR3cCCJK+v8IjtNUR3/14JsYvLFnWfvnS2ZENzMiIdQvFA49gq
0r6YRMWI7g3IWfOAsZwmvVgVJrcac6lmEaaZGMCHIelW4+v06oexJK38C8XMpbmK
5aFYoTphO+JWra9xaw1rPl5BuXqY6sj6enUE6ZMVdIbal9d8Hw9Xu+sB3DrbfsLj
cxff7o0PA7Bp5CHz6CPp2VI5s6lNS3qOPjn2jtZxB4vhwb1F+dmZnNR7YY1LV2Pt
9p/64GQmHK0DS/TbB5MiRg5FLaW5ZOVRLJMtO4pcX2Ut1tJuWDr7aRiowrdo7Gzb
TTD1fAASTaB+8AcvjTDNfD5g8bt45XH2EG/SDdcPFNZhEA6jSFODAmsDXAwPjxo9
gOccPZQSYVBwUbY15ON0/LF5ydTEU+rGHf0fTti1mpXI2n8j1B/HapBGQch9ztCd
Qa9ql2DcU08Yhvg6XiKfyUN42qZHcY5TmLaWNsWIRvMHRv5g5XkG1SIzX/urSwcK
bum0ApW9g1nBHxK13ddneiWxWO4Bq8ueDYz95Vmo2adyPkwXIJrVMJuLnXojlloW
GrP2AXaAE9XA9DeoOHvodGNgoo//NS843c969Kt8WXwIE642Gdej6uvTK4qB/SvY
y3C9HXlnGvZoVyPoj6fi11enTFLnydIrLpACYXJIyu0ydJr7QsAItnvTDAX0HKHv
Stq2wW9oSejWW6CN2OXgohKSlnSHoQkv9eDwnIzlT0n5tAzy673EeoIaZ8qsG/OM
1GCD+4ID0OE5SkLq+aqoegsCQ7illWPhGUVIhC/ZnixsVpjdrbKunrcTWrDRNEF6
jT9RZu1To+i+J3fQndOM4iWiFG9tx82iTuVe5MIUyJr7XEnoqAlZMGZP2qveh3j3
SAcBmCaNAChcith+cL7MfUjQ1uvEP6SF4cOqo5wB7ecGVgZZ4dpbo47CutMqBEMQ
5CLO6uBgtumFaZttnhC+QSEgERcjYiWmII6vDvMP5crHlxqRPHhT1l8J5XKGPXTt
xyZZVQqLLjByI/BIzo6W6jS1ufZQzTD8tcS4V/tHebOLx22yFWngDLHycSDXPytF
YBD+StLDM7+kkmngQGxq8mVEG44M65AXZLjqKdNwk5il7v0QcUPOMz9D6G+8eLha
4dg1bCb5+w77TeAIw+duT58T5RAiEpcLWo/PxjDzQxGQcGG02xEykOySMIhSwYuL
jrMV9s//EYup9bgmMBLZASmpp9YB1uYRutrNEJpbPNd/QonHE79FXSZVP6OF3WDl
UTQs57Pp+SPgCIhm0ZMkEac421CmnLlsyHgp5N5bSGEHa9fpJSCp/VOzfXG8IGyq
xf1AyXaU6m2G9CKx64WHuqMGcxY1K1Uwm2pgYy5bTiDv9/J7RwOMh6p3GgN4lAXC
ymJ2zFUkYGQL9cq/nI6MgBzyIzfEHmsVXnbTiQsDzobXLIwuVzkSy30g+ljjdHNn
sLhNi9Z5nPTdwGWa4GHtGro8t6qZ/ie4SRC5J5oTTkHOr4IgMLgegr56sFSJVr6z
cJRDt5MhnaFyztwLVxswHWajqoemVqVigqAFdAks2kzoed085RlmDrZ2io6xj2fI
EcMx5ZhNQY5WQmmtGWm+mGDmF7L3TZxl1jdj0xGtLDkFsHP7MqYBT4HO6efYvlNi
Afe4c+IhCXL1NWAP2SymZAYZrtMMySWxwUy3m5+/ZfKsZvg4NgmKPCHsduotuw7I
iFe5wVy7/5Y3jfYxX7KG9tcBaFoZZwBuSymVc58OlHu7dFfGToVaHCek+z944uo3
da/nAoLei1msyGWZg/jFOVfQD7KjX/GD3zln/6jFCfvR3++JnFC4xy5RViOYsAlh
8Pn0D0JtPyaH/Okmi0gUFce3ILt1f2V6IYMR5WixkI8FG5GeW7tr/iomenzPuukT
zItRPsREXGPmEdqRlsOGKOwUrfLnv656p+hDp3ZREVNn9e9dWf8srY27nKgEYXdk
YkRuiIKRwUOFs3NM5R8KlTqDi056Oo7CY4Ng73yh5LW09DgkNB4X0kAvX4ONEJtk
Nb6kqyFl8hjhZ5Uw005pboyiOD+lns3G0WEaZaPRTRQnrBNTz6tj0ybRrP0M1y7m
eI8khR9SvgkQZuaLhRp6DT726cSx6sF4NSGRYmTfvq1BFwI0A/v5ZCcvb81QGUOg
C7UO5XXh6CRtw1PkFbBHIdlsGQPKSu0IL2K7Hy+2JIOJbNCLfBaLV0wxn3ZdSBSB
k6ViTuqGDA4eDUjAhmfxDPtyn9uuj0g1PyIYHXd//cnBo1GMLFwoO5tEZbM0rJMc
yknzdHg0OXyymhURhO0gaYAliZIoRRjVtuupiPOgrwHuTY1uDAOcSjOLD+mv9u5H
AI1pTfUinxwgMscAfjQ+M9z6xfNlorj/hdXdq/lXcGDPUNA63O6SYSQAN2PSjcTV
v+dSiTdGLUplnxWSdO+NAEVALG399W4np3lNF3OwDfJ1D0LEgkDjX2q+EfPsDToV
QGnXXIz82eEQ6Z+X0MBygurikJBFi/0IG8r2hp0LKCggVjCbOcoQENJ1YEx9Ox/m
gp2oREP1GLAByohatKh7WCi6oKv3fWHb8MmSwe40VJt8NS9DKbS2XJ055kxwXq63
S9mhQ+f4YBCpoG0KyY5Hm51D+fXNWWaJIJgKGpuMjQYIS+3xm0YDTaLeU9A6HYwc
p/tHC5gTWQdtCr6wmTwJwl+P5JFIB+vPv3RAlMq6ZKPPnQ2BCnTRd6h/nEZnBqlB
A2tlRbHJCEx1ONJOQycEqOfyQETBqE/eAg3RrCxwlwnB5/8sgOh58En//FtkwviX
GzDBiJ0nIwpfg1eIZKiX9UulSDsUT4rA5Z9xz5/binvmRZpjIHemE5pNho6eBriy
sOGPJi4d429kizSLm4higPJErnQH4T1xThW46A1jLmxxpKEWDnxBgk4POBlcFX+V
Ds8fZ/Dj9ClM8MVyGSxA8iQdu/PT+wOEUMUb6td4/gzijHFJ6Yr4/4Hyib+vlLH0
VrB8qA7weRUvtozRgy61KppnvwrwhVswPAYx4s1hcKH2S0DcQ+F5IH51wGsxgMbG
Ovf/Mh8dEOPMYSNaLJlKGuzz7EAEQblUnR+Eqk92epgvWcTPCwqEduVs4+AFoYlZ
sdfPjTCueqlESLcHvgHBlb21GWZ8HbAmaS8955xHq8mJTYhYK7GltnkeG2IJMzpJ
RCTg6kRvSNrsjO5pCgPc1b14wUoFuxUCIWQZ/dPO6L8me8nDmeIwA3Lh8fx18Tpy
FJE9HFX4RVSI4S1bL9rvg3prPFX2T0Jafnt5IS4RiX9IbJtx0/uVX5nKR/7grP5g
O+aYeLTJQH55qu8s8FXAcJ6P9GxhDAkXpiWwHbHWI9VC8pIx6k75y2qAUuQP8Pwi
H0aiCSK3hfMIi5vTTpMMxepow2ljoYQWgSBKIhz7eWB5vx4Vk6vGBXch1JmFqV2b
NQdZjEJ8dqM594w7C0l2SkrXhi2W0TY8Z7IUnZC1QSMomgYIMWE702/TJwpIbFGc
k3kJXY2I/jIJBZSiMbpuaxD6MyA/j4HHnpFEEBD5TWEHuBXEMWtPLXFepBA79CmW
cSckT4TixOG6a0OlSyyPDVx3K2ZPff3gR+27SRrYpzvDrBZ3NG4AolTMVBs6Hv6n
TkGzcA8sY9HRTL1gEUEiKqypFGs0dowL8YvmyUTus8TYNU2km+8ipvG+kiKPahOw
19gL/Zegnh1dX4FwX4zxHc4FOEjsGqki5Fw2hzbKb0/kDpcRGHhF6zI87zQIv8y1
Vj2Lue7Z7srcrvgYusvWSXDQgaJUYxb92xwSugUYkLcnJ3ri5bsy0jDtDBi6bX+I
XTtsIVlqgy+JaEzDibFL8aNcdzJF9/U52w4S7dzwhvfD7O5N0fjBuUu6pMyjWNHl
GDLNIFXw76W0N0rG1MmpnG/jccERUHBBfCr8Lk7IDeKaPPZYsjaWYUSezOqfqNTW
dzNkwo6gnfmh9mLH8ae7oNTqzY4s0y/MjzopCDO0sTbGkaAqn5VlPpHBdhBmcHba
PztqHeXgHztXX1E2Q2R8mR+9Lg4jcIRAaWBxgCQFp53wipkXJmyNjuM2NrZbWozM
4X0C0yA5m4eQwzyX1MWOL0V+3cV0xtl8KZiKNSashm5cQKzvmS+70D1VzfMafk/h
sw5RhP3FbrFYG8y3iDJM2AF7UkA5qoGb1PERl0KPI5Ccbwf+EQYTyR8eu1/Y3mA3
W7F8r2MHk54OFAf5w9a/8kaAvXbLDxLl5APhfWygSI5w3TIdo1gaG79lyjM53f2N
CvJzsJX/Ohp04LM0+Ff/BtxtizDxZBFhXqfJNq8wUNUfra5VYZByKlSfw1HFjkDJ
JqohTFSxZw1tc14s6tbAZXAV4D+SB5saVIAkoAwF0Zf8HABDj4stoNpnCggjDaQV
iXIoIWtx1u/d8LP+HRFZC42503qpkZgNUPU/SM7lawHNNDtRC6TCQWEOE+r158Im
CxFVMMzXFxZVgoDssTSwBAtNFpx4WSghLmPPHieyy2CQHYo2LtkhhCRcCbQOSdrg
K0CcHnkMW75XTjymxUCMHDpGnqyNPyw/o8LZD85WfcLU3gqOBBHERMyJqHBu0i5+
xF3kEEsGs+ReSHZVZm5c02toAu1cp3WzCN7yCx8/cDiI+bc3GZwWhyc8fPkpm4nV
NWTnro1IOyid1wBdA8C6We34rJQgVShEEBnG9BU9pvh+qWXDV0BDKTqssQzb/5+o
s1AgnlPQ7dWcju9xDy5BLSb2lIOH2plYi/OxUh3xTyM/dJNzIbhofbRpKbdU068T
iVUgAAoyt5nWByberRfFamxIZPt0sssffp3FFBLlW/L5AYRE132Utq7Uh4lEp/dv
MaM4ThU1qU2AzgPk5C/vqkG1WzlLG4j10ElbYtJqCpOWeul70znZkJJzFAGyHZbm
1oV3W1370C/4HJoqtiCFUWV4V8UdPx/TFFCpKRhmhzJPSm+D9GkXKnIfA20npMdK
7kIbdoxJmYYsJ3q9ZG/6cyiZ9WugFW36llUB2s0N7HSntOv4rUUXHOGlYf5tTEqz
XSuYSu7MMob+9Kxp7cJS8GLR/RheHlJixXOKcVpl0RI5lQlQhzdQDOdr3pagBUzw
FnFDfbB8i57xGRSPWnag3lqpD1IDgM7igQW8SPmebshqDQlqQWm+23xszZb7l/o5
fFAWoKNJxnnamAq7g7iWq2a6b20CzHlfQa1DNA7xN5kEQVdCUVLGCPKVK/ILT+cX
z8tmRYJFBtrvpYoD4Xt0ipnYqwvF1K4XSwaVa8vdP/yeSVV5ad1YIaovu82Zl0bN
AKXznE4z/KZE/+GH+oT0jSZLo5XKbhdQqf+hrrjYUsfxtPAj3L1/HIemPGdcQFJr
gZRwKC8G4cDFKXfhPR6YSJscTW0i4jN0G8M8oMMUDV/J4LaVk819GmJvnJGC2Om0
lNwqYjb7A5Y7NxTd1g+2gWeorbjE9BinSbFkpN38WKLh7iU5J8fR4ioQMEKXOCRd
Ld8md8C7z3jTt/rraqB6LNrIAumOMkPAzrOF1qt4GdCWS6lHn85PFoiONpmxP6eS
s0bi3gGFfJ4Qo4+XSoi+EJzea+tPzSBS6GZnva/meAroN1w48n4TM+xylnYRIKbX
5kxCEuvA7hLwktRE9rme6Y4xOslHVkH63y4DpSFC6vRv4Iu4htaRYJkEn9ubffAS
OUXLs9hN8mhoKq5pv6yI61kTZBCOrCEfXxeKqI4Ai99VnCQG38+PHYdPg2ttVJdi
qVcpE9VNYIwQTI8lNEjLSVrOWm2mVPUiT8qjKbKUOpG9oLqeQOG2qaZo38/Clggp
FigsKQiGnqtDcX/yWb0cvdbEUXVACxbSUNW/LCeirbzQVQ97YCJMm7YcFXx4dEW3
6CMAAsNxUwekLKa70p8iPfggUqJa6e/H++M8u9IFYxVabJN6uh7uAvnrzpEGsYk9
WRc92/eUglOwtG12GIwlVoIBcpzsmK1eM4efvL8KOqtrvN9ZD5PYmbrW6UFDWQIG
8Beaa9cvMWxfmOwss25aFb+/npat9WXsWvNmrS5xurincuKP4weA2Xj7NEqQwTHn
BxgGxXyX4/qAwm4yjcL25kUVJ/W9sfZqe4VgJEuELK6vg420yPu1pHCzfu+ekum7
RwkOwo8whQHcm6Ey9MjdJKgichfTkUOcdIzL3EPWOen6eS4QNUSKV0SczTb0Zrdy
mcrOzo91qijTvwmwO6KbsBXND2vpPR/hpg+wkAVZuUl98U4PTdjiR22EDMAPDIOH
TiXe4MTjywgdBkYTB4bsrSCCpgeAUYEGNHKprHpLlLixHyRlVoL8lVsxk7sMfeUB
UW57WJH1zOo9jMaD4k0u9ZhD5uMZAOHdg4lbuN6hAxwAsZSjYPUdoSLDZ6iplZ90
rxm8Krgx1ySixB/fD0qQcbxw/1iu1fiWvuA5jbPsJtvHM0l5MqRkl+QL8A1Mvx7T
CC3d+uiqwMQDgUJZvIU3C3KBnFiyCNgVo75a5uIvcksRG1HBQIHiB5iu7j+KhyLy
sSUSjN7Q2Ku5F/LSeHIr30w4NFFjC+fT+VLHwAGCF60Jwuf7vC1pjGLUKNVg/XZj
RiwJ9EL8J9/owzT1k4eej9PwKbypvvVs4ia2nEhsBcrR2TtgJPhU+gx8plfdjmIX
Wj65EUnTts4CM2yJd/UD3XkWZB9+CHXTUquYZknO4yOSVYKTm5JeAOuGwteHWnxT
2ofhv4t8KqtCMZjmEc0J0e2WvT90WINhhtW/FA1cIhDhgUqXC/PkLQIJluzv+ztA
ZqPi4LlHM5R24F7ED3CZBFntU1j29xpI5VXOc7PgEBJbRj17BJaAR4LWLCTCo6wl
ex5myauAFd1PbcJQgibb0LIGWiAdnLBexrFZtD2BWzVPl/1iUVlMjaTBAoTJ7QH1
q6s53A1DN0L7RdHjtM8H2OX9bThsPAp3OadtYKMwiKg+YoNpPXg2CQUx2H8/+Azg
EsaudYbo3xs8ThpnT4cJk9zm6U3K9tLBFdlJHLU2YLhRPAJmiFgWavw6+OEd6s0f
4NR/t1eMUZSaFMEjxH4D0egAq06ucXyB7MQAycwYLlQhP+kWhLXyu4PyKVyf1UTI
cqArFI47NMVrHYk9fa0yPmdnHoHzN2Cf0F7Qxg4iF0Xwg/Rt+q52JPCioR2A64P8
q3faDY2/RxplMjsS3Qevw6lTgsv6sJ6MPQhlLfjzJhvglimXZIK8ob6lygnnSgGS
H8qP77fsAMlkDCTnW3AnZ8MgEJrtBd6EucIhK/0wFXuPLlQuiQu18r/ibunyPoqn
JdlZI0DB/4iIoRC/WdaBGFjbxFkdA7wecmWFunLppRMYeWmyxInBeYijNQc9iW7C
+YYjH5ASyh3g7gjftZo8eRTy5M9fwU4mojObfgrJNcXiR1UFdW4E+8EIjhsj8yNV
zLT+woLGcr68b46f8C/ocIvfv7Fcx2COmfoY80zOjX3Ws+ownEOB8LVNbA+5noIY
Bk2r8mTmHjdT36tfdGU5Ju2wurWr9wKeAWBndZ/+9XooWt2gzYKcCjIx2TR/9nAP
H3SllNEwO+q3f6AU2jMuWC+j8TKsUIegofk7BsngFwh2kmlFuAMKIqTPnH6CjvhT
9FPC19itt5btDBDrZVjLvgK+i+HMZS3mE0hs+WiF39OyH37jNEMOuvexm95t3s/A
5odaCDceimz62thqGMVTrKsWLHgHaYlB5u/isGg1miu75m1tfq4fqN6SeypB1Bxi
VVMNDAWpZ4ugFT82PldNwfD6ybR+f42rDsYnY7a89+JsFfqMPnAVpDyrUwzjrAOI
ObZuYb0qoxs+DuqPYr7fJlJhMs02lDGGq4/kxKAvBtmsbXbhO93rXM1m0ErBbZd5
vF9WVi5cc1ItAeoGgmQOgTsu16toaZe0Av7hnxRjgEijsvUYiWEHyf8aKmTT7vpr
K5xYYzh8pi6Osczl1UbRCoZtO/XKZ0pXVLMX1ntmEIA59mzbh1NfCpKuZa9mxDsH
qEpXJLTxDsW1YqIg9nb99VAlqJ0PfCHIOax5uNyTEkQNCr0u5xL0RifdmBuyx2+x
vuqwzM7Kzzbp0CB//rKg6YYerBKZkzVtfMvJ2akfD6oF5N7qsROQuM5vDfARVrwB
NA9U1xnFA3Fh8dSbyKqJ795d7IVyt7bFWX8Io/M9lv4Xx5fvCDb3xCHCuZFCQFKc
awDR4cXY1DH0rkw2Bss+Twv8N7mFrJsSZMVFwcpbvYuuKLVa4J7wM80C4bKwUb2n
qKwFB0Mred34pLn9Wjhvc0x1N1BCtsjVOZwjAkdCpnHkVXX3Ia6v0HfXYv3ZTcIz
KHw5gl6PRWhtQEZYyR0dbOZLeN2sdlH3PNqYnTGcoZhjP16k4BnJBewD8KxVkk5f
AD9FD30zpu/0is47cTp3kD6iP+qjerZUaSEhnu8QJotTKeGBkgDHseZHq+aMupkQ
gkq8zHkGd3iT10WbvxpIVL0UejTbJgceXF7TFEm16S8mFtY9dTIOYq+d8/Yqd42b
KcXeIqGeLzC+HHgeTi/b6Nc5KUHMuhRKQ6YD6WQCaFU/GJk8cuVPeYEQsCCcgfGe
sAqHNMj+DN72lKTJRylpzy1txF9UDNeoC+e7mzdfaPEZYoI3hm7bq0h6ZWFKKcWB
m+DvaibLNs4UNvLyPrBUxZW26nr+UMxJVZ6VKK/LHGtse5fyn19Yx/y0j6PY6Ypa
bMocvQQtlORMm95+sXhnBiuGRNWoYvwgUyp9AkYz+b51yPTFOUMffk7jUGyHNpFA
eYFHDlNYDqWdiHQD4nkx1NZT6rD7BAi/uzaXH82JFKtNJZYPgkg5Jt339ermQIlh
7tc8uNORO+HzgG0n4HAbn89MjnPGCo88C6uD5F48JtycdOF0x1dOoALC0b9Ca8Ve
UBT+oB8iZwDHvbZEk3Hz1AgRXV008GxJFRbG5x9su97THv/AbqOHU2B1hoC0+ExJ
n3duKWICZA3tNsg1k/QKKpVthYIFHkN7TVo3zHlZBX8PgA514aU983QbTx+gcJ3e
/3+7YVbYC8kMiv3/XqGN4xOaIxDqjhXvdNWmgbzVA0jXVEvRWfJbnaytqBHOhYT/
NE1HPCDha0l7gCtp6GRUQutbZhOjM7/gmVbE83CHlBnnn2PFHD+nlCGeC08Sed2W
QHfqNDstgGDJhdGMtcJQa63ySJuL9S10jikNWeqdwvyqJpoMvF1LFUdP2rGY/y4d
1AXuf5wH5rFWb4WTowitBcvdOPyt9buBwtvUSA5zBvs4HJQmg20zGAIcelQ7QFW2
o+GMRdvXUGMH6lsYCFxP4Vbem6ad1657ZKpVm0sN1XObMvhDr7Ef4acGwnyHvY2x
RSFUkO85wV5EEkg80KGDGY9OYZn2y2REgmI+TzCD1N+QiXvbqDbPw1sPCf34O5aj
ZI6TbtcFzL6SwxkojVE65gIKuv0LFjp88Cdt5TB437bkA8EmBP6kOMsHyBZ8s0Eo
jgyGJdafwSU73ASyBENFl0eJ7ySVcEt2jvId2qsr6frVA71BPFakZWwxQAnVdRI1
cN1qluTdUFuPIIsunpiRYIkqrcoctleEeYqueGWBsvvdjQjiOobieIJQ/xOm8O2p
4RGhEkoeBx667PK240ow/QyMUoIfEOsTrsKn7inGN9lZL9ytZeG6QmkMRumtvcvi
8ZTkyKecZ00dqzM6qzdfWJmFoby962RRM8ZTPVekl0c=
`protect END_PROTECTED
