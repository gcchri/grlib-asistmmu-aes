`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EAT8Owxl+q3Fni8dri+wEf18YjbB0l6kOYHcNPu0qVlKe80IT5w6uttQoVm4zMaf
oCuS4xPm00UxCM9szlG+6bL1Mn2Jd0SqGVhocKCKpaDYVNLRR/4mNnfP6Gh2kp1m
4JxdBlKath4pFEqKQbYnzA==
`protect END_PROTECTED
