`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CQV+6FRiYpJeWGhtb8XBjzdnZyoIayyGMeXDWJvl9C767FQzjPCbe0C68aUFBJf5
0z4PenuFZYiK9d3mWT3aJkqjCwUrv069/GFdsV1akApFd4LHtE+41s7BcD9W72uf
BZhYgnm15lc+AopytXKqw+eJ0nj3f26u/b3as07oUznvyA7zCQPKv9OpNnndQnkd
J1Xl3ulk08IzqdvK+Ll49BPAgfnBZzISPb29Y3tXa2KiCf3omrvc0yWGeVvk7oiP
Hf77j+gqjdBTfTwXUGhPRXMMvmJF4TQJKrnApZqEPuDmHBcxBi3y8odjs8YR3h8P
c5m9GtnXRQgbG7vM8dxn/r9+ivq0tzRlxcUL3egZfK50q3uZHiHPASIWBO/rOfWw
e2g78DJP4VC8klVDkqLVlVM7UFQhVJaQkdPEhdvZZd9xsxKGLJb4ASFJ9R/pBqIt
xeGMH+WNbd5ppA0xugRbDSySNsDBD5z8CQ7+wnVsDSiTAb8Uj0kDyjNRCGgRInIk
Vb37pH3McGtSLGLwP2oYRA==
`protect END_PROTECTED
