`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dbgSDP+aJV3U+MMfkSygdkD1oFe0god6KRs3weLd9yR1hQFdg62LLVdpQdbl4jKu
fFNCESh+KfjgxZR0X29nVfQwClzeZ2KWqhUOf3abq3GRGxugKpwIsufkj6NgHN2R
MMrzVWnTQ1by92lMbNs6HyZbva1sG1jZzlMDy0s/FB4n7L/QCM57EKEnL/8R0uKH
SbwdmVteVh3un5VANWjtnjCe43BW6+A4tAo/Im4IRIAhw0DJqQikKWwbM3xJwtEv
d6HAse4ASmM7i2cO7EN4hNC8ux690Uh3GXidiwOsPK3SxXIPvUa7HEiucPnySzlB
Y5Rji90a++vAsFILS2yiOkbrnrA1AWnel2ZB11PwdaUdz4ndaKMnBb1MZf1RdTGx
8cmZyyd3tN6914nV+gJwpiJ+zIFZ3eqMaf4jSUphyuFPdjfJJT5UgO7tfKLz1UD1
QRhd540OxqRGaxnUsUPR8A==
`protect END_PROTECTED
