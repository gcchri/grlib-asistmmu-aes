`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3lM1FNqceSbKVUDyqTAXsSxqD/FdnmgHAyfoXQorap0YA9S5KAJqci5czG/muXsF
nzAPdG+f54kUkOG6u4AquE4IxPVSHXZPmAC5dVAzav5VNRc7juDUSXey67DYZfUF
RDvBKN6mjezb10FPD/cNcHTicjwZ0FtUfpoAkOZ+wakzKJAxIErmWgOTY0/w3GOB
DtNsbr5OZK30ug4sbMycQriLns1fSQIaIIoI8OWXHPAXd2KKhO1oR29uJ84OxtLu
xWpEzTgC5CmZOQ+LH30oiVMX7mV0Ie+aGIx2c0Ac75Rei3aRswo/1eGAKp6pwAAU
mSP6TVZ2NXQG/Ui63OYgxMa/8KSbwc2LYwgn8MYBDyIaqvLlj/CgUZFm2XtV6GF0
kfFwjyleWg3GlPMvRs+oieRKr2SrjezqguUlPXamgpyCTomZHTZ6b0sqEFGfOw/3
KNV6NB2ajMOgz4cCH5NERT9sQLqjIBq2J1VjyMteZ7RS1yP2+0t8kLngjelJk3q7
J/z8Vc0DaTWkz4G7lDeKUA9bnTy2F8T0Mm3w9fcyu1rYH7gAgErvwHWVOj0ph8pT
RNu8R9RKP1Cz32HXuKjVgM6lzXUl3LFt0TBMJIyrbS+1c5AhzStArucslb2Hyiam
fOLC4a9XZTfnHmAGJAQdYNiU282u0JELxxKHkvbUU0Qqp0u92oCe8EjnjZAuXM/6
e1DYoySymF5RH0/f0StMMbU2+biVArHnE0qP8dwU2xdY7SQKN4IlBNdPEm9Yrz2C
6adhnLswStAiHSrojFL3++ZDf7NFK0czYZv5XFZaXwg3ruVDzdq6I7XZMQICYlgT
tCvidAAHMs6UYFUJswIgP3+L+y0fwLka9UVqgmZeZBcboUahybzOV9SepnGMsmvE
+knOB4JQF6laTnE6k6D3ITKVLxW83VmW0vCcGbk2zj3dTpMMQYhI55y8xLNxcGPN
IjH4utjtlRe2v5WK1L/dQJM7JSv96+Y+S2iOu+KeR2IK4RCm1XI8Qep/effs/SwQ
HVvcajjysnWae3V4DjAAtgmzpDGDYTgJVB5hAcl/6q1W9IDNvk5iEX9ndzze79lv
EezmYmBZMQB6EL/X6H8d8BYcyRVz2Oui+eDorD+fuGtIi9UfZ2ihVxuv22MMj3gM
7+NeOcoaDOcPpHtH+n3cfhL+uM6hdi89sor2fhKbNXopewa0hU2K7+e2mGT560vk
lZSWi6G/HrYntz2A01n47GwzjnTA5V3jLSisW5hYVVdSQLPqVmI+9ejdbFxiDPQW
lzThz/H0rjoho4EfesDSB+yhI9zV1klwFAqO9PPuBGwzkZaDUILmcWcM2yewWoH0
2f3TtFdRn4xlCwGbrNM10G86HbxqIRkodqfGdN34/E3DdFLT8OVtK94EPyDvRCFq
Iv1ziwHAWgWSAcBMR9dPw2DVJZsK4uzTIk4FMYO7qH3mqO2ZXm+gDcQ00r3AB+Y2
0VB7bTgc9xPa6LnSxVV9Q2K6YPLVLgpgZh5e98OUzgqXqFHoPiKfxQqJLN2tHSqy
ENCJgeKCo7nxOogkowTqhcgqkeYnZe+k95qqRgBbUqjlnwZaoBfzukGoje27XJDB
JjG9wIVbcHYsqV3U/yjjCibRUK5yD8rA26CFZoGrs8prjFsplfDWThwcIn9GC2fh
iunT9QMRxuo4UT4bng2zGCsDA1PHOXV1knDPpxihvs/DxQPXBFH9yAcb34h8Xnj2
St/iTe+f1glSy5BhylrZ1e8kvs5NUdzm2Rgi1pUaTfhNVBkdVPr5iGsnMCH9qgn8
fhcjDG3h/d/VdC3lD/MjYYAI7jcBWdtiHT4lWYPLYDT8vRjmrM9Ia9n+jTOB1EV5
LJsSfv+rLyR00Yn2ZustyS8erCb+TjWFIe7l81Pcrgu+RBZh9q4lHmA58UBTFIHt
Jv+cb7Up4Zg71x0kgGtKZPm6ll4Ekxg7xlKeGqe9sr/DnrCxe3xWMhcuM2pA2wDg
gq2st2js7tkm7h69nJ43oqxPfXI6hptEfT4qyml2XGE8/GlWuuff1/M40OA0bJVE
EU6cq6Lu/1S3Ut/y0CxQ88xDq5M50D2A8UhS5zlTRSjEa8TfXy5py5phrEsL6/fl
uofA+XkEYn+WhcwhyPkzc0HcZ4Ln+Cp5UJo9QZJGsNSwLLp75tShUPFJsYOWQz9r
unqCJgRpEamVgy5HX+4LQkO1fllRgi+aJmHsJ81BfOvSsE2aX4biN0j9vyyKhofM
FN/G2ki+YMH1v3ZmYHRa5EUy4gejIjvsYnjPF67yCQ0++fhfwnkgjQ5dmtf+iApW
YcXCqJtwz9RZZapQ0UFdqZJIFyXoqCpxCur+0DFxz20J6mz6iMJmDG79uRig4/Ty
x6qFSj7Nqkt5ST2dspbHSNUqKRQoDA214PGsXZxbFkPO2cBuhn+XNsLF+v0NX4+B
rvzQwsXNNFLqHGDpmBewiTesrMtclilxfI22Awv+tLtleepguLJu3rdOs7F7UwB6
wLY1PC/fhMMsWlnTFEnweDCQOV/7et6hfxp3uMJeoK3dDOti9zkZBr0CoLee14Zp
okJp4Z9ofBhVoJKM0ePu0KbnQPGhVDZ/E1rxU7I1qwPwd/Sc+PSsKs9TVhqARK1y
Zi06+h6tGmYC53XGwH2aFwoPgCoo9lvgSLwEM0n2JDvWErawsGtkc0+Zz5ChyYf8
PIPVi4QgwkEV5kIOSQfqVj/81DPrjkhuP9iRV/qacWgH3v/XsZg3PQlGiPsBVebH
xW1c+qoFy60GcdpyV3jUBhDhn9GuhXHwzCgLC4XYMGkHtcDNxTEcm5eLojTu45Qe
EP9j7afLLKbK7AUPQnNFV+RkuceBcddXc0BB26MTCJKqw4uA/cYsjIEggeMptzXA
ytQIQp73B8Y/pjxOkZ2QRssgadxLzeDtd1bFnfHj/3z5B+qspMPpBk8wuQeZXTnZ
OdLE8yCmlgqPPnzp+B7vgtl6C0hE19quXEPdG1sWtUJcBbh59Q9o+iMB+wwoY2U3
QHWuj+cgOFSEXO9I/DrnAPqzT8AsyxWdWxSrqRVYxkf5TxKrUfktmGtm1mGWPOE9
bC460IciVmfSF9uQtopXvr+yWwzmYzAWF1+0UlgQ95bk+bcjYG/1Lnfd/CW9ZjsY
FJL7R6qoP4kdO5XtM/sMc32v5oDEfz5ehxB9GLGzMZUgKJDRm9z4Z5cmhr5/lcnL
q0gYYHyzHE7tzvvaAXN7sT1S74iDjMULZi5xeQsuO/XJYT0rHwkpU7+1lnHw+0cM
tjYbJ6jaKg/W36LvjFAZKc/7H/RBXa0lkj1HhW73XuFJkirwtEHAg3arZUM5ff5g
OMszZbWUXGGlsU7b3T98dplywJQmnWYjVl1fz6wDEbgRUnYuihXT1vHbS1WWFmgr
dm+Wa9UTfRPRzyn2a9lu6eIRk8c+jhYeNpH2UGWFpj7VOfPopWd9MmEgkwD1JAzu
BdLAsAwRxB3AArvMyOc9+grMffjiqqlvCbKtz2K+RLicmVJX5F9wphYfY1c+FkCB
1W1KbA9/36wPi5uNfivSvpROrGVWVoMQP4s4a9YG/j6hqyzjKKnkUwjj6k4R9K/a
+uzfiobDG+5jYJzIFTQAQLCQvQEFTU7zA8GNvurfJihc1PCpKOCaG1BQvhLjTaIq
8mDyTFLQoQvWN76DOjEm3ZU7cWX5+Nfax4ifudbRBrlozozBWWccZfnScPlOSOnL
/r3J7c66hWrKmaMK32g6gbBDx2QTh0J5vntg/G1Iz2TmbP2r7qWY04JY5XBsdj0c
YJNlHklMAOfu9++84kF8EzZha6NB+zn/twV9Xitlcg2LUQUcMHRYqTkayG2MBI+a
aPxhsaH5KOako5LavCJszkAF798ps2ldSdPS6HoWmvQApsQ2Q2zsV4Etc/K8NJoc
u8mHEUgj2hPzvhjJDQeHpAaYQCnjiAcFjI8O1hkVcC+x0YdaSr/fv4WBhnoHhDOR
wvGo4dxgAJLq1SDPj4U8B8OBSNyz1IenJa+2TyUgC+D6Da9FjRJfuCA3pFBzIp1d
Od9k9uql7UVsOhIHgk+dIuWd2Mjq1LImA/MNwUHbJmitvj7z562LiqGoHQnskxTJ
/o8ZM9Bhf5bylLJkxUyd7abG/hhVCZe0+5Bpz5jvBvsBo0Li4gyItDaeVtfdE2za
7ek6ODT90BhMzc2BCK6LpBFuwC8uAMV2bJOAFnvz73oP7WEZfCCRb//0fRK4MBUv
OiBmtE2NdhgXTglJmoZOvK1QA4KhFA8zEaBP675vvSm37ExuBy5whfeMmKvpV3bF
lpdTTV/D9+cgyxQ59/Exc3ODX1wocj2fXO/FomNKYuoOrqmlgdqRWAZPbwt12sci
MJf6XmN4fCi8r2g5P93Y4p2iig+cZXVIqILhUJ2OSzd8S1BS75MIZb6fXLhsJ3GV
CCiOK6XDZXvSLYHJeX1pp+1yrq5UY3vzCjBWuoG69dk1ZgV5Mv11dDROjbf0i7F5
n0r4uH0WyJcwNByPbrkIWWfVa4Enhqom2C6ZVpl5SzWCXHsqTAyXoZ43nCupE7W9
AX1JS+Nhb9Zd9BNCsVlollS2beiImONKW/DyDXnklj1+gXiMsoF6CbPisHopKQjM
dAhQ1xzCLeGzTAo57pkbUxAf+GrWuSL3J12Xk+M0qiJXoD6ARi1llKOiqA6K2k/w
0qFHpVh0de5+ZzjeF1av4A==
`protect END_PROTECTED
