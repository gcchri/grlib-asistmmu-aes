`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jhuudI87b/tLgCJL9Hzz+ztiQecnJX6DGxLaWU9sP1HQPqjR35X3BSUtehLgthC0
PUzFenzcEhZ9HfOFVHoJOJB+yN3BoqjtSRGOkodH03BLl3Ukv3BkwkApKQ24IyRR
cO/pDWvuL6WkCkIZWBKslQapu/oVk5od2Tx3YUG2vsPniTpcV0dhfNSSP5DTAQn4
UZbQBF4zYAHRjoQInOreLUY9yod1c6MdZKwZTDtDc+vn5x0S3qw79gyk9P6Gn2ml
1DiZ7PJ2gOQtebbpKU+T/5k3y5h1xnBCrxhJZVzKwYZEEgbgBkjMVZkDfyr+ONqp
j4+++XkYc39o4wLz7MSLJ+NC8lmSRViRouHNqkFx6Ak=
`protect END_PROTECTED
