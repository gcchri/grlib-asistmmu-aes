`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tRlH6onoB7YqFhcMUKGA2dw0lyfbt4R9O3njJtykRBHcTR87SPTbTiY1wH6lb3YA
B06Gr9jHNQT+NJ347kCOTP7031Wn58Q/9KlpdNMcdd6FQYaIsC4571xE6kUqSr6A
LKi31s4a6iuBhilENW1kFryBElo7ypgmISH5CtWyc6VsVqoLtRgDeFuTuF/8fPW6
OOGBkz8k6khJKGAALvfwFaClSzKBCeCNuiijwpONtx3o4s7kW0MW/WJiFG7cEpIy
TMxJYYTafqI2LJR3aMHKtw==
`protect END_PROTECTED
