`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iuoaJ8PW9DmtyxAgTp9slj+qg/mKw6tPU2gqmMazbRt4q/Y0Znzczs6i5UhL02MC
QZa3zGzvI48cimy614neZeJ/D725lIc8eJZohGxciuFNauT4AOBHllbd6EkDrczr
jd3IBRvcA6gH1GojHixxChtx+VHifYA7Ou+8LRtf8dbodlvs9QX/fkm65zZ7lp8V
FAu/0oWAlqcLzKy/LrokOmdnXVdQp4v4hucCo1zxo/yP5fj04HzUkAUZatbwWFpa
fV5l3M8lUFFQZUOz3cV2877RFhCdO0Ok55FfGOTr4wgMFwKGGEjtsJId5zyo6LDX
FXuDEps81k3QPVwfaLwYJ5ApnJWQk8HMFknF6D3IgTE=
`protect END_PROTECTED
