`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uQ5UQlQDd8CSWpJLUIos+1IYw+qeLVNzg65WL5joHb0rQ63vBWybAEE5W79LVJl1
t/feJSOUyUxmipUrUpn6M7v33bKo2+J5SjaWRq3xtqpFR0Iwf2jR71TKcNel/7q1
LwoSgx4dweQ8hvWWw7wwIX0W7umU4zqLTYmzrP6ic7luJEAgip3lakmyqyZ5bfYL
YzcRk1/Vj/JLY/u5VxO8nx+0OVoge/XVTi1n3VJ8JlhlgGHIXTWv1RKjp6VlVipd
Ds923SeoU9aFec4iseJYfp1E99SsmiUeosEYTUJZZ7iYOfw9hB1dueOA2Wt6ZD4z
w82RdXMH8POKSdr3zMbrNlhlegOI3ZZ4ZvHteNudlqmLMVKHfv+zXYqKMPHvCrOD
oC4mtli6MY3QVJGBneCJoxoyWoibcDkB4QssTOa2o6Z4fhQaxpJXtojNDKyXlGFG
Kz2ndE/SxkOC5txiW3qR2tm+mi97FaMye36Kxgp28NE=
`protect END_PROTECTED
