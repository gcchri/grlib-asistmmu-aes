`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dJcaIAUGWSOa6FTxzw2+H6QYkHA0q31c/NiNbBXkjNO75WbUuCXB9Z720N0EV7nm
U780m9uip6+vm4cUWsGPO/bXlNxLRaw4Q0vJZcpEt8COCIbTWmUB7A9Ib4h6ElPD
u4BiUvA8hdY7x3Ey8BMwzJdKrNiMF8L4YKe7j3ZhMPkImG706AeORQpiLhu2psUn
OMFDKfnVRyegMKiKcfqI61NOs6fY8HddYTn132q+ZFOPdKxED2yG+QjYzLVvG+J7
7hWdV6xHGHUok7p7b/gSdwmxioImtI/cH51qw9QdHj+W3ncGMJ/2ntYm0a1rUf8R
+V+W0hzXxuIu2o5l7BZdMmvLRHF8d8x22SEfTBhPTjvsa7Ltj7jk2TuNXa0wRaSi
acxOAfvNVao6kRDh0kZJyehmMsamCUWz49p39CjGpQmAq/P/8y/yZRGUvIfwlN5V
SMIX99cp4I7qi8gkIw+vJg==
`protect END_PROTECTED
