`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zbBk0gLgHSaD9C3c25+A1zlCks3rLcfigg1FTQg3Jx3a1QRwkixBJAGYvxCjHnjP
lPUZF0jLJ+LSS9ZH9S19IzqVoaTJWtjhMyHFS7E47L5L6Ieq7t9YOWh5OktsOqzh
gLkvDkLoSwScLHe0+ndfsL2FUd2fqLJ11OTne3ftETITAPP1/iegCLtb3uTSDHuN
maaI4lJzpS55OxEKhp3Cs02bet4mW/dTQujRb/JD2WChZSNioXskxyD/mPKmXIxa
VFQ0JYu6S3I6E8SkGP4y9T1ctW7EfXGaCN/wk0fvE/gPMjHCZEn645V48RskB9tX
dcMV8viZTrfkYfpzKYm+kQ==
`protect END_PROTECTED
