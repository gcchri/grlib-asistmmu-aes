`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
78/HznHluGtgvDLApvU3xUDNqgjklCrufzkzpjLH7la3/day3bHQtXr3kysPQmN3
M6pLukKfiBFg2VK5YuLitcmfZHJxkyBUomlFUjiAXqMeWiKxy28t1+B4Bkq5K8A7
PDNI3f/EQL5wpb4QwqbnQQBCrjOX6MO48vMLxFUM9uZPraYzgaW1SmhbXRPU092n
cuY+Hvu/r/7Rb+2m9kEH//o2Lj+7INDQ+I+vCU/vdj27BOu1OPh0+GFYy7F6Xa2U
m+D+ghPnW9UXZjsxs58059p5BKCKBStFwiC0F6NFyl0Bf53zB2S+4cF0SfAeltNP
Ft9x1xFEN3tnwZAeEf0wPmYq9Eifmq+eZJVfDZ6Ql5bH6ugtW63m+U3w7ZW3xzLf
Z7As5TSFJeS9AwvIXWYLbb6MT2l4jk/Z87weChou56VOQMebV6bulO9hdvdNmSZC
j0bBdctqwp7KuZEo1+cbjg==
`protect END_PROTECTED
