`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0MTv4J0HZtyF4ckwn4buhLWXtvoET5ZmUjsXe73CBoioHQk//DhKj6jIWG+q9CtR
8qN5yvWYvg6uj8RJgqzEg8CthN3q5eqa8CrqguvdNY9i2hYLiYGeop0yo8kCe2TT
CJE6rL6vikzodjULWKARmXU5t8IEdDST/u179yxCjTE3edVjfM+Oh9VETHmCeGl8
s48lROvnH/ISJ+L2i6BM3rlRws6q4HGcjJXM9HqFh75ilP6OPV4/xcVF64Qd1LhI
OqyhR5ksXH+gf1ZOnAtghV/RHCVRzc2di0Q80gjvE3bhEyZ5XzvW86wOEjm0zoSw
7SRPVh6e6ewwKnWwHoDzA+yCixtxAC3cg1FsNWJFc0cRqwN9ulsokznWU0YOqxKK
fSH+3z3Akon4TtOizMBwbGAVb1AOly8exiu6srmGmBGItID9Jnmmsx/mFvz3uiNr
521UqIW2INklPle/B5tPKfyMRz/UdyijoSVgt9v9dt//3cxWm/+4wPTMps0rztF6
5BBazuifRz0mDw6YDS9iPlqh3EDBtlcyjoZsG+6ssK6TgnHd0lVWjah9eTpSdN3c
x1iVCBkl8tVbX9zIgdP3dUZl3BpEzUtaWBRBlKwZHMgLJ0rFTxKoaIHD/NHVu4L/
IBlVj9lJn+TrSz/YQSl2FUnlCyNVDR7yFkq5Gd3D5EDXVjecVT+r2ZXAEP3vLSsY
LTkhq8/s9YrZ89c0nmhSpvCdSM0JLyQaAJI/CTMmbrc=
`protect END_PROTECTED
