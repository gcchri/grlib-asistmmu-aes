`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zHf1T6txZtGF+mjcKf1JLmHVN/e3qzsxrb9HtXNbUX5510Kjw0EsVV8lzK+3iSc1
YyXa8s8oUyiBXPfAw/3glAfN0Wyj5rRtbUc6jlLhbFNQ8MV2PBUmiT+f62SDQtdY
P8NK7A6Jxv2XlaGtS66rU1uzwuoiOsB58fAURNhP6JvnT3EH6ho/dEV6FmitJ6u4
/5AZCsd1C4pSQQvc4zOz813jadj1l9zGLpsMKbVm4pdcjnLTWckWF0DoCIzGi+k/
W/8kBQvtC92N5RiqJjk2zRKP6NjC+UJPKomjDHAnirFdD7FuVq+S9Lr3gfEA+PQ9
I1BGM3YDkT48qh9IakkRZCT36eX2vuIGFUvjCTdwncyK8VoePiKg9AM8VIPMhqaW
LwObMdpL2t/flMaAasspjsZB+cPefgsJSQ3NLjyQgPrmeqQ2LoGXpCQXUsO5aHsH
X4RPs+qev+hRbk3mHlC2aySbQNbH6XyKS8ESxprWTAlpiqoPNx5MzTZKKTlkPLMC
yLiAd9Mt9Nj+f4JNgS4OigIrsk5/BVAwwsR7X9rF4P8I0sVOkoWkjHYnvlEdflq7
Nrx0qCOJLuFKZN7Jjldy9g==
`protect END_PROTECTED
