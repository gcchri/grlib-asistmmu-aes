`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2QolvelYFk48ooJTYOBIFeNXe1KpIIDvqSQ/SXE/5XnbmZiaD93ovJQG5AVdvf4f
qBqkUl33ndEu1f2BVpwfhH3MZHcgpGmwlhTS7+jI6RQMSKO4Ntrs6MVh28kI/jBC
ZVFhK7aZhaySdH4iBRXY3GEP8xetEQs0WlxpsaJHU11XMxH+SvAwJSCT6QokEV/Y
iath0fftmavuIPnv4/LBfN9Q7b40VhT85ZP3Kvjz6Mr0S72FeLLlYGve1Natk/qq
fMjQQEq3c336gvzgX7FtrXbtungjGOsaJpPKY3BavyjB4XnKt8G/7QnGjwISUeLX
i8is1l5Cro23t5tRoyqVGuu2qHSyJYQRFqW2KFn5yyWsWocAr8mWWFbw36fBJsLQ
RjIvv0tYKI5DLDqvjnvrZJ9EG8hOplgXf4agMYfWdzbiJAsycp0e2vOKiHlRBH/o
ZI4HTCsG1XJIjqfWW8cNoBqTNJUYgyjVUj7cbdkq3My0NT03L5yxgoVRUFcvu9tQ
6qlJ0TZmYc8XD0xhIvMIQ1No5/kALS+IJqws5p2CWSWgPFBvi6B2RDiqBX/p7TnE
+qoS39yKJeBnsXVBSM/nQbEQm5gf/P9VUPtVhpMWH1yIrPJp2fYdX7q5kHr+qksO
VfOcKep7uG3Pv9bvXxo1hJ3iSykxiGFLcDkX3ddcQfTWslxFpwXhcsxeId5qdqWQ
nkwCtDsTeGKihs146YoxNlW1eDfLMEzn5Q1rkvc3Z5vVcLvVpF0fU+tJkjFrhD1d
`protect END_PROTECTED
