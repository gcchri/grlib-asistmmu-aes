`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AvbLcRHtcpCjZzsN6eg7kwIQfB//pL1H3o5HNN0274wEJyEZha7LAvknyl3lsdXi
BjiU4AtEyKlJR1QWJLkOrXo7LtLnPl4ERxncamtkunVgZqNdqfCqVmQIjieElxka
gmgDlYdfNTZwcpevPYUZ1My9u4p2z+a+/Tm25ssYYFVZZJn7pZABmJ9sKPrDcsXz
UPm1QQe4uiCE2Qp+NWYuJKJgwoWzgMYgBkpq6zLNTEBKw8XX6cBzdNwYsLp28197
3YTkDa+p7/ZFhVnj9jN9C6CQqu5CP02vkb3dovurK4hgX3//tOO5Nj+q3NByN791
ZtwUUpAJ5tiguyCGxgUJnoAgN9saxgBuvJqBNQiAThdghOcS57qExNGQRX90Tnl+
PvXYUbWgglU+tLmcVobx+XyMgRQwplO2VpJAhGIZn9QD98EEVPFoXmntgkh50lvH
IAymHoIeFYZCJXIUocsicKBGqONvYswTgW3jsZebYP/J0t2slDoEmwk+3RrGbquJ
Gzuv5oFf2juvTChC8BzF8YFKvm7Vrc4zY+IVIFfn6ooSBlEdDc3FDc3vpR/sinQA
acXZ0Ag+vE44THaRnTJwaujnXZXaDI+/CA6Su/Deo8nqzfDGCZR1bn602Ayslo+2
ZBBGpYEODejQOnPnQNC/7C0KstJNcR5POlCPb9/2w7PxVe3zChIVUS+vqAEvuoqH
/OxTdtWjTqnSo24meMgOw7gykZoq7FUvrY1q60EJUlm8QcVMhV7OsM9P7j4GZvd1
vAsUFvSMDDsF1jCwjtunag==
`protect END_PROTECTED
