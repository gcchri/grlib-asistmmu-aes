`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mWebeIkifGUfbH/lIcgy6TeD6ZyaoxEo5042zmAQIvVu4Chc00TK3JBM8HYJmGqe
sn8EJnVsjDhlWSr3Y7YS1oF1rG7cNdsEri5easUQA/6deQ/N6sMJfOkg152vCj18
V+TSnrEMPiaxYpJxxlFCXABxaJjQVpVWZpNHhd2X5ZmG0QjzZaEGmgY50XDkJEvq
ChPu9/SEVtzdYektv+ipGEa5JfwlR4SwFIYXlT30hLakbRWSKfZGiEP3LqQLhJoT
8yTayYGDs5N1bagA2r3YCY94oQzbBY4OnAEfqjj8j9nIwNtDHpk/EBJghsbwL8zQ
H2u/45O6PbHwh0mF7iiXWLyt+mFB+6gfw5yBCulZLyMAmD6U2HjfQ2KIHxGnWCwp
R09D5pfaqKOKLw1w5Jm9OUwbFJaJ/wNLzF5HN8kj4ejz0O9slU5y0kYIz3dJ1fEv
SJj+KCXEDkX6TDPkC90NW2WmOCspgq+pjaUJaJLlDQi8DV+bJhmLP/XS+M39lY5c
0b/b5nQUlyVFyzRSajW/Gzjm2oMZ28fih2OLB9WxtD3z+oSRcX0LaXkf0RtHBSPR
jhqhEcqmViRR08LSCmx+Vf3NLA/F9sTg+x1P5NsyfNQ=
`protect END_PROTECTED
