`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
veWz6b5dkvGm7hSjMZqypxIPvRlbQDK3tOyr4yw+oweCjYRvV2iJJyx6BSofn3m/
x02avVKyof48J79yzVxKw7IGXpg7yIALJWSymAfITIAwHb09Hxh291MyJkXdLVZV
Y3rvNIqJQXdSZRl1a/dOvXg2ISv9I3UVdl5gAKqQHpk/KV6m3nkFyBGSj2umL+yt
T7vectf6V2qYvvCsA3vxlskcYwa+7vQ6rbylPFvF/doMwXiUiYCeEYWXxIOvD41f
hGS1KMg45a1zxSuMovhuRYJB4MnRGTpFqJ9rIHPUdmmozeYNBhnvtDrNXu53tbFG
HJjT99bi1sY+L22EYU1bnA9pcPN7gecCyIaOhOoqb6H3+uRkm3nR40xsRk8QyJdJ
7BuNxDMTDTEcpbrnyCgucodJomM1t/6lrJt+M1jVodHHjoP75bxOkOk1x6dTDc2g
ktNrkmDPlaYrHltJR1lpK7NTeGq1OWXAuRNy09UZgeaEYFCiUpy9/9YfDbixY5ph
hOSQAFOX5z/yOrpxNSm+YrXG1Be0gPVfH9YhO7X3v/JpeLDrVsxdamfjYux7xCDn
UDhfQOLMTBR6J605zx8T3cYumoNrqNvGAObnb7Iz670=
`protect END_PROTECTED
