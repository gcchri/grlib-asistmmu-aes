`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6vLcynrrUZONM1O4tr4YE+rI3xSwFhjW2/9u0d3n1aFR2YobIAGn14x1I/5RZkvv
I0JSdUaIxWqGz//NWha8HrMDLbdJnMLc53I79rYr9wmU/TvYZMYy20eI73gxyAzc
GKXJIK1A9BvEo33j0hUdDXf2QPPhdHMmIF7vtBp/t0LIkB6aFH+ciPKYMkELCN7U
kdMQ9jF8p5ISv4HbyJD2qI5DWA+89sh+JLWWjqqViLFviN3ByVXaTgFL3HKrEYrp
g03jMKkhx/YUGRttyB4FHDgzTLqH60lmtaYR3zqU+H8ZUdz18NYD0sl9PJU+YHAy
fytO2Yo75G82Uw2XKi8Bc8FYAqwydHJo9o7okDr6qHegV4abiODZf8cdkGEmKWlK
x25GEwr3XWzdLCDpSbDw5zeDO3ygCSRjiLKacmKGA/HwqPZeMpo+Vxk0BDZdnmBo
JjDHpoWsIHcQ5p7wGBG6sAgOq07VT5gzRhrgh3yqnbW7bMJ7ygdH7ZQRgk9yZwpK
dVQJsKWuIvuVv0fK9aphdG6ElOzXqzyIhX9Ggo/Z/DVL6XJOiSBEfoSao5aaUX6r
XDAqA4wtLJ3Mz/SH9GvPxze6asVkmwiE0y70dwpnZnhJmMG8aBMxl6r/GBH0JJhq
08xP3cYAZzTfEVs5IcRDukeekPsXsjg6GDYNMyNgHpyl0VXgkccexmMtloW1bo+a
oJwxr+0p3MXE/p0X1/Gb0/5/hOJpahc7D8r033LAlak+KlpKA6N9uKsOOUbzCqyz
i7EytXfpaAMzUAI17yYHBBwC7G1vTZG2oYHDkWvUm9wJpPkbSgN/ltSiGOhq+gCU
FODPqjCdtcfGz3ZdL6NoUDqiJcDFcNYpacahFAXUwfAGHGUoZLva7p4wuyX+1dBi
5rqvxDRMFLbQ5UsPZ5Q6uLd3m1FfVyTQiruGRqXhkft8Wu//QpAjkzIMjeLeygJG
ZHHSB/o1GH7M7EYXiy9dmfEJlgT2F6nXh9M7uAxGi5cnKjVVfqPpibj+Qhp8uLSL
3HiQkPWP0z0gxlYV4yiD7k5nBg/bAjVNhenn+eN/Xgl0YkVgW8ddwLU3uwnQS3o8
tGAjmCZwRXOuNo23O23QeKEhb2+jFI6mSnwCb3d2ftqs8jxNuR7zu0ZuxW3KuhgU
1bRb1mfHLqAqFAMWWMECgAcLEfAkO+bqIPWIfg1hvHpVVv4jiIIUUtMeMq2uHu/o
bYDUJ7ZBdTIJ/AUxGyNXZqdUH/KjxAcOMDj2cGsAE5DRTEXEMjBSA2bUKJ0n5BC7
lLOTwJQWP7NWKN0bOZKyq7SHqg9IG8tcaHzU+9SId/q0a8sCRKccZbj7wv8xrwAZ
H+9YqiYx4U//VHAe/NacDRxjgxch7JUWyVrOhrvtfVP2sVh/V0CF5CzaaEH51usC
6ESYf3pt/ekkNSpPhrPs0XMVlrgt1GEaWkF3RThVu6mOAHt0CXscVwcCxP7qVFZD
JtJyE1AuZ6wj9jxed4vW7kcm7OwMfa8yU6AdJYkB4bJh+8UWmGP2HkCIKvWjfHys
1TGkUwVis/UtrjCTo7Hwm2MNor++bIkvH3+xGsVNB0tNY5DWtm50h+VPUSruk6hp
y6kfCSqZfqgKDUnIK3M6SGf3yM0RpSUBksIbWWPH/PM0tiJj8n/hCQYTW2vCrrYk
8s1LGkowXE+OyEvJCe640E+WIH7ALEviLC7NUvQIBdDLtyO2cRcCFI1xQ04Vsqqb
5cnEyi4sjFrqsawk+7NtnoKODSYFM4yzf/+FPgpVhhL1PjbLxc5I+/mqKCtYmOWH
PxE+BT2g+YdUTDLjhX97b0WLdRotbx+fVWeoxSBmehMuWwBBULtS34QWy18vLg+E
aS5ShG0NFOCe6oqtQO64ws/s+0FQWahdHKwrmt7uZDe5p6fHCFZj+XFmg9I8N7oa
tNJEvFAp8/TVekm13UhlEv7pVvovRiXTVxRZPI04TP3FKNQufnAeq6sfeOTFTh4z
CEqJUgxhiLbhWQh54i2zfzTdCM6sF0eVY2MkIJUZfgbeQvsr0JpQYvqQHTGSTFux
IhPLN//aQN7oL2LaRJCbZV7rMGH58VeOYjQdia156YeirbMA1J0lJMeN8KyRAHQG
h2qNifcVxsAtjip0uVyz2LxBsdNDSKQuVykUfpdehqJ4RNPhlmO1xbVf/ZNr/xQV
iQHX09qjT+iCqx8xGtjlHOfyMQw7+rwG4msuy6MPr1yhuL4kp1AVmt1DAz953Ap/
S9qvILLqCClTKwfJXvPQlUqy+m3vkT3uPl0Tk+GJlseG4iZlgWR/WNrXeywuOagr
Kt2rsUqH64IklZ++3+ecO+aQrFdUIUIFpgJLgZqSokxtUpdQOc7eEp6rTt9HRCiX
KV00znlge84Fux/BAo9ohYngbg3Tc4Uil/Y6GME0EQaevx3Rs87T73c1Mi/qfqVS
zbFVM4gRdXloH+M3cfd1oB3Z3XG6JOPHPYgQ6rQdTqtWetDuELJeTRHvM8K8DOho
gKna2QtSFLYWKsHeiJZncLkbnAi3wTBM7Ja1oOv1JmG5r/Cf6BWzwDiplo4SeUQI
OGlMknlz7aMdx7F1uZN2mZ+58hdpWq/p8HurUh1tu51GMjNiyKIusr18UmOMtzv+
cGEUvG0J1KthDxzXS/sIDLPzRy1ejXWQHx8JLpBXyrLNUqTAAnr71+F7cD0lXw/c
FWKrB0e8yegoveTeJyI+Va23RSeSwVYBfy8MzI6l52HZ63kW2tCGdt5hz/Rw5V3W
5w0Kxt0aHMVaVRbLinmQ+uA8kkVKJnJ1XNqIEPwFqizsaQbg/wYeq5iAWb/ObhMj
sUpCZKGuNsIhW7XTbQAYbmh9a74jCQxvjd5wO7mvz7djIbJVn2qJiHxyKj9OCmSt
pfIFEPuZZCtg2D6pUpUW89MfuoBvVFsll7jw7FTcXmYGNqZvRxcFnUkX2Kl09Hnx
TR7eoe/AK8iCP0OtbqeBDAH7urv9vHh64bErli9XeqiVPC01yfIR+jDHUz62R8Vh
1H6lFk497hJlQ/Rx371Tc/SBFeKghk8qa3+1UpVQuurid9O5nLx9gEoNOnEBJIQX
DqbkrSd9IHHw72N2R8VnR2r7OZzbj/v9dbtyebQRqONXPVkOu21VMmlfRP0BGUAh
OdPM+gU5UL55IAdBXQDaZrDqV9+iZ+KbcCrj48VUCAECnq5DRadQOe5mnu7WsxS+
+7Ay3Nkk3YuEfR7fvDaR9TsEjpyOZaJ9PuC+xaVTR0C+Nhq3q7ZJHmOy1ClE4tm/
qy20fU0eVP9o/MsvneQ2zHkFNS5gunoSAmGX5OiLGPFyTm6c56h/feFLQ8yYcihU
gbGDqx9cr6KQljjTTt7yh67VWaXdC+0Hke7NLMJoWnVHHqASu9/I4I5SHYcj4X8J
/Xqtja4F7JLsigOEUW1d5AsA31A3yOVHjDPf37qETowRstDp5gqo7z0Ly8I0QpbE
2KkaxwRn/IvCIWWXXYhuft9KTP24gPKoqDg3MKrGOJHX4a614VDnLS8QLe7zhoYk
CImjeZ1RxPL0AYUAfgI8Z5APFZXbq2Yi9g3QTflQygqlLgKGSri00ufkxKmVUUTH
tLDf/FkuD0WxcIfrVQW/MMZk8C3Knl3G1JD4PkRFb06hAKtvbWZCh5BDLMO8S1T7
VDalpVJl/E8eQTTz6lMNszuMfIoGCHYSKFJrJabVp5lbzZffpFrAT2NDQ3mFbi8P
LJedYG3mSECbm/hG2PdIyCkw3fFN5ZOqavko4ElDOCXikL1OByVbPq28bGmJJoJi
g7zRkx17RCbd3w3B+LEtFgNoTFJK6FMiFaWIx3z727+TKX/N+G7D4qbuFHfsTD1z
00R9h2H3Kylg6VrplggfWWKaWPX8NAIvZCZFzEKIzdswS/MyTsz8bdAx/pqfL48T
03Q2ENpUfJNya6iaCSI80PDHP8ZRPtKT2t4ysYDsJcs2LaQRONFAQf+SNSsePmM/
VxZ3WeDV4Gf1RM/QnQ/oCLZ0FTmcWS1we78ETuJMtjHuqMLXUEkHW2Vq+dHWI0uW
mnXkUUrzfw3dMaD1l9mSobg8l2hFPEZj/TMKomMSDePajW6nrLQ1RxWv6Ya56GeC
LxdCqFbam57AJG9Yzy0mDN7yiU5nPu7Hm3/DBqBMABKBS052yI/hVZpGjRM85DZF
jYWmbx+dOxY+JarRSYPvX+zEZkyAMxLCZRU9I2Kv6bYOjpycfY7F0qzQXuvW1OZ1
vtBBVKK1CKS4mIQ6J8YE5fMr+PDjpsUPFlLgHwklbWol5BV0lo/jgm/rx/85eEDK
ZuwPMC9MLqF9shyAzYRwkgWIJlTVySjLPhE9ouUonjE8w9WfX7KQe+HqqFiyUh0R
sTpvoFa1cXiDgc5vPjF66JSZm7mDSW+RSRi6WoDEa0GxaWZ/CJijL8ZiqqnZt8l1
QV/JF14pTjnilIfNjLK6qPvlnaYDNURS0pu4AViTplAfY4Lm6qQ7IXOmufDiAzse
L7wIRedQmLglvEhchOcoIJduXE4Gmsg5EuH42d6yfSNjxDSCFYaWKPTsyS0xvr6U
XMSZ0biaKGOi5S2vA498IfRxjnYeCdzRAR4y3G8aNc6q92cSt1BbeGmf7sofM4xR
85f5HOnasuGpEUrZ74zQeRPpGNp+FEiVqmT2zLhEdE+BtxojioSC3t7OiBThat3I
210AUZmJLpCxlHVy5ZPgQLLap85CdAVrjQmEvIjAo+3LuyDFB9fTXyMLIgD1hKwm
cMIhZ7aukPHVLv7EPjBhdUhgg9D/ANAoQOOyHqbvj8atMeOABRA+zXmaSP+19evq
OqIOdl0fCGugHu40bipUge8XmZegbLxym3cDWnLaLhv/nAgJcIAuuYN+EzmhZjFb
xOMGzMlVmUGaRLg3jelq6Wen9ptezlxweiz8cRUFxF5rXoiq5lAClgeit2B0LqJr
9VCVkZx7ZrppRBM6dlsk/8yrLI/8iQLrb53tDyHeeODXC29kPsqv1XQ+ISrBWT1i
wrW+FvVp3aP7kWXj7dHQNSBW1r+Mx0fFyE3NatCje6k1rPvjZAjnAFPPRvMGOOv+
GRHVV5QhI2y7oEOqmzM1CsffbQHVP+FK5ih6q/2TCbaZb1Vua6mvMDBp54/QCGi/
Kxwlwdi6VGWfeG7of0LoZLK5RKWNXJ61EvAI5uyEsSxcWMjvVJZmKPxZj3T8Ymtx
v1UIzMSiwLgqYDUqXOQLyWJQgHSAxe/SrKz8Bdxz2QGWOQbo/jQUJJZC6Mg2Oy8k
45/vmgHfo5OST0+2T0wf7jWjgn9yA6zCOuixeRCRuKLzOJZY2BrKShXXPOb4uZlp
rzkx0HqQmWrrOFbO+9gK788loTL8lbwiRV9IPRQDfaQMScSeCnSIrIO4T7+cjd4M
NP88WuGaKZdcNbFDF8MIIHrAwtWvHlV4rfLg5qdeYY1eya3GJW0rpCOb2UlGiCLb
ZUNcFFbTGsTsPeLIXbSCrGPZRHz8/pxAOFU/h831aDE0/9F+TJLcDRL5BRP5xdiZ
3ShV3YWtjF9uH0xYzLscXX0QCNSAIlnKbN28jXr/juvx3+xFnFWYSvSpOgOvCM3j
7At98QNbKSkIUikGt7CUZp8269sBHvt9dnXcOCj8PjP2fKGc/zjiZWCMCjQZzX8F
K2A1rWKsmL4+XJiSHwvxnck5ohssFv2+YX0n6K3IVvPJ8aJHkJRtUuOJOVlLzQ5E
vvZESXsYIHwRM3rCGKBJu71SS0E3X5yBXHB2t1uHGGCB13IDh8rP27fUlML3X3rt
5R6RvPgmylz/9SVxY++Tdms/e9MD6Cry9m9yGLD977wcuU0K779uUZPZ6bOFvHi0
gx+58kFrpFxqZsCYHJxlbvul+19kGiGMgtA5Zivtz+uaoOD8MnKSkTid7VfQUKNL
VgXNGgDbHw1yiR+NHhkuWqQTcHEqtnzmSXaUD3RSKjVqqM+oOUBoQWuG2SPTKIxc
cO88QU9Cg4pTEypoR0FJBIha/sTouyBc/JH7ktl/6zLKxuPpPvi/NdoK7b974pnF
zPXU0tHphZ3O6+zaSBHzruqDleJdBlHWGNAIG0t6gDFTfmtvxpNckpcmZscmH9uM
fCDtwY11wgncaJgzioXWH6lhSTc1HOTpEtK3yvU3UNUQHUP3yO+qsjOt5t8gV0ej
pC5+uUAtXuCKq/sQrpJU2876tvlczwVUZGcDSmIO5kcpwJLRbRqRk22xW+AnsAtC
FlqoMFVZRJgpR5np76kcvIKSNFIxkQp1XEmBYbPoIpAto64aJHZ/QWBYRoZTID7p
r3zT7yWCNVTIrIQuvHzpTxsp3kXmtq8F2V4FlC0IwIWGNLr33LaYOaT1OBf5nbWK
+VOCkhtZSWDeHaBI3jY6qgi98CATsZAnCUmK9u1TqFMu1vJOTVm7MSb1+/wQNIDJ
CTgBzQWcjAOSNjeNhsNAIS9hqcDjVtfrB6MufvJRABphWRtbdtQ/GNhFL2Exe3hC
ODix+C3NBl2OoY9mvSSqKuSSf8OEMt+XbTp8UyzGp/7w/WBRJPWVR0P5jjeR4Yhc
+JTEy0nFI7o34k0zu7LncOpWCxf5FM8Iq7Gf8iIiZGGv7Dj45QlMikXgs7m4VctN
hfmJB5bDB6gvqev/pWofTH1ogoc/poQfbq1aIBKw0TbeF9CYvLSt2pcH5C8Wed6u
GT/as0Hp0UtZidt8dmcKayZtb18Xv7KwlUl6IIbgiAwRZ8nDfGPPbLJdUtvxaCx3
GDgkbWtcQEyvpi6BrOC+7QOMM/esaPdOBtv4YydyIbJTjzYIo4HlyRsbVcWY/TyF
HTPOyRcxDEzKv6to+2SBrzJT4ApCUSZrOfSojThnKDUBzHYEv9/yTYHJyKNKZn12
Fld/X1gO86qxqdSYDIVuK2CjhVUiVdjFwnk1thjbrWhSeP8TVp5kIym8suraqVYy
6FqafSaBKlvRFErJ7zHETUl4ifokC4etfjw3IACJ7Bm4eyfyKTN8pmw8f4YZqScc
`protect END_PROTECTED
