`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QrX6pAr2lV0ukdh1+AIN/eDHP9uG7ISkMVRkbJ+hBejVKuF82FELs2yZH9JZ20Yn
bc7xgASnO24EUm2iqdLNok7YoL0T401XJlp/ccZD/ZRJVPCPjHNBeZ0xX0sK6mFn
8U6xS0ZrEt0pKIGCeTftDEChet8S+hxpBEDbqTCzc2WzcdrD6Xrk44ZVLeU78rlX
6jAWwpKPBbSAHwL64JLIrcIbQhV3QmYW9543vPrfHHAyDwnLiJwIcD98JCC0aqpn
z2gdp5pcsm+lMgie7XNCXmkdnGKXJWnR1V9yJ+YpofxWXKlEITR3gGTtiCyjUP0n
W2ymyQ/B9y89eHPbJrWcmdMqhLYZG9xb8s8e+gQN7uGE5B10+y+0jfvH4gf29iar
jZ1tKGB6FdGEoK310DfWg1f+PuWEBwoI6axIodgeS0dswKgos2uJ4ta4R3T79xtM
l3eVvwzwjFWEkwdX6sIsvngEQtsbAIsdThNgCJGMRK4NzK+pp3JCPX5w6ACf105a
/1reyJWED4jmEx8djs4ptwHncZl28O+tIY7Sw+iI7bYE5jbAPguv8Yu09f7rVIR2
MrYlXi3ggraEleVN+PpDB9QNtKQ5liqaLeDqCMxy72lwcAAzxZGe75E0puERLMlk
2S1xMLLmIFusReWcDyCNKH1Z3GVxW2JQtMZMvy8Z0usKlk63FU72PlE3sBYZQ2X/
NAH+gc5W466ZxG+53scSwTH0IVINSqIqX2YTyKZozpp3+Drf929om+fJN6HcKwVD
a48SDFFFybY4uG7GU88UBuTZoz7CdEYRnmueA98ghcHitM7P5sTZgZpguTMNcqaD
Xz56nhekO5oxqa/8ph0gmOxDgzMavvbMuZ/2m1KLdrGOE/3edmcY4/9dbsOFDaut
c/suwlLOmMuj8K+i+3HtDb80SFQUrkb+x3oJzRsMWu9ra3T9U/7K7OnYF18oC9Qv
1jRjABT4FhtQULfiXnQRptVB9FLRw+gmVE1Qe/1Q4I4qbzxxmiMKWsCri0MYoX88
He6vxs23G2fyKZbENm9DXo8nSmWW7bJipB757gIKnXO1PZEyg7nwH0Va7LfLLHfD
A9n6ua3vNgEk4NQr3j8hfUlKG9jdjP/16q3J2SuI55NjY92WSPqu+LEICi4DZ7lp
+GN3Od8pZjZAy542n0JMFbzVuPaBfP+6i2x2Zm5FBUYmeCzaoBJ6z6xiJqvIacpk
OK3/vxlupsSa5jWeREqldJwzKzGvwwU2zwfbZZRYOrG7c5GUabLMZn43MecZnkF1
xqFaB+PYMCTZxa0OclGSHSVimufEq3lxAG3/+U4P1YkTRAnsYXRU+3GWZ5liKeze
xvbC8JR4UXfreze+s8QUQOBS/kcjonEiJd3QrfyPJ57S8o9PUw39ecp16wW3LEW4
fgm9Y7zxILATQHF34Ge8/emRMCvrcSurAKffy+KvX501J+a1r25loKzGaA+YW5aD
RF6BRJ7Wi2gU3T2SJMD45OQiVru+OWTKXV7syy7yIsRvuiIL/JLHH5Nd1kj3t+CA
SG7dIZHBixQfznQ2lDKGN4JKP3C3LE87ucM7aNpzGhv6mXO/EuM333SYWIlzARRB
jv38/9FsJrvmNg5rjL99lY0h77q/muyXqW9LIBlF7evR6TlR7X3w97W3UKjeH8Bx
9nN12wCS/jI8MIy2mDIwNfGuIX/PVPyqQKQEOk0BXV2FpXp2NGgC/usdoJysIhoC
nZqpln2XVA+2LAf8/DGmxE9ySzfAI7bVzd1xZ2xkcJA5hNX9tYlmSV4p+0DMMl8t
5j+lgwVl7PXJpn2XVQWEga55sbMvGil24I5RoIsKvhZ2cKzO4/SbZ86X7jM6XFvh
RaBxx/zOAomHzqt4eKpB5Wv8TX71eGkxRf20RlBw3z1GSCZndo/DKZtmnav2Y+oT
kpMbItCkgPHSzq5ZgTr7dMUCma6cb4WAJ9SZcGQCulthCL3fh4/NHEs3KWlNoP5N
T9c91xXyCZYYTTh6HA1kPPeoyWZHJlfHoyEvgkUxsVtiX3JdvFADRAOJSSQfGv7c
JDesH+PmBY1t7LF9b3dKSaHDeoxyowVVhKNIurSuSwpJ0ipd3KMw9xKgsJaDv3wZ
sn19PaToRDOPlAnhs8aHCJ939CcPXM1taZn5mT6zjOnxPHlDYrac45pQQp+zUT9o
3HzgGGPq3l7EWf3zb9Oc6G6qBEfnud81+hYtaIKDMFNNPpwhfudaZuJecepSXJ2x
6hc27jZRJwzXWRNZdqb52dpCP5HGfaUkd36cJWjo6RJP+/YKMVwdfpawoYHgszBh
TX8gBIZ2MeJkcEAgVKb6/jUooXfjowP4ckcUmOItM55C8m4pTG/ZlJKs/nUjtPpy
fpqW8A0iC6pkVegYCfCYt7JJDV/sh1WxkwsClCtPulCMSWq0r655s/g1R2U+WPSL
mrzEdQCKjdN98w23gzpu1wgz9lvUIxBHInlnaCyGSDzw65MDQUiUcMdkW23pYSc9
86qkCy+ilWA4fkt9mSt265TPd/vS4raUw8wNLJ/YVc2d6t0/XW26JGUd0kxAGFr9
wizVsXFvUvm6aGBFzxgUXh1lwaFx4aTc/rlRxXjY3emMhYOL968iE1Ppfhz4HlY6
9p+rnrkdPE8kJcgC/wSElUh7M0dIyn5IJZ0yFA+G5fIdq8rlXRJ40aWn0f/d0btr
VILFlqFcEVMS4Cx5eRnr4X6ymp4KLPTEp+fUzKKzjzcEZ1PQePp5m/0ZL0RSpBJ4
xKjGtkRwAcSVYFu4PzOs/b6Su6glCmBJuBGnKkXiwUOGWQv8nF0Z+IOwld70HSow
b90kUSSDSBacAzvcK8qW+e9rwipXpRvv46lUmy0X94p6/Dtflu1Qc7VGMw9vum3T
ubrtegwkmiPwu18UhrDbYn3e4kXtvqTZiIdQkfa+gsNP+6AV+BPVRU5nBk7r3Eox
gb4qcoqdPqMxzdQfXrr39t4/YaLupp4GotDtzsfhoOWxR6ewZWNHgwoZo4HohGZH
9TjnXvpCHyMIQWnL4wPZDMBO+FRnKHv28IqhOMlFtOgZnQr7+JXlw1dSZCuYqXHx
D+HZIAiUyMAjUvB+2WFQFLXMYv3zLYL4LL6zlvv2sOuu09CRZcJzHABOu6wGFjJg
uZSNfgt6Z5e8KwSNHo3sU1eov8YTG5O4NE7etwgw8dhTbWEFFPv9OxhsoKUW/Rv6
BARgrlAlu4PVIbN/9rmM19q/3P/V8E0QvftHIDvQ137lA11v5ncM2+0hZxGaDMH2
FdrZIHtkdS97LcfQJCTRvad7tjThQnf2DwYATynAREXdXmIMEnQ7iRuMJxS7xxfS
rqZ6/YuOn/st8V+2KaWRI3Nn2tprqXJRxOwseK2u2zWnwkrnunxdefQRe0780h3N
YQlaX7UWUJEhZJK9X4OrpNkjGsp+N3ks/4oX8EmPsRm8eAOKwzq5doWv90Zd+wHH
JgIGbvAS/fI0TDBhXQSQathwO2+uNfZvNCXF7iG+jGcbi64VXqbJNBSAjoEFxzRg
I3SbGZmQDONJKrMzqFhHbTvAxYMEq5rr3ZrEChUTYBBsuiQrQInBrDBHWafBHJJy
MubqMBHtc4PG5hm/k6oKR25hAsyynO1PFXMXjH8keizriqu4CM/gbNM0DOYY4LrY
aOs/+o7bSxlwIlWEjDYMdRtEdFh5PmbVIl17OHvd3gOgsAWnAaUDw+6/nAhdeCB1
LQpLgZEGsXy+t3vXkfRdSpKeTs4Xnb2J2Q8zHcAJ9u+rqw7HWThAZWAHyfZA3fzz
W5Ubl16Vssc13+6cnyLZ5DwEqyIl2aVN74L0VmfQOyAKJbSWi+PEbdnVU1Jau5vd
zWY9pNsXvkXeYklKA6Zy590ZLinSIcVBHpg0wCcvrUnYfnI1Itm3yoBQBFN79Tps
yFWFgdUJsL21kEUU4RDsdcr6AmZaxLHsvrlSp1bF0ORDIZazgqurHC+oQ/HR0ZPE
B9G9WeV/Hih1No9rBVpLcpTIaT2u5lAA5EqcQSteTz96r5sfszcCqmTj9VZVRtTn
CZkzT3SfUmtCPYrqyIvdPrEdk7pUgPaRS2gmBj3y20hKrlpGQ5+eH3o5d85juyDv
XikVIjLuCo980s0fwYuCNEFUYbc1aw0U9js8wEABb1a0vvrctXzbyW4WU0kERtLm
JT56QBmSikwSO3FJErigybq5KeMMl4igK1MWe1+y7d1CuOIMM/U83ABh3iQNWta3
wAOuO1iWzCQpH4fFPkiyFYqZY7SF5F/M07VnM1/H+Ud/Q6IXKYxWUt0qtGXZsjUa
BjYNk/BQpVHM4Y6n3f5K25kqcS6CWq3XEnnRzeV1lkWO7MwUQKU/PQytzSYXw/O9
9H3b0lDCW3mIFNcuAhoqmvbaB6Xu80YHlKr4+/2aTrGXyPEAzquxwaBpd6QicJYe
BDZUsvKGfGueUoLBrxa6K379/YLsg/v+5hqe8pod29K6lalgSLZnk87JcajmrQGj
g5MZpGQG5cwt+CbMQFalJRyIxv0EAAkEe2hkcck10C0j4wGSoThJgwR/WxIma70F
vuvHillxkYukxKmOUfKmGxavTghqIJPTVbbKhixnNbZMIfUk0gNl52iE/mV1W8Td
wsuEYOUhdab3pw3nO37QKtXrN9UUrF74U0hEzkWaIFaYdUHS1+G0BPuRmGnGkRs1
NmWdZn3As1vMiKkajyARfjORZcWfQEEGG08mesRE2VfwvCIbkdA5DJvYUrW+eAiT
Scu6NtbqY9t7DiCojXt1J+Owh5QFJattOWd7fk5v6ilbDd+C+nQ1yH6d6u7v8Jey
srV5pCCKBU36VlGRZLjqs/x40F3MvWbPCP/ITHAEewFcSlalGoLif56eZFR83Vt6
n8/LjkIYM9AGByBC/8rTe9Rd37Ps2u6ATcetrzhtw5qFfPYMMo1P3/9TU/O7DipM
nNUI1cFEnz9Ni0re7NM0yQ4wOyNoOnyUOFZhBfSgjTSBmEuma1ODDiSt5bZIpewK
E5TlUldns7ZZZ6b4FFHhsPDyHJofXu65C+/OvdE67jIRCqzP3acx1+odo/ATY+ee
odP6FwneM6W76N3udH844Q==
`protect END_PROTECTED
