`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UhndqGNWx8bMgfKd78nNh2z2nEkGWFttEbjS/nVVV6BSmm6v1WbR/4+NTKa2XSfU
3Cd9R40HOhdrl+hzlWrgDEOOrZF+YwPiccJSy5l+o1PpLzeEKTeCbtft9L3Y1hay
JKEMQqIUnwVdd7ENL72gCTbTBIx2MfWhTdqZAin6dfml9hbKaWPo3aiLTP8kpid3
hioXflVUoJ6LQaMT9vNXvfzz58UboXBwJrPB128tPHgvtPgP7q5n6KpMfdCOR3EF
D9oaY37FeDOPg2A6/xkAHEsYstBdxgepL/kuvvhRmhq/FqACpCkURgBnXzaikn8C
TY8tcsJsLSaGfCCvHY3ei0P9oWxRQ0Q7bd27/INdqfA4yLdwE48nKvjBpt1H8Zzk
NdOiRzQyN1JxNkjqsUe62g==
`protect END_PROTECTED
