`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1u8A2iya8RFXeXlqpiIdhq1Q0wwScPK3OQ8plDArwdyZdYSMBOdZ5bHDrS7HYI3g
bDcU1fCrHRGGsHJ0ndDFx7RtSdjMLicBv6clj0BpRg43GYxmYi0Eo9+BDbC1Yj0h
M1A1OLFKVr11BdNQ80Aj0BQViAib+F5AmGAY15sEemRFtAObt6R4NQb9zVxDROCG
7J1gpfO3W0z+I0INDXN6y51TvLtLzbQ0w0wZDXEWIuHFI8tkaRSY08lPeonP56Qk
TJKhthLyajvJisvRnioq9LbmVcWfxx7rsSF1XpH98Uo5gfFNeVc9MVRbEL1YnvX5
`protect END_PROTECTED
