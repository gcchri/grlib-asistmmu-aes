`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HuvQo7O1Gv3hhKxfAhLDaX+l6h/BYjSSPK1yeo5RzFGOjtD1GMfdsXfDm4oggrB9
QYccC6dKx0wLDJL9vpifCOq5wytrHCQCgB4r7VPm8Hjj6O9IS+JrQEVvu1I2XCRY
S/aHzYmj7yJwJsWmkv6Y5park3or2Z1mG8pi6bzpWAT7sVg63H5EzFumKrtTAtdb
QfICFTb3F1v1UknqGfmL7+OsW2UatFoZxS+/MM1u5/ncufBfShUe8exdw59ELiRR
BivxAhgar+rYR5fmvJTKddRxH3xZjwzvf/ZnrKj47NKLB7cIKFsbJpqADT+QyQ1a
HfGqMWlrqSt4MhkLvWrfCA==
`protect END_PROTECTED
