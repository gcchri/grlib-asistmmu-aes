`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oJxP7D1OxHbC6EEUZN6vlwgVW/Tf1YmUrCblHhuDYtH2jeJEQfwio2cVR3mHK7yt
Vj95uYaZmDq5i+9HLE2gk/9YcQIQmd5n4bs6aXWSXu6j6gUL+gzLKioPGw4Pz4ki
3Xy0NXRm1sUMK7P3KFA78I665VJn2N/lyPpT+MLdQCm5zexw/3ewo4XAivsWCT2L
P2oHjkFk6N1cPZdDEevVtUHJ/OtNLwOxR8LoqM+BLHWrqoB2HluGypFR1qCRieaP
+3ZGNo818NJ6GPEQlo+AXWakiSofztEQGLeQE+5MP8xqnULJF1rU9HVPzjF5SfxJ
bD2nm1sogbbhgVU+yNC2iY3L1kFgV24jLw3ccHI4BHWCmW6MwOWkDayl0NAbqySl
dDRFLIHuvtFs/A9QLuhAbF/ONIhAs9ozypI9rgqc2JY1mgsUzM7OKvcfna31FSGE
92Qk6FpvDQ9dw5L3FL1BuvstcIkk4ETYRCR4YnRzV0g=
`protect END_PROTECTED
