`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PICzCZbRZyiOo2pGxEFqPYX0+6lkltbck4fwFAFgjS1chjn4pucDLJSz3ZaJiGFm
ZuVYYCvhFsUp38HSgOEM3C6mIVXTJ8vGlrS1T5tRHnS9ly9Yy9VgV6WzXeiKP1lX
8dq2Da/yP6YLZCiMKCIPZkcPn52vbL53ut4uc/3gTlR2VJbEMZC09/xNwYy5n4oe
C1+kwvhfe4FXHkU3Sjoo9aK9I5+huhGrD+JAn98JzuF8K5EWDetxiSYRBu5nUMer
l7GMyXCGlm2LVeilWLeXM6uPYu/EfHKaLuv0ORvhfAtLmW+mGh10eNZ0bcj7/D6c
ZgM2789CUS9UhcnQBypFj3yJSqnSUOh6f2nGLP57Lno=
`protect END_PROTECTED
