`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ulPSmkiHDUKwHf0e5UglO7iG9ntZ8+vI1ArardhUozuM1RAvDM37Eu1jBYvvKXOg
UDcq5v9E1wwQeeTWSKGGVswxAEzCRbLSn6U3X3gzq1yOjtyxRsiZgh0MdgPA6fB3
cQoajv4cxEcTJbcQBnOnX5V46NRYbF7sV+NviNgO/cqniGnprElrgoKL1+MQ+W6v
1yOK8v9Ch8LJ3KUJO3myFfcfXkJcN8Hqz6qHC35BZD0YEJ6bDJDENhGeodPhdW6Y
od4HDFbPHWIHnbcXz9qCr5ioom2gAVuJQxrtW5wEqIRakV6o/e1pFm+vQ7nQG+Rf
G/j70z7dpe7pTjvcd//rXx7WZyz8eFhKBbAdx1qoYkAVDvAOnAcHzm389SCJqUW8
je6px5thQs79Mr9LPjbTZESBiIaOqY/8SpLRFsg0dVnXRRGfcC8Yvl2lp+U3Vtph
`protect END_PROTECTED
