`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AJde/60nTFhFwhI3VgrxUfdKKd246dRkyKFu/CH4Eet8zCio49O+16x1lO+1pU6v
o760ol540B+vR6aBTOzL/0rMQ04SWercR9foxjgbwJB6xRnQXaEl62xNiuFDBz9Q
wDsqNV3ZmuvU581plXIFAV5IVK5/bEGEQ/PPCEFU5KKGv5q3fTvnJq3rBHcho+I7
nnE2CNOc7vn8ev0NwFRd3CNbP1eggtPWq3KyS5DXxf2KmniVCu5hjek9Q0TEXTSK
QKZSOlfG4HiYOPmwFaXDtrigNOE/9TlUsdoS1r9Wjy+7qDQqgRl9QfMvkoh82AiX
xAJUqTuYMt+8BY/JsaNSM//VcnJZZ3wiHY5j2XqMQh0YtgaiepAfHz2doPygwNVV
bNsIroH5oey6bIQEt3vFZT8PjZDs60p1nMStYXVUA/E=
`protect END_PROTECTED
