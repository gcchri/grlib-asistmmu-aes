`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MOspatQZGVdDOqNVaD2f4kUY9mgXWI8a7fTDTRxzPBFpWUk3StcFSpPzWTDB0JLk
uexRhuWI4wcm2lpgGoDYR5Kn+KJgr7NKBGlclR40EOYkf/7FUwzc2N3kj8uveKFU
f66fNaVftEb/zEw3X6QTweTsx+amXDYXLjBGi2tzFqfnl1DojpdqvPVWXiV1H6rd
idAkgpWawCPg2mFL01en6+UGIFaR59khy4JlrzqRuHsJwkjVU1gD50it1DURXIwZ
mfC4z8l3Y890YkkoZ3F2K+Xwg9zb9s5tqvZMBV2P/zfnGVkNKk+9r7VBXWd3i0PZ
QtFyThnEadMXcSLGWSbQgfkjv5IiXWjyNrCj7zXeg9bHu/0oBcjnInALqBE8uqs5
wOH/tn9ZKscKcX9Ts3DKKjitCSpTsM29TRUyo2DwgBSaLyekKpa76ngnyFLRw9Kz
zNd10KvfYNAIL7PbLQ1hpyUdMzzCMFlhmAVtJmMde0E1EG+J6wACJTLllog6mu8B
NR+7pTZ55WCUUYtCrhrhM57QZrf23pyIXdcHcUoPev5bOpQ37KAhEyXUIlzFYeqe
Mw06+2VbQ51Fhe3qaMdMgFpAB2z1wOthjATFH8sy0ZFiMjlWUV32Uqvke9Ha3E2l
cl5QGa63icbaAuq8RxRNlA==
`protect END_PROTECTED
