`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fK+cxK1I4V0yV3LRS+anTF5kyNJiE4Yx0rtWy8pV2A3d6w9c3gMD3XYxBgBwQYP8
TcPQ8EUKjGtrgkFNYuoukc0L9DMbGciPnf4ucdJvhwMDr9aTdHGvINzxAb1vdCzj
oQO332EsQszsq9e4lnP9OYRit+arC7AyeFf5jFbBV4SmXTzPAlYGNPySb4lslJSO
dVZAnh76232RwVNhY9s9Pgqk1FcgjmURBL1GDFIrz8itfMuEiiU6WCsPygIa9RTz
tlRKfFmxP7a9sl9i965mdRod3OyjmRgz9FUyBb5T14EXTXL+M/LTB+C1qIX5K9eK
kO488uPBIQkONevACARg+e2n27FwtsksbT9+6HlSjjbQx3XUYiVdLqgZb4arTr8w
AbuiXMpgnnem4/e8W6/+Rh9FKLuikJqrPxu/4CauF22dhHbFdQ89TIS/ladyo6GI
ufIHP9Tgte8BMiMCf7WAz7bdbWAoqQDMpVx+NU4sxP4Azi7nvhaQCXRz5qglwhe5
IBD8UjTHpWWzt43eimKuQD/ZRYhyN2BHngdp5Fvd2gw=
`protect END_PROTECTED
