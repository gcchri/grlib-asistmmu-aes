`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mGUJw1FlSm985KhhZ9v0Z+yflnqjPH8NwhO+ld4xWDWO9Ira3cNNmCxJ3f9zAt+I
C1sq20Jz9GKGEuJv4m65ODzYlIByqZBbrJWUqh35tC0msRXoNEUFSdatb7N4zD3w
wqe0xe/c4cZutN0q7n0UV96SsWIEumkvbpvUWsmGhUWUk3DkK4raP9hkKmtFwFKc
Bnr78pxu7t6QBJBBl/OCG0WUA4++gfZqAgnHQ79T84Ut1I4tNZWiVsWUBArybroB
S1G8buDUzKFjTNvOX07VAIaJSG8OTqgqNORsZzBuVqBzVFUdiAxToLf1Zeg1+YR+
OVhl1OjDIzMYSufzwFcKbr8vFeLE/FfZk2jve0DCFuATtnq6eCCOWH9eyX6X4/p2
mYmI4veRj6nNRnLexIg1oOwLvHQ98Be2XAbFyVVqp54lsSh8sZrfIE12UBYUSeMq
m0cXRFP2OuRtROUSORT4OgnFc/uiv09/Afs3v2rErxUQfPc1bh53k5ijNWi/P8is
ltdbopLCaWSapq4Xk9VeS9g/+0dAMkceJ1G0+Z1j5mTUl7t9joLYGAvJU2g+vKMj
b31EVsPfh3BIEOE7ZFeXpppRDqwHKuKJD3oUnLPZlqLvmESOQ6kpChPcQ0hQ8XPD
FCdYWrjEnKpJem/iFB7qmpEC+fwWsIouaKTMlpRgIey7YCPh1NwO8cXNKAyRcaXF
6b9na7TaXKIr0ADNGXnXfw==
`protect END_PROTECTED
