`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XGzpwpbyaAqd7H+qiYqQNJUielt3bOKDHKiBshxTqWyUG69mzaDjvtL0m7+HjezA
/Uar1sSWpc5V+7GJqCf39iIu3vUBx2IBW9qWH+ewqRId2l99pD8+rL10USU9xa1H
7XAjLs64WwamlNM8aREd26fM7AGMnmrMzzc2Y0yDSpjhBTTSn0TGWcuXbQL3y5i1
T4SxR36dstpBGvBtdmIBJJ4BWofii34lu5fUzZj6jb2PZGOdbdMOI4WruPc4EnNs
0EXB5axbpETun2ZxNal49tX+84rqLog/+/lTy+rpXYHboUffBY6bLQAdeT2Y891C
KMZqHIjPWmx1Z73uw2/9Hg==
`protect END_PROTECTED
