`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lEKmMVx6bgw9ZKFeKo8wKjoZRyzv5DLdQRlE5efOw9dVjiA4Dfsm71zCIz3iN/B+
kw1n1uvi4KmP7rTD4BctdTMqXTJxW/E7FFIxTVMDay3VK/EmJhuX2vDvwVIxMLBp
Tra5UPRrbMe+IOO0HC3YGQfSMOlMXVN4FRwyKMmDD10W8BHmeWiVWsBISwpkDwR0
vnPR3GJBkiYz6Jtq7wndYyARYwqf7fI0rBwAFmOl5VHb2QBnoyOu5DVUzATMDdUE
69VMJCgfSN6ZymmD2SIakMZs1SADW+0i8PblV+aSlDXGs4Qhi/9xiCRWATAidXgX
jWXkn/9DFRWCrsh9hatjJbrXagRa7+VLfnInwYCx1NXkYwQCu9mJlhr6DB/wxCgV
exwee+7L2w1w/bgyNylpn1O9iwRfBnFmTq3DRFV8EyRXQTcLNop/LWYAsylYjxPV
/bZ71crwHB/DCQnsbJZV1dlpbRUv9/cTrqJbvS6kbXjZCr/9k4mCsgJq6JErNmny
CYystgjps2sY/VMlFtgtX/wxk/srTHmSsIabC8IvRevVP53B5d+ozJGrxsEkcBiT
J6Wa3n5h+ul7WpM0Lu/GmVaIQ+d23njvPaDmOBJP/cNzX767hi2gOAYe4/tvsokS
ZtMO/FijxSuIkeurtnRzgw==
`protect END_PROTECTED
