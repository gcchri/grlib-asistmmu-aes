`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5/5EfLDhWXcH4sOFBzxvzoVs/i0z1m+DiaoZgs0fiW2ILfmxmdMR6gsr5rFw0DZ6
YZLwwkDSABO2cK1L+Rv6740M7DQZuEpchISouh26rUe7T/uDQ4PlISJ/zVCBljpA
jRJvYBtyPJ0PM7O8J0MI7nkTyv19yWlg2+egZ2suDAx9mSNJCLIqpgstU3qGh+bB
Mi9/ljMt5kucUQUh3dlZRPhYrsUg/xfGeQdLnOvP28qtwiKV+VrKahdGGHXKSFAx
ZOGmaQkxPPNttwRdisXfNZ/jWr0Ql5H94vfJ+OluJN78Og8YuIujgrlDwHc1sKuX
XtCl6P0kziKjAj5nbZHTDBKg4IsAeo50mS3QPwDy1NQTwy3kjUNKUMpJRxcl/fTe
k+ColV8qpx2xAHu/+1PG+d5wa0jjKudc/xHPsul35RYfwbBgugRo4p2vvRzvQJRS
H/6CvaqD/JYRh4kCuv6Qex4JnqfXqOnEwk3qe6c6PM08TUC9rwzD+LVH7RdqAKCt
Pjdatusc72a+1XFpfuOBgg1YuuB/BL2wrhP7PE62XWHPcSbUxAnJxHkg1Gw/r+L0
TUBcrFuKSVc1UUyvLeFcv3GTZZ/ERluUPG7+2lTUj2N+qrmKduXGaWmTqhgSqYbo
hIHO6Hqcy3uLgWAQV0rM3hm8DVae1mfBTlLYxRM8DWrTK/gVgdYpJuE+eGd9PBqm
i1qP+ru4DcSx7dujnV7RIdmAkAmpyiV+1PnhbF02VoVu5faUig1IZMSW2CKX8F5D
C8d/zOKX5L4jHNACiJHGiPnvHhEsYZ5z6wC3NC+LI1NxTaO03gubcmK6CYomuD9f
53EfaNGp1Y4Yuin9vaQSIg==
`protect END_PROTECTED
