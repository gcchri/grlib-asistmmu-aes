`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oZwPYIpv4kihQ3LINZvXy6f5A56XOrVQmnP58R8aAX8KOYKjweAyaWum0M9OcZx8
ZKY41enP/aV7iu4xGfrDFDUtq2GDNnEJ6c9sShYssQORDd7xmjePqNghiOfiMNgO
jzfcXfld1QGcV+Qe7m55HRae/GaiaW+ed2rF1BkvSfiA1pWYEG3o5CoPcAquFOBx
JuHXL0MnciuPKpu6ZquoTj+71VEpnG10/NPnAGmkltMLIoVH99SuOTFNthgSuAuX
1ipfgPAFe95kkVXR8uryLg==
`protect END_PROTECTED
