`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nKTIdfWuZVlTr4/qM8DklSVN+DbsUlzSREdx1DWxAOUSUAkDKDJLnjbf0NdkMleZ
VlirkhKMvbAeTQ20NzkrA0vIHM4N9whVuQRSFjiV1uLNF/jdGQEU1QOLWBCG0SHu
uyStNv7klUIz7mYyKDvxsOXayGsikl6LOIHiwYIW6UbIsWyJ6NnrdQRtT9npn9z0
xwkEDd1AI0Ek9JLmUnfkcbW6GS32RIQL+h/ZH57QTsFxGamz4HvY0xEZfUaqCi7R
6RwSldNpv76DWOZpB7C8RDJk8LqHyZcrS8YDOv0unf4KmB0MYVHoPVlR8C9Z5q8Q
AWgsY9ivLKSmQ25LE8sX0j28Bn+f/+EPoRFNXqNBBvwHWMey/2jNrNO+9zf6DsFa
xCwSMBs/RvWuotHzd/LPdatdaWMP91biZCq/RPDtCmriKGV1uegWwj/c1LXce84h
G8aG7y/RGx3Ulx0zdNgk47hDntPMuV5TlPC/FnTE92ZttJAiPYq4r4HVjaxgNGhi
8EzNlOGcxCIN0VLdJvfQoZxXcYd0cggVbfcLtOieNicsROLyxuWMp+o+WH+vQD/e
ZyK3XRp/PeKdaWWZI+YgQZkwYuYIyRw+qcbxWtwzDTjd/RfZsLN5gZ39uvSPSyal
6aXvSLi72bB0wfbtAGfnMwCq1mc+j7erMqeBEKpyV643c3cJBxj5KPKdzxjohaTP
0R5qsc10f47sXYT2shst2xvHZlp+DH9aXmr3504dslRqloQKCRvTTeTBvtoWxzaC
pFIyDvxCZtjjlv5nMcUGpaSEFoKzZD8B8hJOz/LIL4td3Mg0kMV/+4xj0SpQbDti
Rs93DYpz9PkeqvVO8oIIBa65X8TF458xFTPeft4E4ZdtPsBXa3Tmg3EdMeIFqY1U
JgQwjGeD6iUIlsSp16FHJVGcn99ef2x00lsVE4O2K6tZUgqz1VgxtY6/LD8wM+07
DjL/3BdhZXykAOIcFFe/4JBDa+vkZXxWK6uIvDm78nCxpqW4j7wb5Edroc2BeogX
Wd3rX1CoMoCzmzMD+Mpks5j/3apIZNMLqtgCIeUCHmOSg93EAJ8k2nXrNBaAj/L6
BK08C1ZUJYOGHYk4rzLra07/dEHwBqU+1MOLz0IdemHeAztyQAxUFj3lysBqES/O
OENKrVQFdqexZEDbgyF+CLhm/AoU2xK85QAs+TRD//MEJXUW/RtJWdVEnIhZ/XU/
c7mw0JSEygB7+pjwU18X9Vo+PiuCJsSoqRazPC5DyC7NJxETCF5doIJ2HigXIABC
A1S4potWkYxFIxphb6Jf8Pt1sFpUQSmBL1uWgQdcoOGaE/+fbMa87y9HUiujx3Y6
KiCF9JCnJHDjCCEP8q/qq0vh+Jdt06cYm8TtN/+Ct2/dwj9X6PxdRybZl8TGxlaq
jgOacSRp5jseBIRukJlCgcyNZL+NIutASjy/KXEfdGGZj34d4oQVhBq5ZOb72zsg
67hEewCgHxFg2nAdC00noVMHmXxoZxZqLOPxTPDLw+/QCmnfR9vrEb8/dHlnNtLs
f8rYkiBEKZL3Y+kfdOAnU2pE5DY5IcyvMtk+oXg5+6G267KJpsMitrk9YBSwdtoy
avCXCOe28wqVqtL/RFgGSuQ/9bsuLEtTBzqux5jgbGddbeZbigzX1KqSjcaES0CR
e5Ck5RHckKC8P4+QdH8kPfkDZzKImhK7Nnu0q2phoobTbj4Xb7LC34lQmlhcvt7c
ZZatt0IWYct3Eb9J4fdHzMYjMWDrCgu5DE5axbV6FDfK9HAOnoOq4nwWHFZnmsNU
+3fbxqg6EiWLQd0qqthLcGWTJ8pBTirpHprveQAB7f5t/in9tIgbaw+L8FeG+kJx
g6YzQaSzpNr6Wcmq1b4O5LDqQKEdrrz9bQsk/+CiCq9qFf1iBUCXn7w0I/04M8Lc
8IFq9o+CNH/C0FnQCYrQhn8lkSJiNUYYMGvG1zOJrp3jmOYTqiGQX1vJaNZBaPUL
SO4hcPyv+7pISEvCeSoSKd3bxrYa/57/Xp2QroqFc99ObqRq7RX6Q2RFt4KnsQqU
4O4atHrq1U2aBwIM6BYl+In1UlDTVIEelNIGDDd7Dc1/6nc2R6qOiRi5DUrAhn4a
efarppeP4ItyoKXLDBRYDhjxHWT35Etuyp6aXjgAQt+8OwfumQbB+SLvogQnS9RK
BlVOMuSQuOySqlNDhRRxp46mpnKFdeLJyk8SilEqhIsC/9oYCLDtlRclG/ORP5go
q86idD35GydRVdU4vXoh7XdyicqM0oOa5oh4Dit1RTzazzXa8BsqU8EwBWI6Ah00
sR8djNTcWa82u0Za1clpChEOV5Bbb9AeqVvW7or1cG+hVuKBL479Jjc4k/OiGYig
f7hAFjJLjpcQUtBzVMvo8Q==
`protect END_PROTECTED
