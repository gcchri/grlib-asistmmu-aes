`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NzDxjnIhVFYQ65glnbksF09jUfHOdEPsCktR9Hip0zq8k/YzutbSrhpjjbyyTy3D
88WmDpqO7+x3KaicNBFH9ETkD6vCZteqeJR8KJyE3QlYE85ME46ViXQ8mEUWwXYu
4hmmeF2zv0WDZBsdju9HoF9D49RAtcYWd23WNCLcLjC7OgDM+hyP+2AATw81l3G5
Ib/eUhMzQx5OX4nevCmTggwg+cKYVi7lbBan4nR09TrC2oPkVGzPff4gD/k1SJwi
9HBA2+61xUISlZgmcmFDkBRJrzsxUir2/sbkWXJ94b8cAm376Athx3XpHKimR+Wu
pL3OMdQ0h5WnexDSNWfXogcAA08nya40yys+P8d5wc8=
`protect END_PROTECTED
