`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
op/YprIirDpb4aK9beVcAZ8m5copy8xiHx13MkYhi4v9PmFEc7u8m2o07jdam6Zf
5odo72ZqXBWPWMyGS1YV3pPTCTZcER5dW1QMjArwqDT20zI01ZYVFu6CC6krbtlP
vEQXnQyuQ5szF3Ky+k5syVKy3rWgO9bIPkGy2L0aVO9So24pHZHAe10yWhI0wB1S
Ic7Lkzi1MhUgEHMrZ5GiyeuIoaOHjwF7TtikWos5wkV3iKRbrScWwuyashT4WuJI
UDik41A9VbmoXh/mG7lNF/kxwDdurLM3HmURU+28To59cSQ5X2rtD+1Bawbkc6Nd
RawV0KHseBHQGl9xDc42kp5/yS0fyEm3n0dtucmrNTThIygQplcAnXQ/psryZqO4
`protect END_PROTECTED
