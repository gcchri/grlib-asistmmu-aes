`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nI1Jp4g2WQzlssmWpZmbtTRsbcPEIZVZh2FfTkJnJkyXnSZ9RpwVlPye3mKZynlg
CBFnxplciqJjxYXco8MG1VTxbYfUKri/YG5g9UB3PzCVUYX0Y7bhoVmO/hdgZ/Me
epK98AatWdMU8JEBC+IfkgRaok8aFn6DWYWr6TQOcPsYb+ofneu/7U5diUgKY7ri
79icvNcWZdMX2v64lXu6WGem311MMvP/dskUdy6Bu9R218YVqlJ/4rG12DtiNJpT
Fb1uHsH67YFmd7X8kJ7J4/6upc07elVUwEY20kvO0tjQqzgHAM0Bec/7ZxsIXTT1
FrTg0qfCZrS7J7PK/1DeSfMlRp6nJROxav72Awq+gggp29YV9tkz9Kj4NukhqHno
oZqUz98sb8tRjWlqC413v1iFRwGlzJRR3Nps/OnmVCm+jpTMU98/25D0U1A811/n
qLvjRGytRepXq7toB9qp1S+xo8MPyenauw32OvIf64Q=
`protect END_PROTECTED
