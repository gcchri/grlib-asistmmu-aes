`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u+9nxBzganr5xurb3CZusFQtjtg/1wIQ0wC5FgdUTh5bATWRh6Uunm35h/i8JSda
dNWIOLjNAoxBLxVIESWeVzw7LEbkrq7KsmfdrmxAfoQA9t9D7WLtzookgtXnCwnb
IoZlEkZ+z2wFwmi5doE+1T4cahT7yE4MR4mh6SN+MSsVVZweSwYbbfz6yKPgVjB7
7hXQwmOx+PktsROp2bsXmzHfBVHGjLCiOzEVa8+79CucAX7JMNYOu8Bn/YkIWEoO
gdS5TfOTm3L5PqWbf8g8JKjqk2fR0sMGM/qk6G7vH122+US5SFYnJJXwRzJvbJck
1PuwJFtt39ax4Mukgr+Xotuy2LJKrtYy5UA5F/qFWIZe+byNDO46Z8K5aAU/H4hc
qgXIKiku9Dp+NSOZIOJwbHmHkfj9oLToWqLl2ixkZ+bZZYBpbBnNznyKFNz5TrBt
PkQBiqqyLRGVHZNtVMLHTwCiyCBCf7RJnQt4C44iiFRlG1aHyDRIZBwOkXycZdc8
07jdfAJwWtVm6i1+gQ/8t67PNvBTpS/qAuds6xSWcN8zsWcw7hf81t0JXXAaXFJF
F27N7OM3+NlLmbPo2RNU4q2S8CJxmACG/8XLuNS7UotULnmo32t/6RELD8nqUmny
U/3soSMKT+HnhoI21rncgA==
`protect END_PROTECTED
