`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c+l/yS1yEk54iOeCueTzwjoD6t24ksbUM5SdQw51XFxjgEWF25+XO1P7C27dMkHX
tnJzqqqKGWj2dQwGfg/00QzLK8HrHzrxSUokOsUooAJfZHgEner+ZjVlG/R48xg+
kFTgIevIqZh8643bzFJ658ZFEIydBC11oCKb7xikXYGDBhYypXHDlimRD40S557d
wJFJ6v/37MoEwetqUtlV662cogIpOyzgAUyRaL+iApGpFicq3YSMZz4o03TigdHv
IqUR30jvpfE+QCq1xGF7DAt5/aa9i1tmmLjk3ikjZfbArXFtm/aI885R8cASlbxx
TnTznpHhdtgd9qUAzHsiukD6a+9q0PPBaIR/zrVkCw1SPCyZ3ep6khx7Csh2v0qc
T8YsuJjLmo1vaPFw9j5fHEGlunclxvziRUwwfJ6SsKSlK2TLay1s8ezn+4dfkXwp
PsjIcTd1BOi0AmnNrdQrjvMRjlLJaQgPObJ1ww5JA0chJrwijSz9EW+jswBffxUn
hJz+MJqgfIGu9E/aNmjodvkPnjrqmANABwjWNnxmTGuBS4eh8iBw6UGF5c+PJPOm
QBZameuK9CD5JE1n+3RQdCjjxvcFjuUWUEr/NV2g8woe/FbrR3cIN2GJCtsaRb+P
nrcE0/bTrdCF2zA19xEjrTtHyuP/waPTX97tkEC5ssA9o/CZt57n2FJmTmbFvMd5
dsyb/X79Ep8MKEmbNU7qVeVoKGj3j+bDMATm4Xgucns91E4CsJvx8TEdbG7AfZiv
rnnlotxDx4PiiC+IdezzJmN3Geo1lO8iT+5XlOlxtN1vxXAm6f0nSjl8urJEDJTu
hVqG0pd7Ekbzw7/DBp8AspaihhKIoMWdcWUEcIdNPDCA+1tIyAyvW+YVR1SYsx43
FjwC2nzDEwD8ol6S/sfm4UKmbxcXnO20WdFVHN7Hm4ZboAxJm6w5lSgZsf3kC52P
PApa10x2BSISbtqYkjeorN2xzknViG+sbLJpR6WBslybdO9Llm+IL88TQcZ7sxbG
Vs3CIhLftuHrWMCD8FVjEMrPZnM3H2NmR/4RGwFUZnpGUd7QptRXEEaqwrW1IdXu
vFnK2GooTGvUALe8Le7ayBVoGcSEPhxzlOlnTQMCDy6aWRNCSuFXx4+uVr6XJQGp
bMSQEwsaAnudYxYJI4KdvR6+4Dp/5kmlylQjaR5mL+QLpgfhL4s8QRT2vXUugk5F
1kQwyLCqH/joiRt+StLepmXNxP121PHy5wLdaiqDZA9TTv63skf+jGl1byGKKpYM
4hsf1s6dYJ0HFD+jLhlMSsR5ZASmCyWKGoEoh2dOezM0A7sIRqPSOcr0B/siDXhP
arjfUmvgaRtLB/T8SU0bgna6jJvg1eYfo6UlOl6F1mjZaTC0rMzioYMvCTv/m2d6
Ht7HNOTwqMq2D+36J5MMbLYH+LQLG2+LNRVNSlUiFESLpz9SYIPi4OMP3PbYAsm2
AslxUxiuyFzZ1Tf/9OG01OlWeLpC6AdludRBfkVwbob3Glq9kyL/flJYnpD5TmsF
cxaL0OGfSaz91wLH+FbSrxte7LETFrt0u2dwqRncwUuuj7FIU4RWdbQYZYcaC/0M
Z5b/5Mf6RajTM2jrcSnMwkXv6oLeXh/jYJNhGwXQTHEBuYqUQdTG4oNiDimaOvZu
dpVYhd3GuwDCGAeOYlcpTRYGlp2B8P6SI8NBKWdotWBj/LktADt5oslaSzBzH4Mx
9a74AfNSAjp59my4o+1WkCYrVrAqFulOrA3Bx+LSD7NaydQUMPDqeSdu7a7/GfAd
bfcwENklnS3es79Cm3tqxMSqy2P0w1gkged/3CRy9q/HJjX6UwTJvfmatz8UQycK
S78E2PP3OOHx40UfeJIeD+k8km2kvTHB8evTo7UNT9bicGtu8h0Pf49vApwOYeTd
f1J74riHQH5PcHt4oLyjfvG1CdHvE7uB4EEdyvnnp0f8rc7emeYtDWDR/lNcowfV
kKNs+d1+9aR+3ZeUIXm9ZlWQbyr3VKrEU+O0rtz/j6ldFq19a9I7zAcL5c8xX2s/
6vQx4KsSbeaXm6VXI1ppmsNdB0rSLu6KUo7WjZQjdGpKVEP6tFrOWQTuJHsNzMsR
AiVWTv4HD7XfsiSVyRcLbqEY4GS4uXCkMHNS1ja5mR9z77zjPbcH94rFqgVtuDvq
It9+lKdynvaD1GeaRHpnIqSyRE5+9Y+cNSEEfiiGbwEB4zkr92caEA9VDhM1XT6x
eTt/X1UhPy3n/soskN1nPw4RTEPvJ+/yyPCrFLPvnIWBL3kHl6S/q+mCgFkb8mlt
UF9u7SoeID/cQl7X2rq7rgMz5o8s/P6sL1qxvehjaKoPMMNXYQRZYtbV7+gBp82T
s0Hrx3WxyFGrb/mKk3OCkwhgJquajl/+l2ASWbopyGRygEqg4qNSizbZlqdfPtVr
ioEZm+IJjcqO5DFnquzcuAz7I0JJtlk12CXRORt4aRqq4cS6ZaSGO61pcmUVtWjO
zeW+766j8fN59bMB5Hb916VWqr1CZFB+k+PFvo39ogB17A8IqvG3MZAbYxvSyd4o
8ltgLCA9WBHT2IVUHfoZHd4iyz2VKL936+lqo99GyXfI3aR96rlXx4H8bKTTIg9d
WW4+Br7hGplcdewEUq4nuoq92Q0lgMuZ0eVq1WHFp0BNGgffvFDucq8A7dk1bwVa
AusHgiF24JwDSp5g/PZozGAb+qShI/5oSsmtWCDO3/wRg917nHbTM59inZNqOvh3
3oHqrXOlkOb2r9+ic6/e9A5skwGws3RwQdLUUW2b7BAv9MTDQdhUHBbOuJWcNGlY
/p2dmIn7k9HhMxHqqvvwsUXLfzLbxL+8sfg/zMI/xyPWfPfaUnzzYO75x2RPpWXx
kPzH/d5k3LZ6AMrS+EPfwe+txMQVyHJ0xLhGJgHQaHzTNODAFk2xI0ooinHg40lJ
6pxFV+9rgvlmG0mKbl1JLmstqNCoSsYi6NACa/mUIFB1JIbs2u7Ue4XFEbO6H7Rm
qdXSIv7wQGVZzKtVjEMGkwMgX0c1zYPdUxB/wOsD0FukrbDA6ddf8QqhhvK/EkhP
b8zRPUBf0+49SHglO6KaOMlX19ILq6taOsGKRcnDSUAFbAQmZoVuy7Xw3lnTritM
mxrX/QAD8rt/wY6yiSz5QEJ33K/SHoy8nvpqtYLeewdFV6jHkvXccS9oJO4wwN/8
FC9cYkOoiw2Ihx4mbXEk5g6+Y6vWbWPaxnpfrrqaub7ZjoHq95H/uDyPcm4GOII/
TeWeHZpM03wAQz3lG8MRqbKxt9VRRGdz6+VNpfgHd1tlsKSJYCuX7U/RkvaNLNdI
bCWOXf/PBo54+wOvDgAt0XEtgm5EJyB2hfC4eAcOqdMIgMDzCQ542b2kLmeikj66
g0CC9JueQmZLpQUnnkt817FiUCoO2CFq3+pBpjSkbUSn66iFS4lHBrBx4P0hAZ2b
55HCD7lKInKeIcqxJuoRRNusx/TkWUG1a2vW2BVWjAy1/0WQJsLfNOxd4c+wF5p6
2byw2LO1eT8SfwgUC80uv/jfuV2zkUepPPVm6x7cAaMvh+yXclNGyCJBwiIMXuVD
QBN+Y2ujqAyKGLmQAGMohPyhVkwWZIYAEcq2NudHYbLJWgFhEmQsBnAsFtD1ewjw
r0N+rGCWeDPyfhqbELlVpbO9Jj5MCCZA4V70INpCUsw/DvAniZF9FhKuyC5I0Egl
pNdAzj49nZckh7l93TIWbBBldgSttpUUU3eHVWZzq1n42LNL6RmQx6BCBahPUzZn
XXOW2I/VxqEjBFAS7WSParwg8O8euMkz1E9b2YGUYkjIMvyyz7FwULHZPxTjMbTs
wXw/wpfqNbJofkdLYAgdrH/1XaYXM/+tDOKd1ZmAIabk4i4u5PwQNTuTGM0mNYs+
9yVxYa5eaZkzwJ2HJWrfu82b4m2AI74ITU7dyMiOSyRmhxFsCsyuF4vGsnfvbWBn
8uMdfknXLJWKfqTaL0BLPXwALrOjFiPOn7aZWLG4EIw0lDk7VwW+fJwQbDP99jQ8
GkSIwUKYul1mN2lkiQYHLSpRJk7VoiAJp+iM0V3EmjgbSDP7CtxHfY0IbLsQX2p+
2DayjStgoKcgzI6e7lC3wF1aw9ZVZTbNEnixYVl1v96k+RR+LFknEkKhX0Aa7T+y
gKxd7skYItreI4MchxglWpU0sPqi5ZjDfN23psJz4h73LG9C4LIbEpQK2l+M/dhy
XBco3HSBsktAVA8huL6kLKtOQFNlGAAyPd1adYP6c0k0v6UF4bcKtPh8HL2hMJnw
Lior/s/KdBW0ipns0fD13r0i0voh3C+Ahk+4YjhbmjVPpVMOLkF6+vTLftANfqd3
2RKFUfrkgEq9fcszfdkGPrV4xEXgtunEC5VoOgLIDHokhR4FbYGqXSRWzm3ffr1P
g4Y9wT4x9jjyYxB8XsBxIrq4WSvtYnH5ngEdWOdcUxjLQeFgpdB5dWSBlQpU8SfI
+SeLMTjXNwyZ9c5dQArXmRIEos+nghDnlGOvpBn9Z9Mxy/C3crrJD+V/6/x+m7AG
omrfJn1KZr/aM94YU+L3DwqGcRBLwQr5pGecNYHa8hEbvcYZFEuN5USZM3wJcj4s
qK3uB3ED8oxA+OZMvqtQqQj+kYGuMn24v5gGPv01zrXA7LC6Z8wZcmK48yc/qA64
l7wtS1PPjcp80VxLPCicIHZ0WBdt98VcbGFnwPnT5afyNiUODMfKR87//8tXMxBP
FwLfMPD6FrQ4wr1mBgH7edj91r4yoSUKenWqGELhPmIyPKrQvTXwknYtjF0wmADi
/SBhZwQQ/HPPmpDcAWOed0Ruui6PPK50JSmPiQ9eitqrHAOdH/7vcHazpKfzQFWb
Z3tCkjlX/07XOeVtij2gr5w1ZLGR1WZl5lRD/BOjsgF1iJprbI4EtdbI3bO68ait
tnq5z5kXa0/z8MyLNA/Yv97c97RLUmziAv3nvaJn6kLHQDGQGX5r2lzttzBtkbdP
iOJIcCy1HFaNmXnVlv2KCKkUCxfH02fosE+cfDxL6pTLI6/L2z1A7vFN3zz4pETz
T3Ixcz4xiCTlFjd4BnQ4WQ6InXjH0cLYRV82pTvjCYXAu77MTMY+sIdJpwzYCUCh
99HyjQImLTQIEZY53+JbrCrO7royjix0FC6ywUZ300jVUoVKyn0h8N1c6Vd6Tsux
BTuqBLaDYKd2Sg0TPbYp7o/FDM1KqrknWKjznDgsLyhu6Pwy1YIoCtAfpWyTvjST
uBRyHv7GeSp9E0Q8saAK+Kv0hnNX4BH6ejz5o84eVCH3iZewBaioicDzYGCWN6aL
ko0O3C7mN75MJujVVKD47/+0rlTTyedO327QTCnQ9x+nh8HT0yLfNkjLIv4mkfzE
Eb5ic2EMx3Cwyogty5zu773tazmgjp4NNuKEyNWvPJfxnBp5Syoqsb2buk/AjMzW
As7UtIS7YQgMUhNm6ngfJ7MHLMWJW0eqXgfO51w6G81Dpil34dGQbNQyvZ7FA9Hn
fgIxn7yUrW2OmFX9VXON92YlxS6/Dtmnk0hAjZYt29k0ul19r8UUsFDVfaFyvAWA
NLZsIOjQrjbWD1ksKsPZdw==
`protect END_PROTECTED
