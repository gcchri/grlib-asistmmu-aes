`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hyl0DjJy/Dde1B09YigdNq82mC0fprVAvrAvxYF4IUfiecHX2NmsMtI+RPjN2V/6
vSui1g0BKcG63G9LUcnSPRbtzICHSHMjHrHOCwTnE2XY2O6SJO8gEGYoKBoi7/U3
PpwHSJOMxTc24qlKZNeY/uSQBN/BqutjnhtPDVKiady2C+gQwjMtBOkTyXcInuzf
G+SkwnWtxlsO7R8P6usugbv0DH0GsmZOXk4ahJRuXTcUVuXB4p/r10/T6fNWnz9j
yWcSifVRT2IQj9GsAdA1Ew/i24f6uA+uwtGklDxatADSvipZFnlY8l6pjcVVLJY6
0cPxC1SAkziR7syjPZL3P91eE3V0vAnN6WEGQGHvrSGPQRJBa8bBfHMr0ZJVihMB
WzZE1KbR2gr027Q75YjWP/hJcHDWbAbA2SPzxV4AJlStR48yVdOTujJZ4bPU7m3W
oZ2x/eSLqxokvmaW/9Y37DUGs7qFjqMboRtLkNzW/aA4TrU7vH8q2PYlP3+LNNAd
E7PmGUF6TMUxaRWbnMQmNCyKANFHY/O1PGgGZ7Y1mdc=
`protect END_PROTECTED
