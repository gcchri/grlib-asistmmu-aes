`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
noscB9TSyywsmuHu2rtm67JFu4ybb3Xg2HiNR2RJ/piNtUTkCVpALEUZk6YqWfPq
jbg1epMkBMpS7blE0WAm8YoaSXuNG1EdmE6j6Pm9UnK4DLoNsZU5mdwV/6D8HjfK
X7zspmT/9NmKrcmsJjg0MqF6y3VrADtj0oWIbCPhm95X6WQipRpa9hBc3jGVdM5i
OSD7fuaKQVJZO0o9e7wsOIN7dt3NJsgynnwspCWHxfblePDfqgPhg9IwwZ6kwUr8
otcDTRMq30UNUmXmYvRyb3eyKXz9unaXqYIH4fovT5uxqUUa0vLNKgWHtMo71Jl6
5fNlpcPGpUl6xCcDP9wKQhGSR/M8kTOeDA7K8IiB9vS5cMdOgZx173lalmAYIFX6
+EV17PXOtXw7MZrJrPuVKjQOYYVAobHQHQJEA7OfvEQZiSWzWBTAxKc+WgHo88s6
eH1045z+/FTqU+PU/kYhswPJO/FwCeJ3GxIYKvcyo1K0695JLEzZbJ91G9XfEy8Z
dM46OY75fLwXUtqYiYsD0qwdgmTkY7WZSPuesa8n9rdoI78x3GMk3JFTpCpXN5VX
fm6ylhebpqSOnHoqpxzp9PTTP3ircNYU+yHgs4Q4HL7aP8JW2bXEIY4EWxz6xIOp
vHEF6Px5nFctpvuXW2GZK4hAZ6yhi0Zjp6jSqikyxnNwthw7iqCdfUs6FZy8ms3x
6IxukJti2wrOIM1UDh5aJ6wr6Q8iYyfLR+A+8RM56gVV5FzbteQ5HdzgNzMTSmQW
QtGfjCFyqDhGmDuTbwU/tR3YscbYoG7aDQTQVzYtviYPVu2hnuG7ahaW96qy1jfO
o+BfRF3lRNycL09sxeNsIBX4EAjhLG+3LPZ1IVSeO1BtmX6qW71R95AS0ODOvJjl
N7x5gkJ3WQ6QRVsSqQPbxOQ+FBp+jMpKIeje7ea4HX8xnGWeJ7l6Ybe20lmYpBGr
a6g5jqbt4yOCM6kFr+F4oZGe4BxUAU/a6d4CzvMns5JwHAC4eAnTQYsHHQkuvrmn
YAXTofMFHct/+mmUrfXFXm64FbD54hMo0XynumnkHOMsBUG4p0M4/0PmT27A2PWf
YBed0HHQjK9JkewpO6wZbpvwsle8R0htgZeswxqP/xjappyF5nlFaQxutjx1037H
BqzCaRA+ZilnFne7Fhgz5UDhG6sGqJordw6VBSKOr7+vURMUaAZOi0xvo+qzJEdL
fvz6D73R6kxIcC1dWH+24FJwBGL0VSb+yyeptSU4G5eThVZRcRZKoTQs89QArB1j
hgQGXCD9iO0HzeVmBeHOYveIftOl4Cy2fc9gHvX4gOyvfi0j+5IlaCYySKV3FXbt
3hbD35v10+MMBxwy3kZKHHeMLsMV+jWeF5LSX0r75B4pl7NHShXpoocFEpvSV81A
YptPS/DIv0WLNKxgf/zmaw==
`protect END_PROTECTED
