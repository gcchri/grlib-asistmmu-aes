`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BvsOxhhrEzmrpZwh7UMx1Wa2s9V9LvAxr6VehteRf5/ap2uYfAT5QkAe4GzUib7V
fX7Y4qeCjzJQddSs4Q4HhfuGghfqtf7c9yXZhcVGdgTwLzh2C7ph14M0Yq/mHA1R
kRTwX+kboaz2v3llBA2tap36jOhMCmBt6taZO6/1tVfU2t6LvFJKzJvuiDt+BM0r
roIYqd+J0JVL80B8rDAfbuFpTsjvoc2h7kgdXqMvrZrYgZKAsnsgWRJdb8p+uID9
g9/aGWfEESChDjb7KvR42bHLEnkv9hCaNZOb+72Q89uAijgkUFWphd9nw+Ysso1m
Dw70O9pinBSW6ZUa9TkpzN2+BfAt0FgIaT5fezKwIFkV/HU8UnK15XLOMxDXPwB6
8VPjRFOXYjA0+qCPauSeEKBTRERz8DNHAYpg86X49Hq/tShgLfHVFfKUkSYVMztL
6Hqdr4qzVs4w7OIRqmf78Hv+6B1GUxO9b6OI/l54QVIYDcdcFVP8BlIdVG4Mtwlf
`protect END_PROTECTED
