`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XDjyYZxxWhhTH1GSShywOg0tRMUHGSwl2WaKKAjolsOa/Sfxhcicwc+R5HXQLD5y
owyJ3oiJA7nFn1Qt1ZTf7mTLp0/K4508SzcGuWnGNjzsOBeQFyZqmj9hpP1m3aJ5
W5f2t8LoHYYq7F/TiKfWoG4Kgfg0VSW2ZqOAjCyCSwfJczN4UOt0ogWmpW1SIcoC
7stlohx3WfTW4SlD3JCEbik36Jk+KF4Wjiq+d5/PpQAFoEaPZ9DpBVR3R/g5Z++w
SL6a/RBv1Hl7zE5Hkke288QOCxPjC1HnHN41Va7PXU1ZLDbqrklFp8Bpp9hAm84M
JSyZCFalmUX3rWolps/28NQyFL0KRPoNQwBArTOVN9S3n793wL789H8xSWmQEEkY
6t5seNX3c9dLqFyW27uxqdDlZt5CCDXTSi704Oo+Lz4H9v3O6OacuTYnWK/qdL47
kwoWgP7dz36Ocs+Tnw6dUgpBFnx9YhLFJrgeBh/SeMFvTy1hiA5fxghHiWeTcpGO
ezwtoHaLQEd6131NdivmkmDR2lBFDKYHXjty7iHEwu+Ck5QUQ6EHzTEx8Gj9DrSk
o6aTNx5AN7alQErfiKVfPHFfPYyojfIrL+dSsZrBWwg=
`protect END_PROTECTED
