`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tk5URCsAO/EPfKL1xKdjFyXcBEI6yXZ/ph1r7hgJmDAKfMA2SeGU2FRQLJgbz4vD
4456aNLzjt3Bfyb5nvv3gv5VRnA7mikL1MpzvvcqqWJzBSwpunbODcJ+zVoftZzE
tOGn0entpAL6SWM0NjHhnt8LisTuL1txAUHhtg0FG0XsL43oPnycZfTrmkQxbA1R
y2mc+R1jNiuVEnHX1SmOGnvJ0piSL8ax6IvSqS9Rr5ShdMItZyzXp2HGPiB9TvcG
xGiVaEAzm6aOdtoCcwpQX4/XmrtfWUcIsvgkMbLWplD7ID/gIO2VTpKDZc2jIIyF
v6k31FP5m0fwwuZY7ztT6RXHPgYE10LOqdKzxofk7rV9YfVE/LeZv/vgK0INYXn7
IMzlc23z+Wvgxju7ydYqkmo2H1spoIzo6k7Si7p3Zd9wEi/dYPC3ZGHDbt8dj+Sj
fNRWL0kaOTozuNEvOuRl6lm7zAZEehlLlrHVnRrM+US2zmLYinWrpgZ3UZAY2WfQ
4TxSLQHZQxpZh8X97PzMfhG2jh/HRkMRjk1nk0Gz6VVAAnsAe0AlXtTxsuuXjK5y
HhF8M6iaVoG6rks6BoiOobVQ48gWVsTwXgP5g06vex3/O0u0CoelNMcQk50p/vtV
XSLCtRmeTSzOn1guHyFqe+SmAUlMvqgbXCyDP3grolEgoDQJ3kYfWhDx1dT+oMKA
OpH4WbrigmyqebFs5wZT6d06AshHYz6C06HWs+FMcTTtw3Wg8EYPQLBPCmAVYJIp
2QpmRewXQv0WDccKwQfOaRCmQIBw8aIePCD7QGf7Ck5MiNc4Ky8/NGrTbkd/eMtk
D9wHu+9uYyJFor4c2ZAyK05F+t9shA4yelb/yfzPQT+W7rAVxoFHoMpk7XDlAY7e
bufLx9btPJpfYe300uCKD/rTyShvInscw1i4SY/xm10=
`protect END_PROTECTED
