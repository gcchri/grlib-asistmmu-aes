`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xXc2j/0u9Sz2v46zlaG4tuVdoLlbSb5rE7tB+RPx8fMXqst8DjprSFBrGgFwvqNR
Ji4k0T4BbenJaN75Ewc34mIJ3KBGn4E3pGLXmjggsZrkz8skVmZbF0XtzC+WT35r
DJW7QpSysSeMTwM3/nSh9MgSkuft3pPFXsUuqe3aWzH+DO70Iedq0vVmydew29Av
1ZQZ2Ceo4TxLOB0MxEEt223Xsvd287K8hDcuyTPqD1Jz/BfpoUraTlSv0/gkhNI4
+x/kR/JdvHyT6333QU79JfCc7uQTMg9i26J/AQ71hJg2XLofbQy3rlOTBSWiaF5p
Roc6z5LHzOE70kCVZ+qJNuMVCc5k64KfFdgmKlBYgt/mRFTbDzIsq5FfJW0kxrai
LwUtE7fp9UIuVvSki7Xem2qLPvvbCXBYypt3Oh4QiJ7RP2Sj5AcifcXsJnJHgQgK
IVV+rtwV4GNg9S7g+CP3ce3Gg6uD4CzqhvzeRpW0sMg=
`protect END_PROTECTED
