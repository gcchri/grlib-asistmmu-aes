`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fqURPGrIfX3+vqaEs/azW4/bQCk2d05eKlVXZhmNavcOZsk4Tjy9zr8JeRCETyWF
T4zkZADYEGZ9aLHWUy85eCwc4Or6iJRYeRfUhI7FlSCXhkIxWJ9U518sHI7A+cqi
bfjSTpXAXhZF3WhorWK8QNs2GJoKR4ZomBeIcO+xX9tEtOZpv+2hvU7sLtdlrwDg
eVl7dnYJRAxU1mxfSLjNGw/9K3Y+yfDI1d5zKt3k3SaRkXwr1zh9XTcORdxBtO6o
MucO9027/a0ESMjfAvMv4bcs7OdNtEEXwbdKsGOYFRrpLeZhvDPT7VACoY/FbEtV
AMVnGlkvrKs1Hbb/WTdPiYP5vVnjcXljy7tOEtLbi++zFc343gO2XsV7+4eBi1Lh
aOB+ja5OhSBF8ZUM3dVf6yJ9Wyc4JVCnTaHlPbiwcQnA+vS5mEdKMA6mehdkRqUh
`protect END_PROTECTED
