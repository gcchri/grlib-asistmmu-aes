`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Obiv/4T1gLLz1g/d8az1YWQVn1WAPkODcv4X/01GV/jIR/TtHZADY5x0jmFQxP6
Rf7Wd0iwMncplqBfw5VMoCbtHjWiO0RR+RSS/4KxTOSsKXKw8/4VpFLAzbS7pqZc
kMT7UBn3X/U6nPlf6DAONmcS5tR2uo73rwuagtCJcnNR7mVIG/tEoAHiLVtR1uAu
8vX8nuZRelbOPiH56gI1tbThwthz/ST800vTTWSN4l9YqKJYEE/dIV/Cjc6IsEKL
umtx2grWnp9Zj581v8urSXRtEt7Ap78ltw6sa58CEUk=
`protect END_PROTECTED
