`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xttvWFo79KNW1TnHTBF2XIaEJbVTD7rp21EN20HBkh5voyd8yeoLyBuxw4ut6BKu
u9n+llpvJJyAfR7liUxXJ1Qvig2axJLDbeLj/kNDSeqQrlj61UH7WTbN0C5Tx0fF
DPfI45gYktBCLF/szu1Rw3SuWwRDdj/wBNZYT3/+gUhlTEl/dHzytSaTfBT9unp8
U6CMLGcN3Z0vNVar2j9UYDZAM0iQYGshspo6mDL+v15J6WNPP/rZ2p1b6oLUW3Jm
rNDAfp6nnCe/Gqd3aam6x9q739kHFFhQhoPUb/DlaTkWTZcaF0LQmKeoh3LwegR2
yN5ln0RU4FD+zvNnHzjPnJ1HeKN8FF6DiintjlF0ZSxpzuNHm2DARqOCrrIy6Lw/
y6QSCaAZpic/aHOfACqp/H6h/b6xZjDB8RXnIPxpR80fFp7eRiT1LJOW9elXTiIo
dZfjk0jhU2QUI9EEJZxuTCBmTm+oyEF2pkTIcakkUEOJL4FNZMRT4ulY4uBWj49H
AZlSBZKy1C/SM2Yuia/IR78dauz8OvO9z3Mm0WW8hL6YdcE3w2DtAVRNPwZxLnR5
Atc0RLI4+CaZG36wPN9XMxtf850R7qRdE/HXv1UeHLrDrc6v92U2bFYonljxu/O6
CRYrZ2XfuV+IuxKahh7+MWfLb7SJyPiQpQNkdjrNN6xwkGzBx2I9U5TnYNvXVnri
Wi3UOtSn1jLjRZaGrWWExtgmh73OCicd75pbMuJ5+fMI6YKm0qweqIbWAhYiY8BX
MCqVlnfimtzeR/PM1nI+SgOnJC/RMa7Num/9ik7+v3yYq/fre1uzVPZqUcPZ9u29
AUurn2iwCKxxgMaeKoot9cTejUrhP6ekTSPoa6OftjA0N7dlZp84rvYxTv5tnnk8
hsIUuxWbPoCtIH1LngiwQzQA0VHXNWnm/5uy2YtFVJXBJwz/ZBd6H948DxEtfn6v
oY5Q26gts3+mhYLttCQSGQZfWSIA9RjCIVR8r6HtyepwscIrx4QH9zP6OdCQ9JKT
`protect END_PROTECTED
