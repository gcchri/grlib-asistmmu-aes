`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T+vTq8HQWHC+7zQXLv2wNERA6AKE/XMy3b4EO6Jr2r2vzlp+bBwBN9GKEGf+av11
ZvyWm1tfESlIqyDI2/t+n3ZqXv4ys1CDZZaga+0+i+4thy90ZMqz7oUkYWPzWMf9
9t5wyr3Fw5BQ7XCd/92XMvpqLYnLQQ1bT7XksPavqxMRrTb6R0z45liaO46xE3bF
10UlcVR/lccUDgMGifR2q18n/mhXKLsVzTcTWSYhcQ7RxgpwV97+u8u/hzDtgvGl
vp9invM9JeEpnbTI1pNJkbCBKbKUjdavtfdWwRkAGRpm7RPNY/pRoaHWt+w6RK7D
mNfj+adoEglmWe9GevETh+Dc+yDp3kMOE45luXfBcSmNXOfijwUHZp1zAmrXdybk
`protect END_PROTECTED
