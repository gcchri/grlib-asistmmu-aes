`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0rZeH04D23KtFCf7VtJ3kua2PA4nPzx2256DSQLH91WnkxN6f5Hb+pLzPtbKgW+q
K3WEcecZxJgY721ONsnMbbrTbxc9rUXclGQt+jW1KyiQjsfXAkeAt9GUB1WF7Fid
AN+zOBWeKCXwFeXXAlohBKRHGyvGd2jgq7U0G4vSAWaYMisFNntzTSIksCeqjMzf
tZ7HuoCMI9p6F2+J3PP1uSd89aTm+SdYSPuOpY5jSc4eeMGrXB3lgiwem0fa6Xg0
YSfmEo08uvziSM1L+FQh/u8jdzxo0rUFY+aw66IYK8gqICxm8ZqaLkgCD7wqi23U
i2kslYTukx4tSMvU0qUxXZibjQUx7rzR+5LTW30aBr8GvHVMFn+ox2zJukRXEVKI
cnYFN5IzMtkJW3WMu7t5du3RNfE8SoVls63YG6ALzwFuhBzVQoB3VXU/VTUNZXxC
OlZwfFbOSKiPmIXwYKyhoe+1zmPscZQdlSLpaV3c3k5E4CO24xdbXkODuLINP5GX
RMuRMzI/Yq7Rs5B8fIp3rrtZrvBeqtdj82b4B07Olc8=
`protect END_PROTECTED
