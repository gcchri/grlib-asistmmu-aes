`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4TVEz7A/aUssb+rxos5W2d3vSnWEC62r5cW0Q6Wf07ZUst0EjfGKvwynYiSGvgtc
lLcXXgOHhgGd3IS0CmuvjMmn7vnBuQQP2AJbfzqr+nh6GJciYYPf/Evn3v2rz1iW
HCxWN+ZX5EYY7nuwDSvKHFmXwE1raRo782VFt1U5CG2u8CVNjBpj9RVlivUEZney
M5XaS04toqNnck0k8Cz7QAZGlpoFVGJXpeCMY8i7QqxOyMSanz0P5n2X49U9WbkU
zAs2rEbG6JqyggmGM2JvxHY+Q000+x8p3mz9x7wMeJ+gggK81B1tCEciFLQcgL16
ZdeOD1VeVUbHFs0xyRD+Xc2UO6rK0TS2aDYf4AGK+I3mEhGbYiMs3qI8wDVnibAb
rxEaG2ZtAZwgJ+fyu+v+FA==
`protect END_PROTECTED
