`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HcJV7TSoSCzePzKB2WSALKTOqjQxMTualhJKSgXo0cKZciDSpqkUQ0ZPDSn9I956
AQEZo89CDkCk1O5rLyx69rhwf0Qfo+Of9JcSgWV72YERwPXpvqNLn7W5ZuLgGZ9y
JZ5J7T2bLTp+0hIbzebx6FJICaIGbgVgap4F0aboGcgnfBJ8TnPqSfk2Q98ZJWqQ
eP1btA3rmIs3FAv4TksAZcua2xkNnF8Du4qY0NUCfaCweGxPv8jYlxaKdsz/JM6M
r/K6tsc5SI3lRu/6lP/tpnOWq0dwDkT0q68FEKaVZAsJmRxIA4BZMe5lt5tXNF5C
toHcTGIhpsnkZozsS+rbfw50IDsmLK+ETCiA204vYg+4si1MRxJteSZ3SfTnKvqu
fI943tdvl7oYmB9iXVUjEu0ijNd0DmQwXPE2g19b1jAyq34+HHkuJVGJ79x5h4Vz
iUYk+69nRj6XYbSWxtwq19t2f+KVDchFp/JxAJBeAjl3zSRD14UWlTQARX9aYDiq
7frqDSjxbCAH83Z5WQbLJ30icTKRhH0kQajbT5nM3HzJ0hZa8nEZ0JPtZNS02hdc
5jBg9tY0S3V91FPpT+zKDMDIYDqJbYT0qnXhQTXw7tBiGmO8ELUZX6YlKm/moK63
X0Aqy96EhX9pf/BMwPhQBYuDgUnxzwZEMJxPMB5rtNbnT0rC6ODeNo7eng4HjESw
e1N5PPRPha5HsOybmQrQjhlfZXfYWwaUbklnJ1skTjORedLa7plksLMcAzoSBBlh
pgmK9Nlu+sE+Qy3jerlei57ku28hpRGwvjlYz0v6xri6TXk+j8LfrV2ER7Dqir3C
xM5uk0KRGV58q1UIchVTF0vXc19Go1KCkSNjh61IE2wyac9BRmNsBaJpYh57FlGD
VeHmdfPniT77RBBJ3Y/CpE6/aR/3UmWECl106tuwikNGkYv6+y1StaCquLFeJ5C5
IQj24L76dyyp8stVjGrEeg==
`protect END_PROTECTED
