`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iU4u7nd/0/AnqLq4XHIoSBINeaytSquCt2THKm8BZ86sDpajJa4NMaa3XhGaYRzf
acAusRGH+RHMxSOILvbb7qu76rxywAVS4AoyVEDbFbSmkv+0dxSUaXaBg7n0BJXa
rxJJmCycmBle0l1VS85vylo4FytEuy8hk2O2b4F0CvvQw+WQP+vVryq0hrJgg960
W8YgAIjMl54jkQHiHJdjRQrzg/WPSbyXtcCU1/uLR0vX2BqaMSb0TjIOIb7OJSQT
6zQkflrQkf9hSHem/3JXo0ZXCwz8uJ3/IynhgbtPH3sfGyT7FgNnrKCJW1wBhe2M
wezNgpUMx4VFpuTSkLzlyw==
`protect END_PROTECTED
