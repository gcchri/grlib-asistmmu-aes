`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/bw6zqrIiHVwfRU4WeXKWHKjmyakBPKvhDf8LxlSxXjzKO34uSboeyHC1bJFUf6z
dTiqA4aQrJ/SBjXjkpJikQAaQWsNgUwA+6B4EEmOmdqIm7XOByBuUMVs+v4M1ffx
gNKhWdnfPAxeLUy7Csu1kaGu4Wdczjrz4FyiWhV8FdA1skRqcrEng8aDq5TYDEFC
taeb6doQmHo0iz+xKsF4CcHcZWbYwdQ5bz5Hd8zvvLgVZXpWsfqnmD8U8KG7g4W/
ZKtRW+Mjkfu8tkX3yoGkv1CxFND5F+xnIjwsmSZYxiwumS/hZHhYCsi6GWlerFeD
wabrvmuDvoeRjrQsTmm8dMGFWw1YWSJZr3gwYyEtsSS7ghIKhF8zb99N0kNEG+AO
2fwnMCB/j+yP0F1C13JBih+FiAswgSFLkKEgLYJ2kwumuhY68Gj3bDdGT31IXQTX
`protect END_PROTECTED
