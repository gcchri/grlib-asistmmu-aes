`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v1JQhV1Jo8kWMzXKvOu3EZz+Bi141HdonHajymrsB3MOZKAccKiSV1jCN1fn/zXv
yCsI/89W1XWI4qNqWUFYLsUIA852PaVigiR5OU30xRVWnOr5ae5+2J1eg74+KQHa
V2mA0mWP3eLMowKE+bmC2Uqs5xUxzw6v45MJd+Dg735VKqYDG1ZDgvTkjHEPAqxz
fmtwso6ctXTdfb+ZX8qTJVoLg+Ng8zL3iGKoBSItWUQIIfLPoLCx4qeZv/GD+iLb
LJw6tlP/qp5djTy+pkCSONSVrlCgIB8ozFdKdNxoBXwlozNSXVxhQL22OX5fJ+Z+
/+OCj2qnyHNxwaGzV71Rks046SS4AfA4tdq2GoZw1aZdXxKYGJ46dug42Po8V5dO
vbgKdEgAPocuik0MQ/Wy1m6egbApnH7r2mTd3tK6q7IZHnAXzl/f8UneIP8JBr99
irqoQSj5x5vVYdguJbxPNz+9YNkPg6Wu9JV+FMvxNd2Zm1tP/kuU1MxI9yxBY0Sy
SIU//S4UgwnT4XvPsrQaHpHOMRLfuY70y1Ep/HvPQ4M=
`protect END_PROTECTED
