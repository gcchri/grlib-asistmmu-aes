`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6i4wIX0kIOqhoKDnLSPEjlMERsOgboGybVeks860ebEPFAQ1a2JOy0QwyS20N5Ym
gacdq1d+jDQm6vc+FS2Did+/gFnkS5Rg9sWmxIvU6C9v1OomriM0BlNPdYq6n2Cr
w2MxiOsoYOSAY++q6voPey4D+A+tJcHFJ6naQVArQDjuquvnuhGiSN/2b9BrRHhh
ThugTMZ/3QdEx/4EACWGsmU7T9WDxA00wyZEch6cEYk8SUI14o4UuOl0Zk8qbfcL
7vZ9kC5xho/GssXNbxC7baM1FbWh2/ZmnHWOA0kY9jgg88W6/QQxpZvYMgJ+7gyM
cdEaklEveYpMeKpSPbXV/fylhP1yomGuOL0XZHU/vnTziguUMmzXPS9MwhL1FdhP
iWnimHadquzWVkJzkDdfCUN3MJieffrCXgc7EG+ixoAivn4cyZ3JjH+fcyiD86F2
Hf0P7KfAPgZO6xwDMHgjokTJny/8NxJS7EY+y8e0BO9LFn01ujuEtG77pfanIkSR
OOeFTeriFYciOqSLXaWdkZAbAW2lFRfTNTlwY5ITqa6VNjpRULd6KHrNNkSVdcfl
6wX2SB2w5Wiel3lLTQbWqk1ksalTD4uyivJWcGt7CybtxtNTzh+ZWKCr4r7v1fJ5
AZpZ0uyCIxQbHSobRs1Sl3beM2nKqPbZq4qHVvFydH/JZVJFRbsBoAcFP+LgCds7
jgLc2yd9pmfAbc0QuxWnwW8F6HpCzly9P3awiHNnAV0ZKUwcXBSR7qM5e5t1ZmNM
W1eubP/bpZt34VVgTnISq3eySq9rEto3Bwds7pEqnA8HNRnNlrWSFcKawqWiz2At
AqOGYTuwgSmuPfnXRniHvGQS625r6DEFov3FA9d6S/ajswbqXNKiA/74mVnP7NpU
jgRoszq2SjMiVHKg8nvXY0+4fHCt3VKOfTmvhka/WJ+UQCM4gcfYe4Ms1tyCpGTP
11e3XEkbFYzrDI1vhap7Du4tPIZAf7N388oPBIAb6MfVRZwE8i1dNLfO3B9OXWYX
SKA6i//8kZi8nBifWIzzMg==
`protect END_PROTECTED
