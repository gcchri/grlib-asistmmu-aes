`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S4bJt+XOi0D1ZVXRWTQjncyhlWEMNYjgo5HA0S0lCzW/oIAAR4+pFV3J28hcnLBl
twJaolUh+INYlAxb+XoCMDKuJ9iJGgxvFHftnTqDWoK2dJSdVOSsdlGKQIz2hcRN
qVFySsLtd33I7Yp/7P9BWXRoK4X2s69MWgqoUjNEvCfvOAXJjwyfftP9o3zTBzyV
a661WJUmAmIJnx9e+6y0vss4t+kGjooVkHxe/gEqrfII3+wq39AdDEeE02Yl4Kei
w2McZIbODhVv1yIy/B16eCDQaNRR3A1iaFJzEXIegn53UtTZm84e9InQKz3JedUs
HJpkjUqVq2mKTqSYAeLc8d6miEkRDogntPCceiPm5VOBnKy/0kSxWNl2elCEZo9/
zH9cDgSowQAsxDkHhMXPjrWqzZmdKkjiADoukZphnaCLp9Im28FmbepASPAcbEY8
56fTxQR3SqXHFdh0nOpQg+8gPxhi+bKQBwfeiv6HCLTZC0V0dmwwrDu63LD/Ro3A
qmauIleoeT4u2T2moTrh55FLJEkiMOcTAAGquq23K5BPwqdqwTCnKrolc2E/rPYt
PzTq/s0//bPkzmjJjLPqGhtt1iM7qNITvHLT748fscbbbQSv+hCWPaoV8TIVB3cW
7vYqNANn8/8VsMUjkgLU/FZouD1+jDW5x36G6ACPkFvNv9no2+cMM+0xvTxB/bBN
R9Q9zwxLFoHzh9JEnZE5kAczfuguwNL2iHcWQah2zExBro0I+o7b7apBxZuO7veB
QNt44I5j1+v7PYrft4yktuEGWSBb0llSwZdUpQpCIt/sc1tweRSULKKAaE+kWXQL
2OSBxrAkCAOnI0T9F0NGeeMAmK+cVqCefC9dpqu+gPEBeTrBXLMNiXTFAFqbIBw4
NBoxXdguyiqArru6OFV77ZQr19vR5oQvJT3cIi6HLyv1TvZR47fDf0qTzHGMARJE
mgFcxvzPo46FX1wgkTMYfmEeJ+0avTy6L6BZKNkub02+i90gMhQ/bKllzru/5i9R
HEGxdKsoaRj326aoisLcwsXYNnEGcn/FcNn1TXBi0MVZOm0LyGh7NddpaoMXkqQi
b0+Du7tYJG/yD+azErKHJYi2qZvyYhxt6UY3FrTa88VHMSJ0ZjcI1d2o9OfgjUD5
eo+3eoSC3S/PL6sZkW5bZOIgoDb/ySzBpsJcKJqb7U4ot3ri7r3OuRM5GSLQg3jZ
uTjZ/TQxaPUXxl6hmawzXXTBoxcEv6K3B3iv2UHWD9qj4nKXhRElEM42uM3BiDbT
8vgwS4vMXfo7vZtqWaW/R6p6cqqh7p+hOu2Aux+xR6ueH+9f/4O/hWIryWHlAtlB
IiNPPBHbFwpLyhv4CiFZ/8xgw204g0XLDD0ovI3YWZ9DbRYA1qigHhqM/2HO94Vi
xhVdOkOfzplPzjM7Gl72kfQ9VnNf0HGldPRerTTCGX+TPa6qS2zFg2KzFl+y0I3S
5jBRaYaA3YSGC2xTOOY0dt8eFHWr8blC6SO98vqxT+JEsfBVx8VDX/P5RdbDgfOb
BFX2USX1MAqpG7nKdcJUnkhoi5anDLPpZcRB5BcO50rGx/ce7CtPUrGPvXnL4kbD
Mjr+EXtUf5M8dBWtwi269DMrcbK5T1a54fu3fzOXNoX4Do0KQZ77L/DElkkV+6aH
fJxtzD8/5qfsQasq9fUy7ERqYxtwcN8XuDUHgrnjpVdVq/E3N1SlFDFlIolwn6I1
pnsZcgIIJcjgK3V5HSbGnX7x7HzfzRm1rzTB11LZSfdIC1X89X5r/0fPTR2TC3vN
bCyi9o0DAHXlJGZtMKhTFn6CW02cvjLhUYshkxjMHwJ5BdKmpfUAAxfXUhRZi5Zc
t7m/LCQl7XViPPGsxj9MHSgQEZm04wRRtguU+bHNIg4FePGYwpJoIB+MVUzki0iH
6FrzzuckaXImJgeFKtdJivSbASKYeRhlGs8jnjDs9L8lT7LqNX765DvyFgAWxjsa
rf7Hyo/s6f84vCe0cPSaQ4cSdI7B4hdbCTbPHTRoIQNgQAyITgnqQbtpONE3UO9v
uekFLJQOEm1/GByBze3/M99LR/anRDa9BauV4O3bYietujBrGdFVRzjKu9lYzHbd
7MnX6aqU6aYJ4n+Sy9/h0jaZqWF3uK+AQc9cEzF39KEabgPRfpGduFPNCaXGpipj
jRwWz1uM8LDgeem8h6VV7fnB3Ni/wcIyb9ahvGwMcwU1pHKwKIXZox+0S1a9Esql
MzSysaIsw0099NTRwHfl/y5f5ct4wikqMwmTI2Uo0gA4dG4ZhUZN8FNzhvdyG4Hi
BhHckSNY4Jzur1iCfLSgCWNVBDhwYufJAO5ToZpVI9FR0D+Pd23GLGeslra/qaQh
cRieo83CzI//L5d54yh8okWghlf6Yc1LRh7GIHrnLXxJoiJb/W/hvdkuckJKz7yd
dbQEAD53pYPtCQN2zOYy27BUei9kn7uuD8y7qsS7N2NyqpCGEVvrxMYJPj8Ncdlz
jid7nV94rd96PGu6UizH/MKTHiFtvZLs22X/YcTAv5lJNLbIiJCnlPlAQgAg3yMS
sHFJuQfHsLtbbitpbAif9mO4/G59Z/VyWMD5GHF1dpArOphEIxoFmkVc7a+XeZ3Q
1AC3g6tc2UVJpuwLfu/YFcbytlrXob5Jzl9ZGY4e4AZtnkwBCbbSOg41oHWv7DBl
Qn9ULYjRGbCzm3AZAtARHv1ABHqi7spKrnxcJN9/JvCclOpX+3KHeze2fZk8v3tw
YRSz6KuNC5Y/X89Xz9Pqo2H8N/h4NZYa52Uf1T4H7W4zJF5YxcEJQG7sFyWPybb4
B68A94fs4L1L6v2gXQc1dkkThT8fK1/ZSaJHWN0SPP1VQJmQMH9UnhpyQkr9Kqu4
/ixDu9UW3j3MXXoDsccK0nj6iwUQ51DKqm0iA9G+5N4VsldXhz61kCkkRQSzwARl
8dCpwi0wSw5Ep54YoLGWgS2Sbtf3UCvNhKmxcTOLqy4Np2mafMbgqDD+LBHUwNQZ
2jcKkuQpqaktSxyOJIwpO+fZWzOgHHErF+kTc2NZ6Y3UcAijLyDaOA6DprPvzAUJ
BqOJEjQb7lqRfRZSxNRjQcReMebjnbxnc9rOHy4lnPnM/7M1TEUrDaHoO4vvicHA
x9SfFC1IoNOtmKccjkAiRO9tf9NulYWjVtO4ThOzhtu/X+uGuuBLGGlrI/Uqvp8W
K7synrcX9CFrTgBq1xcjwRXHdp7EWqyhTwFPXaMQ7IeCXUJqXfsJ5l1owFlb9WJg
7no2oxB4G1JJebi72Ul8V95NALWtkdnp8WcP3iIr1JOJFBiUwLjwrzGSyC4MU8Py
fxBkA3WTVUELYBaceqMea4qJ00/TVm3ycG0FFVv7vxx1OieMfIoKlvifHuV6mOon
YSpzgFOTg/hp/gAoKYbk0bk1K/i/a8A4FPjjtKrz89MlrORrL2rzpYPcWvt+QjJe
P/uqrvMeyy5vM/01EHRwX2x3TTz/FilONLYFJ6w9H6rpLgiYK4byn/g7G0M27pXu
81zutpg7GS19vL0SWDk6W9alsvoAd9m4IRhTMa2y3ysFeYi0DjVEv+itVx/meqcH
WvKdOpjhRK5dThkfHfbQtlvbBg3cctf2/NkPPNAFLbECOkOt08305lC8LHCYLnqM
McTqg+XpgomiQVV3B8qw2ZrzPAcL9E3ia2fCRse5dFy9ATSTJaMPJ8JKcr7PtU83
Q3SH82BUeAIh8zh581CGAOwbJqaQ7pizpWJO35yzdGTsyZx9JqctifziI9UWKNWp
zKe5uBfVAcyAHDRsxGHpHQ==
`protect END_PROTECTED
