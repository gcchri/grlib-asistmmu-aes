`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WMbswvHZ6jJQbT6ItK6+9gw8dkV3MtKYONYn10firaxKbhrYVR18TnXjjMytcfVo
eC4FtFEdiJqdHBNlP+5A7ogzlMPaPpZX6jEI28J5aB3Y/Da/YBiKuLersEwiPhQw
fpi5zHKGPArxG4Wqdn9qmhCTOdw8IRtX/+XEcQLIlOMAjGAAoo7W0qKh2ZMWOiob
0ClBboidJhfH/HySaGmPysPnbJ9tkYJkLY1Ia75+gKXcFn6UqQnSyVmwB/xOLGYP
sO8KZ/MfJREg4W3rj29KLPfx0pCzWMhsq7/ohUGIDCC7yg3M/f2dyQCrjf8cMTZC
ipTlgsv5duqIB6BYqFbb2w==
`protect END_PROTECTED
