`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UQzT0844bO8X69QnfuweODvh9m+TWTdXB1VWNLS7GXVZBGEyTC62FBwU5TJKVPVu
0iPsOl+LzI4/vCpwxm0huOlV7GGLUHna8ME+u3qufYAB4M8iTawukawUD3MFV9wB
JCw8eJrPOofodO2U0ZrnOVLYFfcvmVYxZI2i4AEIq/u1g4Mi1ZxFi1v+keN49K/K
boqXIMw1p/wriRjxXEAZkLKHXXBJU7XYN7pHdaeNJY9wdWbo/BnjDPabSqlpHlSN
2FeTYbtN5kfWHaXmMMrNQzjQLsqOhiPuIqWDzdCutBREYRywenHBOzaDw2XGnmkt
SoUWdStBFAnxOXmYr46v8RJAXoCpuN9AnHwRsL/PxOkCjKvr0jnpYnIXip5NMQjJ
tmhG6dtp23W3WuyPT3fd5sqzlovhqjhwPHkRIQDln4CLgcjgO7ZfqKElj1OJq7/U
iyPom1G/Q8u0BHId17Cri9kVa+T0CFIeQ1h8XApoxhujrnUSmstHFg7kypUOiwe0
eNo+2kl1ZI+9qDkA8GhkCO6YWEVRW9oDhlbyARmtpett8HUAItGKygxGkextz8nI
J+4F8zQ9Y/YCPvz8WPMAuh0CsnpcO21s7L61lSFtEMwyHUwT11S77gQgtsW4lOQ3
uPdRwsRu9Ii8pQPXNEoXP+OHzj0gDx223skA4D26mQtKa/JubRmiDJqBamgi8SEv
OOjI/zinCLMLpZ/WupuMCIKXrXvfd2A2pPZBB0ZZkuliuBjka6+St0aTz8xDqXJn
3rlSM12skUUZ3umeNmJUqt8urkL9bdB7UHfpIt/lL+hxqQfUvJ7ChJdLxtuOLx/p
FEFpSOJboVbeMQiqNhpfsQ==
`protect END_PROTECTED
