`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NKMmySvCfr+zX1prPxlg2itljaPLhPiIBv+UK+zt/0ROVvgaoLAJuu/7tIKAHrEL
3EffuZACLxJaw7h4zKKaCytFdU3vLjg/xkSKQ1NgMjZNa/00cdlq0iClch9A5TD3
3xGqmfLJQtCyhDXg/rZzhE8fJMsTrLu08+ngegJry2IKFkex54hgqBq+CljzaLmD
4bIKzpRpmgjLCTu+tz3NbfqcYa34aBDS84dUB5hiL6lN+NYIb73k1ySRqcAhcrAJ
ycpKcqhVYD3M/NA1CNHAvSeihBogE8ErLgZIsYPHq3ss0tqrGEUh2SadYRLElqIX
zPUVhqfYSCcMtGUqZNFe5GHOWqVezVF195YiW/RynPnCQWxckVOUdj8rbm0NuYzA
9vM/5iUWGG2ZQpx+rTYqxBmwJfbyhFW7/lYvmgD9Q+Io+gLHTi+x+9LAnEas0NVf
cc9hU03E0xQFjevgK5S0SO6ze6xsK2twduHiZebP1Ko8s0Q3ERM8SQa7Aa6Tqv4F
imR/N4OPUnju6G6DqrWSxIMLuUzce5qAux7IFsKrhxYKNOnjnWOOvNa1jzPg6LHt
lWGtAX0E2J9SvOAjzqMYUm21mvEcKroEFHUm1fp8EKfMnB5MWvsE6kaMpYsigeCp
U+6ZXVAEqfbprKsY5LKyca8FyA0sIMUsqblv8T5oLlkJe1GD7EKfr6fbdSGmRYdF
x98+I6aBqXMO9fML7Jkj1kcUYs8xKy7Jk2uNrSe6wGPqiSvP8qqDTn4yyVKH4F4C
UDMBwGk30Bop1zjxVg++daCbMy9osNq8UU9aL33MVujN7owZ4Y4c3J+q26LhifZn
YRRqtVf+vuPEtyqaoR31N8TgJWl7rW3I8RjDpDpA5w4Y3BSmaerXdQdd+3tk2MIQ
6nrbdqNSH6Sij9taiTH28tkVuVdRC+dPuE5zai+zZnjzwApH/liEddbVSVqZvMSh
QFcREk9GuNDY6dZPxzASW2v1l95rMMON9lSCpVo+zilHxvOAZ7sSz70vgqB2H3AN
KewXTe+3Q293luUQmlYLNXRs9ZDmcniL9Kj7u4J/S6eGyC+7fPf069FgfgPkWca6
lA1oqujrTFHC1v73koiNGepIySMcOZ0Yf/7e4gz0VO99DONtUh1eHH8Q0lHuyAab
DqRPsjbcLg1JOIJ7+qWQj1PiDwgyxfgXaAnTN9WcW+j98rlbe2mbSPvVcK6EIasU
FOTZhsx++JLXrM4tD/uLTBcuBCAVnmYDtYIurY2BGPBPnh5ym25xVV8DqUtYUKer
`protect END_PROTECTED
