`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Byh3wOK4J9/qi3C0NHICkbALxGTSGtuGv+O9JNf0yPpQFLHgozze6OVb3YbC2Ae0
c6lbr37WBBv/LEQyTg+y+c1VjIDqc2F7ySlcOb3cXdCoNOkeTA1dvm/oMq0pUxdX
GZDu+VrY2sv07xt6pDiNCC/jXPAT7/I0w3OyBt7+1i0RrE9nsg4wxNSN5r8gpPsP
CzASsZga6ctc5xaStHpnvxaqXNONHZOz0SUY4g8O8hOvRa7v0+0lqV682i7MEMFD
dx/u2ij/H2KfwHY6JcqJmXOPAjksBKJ4vIJUWuuQqDkln9PS8QtJvYYS0nEizXbu
PkOO3qiAXGlN7ZhFnsTDHdTGnrluqLVsfTM2gupZbECQpj4Tpa21Z4tBq/QnkGuH
5htH/sKYFAmICbQN6stBh+fT4Sj7nd9kIX9pVQ0xKF1P1KdhxZlX/JvfuZqdoajt
ucoj9uxiOnbowleRfAVqnR5ndgLo/TQuwSuCxDwVlFFl3tzSbhaWXyIjECrQydYc
jWnfOCt+UST/2Wa1LwtibszUS7m7wTDj7HWwb51fRlebXpVIGstJvXf3HTz5i6us
2zp2RVGdXcweUzwe0Gi2RkYgX4B/jjFJQDqUO55k5He0tcH2vXBgn2gFvwASfWNQ
70rHdiSIvDLWGJi/MEz3Ww==
`protect END_PROTECTED
