`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7j7CYSN2CnIOzBY7GhqMADvTVySARL+fvOwQc77e//CZHKY/CAkrMFRDgO3TOFlX
BJNYCS3iJV4jPNHrv0jVnmgbrkJWSHcC4r57tFTV0EWrLDX9iHs0Td8SYzbHe/+X
Gw2bKux6OQ6/bzT+uhLsULIRgDUawFueATdygbG6H5EkS883gzZ30gS2pWalOK8n
Ax6iGYIEoIMmhztj0SwfXRzofg+giU9jc9X/3AM3bSLSo4iOttT/v8ufv2Eric4n
xYfwneAK+1K4tFAhuZfpGmF+LFYIivWTcilJt80cWU8No0rBH1votpB7Gq8wqcFe
TeT84Bw5IGIHcFdcUQeIoxPmXcbGWIQsrcnCoRC1vsIgeHJEcov1KTu/dO4wFZO7
BnkLBLaIKsDOZSkZUMKeEg/KQGe2BLLcGMdjbjVOwpf2ij9KUi7KtwiHst9WxybQ
K/Gzl0fRrptwY48uwSqccZQoAS+7umQOSRwobdt3p2l6ZAMFeQWuUN4mdnBFyyFO
VgP00HeL42kbind/VqWDsVQYuDXz7M1LAHcqifwfJD2JFP85eJnvpFu38FretHov
vno1oSA4nEf0r5idBvgZAZsHpVuRdiAZMkKU8zbqcdxe2GKPwzuh7vkhZRiE8m4L
9fJ72QoBrdozhgijNpTj32YBBeENM1SCEhpIumI/0kNo4w53UrXysiqdpUAoBxrL
sQthznfOJM6UGswfp8ranw/+vwLQoE+wc/z9RhnKwdpUfzvT92q1HrhoJQu+HHtC
7GJRd2AvzWqwuAOwJbCXf6NIJ+udFeUIeRaNO/zJHuNNbc5vgd2p92Z8bqdOLjNP
HBom4pR6RfFFgq+fz1JHzk0eN8F2Wk11J1VEYs059M0=
`protect END_PROTECTED
