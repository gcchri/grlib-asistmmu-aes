`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9IZ2cBxdesgERifYKkVo/sy0/+K5N5gDfzV5lRUATgrAQT1tF0V6A10wURY4GzIT
FwknLSG0S5y6CesotqGClnx4lM9T1ZYOOkcu9uMN2VaGhMt6wxs7yNBGXYETsIw/
ktRk60M5QWFSrJ5fxsTwQXw+LwiJAWB4BoswgJ5W8nV7wFGUxrM80DZlzUbjXofs
+o4t8fpPaTCdWgtBn/d3CPtOhb/LcxxbDdYbYdcxk6gHFK98VDvqnmZ7u8zvl6C7
AGdj51Zih8Ilhmv2D1OKeRidsyqdzeHuxQdMeRkm3yd3641evxNwDIXU+BkRowFZ
NcYQWxSGVKNH6fWf+ILlr36blQNtGtWo3U/F6Ti4aGXxoWk+0WSbin7mQ8m4OCmZ
z4b+YVMDLumVE2YBFR63TWAtCX7DFtbVCaXHTn5mfjmE1Gqssk2aWqUexWxJKyrL
mR5It4yX2jRv3AQguuY4XHMaryXtuxRJv1ZtidAVuM0d0n+55Opq3athfdEhG2qQ
GsVPTmQ+kG02KzdXzcW+MTlm233WGgePLNPBj+7bFJiQ0RJazS/z5IVUuWYjOoG+
VxBBEBr9glOSndNXFuI3Lrjn89uheM3pF42rS5y9xEM=
`protect END_PROTECTED
