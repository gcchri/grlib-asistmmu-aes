`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iFFa0M5n4bKirH1tJjYif50UCApnR5dvEfXq5q2hGdhb6nHDOmKfFnR60FXvHP25
LL216BoQebPnZ5u3QoqEzCQRS0rJWnYQvpyqbbpC/gYG/hTd0Lymck5zFMshajgG
0nfmiM/YVwXbyLFu7gGgj8ON7SIDlU01+u4d45k/ZBMwqq2VmzcLMFuk/qRlztyX
IPp427Uy9jPRxb5r38GEG396ImLAs9aWbKl8j0EV/zYC0rJ8xObtZEJ8IWU044Jg
fIPlRF0zv3SqqSSmJo7fS626ZY346fWkKpxGw1oOleAhlykP3jMVX4mUF6W5Yo/g
3rVUYiCUyrFHLAhhfoyH5aJdlGK9VknJ3QCsSjxyOM5K6sAHZg08Gpk5ACVirl9+
WfFkIEl+I5lSPLDvthVx4UT2bssQz1/b5eVObBpKESg=
`protect END_PROTECTED
