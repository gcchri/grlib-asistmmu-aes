`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Abaw8xFP2AetbwrA5H+h7IFzkcnhMNIc8gDA7oHVPu9eaTIRE1oll+GRg0KkwkoJ
0+Jud2MmLwg6UPk13abv8woh2HAhJX1lXcaaZ2pi4uX4ghv/yT25wKoMja1aXJuT
cX0eYSxb7XuoBrNDA/lN8xTv+ZUeVJ8YjaCWzZDmeNe3fzWznSxK7k2TZQwj5005
H0fKEW+0/gj3fp5VTska3xTxvSq2tSxBkpQoAk9MFKF7uV66dke6MCNchRy9BH/X
OqNeiyBr+dFLw/lK8sfS3kX9F/ARII6PuCmZe1G7QO2gfuBTFwPGAoYAZEp5Lzai
4yB1HXbQL2H5J67u79UozA==
`protect END_PROTECTED
