`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VPB+w+mWGkmOmJxBl6ORKq7vwORRGdtIRH06JKt7Ki6UzvCh2UAZxv+g69HFmEp/
mp9eNZIyhHTJuUZqDVLLvOqlk3dHFY+08KqoxAzycRJElXx7O9TKbEGCZbPgGTVG
OYgZk8J2+NTsiyaUVNCUZU8sFB4OinCQBkvvF9gG0p+Ek8WUVybllINX8HTPwtD+
ViMnOKNc7V8rgGpPvda/aFsLnueIqj9WCjKZ8sdeFVDftXom2WhICJ3xW3dbKhiE
Em5rImQAd+wvG0QxBmkzfFsdCPZ6dbyKWjZCW4XDD6URvpMxcZ5vzACUW+/cjcUT
M7Ql5cjohbOUbxdinbnpg1+GyY9HGJiryxnOfO41jCRDTY5AOJqSfl5m9gFf8Xhu
uJDU9hXbL3Aoc41ndT9CZynHPCNekKjPvDYzTl8ODHxzkh1xy8J7pGOfz5Dd3CGi
GNKtas2bZ+i1PI+pyfR0W/EfNbu/H1VA6WbiI7WoV88aAjbLNn+4V4jCRbsfhaLR
fTQH5cBE+XlBqp3pwvVRR0q7ox6J5giRiPCj0qNOodGM2amAsUUZJ76uw/O20nvo
J+n3Qnm62zO3ZZSoTO/G89fd19IqFkno94CQPv64wiyqVHm2Nep+s3muMX+9yp8K
3/4DkuvcKv9SZ61/mFu5q2CDzdqtwJkaRYcXcMl/VV/X1SaV2hzoiaimDzkGZFlP
zyW4vWBiKsc6TyR9JQxFy09+6a3sRRW0wKKkg8whp4G1LXhA4gB8BrNSOCs7T9vJ
oKnKSkwNRqmCoRzKF8IXxkFma9ICB6bbNReXmOrxYuQ=
`protect END_PROTECTED
