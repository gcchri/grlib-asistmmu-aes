`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zfclobuMQ1077Sx1k80a8sH8NhvSFyDtl2LxMtHkHCgoOj8ON8NvaX/d9i8HREV4
C5po1vhOZ+d/da7SD4H6lvpxn6VQZE85rMKXUs/Q4UFkWYICEw1DD8fEs7sOpssR
zz5mrPfVZMaD8l/GjCRi/TfjUdMbtTqEEBbOqN7c62NgysB9ZRTCinDCR9oxR79b
S6l4gqGC3FfsdiGbJ1XbnmsLLJlYbtYA8Ph6plMKpuHA636sLPihdG4zQ2AI2L26
XLNpu+dx5oHfIc8iElWFYrRPCbIm5pox9v8GbEytBomN+8R/8zKpTD+ryAVhtGdZ
TFV1iOFHTbaa3u57/k6I48osTBgHHLK0MdytMB1XG2/QPBWcc8sPl1Rgfx5y2B9Z
HJoA71CFIFX3L2IhlnoXkdgzf0Rcr6rO5m4m54V8EFarE99vZjyJNemghvWE8R7Y
6bDZAYtHyUOUJHoThCypMZqKbLobXmazFZvk1AIDKik=
`protect END_PROTECTED
