`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DYTaw0Vq6CJW+sPaMkEfY+3rmwoyvQ8Zp8sHKEDqfCr54Ysnw4mheDOpA2oTpDra
P5TUMbPM0DtQJ3DWFqkLc79qBbCcTbq/V2It82dh0z+T3/Tmd46MfdBwdrzXsY8d
witibMaCWQDFhNDA2mR6StoR8aKHRQtKBNfuuzUWpLVv5QersfF7ewOMj5hYRMYl
MLCi8Qxd2V8MpX9j5/YTQWI6y5SLz0TRBzxwWy+7lYteWTSyKg+rrhzjas5Fs7UB
FSrHVJ2ocwo0RTMHIXZUEgi/pifBeBZfA6PkmgIC6AIAvD4mtgpHcW264hTn9PgJ
Sj8O+aOuUw6hlhs5MHtm7NyMi76hInhf88w6/PL+EgobNr/OsI2noVPz7eVFvDDM
w2dJteb7wxYxh68+cc1sOAT2as/AMA44xRCHQ0Ggo43cmQZrXbuNKIHKoAzWaGgN
YZ6fQ8031jZI2Gz4/VQY8g==
`protect END_PROTECTED
