`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tEaWrkoO9zGfJZpPn442EDBbgLT3fmCJdhm7dyHQKhjxF4va/rKh4JVzyuUcdhTv
DiWbZmC1slmfLUPCbM2kUpXwsWi3WI3UZyZZD0ZpY6Ce0PDCeOMbdu9MV2eFC0UQ
I2PtwbP51mvN1i7p6OL50hNYKd9AwEWuv7Xx0jYKn0cYzmW/OYuMfqCl1pQm6odf
QtsJJO2iNy7JK5HsMXzd6XbYJ4/CDqduRZQABJzEbJF42wYs7WCo8KJHkJ3o9H/A
tkXGP2rOSLPOYQcJONAqs1FfKKL/5lFjmZDskNdoexd4T6OKupKJTLLn+jVutjsY
6j2w34Tgs52yYReafPUdT6nkeoE4h4GhP2HLXAQXK3LW5YMLVtMxiOv6CRzU0dE+
`protect END_PROTECTED
