`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i9ZqP75gs+g1RepU2kT542tzAyebEchgFw8nkMok30U/JncWs1UxqbBavDzWg/sv
e5zpMdUqRB8gWHppzseBqqExe2ubkaRI9NmxLtZ1hZxRTNYy9rm6706QpBZV4m2A
l9XY2Fsk+Mi9N65kcKKIoJe5+jr0Jh8lfgyGuXgpyVqemQuCjp/yTdVspSoRDpMO
VINUdrzHaJNf2lIzDvkDtk43b7hYE0Rti/9UA0T4h2OjnTcOikuECYALNDam1S1o
1HoYA1L2O13izHfjDkuiE9qoVwSmHOvld2GY9Vr6+jU=
`protect END_PROTECTED
