`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m/W81GOJ8p4MUrgm5jp/SBE6XsvR8K4t6NdcRs164Dx8QMjXtKd2J/sgTbWAF2qb
V9rFlo0RUEIuE1pMZZ9rWNC0HNNsR2rH6zVeopbVKeymdcnttCB9DI9z1NdqvhUB
2F4kbFy7HuLjvWbDbVCjwcedGmwd+suHMB3dp/T6nul/s/2ksu0xwBI3AwDdCmTU
I6FidNc9i0w9W12PaU/tr4Fuqix+C+F/dMMRH+rEAbrBk5Am+4iI2yfaLHe+h/Lk
AzMnSwWiwi9mI7zLlshBLzIbsPhrN/QEEND9ae4CRfrMxZ8rqEHSNPN3zGVSy13U
dAOywT26aazrefcX6XHaeQ==
`protect END_PROTECTED
