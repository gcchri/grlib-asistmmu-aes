`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y3rWHhcZpQgwQiGQKrcY/ofuFt9IENV+5+RJk6cFU0/QVAs6mn/k2QU+iwiC7eaN
KoYjg4CAgDVNHJaaZT5R9EdQZxDtfA7cmUiCrPAgmkbCTds/a4bn7dqPOfNrgHBH
nQzdBibGy1y5W63FmVTm5DIn4u3RavcBXx9nzQjifntDzoZtcsLgUftWw0tvqcQj
MWGNDlcgg+XmhyfepSlTsyrLOIpVHog3KQH5BrlT+lO+faNIqyF/+uwuUfVUBSuo
u1H3tkMdDsLodfyXwHFydz4/fnH/OlvLDlsS/s8DPWUYPlQKjvMcCvx+ukh1hL73
vpJtZnUuyeJvAvCwegoYUS8JxKvgF81HDK0mE5L/FpPRTU9+/o9evFcXuxaK9JaI
DZ3x/e3Y1up7hO2OILpDtI9CnEO+WgJ4SPJi5FEBOFwG8gzskrK+h1LvQE7EuY7H
Y9Z8o2WHwni6W7ReUZpUsiJIX7oI2SRc0yGUfghMPQawEOdi94JkWb3PO0lk6lc0
ry2BcfEXKBmW9l+8M8j5fOSMaxNO/0xuk1msN4PSbax4nR+VqKKdOSYmIbCQ27/P
Za9aH1c1wjiKU80v8Ee0/xBjzuBRgE4iyIQm3mTMUJq5ITtKNNzFtYtPyGprBIA2
vcH+eX/MEUCTtc1o1mjlRMxGkVGsJdimdS+kXq+onSPLQAOUnfvmNODBo71wCveP
6CWQ1t6oqa8vMYj7b7Qb145sMjHX23J54wJlZkgl2ULmcxo2ZnZVoNpUydthQqSi
ykenpYzeIWQfILb5ABKIa3f0RDAVeXjtCqxu1N83ARcCkaXoFt6z9nKsYdz+sSSZ
5qGe4Kh0WzvmLmZQyPvpAIxG0+X//WZqdo2a784WFqzr3w1b+9yjzRFI2Zk3pg8M
6qvA6KKbef78S8HdgDqRTRdSdaaPZ2P8LeZNWaw6RS83HhYcNmB+wAwRZQvzQ0G9
YUj+OtvAPvyRleCWBOxf4g==
`protect END_PROTECTED
