`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lgcp+UC9oBwSfDhysiw71A+LVK2V8tJ8G4Yxrwro/9AEmUuFQoedn/m+3jHYb6ve
ZlefZU+P/YiX/EhbNspC/HQ3UvzipoN/+Sx2jIc19wdNsCzHHH9VVJucVUwVVKp8
nan1XtJRPR3HqL5k2MXeXXFhkiNfMZomg1rC5CKyw/sBdw+XII2GxzGZGrnw2Auw
Qk3bwhrxH37uYBW3SbJ+H9ULWAX0uuxWVC8NzRA92vX1UdrjwR+7p7PoY9/yqpZy
s6t+YIsLseSgpZTIiXU09SNFWFZUbffZ5SGdElaZkkj0nbLaPVxD5UZ+wYM72K16
OUZ9fFRHS1m8MZM7zhwh0NzpfF9YVg2AgBAun8fqK8ADpwAXJG1rXyZgxdHmJJ7S
9vvfI825VjKH+wX4ZE/n4DoKxwDSjAGf2T1ntUx/LnSbG7gSvRa8cHlRCVSsIdAO
f+Hyd8ia1k3s8WEmc6X+p6qnQEJFk7XsG7eP9C+t4QUM0HtCyF8dUPc1MCvr8Dn/
G4AhLc/hmHF9o/fsFdVuC52m6fkErPisFKIq52ry3DZtGiCgkYS9bzv02f4QFlEf
jKlD3m+aJxXPcgc5mG0t6tRTt5k6uOLjkpmKGTZa234hZ3+fgmqGBpdK+lj4996U
vC39ahhRY3RkMcmYkyofoZUozWM9vGkrudNilxAJkqDHHXzFQDdNpJbZqV1TRRHc
wZbe3ih7zWGwh/lpb7S4FVMlApcB8XjCou6BjOezBwGEEuC4COaiWRg0/EjJ1opj
d6QJlgrg0qELnKC2kMJ8mGNdg60il3gT2QdMAearEbm1qIm6ByXpVBFKd25ru7wA
pQlRJBFlCJhNH6YqAgInPUMlf+EroR2Je7YgfbCrE4w6RtA4vNcuu5HNftr5wu0a
E5GXiIMRfplKWehXgl23U4LTaqe7XT/a4wjOq/b8DG9TsVCaqsfBIB4gDCFsz1ga
VauSNlzhzBadIU0kndow4fjn/iy0XQI/IRRKv/Sj3tEjTZE/+JuOviw3xFRc20Mv
s1wJ3fBOyptvmmHIlDQwQUJIecYHnDaEG7uBZwiAaWBtagKDTprFyg9dUWlB5tsC
6QvsX9wzLkrMc/URTcriu/41HAj1wnz6NWR4M7jvUp2FfQ/NRGAg638OrQMUIO34
i0SigvUBBj7f4+qY/udyA89uvDfFPIVhlMuYvt3WMJ6qN0eWTAxYjceVhv5Or2XE
wSisY7Wt46tMgAd85cEIH3LhB7J0bZyNRW1XPzKeWlbI4y4V1V/zaDHEfmQrhJ60
tvUDPZXjwlb6SO1lfmFCNTYZSImpV34rYtY6sjPlvwzxY/w0T6kn9+FPn8ljcLWh
Ck/7PL/9tRnTka21/NV10SOCDprzpbPq1NXBrd3vHMa2SB+mYMMJF7hzMzr9fK4I
5HEB8a9OXcSiRHr3S5gJF0IA02tmscaJGNu9uRv8XxquPPxm8650SAjAkk3iNu72
lwsu8iEVSH26wrBlVoIhcNkOI4AOfm8e0sU6TLa6fotRnQIOgmdi2eIfJ4hetWcc
8bNfG0WQrhn57Nt38sEUo9dVKmry9gkrJyJBy47X9vS+eJ3Qvnn/kGPKEsvyqKIB
Px7LPIWdA6n9C6cFKySmfyye1fwojIbH/PCuNzqwwUpInh5R4U8MlFRvE2PbwNhg
GF6cAtlJQETctrVj8JnfmuDN59rNcKfN9n/8lb1chU0SG96oV2fzqboE24KeUMJA
srX0B1lvlj4eCT1GEUpV60Ihgk3XF+9pJ3MrX7qoh3ivuNuNzwZIr3AE3bHRJ+sL
50mrfYG00N0J297iMDLvXg/gFinE/pMcnZSIAtibT+1Dye5lSQa3t+Qq2DEx6Mkj
4HABzx+2MSL0ISSc+3+7JIPR6v9WTPQfkF0AIPZ9DPZDtnmRBkAcPZFkBZHA/hqX
eeBIYh8Xa8qOpWXkQsLS8woIl2pHCa25UfAambrxIZsoMF5vzvhWOeM7C+3+Lub5
g9shIQ4bRFyr7OeuZVbedUCyvMQyICXd3gTtTtf+CD5QhjS8ycNuyVHuia44WL6J
AXONOhUTINEKUdT3g+i/nP7CKAmnyJcyP8CX8jQdzSAwRr9+MBoCeNkg1iTLxzV8
WReFwayJm0WKIouhbbtaFHq5/2w42/vO3FCFhxCHvjF2Q8OipKBTi9I+JMqz90pU
JFadLOhUYQ18f+qzkNEqzQqueB+obciGVfb1OSgfFj7+epM9+TsN7fEDICMupbnO
BjSB/I515d/Q65JzGGR1vXF56Rw/7nzRus0+bJ/7/G/TLcWRU9FwYmijg6SDmfin
5sh8wU+pgODwbn+vbGnWhS/wduebLFb+1VkK1xv7pWkGIK/uZxUVpAFAw3psa77Z
llRnwyQ+UwgDnxZTXqjx7iiMmvYAlYKKXuO/UkCAXoFKhZ0qZkIWv7Gr+AlozZ+T
0YHuER/ndcZ6iZxKdEUs6namaB+TFFItdf1xN2Cy76jWY5EqjxbwUtfozeABm4Hz
/zJt9wpIKjrLxIRlxM6GNHxM8iN9xCgPeEgRD/TpN9KgPDxUwahWTKxEqKJwz23q
doBKCdUEf+AOk87cygwJeGRVORgXyak0bJmutE/8oQ4ozrcIQNXLm44ikxF9bxLi
diogp76BJ5546bg/4IzWfrX075K94qoRdlh4FXI2NApoc0mvCGrG0UCtjUIP1HxS
S5Il5GtW1Sd9zm3ESnvrF0V5sHBwiUZEb2Fm9gnrdKUEC0N4YQticrRXUhpfmVa7
je6CQUkEdJZQvEG+jsnrlc9wY4WaPl1sPPgfDQybiFy359nYjB+hHieX71Yv3hmt
XQ5MAemp7uV1eZSE5LayjBNsgJ+bnkJzHVOO+hML+wmt8QaPFV+AL4Njb0jsppQ8
0dlpLBVR9pQLqa9QbywCu4H2WouLO+LcvGul24NdTPaSYfw5LCVFjAPr3XPuo4iz
+lpsPA7m9oqKifd4Kj0ni1XLnU3SwDDcIhcTYrbqiufYF4VnizascvvZ2FC6dMm5
0u0v7RNcggcd7YGHhNw7ZMQ2HVH2TwWkLzQ95bLIWCTxb6agG6KCPlAQp6Zjm9pP
M85eN37Ev4KGNsekx40S+VC/16jA0gEQpEPD98WrFYgS+/1rim61cJwJ2D6Yj3Q6
BAFPOuoy7q1gTWPW6PdmbLY834KHTWIKwNum14iTCYqr+mFMbkhNwQKvh3vnKZFM
7MF/FWVOjADy0mUMAEmPPFjdfjDK5N1jpxGbxTnUrmaS3MSDU39RDYtdvQGhNXq5
ipOmZOLnQ2bQtByytwkWgLesLcGWXBVZWevtDAy8QWeJoP+lc1B/sPOz/ZKY/lJh
OLv2fFyZMTWsR3OqTDYQSe1xjwLH3+r9NodeecmO+lb+GpD9tDpxLjHnJy5loGeB
EKopcqY7bJJ/k5AgamWcqRuw31kUUv6fpxzOtSU1zR6iQ4tJ1YbCb9A4SonpxTmP
QUB2JJ5BosbRoy+rQcgfVFNdyM9fENZqzzR/ttb4muvYdHieMsvvWaOBIjVM4Y7+
yURKIUtIQmcfCyNEJDgJyRs/BqKCSmqfiUusSJwbA5XNz6d/PvJGzZHoy+2ht3Eg
RN8BakAfDryen2t3fSnJKmE31ZHTZIjAc/nVcAalQUfxqnHMVH3czNB1bun3hC2i
bPxVHzGqbrnbGlf+sKc4BYe6N4jZWIpwEUR7TdktfpcRRFqhlciZt9Zsj5114VOO
6uh+zWqe/coLneEiEMCQgtAS8163l1xNloAiUW/Hr4h+nYwa3GThLv6HwpDjlMBE
d/VCLqugM+Wz1eZIV8dmKuYVdtZl95xGaK9qPEMhYQD0O2IiRIa4u8Kdz/iFDMv0
ya6+jKlPtpTQfwwNtGIMstImXtge7t6HcKQaHWoWXFHSP3lZh+6J8GypbNxTA4kl
iST2Toh/zYD2F1EHW8QrY6V5hurqGCqvL+B2af1BLl/abzdvN8QCJ2mVlLZXLPJs
LCzdyzZpfBq2EdzY+04KzxBSpIyf3xVfwt4Kd2RoOFk7LZPjMABD4+0IAlIxi7+D
iNoD4gAa8RnBpLIew4YFJ9+OTIXvzK9aWo04bFAX8ZVAJCC3FN1mlp0dmIkItATO
BnpFtoaZf/r85WHebeKczyiRcFDFEzea0X9Q62g2c45PiFCaA8V5K1l2wV+yb0lo
1FcDArSLUt6l4Nl6qBv01ydkhcsT/eb2r+F8pohG60yaICgGaMWWvYrEKC2b1qiy
sxZX2bBZH2+s+fs8pwDkCKlB0ytMPDGdIEmXJ4bFJjtACT8BTVJiGcKSVqI1PPhp
07CnGAfw/9H/4eRGB0ZtmlqcRHa14n/luxv4jaXLK9nswKubEv+IaYFhZWtFwHLZ
qHnK0o5sc9UJucBZQZGLLcOGOQGHxszp/6qCPc5jlWeWhDzToyJtqKC83YUu+Knp
O8nX8eNb3Ns3+FljxnIHPdUHBWVWG5ATl5c5nKmg7HwAJNZZE1Bt9oRpuXf8LmHg
jFUJfwm+mMiverYivPY8upI+Ma9CIeMCRGpITTo4pBxZ59Sug8h4xQqo1U6601/8
F0nNcYvTvXMIBwxk1uBVzw==
`protect END_PROTECTED
