`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8GhdY/4WK4nyIa4whNGUlATvacZ8teTLgmNIAD6etzzypX3hOgxmGCvX3/piKqX0
S+pIbFQPVFA3/CcsngEK67e7y3ciYb0cruYhzX9dzWnaIc/FhIvyaTAVelKbhWYE
kNgNaepCpxVZljedTUgROlJpmU9SIxG2I3NbK8KN69yylJCuavSnggpJodgdlKZ+
7xIlfVzBdxh1feLJhk4PsNsufSe4aBoqcpLveZoSCE0kvX84bD/F4kyR2WKcYPso
ZlcIGjlXntX+lvVuS19YlCoRyzhnG+ZoMT6zr+ZYkeD79uKYMbGxM0/+HzvvuvfM
HCG8vbZy9IIhquZGWOmNSA==
`protect END_PROTECTED
