`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eWOXyHBBU3rPWJP5Tnpit3cb/zHUbX6H4+MZKg0OHYT2gFfL7NHfvQUwHl4PMrg7
LGPczGy4Mx240KE3vcbS34MqD3NgXgyC+OJHfWT5+LzjWpEImqtAdDg7shpBpBwP
5Q8xp716bLy25sXIPIdg+Cgv9wQKELe0n8y9Sgra6ZbdDHCMRCNOjcsKvbPBB5lp
U2AS3eKP8P2qS8F+CVS5U62ywCOR/UO9eSoPQxNbaC32QFvTMpYQ0Ey1wQI5vN5o
H3GSc2ro6pllNiuy1FsX9d5OgzrCLRC8+JYGNKl5S9iJouiklFSFiConsmet5zhd
2RU6oZqpwengl4nVLWY+dh0y5fzsF5jg4pNNqIqwDxuOGg9jwn6HULRugb06V8KL
RW0bGMTRvT7Bxbzj78N654T6WrjsBKvDSeAbSjlEliM7tGYTa1aM9mRkmH10XhWC
Y8ZYYREVimKx2tGucDDjH6iG5cWkxq1uCSo4JtVIAJODc8sRX/oPlbOqV7OXe4jo
DJrGmK4K98GTDsfYYG+Q1QA7IRk7MzgdafFsfx8YVDJZku20Sc4m2LcfEyyD+ZMI
t/eIzhhcEY8vPwBMr3IWwceJ6XKKaOy6DbdNAaFBoTrwtkanpIkZ1Fo5TTtPOsfA
TKt1/QllzTnwHP/w56ucWvxCeQhOazJ7DxIrhFOAaEoJPd2sAzaK3PtEzoKzH6h6
8wwr2cbOAXt66zO34ftWNj2q76s7NWE/B4jXeWLBGwZYJbkZSryRiTsy0YmL7++V
i2jsvdvsuIKQkBkBnkM4WA==
`protect END_PROTECTED
