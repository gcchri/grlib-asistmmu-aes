`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JQwPpFD5hboSR64CcBh6ZisLqhsiyPfW5YABQFAfTH6OCScFCtQHRwxI0IYqC+Ef
H5ZFz9t+1ApU/1E30afm4IexIHlEMpFgGeqjsqna6vuh1fntvICQOfeJTBkZCILb
ZGC/Ol1UUenBHuu264BBFUrOrvRRf/Kexjn0kglL043cXtzx/ItGrhAzwzh2e/6n
40Wc9tvCBulMINSel3ahnW1EcvxcpZ0RZDIcieandKGL3VjoebCeuOLfmBitc/17
oH2ppYao7AWqlzLpRPOwmg==
`protect END_PROTECTED
