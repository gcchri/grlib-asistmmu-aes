`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4l1QdqIDYDN7Yw3kw5AI2JKcIdHrkoywLcQk/+LcfJnIdns4peO/GNj+XXgiE/o2
ctXE0nuOkIQKHHnME+1Holq64IP0RRVTMU0OJr3Zwum4liXdtLBodYwLvpA2D/Ep
d8Mlk3cX+m4dwfit02kAaxqpSpGMTJ02jGR1SMsXAfp+HqGPJ4pVuK5VIgKbdX18
0V+kFbnfDi1yqpx/K787FAi10caPj/Cg20tFt4+FPIuoEm9RbVsgc/9ohbWGAQQv
dKwAHCwDdMRVzL3zpsh1Xg4COdYjdWCXQu7zpLvAx+E8p4KD0PyHRPJ+jnjPZMPw
UF06F9pwwZ2fuOEPXoX7mBc95CFkDhRv76L/pUDLmreD5SLqymsggsmCPkHB/KNH
YPMjxOUc3LJgGBnH06tivnVNalcJUwcJZ3cxZy2Pu5fmAO6Ey4sP/jhBtsJ9KUpT
MuzqB44SGRP3Fwd4PyP/fIUnfUdkJBPqwZ3U7/xoLl4N4AHtnCtlJTfGOxfFVmAx
pdUAp0z+rbZiJjiSszCnQuuxkoCRbYde2qc8U1p2H5LEcCt7NaS009jgm0LenzHN
it5T89625+INjW7bwSpgig==
`protect END_PROTECTED
