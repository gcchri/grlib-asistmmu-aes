`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
npAqaZqxByOvh5xnDKOCZ/41JIpLl/Hc6Fnwi8KqYJmqlJNSklM8xFXjevM4vJOd
+QOqSIG3fQM33TABiZAYX8cRbTYKF/LUKNZVti7inHqyTZHMm9t78FFtD6tPsvup
90HRZJOtpbrVBcLWpZStRajMgcOGZzP6SXG0YBzXt43pGx4O1/VTq8zCH+5JYm98
8caO6RZQkold+2MmfiDzFFtdUNp+gwz7om0um054s+3cDHsX8Sz1XTqHQWUtujbb
W0lcIio73u80semT2V0gKUVtXXqkqSICrcmHse+dKhAzAX5ZDjuRBWu92lbE48h9
e1/qk8EA5NUw76DDZYv+W+g62e/yUR7mltBYyToRDF14THfsiSN7hWngJKq/IdTm
2TLBT5pvhtSD4/dCT+wju/NkDFs+bihYPZx6JhhU4FQvTo0Hwdcgn7b60GjVeGem
G2uqLhZ8PE9TPuArhbIqJqjnnMypzGzHQIgzIKHIkB+J6haTLO3CHpRsSCnyIVX0
eut9JZ9ysUvc+9BtH5P+lFrFHm32Jhz3y4slyMNK+P0AD0g3e32Eqi8WopljaglQ
nwC42b5UF0s85ZXd84umXMzo7rCwFGwqhQJmynM1rUrshLZpDjWQyrFythK/Q9Rq
eFnA0EW88FW38VghRulca7zZBrMP/kc+BCkPZgWfkVJbn/zP2A3qJ3L7yNZYvCRq
X4dooFiJPKW1ZTs9DEybHsWAIzEOZGnXJ1fJ4wYMoRL3/dl1G3geZQlDhCxYH+dV
/mcx0ictYWnvOUK3SquOSy73/hGvdb0T6k7Q9T0Jc6Tpbisj55+kpEvpIZwf00qT
UdJSA3/UP1nWY6uBR3U+zIJgrLZcICMDRCsZtRgGmrOfC5rDtcNs580ymBDYYeTC
lOF+0i4q/70urKol+tq2A611AZamrf1swvwSTOYFhecPuKUhudIsot/CMc8/jjpq
mBuTrKs+10aHF+gzpAP0Yh6fQbGIHJ0Uq28K4DLRWCB/1pAZnTg3rc51Bkq/GRDu
`protect END_PROTECTED
