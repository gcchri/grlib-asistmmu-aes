`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lRQpqLXKAzi1i/0n+9TTKJSvwbkzIqzP/pJRl7SjjcMm7Jmeke0PyqhXMdi/MEfY
ISRo7wnsocov5kX+x7QCSjpdsB/ixkoEzwN7yENOJcyclyjVbVtC2LAEbNxMdNSU
g67hUy8jGEGHsXCyKGUlc8p4T+iG7j8G9213QFQ7c36yNL+cRaSTNVkLqVl1S0N2
J5Uez6Ify3Wdgi1TToS8LvzD+Uv5JlsZM5K+dTqzZquOEc8UvUkxYkfl5Ghr7EgW
E0R8w5Y2iopuS4991xRjEj5vHBVUhO3oSy+eN6Qsa0xP7HiKB0A+Kp3jKqc4tgHp
4NeL/c6b+2zn0dseMS9vbzEvj3JA0sV5khc4VFyq0F156sehRjX0IIPolY4GmzxW
abVPotc+KxrZSuIN/cCXHrcSNuvhwzJ7fWHf1A2AVhmqXAAsVUlIdm0C4SrTIg10
4g3pkEBvc3rpgFpCK4fzQK6RmLgMSVJ72OoYEukSnIU=
`protect END_PROTECTED
