`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iHNljlXCp8fTjQCmFRt+GVN0UN6ZgBiVj3HPbOqflbSMXodUiHcajZ3uRcsYjxhf
/bBFsu/oiAd/MJJ6/nG/d1iHQwJktqOFNveX00XeqgXQkb3cm7NGjK9ctnA7I4wa
vagk0fNJXd0cq2QnNZZCY2ikVvAc+VjsibqnBYX7RrfJb5S73c6lRRi0c7Fcd+4W
3ERR933AKlKKn6m9NGRn/ldcy37t4f5BBFMbHwriGiEdGRhCA3duh/Jpr3peo5GN
2IcdIB4Y/9+8ogxzT84E5odgICFAw5cbfLRAn9sTJKh94Cjxe7H9jy1KoXFNhxjr
hutvajscI83xIi6SJPFH5s3yfU1LWIfPNCn18yb8B6fmQl/NGX6MkhYPf+UJ8fu5
Y0r2h/ITHpyoleqzjiSJ+oI138mao6tBzJ/ePHN9murh0jCbT7TihyZggfBDNKuI
Noe4WP9CH8p7bel97mRQ/H5JMM8QQL7HBK7+HC99vZyKz4LxtWkf65kYhqaGQys6
ODfXb204FEhHAdOyl6pXphUt/t5fgKrvdbYbLsHZiDcwxdLUW7ekaHFM84IMxssK
mLVCMUu1tRnrfjOk376PE35q6khJoCjkFPompxWgxLLjBHMwiUtTQFh+CoNt5BaP
xCQz7Amzp53ByuAKTMME1Zo7E9dtk8sCePpzTlbREj2sd4S04Djm7cRYFPqAzP5d
pEdGIC3mR5DQKpvE3MeI6r6RbJasFpdfKr+8kZcfPaKDf7jQX5tC+uYBCJnao8bp
ly3cAj5ggfCgpFvEMiFa9TCbExis2UECl9L/2/tk5kXVeDLyD+j9BJBhx6cXN18G
Qyjbi0E/6Hbc62PS9fhvdQ==
`protect END_PROTECTED
