`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nkA33VFQhWDFk4ijpjxxhgDjHQqyk8LxKRLtzqHJr6gPGHxdYm1woMJFeNbySSSs
ZKE/akPU73Nrv4XVcthi349gmNzDbWVB39F+1JR1lka1PP4cblv0KnWokT1vD6TI
h/EqUyXipNr9CSrAKgR/0elJceIOEYEJEcUrCGCiDZLQi0/gYeggEBbxZReaZy0i
0/EK+NZJ6/l6pwcdqk16D0mlQ8HD6S/IDg0koDBaZmG+/p2J1O4pVuVgKGnV+cYk
qKZQ9IzPi+K8QAGpVYs+BXBs2KmCuH2e+y4KTuljUT4UuQiyzgDLSz10gEQZAZu4
1dL19MmS8oJIGv3YE90QKZMdWYVhnSE+7nYGEUsUcFL8bZRhQuSaDCa283gLzcWG
YGSg6cMfyXNgiKloc/NW6B+rexRguOFZcYw73BT6HKHNjQjJpUPXolJGxwakMWBs
hXeFqueTC7zc2UhV7oaf3C2ZxQ1A+y1PcZV/U4xEwI+psfhq+YY52k48ADaDKOJH
9PzieCXj41QlrWGvDPGY0twEWeYxD9C9rIn4YmmnpuTvBMNFycomwQRGJ3ef+00e
LF2+hdfevJ7MpqOnVwx4tJN6y7RRak2N4GGbesZgmGRNGIEwh2RdfxSunHb43OnK
stg0VM8obdA2VWT2dKi+RnHje3PdHcalBCkP+EgTv/NcfrYAIszGw3SRjHFjtOHV
ILe7dMwznm6yHyFjFMfEb+ANbNuMo9tTatQ1x1/Qy0Vl5QAYQPGmUlPti/kxytry
wpaRUdJmEJBldwwl9DXhQgqR+vKXqLakGvmuWlBiQWF66gSYgS0i3Yc7OlDwIvEe
Vf4fIHKhRxjLp/nIMFOGw1Gh7tPAO6+96aoge6azRQ6z35LjUabl5PWNGmv/HZVD
GpwpdRHIYHi5sMk/e0bfa63M+cqsSeZrlTQPuBkmHR8r+1X5WHMDB4iTcbGxU5IJ
W3s1KN6CRbp1cmQScP/ClDMw3PjBCUH9RpoXsBPbZGyNmb7MjVBISd3pjjX99csu
RCQpt9tcpQCtZ8E4S8WY9dcFm5IhkELH9Ciio+0TwWftsQz1Pk5uGcuvfNdgkgd0
oIdXjoKSE8ARlXe6FTEYWh7v5Jm3eQELwgtVuu8Rc21mG+EGFl+CxcglTYlT3Y6c
v7vdx6eqntkFNZCqIxleKJHRJ91sio+VGWwJHxfE6QvF40UeKCA9kSxbNosXei7l
feLkXgmWL8V+ZJM6PXssqU2DgRj4FJMg97awH+sNaQ0LwxVZioF48jzTE+tQ8uJr
XWON3z12B8+vSnqao2uoTB0d6E5mr7j/eg20ZIQWx3a7CzWARpvWT39Y/C2i3oew
KJFwjdewjG6ghFZlegn1hStulzVLaFgBpbFwxVZ05J497U4QyhbJ8difultA43qa
leAQNn/BpylCVa1EivOp6KWlFKlf46lERzRprI64RmKM5SqqJzGGtPgmgoC+pkRU
EpoOeHhQwqCgDArdfpUkommwrcUc+O4K6C66EOTnNsMBxsN26B55f+RzyT7Sfue5
`protect END_PROTECTED
