`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XwgMzF3ZeNkzezBMobTJj63z5RV+Wx5eZF0dFHMN1TG6v2N/+UZmbfiSh9V8Eq3Q
ocsOKAp/YS1oLP5LiqkaVb5J/Q0Ax6RUn2dsoBTbtbyXnkHIE2MzCJHCthmwuM4n
xB/mme4SxNh6opeNleaVywDdojADTMwZ9e8BXwk17K18HySrXCQ3FAVa6CipWws1
BoCrana35R7fs+BuS4IPTMGutfO61NoGdCauzVsPBvs2OaI5dSKGiJ3+UQEC1X6c
O1fXPfefKaCZiuWFgukDPAZqCcduG1/KqieDAOke6rKTMQYK0toSSVvavLWolE2L
7WNfgrk0wQ3rVf53GQfohSbTN3USAZaPWV+0aSuTtcdd78LsAQUt31PjdYppBOcr
27TfenuW2j1u2Dri6TWETvkMLmJcLeR9xY0sj/XaABuTusG5U1tFWIZ7sVtDAdJF
0PVQfSEn6ftNtPQiX4uDOCLY4XOiH4xBzPfT3O81ajQZMPZb8+obi2hnRTgmSf/M
0IBMehNAQFA+peyivDf9Bj5lU3ZMMtuuQxTJeLmOFT5e4sm7Weo8N0RsHSe4t9sJ
XkyLbdMzcGxDEZpw+Ybd8pvdfQSrVdqPdyrOD/92ruI=
`protect END_PROTECTED
