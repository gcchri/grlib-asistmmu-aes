`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hr8j090678Vo4aeeltO7Cn6Dut/PbsxVp42kI48D36AboYg5dUwCfL6+UJJ2i8TT
BUl2+QEGYC5JLppdQ6mqUZD4WwwVGsWqZfGmhuBzIbequQyQDLsNHyeToX+xNXiz
sR+C81UOX/2ITpCT2JXYOPZHyJOMopud59s77PpKgqelHUDZrEHPbs+2vbM4/NEF
m3NeWYBVymBN1IVIiTV/lfqtzp/V2yLgzNME0cUEsW3k4S4H0eJFS+aO1KBld9hk
QVXs4n+acqnqwEDtK28YnmvmJTfmITkJ2tCB80Gy2JX3QEuPaulwkJTrEMoRbIj0
bbb5NwjsFQ/RthjJ+hWZ8h7irACd8NXsCA0REflBGF4lOEwUjCPcjrMAlBbzm4br
IzSwQhjGZ7GZW5hRoWYt60FHqI7B5DAlnEZM/wKwe3mgmIxFW7eMkdgeOEljWH1W
/MelsoDXBdzejA76wXv06Xg1jkWQModaKMp4ZoLISY4UDxSidvabEAjNJp3acvHL
d2G5H6e/j/IaPg7UGqjGvURHfatUgt5R+mA+QeYGSkNonu2lU7eiNQD70HAGkT8X
Spxz4KjD8fk1TNGOeOGcm+lbrnUPTnAi4EO4hUIDRJpljqzNwS6zGwalTkwAyayl
z40DvFUaT8wBUQ1Rzwm5d0RG7fzGZi0sSf8i2U8lparR1fOKdBn4R0koMGz5Z2tB
qBryB2cfCoDKvGjKobZoaSbUEqFsXtbl0iIvBsU9Lsz6iulTkdynGVSeYedBRNqf
7nWbH7aI5VwcHcTFEt9HGewyLv5J0KA1v3zl2uGFuU/HrjnjZunxHfr63qjou/uL
D3ilrA9j7SYGOYcIAQSlrR1ZfIcsc7JVy7mYtKk8weF7nmX3AzuxLz2xdBuokDT4
3wvgMpcB1ypdh2jJfN/f46YaHMFKsXvq65C1Z+Uz3Tq/GrTV9hZD5KsD7Lh27TIB
MKXz3kSBxleixbzkPA+OymNqSfvn1q+vlwPqXi/YaDAGd3DwB0HuYAHqs97Hfegz
nA7gPDizpJKkLz3Ce0fH47N5w0nXR3e9GZyvSh4OGBr+tmBQ25+SmcvUK+J1gRrD
+mDGxUb1v7+481ADCQrRlLZaUKpzFiBL2lyob656RzvOu2xfgvGHY4iuEUpIm0xw
XWEtCJmCMrKAuBt25MTO0kKhwz2ienhJUlvOo/0rCgioP+AtYpcpid3YwtXuYTf3
uBO0TduIhT4nshsMz0zB8hvrOj70JJIJPPNWdIzHA+LAFFaBe700DeR4p+ec/c3R
tVGOYAbXGxPLDWgKaQj8IBhDj7SvGjhWpU4TEQJ5UlGKlJe9UzB0ZzYI+1XUJFRk
gDiTTNXcocU9Tq9aT34Ufly4Bev8z0OliBpkcuo20mNE4yYKyojo3zT7vnWY5rpN
zipCaDmtqXmhF1FG3jEwo+x1r1XIeqWfcbDxLXSBljepgoVeW1+WObWozOzpEwzt
uyP0CS2aHVH8+U73+8kCDiExiEMcIFtqValpl+zu27yFR0xMndbkvSBTPKCLm3MG
Kqhc1GgNFopVh0Jleff48PJZ744SqHNEoykqsHrwe32IylvhVnQqpkdmzpYjVNwo
TPzZXWoYSxGbym+ljsQbkoulY9rumcpUT083XM0ioFCeRoep9l4aAal4/rYgmjeh
tOgWOLQ6Lofz2Gd7OV7e8TN8znxaeHy5swn7oCimGhv/b1kSQnZ8kZKc5pBWgof1
Q94qSkZCMa17QLL2k7BaNe4tI5OOLoLkGMWOdWK8GHScblT95kSwmwRWacGWWkHD
NhfamO2rAQLC67bIohxvA48o+UY+3xoTcXqV/bW1jA1R4KdqOPsbL1QYXsygyvXK
UmjE13WQNWuN3ncUzfmZCuV1kkwORtyLZI9S4E/fn5ZfU09qGWIWGdnH7kXGJVMz
7HoANyLAr87dTg2hzciepYJlBkut7/oRDRhCVySSdalurOUdH5BQ/Rf/EdxJukGU
3zwvbCaVG7e3rlJlIMYxawvYcR0cKO03SXwrQcsxdiG8WhwqSMNlwiaC9celL4rF
JIRodK3F1z08vzQKTRZpORmILkAwLAdd2x2EPYn82+DHTBbujrUyDugocEbACjPB
fetERz+fAruYVC6s+Hz2FpEANUF+Bl0HPb9rBkWF5kBh2iEGrRVbn3lcKs5vPDYz
SnRKQpZEmVo2C5ftsEf21bnss8cb+INyi/J5Jdwx14OZ7oHiCu/Cyi8CaexWNNmM
Ve/ELD69MPWSf5GhOTzC7mzj1QTQmTSPzqgpYqU8DV1TLiu3xwS1ISb7OMmYkg+E
9UxeBRe+ItOCsrRugvcm1tXkgv+xk4Zl0xWCvOqhh6Emi9dhFOYK4Wz/uqlvcaiH
OqLtnSKuQT9OV3os2kgGz8l8Se1Pco+KicMVtNwMwTKXxF8OGNTilT4fZJ3CND01
KT0q2qlD6/iCH8rSLvioGWmQL69S87tYimem6J3XzKgL+GeqYXWBL3KwRVJvcz6D
+rvkARHoyUzH+GIA8hVPP9WZuP6bpmME3SpX82ap63a6h8/TbeG3cYb02Lk5vPPw
Utu8wruB8LqctcKSdYqcy1V/ju1pEMgA38IWm2qm9cWN+Mo3656LDWcLzrtarIs/
ueUriF8TGgKy3Di5vW5T3QeDL85D4kT6k0kjTOF4VgSrIjGOaRZ+WwNRyK7cTjWH
EoiVVt+K1THZk+lXwiq/8nZ5lQyy+abizSCN7qdfYE9IVEx7Ggah0fRVhpJcO723
7tSJjUGFgsyhlotKfuIrCL4Pnjx6Xf99yrz0+ith0q6utYsz3dt/bnuVIgQNNBGS
3gbNkEtDlYBOg/D0bmaDEpHpK7f9Nnfxls4l+8A1TrEQq8dEsUPRwM3NTBAon5WT
9ljs3ZXXdu6q9edm4BOQsL8hTbiQiLv1CLMd8uJayPtviGEBPZymSTfCiP89wXdF
`protect END_PROTECTED
