`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8sNSdO8XsK+tUBPVWbK6XyhGt8wmTcviUjd7ped44l0FmdqBJ6yb8LNzhPneef2R
N5rFS3gff5baTjI8jP962NolWGG03QDyscBna/HflOLr4Aveml9L+DEgt9sNzFc4
lCN8DhrKhhfOoolP+oFiNWzsL4ArTF8jE8KNQwdLgg+AOCXIFh+QzJhlXGXz07q3
Qg3JUjbaAf99TOJgNnra+p33kx7oWzGt5L0xIDOtNB9+wf7ygkYlKI0EzgWvoCro
8VqgD66/NT5kCnzlxk8lif8kX/pnhSkiD6LqL6Uc12aZ5Com3pVu9aypuwYODsyG
s3AnubGv63mPgO0zSwts06t1UfEx0/nbSWivKKspg3nrDKL6ftBVc863mYD/rAQJ
z3V4D6h6kNNoQe7nP8JZPmH/ACLPzbU4akIlrvtJFgv/9J0as8FXQwk/SQF+wUGH
R8W/HZAYu+CFrQzUJLpINeh+2vIGG+9PDjm4f6w+j+8=
`protect END_PROTECTED
