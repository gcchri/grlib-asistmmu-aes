`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WwbVLH+OjJbEMlEr3Pai/o4wahIvBj6WYj8FhETVKMhlsoLFQoI2k8B7krZ7aSP9
ccoOW3LY1nuqLUFI6bUZs2gGPKgqIRlR+ElClc1SLmF8PF6ltLzgFQvePVzmC1hI
TP3D5hk1RHPiQzIv5eDnQ7dRAZZIDw/3l3PhoUvUXNKJE3CuFUKPnIlKlkSBsXHI
yzvUV200xlP+uXN0v0iHtGNqiMiwkk+Wc2q4n4ncBHvICeOOI+tp1SgR3wjBdVMT
ONpjngty4NIvR2gcsWTewYJSBSW9C/Aje3fiL9UqEKB0xfZIDZRLKCbO0rLjPVnR
YRPpfk44q1TofQOwgpZ/Zyl90+mYye4PRmG+301eG+c=
`protect END_PROTECTED
