`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mzSHKpGP+fJicZB4oe5ZeP/XcdudjmtrPavWXvWl3J9pt7EJrWXzv9qSStx3Ykel
u6vs2CrHVHCUZXMeIfEyU2HZm30mfxobKRNChmct7j9Mb/bfNBb92GMKfttAxMl4
GIeTGVzv+8ooo42HiDYRymLkagxXrJY9TGsw5jcCXNOPlMVonXIjriUxyrmwoFYj
u/O/OPfm+afFSeE+NL6sFri/N/IzaWk798kkPlvkx8d03UgUQ/0f1y2lf91Al+Qa
+3RkKjQlCboki1jK/o0JKDqW8kqqV1TMaqhglQIHBs9T8RaBwOdax7T/Fdt5DOvD
ttOnGWJftZK468NysKiI+9CLrOduRgfuwf5sjGnDO0v3BHDJJbiJ7SWqSOagGixS
`protect END_PROTECTED
