`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+tbXWXQjWSgpiqn1IijSDLJz+X/cQ8zLr81LKMYP2Dz+hmlzbTkvL/7/Xv68boGI
5WnpMzmkJUzYIYcZkY/MKT58YFPjokvRF1c/4oSshaSj1EEsaHlurRkqqTbaQekV
1xQyLlGhkEpt3NE5OJaDz26QesRPlWXyP5iWQbmm0++3jypfdpOBFfvoztAwYxcl
VotdAI+Is893Jfbk9gHzqFrjdbsCPh8AT6gpJ5aaHNQtlGu4hT58w5mL5NlwpQJP
SweKgvBGcgxb9mDUxbvABWokWWyCPPzSgFeCWYmOHnQfyddsxAKQI+Xj7/30mUf0
6IzfIFO2FlpekBBGhUtIYLpTYH0Z37FWCxYu2Dj9UWbVKm40C7plUeEGMxVPZ+LG
+lC9nb9rhRt0aM/NmsKK28DWlPplcw6nNmjWcHV/GbI4Uxh0UFJ0hvMtk9PneNxW
U5A9znUXM+MQp/QBlvexOWXTclHaqVYSv9tYu7HU4VeWoN6x7vWdobqXotNTaW/Q
D4e6n0cRIstwt/CHfRRyVAEswcbaomAZ02SOq+9DhSi4U64V/M95BGp90nc6v4oW
C2ETMjo2vmkUZcuBQsMatA==
`protect END_PROTECTED
