`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
862WSXs/vsp+4Z+LZeXK4kar433VgUQNXj2BIbWmZkwzO6cin+OWE5jPxjAMLkoG
h8ePokUuFmdGRYjHx0gbblInliAGnn44oT3AgT0U1gEgYuMNUvlz4CtIzv8Mg6fm
/FqMiXzVN2GP8s2lB0Xc++o/OrETuHG2p7WKT1n3y/DfJxOOc5ycoJIgQCwKs5do
mrApEW1B2E8f0DF3c1Uv5XmRsQaz8Keuu4jErkWL9BfCXrpkQl9Pur4EEcp98zZn
qvbKn/c+gqF1uDFlK6GcdRbSWywJ4mJBhwIVPGk6tBoOF6wrdQiG5Rt2y0fYwHs/
Hq89l6KDnr2ruvmYz8xHhPxQ+hzFoM2XvT5RNzMaTXGofWWnkEQ/kD//WNfE/QLJ
bRf9eqdogscVpfJp5d+cjHDumu1S4pk2neI6IjwCgjb/U1jfFCyCgOAYnJ25QQjr
lQhUa9sfdjYo7PuND5ccV9xJvz1b5zsuEdtUO73/Xda4+2HbojaLP97VovXRe6Md
RL/X30xTh6NV3u5REOXNxF2EAGKr8Hy55wG4RFyE0E0TelCFymXbiwbhGC7vWdqf
pAafXoph4Eeh1m1U8HcpuxN1zJWV85frjAYIBUDV0qJ7i0W10350bMJo6+6xHezA
8ZgI8Km5ZrkyEu15jzKaaMtSVqfo7+zATBqHK8Lvji/m0k//0t8xNp0wSD5hJEPO
SdKLF4d3qzbRpbu4rg+Y2J3eusnO234FQ2r6B8qHExup5goJ71CbEgkdoBFyz7Bv
MfPh2YrHti7XZy3sTXwHoMfl7aqC3xNCGh/mNNQiSNWLXX447cJI9vdFlbsDrZdR
/Tfnmy1LT40AhuiN4iGHN+I+vnQ1nPlJ7WOUQ1JUi/sqoOKRdRtASFX619vL4dEx
PbR1NZl2Sc4x/k40r/j6KGrzZUe2SbijloKEL6GitHXHYIIu+4l/vvkA2GYQqSYc
/OZhpTxJ55ztmzH5T2epZ3ZBQxlf7+OIIwFni/rFzWHnpjQ0krg3t3QJ0jgIKpk5
BLvS2E98UtvGnpyKpzEjkx+JQ+FCcpUOpVn9cS0AIg6PvGxeNDbBPfK45NCI9wSu
wZERVdcYEjxhaRHC3lwDkFjVOGJo+9QrMC9wyY0KZu0y0qqoPTJGLD0qWy9ol/8d
mrFfEb4qdNarrIngDJEsBwWUvp+2M/MzeLmhEGQd7mBdZEX2ug4L7reALcbGGX8M
XN53Lz/0/aPwqksbru6DPmfuAPrmaQw9ZkblIkkHZBN6zgCvqmq7eFaTjNub3l1n
YnxnslqrcXXoh7NAPJcX2+q9Z035OaR83slxjyLcuZQ+TOeB2vfn82LvU4Co7AMl
6d5elntSY8Nus4nONV0uACtRLsDGS2TaQY9ZS9ldPHRee8mdw1yGHly84n8/ihBx
O2oHJSn5vfEHOD0m9FjDlFSnJVBmhMD+RENmZhnhTen5aN99HbENWVtYdZrzYPlb
zOr8YyadTrDdD1F8qUx5bwloNzbtcr1tNqqUjXRZY3Q+ZU0f5u+51Fv1fH5POToe
A98X7YQn/PwfdQ493KU/PYbO360MhBljJ3fhKWADDRM/KavAhQxUBljgrxU6bhK5
+1UQeJw1KbDCxHZ0930+k7rw8uXpVS2OVmDlUFrbIB/NN3NhJRwU6+ONWzQeFLvT
h75qpHc9c6rcuwkd2B1WnWcgDTVAO9ra2i/OFwyMY0ZZfV4tSHavNK348wh1RLp4
oPh+y3vNpBTQBvt+6a950Y0i+6a06jKA04sBW4LscOe3CHpqd3w8KyoF+F7Wf1iz
Z1VkaH2l8WNKGD17vnV5H5hw75ltf5KHQeRf8rB5k7WXUuqJsIGbxOCq4qcJrA/1
B3BwZkuWHSD1oh2eaMcxh3zN3AX1zLGQvxUF8P3KSzFHsx01NEuLu7BGDc2pRA9p
JZRtCRlYQUO1jUJcMvJr0Nvh1CwG9A3hl3VJB90ULcvwFRjvPgwhOpHsW58rvL5d
CLy9LTljsTR9iXmyARiS+50AmQHD3BttNAVDUiuRlsKiU8LE/3MbTiAUfvOGFP7M
zaBfj94dfgB52bjngb4r1SlR5hcItSy/mOM1iHTEkNPPusQSMwHvPST47aG/Ml0v
+OMBKItfiN+1iu+mEYJ7Pf6HhPZQLsQpNzosgM8SaT3D4wgZI9aL05Uh3bcl167i
/lsVLnYQ9kJuSC/o23KRiqowV8+2WUzJpZE7rnc6Wrh7GkW7Ow6w1cI4FkSnkTYC
Mi/0f7Os8/EWHvrTDyR+/3//ciLaRfLAv7UWWPv6mt14ME21xtzvWZ6xsAnXwqdz
ziDUclqjW3um+eXMxxqjzSSzoW/N1MX0ipdofb7npSxljQ/4Ys0OLWvYre8iMpcw
dWqcLaONCvhU3Vckwh5tJbT/eebO9RbnzjrVVkfBNjiIg6Uefw1ZQxKz5lX4TNg/
O3BgKmFr+h9zPg4/oZG7szIPCSwS/rbAemQa0LF0wVqyXcIgzyYLNpP5EPEDgy/i
/dKbZIQYR0+mKNSgrbemJw==
`protect END_PROTECTED
