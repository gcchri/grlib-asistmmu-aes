`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y4229Kq/rVCn92OoSGmVC8k00zLhH/9c6oxFLcAUMmfhL7m40+oalCjySEo2a1Ln
jigStd33Z/G1d2xZchXX+rn2Ngc/qsZT2ASt5EUAPUlrTCJvL3+5Xe+2n7dfTr90
w1w3XsOlMIt8NzglrICs/ayMrYpSIPzU4cJYRZIYbst2kr6cRRahmCZPATiz24my
9UnovC2nw1uVfRcshr3i9iBJD/yz2J6YRvO+wGtOdGuu/QuQ3qt3iRMZ0x3CKpTV
RuLqsTeX/drqIeCeJU8cXqNVs5np9dDg1N1my2VJdNVjtsFVp0Prgw7Bx3RRYwhs
NdEPamKmwns9chXgzXHQnYlSHCIWitpMFEhzTkiJNosf3eHXOF91iv0Xmx69Tlwg
bd+blinJzlbTW4NjEWTHRGgYp0NFDkFlVty0B+8yHVYeKM9LDTPRF/SCTU8CQg7j
`protect END_PROTECTED
