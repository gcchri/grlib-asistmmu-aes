`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nACI1fTankNEY9+tct9qdcGJ1C+HKzTGeSKCumynPqEn3wyECXfD73rLRlhRyyiU
hHqfyKBKtYn1ySiQufb9S9tUQtgtQ2Kc/XZRBY6fKp4zPB7NNzhbLl2xFcZqcJSJ
gk9Xx6PsHYcd/6P05hjICDhX3FL3EqSi6a2SbLaVtMT8ggVvnaFw0a/YYHzUGO9X
ELCZ25yv83KsU5o0RUan39IEkSAKmMB1Gp2GW11ukotM1LMpBBDHQkxGJtsL14kF
ZG2NK9Ve1mHvTHiozvodHYam4LIyo7MlWE70f1CxpamF+25gXNG+TBdAAgJLnDQP
bytbsbBBkoADHaa1tV+H7WUY+3Kk9uhHelngF0zPqFsCbpYrL1dAgTkdTTMovJp+
nLQMAKiMA/XrIcw9aRNZFQ==
`protect END_PROTECTED
