`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6j22HigUzSLDUFFNLbnZeOM99IQr9qzVgTEmj9K5vl6+6s44g2wuGmy8pJUrVkc2
qC3QBVBd49VTIs0Xppi9tlaDZd6Hufx/gK6c+twijKFVt9hTZ4mpzBXNsKrfqQ2L
xJoPdhKw+g1y8ag4qKbgK078Tqn44S21SmDt17fDHaeAuv/IQBrXI4FFuuiap555
muKMuYcs5gw14uQXLAsi5AtUo+vLIN53bWvHOAVgrtg5h4G/3FFiIE3/94/azpFc
MrTLrBlq2mogMXHsJqzoaXy2/cUl2zcsMbBs9gC5NfAAGSgzSYbyyD3oSFiOeZRK
EI/YY477fZTP/wYClu0gzaOoUxsaHmKA7DgpjiYIq9LRzawBOG+N0vZIpsFsp6Me
sCND3jSjlCu5+pJbaoFX0NWFGJB3mmAYSu+NwAVAc71Au3D5zrGfW8dcVlMGWu1a
dlmWLSI0fKqpo88bL9VrgWYpKGLJIfuxyRu3mCqfLaftdWo2ObuAlJiCVvjcd2VM
PPosrVOKwm2TeapouR1ZPtP8e1GeI+Qm6hlfzb5O/gv74lCPYYHLsyBOZEzNUpgo
vE+TXa+UkMx8fQHrxDNL/25rv6zNbujNW3GTuaY0WX7f4yQEndeXflzD/PZWwoAX
0fxF+JqRX9egTG2l/g7ggxOkdwTILvHGtfcXyLmq36TplKi9eHblHWPGSUQqkzO7
+av2iXGyW0ijVaSo6CchsyZrG99GCTZRguVzJ9oLLPLzVs6wxlTVltZL6gWaWNJX
PqkvexGxVE4dP6ALGCPlQXuwwpy/qfhfux7LYEVwO1gDTirc+HD1tXXo6CGdmIN7
`protect END_PROTECTED
