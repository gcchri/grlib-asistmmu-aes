`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pmxp8cf3GMZ/bVNirPToXfTjCM9/4Mk9JJTP1KAsf+mHmj0lmSwzU9OejY1Mac0L
E4Oa8lPBm+zeFJEE/FWL+qEr+uCvvWeXa1pcgon7nnEPGu8oNEdz+vUp7qKq3Rz1
1e6Kyx9cJptqKNfMFOt2FPI0p7shFbxmwBpftXthzVDrSiUu6V/vCyQeSIZiEJKP
Q5ZFIsOGYysQBlUctgFIEArshNgqM8Y4/Vvq7yYbccbYDZMXk1QFuG9WruOpFEyW
0PH3/Lg2rXO4LRPBZmaiZd5BFtK6LjY73Nsbb1/6Ob4ZeDnVa721feBteGjsDZqN
AdrQZP1vlNrkUi3LnlDXu/P9175UBsE4SdiZqGtw2L6BDMiPdrZKKDCZK7wfcNth
GCsOhQeazkNTq4zbfNX0rDq5y6/WGH92mc4AOqOGfVXFnL40YYpf0+wGmOmtzah9
JW8V4iOmxDmC8yKYpJ0aCQ==
`protect END_PROTECTED
