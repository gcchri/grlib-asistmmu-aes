`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yKzVTu0lomu6SzqpSwgxLs5zRwhUIhAGo7rpev6gHquoVu5C/vlNTzU3mGJRcwle
FZzvaFvmsyurFAMeWong6cVjLJYz+qrLkplRqEioyKdWbBc0oOHrVAOpqJfFsQ7r
xAv9FJgNPqnnFx1w+sk5Key980bgl9oF9JoKhsaiBVTFqjXtrK33tTLm9rYkbZXp
U/V2LG441zvuD8pvLd5CYt5xvC5685Am7WDy9M+L3qRNehhRbWy0wTXfMeyE4xfW
qnnl1dLn2/8MoBwNdMtmGRIuM9f/s+EFkPzGPi5or0hTFJX+2XEu4dSiP39NmW/T
5HUCsbYTiIVAkY0MQQfFxmB8YvZgodMUtEQ8cG/SYiVhXT/2zcM+37auWkqFzyWX
/QkRbSfaRwwvGw0s+ROBcOyMfBdwAxYaWxY4FQ01WJBz444vRy6vlGmS0b9VrYZP
uMAqBLpMzWh8IhEvm8u7t23w0er3J+sVjAaZ4pRthjDjXbvepzR9F4q2l6RwbR3y
fwZEuZW34uCHAzFG5gAAnsXflsDi8F3gqcRGdYUycYA9XvU5pefLYXXziEeo/Qyv
yDFur2vWyeTfic9AA9dQ70YwebQ0qUBk2Q3I/amwwu42qfcTXBW1cY5DZAEfKQus
XaXdIMcKM/8ybxrH0IwH6I4ThuOAjbb4jX4yj5yDOSBCfVV3pcbmBCQE41QVWcX7
geyJrMbgdOvSfD/maCCQkDrlyMn9VuLW67E+yeqMZxSXzTvYNCZQUSx8F8vbBxcG
E1yWA+ayOEugwupJlqRg9Q==
`protect END_PROTECTED
