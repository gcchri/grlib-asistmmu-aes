`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uDY0DZjncf5ee3xNc6j2Owwq0kZY8FAubRMMH5rE+aoU7HhB/+CeN5EVcX2eztNz
Rg4WW5Z0BhQID+ToqORMeqY0l005NeXWkDZH+BoeBWpV1aRkJC8tqikpvNUDjE9q
0q+bqhUiIXtxwGrYXNI0j9BI0UIzEiut/yR3lsBu//1nWDs9s9BG5iFXAEjH1Hx6
GU5AfLlvChoA2T+k1r8Pl9ovgYyVHd2wsh5nl+Mlf+FEHWG7JiUNCNQucmcq9+33
Ls7WjJH+4hD05iU8phqDZZ5cNKyo/b6/ySw4fMGWExfNmGpp8wErtnP7dkYC08Ik
t0f40TZq+o8iy8gsAI2gg19qQ2Ih2eB8V1uFYbzuxZGf6bDKReTYPrnSPzX0nTHV
x9nt/TequQxMJDbeV56z8oPjuv/qW4LUEl1b7yXYZkfVHq+zOOBXZruoUITdXB2x
ZqKP6U3r23J1RBT6NnhNDuXijtiDAC4Q0MPl9MnKBdRl8Av915VWR+5BuAoM0gls
c4xlUkrRxqQsVdyx4864RAhUz0BcDzMi30nVUDymNF8DgYgJmZpVpil7LaeM5lBC
yRCsETYNterIR3paP7XHYtlYY7Yhn2dbIAZfu/zucSOasLRDAq/0VXqMhNwIR6wv
hlHxisvNABWvN3RQK10AkbKPxyoz5lzh4aDan7JAUI/o6w+qRN7QIo8kc+fzbQ81
PnnLqgFUzQY069yKcn30Wzt16zSZsVLxTQmH1sI9Oe+HBf2+dLuILr7z91Xr6X/1
p1oIbNrZmI1zmPwl9jC6HzalLpljvJND/4JvcxwqdlW4dCwzVNolx0WtoCUVf+9C
d9/hwB5PtAIigpXm0BZG+AGn1WD3YUQDFK2r4VJhGgw17AhD2C6szdvcoBsGWpqC
IeZzuH8NVXToun5CpV7k5ODXd35ucZM5jCq/2WzMXzc0t9bNlnx3wvRBraADXJty
DGA07o4JBVCZujqtkJ3QUgfJhtkksebzMiQVQe2fiUqwHxNPUkuNe7vatmEvVTgC
9jKJlMrdiLa9RU48aiSNgVMQvC1cH+/DlHYs+cWHfguiIZVJA8xOIS5oijDHRH6r
NQFxiplJ4OyOtz4FIci/8B6rtJtBozL5p6FbD1i8EZo7K9w3/BTItraEMEbYlMHC
yePUw8bPAPruyc2xAXvERIK00ZZ9pcZiF7A8/oqUuhcSOvmQxoYsDNpLfKKQ5lvD
vAGmmftHdNYU/CZUtjfbWdCeeVJFmQ6FX3oqBa9uITT9IA2uRsJovXw05E//MjbP
qKFxl7Vw3WndLnxlQp/MMsyLESQFeM/VC0xOIJa72N8RM6unwcsnQWiAnGP1eMiB
Dd5wqt+/Eytf5GQQNOEt7J1BKrRse6vuWbyeuOhXP5WeTY29PqBI/Y7IH7UTwa+O
FAKsy+ely7xNdMSEzNhlvcUoKXxt1e8PeN4QsgU6yJWp+Bodyl5IuGC+FkDJnTw0
9k2D+1BfHaC8v3bEWZyxVUlY/cJ/GQvStRyhOFT1botPF+qXS33tiXzC5b2lNxN9
wb8KuUJMJlumSj19QbfW+qb8vu8yFGZi2pLv0TxJdbjLwnI2k/qzrzNvVeWgH+ne
LlMQaw14h+JpN+coqaZazJ7LdRZuYza2kaoL14RLtcTTqTOdHVlMntr04PRhzGLA
u7sgZqKYEt0RXHRyHiMO77hj6heaES+WApOZR1EjvgJYoTUR5m/ySQoJrUr5+LmN
OvLdCz0vu29/hAXBIGhuELJxfW072NUt546QKzFp4RAY79Ta/EQeRQG7QNs6cvg8
AacK+5nbzmR4rtxnHo73heMJ2VrL7n8nbNighNAimAaMVE0SLklAZdzcwyCcPRzO
vqrabLMrEab1hq85fpZOx4LIVQF/W37XBbfQLSpI36OmZn7UOfkcFXwZfzMVEdq6
RD9zShBYtonjz6QUjot/agirR56zVRqscl9WCNZDhCC0+A2I8AGbaIEGYFIktf8/
fSSJxmrUK5ZKUYCzcG97gHPxODKrVRewmV68oJSbm3k6fcei3DkS5XWouc+YK4/n
kiFJHtNOC051l4pzNtHCGajcXiSGUhtZ0oeNdI+U0QtFlg9QyZmZm+0/1gZWlLEW
HjXxsrDgsgR6uv0d9tkfKROTNXjQI71pl1u7i2iR5dpj3i0TQZituiJAAKd714jk
T4p7aJ7+ELy2kc0YVkh/is0oUqulB9rHKGkUDmMWslDfBKA30YsCAHQGrL8E8Ror
xYTF5AFB95GE2ChlZxJiCD/k+Z/R6Tpx7QnkKf3ZIxYd8ORdyYUYsmm2NFTi+TiW
EJMbLQ15hzMYvAEimJ53gYApHHh19Dz7aSXKRvpKEHMrojXMW7GPjOfZvJgYI4Gq
RkmphBdvRaytA9T6L6k26lYzW+bDft60oQUEgEOkac8YLkRsmGrBqHXMNRF9f5fF
8K96CFk7qE/u/Zy4LVfpr5HREt50E/cAj7ppeJ2BjwVZuLbpwDCFUpsIj7zRHiQs
n3jq7Nv9mg/O3FTzS2J66UBTjMD5OUs5ywUIbh4tgJmB2FKD5mtPY9bj79WCRFKG
wR5deJXywdR5heIW1inpPq+RwVrM14Qo2tZ27aQ6ITQFCwsegLf8f51U91x56pz5
A8JSV/7gynRXBHbN6snUhDPsHdM3UmhKMQM46xdJLYThhwUNDA9b0cLsfmUaBtVz
EXTG7/nPfCbeTXddyeUUn1eLjxLf2xW5JzssF0uq7+BZxbmYrz4IyJugKuDa0pKp
ci2K0XZm/4fpWotigKRRPP7OwRbKq5bR7wn+NUzFwI2oDeD4nOSHSnLiRsxCz+sb
NiymLEPctWwyVMnNFJ1OEd4gGa0P+mURpVfvFj95Hy13ZAioEbl6eCXgrx+4K4WK
X0a4z95QoJOU1CSoR3h46OaIgXba5c078cAyI+PBfVMzQn/43UqIe4nfFuBxrP6g
82o9Y+UwSg6MD49omi6r9fu9vxEMVFYjm9rIKnAKdZhM9nSuDe4KWyhf4hEi8w40
d9FRAaPsDnRQllrRCKRyJtu0cdYOk+Y0ZramhmPHzVPef74LGmmcKWUjMMQ9yjmv
oYhGYQo1Js9z/QngRIX+GHlSH9BB1WrA70W+cj372XtA88oEY3MIew5FnJk2J1Uc
D+9SwWoSNg7+IKSJ+i9cu28YLqlhxHfTkmqHqZQwU4MuIWf8OWYZT465QG8OVrCZ
ALeRREvqJsRTpCbhfbCGgQOQZEsyu5yeYBhuAcMeDuiRR/aouCIQnHJ/tJDoWjGU
zCMGU4LUh2ujIRgyaWaQwNBH40/ogglO8zZfLNAb2Ul54hGblbZ1omYjJ1BVW7Ut
6s6GWOjtAEmImy1DlRJXd5rUSJ8aN36jmWDGmKVIH9IH8n77AaAUHFZlZXs5aMU+
yiYOAbFegrlmz6Eq3J1ct84AuNToLlU5E/jhJQh2Z3DNV8G7zdryegij6Gz0IkcI
30M4gom2d1fa9JAJyZ3boWTIUr3I4loPGOWmGm3Ows5DWCbG1RUjpu9O/tmDAmLV
tec+vZIeWxhZrA6VpKBYKPpM+N5xGhKbzDHioxH1xtyARQ2RQJggfnCDEPoHV41Z
IuzESaftYGKXoQrQw8mD/uTsX7bKSJa/1KhRuLDwZwzxBw1eggcYo2z5CPO8tQok
rCMwDk68vBrOqjoC7MyALPIKtnEScjORhm+y3fOpz0lb62dIIuVcP9PjqAQrJtHB
sDKt37MMA5uwYMU4mDKVcwxokOGszyMTcxRQMstyJ0mZkPzgqyNbaH2EnpvIKNOZ
TScI3Oa2v3rtizqSZB/vnjrd0/SYq6XdLXfovgm7B07ywWJL/JkLtBosewq99Wqh
qROkYs2u4lSlwqaxvcGyhKbK4x7s0VIGzpz5rmxYudtZd0uBS8H2SbfKJZERP6/5
e+FhBeIZgWSWSCplArwSMygzwd6PRN8XAcvAyM0M7T3ahUtMdbTdOWiEkWwJTPkh
9g3GzOrsp+IacSTxc3KTbSuZeQRFZNse/IxjL6rCIQKh7M3oNi87OR53YDeLha4z
PsKMPsLQSE5ibu5w5QAlkO+dKXsvgBGAzOZdluk268I0qIbdxnxbN9yUoOeLcjeW
2wjoBxB4SycRFvkrIvrsznfPmwPwX6xskwOXRouHvMG5gomUQF2WONPmX6FZG+Zm
SQcIYCenZ2GCcOJYR25SvXVbMn3ScbjRwbPa8Ag944gbhMMPQ6fNejHz1EDnle5J
PnZiufB1Y5m3Ehy8rtmPZ8K+hh+MdLIJODN2h9ddfQrlf0RVGEK+V4kMdd0BfqqT
m7jitbc3y4wooD99SS5sMWZEMxxxsTTV57vqGqO8Uv6cMW3SbOyM2bOe2GIuHxvu
wEMjGh6Pmfvlra8/Kgo0nsQs4YUZVy7BuRbQUAQ2oYDCpFLt0C4vfD15MZys26QS
SmbNMPH5xaQazkp1zovIPjLpfgpaiK7qcmYo/h/29Rdc3vhFW1hN7QWCoqhbOQgP
vJPft/hGRJ67xgKe55MJnNh08wC6qIj0RIS+TAa+notVTvPZOqhmrexXeQI98opf
fVYqaJAFaAcV3HWg+Kq9aKJu+keU3FhdgERCDvjX/7peHXnSgudTpSmzWyRq4ZJh
POXMa5gDnrtvmS9lQMeUaqnGOrwhJwtJCXVvNekKf+jf/eC24iWKnEcm1PXyQ0Ym
dcB1iMzjcltpQ587BmZub9GKS0HHNRoJ4Pqg3zTdFqihOFmNW+WixRCGsyFVocpY
dk9t8yGQ+ELfurrE0ErK277cLFlWVCYa0SdWTnRR0sXuASR6JHu2Wm8hZvRpe77B
4h+46uNOyf1eq+OqUaMsuHqgmAKVFD/7oFHOcTb2OmDgvhXrgUTYDnGb64DPp/vt
JPEr7AmEdvUs5yX/Ory/pX1dbMM7YotFN6ex394azxOvpgwMkMxeOXb9kU8t/y/m
ayWesbGEICGX8bxRbmnsqFNHJ0enyLIC19+RMVeqzKjgHKlfowC2vCKi3iiWdiE3
aA3b+KGknAfqFTp+2FhKG2boJ5LephV18FEc4KhaeGWDCeOlbGOfhwTnbw23GTNv
xVEBkElxGE08zqiVLPBe5iXdKzTH6lvUjdk4cVuF6xxWnttlOLyUj/h7iYL9xW0L
zmlnG2fFGwsoxvpmOIYI85JU0XsCEh8BGTOCK1uo9lJ8Nf5+j0f7wBvYQNfSut6O
I7zHuwXQOHxEMspTQetHZQHZbzrJLjmHOIQnGLWCdjQrqQKrMYQG/h9J7d+PoX6x
O/6xaJKTsg2ObOMaxC7BTH2OWM/oqniKsmd5PnQiLYlecQuL/CLmgxN7Q2DFmo7P
0yKMHcQV7Lm5FGcitcU0BztNBpv19iB6R4VycVNphJtW9S5FSAyJ4TuW+qDPZqzp
zzF3DjW6N8Mztj8uMOOh6cAyMdTqRYfaVTQJbr+0D3N96fw6ujPFGAghDRgawNU9
QL0vUmiAAeD2X5w+cPSTMdC3PYqfDiVz+R07SNDAZYoNl1fJfO+Ym/9X9hraxn4x
d8KQoq2prLe6q/+Rn+fjFaug40PlMYIO+WF/JYsddoQuX1OFpmBztcXcRIVxcap1
gN0yNenghkbbQZK6+4g+bhyJ82IOSj5ZIXADVnjBA1KAyOJpzj7C1m1olte4kewx
4rqjnNQH3XzyqLghvXYfaLSR8WEyiwcUqnw3gInZKV51EqF6S3f+kbL72QCb2BAS
h5rYiNlYgZm1TCU2R1ii6WclX9z8hRvyg/0XZk5wqSHmKetNw312LbSm5GeucvYN
qKunbx2P3uab58JUdx9F9U81HRO2PdxnZKHCgzwmHXfrJURJb3692t4WB0qjqi2V
aIoM9JuWpXriYknpGXTqCS35IaO0zCGQdQgaa+6Nwg7+3zwkU2RtuT/5ISf3p+M5
x8vl4tAnF18vHEkSq21AgEU98zLCONSgK6Wj6QFu5y2VlrsZxlgBKSVaLikL9EMA
`protect END_PROTECTED
