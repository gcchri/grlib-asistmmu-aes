`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dUxlIHEZHm77eiTjJQADRV9h0v/kh8EOxvWMQxDkFuvNFa0CphIDUttAOGaI/i+U
XU4Wi1VCUzRmWt3TSz72jE10YpoSSE9P9b1qW/hjDVhtGG8+bLEOUQpHwiBqiZbo
875rYOsh57MOlk4vF3JDuHLTC1o1nSoGpmq87v1XVt/fPSi1O2PnYqYTgA0Sdlq+
rePLDZv5NFeRR5nQyIrVg5ihtVrM9zCiX22b102N5s2yGW0VJ7EHm6RJLh99cQJG
ZwNe0xHqboYsofbTL/uz2ehhyDQa0bJCabRORVQpolgiKZ1e6saNdtmTR2OaJFr+
`protect END_PROTECTED
