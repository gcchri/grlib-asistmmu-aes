`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gi7u4H2E6SMyx6d+BM2GYX2VjXk/ktlCqKzbNTUC2ox4jGYNIa1ayCmmlL8wGerA
BSaAPy0zGQsveJ4wlZjDBcniT+2JE2ItPCl9AadpWe8uGwpWrxCd6S58kbd65gnM
dEY0/gm0cYsQOeWck0hgx61V61SBN2tpEWU8RxOZUvu/+NGppVEJHtJp9T0P/vX/
WRtd5KS72F9xLoqnsp8Np4pMiNoNyjmuiBRNsNa33K/sszABhM9pRFLCQSIm1d3d
NfSYNh8DyT+3onlSmtFHef9L+P43DS08/OMkngLc/ZHaPGkpIr76IhbnAJKtake7
TmnIuw6yETg6PDGNjTHDJneFj+BdpvXP4KnOcCPFQswUsY2rrvQFM3LysDCUOidr
Kym/6TMz1GCKhNmKlBdnjBu+dyllHvfFC3p2GrLdwpq0yyyLlhT+NpNKCgDEsYIA
`protect END_PROTECTED
