`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a9qclaBHu1QxJHKnNM4obyIk73/a7/2MtTHfdtTU3hLN5nSdYJgyklGo5Y9PlJfW
MGfX/aQ/rV1m95OnYSI/jSsdiAUrruznOxLvyuiM/GsvlTKV6/u+ezV6SkLDVaDB
Ye+lH0g1QRRrV8arzmAxczC+5wo6xde75UANZu+CfBtyFOMiFqsTi3ogtgOWHYtU
7UbKqJMPpw8iTRSRw3xypy9XVJ6sL9NNpAnhnTqP/ParW66sg6oYzs8ITxnD/NaW
psm0u59vwVpYAKisuLCe8JdR+/KKt6eGeT8rU67uDvaqSXDvOiDeioHdTmCbnwNG
qCO4WrJJ7Los/BU/9mvh2I20qXzyYoVPeiR+eBa8LvNbkFP5Vuuen36lXDas7Ic7
lpKMR+3P+076mjumlLWylczQMOGChL3WIU9yNN4RTcOZNoWEmBg0OebSigUwiqNM
cxX9P15d8EamhEIc3FGEmnzy72w9ri6DI/bwLopc5BYvnssbpxHkfNBS0EeezH0b
SrxqEssMt8tiqkZG5nRraRbm3+iVXyCgjQCTtj5R8rXNjO8iBAFwHp1s62MRH656
V8O6PcWsWBDxj9QkMmrJi0/r27M3FKo/E5xosUeEChye0ESpwzFN6Rdf4nVCi+wW
EM4cm/Q7GZJDWLxhqPq80xQvxCh/RjuOK7msFLLjH5DMALyEOMgF3f3fQpxZ80vK
B53voOPL4TSP47w+ZEUxeWL9sLinQ1fdlHD9BwzzKLeosc1n2yDXqXkyOsj1kU4y
IFijV2yTchA7CZzRoLvc0ZCOBZpcRU/VtCJILzh0FYlABeXYrTo1d3aZMrELQRxg
F5jMYTMYn/5D+TmMfdgDPRNizZJhGNoPK7YB/dwrusI8QYlcSugFKcuBUo5he+Ye
YJEf/NavyOUDCcJ+yok8KUkSPfCwz5iiL+LXhv1f2hgWzDPd8O6J/rW0C8IyoLhj
Tjcox+AzLUP/bl1nm0gmDehzW7mjrCVlXKAhpU5kk/Kg4D6GpYW+hfD2OTLfwzxA
6MdBAUOkR/MI4Yr6JCz/TsumdqQAuNdg8+l2afwW/JsZTmjgqulLAG28YvFwBlqZ
OaZPG029Sb8l45uIBhe0fNtboSofRncHSRby9GEkOTNcxt+pgjv5ARnvLeFeSfi+
JSrCSuJ5zR7KVp+s++goS0iXgLmgENv3HO5/nBe6je+vLzghTmliw/Znc4MDFqiv
vVLP6qeM8ql9Oowj7d/XpO+iyhpiDN1544Fq9DRUjIDfCotHMTuFZixrTgToHsm2
WD9YOg44B6I8c4aZCBBK+9emLzF8i/wQf0LRU/vjTFIcpemtsCm8vuCX1VTmUqq/
pJ0r314uTHh4dUAM1eaw/Hf17n0ujW3esbi7axvwoX7HmXOG3mVCwzmepo0mu+Ts
BhoGxD7wGk9vxBDBl3KQvBJ8PEaF4t0TKQQj8A+UYXhru5bdHz3eX3Hmj3U5cMAp
+y4pnhIef96AcGmJZI1ZD8TJSzGcXrPrsCiED/hbIMyVM1w8NfLFG+UQMyC8rNuh
XHwxV71eiCsrAvnjkx8VJ1WED6DkmhaDneLuJbNnbUBNp2EdsXjinoW5jZlUO1CU
9br44VGMQJmwJMvr7rV/rpeF1DstYWXd670NIHmsj8hpS4usIJW5iFxvNhW+ZwX2
AXDU4b3AokYKo00mLXAB1YMrIUstkHmQ5aLHw+Mxu3m3bC7TqKhWRDxbPAYQ+duV
d2264dmn4vqg7dkaiS5k9UmfWUf9F08iM8L6XfzdSDPDqJt0zUQsKfgUfPe7zRNy
1KrO45uKq9Bbkzeh7nZDBr69IJLVIDdJg4n16l2kCk4zDPCT+mX8Cy5o099sAFVO
xoSC+fbqUFNMOVyKH+9d3gobHtmPXPmq2o9vYfn51xZHdIwOXnoI3FjeTQ3OJwt/
OSdPgbZiBrNhtfXs4VUUZACGZ+/GITmy0RahQw2bLrzYkxeD+8j8tuaSCgKhi14K
qms9v5mbUzlT6knH5QWC848hoFbSGM28tZFve0L7ZkrhHvlMt8qUQIlpG2xraPdQ
dvd8ZvZxi6rSNxuKs5c+L6eDmIVQ0WiYjcDjUYoNQ6MJ1Q6adTh2Uzk7Gbh+MH1N
RY3GDHjnySXaaEUDhf6w5ojJuTGdFBePPxR9QQX/rUNiiMNxRQ1wjhdmNKXC7bAR
SpCilnY46qCUwS/6+irmtOT6czf6slSzvg7lSoHxMjQhwABN4Vr1nZFcm+BDgogk
xwmyVcXWyOHi6qqdOx/jhkXFC5m6P7jeH1KpGekUbNCgVsgsHZlROLw0kI6aWkfg
BxNHHqBEOCxfXXP1dyAN8BFVOyUGSBLmzVKugUMGwzCkbJWtPdeyaPlWnz37ZBb3
dBc/W07z1SkOJuYknsay4R1bcqgZdAlxwenefQKqVHo0v4MduMUg7QcqxGHKtcnL
caJvnVcFnjUP8jHLhDySYfZxrwpyqx8uYpC+Fs7Uht3y0CCGI3xvPEcENVjDnfG0
e/6a9tOF+cI1fJ+qch6hIQlWqA+2x4pOaUE+E6NRLN+F2fTOzoPxIIV3d2jFXjn1
VNB4oQTQvXKBG6Xo6jv024lBe72Lb6Dpmsjswk84TD4478/zcm5lz+4XHB31+pve
oqaH48cPYXsjWWKOMGu8C5pKzxB4+SX1WS7PdxwBZjC6S4fNNgw9DTpxlmL2uelq
G4r3ojZFwENyu80AzfCwAzGXxblfilMS97AhrVNd53l+2V4LUdzdVNmpmRqiVd4j
Z+6I7fdePb7OfSHrr435C+2ThomM6ZlsoSgCpem6uzv/PBMB4vM5Abs+WOhPObqq
XfvEmzpFx+f4uBHxXDJ+5rVJAgUU4BOi+unVcZyL99zlzbnqhxUxPoTdDQWEoGoe
rp/Qi8g1y2y5OGFkogsr35I1zvxGCgkSlW1d+FSJFQ3IA8zk9FqjvKojTTvBJ/GH
+0qRbhmqoqWMA+q1UjLClj9eCv7ol8Yv3dOw69CNOcLEIAdlv835KYnrOOyONzTy
Atu4KMrxlPNKESF1UczmSLdl/9gFLMCSYW9hj3oHdGKi+g90PZzEKPcI6DWMg95c
3Mu/jwC0+50x7k1GtVDc/lkozvXUtMCDIWEBzmei245DfatX2up5opUGFM/isgQc
7CifDNqfpOTSnkZ47ShUa2JN6ARTkNXM5E26bWKfN+krRx54UelUlrLk/3+3aNyg
GlV21MkKAxnRN0nWvW/YQ9Cc8IjXqNQ2pY1Ak+JFZi/c7fJRjt22I0cnG12jHriH
KGVmUNBCqGbolyOVRhh93x4zjLLZpWr6Z5YABgkcG3KnAMXa+gauPm7l2pMHkFH6
1fG8m4Cspnf0pJuEQtSa9AE/7NaVblGAaMCqhfKaIJoa+nOqhF9eh6MS12+Ocy13
+akdnsBDWg6KS1UfLbyqAErix/A7yytUld894OFFS6/14CXEiLormIbSeJ7V5gkZ
nf6tldzm3aUcdPqm1yoBtQwWPpOoqU3CeE0255puwhRO+mx3/jy/gym3lxcFXSA9
kCu2U3Vo6fSejYX+mIt8kP7ZfD7lhBKTQJsQ4MMRXdHNhzAj1IH5gInKCI8t0Za3
AMJnA5wVxQCTShqaL2zov9ZxAvTMNsOxyj+ZT4kxRihumzQpvCd26ZYkpnakAvAF
bg1dUGX9oqoVuJQYrQdniwrmKHOGdAM3Sf5Fs8tjK1pr50UYeme8mR2GJdPe73Yp
OfkyBPLE2RYisVJDvvADbsjVnX+9ZbhyE9ntwDACfMNEQ5WHKZpbXFaN7X8fLHrY
kEOoH7/7iN95a9L4HFX/VSl0wpygeOBe/WyUqpn9rbKglGJ3xMrcGi87cJ8BmASd
faKjyu0cxYWbevWSEy6ncm6y46OgQWg/1Q69S8GZpHcAK8Uq3E7ywqrQuvPQVyZg
3BV3+3TF2r8OZRKoJXYFHviuijIUXCg0vPlxxj8D5xhchCZPAndvq6RIbpn54dPZ
Km6vtFUe0ALQpNWfdP2udy9tOEyjEPwT528DAD1P7V0eAxgDGE0oCM/AIK/WaEfg
vZ8z12jBRq75woL+rqEbKVSD6arUBVKXm40lNvUhf58mN9VY62VMDuoyWEweZi+P
TijzCedpZ2sGdefoivrPvsGlMEq6MPeie0pAzwwfZEwqZWpW70C89zOBU0UHvPpE
vKPpLq5rTguen77Q2FAJnTwhkXGdS8ag6PblCZgM2Wu9yqvbZwQBEGr4nhskc3oF
CBDh7BnrLN+dCpGoN2D3EuMDxvwDXUB0odqjLrl4Fb4nOAyNTW5uXYGZB4rl8Avf
SJ85/u4Z3BrlYfjZxfW/iQKV/ZjpPR5zrkxDNstULWB1xBxfNNICeLYlHqxb5Uww
iaPQ05+UFjjYRVuqm73fmGOA7Z6xHRajDV3xluSH0kyiPe3nDRFnJuTsVj/a2ML1
e547/1X/x36kQ+cM+Jm0UYZF9svvMlrbMzPKmKWnXYtBlhskAg8fGIGrXv5QUOrP
SWXej8n4jTaKsSSDvBJvFUAeU+18MMx2zinAFAM9TUPx1xnBg8xxqjkSgieJ8+q6
DUneY+WXBxAdwYTASKejC9niJsGorqVOwo+pFx4cvdzk1uPd7UyPawzn2AYiSYc4
l2SFG+Bib/bt8x2G1qzKY5QgHTuBzdEj/I90wFkFewwMMdYgEcFCBhrjCe0b5og6
cMqdOHRPYROnCONpY2cT66trgS8nKQnEUsp8rZOgdqnV/PeOGpqoy0OrUEcSKEn2
48ge5ZbtGqDDV3PtxabGkobrKUn8GViVhaGugGXwtDMudsdU6SJst6KNFcfs2fhm
4WFmCV0Q1RPWiEPjoX3m/gwNfUvQFg359ViEkVi/0LcsAKxhO4tR6clnsgkBdOEU
EclRgSbFlufYqkh1R1cPUpFdzuIcdqUgH2fx0CFIm0LDsBrddRYmg3sNvX02GSPI
R54HWCn8wVjTxn/PSLuP/3K8mnyjenNjNLUCeHrcZ1rA0i/zCLaOv7OUJRF7lDFU
pa1sb5CLGks4vo8i28GHaJCgjpHIKTJnL/w701BiHgzIShpWVb9DYk0zS3OYJEbk
71scURJ25DEetRV6YAZYbnm2b+VTaHBxg/M4eIBuOKlq8IySriPYG4uvCUCuz6I2
qjBHDHJgtDXGaYy3RKMfYXMFXvZ2NGo04YKEa6VkBTCg27JOotoC2KwXwwQ4s/0R
npHuVbAG4nvUBVDUSrnuclnm0Sz7okdSj+E7QipvHqeCxE1+5WgawconJ2ya6SnK
7MpXiuKoivHGUzbjpqvcBv5eteEvwo0eGK95ohTkszB4KD1NJQaGsNyI2yvWVtpN
HQByGNhi1C8K6T5F7g0sVtlXBXIUV1YhtPLqO0jH/UxtAf1RG6kuoGKp4rnXfvcX
AfdWsQANm2VE6FKIFi092aFXZblAQpR2fbp/dfs/LJx7L+m12Zmy0TCWlrTeHVWB
a72+ReNMN+Gl7uzKDA4rCyPYdDS9a9t7Od/BYgl0pKbQjmNQEGU7MqrGNWuchxOO
zIm2aNe5YC7kmxW+5NVUGf6seMsVMMscM9LG5/4Vf3NL0nsCxjnVRgydXL3MKdob
n1jKMfREC8JSp/25OMXPFhXoVJ5FJtHhIJHhE8Q3QudNxbipMHEBS9wTQ5HjRF1l
NibqaICR99A1LInPbhvjnfra5oZ1KKe6EBHavZdI+qOrv82pnCqkmaN0fD36SIx+
PFlSZuQfsIHab/onP5+fTab42yQK3CPFIdl7UcP7jqIUARSEt/SFlf5FbqkNgzHr
rfWpxc3QwWZygKQehWbJCT0j7j1XGRdOLny6CPGaK1PoHslpsw2VBtGdvdWLTFXv
l5xRW3bxK+r0g/D+67LmE8i9PSVs47dYHyuKhBAMhFeU7bkQLhKcA1RcwR21HDGH
C7WHNcY4LU2br9FPldKYE6L723Yzk6dTA25sHgoNjRbPROPh6b8V6Rk7mljZCXw+
dllqk/eRgHEtt9RP2bpkJtMxyEyOflYyaE42vVmA5hJCwgvG3SWZsc43Be9KN0d6
2gM69mxz8a0V9o8fW0DGLIbBL4yLmytX/PaPMH31nKyhgr2ORv7+SjpYb6rtrH/2
HcNnfzOtcJJVkVbK6oWWutey8KcN0pwRq2qUr1BeOEQoAflIYQpmj6klPA/3rMey
1woC4yD7WcYV6q/pwUC09TzcxjdW/w/ST/ghEkS/YxV27vheT6kMxUcsBXLpuvAR
vqScpDw6SsQgx6u5IhsKdNflhnZhwUvXaf5R6nCUOn1iMOt/ITvD+kBSHK7VUUFg
Mm9jsR7nl6T1Q4Jj0hkuxpKhJT4WsdaVihJPEqvp562nukQGpziTUWaIzTkb2l05
H7XZ+gBzgmUym4m9ORIRGkLud1t5tpeThcDgceYrjJC5H3HnQrW8xsBT2y/HZVSk
ELdqzewDA6N2or26i7+6WSYuyNdW0g+VvRGzptcQf2USGzB4Q7NJXhx+etA+2n3L
zXxsI5xRqKFVqrurBLZ1uD1KesbzEgz5IEyOAhyFKEb06nM41A0reWUFMkHW1vHc
5tpjhXYMZ83REQDbACFXwHWD6UO0V70L7CKGD+FTQcNenjaGq1TnzE/RmhZkYtHj
KDy7Taq8qoaBY1R+LfKsluX8WzmbsJE2GjGp9Won9jjq59x5SanW9PID0X+Lm7XP
xcEVFCUWgLOaOt8xUtGyYIHVmHI8gFXNAzmdTbQXxW+1dYVTKHP+JDs9imvLe8ae
ER8d2QHnzu9h8w379bR4bAKayVDgM7Y3LYJA7rI8qK929bAjkNCxez75yVNHrJP2
UA5AQy3J+K4Nupn9gfQrtfwf/B1o7FfLsaX/kzNc4bAnOf+plQXrFQ/rPN8MSNh2
DZ0wFPmjbOMmFY2HvtAViLAsYmgugLHyD0lGSQs18Z3Mfarrg0wSzsjA8to0rLqp
C20A/mm0Dd5ATZIrXB9ydgyGAeipwJ7P03Hg14Bqp19oQC1iwmJf15vTYVes5gGN
E05GW7tDsykZZnurpO8/NxPodl1/fDtkax4REfxIsRrhTsthgFR2FGn91pMXaOnZ
lUqiBi2B/PZZYWQhTl23ZsYLYWRYIt4GqrJPnKXMJkhcyWhYepwDRTFdQcJH/Tdr
+aDO6+Ovs0/rnLpbHdxDDQkADkf5MGMIguEblzpzZ/Lt51O6DRwN2VGm+1Ms4z8u
KUGALDZ4NF+b2YdrGyjJPeoE66gNw0ua3uZE7Mys4XmJLGyaSsPkP+uVWZUZ9YFV
Mz1wfv+MBVuVMeEfbk8J9q+hAlAWmLVFiIOnR5AXq2/evtOiftIFNEglJNktkxav
h6mAuyPX3jOhRV96rUUnfSUGb1Oy1Q5uD3IIH1bbiazZhZghJm3b2V+bERprQWfK
S3K8RLORIRfBeOuYP/mlW1guAOtpJS//s6iAXUtO2WVZqP7QyY6sBbmzZusWPn7u
xXbEQjNKYIVxxnOhYrLQq4lfxi4KGDfRW2h0Tv5QeQldoXGcTyf531XtM3cSMLHS
/u66i+I4HLjOZRkyHlrMjOMRZHrNRYXrltYMTiTA21A7aqVoCgZGrHkiwn4HBZlH
E60kvL8CptPi0HV34YOo4CkNZLFqIBo/JXXuzw0JbyB9NuFFndJf4rqA9qOXREIn
r5qu8m6b3VuKJ7MrdQ37WLJiZMUET0S0g96WHDZmT1pXOnKdqctb0qaMGAzwAWKD
wMKAbjlJAz9qiniiefEge/b/v0eYV/yYhvNr7Oj4oK/cPm2hDvm4j8YIuaSBEViM
nAhNduKqnjUUif+494VEuvsNQh16C6t15ltybxw0QMkWm0UwM3AfTfoetOjuNGPy
NYEyGY9VFv3KyPqcFxxKep+WxK9eyt8VksMuZdRHVFLqT9v9XGzfg7zE4STk8DJy
Crwbh8bTBJbP9r67M23Ls2QRvRZSr6jdr4kmwyevKrzgkhScUKlaK3uekEhthirI
b+QkGhggNvTTX2h3Yxy2DwJR+NZm0Din+Fk8Jurwc2WM05qQj9VaRLk1+Zw6MVh5
zvaW2LGsybLJ6KV6ulK8WAH5ADSE5N2jjSrOUVbMU3fXDi1blTh3EHumAn60bCgb
CQFczKZlrIyL98ttsAI/oIO6tu6zz57GIztYkjkr7ppWRLJC/v3y4J7VUpPbv4EK
JMjBspGZqT09FzY76CyNIozg+2gvDI/WFH/0Rg7S4cxpmnOCM4loKJtb/ntQQSRe
ubSaIY2KjAc/FN28pLInQaT0q2Bd7fpYARtbYtKQyY/WmUZPQjlcHx9ZI3gBHPh6
cQISbN82H/EaGft6jZzJiQNNc5K7BCNuK/qHBPPe7Lf/BEKCT0McaWjXL3Ei5b7Z
HYMLVVxLylobsA3/KRrzHQqp2lSHdRSTt9A/Qa8mXJKAgKLghAA+5HQTHsiw32GL
Q8DYiJAhTrPIniDndOl0GYPzWu5D7huNSL7xQe+d9onBIyWFS6JWT0txSFcyJeEn
n65fH0wkUInN8bMGdiXoAvG7DLBeEoD/VE9hXFPPvXA+CnIxIiArgNth8J55oZFV
CGUetjiAZSyYUVT6mrdOlrYeBA5tdyRx66ajJXwQP5oSooM3JbhJsxCdnIc5nxHe
LebJWEqLKUL8EjQ5d6pL1oJ+SAL2yd+Iz2Ho6DnjYny5pQiHBLn9p0sU7uL8hGB0
1KESrjapGXVpntCSBF9ooPC08+WJ0iu3/zHgSytisGnREUIAY0uV3kdSCwbH/Dhe
BKHO75239j4CDY0khaJ5CYgy7yDrXnapubpw0uUfHnuqLKd8GOUgNtxHmeP3GP5k
iXtUHklorJBpgXVYyJs243Bc2VWKe79+HPhQsVJzNEVAsSZi20r5/pCe9oA2zAy6
upoyiwp9dbj51VmLAt8QHgOrAlkv5lx5DGwdMh7dVppn1GESE12VhzSW4ctShtie
o9KYxbF3CovwKyAb7q1mG/M4RyX9+nd85bmQ2ieaWyhuebtp2YvDkanQhcEAiTva
EBhvX3CjGtb1AsktqfuiHM+5zESI4b1cLD2uWWEM49lYohWSxpAp3035Sfcu2liR
bP//Fw0l7OLzSOHLPHaPuQORujO3uVLc82sy+3PSatiyJROaWbjA4h7gXVSjxZ5U
DpC6b83+DhhXVg24VVpxRbpXTafHaEzF8AHYZmU/QwFL0Xm9XNIiYl2UK24YDgcN
rJhPnCyK58kPc4F3TXmDOvMLPNTABp2l2/M4p9yg5DKOiXKybsFi8L1AyqgVLgZy
R8+sGxz9v32dA0IqQsTcsqbF0yM/ajsrSBXr5c/9QH6GYjo1yyZ9feuTN9nXqfFU
STEyfl2gbMp0pL1bIF3P8pV3CcnD1RtW2cjd9VjRovOfniI3tDvtcdVs+dcdOnJN
gF1/Eyn7U1esAgfgeFQIMERMQEsCDfhx/h3mD1VjlMjBteRffewIB1MqGuQGu1Nn
9IQX0EODEsMhh8zczoMhP+pQ7BerHkU4vYP5/E/z5pfBEyVvTyKwLTBOOGpKTowv
0Lh1eOz64rU5H+gOHmrc78/fj84FnBsPyzAannrVwVD55i0Mtrw5ie+K6j2XS7+C
+mKm1T+GagfP9LLVGazczpGq0sPT/gQAAqZDbDOJ/2/uOAKPAtaR11fGaXCBbCco
9ufMYStrFxqFj2Ag60XsCRqYIEX4CxqDF1Vn9h2Rzn4Q/MQeqi62m7454ojExXTY
4i6sI9vkux51q8YtAZUaYcWh5Oy7j1XNoZEXhKZSvO36dmpP3bMa3Zke9+GdGW4x
9KDP2j5/kP4SINZJltRz+3VRjNvAx5jpVAQACmVguQLCOHv8dyLYLRD0SUKBQN+L
UIWrV3h0NwbXYMq0f9ckl5SI65fS07mrbEru12qME5kQN/GnJHFHJ3LZ7WtwaBTJ
+zVltErsAW38cGMD3cgf6ALKKi2w4PSx4nyrUkT5k4AD+oPaw7t0exVhpU4i8Ou6
YvkIKo+QtipRTG4Vtm6GzqsWDAB04ICI6wRoymE0N6b4DjdQ2wyDJft7BUUN9wcu
PvGYmkq4/uwGMomjJGxIaJ/qerUP6+PrCd2UVyEQfje1IZF90kTwxjJzWbe/qGAc
Jxn2q69IacGRL/OprK+Z2HLar48XoUCs+zZjvIl7WfVUzRx/AUuzCrZa4ecgV2G0
Ggop9wkLYeQVT0nOJAw+ikNDnP8Djl6fPg0+chKZyXDAgaAVwELCVuEV9BKLulMU
ymjxi6rxCck5sQJKKx8Hkc2MTX9R+aiX8bRJlVgo07e3o5LrblhtUOTD/pqTeNs0
PHbDPerVMEz6aKmPbBsaELwtNa9aQx4DDxnSGwHrIU4w17YUs0mqaXzP90sxtgI2
WiAIasxikeRqkSafSCiKfXtnkz6X1WEWhLzn6TFaM42DBNhX+C+wHz8bOLMh8r+t
OhXSux8vymmG5VcDVuX9OsQRpqaS2CDTQz+y3AxOUM/a7a0TiCil5AOcfDjAqpuq
PYjbAN5hSRNE3Nb2a68Qg4QR13WdKeV2K6kHNa1NSlAikBnJD/5Eq07OQD4wl1Kn
IzqKoHPYnrig9+YvsntMqmw2XnJcOgDFdz48ttL3KtlfokAMhf2t67TNhrGaokPB
qtQEjPVLIrQKgtC9VRxjmW/0xYI5J5aUoONFPu4Rpk0D1TtsiXolRpUf2YKcfusb
5GYgRFJbflbp2vdFyG5Vc0Gybj1KmNBH9HSoyUOtnM7jNydkLdeLQefosOKoNEqf
5cK3hAiv+BbLXlUcHnJBja9sWaGeb1jZmxbt6n5C8HdDLo4pcy2egEcKdCuBKCo6
uuFQf9qDdbNQgwqna1zNIqRGI35CiHx0ZGSaVVwmx840ebVMgu2McLYTsLXq4CJr
GsWmaQbbROIFiBLk24HJlhYo+T7ID/EH5xKCbly+a6BkwN9SXyTz2xH0uUQA67/A
XXnxAaa/BUDUCiLQdyG3Dd+rKYbuGgiP7sAaj9qU+dZ8QS9DQUO2WYbwD+yx82lz
DQ/hSMwvd7Pe/HcnYAwOKA1ZBGf0HPYwo0/kmm+k5sxJ2O++jZZ4RUdafQZ4LvL8
BpX1eSJf4xTPoOTHlt9Kwwqz7DcmUF9tS425/j5cnmGwfrK6LboluekMpddUVoeW
TEq3cCRkY4xkPcu69cvOOak0pQJxeWdZI2zXOcvHp+q03kcppki/RddOR38u9abg
93oP6e93+gaPbtQ8JpQu7WkBUf6cTcZu5n7AXlkbLBIuNbA0poKPVOVFrdarZ7fS
btgcN1I2oMBLcUFvEgzbMf0nVBgoEusMxm5m6zP5lpQ4zbV5O+YJTD6+itgy0vm2
ezW4HoTkrtbxe/vgUVTwabL+YY6UsWwNFWY1imYXVsPdAVp/zPlWvF5wstiA3cFQ
iNCzAsfun6zQgrwgxNTuo/Cw8st7UUh+hTORsrmM9+sn/tlFY8hK29HgCkNAEtmK
9yn80ZdzhOk7/LpHZHZ+7ZiwwtPtHba0ABu5NDA1CjrX4nhGyzlb5ikdPlcethGV
8pJ9t4zmqTpUM4xD/tEUKxcfjZ2Rkv/1af4WF21N+HL395oGH6iRulzTqXS4aAD4
ZzXVcocH+PblL9yMFL42qNAbEB93vAj0HCX5UfyZ3VZhFRVP9eXFeDL/R7KZoBXF
fN0Z6AWG7llj7yr0GRkZoIvaqU0Geb+FGRwlXmfwihBmioIhCZa0ibLbiWHm4WE0
Mm0JH1XpQh7IPdrEaoU5Cd3nrev0SNGO+5RYxhqxvsrPp9xBZRxefOAEB6lBOQeL
KWhFYaVT98aaUVq2ymWOQ5JNCvE7jEMGhncD7w736GbPOb9hWIAVklbEgOrlCij1
0Re47aa85/xptepnyoM4wVJL0QXsWmifMwt1VL9D1uMCgOSrY5LEvuew37FwM0+4
Id0zQv344oUNF4Xqo8kc2tvMZ36ICniE0LbdpXOmJTB01vxCjPS9Bj+Q2+EcxvDY
r+ZY0HOIr5S0zV+6iAIu+jff1hT4b3arj5dwDThpfLiDSCLYy7XCXYkHjG2dwf/R
SKEi8AMdLgqIsvxqd4AMNLVDH3BBp72EXPI83BCkqco+Su2QR1L3Q2uaTVlcKHU6
ZMIUVWQ+s/rjA5clgaUnoSchhG5b4HDjbxa6ULHtN9mHA9GFkHbYKkXisCPI7my5
BOeqsGhJgW5GQVC9jeEXHA4ctXdUWwDVvkuSkUeitlqRrOrEPHlikiNMWld1sPuN
qc4znnTK32E6Ij8UaSrFUhc32vZQlTAz3vZa89UVC3EWOeZPYd+8T1GcLfOdYlYe
lYGfOOz9Or9tNap9pFkRKT727TwcrEg23UJKixwCY4OF0ub5V0o0HkrnKCTbK6H3
Rx0G0uY3rOk9sMynDNT1Dgyym/L3Q6QiIWlN0k9sgD16l5cgifHPAak3clg/97xW
MeekWiMG3l8IcNuRBn+qZBmYj+KyzEIqgpXyZ1tnvRsI9oERky6lj5tQYXD1Hbmi
+f5DUjfcKgdcr8EejMLNMnempZba1HVZ0+VUALtUUb8MFAiIpQbd4Vz1s/i4r2Ed
KboD34lx4U5t2h1xkXa64b/5bsa0oQeFAbyWOWODbRpATrLMs23nZapAIMnXgT1E
Uj1OgvgrQ/giKx3jUC0cEWgMzSbrHbxhhFAl/z3bjL3mn4X5PzIf7x+gqjfELDyd
dHqOUj/E81H8Yx4yrnnd0w7u1Ia06l/B8EWrkP8sH7MLBMfzQP8Uj/jov/ZE9U6G
9UZR7uM8+d//adRjZmiX37IBIOEPn8esxy5+NoO4Zud7jWF5Mj5ByzlBRbdzKPub
WJ+b2BJCdOXsbYbfGwu+zPVR8bmMw2Yd+X88dSiJSsSyQDasVwYU2vg94d/GsqdT
waxQW2o2tSU1f7LKkyrUdJN63LXQJbTNDPAxIHgbY19AQOdImPKvJs6oqq4kaZVv
T/u8767/wEFwfad50YfqNd03QjLsTaKm28UiwcOxlA7mt953VSfLf8bXHjqLEO+E
jS2dJ53qrtrPwANOiYata5mg5PEEXQMhbB62Xi+vbHwAKlrvCSefAkqFhZCb2Ox6
xy9nxRsWBlcEyeDAJmeoCNlM8mhE2Wp9ZliPPnbF2wEQ4ro50hOQon+eyoUneszY
CPgLNl7OSICUL3bDMGUE2pDesNOOp9E+1hUhXK+f/iVDarlmDayu6hgLJsEb2RFZ
uLefkAEWNDVFqIw65KhmXRtMJ/E4hRylTYhalg4unElg6psC+j5rXDzvn7+vtByJ
iwLkWKtzS7ZaNM75Eht+Gbk+msFfxCU43FkEr5T7LihpLgcax8EOgdMZ00k0y+/Y
Kz/WoOe1P6lmY1aOKculcFeQccS7uZG27IAxR5RttZsC3fLqm3O7SLITz93gRvR4
jUal5OcP4f+YU1wbZ4tFszeyYTHzFXRUc1Txd1GyDgVIjGrCABtkGsOBy6RyzAQm
a7e8nXAOuUuM+MRcTe8QX3Ls3BWzwNz0BbQMlVKhOXo1bmp7S2ZSoX31rPFguzSK
Fb3uoDQDN1zV++r8N4lO8g6jN5iQ2Ak86dMx211QeViDqZk5xmDbJQ+7ZlsfwTwO
AljJ1J13yG+presuQgEErPmqHWnN1zSnyrP4jf/gSdytaMqvQcuOLf8BW2S3VK1g
nqXqrRQQfmdkA/pxkHpQc2V43p+pg8n/6pgCazOKZYIx7iFB/cOkpDE66kZrkvhW
PRshZEJTixhvyqAqcKxCm4RX+Tiaoq3/21cyPTFEZJpUK5g4h2tvXuy945oVIiWq
EnuBSFLnYQcJ5jSRsYa61i9IQmqsYZ5nLu2i1Wr3cBxQpZwML+ulBP9hBbNuLR/q
ONKbtyQXE97MUJVnFbhAnrWtzv5kZERxT5J0Q//Lky9pM+XvKmpNqVUaqc1Pon80
E20Bj2LAASUcHGu4CkoLW9mVyHpaiy26rkRsEifcuQ7DWj0DDBV+3xqLwtTECHY7
lxAoEsEqp4NGIEnBCRIcmK0z1pcr4hJcT75oRFSmXkoGJKt2bnVNzCuQuXUMaStr
z5lfjrrnGMGiY8SIa1alMI8cqzQfI4AmahotOjchTX06dXnyKsd9MCFpkmOteJVv
MrImVHtsIzfT9g0RdrA0gpc8+s4Ekgej5X6DYHKPvjtG5L5ICcLtpfHNSzA0XQnd
VyeW0RwGkzuHwmYzgqcpQ0sdpN1k5Sype5txt7VanOZ1D2mv5GIAi1FD4LQ6lP+r
zG//fA2rVO44TcBeVEaTIEyimPPOyDPLkR1A77yeUrhOxwLlhUkBSDCMd2UKZ3Gm
wai3t/fkes5axAGrP01wXssrwWoM7n8uY5w4trVOASSzpYDtU17Nw0rbn77Io4su
7GIrkWCJA3RYo5xyeEWMuVdFqxXmg4lETTQ9248oY+BiDoA66/UhyEUodHHZcXxn
orw4PHBcQyWJI/XRCzeCvt+XTdELTSa2olgLH0aMm98rU0wPLIynb/6WQt76Ctst
6YD1D/InyUz1Q+4HwbP7piID8Ue8vTV0LBlcWPUyJj83tlQXB1pTTlo8EeNENDSd
zTHt5JiJFWGdsNVI7lnxz9SlCJwgrY6/TtstQ86jQhGzXyhkFk6BkNc5CAEJ9R9Z
krfjkOjf+pUCtPJCXz0F14Q1Cs6vchww1i8Ym11hiKmebbsblHZM6CJ5D043zTLh
FBu9g2v/L4HWIXyz1Sgv/nc0CL+AsMRF3eTNAYMRSsbDm6QcPIiKnswJYoWB8zdQ
qI6I04wg8W7iU8OchUtZUTMK+MgzgQ1oCFqoR1O2uYxddS57AUT/SfOyUsWKHXax
eoBh7WVzau2ZG96LcjakBOqF1mtTn1p303RMbYVDmxx0e6cYpyCXovcRCytl+2FA
WDUL9oE6Jr1S+lNUqH7MIVK1cKUWT9tQx0vJdxuc1WM2Q1RRWC5peFn/Uzeh+Zx9
OlW7d/l4XIAS880XL9hvzzH/R1JIuPSxpK5jlFFBYLVmVlL0hmL8mLQWlJFTgFZ7
YZhG0bvtbTLiVygUKxuIXrsh/SwqzjYGlXGmqlCAvTk10ym5tE78e0Z5n94HbMsR
JcGzugagMsFq9n7FxTLrsz+GugCsEJCMDCo1fRi8datXyJIygK4F5a+Z8QxDdt9E
eFi+heuGvqmrxJW7DKdBJi1b83/yQWxVbq8+N6KlujmYeh3GFqYOJ6C4LE+U8vx6
6ELq3627NqYrST52zFWjJsac8xiTRlSfwASjqr5crcZlGQTY4a5UqAPyiu2vlej4
8mJIbuL5E8NfYZenl7C5I5ru4Cl4NFRQbI6Z3Gpz18Zh8laESKz3fk6HdgYhuhKT
XyG0fBYRo5RgW2Ijo40ITgi0M/Udd1UUP/+6Ie8j3NlWV1opvCEGQ7ChJBWF7Q17
LLP+qTD2jkCoYRVJ7Ooa6StCqT9F37SxTJUUw0fYgOXR9lH3iHD99wfWJAlHQ4AU
UYgTvaeZNhqUBPE/EVCs4LOAc3SDhhqB1+0Bot6b6xoEjfuXsIQcbzbCcCrRZKOj
KZTMBUXpbnK7+czyHN39UJYzmOunjwSn2+/15KXUDtCl3G7UH0RuauGj9WpF+Sp1
xuu7h6t6KXmFTgIxcJrVGIrkrtUw9SY+6p7hpwvSlfOc8ohbtIlna36w+DGUcutB
V38r7CaVs/fivGQPfNnxKKRMjd9mK+8uktjal7O6bciHkcSMyq5nV/zlKuoMtHQS
cmY3vQ41GGOWIAmVN/Xo7rjmpjKoCKinLD5z7wye7FBT4T3jpyS09aPkuKNqDAPN
gEpb4Lfm3veRy6rJffyxuSjGWtOPKOloOPrg6alUUd07rE0CBWigX8m/CFKANBKd
e6iGoSAyxCTcl82wcuJYR7qyfo+vsHO3FwZPn7zA90VNJpT7GUlSjP8j/4gDIZCL
nz7Bgqe36QY0mErLJnOlWZbP9r4XzDUaVb18MhWkr4DvGOft/g5TdxBESPa3L/C3
VWU7QMEjYsfPPIDXWI+Osz+CrDDptdu/A7S9usJuHd+f5cE1VJ2OtDTxBPE0z9q6
SZ/ZIh+OEiNsgIXoGOzc3guLquNse3qkm79EnsKgTAcyoPr0xomsshXGfJ2kfpxO
+PZu8wnpTcnmXFcjeAy/MQhasvUe6+VBYpDW5eyUTESPOpv/bqF1AYef62zCC+QA
dtUH7MvDVg6c6isEezYZ2csnvhHcN2M/Aly5xOWuEmJQt2fRkzUXagWWB74kJsmw
jiX3ExR/Gmql/S4CUH2oPoV1dRhDy1KKheAFLL6So1e+SrOBZ/3XRVVWZCfRALsU
dYZrlliDMa6cwfWsSQeN4e++acpkx9smvp5uZ4+Mhiewzzl3FpLezWjpMvmwMFQH
q8hteldU02h+VfRj00h6iFHF0AzKSQrAkr9uzA5dJ4nGbNxAr8sRbyuqfIQUlJV0
dvL613KYBNAZyUcRZJASol/OVKu9d9/Fy1PUHiWxj0xKH5pbgumihrS7ecdS3GVD
Po7RgUttRqkpoRBg2wH7UHbWIX2wYRoeXsrs0FMHacmzGVaJL+PC8Bq9XZJ03fBq
j1cK0fLlrWo4hZP5QrtdWI8CFHXmwhmbIQTyDIDdL9vG0w0pGMCq6xwvc8x+03tp
+3lFzg90yAK4VnIwlBiYinEsGvZcNBuIu5v/xxvPpKPbRpJaM1F8fpA2z7LMBmoF
vbStAuH8iVN904ct9FRDfdgRCmepDxn+nykfijtz+UQTnvBkx7MO4bzQ5UrUcrF7
Ke+80zESKvpOaaGiByZUVYgfi41Y030nyk8ZRxJKz34gRmM2E3zH8DCcu7wOcr4+
VBrFKJo14BsKoxdvzh7t3kwbJ41xk2XNs9S7afoeaLWyasjp6ijOXUn4v3j/JJ0J
bATSFfauBmi8ltKMD7HupF29gd/6graYE46ydIQ4D+L8RIzUDQ9HZFok82KVW6qE
xztI5d5SgfN6CoMAnI1EpaaoimW2UGsrYgLb0y2PVDJpuo/fnKgaGrT2pTBrJfaF
bt7NZ1FAEMuFhol1/2TyVam2qI2Nd55T8wrUfjAlp4emsHgnNgbQydCdsetYcwi/
Dy+tHTYrZUIZHPBMDpjTwZXgX7lTkVoQBfRtvzwc7zw53n5ljId9pT8rNEmrVhVi
pxH/Aq7mWIblDRRkPV6BU3iCAol+a9sdV2Lek3F3LZhN8rDwpztpaB0rx4ZLHZWU
qzqphUo0pBrD966HB1ThmyWvbINKN+xj8SPDNfCHQjt2tYNxH5+i4KA6x6XIyPhH
UglDMB39+VJ2wjnRKE1YeQo1gMnpNg1qceopGNrFPZP2SZUnJY2SG62DLforzALX
LcY4EFtx+u6nREsHmS9PGr3AK7w5p8Lzn9DxhI6gKL6iOtnm4qUBgKQ9O3MlMFrb
5Cl2OVQuHZZ3FsHW4bzvmA+cxPwCcPp+lTcq+uC/iJkdQPv2eIRDxmQvjRCGv8R1
+iA6LgEB3nzk0B6JEK9RWNd3d33O5LMcng4AasWc+RllSK9vkG8ElQnMZZSpJ3Xs
tKZ4f+QjbmWzMK20unbH/yRKBUQDoiTULmPd9IkNwrOawA9/J8lD1x2Zj+YWaMin
iAdsdrerfTR+RR/Gu0EmUno8adr15ClQfsHTlWOg7YKdI1mpQ4HNY5Uv4TtNyyfD
WgGZHqS0VmRbJ9+yM6OWUDBdcfUeObr7zgco7I9P9v9zKe0ydZKMJtdWLyJ1fvLJ
NgOEtDxixReehLB62hOJRy0oUOwuqFp8GXJT4XYAE9eOjFACf47+ilN0VIrH4OEo
JZdpbichaM2SWhfuiatvhdEpqiE5sGb9guLRNJlTYGYW/AeCEi3KjVTcCgDktSBF
z0q+RDHp/1+h7ztwGKLJtw1gfwJuukJLBOKpy7OsB01amxq4RvS4X7A+j6cq2U9F
ur22eaMKMQlpK2xgHm1WuEOxRNWm4OHNPqgUASzVItS3m4+r0rO4eDySdonOtopA
mVRXnfKTvscz2OCjNGfPNPD4zHVdAhPyi9gPBMOM6ZmcN3bumVyB/szmnpSQSv/S
k1T9fTKVeVrsNrABI6/K0+H2TwyXJvX18NPzKTXye4+Zbsw/EUJ2K34RP/+Z2/Rv
JNNRA8Gq1X+AHyLZec9PTdAB3Ic2xjVH8FSoeeWTGh75QsVoQyQXSE7zFUjxHPST
xgjiP+xpwjYN1OZhPQkfHbk3ggSu0d6XUgz4YD0S+NYTwa6k5geM3GIi0rGAJY3K
cGJKu/bKKp+o1pRrMgaRVoj20o0VLAOrv9LEh4YKAuVMfckK973h9NIucChXZeD2
lsIa5tcT/vc4gq4wpuo4EDe3D/9rTeSGGXZk4Qkt19MAUbbjrZ9pVjoVZa0wAfg+
LVqM9Kl2ToWc2Z8tmBcR9QI902sNcxFWI7VK+nWYBPjzjezMOzwLsO2VubBAj4WB
Iob1UoiaKcx8h38JVEz/p+Kb9rP+aNE2r4fC7DUKX4TGLstg2QYO4tcpEqgoRT4D
+m/yl1tCfuR05RMTOsG89M629DVtCdPe1zCHGoHCqT0Hd85AeyZYbX5edUe9/zW0
a+qb3kbND3JHC2AvAoyh4H2/VvjhDleMJLMBu4Dgz6GCKbE+24if6zakpF7G+pRt
7V8iePiPuL/gblVuzNf6NSL+13UOBBWY0NtvplaGGjquHo5DvPUMWbFt/uOubNiy
Nq2/sgc6DCeP/a+NQXDqBMs8W11uvEr9jglWH0UPeDJLxz64HdHUNdHIri0WVP4M
93+WD+uQrKRJ6A/54l2FWEPYo97+NGkJfkP/OUZ4712Vn+KOPnpG+QMZOlAmXkHp
h5m0Zxxfr8wV5X3xW6C+D0I8vSzglZrkvi/W/gT3jHWsbVpNyT7CQoNE0hxv7mmQ
6dsAIPI2KqCb50cMzACdtDwRoeh9HuxQmu2M65eOJb0K5EqMeZreOSaIX9PsTqTi
HDEg8FN63gGdyoVBOQqkFi6xkTBO7N9Ux53Ua4RCTPJOunwhLHgUngDsqTCuUqPQ
Qv8R9SMdPURiTvMur6crPJnY3HKeQW9B0Cf7V6ti8LI9/7FqaSWTewq1bb0y4ncF
oyqbOmCn2FAGcEk8LcUelsXlyGxjl+c9Tlq+rqNagCqR+02zcSB2snF0vaLjkyFX
YTIarcEnCrFVbHELq8MLOt1nk4VPUC1fzOzAQw/WujZW1AKQTfQEJbgk1ztKxTH/
GUGKRTyqgMqamemJlauuj2JaICIp5eitCUKrSnx3lIAV8jmJNYvLKZ8pONMnmItn
J9TpXzZW9pJ020q9ioJY33DxqgtXRIYx+uS/4KtqdrhV3rFjaoLaoF8Fu0oH7RDQ
v7/pC5E/PTv6XCdm/FGU3NuH0A3x0/8Ekddu/woU8IOsojuC+RxJ9kZ0wCiPEL4C
QvoVd8dBR5M4fXKi2ai5bFChBd+rLlf+7qOb5FPa4YyexLApAHIde0mS3upuYmp+
GCM7aDD7a+A9VkG/n1DwjONUYFi8qlU2AjXyk1bFEgiSRDKAajr47vh/Og9I1hTI
mszzAKfEuEt3LgMK80VV8fZ7k+X9qPGc/Y/vH69Hy1K6fiTwn90aoj08oTq1cDer
usuc5hyK6aehW0vUVynu3xBwdBNl5ehzcoHbsq8J25ZxqWpQxTOOk197UmLEoDR8
G0/+MiFRdyQrwj614Tjcea0NAyqRBOXgKx6rNIgh+2dZW7Ougbs4EqPYTyOWWBr7
mARymnVPm6YGq3dQNrRafIFGHUO4Ujf2i4tH22qVsT4Wi9XWRJRHPr0v5dS5j1ps
dzSl5TfBoDgxGSLnPcxcQ9CsNffkwgKpH6LNEAF3oyJ5jSvBl1j7yhlaYVyKXSvV
4K89UhXts6Xs5S2jHllDrkPcxAFoOkg5wdnOY6rKMIImfJtgzXpANFkJsXnto8XP
LrepjdlDN8arVFfQLamRofqretyIPZK4yts1ry5lReYysQ+oXWFRuUPcEKwfoECH
D+AL4WINn+9MUmDgjFzrP7RtQVIMOjHqVASKq+1i6FbD4hRz85PFpgn6SkUhgeNi
HTGxpz29Z+6455Myl28UT6XNiF7PVm15CMjhkpK5bCaIhLG/zaNzC1CIxCUGVN5n
aPl0cCHTa0M3ZAPisUVhTH56rS6tfDR89JzFENkgL0EWGAfBphH2ovGKXPkE1WoG
J3BxKiGu2EYeDTub4z+UhYBq5VhQY7DVapJgqI/WtimcbwQe0uIJ8lDhV9vVAz34
yaG6Wme2hU0k6PAdUYMslBHoB91Qc1a+ld/bCk6Vyz/4pCesFVupnIF13o/BKgAw
/73dIxtAgJg4TwnsqafMgix7BxHoZ6FabjkluNxIthESWB2LiXZhmByrzASmcaby
lFIl/6hlFdhLk00/Ox15a6JC12Se+ZIEILTmZrMBVPCuQY1EexH32j07TI68RVyS
fyH9RhZkXBOE2ubkFefos/dEgVXY8078fyJi1fojltOhe/GphZHbR0ySEN/h71cI
Cj1+re+i7z3AJY+rJhKB37h/IrQ/4d74RHVtyENlFWEjUxon34VvhaEtbsuQG27g
wIHCjCptIbU3mdYFfvzGo3T4o6eGj0N8ZBvlVUYfSelzUlDJ2UoXuPFf6j/Thql0
OFUWh0U11qtndNHBwkJ2z47MwEv077+sebMxOfWTa7oldfDvt6/1pIHNaMpod5gJ
08SA84kvVZ//US7tytGXDJ7vr+46t0MTx2fhyfqxxANWsDTcJ00ARZtdFrLxnLh/
aoG+PODt5tVbwjyBXCHI8Wg36+flhj1qeMWFzgDtLWV8fmWOycURubd7XkcGQ68F
99N3v/sQIukRDBv+QTkSc/iOawkU6gUCZKtAZIuSk/9Czd8fvHXr9dtK591j9A7w
FhjSaFumvzURLtuBVtY/jSLBm1LBa2E2n6YQlzcjdn4SBmYXt52L2UqkX5xvDJPY
IuyG2tasXkhaTibBejj49Cix3fr3uYfRLf7/lTmPlkudsUqE4g3OpsoAdmseTeQq
Encb1tX0mbzjHsDQDKGuvjhBBnmJc2dtb5fvOpB3vofnO8fZRNfXMcGZExC+g+nm
iDEb3VgGy1XQ+789N0drC54vKiYOuduOMPiMbjlT8tYLFBQGdQrQ2/3MZIs87lCY
mlaa7A1aGXjBwHBKslQfoTsaQcshK7Ii4hhEqVCAcLUfWnQFcNHcqqMUZKBoKDxB
ijUlCulxjKCrbR2K+WHdUK+GrGqDPXL3hkJnKKuP+y9lv9ljQnG9LMcl2jyfEgJp
rK09P0UPc6eLRycveTRwXq4M3x81/9/MUEzK33HLCMWFM95iIWKiy+bSmEZxB6zw
i/N0MUmqFWbfLVukxx4hDXQoSl7wA1e7pB4/Y2IqcAW8qzCv5dOUARBF/7xZO4Xh
Zc2XMrbeDO1Oc0GScDV/JBByOy4+LlxLyrLNYvjz62sbaK00dgdk+xZfDzmxnvCo
6FOCRCG+dxKdkhzppp9BxxR4kQ/nGUST+WvxVHkyI8LEi7ZEjs8yXQ3M499Oh1aZ
NIneLreaNxR48PehIFYSOst9YBmPE30fExzM/9tSCUJqwrCLw+e0hiEmjoSInSnt
p1wx4kUP4kSsO1nEcgZgWqRgrOxpxOe01qL+L/c+0seI+UjsdqhRoqgihHE1jXAs
o3m199Tvnv8y9TgSqERHZdrrWh4AwYE4ouU4VcXvjoOKwomHkFioYxATH2Tazl9S
jGD7Mnd1OjHKqHcMKexDkJgXOJK3+LCmcGRzoFYzfb484+6Xi7+KoDW9rsnntIjq
x+cWsbx7OU0fOkll7/LFXZGA2I6bfqlPal2lVJ3FsikA1jwYYHzPs9XB70bEQNsx
/ovFWoJbWAex84Tl2vlZoWB+r2RQGtVBhQwLEcKw6eovpPUqtw9xxO+FVg3dxpQC
n22T7Y1UGBr/5HNtXxd71hGmWFGqZaM5ksmTAeMjNzJ17LF5mrvFkflCtx8dV2OE
46JoHnaX4PvVAMbu9xoUSoKCGRxvpfxrp+VgziHay+7xKjxjepHcpdjKDn+MvczB
iU3jnzCMMu/NV6GfT+mUsJzQn/9+WTaDD3ZeNZBkG702jhFbdGUfC48nprJVwec+
7pCZc3ZVG/Nj+9ZTaIg7yIhtWqlhXtPVI5nG0HOlh0euXOIpdNC3GA2cOn6voLyJ
DUXQxXIdlSl1wqt5hNrTMHAA78hn2c1zPRm5bCU6bc/qGz7q8HZc16BFuJShSpTd
Tq9Yfu+kv2FYZqlt0O0UAs5RLjRYRuEHR2csDkICnKkEUwAWMpVfMBmPd6uLJCRX
BY2Z85/vqjf+Hpw/ExISjFtOngK+oj5a9MLygieGkcbgORtXH9C61ByGdU7aO4KS
GSFm056SiyusWlQKzyDly91YRTmyUQRwjamEU//JhfDfizxCicCiycY721Hdek99
ftNd4LeH4wNVmgihtxPMbndEB9LvRFRaEhTUpKWlOY8cjMMWDn+U6vkYFfFx8E0o
eZhreVvFgJSE6grczi+XjFYt0NC8pnipI0B7WeotAOudlR/k/KJYt+A4erLxCtAV
Tc4sZFVO/6c1DKZhskvcn9GozAFpNlhQa9fBlUoI2u1+EgJ1xxwMx116sEwUpLPm
zgOiuF+axkJXVS8WGYGzJfISLGxe6exS8YblRYXeuNV4klBvmB6aFuBbRK066lWe
XjUPRIVSJPcnWm1qSQoO1iFt0SUXJSwjp2I1dCASsnoJQw6dHCyylPkDvfw090Vr
g5KE/hkvbiVR8tLH+7pFiBNxeBWzIfbMOP7pXrHYwy8RthFqfGIz0WnNFkw7yvhp
5obghuGCB7BPDV/nb7zYriY/HfLvAZUTfIwWvqsqqAtZHeoqF+Clw1/MGLB/9yRa
Ooi0k1+WPwYmOpsMKSfpNjT2rHXy3zu/0zmXTLCjmGERQcujLPP/kVyqPMyJXqmm
a2rKHPqOWTozmrpfT2VVwSwSWU36T1FFq1oE7K1eoLXNQb7OKKmOJIG+bJWpOh5K
z8A8xSsYgu8rg4eEyYkYI+ztVJgpdzPbxLhARl8jjLiEE0CyfbWcx7jBEuVciw2u
nW8omhiiub/LQlCGATQzsV4f7TpO4ZE1fjJRo0PHeTNKCg6M3vQWof+a4qiPVKsP
WGjYzoelHAOsbmCFL6wgXtN4kSUP43OOkDf/+DSC2LY8FuMwWzZMjBmtD+IlBGHx
G6ftFeX+2jE2ex6tW0DPBKXjS+vod8vtg8+B3Aa6/et/WTCuNuU/RP65ruQEFPuZ
Dul2aRAtUj5PPou39jgqSahXrP3+vjpB+MWLpfU/43I0KzujNR593EVRQTfPIrTu
XMrEXxPcTT2lUuak+athXDFD233r0k/9efFMLnL4ixTQS4PcA6gVJBm0F9Lt8fw4
nTIfU8+tDwpJbxUKF3/iffjKQ3/vYvwV903NMpVZw9enrOSOKAeAeMM4XPcIbv9X
Rj8/XIkseD0cIPT46EOmtuJC+ioblTMaNWsW/dTzvQu6KxGZAo0yTxVcjYSjUwIs
6KjEDT5EbdhZswqgb0LB6VO5TSxBqQVm05JiiojHaQlKnic/+AimwL29Q/SCWwDr
vfjm+MNSyhWVstaiJ4CdKrD1/bM1sWPDLacoCncO4RWOFuMcd/kmEMIzeGibR+qf
nloyAg40yWkpd3lBMa1SYdqfJvpRUi4YOakX0DutpVrrRNR9PyAQoz0dWmZf+ddT
xlzE1t5OUhNXSPtjqxDx3nuwHsy2WRpN4ux+3ls0Gxu8hn2TrADsOmm50W6C3tDg
PaOGxCUdR+H8YOTagBpqn/joKZZmXJvMdikX0DkKccvNufpwodoZPzK8+LMsQSVj
WWG6/a6FH5QWq48mvcGAaFN28Qwgp23Mv7seWlxeJE9+ttleQL7dho16Fs67eI0+
14e0oYqK9RntRNhxbTT8BeiABb76AWv7rqle2V6jHma5aUs1jrVZbxyWF6HGqXk3
SfX/6/TGZX16c8r4Hlg34Wu/QkjkIlqdSZKWcNYMOTpesy9BuY2YwCO9rxxp8jFB
OCy8mGmCuOLKouvUUx/sNlvc1vLL8Etp2TnO+5CuDMdM+sUfeHRARc78ImJP5ayP
3o/fXKisLXF8UBPl/RIaHzrgl/l0u37OI7TuWl9dJfCTjgiJ5RakhG3GgeuPk3Iz
pTDKj/Me2EXKk+UyTAeT57F/Nw8toNTRs8UhD+1B9fiLB3eku+tpAhiC0CogGWxu
/qn4Qlpc90ACKmULUgeAJMnIieVw+SyGVyY+xHEcxz2Z3LvsAZBEtzEPuGiV9fs1
yQwaqHEKolD4Y07ZTp75NYK+Vd5boeI9l+2sa3hOSCbRv/A++fYLwe0S/V+cA+82
sn54RLmeDMCc6bHOQAF+4kHAeSFobo1vEOKJArxs2WEGOJGr3vC06FXmYtjxtCek
ydsRCGJNLC+jtxJlqU4L9qFKyrQ84l6//At+gexPRsYICIVE9ZloO7ANVOwIP8iF
Ay6wIZW/GRQAAx6gmK0+FeKA258BHZQXUjjBw9HL5eps2xU0UAqNENKhW2cY03H9
WTZ/JAjHh+nbA/ThTmCRIX6KUwSxoOdInsac+xGjMUILMvDT/hhekozNzpiINGAF
8SviWBrZsr+H++jVq9zgMPHRAQtHsJJEh6uuN5hdY43KQZS/B6fzonLPY8UrPBC2
AvzATPzRBgxUlDUl1M8Ui43RsYrwy/JQ+K4/yJ88tbIk3rjHx83TMEoLzDDsmAj7
DKhOsvXdDWBmciq5rGHim3pgv+z7p4YDtHvprpnBYedx9R8sSYLCAZg9pGebvhnj
YqlsHj4782tKSr6+Mu6QaAd+6X8njiRgxJjPQmu3kV0OyDPkE1gWB0iZif/Hiyyt
kF+cWa+u3pouN/L9+skUJakhmB5QLbI1KoXy9aWG9QDLYg3ESo/okoOtb9bkLgeW
ooabmStHBigbtiyQkYExyQrAgB7kODfc7azqqwAoKmjxKbEop/+Itcel4YCuQkGa
pfDMd1sqCxii14WaRbWeD69OA8XByBoyfS3tNr38s7KqbLl2b4uN9eHpWe/1aTBO
s/oggZnEhR/fIbQxNkmpgja7HozEy9vwZaLxDZvXc3AzCmrngxk9Gsg+nxwntRH0
93/HQwhWcMWVyJn337jEQiXYXSjk8faj7nfVaBeXBkvFT4e/NaHIyIgvitlkrJaO
R6ktm/OvFLro2mSdsFAxya4beVijoopSvS7LcNW0hc7aMuRryXCsAB79ei7mMd4O
7pA9nqLLJthQmcyU/EkSXCfnpNScolRHv4oUH0kdOAYhg74LsI5vEAOPu/G65oXm
SiBHYaCeTHs+ih+0ib4qUCNHzLTb3G3OX7Yea/HY6G5y5wgPxiXpBibvdQXZMfXO
YJiFfifhj7xFIKuO9lfmH3CK/gizYYzIe5ury7mp/M3Ahf6ra0FrFrt6RBHE7GQG
OY9l6sU3Y9MYO7poy7SvZHBAZoDJojIYyY3rlMJjapiau9DWFedQ3ONCxATf1MxR
9hdSa1c+uBfg4WipdT/vjaVpQA2LuQDtZkj4zWMXAkxlpSQKZeRttuJGSGpNiAkQ
eBzdlzp8I0CyQVgEF2YWYPttO6IAcowMj7Psnde75wSBrRxxSLfgqnbqwGIY+zSx
XUyO1O9UTWNQEupmj+j68isdBIxkmc56r9eN2mlDc0k28NKGJL1k/NCVS0W2CrnU
72Y532fkhzFPBKoTrh5PPnPx8hB10VSHiq+4LUqxX73LQbf1KG0KZX0SBQI/+4VP
ktrvWSiW1jIOyYCl6/+uS5Xf7H8XRr/n/0sNSS+WNPUmcWO/G35pu8hmYOTX8WJA
GXJ6bTeNNom8Zt/nz1R47CRe6P/UvpU5+i0G5gAX5igNQnYyi/ROT3Jl75yZSjbJ
uRnTuiPgWIaNMes3hWOUpJr+FZ/tFaugFtKDPG0BWA6XVzBmyjHdIbPieMulofKH
pBiuw4ZY+aqiDJwybiw/mBohr7MprXOV0oqWhF7xKSYFApUsJw4Gh2gN0iYrmCko
NUmZALDe8V9qGdvoda/yaRzX0oud5uJ1ergahrDqXFILRgFWdVw/5xsD6nctHrgZ
feAO5Q9hgNnu1uiJ/GPRqrgrEBpnTWMIbnWpjmXuZh8+suQaTFfuL1iRHfBxYdVS
5ZoyG0WX31z1YMgTNQYN4zURKj9c2X07FnAsTJPi+D2jttc/tWJe8erk+nPDVwlg
cwWDgI2JOqoC+vHXWnNL5RJIzbuqAn8C0bjJKTsipY+m4Rf+eRlemqz55jzPKph6
ZPFz3EaQc/ijySQfH024gDsXHEkZSjFACBF2Cdd9W+DTXIrpclSbBOrmMCJbrWC2
OsAhBzSom4mhGPg1HMYiOhrz3RxJ4cgHiWL71S/EhrpSSvWXJriGeT8+jTE493lv
0eEXIaHaotqnpKYxvdFHaCTLT5RPNRKPnUMoLQhKIifcVjh/phox/6UxNf1z73R1
w46jQtcvs00wf6qDPXPbwJ3Q7G3Dusjtg9q7DmyhSTVxG5OJ4fjAwkssno/dL18Q
TPiccBjU/F121z7QYT9yd08T6MO6+Adn/pPrSJ6UEKVdRkb1kjuVI782D+LYn3Bg
0K0O3hah8qwLMnwmOr14uVflpLu9B8G5wrSkxSRNHm2Gh8DoaaV01c4w9CDQefv8
kw1afIp11rpWVKWxLenDw2b0PdRikRRXCwjXIJs/1jF1bquPefX0NUZ5upNdGjon
+lje9XpyAhmXPPYr3KAZhXfLpd4MH+OWrTgjQrGFec6Kdv2fFJYs4DzZ610eikhF
23caipEbLX6lpSi+BFtT3YfqbjRXck+WPVNqe9laIpwz39TjdxE+6BESNy8LWl/9
1DDK29bb4xqmrM8TUc6PQpEJ83suBRCB7dnD4yM7UEJKXttIU5bCOFKSHUAgqlB0
zh6OaDdWi134PsjoCRmnKRfGD4zek9ftyrqf5dCxbvKEseupNgwO8WVfrwt0Hcby
czKKUa9HxnnP8NKvxy5gDFfaJMaNss6YCXty6Xork1U2AqiJkwbxa4YxwmqIWpKb
vH1XM3DGgDfLNCHlo7vJksiq0jwXMJHX8THlVqHOYM99Qmvq2mi0Z7NwwwKOJj/u
InGTbrenquFA4HGX6kALIPD/IYZ6fz2+lu4xHgB3L8VvQ+5inAvA27J/LcFBb8dh
m3QiX4p6btRhi4TjJIkbPJwcbV7TIWk5d9D//wszXm591IUeVslbwib6Mhi0jya7
tofU0uIgTgOkLHJli8wSD34FcDT7V1wlDMl6ZhkCyQEu4TfPBqu8HDz8CHT3cWYY
85cTwDH7bE+RaNASCeUorJz63VuaZ19mLfQ0Wcn/QkIs46ngXP5391FSlubHxLPD
2/DdoQzga6iIhRoddMCMLxnjizsywN6m3B3N0iGmgML3+LzFCmmJaOkXY59nmUEE
MC5wRVT2xVlIi2HAy3ZVeBEwPP4d7KKl+O/6tT7i/orhKcjyYYmI187EIotMseuM
EH2M9FqOfVJnh5nODsSrOPy/u8Tv74UJT1Zmslkc+PD6M9tTfbtn/eVNTYXBu4xS
YpTqvZaO99KesKRvHGwgpUdno5z60br1Z7ejs9/61Avq6W0UVnybcCUe0mMELH9B
2DcgUrl3HrXMP2fsH9Yjq7anMkPhd3I5h33P17rVm3kd48VByS9mkLYW0eobwgL0
JuT9Eh0enZuPG82tF76jHZ0fbGO2PTf0XBVdmy+7Fdb48sVKRxTYe6t1+gCbCkOa
cb2sCJP3WmiaalkLFZhwynukaK9UyKfSo9tIDQ4dHXi/oivIuRukkcVMmz4++y9o
kW9piSiX8bf9RHjnz3CtjT7G2Qb4Flyx6BxyWL8+PAoilQj1leA5pT5rn998Wlvo
JSVh7EVWJq9Qvj/m9AKgHxt4+QPjAEgtel7dbCTNdAk/VkIo4H7ecm7nBgUjlxy3
+QgIKmaiqtHtL7OKvJIUPmm4AYb5Xyi9MLrn4QckVd10NWU9I61j498yLTdQoFvb
8PIFsQU3cmgOyBbOPnUwPPZjBefo5YVobTbTyH3TaDq2dG+yzkdM4NSW9kozpaav
i6E408eMulBidnCMOAlUsmJYPXD9OwLkb4/cWcfQfrTafYSokNuRVc5+XXV2PmVv
YanrUkuRdTL/jduD5oXlE6EfNmecM6Etd7kdaM6Rj9kD6bI6ctSAnSpbWpLbwlxS
z4jPIVL5qPUYupbF+klsPBA84hZkbenSG/y11Q0Bh7EYltpIeaq8CFtw3+zcmiVv
iFtec4b4d66m1UR1/oKdimUtEv8mpqXz20iNqJRmvI38Xra1CA9wmLwgB3JmOIRc
XqvC1pHd9tK+bZIOEAke37v+f402h/A9ri43cumm+Bztszj+vZ+5SC6itxGVmjgS
LBjuwed03Kjwoh1RlaazSI7Uc3R6dA93ovF6Wfxq8e/15RuaHhTeXXnBBUaRquox
JStdU9bJrNvXbzc57wepQoT/aSDH0wnq0GTWE+3O79yPXFJ1VDuNK+a0JN3yR8p8
dVWre+VQnFB8LvcjVMJ9D03kkRErkjo1RL1fSqshldufMXtvO/e3NM0/giX1rDkN
CuqiwTwG4AdXs5v0V/K6A7Cs62FpqblGje9EPl2AUMazKF0PfflUUM/bi7fK70kp
T0eqclrmvM5p91d8pf6JsmB9crfS+uA6CLnQHlIsTgIcBAojh33GuqhNuXioX689
unenh8KVojiD8RSPWmnEMyL4sIZNl4wEMJSuBnQs5OGOgI6Jrr8VRp3CNg20AWMu
rKlBrZIu/NnrRpqqoBnxiok5Z3ysC6/h4hUU2emxCzCSMeGrbpMAn7MEuqN3YSjo
d18asHaxtMQYaLGu/B+ZGtJ7ru/ApYlLPno8fu1k8eHfDU0hE2qQ5erxpqSqHg7Z
fFb8iNycWnJwoXVwBr43VXKVfRQLdjTEgBgDRWGgUUjjevE5QVQ8jsGBy20omI41
szWm2eXYx+KGn5OCtBMu7s2hS/XhVSbioTDGu8GRKe3tgcCiqVuASkkrovVMNkNs
nbHWS2wmsoiHkM9M17TsqAqyllVyN9k3OjbUxjoAuGphNl2rwIZu4lncRCyP5gso
UvcT2EtkL5VFKblnFY5xw3teJXxjP5pII4b6MX3g33nrJa8deHHcGB0ZpSKkjoTu
KL8FdP8IVBbLQ/uiHaeAoEQxZDHaUErYoBQKvRWcigxCcvunMDxd7fhqe1Wo5srm
nURcwNn6qpFJJPmej0QO6DbOil6h7wcpCS/ncwvKBqRFqDf5EBQpsiBp5d6+5yrk
6q+QaDxR1MB4DtpoelwxAU1G3YUKPCEQI+YYawMBb9wdJlx4sRnk9ZEavSMDoj0b
eSXewDkrVsy6U0tnZcPrEj5525xu8xgXGwu2XnfuXurmvEhq16ESrjLYAjo+/2T2
zXhmUdz6OTpfzuYlbCmrjX66Pl6r3TJnpe5uJ+lF1LL0bhUqOX6O++JddkTTDQ5Z
K10Rk80WO6I7uoje9M0Z9gXl5r9r6SnxVXKFP5Bra54Nn7K7EwcyAMJUIFEhPOtP
iCLDEC4Z0ZHq6MH1rF5qEIFnf2Yx+3FEfoQWMr9OcbpaepEkk7t3+UefBo/vznhw
zKT+tsxXSP8lkT/LC4/G1eCmDTeNyD1R7hpHl3xRGwXaTDpCfGr6zNVYNe3J1hbg
/iGp0Fr1qDgGGRjME+x6Q6zySzaAyAsdLk58Dm2zczRNq6kXET55xCHNCqQtkNmy
N6uQf6YyVQMQ4/GZS8wbi7zP9jWRsK/bShosTLQIrOauJEUFBT1T2lTmuerpUmL8
ImBiDXOR+of8oezdw5aemC3AUohFGCsRPsTLRwzFUtQYbJ8M4FpJjK8Vgns4s/FL
EgV2+0QWdOsYnDvZ8hxtvyehoo3OiNAzTfdcK+5JpY2Pp05lBySVRw9QIuAut60P
h7yQS29YJYZSoSpnRahNaEph+k3OKk/C58RSrkhMHQTDspG5Yf2tMJzwffRmaaVx
0LcNiQ/8LCYRzqQ6f3CY08Ezs6cBDIGlfgMF5AU7HsjRDkYFjGL056R0O97WaoKy
1u0yQ8VjyvFw33QLClSunSaY8xluQpQgvwWALM+bjlpj37E2+Ar/+X2BJBX6pUNF
/JSQE25B6SwsjOztbuHUIODe0cIF1qtKVrjfhZ4pIuaVtoE24HHbUgYvVH/sCjNX
GmqdyCFXPF1FDr7Oig8n7d+NVgCYUQ/VXC697bnRsaIXmL7owVrkhe/tRyU+t8Gt
pmjNK8v3AYKMK7ZvwvQcfD4hlC0qYmvn5+y6eRfyIYTYc1smJoQu+xZBlMFEwtHu
sAHTYwUqGyZL1xQsz1tqnv7GsRfrnvhtGzbgcYePpPrjFhhjzFDECvRQ7ZQn0ZXn
3MOFiR/Wtm2Dagr169AYpCSiLZzS0je7WN+JJ9tgCvKnJ0LINkd6mit6vvZRln4d
w2vzJkxzsa5DQymNnnSJ6iV4KiXnLdMP5aInA24AQ9UAnjpdYyExkcMtnZS7gROY
LqmGBQ3yL3Rd6pE9AKTAVL9qXrw0wDj2yk/UKjerE94WLAkSPAJT/et/DWgd5Dqz
y3VevCgxWuGfDDzwNPZ+wn5uXl7B9DeOkpizkn6fWvBVpGmBUUYuA4Fwhz+N76d9
jzuwEN7PtlXWN16Z7TohAmZR2bgUaDPUmRbR+tXqE7g7drFSp2fuBzSR7U7Zo9BT
wBgFvx3xgf5RhxUVBCc1mTjrrzB2jzhWiJFsuLt5F+IoxxnmrJd0kqZ+GI6vyk+g
QjX6Qkxyz9O2BjrNV5LOn8nUG9tQP2KhT6sWPMiZNTHgP7cd/1INtjA/gK+DH2Zk
MXrepr1QqXBBwhQ3YKHIXV1q/gbJFeRtj2FDZeQmxl3Ha6UfBDCkoc54bRNZXOJL
0Q0mESzd/AZ+czaRDhds2byfa6MpIJsiMfWfyqEUwNvYRehdpBI6e8iNpjFxLsA/
hNGNsomNFyT4pt9A694rZVUUdqdBm7hVgRmcrYJ+xiB/7utRFKRKbKELD3kb/qLm
GFIr0hd4SMzS35TiFa/VrF9qI/5Tig4Gfn2mtvJJyBKAZOkXE9kLhD1g5z0plsla
IQLgTz31N3txoDiyVIIiOyYqFPdpjpq8/5zOmHjtMODoLY5hCjXxQRUcGoEGcv//
++epBoT6qq8R8GrgyfrpcFEXeZhH4qsCNah+wPHooyo/JySokL1ifzuSsDOI/D4T
YFFBmDzn+xZFTfdAJyIR6Ses/d+27yCeyOjvXFGyBe/PjEQYGT4q33OPQLboY6qZ
sCexMg/MhFf+PU53U7Cyqitq3aWy3FCotWymXEkGYZFitpiY02/wwcQ518SlN6/Y
qXHzAhBTkOzctGhMR5alccBu/GnnqmbPsMHQDZTaj/VGVKsoO7eyft2hkFFv7M57
iiY+kW5BchlvB8rJKVpnB9Zjwf3LD+J3nt0YmmqgNVYm5WqrPbN/L3afNn2fmKjk
H6xxGzAV4k7dKLwNH7teoaVOSRlYb9vyHF7Y4de/kXpQtIEGArx3msanRX925L5z
lW/JcxNZOmMyCI6oCdV82+plSOskAuwr3z2pG2mPD6dWTCy4ugH8M+sZrQ21Pm28
8JUMMkQ9Og3k0Ejf4dEHC3ppZmOqv6BrC4JtMTjS9UmB1loVMbzGQW/wGhXJVp3i
7fhZVTu78p4Gm3dyqEWNgbParByuSxucE+P5xrZDW0wx6orpoXniV728PQfmh23n
EtW7gks6eHcORHk0CSLwwbrjWaGptyTM0Q4WZqxO+ALOjQMj9YajBJ72+T9bj81e
7FwvRpxq4anLYG4pwvzyhCpiQH2HE80/6Ah9K1JsnFH1E+cyBKSXu/V4cxIVvQax
lEAQkOwoeIiZWANf9QuZBi2mrRT4dXoY4lFk+2k+GhCI+JVEXFLLMdvvyFtCOE9F
kRj51jEegeDqq9NPw+nQItS8zakt4EWerNqP6famnwgcYKOmWuCqmCd+Vz9I+sFd
YCKNSEqVuhFFVrvC8fFII25vyz/2bbmR2unbbAt8djGuiCSU/EHy0LJpZqUJya1c
qpuxAS36HQU47n6dkLzl9a15V5Ju6X8qAJnY7DXn/yOgmP0xMmHtU9MJ9nalj3D2
rfvWhYu7hgDNEWIvdyE340+SkO6mGBvK5P81wRH2usKTwAJwF5LhKaq6h9tORpD3
Utj7L93vAfVT7uuC2a2mlDTFNUy1xxDx222Mq+5AP7CCKFbHO5yFkfgvctx9AzyF
o86/eAS//VELqwJc1JWDF4//UFbI9io1c68KZZhDkcuHPeYvea6LfW5DGj17gXlw
biKM35QFU3rRgtMUOY9K4LsVmhUlS9XwSoYD4rJTQzOkiPU8wWwpyV4JcnYzqg+p
NTG1RuvgUMhmMbLeyycZgVcpQJ1El68RDC8CwPbQIQtlr4uLDAEleVQXsFEoYzh2
s2yOmqLZyhWXKJyyC8tS4CcYgJBlx+pNNEtSNI0cKZWi6eJlK8j1yoaTF/cuMCwf
kEu1ZSREVVXwe8Wwo3nsZWGbzE/LYs5X05YZypwavsdBYu7EKFgFTErNK9M0Ufih
VuQbr1gjVqogyvSL7cTBtAKvRC2YWohBe8CzqD0EiK/a/NApUlq3JNxr76u8YLad
YBwBBPCU0JqVThxu49i10TKc50cNrmjGpdhYQpUKyV9ExMQLPjrMZV3AkOJPI/8L
nOWH0h84f9YJiXrl0x37N8CFsJERFbBSrvMotlcmkUc8SNjDd2DagP72a6S875oD
FjoGUs+WcRVdZuyCODaGKOnVMG/HsZ6PIEgIFRQkPkKyZLni3Gwmsrk6m4ktoN0m
vwZLgKzEONzhmsKC6Sgfw87fivfkZh7ARiuzo4mUjYwq+0D0UwpEVj+dQMi0HXOg
/YU0+FBREsai4dTylx/pGY4DpRTbZaONhqy3TnRU/r5a2ZSA1zFwyUALS/VjIg+R
0JFHRLNxRc74CWnHKy7FyE3B3pNCmH6G5ZkOli95+BynddE5T1b2IZoKBIFs0S2u
Je8jYUr2HUEN7dbqOngVfLrSSNRfqxlD9xAA/9bmK/E+tY9IlW51pUlWw0iFCqti
x6++wdSo6Zsg/h6+knMdA33M98v6RT4a8h6ebX4Swqz7GbgYXAY94O0LA6311DZb
WE8uQmo7WQVZRWGyAR16K8794Abn38xz6tusjvk/W9qWtOR2rNFFqjsQsoVP5XR3
6mqLrNWuzRSy3yZoUfPf3szwqHyVeXhtAjjAOKVHCWdQC6xiqyOV6p0D1WV4Yihi
ah5OrvGMRRStr5TRI7opPnjefRLieBrukWoHL+gG+6nEjGs2e3WMvDcAqHcpfUgu
DZEMG/vdDJYhzi0nm0jut7FOnyhYyBPC//uVftddTNmSHlXg8+3eOzoL75R0ORm+
T46xMNckvP7RuOm7fEKeGtAvgt8oFJwP7rSq9n7dRj9ynUSdCJBSzzPneTroJ6ov
lfzo31IVUr2wcDPFC2JxtwI+BhKSxvsD3FnZ58NYuVSvuVmlN86AvM2OaK5+vITX
cQzsV4xW2pj0vVuPXROCslOTkslbs/AnbTXUr1BQQ7dzah6rFPrczSrGkfUVxgVC
OGl+dy7tOmDho2onc4WGjz6SNoe0MEDe+Z7co0Kras/ysvxSOYX7guyOqQVpIxEs
4updu1fzSXWugVjrwFxKWxE+9VNjtCEA57x152CmfCZHW0/Sg7KKPAFgUwC+V/ds
cVLh9g8/wvYZw7Ib4fZAJcJAkGoq5P43KbYP8qbYpLExJ0af0ZuD6O/BzudHUts7
XS81E+qihiOE0lWZvDgoRKgHZKFVx0iCk3L7EY2ARcio5ApJDhH8uBmex6cRvDhQ
FovcwTxI1UD79mIJw4eHENT7XWq+3Bt1nR48GP3rthwK+NVp0hEHQpYoCmCx6y0O
T8bdog3JdlsuUcPhcl5b/0nbn5r+xJZTgAlrrukYE7X27TOHgvqJkBCEcgTwrMKn
dZaHIWXFU2xq9QtU1j3WHgeos7r5UkVOELJVOIDUjNzNI1ELLRDjW8i2R0Sdup3p
9QJEVZCf7JrI6Fd5STbK0Dk3Vbz01VWPG3RZv7lDVgNxX+X7bN0pi2U5K0QTroFo
MxfTrndJVFE5O/vJ+C3qP7AMmXRZ9Ar7JqD8DxGZTOtwQnDMFfp7+TiZ+peBmx2N
YGVrXl65MUq/l3QXd0pA0oXUlBsDg5fu00A0RYK4hvqOwJR+8VPVcVy/hLr7uvK9
jVHdEcAj9YWlNcI1JvWoQY5c1cXdwQKnZmSTkajtHOuErTQkz+PQJ8n8IbQrKI7c
4/Mzi8Y94Ipj3C21u6GAyb2l9BD/2YDILgocJSQpIzMzzVLVvF1dUF9ocShy3KoZ
rLg4IntZGlAyCHrdUiZk5MJ5gyy+xbP+AIPT2HDfmyMExwjXeURZ9oQ2ocqHCK8i
iiXJnfuwbCQotCikfzaqLXGojKWqEgmG8ZiMIGk1b2Rm/15vrb/2HU6LsOH6VYDk
U94qygGcoCBNeeMWDh2+QBdbFY0bcZHYdcsV+qpy1HC1AtjOuzqFEu9Pcf5hbydd
N6sdUTb6G8IK03moq1OWrn474Bm++YOelvt7LpzjP9KnckzXLySbCAbR2kefd66d
dWni6sK4owginvJ/dwi/D1ZDnaoAuwFs34F73EXtkUOj57sNJ8vbYEnfMk0/s1sV
jf36CJS+iTq19BQSX2oJSN2a44Kp9Yp3BdBgh12oTrabKD/eAXnly2L2GfB8zn+z
Qwe3uv27OezcMZkoLSZVeGbyszvg+ldY/jwBS6HjPwzJpOXU14K856m/rLObj3y8
Gc/VsNlSAbeA/IYXnIrWGRxMzU/i/U0Vw6XwbRATF95cuYkIbB5exX8TJT5qiLt3
H95UznbaOiGLaZNTxyJKaYMrhrKQ0oaeiqitK0m7LQjtDWOT4qdz50QI6vVHeE7C
jq73S8HitQafgJHfCn4yALrjIs3rXM5Yg1DBkDwWLb89RWdALAYmJv9qGK+F70Dn
tV5PKwczim9XZBCDEM8fQrnTnmnD0db45XqunAFKabxBUjJ31wit/bNVynqZ8XBa
R9qv3KkfXvM0Zh0ftNPtvYusWzBRkzuiPRKg4jhXue+7Efy6jcvLuZ8n0ZMhXkMH
msI0Dla2bF7AtYjx1Kmi9GRXkS/BuZX8MEQbIrlIIF8DBdZbwh82sXJFWexWhvz8
iRzCF8SQmpZEE5W4KeGlx9HUpx9Pp1FKui46MTsxLZlqAHAW/U8hoZGQc41y2QL/
6PbFbks0j1IiTW8G3JiX+lFI6w0QjCGWfcOQ5PCD3ibgEfpcuIVJv6ZLU7ouzvM4
lGuStQ+TVt7pjkYdNrEeYgJGN6CHgA1xJUkZLGFtg43H6b3TrLs94eSjgNZTsMyW
ibknHpyQC7n1NhCoQBdMf+PU1g/h7wM1aA8jYH6fPnf4qXnYFQlZmz7S6ex7W87d
U+/Ax8Fu5BxmUiF6xYiTYQH+8c2NwblJWYGtkrEeIqCw6Z9r3Tqzki17bxHsgFym
64wZcbL8bHhsOXyqkMzjAVSnV2XI0a9trMn5jTVgpQW4jjWRQJ9v3a66GzKxbv+6
pWpDHxiGMoDb/P2ac90Sz8iiS5ijOspDnFRHd3/L7bzDiDok0FhVgQGJcOrNfkHg
mPvknXtEBrKheRREbmOc6FLchEhxnM4RZrV6lxXtS5RruF7dB6rXE8MyWdehk6Nf
XgHioZQy1kQqnRTqTPs6R8gOn9/mMOPyma8ApbltGhXT59WnOyTsYvE9gI8Kew8J
h76jlvYUsdg9ALPaDVdQFhQmIWACo1dl94d9+Hh+nUO8oXfEcuoWmQtc5n9/g5Wg
T/BpejSRKt/iCiUOkbJdbui93B2MajuAay74dcnwH9c69PseNalfIrHMeXMOjAwl
CFAiUVHBW0PySmhCjBWgIdVc1eFCWMYFTOUeA4pVukFYz9MMrNS8uMBRWBMwhyuZ
Y/WTqbHrBs1ZXXr04dOWxHTtD7iVX2Tdg95agmtZ8RfoRAnR5AulAaDQx5EQbmkk
6SjJPVQZSu0hcVV3YqU06Z4KMcAW2uU10m6iWnsftoJt9UXeZj+W0XC9cNvkPaYR
+rwBXfT8Q2QznCTxfKbHraIleMAFLIzD88YJ6pAkGZjDAVX3N32Ml1rUFQnkK9I1
FU38+cQis2YBHW+zCu14RPHp2ZRe7O1PGuinl3KyClTnE1vEq6UDr5vGAwuOQhPt
oCN4Z/HVOI9f0Pq8PGtT50Fn+YxRld5/4wOgUDaiE5+yDJonqx2rbiLklxRHRbaj
EKhzXVKDAm2Cy9RxOk5VG2hOlAqFGDzelcIuQaUxhGqxgy+zqMbfEVSS+wNg+ZKK
/rf2i58ZBpnTpNFTwg3QueDEyt6rFZVa7l5kBSFhSdFgikANKgifZdwEr47AVhl2
jfVSW8jpwusoQGkCzck5FhTioAcy607n3n/yItLJCaWFdDHxSxRC4V6naJ4gYySA
oBk6B7WsDqMZLt72vbN7i+SHGy96qmdllbifOanl9MarkLkIsSN3ryQvCN0h85C9
M0fh6IMwFDmbNY7G8HGtwsUBhtaP2Sfz9aPWnNIshkvFL/Q9qq+idUtkfluv1heo
5L0k3YoldKUHeYcOFHDiPCqHkn9rfnNgPAntIjSlfV0sk5xa19RiET9cGcDd4dfg
gcMzMdqPXf0GL9egXOzrBRK0hIB+JzelTAOHJHCO2fr84mv588JatRr7ZNQPT4L/
93AM6etVPA+ocVjf2SGctNpb7dn2a34kfvJ7jw7ckCUcwafHRMQsmqKwTTO3ICQQ
UxUBOqly3tOd8MTIHyuawLlsRrzzwv3to3N2K9t9/BRWtkd6rLucWFBvf1L7nZRS
4/W168QV1dypHBiu/vkPYtMl0mMJkgaW6TEGRCwoMDIK6ybljnRs6rHyT7m+SBLX
bUulj4sEHDToWqOm6/6WDnfU4YEO3qG20LttzNuUwwN7RnlA+eMeueqZiLkXpetD
LQd+mL0UOXFLPyZpEuzbzJc7qdCCx647qCG48j8lwnRQovUn00rpobl2pyY0u34S
4eECrPLci4vIZbo9dRfYIbfSr9LBZZY5WLl7Up3xgET61p+ZAopWhltpSKVOP8zg
zga/Hp93dG+CcNOCJLMKqdgCOmymWyuexosef0VgLuztyglTbyIgD0Cy8MkXKGo+
EFvUuRtn2PNN0hqm8BMKfsPb6TL7iYN0R2Oia/9EJJzOsMeG6QwW0pOKE3wZmJOg
ESUqur1U6KBsSGi6e15b0U6aVOfSL8fPZ9rSAfZGouac4QKztOZ1BpvIJ1JeEF4X
+JtmWFdBEDYj2d1fAqjlo/pQPF9sKWCvMym+kbpWN1lksspIhqsqPQ36zWZ+HeyS
BspLnnA59KE+nJKkFODHH/nUDAJ+WpmXCBkdEqxFA8uEZFLDWcALD2fGU77ak82O
bEbLVnMGpLBN3/AUo+OKY0N05OuBP9GalHXBawFeqVR/QLikB6wen1iUpbnI7wXR
PGIIsVkmbWH3UFFI8Ofao711PhjWjzjWywXy9bm8d4iU2v2DCXUztoRgmyikTAbT
GmTROEZo8l35VOqVqPfLBcVr7wttiSQIRIoD4xAnLQOei0mwk1/gi+BecSMjtwFD
3yUiQI1cA21iicLdfOEnVl4DD3yFK2JhxWRAHwkeiLj/qIKVaHVfC+H9vM9l+j3X
OtxN7916cy5/6e08UJaA8pbtxycu8OIejrPMj6Y9jvZN3b1IiaYGhCmEl8meulU2
ErJj2JCb+fG2rsdyIIfvcfU2UguHpgw/khifqE8MTP1qYFM01841gL/Wv06jBsh6
TEGeO00qFPChO+X7pjwn+2I2hfvbRcJQVQqxZcxTIr2J85B8vRFyQpqli6XZcaD0
JEFf/MzZGvIpCaxo/GMavTiCYVhEXAkscN2vuapNKmYs5WbjZJygkKVE5Yzij74L
l7Om7/HcL7MqvBtF8Q4RCzXHZrNsxGNCqfA3l/mjcmjozYEVo/tuBK42SplJnVv2
Du8/8ppqM8is+wT7vsw8SFNYaUhIHe9X7Vd0YZL0966HbhI+Bh0B0PMp27C4CWfT
p5i2XnnUlAzz+zyUhg31v6QtoHh0DRLPxexC5k3F15HhQL8cr8O7qUkJAGesRG9V
FXLfHKMpnm9TmE4gKkVSY/PwiMlM/Hx6QtRmxlW+3ckkTsMq+3kaiMsZFjMqzbzj
8TaAVjCqagoOz9C0Iokn0OuLm9yrIhd1ceLicZ5MB3tGVN2iQ77xk/2wZuZft5Tt
ZhneySqstxAQi4mqH9b3Pxw3NaDzTzj5QVJMduFF/o7w5Vn+hY4HgsxCTUhl6tRo
QHWskQe345hknqSMO8oHckAhsEX2KvfAyMCQs2gdIhe6wjFbOrhBPsK/6+iebuHW
nPpOjUWpUFl+p2b+5zqZqfhgAiYU7Eq4cyY9emKbOy7A+l4kBiVC3lPOVYtI26na
F6j2WujQF3I3zsHlD6lhGRFSzmsMlif8bh/pKJ/q6AXwRnsAMqFuMCcRUxPlGwTN
CFa97p9GKwqlfmTasQwkCtgMeCSKJ1DXJCoRyrt49niELZii9u0c72ylF4nRdgsW
NoBKCxrMt79NETkNqZHVNofab9D9dvZYtQVZio/QgiY/r6ENSZshtkqm1+JJcwRC
hBMN/1BcW1sBAiPfsPFP3gMZHMok+lDSBCo0bW4N68kyF8+h2V4KRMnOdTx6W5U4
zKOyBq8LitDyn9JUaWqH8XSV9aiva9XZf/vYN6WQ+wMR56CFb7rngas9kdPTXvLK
JNgm1Zds1AuxXfthFGwkwCNLWOoiv589R1OTSmw65Y34Nec9xjhbHk2lw6tm2rPR
DoqkwAaFRPSJG20qBG5HTwNxsoLGjT09YE3oDQ0dDt91A8TJccKWUac0vo5VKHIM
+vVokSch77z8t5mMm65UC1nzc8Hmd/vyMbzDks5fcbP67+pBPLqWq0Cm10ALWKjX
r/N/DfCzHjbKNLv/0ccz7YoEDRA3WzWTZt4S/TMQaaMGqlHbkdEjsFqeYIjZUax4
+acbHUqatWGyrkeQvvEQprO8QpNpAirrUxUg8Z7W8xFsC/UMXGddCJcmgBa3TE64
+K7y7dF3wobF8EqznIoxYjSMHR71begJW6IOE4mlcAD8WYO38MOfScWGx4QiRqpA
JEZ6jtjjvtbyTsOk8XJvQs1CoF9ASihPxBixKDD6CmNxYZ8B8Rx11KEZsTjr/K4h
gTByXNLCXyuxyyfqET/dPtUl0WvDZ/6ROFiav59ry3uwAqSb1Cc+7dWLgSc2UFdb
k618XvE3pGj8LVls/Hegj6I7HZQbCbIK73LgfpPCyu6BgtWLqAnMnG2+xiSJhqb8
tmVVUeLBlC9wA9Et+MnbDeFNd1xiM9QINwXQ5vRRVOjEpgbY01rJBUlIP6eqlfBu
b1dCLr40H03+xBvKJJLcXx5hFA7VlWFCvs6QCuXaS+nqLyO9ANFBaix1FdC5+PZc
kFhNogYx6ppHs06Yrob1BWjBVVWntpJ5eoWBM0lWeopPLmpDuifkcRPYMgzNYwKK
4Zjhu3AJT1wz/h3aWrzCps7ua5SyxBHkoHFtxUFC0wGTgFdZpNpNs0a7clyATugy
lujoZlMTZo1pMsnG7SiMzPTNv8+4etsEYFFX6BjXuGNpaNvyin1wt/T9PFFLOjSi
KUZA/Y/Xqh2tKA6N0+Tf6CiyHho1sbaKL34L27HjfmSKDdyGUEhyDz5onTjHUtay
KBfhEP5MrpuZvMKL4sRukV5kJMakoNxOav7Yn4QN+NH8HHjh3URvDYrAxxDRFP//
j1DxrRB/h3Lyz8z6/w6cyn5uneLVXb1/HyAPXk65RzxR8k42rO975TMvN9KkbaXH
51YMCQAcZO+ob3FnfVAYOFLNkiMYHZKO/V3F0WBIXB3VfzT7+RM99DgyqCYj99hK
6rVfj0ykbLhMgWSfGOB+yqlHzN+NnmDX3ISOIZh64kJ4EV9DV5/kB5YMxJ8ZkCH/
T2cW2SDZQ8/cdO29UP7edRCFznFNVcq0nFPD465ezz8frkwJLONIiiHWQiXNszqP
cAlEo7kUBUicA6C7jGjCbO1W94+o/eD0jvsuxxSh04nNjPLvjfWtADvxOcl9fUX2
CWpnBe6e9woEopYo5mgomLdaMxsKoIVoTGxSPOgRfbuA8A5+m0sUGBeOmTlvfcWC
BvPtMt4LnTTnkWSIjjhrX4WZTCtBsaGLDFmLGzu0iUPhcwj8dyU8uVNRFrfwYqDn
vmTw625unmCj29wAGpoqccBY/iNwotvuL7jRKOsTJVsxrftFlD/2vYPi9VyCS7V8
wpeEuT+rPwTz6YLrE4Bd5XnJg0eDFmJUT9T1TUp2GFLv9J3z9O206poHHByUQhee
x0R210y8hamAcHf1EsM6aUleDeUMfoKnRzkgueIWcx/C/ewvfEUz7eL7LXtb2Ytv
bHzz4M+HM6Lf2ebLGmuFBt8pi5YuCwP7wuWGwfQBwIU1LZjfS7iM3hsHhboLeR51
zLo4QqlwseRQzAuQbu1TENcvqmMYjkpv0wGaZHw4sHlgannWJ/+cdyFCNNr8bG1R
LI9j1sOhZ/G1lK1YR09rsOAoy9x9w87/Qv/34meBQBtSua5wZIIWm6NVHZNw3H8Z
uDOEqr69AMZtOJycxlh7X86JppYzpnAiPuoqYN+RfZFi6AEZA2lUclDxbJF63gBe
0bxNumRLqUCFAwWrxsVo8oltgqpqNNYqgTTjZ/WDI5gftx6mOL3jjwYx2v9ZLZXm
QAxuSGicBhPG0X2L94OxADytXjkLzvaNV4LCcB44qtwwI+vvaiOvK7pjt2HIfAU8
xfCBdzXPYUBpZYVsEzajS3wEg9SSa/0s7X73ZyOkNfRiSyUviRWP7Vzbjs8KgQZ4
wsgdo9627JBha/tmhUP5u3/ZRPbVBKuzqP7lotwu1pF4AzdGb5SgzUGYxIO1amMo
YANHAplyfdiYffbqf3zPIKzEO3qTyqPK8OXrhj2T3zgEBURG8IVOZv9vzHVQcXsQ
nBrCCfGj1H8b9UWzvPqcCSIMgErGreO0NdIyf8oIySafL9qdEwwclwM7QvtiyuSI
0YbtKekYcA//prSGbeP8zZ7MwCSpSJ9WvWQu2TCKNaW+OhVdKRUudSHbmbmjglcB
Z4wFpTvoL10lZqUc2G78JgCvOWqW7/Nocdihac12mxetuohQpW4oDpTPGYKfRdag
+75NFeigBbEMQlCmXOsCJ5xa8pMOtSN4IKiVc5Y+7JzLncwo0fJZBJ5MyhAhVHMM
4JV133W6QTBPI6fu0B38GqLCMb9zLtd7j3wpxe3O4JIOxVhJnU9X0WeyB3eUJHr9
eUAqC6h8PH7ywFZfrgSlKTpIreUsH0ZffD0VJccoHmGDIxd7SNrdFA8O+lSTKALe
/stoWHvE2ZAhtE6zUfWsG9fELUGpJStzw4eiciODbdUaJidQXo8m4oxZAU2txc3H
VG46DR2ondd8VAh4xpKQmV2dlLIDesVkuHHuzh/C7+FIwhKZM50ip/i7ymT3eedz
AbLTA4Ek+zk+0Ybrdn9aHMjmmVOUqGPDHYOKpVbKscm2b7SSIHrQ/RANafc8DsfG
po3aDGvoJmbI6dyuYSLN2dgBXXaCz9laSTdeR8jaBGIPO8VoNuatASL/0qVqlybk
pc3tsq2CIVFph8wXtxCH2LtfEuEXgUS3scSS38zXgEZx7GUyvSV8VGEF+4HIgRij
fZZXXJJe22GD8OLvZr2tPL1/TbDmdlhHgrc7NOAFniZCff/s/IFglkiGIUix6o6t
3pRhvy9V42mZc7qd/RwGtqlQoV4rjvnEFOYYEwkpuv3jMGUwMtQfEzOB8qOetdY6
F8wOZsNu5167IbEQMfGrE7ZeiATUjwcvkOEWp7+otNOBKSRdTpURfv7ZxxEgL5q2
MzZB008bom0B2AlB8EL4vwVnlxQ5uA8N+DboEmMgd7FGzluKRtQXxZKBLPuG7SYA
nSQg+GkyPZJBmGYPZ36kFD9xDndebwBhfTm3u9y8eIqZVy0TZyiN+qhEpO5Bs6Hv
vF1TA/P0kukd0sv9gxz0oUBv/474qZRib9QwELvd+DtF+a3ZjUAfBvuTLdF5sOhK
vwBNos2S3uFbgwXRtjTXS/duRxJxccIQ+svEI3fqiN/7C+48UVufHOJSHeOinLXY
DL/ghEY+HjiNGAELkzCY/ngKbwKnczHoWR6f352PtxlMi93XxlHxldSsLNI+VHzt
anQXO6UDpMBQ2HKm4p6LX5YyTGSP9KUYYGrfuv8afwBUf+MvEcQvoBVzdJJAPuLe
PVfG8A0I3HZqI0TOL1ka75MrbhdlOVWuauTR+rjRx41AIrn/wuqAhofx1gy2fQ+w
R4Wtgj/RFC9EdHt29Nvn88u/qVbi/ZkTDv70pL1ZZPTxWWUy908QoABV4zHNauOu
32wvp+6VHvv4f/4I7DX1cAzyeLELFavLMPhoQbB6V1gfIJuU61MwHjRtn4fCHChj
UJm8bnOD8+6lTcAuPpCFq6/e8kSAHA068O+05I8wvIq72uwNneQF+/eIVfZPkL8X
3T4Im+hZGP179fWcFuQxDkBZy01zoclojNgdxWdH0HXkk88f/D1SVqGuppEsGVUd
0U7jBuNOkBKra2fRNd27lNb9AsVC2zkzVELXVP06j8S58/qg9wo13fkDVeCK+ItO
Hu3Uv0Ki02Mj8hfpBGNxg68pPnvNtygNY18zooRDsoOrdIXb/W801JnTTzEt9EDY
PHYxyil6wYO00kaMmgIp2nEfUdN6k2rQ15Znjmz/OAKwxKkDtrhzv4S0WSF8s5s3
+/FuYtKJiy0XwdHVKbCgUuxUnWDXs4uIkLI8SzVuBT4a1kwYCqJZF880nJEJltSw
pr3h0/d2I8i6yZL5p/UKQKxzm3VC8QoTR3cCyoRrkqI43sLKQayo5fjVZFhIc2u0
u9eDNSNJtWlVz3ofeYhN9+YrSESJiW+rQ7ThCsYP+LJZviKEjggqy0fWrZ6rp49K
2UkFvxG/JhnRCtbFW/M7MvnzQI0MWWxHsi9elct0FLdjjpTJ3mtUD7z0ttkGYwpa
7d3/ibErTDVcKECiNUvoO+9CmuB3I8qq54OD1qYlX0bjMqwUCxstctsq9DuiieBh
sumIpC90KKLyqY/6RoOmjW+WcgG0HBiDXbvKbT4xO/gr1lrlmoZbmNOJh5MAGvvl
zux9S2UBMwcz062NM9ifASaof3IK9PZ3A2J9H4C/cZHqSgDrMEebvFglN0bXIYMW
O4Qqz36PNZHYDWwHhwD60UMuQASP679qyGiv2+a5ixzIRgV3HHk3W4FqBvdqkBhP
SCPIUw1uAbmBeIffw7D5nenOjarVRMGV7Z6eijjmjMVYNV+PnICP1OpfIHaqFwRG
ztUxGilK09bl39Cw69ByD2JIJ64jTeoMudiL1+JWw4s2upvuJCN5vGBgmvShq68w
HHIlBhmHaArjtSNExTfa3c9GYV1oIndALti/PYcicTifNaRBodMk720PHJNRFL0o
kr+PyMaiK70dPcWwbt7sz4euRtNDntfSO4cK94UrzVlJa9FijJ7esI0YZN0CiM4F
geAZHaWHqgp6g3qVfPW4Z1AS9YWYQv6ZIjPcvJqDxTol7V5A3ny6VF0phTzsvL0I
lHfuTfRZ8AbAoDRmJWf5j4gBZvlswkL3dVt/jmD22+r+TfuEvNTaALOodN/TFU3g
eI2PkUl6RGjl67Flzflb+9vC6deon1od4phQizPUNqxDdSqps9o2ur6IezL43TmM
yIffEy+8tubj+YOOuV9FS5/stsiAWTIiAAMOXCnGDAK6cRCcqe1/h0MDo6vb5ekb
lCkcwjg85TifrkaG0k2cII9elzPAjW2EeW7g8kaUVAgdQDms7H0JqyBijZ7tCxz4
20sefYXrHxNjuHjq67RlWN33vbbryU2fIxBeRBbNNx1HfvJ4n90cP+O8IH+yj+cu
G4UNjQFpAYcFaA50Hd0WanBMqmkCBK06D1iVHnOtMttN2thspnjCEa4ghUyUEMY/
ZbZ1G8jgnwg8mUxl2XlGGnxuPyN5zkONLh+aCdroq2y4poXnC06bNjxVIl8BRI1a
19wB+1PPIGnphQJVAncnIx13SlAY1YhN8xrgC72ftNocwpceF1VCVHLcC5m4uDWY
rMkm97g5npJ7cdqtwKE1/IFFtqfyPFCmAYmXZQTfVedTF4GchSrQnFmuLWOkZOGS
LpLZQtNQ1JGJYZKPOpGxUFI0mwKiWqU4/aqGdmxhIm600BojIUyFtn7GW0tuqQyl
eYCQsC10/QJVtPLM42B+QhlsLTWTImSyILV8cK0Dv9hbPBPPaT+/PZnmYSC0U9ym
SPjDuKc3iX12M/dEgjVQEb3volQQ0FhXjuuq5BROwPX+LswFahj6/eSGdSobtgIl
YFswA6ywHCUeEaS5e0J09JsBA06bHYcEbEsOYUY1dT3Oy6aLxiUTcBEOJakJLTnb
LwxA2Pc4N2BrGrxB2z7pM+I819M5PNGk7Rta0SKIANflVHkFP8X931c5AJAcjiFv
pLlOEYVgE46YizQ1FxmWKZYfuqdbC4DKWtufj0/ugJl2zSFVXUNMEtfAItbdmCdl
/nx5+Zd7oNf+fs3L7lh8kPLlhoawDl6zVUYxlpmL8t7y+jDpzS5TcT56AbSPFnwi
he/DeTIM5ScUmFUyvNHMEUdOhYTY3/7PpvaGLsSqyTkSuuLpzR/UXn3MfV2HV5c0
qfrmJQQVmfh30PpusdFloFGeKT9VOaSIE8dbiPPziznaQ+soi74T626TSYXsbFK3
pCa0DmCD1eARPyd9c0k4wnPOsY7/vsGUt1Y6maaRHdrhgdRlLEP8kkgSqwJz7tGl
3vrgqpRln9J2LNvlIcbzonevLeMqiR5lHR0umLSdhLhYUQw/vB0hBmyagMlOMjP/
jSswqCiiW/eQahcOF6K9xgKzxmUJG6RHO4C7lYt2+PzxK9x07WReYlKCdGB/kBxg
SRP6wXHJy/4n8uhfVO9LH+5QoYRpoXFxze22MEXhIts/WSh52emvbbyoBNSjMmcn
fXZ1gaNHe3c9qeeDck4cy6jldLsFIBzzipQRb03qe6E1LGP3rEEStAlfb3ZbRJIe
bXpNDW7252KWsTtLqUhfB8iOZLmXv/qP/sXPXf265JJcfcVrROvSOZkbd9X58y8K
Na6h7220QJ1AgsqGCSPo7K8rF0OfwEjdbaN0Sq2cjhO3dGRXsJFR6Z1ZZD/YM1lX
hqwFnhKH0OCimp8UWQq8chra+0dfRtDln67aZDdsWwFlvGzHrEy3+IGeOoU0QLKN
8/FreFfdvNdlKm1WLfcims0wFxi8tqidA+9wwnPCkdNoJFvZU9hWWX9kt06NK+l+
VAjRHHYgEPVigXQTzv/TZzZvkhsdJc9KGcwlpxnEOfENa3nThDwE3JPGJVQAQjoy
7Mf9X81aZECiFfoFFutV2ghJFqoF4CZT8bseLvI6uzxla1rnm8HmAe892LEeBFc4
BzYVPXSoJzv/YnI9OlKmBsIvjXE83CBygA/ol4vRDT4iL266fw9SNlpnLE+a+KKS
88uN0JRoqf99AGj5MJ9Dnwfk7XPQV71l7VhomgxnhnEgWH6Uj60od/uu4D6TIIe1
wqlMKkWauTSVD67We+vovbpCwyhMkCgANsR1Ra3ABCecbCwKyxgZJB6nHBQ/yxhe
Pkc0KuWmw7UKkllaxd6Wmm4KTAG+7wt5CjLh0LR6yXOnhzNclAZzMkEDEjEGDOEB
V138z9YSzg1K9JiohE9uxQf1QQjU9BdtviL2S5V85+jVG61k28jHPWa7vBm4MCIf
DxWi+yjk3XewE/7WRDpLAhH/Sd1EyL/XdnDqB5mnkdU4QAcTqq10rxHV6eAGhIb6
1i6I7MsvJ9ErsRIJJJl4YAurf+KgBWuoSxeOyNmzu1J31k0Cg3CEuikQL/1Kvrgd
L6/fzsX5f/4hiJZum4An0uZlLSjipdhp0oljO64crztTXgK6uFe54/EZx2KRblu3
i0Z50jS2HTt6nHHlRZrT07dO54yQO6EC7yXB4PFzE6TSNhNb+JXJTIHIdF/7PnzQ
e3mDSNubr+IfRh97Zfp8v1IEA6hWLJwvkdqQV8kYsTjGg8Kfmbych7WgpbTmBGYT
iFAbnylSVOQuMj1QgHJ9Iksj2s8RGC4hVYmpAWh4vbX1e64C2fk6senmN8oirKhZ
HMVSF132LaM6CnJLpUpiZGTOgx8CawopLmjMcY3xVpZivL8/1d4gJ5dqvSAxjSRu
cT8HGuxg57W9WdDDiqOmP3mla7MqPbW6IuB5QDF996N3f7S/PT86BIPzo+VWplar
01Zs+mYhSP4KTJmehHP+wUB6TRp+VkuBcp3t6k97nBiYm21h6uPsOXOzs2nNbgj8
dtFa2VyhdEqmHpJbPnzmQBGjWlF6nivLY/NdCS5Mj+ZEF5/n0kYhi1fEfjNmnrRo
xsXZbjdYwvXZf6W+BKe0MqHavx+vY+hSnAB2zr2tI/MgwRL8e2J1qgBW1UfM+jus
634OOhrKd+MhaoXHnv1CfP9JPD27fsIEKdzu+yDa1mWt8sbzBK7PDDd+l/Fo2NG6
YvXdtxVnHK9yA1Eh5DFdD4TX9X6VaHj1i+XyB1h59YJKIGVHgSckVA8itr9raCCG
0w1z3ORLqvbfR7Pl/krVwfXZnPoK2CoWWfT/07Hyf8wLOJj3Y6fLhJ+7BzqaG/VV
S/CSci7AkNOOPaTCqum7I7mfwNx0PAgjUqNNu82vE0ICJaRWmO1el8C/siPFqNij
u9ov6vXydT8DA3bFKBuzaUzRmpdFf3/MCiXj+BKDRsmQmtLG8pTyDm/Q0kEywtWF
NjgQcf34h4+ElPG6uC0l/1ESBbk5E2HX4s76jH32Wlw/KhnTctuu1RokidmSAo1n
ZWeNa6jZfePM618yDrzLCbihxeEW4571bIFLwn1DWA+/YVMbctuBlsGwozbeIepr
l04OaWiyfyB74WNSjcn7N9Jk0+NkNYI/veIhf+cegV/uu9LVWu4ASTE3ZN7hHKJy
QiunF1y9YeDOBR8ssNAeMdr18bzmxpK1nAJoUblVxXva6CE4D4eLQGVNfJfJLinN
am8iA1PMw0NRvbhlho+T2jcYuy5ityI1G9gbDHHzyRzR6pqLdK336pajYKF24uV3
l4Y86h1XPMLtxqi7qWVhPfgPne/ztiU+5jG/ThE2tyS8rWWIOEhdo7uzMX2kaL59
6ZxnJEoUyLO9e79S00gIUcTwHR4IDWX3TPFP9vKC5/90St9+OmtYrM7Ow+BpybdZ
ixMBysJp6a3aKLoZdCLMtxibSc6gowvgF0/rxBbqIFGl+DsuZ+0C+MTue1vD4JLk
E1MXW5Zirlk5PzgDGZuzlFC+isGlepFYptq1NKalz6DFLuLA3ERwvyXU8HVaSNd6
oh3vw6AmrPGqHI1hOz6ANtUGmuoTtOSxIpcjvh41tftCFCm3TH6sQ3HyT8CboXjV
BbNfKn4cRh67NMGZnVjC3GSk3qIifXvi3pXiOR0C7mXMakV7HKoioKhPBV6CCShC
ej1bGDb5D9HDHdNozRctSNky5IbRqsC/eEbQIXP5sxBpAUCfSNwiRGxA6taJFYCN
PqUmOYwce3kgujKjDRL1uC40IFr4CtRvqSulcMOXRgoofxnF2PCAnHl5ho22IhyM
EROmLDb6kal2//sYpctFRRGF8g3fAXLoOqoDoTAu/39tu0eAdkh0x/meLfbGXlqZ
3reBWThdQmVnRZA+tXv1rCxc1RAg2y8GXjxhtki1bvpVDr0/iAuag1Gi7UYGoJ5z
A3gaCSsN5fHnSjy+hgzF1ZmUs9p72UTcWeZf/mvBVjTtsXNB2l6VaceK1x4It9d2
gYm9lLZB+TKRrvbAjNsdqMka5+gcStwe1h0yjc1UC2pb2u3CYk6zjqgLViSQ+ER6
jpKjW4UhOtUnKl7e2QIb5VlAyw8juiqGuf5PGOvNpFidOgVKXno1nDM9ldPUspsp
gosku9O13ZFVs0/nGkBN1Ae4OtCgFoktc1kk7P5NC/f3/kmeMNB6N7RnSe0Obj/V
7CcdtHugFPuQceSnrAgPm3yMC1D6Ky8i/9FJoIfpCzOLuBCXwyEBgffNZZAYV1RO
Px/5+sAxR/iaFW5jrhTcugCS/bnebolosTLBSsykSQHNps6F4IFVleANCffMjtju
RvOfDKLyWiz+cpCvFqSSFfgTKmKs5MfqxQUzXtHT8ifsoE04wrDR+J0H0lyZvD0t
/bceVuP5Yc81r3i9Xl4oyhexBknD5J3z01jwVC2A21JHgMbrRM3XxPpUZ2s+6o4F
TwOWCD6FHr/ZUmoLkO2+rM/TmD+U0fW5w+LRCbuRyeRMEDtS+LixGyrBZhUZrBrm
7PB0DfrHycQzZSfVD1QwVA8G9+glbijVWRuRi/J6bdirAhHQCQ0kCtLELGI7BrZc
EIYo2CTyVYtxJULq44Eu9obx33r+nJ1Jc8aatepk4nBsw3Gjxjc70woWQQF3ZxPF
ylgboLhGACUfbMXYkNRlDQrt41vPY9PnlEdqvDRYjwUPTl6+fFj0C4PZtKVEeMmU
fs+Fe/IcpDG+TuJg/kAJylXt0+5Sr9JxMLSleXKzK/F1Na4ToUdVy4uzEhKIRUuz
BrebyE8LjwhsfTR/5XXU4RGZE8n+6i7a4HJkkpGEZmdWYf4WHWe821nliswvn2HK
uBoHO5VX46s9Yb4kTomNF83wGAb53AoxCw1wNEkAcmbyf9zU1dP9EELcdZBW+WXQ
bCtSPYbMr8K3E+i3FKYcPldLOd7bYZHa6bMvHVT7DqFzv5UuPoiQCiDDFAVGvWYD
QcKccTVHGRWnjK4UmSv3pqry24l8w1NzzEku0r5PWutbeVEliWA4dUClkUFJKVuw
iqdzb8SeAJK01+5hX5IB+PZ3jQK2UXIfQ85RbuBW80bQH43XLIVC8IZgRSKS2hwB
5wTatU351HX6azWg3c6fC5PTcaxtUjmoNWsVvU+/D5O1Rs2wpIpGxZeStaV/x7DG
KOwcgwKQVcumjsZ0J8G16rUPKM4RsiEE/1UPx3sG3lEfWEbL8zJMaH8UI8uVIPrf
O6Eq1BCMgBv8xF6eqzzSyhb6K8Yg+ixWVajT3lBWkEELJB8EItnOqlsnv/6sKxY1
R4GrdXHq9AOHRfD1XOp3BI+kJTPErq8Oc5JRWetv2KNNOVbI+XmmDcR8gtTKQTdh
x87tQB7nMPdOHzj+eo+dwQ6Yd0K1qnEsR9cKRHg07JVhC47GSEbCm3OoLCQfgzEn
XAbh8VMZb9HhLSu+vvY3ij8dSaETqExMjTtvF5cpNIFqijg4vFq2X283A0Bn8zPG
D+QvbfMzPFJAPiIdMs6UYC0gI7kUPWZmxqt8xFAg6QXxrCl8fqu6Tt77KlP1fGmZ
n8+A21h1mk52X//XPiI54aqCKtyh+JfP6lo9p/2l+seLktWYs5ULy7GjHhRrH/Ww
EZsWQlyQxIvCKW/oGtMNUqDkMLtOsHRwn0Q7hQux9d0ANjwrWciWBD1Ulaum4YQH
mq36lzdVoIRdae+7QERoAcNiZTuFaSKF4jwHWM46Ic9UcG7jHWuOM28MHL2s9OWu
+M5qfEFB8XOJLukqdz8XvmEfQi2V4iLfX+mMfP038V8udb0uY/oyQocggVnXcE9J
XmS8ENpha5qh/j9lxkCHHBAniXJMf/eS/3yZJAMpbBRz7SCGOD0ICdgxtd+91CiY
lAB84tivoMM2dvGgyzxaHpWGz4vSTbxJJuJSU2xM0isl3KOIaSTbvs8FmFNfotmr
eSE+cHpmzfVlycgP3dfqJCmPkxUkmR+NYO3VO4Qi0NcQ3R7iIiSCbmFh4+FlAMz2
mTtS5PvNx81JkzGisC86uUo09+fiVxdAW6HjgNRSTEoODGGZ91LMgaMBulq1lYc/
5K+uY77rzLe6XaYRsbFhkxhLUgoZtMJAilZHAPtc8Jd+V1ZBaR6WR18c4SpkaVRj
N/t6dBc+HDwxD39gD4lh+xO19UpCUXZnFxoP/kFqYfc3XsXmB1xpQxCnFKu6Mp2z
buCPr/FpuQoOyWTIBxfOqNRrme5STRBoJfKh2QHvibccEQ+CGOpZlPjAP+luEruA
6Rx9QZPAX3BPzbQ8WELmUP1KdV55xoixG2iLmepq39P1MSUOaZNPPMy40YBcUq/9
it/7e+Erh4RLaHBOVv4broCwMjHrzzhCk/Rm2x61Uu5jFHsd3MTEKW08GW0Y5/7P
dbT04MT61dFJpQiFBF9o2s6xRLrhzB9Ytarys/eEX+zA0uZWqid02k4bXGuHYcn0
D+nAHqERRLsE5RB+Gi4PiAzNKm5GSCopSGT/YztKzXkG+6LtBaRedP1rzMLN7Hvd
srl88cG3owpUbqv4tflV64N6igPDgd+40XcyR1wJnUEWQ0tXui/r6JgVy2OCQQ+g
7rGYl37dAJXJVX1GZwFuioYdl6kGXpaBdfGLsRex4AvBrTackmXRaCpYzo7bZnPN
+GmUeKLHjUip43/oYNsWSiWo6xnr9g1VlMJNDneR2QEsgEfGYtWzBCYt4wuntvUB
ywC5T4tddoc1E97yy91bX1KG66OO/LrztUycu+yfRhIPuc+E9Q/0WlcuYC11MSIO
fuP3Fmpv/qkt5KaV6XeKCIeit+HrQO4NAD8Qg7pUsUXLLwuiaVfoAlrxVNVSOmvW
Okv9dDkp/flIRo5WojDuL/jDGrrb+lD7bRWQIRtlhLW7PC5iwVF41BHMgTJfPaT5
hNrVJyVTh+qrE9n9VpnF3XIHWwjT4xCLm6tldiNYFMiG8cry3lK9XRYq5uIH5qsY
DZZ2ePOq0EE2YH1W+Vd3elVCf66EbCytvXqS7z5o6p2kP6RhveSZ+mDJ/8gps8aC
0GZLTrQggK4fvHLFgqOLaNOFZ9Y4ACcyXEr6NH9W0zHqyLUSjcCKEQfzgT36R6n9
iHDtC00bwwaFdlU5yxIs30yJPXJc1bkLkn7PfGVdHScmc6mC26tGepF12dzyYxpp
GCj1tS5xR3t781Mrd1JH0DW1sOanU5d4uCLsyeTkbbSIXVcgleQQUuT7Sb+ixLHO
JLSdxgL0DRDd6zNlLVGIJ2b2brtAy+eQH4VZgL/ucqiBpaEmhEpjWbfbpLeJLQGK
pI5QbVvz+i+tackDmyRSfYjomqMNkAQ8ULmTDq6Xy4AOUMN6JmekgHY95sbs8nsr
GbwAyE25RPLVsOYw3x19/GA1I8YVEVy6sTMoMMi+yGS+qteg5G4JVAvny+T2Daur
jEfmr3DDPMz8qPmIYr/g5ZVp06Fz69aggzWLU48/2O0TdO5PG4Lj0e56NMoavuLC
ErWh8idpzQMTnYjIuEtlyPJzmv3S0xQ4GPKv12syrmCgMN/gAPegWyUugTIrYSiT
JOlxMw3Ct4eagUYyPDyWtMIAsMhd4z29v0yyii123B0feBD95KPEmHX0qb+VwRe+
s8reyxjOToJFwDNHomGkAst36cF4IWxMnrutVuwgGrjlo2KQJPBPKzZl4ZEBjT8u
KAHd4xnam3CggVF1HAX0vA9L0V2yAIow05TEAGx67yLJeVK6fvvFf/i/4ahQjS/W
5aqlTvWhwMM96o6zPkmuw9BoTfRUDXMRCjVExmTZM0bXbl3H0jIQswKy6kC9tzpH
O+5O1NT2kLj7qBqYyq7uW702IsZMsOgafqT9NtHDHPciwNy5euOtqQQaMCs5PdjF
vo/LneHaQs8Y5P8uUqzSTeVH6nnpvPpqJvFQupkm9GejSthj3k+uRN6OPh6Kv8K9
6zdlBpI01yMwMr9Ez83l3+Or5iu6msY/frwMjinEwgcCNb5kfUqmO4sSVW4xpgsM
EttI9vwS4tkJyy/Nhc28bXCe6reFkXLoAxhx7GcZaxQMksQ3v59+Qb4pWm4gxPZc
NJIijnC79FdCVpGYxkt9JbmneQlbbae6m2gSbQYcoqt3h+K0w0X7Mn7QlENIjDME
9JLxFT6u0ybsjfPRXMs+8iEyf17Edwbl/ZscC65eqYfyEKAmiJbC3aN3248yM3c7
DjN/mcew5DoW3U5n/i0hNnjub3OlHA0PhLmrn1FGMTVnLMTNpEGOF3QEIKtjzRc9
lrtfHR+D67NLhfyKvc/b/AQDx7t3OXytAAP1sWdlrAfX+oVqpe+lt9/qVjwC0iYf
TNTAtMPMsaW8nE40WqV0kCuUcBqc2NOhP9Pg+8ARGd5PVGYGbOYHWxzK0aqnX0F6
KJecYxmr5JTtk3hhdz8w7KIMgECrNUE1zbyeddGuZr7A15WIlWRR5xMRw2F6GR/A
m5JoPRmFdrnl4vvgd33ojvNYi2/l6TkxoyfcIqAlF5mzGPVPO5MobqkcyXCfVI1h
CiZdvs6bPny5PK54VOJNE86es38k9Y3CmAGyFSz5zUw8yxMutdU4ptDSw0jDzA/s
ylraqE9UQKM1A2xJJRujyYsnXd1M0HhjKnXV2zPkkOP2DP/tVsBuMPUa+Xv6fO0l
Ma+kX7cKwNUuyCf7/MhvybX+W53PJXTw8bwcbgdC66DYLALHMzr2q5togMTr30n9
QMYGONlhIV5NUw8kj8wWnAXNrO+3MtG4u0i3rlcvLExbGPTNORFw68cwVoXfUhpG
rVK/MsBymIrMxz4HKOQQTwpmiECBfdPC3CTS9HH4UCXKlwJAyqOmVimwUdASrdud
NDDvazx7uIL41vI2f89QT9qohEQt6sZgtxIBnJAtEdTGVtb0sxPuvWoXmO27+pHL
Mybla5OuMd+x/LAinb+D/RwJZjaNeNluAgMdcJ3Yjssa6D7CRZdMNoN1BiYn41p8
yapmHi7qd9IUWmAqBtKVzDYrkldUXiY7wlhTg6IWlx7yDHkSIZcOlLJ9QJTKjGgo
4yC2jUSSXRf7kToeqOoC4Kvmx5NWFK5kSXGpzOlDNZbSEimFvjU90V82OHibQ6Q2
eVeiK93hhKB0jvgt0aVVaEGo8iHM2RKiCWjEcZz+Z1uCGBZCKlfM0qOq/nv3dad8
O7n+NtNa7bcMdaIG94upX1GoA0qyKsm728DhRHArzXOsURaLmTy4d4WJrFbJy8dh
lfyE847PNXwcFJD6cdMuzZIWM7OpzgMesOgp5Zruo2vyrVwSV3iIO70uJ4N+NwRH
dz2RoU7m8pDUFuBMC/ADB5xunDlP4kDExc0m1hhz79Js5Kl3ZbZ/GtyjYy0LYVuF
qOK7cRaQet7zq/XmUaYQBtPMYYA4WFHfHr863lQwbgnt5neTBMPKRsKdWkgWsKrt
X5CtaD9nrLeKtHFzv9xFXiuohlNI8MVUJkde2w++6xRqoi0i+ZEWrK4E61rSGsZn
ROgbEumJ4CBimyjFb+Isv3KpIf9J1VZetI4ZQrPeJqL8GG0XGsWsyWxFsf47SJYz
TOl48sEoEtuMEP/CrCzh0sABiaEWLBqK6vLOsQX4+wmDduH/1h2jd2lda1Ord7F5
kCIfHUtRG9D+7MWauMvMgiftgy0tCQEKzS15/SAs2pPQK+2VUKacO07vjEBWywyQ
hJCcL6v6SXGaUyDmZSPfPOeiNNFNKPpv7ZI7AtinO9NnXY5f19I+8Ai9swSF++5p
dvU4HIsUizAr+eANy9ElyvwtRLXeIuSt+0xSmK4mqADOsrStGK0vW9UjQjZ8ZCTA
7PT34LGTOR0exMTfwEIztcksuXh2JRKIMifqnMi6mqC5sP0U/yv58q7sfVhkPlgB
tLis0UyAtjUlVug8wCtK7ObCv+L77Tsw99dE7+KC8GSN5n0izcWU0y4FmZ1y20hP
ANqDe9W4G7abQlittxFSc9lrZmgKngILWWbkLJslNuGIdrGkCAE1Cn2SNSm+UWOO
u5UxWMMGAUTqRHMtvIQzYyg/SsFlZSOVi+IFEFuMtdo+UgGTHYGVigB7x62dwkCM
yuoMm2ePKS9WdH0JHPfYGgbKb5539cbtAbst8ZwVf01752Ws73aHIb9s29fmEXMa
p2mnHyj+e53tcfUmJR/8ojR3cZpuzUgqctaTWtQT7ng+lrIhk9TbgQ6p5A6RD+xA
AwI2J6SXH1RQJbfgv+jt7owyOR3Ftly9OUWfKwpC0T1IQOWwM+NQcgCHhBFShZlx
Bp4q5QT80sLiSz/9m7wsZLhoiNkGDp9qRHeNj/iobBH9n3fhVogrnM4+Bjx37n0m
lM/xn+Blg8UrY+CkBmJ4fMBbq17DAhpTWyOCkN1ufqQeeqKQk+/sZnh+43sA69Mc
Pwt3eMkJlHGP/8c49OfMDgXVXnMGqLvsEDWkMzH3DuDw8zo1SdzqH/xE0rzwMnzy
NMJ+6TzGox7GCVrSgM2KgHWyWg3u1cGZhrmtpovkRSo5/crrqD4Oq+v447k0x2Be
JACEjAQfIpjyL+kgYOv6WQbsyO+J4EC0U+Kvk9+eg09QYU3ykWM3MnTGQ9Fb/tp8
BdouTBCcFta/YFmyQ4QXQ9Z5yUbGuoiE9Yp1TvKQhQGL3XVjz12amZ6eWnZAWOKJ
Zkqj5OX6/y1EN/VErNvjPu1tXW3Mp1XaFL9yA64KXTOfJH8iDNATQ2DfpCTcIUO+
315nD0LQ5AUxZ909JeP9hy/SSXAWJSChF4taqDvA2n9ECkI/V3LY8hEPZaduRWl0
yDiqmpfXs/QB8rcmKKywJp5v9D92+emwMlPBp23OovcssV4HWAsq29jyVSfyCDuX
3OeQpxF2uB3zA6WpY4J4eH8BMiqfF65WGBYyEN40de9QI+RMgzv4ZbvyFIbPYft5
ZHFBQ6K6ts+OJuebW/XTH6NTTGaHZCqnBlLiIDh/NdBJpkdK+qpMv4/SUp6nE3I2
ZPXZWqv7oFtXV8IH2XGT3cfzKaZ523ejsPCtgSMQrTFPGtWhDbOaEnAh9VlpgG/z
bX+4JfE29HGZ5aXbATReAUjGNBgYcUV2PQsfWhRZskER9So+mUVoJUxzFmyIk/Bk
zMdg8iBQv0hWbSoxgyQsO8/vOrNe3n5FwOF7W8cBvIh16ai3kJ+so0GlAobUqpov
KKtQhaatsPxFPJX+aQHaM5jZh7Kagf5uF764hmHu9OILyHwroVVb7Jzf0Gv/1OKr
3EtlopYgPywtjk9VgymuQfnmuJ5K7VsjFnbtKOVj7RRD1tWKyXKgKBZnjMHtK5QC
g6OsCYN8XIZirPJ3lOfUQ0hoLQiVTtOrV1m/gonIFaFUnQoYmRsJawvONH6rc6OJ
leH6dUrfF8NnHPq4EsfkhZIk/xDiXHypiCaOXBsJcJy9Uo7+r8wfXjT2g9lNLmDi
Wh1fcugIvonMf7DaiGZJTr8J6QSIAcJWmXENjwdhg1s+9q9xybW+/6MycFljc9KD
9Wh5S3Ku3EmjitV4Sw+baBmEa3XlEWPHMPWwRog4pfTnzEEcNc9WInzYqeOo5pnA
v7Y1Asq0g10ohrIGQmI0fPj/zBk2koNfehcuwnMiIPd2/5uzy0cSWooTMK5ZjEZr
YDYN56uIb14I6p3hxZLW0/YETUVAZ3kL6fnQ/k2AEWQuWafskx+rSRsM7GCNSJpL
I2h4WnNHl24gy3jM/yEEbbYW2vyfAid71MOB05Ih7iwOZ6+4JfHmlvBkidv5CdiL
ZddY2i2UjnJGYfO0eLi/hJARCxfRe7ZgBLJFckGkFjOmFMOPTjAN0sehVqCquRmK
rn1oSnM6TZOChB4YBuQhrhid0UhTCRXEDRDA9jdMuYyF0KGuGZ2dFWzZgb6AorO7
3LeeK3zjHWdd1gNzjYC2/FJHEip8kWvnySjRw3uSaVz3NEJrrtXOMSbKRmv+W1PK
AixoVleDhXwLti13x1RgGA4lsNMS4RH2CqBZIQyb7poqzu+8bAwAFZDohgGdtCYU
t+IRbKzFU/kLXRZkR5QryHAssNCddcPNn45ZWN0QzYQDyVe/QEaltLiOJlDce3Y4
brRe2gcOq2RXQYlG7dbKrqy9vKj2L50KfqSxwW0mK4W84rjk4mR9SCixj7VbMGuG
X3/7dfvJff8rccoTYJJ07Utb887CKmmqlNvalWLv+t3z5Q+Da6g5LAvlLx03susQ
e8NoubXvLdffGUoeDltqHMUtJwVC1+iOsKcH9cgxjOQLbnsv/1KuZnPan0WhQg1c
D2/FWxeVAuB7ozJ7CXw8wkEWEKzrs+WTx1V6/jLXa+IQTic5Y/UjRpqeSVaGBuCx
IhTv0K7mKhx2zTw6y4hYRWwPR+mgO/dsxIbr+RW/vFcLdyf4T7fg2yl3+BiaK0nv
GCuckl/RST3Z3xMBFK9fd6TqKFmUtf2KRuXM7WzXUSqbQBw8X1CyejdFdr2ixNX0
V2hXZzbSZFf3c9gJbU3Wft8SFmvaX+bitxSYO2JjqqT0TDUuKwGlbk7mc1gDb4H7
HCwDp7BMHkzeQ1NQxf9YGKmQQoN/BfZ+Q2964A8lvZfMtTN6nfBygqSRmpOjOwIq
mYtiqm51/4oCxk/0rBCS0ubc3bpTwricxn+7d/Ksdu+ZCtU3Su5JhXmu14u8/wCZ
ZAgLVryOjSdob078x1SSTM/hTeGHVDGTjxI8IDaEzFAaQsmV4BPpi2lg9XoaSwB1
L6TX1l7SiYGChX5U/ePk/COPPTU7zVuhIDlUXthtltqrDuXTQMfpjFxWqEZUSZie
naUfYO7lAMCRBnm6cTC6dwUn8VZvgIJIN2OB9ojqw29LPSUFKctsWlM5tbbDqENp
hz/1Lv8UAmze2q+QSQk3uhnOv/PjhDSwKVVvV0uKsRFO78yISpavlh5lDT2oMQSa
asaDJQjoS+suE3jRvmiDfCGS+ymjqQZ6iBvTbZGHAi3FBXhbefjQi+V4ptV4ge5f
SQS2e6De3BC6QD0FHwhVaKx/L8F7DB004IkprGVon8bHg1XlqEoIHqu92O4jTqgk
oborSENBNXAvmRg5UwTpncnc9GpBpTQfhOgGRXLr9J3TQ1fp8nPgOnSCsbiH9ZDR
VsTX7ghKU4ZkT7+zlwweqZdj6ynMuUqZnIg6wv0vpmLOc7YzTlch/xHyUCkRAIlz
MHnLGdv0FJxojQYm0GpXbbVyT4k7pWVQRPAE8eMjA0LbL2FSVOLrstYbU0/7PARY
NuqnC35qKlxUeSKj+GN19yOQ3RMrFJHcXjKIMTmk52IAMG2/9g1FxViDyvCOj+kL
HinNUIlrPGeBUtRvmFZc841LtI5DDTik+515qUCwHe+23x6ikLVWjcYAeWM4kZNi
t4LqaiBtjNZeCrIkNmYtWSUUQwpahamZqjNlsw1DCLVKw4VgAmtshSOjv9kZ2dNE
bGy6nTnpfRV9b5LPstQ8VMq9T7s+CFJ3RRns71YMwIm58wYTOkIEYLGK9PaSJ5vi
adB5O4m031/Q80oCh1pQW3b7Kr4sQuY1tA5UgTxvzPJLJoBAZgp2V9/DzMrvmpnU
EUJ2VNOz71ziZGKlTZro30J/Sgkx91eUanBup92u/q2thY62hWiVA+RW2LQpVXdF
saDKjhR1/wq61SGVdulw7TTG+UQ3+7DnU9TUBvnEk8jWl2FZYpnV0XiG9cFJK684
nzWgeF1ySszz5MijS8UCo2E07ZeDQSdthrB2z71drMDoeJ+vZHM8lSzX8Lz8FjEi
B3VQyHip8TuNRUL73vafoZY7lVqLm74o8vnAcWG93Kb1I2722eUYI3JrARLMbwIC
ETbG2njydeiWXpqKxFdrgPahRquWqdeSKpcrp6d+naCU/8GzDLhASOahKNM4Htty
xGdqmiXncHRH6wWan4N5JkO2pdTBFKhfazpM33qOJAotGityCpz6SJE9pePsxdzu
esY4BXXTNTui2me8H6sy6iie3yxQpnazVQH9Qn2DQK40MRKheUhNpVieFvxIYxEG
kaZ2tETMOxjIZl5/ruCkHT4BTWPK2o+AvnEAadgbzsqYL4XVEYEnwvjGKeF5HyIr
A3ZTnBdYRMaAG85mYx0n3cI3IAV5O4IbT48ZwiP6dAGfN9OL956iZRgcp7kDDuoi
VcPPTpqviNspbo5qWsQ7FFNLXF8kdZw2sey9pWKhv+yz6DusNmXwcNakamdrYvlB
8QFA9qZtPOm6mPw55+p5KrJp/FPzbujiYeOjeO1b5X1ZK6l5tRLBJO9D5cTBdQyw
dDE267reVbxo21bYKb7C7/nqav8rBsaHiXxUHOhpmuaV0bqo1wC9aA/7qKqQfjaE
WkUAtCdNqDxGEyIy+bHUIyrDmSAHO1YmLaoMNiRR5Cia2N/DUNOMUbYMeXUAtLAK
5fMZPMYkDxJC4mF6xg1dJVNJYU5UW5AKcHWHXDx8jZPB1C1wlvw/08A5QxUzn4R0
hWan/xBeSsvSG1rB5Q0pVOZdhL0RRdvmwXSkin6CCrhf72rha32inyFgy+WkKD/t
XfinJtI0lenS0ppirRP1KUyQF8rZw8MwUIpM/3GhLa1/fs10W0za34XiE/mrDCWv
2e7wlXvof5ESqsZIAL20MySDHg9i+7+4oWmIz/YYf/55rTU/g/wmxuYwss3opQO9
8S7vaoWrgcGH5wtlk7XiHSYBdd5ocVKq5e5DbmQXINi2j5ml/rA9cs0qL8cWqOau
0g0yRLQyZNn0c15mnRX8ZvlDGGAvfqYfi3A3rMaOLiG2BuMtyTQJccmpFHydXc7E
JZCp6celSz4MtGtpvu6t5Yc9oTsplxnTdTcilP+tB/ZNLMQPnLg47GmqR2AiEo/I
1+pIDAYxVKy+VWU7GAZpCVBQYqxuOPyVCILwjNVEQPIK6tOlidPMIuqWpEf6UM29
DFXDueAuOpqIzlFE/2CK2BmrjZCT3RZ4De0K6jed3V5kz/9AKPP1yQLDwvEi5dG9
sXFvzpZqM/EGm69W/WmY+Rt92HH0xuvb/Ag55gq+TbAS/BYpcCKPmiTEj5zBcZmY
IdYiAr7OAcyLLqXVSS5G1XM9389Et1dk978BuZDnS/SoNS/DTk6RWwXJbMzskW6l
14hdKyeEMMetlJy3C/WNDIJRuwnrkxGflEnhDqNP5QreQW+xtP7j5Hto3nVPzt+j
ycgeNNCNeCCf3TEkpi81RVUGmGvi7lIPcBsJxnRnBTPJaStqLLUlzZTPQG0qQNwy
ZUVydYZQDkSHuAf+6StxuzDYFWPPLMDmdsQgbadGEEJAXjof3+naeRIXgjQzgOjy
/rFFk16+ARqHFl2ec0DeQkHla4U3rSLJNocwVhj4IdGrt0xVmisWEMTe3CQ7+Hqn
fh1EkA15qcEDMZZjZOQKEB8dagw8/X4Z6bkLrc0VFYNiCAZ75TcBztc/HpaGErgA
JM09zlpMRpCpQx+4xONn765ezxchhAdp0602uTYj4FboRtj4jo0lEyzq8282OslF
B1dOrP3FNnrNGXnl8YuKvFb2fhezNtGBYtQuifw3K9mIZgOjXfBLJoumkbkc1z7S
f5M6rsrSjX7UEdq24sG9X1VZkL41hXioAgDQPB30UpIzmRZthUiNNpRkERfPtyAu
CJl4dUdFRh1eTQvEAmLnk+94bG/cIS5WqdPPgZ4cN/ULHKRb7+gY8lb11nwU3doQ
AoxLWwwyy2ZecFIUX/rX7/onidKeX+swPz6iE9FehyxQ56gSHbVnfTGsOhWHSZNQ
t7oiM+4VHdJ9lVheS3WMVtFSDiSnL7oXDdfPIDDNYBZhoTsfwUObLPksyRdsxlcj
6n5611ZsdOOjT1lbVKfO1CdHFObUIE05hfs8WWnlcSIa37XcAg2L6dpZ1ATPs/z2
ans57sbAkGsFZje9lqRR3bxeKoiklTy3bHK258fSHVCYVyd0EAozi+j/MeavJHlG
T9xggph34F5dKX0ZDZAi5qKGTQwyuaZicUJPIwfKcOiceyfkEPyLLGZlE0x+v2oS
buKqixG7eGeX7+FX5HhoGRb3JQNc4P4TM/T+Dhym8tyXYPAC6LIA0G3rosZmWSRb
r9xEIJu5/6xU8MRpwhsDlwEChLEY0iH/6CkwiNe+tih/JuO9EO7W524EQNDCxWSp
R+X0yq9lKVowV1AjSP3VNbJU7INOwEh+kzc1eD5ICvphhPVFRNYGxtn5ZfNzQh1m
AT3QydRtn00bGND3BfwnfJC3F9QR4jyvJSWALCXUNjyoRqsbZ+/qA1jZ1Ku4krCo
4QC5Wyuj9tt6Zb094kTDyx6O0R2RNa9Je06aWQ/8iUlSZVT5vWhaQvdJlkLgbh74
LgsbFXMraIUbZOlkMp+5uvMV4Dr2CZoG7V8EplwJ7/5xTP0I1c7vh7FkQhNxjP7n
eSgJSKP2a+4gCelfGewMeRCreItACi9uo8Jqb3FKT63ClOhVZLv0kOw8/h5HiY77
qqmztxOtLXzvIzDsZ/k4zXXEcEqt2KsDpoYkZjxr18itOUTP1kxkUm3I+dbzzNSN
fybA5l18kO8Dx09XNjinicKZ6o8w/F7lu7OZOER0pCwz0Z11By2jRtM7Fog5yJJG
MqqGd0kbwYPUDAAzgkO8q66taxuxPY79NRDONQoiaIluUz7tFqEd4/UJpdaa+abc
nuzuGHi2T4Fdjut2+VPnsOGqowtwGgm4gRhB0mPymRztu7y/knpOB0aRz3/Y3x5b
2O71imy2yytJ7krhAngshCJ2/D9UVwAl9bQlAYND2KGm89ZYjALTbyY6KSE15dii
NJ9mTBKulwRNmK6QmlXEM1BQ8rEPJM6r235DffKKZZ/ICZ8ndvewwU32hzqxjF6J
fESwbLrjcGz+sWEFA4twXflG55lef/NO3QiJJxmNLHgqVU7dfAhJ1KwbPakH1M4N
4+Y4xjcmJwnPjOuZ27RKldPtBgS8uagpx/1pp7RhUVx8UfU6UvzmO9rPqRMblE0Y
9DiW+MsUlqwJxrMC8UCLp++NLzALani9e+nREIJwgF8GndmKnIUuGbZnUJnMQ2zc
Bzca6bqUDOjtGHFX607mep0EfULFNE27yDEqDTamzqHjxkI3AIJ2Go7iMUREQULP
UYnDD8mNvIXaYxdialQGpKNu31PBKT9Q3UltRRBJwr9TxowQi8ZVWvN4h6deab4n
dFojGGiVpBNtJnpASWHT7+ITsbHWdoL2QcS0aPfpPpZrtw+m10JO4X4E4Fm6JRMc
EXKEIuuiqN4OomPJbpNXqBc0+l53knRxlzmlGDQM+GO91pU5QaE0uW3W65l5IQ//
+q+nONG9qeZBfU3u7v7lw2WpNgJ6JzhT37Vir0PsZIdJsoucVYbzeqKffN+b6tr6
KUsZsd5P28pBaIkX8y5uwD2LC6CfVGWh9QRrDUze+VRnygm+yCBqxubXQhmdDePm
yCdRJjKuIdnqPB17ze6TUQwZYgzGagyzn6Nb9B8vcQeAcDz36V2q2TbKGZ1YPldy
ouSx+pEIPocK43Kb+SOIsUYcWQ6nIv+vsaw1ODIWFTgbQW3e1czfzKy06zZgDHjk
DG2D1IVjF2XKbB9aUipFqcEJdafLYt/cnEllb9datkrf92b/MwAEsyUd3pl0nJE2
VK0QJHU46vXpAIR/Z09+Dq1sKrys80527r4WnxRC3vRfA8fOO7dkSyo2UD5Yc7ml
8OtKpHGo4YpUriwXTEreTBmhpjgqblkthuHPH4VzAUJARtm61iBEaQbm13mCdp+G
RuFENyL8UkKQR9/+B3QFt1fz03WkYNciyXvQynqnZvY+WjvYBd38nSI+WBBhkePm
T/F6zrV0O76puTQw+s7087K5WrscrqSiyw6qG49VOFj04SLNU+o9MtfsHfQJJ1No
vKPQu3brCp0hNUJAPzofO2H/Ep/A85yfErws1tEr1wT60kyaS0h9+5zTxvnquiRW
ok4uF5Nd/lgAEEV/a9Fdvhrd0EKHfRFRzzei61byBd+MgAEeQYxYoqgJgwR6ZO7c
j3wyqiEg5wZOaGUws54ktqzcWyuY+Cwik/vft6C47woTeixFfPuDpD2+gKHZxPYO
7KBhTF9C6FuxVTFS9cIfm3npLmTWqfRcKGTqYXnAqEzKzig95TqAn6dKpERFoGIJ
zMVNdetIZrEWQQtXfkTybxTTxuLaOx3/OJF/bI1PQDlUjw2I67dcgnjCcTm9xbMs
Y2qgMBEqiLWVNKXSGtn2/E+5+vy91EUrVnHqUMnwfD1oKK5Tl0Yi/lkV1hDaqhap
WV/5ewrLc3ZxS78FxNBAYtCiUmXVBTkhGcrDU4DpQFM49hMOueGRFAa2pUrs8P0N
yg/A5dohEs3I0kKVguBofMH5kmEl0w6Wkh9Lia8pDh/daxKtbKh0VUZsLUNMNNJc
xZzpJrWOOYsslZirBu5ZVLsr9LZgOfZinAQ60LSrcp8Y1m2r2n1CKG6Wsa5dv9zR
c1GQs5w3gvs8ZbUlOEEBC237dsoDLab8eXwwDNl3h7mBUIogDY9NlKiXIEBoGsmB
GFdtjOSO6j8KBUthBDPGLtpdaXirPYXdw28H8c6lq97fyT39c5I/hZ4m31trYCE+
cJoBU6VxGlKS8Arlwd9rqWHoMKPLmU33Xb7GanMd2y+KiUTKEjSPyHqoe6WXXKHA
2yHvCKMzQrIfwW/SaVeB5kmpt9fQTeWqwUiNDHGYx9/4pVjhwBzVM/Wfvd04yjnw
3JvexffJjh7S7nRDp+NdB5RkkMNgHDVStY0EUFwVL8BwEWAoTbYLE5B3VLT26sxr
TK/DaX7c/BcA6olPU9XQYKSqrxm5InZnFvjEHCPCeiFLD+vS7vFs+oYdIBPZqOP+
xPhSU3LOs8F6plYE0QHQlIed++nGMeaZGHDoQ9bUIIJ57ztBLYtVxxNmG13Mtgwy
UNEhfRcQYTTWwpN+iKluTiH9Px21ocDKQyiw/JuSnOqbpChf61mtRRwXtyZJ1rtl
p7thTbEytKtm9rAXPygQiUIjvltd6iOqD6s65ys4EFY23FOHchhcexz8x2u+t54o
z5tSvw+ytqUWEQkMZQke5RAHX1DSUvy8Bdm2Dwm5rMk6zmB0+KMsYsh0fFkkVIzi
lZbymnRKsUN/ZA2fbBG5ZbARrX+zZ+zC0vlar0jMUmB3jz7Bv1MdLeoBJ8Gpdsy1
txDKLBysMB6BKUAufuIdj+xwhkmK3a4B+hSIl32vwV6SAfaOviASbq2y46dec3gG
qbcWFjusgXqa9tH6fB8IMAn7fon5Mh1cWL95fO2VK83aFSqwgY2cXYy9V01NN8QI
bOt+7h5vUOWAxZuuBWDx8KJBZx0tXKuWdHdKXRljohhATLux9YxXrXyaF6C9+EI+
XtyXeGWbit1Vag1dQOVzrKW7jNT6M9z1D2SxL4StnDkbue1NtmlQN9cRXU5qzdLZ
wQOSW9PyVyWIWhk0Ojx0p/XfKyMGapHr0yJKhdIuWh0kYJObKt2gj8cglv5pdxt3
/PmG+KS1Kq6SGqyXc4m/FQB6U0ksXC5HETMRiZWHHsRUXeNWoUjq2M9U+LKxGZ42
wUFVbJIZcIP5n2FalHzzUOeTT3hOJY+buS+dOAKOAkO8q7JWKR08tcgj6RUdJQmn
AA5BcsRnJwAtE1CGAat96Ulvsjute3cA+lUGWnMJPK0KHvqYGQWuqvZtqOIDW1oW
i+Y0j89n5IlMbzNJwibzOng1zJXQgdeRvhEeQBI5GFdlrIT6Mu2e/M1bKdZPtec5
2ppHun7t4YqmIvxK+qDAWImo6koSJSac3woz6LWBgr76nMRCP+aLx7sB4P0jrP/x
w3EKujFSogd713HOnM93knB+kUF4j6jNHPdxiAlWlvq8eOKkvnsZniWg7CfeIG/p
KKvJs376LfbzYk8BdjH1kaVu2vTiUJmBhlPJtzbP7JGAMkN+x4dsDYYpgUwWwG8h
e8Qe1a2TlO2k3eazEKc+bMuyx1xllYuTDSdlHi3fzoWWCUFGRYgriIw1LhBSAhWf
QkYvHXN1In/1X94+ZSXZZ+HIJhXskS4EU3NvHhz3WiPRAkgri4zyd6CNZ26VaekL
2odF6pjdGhWnxUBit7vqD2OuBNxhLnz1vgjNjIenI1DWTHK5AOb8xSns9DEcwqVQ
Jfn/y9buFbj0FG1mBtBmV1lcg8nBKhlW6kPP2TAXM0s9xOiuMRCkq+5FwZkVddJb
N5/W+w+qU2Its8npJPNliuV0cwat06q5ZVFwTMrba7OqdVOxWvkj/Lm3AEowDejk
pSAiN29FizRELlS81oB1j4t8Ds1rKvmwOXb1hnkjEjjQPwqW1F95DETOAl8DrkCx
kSl6e1TcM1DMYJmumO3eLlGWRM8w12uk1RVqSqZVv1dbVh0bumcRP5bnT/zIXrPm
5Rw3JjpiWLcna1OME2wnr51uRxMx5Pufpwgw7nTc112I1uJAIR8npIuM2LbzE93n
UxnYbVPpzMgpk4xx0tKWWfxrlClY/ZytSBMS4H+7sXOMOwgFIoNN5eoG7GzLFSR/
Dw6tL7+890FpSlecXlft263qZ/bD9AKVtwWRxMwhizzt76qpCqLkKqAlKIxkm400
BiNWi12v7wnzEPryno+CJMmCSMe7OQ1XMz//wqkPl5GqOSjyrdxm6FL4llP57iFM
VXNI6i3CgXFEeC1OMUvtFv4BdavhUZuaDyc1Ypodz4HKCqH9k9uWrnh+0yCqeNpX
Yes/vvxS9mcnIN0P4S8UEHdTXBqKNyCBYO31XN5vt+S++tqGsXM3nz796AqlGT+M
qBhcw2FUca6ZOfw0oNqfGXyKUDN6PVJOzD8wlZfCpZXg86KtTzUe4aY0pbfAlIq3
1wDep1eRZ+TqQ7s0H7BlD4q1MBJ0f2D5TUDYf0VX0R9n3tueZ3nRKkYWThSOnb+L
RdFe9nt4eeK4f7nKliOW+Bb5IVeuBLSLk1XkjA5/oinWbgnE3w+X90ukmjYpmTjd
8uoyhVR0AMMbUBwwxzG31Zq9+CS1q6x2KA9J3+Pevgy2o1fkbi/J18D/wFBqSab7
7dfFxKGz27U1vxAscnUvN+wFu4i6RKPio4NYTZuC9vAPM/Uz+rE5PwScNzSJOHes
AjHYshJCXQYAmLJFwtZ1XZyDdxNMWqaS+xBqx5h9z9ZVIoweHIKppm8ahHf3yUil
EFmeLBXF/LkDlRAcm4IlPmq9pO6Sg9AzO5OD6NT63OkeKxjkCgxhUsimnGrozsUc
1QkOK54tjWkEtYf/lspRk3sNM16Jjo3/wM4kLrqnfOyooCTqEhd/bzOLYAynHs1d
4Ec3fP11xqRIcQPX5ZhM+2MYlXiN6Bc4+2coE2gElU8maTjWrhqGJYkuMxJBJ3wm
5QlJ4wRwxSrzXditBYmUTaXgv/PHpXJnrfiZc73GaIlH0z/lF1gygAn9qMyn9eXH
YmCR13x4HQnscs1eavB0/aV/KtBwLxRooFyuDmWT+B3GII7hCNszwavo70hmyS6t
B+a67WZq0jk56YALjPJVnZt55BsD8AN0Q3qUB4Hic6vLyCkpm206wFK1f9StPvPD
cOyI2RTqljuJNs4p5DcpHul/4LxgajofDr5+CbDd0RDe6K9gf6LZ5pjI/UfyXfNR
tn8ihfKbbvPI3jBzpjzoa3zqNqphqwoMaSJdHBwJZ8xYy/ENZTpiecJACv+puaC3
d6jOfLNpEpez/V7tYDcrriksGA0Sk8anicYaxkMa/YlHJIzz6zwoQVe+IOOe4lWe
bU/MlwXetWNlQPQ1nu54T7gmmxA+eaUH3NWlBU1FCku0xR3DuhPLlGLx57WRp6+B
+Gr9J0o+dWYzs7CsIvGskPm7sBesr0ZVhfhx6QLUnjypHYNmmu/67i5180aXBZvy
E9JUCnD8qqRtL3j+Y+Pya5RK75bQmdppHNj3S0HnadnZsyr+8uOoivPsX1TTLOw0
zY7HVwTTNJL2OMQHrjSrTSzcMRR9IjpmseTIWLByFeZreYn2QB87N0Ai2LDR0l2c
89XvssOlFzoMef9CUdVqKSTSxcPxPmjufTG7MmNlVdBYwrwiQ6qGSHuoSJDWko2V
1IkqJvTgrAMYova6a32R3XCG/G3/kE0sbY5Dd886JPZPBysBVcp3g//IaA9Q27fC
hvCgCTFjGRamiPwwhIaD1pG1UztPzjzCos4gFs4xSet1WWeS7leCDvdPovbwXF7k
GUN/d11NYB5Wu+uwXtbxkWGYnVvlCwdng+8el47riMDQdXAqA1FeRreRrHZOWO1n
z44kQsIPqMLkzd+uWZ5hs0ppKIrlkzoXkM/zBaNTY1EHBNidS7L3EFsk967dJBOa
5h45caIvY9q5DBMZPvJBf5T2Zbsm5a2fHvEVliQAAutSm+QQQSRpJED61ccS2QL7
3Cm2ENmpcuzKvqNqdGEa9MoJRWrUeZTod4kFirkDLVNGR7BSXywH0zb3Jyt3/4El
spuLDTKsEGj1KPs+gVyQdg/Bs9UaqfmVpXO4JAxueqz63SkiK9rHBWWPfXi+VX30
DGcgXk/qPzqBlFjiJoiDH9dYfMH/ECeUP39zoEIql7I2BxcLBnmXVOuuBJ8V3OZ0
1A6xsZFzh2S62M1HGcrjjHhtbI7fchMOy0SXzh4TBO2V8HDiBKU96XaKWmPqt9Y5
JPWLyddskrq9l9LDD+wIzWSThGjtyNg2Sm19QgKJCRyE+hquqQqyuBNLd/cyK9Yc
/LfcQtjJLLdHdY/2Q5duBeGEJKJldkjJ97C3JMOo9pbbY/+mU6HbttdmEx9Gg8FJ
XLjkAARLRV9s9wpWipfnOL0eV3LAj5bK429xvtsueHdEIf2Vo7fysvPFm4ED40/8
J10vtACauTzz7oobdFV4uRCRvpUbo19wexMBbK4UG4JO44o+grFMKmhRxCSvDvat
qKW3Ew5bpjZjT1Q4UTHsd2594TX3Zdxi4O+9dTDcHenx7SklgDc1y9qGlXpXdJTE
lJCcZbAEN6z+KCVI6jZvrxhi3TRuoQrVtOgKg54WeJ+gXcpkH5tjqzmUBRt3OQbk
3y0BChrwGoRGBEOs6kaVah+mH0p/0fEyAnZf7QqzeHy9/pqt0bUaqnVRF6IksPtX
w6MX0iLwAq6EVfIeN5pqjrv2GupUMreBu7JO8evcFPBPQrDuI8OPU1yLAAhe4hvw
+RfDBCQQ5W3FYL2SpttY2ZA2rum/9qLaPU0DPKJGwxSYeKz5/MS+7CgRY7LVTP3q
5Av3cg/yzqLJA5RiXIowl37u/n9ppsn+qHeRTJlrYhylop3neuyZyRCS3GXL/hJx
nzshy2ucFN1CgyhejnFV0SDOZBDwCd3PT0sK1HrwQo3huJNbbTL2P3HDnf9vKkIQ
Ecw0vnMnwg6I6YappQIPN7GekSPnpjUh6hxYTapFxEwL5IhkZILsT+98LXADvq0n
o8GOKkk4F31R+31tjMV0zgtRmLM3YbW0PaPXEUl/VxxI/5Yrmka6fbYHtswuPgQK
Zs3AzY+Rq/saPJttY8Bpn2bh0cmwh5BBMtr6KFmua2Qzw14DIwD+DI56k+2vK1pP
yyvK1ZNzooX+gtkxkLaMApONlCnzkM9TKeVeGf7y6p6JhgmrcFZtDZeBdsbBn/kA
fYq5ZKUyAXWYFOHYV6kromdhybyMdaRx2p4PFz9RjhZZZ11Fa2Wmi27cpsqro0PH
XDEb1O0ih0Wphv8Bq6PGu5sCQHuD8lCtfATDluTzS0ZWKZY27f1NXD/drMVtvfew
VlzwOaUNF6uyF9pH8eVWCoc2aSxbMeACiaPJXKM9iTc2aY51Lds7wCsPFrrpIp3D
rz7ZPx68Y8ppUa20dbTUNEPjSseUzcml+z0tznhNmOqIPsw4L7CwFBRgFjxi/nv7
tUQ1Cy73qA1JM8JgxCdjgB+XHog6XSF6YtPYF4iy51JI2OewTW6GFwGtmf1mcEcE
amlcMjrtJxlNGUd36HxN6NJJvy82CrbzrHkGJHAbtlTF3rrVDUWlXHGIxeJtcDkG
z0+6y+l4DgH2KxqhjLV56ClQntMT0lESjMCMeQ2NVPRnXdx0H2YBGYVYg9og+WO8
Kj09MEyKfBLcv5tsC9qNpuAm797oy6wvpd5CSLBEVtmI86IxhpKvZDuHBh7OpsgB
vfryLuqyBRQ0HJz6epc98wFXmlAdVoWKIuPyQhBH9aGJbiI3+FhZ/Bc24J2jYzOc
rAoQU6JW/R5Y89F1TA4Oj/35Na/PeiWHpKur2/WMT7rLPjASXBeHQmrgb7Gti2Bv
w3S41zTQ2AOZMcVdzB8+xvR4FCyRO07qdkR/igXE3iArlrqh5bwRDLCmfGww4o25
p7AInXyLU4BOMcHPqg7qvqrF5hF0fLn3WL9N/s8N5lKCe+FVNtS21L0/KWKhdhpW
yWkfVfqxVRcB1KY8sOVtGfMK0rp+7/so0v1Lk385JP2TpcQEBCU7SDhV/CUSaret
UxtBDlsnMjDNDfW0vUlvNgRLY6xocUPJEF1Tebz4iuzwDDnYwxHGGhycg12Ol7dU
2VKq4HPWYl8JNDSVcX+L8ljEd1DAdIRUbg6JB99TfkMkqn3rneMfQup5bx7BvtYQ
lxqBza6tCm2tZsguuRrWrnzFTEBDKFb4E5ysbF0AyP4QvIzHozpLgCWtLCrKjJK3
8gyG0TWn9FPD1tIhNjvQ4eqnXwp5HWetg2m7PllzNdIiR8Gaz/kQZ3pzYxR2qTyi
zs9CJGhdXQax99RjGQl5DX/iTE2acKF6A8GVizoKLh4mKSZqUeR3c5GmBkmm6G8M
eX72zjXqAszTZFWiHoCVXi/EMTFYVKasj+aPnQoensTWpLz0X/9aGwrGwEH6MPvC
2aXi0u1JqnOsOaqmLFhN0MLmtzmxtDKbWnIHi4JLXW981e/IA4QRiJWzK4ECfk0Y
FOiEF7ERM2bbQZVTY6GkSdcxXB2ET7aOhQHfWLVdZCsNvYoMHBQaRJwJbVxVGOKC
C5tKszxAokWEqxfl8kc7zGchkdI8xWzpM9fNXBO/85zpwSrWX5lpxkPuJgLoqL4r
2wcVfrb/zvZQMH0/FImJyUNaDPjX0V+AAF0trAvd2YNgWmcPi2e9wkLNQX2yK2yv
Iw7XJHwTAheluSE52HLueI/vFSFj+ZrYAmnNqwwnLb3tiNoYXUCZ5rucaLuElrMp
d/DvniSwP7y4Qm5K8xw+dG2L6LV03ZOlCbdGQE1Nbos2rFSvIu1UvfW0TemqvoZP
nSckh2ieQ7LK6hHxPir6gn/xnWWztL4TJC+bZiYaPl2kYjodggNN5itXSMfYKKUU
tdyenIIlc6REiIuJyOpc9nzmxm2Y0wFv2C6DTdh5x1bYJr6P9um2QyChvPgRkzwf
Yz9lrLHFeGfY4ukhKtmIP9OfMY7uQziMoH2Xyi8NfRNxBqm9Tug+5kFvrY4DHCvz
CmA55je0NLyfm0f056/2Mf7qeM+m4MzUQlzYICDD8o28aUdodooBjWj8Xs6vuJ5d
2xmrq/jdAqyULwjR0Wt7Il5gBAxJLuAY3WuFOhkZ2Za/NPUHfmhc6XmjKR6QkVeB
5br0OOce37ahLWd42Cyj2IHPp6xJihJaJl//s9+9P06W8TYJwSo5jmCfRpnL7rBF
2dAHsUrGy2UKaVXX2treHrc5CUPgn4rhaEz4W89mwQgfPu5v04+nJaHyVfsLGiMq
yzA/8Mp5xJ9kV/fCjBlsxa23Pd8/vX64VZGLEeKF8To7DnzSexmbA3kZgiMxIIsG
/l/wPpyp45nozdB8JsrNfuMySpZecuM8PIBNdCldM138bkUZNqpDtJHRQufqLYQi
yIrCiW+jjy0x9UeRXLJRRAS8NVDF96OGgOYlKJ45v28a8m05HRHjRKVztZtmuAxg
Q6AvUiK0p15aT57Vve8x7ONx1eE4BzDlXAhNmoWbrDi8QnPVfE4OMfYX7uUUCU1c
rqA3d38fCSy6xE49iJAcTayCYEZ5SDCmU1NH9cmUhkjgvrNOdhqPbny7Dz3TR0Ez
Sr0EG1ycLZMF4LjcYwb3G/GQciDP8YhAc1u61XnlxKWAUyg2e9beieOCLi87TOFe
ryw9D/dd9OS/9sfJVpA2eN2yvoAMaIp3VwqskE8gk/MCmoeGNL4Y3XSCumWsotFE
TuFXL2HAsXRmnJ+Ad/Z7j8ZoGxY7yImHTttSdwuGxuHOtLcQ48PRMS4Er0jzb/pE
0fOKtZgzMF/3h9ZOe9SjGS+I2sUyz2yNJ2nsP1xgissOlTUJHT0DYMtASLXbsYvi
ReHwNDcPPmJ/VXYH6ajWVaRSq9R3qsdi0JAHuVqZHeYRo1KmgJzj9rmO4iKSmBwV
imEFBkI7V3BucFIj5sFwdW1aq73aIt5CGx5MW6jjItavdiAietAnDur1vQ2uaIyy
K85F1bnVhkqH2YenDE1YRO+2IFqBvACVluEMRuyRp3cUClbXo3wrsUXwlUaM7tIa
N3CTAsg8mCasYhHrQnZQ3Cp/N12ayxLA7YKdExqJxVZWQy7f3BOXPEpis+w1M+ZD
QcjR6YNtuCuuOjSO4z6GOB8cCK+rNA+Tzcbhf/nIfoeO37YQoN0aq9OBXOc6DNaN
m+i0uakh9H1Q9//qMh0Ck7V1S+62rvwCrmTfzDNFYrLwm4fYyThYeaYi3hKQ88NI
GGcmhfi6RBMSAIxy0GgkmUsM3YE7CFCKa98ttMZlcVAYIrT7rJ8/+BnF9tZfmQve
QSHi7gp3sEcRoWjaC27DqVvajirCMEXg+uA3l6/gFK122UQ9i21C0xT9/3JMGc0S
j1NWZg6lIdmc6afgOYFdzHt8vr/p3zlaH0V9wUQIErHYCUAkM3xArtH66kpWkCYI
2ltrq4coO9LW0qFwIZqJTA/GL9ZvD4sFtwWwT4jMOhwKos657T5SDC5yvSgOKLm+
QUA2fnStmlxFPQr+SuXWFqjPB7n1TqhIidPyE3CCbx7hzrz5zUvMawsykUFsOg1X
bLkgkq+vuNYVqb3ppIF6PhTz9pwJBzdIPbwXuZXISMJlViXv8CeWftZs10pTIVlO
n0d9F3q7Yo+ygZHHl9wLgKApR021ugfdxPemvnJneogttmnml6YcUEPXhnPG6Ic7
kINHUCHTI29PMmB863dCfO7A4QuUbnNnUgzCMYr1GpMOW3pDALVqnF8nRi3lamly
hTfPvrB4DVNoc1Z+HMlfuhpds6SDkwIc4GHLYFqMvmrfcws/C54HoxrQSPHvwjjs
8dO+kyklB/1VRBFrquxQYZJMExyeVxzb/N5qcyUoj63i0xLL4dWKye9nqx9XkPEQ
GSwF0WkOC3o5rV119WvQE6fXnhpX1fucqULVxww++W5qBF+2Wqh98hxzr2PfCoRT
XjelrHPef0CiBA6B1hzGDBIoneK+L1/QiXuN2vAn18N/Vf7VxSM4BOyfWy3By6VB
CtFj5p8gYe0gkbkKvVOu2gyPJHuPKwUswnr9HVJeQl+pz8HR4lwBMWqbUlqcEVns
BDSPXKPFqD4cxCTGqKeuO/CaGK7wlVFRpJ4W4Dy0JFcXEhhWX3IGU8r/LXZWBs+r
SeYM56aBVGWPK0K9497q2DIP9SCcb8N424mpkE7o2TIv5JEjUA/esrSkMI8c/YD7
U5KwW8L5ZnMkaOvwsAV+Sg7Vf9z6v1ACBY8Bi99fTGDXD/yLwvQa4YF9CQQu8pSP
7eEp2o+o2h4bpbLuHsJVQvtAxPIiQRFIN91jGZsmnRKqiKmDa6aZEGYFaZjsdBLD
XZgWOCKQytkeRFMjXbHk9IwPrniYmSDwRGLimMTpdNq/HXQORQh6svGe7B3inRmf
rbp4kj+sSQMd/PgZjrY5NWUChCvFaXka4amepVCLKT39GfRvb8VstlOulQ4eEfKg
GWYGP+OlBsjSLk75BzRtpG++sA9gPqMsya9Vv9GSjd+jTBwZq9r1s5+1m8bwPWXL
hQBP9kOUsRmrcrcD87VvTMVrgsUlE4uIwSPpfK5Tcsop5Q/rG/ThDDj0nKUezpNQ
X09/YzuaTJV0be7pVi25jZLZI0fTL5BawOTFRVUXJmRGAQSAxTvIhgqu0/eFENz7
7GmWzuzXvFNiTopWpkqieDZ8CfM3alCSDq+5Rl9aaJ8gDwp674r4dQ6V+S3ZwPFU
EiFCCTpXaTgGmM/ITbAwN2sxx4/udOw12Z35V29cGvvV6zemgTy4iDUUG2NyU7zd
sBB/6kHJopNfvxxBh8786MxaaeM8Vmv5LIaIw6BuUpl+NSH/ovGe4FdvUxkMoPeQ
fS58wKtjzOYky/KjTYMbF47jbOqeegP/tFhMY/tkNCIKJ95Vga/Z/eIVpS3/bNTS
BvZNpHGIqETY36HEZl/Rd06GYytA4+BJJusXe8ZeS4EG/KPqiDftE58zQgIUakCA
jdYGQtBuGMuxwRhOZnp2QWOxtB97EychkeYzmozMcgeg6+HAF6iKgFp48Cqq10w4
Ovk1aOtiAcTgTx1QYUm/WxhpEVnbYZck3at7HpzAWjmCU6v0FiBC0l6LdCgQizTe
uJO3XPiLOUjkkoOPLAeEEHxi01oadVXqbH0+piyntzbhLB+wjeH9jtdUKRDkilJ+
Ddf0qK3gVv7589KtCmAMFD3Cjar48jZDCbPk9Ob0NsWFBOo6WuVmn8nsc1U9OMxu
t3nDCdSW5hu4E5ouKnLrYnBPxnouqCLZg1wGEuxnZv7XJJQGUeqAbKHAg/hKx3xs
nu7y79pxQmOAEurN/f2UYr/0ijbEeyugDmN+3ibd90VmeDg4ZPLmVPkTduYwNnni
KPe+IepN7eSYn2GPxgSaAa/9gzqCtSZVTmS1Keo4psP5fBMG1zjOfSjYZfrB5uQe
EHhdciXSc0wIwY2LHKHlap3VI74czM5la2n7XFX1Bw5TNf5IupTuxejEFCqZCmB6
yc+SjRnSVIA1Q02m88IooTh50+nfN/Kwi3pYYS2mFdZX2qQCLwGhCp+F1qN2l6IM
XezHl2q9n8SWSG7JXj3F8D2tE4NmNnfqUcu5a8ceAq2TPe/QMkg0A4wGPBXWYpid
pxtihSAE5xzQ/DCnGed4wpb0eFF1YB+Y0fi4T+EsK3tPK2m+y7OY4wGF2gaJIaFN
YyaBM6Yvi0fFBzZxGSGKscs+jUR4cY0VbGJIEJpiUKOVV9QIbzHNnCq3GhXf259u
ejQUgyoPrV/i04JC8ra0F+PauIodzpbYMxELW5eE2JDGpqfqNlNmPNPTx79bG/i5
I/xT/EXiBRH+/V9bo26h0os5TmvK4YIkYeyFwNdwmJLKtELIsdTZMC3xSO7wZX8b
thGxk0Q1Hn9C/R50nkt5gytBLZUjeuMJxv3j2PdNYWfGspiHOzeQo1b4524i2DMD
HMLgDuQFRc5K7fK9ekqjwqMMasZ+wlBOwELEqwByxbGhko7ti1wmSK/awXthP7+x
Tnshb67ImBJ177VnEmv4IbLsTfW3429qo+dHRRbVa39xlyr5uH+ub6HtvNy2NZ2I
ACC7qQobDBgOQOXRrhvBzJoXm+UV/wAkG3pEfeDLNGXLuEgk/3IVZxhK9+je0f8w
o0RU3xlhKnKPXX0YVKpT1oj3z+7QJkD/FNC4K3Xg7ZxJv0q9CsrykGxCiZSMqKZ9
KYcvBaAEbLMd0c9Ag+2mb3g9Yr30iaI1q/4FzFmpuxulzC4dO0EGfRBh/5WvnFe5
9icUip6fidg9fr2JdZAZ+mY9Xm5KWHC/qDTXqTakQg6R76wtN8bhHmnz/bwsRoxH
Lm2br63AxknX4J5u+Wl8rq93JSeEav45INqoRSRDGOgcmAozbi0owmjPRjnzwP3M
3pIhAPusC3FZLAP32W/uicCPKnpyH3JeKDWqM1mTqGQvinJy1q0Oxh6O3/0SzyW/
gp52OiPEK9colHEEFSq1IJeUvFGpMOk7976HzC2nZY3DUw/xqjeGnM4JjhjUyGF+
eFE8JyCaJUcJzYsinFQHAVM5P1Pphuoa93CfjxCkFv2FEiBcWn6Jx/v9TpmCjvdx
dJ0akwL5Bb8Jp4gR7Q01QwPofHiiQB0yPZjjrblY1Q6/WoXlGTEG39RzoPLKMHjp
MNzk80l/vGag0iIrljTla2cRCd57JSfPQbJ72U/PotImrBsMKjgaodQ/pZaKCGn4
UwWwiewNct+Y2QyncI4U8uUwGn1tDBLWEvXXquBNoNu/l4AyIASUJ2siOJmnvXPY
PslmrYkrWgdDNLHwul5g+Xjz/Iy4onv965/LNHL4pc8sjquTJ2A19LzToweyhyCC
j2ON1Co+CHr8qGcmCd7zJkzr7zv1CdZBPF9GWsBJEBImj1JRkaCbeRJWxZOCncGM
Qk/WVAlZHmGznEVG8cRMiho0q3jWPPjq6CWfGAQwxcHAwojTtqqiSnsgGiQdZyB9
icRS22XDk1somLBhuW+5CSq1kRufQl5KdoJWryu5lT+rYae+qq8ImguPzbCymY2v
OV3QVCc9RxRN8iYkfY8Gvkth1TJbyl+l/Vhll966UR8SFxyWwpz7H322lBKu/SUV
eM8yCqEC9SkxtrRa/nQpjG3L0HRnNRgKf3d8Mh4fLxAul8x7IpCyfpRCCNLFYT1R
a+wZOyaTRxUgDal2kgQJxJuxFdiVm65AqmYrl+r35aG06EgSzBuhl80ZhwMkHceJ
4OIDcfx+b5+u154Ba2hiAk9wHP0ihaik2QiqaAQomKtfDfFwtsrqgqNLnhVfEjej
CuXOs9+XczORUHKGzz0z9ZWeBAL/BQuPdpALn+Kxk4KDslI2EPKUHSg5twyTo3x1
el38MAh2RKqYbZFq2/W3R+vkPCPQfw2phTbMYH8UY1Mab1dIYwK2nAs2Dr/5Ownz
En1uW1QBPOrEFHtlAJwkNfJBhQ8E52JTtEBymd79SfdD7h80e9rI9GyPM9c06A9u
LUYLAYvW56cccpMOoKU/sTnD9EHHYS3fzdJVXagYnZlv9CLoss2WB94O4Whp9/KN
Bd9Xj6ang5hBF+vlPbUwDmhnO9zOCqoKous8mYi3uGcOGNXVDRMNk375u7lfowaE
Bas1sW1sl2fm/OiICIF0gEa9SRXzQ6j1RFnYLw9jI1BA1I4xQ7XkRhMHj9eg/umG
bizK1AnEwTt41ZjiHPkVEGg6O+TuXbw7CEK+YYG/D6X0FLR7Ak1P6kdEA8xLo2lX
umK9jVyjtnBMbNtZMVQ5cOh6aNanQczpre5pq6rXEBfILI6drgL6K11+4pVRklft
c2CrHcgfXEBTEwgbMdNE35Td6ddT3NJ8/r6BsT/lrwSlDZCDSV+1uiZAFX0tluE0
hpYJKNb78d+EmJKcn2TyjkEXBj4TXztwzRzAogit7mJRPZqh/HGPlqx68v04U4vI
biCQ7Us+9anBHDUMT9SG8KXuFMW3qiM8EdiA6VN4TtCBqVST+aLjza0RQlNhW/oT
P7bl6hYlGjvHR01jY2XYj+CqIEg+TUtuLhgdVnPAj0tK0Q90VzfG72vT6Z1BAtD5
JK3cnaJ6no1KYEkBbg5flxJ6VPreJ4GBOmBjLmcCfELC0n1u3LLjPXLVHIPlWX2H
AEaZidilNRqwIwA5NExugTq0Zmqq1h2z4s10HQFBpk8kswKT2tFjMjCgYHaUxHX/
q2DliX2nLgMFXdrqPFYaZt1A0qi5bTJpD+w0NgTD7sBaNRjDAGEwX/Q9IurGgWcx
Wxx7j87lbBI4KIokj/KccUKS1lDPOaxcgRJNyYJv+v9OARf5dQtZKlEjr99t9w29
MlAuJ4c3jY25ohH7hFHSjnIeN9gxrJ9sh7pI7n4SwYBQm0PDI6jPki3u98AFAoIZ
xssly6ueGQpuDW+MnyZjjl03+djCkMymrgd4y/dQOwTvWM/+HcNBAl3DyTmN+Wb7
mQ2OKrpl/0OZ5KQtwYVhO4Il9lsKs+EbnBcdwY6B+Nne+AQaAe6NlCeLId4FOlFi
a648iE8yoEm4+YGmmUEYOqt7PZEtyYt+Z1K17xopkSzfX8CkuYN7+vTH0tYB4QoW
GD1kVVySwjFre4OId0OhjuOXeh0c//VCHf0jC25PbvYuwzhGi/jloMqnVm+vCl6l
V6ggGWYeyaFK9AKEwhOUihlftlFyH24gb5y2dFQvW43GEKCtNC7qCJVlfNTF+/oT
/f56UgquSz1xOr6wFNN7sDUU0OXP5Gb93aacePGpHz/ydderIxpiEYxMMgvzG9rs
HmgY5kGqNQYBJLZkHctdecjCzOPTWxfBpCDYyuTeZ29Al4zAaxQ1+KR46WadAC4u
nOqsxQ425ncFzacT86q53fGO42wBP/dEpnpl8ZvzH0knRmaZBtR8oZf1DZZVQ7Wk
Gp3Xqw5oqgERPYCQrFoQDHy7xDce1dIGXW9IZCVeEP2BWVNAjAdGd3J9h1FGWSvZ
b/Sn+Ps6OSaNp5IsrIxODM0A8pD80QQSV30tanpPsZyiSHiiWRNGaJdB5gYY3tTp
FGei8qQBNwZsiHW2RbInwPWXfMdR4lsnmga8//MBwkdQlrmppKoQ+mJEyJwc0VB9
Ffa8Z5bzBs1egbYcyhJYgcT9Hf+4tDIg/NVOq8h8GTTN7Ul5lRR3/mE1fTd1yg7s
IvZUJ7oA75rE85uBtOl3enPu0bIZBDdZJoYDqz3xZEWZBncRPakcKdbizuHNiHVJ
SwFlFC1OvKiYk12K3l+mmsK4NYYN+NtQO8ActjNZnKKZdg+txPZg2x3iQASqqLF2
2g4EXZoMq3ped6SPJcmQ/sK6WF2jHuHbs9LKLI/jS3zL8n9R9efXIAA7G2qGk9br
00mt3WEcw0TXQAemUQojCEF6IpF6HNvWZoDvCqnLLT3oBrpYRo7Kr+wHCdc0ptTc
psGUlTUSdSw/QWwOov037SuQg5UU+BpNkY7LaueYT9Howfc20h3ZhLbOx90AtX22
CaTiWEY4YnGQkJigybjW0lAv41U7nynk0pqg6Et7bnWuNWV3yfULw0QmBkMRJhAD
fKSTqZH6oIQfSFNfDSHHK9L7L6rcHMOmZabaXE68bIy0m0V/EaqN1WWbfKxF+FnP
zgSavqIb0miPEjGBfOAu1oYfVofR1nF91oKs2ofYqPEMMJsdet0Vm1kI/0qBq2Kn
Adz4+eBssT5u8IFidb51fK784D/Q9LS+anSvULQKjYV0YqG5hFox4XwZzPexYR1R
PokkhrVHLGamEAh3wiyweE2/LjIw8bv/5uoiuw/5hiRCvx322BF661zqOHfGTLof
Vj+tuI/WDmaygrAz43Qtvhh5QPnf9XfZDP+L5OhYPc1e87F1LaOzM8pBjfYwcAsZ
WQzMAPi7LrcTHHTfCsJVlJ0fChUbAlDpY+f4VDMe67nuo7BgyPBoiTWtxVtAcO1o
r85LC/nH8SFb220jb6ldWRc4VPWSZbpVqogCc2pXxBDY23bzIj5AnLMvXdBpHVfZ
cUXkoW8wJqmDPDOTphpWtB6DsIvK06XGu+/akDUAByORnJiiZYPfklpyDtj2AJs/
xvjb4Y5BDUHbVIyLESVm1W77DFbk3a2Ol7DEp0VwOTd31g1xnIKN1AhHWvUzqdSQ
85zQVJ2ZZegyiFZxFQvaqX1EuIIg+rbMbsJ/TlC/Qfhurfd+G2H43m3VrdOwA6ih
VScGm0GubCDngh9odcedF3WgYhtr3P58kbUL6ql1S9yZ1rCBe4wQ999X71WKOlVh
+LEgJ8kcJUN3ziRf7y780q5h83xMSs8vYjQUk6Nnw13yXWEwmLsDk8RnuycMf7GN
wIBWXaAkr2byp3eAT6EVAp8h8p7/ibeuqCLtqyX8z4xz9uivR2iUU6z3uLyIl0Gt
0GsfO3MPzF+ea/9/n7+uTL1YqFyGfTq8vbDg+Xz/W2XyK5Y5iSOBsoGf5hbmcZHK
Dp7dLgVYyNpyvKQYMpsA07bYleGr2afgsz2X7pkTuDgWEaQcRP+qJYRSEt02v0rm
ODbgB/sZaINdLlWEPG3JCWKspYHP/cPZr+u4bShY/HFLAuu2whymlJ5MebtYou9R
WQ7xK3GZ2dsYWsj5NivahkUFc2U16YYN39WFmG8hM24HkqScYCUwKxCoUw+xJ1Tv
yrNy7q4MxFt1jTTYaodpXWpI6hTBZo23RAgbUB92r/7D4x4nCzuAzwB2Geho08Jg
nI6r9zJdF9Wz9PtKiPpGTxGXHamNtrKS+WUxrebCBRZd3/ntzFv5wmSBAJsGeRQn
jT5N9OlJYLeTQmfUcJlB9zcva4HV3KzznItk6k3HkugNyitcyx6whj8m3irVbTmD
QvdLtpkcVLF3LsHztt+Iu49dZUj/oKfmJvbY0Uxgi5lc2pgoBjg4ItWgUd/2ISmw
De6PuyhGsTCEOqj/VCAU8NDcUMSO64CTHaaRnhwW7JI+P2l6MfrMeRq3hkG+sHnI
XByakPA5nBX2XMpR9Gkf3kkUnHTrDqvM8zHePTP5LeaC/NNGlf4ZyNsxYEWkazv3
hmqqErhPp05EvZEYOM+Uo0/uQaw+h+eEfHrieUsjy5oOTbUGBKoWVvTFW7v3Uaks
HRUhj7O6EW5oeZqfDFIppekHxkxkzUGmHG/aD8dct4Vc/7NM0htWamwIE9bVzgsX
MD52YKECjh1EPYmdZUwQJggHdXTWTNkCATm5bm/Zf2XAw3hKDXbHwmyPVamxYwH4
bEjTeSSZxFo5g7J44K2BYQBMj0WCjI3O8qWmMQdFYgmAu/qKV371BTYe/0CEiVzh
GDOaRzv2Lt0vnNPVwDRSpM//aa+L9RmrNb77UtpSVq169STXiHSFa3QsERS6Fn6W
Skas/fyzMOaww1VwdVWVsrw0aB8wUKsqT1IeWAJYXDeoQ8q07wIcZytPpHGbI36f
hWKk0XBacDFteGHArBVFgNE6w9WEBeiCEEmhCJxDRBmZnfEykiCCeNnsShzsE08W
eWqySMRxBBDTueVRHGxuc7O9sbWXkTo1TJJ0J5LzSt6zMKDVB+wnOLmu3vCczki8
EwTv73bRGJlOXxaGhBahhtjgflAA9UwudmJqmGBZKvh2n7DUNHVR+ICrUL8YYxUE
inZfgQ1r8cCR5oOfordd7Rp5QmgvVS01efYXXfs5jXRTjFJxPzNE9H73y8bXiuBT
ykgOQM/XnMtCwyXLaNYUxI7dwYwBz+PDGO/X0SOo9vdplvVkohZznfvf7Fg5xmtW
m+NK6S8J/mRqTW+Qp0V0DG93YtiDXXbbaevY/giQMnrvwfgUkby94yi1gLoINbCG
0VpkJ038cR6RJMu+z61aqfafdrjP/TYoMTdIjHPxxOZYVlna0sIQRO4yuiUsMv6d
VgB195oJS/dHYbGopAcyv0eF5eg6TFlO9n6lgXhVfW6oA9bLlXauEGrwZOYs8MwW
W3UZlp1++ylwhftGbN1d5gEBhDZ6E+zb1MC3bzXNXPFAKct4YYEwK5MP2kpj/kTO
n/YXbWC33hakES/mXUkqxmFJpD6Pa1zLvWSkcN8SIMuXGJuJaSvCt3x5XAW25tAH
4gAj2RzGbrHdZJpPDy/BzW6ZXr1AgA7EZ/pfB33okvSJ3ktkQzH/7Opn5adAVOxD
fSfpE26+D/ZYdmmnB8pRCKncghdZX+xrOCcfzePERaSmjk5IqlbyJ9JkK/TwHxHc
e4Jj/2v6f0sy3UV6Si9WJK7p0jgITyjva4VHePTC69e7qE1xTTpsqnSkj5rVBomW
w2+BvURZCzUtsuENXRhqd6YnoymPu/7/RB5Fnjraj4rv5BPmfnOOOeUCRdUGYy2N
TuM8OkZ/htrQ75hSx34QDEZzrbdU0ROseWqBsyeBlYIBt8zfG4SJAPJuZttcKI77
521oCng2jpUoOr0UaRnfj5GW4NWd4+Jh6PEaB+H8dtpM3SX6KokvqF4+PsTKzP4/
xZhOd6mDXhcb63HKhej/7rW1OpdnRs0VRxShCP/IsBibnXSCKP2jnNTLFPhTBoY8
opjqynGMMb3AkGCWVZvX5+3NmduHmwbesArKJrIOJ2PFSWLNTuJ2HWVZN5ukE9uX
e5SpNydbaHU0R3PjZVAVg6q6iUFqw5lZiNEJkRsVqP+osGiRxUIrUnzoJa+vQymv
yqMMCbsYt34PQ0aRZdGL12tFEFwwzKAXvwfA6nb6nzIcde9ssZizObTyxIUK7uQ1
LKzNfsn71lfkC06z2Pge3Gw5tCTTHaK4Y6j/aIKaOjorm1eNo7AhsZwFVTzoecLM
RPpsnDMNDh6KGiKwV0ITVY0Uab1rGs59pMD5z8K1YVRjwoxuOmkN4Hsq5fTAgCfO
LzWKIC87SlCsMRma/xM3Dzsw7X53+vexkyez/Hto0kmWmCAtYAz4oIn3odCVQH2i
CwB/5hkxI/Ep/r2pOHftjLjVvFdz+lyzehHBfsFEsTYxImIiKVV7IJVFqgUYFKfe
FpiyxF+YKfLnvSAd7P4OTx2zDbkUPcO4Xz5AchHrbHobftDJ/UdnrkjqlqR+hK/d
w4MGSlIiYE7aiuzdKjskrZH39DwUUqgXbsgdLWIrPCABlM7G4Q5hZ9l3bQ50HVC2
OmG1JRaMqKGNf2xTcPhHnopNR0ViBMUXuBSNh9A4MdzIiT2pq6orqSJsAFrHfG5C
H3J83TD4qlUQLY9sldWvYBRGRRq9qexhsFxsduh88x+H6rnawjPqYe5F/g5QfKRE
bRkFy8+PVyXB0aHV9Mw5eL03z9qZItV7AVv5IFAcJXKMa4efZVVn1bdKuOS2bMbX
alnrsdVvQ+djE3GrcKv1aaAeBzFGfOpqKnnpRCuud3zjTlRd6lwq5lDzuNnfnQle
UkSszslaUJ0u4o3oYJv5/PfZzrrAeRSUy5Cf4mUMxBAJ8seVzDSP/pIChawS/bP6
pDbol20C9+KV9boXH/JDfEIz1O9uq4VdeuhImokobr88ovYXegTvEEPxZXy7yyr+
jgPrNsOHULmyikYg4oUckHlcjSlp1guzM60K3tC0RE+9MYuHDzmAzkpaZR8YBQEt
wVQ54xpAOaFgZNTv/QOwIozsfnkCu8wq2q7zSFPOyDzcej/N+Qc3f7/7yo6rgUCz
8d/79HUc6SvnMMO8obUlQeVE+7hmkOQc8/NQbqMQjQyVdRMB2AeFsj6Nivb2aMqQ
h4TRmm1dRia/fKNNPrlTbKkjCJH8AKUaZXTfllwqFBgi8tfN+G8GpPjitrTSp4cI
q4WMGsaeUTGv7KjxwEG9xyvLV1Y2JLIva2y1ry6I9zNEvfS+hWOGuIjxBjK/Rja2
ZwnBmloNkghNGzKVJezstzj96i0bPsUBYZEqpjW8rM9XNqOOrttjBuHWgDF54a4V
4uC2ZLnnarJ1udVvaxybWxA+md0uW85d7Q8YqZLIOduaEy4iio2Czc9oZ2xVZgr2
awGNJjj2kiJIl8qfKWL90jFGM9f6FdNCCWRRJYT/vydxvo3y4Ru2TVzk2dKiWohR
xxDbSi8toSTx7VubM/3kgVOLHtnWkrYV0vOcn/MqM46ZCoztM4yrOZzlgkt/d26w
Mqra+OkXLogbYFhMBiIA4cgK8eytZdyg1yqs1kNkN58fwjTLylUuTVyG/9JLIW7y
vTDOYbiruZTWfmF0RfwCXLC9J+kHEhWxt/N7NujqhuL5oP8svdWp+bFLxJTV9jzN
Wg70+/dEI02pBFHeREtJXfduJ86/7lmWtJn8IQd1Af5tPWFWgt9ZDZjfZzz1VWGi
rOS9U77Oe45mkQEL/1LspB1GtY4wvJty7RtEwkPbFQuwczhZL9Oh3SG2p7JVUiaX
Ec8AcM171vYs/8y9FfLSyCpbd3J+95P1sYEGljZPjOfkkU5zKwXvaa3G1E/AQqz5
kJOhKoBgTJnU3/QQK3meMcnGIkKtYWwU26QboIrKqcERNozdoS5rhBkKL4IOCNZi
og57RFsREFUsY9FAdAGYD0XmY8ap+uDghve5XnlZDQiHEAg4fRHVwM/51EDwQOJ4
8+zeZPWFxGzsVv0tTfsy3LO41+OrsZiOj+wt3LRCeLXlEsVK/0wH6yOgh0DZpMSq
o5XMF3zLYtlooYWizcbsKcWZ18JK9j5mRIXEcr7+uwKiuyLa7cPDM9BQUqCzFO4A
s62goUbdtFKIxSomJANvKZlS6qshCqsQbBRyElce8Z5UsoXNuydQRts1WVUy4TRj
JG+JCnjqmVOV+9S8r5MrN8eQfH4dY8qTQXDlkTzLB4jaZrclR7z+EGVJPVgL8Qdy
R85DBB4C+DwBymp3myOOOJ5t7uQYN/Ay0RM46pqm4pJ7GrLj7lWrADHu7opAegWq
BoiZbrXFTKeOgWi5DryGuA0I5pVBXHB2uCNBgN1CuVVv90DGFr7cb0bpasHDEpy2
xqbFBPjCZyPhgxiOvp0595hFAqRsm3mjrfy+A9hC7MOF+1VuFItaK8ihVEU7+dEo
sRRe3y44fz5rwz4UrvLSD0yhR4Vq4LX0X3mxP/yoc1N8+rAjRyyUvdSsb4Ezi9yZ
78w2sVqV5yce7XCgihioV8NjRNbnipRySrFYVM9B98xmg67fpth9FFNy4AhLnQFH
iLMubJrqoPlzvZSyckhztbYP7CRgzYu7X+GwjUzTDAW0xC27Db4d4sfiVxXOw6qm
Y1VnzAVx5FRwBqWvkyFwxDBvjxQqyqyJe0ow5u4AaOZX8luuFUxmOhJHTU/fXbP4
J3Le7txeEfmRIFH9ytXcGMhX0GS+IWkIn6WWRKNRIlB5bmd6llKfcMFAyANGB/cJ
OU5DcR6y/V0AxQIxNnfnqoaVcjQr/miGp5cTZeCE8LM9M/Unn6pO+5t2fohRtRA0
AJBEemnFaOKfWju2QjaEZu4DHCMYr2MN9ii3haMRR6dxFxOl2zUW+lBkbJ/pkJhw
0GOdQEJTxcBHbOCDlAS5L3s0bJ1EzNOp/duocaMMGqkj8pl1Cc+dBMCmzLmlDQEu
eJRFBaYpzLf0QZDAWJGPyOxqCf2NE9ViYcB6jiteTTyY5mx2As+Jikqsv+fd2mGu
eM4/LaAvl9rrTJwvedflnazm8wS0uYj0YeQ4gdPT517yUYGWdUOWqULM2FJ5zxxa
3PG/s5k0eQHPNV2uJQkxHP5u/WpIM0G3yVqcg/wP5Lq69RqfBGanin65No47TERB
DYA6MTMw0ksOguqNEJVcAdvirDsJJhXKzLvxGeL2WPc4sylO4xdmgDu/6cIlyDGp
UHSLLAczNAxMhxNsfRJWt9h4E3H3EudnIdCUGCKg7lxwz1JJ0sfWoVYkMlO0mAwH
EUwUTKEm+iPhsU6E21xz1yG/JIgSV31/998lrCK4/e4aIZ+EknmRf1kfHisbGvRb
+0RYXxUcUFg/KN3Nc40gUSgGJBaiWtFDUv/SUli/yPOQT2MHJvW5khKAQcYcwr/A
/96OiYUUC1q4IaTblaOVQsPJfSnlaZYdHmKv7mJ0Duotyv4v/bwIdOFeLZrIaKOy
YW3Ejf7ffxZMGZ2Bx+nyNhN44WBgjCTGLdj+++k86RloUjX+5MLkqR0piHhwnyaq
42uS93OElJKBrc5EulUWjp1Am8roXWJwy+81VCKORUN6TdBmBjhPrq+poH+JS4Q5
tMe34ZOGcnIt7Zv8wQ4ZwxIO/1HVRk5NQ68Mk/SCrJ40sigYDJL38PX3ZWCexAn3
3hx7vpv9DgwM0V42J91NYJi9WzQFf1BbZWV7E7UIcGHdrIkvyYrwDqoCiCzJwQ5a
IHVyJ96DEh59nR2evQ/50VJRYsXHSCsPMlGT/EZkmpBdwvQ/0xP4Rg7o0yUBxkt3
0nKbCNLKWx8rr1Q52RbDybCEtBF5GY0sZxyoayZ2u625g/Py9sWRcrUe2Dtv4hn4
QrgUTejIe9NouGopSBK9Qx0xAcwx5jk8k4TwD+s500fkx9rfQMJc00G6Jwf9uhkA
9YpvGh2c9gZjfSKRZlbvs7+9y0dZ49S5MS00pM7qPVytYMHZMsOMbt8V0D/tnby/
l4skf5aXQjQcD6kZBYJJYyqZoK2Fn4Sd9iBY8oha6nXGusdrxAqQjk15TKshPJMh
BrGhcmjGn+IXubk2mDV/s4sdUD4Hkpp6NlJJtnbPznBW8J5fZKSj//OIBKfbEMk7
DDhX24dm/ocbjdCmqYfBpdNxq9JFnf8OXjhH69NvtStFrLMrw/u49PuwwdvaeWsg
uI2uX4sobIi0XYyqCEk8MjU0Fga3N0hHhHEcFTgSvkV7RgohBxSr3rI+OuT/ImsG
LUnLF7JWsgAq5wQiKl84DsA0KSaRzG508eF8sY6jURZ/pmgK6bE7sSSc9utx6gPf
WeK29RX0Sb5qzvC16ji93Te1kLrDCfAvKGpt+5APJGTCDMGmUkShD/FM7f9GS+pL
mfbmw/zFLQxSkd+5+FvS7kcdWf4BFqDvDibAhXORYCPIOKy6wqSF8XKIJS3Ng3+v
9QYrMb+Uu+jfBh5BSzUITihirKL/59rbngsSJxMfP0v4do6O8kDhjbH0uQKRuCCl
sYjLbt0EjtXIsiJYRI1+VCh6iB8Wformw78tolqsadvloQwUK99KA8hYobrWRS51
Slqu4NRwSMLKUMmnYOcGdus9iul3C98yPJaa7oY1dS+6P625nTcYo08m9N2rcaDX
nKZ+s2c80uy6lUC9aZJ4c7ewEdBALfv6+Rma6IE6LAhV+5wqnMcPgOoCsqPLeOUl
vMPSI7bp06nd0EP0MZ5CVO+BFJ7LvoMS8Bfox1QdMkKVbAYT6CmmvneaP93X4gFB
POY96uvI8qV8DiUkuSgi2xwZ2RreN5TD6EAH7P+XV76vTj9kmzaNO/o+Ok5I8ICl
Pm7AB7DgpYHSrlYiXuCQootnWFREf1G15yfn5LjGVvs/bZytkm3YRoKq0WRNvd0k
bRW2a6Z4jrI1mG+pnTmjBh93O1oGn90aMOt+9GOXac5LPkVKXYNYEG3xoNGAE/nh
oC8SA4cK+FVDKXglH70PR3izcSJlXgAtuOdF3SnIcnNeoiASa+VuOznoScDugyjF
aLlij8bXHPgMziBSK6OuTmufkx93ZQ5Esixjo7NOHXfhmTn4MOVG2NVfwNmDPO6g
sPjspizpIsC52VqwRC7gyReF4+Q+PR5lByWac2suaimdjEAY8dTK2Bm/yqnVtPDZ
L6+ujNkeYvOc0ozojXFVkFYcvUA9hmGrfcNbzexKaDZkDwWdU3m4SwJ5p7swY3R/
c5F4tdK5HZgyxqZqq612sguCp2tRATaosvr9i5f0EWwzvMLZL1ZPEIehHuxhbtc9
dpXx+x2ovVqjQkqg4uNb82XtOWN2cT3EX3bPHWqsIhfyrMFz65oq/urdefp3/jRp
c0FPcCqkTwIqNcWQ9aLDSUpjoojnbpuhZzUsSe3KHNZWdFfpFTz0gDOBTuMx4NE7
UU2szUuapttAMbBI28u3Ngn7DuVAYCesYtT484b8UfbF9GdJU6agBmXDPUTUN+OX
BMHcBJUmGKll+E4drXXZQJ6Xr9MQtjMonu+kw8vRzt4/5fTJJZ7B4exKYVgT9MQ6
mqhUi1QXIaQSeWw/gv3qpwEX7NP7bQ4i/REW0CnTPGI2Opwvc7kfqY1kfLv6ssyv
p9jIVigJdUGdxz0m6vMD0Lb6YqbWa52WH9+EDgF365YOtQibUnGKGbXh8FXlzW3G
4U2ib5wQg6cF8MlYat68hMM+ZgpzHrXsyLJFdibIqeSOVmdTBmmngdZAhW8oUERu
dHA+rQvGAWQNt6a7L6NVm9jh1gRryj0K/yyHXrFJq5Ac6U0O7Y8iKc45dVdHlBeW
fbBxUuNItivA50CRjgpGDsiVYyGMYbQZ8C8muvwFq2r7gbLbeApVkAY1ZWJ9k/vo
Jwqfb8TezgglnpHkJlgWvW34nbcuylRqtYvT6JLrE7Crk5wzcRgzJaOI71H22pcM
jpuflUv9QcHIdpcH0N0Q+j6S64G9hBGW5pBr5lJe1UtB1lyS4q7I2akNPmNrc2va
IWuymYqz4Cbh7nsrb6KpNts3TShOkPCx1nMTZ4X+3UMSeyv4TyCFf+QeULw2InBW
JhZk66GTqGwHoQCZGzCd+VDOA2+gzivvGVeI0JHsg/Jd2KmfZG+WJi25WxgWEj4T
VtArWA2uPZZPvInA+jqYMZHsDS6Vyc0Qk/IeCCAqFk5rSzLJ//g6rlHUnPRocMt5
W4qnfwjHv48fka8fDImxWc0DioxhsyCeV+IrDFSnnNtP2DkSerSbAMhn7gE5hp4e
8WJ+b9o7iADnAQyWexlUdGDCDiz4zoAsyY5toNpWKpwmMGPcI25wldtGyBxIlvma
SkW853C2PupAMb7GosEx5Qa8h9eQx8zme+EdNCE8u5uRWToHD+PzC2fSsY0KbDCo
YtMfYha8/5ztuoGv+2gcRX9y05iWZHynSlMp65ofz3a+Rt8ZTMsk+ej8cz7DLu5b
h76rLYg5SK532a2x79KK2ASEf/uNB3o1puSl5KvfdkHm17wMK6Q78OFsfSDbkTN/
dt/fmsk/ySwtGJNkkHwofXrJJNoTib5ISLShEZpVzFrT0lIJ3TH1+/RoYUyoLS2i
+j9zr98iyWWq2yEvNuzSILjVWcH98Z2bq+4KnxDp162rWZcquyYmE8mptT6v0P4H
z7V13Ix9bDg5kyzV+hyPiq2K5V6e7iVkKzplO+rSsVSbmTmu/rWSMYmfyUM2utpe
BszAmJsFatJQLgtDMnT3Ou9SLex3MkVDEBBaZBeLEmHyQRxG4J1H342Il/EY01od
otqhy/VbKEI2HGP2KR8Sz134/bQDiLuXD+oGenQs0t2PslHyrWMekgiw38HK0e5l
7hzza6aiGZjYhOfH3HA/4nSeYWpiIWSXdySmI75t4A4roO74i1twAra97ohcoB63
uOepTl5+NcqnRrKKT5e4OcUFJCLva5ne4F62yWzOrzRB0qyFhvg/BXImL1hlsl7/
7Li7TgWXTk1Lfgmvoyet4lvMd98eaIkFA1OGFND8bZbmzu05CW5kc9zDFOweMBwa
LYJXvMu0lUfrUm467Sh6a7CsNTSyLKy02aLLq2OZ1RDOUGCFBWxCYU5f57yCosIS
WjMo0gGKnYy2iT2WOdV8ZnT6lKGQQKGkck5ojYUbRWfwpqnHUbwPDbn4IaDbMcLc
Z+I68+e4eKhNPFGAyE3neUSFEcQPMtTnO+Dkbf6OM9ZjlGx6r9veM6/2ukhZHd6Y
8rMxBAUyvNKqssmH5EaQhfZ/IELZQ7SeRLINoPHnySJz43+HZHIhQRyBmwwJ4xyc
ka3rW+Gs0ndkW1NL9kGuDQU4eIIJlOnxM4tPmyuEah/Im87eo/36z0hI9nk4WgrK
Qr7WtRix0bkHt2Jxo3caIYJVeT1HVGbfhR2Qh9ClmT79IaIdy8l8LZrcM3AuEAOe
xVjHX3OOAtWRzPC9nQWt2uh7CfCyQ5tgUQ9rtHLQf9QFD42D4hdrbe5AxTrUhZez
rWRu8wiSaXXKHZDDdAWGWkni2505497L3Ez3CoDVb55uVq2VQwMAYHKz5a1fm6A3
fN2Cr4v3DUvTw04/CUDjX5Bcmk1I6Z+7WrgnvLfDf3pEV8G9zTcc8fNPjDK4kqkl
UQ9MxMYqGAYThtw9pNA4Ijcku3CijJ+mtdR+oyQd6ooKFUxPIRMdM0HpF5fnvFXf
95rzfhqgYCrbm30wkwagCEhf3oKf2wnZ2JpDJxr668LEWizRAJeq6gbO90M0Vmgj
44Ab/RjVU/7owg3/dHSzX5MV1fh/R77iaUioCE6SuovrYBlAoQcDW2d6+BFvT9ly
HFqkOBh7J+Z+5QRac/hp/Ax93EsFxYu409YPoLb3BuX6/jeuUTk5zO69pu1cpFjn
TXSWMz4h2KS/+QS06Cc4c8E2eLKioFc7Ok3wjsf0PXJKDLxHjpNjbUF4DkL5aNSq
GFauVcWpIap1Q7CBh0yjviHfPGuLrvhH36uRZLRMBXoSqUSbS2nHWMkmDYL6zKzP
+5gwVQaSAlj9xuHCqCP2UdP1Ihuxw9oxLa0i7ZCkCGJ5cKhxFBJCFGT2+mT3JkmJ
DLn9VdheTdBJJK02s53NJC+VbmlO8iEqMoezgXTgkFYJmY606F3rDa1wMiYawfVC
vbhv3L5xwx4xdDPwO3JUu5P1RZLL621lqagl2BApemuYzyR4i9FOIGuo9x26E+hX
6ukT6zC/+T4Mz4Rj3l6eM29zlJhFUr7XGIBpbVHvyC2knHE/kE/vx1J53ffubCJb
X7ZsVeh4/YjfzLZphJpK34isXVdaoM6LUSndjh+4FZg1+Q0OE9ghwkBT927Y/BfG
fL1f64Uxxtzd8bS2i2K0jLfM7Fk5oSAO6XaBaMNCjSXBPMhMFcYK87Jteeo8Jhck
98n351YGnWij7HaOzV4pI68TrKCwuhBwcjibgwP1o0NAtwCbV4buaVijNtw8c5PP
RO3pZ7VvGLOxRQUkTA0UqmZS1V2rxgerBQ3w5T2QoNUFJBQhtZUdKko2X9sXr22z
SwklL3KSl1/L9kx7W9Q/jxyDc021ZaddrpqdAngeN/A66TVFAZ9d8C4R3CjTiJrX
JI5VY4qiUd4c5xRGr11LyOje3HjG1W/5GR4mX/qmmBJDUv56vAEttpH+qTMkkI9s
PeF1L98q6iMik0xdxpW4g5gfIKSHf7fsJ4K4Upv4KM8MTHvOZqqB4HY1LMXugrzB
dJSGEEUOHGNx9WssgMR4xJKmUmj4WL4/oa3H8DX1aAh/sUeii+ZRe5EH2n1Uocqv
70pU/HzySeTk4A40jdfzgc1T5g+8wH3Jdr06fTz5Car/mEFqlOFMTvkhEGN17zXl
jxP4Dny4pyywPGGa9MjD1Efr+VYPldUgUUqjHkUFHS7qqRxIeQfAqqaemBXAib3z
vSt+lcY4dnDo85iyRhFIPXFGlV3eEVqhqNfET0uSLQVQzWqZmfdu5gGZyGd1A2xk
0Ogv/vAv1aCXbDRH4KT481KTVJFNXc5CxdmPPUc8750x+uBBxeJP/vSo6Gpz4CJF
JLzsLSWy6H4sBwlLxSmYerv8IP9rjm2BI/1qQwmB1jiuSBCBhAOeo1SC+rjN2zJ2
Vhq7oXLkSdu+oD/a46MZ5y6hnQfu+/b3TG7yzPYQXLJZdvBLTMx07kDCMSOXQJM3
jBGuHq1oja3TYlgarp1I1NW3dz1wuOglrBx4+voNjEV4MBm1FOdyyM2uQcqAT7q4
mq0CyRYwweqgqGURuTKEG1tZiMVblbwUGg+c0RbdLZNHJt9T1m9Smr5v3FXSM17f
v5tpfOhu0ozaHIumsRDexqOCKapiKPTAydoqNoF5IK7GPexkuxiTYDVti3gj9Evd
YHPqkyrQ835V9sejmg0r1BVTiMlBxUn55VKWMrYzOVSP1KnlHH6GImbhqLm06Kbw
myJw2DMh5d2x0poFlZX3kDiX+xqDQahvkoYyY2lk44Od/yxV2n+MCBQJutkDM7zT
odAsC+M+UqOBAaxGgAj2fun5iKtvaF3NJwNA0YRsLuBHnq1dcfjva19H8d34e5J5
kZ3kIl6rzt2BYqEDcDfI0J8iabH0jnwMF+qLDfu3xc87ruxtb7iv9N4YvkiUOk01
pRSDnNYhEEWczGEqkwPyEn3E1bojmw4rh++5A+cxMYuFEnyTDKWZWEGozeo8fphW
N0BQwDEtvCUcq34fxEYbYpzW+OM2065fDaU5PMZMXD6CwmfFeHv5Z5uOxpRENsQP
IgPwT1nUmF51G00+RHHQrgayth/ylw36Bib2R/hJaTkHnyNhVbtrtIYYJUx7KSqg
PuZ0Sg9aXFX85NOGfjjcvMiZUPDWD7vVSPeBs1smehsVpn86HFL2HLNuEqCqsUhK
4V45EB1kE/V2ICquJDDFzYYUIzYkGZ2IVEkkkF8p9WDirdFbQp+28wZh4ZcFTEZD
a8Tj9vLqV0sdynkFFTGk+2+lTJmaJWKQTZ/AqMDNG6YQAHJA9x999MTHk2iDOg+b
cYXcUGoeF3l8XcsqdGVm8bOuD4XPerolrK3PfDPKLkrOPL/FPiy4lx0LMjDqNonM
YtvZmMC+CfWEMiU7shaGojpwBbAf82b9VDfwKy0/+denpaSlVLStllIwlvNOINdL
TGH9RYmvaCX/+L8RrSi43UJFshUAYEs5fDk5n7lRqWKgF/vK39p2S+BLllfALohl
98GWLpBQb14YIjKVTNy1S0isH+Cn6IB6dO6f5WlhNI1T9tJxzefMGMVJ83VRgxM6
LpfyxTUdTNapOhG3io5mmF3jHDafGGoJTC9AmSUcrgJjwqL7sj+YSVHQ7RLiHLTP
vjTGtwhHfaIYm98eOHeSFNskdkFYYqRc4JaVM0zFgLgKkVVewfbXSQI6toTurk3d
nNUimoyrEwW9MbwkX41RblwpQyl9DsGQyS8AOuxTYj3tHAXX/q1d3MWXqNP7JqMY
SWFQ5jbf6jWRO/SZmKjfjDg1iXCQe1DWRrZoGylPyVFTwQOfumG4laOJ3jA6Rbm+
bC2hddF1WY2mk4lx14heYS2mxHAVaPK5s6VXFuCFN2ciJpF5ZDvgCfiLP/d8nC2Q
FV7Pih+S8PigRRk/w6Mq0cELGzrCBdu+Svy41+ExbgOp2+fKN7iborfIg43eocN0
jKfjIF0gDehZ6jI+xppjHMIKLIaP+T7sdiWMTNRsRgdpXmZtxq+1cbfAikCrQQ//
ZujENkCZYMi9kfV2DLf89R11LEAI/P1u1e7qOx2ED+kY9AhwyBtwgEqOusrGJ/HM
ejtaL2ElxxdEh8NClQhYMQT/HZqDqwh5dniSNlKbB9O7LMCsQdkx5pzZY/3hWPd6
dGNBNARyFh7XyohK1TQTzS0/SBo8lks4rlkfiqpR/5Kmc4pQRmIieVbnKg0l7H8m
R/ms72VCfN4lB9k2yCV0iwD7j23qiPtsZBwrbkHEe/gjAUHkGym77nB+ju+IyQ0y
aeyGFI1Hzbvqm8zRi3QQA68rgpG2TWEkzSbY0o1+Tv4ReVqomCmg5aASXyYaDtGK
+pDIsNatLQ2aV5zi57AHsODjwYqH7Xx80YqkYzeCMrs7AMcEgUMEsbM7pav7d+zG
8ga1sxtgsB7RhOVcrQV2rtaoTtbE4CsyCAJHsCEP5fZOYagiDrcYMnJrz0OTrRp2
ObWHjF/f5bPhYt8pThHQZ9MXnGsT5xvbXQ6F6b3BN9FyeHm7KKc+6zlD0O7qtqYk
uaPn9xSeUtLBUzlNxMaOYNGH1GI3yueodPZBV7iYnaf5GnDW6DGDY3EPsjUO46UE
5L8vrsbDm8kAUOQ6okEXmHf5vyw4XdKCcOi0s+ivAe15x9/+Pc48brKc5UXTd+e6
W3Q1g7D4Ls9aGlqgTEbxUQDpubb3dot+uvk/9112BRWRcSNQ+AhJhPsogkEGJtIf
Po7U9xmH9iyaWFTHq9k5e8y+JSIyFcSx0QbV7P/9hxWPbU+/umnti/TJKSbhBSlb
yCk6lRujwb79OrVI3bzFm9WfAsKXhvn9HdLdh0qiyQP47THlwGFU3aKd6BWtn9T3
VZ+F0raXMVxCdGRv+z9fMgHlLFeTLQ/YMc0+i41/3qnj0UE9140BsOUlw50f4Bmh
JMn2rfeJUBdWVXHx6P58k5OIcrfNhP11LRJh0uP4fut8Zek72mfDbzDf5yP6jLqI
7mTk4csz1okvoiFGwkU99y9qRtosbEWN3SUxXiR3cCdlQG1qSNel2QlrRJPfBVPq
+K7PvxlXIdyx46Klm64ZbyfQAtVtGyXkDHeP6/nG9MGApWPK+L7e4/ebc9H7UJ61
0eCVD9qjW7AbAjT6whkfBLZEWB/yhhwXHwks57abQTC8wmMFDAphvIWwRL9MHD3f
dq4YyTjIG/vkzUSRGTqsfGonYPAFNlme/x4Hegu520DVWpDBBWd8InbFstLf00mw
xBgy4kBD5DAG6dP7vVfGkriyxiqjHlvl73f9oNYkWu4effu3JNSI5Rn+Kpkudpap
PIVtygPLrkWQi+8ON1pgoHrlPJj+24ECWxlQbx0Z8Z7C/lVEbeF48IAI6Jjz4BTN
mPMyLZwnnhSpQ8SKge9AeRzUVGJqxcdWV07HdjTsB5/yO6LdXQ05K79ngBPRRQnK
9I4SrdezbIu2E924Xn2L/qn4V9P2tbVQKMHG3YQqyHpFxFFrn25FJu3s2GqMkPbp
QsutaeJy9XvQLiUUd91EDFh3o8kM3+GVBM+zr0o44pqFTuAt7D+icT2rcXzxK7bA
d5u9qDNiZkDnr5Q4r9ba4ZjUPuFpPiOJaI9BRo3TjkzClnKHPqNYCg1ILR8mxYMN
njvhEGrcDT/Hocsu0tqlO3UCun3pN1soKMErsc7ZF9tEtGl2ul1yWlFW5DPRA0Pt
2uMwSrCd85vQ5475GS9OOlIFZ35Thd8Fy/jcKlCnKUI4QuENSQxGRarrFybERGqv
paoRd6ijfIX2ny4m/5DAI/FVIpS2lGaGsLf8tR88dieRL5bNumHbcohF+4Tb69OM
kmdd+/AMzOMa/zuO3My6SmYdLbuOtcjvIMavkq2eD4Zj360a9d+ewgiDh851m+eE
Tzszk7j+bxXa6MumNQMJA1qBCqm3I3knoJ2Txf3O6eeW2p9ewkyqfjpIrK9TyDMO
ZLI9d2mXlbMGb1rHXFyc++DShCua5fagO5Sq1APHBpog0TMx2Y7P8Jt3CQcJGpot
uw1rmqTps8/Jc35temmgnckWzThv2Ecxe0MqopH/trWKsHi9HVNPVzcSdKuEaa+G
qOhBlUMpol9lf33Lvt3nDcF/eBfl02tDZgjzK9QhdjB/e3Vz14P8nMPjEqTNIKLd
/aDzF/ucanFZXPIK4PFc/+liWw2ivChRrNMI0c475GLLjRyx6YWNVH9uxV0Auh0o
0+SGQ9aVse0uARX5JhszGPc1YMvkS45LnKqZY+Db4fpkrp6OWIpExGz2otTjo6TB
3Pq7rXSDiTuLPwmOOWLVCLvZrLuUUzUBNrcY6bGpb0cpGXl8+KEp3cEEyz5tErWD
r9dcgOpmxZt+9f/+l2WbhpNy58ycuhNEJvCUvR8dish/iTrEWYGdl1uSkkKBWbtT
fv1dLhrS38UGDbCl3N3reYDem0lHwRBniB1PFo4tLxVkw++SdBwfzUniSqaZtvjq
Obug3Nt9DCvjmnOeKMzc9zko0Ibu6gePDX1CXDaRNlEw6aF88S32VB8IlRhn5EcE
OPuyDKJiSZBW3C+XhgD93VW2VP7eezYLBCHoZ/YyjRTbOACMCM0XE+RhWCK4yqSq
axAZczfhRYok5q7FsFYkFclHzSqLKpAw95u+q+8/hNsQz0P1cKQz4ctnZnSXso4H
m4YLByEB9pUtJDBhqykp0UELSirnQK45nKH8vSG7yiHwQ9+dbZu9usTbHqRKHqrt
A4suGhmTFaNjHJ8GOQPUGd9WGv9Pt9HT04HK4jrXMgWcevURD0PhNygrpSwWHfai
pfchf3C4w3ynNHz+PpkJE9F6gaFY3vCnqauOTrxh+3hzS2jXv5d9JajFgrLyX/fL
M9VM9Da7GqHgBlQwQ5zMibBAWaRzR8zREMcI2yMncn8+L2WiDhzNfEKpC0cEodFb
oOuFKn9FGrsaLwqbpRVsu6DHqbVbOCoSuFO/jQIv6Xr0D/UQCmC0FgSqdY2CUqqS
r6u3CwwknBVi9j0WM2QN5MuhAFeH6pfok8mk9Ufh7fl70Kpkq5CdHjtpo6L5Ceff
S/VWvRZ9gdNjb8P8ESY0OKkuNaBen5jXpRZYyAQDVMAArKHZR6e284mEQYuJ/C8D
N2p5UXq5txzAP9FfxSFlyaaLu9VuqoCNwBx/CmqOOErkOOArEC49QP9uLMekjXo+
TQNbOVSFSPgK1mCV45VM1ixPFbXM+l4dfrSOJadmRJmuvZShyxmyQh4PuPGrIpND
og6k0R8zWktoOvI3ejJH6qXLUsbZNtRK0+Esc/SjCOizJNZrvEGLkArkkcYhLNuX
81vXJYF++o/sW+and7Q2he7emsHfa/ajRS/dsgvsJyVOF4stql5M1rkY+zuYXLse
FXQdEko13iXFH7hlzvJ9GMPWx3Eo13W5N/5+s7rBWULRcGK27nQg9tfbmvnYFJh3
AFNO5UPBW55w/mGkyTX8efo3Zh1ZQt1lPQA/VnIgrgr+4WavRt6KXwtLBJv0Herh
BLagAeSEnNuuxJT+R34i9GG7UmxSCUv7ADFb0slv99fp8VDQEPjdDc8OU31CoymL
loOJvjqBSnqdxY/+E1pJljgONuD/yOdyZ8AeILjCWRbxn/qQirwO2MtNUFaaLJ/W
sS7CCQtCOL/3dOdT1fMDppzjrTs98UCz55dfC3CjOuk04yqb3h+kpm7uoQ1Y3HSU
vEiluO5hPPrlcttMprDz0EuUT0bMuTcecetVEoEw9yVbWn23sVTOPmI89GUykZIy
0KkuWNjzv+kjz/vuL95pLC4M2KFsomzejP9vckt7XLPH5xUkBS5HhS39f+b/e4mW
ODyZT+QdSTqUKpI8vErzOFtYUcpiUQL67aknvUcJKoRdXJiDG2Ew9b2G/VUbinLf
gbye8zyoecv9Jk34nyFpjD/HcElW1vsVn0491JBB8ULoLdsbWDSrHGWUownbDkeF
RrX2pUPdI5vIZM1WjFe3zczLdE80uf9Z72mxqkm3rPb6MQaIP3e+LvewU4c6I4Au
udRPEIf6Z6hA8JErQyKjTFBw1laUcei2F5oARF7HXPAJ77RUapsxjI30BXJVeA3s
yJkdPRZgjT8GYSYOglhAE70MM8+CWFkltycgEfFxqBFtQ/vOU8JbfvXWodgo4gUt
XBvU7zFI9fGmmOfGT7QcvKQK/LKG8tFDAE/VuY2rma9R6KQE+n6Z6+z/ACRqPzBB
yNHlqKPvzxv5oacWbX0ESojQPras1LolfkEDZOwgBJMIcnVO3ThoMwjJpEipDDnW
EalDHWiugJminGt0ORiz9NTiK7+SW6WThdIB90w+pd5vfXmInFEhQhy4Fb5JX4st
hDRZspbzv9RLfeEolJCz91KIpYbEMksQkHJr3TnWqTOaHUcwKCCkzwhdJ7xBSqqE
m8qh5pu2Yc4JeluJN3CgIq1eSKUhmZA9u5FwaklfDNVskkWPRzSq2kLjZftdOwfR
zX/NIaB3VAnE9ls93RdwoGti0adayC+0C+7uxRTOZRvQF50D1WXYA5hzX7nfjOKl
r4n6Ae75NjPR1UCvfsGk026kZv7Di9FKiHZWhWb85Ky+mK/tSx+alWdAICQoh1Wg
kurHnWKxGqXPrZvc+rM8p89FCHuUYpbYmvw/BPpr8Nu7S5znmDOosiP29aqGwQqG
/Gkx9o9JVrmVRtwe4cVbH5N04Uh/EVMFE/6pGFeQek0q6RGFONN7vADsuv15DcJ2
hb5ex9r1R/uRuom2LTBJWdLcuskEFTQX9j9BHQ7INIJWv04X5dUvGZRFN+WS12Mh
Yi8j2bco6riWUQQvgs+HbwqEZi0TZ2C4rEGogulbU6QdMLr4V5YqsXPdoXvShHf+
OysKzU/dXL85Bip0b4ug/f3kWRCwrUfB3DZgWkXMFEBnQqTnUMbHCARgzbkUDO1h
+S6pKxM2e5nJKyWBVIJknwkF+a6QX/mGslXVh/jLZRbSlBRnzNZ7r+GZpA+EDcFw
jLxmUaQFc/K9g2r4yg2zDnwOTmVHbBjdu3gp+QYKT0j//DnQ22tBfGlDz0LEat4h
80ELJbtE3qDjRaJsm+Ku2B6lxKRQIkuNA33x0RiMwv1FiYOsmLtbxaihHE8Xue0X
GWBYydVVA4phbcwu7CknslthcMD0TOLf3zILEEote9MKNII1Q5+luE/Y0JpdsD6N
64JBAxw27e6dZ2RM1k8qZJ4outf0XhfwKCKeFu0xdNEvB8orP8exVpwrSY4FlV9v
vKSPjc/YGs5YyqblsVbDfb7zcZOf6MtXmsPtqrg1azTNep6Iquyp+HLb2QZApLva
aCXBf8xbuXejplYGCHSirHe9vHTOzchea3VV38ejqW57In9l1fHMgc3bGhTlt7cp
tL7yuPnoT/6xcogOPGAdu8ea7dPi5oJeylxu4eP4GKs+QyFTUIZd/znAhuKUC47R
qSD4aup5f+LTMMNfc4HwnirjzR7QJVgI3NMGI8qwJvRoOcwrYkvpmJg0HefISlBp
pE4oK0bQz6IrrY52+k/WfY4RmgnjmgiTT2wl487VhC6IthL3lLzOltcPXMaMBbr7
5KaMQcAppCYDJm3Nqgr1irGlHM39wqbddf/Jba6NFUiqHjrd6hfhUDz3kc+6l89T
M8pxcLaqWG5YzXKt6OrnJPqkeJLxe0GGmkxIma9AREq0K3mTalq3ifNIUgwehoQz
+yBoj4BCw0TFCreINwvi0zhcVmtJBmKl3ZoKcYAxg0pTtI13y8XqODsAhyp72E4Z
y4aA4qU0Yhvc3EP+uANxEKbTGr4U4++8/90ymKMOPAHZ/b5y+IKwVunIEcAQCrUA
mYlbIynLlYcXggG1K3qNVDFOrBhdhFCu2PupXm0SN68cW5VwHQem6az0mL5XWPe2
SG6lMUcB3/U/eEecq82NOqic9WZlvfsyglw8rENjlIwfKlYrWO64fJ3JLkh0A35p
clwE1aAp+kqWRxUUCwCZQ10FFo9En6iBufdi6up4QQDlNMWg4GiuLhq8D5IqNDRm
3gdgncs/I4iyJixDQ8mBFMBTIHaMDHRtMNGDkWvg6OaTNZXvhL1n9ZWl/OXWvaRF
7PAOlY3J7ks2fZGnVT1Y5kRcx3wy+qDPFZaQWDdF9LR0GlPcHxY+8HfYUHJ56kfD
G4AZS1zSaFqp+58NExG4CIZUtM1bwnsMe0zYz9kC2grg/LUVsuI+vNfK6i59cDqY
Mns9bg4VEZKsY9y6+vX3pFSEtuiWVH/1iIGxHBcNZZIWgj258f0fMRtyZpc2RgOy
0u7nCLq6M8MRrcRjighzBEQEwyWfoRigs8C00+G+cuAr7SJ0kyV64mbQRlq0RNk8
Nqby1WdyGdveZoLWSkJ66zBBSLY/X8qj4CaUE0AsOGeeYA1q8ONAC0ERhWtLyMSC
tffLmP7rdzH1IT5qzTCBht42+Uvs3FIzqFXXAX3RjojW+HDTpW4VOlt9UA2SNKSp
QAODPoEMq2BOeOJP+RcD7XhbM/PXcLVnfuYIqyhUmZXKlB2kfNFfz1sfXVq8GTTz
u5vNKTuLhDmniAdTsP+fcE1XPcLmbPQKERX8S/IRaHqYW4FtTUNp6tPxJfYYi66x
mUXYE5H0M6zV/S572yrxBEgBRDxY5DohnzUSxEhgJQ8AcxoFm1xosjkitYaJesjG
mHYBEcELT73lwtbvBv7o+JyyBu3TaZyjU/UA19MTEoZXGtpWSbW0WClDQYid/cwO
UQQgQ+YsPNJtVVbi4XI23ryXhi2JaUSZinTy1Ou/4WeaLpAA5ZzW9qMuP0Su+Hbn
eYelCG27djZUhwIt0r2+aP8vACz4h/SjSQu/HewURQ9bv6kU89M5Iut1X15Mtz/6
vYUrfWT0CdpJsLimiFt+3JbIbD5QCoaqx3nK4DKjj6kp2DVq8wR1HJj805r0IYMP
0wbUK/PE5mi7d8UOvsRUdWKgF3CjOIsl0nrpIRXdtKso2TZCWNOgJa9xXuOHgcmi
VzTblxtPlhw4/coZlBk4Z1VAnBhw39ojYbeizeUqfj1/LxDentToUSl03+9qq2Ou
2WVOb5Y72e8D1whOm/Ntl4S+m5TSTRS1RMyZhtZhGgULusjxl49vzFHMNXN6sj+c
se0blIRh6gt/szltJq33ECrWluqbc6aR4E9o/8qWd9Tv7OiZPFZDad9uRz4z8dtH
EnT7GfwkKy+qXyalUT2OJZSB6BmXNIOvsTXLvJReLnR1Z7uBz2ZM92fF3B5HK7I1
Xd20FF2QXLCMIN9KDF6YysIh2GeAAj/e/a8mWYJSMv51OIF90M914+Nijmna9OXy
g0ZkFbyVwaGXnM2SebcD5IV+nqm/X6k+krzjiSqP6MoDuwu4rGefsu4UKhPnt/Su
3UabEXZQNErHSNkPsLhw4zewNSz3G6E6Gndf8/09REGoDDLBL894D2KEmIzv6GO5
9A5uCPNu0huK9RxsYCWabit8WYIDflLtx/MhmxpKueC9o9OC2ZBPBa4WHduEzm8l
OBpCY7HVdZ3SgoxATKvte8gCVVzceEPZwmwIHz8u40gtgVmMyPGSOiMIbGxq1qC/
m96SMW3eiHLm0vR4+fwHsLVkzH+T/Xqh5kt1X/TQ7bD9uuVrg6bcFSk2vtGOcAY4
faZ4GHJll/6YbCcQg/fJcz2TS15efe/UTWa7TXvb6VeS4b9iQpCoEWb3ungcBbGH
9sa9tB20+jGDUBnI5PVg2c0qBKaZpUWS4NG7IRLpc/F6YTAITWLAkIZRV67p3sFt
eJAKXvMieMvmMhnO+l8cDMMlxIHCdg1U1g3T+W5fBaNPC7nbRGxZsoJEheNyAV6u
vJ7/W21ehvTdRVOYobQd33NETJ2uMRx94YtAHbhIu8peUd33kDeFrjn/n6Bw3dgj
ocXbCsBXvZ7xvY+ZyaZk9I0MSFoWkdDY9AZCGdF9g5eFmLBsylfKoCkzkOgQ7h2T
/uSPljdT43+eZrgrx87+7hT3DYnoNBKXy3ZspzOprY17FPFGcRy5zjf4tZbdMh35
1JxmmgFT8eeOwjr4HVB+tTb7/hSGH7u1bRI8WEuSA+iieKd863I/CO/IhOQG5DOe
rdd3T7qSRO8PrI2tzRekbxsvxqvuzD7mfK/keL8tNr77YacmpW6Pdu6+Q7Ld45xR
GQ1xcOGq/LjVsUJ+D+rzHztrWauT/HOFPXPXmD4uT8+7gH3OR5JAjmrO/IenrbbY
pZ2Cgdu5CX0z0qc+FXIQXpRqHPiPYvQkKOHkUdeuS0OhkgO5A5KFKNq+EQTXTXsF
C2X/B6UYL4yBapHr5N9TiN+dqFauAgWzogt/3XkmKe94t39v5rPer0WJBl8TUTcn
oiE8w08QC/CKOaNGgKbfyTCF4lBJqyGL9/EPiOaotUJR427SFkjIhqPXP/rMGA53
V5XEiV+ubqUfwNDWPhKJdnzH/H7L3JFwYVOf+3EXwsZ3FbD+q+c41K1z6X2zUm1a
wIbEzDZ2XCdS5qVeu4oFWiR9ITa/+BVKcYvNyjD00KgwNYmrjb84buhRJQtgGp7s
x5wOS+FTiOrCW8gOsMZVBKmbbd+niBYdc8OnDFkOPs8uz6anaJrquk8RjJpvKdS5
vtefeaR59uY6wk3BYutzMsLWo1SxvaMMCC5AI4SdJlP3W62qZcdv0qwYqNo4uVol
lUeSLY6sEsAfuKpu65Ly/K1ogTJqADXXgh/Ol+ezLtbRW0QV3G5iL4WfJnVX8X/M
x0qMDjQN8t9b4NOyg+3hEIYEU2vZEGFWJYTe59ub1kikok1+7Xh/3Vhlg6lvm62o
hGDk4TWEw16q0DEG9XzENsrT+TsDSxZcbmSJansBXiK4HDJpvPDTsAqm9kzEVlc2
pCGoPIGGLVOcyhipyJ5Q1eI8TWimmD009pMOc9Ffa/kYcc6dP6na6vgVLLRlmOa4
ha4S4ByiuId4YLUWEoD2arv1mFqzVNX+F8KhDDkCg3iBjISeQq2xvfJafjt8f74I
SogQFsJfgZwZYBo2zRqKj+X5KcjFCmqd/3iDkZLW7dCe8Bp3QNjHT3taCk0CZKUW
PRteRjk3Z9Hb0h9OO1QIJu/vMtNCAVhRw2Mq+UiSgN/8mAZXlL9ZgYsF/LXosAGa
yiFCawZP1wWnX0/NMuoVXFQHCdktw74AJLqUYE13UDeuFRtzgLwc6iYDLQmVAUDh
VAHL/gSkrkaHcMTW28otWImcHekg71Qqwxb/4NRkPrG2ZyA04CNcGs9capbypjCx
hjrho14Ql4QBH6wql3Nw+pqQr4jYBxqLbzR0aJP3e0n/0TY4sjarUqKfM0vj4qON
+sQfqkGi9xDvmiQZMo7qQK2D8EPpNjW5rXAP49eH+7jAN6WwYqYoeqxqGb05gybm
s+1sj+5hGQRWffjTPhdV69YEWgM+/PQQRNv5dBO0rm/bTHf/J24F0lhGyJFUZH6z
AtERmHFaqVoRzXYQWCFV6XFj825b8AhXj2u/VOgM0nbQasTqnwePU7qWQIbmNuoY
oRIQ/a4uc63UR2ZscUyDVNp8BBOYVXjNVNkmk2Hopk9tG5Kjrpmg69WQM0By/K5B
XrFThflPJ9ot8zfMOqDF0IDtRRlN0a6qDLlFVgm8g9Z8NcEnoWireEIdB//OH82v
QW7B2l/Wki46S/ZLPWl11PlMTgNbyw86ZliZ0YiMdyOBkle96oK5xwUzpv4RjYWW
1sjJXwQKRmKaV9V26We7LNTJ+f2K6GVV9k+xGYVNhkB01CKmyHRw8C8zIV1I5/P/
yQiJV4l+ku1nuORxvdY5ElXr859m+7edvtor3765YfBR6/2mn0bRuwtG7kPz08T1
Yha/QkH2oq5Xona3tqxmH3GkNi8FI6JUKf1RS58WiLW+MkKaAe/f767LP+JVRBZ/
t+6628RkZwLIYYU+Mr31Ezus7FHSrt2WH8JvJO3E0A18y5ts0fkme/x9O6Xa1neu
3ZVl12dJxfzS3jELy6tDduHec97j65s4kO/M81OJN2M2uY40UTabz+zVB6jBC63q
BTKcRLB3i++9OS5OMeCnb2A/V39a2Bl+16hvrdpxPOu0pqHOQkmXkc8z+kB9hCUi
Zc+EoPRD/yLOpjde11rvQezfH5rsmvz0uKuAU2eNpJO27giVz2IwCz9udKeALRdT
orPQswlDpfcJ/Q9z4JidIvF7wckcQPQ7LmxPCi9oYq+6aavGVcGjJ+0ZkT+jAIxd
BeJQcPL/SV0a/JrUB96/57jACZ4nXAc1K3vXn2utYLQXLE15dIvuJMuvK5gumd/s
ls6/bZ4JD823RgDj2K5pgMyR03iymLCPM/gh/fG+iEhiXibf0r2a//oPsoP81dQW
1+XEVoZCBLOAufOtui4ZucOZBBVpVjHHabam44G+fZ3boQbNyMSbEAelMReUNOce
49fRrKPmcew3dzRbeaXT/IX7Bt3IidJ1sFxGLCrZT7BKVxFzatz9qgpcRk6eRTDD
PD9JjRAbbJTd5SSLapSrTgnHleEp6tHsUmTcXPrwTqOr7phE+UcOciAWv45sVddS
n9TWYY8N1/aT7bMNsxBAug9VKqsz3D+h6AgSPFE/Q/mA74X7i9oJUq8K3CXU9R+/
YMPKtTwk5EQQCOTHpDH0qsfOHbS9mhRSrOlxanahSB21B6RLq61cuc3dsXpzR/5h
8LJ1BX3LD4I7b4t/VpwC23xn9EXa1pE7oT9Yd4q+8bvE/Wlc3L4GInEfqHlGeAIk
DZGIyTw4mB5UJ5t3stpwx9dMCNEqBGK3nVT2fmT4l1gTRuDYRVqsNkVEJauc/QCy
yGUQOl1Xr3g5bx7oxd/oSw9897XfPd3ohzjMF6WZUYQVxWt86ctTtzD5ljAfUEtz
KoZfxGSqqnxpY9h9V7nO/g5vlXH6iv2tnHfqUo435VwSU5hLnHkIkmv6y0o5gTZF
U4zpkqxaC49uMaXNRLdXDSIi/GKNOAFHrCJx4pxSEz4pkOdCnJnMO7K1DJa8sn2M
g+bNfCNCgG3fyLsh1TUhCMvNMj4ZF1OzDx4VF41QVllfbvJzft9gJ/PSHG1qQU8t
k7FdiL5fFz/kJRyvyrPFpm7aJwi45Sd/eqYIUwRMAhqFcUUTV4YFNFG/XQWiAwFY
5K+ksqLvGfLx8v/zm3IUyT/PHSYdGDRNLak3g82PLzlfvHMNWA4vLH/83Zz01mS1
P9Ceq9Zw5W6TWng/+V3jWG/onzFNWxcmAO1kdnKriJs35MFa4Wt8gK7lW/J5J01U
IeWdY2iliPzfnK/MbNDaTM1iil/2YrDAokB1MIOop+JEVEaC3MAPte0vBG38Blqc
stbPG2/4E1nD+JffwyQDqWaN0sZdMCmCeIP+OOwo8/8dR9iid/fn7rLowBSfaOtT
k3C/VV8szlKWz6hw9DhmaIfT62bYfAZc1bRYUYh5sOmA32s8JofyGpxil/+qtF0Q
P9eZaV32Og/elErppbe8TwNuThsprf2+uzYKT56+a6ERWix3ILtUev6iCWU0RyE1
ep3NF5osKB/enNNrXsoOUi623f5UwX1u10DH243zddTo8s5FIm+Laj2vDAkuDpFv
1MtkEgPNiEWi1GikbXFaFTG0zC7N+yIPSn089DW7/v4yXltVbrRkirNsdrxCWvvs
ImA3zExy3W+WzYaRozXms0XbirqjuO9VZ6i8K7J0cL1CngepB6E8wNCT4CACS7kj
mQSVQnC4rML/2+jjLxrWLELGe57Mpq7rYyggu1HCE/CpDZjBD9VKTaPU2OmrxLt7
N3vPhf34mWcbQg3VpazwyqMIP2LAlA0ONlAJ7VN+bufNvIlozCcNZPsoAY2jiQmH
OXgEkXvcLpimIW/gOknzTy29k46ZIDbSypO3nLoaoFVRltkae0u3XquLzPGHh1Hk
CAvyjORVFlNJmwdjWSSaUQ9aYtf+NyIyi6IYA2dsASOji/20Pwj1apt2qrG4sAS4
FoPs3YbUjr3MuyYrkJSt1PAbY49KDj5KD8AdcRGZD+PjiIChk3s7NHyK56Xgp35L
qjmpWQ/Ik/tTFRtTffqWptq8cDa2FdPCZ7w8Op/IIwCUykdUm0qmRGYnk9X+F39U
HjvPrGcjY9/B4bZlVRdraXZ/XpdiRZau6QmeK31ezvaICUVcvD342Ifi+xt1oJ2y
zOvgj7v7UsWpxSyl5SgILTuOnWSLdTtgH1WxGzxN4qn8z4zk4E4nGyiTdSDd5mnJ
HsiBICtTRQ3D6iEtjKzg+Ex69PB9EyDyCf8Epj6JajGYXRVJOVx1bDcGXSi+xoyN
VqR7eK2zSl260Jo5nI+MLewanDJUk2ipWQsIo6+SFFtI5qd0UtPU9u67WVICmKiB
A5I3NeRgfpLBpOY0xWx+PQWPt8CrZh30UNGwRv5GAimUlyNK82iXWHdWixL4xuzp
0kSBW632iSR9pntO9cW7rdK2MwCradWxU1YV91UVdxJt7WeL3j+G6w58C/bkItZP
G5x0aBoGPn20W+iDzTOo0qdLA68NIZen4fcjYJi2WO/9ncml+a/Qjp2FPCgJc0VB
gwmyJzXedPr+1MRgVrUvhsYTCYXxEpe54yTnhChFHh9kczmDrAkNGeSIxyTFylgL
3uJ6yAWXQVwb4hTZagy+QDdLoFAXxB3/F1IM8yJQupRJesM2F5Qo0iF9ySlYGDJD
9hUlk5Sl4O/lcRffKyvug8uPb8SGNxQKoSdEmKiXVL4wpiYxo9UegjOd7FXUviuC
O6mGzcnmBTSjurujVMfr/vn7PZpDOUhnhsot136D1tNPwrgnIs18uKKVU3UiU697
P0WAK18dzzeNCaRpB/K+ugpVOtEDPhMtDgxyXikKt1VYqafCLv6YVWYTKY/0PFRf
s5g4BmZRdUJRBySD5mOuDCi/87Lj25IqMfQeaRyL4ghKh13ClBYm2vYgrZrnfOR4
lo75oIprglV+gS1A2OqW4eD6w8BVNYbZeNQZEWRCQk7huLt+9U22Nx4oGQ6jHWGp
8sT0vBbWHSCk0w77S++iDd4qhrvvpH/Ysh70H4olNV4tGTjixXYBjJVg4fyiDAA5
P5Z1wyFOsTZcVkcRMuD/jAAgM4RB6+Uby6ydVrf1B8gBmwyYTe/+cx4ML7QL4HHU
N56UM93F17YVEkZhuVYdvTfa8pTJ9tjf0FFpaYzCrwdM0NT2R5GHbaxXglbj+IyA
3CBZuNOAeSDDA70b7uHnru83Pf4RXIICXGY5VFabAKR6VRT+LcAco93u7WgtGyF7
sXew+cE6DRQ0xAFBCfhYYLYEb3AwPZRcooNxFB+T7GTuDGXs8Cb9qBRjo2TKOqNq
NPc1lW/LJ1gjUNuVVTJ5cUqTyulM01iMQ3ZkoTwKn4QMtImRSgfBCEbXqg7UdLnk
OkOnUSqRWPmNP2zx7Ylw38P/ocV2qDqXSV48GGipDH3Ll33/d9xPZVmzzbQxFjjD
1Nj87rkW6ga1952S8urNu1XJZa38kzEXfE4wSTRSPXiqto0QX7/DDJ/NXJA9qPMJ
mxcCkSvozX29myhuF3BNY/wAtbYLi3RmeptA9UGbnIw6wydLuBS/HssSzb4oFfLZ
uoNXMMMkho368hWTcXffvzm6htu3dCSsyyvJyZ0f6h/6PctVJAD4QUbJWpI/Dur/
Km2Y1bVyme58ObFJMyR9ys4PB5p2fQGPCVjUSitxtYSwK2VBziMfmypahHktdCaw
b0qXfTyKNXZOmPRvZowGwU3LFtiNDtXMSSxqLOtGM1QeNoI9wf0I8i6sLG2IAwSf
Spt3vZZfF+Wl6g8HiHJo16Swi7SCp3dmhEdoA38v22W/wRvPBRfqvokTMpVuQmzz
VQKJOHT4plTu1mq3fL99zIgKELc0gh96uUql2d5l65UEC4NpiUix//q4eZWhyzfG
K6o5OpG3hYT3dWtBywmSS/5f0lzIEqDAlsvgSYbcNdU8mp/MD0cEjo6S1swxEIM9
pxCo8/AT0p9EdZBhS2Z9a4p1ZE1cmayBD8I/k8wdasZrX3RJ7bTLB8TXG+KUYrHT
72ZDdVIMFtzMJp9/hhEVH3uLNMVE1N3wjrD9xMkJr61zb9t2wN05FQVcZC18JV0Z
HOVNvw+a+yiO5wKW9Rzex1nHn1fHkEArQro5VIi/7ZkR4h1zyaKK6KUEjVOxpNhG
IL9VgLE7A38aEC+s9+3i6O9QYr+dUJ4+HK0/2ipSWcnGJYLIsLkAlAhW4IkLLHvU
J343TuYMbZchgayBMuxP2/Fp87upDkFoz2sKaLIYcSp5KjFX0ETAXDTRZE0EDQXJ
zzZ6s7aNth4rS/RxMGUhNC/4SKyEWT4n7InFu0fKMrfP9OH+zl3iJvpNRf5+XwxF
LzKC713ttHeBo+kPwlfCSqNbdUyEm2zJtdJMYkem0s6juSn/awGDpx1iFj+jgiS6
dh6riMSf4QuB29UvtJd3ACEUzZ6wCRsoGt6XzOVPvO7wOu04qHNosh2/YrP3mwQc
sbO3ne1aJinc7YxlZKY5rJQAGnOpYjX/sTQCx3kqyUBHB5/oE2l+wzKyeU4WOJ/W
QHXWVuv+htG+kP16BUw+ls7lk+8Kd2KzHN6XPqlFkcwqzvwH9ZocG9JArjiJyy7i
anz2MoNMZBLU6f/82Oz2zpOm6iQarAPi3yVAJJz6qLj1LFaCHkHEh731y3jaw7QV
uhbOE8btP8phNjXZwDqOJ4rRmPaCevBF9FHTpJ6cypvd9AFWW2T6Wc+MUOny5EVm
GiwDf/hQt1Q3SIiE3nRaPyDY/Nkzm67NFzSMkuWTNnXFmq/WsbGrQB7ddemJ1MOH
FkX9SU6RW9JwicICbP4KRevQIsif6dWHQ9v4gEQAW7GJDS29PsGXv/EThueOP4Qe
NwSsLq5/NYTMWCKxkPJs9T7eNY2Gcog8NBfR+K00qlzF91AIM2/B27uR1wDv4SVB
pc/QGOk8qO1i5rKksdFHwZUkMSJZMhYTKxX6za8ukZkRg7DzYylB/Wuwxfe2sjdt
axv0e+b68YhjmgS3bZxX9qmxurntVmR1GG0HkomrzHKZ5g0KXFqCPe/4CIuc1SUY
x8dasvau+JzgENq+diH31GOV2JQgzrUjZi6cotAlCV933TTA2MU6THujAlbFTgJh
GMk4Yli+NVHzUGD88SiRInk1VmoaJVDLnJ40TjPmbdIe3T6QSD3RDUoAT6/O1HQ4
f0rh5t8EXz9hAY7Jmu2RFlqGQVkqPl39zWcWAxrAckNChgjLQWifQCeqNdxFWZqP
OyXVv4Cq89IS4juOAWZtCUVCVIBQpH72qvibsDXmEkL6Sp7K8JoqbaZXL8ZhuR46
3280WYOfS9f958j3U8My7IlhKfeZ5ghIdPXWokqsD0Dpw+lkXmt8tWi3TYDTXxAq
sDnJxEPyxOrMUPy/LJtX8LvMcYjfZ9lCeyXxYcGa2Vx/VFdfAb6TJaOVtOSUWCYu
WLQHuU5dd+GI2GK8DuEWMzuqZgJeeysWnpDn2zGxhjkL9jvGL+xDf/lH9kwYIFl6
TdyKz50eNWmysoou5L+2U3lMPefNUTsq8LFHnFtH22OwP0AM2e+q391Dp59A8KUR
NsNEOZc7bbJH3ltYgBFR4BJkSTg0is1JpTXp283iscdvXBEfG2vhYQ6s1ZsiysQG
LxUIPfZpjaZXrvRUl2q1TasrdEI97XmhzejO4Of06Lq/699N7f+YYuwl8hLJoBH9
H3+2mSP2ItzoFeiGGPSOvzsq3JV+dFv7W3a116b4WGg9N5wA63Wyox57MiexEKEP
J8DlqXN2dYpgC1B3vmIvsDYgDPZJnKQ2EV0GAX6MY98mWM4vqlNu/PlttSHtVhRC
8UokadWP1AqfbaBjMyIC1QwBR/vBFba0hrCGL2Opq3DMRshAh5eFYqFE8eiEA73E
2HiknwQ6xhI89DN/kNuNP3RcZaR07e0a1sX5wE/D/roj4fRutu395SMaaBr5zF8G
ihLs2cEUWlXtcV+/1V3aC2ChpyWCvUKh7TS6ZrJyY8DZAtxj5efUmLfhfhS2k1g2
Uz4KbOAi0hxsJ2JrT1Dabwu1VqnTA9YC9cJyRwKKnkEmxKkRuAiYnsI2dbGnYB1n
ZoQBH9lhiOMVdaifG75lIsxdpOIYMZkYr1Otb5hFYSVNWPY0PTlaBePXgzUgJnuZ
Kk4QJ4t8TeqbWCApmWXjG6SG6r7uSvlwEDTT335K6l6EzLZ3G0vzXN94A8TZ+OBL
s8Foh44EtVHJWi5TOExxYX5g3/luJ+9ZQnYOJGgdRFpSjXr/Uf6D0LLG2RmJNB0d
s1vlXoCxUBulLlS+uP5+zLFxD4bPqo0N+GFzIp79AkYeqB34yisl99Ft9hNVdT5J
n3FXOEtsxZc/jXGX7esAX8hlgYOGn3hBAvh3Mn09J/dFJxpfynhYv/csfDfqAjgO
JyO/op8A5pzn25ixca0DCdv3QXrHWDP44WMzG+qVa0TgXlnGHVTAO64vdOew5JXc
9tpNJxbTYxenhGKSSpH7uA6k+8Le5pddOELJX/zAw/4kjeKF6WMyKO7Kzz6CMaHV
/dui3UtWzogp3PdB5WwRMl2gf2+LOFEX8DN0OGHzc4FjQngvMqk9O0VjErzHmvTJ
qmfc0lf6OE8khCoeamulePRMyxzyDFweGwU42toLIXzqdvscgKXmR2cQx05Q4P+h
xt5jm532eBfiIqvRjHw3oQ5UP73xKAnJMxoIBmcf2SKjoDZV897k0gswPgaWr6A7
QzBZ6YoQcTZ2Fek/XAPdsycyW3Iq4v5Be0MBUUW1TSBHBp5xZdUzoF8IiyioOsPX
uGyFSU2e5uIEnlcRW860HmP1yzZRaYALA06AtkC/SuMGpU2tN5ECyL539Xz6FVvd
244BmzXY1f+WOMBymUXBGE8BalVbWSF9NRDvAiOlUwoRJ7ENnGYWNXKJS/cjjvqa
l201PgGddae8Jb1BhiVkSSlsVMr3mP0N0y8ZGlJb/RR4cTEk5y5IBpGwL8CEd+ub
T1/ce/QRFbij9TBPHinPRXcsoDxywRLVkomcJI+hcBv57okWpvjCRp8PLeuSGSeJ
JDqSWaozY/kBEunPUtBGTTfoVJaUnFFIqmUDr6Fz48FCyjFsRfjYQXR4hjp8I1UH
AzKapo9s4DUxpV1VCRds4O2SHMaL+CLz3LkoUHOPVBHm3MePwXfSnmtVhhniki33
0Sd1Z+B4bohHl14ZMoDunv0v7WRsIe39LFIEdcPUY7Nu/78xY24D7QmT1qCvKlwZ
8oCXw7JwmjRzBCMyBr5cFqvVnwZuAVSo+dSBbagnOTDj9f70JtIgfBDuOzeWI5ix
FgZeEJZqlEk3EDTHuBTTxJVEwc8IGmLc8OhxE/fdtDgKdcGEi1nakEJN0PfaFe90
wIDWjl/AdgJ+7xtkJLdN/J5kupUac9u0kLkWqQhST3Wf7x3FjHoNJUgNoXOTsI7e
9Ov2yWABWj3+mP0Q6bFdezsb9VpppPEvItk0znyU/cls2yKMEklIsyyhB2DIpP3H
nAnKQxra81aDYqsarvgvKpaL9nhLd7keZwXbXVcAUrsv/1BC/2FU/ei3RjSaL8AU
wVSPpj0+juuqUwj3Bpdmuydba6kw72yJZbWycPFuOzY7WVbPvtleM0hfxJD/ErmM
lUtcrb4VyZkvCyqkKqCv2wDOfyYIcCj2FswZtL8F/boLY9fk2usITyHd+aaZLIr0
zBLXwsHQiRHPq1Hvq8Ll9WbDgpTYwfsxXC35WEkC9UYJ3GrO5BAHL6tFhumnofbK
U9LJULSRLsd2mzTSytvsMQE2R1t6UqNVsWLmvRhFSmzvB2s/pszG25x27xQK1ePg
8gyKwDDCGO8EpisQt+HyvCvoOMwJz2lKDnEEMHpDicqlSr/l8e+T/JDsgmaaxk8a
NkCI1lHrv6osW1DPM3045I9ASs88lXFVuhpkBtut/rsqUEGSM5/CW4JqS7ZaYu4M
Eeck/qXgglVN7wgSTv4z9ju3hah1HqWdfbBNw1RtzjNTTnDsQ6lK4JKOCJxo6lre
PzgJVYwjug9zTjmHu7+84rbYTovXj7vf8svNDb29WcjaDEr+sG1xrc2n/gWLyTD0
G3AvwOZpfavw5cTBMqeH03tczz4yMJ8shmGmV35+5uvWAgbHaTTU6b3RRQLzzbR1
LHK1eV/fiTFDFhb3Y10S/Zh3cEXjfK5QbsAbGCeEjSdJnuAsFe8Lc44PmNSr40Be
nZhBq17Vjcp8U73WcbCGP4nr1FI3Ennp7+7YAyTOuclD4Ojq/fO9CUZ0LLCGQzPE
JaNEHezSgHVVAoQQgMzYQg2dzAcckaEc+WIJy2Ll3xJ8tvrxHOucQZwUhAsyFE02
UhHfZfPA01Ko6+BjN6R2tnltzyXyoZ8iyGy8yF98SCmp0+rBYe0mcZXkblbI3Jp/
ezLm5oZuP0UHpXgXSYbErp08t+Nmv1UWoxEsaFrjoZZu5ixLCpK1HzcnREQVZvLt
8ba5MRqYA9I73GE4f8tKJWuCR2EcVKdUt8Hr0bBaahqt0XJdKtCRcfcpSvGYO/XY
AA+fHt7PafpyTSqRDGgOI6UDx0KkFjHqrD1K4AqxFj2kjXy6NoyZiozPNg/1pZip
aozrPRIjq1wHMI1WZL6b01WLl6NHrmc/HBvrTUqY3Ja7sjMef+V4LZLi/ZuprPFx
0gqryTHfxT5GVjzheYKxpbw+0/Sq6bSC6ADK3gK1EdP+2Eyf18WkZU5wTpwZltZS
cowNP+pO2uQ10o0hDL7w7aVM/3XrUe4hITpgIapk8jpCWqJpk9iQsWsvSa6mzXVB
/kKVWb6XSuXzPRBprrKICfffO9179Bo1EqjOOYoQ7cWH0ucnvG8b4hHKpBYNGSr5
AlvJ9Wz8/oFlzobvGT1ROheXgIkKIloHpQpq+uL7l1Hk453F5R6TcxiMbEKb2XzK
zcPkUa9TTz76ksWWlglghajYqCeW78nskUcaC+PgKs1ohOmFRrRJ2U4+JHs3szfW
sQ12DAB95p0Gbt8yGZAaJamWmC6uzm+R3h3LyK6lraUIBdoIJ3OQ3DgLekx6S7Tp
UrvD/qwPJmgj9Cb9q/OfQ2lve2rgn9ombGTQVSAM5VxicH4snJBUjkq2+X2AP4Yl
NfGkyYg/hNIh5TNcSykoxhEd2SLOY6Y62dND7MRgNaRMtV/4k7rcH94x0/MBZEej
fvgoMXI3miOCuK9xIc0vLqFWkt2PLyhOkp/JNL9/EXVtX13I8qDHmLE78dLoNoQg
rPF7atAjGC2PBn+kIGkLxEtaoDpgg/KV4jXkKPM08KAkA+LFW5rBmdbMgRKYzQo/
aiMH3YquQExA6YPi3h5QX7U5oXcqHY4OCCo9SRM5gzk8J4QFgH8j5+EcAHLhwJSs
2KXLtSmaCkrBULs361zR4aDIL4oi0k3Hs6zakolpibd0i0XtVg2zEPj9LEx1rNdn
YTLP+GTXv8avNsBFWhII67Gz2N3Q6LEIaQqDQOl5N0S3wKmAKkyEjAP09xSouMBL
6NO8VW1MlSrR2fg/OAfFQA9kW+DNLiORARzTFMZM31Poy3C8eXuuSv+T8+oDc0Hi
dGDRDsyG+lCaFXV6Cbm6mh5gTSdhql6J/DsRiMjj/lzbiyYDAsUHscmdVlnOwU/g
BvtCZEIpzDesSbowd+PAlpPH1YjqQR0Jv+UFAx2PdZzhI5gRpkgIJ/kbrWHPF0Ki
slsdqqhCg8MVcRX6ZKVYaY/kuT7PGdGJY0lHq7varvRC8z43PXqY2Ner7/UDCG7D
cgtDvTWtfAVVjJxk+CIZxAViJ4+sReT/7aEGDSqmFHB//j9WgClzkvfJgjOAvZhC
5Tdo/rSXRqGiSDy0wfrvoFnXF0+bCDT2GM4MXQjqgxCh5flZFsxnRGxmE0ZxRYRw
5vTiFm/CWsFPkgencIBrae8UeEPZNGDFa01UOuPYvJaJx7G/2ebCjJQEnBfDZch1
tlfGDcq+95amaEQub/DdfMVkT3O1TaXzkwrtMdnyp+4kQtBCA4zocezUCjOUGDbH
AsSRF7RbBjeVVEcx2JaazQUUzeNXHBs76cJnMtAsLVCVbmuot55vKVwbOYEkDvFo
w6/eXUVBvlmbdl/zMosCF08nFB3QCQXizAfsilcBp9wD/63+LBKLCv3RS3FhIHhz
7QmkCyMrhtiG9zPZxmZ/2c4Phj1jXzyGHNl4+p91RYAo1O2r9er/lVVcghxpFzI2
susN/ak1v2CK0ZmkHkNlw1hiXbwRn9g4kuWfVyQJl0mo/qmP2hsKPuzZ6qQyhgo4
SScdeQTD4ZPA7CP6l9mlTIpJVlrOIQY5DUX+/2ailtQBkrlBVnImIH1WmewJlc/N
qtSxqSNgywPEECvr4ddVvvNEF1sDLaNbHg7+/BgunFtg/CZ9FXtHwDF0qu4cSBNI
h7GVTwgG/iO3P1FcbGoBV19pNj8U9zMdwlv2m/AK81bywni5cu0zYENlSqejOpIO
+RJHqo2Wt+B1QiPUB/79oAPjYrnLKIen0vLNmB3XxASPZMgrZSz5L3uCd9BSoFci
3bvfLcgaKQmhcPvGsZr1BtJ07nPwX1vYY9GqNhc0u+Jac1h3qJpiopnk+Q2QAoKJ
m8fjhV/SyXZBk0WPAjDevABUQB/DeYUo4ik6eoWAyg59MgFyeteUzQICmTKNZVq/
frl4C1WTLZrtE7ylaq2d76sfIShp7t39kcQjxk0I1FLeY+elKxV9EkCyVZsUpNk/
i2pGgRcc0MM8vSB3g2Qytc0YjxTm/JJf6fwz1TbUn1cCCvj97UvjOW1HtHfHcRYX
Ur+vZAoQJWjK9cSTwiPOCjjM7RxSO8YHvYsKajFovV6sIW6hgHTRlDyX/GNAU2Gy
+kKS+gniKq48v4EerqBYIlJHv1VO4x/kd+qO+U/j2LY2lfSaS+nDNE96UDGbHVMl
srdK94tbn33k54LVLSEm3PZOVAzFbY3s6d+mox71ohFlO+jF2/feQB3/OfWUzoYe
sxuacVkOauaz0P89uxtQINaKVeum3wTTi9VLDmQ1sfaB6OevyhL0zE8HO6lwAOjq
Iti9T2CzHnSVuT9uQx2atPrAGmzt+rb7sv1+0v1YZbiNGzEJona/kOsdbmTWuKh/
986+5TT41k8DtpCxM7PlcyA92FpUZ6x6Aq7n5RqG80ZkgPgj+2eoVSHUg+i0DOOe
lXp8zsbs5GdcP39LretIACWi/EI187NDbbCUVzy1ADuLATBeI8Ym0CBKqpun2WqF
oTVSYJ7F7YvmJ2FB/SlwIZpQSzeWZ2O01oFwkcsw2ShMinXgaCohLHJvqtG8LTa3
xvqiR580m/dw+xI+lA2Cc3wIheGD+BpvuBKTtXlmjmJ0i8mBejs/0Ld3Sk90MFUZ
qAlW2iMvSWw+YQN9419VB0K2FyQTC7eQUfBRWCgsF+ImSL7qFYNAKvf296bTj055
gENyVNvxmOoeC/4upXAdEp8rviXl78f06bF3IjBuvw/UnKwRuI+BEty1z4fTut20
o+qOh8JD2en3xv60ZEh7SFBUt3320rGrpXa6z5OHYS4ToT1dhNDbnunIZT5JDATY
xJemjN7ccwCBN6muiRreqZE1/183L02wxrktdDrIFkH99yNI3a6/vupgT2G5muUl
7tJMW70mh0yz63TrQVwBRECjUEgVb2Jfij59smHgvKhQJw6ZiAKG162DA1G9/ItX
6MDyc6RTb9UklNSJ/j0IwZbuaI+nw1VV1MMquc1/msahNA0fZ/RwOJQjCfWI37KL
6r9fIeHKdm9b6fl89gFXSbmUiifZcsBDhddPTUa5lLwbdubfSihgsuFHsP4Ws+RG
jqb+M6gzX+JtAm73gaGE0E0MmXevpSCI0AzOhpXn/LRf54dU4KGn6/m6euAWaTBe
V89DYFz17urCMc6+5LyXEoPUBcyUkFnuN7JIXRJLtqzgsXPR3BV8ElqpKTN7bFr/
pHa2445SkUrLdsPZ/3wDtKfWkwoWLad2HmO8TkEJBC3oO1Qw1R6V00qatfk0jq0p
bjRfE8nOUIJHvVRXQGm+IFeHkppv+rTHdmpe5gh59qX6pnD6xxb8c4lksdfTWkvh
vueUghmcO9KGEL/Z8EWFM2heBI4tFnStxfnHUX1frIGyKri4Eck2zq0VS3KSJMBu
3MGn/0rGSCMGQFEegXjT3SltpKR5FhJG7NHmTZuFrJdRRlcCPCECuxO95S7csmUK
W18ABy+3ltRj4FkV0OwUqa5gfYG9ZZdwFX9zXyBcS/cun0VSedyBGYU3859yszTI
iihoyRzd/EWgR9fOPPOsul+klMxTNuKMay+sdG9jbpaUrZsCwQLFrJQopltyYnME
UtWS345cQlFQuRZhezijNaH/yK8mWdgkGCSUlpPpJpyFalrtAVgF3zOC3bNsecKG
dvSykNjV5SgvSo3CKgKZHiojXCrcO/lIcczhnJcYeCzC5NdmEDNIi09xfgYLLMkv
ZmcGJad+i4hjlQVlaSjxoAJSenYFmvY3PTMfbbw7qAvQi2d8HsWdDRANT9kPSgOZ
xPYdHBZit/Ka2EfHkS4qPHRXm4PRsE98tdkV5zDXF/QynH/1a+e9/pTHVcdR49Bs
t6diJETsAbr+HR9lzAkHtvxKTf5VTx/V7uvV5ljMBibN8DmHmoFzdFdD7yrEBb5m
4p5FifnsvRRmT4PQGrzcTVnZB0dNPKG1/IU/W0POQhdhTBuucGnaYV7LsU93po8F
noWTjCTy0FP33CK1lmBCbtDDgQmGGZeu33FN0ETirosemzXW74x3dQQVlsNMc5hp
bMiuUYNo6XZHqS93GwotJK8AvXscw2fafBwBNp/JCreMlsq7BRCRIetT/LDZbQXb
4+ZCHl9tunVYkVltRXi2/D3PQiHbMymnyzA5L9l4fEL6n/delaR2mxxnMYXuMqkO
rrwYPXFYjyRE8ttI3Q8Nnqsr1zvA9+Yo/ZrsoexFUc0CU0SLP8O2WvS9GkYmJ9nF
BqkiMo05OYKkRyEyc9l7h3ZHuhgf0lwsS7k9GAFWBKfaHIkg9ZD5Z3ml0f/ZmRE+
+9Rc26NSh6wjdHuoxA9IDLgUHHgIVKKTAixVFHzDkpn1ELPd4cOx/3tpqZ87w71f
bDM9VEJl1e0y19e1c4eaB0mbq/iWNS3RS7tg19vjqLf61Hd93agFAHvxk2dFAgoQ
jGwlpowTHiLS1nmF5fddGo1jD95SHsv9Irg3ztbb9jjUi9mKv753A0G/moCLQXrr
AsvDoKpjQVkGDnVxFhfd/h/4hU4V9QzmraPjWG3YGr6EyjYgu8xNVheky/WxzGW1
jI3RR7qFezg1K6fuZ+5zOmBXnETEmBr0kQsPa2iplSqvaARe4D/5DCJNJrbhHQu6
h3wdJ1HUd2zf8YiXVs5JvTHKx572D4vykXBaYJLoklxkrfs1hTEnxG/tbAvhK4WU
/VJMtdX+StJ3V9YKHBPhmB7/q3QFT8/JZcUev7sPoUrHcNzW064zCClXpjBswjNK
ugUj2DxdDZgda7fRoYRHV0Fs9AbdQeLzZgLWQDjDi/OVsV40Av7Ao/UAb4zEaUkS
k1yP7r8X/OjxY/caMZLLlhTFi6whgDLxn7wd6Maj+8rHAaZEh1TRxS2I47Osz8hs
JMrigLIu3rXwPRdSB4nJgAjYqYMX4VKqYJrURjes+mhIO5f9+myOSpZ055euaeM7
dmbJWaz1cR6JSJLSnWra5ffMqOWERmtmIB5hGq5W+15GxvEDurLadet8ColkBnGr
5dFYCfKGnmDhkJkeCdkWJw1/GuY8GJGcOhZDtHP84B10yvt0raGE1PZNbUyQkV5E
Jq0e5IztM2IUURCHU78KoqbkluZH+PUxqaUcdmu78duYJR97dLMb6iqo/UKRdiLx
tT+Wf8FH1TMNLe+Bu74ibpOR/7ogMN/LrlL3XK+Fjup18W05PBoOAeb0rTlYiILa
bqBYobEwkV7vk7PBrSVMhy7U9YfDjW160WNC7k/iI6sWO5u7zXnSC1pQyblg5mMg
dzIFq2lyafOstuNB1fupJ+em+dqUllCwj5e6K33zdVJNjlCeA66TJ96KHo8MNjxd
Myj/w2Eb+hIc1fPC3472Se/phincHdAI7nme+/upyy5VpRloz+H/Efycm7+ZlSAT
nJwHjEHuNHe4+W/lZWnZ03QeVw81bJMzEw3bBlG472zgK4nsRjHpfWG5CpJgGXnu
sQosWZzovs14wLuKHygfNxiarJH5ROW3G8CfEjYH9D1mHJHrLHublk8SoS2aLK92
KUBUzqdHMqfdzpiFIJfCXE2kIGAFgnEkNwq0cGH3ViZ9ThNFWZ9njCyCuF5zn4f6
8uGSt4cHFLwdig2zZj4Bpnb58bGaxLgejc3UfBp+/ZcZzR0EzBSkZE83sEIQxTKG
cWD9vmOX7wP3W2YePZB4pHFhZA5a2E4B6z/BZR9IyuOprdllX0odALR8/PNNAMMx
eKvLuHEnQct0Ny+pugK7renKDVMzxs3cR+ewd1sR4DxRoSfiwG0UCf9hF7J9/v+E
L3qx1Dwfy8REq6joFoQZHYFBbXNVEtTPSpzrPa1XzmGse10ZT1p3OVWvE1OLvQyj
AAJJR5yJtdK+0qrvjAucy/ywy+KVxqqqJ6EzBnIOK6rSfuEMYEzLVqnSi9FTboKb
La6ljMn5fgY6YaF9bSxVHNFQZRW40F/mnUVnlIktYIlcH8LYiPqQdpH6JdWZnXPN
no6TlF5LxyAkj2JnmXRHfmzgVHAAxVQ87Yhf8xupmhiEtJlLgjuQDE42ifYfzDP/
03h01RkjHC4beJHEQV4z+X+Sutk54cCb9ptV47eJCWYe3/Y1dp8+ERh2yteG/4Eh
OhfGFpyL5i8oQF2COjw+oUeM0aNCv9gpMnP/u5T0QrL618GP5bjMxJEvL+mV4LqW
2vdKhevxSxkmpoXKpXO0HDPXRLaaEg3MzXmpXrk06Ml+6xZo7yjbhb9xGS32Bfj5
puH5SRwnRsuPCSP9j/W8xWP7e6S4oxJiHr0Mzp4nhMIG3HDhhkIK7Zn/xi2OIwvO
+VxZkJimtVOCdCgX8Y7gTIWQuovpbt4E+wuvcCHL0grUnUYlSHHqDhqohDQZ9s3W
Eo/O5Q7mtikiikruqzfg9P/l8JAi3fcibn4JkLYfcdyKE3Ss2EMGrdzBbmCdnRfY
TUznihzAE1XIPSUILgfMKa7d8c5qXHQjery06UXOqN6m2OEYpBTOnTFPGi7G33Rs
e9WUII7mDVbembMxAOBQBOh+jRxmkJ7raaResMaNm1JKr9RqdjmNJ5TrejEhggz3
KJS3VSHCTM5gYX+VXdbOxqKacDjKc/mC3H13rT5dejFlDEOzEP42LWZStdmnjFK6
am4DhBqToVJG8dLsE0/d299eVmzh/LAp+bMBWufLadoy8Bn5PBQvnXEo+q5xF9nc
dMdOFMzma8jCEY8HoEsvqbb+nNvkB78HCcETJhaSDkv0XVOO2MsEGJXr6Gqiq755
/Z+8djpb3usPNA6MhWi6RcwAl9bMtxJFHztI+jVKxLES6/Vd5Y6650oMIAl5WBqu
6M4HFSgERfQp2IrgeZYW0/txnLruz9ZRQqtStycUojZug0R7KF3wFTSSfVakyKPl
2MwQNk6Bwdj0vJpczCYljaDZOnINp2Iq1z5g1+XXRH/1Ueq10CDwDXTy69yvVGua
6AVLzoIwqPVqkUe1o5yy+E8ozE1VZ6bFZgL78VQOVIKGY78ekaOV7JJPdv7O2sEx
T3rJnmTgwE8gTac9QqzQOxQbLQPHF5mIPIP7ds/hpNKYYi901Y5fc8iMkPZCYQTs
HVjWUVDiR6QcIofvxVnWQNVfDXv0nTSVvEPfLktwf/jGZ2da9iwWpG0kw6dexno+
FCilh9IcxmseIIN+etFOgrGHKY+7GRr1TwDGo18XZeRMQspWvmjV+ctWR2t816HE
Zx6Xotmlw0IpLfUjI9u1F21DXMZ7KCgNRsy+qrrJ6iCNtux2nJmAGvlko5jr1uZS
+LGVZtQrFgLpk1RcHbYDOFcTgbJnry1c/gDnNzCvfUO9Lb0Lpk9YMplGYCCzpNPR
WtNYLOqTN8AvI2ZttnVlsQ3/UVEnL1GdnJNrRLZtM27s4cnCdX6dVX/gR56Ia6Px
SX0Wy/vMvq2pFrJ/PcN14Ua5za/iIAoB0XZaTIKwTb+QvXamo7bncCQiaviIxmx/
3ZOF0bljzO6xThFYrMe5s2Yiv5NEi7KZ8L6uaRNO6DAHIVukcZnjd2pT+TnE9UbH
RsRWbn8t9uRjUA8bbUaCveavTbTe61ZC8o9MgDXtrF5Hd3ZV2x4P1kcVXVsXtMYw
TJjhHvxuv6HO4hRYqcIRYLb0/8q8gngsqG8TP3s57RtTTwofecvImcrPJStrVXpD
wVz7/Jvp3b5Jxle2vBYE6snDH7FGLPo5n0tLaPZD54APB6G+FrVPbflCjj7RFFsM
8cR3d5lI0b1kP7Eaawz6pvilbL//q+ZS1AYIbtVErqVBVeGxGVX1ZjHoogvRuVeq
CwMQT9ZL/3oaVf6lxo8ltTqJGGpCRs3WWUyAGzxuNYPHUQcMoyeW5U54XcRUpmAM
q0yNNHjtrSf4f8kWtltVPB2LTgTOvlY7fVviCLDl7TuUwIzpzfB+c4c4W1BAK/6P
PLHLTki+Ty6FXdMpM27/tYacGwKUsRfAhs+v18XbQ1yBoNlHzTgL6I9atavtjeB1
/7vvB4P4w7GbwIB7JKihi/fq7xqVQFUU42qnA0b4nBZ0b2dhC2mrSeI8o6CE8Rl5
C1dTcus3Lxh7pr5pIgfL254viA2Q0jcJcmwQEvYDDrOEPWejubYcnuiSjouqEk4z
AgVSZ3Npv2RJ2DKYLsZh8ZgBxyBWP82UCXBIBR2w7Wm3SqSz8v6Dfr0NG9WQxofR
84rPKsuR92MuGuxwqVsfd2W10vRGEdAciClbwKkXV2k9YCmTXHHOpkBkRLuw5xYX
S5B+1wQlXS97QaCabchM6fpY7G0J8MhYYRWqOQCBLQYLXY61kRodX4cD5RB9/Xht
1xg9RmDcPwQg/SmzGg8p2UgUXqsvGpGteZrRqCew9JXYiv/fMH1a4Ye0BWCF4t8E
7feiH4lI5TVlShXEfL5lD3W9Px907Po5iM+MrszZlxpS6gi5omucNvfylTfXwuBl
n00Z3wWMxvBr2mm1fTMyIVFhyWCslXBFkGDoOsWmxNizmyeAOHI+tdnYfgTu592Z
Lz5q9etX+0sP8KqJrnBLwKVs3Z08tsQApZdWG1BzlC4Dm8r3C4kj/DEgR7HaL2A/
ntGZfYkNKi/4BG/FYYgIb0+4Nx7rc0xlpLIZWrsMfIilqJ6Ib+sKMqDQgGIBd3Xj
6kT7S3dWjjHbKB0x5dpEp1RNAcLFNf8DV4gYDh1GihihO2OOc/qjCxN/qyb7/x+C
nuOzjbTflghb9eybhOIRDwdOD/k4rDQL/syI5Ab0ahXfDvJDWoh/M6D2lp9Qybhn
qWZmxY1K8msK1+3gtu5Y92SvOTK9YRvZTWNFjmr1Vc4jC6PqOLovysNOuxwrdBhW
1r8h5YNH3YBdqDeket6zE3JA0RZaFARJJbc1Nqmja85t8PO8VGBxUVuSbaboSr4D
09Q7q+2uyawZMg5LLVf6OeBjT/JxGhe/foQqG9g2K/aBFXq+SyQFmUodIXRz+3ry
VYb4lsnSU9uCkNn4KULjezuvFl4a8RjZjTewrUid4Gx6wxvDLV9NoJPMCXM7yLG2
KzmhBeiLjIkzNtgxvcfZaJVOYZO1dmtqVHlSB2tzQUXF++5v9NnK/ctK4pPN/Wir
rNlcQr6baFOprqn00H9NsuisuVCp1p6syvudkXTTS2j18dCBs93Wgy/DutYo77aE
7SeGO21yyM0W+JTpfgNTZfeMizLPu018gwZPQJfvoNPprpo8SJ/ovIS0hCuu8SuM
+FJiaJbmDv3A6ZCk0QxUJ5ofCjEfW9fHO6FXT03ykpA5FrR0o+WI5YwvSC1MPetY
3LrWEwdmdXrKZvKnXq0AnY5fwI5UeamfZxIiMZNtQNio6tfEzOQ9qLcFDMGZFW7Y
NKjSvEy8wNYVbZPnrIIsYgxK0mPwHuaG/YzxiKGJXYkeLhSemXUB9EaE0SMIq47q
Im7ahreMPy2p4ayl1vmSz9ZxHec2eRVV4fNh4BdDxyp0FkD+hem22bgk/+DOHT5j
vlUX0JkWYT8+MlKO7CDKStWRn+YWuMK1YosxmcFDlSNCDdRoWLT5viFFAx7Fadys
go4OpANFhzctjS85iYA0vPP8cuu8zKPF7wENNx/L170nhWFVJ2Kv7PcupwovSp/g
zRPgEM4gk3ISN6gWFJVEjkrFbBrX45K4kjUJfeLclxfU34afj1+BJt2uR39r4U+1
zkM2W5NMShktjJXzyVvS8WFyLXYE8cgJTfIUyYZmf+jBLpdVvv8sMPnHjYkJBeL4
Cm7yYs4zdaI5j1CKyEUXsNuKIzoSiItwxL3KJYwfR+luhfIaVrJFkENuIsEQqAHX
hszO5qL1InQr8q+eouVVx7gRQ7kSGC6AhWtw8w1KeAjm0LIybs3DBCxOuhxQhMeF
/ZcdkhFs1yUgSo8i54W5VMeVrwMBVutfBjk9cWCLbzM7Nv07cNtUyKcT+QxG4fdr
Uh8gFA6WtMdE2Rt7kFfd1GvU+EQSvX6LiwdytjbFDX+DHblAHcZTqdZ6TAcBJ7xW
fyjTN+C+/0ric5/pe3AG90P6Lhe63pTdokNBy8LGMUPh5sqHDYygazYY5X8uNEXj
kSibeBVB4X2CB1RKjxk/JxHQ2btKxr+V6h1S4ougPpuvtN41pnLfQMQmHvY8Rs2x
lDn/FhiDmauTg0iniNPrsSut5upd2tbTZaH4GFCsNuXfjTntrWNZk2rtUf0xsn+C
yAxLvB7E3/uacH8dd+JFVP6zanYTXpdkXZ1fyfUEF3ZWSljTujRkqGrxZXDSKbck
+yvrvZP3cZt6MqAR+8dYIBmPd7a4SbzzrQTKeBgWO6L2sZ9sY13Tbnv30TV3iZnr
iRAQ+vej8BdRTI0AuzJgQbgbAn0m6lxWFmHcyU7RrMhm+LROsFSU3cXH2s7n3BWE
a9hy8PuBEj3gWj3NSaM2VioDXXNVoG0WYwEn7mbc81o9ng6YxdD3UqNuWAb5Il6P
+VjLkj/8TQkYo1wq3Qm7FvYP+owt37sJDqFyzUoYb5QMiWKfXRn/w1+eY+L4TWkX
cBGOxCttfeqCm0ruOr3KEV2MHLOSh5dpBgrXR7varjwK00YrMcrghUtIT2FiAYYg
1l6o0c+CGo11AIQ4tRJguOgmXJo35PGQx6cpJnVzSssdFCJbMH+GqqVbdXS6Vfv8
B5ZqDCdU6fQo/fCEA12j3QmFJJIJgolO8RGZxjRy8YgOWPtA3lb3umH0Kgde2BKF
4tlDR2XEniUGgmd6hGRzAXaqGISNv6K2cXfVDxkQpAInhj528vEdBkdyrDog5c/9
z2yw6uBBsnVmRO8WdBOU27iJzT95PvpQfJ+TanmpJogFWF53xmNQoYmaUG6Uv9+J
FehdbAKY/YWSnaG7ghQ+gTXNoOn076gTovtsAqXzXWKPI0Eg9uiBlXBnihCrg19z
AEmDFI3WZVyhWcIUXrWFlYO11jmZZEq+ECjXki3Grgd1Sst4/6vQVaHX58A63+ec
PMTNQomfuQoCFlm4KKnCGHHs2FHt+168YfwZEoFntonCHGoJ17+D3yazJRQy/Vn/
u1K+rdJncsEYqMaKePtEaUcEBp9rUfXebXAfCF2jB6uGLyTV/1nYYJJrI04FTZnc
wm8yKZoBe/jrmk/wv/S5uXo4hxZb9Lwl7ckgwLshsW6EL1FGP4Y+wIhBYA1vEi6+
nRZ6i3QxXfQv0t9j5ApIfAnQqw375gjUQVbMnG9xXWrjp/pLuishqh2kaODt+ftJ
CCigNsT2n9Q2D3uWI5w2cnBk2kD1Eb5we3vzM2NgNONYRFePk0H6yd2Ff4mzwcfD
mI33B6XVfmszl6LFnp2N92ialR1vdYxW7REm+nTiwovQ60npnki5t5Aw9nHmwodk
X2sOq58TSflcY5hoeBfyHKiFb76P7gXpcqTGphRn6kXlBEYKDkk+03xc8F+HfSCt
KMke7saBKklv4rhKcVLMvkfDZ/LdyWtREDj6K21dwnOazBenPYkb1ioOcjrjSJPz
QXbGwTNJy5KNEj+J0R6I1E07+TmX2mu9LBetqV0Sr1ydF8t/f8nJVLNwh/4r8ocS
cTEzHzOm4oXPw16jd0oWz44UV/wxqMwMDfTQJfKUDXJovoDBbfAt1lIpc5eWQeLZ
kBX2NCdRP3wa4P2ForPyXYz+kPXxduPKqCMAg5hBL8Y7mBY8Q4QEgoXMcSY9hj5Z
yimteLluH0puZMpbcYfsthsaUEpTQjnVf7TSRYjDmq4IslO3Tk6QZ1med7CRvWCw
GAVBDwT2JX2S6j9p0qSlQWOQDQ5QhFyb1YFeJRgcRTT1IyPgdE2N3QmbKTpBpNP5
e3dj8PAHXP8NapYKwNcvfCXJjjhYFUupl6ewwupxsgKPSanI+zIok3Z6M2qr68Z6
a4Y+KlLVtVj7mQhSNpLH4AO9QNj5xPyZ2HVw7ngDFQxz6CmnXdNLmZsvxj5j2twE
EdJR6XlSU2UsGa2XMI6siIfJ263raZvutmmIQ3K57znWB+bG15fvrBME4cJoFPGb
kj8sV92T7eG7e/AgFMSjnGbrKdoHWb77B1fg2MWe1KwBR1/WDM3Fg4ByJmOI0NXB
gZ2/7DOo6YQskQniePhWNViXWHK9HpqheEsW0FC4dwdFBoBg9aMNLjlhAmqHXC8K
K90aX/q6cApaG1bT9Od/87aoPaPW0rvI5U8boEhwLvZ63Sy92aGtEnjLJN2Fz0fE
HOrJ0/7L0JcS8EMNxIy4R5PRrpscQxRSmgPDbxQ7dbbZCMwpH5lcjwZ3hQVhO3P/
CwY17zTqxqKT4nQEICg6tZdQIbxNN2qD4SgwGkmAUavtJZv2SOQTtb+RBffcghOP
OUq9Gidh4Qftehm0ocYEKV+T7qTArQMLMJjrkoPqn1LklQyB1a5tO338tdQhlypJ
eXQUwJF3IMNn/KYxc0wdYIGqYttvDv4LPuDmG6zKtzF9N9W0KQ62vNl8sKgyRNxz
K5ifgTlOytbYp0FlzpxgGTu5IWhu1UALJdIeb+duanaZspa+EMjs9SFbf7QwfE18
D6vgpxaW6j0BmOaJqxYGwrfgp4624BNhSlU9LtZdKJ8ZTKh80N23MDnbzCP6gy4n
W6genhWDRMWdbbg3d+mRpt2kJ5goHmF4t98C4nHIXOwL9sDYM7XCBvQuvrAWlHNM
YwbA3jJlo89YcPoE+nFTumToDki/170eZ8JC4AhSLZNihWRdWkcp5JIwKVaLfqSN
st9fwVIfX2xaPLSCEDh5UTDAWCG6L0iFBAjkegmGM7ouB5lAVAxLYF7ZuxmDBDMs
iqMLWSU/HVwH0QN7QUOQBKD6ywZlxHmHqL35fBH9NlIlWiho/yYyLDt2Jo/VlH4n
JV2WWN4p/ak7a83VUwYazyjSc5n4MbFNFm2a6aSiXvSnG8QMjVjvGPQv2PBvKTYN
/qzkANXRO2+i44LoF4wStKHK69esXX6QmZpQdERhMoa9r2Np6H3v3rVCd3Gwnfls
cqPj59xxtVkEHL/hiv6xjhI7MLAuE7is26D6gmNrIrsKCZ6j1CEOUsdCeD5ByTaN
dqJf62DQ7BfiUbz3Jui9xY7GDY5VIFFxIg6SeeTdlfZqLSFAvW1ASy6W5pTJspT4
IpgQAn5ZbS8Uwfdzy5140GN9cmY9dFBIo5kjsSrLU2AdfQEpxayG15ZAtY/O/HNq
dDnE5+PW80mDi9IZo/ssGzMTT6bzHkMTtDzcvCvz56vMLzljeOPQrcRaNCdMd/lL
4agvdbr61YaegGUkuZrR34XsZz0TnbCrMDZB4CQmyk9/voM6YOG6Hi1wXz5sa2xK
20s7LeXm7M23zQXS0/NF9EG+/41J4QtfAK8wCGzt3wsAPS/DwvN/Z0ce93+RHKYA
NggXxUWcfRrq05FfDTJr34y3f4Eanq+Myp5zG3VL1n+0p9YR+bplh3UMJeNNtd8v
j9cC/uASzxTkVdxWY6EpRcBCyO10qMeoom8MdGAIbr6UBnAiQRNp4w+az66cTRLR
wlkR/DUxU7MYtILOYgxFFCk6OFY0ciMex0fCvkhIvkwLjzj7XmXp/qWCl/DN9Wob
gZMJ0ZXKv89szmAOmFsWGQ09X7YmHQ/QE28hi6vs1APmUzg/e5T/OGI2c545Wl2h
Oht5mHeiXG1E0dGyKfLeNXDM3kO1MA7ZKQksTiKT6KtIjmfLd/fs9QWerxuCRkdI
Ws6bSaus2J7xJoHw3+KPoSLhb/GZnFHZ4hVTdUTIZeglhLFXtDSUQelGCvENiUDI
747vOuw0+iAzNCP0s8dBy/WVvVGUeJao1znMndWfnmy6Z2Opw7CaDV6SWXI863cZ
CbgvITs1DSyqbmyN7GPT3SFgler+XhYqodA0q9WmoQ2xRm/ZNDBfwgFhEwVRcssV
/rSYn0X3N69kM26BgfB75dNO1rf3XOQAvGZCu+RcIwzb5zK8E6US8juAElAYuSKm
8kOSMiTCi2HNMoNxRNFjVzE25/a5SDZKzmz8jwl2V19WVuv+mkWNxP6W7TB1p9+c
QszqCI4OZiqUvGTLpm1uvJnluU9XEzpuj+ATuPmYQwfVJcA/M6SPkgfv6G7beyJg
bHt2Wwmqxu0mSRhis/+KvdOfqdayX1Zhses/DHGgmN3jN1JbfNcLaGTOUIakCZmT
YHGVs0VSrOzhyO1s/jZkFqRnJZ0sRQH/ipbFiuttDfkHwYnCaOnGvJBEWSO2ltR+
k05U/QB5S3HY0VQJUr0HpeHLhnQ0pQWWNTOHiJ76ch8pMozHenL9ivJQSlKiNMFB
jcKaxYfJXv1SvazFwcNO6aP2cKmTSN248Gu8e6jMiuSCRSKGTLI/x39AXZmsF4NQ
hRb8/N1x+VhPWUkOtAhIUteJyv/bBQIVtKtSbCpeosDsPNgGS0IU6aI5U2YLvsZK
SaDYaXOD2O/2rhOtUa7KEAS7K1Qa0kVElEmRq83cJOeTo++AIknE7PHQyCfHg76/
8s9XIqx+yhOiAddItd30vthqg40juY1p8PDG7IdciBnJq+y3VaSPABIN1BUodfMK
JotXFXjNVfHum1bxmOhNeSWVt5+Ug0fyHMML6hwIF2zSu+qp3ptZ8wc1VCPVsVxe
yAySssVP2MO8PX1Vj4N+q5/W62Ef6F814hGnoNbgHt0ungZM6ihfuT9InoGT1ee6
POn5fKJ6XPgpyBgODcco9a8vIHGT1bkENJJtmBN1LRUAXYfh93lkBg2eTRKMSafv
Ccs9c4PDZX+WoM/I1/e6Pj/6/12J8fYJ+AUgeVgs657aWN8wC12TNuvhhbYzSZ2f
hJkj+htGh8aCkpag8V1w6wd8qFXVTc5A8Ldj5nnO0V0QtcgBB0JRWEEakqMI53+R
DeWdYLTn4EYSH3iHP4cYFBDlrZ5oUkoyLs5NPAq9bLu17tRJrUFrJZvUxLGgm9Ls
Yt9CNDzvt6JvrVxfXHk2FlR2gRSNAM8p0DPWNlI/uReuvvO/kdV63kwoJ1KumrVF
77lEuHyHTlpEi4MIEiDmRlOAlWFjs/f5bE5tUSoIuy7ThqipYxu+pqmLNRC4e0fF
N91srutdIgNl0ev/5zPtyB9qCser1o+1vJJdA6vnWXWluGohJw7ffGJCblNaoUDS
J6XwAyhHq9bClNlOVESKNF3Fn/Z4MCBE2uGnfI4RQctJIUS0FvjhQ/4tsBQWC36u
oxUJgr9zDJrppfXwxf1spxhbiY6muJBvx1St5TxysXeLMzmX0rBgJhnWxK/lIAbh
HPo7eoGq1LROhPaL3PNmLwQnz80iwgNPp0cf2Z7yWTsntPKAR7ANjKEB4bkCNS6o
QdMBfxMZtZVRW+pBaGsP7OOMn1EpY4lcT5MtX9C3hea8zeMg+Oa4g9UC/O8UOoek
gRtnRBX9VtblJnYofJfQSYMmuWtdNuoHkoj9siKcZuxsnjyJSSCmFYPhkZLg8Mv9
wklfFDog2quuKJTRszerPwtZm9Z3lO4qtNXGWiWS8d1wBd2Xc/KaSwvyvleef9FA
kSy9IUlo+iWarO4kQP0Mo0LJbwu6BJaYLFuppB2FP2Qq2+t5fPBc6eV5EKkzHaKs
IQJvVk8p4dgGDAXDqjqZrbhW0ovhyPpE9VRBmxMsYVpNlBFCBM6v+PiXbW//t/0O
/gcLccePVC9tjVNZ0RIZJLS3iuCG3BUnv0rHcMApKeu0M9ujKqJRdM5MZ5BOZp9g
o7LPG6sJ5m/jKvtfeV3kuyilu9fRhv7hnKwJJdbLtHMweq9ispI/eWST6kJS9YFN
TftvvA7w6Jsda1xx823IAA0fEj/xgQqFh5b/LcgL2TcDUdhN3hFH3xCcGe6xzyQD
M6QYe7eVdq4OaESCWRQuAycsKqycc0/wxPxOr1FS27tYE7ce9m8bH2GL3asO4Ue4
YPqniv8hyt7ggrC28dQsxKWkyDzeNyA/wIAHjV+5mqL9Zvov2F9ynUxyfgMhaOQ4
b71/xy3+fc5X7580OK/P9KEZdiSMq1PLxvS0yMQ/xZcseVrEtMXgR0UKZrodLzkp
MKkA9t1Gn0BWmy/moLL91zQIXV6WRY0HGFyjs5seUwHXy6R0Q4SLOK5l9O9Nm6vx
W2TvlZ3w0qv+xr0roLke0o0mPhP+FKieeEJovKdSRa//tpsj8a4tFp63SpT++O8k
hQGl9JzrzJVRk1+/zcZHx9QRKnRD8B6+arYW+66Raz4BXMPaqrtCB6FuplipxXGF
lBCcLJe/L5WkH2rrAto7Pqh35hyfYp7CN1MxRyIU8kVKNutGxfK1CzetXD8VHCcq
2hbJwPkHmjgdr5g5xZ9KtokCTKbh9E+o+DgiqnvVnC7DJgS43/9H6TaN4UfOw65H
eMC1oN8zAAMxkRxOd9qc/tYzeF66mcnWBTaXFnNVk2ynbSt1D1bh5QpaIQBEHC6m
N2dlYRbrOD14sJazh8CW3bQ2HebW0pc7xcFa7k46QnEhwgIzcIVbE07gHfjtzK1I
zUbuHJzwdjr7VEhVB9fyZCLpxzYvqCFCrjJHrZC7fBp2ddPJkSWY/5sw9GLUcOFv
ExewyV/czGuQwPKj0m0i259d/oi6I5MfFOpQt1gngPPwoGty5d47y+9JE8bIWRGg
JjsLvYVuA5Zo5Oytr6zYbP0L0P0lnin5VnHnStAuvHi9L3eAOIYY5kx4LD7tMkT8
Y66DYwCulUQvAgcD2Gh0oPa+GXTpbm+Y9FX6UXtFAvcIxV0+IooqKE1kWvBtz7/G
1FaPsgeekEuURptXjvgHYoDP+ZbM85Pl9CeqEvehRVGlDHCoiOO3hxvPmkU/oiXE
WBt5/RFGJyDBIMhIYj9MMzKSr5HfmU6YSyx7lnq9UFPPx2PE9o52yBbF+KK1z+yX
X+XUZAM9bDHdy/NE5fHmwDQeviZb84ZYEDIg2/a229yA+WxXQNz6oDZ0iK3hDtxl
PvMcs0AlrNtFTAqTmh0xXSR0eCkJmTsV4/8bupp2ZqK05nROTd5GFQug6tPI7u0m
XqlRuexGExs8XzSdck+havA9HX5jyZHcAugGzqfaDLNBkIPFq/iZnlcplZQtxYtu
RfZb87Zn59OJigxpIVNobrOntEKXP8wOVeWZnCa1ILSn+U5tbSyV/YQaP0+zLPyV
qpAyHAOzmL+nN4FEtgiJOadJK4JKTH+qBj5FEwwg0xHyBF2QPYXydOvcw2yv2tha
5ZDCUXkZ9zcEoGJr7oDly1Dp5cGoDBo1SvayCrq4Pfbao6Bxr/psaQCEZqES8bqq
AK5dMB4XkYnLqqnUpzcMMtt3HogL7VsbC+eIQRpHHg0fLAwJTGuf2CVcQbplYqiy
5Tdn56oqJElfhgF4rAwzW7gY4Q4C5MzTFF78aIBV2n6ek/SO4OpmsucoJJHDItxM
pGY3FbXJ7jIGvsbHqHpzdbQ3ZxvIPgdlte234qfsoUyPEBjPYlodZVvnGgHEczdk
mtpMRaLHisbITPs+ysGYNWyMfZDMPzLJWLjZy4qOpCQ6zhpsLGi+YnylN11OCByn
VBU4HmiMQ89a7Zv+c9EJ6COVzL2CLiP2bsB/hz/+020iFijmYKawuEYQa7u7BVFh
9lz+v8pGAaaZbnlQm3NrqEQ9VD49rG7A+IqtD7zamBIVyMrTdf2pp6h8uK9TZ9BN
TeOWnsQIkEOTJqELdvV5kLhYxSX3KXkyGJ9PZ2kL+tUFJkHXd+JO5iMUF4JapZhX
x81FcJ2PqGtiDX2xbqpahhOOGrF9WTmFnlA99BSUHlz3c9YDaCnKJF/gAp2WxpEx
ifM84Fs9yez09Rr4x2W/QFaV+yf0OiYxw6T5Kg2uf39DauMk1ZvjR/MFjk71B6I6
sK4iuxf7IspH+KtNE4CNmH0dOVc0mdcz7V2O03eBxs+q/o9ctZXpc2cUmMnLswBa
tHacbMnI83lJI/faK6AW2/RtC1he9c4tWyZm+/+GtMbNMAlQ0vxXRfp1jyd/Q8F9
yz0P5w2Ik5FO/lL79r0fDomujtX/BBoa3m2WfzbJMy0v6Agj4efZoCdQhNLPsQ4f
NaEGyn16+luPadnJMxAAfmBqfxHqMrF4iY4BfIrqVPbMDWnJGW3/gJZWwGd34cWx
z3TSMN9TzgT+bunyon7dNzGjrJlqQ4aWPhvjbfrHLLqAShRsFU+LaPx96KgsEpP2
Df5W4ewk+TGcYa5UWLhupMGTp2Y1YgyHGwfoCrcwMQ8fycuzPfZk5c6PUDa0o0p7
3wKdTeV+OK7x7wFkBu32pxcqcWC8f437QTaBr4jXmhjQZ+cuRNrGSLAGWds+utPS
BOGkTyTh+x6sJ/vsJz6x4RuubqYkskBIbyCst7dLX7KeA/BT6weowwFmhXEt8Kwa
2qhf5TBiuTCR+2WAmNtpFWlLtJQgOOBP122/GugP2oKCTno7lxs+yalxnxceFD1D
SH/jbGRPJw7JSya/wgP0WykkthfoST460cwSZAueqAB2HCfzmOYgOfna+BrVuaYr
aicibR83gjDc9Pxxv5El7mT5byoZADeHfTQxKLIXv80foFsWaVxYVxj+GSzIpK2P
hQg9NuC360qvIReosa7zR1NuH7Y438EfbMFNCuI1ikPo8uL23YN262zs6waUua7p
3+pJvMLFr/FsTiEeG9ZWfPn1DqkdvxH/3dDxkUVnniyI+TJOLKdTH8Mb8qDvMyif
eKHPbeb0wIu3fr4Cac8pJq6g/K7QaFfow3zxhOptU8dpdeU4d6KszIlLT8Vxe8H3
IR4VrcV3ByHtz0K6zGhLK1OeLBNArPvsiDady/uF5+apieO1P7A8PD0VDLNSD5II
sIPBw/tw7pFh+haJ/iwNZlo6xf9lea7DW43XSxKe/+pSH3uKrWoIrZVUEL2EKwwv
Zv1tXtngxWwPfiq7ZdjR4I9jF3KBuMVWjGYugCotuOjBhLJdLYV+1ExBwT6JrEOe
lzOFBUT7t+aCtFHA8z4H5T9EgPq3i614owMiRTgdke9XYZ7qKVAFd5LZflEuUdYz
veAXN7qE0OtyyJqeE1UIuvsH3VPzSaHc/eYUWkJ9xIDyjoaZTSzGYzJknBc42G9Z
DK4Kfa957rSRSq3rmkA+2WhrPVHQzUJlZ6LCIGBwfVAvNwKdtsgwhCFUoYEQYOey
3ztBJbdqG9jM7iGwnBBy2PHXzwQD1lRYdgOPbZ4nqK5l0wQnQz8uON9TuQhVCu1R
MGMGgBIywpRSMmP3yRZJ7jJVCWK3b7TW2ele7gbFeEqoB1KY/joQnszwDUx8UCNp
BlrjZQLWq0pceQkPp3pa+myZaoXw8/gRP5ab7pSFivcj0ZrKs0vC8IND5jIfqys7
I9nbbatV1v1amGmDHTtQxZAy+8S8/s7JWP3YCthH8sDNtpVe71ywU9MiGEv8FbsN
AuPCr621w4rSmvXqlhmuExOp50kzFbqBeatHUKAiX5B2dVsfmePzLUDCJgO8h+yA
N+7s7mu/lxkKspNjss2E8iYMSvCZB6+aAm3XD9Weatfhu1R+AMvKT1CAU9v1A1t4
KItj3iECu6vuQ75cKAxUBGh1YfD6EE5XU92sQwJuJ1F5FXI8EZW+KZhl7UMPXwjT
DKYhSjp46RaUM1SlYIwknTbtY+QM0epI9shSVyfUxPF+MY57y2tHVJ2gqJBrhQHE
8M0yrhiNBWBHghN8WBkS3R4Hy+/kR8K6dkQoui9UWU0d6Ys4kK3LSL3ZhWPFY3r2
vbGEZHKywTtBG1imZmnX64Zp3SMwz5eSVjySDb6Pv8/qSkBNqzBuvRuIOMfv2Bp/
yQZpUHMuBSgFUMJ6mv/XsD6pAH+4DN792eD9rjqfVp9o63upKSpNaAFZDtvO6oNJ
s4o3ivZzbz2fGqZTQ+xetS9+SxKhJFlhPcsd+Ei7ysjJwczwMZxqV/AGCrJOqAw8
orm3kPzeR1ZXr2MEagJMlAnqlsC72+QPBIdxJfEm4fhrPVPSPG7e3uKOyR7G9nT7
ylv5s8eKIR6+fAVNuV6jfM+QmhA5W99Wa74P9Q5v/ypK9ev/v61p3wAEc8IjaXNV
wEQ08oRdTvis1XN+fZCXSITxThEmKxqCZ59/DO6OTV09lyKsShznI7drtkt0htIN
5o+6urOjQRhda+ehssxQrJ3QnKJ1yOCYy2vJOj+zce7b3l6et85WaD0jkpKfZVip
0UWj0kFbG0f7emOX5HtVJE/R+Ir+/QMOyx8V3lj8Fb/EL0zQo1XB7Yzg8tLb+UXH
EyEDHyOPFpTRFsEecLQO0ljO8P3pICLC20FrQHfwx5l1H5T2aNMrUIqMB2Sl4yU7
DVqTTZFjyb2w5mQPIjSbD40TNgW0cs0pu1Nn5P6J/mEABYgOxP3AORbvPTMpEKYy
RzogCR3XsaeX8ca69+ICoPvydem2dhwB3NgxtWmUuXbiUV6SBmRQ7H+rjk33DZXf
DN6ERBiq5rAZykr9BorfjUM0oe0LubfH5DAjYMSX1931yToO3aMXBSlOGSe+vVIP
817cfA/ka4t2h7uuqaZv07yXoDmBUnAm8if/lNizE9KjPaj0ijfj+ie7O2b41Hfx
PfOKtO2uTkpLatZqkRpaI7uNfb+yy2/VGnbXOcCfkBq4IjYSlfh5f0ZAYB76CjuZ
YznTjnksBIZUslt3GJurEB8p67Hwp3ak5nsk8KpN3tQknupV1uWCDCXx9N06SNvt
zaaBfkGZdIxDyzRuSPKYf7IghEhy9SskSFZU9XmNSm/MB66QpccinPSpTtodCAGa
k4nIZma8plRuDeXrW0OozrkHzP7Ipc2f9WGiAW3gDTgnMZOh576i8xiCEIz6GyJm
7LRac7ku3UrgPt9RVpigl6hmE8Nb/HREMCHBLNJoQn15JhRGcgcTTiB62TaKGU26
PbIaSk8m+K2N6Coy/UO4fRkeVeUb6O8Xa6b2p52sTv4eAPFn67X+bPhN0q1mx4cN
QzqmkvGgFqRjFdOOO5UAhzV8m5Ma3ZYIxmTuHX6YBlSelF3nJsqWYyzq97Ad3R0d
kBwriySy1N1qmOoWkybnGIE0aUC4L7whx68G5n8L1EUor2NLRh3V9E3h0+wnC6fZ
ss0oOpAFd18P3X8UMEhRmru8ffcvqU/2BgRz5KAis9VhfcyWxKi+7cKBLDL87gwX
w0jlDCWCfgKGBB35lm+xIH+EhgsTZZe1JveQlbNxD8w/G0AaWYQw6JbljzIISBMw
b7OrK4ZU/62GP4BKPFYNwjSse63aYVbtjUhkVwIyJ1N3Tg9AoNCK7aN+9eMsMQCl
6Es3Hf2KH2OnCpQ4LPhPaXH0HYmKEs2nE9oM2G3Mq7YQ7ea7cGOC66HFrqDFIxJQ
QkoTFRu8ZHAoM1mHWIU2E/WAWfZFRAtlZHsML8PWfBcqCayTZOdvQrH9k0BtACDe
CURaCyTrATFUQCIFhcbELr83pjbVNPuOBsJb0yzcE24BCf/jMfaSe3YpnIdC8Ecn
2wOZz/g77oPrxnkuCmjepS4Myyn6wCbmrmPmy4bMyCZt0q7Va/GoCguupO6PicXj
RZL7rFGirzf6IEGD0RxHhaZDf1k9XJH6C3CaIplF59gOiQoAIpY54rzS/rdGllp0
psqb8FN42yZy79zJetV3M2BPaoc7KTnUinwb3CFgu2hBtyIPjvPN9KpuAX3AyC+M
w2kHcQgaJ7t/u8UDhmJrhfTeB62SLECCwhqt6iuv/SOE1ToyKSoF5ftVnS0bpApa
ozeepOW35h4ALGoudSyo5G9Reb/ZpnWpcq9zeaE1YJdGr4TmOo42ie1vlYSl1Q7e
SjTQNITe3owmoG6l3aiwcfJcFaZawfIlE4v/whlLywBmDxiXVYIkDLqKQMq7py3f
wknIOFDNVJhKNwghPSMqOa828DWoVRrcI/oh5bxJ+XKu5LlECt1+mnUEi9ZEu6wM
IKR6TWd9VZvzFu7NSqPI+ft5RSof0BE6OHHPyDlqqZUR1VyiqpQvsDos+/jUtAQR
4y0tsucXnEIwN5QqTdcP/4S4jk/Wu/oVjSIVoHxP83mYKnQrWaZp5bl11+HJU9Hf
Vqy8AVGbpfjKiVOyTGvS8r/ROuktPvCXbCvDZef2OoraQ6sQgSFiJMf4GdIOLV+P
BGRhW+zZJSzzFTRQitRjG4uEGfq5akolrLvj2j6zvCy7Raw2c4w/0q1XajYt73OL
6+Gh7UK/c/DMICOgTupUi4w5wpkgA1bZPTjQwVauTtYR8S68flA+IWPqxVGmhnq+
/waoXS3ZwWSZmsTgn7Z0lpTB+lJ6L8bRd8dqD+GwG1SUMsjFy5zW0lpCVlL53GQV
eFxleUvIU96fshGxBEQvlgciAkw4esESNwuuZxNHermeccEf0JFGl0ysAsmvNHFC
Xi8mUYh15hpF8HRfh+gttu4F5EgffB+XkOGWRtG7mwhUjIMCu8M0P9K3TFgwPGxL
x5PRF/DuzfFhAawi3yHTlri08voYNmIpWOeysv/efP3TMvZQtw9g+JzLz3bJbdkC
Hvy3ZOT80WuphA6rHCdfhpPs5fN5V92fbn5KURChqft9QCaAZ2+fIJRajcv61Cah
2RjEtIJA10uJYweoAANt1OispG+A3KXKacQvIwFE5t+UAKpfYE/CgT+i9MrdzUcx
Cn8EUBjIUogwJStF2N/eLHHhxwb6T9Bx14mj6PaAPU50c5eNFB+uZ9PE7mu83m5l
qpqpWeV6CRpAHPitNrDemXiKKlK0icQtl/eM8/Y1Bjr8Tqtpl5fsFH646Wj7xMmT
8xtfg6wKtPXgoJTVsOA/GviNqeukTlxUbHRevaUT0V2WGpF/FdfiUlE7asu+ErsR
BmUcjkA3Nu0lnD39QVA1MKZQe9/INqlj7oRwjBRyvb1WKGU/dSqXheNHZvgrylWQ
12N4T6csMGbbpJ4t58hunBpCmgK/1DHOefvEdLe2e6GwM6PtfeEOZRVuCCaNDShw
ItXSphrlR/nRqVqY3Oy9AcU3LvaSMrfgfZK31E+vRyQ4+QSminyeANEawWulHCwF
jHoURwhhddRdQoY9pzXxodHKqaWI0eM22XZ3xYaaass+kgLdglxBKcwdfFQK525l
BzY9SIl1VTq30Keh03+u9By7HsZu8D/WRFkVSn9Yvbc3byyMHHTJaFVZll4DSkiY
ac9KRSEUMd/ImlFM0EL0zEP6taO6UU1GEhbol+XG9CiPWVZ4+0swcxrpkQKTWzNk
hg7FWOosbnHlDNCH/tMA6aO+qNXXYP82oi2tARXF2/T2kMnf2TzjmD/ccnetj/kY
Ixb15DxwbfYh5dmmYQactN3XpJKBUuDraOU73SPylA9+RTwEDuqiyENFXcfoqgWe
L5UGfHaM/4dk5HWbs57my9MK+gJ+2VkR6Lr6k3KAd6ODbijPjzBPjyhxpENpUgOf
XNjLwJXjfBPjF4RLh4OceNqhhWYOCObgTy2ztWp9ebRJ5g9hZNtawcpicW7RF6Bk
SSCeykYmAU5kLXq3HvXBrl0lAB3MImxbtaT7O9bzkyME+f2tnGCMbyAyHqe0qTRT
/ezsZ8aSHF81ewTSJcPAwdE4iTSPK75Cq0tu0nvpLgmhEmbflyoememT5R0xyhY7
e/03t2vwUeEg8Qd7Qg+8sYSLQwDBvwfDJ0khqUj+ob+JJHEtcozjZCowWTneVptY
cB+yC8R4IK7tN/r8SP359j/rQQ6+nWDMLq17PTs3JZOpw+hrpgEH17gMvLe1pzrL
mkIC/BBXJk7bSWFiIvG8QpbcvSLTMqr2twKwIXwEW9D7xDPRaB7/cqhImJ/dia8s
Dxxy+Dt92u0nrCEac/cnYFstj9M0PLDsqnuaHWdNh8kZfBCN9Fp/dRCXHw9YCLYT
0XNg/Fv+QGzKwg9/4ob92Hfyu3BDxIExBY4h4wov4YO/dVqeQFPvPhBN+urtDEw6
sszOjVSLKBFlbyR1I+aiKgP9rFtjKxcV9icCCCNuS8gNXf2agn4cMdKOa5mKhoaK
spJXmXiJ64w2oBjO1CtL+Qh/S5Jzi6Ud1jz7xHcfRqIJafeGDoMZuMEVU0vq2eI5
Jp7+SjasMYltbX+FK2tsUMzTjCCP1QfnsmJwL0UTxbINlp1lQ/8zFcgJKXYB9844
EMG9fDJ0eltl4XbnQL6SFwf9PLb5TFFFqFTBLlCXRLkDVJx+GB+xElfFx1NwD9BI
mlQUoeEwh0zY4QnBi5yIPmGd3wS4wO37iNUqrwX6Z7Ed7iZSwKyPeAwYn9FIzCEu
lgFM8+ZwZtTTCL5Z6icrRu8LUuEEoYVBV/zXRbz5ZXW1tc0NLb9S+Ij7GjYugpKB
YLQOqpvq3V7A6XHwer1vxTJTDNJf81eF/cghsGA507yX3qqsnvHuGKI1tq/efvB/
hOsUjFioCAO/qwAWLkdUGEcmQyr/HD7ZdD1JeaOXoulxuSXKdbIldwWJ4VlDqkrA
ym9xqoql/n+0aqT4joKu8C0B/4J+IaPZLN4ubqJUTJu5jWqA5K1T9/x4kClZYcl1
4Ut162dwacYLR83f5yLvuT16gDSQN5v44cYJO9vxFz/I5vXSVZYgoSOQrHFfcrSa
ZkAA8raXqys95N9Vb2k1g7ozFi2/W0nnSDmQ6J37T85gCGTl750Zfc2eIX5Ol3Mp
JXEIqqtF2lijAPr8AJ1bjoLkFhzFe+y6bC7Cjc8WXNXYMRVGPi49ougy4YCSIrsb
nETOlJbCU6tE8SO2FnJkvgxBPxZYVOB7hANoEOBBV9L82AGYyXBRm1Z+I9lxndfK
NP2glPaScTkwXRfN71DySNEVlTOiuKbHaa6RhL3bZSAFk5QNSuTReCkzjPMATYzY
/iy/2ITu9YmS6gnIsO/SeA7/YBbeJuFUJUI6v5zTMzjMtNqnpPnhGxOCuYKeOEzT
dddsClrfknZop9tm2n9VgThHbBq9+DrisEvBHBmDGsgFBhv+Zh8yFAHwkAaHaKNb
fzP0f4Cx7/rd1rxUueLbXkKluKvV7liaipvQP+I9HHKU6ioCW3K7l4CHGZT0IFjR
jOsv5BcopuwTbX0dbjOVgxCYi9IjSpk9G5RytoxkDHwXh+kcE+k7LdYauko0XFec
QTJXNqn6Rs/1+HtXSViBQCEeJM0Pfprf7i9gPsgrYqQHLCSNbDK0E4nhIe0DfD68
7GxBD8MNqJ//c+QYRzx4O2+hD/H/4/dESGf5+V7zTWEGRPdSRS7Qxm5kL6EPAigz
Xc/ApWxTrLETC/9KTTTK3TmCdWCyhrEbyYb4cEa8ckMcnl/acMKeGkw5paJWdAxM
6WoDaIrPyXJqlhzSxr6Nv5sOiYzNbYVBn0t29y/AdzaYNtr/W5mU/agVgDiW3hf1
PABEVzILXLd6qu4N9fJct0s+Lzclx17+hln93yUz89WPUjwBPXMrn4gox0XEhcNP
Cvps3ypt2AU7tcNZhjO/aNDNlU5hFzkpQ8TiZAnfl1Iqxc6BugIRV0Gb4gULJArN
o84C9+U/m+CQUblkvivPQ6s4t2JNxsVDJl0Zuja0KlL+w7ecqyocrYt0gPyPuusI
c06ovujSEWMUh69cV+VQBEEsHV+t/2ngKQNGw5J9KYv+Znr9ZyEWquMlAR7tMgTN
2bOKLhuU8ThATMY0cNujmYSADUb7hmOPPv1ta+UBSKGt8sz4+Wsku+0XcfBDRCey
ZJSo6H/Di7z6ylK/A+DdgiNlgcnGA0T1y5r9OhVvkqu2NffZhUUZVbT5na5hIHEv
82SKPuODTA2FkoGaWy6E+t4jTSiShiuWbWjUiR1a9KT/GusDVBswX/7WWbdyE7ad
c7Wqz4rI8uxTNuByzayBZ5wE8+0aDVhZiT86AtvFcMP3VSe0rQZYnTxfvTsSWnW7
gOds8e+zRfayykBZo7lKx57m6CQseMHLG+68uPpuu3ZY6UcCkjcDq7C4/53bTSAk
GyficyKZjT4WF6vMkyVDCXpna4jhVoxuoo+CdVgPThQ7FAx5/gcwsQK5zaJqUYE2
jinkZ3PHOTKaIy8KTU+UbXx7JB+iWixE7PfACuj80SDxOKZjShfERxxbQBpHTsCq
0hSylJPygyEfHF1Z79vuWOaw+oXVpFC1Ys9PzA8DwH466Sk/ADTuZQfj5Fkxto8w
CnOCwbEV68ogN0HSZL51PQvVWTtyh7ArWmwmKV8tRknRTpwCDYiDVIFf1PhmGxqq
WN4x7jPTtghvXNKFKsLh4zVlSkPdkKoii0Ylq/9sfw6rUsMwfXR3DnfoSV/iybHF
Zst9DCqOIGk7pO3iovaNSxIdETAUmTcNr3gRmnjcAhvmM2JtcqQ1cnTMJjXVEpPR
UFSJFI4RzrJqKP7dPBEs/7L/oIP3dRxIdkXHMC2ZsRlGc7+9ahSSUg6FXTfNJhKD
x3tUECanGLu9ahdahSnq1n31NN4jewd4UlnTMue3oNK0TWFWTq4aqsqVqaZ3CCBp
1+fy/EoKLbD5nQE5wPKTAFfbCWQiyNQL1VbXMMu/rtZEswEAO3qklnb44qymvbek
jgYrNc0dy40IjgZQQC0OSIYnTNMT0mYMPOiBqfjTZAfyjbhKgTXaQzWxqauFvjZS
wdST+Y+j8VXZ6LWgruGAEG+g9nnGbURntkXVBDSRXlajMPJxyPQq7AzQGV0WZugi
ky4NuPviFImL8p5R6Jqib/YOB0oz1tiwpLyf0ctufGIZyGMu6/uWdrVxqdlB9U8d
TWF/36hdqYllqEVOYhEgbsW1y4S18xmY6mIPcgLEVHp+A4rtiAZ2RiRLYbIZQAkR
Rkskrseo2XcfTA8bd7g/ujY93vfA1R5ftWjhxyCfzDnTKzcsJo64PgLhKq0K7NXR
uAQFDZva81yGPZNPbrGkf5cuDRb6akui9o3OwFMPHy+3ttUUgYqN7Gt3IQQRsbZD
aYS/warC3ylmYXfJ3vrJstPkTeXEjHS0q69ji630SpVp46WyCgx5MDQrKt1Z7cxO
miPkhlloKtUMoA3rAm6bfNGpbC4NULNIufnMzDEU2oFsE4+/GITDnYkNnnzQoxqW
1XWBuc4XN/+DsuoGAKObqjhBZGfkHKAPlg1HTpoG20PBmJ8SufC+ItOQNwCyzZtz
9yeug84eXeVoXec6DSgVHrFGDJrOTR1xnCiXDlXPdVse2VAUoni7b2/hurVSCjyE
RyoUgyWXheXPfuy2WWQhIHm85R6bA3Ifft4dJnn6p9nzM/zEVw2ZUG7jXMZAg8Pb
xUABi5mg5wBsJPhmNTb6OrM71mrzzYhRCEj414LavkSJuEIomTNk8PNVIFqESs63
uPat3CmlQi4lJMMGLChLwJlLsrHEMFmY/01ECJwWF9dSKpjRHGxC5CQGzlv0elIi
rYRj5zG2U5cAvgxjVwPfJoOA1nuy7/iWG399DqCoPoj3tIBRgeNZmVbj0rPq8nMo
5lBv8LkF16Ak25UaZ3TJ1+XTbZPcmCesXxib0b7iw0j5x6zRuBMPOV4oRBnTjby0
aSA5kyqV81rVqdyLreFt9Cyalwk+khEOAlsDLYhG6wqYQoFk41X1PkXHapozfVwt
n7c6Lcu0Nb8NRBAsdNXJc8+weftgPNGJA8Zhm4RcO8N5cKpPR+F643q8zT1T1D3S
/FnnZMvsbCXATTSrD+2HdCu5OIKl229k7Z604ui80V++CItI21HV9L76ZBNaAeHy
82nbiCWagzQG+qJkIinUvbRLr6B2migXNPoN0aA8Uz6xQ9ZV828RZeYCGVN6YNk/
0YxAdmol1obnoNbLAZ1t5+pq71a1ei72L25ASV9EmY+CMnReqGA0X1KBHdY5tPAt
9xX7ahkbQgZsV3DK8aFfS0nAIEgion8rTPwj+sUB6TW4d9B9OpGtJ+BWShQ4jQl8
/Q9eUFUxlgDAWAAV9CaLn+Bukl58IgrbEtIOChIy3yHSOLQ0ZAa/1eOICw4VKdsb
XCr7FDpG3e/BqNn8Gls2UAO893wJwUoN/oq/PBLQw19WUQvsTHMF/XGzD1GU/1LF
rBVgWaz5CuG2RqtChqVgIZmuuKeqYggI0KD7kV8QJiq7XtvrBap18WDDkFZ204pj
d3Ky8+sbYzS9Nq5thqIxtEJlZk3XCey6wUo8nAIqmkQEKt9bfmTp8EhWMhmtrDO/
Ub7qcLWKPbi9ol0zXjSKfb4Jr85+7UjgAqkLETMfS07WcsZxtwUG2uw2vRXibr3N
prvIfM5m+D8DXvmuVoimPhzhumGjamMiOIy9Hys2SNV8BHAorazZXZSgj/Upq9OU
XdvTUnmbSKNBeOsqg289kQFHxitd3+fMQQrB3JS5336+y5ynfcXQlLQwgNQy4OFm
l7KhdSDl4UhCNtxF0bSa+QcNy/7ZqmCRH7sxAe7PfJbe2EA2YZpdKiXpdsXAjeJ0
MV8EhFyoazLNCvagXttcBBu9pTKN2/aW1fGEjWf07H8mpcLl239dwpYQBWtoXSlq
wA/w3RDRB4CE8bLx8vrPe/3k8eYG/gQyul3+ovoQQE4U4sySyisC5JE3YJVRM017
rmdZXgKGxhjz6ZoRos6j3/b5rXN9eLaopbnZH36r2tbDOCkcyJrXpGQU3cV2gieO
MuoCIQgmSFWCPcncmBqwqPM9ToKX734j2YCTF0YrrPAfcCAe8IsMh3yPINGcYTsE
xx0yW9r/Y1wa6rMrC9pB4x/Q5vL2Qx2UBSZ9Jto1qGogi1COmTeijhJHwH43tDtx
6Dte/NzzZIaThP0qYd5hT3Zn4KN/HWXjRw8PGfsZMbIbY+7Y8PtlQGYwZ5e7reK6
8WkrX7yO4XjL73rQzieedG4DSORyIzj1Tq4GjsAbdWhP4H0aVtjh+tZGdmp2ycd7
71UebdFhI2P1VOqBVVh43+rmRLyjcObCdY914yv4UrwAqTiJs3Xs7aSb5JRLYddc
8jMYhzvttGfPPgUwgFjM/uAHmtEM8V4YelyBAgQxOTb+ci7Pa8bKeyBPXRwOOkUo
DgO2w5BT6KlpF0mno8+Lbdtfr2VXTaf1XqQNS88IHfvNF86V0LM2B3iL3OUvAp5P
MBeQrUan+dEYlKu5/LyOFcg5rCeYPPC++1KHpGIFCl1h+cA8AOicw5XlgNbh2kJk
rxJ+ov8xOpK7xvNr/LazDwpDpxmSi42Ruoa+icFwRokX8O3bOuNtGWrFM5tTcHBh
7TIf8BF3pi4TTnByd5K4JTmigoOkSH0XLVuPYWCYNWnwLHtwbV1j48vKvcSpxMKm
8wpgrps9VkJE95XIFxHUWko0MDedEIEuo8NElQ0TKFKPQ3oAf+531hOALDMWXqXZ
5MAgT2JdrzHzg1yrwoSfqOoMMrC4VJ4RwUmf4VTNHQ7wZS8Z2L+5n48CtwMeN98A
iAM3u95Z04/2jRmhapYLoDgGYvaov9PjabTj0EiPg59h/xfyxtQleMb1cga2072g
32SLZY3sPZ8RC0GDvGwkmGMyuvEYk2MK3jVg6iWT66BgdzwZole7icd9Chw2kMzi
WpOb4c8d0eRWOJdGzR/g8Pot2in3ZQPZzOwb/FZWiHfKQsJ9WXM+EDhIcaF6Tup+
Jm0lpsizImw4ioI63lvaSirlma73me0fomsvCKBXIapc+iuvemE7PJXjqoJQ98ve
OPE8TYSM0+5PDygFakW/Rt0QlIqLmcnnf0yU3VQk9EU+ysRMqNYxmJbpELDDsjs0
MGCgolmhEyzaggcPX/LSWgCWwcGVzvbQl7ZkGhBlGjMONamP9bc8IRo3FRoqmJGc
Umjlu/sNjuawwyQnKn5hvdilv3bQWRSQnZ1zlcvQK0YSO4IUhewDhlK9X5Aqb5qU
anjfgHRYLWpk83QF0WRFKyKztM35mCQ2zfqPl/spjZ3cm73jwb2SZP7UHtRBueqR
Uuy5uKgn6f3kpz3iWzWqSB/uWxy6krTRJ0JloXtA/1COYi4MX2JoL4syeC3cbvJO
pcRrMO2RRqHDxE7z6fwEI81r9tT/P3Kl9cgCpPwgfNcjtPsorEMhP6tkW1rMxiYK
KxZPyKEvGr7BX4G7/6DCfc4BxUQZfhu4OBKHr1a/3wbPqnoSKpxKKRxRD5QuIbPL
s+jRAxRL0j4GFQmVdAOjMPupRrnwwmslSoCop6wHiesXpNOw0t2r+rTCCy2D1DTb
cWIYBRLbbQyI3rUTh+4TmhBQnv4DwnPBWtXfqwJsRZSMjIUNvIFANporC0Zrn/3y
jMUEyCt2VI9hvBFdYLSRWJn1qxWG7TFiGXk0WcECC4pwq0A9pZkXS4rn2dQjFZq3
C7s0Etp00XsPv/VXo8fcbP7Hnn3ysbsFHLvJOczNqAMLtOr0QwvSccI9jcAOe3nX
1YHrlKSYAU3sE/jUQH6F3yLAjAqG5y1kriU9Thvlxw6VaserfRBgVIO/bqLEl38T
UYkppNj7nCONbYWEgGGabelD9jrOBR75gzu4U+YFoBsLVK71DBCUxvRMSabL2Dty
V/xLIfRx8rP8uuNdlkWMX6HnC/77O/7zUzTVJZ2eauww+tgrYoy4GAQhM2o68gnD
vQrR9IMepTlMpvedcvTh36jCnfSKXXIbkbbRsqARNDr1uDGuZNNLQiv3hEdoUAQP
xqr54O2MLLC3prTerhoPRtJnT0LEvGXOWVjRs3/Ff3EvFzVBgV8hqdXj1b208IDX
a2DNvQkaWVfoNQLNt5Pie58zPX5aBlYnbylNmuvGdEf5VTZiYXzeHmbQHrMQQGDR
F3x7YeZVpzrWC5R3iwpoaYw+IKhbGs31VUpRlsnfl79koMhCgm41Z9LS6RzvKQVA
UzFExZI1Alnca5Mlz3XfTe5DL3nKFPLfUpQBMfhRUGE1wn69kkilR5CtNXfxu5f2
Q+z6lKuuSzqq//lF8GwYOCuSvP9qMpJWYo2UIN24eInfKmKtzCB4wMYOkZ6z6Dqr
nz6APLvTUvpY1VlVtmSU52xTNH5C7jNBRnD709bWtuaAjCZWrX/fqV2Smi/PRx/m
J8dFCitW+R/1MItbM6v8Fa0H9R5IKcDO0YiK8WzdwnoD7TDfo28hY1haJ2xx9VC8
D42heAyDUpkH/X1ZOMogTgtyk5oRG82RNXxj7pddKmgSbFIAyvyO/bdDGp6M7ydS
n7AJcfybFia1YtnMLQeXxD1IEESA65Sj8hC8PW2NzRwo7X38ZY+mtO6McDBY2USN
5nWBUBTrn5pzZRnp1CtUhFk2W+YYvGCPpzRc5QF/85e9RE843ahP0b7h/32e3ULo
LIgHIvLhQYcCR88IiZ4uxCxBR+uf78bjRNss6HRZEiHWFeQzC7BXQdYPotg/A7U5
GrGj8AkrDbEEL0K+mC8xKntsNc/9HTGP0WjNL9G+3TyLMHdS01bsWH9O38NHUdJh
v64sOD7a3qqvkHCr+QASSb+INwuw0+7gthZmo6HgQzGuEYYhBbtwHgK51q8+qdxU
szHD8vuQdEIklQhzxR6de9skkrEzUaPUrFRCcfEU3UqUI6dSFU/QKaqc0lGahJow
QiTPaMUNghwFTt/DLfbOQ0VxFg+iTFNzK+H7NZfu8rvsnall8Km+RcLbTIUhpOGt
KMqCBpubmheYiQ0/vliSo6cTjlmcl88pyJQ9BROS9WpN0hIh4rombaA8sBvGownO
wIfaUUItcV3Z3T6aFjVePPxeaxHrzcIJY7r7tBw1nPACT35KO1AkMePWkIOfZ9sj
vBQmtkXhPVTRTu9LHqctWfyQPEPdWLCqAwu7OIyaCXR7aEpPR2pk4i4wumL6zDVo
tYfUNIxRoUfYEPuL4VlhM5Z3I6uH/MnS+m+FD9XRfijimeSe4MEHayxOl8ax0Sk4
Lyf/DK+MbKhG1A1EvJVtvPU4Z6bHZmpWI7ccztJPmjqrBlKJo1G8PxPENbZCwCib
YvAYLfeXNkMwtloXfsuvWrJfZ2NY1Ef5/N7ECNS9YU74UpoHV8pKcM4XqUdDQbhM
29askQ4cZcuDihb+YH/E0VAo/2beLi9JuZOOKOfgc/pIjsPXMPBuYwH1Qbhkh0F/
Oo+1eJcjWq7MNTTyAEfVu36TOPW2kAgouXLoEj5m52+jKAMdp/XTU9ZIClYk5ZTy
8w0DvrGUK/IgCRf8tymxIniCwTB8oRT1aIfMR9O8GHeC6ScrotG5cNfnIDNeHqXH
ELQCzr5JAUqzHYuClSIJITb+ThbxsTgkcKD7njWSGDONTrJfDaVE7cVoJJj6sRYF
uK5eVcyAG8gc7SsswASqulAbCcNYXaOjwocpY7njr1H7i2Lq/idIbmkIVlN9zn/A
bFaiqUvRA8XZybMcAItST02D7WAwXoAlsKV+XLPiPVBCWA+WgTOO8wnmvsFHlz44
TvQiIUOuD1lK0pgtGbsheLedj3+0veRW9OSaosW3kKk9LiKB8FG0GNZLpcDV3llY
7WJB3P3GobVDPXqkciagvfOmKKJVTlsl1c61vdTEr4ZdpvEItQgmluEHTzZDo+nG
FBQeEMX1Ws6YUNkRi4OYgRDegdTkOFlY77YyQcFarK98tVaORkkwqI+MB4xsT88K
dAuX1rJCf4eV3hHSMtZWqF4vOFpEkAc0A9YTUROmDXFippNrXfR2fq5hwfHdIdgv
3l4sDv7Qw8xP9/jMwW7GK1ovREdzik9CNj4Z2cJw5rqINK9OFlTIGJEaeLDlhYU3
Rxy9aJhfJAG719D0FMN+/nDb0cP/ab7gwLK7xNqlaxV/g+MIdME0stkm0spsyFkv
EEfI7TA3zRQpBf8/xQziqaqbldgnRpR7wtkdWuQvPpQj6uhMmVCFxUk3YeROM242
yuRuSU0RFpuMITD1puI8Qan+81iaBUNnGTCkSx/CLTMiVde6JaN+bXg+dO8e+bJh
SycR3q4Jk8yWXB7CgauuXieM4X913//kyVoEoGoALAtX0EfvKVYEC4h3M4RFHQc3
tM/SBg+qk2MigKaWJ8I5kLFGkEPbchARup2ur1QcCwK6Sw3dAfbx8bt9Fa8ECth/
kFPRZIBl/TIciIB/+8OL8UFxRVcix25zX3CqNfackM7LfjabNPm4tZEQFA17hFet
Gmu1Fb5gb5BCqKema1dVXC63h6DhJ90Wi4rinqkaHbswPDjLGDC8FjSw/peKP25o
vwb59NBjNwRC1baAo8FEODVM7rPdtade/3CO1Sz6iLsRAlFcxGT4OiSh+nXhSbb3
1yUV2fuA+jYcjNwpj1MOzqj96eMXtSaU2J+zIcDldPksx9v+YGx3VWpkGLo57xVH
d+yiJ4Z1qljgogH9+4ydVZoGRSLKDPSETVYm3q8GecNdB7KrTKS7zT7B9XPJYSgy
RJ6g6M0puujrokRgLkk6JP/vXPTFTISBzxqsFn7aYzQkmfxBFqRorYyfp2QYgnvT
ziecTgjk5oi6gOelgISSsG0RiduvLaGF7TrioPMYMsbBGS/D7zE24nAH8+vAL3Mm
IUPGEtMt2G6ZgpI9b8e3jBFwwemkUFtvoFSuf5RlKkVHm6YnJv8V5T0+sjyzpCfk
R2BeOs8w7DI4eJ3AE7QXxUTuVZYCjmTnkP0NilgglE2fbmDBXWmZVBRa/twHmhfH
PpI0S3BcZCPNQDd5kmYjGJRHKMpAYcFqDAjps4CEQY8r+CEtWKf5SmPms1maIixT
GYGnVaW42nZycOzFgRMQOU3Kw8BuF/BPXWBIm8y/nRjaiR9hbFSMVXITLuZQdQgP
sb8/IU35gZRMMuRUp2R97pFLsTdIMMLsbDVuVfmd4ydRF9rbRqypARx+HF5TuwLH
EtMJGig/jUVrC1oQEUVGHhG548DB9ZiewQV1QU4NuKqKMx5us5/V3MDfR+cjKcHh
Os88oODwCJ/wWRsZwwDAgFuMjpLDpXrWf1798GVYsYs1xqIq9VSgUnMJxbSx1fi6
XwOUkzQiEaArZ8ooMoPUyEMfJivGpbciPZP/t3dFuG08AeKr/z26MW5qAK5Pjra2
ZpQp2jXOa627/5CLX7dyZGvdYZu9GhcvnOh1b3FZoyFgffwd2vhif6DkSa0/XePX
UdVSgADx3jcwQnu7mtC/AQt79hmVvN4qmRT6BEZSjwO27L+i2VhHBy8TdLmbTlpZ
TYRHPYlKFf3kYcBUFeJwLVAXPluESBD+a8Cl8Ys8KAIRHUlzb+be8WOLC29tBy5z
uv8eTUzI0M9IWmvKpPLn6l3Aoc6BVu2YGRKvPA7K0OGZW7Yk28YF9ZPW+YpgeQKT
VEcl6Y//w/dR8Q5k3rl/Hbre0AMYiJgsHgiHM7r941M6z/SW1gNMVIgPz8S2sYBd
nUZnSIjAWzfL2Gfb39AF74xelEzpqM3tvV4Ziw7kkPYkMag2C5HRuTPiAjbXOiVT
tSzGXD8H9jWE7NmCWavk4NeMOr6OSC/xVfS58iyH0mZgRpTfbvO3oGd7ugKWsDvp
Z3MRMXEvjz6yThaVmVgE81Kjza+5xJNArW3vEIQemyaO6TwzJMSO7uUQGzU9IGOP
K3/AAPLoJjER0BVrMcGLHTdIg/zHMDyF8st2crPVJlpMQfdwL3zMhT7cZBnPWR+c
4VkRMPok6soVRaAKDEwWs2F28nY4vdMK2y9mX8iWjmAmSXJMebSZixc85jBohe3G
55ULeCZXX1xuQ/hrAvIhIyYW0VVyrRVGQ4aroq5rrdoW4cypSnSWLCXdyUmxOQb4
EQzFUJLYcVMM7eYSs6TtIwDlyCOaUlP0ZMukmA4YTz41blnby6LHcIr6sKtHC5HK
OrXS/sqGAkjFuLcwDaRcp/ULn3yQP+dOYFMPL9+suR16GYoXJL5/xcoaczlkb/xd
1FG/RPw8iHgusAfpkU8P1H902xoQ4C7VP2YUBh5mk5219ZBR1NLArx44GJOZFHn2
oky9owYluhziSFkdN1ETowqXhhZXyk20BqAEqAQmprTW5BVzHZNA2s9JCDqffRoh
Fojb//mOJULT6XTctlG+niwXi71CYTMgCmLndMj/PsWSoSHEIZbkn3ZPQAUZ+rzw
7UJ2sONE9lMkrPI2KF52/6LOZ/coPRX8kyhFRvpC24qHzKRkZvrtBaDAqLzG+0XB
8rV8qJosuoil+YkyeQznQiclGyvgcJUyaWw+otyNBTmvYjmy5KlCAikVVPefX8x3
945DvVHycyAYENWYGqeudSktiKkPF6Vmp848xyIVBv4g+tJOuczgGvE3H4Nwol8e
oqh5gWET3hjQMMijUj/mNPMZXYMArndyc7EatKj35BdGOaW3l1TUBUmU/uiBG9S4
u6gtqzRmh8HhUAg5sp8zI7lmgN8Pkdc42vddqVFAYIsfK3LjTdZB6jZt4h603U2/
PZ9tWPZOKXA/Zf4F4IuM3Z5aqa+o/g2GJn9FTAz7NhlKw7Be2MeC0y2ju3pD+rFM
qlCsXTStkGNnDZToKkCBgm5KILN8RYq7gf37D1Lb1RPAs8Y2EqPXkwhzUUA6Fuwb
/hjWIB2mfo1mDdpjXD3xas8qoZrZlSoUYmPqdj9Lqrg7RG+WFmDb8TgBSPLLZm6A
r23OhAfuZCNt0evsjniDd81KepJ6bT2l9lNVC2mSdw6pkxVEfaefRzO4QBOocWll
5XZElJ3QyYyosnGA4lMah61ShoAO1iXe9HqvLtweHanLAhWCuPG4xARzNajFgzbK
ngwik4qMBDVgG8cN/JAnqYoTIBGGemBSNjLOVvdK7GC+Aj2vwBoL1fxFjhBxJ/b4
ZcHe6tGvyDFgRt7TE3Bt8i5CV965PuCaswGje07m4htbcPoXxRhEtbBzn13UTWI9
nl0LZjp1DdaXJCyQKIBJkSgJIVVrHewxCELUwNUI0wdEIl9dmMVHq9zmEL5Uknwr
N1mSCRaLfCnILad/LycIlMPS5pOzsbMZPRNu+eBSUfAE07IAByulgF+X8OPynehz
2UbTVaRyNh/E5Qe8WHaqYDdN5PSRiVGRHfTu8XZCMtAxWhEf/W6EQlh+/tQm9jS2
sBLEH6d/tJ8yoLdPe7hb/X885/8uhvCbp010g3f0oxY3LwjUlrstUw8oFqK+lBTg
/4hwX47Sw6XDw1V3vmTcBgxL+O7gNWY3neLPUdgp/n021ZNN6G7NCIJ3WH8nyRgf
DIoeVjk2T7ni2YzB41KKnMuMj4OT5p+QJHZLsp/ziziZk1QT8Xfz0WjJkRtfPEKL
qec12HJZovBVgNpaYDZ5SChnlzKd/zlNAKLaUmx2kFg+x7jL1eIVOCEwosL9Fx7a
iiSUoEx15S2DPIqM5FtS54kY2LjwVZdDGM5zJiQwAimsacWFJwZt3jFhwB0VE74f
eUioYFqwixUgb4ed181AnSJfT+Wv3LWupYd1IDu3GTbAUUlnnVJPV86A/7pYUcGU
IKNokttDhe9RhoW7306uO5TOs2FR8eQb7uqAyKIHV0K5AlEFUFWjkMRyeMy95jc1
WL0iFt6KaurAsebl9Vg8eXYMLVQ8YnF6hSw8kxSHfPjNYv+wUfRJBWrnnXnTntaq
51g63oif2RP0yeWReGvPb2nWAAk10UBpZ999BJJCiDaHvsACzWEwzRvRAGVMx5N5
217tO0TI9Y5x9q3VqSUjIIZE2wvkOGt1D6V+ifT923TXvwgii92eceYWtworkX4g
MSM+FifTDSlWl5OP19iWMgNVu+FspmGoQ/r2N6EmdcH+EfOdeHA0QBFOiaqIYAKB
vSw7MUjUCzZdzCKxIiwgtjnL9wAjN1S3ixLXVCvykfhN7VocxWlnMIBCuKApWvvR
0dN31nB982yGtdFDCD4r0sgoq43PsS1zk5KaBrbTuNjpRuymaE6TpyNIDZWOgti6
F53x5OKPene1WcsCjz2FUObyq4RGm5HQK+kh5F1zitktB9qUwT2MYM+3lEoz/qwN
g9Av1Ld2rCofp+65e8xg/TRliex/sEjiyawcrAX90divVHeAWunsULW5EQO0NOGr
TzJVKe4WdrcFKVmYkPQYsrTjewLAJC/rZUL88HhUK1XuHxcV0mIW3bs7ZOhkORtc
0qsvsYgmMWaA4r3FeEUpLUl8KAdGTwkNb3HtzmdGJvQ0bRZGjk5VY8A7tVTrhSU1
IRyi5+LuK86/KMuEok147SfFrz7A0xrky0kcP+LjKJP1azUG6xugjoxdorXL3YEK
h95RFt4n9pkEZgx5d/aEp+VNYvHoevkIR6lIsqNVheUhLcB9iTxvXCo49vxuBhvZ
h+thC3OcbPUWQDQUk2VYL3zqmhMoQPn0GAwxWUf/+QPKw3wBFFwHeaSk5DdQ1Xn3
YqqooZHnZnRM6K4QXKiZ/GNgac+in0mq/QzacakwQV0x3mB1LVkLhyDnrJEVrSeg
EM2m8+DI75HG2SFh4vxUOCe/VVT192WDqmtJBGI5thT+sI3+iwszzLaKoe7jyia2
voCiYSuzCyfhCzP8Qte0dCqeZ5+XZrYbXY3YEAIruBT1/TIDU9rOoaW/VOBUem6C
x8TKwhvIotJr0hnctetXspaknZQU1B8l58h7TL9tNwB7RKjttvTnjNLJFta48d5P
12M84KHzYm3qKfORy8gYWg/4qfJOP12vlrbGyvfak6FCFWnsjhpK2Pu+SCY3cJ+U
xKlb8Tnkymf6o7+Pnlm31Hvr0dJmtI3LmKSoFemHt2wcMGhYoSII19yKsGPQDLMS
UOEp5TbpZmWTNk4KC3ZtE3c1F42Bc57AApWzXOKw3TWPh7YJRTGBraHK3Us99Iz6
LmcabOsDrxgIfa3OLbEB5Ic8iG5CRZWyQvpKb4jbLW27yionu+ydYLgx+a4o0QbA
fJg6s3Aac9h5Zq0irvkbLi0Ur+VtewMCRgcGXQlx15+hOSug7R2eQD0/peqPwCEm
cX/H12UghuFsjDxeQObr7kQfzk7EESsbFQYfkiJByl/Pgxn9rDskzSdDsgyBI8XF
+qtXKlAw4bKk371+v99ujOuWQdTe1fXDIkCSFPduXRC1jCGoFD/5baBsXcZql8jA
4JBVus7RQkRajpUAHxiMexggTJRg2xF3qBTniqxfbsvYKqXf/RzGiXEVkNDQRlTT
Sq57+oTQpsru+UhZxGhyhx6eUQddNh+luuoIMU+ZXU7xhrQMKaoY57CDYTFTNJ0H
16UjPPc/wVCfLJaEUWNAkKpzvSPsEQyevVKG1L4omXvAS+01CW5P2NX3O4Za6uCB
jI0+7cHYupjsZSdLAB3EKFX4yBD1tK3pIaZrn2KFHbpF0e16jSlpsvJvhMrN0Uli
7bKaKNB3VEmbKc8fUxExNcAaKSnywrlIGeusd+Ksy2Nn6qOLC9b8eXnvXgqEZF92
guIlmuPDG/333TnOec+XUZakExywjsAUJDrzTuMVyakcfSH3DOlg0ua+dM4e+m3B
OmLZpDhdqKe3l+COVoh9ph3HyXWa43KLWByBEx6n70cYTbqNE9Ud7knq8oCPITy5
iu7dPuaZqODx1SaOml4FQvMNxh+EXJiXUdFvZOAo5RxlLxSinXlcJA2D6BUNpEIW
iTGy8sTlqmY9UJbgBMQ4R2sFJJWdvBIM6Fk8vP9cR1bMXzsxq7oUVNYJdkavH++h
ipPz6puvILwoL5WY4Mq3VZywz04lYmMLZlFpndvUJvYC7fKvu9yt//hbpb3vic2X
zXSX5hsCUKslPwAmB3VTiRZvoEnDziqbeJfu4htYiZa13pXgOCumQ4ENs+fjsLqa
IRHpdaZZRiEGmpTLWuiQe1xHD5TWVG8ldIh/5dQSVlEF9BexnFeW1T/3KNLZN6Km
Kt4Szmro8zqdKasxb37dojufEkxLx4Hmy+c//zvI5wKeuuhwudg3xVpfgcMgQpJN
ZIAY+S43eOZ4PgfyhDSdiU7dgos4CfNS1+HzvzJs1n94PCI8hqZYdnUDAf0tpTfG
AJ/5c9JWOqxWp5A/xwu+Ex6h3q1b+gt5kiL7VYEmn8NFZXscntE8JIXrOm9Txc5e
+sedADc6O+eI+h4ddTzpzXKMhAfhciXWsPi+GwYyoLp5MWpEBWHn9IjYocjbBUKB
L9m1Xyph9ir+tGkgobNxKN3WSwfZUcPZ4B8y3JJoIwxPJhYL751cd96PWTBMucY6
oh233eS3zZW8VAbIIb3loT4Xwo5AtYLhPAS16/7LmxIyJuRf7EkPaZuoa5KQtaTs
3gxqvyR84V7CbHQfiN+ZIt93ZgEtk/efxGAFu8FQUCLKltOxApYvYAbjYO1XUduf
AWyJ0Ro1KXfjEdlSrXmGQNhXnb5Zl1Yz4QVgKRh40fPY3Fj2NUT/RhkAmWqGDiBE
AI5geOfYHQWmKOL2/4Yrlhmsoha8hcDje4JJ2yQ8vsivoazDF47bQHeG7/bbxAha
ggCn5Wh4wMjN0tK/Uf2yurXBejEgFvt3rCo/Zb19QQG4msqOc7Ugpz5pRl+nv6xB
bhEemzmJNnsBbyCMbUeAX+/GwQ2fOL7TsZubLfHb5OtntR00AXASYYLl4oUFO9LG
3O4WksrC0kPAAWXgmcuRLPM6mFT8SjXs8OM412/jlu9KDLpShoodsz13ITPDu2+0
5dlSo7bPq5t4sw7UHjXL3GHd5lRt2d5ItIwUpfASoIxUrC7KOzQXYci4AhM9CWTi
LltW8PLe88zPerCTakjtHEtO5Su6WRFL93YNhbr9PEnPkaj4g+fXR+D3cLTeacZW
gMZ4RuzES0mUpfLTWMCuFlNVvgWin3jA7rSdqJ2jXQureOS/dWTMC4arxnPg6Bzo
VdlPEjY6Z8HDCwZwDbEV96IsoERXSPXIKBdEUUrt55miWc0DNa+hJZAYt4QyK6VJ
neYdqMete6EzaG+Mz9mKCDvvsYOS2/nxwesY7LgyDtoe9M6KSDM2NAc2hs0zHRrL
uY64Lt+pTqo9XhBytqwLCYF8QjSOJyFPZf3u8Urv1x8wTQwXKcAWFxCpAfLkMkfG
NBt342NI1KjZit4slw9VRRcnRJ32Ob0WTm8s4VegT3ynbNttlAvLgF0mwKrFEG2S
yd9uTr42Lliq2ThaKZLWRDGT1pz9IwY1T6uKpVOctSNeuzYNSIIAXUlIKNZyubgh
1gRTuIP73m0+jBIWiTcVNffs2Qdkf2sgBcV64VWrBwkwraxlfxNG6vfnXG6Pd6hz
x42JP+DVuMm70ICH+VZLQZC8X+biwOcKaZCIC9N9ZdgFgkg1NwuDUJyLBHJuIzyg
2oGy+kadtlid7qRiHKJPy6ocr6h7Ty87VO3L4mlJ7Mcqgmfn1h+LRkDjp8T3aF3c
D4EjXQofft1/s+WxtQxsZmH0qN8bQr6z+EDzbzt680AV4P3weArV6AaGWtpCTO5n
Vw7FMxjA6N4Q8viAOx7te9WU/pHRirEu7x1f9cxtSCi6mK87psjJsH0/Q0jc5dC6
iIta+K6rhCaHMpK1rkMofMvFdpRk1zTadAJ/bpUAfyPJbMn5ND7YleQXPtyo9jh9
M6sUrRwePwj9GWnIiDTw0fgSwu56M43Ftf4bZHRlpSyGiOJz3KOt9rLsieyXuFyH
p/VbHP8wkAzY9w3TW5Mas9dK/IheE9EfbnlTqgejlOIUL9PjkzklVZPx/rKsRIEL
bc3kQL4dU5vBxj+mBkyOsDcLl9uQpOSafWakS/Mtq34Ycsjv6DWMLT2+nJf+jVGW
vw9OOw1qp6XWOctgQmJLCm9e0qHaBajKc4ZD7Bnr06sPDtz/Q7NrElE7mIJwUZFk
WBKQ7a9kTl+uDdh9mM1WdeOz7qJjy9Ei5SXBiZoDX7mmOAGAz5UltXK9YOy/MU5i
lVjY0buFAIqPi6eAEG3T+tn0BojA9EcCpdDRUhpg7+Ia9K8aRWW3kuS+qW7ImuTW
7K3eaTxE6sT7k5Xva/LljsBpjTx8b2Ejpk6nKqfj4x3dzT8KELi7oE9lqU0hYs6p
frqmLjIMZp2P5s4yKCSi4oFuucSuir58C46b8j9xAlDbmAdhVnAGNnCD06+14ppq
kpbsT1fgzxPSrmhUcq8BtjHrsSjq7JyXge3NfzOLg3rq0f4SGyp67xv4pllQB8Rb
H8PuFKlLoC+LuvwK1jAr0zPYiy8du5vprKhG9Ayg+RVrGcH3i6mut7qySIEJDMCF
p6eopnPmyiXtOxSdnrcgZH+M8keAd549blStLLV2Z1KVhaPHk4kJFVSpvaMzC3pD
fMIWr0wE2/8XneDDZmPffyrOpe5LqeVvR/K8yJSiPb5Ap/LmXHBZ3jmrAUnmWnLW
h7MOriR/oRNXfWfhjasZ7MVC54nIckdYDPOY6S+758185ZNtrlXME6rIFDlKjXQm
Tnxdis/1/vtsWyIA10zFs6xeboxdN+xVxamMFVK92Ln5Ay/jabMTW81BXwxaBW8i
buH3C/hSnGcSkrQsPrD4bl4SCR/S2ws0kDoT1GXEOLfx6mlAEeEXeaonDW030Kvj
Gyxcm/7/v7sojMeVt1pLzPUqHq8lQWJ9EThc3wnMZXRSfPBAVQDZ9HEHj+aqa1XO
hhO7EfLm/n6uazh+K3nBXmI8weu9OmmfhhGhwL+kH3QQaV9jWLqeaPc7dEwqOfA7
oytQVYv+uphOm6ihWN2K7ZkR9VDM6xInPW8Y2ht5GISbwm05Vl+bkflJvt3Dsq2A
HhkBQYLhd03Lc5S+peYkU8r6GJQwm76lKtD7tkl+fVQvF4JTjLHNtxVnDZRvLd7e
1pmVNjvSPQ+mzDK9XqyUTnY7nde1GSO+X3rA1B2ix98Bzw0Nj2is72IGc/O3BSRz
UQhf9dmyeEmHa+sHhx0b9GFstt/YAEuSFqlwV8Wsc+Qozd3KkxSSxu8LyKrN2vbk
vT2dhHqF0ThCnMJPTbjxUTGpXNYs5K9w6PK4JiOWaPaGE/blfWfHMG8nfYI+SoP0
76fjCe9TKAlo8SQDN+J/kg1CesPK1oBkrfhK/TYTCP+RmNjomkBjrOUZnITLyRhr
Sekt3RnNTE8dguxl/yUXenSfVStTEf1cevq3MMXkVeiJBQFFFvdWM4t8jjJR0mEk
1HxjGIVrghDjiB1iUvVjm0bfxU3QHFsZBQZdU2gzk6VPiKTx0qzE52NW3r7vvV3i
KRdGahR3UJjgQFndrE1NZyHuBka0L8prBK/Ryyb2YnPDqx+c1Jn4zFBuRzPVR4LI
UfU30gU8GKR33xD9mC8Rq5on0E7MiQdzYKBdUcpFI8DsT1XuD7AAprZzzQR71E9/
r26iLFGYpEzToUm8Rrenpdtao3bORy3aOqLytnlK5iGqtPjpdTj94KBoSV2BYKyX
JwGzbeB58x3issTm0NE8NrJMMwODtUQLqozxJDTdwb5tXDu6iWR2D8tGMNvNBXYn
+GrHlPuMcOg4qx12WqtUQ3Urc4fyzesklHFzJhCjCQXn8z7EEhJeKIumaY0ltdZa
k5oWC+DWOtrZtIKrMuYSYwhn/usNLrlHsNpQPpQVqxN/rQZzYbjRKBzLsrub9XN0
0ixhghvMl6BKDl7Otq4/jmHgOcoSA/RXDckFzWKTeFS0rpOOn1dLqmTQW2F0JKmq
cm+DZVZGxO3lsGoWWh0pGZ7yVIaEhgPjSZlN0y4GVTfby+nBuMXy+ODVwpo/IoS9
jJ4e98VshAkcSyjSaRYRjUfvYrSRcqWypKF+aCyn9mZU7IexzemC3WcoOPtUCuiK
uq16f5PgGeVp4ITfAlqFY+/qtL5u/CkXJrB2qrTXFOA1eXpi16ZALiTwV9W5ApgJ
33r7TH9sITAKmjtj5Ml1aaMT7HxiChgmiKNO+BG2AQXESD9tTibCKoIlDEjcb6r4
bM4SXHWBSE33RwB0ZnjmqF+RwqP5KXIqtoBNAsV3sfuJ0y6n0xpvWeydi8iCjsKP
7UQqtI1CO72ZUMs4fKgDcDZX/MikHJdWIFHyqOMI5Sx5YbUvyuHdHek36h3v8R0Q
UrM0yuNLrQRobow6/Yrx35l3punX6PtWq49QvW98MAuTEMO22EjZR+kxvnvjLhaO
qltYIDnzSDRpBx9eBZiq/n0zHkQc+tS1ocPdB2sM7HME2tlYeFosKCDZ91woftnS
Em28n3wZ147hppfsTbuV8c4Wy39VcAZ5J7X76hDm7ZDV9kSlsTkrePIU1TkQ2lRm
vYh5oWVNDDvGdCfDqWLivMbOvF1p8GZwXO8k4+efsM9Xu3PMMXummg1tKxZqHQPR
pj6okOWwXZDyRCh8RESSA12wCgKX7dYXgEcxxNiKNqGsszA+YMjMrkJDzUqTZpjg
vXeI3XFuTkKszDbh4zfAczob6U8PE6qRmlGiD0iDdOPIJ+oRE+8dFcoGuJt/OEYr
87bA52h3Zrr9gCgO/of5ImG0ZmtHgKzTPYB3vzTs6mQGeStfB0h5OMSXHahOo0jY
8oT3IU5ftjufE/Ggq/AhnD5z3fhlzqY0BgPqP4/yoDwDZ+ajo6t6DG1ABpn8Zphc
Ry9iZw1whKNZjcU4HLuj+vbDXLnZl6W149g0Yr5vYeJA8BjUIedM+t5q0XiNfwRx
P0HTg1NdwwgUdekcExbFf5N48x8qkFYNSfpJjsXBKAUCdUuiBCLUugvFW6UhkRaB
JBVvw7Eq8ZldgXSyEbrCZb9Ixi9gEQIsprUVvMyVTlKzJ8zyB5bXkn7A0OzPNvem
T6wCkfMYLB3YAAftolStJjua++rCd7WtUer22WtuIg9K6mF9PUJ66O0Ygmb0yu9x
JMswcX8UiEKiMrFOnJU1RZA85+wggMbz9TlYTA/pQ1kT1ufB8E6aBEOw33xWhFbj
3m76XhNISSlkpOOtxwFMx1T3MNp+pe2w/sFg8stULu8w/Iob0SQ1gZPCvDLGs3o8
1wxQAeABQz3/IlarjBIOyliJppT1/umbwfHqOHErOygFLMXCv/bYqwuxnjWMkWz3
W7wW54Sz7JXKq4GcowppmUSmTz3TUARF3MLw5h52smLRzsj/3xhIa4sM3ONcofMs
LIS6kpCcoecnDafWX4UkkaOhnaItIVZ1QklxYZlp72SzJfzPojVyK0/PIzXLmJjX
y9dMeCODsb0cTFFKhqfLsOt5lq9MYMgri1n8Z5xk/5Gxl2/CWh+ZHxtUc88hxvgP
5R0bX7ZZ5zlqIAim8yF568xeU2jG8/EpM080p3nxJCkuO+psbwbP/4svXJO3Gk1H
suLOLicK7/8CZpxoQxcstJF/tS1zjEOtFC/yI3bA2HpI6Y4ASWmm7MDkPTSyzd6c
MqFH3wl/Rd3SQqvGJJfAekAuTeSX3wXBxRHBUN1j0oIDMJ2gqsXovP9R/LceyeFE
SBkdroLfyEST550NkaoiyxyFNpfgrW21pGPogn5yYAKt+/eZRszZqWX+e+Tx0HAb
BZYIiuEsvZXUZMZ89ilPwFZ6dt2Tjg2AEMYq/P1lTAZ+rKEnNgqiqEuJmuoy1qHl
8V6HUgDd+TsOsxmYifj6tepNF469q5BB8XEuOMioezEBwSgBt1tT13JyOtGOJelq
EKYqaGZS5XkekIYtellayNVB1B92teqvvCZWB6srwNLNakMusWW75phqGn+TNX3w
b0hcSCaaWQtlh9pOGxUPKD5IMIHK4s2naN496Lldi1YTGYzhRSomOfpZSRbMGWgX
vYg90esnz1d7nJGSIR7HUAzCs7O+HS6T9tAMoej1WQ6SzdJwkarFaO6McFBE72w5
AVVhjqLG6rtFPBt6UpX72D8hvTa37wzKsb9heOQC3tsgE/3ceq20El0MqKal3K/9
L9Nm07WUlfpzrRCCcver4cWDvDbncgkhft4MuJR9WSdhnxFGEOyRxeraVDpU9MXK
ZzYkvMT1keN46kEPFtB2oiX5oDtkdwvfPFRw50yRNZn3ayose8q9NLi7KntnOEUT
wbsDs5gbdmPIxqelr2UMlYNxiV80fBfERTIvkAHg7TD0oVQxyULBR8U7OUhfiT4c
5pavj9MTmSh8daDDvjyqcmedZTUlR3yHhCKZaGGadRRfG0RNHz8ZCY8JYsrQhiVQ
DgtdO5BO0jttNmGpjjR5cQdeesIiqluCkVhkzO+53jehIwPaxerMp9J3ti4sgHTx
4cvkurhgQI4QCiJ+nEBZKt3v4yt2tr6TuXHEBhemmXnu5kMP0JaSDc8g87WPktrc
zlR+daUXghONj0DA/VPfoR7j612LAAio9LkTzP5YLXCbgoOMB+n9czh8XhkYAYC/
6kHuPOHTJsVFz7PadD/nWVfNatwynLjrfUkKjwpXk2CnuClHsaWO1Bk6776Vo+mm
brde4MkBMKq+okdB/VL2GQbyja8a1JETdeedn4T9Xg3b2/E2cErl5urm9C0QSjFm
8MAS53xaV8dXY6mMER49Keb0q6MWxAjyUgHysEF7x9zNB7CPU2Yg56/SAnCdbDiG
IGsYq8j7XHC29TAhsUT7V1zuF2Cwewegpg+aowP8zaYd18tmP2fsZdGWFJtRCHS1
SSJpQrf/aBr3Y0CPTOeOyB68wbCat1WTifKY7xR9C9CNObARCKoLvSoZPZjrfU5k
qjlNxd1sASOzJCzoamzMfQcDFYvcnpwXIOSIxCppa8UQPaaHMNlrBHxn8cjMAh7I
rUPPk5KhKXMX6tzS7/eRXflQ1q+8OsW8bkJnZByPteJ47VoNq3odyO3wZYvSGgPX
/3ofhXupR9pTjz3GnOVpJAv7thaDlUeDoAb37kLqFpYXynXwI8o/qKdt5Y7LOmAP
mXxF5MFlogEdWxaH1CROAnCjOS7JSjj3fLkLodnRm7HojA/iIbA4D5RuNV74b+j2
rLLmk/WdeYKSe+WDFMk70Zgt4qm/VCmVQrZHrM/EGBl86NAyy4QarwA7BmTM8pQe
aOh9ceMvoxOMM/e2qCnzbbhsVsErKpEdWSIHGgUB1tu27IRl12ciIfD1ZMiihalU
jvJIaPUk54QX3a4MHwzZRiodKXVD+IG9NYZeGdNuXrMixIj7hXHdkIajCQVTmr+6
7bHmaLxXk9F71xpfGl0qiMhNhwBVVf0Qx0+18qwQ6R1gozgXGgk7RGPt4zVcjbnk
xDrZLo8Ie/1TX4HajxdDLqMP2kuoN0TXjpt1uJZI0WtmbwyhJyE6Ku6C9pQc62mL
vmkazrC/R5p4E3YmPxXE0I2XMDtVcZfwQ80nFLMzr830Y+BDz9fYPC+FL02cFTDW
iiSmXDVxoUdWtc+MA6gCMdAXkVjwbOU9iZlALjxRn873ZF1pz+i7XuijrRBB5/RV
vTrnBRbFqC+b/G9WlQFr8+6Pc9DwI5j8lEb75jWCYfrrWpLE0NMozh+If9Z7Pdpz
4imzZvcho0WbbDYcTP1by2e5ACsUD5d9zzRMsETt9b4ZAR18lXkSvsXOYKGd3sjF
ZZ1mnCdC621HG1USKCoqYtwmmObiUbDHpzORffpwc5nX6WMa7Ns2/OJLmpJp57gp
y70YSr4ib7Qtx06R2Hmyuwl7qgrZ+us/5dcu1CKOPGaM4CeSwBBFezftD7qbQ2DX
zmXvbaFvp7u3QaJrM/ljJ8J5xb8enLTOuPzYNaW+2tnDJqdmUNIBRbZO8PtnAk9Y
J/riydC4saH4/rgwEfQq6svYo4TGDOxE5K/RgxO9CxYq0QUOukpxqmA5Q3yA7Gau
S7Aizi5oFQ3EuS59VRAsegBnELOpWGTLGHUp/ivw+ylwwOSS1kGg3JWKqjP4LWMw
/5VuKsVDPBlK5YqjA+gaT80pyw8LOv2sWfqXcpNDcUQX7z46rg3AKpY0N6ut8LXv
nz6yknggEQxVVTRZmKsAWWR7kXcuN0ikKNt7/CnKNwJhMtW1+ildpL9RAsAS4XBs
ejXm7zEx16W9X+IbO0hjufZegookvpO0KsiT9HPS71B2/QWSDHrpjML3zSu4alce
y8UG+EPAWmAy6tXg+tQanViBAfnqCCg+cHyo11HaYUymAOZfSmNjvN0zftP3kZcG
d3QwBzbQxm77lBOKLg/s/UtuY62VBa01tzdbiebxcHb86dcLpdNpIfPW73EsXCt9
pgj/2ipST10C667OhJpoH/4TZaB0sOMJtQx5UffxLTdGbNICwMlBfsKT3G9OzUs2
daHgRmuHvgPZQFp8xUBO2A5yyGoLjGnnMEB8XaO2gO3WmGOk3LGwQ8nj4bAaJwRl
vvsIb/NnCiN4qxLrPxUV3pOBrwILgWUO0zoCFbNcsLW7DErma6Mp+kzzS3D6Lwqs
M/n+K0a5rW1PEQQeJwOWB2dCovWFqTqH8uxf38/t9bMADanl9cMrMltToNnvbweg
GkCwIBlP7u8EyD2mhh+fJ9LqbzowzbwCKQL+3uKPDNx5fL0+WDUhaDLp3jaAhAVz
ApS6hpbJnm/SOPaDYkKcE/wCHzpUZ1N0hDDlUotx/WAD01P/feFVPDHsOxdcSggR
AZ4QYVdkdv5F7NUMtTjheiPJMGGO+xJfUpMt1Pyrja1r/LFarrNQ4z1DTDRXmQ7p
OBsL8xs0vZ149jnOc5QF7M+bwT6Rggi/iRcwpH507/ouiSnzaFcrSC/Vl/YGu4yq
s8OXPRPJ+l4KBbzPwEzh1aR8LlekTzFgHUho+6FwhMdbw8qDkXUb2IYTyUn994BK
FkHmkIwqMeks7DkqrXm6ZtKpzE4Vj3vImOsoZvNyPMVJsHVvk2C9fcom4D70rQ5X
dSX/7Dun/Xm7Ki0WVT8juFIUUL5fBQk7Pc5HQalA1yqRllg5rIAzq30R02xZptx4
nOVVq0lyeYRS3MxbddEwiiV9U+qcE2XkKj0iYmZT5LvyHjKRpHTpe/tpzziMSFjh
+5PobQonpEfsDYv3CE1rKOFH+3lyMg0qo8UFK+OEpf0lW4DjvjOlTrIUeABmQ+b+
bd7InAqJLngNOyH92DNBfDs72+NBxXf+WdAhF2o6U1gZ15zAZHtIjQZ1nCACn8Mi
VxHNUbTBeQ13kFAv2E1S7N9abIGfUc8i5OPsYzn82tFd9kNvLma6HvMqWpnaCtnP
k7AibrVCrYMrKhBATwvnSuqGXiIdy6IwWH7o4sZJqak+kDCczw5V3ur0Wo64w74n
ooRYQ4AY3wlIc9mqWW7HbiWLpVoj2WDLBUL4aDhFBedUdLG9vCfRY85GqM9/FZB8
+feqOXpFNLGIcJi4VFM2dBkbm3VQ4uvbx+XXDlGMkUgQzZyRK0LAeP3xTYyiA3oI
i6WNVBUtZjYN6T5fhcP2xTbVaAHNhNB5Wc00/OzHthFn/re7AKQoQCWrLnadMLmh
qWV8lxJwxSy9uwkirZIa+Y7JjkZONRg7UrfJaXD7VnJ+pNfQRCorctTwxvot1NIT
Q5/4Z9nUCopAm2072GqyOsEXBYtlia/22kzwlyYrkXEY0bnBozri/ji6/wrcm/AQ
BqboYhr0VAd53WtGB3TNgE4sSb30vRg6IKU/DHAktnuzvrDpQm6JRHlqpLGhaXC9
sHUuUgNk7mYZc9qlQBr14/bhBo6nmq3ihZsKly80bOmGALUWfVQ/vBIFx35g2V+6
poaU0SjBZbaRxmPNCAlQbmrd4JB9i9VJZHjIxriP1XjRbXYAJ5t/UzDSM1bbyvbX
0nGhH7zQ0OaDzsfeOCwwnEmoXMbl78aqB0l65bKIRKbXH/V2raQcF1dQkC3QIkOg
dhlpeCF3f9dm8pG9M9dEEvL3zW4xmrgn8nTcminbi1SohJTCg0Q6aHgyUyA9sUs9
6QYZ/AxB6qSiudVQEKqdR8EJHofYb1oZW8Nl/uaCSYxouVyHSq5KEzx6/Pwq1xEp
UUFDZv/aJaoQjGio1YgfJA/w0Ievx4cXuluPkKQzXzN17//BopKNwm5B07YgIi+W
t9W7NvK5MRH1FuE4FOATi2J3H/E940ZYY0fLbq7xgPyluvDd3zemkhCSX+nUZeuv
1Bh7p7GgkV/SE8gRVpB6XXEKW+V2XGmYFh2V0lbKN1NgwiJBWIe1L2SW0OVUvqGr
RdlXLw+iquGS/DhClmaMgOJ5maajiwcw/N+UJv2i7HL4MLJodRQLjMOT/BbktnZF
ikK80DIh4FJt8WWoiGYifa8NLILfaY0zeKoSYFlqGQ/8e35aUK0hp2b6URyyQcoS
XGXJt7J4ldSWI6pYmDQ3V6lPcX1vHwoiC40KO9kkGHUvXW6cMWnJy8gWaTAUba0u
2FtWyAA7N3ss6yhuLnubua+BTRIoczVTEsMQpIiTeKr/AdF4O86X/PwJci+TVMqR
ksgicxBU4LqUpkqzLz71IqNqab8r3SN7mRi+PNyPjHbWxEzjDjhquwPDkMT8F5bk
fOZr1mfkt15Udcee9BssVkmKa39Ar1J1arvGDmvLn2azTbgrJmS4uzw/jBV8FsOz
nAaEEnZjPAdDbKZ6Yf7lGghJxhk7PDRngAUJqtM3fe6zP95eFkuZ3fVWDvArH+re
8SlKzz3fJoO5HjWtVdWpiPv3EBfHmhAOYUXRN2IyCdWNaIZuNDgC4NepLbmwdITp
GqQkr9tHq3mCpOmV3FV4+4XKxbIhIghNFPYv8jCBceu6/rXLNEXITWHPeTMdfoYq
iB/7DLOttY59ykhwLcXW09pNXJpfERqhll/7XiJuyf7VQyUd9pTrvBcFkI2REdMn
WBUc6NdeGlEwQtmkL+uIdqJaOk92eK/+o/FhEBG0S1r8JyWVhyvCpXlDN7e/cAaV
BvVeYO9fhvrUBArw6AVdIR0wGgJSNW7EjWHKSrGiXMKjihNIJRshh0O7yp4mYqUo
E9rHCa5r05P+eQh0fuWVUAw+/W4kwOVOtGBqjGcqThxy7B4+z7RxETug+tUk7pWX
8/wT8zd/VIqFlUzbce6sSED2U93RMrCqnjjLcA51aqy95W2BSyhgaNbiZwyf155Z
yHx6smeJHoUNgBDnGXqM6fBkwBJuiV6aAUKzoEPy+DeZvghrHt8i+NIR/3EP7mgK
QSlzyaSpKRRFnpSffpjQoQPzxgfpPSURNfC056B8Wc5hg4bZHWHgp7Cv8b+jie9S
kFnQFby3KUzL24HKhuAO+zW9EIaBjdZwgV8QFV4zXzhxMvVYV7Jjv3EpQcBBrzAu
JCIDMwEuBan/2HeVo4m+GhNS5/Lrf1mhghx/2oARu572uTudwL/9SYQ+2BLz7EIQ
MVMWlqpsC3x/8mHJTQf12StDYBrRM+DMF9iKzcd6ZlKPTFA+UV6trp5HwMEw+Z2F
Y7FKhADEpqSJ9J9WVeoxVXxnzsL0uK6nQUhN52sry8K6SthzKjprqka8ReePnkd9
wrVPV8+qFj4SG4vhbwnUQYyVVHXUu2lNkfryp2L2NcO9qzceKJ/hzgG0GPr6wt/0
ppB+8O7bvDcGaqaIgxGTTtCq9bUgEyOwUkfMJwPA6TXzd+etRiW2vHt2rhw9gVbp
K6LEY5INnGRQEkFI23KLzlZIhcuRaAO6hwr31LMD6rUoJTZw/Y0JILMEsdyIb/AA
Hd22WLEUSn0B3CY6/hi8azwfkw8I9VFfSlq7Lu83QKGj8H77ZnAA24DhBvxfMyXd
FPS6hEi/LWfK3PJpt8nixVj9O+lrgsuxRWanBF45lAi6rcaVLhCO7VItd137uYbR
9tYWUKXteN4i5WqTYPwhjxY963LJhX9Az3UCV6dVp/JDKO+GsWXvKU7foC/va64a
WKxMKioA9s+PLtKCVc8boxO+ntoBurzdyUDoV7VSdg0w52LuiLE7M6GfdjKMcgOW
bdWIruLBmvKhquOvBepdkTjttZI15HkkNXazCzDdschKtIXz5fF7Kn+8qLHFcjzX
9VgU3KBa4017kTt5zdBV4UGmAjoMluYFc4iLZM2iFmyTxwGyTaRpNLtpkgmtF9id
5XdQZZBXignb1as6bAWO6giehBNreZ6dlp561rtVCgG2cYsDx/GlDTFE1oPn3SCU
TQyPohxfBod/6uZvpSFOJ/7zYhGsOH2GT4CnZ1PQVHao94EVb2sYKFs8rv5ngl6h
R1nPbAFhxg4zN/5QVAAxlYXOinFS02tVmKCIxhDDED5taINpDp1+uu3DzcShQZq3
1S7Ukbcy0J2d6MYz1QLQoiloihJDjLAC+6R4nNBtvupYrW0iEm93YVd5l69zzFZx
a3OmPkA95XWN+7FXny53I5Elxui233FOCEF6JVq/S9+uoBUh4bTTg06ft6fJ5u7r
DTXeCJ3wxw47bDUVfTd90sVSjttjFLosqJqPDC3J6KaXDpqEuaDTo0EKDMoH7PdL
yz9fn5rPzk+b/PNgqnYRYOw08rCsJZyqMExn4AdxH+HJjGXFSlfkHUsO+Lj/NVYe
EGxWzlwPY3VJum6Me3UgybLG6k8TMqTbncoUG+g2Maa70GK2PRFsf8lH0pXr9T+X
2CLvV6JffK9elKE/tb8N6yQ9LiKBRgAkaNEVNSltOjgAroi1Q865yCklHNavB0J3
t7ZBHyabTOnDukLv2rUOmta7owtT/reM6CM1Mi6QzvJ7JVYxP8e3tKEakcRHbqc3
aWAcJjPjPYtmFviFYk1NuiO4mXKF8OsHp7AePU6eSqI4CxD7+TPTg+NZlc8Cgl8k
Ubhc18cceG7IBsnGkPFmA7Jykzjk5/UVnd7oa+RTljcNSyZaLgFUC6f0X7bYF5UH
T6Gxgger4aINib9jmt9q9UIGBHyTapkSmvY45Lsgwn5U02TuZhIm6M8fXis0KTho
q+oP0bdjhzVSrDnCG93Z3DqJX09HJGH47rzn+18ILowxpEUcntEKkGh0nIkIFyni
akjEHnn8lYuZVHhVF/R3AanCGOZk1yoyBZ87k6hK1QAqVf+HgdHSBGbjHafkCrLD
t463a+i6sRY34W8yw27T5uDSUshd4IvoU8Hx85Wv3+/nJN85RJb30KhKXhYRbC4d
wDWzJMx38kK30cu9Dn75wILmiUN7l+uYiFgLYarVJlz7imNfr3y2cE4Q/Hn0eysW
SXiDOrlBtRjfBYO3yPSIr/svq4896w/qHQHSpGeLImQ8ONORZLKhzliLCbNnlRRi
Rup9JSMDg3/JafxrBCMWLyZcM7h4Y+1PptQZ7YKrXZrqvoHPdYXl5qQasWhcSP/P
MOl6Fa6fd3E4MUy3IJuVhaPXaXbAjTzFgDu8LjkG9fsh50QX8jfjJq3OgoYhsKGZ
V1tGnkf5yzqOEK2LpKWuV/0rLIuKN5aHQdP8pYPdhyyvhqlEgdr2O1aeQ4adD0fX
ef303z7IYX3a6vX0Tr+MH5x1dTLjkC/UmiB9TK+UqEoG85YUYHEU4oo6WLdPOKr+
PAsF1g9t88dY0x1/3CHvVOScVqlA3JEX6esr/o7Ua7P+9kJHNbl+r9xbTOE2ZKBd
ma0yZwAdTAjBIZgB0b8NjIPMM/rtmbeyqiLDm1ovJyqYMS3p1wayfrXekjKToF+j
QZmqzuszaG+o8jhMcuudmsAiAQFw4/s6fk8GbeTFfN5WPSr3k/PCfDQywChR+B1e
MZ1eYuPezZVGQH1LwtEYghbq/iGmgqG9FmfvMO0/MHccaU8kydhFkTT9bQRy0AEA
eeuX3o0TV0HMU1JWUlxRVXbHyGNowOJ1M/M2aLBRceK2nn7OZtiwpkWHCoNaozZZ
oUdSDZTddPOlMYTd8TrEvrkMmssY4SmCnLIkki7ZFKILj3Y2XCqns8Ix9gb7r4Xy
2kX3+D4SjhgNTI8D6PXV5bN13G/pFl+3a/su/ycgqOf5wX7XmftM/mjvr2H35IWl
3ovl1u62ob/O/gbS735wt/952l7eS3dsd8C/dsJVMqY3Ufe/zHYvZ78tvHNnCDiZ
h6el2mcXpT4T/O3vM2H17iuv9SPF/swc/4MkrhZT7eFUfYyj3CBwzbeTgx1lRYDo
W8K8fmoIwdcGUvaVuLwv+428Vv//LxwLKSQiNSPvZXzvAtnwKHHDRXrpVxacQucL
ztatrSBqmV++8sA09ImC+Ysu9Z8A5OjlpPo51IJEdGjTzusPoYvdTMhSXmOC4/19
atnJimJ6I2SWMj2bSbueW7E7b6DnBcB1cy5OzuV0WLiq4ylaH5DGZW1yIp6hrTCI
9nqxRMPnMTZQxcPB5FJ4dIKsmRphnnjJZ8RCwxHyrkOmko9RKAKpkJ67bzkv+eb7
gO+yUDEgFEU/d4Q4oq+PwScNp0/Qux6o9/9aT3JocyCCwmLWTw3XW5WRbW97pq/v
BOZ2bLTAzE/MWPrEC8OudBnn49ZogClRKhuLhdtdrAytySynNMwkssW2ILX2q6na
tKnSQCQLuA9HCvO8ki9v+TATLQDSkvxSX0Qxlpe4B2HNLYN2tYZaSAcGSrFUVHCs
bov/fdHmbzy5JDLKOYHEM23pyJpvIeQgTW7OpjBn84dDAw2F0thROXIHB7EqpkGK
qYQ80zPzGaGM+mInMBUKe06WpvD2G5vZBd3ZRWSjJ1y7uUQVSsubAgZ2KHFYgE1m
ghbpmZHu7syCHPgYy7nRQnIKCVGFOD43mxafCOaym4Xc/9cqRvUwmClQ2dkbwkVt
ye8MAtNzb3uN4PUQQq9TKTyaVGKpow3L5snVsb9Ow8x4E2cz4p1hqR5XXz8Cgyh3
BWkeQ7GDL6ziv5TY4qUXc7Ji2fI1cA16nfhv20Wktw64ZrHIT+EJTktBQns1iizX
zjJEnkuu5Q98kjf7YFck/R74g2N0I2u8IEBd3Zu0MCWMsqm8ck062Auj6fqLbIZJ
4gYfK37kKiFMhqzGXv6wLrp9AGvC93zuuwy3mrPDnTRxcEfOLrp2j7Km0vtaJImY
stuZZiVrGlX4qpRc2OJeyckdjF6/sHBnMVctDBGWjfx5Id+gXgJirpaK3jUkqewh
63cK3nXd3WqSuqb0UXiY8obgfj7ejEV2irvi/M6fu/OHDEjYURINvKVjEjA5C4+T
wX3D8++nn3Imv7AibqiRczQfalFMUJz7hekgATZrz27rAp448L6PwZb0z+5hBN4X
NqjAWRC7xcIo/dgjF/VHE+yF+zcEoggSBOm04kc41F2CNkvPRk0yfGTHTSDxZZOm
9wzjDWZpP+kQWP5EOW3lidtPPQimkbvQBhpkBmo307ka+vl9frtNS1Q/mLIxq627
C6nfaosmK8pkHDelB/byafPFhA4XBb7oGdCmaVBBfvQQjDL6fWCahWsXM5ynhZCX
BC96/g+1ORAzsWIMlfz8XPaOwJ39doDksQgX1yOEn8lfTdJS2mu/yqP9GpExKgQb
rPfaE4aizf6oWHj5H7YuoMRKRYb6o3Ecq1VOPhDzEpFn+n7DrdR3MpBEg6aHBhLX
3GUaQLJxSy51DauKdRzpJIgF22mghR08UQOOjMyLRzNUHvZuK3VNMNJeDf3MWQ1d
Irn1G+oc15lTdEGClE7I+57epknZKV492KKZ6Q1y9Ny+njUip0XS/xyb+bC4OtuG
fM9nztEFiIublKgdluWV+wD7jyFSVVKSZPX+GVJ/8gowdEfX91nixFyc7E30V0Ot
n9IYGKIqpnTFU0GproLOdepdX/fR0F7EPZrsAiDXBPlROCJb7LIuw0eDEeOXdGlp
Bdi/loMO/vXnBZuQ8F3fxkgDYOUDHZSAdPT9lw3yriQHGudWq577n7Htn0qxEZTc
8UfpIHqCyfV2J4NNSYGYTYJHQw4k+XVnYVBrSc5lw9vFtogTYyBU3NA+Zm2xibwx
z5kTwHPskz6lLFPRhKBA1qq3K7VHUewuZN5yj7X0lD0jnlMUBpWK1lwcM+lVhH7f
2+eoyvC4WbNEgMqdMPxaK/cRwFlOUUGSKbSgb0TWk9480WByIwVgoF1MsgIkSecW
8BaFOasrJN/jN47BvtazE44lJq8GNPKtAfjuJESD+Ngh9tHh3rxCUlJEhpfgJCah
gqZAznyOkLF8XewBMAGkW5DBPHJ3dmJsMjzWnbJ2fv4T+B4Vky/fOsD25G4rz5Zb
OLwdOVHvEONWGprTFZL4o5PiZNY2uEayFGQ6VkUOKTpyvqvRbuDDnfvVOdx3TnYb
dwkRhFzQq8EiZapu1WjJ1o3wYVe72kqDZsLyNEodcTPFEwpqrLMo+KdMiVAmhDji
8Mf5Fd+st1ZVpuRbGcdQLU3G5PGOTQvlRdZa9/IRlUZyqPd66Z4YQnE1/13NwAbn
U7QZtztfbeFy4TXgKk7yd/0lGv7MjMN3uC3R19aE4/UHu2nfB+6pH5L90ZRBQirB
GwUyEiGE/pdZKwyXwKUwlKwWH9HQZYrN0rwehMwpIwACuvpc+KTthZ2xZz2rRWIo
zl++mrgbn3tmiCgPucB6AdLV2fSbyhglpnkR6vmgpZq0zXi0XANilPllz0TK77PK
79ZkDRgZNbi0sOmR9slN9koHUEX5wkcqG+PnCG/iOkFFud2XC1ZtO56nsRJguzW0
6Nzm5YTIFQ2qafAnVwLdcybTpkiCIW8AUHS0OK6g51+/uMI+iQJSnS04PUP82qI+
mArQJuGod7n7nfhXlDdgAf7hy6hEmhfGu61eX/tpr4jIZXaYEpCCPEsTzAbOr6lI
ZHKW+4vHjyiSPyLsUQhWZkX4qwp38oAV0sdpjdxgK5f1k1fGZefqdW3gK4jQZhO2
LgNM5ZvoKiURypFim4fhIQtmkX5+hfwxaRZ32xXV5Oaon6ICQY/ZVkh760OpMt0N
mh+5uTF1iVlC1hGQtTAKusVD3/o8+vppMFMYjGAQCDY65Kjb2nuDv4vAb9dwaHFy
Bw+aqwPKeCHyO2aT/PnLsZF4SHQldOX9nZ+ecquGhcVhHv4+0fm03vkV9edQIBOZ
EFkwW00zQoah1KJxhO4QAeVKN62nxA+FFqfOtyXLxykbwidCSJ/joXurTMhQpFOs
F9AywVXpa6xmU+huaWoINt+R5bNt0c6MvmQg593b7pyIpQyEXKI/w+34IA8dkXLK
bw9+U9f6dma3Kb31rhmANkSxwb7kemLphXylGB/bZBkKOoIKUoRsZy8lvq0S9MPU
LD4qiZpVrfFEvfitm3XtPuhzq+3Hzq85uJYFqTfogFELNUC8vCh6Go1aZjKqWXYh
PfjS7fn5VIEbiWYlsU/CY/o5H6jFTJ5FF/yOFwPz5LYgs83Feq3g1MDTkK5Bh9GH
sYj9Nik9kb6arSZ7JsymExRMbkinJ9UX14Dj7bXbJ5q4KAzI2NqW7QEKNBz+7lXK
eFX9oPITF9RkOSU7mfZ4xM3kDJmaXP6Qdx6tBNh0ABWK0vC/CpvdqSb1jy/WhIpo
2wvwzPiwpm7rFWqTuoyrGG/PNspUDO3ardxUX81aGTuk+GgtqqGvZWCsTkLD0jMS
awXnxYrph8zd1o1CCTiskQK6Tb4N3sQjUWvxwBehWqrEoxzS1RuKi0KR1oJFBCOI
Y6bsR6tSMdmU7sZERShw4hpuQxp3sJzepHZ3juTE+IBi2rXp9fLyHWKNu7sk03WH
gAI5pb1a6wB+BttbeUcTJ/n7ER+aW4cs11m+/OulOW1cMzLDQYSxLI6DGNOzXgAI
FLuDsuvyPl5zXmn35fvTtqowYOoi3a5rdEFP8t6KHynXLfPYgVs44ykcBRugz37k
wcVT2lZBmGJtZd5vXUSkCwblYB3abDwe4xh8AeBjTJbJbMa58uftLvdUXpSZMPgj
IhlRN0dB2s5RriH3YMIiWzvnb0Hbzjeni+RNlPyj/rrhIv1epbHa/kAmHmX49TeG
E93FnXVT9iKXf7qs/+CgzIh2jw/UUIVtPBokmb7/WTK98KzWqfsv9cD1sKh6YWR7
FqlmOJL5EwRBHrr9dCbul9PzPVjB/nyZ3VZxwMkCF6hV62vS/AuGS7YQNrldKJiU
2C9yA4Z+LmhR7ZG16/lroPlcU6hSdWVgMnuP96RfUw+kW9T/R0+HseTr593jXD2G
gvahTm+yboU+J1sFOPdi6JsMuqiMfe3zhQh3g2xuigdxjcv+SQPuJ/ortveB72O5
5lpNJ2GvHF+9PDJg6AsHp9WDhY1Tzj0ZuMS7tZpxC+XGxf/Lv4ean/c8i99ZRS/S
iQD4pWJog3pgBO0mPY3XI/C15uHbZnFMzkR0nxlY2zRuVDBgGh2BZo8Ai2M2wQad
UEl1AnuDFrOvQ0joziOpxdOmTMB1jEZRbjOXD9EdqrnuDMTKmK1odfB+HYvFsTpT
UnTUaDzVk5qk/TP9Fij4CFfSPLj6T6bWdU3qd8VYhoX10MYFsOGE2eIZ3XUftmHC
pdp1DZx4CZZW6o6fRs7lRyqbG2FCi/wnl2L2nUOfTqUaPeyMG5dzPF9pS7KNd/Kj
M+bj0fx61B/x5XwHSoXnla3fw3CK4a7k0UnRvSaD+lL1xRihJ8kMBOKopBns6Tbu
vh37wHGC4JKHugXkzVAbj/gL7BDDvh9tGbuqxvDKDfq4fFtOI361BhRbw5i1bOPU
bepMDvLPMAxFo0p8E9/Ey2fG5EQAxw7MhpcVaLhOizA3ZWsGILVLI6WZgOmp6K4k
qIrd3LmvQ9PannJU/MZJPUKgE46VIjHQ3z9678RK+EZ6vItBgbBL0gHAh205kObd
thjmwt4LylNzbx3zg+97VabK5dnc3j6ZniSMubG9+/aEtqL5NZBZrtbZ8cfCHK3n
cFMvuBmx2eIRZ7U4cQkIdp/24MiB7jP40ZQ2efBAN6KYTc38ZsM2iqAgbKUP1eP8
obRqKZGqhVNlcArm0aq8NhLZLJT1VTEbwwkvlZnZ5DZviq3SfwtwgqdRWxcWlL6h
FjWfGMVFxDeChphRNQQF6IsTThsynZFPE/um1m1B7E2x+v03LcIbwDcICFWkUlif
Aem2ONB9DHvDgUdCYYjxxUrJaf9ilf0mh0cuarUjtFUhYMDJf6+LYBoCBy9nklZp
dDMNdTNdx2jHMryvaPaKIDZNTYGyK48h8J97/QuVDjeKKFWunrZOjTGdIm+7I1GJ
a388Z+nVnCDPpKC3aL1bKt2fUCbXyjhSvcsj4FxeFBetGimEgQJ/K/uYSq8nOJ/c
bV1JruUdsczR2zW7T/w3ZksbR0TZ10ZHK1xWZrZ/WfSXL/9fensSAMbyt4fiWKLf
znAZWFISaktDTHHOzyeyDNUg79lXODNV4y5hhe39Jjts45w85b0hE7N3H4UMwRpW
lFwKiuNNJE6nGyI4gZdM0pdS7iQB+9Z8DHyd66/Oq2RpYibeN0H6taLjc5JVGYgM
/aHQsqfCh+09DhPmipwKpqOHO1YSmkWuL8jGOWK6UO655gmT+lfYYfQRSjify3rS
+hACpgFeg1C9nJJaBqWLvfCFKdkL2tT/V9s/YZQwSsrU6wSH3b4hJ0WWAFjkgz9A
M9SBgWZCUYQ+YWpeK/KJcTWeFd2CVQE/5ZATfdCcUXYHFzp9t/U5Hx7n4UVOiz2w
xd3OwYsGe5xUhcc92sbtZ8QseYIQs8Kf5IOOzvzyM80KFlOe9GFJo0et0HZYPSx5
Thhfre4pvj0xS3n1j3gbm2e9Dx0SIPakYlJWAUYQG8jtz4LwerL6rtHiGbIu8Otf
3rihPJZGxaGuv8flA6hkg8L6k4hZ47ityXu9f7R6nZIItplZ2ozTZznUYd1PLqBm
Iy6rRYMRM2iLaTMDmqAxCoCpf6tdVh8F29jAST7CCHeKyx3HF5twQZn6fVpDa0s8
IZhpw6jbFIMCijliirNDOlOyTmdpNmAOSpA18+nZTo6BP7gSGvRUuQulpZK6u4u8
8fKKIC7qbLAl76QoQmngCzbnySg8jTk8DARecgBDckjxB+/ZbvU/kyTGNOYWdbDD
/SNok+5yE6YTLKs5/GivNlZ1QveQ6rA91iVBeSzVlNId60MlIUSm2+iEpKzLv/py
5umnw0wYF6M5fCcekjfdag7o7T7eQgk8aGvBv28PmbuuLhfTIBFNjMY4tVw8zjK4
J6phzouFY2NplGvRhSILJKB0jAufcol4kLCJDpHOrNCNx+EYpqLK5CdVMdt0ZCJd
+apIB5nwbHhDP07JhtQJCX5WWrWOGPs6SAnD+ROxTRISPXIxbSvBQ6jiNZI9D0qv
OlOgV5PhEOdx2yKafui+9bt8sfsuAjUKL1oSG/r/5BtrOEowPAs+mJtp8YF0Gqer
/09Q+OHlPZ07/E3Rg8vea6wsRVhmorEQVsUApMsIM6EFkVehj7M56dw6+MdB4b7D
HKTLu87nuRDyDqsQTc8I0opTZ1TUBYnVeOxN3uwtfsZg1vm67cy4O8VcczQLSgtq
83MpCWi5HE2YChvQvY3UEa7M7YAnAUkcBknzb3PywMxfxuNP/SbMkUpINYA/vIAd
TCNumRW2tB8j9OpJgJiBv3Op2Fq0qe9hRixzS7yOInBrUIqY1ysrpPowPBB4muwm
rhUlE/erfwXH2SsD9kMSJV59d1uXfpOyGC4X20tnp3y7muOIb+h0bWLuIiE9Sldf
n+7ltRmY8/syatIFPFx0mlqdOxlR0K4/KgJPWzKLaaMG+q5PI5zH63MFmglBXKFz
MPYeIeRxjUni0QBuVGSr1eokx+E+TbRvWAM9lLPnbWpYrCcjZAuEjrE4crM9u05R
9iKsfBqUQkh9j8bzau3Z62Gdq+qmfEskbHpYVJlDkhrtmatQXGRoeG/g8QgrGc0f
Jiaa6aLkfYQiqUOfaX+NJLhiEE+Pmk09yCjeFUjqCSbVjrD4z89Qcr+UPlD2jDv+
FGDpsky5zpbVUPWqpLU/YnCp/aguAL3hhwbGjJ/+sw+x5wtPctRrf2kSi47/CIRg
X9M7vvnkdrFUh8/QF28PF1GZvikFKjvBdNc+/9UmdFK9uvXIz5HESYL2Irj2ZGgw
US3UsOBnnAhA22DxXN9M3MCSmh+xZOcdJJs3wsQg5ujTC5kY3DD78vleABmiJ0Z3
wmFYP7fCe6UzzECJhwwZcZ5KPt7ydKpZoawPWqBlYqF/7MI5sTamm6mKchrixw1t
0fsEse/4xQkhAi+DEsAvihI6i8Jjv8VgDui/TbaMTCtePf7OfQc9DooxocNEBF/h
/gpl7/PXXlYvFS9g/wPGogmGMrcc4dbOXBk9VeGxoD2qmchuskv8xeQbGFUjWfqB
AfQfsDgOWCeBKz5TuWyvXz/9aCn/8hzzjTtjSQ/b5WQm2rPf/vuVtyNIA6xO8gd0
JjGvStwrMMQhA7zskvo9j/v1jyBNiCr088W/oj+gXEAcl6bzvGMimVwuu++cJ/nS
hBgQdh4dJ34Xze+RtYZAMwo/eXBbrrztnJNpWB+2piXo04Fj7jAZHFQ233xV/YED
FiiLHmam+XWW0yogDuqgaHnZ4snIjHiEePiiZ52CsWDh2RYKvM1KGEon4jtYgAIG
wNIuIJLy6ig+/VFn4MxJu6ydSzOOGXbbU9UdpSG3WqWs1pR0IOCsxNDpf7GF0aUC
JdSSDy9lhMkfgKg+0prLGuhkIQ8cAKI6A0W/mM6jPFCzhSj1OBl4ZWrnJLULOZE2
Kd4vu8HdQjpIhPK3+icRU4+PRVF5FS4EjlHiAZpSnSGJnXe9yIfLtqDXiMR2I4RD
YDc+btVy5hJ2rN4uv2uNPR+9zx7pcMFRLeHenSS30xBt8bksp5J7YzhsffdAxFgj
aG33QCUEZrCXoY/fWvxmrSuaCAe+s+CrjfMM4mpifrA7ZzvjSl3ss1yigquCZ0pi
U+iCBb//ww54hKQ17jWdFINFOGr6esLaUK0/EbKSExRc0w7wwsz0O3oB+0tYoBRF
DRIwZWND8reSrZT9n4C2i/JJasXRLwFELTqmpQv5PMjQcKb4qoxg1hvk/IqZWvbT
hfzrQhK070IHI6UjWvmgNbFwmEI/sz9Q2tBUpVVw2SjZe0C+zzAROK/j8QGYMBUM
OuvLXIVpfXflyD1zlfgFvn8ZE7iSIJjYXLmYLQxmwljlCkxgsVv78Y61MDHP2kMd
9gUeYbGQYM/ZtsijHjZIhVYyTgxqu7xCRt2ZDSXncpDmqPm0jqz2oTlttL7jna8Y
DzYw46x61xnVPO+NL2CtVMaXlw57NFuFC6EegNjzPJi95Jol2jT0x8Dqj5N8t0F9
xAqGuxD9f1d+POGvIZKV3eYxvBy1zpl+vsfmxHXYfHJosYylZTqmsRmkMhn5U/8U
ZPuZkXJliJpOs+pGrTcjCB8eN3gC3XCPxCwnwCJcTTbIX8vzoTjMn0ama9Z/YwVY
nJzLfWd2CV6nC6Evf8M11nelFrL7416awnaUOY+qFJ3yAM5VKqyxEFGiosL4mImR
mTN8xWXGl3iM5xBM7uvuNi+aML9jYtAIbMjMujmKZNiUJY5AXhwK4L85aAZRbbXt
xGgIbSdrOnwmEOM4AFdfYPNXmYh4NcWMmwy4H25mHnnwAfAna2VKJFdBBRCMm6LA
WbGbEONVBg1EvPF547EaESS68Qwm/lEe1Z0H1RRJCEGWfnkUGk/FHGy8a/KAnMix
qbOE6e5IONxAxie5iw5sFkBvHZKCxdl1aj3mZqhAEonLKjtn+ufdRg2XdjZfn99o
gyc5qdD/VItiXTtWgUdP/rHfwPSbqyim8QIqd+ql7NaEPdAHQ8/dErTHnYkJqRZo
b4IWLXy46/ximu1teM37x0hoR5VNtMNemkdRkDyAGTMqeNAkVp3ElRHlhuYWnOSw
DHbIPAwb4I9wr7Gl5U/RX/+MNXXh+FD6+syMWxAKr0+U9c8nrSBuwPS/kXUkoQD1
KIdyO0McdD2gpbAt28FTUfgmLQYRz4jSitDLNpioqzR3H1FNa07pdaLcZ033oCok
iHfYYUqL8z4vKcyKLKS1qeV/ft8/4foBAW7OPmE+kbb7sFcVxYrQikaFn07uSTYG
aJLj1adWCtZvGOrHzas9aUas7ehFUTEvvNkSOELUXZXYwxp6lU2lYYxYwJknLdHd
e796GiC47i2aNKDFh/US16acyEeThv70XqxtizViJSGlLWw3Q/egUkE6vIdvz9Pz
8c34czDtpYCR9sTYYggqArz0q0KO2npxexF7rejK48qO+x4A72T6sOWBuGZcIxrU
7VGmSogmTbDtr1lqhqLixKSOwv0UfgPuZ9IxHAWMDb9ZuQjTqmje+gth47rV6gHg
cbyoRwMmqKNB7NFc3gewUoYagyQNP93MyTfWVdP2ICzDLKBi82taacSwJLYTtrE/
Ji58amHVloLCFwr34/aAVk8Y4cBM2Nm5kFnK1GULBJGqgA8uzZa6z+NmgAWa9QtZ
EQK9u5g5vb92Kkp/LstUnQrqyTNQiA3KebFmYW9lURJLIOPfMHpooiyUe1efwHCM
USMcYgzupjNJCO+FwL235/ou3n0XL0lv7pKz1mnkVlFk9FLJ8tFvApvvvSWf2x+8
ntStBnDqiB/FTsazAG+KaoPvV9Ylj/CmX+9wTr11enQEusKlnlGHEbAB+OSYvQyk
zWTQ2zp5MCTqvBI0eNup2siDyNlsai+pTyxBiIkXh27qrk902WUKO3HIbuqcqVSz
ueFma1q8oLn8BxEqeJwFN9Tf3QWJgxVr8JTHB7i4DYL+bUPoeqBBDgpXcErVmZnD
qFvNhf24RVGf7An5Wx5LMJ7ZDkpQT2/Y6V1GuNVVq3DRx89Uq1e41tqCqLlGZQbx
Z0x1dseOCLAXcVxej9EIFisKUR+SUR/XpRrLB1umJpgSZ5HKnbgX13w7TjllTu6U
kUVsl9AEMg9EJGefTRR3wvouxjaLroguc6YUDyxHZaRlgPKOHDdTikbGvX/saCFc
OqhYoxGf9loxLQ/8EnLSuJo8/nFZeq+/92gyeHmB0ibRWoNaw+sMeb5YPOYbU7rA
sGfxqAbWDQ5Aj+IEBHtPzIaFTxqnNoj1CPYtk/u7m36a2PF5ViL90hXGyU7Sf/j7
guJfh2wK9Jx75IB16hsPq1WE3SMMtn8FVNjOzxnXfcrp6JtHr1yAn0g+kVzXPxrZ
UIoa1xHPxNFhCUBWnJH+ABB04/OkRDFWf4Lgnp1d9sGBH3PeZkbQQ3E99RCA5qxD
73ap7nf6NGsM4HLuNUW1B6t3GRvHclQOsdD2j+hG4EY5+Vk9/C1k5XrRIjVECZVE
84EpFp8wO/4UbmH7eD583PzTf1dmg4q5dnhUZapmCc4t9ESKinuDu4eVCiRLO6sX
lG8hWTLT3mSl8WSsJLkEAARpslWbVyix7I3f8iVx4uYQNj3BsHXlPeeQiFtlIyNu
pvFo9kgAba6XYZEON2qVqHO8Y51IKkewnuAbjlYHF+m7IWG3brG98E4O4w8Zy+hR
6Ncw6JfSA5ef0u/7hsay3n6/SNFSJKOP3WdcmTXaPJubBpeuI/HUHmbd6CJAfZy6
Wwp8FegN259u0E+iD5fv53lPlkFTekVFhWmOIlde+77r6Cypokb5/BpP1pvU18Gv
Q9SAtySDBDfD4fD2HWLUg5qEcfnRQd2YEoMl3RbNyGhdK95kmr3Zeaslh4nnA771
1mYr9aqfu46HF0+gKY9qaeZ/3wwbIjjLg+vdPgXPMIyKs1Vt8KE1mYzNjUCxqjBY
Z6z12fEYC9q/RKc6YzCT1SvJVr4OiBwdwCW4PwCTi04GaLVPMJ7vkLqulLjrE8A6
5PR1PlTyRrZ/ham875xGdtVYMvEqTjTOXyIQWk7Fa9+TgLvNF0Tzoc5U0Mhxynq1
eIdFYLJdogan2rn1/Y4hp4WZON6ItCM/Gpg7w5RBoJL23oXjrhoPw7hKQWAHF6F1
XvZP93Tm3PWcf0MyjteU5Q65kHuQHzDIjP7s3Y9giiCU8H0pAosz0Jq5H153DOSn
vBKXAf0D8oqn9TC+xPsFbzT9LJJF5DgB02BV8lbXLjud3S8q5pBPtbLx2aTBvUBw
gcMA7ozP9fHkd1VvO0jbR9Nq4DrsTIyDDRzp0nZbI4raJ+3CzpGklAYlhiTJU4Yh
ALyzvisjJ68jxQyOAHIY0Hv52CMYNoXofgp6mv9SbsyoyHhn3zyRSdL7OcFfU5pn
uJiC1xA/sygRPsr59GlhhKObERdwoHXbqu25kCmnUH+ay2BHubumKGHdzEHdwY2o
Di6wkqBYzsI48B+K9ZJxPjPBR6V1P1pBU3QxK/u3MxHPuOz0zbuIDVRD/sZXed0D
pK5npqxBedk9xgW/rDFfzkkRM5tYKFCRggvRqOL5/bSfwaUpSTtlDR3ljVjD3YKW
VfWdnWcykg4eG38+bx+qPfec5h/fI4lLu1VF5UQs+xUCL0JNnxxhNwC3tVOpsHaW
2ysByvoZZha8oIhXsE6WaxzLNSH/2wx+8rgqPQ+SeDVXVVi13ICLfx+a4seZqszk
GprQezk5F1+pHsgKBPYAbeRYfF2FgMae0g8K/IZeTTygOh0wEkb3C6n1BCBbUtzv
C6oIWgZ5Nuc6zFrhIguhSIJzZSJp+yUdy/hFSgcaA8SrR1I1lrklqoivbpUG5Sy9
YbOnoSqsukx05zT5VRjEZ7qBwCdJKXg5AunRdQdfSndAvC4A/sAJ9APXr/J1j7GK
qtOfDRuEBNkDtgj4pdb+LfFoYPFV7hGusvFeQEtFnrFwhB9XHlpQvxnIHWjsK1jR
sqS8bCq1vcjrFsWe8Hx+nOK/8+xsPm1WzSMF4PViDPxAUKYx/UavlIK2wlB09Gae
LU5FBzTyXUpfRdE06ZKAMjIaaZ8+3X9EDTs/7lDkR6S31br9nPT+Hs6sMU7cXuRa
+dR2Y38QpOVxUkfPBKHNtGo1s/IHkY/Iy7nuuSuLD3P8Gub8avOE4eVVkZ9j9s9q
WhwNWsO4F+c2tZ+QkhdKz+Z3bjsKcOFVEGbSglusGz00i8/WRvKihPBFUTKuU08P
I1enV73Elez0tUOIFyfMxNG805DFNYwxgW25wKuydj0gJpm+6VO2iQeKD6joSzdT
dOZpl3kzQx1XHBj6evjfPia7M5ZZl625vdi51Y3eAGuKmfM3GUEp7X9BrbiplWxI
8jMb6HQwdVge6RBF0kOn4KnLP6ipc8pk4mLexOKq9D8SULlwjhVzI69/F/0Su78j
SHCHeLFTse782nizoNn61r+oZ8xLJFFCNDv8K4Gk+ftiYi1v/9V0Ar20E81nq1q1
FLh30PU3oXMIGKF7+RMfzGkDHQ91qYJSxWXag51PO3ps5ooTct5maBd+rpKLlSZd
UHwsw2a6mcgSC4BgDafaoNuit7ykEodQy0vk/+FFs6TpQo1+fYrgDFI7pCPdd70R
IXcxATiIbjMK6jtg5a6CxUDy3WNAddRGXOtl/eldVXQMc3JCZsDS48ESOdXYn23N
/DYEqrzxVYDamfEBI2oZgWYvK+g9wzNEi/qv3PF2nz+h5UZ2PIO/PCUodzDXm6lA
UIxlugeNL7tuLrVbpuxmEtldHHejRaeGFOb7JCMS7NWfiLqhz4K5RBdZ/j479Cic
iqab2RmpRbnX1JTr5q7z6SaGsqasc0v3ZhdJG4CGQog0r5rJkEKEUEwXNK97vmx8
D2u7F+YT4xLrqfX/emtOKtHyxlM9RLmPpLZchgom20JKOVtEuOfTi02r/irRf/c9
xU+rm7VRgD16bRUIx6KuXEYkxy9JAsziPQzAWJqDrqgOAEQ9QJEIIgN2Tf4lisB8
y9bnHrZa/TFC4t0vnENbFB0+8uAJ1RynuL9LuAge1ANUt1++wFe/7W+zDwToopM/
BKA2KwUHF5o9F6dAcfu+HUMJiPd/DtiLqXCfbYJQ+q+8Xo96D9M7NlAQevSmZe6/
x8VjXVBicYefpLkul22n1qs6kfTqhP30o7rzr1Bfx9yHyhdA2Uhug3W5iGZvVbnY
2p0JbOms9D1Ul7It+/RVmkjDhEJ/aGHDp8qGRaSbL7As8gMJCottiiOdo3vyjqRh
ZlCcdVDw8fykeQnQ3euewxnZMark0hY+rDj2PRjSJN+9wo2yWYTRT+7AIDkovSFP
iRt7rnjaxRhBJn/t1YIO/ih7Xm9kv+pI6Fz3mYoQ+3bZ6nffLvkSSXr6BkvHaixb
z4MK+365BIu5xMoobWoxgrLaYpk/wQKDaPCvCtRtnNjJHtod9Ciexi//8FJxfrwj
7LN88SBFbmOvlglGKWxazNh3CwLdZBRMaGNB2dUnv+sBNPb9hE17UMkxtZ1DpfEV
/+NRN2DiEhkrI/XM0lJbihQYKzZgAU72jsWo+t9bQbwDjaOg1tR+8mWpX/HDzoZg
n7tOu1yWfeg57jWYowWRKBzq4m6Jr/q2YLYJBM1qv9rfUskYP8mum4WXIlKs0h/e
kgRjFF3CLWXOlJ+qxjk6NCaMHWhxBiQYtZqEhLy1S+0fpL7fSW68oLi4UbQ6onA6
TWGhfEmd8WYiDzm0YQbGAM9o6PuQ1njRUju5PPF1zoorRhwY1xfW73qsn8TYAoxA
katX0uhi1k28T/UkIFgknCsYLfBOI7EC5K9jrMJ45gM7/kWzr7WUp36xj5RBrQQl
BORhSfZLbLZTCSswZP2QN9/pZoloLREFxXRPpU6gHe8qJEZSaDgpLIFIpGs6aBbH
lx3RWbKPxpwaHdWehbl//qTE0WWoyU34kofmnO8E0e8AwEZI8RQzdYkAxjkTwFi8
F9CM7FZMnT+KPBa1ZSWwmND9CZIH/zJV1WWHN9aO2gKFXYE67N0l/pSa6sVrJ6ip
mvIHiGM7WjLB4QsbDswxL0OskZkVaSHtOa46PnUdFxBtafWBe/a35mqyWTCwMCBJ
RcTDF2ElY65d6OmHHppvVzquL/jjX5yGKvEg281oyvcjyA1eQ+bS6rEeCXNYXd8k
B6p+wry+yL2vq+/tMdlMmFPZnnmtmB5vGRx82XtoSIG7IRDufNFP/4jvwQu3rZXu
K3TwDfOVw1ta+4ddg0/Bp7/DeuOt0IhqU0t83XuJp38gk2LUDX7lUNIUsDV6Is/8
9XcAn56bXl3zaijVxPn4ZEPP1xHgrwF+c746hiqSoY8SdbN3Y/lUQbejnrulffOq
GqUNzgXISzMQ4g9nHXEzs1Zy6+JansUWhdxVAcw9NVjGx+KUAJT49qLUtmRtk65y
+NAxw5epAXAsTfPvVQDp9x1qCeD1SLOZXI5/Ts7a50zo7VEUo/wP8k0KhnA69Fy/
ZspNhFsYwzvVjntpvWBLB/IGgUaS8X/BFgHniX8siRSz+050q3LSXYOXg2FAbMTq
0XJAgGNJfaTSP9Mn62HH8WqD3mRO5HDjd5ok+SiNYIi8l/V/VLsFlQvmQQX2nXet
3N+rVkj4ggYMuMA0XVtXGMtJVjhZjWdx29Cx82agb0D2pCwZfZq0VviYcTaGUjbX
VJsOxn2uR3TOOvk7bjg8bFrUh9DOSbUG7cUq9vQNDxFKHnBpC6EyZEUHeVJN0+gN
AA+ap7wfhua/D0oLFWZrLWa5LqsedciqRTfm6mWHgT/gSlglkZ20hp7tASSY8Ye2
A++Kd2VKjDeom7j4QC4+mABAsYpQiGnb3185shk0LbgSEy5XdRS6MdPZqtGCKM27
OCsxzmEwA45CufSETfoZC0r4PbMQfgbCt7onN708/Qo3GaKR7QSzKkgTO0jz8CCd
NSrsOI/odV/Dg88FsufkXBY5aqPm45GNUH2MYGom6SRRVzMZxN8G8pc2ST4mZrt4
BtBye3TlNhDdYjXSofWdo1SYTcrqIrAhCM/BseQojzaBUNgm82+ahrHxdolV1OmA
6gpUXO3Kc8SkmuNBTAW8G17+hOTqhiBlbzl2gLc2TLYjvlsZaErBCeizbCYh5jyX
XThFC+E+Wlpxi6d2jAn7jIzhtQezazCWt6QV5hhvlHxQqqGFHjXhs8tGOF6AUOTV
EWYEYm/oAFqGIP2E32mLTuK0MsKHH1gXjlLZG4SB6S0HzLvDj53SKCzP8ddpD+sm
4LbubkK4sB65U+Re/BiIEzN2RF6RO8SFz/qv+oc138gO9ghjQPlHnWSDG44HvWgL
G5j1A7c/9gqgXnzY7vIhww9aBU1ynKdy5i9x9/B/rGoZ6CsmwvL7jav2toJQQc9K
3FJyjuUCBMIDE1tpHAYPa/2tK8rQ9cdb0RpqQspwG5pww5shIm/5nMDwOGNKshoR
RB9yOjvRNnVlemBrg69lJaWRhtRIQ34+NCdraG/6z1D+uoDNOFumjtGFiwYnZBdt
zEtutNU/bHQJ1OkPLO5CyhNTAJWIVoMEX3zgKOCWnZuMSw17bATVcdVWLtFai1HP
VA+IGkmBSV2w01nWZ9QVRu1K0OqpQFdkWlBHQp8nz0olfd70x9cngVtt06p3/9dc
QqUm3UDdytr7ULtSQ8UeC5yhAY+jw7e/aKGYv2FkAAz5qbApoHIK3VP/faI86rzI
gAgj5FYZINB5dA1YVdWvWbxYiXHdCG3br5oA7p9SZ5tB5QN+Y5sR8xryfdPWLsQM
OvHqu/gHMYBVIS5cJke6A9xv8sO3RhZnI6M8T5B+Dqf9QVEBdgWoChSTTT/kREv/
j3I12uLMXctacQb6arzg4OK9XZoi9a3Z6pRw5PMqLmqyRIBpuyTTy0qHIEUI2yJs
Z0nid3XgjtTzCNm94lRVIzV7vDRTc10PK4DEqyDqrW3QJHtjtoyCcY3PYVwzttkl
67Dlc/YFX1lZmTSiv0GGp9vrlZiyWJMdKP6/8rN1J8RgVjiOUsk5pAwper8zY3K3
cyFnGnKjyIl2rkG/xPO099O6d04shHpsZUpgNKMSw+PtUz1x/zPdmV7kic1kK7O1
BV4swspw59pVELw5UXUARZe81ySIqUtYxMluxe1HnpL22y8wB67PETrmqa1eFYj5
BCUJO8LnCgzUOv7Y6sHraeiuGWJzA9hnSJJnqj4s6U+zAVHhfynuyCPjZCKSbQYc
2+kcwvSSRvBBijDMzBMUhR77wjK0u/A+0wMeOMtqO0g/K7Jh7QQzMphoh1nChr2w
74KaAYqf/4ChvFzXdgM+K53YUaEDqUwdKaI6OO8SIeUpnqCErC4mV1X3ozV2QGDd
i5PFlXRchNIlpswfss9E+3gEkcdD5r6SLqy/wNIdLiWCRhmFfMCXBtK10EvaXtlS
aYA0VvUhkU9ZJRjrQLTVmtGLA4oVC750hG7PcPJjDwRtNGId1zxbE287bL4TXfoW
S5p++/bsas+1cGzZN6umSAGZdvhf8V76wFbCX235uraxN69sI1WfDm27l6q7pkVo
HQr0EU1gvrMx/u8psNVxdFJmFVsoT4ANJXeuFk9bGTcjkvEwZJcJSBmPGVeD5g3I
hM55CRvMf4mtUC8YnLZChONgJrcy9BdydFYX7rqoN/IA1v8JStst4s54F70P6RNC
J7Ykwa7xN4v96BPgUCUGnTOHe8JK1pmD4YnV7KmPo7meOH6tbQ9YZyr7I3ti0UxS
Woqs1holUfZuviZaG/cE1uy3xU0Np3GKpebxh1IUAZvmXJMEpKoO/TyTfdoY1MOY
VuVpbxEkp9I6ZLV4BBOVrTxe9/OXPmGAqqf8UZadWv7cyQhxqFDHmywCMMYSjgIv
lA4ksp4x7sakPGZHFczlAkLuBNYRTNOlGpyV5Fxje14aejOhgZBKmz9zO+OoM4Th
y+NT3kzMB9G9lhhhE9BjAwO8rtfGeMnrlPFnD3XnDVaTn7vRVMvU4VkwoOp+DT5I
q+SMxjK670rXAT6SZQ0J8e2hz783pNG38hRVgOTcZA/MB+xEPDpfdd5EFDHHurLS
F2a51xRmKBrI36ZXFyCOg9VHr7QrJJ8mLi6V5SPuLbU6zayV1OnzV79rqJ5cnuN6
DILAgt6+w8/RmdjKkC4NtAMgAIt9JJGiFmn1z3j72DENU11rKopgsSFjRfRachVh
WDHHHr1Yhiq3hxU4lfO8RZuxLxMzP8nNd/fzSDqUIiScnj6X6uycDOOf+/Ib3uWw
mAgAZ5MW0dM3PkD32eygHm0jn4PinMKGE7ZD0X4f1bf3YzIazLaLI36saIaNKfd7
XuWchoN+O156bI05Y1oyxp/d+zew5kDrVZTA8KblK+oPCL235Io4YxZght/ztCma
/wGvM02j7qYuFEh4H3lw9OoGF7PA//vYZTu4RJUlqGKC6CPjjCs0dNHDCO4ubDHQ
6K1iZ/3kQtvLr6nLMm5kiHuDV5mEX021B0xO/PBzMzJpoiVfBA+FLKLB0T2jz8LS
hMGk+utzvqQxrYAEfIjHdD3a7bCyadkL7UjN0VT3agTtRVnEAgvFs84ryuC+YZG7
UTRXCzvJL708NEtziTPe5Za964iVfvRnu9bFad4up6W4W/WwjqOpZ9t5N7uwSsQ5
H5d/Oq25NNKtxGteDB9ATET0vIooOge22kHY1HWUZU/9oN5Pv5vAlLTyBUWU19Zg
voqcZQCKncXO91L07FkkBWsFPYVX+9jRs0pBsq9Rwld3sWZO73q4OXQBSmMI6HsS
rA8+Wv/2BIYOWZbBKXSXIVt4v2u355egcNnXygM2l/Hk93RzSj7FYWwvIHaQ1abH
EUFywvYB4Dxq9bzAtfOuwEzFAVdxlrCgmJ52kisEXWIzTkVMCch+AF3ErkylpApy
KPQJ1r8da6QiYoh13v5pu0DnGR36oHnDiWF0LtqDj+w0rwQnK+zQJcqQ0bPsrvQO
xKMfndIONF+ugOHHvoSwBODbqA7QyfoickSq4gSrVV/n4xA96Pi6nhB1uorWqhsP
m2QfOCkp76f6MAfu/yzdF/EPT10oNZDi5K4ybXrxDKQxLgNOVwd2uFzugEf1n4eK
BpwUh4qGhUFn0D0nIUnF4nCzqunYsQWI5nDlxgAXS68wMwlnodu9UDShS5nymWzG
m/UzqKl91H4CcVsvPQGo9Pz96rv3TpXw4PCIJb1ySbUX2wFuMKx0looT27P+JL3/
0bTEoDYLwf7/+ri+3fSBiDGif31lTR+OK61MnQsLAmAtF2seK+hR+9Iz6mBTyuEF
xnYP7iG5sIkShI7UW+VhTas4FtHriWZ/KvgvaiXBnSWg5z6Bw8yj031LtWYZVDiM
m8lb/CNrnZLD5FQOJpvUOy9PJ+jg3LUSxHUNNrIomRHsmczVqTcJ8eSfc8iiozWl
5NetyVRlGN6ybcpDwrNKEL7KPB6NlrvH9xDJgduMhNmqGewc6Lay9GTDF3wtadCB
1iTSCjaFhJJlo7nKFZ6dwbq8xgM667fm6wQTauuA7imCVnS7qRmkI+Of0cfY67Rf
PIrL5PS9lyo5og56pyPw2PeVxjyUH/WucuMWP1blP6NFf/zL+dLJrJk1dxP1qhvM
zz9U1NuvvaCRuMIG6QQLRy18VH2mVjb3zEt+GvdmoPxED64eoPympUl9uxXiRzwE
+Scp8zdso1IkU8xIPBzrUsgIX9521fMPpk+238KKLumJmYMssJa1IB8Mn8erCv+D
wkdPCprznmxVIqhYrI+WEvWhShhIb9QNlWQ5+ncVx8wlKZQgY/uAoPfFR88/6VL4
71iMYNjLGtHIUQZOgQkO+Q+mb4mQ3NZuZGRQ8/L64AfGv0dMaCjeZgJABu7pq08d
tIbbow+KGIih5cdHXIbrDZ1nP413OCXiFaUvZmyq4dzHCTWrjtVTieMvM+FzZ+/b
THevOxI6kaWWc7RUfnqnV/yxJMNMSwGf0WKSh1hHhDsjGECOGohTuJaZgz6H8bni
bYAL4sgZVhFNl4sJ9wkEEKcecF5WXbALh3fp9eMyU6f1gaeo6aYpGqZu/zax1MPF
70hnAFBp6z0ydx25udBzPYbrvnZHcLv9lBzwuDVc1npxpHhNlN45jLZ1Z7zvRG2E
9Lw9ZMFMlLiZvSkZQ93c4bd417LAv0k0Soae3EWQVqTaAbavJmMM2Nw4qt/i3P1V
0nyMa5Cc5BHUmDcl06P8Xup2Hc5GyHmSy2NdDiHG7d19mZ4bBhorlFGauj6G1jX6
qlvG5RL6xMXK+s756UNMhU6zHKsezCYrzgJMYxXrdfUnhZDQ4SL5SZjFuh53ks8m
4ygBkkv6euPShpU8nH69QWacunuFHIu+6pqRXAN5eIUdm4aJkzU0yVXSTImQjkXb
AU1MyRZ5CzKzxd48jmgM+cowAenkQg12jgN/bDC4DMyluiq4kFkPFpuRPWCmynqN
WTQpIfdg+DaYNrFbFRicEMRM5np96uZu3mfBbULdiyIo2LIcZYbReNSZpasIqKVQ
KDyWR2leAH7kCqZ1V7sXqN64axU/JcZRw6PtF9A/9Dh3aio1jPpmW6hQMF65/Zsa
cyF12X/WlKDULxJVi4N10t3Pak3GBMBVOsMI9oKRJu+i7HhTpsSkHDMfNDCgkKVz
ll6aypzXeBkdwvfBtmJRjyaGKlQoWtoZ7Us8YL/v7LOo+T6z09okQW00sBccBkb5
61VJZhuONBXEiETSttJS9gUEbxkGmjbD4kWDQjImBtcEeehZmQdBtxfs7lo9PbR0
hR2+2sbJaKMBWuL3g9S98aw10EM0CVaMU3SF6sRpOO/+RR2ugse0ETHcI8OR5ga1
k9LYK39ckvjgOHwwZSuQ89eHUm9aBJ8iWfgZCgIfpHpXoQm9KwjsU5sd1y+rMAPm
THUs+ilgj6X/TC00RQEhuzPItH6MiKqtWqIPiVpeyuu+UdkFT1PToD5kTbZIqKg1
f+Gbv2FhLeXtqQKqEV+zaZxSrl3V69r5WniXCGZ7khNRr3+4v8IqQUAComeiRoON
gd1yXH+jfMa8ScurAMH12sHKnytMAvl6cKbd+VPgDJd0H/kVuBIpSu1oMhzEAShA
5cfYEBqaGBxGr+Hge72G9rJVZ6f56eJ5jZPzPx9KIRcXB8oyETNTK14F+KsNKO9S
I9vW52nSFkqM6tASJs8rq62B39QE612MDbibqSprp/3cx/fpeb520ctmCggG1YJL
H+iXJKC8AvhCZpFLW+JNUkGHEMkIQz9idWJ2Od/qB24DCblKqOlW6WtwIhVGAXPc
F0PcqWgcKTVHD8/JcoqMOYzD3xSg8iZsYKfg+0lXeE0wwtgCPj1fbikYXBuSxRwG
ggcmRErrikXQzaXGrw5eDy4m0C73/0/K/AS01lkopNdZLSnfL5lDap8NlEjVXV33
W0owKoJV3EIjnlQ2KMcnE4wMvQ0TS2LjmqRfzKEkwYlj0sC+VaSnCW5S3nbzpWxf
t2/een8Ux0LPpCWoWThZp4QgPlk4UEUrYnfGTXlaSdx7UnLmimkGUVifj3jOYGth
Pht3wJA4K8XxmKVyGfYpissSNIqhu0qNXAvAKHelKcw0hH0vp6clxW+baNHZ2otd
fv/GJlo78bBkWZfJk4kWKq2myEJdge1L6Ty3fWXIRiGyo7vUZbHk7aJ2p3PrqmPH
VkKGYmK1ZJQpwK6+8zgLJIbeWlbXLhcGDxzwIGjgDNFs/jRtkaqqHxNB38syJt3H
e2Cx2f40OoIljJwse5eVDfIAWdKH4gQu8X6LsORW22spXYVNVVjIXwRGktDt991I
N0D4OEoEXkv2t9YSgbO1iYb1WhHyZnnYo4M5FW0aHJS5D2NYy1z/agnI/r/HIAvv
76wGXL20T0/5BoIkGRdZs6NyQKKfvPpbSxIEQ05OtSyy9KaVzNZUiAvV572parAu
n+MsH2Ut7pVM7wRxEAlp1o8zv5UvDQXIL3LV1iGah5Jl3j/318HhvBNbUsZWVfDG
y6joP4wc1UEiSLUYhg2fpg84OAMGdZ0/7pTPO+FMX4fWPxf5VrscEIG6TeZ8jzDi
icvgir51b5ckfCSIaGZTk16ZXgdurhMuow//uDEY3PSW2+syVmS5tuUzU8uNRrJ0
/ghl0HC8Ky2p9qcY7Ecf5kaQb8LGAbxYXNY2NGCxUm5UyHKSNK/E3pJMveGARn8X
CoPJnNrzMiL2OSdIRT212S13zHML+FgRPY+6drGe26CaYy13LMXbNNzM9NyT6HEn
aMc/h4vN2ZmyMSly7LW6kl281zwyWxNrQmiD3Ntmf2VD2xOIKG9gVIsQ3K804VQI
+VJchE5EEkvblfKnd8+13hw9RhxYEGGD59VyI2sMG+qmfXrHT8EEUbBmHOLaeYbf
bVlpTGAmF8Uz8EtLLqT22qmZObvU/DMP6m7u41FcB/YU5tVT8enZfWYr3vJlrZ9Q
aB2fJaCbfKd/RqThGlu+t25SqLsD94eDYDrOzQ7XHoR+3Y02m5iyh2X1XpEvHl2t
d8WOIFsqZt3t1uFNMNvZZBO/PYjVOCWX9NGLnu4Mvf8Em6P4ZhVUI2YESXTRRgSd
QddDghDcKpptUosamZ+EgQQkNGaqmVaZSe6PY9xGV6RO4lfHjEQhRiZGxD9irnRe
YxJYD6czXchoWzC+6ItOX/LL6NEqfNJ4MTMkNUpSl/sDl9UzOaO4NK+KTBDiPbeH
gdm1cC/7Gw1BagBM9bmMJiINUNrHfmVNJMg7e08TL+/korYieQ9KEqzbQC8NJbHu
Ux9ncM5okb3igNT3cdhGL8ZWciewe78e5+ubB4QklV55PgRuNEhAW0fMsAhftagt
ASOs8GOqBFW5HOFErC4hxPoDVGnsweay/DpSf7A0zTS7m0p1FTGxzlEE6psNGO1p
GuWvefhl8KPSrFF/onFbNNAUiuZnQXY1km6yP6ULFAPxBRFmA99/eAVWk6cPe/Sr
E11g52K4QpGxP5AahZ9CBugUTp4Txo/VtpkX3J/KfJVPq5rdxmoGQq/BHE8hFS06
ZTwHwDQGJH7YzXYpmLVwX3OYg6mqCIqRyYcGU8uI9xWW7S014iwNRFMkxXef1hBg
p65BthQtpLXl18P0I8/tZVbkF7IzoMwuTSTt92bSvd/a5WuJ2TdsX8Gq0o1XRtoG
6Bv3tiW743qnce+tBEwQhD/sTa6QPUv093olv9visGkKL/GXwVlwPsm6Tgc+TFrH
C6b1oq5GhiluEhyn/nzND+00qbDokJfSM6BlYC1arJk5NauBTgEeXtCjbYZANtxr
R1RRKu/p5/a9TxilYCIUj6qL8UGIYDEJ/Cq+EjLkDs71vK4q/HuP5FdPCLSmO4mc
WTir/bY86VLpDcjpZZy3hmUcX23RxjyCew9q70MqpumMsuj7wh/EDoN7NvPGA6qW
CuI1zmLsOnKaOSfRX0HexmOjFQ2mIhNUxaNr+JjBropsBet3FDIgD+jRexpsgrhx
XNrPxiTNoY/uTFnsxXTnQZdVXBc6hOMmgaq2ShFXZP1MYJ0x0CrFomQ+gmFhjGEN
//cC6VYaUCLM9bGAB31gH83OXDc9hWeT3WshQMLmwxG8w2rXtp1L5BCfcRFM4dp8
/WzFzv6BMdCHSM1DEq0KH7x+fezM6DWFeZQRGArHy4cZNfQSsVEhg1dumetZhbbR
I8Q7oWMyiP46809rN9HpD/Fe+TSMXfqsi05NWRzBocKOrg1IHnyUmCEfcyRbg98G
4wYwGXw5PPr79Q+CXwA44YU6IKdG6zBo7OlXmdFHRw+yy40ZTMe8dFkiwd2eQsjb
1+RTT92Xou92oAF97itNQ2FyDCYgtPLKTlJJsT6vloFFUZrzb31eTPbxRGnl5txF
iiohexPVk3uQkCVf8hhtibQAKHX6hKPpkiYfExsGo71ky0KNc2An/+sIUZk7huJP
vBMkvZO9jesabstsFFCXVc00tLvGG63CgxxbG1Z3d3C6CYek3eOohXE8qAw+VyOr
usfV2LyCHr5nhngFWx21WygTKQ7aihFmzQXS3PclvcJc6Cuh6at/FJiiAxVLn1Sb
D+C9u+/ciro9r3nLzYkK3QJFsEaf2GwGnaIn3ik5JPLaGIomDXVSbveZZRePXA1F
8ms02OoWmCdN1st2fbZ39dt/hD9+Pp5DtwtIfzJhj3MPcGlZWBEBQm7F02+UZztx
BZhlPPVErBfiGpiaUnkb4PoGppjpr3lfWMugnXDpI0f6FY2+WH9IRBWaIe0xGGAX
E5zn8hIE5bVa4f9TO3+cFJ0trMb4sks9I+hHrHM75NYJnnw9VbaITHTikfJdxEZw
tI2bWfosXHGzhVwTnsHByB5Q+wcztt+y5dDD6jjxuc28MyjRFyO/enKP687bXS8a
H46NBJImNCck/NMYtlICsOZSu7V2y6qtq8jvH1GnhiEI2PM9+mj0qAcBpdu8ha0V
NbHTnpmVr5YR3ICNgj5XRSgLyQQd7lQSTvzEmWmY4+LDuvqRi/TyhmyuSbER4I8Y
9GPrE4iCjVdfxIkSnPhzB3G4G43xBnwqy3Up+v7eNMTKhcC3iFUlccOhg+B+QKrK
Hdx4zk/AtXlWXIPDsb8CydjYf7oxEvHOA5MYCLf0xbqPdiHojRAsmdxEbFbgyt/z
qrY+keroJx18vTg845ffwhfp1PRcvE7GX0b16m8WkrxeDkeohdZZSVG6tJM2bFci
R8uyme81Vxi5KLYxWAxEXxt4kDh8OPLQGteL7haQrYba7P9X6RbSToMquoScd+Qu
zjm3R55CN0LOqpQRiF4IqipyDJDWKC7vvhLHvEe7iTaxA2VDvtCwRjMmQqiM4fxk
xjsriZ0fK136QM+ABpkM3l9Ji7xm2rSCB9n9MHobZMoHO853b62poME6dyMrU2yU
C1NiuKYpRvNggxmdDncEQwjH2WKEydOACbr+zxKT8BeJ/mzV9QFm07Uno+wjCb9b
6v3bCEobkk2b5w4gQuY+uw9ErGukOAHP5MY8vMSDR89TnsYtakV440Mkd6Lwruab
mvirPIrA5YpaPg/nC1YNzJu0PCJa/6lE5PwRMheoXXpeup4BjA6pMOBmMIZ1TkKD
5KuZ3rXtPtNLmUlLwxW9o2MOE8bocCGUqjjF8UZaPnSG4naxyb5neibQ0fgV58QN
ZZcSjlNGwynfJ8MwFJRFndJf6sA+jRys1Em90HEYNrDL3QkEHvqTmNF/P2XNDwYr
g2kN9LNsA3rl5Q/JaTsM4/O1hoRxscomzAVW4CwOhHX+I8oJyPdrnQ9tMnTLVCtl
k96DrxOkRE8cyqZJ79fmF0FT2tjeFukvilijdUn8z63GkKQpDLetRCKeCewt/xzM
J609gn8TDJa8qbtQHrPYYU9XlUpj6+a5ImiybqjEllYfTFnqhX5b8b0YjIohZWxE
BI3xK6jwAKO2/ow9TpDSxuf6x5LnuMSNccxQXngFUsF9A9UsmG6hn8CAQ+7drIUD
aXsZGhjoqNvkrLmeWu4HPvb3LyyuqkQcL92il3IKowYnydTfE2TCmNnOxXOash8Z
A+FBTRLBwzWPBZscdjgESAU6Dj1jMApcTIGjIQLJoIqILjsJ4tSkbIRlhoOe4l7d
8UcxxGBv9pqc3uozmcYeosSiO4K8Ly4Uhcp9fE4N2wvkz5EnTtBSW5pisxDzdlGC
trUEN6yS2W1rtbv1fjYCWVlAHatX6lHcpVTpoggfv5wVF7yS+cVM5NzkOrFliny7
5xuFX7xTZDw5hIydLRdyUgzwME2DMiVGqutYQmROLbmnKbOm8drzD9Q4ql0W2tst
GGibBOL1Jh95CxZGbNCKCZM/tVeZZsaNUxpoW51L+eV9Qdr6KSs8M43V7YkEliFv
EeYQqLBA/CTSFNnFhkNX1J4iQIMh4TYJ8vJGZTWqzh+j+aHYXLB0qXA59FYjyXoJ
mrTnrsNI7kLgViEgEUtEOG3MAu4NeYQhknYtSM88ZgS5X5d3pdXHeUxJgm0n/Zxc
GeNaiQIiw0I/NKQDBcmuzVPtZPPggJEplN5v39/k3OED4XqpgLosNCVgG9bx/cuk
sAMTIF1dspVmlZagCD3wfosto+b3bPrkBb+3Hu0qtH1nAR93YKekCp5Joa6wu8t3
8zM9dGCWMJ2pPdh71qKSrvfuVRupHKAIO+7GlZKXUxOw8w/N5ai2Etk9xWr1Zh1s
EH5ZvFGASTuYPaNZnxsK/4eaVD0h+R9J+a6ebfr3nHAYP61dfgeGL/jCbcBSQw76
zFWhJ+mRYSKE621GPPPlLN12cfe/fy3HMVt9XLxlsxKFPeQTuikzR502pH5FtyWC
TfLLT4lyni2etx4Og13sitTv/9sSWfpaYVS3JeNZdaeTzMih9G6meQQbtDKaa2n0
JDJ3iMBHIckL3jk/vxcKfaagln3GIokwhUPqOYCRp5zammZiQRaKQckafO178m0/
jhauYkgPJq1yDAkCvYsWgUlshfGobXKGMXuQpM6tJnPtUIQq3DWuWBR01UTpLNqV
XVvBouLe0HwMMCgwn4Thuw4kj53uifgaVIiHits8q3V8SEEFpaNfMybFttiX1Ld6
HTeUEI3WoHvPZr7gEjT9iLyn0kqAZAkB/bIjHfYx6gixGEG4jppV9zFjaZagttsa
cjq76ajJooK2WtVah45lN4QG2tLyQ68gqWcZXgHVn951eFN6LJM9gOKDXcPqFSxa
vLJX7hUMM074Uo52aECfq6RkgJ7uLnOJ++XtMNZ3FBR410CEaW5KPBHGU+wdJxUi
17r6MARNg7gb+MPf6txUCFBufUijYgIj00TVAmqDi1xKtO0+1e5XH9jjeOXWrXZi
tLZRIjved4FJJfXTyy61YME+rjMs/l5DhpPeR5iHLe0DH/wk7tEbdmB9WrkHnN7l
DrW7LPvOdpGpNoS3qL2SGeisZTN4pevZWFtWAMScWmfUWsngbm177ngbIJIUByTc
hearaGSoKtKgceHODDyYc5ASq6LlVhBvtqhxPUj/ZT4z9FWWZ3Sa883IwDFP+x0N
mFBaUL1kVxL+0RlH4pd78W8HaLyUsVojkmP4XEahXagZRCQziVa2NGz5OitxBbTk
Z4eMfgJs19sLDu1PdmWBWMr3vFa/Fr9pVXK6L54bh+CFg6m40UYE+ODKpy4hKw5q
H7xfM/Bl1DY1SjI3K9M4Z2isVJKIHpNS+0PzmuiKUlhKleBuWVhrYDPJbTCQOUZt
GUoL/L6699jHbJmDKdHG1R0Jwb8UEGyALnF61Wy5X9llApxCy2Lfykiw+41DdftS
RL+snLbapknGEoexW+i+hxgpZsr7Rj2FyHmclGhx4WGHpaLRt6TsZ0yNKdaIaHjR
Cx2cHijeogNkxiQ4rF1EoTjhb3o2g3qVbXwpVTcz6bjDgR2eSl6BFKUmwweMvHqa
fC6D6dd11U28ftD8ZAa3BN6OfNJX0zbdw+hFp0UObQPfICQiGndteKp23gAxbrmx
KyIXfaSrYYK4Iz8Nz7t2JVZlmAOu7/YbsKvKz0Uc4XSaAFbd9asVGOeb+NLa55bT
iLpqwyKujrYK1MDD359zMAngb2w6BXQpbP8VIcydsVhHke84WfsMePfKys/V3gmG
tFIwArgbPaD2kmssglTPlsGFiRn98n/nM6VcQRoXZECGY0UlBa4bAb2pBGcucQnm
A7yeqa+6Ni5Sw9GRruv7Hqb68rz7dT2X7I7ybjh91Oh15NEBL6vPUqmChOYjvvH+
Kl7Vr4U9FtL6s0K2zYReQucQRrw4p+z6hE0YiL/My+JpmMCamqj8daaW2O4Nl2ls
WHXckXTmkUDtQpObfJgF5WNQR7aCTaf/xCxjZPbjMGI7YzM4+x/XLZHsd/xvQPEr
QfsnhWNmbatNnKFKD7cdEzdIK+7ZZb62M6GjbAeX3QxzzBCKAn88wm95/doD7oNK
6BmGWRpcc0NvV3HoxhC2y9jAqNGGZTK7vHndhCb30H2yCegu8M1gneONSx1mK+8w
b+MNXTfNpFgIdSwFYBe2vUGSyKF2CO1U5iBeqSZdsobKDdXMrjZVnr3I4ChYnUxi
dvm8VjDZkDYXjTekGNEs2pdFVreTyUcnHyiIoGeaeY2L/OqS9JL+u3R75NgIB34D
M63/fGC0Rp5GhhZjq0ax3uPNmlO0tzsxiBXowkoQuTwAOHz1hJYU8MjeZ+r8erv8
Zz+oHX4UjQmusXbPEkh2z/YHRQM5o3PVlP0kLn3LDxcP2+k2bRXbm1bHoLvBPszJ
LkwtFezJQOZ+sJxhpXx8J2zlp9FHKgczOPmOr1UgBQZoF22siTELOzC+K+4pzVYS
jEbSZfwePGNkwPgG/18Qx2kntJVx4q3xgFJ3t7OwQPpNOxXIpmb7mSS63ASzWT6C
XrQVlcrLfaD3odynEwzV8BP6KF8TrvzeDew9euf2nOjMcjzdyNFaQgp2S/UnTJPW
szSx/ZjbKmQ+qN1NKPKQMzUGZSCExJmTxzO+gkjqrFISs/HoBFeCBTpgCch6LJWN
vTC9+258XQAbdUVIiVT9XpwJnpC9hyJacoUdA+AH3evNiHzMnsXT/Kr3K4nGZbh9
i8T5izLeYG/ZLrFJsRTjj1n4uRCOjZd1ilM+tHqNWXV/XiX5GfRve6OeVTdGHu7K
0gN1fproRaFSmXYDtWBtopMydXYf/zvagQN9/TvxWlrjT8tawAk64FNTxn7iFmvz
aoW/Fta/Qm8hYG0plVJQIY5MdFcAPY1TNK8kyVBXKBEWE7zdoSOK58HK9fMiDQ6b
YUWPQhqTnLAIUTnFVEB6hDrPAc7Weyp2lsHujOKYeVEplof8G3VzqeRpCnCEM6X5
pK6yzX663qTbPoDzbyO3Aj1ZpmSZBxRBLWeSrBvtRnhdTh4jNUbOpuyCLELFl9WZ
V8iedjDdtNgXjT5BwJQmk9OSFTNUi3IeYwPql6M70GcXfGiJI2mB48au/sBz6Jpt
f3bexA//rKEiLLLK7GYwro5X7FWJuebmj4OKrg+Eena3X9Vcxs1a/wmMeLAndMGv
bvwhgtaXTuL48u/jsezhw0kPuuau2cm/kT48HgSz/zWhfTbPQoWHdfGBr67zGvUm
UBsID5gNrqxvlJL9wT2+NG6eqmoDUHFOpplvk7HbC4cjfR/LKu+rZia+SO+lSpJI
Y74zMhQf2zUlBdWHGxjP375g3lysKDHeSlyQCdc4YnSL9EBpkqMkRpEiLwFo6MWu
/ylNCywMNyRSaMB6pvO4iGYiIzzn9IsztiRM0vIL2sYKhnlnQfOUGj7Cfrvn5VzD
QCWYZvXIhZOk6BjoTph/G0PCP5emfkD0vlx7OZSBSLQvZeW+Rdu/WWdRZ5ZS8XS9
MWaAVLllHQca2NEQ4p4oLBq2v6Pqcr9s9z7TXNSd9+28HCdGoTunFIL1EoK8ANAo
WMkN0KEqa9ug/R2wMGlMItZ0kmFmo40uJE52qygG94MC8sAIcHh5jHb3QG8erFQp
oylTAH4sOnECWG4iSSRDh7Elob+7wAFJqA+Xy+KqlOj+1zb5Ms9C5wPwgY1SHjWY
m0CqvfSHH8fNGl8ikgyTKpt0GK6z1utWVsZCtEFwLgXbzg/h0XXAHXOOY2fnfDFs
AAGLRdEH8cj75V466ruZZB3TeTe2wMfalNMFb+dI+yhg0l3PIHDVvA4ZDxuE9S8p
U58teMns1piJKDQWvrBbWs0oCH5iAoxdQjgf7Tvko0F7xnENkqiIqY5UG19yGMGi
3zTPzOgT/f96biveZm0gbEqg/hRVIsUygtshlz5q85D3pwc/02LJa1IGbH1bUitM
j75Jj/Jlycvjt/tUbXjUUhvvUwdOm5x+S+H27x6Z05jMisVOQkV55Yg8arxJ5NXT
DmaIVgTmJ+vzMfAhoWO8nw659DAR0mL2RxbNcWGGjjYcPdscscKlpp+4Ko4iCWCK
tG3W/k9X+C051tHR9fmBoO4CRxo2ucalKOFEuFwFj0fqrDCdDso3YDHwTQxzaX/t
8s94PcJzQzRm+eRqsV8kWNlw0LMEozpe4jKzH+WtFnmi1aym7waFR8QiMSOzsLNA
lPfYeIu99HXNm1UQ7hLLGtxyTAdsWXOKgM+PL/pJo25VZWGU2xOjeVuoFaYPST+b
JBgFrigSerPxPU4uGr8HAoWKIRGCc9oRgJwnKrdJH/vVuj69b4TJCOUImC8L6Z0K
OG6J8MXNgVADIbPJpJu11Q/mpJxb92d/oVGXNg8/oZBah+s2FV35OvRTqm07ifSv
mdpl5Vcyx4J2f9GCZQyQ5MeaCG9gS1hLu4QJvHtRkkzkZEyP2Err7nQeQOlfPW/i
8HdMz5DUwd0lp/4BglFU0uwS9+Sj+4ZZputiyOdpA893Q8OY2Nd7VIGJRtBp+Wzn
Xm59TjAWSKdfMbtOACQ7y9W1aMxwOUMpKgPNWYzjlNxtbXkPkZ/a2bmXO/PexIoo
mzdjahmuNiG2HT3vjrYQd5djGPnIMqmJFbtlGRJ9D0jf/Ycj8u8uv131OyS97Ubn
6V2z48pzFu1fIs8AJCRE/KabDOlia4iO+tEe53D9jDuOu7BvR0neRGUjWT2npVEb
xcGj95baP8Z/99p84H8h7V6OIDem6Y0MDpjwl44w8YgH3WFbxYO3ISX069skpyj4
DtrPCYnvVA5feypG1eEfHSn6fPy+iUBTtlPbVfteOwI0OygOf7aakVk0Ao1xVzA3
UNj4rqmENBe4/N316HqjFeW3kuGhY+UA5vQUAAPxngjAI6kVV2XDltBHQxGZQuXi
aHgZmpbG4HKCH2avABAHp8m1fTUQF2dUQYx7dbwa7AAYuVxbR3fDLxZPeR87tdK/
cM4Jjtdz6b4nPed016Syfp0Xg2ut0s8oeL8/A9xXxgc9xzz25ctH1Bhcgl9fFvEV
3aep852SzvaTIKUmon5bFYEeyckCFE/KFUJ+7He0tp81FeYr1Ua+2z/giXh/ryPz
Y6BYBu3qoMeBCoU+6AB3OZ+taKpUmLVph7LwMwoFCvjWTzz9m8yQh54/E3ppCzCb
C6iye9v2Av4dAHofG3mhLBmkSnxKr31QFl3zUStpmQe/rVWDg53PfGh5tmzA6D5k
4FlQ8nElZwWkvwkRuGQ1s3xHJPjhHxGAAYhIwb1rL10XJR8gicsSy3BRQe5HO9Z+
GIwfODbEkctfmR10a0gVkNORwlbGACCyfj9AzEBtv4gDgGQYG8MCiXiSplJsjmdk
Sqf867JUCm5NHV5XtxG9ZZadAQ3lOV0Bufj5wmHd9hjwVRhK0uSgjZgjlJrXIChz
FywAZ8eXyXS9C6w5cKJ8XDOAE7IH3qUawDpdxXTvGJ3mLpyfX3VctRYBBilae5xg
rtuH0KLUKr+zVRCuMRi0AXdWxCucHIeB1CQmXRBXSiLs3zy71kSVsOXl4wChRyYn
OjEUAU5T/nO3XipS/iNjUfeFeBkD/FmfWBHt5qlDMGKffY87EVnvfWAApkmRaiNz
wtW5RGymb4+G6sZjrqlU3bXZooFProGDa2/IRGHUcTZXadMw/aXbID496W0R44ok
o1NYX7LUf6cL2hPIjTC1NsnZB/UxQARqDOyOe6EmM9T0kFyCBFN/y26LHHJFh2NE
DtpEb9ikSlmGyNZqTeiSCAuFtQldkuOphRki/1xUWa26jsOujmhMw19eTspDu3Xz
wiezwMVB9KsZk+2JJDP5OZdI4AHYjWNXeeUVp3ql+1kvkHoF558T5bwgrSbnjc8s
g+bpifOhkvlerKVGppEwpZC7fM6Nkpskh5J6ArZD23/wTmdkMDWkqqWqQKKe632D
29Fqa43NfCRen9iNuzIU8093QsJ8gJwWAOfOaoLCR961BWv8dwI+vW7EL6lmUHV2
d0+DG7S7nfjScx0Bd4Zc06bc5O6p5aLbPyDtptd9sfxj0WZPdDtGBcbi3KsqJagW
oG3rVu08nm8vKHOwXP3ad8jywr2TL8iaKmjiG21RXpQWwlctDRKT1LtZgqHypQMX
lDj1AS8NyuCQ/BG8yKlEHEQRVSk5zHKpN/N2YxU3nZHY/a18b1EhlD4iO7QpsRy8
Ic9g1hnye9Wc0Zb63ksWEBuUhN+b08L2ckRBsbT+51CAk1aQH7EoCn+jUzO8swVx
Dhjg3Vhc9de3mk8YZk+n0CyJ83vK0YvGfGnY6mun3gC76V4QxjQS1St8zOF9qhj2
oIxcv78bueu8ywOfuQIxWclGL8jFv6a5w+o4iu8cMwIQ2jZEhcJyAgk/ZSu7txTv
gA+Y+F5XIwJP7WeQ30SHUsVXCWKQMuWC6Opo77fX6ClPUC6byC073u3G8AvYRtEE
4omkpv8vro5BPEcW47przr/MsiIPY2qnbUfAJIBEPfxRALKxguYO6vKp2wvsKw+a
RAB1nr6CVVPSCIuWidkmgk6u80TUOCs2Gdyz0gOvxIHdCsEr9pnxBvHxbmb9/GO1
vnzs76IsNr2eBtoj+Gq3qlorCxQbcOJg2jeGkOJACH4BQrwVFmgQi4l4XoxVxuIe
s/UbFN2dmMf4VVfRa6ml5qu6txYBSntVv7bBW9+3B5+EWjS6D7YHrdtqAuOJ3RDx
8I92dl03S/hTwyjGrHnn/XiIDvumzA17upJPzIGefoeV6goCcg1MBdVGbYlqadLh
7Q/RikBK3STn5dK18QBCSlLDPygTEzaMAvo+WfXIgsjEjdwuEU7vgNOpattVskPo
/udehonTYqiMRE8tl4oJ6KotALYGyz1gfGVtUl+d4P42GLdrP6HmMNopDW6q7NOh
DGCTZ0e8w4QVCFoFGku5h7bddtH50De9+4s52C4FH1gOqkyZe82ASLgOk83bcfqT
1g6gPfZwHQmSLk9y3n4scew6v2vkyKNGKGcf3N4mKZGdIJgU7HEO2Im8LVTvWytE
Of6dwuuimbEBZqnddnv9oTpjBo4+rzy943OgJeXONMyUlUKBN6nF4hhndrL/+Czb
Sf9drfL+Mv9NSzdEle5hLnpUex1EB+ayQslTy7pSr2YFdguKc3sZ218Qp2gtpdlK
xnd6tnkK7UMeQuILuQPt4XhwWyV7ZiOAqjTqzk3cqzVVlqDcxyUa1t5UciTboNpk
TIZmFifnNkZI+6aKJE8TZOcTzxjFFtddgj7r/K96qSL1Lhf9tojReEKdKU+2vYQ9
Zt0BjnHgEcAdA3VB5tGQnH4WQ+N2g2bbsWjsb9fA28sxHpJoWQ4X8Y6fOQDg/e1a
uwYDNCjLQA2pb3Acs6a03ITsxgGXugkZbvry9HdQebZD9nOElXc9KZ4iBy7HH7VQ
1fLt5SKify8Hk6U5n/pUqrvAZRYJsa28WW/oDsyLKZmYZ1DVYWmP2zrhvKiM8Ku3
9uc51Otlw/I4CoHnh8wLEb6ycJtd4GhEbDPTBGuDG6n8H5idwb25vXRiDrkkiUqB
01sntHbDTU7rnpXFC2Pg83LCcBjxcrdDLAx9Nm1WkAxj2CyRWWf342yy2gGPFFMk
3+nnQIkUvU5KVyupk4gwM3lRSydN6NbW/VUCw1nkuFfZgziqiQHGZW1B9l/+dTn+
1+YDTBQWBfpk5GMSbkgNrmY6Z/3gHMlgC8TURsbFMfztCdWtUIMFoqubgE+rRDEI
LQ+/X+fwMlXucbrryuXq2b3LfPQV0cWZqN8M5WMSwyaCEs+hW8Tll+Et7KJBp0H0
s01N7rvcaJLS1XJNsnBVBaqzggEicMzulqdoUJYbeebhSwWHPhFhbu5qUDFh0ysD
KA9jAF1QUx2O8CLgIgBdvlb4S5/aaaeEctC83V3drGWBnyXkl2keSPZ37PSpxT62
/WkHlK2WcFfgGQ/W+mu1WXeuXtYX4C/EA4Gy43WxXt0hcBCTYl/Qke4nZF054NC9
cTZR4Kv+UgDTMGmi9K5PNXysCwnTu+wl4XllIgtbVafrh7cgNDkIYnU1T8s40qUq
VkLRYkgUmGd7nnoQv9VsEtFUTU/bUOaTLzNvvqXt40GQtgqylR2k1TEIYBMb0mF8
TD4qQoLDBe25j9B88DimqUkedtA4mQ/NibG/ftqw9xkYlu1Nq/zpFFe5F22ugNGT
z3bxfdj6RsdRg2w1zLPuaRUpWutGfHCirEJfokAP3MDozrYa6mMqmZqPRbf1hysk
7d21iBS4xM6fsY+sOsqYwQgY/O6MLJr4F3MYs1ae1z0Ms21Tg0Jkqs+GA+z/obzi
jL1uasla+O7QQTxpNkqs5Ue5tjMz/pHh958guHsAOwzlbXEEanDLyctDgCo7dSup
3YyV28n8CazC9p6Sa3brjZ8vWudr9wwiVgf95A/AY7FQUUbcsIVWSE4hNfzWJLfr
wAGH/IrfU76zwc3T+7mhNAJ2t98sqIxN4otuNfolhzdbaJmD6UTmh96tRpOCapLX
RLo4LSTXO/hDmtkhTS4/gGpzTRQNtQoxp05dYpqBd8D1Jplk7eMyf4drQeRCpUU8
WmNTUNJrlh/+YnZkW5Q0PMXkGwlgjsFg1ZiXuTWiiXduLq1ndgspCTHw8wQJYF3B
TYU9tDrLI6rWqojQCDTKl1yGFKnvF2hdMlZsDwsiKvZGrwgm93g3tiXO5EzVXZm4
oaFGiQfvkAS9B28aCQbm1V0ToB9J+6T0/Q6gKJhPlRJoXwEHVjvbKK4Gml42hkkS
5Kry2h49zhRFcsc/oax/KtjK7IJXz+0/2g1hg2hNthCJbhpKmnBNki47Ymphuh2I
9bWUsToPBXh3fQMJVChqMdZIwLcbQ0c57blFZYSZxW40X2/ccT4ihP2iXiYTShbW
tU3jloOPDugQchcw5DPDzAtaqt3MyQHIzTvBiFtPbCI/lzdTM5RI4SVhGHsIx/Jn
DHdZJv5GU2lFoCooJfl+5p5No4ZtZnhBjHQVK2d/VLX2CGyUVkNA1i5U+vN6B3IS
ZqRE61Y7QZVT7awCtKZFz/U/H01ETBwmClSzBFKzCe1Vf9ZHwt17BTnsmxOvHEIj
7k+dAXX8LzUoeWnglXBYyU9tZGW/BBFHN86/IXxt9OQaEfvq2KqC87PdV9dLxoEF
V+x+3WyobJlI8SUUTQ2HY41tk2k6BgMM68oh0huUKD51oOocdgmEEfTyozmBockF
uCQJ/yvNpGgOLIy61fbHZoaU8TdFENBbMBgYlL6a00SprhLe0MX2TCZE6ah6oIa0
L7paAKw1jcU6ygH/pb29oujc1JPWu2aI+CWbWvvYGf2zg5nVeG3eo9F0eC9PvqrB
1g8MJQRnGkqTa5qHcAHxDZyb2daknF0cdk26Qrq/l7s52z2i3GGL+0TTavq9fsEv
dhpzatKSI7C88YRoHA4S96ODQ42z5PHFhaRlfOCdNHVLgDJQQt+l7P7yO32qAVCn
YKGkuBMyl3DyFeG0SGEjwZNCX8Z7whMVljV9e1AUHlIIzrenuj2LegZ78QAifSNI
R/Ur8D9zJQEDSsSONXR0NLe+bzu8W/L1eDGp1bQG+92iGzyA+0LU5JpbG0BnF375
C6Znwjlfw3vkIoFntqpKeHsAlzwf4iE4xADkCVgWX5jkgbd9jIAZQI7a+AEjgM4t
qAVS5zRob52Ue3mZtXUQvC2hX5082uxHnsq1BWvFxHaBcQVpWExqfxk7MjOwCA0f
eXyHI4Bwh5ZnhRKGPIPfYAAdha0jeiRSpD7wFvqxmFioRDcAteZLnEk3tm/ictZb
Lh5NQraAqXAIfsZEyc/h8e9yggPUITUwv9pWZj4Uz6/g6ctAPcpZPhGhPeXUe484
v4hIQpUcExsqn0TPoHQ7absyEkrDFHUqmEx5ItwBcG+omrhcsZ3Q2TNTSWQtMRNF
gFHZyThZ0nnc+0gGXvw14+Moa8R7zGJmoV7ThlNpgtfDVpnilHNA54huNX56/yuk
JsyqHQAY+JNvs5Su5jK5LmIq3jqW8vyf43VwyF8XlsnIW/e5VMCJw0k0sa+FyDm8
LhAnvQwz66tuVSwEdbm4GPGzlLp92Xo/mpc/FeW0jnTkNcZCzN38X+YVW9Jo3YMw
ab8aFQnIgUnPme6hU8kc1OmPF6IhBL4P1RHDbA46uJJGs27GWlkyw8LaxgvFtH57
WlTOtZBLt91MEG9hewHwn23r5+MXy2XEAzLRTooXnLpAcyAxSU0gyOzaRRbyhLID
tbECYCPe9R7r9Q5PXtrf/iakx4dHB3nueVUHo6oV+IcT0p2j7gOgkj/h1PBk+Knz
YVJMhPkDdyUhcvrxJX6J2qihtJ7zQ0xNLPw1Rwv0eYwQtKQE4v1EboNIWJ8ujjqh
iWtbq3O9bOlquWdoNv1UdcpGW9VJCYGzlqJyNse7bc4sLJRfWMsV0Htx1lpY72Yn
If7A3X8ExmtLqDmEox+dfZvnwsXZ/5jvma7tAAPm/X0ysVv0BIuWWIHqeVoLJIk/
qBBQHLSgd57GZw1m+EGwPoaQ4NDv6EqEHsQukZVfGO7mA2+FbbUylgk+WhthbB8M
ptd36wmAVd3TdquXSFjHwLkxxZAW9cRQ4cr/p+Fu5sPoV+/qTiWBcQ2q29CnhKIj
16SjmOVcgBy1o9uiv4PBHUXkaVn0guBpEFra6f4BmX4YQdLtQg7etQ9y/6HRNptx
i6NhzyGVkkyS/8sPY+OBVhUvJ7KRWVO+8LeBxFqzFbIdN5vguYiG0XFX2rHWiFYs
XvdUeosislk9++capn5hL50ZHnK5yhBQLkczO5h+A07j9Ef2kt5GSL7wSYCurO8z
0elugNJqJF1DO2BhRCwjlRkfLxuwjb/IM5HJ0l5ZeDXNs5ZppvUz/oZs9bHnwc34
GAfLhJGRSDECtEyr2j8hlaqmyODZxynNYB76AwEWOEn1ETpO1W+m00tB6UiAr5Fn
YzKiNjpelXkoxysC7BmZ54rRwEo8u6SM845Yg0FlaSdmvvkbKF4Cq0HFeg5MMCqf
zg6V8zRIlHIdrxXCfSGXNsCecw4CBTwZd61u+vpEyiViHNYFEaCSDGkIurB0D5zS
KFgYiT7skxmkEnUu5I4nHC7r1ezNQCZ5FAuvwppWJUjEBvs1N6lYArUV2jCnvmOU
jhbLMaEQcIEafuq2bQwPfrhsysOZnP/i/XJrCKd0wLg0wTPlUOeGbDVQBSpN/c7e
XnTJrri+gEFq1qU52BqJoe2solRpjcAAmEDqRuH97xftTTXmpjpIOybMljU43xw1
bt9YU3yYeaXCzNHEAQOGACrpueplsFHy/nPAO3ylPW1+fcJL2HfKO+t/hGgdFFlR
EZ1pYsm+2Hgeyj1Sx3idn5/PGN/pfVk1yg7HgTNiZsmklneUUa5fnXHdJjXIe7hI
zQ4F7x0HeenpURXbp0Qd05dIQqbZamPV3coLPWuEuMOsnM6xCE/5OPk+7yVfghqf
8qe0hKiF2wqWD9yYZJjgu5xVIMx5rmQN9+5NIrdv+fuZQS+A2Ps3sdr1MlC4n1Yd
1tmdlc9avGla5tMnUSP0EK3y6ZtiCTeCn5nl1T7v2tc8U+KvNE3hDoGWnZJSZu5b
OgDnPJsDzwlvFthxdOkyTXmT2slHAWtaUyN/QiSK3H4IAQZHRnRTN5+lTW++IDHv
HSZCs/I2zpMMS5PO1JxQV9i3D4LjFOec1gbC0coVucBOzwCS7fIirt4cflGbN/9y
fU9zzlNXQMokk1MLhWdzpwCgouBZYy9nFGeU7VS7dqFs9f3nD59Hv0aBPkDWbdjo
sE7MP1dsQDnFFzTWG0IplLlvYQuDzn5tAtE6e2/NLKm2IASxAplRGmKOSAQN1bzE
of42UU409IvC0GgmODMUxt3/dCP3/Gq+KdJMkW2m3kpDe6FJlU2DgSgmnKkgRFwK
T3sY7CBkagd6eoTo4HaX1CPuCpq249UgHupgVbm66iwT/0tCat3ZONTkyxOrA7us
ty8HftrSNv50JqMAPyXjAZ6iGk07BvReU5tZXk0zkDpWt2GTJfKjx7gvKz0fAOOL
tdC3cCcNAkmhhJA8/V6Hvpy49dFb1rbyFxsv5rL89aGwsnoCKDt5SGwDfhPTguLn
g4UKLM9Mn1bbfl4FCMPrJlupSqBdlHnXQDwy/G5SXGWGvBbAfiA3/vDlvLfl9hh9
wjdNYjfIt8S6z2tXZSllXFujYPd86pZCcNL80ceqE6yiNIYnWmrOn0S+HfZkmmA6
zlZ85yAOIZGZFLQ52ZP51KMmRPL2BWseeCqHE5hIQ0Jhig3zOr8345A4D2wuDEdZ
iJQ8NF9ftxsEQ4Cuo4rZhDoul0GD1zH14NG2Wc7vzJ9VSE34uoka9/mt3WGx3SFb
5XRH6QxeZxSmOzQUzqtd2t3getBv8ctEP2OpjispzS3cXg1WK21ppR6fKddY0Yi7
f8jbwJVNhBdFs8HRMX71hDlPczMZHqX9Wj+i5HIqJ0YGEY8Qy87tNEoXGc2pp2oU
FKO8skKLgtD4KTm/bZyuuNb2vEol9IF4knJZHrcJnvwW6MvgdDgr2bETL8iBxFuc
n6LT+KmwTascJbuztbCw+vmWFUYq/g++sokTQro+9BSEJgJ4YCUwPweV4/jR5aMT
sFSsmx267TKdhr9XCs86a4r1w238Ly7wToCs7ltmjHKoZcmTBaPFe1yg+yIuUcZK
bwvy1rrt/G49Pm2GNOjVphtZjw4qtZ5STfcsW0BbYaFp3w3Yj/47papqg0n+L1W6
CDtsaCL85PmosL4C6AagsbKgQdneNIhPUO2NXTggtqeW9sr/UDyLucDBPH0XSHCA
xKLakESqyyU01r398LxyVRUkvmK3691vyf/pf0yeCR4UsCMzKADoG8YQWNyddssJ
O1tapE4S7AaJbM0osZajscPglkpOFur0pxRszyB/mlYSGp+G1q0a1g3Zwl/qv6w9
F1rDhdA3bkxEZwWHvN5AtIccuWPZ10Eoklt7q1CF846EsfrdCcIZypF8vQbY5cd9
Ot6Bi76ZQ/BTZQHNEjrwU0dnHzThDJe+ZheqckamXxbYhOXMr0tDwrfZRo7nalv/
eaJzcad5OzC3Zo4hROogB4DaqWhAV2jzO8B/i0/nQBUsNFskiFy/RLBeaa0ugp+v
OSNusMyeU1ud15LHE+AkrA248qEYaF9SlCF0vtNHymxyRPE5aLIBARh2gXaxtlNP
AC33cSLcWH6ygKcOpLIBL8Qr329I/TV3G+FF/zYqjBIz87C7axW/LY7G14BREm77
I5T7yNlgjf/hbhJm2G4FuLyAncX+RH6UhGyGg/Puq4IZ3Lx06xDF3Yuo9QUyea6i
lwNBNWnuvhlv3AemPDBrEGn88eMeeUtzWKOy3bmnaM5a4bvsim/EJC493EVbUhe0
7KESSANqca7mp4PT0WnfwsAmaaIMMY0HpruqmZs6kDRpmIfebju6AYDqDneZN+Lo
cob4gi5GQQpR4a2qIXUpMgKZyuplpatnyfOJQIIYGtlRzB9e0ANmZ3VfGXr5eCgO
XfsHJvOf54aIiPa83ROzPN//IeU6c+rgyD+UC7vAW0X5c5ghP4MRaKaji3b+w3O2
rYTWDzkAfBtNQF7JqPgsULMsTt8Ey6mW/jHlxHo8qs6/7Ufj3P477v4lKTtpAN37
ilWHiquarmylVNAg2+tz9Vu0d3PoD1a0tSTImlzhZbOUlgck+oHXHPTKr32T40Dq
pEUrZodo40+ue69lJn7fNf+rVCtQWCxwUSS6GAA8nsYauJ0M05JDCzjsVBKHj4Oq
cOi0VrG8//VU2F/hEZVcZb06NRqrGENTvG0TjWXy/FFVCpEe476SsZAqz6OzswSI
EDwkOLeyFE9qxsUi5YGUWwRBfBRWVcoShwMNEgcNMCF1jnU3XkDQEFi91Ru/KvDE
TuFjhRE8SYJqDAKKHVQr/0DqsCZeQNGgbYYmn6wcnQqyUczbe4TNQIybwMgpuxi2
W1CHam4nn+jr4SPRnZ4LoXa6YulVgmSMrwyhEhOMCL7rwBni+vhAHS+t1qlDYoZ0
DSoToTTR/z+6pu4sSGlITwScwxhmSm4x6siblwnxz3Wre4B8KDroiVpfODUbd6cG
427+si08AlDa0uD3OMgFwGh8JIxojwF4cpi0Jih6oYiqxbPeAO6lLcxUbcGYTXU6
aoG2XUsU1lXY4q1Z0+YlPK4uI38VYUusZ5ZQ/R/Y4w+y61dAjOa9ty8rsSZkcAp9
eF/NMURqqMtR/7mhlPdmP2N04Mau1T5ie4nZYBSmoad/q0uHOP+OFYiXmDJcvbsv
H5c2kIUmwsnob56IzK1qZXId4EVeA2HkgC39pUYy7pslR/W8hTXQS7H8t2IdIUIy
rDmzObeziIyrCR+kxYRlFe8lMvQkXdexMIbFsfFgr/u0pPtnV3xuCAM3hYl3DDt8
W1HiS8qaymysjjuF0033OTjf1Fww4bIObXZmd94DijNAqLO+kkjD9KqsNmSdM9hM
hTJ3DKI/VlGVNhhBXaaFpOZqrpa+jNQ7Z9Hv6MaeFd9cdzF2Rpdjj4+WOAoLAMeS
U9Xat8MU5FKbcHh8BClU7BhJnTNl7FaFEnfDd45o0DHEGzl3z4dL5Tr6OJ8Kw9QN
g9wcKziSIMnV92Uioy/wTrZfGCbRshBiE1wR1bMFZPwQsh8/2FHFI/JoDTDrNu+4
g1U4B9XSch9KkZ4N1wRSUKTUtMn65zU6JlIWSqI5njZZedJJuxxADfhIo9AfkmTP
rX2MfjqiG1USNi8t9svN/zBCXcPoG5npdG6DMxcGdpKPnzgN0mHByZQQysdJ6Txe
+o+wCUUVbCtQvFTAbsRmmLzE61YNGDz0/lLAfRMRUmjpZPFjqTmJvzDUVt396tJW
S4Mjd3do4M/8YHS8jjRj+ht3Z1fX/NT+oXaKA1poEShn+fr+9z767PQw8JnOJkn2
EHdtWeWEWYfmkbVCmgG89pD3DrHrGZJ7Re3JvhJeT9r8oOpxUq6V9Tz8bcWw92xI
tTk2SXt/P75+IJkdHRFI6zfcpHq2C643cf/9+Yc42uCz1k+b1XCkNXKde85kO6aS
0xHfZoeSoKD9XF7nZYD09lgw2ObN8WqvOC+KsoFqjX0NF8Gh/D9x/UZ9eD03fteI
qdlwMyX2hEE0w6MFMs2gaNN+B1lP9GMxcjNdS9rEfcZNVG2Ix41VsTruQqd28S+E
Lw0HMwllEvBjM5NywUIKON+jFG5H7YTBEC7oMTkbrvXugekMrWptrBG3m5VGTCXe
4zRRlOnYxKh6NtThpKuFPoLs0uI29EE7P2frpPTHk7POArV3sicqj+3f4vWTNnqk
26hf7Pe5rzJ0ePcsUke/K5ksJSyJpmAPA/dOC3vOO3PKufrVJouY8Gry6F8hMv/5
YfNhiLtKezLyvdhgMCy0azfMMRszj4GQVdriHmvsfAW5xB0R/Fh/Z6o7Aj/8S1K7
LLvNd4PZv2YOqbqk6Gq1pQifwAF5p4tlmHocDV4gyT9zr7I2yOGdi55k92aZZi88
c6ilyEAQP9li4wv7QPsRni7THN8zD4vknYgZ4Qmw+OOA9c3LGfYGisUrMl71cHsz
zl8fK9c1TIjtbAS+7mLN/aK885s0XnXrV60PemiWVI02nhUz5GdgGPwaVrQxrAhn
ZcT7uQ3Mzotf6AxZUEWT06LIWeeyGwoh9TObGK7RffurVTBrQcXKkeVQLo/DMT4r
WpjOKkxRBq4MhTHiMWj8tNfP0m/T3ub+FyTn9SKxUUC0SEaeDO20s/Mlu8iYWmV9
guYy/nyJTD1c8gSQhJlT54aeyVuciCu3+xJIIFH4OHGX5jBU7b3WGOoiVekjuUOv
wyg1EeCdd4tqflO8+Zmcstt/6yscI6dNmDgA64UGxnXnward1p/Gl0LmonACOosb
QF+Mf/Ae2Z9JCtUKVylSa04uGfdKDZWRkFsqGwy9pDkzhtpjrtZq6cKAXiGrMnf0
rMdnopf2SyPeiyTW6EX0O2yMTeLhL7LjOLDO6wdoT8b84vgGz5FYHGS9i3SfFXwj
W3ilah9IltdDsLen6h8X4/bPdj75foqFkdD06TA6C2NZJ5QiVcKPQ3VVGra1EEBY
hXcMOQ7m5ET0vBxdoLoSPVS1P0GE/wo/KaBr5o/EwGzF63I/YRjgMuoZFoDKWVJJ
d02obyXpHQqOF67U18li6iDkWonLgYVUfjS2yqzDyaHyES3T1TNmRIVfPFxwjB0+
zkum55ktzfRtgfBrCl646NXvc4ZEd7CLZJSntKSMV/Qc8hYrifR5mEm4ZB9Bl2Za
jMvjipOIVtXex765dSHKv+pl2xgYDmrU9eBhNSK9Pcz7sm6lT3rwRYqbef2GLnTF
twBAOYRtY8e5qZkF6xFV0CtLa9VmPKAp9aesBc0l1kcVmArMPclVXcz0PRTCU+J5
z5vFbtMHS0RX/b+j0YpvwjUph+UCzU9ixaGGFMEwum3AVQk/EpiCo7o4t2T14jlQ
25rdqdm376UGLmPyrUCAK4qMOWMwcOrGA6p0BQY5S06PHAl/8JcZp5C5kbFTWoDl
MFdNsCSFXZ4nL/5TX5IKJX9Da5yzeudarThRaAoCjdaaToY4OT6ykpFtwFzJQLjf
f53k2+MfNyi/O8nUzJOzQWEZ/dDJKJtgxLqwn7reSwj/wq8vEY78TlA8jB687dj2
UTd3pEhBNQDP9Thamlt11Xl6LwirUVZTNTzIC/DLIP9yRIQEfz6KkQFQKhjXkHXN
4eJeCAO1X7uWWnPvabkYBffR6N76GX80M6n97tEopdbtwFoTa64NAxXn9ut5xJlj
p47+a5EEHw/fTWYGDyYeDGURKC9pVFR4GOA10z2zEdX4OFaBBbao4sKiLcsaVrsG
Hj/y3kEpmTpzjEn5IT8vNfJkenLecuLokT2F37Pr9kRySS+up0RKjr12soOVCJ8f
UcIMkIpgJ779XZQ68euE2+/WLdE5kFWxkl6OaXcA/8WnO78zRi7uxnDnVDVtJsVk
8k2vzYMis7lM9iHGUD0HHZLGi0GHU6yKwsFXuRw0/a79utnRPRFDmu4DZVJRFUrG
KUh4NC0CzEJIZN7ejreTWjJYHCoKo5CmlgonyiJi53VN5TynDJmwgYuKuTL3LyX8
p8lZJ2YKSijWK/S5dO9v1o/qbI/5x3r0Pb7fNZGr/EO3iqXtQtYvMTFd6wU8TC/W
GDXwpLNeOr+a+fxmBrdp4yAB4vzrhaq5DOrdIfDwmdCBaEh3M4iyL5Q4OPJb1ZrK
ZIepFC2ZKiqOJFlL2G2Y3DlV3TWn1hP+cndvco9YcuQT3UPD2+YurBYVoDEfRO1F
Tf7msi62W6PAWB/qZOTF9hLCtJvgCsE5oLFkvZGGX/KVIm5oSFDoH/ejNYyBwO3A
xw4pElAdXiNB92qAvjkZkU48GpRI4PfTXWy4EFFfiaVdStCad9bGKUJoxUdtx7NB
9PjL8a3LzyDjap2OVjz1Cw00SvthSYi1yyMi8jZkp6deTXNb7RsgEiW1LPREyZkn
m8T+njLBm8Eph0mvfO8D9KcU3n4PIG8BwBy/+G1Nsgs99gsM2MP8NwGuZYyYlIgD
qYCPYBH6MyPq0rjSTycBE3now1fkvilIcdYtw6Vj1xedKx3BLICm0Mnvbg55cL1v
UUjG2T+B+FeyWTw6U8c/B74jIUq5idymeyzXx116Ow7nvu9SIsIvdnS9ynKnfPFn
iFCmJkJGpUuqdNkez71lK+JLhrVzJNhRm0Iur+Z9U0hvGO3q4xBntC9J2qreB9AR
kTl72r0jH8rz9Dg7lp/fkjLwGuJhzIOUip17sGVKoqw54etcpGceP7TumIvAjbHL
JS+oLb2oh1ly6gdvifdQdi6090FBIbKTmfBYHCUeOHf9Rueadv+hSn3GX3xvGs0c
rp+ZgccSoJEyr2VRETc87clgyvAeuZcnE8tvfdMIqxGlyxSHEidgFUw8vvHCqR6l
XBiEneFwUGTHZw0z66zVQwmxqY+EbgZmRWUaOv8wFTCRTfQ5mw42qWNyBnI9dzQK
5e+rwv9RRl11qKu+QLKUs/HqtxoHilrynixeUUUaHOSOOXkWNfwZsZv2MoAq79o+
YkHhXAGgSjcAmSiaUDZPHYdybU+9l7ySFs28iRwLhr4/lj1A00tlkqM7buIm9pcb
73FAqaCxF+B2Ala0QZwyTxv2ontks4LOZ2f1LqAgLXW+SYuUqi/gd6q7D69GSJ06
ImBwYgRo4fAte4CnFIywggkLElzXzsaM2sv+vNR3aEnrUurxzx121vRlRk80p4AS
GwerCfDeNIFUh1tlIoFqyvuPN6Qt5/dspfggVFBu2IGUxR7GbhPHNSQjsR1bDktY
Bgdxi4xn5rfduLzIG+0xKsN4lb1gXmBSmhIbQC47WaGzvEASyn/hoaSaoMeRwelh
+6e3hd+w/ICUtEBFIggKOabQ9tEklJyeqQDpRgCj6LCLvZP2gniLbEgJ9CLbwKJV
cmvzTMSltce945o8f3M6+bSDDv/jVSZDGaalwDWb7vU8dibU6e5aJHG9DLfUXokW
jyI99SLb46JxFbnlzt7a+03uCHv1TYdZRNvRo2SMEl8pMej6iGVPHoS00xf69CHb
n7pqEhFYdLFlzhSbpcylgaNZEFGvH/sQjLLQbGirbY7fAIMeqBdKtyKPObLuR+mF
wLRYLnob7w2nxI0MsnjxFJbzBUJejhZ4lmOOpKH9XRpJJa4NZ8BOT5guiEzHEr20
QkDvJDeSjiIwJ3Ozr1vOiNbke9wMwYAi2yJdq4PNtN+vGyQn92uGwVJ5XIeaneRQ
CXxFU5kMVSrexIMX7mI87h1GzPX5MWIPp/KM4SSlXybFbgq0wH4d/jGNS1W5urmh
WONOQsVBiS0mLlCxEwyzUqVMW1K1W3DRR8TuJSlqq95OhyJL00SBToT8U7mGGvZd
P1iiEBgmPoEh45k3TpL06R+70V/8lxjQRCDvrY7t/HjD01l9qnnbuW4hZ45JrSkH
WOKOz6bmlG8PvkBuWfmCZ9z9MW2fzclIZtG2XGrTmab+ZTuja7FvCWuEvqK6FcYC
UEU9y097dHtDaVkHhPATpBMmB/OP1R9Kqa5oyQOQVgzWzI66tx18MugF6x/zOZJX
0bzuE2aaMRLxThDqdXPCjqx2vaUXDzkQn23G/71ek5JvSj0vytf8y1xsqEiiUWjV
xb8aXmvY2aYhSuuDcCZ/CQO5y1uA5FfAPMyVIhNHW+JkWw4CZiCzU+yCYCYKbb4T
kWMsiA71pPsRAdVmSCUqqC7JWb/zySn4H4EuHgHLyAynZ7jGgZovj5Fhe9yv0Oct
oQoyd/k9IWaGeSOwUgpSy4WHaqYp8xT93+8bNSdHNNcNO0ZoH3zhVFjkz5n2meEo
1cFbZlbBOu00jBXOBEggmr5fTKP44WSTIpaKcer5BbcFdKLxbIJevEhd2AebSCNt
n1YFJsEndxX8qtPF24LsMRppmIna3LzdjP02ktlttycZAVkMzbv+FNvgFFRMfnCH
R2v3dbDLHa8vWQWdIM4eNPYfOEdt5yG0Fno1ONwO3O4/5F0XzVHROxivggf1c93m
tflWbqi8ZI23oUp3C8J9sSL6SQjDsTybqS920BNaeZTfnpoLRYGH2cTPWXOtpR4b
bym60v8xvTE9rb1XoDKJYjCqU0HaKUqAfJKnQJPja0wjmIY8xYLFS27oE1J73nbS
AznC6QlpNAt5M/u0E6I77+5b/Qyrs9ZyMrxfgPeUltJJnR4mYbydOq0q5tM/LBIt
41jgL2AdB0nJIloa12zRHvWnAlb5BygfOgC5m6BqXvTpX73MD1jK+fnuo5RSxR+f
yMLD3Chz0ZOSBFrovHijLWsehsjVbCzwV4JyCAA5J7mLWURywfoGwr/KP+w+E6Yk
ZZmOXCQym/PLe+ip2nCHpLaJxWVF59RmOpe/+qdz3A0brp3Fk55RhwVQMmlcy7ym
iK/GXW7avitMQ3/DBoy1VQMafQlGdohBAA/idP3rvJ7SbgkC5temMGfkGG4p+9Fk
p2QaFEGh9OpNU0iGqAd0PvOoFhEKdWeT46ZW7WoiTuk2KoxS842DqJdMO6KCMfrn
/dKohOV8alKKZ+Uu2rEOTZGyILHm6f21pfPpWdxpBtY7LSZHAj3OqCsYPcsP8a+E
md1Jy67i90UyAFUeltpjllu+qffEkoQOp/MjYqGxk7ed95GfCT1WR7WujHKL1qas
1YttuyFEMKjQXCwV+Dt1/P3LjKiO/RX2JuJUYvCeWBHthkNc0vCzXVOQB4RQ/aVk
TgrxC0U4zYbrMJrjY37+qYeet9tXGiIzrpVeAAczNIG5BVT9gdXkcTgOo89dzhjH
IE5ISYrnGKIXz0iV79HIbX20/HxDDwJf5XmI6AnTI4JRso4cww3htDtKTcJy/3nZ
jBAkQgEutkHvjXOe0lP5ZbhqFNEv8pC6IRfpy/DN3KBMSXySEN2lkKpWh8Kf1iJS
976Q7wT/5YX+O6tT+MdRdcJ9pYLMNCGjpymNj/E6duaRvsc8JBPzmjulTmpTnyn7
Z2iODnh4BcKyGZNXNXUzRDn+zhnk/AL0XoOYXvz/vgE0SblqD7jPRVubI7WeCrN4
7j2uKxjm8z7xYZHYTjKtyrf/+VeWBtgeRSDCDK5Ei52I4jFhleCxzswEfaylojbG
UmLkjPAfKydNW1gOFxDlL6AmZtsfa+VOyobc43MKX6MbqUg2pNheMx6dXUXqDUPr
ipke1+xvOE5cW3+fZzCVBeLVFZre7InAo6PMSRFcWp/exQTmkS7eUf8jT9cbLeog
cEynvzkVpdHFrKUZ/qAdbR/9SvB1WqTJd+o2rWTbCwnRmJkWGz4dg3e4zodsg8H9
mNSCBBqcCKbOed2pNS5NjnUvcbi81AeatxSzz5PUHpijvQlAguyUYHaqiL8es1xB
RAhjcPtfFk3b8+wIiOI6gMb2Qi52SywhJ5xvkkpdqnewZopAYs7CUhNVkgqq0nY3
GoL1s+DOdqHjmcXZTODFONa8rAm2R7nDIadR2oM6XctQX1IoLehh3aK7oXyPv1Nn
21NSFGWUnTFn1SjwLgYdxcD0sD1a8U7Xx/G85Ly/jTL9v7+kZr6MxoQ9uxK9ph18
qApDQHQn1A4HIDT9wtNlkL6qUeKKGP+nH0TLUbPqAB1zKMQxKiy4kfzFjY3t9EDk
vaJ3yZV5HYORs08IKyLJfEBTqfM3G54OWwCwkl5b6ku5Z58WejtevxGIy0kkv+sZ
WZtleHygW0tfm+IrxPUZ/GOtrt+IGG5rXvT0I4IGxZQ2xCvBkOAmWV3T5XdzUMuM
DzcWPFgTBldG2xdmebLHZ9mQPu06+BCAArkn3NrU8zRqtn8F7Vj4qG5+L6sKmnfM
R8Siao8qXyIvzlwcIKOHAdX7NwSQHnZeYEnC0J1K9twSgHT6FHwh2LuDz7/SMknr
8dJZDNJ0Doqfz4VzsR9vGpjuRCMDXv1UjscYI94MwczuwI1+StBo9jj0kcaX8J/k
eyS+G7Cec+xn3DoQb+HRz0ykyBH3/oQZHydBYaWaT6di5Rx2W4xFtJXNo+uIsjJx
wMzXsFIOBBTVJUGprh/wmILagFMrGzUot+2YGaeRFcGc+LVKv4KjA34c9qvu8HYU
h5S9nbGZLA/4Hrg3+LtxPu01W6MfqkUR6xBhofgR7Sq7tKT092MRfHi3/XpTWgAF
bTPLRMW2wnPeBG+AgADtTBje2uZiwWvIV64o37vFbICNlcjucDfkIRi2d3fPbp2M
m1u1YgtuootxQngI+OvmUEpPBfCWuInDqySFRhTzLCmjPreOIAugGKi6V75A7oJO
YVDUKJE2VFKMYAnKUxz3wzNOrhyAJ1VMbqYifJoZEKSI1f8f24+9NNmSO6YmAXT+
hJhF+boQHwZaHqx5J+V9E+56nD13Najxz3R6f8xDXDkcOyAy/y7B3X04r8wil0+T
FmiKP71QkUPeFE7ZBK/TeMz2UceGE99YK25BcA3i6Ds8Hd+ak3n0Py8wjU5jyjyV
WxAP3lzDRZRuKABCAYiohRRBfnF/bKLCfZUbH4ICsTE6N+rVkca0C5sWyNAghyeo
5/zpIvH9qSLPFdhtAUGPTZe6uvndPxVwt876fN0O4KVTExuxHtV3hy9FGbMDRtYJ
H9CIStNDrPj59quHlMJHgA/CIzNyThC2etmsSlLMs9txIyIcCEXDEkQTgAH1y8iN
pcraSHCQwJmquxDZ4yf6YsB7WXj1qvY4Wfg5S878RjqOtbfIzEkD+WUDPwPVsr5/
4PIPzuTMWidQK8C+ocE5qKoYzH0YQI08P7WXvlBpOTVlnG0MjDoRaTcUrqkxa5mu
mT4futEMhIVssN+2OB1BvYiNvnBaCI3acGC72NW2tFuZJhRcDBnrsUq/pIbFVNIU
mHxGt/VYDu/ADPwRarBFAlpYwcfglGjMB3ho3FIKt0kHVtRd1du2ccUpZOQmel7j
kb4HvuakFucZi8THAElbrxJD5UigCpcawdeikjqBXoNVAHbtgm76KKqI20W4x9uD
6kgiFiKNBLNXcI+5+GskmI6AEMvofae+lhNBDhJkeRb8Aoh41lUHW6FmElab/qzJ
NgCly0wqBn4utz1/rig+246BCHIxn2yhXL0fjQS5PKHPZLvijq+Nh+kjWntwdxkn
Qia05iGE5ICfAk9x4r5ddpzEp+PpyxPH5rdTsHRA4gRCsiY+DuV2bDWYcJCZjPjP
nQDh2K67J77fy+a33JCkhm+tNFFgRFLu2n/2fAMELOaIGsIpQM9/P4aAd+7nGgZO
DcHhAsr1wiVRxhfrqJ1Bx1teiXczlB+SrQeVp86Zr7Cjgf/L3uBzdg1SYx5yBx7/
68C4DzZeUHoBrkahaSXqai9e72qzpQx7ktxZIRRqpXy+YZIne6U9KCHe/7wgonAz
4wmWHs9MtAq4b32IXEP+0Tkj7L5ygLs/Fbm46jS6LxEYew4Znx7dZ2nQPd1G9jxd
3+AzZ9zoSj7fesA9aj8ARctxHTQcT9FQxAr3pbay1lAz0tdCHPj7ma+/LThD28b2
dwi5D1HtaKIrcShNVZMjYVk43vJ9gNC1xBqaFBjGiduYMj1S4G0GQbM4hRBPAYBH
cf+xnNxeOQSNBDUuGljgACJVsyWgDREBKbJavehlxwkZgmg1wjADacjFyVBuKjv9
1UA0oQxKn+wdUgenFttsUgoLuWu5mCn5+8i+jj2BOUiYX+KAWTQEgE6toJlLUWi7
FbZ4LdhSZ5YDZkEDV33E8WRMHyBR+PFkvFgiLC/miXXufZTvKC6dfTIxUsD/n0jl
uRCd0pnpWT1xejpySqjKuMc43UiyqS3yiu9widRZqXyuPfwrPhkbZDETqSMjLgGG
0Qpop4MgaTXglqUy5OcdRcqEW2+/XVohIVZRNjHEAs+B/aRX12ZN0ZiwJFJto2NV
zqZ3ezKLJzBw7hi04m5dsezgTPO3A2nWBj7cpX2MVZ424+vNhIlJggzOXP4v5L7W
8QhFSz8T3b6cSlgkPxNtttPYuIaOau3IHjLQG/PqFvxEAisEkPgGcdZoD2rWD0wT
jDAeMrRkwupf5m2FwP6ChNIi6tyr00UZBNUSBUQZekRMYIKxG6UH4fo7BHpFwXgN
U9iVrDLhpi1U9HibfaxPi2j5AVRRkPWlOImFwQ02HvSI0j69xNbgGrEhDm9E2MsW
2QFb7S+S+HHmc87A527uAlvZzaJduM+OlSAYqatFbeA7dF6D1VIWOzUaCtiZggNa
ACLEUu5xbCvAr1EYCvH95FIczBfHIi0Ay4gCdIg9yfWEXKSEwkKXUxDg7d2czLEN
fZpC3O8JP34t913ua4w0S3W9Y7J6DN5sW55DazWebVEL27sJjcmoFg20BW2vsCEH
7Cmn5HBNgptugkOQmmEAW3Eve+r2l1vNtVFFfj1mFlAnocc3Fiew/3wrl/8TEyYN
HJN6zZNHzY612y29pxaPHD1NvjqyDdtl6sLp7Rc7SfeinI/HQCV9z65554WEH3TR
NaYQOoGfS1kOVOJDZiEB/eQc0JIk7OqvldbMcxOEmquXH4nEVP+OmtpUtoQ9Q0LK
2iT1Yk1QRAoUQpZrDADIzchd3XIl+7Nm3cZgeiWIJjZj6pMUVG/y31Vvv0HZ/t7w
0V8aGSS2QlEuzlt1/qTTxFgSrM6DNFNPto6YsPHys2dvD6pogkidp5hFuOIGKA5E
awU/fNEmlhYcMdXvW/UgokEnJW5q0o5XA4QWHyMgY+tqwR7TTsuaOiiV0iJlBlo+
Y5yDX5EJRwYilLnJ5nFTDUDKuo68GejdUF/bljvzqQehd1HOq837lACg+WTwHjlK
MBMjHUruK01w8Oe9QgxcPV+0k/FvwLV1vVjoo06nU2038JIBVbIKPT18ruYMp9Xx
m80kEZwRZJC6P1DxJJsbwfWIDbJQdW7njbncTr5QzMV+S590ICKCE+Nn5PvP1OMV
snQSlYyLYGaBWifq4oEyfJZiSKp/Scszk+6SWIxAs5mjPw2pW5KNQecnYyUSa6PC
pbw8XNE7I08m/5ImXYu85FD46KMLyiydG80TU0Ql0ZU+LGtzeKengVGlL0XeO6sP
1WfwLFObAX2H9CX8xwJK75a1Z6WM0EX/ceUY4n+0oZYbwA3KolY0Hz077D+LcLUn
XgcGqSmnIu8fikWcI/i0Tc6JFM+xCgax86BWKMNmoELn0DcI7yIBxWf/ZDZIDYuJ
u0wcoVtT/pxjMlJEbvX122kEgmkxYkSGhoM+fcFvkiVPg/8b7dSnDC4A3ckFJ38k
GyG8690AkVJgjDz2xdvVeYZH/FivOPGUyDwzkgY7w8AWI5HBExz20H7KJjCFhB8m
xZX1sod0pZLai91npPyOVMsrbj/Ep970Ht/Jd+zrzz42Jj/sPWE41Bv9XTQDUWVN
b9jYlvY6iUmOqalCZRCY0rpY61OUcp/9nqUw/nJZT4+6BPsoUwCU96lnqGzBsqpF
jcyGFDL8dgDBu4/BSyW1U38YW6A1LCOcmVm2IPBGSA2Li2eXtQtsE7RoR9tzDBhS
JpCtQZU8J/qb/T28cccoVS0xccHQvNegQDIKCnQffwT/3O7g0nIk29SEgJr8HkHc
LbajoLnQISdNCTp+Wgl+bgjiqp6zfwDaLjocuv7fcppjd5q0W7isxhPJaxVyGDP+
AfpbJlJDY1J4se8Un1TAQXXd1/Ytd2H2IxLsEeTSaDoXXNP1rYZkOJ4heAEEIGIK
eQEPrgUElCSkzChV5J+fzEUqMi6ZYdyO/IZI0VyJ4QK9iE8F9DGH/bvFGce4QV9Y
LgD/JoVbk06QWTn4c1H4f9xfNMFwRz64d+3m7mP9R+23JcpdgyJVebnlhuZkvX1a
cVWTrzmWGuhGupS+DlJqwkgDxJ9smwTNWldW5iwIuZWYrf80SzyAAXZhhWed3Sku
rfgfY7v+fV3rJrK3sEgLoda17aCl7/IfAUefI1IkWXbHAGM7MUv6HCI1jtOq3CXP
fHOHqF+cbyaaNWTp6W0ZrlzdPheeY8eI2nILQIXObPvTaUtbltbGwHx1+sqjGuId
w7vKl9Be2XSxrgzIoBWWMSYQMMgSC/nsbZ00CEZvlAueOlRQnu3+H1ewoPFvgEoY
AGM8MPtaAArgl6s26Wlgh1gjRtr0Rsi9HgdBK18FBklSB+w9Iqf8OwO/8m9DD+Ei
43si50g/VqAOh2LxGS9EXPWi4zkPsdkbQEl+wk43AETSRHP949sSYjJY+aB2mi7I
iVZSaaaWzC4JTNNgfFcozRHjGg13d2hiaXZ1vYkU+Pgxrr2DO1BhgrCW3pMPSNqG
A68niyonZ6Hi4XmG4eYRNFyyogLxO5D6nuHaNtcwBUp9d+JuLrTYQxsPG35wgw9o
R7Ad7AlS3rcPxRHpCYrOzmGxJE1r7WtLGho/zePEucFwuDoPB3Ye756lGtpKz6ap
cjvOLsuSriT62GO6uzkR3CURXAY53IjIx05vyh8zZTBmYP161LXB0wwTpRGqWjrx
xuc3pw6W5BTav/kaLCHiZUqDA+fUYzURq1UHWVuKvwx6MBq5ztSOrmXtvOXav93Z
Pp46+UEW7fl/+pGMjbLi8F+WHj3hpVwzDTjbc5cwF7OYXHYvRSlwZWGsktGzo/Zh
IbrxYCyggO9TFXfcvxHvDEpGCZE2nu4jha9NVrprzyeCfN68jOjKbauMMwULmJLz
ztl2Uxn7NDxeh9gljl0zTEEBf7S9uhdNVubL3qOePfTPD7YNDB32ZJYQK/H83/gS
bwOrXTVs0izjosNTIRrBuR5d3oYwZr2hOi9ypAPnfl3S9RZP54QsO2bOmGcbdFCc
/s9rJupAaaOXHlwq1Dkj9oekmPkKI4mPlxs9JK94YOf/1kNKDzQn4dBAX+Sd2C0V
JLiqxqrveDSifUfJIrsslJNGi5U/CbzHBzkXJpxQ5Pof+V4h/pVjF9AxS8l7/csU
oHTwOZtariOlTp7P8o8E11jaSp3SoDjZvsNeibwSh661RbwliASYqxC6iWpiEvF5
itsVIwJGJYhPgB24yaMk7ok4IKG+tlx+/Hq9afuxkXK+vLx4xezoUKPMqtwOjNzK
lQmsZ9OEbGu0g4Vi5EU7aawcjoXAQFGresp/EgM9OsiNKLf0wpmpb3laErl7PYf2
B9/+fYvNYC/Tysopbd4PpEWwafnR8SJe2Ifdu+ptE79pPQo50KHeyiK5jMawIxwU
1Keh+FAxnBa3J9AwawlpztukF8g2u39ea7AEafKejR/1IHHQ1o6C56ev/cZzfQfT
xiH7a2gopilTH0C0ITICWONUEhhdUNjkc9hcsFJ82UAcW9AHEWWpSCfDb7Tj+8CV
Mqw5R4WsnxoxKb1/7DgUP822lJEKFiPl8m3nLorCxaFz6+WeJwtH87JfJbt04IfZ
Yfsx2FKq8nlouZwWbJ6wCs1ux/azSAilh/7YIS/6V7/zUt1YxxO2w60+k8xNkVEy
rXxB1Mwpt6FJ45PZEhrnVpjVu3PuFWJZm5om4q6WU24fFkaS0V6Ff8j8Xh+VNw8p
yVRM0atB2ZoeAil//OCxR0Ld0LIGhEGvk5tcMjoeAnoOvUALlGtsIdBzB2m943K4
vYGUh+Dz8vFEMM7dcJZLfIcjBNZdxRzwBgyanUCvgS42ARfZSr7jVNizf7CpJFOr
Gs6psh5pG14RBqkLlT9Ik7Zgwv50ThJl//l+Io8j2O9DmRxzEN9QLlPWP4q0BZ2C
1JfuFPLKQ97IC2jt0SdqexgSkf82FcTYFqLgGc1Z2xO0hqg/9xu8z1qmipy/UFKE
yEhJoOyCrbvV0MLFAsdEr3ZiU2rcMPz1u9XaRmucyJKz5otsMeTt23antNZB0QK0
afN+s836RhyFu1Nn9R4fGjZsMbN6iWBQKThmVX7KJkncEdxuQVUgsHMXbDlQNSOf
2AgzUfByPz7mtBykNk0N50IwkMbSEb65HSaCmITp0QrkEAwB5aSTIwWIp3/LG6As
oiJeeIAMzARamM3W4UNPMlAY7QtgA4EkA7pT+m44tk5EgBoxtCBs96xV20mfdvv+
q2MUrewo7Ql+4SDq36whsXBl503TmybewOgIuaxFNSaP8plTQNk2ORhfzYl7hSbH
rFrQM5/y6dvxfIQizMeHejMICdfedXxLt3cxMTyweBNywE7fs+aLD4/CICK5Qf+P
Ds5AqBR4GZjzCIATOsTpNAiiVzVE7DbMzCJDr87iyOcbFKLadsuJjh+PjQplFvP2
LPJ1aVVpmFTWSeJepTEhYhUWEjDxRQaKJQHQU4qXBTg7kjZCAmByjQX2yFriX92+
719y5VKM/34HsFRrbjcRKK+S1jP0ieTg6ELslVybdPNQVH0tgh3PafRPk15qmUTb
EO/TY05tq1kB3AnNZ0WRL0qaSUX8jlWiaHET8tGHqgTYKTMa8Ak06k+dPHUt0y37
vbaTnmpNtzZNvdg7vCW83N/QDeTR0YzCRYvtoZieUvGIFV/rWEDumdY5NythNcso
q+Qqz7UHTHBd7ubDmJo6zoMKi1sN96KxNY5vVmtLBjiRtU2ImzNIahycG2BqwqrV
S+uwfLz8WUA2Tym/ihLQ0T2TvDeSujEGZPEyc3L+uCnQYpJYBPTBpUaOD6/84meH
2gshXxPcj8I5nNsiw3w9xY6Dgh6xnx1PcJrLpK/8DNBZYphYs6MeuKYHYat527Ey
2Av1vfQ1TW+9jmJco76TXNp6H17xG9uUVFL3G69dUGPVUrxLJStG5+1BeXzngqnS
p9i/RI/uPcpRqjnRAHKNKZjqu5mvqSfef5oC9E2vg7Zxi3ZVK5HW3Jq14lBqaUpT
b9lWNU/8NXm7umzZJ31ji4SwWDs3CkMYTYIbC4DqXx9DceitYPTsXzjfOIOyqQvV
+O9sFJGotJoTl6MrcqZq/G1MyG3wLc8RRi3jfo+6/ta8uclm5dsB1MfOC7Gxm7hD
UF0BEA2V781H740uRY3oNhbUWXDkM7i//l/estZGf5OGJzPkMdeAJ6HR1dEBrqQe
q6mG3Xhj45cxI8h5tmI69XRqL8vV/D3yx+OfVuGjVpAGANIx6Li8BQKRgctUkU8T
S6uWwfKuxvarwLTM5P9bb2rriCLuoJdep2YIiOELpYbaKd8SldpMUXJkXMFM3wjK
RlN7NJTTBhAK5u1xJA+KpidgSs5/KIwDTHmqzruK8BWaTB4+y7AxnNTVOi6ODyzO
ITFQQ2KnIGqUte6AoCoBD+5nZyQyN4pIAAc6s9u3ZUDNizGYJLJQG871BDBwUsSL
YVHc8ghCk2mjdAG2kTZlw3i4KW+37Xb5cwc8PFhM0A3zdOKxKTnnG+Zif/3gMatn
54bP9O6SyNSExiD7oGUOyefbidw8EaL1gv1Lee19luUNDh8brYL3UHFrpA/+63z6
thnSdOsnFz6PZxMahpsg+JJd85Ssf8DMtr8gTnosPntkQ8Y85jyrj4OrUWNn4wTa
4imc87adDK9Au6M3t58RK93tpzBe+nuMhjvvTasnnT8OXcI/0s3YPPyDmxhUmI31
2ljs0at8YOfSuIRNbAM9g+otITCact+E35VZJ86daJ5z4Q6tAFvKK+R2ZVdnTs70
uoLm5S1jpBrRstcAcyRotpnc1f125rz7edRFe3vUNU/DfM23H+lEKeHIh/YKKrW2
HczupCCyv9kyRbveEjTDfrsT60q0Mm9Akh5UDNIRMDwUDLlurNQVkZcH8f6qbvuf
qHZveJkuLi2dcusuUSdagF3aDTJHqk8fF2OQTbM8/XH34wdC7dsKMjarA1GspQ+t
InYDi40wrxcVbX2O51GH0CELkvhF/viic0Vhqaanz78hXFV90sZdY9k/xXHQLERP
6zFjBxwxNd7+2hSVXN1bZ3sRU47lpu5F1sn3vs4ofIstLrSaTyOdaSMSWWgvH5W5
Tk/eOtNUqQpFQn725CchMa3jlYwVLrfex6kDs4a7d1sd00SgRvVw1E9sqprqyy4N
9x2i7ZPBK9af4EAjnxrVjekHlmbLa8Kqj6A8pVSyR8IydhemAaGikOXPp+ohvxfV
K6T8IUpwUDNLFBSr/50R5FSS9YdU6LFd2dsMsENvsWuVqVcD303YVm01jC+v0ae8
9dfuvIKj2u2YgGv8YHLc7YCf16j9RfeOJIjVT1XYFS1DGOje04mKGlJ6nJRo6DZr
W8WqCnL3aGbZl53HPzQs9dRSPl7X8AWBgnn+wd9AsDjKcjcs2jiQzhoVF8jbz3mI
OYWZN8o4WrvJI1vd9A5kiv/xA8eksIitlU7dppiJs8auSf+lTm61mCRw9PVJxw/i
R979A7lZJzyFsyOwiodGcudddW4WZzGi1UkMYfP71pr2q0X8ynXOLXwpv42IE8se
e38wN5py/dFL+Via/x96hKSOL9+YTatkXK1LZtc5xijPKRLGcTZs3YRB674Ud2tm
kzkyQsJSr4Z74k9rjANj2YJQCG3OzjBrxsg6eRJ6Gp6fKhCTd8nQyLYYLLtNps6Y
AzXlmAioc9nHC2Sd6+onIqrn9GYsuZapLH4hoObUlVUgAlg0koXPviv9ShCoXD6l
zlyuq35Rgs0mMTa27cFA8Z4j+UuCWV6Cix5jbupH6OW+yYvdM2SQLy0TEbhM/5e/
L4syg4dtyAmbTSnmTgouMwC7TkxiiUdmVMzw5OfKKKm1hV78DvtbKpsRP2toz3rW
Pb1XwdWlBeeHeA0wGbyR44Gb9848Ox6odgneBpPj/Uj5bEuL8bjN2tFDr1c/FhXl
/i4Jw0PTnaWAl5xmx5rwMV37Lmlq+MzufOpsUAcrJwOQg/eofwzqMirp/e2yg9uO
kUCD3FGfbfNjP0jddRXnKoiLeFjkyvCTNir2t8kva90AnGqbhSr3DP6f8eDGq9UB
wORiBaXyb/6/7Q29DqQf1MUSIUwg2MNF4YNAG/ZNimx9rDiqMreE/zSvcwQxZyG+
9N+7tpE1m351LDspJ3wo7avyQ5/bHBkIeCeglISuzHc1ZmMySLrJF4nQwpF/Yzdj
TmyGvejT6aPPM1yQE2xmfe/0wWVN/k7QomIzCfWm5I+7+C8eJ0MzVdLL2enh8j4x
LyTO5v1UmwHjuXBwgcGfNe1JEF2+7+gG73FF7rxgbd00mIGmOV1a2ztAPvZC5d5C
8MUgUDtCmBsXeeqKM9iZr0CIurVO/i7sDlRtncwLFyhpHNLy5pRA+Heq5sLbR4jh
eREeo5tvY9r+Fg0LMD79qBjRN6uKK4AbiN6kOfgWHiGEfzhqG3pQgyNsSHUmhuJ1
bMJ/ErIMR0i1UqOsuzmPb2Yc8Q9RF0GKjVgcp6TPEPdRSHoborL0PkwhYnkDP7x3
mZsDCs+D7zOwZJy2XRLbwwWyd0tJF0GxKNGgr0Cnc4y1Mg7vidjh2Bfo35lwC+YI
ePPIQFGHbR4LSjWyIrzdCF5gIKDDreWhYYn4EZ4UvrBI1040n7Ka7vyqTu0MZ0zD
4Oib0SwKFuZOQoxrRRvz7M2xiBDjJjeGb418nJRNrXB6rD1Yck/bBKiDNFos6JCI
NPXW/7DKHEeSKiZEycgFqfOIvmLQ2B/T7Gy1QACSTKkneF6kCsxushQyUirvl1DR
IyxRvzV+aowplZ1t3JTJRdrqbOde7LpEmEEUVJIfbndiKxfN9ZFoOjphKiyLSHLh
zsqXswlgyx/Ofi31qNHh+77KXL1DicFqYpl/AB1tmRu7MVroW8Xcrd8mg82bWXKT
umG9AKbOxI4WI73AC6hcm8ME3Qki3OMxekO+PRacOEa3M5AN0lETC6KXO1Fir0/o
fB3wU7iX4CzAqxcG+a7CDnxcoygzg8TuUFXfhKzzapgRfshsPQXx8L+Spsf8LCXg
mNj5+jQXeL4Gxa3vYGVB2toPRezNBYYGKKJUgcg83cUeuUvSgYDRVytcYJoddcFX
usTo1JEXO/gBvx5io/B6JGIpzp69kKG/bdvgNAk0SEJClBU0zPPZka20EjhMhDHa
DkQoPhAsJ4+/UmUeLmzgyIiveGV8bzFKpdpLS7AMoz5q3zD9vDDVDOsht3Lp9SGB
HX5DpzBiCTaGeAKxgGJvzLdmDIOqWPsO/SNMT5WLPIf6TPyG0kaaIN+jPpUCQuvE
TY07HJ5stF6IvIz/9JazNi/7CNGOQkGXtkRj7LtGaS84qB0Ui7Y/MLT7ILaDjufE
ietiBd72OJjYC241pchMAv7cWk+LXU4Hk+h/Pda93cQo+JTENYfmWWNkHS8OsI/j
dl53DlT3H29P+lbn1aarSqFwvZA37+QnXr/XQjdxbUC7iLjYpPzLXsaVxM9y0/kC
10Y0NpUIRlEQXoUE++LYlAr1jE6Udv4uyY/MToF5TBF/6QkI26aCZi3fJoWRUv9y
10QRpXcgbVFOSaWELBIzfyvHnV60ZsBThqKjnrNkuTnIZ3fLKrx5gOQMd48ZzZiq
ABvUF2P/2eXgQle+aaflHIq6G1Uv+W8r5C6FtuleBxNPI/yMMFbVPa3XrZmx8QvV
DFeJ7+ixDR15wtjiy97oVpAMGndGXoUTgmceu5gLvSoaPeXKdKU4PqpoHoVVhP9O
b5N9U3Bc2P5LGtsunv4F8zxiJyAFcEC/rpWOdHzzcpNiPGNNL01vqLVJFmPbvlNP
nsOoSAtGx3A92vzSeQp0x21/8ihCwCw7xw+W4w6hXnSyfKaY1vZHjUeUmTYQkzZJ
8jZyEbkzQhgoUvH/LNetL5lOmn3CYyLBcMFeJ6H5S5qG+q3XfNFa4Q7N+whm8nRI
dw7Bl+NP0l+7amnh0KIyeq0q5crSv9QjaHQmt2U/c6sEF73gPFdnWgV18jO18Ph1
wz0QcSuXlfaYpqDs9nTxScK4IhNlBFynNx51XePaf1GhnepnOzzQ6dciVc2EwmrQ
0BOB9M1wF3b/KlyCrDZgLXPromazqe0TxvHP3Je6Vi+q57O+XrQu/u6JaETvBPDA
GS9RD47+3owbEwE6M7YZmPqjBYKSMQQlus8XavIbAtTK0ePKmV+ARiJ+5pFklSPE
mW+YiAP9LnBlf++iaatZxAzpyVjcCF+SFawAGROOztt4Zyk/mbeNcq/J9EmJn2+0
ognH0lDIGneg1TKJ0dgHcobWCkdr9busAXNMtF3Ske0XjDF5ISKu/fzZhFHapbX1
APQsDHHoMHglLBty6tvZ17XU47UMmTSO2qo9IZvyng5Wg8UxGLv1ZjP0IzsJGS7U
rrDIJ2YKTrB3ul8DN84e2kIhJatHXDGyUdN1jy96DUJncGvAXh/KPKKQLRqwU7u0
TMszi8T2qaj51B1lx8bzUa1E9vpp8SpOjjdIfEkGvHdTeJ6c+0V27jLM7hjMX/6a
DnCnoo0n8V0XhL5qc1cB1ki0QNzfeMC8xELAccofhKdWs17Hb4uYhYTV+uNEEvGU
OREk4qrH0FUqHT7HqfgxxbFdHQE36k30TYNAIHY5cRG89gPeHr0U9u8tjs5IQPGa
4fs3fnts0GBcrJonF6blHWQReJ08gUc6SbJ86/GP2QWCZHblEDvpGneBUoUjSBNm
4OPm+iiW0ZI32HY+MeTFSCCO4Hmf0MtYaL3kc4UJ5UGg9m4vKbZiZj060bS5Ob8Y
rhHYQoNdiOjfQ9JpovagE8C4Rv2rCZFPGobGQujNCSVwWiOznYCxam7cqCc64wiB
dQGiMMTlKNO3ZBxXUtlJhJsuDxGiqFgbTUQBmsOEddEOOowfV/ts6ESkK2YZbzEX
YBmQBZyOR9XkAhkfPhoYwyXgS+Q9OROCmxsARrMTs/gZWEowViCIev/yq7pOjEyg
BbmOLJrq+JLRvvMYGKnFJ79+zjqf9MFDvofAIVfUHYkwrOexiBWlC1oH6u5Xpbbu
tbc3pn9wwp0+4oYotZK+6iWt6q9MU7flf/F4f1n/pfCp7T2THP9LXtt7hXwi8UOS
pPId9U+UKq6kFjNWrT8QIU7ZlW6OrWPCSW1UJPEfkWYWK0Qc3tqzJw4yfpYuuKQ7
54Zpu+8HmfopTjtXdGDfZVsyD9QYcdhHpAY29RXV3gIpLTNTxIV7bHmez6p335Qn
amclx6grdGUrdLeBv8zi3cL0as5JLVZDBi4uHwgRKCyvbbpTUzBUNYIvNF+bePME
EPBu6vb3+XAQc60LJ/yqjTyVvChNSM9PpykVTCSXG0B5FVfnoyghYfwL7NvaqAUH
ToCxGWUXXWFkfqMcmEYfLlJKYFKKUVA/eYEC/UgWW3sSnv6I0xetF+lcd6baxlzN
rJRqDh6zKdunyF3N2jwZqQ4zevAgznsNmIV6UKb6L6r827shzl97aTE03Rdog7ui
/Nq0oVYp65H9n2BQnDUks/0HNsXd/3ofy6mR0I590RdROriWfQGuJL9wiOGD9GQT
H/eEVaF6S9ji94Ak+xmZaEa9xXc8sH3WX4unEY0XyTKEFr5+RzwwS7N48N72tzdy
PS8BHh26GIDIKdTdLxP2FpfTX+nPV+5C4iQD10+ISYTfiK4zTL/kBtS7/P4q8s50
UOZUR8NmlojbtjMPJhF7oHUni7m/r9NFXHqqFRvzQ5Aaay+dqCc+firxHQoTGjhk
j7RRCA1PGSzrhuniUQiqz+sojzeBoRHw0TvXCyYeh4AMuXkDbK/hR4Y92tzEbVb4
kuzfnj0WEi/dRe+VUxnslMx+s6+SRzygSrSDh0/nB1l+yJ5znKXjkTGeQZ4+GT/A
JzhVwClSR2Q4Gd2Kcfc0E3wWTKVoGrWWqxO64k2o3nIRVI/eu1WKfZ0IJd4dRgAb
6JNmDR9pgKO7cI0tVm3iwWgpIYYVIIXdfeMiVnCw4+v3C1vg9QriL2Dqm/WB2lkV
kBrORFg+F6uJ0cqHnAv/4p7s0ZIbyX3J98dMgEE4Ka0NzxitU2/JPa91sjP9uFF+
j4wGdjWncQBkAFczoOq1IovCV99R+W3C5gRNiStV1uH28em9u9e2XuhNimOn8Cw1
HGOinlJ64uVN2XZDuITAyGkNif9xY46AEaLYJOD5OR/AHexKsfvGxoBAHBaiT8Uq
eXycx4GVG91womjGp20SLE+vNYdcJHvpzB8cDvJALVHL20SFk5/3ULD1hAzukoEk
w0Get2RyiClnofKXnaZMVgMR1MZzLO14+IGIbv/+LpeL35GKlMzzeYsg+DcrWcqm
/2+sWLQ3Xv2T38H2XMkJiKuOsmIBZ4DT00PLnP3mMu3IN3rjtGowl2phP2i5thX9
tDersQ7va7QiFrmVTkTnghd076qdZnALq4icYvqv/ACvQ/wIiLM+xsRQH0JSlCkN
ZNceSWDvQ/n63Xck0Sd7PLF0Ou34WN0zgOktfeXS8BsPq154y+wE/pAWB78OZNHc
/4DJzZQH1IggpCyVO5uVBZQN5qEA0STl8WgyABv0icVx/BXqOlN76jSNasRnjCq7
C9nzRR/Nn1o412F5318v9/lgaEJzbCa5m1WsuTst0G5P1eaRUFNiLXuEL0SOtsxX
staDSn+iqVdiWNL2XUFdPLgI9NXII2CTcF7d/Wy6CIHvBg1Mpn6XX+KNaQPPwenK
bCg3c42itV88IZlxBf8s4b7kKOfWk/Fj7tAJGrYjGgbahpWVbHh2ibErfvDwcfO9
YQj8z+Vm8DVhnJC7Sr4x2jVRnxKfMdZh9rjErMtgYf23cR1pvsay59jRx6o5Pjgk
PFoZEAjXLwJLNJbN1aP4FC0faBHDs9e7clzJvY8OoKLJmGN3GXjtOOF/Ip43QtaO
mKZc2oGzxuIaI/JgsYx+iS8dY8TFxybzXX1cRZFXJGFuIZnCOCvfR3dD09fO6pvV
1X3in0AtcnSrJ2qPzAqpkUxYCtyyUBA3yVKqCVGpvi6zUBRQSSzdQFPusyMRI7zR
12T5dMynoPR+wlugMk5c8SIBiAUGC9Q8OBJ1V3iAsifdZBYFvbu/Kios9ug2jqrx
TmfxqtYJ5L4s2eLCOV1Re/0Qk1kdmvLWsPuPLGnJSOWvDMV9G/ucrLg1GUvRUhSG
QtjpV0/TTHEkdqH4k9Ub0uo8fG36dwCHf8H//pXup70g+rZxqb9Aj9epxxVVXTkk
cNIau2fGIDlOII8CeDm7qeG9ltdiAzws7ZNyFAlSBrdAQDYjNCpF/GLD3ahPiMgT
LwSG9QY87TrQNaA9adYE0QSzMfWNmQk2Hzlc+QsuPcGqTndwFG0b2T/rLel+t3Bz
x7nrlEGeGQDOyFvf+bKbrSIQrZw8gvWU3tQV17/1sQQt3JGUxPKoK8uR/95LA75i
oXIwTS3LTJ7pe4logIDAOh9Quiu3JdzitGdjNMYAy1RT7rJ9iXptsqYMB4oirPWo
0CbgeQ23Izo926xB7MxecIP43YP9Klgr6ix8CPAuTD5afYazmAJ93d/sUWC8Xyl7
7Y27xen8If2E/+5600z5QiyLjv7owGCOQrLwmKRz9QhPrXO5NwswWDCLD5O9OYck
l5Z+GcmDtlUMAD7KsS8oK1YcQEqcxSqace+YKQV8U9WDTwnenSmtzW/tuFsW2bjv
5sgJhkN1d3EhKNuCw24yzV9bJk0Tf+HV/UrlNmC3f+piz4tanRy8uWFOUAHbNVw/
CefhlR2HvCTQPGObJvNxGPuKYz+yHasXsz+fFt8NFd/9p7gRdXvSd8lmlswxQyu4
o53aJLbXMfrP7IZZiBPcCbJs0upKP4qEa/u/eGIFkzwsi6G8VjccrfD7EwtGfZlN
z9502B5k538DQz7zb3whyICksXnM6+2ykY4lQcCszGPQjv4MRaSzhjFGPEmi8bod
X6qzb0qOaUtfjVhVhf2Nn7Xd/rqYR6XHaHves8fozMOa8CEAAZUP1an8rIHjdlzS
qdZcfQSvWr/t0+wvXYUrWHDOupI16jMalBsW2WDsbA41hJ1hCrEo/0Pq9UNS4hmJ
Y+UdNBwyjzgqGaFXGpxZihmuT2uGjBBPBUV/ykfDvWl4aKi4eBiXR5ogO77MUqUy
ZVgCZcKTmqCTbRihDD7o19McuK9cxtNT8SQmqS22NleUGmlc/X5lh8C3DeGxGLZn
2kgXtfWbLoGEOJJ4+K2fIMw2xm0K6crF9xtDS8eNpkd+A46pM/too1jFC1FQWtGV
+DNCJAP9CFFd1pq2gaKGWnj5wWFHexFR4xQ5sflz79LwrPwsXyj1jjhrHFApsco6
hH0YPE9YeOrkdkDiFBpRUzEpA+UnKZLqRYlaC0CmWE/r1vIGCCt90fn9WO38odwp
Qw2i6BKnK30yVT3tlMubsMSc0L3/kcPTsl53zPr5w1FJUQk0FXU+EogXpmfS7sDD
i6kjgNx5JyEh3eNm1EqskQziHVIGisv/FGtCPFuTWiU5CcJce4RaD4SkIhEZZEAn
FtZpgDoqdrOLMeeFa/TQ5QESJY9r082keKCJKiSuyXTo4p5ks6I9NTPvWt8xt4AK
Z5zqedsD1K/texzrnfFbjAh1lBIZ0PrFoxBVBKXRMc3GsxR45PkkAXtP1RJhDx0R
rdkycPJWUHtBjIoLVDSRjc45M1g7pqT5HzDIyDaYi4w8WFJ1pe4mgBt0cGJQUaWC
DuGz0uu9hGhddZxUaUMCQFFhggN2ErIWdSJ4bF46eq2I+x/Q0+LCxB1nzbzInpQe
ktvC3YxjEogU77FpnJogXd3lAwChxerM6+qlLOlbgCnltspPQkpYxludR1XPZBgd
Z/d5dr6cTXMk1gxCCvn0MSzQrvsL/PjaiyCJSDT74ph/6COiGFY+tjYopHwVB/nA
r/f3CxoAxXOQexRl2H2doSF1nmt0pNMOdAgDmvwsF61ZOV/T1bRqBMCqN0A3EJW8
zK7pH6zwCdE2SFWzi+d6GJQ+PlirsIDmRfb9JBOMzMeM3gjmqfh4rTnLUpW6wIfl
65TcjmOfvup600zJI6+sj021Q3fjamjU1hdKcunRsyxHtQLIjb2FsFJNam3DGdqn
m5Pa0M6DfePQ1fG1adpSUmSAjB98BCx2ib1LaDJ1H1czSqoHln52cgpuydyXw8aI
E6V7JVLbXrALVbWs4u3uouy9asmX+ETj+epgS4xyZsM54wkhzfWYQo15yEwbkxGc
CJFZ22dNE/yGeT8v5TTiu6ibrCOH0aXzjyCfGU4trIoZjzIDvbhPXaJvO9md9Bii
HUKnF7Sg0ITzcjMKrAhew/+gm4NGt+MXnnlGBlLTmlowyNWh5ORx5dv3+cwKpFkw
JfNm6KTFAfAZyiOfgsAU1TX5IPqkYBsgPsb5X4xgCE29+P2bHajs3jtsHycc5g6+
Cn2X2AKAP1vntuwgUITtNHfDIqzFCJBadOVzmgTD88CfqkSge/x94oJ022ADAveN
xT7VFH7dgApIKSZTqfzncH5ICLcs7gsRLCTr6Ds0yxF94svKB5xv1rQCPXy1gBZ/
fKoxQxXG6gsppoh6RlzdZTvTBpGggnFQx2Hhz5gdHNXTvTRqBK5Na1v9aM5ZKzx/
DhsWhB5kXyrf06n40qzR9EpcaTiJSjfrUcRdxdn13rmiBVk4Vgx1sWwZDbmHYLkp
gHBm4XcHl90upfpHjsV1fiEJUBZWkTfwr9hp1c7fb+o5VXF7PyyUEK2ubrRTYA+w
vb8fv6gK66i4Rf3wRv/hAIFGPY0GczIAm6Tv4181PEHeBsPJqVduJnj7S9QUW8JJ
z3aGp1nrl18oO6JCO5UaHxOTtBEp04gkhwVxSLXWVojaBg8jseLq0t8hDgOHOiON
KzD8niYkIZ3VpcDXy0bgo56F4M8SLofTDtGkwhbAZ3lNE/ToMR/pCcGaeSkJY3kX
UlWYVQro5seROZ8Jkl0c8HpLzhcltFOl1X4PfyY2AJWPEZn6nDR+mPN0Nqrrlx58
57yfoMnTxKy5536IauLrv0yO1Zav2jWv6AjMKDJTICAPDbwEoMxD4pQ2ZY+CxGv8
I5Xyx+b9TD9G4/0wGRCwhFCocydqkz4rxs7Y0Fg0BDvU2J2srtGI+5n+H1sLMy/P
3zk3naPWvBIKUDYr84ikpD4iSP+npCUxlaKQG9EUCOHYWmBFCuOztr0Jgkin8z8e
KOeH2v8c4DVvHusU3z0Klv5ueXr9/601fyAukdMwvDeHQJ4MQdjTfenIUTXquGjR
tEBAwo9+u8IU7CqYokvCit+LeX2AdRor0Fl4PfpWBQ58i8LCvBZFwXrHKEganriq
ZEPAI2Y5D8jmAJrvZlSAxFnui2NT+/kxjJvjYeBGQVa9UeiohA7kED9NyWzXs5b0
JZUJx4r+t7y/ngYgJbb5oRHLxTbLfTHfZzLYq1tVM5NyIPGFK3aLIfvQ3KFLc9PS
KOyli6CGaxgGhm4FAZQQSewMO6NjqFF3iiyrK9qZEtS+anoC9LTSOZPvetG5Le0d
EsMpJ2Hvjr3n6i4dbyVCDHf0H+v8Bku2V0Bb083RJuIFVhuTZo5EyRSo9Meqfm9L
TR3LSjMPiI1n1Pjk78EgSkAS3lFjBcy7Ho8FBNvx1uxWzcR2OoUQpWumvJvnrWsT
ha256K39oSavR1EgMLQEZDyyW9EwzWHGE2jet1mnUeea/JQ8qrcHtCt82/jNfj9Y
jYqjIOlAmLt3znSc8DugxOcNn5ZE4bqCAu0xD0pItg0MiDakFJr2aWzZ5JuPrtcD
HfWruAEfuyb48V3q1GrodXliYGalw5hdYHDmTY7dItTBTVKUtSmghtW2OL/2kqR1
ktBjnXvZyoc1RjNEY9vsFrzx0mMoBBQ3Nu1+txsho89yvYITYQi+FdRX3uk62fb8
VTCQtcXeYCuzdJ6nuko/PQ10dPmfDgJ5PNWrl2b2LZ/s0w/beFkCExzaaGJubmwT
ajpXgNqyhiDngjUFyBRNrs1r+vw4xV6oaHs80VIYq9v2onlwPv757V+GSpmWWjUF
VQ1O3GOFBdQkqn7n6Eybeh/Kvx/YDEmoN50zdU2eCDOCgGH6QQIeQ0DxwcT7P6MH
Hm7/LyQYkNtb38MVpH5+V8+QGxq/iccEzji8Lwm/5JgG7RvcS087L5aAenwmiWO7
xTf9KLElxsgDAUPe8v91T0K0EMEuzJ06ET75E/jabyMOFYjSXDvJdWDYwuiJX2Kn
S8tuJysQGjXlrVgK4d+wWmG63QcywFftsW17cHSv4K8tRtf4qzawTyeP1XLC5Ug2
lBm55aB5g5My6OsN5zoyf9Wrwi4dC0XmmTgtqbHaXl3UkBT5Fll4+50fkwSp5O9l
iu2fKodFT8ReiwSqm3IIG5TuY+irskBCfDgu4eh/ALZTloC00Y1gRmtRWksc7Anb
+s7BV0k56IdOhLfQwe0VLrHbQh09KjLdV6UxVyrzN0KKtRX4dnHEJkT8g/RrC/1X
sYYPaJQAvyCgG1AZORlffMACmyfY3zEqCUxjoyBacK1qyZ4w8zz0VWbqVMKM3Yry
Rl/LCuApi2inqFTEv5FTdG//KrgQy9PANH2vruz3xOSFzcXz9+zhPgDfk6ZjRDkj
2gil7XyUxwd3I4ZQSO2XfgphcQRaRRW8UIGtY4SYoKd1nSnvflRdRE/3UHhVNJY+
bCS83dE9pBhLwe+GnuwRdk6MzNNenGv/kdAPxt5fYbKroW9rjG28wZiYUYchMec7
0eyjQy5vE/Wg5k5Huv6EPTfUJfmc7me+nMoqxao+2SZis+/PD1F3YEBHC25I8/Qk
cH3qniftMEYt2QFFMShPB+0AM+lqqHCzyL6+WBiCP/x6FhG4SVw9e+5g9IPwKxo2
SlnruPQdzbBNcnYmXf25a0CQpSyBayLnmPT5XxhHXL+EvDPcamUOOPjcG7FuDuh+
tZ8Kifp58f2gBOfUcHyGLvoHWtdhN0QV4CpYMLjovr4j+k6P6d5OXNydEXRhA/MV
qJyCnuCpWSyHWBCtbY3ZZlaJlsq8ntaSznqpxC+jmh1ZTBRlEV0sGNyj2jiZKuvm
psK0gmQ2/n/UUZRb6xMpcbaE5aeh3VwGrEoUA/Qu6AAZEMru+IAro9EwEBA2C0jP
PbJwIpBbdbUMYqlhOc7OUEaIKZhLCTQqau4z51L/IQOaVKMrogbMoNTQc0c2Jrrd
T/wAr48hGgMzwqKD78c8doskcRhEknalsxtnayDH5Pi/O1r9y0QB6XLBehgA4pt6
WNiVzIzutB8yUKjAYjh1SXf7PaK8mnDPNP2ZOOUTRO9JwxWAIbYwJR7GVlOuaz+x
8ReXuJj3wzWLew3fGTQV+EW1Aavx+12Zqoa45iCAA347y2V8aQIctpWkZypwKxnx
8qpc0SQN8jDHgN15XtfTt5+kSG8WTmWr+cbw40WdKF/IsHPkecssta9gpJo9Xt3R
/FgRQOJ7194j16nrtgAUE+hKlupQ6Wflb9+E5pe+92YO3+3yIVo5HefC6/P4Xp5V
KxvaMSCQguj7jhtLihUxaPcpj6z3K2A3UCfDi7/VwR6ZtQl/Ep9Mdmg29PCIcmr2
UN/wX0u89wMkf7N2hAO1IK/9rsdm4mW6yjgL/Tg8PzoAJZIYywaMZ1HoBQ0fdwZ+
J+dECNN3Guym9/K3nbiXfwcva0mXVsqfZV+ZuOHhpjxWmlCLC1UHxB59SEVJMxSe
UwxiGEOsaqSUO3RcZfFUatCFGMjoWrL+6Sy2loMX5mPtBs3fh0MH0+fzwUDuqU/U
02ueCyt+sVXncAQ/i+h6nb+TrOd6+SSPktRC5A7rxLtNBChrW2ZAUojHWnigyLeh
TR3qTjRURlHXmzDaXyzciGWTOAslPkYe1mrrvCHgDeuRzUUlOn2D9zbv6XaS7J04
x+i8JCNLG6hQ/22/V1SG6ELW25NqF6oL7xT6YY754DWjQiBWdI8eRTKxOV2ga7z0
1LE+wlmlH2NLGMqk80B3qD+dlrUIrEM5mNb2UAn3PfZcEwIaH0H/K5gNuUksSfzW
5vo1RILAGYMRpRxUldarzZkLHMRr2gLh8+QB7JLx+Q3ENPC+A/cypoACOOMURkde
XqolQFmRGt4sUyr0ZvniVW/b9pG6hHXCuCHoI6LW4Dm6KOqprBNehJdJ7utqvg7K
t1WriWtbiQRjieWEBfBPWX8v4GZXdI4QjQXrZq0BzESG98aQT5lN1wu+WrrycGzo
zSlKbWO+rMgnoI+NSjIK4drQlllwnbzf0QSAVVZkdXECf/a8D+VutSeFxlO99C4w
oR69H7E/GbQVS/gMyxsmi8+26Avw8BNnYrjE5bTBkIRbHOMW7IUyAmpQHtLGBNkV
dqhoDrSccFxhUfZU1/nMDTiHQcI2nktZrPc7zXF1DCmEPFbRBV3SmOK8iIG1DRk+
bPIV/uu2ewkhwyQA3L25xf9NhXRGN+etyQGkchDSLCzhAcR0whREAq4Tm7hUNlgB
oD6ViRoWdFxaandyn/qcpp6k1Bs6lk03RqWfWa/ymGuoKACN3XOvPhJArkQChwkK
hUao6/TJLaSAov9ahoZTT5eknSHKbzPYX28hsUH5MAkUSUU/SIuXwm686vvfyOJS
iMF+taajn0cJ7FhC4eQwYSQmaKsa4ABvm4b/+G1XwXwCv3Amhy+l+XPbal9Lef1T
/c+onitccboKeWmPustzJYYvP332gNXoxNMO32POjCC065KuqsKOgOCb7XL6zkza
dPqbYQlRCPlNKFfPeh9WELyvw4jmwCgzWPFmB5KQS2pBjT8k1yWy5jUDV663Mw6v
ce/yFaR73I4onh/PRqyLW6qyq1ImmlcTXN6XC9tvMD/OetcDxZYroI9o6f73un9j
G3p5iAJnVzAcPyE0vCE5eJNcoS+htBAJta8wPwP6Xrn9cMm3zzC4ZI5/JqPrliUX
kcmIeEMxJA4wYPQ0jdqzdh3SCGJnfMeq45K6LI1FSK03pU/Sb3EYeVTo/K3JNOVj
m4DzXQ7u3AVvKIe7Cr2FA+MaIGL+boBDU4QGt5bP5+Rm5+9a127RPaMjl/Ki2NHF
LRKl2NT2P1LYssT2Pzt3xmy6b8Tf434ioju0kkZqkmp5krEbxSAreQBLu+IwpdyQ
gbbRs+BwOdP2r1iHnQbLwjdW9lxmOw6oW9X+RiTs22MMEEokGm49plr2oKwuKpm+
Jp6oGLnNST8kcegOLiS0Q5sBU3m5ovLAGerLsWqIlbYIRdAhclq2alDXDplkx0mh
qPu+ubiB3ApLbTBTZyzg/qQVCc+VFI1B5ENVs6q1MqMDfy+QVjG+uPno4B43zTm9
S8ud2JgeEFO9FHmuhZbB+yDIvRFUHw0laBIP1egUtmnSMw4EBL8T8NGKW0zy/y4N
iCGAv0n9TIf46SpKAvr0dkzGQ8E8uyUi4B7+A39AAFWXTpHYR+Sun9KT0WrQS5t0
UmFXMcGQpVN4xrDFQR8ylfFVHLgQ/nHfYiM/+P9w0luZhw2TNhdG6Kl6VShRj1bn
FxpZVAd9PneMAhxU4xDKhYgK+CI7y3Ij/wDfsxA9Z9pQ5uxaQquE553XXTbz2FpE
SfsyEaMtNugEQeakU1dcVxywNRrJVYv6fSRwJy++OLhkV6AOs8AoHV51ihtfpqsz
NIDjim1bnyNWemd6FPClfUJVfknO176lJBfWbVqVATGOAZJzkxDank2z3Jn1gXw7
JwkifeK25C6V2gpxaDpTAPWVmGugL2uUVofFAZiLrfpTY7Zk6ggABaZmJ4I5ZvWt
JCXbIOFOQ/uzD2dwi8eZp9zKxi1RyKB3zDcjPvjonsMaBGM+tqNcKTxnUOr9NCM5
2quYMuAiBIiKDmiqs/jA41tFVDD6/25d5dxRnnIZRfMo5XaT9hhKHb0e8Qfi18pS
iEBZ5/8VlYTv5dKMGg9YfsTnQYM7o1XF9zdPZT22wfi2jS1j55dKcyrRCYQt7LIR
QEHaHZNdroN7R1XqgNfmyWTeRF6+tjcEgL5Xso1x1HC7TMIYIenU98P4x5hcH8QI
cChwVV8smW+JYfPXn9fxfN10AAa7YvCMfjX4AZXor81YEzmzhAt8pZqvRGCu1g8/
qaRdKq4aAz/BBwvIJBsmrBR4FiLuoeQonIS0K8Zfy6Hw26bkjnA4luf5Za0oM5kY
CZEJAW1gNivEIIBS9fgghyZzXkmUgwyNaTYHuKYtrTYtDZKk0S7POj8JvzaoHF2u
PYRg0yIs7m5++bfQ3XEp8V7dEGI3VCPmfUtMY6WACd+WqNoPgxBw5CZy7HFyuc30
lSw/OG8H3QXJvcL/Y/q5rJXFTRkZ7yBLNO9ynBMK7l+ZjGHs1+uIl+8ltM5JWjh9
BMJTSRl37NvTM7lViAOg3upTrExeH7xghaub+gV87CejLneSdX9D1UMZqtbJgMPB
r26jIqETD4WTLHhX9V8S00zZpdYQsV0zsv6MFLe+JSQ+7E8hK8Gt7gQaD9u94Q/j
C3D3w09P4dKJM9T/ui6ZXKUcZHBUAwFxw4GvVtqd177QeKtlqQOQ00bwrUeyVyRS
W1obb26X2OBTQLgKLyd+KlfMGmxmZI5oGOOJxAIrQ6Zd5R3knxyaRjZh4JKN2zM6
blYYw1c8BsEyZxHESCseV+fV2oly2JdOMKBsBVoXnL23A4BFi0iihtNLhU6El3wH
bFz08rebujqftZiKyT/dD/YFr3wqxGxipRMhys7eJFq3lTmH7Q6RZQ3XwNmssuYT
3ux9XI+SJb22aXx4KPe8KvJKWu0ifvKpJXEsHGubH78YM1dilIN0od8v2cyXlx+w
heVXkQS8je/ATwbbOBTKR0lA3z/cXFxWUWmn+fd8UtL8yZghLnDiGKaaZSexSRcW
kuKbvm9etRxORbAIU1UsWNK6xX8sxrvjsxGWCh3ZTIkHxgPhfl1h8Ot0i7IN1qkI
e1jPNwFdR7vB3GRcfLGQKWCOnwIBUnPqDtLbtruRAMtlSqZA3hCwz8QO2mCju4bA
NVFpw6eqvAS47C9w7vC8pC5u4BBpW6eJSjEebtXoMay9SpV6FEF5Z2B7HUPj6ehZ
l8cP7f42f+mtYAujba/i9boC1keOYN2a1+M200ISCQCNEO0GDYfiWl8Lotsl190Y
RslqRVa2AJrshub9XEtEhG/KWqEnEWXtFgQE0HnWnGuFvNqE3+iLKYIcK8d/39SP
oaU/Stk+/2vSNlYNgkp+EbRsTsQtdqIUWKjYzZmZ8DOfaqbEmrXDmR2rN/uBzgoj
YbmTFYoGdfmLe8OvC3CTcdxqd767HmsOlRU5vjkp8r4ozfKCR+o5wPnkm/te75cl
M65et7Nvn6Oj85OTlU0VmDWkTJPmgGdlAUv7XWdUHaJHL8rHaxmzmLWSx6lEyxRO
mD6tMmaPt26mK2nsZdvSgC/xNgGVuhSPBSS/o2lR9yZSHWs/bQlbtW/tyGCLnts7
YcA9wTPEeTvEOhAqqn7r5VnZRDgyPEh702YXuWiQvdMsyiFUP0NT+1rjGrVcRLvQ
S7ye+h2My+XnHnuXPRUtwXpizqs7RTrV71kVJ8S6OOdzvx/e9l4d1SU9iQ/jzB2o
BognZstNjFjcV8qGvburtJKICq579/6aR8vmYRKd61pS4Pvm0eEbQV13hY30GRTW
Th8VelpKUgXRXeAIv0ZQ2DtETDYpSTZ3Ox1UOaHSpequlzYpYwdIqYoUHIbuB5JD
2GJe4so2Wfb68hF/7k16PsMmU9QIHWIEzYWRZb+/ptpG3b2iQCgZQRqbZ5EaD3yV
cid8q8/veFgF+HLSfxndlXzEMk97VepQNZVc/RBwt1SJIkxt8fd24SJ350F3gZ07
+5kfrYdLWWwkPXhngiS6fq1G25cjQvGqYLTqkx53LfDKt+sA4NoEYU/9uNZ1FmhQ
kfhsSDlwvHgYG/DoOtl1SuoyQ3QKLr5AJMfIp1SzemXzuDp2STuPFA+l9PZrb3FS
1e0qacB+KEQfE4oUfTUNoNffJYjcuH+TMa2q73TgQEKCiXDVMy8o+wZ/Mt69c4qi
t+jCwE7tvUHgHBSAebO10IPd2cHf4FKJ1kXVFra6jH0CJ/skR+BNksneYAmufZNs
vbLvCvaAu+0DoU87IBDSPGulGcddAcJW3xLhrvX8thE2mJmYbfNEBpb2liOzh2yL
6neUwHjVeTGSLLQ0KF9ZMiS5sBG4+DttyRH8vpdrUmK+kK6hiv5KjZLim0ePdAS0
9C/32XCBnF9Ok+Q1zMaFNoFP0GOJ5iV+uIqrS+MS+lYAmxYOrE9eJMMci1BHMS6F
gB0tfwcwrvL/uTyMEkQ7opw5dlgtc4bQa4UUqFvGpO/B6eB9W+0eVOdG2EImhahn
zYqEt0jVeWHuDEdp1bw3LFJMyFzSVEc0DCDU+epR5PeIkRmgb9kPeo9R7/N0BHju
1LpGOpa+rV1wSA5QIj5CI0J5YTUV3xjZPmDVVRExSgGAJh1e86HMEg4vKFjYlvoF
7QbWza6OXxMYPZbdRnyfPIZqzzX/5IBxjRkVaRI5aOk8/HXnH+yliXnc+1ck/c8v
IrHge40my3Jm+nTrsOCBPzOR3cU7maXB8d7+gdwoAYY4E/QI7FhwUq6WHohY6Pz4
RuNySk98exUQJ9mSO04Lv7iCOnh9VZRvcdwnhzRDbxKAIyOKrxpDFyukQvrcqYcY
RXodpnfG7F5O/waJ8LCSsoZRmsIm7lzRJAInUofdi+iygD1iRg2jwV/qzF2ZVWy4
pR8EhixfCl4wclGTtuKH8mTCOBy+Ii1T3PDjjaj+EyRVW+Q9PUqgQTFLDLhV+Vww
QI9HRgRyD5J2JdtTAeQDGRSlkp/Bp7Pj+lmY5F4rQWdybz+GLHF1JiRoA9SXo5IP
S/sK7D5Fzx3cvh4l7vyFGHS7rQsU0KK7eM3E1s8jCj00WIw82W2WVgPpnebUb2m4
iWwub31vA+ZvBL4yZiG4xQvPgiIvPlle/r2oxdJ+KBKJvtDPUwWQZCvz2lbukhEw
HCowsdS/CKauLBqu3WJ7g611qwVUkgFzZpyuzr/JduptavrA9MZAM9a/HmSkix7Z
UilSbzphvId4C8ACl0/ehiGYIEVG2em7J9nMeCqZbw/3e/UZl4LFAwDsCbPREWJs
BdOFX1o50OCtuMMhr3q5AIi/bJ+syT0/vR+881AsNqCVwUBr1WEOMD9TP/+42MY+
VuI02pQxhyYhDWjh9T+mjXnm86xW0iQHZ4q75JYs8WOzMXEBei+0dsfxn4CngbCd
3k8WB0ni61vyjhLaNqf8XqU/HcSDuVgZNalPgQWaTp/vT2LQKBOqOrJNuBg+M+rK
9pCXNU9C/ulXYtUHbJxnKDvqym+NXDh4+zPtEZjDzViTZotwNxRhJkpP/R8foS75
E/SE4jV5PvNDM3dRYBhAsHcEKxHdymdXgBrtY93KQ+Pd25IQu4uWEJqDpBXEm+lH
Mw4qBe1x/sxFBd/7/aIeAo5I+G2d1jok66FbhqV7P1Fy1q9Srxr+WvwdE65ELB/9
O/D3IYX6Ojl1HqsiVZV1YLy2Yl3UFbm7mUVvFzsOArLgPDiQOmcPResJHa0o3+x6
u73zmRFDlGj3zY6SZ5e7fpwIZKyqmofMV+fVT0ve+5G77Bujv3jHZHKypMWJY08m
wT02Sma2QDAr3I2gBgBqdBZc5LeHWdTJtgXkwwNO7aclWqFVD/XM7AryVoJ37wRS
sVp7/i+bFX890QrjZMiQYYyI7q9TFA6+Q4s/MaMnlhEeoVXrVUioxB32JArciWkO
cZPExTp6GvARZq8RnyVERZ3S/8TuADYAhBT7XdFS8LqkW7H6+UR6c9tCDqIJfLPf
EWmvdzdzbZTm+bUi3O1uFRlw0+zXBbcyhpNCEVjoUOrXYAyuEtOBF2WZrIFaAmPh
zAyj7k64ipQC0HmJ3qTCLOhT0CEA/OZ6qtuMUWWI1kdSG9wGaQp5OW1BxiZ0uzSx
RlVJZR++q53bslZfktpHI80v8XT8Nigev42tVrXlpO6+gtNC0fu8M4GYCVJPGHRr
apfob8NvdbnniiVr+Lrxdf/hXp1OldXrgzwFVFzr57404YyVDuIGqe0StnC8i1Cv
DyDU8QkGGgx/PfNZ5HjAA1RRoo7vaT27ExS2aWQYvT0vzaCRR/NdJZJba/0xG/AQ
2QZJrcSFNT7QdP1pOI1s/bdUIQIx3PIVQf9zcI0215lsg+tGZLG9dEjQgGmV7ej/
hRuo5hhYKYHHtPojcH6mzSmlO2ItUxcJ+x1TCfyE9sYxEqq+3xXYsfzfYM/EujI6
G3N7OhugFIXtEHjypGEIVISOtjNEmuW//OkQRHICQsvw5zfS5fg0B0KO/UQuaiZk
fTmKFolzUj99CFJS3cz4BI8+hZmijENerS7hM02tMG+ySqn/sy8XWsHUnirqM+UY
EL5cgkjFgsCuUXtgcPCaYNQb5KF+jmz/u80m8CfUjtaduQGF5YsoG/tahrafhsdz
wZrcygNTeWSgfJ9OdkXKwWPMesfCZfACXWmdjXmjt3aAxSaPx6HHMRMObsWLktn7
9qTaokzO21ax+BBufEhipJI+QXO41Bp16lzQII2cxulbJ/rJn2q/yfxfHNfKHfts
XPvfqutTPAlBnlg7JYpKZb0Bh3oIqiw4QS6opsTKNWqioCjvQQU4ShoeBh6xVD9X
rStTf2APYwN9VyCGR1WvY9fNe0zcAkX/ulqqUvv9gFa2WlM2x8T7lxksFoOpv8Xt
1QqpQYxasD88vF8YrKHh4PXjfEhZVqYpCz5NOdEUkHuvYJWd6bKi5gY0Qvc2xXt0
y1SVms8gGgnIrX+kDnwjWApekIdtpyOdmyRysbdogsrBvmHWwU4Rr5b3CHxAfJUa
q1k4drW9SFX4pmCpl1LuDoA9KevTbDkf1fnkXIy+cOP/zUuBHKtTNec61xdHj6mD
2eGAtNz6QnYzBSIuzJsBPV8UVDv3JOS2Dt2iGfrFKC48TNRLMIC3pyRGJFJiFRRZ
QFLor7UMoqVF2w+053FZCF1PfJrI6CwqNBfu9nfNwqVMnOts8zLgnBzPn0z+n1MD
u2D9Yy6SpC4dL2MrnXma5qgua3Lrq6iED5FnctSlxq2KJWdklJUUV94QKo+KL00O
QRX/HDKlsCbff9hczHc33p49StTMk8yUdVZ1xW/1XF5Lmky2wsbjgwC3dyUHq3bt
DQEi/k4218JCUPKm78gUc5pDpuRV27YbYsU6ZxXhiUOEuor5aVmfJ4RJIZ8CYEGP
7f30LH013HOJB+suG23ygTnxzzmaOuGKTi7ZgSbunoRGQYbl9JXcjdQYYL87PT/q
PEIHb/TePiueWEvsYP/UkkiDGuZVc8fAfID3nzwt55PDfnlZYsuOWfQnFZ5CckfI
yBWobO1Xr7gB9w/3NiXHHSrxZzr45qtnpWHPr/Ne9rIAsjisFO8NDDXyTZ3Q8QS6
OGfxc5HqsHgENkSNcB0eSDMrx92gBiSYBPvviJJCW1VIQc43mlgZowZcKAPbietM
0VIxvZ7WAYKtXkp7EgBUl6uJwxdD4BQzEoQp60/dQ823CZ+uGZ4ck/3dj+2ZZVb4
vP8C7ohpXmqA6PYa2wwgMjD0VWEvZ1vDFhb6cZhxMmCLDsllQu07g4GcAAuipNUK
OHv2pi8wFG35fEktLwcqtgPfxgfyVzu+B5SZ0LTKgx9EHO1ry4dHKzNeJFXyGF7v
fd5nNnlif5VVizfamWzMqr2najGYJlUQMMFfLDEIKANbLnoznbifx8mWsLuw2WRs
9io+8QBKKXCbN6rK45j+V0F35esMhfSLT82dfDUhksmrmqMwcrme1jIsHsbG+k/y
3520YyCyCffewu15y9a4BPUOwpfAYiprFHioFkW7WzX1Q00YwQl1AbgQQqu2/Eei
YnbL0XLJO3MyWS8y3jhRGT4TUoslI8b0fsAGhZLYfEIbz7b0XXAdtmNnHbArPeyY
Ex9+f5r95ydZAWPUQGn3YmExrxkVamTI3Rgnl8cQOM3GfgdQaAPtUy9mlHcVm8XS
4IkDNgtu5+D+X+CE/QFj/YfwyYO7y1t6jQPD1aXJ1thfG96/4B7X3GIRPvG2JFd3
CZLZnh3ItPS7qLXt2eV4MYfYs4X+sDAIocS6cKpD4k5ioWcd9tgCUj0E9uP6fZRS
c7kaA6p9xfxF3zqZxQsuq5I/Kx/3R7MbO2qCV5v4gcFN3DylEp4DS7kgb5YxLwhU
O3piKUOGx82yesq0ZkhjP6jlDAJpSLdtstEKUjcUJCMbmnPdqUu5PpYikt1IfUWN
qynslHeM80CzgATz4jmTSbG9M3K07pvgzCP3ablXy7UX+i3rBgyU7BrDR0aLw/xT
gIs09kaMXkcestrzR0Xo5U5gz6l9Eva2F/goazRh6kaBWFmU1MWcIfUTv3R9Emxm
xkS4suXNN9ussVzBZajQo6W+cFdZKtP/nvtKjLxpV4Ec0pYi3O7dGRFJqcPBMCcZ
3xBOUz0mD/ZysG6+N+7A3WS9D95b1qFXSYiTaLgVvpkC838JXjGK/pq8JzvV9p64
Ffzc7RJuRcS2S3QSxhG3E1D9UTzHfOI17ATiOsuF4ky9PxS44i0x+1MzJKEDFIW8
E1hWDLwpJoNy7BmeHRYcxc3yi+Dd1URyj8ML8fG7WMauY+MUqcquQfjGgXdB2p5Y
hxe3TZ1VZwCScOunAa/4um7rEqFARxjqAbMPH9QsYLilSgTOD2qocq4MBEL7UED+
ohSaLienwKrXgu7w2teJIj5tbx1ixL/8wrEfgRKlrCZprF9RvfbubXeJYQUU/oVZ
f2sEtme1GTn3A9QFROk6lzt/f5Omnn9LA8tr7nwjIIRIH7LP0F9fgDYT7SIXAVe0
Pf0EK/vrwM17LlTdAKDToeTWJ5myvgA2Z+cQkwrMNd3SA5RP28/PQuHH/HXXUA6y
Hvk+aOS9FROT5fgX1NiY9Tt9XOo3tfbCS6FiHpy+O0t844P2j6RFD9YundeTp4HJ
fwBcME6yosIZO/yAVOVD6SmLi0+PXE2/YQc5KI4C+LdB0vPhlihYyE6ISuEo4Vlo
tUFX54enbqmFvSRzvGNFk8q21UJ1JI4EdCfKYdeVlFaLThBVOH7CzaOdrXifVtNB
3DTXxRhkpgtn+x7wbQXjiVqIb/qNNtee6dHG2wazr5VWE02DL5zWI2PKS9vrCr8R
sV+8ue56Ze/ykxBHYL7ENBLWATQgMtGK5DLcA1A+sY0y1VyuotsKSnCa7gKRv9KZ
lzozj/EBoNAdgQ/kCrDes0IIQoOymNtWOMeEJ6o/xp99eWuT8V7erhKOuEOXH50p
Uo/+DLjfjx8CPYC7e1eTrGYymx+PiU6Q05REg9a+HOVMR0FLzeHGwn14qm10pqoX
lfp1DeguSQgxMeBAWxylNArRTO1ZUhsbKOZjJT4ZIPmvG6+aY5ybb0N10nEpjAVN
q4Q/xz9FTf34Uj9X4rSzY53n0Zvb1UrKaqg3RbLRjtGIMxSSD3hU1lmiLWnBUb43
av4AVJn/Cejbw/F7kwjtJUtXqpp8YEonjLq1Es2wqBpUKDZm1TmeYneelgRfeKzd
dHajjFrkWr5vbw72hFif2qa1ZoEkzDEai3Rx++IwTREwP8yOqSJS+XmXsnglcMdX
7phTHcZwd1TnDPqi8LGssqRXE34nnjaLD5zu5k+vLME7PFe0mkmnkSVFzfzH0YWt
N/ayXnuQInUT2LX+DcXWWUXzFaCAiKd1B8+DRoro4IRFw4pfJhRdkz49+45vGJwl
RFUj+jJUKVYfbAE4b0sD92Xagh0pFtjD1mU3qnWypMhaMN1paloMN7I6/k8c/Vzd
mN2HVaMXfbDVSWsPznE69X/ry3Mkm1ARq0FN9IgHMgF3BibeSytBq7yzxpe3pRMT
+3c/3Ec84v9zd/rs4Ovnizq1VL/zwjbSiQhgWx+Kc4a280KiOiQfpn6OKa1DjO/w
wpFzlgdccIBfLZgiMKZIUYD5yqQfH/DdiQSuogxpoJu0ltUXU9pDuIiKLkaINo7j
g2avFQHSAeJYCZEI/01Xf8zZTrqIKgVw1Cz45A7RkWIR4xPBz/ov852qNdWIRoIn
tL4j1QGf0i4r6vcZedPpk5rcYRSzYrvhUDQo3aHmrHmqECcNph7xc7H8xL6L2Voz
j9bqAymrcFI/q5LPfycptOcKeooEOXdNb4yvPdVkXxh5ZD6Qk7sMY9baNfofpRri
P/Odo7HlWOHAyEuZAi3EAu1Pwk1Iq40F3/vqf0fpp5O7mPvk0shNYaGU4d1giRa/
3pzacPa2VhgkLrtFDSywHSYuN2uEKoV4Mu0NCW5qXLhQRHOgnLmI3ympBC0Xo6ff
8azQ55IuAHiHWEjwWXNbMQYZ0lnyiwktIIDSPKo5NSB88zEhXENoXJeAw4r+3Zku
IFk6JpdjhwjKELOOb34vjdKtKcmn85lcf5iIo4dYU2+jjSvh1Y3iA9p1f5v2D4Hl
RiQvhyV078HCOrU9F0r6sSKNWaZ1dN4p3gZ1+JfsHGHSbYsKSc5DWrdUGDvHYSN5
fxBtV3OXzfktQ3MBUlXEIWCT9C8RNNhlo5l5BAKNypaQH9AmasEQ5SYNS5mFID+y
OCQ88dICR+ZoQVjaXdMuMnP4Y+bgN9nZef8ScgIl9bZn3oXES/2DDnbED47ZccnM
Zt5Q3vJEdzWkAgVomrFm6qJhh+cVqVZS2Jvg1cNGXggaK3yOhYJypJhNB7MmoPRe
dgsifEYlbTAVEqrPLvUlIDG1LudYL1uLoNTezDIZCDgMYHmdAich1LmdwZLYJ0N+
xiW4uAU3RpODT9myc0qBLIMFexuH1cxwyHXbM76FlI43gWEbOYARJt0wk0qd1nof
LeoKOSgBlEhYU6h9xW6CNq0hQsDXIEf9M0X92mSNmw+7xhZRlLeXkiR+uAqsIfBd
sZkS2mNvLOS9FKqziR7t1YKvSX2Nwoa96xiE0lrVgJdkioqShVk8CrgKaqJ9/SnP
2SwQ3I3F+oanAFFeSaad2H9q/sx4fbyGH8q5NgbmVmnUMDovc1vQ2Umfj+2f1qjP
FHZkCnP9CcuslHDCjropWe263t7LyymQr0COUgqIVup4DhyPKP/NQhiS4aGrUusu
NVujAjlgHnIX5UIYkseYVuDux6xDxA8QLzCOKw+L5/yrFGugmjgszUBDYPfQSrWF
X8t6XF7l4WrPFgJlzfqEaXpj7wO0+DRmfCghiDnhrnCqzRmfXdp2YwDiWepQLWXk
tcRhsnTeNqLeW82y6c77U4kkNFco+Vy3iIhuBRxs4gRmA4WXh0NXs2LSbA7B6Jty
ct5x3tetYMDevgtVKqgxMHWeRlJ3/4lSO7J48ssAwdbqDHwn0JYPHbDa5fSqKSRu
vWcyC13BCpPhoH+iAEZdOxTOlru6c4A6ngjIupl3o2HlbhpCbqQofZc6GYpwBiFB
VlQ+KYBjQJk+llYZiCA9HcTyQS4LgeTAppT27+rJ4uUCvSPA2XTBLk7NIbhwL0CO
V2bG775lJbPTLT7S/9MGM84oUdI9HVEbO0fzZYO9sjgyRoX4WTVJt6Z9bV+nt7pj
dvDfq/Hs99WlsphEreiw4vXFuDS2KbTcIU2c1SHGX7slsUtYrJmEl90bAVBBErr3
TqqJp2oObPj8Gg/4KjyVaamPt7+nEfqFjp1VF9IzfJEcFrIY8ehT1OwHYHGx640O
iJT97oiiUc/hllLCiTEoQiKbnzxzBDxh/X3ziLkjIM0DKQVZ2MH8VORcNbCjG5MX
AERelb9/OPG/uXeuwjY9bjTEAE1sJ/2bg5OsIx2Ek6XFKALpwPDd21Ir/Zc7y/1c
nw+ifSm8vYYL33mK5yMBBd0KEDMiECOAPFyOIemaT4p9g4HOS4wNpMD8Q5WjGZON
XcAfM0SlvN+aL0jd8FdrhbK8aQHskh7hP+X4QAajRxvkCcvm41sxPLGrq57WrKpD
kn/kzaRoHcYLaBDn0/jS9nAd4qGrD9WK/uPCEhJKGaswUb2OXGI8qfagxD/Tlnlg
2NERUd+Ubr0yrCVUgKWhLnjVWCOkUZfYp5lDWxWoUj6oTgIbA3fvxc7jVwp/bIWX
AJKyHwFuZudeWjq73sCV/9hBJwKJ1UE4eu5qZJKTpyb4fkK3CLx180x4q83q+qs3
QgpSxessrWYlnYxJSJSqtGTUAHkq4EhWYBRJOCpwNrud5xTOGlp9IJWw3CDUKMKY
b7EpXhQGCenY3opJ4R0bqapGqjWbONY18U3pEvSSojKdf9vuMMHEZV2nVhsYrhTj
QZXyBxs+xEr7oreoD7rhDpTFWieTujeWGx1UR3WN5Vhn8nyP9ntGLT7dv2f+82Sy
2xXXEQHdIdSB3AIbi6UyKcJs1uQ22oy/ByKpTEdf/7sAQtcv3GE1VNkDibrWb6+q
x4/02jukpCvhUuJ3bpefYsDfh6KcrXYiSW61QvUI9/f6ooHdeek+Kblr0KNme8z5
hXvswmZB6oqhaDURCLJAzR7HVOdhC5CN8P2sg6yvOjH8vpHY3HP4ARsLWYZ1Cx1D
m7ZWNwLCrA4qaTrIg5ul4OVzx6gHt72Qk2DieTkThWWelITmUtDmR8UAg3A1Bmm1
zdrEd78EESKWsPO6LHvVHE/aiLUIpz69sJ2sAqZSrn6M1Rs6BAwylQ59+RwmPguf
iIbnp8iwmMUiB6CqvQ1jlD5qNaDhSDipmBLHxGrH13gt3yLWI9o30bsAhHyf7YiF
ZmtnVUPpM6NfK/PdO2IZVBhvk8cu1d54EOhOg8N3UM30YSOIVTKt7sXER3WQ59K5
5TlOaKy+FY+N4A2Dq4d0d0+l5MR4DOXgq//RS+ZgN+hXYsuEowkxjaDZKOUNEkOx
oaN4tmAjG6xWfB12mdZCa7TWVntYmDAKettkdd6YP2ighol/2T5W4VXipPb2duNi
6JUQ7fJfHBqndvB5fDGWPCJOdCN73nbU9kcJ4BU7mkS+1IHRmRdeb7C7SbNFoufw
Vzx7xyHyBlUyTfldku44M8c6+LVp/kuNHDrpWGuOBDLZ5/S/IH985mVgWK6nky+M
lI8TPC7lURMl8ZwfmBdmN0AEOXjM5HHKEXN74agdh2GjZdSQJ8urE+O11nTNeaWl
fbOF8P/HWckbcd5w4RJVxL7Wia8MQxqD+PcdaVteILpD+sq2uWJMlGBxT4E5+Yi5
9SyE9PvkGdv7o70GmN0YZJffY+MuftuJJnkbMJM/PqUWhcjLnYfeLNAVmhVfKUj4
m3fz4kBFuvb/YrpqSIDlNsGy6nF5el+1n6u8t2m0ItbKfj+/mArJzGrs8LU807r3
c7ejOKgqB3HYejNmZRyYuSf/ifgt/eyp7L9CFdrfMHOAXBhX3lxIUQzUD3ZxEnMF
2UrzSOY5HPl/eMdwz1Dke6c8tGKv61wbYOBkf3kOK5r5n4NhKhcVOUaXgvIMzNTi
0GDeBYelL50F3F6VTwnovO+6/HM4JQBcTdEr2rqG/PCHYu5ehUw+ypAfmP4+BZVO
hxAD7tRXLVGdSrNzoFuqWxjScLcE4uG4eaO4VXkLrV72+AQ3p/OKc4AaUbiN6SYm
bUIEmRYrg9fbqMzju7VT4SHqvDc+7KmagA3pf1ySVfzY1/eLe7znPsVV8BpjtUv5
Rh0PdlMCFa4MB+14dgHKmMToA5O2sfTOkfa+Vpv8vzO2DW0wdVTKqoFFY9BNtEaE
bslmdNT5GmRqCCM83XC80mbL30V9W7G/1jcpmbphDvM19+76ey0xBeLf7Z+dVFA9
WUZFrHx/bBH1zMydpbSEFXye1/6Udir7ANm4WKsk3jU9fkX2TiKrYU1ieYHQM+zu
y/ky+nHFsqkcOEyLUZN68Kk6PgTG4etfBhJSlGU73jeYR9WrruqGcnrDR4p/Hy8l
PLVa/HXrSz1lxou5kDEXhU46om0qwQmuz0smmyDPeSNd84g8hV0dt6eZyjRqBTbe
maQ4sm6CO1/5DIASJuaus/RUBd1NcA7qiWEaZm9/g7mYrdc9nzUM6Do/pK9q295K
FYzEXloUtJH0ug1S5DqHVTanCjzu5SrZQC1RNqmikwhtd9GdQqCYeGKJdJFTj1JO
fhAIxR1rPcwg+9eaJy7+AQS/iMcyqQipDnm+erO5lVf6PWW1qPXVeAwIgL20GXPM
W0p6KKuqOVHfZSeU1QsTSe2MDnuRySCUTH6kuTVkbtgX8i6mlyBya/C37Ko3+qkt
nNrNHiI2zD3n2iAUkXMq4ZbM9FvQpdjJSfXjvLRE2eql6wnsFk35wXrDJ3sFkKg8
/3DiGLfodtFTLtvMr0XXeNqNdS54DWzwlvgbTzfxAZ7xpRG5M0YGudTygB3U+Xyh
Sw5UqJ938Qevxdc/IXBgjrL+NNNNup1Jx6GBdRu8fxgo1r0lOvea8iXl6npnb7JX
+hS48IFOC2foJuAmEC9GrAFClxgWMDTgTaamN4tIA0zLY9unOlhf1dWiK/TIiNhH
DGrHAmO3WmGqydf4+8P9u0gcHj1haw24ABkUETSKUwVhx19nqbgBf+BvEVa/2koK
9GAcPLfQ1/IezhJtxbQAytJ6j0DZHIercXAc7/V0apY5cxNapugyFpyB3MKt+UdO
BEA+PCm3ugz29oH4vjCEBf2QRqt/RUHrPoijMI9LqV5+h7J7uYr0qV2YHMKCRKxF
KR23ZLpi576s5a+EI5EcQRhv1wNJ9UFuVOHeTodtfcWwcxzXYkA81Fw/qPV7JQ4F
MtyNnJQeybIGQ99+yMSWCBgiRZyWFSv5H08QPK2iNyocDB21NU4fkUDxaAxigTTm
EM+zmy//hxugau3ma/Si0rj/IPop/BPKVsbuiwJIPU18y63PyoWeJEHBJ65OEsHF
TuW5q+BOO5NrZYhCO/Snzt9SvlCXcgvLcQfMndz40nL2mNZWODjwqnFwSI5rX5JZ
qlpfnveT3ZjRmmgUAok4ttEzn/ldRcDGS2VK8JUYp7wlTgPNzBVg0kLwHzD7pVAo
xdvM4giMB4wHBRIAWjTX9mPG20x7N0u5KKfSepJ3p61GwECTccDFtjP+Cu0XMh0A
bl/iAbHBsG4hS6r0lDQmbWPAr5s4XSYQMiG67Lf8+/Spp95DZdX3ArIDEnY7/y8p
bmtalfeI92/G4bCx1xTmSvhQA6tsr+q2jbQy08+c1RVlwTUVg+ldKMcOpuj/U5kw
myB24bKX+Ir6IyJei8RutrqNZVM9BvOzwX0Cj0b5hdvX3zba+HG/p7mr3+M2kwkb
CMdBhJ+pbBvQ0Usob92UnfCoU8zDTbengS+Km9xlmalOIuLPYI1fa1I473IpweL6
+IhULIc4Z2Kp/fwwPY+prTxvE6Gn21n2L1Be8D3bAKK4qShYIcjA/6KwrS18fR94
0p1nZ39p0wPdqVGAOavhhxcnNonDisiUeo/ljoACWHFytI8049Qpi02FVYla/VkV
FeIzHSiPHbQ9c9699WO9BT8CrCLBg5CtXEEO1GiH7AQ1HydvPzr7OyGEhOkT999Z
xAgKCSRzzwRsQJ6ReoQjTQXiBPO/dSCBKuVfHCn4r0SHe0e29Q0fnwflMC4nuNpw
aRMGiqXap4A2AYo5c3bmLcHKQnLsdw6A1uSOsYOsM2vEn3r6Fkk/FPOTmK4oBXei
cSdiAX3df0Bv7otp+DUmWdFgNH28/KtJJ3t7EYNG4qz5nIMEGvLwipvy8Kw/HlFf
atfDQzCTO3f1P1Vtp0DikJDMUxWFaq6mTz4fwJ0Ka9+bTeAAF+J6ECbOF2jc9xBy
/eXp26oFf6D6itXMyVVH2b7+gHQ3lqzNuvJyaZxuDHG49nh1ghjZfNbf2FAZJj6v
srTUzpmBO5LxHsH7GkO0/NRm3vYemkEFqxrgGgQ4Up0xTIjwY1Z6PQtQli1ljGEV
nXMbGxIHroc0koIQCu5aezJ8frMc4qgbmYySR/G8myH4zloI4M3z002mgGy5HdUt
Jnivv24/FVPxDWY1FhPrmWiWgK8+H3Nc44LtDWvL+GV6V/3mI9eQaXWRzIVpxmhK
GV0BNjHN34AuEGiL0Prox58lr6TKdsU7vAn5UDh2znRiguk1bYoXlW1tq/KttsMr
Qgkh+UqzBeIbzRlxjTZlqPLLkU9AWzfsHSx2iZug5Wx6wLznWnf+cy5VQxTmGKfm
sOxHB1dQ8X6DYALpkM81RAhMF1kke/Ix4UY7vdNaxr7gnD1PUr9S+4ux8cvFhRKk
77e4xQExv3/MULOeLTPrqeZH4P/9AaLx7DTPqUepfZAtjuI1XgSh63kUjRGyAwuF
Ka5RjqQJV9zkNfNerM/8tuLrOcyuOMtwM57AY+q6hxn5VfGTVJ7OfsjodHGGAxRb
j1bFaYtYf3ZbowI2znpGNhIMcC59ksJqaV21yu6W97ekfC693+MdVoFomhU1UaYw
8BAAhc1Bw2N/zV/5X3kgLOV6Sm6HW8GiSBxHH8410L5mV0OAXsHNlsfBaKEwD/HY
m0YpEGkajO7bvSljOUiWsJDYiGewsCNKqIoCdrhyAn8s/VAwZMqlIdCaL8YWf/rj
KUvrX9ttavMFsz6A0gnoYXtCHVzm3EySotXCl2+hmDflwzI7tXT7G/RQIajayRN6
4UqXXo+WwhN+ZkX4o6OGzJB8UTDs7HaT7GFzYESxDinEKQjyms3M0X0LXeK2YFh3
spm3pJcn90GhvhJEt29/7HKcWVrErJWC705XHOhXSG476FsXBOWP8fGSOl7bvxL8
+kQ+1alGEJCbNhPZpvKNe9xRBuxJor2OwRM6JfvDRGbmg4txhwjBN2ocweFQcqFS
WhtT82UV0mdhdAf4zloCj2J9fSo7/RckaGlNGcpCUUcy7q5Bxdpjcnl85hsgX3/i
Xgn+O5PE6Kt+omcuuZPgBApVVkkGJ6d47f5slrduzqcrRXOO60nAUjQFevvhMX8+
RmbZWeitcTkyiyVxiMdHTDrf5jQHRlip3dY4XGGrN8ijY8j8R7C93d/lMuUqPo1r
u2Ux0YQWBmIqLBwlc8AMLVfrrS+0b/WPYNVZnq5DQbRdDPSL6PR17a9LIrPJEEO0
PqV+Zrwlvh9kK2bNerFKCMauMvXMEdzLdrC7XC5ACoYMrNGZ5PC3V17SwkpXsZiq
0yp45BU+usTv6QL5+ODVldUrFZfsTw0Dc/IfYLHoenXDs95GMjsJM15qaqowMH/r
N+wcEOnoBj9mdApTJzs7aUF/eiM5j+/Vhzqd+BgpGwq4erjSjXgiJXf+6kFB+Vhh
1c4RF/nfPPPWQuxAqCjvy2qmoBh1KfFX5HBuwfbFZ1TfPwqw5LgKVj7XDZCcy4i0
s+6QVrFUna94NuJUbb6muVmJ9KI95xeJRS/PRBeaCENWLSoLjcIBkfqaFgpI675r
k5wXe3/alNHYyl440cKSngeBrzoTtfSEUB9UsKZDKo2Q7iiWWUlWq2naJgnAg+cs
PAHjY5shlYqAPBPjL9SAtJbcI7IHKJxE8NhuQdep4SKekt+zX4ac+BUxjptSwrUM
He//xx4xFKrvKEPWwiQ1ocgrHhL1xUAJr5b/hdNknC3h7SbPImb1b+FYq1hl1oie
cmQKRad2ywZGQBeCS1xhrrW8V8l252AqnzmWLoKo2B2CjnRo8KgXTmLG3WMgOdA1
iAwxppIjE/VGQ1kp+xYoTscd/0mpTAsvu+hZtyFp02/neOp9z/yfNaXtXYrIZaJj
CLJ9UrwD2GS12WPdq7agl6TvtCC34oVLhDK5PxggO0t2+JRn8jNAA7xka7HmFmCh
rk2Z1wLtywUTbwudu/S1ab039aD56Wcvtn6eN4K8cf8X/I0tBIDkm7viFS1suysF
oJbwIrZ4yWuWyjbITZERSjoHp9+ClaatM+iODm9te/mRl9cpVPArH6GxYIqu53uG
y8DEODqGeOPHexw2u7ferFj94hlZmBvR8iicc3ugS6liiOFrE+cIZz962nC435Nj
hYXxbcWbAwNpbAloMY5TV5s6qOJViMYYOqhD44FZB2cFc55Ro/vhXcDlxWKyI97P
r1ySRgZBvFNo1ps5z03WSPU/6CgoN9uJWxikEvYhSF78oTYd8Swp0WhulA0G/bUQ
Rusvkgmkk4IsP1HYRoVc5EOm62Avy7yn0ykNDDad0WaM9GLFhhvne+LLPCyO+XEL
4dSEvPl72ywco9AVvivA4Znz8e9Y0ZmIPSvVMArWNvgKkg0GOul4nlG24+YPKKE8
jc2+lU5q5lee2IMydCCmsCVie1yc1H6KbSDH10mn45B9MO7H0rbJxqaP/xktlnoi
sBdg5OLotDKDhaqMZFJPId+AzvoLHSRm7yPh13L0nru5Zlj1GFkZWExP9Gh1lwwa
5dJWgR3WPNqqXKzt81bAyCo5dcvIe9pir2pdbsO0+DjEsOuTKC5Kgqk9J++xATVE
JZ+vumAACA+m//nENsI16BBL17TBTOr+Q6KUUthT9ZTmzTF18auZVf17JBA1L5aD
USJRWfLMnI2AzYmFsnhum2CGI/EwOBqD1GxfWoCUzhreAruPC/WIU+G2wEUqRb8T
jSMJJLr0brm9B1LwElyiEBWlSLxmn3RKgiqoLdQGzCO1eosZW01Y+VucZGz62lpw
o3iHN7/02iYm00BtN7iNF8xSI5UGGRplduxRRw2zxdT9QWKlCpQSe7jvxpGh74bn
gT0V4itEnCYRXVJ+hhCm+KUCn8xDH/rzd9h/XgTnmCHYZgj7mIwKCMVHCTDbLS07
NUMQbhC9NA5V2q281F6e/tLx29m6hbelh7ESoN5sB5zzfQ3bHtXFjBJE7MdeZH5l
gU41aZanUzxpZ1kCyCOon6zc2dTVFBqagcO2MKh4l9qrnMuugZ+bqTt0rlpJXHg3
Ji3TlbOoRUcEuF55FXUbmXdtxM/WIIlfms8c8ypHBOtwczTQV6GjGvYne+vv0w1Q
ouA3cHcvmYr6my24yNmnNigxmLkgaOf2V3ZXnf2NkJUdkU9drj/TfSQDpgVqqy1s
ivQQY1bH9WrV0fwK/idsJS9nothAeiXAqYAmjqbJS04TqiLehibB5WhdaPImSK+N
njrOmXzKYXbB20ipNwbqVVUt/l4yKQigiE1q7eGKxZmHg0Jcd/cAUIT3UBCk9UmS
8nqdDKotk8FRW1D5nqYpcktBAmrT+cALPQzIufCv0RnrlqQ7FbqqegaZuWsKKnVB
Q0Q6iTYwrvwyVZYTNcZ07mwpYFTLJ+/KgSkAgq8s/N4p2Moa045MkfhPbX3MD9mH
jeI5XMnavSnR/y902CTdONs80ao/FQRe2z80pqDIhkEipY2CXcZ2rZbxkscOnX1q
Evr7c9suqoKbx54krEc9mQufl0PwikgGoqPYPyFwi7LNT6YH3hKCcXC3+KK/Gxqs
fJNIXWv6tBjtPYWHGax+N3SfS/5bGkwSoZuMc28yYjFcOZ4ilwPsU4Ej9/UrQCqQ
ilh92dtFS1XJZs/UTL3U+9/nLT+UahaSVVCrEf1gNCDc0lT+9OoiD/F7huX02zlL
3ZJLwQlfAoHu7GYdNaa6JpJV2KBRSJnylLZVM8Fll/VvhBgGEdSvh7vONEuKpfW3
gHiI5/l0Dx6cl9tZNtPc5Gmuoo6xKiBgn8eMgFM8DwgNuKd4zdudywHMpMvvTBR/
2jWnLGLFdcHEuWS13a7p0toHDgBwC5rrlgx5P1lCl1VL3hJHq9M/ijeEjXlZ+Sqp
tLCkcjt4VdWqROdYcGBEsMFny+YCd3pebXtqumEHP+V16oXg3CXftiYtsqW6BDDu
3zJprNF+Qs/RTO0oOTykyPHSnY7Aae2VG3TIJvcZWqqlZ05jUp7JeFP2SH05qa1H
FkVe5Fn6bW5BaR+gPITNv9MQaAmcv0WIQ1IGMdBRgqB4FrBrPQjRjAwcTC1XURH1
lnSzoiyvy+Na3pVDzEHJrXtVRYP8mAUTSstDhRMswVXlD6K5egA1SKcCO0pSktd5
rEsD1cG6lkpslKN7aHVDInvm1S3vWsIczUr/qQ96hYJTJXLH0XqKN14SpE58QIq4
ymEizuyjYffu2AF14H+xMyrvf5+pGr6XoVBjaeMc3t81gPk4H6xdcREvsZcQwW5s
E8WuRBNuzMQ/5FqkBD1DYqXAVkuniAtOt1QGeGYX19vG5/y+dTUn2K5jaJ9GBGUX
zxw+yrUOojgfiiQIz3dmfw2vdRFjUWB+shbLvbso3uHngmzoyiT8aKqq4WdJ0PV1
fbdnTTa4vv1Ui9cHulE00rbZ2kAQlXLDpihzhaNY1xizUl3IWOVsrgEsrh+pIbvi
Ww4dW6Hwi+3ebK3uUsASE/IaZsbMkdVV7l5K2DDTwKz2wsgeHOSgxzICh8+shOiB
zcrJf1/M4xH8h61tyMQ+WAM+Dwg+E8SogCmtY0UPRCe9c4f61IpDAxj8EFwCdCtp
edXF344JM8ry+Q1Qm1syiUNHcrEE4EuOiLMu3HRhMg11WOKm3msam5OAaS+D+f62
rYLFllpkKqgT5FrqTK9nYloYOvSvr53wQxQI6cgjpl0i7kgO+UtDAeaYTIp72iBK
mc0Zl6prEJhCNTdJCJ+SvAbFIT0H5QiE6brVl6/V4kAlppxet2/3M9DNzYUn0We6
1J79JmL/RMEwOe57/bulF+7x7iG8O7IL069HRN07fZ8zo+meRwHgm0WgE5hV22dP
C7bQXObI/GsG8esvszQRjZvRXxefiqUydgNh+K6MSGHofIXZ7iPDCHpDnjcDNk/B
vWExEEJ8IaTi7piAWCX8HQhY/dXjWMp6nvpDWqNY86vhetvuYmNkPE2TNI0GuaRv
/01eY8ZJYTV+J+qLmF35z9+4R69P7Bn0Eqkcko96VuDorP71igcN7hWULZ5cR114
X3C9/xrVhsQ/J9hswVaX1z65cBy/rBL4nFz1IZ9oZ0QgQAfoqHD+/uJ4CX5sw7Pm
viw2WujgX0ThZue7ixmgyrK+D9w9FPgs90xEqVI/25RJn8cQuM+c24iKC/CT+guT
SN7G+c8hEzaYKkOLwWVmz6AP78bMoQR0RQGtgx0SugxOyqqf4nXNQEcO6n1PmYux
wjhD9uLyVgviMN9Oi7ElIuJI6Oir87l3tvrTYLkMmhWoFco/DLT6YpW+vLzOXGop
mC7Ne7soVy8kf/YlaXSPYQRb/w8gqfelK3v7BJPcZkpqwriO47KmF/VYDSm9AeLM
cnBdLAtiEozhwDj6dPkDwgJklqghVGBrs0VYBUvm+HNmDY9A7JPF67EYbMigXnNB
PXxbbrxoeb0G0vZ+E673UoObDfkWzp/rV9m+T0AXoRASUYBTo4AtGFVV4fCSW+w7
pExAEllu59s9Zhy+IeylNsY2QSU7qJReXPwjQvQ5GJy5KfExnEB12BgLvSWoPd+Y
gM58JNR9x5lztceL5B155RIxL7yQA8ba+aNXXFk3s28QlrLdsqJ6uA/1fDEeO11X
dYNxp+ybNc0SGNSvobToffVhQiEl8ySXnGmzHZq5fpirQCl2gD7OqfSM5g3WuoqD
K1iANHtNyZ1oNPpUpvBu+SwnLYPtYOBX3JEG6nEDnOo5w1impKcGEcpe7UHb7ZG/
9bEkpWoQvKMygg46yZ+BcI2nIjXwWEfloTEdzKTax9egfRG+uXQRD9olZjgMyOWe
kBz5/SMZ/CrWee1UY7o4sQaGgsqGcXJ2yPfQBHUQ45NVE11jwm9b5bHBMgsXjwqN
Q4dVeD2ArUnHJ2//pp1eI9LdvTAdUN6fs4Hd8SsExlanc0sNvED325kL0sY7nndN
kWnJYs6vTY6ArQIFdLIZA2RmuAR2UdsgR4O8yELWcpeqfjRSp1xcof/lhc4T6m/a
bt7IS+JXReYYMsgbOwwohNTqkijmbaSYfidMKkXspn0Atu0tAlf5tz+xgvG/qE3U
CXUE1sBey7/7vfL9LeEH6COO6u+vHktug7dj3otDHl619vXdUVEkfupy6+SfPcuc
6Sb5fAL7OjesW5kycQ1seFvlfX8v0u4/rwz35KoPkPlsrJiTwydjZKCSYIqrIFSj
5de92DuIBFwG8p154GLJ3N/q/lz99hjbfCzWXxBuMWbuxA6jI41tvcS64jBTDNlU
UaUpDKfXbrXptR+lypq6ceBd8oiCGBOI7v8q83qXP1q4MoI2PKZD1y3pz/MincbO
EiVFnaXFL90x4f3wo2EzveObbCSdVhyvPDo5AzrheVna92CMOoXb2MG0SKyepmCE
r6b3EY1QUZke2XB+ACaLDGR9e7Zl6EYMRqNXat5R3KQl4ZlStmZ5P9s8pLFUp1Y5
YVygUoZzC7hYHRKjl+u2AyOtFovsukR5NWfX0d7upkOyDNjnyCDSwlLL6m1gep4e
jk8iCkSZeoXs2gtiBEBwRXjV/6ueoN8coNCGr+Z3u64nQIFzqh/agLfdRUJMZ+Fz
4LKkv1Wh7svCgm+fPR9qU1Y9fP8XBgEqLfp2Pl/4e0nBhRyzpO4hi3SM5bKrtB1V
Ksxdmv+IixhwTMow9t7ZluHGQbQLRCnybHyzrFwu3ikZG0/z4XixFFNCre+HhtXB
eUogMsle5XkNcbCcCJP8VZLViQXc85Fj1JgE28ECJgIAPh0pFUO0EmkzBVOHmRYZ
8D6xS3hPF6oVGHilcwP5ETnDhrc2Z4G0SraOxddq7YVhPhQHGudvhhMe8gLcRGyb
5BU9C8gbPVzUt2eLNXC1OatSev+j+igfZbkxigl0rpT9jnyDM+M7va/BNJev0KGD
+bpFzesJPZcx60zDdmYmXIXiDfKmwJdDCBQ9M53gNmUBxbllYWPaxLvSsCyuCX4W
ugVMsjlejFDCn9QQnwl9LNuXWRCjJzPvUBW+/bIdy5tkIvFeYOoTQyaV/4assqDb
PoMJvwaRkJ10ipJXx6g4TLzG4EbOR/sILCAlb8tlKhPjRE+7yjO+vM9MTyS3CR/d
XTg8Medqx859KvxNVCOJ0WqeirVOb6Pyd4MaBsxHZcXiXvSpzqVWPV9sX8P1mRUo
x6jTi/YLpt+QlOhywiV8vnqsna+sit9B5Q5j3o4B8NEZe+5qomijl8HlMLnC6+Ik
gl3uZEnKPAg/WCOvYVA9ORc6mHESwVsYLuBeJyVsIVivONhjOzNBCcXE4xnuS5mb
V/Utp+dhUkDxWwzOUR7dl6Ta5HG4+3AeD7GuenZnJVZ7iDViqS+4GCSYOMDB+w5F
I3PRuGf6IHZnDXxQcQkeJL7r58tBbP9meXMLzv/7kynifF5tTcGXYX3Lhlv4HuNh
b6JsK82L1+ddjD/r7QSH5OmfgiNCsv4WkxrnxqAA+H1oB4Ot+n1FfX18nqiXT1/B
9/Fy3sxn3wBbTsGF3YklvVLld5l+z664z/iA16hd+fc/AgR9B8JVV3ytfp3wYdU1
mB/8H7FZd8wMgXSPLD+3ovzWFSoBXMf8FXgNA0xsayLQnjjbetHvg73M+oiTWn2a
gMuVCnDc3KA4D+SbIMuCXyfbHTVHrjfvjdLbIXOPS9nGutp0X3k4G/XFKF0i3X0x
I4GkwYAP0UX2sajZQKvF3sveBu26vZEL3or8PyQ18b3yOdpk9dHDOuHny/OWS1Gi
mQFxN4ToUq4ijhm48u8aCQpdK39g7yjF51BvBXlY98rHeD719M3QvtZWpVKb+/D0
B0iaHOI/nWlA4KPlmQeWyjM9gEkzCAeRJHSSPUuvW+hawPydOzaHf/7soCUOc5jh
Hyn1KNd1FpU1gy/prb40E/le3RdnVWkBbjjUfjinPwiZuC3g6XaRRLqyCIeDyjeZ
FKmMsLF/55TYP62SRA9RcZH+JfVIuRKEVUcKj9RKb2BvjTdJ0t3ZNjDnEji3fIO8
qIhFMISbclbD2IaE1aHG5uyYerJzVglmiDyQby5inzkf20+8AWGqB6RdJx7YS0AB
kqOqNIdCBm6FuMZzJYZpVusDc5fARPYRZI07c9pqll+CQorU6h/UkUrAnEkGBu3v
/EFljk/X33CPr230edfddNLuXbF8UAN8NFzz9KztCojvHC5apQk6UsFCvwNulXSU
cbwfFbH8hChank0Nqc06sn6fj7/6OLrz8CODsGJenOYc3f4r6DIuuAYd+5gj1OIu
V+Fd2tDLGOLCmQtA47JzOth2k4R4PbPdmNavbD6IU0YTSGuofL5bhSu4IflZSOhi
2KxB0hq7oAnefYw0QYOywTg5tv31Yzh0xPKQmQORO4xr/lywA+nLEa1p3ZYmjHJc
fPZ6Tpw9nbrNHJ6HDotmTW2euEbyJHvm5ZcYC4hYx8TZQq6GNCQIJHI6WABt1j1T
j95oQmtRvKv3SPdyXcgnaW6ZLL2U6Nu9s2xxmCYl3cJ5BS6bs3Nfi2AX5uts/j3H
YQ0EhjDE4XT193Hk4i51eJ7irXjkdZeBpZkAFumnnrOLovDX0DUzWQe6pR+6Xf8m
FSoxubNC9cnCxkH+kbFzs9ZdY0mLhF3p3NX0P7BbXmcH77IKqeB7xiCQWsOGNSa4
qMdr0QM7NtJ5/0XFRctKiKLbmBcs3ZPWBalA3p1xFCB0GUf6znRnNUroOyq9AsEr
4MlitCOqEX0dLW5yWYfg1C/xdScShqy3iBC88PTYa8md6zIjHTgqd3L9WNk1s/cO
NzV/w5T4lpvKbPz0DxLlhDrIdiMkryvRBfUjgTPl3K2uLlJUxVSl7nvbJSAiUh1y
FI/ZrEqUqlrO0YK03O+sJOqCJsXz5MXwlDPtR00E6bgnd8nmEfLH3sHsM4HoTOq/
LwgHZstB1wKm7hMQSThzCgJc79eLF9GS2ROjRDBADfei51r9cxgk9m7rIh1WRH+P
dAXRGPDBeFMqJQGz3zB7pxRTKxTcBixFDFGI0UGda1NvhbrII2IrrpnAK8Bha0fa
wWe/WqgSXUG8UGGnl9UeZL9ZLIPrK1g6ytWQsAyhWes8jFuHyrv+dbSnh8RQMwY0
pHyrUbrGCZ7ydTkDGDiIdzINnKKUR9bTUo/zoBtL17Pl3CuZm+vD4shq/rLJ31UN
rFyEgE7rzJJqDUEMrd2hOgcHbgG/vOy20w2I8isvz2KTVDQO4xi21XWDiPezpZ2X
X6XJowCjFbTJqFJtHhl+dLL+CvgywGWyypVe5ZoKGc1DvXXfkVvhG4hvn4ulo9jW
OQK1jg6uJNVrJ+9SU6dUOP/4iYcRzokOhUP9wwxA2d5Spls4U7iNvp0MnSG20OoS
Ln9dxso+OJZgPyC5WKrIUvDsbppvkRmtafaYjAQxLuZEugUAzjFD2ti9/y6eMHv+
cv7Td6p1WBrNSKCrKGYTYwLZsAf1z8H1WaAry12qVdGihj6SuJyqT57V+lRDyqV3
hHhFSJeAOPZBANX7nxPbyQbrfUvnSLmiW+tcC4Czy/vDgEnu5lPXjOebwetW2L9k
06BOyEqR38xS2sY5MCOoW+FeSzuSOt1KqRHlpWS2fOCx2U84XXb+5+esQSLSi3CS
I3vglmErWgh0YwmkEwRv8aRKI5alXKAVs1FWpoHhBkB2lfXq9Dx7MEAj6Kk9DiNq
ZPZAv7awn5d25F83gp2gT7Gv2fGKUt9O8q4RFnEpmDFv50ha0MOHqlDx60/pair5
yAMzCp+LW0oMTCGGi/VuWwyt3JGjzW4UFgc1heMhjRl4rT/uj2yxjNccVKxBcTXD
DiUO79C+J38tPbis+/yQb41bBcDIWMelml4SW50jvorude+3Wc1L82Pr+Kn36RSP
N6HhnV5M96QCJa7DyCzT2WNlE/UCf9Y21/ZXRMVvn1/CCd+iuucafJUI4NU3rExk
UczNQZbk1nmxLPz6MC7jWgVW7yuT4dNPnK7OcGBUfrAyz+Ayy3gPakv/5zCTG0Pz
yGlboP/7PjNvSajt1jMZbi2nFC2joYmWOSYBgeQL/X1aj2k0DvzFFvlCOpCzuOhM
kc1jTW4sfZnPtzFphiOe9E2Q0nkGl1hHmDVWsQbnkzdT0JMHcZt5vws4Y/ulMRtr
0YUD4sUXs1DmlN+GZAP2RK9xxksGZ+uNmmPrUPhn40LBKHaoVvSBTG8tla0BBbUA
WYvJ305Vt93RaEoOfPmIQX/OQonL4xazON3DI5sQflbEfbGkKD1rEYV4XmRap674
wnThHG1QXCUfziSKCj1+Vguo5i1noktI4gdVPhgQc75kzklldWyyDYpW1Gf/KIFO
jjigQ6hCob+yjLTbHgLjSj+Z2dOO0az/Nh0Dk5XLEk9mU+WMnU6MgAj5StXRQmIf
fWX5kzji/1d8hzOXRiyOtYsHkNGgeQCx5EU6CARCPVso4OPAAbSlV50N5ZXkWL/G
0wdPxSb47lD9uECzKqT+o3TNLpmzrebHYsERwu81+hU8hMuHIGtny4lRvLfUGXJK
7hAg9pFGsTssE3Vr7QuiXli/4okq51PWZTJiVAySTSzIygkwSTSN9H7qroAD8HtJ
W+xQvkpAcQ85/eTL1CyJy3iZ+0vCZDIc+JJdkGllRKu2pEJyBQkZNz6eyntB86ak
l7NihRHL1tLUrFztV0gHTRSQMhKgNOQMf+5jDe14FoQTrLMVCQxKYzs/wxRZtdxu
0lSu1ZpqyQdZUT4FgHMhUXg4Getsex0tHNoII7LygSMkrulQ4KKHuEGD0M+3Ridc
Q/FVxUr+iuxayxRW3q2OubcbMUY1f+rZbubPQe0UQ6y9fsQtScm4N0lfxTT/Lg0Q
yOwAIqrlixWBJpTI5Hpt2sbpyIwQ2oOCNGsdYJPmAtXY9f75JK1yTubt6VXZzRMm
A506VYiDBT8hqMTYCb7nCcKTehAOyw4mvoccsH6563GHDhwsEmd/dlB5Y2yh1XmG
kMRISAcwQxcb5uimA3d6cr6ELwCtlcrLOIySYOEByNQqTItEoj7ukIYFligprvw5
hNmK7nz2ZSj1sad/VBtRv7eYHRPg9VgrtH8foUG4aqSM4rzoqAl4pUmwzCkDhavL
amLXu8BfqA9GB8NHwHp8GPomAlBqLzYqHT9nVVdSIrmD60BZ/bBKpcqG19E+NkDW
qMK9N8xABcpK7oVC/lYADZkKEFtFkiirxn33YgnwoD0fdWIjjJj6jGwTBpFEmgFK
flgzm1NPfVuFA/CGf6g0G91XwC51qmfxpNWR7YOyK+op0AXiBhtnXukj2gNggjwt
zIdknUFT4pfP52UfvXw5bs8sJHWnc0h58idXrG1wnenHzEHn3d5hSdtdwPurnTTj
io9vcvsbPlN2Pqke3wRXoPViEtxHshDAFAOsjFoRugGCkf+XayRAuwCjSw3rvpLE
vOMmvU24Gala4A+pkXsqIw7XTuYAdNFVZ6ybFV2KqLo0jiGym2lMrOTHciSuRsM1
UzNuKwMJOmpKeNUSOUU3ZeJ6GmvZKFTHLi+K0Vr9FeHSlW3wm0xHun2z7Ka6WTiL
NJJDySBDeNfQpNw3reMWn2IfnjoxJIYCb9cNje+DCFqgqIaHi24ZYXg4YseOxQ1P
MR/AKmJ7CIDUbBloD31Vev1xWeWq1rA0n0Bf2ltGyV/VKeZiWfwsvdSgJETQFXbB
25HQKcCcSLS+yVs3wJvXkjECBw7e3jPI0jyhnHCEAdePqo7qfI8PJSltn+efqNxP
j/XXG2iZQ2mKoGgrlwHaiuIPY983EWrSXeTtHmezpbmbZ31PKNNs7PbXD3nmjcXm
NcuNRXyGHZOqYl8Eh4KOqJSGkYCIaj00y8w+ctfCEQJFJctcI0q64ILMb9I4xt3d
s0HNx7FKuq9BZe5HbCUOTZK2K9l2+hBQ5eqekpDjmWb0empEoiRP7foOMiUxR0VW
q3b/9PfbrfAnJQPWfo3vSmNZl0CipnQZn6T3SLhSZXbzt7HkfcEBbPdRMarnD7lP
kYgy5XvTTngsoWJNGDwWWYaJ9aWH8BT42BogzcMq9tZeJSBwD3VKOG7XQYyogY5X
mQFy/rDdkpWgIebikMqgy6PdizOqvpd+/rdlUb1ZSwImxA3hzTyhoZ/FM6Z1bMvV
6VEMCh8IIWrjFoX2UbQqpM54pS1BfDItnXZp/Dc9Z3ps5PRfPMomoBInp5bS/2aJ
ldNIijYm7jIeErvcgVbrAjk2M9jD/NPFtZ0YOq177XuEjFjOAsddKI+ef1h3u5bz
becHTyjYDDXjjF7P6Bv0z/7/6C7S8dgrlCPNMdSqbh4iFicyNT4RHYtnSi3np7qj
AFzXfuSRP/ntYBp7RTzyNfXbZSzluq89T4t7t7M10T1TR+evZ90gkdHg3SazcR2t
MCqYHC0I0zDcB5anxl0n9wBmU0WPi+2UezaPHVhoDYbjVJlpgJGRM6sDYjUyI0/e
cIT4MmSl0mZhBgjXLKFJ1cKKjUNa38VoHU6bkKLghT3Bj9L8UQhqLhXwP+3Qxc+L
vlLRS5Yupy1ozZOg6Zs3qhM4FoVgjY5na79IByf4wKXkMj/bRcjFaJBwjPsLV7eV
YzzdKL6g0EVWsKCFXK7ZhWY4e/OIbCbjR3eJ2raokm/RIcFUgim5nLh9hG/QZ1kj
baLLW9NVjENzc2D2r4HXEkRgTlAGqpNvtiRLl+IoDZqfLyKqF5eXqdXET3opnpIG
vS1Qptg3e3qLUpNJVEzheCmBcq+2RhxtGUEc2PyS4jDrfH10swwcs5Sdcbc+kQNO
+/XHj3/pZfnwVu/Et0K5YNVqPcKuy7aWA2VdyvPMQ45Jd78mGVBiMryIoe7kj/C6
VhPWIM4hF1wRv46uNF3GEj3zGtiHdJxTsAjCcmMCDo/kCLGThxmGEqOQtIr271Zf
qIUimUP5wVKg4bNbNN92KL/YufBQRRF3sJb7rqGuN8knlrgnEy6EZc/ZD67F1uHM
hlGKnfW8sVB/82AbWFLtYpI7lKgkYyj0miEXtHZvPmpzJmFyVxcEEMhmZc6lp+Ah
lHwlUD8e0Bi4c19AVFjeqsiibddyMKitWG4spUoaiE+vJhZ73djHYJcLkBBKLEjM
558VCOpU/GadCKyR91fnaQ/egolGh107gsOj37Sje20Ce5B7gtaysaVsORUfnaM8
IkXvUKgeKr6EtjhdjxRBUKm7IrS6sismVgh3ndIoOo+EMByv+NQ2OwJc2wlUpxe8
gtLe0pNZyvfJtyr4MM7FyVL4iQUoBzYfBhsfLz2c6I5PrJfvR1xFj+NW9VwWaXHh
tpPrkTIwD9cW7e6SwBNpYAtvHERtgxb362wrEsqgVbNN2cuvWIFDQA0VoexsyuAS
GacXdYzu4ZRLSre7O4WkmqgRZqQLvREWyw/vU4JzUehy1BpM75vFwT2RY7DMAytF
CQ0FoChunqk326+thgjuY+niPZ/bmG2w1vv5xzZ4+HXEmM5sd9RFoXC/jZ3eivcP
bSXK3dPPOkedpLxU6bMBHXU7kDzBJ79F0Vy4s6C0GqEx+gt9VJxe4oZBfQKk5t/5
kRunk6LGBnk3xu19p5bmTguHYVQbodZE3yj6RWicXfAlvFT+cC2XPvOAX3HGUCbX
cmzMtU3SdOvVQoIe1l8shN6L/rJeyLsIk5l101wTGtiFEOORq1VTYUFSBtR2M+uT
6TDfxaicqBF5241cnoBsLOBR41CKyY9L85H/I5xcSbadC6q9J+yucVurgiTTeUVc
aVDfzoBZ6J+hzGux35FkBbwTbSJ1Qky9P2un39NisXy3F1m/nWRxnSztw8iYNyoz
ebMnOdGdUa6sdKr9++3829EaMKMcSq1qkdySkFZLw/BJmzwWcKF+k6gCCRUpIx8w
UBhwxCNarb+H7wGL9FjcQAZ1jXgp3Yh5cCkRMDpOt1BXC8XQxIIndpcno/+LGZnP
aPvdgX2TRTW52CFYRyzsWdlXdWWyFlu4CzrdtI3W0PoxXiqJ/tBwf4u+6WkF3KfK
3j0VPuqEB7x6GX7HemdZCj0B1CfvTDO2BiPm4loaNnDqUjnT6XvPoMwFW91K6VA7
u9dbmYTrh2Ykee2Laj1Z2IBMEEo2cSZ916VtK/2oYsVpb0LkdKb2YVxrqcVfsjqV
ccay4S/tijwgypFlEwFcaUie+MBmMtmkCufaEu5Mh5KF5v/+RIrWSPV27Y67ngw9
yii8fcz5QChHauTcDCe2cCxj3Ghw+TOGIyZSvs/w7+4Ioo38UrXzG38ZvZ6FexKo
UYkbJAO7WJ5BBa/Xgnzvbx7ogv3dF/N8miUbPNx58cwNMm0aK69a8FGDJIlkd9Yl
gTou3D+lO1PZkTyS6SY/dCZxxCS0JvUSkJhYOugrQk3UX52Db8UU2c82Bd/p/NZb
1+ihAqoirLRXP3VluQqp4Spm5KRU4QBh/WhEBPqFmGlHT7Ln7hgecJXK3OOzGCs1
HhdlyS39wZmfW83135IuwHBfZhXUAK+9b429ZSsQDy2q0ldR/ecYEMljIgcrtIjz
VGWv2O4TD5Vmb+1LwTMu9RLVuxlk51ehjtdZlmr0EpOqikSZmsNRbV5j1lDelgxJ
DrBDmJ13us1o6kTgcI7h4Ty3A9FJjLs+d5UzBDR7Bwk39r2lswDBMghGUT83LT0Q
H7LVPXiFNm8CNxXLp0ENFB9GzZNr52SVvf4Cjg4rGagxSADInMDv2ui79wlpZBqX
pZfYWcukTngrpyUKMZ/rgPoOyQE3N1oq0nndDS7mELMET5k0NngtBlonkvYMS0/H
gQ5cNHWnhiAFtwe4YCqtjeh5QiK80QjK/pQSEJxLegw8bNw0DABxhrALEK2ax5oC
CJ34KYozMHDDHy2IqBScTFn8HxXcmTLjcEx3aBMxjbO9eQ/NDMfwiPdS+Jd9zaad
wRRo/Hh2UJmrF0Dr3FM+oN4tjUytPT0mNSFRjK9s3fLViEYQYfoSeo+o+91rT+Ni
TSskUGbjAYTwfGqScn8CJ1Ux1y0ROTAGJ+Cs0zjEHuo+P+1ctpVG/N4OFSAHVDlc
Mt4hyW/ZscaNFHq46sfk9u3R7W3uL1Q19TrVuyKqLsaFSsl/1+tkd2oAQ9gdKcOT
9d+bYOD3HSHFfmhXv2PBurpjQtfuym79+B1XGK93Fb/hSAkmFPL59f9NxVJ8Nz6o
W2C+NinWt7u/oCXz5Md276rL2QwAEg1U6w6Y7JgYgeFdRdp4At1fKdmewAMQOkni
s90qQf/ofiGDt2jzAKWaCu4+2XgHyG4qajG/RZlZayBLSOmvfkiZ4jilVexPs+7c
ufhSaHe7WajIokSElMcrOjCo3H0fZDaK+oX/61/rj6xLwZU2ustXWsLphCVuvOc3
qOUTGWym5DPsZEpSXjGsh2UzCv6rdJva2t94JJ6+G8AMWqvrUKhFjRIEUrzqAFzz
VJviiCGlnFqcesuqoF/gI7Y8n/L4V9ajxZE+TLyoB4oX13yxObwNe8n3PLBWwuWy
tkof5BSPDch/p35qUksbY/P59QJi4Q7HgAOzvE3KNFaIK2S4HTAP8VLNdK4zxVdM
P8buoFvcgaHuGqy14J/PxtfqiK7p7jGcp4T0XSSu3Qyz0rI2wreax/3VbDp9keQD
BVaBk7Mz93a3FXEXdqS1jDDXJoHP4k896w4M3TP+EOIra6G7qC3Cjmltjcv3WINR
82fQvr5XKQgHGwEgtzm13WWViC1dc+RrMjl518ltMZOGDvDHErARsGIiP89ovV2d
g+OzgYQa0LCE+g8RhbfRzHthPpttO2D/CK8Y28wdQbDuFS2gCFPgnbpyHFrV5pYY
dnb6mrEPVwCEtR+V/yp9PMOI7MElrjKBJoPt5vglSwTsEu9Dr5RuXUd2C6wIE4jB
LEyg7Rb9qjmTVDjXOtn0u8+ALWsy/qMWOVh3Mn7tiUEYhaFf77qEfsv09ZTkZQBQ
4bdQZI0nTSrNnbs7BhfkRCUsM6Lc+o0nCVN/YT/7GaATay+JIvhS0fosnWySzgLM
Y2E8CfceJf6Uf6ekEwl9sHK2BE7jbaf43EwPaEftKws8ojPl/KjiA9V6lDOHDH10
yueqS4p51nrxYqfpamg0vXj6dTNKRoFhiWvj4BezLvZlQa5LA2krj6KW6I5VHeky
P3KvP89Di/DIovYQhmWlSTCKqhfX5qIzytIPTMDweVp9eBQ5kJk+QXP8h7myamt5
eU/MEkgBYKLBGpMS9+ThB+Au/FoO6/cR29R56sPtP3ofGIrOqE0UYO1W7guhJmQ+
hDxNNQssNtZa/pmo3rt38KGfL2cqCfSQiOyR1BAPvv3friZHjpWuRHukqbPtbiyM
irzLTpK76B6E52LR0uyh83OAZEDSfgEy1NS1SzOLttN4Jnpe1Qqj6ypeQvoM/6Wl
vqTiy3w9Bh9RIRYGVSeHBs/X+/Ct2e5AmP4Xz3NigZmImHsC0oBPe17k2MjEwbk2
Vooe7QZOplGyPUWx+6bb/+9qSCRK5BkPcgRPMTuJ2THmFUe4AJN7px1PZ07ETXZA
D8CaOnxx3z13Ror9qiM4tbm5wy9n3/8MXuE82tLv/QQgwuIC9xx8PvMk2Lhua2CE
5cOHh9Ij6UektSkOzkiUuPoBkOJ+Gur3a+ZquNG6b38diz8haslVC6lANaL2DW4G
ESECaV0fuNw4N0YKFQ2LlJNRS5e1JMirMLAJsAG/91rcD5pxp+QfrOL1ImM4GvJ4
9iqJX1nZn8FjndZjVaTGHEQw11n3Zqov8DUAl/IGw9LcYa7w1lMHLhASAj+XHLtg
//DdXGZqOHDtsESDsLmdUBkEZ3tQhPBkESE2+1drcHUzr+DKbLsXeW5k795fpXsz
ZhUWxmr8Qq4HcxsrIFFMO5u4WD9Pw/M6aneXaGxPMT71dRBCtl8wB33aZdUhumqs
5/skQtXW5rhNJS9HLVlSub95PLCkfDG+4QV4d3BeNcrzxmB7oZHOUcI0fhMrtE+F
Vlz39PUqy+dBf9vm3khEC4QdbPd55SqBA+IqSVkk3POgbrHfr3nhcORXMf1QZrts
fIz6smfIEm8E8mPEHxddknpRylqDZJxW0VUkmPWNIvh4UGxWfKTui9V+uYPns44F
+hnDHFklokN/CEfXQ/Zzb5Z24zMXg0LsbjTaY86xq7SQHIAP+NkhFGeOy/ujjYvq
5W4WZTQW0QackvOWFsZrj7Cft5c75R0J2paCLL5Ms7BKg/7DVDNuVEvW4cB2Qa+R
EgbIepfXHPSSsmj/dE4YjDrPsoHyV7BV2OoZlFgxq7FILt5L0ufaGindO6wSeh+4
awq9tUu8Hj/YQXHCyvII+bcanQGwZ/C/Rhmx0lzk74b0Uvbp/tLK321esRe3lALP
09VCgmr6ztUVuFFSQl07nhWdZVk6MPBb2wpDKEf4f8to246MlQyOvdhcqp1h2uV/
1j54wg79Q5lfoiCkMxA0v2Rs3jZ+tWyZFTVQnLtxOwDQMFbYy/9s07wldoyKXBZ1
omUDeAmkDoGXQMQRpbUUpWiItt95+dbaxDc79/HC+TD8jon0xlDOyNaY8TZPI87U
66yZFi3K634L/GdqQ/c6LTRZQTJ04wRpBWwoNoCgi4f8ayvBjwzmM0nPmLkX0cLA
z+ffV9wJPNA4frbinT0F29vBAwWMcbzRUWYwLpTsimtUEosXCwshdYUAkVjW0Gvs
TOePHQUCNNWylfO1O+WG04HcMe23Jsz1b1TQy8BaqYEOO7G/cwGV/DsgFi8yAfFu
GekpEZJk204fY2mJyrP9upaZHD9T3KcmJ1Kxhj5jV78beWtpih/PE4uXadfAN2Oq
0vgMgFoo18AI8O6jT65M2vO0a6HiFvyAToMNqD8VfZQJGxv5UrjS3WpqbvNhYFyo
h6y5HYsx5Tp2m0n32GL0pZukgmh5IQy90H7rBz5+JNsTcqe0sp7u1tKMxECSYolI
WObWQO+bm2TsnHnJsHhxnXu7VlDCfQSDPmKjQXAYgK+v38Q03yWmY95qWeXH+ynl
DMKdrvfKKD+S0HhOLoMppUHjpVET7kOD99i3Nlw/8iO0AftUMJ379VdIG2RWfuID
UDjXxq3HRTrGPLldTxEKES2b0eKw4UdpmDDu7Q2MXL8ktVenI9KOSFqYGXz5X/OB
RCEWNlYiBlQWFsP9EkRdzEljqxYdGPCmDafCff0FnTkGP0nLeQLWqlm01OtVJku3
9S7racxEnDfFKhroa/PEX0GRCrOakWML3HHfkJh/HId4SFSydHCEmzzkb/E3WVHl
bo0kjbh8pZ8wGYeW3up9F85k9JIaaQiwb36hrjQQX8Q1es8NA4Gj0lfyZzg0Wae5
X8RXNJRemOZ8iSYJK2S8OMNkPWL4WPexROckMQ5DpYCn7ZwnoBGYsUbolvH3s69O
dOoNbk7/Mz+XPJtNuoEkGcVBun//N8gwtgP/nLKxNbP4F0bXedVQhSmHysQA713v
juhRXxagPIE3x0yteFTKWYwOcvYNPSm8ITdPvOxGl7L5n6HLWthsgG3xAeAD8na6
uqRiAMeIi2UWEtNo43dxl2Ok013qkK489Ts9LS/EECRBbNvw8vSvwNnj7i2cSQfe
6uRodRqZMCi3xkCyLrXDNLcU1A3X2tfp+dPvewFw2a2XYRBvzK3CmhY+ubGbMhzR
wap1goxve1GoSo88GNwKuz/RZ2en5xFTr8gMowZsE8adjCMuBDnNV4YW7R+wH3MM
9iBH/Dn7br4ruEtQ2eSViN3ZVF7tk0Wlzu+5F6IlXmuLU6gqnKl8iV9RlvOyDOE8
PKC2KZvdT7ZQmf2QvxmaIuV7XZneOH/2KVgv/SWGqVmUwO8pOcjznURwUh6hjuAA
Oerd5pfg+DdOdKrD04rd7SN8pRqLhgjqPyUZjLntDB/yvKJkmQQFSyyh/ZaxpunK
2Khg4Ryb4p+edp2eIcUevLYgHhalltkAUW/7aJpEQ98Tjk+bCv4TnNcABXXvjBCy
QWVUPYXViY4CwQQl+ulhV3RZ8iFMAwrDdYtHnaAy0UhfdgfCeAM271sKWnzpI3jm
MxISuWFBZO9pFZmxk+A8zExvZXSd/hsVw2DcRdLA3EbWQ0HX6RSgAYvCvf73CmJp
1KNvi2zvj8SO2w58GT3YPDOfWMwmAHf2eNtOzoeb0M999HpJWUr3xR8wMcgniPH+
uwsZLjJIsokqMec4HnAwm8EHgfBveCKzivnsUOeWItvJbGaSs/rDCVordrlN3jXb
8Vd3ZQ1tPAgoWm93B0/LQxzsgAB5c0lWRWEWAQpgg8bQrDSmFmDztgmT+YaZzd/p
Q9zUJL0uje4xoYmUrmd+CMyozgze7/P9ZnEIm78orfuugpgrbGiC3Tt7kRnxkAD5
fmU2g9HBa7QZFkT7s19PfqqRvwq7XOkMHLUV5tERnAQUebXEa4AM7PR5SqTQWbqB
PRdo1Wg+gqp+48g7W60NFKOQOJIlM8I/tHbTxSncASWXjvHnBSXJWo7M22DnffvS
CtsoWp4Zqo3768jiUwYdTmIPIeX4uYRzkkDCJG9d0u9N+dY16afP+lV+QsVMM2A7
XhUY6ebIJ22pqjlwKBDskAJB/AOreJ2XXIjOQB0F/Zn/xN9XqTbJ2FTLy3XZzWcZ
WQQ65aEX1OlIyi2J3saCHXH8o5li0FckTlDGjhayji1Arqj6dh+fzHM+FEY21fKL
33qi003ijLtff7su64J9ve8ayml08tFwiodOiTy65xWLS+oWyGWeuAGT/X4T8OFA
R7ahuopD7vqjP98uVAevBQOjHkzvSzJBW4TBvQJKuJj+Ga62tn+0CZXzAURGhcLG
sDyjoslY7KBZ1F7vT7ttLGsO6FTr607HBkK2WsjtiItD2J1JPJvF3jeUlCXp+vhB
byBbvAOlVfNJcarwGZVK9bnEgToCDKLWSad5b3Drx+Z9gG7bWSSHFCv3f0NdOtLQ
53gL1RCqj0CBgtR6jZf6wwvLb/zRUdd0RlkRFC0sdgDJ3K+1S6H/QTuXwFeODbEX
nhLn6QVrHqls20M85FNUkw3HSg1alAAtIlNvfp+TvtE7TUpstpM4drfcM8zJl51O
YCOeGOviwmWnxGBMxWkNJEoqHEyvnLTwf40TonmKptzC9Ckgskt7zoO95hrxwfkq
1b4zHtRS3TO5VP+RIbcyOpqaN3aRrqQuiaMiWD1Dki7OIQqdv10tnzY7UsVKMFWf
ry2ZzZhgofkKBD+MgYP4br/NwJOfdC3fXkrnJXHV+KVwG3AthljWViPImznNkWrm
zU6fyNispFvIf27GIkI3R/XWGoNoOU0hnkPnNTYc7KuKvnvKBQqoNOVZ7ah1mB9b
wMmmgH2xGDY4Gplu4xoRbbMATS+MxsrYq3OItebkYmHhhGh22h2rkbc/w2dmbLzI
qcXmso+nYM1jiWmlVJIrEvANYw+82G9uROFsMn8VL5K8XgvDTIEOJFgFWErL0H1i
4sWmSLea62hX+34RDzxiwjXR7wshiSjb8/b9DXNBJb82cg126Mr0k6G/dtjmA7oD
Y7kt/HtsRKz9ZWU0owv+f0LLcAcGBNwrSkt1CXsTwukDW2r9rXiK4W+0qV55B4MM
RUEpgJj6oQvWPnzxq5JQoGdnaC5BhIUXPvaGEZ3VzBh1ey/Hu4UCMc4eHBlC5sN8
VeUEKo2xcDnRdWOdOuSsUYUZUdGOoVsePFW7fKPgbRgth9wbem/0lqtxk3aAtXrG
yLPBds6iLezKShgyYAa2g4f1oxDYGIruTjS8cHDmDKgjZxpFQumSrmj3C6cO2ied
oGpomiODHlf+sbc3gei+/4zCNrqqX5Atle6m8bH7fGJdO4zIjGIM5vHyzCdoCRYx
CW0g07z2rlT0hJ4KTBzf8cydplILPHkk4V7KMmjBVmsAqdxnHXeqKd3tx+P/LZCK
qPyxvSTODwUFPd0HzRQqOIJapGXZMyrFxeI7/inuGQPB8MS9Y2SoPV2z1AwKoNUO
uykt15T2I/p7QfTFKhRZHi3F2MZFKPSWFJff6tDTeh3I96JRVLy7Nuyiwf2MvITX
u5m0TqM6wFslEDxTIvtxfjYsNsc9hZv/Rbo28vYlJhVP4ev8IZBV5Y+Npuew/p17
S94I5omvbo8We5vbVWMOQ0SzXmOqtry/MnytNCHzXLt3sdrxn6DmpVmb0XiivcxY
ratdPiJKBpiVUqP6WoMcUAapzwfbaZZ9+MkGmL5mdYM1hXsbj1hXji084PzT/Jg1
GUTNs3CGkMZOYgFitBJSZ4ouHJmpQrpiVdHrK2d6/7O1bwxlDsnamYJkYmDfCVZ2
yN6Vctt2eZ0h/6RE5Ig1/2fLcZxEHZPfdxFO4Mz9d3nSon+ROCuOhx8hwUVDFDGO
EWrbaAG07JeVhpIZhkuppUib3hpvWjE3s1+ncWXDyOO+enu1nVn+VTY0/MnA8uZr
frqgiEWOxhAu4muCDejVxdnQDsQmjSHemxcJNzoRyhYeSVvR60ZKoozE+Wya+sTe
nGO8FpZKf0hYFee3vAHItaf9LizJPZ3MsKubd8L8MSwGHiMmXjy82oYBt5zFQ/Da
TTP1rztSCAkrQgUQwb2EtOvcHEiGAkjlWgVQvg6rQTWrPIj5rbtU7FdWXyLHNW1g
N6ozNHG1VWBzBysiO45WRWJTfYUCq2CYvf6J4uHW1woNQK9EobznyOXIZsGBVwXI
dnCo7yEAlKbgfHec1YQK0gzl6GAMSiDZYmtBjIh1S/tRdDKf/eZfYoPfXOO8y9gW
9xDC2U2prDq7JHBIEd/jUtQwx0CDgkCjaAQHAgm4c29lNjTV+VUHxfEOdqU2ndqq
ol1QZMHdwa42K2yBc+iYT58aY53tTZIsDOiCXckm2O9R2u1lfrqJs/euQ/oJioAI
euqP18YxXPwWVI5gQXrMk82dBvpYD763mLdKfZToGCjiMTgcBIT8pc0fyNMBg3Cm
waxROpCPlVVCvP4/5xVU1tSZ6kywrBRfz1PpwPrZrUIWTj/6FCTfhhWbcWhJDbVs
IssYOL0TxSOk/Mn+tBBTuzDjSoPuSiAHYEyzuD09sWXvR4oWWnl4LGb02kRQ5X9h
zTgDPYugbR3hlhFytqFi4HGAFYtDH6o9rfQW/viAIJsDee3EIrkiFA3xLKjvJL2y
nMUlU6Trp/AvOSDce/1snVVmiNOL/nYDEk4S22ScfvVMJaz2Jl7YS/lBpdXlbidm
XZ5rtBfoaZ2k5cRz6z4g/g8bPnKVJGhLjblCiy9qRCIGV83YcHViP84W5deVxRV5
H85wLmjHvQDZ0+f2jAw/A5fVSnYaIHbYWoZLIdsENg6MaKmVvFawXhUPiTvOid7e
5fKW0ukutkaqQBOh77fvdC1PJSZ/gMnZ6GGZNEbg3Yz5t3x+GK2kDV4iarvtlE0g
FXOox+LZbNaFx7OryvEMrK37YrQcgQBK3Qa5LQJ3kMmmr3vlJjQsliv2ABemVCd9
O2sBO/DgA8m9txTOxMrdeM4BlmpNsS7jggeLYjoNNRQjWZxh0J9Up2tPKjb/pobT
zfRsYqqI5twmUwjwKIVhyUilnEA5Dl2qGSeWyS0RLHrUGyUxM25RZSNCdzlfIKLL
NZ4W1xuKo8jiZZvsoLX54wlLNfJ+HEiQUSM0UwCaozN4usST6kx3+X1D9Ze/4jly
Qnp4vsErLpzdn13jYtffzFKBJrfgn7rcMNFFyz53bDhG75e7nRBAIgZbj97XlBZT
EtIxmTo9YxQB/m84ZXeuwYUFerivUwznC1gFVwZDaE041DhHDrRHgLCaohywmDLd
WSZnOj6pGQR7Tg3hyOPsAH6Ztw3+DIl6rVrwKD+zMaNmnOR+0zxMmG2G6Jrd1APY
KvBbGkX1528lXTUMqT3TZ48YMccB4YhN6Aun9qy+AZEvx0lskPDdVpvW/+HArd6W
QeA8yfVW5VdlorY/7G4D9oGomlIedu+cXUggZ2xMEE92f7jUx9C1aMXcAYDfj0wB
nuv9Mdzpa33sw13XWwlk1JpLTbQJYBYq4X3aA0phD6dHE4dzg1ubq4uYK03KyPQW
8esvO9wN+RSiXOQ6BQ5bZRYfz2EVROL5mROIVnJsfzGskiocLymLjsfcgDpuHjKT
4YbDUltEpdfZrrQR3iUDeNvjX5rjhw312ipTPBkhuQx43lWVP0tZjw8BAtvA3iH4
um9cychs1XlbkUlKWY8Jh2DR9KT+EBk7B0m0BQRCXbLXqsPxq8VfuULwr53Bkjxi
eWzeokysL91WSEQw1AKC79a3uSvZm1z2U2xdWqHjahGXQO66u9jqBXbAYZabePgf
uCcbHGZaDx/IalzAySbhcYH1Z5YdqxAc0EzLnyqXFvamNBzKOj2ihP0+AFjWF0g4
qeLtd/FB4JgJvJgKHkBYhhjQdZqyP3gMDlHMHfRIYKXdBkpdGMzcaxQpEd12+aAI
TEdRymUBCEme9JppnHwz8gwPf7vZNIY+VzrqatsHNZ21EfmIAZUea0cUs1W4xmg5
l/n9IQhH7+cb6YS+enMtCYEp1CEWFVfys8FzxqRyEJWmTv5tvVzOQKr1XfT5r1ZZ
dJkA19/p/G3I4rFqxTCT5KS/zG0dLXlEtfNPDaXReS/1u6vIQg0Phe18J5EUCelJ
5EvTDBZJaizEDrxr2BO+H/EOD9shPg17GZOCIvEGjenA3tkoYwRVwb0QJpOD/Pf8
u1rOFc44qPwzwhqd0vQwZ4a2fzSHwiINlFsHEKz95pqB30M61ID65R6me+13JPZf
GboDQ0T3/A4U5OpiCazQxRT6Guuw5dSXXCj1RjqUlNo/r9bEFkID4Ts+MbNkfRmu
pOORWO7T0vv5qUKZ2DBXyxwACCKcTxjfDXI+wG7q5USHcBdAxTym6OGOtpqwhomN
/KLFoWSlSxaoxMAb9kA4GpkbBjUHaLu4I0e9R0kyMcgsMKY1Rrp3IlQRhi4ymHIW
dGiq77d+K0waPyCfgeB3bvlJJ76njIcem2c3jKG8QxIF6gwdrVNy1H3OmZlxpkiW
KGIB0JTk/2zoou1MSKb5XtgXLbKUDy0sI+mgebu3cg9DhA+rJmPASYuo0WAH7KrD
/IEmuoHmJUKhSpzVT8HvehA5VwblmDksTA8of9rmI7iwaHtyDOBbdR+w41LGdUnB
eoljfPTJO3xz2moKONGjAqKWouhPGK/w2Z1ZWrcAUVzmiARKF+QJIrkOXP7jVz5k
hlV46DBvBsBzJ5BFUrZTwosP34DKNBjAgQJjW8gAx5KKHBpPQlF1hHLlI/5RT37G
ZD338RNXw0tn2Gy8GGPbedff2AblS/SWNT9vThHbdy/p/OncCUCsRK0RxeItoWfA
7GBSvyWeEPNNXeu699PYAEWTsLjMwmT6p8UiTsI9ZENHfRBSvttX7wmc2eeIZ9wd
ifsTWyLC/Ydnk4ca4LprVHdQfiEa+o8u7xEWEKdVRZOHvGJhC3h+cfA8cEuipjuz
zMO1MsZTr2uZ270wjv6ZStu+XOc6wK8SOQ17Uar2YbQ3luksjOJOYXrJoBdix7bf
wCeti96gdd4eGkPd/kF1OTmqddDQzCF8mldSE1HrDP8WaI+AU1SgOCR6gy3XSGYv
MfQcRL2tkNm4/atHsH5M7adBrzjyAw8UWfErjFwo84EWbsBwQYXU8ZwmHtyUiUoe
I+tf9Au6DBH7yEyVH2cN6wAFjdfcESh+gNpm4CQ8meylhktDR1tzOCucaLGXYN46
rYvcofVoyvY0KO4VNwkm7keZey+v06EDYa+MJbLKIhpftcBxXlamaUaigf9DugE5
kDS9lYkAjhsiYmJWbjOBA4SKrIbCmNDl44FYgnlHZXmhUCkrZv2L/TJampECtmq/
YRKjev3SuKBd2AmSQB6V9psCTDMolCJmQKrLa9ukAcathTOJHytZOjEusVOnLdSc
4hhI89q9J5TzwC7NhWvZFpJ5s3zjgAG1rFb1XO/sVt4R3wFLmcTmShygMVGk/VKF
QwKmXApJd9uI34PtH5i9x027aU+Kai4qMyWhaBSNUtXPGPt1aUeUB4ZgcHBJh3iw
23kajMjW4vFavEgKtVYsTGMv2RHY3mf6cAKWzzxxBXWMrq/8625GDviOT8xB5FxE
zzRpSXH9LStrB9TmsyPwKb+pFgGGO9fbV4m1JrqPSH0brNAmrJdPClgTUad59LsZ
GpNkap5pnuDRhihh7UwSLB3Q+3nO33HM7pbUmfyZfCLYI3oOQP2YGQNU4lPK06dT
Pyzwt1SsS+FEN/quUXJFsVE7JOdTMzHDTLdLijmGQx5hwaBBNpAdW2NDhrOfLU0j
d5mxtbSoWJ9h5wJhjeq2GlSkrHev5Qf7NKZOBcykIEMfs60hQX6NfMm/vNalDRTU
pfIj6mfSmfuVCiZgNW1wdMg8wI7qHFWoCn1CM1d9S9+vlVHekW9WZQjSFhzdTp/U
2K5JQcBtb3CCXdiJDciJpj8CB2rzld/x3vlm3mOgd8bz24ib3SMQDGt4fG4nHjkL
lxJgQy7mr/Rqer649+kv9pmFv4rX9vYho5kVU2f75Kdn5nhsKJ3Bx/PqAKd0b8Xw
ozl/kSR/Ohb/VyR6VP1AllUkMRzPG5J4glWIsvsNiGK8ZWlw+kGsHWcwsj++c4qd
Hzo4CgMPjSEyGvAGbv+kVXHlOZ57g+GLby7964gR3pZZLzfwohYXiQ8J5KYyAndt
siQgXyySNlD5hQvhHQk/R9F4tRKAtLkSBVmx4tI76cO/PBLxpN/36w0NIMWH+9XQ
M+XadbdTIQN3kAgJSWGEhf1fZF3vD4TMB5iOHLITSzCf44iGkoXmb7PsOC4W8ewK
Ed06Ayl+fbO/TD9JlVrqK4WxwHnZVvibrFEHz+tJ097tLVSJDStRdrZb2cEhWHQx
zJcLeH0AE0pldOYPlvzVo0CReWkUZhgTr/GTCCcKNfKP/nzARvLCdCjTrgQi6ZjZ
MG7nWudvgWx3gez/bo+psBEcxlMpYo5Yu8hNRW8vTSH+L22yFIMd7KB0F52log4i
pFl5ZT92k9H+cbxI4LlFPCe6rvNn6IkFYrH4bdNXPjoXOt9qinbdkjdzJnUGmCoT
6H2WsgB22KOG27PVESZIw3jpW5Evl4caXuwrtAEdGBz3bNQMG7ZktbAMLDOwvpUv
qh60UN4ubBPE97dlEOf1PcJ21igvgJFzLm7LEQGI92e8MoUDWzIimBBLzKRqzLPI
p4P3ItB3w90ugkShJtCFlsuhfYe+Sgrwhb/LQwJWU7r6YHmQw4+F8iteF2XtAP8+
Z+M0lquEQiTxk46dphDosUAMjInr/oqjveVLQAEt8wcUjYqpuHcHOlY88vlf2Spc
ZU8CcYAWaHiSyFE/+Zgpr+o0mf6zYDDd8EHLiGz3TbLX85EhJSYdfj5rAYfGnHsl
JaxqmvB2y8JnuicHDxmRwoL8zNJPRh1yWESLs3K7VKSZ+8oRDTRrBxCM7k7sqkXI
FbQDjbqZXtTabyXvkvHOlt06n+RVpG/7yWlr0HadaieRyNUcESoLjqZYO89EjXBO
pAbb0Bj5GgdrUrhFAvlLXtVO7mCA7Z4HULAtPjxA+w0wDmDYrE+OY8fNO3IBFCA5
2iTWYltNTRS1hWeBPI4oKsAIyl67v7BUjTr8cyi1LgIHiYlA+OS60/+0/8yUZTDo
mQsUysvNLEmDxq1X5VMVOASUq44hah1r5ZP3k9RzUz2RHIGjj58HaJZPgMVHX4Z8
MHj1g9w03YSYvHXE1D6BlAG2ewhLewXzVwtHRU6ohq24cXl9BaqQU27jPAl4i5ZP
6yn2CEhqD8zeokBGAWJjySWdIJyGYCIU1tqE8k9hUNOHQiC+bBWjmMnFE+aCWODZ
63gkrm2DHrOD0PGViarqL6eCjuS7fMyQNqMbJXSQWF2pf4E+rBzHWjTMbcGDltW8
4GQ503kj61MCT7SEmIbNtKVDTGUdlbJJsyVkq3eTjRBUa5mbPGfGEZClrdNA1sTS
hRfdcx5DXUDUfbe4SNBWWcxvWr+lkj+BwrCLZLp48WeneCRt+Iqdcu3lbCeYdyAs
rd/QdpohpgBeGHCNsWIcybXCrJeGHHZ0SMWK5a5ASs+j9moY5qGuyNvaK0bmKi2p
9A9sIQTS5amL3NKVUQFRVAJkBGqUZBiaJM4iHHncS8NzGIaZP8mtBAzonCnQ/JQD
EMQZyuXx+GbY7i7RRmQKPMQgJ3Lje4vOg3OVIcDOEfjC9OZKqTUoT8jWTWNWemlM
B3fPdq7Zpm6OtFQuey9en4VGy2yQhPd7NwvzsL0/viG3BPLCym/qyGErWJqkzPRI
ZR4AiBeUDXH5r4uNW47S0lcjF+527h4Ia9NSnGO1rQqYOIiFIH6njz4ERgiRO5JV
aE8Tq9GCWxkvxIQRSB7fIup+ziMaZ2HlJEHOwsDROgXtN54iVXAQBvNMsgcJnfx1
A5svJQ36ES2QJHTBMJQL25ELfop9EzubmwcNhc4XvfUk/abREVuqL8mNWJXPAk1f
QwTahD5tF3+ITF90F4Gp1wSEZj06V4mZrBUDV5kgafPAY4TFMt6iEFoe/A7DP8I9
IhHjrt+BkeLSEQpglR9P0wW2BBjTqQmap5TRHJI6NnDGyS5uRauDC3Leyz2WXel/
V29SH/BzEJG1hH71MNqK3dR9yUgcoNVvxkXLNaVbX+4qyNBd3bRv//UF4gh2WfCx
KFsLity01V2gI2DYX4p0n7Z1KzQNfNRhZfw8ny6gdS49zQ4YhQ0CEMB7ipvuir4c
3G09gejzR6jxrhE8tHI1lilQYBt88ZK9PdV+gUxKG80DIwgx7uUukaw57az4DTvW
4YZ1YAwy7OYSe+PAtH7lCC+0xwtHgbIPlVOEcEtTB5MBZ1cSfQrTgk2EJbfZXh8l
/UTaunehE7mK7y7sk0Q2x93gjj8hR+dqEImXN0sFENr4jiA+YVAC0lZ6RlT5c7FA
xRWZHeTESDRK/Eg8Q077C4yE3ziGaStBNJPEx/XSyExZp5o5IDmjkKaSFlJpGg0Q
oKYF2dD0ODctTJi9PsgP1eW1lWHyBtfRQwc6fWQvmZA1tRQCwFFJ6Y9hUmC+O30l
vj7wDZnhJk6QsYzgENRiPHVG8RE4Q5JPZv0Mzwhvm5U6gxltT1afhpZBR5mRTuCJ
PKSWrdzZ36RMrEnAv2gGsPTsFQWCIfF2Req282xOsUsfBI48mjKe4H3nAFu2kgW3
4Z9KsL41KYvWOtV8YAL5VNsGKp4v05hTaW4Q7ZtY4CI3cdox7/2qhD7TIWr25sLO
IvmYi2Zh0SLooVPmbXaO1eToIzIY+oWM2bM7avxHvGet1ZpAQ7pkyTioGjnFMfox
+ULSIJDGKDU7wz30cP3Rqj4An0Z4CK8Z5AwoVDV/2YpePrUahL1c00QXoMyaFAJi
CXa/dcNhuUSwSN8jlRkZ98jF+k6fVgiHsRQqqpHk/I77iqEGzmikdX9w9mVMhaoa
RnyACXF8P1YJnym6lzqO+5a57lqhrOVvauGQV7Ulef9JnkZL/Mxb7OveIEHegflN
9t8fUqkVki/8OWRbXuWUBVgXVmLDF3yvG7oyRz/NC+5Qzqe0NL4fCNMGnF0b9/Kd
DrmBJKIJz7dPh07NsomLuJT26fQdn+DnMR+MxJgUo+Fo1Mz0E/56d+LOMOxoZiYx
sVH50Oiez/fH8GDMHjIO2Xz88njkTkLOw3TAEV17C4MInaHbaz4kxaaJOMt5uOuY
58nhlkOo3rqH8pgvCYJe2VD/QVGQIxK3G/mnzXJ/qjFcVMCNK7db0HfkWJ6aE8KV
SNF8tWfo/+P+krl25ohGVjCh9qIv0wj20Y55U+CTncjOlcnKiVw0ZzgA1WecCnKn
QJtNK2mBVDNe5+T2p5se4ACuoeY2J2GSb5TgW+w0e689DVukSeEWPsfhHRTOo5EI
sT7wcjlHJ+kILnVatCvdZX+yDr9NiHE2IStFhUX0mWNLnSGewuYrITWaJXQjzrIv
HO1dP8uHnSaYnsEsyeKVBGfr/zhi9tTWmzaYRaibFR+H5hEzQvWFcQ6oH1F2lmC9
fKP8+z+osqI9qyaVOVi+KVpkNNxpUJgrkrkmuMT+Jzyz2VtO0IerLc4G/sJOY8+p
/1bwIF3QY/iqh8em0kKIcJBP32njVqllh9nH0niX/9R1DirvB6Lqs1zAKYGCzm1a
jY7Ag+ESZNXXj0u4nc6tsgP2wa6azObQFjM80ix6cjTS6vnqxO3lPxvBmhtu4Nxp
QgUhlHESKk3x1bE4q0zZuuQIojpXSiyI9VZu5kzlzX+u1CNoPj3g2cN18XpkbykK
ruTS0k3Og8Ey00tT5e7KSDp2nVFDgrMVDvdkj0jrjt9BzgVZRryKKhK+8Nxic09/
HLzf4NH/tEWo1C29JtjiecdTHFg8qUj4KbVseGe2Bdta+w1/A0HEmW9Dq03nBMUw
mj/tq5fcpRDjdsBAsuexCpJ5L5eLRzqNeJF8WbsXk0tJWcaPzw9JXRaJBlKccmJP
3CUPYm40oqGh5pNdzpGfBAIQfQIgNbaSgQZ8Zaf99nL6iLfd3K4QvxAgdHgnAHj0
nT7VH6mON32LJeiwx2ZE5+y47/E1kgMUmYQepSRrh611f5JTe1AHlPXhoGIcLWek
3Rxuc1yyQ8/wrNAVeIsynUG+c9LxlOhr0h64gE3wDAwDTB8ygnd5qY6Rbj3nWkzr
qctspmp1orxRYIKf4kPRICUMKdAyVNiQOdqpg0v6wNtj8OjFeTg6W/QbsVwIvET3
NTzTzvKYFsRHQUzZYs5sGLBSdtE234RPQ/Yqwi/NGverQ8G1GDE0jHO1nOZjnR0L
IdcWYz6K2GbdS1Qyplv78t4PMj1l4nmvjX1+QMCrv39YCHLmHTsdyqvNO5B2OoBw
C2ltvENe/8+Ys36b4BHyTMlBP2BUiHUlS/b/Lr9HkYsMEQ58q4Z/h5MyuPPNONW7
iRXdWRvDoeDutWAaRvz4lv1KeK4slWFVGh3Nx6RAxKpxTU3Tqmcp2PYgjpVor5Z8
AApKMeUjauBzmrsUyasZ53+cnTfnCBFQt3uZVgKxIIAzeF+EkSNf4ownx20w4P6z
E04+TNO26qwjXrOdCvhmVQqvf56xeIQJaP90rCozce4Gl7rI3PXGaE9DEvMdeZGE
v5SfAsAzZ4QmGzqr9VTwzENd98Nn612iTaWxYmxug1uFTiu39dKlR2vep990PL5E
udE6EsZDPp7PH0xcFmd/eJwuMvKMtN8mTI3pUtlEKJcOuvZN2+V8UOec8G09FC7u
OotANYw8Bu0n7zvo6TtYZPkO8frBCMRvBBxVFGVweo8H2cs681dwgft60Mv1F/LL
tOMCO+Jg8em/3/iqL+cSJsj930ioCu/aZqYZT2YLGM9lCcHOBOubKLYT8GXXC9Ds
EjwUdrjmhs2Sm0KV2g1e90cGfCDZULCKy9IOlC07rJfcEL0C1I9GrYHSFusekD26
dHTuIK8Lrz7Ir7YOHKW1NdsJotLtPaY8wazZQT2py7iDXtuMsR61+fM7lH7tkaO1
ABv2qP5W/7EQw7B5xjwrnKdY4xtV0Ufv0XdU8UHrnuXUAnql6q7/G/pt4Jzgw35D
x+QPOrg9RHZ1+OQga01NuZ/P+pSzHkZA0cL//s9sGg7oVqLCawANsOaMVxBVJlCA
1tTyb/yB1eSSn6ggjgrxxMjbSqioEDJX6lnYpiCbzIuLkDbW7Y6o2uX40VRkl20f
1Ve82na2JIY8OSSyI2zOdYZgEphHYTlcG6ZF76WrX2a0zxK8yI9wZg9hf2tVlzhZ
77gs2GPF8Ru2AZ8x7xdZYfCoS1xB+8PZHnklSOs4rqKZvxm6IBfjFFQ77LEr7Wgv
D6nDl9Bcf05rDJXka7JmSyLIHcgdXQuxms3dD0zilctRjJ4+nws/cMvlPels7nij
p8aeb+/3HSr3GA0ChP+dZWmT2Lgz6l50pxHb9LtRsoVC136r07rzS2a+OSWDmhS2
rc+vX9aJNM5RB4NvgulidpL9GU1i3KunEOVFeWmM4kiBA3O2LrV/VfBcmQlo7kM8
f3AZUKjfntkrBvzqQE5CJakCKVqZxF0jL7GxtDmzxRUoHYwtPuv9x4giwf0IsuAi
Ou7+EF/75JZ8Te9l1jGPxOtQPiH/BI/8mhjU4bpVyoqWCkfArxycm61l6UGwN34M
23LFDlwa5uPKj2KDmNQa86COMo99/w/7ueAFviShkUg7lrdlMNDT0cp9JsJ/zCBD
V2kZn0qCZfvNXxcPs18znXkYj0sJpz/6/0gYaHI5FsRN51VRwL/v1hbPuQIN2NH2
q0IEGTOK1L5Nj2TCcO9uzLmMmXxrUF2c+EeXbFYATGpb1oOANbDHItmkao1qDrHh
z1pJwthOQS7X+pxbBmf/6OyQeniFS6d6lMsfLbq9FT3zKNvgP/IoKAIogj1KWxRc
5qH9jn0WaVa4JD8tHT5lPaVFiu6xh0RI8kTn3sMe2TodUMw4oHrwRauXilr9lpJD
y+3HkR1Qf66g4RVy/cbhtJtbGFCKfeByTtY2jNHcNMsZnh1hOu687r1/T+DbMqQj
ptlsN/dqzDn33kBSIluz5G3Vs+Zkg7XR5myMsUuXxJddyYPGTIr8FwWK9uYV7THU
39pJ9zZ0sbOy5GWYmYJq61zRTdXI973lR0cN4Z0tcDytSNJg5fYwsc+XJDHNeXVx
+Nram4qvPVcPLThJOyAdtvTMAOb/BgphhaX9VbCyoRpARIkwrDywU+L6rVBCWY/g
2ul2H8gSPxX1ROfb+8Mx9TKipWd/Nqs1R0h8kh9h2oUJ0GjQtLJ8NtLfNxjCTpEc
pVrYy8vvIvoqkahmEJnEIn1fELAOXFb/9UI8wuJhCom1vkON9skDWRlj4NH8Z0Mi
SUzJXM7XWsiwB4Id8FH7NTlL6IS6+jAZ/1SG+l83uOFba/GtpTla2anjt62bCsi9
SXJ5raBZN3ZQtcJ871YUPBlCdm+STJCyu+nFq9+QwrERAqwfPEkw/nlF5wEEJA1a
+iirLtXDfSgd18y9w/8hz/Pz1aWBFjQPwO3J1AinKDbDkDvhdSfsBqlcMiXqMn/f
9JfwYGxY57zKTLTGFJmU/oyQ9NgEZ0is9wM3O1WWCMIg6XS3UTYnHJLu3ch5FFkN
ScSwsaiEQmsBDHhs7NyTM/lPzeKJJkkkUB15Z/7RWUAWYhzShJWxfU5omrCM1RL/
LCBpugFi4FXSfbBWKHCjEPrNrz0pe34u+dqGi7ZnEfBY319lgQwCwzcsUxqCqxP5
PSRVGNucaTF/m2Xd1MvZIPJk7R1/CJCBvv3iy/TIFy7SnOZ2nyU8XaLop5kiuClk
pQp+jjqh9jLq/6Tt2kmauTrYZZjpWz+xdYmi19zz2hQwPpwtpDlD0BAwkfc2wMlk
iR8pWGbdtQJHPKTZv/wgCw9cErLioNBm+lKLD77nxRiU99wUVnaee+JH6FsM+/GV
wl6AmWRBEaop6vQKbY8nJeV5h+L64gTGorvKWpF7AHI7Gznys/1GnowERUKG7Hg2
f5wP3qBIuxhCSBTH5Onc57+j/MJxqqihgzw8LoBtv/biM8anjAWMGSO5F1t5oZcs
QQrFLs2T/Vw1YQ4IYxrVzzzjzymu7hprzCgHQjapS1twqmI11ACamom9PoELVDp3
kGSJYcSzkrS4Q6srcGeTTFq2sXyWKPGNFa5XfrM3C8MsWJ/aaCeLo3XpTWIomZch
Ty7yNZ9pM43rto8kBIeO3YAEzja3qP1ZR+tdsaK1vVrKps/a+hQd7XZM5LJ7i9O/
kgDz2svElf8hYzDvZWXdScLzDM3bkKRIN8vx75r4qnxs8ECXMUbBdRxRgNWUCrrx
Fml83uV20ARtyjahfm4wLNa+jn5wDkj23ERg4JrT0LeVHXrczesuYOitt0ydPzx2
s4hggUCWryqKA3Lvya0tA16L0H9Ltjouxu20vR3VUFoBGKRWc0IRrxCIRGKWdg3Q
NYUGej52LFzRc1UEVkldroYw2Z0HcIiIS4vX2eO+5/I0/h1eMwlrbFMcK36hVicS
Ozdawog6hM8OLNVHLVJnIUp6ZmLwEj7uQK8fnF9juSgUNc23ndTqa1X+CR+178E5
/ftAIWtLo5htcII3r7DV687v1r6xc79+1RUQtM0N2Q3lZlU1wF9pZrTl2KqoPv21
0z2eg3gDatWULPTossCwIvUKS5Ln9BklMjWOQ4EXPucIXn7GWx6hhQRPjVPcJ1K5
r+elK4jgkwhqZB0+8FlHIT37OfZJRi/I6hXGnXaQGsH4KfTh4QOox9yDoEOKUibe
Ae4ITBdq+FNrWcMZnOCXnZlQ9/BqpQuG5JzSFFFDsjItc6F8QQfZUJ6LD0ZeUis7
QqqGBi3XX5eFAK9u6HHL4jDLfVBfoeemueYgQLfk5FzjMYYAgQkIqtpStUEx6knl
4kpmCbUKmZTwGRH2jyG4G6dVrsXO0sGSg6YTqS5afKF3gmiEVhDDxvVitOPHRklx
GwSicpq/Qm2xsXXuOC5fioVZ9ML29HCvvMx47Q86CwerN7R48XzB+rSwaAaFKV8R
nYE7gH6Fd/ZyehLO8izbkR1tAvUYrTZGHP/69MMl6Qdqak7aqSEFb3Lj5waMBglf
4dMteBG2w2klCtLexrnCTpIuA13zfoVa7LzsBnx+1fDvLuRSsrrlQ6BSzHdFcfuL
TPzrdUCxDaeO+6nxfyG1D2jhQKtOE6RE8lspdDOde0WkXb080k5JI8skLzrH6ORo
oOT7KFGZYkHl/9Mt+tl1u2GdtRNA9frWbvBLtNGEWByFPzmTzVEc2xVjDVLqhI+j
0okPHeBxy5yRCmMkRaIoeiLLSFMwIi1ptTz1+q9oeI3qc+Tke5DuAznbx0Sp0w2N
Og88GNA65dG1Na7N55Me5Fiu2GkalWGk62yxPY7qBXjkyamgiVILaOKYaYjadmOG
n/gEva0r2ZFqKwnh6xI/JcCj+Xc/uABiZPpbnZueId3lSobfFsL0HB58izEFQc47
HEd3x19pLaIoeuh4pku0qDyev8nXFpLqvSwOCEdyUBjBsVfQt9mDKHseEhaD4KBQ
ybuWvjm3EWYchyHxpTjXvavQZyxicJhVxT7smGLEQKqee8urhedkIK2iFsF+HhHV
0DzCrS/yeOJb30l10UaLGxZ4xUVZkj3tFCis7KK78bs1TbXQWwSR1WScC2PoYYkl
UMuISxTMU7L/wRXBbgCizkvtG0Ry2Y4l+KYGeGMXbAOppD+4eWIhOYJTSV5XvEwW
waRxqBBnxcqawE09c8+JUs+1rHWNvCmY2KEdNzz6rWoixR1mUm3jxLEs6KyJyKqL
hx7dhY+CZyjpr80TWPXhOGirkEzlvpW2fomM+F4ofnW+L61SZbFEnnY0pBxH9Eyp
4i/tqyoV6oCfcXjh5luV/HXuaNO1bzWAuw1oyIZhfNlYZ5elokWysMrsFasH6T4T
Qca0ZrSTc+fEGm2QEkmsmb+zJ9hw6wTy4pAoP9uVDUOogDlYtryf20TkiAJU+TpR
h3GA7s5DcvY2/5JcaW6Qi6fvTUURG+xYByTyytzqSjpDM7k8RRdLL4+wpju/3UBc
yY7NNL4JmUtyjUmw7HtuQCd8kkNueEbfHPpujd+0AFOx6M6eLXoQOXcPh98X4s2y
NNmE9oyJhmWwIxJ8dgjnYhpXffzi3E8Wazbi0+VOYYqSAgQyqh5o8Y7xNdV3Vsg8
QxV25y+AqVAYxNFGGqQxzWwncf8K8rPQWmrTokj/Fa3/ZwceEUxG0BkwVxQU/4U4
fRAp7Tlfliaw0jBNcUYWulCbXuXybvFr3DABKtvNZqcZN6bMCwL2KN9rk5cRMg8V
Q/Pa3wvtJ9JPRbLtC76PTsU/M6pRLh/TxH2bBXvDZJmqvqYA8SZSuuzAshajaquP
Q1tKp1tfHhXdFSP2rf+Kg/QdcDcLs3mlxCHuRAsDC9mdTAKPzJkDNqs8L3cQgs3w
y9oG/xKjnLH1n6IKTijVlLDuWnvV+Stdm0+ypBggedw59YDhQyi9miPOcNUy/oHz
N7h+FBvxmg/EJ3/FVWP/ppU9pGcq7DE0wAk6mXjFIfGEAIJHBbtILuYnOMMBhGOH
FqNHVX3+J3uQuDz2tADx8S4LyVQiCIvwqyjmqW6XB8tuk/iAy/8tAaL0A1zSrrNR
z6lMKiP0ARAA0Cz9c2pfEIoNliQEYVw43VNwLVzi3pIS5l9IMFfHSE9WR2LNW2aN
JDdgt8UFLQgEE7BUwW3QdS+bWUQoQcWQtvKumJZpEs7AKpPyKaAB0ndhT5gtILlR
m8h3r4Rdtf2o/5nmYbmg6K9XqCJt/mT4hmfqdYacd2qtsJ1IzrNrz1X+Fxuyc28i
GljRCvAwfskFEU6DuxKZZmPrBOo7ln5oVPUuin8D8d4MlrGtnCqzcmD4CxRW+RsT
72LEVcjJwUvJYolqQYOD1lu62aa1XNlJ4XfHQbDUmNSnS/2MvGrZew1M2Jj035uv
1ZDYO7yks0nJuSDaNsLktX805vCSYZP3mBsa+m94aM1RWa/XBjqBDXl94PHYejXf
IhYBBkJ2g0Ksaixmhkyxgf//rcXNLHaaX15L6puSFS8kHf2aPi8f9uPm8W2zy80+
yRz58iflDyKiAWqsmfG7HBvh25YCjR6o589/j3xPXybCnviHEAEylyR49pAhcrUD
eL/BwvZx7XxMGI7n/dhY/mpGfoiWdmqzGX/r9L++1jdV62EUey6hEvhkFgJWPP8Q
5lBeYQK3gJfaAT2QASdMCJSWQ0o8F+AdMPZbQAM5zH05u53PJK6npO98laWWZruM
70br44cSVKbv//JFLX2IeJN5FYQvFx3lB45n1JxtsCJpIElYNgLN3YgMaBcNFA8g
w4bgcNZ977o3ZvQAE02bjU/xhK6JZrLQVaIL+A250hR1wohiAcBnTGCa9dhHvYxw
cQ9r977BzR7LkBXzRSjKyX2PejG3rl4oNk8Zz3zkIGjOX/MgkKCXvv/H7I9XwuJd
5H8jCTfiEBG/8BdcDGB4d3BA46dCWv6R6gS0n4PpT+neYkzfvznWs4EKIc64dCYt
R2wecJBtRqzh8uJlIkLvC1xRklV8nB0U8tTIHZ6kpCPLGF8xm9WPm3P5IXUV8XY8
Tob8PjTw0xqQWVxgdmfraFUCIsncUUTDl8fRauOFa8ZmBsoYKd96sYvAgrLwM5ns
2eswCvy71qPayMA0ssvi5lr+PHIffTcaHBjY6PXpzNXASKuvOaDF6FrOcMnzr3dr
PTzrFLn30RhctoTvN7qC8YrhJkNf1TQMQLSVt/OpjcoIX3/ntiKP0gBohL9LFjwO
fxMZI2YVGQg3/oXNnfDeMrB67BUcU6Ew6YsKpZZvoS9gOvhE6meoT/nA2jDPuDbg
nvYO/HJjSkpY3pAnRlN1ghh2FE9mQoJdmdSS2mdGeQ0ouA47BdanXqrAJCAxWFES
P/UrCOBh9aTR3ljGwygl4betKK9v9U4PQNuSM9T0vIfAbGXOwfZlxOu9AToaHr6C
jhDnL6dqcYUV1DHnuvLBiqouP0VFqqcLvkJfyGl6htNOIEJ/fWDHO6uSlV1/znTO
8rI/5Ofg5qbhZbqmUN79bY1HtVoihyeY1hgbZQo5W7LZ6u2HwgfkJo4vXFL4/WM1
LQKQyIuck9n4TButxLaL6hzcsrfBy5tVhTP3ul5DMynumYQKNZJVaY6myI1sCMuD
HxCS1PIghNO3aXTwmTS3bH9s6jSDGfeDlC7pEIgeWXghGq37DmjBMJGP7eVEXRzn
ACVQcvcPu9uqWZUYWxS4pUn829o/wqrWcCXRvj+HW4RU2a9P631tQ3F2656AvtF7
ZSN3vAl843f67TW240XRbuibUK+Rw+ATdDJRpcf8ZvrEGlss67CCQa2emIrkbiE7
vaaGJkoOxJU0IHmjUxtc81qT/jzwJQcNJd0C75ep9hn6kRyAak3ZfORsqlyAHhPV
bFxe6+VlaLH2q7dZHzuHADyTjJIwlzxxMwPWdP5zVyi+v/30N0oGrLZN7bf2vs3U
mAto5B78MEuUXjAzoQstq2p8kn0ZmQHa4myPotQF0bVXfYaahVgjiwTKW2fWmyWM
At5exMwJPgnG3WhxbiWgf1kmDNBO5PVMEExMHJ7g4HmyMjCAJv4ZyMwq6tNacbez
/DblC/qqb5fhBUP8XBZ6gj5YKIbzzVo3B9CCDa/WI6/TkLiX+1PjuiVhqDLZQ50O
Bztu2yzFYMwC3iXqvr+Stpeq3hDq04hMgMHONozgataQao1TC8yZ0h016BN50d5d
p2aUXMVHkavM2MLYCRT+SkAS6kqEIWr1kJZ1tMohf6xACm+E+L2yIOkaYnIU1YHv
a7nB95/D1p+D2BsVXpbScxC83KRTS8OxBPGEuSeo7mRUX8OHCG6jx9EBpGg7olq4
PkwKHAQjvvSF/XxNpEDAFib+LSp1XixrhvRXkEseT0UbOxGi0+MqWDj/+kihsp9O
s/oiy0ALE6jdX4eDqSGOUK0MNR/+wy31Sve9Hcy6j52VhqSeBhJ03j/9gMsa3hfA
6IY9u4RY6T7F1d/GxY91KRMa6GGR/4Q8Gm1qgDB2B9+DK6YncMc3yzp01gzp7k0c
dawqkeVB3Ps2uONBG2burnKfLGUoa9ICyGCQPx04m2/MYBssQnhNfXrqsn2fh5dd
b9vDCKTSQSLivmuh7pLGx4/+vXlYZoHm0PjfWznldMx0wR3G+yXtkR2pp0rY5jl3
O5KHLKLeS3rZrtj1BNojo5fbnd8wuc5ppV60sQVmDa3SjAwZDcO+IPzjP6lTOOv+
OzHfFVfaKAZMh54wJ5Bd9WvxteQ3jRcilqFVSYQ6yTvvPBhsujc709xsDG/Z/2OQ
2d9R6wU12SO9GQ086NgEdDHzm9N49dk6JYeLfvnz4gzFoV18PDp2W/R30rteZ9xT
8JM243+nd/X38+PxoOv1ezpfPQIRb4RmiHJ0w5d0J5LgcF3xQPWuigQJcIX7S38G
4bmS5xPFzkDAEPwGmer99Ng+4k3hpeooWF0mY5EgiFNghIbQKqUPOJ7belAIq6NJ
SxzioymIflxSBpEp03p6vOpXrrKmHAkBAG9jLSclo3jfrDyxZxmR/qc25KwjS4o7
UX9x5g/8k9EPZ4Q9hAIizVhG1MeTRpU0zY8coJDRf63DBLJS1xj2ULuUQeIQtPkG
FNukcYc4Z+kxlgmITRQE5UZX2LxDH05H9g9VBS0ugJ+naz9heEiLg0ZDhOLyTL03
6fZR8ODYmRP9RFEsDxYB0ZTKb86CdPHV+6LarOT1nFkOMCzdVRjtU7S+AUlmy7oi
wpy3jiBLBBWjIlSkA8GCUm7IGC9ZEFtXZrshTN1RucwUW11TA9ZpqMggK4xahGbM
cD7BhepmUEbqVkxCbYt+KRn3tJk6ear4itq8QNPMnVWlRG0zQ+kYVQAc0o9aGi1+
ItlGGN/eTVGF+uvCxayeE7lo70OU3I9xixA+6iiqfO2jODgVyXrGefmHWmvCIHoN
6v32bTIjwUT8SNnfeqwXvrG7HPqKIiUNgWJChxf5cgzCL2SjGgyOJm0HrSjj5mK3
j2MW/5jWUoO2JXTu5CJNIixd4ZP5JZPZkyXtiujGOybLcM69vDB1TeB8NUq1WjLu
upfbxho6ZWirZW6BP842dVi90WQiC9MNUV/g24EVd62mazjL08pl8FnrMYIm50yY
L86LQ4JOPqfAtD6yaZwRAJvW1COJRrx2rFqt4I/JHdmQ/FEMdJKWlh3YKaKvITjv
Qd4UayidYMHtWrRadMlKbEFuXsJjf59ivlu3uEX4KCrcXowccBlLwyy8Wjjnak4K
sdX+fsYR3+/nuWYQ0bV5hZ5nCmhptWnbccwduSeeql7dUmrUGl9QRlJZy8Se1Pca
2WV748cvzTn97AAYlrzkpnBsE8XzF/eSqAux44YjotboB1lE/EiMPlNyk/mDr4cm
X4WcY1TaSKYKd6d0UgNT101i60kf8UKs4KGWvhRjhIM5yaxG8piPoswDvBDVT0FN
HRqLQHiZr8IMXYldnuIPvRrXuKg5keAM3c4X8bt6Z/f8uDpOh0Ylx1ni7D6h3wg3
iCKQmtQt0AGxi4xbxOgxCNvhCYIFdgYU1CSXfMwOSaNez9w2+LWXp8Ev/4E52wO/
KCk7y6vIwehLyimXnmtefHtuLNIEmdoAZJYX28uVP7JDJv3a9j1C8bQYSONo5egY
twS+SvA56sEpfc8aR7p8vMYPW63QUqv1dE0EGFicq+H1oIZGjs2+1uH/9aH11n0R
WR5gzcRFxEy/TQnv6+chmRpAp3jAGev6qzgt2HOSNzxqWbI14Kfa3WssIpFkUE/C
CJsMKLuFRLxV6+4BXNH2Obc4HxMrHxm+rzfvWWk5WzWOsgcDDB+wDqUUf3yQwOIt
PqQBZxZazMiChd0VzkVCqHIQF4z7LscTDdCkeIlRtb3i9OnfG2wlIekgd0iAVSGk
J/EUUUTPHMBazZYUnWPw+xMrrgBcYkr7+QlxObEYUUz0FCbNONgOGLS6WstaJS15
NdT8n7kCKjM243vaayj/I1GUQ3FKXypfRsZSegSjZQJWexR/Zy/bRmAu4mXS/eK3
bBTomk3XFyASfE9JmUxB+RKq5alOPEg6wKVJSCuZWZb0i+QR4sgbmWJSf5QnQX3x
k4frk9f6UlacFUx8wMT/4tJbYhtgmLyRTMd6kp+qf3S8+zu7XvsQBGjt0flDePuz
bolBqzAD/KNIpy4QHmQr1tYxpeYG8YCPaCIDDQzYvUpKC5yiQoLOk//vXU7Oxs14
vUDmxxC7NoPsO9HzpT2o3JQkEYzLtW0/lMbTTJ3HoTPLgS8mPouIoVWfCNs3WOln
9iVC6iKWqjGbw9dBCFKrBN5YeAeS7Z2AV+spTf01fF6HWiAtjQbN2R7rT8EpCRAW
JKsgmqU0Dpk34MDJjrfoeJQ7RITH6zVxRUyoCHtzGxmAqSBINJvuj0j8acQREFMc
xEsifNzjh1XfYWUGfbVsXAoaA0pBCGRHJ8WnA1nk7c4bbpEVS2ODspP3do4rRuwD
WRupoBIIarFS6wJwB9hq6bnCz4q0X2B0aKja3i8nLUY8tXW1RA5MpfViX3etl6Lf
gptKzD30sByPqJemmgdphuJwYurfMSzF8f1zXG8vt/wJ/BCUnuv1pJYJtWe2mW5y
KY/Chay66iw4cLLgiebM21nNqANQ7bHb8rOdt0PAHxtN63fajrbFw8JEatSrL4QS
uXXX9j7XnqVowd2F37vmQCfsV2K+LDU8wXZom4oUyKXDIS7bFWhkABctBHZjOvB5
7XaVnRTMBsyqgbu7Ca0R2ECXR64U/9sVBp8YeI3jrsUAlYDt8QClYzNCWbTntNh8
fmxOyfjNU+zcDA1deJSb+CCNM/lCxIFATfBlXoOTxqIQ4ctbzwrIaKVdgvUWSumu
V8Ydr40q6ua0fhKUR/qrwE1igDiAq4yUAW6fYzK5ES1npt49ogZd0lLxmzpOceP0
tGmkfGM4o24AmmYXvUbqC6nRB1v2T/G4i4SRz23oq/ZI/aSOuERENdxxh5bC5JCY
OHgwAd2FuFsnySL49DOV/xumnI0j24zB9l/RNKF2mENfrIE4cLXwMBZ49NWF/uyA
wVp3qEa+P9Qd/jvibNR0t6UXvQH6gInNxYgCb2m2VTZgDKfw9ZNujc8eJNxdJ1oX
4WSRl5vItTqotz78KZzGASiH8spPmDb8cWulAPhKmQWk155jbMkgy9Nz9udltXKL
DRegtrjDtA1+vlTekUbAwFHTYN7ymSY8E7Zmxx48sQlRYnZNELFPlZVycLUfa6C3
L24m5x0mNz7VOUyhJYwuQtQRLkGdHs1BJcS5VtC7Zvrv1omghH8ifCk8SOJ+xjYZ
Lv4F4ZRK28LlSwfkd8SVF0NhSQ0F4NCZ19NXYwVb8rdZOBHPAMkwDJTIQsdPJo08
omEtOuWxM7ykOwEU9eys6C5ElvYgQIWV4HrqGzgqfxmTe3V6zUCbmtq7f0vepOJ2
gZ3ijHvcip22E5baNF3ypSIPyMcgUYjKHiDYleUemErEoEqdZhUPdv35jYkjOdYk
8BSgeyA8UHWasBVnXqfV7pou+BJeVwBPq/Sx/KV4IihKMchgIMs+PrE0Tx9PokLt
M1/Xy8Nd8FSKmE9xVpHjrv1UU0KFK/oA+mtbwmOQyU6O4PNpLWjJH5wkiyq3Xxwx
WsQR3FQajghH5MI8LQZczgjYJOg1g9SCgc9BO0thB/8fSxcTgc5lS5Unl8aBvxBB
N/vvPwSF83UYilJG8HcagRGboPqflxS4nsTOQXDg5kUjbKhFiBHfEWZ9PMz68sC8
Qh8nUzPLFth2IlQjg0Wv5PDGvZ2MZXX+Dmle0hvOQxJ/1ql/W9Y5qVfvMcGhBtNV
W8zBMVNq5/a9fOy0WCT6OOpQT6J+5up9QIS74ZtWkdNC0UL6TUchxHiKfb/vpWyQ
HY1+ySx7F53ko5KlwN7mmf0GxdS7MQRIK2o94rSp2YA4vX9Kfm1wisH6j00ggsdZ
RWTRI+v2dnO62qo41OltbrFDdO1H5cu98Dbx0/yO7Ri5KcT26ZfCuf0egfyQxEOn
u9e3+rvjX7V/WTQijGPUAExWX29Zd0tXe8hTNLLIFS17psFy7nURmz/VpTKMT1tv
il1pGbwcb45ZJC4aqqbiaUw3Cmz1x6+6cgeFR0gaabZU+REaMgkN9oRDh1CmdOFm
bkUlwvylNVNEkOh7gO1y6G8qawbZ0iAlCJK2IR07qGvuvLIpSmysq/ETEb7336T3
Z9m9DpxvDylXLOtm0UIidSgGnrXG25QgtHqFr7T+9f3W585hTC7S6A9X+wwP/KcU
d3Gj9Dq+x9AJlrTOtIhHKNz0IjBHFSVt74uaG1pU8qksdKq+qYsdrU0zh5pOBQJf
Ldv0daMDwBH+0gKt+yB7ScR7by/dyd5DdIUiG5mSeyE9L8u7CAZSTulqGGQA97yr
r7gRf8OzxqJL8PsmKHBZ6gwYD8Pg4TF5cvFnkCRg64gKKS0J36t4UhLp1SgU0qFW
t6UdA3Lo2EJy6h60gzjkMNQPcaIJP1HtsPp7vT9GIAz2+QLpGcCsjkvfL6531r9c
d1PovidXjgjg1ONYEfTtoBWPXFJKWgfCA4ElPdPd5Jn5QFGCV/cPh1EvAa/MrLjt
2mzfsUpDysgsEna06MChDmWkpdaDsmsM20UHSNBwqzoBypJi60feUUHu2kRepISP
SU3kFpSu0a7XjTgUZLQi8zOQMUq4DJK+kHd7tyXXTU71BuRm9J17OofV6yakHTF7
U1MZOPvk1S2hthgxas7YSO3DDBdTtTxb22TGpYvR+Xfjh2s38ewJuLp/YJfYtnYe
EFfVV6RcIpd9oAMzqH/mVOapmU4h1RFq0DgFD//gLZgIT0l06hXZMxxR7+47sjV1
GjjhY0V63PD9f95BwggiLUsPOqj3It5rMsZnBjfNYv/KZIi+71zF95WM3RaOvRXn
645rBBULiF52EVxBygMcJvVUZFkcYM8wJMbd2+fztiq1g47YvzGHkT77wof23akh
IaMAIgV1rO1Ekbd88P97TMA9EVx25/4LdK12ex0KNL6iWYr4Eo4W9CucdbL023l2
YaUoNp2DpX2HAWsLfh2hwywfXubSaCyZCyQ24ynoBdQOfvNGUy1PfgJ7j3zNveXV
twa9xiMeAJyn402BJQwY7AW1MAs772t0Vqi4kLVX/mo7uNh7NmSTWLLEE7e2bC/j
TwvHRTSEGJu5KhNn3pO59cZ1NMw9YDKGwFByURiCyY9uJrCXObswF0ghdiKktu4i
YKkFWHe0BZITQzlpAE2owhBTIGY+QSbQhhU2jgsyXAGmN1akqC78Jl66wTDZG3XP
004jSVBzwG7DilkmX8lZ9UKqE0gCS02JKNu9yfmqJ3xDGcLw/R0waDptkmQABJMp
dK3Q7kOM55nTg2tHnjSGVl2vbjNtI/44Y8EgJNTCjXeweUmo39DKOFyfQgYjxojE
LvGs4Bc+yiqun8enRGJQUVUr3yoEIlMj9jpQMqRxw5/8ksi9NSfQe96lEC74vVNd
np4Ff4kF3sgla2hfXiEr3RwMrPp8j/m9Qv3LLlHTzgjpnghBm88Gmi3Y4exj/c4k
V4EEsrDrrqIjk75C7nFHYvm9JnpNsaBkKprr7ftUozB98uNttd+LD4UYmbFWYHJV
FFOhSI2qGbMktdvOZm/IDWMT44qqyhfJ7K1hD/NcrLFtTevxMakFWgU4q+V6aP2N
SxMH1FJ9b6utjiPRiaqf3rqCrWWR8/VQK57WtK1yAEZ/d3eQZbr4532Zc0NT3dYg
pq01gh5wHz8hu8uThuGd5odJyiD0j8U68ej2ATPrIl1XCwPoN2siWkQT/zU8LEng
GUdLp/G0juVoNE6z4eX4vSJgWNfUfuxff2hxsIf92n644//hiHe0jwrSt6qdOAFW
OI4PmA+3n2X4KVHTz5HjBoT5tDnd5jaHhhkFS1CqTMaZNmnjfmlYEmpEzf9f4WV2
lFn94nYqz62x4ihgp6xbapfxKLOuO8ZHP0QUUWsQLo0SF/jPc5WarKmvjKanPsbl
adqtUXA5+bLjSx91q867WNSo+zn3TnSkod6NwEGbkCZmzt2ZgZVnArw9HKfAC1nC
u7HB2Pnco9LnrK9B2fHh0r/bPZnk10Bm3FhIsJEuuhaJq3js2/NqWS+GorOOqhpy
1920P6FolbLwq8sTOfVfQ9ZmainCfo2/7uudPmWaLn9gvWoKHLoc5yZA/Gzcwdiu
7htmi/q87/UBGFIs5lmAQwBvI28flvm8MMmvZz9UCJegsfjmXK3Yp5B86Gca0q2b
FnghgKbUoAZ1jkHd/xXu2H2cFuUW0doeYUi6gJFbs3BNWW8y5LwHJCl2ZoiQ5VEO
Oopx3FBsoRVQAXYStnj8kehURePKAYOgEegc2VabvRHsLk84/XOPJ9kUFoLNLj3n
h+rK9dfac0n0F1ixv4vSNYBdcCKdsbS6BOx9P23CYYapHYw99oCvQ3REhGOEx1O3
l393llPgAzq0NEPTZdOFY6fw9JbPu+aGgP4DqJhX9k/lq8qDikJlXOKLIHRSURoP
Wbs9zJgrW5oNrXUzuK6WlpZkJryVO9TclWPu+YpZABzttqKAca6fltQpyV96rOvF
JaXYgOso/jSqj/JTu5hTFi5N943sj0UV20xvax6cyFVM5mLcU0JNdzCF6U0virQp
smiAKPe2G7Iioybb9O+ibJz60Ia0oeMDYhXqXKTtPZaTj20atrpjHWbZuaVT8izs
yBLeOySs+ncqB6ETL45PYm6/7tJ3rUmSlQhHrqeb6KSqN5oCdY5B/jZVp4z6z35x
0LBq3jYJM9X+WWuxktqAVb3fHIx3c19oxWa4BRzsAvi0vkjyqcFfYIfLRJZi+CdY
FILaVz8dX4MG2pvfrLh2HpOucCIBSK+eX91+7P2qSuKBUd76/FGcIvVEqa6Zx3MG
BJG7SPf5m1kSO15uaNmGRwpESbTRoktwTBb6dLyNfzOUNLWjW2pzL456/od1gfxl
ffeI9o3xcYX9u49jLjUgJqUBGKTTOpQvfOIIRWwmz2Vxyz28Pt41WjHVfZOYEahR
nC4+6kPLbfQoJQeVtuY9VP7xEeCu5AyVNw2z0F4fnjt8VhUKj8iyuJi+WJfC/Zgm
mcYOsVwR5y3eQmCSZNLKIgJiWsyLcbfCTD4p9d3SXriJU4LPYuPyX5z+knPu6rpZ
mQeZn3XLqa91swjSQrolh4eqM0UFBORQ0DYFvVLBhH2maOZNEbWqXV6wLdSO8Cw0
LUO/lw0CcvXN2xm9CuVUVQ+o/rfnNW1XiIC9DWr0aUflwPHLcG7FhiJ1U/TTAFe1
P6/uBENS+E7prlAq8t2PviBZhDxVcshtqCzpuHmxPMkj4mYjzXGAFvt3k92tfqNn
gYfaboR4OtW5Tz7Z39Q8r91VjZVkMwSMzlRbH9hlAObVAEQCvSffgr6Rhc51JK/S
QofaECRfUjLzo8IT2mc0FtdW0ErAJ8D4gfjm2rFbxUTZxFm9ErymgxIJIbZbgqfv
+g72MTI9BjbHxNc7VaN6YN7IvtjswnMy+dxfKbHRYVizSL8PQ+8Auf3tjFMyFOx9
M1FfcFd1gpH0Mg3bIMFijg/qvL7Aks/WDR2gh4bgjPo1lwG3kvCpngOSn1enWfm6
XkiHfN1IDFwWH6y1bWv89mnxwxr/UFPgzzsQdmCIMM6KjB7kIIEc5ONY4qLst0o6
QzcpLvD8bnL0jJjVfBYmNwBwwgP0kaU3yzhFF39yjJ06zy+6fapEpxwgSfdCntZq
CqCBGP455UYT03svD00FHttst/rqpyizKae6lw2b3Q9/O/I1cshTprbda0aUucbH
cRDBSD2ZKEykdWP2n9hZkONKC6/8l1ofD5R+AJnI1R2ky4cCEqCJhQA8him/ee02
QBb3zNCvPDmHIKbAhbTNUfvtv7DYNDD5/phlck84sfzY/Bz8r3eiDONLoogyVPUQ
8dncQdsx0MUkDTi3NLRpKmcFekazKWYCnvVOqhjP8zJVH62Vf+NTRvcDlWnNEEYV
bAlJodOYOaZ06GAjbpL4SsX/afNy73tbxyEvMzrtN/TrB11rHHZF+oIyXmfDJCSe
gZwDht+sEGIg+1zUiT9bDZ2WUGTQcL+0bj0ZL8eyO2/uq4ssl6WzB3II8N8OMqNL
eSdfn3rtKyF1JVviw+fGY2STMVUb+qfpNnDEk3nd0x1gzwB9Lp6+DYNVC/0wRS2q
Mn56l9EtLDPJRLgDBsLYX57BcECgAuylbnuKjcZTwZlMW2sfQnkDdW0tJ2D4XGxv
Xt9Gu3AdGliKTVkc3HiG8Uy0Dopv0t0YAcRZFORp7+paCE5lKsH+PtdY7fEEzRes
UYERbVwqTwVBcHnJjNJfjiplEhRlH0M13psg4csAKprCzVLYcoEGyDK17eVJ8wAg
sjZx/Fh2lRdCNYA+SF8mTBHAL27Ynn06sKy83L1CowVzNzcaTlvIEiL/Q5QtxoYm
QEfDgKGkFaIuXlnSZyjFeAw1UUxhVU3FfZO4sdfbE38Flcx+yscUq05Ln4fvS+ja
W69P/BTzKGFHLnemymkp8ixVp+TkcFAPfVCJPy6HuwMdGQkU51YYeJWTZd5wzhW6
J/kPgSNXThSF/Hv3lVLGcs+MzAF+FPzaw3Z24M/iErjhYjD7HNHTuCogj3+oD3Ch
CgrNtn3A+xh0vyt0GwzDSguyhULShhgj4gH9EyG/qafeF+/fAuj7DJDgwLVV6OST
QSEZXlwfDEuivYj8CmPSjbbfzM5mIr1oWHWomZloXad2Rj7qZuC48ydYY8dywC61
wER7zO2TXf5L5qJGmuk/o52XEitpdl371cRDkuyePpUeFn4DonmgaHgNUSK/HDrY
yOh08wi1GTDORnV8gxSVbKIM7iB16RwnUGKKIUQzXgWjeetaet1wFd5kdIjFj8y/
b+euytN7/05utx9VIrndaEBHn8Rkf/s3tcnrRogn8fAeUcjm64Qdmpx3/GJx3oFn
r4ApepIfU5viu0GJ8hQTNcZbJ95Z5KFJNjoDqfyzrxoFiBzUkhRmwzOnhRKLjEkN
Um6STd1OA/j4AR5nVvcMQODXUCmA2Qtnz7Lnlkt2+8lmT5/DB/SUafCZI3vZNi8W
69tL/ld5Ji7FK37lHQSB4jL9kB7yT2Pcjz9A2yXmEzYbh2lu0uo38A7Kfh/tAsmi
uU4VQoSjlCN9KoI4pGp2hw7KD/tOFxpj/hujHK4N4QsUNBMkvSqNJ8aYKVf6Smlk
M2i/ikGvkSat53ZzPsiWD72XWddKrD0BhHnbQFbBrA4P/W59LefUgqn0kq/L9qPk
wUA7lEGq9lQjK3iX8OuMPPlt4AYPgTzoeYCQifdY4htpb5NPCFkksJs0FkJBwEkU
lkn9L2rZYW3QhEobgKxMUXyt7hFMQ2Y4GMdIajl6RKFTMzOr3WAKe8OphrbBwPqQ
PsCeWGOKeiGva6kVr1Zzz/K6xwTrtSTX4jbVxVNaO/cTwTHO+hP8HG3GdXuKQ5g1
M/GiolVMnmhe09R4yM7fKrf6tjLZ4bpN1T48LeOAynehbrt+rB/oPeIqbxnKbqto
upVcc0eg2oyAep0KUP8JhnhIaVHD8Jj4of1mFxHIiYJR6QAhFlatPoeIiiniL8FP
dDHTn9yvYUxAaI0tH+yjEOM0Wp5OmFCaqxDRJjAii7vq0zSbrOZ3bgRObGx0yA5O
gY3tUT3tOqX0N9tbInFs1sK37WtcWySWF0uK7yCptqAw9naqH5p5iRRDvm76HLK8
uM221UL8CpaUegaC8JlZyC1UpBlKkIFn5BQKHvldhbL1q/vDq/cs6saB+VbOEVcf
hiMe9TYtLns1+OSQIXRV/cRY+RNZ9ONvQmpQVuLxZ5lVLAU/8LCoAcb9bjcz1vri
+3hYkWfF1tJTMfTMrXvkCDOMO0mV8qdW7wYlHkQAzgQodjspG81C2XjaX4rmQ6c/
JXvA0kprE1m7wjdHFizOLSHSFff2hypFT4vzLQmEdlmnYYAdhnwh+1+rqQZxcF2D
Y69rdiL+QUvtv/6c3ZFqp/DHUJ9nZFOB3FR1rhUKaRsHkmhgrif5ypjl8OZCQZ/h
nlg7wsbiSCeFoadRTzJm7T9lu0uZP+eJFcSw0+A51IhL+JCr43KJjtdWczlacOLy
yIXjazFCCg0TqdjHFSGFSXuHjzICX9NPL0Ur3e1AOFzP5hzRyGBrPXsDnqd2BtpV
sBsMA0tdc3JCyiPLrUZ7ajViNucmFICOcyZy8vRkU3N3i+2lodQFnh2wejXKDpI2
WKvtvWm7IaOaRbca+oLj5HCsEgtzKmCQ8HzP0T/5RsC5ZCp0G8LYcc8WC+2t2geu
tlDxlcl/I72BqnVLk1B7j41bq0s6ScvHHnpt3Bm5VgjABTKJVIqj+tyiVnTv9aB/
sGCa8JLqsLerAO8fX+z46suS7YSZHnKjPVkZ+YdlQkpzRpSHN3W4UlEAOtfj1eN4
S/ErrRrXiBQosCTILfKDHiHqGV0vdV98G/urMvwMUvmpH/lSdzTVDfs1EODhNK00
uzkQauFQAQodHdtLdblaDnTi+f3T0tBIS4Upp52aBMvyim2A08DgAFgbb6WC9EJL
iOo8/hzJjfBPmEqjt+C23EJrS3Kivi9EWsTSgmqZuCf7pahntrzQwOtuaWTPB9B7
40qx+9GM3ORX8co0kQTkocIYsSey674pqCxR3vtuvLV/H5kl6SNns/sDVOJQtKiG
K24XkEtfs43ufTdsk61pDGFwvKRD18SphQwCat3ts+H3KTV4ml8Qq9BBguSyQXCd
bMVS8cb0luu9YkdCxsxFpUNy6y4KaplSSK68K/70OlA+BYUkMVhUzQsoHtg6FaBg
q1DXL1UkosvmQR6z/BFUtttrW82nBfubd2jt4CKv/HrF+kTHTMwbCH1fRdOWjnmf
ZwRT0fzt+GNhBOaH21gUL9FuS6yLdv8nJTuoWBL7XtX3/TAO7s0QwBXfiqBzGf1t
9jnSPsA+3JnbxSeLBlPbus+A8/vW7a7MDaQcRQjlnXPAD48VYhir8BBMVjrB4I2r
QfdGvAkdtEFb1068V7wxqUn2P2vP5ahDxkzSie5vf4C4q7hNsx66cAkf9xZgK8sk
uQUaHE0glFGJMqaUd+x5ZRV6mn8Y/JF5CV3OMFnJvuppWvT9lwj2QqT5EmMgVBel
ct0aN9pOFk/r++GS0kdMxEqEPozQrHn7od0BQzy2KO83bIrvtQMB+cMRCbWelwXF
eut6RtoDSoxJbc8bw2nnmn8Tw3BBkQN5AzBiMmxcyVP+SViLipg48U8nde5PUq3c
CVgWmeGHbvZjDQj2FofN7/sDP4JzW0vG+Ok9mqo8kurEpmSTqlpMCK6zvseZy80X
WYolQqc3pP5hBi4fJI8zYRtG9qdI3qSM76GucttyWDhR4vvz2+MNydFVsgxCFURK
tzyv3gscfwAiTkYSIoogSuJsAexQ5Ty8fxUy12t+0vNEUNIlrGuBHgfOlxpUVzQj
U0w6eKMlFmjw9zuQ1+nC3WqPEOfaTFr8xNqOnfD806bMq4FrC5QAbIQN8zcX6Oa8
sbBwXgJT5NLPws++E1o6aiBhs+w8NjPCnVJPBMZ01o/9Xs5cp/II19L5WENdGcA1
n6Q26HtZcFrNJIRPZR5hnEU4GVTTtVnUPVAI15XVo6xLMSpyOET0Q10lb58vXJLE
psZSSkJQO43XdJevDzCH/h1RyPO8Q0THnDJvxgoWMd2CAogFYWNHDSJj1oe9z+t2
vhei5v9NG/xlf3qe8TEhk/REwsGO9pwKqDaeY3rmmefbsuG790IQPSDz+BFTOnhH
UqEQj29LwLLb1yUO9D0T9bbji/B3TfUXuOXlmnie9yEH5AXvMe112EntpqF5faHm
9ItKXa+FezEnWeHw3GVhbQr43Z9TVuJ2g2+bcY/FVzAQfvP2ZqsxfYpvDx3xXMht
QLjQEgTAgtGlo9YmFQffvh/TttkRZlf04fNGmBFGChFK8syz4Mh1MvQQYj6BYAG9
yWDfdvoAH6RDq3yVeIV4gMQD0K0OW3uIcsHp5sfeKvO328Ytbzwr0fLn3VoItY6X
2eOIwNok0HN5vxUH3E40qjNwvSgkw5XDWC0wMO7S1L3C7KhNHzxpwrl//Cr9YFlp
XSZtZAAPw+rmMn09j3bH6l0n6hgkAQhqAvqWfz/0jgkDCPQDUlSiJi2UigtsQBEl
/EwGd4JpMYMqpbFngkTg/J08SXlAuzryTHCQD7AgQj7FDrWMZSHPsn0V0dwCVXD4
6pLO4urAkvpEZEYoG5qrVCags0BSGF0Fk7LXWhPgepEfPLq4HBhBJ6vwEQPR4Vvg
NmYQGdvX+DZFCAACC6yCIAzEb7qVH64WUh2LrcY618iQxf3A5a/j27cmS44zIk/j
R14CCuOMFHxscfWI9q1XAgXL7hsGhSgq8QOmnh8kT7qKdZJoErAEuHbfWyq123P4
vw9xtWRMwZ5ZQ7yyqFBVpbP9tWtkOZ/gi/DA5wxXzcjn1W5oeQsFeQQ6NsKHDLPL
wtFae0d8dpBNvsDa+bxszLeTnfdZmoyNZeUtSDVh9jOMvAv9HE312gYiL745cmiJ
3txPqJmLGSQkwgLRvikCq2vzz4YNQCPhPb3wkqZupQl8Fc5yt48Ijx+YDzBPTx7M
lnbx4WEBVAUp0IEEZCB2qpBOQb/ecUeHIKs7J7dNH85yteyiHNqP7S6QbOigjqLy
cWgNSGNiXORfD5FoipJ/M6XgMj5s5SpxOLrF+LPRfi5yu/ii0iJQIt3GsAinv3Vj
F9A8156LS/LN2HwBj9oVFdL7POsbivN5tT2iU+rS+aF1ouc+pDvjwbB9oonJd9GM
faHP23v1UpWuXzV00BZgi3r9MQq7Xa7uOEUkZbLqaAV8Iil4BOXVBv/fGRu/qU0x
0o7C9TC0PrS9dZQ69Ssr3hMc+O/yH1TY8hlq9qwulA8QyHW7DPLl9CkeTYY6SBN4
XYocldYQOXgs0M9WqkMNLnDg7LUVhaUB49F2+t6QfpOnVXCGbtrWv2M0uXfeIEjR
sQbALlYrzkUCKRAgEgpxWMrZeAbWYe7j/NfLqE8Lo6uhn7MJPT/rxMdtt99jYw7p
tlEHfNJ/e28bLbKeXOXBWGMaIHA+fL9IoM5JnrRfRaN1c15wqJR/qCAvgaYD8AO0
RzPaE+Dpc2pcwA3Yj4lXMHkUNpMVLQnnhSY9Av++pJuvZnJ8iZukePZtKzWDw+ED
UeMime4775HjHnN0rZy8qQpBXoeCJQzUwnvGsmIL9bK4QSadQQnCmoWfhxEK1kEw
/3M5Mek/fanIRsMfCxLynb39icqM7eYPmFyB/0e2y3pfopprzN/X4hLfQeVSymby
OMUOxl62DI23Z5UPJn46sSJUJYKlq2Xcunz1ImJkjjLij1AzlKbQQUH40iAAWCe3
D69eQq3nVFwIU9mklD335gDejFjePmxAWGFmHQ1wP0lQgXZCHUGmtWwK0iCo8eYA
sw9uIoKTFJJNrKS79aJmtLrFXy8UQeDQWv4X1XxPQSoQoUzz3Tyqytbmz2yZftNP
zVBQXmOu56z1d+LEorElMhRqf3ntWgMuvhlG+YXRoE0NtT7mPOsTjmRPj3mRcuDd
V+BFLmlFg0LcFsV9cfqvz6JL7e2gl/2b0T1WBCWwq4bA4FyxZ0iKzj2JTLUqmaIk
ftdjnNe1+sXKznypNqlBs247bvhy5tBsPL9qi4+kecBURj52olQEbrdIfXWeKrWA
t65YkyEafZADSdn8Oydw6hQWyqtum4BlxUqLmDVcxqOQ952W5OU58PmBs52V9UEP
XY3aXGy38wKASlbfu7YRcTA9Yeg7J5IEjlo5tFLA7i9TxV6AAWFaWQpME1QNP8mA
udN48Edt4+0bQiaAqiVX1Z38xhVNBfPY4oXvhTMeHAWpqmx2wagjrLjwrrE3aBLH
jmcBLhDaHj1aF2bomR6VxvYsAHnm/a/hilwYiaysChBJULaFEJRA9yVpHYSNC/d3
p56bXIPAkubwj8k3OZOFIE2WylUts0hSxZl4Eo81+5IfA1r2KXdi3YBfy6wrLrE3
48fk3LMn2RyLpBhIKhBy6z2OFx8KMcRVXWSYIwlarTt5XSAjbmGkuEbgh5hA07Cu
HzEa+oMkcESwnkjMsuts1lK3qyez4dbdO00dtlvetl5zI0VRqh4v19lT8wB/e3ka
2ikBCUy7sLJJO3W64NqA2uajdOZ6w4y+81wC5UFI5Gv5o0QDpSIbLry3GarcOStV
WMyX/UVevPOkytb7KOCgnvcroCKwiYYhDxtoGjAcfFiQT9KmBCDj6EicLqKGpGyJ
dYbwaXTGXuKPLqaKHMAvquLXNC/6u6IVm07WLKR0nIKMGXs/yiOp7z3fyvVhQCBu
/gyA3olGG8qayrrDfhaQCs7ANSYjjSBPpvC737daLaMZ7Aj62jy2jk+zdIgtivaZ
CawvrCfBAeoG4YXCaZmqr1P8oVDpqqSBGOoQc7FYPBcdX+uW94PWecA85Ooiv+gg
NTErlKEX2kz9M4Gf66xc6fK9ebVH6aqdjZ1pkk46cMMFjHrh4l6dkExfs7XKUf5L
5fnxzSZOTO+iCjgNfAplUGWG3843IEwmbwY92PkcbEepeV4LSjDaw3/Ua0lt9c2U
mZ2Isv/I5TFfl768PadSa7Mg0urt/cgYQ9waCjcOa7yhjOcywwRFgS7cdMhtbVYi
1Bv7Bi9SHtrM8Xv+1W1oCcd2x+ciPO4AcYFaiWzTfvkqnnDuDDcK0hJ5BuLuGXKo
6eh3zGN/6gSaUoqPKjVYYGsKTJ/xAxgapbgYoxjVjR7c6/Io5Yy2R/oRCWNyI3Gx
ABRtjF2oyyp09aPZAJnAwIbbJ9HgIYlJ/DW4vIa5te4SRfltRw5Regh/RFCanX4B
s5sOzShxcKtJ9D6gaRLw/YdlT6drR8CN+J8gtEhZMHNxv6jDbRZgeNqqBow927Wf
umYGQdsPwB5GW/vCY7hg662HLtNNVK6yfXRbQx+invNfZ4VnAdDXC5posSC9bmpP
EWeG97OkWYxhOeRp1P0P1Q3K4zja8M6cmUH/F71n9oMMFd3nBn3b6yTYAT2dd814
PmNzebyR3Y8Kv1/PbIx8qfTfgvt36NSBJm3D/cuaxXX3uA37uiDGABV9jv9rk2hz
QvP6iikWrZ3+OsJmRNErXGfxPAj5XyWsuqDIqCpxWEWjdEeN+pm8h/h5qmc2lEBX
NBLLsWGaKBafL3H63eXDvYMv/306D183U7mhCSaQ+SVItqeE6HwcsuMvf/64WUbv
h6ibUzWL0d+duvUZ9iOkD8XDEPTtbMUJHg17GPm3dsXFy+9mutGhNgpTayKBvmKV
qdSxCmI86T5jO0K+Y09eVXmjaxNbd8S712leSGqR6YbOd/rggX79Pl88j167GEf+
UNR6xTjhxBYWK1IQIAyI53iFOKKwVAae5lPQ8XCwA8xpmyCz86k0E8+cDhNeFsvH
MDI+e/PERL+ZsJt1VgRLVsQbOIoGyqRv7V/7k3mHGEyaxxxniFuNztIsVhGCQG/l
wQ1erEbJdvWluXA8Q/Hj5S571CcTk0r6zrMVy/fK0MZR4ttKpruIW3GPAzU8sj41
g5D1/P93i/4uRiqeOdgkAC4kVIgQ/YqiP1A2vQ2DwmR/sVy3/ri+kmLaK/xfB9E8
nONJ0W3qk+NWnFWYhUuYVXF1Y68sx9CuKYVI3EkZ+eOyGUeR/SfK8nzvyNZRuW2R
PdBjYEfSzc4YmnYs4lcScnBfK0nNvITau+f8o1z2a7Elpw5K0xNcuyiGWBArdMtV
n/7Y8SuRVE5F/+Nhar1rG9Pl4FPDwXehQgn5QRQTMKIWBn4ZdMm0kRxlHyY73s3a
atR3B5eGfW5T7znGgmwcyyX/aK9Fwc/z5WwESYRYf7Bu4FsL4zMi3NEKy57Mnk23
03OWjTY30KnDsf50tlsOxl797j/k1THAcylGAwOEbthmEWySPJdKSp/F1LY8Gche
PkZDuOp0LMsTUlECstb+lOMRxP9TqbYfy5LbNJjzOqRhAGquc+ooWR1BlFt4G5ny
ygaZm+V+njBMJbzNYh/pca3Hy9CmJ+6lxjEdTXgQ5uOXmETUbsWoL/m+S+MVF3uW
wL1J7I2pDJ+n7DjrXZ2mAYTcwqlux47zTRRdeYTRn5XtqrxjUISEPrUzHXHXFSCz
8vr4rMq5bEZAy2jjKcYelz2MSfbbxLERCj0ADrv+2hMh599ky9CNYuO40E6G7eTn
EL61e5ZFEjRMSqq7ODHEfLc3Rec7p+zMsYGo8f1dQRkS8c3yaArDM2m/jvnIeThp
RxrrQN+XCQ3Wyox2iBjnnIXfSUi/4VwXoSk3JSfROlZf7JlpBgdjtQ6+tm1MY2wY
3zcSAZTgPRi41ynKJ1HLmD/nykVBmKhBh75cS2tJ/IUMAIewXnYEyAX2fFMLIZd0
e5QO/7IQ5UXie6Ru0P51ENk5yM0tnFx1gbGIOmmUJ9c8c+fsD/vtDdlICUtYKBq2
y/nHmwWnbEY6u7zTeQ/DviYJuDJWaQJ8zMzqMJu8n6BifToLV1VxcPwtOXhGc+Ia
Uye9ylpjyPLbuiBYSH2Y2k3WdjKXbuK8pggmmmyh+wihqf9eJsinTOxB4EKbrQo6
zEh97EcAcx3mnrdWb/94y1gzTDOWUkAhlAuGYsWUsWRNNlMtcqBlBPEseRl0oTfj
Q2a36e0pAjZOV5jrhgWux1ZdgF3hatnM5CuNP7Uy1Jy0nBCZye9JV5H8GwG37c7H
u9OZyED7e0WmWjDrtTIBb9tCL/3Vqwo+esODcXOcxjO+x9beyBOW9QKHZp9NKWFe
NTE8cBrg+W9UmlJIV2u6g9r1QHnosT9rlmy6i6g4e3mJ6/8YIV6HH4aBgimRDzG5
af1hRF53KnaeQHOs3wP46eViZ/jRTMckJ+TYRtctYOIsskIdkl8DgoeqfEz7ZWFs
sfPtw4m3URvidImlxQaL5lSGTXbvhwDnIh+lTzHytFOWr7qNzDVT//2hoFGfAE1A
ZFn2rqq6/UhkxshmqiCF0iN7q1qvY+LQqs3gZ8Ye0wezLOlnqu7y+CvA1cTqcmes
wyIJVoLRpAiXVbA66x3lbLRPfLk2NM+KYp91jo81cETmKdOXjDf5468XfICljGxv
pg9uZOvHTPKzTz3BbpB5BfggFOUJXmEcF/54BvkdLpEbL9v31o6VxgrR9zGk6e7I
3H0XYba63w1MoJ71SHyV0HRTXiwKMEJEpy0MOCE7pTVWWE+eEYR7pXZshDp3nKsq
sqF3Y74R+woZAHEKbKX3l9ouBgmhGbBYbtO7v6CBYnPu37m68fuR8S5ivEd7eukG
qmVzHt/y1sFOVn31FJ4Yi0XIlRb3WYlGIkVKMKdLu+J2ZdqIHeRFb5/dKv2OhT5p
1R2oK6LK9KJQsjifPFUvnNy7bxFL94gHkSotggH4tVUfxPrn82RXbQua48PkS+13
cvFF7eh0hp3oRJCiaEOxyeL4um3HPRyo3Pu7v+I/TcAg4tLx3Q6YSdQ2+pXj7Gix
eC0t7LotnKQzggeh2Oef9ht47bBSeNKJYCm8PjiKLIuFV6oByZcsGN7AuBjMnsEJ
bv7jHVOuGb1++voGdr0N6L5oOsfl/7V19Jc/dalZK0OLO7HY2FpLfHwgPM6f5Et/
ZccESOT5H1d0i3JmzDro7yo2poVpNioOg9D8lpHP5r0bcmbY54+vSnlyM3hx627C
gLYZqXl+Um5t3QQ4QQLBjUj1vfer90Vz6BQsfQMrDD32tF8If/tHhGAob08047Rq
Ep/nXBcFs09gHAGLmJmpf6Q4tVV37d23QqiogmSIWGdGqIMf99We7l5ERpAJd6cW
OGXycJmPkrwDTsZMZyXeCjEDC/diTGhsqxBnUUOOlTpL1EWohX3DK4QOrObqPUhc
z5RqYDv98QJbu6Yd1jaNgvFFKB6wh4sx9j9ZYfzjOQ7jyzQlRLALLdrojtlnc3/z
VjdeltEgWILVQ1IieumjEGRBfVXOF4v/PtAEjqrNKZLQJ328X3i/DmHRkgqUOTgg
eC5grSHoFrT7kdmPmH2CyJ2Tna/V44YWFrVzqX6v255MCqj289Rpy4YlpyQYer9L
ZhwGiviFjIuarcR2YqRHVHdk2yoWobK+5t22dQhxBz92gbzMzqaGNjgvcaExoV+F
yYl6d60TleNH1UcLIKH5hB3WYhvsA4QuNlLnRazKmzHfpEMV/9a6JNrQPi29xTBl
XK50TyCS2zjoNrrTVV8HWi+gFw/ABussNRBYYuA1LaSZQnCEPBaDxAxlMF9h7DFo
u+POp36LJf42RP8jfNOrsahtfQ3vkCSowNN901sXVB7lpenzMaXG4Nuk+8Au7jbJ
g+D/jHWvfGle/0XSDthWnJaVv2KOHgyU9uCUUe1vkTxNIjmspH8wPMs5qpkVXcNE
picnaxC7Oclrg4aw9Cg0oXIqbhwAZd2zZynG+uKUx7YuD0Wv4T2vfHX5GXTne6Mv
hfbAjY4leZEpimxt6VBWYyM/hPhPEXLAX2YnLwItUpdXOOb1pNl8r56kGH7flkM0
4TsH4tq8nr9Ap8wzSms9UlAaVQkie+xpWzEEEP6PyaPeQgHze8D7xCV6PFvKQ9vG
m9F+la0bhLGlNH2Eniubxcu6ARbEEO47CHgH3XN9O6TaKh0Gz+SMkIF+8KknGeBl
umbJd4mJqrH342PnvNa8j4/IBLnZS7TJq/4FkInU84koUewaHX1kKLMSOxeQhMBe
1VQT3wNk8+/oz1s0vkk0fcJuopkrSR9NFeQtfeFd0hRxibjoqdFaPGdZJFppVI18
PdknflqqyQN07WsMpiY6R6KjtiIhul4nCA2uz6nA7RRLCJJuyMU+HvB4FiuMr5vT
49I4Uwpqb0S2JDs9ZDNYSPN6PUcksuiX/re8m88R5kwrYTQ/JHbSFrufL1OybSq+
Ph5CBUXPwKmuUnoh5n6zIo4JdzpGy9VRHtJ8PjSp4jZf4znCKL5HePiyWJnouxsT
uZl1B6Cps4Hnf5bu7DRfwgu1kKkIOCQT+6lyKetDU+l5D1YKGyDsF8lDshi3dYxQ
/y+a0QVfbdtKohfsBH68t8LuRf+c4fFNIpFGAcwHsd1BQf6OMERKGx94Nb5KU+na
qkPumYyJcmGsQ8QXvB16Rt3qUgnYtc9wCUuN0UQg1RyTmWWsZPlHTLCl07DhzcBi
rmXRFv3X1qHlU8NEzAoAcUYUfTp6eNTIMHomGYbMAezqSuhlytrtWBOvyYxHuGcD
4TIE72AsSFpnuj0e6yCivkjWrdFZDIySlkI3QA1rJm+YJvLF37c87wa0CTx7+0Fa
AVgYiLFoSWJfr5FJIAs+ww+PLNV167RuZFHie+Wt5Dm4ojxLnJxKnNPJ2AvTYE91
/zbMbKXZJeONDXtyYuz2o2ddajx9F67zw1GZaj05j9mVp4p+I3IeFCP0+KEW+Zir
G9g7aO63IYp0lj08UWGJ+UX7X80yakF08fRoB7btXI3FBuz4Pm7BTIGyLCRg714G
iC89pWqU6qkZ7LhGtUI4VY7DklLpaK4pV0KRzC//fCHpH97MAbwCQbF0L39W4Yyv
n04XCXrPKkdTzGkJmJhT/wfyNMnFwUwd1WCL27WRjN4McI1lmeomoKFMfzeW2WiM
vieUZUKuZQm9OSYyf4kHnUN1frv7pdkMZEFFjJaSw4htkoMO+u/TkZ4I6HrcAQhR
jBu64Rss5FrljatpajBPKzxLhBT7GhgT4wkajNDupNR+RcithL6O7zImVyBF3ApE
xb83veh7sqLDFCDk5oq93B3NHeT6q0sGhkC+6zeb1RDIugT+tPBYYWD5e18DXApn
t5qqHnWugFD6TSlMBsGn/cbFQqvdr8mR09La/AegMqOQcUlQ+r2nEfTH7vzl0DAu
S5Z0TQbQ+bFu9P1btCT5wNHTlfL+xRDNHkfMJK+4SeNF1tQPfUBSpQjIM4tkam8R
gAdCMFmbyd7OjjuXhjpvEKHGayU9lcyc4ThOh56kaeXEY+XM0Bxa32GugpWazyn2
L3rlpa76oF2WAlyXPi4lN/pkYDHtyV5XQlzNA8j9FwWmr6cnE3ADWTzNy3zZHimw
mvuylqRfvqbLsgGgVgg8SYugtWiLtQfR+1Cvl5Oqvz2ekVxuc5DE09Mz6rPgNloh
8DKLadyNwyCcq2GlPo4bzsW3uwt90EBND3Flf/3xJwxxpSxrGQja0l7y9zPqArzh
dHM4Ub6xmXvMWsHA39fQ+2gLw371aiTS9Gzz8oGnxKxkNUXr5Si5+WQVkFtnn3GQ
G1rD2m2kDE8lx9N6iOE3kAiieO5jkNuuswNXBgkhkE7ksUN3so4/Zd+JTUevBX6A
PTfbPuvkt31oyYBgCFl7jBM39X2h0XQgOPU4sy7Zm9GXbxKrdtFgc9M+ZafZqgts
Pc1DoPBngpNseR6JpMmO1alSMQ7msJzLP5Yvt89dc/+mBVnObHyXCxj1T2u1L8bm
z8lg1NvPXjtEb6+k9TMX1oILMLq8fLVmM1fzlcZEc0pZC6R6KXAsmc8lQL50tAjs
+mD2aZR7trOrqg0U8mKILGT/i/XTfxT3W+KwBTfgwYSgeGMbmPbFOJ1u0OYkSDbs
QI5pf3HUYNr+4ufR1clQXV72kLzGJQ2NLFnVUREnzCuBzxVQKEIQRAdWq4NAryfm
VWUuGO+jlF5r+cquglcr918nsy1vSjTuFZaJQ9Iwkf63L4lDtBR1Vurk4cJ3Yi/1
pQ/pMaXD2BDPAahxe5V6fxK/j7pMlqvrdt3GokRWm1EvqdQ7YbysFje2cBUvrlPy
t+z2TqqZLkFnQTdLBeoJXzbzJnqh162B4f4ExCApEN6NCeRdMPA6Nd3DMwCfnySI
iHh9rWRjIXjensIHKvbuadyW+5/L21sOlmtceT5UDD3kThU6T+6b48g99SFKuY5s
ubcIRGb9U0PGggQuKSmhgGUrlDWoBXxt0tOnS+zxt9//HZlR/nRuLPAHJs+znmPy
be0OrlIt/WJqIolaO6w39/7XCu5xgA0JL8JGHv5ZNfqfaM6tR+bdTFd0Lv54VGXU
GvH//jDAiC0c9zhElsb/TxW1mk6IoC8Nr/nwDM2A/b96qLt8W5qF6DOhKUJZGNqW
lQ8orpH9JOqKyt7r+OgZy02r7Unl56tYfQrg5v2s5Cq/hl7+3cEx3o02jjmVQiGA
ZcOpuOonmF7t475l26uINOASeIZA3iVQk59dfVqN33nkXRRumBkuL3wKAPgK93eG
h2NANXcJ455xvlSa+C79MOjsMNpQUlNYodV2IbmRq9Zm2H8yfXB3PjiEqPxvCaIK
y7eN4kxjjM42dYtVxN7zlmdm7x+tMa+j9WPlkeZqEKBXeoFKJUfq/zBEPTKvD50z
96jv/7KP9F9XP44uVRkHe4p8+i4GdyB3jYxQ4UnzfDn1+9TmBc7hBNU62eAuVlN8
QuF4/2OQ2A7h/JjR9OSFwK6Ru9enaTXwU5ZpWDbhXeUs0t0VgbyZy3HPQoZcqncK
zBF2pr/6kajwft8BR9dWQOMsozFxu3M1ugfR9RbtVg8anJpYgAzT6hvB0LNZNHaj
h7v6GFGp75rS3n9o3T3v4R0LspnoWIQMNLOUuDoGJSbsYCws0Vwx0qJ7+mcQO01i
NG1aoBBJ+DkGtJ+czVqrsTESdCMv4E+81kWuV7/vdtaTXmN7OLMCgGg4M7ITpJSv
HWBYGyeNm3k31rPcrd+LhDXUfKVjBmGj432kAkYaE+80Aygt57Mz6dqnGLzVwvX7
6oKzR9EOO0Z+yBJWIezPDPiMkTdMcklOzXUVhUUjTMBqL5BiVxRCujbYTRuM5+mG
SIb9/pEVUHYO+EXsdSTbzWa0MRiDqtGxlZ0Bwe1R4RBtnNQ0epdjc6rMkwbFTkZc
OZPaqR/K95C8KDsOinZ5zU7nFSY5Da+1KneZSpFmqcWTkQUwNTWOadex2UYx0QEG
kknqrqATKLouoDqaiDfULabP6FDU2lAJCdxbcOeBIm0EidXesxA1zLkMZLczIhOl
w3VihQbRdb6JHOqQ6FPV96qpjLPy7ZpOUN6oZqmKkQzH6XcA0H4gI6Xf0RWVSIPl
WyFcRF1bOMtBYQDwfX96N/9tcORUuWOrjMpoOs1EoHlIyLEltpKdp3uZhXKvhO8K
IYohjilb9DcGZplaIBGhSxh0jPxE+CcKYwsY4qAt2ylUCVt1I0+tKMHsQw+YZOdl
voux89+3GdxZQ5s/hNFaOjkjPdWJ1MKuUmxM2XOCDUiLLfK1crxkbHmDa9CRM904
/q+2FmCjyu346uK7KKXAmFHn6MTyRjmFwQCCiUrib5xzQZm39n27xKYqDFX2AA4c
ikk1LJf02u0AsecTsUAxzbXAfyvnYAHDk+xacOLtxyZNxdVvc0/Ei/uaJ6QMG+zQ
Kan2VYYjMZV3Qs7A85cR2rb/zK9aBojY3sYqx2Bk7Mi8X0kKSRSgT2uiV6459fP/
x6JWfeN8cZmc3trQ3j6Ag7JJ+yuMSU1j+EAHySIkJE1rZyIWhRpySWVr1hietX9x
y9zC3anQeIYFoSchUlQxZkAp9iToPy5iw/umUdtpqzareGZ/MEP4Z0mxMJ0LB/WF
BK5aLHckH5Yqqh8vuCJRwJzx1OgXH+awri2ZJ8iJIUnXIxZn0QsGcPGlu3jvWcH6
X3daGgW4hHpuHunyOs2ycQQyn7MIrCislXHZIn6jBZNW+drm8cKUpgqirvnoBWXT
k6Eu+1varlHkSugSOCc29Hvm9h/ZTILPVmNbohohEE577TjdfBaunkQXnuzasbNT
dc6guzm5xhz5dt5LuaoQmKDrpvQKNy/Xb/qUrNz6vGStAuXuu23fDJZO9CMTRSvC
FOTSsc2bmEimO2GIuNcMikfEV67T2qInlFDRqSR65jlCYP86jF9fVHRfPzQfNYpU
DqAxK0ltPCflInSXQQDgFb/qCnp7xt9mdX9YekLLYAdyhtk+sBI1gBlI21ZRyPEy
1KtZjpzNhC3CfClhPxYay8mPapBcUqmDW4TrQYmIneGhY6IWmNPMY7ZRTYQMbusM
FFBDp3kyUKJKoNogdUoh3IRvpfQr6r6ufBKiM7d9ev6blArUNmnAQgtwPrwglLrL
PoA6M36Q+moJABUvljN8VHNM4/cm4tJvV3Der+K5DsGFbLkRKQhS6LOU1CAX+fwC
EPeICMOrXXtXaPZf4je4tV0oFxfG36qwTktofjapeb5MAMhj7ZlIRcbMcvwNCORp
LjRBfoUM6p6iqYPgloiwVBpIDwlAItVun6jbbVn+4f14lrh7ulGBFUD4Zzb8Z7qp
2yByL0FR/IPhT5dpDbesTrRKyjmBUh3r1Yrsj7rI8bd5ycbz/3YFx1nKki/RVVek
BFM8TK4W5hDW8LOKXK3L6MEjBxzLLs9HuzXuOl+l/6X+60lOSYB0crf+H+G7Wyfq
AaUN5e0ktxnfHAxRCq4lULF4SY7xrxnr2egA3PyALCo5e835GcrkEBqxRsx8+1rU
mY/NCbgGoQYrrSziFZOPrQyYuchtboJHjS0o57PPSj81B2ZYeSmEX1qhKhB+eq1E
nQtnDAZVo6EP0o5GZ3suN0wvyF9Jj/sRNVcjPoibg2sC7bZcMgm5nCbsKCZ5CRaT
78VehZM4/LfYT+KMbUrSzvtZ8azR0PBL+avpadN0PRcbCOaAHDTMIl/e0t8y+FMe
7NPooSAZpU7+joUd7cW5rc7GkvsB2sIv+UXRPQLkR94SreRJb75DqngFwsO6whnK
nh0zIfSB7qgIKYvD+A9ZrJ6NXioE1Z7rIBa7+jW0fep2+tTr3NQ/OfAm/4HGn+GA
DFN4ln1sn+uyOrauqu1ZwEDaaefDDHt9M+xaBF2BX+5AkFQfMzHRFOHWnXVbyVDA
p+795FF2lRzg/h+XcMYFAN1dfI5jkk7Uvh8reVL81+dBTXm1v4uDV/qf1L0et4mr
R8AWgdHRJyPc5xHAFcHn0TaLPsF1OfiYGsdORyDPNw/QD7/34G9FImJ8dC7lhLxM
66EchCxIvMR8NRSuMQxZCGt3XgCSxalgTy0dRuZg0Pkz6KIaqcocoG2dxsylc3F/
DzGwtAa0bpfzyJvzRuNl3LJQoJNLeBz4H5s18v5tV0FWnAEtACQQz8iFSPaXXay8
uTvpYjcr6jawvyfx/0K96t2DBJE+JAJyqJtMYGJQ0vqKa1kr9ADoB0r0xZYJiUMJ
DprG0NOqolSYx3Po7+kQ59vYnSkimgz6qGMTqCBUvMduvDFaiqWJt+DaK6DiQ39u
CC56/+Gu9h1rRx1e64ykfX39A0mv6q7+1eovrALe3l5WTRSjSs7cytEN7opo5mSG
318yTVE1Bf4HNlzepAudKH1KEJrbCsCyl2k5pxSBbZdlhhAkbYSMlcV1tWU5m/Kk
W3QwvisUxQxnuC6CtIe6OKgl/N16+9dGtdgNyhKwDsVZAkl2Ue9V6uWxWJZ3d7xv
dZsA6yShmgQQeYDFvVB/mMEKF+zwjSRhI2JRTRfF/efF9RqNJo7+cfToD18xTZcf
wOuu72Sa+0edI5UXST9QyB8d1IdGrbblrl6XnCvCCYTDDbKeDM+/+Z0EmTkC5eVK
3siD9NENcYv0gRclJmdTXHf/ocWEJJ6nKUfndm4AW/c4eCIRiDfRTbQnPqgBY0bF
aET2BLkrQo1Nb2Nti6g14oVNrP/6dw/zAnjIrHbWpq3w6SvDMle+lbONepKFRhMX
McMwDAKAvgyy3XFhkM1QoH5/NxwvLnHPFI/RR0c6AyfvHqOqN+mq42aromXzBCpS
zRw7YH5S8orBTLVbMuXaXuLvXlyk4Xr8UYGtbkX8R0/cidLL+cntcUXvTyWAON6u
0o/+EWcTf+T4txssHoU0G1PkM13BvMRed0kkMIGJPi4I5iOfWWOmmeJgG4aDVTls
AkLAGSNf5GllyRgUHjQxoSr17HSf5YG4/OeVSn1Gq1iBm7tMOkTH/GuEW89pKeAG
fcbkaYM/WxsunM8xu9cckn4QBPjACf/DvVjVSv4FVTGCyMHfFGoD0EDXBMNd0fhG
Fc0RfIRVKPXaLefNYBbe7hjvfc8+ap0kk5/eB7qRfcZ9oSBBSbrNEwzaTLtreByw
E67umhgayQxqj//ESBLWHUZT1MyeRd9L5k+CHbRZ1wjbZzjIkK6zbQd6+wVj67e1
5dbzetCu3mJzRcqzRp8OC/TWFg4+pBbDUbtCPySpSYr098tf2Sr0FH3wF2WOTEvS
n/YslRbNnNNsWGQlCKO0SJZTMErW4c/dQQRiFQ8Ck+J7GoL8f26Rfq5zat7vDxIY
HuQ+glC+ehgocf/LzF/XiMrFLFGGByecb3cXP1Ogr/fgUVuEk2ZXYHYUmeCbtu3e
ZsBljMBmBkM3NjAr5jgTtmoAnRWro5PHrp4TAUCYCOiiEgA9aYbT9ArFfMhXxGD2
AHFqZ6FbGuNPhn/DQ+G+t6g9hCC+t5LEe8UivpVUU0t0fZvx0LacMt8kLtqpykCi
bM4QBkw0ghV/0+aBwNyx7n6CILfNVCKtddh4zlomMzww5Zx3D0UeJZUE0p/POPPT
8yvhCOUbOB0AIze8BXnRWkX7tf0e7SpB4cD6m0rx9AWmX4HFVfKG8wHJTnjCKPq2
2De91R7yPBxviaiN17tqHBigk3Zo/bA3QH3S/hDo32Fay2lW6LZqb95y4mAwISGg
vRktQwa/7wBP7vmDS6WfdAzH199IWiIXY12DYtQu6Yo97AaLTGPf60Kuo47igedi
hCox/C40sK5oyz5L9J9UpXf5i/tNusD5jguJHlxg3wnssI8/u0ClGtkc+jHB0zTB
LRIftLEHt30Bt/cJErbsZ80vKhTJcDF3Wc514uZ+mWRuXzxnPN/MA2Nx8EDkOSls
XItPR5LOe7IjsWsZFgYZ2b1cDVoqrp6tenW60w0HQ/Q9tGeiPXO6V0OOeA8MCCiO
Z6g9Yc7xMVTkIa7aRLfPp7bnZ/HXW5yi8h9uBZoTqLV4ReIVTepoFrD8ahQm9uDy
jKHMS3VUmbp9yV2AlMNkJD+QtJVHk8qkX0wn6eIa1SFICsOLWqCoDHCg5vgC1xf6
10HqzL8Aj0rMZBfb+kzyugeJiBi7RxN0HtSDiDQgDYsn92qjuU8J/ri9xS75oy8W
0tsvV8LIdpQ376p6m4CeQaPbN5oLnWvwKusXyA/faK3OgpRt83kASpKnfYFSzCfh
F0ThzlAfLNSi8HLw4HyVr6KX45k0KZG4z/FRHXf44EQNSm65pF4EhZN0nzeVEUZo
ASDC6/BSW9Xq35/+Mbpu+oY3eK+ReFinxJ//Hgz4Z0jT6Jmnp9eXZEsiD5hqHEs7
vg9WEilphxttqYBqqfFuRh64dEjPA2TVbBebCSymY4S2aOzzSEs5ZYtrUEjZ9Dd3
cZOLxPPvs6D+Mt3C13m7Ik5zz2Jwu8az4peOyIB4NURcsNAYqgSW8TJ4lux124Ob
wcFYn1laGZiL1Iw+JAAqFiphcxII1AHQfDeBlT/5pmyOIAyyjSYDtkCYE4m9irvP
px67INZPuRFbZvYN4r+lwR8RgMkGtYNSPn8q7xx8cAZZoJyvdvAZF4qQ/0rVtuOQ
VqbExRfWkpVMOxTCw7dZsz43w+EOToIW/3vKXFOFFgkaE/aF2OFgnNl8c/onfWKb
1Dnpg7NMRFePiWyhbOLS85BlqoRYrSLJ4BRFdUagW7Q4tL4PQSTV6hBEeB1EVnS2
xsDmkFKO0o5iEChf7cykzMbRCRQP2aG4Y7WU8bkG+qcjwbxTOexSJiBUmhlHdpnS
6745TrQiYDnvUAshFgzVGDMs1N2lspUP6bh7hoktZfLdZa5+YT6W8kTnyqQYuhAf
I3bDdiyX+MJfr6vLZDceRQsHJTCSyVhufU7q9jzGw6uqUek2RTJLF1iHKJHKrVHI
eLALLS4ot6jacMz4oxjqdSAIkFTdo/Cd/dgoHf0vH6VZYDW+HAvEddvprr+CbMb3
5tgulWmE75igyAhJF73ltpIhxiZDeC8JI/C++rVUCJAgaxHt3X3E/oALRFUUjHt+
tJ7sa02ViOcG9u4vMEtT+VrBVT1Eduib90NFXcS+1F7UcRgCqft5K7/MjoxMR+9d
reOlmM97uAQ/pkM+RUtnv83ZXlHAtm9NJuM7xh7iKWacfBOVU6XZO6muqw5bSlS4
oczlm0qYRcCqqqxRTzCGTZ19oXAOsiN2tTVGm25YnXYlJS/AsfYcPQZclJo5VRal
hiOrpGTZo9b+N6G8BIVzYDFbMjUaYXcvKEVDNAdhFJ5cEnKl8Lq+hDqozdzp8oye
+cGwzsu1rRws/k/IvAUdMHvoIj1ajk4UqXp+Y8pRx9FavxONwPtScNph4iRZLL7i
TuR2uvQp4zt8zKcJdTgBBGFklJ2eeD9JVCLsXeRMR1OPpHU5RBZWHxJ8kMXh1V8w
8jxq9K+ZhulJRg6sWJuhEGh3xx+6oN3Y1oYV5ugeBpyb46JJ+p1w7jgEwIVnHERa
hXXFMfkvxHHdunOomLTDNzqZxKrSuBmAWvhG8nSP/fASATlegrfbm3R4vzaOhRhN
P+m2kNrihrzrQEiahzwPWH1kt3s4Vuh7R8i2nf3bA6IcPJALVQQlW1wuxY/2hFLN
2gMEJS1tewCDjXmMNQWddPnODoAh8aSO/P2SxRVHWTKz1LDcA/Nca/xMyuiKL4ly
4Y+p5o6vbskNe9yVQv4g+mWJCV0Q3B1dHY1734oVSXrFycLUX4K4+ScBMimTe0GQ
Vyivjt2sqdDCAcx8G60jRsxdqXBHiifUZiSrfs0ppmL/Mqsf0BmpTGvpOmk3+iOn
hwrI0yXiGA4u5WmtIwAmFRYtgbmA8FikxeziignUvsMoN6eFlA4vT7bB41KFh8ta
I1p1ZcaIKewvY6vohi8TLmzCA4Mmf9c3MMb7rYSaHe2xYnfI/X8qUtXgdUacqUll
kpKvx97bkjBcZRM0UdaxIhrnKEkaie8VIrC32CdDlt7jwMJ0cppCRIS88CmkCiw2
SimxiLhYcwJMA7Q0Ce2IEnYmIe+To2B8XT7G8GJwGK4QxcHgeWgidrJoPdjfpJYS
8d+gVO2FVUKqLt1LhH7SRyoB57GN0j19o9AaY3d9LZqwOfnfICR3NlysDo5sog64
fEzg0gk12xuCyJIt4ZwDmRWCQMRcctui/fUQFNp8pJouad3c8sKrqd+PECCbf/La
rZ8oVWrg9LtTuX35OpsN1YKvIpETm+B8+l7UQM5mXq28MYxrNgYCdOmTOs4Swni1
0Cdgo+qlpvpq9HTDMbsF4RY2I2TLlY7k6riynnbXULVCnCzacg5O2MtX/GJc9Ywt
2EOEcpo2qhSIYWoe4Lg25SY3RVN3Aai6SMMWcw9Tn5fP0oSDdrotJO4hW/+n5o59
VNI231Dcl+vyzvVfPY6gHkhB1yb9zy9AZIt04XzNA5scO+Bbxnz05+kwwDDnHARt
4UBMwjwt9tPR+juciWQq0MjuYr72ndLSyvuBvZaxOvswFWuNia+nH8QGB3zs0yGE
OODFDdbUzIhllwG6o5DTdm8u6lw/HOeA0Dp6TGl0KH2xrzvU0k4w8GnWpquLL4E0
JKcU3p8t58LmrmzJWGThd2r1mzgY+6Fy+yg3F+Fr3tXhr5FJXaCMmUtn7hb4mQpb
r4dpFYgVo94hBcq8HjmTcB5eqyng9jOVO1+co6xy1eJu7WGPPtnJFrI6SUqHtI5U
VBXW8c1/aytBh5h9xZTVUii4ekWUR1ZtgdWDDCZRNhjmizYFB8iY9dySWs71zkcP
1fsxADjvvHC7G6gjCoc7XwpJ1ZSmMqt7eQ900mUhGpc3j1OJzOEwU8KXoCxIGEwu
ogeeg962vL+vfC8JAV8kbCk5hfwYM8rro5ICaiCAIeNtOyVFX43s8Ci/EJZfSnT/
in8uoMS2aoka3vyhfV46MCPfX+ZCtE9s29M75johJszLHik2baTgSjaD62FEMQro
s5z32ARiDhkf1UeWEahQE83ERE38DS27Km197o99GkwXQEQVlmYAjhPVmzOuITQf
AMAZGMBSpAcL0SKNIzvRaxOSGV0LPVKm7LmLtxDAtVUDG39EWO3/ZPL43Bom7jJd
gakXhXULh1KT9f41EbIyrj2gloy1gej44YKWwZ4j1Szx2hcNdrQO3XwaEUT6vfOd
EZ07wvB1GFBhUcx/Mk8HQMRe6L/JhByD0QU5tGRBZehk/xMtF7pigXPN+3SCDdQU
tLmNuGt6V0KmxUHqqHQsuvRtsTYAxSo7IzUeHUggipDg8+cMLa9reOiAMawJ8LMq
+2MrzOsMgfdn5qaw5jgJIUa1naD2l8jXI8MgF48FoXkMsxpR8LFP1Hq9LXAOGE7H
MYXtcFp+iY4yMDTT7lLMdZCSrsRK41wk9R5AxXoZ8SohZhU8OmNYKenGFQ8F7vOK
OKwuIMGBL6itIRU3tmlvdZhEljukS/OBITBlVLQ7MDwT2mZgdSMEGZsohkGaU4cP
IlBaPTNNNFpW+6D21mPBLabsrmIP0/k3jU/NfqUVob4ivSFZENZiWO4DPV/og6gY
+EeONdcUAbBwbUex7Lu0bmM2T3fFFEPYpEmdz5Q2OemQg2qoTnxscxWPjELXb+zK
WIde4kf2IoLDjDXh7U+Ivrf2FB1Yv+MxVoqqkfM/qfyqpa0Tj19S8wMOJWrhWpms
ZFZ5hjY3mDqBMdyLPxzZwTea2Bbvh3Fd++a1nDfm+EjyzkeA7s4EC+fFUsaq6E5y
ci5RaTHs0GEw1D9gYez1PzyVvdAII8HURIObIAVYDgjRvJNF9NUlOLrmMqSTfSxl
3druus7PbchrP3XjzeL5XYe+xG4u4E5EN4eo1l/ujgJK4KM7qEJIPKz0l9mNcBRT
y8qHbGQeoHpCQ8n1uSbIU5Rj+KjFGMFQcYFGHhIqsw14dXcEbK6/aQaW0krFOAxv
BPO1LzFV6/8yBLfxy6hEtiCVMde8qDtm40ExqtM2pGmYJ+PC9vYhFreCjfs12qn1
pU4SEznv3XpGbjdDYI0JRJBplFqN+LRrFzu8PRXYnYyLvHnYCgdp+K8sGQCBm1Ns
KYMy5gOejN8j9vVg8uQcJH2kEk/s60YJQY/7DpJeF188Taac9bw9jhtEBoFXxSOw
ED1urjKlpb5u67c5apWXZH125QQOoD4t04iuzFnGbXKaPPRpIOIda4O1DnjlI8Y0
XTN+lwW823Nglu9hjgbCi4tVbrwgq0fBLK4rOtQPYhGtk00hkhHRuptmynB0ryfG
huBmN1cKH6WqsJIKFuiPR/tHcXdqDW8Ng6vmsNZ8Gol7C7yjr0SooPqKqSM5JMed
u3+hlNMxXVq4Pa7sI4Nt/fDCOPoZEdWMFaHoGrvTjSIBClfGYhDnm3awpSu6Ekmr
XG2/qUuUcTtqicGtSAB5UJVrGOYeXOJjjX4WS5O9QLGlR5rq0cG0n8VKgacdeGRh
xn5GELppohu+rgnqhaobi0qp4oFlYUSK0YE4dHgTZZjRFiGiWfpWKXkwtl4BhHpF
LecQO5RQUhR0O9O1s23qqd6fNU/4mSEbDgqWxDXn93eQPABe4PTQXV9sEfHy4iwt
v8fgalVitYrD3m79uxrCiItcya1c1OXX2+xh8j5VbLYTH57rU7PIuLyMXsBdhJLJ
wpqVausK9EIKM++rRWr3MfcQURvVhXIhqR863cjU0vgve/kl+pPJxG4lEfSZYxO+
ZTyLTU+4+NTGQGOcJzk4z1alcv8/AMjGeBvIeD51gMtndEa97LRmDGN8UWtyxK11
AbsHWdfomzkv4hcODJ6sHdwEBX7V6nh+qElXr9LSSbxZyPWi/SRajDyu2oi74o/l
AfSsGB/b1uw5z0sdGxhSrrIMmTsRO5jpSxxdcW/Rp8iI7pHl8rA3LFVKcgkAbLsI
kVEdfOyx3XBn+Cl+29HhX+kgPbaqW6CXkmwDdZVShRa22KJkkWk2y/pvyzZsbxMo
3T3HAn1lVXH5U98ueBrkis2bLrPfIvjcvwCm7cKY9pgeIAcmvO+dpa9ramXlW1VA
vYYSteHcsduorOHfkSJN7QVX+1wdX/KliqgY0ZOziIlQ9qPloYXLCPaLfpxUE8Np
2qd7XxJKFJ6tb+lYqpDoVGdmhqzAcQr5/EtfU3RyqgBJvfrNz4LzhZlXFLDiFyQl
Rx3Dhl3TpvdsdwX0IVOfAU4Dew1v9R4S1FhlvBdv9x48GUtmHyTGzdHN/qd4NsNg
kwizZ5nPkalzw3nE6TlcLBl3ZMF07SL9K8GB3iOT2uWytM21EA0w4Syy6IJNwVFG
dmMaQMzDGvtWak5P/vI7l/W0gEAwrz3FhSnJOmQjIUeYJXPCKhiCIS94uEpGZJKH
BExxvOltKBAEX37FZBhwcVQal9PZ69auR78oA68AHtIOZKa1wSYoA6r7xJMpxUBV
u/A2J2bOtqXzwJ/s1M1niW51skaSFwVfIFOo02NmVPhpwpWVPV31q8ymVSgmZWeF
5RiXLvut+UTeD7sb72hhp8G7vYQfDG+ipf/W4V7uX2zfcemYsccdHPtCJijxJXnA
0FsvR54BWyfx+jt1sFLOuc+R8CeYpADpzDKXtESD8dZd3gMAfx+oSO4U/g4yw2ZJ
m/4ImkL7auvkziEho1pFQ4DBweULdHFtqGqk6HwI2hNKEdJqMi4TGjei8YPWWqPG
6EOMM19h66Thf0DMQvnI5d4KobrWgS5OYPN5s2KqK2H8RgMPKTOwd0Z6E5HZcHpX
hsytz3Z8wU7WQzZwwC3JgbwdUdwOx2xs2NEEFjr/jbhdOFvT7dL46nF+TnVgAqtZ
hnYLe+Ew7MGUXwGpW+SDW7PHKU4BGzvbgnBNEFLkmyuNgod/JFefvluMTEH6mhZG
tGi+Qmk7kz/13J4cpgIy8itDD0a9rOuox2K7yc5QiorFyXPhlkuj6NLJGxPlBLo0
j2UY4vMOZN2FqV4pzqrNMQmvPOZYaokEFvRNLJjDSCKTlk4nVSvJvMN2rl42JTdl
TYWpBQ/xa1dinj48NYCVnez7lbky9ZnFfIb9XUg7tT+xSk5LTTt7e4LqcXaFZZqk
e+s+8dyQRFNJSCb7rg0XLkHSJAnfAUMCS1Grj8QTvFAZ/F2VkAF72NtsVVtzlA9m
X0LMPbAWJSC6xSLjbprBWlJEZtwyoTYA3ss4pnmGgEi32l6doTo9PmR7nAoX4PSq
vdWv+TmDcNPzS3znOZU6RAJfHCD3/H4jEDq4qArZGTuVnphQE01NOwflZHyARbQE
Ri6UQJ8GFBLyw7XtKUiZ74ccdijBh+v1rCutIrnaMKbrtuVE0bo7RjL2yMraBEG8
XD5AoJzh8YWUeU7dJXcJ4CTeBjq1AxL0tDzbQpY9GUm4zpZMomVkesRrPG4tofd4
qurk0MqxXYJfA2mQd/0J0/2nda8cBAJaiFJreJaEYUx+k7pDuQcQ/b2SENP73Pja
nmH3Jw1GCr8PGb3sGkwS0Lk109txOktC4wgXFmVPFnRm59ODEZ7JjCM9FZPwGQ22
QH0O11Tv0uXOW9zW/nrH0caGzIVrt7DzjV3dlRlc/pdDg5YGNrsCPdmZH8KM3Udl
euysmwjkNmtrvXlWUaWJAuu0XMbgMf/wYnb4Dt6LyvI3IIWZTwPXJ4z+lq+Ae8Gp
9azBsBi8K9n0+AqBEOXxQ6AJASXIckjA8PNu8EAmS9BCX6w5/bsU3c2NaRfrAVd6
cNajX4Y+zyYEl6B0ROspI/Jpt0WKwKDIJTNrztmdN+b0leaBNBfarlayRqJqAnPN
J57TV0OAo3stI1mk3bqgUSYXe1+RbbQZEEnqyU93W8DtA2BIjFJ2gx2hGl2JMTHi
RgwPV9r5+jADYYRtvTmio/t9onQZDqGtjvmoScdglJdOBvhHlujj64pvs4qhIPFD
DS54DwRdQtA1oK1+qtGXMvyOUfcFwls9n5Lub5bvCX32+O4PqIW7QA2bdF8qtxsB
fHwJ2iK1VgqVoz9iNHv+UD3/wB3EaR86Lliv2Um8oRovVWy4N46ECTfsU7p7BB5t
lNCFSSBMF+E9Qph6tg8BVEXoEp3ZvKDejikq1I3lrNerAUHbu3EHlv+XgOuoH6eN
aSrqn2Gwfl6sOL9WWQoqV2y1tjAc1dDoejo5DnnRbIdC82Pm5EKJQBeTRFjZE33E
CC0+zVX3FO4LPjz5MDqTSQK9PDJQx658Gh/vYtNLNrbam9hGr92zevGGskADGyj4
KTpJKJ4RfzulfYmjcWtJ7jZN0mn7+iShTaDezWHyaqAd7MZDG4tUFB3lVYjdOwG6
Q+NMD/XbL25l+Izn0PwGYU3eyfVOTK16+ZYZcuO098UAPwzWkDEx/Y/41PtHjF6z
RAvGCPcuZG8dfuKZi6CE4cVM5TakVMEZ92qyvcC7A7cMKXjBNld4qj2G+a3aFIn8
pJqKfQSOvirMfktgFKbnjVlDN3AfeabUZcBkCX56zWZCJuKIX5ey9OEpsLAIztfR
A7ZLvw+LX8WFFhocO7tvarp0vpsbhnw0TQ3KumflEQGLKalN9SIVBMgDe6yIxtOD
kv/aI5wxdFShNGEe5DMZ6vEiTzA5rRoq9D9C/ouBBezoazPxiXjkxBGgk515rrmA
aFHAFcfVMcATOxrMPVmN2sxt+qDKnJmm8itf29lkz1GomUT9Ft4Cq8DHJ3MdttZM
O0Xo7zegGX8Z0rHzmRylLWFrdZA9hG4u11/RHam9fjh8aT/Oo+O5ireMUWocz1fb
yBzaL0aksa9WBaB90uTh14PY0Zt3RNJJZ9Rjpz37y5N7q2HSMisxWj0NksqEbr/Q
flu5YmWtEfnkS0uyC0s/YxJ+iebAhaHfvhydKtlTMHfXpPzZ3yLK5XgFjBEPh1D2
1wAYuozFFc2OxpjMpgDhk5t6sNgkxsEPsEruIgAXxrRYHLwddM1uBlF/RpO4vcdo
SO1KFHS0KU66kZY+gCeCgoYDqzfOitgkahSst1Ld+JJR3wX+EJCyobMpOMaLiDrA
jDE/Mik3rExwHoQO02XremYYVqf7ULMFY9wTBYtk5Gujy4DpOukKvWUB5KGgJrwV
vksE/5YMKNoEkxmN3fRb23m4URCrnOfzSEsWiegKgFS1cDM6wedRiCzA1iZgKS2/
xgUs7uuQkRB8sFHyun5JdLs99U1U7dY6syCJNppnbs2Zcw7sWVtiJhZqABtCVZsE
gfxmPT+RcX+KSoZd+uMMgH1YCP33wo9NXeWHRY1RdnnEbaLGGwpLBpeZ6rZ99I3M
DbSWMMiOBZAevvSG0et0X8kCxo9RUkKeamBX+w8WwMhaP3t38M3f9ucuj4q0/gAX
c5YzWRUeMOACSb7Ym68lqT2LvuSCr21ZgG6wF1BPG6n8lWhtqWbP3Iy6cVtOMtiP
vyLeE4x7bpQ4mI1NoB0x6nL6sqQkBzdCsFYQneKOkWcPN2M7Jjz67swGzQlbEKE9
KLIB0uxDqsasjdKaAyqo3Bp8urHyRt2Dg5vf+Rhj/7XWrUOnHgeJ/Lov9lpCF0VE
UUN1mkTTDcaD3Mft8+oIOrQigJ5mmFojKWmottaXx/nhIKCufkVlY0JtQAx3RqQA
FscnbSPM/DzK9DqePBAHt8ve+Lkzg1RDRRY7b3L9D01Tzj+AWNEKPQx3Zb1gePbK
hwra1/aGL4L7xeFpFy9AE17YdJFLS6DbHuGdOEDDgALmgQ6F8TrzOKYNy5l7W6FW
JwA29qkDAI5M2j6QZEDlKU3gGWMZJYtQIMqGPgFgG7Hs06YzVDDbyzkL93vCZtMr
jDNzNGoAliWp9KZ4sib1niBVT2SoHOvafYw+IGIjgAv9v/7ZvcjrItuqp3xSXH1S
CprfjbLN5naHHNbJNTKn6YHuKYsyC5P+dNDw6jbcHctfi2aPVU0JKFe3VwCqTru/
PLk92L4xRi9r2g0t/SIqF1FK4ro1CPo5sW38CHykXQoTHNam9p7+54TpfXehrtZC
clyVZRjxi93FZUgZVZIY49SjV/eMxdTsqPbas+8L+8qTn8LXhU9KC5Bss8keY0+K
bESdo17tTtJ5G2CQ1I/8jIdDjSVKxFAvwOoeNpXSPv/uGDl/ziczFWqh+u7aOEwR
wkyQeScvDn8xdFFH57lIqTyb/fhSmZR+LxcTQqGjci7vdb+GWUhIyTrKdWaetnO/
/PvQuL/XoqQPZ33VvcYvVY+7aPFfFI2voNm4nZblYgJ+J/93vKFfehMBdFMXpxgb
88w1MfiiefTR90FiUVCQW/CTpEvJw4lb5y7Tzvyywzqz9qMYQ5whcdPqOV7MgRaB
rNcedHiQVhfT2f/uKWk9+1s4lMwtaQruT2pgvw1F+OCKDXIo/XQiZpDQ8LYi+Lac
/2sDuJBr+qFKJ4jtZu5U/vqcHN0YDhTRXslGt+p38MtfBPmnHe1BMLZBPBgPiytB
I5NJ/le3ZCh12HYU9DPU9fVpqCK2I6S9sKK1y7+x4GiUwKYlPE8A7/FgyFxDGVCT
DRxoQqU8U2vSwQ9IK786372lRawxFzJJxpCFRkoth6uGyV7lymNut/bijhzq5T4W
8Cg4Mt+fDkJbRxawI0U0Jt0SjiVaj7odCuFAvo3c0XON8qscCejnFluZP6zj42te
I7J3R/h1iYWPC4i/65KfV0cU9zl+Ys5O6sejgE5W7EMyJfDYHjButD+NUoEL6mL/
vc8QFkqmf4onibNAJ4jAPnot3+aTm7kPeNyGguG8FCfSskkiP1uxhPmficeZMZnq
b0uA/TE8BjRZJNCt6TtGGYH7HjUIrZPl+T7eU87yOUVKkMP2gg7tLVmyYO9mdT+Z
y5l1Ncdz0L0V0J02bgNFlLzqsh7ot+a12pkxO+dSqGjnDUCHNoFXcVkcYBVtsHrS
CbWddX5kLb/w/+wXR/va7B4o+o6Uc9d/pdwS32+qCqPKWQvRHelcpzAgsSxyTLzb
3Vlc7BJlWe076Asw/4rfrnz6X4Isk8ZD4Am9FPkqOy9z+84AGaYOjSycHcZ/J8I8
wUqyCcUurZAAEWvf0AA7pkF8jiALvaT4eYK635FmSUU7vr35dfkQId+MDOXYv8dx
NTsN72WofP4c1ICYGpXdjcXFBhiVnIhTRfMckJIGAz4sjceEv1ofYbFTB6oUcmnA
5GzC59wyq0w8GyLC0HuTqb1lWBgSDigFZOarbcCNJT4s6kMJrCxL3VXev0MoKzrd
RxHlbp+/78RC5eUI8b47OCg912jF4LiNEd5UXrbuLcgITRIpxdrJdymWce5s5FYc
MF6fSU9nChpcOmFe9q8XK83GmSZutt1zWF6tG3T2Vy9xpJtKK5Vn7JLGpja5aP3L
ktjE2etlRjKwYWgvVBYD19JKCdYphUmdOk2SLxIRtFnT9JhYSfmneFMwjgG/31Zz
xueq3ybI/hRkw0WIxmwoa1LBfuieit5pYLKgYQ+uJMMLrgqL/1q73EaQp4yXOt6X
J9UOijm3gUC648lzzuGMp9JojOxuEgODKhNHZ9nOaBvr4Qhij2YUPoN0zXUz8b9O
sXwAo05OebU+qxnozxo5b5UN2FvYJmyDLeereydYl28aOJRsEnylYqlTQJORzFSA
YGKXFvdixviyQ7XHeNXfm43DJd+6osWU0SQ0qLDCmY5fQ7BxK5vo2ZzW4OTEcrPO
LQgV2Jru0C41eOjwAKksClPSxwLBQ0AwfuPr/OPZw9k8IUVB0PjIQuLWRWDlU7Cj
l+mO7rSbSd0ZzIi1uiNRAEfFfKMpgyQBtgkFpsLauQsZY7GUZFW/L9IPgha2vSZR
jXQulGAU5yP/q3Zuea8/fRf2VsGR9NSEjcu3gIEbELKavBGJMGEg920D5+vF6a6x
1Uc22jqxE4IyMmMBMbKki33HdXBK3Klx434GFoK8OHQZTlhotP2HEZgB4FAZBDP0
okntBr6D6XdN3P3gR9U9qTg0rS+2NeH5fZQLpCY/BwQncTcXJIg6U8xpVTLLIeyJ
SoXASTpb+UB0lQDbo+lGEJEvQnkB3SUSkdEmr6HYAJK8ktzccO7tahojkPMINnCj
96rPBMfUAYC4GJxh5mALAIBFuFYNyP7DarKr0ebleuq/Vb3wu5OjwQjahOGAqzf8
QShF1+dWmOwpZkVDMKBBNYchm5pngjxs/lPs7vym/I8akPTQ7dPnO6kn65tNJ72n
ZUwu4aP4KRhToSEy5tfVP69w/r7mfHmoXrVOdAUv/m9NuaT95k+49INc2cO2Jxel
XiHO+OlXqFvgttFUsCmdrNR0TfAB0+DCBdAZqIXPESLsj+qgTTJKDw3+k+llk+l+
NXzVJ4tZ8O7shlFDYxDN+/MdTe/c6Vel4w+XG3RSL9zfpeyjLsaoEE6ItFqPzpD3
GzMHGTpQ9OJ4+JXhN5ZOWaDn+KO5hqpKccswdv8c/KQImCAjiwKjid28NqHKXYy8
vQhrcJUvtW0tfZHucEoEPOfF0oMsD9BII6gEMhkr33MDjvpXyQlJme/uHzN+k9kG
s6S8PkIz0u0a7u2EppG92pQyeFo/tscFMHaPoUcTVJ8ok1y4JZWbib0uDEsVebqn
mggTDaGGDnmR1kkE4SUFGi9aOlRRLx0hQIrUQZ/0QgDlVCVVLhXciblKp3jcUGVi
cyaZiK2WKWxelyDiJUFxwaM7URLR/8kYLhDwG/D9rOtqEXW8k/wsyVQL/tMqsgiN
ZD58gG6s3FFuBgIkBOeqc75aDsV6kBSg/e/18yOjE5q0pwdJAYsaJOO70II2D9I4
4CDOq3YGXdJpcfteBvmUrh2OH/dSutxsqJ970uDrwbH+U4KiP80Y5iWjepY7iIaj
cA8hFqTywoW8KnyEB2RRigY7sGNEFjCCq9zgytyd3ILQotXUCdIR7d4CWglPVEn2
63b+mbGFVyN1vBkiSWyIDXUhS7WTl296m3rE7FbJMIInYjz+y4M8rsStu4F4gQIT
J1HyaRDH4ypaxvxkJm0dlOVDRh+PkIU7Y6cOU+3JdUaoPYQaY0nr+iIxy0QfaMwn
PtFWAKbtJmcNOkJRSKcoXgkmMASDfX5Tow4KXcf3eqras9uPvl0oev4Xpi2oFGF7
jeghwJl2XIwkbxhCJ7CjlaBg0ZvwfmCQI5ZIf2PM4CTWvxOOuF/Tr1z6PpjqH9k3
2aB5cWbncImJc2FjfYy1e4rIDjFtyWmXwUmoFIemRur5OB8iFkqfYlwv3NSEgGvG
OpNXNyf2+AFRTaql1mFJyaO+68RKHr5dE/7mBSQz5n/VKvRNw8M60TS1zgmKzVf+
dLSnV1DwYwzh3fMh6pgp3stL8H+NZ9322NsReQfmUm4yNpHbDstk4cBhoJozyu6/
SB9s5yqog7z3W7rYsalCcUW3V2RsL9mZAQ3m6IzxWoLzVMTzihAwZQ4n4SA5U8uZ
2x0JdYeiVJ9QEPZhE/8z2gHiEvndU5phUhVXMEyXl868jGvQ6B1UZHQWdv+EmZD1
fyy8u8cQrGoWObDWFNic+Bxld0C0zf2+BaH8wmgxIHTC0qbR5x0jIT+EEgzZuU+K
m2OgPFWgVjUbju+obesTg9TV1yyqyYdG8qF18ecll0jFBJpjKWhn62CugEhx/wx6
ZwPA9++87Db+KR8dKmKd6dULm7WiaMccgT8+GrEgCmr2ojRYSXIlwaqOsmfgq5oF
OjSPvPUtIhglSS8XpJo5/4/ypJTrccx+KopjPE11mYbW93kZsztb2S+/WbQWWvOW
rl4sP25PMeczNUUWXCCDQqNKYE6IP+mXTJSXlRrpKKWSiPsqpS61FujOGS0jfDBF
gxSEs20sovWL6b14eP9Ep3lZnnkjLT4wpmyMsx1JgnTVrMF6fWPCUNpeCDCCxmjH
K6SeX+hKn/Pnt9P/3XLlGFrRrDXyXQqlhJEIljlh+GBfpDfIziBaZzIgQLF3OiBy
q0o51R1eL4RMoIUC9U/l71Fdmes4IHhqxi0no/JlTGIl/8A9Nw+aTxmDR1m6Lf1g
FcmKeudr/0Rp+OtMBZfcGmLYcqoLrqNwGBgSbKRJPiTzEgoqRPOaiBGMg6wCQBdT
atn3M+4RAxxJTCVBpETt3itXzLz4q3Em5Olmgm1tKX4tgS1EragaF+A3M1hrfTn+
HKDiumqfGu0VLzzE8aiyKCmyg1U2mAXpKNmNklttKiiNFoQGrSxEMInvfHMNeKo3
lxW3ox7kjPcZGlq8RshRQQ8ELvIZ2P4TTPjyFHthfnDF2xYde+NV7rjt8YoSpwdN
iPW0h/OJoUobOLGXpJHIETy7EHtOQQz8aYeF5MTf6iNd3t5SIA5KdHg3wRNSMvNN
viOusScuOOZQ3QgTlqCvtwGULXP5Xasqawq85dRXrEKeANzALJgGb4PM7ZGfkfp2
ZmSBT/o6lP0yDISoGNUzxITpTdukzgk2pcDqqsPSO2BpgaW3qbJUG2oZQNWEpWaQ
N04GGMhXk0y+4MtW/OsIPGcaU49yoEMF0999wxyHw6AKmBvPQHeTegZ1IS0t7MzI
/4TWu806BnBtBU2inh0raDgLNWlynGAFhCHwUkx0H+nk7RvLULYQ4opvywpXNibr
vvY99nWWpXr97ZhkAN3F+3o8izkPU4uDT46YA8t+kY8teYML4dlfGORWnuDpM4q/
8kNPTsMWrjc9mAUZQFHxj5zu4LDVxhGfPbgG+q7ugH5oAPxY9WwJBYCTW7n+QgiG
pn5Y2ALALDugmv2GzlBT7vmjR2r+R6sg9VYIvRWKqhNnLEHWcOQLU92qW58mM8MT
t8AkvzuhApaQERQPagwYvBY1uRco1NmlptUPmIhnSeuLRx3VE+ybB/POkEMZ2cv5
hGi2lKO6AjfTMDiiAwQH7UImQlXUduMPocz+AKvXJrKAWqS6I7WZrC+CYMdWNndg
xHQn/3OY1goP7mr4u1WYIGSTGu8WSeQb8dh3I6La/KfGLrn7dHx2n27GGtmPBO/i
p8vvxps0hdDe2q9KZsck7cpp+/KSqrg08Ha+DP4iV9L+HNrCg6YmW1w0El2cXw4Y
thi0eoKzqaF41I4QPj4zU1T1KgsyoSlv6ZtzG4LXjVLZk97xBziiQN/7zlPgO8cW
/mqsVTXW5p4fZNXhBrrsE7fsVeNfnhq2l4pTMjpbsoqLkhopv1qSAPkoYKQC4fKG
JC5deSIc1juYtCwmBkNWBM4lPtD8Z0Bggb/70FgVQ71qTyJWgHCiG8r30aMoutyU
yHiuTxVn3rTeMz6fqQ8mkdmo6pvvtZ0YrJLhpxlpizHnbV7IfgofcLcwWff/xH4G
epoVz/NosOR9ym+MFNhVt7kqw1Fn3ifz1jGyxgRZHFG5w0XLXJCZFiCB/vuZjXcw
wf4VxGuj7NWwv/J0oUJPLlasFGn6UbYfxaDyjFu+lGIHzMvo3o17g+dvGvV8FUPf
hHds0W50witlP2I6AWselu4Hwpb12iZiQ5o+kEonY7xTBqzHmbB+DzSoK20gT1Vb
bmifnivjw2DIMHP9KNN0DQauYA3HzD6eZRs7iyRg9+cREzQME7d4AVUvsE8DlD0g
tg0tCpW5RAVjRu309olez2tLbJpFJEDKCJmbU8G0QVWO6maNHP5bDt8c7j5PDnGt
kXCgkMahV0CDwTj3Xiw9Fvu8mNVTmgFhlFL4yrevoHyJVr+Vip1vVQ185dvoXk2d
AgeaaPvIyCJBa0m5nSCMw8A/Gl0RqFMktmJXeshZOmduCbNWQFszXFX4teM2J+//
vPshehma9GIU8mcQP59ev+HNCORVcxcxq0mToPk2g0sdHkUrE/xkzvwrb8SlH1/7
9tQPG+6gYjlx33agRDzQF/tw48bMI8xef/sYgukv2vW9xpBXklAawZz0aTRxAmSN
3aR8RARBp0eqwJHpgHs9KSK0B64fniVN+qKNLkxzSnGa+fgLSW3mf0iQCIQueMWM
Tf1sfHlevlIowRkXTIAr/EslEVTaJPTMw137WsJxVLP6YF2WbAAnCH1t33W7c3lp
61yL6UaeNqpFSTKQOY1+LhsTPjzwHv9JPjQ2VEjuHaDDTfpJoCE75BMROl8pIPZQ
KtqNqsUAK9EqnsukkR3Brbe7AVaVgG+1MALpaQZTlEjUgLKttFfXIsvcwoTMClYn
PRNrUEiABfgV8i+6bKKFPEN3/egPOcgFd3PnvUSYllZZ+2P88JvUcqk8/EmKS5mS
whefBLrpZ380BkSvH2b+93YowJS75N6Oz6gz9EOPTXSyrIZJ7HYzIuHACfEk7aBD
k2s2l4BQTUfhe3Ird5oyZ4ql4RBzz8cqUpK7ChcNB1/ReyCJi8pAGZDEIKSg5nKl
u2/McWbwTcKg4ljaOCP4WIhnVZhflAchxUObc+wDRs0G+u+hlpEMNetebrvUK4IK
kK1t1b07rBpauTX0mdHbD03JxSqE7blFRHOP8Te3DHqzzm0oRAFRQIbzoA8B//3G
HOACIof5T3JKbPAQX4u9LlrmnmkB/eCULhKT0/ONuu6FOuyjRx0qMKQA0V5hRJKJ
qXxyTBGjIULx9mxPXWK16/CKMbzTrw/cZ8DsdeHP+js9kmDrPHHtdiI6CKVUiFN2
KqUc6ykyqczyeUfuimycKfFkNcSE2S4q/2AXvpEBC92bQ/rHYEy0ZRB7kL6J1Ipq
mSIQb8jgX2hdKcgUUzDcSQfZU9OKwndQjhSrDFg2eYKC441JpYu+1Qm+mV6pr+8e
e2EAT5KqI63dAm5rj8Ri0AErSlwWISaJdjpmzvn6/xFabAKk5rcoFkfLo9Gq0jgw
gg+pyMuEia4QwjHjvmrEjTSw0GkV/l2GgWtSl31nzei6DzK7s7n7gdLVb3qTphz4
FBpvZCNCYG6RJOF0eDhxqbRGTBHj7YR2dMU5ub6qIa2pfI2MMI52tgWilLtvCMqd
ZyV6nd44Glj7x3rJriUbXQF0LXtym9Lqf2RQBupkK2zvzM1HjSJlKDzK9FL5+KJA
YTdaoOUAwofMBAkPGjoRZjLASS/YlfDE2Q1/8URC6vDdtCWeKryACyaevaPSUV2J
s4g4GwxFuCrCEePid5+RUM9szmng0WcRNIsZ3U4H4PMND/Fr1gFWB7ey28OCiacT
VJK3SwqU032ZLdC7vbDZEWW9dSPap699IzOB55aJikVnQg0D1xxs1RSBMAhAqva+
iWg8q5hzP/dMlfL4Q1VY5FMBeRzOLEuwXS4297inKA4tg0MT+6eXdIC5RZLJa50b
wOzP/XizsLqoajSjQ3hG0stmKHLTTcySZV+PW+KtW14zE0uP9k1jUCyxYVjC8auf
8G4QvaN2kD5ItCblQHH8C7FXCp3Vp+PwTEN71/rzfWtqAj2UYhrbMGQRB7mhItmC
QbfMCxAjsia5d3VhqViqjV6F+bUkq9wcyAjJgOLjw94cAyWT3U4+azNqh+PSuTjR
KBzA/vFUbeD+rN7J0tYLXOmlHkGRBvYCSPMwM6wd2SpALH1VP2B3vO6aUtdbCCLE
1cPJWrRRETrqUYSefG5XKBvbwkgHxpTOeRv9ydnospK2yn0RsmR0RD1KctPvkL2r
6g4m57QqsKEMAZOqMXD49RmXnETERtTpAUcbH4/4hiKGa4enV4Hb7zfa2wgNcP4t
xLbnJn58e32VxoOkYCT0sGThtx1gwYRcoToUtxWvv4/8W9orPsIm/D36/hiwfhTe
tPWxImzux/nCPAIf0pv1cB7QowgOL+bXc6ehrHkEyBwXbdPPz996CQRwI7QfSJwo
uVGaULghske7HMUOOqLRbOXeHwuYpSbgt7AEpXEKTBTUSXL7H2Ke9FoeGgCHprQZ
HTjbWaESZ6PiUxUkL0BuidrErUHw9eAodbjjyEm/e/mhXoKyCzUTQtJkSgNbkIXa
t/DlifgQQN3Ws0X+pGDmnvv2XAKXBKm/QW92BxQcyVjqsUpi43mhI9fe1KPcAJuy
+PExvdOlAOWS+FeJsehBc/pUvARMzOL1KnT8NzDMsNuaCmOASrqVhFZUxbf5dJvM
I74Y0jb7QCwItFEBNZKOkrg/JBXXQx2x1xchEIbj9+JMmUFu344GF04WczdWFWt6
hYbxsQ9XNrOmcbtMX9EbpuNePM3FtDO41YlG0hy7e1UUDnMWblmG/p8orifJ+DfH
TDXBLNXflc0xQlBilN1jvjadIQUJIptiF1vYZVDBLMLkMlaOOFYlzwU51gAL0126
+RiRgkofmrpPgbemE1K4KOw/gtPv+sVkJTUEZCpMBinAs8W7Q3PEmijWvtlkTkUb
Qu+HoXf4hRtphjpFQUdf101m5pm8Ny5J9IEfEXIUghanl7fxuKg6Jmm/aIexAu3F
J9p/bJx5UHWro7r+V9wMMr8PjVMVkHxbTLDw+Imh7c5wdoP5Fg+Xz7E6vlPYcTAV
mCcH9+B+b4bsouFt+0ECTV0tejUV96NOJ+YCHm/3VQxj+SEljt4gGdDIpXHepAC7
O+W4KF+V/vAFIRjQyFET4DNXqrH3lz4PzSTFLxrAz/oNIn/x9m4bCtM7Ta3l4e3I
2s8+/Rjd8rVpniX74HT4HZDw4KmF+7ZWCFFIYOGK3Q4Q7/pEiD1Ui3gaDN+My98l
PaFxDM0RK3hI3gzaYaQkgEh6iw1C41S5MkPPqNB0qoLF06LgDQOYELhHK+ovOFOU
X86C0Oh2ASKTXMhvRUO4VIy92ulo9cMr0DHpWXJLHKTeIcqccGvgCQAUCVq63xwC
qVJEZev2Z0MomPUM0n0p3HiwNrXKu1wDzB3H4tx2rV4qppges+I3O/D+uKLrgIC8
ttXHRdgb6hcjHQ+h0IFSrsKmrn2M6PyRUlEUNPaJjmVLKROKwFMJWDrHGV9nRjEJ
fho2fdLabpGX7bokLAnph/MZUPMFMIQtbZHFuOaBBuzxe86Z6L01sefbozN8JWTP
tEKbRxG2WJW5DqqaUOI3oClwCrnyAmp3jJGn63sPIP7wTUNkCB+GQmINVx9RSD90
r0XpNy80aMwIGtFfDbSIyDfese+woOikkL4zA0UJ/+oZncjC1tjRfslZQ1IWvqH1
eijmfIictzGvNjbksXvrqa0sPrm5N0qKEZJy3FLSN/41AmhQ1wiU230pauA3wTfT
6ssrrvZlskg0UflYLTnqdihgdwnZCRQKvCi3VME2ttJnfQ3U/8wiLhHv9CW5EjIw
F/I3p2nm0Mga+frr/F2e/5GQXA1SUYu1lirpsHPa5anKr075YqC2LBfbJRzO/RLF
UldT7zOhRfDv/lfV6TqTTkkATMPDlkPChdSBhkb7gORbBjcTbc7SqHX5V9fDPIs6
B2teB54lWZf/Y20tggDV8mN6Rd1HjZkvAvCLQdZBJCDSw61EFjx+CtivnBY7ffoe
sPRGuTHmyMf5cdTbEOzAqgkiNeukpK6Yd8o2zVdQxKfa8TAnoYBEpU4O0caMm9Jb
6aPHYRwB6Z+yHc2pw4fum1JXM+ua9+6OhSchP3II/lPa1A8DSivgeURtjTBwC+SG
LUPeAZ82TqHiUsfCDWHdDE79RvW8shSrctiaxn5HDUL/RUDLJXTJGuWYmMN4np9V
5I40BXj4BfVo0BkgumSFd6S1sAaeVetTXbJXDjhxRDT9bSsYiZMylcTFvthzboxf
OxzfR0C3opjBfCU+CZlQrnG//Zl+NpxY1Y/qCFuhWZZszY9bgL71fia3iqarDrbi
S1u+H2y5XB73mdiY5C8caflgz24XfrzAYjMFEDO82dDYXHMO+Jiujx+5PyMzOKuc
r7uxLDhrHm9UdOKZ046s8Eafd03qEEHmnv+eTdm+NKIDE2AvRIKWPg00AxwkNBcn
wxQeZhkSked7llaaAAsvZJ93Yxfk2HAKvxFO6zeNhkKaYXPYPCHwPLcpqeVqi5a/
d3VpyqCk7FNUGYU6E5p+39l6K73zHhn8SBu+fMHCgEh6m2nT3vQZV+jF4JUG4iZG
3dQQKA2NpraoGidgKoR2fh6nW3Z0yEEfj8adMX59gyQdPw68RbZQ42+D47YDAw+i
xZr2086mkXGg6Z7WT3EliCD6RbU8w7uDppFV6ez55zNUDDNqt+wbjWYaak7H7DXV
fn5O5gfIxzFecyZCesIHiuiTwI/dR7xKCylpeR9wZP/chehBb0w4jNZFB0GPIe1Z
6urVi+4ppzDA2BcjA/2A90pcEm3wgT1yKjLG0vwE769qzuWFjc6TOOY/wSD03Lgy
7FbqP705FDyR22eknn+qHo7u3fEvxCYc3zS3e5LT83KG75SCDZtRVy3UzgRnEAjx
FNr4eHrk4weMxraoY2fDp/Fl0EAVT2yF2Cqysz9oxxhEWvbqgtbNLfHxMFz5cOR8
6DQvwy/TL2iWY6Sx/gPivIsoRTPg4fFY/50ool2vjZ6hqZCd51Bc49QqrJhXp0Qs
vftEXMaZXupuwv3hxle9dsdTlx6+0pqqP2ysmE7wMNG7FpIgq8znomF8mllm2qss
qwzsz4ck0POxkBj4wwf81PaU2WEspaVLeM51GYWxDQhQlwgTycWl9KG1Re3FQAP6
nkUuWLMpN/xKrfJ9i9dKg0rv6swz8x8HHkZ//41VtkyKogfVveK2lFe/Bh9gF0ar
S+Ye2esAvNT012HlSoeCFdKPFUaAZOfC8jp5YqYr2RjsPiuCY6oZyZJR9aANbIT/
naCL0g5B3DU6EuDdxHTZJw7pr+NmfKLfqVLTIjvC+LJDEX7GI0yGWaYuMBkJWlkd
QLLGzxtqw10+srPx/wkE58UrUTHO1uAnt4AQpex1mC+WpJZ4uvpMEQG4E8RANNb2
zGf0o2PugPDCLoybCum5KISwhQYVDT4eo0QliG2smrm4CHXidUIs5dygOjcecnyF
bLfuq0UQ2vMXBRBlJ10nxTCcjXutbbG7TYhGWZCUUQ9I3L4NFNPYLeG346gSWStl
y67VU0SbtVLely5dYXjksUB1x1tPCTvlwiE88qzZa7+RFSjANlLcsvIi6s+dVBl5
CkmJUWgHzqIE3SFTGQQGriMmsapWjYKvPzjZk9XzKNdzEgYamtBK6t4xHgD8IkUQ
3IIyNtfj4jvDBGFCqTkFJ+TuXTPD/RvRG+eqYPnPzOmucxZ/ZP20entCt1fZkMev
lZNEIw3phyj6f/h3ACWxCE0+fx239dVQCyl2vzvmWq/JiWyisPhXN1lIv7aSnAQJ
qea6KzjJ1GVetSOFUTTH5rt0iXgU57RyMe4GSL8xIE19d+5hZcEwlHpbK9XPqU7t
KClGSc+wK62Uw/VPIWEBfLXldl7RW49BrobqXM8HSOYuBaI7Eypui6Z511KD+mjF
1LMhDjfyDhP69dUl67XQOLQIs7A7cXF/wG2NrKajRFgF+C1hHCngEZndO6crpZQE
MD0RZkY9JE3J7MiCyack+fmDAUYjdEAjCD9Vss3ZjU+jfYDEgjd5cE8fm3VsGVEw
FXrnpOJWq5AWKBocfjcx5vPgu6hX4bAvr+7Y0xm38HJQ8eZaGpVIrcyb8WehFbqu
z9SHZxjnjKf3xDXoDuuLWVJ3t4D38JqXVAvpBOmDz6Lgg/N5iv8sPlqeECnemQAm
sXl1Sf8JeGd6mG/b0EKSwOSVH4p7AbtgmWBCf4w/a3zgXkIBzqUjRIE72G4Ns6uq
+zcBjKWa2HY2zimgZkFxQsPmygoHIhdWxtJwb78kzBPu/NaQrHzMGfmqOy1m7R+P
fkEJaO6nAYBQ/T2fLsLsaY68tjHcuf4dR/R3hbHBEjNbhY9EaWee5NN5FJyacod4
oGLZiT5g6d+iLU6dcQae+aN7klPNmBMacjG7SjdvYE0Tiz/kTsRw3bGTlHg0LWHI
euqIl16aeAzC4OTboCPj4q9rcUpArKk5vUm7wPkWHjvxKOaZGThenkHNI3YCeEAu
3vzKu8XFT/8dvWiQsGjzngNJR64Hp49F+aah8F6CFzVMyRdLMfGAeeEUSIQ7v96s
/DVWZlLsqHhyvOlbQPYxE52PU9NoUar05K49OAj+aQm/ct0Fzeu/xmHWTtogO6Y6
MYSD2dbOSpxrIImIgq0NEGMmqrn7oTpw/cJpkEFqvJ9TTgJrMU1/1uaZopP88jA/
mlZdHjkwJyhNCCGNbbGzxdWGhHpOJi3qP7gEV0Ha90hgUtgEGEo35p1KL3kuupK2
5QB+P32aWnytXQSRYsKezM7RgCD33LZfwt8ZVcA7IKWlt+GkQwkF9Q326Yguo8F1
aTsAkd0Gf9+Dd/5ODLZ7Jf2ibiLqMW6xDH7KrrOiFp2GuvMc3dKhstFE5CeuAKpn
`protect END_PROTECTED
