`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xgRyBA8biIGrQk9O5fCai9XJ4JFxbaUrtUoW6Dt6bBbBK1T9lwxytWGWgZhdsY1k
D9dRZWD0k/lDJg01CVFe1f5VsDE6/jqBVz3EBdQ1eT6O/QAaicjY3MyTAfFxgysg
gEGVKXx/a2GAabqWXLNlz86Actu2/0rkhRkTvZSzAndeq8evgdIkAzQOwmPdx/0G
+dYoYjFAyW2HhNHCZCdcnl05ONNbmUyGISBwjpxJv9bJsiXTpfLZXJOXGv+EYkLo
vamsIjQuypba3eilVRkvjDC8eZqnD7u3xUyumCespfqw5qjNC9kpf7s/CuMk0M7s
X15CSZk6O9qwlzga6ciNQ2Mm3TcNuAtCvAURqo5RW3I7oEThZUDP6/5vlGYkIpi2
aqt10NdH6n3U/FFY0Le3yqRPUWau0TK3aF1AhAvkxiaUT1UuKcL94KxuyF2wLTW0
TJeY5BIYAnZklNwLFo1zjLHNtVWMH5Ckgc6UGEJan+gzLshwzkEB9jxTLc8AKrfp
FnSY2x36V1oX5hyDRXn9PnYByf3yg5dKT8gQr5cTkxtrXWLIp9AXT6cQpKsACMrb
+MVh0e89PuDesxb2VtQj7Sm80U6hTQJrBm5VnqezYj40y2J9NWMhVpRcgeFf4wPQ
8Aiii60sQ1137AdciBhkD/auEeblLs/4dzJx3SxArKsZwQdF6ra9ucz7X48raqyT
UWaiquVUb0+1eVqShj93IIAE360cAYl+1Io9/t8Yj4j7H6udMWQ60zugmx9Bz0N2
InoqKYmQ61lO6oCpzIshEf6IEDid6yDhOMg0bu1ZcRKZfPF/HpzeS3E9jbnIy0Je
5tjmNhSFKQ9TMNb2if4JW962u1QUZLblFvl9r5+tJh31Ma14Xx1fptl8PEiI3jMw
P1Q9H4+Oss2bPUIVwdcynbWDEgSoCwhygZkJ/5PzPpV956RmIJ65ZLu4u1/bZLGh
e28G1iMfG3qcWjpJraHoNlnnv/sEaYP2+WT6ONz8e5mTBlT9zfID1cNfq3MRLKf+
sxq1waJk5SgFETuSn2+A8x9HT8uU8m4UOUGCNQSxLtgFOLYwrPZpssfz6g8O2ciG
4h7LjbF4fN964D6xV5/dTnnWsJFSF7nJH6/TtudALRg1WB6kocZz2A5TxqVtRA1G
DYIueMmOiVtmyL4cOCmqZulg4oc4xwoiqyBgnZNyHCFvZhJQuAG20fQfJVQ1ucLq
8v73EWCk8pnEezDTOFAlkFOmqJImqSxC52NFaQqurQyfmbuHeUaVrzz9qBVGsEKa
rXm+Z8lJ+WoWkdL6cn9VGL9sdHTlFQB2OPv4N/dCnyDJdH4ONet+xys8lMhxu9WI
Iv//bYFi0yfH3xIyHCY0v5cV2+SN671iJOuzbfg4TCqhUXIxHuesGqaq25S54667
txlMhX/zlF6q3GUay53BQEr2D5vaCKnwJ4/pQzuACEMv7iBtj9Iu7fKERo8FAsvE
5v1yGPI8H/oDYhHgkufJhJ8CBPgnOzzm+EicN9Vw0BDl3zF3nk+xIx1EBVTnr8kT
D18LVNebGhBbaN6jb4B0qfddYqQWXhiu7Pw95uwksHHkuCgVlcZc6cUWabMliWv0
p+4JOVfmbmmH5Q6uVTec6yZyFSROt1t141Ng6Oy4LhikcYYz3UMAFCmUw6nAIYiw
qlRuJLH91tiU0iTzc9h65TW3qtjCkpC/pYgSP62GwrLW/MY56g+N42roz1wZ7CWg
NBU2tVmx/WA9MVp98FUiCvJZ9IwRnkozXj7WO01/VQr4vXUgIJAb2Vn9vklLKxar
hmMX/IQIdBTMl7zMr3002Ufn8ObtOkQ0oGUfTwi8jBEvlOymsgTKTjDkmbPiOLVC
4M8mbyxC11EhM+jRy07JAtPWaR8m6rbt2ahTN3QNl/KYLcwe86jKnD81sFCqO37Z
BpC54fpBXVtml4tsJs6vof/4XbEasDe6x5DJ7Jj/++A=
`protect END_PROTECTED
