`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fA+u6r8LDyoY+OhCaHVmQgHipGhVL/lCLaApyd1YycLXY5+lXgap08jWeARLqA5M
stU69TXaY1VfZRUka9JXVc3kmAPnaLzkKNg+6cU5m9+7I1ySWr7J+8Rj+GcAi6xg
qzMs6JuRP97UA0yOvKoK2cjDwi0wX7Z6gSE3eOejw/UFdhjNYJUUONV15QeZ66a6
XMpq8gAGJXBXhVIlXWUU84LlE6c1A0MNYzl1pkXmswhgXTtVZFJs9NWDlkxhP7Zk
iMGnqxUUKpLZdbZeeZcH/FZnjvkDwk+V/Y9LkiThA+AvJMnbmlMfjUINYQUUmAd5
kRZEYdLZ3mmGKeBQNUOOy2xw1aQEGaLdZS9nffrA2/uSmbvUP9GV03c1GG66FeKe
cbPVDGXJfOC0gBIhHN9HnsFw1DBMWYW8XfOi9PwEDdiGYE4ntg4rc2Nlc9Trh2oc
8vaR1DoXxgnzzHIFWq+7OHNlCp0DC7+r7b8j2bc3Jm5d7U0FiAB/Q5htE9Z4USEm
DxCoRmgZhpCnNS91/YmIBO41gLz6n6g8d/sNXnleqU9QDqbdXFE/qL5CVb0hFzua
M+22sdNadK9G3lewgpgjkg==
`protect END_PROTECTED
