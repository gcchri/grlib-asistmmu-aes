`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wtU4PZ7SSIhkMMY4dHdtvURq/DbPmxbJMr0JjKaBjk5zd9+vqJQTY5mmlN+BMnNq
T/pkcs9N6Ub9/seAxytRImTeq/5cqhD7uNTD5w7vHNOHB0sp0YyKQDEmhPvZFhN5
ayTWycSrzfeeeLwVGM0a+HTx79ROnbkIb3YFfX/i3j18QyS6NQDCOBOTm0sVvArF
bD0igoG3jZkujuIo5pARoLZFo+pqFhUAfEQCswvVsfw65u9HU4hEbTPQzuIgrgSH
PSloyMr24OV11+4DMDMKu0qeGGTxj5SBebTdVuLhY9tBxJ76/sA3qv5d9WlQsw2t
er5OzWDzF5q2DIzWZYgsWhY4aX/7iAYh3XDl0770H9kzFxE/8qsRttH3Si47aFBM
8isKnJUfN6D6LCEUN17TMki93WN9uNwAlFtFTJMYCSOhn/Vjyf7BxPttcHlZ5NVK
OTTLnEcM4P4cHvcfaORXnCfgbyCFeaJ0sbK+ijLyMlO2cKhJ2jrWa4t5ruzh9eFj
MnqLsICHsbrILTd/+TAEHpQPLCc32ptks7vT+rpv0/TJd/MA/K+1NmxljamYm7c7
t1l8XznRQl56Xr3RsYCzwOESwGAMkxfxfHykXmvAaip8n+pmbsoVCO+zmijGH5tw
6aOymgkuq5W78Q3H3PYtfW7hWrmUQuPpIP0nvQXS2BcrmLr+iHgdEzO6DbueHIR9
8QQI6xCUMTOSPOv7xvMU4zju0eiy1RLC3dL+pVLQafNLU+s8YhqVNAfSSbqQUhTX
vgvXSNkqkI8naPdL9dNyQyggw4K4dX3r92JAS86Ic4LEiWDSlDIyh6PyJi/jAWSs
C6WfMG4TUoi8mBa+qH4i3j4I+8+THBFoZBzJBFPUs2sP2/xiry9E3wGGOoGa6vHn
YQlrVIHotJcqw+90e/bmwBsLZlry/hLcDW0lm9oMX+B9CzByScpwPMKaG1SsKa1c
v/f5yob0UKQ5bgVFm9+IghsJrKaRrJn3tnJkkOTg1BW/PwItyGc4m9K07sYdBYFd
o+mtZU3Kel+Ktsznr6j+aFAwkXt8OFFU09LkhQzvflCQPn9FFbeV4ahyB9yL3r1C
HgehEPBTMDp+tuJ6Lca2piLtoAfIoQYEj/4nK9LsQ7k1tcXnLx26n//EmIsjUxOG
n8trMR61hllK/CQKRjbqK15lxPh0cSUxsXxTbHnNrg/Cifv2O40msscOkGdMLIiW
KC2fk8CNDLSpjlb6oi5zp07w9qO7d2eQrSZbysSbcvpQeog+pFj31P5mSHm0MoQA
NxuZr3DxfrFZcHQVRS9i7vK/wv7E9Nmt/5CS/9NajpBgLi0PkWmvQZP/Cvi2Y8Hi
zZOksxaFp1B7UI2affhhbfZ8Ni0rc0Ybnkumpou1599frkB5qQF1ELA9ZwlHB23t
46znU1XeFwGMvT5btjm6zKOkRUvZIO11inqxPBgwtwVlhbuxnKk/sGNa6CxvAmRB
6VbJ3jATV0ztIPzr81UbNs/mEzNWIheizLRoZds8A8Snb5aLi+LaDkJBxIcA9Jc1
M87rWm43UG2iIKx2sPBfXnLRnrDnp+Sm2r2EegRu0H0UAEWB9nxMfRGVL9ucPHSe
wKZZeVGki+0YJe0kQ9/AAbaA8t8kNdZ7/MXSlWy6gfs5Dwqp4e5GfEOSyQjIqRwD
sk8DcyqLzaG3wUrrEoiI1fcLkKjpzgZb6sYXXsIoy2EvmUTknR/+bGE9++yQKaYO
ijatDudAwCjhv9/52tlacPJv7j3YzFWSLcb+pSiPv6Iwc5ZU/dak3sAc0Qad7xeu
LsbtRz345uI56yZMxDdHloTC96mj61PkUQEl3Yfo8QKEK+Z3BOlVWNR1DNHgea/m
0Z8EnHCK8khK+/DAEjp44JEq+gnDY+tpfh+pnEAub1TAVPCDTcFiKuc/uQZ9hvAi
11QeMcYVqf9FpOoEy37/Pgf2wcSrtCFK+rKbdn9FrthCcv65iyPOCUqV3ukG+cxt
ILVdxNkye1agg1Sgj91wdWG9iiOdAqBiQUp7wQB7zUuVt65TqA1z1UrqlEFFnVGr
hrwO/zZSFkcGmMhLCzEPKbRNAPuJUgqFsqO90AHyuL1l6aM7JMzUhF/XjAKVMdNN
McapaEIveMLJbid8WbAoKSnoOIt7UiuwaImcxmaNmILfnisSX9Fc+0iY6dQ7phWj
mjkSjyoeLkti8THqq0UMYXSnN571nbKghzB+QR9e4ETzdnMKAtekJW4XkhjuoG9G
vTf4U5UMF714EmXngVfgTIZ38lR8FYs/TsgFFirCCyM=
`protect END_PROTECTED
