`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nqXApi33ujFeDKXEcxKoODcG/kNGSGzr+Tf29GwjEJOlnJJZMoCtuRMqsNndKnA3
2Qi2va/oamJjGCs4rWdLxJ+MamDntcbsWdWVj5MMlvj6Hmhek4zm5HmLpoHNeU/v
s7j3bVjpzuzy/X/d2ZQeLMEoAPfYaWQ0AF5mGTubudJnnzNX2g01OByfnwbHYDXi
I8Eo/mLINTtom8gdjwO4Uj1jtRv/PsUZh+ngOYeXer+KV+beyN7n1PnzAqYOTIKW
`protect END_PROTECTED
