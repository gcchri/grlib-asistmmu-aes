`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ctuUPepFDwLrkrrXzKc1Ctc35LSEt7ws0ke4nk3LcJTqCEVtFCoRtioVjWt4NVzX
9nsF2AKc8RXGojHvmEW6j090DK4bHO9qUwKnzkAubfL9nL+kiXYSTCVLPoW6v/bK
1akRy0W5oc8qcqqydf5+tZCQgBwzY1ho27ZJ6tTKqyeOcbeKjDXDqWod2EKcyIHx
97t44IKHx6Cyx/dcSCXBhSRYjvK5PhsgJ4cvOLmv3HCSxojCKQf7d2zoNWfthzzD
Rya2tHOycsls52hzAeNS54OTWPPVdzBjoW4A9wBAwOWNzvjFh/5At0jqLL5KBEBS
fhKicvz3WsmwXJ1ZsXNnnUkHqZpg1RKWbCzldxenTL9XqbdBjLx5MRLhDzKgbVvd
+nxO/hGTsUqKfJp/5Iena3yQKw6reOlIJBQAEBjcBtY=
`protect END_PROTECTED
