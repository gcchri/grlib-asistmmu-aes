`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5zollQoHCczB/C4A6N/ShycXDFyRWr/vhAAkSdaZeSweC4K9RAU8h7IQR/MfLA7x
AssuGpnPTeux+oUZe+Xu45WNYkCrkIEHXcrILxbotOTjQ+tKp3s01XMMJ+CI/Ag8
nZnVF5d8bVSCGgyUAJciPfV6U/930L9f4U2GSPB/EExj9qvXLrA+VmgTHt70EutU
nQuZw7ChSJxRT0hn+IDmRPNVZdNb043PhfV767W77JOw4OrBgNK0EL8+68rAW5ux
ue32MZuI8lim896DmgD4y3/Pk3/c7Ohs2l4E0Ou9R5SbqsoiA1/Z3sKeEzKfG88B
6lBCTZGim/x1KRXHorn4OcEnVpvymC2YAUlIR1t8kVikpI3eXvr7zU+moeXcEbxu
XNuc+kyqPezc21qIoWBora3NrfwQbnXVJmgF4u83/fu61mzqkvbhd3hddwswFIC9
UiB7mkz91vT1IRdzD0KkQhT8CRkiD+11fplKuiFI9gw=
`protect END_PROTECTED
