`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b0VKv1ZZga3IwjcLIASFamonUwyhOehpCHTqzOTOPZgkuB+nJ2d3Zm+N3kuDy87t
a/nGu6vw/CuSPQIRWYbukb9eF0taeTBs0lF/3KwgiVw2LpQY5EWve5fnt04XMtsS
2MliRMQoZHkpB3/+FycGKbgECWHUyRBG2sGNYbclMcVF9/MDbf9emzIKRiQFujef
oIjccBJnf7LoRl/SxQ0QDGKlFfG9+VWtOYKoqgYwR9fIeWfW30yTjM0M7opF/Eba
eX4a7NiSMenVXRYCjPfNCIDWoX69XWfyFIGqHZkP0xudDENCuIHhbv++RsUlEU4R
gp5a7rOAihQSflTNKMR0Uw==
`protect END_PROTECTED
