`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ng2OAxJNpCQepZDnv9faDSH8yoFDF5K9xqQMiu637AJPXRM1WIZfMxcEiORPPTw5
gOElZwhz7SclpHZprwgtz+6EOt7/uuDwZpDptPPxS2cM6H9gUFfr00hao/xEbkH1
Oz07J6dsJOfbms4bN+t8hQmPnD6w0pXdzfsGn+6o5h73dfkYGhSo6zyF/KN3XImI
1XxJ9WkISel8VvDtMJhfzui7jUmecO6bo9HbOBdE+wqFy2ut8MNJJazqDBmoSnov
0GnOEJFMLy7VeRPlO8L8kic0iwydqUf2E8LCKCUZuP6TLBLmE2APERknw0PZSQ2w
SLXKYUXPBma2e0DaABXHf4qv7cS12hnSTJItix74UW8UJ2ZSyimJ+DXDCNCsfp+k
LpXEfQtvyXaDX2i/uXKbfQ+Lvr59f48ouPmivzXm0zGlkwWKammmrk3W+0LZibeg
B3T+zU2CxFiaZByo++/kgOGqeYkIONy61dTIgwCOS0dcuUU/oskKBPNYxIYzkb+J
+XLwSD5UuH1B4SmBsOAfxjRRP2WAQd4oA+DGw/AWu6oxwy0CUY+EK3gXZWWG+7kp
ofTmicPmM4Kug6KvzdG9A1RktT571Almq3ww+HtQ8/bITT0nT/5hrG4BsY8LL4Hi
z2lcVP3vsPXjNDrdNRMDllfjML9IwRZyvLNydJH64eVE29zgh/Dy9pnFOjkjni+D
Vtj79lzj5QCJn3AeRKIcgVXA5w0QiNbVUYBSLo6BYx2Z2jBfTobIyKWMkXwQqQNi
meNuUD8U6zl+DG4odnAu7w==
`protect END_PROTECTED
