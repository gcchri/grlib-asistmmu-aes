`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I1b6iIscOBFYWdse7dhF4TRiYcepbWgtime0qKDtLcQYv00yr2KGRgO8FfDPV6gp
SC4ZcZInqTStaZxZ7IF9emdIdCYZAt50VEAw3yTr4p6eqPRvKLBSFgrbYjNrcL6h
feplL5U2hf5qYdxC97KLmv1/uejQJuGH4MPcifrCfYA40Z5LHgHvIb7SW3uwh1D5
uu8S4QKbc+SYEXDOR00w+uVhudnF6Peo/3Nwk7KpHDxTLF2Fom8Kjf+WNc/wwv1Y
ZZbt8Cp6s+kArQxtCTxacKBpP+B50yORf3YYil/bxzSL+ds5uOKkVkM4fpKGbsGs
x98w6Wqi1/xKS9y79bq1cpfaANFkgATIoaEk55Uvn7VnDS/xbPKkjPmxMQb5vGCe
7bemEbb0TmjtEdNGrB0xt0jDxI8TqlSyMzkuWcds1aGJYcNijrHCPwUgGsXhgAb5
iodZVX0TTj7+YPoMnQHPYnk1nZcdgVISn2ObKVFBtzWswxFeeoU4dmKGfHKvIzRz
yaZI4rqP3X0vXnlS14zNpKxWwlzi8/DbIXxUcq/p6MFP7e43PYvuP1lnTKgCX0kW
Dg26Tne/gsfHZwRxtYYU6MipjufJx44THGQbRf0oEusyN5P1SCKJXaYKPC8hCP+S
nAt2jjg2j1gk09NI3jubJDNKMhuCKRWqUmamXJh7eAluCl65ChsJklxiQ9LMGIJm
`protect END_PROTECTED
