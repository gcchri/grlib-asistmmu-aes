`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jh+jo6gd2NF/L8Fip7KmcSf/ZPQcBWK/ex7TgQqVFN/OWONDpmqt+zDRkUMEdlr8
o4BL7rri44hinl7TVEpUD7fmr2IbnkeR64Bf/q7uW7TojOqojyLTyGHqY6LEKQSn
rsdSGl232aK2mhC+0yO3Aj7ZPa4lKG1B03d6Cj+FujDduHUbhZGq1RRkcxWnF6R8
KUETQPh7UWlrMPQGEyFekm6AgfR9TxmRS2NErv/tVM5WWugZ2ivU98bRr616YCcn
rgZzsDVxzl/qrYoLNhlnNvZ3XONwUpDTlPzlSEadjCaW4E3h0tStD1eAXz02VGLO
GdwXN+tUf4MMtOy5HnutrrMgPP7EnEopy9pCpmpQvA1MtsWsg6sz5mdeHS/+aPLT
+EDytJmhZxBbP8bTZd8evHx+6pN/5oXOFrT0vMQ9Pr8yFAf/jbNAKuCc72i589UC
Jax9iDg55z/YbYGpJpW4WwRDp9MtevHcoK4/bQMu7+AT5v0KwVSLYlxX183H+u3T
EsJThR2p8dBgeONvxmGbAkVR3t6UG+KP4wDo8BebJFSXGl8sLm0QsB/GHLvju7fo
AadgXzxYHkmoarAlbUHlf9SoHKbJNU7y3rzJfu/x/zfP5GT+4x2AUOJ2LtvBsdVO
cyEFJqCHnBhlTAkzaQ6WjqkUNGaa5pvzfVp9zL8wx76X89YmLAw990r5rTc4YQVx
D+Uytvd8JWthYjOyDFxRxsSZKWXjW921Zmqy0G/ylOP7MH4zutKWFzuZJs4ru7Mv
ELeNbhEDOgKvsXMkO9ncfeXSubMXZ5m4qEx6DIp6VRIOyu0Mc/NGILVD7o5nTlog
d2sPiFlYENy9GZIFtuPcc/XF2ke+uaxG/Nkkybj+WPkVt3eEzcZ0BUj6k0LrwQlP
Q/sOEgNM035q4/qVwHD5ZVGf+Nos0r6VpJVNchnj8CJqPCrbItJCANY0ZvKdpCpl
vBFw9U0j/tkqLwo1BjVsmAW2YQE57aTR9REY1qKEovFCx++FNczpd2crzMMWYycJ
YlWMrC1DI2vFGkl0jpLiLjUHpWkVGYcN0+TABZChI6p+UKk/YcsS9yvc6+84zhLN
Y7HxMevXznQPf2BBE2bDUXWOQGJMyontsfLgI+035kQG2G4y13YwIxR5pGX6gxgZ
VHNz2QbS6ulrooxjGaR/MG4HrrXaGBgnouuMC3h6XVEWQBQB0qEPhin6UKJfZwE8
8qto4WwxmdKa8VSWK3yiuiCgbXV7OWEqWhtAn7pfxXi3G47H0cDNbgAG1JCvIWl1
UUbo7IvQCUxbP6SDAuE3mgvCM+Z/xPF63zD5sIW/Fn5snzVyduVvmXxZ6nDgmNXV
CfcYBVWr/fbk2HFru3PoM3gJYdql9vNivR1RE/f9milbwOLznSKSHQruRQ6lVKiJ
v8xys1krKs28gPjkXXElN84phQPiI6M3l+BjWlCbPaD95dhwKChuSHJu8Rj5YNfn
5XaLDbDfX9iBEpxeWAEeGs4+7mZO7l4XopK7yrWZlcVCjy9pcCaynA0cfP16pZ1u
DFxTF65LfJL/5olWY5Beu8FUH0hrvnG78eQZOMej+5I=
`protect END_PROTECTED
