`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LEj3AwHiTZh9dtoz5uAfjC/Hv4cAxGVsKerfg3IKK/tUBm2kfJ1Pn50AjqER8PNT
WojBEMGG5SWvL6G4BcQhtJcAJLa1/KPJZ9O2r75m5kd6tLmJthjfbsGOvNNwBpmD
gt2umL+wV6nxoChdA5uK0jmewQhWMADxsdNp4e6WqzWuBAkVsdDik72LH8p7e9Vc
GoQX14IeoSMZo9w37hzqmK6f8zFvCy8Dh0yWPkd4PQFbKORqFHFUuufXoI/8pxm7
plqjUxgb0tpDwo+X7YVfrW7beRRcpqX2rQgCwl8xBy6Z78+WA0AxE1Vh6K8IgOX0
Yf9LZo+2TycT0/AS7WcaOYulYM9BFGHztS5v2iuWWANXz8g8ZOUIArVMLxvrt/Qu
f5V0YeDDLZZmWasqNRQhqA9ApA56H9ElSb+PnFegc0UE1IfU5pgK4F2/T2JawYnl
P421MomOpT8+qvZO7gPVng9m0QGGzDO7Tm+7AIFRPFyu67/jqFqPh6Yltl9eHzye
t6NxNi63b3Iqo0gsp0mx2fb+FG1M+VnAjGVw51/JyEWegLK4T5CrE2FMceWLrhdH
EviCdAlXHuKKdZe+5B0NJM0EYv7J1f1qaDbInP7uOjXrcbdmdB2udWraIJzFbDVG
w2M25ylRNxECemPZHRqXxEqXKpH7kYVTYG12XcE8zgtDH1voNbw5Zkydq3R8fPzM
mIExhRx73CzSlo1y2hxLCh7P+AYVl+nWIgg7RMpbprHzLnkLpWRrF+tEG04kFCho
AHQLlnLhoUPOQ6rWguTnEOvQtknsDq16ZecJdgDBN6iUvuAHl/RI040l3M9A8/fb
Ks6HhlLWKesKyls+nPzzmhSMyb/Arhn5yi21LjPcL/y3IkgB8mFEhWXXyeYEHsj6
ANOjSkAYXU83BRDGgzZZpg==
`protect END_PROTECTED
