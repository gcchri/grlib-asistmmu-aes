`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uhSNok4uI9QR6zND5f4aOEZzz+RetJoK+LB31LDw2/ltgk4ppsYkI8FrktgwRTwi
6v1H6vYgENP1LTECMnm8f/uvoLIq8+nR26AYAqYhKKPWhgBCGN2wBo9uyB3RrFDG
ORHNFVgKgcPm748SIXf6SMVgugdT7OqoIfgH7IpWacF1AfXTwmUVXLt3tlMZXDQo
F5dlLH36QHE5p8byvLLpZq4YCVoccLcwlPpoYwK1uKVU2seC9SOFnEGsWGTkQ8jO
5WvbrFo5cCZ1JybWGToPDF3V3C0EVOR3yjmO0g/Oyg+g9rbMqnpyNKCbmPuh5Ogf
Q4G/weEs8Sg7woNuD/3ftXE9QgFseu4vFID/42ZoRD85+tD22iZYvVyv76sF4HU0
Xv+WkisFKbhUAxsbNWLcqB7Bjs/4cLv5q73UDAPoMjQ4/vTelb46z6iiVdcVZuiu
8eMSPqKnwuxoo6JFuPBn8YDmB6mekAzsF06zMGLcCS/l7dHO/kcnjvcJoKrhLCJK
ZDmjEYv9E6UFjrX62X1I4Jtrka4SiSDw/HbUgjLcXs4RbihitQUhDKpemE+1E3/l
16F7La7V+KvWGwWhpcvJiw==
`protect END_PROTECTED
