`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F6B1Zu5Vj7ForsVHxH9Vg8pcmz7Z72HUv6qVjGd/NZG+VBHzbc1FhrLtfffXvfyu
7vxlVcbooRqdSIxavF/syfZmNM9HH/haG/fzhyBzmZSuYidRze4KGEon4cVp4o5v
eK2XHHYeQdVlHdn704Gt7kHodJPX6K+lu0qpsc9CzpdqEX7qbB5dvwiYrBuP+db9
M/mzJ7QWfA77GlgVjmn6UHNuOLBrXGwA+n7EoLTul5Kz6L4jC1jKbyF5rOg+gSg6
aUkDrxbzbl323RiA09W58baKcQapOhKQaRLsjRRis5LQgY9G0R7P1EWKk4ihvsD9
Ka+ZGPlmA8RxUSnLgyLOEGtZesS/KCltT7b+ZKOseHG/bys9vu1pSfiBOee375R/
Ym6s+MmUscTigJCnG3yprGt3rK50kDVwck+eUoLgURzHCNJIA6btfjbcsubWBSAy
wvz4dG1wkG65qUdt3vcyCafpWslNI5sfNNq3QZLqRDhey7i5QcStm+7sqezgIuez
SPPEg2iO1ml7buS7kiYuTVV72XbihxqiNNTfkRKrVIECbjCJXVUFk83r25YvYRQS
syEMs+01Rz4Oj4inj0fHGdvW9VsGefvoV5u/V5dXv8CyUbtbGBMSRhrymfzPRrDI
HlkeBSwlSErHprjSonTYgw==
`protect END_PROTECTED
