`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
skvz7VLGY2MsiGG/0w12IjltkPo36Xl+WdJ6nlsTYU0AcWNmtvo6xYyz1/C2w4lw
yGgQPtH/GRM4ZpbEduHqqqxxQWgMAJZwRxwFcoTYT7FziMCHy/glyhYEFNuR5WS6
GJNi3hJ1GJ+TlhQ6DkplG312FOgyKVoT19dzUVXtPoC3WJ2fdvLSMyJETKvmK27P
LaVIP5DOBaObpcI6B2Ci3xrQSWptU/BoCWH79w90QBFkYoYgrFE21Fn8J2pjHs6p
fz28oopDRnRRQwUmIdPD2vmkB1r/F4HcX1j+2Bp0af+TRC2PEVzmRLhzQ7x0SRuo
aHUabfPuXINqEjMR2FA+vA==
`protect END_PROTECTED
