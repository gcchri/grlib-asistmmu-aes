`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xmwmOiNBtVJBHiTjUhTgzwVL7Y9arxwkMurwmNQwv21pU4r68/jlqOiN83MVCTdy
ltVF9RBb4pLIhcapUH8mlXN0MfYhYCiwJfefp40H5dKmRMFTEXFxVNk6V83Hcmwq
n8ACOYZZbfDeSVEWNz8wv0w1mQpZoI2xnMpgShrNxuIemoaQp2LSk7cpuTQ7E3Ke
gLZdLhvaapAA6Z74XCIWjAYsqlG6Vca/WrK3t02y4NXac3a3vgPYINTxSfD8vGBD
fTpUKQump15z5heyrqss6/U5hjk9qVNDp4OuyLmCDMiGIMwKj+BOgk2OMVnn7PY2
1QZ30e8L7DciAeUXG4qyqDqYW6GEH+7aG0FXOnk2h0mESDm9ElRsoGGDBhBnqpIj
HLLdiGEwFE2gM8qFohqNGqNB/9R4ySdRgBdWRTGdTs4=
`protect END_PROTECTED
