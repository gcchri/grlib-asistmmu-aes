`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gy3GTtI8VVKaTSycZ1su0DPEd3Emp5OVp4eNk1XRrP48clpANyCc0ir1ufuqhUsZ
oNhFKFYsblLkrq1uhp9a+sroNvOvu44ifUQfZ2xHSAktvAo9/adJ8osExwTu6r1T
rzvuZyJfOaC7UoDpigCVy1C/62H/JghN+XU5vCVwH7QLmmroSiCmc9iTK0NmMqsd
smMvTNBcYgaN46N0GMF5eGIiSQjh5ovWNDm4dsJQb2GDNAEZzUO48wCI1OgIU4wy
JcsmTq+M2FPg7JeaqPXkaNxL+rBb3loAyhxxJ8I2FqjQe/YiMnIRTwihAMYpPo2e
/bUrMqzmt47K73wjoHCe3AFYJ4aUejhKRXfFvCgn3TMBMy33YOa6vvj0wjAAXmD4
ofG1xvfbQcj49LvZKRjwVYfRV8YCwbLPsO9WgMaxzUrkWU+HmfWENJvR6hZJx9AJ
ida9JmjGfhUXpIdJOZ8kuXf/S+L0HsJbAwsoh/AWL31GRzLUemwX77D31Dfu+Gk0
/Li/uo0czWlo5jRClNG2eChgmDL/lXzh7lPjhmVcUZ6CaP7PPPgnc/GnDsj/rZ3T
47ri6h6KIlRAdp4loAwtiLVVqwj4TTREKoKmfY3BQipxF9jw6BPmwoS4UuWTGKJt
fDby/zfKa6jEvZdko5VxXOR3E5tZHnUQRfgg46aDUhPjuz0pc9GEVx/yvkollpIy
sFUuNqhoc3F1R5R+TAt22g==
`protect END_PROTECTED
