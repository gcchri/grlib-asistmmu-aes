`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
53UIlTaV9OF+VotRH/XdoFIx9uXnBQlREOolgEWvgW49QeQpCB1SedHC8MaXcMTi
JB6KLWmMKqfsEcv6uuXju47zsP9nJdNXf3rNkq7Xs2JE/c1PhJGrfQkYePBmCfJA
uDfBH98/KCzi9bp1MJFZB9/NWpo0uNLr4z2KNw/V7CtJS28SQHD4rtyvb3VCHP8+
DQqvzhcYzYuy1YoLjVV71fpokKBzJf+fVxSyv6s8QvNYWtpniMMEZ7uhICPPuddQ
KcPSHtM0G/ljnP3141rdqvofnZ0GC7KQPTYa9Azq8DOphLhjLFcRfoxqJ+jmGnpG
nU4xLWC3cLniaztImTGy4w==
`protect END_PROTECTED
