`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WGLLIegkr96NaQgkOqJ7smwhVHoW7dOOktJx/4heDWzIyP7AecBOqBxNQZhC4uw2
Hm579iN5Ib32czdzihjGk3ebMHXbG1qOBGxdtIFuYAkfqVtKsx6v+HjxoAZTiiJ1
W46VqYCVQZaxdNWsQZP+0AI/vuyPltGmAXmUxwobFuoUjnOuybg8S9FD7NEwtTY2
R+5Ou3sGNIKdkKCK9xRVzYUnCQb7+9/KaeikK902sDIIPXCv1OApFPsy4AZhuMZq
17M1/flNTPmMZYb+bBvdzT+foX3iiEZbU9xZobf91uVy+L+lhGLOWDHGPToHss/8
LcOZ1sMnhwWNvQGadgA4GSwRqj/0hVvOksxFKll0sikOj1igTz8sJ37VLTL55TsK
ufMF9DhgK3l4rHlBB1QmlIqs9IJtDOW4vor/qA9Hw9SXkaD7o3e6b4zrqsx08NH2
`protect END_PROTECTED
