`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n1l3bAcYfQQ6WRfmMKawEicFpcNI+eNfo/E6UM0Cc2JFmWDiELhfMYa0eqZ0+HAm
UHhQJRVeCbTWCcP3BeboGAkwm5RKNTEiN92c3TslcJArj97aNpvj/FMr4hBnBLU/
qFt8+PVArnoev4RlKX9oJVqMf1Q5sDapw3YLxr2PoIgBTZ8bwjJJwDttbf/ceCde
pRX1AW3vG0cXQMo3MwCWZyaPK0lKM4mz9QAadzHE+zRo1H746mBpC2WbZeWJ33v6
IUZYmmsLr4/WqgAI911PEdszTC6cwQ4y6iSzGQj+o6fZdAWWY0Mu3biUUNKHYAxo
OMVRyCiUyRqLx/oPLUVKNA==
`protect END_PROTECTED
