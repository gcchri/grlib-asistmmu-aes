`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TpdtwOTAkcnGufQJBurTA4ZN9qaG/+IdLzGMDswicO/YX6xKd+aKRIxGfrzeuXeY
lggdqKwoGzn5Z5lmzKk5jx3jVY+bi5hWS/D+tx85dIlF8/scNGhdH9zG9hKXeCFV
9pM0JT1NqXSvHV4CP1sJs/td7mqAZkarCA4Q1+LepS6GMf/LH64yrc1L1hP3XzNC
kz79hlJbGXF4Fln1d8Y2BjB8UF/CUOeFjdrwVN4xbXbm3hdTZpwxPmyKWHKWqmIr
JkF89fQLXeYQb4o+NTefPVf+BXzQaLJqvh0qSms4V5gNRbaZ8tm5EhTd2KPghhDo
h+ZQwLl7NBrR9fG+uKPyJZjE+SRTkO+BcTDNEtEnuwuAs6iPsDKNlshmq7JBYElg
pw5aLhOATkeAeukOYevKM6h5Df1uL5RqX/W5OcaxD1MnpdtqahxpSr5RGz5rsuiB
+rv1eL1QUgrIhQtkToKYRvopS38xOvhe2/iFf/c/I4Wma/YDuVPiuSZhZgBvVW2u
64BSlVkKidGA2RBGXDhY+J6WCtPKFE9JdQjNYHO9rybI/7aoN7tffiD9v69Xqiu6
7fWOihAPsPFrgIIddDQGsQ==
`protect END_PROTECTED
