`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6nELItGSyo43O7V5pJzVbTKLW0f1SWBafr5hsOoQb5EApqTtoHilpixYT46vjVzi
xxqVIAMTW+NfMgxb1IhAG+3tjA3KQsvJCvHy2HkZBM9NgonNgTiqugQxIbaVSmn6
/cCJ9KLnYE1qSkuVTQ7p4wg/ns+v9nIMC1Yrdpfe3A4FKx4h6dBag2ejhyfHyM8r
TkJyoOZ+PY2TvxRhcPS1ObJLeYJUjkm/nfWT97KjPWXYDrNbUCo3S0TBpALDDqOR
vqtwbQ7QSoB4JR3KpauVBXli9Rq4QD9g70xDKXHVq5H4ScSG6P2wzRCHfcgraJv5
AiFVcFiT/vBl9qWDBMfQ0DSdwgPm2XHDqK/bVDEf3rFs+Y4tEA/494fbTrlio+P0
ZtXCcV3BNp1qHruSDdcHD6Zg5SZiY0bH+W56JqrbWRaMwOZ4tZ0gJeC/3kJdbiqw
byxc/UhWEq9s5freU63MZ1lHueOKoa9LT0Kl8pGjzfG5LaGMBJdJRg/jKO6mUM2i
stk+uTnDKHG3mb6iW8qVqVe6ydr7+kO7xnXe+d2zcqOPsuGhBExK4A8swmgsX6vI
FLClRul0OuKwdUVTPmbwcf+PIPkAglMzULfvjJWWOehpEarvg4LTBo/j7nlVe8D+
L+6kemoaMo4LAHt+x2qMy/9RtG40UYQGjnc09dmkRQwxBWltOh5SCTjqkpfbYH0I
4zJv3yZ3lmuN+M/fzhmgigBCZUlIMAhER22bZthAIHeB3e6hlx4hevsSjR0whiIT
OTmWg5zmsYUtDTv2CCZnsTKvroCwnExqtAoNKbdfiVjMdj6XP1QdflwS2zbBmy3U
z4zEN+FggGYBfXc7gdlDkMVXtqw0IDrcIA6SQ47mUSzu6kcbz6r/Ny3gLHREXwDQ
RdH+EveCloy/kegT0vwadsn6WepY3rI3hCAMfL8rh7yCh5aaSbOw/bd1FnDrvHg0
Re4ISM7un6qZI+qCknQM0YAdiPqJycb1u+NbVvkYFaRJcZVMBk7/eTlPHXgmZGI1
ApIAZXb1g4q0kNEKmnvCkHCFh+bo8wVLcXTjjbLKNwaemKM0HpWY9B6f506aqHBK
AeMOs6y6dekUNV8zyBfUdTAiiEn/tCuzJJ05ZUa5Ql/O2BRNCyeMXEQRSJ1XiWm2
jW0/03RbQimDmodmHDgMylmi0bvQiZoYLRDcUfu5njibVMvNiW1NXqU0xw8ccFGb
08KJhg6T2TtMTCW34NuZXG2DbJYXIcVViEYs8s+NwiK1ffbOzC5GNiSclqq81bi0
`protect END_PROTECTED
