`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ue1L9E55NT9kuFS0gQUTpW0SXudqW/Eye1634a7Cu/2jDZr19mAqjBmSUUNXZmpz
owfMRWypPfRJX0jzA+vcOU+eyESMQgyFMJ/j96eN7aevgGVDfdaWkXfZKIRy7H/o
Aa6O4zg8Y+biTF8DQKtaRdTJmdm4TksSZuITtWuGkjqnCXXeEpeQe8uM2IAvdL/x
5SBhttonM3WxXYokQr3UucLhJTpKkfqrRS7GRHvEroBPTmKS7j2MWLuaNxNCK+m7
2BJ8+ZSktW6tQiUXu4nvU7Hb0EX5ISBWfn/Pav1auGytO+hPo2K/4w4xz6EFuO1K
zBks2uFOfa/Q6sXHfiVeJDhz/D12focHAWJVDQGx5lZDbFLZqBJtJO3cHBNtl9aI
vwcVl19q7gR6Q0cnYdPw8ew0qPKZ6yxPXsN0JCViFQerWA8v8g1dLKmpnfSE7cIY
d3F8znhYR65oSQSVC1V/SlD6isejETP753wvIZx4Aj53jNkXc5Rb7pl4DSqVX88Y
MvewI5LCGRirXTaeGy27IAyBqKqtrUbBkGZHi+sTjp/XwklaW4CgJA2hfAjvtU4N
L4mSm2J1iw8Yz0PcNiAZIAgZzcgf08utC/9aqVBtSyCViaF/4F3m57A7wM0sVhdM
wxO6tpqJKcPD7RM5CIcWpU5g3pt7ywGW4Zps+N+9FgVnJ19+KkeRZS9ALV91V5+6
V2wUX9UalsPm/dxuT9dULO5VraZ/LfJp8cPwUK/ETPlAumqlr74CRUh/gy8brD35
sIOSKXY4IVs3HweuqKEifGtpiYrbzt6fQuOi4FPlvj+Gt2IYDEFEtyARpAMZObzV
7r3BL3rke5vcD5rPJjXM2PNgpCiophzQ1b5sxAmHnmYi0aEpyERMQME7ZR+NSiv+
4E8t2f3isM9lAYcRnwlPImDZ4Q93rNrVnSPI6uFso4mae/ZRGr1myDG+JqhO/dJ2
GvFOAvj+QzS5iKKZMlrakdffK5vEgrd1eMgIDPxfizpJLxlcdJiKrcos/5Atu+34
/IsovK3Tr/qSQ4eBGpCYhW4oXNgrGtnAmq0bdIIH0yAKA8ImMyXX0BRLQVJzn4LU
04jc82EU2xJ3+fgY1bVG7YluyhcC8JvH9y9Ca1aT1eTihcbIVA/uO6G2kPB7HJ/G
ZAOTTF4rwl7mpzbY6DwU2pc1P+epM5dwXtPwKHoofxLE6HjTRNMm1wQh+qxs4Ij/
z8ETfMYhrIqhb35Afi8uRC4VAyUCkFTH9NX0gsjI7UNsOFZNbjbU0Ll27zezWcny
XDAFUAk3sQnk3H8qAzsgA05lZpNNjes6DEbqIN+YTbtVDzNt4+yXvLIjfGtB84TG
62ZYMr4Ist9ipkq/5JEBKVbbxKMBOl0oE2tWBvQsvKh76tG+VbSLnB9uq53tw5Jt
NEfznNqxYvk+rMNwrHlvL8nBACxHwnAlv7T0BA1dhs+DbaucbsjTCUYTXzeW8J+0
8R6apC279BWgw0+1JnWvCsFJx1S7AnLFj5j61zg1KK2ZAPp+eXGxlOLrIiAgjfiH
Hcwhh3usBGYkWQsEIK3X6+CKWJIktPd1qBqw4Zaag6/ZI5yFb0rIMsS4R0ZZlmb7
jPj3mCk/fhu+K3OTQo45eN+riwYIjCl9MydyBWjK7i3GfGtDPE9240D20DRGdwZd
sB41u8KElSfLkhANEoGxuXBJLPTNJ3z4yXeMYatvDwy4wxDr8znmRGV2ztnv+VnM
1lOBT3GzYPvtKtknhD/VTEziEjTdvJBBpe9TtUK77sF3cYeG/1kBgZrGtDrZ4jdv
dgLNtXGr0D7gFIPEjSNPM9y/dOOHTXN/lp6svaf+kMwbpleaiTWg83UJXOjD9sLE
6GJrRz7BuMTjoqAvLZFXi8JzOMbwrNFcsvW4XnLim/brxIwUsEiwIX8JeE+dGCUK
K57GoJHDVfiFoqiHTQgAFe+IynfUKG9eFoXGXUSfOu+IY3xdy52xPKgf86VJcL9V
75X8CD25WqUmI3flVKyj+C6pYZBnAo406+okqng01fEBDebYTTslKVUXXynB5QV4
2Bb4UE8ZpwexgiOuMXHMMc2ZVK90Uvez6cvmghb0yzeHzQjT3Ik5YpFD02VorkRG
FxBt5gAk5gHdBrqhdVIZFAOh1L3d8Ol2c7h5yKpEA1zywP95NfUibNH1WLaPNaKY
aC5iNyUrltu7vLTAg6I9QyLT6Jwa7fs2esWnfcpvUI7CoEvD8CpH6KBTIqgPIK4H
m2LBgmY8TpEs4s/X8ITqrE4WF/ucfNZZrBB1vTyq8YJwwUl/P+itl3TvhePo+K6l
4GT94TejG9LweSRgKpKv7Irys1aFtpfUQkPG68009mhTervy6QpsIABwdZay+517
w0ECE0GmVMR2P6PH3Eve5oqkMoYpSJxMf/Rydx0sroKz4jT7nRuyAAmLmhi8Tn/+
FE4gh8phUYm7orXsWNAj7dFGiSyyS4Fz1cJvsHaToCCUBKH8PvlA1UU2N2fP//hB
ZrV4iW2usQTkf92Qh6kfYc7bUpupbeg9hKlJug+DEg9uWFD7faO1Okkvi/wyt7z4
qOU1cElpk/kG+hXrHZQLCyjDr1xem5htfSL7PtHFFr28tRG6CkmSuDmD35pVKtGi
fg2ovc9KTS71ggTwqO4Un0Nox7MFGKyts3euqP7/db0MrqpLh1ma0SV6xHXMYqtT
Q21FBRJqD7zPQoNrtODtMZTYdIhYVsFpaN9p1CQkYwiD8uPjAzKzTBSzXHaDuFnE
gDihL/PKqQwXvsAnC4FubFav4+4e/C7hDR0sEtdw6MAdJgVFbV1Q8d1BGdWzJ1Jd
s5xdalRG4thJ/yW+E9RcKySq5mRW5J5jwbpZ0ve/xS8nfB06HeAo5vmnw6GKCF6o
rVjByjITGAOKwZza79iPE4skUJfnBrE599LRoI5Gv5D5V0XRcO3ZnzgH6ZFs2txo
3TZVm7lNB9L5kWd2RpAkFtWeZIXo6AfTqpBiPxxb0PeQT5ZLwZQA8djgrOve/9I7
KgJ723Nn5tIsMcbf1bueFkGtb9oAaawTKVlRIORPTpeCOgGEJ8/J0bqr3+5dxAeC
XeHGvcRbI0rmJ7i7gNqyhcyKprFbJ36CgYbtX2rP/8Tr2quDN4WdRz898712holh
ZaoEc1He4WrW9VqQ7SpBEA6Miu5VppqQBe4S52e/57R92C0YpO4jrR75Hqj/0AiF
uvBfUPweX6TALOsYaI2gwS3WTyDrLoM9wvMqRZ6W+7d31U+hLaaBDQJyr5ImZwZB
qK2iTi8sji2DHrLNZgIDuruq0HhfxNQW7asA0R9XSJhGgvvCLk9Dz+DCaQxPi9bq
WTAMeqpBRgBuUF3+b03rpfBeMzl9C/6mGqYQZBkF5b10WTSNW80+BJhyLkc4jiTF
Q3944+28634J1dQYuyXvUxUuapTQBiBqM7kiYdDQaKIQUPm16jMHkwZIp2Jt81Gk
toIv9ZAKvf02rIZuEJUUnf1QObT2Z8blu/SmKsQA4TFD7k0kgnh1oQd7ucWAcBDU
ROr2/ObtOlSULyuQvMI3MH8zVhlqERbSYKPUMtjMxbCdQBpkqBLog9M4bT24AuQ3
NpjL9dTn/Io3gdHJqezpFc2txUoIX3kZpt82ruHLSXUqqU1AaRI0FBoXW5kmy8Sn
X4fxup/ZW6jx1LbtU1ZUwfEGIyKQ2unvLM70bqi1/N9OXjdx2ASQ1KzEXRSfWXyq
4SRPuY5pBWjbwtz3kMJaotnbUUbPxvo+0v43oe7qXCMiaYddcjpnzPxJlAI9DrzQ
C1vZpI9r7Yk9tMQgTc7jdlZLfr5RBMEDX8XRtt8bWGd0nfxtrVAo/jFCz4ReefoV
xruto811GgEBckjQ59OtGF2rKadTke+VWKidkn752CxEtko+/0w3YmzAiO1ayMQ+
d9EYBEbNwFxKCzRYhNvxPP2o2dnK7HTBE+wO9ceRJ/n2Hkg7Dsamb8NeOPjaZrhk
aKRejGm8faeFRsex+4U5/H1ST/HAnxmSHnnyp6I60fNvRtfwKrP/Xjdsykkr2EG9
dHdUYOWyOgJhpTdnIxurgbtr9A3ujvCebnjBfGE8kC2D5vLPfG/AZTN32WE6zvj6
T+ZgqfSk+bM2J0yKwNSWMb9mHEvMWcJ7+xvXJxiw+zSB3l83OGjCpWaOJ1dDpGUz
ZW+tf/ogTLj3nSbM/8jVMFGmE/lQr5gOMBxCvK4dNSfUbNAucd7I3AT4m/3VdA2r
jwbHU0mOaoABuCZ/EfOWzwrOUojjsz220bPB2T5D9dNA8OAtjtnY5Zqr6KNVm+Cc
PwCPxnblyDY7JlXZIxwu7lfDWSLcmhwp2xA3ptSOUR7oiqQJE/p3H4RoU430QHd/
Gbs2atW17Es8OvDDWx44IgCHSY19GQoLjuuvLgAi+5EsHxFAUBOyZLPD4dhxfiuc
RCxmV/FtoNijY+UaDWYns6dYqtFYHFPtNBtloQUScCd18N/yTT2GC3CYdskuEX7e
FVxxChGTtcYQeCl5WfYPovPFND45xcjr/P/PMTilx9CLP7GYhOJ+u+pUR/v1/nh4
Pd6qxE8WYDR3ZFBIooscA+A42BJXuyeaCTI/Dd1azkAITA1We+lL/6nVlGSF2FXc
HhJl5K7TSFBIFg45ecVqA2Aju+l/LgvApiYQimXe9aeTTHKMCfU1QTc5JCMamx/y
oTMrCBTl7UC2tHyYjDvJ9nOxLdMPaqyiuvZsE+6Yf1dvsC5RlI/kPImOGNtCHZoE
DVK2eoTElP3vQYLevPoIOcg1gmqi6rv2rzQSI3RFUkwybcE7mt8fz1I8FWHZoD33
L3rqtvPYRhiLDY8GWAh1AbJF7Lo+/DREDHG135mLtDvZaU0Zf8QScX8uFBaNleNx
0KINxOnuKgBY7OPLV/kTFmRRyH1pQO/U3e8VsDfXyvTHhZLKyVSgc8nl0o2/HOJz
116R7NPuAW9KDmpUzoA8DAQ4CxG5bnhnmspvTlqklbKant3qpKWrkEGldEbmv2Ul
DNDN1nPNyYtK7l3/wTnX25R+TgZkrEtDb3F9h+QjWl0ERnV76uYbPs2GEujD9fSu
ET2YL/G732UEToHpuy/IZWq44QG2diIdK+nas6RoNVGjmBvvecYU2fJ7lewTcqQT
Ia3IX1nsb2Ih9dcmBsMmgN7DMVGA+lcrsK7yAKw/yOgfbE68E5RCZoAkKaKB2yb5
uqWBgWznfAWz9yD4UD0WgdZVBdaApFxnAm9GfxJQ7N1+q1fbZY6fvN+U8rJdoXEA
v8CGWBos1o561RhDpkAX72STSqpNmb84QIQKc2EC5KHnzDVILWfBvUfUcE5AcN1V
80zPzCp6736+/PHkqVkjP/6WN4DAqsw7vAwAUuR+IV28ZLxz4F9xvfvxzzbineM7
lOVV/ZihlkfF0I39Xqekuu+UtSvGKk7vcx4HOzCyt1MfjUIegzRXE9sapViaW+/W
TDSPWKoYcJG1ODcNtmH4o5VsJ/HMUIKEteIMPM7sRzGYGA1wK5St8JjPfwwgbGfR
wWl559JePAyVopv4YUC1mHCWnMyZ5mN26PC7JiAihVoaWO63kCVkAFqz8ZSTyrbR
K7rMjFBX6LwilrT8OrK+MVvHNszoJVziS/qIt3Rw9V0rAdm6ej/z2HC0t7Ze1rGJ
xCuL08VFDJ2qxh7Go8jMvbaxtidVv0VwzoO0/9jg9mJTyxAa1M7fpJJXvFAWR3ig
5I/uvSWUvTb2yygX81D3dWOM2nLuSUvmrYLZ6cSE9xhLZ/19m0Bwk2/X/48ZEGXu
Mv/UPhx1y3TZuExtIceY1i26i9ciEnTmhWoDPsJNItI4rmvTbMCOmeL1UbxTFtSC
yLLEIWPqyGlDRrAHg1NkC5rjdlqYBPNykb+B3PevJpURRAzwROPO8z1oOcvcI0vj
GbZLZu6ik5OoLm+frGUpNuTto4P6beiBHpB0kVFReDABFWpj/wL4/9O30d2w/jxV
gz6ZEAaMZc6sTr7rzvmBRcGTFynmGl+gaeL58fupx8vaiVafZTV325A1QbV8Dd4B
52saaWJSamUJlFFDMBxouhDl8bNMJc9bcgHfrYk0m1ftzpxQLAacH0NyzIRG7WKz
IXB7oLLVjHrbxVVkyqVXB6SzN4p7i2UWx/v1mmd4BOS/M68PEj4q03zgsiUw3wH1
zAXWEBu0PMk7JDftt6M/0yJYuw4D9lhPYHspG1ENpTkWMxCvFRevmR+80L/WzPFG
+gsGUuRcLVlVVo+zKNQhsiXmfKUD/NN1lvl/iEgoRRjvixQ/Aa5LkWayqEnv1v73
uDJ+6IPpSkvfcEK1jI1XSnfXryYQwO3kbguWDx25lpdX+4z5WYTzM3LjuqXBiEBl
Y4wdqHLKRNGOo91FheXVEi+h61kwZOAA2OCMa/MPDLxxSENDm0HOok49HE5fmJha
DIVEaOzvcf+TcXrZW2fQ4+Y55fFFI6m4Zz/EvJlkYaFblGGbiMH+5F7guRThwGRg
XPQ0k+Um6EsvJd6mSWRtuDHkHH7987GdtLlsjau3HggQc3xwci4F6ZMfV/kTATRP
jQi9/ffumAZmYCNgpiN6bGyVwY2rpvr+pLceyqnLl/D1QJ6iwoVjqOGNB9iK1hvt
h9qAqR2ArXusbqFoAJOjVso955a+foBJc+IxV4V+hkmpcVuGkAp8qDkjvy6YmHYf
5wmJIA9UcwxJYuMQSbsO3ceS9/3S/t7bk7cG7aswkNRRTx5QXkXtFl1lziuUAKon
dMAIP1hWZ3W9Em32O/nJSVJxXwEdBHax3VZoiysToRsPyuG08iG6MUOBokW8BavK
YBF8w8/uPM5VKhpq+TOdvKB7mEi66H+9AzE6fLiXlAehmpAp02mqiBYgCyYZ2/Or
2xZycuDscfZgW2LdMgc2GBQMiBI6zmj5RFpyN4yX6/N7iSOB4petvVpGq+AaK/lw
8k8VEWPETu09d4aeEzWmNrZbmvRQrDRCpsR3lZ8BLZBSQ4SMYnQobenq+cQOprm6
70YuCcXYA5Kw93j0FKTqGMXc38J/Qv0ATPNqzOoTFE+9g4KOaghugOYLfl0n3va2
rGZGNUdAedSw8s95FtzSffJ18hbKNyQcu3hnYXrGkq8SiD2gUwWvzB7zldhhuBVP
nNN+ZfB0L8d1wimU+PVyMQOgHmG15/7laCfI0RB2RBeLrgBMZEFIlxJr2a1nTe3P
j31A5pQvXyJwVmfbNF8BrMjEGNO8LDtfGdz3o9wZwcsBGjb+rzWo5GjMvjJiIMcb
kJDlbjfQtlcoibxRByavgLvqbrcn7SMck1onGS3upn8QsjvGspNkiKT4+LE6uLi+
6IM5qVyaHJMF9ALBFLI+Bg1eDGmaIqGc223osERxVnKonU9ziychJ3E7611H/RBB
wnWMDe4TDloIzSqUwbMEkNZ3zVX98eqsw0Sl7jQkV6hieqOkPsgcGKISeaOeQf7d
cfL15EafBk/hQjjOtNA9JRH3iQj9YeGeGX8/7QxHRJgbPjKK8FB6Y5sFSOEXgZiB
cBwKpvKt4smt406/qTMvbhxHm3VREGbfITjj53BbfHIUKysSlkYLsGTny1a4Jskg
sQObqpoksTg3xEkeFucZ5G5innAZaG1q0UxO4zRgAKrkU0XbtiRS2Jc/AiZjs5dK
lSEZlOo/GFJ/l7lmalatKjYYok1TIEq4QIT4OzD6S4ASOC7CUMn6bxzL2dd7ZDvX
yVMzlA9xIZfxsy0x2gamPEJHcXGAWBDSHKx7JQ45MWudI1p17z992z2NbHMD4fHY
K0pxGn82uOeFz6LfAm+fCW+svD+GBnmVEwiKNxQgywXPMZkA180iCdFPRQOIeU5v
o+3WkGhoCmHfLajg4Km9vLSEpPt9bfwnLQgjqV5puATAKuRBtaGAFWkhPf6w/pmq
wa1K/LJp9eSFEcuX7laEq8vT+Ie1U4GUZCfL99F7ZILT2QteDtElvDuXsm9YZ1K1
xK5RvB545tfM9YkFTacCdTm2syPIz3NZfVPQX9AQBfH5++ICZjw4NKeXPcsiLbIr
mup5q5sTq4RfccWhyNpcP/0M/fs+1Q3FidzCcGd3AZbDyuiitQw4YWtYIBX6vLYr
eya+ptmPkoFsMLHQhuRLCkP9iy1H6H4BM+8Cm61rQdGi0CisGXSl6JVgZbAluSwE
shlEjZ6oM5cU7z4cysnwMSS7wHEE9mbrbDmszRsxsOh2rk4I69SDAvpX+XjburtC
8JLzMXRZiQ17fO5NVxJOM35uIgo9NBEYsIMrw+ZulwYWPOpeBh2kCK4aKfdnvriY
Hcyo3ANSDb3MDYEqxwNQT2R/0DceFtWJvqiid/aCiKTaBk1lclb/L9Yj9kW+cvwx
Sg7r811u5hYi21FhqGwQhnPis/JP005m/36SEDUIO/0Djnz4qg64u4Fu+UkJbiUX
lBggCX3SL4RrSktObz0KXsPxJHgLz8aPOfW3Cp1FOJfIDEmVWUtfbGMWHTyvowib
nO32F7eCwAsl3rUMUH7k3ord85lx/0BWmVC9Z7iiK2VE4EbZVhhp3QuJSSMHisoI
mDC726s6bZbCboGE22D7qMa6OMeNWA+S9Y+aP31MSryqtk5wG6Z6+vfuSBlWm7q/
4TzAJaBMH7nNdd7xpuLYXRvrOtxMGjl1HKj7A9Oo5MD7lIxKu/erfjGZRxLQj3Fh
gJA1atKq0b8VHJbDKj7GBoMMaEkiN+GXKFc/pvbAcc1LE1Hust3wfnZLNyYd0HKw
dzlp8xCJmCkJD7sa0kU8uxsL3Ts0/1cd/6halisf+lIs3/kiD15zggrwl2aXN4ia
l3piiY2kPnM284yfjh3rsjJGIhSjxcwo7gRk+TMwTq92vd656fnl51MjuNhmxegQ
PsFGVhfEWXy1ndBg8LM/nG4/CjIEoIQk70Y+9nfPo3m7IxKwbOvKT5maxlfazCfz
TLiVPBKH7ABOcQU9jOTYpv2j5AF/Gx/Pnz6RS7XjQYxsgtprD9pwiubrykbzDC12
ebM1614+dHcIo3a844++O+7NJUtrLn8/RaCRLEUlNmYba1ug3veQFn7vSaU+ckR3
OwuYUJFBZZVySBxgQwLc6B+Hl+BlRlr5eDqBtSH5doCrIdk8eMei3Zdykx02i62r
u4QGYCtJOxzArmIh33S+iakYI8deE3jEbIa7oC+tlucfd3N9CGABGgNi87rBexWg
k+nn4hD9N0KlOL4DVmYJeiSt4f32cBNekf41N87Ruv8jkG8XGOoj+8IWiK33qYiS
QRwyF/jB0gSSi5pcG/4Wfjt8lEMnKxVbDx9xADSfWn4p4oo0ZeqMJ+HW4TP8WLji
vfOO8cudK+wU3B8JftkX9n9uWCenbUsf8AR4tpwVwirGaVV44jjJz7TfxHk5MUL7
NaMSo/3rvsUTQioQxLXmOuKLlA5sDkNvVDlMpsCz/sX2N3SDDrgjwphmrwvO+eHs
qE9TW86Lgz5SbTXsLxEQu+43AvNRxX+2b914oX4pQVbwPsQWfRqdf6iatuuwKf9l
7ug7k13Jcmsu5PaSTqRi5PTJ0cQvwNMcIDoxxErwCshf7eFGfzqE+EqpDPpdFs8m
2JQyDFwoIQXkaUzIQ2F1i5V3q17rI3hkJT1SV9udx7cFTFuztsC6psbtfWnI/hV+
nPHLnYti7Wf1e5MvPOlBkyJemUathuYkT7b44JOdSnev3ZwptKuZGXl7349rRMRo
Wm0JeOFPFoMKkumLQ0q8sgLLrwxWovzIJ9E1PRpWwPqV0supFDD8I/hQpKI92WVM
FpcONngatvvB/PLRNw3/bg/s0doyjppLHM9e9mO4Dhd0p4b47UxMqf7ZYEcmTSc8
MVpN3gnynQIu5nl/JWAk/YUD6TeNxKsqr4Z+5OEwzomX57RMItZQq5pZykufMR9J
oErPcN94O+2DQ2fcyqGotlBz9LY0pZ8bygdSBRfikoZtZvI85PPGADCEZSw25Iwp
oZsQ4x3pccloiIGIAL1FAHYrDnevE7zFsaE3P4x1ri1h7h9zuj1zBnz7yqR+WDHN
qHVrAz+b5sLOPGJNyM6V7cN0eR8rRsjsPTK19I+oMYV9eQznEhTgcLqoHBM2IIHM
y+9FDB2GQIJIjQUXC0dWDNJeB+VAdNgjnKRfHJdHXgtAGBtI4iczUhY07qVRQif8
t6zWI06pdlgyJC0jtdU0JeoZkSdkFg+9xaVsSonJGsh3m1Ym80IYlgKGxyzfX46C
cZO5jcPvlSOdEsQ2FGO81t1g2OJ3NUKTMkLEsVh225BOuQd+kJxX/prHeEE/AeDM
1AVIrEu0Mc4kTrFwBdUyWXkoW+pTeBzrVuDRwqXHMpGRRLYiKRFvmy+GL2hD4eoY
2j9IENXl8FYzTzaUeXh+sqPU2m22sma0/TCZEUMuB7NBewUWx77q7b0mXpktb5bI
b5DPPTLXp2/uhWIl86xKxlPMcEshEdCVyFBF/McYMdZE7avuNYYJV2xV+njhkk08
9kacYmy+Jki0FfRcLP+mIgZiuT/iEbGFAlvBiQAgvyYSFH0682ECP2f5iGd6wgKn
v4B5x71L5F7sng4XoRdxamH9QSP/u5+0piYuND+perICTKaeTj2YZVI12g7QL7vp
gNtxfdVOSSZzxCHGXIE+lQqARPE5P+Gw5bANzEgSNMiiQTIKnrVtPcJX8QucpxeS
Ov4S6Shacjxg6r4r0oCjElrR8Wbnjpl81ML14j2jAbZkQ59ShMqTCImZNOr7mopm
ZrwwuoGlgZNsuKP/CV1f5iU0FkSsAqXDlFfTgvNBpQd8R+fgmB6osNA+hXjZPKd3
g8wvWPrv7j0anoEb8pyJxrHfUCTqI9ju5X8CQsbN2NCoIa894svbEaXH0PpJKimn
G8nf5bsb5LqnVCeLNHvWDOdhVANvA8fkDKK+qf0+6DAJ53LMmFKUZjVJtzaFwwzs
ZIHIMVCpbnkNc5DzpJ1/wdEEQPsKBmcOHFtRw9GojpADq/Rbk/N9OLNCwgUBJ/Yx
F9wOfPdKxkHsmFPXqWAJPI7b3y8oBoROUOAP0NEYdklckneePywYjVuU7gWDDphh
N+MezCM1bWmV+MhyWUZVmKVulp2iSbElyjTGKQvDGlyBIAV6O90D5dNCo914ywXT
gk51OzBfrcfj5mJHnE3F6Yp+Yvl2wNQgVg8LDKt7OQYxbNmNo7dKoX45E0Ik/89B
5JtQkQTaYR6fD87N5s2O2ru8YcC1KCM96KG2dpnfIxpTxpAOXqbBmV6vJpW7gT7x
dq8Mkcp1PpbXPD+mWLoMn1HHoDg//mZFKbeSZv24JstfcdmJxOk8tbke5CCRxB8M
7CZp+yhuwbvO1QfIx0Cn56B1wMgeu3Iw9PA06Ni3P+BPmaTBZQl7fePmYOfHNpRP
GYskmjOFAgaUnYjEegXIF/fcpgGus0z4/bVFwjGOLyYv26Dm7xWyVM+zsZD6WeGG
1eZzvd8/6u1vZ7UMWPBiuKyIZ3mpjKATOXYNYyeEV6UvdTknBuHm8AuTSutOOKkw
BccPydblJb5ZTIBAUuxs9eIjAx6o0bZwe2Sc8jjxIODYgBXQn5zmlYJT11/UM5Bq
Q/+k97NbrToks9mok4zwGWafAYmKGkEx36VbA/Jdlqi/pR5LXz15O5ltq5bpMSNV
ma5emFKXsGWCq5NZK2VwuzS6dlmy2HIZEu/OvVZAmyKiz31nS7B7ce1JMuh34cHn
oPdifkYhkr0mInu2O+vQDzRwpvZAxxvoVM2GF8JyGqAaCo9pQpx3AS6bWa44/0BX
1zCvJgr6O+1IbjNyqu1wxMEabr81ENikTnwndsdkAVDRjlrVGcpoyv1g17c3927l
QBLjNL6TTjK3YpFXB3gImk8QH0irt+j5iJHnXJxp6QcnFCHYOFYZ0rXvA9SsYna8
+vs/h8+/Zoa4JGK2vwlo4jCv8M4XrHwgh/AculJZELgY4aEmZA6AMr3Qa57ZhdbR
hqd7MCTfd7XqkV0p5pZCgJccJ95WGKRUSKL5MJa0w2s1XJwTOlBBrlzsEqLv/0yC
TryHEIIfW1RVNVCRCQMdcxF9VZwrjDh1zXkfOj0Up83qqsxFG2EUgzQTy9QDxOvD
EcilMDxHGyrpE3B4N0d0N83axzU29hQezYjqTdOItZrgBj0IpH7ZjH/qmiH1zvqZ
L2RB1uaqaCpcTHaAOOCUn3YFUyPTgM2Q05+UkWUacevUra2DgCa7ktEtK5IQZOco
ZxEQOhBtny9hEJXCkb2QW1+6D05MclBnIvbTbS0xhUZhqLB9If8SKI/KoCImDmaJ
fTu2/Cz3aCcf2UKeW+ndAcPo8N5H2C7PtzwEJGyhOyVfoRLk+22sVtHuBfVafHh2
bwH+H1WphLfOmY+guL6Z2JRAh3SRzC0AyLEwLfhkMJSGbKbya2vPLQYmL8LpoUpE
MXWlLnK+pW8Z0H3SdN2eqWvS6BOUboyifxsJyhHDaKglwNZfKrQHXvQ0F0G5LQGM
gou41EJK/plYGUCcBSVUpYuypkDoVGgeX1RlOzcOdo6SchjCThzDfZZ61Ou/EAdt
NTIcbVmQVNOBq6f9rgaBXAKhnnu4bE/iMpTXZ+rv4ZaDPQxL0Fqe0+OXZc5kHrkk
0iFBsinqrxl1X/P5umUq0r0fa4pQZNRDkIaBxY9VHAWoqGPhanGwOScFu+mdXPHV
3BwPyymvmY0D3AoxqOqlcKClCFchYCy7/isPcscm4u3eGUtLLLCcSWWPZm0Jj6iX
kvSdYeCZRBusqP/BW50JBEdROlT56WXny/AWVZNz4D9vLtdtzlC4S43EW8ZsUlH6
xo57drnxs6L//ZeKAEaa8PZMNeDs+1aeLZucDEbGqS+G90ah+4suh4PM5LaDpN5S
4ZKLn70ZLbjysyJcVRXM04AiJ698U/VaxhC80NetFsEluIOKuICWWyUnwGUFoxho
0QDaowTC3KMb2F13Ml7exvn2OXNfWKmovfrPABaek3AuF0PFtJ38S995gjHWmQsl
8k9nTJhlkhizjhvEPKmmPBLnl8iOSxBcVXOY2iquJk63W0M+e9Gw4M60A9+W1j5P
meisbnwOYmqyDVieO1RBRB6H4v7pdhFKos+b6/Wdwvndkto/Vsj5XWjjSXgO2WqR
bPEw1HWJNb331ZlPC8G/70/XUfedHAfdPNlx/6Z/YCb+J3a0cLoS3FHSozzUx+gI
gM0bgygSWFbB4jH3O6UoXJZYVApyeIWN0DGavEzGo7UeoEcOUA53B3U/cqNpM3R0
NmKj3PLhyt6Uf3kK857WFP8EQfLkVyKtygf6GhUWyXnYUH2YEIyKjPRl/SxFAJrg
i2zMAYWTHnd9PfBnnJsF5bRC+1jnXh24oOT9o0oC8FiBUZTVRstbXulADF9yqjnb
5IVoiQsF+ABToITugzg5TEAQJXKGS+Jir6Xc5arwSz6hdWfN8RTTz6EUDZW1fNlC
Zeg94wJ0nbfAhIlRF+aKB98+Jy1VTWOT/x/Hqx3lkRpgGgZgMKjt+Itgw/DiF3Zp
HJj6lgb5hLGQyjZWBfW1BXmOI4wuK+9LwolXQQ6wRG/IpCZxlRyMM71C+W6BMqbr
xK+nWmCHrBkNOqC9eeu2pvKGb4bibjNnN3YwV0FBXBVNS+1wnv+/SgHTWnqLLk44
GqDSF7UKUlwvGZ9xhQnDV9zOyrVJmtqQoUk5bppqAGNiuI+KSaJ/7oXKqWcfdgAb
7W297ZwSOLVYY1HZPGEh1nA5AeQxbkHnRNCl2HRxEMjKea2Ta93ESf+GPTpByYWX
2uv+rAVRMSDokXoHU8e2OtdsXOD5ENTlFYfUahfHzW3UvS/GdUth9h1Z3iOC1FJF
XsxOLfzlb70ghIfNE3XrR4TBNytHrdanIqaaEC5xZTieDfqnEZiHghx4bYI/j5LB
UMiCZH3n/ScgFRBxY47O3g2UgdRohME4S35wlRs1iP7gYeoIKiD0BseiGje317e0
cen7mFFJWg61LQHy/oe7qIYhlotw/HVUX9rWOXk9prCD54JPeJodFJQOQp6VKyGb
L3WBDuo1U0VFpyFvU8VbM0Js/XRQVEl4XbuHDCqyI/Bcgw9siUiHdd/xLIWN1ek6
puY4gm9oJWFqKZBxU5Fk1matcZEZaY5uNma3MyxLfHgLNr4pqlsyI1H8i0Xyt8Bl
K/olMFjDpeWFBsGqLgvh9m3miNIiFEb5zVutPLL9HiqYCalqd7MjypRL7eVFawUo
cOOy58xKVAQBI5tZN4IFhXbBWp0uBMfEdeuGEvrsVdFq5A1/KL9gagurBXxQ6nXk
/1N0ie2+aG1cXpecCk5SbpmHBlgRqgm979KHDHRlTkb7s+xlAi+G7b0796smeJv8
Ag8xb2vFZsslzYIF7EVJXHO7nTY+fcObUAzpK8hpgn/npuf94R+zjIgBHepybBsD
n5EWN7o5s2Wu582FT8EyXrM0NSUHaQ61UonQQoberahWLvj9tmGESKAOLwLy+iMh
LEEmcc14r4J1YrSFCYXutcouRgOScPVxkVXv1nh9wzzXOGojBjW2dHCVx7K3bVDU
EP++oQqtwYxww1Zen2td2n6R1rFdZYULvdILSxHNeys4F0tO1S3kvSKDhRfDpmvw
usDV0UHv55urX1gMbHxRgt+j0g3yphGncMcROEbgsk315Y+2ZACEqanEKU2oH2S3
lRc0UO+BcEoIEfnHVfAvguQI08Dbk/iYemxjycayW7UmgfGWIzZ6A/kl3CL2nXM8
iisgYscoFNlvwubLU+E6+gg51A9tIfUuJc0u48/lQOZ1zS9ZXTJyNoFcx8vOERQM
DjkPcqC+4q3P8ei63uDecyW5ANdd6E9YeynA36pixU0yziIMNe/cQZQIqtT2zZS9
1rblyJcUnHPqKDmTqe8OKG4tzBhHUj0vIXdP9dLJeSmezpMCzymYvHS3QnOA10+w
WzqspNkh3q9aY98Y69yqkvxjtJ9exKfF89QUKbbEveUbr+LFgISQxDMuB5Aoezo+
wT/cBUy+Lp65kSfccgDg1URwsaCQCXp6+z4XR6NU27bwf9d+HbHoKqVkwr0aX692
XJg/9b2nto1W1AxwE3I2rcfLknNbWNeMpjhKkfEVjmLDJp3y56vTXVwLrmhDaeyh
DNLN3/MK4fCZ7K96pVWe+Qx6acZ6vOinfMnbNPBjg8/XwRbETY3bp90EiqpXIljx
pfziMkn+f2q2YkvRAaqbuE8jJYb242PSHG4WjI2d2ZvDJXMeNlSDtHCyN+dIbbtu
i0cgaz54H3++qaOl1BOBO7q5zefHuBxnhxjfIwOuXu9xMco5r4+gZE0gFOGkUw6S
9OXW4pVL+cGj3mWS6A6iZM2LDNFj3ZpeJstyXSDedxEE+m44ds8HwEy5/o/rJ9f6
0jABtQnxHX2ENMiln3124O4U7aGjg/dtuQMq18aWzJDUN2oV3Gpu84MhcRO7QsWa
+Ywde1vAlXNEnxB4xhuGFW6i9Brz70BOjC3118EcTNMj6xTlr/ScA8J4HOkSV4Id
t63pYAAsY0H6FsrrC3xRFY471lulhuEdJV+n9zE5MkawC/Tnl/Mp9iMRNFwZ74oa
4j/IqC7OqB3iLmQd5C2PptlTiWGvjSmZSjidHHDlKYWhmGbNBD6oXkni0OiFTIy5
cbQtH0jcP7TTt3QH46zqH2/aw5Yev1QztYOP6cpn8l3ze/HORV5Yo+LLg8HSvEtZ
0qX48EYICtrbw1XHwatV5GXI+wnk4BLVMNxdnTQm3kvCywjqqlB/nWjQSi4z9dd2
31LSOC7nDtBMp50Ri282XsT0eMbMZLmtsPECs0nZe+TFs7dKAWHqZ16kUWj0hq4m
FcQMioq0u5Sf6oS/qgRw4+GKqZbga4ahRiHxu+mkCoGM3d0UhOfUm+/GOm9mDzmu
LCCru1rOWbAlbn9S3Pd/qevKU4RmE+Y88mkyWwazGAxDFer29rOKV0RJTqmLnrlj
hqC2sOQLzeSYsgGksGcc0eEyNnQOwI1SL1l2giYyVqWjyFL/yBQlOLWYxStIj+KL
hlJf93Mh+FK4z8s8dyTrpdmZqrc7vkce5sDIdAZuFno9eA7ykFAedA/DPe1fa+7v
gTUCWo0PDxtQhdfMWMFCFtK4ihRRahcdFnwfQhpk0M7zYaZEqlHFMHbgkS/tNHWx
mwRRiwzwlPpGQMPqRRoQ71ICikVA4LHt2c29kftqSjwyY8bNDyOL+T0efTK4YhpS
2e+Dc8ugg/EvSoZDoch+QVeO00we3o53gBgwSypDDLS37qEeMuKoVgGKdOoEffVq
WU+OWCrLfFJsr6l8P+nCN6shP2+ZZ92xVDf7twqeQEH7yR2r115Io/zWuVWfcZsQ
qqP9eklnsXOIHC/K4gHKiHcUtS21MeNXIWtNwXrfkiI6SyoRTj05IPsc7NP/ogPY
hRUBLqVG7zrr+AlMkFItwAKX2sMp27e0gcPOo6la+L32SldY2DfqvaaphE/X3FJc
RFO8pR1o3Fz6MyOEIgHmU84eG0/rZo2PZfWIIf5GqmmP1fTvAoMaqxc11/d1dxbf
OoGilwZVGrljuzxMwZPA3aUupQP43glOHF5CIhmJ4zxv21JL7fNt5JSewpvt/+oT
DRy3qNMwWJRHQ2hAAFPGiS4DNbpgoPsRT6ob0cifEvD2uXLT+FHtWsLi5U9W/eW2
vv8CpRKTzCK/ioPMnUG8TX9fvR5pYBLvl3CmmEL79EwKKin5+k5qEiCKM/6eypUT
NIrvhYhBJO/Xiobn9xz3rwwD5VLhoq2hx0I0YFfRqxtwSazFtkvLj45t+u/BTe2O
DmX1JZyu1yWwHjrLlmXylI5Gu5qEzJ0gV6ioJ8LjKidCRhGPMwVXP4E0/VqUDnR3
S2nhzqr3g4nxfuQj7dHJjvVMI+x1Q9zjciA5P+CX3MUM6jWDm2qvF5sejH3PnWEP
IfNAjyZgwzC2KqjJVjgUB4hqBLYBzxRJIiPf+XCklih/uZeC5W/zqG7+Y4HRdAxJ
EefAKtvmcKvmVYndmbPu6uXdurHvKoBrGf9Ia1TUwvQK1Ww0L4UbKio9p7NqJ9X9
KtF043zVTR3eBTkfKerTVILso9tLpUxMCvJhUAsZafgmJcJlggnxVrNZCfW+guIZ
wkVzn8aE//RtZaY/qzmCYTJzryIzvzha/2DgmQJWBnh5VQGdZfwHZjbZzCiUflSm
sNgxfLCLTLBIRoKYiEhsx7AWCESBBiWN9+I9ckc1aOobIJ+Sohze1b3cFlP/qaHf
ZWRfCDwO9CBcEnM4T0RWqR1JL/iXYkmFMBQm6EccmtW97UxzLwpx5WFbMoaSdqWk
V7OFhL5jNWd6pRM4y2E0GM1dPbIiIfbmRohwGOHApXugO5PlM03ouPlD3F7ElEGf
b+qhm6Vs6S8NgrITGmTKiual65ySiNE7lIA+rYexfA3Ur8mZPud+Sdwm1ys3Z1/4
WrBajOZo+FLauYJbIfIN/JptTgVpoZRZNm839DK6hW63Iw2LBeTnZdgPy+WPrYcm
VmTk2pOOsHbXy8XfceTWLnUHPitN4jm0436c2fZ46Ll8Rp/JOAUiQiUYde8A9KbE
TSLlrBO6dQ2LSfODYBA34BhrCfdCEw+14n7FwhSd1KkKECxQDmmmbc8XoUvv2Bao
M2SiJY745l20goTGYKEeYzWrMedL1eYP+BSqLhWE6zQQ21A1w9mIop0RmRM3HGGh
QxPeCx3eTpwAp4MWY+p3VpcG5UN1Te7sYCUrw/DzbH5egoKy1EdAomy3g5Yv4ddS
z32oRtmVSrr6g4BSJM8ipPGq5LeiMbj051VR+bCa6edK9U8lW5EhnRXGbg+n6+B0
+M7Ee7Xk9vFSgMawc7ZLkYUNeYpO71nJP/iUgWoS2lmaiO2SjWKC5IbPfDOm/BKO
Vd+5P+nysJbE+iQ4PC924HeUxtYHc7aVKq0ju3gm2R+YOfoi5Y3lb0xwbdJwNtUL
OgtOcPomw+QDlfQu/GN/E5Psx6Pqp96SzMlfuD637CVum2RhF9ZPijwglTDAIA+5
o5oaUf/dDUOJw/9Ap959wWnywHxZ7KQARyvbwGQYUYwDHXK6gup9oFk/RqhqPMNM
f8Q092xqrMcevkXP1SUf4NEvNjgsqGMbmKZW6dEGmZFXOBQ2Kn0dpLdNGK3aC10V
3RJpBKHB7dkjak9qGJRsY1RLzYGhxdPQXSBBxP/oE/+neGf7sDUTnP5QSbJH0To3
uBqpMH4q7LAZOwl5vGB1Ek5hF7NQ5BkdeIvtBFOI0aN03uviPkkRgelBCVOR94X1
Uer726/uF7zQd0VOK75T7AmiS2TsrJHFsQ4CbWZmqPAZf64ewtoUhSxK3S99lLoF
s6nQ4o6602BFJruwUIuwW6IoVglu8DiJK6q/YM0zQI4kyF7VPn6riUt+gjriEtcH
fPalO5Rb1Uk3oL07P5CO5y5Ww0/O6ptO+n9VxoijItyoWYGcr5aFoXudUtjacAaR
H08VNGepWUOu+LSB3xD2TScee+U8zavVUYG86hgy5W6X6Kjvdd2QqR/+bycjOdzZ
WbY4fDFaRPHwEWob0HqkecRrpb4GxgQpGQTzEmtMSByRPwPx72h/+knIpsis/pDO
6lFp4ZBNS2tvDnfIusQrdGmvJjNwuInCyI7q6+kroOwjhKoWVjo2y7JlfHD2EeJd
AoA2jq1ve/jayjYo1lvfbZM+8oyStG0LOAGZUQHi5ryQelYGHQTcN4UO3ESszWjK
6SH1GowX9EgYKYrSEIpNFJHHBZ4s5wa07uaRLVdI0DaaNPwXps0/Hn1lXZn6omhM
MtKSPDxtOTX10tZqTQdgcQYKwigDTYv9Q0M/sDgFOD+b5XuVpU0CJWjEC3dM1LPV
IO5QJAwwnlbImOwzSUhmqdk1YHSGk2X0ZmB7U8682kO6yfoR2cSnzLVarcyt/cbw
3Lj9vq83GH6YgWQJDdieRx7vrVr+oUdJu6LBonZ63cat3oAh0bT1TdTWCH+tT77c
ae8cFom/V/IjmBkEdj2g82dF4Jn0KXiMjG5uOQ03IwfGE5psgCHiDFxCrhABki0a
e7THjFhEBT2nX/V47WQZQSmHftQxEVZudQ4cdG8ZWPMOvpb3TLox4vnaghAYA6li
AlEXJufLT8399z+UpJcYb8vtYfxVzajhAl//6NYUymcBUuoyzp7tc8R6nsN/m+bU
eUg8f/qgtpygWKjHJnW10fVt8P32FIMuFuBIuxIrUeq8y6RNnlFzh9gfhTjgDvEP
j010YIkWMGJwjno+pBEo+rXwa5fSV1H6G+sDhUDNSJE2p46pR3DekKFdPfDCr3Sd
xIYB62es3KtBOg3mhnObCDsB59ILsTEcIARLUbDUytN+6ZuhXA+I7lX+D8T2nrfv
5GjKW7OF3yS9AyWHNK2JqlRArJss33H3XHGp9tfrClgxvYU5goe2eEE/2PJAAGku
AIgnGYcIMqKj68FMkrSrtxdr8uzLhRIrxhAQTxeo3XpduPicQcMG+XZI0qY563tP
TWjS3QTOhtlED4Fas31BlZLQ86QFBS27RbNqPrSXjfA0CtzxefTiQ4tROUHl1sfa
um+Dz25SXK/7qURDz/kPGyBTIiBOCl8GoSP4TrEyC8OS7dqkO8av4u0X1/vi5a5G
yHlOoCBNx6E1tCUkez4KJaIbumcl6fRI7w7jlldxPtyVxY7xsWtRPk7lCWoR3uKF
BrB61D8GOqV9YmaMv4zcrAnzye44/AvP0NgZEZCjrpSxKd+yzJVqLBFC1hl3O1Ce
UEiL96jJjlamvRuwcQn+VfuEdOkCmgWiPJm3dfnbeEVfIKgMEvh2yIhrHqY1RmIZ
g2dr82TyZTW2fcuNy/aKglOTgauPQDYRXIWzXhh+c3VBlg8DTNNt8rzt+EYyfjYr
eLEAh5gx/sMDMDfFzZ4YG12lmA6Oc26DEgxLaYUKYZbwfA3Dx06wBJAEGq0rhQ/r
9RTc/ykn3QZv/afRXvBJeqpsMFz3lhpKHZ5Dm3KFJh6NLSgYLBRd5tWxYjcNOd9O
BD6ieIFZgEUiBosYQg4qZBl+ll8BT9mehpKj/EBSycmOVJqO1EpJNObo9WHYSWfG
1xlf1cIM6m6gx/bWWC7CMvq+L9INkia5Z6+9QOOL4Q1FaBnXdEiLjlDoo3ea2OGz
h1bsF8sVscDpxg3rf7kJcf9ZKj8kwXUA9TR6EPRWCg5+Ikjun0zYtOdmHPc+iJfk
5t8DprQ+tqqn9USKB+6ISDKwq/eKofpbMSCLyBinQlbQQjkuOBfBF/xrxqxVMcBt
sDoRHLY9YQnqlrWPUq2HtwNJCeKbQO0Ek9Rlv1/FcBmrWb4GImS0l5AxhHWmf9+l
JREjls0tjTiG0I8sH+9lHxsyIwytTh+Ql7OXHQO4XMr0Ch7mAg+PYUYRLr8uYcJz
EnWXkpExEBZez0kuiFod0fOj96wLDpI9bXbyXXJ/ZIpcnVj2bps+E46KR5yda1eX
f95hfGqHj+BpPfy6BGqCksJBfNrOaIQKWIJaxuil8Auw9MoY/Ioni0rJ8889x8CN
x7OWuPSX+oQ868WHxsFZosYMrtFvxurY5HJNgKSfPcQXoCGzj3dPwkxfl593ThRn
uaiCdCePwBdrgie6lNvMuALAJEiBbFNeamWIqt5O+Jb/GGFWrmZ04mi4iIRIHW5z
HI3NMXwrhAxXdiSrScfSmOrzcr4UocFg7SbSVAbp88QXSQNWlnb+9CLL6F7cYs+U
DgIm4nhnMbRzbIP4WiS33L41/78ekN/z4kGzRxZe2Av/UcezPw4CEqzjpto5MhVK
D0RKsAY8VEKbdy+rFkbPt6f4JPK9eqZy6JM7Qh0XSbCM5MJDHCjr42Y7ZLIb76Nq
h1y2GaYMGqEiCk1gC9KMP6uwIHeZD/FaayccYUEAWx7ZQoCxxcumBOdQGs1aTE5G
oht3J5vXimygTPilaoLsSqpV6D9L1ZwyQebAGhslClngbPXNyrUjeP0W/Nlghej2
9dZbggFZIcwJXGwWk8IP4ThFEHzXNaWzLa675Pq+ji5DcFqFGMtOONdQEkHx9rMz
goZhhVEAToPUMtITdqjjDRrffv0Wp3s9J/ylDIlWSZRQqOXPCZRj1zOCp1v+bul9
CXy1nMp4w+XjiDURa2qWNJ8jVTSyvAOIE57Z0WkdvVGc+qbB5kMSwv+EcVQ+QkFU
EO9azDsJtNJfEUoNCEH1NSmZ7T8StfnyPzvWfXriB1B1M+F6Dhe98guuwMKvKB2H
MCsDJaGuduyOCHWQOYhBWJss7+96mXHTE08oKh7Wds5x+HbcInTvQPVH4BuFFsJK
cqbN56C0An+CcbgtgC40LOdiQz+mLVPURAU76Owb3dfi7ww5sI891ouerUj9eZmm
wMvs3i4ZxKXt/A35DF2B3tgA7HJedyngDE6ErIVBAbfNwjDjcnqi876OYGA1Ep69
R+sH6my9V09G0czQZIhgDMKnaWae0wLmJsctTBafrkscqyeKrF3GvAdbqOM/GtXb
oBWUksAEL04F20XDViUnv2Rubz6OhE+hyKHN3vVKhs3pmv5dfKtWuRRLIbLnMkFf
kW+25ftOjw4DU9ddk7WAJsx/6yTjcTKwBkfCvBLCjeuHBr4q92RGYNDWy5zpDSgA
7atXlDqz90CIK8PjoIKDOd5Pi0QqzuQoChcYouG6Z9DKIojkZ4MoSSfMxgMe8Sck
XCvGGu/7B6la5raxA+Xt/LkFxAXZ4G81P+/4Le4gaVgrhq7I4DOtVH4xaEjXmiG3
F2xcKyJsKqR8ipUuZzjcecTpJqHzWWHz05fZi8WDt19irh78CT2uuhqfDaTUEg/p
rbFbkbon8QPW7PVYwpKGDyfG1xwOgYOrbUFnhuwrN51OgUPH0Eg8+IDvXq0nmJby
87VgoWYB/xQOp1T5ARVTFApHGtmoznJ1lKXQ6cOu4EHKa/5QNQDzypgVazPBUHPn
Izsw+blK53mRU7Z9W7vzMSVC4V+HJPz4My+L+Jw4XJPz0vY0MqwuLw5fWHo3KDWr
Olzz/2/rYMCdmaccIXYOtLDFFiMEh+0Qv7d87Gv4vfH9olqISrh6Vac0OrSZ1JaM
AhmOe4UESkQesvPXUTPo8vSoF4kJ4GW/1a75BVk0AjUD+sCZBxAtARmlqu+z6FFs
aR0OkHuzyUSrjbbM+o0nDq+1L4uZGJ9jPpCHjY4sqEuYNz+fmDDd/2UM4Wfc0Att
5pktBhEacOfBY4JrZyf8Hd9G83vhKhWo6/zcloy5a/Ym+Kb7EwjOIXUCWHksA+kz
Ft9/60yL2V4Rp88K4r3BovPl8OtO8s+qAU3e3lRXU1aa4S9WCcVMFmH2OShyf3pA
wkYbWdnWOncIHhxZcctP5nCcSrb4CyF36xUWU5SHuOOt2UGTx3CveXooJ1oQI5dP
am0SVsilvc2CQDu1HtHw93U/w2+h0g8fJEoQQps1DiCEAY6KeUAVV/00h8NxiMRy
5emzCawjC4mSWV7EYTi350DOVXD6zefyKwXpjWkXg41DKKBv71yPbxBarKqGFq0f
CZukVWpADMcnbD+hi0hcgwT6aRtebihqUsnyE2u7O6mn2DSOc4Ob0TJbABR9K3Qv
APiq5nfEDi41zHAtCoQY0n+//GSvMPEAzwqM/Z0X6/WqasTuh5Sh+SMeJX3Go0Wp
5Ziqw6y8jIeDJhcQX/FWl+lqRDF56Jsb/erKBDgo25gww8JrkJmatM7TeXwe4Har
yCvmupnrZinfeJ8IQmKXzD6RXYUc2DE9OX6rhVRxrdrIWKOYCcvtGKB1STHYu5wE
C4wlUTAuV5X8PqilJ3+cqa5+6OBIKaLdYyfOi/Zr5BZjQsKbSQKrY2PJPQZwPAfH
ovXyASpL+flXz5wxVrG4CN55RcHau0nwbKsAxwlONp2ibdUA/zAGFNK4RuqQ/adF
TkDdWyT8NaOcAkTQTghn+bR5V/08I8GgjPAXX0PXIWYYd5BthfDgJ9Yk2hbfZ+1u
VcK8geMylCNHHIC/UKJiJi/LOaSyYFLjQ1OMjLHNPwKIVd1NIaHDWnXhqulHxVwt
QL9lXgZ80V/maJl3y6eKruvfCIwq0C3Gji1y61Dq+9+YrFtyY+qEUPzq04Bn8qRP
WUNDRapEbDGK5scGGkJBSl1WgH5+8dMKtt25rYz7qqQUIb8Mw5d9mDEu6ORpk93y
1KVo0RAdK4Xc37HrbLHONQV4gp1lsuWfmKn+ZOjEUm+6RmSkIQlYDa3s1ry9BG4N
OokxVKfQA1CqFR/cOzRVy3qz4Oanp3TYFViYEpkIpaRS55f8lTzf2CZJrToGvja4
VGR3p5SpO25TcMEYWaTftzVCVJBgt1T8qoBdFguqA7v5xQmp8dOp/ABgN/Vg+UK5
0IdSWg1TIzfCJ50FU/9Wb/WxWHwEnFh++DTMvym6kCw8K/12XF+XiK9pFS8yWrWN
TFSMmRomuPTj5BtGh4VgxMyDWZyjKlnbhlatIlqhpqou3uyO467z5YGcwrDVLvio
RJ8eoTZXTeqRP26Lp9X58RvMjTGes4EaND6WWNnSALRVZIugI4Wx/iydNEHW4mQz
ILZxihzP1kgh0+IcJUwLqq86ypayQpSz30s/pJQS/AhIlLNFxlxwA0leGhjDNs80
DPUJNUXdp2nsh43cakOjxLKPqGISX7Sy5FNbWBU37RODuIgUMUcKUO51HuMz2Owr
NiYYCYTEw1Z5IDpMVVbjMyuh33YezxYw1WMn+839RqwQfwxpgcoBFXIpb6MyXnqB
cbWaqBW1aclK8L0bjIA00/XxKqweLq87UAjfLnqfA7yeSSryGHvK72WtFwAhtJNs
Dxf6BkPs8UtlaZVQQziv16GKNvutaqKeGB9U8qfaW6zpVg/YWemL+cSI2WpUrfv+
oePI2eURD2aLRQGGbjR0VAhMMjdALAYW89oQ0PlvA1+7mnhC/S/CBlsz+kk7mIdp
DGAY7Pa3lZsN6JK9M0McNuO+BQJRHIQJYz1CLnY7SpYhMiaM+U7h9MlcuLiXFsFP
kn06ssQ8hNSMjzQFL3JrUEb1Mk9lhXI+izMHLa9IU7TD8X1oKPqLIsywYiPuz1hf
24W0k4lOmE4WfShP9ox8fQn6hfjyyi9WsEtOmkHBxYK9EuxVZF4PAt59KFNXCXPu
/ESi8vbJUfDnSuphFYOWn8pZNWxKAcB83KzJ584UF0LmTUvhFajKNgMJoro70bQ2
Xi1WV2PMVd5eUrECcwnOBKwIx9Yehb933wP0oQ/trkRY6J4klFlKPIrIqGdk+M1j
G0xduxv2DVJkMPMX7EWqT78o2FjaVT/xmzMJtK7H2qKLHSirCdd2O3eDSUzVHk+N
Od4eYZBNk3d7lFus6esOzEQHIgapNKk6p+/67Qh0kmZtQUJ2TaWluvzutBauF5Dy
41pRaevCSV7hnkYp52Sc/XYAY2r9juWh6MhD+XSOhJbmhrULLmcz4PbhHCUiiDVr
zoJnt559kSSxglvijvfouk2zrIPDnWvJVVLNvvGt/wyeeJMPex3XWtjDVtLnibm3
uYk0ajB2gL4Zh0ex5rTJbRQFyQUEkKGgh8Oa8D4iTyU9zWByDYYjXHn9viAaWHys
qQ6T3mFcaiqBsiH/SMMzg2Qyj87n0QErS+ebvtlVo2r0SDYXZvAxJp87xBqar27M
g9WMXpKNHjjjyJIm7vH3Wo1g9njO4OKgTD9G/ZrNuO+0IOI3BsqZmEF0gT12D2q2
w8O24E37RFEzT6bYJ6Ld0ekAjSrgWF/x4jQwtQPrmUqtkDEbQKVZsrw22hjtCu6A
X5Fc8M9MSD9KmNy1Te5iuM3OOfe9LOpYXPMBeaL1jZYf8bkmRBQaSouedMwvfRew
qfUVbHWuuoUf1OprtA1zKM9vyBMgXUvSHOASDUDeFO9lt4bpihDxIoLFN/tKgYSR
xcoa6NC+WkkE+/Gs8rDSKqwfQjgeYBArgAnElTgEN+dapRDuWq2HgE60mJwy5Tnh
RqSGVtgeFy/N7X+sAg21nfh0VGyJ5C4Yk6OlzQXEehX8zyoHf4MqbE0VJadgx39u
fDp3ShniSyEXc9OU4feB8FDrzCwAVH/gM8WvwdXMJQcZ7TD1LOhcZ8BoVaj54a6A
QYoH34JxdRNu7Du46ovqL4w45GQWRibQF/glYL6ENaDwhla7UlaOIxBOQRbKscqF
OYEG4ixiA9EEVh5BsInCpmrVkM/VW2yqw61L6HDGum2q1fBQx9vXNDp7eun1e+oY
FQOXJ2v69n5bdxiMw6aNrtBj2/on7rvPMzrdV9xXP6rn4PnkhGsqMpenTJ4XL3B1
U9h6BgVqm4IhnMo7LwozImFIJVHnvIQSeYZlUUDRpNuTyHf6fmP6x3hLhjERgeis
UoNdDepV0yWInxjgqCWmTQ6kau4RH1x4iEvpv1gXPg5DZYpImmLaGX74iO+mouId
LtYSupRG0LSwIzKmbkZS5RKSAuW+hGKbkvvutw2DsUjmmHjTZ2Eo8/Q+nVJJP1/s
W9H5cM3oIlX/AXMgyq/E6Uhp9cj4SNpvmaIPJ4SqXr44l13GdkBlTnHCplwTm2FY
E2izN5S1NFhSjz+pVWijYNpzIz28MeNN8dEZFNFe64t1IgAZbJozpKinF3AdY2e/
fuyFnVkc6vwBGt19q2k4/3iwFgFDtknf75NOzM9+OX9lHoiysqcy9rcSRcAn+IEk
VdjeO3yV7NWRZe4Q1bX//b8ikbN8CMoa248JGvaJOxCWM6IldsrTqnAdu4F9Cn64
xRPZdVWS2c6o2e3OZpU+ot/tjZTvjdFtzjy/7RL2OE5sLrpOE5t6iQaMqf3CQnCy
xJVIPFqTqM2exhC1diMja+j2A+ZhGYtpPbko8ErNUPFtvLxD56PuNZ2GxleqX1uV
y3BSPR7JCiFXkntLXQODVFC3dHRMSCrkr+M+AZZf+3zG/MtUHGuuANcNdmt6y3j3
ykYM+XvKrUm6dc94CSebzpGeJypxYg6l9FeJn8yDYflbdvhR53EO45Ww+nXil/Q8
MqXhrfnfjJFIyM2uTjTSnhssfQ7nXdDdRI7wagn8TW2RBARQzQ5lcDij1ka6ZLK5
2gzQak7aQhjWtwWkEuNF6eARPE/JsRIHU4XQnwGzCbzxt50FR9J+a1lJtQ8y4Xon
S3nQX0uT39AyQnC4Q4d6dO3ANRZIpLeEQrU3Iq8eOhhn1XuOYdHk2T7ctgwZsESd
0ACKD9al17DGNU7ig8athOj59TaBAf9i512mzmE2dJDB2YqVxFP2OdcN0zIVZeUx
MktXbTWFWPRbME/AsJxcvEs3b0gf3JpabspvOGhQ2337kfTnlhJoXZ7jWh33/0nJ
BiHw3RZqWdDqv0BOx6d2ZiTczDZdatPWCNG14dJyU46/QojuwDOo0sWt1EJtKQt1
UiBnPAp1+pOTTWtNG4vRGcNmCpIP+bWzwlaohg1HJWLKgFIjLgq6tKW1A0ArUhWh
yh11ioFV+Fsv8jHj1DzQvUeoym4UqrtVx05IOIS6OlH1BpUWYvmWxwEUnNK8kV8S
mHYxxH2daM/9mdUWfoUzzVo6cJMwZtUOuh1pQ0b9TT07BqC3qXBLCHtU4gW/AvJa
u1He8XodPHMr3IEQGUw72ZbBZ/C5ZeHcZ3wmb6txbjz4wDA3fBRmvnLeYLlugxmc
cOQ2olkic8RhPkB3kygxNO6HeaUfeGxmwxXqWbs+PN7vkWdU0QAj7pzOpgL9xTSY
ydPFSD7fQydf5p911Z39m2PIV7qP+sy+M8/Yt83dlGarIe9I2pYwiMl6MVafbXtx
uP7A/6gZAeUl7cRzDTN2R5qlmoDwiF8eO5sUO9T06ZIqA9f+0Cr9BpI0A4KzZsAP
yFL7pr+MyeMRkG5H4xnMROOa/TrDEdZ8uIRaVH0TQU9wQTJKYLrTpjthnC3v6NOg
a89BcGEomO2hVoV2/PySGfXx4ZyPfQFA2yE5qiD337acFwNT0jRWKkTQIRh0eRt3
5s9zl167lKsquY4G4YV8Dw4gnsI615lFrBt1RMitEzjVWxGSIOv4p9K+Yq8LbYf0
jaY8g9oiclBqhXXMoYLFG9pbaUCa4IXDgPG1ve8cK2vRZwAWltbjeCLJzqBGye2D
3oaSgu5deBWYJnYqfFHbo+uZh7aV7+xpW2XXEPs/DWCIunkPpWgO4qvSbpD2c1jQ
0qgl14PYXnIdcr4g/QU8uUqADy5ikFUToyFc2h6foJAui2XWV55dMYMyU7wpxNed
atJpmin0YUCNTn9tlrrDjfZuPpT5DNEpDKFnHecaceRlC4etr+RpYO4t62U+emZ2
WM7+kpCdmcDQlTdTdYOI7koGtVF4WoGW0JH6BkFggkI7QI6aFGKH2HZjHWrhEO6X
Bqfj53AcfUgLrTTFI1BRg2NPPflLeM9cBWpiU7B5V0584AhcKZnXdCpbD0n+QiRc
yAWpTxnG+6aq6Q/zyafwzZL+iN8RyLZc1pM68WVHrAXuKKN9eaj/+DrKMl8m0VAG
4dgq6wER6KoQ9BRxnKEAXJvJbTLL9kQFjZ0uD+IJm7dXA7HOOLgxONRw5NnEgDn0
JwsBTiiZtMyYaxXx/KrP3s3O/p/7mv8lGHVtQ4Uepro3PM1CmuSZnMXlYLDnxTNX
PsZOOtDHmiq7enaB6ZtwGahINJJka6J1q83C/+l85zkFuV7tsRoXmBGcGCjdPtfH
mk5VvkNOYDblIzigv2gSNKiEWFUMeb++tWEMFGne1MZ0Zrbhs8INTZCGKqrLiJNe
8d/J5yvqhVs8oewoxny4J0ybZ+1SEfxexU1qKHHPBPSUAlDrJHWF7DeuXH88M1xG
7hE3NdocwZ3i9eU2cKjjC8x2efzksa0dbt6W34f3O+JLw9woruAwUgpXcfmy00hu
/O1F2lnkLOgCV+QZSAMvdcxGWa0y1RUH0/Uqn02Q2hcqnbohjzUf5qtpa8NLttrQ
1zj0xwSur6LmpyWm6h1EBaNLmLN2Zfed9qAy9/Ogx5JXF3VD+hx0HYYA5ccCGZP2
n437wC2g2Wcanf+F4ejMC6wLKuagHGc0qr6OwZcAQk9t31ruRhIrNHThd7xQHtLG
Arh75sWlQ1McLd0c+sxhu18HaJeBy4MYrKGl6LDjf7gdtgZtmpsud9DosudPz82C
ilIgBLCYd/Sq+FfjgkB7tuuPgi23MC5bvXQozkZQAS+KRcoi6AdMho66SmH7NKlc
qeRWAc4pgFs/AkkrTc1dZsln8NPnA5TaDN2vI+U896y0ZLm5d26POCK/vfly1/Bv
C7DWtqpmCouMJbGAlo03n7gl/xQ0cY0HhkSgyz9OOSe02w1h7+hynqx+AUo+TUng
KRTs2+wRXvrTVUFGPS1B8D8IaCXjL6PjeY90wguuNIpx3J0xfucybuzyFjhZLOZA
IaJZ/tMjBTL+W6A5zEby9EXkdo+JFnvHR5NTlFXA1pASTxJr+7RYLcdF10XRvYzF
I0dq3TD+XN2+VkGT5Xct6sKlGMuS25Iv0ijZ+pZ4VJCgzdd1lNfwNVEy31BzvLCj
qxZw/y4YmcNL7pgtX5/oRCsThKl10UieDMDT07/lV2Ss05TdVtF50+MXvdWXjQhb
aAnSbHNY5OtT7aQopTpftXz3L18KBa6+IM03bEAnQw4qixsP2PdQINPNC7rvudLf
p0q0BmKVqgxczviHKwFYi7cX+egKVAX6fLHZRBmxxDLSinkcc/4yrYdRFdVGTbdM
CgSpAqQyjNvuB+HKJoOujNFZ8y4uz56BEU/tfKvwUJQBcce+lyQqzQsI1kahm9uB
sU8Ztz7dC5z99VsB/EojvF4DYtxBT8q5AtMwZwF9+s+vyrS3yy7sau5Mfh/W7PGK
xO5cT2bZrTU01/kIdi02arrdBId99WhRgPMgyt6f+hgRVPjJYn6bwO8/tTVFpt32
SkU6spjNWGm6vgRiJFnXEEKr0+hsU+ZEwjuqlIMTTERxPkj3GeJyWnTthQiqr5y+
Ozp/n9MYIzjgr37AFdgRbICT9+NvcN6WurGjFs4td/+3/CRfyfl42ALVHgb/9l8u
6fFKz14aaWbTtXjDph14v7y8jBvGJyYBnBB/oWsx3Hhiat2P+0SpZ1ZhuOGYUjGp
pBsTRldPi4rX6puas9ByUSyxenpt/oELRBpEpsk+S5iNgmdDldmhMpLD5J52bpiu
hNa6ureLGA77JeIT+I+Cvk2Ot+uHNu09t7ydntnB1eD/7eqIcl67ONg8gLx/fVDt
UIgG8tbV+Hgg7QO3rZ5jeOWrcbet6C+2iaKrBUVXc8UwFCb1aYJc6gwxwd8Brf8f
85cr24LitqZ4o1GNjQI3OYAJPuHUmnT1rj9OuWfczSyymVHbBgA61l9fz8MzzFLv
Kc5WV1eLmF24UORjv75s9brMY8b5BiLrnMXQfHG0+SLZwTeMQnKBwpdydi3ETrin
VsVN5zRnaWnhYK/Q56sQoYIJmfPeZTCsCd7lfXtRIZ9H2fx8lLVfD86mmmoHChF8
XpVOjB2/DAzjkCLC74HEiaG16osA8/Hq1jx201xwNd3kGzTyu+6YyAiao9tiiddZ
skyRfNy8kxaUbvki1wrkIenh2lybZPUCQF5C4h5fhsAFahm5J1Xyc0ERvZ0Tenkt
lNSfXj5wodEf25aA4X0P2VESxRCWN3cPLrOSZWOcG6HObPPvom5IWmntQYNcfDuk
f1i7l6J06f4DarSK8WdEu5jCw0okgSlDXvHx2QSrXv8JjHKbKg52jWX7ekx04EV4
q4E0kKj8uHLV8i+84rW8rcsgFJ7FcL6FZdsTu0uC62L0bdFssIJyKDjiA/zhvPRK
EEvq+Y7R+s+SbcBjwwR0mEKgpRE9lVix1WeW1mGhv32TCHFTJWJ/VD7FsOUR2s4j
3Lrj0vgGfBoZWg6K2nbO0r4CtDxZVcXfTpsctlKsRziMrZjd/J696zsKSAo6Fb9Z
Pdo3fjmcOdfR+QOMl0PJR6gFOQt3f233IBTfbkSlz/TcWFB/3WZLGEtgc+jFbaQB
JoQLeTR9zex1zMKibPAe1Tm6dnABcug13fQFOiNmx9cC4GUFFOG0dMvwmTcOZTQr
omu/l3ZKBnNm/v/zLFFg/6IjBPLGvi2tXyUGM6K6SNJRkdllqC4+0Pyqw4FI7ACv
AF52QBvbEuGWw0ZhFi+PXvRaRrkglMBHAPPOcRa4QhpBCJ92N39WueFpXIzgwyHl
EW/QGqrddR06/ylon27Np0GRJFIiTdXIQpaffQHVvjoURoGr3ASXUTr7779HITys
nbjazer2dWHP+6m7+gH88dVj9yy2NKFpVtmWT9dVK+IYR7hs4c4XWKoVR9JExShx
fVBa6o8sq6K/L3dhpyiah7A2P5UeIcwJroaxceK5D0ZTeYc4MHZT+gUn+Koaw/We
WadciRmy49Vy1vkSMz8c9zfxItS+lfSDtigh76lWe67ezIknce+DPJNn40tDzZIx
R2La7jSCy3qFauyNClhqg3lnOeo4NCsxzE+HBFvaLoFZFK+/5udRrH4fTmqLsxsd
l4YzdaN6ujqL7FQ67vgvIO5+kDfSoGDk9hBCS7oKwA8MUSmzpL2/WRYB70Ja2O7o
/CmlJ/FZc6Pi/8JiAzID1JMiJp3nlsh+XKp468n63cMngWo3awNAeFqb9FmjVHNV
WvckgHQBaqZdeQEZ+7oyUrnBmTVTJUp2sr2TJdrLELjKGT4bnd0P4wF0mY/HOgAY
TKixjGvAbx8Ch9X1xtV0lrq7h0POrr4HcuyD+UBHCAEPnIKmBXF/y3XQ1qitJvMI
S+co1fFnigNAmO1iOX8JyoSuuUaWOK2C/WmHgefjchu7ynBmqMZpIpjJO8vmWvfu
/P9GelhjhCpVa5KWxrx7rg7MfjZhn926CyYjNr+nOyxvcvXvEBlI22NO+6y/gCp/
QPIbhzyEPPAuqDGX34DT0HYM43SpxIn2jVttHE+82MstRh9k3bKoYaOkfLalRSLk
zdme2V+Cj55RGCrRra/9XAlxooj8GQXtRXog/88TBVp6IxDTogF14ddF4gp9FoiY
taFtobFLLi25OL98qyydU59NFV0BsvFYPEi1DMA92ST6bahb5zP+F1H+hN2eiT/m
UxPANkVnIq/uTt1hudQXZd46H0wWswg4qxmSWm5yAR6oRRUQwNhRCK8vtEvOLah4
PZk/oW2S2MwswbrJzaL1ioSrMknhnctQrVAbzksPYrMBe5zEgcZnuXlXdXyDDjen
AYQfRKX0qEYJx2Xkg9uwnZBKDM05yrPtv9JXE5qxq86+21CvfF+tmX64Z7onRjcR
fpEqGODTLTGkL6C0pmzWiI1WU1WBdPzPVlw9djcHg4SdpyCcrSprmmKG/rXB9oZT
Z6ainC+LlN4AMBZMxY4V9XyDuGL9f9Wanfdcd1qlCsD5P78GMekTxeE6CsYovBA3
fZ/qhw1SkM9wN/NKTEEmHQQz4iJ//y9BofsFCXYLZYkRoIR9G87c8bFeStWHthlO
GC4Qtx41ezBZnP8ik2A/Vm0MKf9ltN6bzpUioUnj8RqZwY0JDTbUfsdaI0woKKHS
PplWrro5wNloj16XFs6QMYHmd7K42lR9Du+5Cz9R1iNIshBNkSbcOpBOW6PTpF31
fBUYYaMtShHRvtfETcTEAcsqvGSp5P905h71XvNPtQGWIDLbdPWNV/9akzSDrz00
Y5pQ7JcaIqXvURf4as+r4Ddo2tGlBAuz5RqqKphHLzTD1bI43AVo+URfjqfkUubo
bfwrP0Lf/6t0oK0PZNDSHQQIcTNwZ/WqUImXzMefE0WqYX0ro1lhhmPBwt4pzdVx
ITaKJQsRzg/2E+BFpLpU38OZK1M57o2vXBlK4yD+davXorSIJbctyqIOMLvMxe7D
P7kreV2CiUu9nE/rNWfApOZYM5aaywHTFlcmDX2CdgY9QZb4VWn5d4DA4PJ26ycT
UY5DISwBQ0rApcJ8WR2T6SmEQYLmqjwfk90wTDqMdqfXcszTY6o1FyVt6hLfFGv9
EO/JsEr8s4tTbf89UOF2S7dbBcOboOWrw9305+kFFj8FtdwrQfFVTWB7++htPNhX
oUSNeCDl3PpOyoldSQW0NuSIr7ogTm6YCAxb+Cz9l1UaBCrRNoYPivniQL5lBT1h
+dsEgUiojw1vnBimgSDBGDJfBNSDHCy4ikUnEcqyaDwKE3tUxd3JFx+Y6cWq6SUr
SkSPe9gHaXLAS4HPDRxdmAY9qNC3//WRzzzy7IIT1tMck59VccRn9ws4WWHqQL9q
uiU8HXr24tc1DR4Tt8htbwbQl46+1PhUj7NIIiUcUcId9uv2buGWyaVzmGqBG0vB
Z/A0Bnc6IsR+FFnIx7EiQ3ehmUhxGs9RLt1F54qay/TEUaVaDRZYEYqWsI8nAGj6
smzJ6M+pStXX4YtG+H62A/ysQkxlRN2HuC8Wztj4y9K4hACyunV+KDnpQHxaSwcc
LDNcsuAhib384iEOG+nblKFsu7HfFx4SxuYXYBpwJM3eTJw+G2PDWje3GM8kxgk+
ani97tFDJnjWBDY5IJYUAuIAGeTssHVeJyeR0tjaIGptdredI4Uuj0aAYXZmHdDK
6VoNkmhjk0Nt84S5ipgnbx83h4ck6m6j6nRVpn02riSyZqGQ8IIorhV39S3AvquN
79y/AuxVzTmGHQ8juSsDTkisHIiBTwYSGfMPaGeVpcHoKQNb5B3pFegaeY0gG4N7
Qh8krdW2PLD3JfTOR1QTrBbb+GC7rEAz4uRRTHE2ws/4+YrqPli8i+PbfivjLrOR
BMK2ceaJrY2zDSdBf8FrI3Jup3DdCcjxynsAXiNiCgpykgr25+CLELFS92REJ+W1
XXPhFwUPHIh0pizdzD38ZkIfx7EovWUqZlDZrHu7IKKbRVTrYedOUYD9+kBtWf23
oTl6o5AHfqraTotTdfZ2fPdCMOtJ64k0UflxPzSLS9xFnf5hnfGe21keAvv4+ncr
EYP68GHBPixHzwtqWS1ohnqxvMCg/7wWgahyd7kNtohOi+EVixZQyD6vJdmYIwHL
ir62Y7tub/kUgXCnMR8o2LznQoCObrrWMI7aUztlkBp7a3HHMMI6+ypQD3NO8m5q
cSX9cF2UAa7Y3zX91zA2Gf0FA8+CKNome1LUGQRS1EdbZEqEbPxti32+VDbOsqw0
6CHkuBcQttIzzI7FLY/4Embke7T1pa+k5BgS3xMGNOx61ROzU/jA23YC+V3LqCtI
MU6A6ts6tgeD73BnUKfUx3orQqk+sZglleB+xDjblk4c/wrB47uMIMt5hiVCTsqN
zw97ogz01KhVp+1644dv23tSAbGGdlUnaTEpoBkkeCI9XLs8DoRuiyvsAqV9V+8F
PAJ2HJQF2gVkV4cJBy5FT63W+c2oW4xsNoUHsS4wjYvyiCRlIqMWZ5+r0FFycdbH
gmT57NVQenigzaf+dqPeoTrEDPBSeVyoQqnqIPtkcv1poAzPgjKt9RmT6vssd0is
HqU10tcqsqbtdFoHRC0LqLsYy70tETorEkCZ9LrlABczFKLWJ/EH5JVo01Hyg8kA
y48TqsMUToSOfAT2J6u+kfXCxOTBS9AstXcNdr+7DooVb4fULNohSniO95rQGJYx
szseNVIjQe7RD4a6ly81/RRdasHdz9UsfDrPFdnoVHCK32SxXel2QiyL6naRKDCb
rylkhnGGrktFmzQJa+lmFnlfrGWkhoQWcOc43UBsIKsEKfEdwKFJFY3sCHorZ2jm
wlQcR3XS2nT9lKc4X09mDoKWx8DttDBNyUBzDISIN5ewq3BaQGC7epHZyn8d3C3g
8bmHX2NBJeSehSUFdvMA+2np5mKn3iis7WsDM8SlB2DHuJO+h7fUGw2X/0Len2GG
qIyUN0QQa6BrvzWOXKk8U6rPf6up6cvp2hH9OGKII0Oi7XGumGhClt59beyxQcHa
pGdjD+ly4OzCojSg0DU90t7be37xoAr1USum6PSIUQv1gkUFXHFh1k0kV+O6pKmi
LPbO68lTpoFxJnqFhr73DfjeX3grbQC0VTSTvftVLUBO6Vvv8+Qqf8rPTloUMDlj
ostrcBdrlvJZxYrV63aCVz6MuXKWleUGAqbQTqL28vBfje8L3sfo1zvjnlP2Tl1z
kscetmiLA5rA8+xr3d7k3wTng+H+DygLnRptJfj9Ju2sR7vpmlj/Q3dRl0Ta4nRK
akAg1CkRbZBy5r/3nerw2XVvZVWWEL53vmW7hP9DoP8rK7NBl0DsynTPW/1M0Xk4
dSm/S/0OQ1wpt4Nj3d6rz93tj5NnoiQuWa8RG6Nl1kYVPh/z2rAUJiEybTeB1hgt
jFQ050b5MQXpxBZjgXya1WdnviaR5AT0BnwJrB0pkVfjYCAUugm6dVdh9EBcxl3q
PBGwI78G/FdvYR/7JvLZcCOc5+uUqWr6thBbEVde38fkn7Doy+xGPuSYXqo3b+wN
yccLZQ/hX8mz9mW0QoYNO6oxQym6QL6fdvAKYb7lfC9slpVAqOMwYB1MaOPOxamG
h8uI5abHLGVYdZ8C4KalBJqcqPjdJLBfFQMPMPo97zb6zlgN8vbZsCbXkRhxWC4S
75RypM+daH1/H9mpP8xBFzxLLlSgkp08ooi00AFiHyDbDHnMOOWMIb2RNe/jiDGi
D4YtUJ3Mhbl8SsstipgEpJfHVe2ZR5sgbvHTptUM1GyWDrbh1miHG0wC+quRurgQ
08wYMPQc4mqWCMPH4CWUS8uqGG+wfjjdbs1BAu1+3WumfwHm/Grd6wI30y/96oWL
cDNfh5PcEkAq+hKmvAvKYR+jkdN8EGvBg17Bah12jrYxvT7PQ63QD7slT5L4+9Iq
HIX31VHim0qIIa/FQtBFNH6VixDPuWTL5QzQbLklV0dT/zW/jjEIcdCmUBtmLSot
pPY6KEs3sbjp4XC/+L80OdS13zbLx+TwtbMuHFdKk8+SJQWH720Ol4j5dRU6DuJG
beaVupft8O2m2H4NlLd+JKBVaqNgIJZsfRO2zEKzSnGAYlHA+o+O+pc/pWCeZ2aB
v1h7V+suzrw4fm0SFHH+4KUgL5BGg++2hhdi71UEMR2ApGrBnviDi7F9yzTL4vzU
j3EQqUtuvf0vAEnnkvmuQce1pXgQ+5Z38WQinEyx4TtyA5hlN+EVicUAzkRomZk3
tVIkpdeM5dur353TAjHA7uyjkaWeWKf8BJiQ1wt3vYY07MtV7cdAHm8ozv9/XXz/
i+fSXP7CVOWpIfb/3Vx4wzKe7BMca6SlWLR3mbGqt9q7b9hVdRP8YIp/Np7fMfqK
3uI1pfpxwvCWgwt8UovKE9tBH0C5/UkgB44LePz0KB3OLzKoVLdk19OpsUhzz29a
mBgGtVFMbA85a3pmBKWlKyrWJgY7WbezAkQEXFW9EXaU+5vDRGHnz8L4vPJXJNpa
90ODf4X2YbbRuQaK1qm/8A3ly7heY23U2y+0zmOMXz1nZqmYM9yUWhUQvDNoiU16
Ha+Ermm8+G0jnVtD7xun6NzUeyJLJVgh3aKcrbf7Ej6jhr0sDX+5bugsroLKOsTW
4VjmI57MmXpzBuJ9y4CNai7D4Ww3O4OYNHROIyqjv/6XotP0DDLAz+ViSkXsbctd
/LzwstrA5Mu1nctRHMUUZF//7/tEDKFDTZjtuhRntxqkzv6BON/hIG4rJYLbFlo8
7JH4rI7W/FU/6891Y1RbXPKZJctY1hrPt3CcSNzEerKKqg+U95W16/P+u6TzLAhn
RHi9E+RZUxN1+rVkPpLNls/pyPAkw/MfGeBtQGC3CN/zgMa4fJQ5M9shqSISu7gq
v4NWqTV0CauFmf8AaXVvfa/1MK3xPrx8omCwnjmq2WRUNoGC+v57KJrMV1VFJZIr
Rf0BAphKvXncS/dB/W3ZViB6CYY5gNpTJk0JFg28hFZ9gw1+DkDebmg2bkzQb1gA
EEdcM6JzO6lnPw8t1MtnThNb0rmN88CFxvg6J7Fl3Hq3UF4Tp66DhC1hbubclUEl
2rzlK80fAfVQelWYB9ViY+dW2BnVmx2N78F0MQa4Ykxw9qZ6gniztLVzWMW0opX7
d/fk3bcmjkmuCdhSBB6zYO/J+eCY9hV3VbDMHoegXjEOUc2BpXiS6Hl94wATNi3t
h4COWwlTiN4hxB49v45DGG2Z1CqS8bpSZ41X9hsLbKmkWG90zBfNFNHeb9W+eK43
J8j9EXLknPcdO1l+zOBtCque6lR6BJsUT5wR6E1Ndn0fNvOI17hs69UJwx50DyNi
i4Uf5NWSzG91qfVaYauendnrD/pB2uRVa7McrdPuVNw42fQUxv1URN+jC4rhFmRB
YdtxK1/BRLvgvExq83nL3+XSvEZLbZJSDj57wn03Qc9sRbFhLKt5V5iDEwRKfKSY
9faRiPsPEEqzBU0eBU4/HkMepQTbmRj21mHNCTHBERWLAghJeZK/ek8z8D3pvT2q
kCgFEzf2TxtDSfTAL++9vjzTVh0uUAHqxBF0oENlsdhYaRbvGDznK+c3gBUSP4ej
ZxYDn2Mq3esm/QQlVFYKsuRemYKEYbLbZMnU+a7ovXpqjcd88w8qEyNffR1vj8Xa
C8anghFY1pe5n0sORjzVzMAKI0K/spLDPysNApPtQHfnvcZ6HwNBTT2B2N064DGK
IxKb+KBvfY3HgadBW9FGbwHZ83H6e2cXZNB0hqyTA41kr+WY5+3yTSDsvnxg51jI
2+RU7CKslkXQuWyC3bsgMC3ZUoZDFNT6UH9u0etna1q1AmPC2P1VClanNlntYKPw
RThZ/1O2wsUYOPTyiilHBXEf8c65p94uQd2SdmOWEnBopsTSwJPzMnrwfocW0DZO
FbN+1IFHudmO1Jp10SNEq8e5ZVMkns+7sGKXwfia8TbrVx74yHu0mRhbCpQYiD/S
fw+6A+z7D4BM3/RQcrWpCXmS6QJUcvsodufeoEZui+3ew23sVk9Jdwe2EfeIc3rT
Q/mX/5YHysVj9SNg3qtqzEoYkibfrZQJPlIcoKPIMG8yiUSDu6u3Y3Pw288f+GSh
QZMob4+vGg7adNKkskcR//zKlfZw2XpV2y2H0l8YNzY0xfrmqlJfSDt0SalAj2Fw
MBgvnH6ZlHxM4jR4d0aHffFSO0nFdWhjinv7wDeAvxi5h+CBb23FOhg56yj/LmJr
3povj2ydDFiQ/IPzbgPYedOkkB9jEihigaww+wKWBlfQdSGgL4hinzww89wc8+mw
PyiKuJ+omQLrIqdp/AxSm0YDR0HAF7NMAAkGsNpRja/mDZAL3jA4URBqxrPp4ZZ1
P247CudR762HCM5Y64mErFFLmIdAoJO3pjlorpD36aZzd+41LURPV73UdboVhSjp
8tjEabucIbXMLs1rzY6Z3SB/OIOFI9VI0q8SAF2Kw/0OmbavuYiti/ml5aUD+8df
PMu/s7s3Nb1hTWgT3MrMlC5UJ6A1MoDy9JSwuqf7IFdjMea+jlRMu0NGJaKlhD0+
lHrM8eAmoQC3sFqQk9HIF3bkwTeu+xhip4zEf7Yfj0Rr1pGHtMw0hSAK8MhAWT89
QRrCtCRqEIiN9EzM0q2USSuFCfxIkw8141TuJ+mNavC7NDtOAIT5E8kR0DyreEqG
lQQ5T5EvWIf4aVRSMC7w0fwwQiqvG/Drj9oRyJ6gMP7hSiD/+JNECakDGZHnYwcZ
pb9QR36bdfZo/dSzM5fUntfsvwgywNoG6hiCcQ7ZNM9h1ekSCsFzyDei5Cn/5X2K
K+5yFzHwQWRrXqs8TP26bE1StrDjC1FlMlfaaxtfP2KLdcD6HEaJ+R9uZEaP9HsU
4cp2ybZcfIqMCppd+B0Ruc84pdnGOemCKANhUFO2CW5QE7UEka2C2CbNjeZfHAC+
z17s6p+PROKdrQApFCi3xDnzgFx1et7UOHPmF7zN3g345T7LcbUxroz0z+FfkDYa
u8nPysUlouGKdSAZQ3aleKoebRe356iRw1IP1jdJQQ2vxbYMZ6TaqqN9gdFSHFX0
s8XDYiGw9U0dkndyinnsq7EoOgUc1Vh6VdRgd8mptL0LBC6wpAAdM9YUEh44csRd
b+LQX5LZhyWmKRBj3xHjDC7NJ7Jl2TV2xXkBxeEWmuX4vDK6Zp0OsB4FVAWZPs/R
JwBolLCV/jf0wwPp5lvKN6n7FePktJXmfvF+nbwDnAo4BBNnva/rnzXcv3A6t8AL
7oGatvUWf2tOwpI3f9UnLQ6Z0AeOCA4GSiL4sxUII0NjL778oHe78jTVBFjZGvXK
jLznO+rd9M4W9nrZtaxRd/z3FJX8dtJUehR8DrzTeFc+kUPbjTqsprzKmElYSGBJ
kYzRBIk13STQufcnNdWoZ/hec6PSpJinHUyNtzYVoKSWI0fGrbR44M+/CafsQr1L
x9SlQv2G7t0DbWcIit4T4u8/C3R23AHRrSNimXq/pKHLDEd6ocOr6Bsui4bzWIK2
+cKR8vYnkVbnIdH7Ycxj98EVeMy/7HfgNaRTq1ZMLcGYV8BRvJr8XlFb2+C/k+F9
FoDJXNtIPaug7Fj76Nivvxcx2aF5oz2NIJczW9ycsaCr6m+d01liuKbo5+XBL1xE
G8jsHVsSqh2/CtbUnoObO8JRjEzECHNTI9a8X9HSyDCrMTpZfFhh12P3xqXqMsuK
3ab4sWkV9Tk3fBoRcKXGaJMJ5GLWwr+Rk94m5Od4iKi7h5AzkdtImOEEuHwpX+YZ
TobkpeDk8nlAjiLDzrC8MhkSPgAi9jrkdbzTz+xxD+QLTH8D5ilm3YyhOLFg+4u4
7pWgNxOihMb6vzTZ9aEqwiFxLOJPB0GNVeOkGqIo+zJyGrWctq1zcZv9wMHBX8e6
tUlG4FkxcKgZIF6RK+lCkEu8UI260uYigjjW40roEU3RF3fSqi2JizfScVIaxrSi
YF3fCMUwCvxQ+cfDXYrPjn9Vxbig3B3oDoTqxrPp22oBNr8xs8GoJ7mCiOtyE2/X
Dxy7pjgC9hlwNs7Q90VSK7fqSEooZ9zGg7/bku2dSdRFhOqFEycO1Ln875HSaRv7
S/sAGHRBhIuqlWTImxNZn4MkO3zo4KdXamMs02h7c18Uf8fEoVvcWxnlN8P0Npxh
45lq7vfhQZNRl+kpHtLkggvOGkWfGdxuTFW2Qtjx9FqFpRIZHyVFxMbawuie9fsP
Y7crFpEAWEsEmzzW9806XRkXlnAj9qT9A0MoaU9F2VZj8Wgv1r4MRggwJdvEDBxF
QoTmeZoc3e6bRL969UzzagAOP62RXCnvt/EO6Vx3cBAKucBlbn5D4oqlpOml03qC
Aee68hkXzW3TA3SmF9vgwFepBq63VIRCHplM9h68DCGhEnZOZEVGb0WvyXP0xNJa
+FTWQQAQtxeO52sfNrsiELmXqges982gkB4ATCgfZEKTb93wJuw0HGoeE4FMR8Bg
WlmQcofzsJHsCAjNYmi45Pbr3Qawh9EgXVxJPsowW0QjLvc5biPQ1znbzyIH3QyM
Pj2yASSauv1wVxxNQQy9AVq/oT052OpROj9O2An6IqEkqtvXQLbVZ29k3AVGukuR
m9VRc6qudvOlC3+nPERI7IAJKg+DtXhhQVcgNPyFlm+MkWJBrdq5m1Qk5uPRC+VR
DCzA3bf/nTx8Fr88BWcrFjrL6am4roOPmAzUF2GkOLYC2aHhFw0QohpZ96yT1nlA
B6HAkqnBOPHgAbXqV/H3xYbCaVmH2tYgIK1Ety7Jthjb7CHnIAou4/4iSs+xa2t1
MV0pDJPBN5hzsWuIzdLqAVsK7gj0SVj701LubMV9vEceK3elZIfk0xqsTnS2tPnB
O94/jiPzE2oZ0LL51G3kyeUjJtVPzE4srjkoH1HXKiw4heWP28NsFBaBnwnIsju0
3kNrMxczUR9Fjmfx3Q2e45OroA45H+ttZ7q/yoao3oLTkZkgSih7oAaKxPzVQ/p+
xXuafLiToZYtMNQz7q171Sl6xrkpZyjcL2IK6nxWJTFqAFlp2UKlSAbOATn9geHX
QSYZg1rtIET4I0cnEUcnEhJzaBh4ptihsfPb5IM45SwIgO6bz3TJD1h7pX7cOV51
C/Zk7j3soyOUQK7+gPVKf6GQhA1OmHbfS3vgS60UemoATDIePlv1iWo33OPtLphQ
B9PGIAVATWolaccn4HoWcBrX2xhpdfVBvRbXukWeFUhukgR9OPcfw9GPh/KtSQFR
NfOS0M4Ctc9IYv/mkr/4XpzIH5z92FUDuewcJFidoNzouxolEM+Yg088ovk2XnwV
DFfs7yPI23Rf/m+lw4px6k5wsVIb/PF+SK+919yt6AJcd+pRZLnhdkm9S2tmjAWO
1a/hGgaj6YbWoRuZldOpPKpoP1MV1f18X/xPQH/tqJNel01WGKDbSZljokIiZbRV
WTBP9wElY7qb5PYA7rNYxyTN3R/bZkiIaq60L6I617Nn3CJ96Ps+QncK8/o/Y/xD
GQUC9BhnLBunAahpRObunMRCpTphvr3lapHCFVUsC7H6bHA0aGkmTgdv0oZxssRm
zr9SqYVD6Rlqq9/u29zXDAL+cWHHTParqgqj7Nobbca4F2B2YwJLDhhkCQaY4vFG
bBzEvnVQhvCN9ro3MB0m3TU/fqCMhRiC6ZtWtFne2B30whdtinKsw9K9rkabQHGe
hqcWcw8pUk7DJsaLxyXfTCJt3/nxheXFk515gLLAgkjq73B5r7T2Pa0Ib8OUxlcK
4AiZ/yxgnyWKhp9UOR+XmZ3K1iFq+F5RaLqYh95DEgWSyNAKpeHAL2zEW1VcB7vw
vaenBEIiFbJPgdYO2GuBL4wgI1ls1v+lNpeYq/8O9jMhCQVqdCn3B4683zMc2XFH
lX6J32VPEGt58hF4AR2P3QkU6jQH2oaMloDuEIdTZlSHKyvzNCWH36vwFp3QZIoC
HHKzkkUoMAu2NWmVR3twpNwMq93tUJme8ydltscrEmRooW4eM28Unsx/xHefT/Oq
BisMfmTtqhFkAs8CKJawYgzIAiTXeKLycSfEPB65Vf0wfK4YAr4ERcoV9nB58Rbj
9WMXSqyaSjffrXSLaSgF35XpZEYWSUEu3tnlxj6Fj7Ucdw1AXh3XUb1cJ4If5/YZ
qPyxtemXyxL4gSeTMXgRoMMLuqqCeNADEjIF28JIUajBhpQWSaqdDR/I6BbUoik8
eCY7rFNDKin3DqzHULlIrmpj0w5JzYrhI2ETUSQLMA9LXbdjmpCuZKMh5iz/GFjb
pu6qbccvv41ezEKO/n+kSO4B8+P39OIIBvd0j/5f80eC9VKrKIbMNvTrX260+t3i
VaknGhu35xaB3wPv47YNAoDSKgdieL9+5upwYqn4fa71j3t173M/nEZH1fcKOJrZ
nuujE3Z2DQJ5LVtBHmjlh4HE83dBb2oa4w8iTnKU1NBdcq4DHNNHDdEVuRw8WXam
oChnJNeM18y9VOA00YLcjSx/235wIjTMbdi+a1tdyqnJ5N9u9S/HMlCnsJVE4gNY
nPeldNyCJU1QQfvAFBegXvb/kc/mLSo+m1TqYXhAaC482r7L/1bKqRA2ZOTxMquk
w1Qir8bumUT4/v7Vqvptd4N7O5D96ByOGGuccoSuCoFiFMZATFq8HM6M7/ckxu9/
tN3ipnbDyx5ITDPregxp/VcwnAdMXKUOGuxHvwufGzpboBDR30Hsn/Y9DYXcQfSh
lO2oHO2+HSxR72t/HUPzKLDgxQuMEx4xk6+r/oKd754T7ZSWXmxyxDm3sdnNbwM8
67vWMqPW5XxMKE6UiGUmvNvLZXrv8C5Lw2Cp2aA99da1dpbxRlulUd15Ta0+wjb8
wf26FHObBKgF6O9RKqgcmPL64Mq9g1NLzoL5qyVGrd6EoRqOAJxBORBU+yO3OD3h
qyofN83Ja1OlaPccRmqcgEYopVNmSwSvvZcqaFheIIno+RqruFoZr32wwZtT2csd
oNDF9Us4hq2cQhSKc0W1sD8PxGLWQJbDhv2Sg+j7qdx8a/xx01t3EeJ8UFLmGZDp
ostaiF7bydO+CiIxqKi8WYtAg6KLurJjpNTOHB7olCiYbbNZpEZb90fBjWDWlyip
1XC4Yd5ebzMPpapV/9rwGhxOsmi8hc880GFdIa17BmKLONzWqMkYXh9sm4SXgTAm
M+3t/Yl3TxhoTFrp8jIu0Vl2JgYktFfgiC61/obWp8W1ru79uFM2aa3XhPuv89X/
yhWSTyM0pkjDIUgIX9ej1NoUuU2wsTqkrxZRzcU92cinoTf6h100HZxD3ei9lT5G
kJs303MTeV6h81YfIpNm3d2VfjPmPHLKGSsAcidFTfAq++sQtdytTj0EmJeLjK1M
r/CL9oLo151SCu7VtjTs06O1JuKOA3KR4vm4g72eDeYJk3pPjU68sovUqfRC1Aur
IPx56vRc88+geQi/y3zC4bd2LTOOC4Rcxeyin0T+yxyY3pjbzlqHPK+oWE4WHEFK
KmKib/7WKDb+xah5uhzpeKXl1IW1e7uB/7sOshDFVhZM1Qobulm1t3WnpjJicPzk
Yca2WT6z3FNpBeD5ibWA6LDAKZAJzOX7VR0P5p9QC048oIuH/ZRPXKaQx7NmYa7m
+XG+7Sik0fsC/vLpVbrpdRpNCbQbgudr5dZ6JGSzMUBeo6pPgtB/AS+gwregBrIN
LZqBxL2OCvSUKovMTmZIxN3jyony3zzHgre2RGzzgpCQtPQRinM8Hzp6QG9Oe8tu
BdRCCTWlcl61A1jPqlq90qgf6K9fW60BAdn6Qb2GAd4srU04a9tPczMVszguc4WD
fnKLkUUiaYX8j3Uv8hrk+o5IuzL1jd57mBkr6C9pykgQUe7tIIMpUxRj62zlkZxb
LQ+q4QwU2aPgUe1N9Xnie6+WYjefo9sd+nBoIcuBnsWxbsgt+uyGsmX2tsB/bIFU
oM/FUdjXgbEORbvOdKcWnGMJAupv0cohE98QKgu7BdHkIbrsbXDc/soYZhzh9GBO
Y2lpupMvxzKbrjsSAbzfAeO+nCPqC9rVfu+4otJoCTczcHaeg6lTpYfYIkbskVfM
vLgqUet3dpO7q1sKX+/HMqmqCxedcCbU0ZMxxSUYUjYvi+YchKu3em750IL6jfdR
qw24naVjOKc3FqVL+X9GMOonmMs9Z4uRRwoIt2yijWnCnv82pKc0Ryc4RDVrNcDJ
7KlFQaSFk43Y3utLVhmpPsRAuy87thQgPLJzD34K/+IWuVL++rMALvNWCJLKaS1k
erMDR4PuarM3sqO4KYhCbMnmyP4fuW3yeWTtpABc5AsAqP8FuwrO+FKBfqnB0GHv
C8nzqJ6aX5nG64TDIXPqtdrLxqf/tOPj9ANvgzcQ1GJxxUv/tnissxlo2kvWwNQF
PvzMth8Mk+NPIIZleQmK3vuwEpFqUTZq7/m5r2vpztJi70LBo6cefsBsrPNLnV6w
l+cKkhuOsX7i4juHLFePokqdn51J2WwNsHbh3llHjrY0fZTzWmFmkH6ygdRmWXJ7
HipHewfOO7FHpKiOfmCKy4LkWUfXlalMbG2mloed81prvZrnPb/8BcrxUPxrt3GS
6Qc6vg4z0yaMrC3sxSitoyRBgyDSRJ78iAx/KXQf9qA1fBnpzqva0aIFkNM+rPip
+m3JEtILuGlS47nXSiBTlLjqNxHg9ZzZJYGK+achaEE/QiIJFsq1rjjSFJrXYh1d
zcUru58TQIJtCLBPMBHgul0iJy6z4TT2uk/rX9FMIDRbjHrRzw2YaOhcIJwlvY/n
MrPFOADHMzqV4DaSIr4vPKiQZ7vRU3eoS4cPD/AJT7MRZFb7kprIRkYMfMRrAZUr
IfIi6DOJ7Eyh459rLFvsCHLbnTVZa3bxmX/WVAr/67IBITJkUG6JFmi8wAHpp0QJ
wGwPvIC+99WsNhB7oSONUIdfon1DK+57lht9cIswOmGQbdykli9z7REx2fboL1Ir
v9AcuagdO0QT+unsLlaaxrOgF3E5CuxboP+trPC2lFLuy49zAH4pNVIzcs7REDzP
zYJbEEbum1znPZm1rtKQW2Lc5i7njd5/sWDw3cumfgpbVOjD1gsAWf5Vyfl4EDQK
AJ+VyMhGp8e++gxcqoxHNaxiUbcTgkF3i84yuRO4vFb3XRWgSAHl3zEpfcSMau/4
s7ovPWOyo6ESeyBXR/98keWMEm2XL8ZG318WdN6CGOvr2Gpzg1I77GpXJxE5tPmj
KIIYCKPn5FuUq7TSfvSLuikkDesPjqMenxPU8q9IU/AkTRetQfgmu6ZaUSWgGrP/
yJZfhtigY/nMaKTFcwKpcldtcjostDVP3LtgRTofVSICOjZKdw4dVB9G4h1WEQOV
qMzLKzyzAXYBQGbB/ElRSXRz6TDx5LgA5U5/SaOM8G9LE3CYqQAlHzniJCnRVT0A
4rAgFKTGZv20OK5GDUuLqb/vefK8EOyP2Fea+MPwPf11Nr2zhspCRVFUiTDhhxa6
lDPcclDtPDd5k/8o5swwgIneGQpK+giSCjs9DgbznjgHSn1QbchQmea1jCG0I2oz
qxwNc8/rCYhDFn+3eSEryISW7TGQr7F+LE676NlrQqIEmmhoIwQcIlo3ZPUKh/5R
ZOynZ8wuz8kLrGNUYEOjjHO3B99eGJrS5pp9hWxDGA9qoezRJvS/b+qLQacAmwER
w+KH5+zk0B3d1g5OAQBBCqQr7YtAUGHkxgEUaIEzoTQNq0gNvO8pFMeTCi/jpN8a
TuGErWldcdeSihSkTVUUP0iPvPHrykE2Mi9QmQz44nRwSv9nuPRHiFCCxNAAZJQl
IVZYqxnbRMQpsMyWGXgvnTFSY6JCy10EUeRNu/1qapYP5K5HxciHAkU/uefJbHVC
ngyGute99TPo9gSbrsj5EPfzdjKf6mYCBkKCF9Su2kuheycWxlF5cfR0HDhQ3E8q
g3YTkFY2Olj1SrI7sruG6dImv27B8APQ9seXHYhRAkntYzpElLbk3B1HX8v1u8Km
XPqJHBkJz+CxFQ5ZePwBe0hpF0ssDYaET4sN7A/xABTL/rvBp5FZJI8snKht2N6x
Kv0aaSrEnTdxYlL/c0HieBWwCibzgGoDLMTZww/kpo4d5LvLnPIeIo7OBtmIJpBT
IecJoUK/rYIM6hZOk5rO/9bbJaqCR3M5HILuqGdLhsJa6PavNHtrzYtBSJoXfDCu
SjC31KR6jmB1Nm/31K1EhErWC70My9WEbl7rXYZj5ymKd2a/81XPvQjOrlyd8Aj0
4tJsQHNXuoHMvYK53ABRyN1QPRvj5UbWVuxiUP/eOpUOEgnpNkSy9qRvQGyfTj4Z
92/vBSIW5mF8AMWijyVADxv4MceOPaW2OpGyPHM0ThOew+HvMjeZtTrtqNR7kIvx
eRCtKJ6Q9+rmdkNZQ79XVMmVoG/Zxu0THcQwlkZqnoLzI9SoumK7S8+9vgcqzgrz
2wMA2E02mwCMFED3PlTgGPZSiBkfk19/1mf7rgzBR1KKdRREqzhuBPHnRpl3WO3Z
3MHeciBjs6y4h7sro4vk4HplgPVLOQFLwYCAeKdTt5kumD2Jvx8RVe9ntFx26dVs
YjPm0enV9EuCnNcXEvMQ/2eQ0PuJM4brcjE/4zJ2fXHFKqHT2suA0Ioa8doRxz0Z
xrbC26iFxJIE4hRDW2BvV1LSlgHm7AW0KlRIob3U6gliGriH9zqAl41ujOtRY1XY
nsh3C4GV5QrCc77Czw4PicZnZWp6ms71YMgVf8mkraeEg0boFjAdvXHJ+XTOJwnJ
3kt6hjWiv081ZU7IpkJAzeMw+EQH3SJiRuxnWgtvxeifEUq3a/fKryhAjjFYWBbd
/C9NmK7n0h2ZVxPWgrKGfifv69CITWaLCu1QP/yQ/Zc4KjXE8fdp0tK5gsb1XI7i
/s9tScMrizOmZqk3KZ9DzunETp/VXqTqIE50GxkJUnKfOpRhAItWJFocWpFy8/Jb
J0gV7IPyHRzkRjtduysQJ8YGexvQwIxMYI+aBZx4Bmq8g5W+oNowpU6KarohFXBH
QVE/F+ezqBamghJCuDO/mdwxs/nUkzyK2+chqksryFyQZ3CaZR+/jU6hbO7sZq1l
TNmjsdjFVFMRUKPZnaGJikhu+lGLd0XK/G2w7TCwf1hCm5qmajH0Komt1r1r1fyG
vS5NPZpWYYxrZP4Uxk7j6zwaUQ9WTC6O+W3SFJ9J4gE+xZqTAvlVYkn5AQ5qkn0p
xMtdmay+Pi04jWyVljdthUc+/YPAOHoRVFomO3mmeOlpUHYSgMNy7XOxezpDF7xA
I8DFVle1jsRO/F6jdSjr9BzlGjLyPDjzgoPg4KB11ctcTrnqEMHza6qMSqts2qsd
zXeXi0iLgD0m9iBzhMr10YaFI/hbg9xHZkkk0lLQkEIiRS03B8RouKmVNJkwxFA9
ClFK+YV6bFKmC66kRu1MPR3LkszG2Jgw1NvHSuMT4SC5DI4QKmz54Kjy8ZF1Nxan
+l147rzXukssCHUOPyhdohvt7L5jZQKBBEr8/1IlLhvNOLC6yivtjkYXVc+MQIHx
dYzH2ZAyy62lOvmMEOURG4+7rPaCupqo7Fl61evZUO01QW575jAVn/waifWpZyqH
x9OsaZYqhDCFP271Nll32iRXXwmEry/l2kYhJaU0C3mwaWbT1swGMecBvPUZuOO5
OemqoVvgOrFLQOn0cPfr4R8Qgha7plbpL64rSsyceWe/c8DN05rtUZnBuFrVWThu
9jXp9IF+tJTjPtnX/MZicejQ/HFn461sh1Rb2hxZ/lskhY2OtxslF2MMSt+YcOJv
VlGp1FFV7Q4Bu++oKAXSHpuQ1hUHxdHAmObXV5lWiNBjewhzyt6+nmz3u//o1eHh
PjtoHsVEraEgAE7LVgVGTNiOldLKPxaa2Ni/2Fc7cG0eH/FmWf3axrkyNx1PTTEF
cvokr5+1ndXlnDtk38SUuZe4aFaniKsPQmuo38jppo7gTOc3Iuru0S/q3GqML2Je
+Aj8D2ayEDAdPFI8UZhkkMiHgvczQP8ryGftLzQ0vFjqxzxFOEnaHpPsWqvKzVHK
2D7wT8WmLgFmupf5pJDN68J9Y0e91E28yPGmUYABUlSyjBEPWcOI4R757Pz3xBXD
IqT6wSFy1MRVS43yEq0siS/nZv61kgDBkkF19Uss4USbFBW1KDeTQlj+FZTvyoJu
4+wTCx/S0SAt0LKqt8/sOwowiRvhrblkmkPVEwj/QO9d+COB9d3kkxVrWn7E6IyZ
Q+ELBBSFoCpISlAz3ACjQkX5usdzsmO+xMy6Ol5H0V43StL2ZwoAoDoIA6NCTL8o
REpu9To7h/SfZua0HNes1D84Bw/4FblinunnVXQoKq9zCheGSqDVsnrlG9tn1i/O
nfh33kBzer3gYcch+aa7u9EqlGCya7eK+wyicXmFumhdZC+ouxNKJXNDspUxPoM+
p8sV8CUNJWnkY6RxRlOc5tuDtomVqqeDV60CC7vUT9FRpjVMMYKyNGBlsieLyORK
qKvnwZljJFzzby+InFv8oeJ+ix6X3CU4kgUVQOk/r75PNOlRtfHXv4rpQSPZrFeo
vyyo6254EN2Qh2j63iVQGpBDt3mlYSyjoJGujw8A+EHGVKKPnbFm5mTVUwwlw5YA
7ao5vknIWHKua0OiMx5Dn8KDAM38b1v6fpgF98V5vmHQwPE/Hzthyv/3Pe+n/eNs
kEhhpSHCPYciffAyYGjk6Pv33pL3dd1tiFz+zo3+7PhGzFl9b19nloaJNWtgJWpM
plLcsmzgwkZ+zJA6lFQNK6epSmlLFVdNPukwqiu38B7MgbY0sNpnSmue6SLaGWKM
/Q23UbLiA5OWpq3B9yhoMpWOE+bsWSLmGsdPu/qsJivYJeBKGUD2P9q7eo35Ymr6
WnL0r1uLzK4NXBK/eBX/U3pyilaq4BRchQxXot8OWppjTkf8mj9OVKmo2vt00uc9
goWghez5OiuMokRu+0PfZxRthexqtBT88TUIgqj17Auw2hQFDSpaJP5UyrAm7bDN
TQfcT4cwaQErOJ3QP9Yc+ZWFkBQkruZxIgpSJUm1dTWzXe5LWIUHI3sL21nb747H
ef8wp90xnXeZI6R1nN7z63R+sOxlmFwJkI9lSH37AOrZfbQVrXUPrVy5Y7LQ9b6e
hjeRF2ozsGUTyhNIRiHEupAj4S63PP7WSOc2R2aiQoMXmZsUzyDM8/eeP6RGGwsx
ri9sAVWfqARRFtgZ1rps/d898WaDlgun59sbpqE5mr/SOhMmAaNcR70tLBNZVsG8
mE9Tpi0mpQNOlzYXIXYJEtUiQeOMX+cS2+/kkv08VW9+hsLEJKenhKzwYYDHq/3U
E/xjfVEafOB7tHx8dG5aCG7kIqmKsbhzA9TkKVjev2zCM0UxOjpqv1qUCN6VvWt0
NOSszisNarcrSIGSfpQ0PwOORaePVhBMI2PMb8UyLfyD+TdlGwOQSrTyno1JiBGO
pdbyWWaBRrRetHhCU1lMbeynq/dlI1QEQFc9JDEAPm22khE46J3N/6Mei2HdBsww
OwLFRjxartSiX33wxAf5SQWBGp9iuPtKnOyylwt1T0EtwavPoLFkYbXtZfRnMt1b
ynxnEV6HRGcGt1poKGggsLr9bButh5S0lj/fcsMOqeO5knTWn7o9d37m92qX6WiH
/sGOj8+9PAut35sPIy2o8IJnXrA1B4UhiYi/EODDsTr9BC+P03shalFwZZkUzUWq
XA2RA6tnTEcPzf3trIcmdvwmdyOQ9N0b3i1fVOHtJNSaYFQTq+St5PbNFTnVroJg
KGPV7pDLz8Nqh6Xs0BpY6XBqZ686yb1DnXoB0HG2oLs4SwEPQFbg8y1RomWwWolD
yRCWeh8KY/+9KZxP/asL5l454eEP7qK+HOn7UrHZpVgQp+dYrj9jw1JfA6Z6m2TC
f+/kNuhLTbR50FgfCWBL917Iv/AgZ012+zXd02ROG0Ljm3doZgCEem1E+loufUu3
h/RiYhrvjXdSRPOzOXBGo2zTo52PKkwVMWa1Zdn+tgJv2U/JuR2eNsMyrpJqr4u8
S14OXwjqwlQlL2XEzDW87cbklKzNXpsk8kAp8RRg+oV3vj6FGf3/WRWExnM6K5T+
48UpETlmX0+zIRYzZgdphXkyt3U6hjK8d5n4S4W5Xi7B2YTtTPJhaJuD85gmfwPo
O+HSHN9Lsrq6Qw+9z58xACO7PHpVf6WlBlwLAlXNE9SJNsR5ejgepMWtADRsyR3r
MCksnAjF6Z8ystB36lipOGLLWWEgHTdt9GSwT2J6CAuxsJNn5AQy+Vqu0lqJ9gGb
BTAY3nJ1z1stKAfmrRZik+Kasflyk1a13FFbpxzBXAhMiuevlTwHqIpYbZTvV4Zs
jxsQ9IQoUYRlhdFMjXN9Ktn4sussTXZvjLka4dGbN2kZ6567yjuegFAktSb04xbp
prU2YdRAylsLQi9uWj0JEdXp5Y9jPL8tOhvStZtP9Q6hehQlV1MrSLYvYgkiVOqf
vwQraxCy0uSSLsL4LgwZBf5qeFG8sE6yWCjGsWEd26g+JWVCTY3C6wLAgzcTfw5z
FhohpDbr5ANPRFj+W+FT8ESWE0eM6uYpax1sq3rldKH7j1bVzEolAC52sD+xCP7a
74AmQGzzP3J6KqA8rHj2L2/l2ZDriGx9umIvxgeGGFoyNdKbpVbzJj8GHn1B/XnN
gfFrkEYwTAjT+H3iRbq0IFU5OJKiXwbc2vVgN6oSFsRc+YyVjuNVxDOXcRI97ddk
mtXmxN1y2Ew7toyfdaTSL1wAfbrsQCOLjQQTh5uqVMgfp0qiasfNODTKPiRZSp0H
sfnD14aryj+5kd6r5uD7w/67EdeFUA/Au0sOEFy0TtmJfXbC2kcNwoqe1p88HX3s
IXj/GF0RrQfM2AzhCdJg3p1fEEHz7kKjudBQ+JKQRdhVd3Q0YfN5rubeiFLNxC3r
Kjs3hqF24rcPHg+gY10a7oGkl8UqL70raQKggSDUfpMJ2bOIuKEsETbPVPhv+nwl
oGkSzfpK/KrKBHiU8JLkIr0fdsn5OjwHHZ84AhuSgXdBFlBiYIRK39sd6zPYCloe
HBznRAco2+p1V5edOvi4ODUaARCp2r8XM/VG8+VnV1oGGzgjkb3IrWuLHQTlKQW0
YgXdV1igIgE6QtAf8dJ0wOBrlJrSfTgujza6eA6Osa67+n06lw0P+grX8t4KpdFh
9ke06DBy4DH03st1z3vV0eA1FnKcgFzmYGljo6UhTWYi+P1YqYtkLCSL6UC6YFKV
U3d//deBT+ou3ZW/7yu0Jsj0KhWAve9Co2A7jr0XCHretPPjZOQpxFVVQQYW/cgk
pc3gtHZip6kIzI157k1BbBX5x1i0QkVIm7l6vmG5GEnNS1xmHNvTjWRGiKgOg6Pc
qPswtUVWaZL6UvmmukGuCrRTnux3Wjd5RyQkBIy10KV7SxfRMba+7YANIrmHbvDq
KuFB5SZMNWELI7056wGxVlF2YRoZb1/kQCvqFlZuJwOLmsWMVpg2xPo80Xgva1/8
W52gdYup+f6UzBejetWqllP9MYg9f538sQYLVB+hshUjrPDXtgtcdKfL9LhL2gPs
ZWxtGFN6CkuneXVw7NolWEf4rDcw7qgZxmsELaIQGC2gWKnjlYmYn+XStxkD6rpT
gFw1H/2VDBqf2MIrf3R6+doI+ylI0zxS3zyPJaykhya0B6RYaEE87u+5tnG7z91z
yshR5LA+DnPfMGu9ZxSsrQKtdzi2hPmZDEGeURvdHd54DZ0NgVVF3TZDzl1A1qMp
mFwavYZqbS75EhDEaiVEofp8/XBIQyZFvja+gz1VlkV8GbTHBP3Arb6kiQbta+cB
ohvueCsBM/xXWCbfH89YeXsiMvz5TipHYzKWtJr5kxYSefzS4t+s4TvMYJIHw3mr
wudAE8nDUKO9HNbrXV4vE7f+OJQ0eTqMFdcB0VV/qko2gLawvbLUhUDVSKe9jV9c
cSXAJDv8EKbtukPLOq5sWoSshhmrNjPCafMhQpnqyrnKyRrjGWKaqlLB0SBFL07L
ed5rf3FlCZfO137sluB2v1l11TqKjq81UZy5vpumlfYBkvxfoBlLkskm4Itwwr0O
nToo93Z6fCPrXrCt4sjRFkUtH+LmSBxRFUrIVIIK7kQvAbavWqUQszlmr0KTc6Aj
xjtM9A1oi9GL8xfNWxldyJWd3d0MLZysc57bGIfMjQv1d3J5lchAgPYqxvV6aqex
QFlzMJONdEn7SNUTx5+K6f1lukeKbSq26+EscUSaGcLxi+o3ACWXj49aIGZIxaLm
csCCsDjs6e+mjbyVRYJ9ow==
`protect END_PROTECTED
