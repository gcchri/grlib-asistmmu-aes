`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+1w8W+nvup9/oW/8p07c+1oCE3r0IJCxr16cL0rt3Zd4Pt7oZC2t/v2Af07rq1ZX
AEnNTClY09AwmUGBalwKcsTM3DnKdfnA0OdYEWD0TuV731ujMHI6QsmLnVLnd8ew
mSD58zmrJn4DClCHHlAAablv4T6K7iJr/ds1imkyxA6jh7PQnBwNFii4RcFDaEas
HDQkYb2nEplZUwxs09/oAvRHISdr9BiUHpxHvrOBn/XIqAhZmw1fKXxvkqSHrSNR
eXpyRjyHT2esukNe1/JUA1GAyF6whN7w5WCVsM/ODxRIe4oh3cPetUe0ar0nCQFQ
24xOtnA6T6k3CpTt8TFjvA==
`protect END_PROTECTED
