`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BEyS1OSo+9tVAFHfpmaxWcM0X/KoYozRvlT+QathaPapbnlI1iz5xTYRNVQug0GG
ufaUkFOb9AKM+6w1aIQNWtASrWHnWEfA6sN8SXTEAqepn4dFBibs5je7pWTd9H/4
I+wsgJzqiUFBdXwisvbCN2oESxEHbQC9YtsHDCNQhBuvXXRaTB9QUSeJUr9eQ8Ti
2UZNcylCAllChqGQh9p56cy6VL3KFAQ3M9e1XoZy9fP6FdCTe5rpa3NxrqRYjvMk
ebj08MkAmaCb0qGyLHIgfjTQDnlmi+ZNecgQLujynkFGX2MP9rzQo4TVEAY6ekHd
eDfcJLAnLzaBMX5yQhroWr4tF8tX1u0yeDNGUaL8l5J6zJEtSxWyjqeeWkaUGT2o
lYVnQAw1KkBgN4whETbE3+b9T+NqBkPydpsX9fiiJOo2rG4SWfLB6KLPI7hvzQlB
cj17Z83VQ/6yNc6QKgWWCkjKcsNtZLgEJX/ZSee408ji4CmAMe7F1ahS6VdCLGdV
AhwAwYRJKDJdAA1WYx3yMX4Sd2x0WiVTWhaF3y+qu2eMIlPju8P3IsFmDkZ0LpO6
cczRogov5ART+f8bUnDQeQqfNsd3as6Uvl4EBLRAbfIV7Uq6882r9LtLS8LSmPRR
`protect END_PROTECTED
