`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NIKF11xoal7eIOsSUJbxtWSLcbJmIxctuAyQD+7l87R82t/TuN2NBctKHlHDhiTA
x1MRpXwFcDTjA7ftuMrfttqoqrH4gYCwcm04tJhe0HCsCa8zddIodv5UEf2bNQTR
tog6if3so22IAGUw+H4ksaDG5hYqsDOgYs9J3q8i806ZkMVaoLZBqrqTQc6a4wwQ
qrlbSX+i9uJm0B9OeBIwycQqolkWGaHzjUXyq9lrTdkzZRSVzFUb3bzgZUoJeqvS
tR3IS3j36ZVtkSHi0yQIT+i2+sSl9HC/CyDvrnQoxJhdGbblwPmY2Ks/IDOXNXVP
KdGX2YkM26zTsbolbPsyKB9PqH3hANLkqErtj1wdCmj8a4XQir6Vdvp/jqigX9b9
HRfnAzMbVoAo90KKTuAdJnQ3+T/Mg3Q3ny6oQtasdVdWmE3F9buc7XdIHd19XC8p
Hqr7UpjJbUuw+/rpOnBfRe2POsVChL+rEmUVQI0xrU2RQtQRy7Z7HlctZ/invoqF
Fd/flVhDi7D+V2cJR53sL/dViWCweZ5hCNrlfF52u/vDT6uBDqCH50JkuV0JZ0S7
KxvWmNoh/EkaMAL1LgBm5aFuzF0joEAFkTJxpBJ1AEBZbhT7lgk9S1sAQs/BQdRW
gy0nqeu6be6HFFBJqAwoc4YkFaEmsP46cPF7GKXSQLQ1G30MvJ2KA3dBDpRHS6Qx
aOkgcGc1q57dhQKfcOu107q5f4HtM51IuFZ0MsbFr5VKe+YBeMw1GsayEtOFUy5m
HzRmg6IfchAieRPo9/5ndrCOTjxiINdqIrj3r9AA6pjldNh5JmHR4teKMSY8Fnmi
dkSK+AeqB9FkQNNtn9x4CykGV3zTBIKCBRNtUjNgZ5GNAdyI9/xGd+u10L8ETTOn
UIlMwybAogqrRYMMNhC6l1DaLhplFiGj9E/rC7pvfAA=
`protect END_PROTECTED
