`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DpGVm9ympjDEK/0YYHPhN8bSD2LzABp7jh6I27D5obEnJCQQY+K362ykyenLO4Gf
NqbN6DnyroAi5f2XUaoz6ngYitKH6OaIqOgpsLxZl5Pg2Qygg4o7jmnNbZZ0MrMf
zKo1N1XnGPHjwiYHYxRMnCAVqqt2wbXSTXUScpv8Wxz/AiTgaoVAjmyZDqE4zpAy
3UvuutkTPWl8VU51f01GJ1X2fd4dqEMxAI2Ypvksnnbcz4UR4Sycuz0p9MEnDv1W
n8/oSvYlMh8Uavx3/2/fzSNS/tJYc8AmC1s2COy6p6Dv9bZoRYpXFDd0vc36F6vp
4uxqcOXH/blmiYr3onYhVMI7fwK2e28DdvopRlTaNiyzyWwWITz1ONrDJ6pWrZ/b
siKMNvOY/4H+fmMJl5yuqQ==
`protect END_PROTECTED
