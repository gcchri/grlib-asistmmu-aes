`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aKWnL2HcwhzrT3C90ZFCgWEOv/F8/tYQr/mGnfvddPGM35FxK1E26mER0A4rm7PG
r24wk52WjquOov4y+SORqZMkWI7BNjWGG5+YzB9Ej1h7V44n3JhSaQN9+B5AJq33
NhQmhz21jNG8U7u2nUDSFx7hLe7bQs/P9dcSoNyq+ZZB+YmWsedzzHbeUWAQGKqZ
QKQGB/fi9AMOhJTCWXutrS97XHVG3IXMVsHmSfynQZr9PuWekgnmx00XH1UmJ8LN
VaDYxEMMgQew7TGom+dAvMSqyUO2gZHm2WPrCcId5oDjaIBOQCfI56Sf3b/HX2j5
vIfDwCkKqYE1FcgwpagwwaH9vT6EVR/g+761AREefyXdmoQgYiHca0oI0F+VDhiR
wHXIuwb8I6y888UmhqbN3UvPRT0nHzQ5kVsjwhhkiZz/ePLfdiV7xsoa6MCEHMl7
xuIrozgm4vntnTxsa/BYAm1ujbY/NRl4X+E7hQpIF3s/MTjqXlAtiMtxp2uWoURv
FteT43v63NerIRtebpsxVpkdf2vhwEtvAieTkeau5/jjMF+sfn472s9ef4bMk5ne
2QGzcH8r9r6wldDoo+b1A7ht0N9Av1WYokgizat2U8POu68Jx/TaRXG7uYnzZlGx
tn3B5XeZngfJbXbqYrM7ElYaMXBvidd1uZrw3FLupVxckSS1QsB+ltMDrhwoKOR5
a2ESPaH48u1Q2mEBXIM4s15e8S7eIUKvjdFKai86C+HbCvX8krQ2/QwJh8AZZDNd
azgeqbcFJ+8hs869HexTtolV3LZTHFRE7s7wk6TZBvCFZdCUqe/Dww9DHG5snt74
txJ8kd1owtPEDGVahb22J6vDkFnxvRyJ+FmeIxK7ap2kd9gk9B/AzxtOvOQyXuD5
6EvVhK1HyUbTY6Ph2jQrWO3MVHNzbb2TqiGFzD2QFIwxjoJqnMlTe0llcxEC7GrJ
`protect END_PROTECTED
