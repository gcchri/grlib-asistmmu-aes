`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GRXe00VhBJt4hRxN16r21kfbS3nRpSjb8+YNA8ke3TwJq13BtIhFMIJDATJyMQaI
K57xtW3nHLLmXRbb7Gm/agMjDUzXOotAPJxcrHck0yX3FTCTEaOS2pfwwJu7CA4C
wk9wXUQEPtLZnotZ62NePQOW+Iuuw57JZBQIrfJbml8VeRbdf8EoEK9wLfMsY/q9
GGArANEuOS3I87BDOfW2NkIUWzYHtXPcGUrVdzwBzPv+u7o7zEzp4iEGsR/qu+l1
fczwxiWjVCRO1vSfGJYb7htlwhKG+m+Et7MawC4XRvU=
`protect END_PROTECTED
