`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
neMP5FleDDTFrbjRJ1BJRRK7bNOP5iUDt6S3V6KLb2vQN3jABonXg3PkwAQEBa3W
Nzv70q+S0vTxDRP33c1B+pBx5WABK7WbcN/VxNm4mYEacmb9zNptOgRAl/OE96WM
+X4vrCzJ+Czn7wODZTQl3Xkj4R7QGwKTFgwvlJSGWz7mOO9cRgDscNxY+vWCN7ol
nkhh1BVYKOg6rpaAp2mnHY55wsDfmCqYR7IAJeFjlIYsmbqTmRa2fTq+ECcuyHpb
JNJ46IlnmH2T2Gg4mbFqKEzM3jbJPf3UP9IgpEMcOpZELyAvDO2CreLwur/bQLJm
eF9QapYjGYpHMeJ/grcjue2agJ4GMsloLZiOD4BspMsI+YZbXn5PU93/F6iO3ILt
esvwM/64PEqCpCK8Iz8XlGuFTGqTqd7AM11Qa/hdMExX080NmGUEm506WBnEUfWK
y93SuvBYo58K6qzfAMVSQnPtWk5izEPFPslap5sIsAeEZ+M04Kwf7eevAhuasCIY
CLGdsTpaglcmSdhXphaHtSbeJoXu+TjlX0pwpWRIlk2dj1Y2H0BHPv7FaA6/CBj4
n/FTyk3k5PImCo8Lgn7H0KzebmqVE6AUMVa3oVDI1F5U/1pFYyK4WTUBBHO/BSzf
avyr8ipeyorqwL9lCmDXrmcv9NNKji3Ha9FgHvK0mkRHSWQ2ArQoedqZ9ZaundFQ
76ixcNheqsWK/a/LaWgw89yXgoesDqr8EPt3eyysY+U=
`protect END_PROTECTED
