`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Eb630TGjyM+CGgmLc6TWu/j9j/M9HSAHBAyMNNT7f4fnhq1d6XavziRujf1qk4IJ
1uLFbvut3DsVj5U7776/8gUBbITA8Ntiwak5ZEmViSglfWliE8mHd2Kp9j7BUIvc
2C+efeavHZ5n2neHqIli6vHqG5QR82I0+ZWi5IbZTk3FaiX0/ndoKCC7ytRNZcP1
6uJ7ygX3mE2NRHTVoRLGGtY2Oi7h8SNrBb6+NNS4+rVQ2WmSbjXSlAzpMWfWZp8+
Vqz8OGooi7tslBqrLoKkFAx4WWUrBKmY35BZaol1QpeEdCoAk24KyYVbvA7MPRdF
vRUFlutlTFIY9yrItRwOreZiPrKMcCSdCzDNMvQu399JjdJsO20PX2CYjI6rrH4T
g12p2BZ89CR8YM7t2Urk5/kUyn1BFmOZQ4/TVZ9jcSpUosoTSZSn1NrOkH8KDT6D
biMbkhupdyYKdSMileFyZGbW3ErYymDbX24l1Ib66bjorEUxZNB8mU8Unv4iaxh3
FkhpWEnsXxVLjzfZWudG7qCv1gpoS7IGNYCymw35BzMzhREH1nSASrZmpqDpRqUn
ehPyL/JrVg2ZdLkhHNoycKZYoMvSyC8ueqhq1ne0quAQ5XjqfQ2lzkPsweJHnmxL
U2+cmn5NIasU365LnIZzOw6tdx/XWYjn0gkmySQSch2s+HZR8gLQES1L01LKS3RW
C6KTtnXP9Utuvaa9fMFXdW0j6C2koP29Hg/Mm/Vnb/fAkOXJpkti6TkyyIkT4qZE
VxvFo+I2htjNvpUu2vFhdev7/eMEgkex+euUch/JFvOrTuyMDizOU/hvJP+OuzMy
oaYpWFAVIoRpKWqWUxFYzNeV+/AFdG70AvQlq/FU6rPjVsv5hrio7UYw/5g9OZKH
03h2RW4EttiE3Y7LeUNGIQcBKNU77I1OVyzZDedunAxypAswTCIoeK4zwR/d9J4g
YmDTLq6v4NXnF+8NZnh3dG+584EmWMlZNfwYriCjaQFV6hQisst3e8bGSpF8sv4N
`protect END_PROTECTED
