`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yPMVna7lHwb16HdAUx1GQ63dDnyh7twSfVwWu48dDkKssl4Ot7leB74Feflltl08
IKesrly4qZbgnJ7TAeI4ryaIija9m8+b1tyIc+/Iv8T3hkkC26io08QWNcGWmHl4
onOY145oDdEYl68qxRxwT+mqXeVtKwiLwq+Qpv13REB+nhg4AcA2UK2I/2q5mLrn
/MQWTySJUODeq7TDKvvyQ6auou7gVs3TzOejmYGsHGlsb9+s7H14giV2alYTWo7l
mvEXRM1heVAwjW3r63uGLAngPqghPigwDUmlKt7JfvLF+7caZLF3KXajnXyG36b+
qa/FjuNBDKjZ9njBuk5ppBKfXT4Wv1O2JEv+6RnjAJjlJBpGZ5kwNJrJiojreHyE
2QL+jflHWk/ggbChi3EPv+CAWIAShwsVDLS5UlgbRYbRfwtcn0liC20eryejdTXs
l4Bx5OJs/qb6W1FXKQsx3Ei7URkNtZ/TW8qm56KVw1NJUhQKJSMfaDxdOItx72W+
XEsohLTwQ9LUe1WTHVszUAv1xF7V9eUy3wyIJUe67W3morlMyV3dhDDaErPlllhk
SJL25tSiPW6mpqD/IH+VZNS9Ym1lozxHTZAjytSHSJPqvolFLT/Y4BLcnuwqdjui
`protect END_PROTECTED
