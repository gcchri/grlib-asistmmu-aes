`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jb1ZRKX+DZllqYbCKgZNXeUSRCDQRbHzpMwVXKL0izSkvmSDuJO3LX2PbWe2cFvv
nAeFmIZ35BLufHkWyYyEtlF01u7e+j2jrMG/gbClwf3x5Kr2+iBKgjkB+Kd9QH1n
lN04m6kZnhSDK4Xltzif1//Wv/221n3H8x8k59qA7YVj3Ty15lKWH4wRUZq1dzF1
2Hov9xl9J+OweIKPtKfpN5PlCzctpESU551INg3ZRwt7JH/ALcHbQbVncDN7Xgpr
lzn+tPCbLSfgDFXi0l1BLQ==
`protect END_PROTECTED
