`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KJ8SmNeAq2rdSygtUozmHUyYPE009CsCpqvWlJjSNu2Btt7D0NesTE1RDW+gRaRW
lpyexQRvv69ZKLCl+dUX92ewOFdT1gtRNBmFPRhEeyKbwuhx7aTpcnTpnQ+4PhxR
ppdLDqkoJU1GUV/JrxlMKHtfd1IzxjcVD/Z/jxWyAID/545QdSOU2PH8AWdyEHv5
+wUeH9ktoAq9r7Jcje+gJgMzqmWRrsRb+lr4keTGPEfi+sBz2rmnamXGOTKrNQKs
27DuoXGo7/77R/C75WDdc9+d9sG1ucFc4PCK8D5QIY914JX4mUHy3np4cmoSsRZJ
xuZVntj8seL8vJOCcC7aLXTmSmUqTdWTYBRy/IgvYwI3qn43+NJsOniWKAspfZ0Z
jqKpjv70I30tCJYH9+cueND4o3D9bt1cAToe6lbFzirOt6m5L2dwEoP3006sxomJ
4/LHENWW49mVLYPz6eCUf5cKXWyToKiFtk3AvSJzNCi0KfmGFfJLe5eUW1EUjgzV
pYoqrwm19paeF84l6hG0MYW1RpseFCIOZ3AMctm2q54seBQtYE5PawZMkF5Ypn1E
s0A9HsCQiHYGfgRmbqvSoyoHxOulvh4Lq7mmpZtJ3jSfnHYp1I6WbLeQ6z/lk2nA
n/Re8qJH0Kb7HefPw7ioNptXk7mGC2va3bWk4D4twSC0Kqw0jXYUlwbA/06G1tkf
QCog1LPKbyYPf3Ru5JVSPDOf6lM9FLU0hduTWHBhONnpfAjS4lmXD3yfAXcucLjG
Zw5E6ZvG2Z7iDRJ8IwNT16gRyF0g5XpgTb2Qf2AezR0hkdCqfMRgdwBLaLS8pd8X
CWCXfaJfgKeFCf6aNG1oILvfnBVrItuH9e0zViPgfPVcVkRTJWg1rFIuUivIkSLl
+bHQbWdQQSJxjb8xJbxwgj075EZVWAmfuqpKRCupdt7abBzBOEMIrikBV7KlSvwL
`protect END_PROTECTED
