`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KNJJOjR8pPBD7gMfYuRMKh4khGCkoD9e3RSov4CMD1wTpBumID2rGtG2xnPzvPIb
AILmf94PIfB8aq0n8369A6Max8O2oHBli3EwV08BelOh8JFkV+dzEa+kBWu/voRm
zyZ2uvKiu0IpFKm8WG9/lNbJ+08qBbhNhq5ppQ3c+o4ZUEiSchq1ilTB2iMdzVLX
y2SX93jtkiBiIK2OjrldEt/Ab7s1GSSwHNJMdXDgaezAQ06uSs77kyapjYFynIFn
pt+NQmNE0Kg4cuRFtfpiOI/G+/oMpPiw/zrpxWjPCW2uAe+xivxEV8QDc++DbVOF
GObEeJGuYfuuLf4cg85TEavW4ZwjeHKCcNmoXrPXJam9WgJ4zyImtQKWjY5K3Pct
ymEW4w22ZUNOtCX0mi29klpib9mNdv+/MXJrsOHzK4A=
`protect END_PROTECTED
