`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pwPwRWxra+2rPvLljan4azvcwvjvREHChg76W8VVRki1FRPmOX4IxHEI3lxSE1R6
flnfqO2KuGwByIFBOVtrSh63BX/o/Il4Iz7wQLpkpkt43AjT+dfYF8sxwuyXVyEf
KCZ5+hh4Sv2sLLHMihnzSDMSLwcf8NstQl5Q0DZs51sNuhrKeluAYoIeURkayZAs
8BlyeH6A5ZLX5vnUm1GS351mcSUSROm7F0lYzIkOe0SZPNP204PabqnsAlh/Gojc
Z01vDPqSovv1sIW5+ZA/EQ6mujQKy6RoO+izdzlI3QRddmg5nOa/rqTX5KAqGbEW
1V75Nr6qCiOuYYJtEZ6WnpAZYUjZtvqDgEjtI5NgH6lmvFEIBlHYEyJAbgeOXnm0
cqueOEKR5iK28bsx4xXyf2iY0A6Y84uZzKX+lIDNvOL6pb7XICwJT+uNo4imS/+j
m/uLhKrW0RRa5ykjBpUQOpMJTk6a8G89anwaCoHnSsTvjWtQLZ+4rpi+TOXApCYV
kSvsQGPhc0+MLJaWWzZjlPRPG/iE/qG5vRwS9rK7YCxyzAjElqkli9kZornEdKkM
0GSvawxaAK3VX2fF1RBxSunWuF7zjNY+x8jcGBgclgdhhcvER7cb1Z7uVH9eRB9D
ZpvoNItkp08sTixD0I1tuziAnYoZKO50IYo5OXieYeEY8QJei6yRmxJC3W4rd2mr
wZOD4zsC2tBh/++n1yGtXaXjE1fUKRM4qyyHRrvgSdQ=
`protect END_PROTECTED
