`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AbbWekIc//8xp3rwT/92F77jx6uSRJLUqtrhqSAUxJHWroe33iaRtmbzuw/ex/SD
2kBlymydS/EKDqkVtL47Yy3HycSFv4F2eqZ6Y3hjRIjLnenWTFZgg5C14gVVDUoA
DaLdO65m/ZUWcO+iSn0O8Z7kuoM/eyQcewOmzunkk90WLsHaVCVycVGwpp70jFD7
sgOLsMNRiAcUkej7pVGawKR6TaOzRfTwOqhlhCNnOTjkguhRNNMFOh7mOEnRGBgm
u1yz199PaYtOF+TFr1l2a+Tcl09g4tW/5FIYafvv0Is3CVGkUMREoGuFi1rG6IgB
wli8fjfvPWetH4enNonGjw==
`protect END_PROTECTED
