`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nNcloW3zRfQ/eKXTxsolrifePQRhT6XWJkd61noj+Mv6v/k5oGD8dfTZNPRKvBCd
tDy0FwMdrY8D9wrV6T3RLG4YYd0ciRlPs10eUQHLofQYtsTZeeDrYYbyygGjMDxt
UTvkE5X/cpvlHMmNLycV+9IR3Zdc7jrrJQq6OXwO21aGMesuAYietFX/IOGORKes
kbDe+9mtmaa1DHxgyM/y6VQQoT7Z6h+dduk1FZpbckIy/i+PS2SLlOIZLiv4Zp/7
WT7bVxHFHIzrGsCabIvMGZdQ9tFuujfr+0saMFJfpaJknO1HQRIBq+JlaUSXUES9
189dOcCL1DfsUO63RAhKrwjYWShifIUh6k1voCY80d4I2aMLyzkHA9mUgWx2Chw9
bQgG1pQ17FEcjkOCMrHnUeqQweaa2l8IITCKfJALFds=
`protect END_PROTECTED
