`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
si8ILop7+JmgkQtUAXKovNZq7BsMhILVcOp5LKKVL/ZwEJ32spQfzxkhmhcaf+3o
5H6KgE1qdSOPARM9llkhcvTF1uBA89J47v1j7UoVssAs66H2Vd+y1GFe8UrNaVqV
r2QJbMQ/2m3H0vzS6AOuF2NCbgMwaYNUtB9WwriM3jrj5gf/PT5c8rkQbbJO9hnQ
QY3bzfeW8XaLccPexxxiwN91aVabzC2S9DI6p+78LDU5mbTBHvxsUptMhlHssypn
UFD7sMAiZbtSy1D+aRP1llpF8x23gKKJuolONxI0RkDRSPkfbjbYwcxH3EecaGGb
ch71rS4XwoIPkJ69PlHdsMSpqFlstPnIq5xAjlgNH8J3CRR4gkfmqzYTsB2cRIWc
6fSZXJrH1vAry73xmFEQu8FxQ2B/htPREp10BClvLn5nhUUgo/bq24FHwpmchG3l
FUhq2DcHZBzjXKXiECtck/w+rhI3sfVxEC8wp3aMWzO2LFgrTNHvEdx5IjqjIsFi
JgmwPAwOgU42AVrl8Qj/mP2NC7ZSkp7DfqxEWcbz7XuVVyzyUtynMxKGfeacXnyo
sujzhfNUA6J8hFPVyKIPMcLVGZJtJGhP0nRl/KtPOUG47HHUDZy6VXYmUxrLKs1b
W/xtb5B11nXclOPLr1EOvDnq4UhDjq18c9dy3sIvcBpQIhs0QzIj7KaeIhFJlF7y
`protect END_PROTECTED
