`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j9O2r0r9Mba8Yo4wWJx9hXDGHXV+s3FYKzrlrfpAZqvJYaBjEAYxrYGInc6YFHw9
PmyoyYi40z27T+Z2fvdW0zAt5zg9JY70JDVUjBwI1Zhzdt1Kmtwo3R0fEPTEgMtd
UB37s6oecYSYb9fZ6XlyP9e763vVlyJPGsPA6FCEyvBdyF+0LI2tYEDrA5IPi0xc
Ff4QHseVJf4vJkuHRAkxixZ8HMWwyF+UBiAlj6ngTx7IqLO70+2fr9rZS+lAB/CO
MjoH51HJYdvgfd0NpXcd3lRNrad4Gf9bmRquI6fMiNTaufCyfIDxF2T11Bhwehe1
eTc4GXtdI94WjkGQuJyTELHCQOw0udcs4xzki2ksDF4=
`protect END_PROTECTED
