`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jJwPUBRlfLS5qW1pRp4RmlX65KEc/+8ksjohdJS6NUSfMd+RtRDRO0n1VJYF7Xde
P1Y1e01Y9Q/P+pSClw+8MH6KoRxIIbY+DvZ8ja2z9hGWiYh/m22dGeG6ZeR6U6fA
+JlUbyHwD5ONj1lrQbMJgxCeb/OeAFSqRx6PXO5MfiQ38gKnFRa+hp2TDIFyOBNX
OJzQSpcI56iCWdEIe3m7OtUsEV2Kitg5w8SOlEGY+ylfgSwJNc9B+6btWZhq0I8f
WbUOXHJReWaltkjP8JUZERSL4p3Rf7inF5EMtNvOJxjZWrssFO/TSFcm+OeeH6Sl
iDMCW7lKATqHI9pkCN1Sh7/A5jfTCjjmWSvon0U/i4k=
`protect END_PROTECTED
