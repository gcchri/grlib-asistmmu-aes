`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VlKp67icVmyalcKUqKPOUltwOO8UN2JQZo3lf6fbxH0FEqzNYCDxYEzgrw1Ku2zj
lV5n6z8thKYQniFa7FFed5tXloeZKDWNwL3n4JsrwK2nQOaOGGkAg7If8uupvkVF
TQ2eSzp8RyM7imjladBFlBkHsNLojXAsddEsnbpw0lqJjGCUgkpHOM+gbFV4MQhZ
scZ3KRmg1JIAAAUaxwR6O5PRbaD+xfxUTKE5seXKGE1ucDTW+bC/CyeganCfecb6
`protect END_PROTECTED
