`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O+h3+Qo9lwplGN0/OQMs5pHiS+V2OeGQfkZQv11It7xlCOWtEXwivczke5cGymTX
YtWEiRp2Rg15pPbExy/7w6tPw3iX79F8SaKVZsiCQ+I2WTNg4ZYF3XmlobrptuqO
AP01UHXpA2o8ez5BI/jvl87b5zTZWH8neB2IlTKuWh6qLzLrIwou0EeZAvV4f7qQ
scpi1+5w/50qBVALcI7Z10IMtiiLCTZ8AfCsQj9wLINGHAt9VTtNr2pfgaGgTl7E
017O5hp54nElWJA8xet4MPLBfkcZnyA3GJxymYTkk0SuZryDMn9v1/C+C2lYq9uk
slgcjazxuj12W9LyrwhZdHhmGS58GcbSRSMC7lHiuPxrsFLwaQEUTliJ4AtejsY0
17zmkfpziIDVeylQbFydbzpXKKWwyG0jDk5J9RqbsKsrlokFeh6pXU4XVPAWEfB2
M1R95vHOniJRopTrrP8U262sp6sK7zPV+EObf4GrmJQUjeRdOYZLOVqf6VWaqgaW
DqhMr8yix5JXy5v59gPsgWzZGCVLeydfFajTLLV3Fn+eWoGufe4ITMR6eQdZlD5z
DWeL2yzDY7ERx+swwvnSY5pr5pEfJuy3H+wbhx2XhOA/i/3+dlbVX4N1mu88qaPA
x/y2G7kqRkxxyXJQSE5gqbZE+k9OCy4NteRCJ6xrcs5I9Cjb4eaSKru2qlFMbm3A
FGsw11Mb1jZGcAnHa6bii3T3rIiIBgvjFLeAGquGC6k=
`protect END_PROTECTED
