`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t58cnTUpPRdoSi9GtBy2+e9lAjjSoYXJSvLQ197KutZowTo5ZDMofd4fHqZ3xxAb
9sE5v8Mh+4caUGz5WmuLZFikzk3b8SYtV6UnZz/cdjHXMMgIn8Bhz1osPm/1a3WW
OH+v1EBYnqBOqUfgKNJ5RbtBPx5WpySs87baZFAyAHnYYtAFUG2umbHsTYtOXgy6
Mw/xknl6UC7G6Qa/YpSOBTSg/tTDRce/kd5J5MHJ5xSJ3g8XoMTAy9l8WOfAu13s
3rEDx8C1J8uy77K5QsHBZmL/vdvX7l+jRWhqDt9RdufG2Le5UAJGe/l5anf2Rx3k
uGFx7O85UxxWSHOljSmxNHsrYy7Cnkl5//I3I+c9lVvDxOrPrTqfdqjDBAVXGLZM
MiRZKp/V4BM+ZF8J0PnSqYkwYLT38KKzGHE/+Gr5C4LK1b9JjEz7y4bis53onDki
f7pQd04bk/nuZVu+/DywoSaoftqPAfymkg4LvEBPDUh2m6dbpqx6eBTjvjrl90oD
B7HPWO537ifnHc25kxV3AknrF7gTJ8ZIL5Vb1T6fDqiw26oE0bBjZx6ceLSH8VFF
TI77xYaIT3qQHgKAHn1na8Jx/S1hwOdrEedHtLCRsMw1m1SSyAtDMNuOWGx9GkAg
4bJCBekpmsKHDXp1hrLl6vk/Nt5Y/fWRGkR9avvDI8qDttWdtuUmmvZmh4jeW0sL
EMQBb3ulidxfvjwuMeFuCOLgTxB883KXSUGe6VvzcP8JQcON6Bx+yXBLo/TRw5W7
8hOuzLKnGABm5hux7pTXJMnT9voG2gNrZAT9CAa+WHSxEez8JHHKbPnAbU5kgXIk
+/1JkJ7YnYmZEgbkgJmWBdHgdnKQI9OM6hf1+HdDjlfLq2e1xO0xqwUKsqUsJtHX
BOw8yIfuMtq/PcsWLYJ+OtTwiyeKJ7omheesPrwVEFk3wOPdmE0/Tb2+bTb7+RgQ
F/y7tsH/bWzhRZhAv73zOvcz9mlBqntIT2BValmxyzBXPG16pUIgy7FvySdXmIbo
`protect END_PROTECTED
