`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yn8RSFpLGqRO5jIWRFwxnhnrnDAv/uqgXTJvQgjTMwcYpSOyRWuxAmCGzUHiRxzE
wONsnTjOiSx2LOMpEcPItXi17hEbCGVlsIjub7SagZw7qp5YjenOkXUfDK+zdbae
IAP7Hb/5PX/E5eCxk7NPrFoOFphauMpEXbrZINIkI8EONOjQJuJG4eLQXt/dzw36
hOnZ/v0gMFHMIuN5A3C8l0qj5LdkkUOMEIv+EJ1WVVrEgfi6RJGbiiWd3GBUhDKu
vhwgz+cSGvJBtAQvmi14yKWUrO0mIKjyrumFBCBGcoyHeEwSCGaEH+uEwPNFW3mQ
A8aX+EsLo+Koqm9kotGnu5gNEGPfU+7I3+pbpDdCZ5GxQNOyqYJerb50fJaEw62F
2xD9evQLqTWO4YlRA/8uWzbFMzK4U9cgpqDTkHCq2rxjLNIv6vxRadZNr7FKd90V
VKCpqkA0Lm89mO3AGfhIq4hAO2xYpKWHjgGD0bpMLbt5p8HPecNID9IK0GgSJHkH
uFzvoRgH/or8wN/Crj9zeJLMfTj79/0ylxfNZbPmk2GHBpWN4JyGxAZPcAuobtM2
uo/81NPA5nurKB5FLa3Fc2UgH0bLTTr/zKxu4ifU7dGBWi9XMlYk/MrxVGWzf3g2
sQ93wWFgxAoTsjZPWJlULsubS7GPpryyfCOu7moDsdA=
`protect END_PROTECTED
