`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MppYxXUGv3r8AI3dqFqqe2wwoUodPlPdtDkh1g/AaYmGRipCo6vtP0fYjwItU/sX
SRFhqjzQBqKoY04gQtHTZVc2C+BKqROW1W8ZPw3oOUIoEnS5G0L+BAEf56d6JWCS
yPOPAEkBA8e/C5pQiaGfpVG0kul1Ih8nl7MplFp21DWDmIbHtStsh5AHVrnAxJxi
F6TdufrTAHPVjVlqRmbGwlNwGRWRZLpNSq31ngK9WTpjr3xAWhh4Hjmh4A6jhlqp
JoTwlorGfpVhvugP7xitdJb3jvYKOdc1xevBBAYKNhve54g5zyHEvKv8fLYsrKk/
Y+zCBZsqtb1gulCozuzxgRG9mU2bYHHMWrGsBZ90Fs7sjUwLMy6lr6GZd+S/BXEZ
6AVU/YP7OdZjLIKu5w6Awn9axjIWGiK13N6UHjY58EJL52fuWT9tFaCV0/8WHDLb
h8JKtZcCbD2ehWdAmph+57YiuEZMZ2myC02qxS5l6CKiK8lbsLCyH4Lfta/gSmD4
nSm+EctmaLcCMl6/ScPCMUaVvyRwp2SnCzgJoIv+M/2oqT4XyEiKMD2fJ66tfncp
y5OKM53yf3KMrLNh5+4TXWb5m0NoLNd7cK04UTCF115iSBHCEgzuuzzO2ZTZjAEn
T3htGtlnHNYmufxSb0XLdKO5OOEMZTO52En7nkgSNVVg9KFENGir2yI/XkD5pPp6
yQHncyiQj5ciWnQY6Cjiwvq9A5y3vXY5L9gUlbcUvKh3hRPfn2A2iBhJIWIiHISg
ibFfv37/de9OhTc0knTn0POTs3BDRN+6+zo2aGeLVR2SWVGWfaWwwzzm2UkQjUVA
NI3pkts3PCdJA/IyV6BunTCQWeJ6pq7p2F9DhCnkCbIxfd5ShQ8RbRWdGnf+2dfh
QHKFvoxte72nyNKDKw6hbTyDf8YhvvMaC3ANeKjFW735GWqA4qHTRG7T1NLSxpB4
RtUQFgBZgwY6Zk6aORQTrLJSrgjtWKjCTihxmO/YlAqPmE5OTANHDQa9N89OBV5u
LSEiYW/kOoh05OE1HbC/L73/ZoW9hIqG9nEeti6unplotAeEgS+Mpo41D8a5ovbM
wjYcvyl4VE1b0dv8n1RB9a2GIQvv9sg/P5MmPNbj/YHq2RZbC6HULdvB5X2BC7KR
1ARJzI3CtvL6fK2zOzskCrZtqz7DPs/9YnY3luNG1d8DsEqKS62VJ/WGpH++uEyl
Wk5Di9LSFh5vK6VYUyEWlTJQOtzEleRMORWEkspAmgvWrx5hRvUh7/oTABjGTMgH
ysphfwNv9vWUErX5KDp2IIgGcw7t2Y8zWgW/AGxlgrWmstBNx3pspBwY+vVMVMZG
840GSoJaSXJ++a1crTPwuVnRdYZ9xSHf8jgGVmoRnWacOmfST4BJnya08jfoq8HF
RSnC06pmy0L3CmFIdkkO1Si3WYnfFsdHArtyN3cHtcD90SnDj8fN1fi+ZvCAJm3o
AP+BC9CS40VlbcJ6RvVw05NgilORcYcYbNY+dtAlcHcj8rAQcfpUZqCyDxJfUhRh
Ejopa/eKRzud+fzl1a1cmL5rgYMwa3joUlknAfLTuCoLjqYjrkQ6QOXBGdOIuakM
8JUMsXBlOyMkLLmK9G3nhlsWD7cK95Ngc1r4LevenAjJlOt1yT3sixM0nAADWRVg
pmRyIy0ThxNh+MmGoYPVWWV/o6JzDivbJdOgfa2EygXtA59cyJJ137DsgUrvH//B
Qwy4TwhA/PETdm3WE0QN+hRl66XdEUbD7tivZ4cwINBZ17zPa9aH7/TiqVYXrU6l
BmDtcmkJbq4F/yCg1EOrM/3+jRQUGJavkt1emXafFIZCVQU3eoZ1wMSHIcQi9D0o
gvJh+a+Ga1Lil8yF9e0hPt58xP0IJPgqL6R4xwCxhKMKmz/gctTW5wqp9XNzC11/
miRpdye1yhQE5g3UY9kmL+uV9fuH9P4ib74f0ddKqqCp3Edo2DTLvaFKclaMXpW2
5PPf7jIl3EPoBVa1UGLHJBPK4AfQ1LkMIVytSM2vxjQskcjA5ELzCY4BXpCnM2ZX
8BPOGj1Aqjt1mGk9RaxvKRKJkUVTGqrdCuSp8Hj+oqMiUjvQ4WVtDXDZpxObyvpk
L/KRe5R2kk1G/QNmiwrjFsr5BE9R7L0/jZZrfNCTyLqgUk+jpGatg4okIV9R7RY9
Yw3mcGmz+YsS5mu+gOfr3vyhS4Ohqk22dMOmTUbRsqRF4llPLrS7btiSz/kHZB2W
7lHYd5YvlC75l2/QF7j2+lkTLDaSMF1bg6TjGG85k1Qgr0uasatl1x4f/R/pvR1X
dftqU3jV+AUovoK+NYMbij/o0A3x+zd3xLsIoTJ+ZnHriNFODGYevXWDIoKV14y8
xrzPftXh8DaMNC42J+iMNaJGx77Uy124y+i0sOFQ5Ta8M/uyRiZAfqWKPgh0VKBR
gclOHDF7uGHYGN4yK8Htjc+kEyjRh4dKQwtKOd5PvgR0+7g79BsURHynVguNa7B+
4DwTjI0wkyCtGWm22ptqQMpjr5iOeMih2mvxCLsKZNLKEZZk2wNQz1KN64tx0Uwt
ce3g6XLI7vhrKPD/LcAHqCAD9POjGMf/oGnpVmlAvvxeO2sFSzH8P2PBOq19AOso
p1LQtuYw4DGh1pZ2LKneqNPmr/pfhmRuRIn9k2cOYrZl+sqbTATq2LkcZAWxlb40
74fxAA2eqlDjXhoZM8tmz1OdjBaITE8t0Ha9xzbacw5Nko9fqnqevC98gWVwUYoa
EZ1ZW61+rLKQl4MEIEI2HQG3uwaJA3mxjh2jMmN5sNJOlblb6XAYdQ6CRr+6Vkxp
N4BS5+o7dpfTDAF3rgKHn0Du8f/3DIdoEMIKgsgqz4NbhMvXDFtA20FfCQA4sYk1
6UfG//6VFoDgCIRq2gDePBYbhFv8j9BxxpgVx5w2nHt2W3Kf89oK81TvcHlMLX0x
QvF5NOP9gM88JzQnFDwgCgLcFl6kkQqcWOj+BIFq790s4hyerjdvJT4teL3xbPpo
p2kbX+4OvfnzgGb2jA0CfiDJv11qoRRdk9dARf0y8fJK15C0YGd8Vr8QNiTFNNi/
8WQL0OtuY6/iq6FvHoe9sABCxzEPKvJokDUynuBgwcXcg+in5aG3C1OqTB2KhFWq
4uIRQLlfuXycq17ULx1g9t0UDlwdKkXAdPBOgC+N2X/AEDi6XSIO1HPBMU3IU+ck
qlqx2vGJsJ9hEZ80SwLmnNTqsI7+iEj1QePhhiaylj2V2AkKndvzt6QkvHE0g8Wz
sxltBRPzFt5Srnc/uzRrCMpjQ8S37Nulv1WmTJ834s4WLxuueYb6/BO0vxCSydqH
AyjYn8FoTKeNuuCQqV1QLyu/iAuRrzclBN+TmSri2zlrsPwkT08nw4pbDI06oL4+
wXC5zUR5Y6196PpAHXCxANI7lp20guOjLrUO5wxfpl1FjRH3ohzVBCjkX7C66ZVo
80aCRoiMPSyj12pniRljCJ4QqEb+57fmdByU2K02q4354jYu7S+Cx3ommOiPLD8y
/kCV2a29VCxULaUdulopUb7fzbb8O2EG6devA2uXiscDIOmCL1HVt2fzYhhTBGzu
8GPSJ1MxpvN+T91l+iVI5lOGsK3SQv6DPd3aaSFvJiOIb7nhe96s70Ehv9LLE2S4
cd0TQx6h+r704/heXXcU6JQ3Wlc6z6pO2KvtBquEx8Q6cUUhQHblZH1YLh4tiCZG
/01VjcoYIfq7WglODoRv2UDo57UyQUXA0vTS4SrW/+VWkkjbTf5XabfqDvOJEC/o
RzZgPgFfQnMpRzk95z1ms2CKdR2m3FQcTNHKqjLTFmf/SIx802eVa7aMf6q8E7CJ
q32JZYS2r0FEZP3J6gaW3How1wVUWr9+98f9JGb8sioYR8e2x3wGHXSZtX5CC1y3
fVGasd63bzi8ndD3sGvvpt5hZ5J+SCdHH/BwZgz3O896ivwMh+CRmokcfbpPuCZF
hDwyePyELxbvm+6Z+zqqbrsbSJ3Y49wQk6hK56zdAMWx1Ml9YVYaKC2U2ClX8A2h
lNtH0YA5zlyMz6UY7Odn0Jjj9xQ6teShYsqQN4mAkoWDuG2SfiOS7XnUiooA6jKc
ZRyyyXZPEr5KScRCQoyBLyta9H5qXq7ecxtzewYLwKI0jJTHwYZoUcMP465M1XQ+
ld8G39YDYmFStfUrjTf72h+SiQLtTMER+wVJpBKzCdacDwtyELZReRioVNhUY2Kf
Y2dXGMv7/eiPn7O1O4HtnR8Tk3XokBl3wKT1AvPcf5x2+9IUkDRa/pJsb5Tg/tZN
CVFfpWchnShAUDuH1B2cNUV5SGqN9VgGhI/eTMHRMRLoii5LtitxFoSzZMtT/YaH
HzHYh7YStRmD1fh39YuT9AEdXdpVy6O5OlrTWzqDfTVZE2re4vwbeLviyS8HpjoL
dL5bm3ZghAc347DsS6fQAdHGwRT59PRtY4LLMY7lg7LggbJVK+X0nYSJ1lBrRjrj
s1/qz+S+OE9+ENEow11iHkprAvdPPDGW9AKUIOd6raTW3RJCwFp9Od6PVUwSfsMT
GMCUkLrGvpJHPj1C8HHK/2ACFjsUXa76HE828QGgFiLRVTUnrcnrXN6+OCwO9bf+
cipBRHqI8ewAVeJ1U+rLzjJ7HiDypPrJnCXhLl83fvaZx7x3BMnqATfzSUpR4OsY
o/aAyG45tS+vf3jQ35WFy8FBQFLnEyduxsa3YYkjWsB0EjAHQQ7l3v+gSvtJSaOI
ubJjhX0pVUEpE41oU/bGTxUm0b5nIonxVcOVV+D2nXBd9aeeTuRaBnLQ8aklF+ei
WbyZf1sVHudaH5bdUotpVV2wBeDkRsAB1ukfJj72cQ+PF2nnGsMRjP8jF9TebPw+
Pv/Tsu+dOc19i5s49NHcDwUwwA2ya3Obn5OqvRINVZw2/LELpJ4vdhFawUT479gn
7FnMk6fvPNNcFr+M5mhDjHSs6wkp1553LwJnu1ZMTD/cc16LCuLBq9IDdcs3wF7t
jWqDhX/A+4ujT4nwjOK7cnpS8sBFVnkI03vd8rMVJVYL92wLW18cOSt8KlaHGyF9
zVy6TqggixAaMg6B4eAt31WHwOCh2B2hebgXQ6LXsF9gO8uNlh5J89c34rCD0ekZ
4b3tHG76/lDDCJzQnCUbfyBWMddFsaRp9OdE1DjoEpA6ONkpZz1F6XQivh61eArG
u7wun+tAX1Q7sGLz/G1mUA8+GtlxEFwRsW9VhvQ6qyK77WhWyZA2rIR8bpJZD8ZS
axqWECmB12uEuxVm9mM3tIShp85p7ERd4Bc+tMoqMXhgkNh9xnpWxTXP0c+ocu/E
HHrl11AEEtbxdz+saoF4PUoSXERgSXdee1mpIMHzHOUNtW/VNbjH/Li84gmvYuw1
WyBaMm/nXgbOnueVrFQH5M/Zoj6Y6nEvgRQKzE5M/y53Jkd4PCZ4vXaoKruk0pdm
qeh/231Y5fr8jC3RDczdeFbplTDAPUpgxQWTuY+a4BQjjdfGnIXpMerAcJfwhsfe
zhA5uE+Zj+fX+5EcEmSxo54+OSa3V3B6Iw/7qBabsB70esz6y2fCppcK5A0GXqrj
qwPoT/cm4LWMEwLm+SPklZK8M3gk+Zw4R9N1xAxdyM+PEbf62+AnIp9pGBVk9fBG
dUfpxEZrmUip6uArTgk5oes2gsJGrFvVkR/L339EfdOV4xxINmdamfxkmNA3NI6d
OW0ICIzImtc7p6FYj7FQNMwQPNN8NFoi/nwbZRPIbPwc0nvwcURclu5Iv2h76Aqy
YzsE8vbgNiggizLBoREuEOHDlW2r3o7a2UVMvYhmDkqawEEeZNehi3wOtdUUfX+k
dLwfoEqrMXdJbMkKB2Ec138nCIBo2NiBqd/Ch3fzQ0OzjZEuJu912ibUqPPcIijm
RtVU2F5R+x6sQDo6t9lNr4i8ABkyjNORSbv5Z+Gfh1CSvFuFY+hlqJuo5ceSl+vE
Tw5yjkXyMB4gQDq/XgDd+iCinbud1M0ZNaGc6MDKx38iftu6lBp1oyUFJc8ZUTUs
jbhNdTOqa7ZcK1PL2eh0smhijOACPoKxeXqPFjG1BnoL6acYalwjPM0vqrRFNQ27
W4ReSegQzibldNnC99TxMiCFs01IK2hBsxJ/g2spSN97Y3/aiKguLB6e/qLXIpXN
+WrNXMxxtN7bsF4qkgrrtRRBISP2vjB5IOciY4fzEEWtyFkFE2d8X+f+VAO81Hhd
bW/4HJeNb8GECubFjwwhhYARLdAnuc58NVQY2ip7ZaND/0xLiVCmUoiDNlXHqisB
wQ/UMiqwyjF5Ngf3DX2ZejfKvUlz3yVjPja0lmTeMPtAzQHZDV0JMOIppcgjJ3/0
1Q8bhLvuslc9AM0jAmR4nxjoKQzp/v5VMIjS+PVxLNHCfTOatvbNfG1FrnNq3RRM
+KCqV0PXpD8mljaoc3k2bLZXOxRhoRw+qfjfuB5WyozTaejWhhpY1mrBIRPXoc0v
egeu3KZOE/HuRbo7eMWZTrhQ+L5WO97XDlt5P7CSem36RKzQbR8waTPAZFCOCQWV
VGRZk8sPX3QzqGTTJSCfGPef9F8hDsxlzYUAZ0+JUmtzMAx8EBbGpSa+6swRbsrl
pSJ3Kdh0/rGWqwY7xHCypfsWYyk4dLbB0PoKEXlZEhPtF+LDnqJQ4GU2aL/c5yJG
/TSpPsPAZ9ZaYHYrhKB06JCu0iCzxtc422Cy9WlIKcpGtW8CbJtKIVUqiMHvNib7
SHzO032MxazpzE6TkEP1xvLaomQX9MzO2Ns7e/6NIbjt4Vtf2sx7By1q9iEVlsZa
20HsuWyoq1ERgOIHgL0E8odWN1vgSdT7IJz0SJE34om+CU5D/YhxpnDVp9xr3wMx
jqtJaj1D8L6hDKPPskIAUiMKZDaSe6lfo6WCsMhrOOf61vD/0GZcSIgzHfCrG4sB
IsGI4Sld0UvrRHWMj1+rwp9ZyXL9i2LNlUBvT9s325OHNSZGXYi3CuLaUuJiDLc/
HY8NWdoR/z4zSihsklrjUJ31G5YiTyDashrkVi6e43E39qjsn3tzlfSst3zE6Ssu
o/l5oJlNfs99rEbgikjUIp2Oxk3GvSQb9uk+SJ4EJQljL98kxWr4yQKuuva8qFGW
KxuVr9/Gl0RQwZgW1lRB/LLUX+So85sYJBe79BrtSWZYW7YI5IxQaPbFXK1LJB4k
6XrXQNwrRISGnXvctixHTzgaN5lry7MI1FWm/zhbifBORN+6cHDQ3Z+QIXqIs0J5
D+/PNP0RjMhvOr6MWk4ezJg/zUeBA9PaKtofVoCYbwp3lbVcA2XNB+GHGfx0WhIO
PptTfDadwSAT+k4rBjnqZTIccK3flFzS0awAOFAic93c8w/vjX/JaxE/XYVutXba
jjiWdwWiJ7yhrJx0qiBjsS8FjAxwY85HexfoH+6afm94Nt8yGCqpb7pfm5efzUrT
h3PaqiJYSZDX1+c2c0Qw1n36KmHRGK7owNM41ZSDLaj3HGyO5PnrbjyC3Naxpu/j
NX6/aQufj9AhCU5//wn125S5CwL7nR22OhbeuTIK6MZoH+EZhtYcfOKmZmCn46tO
QAkA3OdzSo41+yjl0IvPL8Jd98Iay/eFWk6PVw56Bw0Mu4RifnIyURF9iFR5jR/7
FpzZbGFT/DH/8Razl0W9fSTSGRfTurD2YQT6YMIytNw2CcdVerezis578SJzX/cO
NHTiK3txxR0+zPwE/bCSUDa8EOjOUjomrvKmyFaN+p/fR4o3B+uyvS3iUQ2jVImg
sDwTEzPyobdKhdHtdwNx2ff2tPdiMnq6IOl8+Wx3X5UZJH4YOnxsaSUs0N+McStA
6rV2gK6oeOFoTtnhhXPsHCZFE/OOKopB0eSMe3iUL+MdQCUTCotTlHriqhcxwLkU
+xTKENLZW7/jlpatjnM9s9S2h+id8xlh62xeFViDnI0WdzHt1m+itu1D1X34t75q
z/BWEVbvwq5FET4TEixaQiplAfgIYbqF0Ee5ws+HE+wj4vZG3XVTutmXjPi+Vsep
81BflQvNAieAFDXpjw7+OKUNwoPSoUxjajw6PB7c94zTOeo9eIRCnoPaxkVKeEpm
rRrjB3M9c+W7KmxPZpTpW+OB3rekOHydJtofIPCwnJsWw7BazLyDIyw+Zw5xN/tf
6GCSvin6I2JMwHR9Ezw+rMBGQwxaWi1y5WRkFf9RlaonOLsCSIScGPgSMxdWKfGE
54E7GnnJjyrRM1JOXc48gYX6AAkYRJaM2Ftx5P1oIY3raJafuP0dIPmLwkz5xxfX
/mkSzTVR4Ge85NvvEPBGihWCPwho7XXBJtES41XfFx6CD11tjSoUk1LfAiAMU+pV
0JPt1n3jwTLSoITNq8tcLKNma5gmUcAqEwEZ+1XjXy4lrwUyOHRBgFypeHHKPsGV
AeedlJysokqfwoKjRRHlctOr3WixK4t12Urma6pMtwX41HcMgf1xly03CPAw8Fqg
t5y2fq46oKDo3zHtOzC4PO24VgsovC6yW4vDZcHaAvwmEkWZPceDmRHrbScaczVl
KcF4NXz7z+jAUNpplz2WdYW5xlXNUzQZGCqH0NhHKznayyeXpYTqhbE/rTAxrzIU
jkj0XWlsm5DQaNmMCQdcJa4s+WpUzK9V8wZqcV7ut+tldRqEg92+0X8MwXpCAMVo
PCnxmxIhaltZNHDGoKIWnu/Tc8tjeI1G5engx3mtZ7Trg6deVeFgtsoXPfKeP+gp
cFsqcigZWdoqJvqWcmrFy5gfC5ciTE/V6LwfoQNMR3Dz+DvOSpDJ2BVsiA9gH5N6
vDRQkGATAEZ43W9QsePlfQ3Mr19sy/m1dZdmUkxn94zImi2fY4Qo1pxxBgY9LWFW
69gjlcDLtyAeLKgAQHA9a5poWkq2iCG4Bn6z9RW5J79Mnk17lPKJpSYaqDDYgOfx
jpzXHPcVbybQNjuFK/AeqqV9fotjgpau+6kTfZHiz3OUzdViiTKMAc1WaCr/pJU1
coyaJ19zvdEW8q0NJ77cenE8zsfpBHutn9F9M/4XEOe5mu8h5zsoKjH4OeOUsJB4
iszCeFdRfUW3kKcr7Kr0mWFDuN5MYpkQ+nL6n0qTqonbmXjGvRXGcFhNxuZwqEHp
+p/qXGSLZK4vokxYKN2HJzUN25+Iu5hWtgkX8BfCHSL/WEUgYP9ThjAlUsxe0XSy
1CqGSYp/4PnXdt0yqgmMe64CokrF6dukB+vm4yinycFU8H+xBziOCtZcpPRq7BmW
EUkWGPmOxoQ7bWQzMqDghXENGzl3z4sSYRWihihBt3YoiHQo5riNVpOlKYJI1eqE
+V6yRnbmz/QnukszPjCyInhflCAl9+IlpYBScLSf+95B7lqjEbLdoAZxbgfvVvL5
b4cWb5pmy2P7tKZmoSjpDT8Dv0RIXCMN06ZtjXj2krclXWytrxIi+3btlOsuzgw2
r3koEBdC9D1bVwHFqn87vZay7tbDFlQLMxql9iQX7386U/r4QxcpYI8tN1+U2gDZ
YaN6BYLXeja6ZyqDzkc8Uza3/78l0jRHq+O6hFyfovj9L7k+IIL689DN/GVnuqp9
Cp3aEO4fF7EFeFwa4b+BtXdLTJ2uPrszJ2Yq+ookJwjLU7kDL3lwaMoYYOebbL7C
ieWzL2LYhmIysPRKDpk3FODx5aqSxwBBsVlhDd9nWA80RnZTar0zdp/Q/gVh7P+K
89nCDrvEQ/QhKyNmPHtl3DYOg2vzwNFNtQWqlXq4zkllrms232XY9Mtj7333aXdv
1UK3OalEJjpI9MFJhdp2AIFQLt4A2FOun3CgklAr0vI1Z4kBdgJdrEl7E0vqrjeo
v8d3MIReJge0D4koYGxuuhgSgYMa6YtcoSSeMCF0TcfzQCyQdn0Gvx+Ee4iYhT7A
sCvh862pe8pvxGSRgG1kHyZgZXvkCAhHIlMSToiNlhpnerj8UGAeAepGgO7ctpIY
xQMLN8ymWbeBXExYy5V3q5rOw4jiTCekA30AOOAcjSKEMoE7eUqUWh3jkI43Zb4y
T6m4a9mk4b6LlFbAUcWB2GxMGFSGLFHyhmimSMJrzXxTHB3l8fDgY8urSU9f14Vj
TWFiZcCfSfwGfhzZHZML5ZrnuqMrdZIyjNBxAhnhsI0zbUB+AQe2I3yh/EorvJ89
2krIuBWbVhE0gJLSprqAt7eQXy70hNej32a/mlLqLeKqmpYunUkBYalVovk+ejxn
ZmCNgDKFy00LsjKy7w1coCTeUxTWR9L+6nQ/EORwJpIDUBVFxBGK4sh0G3Q2aUpJ
gm2uxmccmuuhzMbdMpMFObJmxntvk9mQZddzdUracXBqHN2MGTZXT9QWoAfaJhP1
WPOIrvXSnNbx4esqtC3dM81NEI0xWsvGf0zxwq7mjqHiVdssYmZftOyqF4V9/muP
0GHWmU2kVbxjOMGleABkJX4h0SAD3B4rL2BiUbfiunBnlc/hoqbWjtRtefy2FNwu
fZr+QVN8ymhbW9J+eV7Ak5PoQeiFxjNFWBtMTkyyHQKtVXCQU5Yktj0e6KT3Z6dK
qpxVxGJsNNryxJ+wAIONMLlp19QRwMfjGq0gOFV2V9C8hTSB2A8S45rsKJ/rhKF4
yNJT24K7+82I2XRUjZvgIWusUV9JVog7XuYuaGbFpDJdUTBg6Z03A9xrEwTIKFLN
B6CdYSzZvKybaUBZ23gT/66K+MdjKtTZ5Kv5fRiyMvU3E46h2PwGQlMgqWLqKfq6
jciGvJInENRpZjGvnKtmko2lgVXjC6HlKno3J5QRCV/mcoJAjIMs90up+GrYuMgy
NnguZvRRxVoBMBrAmOSRFeb1+rOy9xfEbnKT6wvTIQJIuxQDWzRdA9osi+uOJxlV
54y7F6KiYy5boT7O8Vc+16MEdhBgPhcFi6vB5OcftOd3DS0JxJfHNVhMi5pVUsmx
KxdMw5oSgqx7hC4hwf2RkTLu+sL3he8DCaOgnoAVkFPwarrtOGLSTBf2s/VQIP9t
badCDGBR6skvaJScKkJPi++dYDGkok71f4Ug7SBPi6nG2Gn8VyDhn/CU2a73rlmz
WGh9nTCdWYJXy1X9nI6ujTo3D6Tk6/35wf7Y1DPXRYAhPxomw55nMyd4RdwZuJpP
7lZdANKj470gpcwPaVj9ltkbSPxC/vJmT81nkZrSK+D8612hkZXC45UdycW3CMQ4
nAoeWaBczECBRMpQJg37AhIPX4Q82qo4gl/BewONbR58cnwg/8Mv5wAYOiYng2oX
6Mxw/rgJPRgxaQ/5VUH40SRTIPj3a47r2dkX2LGm6Bz3VlRa8XJCR5JHk9HF7m0i
+lsg+6qKjCTfuxqvaNKNGlxtti6ySgSc310WMjDzlj9YgknEMNJ6jH/LwE3WQmri
zBL05UNCD94NU7MPKFOc7CUuDYcinLwGUyHs/wF6Cqv3YCXDtPeLUlLOxxaxpgyR
3NvTFE/L4ocOnzdFslQaNIoiZokF7iOzS8pqWpxg6NJeLt0aXXIo+/a7I247sOUl
Au6aSltSNMYVBIq/tAzqBtu8skqG4QaBOAd+Uq5/ZCA1gBkxhD4W+Zt2XDGbnn00
dsNwW8ZFUG8XXmOAXWxFpiRqKzn7FLRdK/tZ8nh6n1B4XZn+hC8YhRwC7WgyWCvs
noFrP6/jUAlptMUlNmgcjX3HG0AygWY8naKYRqb6Yc/M+YDl3X6lP0NYe8QwmUE2
gZHj+DTbFPTwFaly1TLHUIAYRK3Qf1djXaz/wS7QuJ3YMmZJLfXmmqh8JmxC74Eg
uLZJypGoPuTGRkA4aWAp9QbNdQ0tvBismJv71XwstlPXifg2GiGC3DJSIpjIdGvi
NBWH6pV0DxwOn9hGCgWGdHM8f8f4zH7cUtkDAs3yLEhNyl1Hx+bwLrdwyEUJsWCp
5+K5rhJP0Ic0XsYFWyYFvpgWII34gIbUCNIQTX4GUgl+MN9pao1C/1yKcasL57RQ
wWwh2zlbJHGDoNdJTkhpXUUYd6KXn9ge1ZiO7/YhmmztxQ4xz11LTtznCs60Q8JU
ydqOJZDPsFtIkGX6zpyS/IrVTOTwYxdkLcR2BTbx2/kRB7yKARbjI/H16esiKIaH
m6A7FACC01HuJ3B/BSmjDog/Nksq04YSsupejGsIMYdAhtuQA1mm6CUT7PxBoX11
F+cby/MaJ8gEYZZCs9o16YN3pIyyLKIvxiQoOumCaC29MIaDOe6R+fUdfk0CRXtu
07nb0QT6rVj9+5cKbZ6s5p52HC4JtZpCgI5Ycl7iIlN3WT+0cK8Afmtw7Oicg2S8
3YnJmRBvhh0PMjiUiHT4ulMZ8qoFe6lzUjsHh4FcD/AVZ76Ehs9su34ljcclSt8a
UmLxm3l7VdFTgpj6GH8xb53jIWUS770CvEk+wdGdhlooe2cBhr0oIeYv/wn/wZZ3
m7dozyRSbsWKdx0GMLvPe27b2/+d35WwWm7NDpFaY1HI9kEXkSs5GZ9o5euQPn5d
VWOTNDStC5y0Zllfyqw06wYr7tnku2bJVoXiusy5ZUl3RxifKuC+b3OAt8/zZXk1
s5A93UUgtXJrrc3TVX6T4WLkgevpmzt5Cxk36rnifkQ3LHLpkfVykYJ81OBIO0qO
/ZLZrzSfCIf8yHDOuhDMuLjCUrty33plWhOjyrYn+JSUw6kzIvdUbP73yC2+1612
OplB2AeyZBkBdzPH5qIwh4VIPaf9nK+2x3QOoRu5cY5e4RpG9yNCtyNsw51AswZz
JhdM95wSZ5G+AmRO8IbOmWxnDNw34YyOScqPCOb0SgESpK49t/7eCiy5ZVACqfYr
dg0StYt/ChXAwRSvB5j1aE3/r5x9mugkzFB8iv2sl4LRjKBD1OcImQLhToF/mXLl
95eMQ8OeiUuaPXT4r3En76Z1MKHs7NcZAPWXij6+SR9qcii/qw0Gi26rBsErp4gS
lOhoRBwySPYiVGEFGxtfUr3mJoeXwgX/ntV4Dh0nAMAMSuu5sakwV2YCEkbmkJ05
uN6IEbww63HFkA1Hr8CgryTSkGlzl+XhcHIk1plJARc4LXmFItRbkpVNfId5CifV
C2hhjlYZWsvCReHi9QJhyRKQV2WuVeJPOO8mlmutPIjH1cHlsHGF50dX0vwFyNr3
6SFWqDLeokcQgK3Nt6sT0GvgJFcQnIDtBlik5/XPPf5BCqUG4Eh69K4eTOjjN70F
44mB5TdYK5HKSrSW0Nr/EabSJxon4OX0l4pB4ee/0fk0cSB/iT6f7Wh5FLUDgxp1
D2XNfAuqIJLCKGomaCJY/8RyniwMF+Kk5jP73fS8DjhN9sR/CUdrc6xUCq7nFuzi
XNtrQCviwAvVp2qMqOVGbM9C9u6WLHH6DPqt1etMRgcwbcUl1Vqj2jDZ1CTdMnJd
N/jueCipH5nH4/0AHdMH+X/VCiCVHewe8K2dgpqktnzswGWyFsR0zcreTWz46RYj
zZ+f8QkIszDThZXJKDb/aHj6UI+/vRPIywmkvKBAK2OaZbobwBAZMpKUNktAPLJ+
t6+NXV2g7weZbgPEePFsJfQ3AS34ivr4pPKXfMZBLzKRucMCXzbWATbCooIWcr9X
O1EN+iPi1ARnDmuJCq4PkMsWb68bRM7BzSu62o2MEy+Pe37YBASv+DOBqcb4bPcU
+whhn3908zN/IEbsS+NFFZ4ns4Bc31y+9WeSSOGE6VAGlPgTiriakcrWrJvNbbOA
Jgfm8tUdlZrATTu6SiCyGljkHdDfW2zS/KKtC0rWlGDXG6tJL58uNTMf4tkpgFrg
PBedFrIBNDS7Bd08ZKWGbAN8Iafg8wGmR9fndFMpuplw9TC7UQLoG/Z9VZfFJP90
26sa10a9DQGMSbp2cL+AbDhe6nJco8aUBLzwACk998N0tv8VPR3eWVoBT+Cz6Dfp
OzpBm6nPVnpOw3mYiZrpgoepKKuJxlNbZy3xjdCLaslDlXb+oPoncxGkia8+CAmS
eLuc/zeJlAxUuOJa24hLDGvv2QkFtIx3OoW+66zaFMeJQE8wXZp/LtUPFQtC2dJE
CIDNB4bOGDg2yoOHfuBUN9KvRZYewNjq7ai5ZWn8uKrCvQREFd0RDkgcnym8/sYv
ixKvb0WYI7yvfVlzb0LOBZDrrP5RfCUbNsp4Dh6DFSaftetSLQevmxdcDQM5CLtI
M1o/AOQIDeTUJO2AJYLNxL/SKe/K83zCXhrdQkz0ASqbnEPpeY6GTOygzwVk3yuM
2fljfxHfft3iiAOgd2NSFJ/eFg7vtlAO7AB2V87NdtxzXwz1HRs4pU1nvjuqjqG9
txPLCzumyOIUoIeI2IX54dCiY9LKOedmxHyKQLu02oeoXvK/XM/JmCHmhetFJOv3
Kh3sJEloBjtFX7nuY6dbcUQAy3WqomL8lCszaxrznAFMY7/ihIwZqK/67c8g+MfD
aG/s24Ex/5EoMuzdE1BLm7nDgLl1Db3jJXl7Z8yr1HyjFuzg2zsEKUu14u/6efW6
QT6nERReeq5Dg07ycHiRpGZnQ49d6jh44bYDMfysmA61qfGB9qOA293jIi2OCreJ
R8W0eWpLb1iz0S3ii7Fdu27H1siavtsyiiBmCy9AasAV8Dq4f/PDWIKPR23Ik5Hp
oKtRhbloT/CypIyyKoe7l+wwFKsboBGyIBVCddlKF3Yq2AP6Y0inHHe/CnT1hM0R
EHlLlAazDFKj+7ZtIiWDPn+/DaZ9ItZOOANX52P3iTs7NcQ03Rnlw3Icy95XMq5L
qEz6N9Qv6BDxvT0q6KHUh3gIE+2UxCDzbfXDZENf1+Yx7jQPgwF8RV1PIr00QUFo
qIjNv6ByjNeMnSPgkTxOZ1ix4ewHiO5JEniFQnnPxoKBxIyr3TsiTZi+WbIRZlYS
pM4lMfzCd7MD1KaYUZksYr+ntT7YEry0QlDOy/DdjhEYpn7GUnRAVrt9bATUjfpG
0FfqyTEMSZ2sC6LYzUTIrTLkyTm2gshBJkzNP39rAPoFsgbRYNOXAhLzNj+7I1bo
UXz4Cb7PnhLeM9Cxobu3iF/ZiVw6Vy2LUoTuGvuEJzndFoF9KM+IBKNAG0x1ypz4
mWYtP2H6XwTMGoVh+HoRpQzN9p2DOzw9NyY02S7DYjoEKBSweZLR9S8PGJbmOktp
lKniLa+E2em42rSXWbD/mVHPx/V+D9ItQXKMS4W0RaD7RMwayrcdfv9FNce8mLFo
0KKcvDCs/6pic0+MM2cSY0NqIijpfKugNpUKmqg484fBis63H5Zuhu/x5EnwJ40L
Bnvt7OzFWHwYQL2Oc0Vvmdlcb7ewhU4JiovpRzhQyRQ99W89ITvLlE0BLn5v7S+0
tQyoCBzVe6dzUaIjDBYnhxsl/j8MlEwVbuFpbSO+5uYQSg8MwnBMWRW1+P/U3fs2
Nv4nHik37agL23dDTMXwSSWyFwX9VG3GFaDnG0z7AgWBn2QMM4GxHAOonzQTGqbw
RNSZHLjCEE53TOEd0mA9pcBp8eZ0uI/71QHS/H1tdBYQL2DsR8dWCLETXsoc4MAn
YzFGbHbLgXA8pVSGSQIYGDbYiTtT6Ir2Taw0UEDssA2Ee7cAgIgUFjiwW/5fDEnw
wYnHY9KlKGuXG8OCWgTntAQUOv/XriB/W59EYyClTIGQVYCeT5E/yrZLiyVKHV7u
G+Ttdqho/EIcO0JunTVdruDJ1l74qT2XgioXZqiAY1PWpZyrmJvE36gSneVfHbLm
ueK3y0UeF8eQ3WJTys96pAec395pYJQj2A3BA+hRtGqQqMdfa7jyXpUKgF8fsmbS
9qQDwIpkKqneWIxkFndFNymiwHccZsP80W4bP2EsSCjX7rqezjxHaVsJgrtELJRV
tccR2PHT383gvxJzPF7SSTK2LGTXFB0qluhYxM09YtSVXTQvBhBsgKGSjq2FUMvh
L2MoyXo9r3Ny8e+01adPxGstQVGowFKk41kSxI8z2ZHrp2v4b3YhRpYYhBijzs25
LXMWaVuwb97rBmUTeb3JuDSbg64FR6GzNgK+n3UcGG4F1hvn7bKRcKm9M5qg23Bn
zFy5oNhXeHgUAkSOeiWL9BXc9E5XqDkCaCMamwn1di6EepKeb3jDczlzClsUaHjR
9CSONskuo7FlhjoyHN74FxAJNCwyN8ooBpeU8aq2B4PeuxKnqX6JwPzujq88FJ7k
FWy1olJN+lVaTEjFY51VpQZC4lK2JvfRqONTRjidfXxG7uLUFLmvVn5HkqAUHWsz
0YW12ziw+D4o5/NmIEiyHr8SXbPwdpZzblUP3KCPkBaSbQpmXKZlnymD9YTt4Gf7
BOvSZLCN3dgPZ+PDBCUSvYQKyTlTRfwD0ywB4n7rbQeXscWYXkT5IiGkzqacKPc6
4B9+lFBqZgR+piovwkGDZ7edaycF9YiKkFJ8IrlNxGG1qdnhHrCXnd9ZbMlvoW/7
xQ6YExpMmEgk+t4ogaHpKF2zi7S+5p5RDm2Nm2WkMsoZtyETbqITq7uxwbZpD/Py
88CHl8puYd4pQo//q2XbVlqOKNZxsoBAVO77XcNY45WAtTnjqIM3iTawZBwhBkeh
w70Z3jYARrcHOEvn1cUil/g6cnQqEx/2+6CfHKUPAmO4+KVHGg3p+LAA2tnqOy29
rAiOSEHOiCbDuSVLm3xYNtBolmcrZbEBhht8i6XNww055eIAOAMaZIan0Pi59aKQ
A9nX83rkzvd0i/TMG18AgLsYzW6bbLlqcnHURjj6ALF4DtDNtKvUroxvaz5cp9iG
9UDZ+xnJ3HkShFqG2yl5F5F7wfGQKUZjyXrvN8p4UI44HLS3hZcserm8Z1299G5S
fMjMY8jdYRd6ucp4FZ7DYo+GC/LfvQIDYncRDHvErWNZ/X/55/JZUoCKc2UMWN1r
I+4Q61TCXda2o3cP83kjTmGcLOOolVCyH6AFDNVp/Yv21b3KK4+98b8iAmtldcYs
UjskccTJUlBZ8aRK0budJqLRq1YrtZ261yI2g+vwz/5fhTjXwG2Ulpuba6c2D7I0
93j2bcCJw+XYC2+rkM2Xn9hbpcCKtgaBTCORbHWIAAnDwT7IFNNglqaaPQ/gxu7x
BJUx6bpvVhqWvMxz/GdeYE/9PsynoAS/ztpVJC/q/EEwrpkXBiodT0PLDmQ6oQHA
8LrZ29EYjUxJfoAk2zMDE07tq715It22KBheWsLsO3UUoVmzK/SB8oYHIG/kQ6tY
8CI3crCLNfTXqundM08BVNbHuf8xmb6G+76pQxGL3zUqTdc1tpkurDVjXT1YPj2O
+mbGMVNAFU/VDUCytJwx7+lLwHWv8WGmq3AjxBMzBiujaWLaTJtWB+lFRkb9W9AK
VjOju7Rf7ayZFGs4aRGfZuArvs1Rs/bR/rISjL2U+gfON/mRsSM9zqwML2EYPvPt
yj2odkQG7xtC1EDI8pvYf0nZz/kfRybcwEaq3GGvVhAAq35DvHR5DtivWhYPbeez
vsWBWx06PjmxmXyo9wkbgzpq3n0QUI8/0CxPyJuRUD4j2BzqLbcOkAjzGSNvvv9s
aoA0yKUP/bjaZXcHR6LhiUclF+lvaItwSbdTKhh6T6Tzm6OALG7aAeu8sKBENKEH
fk77er9rd9Zm+QLyNR44O8lTd/qxPEWE/zG5uf4sRgYTOvrVHevp1IKnGKgsz8Kw
`protect END_PROTECTED
