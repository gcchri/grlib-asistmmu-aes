`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MuNHefPuZNhavhaMClDvSH8uTJdjpn8+59f8DQQnpOES1Bc0vndmHKBw+QpN7C+y
T37icwquJRg/m/9p932YUSmHHjq55na8RUbtzzfQlR1xDd1Fe6hes6Lkl3RlJ88K
V+55l5S2Y0xlzHDhQar2CuHPO/7NHJ+Irjj74VNJs8DBAoNJxYp7toKcgrTSnOO3
Z3dP9D94le8s2i1KcIwfhr7wMIi9Zbmge2WNlG+taCAWHH/aEuadYk9XflaSINtR
ZomjG5T4+EP/d2TIoldjAiVIgGlb1elwO29LA233E7PFfoKnouEt2puqGxxyuxh/
XbharulNXZ14LdUxsPsQCrWqWda31LhrpIyTsD8vjD9PHZ1vZYvuUxDHLPD10AN7
z6cXgew28msfeksAZMXABmWw7vuTzSe+MIyW3e4pjNEvuJpIs9acsrzefo2UN5Td
YWA2YjS/V3NqZVQ2V8qXugoT6Q4l5vK2W349BXTOeYGt0GBGJuOcHpGxchIUCixp
Ro7xL5hka3qtXaEoClzuhKOKeEeRT4jkblsi2LHZtxrAQsFbAnbVsXyA0MTSHqD7
9PqImcUDRh0ytF+/33mHca5JLE1iczfsYd8zsfZ4QpEZQA9vpFqNEO7Gsbymgp3c
3UxDgKXBucS6GSL+kYN9vw==
`protect END_PROTECTED
