`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o6S1g4Vatxl+Z1iWeDvHHnl39I8tbNJuViifUwo25THgRvm/z6ND1RFiJvcNRO6s
mZkjuw77eQr11hfRgWNRUQK2spwVWCcSZpB1BhzrdRFSfS9lY7hQzbcKzIuorMZL
LhxNUmXdLWG0y984SuplZAW5v6h7HM6CGi87RiooWkBYjF1mFjyAG9exZqm/19da
KeTbUn7OrIbe0tJNox84ON6Hv1EF3HTmBYsZDBFGMZQrRSyFTh+NQd8dvUDocBOP
Q/r7+fOPP9d0o9Arnnlm0bkD/VY/nPJjPBtw0mpAFG5EFBuU40YUI3zCVsJSEJVy
UF1ASuepZYIpeN44Iq635IaCKOzkLAWwaaDbEKktT284foRZHqXLNfjEP/TyUM/Z
LRFAhrLg2Z8DsTYsFjUxr417O8c4hs+0ke2oOT2ohImnXMNuaGvlqyDC2D6ipOPz
WeWyzyBw/GqnVtGXkY6KqmwrvMH/lqwmqDS9jo606KOOEUmS9B8s45aCeO4olo1C
`protect END_PROTECTED
