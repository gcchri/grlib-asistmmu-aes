`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ix1+qQyxjdLMxJhO27dXvI/d/13z8f3N/ct9uu5WxTNyv0KHd7d0ZmRn+jqyGJ6p
JHgJ9qUUnro3lLw4MBBDBWqkGR83qJWeXZanGYPxLJBn2+WcJ9HHwpXN++7xemvl
Y5rKquvAHgG9j7VBgq8+HISUoZoWYy6xZYQEmDFdG3IU+PvN6xeXV9ud3CmCK907
c1F05BX3kKIOAJKLIzgQzDBrh276WZkfTZChEEM2euACG69yj4p+ea+M+R4uYrXJ
JuCuy2R9jdqTIUg7WgeL0fKCKmUDffSGKVXeMZO8E8OcYWKENUuNOBZu0I3tviU3
HkWgWGUGlxfAK46zW7jbL23KT6ThYwMU13Dil3pZwmI=
`protect END_PROTECTED
