`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BVwiiNRqwLNtEltYrAPPoNBwBqyw3Ff0quv3NzYUVay5S5fyV3o/P4ASX5MrAyHy
2Tbzv/s97pHDge4thdb5q0vaNogo08d7WliPec7U/mfNifPiwSrWQfK1zTQO0yHI
xFMvZ1bv5hNGeB3Kl/OJ0OYeGRBkfy31avRtqe3yLV50/cXtOvjoPSZX62JHF1gt
nc9wX0pkrtUPIBuI3zPANFYLaaqJcd0gY76N24cSUP+YAj9x4zOtCJV+cmYO0yDb
lDdzhOQXzkcWWoXlSli9Yf9GIVDraSfZXLcLhG5ffILaxs6BcXmdRuY0VhaXa0lm
FBUPV6saYH14giLWfL+atrrgTCfOBewbgypngldGI8OaRoQLs1xcPvEQSv1ah2Y0
ptNfPQeISvy4K/6H07bW1w==
`protect END_PROTECTED
