`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1lG1UzxtiOVVuHIAKxE5GRs3spFbpgTB9TY1ZVHwj8b3iQ5uXT0t2cuYqq98LI73
qu2Zr3oPez03SUQWxsXXfdfPxCIbzStVLHf6g1TWvldwdBN4qALjSqBGHD96NYWo
LDXLUXFBwUbyOz4WzWXGuHrzGqboNJvNX6tq623eOYmbxmLJLZxjNFYyxUOXUBwP
rXBR+RESc+BJXefnBHQ79mvRqb2F4cBzkfKOY6mlGu8GDO9Nrnk+GBMnhlTQrk0q
UZrG9BsqtSlVYmVT8L23IfZZ7wxUxHTo/5AjC2HQgCdjaUw18/k51Ugu50f3vf0c
kjPCyDQ/O7Swznr+TDlqUOWF7qggR7m/AX035ZkzucNuir2RDMpyOWCXyGV42fp8
`protect END_PROTECTED
