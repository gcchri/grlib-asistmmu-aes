`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LgdP96V5c4g2MJzWaqriSF2sSPJEot3YBDHFwyTzyKpHqWbqLjv+OSCRTtVpWUc5
yjvzQJXkvqwBTUyRLKfNuoV85aH6l79/NOZLQjWRK1Yuyjygm3t+W9dZChlWjTdD
La60PJPhK395B9Wx3CyqRaHzHSS1MrMX4ULOC9y8LS/i9J5AiGtjZpG68pohewK9
4wd0jYgVWwbJcDv6Qx7HkomG0TNqLbLfiy1RfOmDhi9rvN0u6VTRQRp/ste49Tt5
6ptQ4VbTLhW3NHc1102VC5I7vopwqTLvakbA5OplT5Y=
`protect END_PROTECTED
