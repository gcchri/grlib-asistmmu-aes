`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A37uBYRm/VPuxFfFyJpYWo/FJOb3IBTLoEVIBG+vlvce2/lnuVYHfplZXGtn7n2r
uLJJ06L2RNKrU851AdY6AvkynkKp3rQvid68PA6ZlP3xuNgCN0XCMmm3roAAlvdx
X0W+q8pxYh9XhqLsu5DF5lch1o4cLOZZq54EINmMDWZIhhaTwGWGDz1h5QxTAyQA
gBUoyLN6/Q+snqyotv0HTn4mIGFjIvcW6ZlkRyfpjF9TLzorZxRD8m/Ws/vKc+22
RFRnNvIldL/27BfQBlAfAlfbHWA7gBRO7xMv8iys6SZiBa8DB1LtrNjA/q2jR596
Eo3mvEvHDk6XDVvVXHFLKUJa/F05bNPUhoK6wVeUcFl9/hhMk72OJqIGDOa6Ix7A
7vnz6w/nz6xtgXSa73oxd2M/hi+OfHx9pQpQB/udZHrQh5Xxu7DcOr+DKP+H8USl
Vi8o2y/3ZFiM5Gnfs2FSMDTk/CJ7Ml5I5Rs61R9/cQWB8Z80euEBN2nkW6+8kwD/
yVB9rX+gZYCg+U9HrCiVsprehuoLAmSIw2/lF8dFxl1C8c1ojpN/wHZtSPIcLqZL
+6R/JXaFbtI0eFV8SYMC43dTQSlkmhciTqyDNkeZv4l6O+zCstF4pwkihGvaerZJ
E9hHssmt2EOnIbQqX/irZg==
`protect END_PROTECTED
