`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gG/0pcmzJLLeCMR5kcC7AikXL+Bhc3QwCaC5y48St4evvsDi2UYxUEBYetMho9Ai
c99aBJhnPuej426udomPZH/V2ViMIFMKT8qkx3poKO6wSBlKRfGy5EC0zeRDUvLC
TAvG3lNaZrwUUh5+NXc3ayQTfVdDYn0eG6youX/CfYnQbTPoQicYPaq08IEqEG6+
kj4afw6lDUEIMvrSyoAjTE1HV/ZcBkgac/iZ9aoQggcV4gXyHms/HDp1fH14PsGT
oT8fKINGTFk4uyJ1kfiawPcxlFmvZJeUgjqpQfJIezO+ovjRZLVR8XD3kT9nccea
M7+C1irUo3on/+w1YDT30OFSL+PjBUkGDf22g+x/ar+Qb6fl7Ur6gjNjX020vCQd
hAyAtUfoGwaw9J744CnQXon8mcO0Fg/c7KbOT17KT4qmtXLSVmawA8tXG2B9vAKj
GmJo72M2RFb2D6WeANjB3U3XfTP/Op/4CEOTAc0J/Pd5pTEt6ZQlkFCtkdoRKlKz
aSvt3DSd6WgK64qMqzumKZxek0UHfrS78jwP/lu/yvrjkOZA72DuNRqax5AC6fx7
m6kX2ZqtXbXUaOSki/MG4sSABXrJRmgXTlpXlJmvMkwXPTy7gWr+//y6EdqK+nkS
j7781T6TuHI699Kcn+ecdjWVwtLjyFULJW42lV3K4o2jabLX6x+LaBRsg+57GWD2
fLcW74QeCM8HrdvcGnxxnn+exc47wWtzW7xN6H/xu83OTNwr+A/byvhAq1m/86mw
`protect END_PROTECTED
