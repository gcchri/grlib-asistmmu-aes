`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xe0RxZA9k8N4XSlSn19E4GOl+8818R2fM63wxGfmTMvXA/7ZkEDsNAxcKyXKG9Nt
c/a+8lOpDKqHYn68eTjse0wYjJIMgadoIDEMzqekBLSneLQ6hrold+uKVLzk8Yyk
w/r1qg5CzeoQ/PpRYqFXltGRHn3FlvrJ8bSmlSI72v8m6v/0xy/KrvzoY3fv3Gp9
SwITZB7WwjzaPwOG6fLXa3TG9j/dClj6/gozjtzh4GCsy2TNx3smYXAhVwUlF/Wl
UdMCLvTYQtMMB0CDSrSlmjabA14nSLVFqOSrEvLQLw3O1lGSKP4C7vAVTfy0PXJd
a9U2BJJtI6QNWENJHSrYK8RX0H5/4VNU9uRvQrSlZQlz+IDRc3tCysfY9riZfrmy
cz46wd2fK25u58+N1cDgvP8GvaTn5M9rds4CM1Kf+/KUYMK2KE/VLB4C2gO97qhF
NbFIs4DP9p4fq8wQ6VIy99J4wr9irDCMpU98ll5hpqqzL50OW0Atb6+pz3BmcPD5
KBMQu0BTC5YTazKA37ImHNuVOhQ+czTiCcnLvjYaVS/6LyhQ/7MGzsbleKAImE/O
NafmttegZlNbeM13k9XzJ5KPfeXun+v2nv0SoDvRZL9HlydHRb8J4Q7NzrxlJScW
u7qr42YzXgj3r/H3pE3AI3mG/TXIBmTFHFjxjoVy/m5cb86JD3IeYXrDBqdb32Y4
rNyso9KT6uhxONSpLgmN6PLDuEBTZH+AExVCTjdjy9EWSAss3FhesZfZJaAk/Q0S
/AcEqE1oH0UDgk/SmU3l4fupKs8wiIpqmWgame3JdTnQHhrcMOQ9dUEQI87cdcZB
F52hNOhxpCdmlc+CP3snXttVbatJ+QtO8DScYa9tB7cMvmAB0AQP87K/7w3ED0ZA
rmKay4tMTrN2JkK7cdQHtG1bg7e8wcMcPox+W8CKnMNg+MBjFVb23+mQJUkQsKit
ocfz72SJnTfKbugoqXQhHFJhDfwDK9q+xNbppSmmCPyTlNO0eefj7iGircOSSULL
xL5FUTVvXZy/dvNinvcl9yqkInDtpXHbPNH8CuYbFulAvStrfbkaUIeuecrErNSp
u1O8ySxrF8FbpGotrQD4sNMDL6D5/bhBo3m80DxknkuHhEVE8pKWjXVtbAP2sLDZ
vCRum3cQKRVBb2rUqKsC1XokKnwi4d9wOhBdbKr0Y7YOWAvrS46EGuViCekvPxJ3
ZsbGLJmFaQGOg8AGq5rZWbvrc8Yr5ahXIGb6VN4eHoBVDVI401b0i9AzreNwQe1Z
qURXNAX6JWYB2aY6FPHjWNdfMYJ78pKpeqxD+j1D2nj9vMozTjfjQEk9e2mb+wFd
fEhT9hQKHkEroRcYhsvU/XnzpDfZZ1C/Ft4l24i+JKJ1wbhAc3ibTehXHXH42Q1A
J8iyoc9e0sG3IoHnMHixHcpoYWuQhx8YFhTu5NRyDLXEmD1b+IbtfHTgck11AzDQ
L82H1fE+KzaMb14Hs45IyPtlbfbPFxTX0aLoFud/Ws2zjLgSn/POL197/frGVEGW
1C51TtW8fYX9QJWXKQsJPPFTOgFayfhpb7KUc2AR6SpGmKOHyY6/HYlbnFfnW9Sz
xtzNnU2YFxuRrOnHRCtbJWleIBbdkcj15fHRqFmYxufMIAj/Aio8ZEozXlj/x68Z
MLENjMpojqT2ls81YrRvrGHyGS8eFQMvoKvOl6BvZMJ0sREYMpCaZGzuF4Mslh3v
L+PVrNulDr2IaawwlnF+8lnH3djn+wQPWpWpoRI1NQVzkFua81TnRSzjTRw7WYGq
mSIpCi+g6IC5UjjPb79iYQDmGgrxpv1ahPX+GIZ+uB7UNbxEkvpIuSGot7r2gtfn
I4/BUJDdb8KN4uvR6SlRVb3ufrD7QmNHJmyo7AdUBquY/PWG4yRnf4mGCU0GlnRw
09v2k1TTkJxfq2Zx5h8gtkMxcTbYsVSqogCCDFchdNLi3UTttxHd27wwx77aGXSN
/JK6xr0TsasA0gPUvwiP9yLRG6l6QRla7Kxc/tjTt8H+7Mjymceyv0A7yFXDU+vl
KbUd7OZBNkCnDpP7f7BoQixG1l3axt9xHZeHShsx1cXbKQJavrymSUJk3NKnhhf9
XL/1zwYydFPzJs9wxmi9Q5QIW6g3PXCTXoAF29ML5to285Bn72FzwgTz6Lqv9GG4
y2PT0EyaasElzs4LgoQS7rP7wesFMFo+//29OCC5QaDqppl/kBIqDKBD3NDprOh1
k8Xu8iWdjtWmnDOOPNo0E8w2efiy3waPfK6ukMvn5lOBgaKGdusb88WFdsYCtkEh
HyFgrZ/jrwU65GDxNCgw9O2uNkGvJLq/x7ikttZF3ReRisDcsJIoFVANuyr+d1mn
UptxlhkGWhjp0baeRPRznLEAJ5teD4vTyb9v8U2TmbT8o3r79rSUuNPb9cHVC8Xn
EJBooNtkRem2963VIpKWvmUizRgDkZnBgisGrudI+cF3swrbAJe4hPJokYvZWIko
fqaIfH4De5QjXl/xBymTfTuHJEbVQNPcq5tT64irLv3tzWJ2Z5ePPjOipeCng4Py
0yUwXH3Evnr9MT6j/yBJGR0TbLDsc2s+0L8u9lrAr4I7D9zjUMNFz/PLwpkn8QIt
7LpAdJA3OyMeICCvY1fpLU8w1gvRqJ47w+WhH2CEr5D9ptJ3YfLg6+7oKzSxNKiD
dsE31uRHhyYkSGi+WmqA6Gibi4EZIIpsUHDFELuWDDN2dFq9W6Psq9aRKrCJydA3
sxCXIICNZfG+FfygXvUYbVKMY5lsmV7n+9z6eH8DeaAruiugQiyhaZO7CNSSr9mr
/I4qs04Uo66gDy9WFtoAdZ0IGwmDjsPCmx/luOeBW2+rMw+wpo0zrnyM9Wq3g81w
LANfSIz+sl7A0x0BNgmDqv/6YQMnB+eRSGPr48Tybr++amAKdRi8cVgPUONNnjOp
AFK+QmDbv7U+oveknMJvaDiB7pKODhSyWtq2enmdEpA4Ito9PxTgvhM43jUwn9XF
tr8ByOXo/Ox17MEPHH0sVGpu6cwH0Mxpvv/xVOttFVNdVh9GvEhuz7Bpk4EcTRDL
1elX7B9SR58UtI9Jednk2V89zEdUjwgz5Vwx56zp8nRdVtWGIv708wcm5cv0XjXC
9Z6goCKzKyH6tk14eiAKRVNjXa+Jo2SwLDaXKCCBh/azqMh9XbiXbzG6rBGYm1qk
JRIvJD6C3pogn40+NGQxmHaW1IRUiHc79us4849CK7NuIAGo6bbnSiEkqIOzbg8y
Ges7tCW12W5stba79oFdveff4GMq6f2d8y0dwhlpFxHihVV7Dv2Jfip6+JDhY5iC
gVUb9oeKSdTnOpcjitr5HzINkCW2tpRkpvu+678v3QxnN0eNNrkYHnpddaoT8g+H
fUCMc5B3LXuAIHOr94euoZfQv/tqpyJZbU2trXP2pRloRgN7cCPbpLXj0CVXy8uH
Gzbabu6lSCA95UnCB0SP6U/uf8T7BrBNTWds/LiH0m15YJNUakWI1s2Qgx9YJcy3
vmDAzpXMurG+hm0CAraqya4HLkqhJB9CoLcva948A+ZHCcgHmA3VTtD8oz0XWfGw
0bWsmmwcPPJ9pIBWeYDyhiETwL5EUhnCvzpnQUZiQP8IQWrwiD5OOYWJ/ga3wvpV
RFmXPftv1C5Ul6/UyQI6cDGfHS46TUM3ynP172LOuG3dkWWfx38OhD2kTlDZlcA8
ukUMoLIgDquFVp/Z5A6ibxg9n79rm0bUR5kKimLMqxdtCwPtUgBxX9xjwdAm2+EO
K785VpPTEnpQnuTumdggMb0YIrBPJpb6/ueeUV/UhoIGdky8P2Pn5MpvvmOo8Rhe
TLKJikA7hNh42p/DxK/BdG7/+SsdpyqnGxbh4tfOEV0JbAtYh/N3cmbBV0iAQwaW
qoOQfQNuZeU6dH3obREFnptEFCnrPOqHndjGCnHK80rSR6TcOWVC/QMQ9F12ulT0
8PqNUMgnFlNp4HoBYycRv1GNEYPjRZ4c2Po9PWDIXtLZh6F8SoMhAutiboFlK49U
GTkGdRzgvLaeMNPATRguOxRX06X0sn6AgBrY1lCflB1QmR7PU4aknWbOU5NjImou
RV8OM5KBnna+5Xa0E3zi4TRcDlWM2sJoE9o8aKIdlwGFUOIMXjZnPbYOIHbvJv6y
+CkQ28DHY+9zISNCRWN5jfPuhyKynPUVft/MDSziIcSrHyqS1PSho17o/WuGukIw
RiOk3A7uqxxmrsgNmQO6ikwtV6EGcHNO6II/fSHSFeYFqpFpIugHFX+8aBX3K7MD
5GylyWNfrD4INAwsoKjYYtB2qxcLC2iHcX2PyYOiXo9n5vCXadQ6hKxE40TbmGZc
/AOO+YoVu5vERoVSXmoy0P7NkflO4fCweR47rLJ58llf2gQAY4qSo7Gdl80tAyE+
ie8mlx11y+Z27SvmMhB3g7mUP6E1O6re63efToiYn29RGNmvFPGMeEI+2BZvZCV8
3X3J0gQtIBhtIXJasOvdtcvcpMJ5C9OpCiERiXspy/ZPgYqXvRAHBH3lRx/SyeLZ
PbuDLHIuCsWYwl/jl1Y807JaEweua1zM/Kh7WaRM5VnZBuh+0ekhqJqyujHqEz1R
DcYUYHYAoqMBbrp5YUTmO1ptq8kmXZ6FxTs9Mtph/aWIjOmcaG+hMOXKilPXwH8F
sCmaP2C26i9FRrAu//6gTu0aDZNV/C4nvxl1n2C+/LgQDdvaPMWz3YTcYukCxE5R
KXA5R35bgZtcOaDEcFO9u1fGVdYCfQMeSNt7XZgdNYkVoia9M5R9Qeedewce3JTW
6GmF7oqU7vOoFpm0IFfL3p3ecCiPg40rJUf6kkPDT+HJYTXOtkJqDW7yx2f/OPaK
xqmjp+v4RuOUsvJqXKqCx5q8yt4+n5WeFUB8CdS9b46m+TXVr4q7tVpaRvM8jRs7
0XSEn3h5YQHG3F1+Ovsy7L0JegtwnZDaGbbncLp6kPNJLbrEeP6zKbpJEE03KSCI
g+IyyTKfAuLaE+56DeM9oMIVXV2oFMvTkoCDot9foFd4hW9AAUrbbVgNCqXMj4Eq
8JNhSiyN60vozbOT6sCevFqZrhGITRKIECdS0uiQgHyOW3yfaEg4jTL8KBz8PVvL
nOAeO+nBOwsN+8DrMFFApuUQ5tnyhC5bxGm5KnWoFCRBeAtYtgh53ZyDXDWprzRR
2V6ySpubHQz0G94U9xji0zhAGLlmGWOX3OXSFoueq5UtRVkOAu00znXMIe7WKaqA
EuUcrmgsn2Mu+nxU6F36Emk+6EG3LUa5lRTqDh7+MN7QzoFrjyJC2wg1yjVnhv4D
ohN/Wa4cdE3lA3v9xSHDG2LH6wNvrXH/uSlhiBaeopdeiclUprMvHJXhC0n8ZANT
/Uto0FoWHwC6QRB6AnfiG0rUHjC6GH+ZmsoIU7VlNHESFl68PJCIyCvGNzlKkJKh
xzofAP92PJNIwz3CMwTIDzTn064nC9dqQ/sIsdPhq9LhQ29KWu+Ff/mqs2bl4RFf
uOQ2JpZsAhzooMJmo8jtUttrPCN+mAxSycJFYAGERgMJjUXickEDZOwqKytRiU3t
I4u4Vtpo4NY+GRQSsoi4K+ESrjvuV/3jnQPp2uXZ3y541C/KfaukXWtNWpLr5Ef4
r0eid1X/7TKEOpp/RU6cV6M/vyX/fYK7pTY7i/B8eII=
`protect END_PROTECTED
