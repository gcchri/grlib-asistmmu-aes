`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LGPuFThLFHkXuhMjbBVuMW+ty6fsHSgc5Ev/SJvBhReJTKO02zpE6w58O5r6KpCY
gSD/NO1V329cAiPrtyHcwajbOa7pZpiFkF4NJ6I7l4neyfouk5nGv52eoBlrGgBL
mkCtX+6jiWm88GwGaKGFREnEGivNb9RI36Wh4XXgk5kgdvOwcdQJHu17BH51Kd2d
RdHH9oByyabtq586+B+9mYtsHOG3fH/rwSN3Ayw6B9dA4AfSQoyZVmW2ItM4rhbr
sCLrGvc54eQdQYWvu9xu0jmiyAqImljhz1kUaMGKr8ywMIl242HxKy31+fm7QBIi
jyeBXmvhkAb6vLwYKk8geG8jI1glK1mH5Wra0Ns7a1x42a5eoh6GC68ptZrlVFMl
edWayJ4cX1D8v6oREySYA4DsUBbsLOe3PEbJ9nwUAFM7yRbIKcQ9PdstvletMveS
BjcXjILxoP1K+immqF4z5w5cfCPV6zEohfQA1RLBDHWDb/mVcv8tV09e6srsC56n
rS7sTGmThdXDFV/rQv0WkA19CHYfT0OK2ymEFrJDxl1dWEc564lgnHoFUh0vziTh
RDJyEjuy1fLtkiMIgk+Pllt7qJJv4VlpAvopVpCyvW0F/43x+j/rpIYwyBVaPQOx
NO4W/88gGfWzdSodSnYQ5GlISw24RGtG3Ikey35ZfS4umHlROdL6vvaX/w/7pJn+
`protect END_PROTECTED
