`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yfRnOO5UjuTGvMmnGgyNo2FiWVuQ0GIRjwagwGLdwi62Rx6X0Sf3YXJshSOva34i
BYpct05mx5974si6m/9Du38mQNvrFOJ8eqfe8JGswm9YnEsohZ4hKhUYMV8HuwlA
iJnoOez1EgGKVqQy3HFZYyX0gLrOLNNjCUatbaT/TlhtbPj5F2YVPHI2Ly9dUkpU
+yM5TLNp4BkSSp/qbzEdIqrHsYFwhFR3nHGBKC9zFglBCk6vz4yrCWyspw+Q1WKQ
Ffcq+noAdB0yuVNzS4FP2gvq9rSQ12P12vKA5wyXNwWqo1blhl4SzxTGaNB5N8Vu
X8nT3gX0szxDgCFyy0ZChmp4OebCDfTDIFHIL2Y/QmVb1nDz7GQ+Crvg9AGjHnv7
+prNV0gPioO7pzbaRSr4tvPN4bXTtux4TSL7f0Xo/IY=
`protect END_PROTECTED
