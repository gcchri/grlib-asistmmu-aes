`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kZ1DbSgZgw38EPKKJsaiQ87LuIJWRTkYA74pG8/LUzFtNtDdOKOhT6Oz3TQ12MxH
nUxMHEy259mjD1+xecMos0jwWTMbXN8DmRnPBXxRRaDDZjV/FWEOAmBormUf3OBj
w8JlqLlEN4ajyt02Q8fVu6TTKJ3XDRc4JhM8QARYYQ90n7hpHiOEjlcN9evtyCKk
H9hyzAGgARufFQk+XTpKj7XxnPnvdszHOnn2HAt/LIHFlv48LAAstgoZGSft4px1
9BnSU8RIb6s+QY3uI97FiJ/Zxc2MqemRiyBCl+bccwWb9zvlXjM88W7nORjztw7c
GsS00+URXNyACJXxlC2SWK0Yx9R192hSWmkFDC/lzZ04HhHpXQaUs9a5pQDcUJV0
`protect END_PROTECTED
