`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wNBiMbikarCZBeSQZij9a/OIsUmyZv79YHUlGHJTbDmfG93V6lG6yuE3PhZxWIrD
Hc1cboavgnz5abxmN0QbBF3suBA6mzh/bkpYRTJIzX5+c1E1mNArriRJThRp38ft
S3e9N0mVPWF90qnxckrK6MSepAm6JjSvPAiV597w3bNrK0fikdVOEFGD2scWsXmL
uLbe8ufocHes09LdDQD9XQ==
`protect END_PROTECTED
