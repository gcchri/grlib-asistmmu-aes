`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ctkC5Zaft8iiu7Zi+bZpVSY0G/svzdl6RpQrXmEP0ymfIq57I8zoLsoFksFQiT9P
1YrIJ/g2Ys8Mhn/q4euoNKPtl0yUCu0MOHv2nTZsKHswkMLVENoNuhZhPN5Q95bo
NXUAco64L9QNNGjwNgagfM2yXBMBGO2gPlx4dxAVJJXfDwP+VGdV9vm8I7NbquPn
slWPBQGthivmD7rp32nEXw3A6DrFWj+j6pTABzD2MA6WuLbg8Tqfo2zy8yO6YQ7e
`protect END_PROTECTED
