`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TAyT9vB8MUYfCUJaXFE5LI010GMkiTsHuSqVnRNJcglB33qTgd3iSxq11IyG3okb
PLnKuZBlOtV1sdL3Oa0r+imODKPIynHYnV9dK20DYA1Sn5i5bl3auG5fqSz5Hv9Q
fv8+ohEWyr69ep7dv/N/WNmfRixlk6FTw1tOHyJ2GfH7FblNhloMgXdVdDM34KFS
vjtZM6ZTBZmerYTNQIjkttm9sFpWHG6ZxoPu7c7mHU/uBIlEM+O8UKcOlDLzq0ay
FaaLAbaKwX3UFqCfQ9fiiwl8Xq7RvLt7l1d5y0FZvaT1NsAyIKabT5THn62uUpPp
eWACqoSkFRca7kk7CdpsmArztZjRjo1YXDOdqpnB1/1dEdOi8fn7K79JTMfurdo/
ipS/QtP9YEUXJERQQRENjEX7tiTr5YEvFI1yXvgmEahX1BAWDXuIFYLXoTgHcI/p
j7srTM5+v2R7rk0ePiqAwu0bw4BSxtDU/tvH5d14EiqMze1FyLbrUjjqBrTSyqXm
QmC5Qj7NvavbDev0JwZ173d1zCro53bk0jdcQv34AgYsVZeaV90AfUe657Lq/wwK
3khhm1nGXM4eWH7gPGGfJdNm1twAVLS8p3zlB4nGDBi0kxNmmia8Y5rct0Cm7v/h
yowxLE5kgn1siZznkgplNPdLf9nERWkgAOoabbAm9MEpLbm7/qQX3/7EEXQmxsef
pbRnJffNnB0PMv3PUsTXyYSEoESBKxUsFbjn4bE0YXcla7INKOGNygLQK3fgpbWZ
w7e8DsIoUuRzONdA7TbcMrytGOD/+gIYFOIEDNQBjOMYZcCxfYqNtMiGIE/m+3dH
c/RIC7e8rRVW2uH3XZAK2E0BImDeu3srLdPkhg8chzHBD0Sbnke/zweA9gEuJFkF
Z/tu02daoX/8JFLWy5OFpUO+7oqn/7uILNeajZbc2xk=
`protect END_PROTECTED
