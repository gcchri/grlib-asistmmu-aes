`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+tE2SD/QYyZvSEYc+J5WD88aExdLVlNMBs0xAzRGEHMFav6hkaBxISzsvd4MGK7K
luDHVy7j5ZDmJEQCUAJWO9yaNSsw1iy4uEPYp1CjPZzCNi4w9kAcSSznqJdIWcxd
mMd8Qjy+ZigsXKcktYoEwG3pGxwqYkXWBaTt3CqjJqnGJjaC1DlicofFxfISC4cF
pudJOo6ywV4yluDk8rYYoChY+cO2TBkhe5BMfgQxotpMV7om8RPf9ZmecC6EnBcS
XpIBwLABWPTUyndgiucsk2og+zSQhjFBm7x8ZhVtgtzwmMRfnACTFtJ20FB39xcv
rQN+7UawTpxwc5MLV3TU4TG12+Qhvg+GuSlUAmIGUtPQNuJqYyOlMVrXDysKTRDP
aYfxxD4hmAyeuP3nmhgtzVZVM3jy3G2H6kmxLOVjTiLbzo+4mFnimUcn/TpHpSkR
TPKccpzIGyMlUW+zF4MRrb1VHFzal9e0MmLIHOrM3/D4cIeJ70XE2r7mBfhFr5pA
V/JVfAGY5YHNSuMhHYI7vUMn34EJrX/DO/4RpPkK7YqssY9qno1PhUnghSHMGOnl
210aAWh1BUIZQUD7ZrqGNXQ8hnhHLVPSrQMNsnodTNN68KtECG5859y7ptLtLgBm
GrqoIxUfcZeNPp0FMY0uOnPZFPPIhG46zk2JM282n/VoToj+uuJ+JlQbS4DOu1HL
ruPZ9zUs9Ue5Hw8grQCBm6nIEHax8Sfk+eyECGQKh4RA0jGHjYf1t7/Eq6gXuz2T
z41O6xCtPDDuS+NPafPMykg01NADLfedq1kRdL4hRM/G4ivDTFanSKhtTdZ9vsLV
Qsu9omlzs9QipNnBWYTCgPKbTOx3RV8E02o4xGUH8s0oGFcuQKDyPxEsNbdPEq92
`protect END_PROTECTED
