`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b7Kwj3eJOiP9rZIOkCIGfubhy0hqyYxc1ylimkIqG7PbxED5DLiQMobTAC+w9T5z
Zmpor5/3rmm/wVq97PIekZZ3Dv5B4iIgqDvkxUtEqp6qBavqNjIaKvcoM+o9k15/
0G1xc0TAss5JK/Mmqb3jhXULFMBSb+UhyB0rgzl0Ol5axMMJVH3HrXx5RoxX+UTt
MpB+lZdo4Ylemp9XxPPkhNpoNo+s7EYJdiL2MdgrHSKkjFMXGwpcZohOGpqcN1f8
X3XhwboewvwM3OrZhn2975Q0M4c2n6rw0IieuAZKXT4aLW6gY/7lM/80BhiVdhal
kw4Amk4f6slX7ge/49PgtpYrOb/w08bQSUVeGqZpewcft4L0qGqsxpMTaATRG8qg
riI8wGMxPd+iOyp9Ho8dwFMutEEEUqaLtxU8r8zM61wmDoU6c1nT+ndotbsGD0IN
Lp77HYVDePliI2ZKG9x8RRvzf/1KUCIEe6oUPijquoDJGHa9JFrOon4ZFOHg1V+D
APAqk3qC9/U7kViBqWQFIqBHRFccQWcT8kUXy3pYPaVIPlIQ9zfzf9HoRqMRJ5AH
uNweExuEi/Mi7H1JHKsTsviBulBAU0NCD8l/uxOrneyvALz9i3vhZab9O7YyWh+5
EyLvgKsC82zUKtbZt2OEQQ==
`protect END_PROTECTED
