`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xPTvBOjDkyiYpHyRbZWocMHOtCvEoDCNBa7hfmnNfkXDu3EnxA8TBIMs9EBBt7VA
x1wMWDWKnTkGUhZrlAgM0BWVcq12C77WZObmsOJmYhUCkRIduTACNK8nQRjScHpk
U+bkdHYTYnlIIfEXB6dZjKur4zYy01lfH5D+Rv6zAyP58Y3LlL2HQLL/Na3xGk4O
uc+Vxi7eSm2XBM3F9xsBF7ctHcCRKTClkO/74CZasarzHecRs31gxA/pBb9ZClst
0pPXYkGuaDWGO8Dmug9D3mBg2D+VtSmlF8wOJVU6ekWZrWGJOdSIaaO/PkqLyYZw
nLSKkyu02t8oNkVAwPewBZlwHDmHf3o6ru4c/N7x4YfoeWwen7Fv9jffgiLFzsBn
AuMAPn8F27FEMIDXhVR86dB3Ei6s/sONxcZSIn9ZzR1RdRwXGbnsl9+l7zXCVPuj
IkZaaJ3gMVrZL2OXvWnNL4Py+yPFpRf/tUNVYk47S83/zLX9YBc5uoudpZhNpeGQ
`protect END_PROTECTED
