`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3IJDar1RUPWU5HIQHxu9JzfvXsAVoywtQpa247GxYtwnGjR3QmZJzwjdLnErJjhs
znxInb/P1eU8YCSPs0LmZPt2eCT7oy72FycAGBLSLTk9VGlOJsAmPKwGuFX6OSVg
QK1ZNhBVh2bQ7z/sHSYIwMAAJpdgcEkODOHhdfwSZ5RE7lZU0If0XU+tsYevCZpK
GcyybB+hLH/z+d9gRtuOxGE+AMTPD8gPl2L/qnrOvtqZGdIubjHOHDOtryBfPBKo
MtzDp6ozQ+/wX2Eo2AsY45uEmOayE/9AFPazoYEpk90mqMRAsYNznesrma3VubHV
ik9/47m/lJXc6HCky3PDK2a4zyojrLCcUOSj5t+EdqlVf8qtr/Xrudy5wLsQ7azY
QLvpalafXg5oR5+paHemH5WhCOsM+rSB16NJoN4HYf/FIAy+qcPOlTWQYT4ahDXI
hE34zu3ocuHk+ib573CBtKZn8zh6UWMngJ4K5F4CfMy75vHTYaK7TBLzIFJafVkT
pVZtV8FHaF3CpqWflGNlKDlStiXPop9fClavqxW1WFcIhwhySI/3X85szMYh4eu4
qVyf1nHYmPofLOA+QZrIIK2EyWOArsWkbxXfxLYBXii6BxqL5k+5gvaslCKzlRmh
k+RjRuruwp6sbEQ7G1yPBPJWhoyaTu2dLAxg4p6z9njhxmBOLZpqx4PCk9puvWbK
wRyfnj/OGnni03JF755Gu9Q96FF/cmRkzeLjqMyMTEnHASon9a+hsbTihh7BwKxQ
p8ikzZTPABBp4juLj4CBk+VJoI5f8xDtQoToUAUVThEo+AlU1a5/3T5brrLzposT
wpNv7j+OaZTEqJo4xuLlM3XhVvNq2whvSpGyxn8E/yfKtSForXoxW2UE8W72mjwj
/n/UbAEL1bHSBNj5hwUkhxC8xtXHlsjyotuxkK9sNGahhUrW3Q12rStOlN+L54yC
5fNO6e+E9Op7AJDhEaOdVhIHcxlSMaHnW4uSkC1FgFfNyvCPHKtWTIwPuFvJZE0b
WSLOQTWkGFYg1Jrrr0lsJvQg++pLkK4wg+reEIpQZPH9doImTOIHbt6e7lHsoIab
ZBREajMEsz3/KwYOlopySQ==
`protect END_PROTECTED
