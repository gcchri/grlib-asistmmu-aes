`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wPPz3+QMktGw5blhiS6i0AucMcGa9rJDO0pHPAqPMDC8PtcETJ8qeaytUerzwody
od+sjx53fvWDGcsFTmmsB+pCGYNR19P+RbNKKZVd8/SCYjDxVqIgrCt26TMSsKF9
jvE0wC+5DPZkJDemLxYRJ5aRwpQ3wF023A2jwrSAKWCNwv90cPddzBY7nycn8vWb
umnGoaiAVnMlMMRp3IDDVsUdoenTp9Xrlxu5KgJO2KTZJiBcogcwzVtR/ewYVIOR
4Q0+NSX6aTTDjby4BkcgkLxWYgAPySw1b4K3SAZItp+HoXoNU/RuAu6rU0GXD2hj
M3dFCfBfxFBsV4OPqoTCbFCc9HiBrasSo9kQmEVD2iX6Y4ZFP4NkMMzTsHua3tt0
sCPth+3vzEjLQiX+XZTuNd3RJiEPXCRORaU7uvSi8ToiSgST9tRFuF9Ihxo5ijIr
1kGEZ1cDAoBiAWuKpCigyjLTEGhIJhCmtwUcGQOuklxOk34OwrJ2lLuA0U3mtlYc
uY+hAYsz4ppMZ+U99W6Gxm3P62tDxIuukTP1l7lv9cAX9LNqW6DNZGEll4PUlpwR
GNqQNYOpRx2wZ7zZM/WB7Vm6F9ftfC9Thx9uMMSsKSrSg4MRW6s20J7Dto/pQw3r
KuVmsS0T1UoKvy2/00S/wzNoPQcgf1iBWO84Kg76cw2ICfv2jqprsEffY4L84hSB
xNtDjrx4D80SqgpzzHuUglEbza5GE/iGerDB67jci1NZHLB2X150eKbyNg54jDEg
yXH+mKDj7vj4NZaA5Jx6GPjS4xaNAVbCZLAPKkO++ChhzLhwMtbVM4eDVdmTIAPl
IQ7Obtorz1pxyx4cjZO4R2oLRusmuPPstmCDh04WBQYYn4vXydcTKoQXxZr04lGS
rk8k9XIcDuKXNVWm6RzQiHUUu5TrHYj2kycpSZwAf7p5SvDFHydEfR0gjjXceUUR
pSPH5f2gXk0zy4FicPUxkOa+a0IzvOXji/ywfzP08tHcoJToTXgW2ZiXv9OP+9nN
U+HaXzdrzQIbmHzH6rvKc0d6FIco2t//1uBNnTd+F8jQbbb3iati/glJfgw3smuQ
lBvSAvUyxzQ0ZTCMnJxOfQAqKs134b+VQ18L7SXxhX6Np0fRxOL/h1g4H6SSETWv
euS56vM/C3oDDZxSLH5wlA0soVgxMo0myfZ7P1dCuspRvQoLF95TCtlRAekdxwvt
W0x9QwjP7zon6nf2/7HndMsdZ5lHgXRJ4ZgxB8Hl84+fB1yBpDnXD7UJsWVRYeAt
6boO/YTJN0SoSaAW+3tlmMbRBJYlaikVwu1VpCfby8dniB5i70AedNP1G8AGoHWz
4ng3AFwLQVaqM/hOKi41bE1rTmSXW+kR7u4Ic3B46K2rIZ3lpBr4ZVCyl5BA+Meb
8FGUVmGAPKF375hR7iiaFj/lAeUwiBTU8+gUhGAJrVSBA4MnGPL3jTUEFyexi9cW
pSARb3f2OQjGyn9Xs5mBxRcWKYsFZyUNVuvMrFwdc/ja/3C5DpC4yjgOD+crUhVv
zhESqAXWcDmROqF0LVR4lcTt0ZbFbdBcF+WMWE//uXGufGdhJ2xdoE47PLE6jveR
DViqINwy/6WGGik4OcvAR4d5JUUkIkdnwSPFqjKMu8ivZgtPOLgaeoOKF1EKfMbE
/qvITPSJd8JEvB8OnOtmuDa2mGmcUsQAIughguo47LHHV5y/2CdSO09NRJ08AXm1
6FxmAjqmQSB62p8APIlGuUIfNzdZt9nFDCZg/jdHrHLbOC+pvvQrskt4hChdKHyN
I+cfusEYiwftP9e2+c3P/x7068jG74b4OyS50WKTna67CO2Y9ox3oPh0a/ftYtio
io07XcvHtVXA8REqqOHmx1rhMbRzyD/mx//OTpGz06lVzl10Y8sjPuHbFlnw8LdD
x6S5nkRCsBweTblN9a4pbINmFhoC1UYFMgDGd7gQPOCv3iXW5LORcGjqVAL/KiPv
KknLGN/v1DwMYl9uQi5itDNw5FOdvArrCDZjoiixvLsBwwjGPxOLZ1YV/Z9/1bjy
S3ZrM1ichQvYHslOGQdjAztWnCOPAZxRequ2PIv51AVuKrpiGykSKbkbeA8bVJbW
r4OxLTagUsJorFWj6wHaYwkHHEN4H5mHENI3/UWcmCX6cSNLwv91+NtBg8ziSeG/
+2hx1XjIe7qMjCioFA9TKV9QhuzIuXroNdDwNzBhbMbFJiORNdQvqZd2obALxloS
iW+OQEx4ZYlZy1t2f4NY2THKmf4tayTIQ6E+LhnhJUtxWuWrnfrWqQ6EjXyRtqKK
2XkEHvXGyJmUMtStFnHyQgIX2w6z2poGFGo+h2jIrVx77TreTxas+kTocSRK5E5k
WzA7I5ayIqmwixms7oMN+e8mkGJYq92XPaevREFtPlTSeZZejQK3kQXuPLuc1Q5Y
dk5uL26W+bB2Rec3kTlWR36ykTxdSD7amMvbgUF/6zwkfM5iJqSQNvT1Ve4oyVKr
PNyiPU1P1X3R14xqvqZCxzy2d4b/ETbC9N0cy+Mx8gUHJo3GAvPS4cDu377I2sWs
mMuhMrVmJFpQpfkwgDaUGl3UnuPKIfswIFl6lSisTlpcPLFfU30QcOlH74jEPF+8
SQA6/X38VFIJ05/vg3KD0ckriJFkOElk0cjgXrBRLaDARx3Z5WcqhnSfaSxpwJSa
zgy5Iir+/Ya3OQU41QVe/IFV0rVdDpoe2CDk84eUevjnbpcBFEJe7Yvs8tGMBnEF
Rrqrp8VuQgtqL8EClN1vMf4jUGDQOPA4uo//4hoM53KO9U+jjep19wnnMk0GXBdB
L/+7WQ8FxZVOOR1HsUwIGYKkX+DP9bIyfkrmlfX5C2sevQzmynUiBBXUx3+og47J
IWoHVxFiHW2uMRJM7ZjMu1XknVsa9GZanXk+dEbA73z0ya4ECjAbtgk8L1qGg2TC
BPpgUa+58HBVNqKjGGqDUYlDyWv0ieP7vvERlCEuHx0gshmy26t46EEV4Gp+CnT5
vW9phxYMXCT8QyClN9r37hRJLxfln3U6AYe4mUHyfz7NTpl/LtsslAqsFHTAT4f9
FVEXMkK1CdgycHYwRHbfyFx+zrHIXEUePjcdDmwfBcjTLoxMMTUmq6Q5xv0IOlvB
bQbNOVqOmnXHfCUvU3VYVUYd3MVV0rrdwmhEhUUM/cnNOL5DUmO3VGGNMcXoVLgJ
GNFaadNPltKytyLjtu49hCXnTCOOby6LFLhvmLZLHPi3zXL3G/SxS4fG7uniEZW5
Gnw9vU1U6wOd/z4Cagu42MNG9lp8vWpzRav1J9O3dcdze9RIl2cWJ1SKMyyCE913
fXySTAqwIwAVrRsYJEVgen7x0n8LgfrWJqX/FZ2YkovVEKx37EtLgXDZVpANRyxw
WJyvYVXQ/enA2Y4TI+GiZ3UFSZrKYKRgcPRTZKzF3Y4FHtQpvI5mffmTvLb3Jgp4
iAsezMa5q47+DZWuaqeSjtyhIBFpCE8egcR/JLg+PKunRt9Cb4g0W1gc4X1qMmqH
MJ3H3jv2AghDFCHMkwJ0CIhAHGhz5inl+q70aIthCpg/UszFonS9+9SGH9BHtJ3q
+GFYmd3lpjMM+wFxOmnlGchiRTcaBMXHK97SLSxeVcb3YrTU1rm/fgsVfTHacQhr
nLQNykhJD4pHu93diysbYH8bPbO3Ucqv/2ZLGNtwJfMFCQSMcD2pRtjAG3g1zFVK
c0w1/VPzzGi5PVl0hKllcpqayEGWY+ew7llqOuNMkAq9PpT2yqoeSJRT8Ar4R+DD
WMbfS4jkQeMNVGp4kfZdSrJCmHE8DV0VJQCMW3V8CSMK3VXyhrgkWeoweHly86FL
vJV8o0iET0qHJu3qVFslm58tAzRQvGkZNk0xfKW4u3Rci9f7vnobzshoWnAfkBdV
WEfRViJe8DJrsD52aX+vfjG6cIs8/L0//quMyxibel1xdFMcG8L45VT4HdrBxSO8
W/wI+6UPeRC3D694r9BZ3YhmshjNODReUQBBBxqrrvBaAtvHbAwPVPdp1GAi94vt
rZ/LFmRlAthOeqd9Fkrz2HbWwXUwmM1EA42E83Qj34EVgcPY42U2HgA/vcm7uUFc
wMbvjE3oU6E4RiUkS3oi04IjKEE9STvXz+/R6wAMvgugniRmZ3p6o9LrPOJ1njhf
H46qL8SmzglGYCGFZwMW9pDuF4K6sUV1Ysjn+teSH4qe4WzP7rgrBRx/nytTp0nk
tK/22XpfzRULJrPDZmiHIy5YmvCXBir1QwPWlM1/f7dDIYZRWFRMaLVVKmR3Lrz9
E4+ku7U2WbOUfh6bTeZ75Cs9SWNshwx7IsAVBCZbffirWvh3R5QHwZktUbJm/dNV
CNAJ962ZqmeMhpbRZfO1EtO7d27hycEbm6POBMhtRzDrSy4cmgB1fv4HBB0SnmtS
R/C/UncJtmQq3TVKTzNifrvJ2pf1wP9ND0dqaKqI2bYnznPhlVWlnL+ViEIVhJE3
N4EkA4e7iqB80p7gFWcv4z9JsD0veKbEpkhZ9mYJ2oL2GsTcXFDj5u+czzCa/p23
McCfWm1x3z4FcUEgYpN09xC9G5o4eEtAPIm/tiEW6KFH/GHpdQW6RiipHL0EszPv
kdCMmApTQZtvUrXL95+UKQbmDr7PKmfy6BYElVDkCCRksOjUmeIvr/n2+nLpK9HJ
tSaBPPz13m2Z975KNfZJ+EiHVHq5RZZ2E8ecr7OviORfBs9KZY0oLk4L/kf97abk
Nj+RsSANGSgv42frj7wCzkw9XNIpAn+Z6EvAPccotjaWoc2i2glAAPCbU0lx4t0Y
FgVL7ScDYN7pR2AY2mFg6axr9b0hl/IYqg1z+3Q0djRIBQ2VuaCxGDLKQ/4ySB0o
H6sFYclKrECYAwb39etuD4m+PhLy3g6ZhSmWQm8vsL1zjWxEEPcfCUPlWD2Aw3zS
x46taLjbPIHbbqOIiMg306TIQDEKtJLNjE8gUvx7o/NiCEHmFJTG5SYhuFAAEKmE
01QAnNQ3PKWO9vLlErfVPSIzN3UfSxZQQ1yIUJvJgR8Nve4zK3EXDsQZND4LKGne
jlk6ro653s9DxEeXuyItc4rmVTAeemqLwrp0sOrD909V/dZxWW7HAtbdGe8SvNws
9830b+g5tQSiAZKd7+BKvf4tmEaMtkm9fI9y52znnBrMnJ4jfmsS0O/UQ2Gf4ba2
DaTF0m2ubThzGMo7wOhiH29sxqsarOAiOSQoNc+OS5eM821sjtnlrxeXhDNV7h3u
404vUwfzcseoMTi28ALVLaUCWaBQdg5Y6gpObZPdflgunNQF9slHO/BcXUYTUDRB
kLckfp1vAMnrIfq7uHN+4PM4DpAReaZR1A9gkXbfUSKkihFMEyZH/NdFJ7/f5gT1
Z3NLDtwad13R+EbaMNa0GdmHpMsDpGwSlIwBDkqFJGFewEgr3hl8F/JQVGfH3wAP
B7kCciF7e4bV4MShiVGs93BzhMun7jCQ4mDEVg/FN+sCSIXt7KeDEZ0dIeUnY74u
GG/z3FLnK9QYyHlzhL5cQgjJlG0LvoArHMfZYmCbrxA=
`protect END_PROTECTED
