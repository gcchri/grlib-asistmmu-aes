`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/MjRlzzEMO4RmOvR3yJ6Zmn7M+4Aq+baduwqRhbYw8cd/hv0HiK/pBk52hJ9rUSG
4z4m7hxMMgyT3/cAbOxymJnpPnO/FrGf+1otWTjDAtUu4Rhx7gw3GusSIPx80jE0
nZ3yhozwcsT/CJeY5InIHy6qCSTxSOi4xAl8++SUMmo2OQIzeS8b9s4m1m2ubPA9
xFEW3z/7xebE3iNpEDfiNCkER5FQkNImyz0ejbCvKKb1zClcB/+BuigGq2ZUqhK1
tFkGGes1LA+XICcytOYIigy4JYY95TEaveYIUYWtWjbzAupfWzrgZF/MG3U71+Ux
mWe8HymUxu5b3J91cAtdbdwyIJl7aJ/DiVmkvhAYX62KnROnKbKHkY59WMMuCQhl
/35Omf4cE3sKtuywh9fu9Q==
`protect END_PROTECTED
