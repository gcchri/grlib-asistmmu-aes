`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZBFXnn6anDMPd77qBmQZ3q7/Q9h4H0YkRcIfIc6SbQq/LINjfn2B5FUBhu50dCMs
ICHkhd4zuSlNQJIjT1L3+8IG1iiVbN3NTNs2/qt9jkRScAX6eVDaZWJpfV6AB9wW
7rpHEyPliSQ24/2kI7EqMW4pmq6BXY6FLypUnUHw9CBgGvZcesoxODM73yOjE2SB
pKvMknDllhMGgDLl9hOFukZXK1MhN0ACFh+HL2bHn1OxMCdQ84VGCK8Vew+clSk1
SIG5Qc4IZqd/lWbxSJTS51h11bi1vWoSs2jVEPY9yDEQzaOoeRoDwXgTzmuX4OzD
/mfFo6SMAak0AdYUDxHs7FgrRb0HzIrUM6URJxc3YxYHmF2aYVQ9o+QgZ7bWRoYG
S/jU9vqriYRg/RpbdWSzE/8h42PMR7XorFkpck+ZMXe1FoIXf3MVA51Wa5wKbupT
e+y3qc5mk+/j8drWTK1wjQlE3PGXRcYm58KB8rG5WAlXLJHFjq9v6vQCf11dD4q6
l0duRyvCvNU7p8qETvi3QVbFvmKeRO8Y/2dFs5A907g6v0RcGr4CyNzxfwCSreG9
bhKLubIO21sV30RcomJHrIB2n+Dly3NUEiWkjwq3xh+0nn5gj3u+yEKv+jQ3kw6r
Yay8JOVzJiSzbIP0BLA6id+eEodQwpR+3/DIdHOajdEpMxtmZDIqjlXKbFXwEH+9
rha5789W0PEACVKbUCjw8qyFHrT7ri6w/Teta1Aqf9r+tfWAI+0V8r7Qyh4831EJ
XaSJHtW7aBNQX0PGSUeibvUeCFHVDHSr0ZjVjJZVizvrfDunYK/F9OBHb2nJwy8C
WuwdpLBVqoGjurimkiSJyRrZ1jNlhna8Y40ZvCVcJlh8touBenXN9EXZQnXOMiHt
LwYJywOvJC0BNIa6BqJEJZWGZFp7r0eyzbK9M4RW+5Ehbb8ydifXosYiin4ukcto
`protect END_PROTECTED
