`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pe2fuo1Kv4IGZhVrcDe1wzCabQ4Ut6H/c9NdEUDeqVwEaN4K4buMukkdicTrBuL0
+UALcKa/529Ct47lnMwAyfmNoSqwRgmG2APjxCWmHcExvENnDtk1Yaj7QjOHX7Xq
BQRQfbGDMH0Po9qqp7cvOVZEQKcSginP+aGGbx3YuPsVbiAzdt+IPWv4JOXQG/g3
oK04xGyxc6IyqrAn65rRltRESWfsgvjAWtNB47CwPzO6R89qa05rhS0oqv5teUYm
OL7r0mxHzdg887DJ0aqlNHbxmzP0Lu8W+IZl8Z5SEmSvRiukFaos2FkYhP8TF0I1
VH3BHRP3vQ4EnDX9d5dAE6umTEo1BorSkURHJagaih2C0MIJLZE8c5UrlsyTF5i4
0pzAnd6/JCH+KBeL1p1zsC5PKyJ7culFAzcT1F6tk5j7LKtDC2Sy7Gd2IwAv2Lkr
S+COEBMiNmysLBFGNro2ZjAMf38CYroCMIWrzMVnYq3KaPohvtdq/KjPKC6FlYB1
J7KeHY7jHVE/AV8kJhAljZ4WzO3u/veiAvY++MguVAqiKxaD0ZtHTmuQz3J9c9VZ
S2HlQxMG70+pMU1MFpVAC8AAXajHoZNGeYMRPd1RvYP4QIrAlIfpl0Ry7V1SJrOd
h9amnbM1rzkf5vfM0f9jGNJSWF6iBkVmX4dV5Fk6ujHHAgYpgbwtZ8cAUZnk2wAd
dDy7il8vCxCxTbtEFxpDJxMDyBN9kZnQbpdOxjUCARsjGlEa7k7KQkgZm65zIqbd
lS9tufWH5hvtCNNDhxbRa+yhMxaOo+JAQ+kQGAaSSvD5VncMgQqtA2x8KBB/ngrc
yQnebb0drbaTJRQR0Q2vfG/8Euj7ta/rHUC5hRCc26QoGvJmFKDIh9zO7bQpkkzm
9CqWg4Bentm27FSfoo2pJETeEGtaVq1sb270R/fkZl4RFmr0Frcw+imTvBfsfzpL
qOhz9839zbIIykvSDU2CcYP5ChqgYeGH30YlDLxcktectbWWyDssYnesTRAzX3h8
7xnBqCLyjO1TNo2lTVCx2QmfTRg2hJiXgFp3/GlebZ3oBXew+297bH+HHsxbz+MA
A6KQlP1Kzugebb5uVmdob9oC8D7z4+23SHDqh1e+CXO/OLQzx8d+znZcSpukqsGa
lRwX0fdDJ9b/Hhknt0TgUBoM+jvxPvkwrD5dOVBtp4XYEtGK3jn7+j83FvbM8Wae
/ioNItQUhELAjEUY+pQ2OOkget2MuV25PsW7w+hXugpdced5X6KnmylAhqUvwe6B
RbrCDKX7klcDKS+tPD3jjPEJPfkyhw+/BXqWDHT1Jn36ZaLx00lFFmExQztEjPv5
XStzu/V8B9v21SxFrNSXsiMbYw3GgW/btMYKuuTB7iVMP39u4+WoxjosqZfPZCVN
NWOMBwe9IkTIbiod9aqT4jAwFj5HndI9Fl0RCkXxFIw0VEniilfFsqP6SoqRDvCO
7djFb2x6D2/G0lnEviulgubJ2qqam/8D31otMjt8A+fyDy4cqVB9hh/s0SB8ZOK3
7Y/zx01ZZZ+qSdSmkzjbiG9JlNaCiBsOn8iyZip1we0gFGHZmTWO5ZaD2ykMgabv
kuyLhJQqc5sMI5YMnY1uzVjaGCoDQAROfTRa8T0iv8y0tflcKX0nKft9xNqnbkQN
WHJfc9Hf9TAU39YpxPx7mqDk6dnQyu1+kxTdW9q4epGWcwrLZIKGLac5M8YBmwyc
TNoqmLoghpbEe1gSuKOVUXeYDvMDe1ofxAux5eEn+CbCjPHPtPmUUMLIEQGciePF
7u9iFjF11qlnmGr63/vocpwfXQ+YqLOZtlsujsMHtYBoAOoYvXm6ZVezGkCKmTWO
ev/9oSv37hkiLABHlsgLefvS9ob+lkUh3nF3OFgEtZgy4XZz3nKbLMwW6LnKIpAg
UNZS+G/cOHgXY3D5w0KBGBESJ5ZMZcxT2KpSIZjVqD98S6cfY+8aBp8KwGy4PFCY
nJH5Hfv7ntSnz1NZUObHe/+Hrxaiosot8YzRd9gIUHHlee5/46O6RG5ArUZkcuXN
y1uZUe+cmTwVhpTFEGYKe2+kgLC5c3xQsSeMWlokFqdpw2d7siVKvgR2r8mtJAPR
fXmWtE7dMGWVQbFj//y3yjPllofld/NaH3/TTlX3DOpgMRTCTaI2bcKcD4q598nb
LgkwCDWMPWRbht+2Pd6dzOSIlwh0Is6msCdFmqlMRl6d/LaF5rwiLyqmxwEcnI3r
oDS2hq783NGNvQsPEtsQGUCGu08ZfE7zgFl44rUD8tUlwUH0Iuq9Vt8EOu6zHL18
0zNZPXyTXWbu2zquaA8kJ3zU0OnE454gKEoACP8ypeouFM7PC+YnjzOi9GSXJw+o
9NqFWgN2A+gkUW5BWrD1uGOBJka5xwgm8SsDbWtTC+UReAs9NszBBh/PV8JxlF1O
S0EB3sGJs5D0ozHOnFXInQXSElYwvvus3QOVk09i1X6qL/H2GKXqtX3q2fXSGGR8
M/QOe7A1BZ6d44oL+n7M3lDL/zT2ijBclcjkoJT9/8a1ejCy7V3xNvF6FkniWfle
BvAeY82EOnzfuoLKLMU7mpGDZPhPm/ZypIvzFQt9MPLPQcvEElVwafP2s4Lu9PNP
`protect END_PROTECTED
