`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
82+3jNI0KVY2ZH4gmSFqkJqPkstrXOYTpXWZwdsnjW8TCC+SsvhlhQDE+wGCHEQ9
+BBm2efDt6NmK/tWzrtYW7gxxZyhpKdS0T0wramTT4B+G3IxG5OyVSj9+SGllMJp
dJOfCSiKDRDqkOmbSLsk/qY++c6BOkM6OlFQZhxoZChojZfaxbO/5ZEJiL5Qo4za
YjcxYo8X42Poa1DNtrGX8B42ErlLWWZ3fxNLKRCAL5ItLz3x2SkjeoTprsp+6g3C
M0BkgHGZDJgVMRfA2bJc++79uNGYCbvchUXsdQVaUYPpCVplAoveWaC531p74M8I
R7grUiZvLTaY95hgXDgYBA==
`protect END_PROTECTED
