`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ibMzomD6fWVWx815CMmNVZRRep0ElI7hOZSyQgFPVUBEwYTofsgIHOPLoFuDu9jU
jUiPQTTlhcyCpUneeml/Th15cEsYBG/n2H4ZoT+3n7jbDbdBxzI49cbPAbW1yDAA
D2fFZI6kJkx+wmIDkd9CeJXj4jpffsOQ7FXmGK7LUmnjsZl3rpikUexheEiwK4ba
r6j8tSN4ML5m04VEx4Axu9/zFYaTf5Tn7y5a6qa562NweEdaqgcrF9TJECE5yuNq
KMgJ04Xr/SfRTCDLLyOIxg==
`protect END_PROTECTED
