`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7FST9/5mKa2fLoUWDujDhDB45zHctpPMiF1FR/1JCPKC1hqmErU5L2tpgQGP3Hr3
oJMelVL0xSjVXhrsNfcECQEAaa8iSukcmy5WaLP9HKcMgcqtO9G/Ptx/eOV+C+1V
AnEqHcZIpfH3CZT1hIbSeUk+gSZalyGx8FmPqhMQKher/DfrHfoqhlVchaDkUCCI
xa4yRwdRZTPsmhyY1GUok1uKXJ+DnyfLYt36oVCWRenprkTumFZqwxVDU86IoPke
BMqtMxGdC2f1jvhgCgBJulrBBAqYrSA4+huGMonHtMl84MYts5tuxyzbYZtdUGP3
XC6ZBlXuju+kqYB2KeDFBlXbJWDlN5yq/rQKHD4Bwa2gBxRGx4BfQVJJqU3zuuid
uVi9x24qUmiTDg744ZICtcU5C62RV7aHoRPeQOsI8Os8PgTEOM/8LyUT80i+Ekk2
DX2l/4zxjs9Ksh4uDFnU1RVSdoegGKwGy9q755vwvG0qzudSs/h7184XvqKBUMTu
0P2PAC70RqFGS+2pS99Bp4OmvZ9OzyhURt4vLnEWt/HPFiyD8n2ESc+iu+Vum1RL
8BfPZL7qgNl4KylN5tVqhA==
`protect END_PROTECTED
