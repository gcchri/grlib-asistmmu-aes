`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zm8rdkYcCrBinPEDaIw/NaIFjJO0JfY0CJdyNOkRK4+rf5NS2kyoH999wBKAmh3C
AOJWxKHMbNgcqKhxbibY+3WRPK4PwTWy6lTbnsXynTWi5vwm3d/PTVjezc1gjEuX
OaXvJUGqZ6qT7SCevu7GhAzX0a77th0xucNlsrJOZof2em0zisP8keGHrSdeOM8y
Ri1gr5muHK5olhFg/drYR90Zj250smfY/nEH7Wlcoc1MCS/IaK2WFyYOJxKyf8L8
oeuEcGlFENGtVss6QEw2mgQtHsQPGmzIy+OGD5c7qWd+Im/azE4NIrJtDmmvc3Bk
OTplYCLBvMjVT2R60J7q4o2seEQjt87mdUPCBnSF+kWTiRI2W9ygzNxQ6HVTQOgP
zAI3mkNa+oiZUPilgvYODj1wVDjYUTNKzxQ4j5rqZ5pojqhkdMLwqKOkWPLatkk5
`protect END_PROTECTED
