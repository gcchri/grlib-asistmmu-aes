`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1OljQ06TJXH9pNOdTtO7hlxKt66tm544JtJttJvpehDe5j7qdd/0RZEOSG2lV846
zjLfFMHC6CWdnx05GnfBBnsT/bS7tMO9FYNakR5XaPwODQ2ir+ra7R+rJ2jHN0pL
HXdikVMYKCWna6xD+83WNV7FL3svzv0w5Y1XsR09FJQsvphtlbPI1w6BBqd3ydoc
EY8QAadJZgmKi7UnaxDkxFwWhz0py4lfRe7M6g17/QCEwKZY1J9qBp8VFicVsRQS
Izy+vu7+pHdqSJ5tZNgzcPy8sZ/rzG2TC/hoFnydTZbSCYjfwSfjUX/xbu/R69CO
SJHuIYu5FFLGf66Tpfqx3uTVEpWiMkDSQuG78f9zA/HZHfsQd5J4ei4bXJwsE6w5
7/WEBFgKafElC+HAk6IHylKnB271PMXW2u0vZOIyUFCyBUh/YvXVIurg+uly1j7q
Sq4hasJi+HzSYX1damw8iy1jlPmGau90pRncEq8scjLRQuhkTKejc5mqtPYnUiiz
Oh24hZKzhhnbXBNzeAA95qAO8wHkDL9giH5NQhGl23v1qcd9Df5XO8dvwgkqYRfE
hq9yVkPBjl98hMjuBKu153fRQlgmNTGVM20IFUUvDy+XSVermbPHdj4CjrSt3xYl
Gt6iEOW2eUcFE14hrjqvXOet8dqzLz1LnlIWTqMKaOhKcORPYSXJlfZ/kqG1eFRc
V5gGfqIQdmeMb1PaHs2B4hjlzIuQP1Gd5hT57MHwvrJ74z7hm9GL5vpk1ySyxfIR
r0jr2Voe8wgkmuKM/Zm61rItR+TJSI7Ch5tXMhs0nDlCwr7B8FYQ3HXnQqndftTr
opQYC5sa2EoAQ5aMrwRYJ0mFJyavD77pc/lSPly3GO82LSJRToivCsBP+19EZM3a
Lk6yRDr/A7aakBz+ZzwOgsZt5BN2GQEKvtKHLeFTYLbbs33H3ULcQ8tvsBHbC7VN
YJ3C8wVVBRpXFnpGVIBmYMxWsDvjkhCU7jJcL3N0Y4EJ9oHSLkz3BlsVyahMV5+x
nXA0PUeljDXzj8pGLbYQI6fca0clEcYFR+7LbK5ACg9vJOwKL/ByXJvqpN2z7CQV
UcCDgEY/wwmvfl8b61SrIij/hQvQkaeGqI39SyaqVAU7gqb2sFdoFG3AwyDvLCB+
3V5rj08oVBh1hz2Y5IdM9StAWOIMaDuJ/dT15aZB3tF0buWkgPXB9jrdvnmj1s/W
rZ7DEtPYE2gcSNvHfLzcC9O1LG49wvgVzGCdRlraOUo6zVHyQdJQgMUMKn+dTCLz
TyTS93Mono0/+PfZas8tG/OD3bwDRrih9+tjyKxwekzgByWR1YNdpQDEOgPJiONx
zUPvq/Rl1CtrKYhPRG0sxF2BFElxiGTGT4JJCuSys5EPEB02esIguYAS14Z97LK+
rxVbBWegByEfwPYdvc/eveM7j+Py51e6WMSju/yMATI8vvO9ABUQfIGw++r2DZBz
t8raJkh9vgFIIZqtIgSNCZIXkAfx0KM5lLPj/MDv/98bVw0MRUV0vK6FCKxTBCNK
Wmn9wns8aie5I4Izs4KrbHx0WwanW00Hg4ujnWibCaqcqi8RYN7Lnx7eqCbrUhDM
11SITOXxQu14SKJfTxNNDeP/Ivq2VnNeBAb/PEO+LafEcoPxKENfswFCyeImQz6H
uC67Keh5c0Bu8jquoEEtyHnQdgtZX2G+W2amagl3vh3Xo2xFeeZxd557xRN6KT6l
`protect END_PROTECTED
