`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8BJjbSDrxZHYAaV0jYa8pszy3FyHKgc9EKTnTtEfMOtjK6arx1OBK8aFv+yG1Ob7
eWcQDq2xPIfarpUuNKN/F8Nu/OSXPbgK6arKMoEmc8W3nVEu3V5gbtnXTcu9DxwO
olZezgDyLzjIJcB4K2nfX/yaKGX/qkmT/jm7bTsAjiKVJZp/uAoXachHbgQSp1sf
eN7nd+K6vY74t1WzY8LOXh+H1gIbv26qg82f5i/XfCzvOBgV4KU2EtL5ke4EERBO
XnTvL5pBHfzKj7Lw1wsYmftIxxBhDTUCwe9aGwfkNqdSjykiNRB3XGDULJAgqhOa
C4fV9+74TJZ1O+rtriUOAK+q/YTuo19SxBtyey8sqrSU0Wa1X53lTmjl1z+tTq7T
uTLTAdZHt4p1awNMsZ1a54AfVtprHoEe781F4oBMU2ntwGh5KG9tEG0WUI4Vuxkk
+dWe3aRXSgB0orfWrVCzgg==
`protect END_PROTECTED
