`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HsLZvyEc0BWGxCQG8vl+WTFuc7ympHAApQv3gaff8r266U04KUd99dDA3w7WwfEd
P4zRuUfSRCyPt0Atp+oU5bC4QQa1kvxGNMBGPwt8nXjINZlPVKW+NKCZMO/Z71mj
WRFnngCO1FAGaNek8uY++UxtkBn5HLsT86JX+trQe+7RUZYadEJMPjfoob6posU4
sDfVEDJktcmxSLsMW2Pt5BUFcFzi3eRVdw+ESHUohdxy5dylqtARofZn+8XsAIrB
lAqBohJ3lkNo0j56mWb2OA==
`protect END_PROTECTED
