`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EkW02P5ynD9sxcUTciPuSb+d6v9imJHJTscYpWVyNQ3va0ORURI/ag/e/49ZnGen
JrfYMkyFmhArnyUXsgx2hruNdvlpDb0rQsKpPmn2t+oLvPDGo+HlQeREvFFR3Dem
iV/hHE0uzaVvswvzagjq4DLKtKVvoWITJy10F2P1VM1O32a+xMt2UFgLRUTGSaQR
6tNRz8im6vm7WGh0MTs+yByoTlB87UiXdL72HzNhwQKkZ3/saSvcqJ2BI5u2QSvO
AW3bckdWhCkV0GXWzLenjgDJL8Kqq4pFXfF1Dtu7lSzWIia+m3eYgnz192bajM2H
DTiv9yW0N+uDBw8JgUUYGg==
`protect END_PROTECTED
