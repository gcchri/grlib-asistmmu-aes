`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2zJsrCZmeskN6KBwzBN8kTBysaCXM8wTzgZYMeLXEg6UkqQ63pGUDvf5qb5/Wewp
3LgzQa8h52ZMLceC0p1EQPqDcoeWy/HacOS3njf5HpDs7ZSk5nrjH1efX9yWgA0+
OMd+4Q0drycjLXXekS4KgkfqcDa2s9QOwWC+ZiMxskIok6KCBfsloVHJAMfzCCPQ
RAbGU/OUGJqP56688zQ8Y8ToH5lS7QpbjupIOdtSnaQnevdusGfEiE4N8qZV9b7V
rxlxnUdaWxgfTPWZcbMFQtdUfGD4RhuIy0iqBY3Xw8G50uTCaw9YT/Z7R5haJy6F
ByJAvN/wAnFjoUzW5MZOYLaDqPoExbsb9p97bAMfHZ9ypKOGsQBYWuZwDov0Fmk/
i27hLgxbMz6iEtZAonAqpe5EoKEuzP2YhFWvfgSGCcxYzKiloO29VIgjXG3uiugo
/is+R0m5C+qeZ0XZ/fAHzFxnXU8unZmTeewr2+s61KrIuHJuR1rINDDAdyS/o/uX
atH3N3at0POFEHNUx9n6VUs1gmbvj6NHNO0tcpAahf76nmgX8dnlAXVuxb4p2d5Q
sZNcU8uLDB0sMls3DmnM/m76aUSJXT+EYTZRd5EKdrsZwKJPK25QoydHSNyNN0pX
`protect END_PROTECTED
