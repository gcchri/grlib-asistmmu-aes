`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WeuUe2QfjCgTwtbuDyysnym3A2ZjvqVSLZUO3OBxSerwgg8LIL1bS2o5V8M9KfF8
1EpZcrqT841NIKYmfyVnxyCcZlBcH+3Ol/3/H6ljbX8+5e+8m877NGdi7oB63gbq
U6eBA33tAWbmel/TiZv8L0SlQtZVbSJjeT1v8m2zI0fb3sXOlnJhdNEsfXKr5pi3
OP8+qMSWY/QPKy7mfe40gJl5Bxdngsf2W1CySH6eyNtEutBB55sKMXDkUnv9Yk2A
qjqjvf4ry2NcRUY61YqcJ5A9LMtmCA1oPC+ZlT6cmJgu6RdwOQLRx812cueK7fm/
rTTHPBL/W27hbXkUnJ04jhZ9lyz1CvTyNPtckd3/u8C1bVQnrbig9N9W1GU9Z2Fg
+B5hNTAARF1UyLqHYnIvpvsFzwr4NkWKS6BCt1/JloNnBQvZW+SugWO6b0PxO+6c
Z9T/OidaPyvKzH5gKKfEEfXgBXMTRkSUXTnpsZF9hYyKTVWp4fjpgj2D9CtCG4YA
5lFy+Iq9mbFjL/NXMGoALowpdb9aG2M5TNxONzshYLSBQ5VyhgLJjS0cDt5jrPKL
31JjdsCZSKtM5iLMirqVtAqZMM23LZQMEWylpRfyxp4J2kP+ZAEh2vXISPEx2LLX
AvIfWqOpKVZdN5o4jvDacS7RgSBhlH/vaNE9ZCnUD+DhngET5luTCJQGq9etuC4Z
BhmSw6iDTBhYJwyzJtMJAy3IhWGXLDJ4QbVRyvd72ZfxYox9AY0DH8hSoybyHmB2
153P6thalVKeodbB68B5JodDg/aMKmKTajhYUSg6gbTFyRGuJsONgVTUyZTp0/PI
QuvbTE/LnAJYcicDCPOH6JWeswUeciDYRtJVccCfZ57WYKaFyfSWXZ1HUJDyA7uw
`protect END_PROTECTED
