`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dzzb0P0npdlgxNKrGLJjZFxu84U3eAW3ztPp/mrlt+k54mP2qbKxav1Y6YNPpd/K
cJbJjlUoWAYY/DO8Nr6KkBZZEmpKKoBPWp9hrrkK/6VTdcPYFuqZGtzGvGuHLt98
MgtwFe8bg6fz92IvLzGKZ22c5CGcQYMFiWrmOpFXKm41OmEl1HFMOJLf7KBHm6/0
lfrxz4zM/BbdhPfpvDvXx1KH/yWexNdms2lw0D/QsfCB6HmWQY5AxlUsySt4h3iF
dhPF067gvZVi+Yp+R/PNKPUJ3y2KV6fLNhgF7mmBgot5Su0h67FNVqTXAN6ACkUX
z7fTEPQMeGD4q4N6M9vPW4J/j1G1GDXMkH+R4WmwvieE0zJQSmUzfCfSonHbvn53
qHFPVx2tAZqlVeYp7AOWdFdAlemLtygNH0z8tDdkHeDOX+fOoYTYIYs2DnOqdP8P
6o5frd6na7fd0ocrJF2zAQk3NES1cct8CFeiHIRnnNufou8Hgd2ffv9lwWPh6mfF
/EGpOJXIQ4yOojSlWVTdgWReE+RZUhCkyQGTAP/JSxSOvAosmGuA1TkvH8HLhozj
vF+bKamfAh/yDIZvyWE0xDHnopSWWvbFeBoaChyIBeljoL9RlpcOrDAY1n68vXPY
oM6ksYlq120lh2rG5tk9ZQ==
`protect END_PROTECTED
