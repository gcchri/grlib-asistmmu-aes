`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3b9XXB6TNyTKd70KiAVjfNTaBKyojaD3xaEBdrVNJ2CrlzvOqWJ5XXu+pv553NNR
Cs5vctonWke46Pt08aFLjm0wxXdY6t/g62ITD/0ZvnoPomi+5GsAJXeJwovJGfCh
Tu1KwwEuthWCwW10R4JXXc/21kGLTj7JCyZ3TQi6jgJY6xNLMfTq7ugaZxKoSErc
Bt0HGJLiehsdQ8O0gzVSvCDq85bgAmRg6EBzkuuoydSPgU9ZqMzJyX0PBEJzhiOi
`protect END_PROTECTED
