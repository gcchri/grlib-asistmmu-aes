`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ci6BJJWBvWEXh60Gg5vXm+SFmXiN8pFDUf3TKll3aOsFK0mGlbZRVPvfUitVaq7U
r27WYpKrgR9HazOfQpvkx9Sj8Fb6fBo2SqnwW152RMwd/DJbmqsygWznJsjE61PL
t1f0TdaWpdifx67S1ZrM0rOBTIT7VRDFg6PgNzQFXCLlJCcOuUcLbA9AgkuVY5FO
tJMa34ebbT3XJA6sKARDfIbC+LKn4ZCEwvwBL/e4MALfIwD0oOdqECm55kkY/s9t
wBZ47+cOlpkGIK/Ii/lkqZb0WFbZNhIOjr1V7MXKYluOurWhgnoPupsaWY+nVD6H
Iu8yDKNr3U+0le8ARna0OvLuwUqGhzhNtJGkUk7Jzg3XZoXU62aqpQcyFE4nS3vy
+4YB3L2nFaKSb4SjsY21a/3GEeMkv4DSkOcO8yMb2FVdEfxjuVlZhfKy2zpnlcV/
r/Iw8h8rQHKL+Y6Xg2pRRVksnBa83Eguz/locByGhE3msV35wwldFm/ZVlNM7drB
n4WSJA2Q7oHalqnw5/m6nk9sNpdCq7D7aJ2/vroBQIt64hHv7xoXkORoMXqP3JtW
PlvFDhpZ9rVhjrHkXv8Q3l3Pquz1+5pQWaSE6tOE6kSKdM4z+Zc2000CITN45fsw
jJva4LrQ++2bjEzWM7PGo2YJJxBXmgiI5dABNGCMLyaZ9mF1/LeyXWj5EZFwR0dt
zlGaDb6Nf3qW5WSxPq2eP+E6aQSeF9EOpIy6F2/xf/3AOCe6umJP0RglqfnLXH5E
ag+YvhF8Q+/BCprBGksfcpx2v1INXPSYSq+0p0+peHZQ2U1xJvPJPIht6ZF60LI/
iz2F/FUxV5Gpwd2e+P70CMlKJ+4y3bTKx+NPBPgInL8=
`protect END_PROTECTED
