`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l5z6g26te89CMmAEy9Txu9vWdBvAYyDkfYiZ5PzH+tWFHi9/WRWZRYZV61VzK9Jk
5RFovDPSkf1s2i9rJB0ZkXca160HeKvDU+R3YciKT3JDQ1/ghHBgU+voRItUcquA
tlVf99l80u2M8sREVoGad+lhNsFXdvcNOfg0ely3BfuQ56waKkxnVQHOeSdrUJTV
nkJkKkMklX2zlLAWWJxSaAwtHomJUEtsTOxWy9Aw6TGkBgAJRBdC3MG0/9RK+3c+
wO/DS/hZpEZd+27JNomz6bCsAKc1jKlHZn3jqbEp4VPIPQC+BaomiaBdAttNjUg9
uRsFD0IU9jc0uGMqsdy6G/TOW+Kp/jj3aNYChUwnRdABJ96jVbOIB1L/3ancQuqc
1t1/lpQ/Ks0s4EFqjSR/dwHONt5TCSwC+ZzyO2Ikp+kbhrI5RAiMqlklo7lx2tvg
cgUGy+3+J8tBrt+WL2wLVgjc97z4LsVS4UoTM+sVfaCk5jcy8JpeHRXQyAQs+cqp
5kZmHc7KzcPhuALNP1degsmej5SmMzQYyNQ8reMB1JZnOLHikZboPRWuUUlXisJN
D2kvS0uQMz1pJF4WWEnVmVGPD41NOGZUoOCUvpTOttDR+0IPa3wnNWhcFI80338a
nJCLklHm5KT6oRY0jlU3z17Hi8ahmHwuHAcAA3mbVQISSPnGd1QvN9LvlZGx1VE5
vlSF0tZVQZdgHjD8ncBEjNsBIjitVR/Svrr/kVP9FtEAcIz0C1J5VzkSurEguJwg
SyneEu7pXAENl0o/C8aA1yHtlDkeQS7rhzks+g5yXKaQdkcR6A375xdco8TR7b9h
YhhJeGcaTXSKoe3DOmXT4GUhijDVqgegMbguWuiYJ+gBRqql3/n9bPIMOdUOlra+
Fn2BAM2em+zzZUPTTnb8LdXSq4VQWT60/6sm33A2fqYwkT44rP1EGKDe/FxVEbcG
6OtJmtaa5wGrDgF9ZW/hwdoCv0Ej+1vERfSY0jfOHB8W/Kuy9teMFcN6/IkNEKj7
ye8BWoCImeUDLbdhZ1FRGSfnWvUHJx2EVmINObwZWXnmKLC6kSao+jQMLTr6tuVr
IcTwgUQBtgEXeMnL9VzeuL8zqb9aEPpl+qL9mCh05I8dPJ+aE0wM3+pPKubdUuwV
m4wwlE6WUrk12wKJxXtbxbW/RTXsJqQquREGRi3QvqBjIjh3D+txpjNE0h6doDla
0m6pzVbkj2xGbtXSgp7DRkhjC/RzmChsLjqpMNCKw74/z2LpjdokAZScPJ/s92AZ
Of83anvSoq3L2ns0XkQnsL95cG9ab8EmSkvNz60s7/Nab/DUCO2EBkSoIsNDpKmC
ZqNGG122ojq1F9E7SNB6AbMQ1kVGKxValwU5AtVjs/AzCTf/VD6FMwupqoiaibOu
YbtX8t8egvHByww/4ycJEsi/ltsnpcrNcqaUjrXGJsvNxBQmmR6sBkGatT2J3DoW
rKoMFlgw4fEl0ZsFlmvBem/4ItshzWtum9d29c6TK5d1Vr0tUG4PnqZizzFeC7Si
cGDn6yfdH6+HcTnMcerWSOsTDv2DOgMZT9E7tuwmIletrEYakUT0MJHphSo40Kr0
qL+CTd03m92fqImHLmzf2Rgy5qd6j12hHA2KUZhDHkMdcntjnGc3sbjEG9JlLWJY
NnWoDiqmAKFPzihKrR16Nn65nb4ezuzaCX9YvrHlMCan1TJMM54opR/kG7FCogEP
4zXOmqus3gZp7hYZcChkOClZPyHFIqlJy2qiYqA/o8efb6z1BBz88WMXcZqmOc+W
f7MmM9Liv3PS/OxVB66oax9fE6zllutfwUM2ElyNivZwhzp7gqvsSBL5eo3wFpUW
JkeWM8kWzBCYqP9rkfD+dP7L4xbPLtRQijKrBrS5xBYT3L29gJ47ElVQcJIGIa36
rJoF3E6/1JQiIUvPPzHQFNmPHqQFzzRXyogKkeWN/t3Ml2+m5qbO8iVqAghBxslg
8pmQxyCuV8LNYghuOeAd42f10AP9DTmOn8lGzxw+6kRrMQw/Fxxg3YBSjk0hK+lO
GlZQ2GFfroz/HW9RU7OZnKI4039WKZj3bAZ5vTRGv2rMDprKf94+ASBPBTADST10
wrdXFNWqMkKrQ86f08bq92A3Fko7Js6n9VO8lAqv/eadEU2JSaBimaaTAaZtSRoH
K/Rb+U1xBZBrfQWLrOp0XizY0qgWbVilhgCBplQbVSGclm08Ql8Ut+k4fumXA89s
ZGTAlV3TV2LakOXmWLO85RtwLtEr4z2CYfRo53x2N2lNkQhG2zkCqASp7zIkdEfZ
Rgp7eX2IBUq+dk/0GD99GyWDtv/74Rfjdj4hUF01EszXQapx6jH4spgT8ZOwEcds
/4t/5yOC/iijSdTgcfuj2k7BLYbjCQm8Xc0A5Ucdn0rB1SKcmO8apXUOcg6dqX3B
AF463JPrx1xhdRqcrmzb6eT6Sza+znUd7t6zgHkA+htMPVCcAfJCV11W+bX/rsqX
ppfJYOqlvveTSCG0S7jmj9C0LujAb78LXGaiFaxpEzkzpE1jfmZXGuxLFLPB+tWl
RNHUlaUqp4BMbE3cCOZNtbWmBP1KBiQ08ZSMkyg8SraxXZW+xjYQzaN7zZOHoHhS
np/hji5eb31sKXDE9l27GrQQJ7BDb0ucTuSQ9lzxQHucdSFU5MBDbBGyhKAIe83Q
lQfy9EW8QyrOgARE1W+ei4MVSqdzDkkPIqi5F0a/eelEEM93RAcDB5UW/qVGD9jB
ajH3QJSkfQ9Xl9/QeStV9qLgrIk2Vb1YWkufNFoURu/Nevk6/pyhuErSOTyy98Gq
HyOuc62t+lOZMzl8c8ne/4f+fmsZd87sFtoDeF7+C5bg7bxdMNkesRyiKXmLvwld
703fsTOdBdGe1+qSubMgA7YEq7Mod/MKghiCpFuZnVqZG/BmuAlouHl2qm3bm6fF
H6FAqjeylhY9PiTYwvKC/Z5RdE4H5Cm985mTki0GoaHfJmoyLbfP8rjqUWFlKoHR
AEtF7I49EikSMjoCOIQwCTJiqtOra0zgxvo7Z/3Mqu//IGHR8bhm42ZRLYA7yptU
gVGuUKw/5unSXarGis51iIG9n1RsoLja9VqbC1Cb0aV/ztxvAifhliaBwQUEnQbZ
CFEMioMhXAgNMoDsHAoNhmRCenk1dI4Dwr/pUTYs85iDaI9Itm0/rMvhOWhvU4tn
bycXA5aWg9vwWLRbVzDqZHH7R9upEChCGsE4t4CH5ArER8pojsLpxa05wOcxriIT
+i5fwV0VBOnxf/pYPkIc82lQ/x3R3q99+iJWGh5YCth0Q8u0v8ve95DXagsApS8v
XdEcHIeY/8AsFn7sP/XM8DEllJqw83DAKySLT3+5ID+C6dlJjJ5TkFZfQmxIwLYl
aMy/MTt5ucd/PzyzrIglckG4U5xJYtUAHi3f5h5p8GZhPWgoulzdgl5Puy5zDRtD
l8TYa1rvuzsDbEvzwesCC7IMuSklfKG126XKwQCSm6AtV6gE1RkZuHZ3aaLWk8Ul
K1lGFEjl7+eBqQarIJmFlfP/XQQI0w4tPlvAtVMDqt160YyDHUpxFdvqCCZgxYkj
qdh/37HmlAE5UC8UXpfNgtXqhMOlZoTAyMUGLd3BI/3AimH4uanxuHLfPY9hO0iZ
RymoVOQVeF9/bs/GROaUV7orq9IHu25my6SnFwi2ooDXZp8e7oNTwWXEsUVBQpNS
ASLWJ9PUNxe6Lv1eIYrn+qhTmUXLjJ8KXYBz6sLR1ak=
`protect END_PROTECTED
