`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2116dDuBOoPgOXAguAL1/HyItq8opBbu1OXs9oO2rBl8ULVE9+gT+EWsSe3NRupZ
wbeTe/OXLxmbxy6hWceSsEtsfkQR5tYA6TUeJ8COqXwiBnpE+05aimFkuSnA4KmB
KTP9dufJm2AsN7Xdkohs6jQmpfZl/LRGFHXKEvYyxerJwXEMI7r7RVGFr52FnBlA
1L5Bvg3hNlOVTpNKpu35ANnEbhdFV31hvIjESJyUga1JNkverqiSuHcK9sMcjhfK
CoMQkUfBN/0H/BWDpsWEkoybrx01iUJ7MeWxHxWHIYM3VMz7PfAJUk3xc9wINwht
rr7dA8e6WbxTm5Ktt8oljYn4+WN+3jrNmvdJLlS8sEN6OczoS6UsuNsrxYUjE13M
2ViNoqK3+vp66PZM7OytXiYzNjafXSry7HyjZiQCk25HUPt8279Kgu9XEH75+o00
`protect END_PROTECTED
