`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mSeJZJ9isBT5LsOuBS7RTt4TnPRphe6LzD6sUslqfQihaN0a8BE6NnDCPIsNbQnE
G5RRM5qbiHmBUwNotj857cxXMTmIQR0TnGHnZYNTWAO0FC3UHsjlydHnk4zROqcp
tMB445dd9//ltKRcflrQ52Y+JjbUIpAL3aH5L8JOOFFwrkoG3l4kLOUM3AMcGwic
kBgQMYpR1bxHabsd2Vf3pL+jJ7zR0eras81rNdhX0tZAurNpW2nRFwas5jVyYY3A
efZluognupYo1Gf79K9Z29bkhkm6qua0lp0/dD892upKCEDEZrW7aFLwLr/TF4a8
QzmDc0PUTHMOf9q6nORKnpXcpgaTKZO13KnEiofnhZ/wPmoeE4G4YFImILF7YgnR
CVYylwBmrKBuapnyKqoXVZ6ch2EUfRVDEwMgSD2DDkMTKDtKTDKd0K3TWxhzkyRk
`protect END_PROTECTED
