`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3t3k/7dgnMbicIn3LePO1C69U/mvgwU7d0XAU2L9nt1Xryloq/5+H3XTMs+szAvn
k5TyfWd3xMBjNAKNPyl2vgaVywyBrWkB+dVufry4F9jheFnpjqVeHNxClFuiSuuL
bTwzHdOsOT6LoesEey0nWGC49CaC63Q1KRvySTH8RSUHZ+WFk0aMrCF4BhM8HV5N
chX7vuH4wqOID3j23yaHPjbyfbYoswDicocOAYkSkwrRZ7i7/KpPoqO6eXjzYT86
mYAM17V2w5XTFtNWLACCLmKYm3w+bY/pjCiLGAlZHzx3rT6FvApGDOAwxf0ayhIT
D2U4YxBPR2+yt7x3PsWX1Srpb7fFB5vMq8/sI6IfbY1tLv+Eg3OmWA95ym+Y4p1f
UA7y+hizqnputly/H9bz07GFO+ETmeu+3s8ASB6ZTFYv/KPeIk0cbvURCZ6qjmi6
LTmnALeinmxuqUZImbg2t+zPmU4+qpmG06WdW1CigQPIF0DajjbHNCn5ARa9ioox
3oOFL6j/ampqselbdoWcc6wH+hz73CpiyE8kLVDKwi599t7ukMzpgZTOAmq9IgeU
wEp8+kDtC1voLo5J5J7DVC462IAvzHcD5XoeBkXZcKV6gJEIovct+dmx9kzUbgyM
sVozQzc9hJXzZVwusQO/o9A+8L8vmLcgOM0upYoHtLXAGaYfUSZ+aZ4vLXDtxKmw
mMY/ph6VuApyjxlvrIzXstaEjIlHXHMFsU5euhEQOsuTht6y/V9EkVNQ9WVFrBNz
LfgWaej/2vnoLN+HQ3cb4ZrV1taWdvAQaF+Uc635xO03M7uMr6X0UeXT2CFKROTs
iSmhphwjnD85z/jIYGTXIqwMUmX9pZiRbcZuCTy97xOXc2ilh+onut9F93D1yosW
gfUbTq8V6pMukIi/tXKbbsk050+awt8Dg8oQf9azjwUTNCtQ8+CsOsb+1ZG5dGMn
8Y4Onv7gcTR7KNJnDZoJ1XLLSGhJr5PtWg2A349ed9qXyCJCeE+6cQUbHnHrJTzi
/PdqEh5ThXORpGhF2M4DfTmVtUbR1zakwERf+sKQs/VB6CjL5f8wDgQG8dOrtrTH
U5RNvOXfyZlTZYn64I0Z39I9vl6gwhyckBLJKhn4/5lKVMuw2WrkoK69KddaKu29
gzUksAX4FhZo22JLmKvxMAiFPS0qUNCTRHzJT3czaPoJA3do04WW1bd1nWa0Q1Dc
ce4NcXD4tD3lh32w6l3gl0TVE30oNbi1V+yr4sWEXcyPZPzcZX8P4WIbdIH+6B6S
FJzWQr7U2uULTxKkGpGZYO9Gj5ISZRiPrWKmcFqnFjbE9z4Zp6NTrga+/ErwkWmV
etkewAzR8BLHfQME1ICdnrojCeqBSySjx587kTD5AgaC2HXWLnTmZiv6yKJybUqm
pfgL347KoGVURykGGrUM3P6Vw8REgyMic7Ql03UZU55IKiU/zQihK4x1eOFuTVTw
h+m2Vek7kqFjsSOdYiNXNvGQG2KUK9w+82sO0dOLZC8VJBxotfD8Vqsqp9LubKfD
3V/STtewf+0s2KQT/KAoXNHidkEpovQnZ5PN47r9wCQm0/gcrjux0LmIGp01nDdd
g1iUXvdZPog+PGw0KR/TQQBHVXr8IE6T98T+rNW1tFTOUAne6bSme9PGn6121BxT
G5WBI+B2eG4FWrOZzxk8kaLa1UkpZEpyKDce1Vv7iGCI/CcVO3nucuA/PuPwYzkF
NmcQcu760fZBudhjJDMNSRGN/3m2AgpoMef3+q5X6mBk+f244qE9x349CVHokZM9
LPSBys8m50s7u0N1SpmmUXlk6JAY7bqf713oNB6Miz2Gqtl+/hPj2IcBayMY5qJ+
aKphuFGT6zxk/MEJJGKJpJgtdd9FNjJptUewK6oJVCI/2ucGg2uJ4yctVqh/p9/J
Tk/hkVqCASyW696nPByiirBaeuI00tPFFV0WDDeqPX/PbXNGkCVxMW9tKE1xvOqy
4EMT34m4amoCC6HS6Dv8fv/skRUu0b0cjY/ecM/JYG6c1NDZDypht//3xfHn9SuM
QpI6m45Qo2StAUY4PnyHE8lgzI+Omo+2CnvmSzUxFPPbrD5p4AV+t+uqWoUP8imu
cUN8D8dlM+ktLVOzohieHaicjRoOf/isN0d3cnfYB+VlCgnSMibFYesA8yHTqC3Y
Ap2npmFSdo54EPFCysgbJMMRNjbnulPH0lCbbYnVKJHTbIiFOS5LrSCLtTnDjM0B
zgWb+qFx9fiKnMfDRi04wlKG6/X1EDtlkK5+VY70NPrJA9LU6vuD0C1sHuowMyDi
LDNUsWR9kgbHo+vgNOpJnNJ+ORyONBlv06v8ITZNboG5MtWCgOrf8Eaj6L00r9c1
q7UijS+Fggmx6vPzwdGH8KemrN+IevW6hpu6pwV9nDWeyoCnpgd5koS5hv7zw615
/JoGJW5D0/dv9fJL0vHQoUhQOMnbvaZgTe4Pn2QszSLDzwtC8HJJDZaeBapaNGjB
nuEFLqc0UW7XLQqThlSLZyu+0y3yH/OTWFZYl5ZbBHQhBQXWlmMjUoKsP34+VV7w
CYC8IeHiMl4dtTzQRYKjwfpp/9E184cJmA/300XsFi1jh3fLALVuNX1xQzF41DaS
tkKDiNdgq7SjhTcDpkLHqenkBr+lhSqaPVd72z4aUALAs7QXMyAdM/Trq5YC74wF
0ihAyC1TTTEEJ6fI3sUZd+gUQ0a/aHp/27ZRdla/mc1lN88NzWzfl02gVCxSzwl1
yFJTCZiYlQ3Dfunxj7qzOsYZmXy3Pz80kjDOWoulzomL6E541p93+x+8evsDUCcy
rrUJptwHN+ij2CTy4zG0wOcrXSv5EbsTBnOQezCvAtxMO61Ab3QW3MviAJyMwObg
w9QVI9mw7CmqSq8aUQ9Cj7mYsNIAuRtQbDcImVZItJqiKnTJrhIxqZMqdx7XZK8B
OnRHVAe6ucfy4/nv0E+gZyQxgriaMITIirD1U27bUn1OXElgpa+5NsM97E2IjJlX
F0/L3PWBPTntUnSc9byr6HL+/dExWP4jiizXdy7QidIXx9S3O6N0TGWn/8sQTNRQ
0/GJqeKt4XYX6SK73Ad+TxRAB8N2pNt+suGwYizk1xYTwndXwDLErjZNmKdCMWJY
9gT3+iFD6cA8Ui3fXJDFRlReX1snppfFP1dTmcTu30GsSlA1/4VGPtP+HdLX5iOw
6YJP+uNNGBt7l7jTngCUqpAlTLWYaY6l9x+Jm4/3SeiyaWEZd95klEfpRxeAQS5S
oPnC0afp9HfLe5Ux7WBvaS1BenL2qOm2/mTcVlaGnIHYh1EmCrXUYSlGIrkQyQvz
LZ8ANnwFC4kdfno7S1uRO+i5jKGkKam/9SBz4xW7k/01oZnWp94PvuD3uU8OnRtI
jhuBUjhZH6kw/AeH0oGUCsWoiNyAnEWhiIaFsSqrF2qDEgNOndPRvtl41FSEcEtY
anVrvwyGr6a83g06Fr1eJ5R2TPlxSkp75t0M3gAuR24lRT2FJLUkAO5BeF7Wzx+X
ediiiHVCLeuqikM47rWbVJppukwxDA1GscY6LYghObAYrz2YjpBdHR4MQ7z3gGhD
MK5Av9by0/LchEmbKUhvz5SQfDnxFEtES+ZL0N58Mif7OYtWwSgyfOruc/J9VIXG
J/I5zz14us/ZtahUwMgW8I4zwhMfEJ8xv6QY3oLDrd7WZREKJCVDCKPPYBh3og+H
3R6RTYyQZAWqGddUYb0cpQYsvSMt/Ebw5KHTJPAA/bKXFYjLu2Y8MO10TGyXZeOn
Er0qIcgAUgHied2gh5oK9oCwnVU7hlGqPa7Ab22sh475GKntUPUyyItlI+pQH/mW
Hc3RsRQSUuK3e4xmEjNhO5eWV5nW6xuNK3O5MtrcZ5WYvjU+LqlwcAiLKeJ6SvXY
TFLcb4ZTi+MiTmXaNcgdEauO87+a/LnDoLaJbZkYiPuB/gaKoWsyUtx73o1sS7j6
`protect END_PROTECTED
