`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gp51m1IEI+Y6Y1/Bp7rhxKwx6YyxAWIYunhMu63Ts1s9IdRbfR5fS4CB//1q0zKn
i/0TEpfgsuKg1VhLTGW//Pa+MhtQwojL2IN417aUFXl9IyrLXZvxq4x1B9YWbG+p
FlY0peFXD3cyvBjC9oOqV9AUfT1xngLGTiP8hf8ssIp4j3ZKJqZMcdOibg3gyhFR
olUxXBprpbM4d+rZ7LOt9ebMpUwN3ZhnEQx2VT9aU1XmLQBs9DPpynlmoNUX7q5/
1+NjB6EwubaCmi1p3guweaXrov0hycnrMkNaw31/xdKRRfFYkGG2QRGWRPXC5Vp5
FTXbWBVIWKIox/Oo0cl3lw==
`protect END_PROTECTED
