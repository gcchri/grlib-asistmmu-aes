`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Df6nFebb4qkBe/FtEh4Cm1aOesg+m85rfB16LR0dqCHg6RAOqdhY/JGH76Ew/2HY
Ypl3yeEf7qaEDlqxmkPjCjLcauOIpSCfn6QH09y/YaI9oLXrnWTYPTfKa/Pfdmeh
OjM7f5wK3YPBKbLyfdLPU0jMIxJH/8LGpDBreY+AyuFW2Oit2j4fR+9BvjW/R2QI
H7U5UHH/ByAthsrbCWiYWwYEcLGci3jaVY+OimY4ZVV5onNvEPr0bUsEg6nhm43Q
+BhLMUrYoMfQL3eEKuqHRenCBk5hPJwxmjqmtHLCQOlGaoIzL/4O2Ae8ZDuLdVA1
7pcoMxq/BL3hdrUADlSLUJ420n75l4BhO6pBH+O2Ml2b+OxEzN4SXJuo78R43HWa
fl55iQJASD+iqOewA1r6kxfLtweUEvC39NUaZPPE5GitoBUxU7A1RGDXZSXoJBxL
L+achihra8nsvFG5RwN7K1eHvWrM4A6Ts2NClBfH0wkCeDrw1t6yd+eEr0bgv3dZ
jjSx/bq0+uxsYkp7WGxP4p0+4arQPntMxY3wNj3DwRgf4/0Yv84IfHB0zzK2nlz1
I6gEEbKYaGt12rOLkx9f7+esqfbgjRW6CtcZsfF0K0DfYvMtjFtqjvltFrE/nefj
+BM3H0YBWUZbKMOXjxe0+2AgdjCK1dMCP12dxcN1uTxNV/qs3xs7Xwo/mOmO+HZB
EMMYjS3yYJJ4bRbTCh2Pr613vFq969c0a5l1RZpG+aVc/Tv0h6OrcbGysZtFvxEG
aDmR/QW59EULyJcV68FVTy+NIHldYRSz2leWVP5VrSo=
`protect END_PROTECTED
