`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+yDRO+jKj3gawkiuwmmilEi7K0kZqCu0a5jgnZeK8eR3rZxtll+cwyXnAJcI2k+S
wT7mtbIk3vvihwWFi0JE55Upoi8VGqofFnWyOqTR7hns8qvbu7DtZm1Q/HiRhqqj
kBBxlsvfdHaBUDGQc0EJ/Fk/HSYmWU1UsuSDsOgZxnpPVSYn76qpTIsW6sR0kbDJ
oYNOA6SZw9X4T5cz4pFSQnQOvcAu4bArOvGWnDac6yCXSStDYQIMiHYH8JpzldV7
Vyl4p1QHwX+LA1Cr3eVGoQXSPvCONzkR4REexml+m1LvYoqoHkchzWW/uW55UZ9R
43v4VI1VxIh1WQ6Lm94ESV7hSwjVLIC2U9CK0fDBGLKIXdlBT4OslQlrEH+cpo7n
hAXoBG9oIzk00i6SOa+RP4m9Z/XKruuOt9EBfQpIsX7HocQ5oU7ZHY4PbmA/Zm+7
WgVRnbhMZCtNt5Ro8BEyvdvFwCz+2Dj47lcuYNmSZaoF3+whOXa990LWA0rdyP9c
Qjpm3hGcp7HLHMHSGAQaCXDcjAcgrG4nW2TSP/fs+eOvI8pHZhYRg4sSNhX2FK8c
jbr3T3t5FJTq4Z/lbTSrbrolEcLlxmXb6NCMnYp+eq4fIOrH0YtI1dod+TcFUHnU
NOLbR/XT+x5IMVfAlUAHitxT87TNtKudI0ocRNS1Zxk7G8Mie5kZ+UOyb4i4dZNW
5L3gaYoGH5UvxJc5zJJ3JVHfNDW4HpxNQpYayC8mFP/VoIOldY6hYNlV+aT/FQwt
EkuoL7YjbupWag6xUGAt7+iVmVwmpI3UCxMJADdSOPPOUJ9JCNsQdrnvjJoFCqq8
35Niup4agw42nHK0dDKzJSYFtewLH7lmw0Ji8iCpi67nS57PEBC1SL+asycTJmZL
y24/ZuMSBLX0CIByomxeKuQZYV6NAYshY7/z99Rpq2q7mJO+v2kpnm4OO9h1QKVf
qS3W4u2G9/z2zUkd4YP6woxq79uT2E4Bp2O7HSdo+2cTXdAXGAE/hbB3dHBn0LS4
ciWoNjbJiFPKg6TS+1COEY+hBTOBQYy2lkYEFZCzjzmNYgV4b3YYEmy7H0FNY/0p
ON+IO66LnxTxjzgssFuwBuC5fhebtGn6MF7fr21bG081OV6JOokrKxmx2nmtYuTK
83XWQc8Aqw4Pp8mtJVd7Kh5wVh0rZh07c1b1yFKebeu2YPDnzPGB7D4a2PMjJ73Y
wenPxhz887sJYkaCZ0OPzd/RYPKaUNkzLjt1vU7u9bTF+7+Qdxito9AmYng8b/kI
48VU6KeoiAmnV2B4YakibgXGGKVOufYFJn6ZHuBX4EmnTHGTIjk1EATSsVR4A/zs
rdE8x3Z2IBxc0X8j6ITrtxymaUIThRvJSPO5m9vpJJClxzNq1Bsk1IKUQ378zoJx
GWaUkDu77TSgdn0H3qR39Br2+qzYucZv7aXcwNrGwFT/oYJdrSJXMy0aVeGN7Sz8
Vi3IVtn/yv4YQhRuWJvYRAqJruYcyveYcec9+Kuch06JfE4LhtwGQO4URURVt+CZ
qu+46fDDRKlHfxJvxe9keIQT7sk1pnP+X9DdXjXWCOs=
`protect END_PROTECTED
