`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4naIjt99ggNMjX4S8IQMCmLw1pY0K714yh2dVZO7qFq55MbV/FE7zrAdRXKbQeQ8
zkO6oTZ9vcfmaF+cEPHMlFZQxeGSa/B1ErjYzQ+JN0fk26k5YfHve2bDVuJv13T6
Ye0xd20n896rg0eFWuA5o37pM4JAR/SSNzZNH5kPIWwKyQu8hX/ztqIX+Dl3Pi5L
1gF94D/e/niH7yBANmKelupctZgrq5MOSCmUyQRwkrMdL1loQPXMTvPJ3vi5jmvJ
gM3piFEWaAkW5G78+7ZlFZxj83TvXaBkNIDkcFTeicp2jZ2T6LKREW1hI2g0Z7Sv
Rdk716lmWnW38ECf5fp9MWu5OU7JD3EsO7TKnX/+NQJ2Oe5e7szuSi9NIPV/2Pwo
va5bPPDjvls40vZzPP0bY+zX9x/zWqtc5fbGWxkiiNiwyG0zQlA/QwTo9zNIqGo1
l14bzjfS7h78PWrHEuJ0i9rGhpizRxW1qblOTTo0KUgRrR2VQ+DYRVSXS04u2WkV
NDA4MlEE55pXZAmLEBoAZw==
`protect END_PROTECTED
