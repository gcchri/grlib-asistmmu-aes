`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3in35bIa9sECButXNvBoDx3TJubUDwWNMRWJZ1ANYkSgiCJKKcStgGVmmR20xay2
Ppr1u6+eK9c6aNKJbxU57WGyxs3l5CPKKr93cguremWR8L5LO1Pf9HNoKHpw/i1B
wuhyc6YqIbUERaL5vfeDdMzaP1xHnAcqkJNYSkzhdHLXphP38ppxg3/jt5h8PrDA
f7lxcLXH4okD3EdACefoLE6jRSBbtZO6vygriC6M7HtWzUVtCA7YE0Dv6eOB/ixF
XiVARR68xhbCcFw58s0stmjVIUEcngnKo+rrl9T+yqMcKFQDve/ai9XjJRC+/KTQ
uEREMkqkNC7VYhtDrMMPhxgisKWgsTPdnomaayg4sLboz0BNX9w7q/XIEX9UFbCP
nSAl+J0mN5+XIfym2eK1Gzp7BG1Q8jniu4YTTZ27u1zFW1CFebAom2hhMJ30MSRa
u8fMHpsvgXZUghm4onmP9xL7SR41cHfaast8Iur4X4GbYqCMNqfkg37zPEBeGn9n
EySK4FZwybrmpOvrnm1qvBa/VH+Q4hTdFb5ni4HFGPMf6ZQIDvS7gYd7+YyVCwD6
54elD9IWzGYQesdqhPaBNoq7a0KvRoIP5855tylFqsHe4wUB+7feEmnVF96mV1h9
MG/O4reQ+0/Aj/qPw+v1crgc1RUwSdqQkFqsbFCFfNb9/eVqIBP4qcRNKLUAANg2
N/iSepWAW1ToMyFGP2wHxw==
`protect END_PROTECTED
