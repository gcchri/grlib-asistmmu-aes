`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xNu50+w/qTTK/Enu0GOOtWSlOfKSJlMb46Z6O/BrvhLphIiRWFL9IO8mpqf4fYwI
IYhlnfBfbqyw94jIdtY7iTAzbTaUYo6nu0B2yL7pfRsyZwu+HPQtuhzixmjehAab
CsDkFUm/DQG9aWj7NvNzlL3xIhzhkEPnRPqTFEyOOKvMoPO+lAKf1AVpUEB4g6Iz
+O8dsV1GcTWSJdIDhF6+IlgUMiNDCm1hrsbra7jWazK39vyooOHmHDuJ8EBOJWTU
MD0SgibZtYpV8zGekInT22hi2GJxngy66QUbeVEBsXGeDTLOtmq+LAwwj472gr3R
qM0m8shJysA06LJLcz6NxbmrFBCovsJUPSM8NSMMGXnP0hLE7V4UwreF5G8MhGWK
9OtKaLd/BHvXy6JTQoX9WS/aR06rnCDo3NnJ5sPjNUvK/2VamyzkYt6p/7hpG98s
EMMaYYc1V/mfzVXWv24aYg9ddHGyd/8v1uwRz3jPQtWS5zam9TNWu1tnb9xHogJN
taJjDSnPIksIZiTYvaGBsck1mbRBMR61H9OSuyrQoKniixggXhauCpgV1kvQPX7J
GcfxdeavkEHGMboyla7jEUjf4v4WcoqQdZtxyRKBG7j8MbIRM8mlz8qbrxu1QdkN
5y48f0E4q0jLwnl3cn4+RaqhVBc4qOZGPyj7bjx0kjglM/YLhvVo++ZLY5LIZxFQ
MXlWO1Vn+5PzLQomDIawtg740WMOLjzWOo7+GWM7DzY=
`protect END_PROTECTED
