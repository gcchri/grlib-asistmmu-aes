`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kORbJrJMYauzPbnwsoDnhtKWkSzk2/K7PS0gzBmWx9Lsk5jIXSrz6sCmIFElik9x
ksY/ztkhnrc+3O/zaAHscWA71JxB9xO+IH/dMLyckRgyTj8gsuYaULjvhbVweXmk
VJeD6Zcbg9GjKQ3R1soVMg+byO93WsiHi5Cb3aCs38m09hQCFyg2dx1w30lOiATU
F0bZaheyZo5BcX0ck21N1BGSToPno3+y/hKsScGiDFCDBaqyoZ/EhpO87N2Jh+jW
5nDiGb6M4W2ttcapxwlcc2qzGGsirQ4li9WITK5ZU2Fwafxh2w5FO2xVYOGIshp/
BN/wqaI5sV2vA96yi83rdg==
`protect END_PROTECTED
