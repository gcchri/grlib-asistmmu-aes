`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uo+SF43Zoc4d5NeWzGgHSz7HWFpkTAkf5x3SfvULoOXEQGW+shyJssRUyopglLZJ
yAqOMzp85AwA3+9yHLZfuzQgtz7p2DheVRdg+E+1aDPscrUK8UyK10/G3QqcUfeK
eDXIG1G3PzrP4ygvAdTLDPF4BPNdFTGdzhRZLGiOYlwpYyk/+xro38LlDI4PSPki
F+9MDO1GX+OGZRDEfibH71TaOyeqS7XkMnLkHGsRXbnlhoxpAaf5D2sefnC3Mmru
A9Cgl1cW6FbfCkzPb/i3fg==
`protect END_PROTECTED
