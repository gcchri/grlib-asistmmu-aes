`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ek7jmICmffKcSFzbGrSmZFXdqXRmkfyx/ZaV1ZUnSHnOkkTpW4/ed44Lo1F1HutF
k9NzfoffAcPmKFcv07E0xol/uQVkxmq0zmk+kTFxEBwiRWX91j0NqlOiQOnnVzZe
cJySHqsW/Z/U7Uo2avV4f9kQ4ZPTuh7M5qpLyTpVeLis3/lOJV0s6oUvDJrkoThs
QQzv+uKr0W5W0I0EC/OZf1LXeg8J3eM8fckrxXeJKNCbIbRUrE9rnkd/MOubLO7V
JdEARBZuQaWMehJ+C8r3AEA35TNvQxrrWrVMiBUC+7Wr/Y/Rocg0WoGOLyrn8P+j
`protect END_PROTECTED
