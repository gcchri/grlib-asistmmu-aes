`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RpqBWCmulTG6LjeHWD+yJRmDbu0SxS8OeJo9TT9cDq1oTMTDI7seszyuXvguRNIG
WY287uPkj9mXt1xOO5XncZzcGNGAUYiY9u1VwL8fma76I9t+4WAtBwg4boM7la//
xvjs6z91zxeu3i8hBhPTlOZfR/tR4J9fO5KKgis7+JP/f9lNmZ+cTbfeWJPNCB5w
9Z7jywZhp2yxo6jza4AYNdfg5vKgSO8YNU204WrQoQKRtnRO+TZaqFgIy+71EA2P
vcxClbKyImC9tbpOdTubVuPX/Ir3U3FnZLCN/8le6517LsZkykNMcVDLAPnHeUiL
RtxKjL0gz7KC++s55ehWv36rfw1pPGAuiPK6qtVqJ/8Tz86mpsdcDoay0OGf72EF
woN9OSCQc9BJm+2haATH2W8rrVnsqiw20GuPLR4wwiVlvnpHMm4o1waUQPWMa4HD
OeppvuynXHNLyaSEjMdawsgzWxwmgLGMefCRzrMTZSw4VqX3d5Cu98rCFTntcy3u
wFEQ2Ym9E+at0/EK1bZdmMNj8hgKYpfIsX/qO82DgFGH3hCddcDTijaJw1Sv7gxN
Ah07UoOym4EN/oVDRbSwDg==
`protect END_PROTECTED
