`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yrCh0IuykVfvmlTqWVzXhxDOzqL1mRK4zXuZFW70iWvdNmB59KRprTBWNup7uHg/
8pZtuIy2g2bA8oAb1JrI9aUg/vgeWfRr9MvrIC4S/eR7B82s35AdezS9Xoy7h1qG
WGz0gDpjoiafYvm3uM4ADv6KLwZJWazzOdD1VrVAChXNNfaUmnZIGv9OOWSYVwD9
T9DNKIuKqFxpQsPU2dcGzXNRPtc1r6UryLJD9+4kb1XrPifZGq+fyE2bd21Fd0pV
lvTDBexFDN3ggDrrOiGc04iB7w0Qf7EMoxhYupEXSlf/XUuFAaj6RyuWQ6wI+Tww
yQ0e9VvZRCmlORGVOPjQHnHx6p2RZYZdCIOj8U9YenYnHFaN9yfBIcVDmC2VpBly
V9q9Eh4jcy2RWH51cgnpyvRUjknpBhfy5smcfQb8jPrPjYd0fmsf8UR2QEuj2AiN
CWCd6PS36tEatQxOU3Ys9f6RkZFaBEFHdBiVOdlUNLv1vrNUjHOLwVnC9laW6XQz
jw53fJxJ9fPL5VVNlPA01xL7Xj2gJcbH1etNMNjkjPgQFUkKwpGjd+FNXuMhoJVZ
Sbu5I0Tl8eZ/yUUSF08Ccy/kvtX2EWsie7l2pvXeKdw=
`protect END_PROTECTED
