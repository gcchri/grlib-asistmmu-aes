`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KzY1uabuz0wl6KvyXuny4jWhesZ3uLCxOF8n2e0WP9F71RfNKYkg9b4W5mJbaUKP
IFF8RrvfVxM2UaN9e8IOF984KO/SFxMmv6MJW4u3NlcHEkKd9jiYbxSRmgbHkjY7
co2RWrkfeJlUlpa1LQi7vHabfhLJrNWZ12IyWycb3kJgw+AAetDZ6ZJmno2v77Ud
XcCeAkAzKBy9XpwTAkzfTA9GXeVjg4d6+bqkPaZdgx9vSFWUWy/sth3HAE5cunh1
lymtaZ5vWLo8eumkqzEi5jhvXa3Le0AKcisTEls7SE/3ofUOnmaEiUvc93dyy07U
QnKM8PggUMtFAxCvixWbM0QIobf6mS6e7Ze6SGIYrbl9i+/VUdrTEF2WRWqjwNJ9
dxW2Hy0Wty+zEgAgv3p2Z5ZTKJkYHu/Mlv+4C5SmlPBugUHK9e4GJlarWqABuWRW
IplfiSItH2EDitu3e92T6n7sv8h5iCHrd+y641/zVDmBjKMd7Kt0r/FcOhUebsja
N3BiY71Eh1qQ3abqXOJb04cZ1F/3bElv4o9PW0f0I9vZf/mBJ3l7aZixAxymr1wk
udxrkJwv3d8OAy9VzP1BOcpkHo/iaWRzXYhAjh+mjOskERd7YqTNbgXlCLQmtJ46
H1n6MiEuxvFjmc8W0wkjbW7l0zj1tiF9rHe3W42ySXkYReYF5QuHfEM7LegVehpc
aeWh4BumNQVVB2RCHVoieX99OskiiO9sSVLj+5nyv6Gw3OwHKlRXSyz2nIfi03Yn
sDvDXhmju0htIpyIoqXehmIffSJ4fZzCGTjfmRtKFgGbu9oyutvZOmko+suFYGq3
zgnZlO91DjHAjniu1NkMoWOqGtUz7l/2RI9IwSoCiGufJVaX1vti9/PqY8CNTH2g
CVkVtdoDRPxrhlnWU7Rb0i3iBCIoJBv50wpPM57C2ceTjhytCLlnq/bCugCgViXe
gKoWb0oNVEeppkB5WIkOxIfkj4VOoiRGdnI6x8nDxUBGvrcHdGSJRO8518TUyWe/
HgU0M5naKIg0CLScaDpiE/jtbpy80/hI9y+60sy+it/+qXSNO2CETSuUc+x/D0sz
0a3eXlirFlsvOfaG3+1vABmiqXHV6g3AZcywVN1GeYrN1BMhmxJiNItvMWg1Mo5L
8HPC2fpspJaEbeP5v5ijBjsWvOKsyZEXCnaBCZpFrpH1+weSjmQ6h6hpKfC1iTYm
Wj3lAhqK/qBW8SvK+aGDsg==
`protect END_PROTECTED
