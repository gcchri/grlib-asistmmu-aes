`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pjy2XddRMWJjSozI0P07+1PWbcGk84v076r+aao/gJ/VAkPzbO8ehSiqNTzMfNBq
Ts6E/+0Qll80X90H1CivL3cxcLp2BeIb324gegpirBPC13YDuPfVq97ncOcILxpQ
brP19DNQKptco/igHA0zPRSUMCW51bDoPZmfiSHmUVQkms59UCSNWTGTzpdcmz5J
uvvxmklvIabWzzkSW+M1JpbGYcMr8jcC1kkAbnX+EPrWUKcnokeLy2dJ83wT86Zt
EGVSDS26bB9zkywCS3CW/Ij23M7pnSYwKrRszmjTMkKACGbywV7u8GU1gc5TbjLR
S8a5fmARfOG7sC3xZ4fbpQ==
`protect END_PROTECTED
