`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MMAREmS2HDYKdeTw/79KBkHtnqWZvp8Madukaj4tAxci+JvEeAklq3yyzdrTQ+6u
WwRY8e4ZVDAXfD7KIcaRuBnlkTPBev8Ea+0Y4sNeuIdZtYtpe9B6nu+JRaglXiqx
PTcaqh7H5wE4SL/43uUhcrkqq0UstiO6uZlIx4Vhc7kReuI2EqF273GqUdJMnLSu
kRMYVMI10AHHQFs6QBu7ftWNwo+KAw2h6U1wnOezny0aBmJ5j7MAqXTVqazMo/pe
fvB/PULCIfA4QCJ9FpgZBicp7pSoLpvETZ7PmRS4x3ZcvYKSA30FnHq4jHnTzy9E
jzuPSdqYR8hp+1hn6xR7mj4K6eUabAXVrjg0OCgtsdP48f52RqFyaD6R7Ddnl2it
uxJGKxD6REFEPjDSZf3MvzWEKNK3qjjxUzXRSQkpiR6VBWclwwTs2GO1+yNbkcMt
m3wECD25Y7S/iBb5jZSQr9+U+oN6C4qke+13GlXKn1JiePAAwpRAes7+02rcqBok
svfPVHvp4INVjnJC3EO8Bu2FY3pKGJEkrsPsNqajDvjWxpjLgY22+jFlgN8Xjiad
kPaKhXj4BZZCAlVHlL8HjrswTVvAgezfUBpHjFf2IcOjlemHSUq5lqVKF5ow7uV1
bJ1ZeX9hRrsa8BjBsdu+Wm+lkrypCbcTxdJwUl3C7zxlQ1sB2hvw9vG2hE1gc+48
8PErVMHN8ireeyG7wM46zivw+NmOJ/VP8WBULx4JT2tmkmalxsprWR7Cjzx6zspd
OolNnpRKdLOuZaDuNC0M3v/g0/6UWFA+238lYQKQ1TGu5JwtYck1e4Mmlrk8l/fF
sM98bcT75MZkUnBQ/T4rBhl8xSwRNiLeJz/5jjav9/GmNPsl3OeInYee5CU5oF3T
9q+VZ4EbbEQFJ27w5lPgMQ/OpJ8vQbxnEmjbtg4KQSLIWbzd1QEvnmCDagyO0D5p
wnv2rVt3chl0mB4NjXud5KlaIxXr8CBLRy049/lPDfbJ/1PRLwsxEf/5o64nzWOD
19sHWAONcrqTLPIzi19MpBdfJBoWWPHyoktRHOMK9DuzhrEvK3Kh3SDdP0V6vzc0
Eu1FerbkHla+69QPFSAR6BCPTKjpZ5vp04RSFzEwM2eQ7Z1Udjwr1FHYAdqR2iPx
MxkYrqlAG3OOMZeC4Zprz4w1xWVtLgaJbQKjUr47YsuCeNpX6FugWHNmatYdBDdg
s1LrWte88V8+B1NUOXFTjIU1+PStpM1iNvHOSlSRmph9FILFyWWzpf/nRbqniNki
YYhP8lLsY0T7TWWA7lph2z8yO/EdHWVeBoAaWSO9sk3DOWpdJU3Whj5upH3T0JJ3
keu1Ng14KCxH+etA5wzvphF5IfBAgyvydhlg62sgwBQIZI0l2Lf3BzkNr5VzEzFM
Npnav3gBZctjHPE12YqaiBVzb/nGYBdypiSSnlcEo/WccEkZ3Uu3lGtQF8A9XtDb
`protect END_PROTECTED
