`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0tcxdpylvTfk+U3/iRDiDXEExXHX4i/Gw+y9gNcyheCszvGfAqHDc9u2n7O4G1uI
3eqQF31bUsKcWVUE0D/eDf7QnOhL9lIDBP3XLFK2Hu5Dn73iFquOI4XHzNa55Nn0
2UH17vq1M2JBw+XF4cNzm7N5/fW207NGBSRxz+6lTGkfnspZf8btt107PX4o1CSN
COrBeSpfYqiKCAnoaNe7VDpyHrBqm23TEhDji6ZV7hSGin1OqssgzklIziFl4DKX
1p+6ZJZd+9/yN3EDb/LKIgDs3z19+BG+PilrXx1VdTJGel7Ld1qTk/rUP9IF8I4p
2mr0QdBNWMSjZzstM5rBLezIt2cNVh2F/lzGatLpreBPuKlCKWi7fWvdQ5Pt9xVj
RzjNEDquou/TDYFtSSi2BMMuETZVNLIdvW/QjebHMhuBKhyQy8UC6kkq+HrmU1Et
OzSMdTbS9BYMFjTQPBvenBhna977neHseRBTumkuF4rAn86v/ch6zYj/KHJ1ItSp
MMupN9fSCHCpEHEf6wTnbQx6ZawvxruLtlL2t0P9QyCuG9Om6o9t62P2c+ycv3Fk
VSCfXpPeIPOAXmMWwUuQmZ9+7zvY10Cf++fS0QZc8/mnIMnYG/ZkUYAQ5iB0rMDr
7rAIjYdfqv1OTmy63KMdTuW1SWYlMc5btam4CaZHh0lTo42OCIRNw57/jSnOSKZW
K3NfDN71TNZWTFUjsa+h/7zDGiD3vDFZCTBiqe2yNmqncOQ3T6rM1YavKvWo9HAT
texwRf5f+ChqrR4pUU6K+yZrfZn6LZUpvyAFQawjr574iCTi56OZFDmHAAHRCNd1
qNkByWeGwG0DhlbHD8HzRpUYlPp3p9Fhxrvg7Ym9YymdGWNvYNF9dnetQ7cGqQsA
SYB7nP9vjvhgpYJYDNOKOzEBb5vGQB2aH5zfecCnaPRhZPAccGDRTMUpHOpY4GLO
fFdt1uo05krDIBjYSVfcVl9bVwufq6yOc4VwBT/7ZIJWZ7v5udoM71swagPSByD0
`protect END_PROTECTED
