`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yvddNuC5tGYX31/JRZB15YBs8cV79i6eK/8ciI8Tv2oIVlLJIglcxPgHlUBhEUhQ
uTSSm1sJT9FMP8pA9WsKSHh3C+dOssoTBR/gJonPLLo+pxszRge5P7e3kRKRxtCC
NxzgfDYKLKf1biZ1CGjcmtqszhJrpfeRt5dNwhe02GXHAgxEQMkK6weOgUB62V6b
KKejRjGUKmS61W2r6+mg9kpqj6rW4fHChFQb6E4tjHWM47sWOvN65/qlqlJWrf1z
EiQOx0gzf6ZNvvwJDH5lNBv0LsYxOJzh9TRZw6Ww+G+oBToCBSawJGDaJrd2f/Ld
yFlSFuH6hFtPnvEeJgcR3j4x0wujDyVlaOnlKVr3VNXJzJp467Bu9oBrCWZwmpc3
6D5S7gD77sKXU4YIvCaNZ0NeDckXNr3JagHy7vFtC46qDlXpemv/Ink5yvyxhiw3
Q76f8lo4lqWUH5k3PTv2MW1vDbIrv2V2gMLPPKW6YgYRQtJJCOpLRl+Ezi8zInCN
M9ln+OJANzxURiqlqlHkGb6r7foTh2hEZxgvt4y9XkM+EJ54WafUodG05yTlRbm1
Q+daj3d7NJ/JKFoaL3D05xd1SDIgE/XwF5jyp7Icec8hCB6CEhbhYV/z7zY1le3r
fe2DM2d+KGLtlED24VyRW3cHLhU1IESddDdE10/agPo/hdWHyupsKGMLiqPuZLpJ
nMru75zg2Nk6UcAuRup4Tgj2znleTjnfUxTKvPNm+34MmiSFxrUJOM+MTKMgN4Ff
nvCC9DQTvia5nWwpc1u/Snjtf5VYY4rGIzZFNlvm5HP1gmZq8ALSl9UewGRuzOmF
V2YTsoqYj3OuAkUb9i6zkX0jVQpQtQu/IO3rVEDQJ+KXNnhBZD1wTHWzjph/Kx/8
oOAUWiFKcW2TA4m5fOqD2I4atvdSg/zu/e5LHDw5je5e/AqWU5jBv6AfuTx1wPK6
j85AX+KKlEmeauy8dlyt8PLGq+Mj78N19jPUbmOdSTdXnB2iooV/b6U4U1cJqwoS
ZKVGdqyPqtBqA92Ih6N++CotiNx9SxsMBcO3ueAQ0ndkJg3V6St4CVyEjjmD5aRw
kc5wVO2TXbFUkm1vp8B5hYLPBe1RBi7mzWDVi/NVAo0Jnrj+/H2a94Ttl2xT/QBb
oA9Sw9qn+jvRIFIU6HY2uccDRZaVSqlroE2sxoJ+8dukDCmLgQ2LXHmD6QQj0HL5
7+tzr+MRFm6fEPCQ1DA/UH4LZkWbxYKRwIILgM4jF4BJhbLPwKUiW0HJ9jDvBXvQ
Seu34WB+crTRPQL3DtmsYwbwIqbZuvpwgEqEAdpujBFQP+xoeaZ46IYNYBCPY4JO
Vcb9Cibq1NWuEGL1GQYLtXMB37J31HXD0+3jWp5X4bjH42iCWro6WMkyGHstcoAv
zgjMjd7HK50JfFwD4BQ4Z1ilMM08UJ/nvSDNS/EZfMsT9u4+aMZBoD5gnrSxxf3C
17Cc4B+rOJWYdv3XRrkfqr2yYkQ0nUlgMN3g48GafNYYnYKAyT/8yvsHnkkMPA3s
L3viL89wmqapHWNev/jhC/f4xoDD9L2gxDhJi7tbXjKwa6YQlo1kEcDPPS2JKuop
VdEEmjg883YGn4l7x6GnvLEpZuZo6YBSVqGwoA7Zg4NczZmzDvcMYueriD0XmvJN
PecfREjgOT9jcvNpdPY4M6AhEhT7dT7uOrVqBbdVkjpLQ71PLXuOGB6+u91AVRjl
BjyqJMrWG8pzbJvo7JI27Br1Q8I/TwJXZiyIKcBxY/855Wyx0rJiTY17no4mH/v/
18hAJdcWzJfqalHTSN9JZM6PPNq5jaiIpqppYCF3IUwTyGEzWlqhzGUDCXG7Xsqt
KMZPuzyG9xI1UtFtAqfRO1SvMRgZpaYckEZyT9TNAsoxDFrLr27oOIYGqpOkg4Sa
gi3PeO/lUMJT51tOyfhkppHViE6WTUAG30SYlxLc+mZprfJ6dzkwNEz93IGfgpnk
o2jX4yGcMNQgSMUzlKp/1b0LkjvOrFUm9aimzKyfpeLlDs0nLpcVJt4tEW6BryjG
PnEPN/6eSQvVBleMeA2aTN9Yt8RnDuM5ElvtgS4WWBpnHfiv20bPSTFlAUJyO27G
91StscpoSazLa+7oNZDjzIBY7upPG1QqhxxwCocfbLc=
`protect END_PROTECTED
