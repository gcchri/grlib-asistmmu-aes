`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HJeRXW9MRXvJx9kKSrR0aniXlf7EqfxwtPPInrK6xJGwejgf3muJdM/zZ0HOwIKH
78qtMoRbHwZLFiM4gJbxCPBiKoVo+NUgdf4IvGe8ks/K/5dcWmP7bV3IDbzY842G
QvH4h07M6rBpVeoRoexkAcSLJTrkQROzWrBd/1WON1rwurpB/RA15SoeFM6nTOkN
vNuSS350xsdppZdm8mHwc+uiOTDJemVdocM/WZrwJoyKmy6W2CK1xUCaWhUNkjai
vlWZ93QuSlfFIybNh1tcdtqsq4fHZ2k4i5S8PRfYWS8tVcUZmhmI9qDMQ889qmhQ
uJ6tcuGjQ5JkDht8wL19OhQ7PLNmbL7OyZjvU/FDs6J8Mps7pnu0XGdz+GYkhG/y
lnql9Xs7/VMGhrEfgzAr9g==
`protect END_PROTECTED
