`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eUBBYN1Fqe7KkPqbVi3Uh4Q8g4n/0KDhN0JEtluAtTYMtWQfIxBwsZ3vSO3A4pXl
mgjIIV1/LLRXDkSjRKuqQxw+tJHYbTboy8vM98eADMBXTagyTrUjwcE9XylCW4ZD
an1QyuvFL8lTFaPODxQWMe+rQYnzcjHapSS/N09VTax+0ZmVj237/f+sBQ7HOqF4
PFWPwN1pV4YxL8IAm4uuQQdWNwqqSvIjDTY9FiKM/X6Mz/8ncLB6IX99bx63aKWC
POmo7foXOwgC1Izdz5DVQfdqw3y+TwZibZrp/BLPo6ehqyJLFLlRx/Tw8cYuwhEJ
+0PxiHaiyNM+8JATpuM9h62IhpNpTh33tU9fF0sd6+bu2xumKwZsXfUpeOYzJ9I8
+bOZuMGtqM7sKuYmSWNySRb03POGMIB1BzULQ8qBGOdoaYpc7WG4K7Kcm2nlon4L
7cwrmhfMWk7gAcxwV19xZHnEyjTvl0qjVp7Lci1u9apxqlvbn7X8Z3BNVS7EPKAt
ZT/vaX7SB00ATGnexSneKSd97nLbrlaL6gy+V00mNy77JpfOo9iJMyXLr7BjdC/9
O85jZbxLb21hvrSay4qlb1g3RzvZhydC3XdcQvzd3Q0=
`protect END_PROTECTED
