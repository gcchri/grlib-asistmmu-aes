`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eR08BKwhxxOt8mJqgARMTCS6k56RXXPXsApgceEagjczQT0L+Cu5GXjLas5AQtwH
SMw40Ccw5ZSWh8lqZD9PL82Mu9zPsJCebiMBmS2Yg6h9/3RO6J0Rtv45+SI78ZJY
l7JZJesxP4TG00/GDmwyhrz+8vjVT+apXt6/0osd1CVx5XXoRUqiekcnAt16FXab
ClB/GVQaTSnXJjcqK3dSciEooB4wRAntc1+tPJBuA87moRhuowdUB4sMI8iiFS3G
2lEfsAB9V/zY40p2xoIUEg==
`protect END_PROTECTED
