`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rK/qQagfUxX8zY38qJjRjsGhEq2c/ReYLfyOkyNCmmOyQItFCWQQjbq6svfrszvE
jX37rNm7tPXQc3rNMtOUUApRJ9D8/RW9LTtvMX8T7Z3BT7nD108xCzJpQ/95SGfE
BXfDyfpFav/ON2jEVhWroL623COh6dtUigAA0VNfzmrJAZ9JP4QjUxpC8wrFyA/C
iELD+/YNUhuX5QOE48dic+VlV2qZPwWOJ1r8sOtabzvkZl1GKbM+PNyeCweIwYJN
Zaetp9Lxc8H8BdoT4VojJ9P2M2YsciZ9r8yBpWpYOQ/L7MvBP9Cf33MoO9eg2AyY
7i3ithhN4pt16VZueTjIhcAw+GprI8LsADDgwAYabkxdq0c43zPXXc+3sE8xSb7l
t0CXueObI+UCexZWYNFAt5cr3L91oI8snahBM7QzsuBB8sVxEJezKSZpWhlphoJl
lBqxGZRfXb/evg0w91eBcXNW9G5UvqbF8C55+Nbp20zxjvz0dnLec7TrwboTtXQ+
6y4+NHsCBSYSCm2RO20CC9btIaLbKuyK2qkDzoJWi3w61j3TWjknS5Pq2eKkSI2p
dmQg0rRk/x6fxrXUKjuKNU/GKuufG17n+iW1uBucnWVtAOlAQMgK2IZMdYneAtom
wYJ8zQN/BE2fGNuKtUiw7iQ1wgxFzBh1c7Pzkgzc12FO/OsTrV/DdAvjj8QDneel
TmaysuZ0BregfkUPvW2O+kSwE6pPF9LDbwLz4B6age06SN8hxrRmZvzeIgybDFiC
liKE9b9qS6oYteMOWKYOn26HsoQm8KN4P+dS3YMVOs4nvK/LkFbSQk8hYH5Y5afc
H5+ELaSX0ys0UvnqcETxxX1uU70Khq2wCdpeQK5Eqt9WDsxlr3qys9ry7PqCBdq8
sNf6cJNN5gRdFuqG6pIDYebinTc1J7HFnshqnPo1+XlnUXIi4EPn2x9yq10kurIC
+4VtrQJvrFVaPdm/+7WRHNQEJ9UdRULn+l767bVasajFbt+uwkGvk9Rd5LJP2yT9
cOh6Ggu1ThvjH/IX0B0TptSdxjbz0eJvQQ1i/k3v94HxfnWJNlgRU6GE6sJugkbL
GEIRs/c4XVUPiq8W71qMVQZTIaUxjekfLucoin+39NhthISIfkgtRP56Xeu7Zfqk
PVzXQwp6fbjVrhRV6FLT5NgfGZtAd56ZHUYRYo9kEuXeI1fJy3kJHDe/0DQOrnSY
8yAbTx5q+6pl4vZyKAfMGSm0GPu0noBpBzFckOWuF1i5gjErZOyQLiRduG62LPtV
iKbGi+QX/FXix7g2H4RHJAEYwhgLdzNq+jX9V3SyjBAooTF2woCozTeP5YavdVHE
5ZUGWh+HBJRe0JQNLXlKXjMNVF6343O14X4ARoJ+REgAc+jLlOGY6uZ/wArLwl44
WJ6nH4oPpfLMsStHy3MANtXOpjO2or1nEU/1dFR1IN0ZUyIdbNSIlf/3NSNY573X
wLk03tS90s6VjDC1YzdytMqwvH0OLES2Ytq293VrYHggwd3wiAHoIAYAxZVsBcOs
n7MfWbaFqt6lLKyWW/m2opLDhonxV2MakvU0mXKu6OZmzsqoI40G8CfU63xVigX+
FjWrA45KeYI4V2Nc2BvFkO+DPKES2lz3PSeHhvnrgdHq3s2y9ddeG8iIEcE0tx7u
hQHI75D9RAQ0asFZCt3kKasRf+4VH2ScQKW7TvV3+kR94WyLASvN8w9Gh13Tbh9n
i+HbrOGBoGjZ/KZ/ECXxX1ChlwN+tDG0GOUjEvcigfwpgrCg2TP9bWQM670PXwrI
xRH5xGNUgVouf8bw5JVyGlMmzlaE8th0jHs+wPfLWIgRwYdyAEQjnXat6hB8Z5Ov
GPS1W+SEtxTTEQa6+IRBYGrbuig/ZzC8DO1c6VW+0J/fLbzcc6BcKTmxANfySafi
5UAsfzD1ZXqPkbGKdqg7fEo/llBC0gCN3fwNOVHl3H6k17DOcEHwdf4z+yclmLw1
b/H6k+4SZ23bkwQkoBEkzugjmzusaDSSo+4ESlk7rSQYdziUnY7TNtN+gSJmyZrG
DO93odMrzZU/SoAJ6xh1gln3Mnia3eBIqgH82oWN8K8i/oiR/t0z26EbelXGB1Fv
weMghZXIbcxfZcc1nAPpGEXaE2XATmifoJQQIzGznLG3HYo9liK5FBZfAB+5XBoz
GcPFlQuhEPQoIfJYPPdCn3VphumYTdQ2SWzmHA0e/uBTwN4Q2RspKTPbqlLmMlGI
rShXdw4bfdTxcPLi2JWCKhC4x+8CdcjHq7/btwXykBsaDYGOBrOFZGF8gD/MuiFY
w8urLH7diMOykGASFrE+jeP0GdRCcKhTzH8tWni97gcUTOJFDrU3AjhYmeXZWDxS
vIVSkrOXoS2mOs/2I1vmY7UBaZw+Q7u6SS+rqsKyACYCrt1kKGjDUyQj6/9N5Vrs
6lVxAgFLHUjfTF84xYZosR+HAdD9UPasK0qE4refDtLW9J8yMtKnW5YTC/KCBaOU
D1Ng4bninI6C5GCGtdsw7BxKYNnuYAEVSzGF9DkAyANA5g47HK5KB9qcib6lRaLB
y4nnwcQl9rxXp0dsKOU0mDTYcpRdorOmII0xHSQ/yIauWlE4wQ4kddLxWTyFwCdB
Vtl3+pgNuWK33E6/PmRYh5AYHW4aK9b25pYs04IA5Kp7+ChOZyGI/xQbVo2ufvTv
EfkQI5p3+FdZIwUNUiUtD9bOKGck8EhXnlzSxy6BWMHf2r8pla5awm5vXI9sm/DZ
vGI7qAoMPUBiNyTYqjpS29/jRmptmYq81kJPX3ie3Vk8l6sP0qgzPKaDRcfdDAfn
2hNNpQdwm9q1WkP3aVqE1N9far9dMD8Ve7AHfmEAFyGA7EXzBzkTISpq/dlYiboA
7vNhs92sw6sniWrT3cKbWlMPrLyOSvXH5CpuCz9AhTtA30IIoHj37AmVrt/bxVLz
ISPoYR/3N05xa5WaRnGND+g/ll97646wqCXWt59rVtBHHupKPZnhzvXdoWbBZcWl
IzeQqhT2bBe5L+lnZlwmauw+2PZHEaelRH6n0DCqQi2xIrT6q+UaizRF2ugs34iS
bXV/I3Km/ZyZ6HjDD2E6pXXATqCSut5Uwc5x1oWwiVy1w64hDwEQFrFBCOACeCka
QwDfpHE7eYMkAqD6zVKGGHXdmjcoLEj6TaSqf/spk2Ud9bulr75S9qCdH/C0A7J8
c4NyckloVe6SVAuhCp/wm6Ad8DlU+BdHvWVacmLK2UZe/T4wqmSmjfgWlLePdFL0
5KhgohNFoJaH2ViEho+HOPQ4XP+TTxk29DOxIXR/NIIMCOsNU7j4CqJ4kmtZMM7j
gw9n4pnl7ddBl1mBowaDe0Uq87VE++IRL2xrIhnWMgbKWpK/Z80zHr+LYUTEYGjT
zb9UQ4mQDvKWdENemBJJRlSyhtvQXgYDHoWangyr2T483KY+XMVquk3IhfrGFjs6
dFhoM07aIuR8sKg0P5ZGAr6UVHrOtMFRWFQlm05dvikc/6VyyQk2YkKoDlJfBigv
vjsqfMxIiJCH2P8hI7bxAMPptlf0+Hhytabu7Z2/6sI+bV54f4WtK0mdRQfD1kWI
s9eaQzDVaMGE85iQgO/CRq6WoTvNdUpT3DX/2YERKVamdNNZwHLdeBn8EKgxdFAr
yMC07vgcG8L7ZfqfQwvCJhZb7NopSyrQpUMOs0z18dMHMLgJthHMa0zBRhJ35BmN
FiriDQOQ7RQLlJH6V4Pa2gAZtdfjWu89o98SihBLuMmamb4HX+FtVCq7aWcR3vIX
JBbFklGNPSWb0d9Ta8i73Q==
`protect END_PROTECTED
