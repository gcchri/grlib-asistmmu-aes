`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZrmN66an7aO9KgB5ipjH66AHB1Ya+sS9i2m4LSBviQJlOgtpWHXx8riA7CH81YmJ
odQWTtEFgVroLKrjON3Z2duXWWyEuhZbOt33jjQyu8dXK3nCtQ8ZyNnCd614wELy
2E2DBznW2/Fpul5lxJ5w1G5t8/mk0mrrBq5ow4FH13qt5MVgvwG+zw18XDxHItTP
kflomCjz6NDVVR9E79Ju9R3MgytjO/5WxPA7B4cwE1DtRI0cD0gkmg++HHnHBIOw
QtD1tTkuFDbNuCaG2ph3XSIS3SYQY6xW8bspRl2lnXrQhbiC4nlUbLeLlr11qf+5
2iggQ918kY8BM2EcUa1nPqbJ2nQM886EWQeb+p+fFya1PSm1kNcIU+hkiTShKpPB
Gq3Iq0+btxIPOpl1tym0XsIIcNOVma2yqC/SHeWxYEM=
`protect END_PROTECTED
