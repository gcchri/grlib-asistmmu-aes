`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G+hgU80s3LeVDyANSiBdZrVSn50JiCW/cRj6xsk4w7Ia1djOMLZZSrowcH5FdLnp
2VinhoUqAncT+9FirdMDk24H3a9V7U3uOAPisvIfie4+36F8rWPA7HhAP8QFLJSp
K4HFAHk1tu71cKFk0OOK+O/rHGsVA++fE29bhroPrHFtyKigdDZgWbWTltjb01b3
eZ1g3x82o3kIo7jZPjPYgiBfs8z/Mj8nB2x9hXSSYIOGDcpzfQjDS2ir4Lof7U5L
JP3uCqUt/4TG6uSl8igB7FAOCZu8K/W/E5PWu39+vTAIh0guISZMSWZnEDILapMk
pObY2rlKZa+29i5gmeIF2g==
`protect END_PROTECTED
