`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W/xIAIHc3UdYOH7jPYZF/cI4GzhD6TVWIV8AKTkUSU/FmpDGT3xWB940ACa5hEb7
K49iP+WtIUXnPf/KCliRil7YGSfYa7WiulFsS78YfSqWWc+fOYJvb+ynt0PkK4hk
f5mnR+do5tB3Kc8u8MTv/bu9LxKxho4jTfJi61Jdn6aDdd47e3aJyzbmvQ5Zhh5q
k7niNCs3RG0XwXOdIaQUtWnjJzOvlXxBGPGTn9nGNCUBq2aZsKWefJ03ymmKGzFo
6DTQxuk8NpUuXqKP2j42QDWq3YrHblFuxdLenCDLh54xJl8FhyxYnDji9CzqQkSh
0R9WfrjvQGMB0YycJIXFuUh1Fgt2LfCdE/k525JoT4IHqD6NOf9JFR+uj4LuHtwW
aKjwCzC/vUtsreyGaeOOAoojGBDRqgf7y2uMjIQiiP36f8b3PihzmavcZ7hay4li
EhH78m1t4KlKNS8UY36+JQ==
`protect END_PROTECTED
