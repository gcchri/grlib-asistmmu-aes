`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iMgMa/fWpDYs6YQ1fmnQneGCglBYSHhgDcqvRfOl0zZ2V/Hoza6jgLXwuzBg+QkL
kYETVezmVvgFRN/W32xhvj2jN/TeyAuDjuWg0OWYkbMVI5DCGLJth+ogu2aGVV9Z
NSlQHEysb0fx6LkEChzxC94uO2hRXUBAhdSV+Kh8wPRR/crc8SehCYFq+Xqz1+nX
bbUPET4XAGiY3XzxRR3Hneo23UNVcItEuRNfc6Cj9NGsvmZ0VM6z7m7KB543xEev
NGpvpmcFRkRNaMYbLx/LbgHLtXDUuqEeOVLth8NMybOuDAUMOyogK3XOy15Gsc0N
Y8WK01GtRGkB9sIbAGCADooRfGAjBIp32h8M+p6wzi8nkc7Vz7MCdPgz4xcNiDZE
VzXjjlRAeK5thGQ4MLF0bnHUOxp/T+7PnZdmfaoYqReBzHlPpP+lsuGVc0hsN6V6
WPcHgsqwJCkrhrg3mtu0+d0ow9+1m4jbeeTq78ge80tsnMoJ4mgK2hEumq8SYOvk
+4UsZeBnsWNq6cp0zWT/ZwEIdcVKCoetJnxqV9wbSLJdeSfWfQaNUr7DaqzZahVX
QWDDHKTMnXwtE77sJHGcG/i7fZ+pfH1mixCm+YlMP+SJFadE2Cl9yp+ps5T4fGkF
Qow3gWYJ2y5yKToRINN8dA2ZFS38lFwV9qo+oAgMEqJ32g1zJKzmatoCGtzeSCiK
t9Fekvvbmtdr53YYvHZoEU1hXul/uY58ZZShFcff2qcoVNo3fI/gwUGzNfh5F+Sj
QhU7uak2uAhy/eehoDn6AkMxC8vKsgInlJfsxGhdeHIGdn45qiwAR002G8zGx+0k
DOuvVBVo+8mcSfikI7dz5V1NWYgmerWlMf3kUf/7MAo=
`protect END_PROTECTED
