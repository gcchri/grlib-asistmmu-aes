`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ZIE0dHP+gD0e2C26r/9QBlWSM8jhv5zGJykLTpPaiZfXnXoCU8j8rLdeRlE7pUL
R5p9J/V3uahDeD39jB3qv7PL3u4Dy1UDHoOrONOFbH36QMqzKXDlVQy/LSvo4zxg
8t9FWck9IndeDptGfGuyuvH0d4n0oTTgPQkjYcR0TytW3/qo/3wFjr2io5VjNi1S
eMJ+uyn+2hgKSr1oUI3tSxVfxCe3QDiq/FK3PLVsqJgFu+Xd4xgy6ghUSUCcbeUK
mG63tWdTaoL87Jioy72OqqcB2oCi1Ltbletbj3whTKL6OTFuudyxQjoFZr3eXYYP
`protect END_PROTECTED
