`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9cUidd6sNgD57Rq+nxpI8Ossx07lggPbRwE7lC5U0Feo9ubwyiI5+JhAQrITkzEj
d3cnskj8Txpn6SdR3I5Pgs29VoqhfrGqy7gs6eBGXqiRI3F+oXGOQ48qq9cLeq4u
SeGczpKm6Divk6wAwb08QqbRTQK2x55pwA4VmgOOS/UoxPfNW3EKL1hp/x6Rq7Nk
vezyQRF4Vnd9bU0EWqwZJvWpjJTrDeBFQc3IQl0Oww8d+UdlWNxjnOBU7R+S0CbJ
/Y3mL3ELbtKxfleRq+8EK6t7QtxyWK95/KAxubusIuS8c0jIiCKa/YE3z3pLr71o
65xUl2EHS327iMvHz6M5FNk4rqgbFgbzXfmaB7JojbekPowflKxQTPngZPq5Tl+R
z4IMH+/h3iNyGMMv73j1P95eyIxvCyC5tSgZ3/eVRzjcpGflDCurlZmFiVOQX3k3
BYAwS9QDmTD995nV+r1bthYRLC01IRNuio5D4Ph0aOSmwFO/6ATg14IIPut9tW9A
U6iQDdx6XeaTkVTYVyTGbnAaLFP9Va6mKLxAaUCBb/IXU50JVUEDKud2ZWQH+ls1
vBH7wKziYyyqptSr7+1wo8nrt/B2A/9gWWwvKYBazLMd0vtnfauwLFgJuJc605B8
ruLhXfV+YMdO5GAYjs76tUmYXNWlMP4q1iErKxtEAAL40aYWjVtrKclQawVBKh0C
ZBHkACagLhwnPj58TyJu1Q==
`protect END_PROTECTED
