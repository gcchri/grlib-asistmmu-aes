`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iw6gJM156nwxINkJOMFWl0i2gYRscPCXGveuB6v9iYvDqNPzi0rn6o83wKTtnx15
oCmQbqJpSqrpMWM7rd8hUtHRZxw6iHjkMrdfVaoHrM8VInsD0G3bRGIddiSvdwpR
/0MFFiCED+o58O10gc8jai86DYuvsBc3kSeBRveOQc5muUJElvDLaSV7+FBvh/lW
tG5tUgEtr93wAKowrryjJAgbQuI5EJ26yeAD6XNnnQ13WgZvJ/JTFc4Kxko1dmAR
bCw2njt+NknNA9H8TVpAoMow47y/QSnJ6BY23BXh9QlGknasLNAqs7rDh/iIHMAv
H+DlMkrbdEIr2GumzecLIPUe2ZxDspqzfgNzwnXwWmHQ4Q7aGsjwj0p+hMcbETRU
GIsSGUYTkLe1MAAfIbDC3hYlSfGOoF2B0TR6fH1gziNR29cZl7C1hovco1W3OmD7
ZK6N13T0rpfTuRc1miWGBkX1l9wRevCgAxV1ntQRbi6gTiEi07EQ4oB5dy8aLjfl
kXncv5ug/3TVwJ5Nv10aKMpI4dzjNcR+0Z5p8rXiYpdGZWhTHE+C1MKHnSmAnEAZ
2i8lbeeW4kZtC5Rc0xy9JTaU9dPTxlGl6ZPvxmcCT8l4EhjLUYs/VlG3lKkaKLSE
LCJGPD1vJG7JRvHMoHjcjhjMjx95x5NLJm/w+4TgpA81aimKyvzgTo+zcEpU1EaT
VAIGGcGynIV/FRXSnAim+1RBlO5CMxLzF+5YasPuxjounkR4Jq19j8bDUVG2McpD
Y+3SpE4Dsbg+zf4tOKosU7Kipfy1XwWuxmOzAPlUBbYdngFyLAkG4jLsTwBrabR/
du3WS5KIEa8rb8KKLMZF3TtJ9CV4/pmrcDCqfqXsQYxq5QlayTi4jL3wjBAYaiJW
tIeNkK501QXkAZ87ff2s/e3KufvmRPq41hPgGBtMbFqk00+GEUdO6P7o7eSsQhqE
UkRyTj6+pOA+mUIjPe6Dte8knOzqCpAzqW3r27ldkbgYPIg5uHs+KRyentfRJdhR
lvM3ZCo+kQOy/2Z1UYR7Pn5KJsMYSaW/jDNlSX4yJM8=
`protect END_PROTECTED
