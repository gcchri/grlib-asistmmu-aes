`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lFj1GxBch0Z1qtGO/Bf1QwS1HgPRHR5dM9EVI8F1zKDlDyyJVcETx6LzSGZIWMdX
bzBrTsOcloDkcyCr2bepIJ9jK8S12d/tlAxcIEYQz+eucd/vv6VWmTJfwyibMMF0
2+12AwHpA4Zkr3ksSjB5AbB6oTtIx+xIg1RKEInOz2eYxQt+3vwGd/7CzoIKrk/e
Qh5ltwMfQz66Tb9BQNqoft9BUsyjpjMEtto2tFWidAmkyqwLqpXNNVxzLVNEKEyI
1kiYW3nPxWSbIPblH+SpzBhvzZtiaMUxH8vDF6+daKkDn4Q8tUwi8wYHI/7Qd9s/
nGDKCsqcLU50bkQE5GM+BH3nZhNUcNnMMIIbF53KLv92klMEpQnzzcVS6kzGrRMc
osZgJ6YnWCXHgoGYgBHXqg==
`protect END_PROTECTED
