`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ROZfXo0XTdFqIKMxopKV+gtud5Sew9hEXkDEnWspIWrfuFZXzuZ62Vphvn/EpUZT
cKYg/PHanM34e+5plLtQ65+hVX5MKwIO6iiYnEKWF4VhMXMRMr2yaastrHPCWVrM
wz4TI5OUlZMW0Y1aRPTYQt33I3OtHpwXAsPTIqqVMp4yWkacV5/e4tlSoUYaPdYY
bWBJY0PP0NsYcr1/Jtf2MQf3oWj/nnCbNZndj2DCvx8h4bYtvQSD9l0qgwSC7Nju
a3UH7HHaPyiVDCcldFIDYVVrJSIQ9o5VKW8yaPRzpGj/p3+PuB4Jg/6AAzpLSKYj
0cIrkljTzBJRkL2HOs887xoh0sjeAfE3vSe18hG/HqzGmTfkHremo4IwslMUralv
G/qCynsBrbCm6WnXdU1xrLsq91D/w+HfJcgGWD/jwZHtgNOd75kRnTwX8O3cIcUy
IfA0AAG+ZWMfkSmb4bYfKG0MVVTRLShD2hT2b89PGGd0GAaC35sVqC+3W+j6F6Rm
Eauo2FKqy5yy1h3ODsjovqyuL0yTDXBhUeDM8tU/ABmIQy+T8HqSnFZOxXC8Cetb
yT9XcjW6/Ca+Uoz+ZEblvcKExj+OurPJVs2mJXybl6Y=
`protect END_PROTECTED
