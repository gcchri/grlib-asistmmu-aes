`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b1AB4WcNoDSMaaTGaiCgl9rEhNWneaV+sM9+bUMD1+I+9EBfpZOfA0noMNgYvCNB
oZBmtFRNs9/EFr1/wqOVcOkBkntf8H9BqOOpBTYoQYQhmQGn4V+KBah94XdCuK5g
IsfZOEMqRTG4bJkK1gyWz6vBK0C0T72Nn+annhYwP37d5XW4WK9leO+kjZ5tORxZ
88P2HzCTNLKEi1hzK+1I3xDiG8nD0KFcPdwgLl8kbpNJjCWmV5kXUZflWnWHbIa9
oxQ6of3jceUrWOL+ZXaKG+OTIRpGAQ6Ukx4D507nh9Wc5l/7IDDZ1EjyCB+GICiF
LjIp7np5APq9nofpVY5ykW7OYGM0q/4d7XB8xOz2R1nhdDqfn1mreg6mrjhGOnF7
OaVaPdrdN63wBp9x2sU6iMlTdAJUQP/v91frnlppyl1akwMg8kBrJwvD8FfoNByG
UyMA77/pUiGNeu6IQjgorc7i2UEo7RXeO3D1UbaDpMLZwm5XGwIz/vHK3ei1yeSj
RZZ2DwCGIE+mdb7oj9ijzTPDjdR7V2YvamRRfevvxM8rMe/lGUWEmp10F0J6+0dc
QmzuvTT+rWrX4vCOpQrUlWrva3hxfYNuA3Ea4z/7a/c/IRUYmUZuzsE+39bKbe+7
Wt2cnEzg4PmDboxnp9+uWQEa+OhDHtYEFSbx5lDugVPERffw8fCv3BbTfLnTTlAg
CmW7PTOemJHcpgYse9x+Z8Y/WIJspGKoK6u86I1hqcRjRSw23k7gueoT7SlqLdjm
jpw9iGFlmssjcNqBlIh5TGhdkcaO/uVfA42kCT5+R2QzSGRbD9vJztbCD1fQrkWd
gvMWaCW8NhPZzdwfekVBPzAVt+XmKQIE/0Vtd44zJdcAWALbtJFBIw62+HJr61Gj
ZEdGcP4H5Mk2M8BRAfMaejpk7cBoa1JxoNC0kSqkqbFHg/91LjpQCgghadQeSws9
`protect END_PROTECTED
