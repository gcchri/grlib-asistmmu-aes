`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZARq9kZ9wTnJa4X+3YYEGH7vgCXr1dGZMDuAlyLfiOWlL9Gg9/S+osSg4dEroNjp
2/aWMPlwzBkFgXqESoXsdp+S5eirlnvx23TpwjhpH4eazh3XyvO4bI9kLTvO+CH+
CPIyO0Rbm1E0wfBS5ddOlXjKcroADvhOF69xSkbvoouvX56SxYO55exTNlLVt3wB
1zZb88s7HwZloG9TliNi3zS6r20eaTi5WjYO+kvX4VzlgGpxCCFZagGcGHoSWgm1
vr0DoSQqTQAEy64h2ow4zBc1w8w5kWYvtiw6VL/Jq3vpKTYyw+QbFyy3Kww4qR61
a3i1DYo0Zp2MKWQAgASsRIF9RdebQyJIjL2curE7rOaLtj5URGGkH+VZ7XQQw+0i
yW80LmIH+j3aCi6BMZ4zyQ==
`protect END_PROTECTED
