`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AlU7+B60ASmP3F+4h2lJEARovp4xgJTxuCL+3BMUSoeUfbZjxFuG294EfWithYzc
mYWmmW6xdriMNhnWlXkhUtGIvXHM3MBauKr18BN2Ayag84u2LZ952s4Ua1JuonLx
a92VlCWzfaAx9TgaBRYt4WRgqzcPt7EBRmB9yDzM75v4FdR0iQVFGv6a4EcpuYZm
R1bLKVcA0F7cXtz7OFaWiBffrbufqFd/WUOhk3A4UFF+wv7l4cgL7jx9EEVhPio6
Dto7ejqcKhMfNCi2GEPo3V40soBXkKd9cf1GybrAR/usQ+LyM9xwmUjNg+p478DK
oDG5Xkl0uQLE0CKlCtWWJJxrrxPWp+wkqhzai3wkRmG7FBLQqtp0xis7ED9cySIQ
ffh9XBWa8lahIeFAKrRJSFOKFCIX+rJTALEMheiYDosF38HC5hSxNNaXRgE6MhJX
UFAAnbihGg2j9ZjHu59pugk1tjXLSWnim1D4nuXdsi8ru3ALsTf9mvQJ4qWFay9H
ckbBJAXPdwsbbqGeFAEibT9azHZa/kHyNd9TYIfjBD8U/tAtHGaLm47givnrqFbb
`protect END_PROTECTED
