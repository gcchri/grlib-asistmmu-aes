`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CytVcQdQBQNlSkXv71QN2sLlO5+ROztjXOOJmpxiN9zHSkKGRglkaqUE0qSef8X1
73nz3StrUfC/9Yo27BjT+RXM5SUu4tS8N0zZMhPnquKyRbT/ntP5wrxvpRPhS5HR
si16LHQUm2EaLGEsPv7pcf+Z5d96R5fFGuePmywOp0/B+W1UrujQePAByXYxdMF5
t6Nv9N8shXOoofYxRIG2GBCtaaz14HyD3rS0nw87dc1WB0zhi51TiqkJbx/vJMsv
HC2W4BLuRjAT+zpw4RSunopLNpORXmBwRgUSOHUIjzxxvulV2+zKypiQWSb5KpwX
deSxTN3wJfJL4wHPlNq+2uuVCRrM2uCFDf7AkSJaBrCtbjDuQ4kLgXgZxKnPF8Da
2GTBVqgQWE3bwNb661SJsrR6Uo/StGm/evI/K34eHxuK2bg/HDN9u5/YCh0Qveeu
kbgjh1l27W1henJzny2qz5yV8tRWxOKCEALhQ9VmfN7ZTqav8/HKIdPozIEwuPtx
Cpj6ZHk7kFNvcDIrp4UWnA1c4toOPIUu325SxXb46IVktYp59HukTAoO9aX+c9+6
b9prxTths04UNFwp3fIZ+E3rInrPrn5VCQtA7T0pnptToTHEkdxWzAyzVQsiMd3r
fS/OrWGhudco8hAEcQ3oZNk0M1N77KuF8T0CPliSV/9MU6uLqQk/qDmGYeCORPXk
6ki48E49rO+cwpmiR4h8+gjBTCOjI2dkDUoMvshhzxM=
`protect END_PROTECTED
