`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jz13gyxVYhCDviN0gO3BqyTRPRKevKkpuumL15qfcGkAlCQOhZzEMTOZE2MP7Gqx
E7bivmItPDwToAyc0qHZnbD/8fzvPld6AfwZ/2iClLfACsbp0MG89fq1J1rMOC79
vYygE7/h8iiyoSEUpR2LWbcqVht12F6woOOE9CS/Bazvnc7KTgaJ845nHtZhRBjK
6P2NqMLiJ4ATX4mfl18dDiPu9txUX4qm8emTTCQHeBiGYq33mBQ2nHk6KkohxAg3
m9i6qp/JGqM8+RpB1uTASUh43jR535pzLI6afvdfXh487TYxBIJfIoVewWxVVIad
OcU6DfxekQinAFAD8V1aerB5ultW/7wkApBQ8tis9gH7nBfZEVsXgYS5q45wtqJP
Ync0l7to2j/G9ZEuNyZBsisroPtPLhFJ3BgkxYchnYUxsUGo1/H2dpWJ/7iu6GeA
nO0TNIXRB3FcUVFTRnqx1lww4igxQSuZ0kpEVq3zNT44F65KPCJQmZVCm4UQ89SF
PY5egvv/jtct/YGAucMlQ+uHjhYGy5OMT0rcyQLob9/MRYer12vVWzb9WNPzy1KV
7lBKQpiYl6HLzEPFdes9wRaOX0703f8q62mveEsnlWk=
`protect END_PROTECTED
