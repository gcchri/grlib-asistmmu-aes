`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1R3ZDnnuffISGBmtPDH/B3EwFBDeM1E/bslryFCYGmFgU/hcL7cXON0Uwd4z9zg1
qv9xHv0zOiCCbqpsl6Jvbj6OFqKvbEoHegttkl2UU54PIAqifWJksy5GDuC3ZgkT
K4SEcoRC6zGXpQjrPR151Ry1AHHBpggqtnd9livtQOLXjQXplOuOv5CnphvPn+YK
V+MBTzp59l102xvb/qCfX7jBy2JjV7so6w9V688rTgKXMimW8bEOkKSRSY5aGtTg
bpUsP9vif/5cV9ReW2x3uh+fbeDh9RGVvqOTyZdjoZdra/vNB5tM9Uv+rcJt/iXb
ngBkVtbj+ogYGCfAqjW4vBGOPoERWG0NdI7xw2w0Ef3OflZJzzrgfGl0h2T929mO
/2CJ0pbZgH8erjYYF+74TP18LBOk7tO2y+HXG3HoGqe4NuOsj50RY+TrF/M0RWIS
MdxGS4t/f51iVV1vWE5dmZ5xfstPRrEhmfIT2Xga5/mxgyIMfNYPEL8kmEtVBmqs
OzcBEsESuAaPfcg+Vxp5KbBNyRpEfaqG86tPweDOvhHSu6CR889LU4GkhrG4YaSQ
cjP1rbrOm7FXapLXzxfuVtsNQUy3n0dpBf4w+e/TGqcN7uUaiIPTbYWtiSG+FLbV
VfPVnm4v9Ho9OFvSKap38a7DSlrb2DwetSGKIwVZ2sj4ARHaAPARuwue9sj6DxYs
HfpM8GT/sh2JGnI9FU1CA4kEDvHDye3eQtPAjuzjCS1GYs3O240hVCQ+Yl8twbrZ
oXUQ24iMh/rAL5nUSH1QJ/KM65ZRzKmyywcFvJev5ajgehMjYYUOedxWJj26lxk0
pM+ZECvFYuF1uIMMi1V/wH9pNEK4R7WY8mFkfJUIypv8CpAgmYdYWFGV382aCtAg
2y2LjiddORLibWo6KayvQieMFvT4txJJWtst8+lRtqe4aLysvnLrIvGPQfQJ5oAy
IeDc58IbgDs4cRXuKvc63mQ1JrJCWeN+02AALk2P+/hjIIhSYEsniZCfdmG94ZqF
Z2Ll3yP3TrsLv3hQZ6N8mjA4bMi5vhC16H0BGEEX8vFR2ZPV6onYqvvG3rw+9rvG
l0lE63ID1kQS8LZxcHw9+dzdoXsiswqfAztEPC4hnbQqllwFUsEXw9wxOhs7Ah8F
cWVj8YKMxUsy4ccyrMI8TQOTmrmUagY3vZoWGoeXy2H0dX8DqCSjHVvF6Mmy6JgJ
3ZwlCNTv2C3lUaDiduuvhTDbhVKWl617YTiRHp9jZUzKpIDRCMlcfOYKBZkHDDjv
MMKVXAvBM3VsAkpIfkNxJ9rCWgop066JaNcHHZWDOj9cwK7SZe45Exh4Ja0vZQOf
n7lUCs3yYKDM+1KyZp5t9gdIEfvFuJVs7z2Ey+EC17tB9SJ7GHNjcI8yrn4nSjca
iLcdkpp8/CepWQGMnkBiLaiRYVJGJWjugUMUrDR9s3wESvEPoeRsi7SuyNhgJJHD
0dv7s8yHxGJ92hSp+MiiXbcUgsjaJFQ1uWma0/JT0EMnTBDjYWShlU0bEOs3fQqK
mZWrYPiyxCzgRJn1/28atGxg+QBEAIpvicOK0zW9aebbem2ZzBFHgH1hfJyZlWWq
LwpqZLz8KcRahJhSRj8fUR/FgimMDOtJy16vRFHE3G/LJPFqiWkoaHTJ3DwHvOY0
nlppL6Rbq0OEgbiis/Q51fpAQJsdTKbFEXv1D3MMPYqZEHOuOYewwZcvkcLSxljI
oFLmAC+x0XS2/qN0Y5MX+VF+yrNdEHLOZsfAYQ7uhT+TndfxBJ0dHR1wgecyXMjV
yYx3nqucc3iQpm70XYTz6yLYIv4uZSI4rhV/RQwgILISKChDLkvy0FwsvEfLci1y
kz7/Ad5IGdJBh+sLdHZ42+5jYvMM6Q8IGVRhY8LSSK9Gc46vejsSV1S8K4L7EPnx
nLJH5C0LvRSpvCjLUzgjtrcE2SOGdk23lt+tE92HOenAMnspeaCrfjDetmm7wr15
Hs3c1RixLFgXamcB5RKlKiXAoD5RguWNS/Qu31RwbJI45oPVCRqiBUGcvpzBapeB
ZrSQla/q09PAQapII5+Y5SPEYo/0lQh15tWyR1YRow3ahk+nP20Ru6+gIzhH5MRM
oAkWHumC09BmmpHQRRs6Fsg1LvrE5H+DDXfmaaVbbNJiNOyU63hIEASLO4ghihli
B+OGdn0T4GHImkqi2xqoIOTKYCnEsP/nInf9wKNBkVA/9meuVtYidHS6xkFTl11L
yFin+GZ89zbxKCIcGR0t/Wlgzkr9It1vVXg091a6xVa8rZHQXMG4a+WZMlihE1mL
JbjRSook3B51wo+Uncu6jbOr6s4i21tfAu1SbRaGU1hl8McAspRjA+uTdt/bqOLS
/Ok8VJ2VB3OziRq1yHtGH2d7VL27UE/mQWF7NWz7U1QQVOt7TcZn8ZZ2qqLJGMtR
kpDlsiXxNP+fxMaGhAOwwHrjijq6hs3JUrgZ/tGzFHjZAcIyw3gIzU8QIvu6S42e
O0hDRgmzMIfyafQp960VoyJb16qDWmNOBkvrwBMPqrvuvDH3CHcDzu1GHK3sy8PN
2s37c3PPrQZ1G3MYyW6TaBwHSgDtF0N421eIPYEBlYugTsMvR4nQivPmYWUHcioC
lCcHz4VVQ3c4KFCQ8EL/kfvKrDUj9Ots3Jsd1HKaOpY6frTmAu97ePSZV/iTK4xn
rw4rjSlzFCopmzBU0gxawNRHgX5yw1aWq45C0vV85kXLveZcpkK/ZNPDNclUJgXA
2PPu50RBlUDP2GIMHNMogSzC5LsdHiWq8OCZa83iGPWH9LeBRiHvJYzjAo2Cgk29
X+H3r0oZ3P5+GX1qib916XBKtKZpBatsSaEiTHTFo0JDMyUkmZ8h/Mxk4h+UeugM
UxJiI4RNLcI3MP94I+CrcyWAstdgkuTbIs3hT1SAspKoTqBAsxWv9m3kzznEzjbg
/XVZ0at2Gnzlw1p/Oimj8pexrUlqT77oB1eeGwJ2dEBa4DpuqS5gfVw1H/AGWEch
57SwibjSyf9cmyhc+sYYXolEVKe0f+PlM6DK+4gihJUZnfLVOLKMrT8bsBjzgNYS
Cbi3NwNI0ySFt4lCCbUCo5JLWDg3PI+wIhS2XHzIxw4dQ3MbPYtQZI6iMOvJPDjz
2d9JLUcsu1V0G43kOAHbaPpzSKZ2dn4+2GmI0caxKBp6MQCXHEzpWW3OhPTWoZdy
SFl8206a+1/VC/u8gxF4i/vdGZcujGrMETaTj5g4jm3NDpzTrtN4aztVw3/BTJns
dI8KMrwSY80gI2U7Om2U0+JI56mVyKelBYX5e+x2htQLpm/F4HWLsUZoiJsKvMnO
+XxSjLjr+msUUK6EbDe86mYkyLS6mquhWDN268txS63cwhpRq/PeJYlcAh74+D1u
IYwRDZPy9W3YO3sFpax755wVtJSwKQIGptybBaoxZmrZJQCGigGOMjf4M+ADMR61
1E3QRoH2bSW/tfK4LeMRpL/uh2UBSB3kDWcUOCq6VOLTNBzq+dIbu4KujVeMlYXp
mxZ5ViqzfMobPhzZKIwUZdi0JYasDTYUmCz731LSltdBFprkcUUgCfUZaqFMe8xo
sHzKiWQSe68Sreh62m88yK7bsF8HpVNfiecd5lKEhoIQs59d/MqTEPoJ5t4xBQ6F
tDYsg9NghZBc6wGsCo4O6Jq2JBYhSB9NezK/6WMzyVLbWdqS8+LUyb+XF77g44PT
Ds8zNuUNKJ6koAu6iiklcyx4V+QKf5lAOY3Cq2dAFkyZ7aYUJHs0KQpU30scWVlf
gPzrz0fB7iWclK3uUv56gHSl8SHSAkQhpzM5/w5XJAl3AHRD9hyB0UB6Pw3NoaYS
gZPNH2e4sBgLYas8v05LDMNdc/tGUlTLXaGp2rSwGFV5GXS+JQyY9zfpeRzCn5Mq
LRo+zR6g6ksZMbYY3IQ4kcKGbpqVDd5BfPdHBHnGWtVlY7pWtUvrArDG3Sn0RLYl
qVAqTjF4NVF4MzEFlFqRWyfS5MqbxNZePYjbIJpTaghIsk1v8jN7/khFsIRpkKvk
z684JoLHxDO1c0Fbv9TqFDWMO3K3lKS4VVND5eeJO2Pkdo8CRbC8V2Yi4cMp7wIJ
/i0WfKDFPAy5boF+dDmz6LxchoMXTcVnL7eWGhJ2POmzmNPkecbliRIN3uOKWRyL
o3UGdKn+Ro0/hhQaliMS1C0f+TdrbjoltWeJbrb5P9AOhnMpiYP7CroFSL1dY0cr
V6Y+pUikysupeOoFR66Nvvc4dN1Anod7410csIhBW2gC+daAhhiJM50tlGfuikQq
XZ6gsAfXDZhY1XUMJyb+ZEfGa9hbTlMtMb8Dpfn6tXBeUQH6DGeluoEqmh+3ccmL
vzDHAFjlDWXFKgWWGIRcAHNyo8SOBAkgBkY+tfIo4iDCh/o7nJZr+mv3dIjArHuZ
wcGwdX8AN15vpTckiXj6FB44+5hiLiofDUdsae/QGySd/FAeO16TItT6vhsMVKre
0+KFN3ojd6ueVKQClCs2O1HMhlBd51FpB7pZPwlBimRwgdLsokuhaTUbbJa06G2R
Xmj1XDq56nnVw6iILyl7+UBj6cnzmVyV/lCeBxUIjU7wpZt34H0Kb8zUeIFL6NvC
58Ijo5cNjbpxf+VZ81KZJNtsvJQDYRD0y9pJn8A4lqaPnu1uTyUP/n22fTlNuys1
CnQujG1LouiUD9xfokjnxPR6lmQJ1yBos81Y8Hdx0Mjwd2A4WLjvGIUZrkNc9cIV
Qiyq4GzV0ddgehLFBvfFhQiauf2qWOQ3Pu56zzu7WvgqPdVa+WSAWPBo/HO9aXid
qNZULC84vA0ntHnM9//aJqih5p5oMkvuAhC4hDADHGRnN3TztVUcox+dWVYKUvM6
QvQ3BdRBVHXEgFxZ+4fKY4IHhg24hXVKnzaVDTRQZMD5jeE8yeQVsHoJSyn5jkYX
OOWLRuuBysHltmgWqWYzZG5Kps1WTWVMnwM4rWFxS2qocTx3MriTIUbEcwo2XMLa
MAj37K5SlDCVB4zjJLTO1kiFVX8fOMPjjdq6wniwkSJjdrE815Rl/acYpye5QKu7
4wk12sLFL8FOPgWII67WzIOT/6nUOEQ2PiiPXf5GDd9VP+hM+sYS3cGPtv2ByhWy
/1yeJZwNIUC03mFiV5/wi0pSTPI6mfqN8OgMnkSk5o8hp6b3e7HHeA8zL7mQu5Vt
zABCjnvwt6DnJeyOBWnVZCNk3ai22qc9ZM+3d3D6xs2P1p0zCmWfxU/SdqEArbWz
Go97MpDyhG1Hsmoxg+vugWuVPquRUCvk/5BxT29dm+HC7DSkrWJ/haFT4FJX+ibm
ZI4HsTD8QF5aYAkXJ2ukaIXM9mZGcKdwCouUfYCRmxyvnpF71vZU9AR219xES25I
iiFqB3HEiUWLQhxt0Pbxc5WMQ9V0Vyi5VPmo2F5+UK15/c7a1hS8NjGQgzNZw+A4
hy/FAoTsQtdofeibprkmjyk8UD5G+W/7Wi23B3tLFYMJOD8cU+kPcxG2Tblhe8nl
zkgrlntDsIWpZYBpObujKl1Ta0AyzJSeaaM6wLkultGZDaJH0kf+56nKj/bQQywL
648WvnRqZfxzRectcCxSUdv4WnTJPXhKJxnN8i0ReBBYUB4YyDnZA8t2igWV5eg6
GEBtakjAx4dr0L+3sIHgDbGqcFHS1eK9gQLqmKCHCeqxQ9eDJ122GAw+I5sWyVXd
nCEgufZoN1N4AshC2mtOECeKyRdR6XkARkzocavm4ACCJd+xFIUSLVsBTgry1UJu
w1z2Bg9WebYgW/BnzRzPWdLcMGeg/fPaipmWHyoXzE5FFma4SVzggdJmjhFRz23e
cUZwnhMJ8CyZiiLJtl7H7CsNxXUDRo+e63BbKWq9Bcw2G6zNCav4e7PHZALy/7bU
9QMSiV5PwH/rslHGFoLrZPOexywFHSS8i0XxWpgyXyiOrC/H2Wn9aXJFvMCfCCAZ
4+tOpS7mKtpsvRoPlWPnycYxXwEvmeSo1bY1L/p+lEvuOK7IAbLxdFE7rKa2YJGB
OH4o4mxj/Dq1nkhNp0zJBoFenfBbwWpneZBZx91jAR/STuFusF3MM0SlebtGaF9p
m5ELJDGAkuMgr2vPpP4A4W6hbx5gcm16yfKCYN+p2wMUfIQdJFoLFmy5Otge7pzi
USwrhN7MjCIeUnpgPmD5XEe5CJC7F/k8iXezNJGcQmeGO8cIt0l5P0mLxmIDYAbA
NmQtWEiDDg7CdYbjK9/5WoJeYkDgrQseAEr8KS+8rLrDMuF8ZvwhEBiX8Esqei0r
AzH5OIqpnjZynfvO3T1HJ9iFKKvhJU9iyWWrhNgcVwqbv4qbhlFc9PlEjCD8cb0D
AFL4oxOKK/fAcxnV7oWVhm2T34k+z9tkddrPqWlkiCtKUgSYXwoEUrrpgkW9jOhy
PVLpJeMTeNqEuvoUGej3JOTxeJEwvoMbOrM+Ua9i3zhmEB4hrEDfcXC+iZAfHgjY
6sqGO2XgOR9O9STc2fl+L/MMfw0Rz2KIOgwQpCBxIHCF40xXPpMFttRkGDwoLQio
FzyHdk8twj4nQVOA3VbDa7mmXWpVP6FNtoWTaBFnRHqzMmLtfN2Cpc23SYnfUZ/p
rgTG+Cld04HzZYHO+mYuJfM0QFpAMjQA6kCfKATuORWjSKtVjTU4gcCQyINa2ND5
Dc7MPozRfE9jkTG71fxsFHtk8WsM6scVGGrspcuRzR8I2yiZN4uvIS0NLexqhZTS
QFGh9C76ej2oc3061MRnlOTLBVCRmvZDemUypnI92bwVrBNcURkcO1ENCbu09n9t
meSV4CIkU4ohKSbj7ftuAr0I548ASKXkHEU+BoOwbe8VvA1aSBGGsWtFYKOMp7t0
A0Kl/hBRGmmRO7oW1+IroqUCwF+YKWrCwmCJTLS8jbL1YMssD/KTwG4hnkkSWkA4
eu0ZLL2e1lI+IOGLJW9ZZ0FHFGVlHXv7mx/EZFUXdlueDQIT+oCr3leFpBgcgcEY
Tj/4qnHhlYdzV1qQfmvz7LySMUk7AYYv+t3xTJ4i+qKhtJTw353EG8ATDDg0hfMH
Hcu/BJhPQafumEt18BIgRARtQqbqf4nQpTlD7Z0XmXfU98yf/b/bmVCErUflpMT+
9PVsWVVRPr8069M25RrjJN5SqQjTRDWvToJRof+RfjlQx630DKPUKkyveD4qfG/X
XXLSJIPpyI+vRwwJsggviQQMxg63ZC7RtNYJf8XltxDVgXPy2XJeHUsr/PnXzy2R
pWP5lUydurXz1sVPPzn0lOYkPloqkOSY1jBdRt+HHcN8ww4oofkD6VMB4EVRPLH/
K40/NmnZMBI/XgaBMDtBEmtwiOujrCDTaRI8bTIvVMpS3hx84PRVpg/KYcW4ObKg
Sg/lHY1NeTWHfYOpi+7jfgfGbmac6/+5pSa7WL4PMmvjbUQtZs/W6VLhYzmXQtBc
XqKtzkK/dUu7EnieozNRKiAX6oTC+zr+i7zraAAPGuOA+G6vW3QLkU7moj/FfHNJ
IDNnDv8VnTvUWbLCJw8NPPa+WGe6MPXMKOGGwksKeRkCbHez08dY9LVFfiRK0diI
2pbb+/5bjaOGggNh8orMaK2NwvPNR7pPgXECWT53sI43qt2HGEuo3mkYcOHYLBty
G4JmK/fyul88G86ocI3YKSo0DlFXeEEIZ19A8l7FnIpBSLDtsqw3pmUETcIt/Z9K
ZnpTWsZ0cxBHVaGYoQO4Fm4GvudYfOvougXxhiD+xB7Kop/DfG7Sek75lDa+1dXs
4ZUz4gBFF9y65kssC/BhjN0vQTigMflqJ7TePohE4PRKWgQUwL0iA5dkfABF7f2Q
6S02SuKHrfyQ4FdGSVv2Ms/VJYfyq4xsl43i8yNkzUiDArhWAnPc/NfkNTazh50Q
JDg/xGY1vhE18Q85TfxtV4YXYarG1sE7xPdL9r47p6SA0k84jKWxXMMDF6vEsoeO
lXR+IYz9fEN0UgFfrVmIRIWLo1cAL14B8pdC2HqOrmOElUXrNVnSYNq9qZM0mu4r
kG52dZa2KcYtTLCiVoYP4cmjBFHhAqkt+IB2tWVicgFJA84S3ZYEvtENPXIsZHW3
aJzuyx/Tg0SpyQlZ92D2ZgqyncqE/w87t5wTMiTIxn9jIFGuJbQIx5cWmp1ukua6
onzqusmxBiKnIQQh5albd7HBgwUodGJ1l/Oew5kFpT9nrI5AMFLxJs0mowhh3BmM
v8qcMt6poDeKiuGh65s4Ah6A7P78OONI8kkyjkeD3m4bCMaD30MCRTviOK+gCGNY
8YZXG7KoyqqIiq2anzYeAFNdmMEZlEVEY93pY0L9XSZ1vwDlcFQhMNefTjGYwWOA
fjJRtTBcCnjVBuCyZoZTITX30iQWJW4fAsvhoSRPvc0okfmMq6c3XDjARCNKi4Af
TW9HfYlPtprBwfsnMZdbJPl7i5cgH6heAJQavoIlfAEYR+ionkWrJ2V9ezserQbb
MDTjttA89BMmBwxWyKpBIfZ6cxeOEa3oYl38TEYe6WhsKj//sUDVW+qvdn6r4fHq
LyL4gcF5psK/TFlL9dKEhArjcqu2CjpmtQtfjm49U7uNfK5DWEXXTJ2QlIgB2naK
HRVTnwddQqYOB9d3f0TiqA/COXj4ymkgRsu0dFaLZLP8DRoR2hPlD4EC07F5fggH
mvcv6vRytVvGzP1803+zQS2i/bUp99wNrirAdMXTe3QrrSg6YAil8ghRHRT8jjmF
UXQJ4nloCrZA4Cjnpcwph9e6V925WaWJxDA3pDmB8J++IUL8Y+5zloYQ/lVhgxk+
shibJeAcFkKCnqXjd1ITAF44IOZoaZMkmKJWnNkdS88DZlgDhGHXxRzzhoY4NEro
8//zUR5pdwFkfX8HTv7SEemBn4VpFQNNhPzHxvOjkh/8E21xNRpm0en7NuPFqw1F
cLqN0T5lfC7XTsfIBxRNL75jwKPBGLj6h6DKZSSbC/iU99zmE8hcfIxmsLetk2BK
DWtoPrqzU6jVaiSIHzcvfS5s60EU5x1cqqmxFFukla1EAvU062N4qjxqDU52Hw6n
Ln6c05ZccSrtKaxE5hB9gDMYGQSwvMTn/4Jf5mNJ0r+gjFT2YwagjT6zo16pqSQC
zCIX86yiea2mOTzN4NB3PfOEm9Uq6Y0krC90ywQaEBD21bJTg7GGjSHoKbPKfKuQ
IpjqMxagBuNOpQAUV9gw3Y90vSY/n7ehQhVVDP07CEZLEzbUb6zZFXlngRmHF2EV
IYyg1heMxaYSBlLdOp4v/dIc2zeTXbdE6zTCh/qklCdGUY+uk+C3zmfJzoXxqpZo
6a27BbKloASMsjXdbSsSVDaAdcJfa9vijiMJ6eTHK3kk0aDvS9keYp8SRZf1S0+v
PlLdbKqHK9E86QKb1TYw+BYMPRuO7tDNk++S+BpGhAl27b6szYEcjMscrnl22WN+
u1df8jmd+arH+6nHioPj/zP3S0SC5c2I6vHtOMZ8SPql5eBed6aFJ0tFezz2GjDC
L2/RcPWFEvIYYNSnCCpfJubC5fazYan/mk/hW+orAU0CiRAbvDKB4Y/1QrEGdghj
jrkE4oBjfAYIeOU7U6je1syfY/ipswwgjQ763gu32YbJEcL5qzyLxMKvhvjk8enu
w9omn3yxbix/OewfrsVmj5Z65rg+EXev0BWePsmdld4oxJS1Be6Vl3svs4k2MgOX
AR8e8avmUOEtoI8l+geiIMqLJrBEUjQZX2J/egq6+DhyMhGKaMcEi0C3MXzOpe+4
eZghf0LaKrU+zrLx1NIFzm3gaBz/Td2xcKrfqnDLv+Nu/hnjV3yNFeUzoqCV6lsR
Bd3sWEo4/29uSqu2UqP/Lddty7EWv0NighewxMsAy+Ea2eYdwBKoIHug2Bv/A2Sk
NWgxlHiK2Mm3aQdVBG5dY1Xf+KPADshzkucEjrKqGn19IGdE3i6JEFSFW48gFc1L
Ps3+MqVsQ6o/I6lhO1PbpXeacxudvMAZIdXDMr6Bcn/D2VKZlxn2ESI5vf168MJO
aaX+tkRtJaNHwlgay9TRFXyohZwMCOCUMDn4W/GmeDjwhtNx7Gf4lItP4r+XVrtJ
7hK/UhWUr7E1DfJCi5cGpHTQLJTNBRSVthXxFF01heacU7MOaDXuUW0D7o6hT3L3
QTNVQ8ziTxmHmftCGU5qTFqc3guxbB3R6bHmq9ujAvsrUF/7SnPXA5FlnxMQ/WK7
q9RILpWQLEyGEN2LZLVFtYJXTAPqurFQ1GXwgAJErWxkmQ5hMSsK1N7rzYi0GMdq
nQ09Att83FSyLeA1BWHHtg/taCKUlaWZvE9Z0n2aYNoNDXLfOkecpRrx3qKpF5sx
+GMMKUcE9NuR5p9S7qgvWYF42BTjDUbVIkZasz4TJVLFeyI5VjHvc/vEcidys6ok
VMUnXaqc5P5tv8gkODm1yvCCWOiuNxqLzO8W1tnCcOVKoIqJo3EAWnFQ/k/noZL0
vXsYL34TcTJlVfK3BBGnzgFIx9Fjf0djyCB10VCsMlzJZnbMFoJ5kljhZ0wYfKDh
arSXMNewStb+/Ycdrx3xDfAwwAWY8EyOld9rDXqLnR1nBe89y4fibLPAdaTaUg9J
ywqJ7jZ9bH2CcRSbQPb7ktfqr9ZV3nT4bdkTj/bpxw5jEInrGe5QCqqEzdQoQXkV
akFSOGMu/6f+DNnUtKWJKOTP1d1nSXLnfxMHeIXsB0pMr71y/nnkUchM6L0b5Tkw
mAF+m2tpCV9zfjBjfM1/A/Cbr0HmsBGKwOA/TwByzxWxtjucRSAPVNhWCymMKCf/
iSaP8heQc5H+pFQVlNACisp6kj2OEAR2gttKLsaW2/O58X0nJ5dfJntVFL9uqEaR
uGdHOPKOye7mk8AjKeqEEzWybTb+WRojR6dHq0hjyVuTlv3eySm/kW3ITYpqCDf3
TZ8ZRMK+CFLTX2gaZDOyBC+JeJCFRb+wiZjSyszKHwAKVyUvGET3HjqdA1cJtcyG
oU7QsjTNPoAfdH3WfDIPgjFlP7vz6P+o+apux+TsHoPh5wkwI2tcb0Nwg8mEuJ8E
d1v7hrQWzANouWQZh3hnYDP+A0rcweuj1YQ382YRfxzwlX+bLbxqcDliYPr39hhi
8f0eky257yAlNis3NdNMbAqafpjZeYzjdKkIhZhr5iZepuVE5PtPQqpS/xA+CK+r
9lzu9zPtc0S5pKDO2LcHyt6wBY8auu0WonIcgbuAAVhZqP9XRQhNDn641wB93o2N
nsAxvfimq1qv+2WDdve+29EeyVfe8wA7uDceg8rZLq2KTw8CbwbcYSAL8tfj0RtQ
KuB4oqTKWNdj5CKlSlyHfBklg0UwFblbW34A7Rr6+1hDHEegSeOzgI03K72p6W7R
Cwgt+9KNWs3Sld771F7u3BNZ50ZsaL+9WaOHUpU0AkqYt9Wa7TTqxNm3qaP3XWgz
0WBawSdhnCEgJU0OlWBK2l5O465gSWwV17zHWaWXRmrfHvkRCcUL2q51kNUNkdS4
YCq3NW/GQ5jMpf9pnWc+P0G2JCPkknUBDecTFRdnFIT4X2N5OvIFMLy2ieH4c8Lo
MINFMjg1SrqpY980jhDYimGEygu+CiCIT+kx5hwXy9JND4ZPabdnNt5qSGNvZT9K
m6QlX+H2xODQyBFC8zQNzTXhrFBNGmSTI7hVpb5hbPVlcZ2dKw/2TOq2KEhztZFJ
AI5jI9UhFqcbgN0FAsbE2ZTV4iKMTnIBtE+EKZvL2LvVBJlsuDsOczNoG/xyYZ0e
dn3esLJSzFFQQMepgHhITRhh9ZTKlEgr4SOT4HceX5xzVjI34vr02bzFvKR8iodk
5+aNzD67Q8j2kxuujkCDKu5iEHkP+3fFJXyqmo85wT73gymfWSWEWc4+Eb+qI8Si
h5iTPGglSqoab6sZ3HvVuvN3nCgTGnzXAhCXUYLn0q+kAjjmG6crjPfjLxeOdZP7
GfXhskWvnXyt5BrLGrMQV9tDibSuI10kOJpGFjE6a5aabVOxMbS3r4Fi/si7T/2Q
KKbKQqEsyH+5ioCbI7+ADRw/0YWWwQhTZR4/8V/Gj0NhFnP1STFBGQUI77oCqPG4
VqOUvdfhJJIQfoaqejlPldYHI1t/yDvxuy0m9IgIQtIC7dYvODFYh3mxbirsHBdp
M9AaaFCbScvM1NsEEZxwp6ekrxf84cvwj1V/8kADpuLST9fAZaW1XBF14+bOmfrf
eapefj5adeyMLH2MheGHcugvX0jlyvpPoR+QRlwSa6/lWQKo6VFjQS56bTaH6TEC
UR3k1NL9C9cozKs5ZjEHGevbi9TRsihVpWDaAMxIzHbkEePR0HCMqhaGYj8yai13
94wvmZPvq5Oj+9Jru+S6V46M1VP18FziAWx10KdFkXfnsz8gTX3s41e+U1zwd0H5
nhqsnky8Hx57yyj4wpUBj3c2sSUMF4mZHCsJnKNxKFvZ6YjN/bhWQaA4shvX4pVN
ZKb2R++4l5NTKryqitUSH0biPqv4daJAh6Dbiobkj1XXQ41kOdq/QFwitNd1d00X
z82rNixmfMjNqobLS7aD3ymIh4XbWycAtao4lbmZUZudUpt9Ek3bYcQSAU0f5qNB
JWVXIHbGNXWPA1cd6EsIVk097ii5/ycxtm0E2XsGw7hqh0+qhM3YqXZfUfEc/Tf7
APbEDlgsX6LMEhx3OE4Yus9It74/h4Fa+Ap/6bm1z1bPZbSzqYMILoMbtDvYUpba
NNOepT5KO4XJhFFZAYBSNGFNB6MD8D8OzfijbohbKmfT4yhdJACs745R0zTA8bqs
OOVqFToMZ67rdhUXJZk+L0o1SJ6mKQeJIEZfuR8CxcRQZ7/oAIObDWvIpvW2aTzd
xmfBKfQokXcxmdO6NoeVaioW6VcnSJGbO5mGmexY3u4i/BhipVPXX0ub7m9VVT9Q
vdxZlSFS3sMlWF8+CXQ7H0b46yziDKw9YV+ngV49kdx2ekosz1lff8/Mr/x95337
pazEhtIci4d+aJ+587kR+dsVFyKfJ+TJscXbHtID4IM12AqbCyOApDYNW8VrDrb2
DkZhHU2kKepq4duenuTgZCPCWsKeOcMFv2C9FxrfZJKmXwaEkKtF9I1JDk+ntT57
3q1R+exKqKx4MLf6nhWrAhbDeS7evmGVFUt3GXiBKkWJoJhDm2KByj7Su9MEwyI6
un9G8lmSTVW3ZEs8ZxAD4Aw5pmEQkG1iNlEMsZ9/EJmbvD1BqfjDb8nBrfiyh3/n
8kSGOjSP7rjaNZimkC1fVMcRUMqRWqNOA9QETgfQDTnkgODZxCPWytRxXUBQSLW/
7J+JF1MTIcnBPHy+o1zQLMeXrgy8E3fdPCVna5n4x2mKCVpQkmz7qqDHTdhvUDlw
GDD7FHbzWj9/rSEBSQUB5tv8/ZskMvfu0nuOGZtHrNi/3RFYfQhsNgQF0PvXegIQ
`protect END_PROTECTED
