`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OiPM/I+LWY9xC4AsAimMM3PUfycHUKnPkEDHihfXAw3/FlcGIB6vAAe9BqaoOAOx
yvsoDTZkOyDpMlwVcEbFzvXbAFhxFKUG2zePRB2MXBjXXoTtqcWUKOnW3evTjkOC
DaybQL0uXkdrEvdPYKeOm4vSgdX33LVcoaWsDgGV3s6nLm7o+XvJgSvyArtpNRqu
4d31cyJX95dY1vaaBMHEzYJbWWiKLcnDUTJLrvSNdw87GoVPOtojD73mt2A0DaAW
BKOci9U6WN9DXm97XyvbGc7k/SWh8igVvPazl6z9PGFmQVttREM5cssT3vjNi/KO
5TSa/zZ3rC2d8JO+Xj46AbdxgtLnDPs9sni4manPLIR1i6Ewq9jNNNiWvVAhi6c1
ZbzwKp6+wu3YFQq/YpH4b1YcTodzzhNpWgkfOTnDmlGmvyEGb07WACLlhzzcav1O
rDuZ3g80cqJw8lrQGQqi56bfm/mGXxda6vnYYi8xiTswS+SNdRpeUG8Cf8ifMi3J
UqbCVXjuuCnp324dW6AncSHtbuRtrX+j2S4glhFwN7rj0xu6qSpM/+RDpWe9v3Rp
YLbi9OT72IdBObj/hg9zdDEJ3kYDvPjhUpuV0Hj0eN6tuj6Qgk1LgOWZW4xtl7Zq
jeY1P38+K1XkWugbYzrV4EzooE0IbT5T8Zu3oMc6mohke53uRu9onfnScVUMG15E
1PJWHOvCSaKqGT+qJK6kMBl++UiU7d9M907D8LGJDaP4GkyM+6VZK6fDagGgZ0CD
wDyFWYK4GsbZVZVmWNaLha937Sjyd44CGGmxzRbnd7QYEatzSdlNXPllbVN2X306
3te4hC+Be+oIYXCWggTPJn2GBSH5gaUv9pnR1H90Esc=
`protect END_PROTECTED
