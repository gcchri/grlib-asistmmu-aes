`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dKVHhoqxpBOxFrUED0vAaz1IvbIbc0v8Kl9wLdRE41CmnOsVT595FALbjSHC5KKV
MURxxUjLl7hXrFR9ECfwI0S3iCbV1nS+HpcXbVFkJ7kXJtwFC3HvxtlmEk5qnFCx
U5/ZXwsKvAm+dYhTp22WpQRYp0v/jvm20FDemxhW4YHi/oIDFaDllS7sDRPIAaXj
0Mhc0NRaSa9heK/e2IU4ipbkqUToloCzriljTc2gvxXHFK0ejPjzFzdOmtH+CLH+
cvCni94FLfW37WIcLYMtlQdz8FtNHggrmsIWqyASkt5nSuI8mZx/wk4lY8OhTdg0
vGHfQbb3b9YMNDfUjdN4tFccH3ObTlSDcrY0qx7WVP6nkmuoEOlhEl/J+pjXBbNX
6xZZbGjczub7FYC0jQFFYUr8tQdLAjTR+cGnk7FP2gtnMpcMJWds9Kd9MM0gNmUt
ep0Bl/rQL6Bbw3oPb066f8XAE0/SGAaRZhnA6NnOWnePCcndBu1uOrUlqHX4/brz
`protect END_PROTECTED
