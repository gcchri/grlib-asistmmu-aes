`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gL2XIHeVlwobpMbAG/gyZcYSABfHkUS54XvYQyqlKUy3MuVx7rYXk4fNqLmPmEA3
w6YDsdvG/DHY/0cgNHMPR7GXrSzpUf77aTFRa+LHlH0LLEsCfkyQOsdD/dfBGahq
Sm+bErmaV0ML1Nl+nyh+sROL6jTF4RjYquvtedMzHFkE3ZaX4mPJPybJvT6rg4uD
cUary4Ox0tfB3pHQbBlzxNeCKC7imHbJOF7vbxVLVQl1VGAaVseNYltdNhMBk+aR
2YTkV3L0rH+Yg2lCMz9VW4nYRV5ELVeaJuSsgXv44uJN3AG4kvR3blYOF3ccDNbm
/7ynt4SA+7JXHmEofuzGE1eUAOaBQnLp6cb5vkUGlxTHQpAIRqFDUxEsC5MUADbE
`protect END_PROTECTED
