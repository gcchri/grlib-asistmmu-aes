`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kPZ7JvT5F4Ye/19cxuJ1FcRTHRmZhms1vQdDXSd59AUGHmNulZqACJ4VNc+zO/Pp
FQvCUK1Xpli70DfVrkwJxsJ3IQnhoHWXCBY/1yk3MySwRvE3RfhVXyOhqxSZ0vW+
TqdoLm5bnkzDOMVVvWhRLlXOuV/SnNqQvQVEWh4+OuET4twFFHYAiHSGi53qhi7w
a3apWAfY5foYf6RdbRnghDR0LXg6Myycd13gIOibvReWBJrEkNrzNUaaTBBkEPKv
63rQSdHT0nyM+buMCqVGNUcVoFnbcPpCFOyMflLPBbeP35LItqMUgLkeW5MP5Bvu
uGlpqSvDVkRHedgE+uxra/L02I8Pcr3Uj29dMN/dD2crithcm/f+jmx1fjiytvP/
p1lOiL46nL7Hn3Pvo0IIUzO//dRo7v8UQBER/+BXUpzrRxyNs5EioTffnAIch7HN
Pk6Q0oEK22/O+ozR3TJxDAxXzUeftTs9bss00VmJ9pftDNPFZ6F2AGDZDw3IN/2U
8rgeDRMzaTd1Dhu3z7PC/KTtguReu5F1ekxjmqQnr7BdD+v0hp5/p7ga2TEmO/AS
5oUH+UOKnYGneL7eISraGT3PcXrGb/YXSTzyEaM+VZ48hT2lHOr9X0d60i2xT8fJ
hOuelK/58/ZsxPyM6ZRmBgnikACONyaN9KG7LaF2WfkHwou6sUtr1Y8zoYGuPK7T
cvtuyyC/w1DTEelG/fwy7lJOAkrQG2OsUJRI0jN92bmkeJNXDgu3kvrIaRldPtqv
AyI52jrhemWRM5+pf7OsyAdIVJDHAEeKg0p8gf7X/V9uLqd0h7O3kPCgpdcBv4e7
Ph1wlMgH/XZs61ZE+hZFURNZjzx9yW10NxCdaEyoDPFlMHxerXkeayaHzS3ge4yp
+DwvIvUdcficCybVNbVI5xg3S3TdobGyGWhoA6LGusvPbeb8aY1fKJPNvRloEISH
MFKKBY/plvTTqgCR/JFWTR0NFeZpA6GrcobvmujoiDLd6AvqxAI4rYi+4UEmyZZK
g3Sd96Af5qdud3kT1bWoVnyhTyRDZtpmw31sDs1x2BkkBXoUsogEQPadB/v6G+1J
cM4XX1y8jec5Zmkmq4ddeiGiEBCH7pOTbgBpJNXW/e7B6G+qESmcC89montckm+h
hj1WirUv0Gj3IEc5K9kuxXWtcrcZ6kWsj5C2Cr5O9KIRkUjZW1huWVE+yfgYysnw
ykcqYJ7SZFKomqz4DK1mU1XJj4gO8qXrxh2VKvBgHxddkf+VzUZKGAC6c6qK8Wmj
wTJm78ET4un6jTMp88pxiYwqp6cZ9GYQS6Fnz87s/Sj6/e3Pap8CFxobf6+YT9QP
Y0VAeCgf4kDsUklibcTOWcpEDoByzqwJuYnClAAPrNvJediPGEednjxvYl5Gb92C
E4Zh3fjQeGvlWprle8INILqWM5CXvrUQ0aQnVFvgG7OWFdVGV8iQ1sULLAo32HTp
8PdftBsnekPLXjuz1paae4edG9RiJPeOQJobx8sJSE5vdURuXFjiq5lr6MPCictE
qceXfi5GTwDe7D/CDzV8JAVXVvpfDF0Vrye3y1Ee5G0DicRvsHqnTADiTubkZW7L
M0GVa2dynFtdfieKeL+oacMNwZi7buyuXtuwOoriInhiV7Dghg6RKye2oRo4RHgb
6kbhIgaN/RG7LMAMYavbJLG0nlIyfWlyYu/uqiV/L74+01GdkZoV+EkmoY4W7oXE
q1FQOBMpYE46uPFgppQvt+SDufzXtTRiwFx/Ms9SI6LzJeiYUCU+x7WpPaiHw/Cy
kO9/Xyrd5uTi8/qwMZ9HSiDxymWJlFvfwVJ6BIv/OKSAlk2GL6ATPJUnAbhFgm89
i5FAfedwkuo8VmVNt5g9fzzEnxR4A9qTTp+pIP43KBkUgCN+q0Hmb0oUL3bV9cJY
O64pbQNPmwAcKpc7oBMVmNE7GrVVuuTMWH3+vcs82wIyblBAwxq778tBGVcmQrwH
oob9bwwQ5vyotzWDGUDPOtICaAi9TAku7fk1d5E7hHQkw631Y0LdqhouGnW4O+VE
WFhyKwF/3xdTkq1XsxnXCVfvuQW6sQZo9bl4elgegoZ4hp3sNvngHNFRjz5GIej1
L2+dlBvwo5cAaOFEyymBW4/4krKSqK9Q0k5rQP0bDdZor6Koer7HW7rxRakswOUf
7VHhFhbTFDYEnzAz6+oC2oQBVYAlqKU7y4dSTdbrSoiP7z97fzPKa8Bf9Wrnotyg
+Ctgsrlb+K3XiuDn3xLL60T7kr88zNrYAk5ef5ZNZU/b4OtAn98/51XW0I8C2Ypl
GpsA3JtOIJcl4lthyKgrOzD7m7bi0cD574KH59Vog1KL2+ugx9/2P9jgdwL9wOWc
/rjdYmaoUODw8dq6p696OSXoen886qewjvPBMbHovq47Xz4uB2TO2fvvrez/qvLV
kFyB+Xi8zEua/v27h76uFkGFO9/uGCosECs+BrnljxOpz/yRrUDeC6kzzXt987Hv
iOHAMgZQeopVDE3odE03vIKiEFp4TnNr+WFc8Cdn8mgkPSUoX77iapYK4P+CbX+p
8JvY+3R+Drg0YRcrd4lt9WFzFunRXtW+saY+zrWkpS7nmDosKktiN4Zh31V4n+NI
9kRUmF5R3s0O089c7ZoQlVt381xTK+wEao0KNkrGt1o1HPoyvEG2KpNbP2VTEEa7
POHJkBg3+KmUOPGOsIytsiDrLdj5L1OnYokG+cv+4sJd2rdbXZVALAZc2IUyNXAp
OBX9ssWH9Nrm3jqkQx71WyExvrXGKIwLEffZzer1982Xleu7BaJUgq922Zkr70MP
rxjEWyYx1AOvNvoC7eFFJqrI9dBaGBH/sb8avOG1834FvJVcExN58Zil7eOo+bjZ
iBXKONnDvEKKapeH/lZKqj439EhCKp7hHD7XszcBz+YgvO4Z9zOmjGexURoPEGPn
CQ//nHxMxRBifRnUkNOqKXP+bINWBE+Ew1ReMEaBpx+E+7MDPZVJvym2jARR63Iy
l8Rf8Dsc1owwb0RDDGI8mA==
`protect END_PROTECTED
