`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ruR1W3TzxS0J1mS8ffQxTVCl0xUYfCI+H3kneVFHagiMLMiDIm9a1I3Y7eeMK49W
oE4LAuFIFULd/eybmck2E9PzfB4SXVSAAFQ6UzHj93iIzf3YYk9MBC1QEGE6pz7F
8Q4XCM5QZg/rzMedoTVl0MjP36C7VX6nv/dFibET7UvSy2ar3i7MWmIil9QgKfwn
ITaCrBizzhhd1k3sG+qsCC9eae3/OgyedrKwfK+/dBGt5tQrr6HNT7kyoyITZ9uy
JmLNDKsTlJ5BWe77y0sZW8V3lBYMn89oP2fzNCxMTsPe2E6U0LAjh4P0qUf36IVd
SzqY2KzFFlSnrGuVivJVGM5/ewCAVQb/iRS7iU6y8DwpOf/PeJBrEiCvluwFay4W
Ha/809oisq/C0AONCzj4xyP2J57lpku9w5r/zmLcris=
`protect END_PROTECTED
