`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ix2xrda60bGbG0NCpAjWpn2Y6WZXhayGFQ1V19/YyXkYeqUPi1yr64AD3o4cDE91
+PgTWPIF9e3Hm/Z2qTrxCDPs6wT+SA01slVXlVczPzmnsyiy94JojL/Wr7iKWRwJ
B45XD47yHjMkGi/IGi1wunEe2TqnZtvE9M37W511u05VYPNuferi8Zxwhv9C5KwV
eUl3BoZh0lEdCr+owvPnP94y/6P5kjke8dAdksEO6D8Cdi9eN29By1nHMzOH5kgj
qskkYAhouaQlnCHz+cxzC9GIEVOC9TwCwB/IAh06xykRoKIGdvgMGHDTf2K7Th++
zT94xkf9SMltRGx+TTLLNo5Pjlo3lpz+1IHIVoABnznhmFwqkaxg9LoOxcIDA3VP
QWDscKqgB+nkRqqLU3fxFdxx03nyMp1HK3RtWzx4AfiLZzLHwa+tSZZ72iez5fg9
MzWRhp4DAtFYUGJuWIeOHgPInh+uEr3EXCg5xAy4e9lvN0BERJRrX5TeJgRyUdZz
QHDgDrIrzYnXxzMQ6olPpcDqCU5hQEsvyT/t+tbY2d26+mk9wIyT6x9B1nxMOQ+t
t+ZZwHCfaH/jFLhVj3703s90MQfmnvxVmj2CGZVFALY9RlJktNe8IIjdVEv2u5rY
PAJo1bnNSLFs0b0sqVsa6OpxZEmDD6OJkpnVl0q33oNo0ykBDlepvODP4bMc0Byn
nzKqFndjzk3nOCZjpg1+PJJTMNnpMDcFTpWAFQLzPJHM1e5q93C7dZxSS8H5Fotl
WUVxfHxt7uC/EzneFfYdCl8zsrVIKKQp69MN0XF1nVYJDiFxR6a1O9tHGQntQw7E
99V9O45shw/bybAwrj34IK/WbKzYK8iMN68UYQQx+/k6oO7PFGQ/ELToFv58gs2U
4WlXE76rUnuDAnh9LzX5MyVnxV/lWDOpIUjDqya4imoMIZ0emGWJusIkFgrVFbpW
gOJAiG/nV2CyfwchOVfmWhzXPZclyqXvYGo4XJHWHEf0KtiRWsG2ENBy79gVkee3
fPtyhvEfIJP6MldZPberiV0fohQEdsXPKXznSZ4hk6Fi/nsuNaBmzElgMSKR6bDG
hmNYTF1BofHD/n39xbrH1zjRuNL87HzjAL7PxslnwytdHUfUYb85FMt/vlCHcgey
Bcm+bN7qfDMg/IkhQfVunIQS0IiEffDmg6x6SE4U4MGBFbH0w4/3DDQuHtpf2sRz
b4Y5TJyLtBdHqaPRqz012nUMwf4EAOjjmymTYxCyno1xl/q1XdAqYMNJCtopAAcd
Z4Rm/ddfsHfjD31/ks7nsz4402EajLsvoQbU9nqg2UD+rLFNVsqU2B7iCrLJ6E6s
U6RQpBknwObpfBseHiqnLQUMVLssbVTgs6Tqhejg6VIK3htyU6ycckAN60/w8KhD
VqpagFZ7g8crUXQpb265p0bZbsHU7au2I32LgKTDWpTRqq/FpPwo3/U4vVVr/PJ+
3l7GSIC16D6uswKMFd/jOm403x6puzfAQZwOxHETw/ktLU1U8cUs0H15nGkwnjbO
HIsCiImO/wC2QHCmkHnFfG444eB5IAt5+QTLRPrP7LloHHne6JWVjvSl/xa+Atpd
kHAD04l+akJRXvdaDfeueNb6LBwWKGne2mf3YBLhomrIyMuVxVBO3rvhkVQlymqi
C6zclNsjOIZjmUb1nf08oFGLJWOfz5gyK+YxymyiHbHJvJgjYA2PXPCVAvP9VbY3
qcVPnGeNGwggiU6GXK6LQi8g8vxHpTQbAY7WMkmG8Rmq+2nKwL8lHimLjsWzfqxN
lu8CKRyGpyzLR8n8+QuDDpYblWKcpRuM+jrQAh85R2HKzzS5mDR8HkshKulzz3fY
CmwEL1FV8DtZpMP2b3S09bqdcVoDX3Q2Lj1Qm6pWKy0wndrfiyjZQDAP02vjzHGZ
NzCbMTzOIXi2D1eE8L0Dc/d2b7x/N1zvIoqc0TUFE6v81D3PsyiIZtjFfjvhqYVn
VpGQ1BPjdb3r5hijPcPZghE2Fm5EzxcWuHyaAs/iQV0lroZI14LiYoHF+ThMacUj
6AUJyhAS6wPKBzzodRzRt+BXLGMfV9DcoTrFSg/gBMqwPbxPgP2XcLQXa2gZZF7p
WF6gTUZOcd05g98x0cxA3nJObuMVEP1O+z+SpoA32nof2l8AglDv42f0B0aEXEw5
WkLYiUc/K7ZbooocIVEJ7+CAyuevwI+eiqthgCzKsc2e1fxnH/NBkTaqZ5gqACZm
oSZ/fyU56lACUKmdrS7UL0A8hYIPV+vYw4i9ejblu86NrjbAs8lFoN1Xu86JYaub
NWR8m4kAfceGS+EIfwepflaPCBxHT5UM9T8/MzjUavQsTsVfuVva1Gr1mT7nT99s
34UVOn02XKCS0gp11uIzQMTfAONlNgBUmAGE2K7qGyofILaZdCtS+rofLZgipmfe
KHkmSodh43fTnMKMvO/+REQR/Ngh3WjcK6vyDRJOD+UeK+mcLGLYJt1WtrXnsTxe
7b1U35IRpz7vLFEYuLCArhzthD4epmCcA/uIkEFlBNo/CWPp/Q9hfFljKyKQrB74
cxYXphShi4ixf4h+Jt2DS15Vs8SdiZ1u/HMUWEP7TgnswhxZDcsJ92H1Zm6ghO/s
2bMN1CxPWvLWHkoWwcm6nyddPIfycQqNVyKd7PqpPgLHGFueCpIF0oRBVZv7yBwT
nw8U+kRTf+OyS/CQSKpeOG1YmY8+oY9m9EE4JdfckYeGeNUdVwp/+/Ac9n+jSQrn
iN830MUv0QzFTMWPAl2xAzIGezDp1u0dqYVScwAKeb0lcxDcXofv6O2vHCO4ZzzR
W9h0s2IjhFmYYv2h4oa+hGprYkOD+XxPU24Mvj8C1yczTpmcBxVPI9RS5ngKNnyH
hcrpalNpkWahbJCwC0/ZBfkdiqXQ3ccGbPdxhJYmeV7FKQRQXKw318d8gy9ujfph
bzDewrADTgud984Xe/jkYhdAQDwBZTwJpDnu7x/mOtrklbbFBeHimO3pltchx/Nu
MwxUc66JmGVtxe22LbcmAQ8fuJhnvvMQG93Ont7/gBtqCNCDwquGIlGhxIzctvMl
6/R2sZkwxX5oW++DT3zmbfCfQQ8xd/s8oLkKrVbvEDcGeX/oPFPbYEurdvdgI81H
1/kiB+rQBB0jGqCcobiUVSnKUFzAg/MrxcAkiiT767kP3C+FaBKRSGnSerQrP0Yr
ddTCnZHmIlogM7wdbPLZuNPamLsgDMiAco41j4/ltAeNAqg4sVSGZFmFrIgfudtK
n+ngl5TN0sxi11/OhwkEIZoWeUZqRq+c8O5AXEtuu4Oezu224ny5RHx83PSaZHsS
iklJC5PPvgnW0XuoUqJGF1dzWA+lJq+n6rPp6RJPnLVlRZ9JX63shuX9zdt4L4il
YZlJ+ap8WvXtP+GWnifCAnOQtRosKlReNK1NaAU5TNNZFgzHVzgeQfmOVgmEK0XK
WsmRBtdH/qrztwLXTD5dICC48aWyogFyzIrvUexwcM14i6/rKmhdfcV35QmGqP0J
UMSYouXkWKWXTwkq/bQ/uScpM9s3z/TBsP1kxh0WZyVD0fCz0NqzQQlpDk08H1Tg
klbx4z+19CQmk/U96anTrACxA+Vcskda0q5yhnoWk5gBWlPShHPXkRfHjxGkHqK/
0QVP+AXtHtvlMt8RNreWfVClkEIY6oAKG0D45kSJpPbGvHdUUxdGMxz4lgwRm9wv
4ZwpsM8vQdPHxaKLVlC0noFMVo+fLNLM+OrLrsjmddjEm8yjXhW1AtqJssH8zZdE
LkSRZ2CPq50R1Vd5xY5BwMKxctNdTnRYF+dfY8UvwtRRyy9Nxt+4z6fbdbIhubVU
i0IxOXZaR6XWU19CF9E0gQJVgrFGVdWycr4A+VCkfQNHgiEYm0wGkJCh/modrEAC
I2vrsvfHfin2Gp5nC8W34uxCMlFmeRHoPDWP5rLKHSuuKSQ4DzXZJyzsviAd9mmt
sgSUOOwVwccShL+PxB3CkQaAe1cTFASaDCH43NpLhyd/USpCjtCcwk8gWvodc0m6
Zpw9hnodDMjou510P1p3eBHazNvoOZ65IY5y5njy96DQPMROsYgPquhHD426Oidf
skmgA68mRWN8yzuTzAZdB2yjKNSxeaTvC0/KfFaDultR0uxX6GJ7h2UhsVT7AEIN
WUPvavrSk4apiq3ZKYBueQUfArHsv7+ocvh4ZuCY8rd4x8BdhCHxOxkk7aJtBots
oillIQd/3ylgBpteUf8sa59DLWLp9ZpHiPs4SZ/r5ZMN/mhBI39sKomF2wkAeMrw
LW8XeF5cupvjxmqZBONCfZCVTNk/SoyyL/kmKOWnSQJqGm7Cv1lNaCSr9qRpSAvy
K9aej8it1+BpSuj422uB04uQQBFuTBGYQ2vG3cJDaNbWLU60u/7Q4RdXIn0syBdr
aCvmSTI4F0eQiKeE4gYtJGGJm3ixQ4zYYie27/mRTUTI1XvozRl1R4RDcUv0uWIx
X25SzKdnJM9iyWf4L3BupTvLA0nP3BeRGhiR2qTBK2hwxqWeLed9ZaiAd4xCwqPd
ybsB81C1PPSLDZpYRw1mlEptMM+n13NxaF8PDNLXujng1S/sM9UxxmxlL7ryPSE/
B+f5KnvObdNNWD+xPDPhxwTJMVSL2VjuK8hf2N9saiGp9+K6Z2JMUdn7e3QTXrwr
LsmLDN6D2NxenzD3NGbIR6XyTD/fitOJouYGaWw0jGjE8mz1LDijjt5xvIDdP+7f
uCHAuDhBavogL702quj/Ul2xYOm0UNkVCuXAsbbh53k9FnDxfL0gB22r9CeQdR2b
RQTi/qpe/3oUWMsscDEg6mU65qn7bIYDGOSlNK2MlYrfqND3jIHeg5AEb4/vJLWz
zDBXQUcU3Q7B8ZsuBKYFOZtulJzzx+vNmtb6LPqg6+HTTxuc3yo6xwVyXuNV/eIo
67yqhyQo26DirGczT8XlxiM7mGyDxG1jZyRP1cKS0/UR9NNAuLHT/iVEaU6aCBPA
U8m20IrYzXDNyOsmo5UgtHzQqJXCRcN+WWWyHMuxHPp2B7v+U/yfNhKPZWprs/xZ
/7AVGNymowUvwMkR4gSYG7rYQ+ulbMbyADGZ2monx9s9zdvjujOK1cwWReMii/d0
OOPYK6S7o2OLGaUH0R5K3gnOOqlWxgu49NX26oeK+22yE7Be93U6xYcFNNnmD9oK
7kyu4qYARgx1kCPUV4E8+7vXOwDt3gMGr4c22jxR7xlOGtN+nQS0Fgia05MWNMYu
PIM9qR0TyBMXb11e6yQvqxluWt9C2MoREIXuXcqazI5b3QCyhEydJFHY1QfAALZi
WgWizj4oICCoXgepqMsxSSzUQJaEUoCVZb7tCTarcq4rQQly+7vfJTrLUOvJSCcF
nOBR+wgStlGWAiMIWfXT3g9BkWCH5AUT/vdJDTrPVkpTgR8yw4WCx0ikmBMZ/ib1
LqKT7tmEVlexHCWS1Mw6GjHm3Zv6BKD5QpeygQtteDRw2bRrPTBCMc9MwOswrH4h
v3+oLB23IcUqEzmddiUlAGpDNLVyosHZmc5WOZPU7pqP/PFg4M+J+e+Z1XABQCcB
89Exsi1XvuG6p2oEgnMs4uaHmAGLFiWLhFAlso+AEK+e7Yv7RdMhlOB7c4kglWWW
CHhJVAPkt5BturLLNAJRta+ylkqk0yQrl4vVnipYp4zjftvX+LhcrbA6TnTqxPS4
OFAjTQWHqNCMhtQgsbiDwV1H/uXhey9ia2g0mqfaMctLPZGEcnwRbrb7vNi8cnDS
NY8XVxl7f22+zM+/WgEHuOb/YllX6Wq+ew5ipVgULvh+/B4o0FUsEFoGVseJIsmR
JyTfoPBjgbNDUDR8+pxhALrCdjeLD+IWvuAdNLwJw/IU6w6bd8BdBJUYee4IKdpG
iB7dNK+1fS8DdvcpRd+WACaoqNHdKWK0DJZnk0L6wafAsHgtoYhXV6p6knGrqGPv
ZtZdZkY9i/1paPxLgO3WMBQrHpGeZh73bry03b641yXd7+HCtkOx59lxi58ckW4V
DeoN4ZAx5Fb8DoSeVCSnZsEdxmMPbPbZ54w56DZG7kc6dMHsOtHd49ylUBnu/irR
bCgw1A9x15QW0EKBl7GoQhg55wk9a7CMB2RrOklSm4uHtfPc6zmH4QTwBnCzuVUX
je8Tc49ajKPH+MeoQ+TZLsE4ERNSkjIYoAR7fhSkTB3+v7enpqw0FhjFYlcWHTHk
KytUN5zfAxUyt3zZB9aiuHqoVxi22WDsIZhKpAT5zu/gLNLrdm4w3C5id2oyKgW4
A8TGKZdjAcm8/1jkOk4EzkiLGjBqPfdGM58WdL0zAf8+DQPZ6aM24/D4N9QRd43j
zWBSdidWNox370v6J2tg5RHU9lBxRytW3Skl5w8tckwBWmUgHZ/tgO2S2sQfBdQY
CqzafLtbDsPV5XFOho4i7nsP2TFem0gSpqM09ZhO2BekXk8Tka0z2TEcb95mMOrz
43E5qFt62TYrf4GoWwTI2xDC7dQmf556LfB0EgHVNKBbpXbaSUMUJJ6X8bSaXB8y
jWa9NywWhhWZdPtgzcW+iPkPX31z3P9d0OF5uYhNKdFNQoReTYlfYjhq02HBgK2i
c/91TpilfiB66BgKt0fcEWCHVu9H4ojhu0Wooys+tcQFUiFiCn3vObUEA10ahQ88
sy3OIYXP8E+bV5Oc/V8t/hlEfNHVaU8L+wu9wYkzcxVENIspaoNDaNKB3Xwvjro2
BV3liFxE/Z93PnrwJC+lc4EToxySLzTWUboD96neII+Zq8Ik3+Tc9GiyLx9BYvzY
dtjUsTZlbhQAcFWjY8dJdwbwii/YXHWqiod0C2AA8lDmAtb3Td2l5wqrKo5WTxtU
MeUbV1quAo+INO2AHG1yIh6zZsSb6bYD71ykbLBE5Zym42ch6PsQMyh1yuFygds4
PVFD+9mPntEUNJTlVRE69aq2tb5hHTQW6yTrIbMZqfhxW3Ggiw/j6+OsKWkLjymc
yJijqGGKBitOd2Cxo2VBgVbQupyWAQ6dPxbJ67hcLKEaQ6ItkVtSEhZcGNftF3LB
KAujTQjjbPa4gN5sKEkLsJmUbbT8PzX+SEEljYPftWPWXs8lc8Q+P1PpS7v7QPFk
`protect END_PROTECTED
