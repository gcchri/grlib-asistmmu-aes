`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fAnnTINNkR1APs6nbPE3gIwTajmt7iPpGOqnzOXDug53fTL0MUIS0TOvmERY0tdT
30gMIprnITdsphX6XmVOIHNV+srNecP9qeufqUgfkTTKgglkzzBY4jVjRRDsYthO
Rn0dnCPOvFR78iJK/iFK//hTP4y8ivoI6wjhSTFdNhCJouKHJ/JZTUftaY4v7zJW
kS9WRnMRv7YAwphyOSmXr2hI5oCBfzfw1N7KUOATKYxDQ4RX7yO+UmLSkA2XCzwY
vfhlPw/fdrNTov8dpRlX6lfpxs7KmZU6qaQiWxcxhmPcbhBM2ZeqLWG+JdNishwC
SNH5M/rmXVgQhp4X/fQF5cQo15plBOOWy97hKV8BX19uaF5xT6PdAv5FmMAPWXZe
g5ux4ocabPgiCqB1OAhlbU0fUr8UWvXxMzWQNHCqpB8u0bkWSyIUGeg3eBsSS4QC
YWhl0/xYIYVOq5Rqn6EeFg==
`protect END_PROTECTED
