`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cqKkcIshQfWRwMQTEsPJSLSZWlJ8aQOZSZhR/yg5Cf4ADbcdTtmi1BhDWt+B9wqZ
TOl2g3BVZ+lSNqtZ0GkEQMgemtrYL75tZjLiWvVNbC2MoJbc7OJ6S6rP2oD6/yyO
1VWphOSpQfra5bOVNAtrYeG4fEC3dCBIQtvTrZMs8QOd6SUbz4ybK8dKW+4r4Fh/
/0UbevqTbELbkTkTUFvs2BD+fM3NLWfVfoAe0gDC9SkFq4yv1tiWVRon059gRDi8
LB3t6EIhchbzYgqwNZ+F3g1e5VjrUa/G4kqcqiaO0n4=
`protect END_PROTECTED
