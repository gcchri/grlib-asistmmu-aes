`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BefH0yeh3i5RlEQzLXDknp0aDcqKbznajeZyZuef1XxVw+HPwe06ewTVX+/S7A68
cXnwsxhgCbrTon0NkHG1gbvC+m/3NJGz5tucQKyY5YJMUfWU/+/28w4e2Gc/zSaT
psH9SKSGtLsdgVqE5vfo6yXJRmxLVIr1/TSBkGj8ikevUA43lUxR0uN0E/hOc4bH
KeXSvUDYvJX1zWmG7B5o/YmC4msqI3pEI08MopSvDj7bKodnHogMaBEh8x/q9zIC
Ci4q1Uu73LqrE8UxWV7Eg5xuhF2Xc4vaoQcV0b5d4zrJS+8MCMz62MtSDthmxthy
az3RcRmjJdXQf5wMlPWpzAQpinX1G48orLWnHmrUQ39yi0UBOM9lcCl2xKbZyVwd
VD5vEzULOjuzOxZIczvtyjoxyRHCo7L9udFG9bO8JjbeyIbIyuq6FnwPjQxcWeEr
XkqeDNWY0aUfr+4dUXaeirLh4NRM/6RHuH1aLwEs1Y1e1Hpjb5PHvB7AnT4hKmUU
uYkBSy1SwpNTt/5YJnZkRG69PIkrePwwwf1cHfzUK1mOwEZM4xrh8Q/Ds3sQxq5I
vQBiun6Di4IiIpQLHr+3p4ZDlm7GdS1nKgg7VwpprXf7Jr8fmXPnXCkkbVgD5gqc
LWgkv7pwo2Q2INxlBvCiClpRKNPlUbDbKkhOAU5pfMMutSUq8fSiCrKRn5+XLqPm
O4akBY8QcXHsSQP/+RbTZVCcvMVKONGT9EjkOJlFJRU4iOONhC5zAws0KgHlN3d0
1cUHfQHDzmbwfYXvoTcCriSp87DUU9O2LihzfCAMFCHZnDptru6LEsWd6D3XjWIe
/Ke+A4q6hX7uloV+r4uxpOdm9BkSfuqn3sgME3n8QwiobhygVHM6PHl0YcJ91Mmr
WlDpM6F1dOWCaYo/4U/5XkXQASNOFLs/U9O/z5Fs+vPGe3h6EZM/BmPM9jGjEwzP
6R9gmHU/6LJv7a2lALGMPJWAJcXGXLHNJxm39Zl8m0lpQFRW18dx5aaCumvb6Ltr
MiDNxSRN4Wl7KezcOPLtonfGVRDrauFCaJOd2Vk4U68YbF1Ot/jJ9HSX3bswz/UU
T3cDXtViVsMouIEcCjegRraLYoJoVB8HfRWKZR6R8a/z+azpoCl5syyH/H3xSZ6H
cnvCsBH48Z3LJLcM03LJgWHzniw7V7vgLUS8uBVvJ5ZZcZ5/m0vzjPQn6VV0INIH
SydpKLAoctqVjd7R6Y2QOfsFdr42DWV0XKfNRQnz07hgxWwkklIhVrRxqCjPKI6c
vJggpiDL0ceK4UoSAb2Cyl1O/scVwQ72sO+KEmUnxDJWjR9Ycf/0A0RflHR2IBNS
T0JHTnZPzzE/ceI0H/UkeLqqOxHKNaZbD/mMjorK0NFwmV2yoRbLCbO4sN95fbz+
yV4DDfM7HEC4fdzLQ/W0SAazfPvbQYLFqvVtkLVUUW3QNfAygXEhC/urims90ToG
wu8fnDHJHtmpGwdAzGSaXwH774zDqclNdMkjUdOpxWaRV1UBQUpkGA/ua/66m0qZ
djV0nTpeWQCV9pgo1EMv3Rzu2jigiHJ+ZJ6vZ37KEcSDyNagMt4al3JeTGGOwLn8
noslaWb2bN1Br0icCQwVZlqqXEIt+PbR15bNxrehh/qzmFHFWZlV/yBV2tziqwdk
ji2wq1VY8UWWFAcEcKLkyPK5auVKg+i7Yoj3LXT86sTAXkeESBQpZwouTmNW5QsV
+89NMlLTpMxTQjh7/kf/od/7xBYLSACoKbpDkICj0AqpfgxkG5nveMSQlCpEBUDc
TL40ph+41pHRjsyZfE3uDyceo9zitXGoy1kRZrhVFlhIx+BzQsIlM/BwnWhKjMae
uEIStwHnbeFv9Xgr4HEfOXVCeAePVivlNsCYthAojCEz0gA5mrqvo9Xgyg4g6+a5
dvfc6IiIlsIjAueuXpTGStuOPGEeJ32ECtcePWZ7DQ7v7y94Iej8Y2L0oqhldohd
xdzRQvXsocs3ZRhC4nkSQjpAw1p91GMVM6znbDVnnnZVViqHDHRlDOk6ubDPE2qi
dIU4HBb5yWsQ7yrieyFzcGi08tlc/YGl7SdzQYXZgfA=
`protect END_PROTECTED
