`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4nn/qRYwv2EGhQLmgB2Lf3G5o0ktFhVd9uKw7dVB7tgSrlyVCulCM/yZveEHlX7s
FIBTNuvk/59zoX3Xr72x1yfBYKarq7nEnUQ3JYiDzw7Pt/AHZN7i0LHCvOGbFXyD
QJVTyFd7VyT+RbvZeNP5zp1M3XkZROqXVCfaSgi3pstBZOoQLkhC3RMXCLVTbdcD
Jv5408QHOpeeDvAiOduIoqfG4PaOghrjMsFDwoEKrSM2WBKQDHmfOndW8y6mFX/X
twJdMVgAE02vmopzUqJp3Xqkv95M9K1v6+yT2+XNCJorbVoz26FsPlfr7Wc9Sd94
nZWn4WnXeLuCu4cZiQNwIto+C5hJZBgExJuLk7kftQwDV6xu4/8VbFkx5O3q5KtU
cSpxDnkOF0VEC+xNafvxHA==
`protect END_PROTECTED
