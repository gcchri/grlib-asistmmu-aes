`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OFBAc5B+MgWEV/6+arB3CUQCkt/vE335iZgRN/3DBEOAPvVPvDm1gK2ggb3QSdEb
2qyyEDOMSHx2WepX8Ck4T+4itya4crullTdL7lTEVCjprJqR5wO6phDrvAysLCAv
OTR3yiNyu36m/QlDHwIk2CBnKaSn0OmiY+kZOqaBqkY9McmQ+2yq70fcp+nUDDWx
Pc4OnNrsMm+eyo5K9oITryS/CQc4MNj9ZOoCNY13S492l4sk3eGtoD6bOF0+IfRq
dcLmRBQDCU3Hz+j1g0CEjrNH0DqyIYC1B+ekbXOImJXK4k81XDCfsqeD55h4LYIA
UuljCLuUxljoTrVhywzS+OBO/FQfANuNIi4qrpTVsUeJBHHDdA5jFwBMPwj8ffVJ
0Urk4q3jRF4o7n06K1mv3bTDdBSU6pywGUscXG+e49c6Xoez4h+qEN0Kr9gzR+Bk
XG9QHXRXSis2ssgSS/XSfWdG+VLkpryDhn/S9YVvE9Xth2wZIXp8tn4ddpG4g7Kf
4CjIVoyCEv/M5nhloVuxw8g97u4wGLKqshYuLyfAi4VIcClnMNnkU6EuP5To0EpD
TSPl6NHvvbADC3Lywddfpz6m+7no/t1a8Ls5xFzkPsABCSLi6g1PoPOkoSKGRVcH
OymeER+Dg2C1UWCv1GPDpg==
`protect END_PROTECTED
