`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y+T1Vio9VmwnEc6obgIivl+kV2zjPFeIBTNrHhlz96gmt15A9+qpQUvAkeg+16QB
9qx24H7A4d0iy7VgXHbQdIAMPDej4rqYd/YFBlsDwRye3bYkhVFIaLfHmCvEO/Lw
WeOEUF+c0yy9VFilgbh+M4MABDOKIxB6OOrBELuHBlwTNhHJppnbBJcv43+Fh7ar
XGHX8g9tWovN7dpGadw1ac1rcM7BlkYDpr2KcVrC0Ky79logKoxW50ot75mByyjN
XbLeMZ1J3J3w95LKg6KSGMAT77YovTLgf9xqSUtuZfyRKzO4qY+n5VwdI2fgIYsJ
koVgWJ+EPzR8Au7a0QChh/tQ805twBjQPvHSwHYUFNaEYltUBhVqQ889x3q35/ac
5bM1ZCbAKcO0Z2MiV/Ri/6ooabTjnvyjlLg8BntYdwXEQM4RXzP4lsGXtKG4SKss
`protect END_PROTECTED
