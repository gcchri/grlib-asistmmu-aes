`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NbzJOxkdbRojIClNpB/izjnLjK737oZKjqInATt0gdM12EbZE6NiFAlMnCxAIIH2
XSdImgTrCnvfNR6VMtB5s1acL5v2h6XunpfSNYO4ZgG3BnfBQ3DjJVTuflf6vmBP
1GEjn5HbWMuYYfakA7j4PmlG4Ts/csLPaOny3dFo0HBhhurDG4TKJQkUZ4yKX3AD
hBIPeGY4eokL4tNgB6AUG8irHmwQ1GNUOvYGdm8hSYch3X+vQgvAqHWRxvT/X/Lr
Pshr6vcZl7WGSI7sXS/X58cGsH8syNwL+PfOi3E+uxKuj1arlueNPkb0g262XwVO
TQMEpIJA08TtpSjDZAY+0nK2+l2m5/yj60QijDV8n1e3txX6tuCddYump+dOaZqu
kejIq5CkUqtpLie7lBqFV7xqTlrw+2t7YZ8cefnAxxqU9TcepJGyVlShWglP0G5F
hiRo5Ocp4Zs+L8lP6OR7hXv9rLkXYuB11pRLJMtx6txmv9EQ6o5EpqI0FcEu9d/4
VhetIVbfnz2SP6MKC5SojhHwC+GkzQlOF3QjKYN58wOPdvvCKx7peVzCowsQK9T6
ULXDvhvPanw3hNnOJmd3KXE8Cub4RcN5hntH90Fo24FUjM6so8GArVW+xm0ptzAr
FtQsJfk1U62YYQefnBNtmU9CnLorA9cZLFrq+QCDxlBzaX9r9wcYXRy/tqpMKNGo
`protect END_PROTECTED
