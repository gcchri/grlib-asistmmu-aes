`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xdt0J5rEO2NV95k4yG8cCKcm+zYdTZsp0RW7lbwPAfr6OpdPfe9t2iUbQeODkqKF
Uizv10P4NWwgizv8ZRHE5x+Lgfnna+5wsmT0qp6nqyKFYmx2E+vUS2P9WZHUa2v8
zypAOEU8/RpnZFj2LRPECKobuULUPFM4SJtr1+NFgTb42Ere0KPaEDtIDs+sOU/W
6rDytvwlB/Uc3z049JvMzzRUn1WXzsMTuipNODXxzaVEZp5US/LehBS66DM6GDV/
BfrQ999y6TaWoRVv17uXVW/qRdueiR8qPGnxGjA5nCKsoTpYAlH6e5WeeROi7bpF
7UN6vYpNZQZ+RrDktudg8dR5dT01Yp7TAUnar+OvxBMr9YSls7uB299TZLY1pIzo
OzbPU4Q1mEB//YHUkJt99w==
`protect END_PROTECTED
