`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gAnETnElsGf5pVqchw33ckcCG+NKn+SWuZ9SBKyns2Y8gdavCjD0bVxhn6N1UXv3
KUEF37pDXOV7Rm6Z+Cef9iFjjFSwnV0F7IX947kDcN2hwvBM0HkXl1Q1HRvd268Y
rWJmy6k55LPHXz+v2aOmz5CzH+t/LhmV8iZDu7I19HZm+kd4V9ZB3AqL9y1Ka18R
FAeHFVmB0ItnMTxjtME8LhLTRZcdrbxYRc2a1hDU/dCdpMVmLU8pbl5DCdf9J6o3
3uuDnWsYvqbioTH8iOJqgJ/87JscIC0cqng31xOoNz49gT+zaB4uUH6niJ/0MsmM
q76bpr67z0qsYZgFV4cNjGhnrnt+o6lL9b+X2oyqLikefD4wo01FqY2bdthT6u1H
kVF2Hx33KqKQmIrOhE1NVEfCz+IxeEHCPR9/z9yhBv5XUT0yylxaOg4oFzV7nv4n
EMSeLRxMSwWCSr7jCqUm45E/SYlzDtDFCyUHQ2flliImq7yjlHifktOKASKmgJxr
`protect END_PROTECTED
