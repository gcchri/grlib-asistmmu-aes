`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sAZW6xGRDOOzghLT8T30O60FmnCL/l5+reDu8CdwFxWkoSCI61IU+Y5E4Py2R7VF
eyFbPTjtbzso3svrA3UpJ8yWz1G8xVhjjM9WHlU9g8n+RScdwtp+v0gS64ZiZbw+
2udCJBJqy58t+oQ4fqsbsMdXPA8BNaU8tJOrs03aOHxpmdYt3/9AxOcQGWbP8ffk
3vnPjwEhQCHbsOwZ4khEniaGR8By9GSEhYZsn+Z8VByXJVl55qkCb66PVobRuA2f
MZoLCXN5jUxmofpYMdvdRVbsuUyRE5AgETnf2rh/980EBEPOMeN1cR/jbyhbbwg9
1H9Lin5lOUYIaxxZ9iGVXw00nhvEzcnYnRkdUOrJdjDvm/EYW50OHKEVKHOcIVcb
7YDrbFYnnLyF+tZu9fGOMjk7aI/fi8ozxdCu2rPEcHfeVKcVQS2zx1xMFKFHrG4f
MMp3KljfSE2kY9JBxCKmxx9e6FCjUmfDuCxu85S8NWBO/k+xfjxaHJNQWgK6KyPe
HQJblipg87vNqV1b5VHs5wB/cr97XPagMK24CiSLGQbn2GRAKZNfMYeM9FWa2eYi
xJF0xo3hv1DHqhBM44Ah6ZtiVmUhWo9OsHhC8AmEmcnt0QQQw/JmGRa+YVwsHnla
KS6mtL2p2+SJ9O2wCBPZ8Is4wMg1Z6C1WqBYMXwZoW+LpcF6UecmQxtoZ0gP33yx
7lcTP4fc/LqT8HptcGj0N/XY3V+tRbksiJxBRM4Knk5hkWbHQ04E8/Sz80mmSbH2
v9wePe5HfdszVxZQ7igkRvefpNU/cpzhv3SljzWb7REIJcWw1h+fEos1m+G+Fpc0
FGuRTk2jSwY8LL8P6tXz9XayDy0zlLJ8RXr/NBWMLpUj9RJkQz6cKSXjXk3Ui913
S4YUyluOJZJJkTPdy8VWAzrI/GDCaq0lyFXHBi05nzd4h80R48ENDZtqyQt57eOl
lXtwwaV5Rf/B2cwjnEQzG1Rsp6p4txir80jXvuUnqDOCZFyk6PP2VZhMKjV7zo3+
2AvSYfbDnU7Zn6F09tkScWcQbKQw37DxpF8FOHwwlFsTjig6Cug+wfe6k0O+Bf6O
Gj4YnMBGRrbsJNKnQOzoqgGZDBUdv80wCI1FmC4bXFcnmRdKSPzm7l+/3xN463vb
ZCOCJAm1VAavsFQUmZQRiVymkVJt54mPO48XGBH9QjkOEOLG+TTB0T86+N2sKU0p
2Vb6gvJHumO38NUhEG22QyY+GzXETuBV2X8G4eit16lmxdKnJ3/t4JdG+KN+AoyH
2JhJJLzYxr02ifquJvL1td11ODpQSriuyUNHE+1vs1jE1Pd7WDIsiyRb27L+p4+r
xuejh1QZEd3wnNUj9mEOVLKZ2t2yTqCbg735Lo92RRJebbSwhew8AY3+oJMvoP6E
SihsmGGmrtI2a2hr94+cnh/m//Mx12Up6hTV/QpY4OO95Bh//HE4k8OprtzKPXcN
VtkeNupe99jj+KthaR+e/eYdG5yATEXd1O3/F5kriV1vGdhjQUDUfgzwq/X18kBb
d431vpyixwKXwVt1XjOWsg==
`protect END_PROTECTED
