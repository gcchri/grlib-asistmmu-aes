`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5rvr3FpqPdw4vqZvNegP8lhm8S5aosbRo1RkmmCmq2vBYSCmgeMCTIIV76uVDMM5
QpCUvI/W+Hil6+DHmh4P9WHmWf2fNNOm12cd/l9NlB2xG+hhBasigyTIMPzo3dqy
SP+jeiieEzYUDnJVy0MZBr7L9RHnvGf0N9j/r031XpZjErTPaYjQtNrk7L3yid5N
fB2ZLqZrNdiygnVDO75DO5AGcfphluGB/QmanaECjf8B5dJW9sgxrfsWbSJ8yCDc
Ihda9BXlcuA3txDLZy4n3u/kAP6p7rZwCjGwz58iU4Dt7CUgKFEoONh8dg64aDxU
S3OKiXf2Pu1MM81VIkR6Oh2RtoJyBYhMN8mVLhVZ9HU9ZZ7hzCkjuzbe63iop54D
rrAHiM17mvsoAtqSYowzZiDJYZ3ieDSobsvclextpTpc0LF8sUtDYY3xGQyuJpea
pEMO37PyDHPBBAbh9IvxlKJKvH2Rfx0ov/zRurH5N/+ngvdWLTjiEF7IOr6uOF0q
FD3QoALejBnrAK+PKgdzwHn4K76w2JPtrLYWDqn/3rT3UtBfTgZg/Z9+wWJhZSg5
MdLIUVde/bq17bvPxuD9coNvSyDfoloPBr8lX00Vwx1QpCR3TZJEWOwiTC75PPHU
DoXW8OjrIR5MxgnF//vPgwZmBjn9xNzj4/qkCRVDUOGPBi1TgWzOIGxddp6QnkfV
nat3+4/pQppYaPTNGiRLBcH0j4ckOeXB9/LPjHJFXSckl/seIyuUONxwF3q1ZPx/
wHu9SO/abCr1TrPwuVKo2qk2VCsv+CFlS0E9/NAmo4Z+b1hs4ZOBHz0E+2KMCKu7
0PH0ugJJqBfKhGjj+t6nULO0GKyHku207Lc8i771cJKGGkAiRXc0n3TJokpOzKYD
lSTVNJo9xILRrqDCYChJYzpUxo1aVbvKKxagbaVJfJsJ1klJCWiPOSyxninQYt/o
L+mQe9Hd2XHEm5pKeyzPIWKlfwSzEiqhZ7GxHo6VcagGkab9R9DRsS5X2XE0Fv2i
KdKyvsNxtQzEfxrKGqhwcNtHFW1DKCLLCywYO6zKf0wvaeuEpyM2SKx8JOapl2/w
POkFz/4pvYLQkUAErYbnjygCeM3GIJCah7afqMsUyRE0xl/HRKivI/sW726Md2v0
TNzIZ7RwR6134xLmityouS8r8KusOGoxwyJxqHeX1HXieydjmCeJxUElTIUYNv+J
g3c5bGdmtXmIJ8/FS0AFSIOpZMzakEzlKYGezzL0Uzf60Bt437TTx2Q/EboBXQlR
yiD2Zok5gfVZFnIjcSUfjN08DkpXmpREiIrC5oL6IH9A1uqA5yqd6Jgm3sN8CAo1
acEkNLDbho1g5FJUHqFw5zk4OGhMj+nVSuaimn13+2sf6I84g/lZjnbGta0vp/uY
um7NN1Oe3h8WZOMissLgOUEyoa9e1FwAHa4P8xrtefodVzcXrmHyOB0Nzoatdv6D
XKeXGP1Yid5EFyiQQuix5z8fPR+aL9MQMRkUuPXpZC9W9vTj44oFOwjD3l13ik66
`protect END_PROTECTED
