`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WWCB5NsFjqmwATjZ9tn5kuS5ovVStT3fWsLdaNO0wvaWRQMwgtkPNPTlr5mrQUMD
ITbQj/gSD306hZVqkzl1/wiLA0gLubhFGNu+jr/uDbZ0LjgAAP7NoXNuzYg9lUnM
vgQjY3H2GRqt7SDt/qcZwNuKcKPEGqPyQ1+LWDiKVAQEIxQmWt44rpZ8oAw/YpXF
OazBqBBpYr+FvfLaeLi+aC7rHN5GTVueouTIiA/JDMmqmQ9lnjAU5sZhypgaHu/R
dcxbXtX7siokQi+/EaTPrN3qb3vffh5Mih9hE91lXPYbd3L6cbBVn1Pi9jP8uK+q
BJIIEifduHROUInKc2bZJMQHFqpL4BMx77HfUKEr7NghpdVCX6AeJg6qK9z1LoWt
dYc/y8A1lTBXuE6p/alzcoxK4FPcwNl2Zee/tsjI2WpcXp+DYjZojU0+OB+5jD9C
yVFb28069W3ppousVGZj7gliLPDunPACnzK6OEbzt+ka9Jxm3ogA7NOVgyXRpxRM
mUU7O0rkHLmdE6gaAJA3cGnR9b+BMwJTPqhQZnpIVCooYM1rVdl2yUPLFRWFh6LK
Kwb81ENLu5Lnz0GG3FuHGXHJeqNYi4eDguevBg3jIyCT2ql3VQB4eXBGzGgIIMI5
9t/IUcwRYXR8tmlQfJEbEvHd2orXuLz6w32BtE5E1bo/oSVYaNn0f1e4cDbGv8pp
s8BIaQ5RXQCyunnOE8C/+i9YzlUT7cPgPG51e5VVa87tMpucMvYhMNZHFRBrZDpV
xQij2t/Dd5UwlZcYpe7+5WdWqkkjA3Bt08wL5KxZsqGRGkbbNHmo5n6D+lJTwcCw
0RnwtePf0CZXVeucikByyyjbUm3lq/dcTfsRQJUohjtgztxZFRzy0aGwTNw9ZebT
rwZTUjBOYAYLTc3Rf2Z+GrDOaHNbeYD/zK7bISUtfuwD22IEmTDxlu+PKrlbCwyH
a1O3vBjL1s2LlcNdnP/oCSLM9ZtBtA9Wm3HrWZ7YKzjro/m5VMcoJF36TRfJOwTm
9HZAeUEfb5CVk6jfE1GDbxxTKz01tj7HzNdKL0XuBU47M2VJOEKQpOZWJm14CjMd
TnaYCGEsEbvKcndIBHEmoQToSxo0tSWnB9ogWvDMj5r02D96dAKYKYsVmwgr7fIU
tMspcGSbSbTHU/B1YYFkOALnWhvVoWZ7+jd8WM7cqH3OwyYdaRaoscjkA3ClygnG
tDm1npBgLhMmLjN6wb5pGyUg91Gwneijjwi0VVhPKnMmrhS/7o8MY9EDqbsu1N1/
C4cdv3w6EueIBSXLqXwDsg2+obAyUs74I/qPbBKeRAwSW7xluLFe9Xoj6Uvw5YOS
i21IN4IM6UBo8GIffRWecuXquhqGHcwtf/lYiJbgKIzPcLpIFUpeE6cqacQYKmU3
7GoDFaZklYPldIrmKN1k86wv5kg5a55q7YvDUbPZ/IUcA6NI2zhXRaNiInWr4aeG
k8XJWpduJQqgFuqEXuUVknkHuXCHx+xrJR2m5sLikU2Grwz6ldnYaXbDzoKPttIR
e1Vohxgw4bwFpIuoM2krs3bGzqAF8geSrQWuWDEQbhyjeDhGxrZcsBtgmrbBPrO3
jTvYAILdHaOU969A3WUdk39qMnYR+vaGar0aiBhWVT/uBamfgzvTqxASkAVXkhV6
oy6AwV2JcmAfV1h4pA6gOSQcDAWDGTHnhhlb7Ggu6NVECF/awt5RcRcUv8awr7HR
rtX63vOTfLw3t2K+AO7kujJ4+R7iTIfZwt1rfZEnWjcys/fu4k83KSr/Hc5ZnKok
vj36JYIyXBm4xU3atbHKLrlNZN1AOWVDcw9IDtMJM8pAmUehOEqhr4m5dGi9lHPa
IJyB7fIx+p2lkXPP9M4mwO7h3069+wUeiqC5id1X4aerZEq6FUPc4Z65ihB4fOve
vXwX2XlTI28R8OZs3zuONC/GPI3PIBNSvcaVf2Fvu+JApLehn0V68BkXlvHkxG16
DMGbkC/xLiHabiuUcNLYZ27hhiE0jNGMuDCkPG0M4NyG3I+8lTO/0EP1/5YdKOgU
OP2mTpxyrE53OmWC6QNJ6BppLR1QHH1puIGARy0XNhAjZ7aNO8Y2G3atlOM5u+5h
iJ6l3fm6ybr2sO9hPgnDPmSQVFZmpoKKq/siQXIAruKHvpekjWN8nhQLgwOZfaKH
`protect END_PROTECTED
