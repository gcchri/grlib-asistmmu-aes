`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JpP9KkwlgVGzyvxM7gC5w7kHCGm8DaCLrLSHYWh2J0zpJNKce1UaXurcvMsEdIGo
rNqWSCJt8Iv7ezfTwVsm5NBwPIy3HQRbK8iOzzEzNGxFvLV7WvG5D7S5cYPQpFtG
jitfxzk+HxVCZUpB2bPvx7kcfhwYjrlAx4uGYAlAMj6TVLdfi6s1FhdSai5hm7nz
W6LzMPoqsXQkycOkoqoIgWwtscnrGsnf6T+hu48pOOG6me+GTEJVJYkSKOQsxh1y
MzOj2cUbNJfIqmjz91swZ/VwXwyTcz39+azUBiifOOfjDXKu7Aim7aPrQ/SzdnK+
QK/6P5ANra/6fq6o+211q+e2zDQUFrzl0KDOQv+w4MA2gaqrtPrDLdEPd/Lnb9Qd
F9IrZZA++baWxRaMr6gmoXy87YQ+AJAHIF4AjPGnxVU6OW96PWMs8L6Z9m8TjK1M
W6XWhyKqJijqN9MK0PlmuwKDC7A8Zu3GBPAOWPlHIjJk6qprqZv8MzMr49jlt7sT
TniC8XT6mu2SdcuuyL7+LXtO8M8w1ARm3Go8u9hOuIfrWae6lUlkq0s2sUnyvuys
fO3l/7cRkPQyDB8fAiSVBATe5Z8ORwp41RH12uHzYBIFqZyhXuLUHDJ5YA6yw2zO
/dq4no2tRSvwtzo0S4B4ZCD8cga3RxDgW7rTy3zhgDg/7GGo0/eFDxOElvw7Jcc4
nCqyZlLAP80o4jrQIipIgvZ50X5f3ZeIEtKpFh6W22c=
`protect END_PROTECTED
