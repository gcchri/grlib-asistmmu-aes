`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9202c0pWJplV5rz1mswPJPD5c/gyI/I/Enk2RAkwy8Lz5R6x83+S7QglRY9PwdnY
nzO3/fk+LWJn2O9PVPBeu07hjyWSibNmzbAtiH9ZQwBtR6sF1Ls5KRt1iS0EkxvW
NEK5Z07vzlkbtfVswjmc80p7v8aerpQ4z6/3t29yquwOdXK8pb/xtxVyv2cCOK9M
QHP25J4w5r7HdT8fZQUHqCZ77znQUvS2aG8OHRi4FGSksK13FttyqMsvLjxJHtyd
EvHA28aFGjhuuvrOqyETTQ==
`protect END_PROTECTED
