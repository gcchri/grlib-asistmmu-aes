`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6LzMCqluvOqNRm6BoerGH3MeHEF/VwmbIC7PHHD5jCDpa7l81JhTeiHV4uKxyZUM
7stFr3V2IiQ4E+dodTWWJVNbswu81DgwuV/dXguxMA7DElyc30Q1vFkhw51mezK1
NVjk4WKDf+t2WAR1Ua3OawOn42LwmRc5eeU7ShpOzsF50GSaCHHkzamHmyzDpKeM
3i01xarBaxNJAvMAlYI5ESiP8yw5vzbT6Ny8L/9G7Ii0Wl4kTnNZuPezv/f9iTKe
ynvIHdLFJU+HFVSI0pdczrQxulqhrFAUBjE2JQ8vo5WzXX2wnM5a1Q9Wbv+Dltpx
l/YZ3ysnfbRI9pkoHcGRnhUz81mfZRPhyIEJroKlWLBDsAqthvlDiwucnHFMG+hB
60BhbA9ZM7jcdDrVnKdpibwz4q0s+5dI5xyDlscA0M7zReEtMkqKmrTOX3WJg59c
xKupTG6Dy9VUwv0M+IA2do+hFv76RFy+NtlokCvhxIkMDCFkz8KIhVYKPpwjTs3Z
F/sg18lwHzjnf4DLH5Kol31Bkiq4BuvUEZxNtCH6htkc9IauEG8pWSO8UiN+U6Yo
/mqRtnpvyUxgtl8xGtXTbRou7X4vdxxp1AztmX59tukLx1i92XEx2DI0C0JEmVjD
V4ZxeTIF3MuBLTbkiXUYfEZqXZvk8GbajD34yjeIisKb33Tiq4r78q3EstKhX9lC
DgLnKdaKuBcniHCmhlyRYZagb+lVymQl/GvRiwlh8CIFKyUzgA5YHVvgvhBNqPYM
/s2ZiLJaUQJXS3BM2c36rJ2INBvML9tO04pH+yfuH7bKiVDRLR6P7oCc9ZpEP+DJ
0oXAXdegwIuZlCTL2teLiiFD+FDuocIrT6vUZobF44QB26xjVufe4uhdqw1pZ606
iGV1tqYPiCxcFKCNd/PqPSMu1h90u5m8zUH6WW0xn8pYVBc1t+dSVsjajWlRBEya
PSsVqZhz9NAJpt7VHFt/cTdKvUSLXKbbn6Ep48Nc3zJc2jLn1BYIAG06c+PEIJI2
0GBHL5enxlU/tndUonnamOXHM4quYOSJuu4l+deLhkJQQ2CEzzph7vB5EuwHkDni
vk4Z0T/HL3zr7oUTV/S0GL5aQCgWjtCfq0Zt2/wFsEhHQS2WknOtkzOc3NBS1zhG
GYxFLWYInB61wnjJ8KLZa+lWAgSWeMa22iVN2OKAeUHinRcXUBtt0dyNy3dJCpCC
7ecCG0kddpD6WmdYTcbPiS70QPASkOaMSipwKgOz/EB9dfHIMps14nKCInTA4iS2
Qi/bpNfoxXSWLalODCNrrfrPzhTeKO0gqT9wbN3+NWNJ+7xMSliw9FnIBnib0XZC
utMu4odSMo3GDg7VkRW/j9v1mG0St9XmntATdHsa+FlnRVoJeADvkvVA6k6hCvY6
Q64Is9BZf0LUCbw7jOaPBPyJTSfZjXBsKGmtXk8Fud+jxHSHHYAxo6Jk6xM195P0
tmLT98xrzouGaAJw1sUz3wlEoIZ1Vppnr4fgfDfgpjBjHaiUD6Y7WkA0G3WpM07d
ym5dQjYRnA2A66zrqUmZOmf0zp6fP9TDYog+u6oHBm/4EySa+8TEJes4bssQPvbC
XrV1+ww0tIwJyKP8UHPFvNmPbUr/CxaNPZym6E1YhnN9T9/ue0qsApdSaUKdXK8v
ToD2yStPEIwJ9jCSmAoVeOpJ8/Bx/bXVMHwfeMk4nLp0ULGrFSN/1mbWWEwB1Llq
DzS9syoLUSzbgIwxpFjVK2B8+MYKGr/nMVYxrJv1GApccaN0W9ENTnhI6oXP5/hu
sK0GfmYpZAa3XV+M5/Jcq/YQH8bnxGdvahlK8xz2zcm0dshsyhfzstkZY+pKN8xr
MDqh2iOLEHoqkR/yD7sS31OQJ/qza1u1wRHPtxppgG9unwZFF8I/lW9xJvFWdNlj
z7ZQagfTLwFG/iWJYftnZDg41ONlMe4RjajGpleUzYzoJT1hU60hUro8/t2jgzZ4
X0n73p3HOVt5v30Mm7DhzTX5ZCVHPTlHF+5epE2DfZfXAmcMOV8XB2mgdu5m8ECF
fmLMrRk6Ylld073t4pUCsFjrkVe2xb6bVd7a+dwURWt3ARaO0pbmkIMogOgLYhH7
BfYbaRq/PKfrbjv9Er3qYLzffsWCfoMjzetK/Y/NybjkPlA2boEjbHcHHInJ/qXW
ky/CnjTHm9nUDisOyybbPf9zYTilv4pRs47FGB52Wjx2vB9TNbk/OX2mCWseigUt
I/81cuO6oeTOWEkutVTUvRPRuPhFFrF+mo1nGsB6abVOagmfq2CHXkXNIK4pFjTK
GG6k2EA10UPubKL9Sb2kIzNmCsOC+TV279frkzMZOV/B+H5BCwqprKHTt3EcQrmh
PMjIbyHeJXxQzbykuUqE3tHKEJNQPWs1N9FHQtKN3ITGWABI7cGU5t3S2L3MkdXc
h9g+zZatqZJr/e7L4edtPkdEIA+k0N/nNCabK0N82QJFOSjgNP93jPT0k/a4CiQn
YLHVDBCg8A0a76feayQchk71gkweHxg90QmPJ37KTQkMl15/m2dHFTOfp5QTEdrz
1tE4ka+vxn7JwUcLFWpTMxCMgnO3PX6E4wv6rXjQ031mcFOZTnog+NFBCUAsu6RT
mnw73kOnl2SbzJQg3MbtUojyfTlLUV7Xh2QQIBSprwOoC3DdibzQuAa8EwcLHEun
63TX9fphMAcr9ywdECO45JOLfF1pDl8og47u12ydaeswLD6PJern19W1ntfTeBf+
jf/J0b4MKaqnTZulK/ggJ0uyPtIC8TjpmQl832fOQuwydGGceVShXhR+IqMXQyGc
GUavsLUTuJNCag5rSDSUof+qA0LrrfvYQQVlnSVYvGWNKd4R18IFryuTJbsSESKh
ZhHDyHuAzV6PxRwXUhBjSZc5x9lziVN4bXOIobxnodawlqrvyJpadF2lwgXQ+1OK
XT+m55axd1ZtiXa/US+cpDN+fL2FLAciI3MmMxbqfCgncZAzU7jsQV/azEE51MCL
dlDEhoaKSuo9VjCtLcLNo6CUFQemTd3wmrNfFv1rX5paTtbdhS+mlQWl7Grri2M3
mF2K1auW0Xc8lme+gujOx/E90o9n6BylhmvuNwz+P6zWoBklFW+pvc09fJPK4FVV
ObBmIYs5WTi4u3BxZcRUoMl+4KzvbdIQqggJcWxzgMCCKyeYVD1yL3DY+w1+Bvdi
XdHvFaOGEcszLeM/xIbY7Itxgvro0MKI524UJpU8Ny7wQyOIL2yH0vJksBiCJggU
WddKIIfipJ00DunG112GspHdGA++QWLmqde/7fjx58qd/Ovwi1W2NUqLmw2lZzXY
EZqov5AwafMSGBk0b1LQE1wyGDdj299Vaq6gi24Ve0V+tCwMZMyrAyK/1Y6mUaHC
nfJEXqs5MzkCzOnFv89hmW03Z3XUTMbZf3E0V5UGDaGNwJUW/o49sKmu85T2SDYL
3n2K5fbYmn1P1UWEeVApQBBzqupGLBhNHzg3PqidKqp0q+ilTyY/n5k2UIfg6JY5
GQ7D/fXjVwHzQfRzQbU7OZjmR1/WKvl+vwhRI2qZ68HaWITnV+0PGdr/aJ2Ni3eB
xk1LkUPfcaKSLrpedrOW91HxWD6QsfdEKJmUHWIaRRZ7JzlzCq9Xi4iafPiP5RDr
SrHAJ/FAfhKlK3QkztZZLU0H/7Be1jyiBtmgGGKOkxSAAiLcvwyMlnawum4jJWU8
pewdKm5voyIshI6KoCtHrDJlxctbMxrsnfw8wuXEhpOKI9SXfDSSie3hTcRbFJmm
+UfnZTgaW/iB9tYvUXIsDu5kmKaccKoRI3QvEyKNkNRHJ0osHeLdJyXHlIK6rmaf
7K+4zTksJehW7cLsdbv4EvpcP/IJWwMeIQ9DG3117XedY+3DxUisqw+ntE4QOOqz
xulL4hHsKaf8QpAoUeKXzaH76Xq9dNn2SYpi4g/Fhggbul8O4VChFjGA1NSDd9j3
YHnLhbzQZgIfkf3xAvsbX7bIMJh3TnR81wXBYu4wkXIE7/HbrPmrioLUD9BmXB3I
eSztzRQ+9c97HjybTTgINkjqzZcdBQJx7aMm3uEEs+9wiXwVo416z4ZUU+2TFBS7
3sRQV9bzlVw2VR6TAh8CleLWsc4tmjkxAjJJR6mr3MmzZmm00gcT+IubdgJnDA65
2JC5mqWkgCeFdTxX1SWrv1/VNZX7ga8ASx3ujQY9I9z0iVy7mRNouZmFlGKMMYhV
eonD8/O0IxUokAgWhCaBNzidZmuxk0E6M+KI3XHvfshGJr9ctW48BNrzlQjmYrgw
R7ClI1aSKAi8VRyWhd+lXyUgFA2RT+HQ1IkKwLMGXFajLj1Krh+ev8yPgunK1iY6
oTdwJc69W0SL+k7MSx0kHNwa7AgHFCwJ4wKJbDLYhbFuO1guZg4u8gb4zBr1bIla
pVPUxbFFP0929c8q/tKLL7kirmClVxCHBGzOdgRT5dTD43Gv/QIb9gFJ+MLGbKsh
etm3XcKj+3CiKacOcjiEbkv/gQDfUOOmsqoUKL1fN+hT0DcCUIYyh98XABUwa/lM
zkeMKhrbGM7LL8MxLlCva28JhH5Ze40pPe1PTXDWFky9gpsqRj1yT3mAHIOc9Mim
m2O7ioapoxsQ9v4z/e1W3SjSJF215wnMEzSqPKvcVR8aTV+uPm3S5/NVtNvM4NgQ
jNZ0g4Js6rJel60RuVDnblEKshFni+z6RCpP9QwSa5GtMOW6jRwllb+LmK62MgN5
6QELKua6hoGwPTjXyw6pE6txZYMHgzKYv2W3kloZpNNUiJDyWyrP1Ru6NYB09AL/
wPEhFOmeQ9+FvYckzHS74YHuR6s/iDJtVvg8BLDFeKsZx5rOGmlCYSDkbjyD+oGA
8LT+xkWrTiaJQQEOEj+xsbyDHkk/PxdDRXi1I2U+gIzBH6k+qHtPl4+tLx1XEfzD
OsUFykiZwiRmcpBU5HG4gfOvcLxUXi2yZteWY7j13ICDVTHeWFh+vQDqhCOQnB77
4x/3VP6SOUH4KytdAURbkoBE2oszf5T63q9Cyw6v/bk8yZTcI2LXHb0PqhUipEtR
bsO6DpENyAR4Kcc+PKMpG3UIdac2b/eiOoJdvWZtW7pDMV48R6Lm96h+YFfrzdpg
Ppse6T7ewFoGtPpfgblmKcgtpPvI72nKGA7srfVZ+Jyg0m/Vo/qtbU+0yt8RGP/3
rcsH5V8XCwNuqO+nNdbToPMcjURlBeXjboUduFeOsAj4EkmoA4rXJlaTEwqN4Qzs
H1D98OVhZKyNFoTzvQzCKBUbMb3Se6cSqgys524cx/kfV9C94rD5MiKvItAnpWqF
eA7lxKwtCyFYq7xFEb5FLz7Jxzuz3JgfrNy3sxI9qA5U9JCOk0v/4n5HTTJaNla6
4xggGpvzFPfeSa16nv6nxuTpfhOXQyBTkJeyypdxQeXBSTf20I6l0PjhYRwWD0Ow
DtsBflLTuqX7ic2fjhXkt1+vIBeuHQubkTeueN1iBZ+Qs6MMz4T/fbA8o6sPttrF
ghs0oxM7NqcKkfgei43+AlE0ehyV+9W1gbOGogq+01CSgpgfb/s90Azs1PpJlre6
gArmnSF+aVnf8wneGPqMRQDy/dRFF0nnS8S8hC1UStKYm7ifl/YubMpWNfbwisR1
DDg6WMfnaiEDPdetDJ35iB3I2ZjBuAbZhf0Oq76q7dbUY8OKG0PplVq9H2WZPK9Y
YMChHaiIq/YqYgmJ1ffuu4b7Mp9iJ4UExxg1Qdc0HnXITtnrt44i7g0249lumqUl
ONlvMamfTkgAlWtfqSK9ddgnrtrwzgyPCa5gqcSpnX+1j/aspw3anQci7zYO9/Tn
T6og0odkdCeIk67z54EW35nR4lj0Vd0Odw1Y9F6gYyXpkdaGaYQfUL3VeHBWqWjv
WEHuLOd+tH+Mp9eZT3dLeDmPxlNn/vJL47qQKL+q9/0df4gFIh5ggYH3315kr0py
nBHlL50qx+FelHAq82+9IZEl3kQB/Oi1alRUEFWpeS2dwVIEKJS7HNCTsLox04bW
Nxg5orc3mWMcfK2kBrTNPgCsh2aCeGVJ36hvxLGO6PGc96V15zfOH5agJtG6KYGW
FfRQBYuSbVx0ju+UKJLOiAx8TSRSYs6UiWnyAWxpUN80WTjOso87kjDc1V80Yy28
06dsp9uHW+2WQSj/a62NAe2mNfd0tmrOjnssA6EXNUUxPmxmVvzsn4+SP8BHcK5y
ci7g0BbPeBwTsfe79Y9FI2erBShhfc1+pYhMWNFp7+hYdlKFoo6ykdwYXEpOciGO
cLOrsLwAQB91K/EbHJwfFGkpJpuuFaliV08itX9ADZ9Bk4sHvGo0q9+Akh/vqpSL
vqiihiPGukAzRBYnCfcM8j5/coX/cAfqe7eKmijsHNLWoEwxtqLQob4BJg96KKq9
EPnevTYlp3IQpGfZmH46dFzecumJtCEzELUPAMbhpByDf0vwozAMdr1PqMMK2W+o
E0Kz53cxcJu553Xj9teFRwNGymOoYPRMh0pyEygkQt+AgJ+3u8nzZSJjip9KbOhJ
FSAcrGNgn6dlea4AEQ+12Kxovsl9hcjzDsEQdAeEpMNFZOZPt2BKm4avWhMo/hS5
SMFn1kUUKSmlmMV7bNczSUErZE93i6cpGFmuDMETva1Xe7hqPv/iFrhbKUwH86db
xxlZDnAY2ji6+kdx49E0aR8FchwjENHJssw9Ya9hcjYIKDkOXQktHIKKFQUCF8mz
DDnoKHfsR7JmAjQz+v2Jijac6f1RwwVrQiM17V8YNWbGXCH2U/ECrCQbRa0Vllu+
ZAHhmcY8xzBOAc042KNBZqxJrUUU1t5nU3EBlsgoAiiDHQzeWU7o/4o2AEH7izKi
sLYjCgAhyFae5uNdVH5s9MDX7RQQHM7GhrbFKYfOQ76NsjQzo7xBNCBGoH5/xcIf
wxcoKrVHxJzyjg/qVQB1/eMvjfV2epoxyXLdf992HFbMm2Wa6UVU/6uKIyy4oUBY
jsOBTF1F/w0VDbolF6J43rVIBUn32xylSAZ1Ayg/QZsw0lG5229HSVd1ekMZQRSp
lAAqMD1uoOXBJPvvR7xF3v9i7fqAhlzM7nXSpKPohuM76dEgYuwFHHUF1hrC679U
nW9yqMKkH2lGB3aYt41UOkymaU+mAiyb3fEVO7vSGDsRrVGQvIWr/mjdYYJh6K3f
+zqIR7+gQLZPpOggFggrMlOK932wDwvY8gJ7JyUr7/SkMyoc7/id0ZQ4SwRA92Lo
ZSUyrMt9A3q25jeqGhGbVRcDWWt04LdYcOKI2y2XvwDmuJxQAoEqZXfkMMiEi3nD
AVEDHPxARrcqPBuDX4mkreLE0aqSVuWdYAKDAvdB+uTnQP7TDzDiVCk5WujCERbf
MGuyyz0h9Zs7i96k7zFrTtFNCPbkQliDlQzN/fKjQE8iIPq5q2TCWLXy5/Z5Ed5D
HEPH9Nqsgq4LGi50TiRDbBTD0mXHlOYy4CsrhMToNv47idF4uF5fSR1polnoOOeV
Tlr+xWiXlsEr6j0m+sLl3TtFxdkUjWPAEfDQ/dFmL96UJ5d2AOGilBEnj0X1ELxG
Xza4IoCUA8k7yV2EHmQ2lE1RVbfWiolr9QAyWyClx39NZSsNrNrI7e9rt3aj5Ua6
Abb3045/+NAOSsLQ10kQo++I+55KSOWTYHESTZeH5CB2T9WIkub+fOXzNePAoYC0
VkLZSNWdDKUBL7TCi7Ez2JcDcn/Ea40jGMU1H18k6YJ5oWHPlClU2eeE76eFkx7O
mnBkmptYAGNXIMtTS6pPMtOVNskx8qJBb7Pvy62ePihWs4MCg5pKoZaECObwkSk6
FjiF1zvJeqgJvmdWRCSZ+npYHcv8qurEoGkMYS+VZM2GO4WR23Dhbv6PgTnAtdHd
l6fGmVjmAsmk6oCiyqOSW+4Q43bGmrqIv+zZxQcrUXGhh14MmdBrmdAtAgKbal4z
9nxEypZcc+rcmxGhKmMLHI2WEAF/otnjiQK0G355n/H1peH17e7OVQBYwZyuSN1y
TnER8h7xThLZZuLD1vDUIOPwW0bYVKYa6K3lwZgXtMMwqU3M7jKW9rR3uiQZvhp4
clp8EGhCUkqOY93wjwO8dqUuGfnD6mxcaOmf0tUWyucA5zsPM0iubvdH7/QBSn3q
PZhBbQtxWpx2TbqiEJHP2fhI/8nUbHhWTErRyFV0bIaGFNgxsyo162ORsMmC/eP1
dxyMgF0f9D2WuJPBaXU2HUlS6/KNiYrF3nvPLdsa/qgyICFrnIs1kMF0QsgeMBGZ
rLoe8EfMcwcy7NDP94N8xBypZQ5E+B8no+7/OZZybi/iaLpNo1vJr1R4ZX9j7mq5
kiYHFIat2hBgrZVK90qpy0eS/ZW/zn/ArP5EidbrPQlMWNAcesQ+/Bg37xRwza0l
lQBHmWxaO+nOmK7z9z0BFIKbLcr9jDa32sNJkLFWGowPe5OfTE2LvOD8Ih+aDWJm
2AY/jQ2dBNVG3PDVBe6y1rnSZls6dsEEJnXRObdnv6Btw1GEIU1ehYpTDwd1ffYD
Y0jz6udWvoqq9fAGIqsREioThocvLvoDaURIaQmPzrXE+LWaarwL4fFWSgAaNc56
9wRqGIhLJj9xk6O2aqYFjkLEJu9mI0dwjlc/FSaRjQE9Voh7IZERD3T2EmZA9wUJ
Jiur5cuTJlFQSW3iS6lTOtwNi5WGzfytOYLJIQhd3PTh8ftMltNjDSTKSxoz37zd
F6Hr0sZeTJapMKedAEu7pnI2al/O89DzOOaw4rBdE8GPeXjfqx+VfJJToH6YgRkU
BjAIRLmTvOj3YQXHnsNXIMR2zZkF/yOVM9Bl3iS/nrOwVuDT09zGRU2KP5FPikB6
N1i946bKXDTIMpEUcKAeo8Ap5I2hmp+CDn6aO9DX3C7hrVXTnnLcQE829Uz4Es1p
AxElnavlnQuJBrizirH9+qZgjGjVFmIx0EgH/CYMGOhDzdlZq1sbQYUdEVOsotQJ
n01dqJW+SXEPJAPiRPR4FcRwzab9IuU/PdPQEHECKL1rSClMRw/6nIOluO/nbL3D
e3tJIDmFXJ4seJlAJMH8KYb6Fdp9Hu1gSx0u4Uqdj5grgWZpBah2TPc+0JYH+q80
2fFSJW926uupgRVLOk5u+Qz3qUXyID9IUBAtluPlqdFgfnT6PTZY3iy+M7Mx1tRO
VDN7pwq8cXyFO6zS0uvCtgoE4NNCUuZrlEfbXxG3tpMdTCFK6MT2Tteh5k1Trv8H
Ewpr5GsqriuAyINlDXlH+8hpuyUgzs4OjzGGReddi2XRWEaMOQeT0UW2scYjMGkx
8pKXRCCJmlCv4J05u0bzvmAsrAXeID59L0oMidcAMqurBFELW7IJ2rqNRvTiTIg4
/5dnJIM3hS8xnKNGwH7C8XJT8DS5GXvrOHIX575iP/T5IUcQGlx0b8JVNWrbui4l
gNKrveGOemarjW0qZojM8/byi585ZqLb37/rpyGbTkQoA2sd5bxS4ScIs5bPMTIW
IjIdLnuzDJPtCcvmJ5qWisQJPU0A8tfRjB4vwa5Kbd9O7Ysz0+xiID6heTL4AsGb
fKsZY3LR3lPYlOoN27WJ3gBX9Q90lhUZMJPNM4nhomfetjY5yVhBv7w1qd1BH6T4
EIY9cCBreTl5BL93jJhzS//uTOveMk3NPUTiwZmOmyB1PnHGqozHPmC+y5AhyfxM
CQR2V215DTMoqgZcXSAQmPlFg/AP5pcgkE+2B3091yFZ3GzwW7jkYmsXix6mm+Fj
8wxOyJiH4f3OBoLhP/7eGEZ20RHNByEE12+mj4w52X4C00X50RMq26HInd+p+dWR
T3E3pWIMXeAT7kQxXp7aakJgiARcIohCQoB2wFaTr0yibMpViLeqhUxF8/RZz1cI
B1p4b6b+j8l/UuQyN5224EHXuSw7H9yHW3EhDzuvp7TlbCn/E240YqXU4t7b835I
XER2CD3j2XSyCGCchNZ6EhJzoBtrsixjcbfAQNfFRIRPWFc4ri+4rnXIVIs5WpEa
WzZZgLrU4p+pBqEJEDJNBxlx/nm3pppsNMBNyQl3CeqnmvSGNlxJUHfSShVZpuil
UmAQMNbxR4EGSH1mhir/oup5XoTZwztBp6V1/w2+8htg3ODkYMV2vTe8Rran4/Yj
OOgGg20p3ZaHsXnCTxUEuEazzPyO6t8Kjd7N51qfpp7CGqV/ZMaiZlLAwp+Qnn0+
dNNmaHhY7UvC31YAUFKWuqI1e6T4XjegT7cVEO5HkQigsjzjTHX6Sl+lbWjnmktk
AIa3i6Y8tzBkftVKN5/avFHXVBHhQVX9XfiXsR+vPYlGVt4b60ISzy/LCvTwufNI
yYB0058+erS4kR6uNizNa4xY+DEWslNcR0guAH6H7mJVlk2cKdWQjPr0hS2bCDWi
FKZ+pO5mE0ipP+JTzD5yDikEdzWpLdudBWHpyh0Pj3cDr1KrwhrcA9yNa00Bucb5
LiNtSSjEIgz0nqj2a3TWCZgZM9GObpew4Ptt3kCPXzbjm4n49S9G5mMRzHtjdnxc
ca0XIbjCtEWZEXSvfNUMuSlv7+/uxigZWFf/1rsfTJM+iw3bO0vPK69NsLDBWLGX
uBhlSKK451srlERW3MMXWyLgLIJfFJ6hNqpw6NEvhHJaamtgoEfAtTMwaRl30ylv
twkGt0UfatCuf6ZeEyRNbE+32RfLs+IZskgLqcyqloYh8pa74zVmLeJseGG0jAUa
rlVQdc0mWzNzh5h1oVrxo+sbpyoETFempHrlqkgevlu2ZTbYueyeXFwpF42vBSpb
MDAa1zZxk7WO6ZdAsfKWfY+h3PyMzFzt3TudY27dGc066YxYkQWSTSuf9IvLN47n
DnPc44VJbAxOqinIm1wTsxzN2z5pXHIHsLIMW4pKHWhCl4oY8BWSkdjx7KTXech+
KsM9zutzffQATnHpvvRcT4jfQf9k+By/BbAqniDfW0TA+9Reo/TagmnzUEIxX+a9
qk3C4xQEPcp5yJJIlwxXudL3l1teAJuvUrgtdk4YhXpBZIW5A3Pk1hpNtsPW30k6
YuVb5kRpyMKo1QHGjGOfM92tu89/Mi8gEBBePLwn/SzQdNJR8UO+aNltFH0Yx5T2
eQGiPvjMGowlLDUGUlhuDm0VNiX6xktQinqes8JnDc4+X8F26lP+K2iH08d5DpG7
uR+J+n66YYTpFCvb+n1UtZs3tElTEMF+f+tu3inLDoVrRPCnbsoqpkmy8STBePNR
5xlkfd1QL/rjvLPqlgzHurHASzUhkAdYgOjno4wa9zPIOtM4AYjK3092Sr0NLp6O
Tpgknexx6/tFz6dCEvSVRVqWy5BrmuiOpqquoS4+8bIu+7yJunLy+g1ZManCFDwD
ABR1MIBmvhTufshS/BW8HxlXXb3tzTakxf+Jf0ADv/ZMnWGOnuwjhzEIyqv1ewgv
0c51B1g/hsUC/YPTo757rKs2sO3zi7xTfBq6dCmV3xw8YX0dhKtsXuO+BnC1d1ce
TDBFSWY44ITr+h4EsQryEFa/7wUXmMZxXEnZqmnSbDA5/1SBewCmVd6kBE+cKK/x
9XDMslap/OZNaG17e9b4t8sAtWKadHzH8+6/d1hKy1tegLPUlHILJ3ZF3IGQQqPU
wSL+ywmwlIqoFQ/Ibe8yDl0juLnxBhSj+0rZgDpkZO4L8YGLu4euurtJHNcg24kJ
e++FX8CNEnkkVB5R8PG1YLXBg7NCvrLyBYDR4zkG8gnPdk7jcCzh48kI3OAbsbym
whmCi1PlTYZYDmeH21MZO3orFxLIf9ybNQH2xoiKgnLNDwF/zM7c9NuZFyxwnz9v
5uiuoD8/AUIj3i6RIIJExn4OnsUiFVTHyIaVeySh/qkLJN1/wsIwvdIW5Go4+dam
PWI7yOUiRwXSAuYVN9hKqjzTjP7yIZZIlmsSyZZJhtOrl7ROBW+iCE6+S2VbBEwG
qyylpJ2C2mcK3vUZxe1ZRpXEPyTILGd4hirVg+1uuuKaZR5kBFOTIw1twU8/tlAE
lbOA2LYXDJck5YQCpHeFmkOJ7CM0k4G1mYCZ5FIXtnwf5rl3YsuKTMwBZfsyNZ71
ImKS7x2xRj7Btzhji9OHzu3Ylz0klnU9tB0IgefRmJdFghuTZ83FfMq6ONptgRLL
HxKyKCyk+w9+ynmH6G8gnqh4X6kHjrA1Lxk6fRiUF867WFMU7Twu30tHF9FkflS6
NBJR1rpkyna/dHmG5GwAq6gg236TDDWQUIYchVatrbFdR+edXW6jqGpn8ns6rD8O
nXsqD3Ek7w/3Sm8I/0g2JXXj2NRkYh7h9MZF8iUrj1t9HOUtx0E9RWZfylJXHhse
LZk+OPvw3gPnFOlCvgpz5wa8lQmfkfC70aYsm3MlJtS4LtgPfOXabeIVq9jrjfRv
KJkYwn8y3f6+s2CWFnS6PTeiHjwiYV/EzWjpnW3NAAsbt3ytKREo4j0XDzR9pTNu
J7B74wJRO1oBvhI4UFFkHDKWbMcSpVk/bh5e7CRIUfZnOamNIqI8xhWPYO3zgywp
9EGIezuWtxyYylm8rrF7lvFOlGhB8f8hZrhOngJXCriHt7JgT1utQcbz3iF1FVJk
vLuEtgsWPX/DrADF4E3dQVh3G9D3HYoDwK37Y2EhNNu+dMc5nVae0eo+TC+PQPpN
vbeOhG+YlN2nRPBDLM25ZHLFWZsselZeKz8Co8/Tv8+FFTN2lZvGMjhEIXBK3Sb1
fWJalVN4lEP27Kbg4nC6qz8PG07xGnnwAXvQit8NoROdRYNSzC4xYuTwEviWku8I
ajVlsZJQFaZmAMTR3A/iBcTTdvBfwPfMot3m5GXHOCgFXVL1XpgsSdIxCFeF4O7F
Ws0p/dKiUGY7AvKpFnnowXlxkV4Lr0tpVPNNkQc//xPwls72F2kul93TsC92ifkQ
1Z8dOg7tbs/77a7g1o2G7OsnkSbhxZ78u8dF9+tQN5NodChpOh30CmOlTTzww2uY
ntDPiaFmoEWPlBYooUfJJCsXoRX4ueeqUq2w0XByPstrXro3EwM2l2HZBrl2Lxzj
SKbH/dBBzJssDQzKfYT3bUAHW7cR9zUAWuvX1z+wkbB+W1OjEdxApDgrNT+FsX8V
RE5vTAVobgMdmREH/sO+o3TnL8qhUrtXk3Q16B/L/ViJpqwt+g1OWDUke1BYu7Pk
IOfL9M7pW7bKsNBQF6nXxvudxor84PATZ6zlRf7h6lJkgaIdzumz5T7npV8i3WKN
6ow3BtnQztgZfPabj61Dh933+LhMFmFMUtjOZSdMVNW+nRQtbyn72oOCZyKjhSVq
AZW0D1uaR4N/KVfvBpwjCvw6MuXyD9Zi164fLppWVHkdYGdC4BNJzNF+xLihOmz9
WExvnM2X+aCwSv0MHdG/RE9ZlrZ/Nqb4wBk4LEAgrORfzyCyd4I7VKwyfnSlffrf
CJfPlh0C8bErXQ1kJPdYf1VNzkvGqEydkelyo3HBU4AHQclwKquttvqj+ll39UuZ
eQK4gg3Ge2U3LUSjfIkZDdS98MZ454H2H3Yavk9WXH9pCezb7pukYoEcxL2VSiir
otbcNKj28jfELZ53s3MdIo7w28BEugwKSDgGQ7kC5sU5C/41o28m3ACJq2OmwXH2
IzMZeHLlKfcB1R/6SG9RNhYz7NmowDFXMwaPQ+osPfpLCUfo13GpPeFvHFWwPTT0
YH5A1oKus2aabIhSoNUHm5Vvgiu8eYQINJVZKw49z2sETfO7ALtQOiQZw/Q8lf+W
+92oA+iFI5WRO30/zWqopgaO3DAYnboJIe46A8LUHkHZt4BMfeVLp9JRAnUzN2Fy
IFjajry3lZOY4272oONns5DB68CGTYrG9bwsa6leLSlF0BNgm0uO4RZVA8t9gmyF
cTlSskZRsBj/G7VkoCHbO9V7U/woboR2NztJBDTcrKtOaQWffRDPqSmGUH+LBIog
CAyWd+impJ9NM817iDArQsDcQQizJ9yP1tgmMAzerq13rxG6ohkEGd9HvNGm+Mj0
aRpXblgiqMai79Pmno+dBKYY13eFACoSIP3vmvZxJqiTEAlmVlFeJcgeDFtwigPh
BfsK56bvGAYeTxT17+Alr0GYwgtAChBdksur+SypBjGxk0wr/Khj7NJMHrdStdp0
2p7QKchF8EntpZrmQzmEQhLKJULWVDxLg4AiK9QqhPLpn1aX2ny+27u/N0L+uDLU
yJswHu2HDeQ5horvv/qW3LvoeJ7SxS4Szh9UHBggjNUL12jh116uSHsBY2jZqAot
3OZ7EuItHOyXCtwlJnaF0viQ0IHY6OkdGXsuEGMcAcnAhjdfZg9/LPNXx7xiY6fm
mQ5zpC0BacCvIfxiJDFL0c0dFfqYoo04ftTGYe7xFRudVWyQi7XUQYeO477QJmwo
Q42irG14nZ5KqTJwr7CMVgIXpg+gPZbHOks1Ch2LCBEBvwQnCH8ZqwvuuVoQotGE
snljqUr2RK+boT+HSAutpEfyOywrGuhRQAz61YT5O4N105j41RGyp/6xNMUzBzZz
AQhWmHQMc7sRcKjejbqeBcbtIt8ZTwoIF/27Fz2yZpQeGIlHHV7Il+y1b1ts7pg5
IQWsXvDtcdQjV1D+NSVUa4sgkvLxfF0L+cPXogxsq7SR3vrFbXjaY6Mq6oE5uJQn
SHF7ZMKFArP0AJgo5KlOe55JL9XjcCoXxtf+mTQ6TY65mhFGiLIleT/j3B9g0lZf
fA7TeWMhUIW0JO4fftTMSaa+qu4anoVdeyJ0JPzOAPskCVPrseHOydrYioqXsIzK
zubmdZqR5jjfz3uRUNMB4hDxOIZ+5d4bMdiHFMYIlI1XIW+vsRLVMOLedf6WzbOc
z++jnCo6YBkkEiEuO7yt8tkRrYCyewAUJ5JfthrUQMRrZZzTOikyByFSZj1dqvvG
XLWfizNbdJAIr12Gb0UX22n9KzZ+JV2jIrlmTmz30eDSMKMtV91NLUaRfhkuvAuz
hnHDv8KIwU78QCUGySxc8u3RCswm9Qj+7P5DAANXK+jqe+WBzc4s8aNxwNFIrXoU
EBKJ/7LWCp/4rSmGHjoPqSdHY6glUVN7jpsEusN7y9YIIr6SBAAXRfRDcrJP8o9B
mW7PLRyrcIzQxW9pSR1oVET20pEfCpPzI7IiSjt0M1t5KU09xMD0Wc0jS5wD9sPA
QAPD6SIWH2zQWZHQF84Vbac9JZQ6vVx2vyIfrwprKIFgE7sxnzes4d1AmUWjf2ci
nPDcg8h/1yhk6fwEjEzizaS4KPq6DJ3vaybOWgX/pw234q+FN4zACNdTKJbB2ACo
Ibz+k2vVkVqbs6YhB5dIo9MtviTdYXCnkNfHJ1FadaV++xLjBgNiLeix7z4UK6m5
wacEq6zYzCSXhKuyPgcpt4QkAoxS7sItJGykO+93RXIJFVAM9H+8Eaf879nG/GPz
I7+8BaAyV51udbQPxQvYbvWLzYc7NKHCnLBxlqvRJFnXK5JuO16yuDbPV8Rknz5e
q307WM0IKKOu7gLG8xoSuYk+7TZhxDYMTZXjokrbfee4Oo9C1JGMbvT0omFCKEki
+drCnAOJt1IIHI35WVLV10MBmk+yNmyJHikvGYzyC3eUuvgZ4YY1trAcsKJ3VfHn
8me0oJVskHtLSeCmT6kIcbeBuiGPCYc43O21oGBfARzwvBhDfhcXSsCrDTNJUG8v
EZaSrwWNf8hymO0vdt1sQpUsnSdtHm2umIYo3blC79hyAe/z2bxKF4CAZADZurC6
Akc3cQ5chkSjgTuLRS6UINHyuK0cOD+h4HZHsuzVtSOAutX74VdUHw6eCiOHI/NZ
TSMmjOBfVzQXZMN+gJX+jnhL6/wAQKIWAxo72gIi/pJBk9cApgVZIgJLrKYn4Fs0
xl0aSRiAlNLfRKl0TpktePfywlYoBJ3ua5QnH3Owl7S1P97qOKdW3aMdhm7veAVb
hDWcakMs+IpPRFVpl5/8tmmTZyfqwekJBkBioWgjsnYebqQwJf8nZ8bpptlk2+Wu
bUmvMZicby5xEcpR6AjbDXlJGuVeIg6zbbGKKvH7SAHgNI/xL+Mfk1t6Q+UWDFYo
dde+J2Idi+VBu/DNl+afz4H5s79Is27izsA0kuBiVP9wrv2AAMeOAwQSSAySg/29
gZljkhKyQcOe2OZWthWoshYULEN07mQIqtH6u72OWSf+P67Fg48ejjq/U2a2CAYP
MRfo/5KusRjczUUtM/MUnRTaBdI9IvejD6hwBwa0IQJDMAHrsvDM5usJ78VUsYog
VO0shgQq058/WmcN7MPE1BXLDHqdykV4Aa0eXSt56aHnfQFsWeoydvqasY6+tyRD
JF6EC+TrC0rHzcxDWE2pTaO4V/fFMWnt/DrQw32iRTbnJv93AztdhELOwxZhm/5X
igyR0OMRegEMnTEpMcyzlltGXKgTxsIi61hZVY+cGE76O5BzPvZ+m9LcRpL/OYLB
ZL9gXgmTk2cNFmxBNdk+/pQZ12vIBhHAwo1U7k50suPvsh0A3XYiGCprYSW8TEdN
RwMYprq/5kY3Uf0iN+3Q8NV/UhNP6zqI25Y7EYQgvLsAWFVhDty8flp1DTPVN3GH
0g6CdyFzyU26E2XcX9+qIsd2jQ7VK6emLhRjw8oCHy21AQZSM7rbXSIAIjRUDTR+
8qO4C4aW3w9s1NOKS469R5XpQhE1s/5i9+ow67DjSFYPKRYOFDC+dYbT0v7eXjMG
YEG2FLfnthw5ASDBOPdrbGlaGJDohFzwqwNKdT/K4nenHERONipzge0q/tmt15P9
sXa9CikH0ma+KzXNAf/wSB4NO5kZ62BFJahh92pQt1XGIn83r7orXmNmrVzJ7ajQ
3soqXScXz7ETIW0NjxgLQYSm/0BbhA6eCBCn6MZlAvTMjjC0a/f/eK4K1uCx1XFL
rof/dP+0nZ/0d/3d5A3c9HKLyp/oedxkNAVKxvS+DnJATydRIS/uGmFVbhUmO8ix
gD91KlThOuDEZUwx4Qr/sCRdwwhVJ3Zc/d9m43U1jHtrzhyXIxZMwSz7TyCqB2lU
E9c9gVhxBWzJSWPLO+TXdWk06VSMGqooxpE+tocDRP3dfJ7EnUv/biT86AwINiFI
IG2o/fWy2xCb58NU+OR9jtS6Hw6uMBYR3ZAw6/LxjlG3R2QH+yUIxy1/UXqd7Z7+
3967RwT66XilUNayvM7qjTzqgmUgJDRPhETsQYBuwuQIG8n7Jt6u+l8bzwmdjLsv
3RvPNsmUf0FB9R7U2lqcLyDA++2NEXjXrnXLPstSXIEvhOhVA/5vcPD8IVkbQXyU
/XjKl3O0ZPRwqZvCRXg2OEMS5G5V/cYVY9NsuGy1gX4eZM4/izezXLQJcZHCMvA7
DjZdAyeLoSf3DvGRl8GTGznHEIMKDEUsTbDiRSuPqSKEv/mXnftaL4UwCG0LM3A2
Z8anE/ZxoQQtjeBqkCC9JbanjdiFPzHd6iykfUh0P20t+ztkkSyF0m8k9eJRbnPf
UzK15WvvqSRrdmErbwlmkNbZOCM2flkyq4xJP1TafUSlDb5/3nlop1NqDFCkr2BW
oDZaaZS4QVO5eBFvKfWWDIj6unOHyoO7BXDURVaSpsGCGatAzMi01wImOe9ytnWO
rPM1cIGeXMjcCvzeL+wxOukD+4bjIR/F6L1cV1mFRtog/MxLP7ydXznbzHwuIc5P
IhqpkhN2oa/mWj5zsku0WiGizY+4iBBf5SCOyh7DuyYYBn3eMy06q0DfB2y7AFmO
9sOP2YkcwlhHsHtjo21EFIYkRIg0EW7nh/mEjPYU07C0tg2VVoM6BmCQKsqnjXIO
0C4ZI9aWf77lOuglUFJ8Ks1kBADLJDqvMsRs2I1PNk55dIwjNXznZHP/tjTO3Sgo
AOzlIZs+SestaXNbH6X16N/hJYr2pDRzMkospz3k6dq3pI73dUiVZoP1rBchzifZ
9C+ZBb3y+XkjhopNRVbRGk6/BnRPdFbYXXIKizYZ2M1g8WB/hkUXi9THE65cs2dB
yOleBArPcXxoyPrzeOpA5hz0Ux8GIQPo/9NzOBrEg8BYZu7xhuP3oe0qnTnuu55W
+egI0nosa0MO/RFnqNGVE4jVQizlDtca8oQyAbhLmQK1gyczgouAhCBA62kiQszC
s0DtFG5cyREr6Mnqat5tWwk7EpxTsM39h/4uWUe9qs1sOwKom96F1Rfqmx/p9Z/n
KLq4LlCvONXzTuSs0J0wvP0Z+D936uKH2djX/WP54Uv5pKJlFufQInbrL9hfhcxV
/iotqllcOPZWWV6sLgFZIicL7iM3HXJFvvQtO6o5v8IbOayy1LGcxUo2WhexRpoA
PeCdsvpnxUDqP06RTRHJr63TmQI+3Xt7hm974wcBV86eNe0UQ6sIDRIW01ZWo0Kb
2bNHo9zPpPee9Y9Jhzmu1r3Tw4nEHCy4kLqj7daJCCVolCOpNmlDjEk6ztrOv+Ff
zJj9EB6GruDygDZ1P4CkcqoqgBvGEVXFaG3Q8+zggs4ZP9hoyzRRz0X6tDPPjRqj
0q+qcQF4Y5O24ZxAw40Pv7HNkcTlMQeN5cHyX0AWIzKZ3CfqnQBs6saQ0nJSAuu9
gcht3Msuvlhjs5gmOkA9LOoD1tGp/3IkX65u3To234Kuj09Je4rScaYeds56l92S
DJWELS6RU8gNTuB27hGQsq4RdY/yJryOSAX2flTiifHClTpkrncyG/BYJQpXGKX3
tVW3gOCoEnRMNUrSzl+7vAl69TmXOWHAb+TUiI16yLc8kV5tVLAVIvw54fd9Wznl
RlvDt+ZF0FxIsBqXgUWRTdH0XJWBOAQUOuy/S12dmcR3a63Y+TQxzJgrW80CNn0x
PETyNVTRdtlLTMa1cm7geZsXHLRauRvSH5uKKLRJGuVt4IAnat9yBwEQXVH7QU/I
cnsi2tH1p+OCS4QwAVoJdFJxgbFuzl8U4AOLFPkMJ14ifSO4ztvIYD9u/9I0n/X/
cMigG4nwLt3QLzRPHKR2M9/RibNmd5nM/8joQ/Bp5xcKp+VVV5qBXWVlKTT1fJzj
w6h+6YAxpDoSSV8hUnor3awsProfyb3noHwXoab2GygzN2NjyW2qDwCKoCaUvT+w
uyi4+I9wBqUZnStazCnTXuthfdyD45FACUbCtnWQbOnUgdNKUPHmk9yf91w/dm0r
qes5N/f6y6L7AiDX8D/VzNOFxUJZa2BDiEi0xvxtQZvM4mptMhFd2cDWTtCOTy1L
ai654dTmsmtErPA7SMlC+GyjzO2TvEW0nz+LNgXe33EmrSBTNZw+OdS2UCQEYZR3
D5bN2pT0kH05nhImzf79BUw9+2frkTzH9sy9dFFl72Vyh2wCuU9pomSUmCqLeT8E
KHaerqCeGUIbhxQYV/vuJB8Q6VqRmX1oUT00J5UeTknSmXo3H1qwEujRVj/UuG82
sfCIAzW0/bNuFO72ameXXhrq8XsQQBDwBoIYZEGZAyfKWMdvaOrNzmDgtytW0Oit
xI5HBtIz/lHXmUaiBfYIsa+wMqbqSJaXTH58uHG10y+gcRQOaqX8DxZrSBgafwIC
nSz+xw9nVI/HmhBWwua0Uym0TD/d4/LP2adPbfCxC7UzRA7t6sTHsgwwKxpY2js6
8l2eUZwOUKH+VM5wjh8GA9xztAwaTPOO62eIuYEk7B650CbGXZId8m9eaXyATdQi
klPwmCLlswGzfhut5Mneb1hOAJ4dWGLaV5auf0wUdvv2sbeefFWHJTJd+fXNSN5T
BwRb3CrX8mRORwjUlt/TBDXtiWHA8mD8rPrUeK5HYsnOQUaSr9G2BfI6rcxG7RVr
Oeci3o7eGfZFqWH2oYSOev2hnA+xjVm+/hNrUs6GZYLJKyMMW70KJIhaBCr0L6kz
MpJM+9Nx57czV0wCwuiGDRxqfV0h2FL+D9fY4RK0zhUL7JOJx9nWGug29RjCHh3t
T1TULyuzUnXK/7ktoyx2qhk8QGvu6aUlJs2SpWRgUpHUzAwcTdQBJ4Jd4oSqLdvf
2kikzQ7/ssnvQJStYTOCYu/ANKvvGKfs1gYE06WOryZ5ew9cy+qnjan7kyhlv+we
OvGvEZ8YwgHCyFux0ZE9wWknl01BwQQjl/3AdvCWmw/FCoTYqqCWGbYS4lKW9IkR
hRLrdWQOS4Z1PDAJ9/Hi8EXt+jt7SmbWNocJ55Swji1Y0Vzr+lBSRw3LVULjaA4H
SbnuvGje3HRBQ5E0Tt43f1cIJ4d5MKhlpX3QKbWAfEiE1gzjMadBLHrqYb906vZR
cXSNkaEc3ob2FgbriaQP9ukpytMhF1hIzMnBYn303fmOOw9g8S6U2n5Mj4mjUU+7
6iEfS1JoM7oXrwOpPmaFEOx4prpre8Qx/DG5SYi3aw3XIhT4zO3mzRndkGyVjt8B
CQ/eLl7hwY30mH2ZVrfUIrNsZ2+64wxKYOlcMoULmlORwvvrmDZRNpxZl0Y2+bUZ
ye/Hm7GA8LL7UO3rXbAiO7D1/VlNX7GAzXmuJ+lcq6aNIhlkX09PgM4armQJiYvN
MM/Ye9/4eIIxEz8zF68h1Vu/X38xciuS+mN7qJP2Jy4divSdGKN+c/BLg1lwZan6
ZSRaTJztDjqz49hov2RWsAd7iUBQixIaQQrpBjO6vaSk/vgisHwgjsZEPqU7eppi
MPOOSBBddbqTe9m71PRCuOhMjHDaDDcz57h3TWuMtNhXSs8naGyeePtf4VLd8fMD
spVfCc5FZgo3VUgNqBWP4z6b2uRGqZEyV6ktRVEOfmMT3THiiXR94bRIqKmAmp/+
DW3RskXRVsQrSGFfjX1Ex/uUgFp0YLkwWxCCQ+Z2rZpilRzRBig/kI35MMl5RmZF
/y4vrktDelA0o+2ka+A2EMx0on0AHeNOUNFc7xFKuib3zhV9kseLInQKFZVoAxJP
oUyo+KHSSi5cFWya0OruLdYZmM2Zjr5DnkpRm6vsACnheKoOrLTrrGVdjOFU5S3w
KekUqHSIH78NOsYFEHhnTNaGevz/OER9PdznnIwojFaeTTTF0YmlYLQr70wFQ4v/
CGttwJrViaTHmurWZWfPNQmQ7Qy192cJySEv4coeRP5mxo+c+YhRuUJ3O3KkFE3t
Dcza/Z1Xp+fm3PwXbNOyY013mUaLrDxMMDXE/Vm5CYpHOIxWoJH35ouzzlE0zHNr
3NVuapK4h2ZhBE1r7b3r77+XvTmL9O04aD063QSrm/WBFCD7Lx4f84QGyddd7mq/
NC5vRSvMNEt7zmld9Mln0NdOGsbTlVh8HCBlPR4XE81scQupHGej65DjDsijihOU
q54pYC4VuKYhqTmRJdRrT49qt9YuqJn91/NyDpt0sdyIpwfkdOzr7MpB0oc2QQsZ
X218OVjxpxk3Q1C2PvFe4Qb2s8SGe0JBqM7mJfbKyUxXFFQUFdbPWDUQOUDF87zU
3hUF/J5tpvXmStxnUXCBX89Q+vHiGcpyrfcf7taAYeJ8N74Afv9isOfqoAkBexCd
YKGLrAHX2qu4b1C8mAAahjvbjlEwkMw5yodVCikYECMm/EyB4WiG7EjT7/Qn2yNY
7pFuK1lUsUPEo2MpfGDOpyyhSF85Pg3ZMbyF/K7WMcU6YzKgavlosOEoMhKhrRts
zIsOXiI4XXwePxRkTkLoQVwj7BiY4e8XPlaP/5wPcrwBbE23hkMHTg3bwiJhjfve
XnLC0XJUMH+/pT/uPFFubP+KDl7/E974P8JEirHe41/MDAc2cXoaBKfdu5mkNWA/
zVYxzyDi7MZr8kICXHIMnNh+8yTvB5GirEb2SzJ6CvnxRlJ4+STg5Xu2nlQlY6jy
NVGFIR7GTxZFHvBZ8RSkKznF9ZNVXpggCWGlgmfa5nRTKHtlG6TN98ffTR3oVIjN
0OycC2kQrfIu7Rh/TckQ9plwwJghQxrNmxfCQbhUYlGx7ZFJH9r3xwB/t0ie8kie
q0F7lw8Qm0O/eN1buGmf1TVhtTDAp5joZw70jVfQX1D3Qz8CA9ijJEMyIJhxrM/R
tzqk0s4nONlK1uB8VCHzPE1yvrqM1hAhHhzovWYceX6CI6ZiM1yYqmfrVag6EIwB
yF39XuT1y8pB3RJ365tzWkybD3znJ6zH/fFhO5fs2wzqhcHQATgI2CcTTMaKTG9M
1jygo28sYbPAF8nuMvQ4zwMm+TTN0iaxAI7F8YZSCvnMkAP5wkjQhoHqQ253tb12
7SElG/GMlLwgLH/G5xfwP5VUOsOHb0Y+RZ7GyZrr5qhWMQzGIDGkWKH6/EgWFGCQ
0aw87fZXwr0tzErpoeVbPvahEuSGnHATYg+S/ZkDJGtKnRDoqMG2lXFB8vNMzxT5
ifYBnFItAhITd4dCKrSTuh6mygkTCgzQkPpzGFO5QaSjggRF0aoBQiG6WHqS0h6C
AOnnVtkwadyLNwjvKNswReidW5gEex4x52MuWKy9eqjvjqHmxE5a/5XjVByRfenb
G9/vodj+p3FX1P7lrRNpSQCWIGzPa1MDgjxF0qkeTrAuvPFR5C5jkh9dQ0R+cUKA
a7baSOWDq36k2HAJKBrkytvA8EHOAbjlW/2oeBBk0M12bNcVOEVTWgu/FYxJyol3
RIBmBeXMJO27Jz0yJCCJsSsEFTcKpgP5xq9/9VgMDqsS97cy8oRDlvP0Rp8PB/0e
zQ/0PIzwYrImM/q6E1oJ9Ti1YMSgvFT12eVOx9uEoALF8xId7aFDG4tCa5fxdZpN
7fq5pwz8rbjqcDCWLgzRCyR9hE8Y1KPS6Abl0EASqNGAU86m9mgWUrz807zNAk1G
s+akIMyLRJBrHCQV2QfIQyJKkQFjx5rOew5BPD09uCePRbH9v9/dy4qfkm3SYD14
n1Zde5QxTyPFtH3W85v9MKVb+EcRkXjQfzf3Gg0kT7fHjYqjLZhfmNxYRjqxLuUW
UgO8nIsCn/qCq8v2Ir+VdF1yMi++TeYDJec822w3N0Gevih/tt2uQd+a3qi4qSgH
TxIGjhH1tD5VWJNlcnBpjTSDSCvfDv/r9+XiTTkgZp/oRJQBoo4rHCvOTW1R7NXi
adqMiF2NgIedP/JvYonEfVh9hQHayW2/82PDWsq6blWOsZIzQF1U9lIGJhttqsj0
kyYvfm7+wvvrHpAhS9xMGSHMQGRVbln42T54HMKzOFd6I2/g91ec2QvP/rJY/fjG
sk6zRfuUfXcu6uWpDKtl3ZepM2dkOnPnR1yYbgAgMjPzMBPGwzCTO1zwaMzFVs8x
I0eX9akANIuQsTucVYpA2akAdOG4uiC16sdAWUgU/ijqrtMSmcEofY/IG2kZMzhl
+DzduvIJl/PV2LSzhqpLhx6Mqk82i6YlfEadCl4IGHLnh2PQKqA3OdQ3Kr34pJiQ
LhCT1ChqfIs62h+nn2M7sVMhwk01pV5AjhtzfEM2eVWx3aHs25ugyclkVAAGog5u
NfLwtkKgX/UMTN08tnxtNQyvFf8Z6wgS3r3zF/9lvaYhUXlVq1sNAZ7SxO2RYXid
n03HMfTnUp7KmH0QmC2MeDAhpz3iW30QUYjD5g5eF7gAAJKZZD1DmSGNRuD1MmbE
eGnD9piwp5rNzdhSsOCmE6X3ytGp1OjyxHIvxROil+OX2atZ61h/HCuHR7qYUva5
eoF9/bsSK7jQw1oGrbRJSyHLm8B0FkP2RuIQZorC+yjl7JaJ7WZBBbilIbGYbCR5
Tmu6KJgVTxcxMY0kYVv3lWfqyWCt6UMu2CnuiyRCxrfzAc9nMSsxg/7o+kPRfkP+
8H0TY1US6YkbvsmPYSUYqjo3WNPAcnVRGXpPl6bp5wYCi4pdTPn2i+oqGpyBwV8+
YuKzEM+mBHCtOpQskXd/oqY9JSm2ZBtXYkN6PsLXhQQW+/uHlNtzAs4ZsCSca7SH
+5f8E8yrlNOKXFS1WNFcAImoM551ElhpyWOxaQoZUYvVYRkmbHbJvR0Yb5pshWGa
kBP+x3cKh5h9+eUM4Z3yL+W372zKLzxhKnhPxACdm+w4S6HC4m8BZRTXBkEORGxS
mFrRqRrFhOBFiGtF1tT8guZ9M7UWlxvGuZEaXM4YFLQsLSv9ypLnOUaqRVXignd8
6PM9gudjn1GxzBX6ewEx+Hx55N8vjDm+CkxrLm3kPgro1H03v7r3GCRRwDMWWYrq
W+JFHMzrko3oYwKS2SI3iQdZNun/V/VEk1CxPUdHwn6Ibm7pmwQ6RsWRY+aNjBpA
uu07Dlyzqjee1mRb3Iyq3XL7wEEXBsr41uLbhmtVal/csbirOI/ErPy0hN2mLwfi
9oqcreBYF6Sp4bvLJuvGeu8i+dEpwAf8Pdl+lmk+a7+UOFu0fDuYAN+Vs9ydZWhC
mS+V2TZshVoZ74xzuw5At/oWMJN0ybnAaf/ADLLtIyE3yJztPOyVuMHa33aukgwq
Banl51hmnGgPzQUKHRdl45amV1YpYfuAhCOhX5KWU/fq0lES7t/39o1/oU+fJKuY
nP455XN6iS3tSScuNocnEvq0kXLMTnr8+e4TGS6stpYrCPDCJZ6XmKcpD+Q5URBu
9MgKfumMIecNRzeSF3sr7Y099c6wqXVgUylJH7BlRqwhECLEL4VJNzjFKPVWSQuL
4CqMDgKPcZfvZ4LaAMLma5/6p9CVM7pxGItSfQuJHMjOrDmLc0mVj52QneuAtT3u
s+5rrwrSmgNb8X2tKgO26hLQDWq/iUEALm4lhCNGsG4rweQAVcD+Gs3JJqa2WGMG
yLlb1AqPBSxj7WeUqqDmOxILe85123gUOI7KsvfsIoV34PTFaUMJHJtNAnTTatLQ
ZBWHnxgREUaz4xydHLJe4A/yUpVVdQLlqtUlweSXBaY7dtsmw1bzak9jdDHs6jBp
wK9smzxaTIYt/Y5dGkWEbAaNxmB3HlSd3hgshgbU9a4wTu14TtXi3fP0YPNDv4ro
ypMHYCuPKgu6a6frJluUmX7joHTPc+wPET3lLT1+YZSyN9mDbMmhmPcEXAemYIK8
WI2Vg2XLKNku01UmxrixBo6j28/QFRcqdii8lHC60uNKDJLn2EwZ5Wuo/C8HMwpZ
rmiCCsNkvkSZ6Vq4EgLzhlGcIDOWKLt2HOwaPajWZDawguJ0nnUfznJpRMXL/0FB
cQY1hbXAI1IFtuhXjEzPTTOUCy+tkoJMIkFF7lIgoeYakrVcpXZKa3EtVhG5wcet
jENuuxg2vDK49tITSffvjjgMqOZKynARGNSNgvXOX0dRpUEzEcH3vc36ZJs1SuP9
4BgcGeOzyGjiuoGIHztGAMTu1Cdc3r+i1WCC/7nQEieAHtZauzkBh01H/bLY5KsC
LEuN5vQVqD111tx/CXJk+IZiEhfqUj48a7RK0HuZOFFrzDDjdxIZhDkTxP8zYetP
3oyKFfDeJVQhyfBUy8tuToexT8FY3yepmp0vDnBiEM2tGKYhAxZGWy2OAgCA5ndJ
Yc8M+l19h/6CpxhOybY7i3DpPef9QXg7BODwDmU44L4+VBeftLUZ78tFIMMPdu6V
R1duXoBNx9w6g1zwq/sivXnnIuV0edWtjYu6PIiOvH15YtjjqbTvWdRfxaGtrhkV
NjLDqYzJUEIwYt77WNnFmh344qly5xKL8JlR5W6M6Eb+Wd1sYhoqBpH+MgMMpGwN
TZWCFtMpz6wdUY9ZN/1FTI5n2m9Fa/ytYcK2urNjDm4lKvUVbsNqG0Y5tNls4tD8
IOXiofHOxVTbHIWDvSr1q4Tx8Zy9UuAnBaVBrwIOPz9WQXBmMbBDaQvK0Rz57ema
SYjzcIxxbgIHynTs0MsOrzjnzPWeN9w/LOTZjdQ1uYVjauOrk4l4Cfdjho6O25n8
mOp1eEtnxNxSg3onCUadCry+PzxQH8hzqrY6sJ7OTrbLVjILUtQCnSJKSUUZMNvg
ajzFmJFIN6UkWeQsZLIdPt7DedopnM/eemtSAJRjSGeTPdnnhI75fd/c/W+uODAn
/gVc++dCvsYc4pTrk5fbi/BWnkcUlBycTmgVIYSMF5+lgrdlU+Iwy7xPYmGXmbV3
u+7PfaY0yTEGxF8igH2ptH07cY5fXGEg/tPKHnkJaCcHAk7uSJk9Jgp20rqrJmOF
wvJ67KMtu11nIpSgzPEc4UBdI++bYdJBUG0O5NUelk6PDcXbC84sHuG6ubQEhlQo
k69sAUqfnueUGxlWzz9cFYqAzczDBKm/Rnb20mVgsqqq+hwr8CfCfM3BpMy31/Ef
Anf4ImWJN1acEjve60pE9vVO3W1msCmVU+R2eMAPDiMnpfQCAD13deg3oPUtHyAg
7sKxBpbF8xAuLOCLY96ORFR7UtZCPqfcS2YD17QW0bt3FiDzhFx9KceEoUkM6fkP
jmMtMlg1+U5iwm3J0AiuXSJe1+3ikKKD0racaIfQ0c6AYbzX3X6hqexs5/NuTjTd
lBw26Ym0hR83T2AYHghrEPLAiS3Sfb+jrmViBIs7uybcZ2gI+4cDcUQIBfrwu0mt
Kv3iIbuvkKUpyw23WFdT+wIqBe8ZTr28u4SjnL5mLJu6FOoQ9+wdXBgP9ZWQTT5M
KQpwaCVfiL5RXHuSmyEU7ppqgS4MiWSt8QsyW19XRgifSswfQwZjVBYzSgUjgX28
ja3Y2APwloeISqQi7nin1tBV+iVqXV6ABS3BfLkAOKCO19EZ0AUYJFICSz1p7QvN
z+IJrxguhGjqZPwoHT6Fgd3dXZ6bQCDV3ieYCUVmKcSDHRX0a1zD2NXDYoC77fcx
3pH1OgA20ggyzvPU7dYH/o5/+WYxmE149XbxWIzf8bL6Kg7cYG1eLURRV8o18jRu
PYVyLfBtW4trXFQnNfHxaGaS3bX5iWdqziu8fuI1JVpDOBLcJcjr7o0PCMcxxZnP
Gdsneu+pFi6G86TwowdOXdVN5bvN55VCTfyHY5cOlzF17JCX/x+V+XqASbbQ+q0N
Wxx0+XCJii1MBpr38aG7RvKYpJTqFhHqsnzWl+2fEcmuE3T/KIa/k50IwfImcjzl
qr6naZH43laIQDy9H+hjj2oarCEdAOQQ1TZd7SkOmUUQIXDuklBI8V2y0RGc74zT
erwxqiEbFZt9WkPtW0/X2z5+Pd5iB9JfHKIlFJiDo2K6883I57xwJkluyZ5Zvbl8
LrSYUmrs8R+x9KbluE9MVV5y/vWFAMZrbVnUJt15OJ9SHC9yr/qN65PdeHn5TLYu
FEyW3KAykyfalBWBh4S1omIFpuQFShhaQvMHH7JCxeLkXmXgi6PADX6xI2jdq3dF
mFACn3kF8u8k6e8pQdvszneZlWkBVm1G+tuLwjjy0AWGgzopHV1D00f3nfXkrZiL
ppENBWoFXs6BOTNF41NnZWRAuSVp7C1tfhfT+awEjX4tZ5WUQ7qwi+LP4a5RHd3o
zGIlVdIc+vZuzwVzv4GmtFgSd4IaOD/eAjLk+06RkwcslpynKTCHhPdRLC4feM/B
tZ4InHVQX0giEc3uPfkEQvkQUyuLZVnFi6bHvP3mHjUp7cHeDCfPOQLvLuWokuQ0
JSgLPt1WBk5QuH9vWusmrq9nsaMGjdWHt6kE75SWw8BuxEGAd+k1W7cErVWLC4sC
KL9HoG0y9JTZFfFtJRoX/KCFLbMAjq0bOgFfjW8L8Hk/h+cLr4NbHQn/3g5O3oho
fLZoj/IX9h7DQTmQgVeZ3IpnmBffCc8JpJB3REZGn7sUGVsmz0vZKzY4GxivrtJY
wT7GDtpBIqkL0kVf8xIBtoBwg56b/vpdWW9X8kVVQIH/ccz2U/KGzPbc8UrtGtlH
6ZJ9i6L/hDiE5TF0CGedVHovOzVwLo9ZtoobnGekjl/DWzsK79smF9R/Tp+HPf+d
wOyqSNwVTeRIk594HtCcenVVbhOVTNKZxGSnvgVbZvy9cVL53o6/lidq9VB7kebK
1AlV9q4hqZHQDu5wpjKi2Ax1xByE6Vmva+vjoQq1WRZOdTITwQqouLeKBqvJuyzd
POhIzbDZu762bD7ghEsyTFVVBJTppcuyM5Qau83egBGi9+sbGQYj67rtGavE77ak
2jee3zWdIkzQdqXoOtZXUwHjTpkbAOVBu7hcCB7epXQi/0gz4k4aoq8+smX9Ro2y
cik804K6mF2UoDCyJT/nQ1f1YZ3bq0xFfJEZP/JBmvCOM/0NGaqVxedUeM3vm522
BLq0q10zcoMyzbyMSyHwuk+CGDvzmzqmUHhXt7n1QkAGNpbst06IBaWtVanpIK+b
Szo8aKyQYZ6RlBSj1hBnpc9ffLC0IUbZ0b9atc7f2yrTUGWZjFmdGYd3BlQPLyFS
CZhC4xyFK+N/MApupibrAakGzjT5UM9P192vkIg7ahRZti7VNYabmy6MAT/9Q1yR
+JPIA9tGoMDuQcmfHeNM0Qb2QuJRQTnhwVQ+yBeFuyP+sWMdmNyKsvA6VktpfAsd
Q+G1ELvMExFI6Al+Qs7UxPotRCUTDhFxpZ/1zrwpLctjSfUfZXipyIlYPSj7JC7L
PzsJ5u7sqIeE+4X/zplCD5EAgS/k8HOmLSPvBddjQxCwvwLM+SbbiL2Qgp6ocnJn
j/VLeGlIjCEHYFwL+mdZVV6J2u4d5EqR2XMB2uDrKp2Ae42UGdFNArT4F6Aej8R4
bplEbxFcy5Aih8Scjf7mZyvJJlrj1P8ZAcD5ye17ylWZ4VX1niQ1Xhx7gMbEy+7x
+HnnJ/OUau9+VaTWny+jiVjg6krYv9YKCvi9TKgmzhwYCvDZ4jTJv8FlfgX8tvEE
PFVx81/MiXtWMgPaZ9HrjxVfSCfmPUcdWbLtzwHHDbfpkXG1q3XZPr4MtXGFw3M8
uus15TlEfXikaYOAB5CiPKVzraamDlJmaaXzNaQvKARVn0SRZBM6ViiGOzJF7hL/
v9QNPJ9j3uMPxo4pUFHnj+zqZITsnC1a7cnwBUq0em1DupVFqGs5TXRnWh62qBGK
FfKBHcga66q7p7WW1vMJH+MH+xpvNzs8fuxSCI4frN1CfrulmF33M1ggoIkw2XRM
rlGldCHTdvfTD15XDVVInulTLBITbh/Cwxxmc6nd92RY0JMvNN7FYv98Ow7lz9Bf
J18O2O24L6IMTalfXsrbnzGFH3Lg4+lPhXt0M2IHToFrf0SjMJObAyjP5r9VSeEd
447CzlMeI40bcL9ETPyC0d2kTP44HAh5sv86yD/KpjowUD4Dr2szGzlHu4Ispu7w
Rcx2yTJWNaVtEsI1a4RgzGzJJYwK2GofaZZtnC3PsMIS+aXqBcOZm++Bxj9EysO8
b65hqE8N5GQYYbJNB0IdJNj7SLT5PHcR/FgFWOCRgWJLvuVlhP1Pue66EJ7G6ar1
ZaVY+JEZVvblgoyL7Hr67AvLPGBhwJdPIUl9RAzbLScJVgLMYBwEvVfc4K5QV76n
66Xfz6IVYkhQi3hR/2OYnGhObqqPcr8PPxCQnOaKWukbFbxK7OovaDfdzCQJklai
7ekPd4TeQesBYStSyIaVyTgYX8DbAYXtWUmQLP95kvzVKaCgz+JwQP+GFGHTo0j8
ZbBuAybzcjIpinIwChfx2QujkVW+mnz46GxpBWP3+52Jx3lEzJPOYa9bKps5kI/+
qzNUadVdNun4mnRV7meXV1P1/ZZvgMuBE2GdOtcyjU+PJcAA91AZimhgKFR+VEOw
tUTqcQ0EFaZdxYji/8nstnyCOqLlD9zK5YBjfn3oFE2fTzM2iJKJUH0lH6PWkevR
g/7uaT6s5nwlk7vvD1CbbeSwofL2HjQS48+E0VaoKK1IaHTYfjLX8qHAstawbLKX
1rpVNylUn8bkxTjUQofoEnS7srMfRhDisbgLmrdTrJSLWdoUvY59grCh3FpjL1HL
O1Ah3bZkJseMb7ABLvVtfKBSMwkXhPqH/vXkuw2QF2fYgrJvtnLSixK/kUtiOF1a
7qZo57wzdbCp/SKRZFKEFHTzGsFnk4IBR6ip3ByezRdKDmHgc6GkrrpK85nip1KA
0MDABSDcKyD8KJruwht5Uo1B7iyO3mhtFYLo2uH0+LhXA+FP0AEsCZXNM4i2Q/MG
FG6NspeCBxETXxj6P5x+fmEefDYW4LePlht1scVHFEFwLj/X+zkJLedEdPofirIt
htIeHxLX0oUeu8is2zaCcDQ+Z5lhcwyn3iasoihGhq0OkNVl1QVywoKC+mcRRVXX
TOFi1sJ4LxAxAOMpKyHL+3lBIU6jRGA29FvnGVka2/HiFCYmuUireoCm9nmcFUqb
7MevJqsQg+AI0sWSNg7e3vUoxuZnI8n4KokKS9GX7y5CBljO4UjJUba7G6yUYGh7
VW0edLqQnaf2rmQQpCL0+62pqja8UccbTBFRcKl0SecfJz9/ZHFyhyuMlB+PZI85
OaCqCHod4GlQQziRYWXQDKoa0Ua6TMXiqp7oHE0AzFGuBeSrhKCCBdD3/HI4nbpP
xPeWnIlrlEqwfQ7PExpRpGHi73qqYXSl9TsD36AZ/E5h3z+S/1M5janKzLDRYXSq
TVth3OLqTlbobTNwUzknoHeXwqevjuHPYYaNwksdIWiYX8Sg1MlFMxE2e5ZQNrTn
BQ1m12pVtffa921hLebFy4mt+LSweE3LIwAQRKItu8wNM0R+vJUPPdTUgiaFsG+4
CEoWiL5xvvJGoTm4nO5pJgii7cipvKWOBBKKYXTt2E3zhg8QmVYhrg4aDF8lErJZ
ukRNET+634b/wINwL4sDpOJ3deLTvggebqkGfwlUL0XjEt46ZGmLZWhpcUwHa1Up
3ZRM/bncxRD9QHJbbtAUf65bQ8S/rkEsIW2BuLnu74LR25qS7OVwOwsY0HuCw4UU
JPeulgHMKWpjNeR9NWXypaScppbURPp6BWGWnvL5dZjCk9l5iCqFNG4SzCi8xwmE
toSv8LpsdpJnw0avt4OOzmDH0Umt1Ar9XVTMXUXKxXZaXPGSlfFH0y4YsZZRVIeY
0VO1nJxs+MUnb3YpebHNf4X16BBgOoL/1cE/SWcAoKjyNAkj0/kgHiSBNaenr7Rr
uZOXJXG5v6wimM+Mo/CcXAnU2HEt5TdmKRj1lJkss5AXByjOkstQll4LGaC90vB+
qvL7UqbKeYbRIGZdbcp+UAab2ZT7CDHOfAlE01DQil0x0aBumtkx19h8k8Hns+OU
v3Spzpi5o1HsAYNJmN0NvETYvL582wBPc99cFxEFPkeKzP1KpsrC9b8SXGynVojB
+UwjSzFKnP/DxhTW4SlmXZpyrbC/8CkiMCYBgXGKjZPpr7jo4RghV9GDjGpla/Np
ry0HpNxBKlb/Czlkr3pAKKWExdKHgq99X9V+olcBx6jfVFkEfthtydGB6Vx3JOWu
m8Tj6JO/0q3+6l1b0GPbcfx/GvVz5UQvhytAh895YgH9tcT61+GCuPmtgx4hndV3
JPOuhoKXSrxdBYBKv7GE8Z5k0X3wXTaRUTVI0SdhMqI1OdLNRGNMMT1FAH3lI4TS
xtFKx984VxUNA8rjc2AzXVmnT/OhhGAeZg2w0N2yHW9Y4lJGyE5Bi67yjDUKPgHo
gTGkpf0fS72+llJSBYcGh9ArpLDNWjRtdagzabTJs0UDIT8g3DkVwZdIa7p4S5R3
ok6ZDK8RnvNX+QttFvG08paYPxmMWJJV8AHM5bKf3U7BTRaQB4Sj5IHdrd3OC3P4
dqsQFMkIlnIpsxDyqfi5ZpsMr9DIunNNqHFvKvkoUYXom7i6hNorpA4vCFmh0/rV
vwolsA+frzq3rus/4der9KGa2n2PPCGePtcVTxPwHn88R+ImLy3JuPo3uw0RrMBj
Wow0lUgiJhGlwfbvIgfh6U7JlpDxhFrfhlCVIbTia4ExVL0BpOYkmM8rjnNGN+nm
3BkFy9Zt6xqcDCkE1uC99ApZBEmo3jX8GYcBNx/Es4Zn0VwHrE8OVcQDVHR8wIeL
ARmKdYMJW1HBy6EsH8P48XsEB3Mjo2do+mvzkgYSr5dSRgjfwfKFMGPZBHs8H6qQ
772IjOHEcaCv4TcZW1TeCCIDNpPiXs5sd+YidPsaSwL3eAbNqUMAqCU7QlSQORVP
lTRd/LkQy2MqSLIDfbewcxuv47tRFbf8Ut9A8T+fP6qw6upY4IFP8uNWZ8vFqG4F
DBkST8ciyFoxPSkXL/7LK5S4Hk3QroP3J5wdZKeyB+wDPduQC+P9mmqUNQHSEZbL
HOV3i6JO8gQBN8ZZSQ6zF/i4eWVW25eGjydaBi/m6brPT4MQokT8evpPfM3c4CJK
Zm8NA1wplE6bZV68OyRvzAeteW8LA5UYxZioto7Tkm6biaefnkcnmnR4e6GoZ1ut
Bm8JQ89/rQDVJ88x1IN6XCroZCdb7vCHQXNJpLjmWl+gcfw8sZ++wszF0juYwHJV
/fN4WgrWQFa3Ywg0QZ0Dgtjc0fpE4fiNDLJLWgGUM/IYlU83JZUDW4NtwYdOL1Zl
OiuJx5DqekEWA+gPyTOJtbV12YLvMEWeeB+kVfZUJr0HubscblViUsOLvWVPEMCy
sz+YE68i8aJJb+67H/2Q6kl5p/v9yaJ2/etrqlz0IpHnoyldTujct115Lba/7tdt
TWakTwfXHFEYJQoAvGNcm2SfIJ38kLA0rtO5UrAmIoQsQklrV2PmNzcnth6PJ0F+
5OpzssuzhocfZl/Bb9zMJ7zviqyEOAsJf2oRcjnUNA4TBq65fw442pOyrlsLoM6U
lkswZIQ/zi0GIXfVGxADp8gF2VuLNF6rfV1kUfX+elcO/YY2A4I5B5v8rT/fqI7n
7vli2EQUtNuGqGCfkOmjI8WcqwN10Q2u2EJksBoLKE3j9GXcMVLXmXfE0J0Yis2e
5BZVMw5tMf1lDUjmqbgJBi4VqwOFL2eHpVFBocGV2pukOBXiRBWOhYur0WFMvTmn
obJOeWJlMZMKnQRINSBnKCgfwSDt0PnQMfg1N6aeaaCUM2a96AH+xKxiFM3gCVDb
tduNEAKAj0j/F6t58pGMhmZGl4nbE6kuvDSbKIb1Jlb3k54HAU9Q1dECtNzcZdgT
5M3p9krTKNUFfCdJNiMqh50NsZwgZD36mwcUnqLJP0H56BxcjALV1e1ruFLZEn/x
EGWYPVbFIbckcYzj0AFk8hCMaUef3mYtFhGQjfb6uR7rx/3II7NWWsB6RixpLQuX
4MN1ef9PnK/N1d8+eZq4aCHqsRijmRIHuNX/4RACUau042aUyqEiwB69LLvAoymB
JzQtOMt0tDzxfDQvaMN+F/SVCSP3LaiiQa5uQ6znBUIBoBuqX6SZhgk3c9BGfu5B
ROFVhYM6itXvl18Yfv+btmHwwfHnvSIpK0GtIXmgDuOGvBcudcL9OBF/yl+085Hi
risXZJgU9F3+mUmGTqouGRFVB+dpe4vRZUeHLV5uykl5FpjEBwKpPEXqgoy0MwhM
Pa7DGWEiQIyqjsJk3xPFHdJpVEbCU3Jx81AhOTsbod/LVbJD/a6sc5/8s8XeclN0
MfxxB4re/c3XK44l140QKLLOW/xOJ5Aj52h7rKiUYbPxAelNx+rx1sZaygMlcgyv
wjT5S/k7bNQhKbJns0XygcPzwbCIHSI4iqSLhi1XnAUJlk49ZQohtszRwHJqCkMt
+gDAIS3Q8od9ZXqHx5mzep3PF/235hVUzsnfFhEwB5SF5mt6bHktWHg+8AOwbM+I
JuV+zNPQ351VGujr8GwzU+ecWlmUp83GlZyVzEbc5OHcPj5SJ6JlpPo7V7Cihp6k
+Y99+wYDC/OG53opsDKg7NTuSw/nDOAh8GWBx7AdE24APjaGlr2lsQ6Yzy4Zq0cH
HG1Dq/5ObJq775PHURQisvaoWeO/TZWaRVnE76O1sRZxArsDMeF55UkEsuDrATWl
d0T0rzmF06vPXE5oWktr9w6AnCNrY3ym185u6ai3VkVimuJkY/dwwp+YyDEUdKaz
WVQo0cTfC3u5AAi6/95jTmyhksHB350wIiuvBhTNw6xyBwgsqFJPhfMRmi5CwyDg
QHJkKCmePU7WTXEw8fD2rSxIWaey9tIh1wELuhRTT5VbATwk9mrOL7VayRqOooIx
AMqqXiU4ZpDm+0lZXtdA/pMf3gTMrS0+kHiXPwGzBUhKb2uEO788nqOFf98ny31U
bBegag/MbEnqQXOVbfo5A40P7kk9BvrbTnKlnlkUyqlOa/J8n7U5NSK6jDs2cvUo
AmhRgd1CIagLXQi5arjaAmUvaBPcCj5J2oTKb1R/8x6I103ZhITWwrF1BDWQLCF3
wB69v3OQW9csFNSka/FbmlTDAuP9wYwahWETg4EJ22Xcl3jujK2qe5BlTU9qDXXj
6rHFsFT3Y3qC+V2nnPE4iegek13nljjzVGS4LbkGoHLkVAdpBiXPRpmNv+gwVWqd
U4q0CCCy+HP76Ukm3h/FK55/2O/MavOW1YKxd4tA6h3pYPPhMbb3sdsdMxPU9z1W
L06x5HmTHvIMFhRK5/yj2IfRDy2qTM1lmJFM6oDbHomClGpesCCQxgljid1RrlEu
KIxBiar5J8VAQ3H0wo4crvjEuycmD/OBh85m0qX3fi5xV2Kll34XNTTBl7WHD6F0
8IiWFKy83sx8VI4IYMN/ka16LLxAxgQeU8yZsSD23YA9I/sIzQNg/YZa5h/CtfE0
Y4Kicih9zJebv7YcK384M9AVjYURpqU0TU9lDKS8vEaubiY7Gfpd0tYpDuP4iBBR
kZ0vdA5ra8RfrpOsf3AHCn7becHtktl1oI88RuaDeaP5OHAQ/Rky7vWwSUdrJ7Yk
m6ajwahQpbE9h/HZPUzaV6x7cu0XcbIyB1/2O9KTjnLCjRc6qgiGyo7Bv5/yg3AN
16QRCiGC63bAalJCK5xirGOhF6ch1FIvFs3tyn+Q/jVZz5irzWIUCREHbFvjCfpR
9ChhGWP44pXBiyIOyL7B/dd00bHxN4yrPmvsXXJouHHbfJ7D/pAlserM5RxXLBDB
bMrEhhGNyqH0NlCBQiDu8b9caZcKqavw+2UyAuc+mxo3n1f6OZY+bk6nDvAMXGxr
jAKEjdyKBCmNq39G1Dga/V6UojaDnvQDSU6uwFeVQWwjuspnFZEDvzdUUCzYJhab
R0QBoa76/Gsf6Tlxm8qQ+oOjQOC/dvNyvPZHEpKpofObx0FAEoa6ZEo2KGqrrseC
l0XAV52Nvq/N/uJegrGOAMg49/yWw1Podzv0b0j7lmhEDPO3tccEejRQ+LzRs5oN
L3fAe+ANf5i9qg5vtzYOp03l9yLyE8/RP2ItpSu5o+SIk31lz9FGaI5bAgX94RKb
y2oQ9NaDqWcjPjqe2AuyYdyVpCS7fgHooLpN/T9NlftNWlwU5IMD1CxTjBVgNtn6
x1nHItnlE5Fh+P4zElE5tMryIJn47aMpmL3KQxbmgLcK+gFamKD96yLIwlOt8NT9
PAjnS6ViDWSULg/q/jbvlMaVJPiUjKAsPp1mMUDwkdjw2mWMjHG1OsFo28jXlbj0
s6Y3mCHUOd188j1zQVpdMQV6OcUbLwuuU2IAMYrIFBxRbbKnSO5gML3byjFhwqW3
K+AGqrC2gxWlcxfUpxUezHx53nEGYxkDWb/iKTdtY2hhFJOGmOouxsbLkMnDGhkH
mtnJ8gkdf2vXrB8P/D/PrcSXuoqhl+1pHQ8B3JM/gbu1JnOmWAyI6MDLYv9hEdfK
cuVJn/AmBzHGWJb4qOYRO7q+j9pyvPDY6u0pBjPZKW7ysG21SAzWd6W8FZ6TDQhr
Ij4sKR817mh2t8LgGiE52Q4++gqwg93SIgndDSd4ZZ454Zk2rveck+aaAqnxGTbA
mKnOSH+orZ56NpnEoyOEVHLA9I1uE94ZviGnTiCo2AoYF9kREQPOHS6KgJ7wLMUu
tbENHNmCNAoXoL3IUp1sSr1pgptwLyAzk7GUbUwZtBHmgmJFz/SdWR+Gpsi6TxQ6
fO1bYPKEcJesY3IGT3GcG+BfeDKh/JTIt82DQIt4JB6EBddwKgKG3ogy/pGwnbeH
eu4IFgeZxJgxExkR20KkIM0kju+1tovvptN+R63I7g80BNtHICg/ePrbBqxTmEkZ
vSdZF+42UhJBzP6Vo1fTorS6f8DNSy4/E/43ermXnhhhS3lUB7IxzWyG/T86JPiy
6JLAGY/TNWbKa+lrlQXyux4qIUiTRVDm7v0iTgRzturudjITFjnd3PshqvWd63gD
n7dYU8c+P9aZYUgiZ6/EA/MB3ChYF3bJuJ8n0UptkCsmISLA+mGQe3fPlX84MH9r
LGgxqzI7/Ql9hsl8PauDwZ8kE0Xa2S7XvOe29BLtdENS8jw/jPQ7tx1lrfpUUBkq
pHQusZzcKjee42TOQsjS3JBiTJ/DMPEBto38i3gQt8q98WK3inFw50bfY+huc7+J
wEJ5rF/0HkoH5W2zCcVnYKLaevX5NBxe7QzrPrkuhGGTl8EjvJ2S9JAsAWgaZzhe
esSAjok3b2AkLPmFErrJYKiBqvf+0qRQXlO85pdwAVKzn6z13FcxuisPKrkAuGtz
mEw4lKGmtmP8s2SzR/ti7vIwnZ+2GAlymd3O3NbP6jNWBUcjw06DUkWfZWphq9pg
RbhZi5KZ5/iOEX0nB/GAGkBzkZqhB0DYwphRrD3lIGRuor18wOuRAvcLwyJ0SdP+
+fssdS6lrWNwhD/sJ5ZERHiCwfewtJ8VTK9ZnGir4tqmSIZKzqOIB3Wge7UVMihk
+eJA5SWB8E1k8I6UG/2LJPPBP5E+QfWkpJK7pdULKNxP5cpjP1FuW3OzZoTo77uq
DPDwViMWt4n9/r+eZt2bf9EXvMHgtLQBocPbwZX6B3RvDyS/gJu+9e8rxUorenVN
YBngob2+TC/GUl4t+Sm8q+G9V42Vu2GoxCNCv+IRzD6zXitdy6gkB+fvJ0NasIV3
v5YxvVGOp5rNXnOe9/piy5Z8EfNbUMeAUlf3CoTex4F8fw3pfR9y7LERfulE5S9R
Jj59/8Ws5AXjiWOLH2neyTEMvrzNZ1LDWKZPCGfQABaZHyHYV4RrdFW9fQBmEdAd
snntvXFiccKSNdwHI7iHheeDRnqhWk0Kk3vURS92lZW0FE8gfa67Hlcs6usYj0kl
fg8zQ8FyO5F0iBeAp8pT3CyNF8miFEu5hhqNObCTR6x3FsjCkNUy2KtHyPsfr4wE
60NS5gn4L9E0Lp8PrfMvLzuoWHziv9wCtqEfUuGSytQXf5QZ2q4F17uM3IVPFXb3
e5UEKWxqngmlhA7e76NdZVHUB97GU0gE1GrhTPzfiTnhGncceArlRVUr7v8JZhh3
XeB5uOlpgaO4VHQShJtKe56+971Ja8GAuBT3H8CQYdIFuj2vvCDsQRNql4d2gOBt
xbjfhHicK6eSIxQnipbEIVgq8cdQCYaNSeJByqa3zZsI14nHuIfsfUCYC2kUZz05
pbm2JMwl02ghOyATnZq7ZSbDApx/mjsVdq3yZLCaeuRrrupXey2tmGN9LISP3AUa
/6KOw1oNksywJCjkzyXqer0Q1+pfl/mVrDRIik9ydedw9U+MBIvKItqak7j06K63
aQTe1mmI+LhGTWQTU/h9dQ9zt3ymkghehWcWtxvrnRzZK3JX4XbVRNaF9fG9hk2U
rJnl+bXn6HPGdJWNsUHd6FbpeEAMtOYJhIN0JcCrYqP61FUkf/Qg2YjWKCYKYap0
z8U8EYJUdljipLGb9bPWwE97/sAObiCDp6DksGh0ZgA6potMxjd8xBtY03Fo3a1H
EQB3etF21sUJciUh2x/DooRcIc0cK2pA9aPtkzIveMeUcY5omrGbdUVvB8WLvxS5
cnoh7XG0m3w18ThsrfFrBizz5V1FuLn7k9hJKIw8uS2L0spgXVti2Aj+mCs8OwF/
cYFiHrhnbrolT5t0Ilux5eVaoK+Pcip3lRyqSVWjHrIcYXuxAleZqY83Ls53JT+v
B11X3Ox9AYpYXFzcptYndlahzt9yUEhF2gMzzOOOk35RI5a/dTLmk+mjRypDqC/y
FIlduLgmaicmwmtjgyN867qXHGhCHtQlqqZndNxSoF2v1PrNVsVwU12/r1UHnis1
0rdnHruZp81+lBbmQJcP6LCoFQk7Q0UR52FJiRSpS8eAKu5+zG62dZP1k/7b1XpE
HnlGMKlXedn5QMCcmjZPTEps6xH90uvpEvP6gVtHzoHI575zNJlkI6Swo6FLTknh
ceUbD7XEDN+4CXoqX9Gp3OgM7zPTvN6zI3eOdlr0gX9C5x2bEWNIvB3Yfo+qTtlG
Kt6hw+YHLvmbetThoWkklEiBeSlcMPCtsR4WQfpif4l04dEenL/IXj3++V+ctXw3
TZ2ws3AgZbyhX2fQVt5kF1eEsweEhk9QsUotB9d1TmkDUyu+Jv2QUaHwyUXfStwr
nAAQUVwpMJheZ4S5zktf6bGm0hYmGEC/fcN60vocnxPeOLs85FO+BUP9I5QsEWYA
K523eEULv3v9BqjMp5LqBpxXqx3ERQ6nrPAxrFIAB12KSgdcVwDm99IdpM51V84f
qqRPvFiQ3glFa1mrks50kv1t2KklnQlw8sD3neqO99QG2/aX+a2UW7WkGrQkPvoX
chCTz/bmaFeFgtgNuXVlnAFwM88vStN/myoWWHrYeayPCQMc6YYC9XISqRKb/rYw
YKKzjVPymivjKms5NSHe0akXIlHQdtA3PpL5rhT9wpktlfK123lZOWMLxBAUVA5V
KGIez/3agWGBAlPr9scwsDQj+b5y1Y9VsGE0dkUe6Ibww/+yiQqwgl7aXhSr89mh
NoJoxW3u2EbIXmLG3E5KYVjbxGfK/edex4RKldFZ+5z04t9ASFD6Hbp62yW26hwu
VZpGkguD1cvB2FD2zfym+X1lSBUYbpwcjrgcZSWNO2w3wkW34puVVFz3lYjzmTF8
wUS7L2w1zDwRdL2LOgpe0uq2fjodnDnquWug9mHkfwCmweyhStE5NUk0WotTXQAG
zXVgbbCtfAeNGb8MJpX/rbYIXc/bobWbF0atn9niUDSAfrfMOlBkDrP2CbtuMW0z
qOAMYPHh5WBSFSxLS5Z2KJcW/iEzDbVfp4XYrcQOEVvUnJUkky11bK8FHE+gDpEF
5KZVWUDmMXal64q8kC9ywUo0fDyXhoKPPEwHfPf9ylNaW+6IELkR58E/fUuylE+y
KsQGoIrFPrmtzr0f+uvMo5CHiupbMEgfRMjjnTeRHb3GlEkiXV59haftBIWmQfuJ
Oq4RR1RCM3VCWxmdyp4+fuZ6fKitEXtI+8SO6tI2Mx6V7h9Jpv7dJsAvXhD9k9PF
X6BTKAHThM0Ozgb1WOnlPIWiLnSqvEcR2g9mM9kfEmuFp3CLZrRMl0ucWgVybPpX
FKsKwn07CPQPEqJZBNp9gKSqrh4XfxIoVjaLM78R6wEiHz+gNKjbLrPkt0LMWy/w
jOCp0qC3KYxVJ7DPPbX8MXszTvOYNPa/iDHQgadda08DER+p1oGQaG9yS2j0H7cq
6y4QDMe8wfCYUReVHL9FK41hyXv+L6GP22frSaRBPN4/gXr6h66S6rcEnaMC9BM0
rTMyFX/rLRMIeW+fHC3MKfr738ncYTCkgCJdTcx9JrvSzROqX10ePdotNONgD7ce
jDLbercO60PXnqHpPCOeGIecRAcL5h06WFMMYn4+cHKAsa0Tfcf6JlJVAbhKeVSb
WgQ17mIGvqLFwEqXJYFi0TOVkpWBw2KI/HEL8R8UXTp+Eh/tZ1MdNS31s8100juW
o9j/VkhgjIdTONX7Ss9pujImwN49wAcgeII2auchqSyLqXXgI7Ze9DaDpPgl2L04
JMbAr/e9kC+3FHQjbxZDX7WMirPDxkadaX0k0THUs5Cl3M5PWR/4+kdAbu098p01
b6St2ukNLLVAz4aC3RsxbWv09S0b5rpkUFS9u9t7uI80AvkYPAFtGORTC3z62xTZ
gQOt+/d1RPOEW+/s2/s6rV3QJ+sj/0+jp3XacBZ8FWuH4A8T3PGfCZhCN5im24Hr
ofRz2ONzHPc4dA2El0ENbQ0uTgt+21zGHp13CHkL9xQi4GAgHxXZuD8ImdXLbEp4
wwCFdxEIRJeyuqYn5S111aRIqZTBAx7ttrjExqga06L1Zn+wOa5Y0SxFWNBybU1c
saTo9cr94fP36U31cwtIRyoUrTI8z/vlXJwqH+aTLX5Mpfv1F2yD/03Y62Eb2ZAr
zhc0LQUPxmWE/BBItKzfqM7zqrcfyy+KPjaPfum+m6qTCanvZfs3Lv6UL36Kk+Lx
T6BQOwMgLb1ZIZIWXaeYEVrNXYrHAQIxvY2Gqs0WdF/2eYCNIaCUCXaSq5zlYJ3S
bYVcUtZZHVWFR9cytE0A/fZOR2uu7Wlz9QWm3GsVbhxZmtXQ/FaNq1WMO9uaT4dS
R+CGSgdMFD32drKkpwZdAuT8KIIkuREVCa3W8qqb/qa7g1NxoJ1N/+r8R6zAdBLX
914+//emfmnyKLy7tV8Po6dqIHMcNo1EMOFbYKkXd1X/fy+Tnfds4obsWxuF1CcE
ohK042xrSvgyZCEUUCBLThDOzHGgkBk9/9F/Iwyq8IWzzn58LxIqIoUpgHac7GNy
ykW4J9Up2FygDEz02jv+XLfhYqpl30cdwDvbUMBeECDxgczCzWiKIDuTEaJX77Wk
bp3DUXBZcKKUX55brAOIShZG6sYohxPhMeWNoZ+wAVsHuQskRMMThuoYE9ZVnN/F
NiVf3Zphxc210DD5loWwv8aRdKg0nNu2T3gktEx4vXMi9vuOUfytUp+qD2z0GG4y
GvWDZuDgzuApoovH9jIZHtZGDdahsGwCzKRAWYBQBpDJQvRtIODOL+ZTjH1gfKhg
ABwuLC9uQEVdOrfGRNqV6uPt3plDPESzFbU5Umt3xb1PpKdSfLDJakkF219UGO4t
TUdN3fa5JO8y3ZiYZ6L1DUiqFbidTp0vao2MAm7400Z6W+AGbwCpgj1ATxhtJhhx
spQLfWwFLcCLTLywUONaF8EtRfrnxbY9EZ2ozzG+ytmZPSakL4n2cHREg+ExFb5m
FDGSfVpJAHbMRaSib1Fi/ZVSBvKPRRjCaiIwjJ8BNLJdBrgwqz5Auj0UB9IcM/1E
wvuO397B+TOkisnMEoSSOWq9Ixx/Ckmc1VyPMY3NQS4M6c/9zsdu+g/1/SiLg5xy
ohGm4X5OIYH/+5aLOiDJaw6+iDhm3rNYCXqJUxTPBSBvHcgjyzZYJj0ghrrJ+A/e
Bqm/ykoWJwGrXgO4KMZwECMJP+NXABhA+u/mfaPb4zgYH5a3K7Oe6wCPBf06jn2R
GwiEM/QrU/ctj6Q3hS1PjjQX/ORuQzoJZWo9wVUEHigyRI45nGqBdxkLKVzVSe1E
w039QqXXCmRu/was8MqTm1YcUXMBDvqLMegfDFFbrnPnSm2TH14R2PwRz5y6ul/V
DvFMQ7QIR5mlxbuSrO4X7cMRZ4r89I55xhzLjHT7GTC6c1Sw2hnzok02o713ki6S
+djM5UI0Ex5E5W47cu/cy141DSLPs0nSP5kLrrVJtKPEds/deOsVnCQgB09JZ9zg
Vb2dE+3WQFzqXf8hkJTmPynOb35wkZyhgonJ2NgkbmSGN+aKKusOwJCYCYvPkNjX
Sxw552jn71106c8ohovzySrLyZH6e/5uzeG9aQWO0sx5dVB2aL6JCGM7Ud8FinGU
hwKuFKCkY2PNteavDS7jyqLZvjvle4wmgOaotNLQ0D8zBShwWp1TFsGX06pfY0vx
hUGh4lY9tOyxQ3kWLnMDwYp7TsTCO4F3Pu85dInk0Vx1tO3eUW9BmbdggeRedU4d
Hxt6unbPs5iiGLLhiuAkl+Lsr/sKvi0BS27cRqk6orhvqGVtZjjG+CNIhEzUDLzF
Xrf1KQpqDibVjErk57gBDWursgVkSFXoa1PeQkCJa0Fd4Q2oRXf5+w30NQZHlg1j
SQhl4d3zmLqtMcrcpj8Eh6K5LexLko71H0Y/N+mkouiZa8XdINn/yCijzIXHDHJ2
/Y62wr+YZReKmbirIOcuB9aXdhr4zg5cEgpA4xShYdNe/GAJKMIK14zdvhVSAfA8
99TVdoBSIow/0uViEcJ8Qq9jboweDsmlM03Vgds0/77E370PeJZHkVftKz2ty0Vx
CGe9zQmi0RfCogsDskKPgW4+Y/OPaKuRvmydQV62oMP7CJs75w6UAKtfwgM0XnXW
nCICPARrieMIQ31A1q5oMIfEyX1qBc0ulloDr1JzjkP8AJ860GkQbi9T61MTCyf0
ux0VhnNsophHjeIeCuoZEzkJcYe1qxfIXHCuQlKgX21DmWBuoF6UCW68wV1/GIqs
TpKYc/b+o8GZNFC2IhagB9DCk4wZhvfRPZeb2KdUnXrPrv3sgvHecvVDDrG8pKxh
hu3Ls6QUws7ZKhsfIsC681ly/jVeCzjnmGXnA6LIS7M27cRGmdqfaMrLSh9P/py5
Kz2pb+Dgh6dmPocXWhQIVcYMIAzsL80s9kLLDzBQ+PEsVvG8J53ElMi44oex/BIB
BkYjEPSRdNnVkYioZIonRxxn1f9fIxzXsfIPQ0CueWlJPfUc6lmr0zsdbfOs5q+b
0NPpbz/G/ywapN8M0nU5sMvYEuAgi8f+wYhHN6ruDoyTvH2xBoAy9wJCis8FLFhw
3titqulS+hOCugHxUO/vgEBZ2HH+241Hrq52HuFQFkbOr4qLOPheeE7KjVDSa6c9
HjO52VTG/OD+dZFw0FcDBHQTM0whorFDnEiwcZI6lLM2XSYDqY0y9PJKQhH9qAxi
jAU7fadDriWw9aKZ3e2rswRrdpdr3b/6lah6+bDcgVynJd6gcL8DlUiRUyE1nlDm
xvtncD3CSdCeEfw0Wx1lQWgkU57HCzVxsiADRW2CgoxEWbK/9gjWBMZ8cwU6datH
54Y39d68Pzkour/Xa68pz3djRqT4ny3KshjE8JT2gh4j6DzBz0ShqSKLrhAIp8LL
NcvwhwOubGiSrregJ72J+gxnBj/eRJNbQVW+Dfv/kDOCH2GmbiCxW0DODDnLWGLt
uU5Xc9uDCD78Blb/jx89/pw7+mbSZ65I6ihjo1SkIIP/hqvnx6Xno1/PSVs5iYr1
L6mssvu4g/X8Uq0WvORDB1Cpx2+41craTA0/zDwAiKN+wpmPRwZbo5vnh4h8+zLO
Omh69KmFIK7zFpx6nWZM+er0QM/e8n0jlwUQs46oqxkB/Oc10XeqD2SEG3wDB54b
ISFGMlSyEKRiYeTYNfc6CbI8Yfnz6g3sZm1M1XATgKzlIdQN4I/kC3mtaPfzRvh4
4s68pByyPvvQ7z3cWflJkJMhY95iJSbDsmPO/0vuQ48wWHPVMCveJajGmnqeMtvp
T9IQWO0KkWIR9X7G9Ap9JuifUZ7h6DQjxJb3kVcLXVqb6q63TKOyHLr0UF9LJYSQ
Iha4Bh6Y2oOhdvQhhTR1BF7cJUzTBlkrOZ2ZPkOuH28P+kSLSx8OjWt4krRvR1vh
UYpEIQgwoBQOdD8+fwbMQGDKK0qejPZ/02H63pQeh50GwZhzoxik/hZ+cWmpRU1I
fINMCqwVatAUoDN6kLiGAqlrav8B2UjqsnyLEQ/5fXhrQW4gU7XzMZQ8irhJ3ZXF
kuXIGkw12EqTIV4JLnTCQc5a6NhCmZ9rNWNqeyfnQ8TRciwTDn6G2+Qxc49/Rsks
nNbFM79p+2fTGNRZ48GJxAX5oasNafGrRRe7EP7d66t8IPoO4IgXg0HqAjbR2GYe
rWx/eWtsMt05ih8ThTOI8Yp+nBmAJ6uj6LVYp3Y53E0UBErgpQNScZFoQVxmCl3d
Js3ZoHQ93YH7xMk1HxnCCZ7A2ttt+Kw99RYIjuRR8fMHlEKW01ZOpiU7w1GDhpHw
Q9lCHF36QnozYkydsvvu2pr9De9lrMjNdgvj6AdgZ4WlhBirSp4ycWzdvw/zBih+
67CFiYLUF1D7i/zGDTSLy9SOnryPpyKKHq5oPzctvJtgCZZT3TXWu4pLYZbBLtUC
GY4f2mJNFKhw2vYcAdMCMa4u4my16lk1M2bdtrQ5ZmrhJ/a9j4Kb2iyYRqf8e+fv
uREIRw/6IPH+pzf9fwVQhB4l4Wb2pSRhsVU+ZV0F4P5H79ReoXK3aNyoIh6og2dz
2dJwUZyKYS2tjFftk4WMpSASUltWnYoMUjUyZnutxnv75sxqu81DcKHf5DpSxymh
GDucZ6P9Eb1mZFQXbvpSaeFiU8eKQrUmyrrAGke7Gr4EU7B6EwR9vK4Zim5YafQM
co4J9RS3nMH2X3OurX7LI2aA6x0ixDRsFoqQKZKzpwq58ECOW+j4QsdcfBCRtysQ
w/YAkmO14/pj16c1vC3+SdO+cQ72cxKJR9Og8GZnrH8Cm5MQBQ4Zv4ek0pAyMUtM
cm2R+DtuFwwN0JjzvGjv3wTAJVrUj+ui5SEnysz5QZFEDSf++myiPVGzriI7yaAw
VPDrQdz60/U9O5lAh97eFOLpyB7Bfhc9ZRmEplhO7S9QpGFDplRU/Gb2h+S/AtwG
qUfbnLGxh3hsTnKaoRSCHU9fx7DIe093qC8tE/R/RhqT1ORo9TqWShERpuCbuKvM
qOGgbbvJqoynWE/kXqW4UA401KgTjS5c2v1XT3cIJor6ZOhGeKTXqC5RlCuoAo+O
g91JQaVGLyxxsLnFcd1E2TsKWxLHpvbQ/SaTIr2lcd3KSACEU5vdAEmlS3/g0CQQ
CDK305fhfPqpNAHDibxUjE4MdnHMbtkPUzec5Kw4ETw952+KagXZzQtZNDn97WYZ
jXtIzvdPPImmTLi3oHh17AdpCHaYURrRN6iddrpSWkcqFoS1SswLWrbxbxrmiBLl
5xszHkI3rPlWN59PVUMEZGdvAC7MVQGy1bth2Q38h3PAK8/n1e7cH7DlcRghZy5G
h73zyJy1cZI/6BYxM83MUNvFBwNmeet/RQQqtE0XhsFFi/vp4IzbkStAHZEvxzNP
nJgxVYJaj+HTVkSQuYgaPsCXDrdEPsKTgY1WVv75H0gOkfFVKzpNqOSS+FI9tx6A
EBEz77wT2Xb4gSpNnF5lnA+NhvvdEN77kwmLG0GZbG5Bh+SHDG5/LY/ilTw4Qhxy
qt9SDSgVtyKznCrqQb2W4h79t/OnICm4Ryv2kY1fWrlGKJrGf4fyPV5l1jBUH5qq
lPSZ1ySzMN4WSSIxOObqyhbi4WJLHeWjoF59ylQj2spkVSF3DZRHyKlyNFEL5nRK
CXFvjpMP7ZBh0k5AUYQe7PpUcWrVy3QGOTNZVcY5m+62+4w8Om4tLf/wiKJpfFd5
8WhIfLRtfgCHlcOmO2g/TISQZumQovxzeYS2ux2CfI9RH6UrUZGhsLlyV+r+Iwo1
bFnV1uwz7o9KMgAhw3mFIiOKkro6JzOQ+nmR3I5RVUKTHsu8zSkpwbbwcQ4G+qoC
U+wjkLR+fGSXQkPBz/DrwZkggccTWIaGCQiIxcvlCVX2yqNNeTTCBrxWWttSGxr3
PNcTMiE1ekjHqojSXcch/4TU/7WYIEHZNJ16tYLHVR+XpumxZYvqltnq6NtwVDak
TVco07EVrz0HoFB9E5GTNeJEeaQi6DO5mZ+VmIBcUklEpEcAeToVYsQdyAYqEfq9
M/pq6bLTrvs8207IyhuqhdbOcalT+dPXMU13RBBZqB05HhsJTusjCM1Pangpy+gZ
5OtWhWVdQkxyZCo4TR2kotgnlayKzquZjOolON5gr9lM6M7D25k92RB4FwzyFyj+
Oz6ddZdEgUphIa2O8VveaDpPmWBy/wfvnKmMtVqeQ3Gweg0wnQP8Qm27oXYxd6lr
n0+Cc/ffWAg2UP+/iItAXrn6YWmk09snyuY1/3bRN0xXw9LUrPOQ0CMEGc4yEvAP
vYxgnF7kNb8frv3n6HbNcEV29LXdVfxuGTyqLXI3tpE7Ki0PZPC+15qbYgz6gvJ5
0bRDikqWgthgH5LYsXWPDKi/7yhL4upEueow09JT1hDb+2SMzvRz+hOT01+HqP7J
VzRbzUwYw1/hDgTWhZOLGMSr87cm+CGjeIvu4fAUlxgrSu8AQC79PKgcFzsggaao
9H8843QyWZ7IlYAet8n2BGlM2GQEXu3CxfKCve5GAhaXKh9tiYQwOonC8rxyuefz
CUYLRdTSQvMEE2aBC+6uWiXxBWppr6sJsxnJHrQLCXRn3P/P9/FASqXVjork8Zy0
iZW72BflPLOaJ5mzmHLK8U1IQk7ngpHn+r1uzt0GVX2qMJ1AU0AY5K3k0gF0NIqC
lDvchBYl4P1bhDI6f3QypxsSf0Ubxnidjtv99/+3iUasl99b39Y0sMES9yYnak1s
jxikt3D/mU6jNOh3wPhRehg5ZBZ/F3tio5NfMnJCcwondKzSEm8kdmYtV4C6TcHG
1MSXqvIkeyoWEgv9oY2eB0XANhjUEuNkfIJysg/7O09I8ZsYw2s3zeMnxzdxZ2UZ
bqhHH1Xm66VacSYPIGZORWdcUjsbig1Q2+hk4uuCYyKyPQI9c86WvNpzuX/e2K/9
tIgjXbzuq5HAqWisF2WW8J2Xr83TS9Q8fmkOrHV0y7k3yuZfPWcwhT+z04TQ3Utn
Iy12Cv6C8Z/SGeDS8rd6ECc9DQEgrBOYTpNXITU+rPibdne5J9Fs5ZOLORINBMTv
jCQbFKR3wgb7jRvdj0muyGmnmClwNKBoJktnNmec7L8Nw/OXmtzllk4t0fcOnpdc
yjW1iGv9DSs9afAjRbwdf85TqxwLCdv68h1iO+1jud5Xv5J43TUlkZW0dhWWSG0a
7mPp67AMFcP0djLDhQKmzZj67nr9OXxQCruJ6zzASNXvULoQfN8YdoGPjBGnEPMd
8wWbkVZe17asFTrqMdcfC1XKA/5Y4uxgBfWlgEiLwxvDr3RowRhTXrK0GV+6vWAK
lSzcwGxXFUR4RmsZWbJlSQfQRIDQkYa+ZPmvaWpumFT77HMeHymI0vUYe8o/XLhK
ZdiFHnlZeGghMb/XSyNBW+2IKg8//KSvSzz0upodnB4x16qYZ2bSpaFFyoqN82yG
t5seo3OXE0sMqiHg6Eg6Ik4vHlOCnBJ7/iktpDayEgEy0hu6DZNqgmlfJH0IfTXC
rmMPZ0Z/U5vOCFOtYRQFjwl94pKtCZGA4u6Xwq+fF2SJPgs6adrKNygmiemjLDWv
f2o8CkXkyRP+4VhRrQbu8B4zubD6JJuzV0Z8KsX8doHpOVI+tVvcpM8Fai8uqAr9
bP8GiDVMHhtKSiEJUUawlWcMAbU7/dPqiNxAotkAvS5izpxatorRrUm1XrXr91Hq
YMbHihRBv1qGUNq11zs/YU9+aGK8tasCPM92nR/I+xFFxrdZ+bbbmG5/jZ3G6Oa7
RE8FHfrNcG0axx7F+h5TlWq6wDIJ4OABmcxMaTyQupAUbcqv8ZXG2zoWKhJbXasB
zj2RrOtI3hUdS4k6hwSMCYclNUJbIMB4cyDsN0GPH1JTqqOntvHoSIJqxMUknUYV
A84JJZuootyzGzgoXbUBfYh61lFT8DL2uevjr8nWsqMne0BCU82UpNKUjgdwcWcC
G4cKSK5rEmYAASlP0G+fualXOWFABXUdywEcEgYFrnKPLRbRoDPYU6mLqP/dJV3P
ZILpJK/im/bZonLgn9MjtIJDnUTnI1c3IGHyaPFNh72jWVbhg6/NHka/krs2QkGD
WM6bA81+ioPcx241EH7/h7Ih2ry2f8fx7aDYst4lWjUQ9dVe6W4MWmBFrc4Tpqc0
NSoKW7Q01CjHX1sqa16fTtvjWuje2tjHw4Aj25nbfnSOfDbR5H/ucSl4K5zIaKns
9/7OFO/DPdk93WdfHq6qvm2MK6QbGh3KwFGJ45lWVnDbOwyfXpfuhRN2EWSiofOf
YoyqyEiCbd7aFDK1VwBQr8jbDVAvw2+wichl4ioPOMlCBDMiaxb/FzwTeLvbW47o
QpbmewTt2M60pNqsMLk7afLcszESViT9IYXypGNNtHL97S48pv/J7N9Rwi5B+KlZ
ieF3dk4uF2tz6qNDgfrXaG2kXA+xT8iA2P4LlboKuruIlzSlDAQWhKFW3p8R/Ldg
OtYK77Jb/UKGt/YJNOGn4Ncx16gEEK6lXOpdOSPbvBEUbWevqdfC641m0fbW7ZWP
rpMcTmDjJiI2sGTcWKTwuHE0bfCYVuySIAQmYn8U2NG7lC+0f78/ohpxgsYeiqo2
YcqLkeAw0UQlah8crM8lTHpb9Ol73jSbifFLVsm41IFMJIf95VsOa+0Rr+0Bu62V
QhX00Spt/JdDQK2+xDi3q1SV+NGNcrsk4vo4lcAZoKigxkED+h3ov9ZHWdr123ta
A1andRqQPNxw9MWLMRXIZlwORhfUlYr2IAkmepB0yFJPlMQX4vPD/3JOqjhvTlKq
9Ej5RR4ZIatTDWMK5D1UU4JZUpSpi3KWTwtneHnSWwOJopwxbUvpJzZVJ2TKyC0M
OEYwFxSUpCLDjnjwA3acTqKvewCcOAmyRBEPVBzrl7vWaHqICKIevSvSojL1UK9h
cgYtMYBmEet3nn1G8n/HDK9uWjQiASp6xX204A7KZDcKtoKjqcLAHaS087tWiWei
9urzpg+uJXPqmnQ3Yc2xbnmhXxDL/XsoOl5bTZZTYOPD46DoABgStOPH6G8iV0h5
IyifEYpeaz1wdmqxSATWmfbROd3nuqQeSuilr/DPKb2zCAyHDVa4OfZDB6H1NIrL
c4uJiHTJGxzaZexTCpbhP44Jw/E86+iziVnsXEOnQoYekt1NPtHLkPCYzQgi8bVb
dht/Ce5Z9P/blGTBqKopueUZxCW6yma4pPPTY+9rEK9VfCQYT9zO+Sb5mhiGDPYg
LS+qxfN9OkNboXCLtFem9w7mIzalDWMbySDumJkN9nHLZ3eQo7J1nPNlkvaJWmfz
m+OUR4r8RfvtnfPQLd+VzIKC5kESRtLwW3fuqG6DDgf+cpbrpOcOZ+777XQCEt2z
wNQZxolZiU2hd2fmi67+dmbtWlfQ2FjpHGMdNTLw8KRpRH+19Mt1XwVmtXImEkB5
MxZLrePN9/Ca4f0zHVV/zHAQyRd7+tYenPk9Eh3CEVrOHD7Ss9IgeeZxmX+Tukqk
qiOelw8lptThfYfA3ggvGN8OIe9rAFigkxQ75rySsd+iOKvQt8y4NTJOjLL0rnUS
TPO8Hf5WPOPpO2+5nAx0Js2abJ20i5crQuNEvXKaL1EdBKL3F1zEcOJ9Jfktw6A2
5tk6wcrHtCns7Oi1N+9FZKRWpXSomCcLHUfvQhnHiAXD/sTaAqSvSEBnQcoYruGH
JQBfyL362KOarcBRpabY9raVZCgry3lLpKPn7h2Mp4awzeyeJRj7K5DpkQx4GxQu
skdN3TmvEgFzwCpWQMO9vINYhcL38de4zZwWxy+dZ/c+1CsBHc1zXJTr62y0h5J/
VpIxXNQCdrQjYpv+D2tTTYivlTz+lZuUQXbaKwlE+FZQ/NOgV1/BMAaqa2hVeCXS
9+L+q+nOY/jJMEH1iwnHGw==
`protect END_PROTECTED
