`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3WKX9qWl/P+Y7v6+Z25izWvI802L5qmQxv+8MczgtTP+MYeWywaipr8pZKzBSiCK
+KylYDwo4Wg0LKaV8uYABFPTDJyRXabDIsz535GZ3KW8e8lKIMHSERlGHeH8NCPV
YOxbM26fvoXJQ0uVSlPnqvXZT4mN53igDS6Th9HZXrtkQgUb1onxZFfmGo2HT2f+
DbArNkaWRTo/22Dmhg+WpnskU7GGVWccaNG/bEJv0rFC4Fnevk85dd56K/Q+rDy0
pWJ6pJA8MJoPoGMrl2KByV5HloNVqx3ScNIFcAnRT1WBo4rV2Aj6Mw/DjWR3YQwg
T1iy8qm9Cxn6fnOtp+xHyViG7Vz7Qxu1r5Z3VMhT/M74AdkdIegpkAz0YoOq8Ju5
wjbXJp96NkHUELHbOTAcZqITF1kD5cHj4duMjWagw2idadIY/JTwsR6keGbjoIf6
ki8rJMrPaFlRCU5QTw77yCU1diKpRT1T/B99pNuBQdSawE+U2MVgPOGtqB4meO44
`protect END_PROTECTED
