`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DJFraS69xTWDfViBRQOUzQ6EFqkPsU9ctJu8JgCvDazBQgnZQ51GswQAXLhly2+e
DBg+vV3yI1UQk2oBPQSXjGug1fr6dx1JAmIArHTZeqt8gRLvOxUTT9whixaAVL/e
H7y89hCbEPKrrjHJt4Mn4rpUb9cAK3k7jcTWY8BXuwkjEN5AFv/7jNfJHsCBkoMZ
5m+3mn3tqvUWWRFzbPEkSzHR4puaw7j8EdJ2EhvotehRa9ATrA5da7EHlfFfMjOU
1DGz6XnB/m+GvjJgqUAxv1Yuom81ioFeABTGOG7r2eYe75NDRzpisG2iZBfcLCdO
qamr3yvNKPQH4Cx6s2+ket0W/me41nbjI8ewqq1fDAPHB51ej8j3WYvdyjI4vqXT
lJj0ecNALlHT9xal9ecBTN9hj5iKVkxBdaqbcFgAXU0B5p6oTpN0e9zkf2ZOF3pc
VGPW8gQgFzviixmRo9/lMtUjEx1YNxiDIYsqysmAFJwMZmoCOV29Ds4Fr/erw2Ey
YqPTUtUdvvSyiTRLw7CbP35YgbWC0cmDjxqIO0VYS+d5NoXKJ8rNMtjfu0IP3WvZ
L/IeL/2GRUKd+FVuTPxk/Ctbsy8+JqtLjK3umIVTL96bZmLQgQLVyJiKLDNNC4do
7Y2iXHXhboicD6u5auM3gjYy6MOqf0dzuZ6DnPdPHjnDFzI2uvVWG+ItK5xmFkEz
8Q8uHElw/WoMVmxWzucwbNYhGrsqp2MYABA9IfyDgAe771xfjDTPcqjCruV6R9RA
dIaYz7mUsJoymd/OaPCuxU4OpGYNq2o3Ll8rXFy1AFyKrF8CmKwssYrO8xQ6pg4K
OTXkezR2CR5pGB70T7sb58/g9wsIeu9nz43GVCgQJDNA4CpkCg9wnyF+MElLwV1y
BxEK1tpj8nNUF3D3/Xgiq+lAI9jK6DW0pKdvpR42dIOd7BUAseF8mTcggj3c0zTY
`protect END_PROTECTED
