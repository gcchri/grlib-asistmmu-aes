`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GbhZuuy0kLomKPvPyg0GwoHpmUCp2acBiF6u0kYiCtr2xNY2Lf6PVhfBvhVwgTfS
NKNH40qWTQOZ8bYZWYStvx4+CGOk393mvyVXGVGW94K1MfOtVsnGTuKvyA+HswLI
SJ9Q8848IP2PdINZ91Xi1MCxtVuQOduT9RbpVaK07rOmWZhqwOUebXo42YbrHr6p
Rrt5efqLDgHLtEuJE7WK3AdkQ9Dg/S/0NTLN3bwAH1XvcLruni4+yZdiLu/0pdO0
J5uIzDn7oUyciWh1bWeNJtqURzsPG6FlMG03PoMB3wyr5qkWlfI+vTru9QKwjxJD
MFybar4UN+HWjA5dQSed9TXTRelgIaOCdesAYj5Sz/G9Zlqc8aFvxk6wtaLAilqE
IwL2mekaP3bluuSgjK8sIxA7KnXRed6nr3rX9+5mwYbBzTXVtrdcpcoxZrd+9URz
5CJdXwu75NsHJNpOiKF2TvIaY42g3kMyUYn1TEm39+vzNrwotIxUchjqXDXPUnMs
8Xi/FdNo4PbKwaZb5j2Pm/5OW2/ggTbFGzbJNYDmGYcU8maNGsWiLyoZcxADbB/m
`protect END_PROTECTED
