`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tts3WidFjhzhcbTtHPaUak8jgbaxB9BnFdTTtu9W8SmiQ7zZXLE5NCenHi2drBK4
E3fKXnDilk+/hyb1RGkh2VLcmcy7yAKMQ4EtMCH8c0JSlwewSN2pCsOg2hOjVUUK
TsdEzxUEdWuAq/1IzaOAsN8ufucSYbQ7PGfspZPp/a3W98qrXs0bDw4nbtnGcDlN
B8IgwcEuxMiyQapzY44wIHlo8vnxBtXAxqnQrQRq0baEUi2bwftAdDEMR2UeVDHE
Wex3tbBPwx9ssvX6y88hUs/FPYH2smleyCuxDxnAZ7PAZ5t1DqBpEyq5O2whwRO6
onXr4isBjOib6KbL6Zoz/lFsVH3nnfCaW/4a2knxuJUD+DTNu1u2wq3Mq4zmpfG+
`protect END_PROTECTED
