`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UBg1CJDPuvW/UYXF0k5TfPXEwf+EKbkF7B+edYReoOHyFlYdWHvNVbg12OTEaCVb
3fNfnAueqaiKYenThccwt0EJBIcdApj6fJmECDmqWpMNHY8NV5kM2mKF7vhPmYzQ
F7I2AjxZtoCntqZDS91iQx2fxgw/Pzh/EeXzEV++m1IEyPgLbQn9VciUGKGWYCJ5
HGSzTLbe4u1jAayJUXvcF4Y2Aea8BPFeIO6P2DRhJKdJ3F+n+P0Xve5O9PFnMnCT
Oph7ln8EzfbSTdQgNCvTafF7+vHMSVAiuZcuKrhdjYl0I/gWf+RP8+sXctCplDBC
Z4Q7Xg6A0PhIcfF8Qh29GUqp9RLlNKLKdnC5UR1ApiNI85b+l++F5/BgsElq7gSD
+65xUFoblmZ3lgYDwtlYZNhP2kkeDvKS8Xar0wUn5QKFTkodwXFTy6czrHPuOFBI
em0AO6egpmPHtazIHfKI4NINbbLUKAvYmLlejjdByhcfWitvETQ7L1eLVSfG7uJn
D18I1jpLPJ7/tjord447P23IEuZmi/EL40QeaWS+XJiu2NdIELbDPRhfDilsiMFo
pOfpfJEfFGr2xd+3k0erdVPqirOaA1tMxjaDiG4o74+RkzR2y/h0+/WOQvNWQrPO
jj3jxGzWtUI/BCIQWrcNiDG5mL3/rtL/xvt6q5exx4O6dL9L6+w+lRMh5uY/6Feb
avUmUIG1GoK+64xagz4DlXnSZDOV0ibj1rb5ni3p/Dkli3Bx5J4diT5SciABIHNC
xPK2VyJnQUGSjnvTPvYlpn6rss9oldSzU5L+rSUmY+4+4NThg6PZsJPSR4C6xv6u
6D8gCP43jQ5CYjKDi5J2M47qfNpT5vPLXzN8UyqJ8xZqsurlt312pG3o99ZKYNwi
976xCSXca6RByIGpJrZ59+rp1vWoAH+vviKyBUK9sjYx7pe42HtA91NqnGfR1cL+
lvlRy4rJdKY0iYydLZ3TzA6E8dKNCYDIJwjS28Xr1gRCi0BEu6/EG033Tb8Czh6v
S/rE1AZtdHBPzCh4SERy0A==
`protect END_PROTECTED
