`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KdwsTRZOx25k/gE6CNC5SKOnZbMNAXzKGXTf/u5/MQrZmwVrvJtYYgg+adhDrA7t
V5BDW1vuKtSTnx5Xw1cnhPt4BcnzGFwRK0uoWsAyuBEDzB37/g22LGWUlKLijWCs
pgMI0nJh4lktgGhqgRe9kIj+zxMnrJhkqvriiRRAVYichtNSlLbIUPXu0MU0FmbF
b0AHdcKYWBNtUHNQGMnmGN7bjVRbnoVvujTTC6fFaRJkqAiyrKQ1Lnzt9UeASQF2
oxObiFbNteapTtYUFVlsOF2pVkLcCEiMSXI6qQgZKj0UdAt2hS7t+qUM6xh8Nbvj
mZg6kG/2tPeB6LPo3fXSD9lzGgRrNAu8qxWssc0owbUHQJGETdtSXQtKygyXurLw
eDj9Em97BFEImPfYD1ez6xLc1aZwD9jn2YDkbGWYdG2MKN+Zjox/+WP/2UG/TLNs
jdATi3ycvxJMC4ng8gBdJVGm9stM6/TEg7TIgdL5FGLPrxOkpMZ9Z+shphSPMcOA
od4iPIK4GO5Bm9qgg0oV/T6c4FyKL5CRZdy3dt+jarwUOA9Acs0vC9En9I3gH83D
8bilQ8pQhBvaLNsyzHkyUA==
`protect END_PROTECTED
