`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U4xwhdXbpVlE3+ww8/SPIBNVHEW+PztPGmZpypG2WIYf5/z9JSyDL163KwJL3Y5l
LemM5HL5u4TpbJlcW8LDVaB5BAgKQLkTA/c0iE9IxDtu1q6lQXJbiY+dUjjPtINh
tpkZMlREfzIZPrWoQvM9/p2SjSFnNHoVD2LLbbnHUT+wBfg0L4WJgeRf+UuzoRoe
mQM2Vc0rT+JWj/D7FIZxLvkkjkCo5WnYBRb6t+arrsH45JrdhILIXT5MBHfIm1q6
SI9nw0Imf1FZkiKYO9X7ygP3oprifMzVNGJ3AaBrtCNOL6k1GmSkYcTJFI+kEhdS
8tYl/9OdDylWGS7P43aW9R+YFJs9nUydNDakBU6aYOCAeiLR17QJOLn0ElLK23VI
eyCrJPLw4tdZvTtLiq3NbQ==
`protect END_PROTECTED
