`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AhJIL+2cfzypa8SUyi8Rg3xkdBSGAZx51M1kTbBC0PNP7+PmY7UveA8QSTxHKnUy
HchD9AT+FiXiSNuMZmd+LVUpYG8+WkSqMhvPo6EfxviKwOJPweIEh22RYFwWjuBG
tqV/ljPdaj6msZc7rha2prS5LLEhMADEl9E1DpExQxzekKpQiYdcJLCQKXgMiOEt
aA/2O15+d/nVXyK2QU9XlFwbMIp4WMlSfba79g+YvOOyefKoYVDY+kqZqomBo+NZ
p0aUDzzl2vEIDD+Ec+XnQ4FTig8eYhaWLO2HurMpCq7h72pnM+cqu90X/8LmJJlA
KSR2eaMFGJ8X/EJkGIPKf5Dw83Xxt+Ick+CzassF2Sc4MpMP/llPr4ki0KIKF+25
cReU2VSnSGV58vBX3dp4CSIY4qlK7BfzRLcSLfpSZnlPpR5a8WVE1tDi6th0jSnY
o1706bHMPdkcP2YFyigg4Q==
`protect END_PROTECTED
