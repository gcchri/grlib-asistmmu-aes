`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6hSXAeVzlxaF5772eUclLOhnWVU1cD2/oL2v2nsLWYFZd8xfn1ir6RbnvSy+A06E
aTWXgeBpwSc2wpXN9h/qw/V62K1M63O8Id+APnzGjg9rEuHKEp3cIwDiU/JMZtGq
swZyERhkVfRVtF8BIa/Hu5MDdCBzbGuHSmbGTfo90Qc/5Je1DDf34F/NAg1fJMNA
o3jY8LJkqgbWXi9y58R2NQ3qbc0cU/nG5Kyrs51oEKzub4IH3/og6TyeGLOXfa8o
/iGLYdpJ5MhjtvD0ylIzVOgfw+7eZ6/H/t21cTzWRxdxNj4hSuF2oETL74IQsshW
`protect END_PROTECTED
