`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qvAhAWZSEKO4tSaecF7vFE5xDKTrnghQxbC7QI4rRgs08wH4riRzsgPriDGkmlVm
vHJRm5oOLxFXBj8unLy73Xe63uSN2Vqv2EEEQaD5f8y3gJ/mOvOxFA6jzHZLTIic
2N7th855fukHJwVGlOhR2loX5uPS5bTnw7cyTudUKO90pTmHaxHSNXYperayK5VL
TlFHaC/A6GG8ScGddO1e/w7CbaJFFFcy02ga1F/JbDMiRcpRAYbHURrsy3kCbifS
0TTopQzWpOTZKuog76GO4oUk4+cHjtPsisiKOF4xBERoaJT6Awf6TeyMIp/0Yv8b
rX3Ldh9Qic8JLRsBvHsluSE7sZOlj+6XQ26zOYMEZHXLCCa2JP3zZJuLeujjy5el
1XBC/7hu2QtrWgPBQuJIWQ==
`protect END_PROTECTED
