`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zRUzUceFbYCVCBkk2sWmwcueWlua/iKwONnvTdg8vAa01FoTym8BECjFgZDSgxxK
TJQ0jlHW1TersQ9UIGvxj6LM0oh2NqDV8xN6bof5hj91fuOLc8q7TPm0ZGYZ9HSP
SJRJJywFFLomqXIloz+eZ+iaNM3L2CvagzWBKDxlXoB91FS5I6aHBS0P6RzpucLH
3/ZEvpsbe8K4XPyTFAI44jCQO75k8HLsgvkbyo6kuLwsaSBMxyNtXvKJFDYUV7Jb
5m1IneMOymTjejg3yFVG4pWx1PTIVG9LcCSfh5hQM7Zyw9jg4wVTmK6T+Ucxht3X
ounUNK5H+RyO2CklP4hQhRXs2EEJ2IEoc2XHbyfSoN5sYcqPqd1FX++gWqeBhLPv
L5ui/Tfv8uzZXUH0X3XndtDIZ1BbAxjvOTYR5wYTFCOCUJon53tHEg96zN3wu4VP
xXNrjphtOhdTL2x8cIwhz91rqORbvZEk9+Yaj4r7FGW1wRgXOD1Z7KoLA7ZxZS63
aVCkbfGFpYR2MhcIAqxDouJXVI0QqUnKFK14jCA5cOO3onhkZrPJ5UnXgegbvTR2
OXNDjBZGpP6yc91IkxFXuZmZu5tUQ2fKxk3yV8/Ohksi6xQl56YTJWG/Q1iQA7XJ
C0wk79DeH52DxAlliK/iZA==
`protect END_PROTECTED
