`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ItVlg3PmL596myzhBU1mKtjIP8EDU4qoOGIXZwt/SjI9no7eAsZtdmHdKeY9cJ2
O1JIYQ74agl2lZj6OLUK3SacG/onaQg3O1SYH5gH/dKFskT66bho7vBFuRSvUd8v
vvy5oeZX+wKy8mWTL21rzx8wIycKwLO0TGheiaYz5XPmWjliG3IlZUctheLiA46X
oMf4Lg3xHPKHLtT2RyIJk9plaGzpYlJnU4aPp1CcIvRABM/dO0cCeaTeT2ksg2Kf
9Wz/6BTyTSr3s1Xm+RF4oSy9DDlngNQzvZKyi9Hb+TS0tmcO5TGUuRlDKUY1HYXX
HlI8K6dSSs2on001m0NN0HqsrtiXAYU3Ncj2oYHsXQh9u0+GwZvSCgPVWns96PjD
jyG2gFPFEitcbV/htNlkBOElz0K7ZmufKTxn/Bcv7etE+7NS4kjV1nSVD9QxH7Ri
XWTvAA2ldG/5zWHIfq+qpsOcfw19nPOfdJEKXFxdfJC/7tXSngiDXO8AxdrEHMMx
s+mcPk4weRb4Nq/MiM4lviA6tBYr4UEcpcBAF59U8SKkmqmlV1tFy9FYOboB1DYo
OjvzuPL5F079AvfeUKS6KNzVPHHvadHtN9s6bjskCj5bgd01CNYYtezk87cG/9Dy
E7MhJyacklr/uHjisip0jKAAqmKYu+JoeYG/vlXvyLymgd9tdRO87rxq1m7ULs00
Q41oRZglsMBfMxNKWwWgQJkcxHLmLReTcf7p+w4iuYDPPHyvoh5pqWARap+xxX1U
yx0Gyyfd5Vit/9jM6cbKSCL0ePa1bWlA7Fg5PK7hzvCYKdGAuDAezTzNpQNlKfkU
sRYOgx+X5rgnwAURbj60c6BRuxbh8JbMcAUUG6daMPxnD52pbHzlSZvLtz/nqSH2
WuJYh9EZjOdtGqGLGw5MYIQN+0VTMWo6/Noh5mh3M1w=
`protect END_PROTECTED
