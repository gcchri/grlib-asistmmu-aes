`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f0+5h8uafaLHuO/Xmekxmx6/YKHsb4mdO0S+DxUZOIRxGrtYG8XAwY49yZM9KHXF
+GLTt2qYXbRPyMOBo55zJuaCmBsKkRulBeWryBqE9mUlqttHHon/BwGFFAoJ3Q+n
HR3PQVSCCZJgogvPbn33+8hsW1uWPN2fyKP2amg9bIpOAMNNqiZKE/CeCLuG1c/g
njkBRCJl87jVkj4VJ3z8S0aSpIjsZScyFIIp8KgMviMFbokX4Ef7SQKi02tE+wRE
f6GdpCNh66rUZ654EUL3hkc/y+RRD+/nCMxUoXiSb+ZFf+lt3COXkUxlgH05z2js
HcLNstIe5Ague7Yf7CXMJ+tQR4gTvZHbDkHN77v9tOZt+PcK9Da0dY9koFHXfB66
fytIPhB5HPyzl33czUeH/99LMV5W5K5iTPjYnfpkYzw=
`protect END_PROTECTED
