`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
phHnPGgUQAwKwuIlNCxfbMpga/pLrRICPhmK3GErkCvfnG2r0bmlSO7EMNMY/WSl
Le2dIJgUUDhU+1uPC4SMnr1NZ4eIMvvroOTZ/T7C8t4k8zAuF0XIEzDmvHalkqhH
cbkn8itgygrm/o//rCnxPAUQ5zir9IgwCdiuNw02oaPdmC4w4qwINPvCRLBDqjJi
Tt42u6ICqlEy2OYNMNWEInXkyFIgOgjCsGw2riI9MijrELhUZ/MuL2gUYJnkHReQ
s0jd8YlrG6Wx583/oFyfiqBbTG/oLgoyCaz3ke0NG8RcEerDLi+/xClgPysKv4yZ
o1IwhEFCd4B1HKCG/z9WlPDLdg8t9msmJDuRTgScbqT4qywoELBoQ3d/l1Q5aJat
zCepEjD0Yb87hlmErNZggqxdluV6YITVw29mkPPYdGLIGDYm8EzkemzhTawIXT4S
B0plfOjLKK5Tzp3xY+8LZV5kf/87fFE9awmXR1il8ElYI9QWmIsfjsBj0JaHBU1R
GrAV/9mlisHc0jXeNrGStJIPEyFuygeVALjBEIAl8otIvx1sHGEc0raWwVDZCNMx
3WUaJlyurP4pqwpRwSL1ixjdLBHtYSUfGXQUBWVDtax+HbEgzwkHDJgz+JyNnWvd
AvYq8i6vy7SuMViM1ahU77+oXX36B7tnydCxxBCoe/A+Ykqrr3UaIOmvnZxC6Njs
Iu/+HCKm/lPoXwuEyDYI90SZX8oPtK3gjrzj8JmNnv0ZvX+ugDZjnkJhnnlgCVzk
HF4gd2l6rm4GmZAcLxY2ir3PuzAzrK21VVNdhpk/qrEOn6bwdmfYJreHeeBAacnq
wMge2LL3Mxz2a+6VNspU0anPsvG/LPA5a4R/6l/bbeF1dRnpSw4V32TCGntWtne8
BWLYQe4RdaWhin5FIkymVBemwdQ6IbcMlf/B8u4D0cS5U7o+39znJxW4wg34gjOr
TivO3Wn/VebXuchkBJOHOxT5FGxaPkwqw6Axk7+JZJQg2AV2DqZa0xRjd8DBNecs
fP+6Z+e7HQQ0GpgzZXAjTvqNNFtq3uO8KmPY9arTXQhCuMmgcle3zwRrMAC9P78j
stU8eGt5Dbj/V53kN/YVkHYOBx6DR2bmVUUlHTlomz0qyar71g6Te9N5N5mS8GFD
o8rfHDv/tjPaE4QmVH8eu4XnCTh02ji22WGyxUsh8DbyndzTA9Dr31ZZUCF9H0MV
0FmlYveWD+pOXSKzRcClPE6ymw5g1PC0hyv2Rr3RDfFa0Z11runALRLzNXZEK4qC
aQvYanxygQJ8uauqQ5TxKVy5+72PSmiR4Qf9OX8Rs3/I65eqOjUnt6yG9xg6gRBn
sMkbhV6HQoc0mBlbQndikvctxdsBVaPL2SHRVb4jEPb568luSmlJp0ZnpJzqDxKq
ZgFp286jA/EcEMDZNYe2q9d9HKTIUZSa9cYIyCEWQbwmhlcXlTR0+CthDGmniqkO
ouwFEvi4U6VtNaAAK32fFrMAZ2o3kdU0Y1FwRxQ+fFIdbz4ird0yNCU5n2rS4UG7
7nLcWbhbbaFz7a+NAypcJtpxQbIyevxnEndJZrFDiuZ38eLvD6w1NHvAaajkB45u
oZrZoun0Hceer5HfDz6/t9UQ3oBd1BSW8HKiTx1NZwvpf19zjWFnMJhyDZHoWOOJ
XmpEdncJPxo4LNdVtl0DHQWmr3ildE8UhXHCJtf/na6hrbzey+1bzB+ne9keIuhQ
+n6SGF0jc1ej78EkyLrTUOwdTW6DPtqiNuSPrJN5oZgsIzghWB9GhGCUhVFxoNSQ
DyRXkztNIIeA4P3/Kt6VNmZzpZk5HnnHI/ChvF9L/fShHiua7DYAa2zJuIBTmHf3
GDMeqr2/rz70J2kBObkIm8lAeqHJ6EXXhs/LZohYyk8GLqbwBF1zNOgr6MxOAd+L
fT0j8RrE5spGkU7RXzAz4a81Zjnevlhmkpz0XH+CAxYuFq0WCw7U942MCeHvurl+
cs7n2pKqx6g537+gIqR0DmfhyJyTbbcJrCDgf1GJxPvYI07Tct35HnP4ld7hjx7x
qcvsDP5AvTzyPNj2FTiGWLZp6/vIwXXR298k7kaoA9I/bkl624ErxPh3q47RPt/N
MnFIa1FE92yF6XYRXZzRr9qiZSrxFk3AoyVEBhJ10b5q21foxk4jtQbIZ9C1Y79h
3fZlUUPFTSweeM+MTOVstSyzbzhWFu2d4PYrTdKXrhWblIgglWFGVcIlbxLtQMQO
cUT+NvfqDQ9xYC/2o3AMJKImQ0yI5X7aQJ4AcHqvfiQlCBbFi09k11uOpvApixLZ
bSFD5zb/3QvUN1k13cBOzBaRU4A25megPIdBcT84WqBUk0wEMmMSbY1r+6aDynNV
0bkK5241xPbQLSqQ8ttvVNymxMnVDBBjMZRW9ZQQWLO8m6ntyWtHqzMGuDdigAnL
oSUipvCNBDTicewtYBWYj0FQfVe4wrYy/RvDUaXSAzjRiL9SQCjhywT84Qbs/q7h
oeaG7A0fWvsp1f6A3AhaXUj5TDge25vLbeklfgwUUoxkch7fIRzBYurgNxEc0Z4x
Jr4M0fTUlbAZJAXesV+hera2GAgvRHYPiiYAIzHG6NzDjvm1pRgfHyzhyc3HiWHZ
hBp5af77sgwJgJOJiNcoMVI/C8Hlp5fUWomP6+Z1qY5+IibcG7z9V6ah721tM7wr
kiuErriqWnYJLDFnIcaT+lLYMyfjp8WI4pUYzq7S/kEd1UREyg6f3tcHrqEkvyNl
BQydrPfi7tkowuK9NrCJeHHgvkFfaoMHBWxT+UQCUmgpQ78cTrGKhf/g4ZZG7OCk
WhrI+Hov0tTFXq+A0nd2k0g9P+Zc6LLHLAa0DRfHdsGMRQrqHEzGRL/lJTo2WtM5
2Xz5tTU2EqZFR/VZ81n5cHHOa4vW9Ir39uRLVbbFup2aHBBSB226wY21xVAJ7rTS
dd++vfzxCmjevvIANNqu6dHRJZqpZZskoh6MLu71qvvLCsZoTICXj0l2nkhpxjkd
SfiS+94DmGH5VKCb9W5AXXMiBnWUB90gYJnqcmRMrermdmj1czj9UMPyLsP3Ifhj
zVQpnFkE5RPnsNPXeiHIWd6eU+TS3eQF19ryx66vVd6B0BePBZ3eU9zCyPr/W4DK
zX9pDXssTIQHvGd5AJJXT76XU999IAgPNaeDStNj7BxzEvE01pKyfAsod0QT1V6J
frP21ZMUnELBDC3KnuWjr7l3d/o/CLUUNK+5t6H9mxVYw7A0RoGYlRdmTlJzd45q
xiA2cGjHDxLXy5P40/fKXFrYl1355+ez9My7z28+pAvR55w4lQThFCTtLeHN3KQq
V4pAJ4PYAtSA172xikeI/Q==
`protect END_PROTECTED
