`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kfJCxh1B86fZErL6Y0z2Zk7t+1xdA7aD7ifv+GUPstPn51UGXP985YQqyqEEyDr9
k2CfqBmgebc+rTegqsI7nCrduKgqSFopz3M6RH32cWH5Ce8x/qunk9kAqzEMToIq
43ElQsmlzIaD+hHVzQPQi7ZXO0zfD/G8qL+FWd7jahhPh8epJ1h1kzEQaKK9UYs6
fzfgjamgS5GJPSlVZzfV12vGbdSjK0g2Nw+oVrm+/NJulOQKOpEhn+nxqE2/Qh7d
CgthOW8jRGvrwpA6G1ljkTienH6izbDNtfY+ju7XL/3UICJa333wB3yPmZ8JxXiV
VT10jA6ieOM53x9yLbp41FBVU84b9gK4jo0sxg7N30rkNZinHrHfT9mnSfB4kaeL
8baWWgw6Q7SCsFi21bldJAxEywpHmNlBS55aq4pFrqtA1b60h0iyfb5Q/NJgrwV5
z8NDSv2hFaPmCXB7KkFLVs95qT6PXcYvNMb3dzlm55nG6+6+L6llLhZT6y+ljF1Y
qZFcyQmR+FD37upsJ3jtIysTv3yxSDqD6zFPq1JlhR4J5YZBaqOnj3TZDAfMHJuH
NkkbOLUdwOyDKPblt02JFfUK5qjN433m6W3KPYZO4lkzBGehM8trmHGQwGWnu/8Y
yKjCzbp+NMkP5/PKdkklFmaH/OGH5586D8SLUdQInMgDw/khlIzCOt8Te140tc9v
`protect END_PROTECTED
