`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UYaC6lJnMopJfkULCNxG7yTfJw+03A/uryGOk3vIe736sjiAax5S/plVbhuxw7qA
4ie5lZjCSEhXCxbx8lrnd4WEcQEYjJ7d8r1lbWrQnwvsJM1rSBW9rWy6unmiU6jC
8ECraBVT3QPq3WH4m0BJtBOy0R//XOvhYAGpAG+gzX594U56D0V67dzrxVV/fe+J
U2l0xhA7VNcXOTl3PAl6qO1AIFDSTGy10qoryGsy5+lX2JTjgWluhqetM/txBs5p
1Mtw2GKPUDP8wR+td+GqhrwhpLX+kq/MbT8tDAQdZ9IS37fmJGsp1HkAX/KAn1KH
U/AzNa8zFEh3kS2H2w3nvQ==
`protect END_PROTECTED
