`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xPOM+yjyUid48Dg76rtXl9t6+kOAORDka/WzFhn0yVNaShDPQDGa/ta2DnP0LPYR
qniADQHAlqXhQi+KrVVYLzmJf+Fbg/FNKa0Yt2w7AT0TXW5NC0IPTc7enbjapZn3
lqvqGrj12AVw6tW+xY13no+79MZwLHCzpTgoWVuhGV4r02VhrALcnBxavrSgWMKw
RMw3lCiozLwGkBsHOmT0PZ3TQ9bIS1Z8JCEotfbt9tsVVgtrHJLGWQgR3RRLX/Az
lbAWVg/1MLOaLZFSU6RvRwZ955flpQTLeuc9MbAtgu20dG4dBAkvWk9lgTldMaYW
C52E/+IctGmaV+wS04nOErdSsJ6BKhgVoVBl84JP1sZ2N8qChtcQOJZtUpnJUK5x
KRFct5qPy81LJTV9CJc8+0/fo+KDnMkhNRjFqnkD3aVGjJyPOwwOHCE2iPzxKUgh
wWEhMYahYTQJqpvJsgshjPMTYwRAkgmeXYpj4DgIpQNgXEDF0/cT1JgyFBHSRqof
zQx5CrF52U0zMlbacIpVT2/61dARRs+Tl8GH1+huesMFX8uQQriLxmlHOkjXii8B
Y3FLSNPhzR/Y42vJJiARkfL4/FTXSWYSM/mGS5FGDOBivrn8Hz1KHSGhPNx2OTfK
NVf40V8y8VOo2q53MODKlOObAA4s3R7YQfpCGBuW9wP1kG7EkcfqoWlRUGpL0kRi
ThC6z9ig5XIGamFVmg0q5lw3kH4YlDGRYVyET0BL796ktugCy2xuUjLDtHhA/WSP
cP9CUclscSEW8EE6UnCBSOvPHmw1DoawjxuEyp5a64uvfX9vX2KuOH8z8WvkUnji
D+RNKibPIKnkRUKF3k3367KW6nCvovxeWtuX0OxzO6Xzz0pD7fTEPnvnTZ8sbwmB
Kb8NZRJ94TThRVOS5iWTxrDCAO+G82kY82pzV2PaoYwQ+qAPcQxGsBRnGuuJ/5XS
wKvnFQOMaCOiKI0T4YZ2RhgxLHq/UlT+dsDVAjQpFZg0uh4hqMUP/Bv+FVNF5wHf
UGyWxn/rvcCq886oZpRA1c0cjNcxcHjxby1PPYx20hsr+ulfUovovsFw+Ho0d0dZ
08SJKHIp6i6CooPJuhWR/y2jq3piMvZSwbFwBFX31ckx8P3n6AhVGf1xjlFMKgx9
g1eakJAsLnd9ENN4Ye3Rafbr/NOXJKfJ9Hhth4oxrjfmqdgFGwnjBRS2JGEw2EWn
3U2dxUvlwCLiZMFY4pMJyqyH21FCMW14wcQ00q2+dIalA9f+Y8HWJkWgaeLeGhNP
DazcxdUuzi39SsyCKBsbvUsGRfpOj6cC39f2ZPC/ogU+DorpKAzffl3+FBXYEfng
uJ29Cn4VhdHUMIxY4cCTTSJNE4hfG36QUXDrFMxGQsWg4p7gsRCYQA88a3lOCeNd
4y4QAYv5bRS79vjJDtVD0uSNEKJX0ZXeegvjhy8feg3CyuL56hUs6xJlB3km7uXX
8qqY4vBUBftTdVaO+OJGgyuVzEKUtqoDa7P6G8TOyvICDWKP71CGHZSLWayXQ1RV
LlUv4rPtZvj5kGFjIAclEizeGWOddsnPftP2yN5L5uiRiDw15ZY6ZoaHElw6R4CX
FK4aDq1XtUq9Bhb4HoVtuBE7OGlaqU7COQ2kfQZ7i1Ax2lNB6a8UpTeTVhDLu/9B
SSOqt5a34Tay25Y6nFEGrh0h6ql/Pi+8BCY6TxiJ540wJs575yJcTkULVNPJJCoM
kS8dsCJVjd7nv0PHOezyaEUVVaYmjRfJs5Hi/J4np+Ig/BZbTOldRODLOTb/CbXX
NaUnBi0YaFcXvTAWOnRtthNBmF+NVo4c0s82op2jRm0DRcuLsvIg7B2KEATTOzar
gxOJvy/3Voby3w7GCmp4GQ2zM2nBzPcUVH1X62LypdnJsPOAAKYrpdJWf5wnlsFS
d/DDfXFOwnKSiQ1+AYDtHoD1+p7Wgfv2DxP5utZl/MvypYBn/BMe9fOL1EAH1OMD
djOCrFZdXp7lr8KuOGLyIV291rgu0uX2ce47mRkm3nmaR4+WZcvgZVwS0PbvXday
CHxBSgAlJtbcEfwNyFILuCjY3AWhdg1dN0Cll33f06rJjLdZHHIPZjBujHjBF3sG
SLIjXLKBptexIvsJJ8j/RrlIULRpdw8T3+9/QWGa81B3Tmq/3W53tL8Y9fkNbPTd
R5sTmaMcDmF1myN56hkX6gL3y98ZDeZZkwHu866PuWNVqH1/OE+xILhQsji69KXZ
PSoL1d0h/5wYQycsJHL8EiULhaKg1uilJTevnvdTat5XcVQjM5tQv/xeZSRYaeuQ
uMhiusOurvFHWzAitDREE5ImIR01rpk0EOeKt7Z0OYAS3X3j3+P3deiFdTSVy/ux
Da8l9M9vg8tiBjf5GdpYoOlN4tB0Os6cIiia+j9LWWwF6jTuOhFPgXjWuoXCH8rQ
bGiVApNOgu5DzZobPLN82D6s4v2/RZOrhV1Uq7FD76uCWKIVrQC8y/yZI4KlGCEM
Mmm8g5Ya2HnfkK18EIhorJABRTZQPbqR+QyyLpg3CiTRYhGGkVb9o/xJGyIcb400
gqqRrFel2E8C+uhpikT6c1nnDt0PqP7ZDTRKMKco8Rccr+3oSUvNLHSAsagTqAMB
8fFTrXu64kFSEl/z/zJs1h1jqM+Ar588SNFx8Dg6mduF2eFtrH2c7ZAR7FzvyVT2
1L5z4vtrP1MbBlMZ0Az7Ctr9/pd5knk3UPPt58MwtKXDZdHykIf7JRJ2B58FZIMU
DEzr1TUOn5dASVQI7SSzuejuT/CzygrTzuN6ImGzzPM4TkotCBpmhpQ8Xu6zvB7L
Qaro/fY9X8tkyciH+LhEt4gA/WWIVRMjmHizpjemjSuq6ktUqAfYhtuVP2DRsegN
Y0lxNahuviD3ucYVfbL7FYFpZ/Hzwj7DQoFo36V6cJ9mxhv0Df0xtE3drgkXqhZI
cm4UUmUAdWKqwo3TRZaolfmhNNE4jrSws4DIH7feBmSex8yWja2aQ5vhzIEFsz2l
H7lhXNO+CJAQ/4CQ9cXi+LfI+7DM/4Qv7oCEzblJzhU8nwbfdFyBq1k9vZRN+qx3
U5S2KcXZ/4xyf11u/acy8hFMja9sG5GNSILyoHRGTWU9DnLNGombXF/kS2Hku5b/
4z3BxHPyOfZQOasRIw3DFqi5k0p1oYix6mm6Bl84H38lAlDXgk0he61ycS0eBxBv
MmOn7AAfoS1+v8vP3xCD+j7KPAvFlTenAEeFNXELOE6OUqqz6fD0ii+ikZP62Ezf
rxy36K1P6IEu1/hFYJnOlVnfEGMWM1QbhIQKRdrTm97L7nwzBB7N+ZsJ4eMzkuZ5
7Z99UG8ED8+/Mse6PTIZQYKvWAk4mOZ1un+W+wDkiEOs+m4ffBnLGdOB5TLvla2s
lO2jcnw/CmGVERk7b5D9z/6bM0/IsRg87TjMuiQVIYg7uay4N8HZIbdkVa0sO0ZH
YGpfU1KZF8n8nb0QiaPULeyPEMnmGNnwb/v8VWPPGWtxI8w6TS+5vDjHX7dlaZUI
OAXrxzMDyyBDfhqrKLUtpj48geSqDsdCzaEgwNMGrWs5ym72sPBasqJTD3QTewOj
6lK4uJuVKxVNRH4RTIw2a9KhR7yVSraosxJhswLjVhAUfVCRndDwSbk9FowVA8R3
rau1p69V1uctfCDAYCYPVZWgXLwyQrE8Oe2OYmX0L5ovkn+0fqn+N/0YHB0TzmLq
2r5X7ND7YJD0kZKBzb6CY26gWsvXINTZjYJoNfXQe1Pc7kIngTMGcM3tRlXf0eWK
UiCIImRXq3RnkiDIg4ULL2ZmlWZSa+SrVgFEBmG35XyVIrH1MAGVEaETN+88Op3Y
upzQOMZPL1qzzH1ziKgbaQGy/Y96ap7ihWWNi35vxLbJg0NraV7RPRVS4sSpWtmV
+Bj2drBMpBCVrIKVTQD+wyxV4LRizOzLE8LBJ9uXgOcAOG4/WFeMmL8j8lwk4hX1
mab81jjYBIxRqaQAbTloSYoBdCxJjMO+T/DF0t6K8fgJkT1+jxnsnDLFZIrFecJg
HIJENfuPCdaG3BB/54xHXGoOjQuf4z8qS7fVJze5mEST1Xgx4gnTqaqa0rRH1Cuj
W13H/ahRSoRSskHXgVhQLxszTQSecB+3/hnLygFt7VSO7C878uBT0pj2PK5wvGGW
46QstewNZJ4lOABZpJxBchFPf6g0fZvCnCXuFRpnHlV/v4XUoUAVG375ZCgZ6+k9
SZ7qvSmJk7htCFeXpa5KaZ3gKPvOMKEN+QcC4QPoBBROQ0FCWVcJNwEnC6Ke8aua
fxeWb+VJcEETGW8Ih+7DVuapHUS5cnVbjGcjDKIjp+C6Z3jizkv3ZVr+x0EF6vyt
H6CS7gqLRc945ETFBOI9e0Djd87mgdJuuiwv+iYcsSMUewkL0dJ5NtClXhHc3NSP
52EZLjJp5W1Z2PhwWn3wLHbFq9roYRhUTcK4j4qNXsV/IHS+Xiy0/E48+YFpoNmv
8NuA6cEYFMtYUoP3zr+bk0gD/0+DeQcI6qinY7tm+lRSgM1VHZNP+sKyJnktMASw
SDKbZrIbnwMgulXuLW4PPXLOhHcBJ+sw853cGIrLA8n2z4xpau5gtSKL0jM1IODf
q+V5RnToILQSwr2KD0Vn/qjIo53sNT3xO6+ykczi6kEPWZpwR4ey76e1rfbTonJK
OOoCycLgukNIVTxfIJB0wBFeI6F94LumC0q0nLm0zw/l+kzeb1IE4XO/iCdXITLy
RFhy4nwL7KSnwgLRIMsM/vBbU4eM0F4xhS49vYJUxqgYsx9Vv3wSs34X7RtOO45Q
oq/R9ZPCLRtLN0Uw5gtByPh9gmYyUGEgumaAfSd4xUVu/6u2yuqwchKh3fuCP0cE
IyKG9JYRw1CzzrKy/GPzgZ+JIlfdBAZv+nHvsptI7bb/YHoFhKeyjXqSniMOEFQD
fnd/ewzDYUAHSUdd/X79RQFK+jEA/VIkb292uNnik/x25UfILYiVTrU/T4kht1kO
Mlc8hJxqWejgIclk+x7IuEeD7/N5xnxu1xtDxNP+F7Wsbo42koeRTyMhjOLZaGf+
sOodMjwBiiZuGQaQCKsnvfwqBgIqkyJpoPQ+DEWAAMD6KBR/jnnxxUjNPzYiHraA
IHD0UvIVPg+WULlGY92PN88tktm9qJLn8s8O7tKuSU+uj+j0O9PRkTM+xpEZrg+r
AcG3GjDB46oUhXhEQByUpTRpwgHjEmNJ8PoYr0SbeFR4YPT1a02oN0YbRnrzIioR
czz3+cc9kSJEpOQoUn2ehNkIfVJbM+u7Rz4ZHKAMcyNIULMSHGov8RhU4P634scT
AhXw0AnXiv/fe3EpY2s8bjFzx81c+c8viacJEJWYn0eqTbZujunFSttgOFHjoPqE
DfPGedwx+5K46TTVhZkiY4lTI9JylSSuDUT9epclNCRx6eEuAsdj4aDgOvnI0kzN
wDayocQOWSVMneAbStyeR/OBD90qw/OqFVj8Ot1uvHr+EvwwnhsT1We6y6tw1RXz
brk4hZkmfyUaf3YM8kBkuboAEXWMjgBZTYUqJMIxLfpSlXGzjPEpSG+sLdeSuO2D
BIqavasIJMw+P2kdEXU/bTYL5zNc3VoWigpBjY+2qrAtoxO3vAbiCfCldl9964tC
9yaDUZqoFyIeu4qi4Y70bVI1HUFm1r/ER/4RTuwIRYN5NZaGRzPy02xGzuyGBnoJ
3F3/QFrZCZwUWjYnqCoch6bSPnf/pbJpBhNP6rJj4ZRbKq47ihOer35AohXllf85
k7WnOYRHOy6A74+nAEjjgkOyEnu5wuTUTXcWppW/ifP54g3iVQQxKym3YrGi7yWb
43ajQiCM+bqXGLZSKg/IMvUx1Mqq0JLYqsBPTzxRnaVpyiLaIjJieyl/32uhDxzT
/XCjOUAYSc/fuNt9R0endkDvVJnusZdPHpiPrrz5SvYAP5r9KvxfT0VHiEUE2VSm
ddrlNtQUm+POql5uVUwgzN4tw6s4XKsJKkm/VPYQh6RwnIkM3wDZzFHVQmPf6xVf
wYpeL98LOPth6LSp5/tghMDqpo5WCU0cvJKfSGU6V5wp7ECO6+uy5FSuzsYGs2Kp
krBrMw+NLjkeEjXIYw/MUekr5UYaFchhupDkphewMY4xZ6byNUY6CLvlDjLjup8G
n76HnsFyfmOqw9bP60NPZbc9uMmTtCQ2Hn9D8I2xK/3BuMiS89fZcNOX4weSqWxE
fZwaFL8bQDqsw8IW/2zbjIP3uIqnpMGK6RnL48fhLdF5TneZaX1VUY54wTxN0Ckt
pwWEP1ebya45QUcMATyTavosRY/2dDH6SXRBarJn0CFrjnYt7gGkflJB1wLumv75
OIxlEBCbbn/7csGjQ0UgvW9a0177Rszo5Mf7jmdIxQB9JzuJBxyz+YlXUGCdiN/g
Bw0lP5tz4HZHT2oDb2LOUME+A71uqqBRVfSZQfb7eNstWuXk9CPRxj4Kkp4wkrHM
6NOX4rNNZW+plqSaR7dnon/grUIQqw3IR1oohyTh7Ud4reDmFerlbYLwhdmpKtCl
oQSS4ehmZTNetzDrNkZQCuGTGcMYFMUnxI9ORmEuyO2cTB1Gi0MGM79UF0k1Kh3b
WoZ1OC7tMIWx+ePfWcYN/1diFhmke+12mK6OjKEHJwpfTtIHTBo/mA4R2OMZy9Dn
cT90pUWYa9rCvFz33+e+1zYh1qlw/PAGK5fB+xpOWV7XO1fSvLOueoWDuOjHhqpH
WcMtar+gGUbD84UsxJWJNxdn6ghVF6tonA4aPyO4MsIvlcNSZEFXd1U6+if0BhYg
kLwJ2be+GjHv6Q7p/SxcR7RR+GkIswdG1xRv4oHSP2BlnYNiFwMO4Ihe1eAfDq8C
gbI5srD01Y7jYAPUvoHUneJ+g65rCkVF8sYItx0ILE/SFJK88nwvWUazx2M7g38I
pLF98IfA1uT1IlzY6eRFWq0MtKXaecnQ1EsAtxWiFNkd0g+Yu4NEBsuHPS8zD+MG
/XH4MWgMb3B8UXzTgfe6zldEM3n3BxKZXMrWskk5exAvc9X84De2o0Aqz5TzOtdj
VAgqjwfk61n6WfydvL+jgsyhqieJtYUdqBrYLxCxsBDKnGCFsyMLHHLrg0jdqK1W
EcYdNU9MpN3dhYvrsAqrfDNHMNRg5v9iVtCiY1w2W6/kUSA3gopQPUvVimFYA0Xp
oxNrWK8ZmLK2yt+xr+Z4y5RkdexNtPycKWZ2Ak6pNzWGIN5Gis58RTOMJEgX7mMy
T/Lqe0dtdhkPArn1ptNx3MGa5A5S46LVNuhxIvpVb5vHtNq2DHHym7eA4Lfasph3
CcDJuSTtNi8D+ZrMr1Uh4XkrLGaOBMfRpAHP16+3icxQZr9D9+aPueCx29QCiPkh
TKZbBXJ2C1lcz7Tuol7rUJBjwzGK8aj8hayVXizw/dR5zt9PMIYs0EGEf0zA7CO6
ETvWebcAtCH0BixvdzysXpyC6on+0xuzN3sMNjBrfcrEQGQe7uX/GKpFI0ExYGhG
t4UTz3AqXL6QtMJJmsqP5EUSVwji/mgC4eYn8EkkiK4z0qQ4/0cacUpx/KVa7BIL
TSSJbzx0xW4wzBeJehRdzwPusZg/7uLg+mdsh4hWf2qSRtgdfOUrGeZKjn9FGDwC
Yr/r36A7kd6wKKS8OJtn28UBZHr69ae+r62OEHFGVCD/yrhpbPE2JPMrjLom+IQf
iV1+xQDJlvqacEJeMVem97K7QKeiJ/mWd521GieNRBbPPDJIADhSEsm8Qi3eLq0i
MK0sMT9kkmA47QdPxvRFN6t3sqwOpcFc1e1EWAjtU68m+bMqKflGoJON7DgGAmJ/
beScJiJ1z2lUhOUd1KuK7oR75NXanNMdLWWSOIVTTUbBSKuFTNgk8gemBSUvP6Za
FnGaHxD4Tp1cjshE2kwIX9Bj4yl2+Dz6otcLDbTVuXz+3WISReATTFGCcM8Y7rJm
+//0MmRBu7BMaBFzvz4i3JaBSAjN1bNDIQgTuROqfYYMmpud4MRFLHLknY2RLfJD
VUDfSdAhFm7mq0GC0a0t8GiTtpcEJF0iLfrfS10kYDDFNqjCGWQrXOLBhfHevp8v
IWB/ynCK959gkURah7XLV6hP2k2EdvHwblFZ6f3KtMFKKMmV6arwdXqd8PbTWmab
yxKI//O4TS3LfSthys+H748D/T4V51YlctO39lNWIQGr3KKAPVccywWcbkZxKRXG
9BLLP95+2cadJtbSxTYUAgCuXp79wM9/dmJOq+eZhi7GDrymfE2cD2kEB4PQRLSd
VXXBEXT2sUabhEoMcvRjjEwLlNR1Avqsz77HuPx8oJ1NJLQc9/N6Mag40ppA35H/
JGsmv+/TJcCVn2mv3g/V/jTep+CCwRD1MCSUnuwJPtCiavsd+bWLXKMiT2XyE02i
pgbvno7YFpSAWby778GR1xIbMxav/r9WSmhLG/RSnRMILpgbw5xINNbpS9OsOBgD
fBIfK+RqZ0t6lt1qqK/tAzhLll2Qq/wIkY6V7exWwRVJQNTIfYjg5krcioNPCVcl
5fCkVhoB4L3d5nEL3FXNEtm0ZwOJMlXpD0I4kCnyJWzASy2VqTu+tfWFISbxTQts
/F1qJbZutcgcjJNvL7WTV1xFvFJaePoSi96kLre5NYSnmZBfen2POT/qIxAJpBpv
Cs1n9fuZ809Ez/SCCorvEQjAwlaZHLeRqzjYFX2xY3+1dpgXMyd/URoOpGuvAlWV
WT82rAswIlwkF7JntFvmR8grp5VubcJYK5nAb+cHtPgPyXk6zvP8+Ovor4PdOAP/
6rbkvauYV8HyikMT4K+C9AKybBRswcPsyDFDUgueJknSCAB7kQSCMO5Ktd40oJ/+
Bm0tQbdB0MNjxJ/A89tHmfgs2FIbqNl9hxnZqlxtmX1OlEpQJXF+o3TwyQOYIcJ/
1rJFAk9aMC6uvUYOXglacDYd2Ybf6SJD/TEtA08Fx+qS4b205qTLaG0tQg03E98K
bDue4/b2SXXVuOnQyyWrd6V58CQe3zgZ5VkrPl35X1jo3zuGe8B0chQskfPKXgFv
kcrwtMnT655FZbD/S4Qmx13bIcugYK9M+5GOB74MERfzo7gc0MVNwzjfo8CzGRya
yI86Txxx2UjaSkknxNOpXLg4WF0zHk0aHSm7W74zhwE28CDwOCxXBobhlk3vUB1/
vmyH2q/7lhhTDJ1s15tSg22QRBWF6IFv94e42kd5nVWtt8dQfoYP0n36FI1F7Kdf
dq9HB2q73Cpq6E/TYWEzPcmSLq6jovAHVYnZSLlAAmqLeiutnig0n2VXsDjzxDCR
briXHgn+G/MHTWeEI6mEsfvA/cSgG3NL7Ji8/RBHFDAyerUKkQDFdQjpk2fkq61g
zZaUXqQ4pJtYAb9SVeIobSl5uqHb0fD1PlDU7AydOSwSDdU5MUfkhK3aYqcecgOX
CYhSNlFskk6U0sGSVWyKvWJAuQCwRDOSOBDpc4Hq966iGWW59I4YkqaaC81sbSR8
gcNpsmcpPf4sCiVuIuwHXgAMGIeaAAFb824aOaDuZns=
`protect END_PROTECTED
