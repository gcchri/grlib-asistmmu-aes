`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+jq6o8MrESUYtt//PCmVOWeO/f605gMUu0AJ328xu71qp/QnpMPlzU1jbAHOZbgj
g3CDmAskynDr/Jg90WAQ8XdjCexlADU9YOWpqRRF4sD/mYVXPaBFWJi3rohgl/e7
8Pg5iE4hpXW+ORJ3OsDRP/taka35c9kp1ZSVc2AXKmWJryoxkEt6AmceUl3/mZWb
v0xtBwpMvR9Tnn2rgaNxbbkULhnrSriR8bc/99Qy6kM4YeO+T1KrOsoXNCX2WtU6
HY9baDXuv7U7wnNJPCdwVdm4XeWkRZqqMB7lUUX7j0LCNbXAIHKr7Urh0CJE3+Ca
OGgKcKdGAxiiXIfikFOyg6pl7GX1B1He8opbfSyQ7urClYd2p66EzJDSf6IyGIqU
L5SToC4AkubTnyOR6RBcaYu/FFddb1/uvbFHyWeeUn7j2vIgKmTwacRi9X10Wdlv
Ip3kFegmRQ577oI9mVcTczqn291yphvPPcOl5rGPjePStQjbC8X44sCdDvfC117V
DnHuraKCeZKYJBC4y4UR0BCngmm8WFv2vzyElCQGWibGn+ZD8HGZSFsydsbFzZp4
p0jyRoYfH9n6hRtVn0S7u+HK5oP3RoCR4MraAh97V+5vtx6xEoYlyLXWyyUzv5Sj
abzcjqPhqjLSIFFSm4vdeDVJE9G1QND5g/S+AuEa49c=
`protect END_PROTECTED
