`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AB7uM/nftlJ4q1l1SCx71GanHefVSttemV52Ut4LFkM5DPAdhPnbCL222/3mr7Bf
gUr/3FIfweXN6G8HQMwnOKDP0O6IhQasa1MgmqzHF55vavOHp4Do33qs12it7SR2
egJmL3M6ZwlBA6EIYl1KIlP8oESJB6HiLl7SVTmTLBJK4rT+K5bgI/oAM9gm8PJz
djb9pZqq2BcF0+KdMfDS7mpjq1Y6wqiqnJeU2s2yi3ijmuUhZKrdMgIexYzVscip
FC26pW2Ecb67v1Qw+Ewq3g==
`protect END_PROTECTED
