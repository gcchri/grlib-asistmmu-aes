`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BugBS1Qb7Amrc8WAKqJuI8VYOHzNByFAq2mZc7lHtNLplanJThs1LVtE9W2Asjea
630WNtGEkpO84z7nF/BmXyNm5DfRIC7t/49QNcsbN4HamFNT2bQdV8APie1W3/PS
28lsm63YiHGiG8JJCVB55iHzlxbAyNE18Naa4PkGa1Tcp2KrkSvuGXU01oBXauOc
WZiYorb3fkKA+ktuxrTpwtCwLMsNk3JzHhpiYeFU7f3T5FlJaxmUxgsYJNWDvGHy
aClBoIJoARK80N7+Eea57zlzuxOSerRLgcneDhPme1eojiiPjy2KXe80P3Pmt+Sa
+qYsG1jLNH745M9FFwkqWXxkPqY1PnQXJGRB8zaVDfLwfdknTvMoSTP1xofb/HuP
ZwJgsmquqkvRwjzbhvJXWAiujbKcx3QedIUoy6B4BChtH8T+ARclQhYptSChxP6j
JZXB2xSYa+TwBZ9BRrUE9JbM8i1e5sQ+jBItQlMT2+99wIFfe2AkNcyzy1PJatKT
IfyNX7h2WDB0ch5Jyu78inSK8mtOwoA0OZRH5SAVohxTfg6o2DmE6deUOMAeIR8d
PO8mh6pgaO3hgYYHPQTdLHnn0wuaO68nPWmLM70bAeuEICcLDb7s6m2n2rDgPpYb
lDnXar1X6sCUM/mMjSqKEqJCNQgzK9wfQxNuiT7MDn0/3l1SZesOi5XRSszldxvM
rfAJ2ASrzGYrIL9l+6c/2iVFvocmB+6S7luW0Gbs0uqwZF6FcrdaEpuMyNF/nMkl
pxgoSGweGB6PY06bZrMhzHCeC3p5diwY2onZSTy6/XgX3rRugMxA6r5k/x4RpdGd
IKxKBeDfjUmBNSZkh6qk3SH1zSqVVhHapUTwL9Lz1Bf8gC7UTn4KZbX1hi6xpVPA
6jgXBA/9iSeNbmtuYbUA8v4tKg6O4HWq7ilMYfSC96busRpmmzcvrwKNOKT/Aw1E
KgjnJisaS7ehoSFqx2cofFp5fg/UCivs/zQLVLlmI/+NzPt/IzMSNrB4nGlBvIHg
pNSvZU7vBWtKDLP3WqgvJTWiHa1UJPv2YJJEutjr1fdUqiMphh37zF153pCWu/LD
ofjdJ/jacjblKIIN4J1n6/Zn93l2qkwsAInA+VBlqUQyszJdMK63fx5tuRKhHq46
W8Z/mVqgq4bKle4G1Q78fu6ejE2lUfH43iB5mIRFJhS92Iz8NlAMLPdAzNU8zWIs
q3fB86uZTa+d5Eh+p7J0s0GWeua6pHUFBrz5NIpneLHSJp4K0X4M8mJ5keYjuiyu
RY4P180cFPqDte4af5aXoqSCtybmzM7t9bCRzI/MLd+i/lG/uttaW784hXLSt/zV
RlFSng1H4NX4z/JaEaSaEv3GQAS1pJX2HOpCgBr9xu4m0A5qWXMGiiOjZBPO7irk
GdkQ8BMkCT3a91L16K1Iz3WK+srTXRySr5gaPHFl2PxbE8H4IIK6GWyKMPnOfMsE
m5vnwmWGtU/xxy2wgELGhr5pNpuVLLP/5KZsIf2U4Q13g/xQU6q/he4MQSCNlzUc
2u5fPr+mNi5gj6DgLGZOAAGg4yDOYDbvTZEw0Wmzn29ceKbQfb0ufe20fYODqO8D
cu3Rl/ynXhEXAVk89iWpzfp5aRqC+xQ5mPKgTwRbhqfJ7dqE1+/ADDnvneRfvmIU
jsQlyJMvB3dSz+gv/MJM51jTDoQ3MlJgxuczmdouIg4zQtXwPBQVlKCTlKgQt9P/
ElKY/1UCkCXrQZ6rwPi68haHdGw5Jjm9vOLI/s974l6XNJdtJ/r2RBAmE41Vv7Tn
TgSiUhbfaPPeW0tqtBO2vC5SPLaOCpvyixP85AyfcWf1MJqJazVRlEu61c1gPytK
OpK+dHMRlStiFwI27yXneOtFeJ7be1LAuDmxLX+LSboGtuyrFKgakHSj1hlHTWwe
kMr+W1QpP39sA3oruKWnLQbpHQlje/kSWBjhbpnfyCMvnHx4HWSR+b4g6USbW3vK
avTodFNLvXEQj672yHyX6TO9Nd8bzBf0j8E5aKyUn3VUbjbvZ02wD8proodOqWED
o6ktxMT/yhCzJRClMw1wt3eHeiPhYERId2g3tMxrpOi8x3Q77Mtgco4P1v5UJZ3q
Ua5OITsdMNQmDasUTtuBKq3tz6pFRCDvILzPJyOf4uECZZ6tbNliSs2YZm1i5g2D
KSH0X6KKc2a58QXNvBHNU0vjh8Cpg/lc6IA6pYRhmycMxbK4jqJA/y/3J2NBpSzq
Y9qhLf0qSPhXWyKGlXWPbrX0bvuarHSpfrx7t6gz2ACpzRL+ocZpqJ4oAFABrI7v
8fjIFiQPgg3drdcSv8r0qacvy4FA7iP2gs45qJP3PAEbwj7zY7MHJ0fF97sHdfqP
Ad7+f4x5DPKS/peZgHWRw8m9vIj4Zt/5C5qCgqGMUQfKEv1xien/qxbgbBBpyqDJ
HX1gnSOKvr7apbOn0d6Y3lsDPXfJ3l0GP4FG4PqKQg3lWyNNN7zouLlwI61tY3QX
tU5guS1PIj6Il1C9w0kdmA0mkq4lK6vVg8LBnvH7DJteTgC6UjbRekP46dTZfcQ5
D9Kp+8JyZvvwZJscm5K46lGE3CAsKOUjr0b9FS6D3V8Th5lS7UG/mipHjSkkGq64
YF8cpsmcxePTL/zEks+Bsi1bqQTAa0tdICM4m3uASj7HJhWtSK+hbDb9Iont3SiV
8S8LtMKOxw6dUp9pWbYlL41UQAULq2DQWXJUB8p/0/Enr6eZ3JpwiIr/tWdxvSCr
E9sB6U4j7FmwRLwxiJvMBKc6fXztCxPzGDwjVdPnpE3WZiIR+CZpsd5F7+5qjyTY
knH8NhL8xGjU4W3Id6/EYhr6TfRruD7dNdy52piL5rrXhacjyJN4dVCVY3b5w0oc
ogNpad780YnLFXSGov4nIegVIhZa1d+3MOwmRMYUd5i3AZUN1Uhauyvt6BKfug9w
XFegLcVCoNJTE/OS9FuEcNJCCTfMLQaCTV7pvC/2AbepuCsmJ9TfGYY+mZjVbMy6
NIdT1vxYpkXbV4CR8Ujuj4cw0c/3YN9BdxrlNvcC8sY4xtD/hvcgYM5P1lQ07QR9
isDLjDc0mApd0HGHZapgxvLC5Gv8JnxKaM26+YZf6bwgFbgmd67KnWz3r8uSXIWS
EkYEaNEizANwnfVjGGbEnTMaPKfi+d6tR9avTdbvG+HtAdiEw812gS1TjqXFxNjC
sgKhNOScdqAi7/RSpxQk5D7KUpldxbv/JhewUAZr+XsjzXu4UBXXUzwRKAztQkVi
9xcxiRXHWFlgbNrOdJJ6/mbgog+fseJUdUZyWq7o3IftdtqlU43xice8EJeMjt5K
c4xrmcHGkkJsBFK6eDQcZ4FkxAYzgu6vMDDlLnO0DXsP4AgrL6GmBLJgXb1DdOSL
wj2ccb6uzIpaSRemkTkDZycx27nuqHL2iCrpv4xm1GZtq7AAQwiZsqzgeAtoKigb
Qeh5V3HeSpifCy3Zeeil+MtBpq3xcrEfl3HclVZELgglZ/z4bClyUva0FFDFaPHL
PwgD2Et5q4w0MHdFZlBlE7B3ShiM/SuwRLYXulkbrWjSPwquGmTTRQ+HT+Dh4A2k
LanAHZlv2jRSiVOBXVttW/IzdHPrFwWpNsTa+2elih9V3E5I0rWuuzzeW4SNjRDG
txDLg7ytVocxc6IaydarQKz15AS8uwoxobairxChzsauq6s0GArnsz1eRqPJA1Zj
WhsEopK2I2933N8+jjvy27iLq9kJeAl8nqFgZWCaadrm/WFpbLnXGt0AIhcK24Sg
uf4mZX7Z4WhvkKc/d2wWI0Qu4WgjkwPpAdI8IpdcJum4Fv1wcvwetROl7X4bVSX4
K4MIsFuGf4Y1fd4E5rxmsvUf/wK+TRFHS3Q5SpV/oWWQbahA1cI/0pBrpYiFIDP6
glHoZamWrA0A4ECUMFuVARCYBzZB7RtHIHJ3JOAuGMAScdrYamB22GnaCvMJt4zL
7A0TRQJQZPzxowcYeyJtuv7guJHocW6CNsToSsKQtKXnlMhfmAb96v/942tf8qoS
4z7XEGY987KnkFJselsci48nMv5LlrlvJuFTx5U3creYXAsotft+Lj+KAZE0iJfY
fQwGgCuiOPrvSB1zb+QgiNjQ1CrzLNOLfYyU2XA8au/ogyfF2fEDiv2VNTi8tEFI
wfPgSTiFRAtq3HC6oF4UnMK9rid2ecldqW68oJ5LSIeUNyC43phjNNzY2zS6nj9f
JWX9B7sEXaKl9CqyJag8Mkzu7sXdgEBDNgf/yWvnxCs=
`protect END_PROTECTED
