`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ka4ChKz60K0IvfB/737uAq5d2RwQDS6OdcisQB0aMdbD0HJXyj/QY3zASKWNNBby
44Qq4YL+nXh8JpaMJ8iEAYPc0zBgXZ0wh0qtiUhnJNZw7to2xPUy623PzGlVxgHH
XsGi8H7/fFfxB/N/bAet+a5E0t3d3oO/WwC5479WbHVIcmbmeLPiG6wEQJeKfbJv
tzKfWudJW+ArbR4/sVzZS/0aPeQVOXbC8NROogQV9Mkug7H5rAfWfeLL2U/2KANh
CiWGcO/7gchrokw9dpgiIADH5WWc7jMF7Pmle3wfpNII0SZeomsQBhQk/OIaf3JN
igRHHXCssgclgouUeSP2kTNzVU8B4J1tJ/72pXExV+p8Fqr4VH/ehEyNpeno0nmp
HO0Yr6foYai3gApcJciUBRxok09kExovvJS7zSyn8VyrIvWTp6Edr2UxcvfkSutm
bKfleedBv5pIGsU3C3QUfG8zQG9w3kohrKqFsRT9m4JNRQKXpSaXQhiR11QBCgVy
`protect END_PROTECTED
