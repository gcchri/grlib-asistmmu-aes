`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gn4LK+MJlwYY3Qmn0AwV3JxsMdDmesKYtySnprMxml1DVj1ZosrKP3PZ/3+R3hi8
Fqq9xVXneosRCXRvJ4LfUCNWUGAXjvYM8ZSkd03VAbWYdX2VNfeT/WNYkcrmuFck
aW8i53T7y76n3JSX9ytOvyxpd/hOYSswglw2H+T8u9M3Wc24K9b+8Z/OGyeOH+i3
YUitclTeuTm3dOnnPcfN3SLSwXqdoD8ALvIjv48Zigj3mPRjnMX+mlAWwCAe8GbE
ehOg7sddTmwmM/sY6TAubb6JlGD1m8/joo/c3DM6JiZgbupku+CK85+X5Uf2FI1c
eNgHinuEEPsqDKdb0SuJ+DV1dabTf+LjGkE3bAMB66S4Az/j3Ku8axmGObK26WIm
fpqrO7mFRruEo+FnpLlJ5MSqC52+aCVmwMrlzgFqiPfJL7J5RZSV6+pYm6vrRw1n
cu3B6lnGKSIUjmw+ZxrFUEn9+dzw16LEWgDbV6OFbEIXFs3Y39uuehteBCbGGDRe
K+pR+49aNOxIz/pNVrYq0NpVhKz8Fj0N6iRsWTQVWEwKQpDBtEdT8iiY1Xbqkznl
t4MN1nSkePr9ARM/IbaAygNMcdR3kix0H4iLlmlcd4xomtzuDEi27k9ltm7tuM/1
P1J5YARefsOfhwLVKHZKMPLTpPb5Eeq3S3gL+Evb4F0wS0qvg0b1xf+UHlF0+fds
6vBBzDDpuaz1AeXXgwBQ7OYufpIxq2GSX4PZU2weJuNOZ5n0pjXibZEktH429Tg2
cIlEhsABULZZUtlqIInb+IImPMQj289BCS6zUAXFGLDfEqT7htJADnWVf1o1iEeB
mnp5JLKsw4dTEDyQ997uWHLdslTAMoLqcXDGQkoikLHkfCJDJOq+2Q4Udyy/bUpe
bik3sFmwqPfXycA5XH9n06AtF6MI1L2x2Mh0f18B7kOiP0RjWCLWs3zF3DpafHFm
71GJU2EV+afhW1kLFjubQ/9DTEbNtSZMJleUjQWEIRXqbjM3tLeJm/RAwH5yXhmf
wVL0HZT9RnfrrdCU4aqv02i1bhtwCWHwxcn8PQBXtxSj9xYlbVoPNaWkWpfG7cy2
NU973xA8btYDb4wzANJD0nZPJf0L+EjfMvgL6UPXIMLGS93DS+O2W5fImerYhjb+
wRt/+sLoQvqcCzpXM7/HJrpsvqNmxgMvAQ9E2jC6VE+m46ezAuhY6EwHIBuD4+hX
PV4mYKrF2uZV1Rj4sNUjwlX6NA9OFDP9Cirlk3JklzhdwdV4kAKvL1Da5+qa6l4X
+kdhGRWR0pJWLzFe1pvbWoQ1Q8zWGtaMPDAcJ6slOepVyex+RFVoTx0wV/c6INS2
n53nSvqgf5vOsDB1v729xFZsTkdhNlfJt5LVjfdoZYVXLlg+JxLqx+5F4GXLHPx/
vesSxg77PUcGjdB+A7f+izgtj4hRwfUkyke0mEPJa0FmF2Zi63EDUiKQaIkScgyA
tSMKkTQVLV1na6SoAyMoxpDyupJHVllJtpbycdkwyNtmqpg3YZzMtjOxRcZ+Y75P
2d98B/ewgcgRRAN3dP6pU3Z/VL8cMuSxMosoiq5n9wS48B/4NKm5TfDJQRj8ZcmJ
HxnGMv3P2jLqilIsW8Xu7F7tBlCXfmTYoOnGcmYCQABbs3oe06mlihU05GpT2CBY
zSto68ROjQ5LCyW1ISAwFN61iG+zchE07eVxJsArwJEPmQXa6C5zzNDqkcLlK9cc
Pm7s64snIhkpbroZSD7U1gKoX5LN4wkzA+nQ1g9SpAn7UziCHUaquxkd5FkZn5Rq
gZ04tCWSm+XgF8Z1d+ogT3ZbX+rNIFWn4eJBLKvC5bOJzbr5ui9CGcpiiAlzyLrx
HnSFQdqX5gJ0Wv+K6336Ae0yD0jzVNqAuF4IFlTNy7v6DlJEbvAR2kIlzyI/b8Xx
JWAbhvNjTey/HxiG81D5t5HUelqGFnoEctWe9WuEcH2J4FGIJqyeG3/1dOsJt0Aw
iwFM6cs/CFR4UWsxkojBY79n6RvaADnQOt6fP3P950obR5nDal/hVwAzSmcG4r+a
pbL6Ym6Qd9A4PuAFACb8uGbYFOfpU4EG6Zy4u1MUdyUNb4rsVnoTpUFBg0w6Z7Jo
Ho/pmEHgCxbtRaw32XP0RhhydDBLAcuSe50L6JS7VkBfe/uI7R0dvzbu/y63woFz
WVTxqgbu7b4Et83ARMpf9Dxrv6NDEOrSy6DanDJZfkVtMO7ozNd9qmyGOShdDDjp
KYs6FZOoRFfD1v7wQ81xXin2mIQHS86O0IRwxplJSJaIg4jjDcDV5zINg0aviOK+
Qa6Rj+V1hENlOfrIOcj//IIr5NYZPbp6Ig18OdhMHLSexEbzz29TAW1glydgSxfq
2r/KSruz1anb3X+DUdxllSjGyYMBMOL4gXJrctIlxtamjvCIfFEewBwOGrNqgUh+
+rMClp/YvDCjLuOD4of6678GMA36mq39PduGXjIfYRm3EDts0tBKBWq5ZHCu9mJY
i7hq/POGcwa1k8wfpzx1wpumA8xGH7WvpkOS5UJebXgAK22JzUdTFOORCN/+Ntlq
FqI4CvdBlKfTTZ+gxE5yXbgoNXCQZsypDYwMuO5oOJo0vmmGqzB1PguY4lphkiTe
5+Naf1xb6/li/Np62l43a9IIpj3pySoY+x6F8gpNQxLyno6l/X/JD3LmylmYb5s/
wdI1EB0J7I9Dwtoorp7h5dd5hzSAaV7IOFfsQMuR+MFIy/ZO076Q354L2UWN9tO3
gGh0NIIJHjOPFhEea0M6puFmb2U5Uu+Vyq6R+8fP6cg1rW77Rf1VAb/7RIL5t7n9
WQrHifUxe7elY/h6em10aVzAw3f8S8r5qPS4frD0HbZTafDcd6v9IuMbIBYMiIWI
7u5/GGN010colQtiECX73b2Ti7Uv1GNRB4XJaOTH22k9AACTXMC9b7lkadldz6w6
peHqwBSrp7WeoTtUDpvUK1rdLhEdMwaip1MArTu3jch42zpjw9IGXdV2Q7ErEc4n
d7zqGETb3OK0s9M7KIlBO7IeQzEkR9ULTQviKO6zcpg7O+QWFc3hfJu9gmXhNmab
niAPyrPdlslePsSdjDK636X8yaJ4h95jHVz1xErxp7HbHSGKUYMj7CcWCXI33bya
L9qdRafHu/xlrVRl9jaha5brTxSuD5SnatP/bJcYy53i9qPM7NBe0vko6SZaSKIZ
CmdImvYPs915vf9YWarvEYtVhmQCcxlDKmeZ1Our2oQNNc9ZAZaI55lvMxJcjWbu
NVMkguNqB61n2vbN9CFZ+C3dSR73CyFwHvOPevBL6sMjISbBABjcTDz2SP05/6qE
jx0doI0I/DdLuDRZ4Bp6Pu2obZKe5GtVRk6cJ70XHpd1y0Emwd6c7uiZQQasho1O
tF4XU1ABbOmQyrB85T66z+g19Z22cGtUNp9X2veuUemXH6Ekn0UH8AwBOLhjFwk0
d78COOCxck3NeOJVXmZoBCTUSYxpe6sB60X71RZKoQjwkC6AZulTVs4cb0zLkkPq
JlGf/eVhlE0OqF3AAa7o9DBk9v7q/idpe3RYnVAWVkbcgOB2aLlZKX9g9sEX9cre
zmJlKxUB/f2Lxx6kLZCpG3QSLJnbREswktZQKXgBosGeWF6iYPRx9+OeUgrr8b5E
NeAEJHWyFFAAkfxSjQiTWuw9jRlf0as19jM6as7/2mg8hDHOrZezaUAL7GC/mm4V
e4pIr60G8/8tL1iAP+LmssF85/Q8TNQ5KrrdOk/6oHdoO2VS2DR0rGS+9SlxBwiL
/MlgXN8cQhwQzAbOhIPdKISDknJ/BkQnjaCXXzQwbhFR6LMlPwTw07DSjcLFZZE7
osyg2uzpvZkBgX7DpQtaW22pTSw4hM38hPRGL5H95yakUDxcCVezwmKC6NpDkVmp
kXwdU46aPKkkJ6KQRSrOBQ4iqm1Q2GGU47KKLUlXD/srH687C/uhs628XY4g8gWv
GYB2gk2+mtXSbPQ/mKbMp/s1GTR2GsOQLrY2a8jlYvQ7aesm57j3+0OcWDv1Pqgg
sCB4sjaIiBSM6mUz82md+W4SCNhKbWJY0h4Gd9FGQc6o7kht7GAZvxbPKnZg/DWF
77/a4jQ3tPAHJe7jJ/warxkCXp+uZbebV4qtGUUogfaCEpKDPskJ0KPm1CZoPsEt
gkGKy3tIjai81mPGScfpUO6/w3O2khTEeCsKQW0Dcv5ieAyr59Nzy1GHs/PJEg+4
ARAdHEPMPw1S0y31nBriEq3MU6Chx7pbxqh+kSVUrg2PvwVIXUeSV69PPy6omtNZ
EDKeXqS39DsNKyb2ezTp8rspJCk4u3mToNDv4VNArmU6sf0d4g3Dk7bz9JbyWDmx
1Qn/gmCLJ5dvwsfiTjwr6bcXvSClmwO0EVZPojrMKYSLXROSx22Y6mRJdvc1PFpA
NTI8no9VjqGKLtrZVPi9O3wMlDEcP5tHkwhlLkk9L+b5mIXsl9jPdTqL6pF2EbGN
QqPLZlwS//9vLk9dTjY70ZKirxS2JX2lzVBt0q7nYqb89tIuFumcv97o1ostpteW
HKEHChuXv7V4IAN+KMTrlXunyOh+vFhQoqDZZy7nigGesJJvz+h/gGt7S3LniK73
5D5c0zmNMUorrl1iSiu9WJfhlyx1pZRc79BPOPsZ3PdHjLV/h7sny77L7uj8ASeL
tXJ469CZ+1DCeTRBORQct+CwsJsEMnMUo8P13fB2k3tAwicwk1m6i82Yg59cmghd
oktIiq4OfLbwpmDJxMQLyz4TUEMzOImVMBvU5I43/S7gb10OZETzK+LqhU2EbOF5
v3rAEhCCUmvfjec9LkqLzEtcUr3QKlYzsEhaMRkFWnKorDMXV5dVqv9Vo/ega6oX
YQU8OpEhUKmbVO7yTO2kvbANoMvScVWKk20QZKbdeYRED6gukJj27JG8dyUihN/u
MvoiyoQJrwpyBEVQehCfSRxlma5USPYxf8etPjLI02X4T2gOC73Hw/HLFIeaI+9d
BBtgmY9uTJ1Ii+8SgY/PS5ZwhHTICBE0KFgc/CYOLts1AAoVe3Bdv/OpZqHFqC97
EMZb1lYbq8t+GBWdrFTifj+O1MN8ZrUFc0+4oGxAgK300xqm2Y+KAHgbWXuJOw67
L8X/JVEfiWh18Kr5X04VF7YIUFxksLXVMA7fjq2DzPNuu1Minq9Tat8LquVzUlW4
VZVz7NREYaG26jylJjyCRqVwCHh0fGbZsjAl73dqiU+vYZp2QsC23plMENORl5vu
DkxSLfPDn/dGzJZaxk/bILY2hd74I5AbF3NTuegwkwi+mPbWANTIEm+gBq7v9z9x
oJLsJYZKH5cxWp/jXsk+APD9fuSEnEUW6kZhDg7Uw8C3195WlrNFjlEhhg97M+2f
N1NS/X4Cu388urmFlSEZ8x1Km8BHJzJifShdTDkCb0GrscWnmUsbxtoIm2+r+0aY
uU8ZSXFBiAc+7pmJRZ1TMXXO2e5Y8YxocPsMwny6PfBStEaN8T+6XQhxeAKlK8v1
ejCMo4bpoV8Kcv4re8jLcGrpCKce0z7tiicsYMoaRZn56GVSdtaj4eR03W0IRyYc
PNINtnwQrJFosWPd05vusCbNzyYkz0fJY2P45KDZYpf656xVM7uXlv9Tc5dadv/b
qE6Ov0FokTIVhm+gsKQghXJG0PTZDUWVqQZ7Hd90kkvGt+KehuQYqreogf1PUh1g
nlLvnLe179tM0Bxs6DJw1dOpVYxB4C8i9X0u9VpFdrJdcHZr+/YU3HliRm02M03z
L1pyefx3/28Af1HoRS3j8odx64xPUQXddpNfwVwgJfA63xyL05eaO8sKdWqwY3TG
lfxmBT+vvvCibR01IZa5Fv31nJIUdXZnQQWGrcrVL0EeFatRCAayGeQIBeKaOqOl
dGr4MRdhJ6TA1341YbnBgdaHXPMgH1nY2Lo0TzCKsI8MCiILj0jv8uaS2mgUTc0X
NXCo+arawjTam0uIuf1T4bsNuK5t+ps7g42FyTEKi9s19gLbbfJiyhX3MdVzYDl9
Xn/xqwX20eUUUwoaLPQz+Cbe5m/z+JQVwBn7ieQusrMTmajwMsQeZXAGm/+zp0Pp
ebk2vGQ0qXPi1S5x7uFfal/B9p43Odrut96oVnZbsm1pF2vuIa2FodNF/HqUYL2E
Waclp0Eut0uSsOZXjMzYxUfl7szZlpU+a8czl9MQrH6fyYflNmV2e8ULgYgM3S/Z
bEEgmimynWPd9KxSGj4WVKyDUDSq/bSbJTyPMvmJocvb2oWVOH7LE412veM4qwGP
iGHLJ7u7ZEfVmoC0k7PZfOvCaC8exuWWOcK0O+k3LQt+XG57pRoJEzz+k1Ljl2ST
E9hVsLZGI4dv/HHcHZpMy6zOd0q1tKUlmEWQj5E57mYgQoZCGyPoKQMYSUb5zwCZ
gjf04sH6ET2sJ/BCjmaxqgJjg5MDIp0pFQyZf+wD8emzOqpIsxRhHx0ZQTP2Nzgn
tVVrLb9BPiGS59iSlCit92H3OgXNNsBGWDvf+ZxUSghpBR8N+cWedfpz9eG3zXTX
NxF6A0gj6+1VgpWn0+bHvQP5sSkkX7+tD+ex7yOqsCIWwN5nvxx/tjXSGxD6733k
nsBxIxKmiMayqWxYDKq8yyiCGlmDYseeRNyspZ8bYpbIafML+2tEQejzvYXxiMPT
IHytx0wlyahRwMWx+EfFFSvpNyTBngRlJhjineEuDF/AKn8+h4IOdkcTvmI+V0aJ
mxIIKxSDvfICh1AQTRpkVWyxp9QZ5NQAXzd+mjdZ/1vH9GbOuDQQTTeb8vITD52N
YxVwAebCQIo7pGZze/oPf7X+p7AWem3+ZD5bZcHSFynaqazTbwkTFEK8XjJFg8+4
hrDclTursbvSZ8Ro1QQhb7wn1O8ZsWm4WSNzhETXUUf98BqPii1eGo7yKMu0ye1g
Npy4edsnZavQSEF3svYCa9ellcSa5plhXf8XsP4zb2HJPcs3+GFpzYVy1dCYv8KH
BFxL1vu0TsQ3z2KNbOUzjMkpnsP78lZxPnu48AQkP851p1suP9FdWnLL7YZSQiKM
HGqowGTsnrn++BoXezwGggg3njBVOzL8iL/4eE8NCFaeyNKl4t9Mp09DoLTWXh20
rpi7SD9LORihoguJm8p0SazpRRKunTU0IaSC/lq2qxUFfMx7/xSWikegblOCHE7K
5zCL52EAgtBdA6XU/Jv/w4eOwG0ELpH98ZmJok5Mdc6s+w/ugYlhzQiGJmD8iIxM
WcTKN3ms60CP8Dct+MsvvVVOM+FJVOgoedse8RAseU370gl0CgrqKsVHKsw7cGyc
4RnJDES3sQwrkDMGkySqJ5VwFxim4PH+6w1diyhbbKcR8mKRGodWN5aEnPz/pasa
TNxID/Byl7hmhDgkH/4L5EmH205WNGgW5WqHcbAP9PH7LDlRbi9H47pM5y3Tv124
R4IoBCwrkgbH6PUBFloidE52uMZtmZkDYf9ia9YblGgT2Bw2v9Tca6HG9Ss+41zt
SQxMA084DGFlCPtE64livsDuWsFmjSgD+CRGIqdz7ntsn9pck/RLTi+1WZ1Z82lM
yGYPyvjQtF6QpLljSOHidQJEmRBTonhNQQA9hxoDhOTGxeaPZMkYzQd+cFB8+OKE
PFKsrqQRBcq42cN67PxdQzQQ4vYR0TJ0wTQgkfT4Slw1RADnYazoAKn6d4sXF516
wtqZpccd+MNYz6PWdVwBBEhW6ucy5ivmsU2qgZMw3X3aA7ttdLHxoMGHmuiSnXNi
KU4qeaqxDWXea+xDF1PccuE1EA7YVrTrcqFVFmrjzhHwArTS2PK1jPSx6qHApi1U
3kGpMLgV5arpeZw/HlXsp9AOjNrdLsZtGoAISF2fkdPAN/b8vDWV/WXbNcQFFzWH
eWUmfS3RdTzN5rU7YOlTo2bwKG0+Oau5Qm8GpQ5MaQBB93egR5apGkuWBMISvCJm
gtUtaKO2V1O7uywUsrbqX0DP2jFK33eEzlty4qo1zAIjP1EUaw++yqKmL9meRMqZ
AQKiUx2vK3TnEgTGwd0OZZap2H0CkDH4rhsmYLI/CF392Vyauxc8ZQ8CrpHzKMRR
HSbEznNs4D9o5Nae0nGBetJXyl2xZT5HTjuhbsR1WE8C87uMRrtmzc8UIgNvjUZU
bkU8/CjJT7op/K9+E2rxvgnzklo/hjKhw8kCuzRoARnDSIKBYOxn/cTN4e1KQ1b8
TbkRd90iQZJqBFGsL26EbaXjmeY0/qDkVRHqtv+RNhcZX2jD2RolklM9gnNJcmgi
Ou1W4fPNGnLyrPqocEuKkLdv7O7M0d63hMrk8Ojyvjub5Fr823L8f/aCCSnmpOTm
dqwxQWJxGch7cZ/W9KgntVSLqIEZAqlItKjK+9JTOlODruQvzN/X11cwpf93weD8
kix8bXVaL2uLNgz1aE1VBeNEcJc/WuU7+0rPW7DoQhqWXJS7T+Ol/0GKamxSOF0y
lBAsExpFo0Z9Rim5pZdBrVaXQGxWuw4bUp/AOQykj6BJV/pZHWG17Szs9VODaLD1
N6XoKE7lmtLBQVrvaF8ri1dq7jhStwUVm8Sjfvgp6lmc2ZszjCY8Pe3L0WcQVhH3
VAdcev5scj5VOx6LOuXAo5VSOcufdpviaRoS0H2Tm6fyLGSWC3SIN7DG7iBYxIaS
ZApaHnEKuVZr55FFfJFU+xAIL0jn6dmC+H/CpQkPNUiXh3GhZ00aaaasDw+qg/XT
iSza0LUUrORiNvBtQADfoLOPxejuLDCIM34mFPhRJ5CFmpaop6Y7nhXt2xzHVqGy
uqaxew9Y9J9v3ohwUfM2avJLuA0a30tYScockPGNeNQoQmylpjyTEPvJv4D9Ngqx
TWQ0OKJ39CYdOYe+w6uytDsjFFIrU6gTFTeXMtHrHmMx5N6csd/H0coot/BKTgar
ZYPvxxwm1PGlWnWWKrqS/erl6BmNPfT23l9kfx3//fFVzcrOAYmP/X5MehxInUFO
514UVlEKSyxNoHBH1tUWNvsFlVFbm0aPILT0pYDLWpDNm0Ag6Ry8aIera2bGwbZv
0/UenWMzdvWLaxGNFWhGN+lm5exj6DOb7gLI8v3MAZhivaZI/LP4ff7nWHezujwz
4Jey9AFB5nW2UVbKMVz5j3SAshnKbxFiprGKfD0AU77FTtPBIUroMtAqwPo55OJR
itJssCcGIWaqBWojPE/7QmaWnI6XzKPzGzEeqtl73dG7/s1bpxAGGwc1KCQOKWtT
sZTV9vNvq3PcziFPN1yBac2Y/phyYKnLoTG3PQcIzLMCd0O1WPoG0SjZtkwAn6Gs
zweJeqyk57zYs437b9CCyu2buln/e82jQFmtIupibCdC1/vnwOwIj4/nEQaFyMUj
icU/NQXA2LiZZfVWj/tMnYG8ab3DGEQXEgxLBunuwZNl1QMIheM2nYOViqpYlhIq
gqorVkzSYqLVHFuDZ7/3gGJAj9VzsSX7xZyKjERHh0BzOfG7KIEbqYmTiFjJnwJ+
jIDS2m7Jwz906+HqYJpiszP675bUfloDG0U7IEFEydN7t6Ik+l1PyExx45s1dIYg
1J3Xt6kNnpNRqulHjWwh4q8hMx/R/q6SDrEE1hESfpvIkyjZP0iyMzYW34ebaqzZ
9C4GIYmJkKbl9TtkUounsJNiFoP1N83ZiGf/iZ7XEcMZr06cEc71Oj/SI/1KY+Bl
oHjusjSxezlg0aoyJu/B2N5JFFSw3HBGz95bKD0uwbkdwVw0MHjztNxeHDDFvAB8
4UsVig81j3x3QxHE1lNmROyR1KLCHSdPNPwwIZh3+cNm+3FoQZLCGAOiJvsbgXKI
s7cTFXxmIG2oJRk5lC+1GPdIhG6fetbPQZ13/zg97C9jyztqFKdLKXyidXz8oq4X
KGUgxcs52LvDuB05xaCafWaTZl4S73c8vqtdH78T7FBSp8MHl1B7islZgVjqLRgy
0o+GlJ4LD/I6KWNDg0RC8xuSXr3eWkEogZJWV3KaobRhGbqMZVp5xI3427YLHAW0
EeF5qItRsxOFCpqXfIRwymbFmt8VSXsZfeIfodLN0y4GVcFCewfdmhp7pw7D2APA
JGWlzmOCax/6++yPPJKT1iXJwfwDJ6PhtbkoSVk1QLCJTDw7xuVXAgTUiXUSMb6e
gBuf30bxUOvrqtIo62iT6byA9d6Q5i9UFvV2+pMO7+qnzTNDTP9wOAoiLXBYiLK6
BP0HSAGNjVgkvXcAFwILLpmIq2bKoAMu+iypBGDCsFK31B6mk0hi3Q4pRHx7BXMa
CpmzSKvvRijZH/CAJHTda4GPTJwpHB5qWP7xxD01pLUSxUwY6FbR5ORxn+96ItdG
fI57BgT6ULLFafNykhisKpYiZuwvK1SLr1eH2cw6su+JGEAMHNye5QLFTA2hHeyv
JvwizB4J15F47oNWyS7QkCDaBnVTX1Ytzl4E6ICUi51CCZwgtTqk1ot+GHkkTj7/
l0uACvAeMfx1Fp5MNfz9sQPSbgU3OvVHV4pp8etJSUuegG7p+9U8N81gj7LhwgkQ
O+U3N8GWUapag/BQqzMWZnikYAm1oFbxyoeSRH/VGtydzmkQpzB1aMEyQ+9l4mMO
GQf1NGf8x18d/7O0O9XLQkFlExBWEkY5aOIapx21DPuwVhxHISqVdPUyuEH0ewF8
0MrKtxNwHkXa5MP1c6hsJ22NsnqgCli0tNktR9dIu1Q/XURchwGHKPN/2YtvjlUB
y8GNmFVTDWse7d0Nd8MRnt8zE+RCZHPADWvX4+dmZdpn0BBV5SvOO07V5pQbhucq
/cvq9Lq3nCpwl3zjyX44/z6Yzjz5J6yEkk91nVz0b2le1BsmEDwR3vPsWGbGeOug
2Y1rQ9RykZ3BJBHdLyJNQQtybKnnr+AagaOoPpL6iv/EyuGmmyxhM2vl0WVKbiko
vrgAfyqYExasiUG4WJF+MAcvwirDB5ZMcOL85JyEgzSmY0XWhBahIgTVHKvyf4mq
A5y37x9HnrNgP8wf2vn3e82SEpQ7VHxYJBiuk9dLt6Ls+oQ4DV5W4H4CG0kwva3Z
NsQhkxuZgDSX2oEsPijJcEH7M4jV1+QNXsc6f9KE81/ZRGeQtRXz2iFUsGPzEsED
Jta5ZiJvgSD5kNg4s0lHj/c5tXhJAMT7buUVAZiq/u/HuHNUw6e9uyw4DPLZPXzO
p4ST6ESB3d2N/a6epCg+ALelkX1si57jRExTWcVLk5vrb0UYA6KJdErYNeAs6cuR
1nxKTpSAENrcqGI89L4KExqt3wtsf+zmPgcQi5FJPLwXzgS5hjBHKye1/I2D2/pK
kNpmqsZ11+G6rou5gIYawL4uq2bUK/IYUbJnu5DS3FVHPyhuMyh/kwSWUALqZNXj
3B+OkBIzhXO7z5jiq3WVSCtd2XY9leIf972tTA1emocKBFo5BrdoY4NRIthCVtUp
k2wbyguIx/CJFwLwQRHF2f6LwEoPxA/oxqnYu8GaH0WnTvxWVuuqEluKWkqZgw10
gKlKcQuBgNtdO1vJhh1wMWjUAMPl4KskKdSHECP2p426piF/lJ6ugLcaFqsOCzOv
ZT/KOddRlgRZwe5ymDDFJr5okWb/+MM1fcuhqMg/zzWH4eGENXuqqVtBxBgIgyft
mvB/+cdLdFyEQlVLy5YH5GRSwsj2pJTTUw/TOA3H1sDMXWbfdN5itjGLpGnbZr49
BtuLucmluJgFIfBIiyrD9/2vVHT5gjX+08bJ+Q5ofkEYIzl/v7TClbinKPs17R6E
KirPqijDKOJrhJ+zn8diowufYWk8w2udoaBR5+eaPjmckICVqeMrq72SwXxrtIWC
XeszPS4i2KZnb6Z/yMS7hEMGbdLxoYgSoiRxu0P7qp82Eeqg1dtxNeBr4M/JJome
i5lMj4j63YX+rvFvTpikXjx8ufZYx7adOJP5VXoFvjs=
`protect END_PROTECTED
