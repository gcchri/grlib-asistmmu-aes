`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yT4sahKF1HFLqkcjCgrzrx3Yszkb/cprQPEz+wcMRptMNjPUNXoVTrHyccvgNVwy
c6yQ+/RIIMGPQC55RuVioLpc4Z0HTzHU/eVpvl8jt6pWX6Q13xicWuuOxMV7OhZX
ynSigOo2TstI/HVADhWrwWhXXJ992pVpTHKFnSqw9ap4GCL4bCdY+xuL0Jx+55oa
BVnGTqBAxCd6JEAI9KMKHj5ts6P1w368zy7eO+rXNY7GWKJs1nQAYQnBdCmkDBzl
iIDHGh9O08JLL0Fc80iOAaxjjbEFvVoRKvxqnYvYo3AqIzvGmNE65uUp3hY6wlBf
DzlmEGsE/sjxK87+TqOLVL0gNhhAZ1HMVlgzBov2xD/U5V5yKYnBgW9yPdNfXHVz
Au7KzvIrkuc38ml1RmV5La78CPod/ZRIpyIVugXbV+drTatrTyITn1JkMHL4/REz
RwAv7+7YNkeoKwxzTiAv/aUdg6Td/DnNxkwsy1jVLGlK4u0YdII8KqQT6e4/osKB
ihVn4ZsKHnHRNPlGHtu+/o8S4CNAOBmhe9ssl3bHZv8ncQJmZg5sszMqkjQ99DC3
HpN2iyA6t1OT6oHO0gRQeSjspU5X7C9Tq0nnBDSVOPz2UbpgkSz8UCUDJTCNhKzX
iaoiSy/ciKhUC6Ja4hZOzQM50kmSNzumYZVkbhyYdXbKu5avoEFk3cuan7SgZe0M
Rrsc8pRGgHi378ZERV8w0o8+DEywN2WnM5gGkV0OXTiR9UfOBuum+OpDc+6COFGz
sUhU4/MVC7NJkeyXWXgOfy1MGiHwYPyZZMeBYTfOQM3Q+01dyZGwY1bs/7PCi1z1
3utIP6yvpzC1YymMHSduwP3xjptL1SNZqSrsZkiawNPBlq20YzteSPA61cwPVnhV
gq/9uspUanoYAF3tbjfkQhYajTFC3C1yeNw99qlC1GyTD8bG7RSlk5+jgp2D1DbH
8clgQkvrkYIXVYmnIk7vP4FYR/tp3KgHNN1XVUnQUQXitygaxfyh4ku+MV6DpE8J
21COCw4+kCuFAp8XfYQfxWpNEmDa1igRq1ph9jbteJOWo8H06mRqmEmUNP7srFWq
Z00AYOPDffuZ0t76LQ0hby96fTXIvqJXOkSdNqZb8F6ZQ2u1Q2FUF+vZUG3Pig4t
ewfJz2+Za0wwcuc6UUQafjlZXglk6qAJr6s0Pg1arhnB5y8tnITxbS6f0597ntys
yvQGK6JuD53KZyL5SHLkAKWG/H+oZj1fxlbS5E7FUnDUkTXJ/RWNxywHUx9tdbOW
R3HUsHJSbHpb23jullYMa+PZZEl2GBGnNjXQ0fewCMdX+l72kDXD+74nNNcEDGLO
DYJK5cSUPlslp631KoOgQpohwfiL3JAJCgq8V2lnwjZsXkW2wb0KDyE6jN0FkWZ/
3aozrTaV9x+zXL78kXiwjp9Ou31HGd0HfK9WPEjPmAznYRZ2Uf9UXIQZbS2+fXq+
Z1Xgi156XeaZwWYkd3YQbLmeMJUxCk+oS0/KpIG07D+xgOplb/34haIt6HuKHBHf
bN64SHucHC808Ky7H9zFeBRQ+umcoh2wfbP7Vmq0+dkxerjvFabPgjAm9m8Ly4aL
dAVlp2aB4dUl5TyzOWoAD8tIe/TPruPrzMOcIKqKk4OKk0OPSU7kHG2zMijdkRmq
Uh/6Y20/pcBf8I/+CM0usUweWlUMsD+rl2sWqWyTgQQLZie6eeJJGTPVS2lPZt7w
+IZlSC1WnSJgopPF4ot15yYf2rnk1LCu7qZoNK+fdGo5CAtDssmYPdAf4xXeAlrk
MQ0lxoZc3ONndFWgbVZFSRVpg49ONAoWRBWWLay7dQEcl7UQKTTzCLd17aQiCfAc
fDIaLNYbvf06eX4szkmYXcyqKI32eomP/TgRligvh7IdCrw31VeP+dSyHQMcjfyi
NjTDeHrlIZhxvMFnPJAvA475i8EK7zcs5PlbJbpm5XtyMv2I9taRmKx9hJF3tCsy
dcK9nYWd8s66leJtf6cS23kp+CHc/IsJ8zikj6iolG9O7KZhG7U4gRQFdQnXkDF6
wDIxux5XADPmL3CNzn8v/+P0RiM5OFy8HgbPZJDpflSQklADqIn5Qsb0SpeKNp6X
o2jv9nNgR6kZdZc7ke1n8CXhkfl+83DPsdw/51L3nL2mbhLDVQA39TgDO6iYr8B/
uWs37YEfb0/vlrSMJM4nU9ekhX8WpxlEm89m8UXTuotk0IoEDSvLqa0l23RVw7LS
BLfdJENaCd+rYKGZ41hwJjrfcriKCSddnctfynfatRcHOoqWce2/Q3sys/nAdqqb
YXoPZluRYSp0qeYMDRp8FvtMW1Q7UDjk7TGtPGc9DJVVVm7rQm3jn82+7FpyEPe5
8RdYEMTpMN2BBn7EHCCDn1EBsr1vGrtot/bqfhCZr9r3/YGi/T/nD5B0YlSWUoRd
IbO1kM+XJAu4KzJcpacq303fE72yzXqTa3lrmTouosZmQWxxzPtyOLm2z6pYbFL/
UIl3oZFqObPvC7R1CJEu6pxJKt2vfHcgNnTv0AgJmg/0AeJV29hOGyJyXjbV4JIO
MCygDY9c74xVqs4mOLX95J3E8RAo7D3sdJGkbL42pzD4iJHML24+SU3Hs6MJ3B0I
gMjmWRSigPRvbpJxgTxI/pDS4EmHfiFAR+qBdqHlGQIRKnbYiaQsH6kFJdugtseK
g3J/djXa3XyxcndNus73Rj2lxXx766Npn5HQoiCTo93baaL+gDZYqeM8LTubKfuZ
5Z5pKcm/+CpYLwS+ZaPez4JtjSNgCWhH93t9K7sWc/o7CsKBxz+N2AayuuKacX4z
chcq/fpLHx0AJEWAFCbAGXD9LL7LUBFXjEYfjy62dTW7KOjuttnGqBfZdC2oTnib
W83eU7shnGUN+vxk8Ai5hP+Ncw0uZ8a7WnFodA8K9vCrqFMUtE0Wqrb+d6Js8yY6
3HodhKnYCl4vajom/csYsazSqRJSdHo1k48DewtTH6GSBV/XSh1tt0Dtz7SNuAlQ
xEAFkGxAxwUjgnjPKaz+GaGN2BRPlnEikQjAlLGiJG2PR3MtT4bLLWrVUORGmOGf
H7qdaJyjrKuhFmHmIQuP2jpuT/fhEEgIFNsur3MJbqKo96iASJy8EkyXLNiITU6k
YOTzd987l+eH2cP49I/7IrMtUs/TA/eYFSJhepBbTMRG1cipdRE51XLQGbW4c7CO
VyM+cIcQr/j7HHJ+U4abJOnHuB3kfb7m7PylPq05TKmv1aTHQqjZLs7Am4gGUMbf
G3+45W3+xywzeNWV7aihVjdDjh+OYy0G2eRuC3W6ef8WNnF5KPy2xRFMh6648nq9
tLI9XLEqbMowgsPjKcZTabvJHN2JBJ9MMXi5GnBP8zmYC2aEzzYkGg25QD+bX33l
GlUFSdgHnThgoN0LXSjCDDezBk5uIol5+zhRmCYrwnI2+/W8Qhzc7p1TyswngBEr
+Qnk+9LaMfyjBwhBcw7BVybddY89fpQ1HZWY/Ekdmcv8+iCDzIoWEbi1f8kDBd88
/WBuKRaH7kSybv8+xXE7p9ErL/R44f3NEYvxiV/app7zZcb8dEd6Vt/aIohHZxxC
N6fLawBTfM0+Q9qo8EXFYFjQUyssyinBN1UuJjGPNtc2kSpcTQouhuao8u0yqX4z
xAwrnD3l27x44tpkAXaDIClOLJeD5Q90ITkmGCx+MvCGw0bcYpxKI3pfyb2CTuua
mnSLP9SAAB7vS6BlJpU/HFsvnw2FVMRp7SYAvUS7JdHdEnygbHduV8LeoWgr4akO
rSF2uVmrIfEKsIEeSUX78ytJyZhkEHwq4Qj4G91qb/M4aEMbPB51ru65+3qCmVHD
9RKJhslC+GC4YUykclQzUnWS1/fuWPYnWcKJiz70nB1xNr6Nle0k5GnwIGfe6S9b
zrfKYC+c9rZaEklq5jnybB0Cu7OSXFoDIUSZ3COAsgzXOQjOf42/DxDW+x51vCQk
0oLoVw6DZFKMvED9/+3qA/nFs9ynOkouk7Iwu0wiVbcj3Mc6b1WkV6mXFBGqByTE
xspdBdoldXdtgE7BMFjM5JJXSZntWwF4hFG2Ff44qAuGSnMnbOYSdZhEQKSyx942
F+jNydB1u9q6+EdzP2qeADk8wGqjLKow3DH638RB2xKrKWvXplHq8RbUT31upXeo
mqVqZJupGkKX1BmTm0RvZErTJIRCw9tOE2wiIIhkXoLxKs8YVZZ2MADXpizxVeJR
f9Sx7NaHrWuEP7XmAI5ch/Q5zuPpRQn3yd7t0NupIp6hLihCR88a9DzO1b6UNJSB
Z0b/GItSXWU/LUwKMZDBBrITN/hvNZ+CXU5Vm0/V63+hNBpZWKHBEfzcxoBNeOVe
NC2ZuCSHBOSo8ND67OJ/zKYgUQpO4dqdUuHFybTx93hKonhc3n04XdSwojp/TeYr
+QjVwxLaQ46Gb+QfIOSr/ys8kORiGLMZ6BjLN+OxWAc1irk/xVWeRxkFUn6RukOh
W17SAAs78KyF3gf+3erzZMugMuWDWfhYCJnD2BkNDlwGd61rPzsY/TTGpGzhDqbg
he9sta2/zwYb7p7iQbFx98S4Lr8ieEKT9cw21AYGsMMfjI4t2ETmWhUXt/+2ajMy
I1+3I10HUno0ari744bGwrZ79ut0V4kizDtDe1A9IC6GJkSd5/Le3dn3w7NwOQEY
nKpleuQA2nBR693ckD9J2q5i0DGRvy5RoJzKCi1tMTMhKlcIA3SxT8qN3h+H/K9/
+xD0RF5Lan9BrV/fbh9v7fVqDOKpTQov0LwfCorb7s4RiTYECWKq+HzQ+RRMlKLy
/ROCNCEQU+K07Ilrc1BfbTnRXYzsnzlFza2oUyyK7y9keHAMsxLRPha8b65M2QPT
3gJIdAXLHhZPt1x/RHdzaEgVmTSFCAmwMRQDulv8HUg/8HtEivKQa9PUCtUoPuga
WfO0M2TCBh/Qgf0ft7KEGv0b1iinPQArFy51SGfOHHQyIJnIIk1EQGIC8ZaA2GOR
uo1xYfRu8rtNO2mHvz3AMjM3Cy0vUv/7M80gnpkthCc1zXkLw0dkoujB+6OV5Hmz
9NR2kAs+0/dWQUKQ6ihQMem+dvGCDliX4IVfJY+zFgdvxMF8kIi1gZdJZPZb34hw
K7W/bYwbrN+CTxK3Ko4dzO5IEYJVBH8uP0JpxlJaNwtJuht0XpUMqIRWdpFAg+ke
7UIFEfrtkapg66ne69E7QSoqsLNW9YNkuxSElc71LP+1OkEXkkQc79QIiXZVM5sa
nisgQR199eniu5F3OGj7oSuP/m8uQl2cflPW943QbtA7skmNYahB4oEZN4hBTJ+6
2ESfgsrgYLS9a0VYAPckjYjN3b7+90E4OI3dPg1CdP4LKbx/j28Pv0+d2zoHFlEz
B+h7HA2qOZcUaBeQM9MeUOCgqyB6a1cmY6p+H1Bhud7Wlij+Md7g3fVv4zavTXd6
sNFx7Yjz6EOsQNlvWeoRxHHF8ZBOORQChFzX7DmqN4ITDBqFYbijZDaN8Z20Ji/o
mjrHh0ixwDD6cssUedlp05pQW0vdRR0CcYOakqilQu/X2VnfeVFJri2ZtlpgpBGn
NxEsyIynDmtoI4C6jtLDWzVGMtauX+RswXACbbrO4r7XoqGVJptqbFUzsvEPcZh2
yBNxStl4LgGHtY+2CFbn0jhE88K9PCp8QeM7xOi4JXH6HHFf0Cw4R12VUVdv2GuT
uKXI21a6bt5H5k7DpnjOWeTt7e6/jdeSOCNG4cpZ1XHAyB8D7oANHbJNMpHI3TsN
u9fBnVGiAud5ZbG1P+SWdfNrfEuFy0mKVDLsuliK4uvSDMdem7zbOvHouY18wGwX
XfFMqp1pBboGnYTvxEQ2Mz4XdC8VCTeP7jCQjpNuO2vEq+beGJMsc5+U1inSzWu9
88gHsPY9RDmXGNX9YsXxmcc1S9uOfvSe2NI3RXCUDZ7gAr5LKv/PJaQ5mMeW1D1N
Km/gd7VIIDwbcWqdIWdTX8ZqkCcL+NpPRbWwYQOBkiQo9gZ97dOUrgYImQBP0ppd
a3KphyWJ9aOR9CqPFdohNRfXGm2fdjbD+hoe83uO9cLamwcu/E97HwGMwGu+yav0
n6jHrnxq/VJGwv9cGm7awIvFYiU3lIQotWQ9c4w5PpojcVC6aoJDH/K04k+ihPSm
yHup07YZfSn6+PLwF/qqmkyNUHAHmjoPwTadV6TTbaavhAVHbp27kg7z9nwKrqpi
3qE+6ZFfVLQEPpmql8+UmWWX+MabdbjyC4XJKTR1XQoPKWcSTlbfNiG8x75YLnBB
sv7s2Yl4anYmykYncxJi4SvQjzwZpo8vbDYhgK+D+UgZrlwQUAExoUgdkBPFkExm
IrSPQlSPnTQuRy2m5bgvHaeNd9e1kLeOsX7Nrvr8KjFff70NskJsD+M1iqQOxVCX
l9yVM5zluqYWkgz0p5UJPIWb2l5leAfgcqKZhD/jCBjEv2WA5BbiaY747yQT2p56
uUIX3WmB3iOBVl0uHWilCZEWstuTy6cNGsVpdMdjrZEXey2ekQrCwuYQ+3FpSpS9
JGUmdw9U2IW9aOsxbvBBFRycgJTi3FGRcM7YCJD4COQTzd36In2laYi2hZ50yMxD
a8rWlSV2LxpOOl+9aZ+JrKx1BlQFcWi/JW2SiHU3420WD8J9LNuWQ0WTZ46zsh6M
NLhkD2QpUZmiz4kpOcMXiWcrEp5tAIdpVZZ20Za7WO4+tfspvW6Ho0DPg2Rm3Yzc
6ZXZATss4xuYOQzU7BOZ9K+K9Y/fYDjcUIUZIpxoZ+6XIQSiM0v+a5rkJzEi3CI8
u2y2dLleeZrHzSyHYKBENBgE8Xc9/KQqVLcacKDHMozjV4JkAF+krLdsXwZU/Ik8
BsX8GlS179J53A1n8TWZ/HZ0ltfHqmTXCQ7m+Llu4wIEz6DKGY4sjHy8+oOlCwHO
iUOVrWAquqA0JFxnGvmfnjMUEiZtEaj8jWcC44Os4aCk+g5BWtcOXhkIXr5BK4yn
z+jelvpDdS+p4wRI6zNqxW8ltalt76j+f2XXvU1fJuLK5b0GXlKRuO0CV7yfw87O
x9gzooRwoyI7Jd0zcArNzCmqzVUFYHgSZ3zdgKNfCL2jdETfg6khuwXn9MBXbR4m
mewad+X11lCMUmX6RN78qb1pmpGrBrjmdFJQcKUE0+N9Dl9L1baiaYjHKarU231F
UrvFJBgGrUbdipseDogWoaCGjZLnInxnGi+DqZXv7QVC1nWa5YeaHMhnROpt2nrf
oGQ1Nraw2ztAxbyk8+lxpBZaf9NMv0cguZfz8JYP0dNAxsivPA5dqVQCpFm006xl
sm26B0mjEWvexewkHEdsY2oP1T+9ll9HT9fWO/CSVyoRbhR19EUU32jeUCkG06oC
gkHYPNIROHEMGONLgBoUoPMHYfNjfQjEqup4l61sTTYFjiF7Z+YV+sAOxUCJR6wR
0erJ9YHnXvW5B+Rd1GCpCnPlOalHsn7edXBirUVhJjhqZGUrPpA1pv7Y9fWDwScc
jB/XKjYohD7gFBQJhidsxPIWQD8X8r/GYDfFTooS4yWJTt/Mt0z7OViUSJo4kcKu
U+B/j2BUaiFdrdXn6dMRDUlLitZ5qMP2FL54OjrBHLaEyecgNRlU6Fz72xZ5oQ/Y
QNypZ7iqUOAYkKBKZgIFP3ljU+Elg5qPAgJB+kurgvqamc8jDDN+0pJZPfT1NfKN
ES44djAeAh+W/RRLkM/0h4A2ooZd4wKhdeJrOTnUy5XSW66ZMP5kw2+wq/DB1Igk
uHwu6dx9FmZwazO1MVnIVQfGr0NjIJeA+/BGHeJFmJNYb1O8kETZaaV0WF6nEE2c
CAckJ2Da8mo5Zd/IBp5lp2AC8J/7zYbSBbsxBocjqVcK9pxxQNABK/XOJQw87bYg
vSWvMM2juimfwFIhN9DBg1xECNNaK4Sh+znd/JghwNJ5lytujKTefjhtbMp+gM15
dPe9KSfSZEC9iG+HP7ksSEAzcXbiv62jdk2F3cUU7Pa9+mkaMXGS1v2Zpwbgg23R
zwaLuiI73eWhcvQ6E+5FrDEicJTY2Wq4nZ+AqqP+6A0E9NKhATYCqqes/7u4s697
1gkLEjOvO5p0LyEkrd+XHpSStWOq6QN1cK9NrPct49Hq3tgQGFnLxfAr0x3d0Gww
0Jhm/+BFQ34RbKSM/lgUtGI+Wuc7Z9yORaJw7Bsl6MDK9DJJ7pskBBHTn4udmGLE
emDxKhLigUSH8quaHZj5d+5Si8lsKn4GjUK91srLSpeLjeyzmzg87AbBf2azupF9
h/WNbHzDH1fNL+yWGLH3RMft0GnpAVX5jB11FlNP9SZrb+WmExCfChpNfukhSUy6
xI783BPtbRqBqa3I/Cy6fJafs5vjJlb07wkwwGuhEZFOiotSdrTaTFdRZM3ANpML
Oppr6XKw2YHnr82U/16BYc35z03RxV8Rsnfj4AZ9Y7k28HVlMRr48T0vICzp5nQH
zMb1PpbuRmSfsnvb8gepoFWPSQIzuHd+rO9OJM8TGKUcZvYz7g8F5vM6BjJQAR8G
ssZZx0ya9BB3LOLZE2joFp5DwF5LAAs+KA0agTF6rY6vNppavPiipsVfeBqZx6ST
SUf2L8PKC7tEjMTvwNY9TYZWKWvrMM55NcsoMi7CjGmmdmP51tXdpvTP4TDqRfZ9
NB836D75v4fLm23a+VLmHplPzuDiRLVWXl73K6HgJBTptewWKjaBnjGpN3y+rl/n
a1w3QVDYYmigePP5BV4u+y4buWngYjE6em676e9vMfFBZ5Ec0NCrLAOU4KKkx8vT
AZfsrr+02eAqefKt1PtgrkqPMtsj6Voa8UDCrJsXrok7yx+zvNSpExPthFB4YqzP
Zf0PSl7vm7XrZNkv8Q7VFJJa97nMJpgAg2Wxw11XbnpW6vWpATWjX5LKo75lpXAF
xe782ISP8ZTK7PJCCuAHofihVtwI2KsBYQwPbQqxxJ4x0Yx3iLafbHPYmw5lqbM5
M5Mk1wuKjSNiJo9JxDfzF0thXi7Flp4AwV0SDGyOMqgGhheXOC28ewCbs6TY0wkD
RtVouyC5ekp/OAof76sJ4hY+GDMgJPFiGdCOD6oDE8haFSs+nrdn3SwahIE2Mqyi
Kfk4tG24SfDvmZhdeWpAX5HdyBXEwlVb/LBBxZkz332On6V6mCc8ioa+1/MVth+X
BIRGRuLRElAV71RshgWwqd+ohP99yWh0WqnSIwWKVmm3xC/D5ItZ+JM5NE7Clmat
haCweYq5YLdTNYFzVY1esS02UwHo0nkAQK96NKOx+2HsQbzHCvHUkb4RIo4k1rpa
x2KyMbd7G4pukdtEK4+AzrY9/4pWoTWaaMXBTkF/YpUiHHzEyQMmGnbV5y4s3Bna
yekYnm0SVhUwgFhj4YnG5t1zqujkHSAVtdNVm3m8vtH4TO3/LnS0OxsPnz8Pt9tW
q12OPE3CNxtOs3R9xKJcsJ5LEwch38l86CSYEAevEOoQuGblJTz0CzuBUFWMDqVH
5+ZlpENYMDz1eBZJF8h+2ASi6k5ffF5zdfxkvDd9xTdLno5dMxfKVg/fhKKHnySS
1cejIQWTyruvmKr89Br8kDsxp96OH/b96uMnbviF/l9u0N47D7NPs1s0PsidNiir
msldypMAW+BBT1SJp+33rxbskcUk86JXES/ZXFlqNwEbKBg7wKqhLIOfbxqAlEpC
owtuqofQ70HU+An98/CwvqS6v4qRl/uKDHqBOZPwnBLIGdeE91mM5QSCGHWi8/F+
1291R0rUr8osWqYEcg2uYONx78rvs6LK8C/ZBbFkZIn6GlL8P83hiAoJjDkrtldR
6NfELaCBFhTyyNfuu9NRuQPeSzEFQ7F3cQVYgZhpTKA2GqTyBnr3izRN5EXmhzpL
hq805pZrCC/zDek+mR09orBvEF2qgpC6jcLNNUE0Ka4l0RMoxkpwlXykFKCjT+Vk
YTARGIve8yL6G2b2w8wSMw9V5dFrMVACQjNpj6fO5RQ/MTwzh0gNSLAAlR0h46EC
xlBbNjzgRWCn/R1lXqyjPdNcWio+ZC2pU0S2BxOHdqijQp/ecSLfwr/Sn9fMCppH
fObD9Yyex1wsR7nR7f1rx1Ax/E4RgLafMzsXdK9fuJoK8E8FwAAt4VajdtzE2Ol1
wKF2N16EKYZgfZ+ESkx96ZSj/b7fv5k8BPJJlzSKPVl4m2XBdtC7Yf0GG05qdaGY
hR57m+aot4ZCfHBL3sr+hYR9PGUh3ZHoxGJgfCHQ68v7zR4MjR+wYXcfoDNvEvkN
f/NluT866UNL95JwyR8Sp++X0tVAfEys7lCMD/JTrDeY+OrkMrLbpD199KGsnoPj
Qcf8FIBM1ctFiLIAhuJUdxzmplXJEfjNIJ1s/qVhCRZIGUJusoCPSdev2ms/gTG7
T5W1JcfRDrzX6dBrXp2wT2lQCLnmUDtIWBIxc5i5YnfNMq3RhrsRC8dgOWPq99Q0
F4iEnpWML61OHoB+m4Q4TOucn/6+XZAEsY57w0gyiTENn46OaoInDaMeVi5gC8mT
ThAUQRkpOmmSeqrMnXnksriFkQJdkzgB6JDc54Q8KFV0tYfpHFc0pki13bkgs1Kd
7f96f85KqrcN2NPBS/tqTz/26acFvKq1YmQXsjAdv8wC2IfgKF2zM5SCBo4fSlca
3PlLQIXKqMWbLgPEFRvWE8qpYfo0BTSeSJX93M68wZGimo/jUdO+MadYO+7KfcUg
lRdLcE1Oegy88oi3oWpKOw2EQE+TCzmxDaLRqlbg2iogOYwKAyMdHGXWmc4T8MIu
sq3ZGyBgC6/xCuaiuNVNQxZsTd4Ye0PmZaKDD0JBEXoWoOKYImCtxq9l5pfuVKv2
Vv3HOBO6cW7HQ4ewFIEMHjtUzxFdvWLbvVwV8zPh6NdT16kDgN1vem5zMxeoCbXY
gKq002Nkp7b3eRP1ZJ5OyWoyRIPiOfoesZKHKj/SXqxF6YEeCW8ikuFky+mAmQaH
WA+KLVyEGythg/gUBxJwNIu//KSm2SGag2azZ9RtQ6yh0qEVjiGo3p0HJT1bL+KH
VEv8elhof8udHg9Ww9mJq+USs3sXKpEVAWAcXEg6AjBiajOG96eN0JuOb0KsYc/f
SkCLAln2/aO8thU+58h/lZK1GXvRAwRrwf1O8zHH4fMVciEAs/Cmog7U4iomYziY
rEww/hwvG6amcFFRg9v41qr6ZXbEqCUOPHyajp6BD0ZGe7cmK9tKsCzy96YEWuas
E8Pjgw9Ca0fYmRLCciyWYzs13+KSkDAAcrPfS6GKBe9f3mjYIBFTaDd7F5I/+s9A
GkFalIQ9zDJsQc29pc2gQMVrTV9sAB7NSE6REfTUig8OMFouhLSv/mEfKjnuT3MI
xhJeaghBKGK6yTYCArerAqQKrYn5AqlqdQ99GcUMNNcbvbF+YmeWH+yAyATaPRb/
0OXucPIG0wPm9iDQq0Ib2SdJruGUxqL5q4LMezyqQ1xn72AC1z0YrpJG4zhzpVnb
kM5CIjmbcHoSK3xZt8jUbWNDKeMvt6gk7wKYgJ7Cha6upnD5ZjickxG8Q0V9GPQV
xfW0TfyakFPVtVC0C7w8e8smmhSKnA7TuuMYoHHKpl6zvswE6uMTz/4P1xPt1vzE
VUJT6xgXm5zeqlE+DHzZk2ufSlcn71HivRJp1p3AlVcvDnyZNJNX9h/qAtyniheP
CMYpGIbAmQDNZLgnc/JdYAz3zK+5XOc1Obv1Jfac89e6IXqjCaelgYCIAKYtHcN2
pwK6S2vxQ+oyRSxT3PTxHhOEJQeF2ZBk3b9/fxMqab1BnA/Za+t4/TEY2nY8yQLk
HPcDuA4zSVryOeebGrthzwXqeX08MAMT6dPGP6fWAHqGERttvnYgcvULp9J/VlcF
HX+TOIuhl8zPBVRljKmXm+DLARvYmeL8a6guZdj6nJA8AVFrzrmflxDRovJ3YiJ9
sdUsr9mKtIEnOX86dQVBbC1OYTP892JUPd3MRTzVU8BdPilBlmZVe1lZNslUleDx
ztrtk6xpq42HXsHm4StdILFGdKAydi5mlnM7pz4IwWyGv+gnvQGLmrHnbmHWoAqK
OjIRFLfnEGfA4CCaI330POryT8XrjxMURhX24ZyDkMtbtk4AlZwuLG04fYrn893L
RpGJmhIZAft+SoRMVi3TyZVjYAa1M8sfahqvfFdyME+RTX6rRfx2PyjLCqyGghpI
hN0wxY0qiZAjsRqOXE+gX3YZnBCT1Vrcgptwg/4riN0CU+rjtX+UN5+Q3UiyjwwZ
+ByILtOWXbvOmgG8K9fqSZaEiuO2+J3tOyP0jww62H2gnjoLO55wGa9EGh48X6yF
mnAOSBGI7tRyZglXsc4BIoZWKEbb/ipI/eQAMVczg1gKoPDprWMP8CP+hY9+bIEy
aZIMQXT+4G8KtgJURPuVlNd7/0eRUZ86sxrxcuaztdTVOfsLQEEmBY35qdLQEBXf
v7aKVIfq/7alUmfGn9RdkCN1SEmS8+TbouVjt2uEpvxVsGrKJT07sqCXRazAULis
sWg4C6Qb3YsTtLGSZ/cLirvgCH1eGLbIMMLUHwRu54iu7hwW3OwqXOapxbzhSDL9
pjCmNG3weZYY6dSBH8asAKWMrSwIOJGUXLo9CIeYvn2BGSnx3lpNEXnjcCUnRxVg
LuCcxX/pzLvdYWqvk4paFEXJD2HwPpQtQrr6bjGDtc+lx4zV6aj1U+IVsajElq5I
9Rfn1tPCq7Yx3zX99WjKGpSHahtaKN90Ixr6/Euaz8cS8k75GrVfHFt3pHGp9Vcj
ejA+MzHT8zWa3GkBTqj1nmDzDMDA6caywrQQHf4egl7ymgk44lPG0KXBaBnhPdnJ
XSf6oNOI4xt/3BF/d1CkELHLfgRhejVYUxK5qYiP4dg8uPZaAsUK+Kg1lG5GUMZR
eY3fmOeUbrAHF0VVlc4Gv/NVZCjL3MVBsDxBEKunhOHE+cdyWhqTH781hfu11s1/
zUQm7DuN7Zfmbnm5+EVfMC1GhrjbpK5Sqzc8DswuO3hx7dZhT3wodpec5fPuICm5
QAcMxqknwHtjnlD8UfjCH7eaZv+O3DijKIpbBLA+pta/mWmRbU1VO2BUomqHzVOn
DA7xpV3cqnH9XPLmAFw3ZLg2J8h9Ia4i9qnaDVrwm6ujqgfOOGwjCCkZh5zoQPGM
9ZHWhzo5WeJpYs/83dpqaEj+CKmxrltyk4+65BCf+MuVPo70g561eIkbJfCqlNx3
VRGlUyfVjPf4RjzN90ScNFDYD0wczTo/Y8qRECu+pIEcEwYyUGd9qtvvmItadGgZ
NaeulmBbsiplNMQmZsf5HkVLT00I4Obdkpq6e76+2NYm5GfOldJMY5lT6GHBnxAs
JELe1TJGaFd/dt6N9LJ7Daiir0NdmY99vU5Qtt+gwRw+HVEaw/a345aYYHERHp0g
EWa8B29K8T+oRskT1yc9bjqoXwSFp+pFRwh3yLmD92KW2+sk1IMwNyDABVMS2qXK
+bY6rLcQf/crZ2jrEP1PmUJRWA/sv9orMg41gbcRCh7VSjxkFgYV+qj+tO95XUvC
9FUijqZn0Rqsrm6d1aGi4kBcKHPXViV46YAUc3Z+gNaGHIUdgp2qyJ+ke3p+f5vu
ph5mxqKItH3jdppoI1SJdvUzBmJLcmzE0l3XHQGhOSHG83yofk9OkEkpqL8UaLQL
IUzUI3H9PLjsRr4WARlIuRD5MHn3lE08MhcaNdgMyLGnGt/Qf48IwmaqncxF5SnI
tKCcqiTmVJ6J7uQVH9QtC4Uk7SL5Cp+sbjiX1X9tTawby39dIoFmaB9yVmV58fC1
GbEr5x/Vg3ZIt9AFImr7/i282/5A9Fk5pPEl8lZjXm81rIHidB+vGIERUWIJjCCK
RmPXOEk+19/99ZojqZp4u+Duk6L0OZbgS8Tlt7g4tcphKeJtD9EmhtskCfJXzaoD
vfuY1ijKNIjWfnf+thfw3DION85/AG5BwHv4e0iQFUckCe5fZ3VDNZEhDRzy7XvM
AhW2su5aNuLl6rWhpaSevYZJoJqUqN2Iietc55INwhqsQTdvBTFQtsyWGtpafIsu
F9NnbGsL4+UISn+k4oL5j/rX0JLa8aOMXZ12OHYPaY0RG/5FFIDLEzqwWM6sgmQL
vc7cJRIH+eTxmjJQhZd5MAOT/B99KpafeMih9Bdns5gNE0e1XwrzOB+fJMLPGkqm
WwhX9hDgvrFG5/A6oOVO4uYlQQ7GkCAGi4PYIyaZzXDaWm7ErLlEFDiXUqqFlC30
seh4lHCBiBNj+cx2w5BaqZRZddJofNmBrw7cemlIWVR2knBQVM7xK+NOaUiny1rE
cLSzUK/+yL6vyoh9r2T2Uwilv3t0I5YqE+h4NpMVhASPHxSlFlKHeFnlNoMbW5ub
k1FLYr4yHhOXPQJBoaMd0yMBeN/pehvs8VqByz2JC8pjdRvWt7TWXkyDf4jTLz0z
RgxPWM24by9jdbWVoW91yJyKf3HKXNHOtTcBRb3xcn3ncmZRNPyuDZZcIs4Pcy9i
Ot/ZSTEb9cxglG9bFe4Kpqt0Z8knASwPSHJ/r6DHbNyfiSlbAvtKv8IJAioJv41L
gfJad/OryMYk3MDMHdyIrZibD72RCdGHKwBEyqoUpW1Mj88hGvtus2Ltp1SHDJSj
3BBtZirSILcM7XrC8qOyFakjZCJTLI0jc9VRpXtleW4wyIZqDB9mI56AodKGR2o4
YaG+Oq0z5UHFoxFZPd3PRoYY0hUYRQpTj+dvKorCltAAtibpOS9TgSp5BuSZbRUi
s1R3eGvA0OPoo6ylWpWvRFGVwP3ks+yM4x6539+WxoAnnYefeDIOg1/R4illxCLl
q6KPckiPTyqeVEgxIyjSDFSpwuAiQ7kvZIBc+ooAy0bENxAPOKjBwFERP/hPrUF3
OT0A+FKrZIjf/MJXTzz9VWrMxnbnwNe+9inCZgWsvBR/MFmgJM2cnTcOcOa6czzg
WydHd0cztWnubQGQj/SkIrGZE05LklGr5OWFiYIUOIHMHVlAyISMEqeZfbuygmSe
Qkk32RvxpG/rkNfNnkoeLhLZIEBuMusRdJnVbbI7D0tT5Li4lju2oIsygyJMMXZP
h75OumMuHjZs+DJzFEqZfsr7KpDnFqc/wEAbqDY7o+IQ02jW1CYKCoxFGrBf3kfN
KCDZdPGm2OznxUXr16U16k12XOMtIpbCtL+21pqP1ihDdnqp1YPB8/sb/iVTytD2
7ikUSRKLhXQHgdWYxDyj4m0+q972+cJjP/7XLyoL6J9YwqJm7QkJfqiN99BNJo17
Io4fBH7mrvdem8bwyhX6dzHxBQXyPEOq88Hlu+p49yTWoeQb8vOhNWjAl5BpACcp
QJxNvz9wLQwvJtYGIb+bb1278O0yzAxTNsZjzkhUcsRyn0qMx9WMa9Up8BXKEg3H
WK6/M+L8dYnG1nRz+bfcA9A1Kr3Tj0mg/kB8MpJ+7E8Nyx/kPClRfXvNPW57URMC
ESZUG7AoH7eKnc3DXp+B05F92YR4IzWaxGZ1lx0EvOdhuNxCkk2lyzAgsati8Nle
rHvK05HV1oA0MUxLyt25tcGReJLfzfapMqtm6Q7OTnuou22+ew4Cir9m21N8XnW1
j6YxCuv+MAMrfzyT2VIuZ6G2AMbgMhtj4as10XUGFXN4QXuK1EOqfA4EzcvPcq4r
jB7wOjgp21bOnXBxBl1AgHYTO8cUhQbZAI65Ubgw/evcjKMGnsrHM9qpLRrqW+I3
dQFneS4k87yKyuVjRZ6EYhS0wEw3ZKTsuGWPg6ZSCKE1JfZnUESVdjwZXfTPxYIo
MBGJIoUcgw4uXekEybycYAq1nKdewBQRBI8QjoLiGhOx26JMNtcThihnna5baoau
47kG1Tu4xPKvtRWzTcyi9WHT1HW1/dfyYQLOVtK39o47TgnqKDr2zYz5LqtUpYpv
J/XeJQm1ywBwKte2Lc/UONo7olTXq2Kw1dqMT1DFxnEDb3vTsYC2VLAcQDNoRu4E
8uHE6ZMFs+ZYcZUAWFp5TBeUewbGGD81Sker8cr8E3V2fePXUu497fyqRvsEDjkY
NnrAca3qviT6+ZhR/ZzV3B8tqW65pJi7TF7yPqHJ3agn5ipAulxY7fB5GzJg2KGH
LPxDgWllprHgdpxp6n+W5gzgB98pmA6tbIv05Sn7W1zb90u28JaLo7D/QObmCX+G
n4mhGRWB8zkqvu3H+VkpeIJ8zimZAfl0QAzXkoXFk3I4HssgSIOEoSHk0901QIEQ
WGYKXlhDlwe/pXG1TC7igecsi4qWkuhGtLqhVSH+anOn8ghl+Cog0cwgISY/MhdP
hqEBybTJVlGG4g9sLhBr9h9MTRoO+0TENLZGMOpwvOb4R4baFiFCmiHamtJplm1f
Y+XiV3bIcaHoLVs67IjiCXHvxn49TEWSxs8BoLjXfwQ1i13GIlNXuZBygLkdNHKI
rj2mNZE/nPeRjVs/Q9mwkVpdDwHuyLn6vhYCPZq7KC5h2idOG6GiM0L3al0p0VSz
kxnnxJoxbl74TM6sGiFmSYjbidQRvUzD1vNEh4SF//1aPMPec5n3H2t1oLoeOTUy
3/euRwicuDb0H7GvntVhwWP/hzPMFjGUDpl8kQN1bPhA6zw+OKbYk5KS3wXSVllk
W3ZnbPoP0DVrXb9mSh/cS6h8ttrSUPH1RTUDxwYhTFw7hFW3otB4A6MM701Gk4eq
XeMWZtEQdd38LaLBljioc6Bdhsu97RcvKMRVHDTUJyNI8rRY+sFJkRDhLNLFgOYB
0Ktf6YwoA2f3O9+YqXk7U0Mjsuqn/jJmRLsM3PzIFqKa0PsyuNDC1ezX5GqJ+ctT
NN5nKpc2cCUdGU3NISrvwXbzOGNnFTzmCc+3YLQEqf2AMIs/atBNnm57Pey48LPZ
GOXwUpWbOv3Wefmo5m5T7Pobjym+2yJWYvNXd+bpeT+eissisVO2x3NUXd9BZeJT
a8bX28/Alyj4Mjh8QaUSAN2thcDerQ6grLtGO5QfaMQBA8o/mFqUkdeLcucak/5q
u+hlg7hE/MoOth4L7wkQ2d1VwCgDDieUIydMT8lVLvjT/OjZUjIiO5xAIKGagQtG
d2ZgW6ohNGX7l4BNWn2bP8uEb0akGnHaQmjGVOpNFiAVlLWjPC310ciA4FGjCMi5
DuxWay3sl0XSCjYd90S5Gpp+OInFxmmmC36eMzDAUkGs4oSC+yRqOU71zIpQGers
nZ7ZqujcODVIv97fWSZp4glskTS/TUVoAEvjhiOSA04aGdQsE69UeyYuZ65tqTNA
U/RKR1owCkuql7dPQGWuTnLIpQIgwymDIYIqKDows4qYncveuTEb1sNPzLURE8Xh
ZHgNWr5VAIjyc+H+akkiGA/tOFN22IP1lSP3tzh/ZHiw63i0UMepmEQEsEWdl4uu
cFrEY0+zFFoBPYg4V/+bJ711F/HLPCg88KV1LzlmguOsgp0qXsCjHh0e5kgc3uLN
zwEVqQA0huoqJYjPS0xRvwJAZ8wvQbmeCPgnUu09EMRIXCXzGdJRS3WdrlOHWpdx
zlEKlKHi5q+J3tpVSyolm6bQ78aJJKwFuigNHfr75sgtFm7MfH/ZBevDld5Z3RXG
BOLGnF8FqnW9PNoANwdsrIDQdy8P7YsCQlrN2SC2QVLIYt5yBeN+mAV/ltTCAHiR
cQHnnhWB8zr0toGTBFCz6NI3eaDpX6ZX8sP1fbQCT6wWTBkU6X6J1tnd51kuAyXi
V71a1R1Bh2CIdhunuqgsAhDOhynv2o2MO/cC5k+zArg40O7dUEVZ3lbDeH89ZQ5S
zVVbZxxDKrZhnmtKARhVG2/Fh/uKcjUQw4Ha57fboxLBHJSUVF7YtD7CWdT+TNsS
+OEYpN1cKKKgSMEW6uRqUzRlUG9mxyxFWgcjpbbEWoYjSyc0URbuyZjNYOn2Rqow
adhXWF8FO2KpanasQO2nkH6X1ECutfnVaM++tCKD8z4lYBtGdzJzXu77BO2jLcce
WOvGpd9zt0RAijjLjHcj1g+cQY+GcginwAgn8DL5HeYSf2AYXvipFfn8515duiqI
nGrTilxCt20cGRYQhBId1LOi3NQfY+Wh2SxRjnD0LVlFRmvh2GDwTWw4xISsLE8h
GP1GltfqtMW1aBlUQzEyVQpyujU/QU22VRyG71cSsL5mR0A5+2nxHTnxE3EX64Ds
0LKtdCuIPGukuiBrLuNh101mxppwTa/Pqmcmj8Uw3E0RiHX30Sw6BxOASDWLN9X7
jwJuTYMDCMYDakYMQ9tsoR3mMtE4E9z2ZI0qkTo7gwNCSA+YklfRFWHV0w8ikMCE
ARCCst/PzPOBhbUdZtqNFmfZwDrYOhTqWYQghk6J+7IEAyEnLK1CntRrqXbhATJs
9FGMUzmKUU+kdCANeo2oZQOD2cXydhHvXyzZHeQgYtn4MxZOB8e6VgMVX4KDhqqo
W4gMe+szK1Rrjq65vrpDEuYaIr8EpS65aCG3vjzaUkFFOd4oUBUcSt0q5AmuVEOs
QroUJqKdGQD4jOVBt2qV/PIG8WZTZiGfQJJ4JaMKhRLQPWq03KOd+JhwUNgbRsGA
XwDkhyC3ucdcRBOu7ICZQEGL/TQo2Bm0zYv/0g2KsDTMqJN7LzvoCNfa0kHSQ4R8
xi73ie4cmeQ+BzpNngjH9MSyEtfhohcIXFejJ7e8Y7ic32Hb2Nkfk+bD//0YI6xr
uD6cWDEae/oT7uKSlRa29ePFeIxem6fX+dTjTtwPlRzzb9grIpgSPyFGWojYlZrL
/21pn6a+ThbK+aiyhVNq9bUcd+N99xm6V3W+GUfEme59vyIX2/3t6FytZF8wijeg
RKS5BxIXfr7tL1tWzz1cJuQoXWKjjdoqp02XhfwIrP47eNXpsUhzl9/WVHRD8KYw
e2U9OGYOdZ5OPtohaMlqibMRLNNNdHqJa7HnALVwkyKY78nV9JF2b/6xDFyJDiY7
ykfcy1hq8b8OoPub5xx3vK9m6PbUdic4VPjlW8uQ3JFHcZF+O72sb0do+aakXyEQ
67A5CeOlt1sS9DMq4nl2uOl6ONUIuPbME4Xg2p/F9yg6k/yoW39toUyeTTopSJuQ
ppBfWtWYovoyrpmToBlsqOwcd2StMGIkmsSKsRsAW+PHL3MyEoKy7+R9XGrPCo3A
31g6nXtBSIIAv6chwh7QxBzE5DYnRFQZHx4dT2Iw8YcxAZnMFnA9jNYgC1ofoiZg
FVvEAyWxhudEWSk+uW0ysNcdioa5+aC68LhHPux32WxCasWim8VCPNrJegvuREan
rQUINJWkYpz+fT7GGz4CXDgYj2Jn99KR+Cqr1rlz89QCIADKOIPXLs96O6eZxUIH
MO0Qekt2fuJzo9scdtqswsN0WvpIQN4/J8zLuhvyhTi72Y988ZxWDm4XnIpcd69n
Qejuryr7iuiUCVzH0Xz5K9yiMexDGeTC0lXdSGfice1mmJ/+BHFqiZRu4CDJKoeC
Nw1ovjsvQUscsu0jDKB8UoGxafBWlNBr8rh5SCkcYLQlQHFSj9XnsyVZDZhEHBEL
MzcyPxGVOBcC9bJQO5US1GsJ7c0a8ubYvxv3I7a0e3ZlvjnKQqxNm8NY15sIodBN
WexNKuRWvpPZmA10RU+4j50tVywVrE9xKg2pMnGwmIQe+kVG1r8jJWu8nu5s7MRk
OkoRqrKp7EBWRtLN6OcHhhCDqabKAMx2Ow6LCZwlHBz6jPh6qss2l603Fl4Jwl3a
Mmq1+QiBfb65So4Fzhw9eTnk9Gl0YiKV2mjhjbbOOqh4/xW5rS6IKMxQTux41N2Y
+h7IT8uu6CANo+7FoqCmGkdvbC6FcBxVRo/DfuhiEWppnT+xPZooSAY7yRerbKk+
tDVf71ulbbQ5Aayxt56/BAZZkqR6eTxihs6iWMp8poq3sleH54XLARxhdU+drP11
SLsk1hHdvhe1oTZngmjXzOcC/0OghJq4ueGuxqbiV0flVDr3EFdjdiv+1AHp4Te0
iSCEqrSdBYpSaWG4sOf1jdlfkTeKhfAaQC71dgaD/QAr3egHhOJ6GUGHpGVNvoDG
O3g2/uTGlyEipRHTzX5Cu5OJ827TLRK6PiePvlmYuhvaaL9hGugBlNrlzGHpgRVg
rCWuemXlOFuq1UA73jf2YTZu6unepZlV7v0guKyYYhHXwQHWEs69y8NkuNeP/zrM
tEuTjWkW06ygVGx0kDFRaob14++tP58+F0/MsLtl+zslTIUA910UaFai0cyacTzg
W/y1xZYc1GTcpRkmbKBMscWT5zzboq8zG/sjO+T59K1zbyNCDFH7vihhixYvaKSe
PNOq9O8zKa1zayJkVVC2Pfm0qBfgNmjD3waO8R4iwyEyi/VoyhkdB1rLyU2qIDo+
MIEI439LK2V+jAKADNuwhx/pos6vAupqkaA+GPjYMs6fr7GaU3icSJ1FFyP5v5T7
YydNX4eYYSABbFeLQDTI2PxRNboz3s1sr/P4L2oaExjx8odaimZ8gCNbEzl9NR51
DlQYPY3xVGz/fHXMugssO9OSPW2AtelttpDSp4TkYwNEOhHoKY4amtyVPq8swEHS
KxxduiND5W8GvLq6octrAF6DwbDunstTfDLbRt3Osn6nOyFJ8RpsKralAWiOnNy0
FSP2c11koqO+eMaHvR1h6KToPZkoM6X1In5vkmjDtnBhKQf4dHqdkWx7OvxTC5C1
4osI5j2HuKRWFXTI0s/LfYE1UZW0D9zdhyz/74yfnxmMOSoJwYJbaMWblpw5hYyg
FWmeJDWGhalGHgU6zYCCtGI3sW6AUcSeRa43gZT9KILvQ5cjBwikwo2bXs5DNGJf
Zckf30EEYUT8NWJYh9AtTNSioOKcGmsVR6zlC9oZFS6D5QEUpwxHNq/ThvPf7hPp
MUwIBOKXvdAq4GwjCZV6y8UFF+em/QOv/cr0lfUJ63+ajbKULmDxcjdFbUIccO9g
xsXYG0grp8cbYWiqmRcBkxkFFV8xqwqq52E7Q9KK55DloYbqkoY7irg511QCQ1RO
K13qmv2F0zUJo8X3gD8FXWeyPNkQBpkNW0KYkhY0Chkn0vJ5LmbouQEopQtHJToY
UWupoAi90ttVvHF13NbuOaHLwYe4bAk5ZCSxCKL59pdvI/f4cAJxdBojYSm4ASF+
SYasRon/CyVAAzdfxsCmzc7sSTBzXno2erc3AsgUnQpgYxor+FdUhvDMyOz7b94o
DFV9R8/zc2YLWZd17o3HZXWsqHtQ6+qMfNeW0MBZJZhg2Fee1BuK7BwEGCJGJtki
MxWBl7dsC9s4IdPq8Tjm7Kk8awd3XH5BctOKTb4nkkwHxkm9o49zWlrsXErtK3qx
XpU/ZshyhYdX4hwZxtAILZgOap7jzpDv+9vnT+LOuSQE486txgBHdxDKo5nN0/wk
d7snUeSzJQlTOtgImgYf2aOyH6LWXWTqB+2a72ftm/frEv+8pawsp0V4FatIxfHN
KqeJLIOrFLcSTmhQsHGBN/RcDvBfmTFOwRQ0caBVhHE4QhSk16Kz1v5+cbWS2h21
1BZiU2H9g3cuZIJC7zYM4J+2dbZW/ZlCHxpS33nDrGdtHsP/KnPU+Z6JH4M75Jsz
OM/FBBJdKu7s5hVCoYOAM5J9FtZYp2qErTNzgOQzQucBPEA1H37H8V+f8P18yujk
qFs1yWgokIv7F3p1/BAqCYCpS2xWKfa686SD1l8vJwAwg85YEFXGHZZiqAlAqr21
+z+vi5UbXxDyWXXSZXvd0BoNUQvYpqcsl+T3Rq5Mz5QAwvYQBO1itcv0Ts3OUaSp
vl0oMTWPKD2XWkqZjXfjZMz19stx60+Mfx63i1JQbp8ydOQ7B0R3DeOymK1/VXZU
O5Dbk61gNqHE1oCQECTcMMzEJh4GsDlfORRvfVh3L4B+a8ZhbB+IxsnPf3Oabba3
Yg7+B+ehIEDuFqkmDnRheVIDUtvvNS2QzsESPpO2OAG0uMOD3+wG7P12WXUjiC23
1hmUQwt51H0WGNO3zgmSxOAPWLgG+9nf6pOllpJcOWr0fstx51YlZioO1XaHUGbU
tavvwxGDJ5EG3m002BvxprP3ka+WrCLvhvMkEOUHlk0MQoSCLWSS/WxtXMnePrkp
lGwsA1WWIYSrwsV7ccceQLA1NneO1nWd5yRKcRPMo4XxAyGCuUETeSLmlBYkWTy6
UKjkeF916hnO3E+R9C1TjAMiBPslPv0clzsJ+yz95FsJz0oSQ3Qgob1CJYY0qcyB
mJxxqC6c8D2Wtz2ev8DARi9AN3tsYEaE9HSm9izXT/0UyhdVF8LVWKNpudGO88nB
vXa3pV2LEucE0qW0V8usxIW/vio0AiHKTV8M1SIWGW3gehErjiKsiOZuguHtEDkA
pGjYU5v+Wds4isgYDw4mlS8184Yi7ifoVFzilqeVDkDGYEv+RaWoV46XacsHXKB1
1onak5/Y+yANAQfz7tvoEgt3kSIf/IY+lxStIbJg7WRNkjtFC9OOT7r8jENm/XXK
YpFaAtb4kmFiiKul35Ft7byS7MmRzFn6a9c2tsleP95kzmCLzDxewRIgpAudVpCH
JwB5Xydh+kAy0s+6qx27rABBIuVgjG1XylGQaYufOadl2kBT34I1xzZu6AO4+GLn
o+15UaEBVn0fGgX0JoE7UxCwzJlUZSvrW9OC7rEp6343yBs/GZP03LHEq2QfPydi
A4c7wG6Y/9iuvpgtJauWFdj1PYdoZc4XpVnNahsif+d6H6YYQwYH/OKCNcDldC/O
ZFEcAjlkARPi33UwI7xbPbyaBDZhGr8DYAJS4idssJ9Pl9PBeCYzT8KWOc7zbTeR
iFYuN0yeeXuh4Ym50vFnt5rT1EuXFL2aWRgSnkrirXRrZx/SEUbeokTlpyIjYXzr
UG9E5blU+s5IIfqTqZofTGid4KC/0USsONnKaKySw6K/6asmMw9p1j37mdwlbX79
EYx3WkmhVay4N/X5k40c0eWwySrH00yOGrgmjiHAvE/LpPo839Q3Qiq4t/6hlZDQ
Bnd5JCEwR5VoukJe3F6XlvfUJBnV5Hcfghc8UpRbDV18I0h1rS5DKFlKtgk9I1yw
/bHu7wCPIVa7Un1bDDkHXMVZTq9OJHYmvzBXVVS0ANhPX8V+4OWRV8kkFRL0DINP
gCr3d25i0xTlMx06ggInmhbx934lNJ4sdd9lD5cSA14RoTRnxyyIXqF0+r+2CfKL
8pMCaaDqXs/CZ7h9InY6fmvRauSi0zBGxUNbVmSNOVDHic0UzOlU+KiTL7KQG5h1
qNVzYaVF1kabRnHz04UEpwZhc/A61mSD5mkjWcQ8OsUo5F4cOo6h4azTap5DdQYS
nCvzHlweWO+bbAEcd2TSSJ4N4zgERZ3bIgMMZAWVCMjAvlj0T/Xq21rfuEo7pGSq
GijXD8/Gr2FnEnq1qCLTg2ODbKxQDCFNf6OiVFdcYb/FW920Ln5GNZ7wxOj0h8xL
04wXq3AHptlBkdqeFsJEqTAZgvs7K6L1Prb3yYJ4Lt/qQ/GsyRxphCT5mjMGFj72
vUm08SAA0w1qM13Kk76pQfrCzzAJJlZsdXT+KOytVov6BBx3KeL9tpem5quHUQCx
u7pw4dsqz/s0WnsYL9RmcY4j8R6mCrwzq+WYlVNvuXs+UCZYUSzvlwR6yWI9afVS
XZuPzedTbXVvPAQy0iKd7UIaERzncBfrY9ORRrUr4XPm+wqhQI1u7xMhUzXIU95k
xnYcZWDRYclKAcVgtyaYwSbL1L62VYxslGJpF+DvmdsLNT6hPF5RGV5e0A3X0VcM
N3cr83CJjtWUfz/NFqQmiA2UDeUIks9cIaQGshTwnpD0qFYmQybshuj3XNFRa7tY
LN5UgXiebubHOIsLIja97mDSTIYLDgEwJbLfPFRCyGFFafb7tbrI+EzK2fk97HkT
vbltqKkjEJoDSxO2lPBg5hvHvY8hUzPwB5lwn2fvyjRqVCzE+pj/BnzLlJDJ4gvI
VtuFSYuijtqVvmBiN8ATdIb/MbDq9K/ptzWW3R1LgSovMUDJ9z2vXn6OdlwXvukH
Y9jpPB5cM2Mf34oqWGPHrsqIUmue6m+HGynF8Vi/MnPvaIaidIAgEKjNuLRm/+B6
WB5hdv2e5YAmfl2dWDPAovsQ8OgW8dTig2uvVcC6K72NlbZgNc/g2dBKCFoN+ksq
Ss6xizNaiL2XMntz0jlJzsWBd3b8+tNbusWaWjSOTlRIbEKmX5dl+hXr2DBGEqS5
OYzZDhVHl/zBMu/Td7jatvvSoH/S1rt55VulcyF5di7AUvw8QildHXMyIYp13FJ6
xE3UKp69isKlCk/6Z13wd5CXg4WynEy8QGhd6tiTpJN3aSJ/8EkaCyfnWWMqktpc
biKCW9bz+51vu+vESlTvFeLDfCQofYH/0eC2NRE4EGykPo31Alz6dnaA+DYCj/E5
DxG9BUz95v136Tny5QhbD3Rw8qBSJ/CgDbQGmU69kvkZpL8iu3heogzi/X8GdPXP
QSeE8TRejt5taP2LsdMUActLlzwQoasiOpKmT+G6NP8c2YK39svheYhUk6AAArFV
QJye0GlSt6COspVHDJzbzo1E535OISAbtoH86fwIlePR193TtL8t4aEUTVPIBaXu
JSAQjKflZRdYaYdBUf7erO7uPc8vTFODKNirU3HbxkbmLStrxO9YXeWADqrpx6yL
QBftU7HyFxsIg5vBiasV6xvQX31A05YOYiwT6LF0o+IZIb5sulIGZFFDH96cPe2M
X91/2aL32AbXIy47wUQbn5Suade3WGD5w5ijUwaC8LGSnUxGXfAiBKHBoO+IbR1/
n6/QX09G3X2WQyCqx4SgmbAYHkqW9nZuTnFtTRecbBzL5uPcgtPrrAGg+itxXaT+
XVn4rWCzfy9E8uDX7C5UOheVoQzKgqYwsksv4+ZW6Xitu+1jxg0tp3wZEG2stQYc
s4FUVAwlW2FrSGZ8y1hwhN9n9h9GXKSdxcjKP0ZwUMIL/ywBtk7DbXF3/XQx0ES/
YPDrhM6nywNSSsxvqXluspLtxIg1iJArzIgzlBlQ1x/HJWt1O8o+Xy8g0ruBkoNz
7OrulwjzNi+NNBO4xn5GQ3DjXkfYMaqATdy3CqzpRwVFAIfvWHRP413FS4kTR/a3
bE0Drz7jYoQ+obsKRUYoGhb6iX57SzVUL4cDK30Kz/Q1KIg5FLdJvLuApm3XiRgF
QeFr4d1Hkas2pfmkmEMttQGydRSTEMh4I3OmC39cK4ZSwVXW9xoBNi+vtuWUGypl
d29se2+WOpwfILyPLaeYFJzRlGveP7MFpbhitGbznRtXvVpOuZn0TvQIyZoEfnFy
18nSZA+XA5xiVA96QAEqbPogN3ahBZJ9OukVcF6/fz4yIR5ySyz8z+Y9ZqH/qy/I
sdExZo1V2TeAE7j4AYbdsP+1DEE/031G9N7jD/e3li3IGYRC00rSBwBL7sMGRQP+
ujqhP66Hkrs1vVYXwiHy+UFCuzw/Teyj0iYoYRxxgjIl/V4ppqpU1GlML91dODZ6
QNyI0PW+6HjARoqU9YPuLLYL05O4jTVtFpySs2I3Cj6AX2ekwdG+xRNBfMjLRZBH
nb9euskAI4hQxKG/CgicdLhKQMxdoI42iKGkCgIPFznEfA63Bz6A9Kwk4XKPAtuL
8VmWmj1tguXkoZNqZREZ10Th0+zQ1D4JWdy8TRgBeiMY3pMNUybRTsLBYtMwlW7r
gaUZ/aAqSbVQlH7lVSDh8w3DCLpOSfn2mIulwVCzMe6vr4547tp/MWiqHnbvHxMG
qAcTs4l3LTnQ1VFPyuJLQqWqLLDA2ULe7qmvkgpYhhmpfZA64ddMsE4T/iAHMKe1
bAnOC1dTqFT4FOyzOEbtFlhmeIC7A62GWkO5CqBJKhIL0yYWhwpv4TNN9OZbM+EX
3VSBBuD98kUYEX0PAxFNjrKsIR6DbEJ1dnFyUWjhhCNqBFcDG24z+WmKNKSl39fS
VSCfQJ+Ebl3NhOFTW06WcxjWJcW5B7zccyCALMRB+Z4edclsDouJISAhmcaZbi0H
tTRoyetbaKn40LH3NVdgKf4as4pbPydIZvJDnB/JRY/av7T+7MzlbmA3SiSPThl2
xEAyBVxPGnX3kghua9rwSMyJhfLgJQGOjuDMbFhlURHz1+ifU6cEDa/OxI1fbzCJ
UiTTIZayzMy78sfNwFAFC6AHGQu020L236ZREOlchWM2nrYIt1zKhFjzS+hZzu7u
6tjSZyRifPdSkAO9Y2EGlnLNqSFPT4SvoeKjyN3K+iA9mB3fTN1iewpimT8MTRMe
QSeaMmRyxHdC8Q3IjWPxOdI9KO81z+DSedWmi+uPpKyl1TiFoBeR1u6JOOAZnrNa
/87bjF85M7HPlfrpPGi1Po9g9cFyn4nTUl5vg9nZ+/4swJYYFx5dDghoo+dg2avI
4gJlbw4jH9NobYzxOhzzsi6gGqy85MyCtRNsr69N1jyvdBAZB65xyraMxBgy1gR6
oHX4aL2c5QmWZ79SwPvmyV7DdxbjxXB/YfYHYulGzt5VsDjf6315QUL/JYX/lHOx
e4KeCjyoRV5trcsVBNDf5sA8YGzAJj7zol51+eM1fIqEyInscGzNWZyGRRQmxRVl
a8RdkG5604EBhPiISn87/JGBleF/qWUrD0oIBwWd08vp55UOXTRvpfOGkpTsCzMp
FMEadhH6LY3SJ5dlhsuQ8U60uUhCSjvzVT91Zt/idUy+cx2FvDxSNYmQEMACGsE/
6+Blseorzoxr8dQuwQp72Dh62iOcxJOAVBn0i5qq8+cQM+whHxyjgkdKlDOAVDjD
s+2pmUTLgjf7WvbE8AjDhV6bE9iSF0ROlbKjDFnxSWHn+dD+4EcyOHCacoIy186R
1IURRm66LA7PiEYw/SPECy9i1iHXVTloG0n9OB580rUL1pBF2kA3L0/E80GErSl4
+H9fJl0cxap62a8vyOm4faFQr80G9cazMOa24qbf2s1l+8nrCqzaBXJ2Q+fehbJw
enZHXxJofRUbKr0jkNBlTnQs6ygP9j4HGJwjBeOUFWokdHis/3u4exnD6y2cOmg4
SQtXVlX/irUPMIWumhF4Kh8wWPIreynXZWd1uiEZocgINt+o3bpVs+BIlLi73iSN
64/2Rag2eWnN7H5wP6EncpwiZUuKFDrlyxw1PkNOfRWqZenTM9G5+kRA3D6MWIX7
breNvKCcBES7EY6XdLvfFP2vKJCKB8v4z2oOjCLzdyV3VpKnJhcRsBNBKzNqOkAs
UiE0pTIMDaXLKbClf15/O+IO4MMjKWqzkiGVBF3BPyjyGuSuKAXXZIiRW9BivMlS
JkeGw+H35lTjmq6KoeRfDFK6njZ4sbyoCi2P1k3wtUZn8/Pqjm51SF2usw0F21zB
92A79Ed4n05sJvI7xLkk6IerCyN7oMISilZhwpg5hOJaSdAbwu7VVsAyBvKyoCBF
fYoDuRhzKIkOoZofDd7tNMwQBjJPwKojc/aEfCBZyAEusG5RxGPy2z4berKr+Ebm
vi5AeN34DHOBi1r26WS72/eJrGdTTvk1LDlHTVczXVNN0+iSxGhwNz5il8kjKwkd
/zT8dWXGZhoXzwdARjgmCjf6F8a9TbbNx05WuJusBvuI0haLUAAaLwmatUZMA+pf
xJVvGJZYo5B1CaPLcvH79+MBFtgrzTY8QWoaNPgGxWz18oLhgc5Fz5xtT2pxhBD0
k4bCEEv6aO9RdJNcZpLchO1NJQXzueH5tMC7B7BK5Rts6IVnpcxbmCGzAKkLxreJ
vwYYGWOEdk1n5KPksnxEbu1y8HdazDgSBViU6aHLcQN0hapFMcCra4wwIAYUku14
BgL178Wv1OkmJ4kkTGULXD784cxGtCo06BWzKgJAJl9VUVuQkwtIBcuim1ToqBYY
RlygVNvyPsE2oPMuE9bwvMhN1vgStG0ahp5+cIIKXeppDvIyPpo7F8KseG15Ae7Y
WSjwUcFdLQ3K9QlBNetRRlasroqcdcs/Z9/0Y5Hf+f1vtaVugCjiaBQg1JGFzozS
ZHgVGfy6h1yCouvBYag8rChioKCR+kgZELzOQ/P4LyuKxST/7opcWOC6KIhsKHMo
EHZNgA2vVW7rFWOjsXMQ3swW0YZpe2RUCBB9al7pfSKuKFrTYGxqn1e80p6PkrTb
swNqT+ix9A6h4TnY2npF0uDEP241Drdle+wB0m7n2V619mqyRBDRp1vrgWGMSOXR
8w5Ghh8eFBMP7JJbDKTA4Rk/e4Lxe3PcR6f5XfxQxksTWN7GmSKAqKqVFtgrB4Bq
ZqFwgOaLG6lhZUrj5sLpZyOQACETd9oapvcfWbxq/yQE0TSdVocB/R4T0gUEpa0t
1PG6xbbRyl3wrzZD2rmQ5GQlJ1DUZkQ5Rnxbz3jypPHP/GkXWBhiUDINISu6QWPI
XbedRq3tJwGG9d7OF0wLqKZRTMzRE2c3XMoipcw3zY7KJHIF55Uf4W0i0KzyytWq
fddnZvy7BA/F3eSJzRPHdej5wAitDAg7BrQChpjJHcQ2W3FINCUhJ5+AUngilB1K
iKxCngD6/B0Z6zwq+e49MwJLSIdPf8IrMGUDAZCAx1St+1itfMex007PdGm7/h2w
7P68IMNu0i9sdsqJKxDKSFSYxp5KYyIHI80SroJnZVJhezjYVONItiW6VwME+Tst
ko3LmWaDR/38LAO8yrXptsWdCHqqun4AMdW5ckf5Xj7QDP/RpOJu9YzDMr67nTSE
biKODicwBq0wApWxfGc45QYR9l/0mg7jZE9gO5mxylQX4C5PuWUz6CFddFDamour
uy0WhOeCAJkrtVdA7i8G1y5X6pgatonGBMTWlfwAJJmnpMc3w2x8pgXhO6tBjrNI
tX5CX3QC7wMEOTfotypv6nTN8O2ZSj6bMr6VvaoVYiZPFywTKK8D64HGnT2X/lei
7yjgVSmAJohrvGpm2xt/ZcwgBVCCFsACHOoRY4Zi8w5r8YIch+1QaOp2eJQdP4Vj
pcozMyUfKXtYwl7+4QW2pZJT9TjKndleuKjTLoGSSxJTQhneM0oMLqKdkJoDBPAM
CdDdEASFyG4yiQ+tGCxRWHsGjtgIAL3X72T32NTHUfqJ72bQrezHOF6dtmotRjlg
CKZWP5TLIrQAgxB01zBKgZtnWfu84Pz0zB4MqXe60mVk0m9gd2pff2hmFktmXfYm
1JE0ryVvehhsGEMLHCSQi6hL3Wz31kHCMsV/Ur+UucjhAWqZPLzUrI5Ye5l3dzd5
GSj7XP/U7NMx8M4zLJIbbh3n8IsaKmdOhirMzG4Lb3Dc5YCtAzVuPOWJ7NjPZiFl
n/XjmacFw/Cb8z/KRUKDAWhZqQQIHYuyXMB/N9RqPkwkr9osZ73LwL5EK00wOnIe
4IL5euc0A4EAdGY2eELHMPCa8jxQNg4zg8aWOqcwC8iihv7Hw/cTEnP364k39Z84
vkMa0BZ4414B5tk7G1OeF04HQI5HUAC/dVV20784beNg5Jql0f7hnXrcKz7n4Sgf
MX6SO+7A5gTkPfb+F+x+wq5O36rArl02N7oRoSuC+FwtInbOx9rEDqQFkZQQm9WK
CMm7W4rC+sDrH1UIm0TX8OLm0WzFHXD4wdi/2Y45eWQV7e+lam8MdJxKmY4T0FEM
ZT2yvxKUsYhMBcjAYS8yk3/t0jsZ6u9PQBeP+ghBhNktDhqpDUKuSrUAbPv9EtSX
TnD67hPI4z6bhmjItMJ606ObrNCtcct1dx7iT/8Z4gm8/H5SkRip9gxtZRSNKbhq
uC9OUuhBDI8zEUdlo0+nDXK+O9PT887Ao0P9FBOua4ZG2ni/JKvSc8ZzoL8EpytZ
lIPXSmHPkGk1Ui63SfOxuRKyjkYkZ8VdqV6PI7QVEPysRvvLLWN8XYi3rwZ0WEhH
1c0k+PqZR8VHFph+V0IZ37Q+r06BN3ihDB0lrAjtFM1lYMKhPSRaAlz2+FxQfGKB
d960ydUiyalOqX8mHpLo8X38WA0ncDeyOAzCBui1aj+jM3Or6agt4aWlzY5LTlsX
Mg8Lp8UHp6gfNfEmafoZMsjlYjJRF6m3hmvTYJhuFI4jxgktD6a2b+idg7LEdfjU
AAKhlzjcZQtB7qSwXB0WKZrIDFrBzVMD5DH+gcXjYXkwvpc9eiiH6SW0sIwralXw
Las1AxA1EwnLggntLGDYLUCGVria0ubXC/aImq9Rl9vNGkPsjl1P7hG5/lEGqyyD
x3G9ZXtRnYwzZmdllCPbtAjsMR1ceAFGrs2GmI5krpzWMABdssGfRp23Y4yyVUea
OwkiH/ZBSpydQXjrNMfNie0842SfEYFGopMjTIJFOQuozZf4NlyYRbULFc73XSBI
hV9ea4EAXXPh9pSPDFkEPuJpp8jDsjUONq+gh1HeK1tiq0dGt9Yn9B0OhWzP+SbW
QbEhF7Mybvn0TUtOhcW47JK0u+Lt6gJKVXqwty6UAnbqSR5Ve89XePcJW6ock1KY
b/d/BKytpwZdbMILkuZUwJdBVddC1gQn5Hn3IafGLoiZDWO+E1kEMfzX9EI+XC4R
GKK7XU41rPza74tpllYfuUXm5SX5WW2aqnvPoitUcB1xqNNBmAlufLMR61H7hxoc
NCDXs89QCmqr/rUDwMeOKKZI1A4NFUV/Vqf4MWEbZDuWuS2qU+0OMU0ja/tppQHj
MMT3NMl5f5cAqpUi13WxfsNtGxgQwbzdBgPaypScCC3f2htjKBv3v40FHudS+ias
kr/GecGDlXjfJTlxDyK6xjJGQQSY7+cKxv9PP8Kf+JDQGm3yxhnPgQ984QaKE4AX
9NFcS2F18eMQ7/1t1o/1FiGWY0ZFXqU35gL1mI396DwA04n8Unln3a/aSL1Wm0mt
mABWJp0wkFmehFjqon2rCXt4T+9gjssgX6mM0kqJezg5AlaV+nsgksuxr+4oROTS
bifWEUZCv0ry1Klh78ZPnKIutnyahmbQJ8belXDHxX0C2GY0DIiUGEDfcTiACjkV
rMhplcXEBcqM4fIRzGg1UukD78o9+CGUJS0byf916OrIlLmSgtpoAZUc1pJrngBz
P8HPdLka4SCvheHt4x9wbhSgwUUVRfdS38MQqkdMWlK68APz8u5rV+Hf+FD7huks
K+BR7v5lgSS/35R4eEuCQjkWO+cQVVG9z6BdfoLoCbFad1RScU+81dEWsrO+D97g
P6IP+NaB//1Kyg/0ejYGggU1iqlFfqyDo6lCUllZe4J+cfi7O2D0L2j7Zjn5z3Er
ANj50ib3T3jhmTtUSigeqVbpdNV5FSQHrNDZZUaBin8Cm5aqmJldYvt2k0AtuTbB
rjueOH5HRy//mJI9b/1pApcXNefc+TA+WnZnqQO3sujF+WuIAtyIEZhfqGbrTYvX
uyGxTBCIG4bTIoihgk8zvKOiv2Sye9v4U7V1PnN+0hnDPKq/xpXEk56t0d4fGxzF
ZO3LAmrOZBuJJD/mY1F7nKKs3bnCq692z9yuZpyCERof4U0DHMAnzj739T4YkkAL
OQ2j4R+/YsfjQsWwnUDMNBiZfgtnD1SDuMxOiDxwMCYIonKp8ZwqKv7ijuBwu9R3
XjfcQjIzKdiEk6b1TwG13EU219VJoJbLUhYHLA7QyharwCJjfzMXdL/3FI0HTwd7
8F+JHOoTr+5UhCEGnyzCIlM6zPIbhlLxwpoZddA0vSrcCLXPzI43oQO96b3Hzdba
KdPvfPKLSHAaRLESP1Bw1STIb56PCYrpB6juqKhphrHdlugvRdKNhETQWohohqft
Pv/bReObt5O+mPSnblOwt2vFc8j4RPX2ifC0TjvZLTyDR7i6GHEwd9/wBIS8utEo
WLA6yxD1MxDe2B5or+u+VD6PWuHqGIbzLG9jVZTyOUgGIKDJCCoBKjW5/ArtRSQ1
Lhg63zupR2dtyGnpgCdngl2gwT50JcFCIfLXLCXjNjC97RjJlfYqGvVaQFE7JCb7
um43j24CfHHBkgxZYvAAe++obIEaeaHDIpa4t/ftHaUl6ciXukZ1GpSW8+CIoz00
vSo1COFdsVFLn+7bVwxnRSJcrE6ngvndPnod7FakWnbMZo56l7SEXMBZUFIIG1hu
6D7tUxCXQMH9a4sh5eMkBM4/YVjOxaVEAcaYAz2eAskiOr8da0B2IYTln5uez0J0
INGJ3F+HR4H2lsFbPrbAoHIxiJc2ghfxEenZITrhB+EWp6JO1wOJaLXyq2HGna7C
FCYQdB3KRdYdQ1ePcj0O7BsTe1Q+4AcymWZ6lUUMD2I99fiJhBAMvwJ+E0MW4Bqq
VAWSnyNwwuizruYn6dHAVsYEEr55MZEVlziV3A8YTUalpmWO+6BGtBlDcClM951D
hRXNIAY/JxxGvlw1UivT1Ve0iCIbZEEj7PJi4ApiSPruG8b+dygFdL824BBYkn94
0XIU6A7iCrGnjCcmxxVqMBfatKGKSZBIT+oMQOiVbjm/Si8IJ+FfUFF04PfQX4Mw
+Z/i+Y8btXEYOUFy3dq+/tNo0lnzavkz6vhNy5KVs0d5iEhHoBNreImZOFIFmOmS
6eFzr1L7cxYCVUUVwwJPhp86b16TO7p3wjR950ehpuKfgVoTXrcNoRlZcWIvXUZ3
HRPH4HUIgOQh3oYSpp3XhHYhwBa0Wh4tQqUlwwjZAOC5Zv0YDP7EdbJnrL96KGk6
KweDXA0zg3h69Whff0rEBc7Xspzkn+khpyD1u9Suht8UliMDBjd5LJ7X8U2OpeUC
G/ga7UbAT5+D2DMqqQEOq9gzYXhClyfWbeRaA3hSctqYkVBzJcKnBhS5eVYIJC9W
V8qzSfiLc+vTcGdoZYVAt/gUPsrXwpS9mk+CEX8DSuTM/y0y3E9FwDxUS1uRGr2V
cwOMPrA6t7yDxVlOaR7MnaEs1iova2NY/Y52SPdBWyrIh/duTDB5HTs6UWGLz5V1
mCrhxRqrAzYA4jafdZzYEoN/uXApb8iwEHHNENL6h1DgiJFUn3nUs6L8stHVvvRH
yHTlj4T/Bq5Hf8ixwAzjVtxiPnJdPo949n7Uj0B+N7S4CTcwkAwxsanIcfoXMyCT
KgJelzp4Xn2sy34rS1pIu0z0nqxqKW3hBDhoUGSDwXUZr0U9JG5G9oQ3bqwQe4CE
ty6zYWVuQkd836CIg1Ye+hr1o5OV2kFtRn35GNmwjiP/pVuxI34rJF6x8W4wdITm
FkhvC8ur8P1TxNBGhbut8oqno1i+OzDZh4EuKMQrjLFYFdYaO6t8R1enuWAz4dpJ
/5QzFKXC580jQJzsQUMYtrP6LQXarVSCrAMr66jkwI4Sg996L/2qMA8kmnn/zGUd
dV/YP0iA23/tQYS5ZsktSaScmXN+M/KGjgjjSLdv9fPg+b9593krGEC19A/faDcS
X8spP9xvjDF6UUBeuHI8Nc1Xd15jzu+VUfT/bMH7zINeEpesGa/CygHFzV4rHGwu
oCZB6f3NUFkf20xq27z80wwNt6/hPv/dZdj+SgBwgbV5C+IN6AyCYopGsX+B0l9M
PYQFB1gqwMfxZsBBz47TLs+wYWuSa0qgknadVPuhWrbE26PD5dlYGnag/nylqYs8
kJsP4Hn3uX78rq/UyCkh+m1MVfu28xe7A+a/jsAkFfsMynxlK6q6Nq39VF3MaTyn
xifNKWNHKa8XdwM2GN24rFaNMuqoCjaRrxcJ0ew7Ugd+Hl0BfijqpFwG80dxWXff
NYQqpHnE3hzbizz1Ngtred2Mki8v8mQwdYCC9Y12MnDa89/hZWA6u72kigHcxMIE
Ts4ju5qdNFQfbuOA1lpqeZe0Nbm3LZOMAw7LGak6nuwXvvTbcV/o24aPQ28f8KV9
zjd14h6WwAUWyw9W1Qsp04+kCfw3iPHvTgRypRLLxmg8ZeuCQu7HbJPE5Gid+SD6
SmwrsHi0lrIshRi02CWNbkLyTxCLFUoOwhphh3dkJTQOVWO6j3aLAwQKtOkH5UqA
keK28yUuzKE2ycjiDCkkZHIMbrw5uwKt2oLB4PQ8gzJm3K0s54sboqCSAGfm4qcf
hpzAkxp4y5T3LSr/N4KkXg9t7XNOwupau4p31ISLFPY9J+Z1ypqPA4d4UitVPH62
23pvEt9pGLikk5ACzVPCj1ZyGoWpEq0aDJcnUAfxU7adjw4dSAW0iJEWfzHlKaFy
+4Uw9m584YcI0V3YOxQpojk+mzqRKGd4izctMq+pepO7qr53deEpM7YP+b7/LHk5
Wg2sUQ9aDGZuMjziJq4rzI+Uu0BnoII6M3OlwKaYk7dJ7INkwvRWENXmL4RJ2kX3
AX4uYDqvM8Aa0WGkfgZhxZkPMEx4SA7hw27V0uLzXOOKQabSbsfCpodD0TAxYjBj
4Gg2O1f3wdTEskr4ZRh3UL3N32HQiK/fHGxbWgDjgJJMnopRyOKzgNIpej1QANDB
95ux2vZknzA9hodEAFxaWCvIfJ+AywZZFazbQfW+vJpOH7EHDFjIwYYAQvUr+m13
Vs/kjJ44A0BDMnq3IA85cd095XIem6JYPbBr+5tB44ox0ilFrlmbcGmUN+mzsOLA
FnW/o5lMYi3uFH6tHh95mrEC3lIYExfRl0Zw5oxOJbG6ghUw8Gr10pU+WLGfKPIl
VlPmOAGTpRs5JCLVE8xBJuuqJxpGET7EO7SuF1vDWjUAjXep0BlcrAzDsqc4DeBa
ou77h8qc0xOOK3i1OAlOG6i9VZ/t4wKnvlsEdiFSH4XiwUkQn5jSDKJzH9KVCnrk
UgunyxjdVXoV3W4ICz/XLlm3ACsQoQB4NCjxwAhRCX7p/kY3TAxnwATJcrh2n/TJ
6se6AWBSb5hCzQ5pEnB/UhfFA8U/Z4zRX8B0EEpSpRxJR5PUmYOQ5kqJ7BW6G/Az
QOoXcSkpDNb/tq9Z5+IQyJixrUzRmGYmwTdOc937QUp/bLD3fMwWTdYcjfVocsZn
PCo5Ps51CMFBDj75sRW5CA1cYKWQzK0R2tSlEg78tM5zbckaelCGwa+13Z1nvU6V
jRJ5SGAmi/03suBnzJ8jaUJSS0JyZtPjhUZdaCBNuQE2o/EWFyD6XR+EzI1g2XcB
j/SUcqDgGHQ2nbYQxECBa4mFJUZKXypzkZhx4Q5OOJBHnqzHInKoeTWG5Xn6h5GQ
gX4sf4FfWAcs53PCvPAwh5pbCqs+G6Y73hMMjqaUaDCx5GqT3bGW0WmF35Ii55Ab
+qcbWhU6d2geVveS9m5Zd2vJsS3KK3rzVBldBe/GCXv4Tn+QktF9URXMHwks4l1S
2x5fNN7qO+PGph9I5sCXxK4HlHfWDMwyIZazs0fTLjag3c4GCmpGXqYPFjRiwP1f
aMcAVF56XNW3KSm+WhzP3AOSPDbZmuUMFATL74lTV0eT45C8qoF5d0Q7czcu7srR
39/SG2ltD+XcdxALCunIiKyocrn//lDo0YKyQf89CYGznCHoNQqF1I/Db+OeW+W7
cIXEIAYyWSqsiaCUu9Om+zU6xYqed8sWV1gnYGDeOhZIO7ro/ScZBEk7gjOcode6
Wp+O8nSyldP9nuN9C8VPDtnDrgHU+ReemdpyMrSShfhjY1qezo6kDsFH5/kaocur
cmIQ8NQ/HgGJk1aWsP+XLBwIoZuJKAYdkRDLZJS58jVh+Ln7xgS2LPUQo8U+rHmS
JRAVO/xyF4gMaFV68/k0hPbWiBccv60zdlDwj+XQnqgR5pMnx9GyWpHp7KKQUOsm
xuJiY2kAtstSzcCIQnlujNBqbyOvA6vlpM7oOXutqYITqz/4CeosPbQTU9LYFJtK
CaDLIwd/5dwEKeHtGQ5r97cDWUSkfadbNYB4MPcEvFEl+M5oC70C8VNYbl6oOY3B
77MdHCHMI0aCodaL3VUATQ6MB5DwY6trYqC5i8njdj+laT2bGrzx+/W7wWvtTFDt
raxLxkBb2aFqq1b+gicfqT0kvswpM+0qy06v8P9/72Gk3misUxYipUtkYJZ/xtTt
pF1m0YEr1pfAc+KLmejrUq4fMjnYRjFeYNTG6KNyKMiNheq5JLgQhl3cElwdqCUv
mRU27D5P/bHlwFkNCXl+a1nrTvd0gC4ao5sVtcRaw91aj4Y4ESQ5As37HkOOHS85
7rpsHpSf4/7WzfzwNywXA7nbmpWbeaj7hHqVghbZ8VpO9sHQEuKkjcJczbtZI8zq
/9n3p+Y5vJ9ISs9lCaXA2WRX1uGheTg8UFrZ++6ie26qLeC69jg5qlkl+xAFy2Mi
RbqwYeiNAFhrCIt6QwRZDjM4cNGj9gE8uiz2dl2qxGIhTWYFme4ypu04MmSTgfZb
DT+WQlYWXdxrxyoVAHrndrmVsghuaMMHS2ethNRkXZe+L8/iIXf+w/RvsLPFoLtq
B1rQx6du6ff8A7wrOvVPyCKPAhYyRnl4xqwXNdQLUHN+xt1sEchweXoIu4Z3jp8G
af/G57nbcjNfBmkoWmyjNFMZATxQH3KUoyVMF/ztKUpnT0XmAE+A3RGjbnLiqpYJ
Ge1UdyTVBah+S9nBO5xskMA6Jibr9GVeXi+I4SFebfUO2Kri3xJ9OePaCYZhcRrr
9G/P52gUX2ZFuso1MHooriv29wvRDP7IuIV1oraLGRx8eVrL48KdIoNRb05a7Lcw
ec/6uQ3xmpi5AaiYm0KBfkOrA1BubX9wFSsmGQCvx6WCT/9S+o9P4E3OB8c8HPS0
jGLuRlmJSy6JWGfwGFzVaxuEbpOBFWvmYta4WQrkDqn7Rv7olTFVqq3lH18d8zD8
LF4QQS4/YDWbIQh+LgJvTXXOx/95ezJ6zKTX54pGOJO/37TBH7lPaO4PhEsOVFA+
tSGS6rGZCsiqW34ls8zqRbBUdNvjCpWYmlHnsBBKAF5mdHpT2qrDlSLZHzN/02Iy
Zf4C4JiGhaYfYni/pxLnMCHzI5QKjGvyxUQ2am/97KOCaUeQXxArQredOyKV84DC
2opwLuB6G5wGVjyiPCa92wgrujitdT6e1FT3Eg9uuXioNw7LlKJ8Q824o2q8PLYc
YJt698G97I2rQSVOR4PgCpDmeiV04nxqFvdluJHXvQ6x9ZkEnjzkspxcuUVM6NJw
IlK8yMhkly5PlZ5t+dQblS01feFMyflnh9hrJhQLJbmM1b9eneFIiZWJeMIY0C/y
qZDeg82mjlUwujzTGXLgHNuMosxrS70Nwy1TGSKj7juVG76e5i6Hlc+ITUx8zJ5u
F3WUhQhzCiooEgNxy+lQNz/H2pzf3+iRlRDN/RCPoNgHcW7qY3reK8vtsQIKB4/v
vd0MEQGpOK4BPY2hc49cH9gU+xm+PtBLcdt8lpeYeXE4jMYyTMCWm649eLXGOjz6
/PkJ4fZ8SUiFlTlleQawfCcB//Ze4lBnQ377FhAKe2pqFM1/j/Y+3pqqUY4GhTf3
jVl5lB3Qb3n+DLWu4QCnaNcSSXjJpLg5lqcSLssRtTQ54Ix5351Kt4GuPsNnb68A
cql/+4vaof70o2OjpNWY9WUS3V+ZAV7tiAJhSw9kKcdTePFCEGvO4LXL88CA1HvV
EjWSu+1p3vHJcIaOGKMUopJLdPOwpQ4o9rkrft/gewtY9Yx4jot1B3teRVTv7XZc
Eh33LXwAc76Gi4xEgJ37t7ZfqeKtLgOHflbAHnM5orwN0fWfsmNSpBDOFxufoH2H
wfQpNU0rKeie4WzhqvkqE97XHJEz3RFuucZDVp/m3Vky7j7ataf87LUFPSX0QHzh
9hWRQXsCDfGv78EAhpgC09zNFG8i+vdCIi6N890bdUHjW+2rkkqvyMzVsy8x1vMW
LFFlEfbFhgQz98sTrl/gLaqYfY7xZ8wbUoCqNziNYskv/Be3ciapCHRXlw/6xoeM
ki+aBVERplZPHVji5j+TjgYxVjlv2bMozEdAcDVoMYU5Ql51B0QIDQcNtofeqe7H
EdArkP4hj+JqCljR3Knf4qn/Mh8igimwGCUHAuiXEDmunSTLsbAGJDI06Ora9EbT
BA9bEEPVdApNgTH7VAnYHRzWiSEObCi9h8ZHMSQORms24SMcZ0jX2T2pOk1bFHtm
nVzldDVSXHLyi1Mu+Nl2o7oimBZjz1SGI9FUHVvbpajqhV5Dhiqfei83v8kM26uU
T8BkNSzD/PCAovaSZbsPqJmJR0kVP4PmPAWZOM8eWOxMkxlXTRbV12BeK/5fqKyx
d0osdqbPgT/ve9HUo0bPsu/HSh+0dzwmTp88gs9v4TSBdwoLv0+iI72xO7CPQdD7
soUWeXikzNgwIN25a9DlaREvOYG1a2KhijmjGPm4sQ6xsrLOWriwIWi8fXVGSsxY
5D1y1vq0wOhfA4FmKonbTAhvIi1OY+V1do4kbMrWPpzOhm+PwlOE8uX1AGeEAmqJ
cDPb9axuOHzIN3j+HVHwANAqWFPauY8LIjugby/wZrlrISkUcOOOm0hsNgJ6qDbW
CGqDbH37bH4099z5NdwscNv1rXe0BI18l5CF+/sckYyDEpNvn3RQZxbfUlGvr6nW
N4Plk6u6t4iOjIdu3gch1mAq4C/wTzdtlqkNkXHR14LAdsnWsx6dsOYMQ13KUeD8
0rpPrRCLdQHHfFKwVo9GUU2LP1V7s0eZOoxN8ziiJltC+116Ms0cdebq0oM7doaY
JS//Ez3k4U8cueSObTiwJ2CqbAwn2CMX17W03W80HH4NnebPWnQoV5mgCiX8xGSt
tEkrA8ffIORTvWwLjEqsYGVRAYnrQTg05unDkU+LvcRzAg1040QtJUFMvHRF6pi0
/K0KoWNalJGxvBMfPEqmfOZ0xEaVjeiVJYemW/+ZpmpULSHKuIIDrSTtYAAk/SwK
G1OEoyeH8GxTmE6FQ01dVLniwtEBGS6T7sv1j9ToT26YRkJ3N6vaJKhqq7k7PMbc
P7GZ8C4K9UxtEAqNBi4vmEvnQCI5YkWVdEKD8SHoAv9peSFwV+RoEzBfxzsRdjqT
kerSOjA0g82OjOzi8dWTd+3Dh95EG0B/qfrtMGfLoJGm5OWR9IiqEza7Ufv4AzJP
PC8FiUJkiIOOaHJyiUt7p5kwONP6Ays20Ee1YrodjcXd94L47TfWLJ5mqlEN44wa
vVnIAaYlCwPsrFPq+iwHwyRfciLMTLDnbXyBpRUz7yuE/ytbGU2jI2EwmJ589DE4
kfvl7+PI4oQwbOEwFM84d6rPntVxZljQTj34O5WwrBcEorvk3lFCEnI1MtusYvA0
+j8s8NZGw70zE6vDQjjjF/ArsO1UOwofQKR9YDNG19vUm5xLDP/1KGodU7ZVpU26
DBW2qRAmc4U6Xl2a8cu08jey9sB19b9+X2nj/Y1TJUE6Kd22KnG4pWz4BytVmWMR
Z4EajYsmw3wylNMSPrdkXlZ4bpcy0CO0pnM9fx0GtJeOQ+YQM5o034N1DNV3H3N0
LHSx1djlu//5cnT3eCKSi0c/XA9s2WKiIh/osoh+fw92DmrQ1wMDsO5Qt2zeU7bh
QDy+owutp5H5DGL4E1siFXwst6udJA6w7aOwHVQHdxxF6PcCooOezj8GYNteAxvg
AEnviS7ckkVMikwNc5brRQsmNIYuEQC5dBGkM2NhkJyWI2g6exAXir+pQAYPK2ZR
3RfY7PtDvOd+3pzzYu/MnExJyvalCuhJWA8VehmHWfNOKx0yQHJe/OqlJF8xGSjH
4wv2lGi3l3tuxxnVRhuM9PtIDp/Hs8sACkxlw2Vow7Z/l34wxw09WeWEKBYyz0wq
lo8H+nDkGWcX4Mf0cdb+weLwSut4i2BE84vUdBxk4sHFa4EQGcCtkIZAKtvsEKuC
F1x6xXRT3ZSZGprB7dlg3G2SCh0pmZGTOvYJlcWL2sZLjsIurtAtiuK306zN+cNX
DO805V6YUPafjMzHT/MMfhFpyX6weZvVTHvTobyg4TFDLaaoXqzMf4A0P/fcUWJF
YbRacboTRH3MkC1XDA4M3ulqW2vtdFfM/PbOG4ulaPN81dRfl48zGJHhZU5u5IY+
SVNEIGAwzyStzVgO2hVrBF2//OevveLMBDzCelKUGxwQLaU4auamsNgPnPX2/O89
sdOY8esvpa0jrp5U3RDSA344rWTyxPvxQOBY3YoU4dhggO7WoW83wYo97I05UpDz
g/ME/jwPbOVqSqLfNCFM3iwy3c04kJXGUHw6AQi+yJCXDd7rIIJQGiBBD20tlDK4
yw/H/N0hlvDjJgeo8czKYsCtwhx+gMZRlaohlSwv94vhXCyUuC4zLZdIJfxhrby3
IX2Uf+LGwTEWyRxkjmCDFFQFdrKAdkAiHdKXQwUYW3h/O65rm0FfotWMYMq0HVNV
BRhfN/5deHXXxa8TBtKUvsCQcwjrPIu9l77cvrRyFo70iCFr/oEo2vcQQnMg5Gm6
zae5/mj9YxFEQsLmQqls84/qldWbRivjq44eSCrqQuk7w5N8caXsW3CAzMnQvcxN
E18Tc1x/CGiUJzqDawmyfyOA9S+aeH+clC3Ek4KOi+GaewX+ZW0UqOqdHDsBxag6
mkm+iOryjZNanYlDF1jsqjYk6Zj22uPGJbi4n8OBH+OzDYZih/lTwC0yF/gV23Er
hMOGMxI6RfswpKkXKxpCCVEdPW7fdMBHTKdsJuGlezzhpqKwSlWprLbLHYXJIWxK
sEjcGAVgpJJ31ZTmY/4iRomuFUSHfpD5PHicUuu60nvPq/pyn2O4zkTpOZwTAV8n
u0xqAI4ez6akKGAR4Rke7Dr6JHafCiEyxHGTJ9fVXEd7DzZN6o4qpfq9XEKOpOk/
HJT74NTNBtgXSm0MAww8N0TnvJjE25hx3rIDTNYW0j9kQN8fIsUy/cqLs8Ap/hgx
vp7o6k72tLppK5CQT5Jn11ZsTgIiKuiV6G0AUiMNptrJqrqx+5t8k5aVUv5tlj8h
w+jkvJKTR41za9aXjAlGwFQ+TTbMf69H7Dy1L8BvZyf1/sWZV5ythUKsp12uU4pC
KWEAIt4kPmHIoAkTcKmsy5+IXG2GJfItNBR9499vX9Uw/oB1V63bfN9r3b16pf8Y
noXmlsE/od5VGuMeXs/1rnf52pGZ4/z3Fkdy1oYwTXxmvMFG/McTe3U8qgyHJ/uj
G3DUENjZofSggqhng8w6f7riKhp6JdnFx4nsP9zDcUUp9dq/o4x1JGZtGJMiSCP9
j8DZE7HEc3GXkIBH1YNej0j8wjEaAG0aU19DM8wSUPKwrytrnL86BhyUruSbvZQz
XSm9pdXKSbvozhywYpyPWNKn97yjwoCRZHB4X6tOmbxS0sKH7Kn8PBOf4M7AmCUh
NE0hVN8bfHoUgTmlpXyD4n9k6CDFnzPmKZehOR9CbDaDF0inJeq2A2m72cvYTuuR
h6XkUlPOgM4XiT/nVZmHYiDLTPROl0j7BUHXVggNmCheQa/i80Z27VypHy8H9wrS
iLnYGYpEaban6IDKq55ajsrgPrhR1f9zFdlarImhtyaC+JKS2YpM+4UgtNZzoeSC
FZdkDh4pk5831eCDRO++nUUiPqo2PCyvdzi4jBwDL/RCfEN6h3A8lYvq3MkpnrGP
83YBWT0BxnFvw5JJvTeVOnDZk3hTYiVUvq5e4RrWAwvWtz6C26F4OK2kd23SPTn/
fKqD2yc37a2wg4BShehiOFRW6b6kePpU9JIh3LYQgexz1vIlVYnjtfbbIC/FR3ms
AM/xpHr9gEJfONsDpW+2goOrw7r3q/Xrv2TBez3Q01gUjwRbCOdOegI8mrp3SZ05
IXBSqCvgi18BCUa3aQ9FttKp3I37x+/n/GjIe0XO03G0JgoHMVTOA7HHEhDF7/hJ
fbL2cVd1eRTe9pAKOZc+TGiWW3DNeLDrueTf+1wgl6KXL4DUQNBzPtxOTdGLc6fh
70UhaVC9FGh+cEPKxvIUlUCqM7s0/uqoxEOJZgUgm8xM7FRVHKkuPZsCbzaIoEky
OItNp27H3Qk0kFmtilmReWvlUZwEqE/1bKuol5/Yp5fduL8lv7gduNAa5OhlK0aw
x+KP3Eh1BIp67s0HGakZj10c/8ym2mGni7HnsLfKyijKbAJ3CFziaz1JoJlt66jP
CLZxh1QO/EGJDkZeekmCAiOYQ6Umm9JgYEM9XVwGRiyq6U3aXgTsQ3aMdZyCjDUH
aXdkre6XT0M2hCuzDdjdqUsOt1a9AYvTWi4Jvpv1aNR/Q1QYuqKxXsntWxgWfJrW
EsmcyV8d+RmY4/bai6iSdQmpgkwrutoEBBrYY7uRuHTJW+JHMUcpu/BmZYRtkvhX
TYIuDsA3v1VTGNbyuXCLiWiP9C4JU0VYEQ/iDh5/zxF9lCl53HSxQcUrEZjeSdQ5
YylIqBVmeUlxfE4/6dyhyii8HQRUo770AtcrAxMEFIZcVU1NgQQnsqMQoUV8Y2cz
z9SkbQ8b27HgFiDzYFaw+2Uw30iIKaC4FIDmstFYEGFQVVv9r/0VOwU6zxyGvo0x
5OPOwYZPCAXnl/iVVPO4pruDfNqWh+IrnW6JtLAw/GcI6DA2UX477D5nVdCjUr87
hDyA6S3z486cMUCJsoQu+lQHeJZIB9/HKX8ZOk9jexXEjMmeicNfpnu5+OmWp1BI
w/vQeVl31Fzf9GVOUIB1yRst5MyN57Im+AZetfWtX3PeFPnjsyw3zbVC6ANUwFMl
CNX36cIU81oWJYbPKWWkfFEn7UtTwlctxrDH6JCMSfGLIbe5QX4IUJqLv2JcfY1i
1Ospe0qw+u/3qoJ03ag+7MjhNo7opVkegHF+Luz1DlYPhXlNrBxtxjKi78erA8oy
xVKUlHMf52F0E675UeldOAJCpFkl+ay/NFdgmwW8ezuUDgD4IqdhPHETaWz69DKC
bOGnlBo9vX9TM/q5j/dKOsQ9pGI2sJAsGtxqFZzkIkrnrmpSN1LKL+QGpOu0qabc
Xy8nMAoJABLgReIgD+vR2xU0CUBOkP/LbsETTQcUtW6v8xiL55CHTjuynEq31AEW
/UW9HShxhrIs7V+oSCP+UqEua+kkYuLedT7JnW4LA1KArdubi8ZK14S9BByluTeT
stJHTmpzhHsBOo01DRPPQMF/0/8LQz0hA1JwUuKg5Jwo2Y59s+459OFMh2GzDU9W
McTrITrTz9qtH6MaA7xtvfsQcvqBOy2u2nkz5j2AVKXLhzsJkVMsq65g/z6ny1rj
WLawOcxYm+ERcAJiz+whcyHMC5nunqo0qP0/4oU1SdxOAr3ZwN8dAiSeRT2c6sRd
vSJdPJDFnsfZz3sUGy8ZMznL6bn563F8kRnYebHoQ8cH5QlfZbsX4n4/6xvt/ShN
q2VphmZTIaPVvjQJ5FpWMrLwf4pRH63y0z6I6ShqrKeqrgeRhPTAIgH39juVTqqJ
sG08kllHOYwHV6w2VTueoTR78y4WReZzmde97yfR7jcr71IRyfalVZiWSEPl0/xX
FN+RMwKouKZ7zWs3gfC/J7QArUSN+sGRHMWJEt0q1fUvJs2oqQOIYakefo9zs7vx
L7ilEymGN+qXHw49rvmleSF3Gx922po1ALbMqyCUbirt2qMYxReVq83kl+QGWhtZ
k0h8lzpOhGfa7wnjmIcykqU8qBecJJjONz5XpznIgZ4uI91yGn39xlO80tVPY80d
H913NkptwO1dgH10tRVS+exdZZoYhInX7Bf/4+5yij2wgWZnXuMjXAfq/bUSOxqC
Y0m8N1g+Af88ReEgcFoPJh4Pg4QaPwpwL8PseDzfnxE1iGzZY4N0MoiRLN2qg5ss
xB2HIeEEqqOL/iKDCyaCW6ImybHPcHpcApIfQg/emqWipH/PakMPQuVFf0mHgwMy
1Tdi7z16+mIdO85RsgWvxjkwe3yxbhffOWBmfw7F8d9Ueh/uzMeQ53oJjWUzlDuk
LB+jx+fpmweYQKj8rD8GVG6HYpjKSkc99LdCKmnTIuwBWZXLblexTeHutlVMddzF
bqGI0/qsCKQwTJfBt2Unfl4sgR06E46F3tIO0Iom6iVUOw7fRLHrNoDy28YFuBFv
mJOoNFh3l8Kc0n+974vqtJ+zyFxhkP1vLJhkIJJwvGTwijri2KfjxlHazBoCd9We
oMXjeVpyJBMmK2urLwHulkmZ5snmtKGjua6n10qqQLOD0XH/PypAKZkPcC/9PUcL
safHlk6T/H/bLtGBXLksJdCEGHlYLTl2TCbg1gPwqNpufYU1BuquwW+DvqNvPvFn
QugVY9IXaskjJNzeYvOOXYO+tTMqI+dXglGoIhC23BSEoFxZs9VI8S4Y5m46K1kS
w7vWGo7s5dTDlDk3WmsDmRmXug7KHX7he29Tn0WHB09XvlIV7lqAw6xu4ZtjFZPh
6pjdszBAsfiLs2AMT0l/0AWbCDSSiSHfJW/zgTUi0XBgdndHZWo9dFm591z8+zLl
y2xUxLn4j4hd0cpb88Uze7mDOHDMaVvoQ8X7TtOe8SIy+72Q/6Hl059780b3iMfE
8cj+hhkxtZdHKFvHe/lC+j8SqETap6bPxNVI5S06Glj8ufUnNedGwFFUbW99ycbt
BaMT7swPUfuG89jS9qmQL2JhjJnJjcOxLcoCVqiUHU9MplVUBpkTxYteNife6Mom
zizMEvy9Yhnn+zqHKPluvI4v5T7gLDXW0TC6io2CKLulEVva0abrNuQccjSv86Hf
kn89MoF8UuVv6bbmDnJxVDYGEPyFiTd/sf6EoIA4xpTxeYRIWrcYTkGCIa51HV+D
2IUyz/IDnI7RT+tQZtiT2awEKJ3Ld3XOOzCm+rigbLRPNr6JwAoXYOdK1FMy70Uz
sL89/6kXRNfGl1UOGveqbxO1OkZwS6vZuttO+QARHHZKyvnD728w46BSYl5XvFQK
Gjojh/7EOTlIi61W9Nbr9P93KzEkK8ENOqoh/WJBToFqT4XRAEzfASaSPsJPHSI8
2CJn230iO+8N9NjjigG+UkM67THk1bvTCh7xHpy1uL46HSpKIgfmdIt2fQrmyK/B
U6YPU2Er01l4XX8AJSglta1UJE8uX6hRqFA/aAMQLIKiVbCcQ6OIKXT3nHs2bflJ
YaZD6z2lnAW7gBd0ttaiCD/fR3FK5t3gNEUF5ri5ZDfgOmOBrVinHwTShjqsDICK
43+UQUdwXp4U8jHWekdyulg4ubA2kO0uKo40Qb+4OtBtbPAXxyJvn5J2Tcc+peF6
4aTjf0lw8dtc3sGsybufqoqjtQFqQ7FhM1iID9X0plX6t+4gZmnqBfisA4AjiSe8
FP5ysVtD2AxA1Ysqz28oijWY1FhuOIrfY/A14fhnJi5rfMkQ72G+He8exqgkVHgi
xkJHu9zFCr5mxA2SNHyfMif7aiuRzzwCSKw01tmHq5F+Nf9D1w16cdaekdXm7Vt4
H6QAw0mAw01jC93thfVPfTxHSaU2O+7ChuBzDYTULhNcN4mLcL3bpEPZoKn3zLr0
xadpS1BsE2MhBNZ+CPWwox6t+oZv/Ql1MceDgMjPNNTyY4lhuMbN1JAiY2mRin8H
7jWby0YvS2GFUDDGWq+DbrfQNA2pEc+P2O2oThbkP/SQvd8tHhmQjEnmC6y/h7Zy
2/nQdXk4YqFjjSOFxj/vzRSqNOkzoCkYb3Oa78pSu5ED4Yn2KP+D3esqDjRA3Xi0
rVcN0yaWaQcLNT1hVy2djd15cdLWmQojEmmZlhlDLAx12n/UXfldfphNiYDHFwJG
WWinftA6ImLcQzp6Uf3P3WeNZVXr+vX99Wb8m7EsqKj/+QSs7PyE3xKn5lACIlco
XF26wnMtQHtbYQKbf1jw41MHK/lv8FmXdBMc3SViEAaC3duzZFCIK66HJDssriAY
+ArgBtlHUXV/3qBBWE7+HdK8hJWMYFHNkSJZBzol4VHE/ozn+55JdREPyx8C+qP/
pH4Yo2FT7LnspsfS0OL3XEVAForOc5o1tUcFA/COyPD8Zrhm+yPc8y4eGBcS5Tc0
gwqvIAUvDvi8rZ8+7nDNCRIyoNX0/b0ZUOotqQq+SDyzzUBOdp8yzWwiXIe6+VHf
PS9n+uj+S852qMMZGY+BtoqhMAX/xMxyH7+WjvgFTbyHv40gfq7YYSo3+mCF+6yX
NHif6DQBTmvte3zGs0uNA+Itc6XJSai0bqSdQMFy/etPvyo87ryPVgLwrsf3uPtL
6m/gocetpRhmG6VHxlKvRqoEIW3ntq+BhyrX3vb0CxOVP2Baj6Qmuo/37a5/jRjD
rCtUMpQ24H3qV0O5MxaeiQrNpMH0JHKTlZuwTA1IvPEt5IYXBsaOyfv88IvC1MK8
tfD9/6a0H857SqoKK7L/riTLOtWgqTvQA0dbiRNneB2l84j2LaW0crf494w6Ho/i
XBpEVby5Wdhh+4xShwBJzc0f0ApEgHvviLEuh6iuCJBejCgx9v4zWCI5VB2wv8NV
NV118wWwUysqVitV4lr6puxgQMfu5bBpiM+uMRW9/qACx7azLM7LMOzYAz1WK/JW
x3J3FDefCEkXWdPFk57JLQuFWEGhNWWvY2FKn4QsXvAX/JLW0aQlwTwF1oxHP7LX
E7JYgxe9e7OlhQW4QmrBKZpMeUIFV6KzxFLt6nIvcMT7jcelpijXVOTlwBjppS3R
oMNW126+SvFCSlEhP9Gck+yOfE1ie5aymCs6nCl1ZT+vm55TaUf7ODG7b/+wE0So
wPWgtYmrivQY/zNirfxJwa81sLEQ0/YMawHW2+IqVn47mYzliMP2CYfC+ninMyqp
Lg/EPHzxeoO+iVvyfsduLch5tpBai0owKsJDqDCy/6O8r2HGqPgrQ8uZg+DpB+qN
YyYost0YRHlGz5px2v3unM2k4PIZR1QWfk4qOaRaFn0vOeoGMpuIUvqj7S45StbY
zrpcrDFUMcdEs5cQqxLIX+AwrSfAU+karsdLawLbfZq9waUPZcEdz+FV42dPZmmb
7V9o4XWefh0NkZmRtKR5e5mwENZCctcvIKw/WLt9FELPkJoCK4w1BRCHOzlBaLwi
opN7rVOlijF3lTO/m3cEePyGd3VznDW4uu6z/oK83a8bWqRH4URMr2fVoFzuRw+Z
AEuSLwDeAAi7sryf6/vsE+Z838npZGYybhKr8eEcoqMo5OhgQ85Y3ZzFUPK+AsYI
13oJN1XooTz/6jatEbz7DpbHdWnc+2NCoX64M9xmZ/5XgtIATk2TBM9DvyvdemGg
rY1i/XX8SgHyPqmLhzGxwDHe2zYwEbDBD/64Gm+LRcW7jGq/jxvQWoGRDimemXeP
T4cuDPztL7QV9+MikTiJAsYTx2V3SyRChg9Pj4BIwZNLz7kDjWQH3Uh9J0/GhxjN
X1vrqW9KbajoozzTai2Mlw==
`protect END_PROTECTED
