`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J2Q3aOgVNe7ZjR7p9FvGh+bm0T9fW9dNVxkdpYT1+3/KbCIY7J5T+oWtVBxQhXKl
UDa8Kf+XTaQPkV09IqGjVjnZgR6q/xD1oHtYguPVnI5ESECUj6bpz18eazsSoISd
IzNt7yH+wTeqOzXuYC2YFEzDXQChLxL9MwkDQxrK/unmHSVBuS9bMg9n42xZuRsv
g3e4bZ3CGFeBkjNizaTgdrLc9BuZV5OYFMfF8NpWb6Y8NFedzY49khAJOXUNPpr5
wOICF4TITWN0jtF7DiB8kQQ1OxVFAyHaAmcE96lyJ4Y5oNbJnJ2W9Uyt/HXp8Gwq
bOxxbeMjxOpDG+GK/sX/gphQ/SpEcL20p7loI++GYB0v6NYmkN2BJQq029Hd7U4c
n20EVdIMCDw2+9GkJy8HncfBSdzrgR4aPtMN9LVZrWUJ8kefV3ffqDX7ZcKahGHg
8xGfd7pp3+/4aAdrhEjdXshOESA20KO41cf5re/jh5LPiBAwbDrPdX+cA3IboS5H
`protect END_PROTECTED
