`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yTEuZatCgIEl/ewaclmzNRllmjUO2uHJ+gZEuCC20jNvXDVB9UQDBhJTNAJW7E2v
uzEHJAAOOrC/XsLj+v7B457r3n8ey2uihauGcoNfpETmmBq5zKun+lMdZ9BGsKch
W6BuJiOPTiw/zqRW/4iXP8Mt/8KbMTp3DxEqx1qYO2MG2Q22henx8G9ADXiC19UA
E3R8PuzpPWBlSdD2VWKmEW8Z2rzc4v1aoVKQw4mRM4FMZ68EExPi7os1hvejrVog
a9YnjNsjp8bfigQXPsHKC6x1f0UGiWycXRMPzveRg3w5dZQQxT16r2AoBBM5xI7w
j6wYx9bf2PZocdOzfx0VIU6nIZL4v3CiJ5nlFRrL/PfROIwPJTBcYdbjVZlr6x+c
eZ0C845gNJZp/3u6mF01tcpl1Bd6vhtmdzSFThOC8nc=
`protect END_PROTECTED
