`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
026nOwDsCW0qdAmOO9JxQByD88RGZa92Vc9FOjR3jsAwA25/EaZBGZQLk4ZT+IlH
9m9Lx4wB4U5are9mFZ6p88vs+IRXgRw+VRNY4PCgq/W0V5eFAaMWiPiULEZED5P2
zTuYzgKQjrReM9t2hN9ZPW3odUv0vsS5y05//HQa0bgKAtGucsv+xKwXALrV98Yw
EVJDZhjKIwvyxxS038C/gIrb5JSFOYsELo8qy/o7yvuGWAjpU/p400vJzB2cHYIh
ws8Z8AFUlcayzlHDVvCX0X46v7OoYbymXfeaSNP9vQdgCZY+q94vksdW7fRKwFFb
GGgAE8J6zFD/IeLEuypInZY7HfeneI11qjDx2wmF6KKRJUXDNjavaCYOakebAvMA
VbJba+sXl5tdMp0B4hvzeWbRzKmoCNB8fSw5GCiS1v0sBbaJ+8cA5A1W2j9JHhaR
7uks6SeftF8lOI2tsiWXzLtF6ZO6RdjteIw1OGiN1xuMogUn4Fbc3V76n02LzIPu
fDHshB6NgVf/GQ0dFCruPJt5wDfVnPqd++9zxGw3LFpRinEnYgFcgie+av3a1XAD
nyj+YR44g8pG8MGbViTqhwd1G10TF710eX5YKLrisgj1Sx04uqKQIXONecwdJtx1
1XZ6HXKZZGmZlYnTZMfD45lG9Y83SgmRnjImSg/738hnAVJFMAj7Mc0Kk76xR/sH
VpFJKvNWrsYSVRIOQEv4lqg6UsCaRQGdL397jJj7dS3mhbBraB5Vc/3gKsQhkH1Y
uW3vsJ/HkM6fDUnt2brhbBH3o7ORlM6PkZqA8m28Inh0Z3iS0S6NJiTtEnHdf/+s
axj6MeBD8Y4EI4pH1dF4v182KLPSNAKRxr+2jG8Ix+ZRwv3R0IvG0U+KWXSox7W8
XCg6/G3L3GVRAI+ttk06SO36QSN0cobhfm/ajVPqfKMfmwaZz+41buA8VEnqTTuS
IAZ26TO86Cd5hL6IghqzgxAjMr5UyWLM8gV89WrzLlx+7IK98exb0fhkmLFHcLxx
RBT3WhoSs5AGH7odOudF7e5dURlyG/dCIdbteboji2HPa0XfxiUv8pjmPULuqxw3
1HsnVqZ2IhP3o6vcTnj+Wt0a5yhnlKNiEPorUppe4SN5DQMuv1wF/1V5dFEuqN9u
JFKUARm7OJAf/38SrcOh0yG84x8w1cn2cbHwEu2p3ehDz8N6TBXWzpzULlKHwnIE
KIrMsVgAdE+i8AypJpORV2kcoKe5sCzMlTGbQDy2QYvWMQTBUPWLbKfJqgIlCJUe
s4n11yviZ6VJS1WsrtrNKb7eClgqSisn9TBM7ejzq9R/jKPXZP20Incgwmz6Yi/f
wJmL9sxkuifJ/Y/Oky8WzqBZaViHjDA7+0hxeUX49Xf7BsjBToD3bRYHAeVPrX3Z
LdcZTuRMHfUh9Er4DGaAtOpRPbUQyPxo73TZrbkfIR74IfGZtvJqfSltQJgiAicA
kVpMsZ5kVVgwox4pvwO1vELeSqPXj+lQbgfKM00e/lbcNdIp10b4OYJhsH1pbsDw
miPyHxG0YR6PGQbhiZQ9UC0UTxRp2tcd2gk9i07am/aLtLF9x7/JoxG1oidrt3nJ
6T53hAUNWkQcIoNkcU2pmyDHI13eAb3/au+RPF6VK4tVTXP7Y6k8A0B5iC9RU7VB
cK6fyfSQYFWVil1PiSf+zfcuWWLwognB7PfYQxq1Efu5RUKpFf4jpxRyylSRo00x
fCSwHbwa1XKyBxl1iVy0XluzcNdoagXgoudgxCij83Bjd2ByuLTea20nCLJRS8F8
PGrnl8M6eRZ1zPPkSuZ6U56WG3tiFqW8vwcvfDy9bfWkV1+4eIA4RPaAt/bGevlZ
KV2+NZPw4AcWwrjCXFb7sw/Aa2k05RggCUtCY0C+tcp8btOgPS4VBM4LLZRS/nfx
mCDDDr2UiQxAvjbS+rR/Bh2EpvIlZjYHS3Wm+Yp3iQG8r9ZJJZYoAzh38a0IXODB
PgeF5lT/TgIcPS2IegOnUTGLw+wMCCecyKsSlxfJFe32mZGnudpuUC0DeMja3MRS
Hctt4fwSaoowt4s2A0u39i6dTDUpuel6scBNK6xDxHxzbmp2fFgPcU9N2bRS23cn
O8FyfrP4jyPZ8Y95oV5+ICE9bxJ2qcXFSZivUSQa2wbY7/tBeIk/ff9FRdXQQfTw
SaXWNVGMeuxw3w/KQKo+Gezcf64FzyxdypX9fnvMNNlzJ2OHf3eAp7W5COT/DZls
dI6L+cymIMrD4aYj2FnjutBssC2WfJuomRJGQtVQ70Q5M6NtctgvDQkUKn6Hqc//
TCRXjgCX8kBtTwudqLAluIBPS8IK9rydjmjH3kt7fWGrXfkDOv2DjXEFqmZLpVeI
nUDqEZvcRffV5rj9Wcb/r6faxqDQ9TZxz5uYdNW6kKt9NmwzwMZAlbZ18M+W98rY
SqTniKVNlqrpNSZ7Jr7rdmDrUFFW51OiT0E6TTXuYAAVNBnhKFNT1XmG4Bls5he+
8et17RaRfJ+W64VQONMieiIm0xQvRpzjzph1qxKjwZp5VyPeoLok41neqbfvwl+x
7g38TnPKWhv+4eR5gBhdVlw3kVLq7fanN0pR0pgOrI5DUeVBH81d78MI5OVL7shE
tBT9/RlSxPSxfar/fkJC6IxEvqhguKxDkcHApsPGfZjGHeny89KndL2yroMvyYvq
xIwE34LO3CY/OUUkm+vc8TrRY/MASkiaDZmGYFt7ACygjjNrLb3s+udA3EPSk49O
kO4xJp8QVu9XkjynervOC3j0cw7vdjhTn5ccrdrobcu+/nKBvy6xWnGJ58vPGl7f
XWr8CxcGwjtMT89Pat3g5JBGyF5BE3CPZxc/IIwH7ql8PPlRWNxINFjL+birHaPb
keBWBT/MIcsziQJJg7nWlyD/vxtvPNtw5iVMfPZjMkqDJ8J3YQJZh1TOKiyJuZFD
luIJ0o8dY8gkI25W7atiAAf/28LpqtwK5YtbvZkwm7DH2RUPNH4UO7usl7DSmtTb
r8R2LCFdNq7MfnxbxkJtmnGBzdtLvQQsNleAnLiiGsO/ZMrJ2khqQjWI1XdLw+st
QWJy08romB9F2dO4f3hnxQZKoiqiVVlRQeNzBaN2C6n5iAVbxZAv5eyHWgn+Idyb
xbyncsIqBlKSxy+EmM0f14SbT27eCDVlbZ3S+zYTLh+F/e+W72o+6qnQ5veTZHS8
eRgM8HiWD7m/amW5cQiiVlImEu2dupxb1Qk7KEg7pFtEjJJ0EPnV/TzgcVze/vgS
eTGBwuqFGAOnYWTu0tkgU4wMHDys+znZ8aapsWaxBLOKMsRPyaw6h4BbLHhMaBbQ
q6EhOjPOmtt+GIEkuadseDZUuN2+QIFobyBry0UrtES2JA518+okNBMs8mAM0axo
SYLtlNgcs0TWUgLQKbA3yKdKDDcNTeSKWyD8uyyb/XSOXibIQeAnINwP2JNU9MHh
Wti/CJh3Ysql4jMCboqDZ/kfOfkLGlRUEkQvTDQz88t7bYcJ3dHR+y3/dS1vU9pm
r6my9sVrBAynoVNs4igl9KXL1AevXF5Wj7lLYn80aev6g7/atVtU44bir+6RwQA7
hxKAr/YHSiTFCBFN/Ycb3FCUh+Cc98n15fy8J/uOaDeFqIH0cHibPTduz8d7XkoJ
/TMes+PF0GZQSfdMaEWaAzX37X0AupJnnMmGc2LzRbLcxtqf0ciH5B2tr9dLgBmm
cEuzT4vabaya4mK3aG1TEXaRCRmORtnNIAXapQ7bRsd5U0UG1QjLTWldIhw15u/s
sZEgjgd+N4zLPMNS3n4FrpY++rMc2PcClKD8UTyxNr0UsLAuAnVgZW5VFH/9UBrb
8f0QKDHvV8SMVKLlWav6VkBwXA1uBGPeOiO0ysaOUEYBHRAlEF5T3Hq5iEDaXaf4
jDYphO+9oRF0iansAyiKRG80vnY4Pvju09vjm62yaCCKeMXND+idFUm7uumqLDjr
X0S6ioC3k0JhvurTrmO6Vdloos7SxlNZihzTC4+XMbRnS5T8uU5KQJc+/CsI6yTh
qdm9MFpiZqPOurJFgVKmNvg9ahj5FsLcrsmJkBnTZ3JJCz5jwfHvKhKvZz7W0Bk9
3KX4AYdPqwlsz1W5R0DQPIuG9dmBqjf/giBsspulhSoVEJ0KDYHsrKR++XMSc+j4
/rte6dSzcmwZUe7pvocEIZCA4UWA76eCUJGSF3YsnCCq+3tcEgapmw7ftLoSRHzo
pnUOAnv/vT5W6q757HEH5M/wSG836YWVIfTlbXhj1h9+THjJNfTuD+Ir3G6TkfGv
H/BTn+CraGpcU/jfiGoloxTBw+FLpBF7hVkOfk7eiqGv8vyQydOsOxda8HPUePWc
eXu9DmxtP50s3nUMgF1Cm7VbwN4iOer4D/trt1zbpY10sFN1oYfMwJWPdFR8b9BH
8VTjEtaT2rVBENPWLkjWcKg1dngf0dy0xIUP/EDkbOrXJzjloMrKznh8u3qtgbPs
52A7rRUdKn+/rWJqIYdIa0+FbN/9nqb+SLhsvVhJcgtHplH5MGhAQoQrFHFvkk89
nWw36sdpfkc4B6fKmKRNyIJNUy2jQG+JPHF+f8INwRx3XA0/YWFzUee/9mCRR4ZL
O4hVSTshSX8XkzoMwcaLfsKNmuvJqSeJuG6RWvUeg2YZmVovnPk+x4Hs0CHaMoSP
Uq3ZHojhirZuy2oHRWkAlY4SiBlfp08ehPu0I3Xa5yavtLHQmELYDSOzl/ntgZbj
vJL23eElX4A1oG/7P2ZzlpUIKX5jML/XkaxO6GplGppB8tsRLCfVGA8Z6OfnvJ15
TMnnIqNb+JLEaVt9tjI3M/x6SEKb1ZnBFebN6yG8gOnm3B1s7bCdv+6vJPxAA/Q2
xiG1WVqoSh7cs6GVdjDvqPZkBxnNVW1+zQDiOYA3h5j4sXHaahxxVC4RUAE7xMmc
Too6bbRpuXvfFZKRo4u0VPLx2Qo6K9p75WQ6l5vYnxw92GQz/QUHgl0sayCJVvW4
q3z/hG26UE3Zwxbf8szhxlMEqEruMcHr6CHX+eQRE0PtAEwr7R3z4mGcLFIZdVqN
8wSjX2mNZV7W+iF110LvZD6lQwVPpwfvm0T8qt3NbPxT0mf0bSHgzSllxo3dn+qs
7Kppby2Iwdr0ZDmDxi13GokppLcsNM3gnHQQENqkxnAoigJgezZ8LRjFnLJpNcrf
s6zpwY3CoAYU/ZTkVW3h1fhzKxrXkixlTNPSPEuZTmQCyX17kYVGEt97Xej9NW7S
SHJBky15nOtwfMED+PzY2ne2ZJ8PPiI+JahHEjAoXoyDYCD26FUEekc94Wf97KWZ
ZaGGxxeBE2PVet8gwCKx8g0y96qNUP+s3dWxE442o2XSxqXnpp4yOLUATheK1NzC
piDhqbfClwvxn7zkYGpFpIvtW5RsVzGdqMiouJIB1xq2KUNimlEltb5as4JWMRhN
DkD9UHLRCmrkAgZE1aA7hXDfzMqBPFKsGjKNkEjgUzFKiQgMUCeSyG2ARzAFhl1u
LMRQsPG/jRNoQbfORzxeSMumKrzdHXlUC+tUbBuktUEon9bYOtwjgbr5cGTTlPj5
dQgMaSCLnjVq5GbzCsO6FjBCTN7u3TC/XNjfdXhMyfmA6Sw5Djj+rwnDG0CYv4yN
iPTz6IwXEiIJBgabaDVw6GpB20sfN9HkUpnUdj3gTyQzEdiTIRUIr7abBvSEiiIQ
F3ISpvz/5vH9fnK+hN1Cq/unNxC3KHIW0t07ZNGEeEJxZz7zo+UQsxcd/2WhxkZH
79Fm9GCmIHs4AnJ/nvtyKXo1WxeDUftRLHS8arGENomeNQLAX5Rq+cS+bdwd2Sq3
o91dNu+F0LaeQejgQW7nemcS+Gxtv6Z+NOx9n4Bo4Sttnnolz9PPKOZjqQVVNN/6
O2XgzTB/SRLCsPFFYervPuzoX3cCRuoXndpkgMRgXmXjwlRbMjxTD6bQ5uv2qxI3
650arBSzH5lDleiL3ZBY/kteu2gr9oZEC6SL0o6Q0+OJU7EYsJNvTQaX3vkZRtj2
TuAUEbvzd6GwXUfxk4dgkvH66YGGZO5bzOJM+xlnsZs/DhE4VulVKnzxwL0p+4rE
eVWn5jODfQkJhHOMZmQfX5s8/9dA7oZJYoWYD0VHVNAa1RUoUE28NrkLc/P23om8
hrUlNRESDy9YfoAXjiKamothatEr1ReDQqwDbqsiTQslvOy2Wf26dMlf7FIeusjW
L+ZfeCrytszUIBELHeXcXW8zWbK3tM7d8Z+aOjTnCg75pcH5JzADwfgVlUq0PD/K
/p7TjaDGlR5wcl1Za6winY5dPQuWZZMSRsyuAmR7YzGHpVlXVF1VQEjCshA1vtTq
6MfebFQjW584A8sI611zcEG53Bn93ibcNmE0mcI4F0gBUlkrBbF9Lk548eLQLjst
rvknvL09rZutwDrRsIXzcuGPkPHCCaIHnFlE+Q8fSymxJk18ZOOMTpfPwmKMhp8U
ajfVYuKS5pSg+SwaJBKZ1fRz9l8VSkIgwhCli8HPLlsztJbQrQCsNiMf7ssi+Ipt
wTar8YyVXwrFfX5MxPwlPG/pfc/mdLwObeYsLRXfwjSpFCk6R2vnM/W6O/KT7xMV
etW+WwrgBKeTEsRRfFogxnW7BZ/miN0fY3uVIVupWzcbMteG/sjDV7k/NMTM49aj
l6oqd+9tlyDqWjAsenz+VskmiHHl/UcC+sW7cCSAzMa2IZcQC3GdjsbUR7KFuiC7
b0NfS7WW5DrooIjNTiEBq9YZvlgouI4OUY4Vx8FO2ZMENbxwjjgUt7LdI2zkc6Sg
cXxbgzTndmbJR618i/1usBIPOF95Qg/4bsqfORkfUd4TZjq5kuik3CwGtKgS9qBZ
O5WJKgoaIO8EFDh4ShSFEAtfLPPvYqk5Z6AEC0nYPLfo8sNg31DUj/faHBTnuaWm
WdMh6q7ziVQU2HoSrMuxCp3bbbytT2riZmPHK/X3kGScmTDg9l7Ks86g+WcHc2Ci
9g23ElWq7U3RDy4p6vp7/re4SAD/vFdem4PIa4O/3N+CSyr0ErG90YTk9S6WPROr
JUS5YOy08Idf4rZdxBNu4Cluf3LDKk372U/CUomCPAHDIzcMsaC01NV22JKJQ+dt
jtvVFuATB/Hs7PZj3G/Fs3/A0eczYvdIfIF2KHO04yFMK36X7l2wQQVkaK+SWMw7
10j3aN0w+O+C++5IbnOzb4pW34ko4nN+ttFhJzI41KgAE/X24hlaiy7F9tuv41kS
6imx+uwTyvOZNBLyVH/FuJMLtsHTJRQj6gUTgO7MF13Zm9ehQTJbny6WNQJfnNBM
+b1SkYK62e+Cjgrwa2eRDe6hutLkwAJd3NxL9umemaUq0+TnyODaQoFK992YoPpB
oNPanKOjTVyyQrti8nxIhPCBV2dmKbp2P/b5KJqVe/2gkylSC+hIcIyUGKbuy8OW
ttuuR9q/VexKLSaZXd05ddNPAYA787KkQ7L0eAfP2W8dFbPzDxkAVBbsO87VTKNm
z0EUIKKvoyLeZqDHaqjz/NLs3/MKR2lesEfKN8WW1afn7Hv31o8ScS3PBE9f0FV1
GaNO9WHJmW7oKEOTDUv6pFswl8994n9ld0ihNUsybYYvTqDQ+YJYBz5qHpv2eWc3
Q/4jQSYnjTtLNte7oZQ6lzRNI7pW98t4r5FAGv7lHA12uLkYnrx0P1kGhJr+8o22
9plnCw8WnbsebTd/a0g0nf8uz5jt+D8baaFDOYtjCu8FwnRKmG/xLAQPnZjgBJKh
5OwTMe1te16JGY1OpEE9cSniwSlPUpzY1CtG2mmFW/KYLQ0tBYF+01HCuw3OQmDW
+YqCg0H8W042UdxxskXlUMEIcRJF8L4GC4DR8wdAQjvge8WcLBg09vUH+IE5Z92g
Kd2hwMMrxotzo2eYsGiUxAhhCJGvG3DQ0sqXEESUDPdS/BQBHQ4qjfHh2rQruxY4
2SrH8Y0XO7568WXGZZ11d+cNYIoeFog4WUVlpy6pwFRMiD+nKGc/hz0w/Bwo/paD
mQjaix4SDncXrfdbdIfFDIKwwTmLunlnKDf07Y2jr7VsfmnJC41Z4qtDuVSAckwV
7isOtLDclvzlIqTSV5g3eLGgSONXEOhpWX07eLiiDF+FE51Kv25dBvgmjvTVs+JX
BPUDVmcMLAjkTjImirGmRg1ABJ2HvLNn8i4Xb9HzSGL8IoC0E+ljVDjPMp0A5eRJ
vXm5rcRb/Nnq5ZadyRyvpVnRz2ZmE86XTVuQ+MWuxyUbT5bzKtW2VleDcx8rQY0U
LoygsizoaEFtK8UzSTjOco4lRzFbl/qM9f/3vRj6TURQGSLxGOQ8oXwECk6dUic/
apbG3XXxpt6snS5zLETn8I3MuY9j16HYmLduCMOpcV847a02TBu4MWZAB1to5p8Z
s5TuTFD0li/+1iZWRh8R/e+QfULbrYeAmEuydegJPi4FafTLBuY4VeBfMiqKnMo6
pCsDaPCyMxBrUSLRP9cBgW7uoyaL4/ck7SpxXQAa/gGHesNUv4lhmwJwXRN3Pldc
ClzxlMzfD6NhMx3gegVGJsT5KKwUTXH8s44ij753ul7jDHyT9EsEsR14EmBaUORz
nGXMpIwQpH0624zo8azVP901Azf+omZOiTVjP1n1r3wT1jI1iElR0LffWTx1X4gd
hmkfmgfdJmyhdEOydQu/Z/zzkKqeEUtSMwm4GVZ/yTaEVFl7y1jFGvIOHelNmmzh
N4MKpSTkAoi5u2QFgqk8gT4TT7pMyG0KUtuoHkMh6ReW1lkpTz7LrYq1L7gpDzES
gJZrdnHH9s2Y5zCiJMuggPiCeVQ10PXIL6naOya9kTisusaP254nXccqQZc1BcQ7
YBXhQLEUpxg8ZdJlawnOFk0tBFXE8lhXyXsEPM3pw3xixKZkYtrs8nlVdA/QKIsO
fBSJif3sFXQroziK5ZTvpKZhz3XIMCkQPCSLNyuc3H3PEhEZGWHMG/fWbqgj5mm8
UpMvtn+WqYL7OIki+Vl/oZsTqaBNp7eB3FJhuY+eyllxGdJz9ViFfVadguG2EBQf
iNshhGz/9MpYs/XqDzlJy54Nh0rcbpVXD1EgIhi35t+ZecZac10zgcL7P/sWh4AJ
gd/io82rSSUzmXlalmtBWbK8KQV4G0FfEoblyq0xjVV49iKqUQWpRKn6SCrpOHQb
LIcq6A1OIVdXtdRawfZx7D2kGNVumoKUn3n2FD2vNnZCd7/disa35K9PYaHeVmzz
OaWCA+1KIO9zNKi4gj+ROQRx+SfH2DwYLW+43Ma5cvt6UpbksujWikTQZySsG5hn
F5vfbalhGbJ++rNdZtkK8R4gYUEutN2d76Kwj30I3zyp1ld2cov77fxwbnpp5V0H
LFxtkDQ/MIy+yKB+ExoqhbmeS6MDTXSsmaqb54AHQORLQXFeSDnet0m0GP0zW+v5
Q/Emivn058M1Uv0fGxBNb/vA0eUgq9pv9JCIqmqw/HhtA9Q7l0ICZErT6GJlEsHH
/c4I4uk0NrnqvDz5vjwEFrldpK9t8veRzkGM3Jq6S3HnJyBKm2pnzTOKZ66R03Ct
fqtqlAzDzc/mmrTKCwBYQNflb2elKc+y8FEv40xT6gDVwOOY4G8Tov+DCa4ZlCdl
Lijnpc3uILwbshdZQ6SR6j7bnoMZHVMbWvTVHpcNU0GNt8EWwMt0u9lkxcVAefzy
VjOfbahhsil+c2CBdYdpXWGKiJNZ4CQH8FIgZe6eIezPKAAnaPTHvyjxxtXCdFuY
S7txkj6/Jfl8FFRdgkU7RF/st+j+oXhqBwEp6r12aqs6q9baSVUANdf07YuQK/a6
945Va3J6+hW7TsOX4awGS54iEOrWEEeu3blKhtnb7Lh0Pm0yTCVpn0MIIGvizYnd
oJnn1fvjpOJQLo8MLCXHwGqDU/iruXhW2m6tbTcGvd9LFQoTPS6u0RjJY1VefE0E
ehinGeLuLl5ZvVYO2iPr2Bn8a/cpFwt95TcJaip3oZLnW+q0dmWaoYHY8dtG4cGt
zQBLIXnDtinDbV6pSzGCYYtzA994VZrCx+9XbKZuvbjdM28nZY4tT+teemGW0PFC
bamGleYOdiuibYYlI1Kb8ma3KKo5hJEcx/0K1idpDTjIL2mCI+r8gO4IikeK7vdo
vvZz++p5HmpmIILHRgxcRmmeoAE9t/vTFXxqMVzJnsTd+vdd8y3zf5DuY+XU4npz
3yTRPqf3GSL83SPuYavF9MI0WorvgGVghjbXaxrdtSJOxjeRo0zFoHfgWZ5K3pzt
RaVnPkP17Zx1BiH5wtLhFCVeP1sXwK1QUkUxVx2S/ATq74fkkqP8HW8jFEiyORlZ
5PBDmvCnkVSNvSacEMj1omAlr+5iFSmqtYAXSJNcUKKFD7zvMWvuWVLg0tyHMMlC
/T8RNkozgqVV3C7mFWEyqoB/+9HGyWOEzrePVXmZTffYQ4CdxJR8ubBZ7pGwcdYb
Z15smBc4zmjNm73F9vIGEdi/2hs44hYTeYHMH3Fqygi2hmJO+5URKN2Ox32f0x7f
4RXING95T277Fsvz7Qn3sJ5iW0757KFAcsDIhTDQ9TXMbrHvrl44ffIJDlHVR9Sx
facqVQHQ4G7fyS9zLHjq7CC8CND/WeL/MjpifO6TgKccBe2sSCWL5Xc6IVdHmLZs
vzq3A6Esvxusr/BpCZv8PNxYx+BZ7Byce3gtGD+IRQyqRnCuhSSIX6qh2iu/u/0H
vHgADuwSKLXf/XpyA6Bnhjwc9cj5WP4NAR8EwlL+fsDeqwRPNw+OJlU1lgiYwel7
zOrD0VzIBF+tC9XNKVug3nI1GWRMzDw5MRmihKfcYEP6IM3Djpvte2MyqWgTA2gE
SuIoy2qPOrQGWAZ0bs9gHWLioPaqlskOnTv0Lfsn8886R7zJebTMSxJzl+KG9iJ0
XRtcChCQoZbs1Gd7nnOBUZfLnJxSr4Y7wn13vRty8Hb0ElOVITKWNCUCtmWshm8P
+Yqi/ja0Kjc7iDz2XIWqUuv6NehYorvw9sV1fUOd0Rtc1VeXmDo3Adxt9JG9iufO
WNaNQ7WdJ0Xr6aGlOSrp9QLbh1y5Bj33SamhYfPUxoiusZeyu033GD1FXxfZFnZC
sji7U7VbZi3f7mCWc7Qi2xWion7z787qpfZ8wrLf6s4P+XPmUjm6lU1raHxETC6J
HrF8AEKpItH32RaopBXKUb1GlajqxvoSKyAUfOYjcUGAiVydnD9ijIQ50TTE6gvC
8V8bGHEuQMoCF3qnT9Xno3LmuVzUEW3ZR0fIvQf8AMDlLenat+wCosM3+aUExxvK
43mcdHPMtJZubwuovP+8VP1HPMXaHyanK/kFlWNccYspljv8Lf1lRbw136MTFH0u
gRw25v5q9wGcJhUm7jUK8EbuTitDncH5LoQXynqrNU7CjI8xWjotJ1KwEojWKO/J
7s21hJRlpzakw4EuMDl6C8bW7ccO0vX/ND80VlBVGYPW0zUGmkfjQQVElB9q8uYz
IcwtASkpPs7Upmd6c4c3MFZkv9MEQMsFIRc9zlJeJLEV/82qQ/5NwDvVJ3Sl6NuD
Zea4AMyxT2+Z820wJKvpYeFzoq4wFZauRGHqwzP9VVf5ahh7Zj9/Qk5c1ZWsUUpC
ofxSWs5MfsRYLki0jy6V//uQ3kcuUciwC9YrpjvJRBzS5TlNnBIc3lwTDqAFOaK6
iuWbpBnv+xRsbGAipBHdqy8JkWggLF6RF53uBEnbV3VwDm9Z8AYMR1YsQ3VsqYOv
KzeFsia3HLGdJhG2n/CPSNZF88pZmSN2g0enAhejRcXmwSozYDzNkHJKV7qodD0D
6zJeEkESjJvGQNd7Nc+9mpwZBeBDWtFmsHbrPlUr9Hrjm8XyQCgj7/yoWeckew8y
w2UFJXo3hLKNzviyMGgrJgALtMujnPEfqPxT6Yve9bZuMJjMzmr32Wziiy5zljiB
sztxQ8g9aOAQiIFoOktYS0qgMfmGh7t3v9x731vRfDhDd0TGvVLwGie432EwSZxU
YRKoDqbTloa2BXPY9g3h5N16noiFsPak1lk4dfcDnR7j2hv/L8x62hgm2AY+FzBo
597yi5idChpS0UZk2I3ss5o/zMkYW4LOWfN4hYZC181EROA/tZluucjTaXU+TIQ9
84Xqz/UR4I/hIylHrEFJT97jNfFg7UHXpoMiFADbet2U1+HqSeDIF8O6sXP/ZmNa
mSW6dNX39Vnq0eZlcydgqVvu0eCEIA0D9TDHgPxnirfC1D7fisyrWWBiUlMV1p8x
O7CFUVvlpmyPWQOUP8Zkur3p7iwDU5kyFa3dUYwO8G5FPH1cjMCP+9P6sxI9K/HI
tV1HqVJVOyGTdhig23b9VO5UAi4exNaELqRHm5OR4+DHjpLqSIqDscUVu9pZb29b
Lp06vlAG8uAdqffqCkYR73ZwK+98CawJS2a5FFOrgxp700l7LwyS/4hlYAdZgBqT
ZWI901gO38IY9l/TqieEUVil1bYpnjIiADaYPqH1ldDAb3Gv25YjgNhYHMnVOF+v
kE9l3WQE04l0bEM/ssW3PuiVO1F8R1uD6ROqGiWGkj+gXXj6q2vQNcQY6WkcYlxX
M3x96yRGGYBaWj0AwfKGCKJr+atUHX5kHzQp4zfmhhfXYDgXG/XBxEedUKjeqd3R
2c0oso967mr/99N4bVerj9DPjH3EZLEJYcnEIRjfCdOvtn0McjWVi2K+dRm8a+b1
aSm52jmksZQVAQWLV5CkA509/oKUg4HJLE65y0JFr87tg1yGvpgojLDPKnqUWdP6
mOpGF9mD6cj2BJbyV3uZpLynxb+2IaOsBq7e0RpzV8noxjhM0bBOmQlkui+t3w88
tWNvOz2w3+8PXv9DhhsdoXfE2uI2AvbiSBjW4EEtbsKFza7iGk9H58Mtf4bd8nbX
Zj4ABmDU2BHDLZyAELLleF5+qpImtO73J3oF/z/x2R/vo/45yRLyHVs8OZ1sx4RK
zvdlr+xiUUjb3hcg1CR4KhkVlwGi4JHaiqNA7nFyf86Tj4uMADngpdj0aZHGXlL+
wso7QktEQ3TSsDNQzGTFHE3RtG5snw5GyG0mk6YUIIk5lUtjAYuwDNhUfikphU2p
/6WDVmZqcv7VdtBmVKVvDRlMSETNlL2geu0Koie9bNs2CPRrlpi8nKOEwfmO78HF
mKUVg9ud+dbMiA987ro9yWwGcVxLpbbKQKeUHDtlv1eauRzvHHACnBvVgUiYWt1R
Zw9D8B9nmmatE7yy4MJKWVljPB33D+mgXPd2+S57tCOPFHyjsiKZRvP8iVVc5z5q
EjHQ/7EtiWkEXLXGeF9lcxYWM+vJxfLJ+9u/fgGVXM4lycX+ToEBS7TeMqBR/BK1
Mor+EnIhtse1FPRVz5nDwDaa5vAoXk7XaJ7eHtju/l6KwvQbq0Q1al6iABP58iCN
ngI69slG1+oj5gO2QWmacz2w5h7sRbEKWn36vCfNIj4A62vjvrj6nOdrneV8Q8F1
TG1pzpzaab018Ay+bHKLkkRkR70IxtYW1sZyp5KLi8J6Rfw5lMIvp3GdiATd6+0N
C6lmNdJ42qTxI+eLxCqOG+bk1qyGPMqNpAIttQYZyuqLVOwpTALdhr7SfCpRqrdq
ywZzCSQHDjFWkuQIeI9Ogl7kFD5NhtMuns1PmWMFNXz/w+l0Ume/j3eD0J+N9Ta/
1HgLyEpf8AQWucHqOEz+xwBMeVMvaR2KtMV6SslZo/W1A7jqN0RJ4hs0TGxsewiL
sq2KzPf4K4Sk92bqP2hHhM1H9uj1WmJGeaUNVdl1f+U63Ujc76KG2/69vG8OS+8D
K2Bqowpfiw+AtzhcpsLFy7hW8Om2XX1XuQxXVNXhq6PO7Sm0jC8QZH+SvDBYgLF0
f2s6ERyEa4HdxIf2NL1LlHBPNYWMzz4rt08Wrg4Av0ycitTxkXLWvwo6uiCi/mBX
yCElWduZvXD68Spm8RIeT9Lt6R+lCQ/Q0N0dYu+n/skIFONapIzJOIFx083Sp2cn
2z3LGDNNgQTGy0q8aqLEC8GCvaWD56ATIhpcp9la0moKL2KpG7KRcxgLP6x43v+2
8tYTHOX34XcPKY2mVFCv5hgnp410hQRDFUz81bub3PCZeLaf3delSgOydEUvPZmE
xCnwQtzT/C/1Y4PrZCnBNxYbi2/myop7Nl/nTdFKCODGlHsm8/qZBZ7VL49dJVWN
TnCdEh3M+O07qU1lnbCaEphdsulp0LOn24zmxl9NUus+MR0SR9SlGPtufgvMRHNh
kgqpDT5TIkH/07hUu3MHJyaG7wKux6YwlZebVsQIDaw3TleEw582tE8FsiN2bBMQ
mVW1zBPYKHOXi3zuDJ999jEm/il7gGYKW4fquoRFpr9lunVizDrFitp4KWJlL+3h
3I1OCH5KfFbq6udEhw+jqn/ozRyTYD1MsXVOwJjyyHzsbDNcMpzMKQ2SgdupLV2w
5fgI2swHU1RZdfQiY0ahAVmN6WAQPpGYeZU3Nlh+EfqmKQTPWIIl3/ipLwotl7DT
A6VK1IavXyUEwY7Fu8ThyqMe8sbqCSzoDVTkMAN3llRJ3JBrA7WAsAvHRRbZ3GrA
PFnYahlqlIx21v3dzMJDGywhQwwf/qyqCaUCyp8+irGlhcHrJfKpMLov0r0yJA/5
1CDcaF7Pg6Ry+jtR+9TmmpbvM5Cb97TYV3YRpw3BIKYAKy4+8cFJXZLQVauPgHzC
hJeiB7P1kitY69X4e6BwnHhxw148Gjed5kwlAI+/BXVYrWu5LcTUOP5KvWTfGgzJ
JfIBgZdqeVzmm4R7DuBiFxTW64CRQsuZTxsQJEDKM6L3/XyZzzPvqW2pm/xu+YGS
f7FvQ2JQ2hOiKq8kgAbSI2HbTGmY8cwMuZN3VHtDdKQO8xrTSkRUNOIJLc2+I+YU
wdbw0NPRnwxTiwzRKBvgRXsRGUN2MCd1R/c9vDlzUHOxvA6mXgIcodb6HdjvQ99b
6pZLeredhhupwq+tRp+nK5TDO4kczHgU6tq3joGBkEZ1oNBtoW8qjX4OYIDAKTTm
kMBqJLeCDa0CjGzSTFHrlIEwoKsGjewP1uuDuZrThmF9tX20g5KiPak6DGNuIUUW
UL8yYHVuIcf9J+4zev2e3XXQLCy7vnF3Ycg1gs54/AdVwustbfQlySKbQBFu/ZUf
paO6mjf48/as7jRSyS45rRe3baK+eXZ4+AsAevTkED5u+6AQIekThShyaGCJCd1V
G76U4RRD8edHFjPvaAXzCdd5yJo44SCsCoetpYuwRL6sTdValXdvmV0hdJEwj/AT
v6GKqgbr6orp4JsEGMo5QDDiS2tK6Wtj/DMvumYZrlRfP4D/wondx56d7PQOHQMX
mJJj8azlDvyi8WOwWxtVJ5kFl7XYKHbCQqFlEcWH0e224ZkWx4lj5Wi1YlFS8Dll
L1CVblQP4vdUcZrXmfytz8pbDs6Kwo/jZ+e1DT6QqhuzeJmZO6Ua5/CXfJDbbrIv
DaHX7ewl/LWDinjZdaDgCkgn1p/ZkZWH1IdzasZHEDFo0gK4CtlvKvh1JdNirZcD
xYPVtsSTmr8RiCfaWq++E/kOjhybAxe4AQ9ugcsWUwFzqbn8vOJroCbBfePRlain
yQSHiA1UzTYlesjavzoEgnzBB8SWP3lmKQ3TQJdSlzzEI87DBYWmODfOLAJ7p4nP
EUsQCyAkR+xhhfTI7asJq4NsWxyqTj5kYU7NwTEr8kfO4Og7vBhiboQLamMuJBKO
s72IA3hi8UD/NmoAXy2BpWMAJ3zFxyhp4vcgqz/c/vkv6m61aOzrFrk2UhidrTNr
DCur+DVg45TWc/UY62VpdhR9eC/cutalQwFPiqm3jAtUqlY+ZRj0n2Q2DWEiCEUC
k4N4Gf+ByItZ/kiIeth2ZMttW32z94TFauZ5gkMZqvUD213lX2KgbhjvGX7QafrE
V5EYN+uh502WZhZynkyIK4pLIPFdrsUpAp/8NwylT5EqGOY3adUv2zqvaI1kKJAS
GOQGe4XeDnwkK7nIpr+3UVBNsd4PkB0tFMyFMKLqKno2iTIdP4FJZYH20/9s+mMO
5KzvZYt7LjuoRHfOtxOg49JUrvHObbWB4pEdjzzrtolAuBU7q20IMjH1YEQi4281
Y2xhnMBvfo8I4D6ClpmMmqmNj+vSx0Fo/aDaF/B+ULHE5zZZn/RhxUnlzYKhO3pm
ApBC/1HML9IqJ1yqfaYULaKF1la59EZy934s1RFHzA4vNZG6kLyIh2Izot5/NMHy
YY6kYAc1h8RLVTB3EREA5hhZYvl5X2TYFgyIYPWn772d68BOMNQc88nqBdDXhXvM
smVUn3pzoZ7yQTvYd84GgSuZTlcEp5Bg4s3sBC4R9HfD0W0gkt3W/KTIESnKICEd
jUjfOyaO/sdc1M9vAs4NXUrdZj2d78frHDRkyLzWfjAcg9Lz4xVGwLZvIz19pAfI
UG6EXzfDh7bp7SffwTlWuVGP+XEZ1BTQtBCNI16HFFeDx8WnIEhIa2LVyqMiYiJw
xuwvCm5+xDWrsLP4S9qLW/9SoFT//pTGoPuo+Te8Cw9+9ll7thwHrhv1RRKWc4mD
97oLsQqRwTC6RrKxa3IAbbWaCIljFpdpX3bFcGuT6dyaRBQuFf1oiN6R0fFy31Vl
EsFJXDaPiDQZmA+srtI/7y2abJ1lBsvu7tkAauUR74hQInyMpkSyoLwttQcnr43q
DWxt6SikaT8OEmJe+O8PBI4M9Bq3gMQNecqaOv1EFU4JKZHE81Zmvm4KBCSvyArp
LRJvq1ZSwRxwUP5CgwSoJWigSPmck/4W053Cch+Edno31/cGv/f7tnFiwOCjVQJb
QG0OqpEBWjdfR5+ZAEJgkfyT+4qwuS7HQDCvi1709C9zfe6yCgKhqzTuh1uRsukd
0wJzYaCaQCw0omZSzx7IC5NvuMKfL7FtwZJia9snBNBEaOuxwPMe5d3vw9724Sdn
yVZwZdlm57xj0W4L+XaFEVOzb/k7N22Sm1CDjZ2lxjg11vX19DDwWKYLg6oiXdIZ
QvI323uV4+4QAXKpZGOxYn3tFFjcDJnCOLe7/m6xOJJCSCXB2H5N/t/gWWMgPaoD
umKQZrQa8DFJudpiCGSNUSp1DNB6sQU6GpnnFfYvlQ3HJ5otJVaFG2GSR0EItLE5
HHAu6KeuI233vhbU0ag0DeHqGgHbr0E1G5GV9fq233NiAp2GZH7a16o2tMY/PGXr
sgi2pGu4JTMWrDFFjwV30F7rnGZ0IMCpKrZhPtkrqBMT/m+3BMys3/sco5Iz+7bs
oG1YA5g90zW2xPJXtNokPc6GM8z/9smm/MN3IxYhk30vyE1OoyJ3WNMMnli80+UG
PNLyCRiTH2+Jft4G+UHVZTYTwYctHL0G7chQOHP9zSlYLr2ffNB/zt+CqyzNaWip
w8GCHOuVGsO2ZWl5USpAxRpIdHd1Am1nHvhLmxCj06blLBP0s8GM4Q02c364h1SL
PCDeQkci3SwwIhiVQTWLG3JkPQj3LHAl6JbiGvYnTYuAaDB9XLqETbsJEnFikwZg
kk/0jWQ4oIIxPLP10xoEWopDUTYAaBK81OPqS+fHIDp7Yqde4gwPIPsJdTCDOaRj
/+Q9BUoyqoACAk74UmZORa69b5uhtIS6s7zP86yZ3GGWjdNqF5lFqcf/GG3pUKeX
E6dUFAToxVqtnwl3dfKNvPfOmr/UDI7mfEXpYp6vrMfQYNWIx892wYaulQtS9/Ws
K/2nLsCO+uIq/vS1ISAMp7Ml1WUBf588bHYfUd527ce6grgICLpiVVhlLGV/oiKw
R/rpBWx3sO5ZIaRC7/UiQ/fGptgft8Hz/w5o+5lUK1F7l5zZZTpvVyimcdTaigLp
TAgR3yYO0dm4W+Y/JNTgQraCxBR9N07uycLGwsV+V1I8yfgjZXZPPKrygzoMmjip
D9Bp8MTAFQRR2wKPyZoCQXgTx8eFfQwZCGruUnrNSu6prtxm6BZ9onCiZwPIxC7A
7POkMS3e4rjFH1+0j08K3igZuDAtN6lDYxu7RS+At02lOK/wUIwmczvaCURXWSyi
sFf8d/XDtfLr22QCPfbnreMh4sjjllKLDsoHed02r0tLZfCS9kitJf5KjaHsjZtJ
jTi8qHlsD5m2crixeA2cvQ/lhkkG1B0NPe+HDCqGtBQTlFkZE8NR/k5aCthl+2Er
pLh8yXWTjSg/ruOnfkY2iL1fhJ6GB/+8KHjCQPoMd04IOYWbKH3O2/8yDVAp8x7S
Oro+YG5148HHVXnutq0O5sbaoTYDqVn1+Cc3Impwg9nVdYYMKifotSD5Ks+rZFlq
rnKAi6OUnWZS8RAHN17iHcF5hfBfIy8Ner/oe3BGEhy3gH8tp0zwk9gUMDBxlBZl
bozjaSZAGpqtk7+nofXmY5xSenwowjWLhSPRHWC9NhhraoVSjOUgsiGLfFYEWWGI
iQNdCz155vZZtBb+ZFOpmD5O2QS3cfAv8Pj9UDmR3ThJp0HK24NZVnx8xvsvqn0n
acK0NzypiYElIK4g49sKPAT/N0Ni2kHKpzyi0k3NoZHwYQsb51Vq6ZQdHEq+CGEE
z2H+0y5xHJvvaojzJMmd1VXCw2vxZ5bt1MqMuACCWIZ1qcctNEhu8TlvFr4/QOaP
BhPjMgogKFdm5zbBq30mapt+TdmyRTgzwwggy9v54kZzDM01rzQmxfv8zfra5xjN
06twqBnfnCkW8vidhe6keOmSp3PziP0TVitPM4EI5F2pih1jfMjxBGYxTI3n+6qy
a5iV6WWtkergKrhU3ckzukdhnpWQP4iMRfKPlPQYPtdm6o28DccnagQQUVfRzrkv
h3A7l9i+BCbCbbYdSFgBVyX1MtTxwbDeCutIGWkrkR92sDq3rcOFQ28oL4f3Jd/m
HI+rBFsyRbDXGVYHvT1pX3pANYqEAd+ocKujxm6gc7I6/Xef/OIrM/ECZTTGtUeB
LSMQeTLJ3jsaMXXCKSZfC/czE8bnzXIWshh55J6fZmflUY7cHCHNv5pPU/fGXWNW
+8cPYcl+UfagVLccAloKKV4T0Z881rWAtaQhpEPdaj1qA6GKGg7GpBs22SdeujcB
rvIELTTuuP8FiVHGi6oZiwtTAsQq4AsparkjaM3Cd1o8Y+XsYZpqTGMJx1g7/JLf
uiqhduAVK6nJcpyPCpFKTHcIMjo3eiozftrIZItu4krLoikOM5Sxk3Qaduxp3hVC
VaomWXSp2jfcHnAu9J3wNfyn79Q9io5Tu9Ga1PgQ51lzu291GKPoiXgWMsRDtJt+
lLh0A7jdRnDYUvwM5j7pEEzpYhBJ2ZD7UpbgQ9PXuxzQrtgfZOaA+q3Qp7v9uwNI
o+xsN7jBsMN6inmZnda8+GFL9fGVlq5HpJ4HhgRshSaqP3mWOsPMzF3nApoyyM5m
jigKDBFg0Nt2WdKJsaMnB0d/XWkp4SqU13s2ODH+hFEyDNKuYzGwEiFGraF7mOI9
u7UsVsPD4G3xH9ev5QkhoL342jKEMto5mfbAKTztBDqWYJmLVTuIsKhIFPLOs6yK
izJHQV/7PVtvwTdAhVm+lFmXAm4+VUnW8RdjJ95fTdXDypa15kkbR5Ks2npitMhd
nLv9k+FPTehkmlj3a5pCCjWXMMrfWKPaYcxlQ7ahruwoqz7pCAjh2h5SgjnPfUoJ
IVexKVwF6nAUN2AGnaPnTquEwmJkrO/Gu7T29+td5k68fQu7ImYTkdQhIbQsAI4f
KFOFLPmDjPuNlfeU9B5cLZJIgYDab9tjKEYwZ/kGsb70p0drJ45C8n7dpoahT4qu
RDgtuQMy3TLX9u3qKLIzIVCsYFUG94sQZ8UiYs5iUre5JmEeNStDWLZU3rwCLOlf
z5nEBAR2F6n0vuquDEvpXe6Xtm0mVxdJcqJmfItZqRPPJI8BRBag/ytR3n9W2kNj
5MJ3DNrRy9iDbdIcvKMfVzFw0ZR2EicXNjMtLIadBwrHDw7CFfEmCk/ugOH0ACWt
yJgQL9BSkn/ANWYw3nBFAA58iI9945mq7lLt9CIJNf8cZ5VZ5AQsQ6cUR5/yT1Ql
6A6SvLTKsTjl2P3wo9th0dhc52qq4MBFMv9f+nAD7XJ0Qu6jz+UNzseK+aJyTVGJ
/aEqduTgRZKnzVUg0rfEzot7U/734nBQ6dgK7JqnYTLtnVrr2s2cC4IQctrBie+E
nuUwXV1+EnKC5xQEpFXbghR8DS4h7diuNYduwd/OkYbkDl/dnluwebZDEcOugB5o
YDW3/A8bnknceOLnQsldm3TO77VkFzcAG5fqLaWCtlwYV0FPTQf2xCh1vHdoBVZD
O9cLinZN/nRo1sPNQsSQK2E6JUGkkvdpbaBh/yT6SmJrgjaaH45dXjIeQrAe1VdM
ynmBTNHiM8OYc53LEzMm7LpF1Thhn7vF4RfWIpJ9VXJh30qak4hfO5pvwyHKqZrp
olGLVe+ddjj9KZuvXhVS8NP+jE2T5PRQdyhL/zRtDMjap60psHuYOKTbXjpUtQ6K
asYD0TW7icN7oPj0krn4hhclqQy7d4PKDTlr0d34w2HdAZqvc02z8/GhN7gT6N/B
7nuCGUWIsYfW7qFa8yOoZc96TYPRTVUMRZC92GwhCGZ+AXu60hAa8TVxbLnGsgTy
kg89mb9G9LZJ2GuFVvNtVxzw5XxXcjrKmygypUxj9Sjc0F2XV51OcSGGSNheDuyl
NYY97BZiQg676FBLpP7MXAlX184jB3O1t+QeI8+DrVQzz1axDF1vyIXlYBVx0ODz
0Auex0V75cX2M3bogc3B3EGPn7tqkn9soUlLMLlllBjDfOr7f82t+9O6MKgRpxFy
WfBlAi5lTSQ37xGBanXb4JW+d1yoCU3bW/xanEAYFNtAbVNhqTR5XFEqTo1Vjv6m
DpVofJeZGNBEqpPzy3itluQjfN69RvTGRvdAJkoYzfHC/PUUm43hzEmuv2eHHvD+
Gi4ofTk2UMFGqXhGaGmq22w1gxqbjgBy48MVdr4ZgOCrSw8ZeAncDx9S1TePN8NY
PwYFupmZcsdcKD9eE28dLzyYflWxBaX5/xbfk+u2nPs0EYJT146jqT5BXYu5nq7z
7cPdm7gr7eus4MmQ1Ma+QwrTDO6slxtmRom+XzYUeJ+cHzWxBNc5muVwDbpx+7Qy
sZbbqlLzLcG8bTAMpXD1pb6xGIsWPUrhM9ZbSkaHYsX8S6+RHzlavK8VmdB+Buo8
bRn6GznKAs4ZPPgGNXBkYHSg5Kb5975R1/r48li5eYTCQ0HhPiuXGjXZ9Bb0E1IZ
e+46A8Zy24oWmoCct4wJXUBbNt50bweY7VPR+2t5UBmqcOkCBLmU9PiLiar9Tlgo
D7OFrU/N0NIVGTgQQEw5ZLk0q/LPZqOPnwiC15p0mJ4jtXnpD9xUFgQvxfWusjQo
cFHKO0ykzWw1N4zRRbrPBCz80kqyhFqd9yLz2pG3bOtXRxRtkXy2yZwLAIon5T8x
gsRRbYL/3ezklGeJxfBHqGcEGJi9q0TZYXSEarqmae39iMxOX0nLMtckK8rpWaHd
umZcH7mA2zu0GgiE1BUQI2ZIryTXTe2SuxDJ5vQK5WwBT/km3vYCn3DvIoOfwAVn
f55udBi1Mi8Gn8+dLf90IoPo0i/Vs3Af0zsXG6Y+q/SMx7rbQlQqcHdWZL0kgD/m
pbRnywuzRlRaol5103Dg+jAVqyt7k8yBqK1K+3zIdVKvZpTPL+izxvuSUZrcgqwg
kbqlguVkaH62rwOBcPcmkpksckJg5rTccenOPFgLhDukri8Ry4i9eDmGeBF2FwPW
ZG2kFZ2CcmNc23F44xoWHl3Fxg8+CmrXxYbL4RG7+jivleZkpnJtKsMrsNT8JUd7
JdZ2jzWuuZLTfGMU2NdjWuat5B0yCzMe5l3+5xSLshW00bPrLHTJC4Lb2/b9S99w
S9FlCdkj1yQFQJW2KgYXpjyEuEl5BE03i+GS4AD5TzkLJXSXncyIFFNwewnHdqN3
/dSKgxp49FJBcNO/iLWIjq+PlTZxVITIcAmtmH4pJqtpMlod3GZHC2sNy01SiAfe
aCkbS7WVrxYZIhhWdNozHTMEtPm8cTkTPJjh7ttFkJxMlxIHVgG6jCSU22QypAkT
moBDlUnG+cEWPdSZjH0AtpM9twLKNIPKjn/lJ9uLQgCIDFeWvmw7UW4DSd+vZH2V
tsabr5gsSrVPTGaiKY1qO0dz9fhZcdR+uSW5sj5Tb+wGPaumDPDXif5cVsGv6Y/s
/nTzmrxZuHgVe46QstwNrPUplfYEIrEa70qHRDbWm7GqgIDJ1Urle02cK4Ul9lRb
6RifuT0xdAE7pHGcPwdl76QxS6cxvO7McX5s92rEJK/+dFcrkbrPS+EV3n/ukYQV
yACrZIywM9Gn7SvMA5a4Z9xrZiXmyLH6IdZOFsuPqHIdNbN1c4iwTeFsCWMOWnM3
+VPDtgNPq3PKgN5Hf8laKjPnPaxuXLEdOR+wEkavkJYJLJtlOSGO8bAbpvYDo1aX
nRDi5lHesj26Il0x70eEYqnUeslaii1yms4eTZ/pVSIPlBzOxU81xLn5ocW7p6cu
G6d8oeF9WZlyE+qHdf79ss86Qq4yDQUnhEKoIgrU8cV6RqifB1L3/dnZfa2LBy4F
9uxhjtCSWqzhLmvtCZfmjxRKOdmm/925da5Hvh/+MIuCL14ZU1O6bwcArOBradCv
3kspqyaatX6ZUjl6oyZEoCLaC6ZJYC5eIgaOG9ZkJEEb0lQ1tNyngeMFxBo97oED
4Bo4ko4kBUxikoXkHJNfAllNoglynj4IPnUPMT/GEZjLWiXaGXrpbewHnZIFJhyb
Ateo7uXKSCYQmZWu5zsd4ZRcXJVkM4AOg9SHQ4KMPyYWN5B+FGqIro9NgpaAoQAM
c7vPwId8qmMSmFTWB4N18GT1Lrb3CUCmFuNgH6SwN1x4dortRTPxvSsoy4T1SLoY
VZr7/WIepejOYrX/bqpb+mWdRnoe54yve5QY5CpOGJT1kBgyNR7aQx7nvzVl5qdl
o/O67WcSEeV05QV3P7H72Sw7A8cNy2+aV8y+mfe1t9vlw2qhxD2g1kuwd8RHa3gQ
12fTqb095g85XumoFUfrj7r1UgzD1kGxR9234+Qqplu+x1Zr1WIB3OhPPn2hJ0jT
8hkmI5AG5aY2u2C5chG4BX2Q3tz1197z4FHUovd3grXv+Up62mHjqlqwn/V+seeD
5Y2z7/rQmyGI1bd9dhl6Mry0ikmoca6+QjaoJXDLhrJ1nVBw1/z+rZDfksq62dju
pTdEtPAWpJqF69uopIXwBmhyROIfivRQvbPBmuO5XRSCMjk9DfKLWY+FSqUFDRdp
7EprzuKtzvs2Lko5J7AWKKVdpnfzCjXne8YRWlnilFnlIXrIk7kmP1s/TTfiZ2L0
/3RmGinnVWcGZgj1uxI0houad8LFH14wfwknW2UNnI89E3aheRkCKie/Qpj4mnFr
EXD+tZ7e5fXiq4/vn0fMIz/hvaQr4QBDZArS76S4IzzBEwkCWh6pgcIlbCDfdNB0
aakAiTLbplb3l9kO9HRn/HzlPeAFMRHcWwZY2mqzwK7EZ0F76LFWEn0epg5kRLYs
DePRZqJmYNItjqEHOh8MQwptFv3PbgWtAOTDGF495AgvYobsRLnZaseu1+5ElJl5
2PHnXguTLCp7k7ut2v6S3V+mJkhV7+sohLRQXd3crYvtgm7lsQpB79/pUys6sgaO
REBpjl/9tjlWrBUCjGAG0QblgJu11tHPXpqqFnAq0IVqToXthrx6hw9FP+o09fJd
vCHAxjhRVECzA7VbFWLvV52pAY32Qq4iuf/b1X+rQmG22566GMwy3VjQQUfKAmV2
j973IS1mdEHPag+RC49neQk8E+5Lgv9zgw0ZxM+/4EjiuYb2ZtnWZ5sglTzXLV7u
GYI7ERSUDiAkVAe30zcaMNTwW3yunKWD9dOOtmFNqBqO1tw13Wl11zn20+FK85l5
uqJiVGochg6Z0+1jmfukPLhWVo2pzyWO+GIrlRCG2wCRi2EoiUpjX6a+F4ABLReY
/uCESFoG31sLQ2zLfX5lpWwysILkKiuM7ohbnqB96FvnW//OfqHJvzmfbl7WUQaZ
vx0BGRnxRcX35igcUSOT/DnWMPy1DV/9NpOEYsArKyPwftQKS0IcrDc2oF6aFdB3
U6F9MzRUbRyOwU3DXB5d+u1QnsWqehy0E8VAX9iiDmiI3fLDx/6suknhqQwJtJGw
zol4jxICGSCciJkspLe07dbJvBEG6eO2wt/5YGV5jzg4IWo1KWAPgBdLpVc9Jqjl
x3w6WFCjde1UrOLPBA+lRsLteOWagYGip+3dVzTPHLqF/iszjaurzAXzxwK+oZ6H
qZzYY6DAPE6sOrS4h64mMXHC9zvkRsP+SqsCWlS7UUTZv1t05aCxFWYMFzHi8FPg
pQplVchxl7xAuC/A/e2fEa1oCUTO7wboClyAtqFEjY1/Fu2RwInvXKJyncdDXTJU
wKWmIcK4qEzVwWOTdmsqFngECDrvHQiHLUfnYSKygyiOsF7J+RAiBBMrMSR/0/gY
C92JwEdrfx1q7XDmX2bUQPMEGO8KFwp3uCiNZ0+wa/MxcIzK/va0O6sVUPR8yumd
qwpoKMWzsZdtAAYN6vfot/LN9gQbfZ7jevFgOSSDX3N8QyK5Wxs7+1845IyUuC8D
y/t6Yt3U7CytgMjZZgIr/yXYt+dREvKzEz7ZPozVfeMw2exbQmrW3PWdzhCOWO8k
qokNsGJr1r9AocZxct5JcZcJJTyMEZqG7GOoKLyiQfzkoMMDUhQ7T3aJ//OrvsiY
Z5FyGK4Ngt+4BKkbDpoaWNlVLsbB9kl/Z7JZAMCbOANsavwsKVS63MW6YpcV6fIt
XcH18PSXks45WXtA2yyJThe3bJ6jaP0ub+hf5X6xUP3zv8a2c73ocgpFLkmx6M19
u+goLImaMjkWeKH2LymAa/5nMfzs74yYpJGHv/RhoB3fCRRXAG6h3HSq3uEy0F9L
Q5echpPDM7K921oSeUQHXcUzXAV0BoKdOkK4dGnxg/CHo+bLcB3acYg4acMlBANJ
5TqrvgLaMHXGCUkr0Qn37UifgHfMq528Gme84w+demArMd66cqIZ88VnasP2MFVK
oDKPecJaCvjINbmFbjQMN5zlgbQ4ZoZ6YCMA2b3M9M1q36KObiNxaHwQoRS2bS0W
DG3YQDg57vlbQMhAUH0XE/Q+OjwTVP81Wup8fER6kJN+Dv4pRKcAGIjOglM65pd0
qn9XxUWrAebhHg4b4T6ikIVm26ib/RKrHENJbxUD1NPOR2ck7Yd30yPvVFms3VtO
bPRCtqLpuzaNRIuO2tNnjgs+xCzcEdwhy4QOW/DvaADXiAMbWNNevgXTihAxDNnf
TpvYWZdrXhT8orn8PdFKYUixMDr9lUBA/LosQnHbprGGL4It/fjh6rupDmoNgj/X
C4G/vXOGGTb7nvUg0uuslAM348eoaXwGEQitTeub8ajCQKs5b1TWg1r1powyiTVG
P40DSLU0o+51frmGjgnZsxByrOHWmBhqJMaNck+QjdaTr6TBnIDp2Ez3JmlgqcoB
B0FHGBDO88k8am2j/lBoRA9ti4BYMp/qNpooiriecEt7bhW33vCOG0INSa5FoCAS
8+3JHbRMnTLKkQQWZagsTu3uNduxxSjJ2MOkr9BDUAP9akvhMbp9oJIXM7GGX/IB
otK5SCWQbQyOj13sIpbkCXH9lyXPziG6qOAmG2vcgGVaCQISaS1PJg2X3O+RAVKM
nIAKjpbHZhUjZ3JHB9nvegn2dpkQomXGjOsmKG+7wbBHfpuUcJM5o8l8elbjPMcB
sG7fSemI33unxs/PffHjTGxmtmjFnOMs79MLgBWtcZoukgTyKm8v7lvEtDp5QRL8
txT0S81EYTPmzeyYltU1t1ZATVP/5LlwqJt1ZksosM+tTyAYq149WkTK4wySUdVU
yCv81kKuWiI+LFmm4WMf4YXF+EmkFIpHQC+TLYaZ3Bb2uo8OpNtKnp0I5YKlzOz6
PR7IKiLGk0I7R8AqgJFgfDxRmypm15RJe70aoEMOyAPebw47hlcDUqRV4UDXVIGL
TNv/+ROtoIns0O4p5p+uskcdxX0kt1xBYDoIqa6fR4fnKFax6PKy39xf001+8VBV
KI/nu8EqdSV0eQ7G9ojmpCOkh12CS2qPXbP6z2duKX5q2CvrDfi27/S2Ba0zNX/O
PlkrK3nUW79nGoVziaSNVO5o8Dol6/F+1EzNsIQPu4eweAQRnnc0HHYNY2+qNk0b
PpCEgzM6uLTbXfFeZZjMO3YXwDf5jnyRhcBQVpa5Z3yyZyVrin9ieXFy+Acm0xSx
dLA6JGD8F+rCkH5KIKjnwtIm0lnVNVDwqsBc9wEkwiZj2RV1YekDvyH5yOC/xsvC
wlagSyTTMk68DGOVjIEDmb+pVg8mSUuv5wYRzwdxLJZuFeXL4L+obf1abLu5QaQN
uyZuL1n/emFD8bhCrfEj/L7/3RVc1xnElMB01mAxxK56+yOp8/ps/3smD+/BS3Jp
YYU6wP8HtWM4rl0wuBOFSa1wWK/46T5Af2Qt3yrQK3AjoZnV2brPYGI1wKdaaCx5
FzLzyr71aFOn/hp5lgrHRlC3fblA6/I2PiH8ho74hvkgNWUqMHCvY0iO77ye7DVm
G1A9hUX/Dpdc/oPuLW/s8bsVR+yvb9bwMDV+vRqlcy55nYbaEdvaiPeYQup6VwxX
jVetOiiy9EZvntFQBReUFHHXMdT25EzVpky0zIIkygAetOl54Q3Oj+9XMnFSvlKO
g8sabZj9ldWEvbxhDWJ52fnDbMqOzudoYx01NTakPsuslag7A9Sg0QeUknKG9T9B
Cix1M67Nrd8RCMMVhvqBQvcBpXCAHBZ49gORjU7lCnUx9GmOzftzuqbu+qanaM1T
NMRasloZumD+mJfs9Isvf2yzCV0mOQvsjSY5nH8CRIOgbE8GIcnFgWjfc+efFDdD
VJCXMt08gx7XHJ/QHlxY3za3mcBecSMhgz06SA0kBS+SwUWlt6mm7Hmd5Mwz3MqE
+38tqLiJBnpC+BtFSf0dS+EOzVVGo5El9XdpStGmpYAmdfH2YNF95RseOBWEezCY
3uz79TwUPPQEMB+91XizJKNqqyzOb7ldtTQRG+4bIrLv7y89TPlFuwhXxDrw5nQv
St9WiBwPnudBYBUqklNEb2O3X6iGgD73ork9PtmR8AE/MlPHMU+EdBU0M1qu+uOV
+YLsCN1hQIQzI4cD5Xs5k16DwFJYtkZ2mELW+z4QBBEKEG4VVY8ljs60RbXFZFWv
4WLRnJiOdn9lrvAQr83lDKM4Y0LQiEnz4lIE1YZ/m/wLZi7Wc9haQun1m0pa3Vxh
F/d4+citgT1csuDvX6pBWw9V8gcSBfBtsDPnHooklA5LZbddjuAOFgbxSrapNHpm
gVCe7Co96dUl5A0rRT6I8vqeHwNmqaD4FjH0SeTKK3titSWk6KSn3AxYxWDACuH/
Xn8UoFB5IFLw0HM9y5C8F3KFctol45A/T/HK90FzJ+BKt6SbOI6gqx11UR3MENgm
oTQCtssnOVOIWdUa0W9x4MX2zSWL9zEfNHcFo2CKUsBk3y7OWmUwVb/gVhBiRM/r
MzCZt+ZrNzuCOBSHN6Dr0GHOez2N+jC7vfNHx7zHIW7hF1JMQ+ZSMXNx7N27/afP
hfJhRZhBjf+89gQS4QP6auCTzZLtnR1dMFfCmU+XG8qgtu/PeVWrqZtv20D0i0WM
nvlhmwPd90zvTmDG7c3rrodyFuGpDcvjUTLd3WTSpSkvVgkWung58V/PEZMIVCd5
p94BsHbNy+NWWaYH+oP9FTywzlIEoTEUGX5irS84ZxuA0Odz7llUpCi5/vqGKLwV
L4vvayaCGDa/P8WutcXItleREsupZmi3kvjLYBN0ngCAUvForwQPvNQcMPOMHMaE
MwfvGZtl/I0h72j7iRhNLj4yogYzx/XdVlW8+Q4ef9wPRg0FGfMqZkAoIOJ322Yo
fmOT2TJsFyT892Vby0rucMYkKIV0rqAnikWrWh2oloBPfhi2WkqSeuOHILcJWSiI
UlfxGCzEDYFNJXn0wjBpGTsLVSfFyJbSaEig5awskS0sn1bJBEuN0isNrjQNF6FY
CjEVVuZMA8+fHR4gST5o1KiTj8KTw+FuwPDYvZrUcHYPb/Waj4GLY1aRuhS9gEBy
KnjkLE8Jkcv3OJ1ZUZWb7LzBZLTKnlMvIabujK0LEfzRk8Vg0pEl0rkxvjGu4Pyx
7B/1fCS0L8O5q7gkPXZ083puMjR4anEZe9OLPlI/UGFtzGbMHUMguuyioOiOyqtB
aogGSBXnayZNr/Eyu8woksiGgfn+otsFA/1IN9sLkH3plHIAw49iPRwhhQ2VqBh/
e4nemHxvzpB/tAOR97VKGvPZqNwcdNjrYdM27PAyfoaU5KlLD4H2BC2LvazneFqL
qDOdnfRoMj5CtD3AnxxMDWvKkl2qpm1EtnekPXL4nG3HZkkMAmfqlWLhCou5DDi5
JaYzcCh6UorMYZo2Gg/UWyJEuqzidloSLVa5E/lrq+viGindrsA6Rgl6MiryPWKQ
8m2I7k7xf/JD5Dj3J4UVopR/cjkmVbTpZ+kg77g0VLla1dw+SIL9R11I33IUipPG
9xM0Et1VFezyNflEo36i0EaKtgXPPgvdPLzo1ortFsFZGF4Ya/FEi9DBoTc+iPrW
4nbxg5GppdEC8yQ48By0o/6OD9RKFoyTJxss6re4lfn3acPc5nkKOo+UpLQjynhn
j7e3sRa1Yq/LsS/DfFeIY7KHQ3v1g8GnC4tyrhR57EiEZAgOjrN9LNWyJ9sxwDL2
mVrmM2UWAfEd7H9qm/ycEXsspCgv+mFpRKL6Bk12BRdg/yuovRZKbpQ4YViYuhKm
Ym1ljMlWUnzXcb1rWdgACKjhjfc9EJXJn0vnkQ624ApDsru9yw5JfNdIcBPdtMYb
a8UA+LxvTwZC/hm+PcEbGRaCurW84xZP49ZWNnqV7hNWIADbuAB5vsJOQhcPmObb
+pLyusk9aMuJ/UIgmYeMSsQeY0qNevVDdrft3bwn7D3RUItwPj7PsQ/K6PBo1byF
IqwhqsEveGeOtyz8paRQaXZaFPMW7WvIv19Pi3LaNM+4wxMGnNhVCTpc3CdLF2CC
07EGzgYWR11X5jl6DDHOsMrxK6vy3gDPABbJe8HwO9zxAn4XIzpUgYvRjPnn2nVR
+H5q0tmV4NoFCnrozbPSvn1nBv676kMxP8MweJ7lVy7I0UC6WQIYaFqP78ptEupA
nhtaIPbCdnix1wcIj/KeupKDyNW1g2nibMvNCNevRCYyIjeHoDGQdDsWMBARwSxv
RNTSbr3BYNgREN3+lxDY5Uc97Tgswgsv9rNDSlqNqAnVxZJdyo0mjKgstoDdgzPe
ffmUCEp5RcoJwkjZCaaJ/aIysgjQfchS4H7X9UWIguSSL1wRsCSMnd97sowOEesX
o7XyMJd/TQqWc6IawoM/zS6Nyohxtg22eVDDR/uw9CRMI0jUtz6q+xXFD/jT2ac9
Y9afinV8P/eDaMD7B1bbsGaEGskt8w3ho+WsnIvatqZlmplupJDjO7F/gqdIhtDe
cZufWm4X7YZt8hhP6InWlNH/T7FBaNrJ227sbUkeUWf4pxURGBNgBQJU1WtASpnT
oVpZ7j0Xbm75lKlHCKYWUQa50nJEXObCGYiifLHaguGcv+AxFCm6G/aO58XgGQGp
wRDoF+bB8De49VVsZnmwxmMt2VFRAx1SZ3B3qV+ZHogZaQQn4Q6nnVYNsDNeq1Sn
ZQZvIObAHSITbcSYaUQ5VQggPHAlSdFBNRzC8AjYg3iHLWhGnDqCAMkPEGpb4iUS
TPKWQU5i47CIkWf9Aq4HecxdThxmeLVZQ4PKZKlvAn8SuBGEuG6ZIq6KPPJLAmfY
G9z/NlzD6u+dV+bDoicVk8WvH2LosqWnl7dlqVFhOh7ERxHsz9B1POlca22wkq2/
TzfsWFAvRoOBcqS+0vC3y3Y+2s25f3A/cSSsrHXSl4KZ7rkGG6/t67zal7VXO0q3
1rTtmU3womBEpJmioNsenECMNlK3dugEmHT1y5YE5QSA3tYWipO7lvPsnE0/uDeN
27S0REuBQT37CziyHtE2IzoHHb1mc+GUk5Ws5+0HuzifatRW3ZgsrSl8w8wzJ1Xe
UGitouFX/lf3IggSzFyNTjF/dtO/73zCyBgJkGvrECGchwGsEfo8y4G+6qRjQCqi
Udf7zBfpSifBl4M91hZc0qV78gejzKsbnaUmd6feBtcCUQRGdIiGLJxWQGCWqVRV
VTXxmQPTTjlgJWqVES8EdqTk0K/WyQQoTyNjTY8xZYr8MYU0L443qNkDOj90dC7E
6Yxvu4u7CXzRrla1MuNTdiKUP7w0hNV+DqwjEkPLrAFxX+nd17JSzc1pmGw+5kk8
OTY/sxQgDWCoIwpcXR8xV1Mqu6Ix2aW1NZqEDTnvt2aUH25bKp2mwCi6epE2DlQ6
smWYb1OUYZidO5fSOudG3zEul7qXzeoMCKBRGDqvEcZ9QYql/Yjs22Zwy8uEIbaR
xFOh5xV9XNV9ERRYRB3OfQcf82Oh5tmqSImsnehZ8zeQeXWuXBFcnSdg+N6LWoSW
4M0+L6YA6Fjn88NBDJP8QrXbo4SEvjwwC2qrO2/qHkLVPGUiQnERcEGAKaA8Yy5q
scRSiL0iZPr14ofHqOHeyETP0csNUlV22GhrSD2G57UqD5BPdhBmBMIOxj0zU5Na
ANUfF0VvpYzUwVL8b0AnuPs0zx1wUVefPbpGYnFLzcPJMwPY/+oEQCftDjCDlZoe
f7iJ7N09vjITEnwzBMzWJbLKB2udfDculq3FKb0aYRm/tt7FcaA903gWkbCUwWrN
j5sIKJXSMf3W/80hEPFN5FdZ+W3SVELqUD4F+H664Qq2/mPipZ96YYsn+MhvLkX9
VRPN2BU7vWNxdg2h3KvA0cW/xbh6M3+QI/8UondH+pwMQWdz12CyU7Tj3YwOq4ax
fATqnGx/y7GBR1T2O2dsWaiDPKMNw5YfoSV+HqMArqXnLd2EhpDwH4Ol7FL9QTYU
v0RO5PQAuJsoxukQR6kBnUMXOTvqfa3e2LbiiDrEKvi4GqyeGd8H2/Joit3JSjo2
zLxNEMnGOotKnBXLknKZMxGKGNVobyr4oGyOUYd7LJGFftNbbi9EsZs7Dhq6hQiu
cq0V09O3eIN6ZbumvebW+f2S9lF5urAJgx06ZFPw05p39F5L7uppYS04UEhWVkpz
c6UjejLK4kDMV/UWSuzeCxa9sSENkaQnukusuANEG39ZXkkl6YxbFS/hqaQ0UYEz
WDuz8dKbnZwXchaMNqrjSKG2XK83wQK9xQP78TJjQbLM1Hpx2lphPZmVIEP4rkOh
XDDkwXxAtFxnpQzGbtdBlG1hDGd650v7Z1QxWnM6xFlOr4MzViYDExwm/LpOZQz5
xGAxWvp4LkLriHol/oGEJ11aNXzqcS22nBgXQ6gIqOmeRJd6ms8CqSnIMxpVCT4A
I0vYBubTdvixghKJZ9VmTFjHretE2P9l7iHLGAA2et1VwUOvryyzivJEIhX0vOcE
fVKjHm1+dgz69ZULQtJmHcqDHMrwmuow+vCGcm5V45ILira9jmVyePQ2JSwarjm4
bveCQpwYc2kPR/mTuRCX/iLRkOz+WMTKEYC7wM7x3MKOY5+OpxVHPUJcSRcs64dW
8D3AngNjjJzF6cwAWo6QtgC9sDJ6Ejog2gU/Jvq9jrtCTcbIkEaQE5peT/XjimWj
g4PGbbtOnhjeEXYuOIsha5fk3lh+KokGytAgMiQuvRj1ip7PoGCWC0+7cczwrjLZ
luAPoQ3BhHRlgPyyGRFqnYhy+1uuz7tIom9zAJc6qA5ASmHnJP/N5X7BPcGYicFY
G/Ts5W44EAKJ5kHlqd7hW9usk2N9vihDLdGK9eG5zcRy8PCcNgJ5dK6t1pMN2t08
/uFiRlepQA+pXSqKil2WoXlbOw7+qh8/f3XOEadciMwJRWbg2agh9Qapnls286tJ
kuMuzS9r11GjDxa8wYp1UUjrqiwAg4fpNltVmk4aK6uMy47SLUPqDS5j2fA4UH9I
7lhAX49kJgYmmRdJEwpQaDcyautznQ7+hhM/Jru3+2oZc9OL7EZiFEgTPPtaoD6k
+Q0nFPcnKYmcF5NK97cNoXi1ApcJy3VjPVCv3OYf8tJI/EU0Aaf0MxDRwjGtVQB7
n0uub9LX4ZxVNS1EX+GuhXV/G9BYBjJTyTbxOxbVQV5GYTK/zPaKtcDpuspL+Ynz
4ZP9U3mNlQeNX71Uu274hMuF2uWyB2JCsqzdaBuJfr6EU1nZ7dHiSDqnvcom9PJH
eEMHAwA/5xdiiDXTt7Ndv8wVL9t0DFTaxkIVLjL9e6q3nhTIpHsD2DN18G71qtyN
jsELln8YwVJqneSb441saUy7IeyTUSEq4Z0ZLKVCLT+B62DDGvPSwwVpZJ2UlmbZ
4m31f0Wqv+ygxkqNqdr+43Vbna/dVUeSnlcSIEFwOFJ07fI/97Lvp6UeacetpdRQ
e3nZPm5wsoJPf7sxYkS8PDeMUwa/pm8a5iHmO8U8YJP06HNEYYmAlaoNPQguj4B0
Xt0PatbD+A4PbIgivlyRynywfn9gkIGDX2TgLx6Yup83euj0kNY1v2p/CtBmqbFJ
4MNUcPy1mSjBhWLPVPYBZK0HC3wikeahlxnQrmbU6OsOIuL1kcqvR/zfmA9oGPbL
0vBUn3TPbvUh3rsgu2b/3y0HRG02WVZgvj3yQJEVlUU2WNpfes0QQ+vmHayHt1Ao
kS4OHz6WlZxDqcj3BRwAYCYTDjYQKeviUZ1K44fgJhHRtabTMSw0zIm6POq5/R/n
LuAkY2wozq5HfHFkyNK9TeZOC26Xr6/NIdUgybhTdAbAu+N5Z0UDKUe+NDMFObty
Y1udA34itRti7GUi51pNMoXamwmDyOW34VFq2spYStIWL11GB8e7UWOp2XZjAfD9
iJRfEGW9H1mD0h//dRKkX0CSb8J4GeGCitpSSikMGpP7ysKgKwTqlqY4IakGS7YN
z3TghQmHzOZP/bXABcrrrgIvA1qYBE6x/wiC9jXFyAMdxn1d8BpsiQByKKHlye4Z
IKwHkRRxw/lV134v/BAH9FP9pqzklW8MOefx81v/j8gDSOWXQXfFwK4pusBkgVml
+IbjWAhC/uZn1cUzB06OLWGpWUCgEV7KUm3hLL2I19mq59a4oAhlBNMvVUngyxyj
yt8NtVopMhe2W88Crmn2uZWkx1RzYU+K21mpVpBjY4QBuzdCwuTwBxDC6HTo7HUI
ymwhrsrF0VR/592YL67hlZE9/wYYS6EaEfGgcavg2aYLSylhSmdK+HnI9gZlZEfB
8sb4rKEFP6JmltdLqXNXdisLqSEvL+tKwvZmndCJO78OsS3FSIzolATb8uofH0D4
grZTJvs3+WUgJbcQTomHYtP2K/XoXAEHRghyWk5372cXCG4Is0JMehIx8SrkTEWj
iIrIuSYMXEtU34uVULAkyu5R21h9aFPmyt9nnbsWqpOYh51lh3+fLQwAnln7qqUI
+RvAkkyBZ+RQiAUHlFdV3eADLpp0bnV6n7wyUFgFGr8M7EWqyE7Zbk5KG8iqIAjG
k3/jHyT639QOHStgMkKXEbnVMlASv78NeypQgarT68yAsLhVONi1+ETdLvk/0/O7
X3Fz925McWGlyy0efdNtqacGiTdiLmk2eWELIgFvErsOu8JGEbQbmINvBmcE8b8f
azfG5CTYXcFq7HIY6SZkrhbUZLFSRUu+nxqHzu9NQoUEKcUMmpbT5xvBRC4/jLla
nQAzJPGPGTzIQXNs/H0jSG9aqx5I3bSY3wAg1PHKzz2vy2RjEL+Pm5BSTmbWTdAO
YvCJm+i0XT7hjnaknCIpFTjXUBenl+LT0QkcHUQFRoQbNRR2S1PbiKEi/2RlGZVI
kzcJDVW3WiY+T/GXEjgzBXIEMNOjWCEUxiNG9mpnak44bAZfzHMULG3TSidd2aBx
wBxpboPfQVJp+XVSBMauZiVo8bwtI3M7godpEZYJO58/2DcCvACEslllZ4HhqoUS
UG8viGAJyh42uiFqK5XfLdQ/Se75IIZ2GrBp7SULfwAmbXhDNY2CN0GeRWCk4FOD
4BKcnu20ho6RtZT21fNtvocwAA71o65Z3uKk/5RQgdRWx1PYkbpyTRxcHegcX8HO
1mxHhRsjbgO1FEKw4ZG3HOorZj7JPvbxjUzm0+IxN4IePomjzCIB/3NBHXXe3wBE
CdjTS4XLP6ax9hFjkttBdnocT7jv4Vkgl/Ip6gWmZDl/0u5N2Wu0v+E1uSPW9cID
n4BPVu9mkR+1hvtNGoFdjUHsCtHbHXg2LWTpGk5OslUaxAwqGjMYCwjNjnRx4LJN
tZqVCyYNYXUWiRzwRnNUJXOkj2za16rBfBnTmu9eoie/EenrojZGgZYeOcG2zTVp
POHBYVZ6Qr/6qZ/kSSob37XwoztCcnsNl4MqA3te+nlaFipQ5dW6dTNMP2Hg9F36
fJZg2+wf51KlpvmE+EV25ODFoXvlk2cBbNyn/oLKPgqFyzfbEEmumAgF7ibf3+uE
lJK4GjQnG1683iqm4anP/Cg8BBRyh8zUNtUi9FBoI65KbufgArmFdwpkgK4rQZSB
BP0J2uK0GqcawRg2k7sBF/7uFB70uqDWTBf9w7LonE8Djzhlk8R0YGCj0PFeKb1d
CHqmy27Dq+p3qh5N36M5zCbCo0vEE+UQKLgqDTkO1y134tl5e61PcOyjlLewDiFG
ascjW2zg7XXgJUdfTyEo3k0AroaKOZHLijM9QemYCIqhFw7u2+e53iTZ0Fwe/tBR
CfGDXHXF86zbNgFU1lcYLUFEGLEwOxouNcgedcsFRZHNNKHq4MdIthYG3cMP47tf
Ax7KsB4FnJ+ZygVxVOtfs5j7wH5HGyKiRiRr+5MocB/QsoEj0QxjlE1LtfufmjOl
3k+ZpNKZE3Ri7eXZ8HM7sHe8ZpVYTdzHaR2JOAc9oGa6BalbpuZCygFP7T78qH7f
c4P9s2h18r0dLzAvw3zawlkvlMij2T6bliND4xL/c5+Qxmjd1Q3JulGkQjT7MR/+
KLtF/9MD6k9S+r4nIvkGACezcLc22l6tw43vH6pTPAx4yP4PaIAwr5kcbD1SaBUR
S3RQ/Pp4VsjGW0DIJ/WhH3ov1OdLSgVKbpsGl5JEtotSrG/ngfayT2jB/Vf9h/bu
58EGFFTE6CenUeHxpOs3qYIIHTvZm+bbrVvtal3LpItAwgO43Crjr2Fp3BLbm1F6
UoWjRdOR1PSsXhh/uf35XZPbLyhbxsMthCi2zcyj+5nXnxBOJml7y9r0N8phNuid
ubcjjGKLgNFgMeawJQ+az7fO97Wetboa/dHhGQmW7KT9Bj+nPm0i3ZKf+V/c1nhx
XNolqFT2CC3GkjnjKG6ZnSJBezm3mx5oT9MwRnSZ4BfSV8duWrXsSqBylOIlQsBf
TPQeLMLkvkPtAykMKP6s2N6epim9ylQ66/qz2H/648CoSW52Lowiulj6cJN5t17X
zqrxqRxjFpscj08UI2k/ycmhbDbFrPEvXX3DgfMys1zo4KHuD8swRvxSynoh+bno
dwYdw52tEMU3X3x2flYl7um4l/9dRMmDyfpvgysWsclky+2LafjB4ZeGJdq0Nn2U
ZwKjxJ2h0z/xsNhivaaX62K1lLH3D54wQ+wRU6UQYv54bu9lymKgCwdD+oqleNL5
UNCtYn4etFa9lIjtqiiJ1jwFuB6eWEHbRQiuq+kWUpQ5rBhUo8boLYuBdUcI5Ofa
mjhwvSDpShTwj5FNFmmPoPh1t94vmy5XUod3NMnfcjmTriYpNHDTiGrcCJLlCG3Y
E5m2EP6bjkNTLfz6DdTn5mECo1UP/h8dG8PunWshV652lDteXjb1QC6MfFOzb5Pz
/5DHwyhU9YlOykuVVd+HbogQH3ieS2N474zWzk5wXYF2UPAatjxlvuae+dwS0kvq
Fzi6ism767f+cAp6meBid32KPisspSNJinvCBAyQl2muUZ7t/al+AHMkFtX5Wp03
JpW9/a5J/o70CyhyFmy5+BxVoAGJCAAV8iWxmPdb02yrcArFz8CDA7kegFXuTGiu
gQRjNmz2PRhwSmCK0LoJ7UXKiL++N41P3+9gzpyiWJfM4wlGcvD8Uzm20uwMud/2
dJX7IdOGryTzh7tjqkWZE3Kk884AEowWft7IY6G/PcwmDFn/URhu/Ymsp6SrRetJ
yEulKEzF7Vv72fZs7xOmJpOqWni7Rb8REcTdw+uU05+EqouODoaiLFvQD3CAEZrX
MRQqTwVbB++pnlu9Jo7GgNmcSmSm4M4NsmW8APd5y7UAlXNO4xgpSrN9MLJ1PDjO
OXIW3gjSo0h5VJm56aoIVYD1/wB90LZxVhvwA+HsokTa0m7Jd9rU8oonjLWor6wk
8ETQCA7tEQIZIUwNX1uIcWgASUxIY3pFjBoAYddlOOxk8UFfvZPLrLcbd1BUPSnq
mlcEpY41gZyRE3z7tv11sW4GR68DLDDK9F1rtL+VLjaaUc5qMoEREsTVjsEW8fra
RzwO3Yq06DlPMsY4dT9DlH6Gynf/hsZipAd6sV5VTT5ibiVR1rn+upBgQoooaL4C
wjFY5T+ZKGflkgjiKVSEIC2LpiTDyYPnrC0gyHmdWNo1nK3aP9oJrwwNYOjDDiSb
4mkNeO6wZKMScDRGAnSM1mHPek1Kj4q/tOoKUcKvrDfkhEO1F64yAJ5KaRAahBHU
7bJRMIq4avgSPywFlGpdcIOneOZI8D5dc19uLQPAF94F2UcK5revTqAzK5GxNUMO
jtjThpiaXSzUMM4TJZxLQd2jn63/i8TRDgQaKFvzK3jA4EjT/K2qoI1rRnsPxdL7
hiU8e9RXeeU5tIJhxqDze0pzcDNL7jn9m+rkDMvvJg3uzRM9KGjcZrU0v2+iynVB
dqxL21pQkwJTBWRhJ6VPiigR17vliqaxOVuE4iPBRrbsHG5Yx/pETrJJSwiA/4y6
C9QRQ4+NCnkGLNaxKwM81JZl4GQ/1sJJvSEfA1odQxUxefaS+gGlCNVIyrtNIq05
/yAD0ujpzgw5Ad7DPFBibu5X3F5hKgZMIvGHhBgmtmpJd+ei4nRZiUNuoTtN3SxG
nlpUYnDhs57v+qQ4D0/SZ1d32UaZGA93RQZaOCZFP1h00Dco7UEoR5SF8VTiQiu0
Zz9S8IlrH4VRjU1efOiLcOVyoajDEPvSBR3rx2pIHEHUpvKbaY/VRfiY5wLtKYWp
Qg6vFd0QcNR48XGqLa/U6EOYXSsxlJJb35R9SYLsxQi4qlLriKRsYvYnLGTnBD4E
JwRoFpquG2hW2HEJYjDGWNyTkvEKJ5smtxKyaeEUf2oZoUO5ARF3d+JuQ3eE2ACj
b5x7EghdP7aNlRr9Y3mXysHPJrybSP5mC5Z9lDec2XA6tQrQ3/WYBVo7JVcjXyoV
iWqizWKgIKzSdQLd06ZWIn9V5OjcDKrfGX9wRSCwi0uOVeLv3cpL7wgC5KauhEa1
LdwKAoWpSTclwMzTjT2cmPOf86ASbAMqGi+Vz8V5vP+F6+F7HKdHhI9nMQdeSqYF
bfwyXcgwLzmgiLT5yX+sj1siwfBPKJkSZwsKqZoeOGkZhvAm/8iKoyWR9SPzCmJ1
AXBGSGeg1K03OT6Kti/mr92ef/xtypBYr1pgN/l4sK7QrhjaGf/E0ZrAfkwP9IOD
ilPWVteShnStPFuG8ZYOCzaPC5xoQr0mQY0bq37/2gfkw041mB1NlqVUId3Tnlii
1NNLKiWExmklOLCeZQn4nCTcrWmqrYApOhf673GV5vQs6l2P2O4IBXjQxAG9VpIi
WBjRpexa0qQ4sPeGlXDlOoFFemPmBZJd/+SEnE9xQfZLugUaT99dchmJijc41/d2
LVpyVcdzYs56k97FjvvT/POnjbeRpJofI3R5rq9Q6HqsgwY6nCwPjiThTwXz26qG
9353VzTlFfqc9K6s6zl03zLrF5EvRDEOKR//QYRVycUzX6v53l3xTVw3GJdmhNOM
egNThli47/wjiqW28orX8TO+eF7l+XTqm96JyKpXo5pjI5O8+xMnjSjb5RhkTOxJ
a6Xfztq9zdLZq8eEa2lpMsf0ia/v68ian2BJKRqKOSK+R1DoP9IzCLGK5iZcN/yT
WII7IG2JPXCCjt4sTGb69uoewnrNjMhgqZCz74PUF99Nn2KSZKNUVOZbDQXRdKqG
kOS5r9V5qatlJAolklnzzLKVLGblNCXPA95i+ZdhQQDPF2WkRQiFrRzshbPBgClN
JMm5WvIZqUb3+oGtL382ldXGZDiNyL5NbfQzfKvHNJrEc+MWMTrBA65dR/vtc04g
kWxrya+UJ7yLcSynVAGzI6iFDkpdjU3H6PHvk2W1CqFnmeY6j3llKLMhB0fPcfTR
sI8GRqwiOLjSqI0WzUTOWQfwKiqobR7a1rOn2I855OaP/L1Ft+o2XRXdnx/Y0ieM
DLS7C9WwdBjJUJEVFQr6mu31bUHQIHcRLCIslaZ242Pv9/l1etPGqGAIEmTFgilg
yYFrs/3Pk4aJsZphz7zuG4eTPzSwg4jixNLeamRWK+0q822tO6BZCo7mRD1YXYrb
Zv69RqT29Y3nj3FB1pABlifN7qrxuqNsG5azQu+rDmh6RTZybFVjfeFmKyruYVan
jc0jTCeXtReql7G9STJHPGx5vq0SPvCYC5jeo5wxB59k1psPbJsB+TINTEmlZFiN
VrpZJq+O/TvbYbfJQv01BNXVdrvkP1cTRGOvuCcl2JfRBsxD9o79VTRmNHewuV9f
SIHNpEgxG+sNV9++rz5OE82oqaI/4qZmurqwShE7OaNHf2BiTJTc8mF7I+2xOP+2
nSDro6l7QwPCGOkOLOTsYF7y6iN6NMpgalyvWQ3KVccYyoIekN6dyk09yxJAl1su
iFCdm5KRUwWUNDpENJKSf5U/iJ4riQSdEE3PYwETYGl7KOyQzDpsh/riNocvvWcz
aAfjKHZSrrnfieu51Oy3zn+NEC+IaKE+WHTQRMDobS7cGeqjZpY36tK9r1B9xHkh
GzIAYXjj4Fh1rNit7HPr1oU3WrvE9t0nIxN/D9u16i1mTDgURmQUlAhTD+uhu9d1
hX5f0zVLgEWer5z+f2QDoOAiLB03k2NlGqacdhkw+eMW2wL6Qm6id4IzxolMw1ZX
AON05KDOSRMHIva1IE94CPHadATrH8mCJcZv3pCK8Y7pAuVLuCeCFtFrgjyglji6
C5y+Ofi96iR0OBBSRgI8ExB9Hjh8tFE05UMunYwFPw2mfGKaATdYO4f4NgeHnzpv
QLKQ17zMa8PBOdWOgbgwbNRlH2/qdyGE7Ruo2nNKQ1ajGRGbY99s3g3Me6PXocBe
3YuIfDI1UQjxANo+FTk4A15TEh2gpyTWq8CENTT1SVg8fYsHC4jr3MRtjUoRovmR
3aF1RYqRIAZ4kXrYGF7uAk+2IflDtage64qzopvXhnTyH9esfb7HGdxv7rpni4XV
FLs0eGYa7zuPY53WAlMrr5vk5nWRmhmsw2qj5trKk8B8bSiPI7xoP6duQy72G4zr
UH77mBtcARg9Qyi1CJ/+JZ7DmwNynrLV0zdj04JzHpRp8vTPPfMVWWkMutpcFOWM
vgH19Mu0AZ7tnCyn0joxY13MqFsYZXFvm0K9OzehIvHlQhNJnwPr6xiDPXFPI3sp
PmACrVKJeMGgD9nfu7dn8mY5jtIYNaiVta2HDstHH95oCyQ1ESwLn869aqVujsQP
jxFrWCDY9tOgLu8u0awAvtM7RrVAU1ocUHKnEjlCuggSCYsVVI8hCKfMntZmPc7K
HynW6YNKRTE+o12VwVYiBf/8YERf8KGFImUZHaRpVCQhF9RTbZAi2+pOxtUBY8DU
CX9WfX/WVnVQE08xL5ZUNu6k9wvImompd2wwiqdEnYNWGYv3NNcehQMyR19EXrd4
dmxi7d5yekNAlQXOc7GV+BTUAQWqoiJmQvVe7RRkNaABwWhZZwAK83RZ4oNy5tfH
8dfz1h/tRiNVTsIMZ3IyLquTaxfU/QMNtxsWpvjxT/OQQRK8+WQ+8U4Dqou1+nHE
eSRkzv2rPyMtvKJB/ILtjWAbKERkdgMYos10ybciQ29ThOdi5+Qj9Ve6UW+rgfbq
4iHoJ353/vkELGAh8MDFD6YbszJTMChfQylV/0w0GDmTZ/KO+kDe9tQ7XXZGzNG9
xreJU8uPadLS53MubZn45QbvqR3nn+CvknDslGnhkbsIaoalAWLWDfe+wgEJkhiX
VjIhW0xPwtmnxUJ6gSuuBmQlP5APHz3QWbPCKFkoLLU8jHvjohW+O5nSHH3ve42+
iHIgEssvYIhKIPLW6LC5654k2QsxL37/r3fqxKJ5wqeafI3YZdxXv7fQx5G6SRy2
2QFxN+njlAO9Pe+Ey8Untp2QvvHBvK+RHUWc/NLUqHJe/FEZ3m1hw6VCbzTDkafZ
RHCdyzPtd+LRdcK5L3ovNtYBdfHhLd1IyzXQTwHajdXi350GAKm4ZkLtD1NRJOkC
ovsupMu6TEz/sn+lzjy9W5bn2b5TY2lGmPSFOt91kNnxHnbX0fWrHjFFRDZE7x5m
ZiVDLjwN//Yb5d5vLlZaErTB61t2pxevDGVrHymyYvPexaec7zJYX5gii2Qvu6fC
OOClr9dsrAQx/6BocwsBco40NfawKpIJn1crmZKUoLQTKA5l0NLAgIIrp/6z/qY1
+59r97KTjKfehqn6CDVBATSxckeSrW217x3MKzbNgNK6j1XVC5zIYgQuVUqoEhWp
372Lf0PwuJclXkzQcX5nmdWiD45gyES8XWZttio336wdNcpQk7asObpConx2x7lZ
4Tp5UPu+FJHx7ncF8++MPChfN/bsAaArg1ck2OoRCvDAJNZet2jQebIoPSiAvVLQ
nnvxcnPqNa0D1CxVSi0q9WPVn8JjOphBz/Vy1o7GnIUSSGi+1aBXlG3xdiCxgbHj
CG/9KFhisufT/x+rdz+H5sSvBoRS4eeX4yubSqIpKwUFuaL5ivg/iiPyYHIW7MM6
Q13YItIyyNgvKHoFFAmK3bJasO2Bdm/iwp7SCW5IjdXA+lL1V4wgr2YnjRfM2mbR
1sld1kYru+6UtlW9JXa4d1pMcKLBrnANrFnkzOzGrwAPOV3AlrJO2QE7+LHj3H7e
Oi+7aGHpKZLIjJJLhbeDJafcve0EMkWdjhRaOV+Yd/5Odyu7ZODydTvrr8nLjJ36
WMRWsPDjFCWrHPbK78F/XyOZ5n2jylbeOFRGCfoOsv8mF/1fjZ5AJpmUjaOOGHam
I7a5S4/QqXAIZZ6Hl6Msb8nqqRKFJ4BjrGhqcuj1YsmDepQAEt7ZXxIMyC9BGIvL
DFdyUslaMlRquUYSWBNujEpWSI4lbRUHkwGmebZrwfRrHRolm4S1h4j72/XxYClC
/dNb0lfz5Wuc4CmDlA1f6Qb5ZjFuOR+akA/C/hMFBH5JcMnH3gB+RzsArDRyWAaz
W4XFpeGspsq8DMqzB5v/891hNRTra75GyrrpZ9pY0cM8lgLxMghq0zwj6kD9w0Xi
UOqmq3XkiUlRGlAL5kfOp3z8zVcybRBwQQySviwVoYik1dbSANZY1UGXeuNcLFt/
DXJn6Y9u+dYJB2R5JDfZnLxwYCabNkThAddTyAUPOqOTMlw82wHy/y1s5PTTwkXB
4D70Hh2YiWE20UHRw58F7Y6ciQ/qCvynBQQdRluFx2kr3M3+ZDmXGrZfKjzWCPQE
jj1XR3nzIXx6k7hHQ0uqsccdyg6bun2vXMOWdvmRkkl75H7nNSvYoQCROroirgrr
PAMKk0EjI3jl/ppNdoKTaEpq3riSU42CVu2zzuJjT6GEI0QtnBTIWNvm32G0FMR5
T+OHr7U+ZICV+zTM+mrJVLCWJ86+DPHovs3op/mZY1eyy8OfHxnO/GGS5QmvQ6yV
usJdABJEaOPDWnkt5C2DoTvwqLuVeQBPk2tuClWNzP9ThE0kGYxbv1m5PdQX62He
lg8jq6Y3SDbCyxMkc6PT82ctmFqfiMbt/2rRB45cm37X7ElCvo4LEU73cLaHSfcN
BA4Kv+aElt5jAhtFNcMnGtPkV6navC0cN0zXma/Dufnue5E+5ibeFpfkgDX69Zrs
esss9hRoUxWomsubeGZrFdo/Ct0D9Cm+Bzc01zOueOOz2a88LKLR7IL3Gsy3jUBn
LQoZZ1MpYEo6aWUi3B8hWelTpnz/bD5HxSxLtjfperyQ2ZZwSVk1sF7fTThXZjJT
SbF/ShrBrACDhp3u1WXnBnVcjy0Cx2gtQIX/YXdjZbY9+hFT1odylXA2XyLCWqU2
nYmxqEqkIVS81DnGjFFB78bkwDLlAhfHOZkdCZJJO8dht/hPfxdfLHh31DMO4om8
1LBeEHhs0c4AFAlL3D3qDdnUR6h69fipqGS+wmWf4qvfoiTXAeHlSgNz4PIqj4my
ETE2ytwNqdqOuTHmLP/FDATHTjBfqXcAOSCT8+I8BmZG8PeaqPJYl+2NO/h07278
OhSOOoRWDqgTgT4NeXNfI03yHxO2/CHtgQu4BJ2JFMSBnjD+lDhaAGNuKwlkcQ+H
WaiDeD+rE7NsssNYU5+y8OYNE2JN2Z+fXDPUDXIimJgVWxYDYr4d2PlBi7Yf+eP8
JmnYvfRtEXw+8ZgD0z/mRf2GvGxzHbUDw7Mr3C1LGeWrtNGBo5dEf0/JwVkZBDBx
QmJo5OyNQittyEmGmdCWfTjy2E2qf57K6b/jF80fPltMHns/zXOjzx3viy/gLH8y
zOoC+yaa2JU05DN67thaAPfc64/Haei/yZNk9mYViwGSO05etuC1WN4JB2yd1jAP
r3MPn8LDhpzThJPIzBOzEW3qXomOpbsSt4n+IJz1+iLS0GFhiTl4KP5Rrx5+pjfi
TzLN/juA/YjpraG8pSdKSVMaCNgKYC/7Yzs9XQv7PQJVcApiU5S6q4IfrSF3vjoy
WAmqhqYaeqFkKXZFi576KbTiLOGV04EnUhyAt/s1jBPPZGSAxxb9vEmkKlKuYPuN
SKzDP3C3qXBDyqiBW4pZSshhvoobWMh+a9EOGjmqQyjozbF3Z2j5f2izFUPEVQRm
YYQo1x++ZjqlgAwu9rWOw9dR/5eXyYzms/vJR8yMHiDIHH2aM6GjtyyrOyxCLQg1
ismTTLQul2KgluePMvB/X7LC8d5TrRhfxNyQs9IAceUWK0ugQGZdmjwoBl8wBmB/
38T48cdHpQ4tYf90POXIm39bnXel1E+84cWUDUlkQd7DEGbFXYF0ALkPtd3Fc/Ec
OWm9AHdzAZDuYPtcgGRWYMwfJQIrHYqHmOSBYgjsLS/QV2KLIkQXMb6XiSWkTbRF
Q72tvOMTSY2jdbXtobH1OSp+yo90GLAsEtXrnDE89ozoYpspOTBL8NosFqS7/blQ
T1l8Jw5WOJyjB28LBIuDAm08ypHXVbXRqAmr59Gh9ibBvY9mMjSo5sUTEwkO49Os
h7MsuVA+LZZtJ2JSWxuXbsbftIr5yiuPDTJp5hkiNv+DBIM1ml+b3PGms5M/+Xpp
STRqZoMDVUNskNIU71FpwqRz85PW9QGjFZRJDoRJE0WMLFSEaLA6c6xjfDd3fnUv
7TN+mhZ/o1WxGCnUghXawTuoNF9OeTCbazDL0teSNO1Im/08B1wepqKbUw+t96WM
ScjTmkT8opylbPiBk+/fvr2MkoLcusnwoEQeTQ8ME0WaDKLa5PF+pljwDDYS2hNu
SJkCJtoZiF0dSZqjCiX/y+Nm45kuLI7wv89C1Wb4NLS2dLAXqj8tsbwHavQ4M3z/
YWNCOFcyNeyFnL2l7NGj4y1M3wN9BMcZpAMlgTBK1Sn2L3dQ4p/do9XavAjqvSzu
kMveBXdn/YcTCtm0e+Mnyn7ZJu/4WZXh/8f33XWWFlNFnS11CX4aV23zBFZ9F03+
ckkHT8CtmtvGmwJRx10mOeutU2BUxHUZjxbTa2ZMzfa54SKYM5orwcudKdeBHw0/
dBzNR8RuY01u+l+TFUDRdTMIVZNEPxFacdfHZwkQEDcSFKtSHPasFBpeVclqxerz
KVrkcuH9O3Qm8Jmx54erLuCTuC+Mbb2KG/E0p9Y6NnRZxcOyxcDZ6TDpoMSMJ+QZ
CEA8XnjEs733C6lkRw33ZQM8NDCocSzf8UxedDd2OLmJn5mZchGUb3EbBYJLstJY
KSmj/uTDnjvnzUOJB5lB9CDLL3ldqikIP+UscMUHtyMpnW21hXuHupHrpcyCTpmy
JZVLhEWf0Mbw7Ps1rTbtHUmQiL/BPr+J1oguVtNwyoN/p5BR7FLPSG4LkXKID084
FqxvgqEmLaKPYHi/endCBVnAHHKDEAUS1ezb7qRRiiDrOE76yDYmP2au70TjQ5RR
Zq1kmfqpoRW/QzBHFDrjfWBBuHEackh1Fo/X/jH+fQbJWYpoCoIqBNunsbZsomJp
VcIwGEpNFMR+drTI1zKUEjYrsBjDycAghAy1/xoz8jQFD/M30DLiFsEUe0quFlg2
gnKIgNyb0uOxUp2Yjr+nHuN868nq5JW87CI8y9GGTQqGVin9vPDwnDQJwE2O7lDn
+SxpDTiYVs31U2f7z/B3NO4kb69riipn4HdZXBQyucAXhu24RflX7Gh+7/+ITp3k
9TwRFnHsd+FN+qCmFmNb5eBLIEE/+kcgERC2xwXQpI9V4L2zaWrBXAGUePoKBPLe
5/PO1eB0opN64Vd/SE5ioYsxKDFDzP726eIU3OksPGLH7sAvu7yz+111NQNIxV2V
PnRIZFtaW6JX6G89oTqZwWfuHlU4/cPFA3wfKSopuZaawl9vbbJVCpL98s64E9LL
adHbKfCFbw8kPb7JHUCyNdETKj5F8VRa/DlI9UcAsO4/m+vbiShk916eS8cBqyJR
mE4zOcxhrJe7AqS5W3pYaISt1fRvF/nAd6/crREiOyWxsgAHxA4c/5cpWL4ZOld1
dzM5mV5pBRabiT6cky+TR4cU3cKBDw22Nm28J7QAdDNmPJoCBgqu+GdvWbICWakh
P0UaLMHbTYCvsyrn+Je93zAW+tkab2flCF/VvwZ5a56YvNk8ArLwPZ46InDEcp40
B/exq8VbikD34pVL/0RJIHRE/Z+Tw2SRVaNo29Bxs/+KCp6A7z8iNyLlFMyVTi0B
OHuJiOXktkX7/Oz37bLQ68iFoo8xn56df6dXP/9WWx9Dlwb0rpSpB5p5jCrefpxD
eVcdcVV7Di8LOi+vM3jzRvhXoc4d4H20CwP5rbryBEm5piWqeSdH4i89v22e/0rF
vZhKDEJdxowenrUZ3i7BDcWwEzvAngz9IS+Lx1SHgpyvTrlsIH8UBkBpHdHBiSMh
l8dc2zlbXM4nFa7V8E1F8eqz+As7qzXDkEGUa6XDn0T3/mO1suPVr8Cf+bVM5qKA
+q9zZLYy8zpgfzmK8zg6zRplR+9BxHB6De/FB8D4IibHRy1sxwRsfbvLuvE/CtSB
b0Y3zQBY5jGWayyc0iFfuW9Yb3faLf+cFpuCY151yy5eMBs5YPoJCPlnU2NNLjIO
8qXP2lnu2k7pra6suRnJxvDANay64Ltuk/iyHDkPwDaQhYt+2+SXlJ+3AmvkG8yH
wiqG2ZNkieo4tT/46campGOQum5KUxjCYOxa4e8U7FMflj7J42C63MhjSXYJHMig
X7rAq2NFCpNJLGxQtfczXBmInFSdvQTWAl52zc7+PYWnBGst0Zau5IOjQzm2xv9K
vkvYMnn8vXFf1ZAZfINM17nWRG3VZ+rb3oDQQxnwCSh9Xr2+la6vHcDuyfya0+IU
eupyqJYcjZRPU1VX525zFTjVBbEV66lS8JrDyRqLyWf8WCKuOhWSo0FWUF7TDJxm
APShXTUnbuJ0LMkl/MLRfAYysc//Mbp57+4aTPu9PxoyB7eqCFPQZKwJbtS2kQtO
deLieRLDIJDq6jNp/gi90asC5A1+YIaCR7aoA8/b08Dq9YtuzcXnjdkCssDvBodd
VPfNV5TLpXRke2wAy+TNREFUCws3bBzoyJ57Ca2O7j1J9dx0oHCyYlNrxezwJtwa
EVvsZYzZfejk+fxAwj+M/aN39ADqtDV8KtzIvdXDxKD48UWFR2y0Zw0lRQzsnAYt
lN4KvhxGfnW8xv0xXdbqzDR1pv3ONcCuVb8Ls3NKJgRtyGf3uOja6HXzZ4OcQ+jx
ErGTf6kpfBRp8TwY9b4r1iyR2OQJgvBQKqJLM6QD2bLnyyJASoQh5HHv92xgxcAu
D2gBdIqu9lTJU1HHPBxsuVdUAtgaIgEFVG7qYN5wEs1QwZpintH31DUKNBch1kMM
BeuryEP1sbW1optN/aS4s2msrgTO+3wOLT0mDvNKQJpr0me8+XvmUO4eS3rTNDc5
+ar0+qmQTkt9EVp7HuXWQxUVZDf6bGBQ1jC3/SFCIOX5C1ujI9ur8xJt5uXSo+CO
Mosv1wMMMZLpOGTWExtSdar1uDTwR19/1BUSI8bL9hhgaqn5Dck0ZUTbU5Y/WJsU
5WABliGGcYhM3WVagoyPV7o9+r0JI823om9/UDCkQ+aatRtabv8G/9FEqW5rFGkb
K6lIB4tbb9g7LcYg4rA8wE8hvhmat9NJc9dTZByqiPgJ6f+++xesZwbGartTHgCl
D7k429BBS1Qv/ujBMFbVcH8p7kbYIrYQ3BaMyumnz/uZrb2DQFZDi0tcuh7cEdNz
CoWHhK3tC1BK526j4/Zgf8rCmtt42Od+dvI6fsFhPmxzVvAmh4HSfeXMjA+o6QuF
wSCtc1LThhLjq7qfih4asW/P/w1/C0gjc7Dw2sxkYiFPh/TPTcgx6EIVJv1eiDXM
LRwk7Mu3Bx4r7H0I3cnBrCSQ9DISUwbXQQnjigK0f87omdgxAjKAsxfQOkKj+8xL
RS3+vpaO0SlBk3Xa1T7jW5h5/kIMXeAo3aABlkP8pIjKxjqhA5MV5bWGfPLqHd7u
bvqWT0ferqkbOtgZvd2nRmMHWW2VjI5rx5uDlwsMei9um0H8pRzJOTgCiYAb3BIZ
dSGCxA0zvxVFTLjWphWbR09b64Iv9ngcut3OuF7FmhddoOsqJViCcA6JvwphLgJ5
skiU960MCX9xwcb16ZFhR18OL1FeFkodRe3E38n+L+dEe5rNqruiCA5K95e0oNLL
E3NmngwLwqsfSTbKp0+yqWjFSJO3VLV4PyU+qM5Xm695gyoYNrtpfDKlD++iuNmC
te9UWUzUM2nLFpI/crAIFHhQ/NekQtlPNkdrTLD46zwdR4RFllmR9nq7uA4SBmY7
qf9iAWlq7d5+vob2RBo5qvcMfEOIKY9y8k8rFqU1BnzmdYJM5Ly9rQzXBD2gkXAS
HnK1uWS+RYXZJN+FhHi5t/UoVO/VihW1Xfk/XCCFPODv3xTyI1jln3WWUrY9z1aG
/tX17SiYJy6cxb0Mmi9oYJpAcmRIJ63kStVoUwzWVoENAbSScv+CbAjAAjBY+ST+
DPDSyoDxpJDrKaEiYh6zmj3BVx/TtXtyTh8mYKPerkRNs9v/hBEUUV8fSTSIaG90
EkGwij2oJYNmzV4cUJ9s5E66Pa6bxvjCLSlx4fmt4HD7odQdvNE8V+Aj9fk/g6Nx
b70cMgWsaLYzxAXfu6obcLRWyk13k5ssz8TqwhI/fObzKVOWHDK3lyGN5GiaGQcX
LZZhZ+VoZipDrR476oR6lb/c3HhFrMShcBgbYRh6a3u4PDel8TjOXLhG90uMPZqy
bh/GDUnugcQKKa4PCscIw+QuVulXFUjTMfRu/2TwupWmuMJhEvTKZoH+H0K/PSif
B/9jv0htDFBPTAq1Cr6Iws5+q//8WU/2c7t/dx9Vh/qvm+ZS4b3CIBrH/aPaO/kk
AudGqPVBpNFirHDH0Ci93Mevt5jWJ1fVZ5sHBMECRqGTapMmnes3NmxdhPyTHrga
VTzLUPtRChCrHbVeQdTSx4YNdLct9BodOmOMhiUfiG3/eMmueYmS3WzH5mR1LELS
NerzeaXlxvY5yqMAONmiV3WzOyUKnWkgnV7L3QYLn8FRYWrMo4z+rzB5KurjLgI5
kfD5hJ4jVRRXseJXYRHVvLeu6oB8JoVwySn5ZMdWRo5psm1W08IlVb2E4nxs3+hP
EvKZEPLHdxtp2BzVu/5GqkQsaUO0H0mshsy2egCY1Pkk7iaNyzvZWjvd/O9aK5Ak
80drkOuCm/pdE2t32/z6OIFg/8M5C+4E4tQZK6+qjOjfgOe2dHsMGjqUOLa41fSA
sp5xOBaXONeXRPGOA7oQwMXeZTPLc59jWimOtbExOTpihIkJG9AYhm+B6fKdGJ3X
TCeiKrecVvha2mCtmO5zAvbUnSA2PLigWLn823OjTXvXiEnKQL5/ff2+DdWwjv5U
xAJpj6PgyeVzxyUAXvhAMSjaqAKuQ0ll1++IxhNhUSdbsbcYULExxrFbkGquOe8/
6lN6zHpAJ+AjtTdomVYyThmADUZkfd+H5/i9lKpuXw2EfrixlRbRGgSm6gTlILMV
+YjYGZRjVj8DTdY7MIoHd9X2OPAFAT6FVY16O4oc1uXCgsD8xqJWOP5jsShxRxWM
P7z9u/0DcM46bO3fzCMLO6QGEE96TxID6+K5IvWomjoBkib6YC9UatKPef5ghhCO
AP6ZejqeexoQUB+FVWsc4Lt16ed4rpsC19xhmoIRGxepqq0ISws/BTZ/3IvkkKQ7
4R4w6xYWJhKJo+X672Y6UWEOxyPIo025LDeD7J5WME55T/XNelkEKiy/Rkudw/c3
wiY1ELn0EO45+9agii4NeSJKn2hUGBpDgwxNHaw9SixhWoT30l++tQSGl0YBNDcz
m/HXa7eO5AFv9/j1NAprh1P+v/MeoBGj2Y4SaYOHA53piacGWz7HBZdkgZ0UEiMn
UnyvlVZ/BpknOuHY2oXtTapEiCElJMEuF9oGWhh/Pfczt7FZ4Tbazs1cy0RySKzf
aRIGfvGXIRa5TV4HSS33El5nfCDGe2/6xaxoQ1CwvV3Lum7E7AefpFzSaFUTi2Zd
yk/onbcaELs+JWg6UX5k+4YqyIGnaTb0CdFLvZImr+uP4LGWbh+8YVla1USh8Us6
z18niHObxBgEXZ4VM/CAI2RTEQ4TOUpDxWW1hhbCZPALvBrfhvV5LBDhLZV3I2Hk
CcORTU5Pg7/EsI64AS52CDowklzVOSzs7EbQPJUmPiTtYpOqpqP4U9fFY0erHBC0
TRLOAC2eyFyqxZdrb+OyOsG0LFKMpz1hm0pXxt9uWiSrMQFxdttIZOYCisYZ439U
AQ79WKEJTXfbxPHxI+Tn+eM2JRKDnOv+LViv/QhjnWgtJ6Rsm9H/vdfH7Ugw/mlT
GI981sENyueCju4xucVpCw/4LWUkwz5mCaC6Lv8htn72Fo/X4ZVXW4oTP1Rmf86F
6MB9+SkkiIHqHLoiZBfoMfanj1p9fiJOSeCaVI+R00IPgluri3rs/UcKj82XTIJY
7CxGFpX6ye3aKfgsjFn9TWYmc1zvZP2sbeN6hO9rXUWlSX4krqc8rYm8f5nj+gyZ
n5GG+MR0v6N/HTR4LqW5TIi0EQRR55L5ZU8DszD4Fwnk0g1VquDmGiWq6khD9pO0
7jfcFmxvVIgNlttrqKWIsceT+ifVx1HTKupwzxerXNtKV1vpQUedmye+bJj/1AC1
FVW0u2U/cdnGLKeLbGQNhtIv1q1fqvyoDDxeurVCZf/HeQOBC5M88/NwAoD4QAxa
xbr/at/65IEI3NzZFN4EVzrriUF2fkVRdRElUPhYGuwzgRSl1VxrrKn/Sv2WC+31
WSmiQTJWkjXUULr3075hLCFvI+qDcxVdv5+gEksl/CBSoU43s+WNj0u8M2dmIHcv
e5/ykLLHrK0EoA9nwXEWLWRy0nJtnpnTtAPUf2ZDP3ecLE3wn2TbiLV24w+e3n/K
KyderQE9ixRS60K3f3YYsR+xYZ8fyX9eQQF7+ePfN0bdnB1K39swCcBnoXv6FO8n
6k4TuCnrm5JvtTmhPwuVduC77PhZNg8WKDdQfB81ef6YFs43hioHgTul3f4gaOIa
Qo9swd4CkTAQ1sDGl6YNJR+7DxdMCkdvvOuTeit0nQ7xBxTBxRLKSEMO2Pli7hl3
k2voW1964J22fxjpl+nnabaULZnM86RdsMhS10JORob+45xkXZh8vvipvpkCMIO6
DbQoDq1b1MTwBMRQ4yi8vSvdG1YbEmF83txy1n5BGSIcjcG+YIssPZUbefezqWAG
eBoBJg/2Ad7Pszd4tgKCPpRu0nB7VM6eiffx2+tVJEaxpwLZ0sExBk7hk1tI42ou
kaOdAW9Q3vu92KWt7cyWdGPeH/n9YZs6yWrYY124wZh0SaVJvkiGBH7st8SjUVa6
+0Ts9nvM3c9eIUuOrwfsOYdO3hn+zcCvgP2pPms5Zz9EnuC7RaTTq0m+RnINnq/5
pPdJB3cq6yABIvScMO40USW9hqP3/xZf+JzfQz18mKmpRJ154/KMW6IIs6okswrd
cO1TICIsa+WStPwsmKG20LdbqH1l1ClfwLzXUIyzJoNdx5rXrI2f4wyVJqWwIAI/
POtrRChU0VZ640e5T36NoSLExOqI1jZEbgjMUl23odIGL1MpRX1fCnxkTA4jLuVg
9s9cKZu1dIMzfxt+4UaLSH/qF5qQMwaZHq2+mOVkxhk2QDzlxfuZvU6ur/lO3mJP
rJxsK2YBiPyFIawE6FB0xnIHr1aKm7VIu+K1O6CpXFFL8ECjzk2TMaK55l4vul1I
3l4eMgA5j2iDK0CHf+GDv0eBBm91whhW0Zz63h6MOYSznrlzJKd1ZCsYHeDEXJ52
GuZTCnmrGvq5HUS0JTUdKKdexQYWOH2CkT9zki/7tdz90yfFSZhyu81ZsUGrb5I2
ewD9X4DhQtnZyj1e907UBWHMhbnnLEiANAQI9ZhZLRG0AEX08p5l4nX5mwlFMXWy
Bh/WkuflHvl71cei9ju4jw+heLPUFvUcfVM9kwkIlj3/kDWKc1sRmmq5SlGb2SvN
MSwcpykAAOkmmtz9Lp/AiZV5YHVcZRlNRFIuhUFrSUaXpKtIhccqhL5pidUeWI6b
mT+ukSthDxK/Egor0qik1ABzaAdpPIQso7PRzZe1qPO0QsDpH3bxn83Xa8802kYQ
diGfNFZelyQE5P6pSJVOnj3z62x5+VWG4Bya5dHd8zZcY5Q+1nML4BFIIXn0n1vG
4ru2YJ47lZnLVAH23ZUw2uMgwC+wDjrV1kF/nzaO9aPpi+tcqh6ddltWH9d/twOn
fFSVpj/ckVrxYwzf18w0gEADrHBU54/II0HWwxvAviq4OJKhBA91hpvqNGPM6cZh
V5mADEfY44FrnsyxH8/NXZjcaQjHrS+Of8pwzfDVUEEzNc6bJYP0DZWNTkTdCIDl
iX528th81WV6NBzKG/gsuylmF7k6PC5H4kIYfBsV05HgrO/heQBLcSjJzTqS37Vd
AEoo1w7iwQKg/UWfeDHOXn6XkVftv8Z0WUE+rBtIEXgSZwaRQc+7MD+r2upRtrVa
WvrC9F3n1B+YohRPnmFiHrEM5Qe3uX0vWHSmCUJcZZXR8eU2eUNDUptfH/+8XaDo
xeO2uAykQkABJgCv3cdvYV41eAKnFAOGqUpFqWkDEkVi1MBM/7U11yqVKAwv4NC6
ZVly6GJ+HG0GcDv7phhmLm2TrMeC+u0Nu6jJ9+ptoS/s9ALEzslB8wV4lodCz8am
bG2/L42fKXkQNuB9gYdk629lp0E98FEDQNrkM0IglxS7EPlZSCq9cX4jlq7SMsah
Cn0pgb/EHQR3Er6RBQK/uyWz8eFEog/E4adMnuPdlrr4z/mNdnOnXYWirerkw67/
1rf6Js/jmddquYAjThct78Wt/2h3AJMpSotB40rYuTqMO6wlAM4/RyjnS6BRgCoo
B3dOdb45k+b8kjUObSdmm5Gg1d8uLXvJk7dVGN2sp6xvl9nXgHBSKgYQVhfdDRs7
KUkQ4+UUIv4nPsIMAnf0KrK3RM1jcxWeCQNMzpomwM7gDzytkJupxxz0VpGS2Hfr
4vmR+5zj4H7p76c7nh0W2ZsXjVfkHRUKmI1f0Vxe8O33oY82uJa8JrsmvAfgarta
vBw9fLpuAMo+tYUyLe8mR1nb1/nQoBS9xxFz5CKYYKVys/2B9as2ze6FPTJ+zrGP
3nPk6/KZgfRxThDtvCq62VIPeZwuATVcEywAsmYXShB6e2YA86Nx6vyssQd2Fjos
njZ96Vd9mZWnhelUReFOm/LQAZhWMAbcgO4HAyi7pG6GmL57CGNjq7JXam7aTBS4
yLnZSEZWWBYRD/Cvkbl+NPZvuTucALobiu/B5q7BMTTnol4a0cBtWyDRr/noZLGn
KiQS+ZMXz9sVDIirVmg5YUwAJzb4wfhtOd4so4wzPlEYvqJXkxIsEdoebZ8q4JWl
ScL3zVsq5i+DfQfMg5O9BhJ1gh/AnUsJevN1P+devw6+4JcojSsyDRVZlAae4scj
oSV+W1YAFo5Z+f+TkcgGeyVNJXvkx0Co4DL/4zLRWieCkR1dXE7FKbQSNBVZfTdk
08Q63qocQ2gzc1CelkpoZepkjhlVlFSBvG9wCq1EL5n+dI7HmZbTG8b0Ddr+uwDn
CNLaRrYoKK3HGZGBT1Cq2rZMfxdMRUppTf5Ori+Epjg5woUgoffwDOFT0XlIg7ZD
jh9nqNmBwb17OsHbbxe8fcDmAM7tO0cehaQU3q0SLdeGlERf6NrrE0OxrXWGeLXE
otcgXfkRG/8H86lyr/41n5ST/XVyqS2INg7W8+ADZkZAr6kh9h12HkzoYbm5vj2H
AVrQiX/Yty0gNTw8lTBNIr3ZsNlA1vj8icHPvkIeo1xIvWs5ipGIYL7gxl8WPEH3
m0E1ixq0e0MVI35VL7X2OfHBoxXrOK/XlYpqKo31c/GYKlV0yXXPPMmHMNDStXio
1u+QTWXlfSTWIpqRg6gz6FPtFrR6UNWYaiRIyKshUv1LbjivmMg9/wCL07pcSpr4
2ie5VDn9/Ff90BWhstbHqk2pzgEGS+ZxzVtE8lM4yqnKUI3KXCNWYCZtrJzmJ4mZ
h4+ei7BtsGQKgwtJnDqV7btT1JyobiA9ovoy3yE+ALUVvL7KX6bmNE1PYMRjrkNz
/M9zMhecuPZhNJhnRCkAJaRpKRQFL5SXYXAEYgrMFxMa3wUooZ9vBmBCKOojjzvT
xfAWpD8/CVVB9VNq/YwMuTs/nojUk9GMebAgigLs7aHDKseovjYQKI6C7Oa3rEMu
O2aOKy9L9HcsQXFbcas+c9B8I6Jrk0qXFAUprH/xHT8iDfadfZqtSrIqiDvFpHci
d00gtXWiMvsf14bZH1vNnnVODcqcfLEwKc2jYDrveP6unQpN7YVKUoD604nAuq4n
MbbngrQyphJNK5lBs2c+5+zvYqUAvVI8TBIkFMhEe9RWbiv2dqurRiBfSwInsSsv
NgwxAoJGssTzR7aqap+URjE7HU3upOCYmtx248Be/q+oN5Wioviu8HwMUjTOCXO9
YZooR9t0KWCiE0QpdnUCPeBl/zKBKeMlkNJyXi9bNT+P5LlT+QW5dDP/6WrySEgn
x8WRW6i6gDDMCN+BxgmBw5N3YNNEWfaZIbnqLvSbv+z5IaVjprxklj8LcQ+YcTI6
rgbOa283CAEg0KScbwJ5mAsLEjU6l1gGLFOEMBJFYKxlPdr01W7g10ma+rezK55c
OFn45gu2yDk1m25R0F+t8cpMLVz06MI1vftisOCeTL3FJlxOAK6I5322SGszX2vm
9yV97w0y8ljlReuFv9Z730ZjnJ5vZe6jfE8ZCFtbCsPkKxjBWYI+4wT8mD5IbssF
W6xLpSOr9ELVrE8Bbf8hxBCTD5rwkisJcmVSvOeDZHwV7Hz076vzzRh0xjtIADAh
KwdaZjSf7yFL5Z4634EowKEpH0vOxA2bYBWgXiC0rmCBMKfRFhp9DxgL0olEj398
2s8akueg+60RPLWT3Kdwhprc4NnK70Ea2/QTX81GeSZ3NFCWRYvNGwY88o9T0u0l
zNUTP677c78SPriHkP8hVNu8xOz3zCjp1NzDak8d+3OqR8VtWXTh6SUzIeOmIAqt
AXMAMs8ZZCSGO0ouXo99kKKwEWhi2QNXAhOt7P3m/n3eHHZkEM98/4kstj2YTSWZ
Lrbc1xOtOeKrclIrhba/i41ZXi0xt6VBdfPL+y/pXxpmCbcWlVlJB8y8iKEhrnVM
q7eqf7xSL/hPDwNcULapXX0LYzsn33hotFnlJXmPxgVwTmSfToyWK5i8apPN9b3s
03Vz/IKvZAbcxVlIx/aUYR+puvL+KFXNhE2JHNfwqnALAYjMnQQUXjnhhljfJ5HX
c7UqijJe2snAo/znGDQ0Uf/fBYrpO1N1FsHNNwTFNQYVpOxT7huGnLt28VhUiyvn
79in/OL2ghKDhI6NGDephcz/Y47TjOYMSSoFqnOPlZkAAmPhONy0zo09dndFI2uT
5Lw4aLfEYB01/IIlCUd1CxG3GkZTN7hTImUyxoSVvvainQRdFG2e9gP5pa/N1bmk
U0XaPAK4Ez6pb3husmldDEXUiwBqKpiadBwlVqqFomLoqlNix9OFOSGurx54lQPQ
n622KHqQLWw2nat59b5M6CbZkR3IEePOc2jn8FK61BevgvOPPZPoEeILAXXjIZWB
SEXj+/93195Ax7G9uo+Q8h3/GJxaHxSq6pPxM8E5NiLSKIt3dKB7MoGyeqflirDw
R7d9AQyYIRHUa6CrZVmuNYlC+MZBoxe5zkDGEsieGvyHbEUBgLHToBVA7yh2Kf97
ifKT6lLTOWWbP8qFd5uWp/sqzhCkPYTdYsPRmAI7HcM/WMnpW4tJNDrGC7MIiHYA
zFFcoz8SKQiXeuwFdTHfCyTa/PFBxuyc5hKxVrZ94LCNtM69JJDxNYnINk5dCC1K
GFemheObprem8KiLoyL5TRo62WZBaePbMZRe8MKlSEBwTf+/gS91rehhlyYGKsRd
Wu0Yv8AAdKc2OM2uGEddUQm3zMEJpctKxsAyYnxx2TQmgsk0C58cgbNi8gwSYOL2
K4eDbfUZvbc8AVvPv5kuJdWCkD/Pptlb4TIFJop1NnNzjKGRRF4/Oxzkgz64kEFH
gkiOHNnvlVIRdkhxl8QPOr6RSstiXyJIDGLKbJQZPFyRbnNLjbSdjTIGE84xgoXs
iflQmkjxeilDLqWw87pqz4qrDOINn1ryhaW6R4FN8JrQJ8Eb1I+UOcE/D54pQC93
c+EA7bue8Rdk+7wB8ieW4sfTuXoBI+tKgv2mwiCpFtBhBrI+YqHfH5P+qV6owZ2K
3HOnH57H4K4BVAWjJmyncLVPhpCNj/LuoZHmLx2KxwyUpZ3lQj/z7ddNu5omsTp6
mjNowiYrm/WoZC+Z+ycO5hoKuN2ss0ijj5RTr2zfTMTmsl/2TAxlh2NMvbSSGb9n
QJkch69NsSwB8yiCdDVi0+i1N/L4LBv/BrcW4YqvUgA9soDl7lbBQLVJcRuVSuMV
fQhmwEPjQRkUyHUe5kNpxKiOrfsorRbW5OBeP/aJH+OGtXZ6X/bfwgdCMjPMOg2/
wCqWR0aVyW2z+CiRmioSBUmN8EZOiXjG0SonDIkhCj9Gj9pwXvWpMnzCD5jgeaKz
t8LBtf40zcHFID3FTaotfIotpluO77GE3zrXdGpkgg+mJ5US1Fqjhk66y5QKeaYn
SW+WZg88vjp2DHS2Kz3eaVredu9YXrcjZ/c6ICd9THUTBcyv7H0/h4mLnPgPmcoe
eDCBB/2Hrgi+go8qb2epFFWaJUvfm5WbwiaiQLZgIGTgmX/eVGB+7eVria9xCPzA
p5Z62s36mHg9W2coh/jzKqi9bYCWtU4H0IWl6MhwiiWFY9roogKgVj+n9jqdnPOD
pPH/vp7LyyVaDtGiMLmSIjxDQAS7fHmfBioWOJFrvNdYAiMctXMnHX8QhV+WHPZk
7OyLHUQZoFxd5S3skYa8TAbUx3X9k86/AzFqlgfdmYPCN9VFtJOXFlFZSFXF6yoc
bN1EhVqmRK9trshnY060HrnwuIV8+1ejMpuZ/emqTzgC+H7nwJMG3S3QyC8q1FMU
iFGdn4zPU6K1SoZNcs6ucgAZHOo3PcRAMC8KeVzE1lCtbQh/gwdKSQAPAVS9766t
dmmulqi//TwxRRuM0ub4XuRMcMWyWX0/ib7ynx6WzMIHazo4iV5NSC3wkvVUoiSl
h5+zXFeY01PSgSJnyA506qjvQRTPVqGdwG7+Z5B7TpxdJ7t4Uwf12uEcGbrN5Oib
bsxChqszlyTTVNWca7UrUBoyYhB+0M+whR6gNSLmjyCSHHuML/ChyLilFgEqGrfW
cgg2uLFJ5kICFq4Iks7V48nVyZUzsvVUo+ljuDd4FRK12anOALk6FsrF+XxID9kh
O0ibVBZKKKiwF02VdGLKMWK7Ka8L2qMtqtsfdPDpTkqzLdN8+SCkPHsEwUi0rUI/
wHqOC+m583DA2I3sgH+dd+wi+/6L/ud4wwA21Qd0pR6CKQIaJDYtQY5S/dGdYE7i
dj34KaU2Ak5+H41z234X1v5agaZW1u6qbLMqufB0aYCcCnQ6nbPbBcQkKOWstA+n
hRDQxL/0Bt6lx7qVxwllW+w02QNXDnPz/Ec8FApoF5rVDKsjBvr9ndI32JE/Kttf
d/nMCaszH90wtpspmlX7BeiLeB1B7bzn1TSswrNXCzlgRbtMf8zG/3K8fZ0Lie0K
lG9CrLsV3Ouu+ooNOAR05Dm2gKZG2NemtKTMAV+MxmrjjObu4K+asN1f9RypIhtx
Fxkz9YSUZ7ULTV3d+E1wpMYOZzt6BFxwtbuAbSTPfVlAGmrRrSY1g6JvvG0UE8al
cGd8yq2tIy+qA4J7s2qKUZUQ2tyfGhqCGpYZExhpxJXCrAUQ7rORUj7POsVsy+im
V0l8QCsN5hJHZ6e6G60N8m/zXvGl0f+IwuTsIFWLlouV/x5x7LuKUwNdSn98J9nG
iGtE+gOtYgaYDR0jonZUJu0bx6AqS3HcHXkrw1pqyDLP+YgtUTS2a9ZjamFpHCfU
Y4bAdx5jRq8kwVuZrrTzIiLf8fLUgY0rcxR35IoU1faxJ7c0BGWWeNodyFUz8T65
vEy55xEJfLwA8jyx9JJlHm9PTc9lsgVbePXIm9iEUdIe0R17v7kwUu1bVGGytqM7
8aDR9jzJZpDPj6RfugRjHsmDP+DmNkzv6MmSc7t1kSmz8OxDPHZ4e829P4hGRwTx
VBJc2JD28gRSx/yqWCedaKSxRWrsjqY64SVXGTwnerEmKMvcNRRAL5SmvQKQ8Z87
QlOro/fls35yE5TGvhHluaiuYGw9xjXJHAwgg7qL8ETW19q+ek5q9iLjj1/jvr0g
5M5OCTktkY1FPAxsEIKyx/7I5vEdt3bUNIn0LyzFr4rwa1+lhzW4fSd0boN1mJs5
fQ7QXGlvHV0c2wS+iF8n8nz5T8gLt9neqRSjP9RKjEvVAaNRbIGG2vGtxiByzkNV
hjcx98ovMEcn3YnXgOHhitzMiSl0HL23AxKUYXPbe23H8hI0ttNdFHC4sQP7VjyJ
mMh6hu/XtBamgbyYiRo4Xpjrd4mp60QfFL0OkIeuwx8R2/SAiOzqj/cnJafyoYtF
5b0Tjg5m6CqvB2omSM7u9ITBS7ZAFfsQ/y5Lf7dNaSpCAqzmdDfC1NKMfD5J3BcM
eqyPCyCse/DQoRfYsJfc0t//dqvD57DiJHtXchWxKzn6VWxd6DxLwCLrW9+UX781
jgiOZa6JqxdUmnFsFgNcpFqRLd295FlRvlfIphPodrGdf0kjwPC/av7VIzCFZgp0
4roMXbBvmQBk0gFn36LjIN7blUiigW0h0X1IW4WQE0BdE1pJPSVMRnGzYgnw/21U
ylCHHHsH5wc0QX1NIowF0peR4vnBbsPr13Oa6qVSN5hh1767Q9zN1rev9Mcdg890
yleYqilBo1SAG2EPzI/SvYR7fbrQTuBleg88IrYQ8fdQGz6ZYZmf7QPy2ft7/vVp
/zvUnm/GhEevYqGTL4hoZ/jBaGtuA4I34LkQjAP1mODdQiRJmXzD1VWSC1nDQXkV
OxA+5tp3TBBCoeONJxtRZBC5wKrkpmGmy46mT8MRR5DM/1NEEGuqleF2cjqf789I
dqhaE/5K6TvSjQIAjkYK4lFBf6zRo4rOo/pvaLwgrteUA6gHAdWWbCmr9N/F9zf0
hEi23e1ZLNLEj2p0G+4Lwo4X0z04/t/1wzA3XI2W9R9T+syvoLd8BLBUOeX33j9o
oSxd/hqWOAZhYP3WsNlE7O/0l85c0QRuxgov43ilX+MbS74t2VRziFwxMdKgujIw
XRNejqlwPZbKSsgjDqDdAsuEZ7JGIGAUS2icWh7LgglMleMuVm5F74SKRZXV34ma
scVfw0Xpa/TCYNPCvjbYwSnW4Huum8gejE54b5jQTk8Ery2PFsoHtU5fQCAQzON6
kILC8f2RoenIqv+DiGYIAZ1EkmsdlVJAe6wL9IICIGwQm3by3FqKh+TLwwd2T0zC
BJsVOYVukAHoF2btzk9HTm75XM/VhXoIGABRIyw1jLy8kBGaRAWZph9CBbLCi+IF
Ev9uvZazk1H23AcCmqB0C7uwqNL+F3lKSkaEdtNjMEl5RXobnB7zGxFsi9MKBTy/
UeKaVSks61eFks5mQneon74XNeDPKFxjeqlcykDo3aLD0AXj4okfuhrCynXzoyWZ
NsdOl3d4NyxZIgli8PbV4HKqZzeGAb1rimzDqJUOu9JuoVY95I5CMpp8JUp/fJcb
+8e19TIPPYu0s2VEkW0Tt4mrRmCxupiLZuhoJjf/OMGFU8dqgIxHS25B6EDDY1Mr
ZqEla3ppXHb7/2qZkxe8Oi2LFEyqd0Z9Eu7vhomRF2Q=
`protect END_PROTECTED
