`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PObOVs7xrVQR6lW2oHvU7H53CQbKM9NjGNJj8Gb2BZ0zUJys/uh3rImXlR33bP1k
baoD7txZFUrbenvOer/FXS1PV/ERLsR7kT7WfUY37ymLwlpaKEFfqOjm/RmM90pk
hy8c8sUzvq0OKT9HvJj6JpY+Nnsw35Qnh162CcJ+ToY4XU+mj6MzslwVP9TTYDNB
GxEAodRJNakdG7PGjpZ6LWL6K6dex0USj3RpwwwUoMND7P9mV/9u7xVQt2vsSar2
Kz/rbjJJV+6jPh1gWfcVls7w+IUWOTPD7eEDrL4hORWjGACbL78i+JteFXoRzaUu
0UsRpu8JQBWOIDkl/kz2HEdLfxUuJhpeBavRTk9yCql4koQo9DNRmQ8xJ94b4KCV
P7niF4WacKEKxJFohUjiZOqXdiAU2OweZCfbcloWBnV450P/ug5eyIPySfT5+/S5
5SrsDJT4EGkpYIvvXIq+0cdwGrc1Evoj1hssV5rijdegVhGMc+HNhLF2Pdp5SZyq
AOGOdSkMs+JMIt5IFdbo3AT0xI0IInvNKbvzRn6FE/dIdFKaKlrJEYm2JmIKPLjz
r9c8qWnfA+VBpxe+GLxi1EWO4hIqXTFDWuYtPzh0bZiPVNEzK+/hY7jV+Dwap6RB
23UXF4hRMyyFQ/PCk60liVKsyT1u/iJLBQxSracS4BLg2iaU+CfCP2FpmPorbvop
fkwhpkduRtH8KkyPDqSJ/1LoEAnXB42eraAOXJjlw9Y=
`protect END_PROTECTED
