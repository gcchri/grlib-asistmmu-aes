`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5GeiqIKTFR+CdRbCqeRPuGbByuDZYREblnTmoUaDu0LN/zNN2zn9UYqlfEJ1ZpcI
Zj/Zm6Op3XX7WB4rebgzQWawsAQL6s7zkyphuvF2+r1KC7I86KQelRljPxKb+ama
KcJ4ZxEP+kde3DmQ+dBd3mLpJJ++9zRDqg/J7bTMooKcdnoaZQfFc4ulcfYNSerD
9rloceE42dK+SoYHSe9WpUyanBEvL7ZLIu2lFixPtb60Lsp2B4vZpl86JUnrUpc5
kBD7Dahx5GXT62NHrgR60q9ruz7N5HFooUZPHXa/CVp204yVINYRFI+/gtSQ5605
khY3TSLKLPvyw71uSa87Lje0vofHWz+CWQzKFd0UtIt/im8mdRYI9U8x220H+//F
QKVmkLOrc/82yDtKogLch3thO17BrmQ6p8mdZWSfukgYa8bYpShA0Q0Ydmicl//5
FlzP6VmyWn+GqGvA0a6Q5Q==
`protect END_PROTECTED
