`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q7Sd1W/hx2q+0P5Ukf32G4jeJAon3S0JKwQYqjNcRXXYQ1tjlO7h9eSuzuzs9YNk
09rU2Z850VpzHjA/6sxURs8Hh83710j2iE3yxVW8PdeDgfTzHirbVGTjYONTkbxw
urqX7Mqu1FaeZ66+6CXOmglmgQNyPW9g37g45Zp3C8DU8ElmZWR22jNBHwbjZgUr
HVvNFTw+YeXedxEVI+8J/1l/OqYYXIXHv9uldswz9pWjK+h5deT+CuwLaG0B6s/f
B73uLPVyI/hygb+ltyfLDE5AYRdk+9unj+jqvb2xZGY=
`protect END_PROTECTED
