`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hWGHTux8wgnsFvtutoxr5L+SxEaRuMGNINrhZUqBqOflg5RaMzxDIsOe/WhQgbIR
yBobtWDvdpn9qUQDAX69/hVchmLe8ROHz/HJjxUjky8BWuzczg6zOo1LVZB2W99l
tLRItRjdEeXQhfJ08wnuAyYc2LMN70eYUJCKmNoxozsalTSoXOAuiq0iBfUyOO6g
lyEcpmroF7BLTFnR8TTfyAvbCNC3Ffqin7sKCjGpuB5vGOGn7iAceQsZ4g9OQg2q
tSouJc27PrY4x0Yv6ac98YfvvY9VJRNQnBqR4jiiATcN55x63IlDL6yB5nRIiHR5
Qb4/zNMjsJ9SvcUEseRfBxwflokQ+iEFZX9/pNrkYYspLwKNS4j2vnwZeCx7FawU
6kwxm3Ets651+qVbk41zOjas8DCcnJuaAeqCP7dGoRL7zvTgQCFkFLb9qoqPPoYA
`protect END_PROTECTED
