`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3W+QqWaJ+iVatrcOXVnFDBO7cacSLNLq9YSCEzkx4JxcPKZDxP3i0fWtTFWbuIgB
W2qi+N4s2AekrEcJGfedam5hVUtldGeu8NvD+wHAXUcyLx0Hm3Wk7YusxlHpBIkL
LkzPopKIaw/WBqcidBBAYLAFHxqOgE0i0YEywUB+tOpRCX6NnHyCFiBEh9MSYwgo
VFlYmuPMkfY5FbiMx7APwQoNAjBL2QQ6QRv33SEJHsicAKS7Eg2PcViSCm7XzIk5
DtTxwfRTSiC3HE42Iz/2GdNd+WiLZXYi8w9nSROU/sDU6EeQJBJ61D2gbd01qSMh
Jwr1Fsc9kn4PLekTaFSJKyCsaH6Zbz5K1Uw7aTo2x+mCUcqLzmN+oU9dSuDeyPN9
p27fgTsnZm5F12lLuTs2lhAH8nx743AI+sFJMzr29+3guRnghwbgBZGOCcah+4R5
zrzssLcUVPOwNiqesGu4/2vWzR6CKDYFWpjHjvpXj07jP3clDVQk6zCTv4rSYIGf
FtZSv1AxelcDkNFJ9pwLPLsLuWtJkhiZ5aFzG9HPNsajBVSXob9EtYa8K5KzZb+Q
2I0g3U5JGsW04pHpmNILxKI3WJ9uio/fennbva7mG1tXjY8nWRI1jiUyMFkkhEHF
v83cjEll9MSfCLdwmeag0vtxdm0kJ9Yov+zhOw/7Gt73BjNhiSzfCEUMRX5bLWYW
plIYpIM0jiOBdYaa0bh0BE/R2BEHOnbQrH1/ZjxgfzU3Ta62osGJbPGjwI6zRu0j
4hbQNdbjW0VDRniAapH+WHina0mDZJu7/GNtH2fP4wqqZPItuBkfTh1azFm9voyu
lWcSWRhpfy16x82E9Xt6N47kszD9C1+v3V/oP5FlbVyVl6zU4t2jnAln5Mp6lIz2
WcmpbG1/0bsyctsyZStXj8EweJ3lKR++draOoaqtRtXU62T3ML8AYcfyJ05by07D
TTXRf7c+7AxLADBlWggdqs5q6GOjglVw92Iv3D0D7mgFMsYbT4cF5Rw5F1kZU30+
STaIUaPlST9UnnM4cgN04z49MzqBNw18ooUL98JUONYgj2gjUsR9U0QFO4epndtH
6JIiqYra4jHBgtIYH3JHS3rRd9QFB2OF1V94gp81XY4GyvAfcVLHglaB9NOp7lny
sQ9LkceXmV2Tyk9+1NVe6sAgmIGplQEY6hKlLGL2m3VYnmC6nRrr9QJmmw9djIjB
NcKC1KY/1a5GMo3l6Z5KQR2jCxRKmGfz4Lkdd8T/tAcbXIssHToUk/15j1BHU8VW
6vacIzprVX9s1ft7JT6iN8b0LVvpIA0Y8nU8kMYQby5333e6dZsFrUdqLCNv+HOg
lrN4d3Fyy7MdO/FezcMr0oPvVl6umWRWhrAtuHtY5Liy+LvpWW7qjSsDDbtwNKTC
mf1XLS6+P1Xqag67P1KHrmNiiXWDYjyNnli5RIb1ZOVSliRB9uBMhN8cfbFQDWWe
hGS61TSAmpPoQBZ3lTwxcvo1J3AWc+Hl+PCA0r2qhOk=
`protect END_PROTECTED
