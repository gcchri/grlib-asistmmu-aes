`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5s8Ttb67pxGnYK5tbofqMoSpBd8R43zAxLbRy3KaGef9NQVInUiqLhG6q0EOdgFk
gJcaW1yLfHZS5GYTKsMRa+tAbV7jI8KOHhyJpP52tkMprtTZ+1xsS3+LXGrzDNvA
wv17VzdIF7CkYvx4mvCswbKVuHhzuic9vZlFx0ZPsRNwRHMktf01EiVrwZ+gtWUW
iPbmNUHr7d5Mr1YAnEc/k6fmRYTP7Db11NRWhR7OAg47sUU/WWg3CRt6FodwPHA6
pxAaLT+LlnqKcgK1G2fsNIvsWGZTDmtDkcjc5PLuQXvdgsaZdqECuK5fb6Y16wJi
rRwSC3aPKLGDwINd3pTWdXQLIukv0hTCGENhXt4ef8zQtbrSuip9Qap4XLV9Xv25
sWXX4UWXyWsS/GT509NzwEODL4veEK4/FumWvdKMZuZ2Y6mVllid4MOLg5AbRsXa
BdXTlJoIxaiERIiGueHx/MO3pezTzXdCj049kqXvz6XtAhHTZcpYmHfSVhjoxRCu
jJA9VRNl/8iBToJ+1Rw8iSHcEsq7Pgv706Ru+Gv5sNeUy3bqhJB1tMC7Fa2/m52n
gM4tHwYUrSsB6dUpEFxmP5rOnMGgq/zzJ8zMMh8SAcC2QFEPGNR8ITwe4bsJAokb
vjY33TIYHIMG/GU4z9Ih2UAh3tlm6tIzUtNrU2pWtAs2ahVXE5aTB6gMG0/wVA2h
GsRwd8Gf7exfJamDuEnvE18GrzuPKoo7Od3gISDT95H8logaN/bdbfiYyKm4oKBH
WqQJpHOs926RfVCVEcDwNCh7G8nPiSymaxy+avKOBwrPls7eK3L2mGUXU2ElaeQB
vSfG3WXBqtU+P9FL/swJu1i8Wnws3bToteSMqZYEFgPlTf/IB7D7qWPtMtpnv4vD
DXLU6s6j7z08NdxkBIDZgoTktSM0OjV3IxZx1EmOJVW6x0z2MZqWyQ+e5ScGXRLf
BgVS4u/0gtHpO74+l4bpRsknL9dGKActac/WijpvYsFzsNjMmbDvA+M0sqdL9T1V
gEVi4uGe0O/lGP+pDUGIj6CtPrmkZCyhT+d5hAtxZHQOfYTpvlsGOOw1dw92zwbv
Pfh6RjoptphCBnv0eYGQBVckJAAdupowap963c+bPUIDa/SmzFElpXv1X095p84w
pfl8cuChNeIZjyBn65AtCXYknXZNYauZwzANbXHCJpn/nClsFJSDfZaY06psDlKt
NtQFkuuznXkZxkjfACGoFjQAEVtacBogDqbBehmUKwGrV7iNbiSdeUJuKIFg0cI1
V0kL9r6/Tctg+VDBzh0EFz6QBDOIRDtaxfNnF4cY0V/4HogJ0iPirybZ78Fpz6Z4
36b6sA9Gug+BWnej+pemYXl5gf6ciCAKfZpwSraknLX3al29M0vGNVG0Hz7CItlr
w2ou1g3J0H2+700ZtCSy2tcCXGhwG6X1kZEvKaLCbuVKv4h2lAuDzLlnfENZ2bcX
cSu0lWMpcU0YtjlRva/9ES0aRJRcrgoxEAchdzmISsP6oWASYv/BRvd+Ckuowj4x
1jlu9W9a/DHQNZcsPb8iJIj/LoRpbWxSx1ybGZsV3hW0t4wQYfA2lK+AK3JsQKPb
GRpPdTQaidMh3H+UzHNTt+e/mfYPnt74DTlFgLOk1ltH43SoIePFgnbrEmLhSNFT
aI+VB3yWaLQPHMMja+JXorcIANDHaJC4HVPt6QtrnjsNajh/skb95AWe7wmt3FSv
sTO+zE4rxQZu5FOscJg46slY8crkJhH7xHaL5FKW0UjEER1nrUafKhqBvEx6EVob
8noxXIG7nHuc/hzDmuKlfSE7Y+CNu6IRwOUjLEgXk7zN19Mh3ImGAy+zLqCbGxCZ
lw5eEPAHk8+aJUV+NA0RO8b1cR/6HBzdVwChRPtfryijY23in1xYoGmWUPWBX6oB
N8DNwRY7FJSlkmJ6xN4Hhf2IuV4C6K9TUcSPRYQcjNwY1vHY/3c5Jt5Sq1Mu3XTR
zR5j3HIEBGwS7hHj24cPy6/2BtUF1va+2pGRqhyJ9oN1YxITThE/L6vj3nzzDz98
pvmC4ZIdUHCH/NoBo7/eC/DoJQ14/snX15yVH5vPxZKWMSR0MsXy0slQqfGPXeB+
mVEL3qn3BiXLXdX0AqjqOHemQsv4Pp6l8xpdaqRvioTdY42yHFo08o+LYwWNgCiY
JC8oG5pqyv7gIfE8ti50CRX9bpw0Iw9kPPqbozqFsX3ABkDz9Z9OZqo5hMlCHKoC
cy9p7niGqqGLyhNrErVf752XJ/Z/uKo1+ht/eaG7D33D0fS16dKlkxad2nTp296R
+6S5FLfznsKLJg3r+wHtILiTU0/zYez82Zom4woJsoNnEHSLifIsE+rKNPbzDm48
zo6m5yYcEBMcurS15lubpT+zbswOzqpeTBj6xpYOvbABcc6J+4vSqB19Irl7HqSv
PjBcl6vVkK1ucEoVjQtoP7mZnW8ZaRRYxfBy/qv/mLsFbSdmAo8tMtKcqZH+8RRq
kMipN8t9KKXcdFVOqsW+kuPGhR4ukSFDWbqoVDaGBsXe5pcqXlI777+sZ+9ADb4n
5cxAx9h5hqYzcEzVr/IPX7pvWn8OegZOh9y1jZbt+prPKk0nvV4WS+jFQpRO5VbY
ILCGhtswugISrAlyUVAWMjK3E6inkmT5G4lCtocAAEhCW6Avwo7P9cygm8tgJXZv
cUxi/NIYe5G2xJg+K1U+ODkDbLfUpJSFkyFflDkwri4HL0544ID4VhePA9gd1jwH
mq/NN9ncyX1XLsr5SA7+oxYQ/telca6ngHo7TP/EljFlq+Adcb1vZsQJNy9JV+bg
snXjewUW5knHnGlYtDc5oh2+CDQ/Q8tIFLeeOed2jyVSVYOt551B0hV9QqfAN8jR
W4//nns+qi797AA6krAN/AFQNOy/lLoW+ou4+fKTToPA/IKgM++FckerzzP2MC8Q
+u+eLiif0WX2BXadPFKAXLI7fSgHWhSTgFTzH+gjcOm5vSu90NaFLvJK7ZCztAfs
DaNX0DU3EMz2LhSPaTVBT6RjenlzpbB3qMPwcsOVMeFHK2AIrncw0ZVRz7rB6dss
MoFXB2FQ7L845u482cfLMfbs5m+Z9O0m98UyLSKa6+dT7ppbKedFU48OMYay3VpW
wCWrOc9/sW1Mohi8V99yPWTyIozF0KzG1xkaahc5up9fVLKuppHx3uwVkVTleBwR
WB4roF/2+jPi0BTxS4w7jh9l2Euj+1Jvyb/OdSr6Wl7PZ8PvpuS+Ban+zA/V3JXj
hVbjpaWFCI4Zv7QsTXWecC3t7Sj2nQsPj9N0FhlvFbddfKzd23rwUnqGAMFrQQfM
o5jQDYBSXRlgeAAW2gPb30SlKzFx93nNcLkVn+Hm73x+BprCUUJYNnVz5TDFSpel
G2R5oEnvR1BCAZd/Mux22htFDbNkp4h/qxZc0x3PNGIrMwr3RSX/mZ7C2cdqu9iC
6HL2RXOyaC5X0CiAxNJjOGzDLHtHNQp/jx8pTqd1+ukFxtmnbzzVmT1dvTNf1L9/
i0b2jRfQpHiAvVNfSXWPf+AXbbp3RHI/vCuGuYpStoh9IW3aak60MHI4qXQoN68V
myNb3o4zEvrdUjBZZAF2C09MlGFYCep34NGIf2LZM6zO9cAaBqK334+oBS3G0OVq
/af16gX4SIs6EXZQ0OWmhNo+jzVhygmV7KJrfYRtxw4OSHf1k0HcRi2uen6qN6IX
cAyhQPS22o32BVgR5kBLzcJSpMiWKULlf41mKLPz18O49HyV/Y6G8OgfGKQr4kpr
tlrzYwKE9eGcISQ9D1yDmkv0XxRfEp85P9H0DTssdp5oMfKjFYFc13urF4JT7QTW
EA3Gfthxv7ThjQ2p8MPqkzNFRHQz6pJzASH8bvgHs+ZYnvtxY5ClcPsbDZuU/BIf
rDmDTcQ1lWH9Jk6IbkNV8NkvczWsLwEfx5brclL5CHzDZYVlPTbSy+YnpBxJlDjR
GtjTEt0Qf8Fj23KyYQyxIM6GOWQBG8HrrtqFmcNRRvail42JYVm+IbAYfG8mOgRm
Y6jqYB358qtdoWBsg2enT+Wtl0MX2NKIFAhRfx7RAM7/V2sw3dsHt0Acr8Wo5AnZ
ZyXdvUQ1pN8Z+I/o7QILEiTNrJ5OKzRh6Eo1cxc9U0ZADfOf/7Elw/koOBL0PKdG
Y34Ko/5x7X+ie4sKJFlqfOKnrcb7uR8nUyUAV1xmGiLWR0n3BTOHHazw71buX8AF
4IcPX1rb+bigWn6NoyRr8Y7siL/rUljndErMkzyeczXJ0yLclacTA69e8pJMnBUK
96O9kiq26jM5SVIuzMMgUF+u/qPZJmeIIf83crXHX2k=
`protect END_PROTECTED
