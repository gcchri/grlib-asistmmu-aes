`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6qfNAKTtGCCRWsU1MH3hmq3pHWN6Y+aN8Olm9F7CSgWxYvBCeJfHuyxOwzd8dBbg
yH8TQ0+aWiaDdbUNN0X67P79/3T49lf6iJh7dJO/UFxQV3CPJeJHxo0jGBz9++uq
aAkb9kKKBoR99uDcEgR93HFqukK24YhwO/cmHHJVSPEkH75z1D+cR7jBm6FDRMp2
9F0Bu54QrPg0H89TtX+WBi+EUy06t+46IL+dsGr7cObmgmYFNny6veQJX0eiwREq
oRWpbfiIT/AncT7FZKgyX1o4kMwEBvfKN076IkW8eGfYxGrG+N6hAALRMxk+l1Og
BVLLz9hEHMBHossJql0bOiw7AHLXmnHzL82GESLXomIIuwX+ltm+mmLjF9BzRvCt
uGXmkhgpjnjHpe3d2B8693bexTEQG/mF69liWkG2TBlC2BiMutHmjV+IhVvQSQmI
txvQyz2g6erYMk5Sp6Q3IjiM3QwBYc8es5olgrQtHVVeNb6e75srKVmHAxHkGqo6
ijIKYFRBMhjUQFv8avrHpu52EopQMybXKck0knViU2ULcae7l21O8HfSTA8B83ns
l3lnfLGoUnNHNr1Ck2ldrdtMkFMvDq48sgxVhknPOArFxM2Ln57U/fOHiqx4IbgU
JsoOLK4vbImh328nWOIFKA==
`protect END_PROTECTED
