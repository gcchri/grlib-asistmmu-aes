`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QQ99wiUbug7ysFlwoEWLeWMgF8WmeOvT7emotWAYwlmHifjovjo8u3huVJ4nqPrH
BFv8tpmg02LkDmobgrhFY+DcE3I7J4nSt9k+c2MEeuyUx5+5PwTHe3xPq8RHsLgX
hapDShCbz5ytHEyil6jCNlWE4kNMG8tLggtH/lpGg/R5vroHDYjgPAhfH/OwEfEd
XVcySru8Pxi5QV8E/HtBbJ59mIZdG6NeIX2SXcpirEf80X1KAIPz1AKjSxGZDe6A
5jQTsyE1gVfLDdDGmqdBCk8qS2j3tfmb9Zafi27cMjmrzFYshDDNjNH3aeC0LQar
GKiWs8TKfU40ro6afEjF8Q==
`protect END_PROTECTED
