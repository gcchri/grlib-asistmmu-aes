`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5aOt0ECf4ALxDW8cT0KU2OIdXV/piSAW2gK0D9glxaotS8lgom5LKymg6U67HicL
9v3AgsA1Pvt742rdl3WrC++HRSt/B0F5P0dGb5JQUE0Hqm3wpdyothh9FzJjmlHA
La2dnFz7XtW6pUVAzrb4hwc67YLQzxYQdBkSmbLVSGllRrh3BAoovOi09iqu1QlQ
24IoqTo48UPdxfW4x7yPPCouCH1GVxec90OGfl3LI9ogneZ0FNaoJgQwd0aZzAy0
uT0r8xbgP97/VkhXDGIPyGO6NOGTYzqcGDMEOHxb0/fTBnVcmrWLILpjhuv84J0n
mL69SYSoLeMUvwlGLRHaNKgUM/d+Omx/NMB1s9bqDPtuokTcdnCtA8J25FVM2qs/
5qp6A+DZdGLie359fuurtDFnFQSx4Sr3/rPLAmtEOuOZc7ExhQ3N3U19p9W6h0Ti
dVqU4pJcRue096RLFLAm4F5i/ywXbNVtiWZCVVZ5cBIpBw/xo22nxdPKrUsz93H/
ouEaIz5nC/YBp1Heq09kXgYiysdh3Dhq54xC3quHBV19a7hkvzBTqKNVqqqHvoCh
+XbOX1zloDp1YIncg2bbylD9dmSaPlY0NYObrh3r/MOQpn/dIvb7qgJ7Dn/pVZ3v
+/lffe/2e4ygn2JiQrajdAyaZU7Vjifc4UXr/oSCwf2Lj/XfpL66sdaJjpRFsKqC
0ZbzdSg7kTVqnyshzaQHYFxBBE+qB5DT1EHoKNX9VLjTDHRAEK1ngQTCsoOchFyI
TL4XXauUgRwa5594Q3PQ7ztijqMgUgQftiycn4KAgivo+jZw6tQAqLVIWHnLsVXJ
E+Qbcb2dH/Hx6+KFimWJbvPhP56SM8NMOitWtNhIH8tRFqcBwxuGlBQNb8hluQZS
y1mHNMhYnDdRNQSp+VDWNFaLC0neYZW5s2KYt1WsA9kOmuwWpy0Ig6agM/a1OJGI
5MQ8gjvYVdPZyB5IR5NIktlpmACDeIbTg2jdUlNttSRs9HXNpRtnFvMP6pIZT0on
kMk6ZOW4cq/yiONt1db4/ai1rZ+JZK6brtJGsI31YOiQmsq7K+78g8WlstcAt74f
sx+jLhQrzBCBD9p98T5lqR0fTblv5nT0/8unkV1o9DWL6sp7ztomZWUXNe893j/z
tD/FEyXaM8cXjRmcmRrEJPviOtNx3yT2nEabWggmGXdKrQhpXU1wOMqM87+MGXKb
vgvhAAEcvgylhMxIRUIpg3DmsH16KWq3slFhHwLK/yEbwHff/vrWuHdQR5hf+rZD
tlekkp/pJ7fLospMoLe1u4//I25giu5bYbtrqtjXu1hUenFjJ+dGzcetpBWtPoPD
k0WYTLm4A0WP2287uhuZbGWUWQ2a4w9Aifsy1OhZifXClXp5aV/+JnxDd8c1PSRZ
wvOmlInh67pYCLvAFfNP9Tz8WWhKl3Y361hcoMEeQq/ZF2OKAJMqoDhDZYqsLZIb
iFIYbwBq69FQ9Qvlp+ufdBExQCS5e6hozQULHO35PG5MuMJMBthKXjR/QjwseF3j
Vy+GSX0Uq+yBLhE63m/iM+D90vsQ91Wmhi0+4vnUXlSXJaRfAdkpu1uBFC8dw/Ky
Lndrorsoryg7oKikwXBJ/DILteytoO/MCBMiY3HOWvubOU+F+9FXrsbUODXx2zHY
h3DAr3z/U++gLKlWwROn7abuA2Q8T0qxwjsRbpMiJujaSom9mvbLUWIOwCsMuTKW
GmKy11h+y2olaOk54IYFrx96WuRons5/ftv04g/vuskkfB5cj77I1MkqnaZ4vOSo
USdu35uwcyfPruhyQYipdeJgROy3eIet4qT32S3B6nEO/lM4SCv8soXbCgygQA2x
kPbtmaBn2eK5BxPVD4LZ7krcIh7xAIQ6/+IKCG3Z0LoDth1uGMcsRl8FAobIikkt
LuDpRunpCr14+zf2lJk7oQ==
`protect END_PROTECTED
