`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h00VNBwj17dweN6UN+BV7nq57ZPDlxPaVJtenNLMS86M2CJ0v2R5pNferwqkgx9W
tHkefgg82Ga/OXO+cVOp6fUKGYJKOVOpqJZ3mmrHDsHtlNIuC/NBL9Jwt5xZR8eZ
ocHjQyIuDPoOjY6zUPgnOej5jZaS0peTl2dZ3oeEKUDFFhZlQIjgH895Ra9Ae6to
bPVg5b/xHS60fd7av2IkP9vPFgHadu1igKAPRHwNA4FzulFaw2q84PoBaMtKPE8x
Pzk+92UiLS/KauqTHvBNXIANMPjVeKRPXv+5nEYpemrlN3J6gQEUajo+Ip9SRQnX
nswzgM06KfGGpo5RS8eVQQmYOnn22bhGnwCZmOQ2+7gzlin1I6BCyrfKjHrdyst5
2IiMnCnnk4N/cpL9NElLWQnSEiqzDBtzLndRyDp45DZCKbHu7YuoHzizk8WSXevT
LeLldl2k+sGN/klqzFgubp7wdJCZ9dnMRtTGA3CjY0uS5dNVd72kdvu3ZHvwE5WY
hGAv33Dr0klL+KOVej2CdhbB4KwbCsI6shUwIahbDDf5579Z1XEvx5kIGWIIF+0B
EHdU2F8tpMiOGwpXlRBkZct8M6WrIIGzW3oYeczLJU9YYufbPci54gzi33EicXWw
zog9poD6ekilMbMg4pxC0tvXikhDNO7+phZXdc5uAJmlqOJPbwkfjU2lqT/pUr7j
z+t7kufHUxl7BGlbHTbniB0jW3O2OZ6tqq8ex58+Vg3WSJdNmT1tmvMuKqNfXmSf
5llrXh5MO8pXFjvyUpNButfWr9rSe1PwpVAxGCSQg10YGc9ZPrjA/Xm0uNLjbgyt
jjHdEFDn22tRE0BusPBm2aIB/EYhEoG6bPLTmzpVFYzr7pJWiKYQgQiGseSziOZP
6qTfmK2BvB2tWKwpJJHo9tDLNe6mrHPmvk42nHliVyKwXsc8VxaJKapvLG0bdhmq
P4voqj6FO1usBtq/fQCOjGUHhC4mA+hrpMsDnkmAaF0JjCA7fhzK0fIu9d3oat0l
/SnDG/C31W1vvWByPyusmNiNtt9Zh61CPE8zGJ4TdjSN0s9lORwsw3DxlyG5445N
U/nln9IC5WGw8q1Z9tFqa7OCymxGY5EQfJHYZxijMzgKwGqZ4WgvF6ncuYbLpo8d
RjTwEHYi5dB1Tia+hxG3kghJVFHVVAgdoR19RjWFaEyegp/sMdgy0ehycu1wAeXe
/65IZj3rI74azu9thP2xY3K29lYIUSKticJyiOZVIZXjSMOyL9dUzh2DoqmvvKkn
86cyHSkEEOozsPckwn0nBLqwU1ECombebj3S6735CBfwj4wIpjX5GxLvQ+rIWasJ
Cb8LmJKOFUfkgj13Onukuihd7A7YuDNqoIdTnb1XBVxA7ZAI5cgR/IzBQa+tJY0Z
9OdhHCDC9OuKlgFkDF4xVn/XCha/jsNOCIE4Yo2L57fLbo3BREawfPJe3toXytLt
T1i+vdATpFYUHN9dScc1DXSq66VQseIcKW+WXbPMRgmbOmizi6zNfmn/Gy/p4358
+Ab0D+o5KM/Ezw6Eo9JJpUqWyzYcP/KForbcoUfvNA5PV21meCPTGm9/zlw3bQ12
V/yWK5dc7XVygvlEyPgwzdwvMK4F5KQ/5Olyq9VdB6lqsiCq0lVJxJMmTcwfHmza
ruVfxV8aA+JcsGvMlV+XQpoMJQ9P/xqqnK64/uArTukjIJaKI3JKrl+B83lvmXvZ
Djyyto+Ld4HTI4yQ7M50mxW4JDvOHnoAoP0VIPeWtmXvqe1/gi63dGPHl6nFMVIf
qypxRs23OXPpaN3TO1QkzRuumD0k/bJlwMo+zyQ1yIVjpO76xJ7gKj2dYNeg/CXl
g3goI8o1BMJLyRt4XkIEcwoz0comdWKxixBUZpqfbixdFCyAb2dEUaRT5Gnsj6Rg
RBUwsox0ZPYzNGN7wM/UUwyOVKJ4q9uPxNTdpSqgE2mzDOgY77gLzLLngpSI/Fq5
GF1UDZ3J9rj2bIWILQldK/nKF/w/i+yKqXcTzZvqotD6sv+WIkjlaeGzMkRQrYRJ
aYGB0gOghzPeBYY21IXZWZX7AzGC+sJphAw/kt2iFXF2FA/WWzxSYL6AM73+Kt0z
Tu2/usMggBcrdVb0TxeA2WOlsGkXfh8Ld4aEDwPxIfXZ+qRMm4ea4NFttcpNuQLZ
Jp75m9h7V3ESXQv3Xi1Rc/IXH4DfbdhanYVGXygsCyxtIxMRwCET6gbx+zrDmd/W
ywcgsg1Nb0cy60ZMnllu53WIOy1G+MaX92iYXe4OsynrogVMqDEjGCzNtu6KahUd
INfsTWNklVurZxc8qfQ8thEOhJwf/XM270aYe94ttx487CYheqWDhlhfmTN6ZKkN
6q9CEkoZ89DRq/+E8dppBsg6PBzn4YkSiTwLLjzWdyOpYLwdaO9JiTi6vvuAJAkr
cgQfANww1AjHF2VRXusZtuWxZXwOXNt4bTkS5Sby7iyk6WO8HiBfcBVKHhwQQebe
eRgrazk5mPF0ycMHsRrVOfrNtejwPvG/PFXQpjSgHB6RjPcUVNGTC2ridyek5F4n
Ljw2l3E3LJ8JxgkQQveuxw1sHjr66sb+l8xuPrcSPuq1c1U2mhUG8gpNieM+Sgp/
1fLXFlLkRzu6+llgWtlq0BJvVMmQAwdgEyr57fR4AoFQ66bbulq6v61MuyR8EyfC
YIxsuy72Q+HTRh1oE3Wlag1+hhfIGoXkMt0OOqZRSnyku+Iw6zWTZ17jCbe9QiFd
dJbckpVu1lp8OagYZbTIzIdUMOSFxwGgKGvuxUuHngTA2mJEePrTKutdD9ygXIqO
g6gO1NTfGNrXm4Man6u9bf/iwLR1PNqoDxL8I3lR1uSkZ7KKInqPv0l5j+kLc2Z3
t3gNibO7xXj1hXoGwL/opaabUierrIMX9F8XqgwNklVXiTV9DVu77Hi9Zj0k2+lx
onvrTOCMD9qMJ8zqVn12r5WqgjzHDAAKBF0sB6EZ0aAdq5yCRRZHpoCUwPqL75lH
tdwu7vRkYn6c6smDlVIlWiAl9nu6LiwgmYTsSwdCbEXhnopIsUdT5rcce1aFa2Vw
mvNVOwBdxgwOGNv1ZyjKPpbae3ZdJdNXyowxNOJstfcM8acDm6V7z9smtW4qHXKD
5eB9hORkT1+GpQsafY7Dr+GBBFyef3XJGagxKTqHhWDzcjv3SP/VQezFid95pVFP
Q/MWtZk8vWQW9VLyUVYSpQqHKXz+Hy0I9WWqFEtujflZLiC40Umi8Xva3G4swrtG
yVhRY71Y+ll1mfMBbISgAiKU1fhd5Vk9Z4WwKEQzUc5QkZamuad6lyFLdi3zwIYf
oOq9ioWnNGh8GzeVBy6DAH4+6LrSLJ3Y6SYDK/kml3AK0f8qTYn1jH+BxUCz3FIk
9TAl3L4b/SqmEL20nj12GJ1xGEQcwDK9MTpsmnDDc1KsnMC6mhUkG8wDFLuC2QVN
jBrKzGl/76HrphKWJek3Y0QejsfH39W7k9gaVd/Z/1HMX5y64xk4dVAfGs2q7WsD
iXNDTkS+W0m0id8PzDbw/S1kQMyW0LTQMiuXRa/9Mj+5h/ULK6eRuSOoGBXbc4st
OPyoEprkMXrM8OwM6xbhTrdSGKQttFFNKS/c7eJFbZSWHzu6cHzLVvLZLiaPKYnR
y3WCHRHjROI5AXxSaFkNJVk+TTGdbsKlCo0rWKJRRT0RrEWqyTTmV5aGWLPH+kBo
Hk+KiN2UElqbC84FEFPFEBkK/MLDf1/9dM2corIubf1SATfhbFsAq4kZpk2bWbUj
WVcrUpj4hgUFdr9WKPB7DZw/lLE/LW7FZUn7Tms93bdbm8N03cGnfwYhMpfrn+LG
BGCeJR2pcZgqbtSE79GksEPNdNKuA1iKwovJkOl+sJZ9xSXHEiSzMsQbYAAd2HgK
GXyPo4NnKN+dlH3+bGMO2REm2vcQY7ezTSOaiDcjebF979Xqj9vU4yyHm/wZbwOZ
z41fJcSQ+lbWGA2JyXAxA8Tz+nnSr3DkwvosqGwJXesYwVFMENOvHtkv1dFuw5gp
d37OKkpp00uApIS4Du1qddpcNi3i/ADE+rLie2IzYHIOy1kdDc9DtCKrkVYOO4z8
1R4fXzSnmLIXDzfMnEqZfbd3N8x2Pxxhq4TcwVN4jNRPJITnen3TFnhb3opKUcPM
75+EzyWZhSfFGJckVCJ7LnbvUeL64j/XNDMa6bEJqC3HlNvRs7V2QruOGOftV3qV
SdFXvCK/B8QVJV8b8hShARi8eiv/dX986PWbwG3Z5/vdak1WCPo3vorbgZxvNu9M
0kt6DOjCNDsqnWQ2Clq1J5urUjBR9Ox2ir5qp6lA8p5casbxsDYaFQbgYtxZGELX
jtx7rX+WdR+xYa85lQqwCbKAPEwkSBwEXS7z2jTi+gnxFNjFd6TER3qbMd+NSctn
ofcwlAQ3/SY16zAlkhItA9E+FWAH8zSJWTZlt9jtmq8GkW4MuExjBy+ZlWCcrlmi
/GuVjiJRHYQRgGrYaJA0speqD6xCLAqbTF5l36KOkmpdD/dAt4EAKqGI1+50lufE
6AuXPi+AolIcXRMNSwJUkOkCq7rHDyGX60NCR2qlbniWGRekKaeIbaOQPjWhxoAh
N5qTUhhNvRPRjXt33jrDOd2+1kRMdLXkBBJnS7Xb+u2rIzRXSb5SlLODW7A9oh4v
BFsVTBRLEPk7p7SfoA/8aNz5wY6H7DiWmkscg97EXUVNvdLPXAjp+N3rh7KnnRmc
3v+F3AvyPrdFSM/Qy/sJwAdkRzBCcCxVbDF0/6XGC2GSKV2rRgp7IV9lNnteP0IL
gqEYauo0GPhKqJlf4592OsHoAVSR1WZ81g2+YcvuHEuFHQxHXXespSN88KsZp6st
zZUNrqMIaYUsg8QLIzjL4k6mPWmbvYDzwM1OL7EVKzD5thyDDFH+f8C4t+SBbhWZ
`protect END_PROTECTED
