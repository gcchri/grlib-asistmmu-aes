`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HevJ6SxWIB5UswN0PhcHNGnlHJ+5ZrNUitMWgPZK4HDKfyB0DB1l4NtTKX4MF6+w
iWCj5kGRTiB3xRRBx/0bCwgZ/JCzx9jMiCfIewnfQZPuT+2SDS2jNJiUHCZOcTGt
MNweaZ88MDkHm4jNzlvsPerqFQ+L9EfNY7Dk0Cy1D/4Klzaj0YUtc0OrX9inb5z4
V384Xp2Nd7hZ9ucdopBeQ/bMd8UwkYAy3/aaEdbkXQvtUnsbtOhaJ3+b+LLNq7i/
95knP7Ui67beXzkTEvbZvszLVHCwuKSHF+ODW5l0GLe1wD3MriuPVOycc2xRrnoZ
FaS9uBtnD8vhiKd07hF/QqdB7e1ULdmAFiANqUkWVkSCSR+zNwiGvOUP9CqAi3yM
IJT+jzalk02nBCqoDqAAxqkSjjJ7XsvewrvNnqYFLZegRabGotcef1C0V/MzHTxV
otwQXgRrWSD7JEvp5oYzNJRpTBqFRyZ2GLuqm2zq750HXNS9LKT5U380N1hWCl2L
JeHM5t3bB0xIDGjZZ8Kee+itQXyncv6Qhzq2Sw9haiIgnrMASXlcAlTv1fvhmGL4
DlOfNyuv+nZRkPXvLhX0pu8qDfcfLPWIud7z19bdbIaJKdGnUnVvcEDb7WF+IdBh
x5mfmInRDibcR0uDUWWj3A==
`protect END_PROTECTED
