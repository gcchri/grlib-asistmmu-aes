`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RAQoIoja/0DAIpOJkm4GoXnYQS6O3lguVCjsg+dMurU7yjIAUA0xTKaoauSgBPas
JArKc3NzLrzArtYgT4gvnTcNd/+WPAskPEvfnSsOpKmnBIPvzxDlYXeQwQQPSxgq
luv1yxOQLGwdMAkI3DKp8Us4UPg+I8UUyKst7/V6MX86rwE4ZxHWlqlofB68x7ha
TArUZp0pTP1O0dh6SGAwu5huHGM1Ys8R1ZhXU4P6GZeWSg6i+RtXdK5BGhhgmwN8
ugLIZgl3kT53fCLk1JhihAS7zGnGs+WIty6k8VsjV/4hxgWjUqGjmd90Svf+qxHf
dYk6OHthyk1ZTncCa9gMXFPlJ1ue8BK/NMaQvWV4KBnWZBYgRB1QVGmjV5kYL6s0
ArlnbE+sT1lgJjdFB1FxV/OJn0Y1tvZT1XDXsP2ph+njnm1EdBvM8fF4y0zAGQll
8zvt6UKe+C9UYDqLFh3KEPDcHKX7X2KPqY35KrsA9lLKxaG6q6Aq9pJfZmDRP+re
7YaBnQSdQN8EHgawXO6BeiQoSoubAXBJWtRK893EdKJKw53hWAw8OnhqEJykoziu
iDgaEfL9Dtc1iLwNWSUGLDNfc8Ops0GMrPRUhaujuWAC+WBDQbLsqxmfqOln/MCy
O0x95CPFEkq5vXqbNLwUqzJAPocAx3Z4ZGC5f8x2PqDvdXcA8FauJDs2wScIV0QJ
CeLRunoY4JvilKWSYRirWHwEku+ir/Hb6UYfUeFU+YgzLRTOlV7g1k0NKeQtUMpy
E4wwSy/nQh6OP2lcKXeFgtswAXoi6Ccwt2eRZvqOphBvoe1X4iEpd6CM7X3chxcx
6d0wok/6tmhlFiO2I3AajEnJz49Gb9lNBm781cjitoF2nSqn9eiTEYf4tECWRpGN
D8INhIFSvCEOfIAz0RoHX2YkSG6WENNCGimIoxEqoK3m5H+kmdN6K2kBF96uMNgw
rtECijpDvHuU15w30wAtkvsQikSG2PMgQ6D+oUKYFch0ertn3XLjPN5CpRC4aFLp
FlHGY09KblhNMQQZp/2qOiLCjfuZ4nEas1Id6dEE1HkUrhMoWZ6m8mjtgHrOqPPy
3aYgprB9O2qIMZcgBNwpIzAUsH4DQ1Pwm72an4RVnYZuZJ91kDbvjmH14U2pBNsM
d+ClwFKeyD9C12xXXIyoAh0p3phtzwncxImP+wSwFj7ms1v7TmyKg/z09mzJrvOQ
D16Mhcwwhx4ihlPSb3grlbSbioY6/ELmWV32BZTv3Zdc/EwYds3aeXr7v1Pkzz0A
tjgs5UMh2jNJlGpN3FgW1W1D+R9fkLO7dAJtuH0AvASUEJCBtFxN1QxmJyN4YSdW
xnBb+wbORFHg/Kgs3Z8+7DmKyaFgJ2Qa+gldY1s+aN4NRP9H811CQszZiaZazR77
p/kgx13RnMZ47ar1TtY0Kt7XNXfYp4nREhfGVxymg49PyB9qcBcMClhXrES5hzKg
sn45URcULgi2xbvnZ57MecoVbZc3BGMzpF/RtN/GW7PEPKngPI1UQ+xTd9kLxFgz
SeCEfsCD/mD4LjRqEdMbpm+YcOHSxaErt2ZGi4+v3nA82V6YgPSA2MTON5Y98IRf
uwtVV/6OBFFZY2pYCPirhVDMMsVPX/qkr4w45XDdWBIGeo3dirKR14JO9YYqWj0n
0WgbBSDZNW55OjdwKTOCQSJrRrKqlIDdmpbII0R7ZhQ0KRpZu4j3R+sYxv54ibSO
D1cFMYnagqSKW9HLkoYGBQQILbIK79wNIG+5ZBlYAkhaevs0miw72OLPLhVDZtua
5PhDgGEd5j8ureOC3ZjlYiDaGgmyONF9DT1pkWpVkQ73l0RMGWZPv0Pfp3F9oqoP
Uh0NVlvuS+f6KlsJVSGiGY4oFv83bDkyqP51eNjP11JoUrdhLsPZYrDzyMQP1sed
dt+Lnq1vLCUaBYQ0eTiclUt9E2aV0SlyjCzhMHt0k2Hq/JlgrxXVYVdxiXD/Ju3L
3hS6EXO59TC4sozRoUtidR+Prc90oRnFcwbqlLEu7TEo/m5qJcQUcwQL0k0f3quz
LLOoWHBBZ+zH6E8s+yV6K8jROS67fjihdL4/vqlprzmcuNPf5eVLrCKY9D2yWvwr
jhJxq53djpgnDDYpwsv454Tyha0W2cVMxYiwD3MsCOAKj7C5Vb9+rmdi9QeoVu4O
4wdYUV+RiMrBAYLbnY2T9gEEjoD3bkKAmSPEvtDFP8MAA1gNIO+0nxfUBH+ib1k1
z2nU3F8E0dzNFPO0EmBmNcVhlyqtumiKc7Pvj5OImqoSiRnqsEyrG9i6KLjX1A2S
842kPbNxp8BoMiZHbRvNxfKVKu1qWV+Bvo5lWXwkuKiNi5J4YRy8NyatDeYEQImp
qDKpjDVhoy9A9HCaV7JCsQsqkblpx4RLjbL9wfGD/OibMm79AN3osKtaPzjZtUlL
zNtOmLNMsscJWh45YWDCCA030UlJmjnJ7rzeHvZv0VBimKYFRjHRnoN2aqWIuc29
/PFwDC6SLPkbnyTNTqOqihOXAc9bxdlZmNwbTWz/pxCv0AOiEc6VCMijlikvuFqz
eswZRslv30oQJU9hGkzZkK9YShQIDVKQl1vUkGR1zJZMv8RZxApfhQ27O9Jvd/WY
ezleO+KeUXk7QgXTpQNpM6HOrAyIYorW6hVoTKzLm/ni6mYkvmhEwh7gebeLTr61
guHlLZchEFmNpxEEd9fPxILydO7szIz8/45SkWopAOaUgLzBrBlaNyI4QExpQ7eW
ju0EEYLi46s6Cmo7ccb0I2pm+TlcvJ2HsDN24GhGJ18p0u5k8DtKgHu9u6YDbpVL
p4TcvvYrayeGKhwxRTHv5hmQZlZHCdC6VG0CDBVt7CLIfk6ouEvgm/cYdFumgQMc
B+pH6tX+rHN2PJB1OZcK8p/EdxFmdZ79q6qaDQFm5/FgWpwaehf80ues2QvGT0KU
GzUcWrIqmB73DhvWXafmSwHs988kudBX+lHbOS/KphCfV5emgnsBvn+6Hl2foyIu
Ix3X9Q4kHeURHjiIbm5wBH/HcuRRNVQkihab/gWqxOqnjxaMUpkjv30cgogYTm9v
sqrMJZjlHUSuNfRQtJkCdDVjBztA8GJZz2lcDbABBefPEBQcl/zi2MRYS/uO5bk+
SOOeTr2LLNoa44QRf+ILxs39uigiNJfHydB3zWnYA29EltmcIL3Gklxoep/4c+z2
BsastYyufgMbBVJc/iu/+b7f0Be7SgeWsRy86139Gp1yqbeY7LJZPK8Rw11Fp0Pi
Qr9/Uk22onpnUsQraqN3fMfGd1/1M/Xm8UnZ3ZzzlmOhuZWsNBG1dXu2KeT604O8
9W3b4KeDGSoZFIDaHdHU0YIh+4PV8r+0YNZrTKu2Va/lgGudoC4NCe2MQJWjeTW4
lGNJTkFA5bniLsLEWVZJWfW3dXgqKjqhuHtqT/B2+JKESBWY0dKXYCvgFDXcv+pI
Mxkd99IdPkzYU94MgNnmzDVTdcBuFT3CWi308iK4L83gLJkBF7wAErRaMAY74zcq
CkmQWt/x5O50gpzM7XsleaJldtUogV08hiIhpjaWAhniCu73yttB5uMna1mVY6Om
6OeGclUWZkvOqRlK5s07UyoMr0I9X0R4NdQgkXt+NYGcfLgZGWi4UYQPegpzQXmW
u7+TOAl6C3Mo2aXX18XWxicNGVk4NoFidvnwkEyPs9YHXY1bw8MlbNJ40Xi2/eBc
A5+lUo07NpCKG6xpoDy2Lt4Xb1pVY6vpYVDxclNCkyWExp3tUpB9az/vgrJD2yLP
ot6dFpqTVWkN/Xv1A77RkR94GApkyo48dbVucatQPKgnDL/Bcte0ZXVmtfq87rhr
/dTAb0B+TrsYxZS4pLhs3pCKqt4jgpNC+cIk72tZjc7GQ2pLG/3nYKZNUWMLi699
JqrbcrYtENW4YOhAq9tE1lJrU1ECYEJ5Nywcv8T/Pl6iFGMBLI1qcVku1Fhc5Njs
GRit1MrxORpVtPFrDGtlUtkJjhH93ufxyYYfVrE9LpUBc6+AjGgfW4IyR/mOK+of
CXX+/Mmq+zBmKdW7UyIJUc2otq/xJh5yE9ILSapsPpijkT97tBNTjn22+0e3Wgzu
rSL9mTXtmqxy4hBa3PkpkSZ/+FeayW0re/rWRfGI+XO6iZrJyxTF3wjdj8OCpHLs
L658iYcndLxjcNocAtDu6qWiCYP8r7j9R7QrLPN2WxTdbWTjoZ/H3sz66/nqOJ46
gNvHFERtS2m+6lSDAAfMulZzBhMC9zpg/8waYsgljdCyks0zrRV47tz2YM960KuB
OKwC+5Ty3GbVsaXs/rxJXeK2hPAy6xrjvHTtP3FU+GioZcSoDKidvOjKwtiOX8Hb
PfolPkUDBH3Ct9LClLFBQk0JilJtj7JVv+IoqL7suxpWB9Ciz4ik7Icw3AB1TOqz
SmptAxjBdGbglAJjq6AIzHRofZtxBc4pd9xJJHX8L6mHpf+VAcwHn+Hm+DF9ryo0
Q4p8U7e+3T2JOzKRwzvnq4westO6fE5rJBhEsAOFcVFA9Wb9gIdEMQR22SUx4WlU
Yn3izEIOZQkqTDhF4VD441VGoF83+NHaaWjYMnVJqcs75ZmRlKIS3wOUstSNe79j
YYAmI6vALSIVQg3mKckC418im2VqxG9Skzm8CvBYruNGfm3qsqY2hcCEqiTxNdP5
fv/cYcHzgXdbFetHishgS/Nd5SnXFJ/KHy84M7i4+l7Cfkdpxs6Ptvuwyt3TR5+D
3z3ACeOYhHpuugcq/vmG5zFjCa0QrzxD8FYFroU0J6wYudl02F6ge+KCFFYpYIDQ
O0VHvB4yz46SIp0jhcAomBF1CDOLS6Ho4Lpfiag40cPcglhQ10q+Sr4NFP3Qe5RZ
CUZ2K4/veXkGHO/mL0GfrrWnbjeZjETuoES/AkFcPyIvh0WI5UVVgtwK7v3m3TJh
YxMcnIAOY9aAVCz4EkwHCgWXyJu/mZGD77nRcurOJ3WReHALdMeyrV73uBI5Hjds
T+0ZbobZZpuUAJkVKi9eQ03ER2VpV1ntfyuHHpolVIsRSryz+PxrqWHypl6fQSbq
Bro2087LStHvHms+vzoVZ4MlPj6jOeBl7SoVx8BzoBf+DSv2K/IKZdS9bzb6mjJb
mS0+kQau+8AEndSMSnmmIUT0xXVaDvJHiV4p18QbKQKHeB204mwaW/TG8UqEcc3R
zX8l43fjafvZ708UYk5cEHr12dNCE/kdvD0HeNp3fPBmG725abZMrYnE9JXPS7iY
9ilwYBSjdzwonpKGocd0yJw1EWS5seZ1ew9BYp8UfZ0uBMp6k89jjle9fFxHwtpM
iU/10XR7Vb8BAnudtpLTVdLAOjZBJ06dqtyaqGDVLezfjcH9d8ihBgILpQTnyN5M
t29t8Nn+eTPXnTDANUhnC8MVbnZFtIhb88wS/+cD6RIBl4cbus6pp1Bv86V6aC0V
+2LXHmXwVWsuys6P++h+YWQdWMo2mGYqznmuGiv1Ma7YIAGEepN0y9CXs8kFfUuQ
UcP95Z1+T4mdt+0jWlMhDi62CSD5K5bqHFBBsl0bTPt7qSISrpRJGWzH4NKf6OPP
Oaq5222MPqAU1Jx+HhNeGtcll83hypfyHerY7gUoTorg7YTtCqZU/o9Rgheqn87b
pNtierCgTo9/ox/AmV+JS4qVYoj3Zud9/+8zYJmg0IroxFLGXPnnQrFg8mWjqRwE
llCfrYVYNVgsDIRdjKtoRdF0RKXUfP04vlq7NUR5dyStlIo5KUw7UnzMV5cDdmfQ
z1WBQcJDdhDStTonpc5BpzAOw/TChlA/VelcrcQnEoWQyQRm7xO8TFBKIIih7RBF
foMf6BZjcRKn29dQAIdDHZBE4FZ4sSJyd3MDurO5XvBqYBEdPUqcMFVbLCHcSVci
9970T8GsrP4nTpwXYteTKilITETBgSUXpCQAtuMoVzZRUPmaHYYNRnp5inNrUGmd
6gMU8YgzjI8K32DkKC8ZplPRPYWnU8gL2eLpkAuQvz01QnCdzM7l0qNFeURyamVe
39l8F7u/SY4BHUCI/zO/GK4+RxGxGTYgUbpoUGac/Byf21QvhC0E3kQKQggI+Tdl
OgvXgX7YoaB/0/GvPQnkfzXl9xIO04FfZl9fuZdvtOe4vYQT0uoOK574c1C5PzFp
mflUaKVHbWTGw+TcCqrTElerkERgzBG4Q/fLzVopykwV2cixmTZK5A7DV1DDBc0f
gs3Yv61LvUkNl0qshtacIQBWwA7RwWtJmyL+g6u/AgyWvkysP85M3GFKbyw6/FhT
2IBJxX3v/oUlWZvo2ZBHl66qv4Dk7hCK2T1oY+F3tqg2IaZkkSmVZVRDxohZZ2XS
/COLC33JzP4niKD9WfFnX3G/cRDQ6V/JXw1nErzCtiayjBG8MK7Gb4LVkiK2qHUG
d2ZszesNFGkmQma4/NaO0ygzQiFYjliX+FHOIJmwEDQFZLyqSkS3iSA5YpiUjhOu
o12Yj+S2MPd+4G+o+YM/dtJjgaPdflI+khAdU56h9ssdUnnNiHHmIyKFeqcyf0AH
MMpCM5zAzcMGmqRvyepg/b6cACPH6LXJfv5qpRbEib0SPssNMOSWwn8GngxO0o6A
DRUQrkyajyaq3T4dn+S8sUszSetabIi0xDRmtNI3sZoezY5UlV+1yvAukhPq4EnP
JQmO2CwvgaluATJXU6RoEKZHY8sWJJ83tAfEiijt/jNPlq9tQfAqln3d3TfbNhCc
Yi2bmMTt/FBbo293g5YdTcBOQDV5uEDVT8Q1XeXk0mPQ2+qo1HaXu3Lv56yMQ2hf
ZzVZHts1ZudFupVcbM+kzfDNpdBI1gDTLtgP5fc4qYuiiTsKI+kILVLtMjags1JJ
AKrTn/KKWfdaijLKc1NtrSMKY58nYAh0Ud3oRJonJgwJBXrY6WP9r+Lg5dlAQsU0
AUuhtVvR/825bMoa79YORm9MLXYCrM/yzExWqYKliW57pOFEKOip23xvdWRK5zP4
DT1voIMyHcy8R/XwG+ixuJsoAmklqknzk+reVzp+6xRGWZk9WAY1Xa+Adq6cC2Sm
4mc7AyyuRyksFXQ+AT5PHUkGghDd3PfPgS1eoyzdQ1Rotuht0EXMOUQlwAbopYe/
YPeFssNdCbiwy+J2nz8E4Ct8xoEFA9UxctHEzfz5Mt+ZNVtsZrqdu4PlU6Xham7R
6D9hQDEfiDQ0nEspZ6whsGcun4UvF8okHA9TaJnzECB6A72MZvRO5N0gqGLWfAKW
rjrPqc4vIIDrlydzdVRw48FVBvaQ75KfD4PLExhBPdomSqaUUASF7pf/G33VPD0K
AI6L7+hhn9Ve8tlTfXZ0BjyS3hFDzw5uISbjpXMwUs8mTcZIhhSfSWBTv7YUzDC0
bGgQvHsR/bBVtuv9NsQDTS/jDYtq8VpM1HUEtRWO8LzY3teSlgh83Cke8NLVkrur
ALRB3v/f/1XwBHl6M1gV36N8F6l7yOsvqTztziz75gUyXSEyHyJ4MGuDrfQfwHYR
9yKhMhTWbVJNvoq64Lzivi64kPPrKq2lsgehVwpAfa1NS8EfakhSQDgUCUhD5zyZ
LO9nXOQdZaFCYyjY+o+ayU7i6PoBEBw/7r3d9RVFjbBjAXG9PbeSamBoJGrVIKfH
vLaHbCvv7UI3Ld2GOCAJveuq1zKBVsCXU9Tc39JdVTRUG8GUYN0PwByJFa43XrT9
hiCvPGayHWYkVPG7J/4xeHgfhl8j3fSaQgKI8vY8OERhRSOzP32qk3/nXrAX4DU7
eiOX3+LfT8kaUy9BMRv72JxYPErwmZkS9iIvVkaYyhAtK5tyFaVoP1fK7Pn56No/
/RJNXU//mrwQyT3XxoVJY2e6amarsirClyeRtema7UmUiwSUzaAhOAiizDOc2ihE
5wPs5vvdMRAt7aJMKtD5mLw6AMakSY5bGnqNLCEmaj1R6C5qk4DlQpmKqSTTY3vo
Y+My6CM7Yx6Uzf5kXlnoKpSrVrFYJ72JxVZ1rPY2hXOXQuAlGL7DBoXhYj3sgQi5
QuVL/f5hcp8pZ5Nzhy5rbKlTbVOuK6G6n+7DW09XGsu/lHOPSt2pW4SuYBjpkxfs
aN7EBF8GpM2+TgHITlCXP8wrHcjlMxvnY4T5XcP98W0DygEcmp7/WtA0ZAGEUesV
KM+Kct6xegE1BmwijUwtLfOV4g6y2VJaKp44UFqR01QTz+S9++h04OGozfnXzz0I
7/ZnqDXNXzfdToRai5h/lJ+jgnrLykg1dyuLLfZMs7XBTOi0/HO/tNXH0cSwv3sy
HzNXsCUcV0m/FnNZERFy4M3C2jHO459UDm0NkIMzAXHru86CdDqPujZD41rHFkg2
JgUsFOT0ZtutDSoV5GcKA9cLVEbRrwrtcl0ko4KsBUy0m7mU4MIfY8/8Q2vsvKO2
t/wXxW7hvQcQaQ7Kgry5kBoWnOP71if4tJ1sEURYwdV6EllpHoQM8V4ZmbLQjmZn
Gc/S1Dsx5tLru0ztgsgi4YooIg+uYPqrygCZ+hkheswvWYiyUt4tlx/4lKQue2Id
EJeLFgrMmmeXTxzNNkmaeg7+FW/CHmUcl+M3wOuLjhE3Lnb3rTe0SAxbzvE9nM8m
/hvI2aQL9zGBxEcs1vlLmYLXFQF+yq9pl6nJzb/Z/XSqQTFfSe/hAb/heSh/nhGF
16nWSo33rhXoV5hA/ODXhOmPZww02iK7RaLfqOCa4wZRHkGvWFwwspbAe4x+97WI
j+8XCRVz66qmZrQFs8YzEJNVe5qp1b94NnT1tmnPxA7eBGAaSN1ouoq95CAKfqap
5zBViOhjVM08R+eN4VyJTOit943HcTdkq2sDc/+5bcQC3nK3lQ70VWodm5hnU529
qMaUes2eZI+5s2M9qyNtC+RsvnFQzZcmmBAa2pQQwz6vap5qVWJ93eHzhJx5YvnK
BQP3FOezHQP2faLeMAYs0CzgixmNG+QFhPcdYErx4WgT7az6jH4rwRiDT/9+HW2/
N7e8ho9bg2YHQVjhREKN/b0snFYVXF4bQ/08iHSbLkxI4dxCq4s6q6sVP+hsObY7
0SGsIIRwVI9LqDQgqDv1YKuF1s8CBcRIZhFCbkA6ohXQTtzfJgPhaIHfNWjBKeIc
rFNR9s0QQqXHN9UpjIroQBIQXrOiA/ErpsQWUVU7Ui1doqbUPaDJiRWAaKuwRrBh
vVnVCmwc7/OwfjlXV6fD6udDwAaz9gaVzzSVbtVvBXkzeMdwYzX4WQUx3mmvyVCP
U42SiumjBNj2IWWGw8NCGV6RwhbHD1K72PlznO8mq3IUpcWPDryn+hxF3PS0+eMq
lWgt90D4JS5Befh/DUDfamzBOvJJj5Pn7ApNKWQ5tDQIJwBhwQcyZ5gcyKPc+t3s
ifl5I/NMgZshTvfKU1/dKjHBvvwZ35448pyikLQC4WEwyPrQHoAyi4OI9iQbTcpD
IdcAUGDSbUPZF1/RgNaGi6fMH/kRCuDW36cUIvKIS12xdcfWHTQxivt6N0/fZg1B
0GJGM3P1+7R1Wo+ZDaKog4q8uDLMY1zhUY70iHxjNvU84+/ImxVfrb19tbb5aG6M
l3+zLxAL5BcM+0x0/uzfCwezMmyNjrHFO5mUA7P7Gy921UzZIcR/ZxwOjQk8Ilfw
4DU5ThsL4lFZsJR7PleiZC5LCf8cUIheHz3HiUulroSOoQftbGU5KGQfNL/QhqwF
LnH9qxyapMVIKErOiT2l4pRRQ8wfVwcGDdkg7TxMtvPax+vqTM9IbHWZ22Nwldde
DmOSN/wLPcPZhMax8K1Vaw71SpysWQuCM+U6GnWLk2ZlSxKzMrmzPz1gY4dwuNy9
UPSlax0DBbUQbO433ITaw8KmE1dKnVmkE5grHNbz/K3n5Z/8Urc+1aJS1d3/Ap0n
NEiJ3SgUq7EoxYj9NFiTNa4+Z+5uqFqinZ/WlU5SNF1dt1/U90MG5IKcOb4vxiCg
SirOty/mNWxRHESDleflHjRNuTOKbNR8VBjxg9Xza+fA1R1jWSDH8rEsqjWypBS1
hkrC9O7EzQ9ARHsZiYCOgvWSlx9ZDADoZdtfFSWLRhqtzDQvXsOXbWVp80UN1s97
iOydh8ar3r5t4QsP+mb8Mz33Z3Ab4hc8zQzikHJAomYh/fm+TFIcZgkFciNLJDMx
tqKBGOJ4w6IZX+2zK2pet2q5xuAw82j1f0HK+tQz9Uv9BuAdse9YQaaaCpZWfWEf
qJddlDlF0tyVyJUZrQ7kAgtU8AsTzu+vwjWym6U95YXNeNmmFk5Sal9JoQXexPJ4
azAr0lcswy/nT6tFeo/FH8B/dP2mZsj8p26yXwIFeLwXQg0HaXuAZi3+FYHsgAOA
WjDY2bnR+a0+7UK47YiTN8ju2O/32jJSVsMyJA7+z9wTJ6K93dgPyd3GjcRhN+M/
c4Nz2Dss+qkEzBF/sJIocMKx36I6jR2+UV3m1psEfh+ciI2wCuFbfzb8pxe0ykF8
G5F1A/HC+9JH/VUf8JrgSlMAOzdtPPI+k27mXx62y6fjcGSnD4/btr6M928zCu+6
GkLaRfNO4157VoNoOnlm2aunkYclTP7W/qOp+JH3CMITxpQ69d9iQTH+6CxGm6/7
envovswhktOdkXTb5qdv1mOUC2aJAa3k1ZSbEtbljt0OFk46t8zvJoGXSYToERm9
Upc1sq4vCIUBXSWmBkt7NdEBhmAnYEdgk+KDect8IRFksLrA1kshAzjO4/IyYsZ3
mgaVtlODAFVWjkoj90eXuoQAMmrcBkwZJKmaXbcV4WDJHbKp6QpBSnFdpF4Z6Ym3
R7o/Lv7vgg+2A/jd8WQNaW4B2oCaVLTAPouWFLm11Iyoj/+S1iBZfmVXZTusMPoz
REsS4fSaodgwD/BEyQfnZJEwcil1P0wB1dnFdgP/DMFNd12oLTyMUZOwCXNEwhpP
k5uRvFCy5XIODHLpM4GbQL9K+n2GxJvgBmdviiDtjiV2WN3sLv9iG6WhNmPU38G1
+PJ8Qp0Q6b7H7gHTYa6LtHbcSb+NppFKhY6RDgS2twFMLqqI9uwiMdpCTtUAm0Zv
pi4ho5icbV0+Haf9Ue5+v/9s34gj3oVUJI9gwhpIFyv9/pRriL3f/DdFwn5DfFtu
fwxaZDa3IDoO7YRd1CpjGODfsifwH6uvEz7JqGNxuerR2gknNIDUDm03j4408MBN
gD4u64U7NR569+bbUoAIV5+9oRHk9KVADw1KcBSJUamQqNppts3cc0MGwT4y33p+
s/WJvoggU3ZMnTg3WzFNss7JNrdjwSVS/FHBSnnOp1SHoNW1NN7RRvL/YsjAnlfG
8gCxYytswXU/BO9/FhFKFoIpm+iU2ASZtLVaqzSBRd+bmC0ZsJSANawJtwyLHOxS
lyGekcQlfVeEW30jt5Q2KcAkkxusUDCr7XEnmIqoniNeiIwtPSOFnN/893zHH22C
++r0acMLMdOTM9UIPi8lTJk3jFlkXIs1HxUH9KbaqMzEPSrL7LPYyNQsgP4Jq/iu
xPV7x6mGK5v5Vi4E4M73cSM8EYHXe+y2tQy2yWbk5tuLcdVnb4EEkM+cM6J1JOCG
zKDGeQv77iW6soW0t+fyJHVY5PRendk+P+uaQIKvyhWG5NrfiZ2BAehs8cdnhUTn
J7CdY8mUkS3lZ1bAVoW0qwlrnqLpQ+9wmhA5SpyiZF7rKRZvVBcEoTPPV2mlyoo1
FgYKlxXLdXwIS+h11ls2y8Q6FSbzehNaQAG9ag5e28dlGhlKyjf7WDEyEf5MIwdz
4QePby/o+QrBPxXcenvPpotjgRRw+c00XI36lZDxtaH95sN9mAz9d43ultSTzwa6
IWwBrgTGnVELU3p4QXq3TpWpFlRpjH7F1/DCGAokRXg3iFf92Jq7NPtt2MDWI2Bu
vfyZtlTf4bJBDEi5jfuN8gsEp4dlprmJ58eg1iRhCK1PIriW2ceP66L4b+ChlYVh
VpbDdahIAxt6GaSbVVevhG6N/QLpuisJ7tPZ5za0zWBFaDHHNe2kARng2/RSugEA
zDUVjZNZl5VMkFgg2Afs3Bs/wDNSKnnn6vth3dIoaGCJ8a+KNppvZOlq5mI1OfJS
q/ucfzY+g4rwJlwjjWbcyzHNbZXHb6z746y2GYNQskBb1mPNu8RJqL5g4EYBeYvo
01MOF1dx633qsabX+UGPWoYCxZ1NgtEqZRV7LhSm/12kM7UnLg2mUDEn2xeiQA/X
cr6N7MU1Lu/Vg/KETrGCax2CL4n8hEE9THPNaBZ4r11STxioGb/MiFOwHk7Vrn0M
ThmHrHytFeXRUkwPZwb2G22m0jGGtPn1hjxFdvvNvQtwOLZRWLmSgWvlyZcg7C4Z
iBU29KzVm5esNLtX0s0l+8cOXopji9dUIUsLrnir4rPUpZiKolxWO7/SHDjZqPrb
nuH95p5TMzA7yC/widAGixPDEHFSchL6/TVaZhfv2BTtSG6e9DCvKAap0Kldzba1
+BY2LE51sNCjpy7XyeLXc0609t9ofV7JMJviRUi7yHThTEAFwZ0E7Z9CI14Oq4xK
15FTzddwhzxpZH5wg7Otu5z3pQ+UhLgoRVGUj1cJihLIcReKYe61UkK3JQV3objt
SnD+x03jZAykwA/XLVjwGWUdXrwskSDSg59WNbsQBk/8VY2LjVkIRaY3l6m0lIQ8
b8bZXibOJUBvdRDn/4pOcwVErGMOHIS8UGCZ5afy78cgYscTXIQIlfbSeAy3p90M
RA4/PZhnEyoHBNXXF3S5ixczHYTjOQ5ZbPJs+IaYeDR0Ju3JjdOJk/N+uh1IOnoz
uPUFIHUKv+nfRTgZoLn8tyQF7j5h8HBRLjaFhgk2qUkIbSzmdiJP8iQhdCKvmI2f
BH+gE8OewAgmE39BlgqEwZ2RpG4GllETXrXjrIX5+MdxCMbsf68SPb9X74BmQ08B
COppn4b7Gnq3z8HwlEX46s2Vlkddn//2tQe68Rodfe3wsGj29JWg5DcP6OK1LaGU
cerRnVGQlnu5E/8ZHs6NRA+zieCBjIVqHQfiP6nC7sbJUMHoAOH8wQgcKYIZXsbd
daFMWg9h/xPhUahAp0i3VfvXal751dZqB5mjfuxlWl6RXQYKr3wqRBxbG6dxL+r1
0Pimy5ZOc4W2RTOHsHIHMFOzXMyUmUCVpCdSQ2xTOcQAIQwGUeY2Nq/iMHV7O9N8
1QyLY0kdZsNSj/NwNlqGQaUUvJAawmAdyjzDCieNQvlMTxaxRvwCpLiXlL98UZ0b
WM4Q43Gjged3QN2gPsOQIOR3hS4+HaUqDPp00H6Pb/Eu/rzSVo0S70zGdx6OxHn5
CacBjp2fQDjzSQvt6uBvVmV9CfzvkW69vWPQsqoWwhvbiRwj46abbNJTjrKyPvz+
YsqG1Wom63Wd+iFVranSlDP7bYrJUFV/SNYjbNXJUqlJoNlUUV6vf9fRjhpThqF/
oWf7wuONEuqbJWej1pyXuG0GSsuT/msMn6/BCFBI9fJgBBFhNzPXZKl8PRNeYS+f
NY8Eh8I9BV6fFTWUSAOi3JZm/sX9RivLpgLYvUkvDmCCLSLtD3HvAvE+/2eUgFsy
SDrDJfj8lOgeXPWerk2yn2AelkhZKXzf3/4P/s4CDSIsJO0eghukZCuHsg3B4JBU
K+9DUgVBScZhqrOQykPEXALkO8OWavZbd70/BX0gKoYDVDoO+1AltAYMTCZEdhta
NWnFbZmjl8NCgRcAT/qssF7s68KJaogn6jzu7/Cz9X4ELqrH7X9LKFSOaihbloB2
+6KObCg6vEA4qwwAjXTXxNpeBp/yJJUgpd3TzFYKsV/4D8HP/tceP5cf1ZQQmnWs
AQsOCak9kwoaJnwo6Q8PvzZ4OTL+9fAfM1w2E2EVWZFiUWIy3GIFgbvuZzwzjteI
moH2PMViudfOvngLDGFg1xRdE6TRKqnk2T3ukO4VxLmFD21/PjHZMTp88pHiQ1nU
JzQvVQ6O7wByebTuBJu2sW0CENkhMrZrgaAYzZACGhszowoSKmbdCRmiGN5hNo6v
X1FlestM4tVdVE8I+Q16MfVpI5tLzEBUI6pxdUuTNRhJLFdrtBO0Luetttn5WqyC
dB1lQ6JDnZ9Q9/uGIpqA9rRFs5HDP/hEBi5PPoCt88owVzfnWRY7Sema5kjf6BLH
rWpex2rvo7NHSQbLutRHpmzJm1NdkrCT/mO/OOd/1ofwImV/7kOZgFv1403XESIQ
kdfJKbhMw5ifxe6npFWvLBToh5Wxvd+gITuKt9nQaFVSyfASDqHtEr90gq6mGOLo
SmB3y54Sdkrlo1HMn0Weh37IkinLA07uAbsmoAGnVRiCg37XVbT2YS9mqXIK0RKt
ZmBZNdcMEPlp7EmR5iZw0gNpH0mjGjAesu01oNU2dwonrsl+zMr2PwEvQfxE6hLJ
MD82Nj8Ap55OunC6CfwP0mVsIwlcNRuYk26s8UTaiIZyVVs8iJ3ZcLsdmj6gsot8
07KjLCXPgfm0wB32oQ4v3Gcc3vPObXRmy1Gw4sBDiLcvZoUjq08dIozLDlSdwND+
2KgNMuLH2OAnMJWWcmHEYUqlb1RQDGSxa8v9teqTT3ucWVxEmSxeYcfgjhGWUB2F
TMdoHb3l9b8jo7Xf1hyDN3cNygBLCDyFrlnz38Xxoj3M/vSbZEmla8cBWJ149Fit
Xf9zJxwWJkuiYptdnySylJxQ1q4Gx2b4O+k7nRog7CBEzyJerAImde5jIuwqSIif
rrXhzPnS7WmGrlaMUHBdVNtJNFNDo04i/ajQ2L/puTWKadYoWO+9CG1ImawXD81J
Ise2rGSCQsXV/Lx1DrD4EI0x5Wjdi6Is1vi00ga3H0jOSKqTBXTMWZPOyFTQn9Vs
QJ1jQCHj/nI0iH0ICEeSSR6AfixJwVDpH5vroFuzb0XENuehtq+vKX+sjQUefNUv
07kmU+Ic713xuMIQVs6TqBdGi254SdOeLQGOWI4L4+H54n7bAxhXQcuVjOHTqPM2
cjPDQb8kzZYLUmoKAjvl8DGBWowIGRluOcsboInKE9mi315cdxm9zCcUAxJP/BCv
doBW/lmgbQc+unowDYTRVcfhJbZRHbqOvpMpvLfoLEi5Zy30ibaoQYMYDJv8S6q8
Mla6P84oMyw1kZCeI6U6beqPm1oB5SZ0ykYBU/+GSHLFyzlBnxjQqDfnph3Tl28q
TJ1qRW0c9Y2mRUU9IJqFVymfiFEzMjHFcHvJahXJ8YGDGjBlhgRf1y4gYbf5pFz4
os15Sofm0Av51FAXLfEluj4Np1bOiXEKDay83L6+dIw1pLUdKgz1GBB5o9uA280F
tjX4hue1XR5TRkcYotxpmmwfrZAUolH0Gup6Qh75HOEc/jkuG/k04PSNfepmbeLq
ba2vHuUoiPr6CSJulzeVW5ePED6DjrT8680tqIEcgya1tPEHNwvSqSLA4U7VMN+d
Beeq2u7wnb3z3WhhiRrXFk2SUaQOGbTCDIA27Pi9O+39ox33N4SkDM6v1fotKIXj
vyGwEKeYXyRfc39oovI10jYyuNXoi95KllQfU80L+N5P4fjveY47nAb03QCA/66D
ovvs1hCY2clno2awBsIa+nuuDF+T4q0JHqC8Lu0WGemZOV0Meb4LoRDWxXhJLGBG
mKS0szMh8fs/epU7XwMWeSxv0yZ+pRnWDEXQbN87ZCUWYV1yaQNHerH3WSCJApm9
NSat/JQlvK0xvPU7sEYi0rHB61pglJvoNdGqTg0JNujLoPYKVesZ435Fe7muowcY
ihcC4vbFMo2ZHY2UGmMm/0RRHH/gvc6t/3x6tC2H91rDIqv3V01oTp4FZEmhmlTS
r0+UGuiX28HrNDN3cx8jW/etuNHjPoO0dhFaVN+jDRLHvwjgXEG43zTC/vlTihUN
G3IbLuiSce/Shkx2e0rf+qZgpH0APr27t0+czC3bYe9A/iqN48opzKEa8JozlVSw
FBFnDpTVXMbZ7CGKe61vi73nmVBcQLJ8Vv3CmStXDunql0IpyM/dIPdkf3eMpl7U
whBAhi29h/K8nha+oIUDgcqV/lbKRpgABucl/xd5zz21Kbl4KbhBVEQbUkQLz3De
jq93v8w/SUZMSv/fMPtHwQi7WLKT7BGhlXCU1lfvWOlYGIoKyeUkzkPiu5RErLt6
Z21pPyRfKvMm7LAnciApb83tXAqvFHYGfIT+B2ubjGwU/RVybJ2n6O9OwU8csfR3
vaeZRQB8Vmt/aO7wx4OmSI+PuWP82UWYE3Gh4RQBpNlu0of/uWKeFBlF6sHCQ1xf
b1Y2LLb3/u+GZ3fZ8zwhBGwlMbf95CgE7GSBX3vVBjM9+UNplqRRx7axHGBGXbnd
8o26UcsHd67i3Cufd246L+C9MWSe9rz6bv/TNe8NouquR+alp4oAwMQkhe6lxfDM
Df0m+tR2qScdf8elfpT29hrOY0BCWdLSUAUE6a0nGB4Fw55VVq5knaTYmqA9aaNg
L0TUUCyvupaWe8FPHvuEkXz3qWYj22JBnh0oDHN2MGOH6IrRAsTNALfb3ACvOOV5
pe9oESt6Chz6ddEmyJojeNqUeX6XvlqXe24k2DSZbTbHMMMMOCDaOe8QnJa5ErxL
uQOMv6o6bpDpLyaauBjOdz4/4u4RZEXtjR0DCNngjNDFgLRs+h68kw3eA20Yq6X9
tfhZyFCnKRVTe+b7gGJskx0pMChZZVWJDrkIhMO6taxeAmqRGEuSvS/R/coLFBeI
pHOdNTCUtpvRwLH8R3rsPnbRNA2bR9LkLnmE04CeT+F1CSNZMP9ok0OOF+eNNzyP
oHD1+T+LkRJD5w/1ZjEJ7FFkcLFA3JoKBh7acqT4olao+nE6hvVHCK4lB+6dLnXn
vfA4cD8Y4LXzeqDC/EG4HB8kijswi2chEJSe7dtD2jGR0lPr4EpElDzSDLkYXDNz
Uf9Rzc+KQONDN64Y95Fp6YuyOMBGU1fU8QxV53grJxPBSPQAZ0h4mUBw0OSupqZB
O81XsvTXqMmVwzfJEG0/ZryrvVuTAIgyZY/FEy15offVN+Mz20YOkSciQWxoVkVw
xSnmrvyofwWTtC0h9dldBQOik636iRjbt4p3f5NwDeXnKohiUJ6+MK788pqfueKS
zLbs5QiWosRb2V/kIbh8dGVJ2/RB5+GsUHxDoqwx5YePWxhnPc6q0Ex87NQAy2sq
91UBcR39FDcD7j6H+LalB87OA2n0SHoHlBJOHFggswXeeFdALr78D58XcGuTsQ0G
LXBTNn2Dx2mjQZl8pEC3ggHtzgyw8BEDOI6VFq8UeTtnIpdxb9+3jDS0BMQ+GJnC
7/2CUmKMS53igExpII+4vYC8FvyN8Va15Lo9TocoMc6FdNsM8X6sNoDhAjZronX6
BmiIa35cj5YP8XuHYeZJ87glmiVNPwoUc+2ihiKYfz0/IH8g8KlTfFfQ/Io3QSzm
9aw/PBbdN50jlFVJGPoWfQ68DN0N8P3H8r0YuLvZ6JxW6/UpkmYJnA3JoNV2R8BK
if1ECH3snmcKZ5NXkLO++NL1Z2unIY62yVvLQsGcNIEHTGDslg5yZeE0eFuIuj2p
2FzGRXYZP36zSSy0CmeaC6MaLBD+3gOW9IDTtfOqHGW0oPxtNVs94BqTYtmCGgHF
IP/veWsN4AJJyf2ZWeP1p8peTY52F2Xj9j7TY0hTWE7fFrr7YoMYIAV4vdH+1JgK
ahJ16fUX+7RIepmKwz9mVSYPRhXCwsVldc6L89CuHIWzNd7R+lSpDbS8XJZHevmy
PDlq8CPtg2tpRyM4CWq+96y2cEiaExImtedeKdoL0aG1n/rPqrXY6RvbitdsSMs8
GEYj1H+ZnWN90M6R15tLAp0f6o4CTlVioFIb7cFEu8fDB98XkVKEcfiWmb2Nr+qu
CKq4ah47zeC0HVwgMBVeSFHu2mm7sDM0p6Q5kvPGWoyRPgpJjn0mikwZGwPqbWAk
xmCi0ZySopYXcyguKEpX9EKgQ/qSL8Phkv1eWmss1JpylnwBRu8dZh4axKL8rlAb
T7mTe10MN6ybM0//9nnQhC2d/O2CcKHmsEQMYCterfVtL76JZ7k4OmNZT/h6UFfI
QwcmM4QmJVCTec9iPGsMAfRe19W/tYNTo0i+KYxjJseIFVASczY/TfiBLNgbQKbP
eTygcM2Qtww7W7eolNmfKuJlIFw05H24ASWDvuPuM2Bx5WHC6ZA+q0GicInldQda
NcC5AVvoAveg0bvisYp+kqA0dRDg8zZKG6vliAOzgFMBFhvoCm+TB7m+i/cEvHGM
86y0b6MScxWiSUE3mFqGKtwGg0Lnti90fvQR8O0dR4lLlqQJUR4GpaeSoMFSCewS
9jdJ4qn9GpASf9h8E1iWFB+bC7l2phFirbr9mQ55rYmwwkWE9nAzYVLsO0/3b4vU
dTIVrX1OI730Kxf6lJ22IJpXguX+GWwpnlOaewnmYhZYEyXdwCvmVJ641FRwbbWS
OHdl/c4VthSVImiaolUr15IU7iMGEnl7Fhl/+vcNfvDaqZg/UIWRONLKTL1fna1O
aDhJdlk6bZC4wrTVINlhP8teZ8GExIE3i9sXq4yPcb9sJgvbxiEb0p07o0Tr6DXy
clC6SVId6BCHZIkuDX8A3XMPwtxPhbEIytq51kaUSJ+Qn/41GPAvqlZm1jYhuxLV
A1qm0y9YXhrvBS2++mFz/rjKPlRTrl+JWbzzodqIEJELdfQEkTCUUJJ94QGtc4T1
VaQpMFqUXKfiuODzCfRyWFJLIZJyCueEvz2rC+BF8dKRTIc2wtvaXWsun5Nnlntl
DzddsZZPwNhUsRCj66NWqBn/SBFgr0q7N0NG4I131nR7YVoy3mWZU+YkYD2Z6GWL
6nxdmqb8dZ/qAXXvt6fLBbpk6eRtozIK4UNTWUhbJCZf7Xc4LsasVlQprv4zC/Wg
tVrBZ7uMT3AC7JAJVdA+8mXRuIWH5Pwgf47Lmf1mygcWAoKbFL6cY3dqr9PIHi2h
ST/3X1ES5jLZ8aMUoOIeUQAGhDGfmFc+BZ7ycqmnUmEuezqPEK1gqj399PZJIPSS
vLTo4tcId1hLJugV2izXNBzGZsV3+1pSr9fA0I8G0lbFTOi6bJihmlrOYzrXmPpu
fdbG10ZmGdZr+PAIH9SwoYIpDHRQfb973yALlHd4R7C8lx5hTOS/nTHy62d+fVUb
2AT1pyGi+zWxIkAGqWrRp4P7Sy3w1qyi8qi6GoRW9GCCuiFB6hP4MBAqQJP7OGqi
sTxhC8w/qdzOSwwUfc+LyNYIT9x5A3AaAxvWy4ypzf4xYP63R/TfuJGXwlnl3n3g
ZVr//ts4Buw0iJYiFQQ5gskQFFlRa12C2efYLwahz5HlAONh2U6a5d+lC1hBnSL8
fh55pOujFoYHLqAXptC0CYCG+w4SdirkOid8n17wRyTRgfspwYBEv7KFNm74xoA0
AMhJT08zTJtm/7+L4U1wkHI5tHr8fS89y3/GdhRGJHLsAanhGgn2vzeXKcTA7hre
EmdQON1WH+j3dYhW6Yr8O+gpEO71m7ghaCBFx7uoMa2ZOTBDdy3YK8iUrcMGNr58
DkrbZmlsZm+e+5+nzYuRzOMdOGB7w7gtR4y8o02s9QVOilVA6ihzWr4TsVIkPTyJ
XirAjwqcJUemVVLHowmW7Z6E7fIf3ENFCwgfp+8sEo1o40wqwoYwOEZrclw9QqfZ
VC1XruoJ8LjgGrhqK5XVjafFumvcLnhJ3jAnTtFwQWuFU83pqWlhMYs0AKNPF5/J
kt3OQtu3VQ6jAslci91fGVmiiC4rG4M2nZKaLrsIrJ9UeN6yyvigDrGdNnofwqn2
1HbNP7gpdTX+oqjeB3ARlmA2at1IriJN/GEYEngEmbGM5qP938zIV/LUKXQ9uP9r
w1uRGsb+zBXWEmt76bOrhZNyoNcmJe26Te/LaGaFfqKdysHxkkRRYVqVff9073GB
adIAhAaPQTQdg2RfexW12iTfBCWqS4Hlqw4WqQ42dAAUjc/WqB/n6d1BHjWnm50o
UeHAu6Jedj9cwxUGbfvTjTnBQYAOwCN8+a4bPjzKBbj0xjc59C+th+nxl29JRbqY
Dzp272n0x8qaN65DFt0SsV+p800CxmXT+MZ/C7nAhX9wZn+9LLj1ICpT+fRfO/Hc
uzUWKRcEcu+p3fjR+nvSQx5cccNJ14xhhbJS0zsJBPZ+AiphuJ5rLPt5NXCOqHib
zMeTyMNGkoRtG82yjgzPF+GI6TtYMZn0Fvo7k84AljqCFVH58ENmwxhO2kJrBeuL
34J+yemDPBW4XO0B64BXxC3SrPezh2LcEcWPT7gwmRBUhGKKy62QXdHhSiaAPjZV
sbyTAccxs1U69dmVBs9/F4bWpiQltVMbxpizzob9lwZL6L+9RTTvWzY8sUrxRi0E
KZAxn13YLaZAWELzN2+qt1SyxC3TchkgZqvqn8ArTZOX9Jfr1OQlTpvDzb7fu9Ue
npWXVslDNK+euH/wG/v9s5UvZ5eY9J/tqjgxkc68YoVZ5AvLIVSnBM6h42Xl5luD
q0w1enwTTCGlEWvAAuJ8g4Gj3Li+IcVIpOuzRBmTEPpm+tnBDjNjV2lGxrzvTkLN
6jS5Sx3OK6BCtTS8SwOPtDoqdZHcOUP1mzgmVlLxZaXDYc3sbTEy+5dhLZtQxxZY
XfKA2YrxKzq6xWi/GDPcOIzNYDVgjHFR9EN0Hu9WVh2zBNbHxwK1U9M0WKuU8Vor
zF6YgtPgCRc3dQrFLTqePCqprTFNi191F2XX2fQdsxBYGNAk34Q1KY19qkgAIOD4
Z5yDZlQ2jBAPNPVU3nKDzREOqfbVmYbHNYQHWnpB7CPCjawg3LJeV56vrGUP0Nv3
AIjBPvpWpQ4x54OEA7H0HGPrs46RvaARy142kyokkAT2j6K1JmT8cxt2nUo7/Juy
G9CxoKmm9hcBXhXdGvVpIk+Qm5hVg4VdKaUI0x1LdCbg4OlIPokFeQiEE6F+PYXM
Hdo2+fF7j9Ep5BJszb4EzWYIr2HVKfWugGZf497FCb9FfRI3D6zy8caKu8smY74d
uL//js0PlThmz+1S7BK7vSMi+2XxabVy6dS+90fpz8DIbwommqFnEn32JE53SviY
JBUhHKo67sVhgPFKa84n+DpS0M15bQEoHirIJcfghmo9z7ioPqRZ8vkTNTOBeWhB
MOkg+ghu8m3wScWCLcxCg+pzsCeI9D6g1j3+qDr+wTl+vwv8JhoJl07ilh7qfYXj
IkLe/AJEGe6A9s/vPpfN4xBseMqip3zdP14K7+gjJwME9XjFQQLNEOw9v23Hgoq8
vWv6ofdaX1aXL2n4UMcZHoJf1ka7HNic96hw/K1keAg63aZom4y4QZduUv9FPKg9
nbmiZ+UAL2Cqwp3h6MxMB1Nbs2H1tORI/y4KFDJ1wGGQ8TVG6yI36M7YPetyXceD
FM0Shsj3wfjG/QkDJ0xgHofgm9pZM+rS1VoQIGuL6U52VnY7eQBh9HQartUhzuCB
gTZwQ4+N1wcGTWj5kigERYrJHn6kcRRXcbtalIuQFGUpn8rKdg0OCpuQavUA0EnU
W9ogpcVZWmhyBZ/AlJAdaUaaDBL0DAcxF5GCSfWe4bawcoW3A6JX8sx5cDF+Mfqn
lmpYQdaRMNA8oweoX+Y+L9xdcdxBUw4pcrjAzem0/bZG4XUpIQEpIhUZoNKeCdAd
w0hssdl89v/rhjSG0qLdg4qbZBhWeQx1mK7523PwCXqtkkmBmgTwPTTofLVubgAv
ueaMTNp3dJtC+AdVKlIAts+yEyeVBWnvrQEaoHHPaKomGJG2u5MIFVHCm2NXjGdq
FlKkWSn4UbU8q+ar2x+FENMX6qOmToNi+5k70KhNL5FFupCQWlH++EgV2ulAdGNm
onc3dU90Sa5+OEClkmERkf765mTMfQJkkbVtbwQ6sptjU/15dAwUew8HW1z1DrBd
mN262MRh2sAalhjgSQQy7FsoaFcjikmdghGxqhau4zW6hOp4DVJfYmbtR3zjLYGs
TOwCVwQ00R8rAkKfWSl8ISSUukkjTTuK7BrFhB4tq8Ydn2cqjJF4F/N0Mto2PWoG
pmG/sQ+q+ygNK2oBOZKVoXLA2gxpwuh6qD6Ofr4y0LMuwgXtthZjH0YOBA/cTjl0
qW320Hb+n3TXYATOvygV2pakkk9t52uJGgJA/SYRAVRa/pOAwDqdtIsmSWvi7tEh
F8cItX4l4uHfX5u/mepJIXmlwVug2DRBRkFJIUToDFRpC1jX/JGtuFVUGchUmCjA
MMPrCiSepEbXRyGEu6cu1mpJZmDGz1qneCfLA+A0AprCH9yDO0Fb6+b3uJQFnIuH
2yb6JvfBEAOh8dbJpvsguJ845V8uR3tqPw4LAgcq0vvoVlyERALE1oXiQJzXX62a
YshTfWUSZ2JkuNnlqj2c3iRD7UdI9LQ7W9evcf1sdnl3zpIJMzN75Sr7J19pAj31
vvtEMyPsbAfR7elbjzwWv0DsZ0vEFpXHvL7POrrW5BJkuxQwU6jA5iGO1CpPI6R7
bk5UG2NnGehcTW1tR/ML6CD0BB2iZSnk8jE+tIoFKGl1y3BvrXaQA1G40Y9VYC1E
uS/0dlb7azQglKU18kSKUaiKXYu6N921nt4X556sSyuPHVZAWwy04ppRmLbtaWZS
8Mlbz+CKDAgHvLuGpR/+QG6dbqIgp3ghJDi3HG+35yVtCzUi7nhhZqpRclGh8d8X
4jdWhhIYO1uubsDTnI2bKbVQlG6eINTsi6wM4APtpx5lekmkxz0AC52+PM5j3BIU
JZlc85Mrjbh8t4BYH8llI5QpIYNQY5TDPxsZ2HS6SjIS8pOw4Kacse2ql5JcWUPj
8loyYvCjfbX7UxTJCQ5sAErSNmCveaeI3qN7QjnTzTAw9jC1X0OyVp1CBBLzDfnX
GqU4uv4G3j7gMrMm14LVK+lOjN2asUGDAG4e8vyKICRYL4ICj5eU9Ow0/IMxOkqx
BJNsjDBfEgkDLlfN2G0fbO6snoHE9hQEJAuzighL/VDTkBFrpQOE6qi6Wl/WFx/Q
ejaVyvXmGZZolch6prBYLQxt6/VYjITHbP9R1yW59atLl/jBYnbI+caW/V+pCYUv
CD+K/lrS0WgE5V35AzKGhgfckdqhO2haVDmku08Z3+bQDbvxr//49Cly7GtsCvFp
0pQALTvXknGOWKHQvsyPFSIg9m0Eq4cMNu1i6RY+f2ccGz1aBHOlSCCfE1ohlSvk
qRz220Teep145jz3mZ75KURmOHig5xftpC/ugTQz/uZ2drCkw5u49Df2WPyi/pTe
DhnPunI8eeWEQeL7uVB9/2vkZPWyA8LLpRy7IlvhabjXVcfX47DUXLdN9VzZgceC
6hR14bF8AtQWl6i9diak9PxVVul27fAF0x+kKTXA7UqMZKjyDhxaAmiaALdbOGMD
GcEfRL5JJxOUgOjVUiE/1LA8GZgm7SKKK7fJLfpqQxtrPM2L9DnchcIcaFm00K5c
+VwxZKnUDcOSFhhw3K54cWgj1UPcUZZOcaQHxuZuTprpEEfmZ4xxsAC0071VvNe0
GDAMSwt811VNxZ9Hw/9MqKSVpRUuzL9l0ywQmfwn16ijxkULQoQxkza9oLO1VGPo
DQIyTntcAW7RyhvLyO7R4K9qY0hd9aL/yZkAPXeMrEvBxaUiuawRR3+hU1mQkd8B
hJBhmJEV30BTOe5ucOiVF5ENXAoBBrmdClgVCq+DcerxxolvQ/WepwUA/O6c83ZJ
QskQJuabHOmeEnnoABJNecMS6kBz9bhJiQ3GYzGObSUkO72bbgVSsTxUbIs8GlZA
fHvWDx67jV3izVllyhKJdSoC6ArVukOreC/h4pKnsVzSxgW7v79RKVH8p7b4SoM2
h95DdUqZM2HkrFkSMzZdlqNF6ngpdonz6SxOVw2e2i+tZ568oVEZFrlYO6ZrO4zO
1KuNJm3RowwUcWjgRROfCpQkFsUCJ93BdflI4gUrEMIspLKiFjvrY+LDWH9raPb/
k2So39FdMGdABMbrBRQIzEWp0XGBnp1HNnk1+50pbQSylRINIcI5S2RAVXtpx7dn
WGEmrX2b0aiKxYknnvNiVLsx/3jMqfZoaHrAEAFP0D3QhjTy06ipA+PcoJMgsRGP
Qc5uWdRfFA/p+lpDODB5tj3VIX4ROTT7yN0Gbc6SyzSmIfQNLoqzeqZeha9qkmkp
aCpEJhWA7LwVA37ySZwSIXhZGN4uXxyvzifu6949Lfx2h1fkDdRdhXoXjK3yzDaC
eInMbHzRNkM6uw/lHPo5MNF4AmJekgdwrRciOgPMOKIU6kDxmI7+DSnw4eaAf08Y
HSBe9kSktcyV+8fDQ0XZcDDGhmy7JRp0ffaipKe+OlhQ3cb8V04KseCPLxB5fk+O
eTlRWrk00xJs/2c/xdQst5RkqlgtqFO2aEqPPvFcBw/e4BN2Br0/FEtGYia7wZ7J
Z72PO4wtRnVFqAnkwFvrm90tT8q918OUlgs3ijHcwV++O6DS2qeJXqUGD9t3P/xH
d6qUSEHLkD0bFVpGHFLLddgO8L4HtXsarQEH9jXVslLqHI6n1kBSkPxyG1MhIscA
HY2nsh8taYC5+Ij0FgGxWOVUu9iC1Yn9t8Eh57xtrKWwfOb1Z5I7Tahy6cO/cCNi
iV1cFwixwtvQE5OlqhZeLd/jPsjTeHSTQpFjyTq9JVqHC7m5pUWNP0qvOyDDelPM
UW20j9b4SNgHOAQayHur+CXUFYZHYd/bqVMv6dklkZsp2a7S+1fn5VrDi7RlX9TJ
tFUE1pHdthPyuFZLsn8fxJRbXUIbGWbCELShxRXSRssheXh5Swqy7IrJfoxLX2rT
X5EvrhjukiBi0Ytoi0vHiGqG9yWKUkpec2XZfDu/jHojxiwm0pzBW3DItCA2SBDU
lDq3oH3YgrjR1M5Ljl9HwaADa/ojE0nWTTolmcQgWuKVGJkCZ0DBEapYAfsntrB0
pbrfqQOq6Tu24PiwtZwNE4iYNTkpEGyRL7aQcWAzvuEQbFvEhg/1x89ze6hikdHp
pEh9L2IK59sPmaHkm7dPo+fuxvFpDSQxvHHjGR3bjWX0JPJTkUPoNJBw43NVxCf4
omXb/Re3M8+N3/2UQmk7+ruaSY7RATsCLh3Ciw7lOXsb3qAzm/Fol39LRPPQR0IZ
RQOcr85usoFUZa8ykTgdghDgAp0h2vG2uJGDqnCINkY9rJST4KlztNjEss9k/jGE
vqB48fjPyvwuF8eEV0L2ex22fsQKROkpUxgUFackhR6JjteSSs6va41n+/Q/JR7/
E25vqlwlTZVXp0QZRbDMYN97OASMOS/r5xcNg6I9oQay7jpfwmYXd2cEZeEYNE+w
Ik1to4PCYNBfNE/guFikwGrwfpYK6CDdXNEuzeSkR8/IOP0vgvYI6g3iSzjvPIi6
qdW1nCfA9AN/VBli77Wx3gMpyl5Tc5vvXJp1YKUBigR1x31WlZVU+pHCRuYPRVa2
wQ5qyMPUuoH1v+3ZYHTQxvE1w0cwWf+lvMLBUrMkF3dEX9ilnrJUXRvCp4mF6bry
/ILvxE7WoKGDAtYqOVgdEMWJe+icL2xtCISPLch8heGrYm4TtoQwIHuuMie2989S
z780KS5i6Cg/Ry2gAFXQ2EjV/h7Yvx9vFxa3RSR12Q4lAeYmg7wHNRswsryhU9G4
YkEpAa0Z2ORwLL3wI20q/koRZ4W4ejUvjBS+WO8vTbZFyi45asBNQpyuGyO+iCBm
v8msn7gQ3YOfA6/5tonydqGdw6eIyzTdPxP40i/Ci2w0FdH+YZanySeuxQhMWTKV
8Y2zA8nprQL9YakEsYvnB+V7gN225cwhijMXgTQdBIO94eUMavbgg0xEO9DqCknx
wrtui6moLYkZHP91/1QlvlRurbDqVmQJtSWPyk5sGm+ygKGVbGUi1sfuLRCe0haK
/jmte4DyFARzywI52bam/Z9N/rGzjC932y1e6g6s4QNh7IN5EICVkJeBl36JfveO
984F9+Tdd/eP+y1NSxzBVfuHmRWqWK0lBT7tzCOVx76HPNwdNoN+xrwapfE3tNSR
txeIDIMBCGurZ/HCoNm3X6Ux4cCUVP+8qacOIhDjaEsUr16wruAJK+oqBTypTpIH
kwAVd841x1UQLnZTMfIWzOLy7W22Yzj0nTyNCbhtrGgbsJpJRUGZwMFBf6oQPsu+
QbuHew1GRWRB2TOOGz76ZEQCg58kWDV6ZkbFPnkgbvX1LSIPYIaWJh2LHTVXrxqF
NwEi7EcvN3jOY6LyyIjxelUCgxyB1vppJnh+L8vHgsaBPXsBLndj2Ys2ITXHJ2L7
ObdLSBUM6OhjD+02EXvboorPqiKGdQX3vdcBC28ZWjP4LAaqiraBioTbgAenI8Br
xGtHfLc9YAskqHfXjfMnhAudL71QBXkf0qF77giXpSUrQE6cJDjdMtSye+TExctP
Trz8NBEVV0JG/gspUxgfxNZOne3bfD51uFxl0pf0Zq5GsBfBFrhnmG+Ay13Yqajz
SkYqRpODIwZ2aaKk2YKbu8H2b1F6JG7gpYFPy4Dog0yHdbcMEuT8qsZzwFSdU6Cp
eYN+zisMR7duqsbaNfZCBrjhqM/Wq9mnDpTG4076fmzreNRdjyvcSHVYyFvtgbrb
pwz+eYKYyFDd0NH1fy3b5GFQ+Y1Fam2kzjXZ83JU7eDrCnEicRu8nOnUCC1Cxmv+
kvopAjsGo3jeH7iW7UK3NTacaLhXM5Tvp4HeKbfejFgajIbtQVQiOtv5FWNspsgw
smGFj3HW6yiIWHlqlEcyXg2Wf4Jv0JG0FnUXPk+etcQxaOsZ08PjA6Yvs+sM5r8o
CYmLivSTKkipERB7TqElwfJNxo62WQ9Dq9uAN+ierGb2lDzCtc6H4U75eCTEzlTB
IP02xZ9XltXbr1CYaKKdp7sD+kpuGfyCklrmbDJOeNH1vufpSfdTNQrepn1x22RB
doWetljQ6hYVbkDOUxj+H3ezE66BAgVhGr4AwDK6IsubJoYXJDVnB36FY10WxoSr
L6ynmlU9VfjXF/Rw1XyIrgRTDWbI+nDfohPJKXCw9W69w8h+IVMXQ90qoNyHxcmr
toPItbpCoxTUezHMOj45/vycgkTUUctFWkB2Z0eXYoHyqzK8222cnqbsT4jERGCR
4Hrny803ba2uvQVpJ/ceYqVlvSBD6zQFPlrik5WeeJqVsIpJ+73tXzcesdmbgNEK
6/7Kb8FK+FbXSmGZrKbC/255uZmJ2sJJyAhMEwhbILr+ZjeASWfSk6N5LLptftxS
CKoXbYgkCDSa+lhd+ZgM5hOOvd6ExnPmIwQtucJBdelkpbqYGGNrfCtKXjiqukkP
vP5Xb4zLTJOT7RGWm17eFgOEukl3Ffw3WMeEVG8z9zVUCdmNM7bS+V4vhWuoWkai
00IrUjrzwsPJ5/pd1tt+OsYDePoZy8I+8UbDRkACa/KecvsG7atOwij6Y7Z00gPI
5cCLV9EljWxRCDFZR4ljA7HRmRPk5GrCiFdtwYtaB46BdsCeWYwqlN5nDuWy387e
yWDLFUMQUM+sSAkXHXazwqpBc+dAHmxrgWujgOqqlEDCy6GxNKdPDIumTSFdqWRF
ndUkujis/Nhe+oK6qBOqrAFtktvg2I+azWpvuqDJTJeHmGIRF/MhvmUoo9RYnFPk
6Y4m2/lYukL650Kngmwte4EvC1usUrNQNGUoWEyHP+ODBaa1fvWeFEGCuwcG2P40
YDrFx9VZwR2FsbgFYEPwkCfIMIIuWWC3nB7LhpQGNgWY0RXKYgV4K8XC7JjXUYmT
203XPzDG3jja2FPDEuUV9YfvDZVpAEam+F3G669QNni9rukFljKH9y7bwcctTtDG
VAUMrc3yRKvS4bXiNMPwpil38d3F2msBpHbvJZ3OK1a2U/EM65BBOWR4c73tsZNQ
Da3upi8UjrKlt8myAA3lekBTO3komLyYP3XrVcqoRJAq36n8uyMBB9Qtn7pCwrnk
8eecbrF7rkh0AnMlnGaG6cIgXHXEOEm2tM13batitR5VsVj1EP4Od850ZNg8VB+f
VUZVChrTocAsbFJT32YIgG2Aq5mOpYyg0Wuq2q6gFoqv3mpZqh2ithbc48pT+y4n
GyobuQQ3Lvyte+9XD4mJ+3/H+5ayNLv9+okPGLUf308ffjLLSfXHn9LFa2R4xGJ3
WKF4MUWMuUpEU6QdRvBMcWjh4yS/X3zp7uLM47zXF8UTGsFGCTuGCtRJWAYYM6Jq
63UPfvgDp5wPyinCtTy8qJiX75YB8pz8m7ZI1vxecE0+5tghWG+tPV1E1vmLpTsh
dN3h+gznu6fTAAiRaWHJw9L7aes4yFKr30tW95KcPnamZsFPdEinUmZWZt3QuAn2
hoTDbXCxDAvXda5OySwb9P2gJKuBM2V7dGLPjwbafqg2CyyIE0ae1aZDVJO95E7d
opTEoOf/p18HvMgEXxK6SopmzQDXc8IH83p8CxH9jMwbL8JljUI0KtOVgruDXzKU
65LuuH9mfQ3CK+5E532AewvL1V7vGkxCz+NMBZ8LZkNYfHqeD7lveWh/R6K3lV4S
E9sFAhtQWxE3R1hkDo6srPnC2Rh1nnfxhDs5odiqnlH2/O57D+8W7OzlZaCC/aBG
QldaQI27Viia9mYuft2lSqlP+pZuswSlI8qMcvOlaVA1AtfWFmlXehys8t4n/sru
qdCRItkqyc7YW6babe80iU9Z/rB9Uk0dRlbkY+stwKyLgJ1ulcPAAjLclgzHSItf
nonK7X6f7pM1K+OjHJpC/ODMR43QltZ5IZtj9qlp7cRMaEK3t4kZTcBfK6F/hEHf
xn4HQiemQP/OkPkzvYDStew5PLrNOZqI6j0e8xvjaggaUuh7dCzP80O8O6xA4aJc
+MikkHQRoY2izqlBaMcBQZGfxIblVudSwSBytSjGPt7UimbWMghw222v2VzeCZgF
Sf0iUikz07aMmXUruxZheEbGc621SN1OkER++AwHgD+r7nW+eHWvHz8BJZxHJ9Ol
J3R9fMZWnLo+Bw2OghHwnF75JzFl7ZczYvY2Rx+c3a4iw6w8HHcHz29cFciy725n
LjwUJLnKYvAxbycPuc37CFFKKyyMTI0TEsqv1GPssuBD9/CRZMfNiIwdUvtA1yVu
2Sad6nK+U/h3PbcOefjIvxrvaI2u3jRAw0nrf9t/dgqws/PhXpPJhx3k8R0jqO0B
kCXSMiBs2B3Z2vu6OoMaBZF2lrimzDIowZajS4WhEOL8vkgwVDKr+TuUUGbCMPK1
PZQsH84q6fOl+7MUcApsMkYWH7sOjec9wONQaLC5voaI/k6qiuMgLfAFwPHVQv4a
Vy/7TUhHlVk+pQdzunLEZ67Fx7rtEltMV89qJhxC7zVodBjlPkhEsIHermtFgILf
efEZ8seGuowq/gdObhW30ZrlkvnkkgZenJPTz7fRRXA5p6R9QZvdjacNX5f6HdW6
n7j20ChBZ3HP6mFbyEwgO5bHSFJSpB+MZRwlGi/vF3lx1j8R/qyX+x5vDV8xeKBF
qFy+XM7ArMaWgH8ahsLi/4kfIo+4ZHOIgEQPhCPoFSJ7Z3OqrKdAenvJiNuwvVa/
2ZcUjTwq60qyAGWcJnFeFMEJUGj1JGfRUFZcl/9xU9pkT6qB52j2OSrYp8ENcRHc
GWXx3OlvMQ3nd0/KCVoXrMD29oeiBZWkLYPb5ezbaQ87xGlkbIjxtU5cyEkNSKZT
3cORM1l1kHJZ0wIWla1WsE2lK6mjnHeS6sxJQn76FGKQdkStuAlbig4i7nm7dEli
Yfo1WyNQdmMY1xrNFPbfNn0g9Ktfo4SyXo1Xikv/pa209Bd8JKixPHPyJc4BWkAW
50WZFGKyt0h3P/g5U4sF3H7uSqE/E3jj7JHDc3wtuTOjXFx+VVmzc8lkHVO7cDy3
J3rUg4LG4kgwluGg+zUkTgwqQOy73JXfJZu+wVET038ixI1OAPWdURYHyQI5nStr
eHZS91g8pOWTJYeu1+EAx4P+Lm9JJ1cZ6mNjdBPnpQXxJsqqFT55FRvbjruGCwV1
IEmWvqu87YeJeCNtHYzwoP0D4eSyG1NMaY75AofSThoj+9CBf7ldS+BdnurtguvB
erV+/Itr/SwSQxmC9fR7zmzM7Hylb0k6z5ZbwZlKpoyI0RgUr1tMhvcrSOVOrlXz
bMzdL8+6QEx0QfU50WL5NXLAKrZuiRLYFhFDBisPpT1g1pGvOOxHVZUXpuPqP3kC
w/7GjqitCHHcqmfSR5hIKyTdtOMXdNHRhvv5Kg8jFEW2zMUBxZ/dRQruwGg5idyc
xlmXjFUBaFMKNNvKCUoZ8EbscRi2CD6KhpNQAfCxv1N2G5pcPkSMKsWnH8TUpXKZ
+KfmwG6C2r4xIs7Wjs8h8UVyIZzn2/STF1M2vUkevWzyYZc24GJIi1hvYv0Ro7Jc
mPuAOzx8t/1mWn6kAwtGNDuX6zOgtUPlo/E3KqlJbWQLRECehzp6ZgBtNger/OnG
GwgV3th3q6KhhgVzv18wwqA5or6hDq/QCLMyMCOeNuBnYuNKjKPtl18M/K5zTLBg
eM0xazX9yFAij7SbY3l3/o0OTYY2y2ygcCa4frTUUBRnRR7EggzmvzXczTBomnCb
SeJ0gh44jTa4sHt0u1rN6ft1+6czlS7XDiicvsi73kCET7VrFOapM/5FUEJn6CKF
cFCY2unNYSoAXDMlE15mP5XgxosLZ6HX1J5R4FD4Z1+uuOM80pZWVlw/gCJnAaaX
ziOEEuEo6Z9xKBriY3ar6arz0fBWvHINahBxmQOsnraoIte+pT3weQoiEISJF1k/
h3lOgJK7M0jtFim4avuiXIqs1qhmGdmx+ghw6YjtWTMD++D9bmPB96mZdkV2s6z8
hg9cC3vrf8qsXhARg2wTXEHg2BvZkg8ofEtxC/wWgO2K2v1yTQtEfb0oGhY6GruT
jQ3UnfCycViCUsxGHqXRTqvr1NbcW3Z4DgMl4dYq0cpg3KQPdStHHnXhRgyuGO+6
0NCchdxFCQrE7NSUenK2uonK5pmyxxKTxXpBWqCK/SP5HJ6WC4HT+obs/YNjSzKt
NZ9LzQfzJCs5WBSjGNWN6s2U2lH5aS0fBB6BdtxrIEsgn2pm3QYUBW4xXKM0XLvE
hZqgBg3H3v41l0LBicSJcRNCWm6CAavXzZ7Xj99DKfP0V/D9RzNLt9JhE619uHZN
4eUK1nnNgpLwilzAjoun5u+v7JjZmE3HE8ujoOBwsdVq0XKIy0r68PID+AnKfjBq
N0teBhOl4zpw/xtZbeH9OOAC7iuedr/Kdi+MFAYlrjm49GKrTzB942AjCp0/BwPX
3Kqc3bpz4ik4bRGx4IWohI1CsLejhJg9j1QKlhtVwnI0c7lKNH7YWNdOnOT4wpxy
LAaZt9gLGwIZ0lmQ/eF3M1rxt0eGAPCt4O9WFF9Fkykh6S63AAdnpjfXctCzwCzK
4L5FAFvrnQOoo1sR8iczUic+BGhifsWQpTa80iKzNH4A0UzJkfw90ei7azg6aSLS
kkqOS0NuurJdBey1j7Bjy2++vPpNKaekQomqQTyLTQwelnZgw2AJPgX9+QaNjmMb
uMu7rLZotmcv0+pyZVuk+q+tSARppDthX53Pf2WnThVV5pV0WntZcm6fO62SrzOc
xQ3AUZJej+lZqv9YAjz3HWt4n+tuLHATeBj9/ZdFqV+WYVIt3IAp6LZBQYelbIc7
AQpE+Yng74dbPgyW4KAByOBs2MDCV1LrXs8TV6q8yVltJoVeI7oBBWC8js2F1yef
Aj2KuItS6paDlByCeq8NSE17oMWOkW1jbQE6xqr+0RxKjg7X5lOpB2WBerUXQ3VR
2ocb4/QYndflOt2SkESrSUT2y8eHFekb+gLHEiLxs6voQft0h4Pd1JuHHYoxMJRJ
uHXthAweu7TZ3pzA7vft2L95HZNMdhaHPWrjPP4ITpgN6cbRHmbqc0zpn2EffLmY
rJ9ckZ/WkEX5R0YXiBl0TjFNDzEeyUIq/fqT7TzbbIQ5uvUHdWOd4Mg2OEpZWGOi
kOAdcubH4hrvr0lEyMQvngOq0ivkhYOq0ILfEGPjOzkKO6qg8sX9DR2xXZR4ownE
KHGlF/HbfGQ/FRnReLvrIMmrtyof2sZJaw+fx4q8WGNwPWP/eLo4/ttwxQdvyd5H
CWq8SUCBW6s67BcKveaxYkk5Q+p/d/hk3QUf7/NC8DtGDXAMRG3df3q9b+PgIVLA
XJBgzAqd0MQ7XQwfXL60a0ZzlzFAQhCHN9PWiVIfUJCO15V2FU1alWOJhTL9TML/
rTSS0JtDnrldSTwSnTV5ur5oQhxVyaR+zziqN3xua1ep/opADUaJXtm878mmsm/u
s8n0qSez9sadTgIux5nsoqFBbrGbf59v8BtJo8/iUPsI9nig06rWsCqnFWRN6T2P
wrMuvrI5DyINE8YIeqpBtAU52sIiCtp2uIWovMH2JcgQ91jvrtRtnW2kno2KnoyZ
KyIqoMnokH1WyWQt40i4EpD1LlnMQXo7sPJXK6g/btTkfsQsDdnpFJoHjEttdzAt
xqma4CBj+aCO6p9Qqhh2TeJ/jjyNcdn1DPkUxXg0ng0AnDMiSlzTQoZp06+A3END
0z/ZNa+3TOR5R3aUrxptYLBsquc1PpGVosHJ8sCUga4+Gr4dK5LU1StRZ0b86WZy
g7aoJwGOoX78H0t+fic/5naJrayCNc3Iam4gXDQW80B1VLTVnm1CEbNbmtspTl7P
JP7E6VS217Yw2iFzAbuvmixYni1WpqNu6COMWmGaE+lx7ObIaDcV0Qj9FsiR8KEY
WIycouoGAKMh+rLDGrWnNy5QpTqxP0cV65eUkavyd+MF6wJln57O3AMA4qWOaq5v
+cvePrkMHUeeJj6sVRS3ZhKe3UmtgagXch+kvwKZBKHfbkH55RMOJjDoGt96/N6S
KQtA4SQClUIkE+RTYhQqwUcet/baWorQbH+G4fcJ5NyzWkeTrWGETjgpu04xJirP
UdqhgH8r8njBFLkjkrUErhyZzjPbrmwmF4qacfM+jGSehChlawwBQx1DbKhwT2te
dTAbwnOy0BKVqp1icKRkkbmO0nNufJ4aBUvO+RzCTXjGVrh3thEFu19kFi+EYKNm
laOkhGMkZI+XgiWT9UVFjRplTT/qnHe9mMobWGhMH6+ES5ZIPIflFMOQc36mIaIJ
Bb5RymULrhPRyeRJwZIL9gnouGbml8KYId6mPbjS7izCKpMskUl5WH0+twd1bRF7
YHqbY/Hr9Ggy7lP7C/3xgzp+DzJ9oBwsfNbXD/+itpDfInIXVfpVWa2rfBYjVjbR
k4YSUE0A8J1XZZDvf9ek+hYMLqyfm0NZqSaxPFH4KYdSuddK1uEmmKVgRm3NVWYO
TFJNqDl58GKSho/CRvofqTyJRleyAOy6BWv0CqIJh77tu5VHsAsFNQJFLBeX2I7b
FtVktdVDYEqDl0+rg6JYsq3+VrPX0i+Uz8monKwMa0l3P7J9N6jIKaSKsxM0J5j8
WdPtpspnkoN5GPv8sgo21r2IuJfwhoLjFIo6SXxbQ0Z2FlSzwf2WnCzkFv1xG0+x
O9CCSpk79T8rkinQqIqKmb8H5PCVE75nSt2u2JetzzvSl+IbAdrUfRSuiK95sG/w
3/W8JCqR1/cQtx25juxGHLzSwpKUezJ/l1TJyb8EXdFjtIV8F4+0xkjcgPAAaFTM
rBgNTTuVDQIzQcvRyydGMLgrIrwf4RqLgBqzeSepiXHSCnJiu6OLm6mqvlMLiv5Y
YPK7ZSlFn6n+ViDn2PTrLqeQVsCvD5Mw8NqzIc0agLW/h61H9xCtOdGexCStCwpb
sOcT1ayt/nilJx4yVLl6+taxwgKdv//ntQwCOHAxwXIHPteR08i14b3G0xHtWTyz
u74JRSeIxJvtSnful5ar8gcaZEaY0yUWux25RBTWg1/8wgqrRe6bCm0TXZwZJTdQ
SIEKUfnE76Vr91bLbY1RlXaCxBsSA5tUpOyGW3fgjlRPEC2E8z7WKaThiLPFj1rt
15Zbw12FA9JXOn0kvNomaAy/YlkXgkTPB34z6bhxT9EAc1hqSe5vr6QE8laDCjkq
KnUaVDFHFXFmWpis4mSb957BuFupyZbNCByB/3CO/0UZz55RYHvAEmi83v9TQKnu
hOzHu2nd0b0JlVnThjnCgnVX+e5N0kHGroQRpmdigr2LlZ+hxTIlP50MAx+1uY/A
LT/6u8+s6EoOfwgVxN2/GDlpBBpMJnVl5/rAJbsCcWrfOaoDKKx0JOeu6d9wXAXr
hULxQcau5Gvnd3iXNGf5kDjQJWHZGs2it/jc2Xc+5hjFaRdW4rLxVre0MOzlsvRh
D3MfRC1OaRSEHYjk4Y3muJDbkF05qN5fWy8+Iij9BNAaY0EuC8OxcN6KlRYrqfcK
gc4GFXQTgaHDI7CP3ORSOrS/1GK4zWsAGODEZ2oTLpQWsYUXJLevuMm4WO3IDkCq
f8NvCX7YvM/GYfg4LPApFdX9Grsdm8Voe4ugTRAak2qCJjFd/gmde6Y4p6m2TPm2
NYryOHFtpWCx5SDHOC3dy0jcOURVXKF/Y1rV596aMmM8rNDsr5ErzAsy2v7dnvkG
GMpbL2fk70d4rg0x4LR6TEajfCluA8LceZWli7KOj8sruTzVTTiB9Wq7ooPo4FIr
9GniS2/zzQbS97EnYi97iLUfnStJZO/QxFzynnwZ1MgtVYuOxGte7Saw5g9UDjZG
FT1VYCQ5WnQalJyURznoWcMOUlnS7njEznQ3YmHUq/r4IA6FWNeS3elhuN+VfxZq
pE2oQyk7Z95vPqlFmuIqJE9HNyZDvFkx0Z0xRBWEJNAjwiIaYqhE0QPrWSHqIZvb
hV3nnBhsIFu9Sq8yvDhTnxnZqARrNh+8zN0t7sPxyBfExuGqm7FjOtS+35E2x3RV
NO71TlcINuJvD8E+OmQfWLpdNTlxa5w9IkKUDW2SBsAkTbrLodnLiIwYdwm7IJpG
CqbUlRRvkHXIj15HxUWdAOpJnxDYCfPiwKKZqO0WgkUXm/in+1cXYOeY7MpFCehy
AOT+5srFurDca1MX/W0gRKYqr9izKLR2DfnfE6pl1VYvBC6TF5hhgACkCPITl404
IzyGmJA1KrsLmYmQ7V27k52I3r/yqro6Xxz9HO0X4AX8tWgckZFLULZZ1mOIOesD
gf7Lu1haQiwTkIczx/OePfkb8QMbDrCYzKSTsdhFL0IlPSkcpEgyG7gEjL1fmpVY
CM9urBY0olh0SwdOUik6e3+U5lgdKkdng6lIICPcdWDSA6ubspvhhOFKh5q3Nh0/
192qCMzR5UJJdT2DpFGfMcFAJ3VYPy9dLdfqYK1HZx+1BoEbD/8AaRduHO2FdNY7
EnrM0wcoKYNmJwzCyAaxWzhGjgW9S5sFpWea7Mt9Ti6OCBY56yoqoAEksoO+Ah03
cE2b9nJ3tqpSGBYZhWXEsOIUn+nVHTvSY24Isc9E3HlgBmJv91lwOUs0Z8BEJvUm
1cSP6HIdGWyqiZ86OpwrAuvOoHunJ+ANtdLGHkaHj1TBZQbr3R5KH43cTSnefbdS
/aABQQ0Gu09+TepqWikgnhRclIXmEQE0oZRi1i2IPT0QW1XlxyrdnXKFhEdgWVMA
q68rzUdFSGETS+zvEMpNb9SVO4RIY5QaRBWGHhOSUbawGcT2Mb65BwJMIJiShe28
e+mgEKApNlVNwG0aYpbxsGYrp9B3gdnVgGI6LLmK1GQDiw58CrKfRhouIFsn9Eba
8+28hh/fy0/kgAPg1w2RSzPSF4ycUfKPeYY3/NLFzJZ6Gp+qRsk2wY7ia1dS024W
2qiyUVbQvG/xZ7rqFuSB3MPQmHawgQJ6GZzrswRjPaup+YKZFvJfdMz27XptB2rB
IjWolCs6d411p6FS81XR4UfWJ5Zzl0hOZ+zUfc88niFxrbCebJbeg+gAqyMaQtq9
6ptCWr2uPL4s+SPlOln8SY+riib7Do8ptBzrXDR+wg5xi1xNXAgypeVKRq8hjBhH
STOTc7OHCXNo9U00IrBK1EqH2mU6SpHDYtjANXpMijV81IxP6NwjXdQH/oEnkqcn
RpUL9fKW1Hr9jX3cqV7EaqWhMohUJpOmzcQ4EtdivfUCAKcFMlvsVaVtled2+bHC
ZpkvPyfTwFy0yNSPdHcB71LbOxTOGuGmTp+BaMobOGjiYU9al9z8hp5CGN5qtHBm
U4wX92R7BA4wiCzB8Rxxpt209o2i6tuFXg4ttbXyehH8FmQ76qt+mN0kCj9lWgr5
oZ5g/pQgbWxwuC0VPli2TQMP/HBc8HeKfFbvlbjkGKxHG4vZt89hnd9k1xRz/CpA
bghXPt3ppxNyXg0P24O7WVS334bm19UgjCnlvoL4rD2riv9tbiHKaUu5Epr99ENS
MX3IKZ9cOa79cJOZgKgOGdpBQbtQPG6Uf6a+Ztv3j3uEdvAzhersZK03yWjknR8B
t4jCwrOpt3ofUu4tA0v4CdVL4iE511uUSgvDxK0J4GoyLlLCaSnhfAQAa92hZpnc
a2uj1n41y3PfClrERzcez/VsWrZmw3RvmVRYHUyqJce8Atb9fWbvIymNaZBC3pDk
eDU1gurGLyGEp/NjMKy3XnZfroRXHI8a4f855ioCnDrx6X9B/jRirCahwSthtCMT
AOtFF1Wazn7fKz5siQlqGySKxpH/0N3b4llhA6L3wzExw8UjSP56GRwTEk1qh4Q/
1nBTT0oEW+05rrYtVy1z19jKpWZIiTlAHpvJuO+yTTXm9DfHgIWVYJx0CdeZA5K3
3thRukFZC+EZnUyXJpC90Df3j8MkVzy+69c7NheDyxurUjXo89gR+Gw7K6wXlvnu
6IRDWt4x2FZcDq2uAZEb2GA/N8uciGrBJnRLbcllKaSEArDGY4kjguQwjrUQg8+C
wpx0BDpMBZXPsiYlayNjSGlBNvHIzb2Lb64+FwN4FzvfTnT1bdelpQBALSj8/MQy
vCGQCZ86pdCqpJQl9yHHjMkVP4HqkCLwwNEK+l0uf6Z+Hwr6uiHAvjqVE0axeJ0V
gnl289AeJ9lCXFjx0woHGRHLbNeMaykjYPJhFQgx05m5lH/zksRDnwljXI+y97Kl
O1aXeU/+m1aCl6w2SA9dxuAyaUztytq1UTPyWFffiQkfN1iaCqJJfv7un9A/L9p1
W6rs7rYiRT7aM5yyx6JEi0BiZGDmjdIeA6aVIkD9vmyIcGb64J05WSOckyp6g5AJ
7iH+DOCPMDGQy7/YIL930mtmo6fCudnx3kZxZnwLFVUB7aQ7QyeiB4yGHD7NWqVH
40SqhqWHhi7coibZcbsEXhjI6GPDHDITzLtRrcpgiKfgy0gWA2cFTRFDPPRFcZQO
hO5EA02K+7s4tx6iDDMA/ttT5vGxuSIINKX1rSa1D57Y0gpojLPtoS9kLzyHc/qm
t0evD2VHVuC+MSsZgyzVbAoIj/ZZ+zTaZVYT3ImcceEkMN6OCZ4vB/xmQhteublH
G411crKpdNqObYLvsZx7fEk3L4OdQyTsytwM5plEY5OVSKJ5IEaRrbz7Bor1n5LP
n8yXEsdqmsjUEbmun4h3m1Eb6miMBL9Z461DWGpWV6s2JSkDxF6VfNklBrf8rB73
Tiz6mlMzuUQyk4rn4tVCQnBkkw2RazfsGAtOScNb2VuVmOp8nTDapchwXWgOGAZr
0K3OMJ1QnHDPklkSqfrPDpFJlYnYS6Z8lknNXHVBn+uvp+3Xwzu13pbsBrFLwVN3
0IjyPY9yP0lu+jitcSL5tn6AyAN3QmAmMCh/CVggSvWsXUANlk89KfXdIkKDNa75
OlFafGHOJ1ildXJRdZ/Y/Kk7fsxe+YCXREcWo8XsNBno7xMXRW/x8Gmx21aR2v1m
tebF2m2HhUjYrfjK1NFrket3sDyuME9sDp8VD0Dp8Tx8PcN62k++T6RMdVafpeDJ
sN1TXBlmj57bDg4+Yt4XIm2VsWyqUHE3bpyagcsI2Vgr3yz9VoIS6zvRuSFcUXTc
68KNSF0YjIPgQUZRxbvQoeD9kc7XI3KDWLf6L5p52juGcibOk+EtS08GKMVsuBNY
poD2YRh+yIYFJu/XKTHLQfhb1hTopmdEhDWwDWwKO9xDHQ63ExK5cbi3ev3wPLfJ
k++p1e+yBNxMugIN8PFTset8mJQT3upDNJD/hBcS9L/OGpClNyt9FwJyp25NVXX0
sjsJJOcxRbpNIU2KYMPg82qzchi7KqPffctgvh6/UFxVtJYC9CKEk4s/+F2nnSwa
cRLcgipl5M6N7Pw388fBxJRKYUQiZ38VsuggQGDDIXQ0otKM8GNtVmo3hJS0nRvY
YxNwz3Pj7UOTMizS3wnE6Le5qZxLA6+9I6F2VnNqKduboI43uxtPmfJTI+wczQco
5Nl7NJbD0eCW3izg6j/gD10V7QIg/Nx06S+zc8vbmpKoUTE0NRbyoBrPxXBam4Ow
ksYnEhx7WOrD5yCf/mQOH56pP4WdGo4O8K52Pwxj1hqoy36Znuf7AzTewdVlASIY
hnK98yTxbV7zXmMzsG59+WfXz7uLbylFC5zjGp9FlWAxwEzNt3o8kNcJlWc5Sk0H
YCchZdbIYvZ0TztWQ8HU+xVHYGQdMlyt0R5MafWFiA5i+ORgiS7v1kgRXQOpcgty
bZYDhsCILBvl3huhn2Aui1o/3Md+ncyX8RjLokR2fliVxSuoTa//st7tl/YXfoym
4n2vamGm2eJQowa6CxLJ+a2XGifAhrdvKAu5+pRTbycIS14XWhc0uxoNXMRR/lmL
buYdPcIqgjzRKuGk5CR/3t2HURfPzlWzjGNBn2kkXvXjvsG9MmCwsFN5fX4pEgAK
OTISEQ5kNXy7TLi0hcZ4NO+JEJIiNH84iCV8ktOOCJAhbR2bcIdHoc9Tsws/lCSk
RwjRKG4dyqwKxoKW67VP7auSlHOIqKnVw8JKD2gbriQCWOtOrnvU/IWPVA/FW41C
vji183Xx8y5kQ1E+Cy7aOQBVERZbv0q+oj1voZXqNdjrZpBDY0TIg+wg2YHAtgnP
GudGss7vX6BFhDoZDVXFtq0kjGYPesVRW/b1uYOrIkZTNPGV1KYDu7O1IVIr5xHn
843XWPcdJ99Dto+sjTJ/Muqsn2v4LZum6V6nhwxdcXT535EjQ592slIKBfhdiW8y
bG+9TJObE6NL4kPMGkP/+Wnat4PSgSf6CPZfQ5PKrVsZyU3qE8j0DUCbi8IrnpM2
t28IaCPtzqqYbOZcYbT2rPhFScQB/N777R6J/WD88lJatA1Zkgk3uLhkdW4YnnJh
QNq4oaFSm3bv+AgZr0D0A6LiVZGpMpd3+dt7gh6iZjOJxs2t0q+bFZvKlVPBCqPP
oV/OZNHVuF/vxcV5mVfr7r2vzC5piU+oB68PNR9sHrWX57rP9AnxRydoy7KpcjbS
Ell2JEgFBp60HHbs8wluaohl5YXEwEyex+/XtLB2L4xxXWpiItJk82Y4Ri8NFJvu
sMU3CfHxaPanTi+m8KVt2woa2xSIiR7r2bpEwZxGGP79+B9980dJJE0OUmkbGzPn
r4dSK5D1t25jFsZvVMLoq/v1r26z+I4NH6IDiBj+Ds8XRwEGT4/EgSvWDSXBEv8r
HYnRtWBYBqR6s3WJkmTq4qzfZ4sIb/URFU+Z78XuTw5erWuFnr/lGsxZrfL3dPvh
ZL3idexHpbtupP9w5cdddeREPBXUM0VPpmE+dLrhDuTtm0dx/7JufrnSOmIe9ox5
60cmO7oc1St9rFvlVicJfFSJ+fk0YggQcljUkgOpn7I8Mjk1iqSHujBEttcHf+5y
3RpTTDuGoC6jC4/xJlAIGcQZCDd8bx6uUAlm5XG48y+rmLw/07c3ij+Zyb0DleD0
5Zpbx40KrCKrBQd8KpM0uN3ataG+Ik8pr2K2VQQKJA/p8KSdQx96QU++flWOnw+x
qqjiql4Ls2awZ7IWsYGT8cA5OnMg3eXdiMe/bVyTos3ZA8jObz3GGV7IrcMeB9ss
kDgTQKd1/EezsRN5QfE3dSAuDh4uBQfLCpzb5hhnFGGu9meU13KbBoG7kJ6//ozL
CWrEmYHq9dyxsoAbKw5GiOMUwcolCaxVSajTrTjmP+f+TelafdYE1Fa2SzMYYKMy
Inix5ziZsQHnGkg4L7WCevzCEkYdusetQb4BapL0VyYkFbnB6psBalBVV8KWDMfS
OumqP0NFgVi6tBQhiCMI072N8ntfSZghAdZe4dXKvPmyDcTrwVLZg2VicuRLzgU6
KBvqpDtjJr1hb4SlxgOi5X6qaxPld/a7++e8iaibidkZQh5GvmXWPoJwuANO61N/
IuIFc+FS+cz7D5gVDp9gPVcV79RVomoWqbap6HoXzvwBdrmwKfb7+DaLft3/oB1Y
XQL1rSulVwghK4zFvs6Ak7xArc3i7WLdGdnmTaquUKH/bG2GhoA0qNQusVczOFcK
u3ahQpn5EjD+ylJ2gmbRiAY3YzZf/9t1PK9S6VPJLzCVUASnlWGJhFt8lz3gYUNk
DnjMaTyGkVFC6DMwloo/1tJix3HlSYkB56d4GMC7fEQ2E4A4SotFqeBXOLV62Z6K
ItkrFW9sDYL5sfJdntMIBH12CnKn+mpTqb/c+D3JQh3qnMiEU2ci9LiO9Xsc9QME
TNml98uC71IVsXIGep4PQCEIVP9+tSlkOzWs9eN2iqq8RpPcnjhTsxEY1feISj0y
zbXe8F7vxQPBEszZkRbrdrTf01FyO0XGF8YF5mgvT3ClwAXNIxWtX9vul9AypTl9
6nStO7qiv9mGNR1XM/ZIQeAxYAMoPHEDCtUtEKmuzUFXksyMKDPKlMM1j6rl+uY1
ZYjgT/tcPg3JeN3v8xiIVNFj9A4A/V8IkoLpNa69ObjXIho9G9ws4D6kJodM3Up7
dpGdRn5AV3l6Su5bMy3udN1z7sVyQPDixaKscql9BbAJKU3Wu2MwOoh4OrMbGUPY
ba4/J2g3/qf0WDs5akeQhrSrY7Cy3m2sH/kaojfaofSjsWYfsGVV7Jok45xeeVQ9
4W2dkwMCSH96kRy10/p507k0agmmapto+u7FZKELdlKC7QizZW7YBe+yuPCHHMFu
/w2+9ippyZ2COx9narYCxBK1qPJInjwd4F5dTncrJQ6ovtTp89jxXIijL3/nMRtS
XdRTQGyab8ljWhkJTiOfjUGb7K8W3KWRBK1R8weDUlW445S0Wytk2cDjpsG33fX4
nG8xVGgJdabFt28usWXON5xBZBBOyUF10kv38JNGSnScjRCZRX7W0E31OgsRdung
XxSzqvI3js5Rbfw1A7F3gXXzfaczt07c9a71LHhR/+H1xCEoxPM7eOpS+8BwMf6G
WDg70fAU7iBELfJgfG7/AycTPmbOgnbeHB7Jvw4zPR1dazvmmvl+XBKOR/s9wzNG
QZga2LU+WIf4/hKKG7hGtj30+q/iaZvXZyEG3SyUA/FolvBjznqQYMk5Mbwl7CFc
lHVk2Tn7zwxrZ14q7cfKC7NPddB3JBY6Sqh7m1HLxxjmQvdQjL3N+9oKPtHu8Ymc
pZZHbNdnQAWAvX271P01BaBJe4TkQWrp2Mh/nmaMqQmSWpb74SUXqv7/rukdNnkQ
xmKBaxvf7cNhKKdi7QPShPalYyu2Q6D/LSTx+bU4QANA32ZyboJ1ejFVUNLxFXhs
eOPdWlm/9lgecx5a35sgG3kohHDdoSi2qIqI0LWQ0cJrBTWYkCQxbdOsRZIl7bsl
WagiYJfeYXD3lsyxqitLXVRpL8vzfZF8wDVJlWYMaUKyc1ZTrn4g+okStcXkpdmL
Z+Qttkh8cyDRw5QgRE3LjbAaJdUqy5NgxCyUvsuKFRyiSFfbfcR90BTL3AuWoKhc
fcjvGIg2/Rqj2yTw17liWnVVygVGuEl3pXRzZURaR5+cyuLnbmbjWPbDIV2B8DAd
zZ6F8N90VjSjzvNpvPGh1GkvCt4xErliRSZ2MSAJcTSk/nz5SzRfezfjSe80lWKd
d50lJAb5y0AW0bZpcApNuVwo3CNrD/Mxi3VJdCBlC+Z+Rxhm6l+v87kT9PTtM29G
MjdCRFITr7Ut0BMh75OBeiKtswudRVbWmfItQMeDRoQ0HGQaw6cKKNfE0FAMNOM5
PuwRbwAYrUjmR9b/hItu4+VTpof3dx7PFDckZvc5n2Eq+ZeMyaY+S5KB9y1Gz8AP
qkm7096dNJmgb0ZY8VkZO2fpaAnTeTk+5chc+5QEgOIjwPQhUDgqTM5LcOVVzgCx
zuhBcoyrRZXsON80gDil2XQLBe9ic9K8dG2KyfuLl9fTfQwhDgAhEXvT7jFK0gUg
1+VTkSPoXfBlFa02TDzWJr1ot+GHIeYd2UqM3RAg6rzwhB4VHjQ0eQJNAP3QU+8g
NRxr8ddGlzqi0HVHO3iaDdfQlfOe2jLbyR78rYkIFAT0bW2tPQaaA7nxd93dSMLC
VFEE3xZPvjpT+EBrsqEqdxvcu8fUpUcWPGmnX56RMirru1ZDajU49q3ImRB+qc9U
jbUAgghIvsKYaxcWbqOShqjJlYbLZ9o3L40eUDXAEslal6yNI+axwxL6ZVzAZQG5
9gXkNXwxhsxZE4o3PMyV4atAvr0PqgPZbT7MBeLYp461dLkvQs0UPaYOMFhRiAO0
bg9p60DhrYhn9iSxJRq1569ah/jCpleBznb7D6XoRcUgObY85ng/AYnebdF2CkCU
gBaxU4OAdpth0JRpZaEx2mn2pi3b0WB7+Y0iowykqoqqGtC/BkDXrraYie235uU6
H6A1upuA/wXJW9Ptw/lCXBcQnNOTWRRoHfQtY/zcy9vlWJ+llyeJKABIrVPf4gwa
ce4SzJDZEQbX8/f6e2os+YIRkt9y8hFLe/JxOFwLUGtOcmDy87q2o7FyWophEc5U
FpnS/qLidznXanvJ5vswBNLMoogHdTM9ydkayEZF4uBVYaW28/DIiJHG+g0z7VD1
nyZpBTnuDNG3KvEqyU6cR0uBvdgId9KRTqdCNF8qeOc0KOGYpLlQSCpgzBHYMdaz
rZHSPQauCz/mkZYoGStkyWNCJTOLuXrDjo8Xn0qHA8CyTPQcFdaQpbcO/j9BLc9Y
OtXBzvAui8nBGUNJRwAyZht968w4MRBjv+wwPhvGiK3S8SfMP4yZvy84oYoVdd25
vz1e0Md0rPyyBYQwWWnwgsQjcvZ0tw172pfZURJcgpYU0Ip8md5QJdBLaRWdvEm7
SgFO+QMSmo9OhU48vbQfCUiHnCfCuWPr55hN9X4yo6gt+L85AaJ0dCkUgxCG6SBg
H7Xouo9VuXjlkdFfu/muYxm0xoxFg73yyhG0nrYZex35bjfFlWY9GQQ4sbzzc1rK
vgOxU32RJ9T1j6f1dRtlzabpuixmA+1+pRLNsFLCVVWJHGoXoC5sO2z/+ild3JCw
zRaUAuBK6eXLF7PKNdYDTlCMImmKbxcKV9VaO+fVzndZUNxDaB6UHlkrJk0TLklL
pbdBTG+5eiGtAKsFd1Lkj1HHcPeJeQBHUoJbtbTbQuxmikURPUWJri2P17x3vQG7
+ev6i6PylXxi2OBtAfWHP0zNyspHay+qEIqFsYTYbHLDgrlZVHOOZa+1YxHgT/WD
AEJwGjF+0TiPFVGhx+N/JfDGuY0BQpwtt8sp149ezAmIQK/FmjQrVz/Bi6pH+c0z
LmXwGuzfi8cNXs17nL2XMr6tvk16JfWtUnfv3fpYAIv8aVhWhcpnpdsndqWcy76m
0j4o8Uz0MxkPuF1qzNRiEyj+ctCag0glVl3fms33itFXGrSK7GvLiYceGAlCOK9F
TwmfevZQwXpNPvYtSZmuiOXZ2AVFbwKO6+s7QmZFUk7XnPCyKr+w6Y6jAVGMoJO+
k3sOaZGHi1PoS0lFzznTvWnmK3XQhejE+z209iybRx06P/MVOhfRaqxk8o0AFvia
fujJKCsUMC5YvEMmLeIYre/sM0PBuZNBtn8hG8NxGJLP28LYqAEVPgHEEpduAIHH
fM45DgJfhSOwII4ebzzHSRa/9oyxDXZm8BR4zirqXWzruoI2lHql2pYJDksFd+Tp
0HHcK95xcPYvCamGC4vgwLAb0ubTsymw0i3ixniHzbrwgVjSOLbu8H6B4kF+a45l
JQk63ZQnTIf/1ln0HZPhy1G4Wk+DYC8JMCULXYRuSO53cjtj3e+x1rABTBYudMSr
d6HjfNEAu6vteHODr/51AWoL9l3Rm6SxkHpMZ2KipLk/frJinILu6Kl2vqzDp94/
EFZbjBiaC2+zFgjs1QlsKQ59G4Bt4nSgVTwDacZE9+pcKO/L2ekqzGjxhHtzNS3n
mPPHB7bf/n6lLpN8WixtayN1qofh7THdt1XPY60Rys07bVUjyyfV2JpsIgbGa6pS
bPfX+vDngyiifeUQOXZWUXopEMvW4HX/nGok/Guy1Te+0+IyLl3V/pXZUT0g6xRG
tJnO5HLuN+Fz++DJdVI5Gtq3ejqj5jgK6A+UcFpk07KB7SZEvrB9rfntFx4RGbjW
Us+JBoe7P5S0+vYJ508oP/yUfWjAhfwv+XUAkRallyC72AtVXxwInmHp8zl/2SVT
r3W1+HQaNIgDxj0byciXeCotQalgIFpXnUnj1n57FWk81oYCoCO338bI/aHd/eP7
K+yIp1D4KHnlF5B7foSKtp1SucQFYowH2iMUKGk665DhCAiP2v8sCoj0JRHUptxg
53IJIPit4p7nTtsmaDpy3hTXWGGCDB2GAZrAd0Lmxo/MzoHw3JW8fme382vpNfMT
/c4oOYfTGRcaqVki5Ie8VmfHBnrZZ/H6XjUrxfgGdb5Pdr6S9iYAcdTKsOehLstq
qf5JCEhe/VlS17QXRHxJ+Ntl+tGh/8LLXmDdmgcUVQZHmJTffp+CQknxNBAvGUPN
IHCGpsF0yhZa3PZc/DPHkdxDxVRYffA5NHOh/RIijjEIVPGl4P/YI3J1vEhynJBV
Kb2xgPDFGSIh9znb2kKAh1lZ6Hp7sUih7kNG3a3upsqlRi4tAkw4Gyqo1nclev2q
IGVuwTmVUqmaTO7iYLnV5FMioU/q1DuhHCUWxb+GHS0o9IOlBaqwtwAr+U1ZexbH
rSM7XvttvawkaBCiJ0Cb6WGQpe65vVv+4R/ZaBEYppiT0rbmUZ6FKV2gxxkEnFVM
L8+ynIly6mOEgAGw0QV1ASJwWdHv+NtPuumPRNEsuLUFbZSnCd1PRpI5p+zXXTzJ
3FUU25gzMyLl+gEQqwcEpirRmnWGk/GQGI+Nz7z5i4F02zC04HSfb/tHKU0ZJMh9
raRS0QI4H+PI8/xaV4RJSK1s+Iyw0zcs5LbIdp0ytg5+hqAoniLneiydilc3dJXM
/VwD4ShpOLKQ9pcNN44xeHgzL1R1n8d+opviQZlxr2XX/lN36GQwD/75zT9Uvs/r
Ff+Ybl03SCjj4APM8vpb3tdPFVfv3VuwlsD5Yz3lFcjlIvVLFe37ymEai4JGIfL2
2s528ouabKFheeLGyAxv/MCaJPINDcU+G8rV86QjUW7+7NEtRw4olDvlxp+7ZUkR
A9Z304PHXu+hsfVFs6tSvw4o4dUEBj28mlytmWtNazt3SrYauV69jeaLDdTSX6TR
xaf2Oi8+cxf4U2EQmYmtE4QFRuTZWr/QyaN2qv5tOlx/qMhwNkOC+VCajeOrflUn
oaweIaK4MbTAc9duxueK56lmamIDJfooBrRT5gF4uoOE/S63KlW9rOzPE695PHCa
43RcZ39XxNypjNoS1yNwn3lB87x4RxdOP8JsdWcqlLKqYYFrkEo/6EszSPSojfwV
iyVzwR8sjHwPyPrgec5Q6lSjNLiy2S/0h3lDg6M/cC0sOdstZfx5c0ENs9oIbfn6
JJgQMHsMyQcE5aXfPYOiFSUAVSWR5LD6rnZn+B/0Q9PPxxm1HZlRkOae40PK3521
p8MRQc03Z+5MiiYi4xV3NbyXzwiq+R2A03U5lvZDjD2J/XkqQ6/oht65W16lY/kx
R03VUdupTzTbvR8IrMM2VzmxtExFujbC4TZp49t0tUpsAcq0qFWwC7lb/K5qCJox
Smcx2hh3ZOXJbljMqGtlLSdJAUJ9oLnhVHIFY5nNDzrtVoeKgIF/qnT5syVxUhru
GzR6xH4/TSXJkZ3IL6ZaqKHU+dHfzWXPwOSdV9P0ZmBnOd62W0wUqrraff5NKF1A
n6ricHrrAWPooaeGLyesTb5qOWZZ0rnt4k7JLDD607Gees/OTc7HR2apSNqrVrN+
DTZ5QyAWIendVvNBaXMi9MlgIXbcce8Hkpp2i+cD6BKZC7Q34hEFIdHzpL0yHgAW
sgjk4+awgq3JZeDrEh94VPpE4ZXu2CtD3kSRc75Q6dSf/F0Q6FLVTPtQFlcAbuEk
HXBtlcZELFq2rlx4I40EGuhdbIb244ku1XvGKjHEBQFX5NgJD0fok47SpDQM00zP
RKZ2RNyT9BodlmZp4udNtv+SYloS3HQs8fYo29h7GJuhqCypMHVMxCf/hcFR1N5A
sacY9u84rmimnd2cslfzPINbGcCTW3x7kLBArBBrbA/gkDGvmrOwRa7DOZMVUAdp
+zexi3eDbCvvYTVZvYxfB5tN1GEFIHKuSCqcCeyEdXHg6fplCrDIQqgWkQa+EcR+
kilLRyQEy/iz/lCN0KvvBNVon4sOZhKKJBSOoqUmAHWNCd+cR2oKRarK6H2eL/1N
MitqcNfWeNG5/TgpGry4IJaLpKElcrcl4eRQdWkfXaoFAusCgBIBO4kr7nrvjZN8
vrYLnPYLjLfL81B4HKzlU6M0BqhGZhzuxuyTEq4C2mb7kcJuvaiK+OjDBZXXipBp
itd7z80gNr5HCZqM0BIzoC2pm/xRUwc6iYn/mT6EhI/Dmm6ZxFBfGYKOYy+F9h4t
IYCaKYbuCXfQ2OBlb/0PIkulJk+UEkTb6AtPY4qYRcXQMaMVAt3PxpoXaoXBn7n6
BU7DFK+acBRJuvFYK7mWoPax9sA0k/72a479kESXGIDakJmjMVN+qa3a0MNVw/Ad
wPEc+8kzQPsgDDxRbVyGLfJZzwVOu6JFrTF/Kx9yNWVYIQghZPaniNC8v1vmIV5B
a8AYgjVa8lqJGuRHotFSxfthCONVJfz97jiMz8tHyyZ1gEPvlqJp6H9iUEuK/WTA
jRqMgCaSIV1m+qHdCP8ejwoSY0UlVXAAz83ttThIYoa33cSutjhGT+8xL8bida3B
RKZwiruCUT2xgdLJlZGJTE+/PW5kHPenMrwbE2rbaZXXNNb0Ov9w/onGVt0LJUMH
SQeQz2EJJKdiHhFsr52EyhnvkFzP3f/uc7hNIE3aGbF+U9S3RbBHIxZUzjUyr5Ca
CmrdUL3csgnqX8PSYQ0rNXnxNBjFkxzO5zOLPmqWUXqluuXmv6ZquuATr7aYP7W3
jtp/+52OjlKi1Y3E5w7mC0EBo5GmotHJfXEd0fFXjJ3elzGpEOsgg7FyZ+BiFoSR
4H4xazYAb5bN7QJfDEXCVGDF5m5Jigh/oeSSYijdIOuuvO9ZCyzy5O2VtelfX5af
9LhjRBxvMQLXFlIFwloWozS1AB5vtvsax2+jLPpzi+WQZKYCDTMnxLIAyq8O5JPP
YTvr/o9QS0wMmuG6w8t7ofaGACBjAzg6SkVnUyEdSOS522Xhjt9glqiFg/UC8rge
/O44KF3tNSgJY9edg0aB23YhSMSRtrcIuMTtTG9l+iPyM7JeyN5BhE8H47OPDcSZ
2lucgCYJr+KoYahkKtmCJUMzODLmmDuekeJc7WwFBBwlK61Lxz1CG5H92LcJx2Yi
F4DSOAUs3WnCuAhS7im5XP/sIwklScbfclddwcgT4rBYNqVRWB71gLS5azM+Yu1t
/rTq21bmsIKzkSgISTdTGkf//GdNhVFvrqdTOw69C9NtDErpkulS8aFX9q7gcFSd
C5MpcSlgDBq7mWIRJ9ZpAMKjCq6cQmkI+6Hjr/vGOTf6IjWJW5H9nuwtyt1dINSh
DZsid6uSQ5ZfhYnIb7e28gbG7EgJtW6cnAtdiQtHCO240D1UfvsUZ0zhfqvdsbO5
HCLVm19svalgM7QxW5OZG+9mQWJ3vmLGg/QTcreazyRwV7H2wBtJWtMX31hF83b5
Zs2TUGUhk9qeODBrMK8hCVySDKkmG2U5rZaHMlDl9wEsm2jyMpdPbUTZghofRkS5
TLFdlmY2rldhnJIjBpex2XVluyXohaFfxhEcDhpWBg4mFqWGbPLTTbFSQN7FS8uW
m7IxhWWeJpeh6/cgqXQrc48j8WCYqfWB2AafwittIEDn5qdEXV4ESqkYlFVWtFq8
YLnzJ6q9+sYBeQwQ4wp4pdOTcNEVENYGHNF04pWBmAxyxujghD265ACMMN/Apq5z
rai/XqrNyudCtaq7iLHSoE3AGGvavMrF/Z7JY2bPZuWTBaJrRmqqhUnINm4nNkSS
U8laz0i+0+2+CrDWeYY30l7yPeSqZqYqDvsFt1+CpLo2QqdkkfBSUf2p3Rw5FLpI
5tcNTFmek3Ui55RE1J7jie1m+gTNVADM6evXXeb4saYpDrGPaMO2LMK6GnDbHUn0
Dzma6fk5gMSRNxR3pR34bKrq0tYw0SSlnOCkuKlWRVNAaZyYRCHbqwSc45MSb/fr
ntOQ3JbLmsLBTpX5YREYru3jGjeRIeOZ8bTumSwjyhXvCZlXm6chvPQ/WKKnwqT6
VCJvvrCuEbTtvuFfqSneq9wQXnNb8wfCtEdiWLpuLcCyLIo8DlD1d6EUbrsdcQAg
puzhTPyJIPylaG8tiKqEk27W8jKV4Uv9zzByfuV0RlGD9aY1/+hkxt1+hfaiBn4g
R/O00mMSCvwIGM6mLr0eHv8jDSD0Zvwir37he3ELvJhtkHvjOXkiT6ElG3/tJLpb
fmFfhRSz0oK3o2jHfGkk7hCs4aXA6J2TqjsRZHyzvC2iAtVKUNuuzx1UElT3lFkb
z/ENWbmLdQZ0fqENlex2sT4XB0KaHTkyNjY1T9P+aQ6w5fC2k/Z8rRdpwBegy1nr
3KryMAsowLSD0821Ym9XNBD/Afwa85DxveMw1OI1am0MjUHMdyPiMfE1tRN9hn73
qUi1sDCV6gf0PGXOO9uH+ObEqX8Wh8oDBKVDefGbttfJ9rj4o74eI3lyKMLL5v6C
2e8StQCAjKQLJ616JZ22gtdSBayFhx306KGk0y/cSHJmoYpv6UwiYjGrEMpszOSr
YUbWWwck65srzJl9q8ggIi2yt9Zh/GH/9CDrKvyC4Mq6k+BaMCPhdIPtj8bIzHxd
MFmcLwCQXlSXWdvccaPC7YnrLlCpzaX1Y6mQ3VuQekJ9gsah00OoPYGIdH5x0/sL
tPHyt9sdzPYONvTmdK4eSzaAawecQ8mLx4+tdeWVSND3761xpfKKMavg1ssO8iZT
AWOEBZAUpgv8Bb+4ggqSGQvy2RYuQ9YdRu0wr356Q/MYl5ATT3ToFqqeY377/l9N
oEHfTGvn2H7V61qDkwL8dHicoANrzK9ZpcEliIWT/a+1NQLf5L3izxkikcM/6kzt
QOlEvf6/E7mr+GvOrp+nF6x5baSo+Oe7Un7zZ9I+9bMwPkTWDaxCdKyJPFV/Tm7n
Jo/u8g9PAHQMrZsxRUuR+R+CRYQ4BZySL88s9bo3i7PI8EU/yjO6zGozTUPSUeyc
Lv+9O74doagD5MV8icj7jAutyp5NSjhmtP8M2qcQPblzVRMdEi0BFdFavBjdh0l5
rmgEYb48eoKo6iTdbpREzNNfyayvuCBEvyrQ1iyfmYQ27UC8PEwjxxb9balMo8kH
R3JBNDMrjkrOu9J8reNFdSzuKBJhE7dDkOeG/PGAKtWw7O3nolOm4W943P4Q1D8k
lFKyOVU4Ks+X6aoduVH45FUi/0Zg51Zb0ZUm79aTGdf3zrqEdBxxQgonGuiRr/3F
RS3waubwjBOyQ6GBJhE2goryfWdLCUxxBrzOpWXfJAkPw6ZrlJCbVPxJgEZ7EvqX
XAux0bEWN9yKaEe8uBiajSWGwgx+RXNP7Jj1BpQEuJ75eVHeO4YIn97wnThVg0t2
ajRH9Ahicb6q9uu8tKGeJwNy+ihUdQeIIos3hLuvInvWnRs4V7lYYzyMLxBmU+hH
DyCrlCXg/J+cQYAG+rV/oG+GdHoQIOYzluS5VX3Q4U1Bo0CGE0P1vvS92x/2Dsj7
9FWbvXqHQpGnzAucflTgXTxaNfjei4PqJpISnlKhnf+3kOqaNmiPTGIeyUyHDO2+
rFC23awA6S054SB3Ve1oZT65gb2wYZRDl2aI42bDOCRfIcraQVi7dD1l19b1l9ql
CdnUWkESvFBv96xXei2KeICuYGf8Zj0Bz2r1pYS7eA1dEPmg12hJYHyHp4gQfQyx
TLnf2SsQwETD1/bB6eeDmx91IG0L1I6sQZ9mq1DnB5q4WqwoSetoIrCELkRQ3V1C
CyDtYUVfVsZniRXiFJ4CpMFwrdFqAVxE2dNOAY2mM/UDRXD5+BnTz5NcSLuXl2Iz
XZZHe1xIOH65isUV2yD0KVYNkc0YDurxH9whEduzhxNIJvoX4nUMjWtsz1tJ/QqZ
pze70p92fJn9Q9Yfnd0bE0DGkJvhft6UrXLYqCMl71CqpzVz2X0GCE0Z5QsIqWta
fH2wEuiXt0M8K5e+vDqs6Uj0MgbPehYpb1EkDxAkI05OXTj5dNIys3Fm/eBedM5Q
uDrJz2vnGnmnpuOOE5WxhNa5RLy0g4LdRMRQfC7juZtsPj5/Xh9RzjgxttIOKkn5
7nbgbLwQtLxk88hvYwOLw97dUW5QGR6eBbdF6V5dyZW5mGYK1nC0hhmRez/t+nMj
UEIBqUFudEP7/Y2doaeYm02TP5CBJpmgmVO9gr/jINv9+JhImAQNGi/uG69qr5Zs
NhvXPRmHsvpmZJ2PCX/u5xtD6FqroVLLkViXWWim7CI+Pum3NvaRaxcYIPfwhB8s
5QfD1COwDHFbaMoBqbeIzlqg3AfbML9v5lJ+GmIBAELs3RQ0MxKAYEmoeheEt7QL
PUFXC0eM1dIeg2e33LSCq1KjU7GFwKzHJOrx/KDC4eXl5jbvj03d4mDP4cWa19kY
jUXDrFjzrHXDT6DoEMuysEMp6OF61y1wiKgJWPfHQr7wnQIeFuVTILapRhIiQiUT
93wvF43IaWXX4few3PcrF7y7pTQorlj1rxf0bM71M3+4BoUoiCDo7Gk3IbAjWdcD
ES36kk5JURS88hdGyDRk57wARsHWPo5ipRMCdBqJvLOXSA5qc8uSCPQSv9QunLOc
PJBBQ5B+rhuHyCLafMdfU1vfHIn2UB32riabSTy/4XfJR8wdehSdZ9Oyego76OPq
Zq7NZESytyKHf2W9Uqx27sR6HoGlwfp7D0vF3nW7Czs6ShNL3Tw5qjKWY+lLy+p8
qyRDiUrWLqoMzM3/7MSPGGaZbHeF/BHMAp4M1hxUBhLUvfmmbNsf4iVcOfbz7xqZ
AzvpFnSvWhv14UJiaJZh6Tvmykb0DYj+VrGCLauKhNq4OWqZEmc7YiRfbdIvOVAy
IOb3dH+J6otxLkHJo0GhyRNn3P/sUMl2mkGbpzDaD6aTdlqdlY/0yTs1qs0fqEQF
Tjm8U2QCLb3R4QtP6B0gztUeHauEpHgy9Ktgm7o3xzvvTttmXa8qmCodLy1vOupy
eACgCVa9A5ZRTQSxzf1XPZ98kfIDip5DruW/LOibFqM/fWOFC+lMoUAv73xMN8HF
y2RK3fdVbsXMQAsMGPoLBqO7fE+3Duie0XvUQbp6sXHu+1GNqxBazRF4rBvZ6KK9
7AI69RkscUECWGIl2/z10M5ZX1WhUICkoI3mqI7uFqBPm3KtlGE9ehhD/MEq7SZm
9J7moWHKpBhugbQrma0Ga5Luce1NW1a9qFFvOAJhiGdKv05HgS5A++zl5Vr6CGZ9
QkvezgHOJ8bwUu/KExYPYx/a5E2a3ftxchBIkk1LrTSKrBjUCEQsg2uMJCiywyYe
s7ODOm4uoIjYqQL1jTLML+wTLb3IGj2+h1H5Pk4SPvylSBVlJ8gJTxzP3dguFx8t
o/5kb0oQZBMc/fLnjnFexeJy+FkMWXtR6pXxmlvaIlU8220W0OcbdmGX41wJZN1z
6GtgO2Rhe/Acv+VY1/MGWA9ei8YyO4dA9uBkb6DetSYtKWY4IDsfq7mrQfiwnB8h
HG99qg5okJHqHTS3Bu/a8AvpQmQZdBJnfNwrI7m8FKCOKVuZzC1GaGsKou1zilG2
5r3BNOdmnxhpjKFo3EnSPpALCG4ot1xv9Capttez6jZ13+c7qho2wloECUFZVGqs
+elvjks+i6Us8tAtABFxtAurSsDtVtkT3oEA5+HdhdCaA2hjihkRl/2XDqmogLxQ
oEcksISvbs+4wY6EaBki9NvEIR2/D4gKArM16VvNEYfqV7MrSLOdwbt+b9b9yEK+
10NPPflrahWN2b2NlcN++BNUsqwi3ZhlFjSwphVUVgPsrOViX0v6RuCo1sm2Hkdu
mnAvYYZaLYEN439KK4f9IG1GdGtYXg2UMqtd8J8QmRY5eyQjlQ+WnN37UfQ2XS7H
kEH7fKMFS0ptVgSqpoh0qADR+3krv+IbzJ4Bi2M5fJKMTxi1OCrwXbbKcj6m3xQr
eIt1KYdJjwq7lRINAznR/A4/RgV4GLbz09D+5tq5gHH2mOESAv+9nU1hMeyES54s
35gP1Rf76iARl6Z9eVwVOdr+MaJKy3e3fVuFChg/kMDgcr5yy+JUW5fC0ueeLYxr
9xW2gZ/ka8zr/61JslClnPyCEy2iqTOSMp/070LYcyeTDMFU8ni1YBmIaWsCk5NL
tEOaq63tp3kzxbd2J394fNUkwO+IslGCoeMvpXE/O634nV9l8tzgjOTzGf3+WeRv
amrW3/MUbvF/QuDwrI6tVeY/N/uzHUmVW32rbgIQ2fJ99XsuhOk/99DOMxIh/yTN
Iz3bAogDXNgEyQcna5JFKRq150vexgwR/M/Bfy+/A7kFba6m1TfqCqp4zRQA4iiJ
u7BnvBGW42ovauJxLWj5eW1V0HeWWa4X3IgpHebn1mt88kxWlkQKtPPaOe736XlB
8SBWTzm6bF33v0sDzhrwMIDBrp7nwCbYM/J2PtsZ55YejYHSk9QL2DF0tMZirbOC
kXKII71KPqya6gVgo60zKwdXrFn2tTCNoV3ci5EffA7dwnkxtSOLMkRjovHB0bXt
8+qR2C1GXBrDo93RSzpZcXzm2vTSZzN+aJzLnYfdE5QTP9zjbyg/lEnRgFdB/I0r
PKDeiWnEtaz8jmjPaP6zlMHZWip6MSuP2J6fP6d/QkbebxqgOwhMB+PsSRnKEEw+
SFEza6+dtXHo1YwO9imfcn9+Tc4tpKIVdoSPc4CHS3/bce5NbRJuiXuBFQYLr/fq
rm7Cdi24ejZ958pD4EbYVdKz83dq4/8kaSZWaFSwkYPnkJ0ReFtzbtggr1oVT28U
sdd62nNh4IJgJPUuvlZq9wFYPF7W4Ljg1zqihTV3QgwHjMxTmzl0dLXoZUlBezoa
g2Ktcty4cWMstogrEdhXeTJuI2Toih2EQBxvuI2ht9xEM2x2GCK/0Yb5o22V1KAY
07gXvKZ4Mdy4J8M8mPpZ8kfEUBSIFg5zAOVO6eDJtA0cnzCwXJT9yMoN7sx8q1Wp
WuNEKZ4a9W7Bat2uHnA9rTbNrPXksRZNWYJjY377P1P/DT9RGOBG9VPsxldyv+zT
QA5HTHcnrf7pmRecx4173KkFj0eobcgEmO6wqibBMQXBDAX1vJkAsqCb3413dPm2
Rarv2yEXaim4jhKQb8GB+1LMBuj/bDeWHMleZzf1w3sjDaupp1rFczE/96T6qSwT
u3LXPRvobeE4Ub7PCNGDqBcC115qsFBv/G/YH5oADxEBfeFBCRB2iAHrirpa13VC
hlRhL3V3sy5GN2TUrJ8kz4+3u0aOrWNGFVn9W857MfxeESu8ey8PvHOIrDcrFQ3z
U3G8oKTZ27HVTLpOOeXaNCm0v57mKyi0bxoE1sioFOhDJIrw+XKGW1XVRTbMplM3
SbMkAmHvyXdBy1Z9qkuSwTtI4a/ABvFX0VvHgPN8+3QWrI/dTUAU6Y8inHwTdy1+
YdnP5hEgzPZPS/bfvS3XwQ04IQzR0ENoK/i/FO5pgwOQrCluS4AdSsGQk7BXZrso
mLJjO+WArUw6a/BmYhrdVfZ3OCjHtnyn0ZmAS9/tkZIOSJrExV9KfnORCz0xzoU6
xQlz3HiSFs1LEJ9vBUGc5dwVpclTgdjtQQFEGU/Uod4J7ctQuVDFnLOAPESmDkMI
Mmv2/xl2XNX8NbTOf0j02ba4ceSseQ6P+R3LR5pcD2Pr5rynYg9KlcbDv5/cl33h
yB3E/t34vJNVRV8JSQlz61LwYoB6BYBAeO7Fw7MHbMcspmWFTbZo/wagg5AWfLT7
yjEL+mvkRPBg2z99btH3TskBbUbbiJ015dZAUnZxaKqgBPVDrazoey5MwS/aDEMm
SekhHx88LO3DXDzkH6l6jcVeGy5yUqY6mR87ghhAR8+RCSYb3R/YIzUmv/mmHRhg
eJwUD43aXuQm6Lui2ibjD06ZGZnY4igva8vj3Cd68tCpyMqx36/8akGRUcOVZAov
rIkwDFksA0gTDQg412uaCl7tcB45s+wMupqEBljQwJvI8tn19oMeCxNvjqnRxI7d
DnBL269eoQB8dgdFWTXHgUGjZAFVDIOhhukNS4P+6Tr6Q7m3hLIA9PKDDlglh6vq
C961gqo6Odi2rco0zWsPGue8eJ9igevKsRFrJNIvALzzmPHNqOupmL+W/vTdk86K
Y9ei0WzM8ZGHkMUnwtUNFcp4RfmEnCYrbaiZdtqJdKwcA914U55RYzu3T0+grbNT
Smzxj7za0/8OH7fIlX2lO0lehUYm/8cU4B5qROl+lLjj5YaXnbkYt1ha1u/n3xs4
4t7/X9elNpYSIxj/JzWYWQqh/4QXpXm1FJStW5TrMKZpgB6xUz+CE6HojYp1K6g8
IeEd/hOo4+eSQkJl1D4vWuTOGYAu9mIa1mGHh7gb6/++m+rHpkBGOukKKeNeio8a
IffA26qkKBvUHhb6W2HmpoX+yyrEz+LYREynP1IwmhAyUHW9qaa3ZHieBEglk0hh
RQFfE2nKFkf/iwiAx/e+Dnr6XCK9ytxGdErKhWfVpfUROauuFJ21W4SqM7f8vy4J
IJwvxS0xuZSWEgnzoagwUTYo6yBTbOsd2hcvKIqr9R+wAd4d7oH/AVo3ffpf3KkI
MKt3q0P7T+Ug12MDDJgHTPmlKhwio+k38F3Gq7pRGWFmdL4zFG5P7Sac26Zgx4LF
Bs2FB7S+L/MkL6dIk1SxDvC4vClbnL3bi0Yj46hkatS/DRZHdXk0s/yflPWPL8wx
FDMxPTm/Lu5sEn5lI772BH4Mw4scPmuzOZzTJ/u5JSNw+jbmz733bP8cYjPdZtTq
OgemZ9mxa8k0n72TD1A5orEMtqpF1TJn3fyyFkUnSq+XZJEwQFbx6tcHg7iu3nPS
eLUb1FLR3ZaeRRB5bmVukz67G38IfR+QslwVZI5g5TsdINbFXCWT3i87GvxWCC3v
WKPiSZXNBK/irWYZ9USw8HHJ0eP265aDVofBcwPPHH95zmpV1krxo9f7aHf4jZwS
c72FdjNznDLdM7/brYiJmqdVcuKqNMe2DzxesvnwHNi9/GPxW1zMjS4EmkTZIgs/
B757LPHczVKRE8U+0n55/1woM/JZlQRNVj9HO74eAslXfCZ/1hZYd6vYDRfrQFl9
DYsAZTXvMYb63iuZ3VIae9kK63EErVVix79ikhjYabbnGZeBY4KKAsagLuGv3/32
zXdRSOsZzl8259lVqU0YPltWkgpQtIvD3hmrxEjlsRjNQyvjnX4Ab5kYt+Dx/e0t
Mis4qDP7s+PSinwfoW8pyJk9LNAHJagshKJY0zGI/5QeW/gx+qu5JMLFQ/TDrQOi
fDPPGk6IOZQ3RR+mK5wBW/puMvvgzQGVn214k3/3lZpktVdrIVioDfRNKfA+lfGH
8O8gkZC0hxwT73abOVmZM7rX8czexC3hML0hlhjoo44+ClvgAj5+gi7NSsVJyxxm
z/BlLG/cNYgJijIyHhcC8n0Gt1D26BXTkfyIN4oHnBwBORFY/NO5PzduHrbUHLvC
1b2b7wm1AOcn3W0zXaVVL6CriJZ0V/LE0GlTCaSJaPocO27e7WZs2zmCY0xyoZnv
CikJ20xKdJQYjHprN0dPFcT48AoGg0LQ2Fcqhjax070CbSbk8Tt2JYiBMSmg5Vcg
6JgA6IcyECAprljUUthbK/QyIJ6FQI8yjObpaTov//TIOLv/e3OHfL1ONYC5/qe9
LU71bZSWoqAxz8MMhAtIb9IVwKqVWynWFBII+lNzEgRWPg+0wbUUaWn5I49eSazR
4J3fJhGv+c1vXEOhbu8fiQPQszudSp1Wwm0gYl8TeWa56/2zxzrL7U6MVeloB92e
2uA1Oe6IZlIlVModtH7zFKjFEg9wNhwgaPmoJyTyhUmsGM8sfIqqnwdjCw61DgbE
gEcu2ZCrTAvd3X4KUy08kTYXiGAd5S7j+C1hhg5hgcC/oO1AN+knaVMPePOuyOUO
EDNBIF3kOy6E5TqLYWAcb89id6ZRDRBgtF4uGLeL2gWJxWv3BlQDGZGSxb1nb3qI
fPa1R4JYw44Q1nXEDbIoU8sc46f7zdtpTAqlf6cbDlMgo/qqIhUK/C6Wq4yhzcum
qB2wwwQFFfhiI8MRiFXOBJkGZbYFeqQkisP4xB5XlcJuv8tMlEBw1FBNckji55xA
KG1gOjTX1fHP5AyTUah1SRElFSpVGVGNp5Q32Ey19cTM1eiL8MWuDtjTvonsRuP+
korNsAUnL/zjD3O9AIyNlr9UdWXTMz7/PmKD6OAlyVxJG+JF4SHH7DKrzNrA3cQK
C2Fkn0jUYpoawAIuQy1NYYmT9QmHqQrGVuUKU5o4CKxtjWD932ONbUxd1/W0u9s2
aent8nlpoD9OZ9ENgwIXLFPtc7nhblo/sXOpxisAgeEL2xOXXxCYKcWKBZr1Zcxk
1GAO2cMo6QTxzylrA1ltOAGEx0KAJE3Wf4NyMfemjnlIGhVEgZ+RuwQ8eWe1O5QC
LFOALpaxp9DWaPQtwGXLOJofnt8Bi1PyJqqdso3ACNwZvsw/NqSmbGW7TVMIE9eK
ZJARWX3frkriygQOd4f8r8liXOVxy/XW1EGhm9g4GD1XzYxDuqkhhOHGN5jV/II7
wIWAEgfIG23W5MxRc0riywv33xbQoBPp07/KNLEnHBwtD9A4WIdllfMJlmSfIDDQ
dJAe6OMFJbivFF54Lm62W3vEWNb8gtgd+sMqjCdcTQlU5kMf39TA0v4Zekow1DrE
ocfmH0ZhxkFaEZRm/W+rTFZE8+hcVatTQ1sYOtjy1PU35yrEcMTsy01Ig/ngd3Bb
51gxotzmib/nYrVCuuD8yv7cUORD3TVcK20gaWzp9M6Qqeb2zXwEqPFviDEahh3K
jIvs7gN3undsgbzv4XkC0rCgXdP9+hZ+/Kua77jUepSGIFfJNsDGDBYALAvHG3hH
aGOrmROgNtxAIdApLUfLH7VAQuNvxvXFx5d+YmM7wm+1Dr0oeNzJhjFk1/3+wIzM
Pdc1v3dT5jUgT6dLQ47LgWIVINFm2hxQ8+P7iD5ZJcD2dU7OnPM13pqLnBRW+7BJ
JGeiG6xBVh5Nwi4RNG3RRp/rgFUbh6DGoHLCw7u9nlxDPEnshxPe3O6563GVLHhI
WJrQ0Taqf+531gyRryB0RI3QiFg/Kw3rKN/sB+TNirpZtOJY29yvb5BqZc7cIIUW
3ry4QGieWkiN7d/mf9E/sqHm5J2BnywOrPWR8gIIjhBQ2Uc0A/tCQaQIpkhA/2Ae
qEThiPsBE309vJGDBmO31LK23d5WeUcSvr5NJqjRXFLZQHpf6WE4T7VvQCzfqVJ5
xS21JbIQu5TPBe78+1HJv4rTvN393LoRJAekiAqnIORa0TjLFjxpF/Xvn17Uq/oS
qgaTygCwGL00ahlTboK50VKF1YpZMFKxS1H+86ukZSq5FC318UrmdIF7Ww8PGhJ+
axDL0RicjV59Vy6f+wO57mrS36MlUK7jfzpQWhgAQXAzD8zQqfNJ3rfUBnpPU9ld
A6Ui83cpOk6oyRdYGeW5+Ep34vQRHXKAAqHXgvB5ijavyJ9KCVcPxHPUqxW7Xefj
nRWoYUaF7brMXOO43D3Fj+NdlrDnD8MoHqNK3o1WQiWotTij1mk04rKRQstUpogT
2ek3TJViwp10OzAYAzUxGjj1stjnQXvJLsx3ViHZW2YJr+tzghJLiYMj7iYW0CtS
4XQ9TtSnT7dKQuJItwyXndZt60jWjX9ltc3gurwgxmc86mL3FNdWv5d36aNT2h4D
HguKRPlt1VP31gFT2cQtiwjcZoFA6JMttIzzTmQzRguaAJqQWvEQ71yrRVAsTpVY
`protect END_PROTECTED
