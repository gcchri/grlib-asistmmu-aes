`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V0qbmk2lvoRYvr2JQyWuu/8clFHrUZjX8yls1PzmenL0ol266a0FZ5wEZ4SuzJ/d
hRAg5bGIDfsQX883odx8Gfk8ZmUnLP5u9k1fdUA+ynshpwRxR/uzgn6fBr6/ZC64
TmeCkKJlMBpKb1z4rfdSaSiSRfl3/3qwVKyvBBQXnC4AUTkAEPPF0MNhuRHWHI3r
KtEHczMtpQjnzAS798Lq5Sciq/6SQtjUEDiId8qsSDShxuAJjFBg1OzKyfK0B6E0
no1HT/kWyG4FwBQyFMmfWz88tORohbBvWdwCfn+h/3s=
`protect END_PROTECTED
