`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MIsi1SBm9vUK8eXs9GKwbfxgjp6I4cHAvv0tVipcHi8mFnXj2aJpD8S6pVUGJqCb
3vPKq8AkjsovGl0brebszsRKT3fXGc0lXQutFImBGWAmTLs4nC4/KjNknTllYqSd
kIzzogOHIxbTNS1e86h3B2WHqgBtdKgvoQpxkyRFT6lMOcfx95FJ8RpzC2BuCrh4
pXCdKjIQrz8UaSPZRutzAEDqtvXpWn8/r6xtr3Vqk1usF6a5b7m7Sf+6TzkoZIwD
Iq/BE5gsWlMmXUhUlabZm18Fi8Bv0TQtqcI4UXwPI2/Y3x/uy2LvXzTL+Vopx5Pl
DfoDK6SjN8bbbA6nrJDKkJ4NDJkFzZ0+m7TUJqvXlOWY2sTqAnyafTti4a3TBGnF
I5nvfrU3eLacafWOGXaG1U4Et0FnEvLLQmA4rKZbo9Ki1PTi+89dY0emnNAk6slE
rluBpDlS4TuOQftDeat1mQ==
`protect END_PROTECTED
