`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Nfh9223KGerhAEhTlQvcgvs7QW3DeqRnW2+iUTeORpwUgQV+oT26caUSh4Q1V4v
H0dFKNrk4yUNQWKQWZk6UcF6UMwBVNtNh5uuB7AfRVNe2cO4k9k/LOXew7xGkKzo
95LcdYuM6dJBKSw19koV6mRxu9PmylFl8gCA8P/R776+CFjFdNoEdotLquQmOVT7
edK2t4dW+f8lOD5B556MokJh1fZqnbHGb7bVFgcQCimBMonkWaVU5bjTOL9pnGki
4uaEUEOqvaEwV4exI3TUVPAZQBaEi/U3vwvQXWPKz2JsX93P6b3+3cz+1oI/Hv59
onwHfbGDuMNdPTvCnFLEXLHSUdl2SO4UYqhY7qQivh4n+xIFn/aAqvrij67yhwFG
8KcLlVA4mD8v6vilqCY2nXTAjooZKFQykqMKWdp+LmLpngDOpQvE9CSjuakC6xev
sJOVoSlqYp4MYAd12q9CcPprfVNDwlrkY+epQLF5Lfwe08/u1LeqcipTXlrM7gHD
h/b+btnpYVo0X3iKwgBY6AePpWmR9vb5rZyr6uIzKPozriTnl4UY7g75oti2wyhj
umYzAeA7yjl5DJ9rhktF5Jh1L3CATNwRpnQRcpy5+hHVAm9quDfqtcMdG1uhQAh6
Hebh81kMT7q8e+i+5bS97O3qOaF3JkkQHmVh9pMgPlexgA8O5wuG5Y8OWNRIcWm/
RBeNvTBkPaPoRfyul5GVGn500DpZGu5fbq2KNlBXBiDDkastxAPadoJOlCyCwGy+
0ix9yRChv99sTx/NnVJ5T8p8Qir9gb1M30WJLqt1EhzUZu44K88922yERrjbseM+
YdnySKb+KHl0WVWxTqS6P3wEkr2sbNWyVHmBzEB8cXNrQBhCQmeElwdgyFrSKzap
MRL3GyqVe600xUJU18BytohtMUMcbrZjmfkW+ybQYi+AOWXEshCrIXgE2WRxvajg
pc51FUU5UvpBPEa0Lcjs/IAaCJa60Vaoe/nUqqNKFRMbFzbmTgMO+HlnMn3WKO0g
g6m2EUXn7I1+Ruin99p0bs22F5xyy3RV9eB7nVuG4ToaCKBxhE/j7OOPnK5KZp1W
BWloEdO48RsvHK5ktJtKBFfxinUX+mlxWg/tgPG8ATBXRwgzCKgXbhECHryXLhA0
XqXPiMP3pAA3n8THmrb6522d+3bno1fxwgZ+Wi9945LcnUnZSuGFz/v8NkKe1UXV
kTJb6kHVbeJKRIadb6l5RA2hAKXlwerXz5pF1UqOmgr3LwnCfszJXTLqYmUrv5Nn
g1/bhEV6+5IyRjd1MEs3F/W45Tt+SbcaiGDMyWSh0qyXP+0O7YGg6xaksOp8Y1ky
wSu8yccO06eI+GZW8wDmqkpxhNL4rgoEbHuz0NXRtArnMa08r4fdzxn5UixNvPIX
dFAu2Vm82XKfBvGxw39RoJ92TE4DcE+tL/Y4BmOu3Fe6KZCG0wGykYQkboXFF+ON
eDzVq+ld6Jn14S8RQh0cL+M6HKeaUz3fhVR5e6qlw1hW/bMFs6xocSqwrqE29OLs
zkmNBeFrLHwKFeO26hSOSmRCqsVBA9c4ZLmNjGOzZZvYTsUMvG7W92o0U8LyTLCu
eBqQhm7nW4wAd5VAAZAWzzVjvsCP8GTERlvOhM+rb+lexoF22mzG+TYzdZAcZJba
QCVzUMQaPaUmTi+YtOBqZJ/yXzECxGGj9OlDWEwCISeY7EFfvIHrOZMTn/uoTjL7
fjM8lBe9gzwPMjjEhMXE3Q==
`protect END_PROTECTED
