`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s+doFq2KXMHVRLq4KhTlVrJLXVN74lxIaFGz5g1G/+Ygp5Gdj2Vwo3EhFsWCYRqa
AMoXBaPvphD7va3wcPCbQcHesI0vYjjUwcdly3kZtV4gaUrDLKzhHvZUxbc7puY5
IwjOMPMnhK7oU3H9As4c9ZolELhjP0Hb9rwPANv5gDXcaEj/9BQbSXign6vk2VOg
cK94q64tQ/1fHMfeZ7vhdL924S8SRMUaf3VbmIoEWuQUV2j8PzXhSOECA2Y2FRTA
mY5SGF+JMormE7wVCT7l05ZF+XJZTsnx2+e3/h3nXOIGTF42E7fPgTAnVmf26j98
KKJmPU3nwxTEV8RhtdvsVtFE8ThZ7wI7Pwa/rg8yyOGvWSgJ7uCTiditNrGZL011
gifslL/rUNiF0Mfgq1xjNcoo4EqK2NlSTkVmRR9YSjqLYd3iNQcBeNqTWTMPDE7j
KK13fkpGvilJLwKCL+208OyVzyR1CNgiFhJdoWJtvwWccV8M4Qq+I1AZpIFD45wV
KdK/Lu7w2prHkzmibvXN/ZJccsr79TT9P6O31mraJzUE7zygjJO+R4FnOayxZk/3
/ihWFcOSLtzpHySyRJzyhGdzzqRqT1hgJyAGTwsiWkw=
`protect END_PROTECTED
