`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OL4FMAyR/Ky/6CkBpTGEDswj5NPwpIi1d7eLhB4wi5hhE7deDgmSVDwsY1GS8a7P
woGd7PYeD2Iy1jjcw/+SsdenKwXVWhO08Oj6NKlaPnQBWZ0Bn/7q+jGsay6wrda7
9VjjXT6CenT5n23hC0eclPBCA9zefbW57Ts3I2X9M4GiFjj6kS3LTRNvDx5oaXwR
qGq7wsW8csrT1iNWxw2Ifo+GlYtrf/kHtf8wOvIHb9Ljkx9cPQL90Ifc0zmuQUgx
SAsYZI1IMu5sOVzig0FzZq7WKPaQjm6PZ9zE93eTSBg=
`protect END_PROTECTED
