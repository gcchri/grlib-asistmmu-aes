`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RWmqDMJ94W8H6dpIDFmI3jewXCEFHv7OvpLnwO0uylvkjz+u5/Xh8570nW8fZWvU
+1eEz2+u6BjkMg+fwgzTZSjhQf6TWReoUoLbmkoV7zmcTzmJN5M/O9Xjbiw7P7Fq
k3DlXddFk0eIM0tNouQDkF5ace8raN9SziWYIsURrZNMMWtL1szClVb3zoIzHKk9
5XS6Ubts5OZCnaJGihfTJ1kfyUcPXPvNu/iMZobngBeLCCHjz6HvMOXV2xsPiDht
vnaF/ydyegvbQymWKsLzFX2lZaW3ZQ29mqf8iNnY3j4d5eKd4nhHeYXmuFs6s8iG
i8VCESEMIwqOo02SkKiPyv1h0Z0pdeOgEJh7F6o9kDpRIkF8L1VmttwEUUjSDIVj
vuEr67pUjbMbN4BXpbZdZGVTvckW8WTUDkVfupqi+4LCgW6em+vSIhvkzWFT5OKV
EhniZKi/B9qtBAhqAD4gCEE+mKD23y+JyrEmgxQG73YuVUc5c96to6sdIhGtLUY/
h40v6kl40cbors/vwh95Sr5wzNr+yz0ccVeX93y+LSh40sKgT0Hd0HW7QeIkbss/
cbg2f1DtAqACRT7LAOsbq75askO3gx76BbW5hE/Q7ss=
`protect END_PROTECTED
