`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XJ7gesqWs0P8RKKQAC/5obuZ3iruHgmiycMiu1ROTInD1N0UPpKUz4iMd0UeIae8
nkyZrTV6fBL0nXQTEccDCBsHnLmVNGy+9WekkT0afTF+0h4PNAboSYDJ+gsaL8a1
UTdXN6QU054xocYDooXqvpKGxFHrHBT2yWg4fYBwa4dSRKwK/w0438VU1AQWu7aJ
02o8YToQ+gTP67dS/AORsvXIb/JV6rtzLulVkbByrJCMZALDCJFUJVP/Ry9LIDPJ
FbiIfKaUz6MgYXUduaXakJL4lqM6gDnfIw05ybYIa6zhJCJs5Ym6Y4PfJ4V+gAGH
Ho7ZmdDBsSKMIIiRLnMb4+qosFsCrPTLQZ45apZhBiBg481G/NXMUH++k9OdpGjm
iiVGNDX7lHRdw/wnVil0MwrY9FGLADoKyBI3w8f9nhSWBkaPesLXAVmUKzU5Vm0/
w+KMq0txlQMjLes+c/A+3Y8+Ea09+PIExJsaqjVWrqZy6qnK8QRLvzQFG06swq37
UWEFjz7bo20GyoF561yjbA8t50NEA3h6Hq5aqAr+SoG8hOfIPscEJLSJc5WKMkqv
0BjaxGFNHhFW4MklltpAVDThNovsK14qiWfo/MsbTwKPb2e96/7YZqB/p85pMYfO
GQ04jXgERJGziytPp/iyTFkJkFSiZYDQeU3fPFB6iSpwS9niggrb8UTFmTauinBx
NA6rDom5Vn91pG0cgXq95R/GQpvYkNhbYuCyP+L+Y1OlTRi9ZolDY9bqp4qBD9EM
1FbmHqCL1FbCFfLio0O8RCHQdMb3cewq2fbxn2msXDLpxQpbCwYGH0XsLvq0GWNG
xdiunqIRUj8N0UlduOfXStsyxnM/+MO87eu70GfhKqcxrinNtnWXWVc9PS+mGhZD
r4yRoYjoGG2QNHDw9lXxKOhECed5n1M6nROueoKc6affCzNfTfioUFgkqZU8GW/g
gV/U0VxOHSxVoOzxjzOAmrS/ZpdI0u1vQ05cQDIWOR4NE+784+v1OmR8MrZCg5jT
4gJWUs8GEKSJBHWTHedUQF9+1zw7qKvS7ZRoEKNSH3gPuQwbRtu98i/80kH78o8q
3INPRFxNYWcbbJ9AYRXhH936CCKBrvRHgrKuLR+wcf90+AW7699A5eUDJUr19AJh
5+9Tz30XgBKRKq5iUZLWaoBlm5zpzhuDB2eTmmKgVur8jgDRVJksqswFGnXY4yam
BC1l2Z1wzpbXL7eS8crDoXSn36ipCU+l1yllrsD2o95LnVt69IvFj/rvgcPXWhUH
NdL5rkjMZWMFzXV+lPcsszRifMgDcVunfFvZNvtny2+k/tHr8iESOcFmqxy+ntWm
5l9nWfyfdwrwCAF2jXhIIHrdjb3Z2hHamKjJmhhplM/yTSIdtmKHjDtOO52nZs50
pT/vr39tNttNvPVWWgfn7mID8oDbzTiOQwc1u/7qV0a06ZB8+ASaRNZ4Mtkhs85z
MR6TrY7LtY8h3YBn/CHNju0jTxQZjtVBeoviOUNw/2k/L8c/5vyjMyl5Z1zLw9Kw
neUXetRpAoGL5tl8qCVztx0J33Wpqzg0Cy+eL0m051V0edwo/8SEaRojxRETuttC
eOb7r61qpE+ycbQ86Tey2Y8MhHj2PuSNOKzraY0wnxYppuxnT3QszUrs7t+4CXgd
9CX4qmPt9Fhms7kJXVelQS/BAbla3VzhDmjjDVf2xJIsPnZrWpg85DmjJzWfPGGr
7K7BtRH2ir3jH12c/PXqc+xHK18mUMT/Kh6twE0+90GzxW+5aC1UXL6ExVpTSGZY
EfC8EV4Pfs2747XUK0909uz7FWnyAevAQ8SBZOvPi3ZUEYt5yFkH0+ommmFVd1Fn
iJtXBZD4+8tFmiP3UtPu/do6ddfhl3IrAze45J1hq3GHNI/NJ7363KoWQhv7PsVK
1BXhxu94YFbQCYAHpyZ7wTRouK7ksK7iSF0wXNMoY1tI+bru+0j86JE+BEn/BUvm
8H4kqavgsDm+Pf2EXbqtxp5YkQh84GDrMsy3DGQHWg0AaZJcs42Yi7ArYel9Sh3r
AuJ9ICmAvzu1CrBH0eDPY9sSxkvFZcb0ljXO8iVsuo78TGdz/BUCtFkB2nE4Xr5j
KMxmvTxW+RvFJcANcPTUp6HTrUwRTQG0ygYFhgwaOm/zd1Tgr+sCiw5V7JLDILiH
`protect END_PROTECTED
