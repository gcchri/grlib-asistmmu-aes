`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
47EMzJWCNinWeFlS+VAkdQJ/ZTZAMiy0//8Mm9iiZpyw0HC0THa/NpQnI/9foVwQ
913W4fjbp0h4NMRdYEOzhrGCYeewnwj/YsGQrpCm60IuuImpzSlscTu7fXAH9f6S
Bvxk1QIF4dNVoCNieToDSPfsVpuKqsK7pWFHyqJzduARpQh3yDrWtIn12tpT3I0v
L6kxZmTUMe/VfHLcpKcOR0DsArdIWkORQD0FjDjvcLhO1jLR/dqoBcf7aMCx7pU+
boeYgOlmyHK13d4rmWT8YYs493K1Q8PKtR1Emes6dLMHzKuE6rm0kG80otNRVRwY
BLWLQNhtsHEHpL515OtC2w9pkyNo3XVUUsaPvwlOLlG+ui5p+eRyMMo8KVrxNPcQ
jzwZIW6kRFXA45so4MBiJHvW8bWCE7ZgiSfAWIRb32uD3O7kuZ+FYbteO9JGFFjU
`protect END_PROTECTED
