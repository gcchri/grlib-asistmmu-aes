`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AROplh36owqWVccBCRuugrk9ToRUte8i14SNPqJ/BSgmH9mXLCVgEaGG3FiUknqc
CQgSPdf/r2iVvbO7Rz5qZD/rFanoMDZKj6b4LX8FF86DxaqyUqFUCLHegGYGGHeV
Ys8Pr3MAX2Y6hl8nU5EPU7gjOyInIZQPDUdI5aya4OgkreD2qzuMHVK/k0WvtgC/
IKX1TnxfUVdhX5L0dlDMChqotH1RZ/CRXVIQL7WaCvrh7FyR+XjCD81Lh3Ynkmnx
Nfk0Aw7iZSqSehA35anvMnoof4s8xvnou8e/+tCN/erlIRoVWHi++ASvssfdm3qO
R2YVkOfs0uOOxKSF+MQPVg==
`protect END_PROTECTED
