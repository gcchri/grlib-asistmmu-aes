`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DHAxguo/W0fuA4LUAeaK9+jbMrBoW/PHYceQC63avx5Hff0HJwyfnP9NiHDSpAg0
yiuHccJYTTn0bUy71ipRKFxHKrNTZLLZc+p4SehtSM82nkkp8PYx8OMNge3mEM7j
gckZfMiozpvdBsq+pmdH9dVYH/wRmKSGispoMS+qj+a/jtD05GaQV4BZ6vyuByNU
+W7eR3knIB6/B7Z9RgsZlS5wrHrzkSud/rtHTc0duJovmX6PJyU6RpaZn8mJ70Wv
0YZdwN4Qsn63YGXxNnFhZTzXfduIt3QISF8XpvLfDjI=
`protect END_PROTECTED
