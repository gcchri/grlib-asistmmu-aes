`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+HR4yktbwR6PIzCA3TGFNpiC50u5UqZh27yAttG2ZUaC9E2ggQ++UXK1uV8XOaf0
XAWug4zXI8Yj7Zcg86opeUebDm/sb2im7hZn9PCPLrK/svthiF9NVwyBx1TYKdOh
93tGtiHFFXmtX4TKPU1ARU8jEyNgU7zlkmynstxUnjRdYScUdS8EogOUBRDmEO2Q
YAGOp0XbxXjmtKKEZO3Lj+cRR11UXFRpWdMYhKeX4ApaCqUeu9hTv23eCp3BlvCf
fRowVg9t/lfWad5QBNv+rsEXFTExH77lr09TIwHQCKY0GNqqDW8/Dj7ltj+fJmdK
akrjRQYnSsgh76Bcd1Q/i/cvq8VfFPwgATkqg4lj2WgPqvzUgWpKDATWFSUt8Bb+
Lj/2oYgcOuk0kO9VeOoflfeU+u/CIq0O1ygMksV7ewCFoNixdxlXaAvviSNuiCjV
5RG6k4zGQ9vNRetQHZYqZwGJ43balr4LKI1PqMxX9V0YfQOAFXZ/5BSqqjMiYYHj
aD2Wnz6JiQQ3fzAuRp3Jl0Tv+OTkOyAS7rZaK1UU08LWM0QdDoKQPRKvMY0xzKZX
vR+Cxdw4r6QJ8ap5n9I5jw==
`protect END_PROTECTED
