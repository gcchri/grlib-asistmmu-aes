`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
abdsRK+0BAhqmBFCM3BtvjcqEq0Md1Uxyz9cbZ++qzm5TXjXVWI0zLeq4o9fZdjV
24SXRUbF1Fuo7pVJV8oL/NvI41oalupwhbygs9Sh2ULSIlzet1W58Z8LHnuiZFy4
ZAvQY7WiLFElzufFFqKpZUJgjPtJ1ntryekKYmagSawG/qTKe30/4a1qdjZetQH1
JskQ+rJ34eJK5Hy7zZmmrrLYpaggzKL2SX0uduVB+FflQl0vYyHDwiGpptE+7F/0
8aT9Jn+iL7QBbKKBun/CEcBC+8tQ3xuFhgGKlzuWDSZeYXCMc6eT4PncGTXss+/o
P4KTPyPdSoO5o64J54lYHQIq0Gwd7KcItBUzBU9biTX128nZHmbVEZn/7iwvNBol
kkkGyzpxGBjEMmUpt5PAk0UQX0goInDT+JoWxEHiSl71apnynZ5b1WnhtD2K+dhy
Fc6TQaZLej7qOov5tLm8COoPxIzln1vQBmh6v3VUQv5tb77l5yU8IH+tXOJJoljo
rzFJYmCBJPA4Cg5+YbuRvJy/W4lnNSPjvL+eX3d0d/6AwlBIrBzSLDQkttUCLcv1
PkBrTF6wHtalgbs2khdFq7zwT2zEOTyNkEQHi1L4Pu+WpfoN1N9f0zNOh+ZySOOW
Dx4LagUupc21fEvS0ZSKjl5DjKHiAeva8c7AxUeoUabi7FYP+ITXs6v697ljnGB8
3R5nZWR7qI4YS7Jdx40WvXaE71eEJepSkGCOaCy3XONM00UXNiLOc5dLxx+GUgnT
SB1wZZ5o2vCAPAGj6xBzXOxPq+PyeE2ZzjN3hGpL3jA24tEctdtDz3GY0jTPVdpM
GB8BzYseFvm6E6caR7vIk7bqR7Qq7Q8s68xiLX0pIHyGg4g1uXtBYX554cr2GDPs
RR0iSs6si8QqGSCxQ6xaZqfNSkGfZU3+eGvTBh24Aphlz+49guxws8ljxOTgkjbK
qvzz2TSHcwQFDswSFY3AWlW/tQDde5Lxyeo4iX9UPryTnpBnqT3n2v5uRYJ3PvZH
QDnkfmuRhrlvGJPXUBmOGt0efA+Q0VXd48uvZezi67TP/QKQf+BnAOiktSmf2cQq
rGO0sDiNGjvqNN1PD3eCL66fcmfnofvd4AILyKSlAjFpg0JXUT2qoGzyWHkhSmPt
Vd0iF82i568EpO58NfaHnMje+J7goJNnrCvaDDWq+fWct1ix+Ugm8VGYh7tlqNLk
19tfomv45uL4vG3zVIH/FrsJAHEk1SMbmfJtpHa44RQfJy9uiPQilAsPMwJkqqhO
kSXQk/3SQL9oaIyYufigZNVN/Y0c2ldubHaePBCO/qjraIKxnsJUhmDewyztWqDH
wZxNhlu7dSA/lJTaVc3+MrjvEfogGpVBJG8wDGYhy4f5DJKrC8CSPViYzVFcMkkW
+qvEybQRg2q4cDUJNyT0gC3IDbLKF3xuAcF49H7IupXsp7Fv9fVaMZfyXnXdAWE0
5Ct8zuKsCl0VcKQOU3iZYuKx7EfQPZANsMiPPz2pfmrLwc7AcPZ/uJGsykZIuuOO
bZXRxR+QwAvcPnxaR3P8yjXShwoy4cLEO7zd6OkaiDgeDjechLkUUL53WIqTvEk8
4bpD6w1Qrr1etrMYnsCi6yiV/0v77KGwDOLguqv5fEMK/RGLUx1jydhwqxNAm0fP
hT29wCBcBlp1kBLwW991e3uCJm/8hSyNtXzHCOF5dBQtKnyMOk2IG8hW0v++qw6Z
t7hOCq+/64204TsXsqwUwuhK3VvFov69NDAmi92jbKRVGdTbP0TtAM4X9K0eSvKj
2rhb+dnqgujkSBsZrKHPlPuGA82ppkxIwCBPL9iA/6MQyqq9QAtip6l/0ZTtSOZN
s3+n6pK1Vrt9xD4HuJUV+UrQlEtQW9ePwDzZTgTcuej3U9bqxzoa3m1+Gc/qmNQJ
pmVyYkrSVuT334haD1rtoBWStEcdfYif1VeLtzIqOujM4WBuWjIh/fKQL9HvrpFR
54utMMVnSlAg7nEKnafBl4mDUf4xHM1iypV7b5h8SBlUzdjNbuOAMSEL78TEH8q7
l3RPn2GMaac3qy2wI6SNkK7MyshrYhFHkPSteIJqTDK5IXlKJxwp1lTAaxWdIhqx
jWaXkOhR8F7xeqklfm5XS+Q4CQO7yuhU3m84hsOvP1/fwqOCLsI7wQfRx6MZJoDd
tklJXwjJKAGItQtfiUhmNUKMdFYarglIvZRFGARNpH8RLkEFolBQteCgMWkvdJ/f
7hlKNAhMV37DMa9o95u98l17DRcOH2gqNuuc0wjyFuOmQ8ivdQjDgLzXSZHhnTgs
+9Dx0IQVqU4vO6QhVgCfPWM+XJPwLbxtalbinInfppR2VwAbwuCuPq4NYryKn3vo
st1F1icap7XV63MmxIVtiKFq2JAkmzXTuZTbTZTRe4kXpVwUVFdYmMuL96/5S6C0
Y+UFWdSw/Iitg7BOZZueJR9OeWaoPvPGQz2cJUWW6gIOcoNYmu+zH35E4PmNjfeF
Cg/WHTln5NAzGxOuP9MSRAYiS7cRLxb+IPbv/C9Bq4ABDRmi1+SB5fY1M/kqQwXG
VzX74OA9G3csRJG6rYI2waRGoEwxYSnYevcsy3mIc/WEaWvHCbQlScfnvgiaBwWX
+OfD1M71CYsiyZW99gKLZHzKAeFVqAgLg1nn7hz8XJtWellHwqcgTParTPb7vGbl
PxX192FGzX2SWVb5Ke1C+tsW3YtFIEqK+9NgktsrOtHCYFr70eqykx5E0OgMFAWo
kYE+gp1zmrJJ/0IuTpTRQ+A5AlCps6aQEGwZCv01Y6B0pHEXCUmv3FGq9nrSKtbV
BHnT6FwMX0cxuT3lDATuK6RC3tTC0BcH0ElQc/NFe0Xhdj3kSgKc/6gCrAPU0ant
kr3nIEgl+gUwAZSXtbds9sekR634DEX7pLo1tNUeowkrCZ9KdybNjS/X7MPetDCI
Kd9qsc66etctw1usxSW8gW7VNlhk4DwiatSnzFHgsw+MyOm5eLr6g/kjoCioMAGn
qvmAp73kKJ/mqoCx7do9OcHTK0SD80IKAiQUiGfrZkYL+mxIVjH20sh80cwOl/ef
dzFxMGvvvfU0to6KAc2KS8VtuboifG03wfays3/FaiEv6RtoIYWznDrSRxBqnJXu
2dgdtAdBAVFxX25SbQt5L1Jf19RlpWsGCjr33hH5/oOdS1ChNLf7kx2E7j+HtY03
rEuvKZ8P2NkdyxjEk26M79S+5l147qHZhYhsk5i5xTLRzaMTHwBbnnS5PIppwYLr
xh9qFhvSUSc+eqnYz5yfXKYEAlxY1h0gjKa3t3Z7cHK7MiY7dLyS8yQFc68OQWF3
hytlX/VB2+9e/FdQfcgZ20PqrmV6nUyYhRklODMnzO6bWexH2uDCyfdBpkBMHbhS
sU2gRooSh+qnFG23IZtP16Tq2QwGcCUn9uGpuoZyyPn+Ze9axlfPp31Wta9zBntA
pTJ62V3BT8RZAVEqCIMMDCafk2rC1Q1e7/h9Zw+sqwBEjTOwP5vedVorK/98moKI
3Ove/hoqmouy2UA//MoHljDyX/kelhXy22+9PDN/HxeFL4+w3vpT/2HvXlFlZyR+
1xZJszeC9iOifeMFVy2OzzOq6ULUZpJKLP/YCrAKf933By2IGhvYD4VbdOP9Cs5e
Uw2hmx3D0wCUHobAA0qXgzNDN4D//wq5b97TmAtSWpUN0CDanqaeiiYkBiiZT52d
1nlF5MPAYY5+AE9DbrTDczYi4iXRNHYoibKBkwDWzTY0G8ls4Ew/7sHrV4styOAl
og1kdEWFiIpPN5rgrrXj2qjNuwUftFFI5fBHEylWqmn/A/usMEOEL6ZsE889wTBt
gY5hVNYQnhCm8z1mi2Bk2MGI87MF0fTTf7eawapq6ITYyeP7jUoBRPthTZRIQgd1
gzQWIoJ6lg0ojQqUQMV8ankU4IPhPe9kqWqNAcul0+LrZDIXYbLlAcO+8r5DHXPK
Iv8fj+ot+4H7+QSaDHVNsudKciFalzEUN5wAKjBP/PxUu0PV9ig2caPcu79fE6Z6
vMxBaJ1wJYG4riJu+tOrIvUqmThztrOy9Qh7hKAvH/hTVdg7tQ9XkQ4bzzgq4rMS
kkYKdOiLTYBoRxImcO3azadR0oGBO8H3UvDWE3HzeLH0t8F8/eajPuWLBrD+A7N6
AsAHPCESeOcKDeb05xMvqsNpHJS/3eRQX5oL8Z21onthfZUmx1hyiOu5/kuGAPDc
4s/+m5ogip2oiz2Lg5Nrb1/2Kw6we5Rky/jtTR7c4Tuk+LfnI4ZKgzi/5s7jNegZ
eqNrtyWVucsu70uo8LQQPXCtg9Y6nJC4NMs19GxkdLWE6hSA7fsO/RtvsU974kOX
BgVKY96VVDR2f2AnGbaNPYzq5IQn8kyKa78MIdw8P1EIrXkVoh8Z/WIZzcBMxblc
HoLOy2kY/ZTPO+5MxUX5aNKq0bQniqzBS8W1Si4VnbJGI52T7QRk6X1nzbfQqm1Y
ptb1YcY8FeFKRMCbCamrr4y/Ss7p1dv7YtCz48Be/ZtOsfi8RbDV4gN2ayT5X/08
MhqTrug2xW0XybO1BQIRxVwE79Xt6zQN06QQ2RPIYD04CeovyZG9LTwFUbRMT+Wg
kCubaeU9Vawe3e7QXWPE5zAebUPpmSKwtWrdiyG3xbwSXtglJ5f7VsQe21lGM0i4
vavrQNkJF5EzLIwfDoh6wcbc2RMV9AgO7CtKwrQ3YqaL2ArpMcPN47DSmmaYk7yA
jJZow3aV5c64kPJMqdwEz8sdbdwAqzlQ1+DIbdn8eqh+/0i1SNe1xfHaDsOqUaeN
VAYlm0Y58l0ePcGmAgWw139UUbjQQqks93R/p0qtXeQiXHMyiZK9hmxmkjTuKchV
hZppSUTauuARbPAqIbeDisxSDRekO2PUsLiltngzyDhBNG32vfvYoKGC1cqmRfCh
zRYGm+xncK4BPw1dvGBlkAyqvmoeNTdo0N09iv4bW7T87EET+G3nHiua2HQ0NByR
umEFp34z8FXnORjfOrcd8ZGpTOuRoKRnIgXJQmgUwPYdhjCUVG5lSkJSp7dAFcOm
9s9bRIao4XgI+AEVUFP1Ebqb8GkL2uFJyhNorNyFAJYiG1+UdA6B1Mli/vKx2Yf5
FInCYU6OxD2Lts7suBmaER/MDWIc++solBOAOU/UJbfqMrStHdRWJP8Em9dSFi+I
yvTzxdVv3dYVsqFgLv9rs//dsI9qYv5CO4rRY35ZXttWZuAvWSWlS5OXEr1Af34E
aMi4w0xsE0YFRtvF63/yP4R8He0Za4ucF83CMwtXd64y/hzc9F/JzwxINNid5RyJ
phV8Cb9Q+Ejos6am/vf6dHredRw3mzk+kDJsRbgVanB+mNJJOtKqcqPJmp/fXzvW
RLOMdvLAuWZ4f47LM5Bv2jTBgTb2ElMtpWf/yE6ZifzTx5eVDKi4LQcSsrWu1t1O
HVShIV+0GDt+tH9lrSSnmKSyC7exJuvZX+r0NXloLSSVvZW1ZQKhCuOOGkOdCITF
LRO8RlqxKvn3QeIkYzh7OayQJpvBSNjQoJsZQ7FfXVAr6ea8SIJ5wBfZrx5LoTm5
h7iI8X4V2+FQlb+sqTAddd7DWt1CxS0r+EYWbP73jSK0c+s7Maln8xQZjDx7NxOW
UlAPYjl4k/MznJGd+89+MzlCQSXBLqgySQZPsajIg780MxT0KKVJW8eoXWYjawO8
Z7aQfNubdqUBgJbHAThSR1jbJod6/iBZtsR6gLWgAjGTUgUm2Fi1tzNgVJ6AlTM0
fD/U+tWVSDnLP9ybB8ro8IQfMwqtfZFFGhSLC8vj9lcgXPJV51vkk0Smu6HGbuox
vTUcHQAnUo7tcjekP9345sS3J3uGEcViDkxPqiK3AqkzjbEvUxgBs07QbAYJXIVE
vRf/0fiI5sdsvurW0hyMbj3TkMxMJV/X/T/Ievy4g6A/ofqMAHgUVCsyJRZXLYxf
AUjjCA6shqLOB88hogu4JlgNoYCvaXyujE0S2LVv68cFBWMeg5MsIQ9KNunujiuK
JFf9eVh9wGByL/2iziH6aGVnKWGuo4TJK2hfq+CIoER9Ed0nsWjIAmzocofRpP50
usHhnh4YhK2Sq2CNQndyXvZ7WNYNuB8XgwZH5beOb7ImWbbzsgtQ/78LllAx6tsn
iCq7Dw2BKdOYMuVHtb2x/y+elEYadVBoyEMc4Z7BFOZOgI/Mw2hyaOp5+P1ZkSuM
0b5CJ30I3UA3UW7Xfma2yRK4fnucJx2o0gcJo90DpSEkDP7rGmkHFVUc32Vm8lzI
i+igB7kiK+D1Rh2I9/F+qQGMgoc6KiHatrpfAV067nRkrw9A8FdPOaUMhtxmfxg+
fdUjH6Lg32FyYWMZkgmNUYBWzj1Tqib+DdNLcPk5LYGvk7lZLotHb+8GPeajjevC
Kbp0QM9eF7QwUWbQuGANKartXPt9IvWkkYZ/XdOczOPxd+NnktppDWDZ33G1iXYS
ho+4Lmm8TvNb943i3XYes94sT9AaOnytrDT3Sunb+Gt73GCxwq64qfKxf8qJcTHD
mc2iRLjQc/nfXG/MwmBItXWHBXDKbEHxdtaYJiCsjzHHDSw+SKUrKHN4TxVp1Pz9
ma+z5ozt7hVCSjYo+iwwenSpmIJxTqqW1LiaxNgUdXjUYgwJX4lA0KYSzG22MMVN
labHaBauYKnRB5tzZV0z+WiwdCDYMWh2k6kkjb7OPy/swpkNF5PgCSUzlYqTDGPC
6Duo2I4YmmIXluHX2TVUyW6Ph5YGFoqGHvoWI21PKJRhWCn2XzUpZ/aQjGJg8T9q
bXCm2u1IeX8ijC/gbZLr0m7isUoKUmU39tBtJl0S7Prrj2xRswdGQZeSqgr2mtSc
w6v+YDaTWNpMTYrgMN0hTchAs9c1IjQcpxSqwZV+MYZjW4rYr1ZDsWKW+IwzsuEK
bQAU4JNjtB5jwzMOZ9/+DGKJwobDLY+3scHmRX1LANaf+n4voOk0LXWaiYIbQLPJ
ly+N+r/49QhccPoKkD5X/TTu/qjyqBRnixJNWN3mo+bM1JwGnP63s9NwbIlp9PJN
nOiBjuS6bWb9H/Rv4LvjyfnWZLIFNyWQgCRzpb+R9/I2MhTYlNA61d/VNlZ5fZPe
AAkgeR4z3GMwAInYZwlYJmS+P/VlBVueg3xX7r+SGiKtsC/K+XBf81lhj4s3aYfM
MPRyQOaw9RTDe8UmC+UiXwPh3N7/pdiHxi2W9hzN1u3mRHtWogydj5lnJ0Wvwwuf
q9q+9m8Bx7wTyLhv2rVSMEc+x13cRwboGRUEVcSr3VRRzGdaORE34noqCbUQvSNB
OJs4IWqj8uzcGdsSd+LV7MUcRgfNFah4Ju5GCBSyzMuTvZ/cx7uCvjboUV8uX+AH
YMK4oV0/L5IHACDKWb8tUg9FKpD+0OYL5w7jkz0fbTg90ZkUwpfHS6Jp8k/Xaw12
/DpEbrm+NZzdFEevGSF1U1KI9UsdlGQxIcEtlEcfgTopjnG4CiFnDcdWd+uBKle+
DNIGBOPpjE4QlXQ1PhGNbr7ntRgMyeipwGXM5EOO9c3kduYQ7UJWXBhpBjLuqWOW
UIGJZ/KfzdOyWNKzhThabTWFe47TYxNQryKpbJWfoafFDVAu7ZY8uhSa4WDAlvyW
HjjS+FFZ5+LT2cSwRFH7d5Il8DgxU3orgg65rzV3fOVeziCh2JWF/8TjqhHPlZ6X
2OH3ZtdIZywpC6oWAmV52cL/OBbCgnRRvz+rdbwm5f8B2D6fO3eidk7FqnzmYkZM
Fowz8/iqYOHwRp3MMWI+Xs9LZ7HYix41BfdfGkYg9JEQjhSM2r2DyuSOuJKIO6xF
pOS0JHuefi4SIwQPGc5nqKkkNFwY0QUtlQ32PavF5gKRztjx7h02riG29nVC05qc
0rjnTfB33FfAkO4BZsJkWXBG4xOpMnB6SXDCxN7aAnD4Ih88KBoMv3gyoJ3nDxlE
v1PVL+jQ5FbIQ03g0AqiQMgZQvF6bFV7r4fwM2d6VWXsYWmil+GExVsq75/Aeih4
LsG8Y3sI4QilwwbJL2JyFwntotgOvuPum9B7qGjV1EYXnDPcUmg9iBUoYpTN7Xx2
yNBKxZYQBmt5kTsTH35v+xscXdlGvic0UE2Y0UDY7/1YsZCst6HSPzefiHj40IRz
mbO21JI4hIbZNNhfBUOsFpchGOyp/14YSJymIP2IadpZz9yT/YMQsfRH2RMBm75f
/xNtdFj2WILCocseZBffUkSWlnFRUoYgvBf/TxIlrtHXkscrM8yvgdREf26ZcBTS
qj08mrEaINuHaJ9Cujnu4kXBKX+yG2656xtDZdM9y+f0fXbnrQqTVtNEcDjle45/
o+UODanR5o2bbgm+Af2BMcw5yGmQ8S72jaQDRrAe9DA7xyRYBhgZvySqQ1U/wyiS
d0PLvJ/isI+TelV9aFegXIido17PM78qFX6lGlYu9Or2VYX++WWvJTcrKm32Pngl
OaqfDtOu3pYZp0OagIW6GwbiZKLDqrsZdHx181F419J29QtwxeiNFQpfjheJ5x7M
VTHNESfmQ7gNclR40OLdszy0gYfpPF1y2iS9zl31cYLp2lkIHp6wQTvzgCE9+uef
Oyno8gGo2TuBWH9ihNqETsx07z501FWlR2222Ow7wVMqRvL7hXusDqEl8buXJw1q
Fb+wYVBGTA80UWt8HdfF9KQ/OPG/mO+xwF3fTaAjsV+L7kJBGXY9uhr+p8sjrZYq
ArD/0Bv0nOxontjftDJNML8ebL3k3hyJeCox3ocUj0HvF6z/tR3w6bbPTssO9xgj
MFUwyDPwuVUAqsW5SmmtL6AH/KQUoHsf8e30YLfQa39yTl8MO1WSYrSv+PfMmBD0
bKtyn2huuP+oNbK+ZQlJG7O4PNMwqi2LaLhaHNaatIWXbS6X1bc27WgWmkU+cu0T
Tn9VdydBGZpzImhgT9qqJFIjkq4x8Z8xO08jZoJJBBWmBelDlgzW5nmSYFMLgsNq
eBei+qpmaA+Hd8KQnYBZgHSvFexN0CuEp7Cokz1Q+avT8eYRHCmcy3ywvL9Vg/NM
wU2pzliBZPnGZjhjPKefIZ9EeBetxP6oatwP6jxlZpVRMDzw9c80EFlKsPxnongQ
zIb2+d6N+JiU7M41vJUG2D4uaUCY/J+HekursVVaUHPlLQhWO94zWhzrLaObtlRE
vzo1ZIsmyjsgg0mcALLc2+FOPZhNWH85Ko0dEEUieiBbrdgV9Wk3iK0uCO4dG0s8
pizuahXKzXrVEvn0zRPgJGA7mcx4wLhbk14KSZBlijOduQlSv/jLKh0acNgoqqY0
AlCjEAEqwBy3pXI8mJQgbD5JapC7Ad8ypuwyLqqoKmawe4H6pLTEROUX6ccTWg8K
ykuprfiWmTSLpY7PqHRk1ov/XUD5mealSIW84tjkbpuq5SX3VbCYLiHeJr00LF2a
b0GvFeWEq4lJqKZ0JfLK90wxfbwWFGZ2MbKyX+xYRgpaMeU/lv+OWQi9ghNYRzBz
U9Fg82Nxh6IHPfd1qbfzpjNHtogPGwyxM251N9QwcK+3XCedXgNc8caGrfOvK4Ud
tVqt2CMCKWaLXhvIxTc5UA==
`protect END_PROTECTED
