`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0RRsBBvQvNygYMFrMf8wvbUMBjDuEZCcEZ+eKJVJ/HKYvkXGTtwjG74vsVk/wXtE
R7USpDcJhjHEkSulrFFV5uT2RpUvsv9v3GomPw6qQRWS85vMV+DkiRjDM7uEaHG0
NXDNBYMeStl+N1hAMdE45Rk65dtKM/4TDYuA3rkiko7S5pikK7QiMNc/fG8rhd2N
b463gpXtwZ6zXsdcwNMg/livVMTYzmdnOnw5pwOBuTCYPh2LdHPuEZb2pEZPzS/Z
HdpCdZFQecVhDRV11ngAAn8bENvP/WF7D4z1JwyIGX0nfoLgfG2F0IjQ+uuXJd0j
rPs6s6XTreBk8aKOe2tXRbmisU8IGyrNVFp9v+zoBo+yJvm9fHnadGyCn/ft83ae
gvWaby8iv5XMU6XrbeMs7RSbJWlEXOcfxtkaFAm5SJo=
`protect END_PROTECTED
