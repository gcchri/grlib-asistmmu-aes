`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8LpHSz0or7DV8+K5FwxsbWdIYTLJLrTv8UCdad/+DEoI5tprd1nCuYor24IsjwlP
2uJ24ii5ftbVBF6jEhXV0iuxTnbQ/bapzZRs9o9Su/ChA4PXcV3e+6gAAOlK6Rqp
p3teRmqjolYK0BZP+7eP0O0BiD4/UUiOxaTgt0SEbPw35VUpOVME/GNXLvoLSBwK
PQeaNccRvlULDr5ZW2EPXSf+Zn/78W1i/k7Kded7TP/izMmHCXGVzotP1VgwoE0V
oPn0rXQAGne/KehniK/Zag==
`protect END_PROTECTED
