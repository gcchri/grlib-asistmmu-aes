`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q50GfXjewpb/G5zy8UiY4tlI0UrG2uPh4BvuPZxFH+dKbUxALnFVPUeedvy7hFtF
RgEicJb2A7kWi3jZP18kwPk3pUA/rAwGGllEJw63lGQgYsetvBBnjjq2aoOKoI8Q
BacwHjIbBy9FxXfDgY+vRcsQLmti+9sIksN3wtfDVkB6CbAU70aKTpqIvVnzioOE
YDn5WwqW5kt99nBZMqPkbQYysGaymJAwQ1boAqOx67M/DLkfgRS5BEJKshm5AnbJ
0W8i1H+nVhEN5P+ynG+AKZlc/ATvtfhKFdwiVFZ18mXs+KGqS86byKG6++uXV97m
6FktibDnu2KXIX4QHqAhHNLy0nGTezuk3Cgh+yd8vodImYfE04WLY90pMs4nuGsY
0/ZhO7Rwvn2c4eKlAMQdME1Zb994WfiVG1RHKdpKl2F2hNEMQkpP2SiDPP6TlEJ9
gHO6JnKJBbPIAmSqliYzT27SC6YDGjhY53zCfmUIAHYG/hZ143E2VA7X0rYzQ2Ws
`protect END_PROTECTED
