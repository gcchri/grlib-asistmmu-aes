`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L+zZ3TwZGSA+gA8gFCEHtbDPbaZlJW0sHIX0WQadBNojJm9Q+29TWU/4TwhpseDE
+wZAZn17WFFLdohXMIFZdURn7WgS9uey2KMJP+uGtxUmFED7dxiO2OFXmL0jw8YS
64sU4iG69itxiXP2ExH3OLk04bbF2WEKrZh9U93K0GWbsQSrhG4hxRvzJUJL4v1W
xt77tWhv3rcaMW7AtfGF6dZmfBvOanBqfXCpGVXFSuICzzVdltW2r+MrTgtQdqQY
1gels+kQ9m9qgM+Pz1mx5CKdywTjdFTQqH2EpJQZC1zR49dZA307ZFxgtPmLJk24
ygQvtvPpQj4gvan0Bhc9BMjHp6pTVuM3pY2pPRIJF7+iK82Y6X0FrumyOtFWE0rv
t+Md6CS2wu1TBP72ZHH0xqL7NgNKLfT+7Q4JgRQr8WIBaVnHYjwoPNY4USz5QjGT
Qofc/I37YC9f/c0bJl+Q7gH1N/EDJcKXjLn2bvZcw0Q86E3ji4Cq++N9Q5gajEfR
EMI2iv1ITW6xpXqQ+b+/8B+iIK0cLvWCxD9wfdp4/tTgIySoiuUPtmAsZKnIX5Jv
xyedkfy95sluWbAIxbs10eNm4k23lDhHHFyPFsNRwBTBPL7PEpfE2hZI0Us2lzQ6
ZebU/7X9QIdMZVH2o9LPZ1pNiGrW+760VyOgw+7JbCLBAYhxytLKrdpMicSI7bg/
EX/sHghIE0R90O0R5E/xnaiXhob0xEyIIkNmsmGfHQcLWbF14grEhFTapbBHAUUs
9Evv5pgvb7ZDSfw+S5oU3qlPx3Aitm1cxW3zGeQTz/w3tIeLoHZ1Ee6D5uklExmW
GZmlvnugY2kIu1rSQBe7cS1JnV3NWhxH4ChRCF0nKvPuG9zpRVJor92hP3/RiD+9
CJ5pDvvd6AZNa6K8FMXPpUXvByywHBC/NmYjZKGbeskIJyyk/R7Mk8fJHEgx6QLM
bBVVGwsMdtmnJbXcBa34B6lnNgc0OxzsRQ2YYJ4n2lxNW5GYFTFjKMo9QAa0vTlq
TKa1NNbxaceH2v62DMuwEQc7g+kHTHfFuihKuUlVJ/ClmZxUsDqAodicrJ2TJPT7
/dunv7Ayb5gjLIiI/sP5246aV8derGEhThXCxZdzVBTjuPQYU9QOC6mzqWcqlnSi
TQm8b525XUvge9mltIaXPWPxhQd6+Tu/6NIdXx/pgHJyI73PTJ5daUBoM42edRrF
lliEkhkQ1yN29JXLkI2gkbGt8nZZcgNFUmc0o+9f808fRgqmfU4+urd9aEuRtYmt
MXieMr8ojV/SDmp/mpjpz1565lQPL0i0fwrVvW67SN8gLjyGsDVC7IqQT0+wKMb6
nSfVmFkxplsD8+blDVpzdL60OiZuhKvZs5cRQkk42/aWuYMsvKXut9PxBHjMoadZ
zKCV4CraSffiZ4DBgWVwUgc4OPinoZO4J7+jk7pS+FijgMD9+ddQ7wXIsb6TJujJ
aGfV88Fdqpl7AnGN0u9DSWvXuAQNE3gaeIgLMHJ9Ccl3eg/zo3Ub9h9xV8OnXoWg
qMvBMhNf1BVAtBdX7cF1JLjY2NM93jVkcBxbIQdKw43a3nbIZxXqKarK9AEEX4jq
l0n7tbxw2BiqGvfschHvbHUunawQatO+f66Y4Pb0M3vjIZLW7N2YL/Wf5jpNyEtj
1mrGLsHIoizViY5HvwP8CuIDspBmWhCv5bywuXn0FuVsZ6R8smPUatFt7u9Dgw04
oGcibcjJapL0LaRMVLXLoyanDPUb75pN21q9kthnWbJsesYDS+i94hc9SZgOUO4Q
UxrAl2f7WDNAUmksbumH/I7BAhi076XgrIlxQ2IRLnsLKi1z/khC5K6z6qWatGss
6PD0Du00u9Eems8xdXGLp5N/SZMwSzQcweUePhXmxVFnBfFe/CAhhw5HVnyIg+U7
KVYqBjnn26PJMjUvD/oZdqu4AGQ32fkRlSeYU9Q/GCaoGBzYw84PclCo08n6rseS
BmS8jMQxhYmomz6JEN6dzw9uM6fZz29nzgxnGUfskCp2A/9M7s8F4AN57Cmj732g
xyplnzDZ6EI+74NzNekJzX3OxKrOQRGcAh+ZnmLJDh6aNlJV8EY2OxKTDV5sc3TH
z+FIU2K4MbSdl6/WkOpMlx7Opru7Kj2mfarnDyNfFzHmWvlAvVKIcEuX1XDHgdHk
yL98LBPZsEwbIf8ht4v5pSKbWB6tnHPERbQI4JsOmTt/UUDXU43AOSqvIaDv32UJ
ODAmGaEXhYK6JtDH6dc3oApa14QBGI38vO4noIr9EjbCUJKJrcFYLgc8v2/C1hHf
nDeq/MYxceKv2lETuJSTtA6vjtFcjjDPA6shTlCqhlcGJ9oyxRULE+E3Qo1GNauu
wKWZWVPpJDV64AMu0Pe5byurDpY6kmjM2zx0amcfLTUb8ibhjl4NX1fW4X9Sf6AZ
LoQmIxuCEX3bfM78G0FIP8WItM+oq1lzyFUqc0eJoHuz8gF4yhf21e/z41lhgkwL
gDrjSYinCn88M86HradC8dcnTnyaIGjqoYc9z5sjlpEAb9oOl8j8NXI+J+RrfJWG
d9XeanJ+Gs2ynFr0d8LBmhAjvGkPQCuVcIcmBqoWuM38cPVUAjpiiDJ9lstAU2GB
BpJKyrTi9B+1QfGWYSBZOxZZ9ujugLr7Xu8FF3HZcrRtvHXd1Zqt0JGAM0YGtKJx
zjImwfljcQMJgiKC4cmVgBv0SpsG3tjIJB5CL0k0dEMLwQrV8RnVP6DGCG5GRQTO
3Puq+boYGos2a0sZmqy6bFUfHLANFQNe7613/5Hbv90Jg2IVlEm9RrteopxAmYpF
YxwSjP/uD49FkgGv2MlJhewIM8UPq4kM0b1MLMBmZbVK9vNUoy/ZzZFObbWN1B7b
CFDL/f/c5MxxO1RUss9N+yj4lOWpbnWTUe8o2bO5bzYe1p+ctiobwx7UJHxjFyKf
fQyWdWZLSC917Ji9VoJXQ7av/AyOpIsyQFJmJfwtxEjQrFnk+hQsLaHEuZpxHCL3
z7ggK3szv8S2pqx7USdDAMKv6ZiB58ikZjwywTn+sX8D7Kkk7qKQNBGv3H4lwYrG
TpVG60H9mXHe8iRe9+0GxRgDXR93GSL+ij2oxwRD+hmyPZArLzDiO/Oc+bWOGWE9
EON8DqrbrRXv3eVl7tiFKtmdHDJdYqnXjmsFby8gZ9/XXDuFjCpt2SGaN36TMC0b
J0fSuLiABOFza+JYjpNfgEU+N60bywEQBskHSM0bm4ujti5XN8RH99ZOgBzJLLNZ
AliK74k2OfKQSdY4XZ+/vR8D9SNgxwyMK/QYuC2qHBEDq3GRuvOBCgEu9qaZpKLR
LUk8B4XpoesZIenoAsQqDiKzcpSZz5EINW07Vj6GhT5J2FofQLzzWFi4eeDEOLF6
Tnmb+6WE0XPw+BDO1olA/xKOh/ynOrAAJk6elfZfRTZZCVmLp41BWp0UNxvUmUTG
W7+UwzrCX85LqT7y86fRx1Udw+6rM8wXr4ixZ45tLjHF7NBzYj7DfjLS35dJqX6i
CrP7JSajOVlNbMUIQGZgy4juPrB5Zg4jrj26aNEPkZQ6gQZ0zl9QuCa7r6J8biM+
ONforNP3BbGGOcg3ZyH6KpuuRNMz9cpZXjwa2z/GSeakBdJJYWylvbgJ+DckjrFK
ws/zmhzlf0NTHv2Nh3KyHr8tO/Pvm9+xq2KYRb+JJBo+zwtQOOcigesE/vIwDzsh
xFhJudwY4WOx7ZsJBOrzIz3z6sAFTepf3c8OXGj4r3MM/PcJouUWS0MG/8MwA5kK
uDXE4KvI/Dgx7MylwY9DbBAho4qIL948A9ycxPm+FU9aqJ0Utjpy/5b8C56MWKvi
VePLMkomOjahsabzQDEwH5yIw9UoDDOxKsqpNCCxDmscFnGCmHSyCz4qJQDP16Qb
HSlJ5TS/cBuO1oLaSW3z52yr6RKT0FGrQl62gX0r2bi5g4YwpfwRHD3HRlQjRxy+
itDmyN18oAoYMXvoby3qRK8IEYJYATU9fBg9unCSfn0oossyMt2O9SrnvJ5SVvHP
LJuSTe/yLQS20COahihyq4Q/UNcU06p9MB+KW1bPRSHzOrBLciouai1lBGDHQSyd
EdIpodp1Y9BgiBkUIc7K8WtAFzuc/+FCOGkU0LxtN1uaC+czK/v1AA7hTLw58BFa
Wsxt9Wxfrm63CVxQEzuoTp3qwDel4suon4EvT5p/OdL7EpOr+mAoKqos1+mPPzMg
X41kanN87qV6i4ZPDQFNDoaFpaKIoYr9f4p8RaGZyYjHZDpc7aKyQAJJZ3cjM0z1
N8jXVODJEGxNb6PcyVojqngdixae64HONRLykMOItBdSHOiaAQJiEqm4jfzXBOO3
oakcdW4QRLPqKtblQPVFJN940klesrMOFlvSPWyBdvGhm6AwYhReG83QfpB6rEWT
LQOtfG9A9DIdLU/ickDC2JcJiLu0Tx+2H04w/atCtz1yrMYDNiDh4hl6ruYewpo7
Cc171yq9Knp4QWI+Z8OCKffxzwcV8rF57gFg0SeRtXzLeTbBo8czMSi339aBMPeN
1NMzmnL0r9mnt7cV5MSKKLCrvJDduWYl0dxopfyafjjhzTQkFM1dzJfGdX0+sGp+
GiLFil1zUUgI40OKQB56qTFOGXQcCsZKlYK2U4eyOe/TArEd1VtTEou07hsKziSh
p98m8BPGBcIsz9+VubXfY7jomub4CM/FcIvZ6bbedTXlTuK++CclgXKNhQRFGvkW
MeBGfbzMEStIvJ36K0PQ7ZxKh+Jv/r2gIT+V8hbMlK9ZSj4wUEqtSNZwFvFZY4Sn
uMQan4tWMjrj6ZBlwJ/xYCnuCZrFQcXHhyAvooCvN6frxwdK9draGuC7bjulNgag
vh7lfFoT71+q/A+k+t1l4hJpItI9g/tTwSfYY2Eng2YU1V/U1NN42wjjCj74AYFd
xcykJgM5WpMq8FOjXfmnE8nqZwkhaLaMCE7Eo5C162cPV8l5JS+BSimW9/ZXU31o
wGQiNgUdcQPeUsvRKmv1GyrqV9qOgSxi8i8wihhZbnAR37srD/Bex0dPL2x2Ktk4
eRKrrnF4qlz0Hc4FHpwU53uAVbS3kvZy4evFnFm0wMcwLcC1rCrInZl8WmSiPqIb
0/QqEzcUStXp/nS7TcXxCCBDq0Vi2Lep87AaqtKZ36819G6sypvF7ZfdJzX/fj0Y
qITJ1WzFaeACJbrYAByXl6lLVy1UtXe12zFPCx/hCi17I6RDgOPbGwYlVsZ4/IYn
KQmESzmHnkSAq9feyBeo/kAk5FcbQcs5FiNv77cILnHfARFjCkBt3wzOCAYSV2wd
GZZfaigkRizxqWC3prfarlPLU0HEtqrSpdGZ1xMog2w9gCoVvt0Am5+nU8ysp6xy
XHNOPSJMhr1Bu/MaJcg+4MxQe+cDnlSeYK/5x5Q0p+M4HrHCiSKx5NR6CoHczjZT
ezSO2aCyhQfKRteyNKIRdMSf3DbXgwDBgBe20sjob1AEz8LDi6naSU4buZfYm/Dr
oq0MJ1sDHY1iqvp9qGQQH96BU2+TyFH5ifiin/psB0uvfHACT5oIUWx3/YjhL6nI
0AiuAXZ6WhT3tU9/lwtoDCst88qDswOTclBIF2vdVb1/tAQabLDCiG7CrunayJXZ
j0WVzutMCQ3VUvaboy5e0z7fj3SYwWNNCttk8YycOPsfEbB5FUqbJP/H0xkTKPZM
cMyzBrUVA9FH2WFsZ7dVsDtKn7aHUCFTvZTD4xVf5JMkPqHpi+6dGdSgBRM3u4P4
l0cdX8lq7nIlLR2AiFoWqn3zS5co294FCbVEQIWLD+Ju7DjJk5Aw5FMu2wmiuwQ/
j7NzyXSLsYkdXko9At2dQPIAnzJ9z+yQAiqHf2siTJRCPfp8uVaMzxL2A+RcrIsh
LYrDfR9DdTrAbJR6zhNm+oRShft4AhB9pKo2yGClbE06jOEK+eFu6GItg1m/ep0A
xSnQGX0D2QXOv+e+9Mr/pOtd2+DUAXnx3CThj/2LAoLMQ/iAefXHqcrnfha4x7uU
PpTLG6SgcNkLrTGFawF6vl21SsaWGnFtxk2z1AlbC1fQFOM8THYtU89MhZLaKuvV
QGVwnA6oa444bO84BmaNkCqVzDPDS2RZ1Xm50ImF07ydg/UZ7qtQNBWqs4s++Q6a
vhvnaf2icUiW7PIJLVPuDe72bWkWSqYLTSNQX7sMHMV//IstBdYpcx5GpqFR/lNs
RAjlP9bH5u30+y06VJ6meXhOx++jcH+LFGrSHAq2DR41fO5IvFMCHdxOv23eZEEp
fGSxdG4fLekzZ/nkcxM834PGTwFkHB1loStZ9bPmPUq3XUbrCAhEWv9nTCh/HQdi
OsVyeQdUXZWCwOlDIruVj7gQAPm0vlwax7caWrV670vogNi94rTNlYXXlXu5eddn
nmK/bWa6+UpopGSJVivx5g7/sSMKnessP1dXkXDcDnuAxRpDjYCuA4N6CgFrxoPU
FKoVlRSihmj78FjzsW1pjdBSdcrnxdQEge6DegWSLtEAj5d++nmt4AJNSKq71yJp
cuvkl+aDCsz6+VvTaPVdfNq6FV1z/4EKS1F/AvqTDQN5F55JTdQT/IxMDjfgepxz
yrWJUvyRUhS6jnneuWNWt677xQsYOcvQBfkxL80vejE1W28m5zV9bA3pe2A+nf9g
bbWm5phUJxncZIzO7FPZK4YT2VKpqWdv/S5rplLRF2V2n2lLp4WT/nMBVsecWZbw
0+suy3hfaFqWKmIttnyimGs4olJgyvsvLVQcEYSuZ5ApnezEJtslKZ8H58I+FoJK
ro8yWfSC42BidKCIHWWUPREiXmLMzEeuCIOwit66+Cx7CF1g17t3BNClRkeHCT25
DO1rQTe7a40KlJDhEA9PrGWDb7QxNhosaI1QOdAKmuy8CcQMxPek8JZ6EvMxfz9M
C91fsXoyl7hUA7+E/ZzH10xr3aV630FDMpHFPCWOzPo3NVL1a/OccZT9B97vEGQ8
OqywMAS3/oQO4Xhw3K8XxXUfTL3W7Su64vTR85j5lGzijEu5rl/p+nNoEdKUokl8
P16NBK/VKAj/STXEL03qEWRxFlwbWGiEWESyhOFkiaN4NJhfUXEjvpUumDRj5ql4
oeWlRy03uH3OLiEmaZlzJ9LK2NlaV52V0+CDV6m4dnm6FhN+ZfBafzUc1JuFVCz+
A6kUBlpLtWjbeLXvCQanBXnkBnFklYhscQpy5juzU4GalAohp3d3iNo1lNzq3b3V
ILlLLAsJPkUwJPJn7NCJwLicltovQplXimoZjPZrhr6ojr71EqPPh+Hu5pYnZ8fI
NYsxf+S8k0IvWGWaCRM8iywDalrPk2bnKUz6k0jXL8TkgOeW+nlcu7gvoIIvlTGZ
hQnVrAnh6pDfZVaB5zMDI6fvw+qfsyRkcfe8COyLCFGVP7tEJyM6dhEr0g+FfX1A
3/IeAnObXMIqoYyjXKIF1T21S4KF0/MPMHUaht6UdxrD7P7C9tklA6vZiquRGYUr
m8cPNaD3UKVQghEyk2QN9QjnE3DFlETIqoUHOc5zWb8dsfmg1La9KmgqdB467D8P
CrrNnxjIADWj8SrEteoKmFdfRPl2w6fcFzdaHtwgASvtfsbafCxez/fkZq/HHNhQ
2Wby9NVvBMwlOG3iU6Q+01+KT5Sl8eSBeIrB4u83R7xhiYXn40ZPHEDx9uwcH+Qq
ON7xIXPVmP1C0fLr5Vw1vCbhRENCjHeOs2H/oMivYihqxFl7dakSQihc2ITuY9+s
ISYve0Ujk/Hj26IY7szTNxzW8fEaDOgaSevVmJQUwbNZ1qLNaMjKcdLGAQEvOjUo
68InJ7TIQ7A778tDdxn39G5/xzC29Zxw+HlCjqDt8lXsHwmopKvGNyXTtJ4oZM8p
q0fLPrDGOoJC+rr8wIouE81AOC1OrOL0V6HzHv4LAQDu4KITTftCiu+Z/+pQe1i7
Wnu2auddoqYRvZa+VMa4C3Mu96UVpJkBi/yy07nrtxv+m0eVlGkBuGjNiI2gy87s
KYqp/dsO5pGLfR4b8c3DYkVBtgjQrBh3yvPR/fpbQ97IpVNj9IPDnXAMQXYbqM8q
QRxlh8HbM4SGuDw8VEU6bM3oj+IlYUt2Mg+vysIfcci2rsl8OfC3b+Jesf0JqInm
r/zElkUtzPwVtvo+3XgbfXTKAx4GobclWNqNi7qZQ/O1nuXkzgF8uBz6WwbSBqy/
8vxromjwAzjigOVRvJsMEdf9A8kjvHMODZFYCgDmpsmx6l5p8TILaTjcDLKqp8UI
kEL7VaVsMHp12PJZAu1ZxeJvHXKH6lT+4r3RIxH2gherBNlBssuKZWUqvqcI60b6
jTkInn6vMA96yCWF5DlRUdcgP0Md523u/gxyDRwXQOHG8MFPILkSUzdLdAfc+NzV
+C2idGDwDNYPv5VA5+1QE2nwn8u5k3BABKCknCaNArfjjZ+Ob9atbu8yQuflT7au
i7DlVwRsR6NWky1tFcS1D2z8YZoE52RDvoDXwlqi8WX0mx/+cIzkHAtasNAY8Pyd
wLXfSRQkpnmdqf4ewk9R5k5HeFLpKFCvBenIUX+Y5qo/gSg1MF8eI8R9ZvHcFO0B
OJh74+IF+92UGNWFHb8srK5+VtYge2qgFBnFAVFn+xD3iqTnY6+M5EltdaKLhyKu
N5IGf99UjxDIX0JdS9G1uC7PG7aUmZMY8Jwrmhk2nYrYZQHdU3hfgg+aKZUnElSm
6hSp1ZIKhmVvYpduftZUD/SNayWCKCtnlFJ1ZcpCt2Bw80rj9cEA98TvgWH/nH58
ZIC1Q4ntN0smH5Kx0bwc6pLsKLSj6MO71Vjd9D+KDQNnxF+HU6HXhpuJGMpx2b5m
sha5AzHGdqpHHWlyLwwTdakRqMxs/cui6oeWGHa2rtVwqN1AIXehF6IfcpeNdbWq
7WO3h9/MH4prfngMzqrdT6069D/4d5l0zexRqLegm5+wxzLuscNHaM7bmub922RO
YNrpw7IbzJo8lBI3VXcrT3f6An+ziLJEmceM7y3Ry3V2CmBANEjQoauACa3QUt7w
bdbI3ldTqlExtyB0WWvM4bV9zIxJtq9zIslbSjLIHq4zT6AWLPqwcd6vkBEebEiR
8b6AI0FuS9lW5Ng52ae3+sERacZSpth2/uTiy9HxfMp3h10hdUBxP3WylRlsYIEc
yOke79gGJLZGQQOy9aWWOh5szuqnEAOAt19z2Z0Ckk9mJ5+oPzIRa/zpzL3p5tqz
psmDguApRY9bb4FrmZ0J9zHI0Ju2BO9/3mFIPWPo4TQR9m/3GziGrF2axexrsZiy
HXFJ4q+FUd3uqU+kP9OMLNyxxNAST4X8m3Ypcz9SmeGQ8ctpRp5ykkXIeyL7oVTA
wIKWhxu0zBnmR+lmT++pT5ZIJAkqYjBAl1qlUckbzzHm2g0k7+FsIm5DJDj8oA1V
Tq4arYEbV9We9hu/0V2iEnq4j0IS3oYIOYEuIoV9KEKEgm8vZ2HWET/sPoG256Dl
n8/lubxJBAzF+SGbI6Vz5tSiy2JUEauaMM4ku14i38fd37XVPueNJEkbG7Kj/upk
uGXfZ+v88BeKSo2F/bE8q4MUESRpV3oy9PkiL/4WQXr8tH1bd8yJbTxIshLx8Z52
C6d95Rr7AQo+gyKMa2j6XejuYMbwJ/wwUMUleuz9f0aP7TYqxHWHZXnm0A3kXR4r
o+W0nOz7FsJrpZITIrXb9mOXzkgPSwtzFVvSdaVByjiH0CzBeYfk/CXD/7QNwJMZ
PKrqjZXZpjX+bD16qdFYulAiiirUOk7cf5DwcDIRqm7EFxhi0RueacuZZw6dOj3Q
pwK5kZdaX/j2vsB+vuhOYc9u8O1hxYjbpO9fYES09kQvxjxcyfScwM39wnt+40Jh
T1aCUd7ePQJStA9Zlape4CUsfHawYBLXoxgQWpmHHFKPbQfXT5YRtGogynWR1Lej
G9F7Ppy1ty+Kunra0uI6gZ012vJS5Q4wqAFXigVE7Wa9XCI7KQK3dcHWQkgYOfyD
MYfbSFG+qL0oquUkQnU07mIt8gBoNxyToRuAfJa0jyf5hM162nFNlzMCvAyaV2hb
xal1lJP883PIhNW7SzAUoH6bILHaF2AS1/OsGswA0eg4KwK2xWQfbTrtMAUCxu/7
SXLXbcMKu0xm4bi5B/p2yrLsFjmVpuV9b/JgvIPoNzwczOt+Ykd1hG19Klah+x7t
NQMo2Z8TU1bugtOnhHXpunxFSQS7Kg8Y6vpy8TjdLKjmQ+/XWrZUK/kiyyNH154C
DdllCpkw5uK6le64BfFWwA8QwDWamJCYKlEjTR38LNU4vsPl8SASI2MsYIZy9Zzw
mw0y4/Ocn/tYrFp+T/E2p3qWmZcEryMeqpV9DL+rCNagyS9+4oh1bPXNYs/+naCt
5F5zeRXBpLW7VRagcLwzaQsjdPs65ur3Vsqyppwi70kg5ruyUYWzZzUroh7OKzUa
M+4MDJ/EWCO/Vm0wF98zV2PMi0Icn5hFVFVRfda4TG3TVFphh60FjKqZLCdh7K4a
OB+QxMsB9YW5tHfucH1hs2ZT6FvJ1AdHH6VYII1zV6iVDkEkmoA2F084MpLjcwF4
nVl68OM9eVl8il5AxeFSnhqfBTQUxVNzL9O5XyU0IVvOGYuDC/4gL9GTXIL0h53S
s/7rwJx8USf6aVdzKNR55mJ52weeee3Fh/Wc9KZSm1Ug3yBpCBNTRqPLGIafMj6k
jVuO4Q7KV2Oww2B50yx7wUOeIiLNHOQbFFRzf2vcHqJkK4YXnr8bHyDtXFIAPkQp
h3nk2WUeOBIvGjzkvmgX0D5sFFH1yOhbLub+ghlkbkqzBlUToxu99+c++41Z8BJL
38hamKdCoSJpMm/KLUv1eOUg2Iwq1L3bgKl2DYSyfHLmfRMMwW9EjksDrwTgKizK
O0Hk5LX+v7mIpwWH5EHZ2YKLYYsOUte8BdXlJShAQv7can5JIbjfltbgDz5hl5WV
QZmm1HfulT3yt7OAfFCYkBKajjsdyxNF950mbLTlKhw5+3uVFBI0/cSGzvPTyf7Q
AaDraXvLYpW9eE9yut1nWApfXAgerDyi45fzCf18PrSgY04AMBd52bFSGqpYYMuQ
tVSPbz6yayx3dRxe/836/aFFlMVewvuNSbhLK8znzQiCEp91+RVD+xxfBFjcWuUN
z4wD/s00HWHbt30aQVZ4Zj0vbrIx0AR5IAvN7Hpp5kIEsj94QjhvZLQ8M2xQHp7I
p9lrRLyfinsBnFCQTgoviBvlwJTxfmv1IMiupkYabmye8WoxMML6ph3hqMuTUcBI
leVkeGtXnO+42Uz2nyScrBZM8lpWW+nmpWfotRg+9TafUMMUrZ09Y41nUPg9awyY
9411r/UkFBwdMTaMigq5AS8VTrSQmHT4qJciaydKV8ar0e5Ius/owH/BhfoiDlb/
plknMc/eTvcZx5dB4jXso8ooO5a97TooEQWsqS2SgaRxUkof5GyEreYnhv12vNsl
32vjuGt3yeeJV+W6PvXNbji0S9TmoLjOARBSbTbNHy6Uzs255gxKLELZfnxKuQWw
2R5RU1qUpz9Zim/SpzdZlryVlFIfSuq9RJmo9GNjkmVd1wjTiSZluqQQ/gJw5i1H
2U+xkEjgII1F+2ObBAU8lD8bdombTkoPXT8o+ZU1R9JcV2II8Ttud5N9dz2nh/WW
BpStHRr7unv84LCi1q8WmSqb/R1rk5WqkOK7qA86DVCUel97/ddbW4XffYn6SJaH
XzfS2DpvJiKeRlfxnwRkvkgO3X+F0sYTNh4na5ALWsRDRiZMXxfYPL/6yuNG0Y/2
UBmL10ptGC+8LESg5erKbvvcafjjsGD4NgXFME/y+rhBRCIVs6eJPheaHwBMigGV
Hzr2Mdv20yLPa67Bw4YRh9LNRMbTm92uOpwVL/kWuIXPnhCfUbmutCq+fNQNirG3
sSMwhD5xOvn7YzlPyzsJUGNrGGQT9H+mdXEsoNSEG7li26FPRryZaTYpMQjUdyDi
+LPFdrWi8O0qepm0eUMCl1RkhLvWvf6e4zxw6+hfV9tk7DIWNRApzioppa2wLQK2
dzDs+mg+mNhBwY8H1s4lwFFCCO0l5sMoF+AzK3LBJOLbH6eJomdznmlOyR446EjL
sdf4PKFWX581dvcQ8VcA8O8kJaV371IOFe9ogg09ERKFkIwgWThc3EDGd3z+K5iu
vlVYOK0Of5Kyr3hZUTR5p59HqjcnpMKdgHJ9QYSxRuC8UDcWHxUTRLX2gpxuG7nL
BUUDfh6MdMOonY39bpawlYEMvKbr4LGE7qk7TnQSqgLY0A93hCzC2uJX+LgCd0Sq
jZSI1n9GzaBIzkEXJdQKm/fxv/VSJqgHjoBJh29G1wt/AgGJkNtA69OVq3fKSwds
gKvLIba5O9lH02BJfU9Cbi+u8Aw4+P8rDxTapNIf+ea9ziT0jd17wCSoiwcS78yB
Xp5ESnvYbPW/2YfimFnk08hnRRxNxkKV8UYsK0Ejch+Fvntd4syFvEtoRPlVYeh4
LAMCXI1WcDfDC211kTg4hEipHPA5FMQHHyVHrq9BiJ6OiGlBYmae4jPpylZ9b3DC
9qyG9GYbv6lset3XINIT3oALryXHCwoh+qjdMCI1jRviduaHu2BhLIgmXtQMHsBv
X1gGXc8JXWSsNvAbKz3LtLw2R7hXTgBWDIkulubqs/3/VeRzCLxJdVomqLiEYykC
d7GaxQVSSNFzAsbNnB37sPwm9WpdGeS8PYSk2dpD9kL76r+LjUOkDFcSXvllWbLg
Sn0bDUW5aJPjF0boSnOasIYqk+mqVqwPUxldEcKTXl5a7PWfD3kA1A7rWIuzI8VL
wfKUfiyp30e0329JxgZqMPeVDuyRZaAhhhcK7CfNK5HIE90QzQt2rZFQeoSwZgaw
zYZla9F9fL72feoahIT5hZb3TiJTBaPHm2yJd3Xfk09fPpYK4WCQ7Xj3KQ34eBiX
Tg4xTMjhHoLhOMuuBLh3RWtFXzBCRTkeaAvQVhif1KtXfftXiVwkvfvmQ7NUQj4Z
DFGsbqR0eblVmVKefjYchgOnP86yALMDghOsIXHh8cIPhLuDwoHSOb2HF2Boq+sB
tJyvVp5hI7hkzKgX4SjlOTk5/7LH9MQc6cMRtjVmYSg3/QflqhaRsb4CA1xScpeB
rMPutnqmmQlDOgKXYxhNq0OEcO6feXmR7VpRKXmsSpyzm3claqQmEvFxfPi37ewS
ixbiH6+5CjRPrnUSA8hZu5ofjdF6h0owVALJ8EIvJOuBELq438Pd7z/DVYtt75Jd
OlwyuC/mdLgm3/RPCU98ighBgcOy7NsrgooihF+K2fVXmAExh44JxnqkMnfLcp4e
84oEUVY6BRWTmuX+NoA82PTT+lNsSnKyugN7v8LCG2djYvH4/x1WqPziW7d6MhQh
eB9HO040cpNTS5PrTeF8tzzDBEhN9cm/So/f/acPYHe73svCWCaC4496pK4ccgLY
No54EvS+lKB+ueBsI/0PzX7I1ybUPU/1fo+he+LAfTnEjdl9EntRrshNpCIdbv6+
X0iHK5oAI2i0zwHKJjJh1oUibs34QtA0GlOl55zyC4CwDpTXeni4k7OU5TY6WZvl
blDjqC4U0b50pjmyb+SGRUPU6NfvWd1HuBLMmsIw9DI0rKdvLK8/UXNGyHJ86pSa
LpYs6pIGO15htKrnUJoHJ9z3rY2uzG3ZqnM/rtWCjZ9yoQU3fcI3LHPOIDA/56IY
XAj0IV2lA1ND2pEE30pNWhmqSfJD8OfZCLJ7AfVt1VqQNBTan9JBn7Z0sf1aBx3p
xVEzGJv8GraMlqPi9vhz59tunetzqKmYiNdMt/stCv6/ApbQCb3NB67VDBFgG9wx
dJLvjyNTFaclN+6YALlhjiv545GGPdXgqAj6ERJ8j9QlnBLM4loplDQ2S9xYhEU6
pjuJv8snRL7SepMscKGsnm6rdsSpcO0/N8qALvNoywuBTDbrLGzKsCGp89otGULG
jjGRm0O1ZjBIX1uNLxQsTNRkyiXFAlnCTCaXGwz3Uoa1m0JHQK6N9gLxvMPLP4hN
r1ClOnaNJEmF67L3G5NqmpPSoJ60LsLZP75wimYq2IyawmR4E85cJ+qE57xnsdfX
HVjlkrMlcMKT199W+ylCycbT0AYVHZScSPoMX3YXY/ogD2A/eYiNxVILx9HbD6O+
OVaukQlzf+EBwatsfNnOSgUxlFjb4XeMu2IW9sCoJqF0NKSJcZgzqbCk5YoWIk7r
pznSUqrkLEmlz6upn8E9evC1eKw/kA661YtJoNpIcjo+/EyMDwqtFXbvBqMJucfb
`protect END_PROTECTED
