`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hY5BtE5wz29m8GnVYto4TTlRXCYjQb0O2sTtlPeNpNESQvOeNS/lctXbhSa1NM1I
KshBJA9EfPfc6fbP/QfsXTnT+Qw/QPKpJLc2ZNgC/3dT1iSjAEieBqnctEwU8ZUA
ayQGGaMpqNaa7doQqZf7YT7IxeNQR6kmBGTd7xY4/E7u9+VDCqPSxzNKqLfsBbD2
eoqs+VVBtfOiL9WcyroZ7XN0YYhYzLZVHK6cdXo+99Sl1Utxy3XQp6AqEMKdjTTv
lUbYMOfExnEMrFdnOxp8ik9nwhd89X3Fmi2BqKhor5ge+q13G9lHaLtB/uOBlCSh
8bIfgRwg3RLuQWoGX+WwIakPXPst3EWHIrFV2kOMRKfDgbTrx6+sytObm6kNVWO1
ukEcR2cyCq3OryN1qT8jTwljizaAbpokh9mDgYA2MzEJqI4eeuf12DCgetS/Runv
nBQz5Z2GP/TNyxzwu7D57A==
`protect END_PROTECTED
