`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ff+y/V2E1ZoioWZ4T9rFdS2X1EB39mDlp2Lbs/oS6Ja7kUF6gi33BqvUx0ggcw0v
05s27cvpO/y1eal/0RqxxXm0hgrQTx7jdYE/dFGmerZa6E0bLXaOdKOCFfqCaf+r
3X0ySxjldtKkGu+35OHsfXkfMvgos9EEvQdAieSBDk3Z8bm5d7VdHmK833N27nzB
7TUYP9jiPTuEp4VV0iMn2H+wEav0zMOCILmKYSDp9zpQ142oQoXKTbrC3xIFGYHW
i+FwNDtqcWoB290jKF7gX8U+iRWgdPXDmpFexigJRSyqYvbe0VZsNZIO4P9R7iOx
i7oOxQ21BBf0O2wTUoCGgGWf+pBft5qEC3fo0ENhHpq2gQmTCnDJEvyXuo2uor5t
XaaCipDl3ZcLGTgfp8Oe+9tfZ+SK/vUNAQjgVJZxDhg=
`protect END_PROTECTED
