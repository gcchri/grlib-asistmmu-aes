`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+0wj7AVhdkeMj6+DcDl91uwYqH7xi2LQba9aSLvvu4IN/X1whDvF5v6qzVR64hKc
DCgbnWX6xRljhkSGimdnn4ZE+Nj6N5lnd+hF8B/XI2d1MqMyeoMFIHV+Kt2n6Amm
qVDlIDoLvSn4CmdyOWG55ll6OqOtvRhacxVxR+3yHlDzIJBWNn431X0v1Go8LnGr
xh3gtBe9aZ55JeQg1IA6zyNHURiyquOMJyabQVMlnQNTETBzL5gjlrLEMSHFl5Qb
A5wAMLyAG5nApnDIUGsXntCt/fvr8Ig01oqL4GwYjGaVGe15YHNp65M3sAZY/xou
jYbTzXRdoBVdPb86p8rPMDOt5j3oVvSX7G4OiAIDehLH4qLJ1Ik6Y+AvFiOiXbue
4LKPj0g3DrzVv5cD7tSGEq1VZ7fjkJ9JyjYUdRDk9aM8gbRrY1We8RxoxMHoLIMU
uHORMDNEj1ojCz7ra0/PWwbcg7z1tHFaWO4NAx7ur/W3sXfIPTtq94bWGwTORM+c
w/uxyehxP719fSZ8KIlZdd6q22ZQfmCw4YqKailK9MUSNseh7+SL+eyoCc9FlfnG
hFcDAMQXNiTQNd+lMDZmA30aISgNYAvI0odwEBgDXfLEvoQ5LFIz2j3GSoVvOG8o
y9t0F5K70yQsLt6CXVIXwr4nFX1bUK//H9kVGCDZo8XZKsVIXqchrsT1O2wB4Wyo
AqpTDVejwloKM+rAl5/+VL5yeoLosWWXRuhf5bF38Ex8uLuY4gMgTdAmwyQDYpxZ
nO4sE81EgpmD+CZTG6BJoxdHvwpIZMoy61T7a1sh6Vx6ToCXCEzl1FrRoFsyt2nk
k6PK/wZdoY4/6cYMh/DUWNdYlKYf6PF3pgg3y3QO+eiCt6EOUmwNz5p2GfP3UUl+
AFKtpUssvyA9WthEdAXZrK1oQKDjRD++RqJSQSRyjjK9/7lI/A0qjYROB+ihvhZc
GFgxDZs6QiSvMS9EsP2KaL53/1Oaiq9y5xR1UdnI1Ik+G1uNEZiGeH5cSz12UWMH
mXI1Q3Z/w+FpW0K1AioC2A==
`protect END_PROTECTED
