`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
77p17+zeXHzfP+u7kPs7GcFswvCCNQ83CXP3k+m914QHOmIi60gLAkfJeXpxt/6j
oo5AwQcg1vPhQiyBcHmpM3Ok+zbYGZVbl1cEXE9tPv5p/NjFONDTkb7vm/dnVOxJ
O21B8lPE/y6TJrki80zUS3J4oRdLOfjqkzYYslz3Hkz+2w96ItDTfKCXi5I5e2NZ
eOjMbnhm/Om7KbHsxgSDOgiiFrs2QrWIB9A9g89QqKvzCDHG6rHTbcVmRW0vQDdn
83ZGD6VIOcQ4YflLH2Z6PxiHtftw+DhSXkSeupvoyk9R7DBQwa2vc6jYE+N51/d0
oUmxAX4W28a1IKBFMNjvWcKz38pG/D8wPvxHKBZ9eqAqdOCEm6vwBtYHpf5PSXFk
8w0PeEUzLlMvzvI2ifWuBTJi2jU6LiheRoFxXRWNDTE=
`protect END_PROTECTED
