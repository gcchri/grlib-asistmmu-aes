`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5QgUiJ5sAJ0A9kaG+aPlmRPOAsW3nNAA4KW7ipYhrfNJQuHhXF3S7hE6KhhqlQlS
rjEBausW/+Hunah3gN1nFq+C2mH0zvhpxOWfVvCe0s9XGqNf/W7norWYWTn1/MnI
Yi1GcJi6sEqWz5dsMWN2Q4rtGUKfTxiBnKNvs50hVE2OJMfAZdoH8JrDttiH/PgW
vwCwLD3Vp7UxqCPyl91B/0tgjJattcjdXbLOEOyjbQha1UCmS4DCUL3Izfs+AUjz
bZtah1esoKbC3O/ogwEgx0xnc6cjpwxFzy9DbTwS/i5eaXVwwKwIGNTSUKjSUpFW
A5S3Zg5Bs4XaZbZlxpCjgA==
`protect END_PROTECTED
