`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6VYULjViqgdryYHyxlh1qXxKdYgCqIf8sLX4+M708JzGwty/5oBFukiyohAXQliP
bpYIN07uynPoufRr9veC+EsqvmclTYdqIeVIQ6NUg9Wirb6q0bdO2LLYaNwHQ6Bv
JwZIiihhyidJGfKsg/EYFgHAVA2h1ztcTiltL513wb8njvM8jrRww3Xm3dF5O6dD
f6bhXoY72XmmTTaHwPTNxIEVPinARY0wxaakbmX2ogMh6ZSk9NyGTU90fXQ2qjGB
MV/nx3gerFdJsmCUdO4mdOS6hLC1JK8K5M+ReqP/ulalpU7Y1PBl2PnIze8//lJX
gimSnc7PDZ5AtHNZyPc7jhFhOyd/EzFdh0VJ2C0o5ZPAHXvXp4D+mX9lyfblOwHI
de/qxyCMIaBKuNlNqsKhMGH3VmKxNXeStxRcxQM04/rjSnWHvAPWxSKYnSN1Y/IU
/yP9pS4rVZt+cqziobUpv2lLV2+P6GGZEv9zntWSHqnitDvDaZ3xgWUWlx/XKsmj
ZgEGV+4WL8kGxur1esrjFmyLqQXTdyjR5V9aIuoxMzU7UqvLsUIk6pXBnCsX9JtP
5gOPd1r8O6kYkqGRu4wdJrlqtuxMgPNvU3U0MsLyLsAHOGa0HP5eer5C223wt3SP
eyQFaS3BlnFL9BsRd2YBaHMBZIKgHsK/KZJuDaWsN3j/ZpwLhV10jN+sq7QxHy89
XyRuU2bFNHsHcJfXNCRH3NY+tt5dyagXYlSWWFFZcrRUAc4hV1KbgrKzQE/rHB4f
+oYkeE/oYvT4XwCEuXObGaL1KuL+2SJelYF/6ooAmTE=
`protect END_PROTECTED
