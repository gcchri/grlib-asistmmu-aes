`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g1oEqLtrI2m2p+cTgYD1sSFwLx1v7/4IyDRTGpJn43nEkyFJJj5u9XdLRzxp4z2n
23O+k6mUEW9f0cD6j2MCONap2ZD6KAiVCDPMWagB38uBdiBA6FQnauS4VHlFuVfB
CR09+Vo9gQWT4dbKsJqeCD48PflAmJFNNc5Eoytkle2Snb/kqsBePl0qYfTcoFXd
dkXFnvLLgp5ZCzWlGv8fZvS7TRaVpeJeqFozR7l7SRFQtFEgE8IW0170atGQdLuT
bFZoXk/GXjWMOyH1oCh5cG1qMAsGP6yKEVALXHoyigu2Q8dhu7eZAxEswu9AdELL
57FMwN/im9uyUCY69jNoORZahOK9b4pnsQnG5NcY6BPFiDKFNZg0APZQ+p1tKRBb
BgeRT48qlEEPjkeqy6l3OYbEEKe6YTa2vLijW81DU3MURLFZatp5UCubgJN8xDR9
kgF6hjTkoGrsneE9M3I74Lv5rPS4BH/QBghlUmGmN8eWi8UMWVJAIvVFxR/mWRYU
gyXAtvmS3ygBMqzVLx5xIC3dhG2Xv6m5eTZA5sGC0p+B4zqYd/W3M73WZZyqLK+H
yTfQauc9fLdURrvP9pOeh8X+6yRjYBBJHh8dfRrrZnyrtJmOD3epN2EEVtcXqFTA
NJBxNItQIlol+31m/uNdlw==
`protect END_PROTECTED
