`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gZPexX4hE3//ciEMK4IjSvZi24LRG6Hr/XPxZpd34fy4QXJr3w7wmcYSOA2xwcak
fd3kLAv9Yn3u3E12ER08jkquZ4Iy9gFd4IzTLadXQv0m11Bl6PABXsMa7UaqIFoJ
4THAH64dPr2CjLJf+48RncL1kcQhs13+E0cK+Q9lFoV+SyL72GWQt8uZTKCXGfoU
h0NEfYtXwnmPiWkaE4OP4wXR4v5FKX5YF0sHxtvAQvgZOKe5+RNeUvCcIIgC6amT
Ua9QZ77O1yDP1Q5aDesNv/ba8um/6/ykN/hDAD1HfWHGHvNOr/gKUn4Ke2Kg4UQu
EmRn4/6cjnvhpHmtKlpoGb5fxin0UHNq8hyOcEEeT9/OJ5LiwK627X6N6B6m0lB+
atwT06VfhS5emLn0w+MW8bWuDkFxqWfOqI0fsGGBXRaA9B40ypDPDvYODPMvF8Dd
+IiUfVi6YNfn1pHQr5/LDXVy4dcbZYASL7c4efZkUUDBug6t57HvzDpaAPyqZwK9
xQq3VCIsS/ezrwrY3f1yiaX1Ttho/1TRmE7XuXYDT4lrHa4Ly1zqLYXD0pmcl3lU
`protect END_PROTECTED
