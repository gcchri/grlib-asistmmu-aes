`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hcz5GQW927Syr3RLNw0k8HkAOntSjIS56f+rQLWeuX/CD1TJpX9IfiCoTK6ggjmP
pZKhnZGwvHtiTUckHh6k/EkefQTO9D9MOm7z8mcAZFa/THgBb+Y7vvsYty/LMnLK
zYMdcW2lsN9g6jhO7ARqfv41BMbP1o/+vEOJDPvO84EKgdH5xHC8BynZyqFamgG3
3Wtt3VjQ7QzronOwP7rTsQJpiilw9IdlZl9CQqurRLoyM9kMGm3NpEzukvuzeQWu
Mvn7/qhFuyJ7I+9uraXB5FUTbtWP17FDr4nKKv8J3zs/8qoohnYHnGrvAuKT35nP
vV09j32KCfV5aOJthbQI/7ZeGt+CrDdyCY1mi8KzU1zsVaz/mgHMUieIPSDjFOqI
0z2upXATSTQM48KH32FS8N0Im3kbQMYK6j41EX8cH13+O0zOna8ZsBokyoLm1dEI
`protect END_PROTECTED
