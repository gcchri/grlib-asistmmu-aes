`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JvlvcW8r9jlNxA7wyU2FZrvr8Oi4VQ/W/N9Uz5rXeFPI87sYuGsoAUAAgCiDbQMz
XERoi749GAhcHD/VNIWMvn6FKRm1uEddQ7SYBIWMLsWTx0ovjioRn62UZiBxAcqP
h8zmj41h66bt/rOi5nEWVGF6/T/mjAN0mZxRJfpCDKg5C+jtdOVHFd2NI8hP1T6R
itPdWctvtVYLmEHUG89HhVjgqddUc5xyqkZ/W2pJ/8G+TGLJhJgOrBIVML7+KGeP
+t5hBozDeTPAj5LrnCZyZX6uPHWhw7w5tjPaiso1Qa98wqqnlT1yaqGUtYFISZf3
eoEQm5HRaz19PIZK34X+vXgqgX9+GqMujsH5UTWckmXm90Fd6SPcl+c3H3lbkqlI
wBiFansOo1DmHFkZh4UiSrWFTrndtJkWNUxFzZERrO1z3J1kAd5Im18wAes6JwIL
3z7eL6XK8d7rhMNXveTGU1ejiQT8hnjhe/E1ClNfkeUbH3KzoIPf1k6xunYY5fOg
I5RC7++fFEUftNQcybNTtdi+h88a50uzT0uNoUK1xwAjzhXGR6otHQUi+MCXcMiq
Bi/JcSdqO68WYsjcAXwCCfPFyziBfu7X8R4SRPN8VBIGTQ6raWzx7dfoZesbHlzF
MK+Zs7NtReUG6iDe6rLqax23rowV/By2tiXWIxVVad2+JDQEc0YVaLOaoE7YXdwq
p875/4NI36KBJ5UITBUEx057nV4rDGPzYkOvLjNY2DyfzpWAYNo7EJOj2H479f94
yd0Y2XDejaQmMnmMiCRKpwbt7vxlxewcO/+INT5ycI+ysPz4QodTVqBvIesK0Rni
9jxDrsZ9hhMPR2WKU8ztH7ZPlEj7+RGYPlMXbgQL3X/wjwf/3xqrSTuu+qE6kUou
Jde5lsCYApd5pbKziFXIxAoGB0Cf9fE2Sj88dm3ZsygxkkGtsHeqOjHhfSZYS0ei
3SHwiSXEuEMEiGrUqv8T8Sq2W054MStWYL6MLukhfr+Tid8yFFGtmYxjo8HWDqzO
C/66CCk92OGt0z3MubWglqqXXNc6GYX5C7BXMHOnsQqgfWHN0fy6+ux1L4ThKsEm
oYO4WOdQZ1gJLPoYP0qHxzsE5zToUOFCNyeTma6RdEyuY6dj92l5bAyAco0gaaLv
uKYNcaFUt01trgZnhN5sCnZmNPcSdQB4xfL5kaGEkK8ffIzjHTrxeFL66kgxIlyQ
7032SVhebPsAuVsAbHon8ujqPG7jZ730AVaHuyk++5TN46Kwv+0nIxOpb8xUmefC
lqV0G0ZtjFEWLQ9Jnlo+OQtMewf0TqKSkGPKvk4jbUGOypHBFuhMZ/ZTDiUbCPTo
J8YR6SGqTaKW5mHKo0/0N4xVp+QVDiyiM/D+At/BAwCxJuKCsFCtd+Noa1BSobBB
shdh2iV5UPlMlCPPh0TVc3T7nzh0fCm5zD45e/TFbiVwCwKoz9NPQ4rfLq7oqsSS
elWYsD2PNKD3I+imXoImypi63asSzbjsixUGVPF77Mpk5ynV648BchYfW4v99zk+
`protect END_PROTECTED
