`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5cRlY0OcpjYJWPE12J0o94E7Rc1rIxnPls81jHcQRbP9ElK8zXbXrgfqfZdOY02z
NKHQSZTt4ViuaT3kJDpp+3LezhxCANJwImDaY1WPr3wEeXm+iFSlH93qvqt0oEIZ
cGUv7vrTm2ZtZpajXWvo+bP/WlhDQvoRJfz/8k5/MlVy8EBAZd8aht1lkEv3UemA
0DFP9NpGlRhWGrTdrz9qLKdQWDZQpfIXM830ThOGgYxBriN/jCxykGtcpiLDaDKJ
B43D0Ybf6F+fgQlPvaIVFlMQ76bg5w0pAiH1bVpK3au2PUcpiQwNFGSTX7Yb9MiL
fosVq9d4lMAQ0c2fR7rgy3pwbIah/T9wcNbkdM5Su/pvJ+PoF/mUhAI+fPkExpjP
Zc1fKdrTtdGpQv/bg1Rtq5yRFY6Sa1b+oKg1YIrYfVZU41kLcceB41GvaZwaiYIa
J4fMH7mPzvm+SHqVGkjLae3ab83q24eUCT2S7vDb+xGibmLvWA3Bswnrr2a6xdf0
bQxOPpHpJihv4mvEUCoi2u1c3OTKAv8HzuVbqCDYdQJ2cO6TEd/wFSso9QN8I1xZ
JHVIYhWzYFvZRXxAeqQhYmv1mZYoaUkBLdy+SSdr/zcJbcyptqa5hDfxwRgFIwYm
k+iaM+brsENMe18EP9LKvG51aa8Uucx2YvPqIdJSIfTYcctijX9jSdYOY3X6bCvq
Aw8THCYHiPAuMz+e1mRyiubVV/mgKzOKN9ibn6cw7efCCimvtBFopXYeP3tTcAd3
sJfBRpwxKBBtlFVUrBRGet1sLGe0FcgJqTxwSxpCTggm8DLlY5N7DR49CBcMwYRq
O/Qsdwn44qpKEb09p2z7SM4QdKa4UTTJLyeA2LOAQ+pQoXFYtXQuqRSoQyd14uq0
CGMZ1uEOSsQg0FXd6UrmbX5ccXeH7iS//lWrKr8zb4g7sOU5ka4FXpJEMxmsd2/t
1+WPQ3lKPf3XtwtCbLAE2qO6GzUcYoTdtOro+lRuaTsj2YAg9Fzr7ITK1Ezhn9KT
eoPw+EgJnG398wlv3xdx7mX/ZtX9x7T2cJUSCvRJqhH2/0c9jY8zNR+CXCNM2R7+
irSoegUvmxeulGMnJL+E2e3wqJjFWq6bw0RXU9F7zN5gFa/ihRC6fkN3jOAWsndo
HO/H68Zef2QoLRKLbLwJtsTJJBxR/orJWyMesl6ebecWBRjM1apMjf8NyKVluwII
G2B+75qqO8mczJ4yYwR+XIm+gLKYvV0JPyr2bTGQXqFyFGAqwZLFNCInzqI1GJ8r
hF+N5nCcZkYQtrP5Yb1EjPtTrOrmBvAjg0guF4WrVpHt1Y+sSoWXmV3aO8cDFIXM
SU/9+Bvj2fLhF2Po11hVr/GXSh3J+HnQlH8sDlH/5zq3vcW71moyCL7rA8T9pxwW
IgaZuMirCXhEkdkgsPFiH1s5iynS009hYG4ow62a6NCMoHg5tG/Jxpdkt9TL8yP8
kdCa5ZQuuMc4MGYILAUaD5qnOBSRRqNKXqF98KgwcwkBY72yPgc6TNKbLnyDkN02
3wo7xS8jly7b/tadwzzc/Ki0cQj+FJ84vvPC8flVY7P7XrFjlZV0WZvWaQgDpmW5
pZr5uvOrVt46CSJSjStAAh7vNS9GM5g0+BYOytuhWxufF4D7YFjWB7hlNBRUHqdn
0gXHXEtuKwKnIPUjOGQ+eGNKk5naoqEieHG9t9OQjmMbiT0JkpuhDKW1AsEYnSBU
7pnPcHDX5Xu11/S0mTm0XHNk+02Mm6/0I27IJgJheDUzafzuSMxzwRrmcsiMakKR
LZ+cuM5sgNkDkvfVveRUoKzWm4rQPrKpnBOvebTHmIs0s7M01zzkDD6ucvRWIywn
KdRhQ0lYstBlIZYWHNMyNdkKeLGjuZKBX7/eRpEYFN5JyaGsQzkrZWT+iyoyX39k
g5nduITP0PWzwj6udUpUY0Y3EiymZ/3jn1ddiBDa2v2vgEPt7gryH2Y5UF7ahCle
Xwdv4GzWTVLB14etAT3bIYz5ISRxMBv6xUgjM9ugrlTxnHOdXZlcmD/Qdf3zVWHl
PtLylfqsmZbxnawk3+IE0w==
`protect END_PROTECTED
