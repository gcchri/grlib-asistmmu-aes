`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZsZqR1ADx/5Tky/Bzt67ql6R3BrXtMoBTJpK6hqzVlwHKPiuLCmfdD+kyK+cGVS6
sK19frUdOVVgGRXF4tYvLldMiCdpf9PhHUtpksvXr6Fku9Gik7AjWsfShnT9wi/a
r8egatdBw8trORJAcJYI2fLBQDyUGw9/+YKSttbl7Smw3ZfHVF6nPx0YUVXN2M29
rslI6zBSXBmm6I7aQR6reqqrFSHNhkSmUiIm/nC9nZbEL8n6VaHCU7NsC4kumacq
+p8DRRsfRtmM8OCKmguVsAVLp9VW3piNZqKKZ3KhDI2dF4aa8M1IS8ZI2G4VoIGn
HFU5nlyKPvMEd+glpnXg04bwI/PSwU5sKzMKmsHoIE2HVueefProP43kF4n0Chj+
`protect END_PROTECTED
