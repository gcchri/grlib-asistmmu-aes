`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZJVN5iZLf+EOttrbhIQtEEn22tj/VUim97mnmrWDFlumWDLp27VyNzpS9EQ70OyC
7xl801e9YEkAVxeNYjpX8VNni6/ffiIHQTMxQVDHL/m66EMbT5zYswJYS+q48Hld
6GGOQp+YYBkaDK0WqNMRyBcEWxElgtYXOXapYEZPMDeKS7qRGH+KrC+8bofA5uNb
fdCcnx/Zx/K0e38HRpoCTh5PT9ISMViEvdAKGp2G/uOy2g+qdaZ/J+tAkBqTRPBE
wP5uMhumgKtkKpM+ftSblD53waICDY/2jYX6BuMN4KCqixBo/Sp9NQOsJEg3GOHU
upSEcvfhYay+hKFRoWi/rKcrrcPEGmmgxjfsWHWx5l7bXTAYzx6I69mfYiT0h7Wp
SGmFLqTdAl/Dn545cEkG2Cf7znVLg3DqBoepnPWFyHXHurrdNRFiNQvvMnrA7A+Z
Ps3w87wLttG54SngmfaAxwUeSPYOIfa2a79fCRkTm9KyqhTsYrNPCZLklaxg9yzq
r9200EHBbGNG7Fw/g7j+3VX8IMeTDsUdXnt5uEgQT7HKVw8H1DKTw9O55hDPfh64
iP1hBMJp9di+T1340deNRFJ+mwGVUpQZ5c5+W/QHsU8yhYzSOzRjr2dG3NXbl+LW
EyyGFdOMiQA2JOaGj0S6IA==
`protect END_PROTECTED
