`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pCZUHzoiP8JGZn8+WqNvTHkH4OF1qB5x6khR0lvjwf9JHMW4Xaat2eskqCh3C7SR
kmIP92zvsqTqfkEI6xnfDTkDdhDamUuMWB0OaSSW7xZlT/jhT1hOmLAY29V28BZ3
zCTikvOs7q/nzvOYJKVuptgQc+jccv1rihaykT1eO2PR/lN/AfDg/JtPUi3vyarN
yQPsUCxqQOuSQNWfruUjAf6I/rGrJO/vCjshYQbw4PYTBtYN7fJrH930pkiPw582
ZmoI5FLKHSozJG0TQE0anA==
`protect END_PROTECTED
