`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2aIxpIiyy0oXvjfrTJ1z1AeEhHpRi8R1k6pQPk+jGxOZHXwDG1Zvh76GxDfFZiwl
Sd806oCskd7lHR7iJnOQu7WmcLUh9PT5zIn4pk7r/0VixFWQUR0d4aaZcpVnSR4t
zLFgzKgLdhV1m/3On8/rXtQ73jXTZ8jmyqlr6H5hfM/PvxT9siUZy2kReXcEA+Fv
4V0uSHuHsre6PqUZh31UnQ2vuWiGis/IDbJ9hso0uZTwwhk1r6B8wOUaRz02V7Si
G8e6NPrH+lIgSZ9wW42kgfzoPkqaH3gbEOTeoomvVP2YZsMtut2MKWwMOFOnOgW/
/DL+Q3/l+Dp4yJOk3zfHkiJfUUlWzxinOLD7D5QIzaQ=
`protect END_PROTECTED
