`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PmN46frbzMVvWarC+lo2w6zJ7bOzXWML65o8rUCLCbIczwwU3NQckOMgPE2gsYcz
uemJdJx20SanPQQEGbNyTxKKs6SzNJvS6SDLw4+jVhG2pt1MtIIhSX2v0xPS8mea
MrJP7rdW0nl3U87/xNfcY2T9Fab5fUj9Sbo6hbF2PvzoVu3/Q/bX7xPHbs4YroPY
fZutm0WQbeRVwx/oCK31AKMlFtybp1/ToxSEoTPknVPFfiPKftgAzGgFxaS97DpM
0h7zk7afrSYzxmy66ehYuQ==
`protect END_PROTECTED
