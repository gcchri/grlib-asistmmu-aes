`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gyNDo4RjG4zzsaSgS28lnK8QYFVt9jFKaQ807Z6z4ba9BIVjkQ5JfzneuXNACfhL
fBsl1pY5DHzFNJnGTy+hfgUa01RLJ+/KaCvuO9AOHlgr0IGV9zVKvLIUolUkltk/
EHsux1Va1JMHfOENdU2NYyMHEZBym6dZ6KrrzilEOs1bbdkfffoVH4q+otIudDKZ
vCxte/2+dnGCsTbZQW7igGkrBFvNY1HXLi7w3vy090V6oLUfpRwtqJBnF8KayVlr
2GC+Hzu5NOmARNBVvku/ZRa1VIlOimmKrjuRVJK//rAEWduSa6OEzospssjxYvh8
ROOYY7zkQjb9J5G/7kJngAMlAMjIwBeo2nlsOUuv62mV8Y0a9mbQoMttzsLn2Or2
p27G1uRPwYIOtBgv4PhAEH/Q1hWa7wvc2HeWDlNZmYeERly0wuCyNNiqX/St4Bag
PuhnfyMN/GV99AJeKGdTqmdcn2JWroe8JyKSCoA/GNxXLlxoIIwRDyaoyWABYt5V
IqwGbUS7m32/KfJGSxxRYtoURYgpRKLlgRw8hBHuljGv4TiMTeB9uqGsj9zli6w7
an2oqAqCKaJpt/XoNqMmsibKIbykYxVg9xNiXlJ3JvUmSSPZOdjCTDmZxWiflFuc
QTsQG0yMibD4tptX47qNXBg5Gf4TCEkQmBmFx4tij48PJqpESl7ZYhXCLMw7P8mt
GNk3aFMduc2tv4Z20JPRk40kpSkXZgbDYAOm+M+zrexBCJNZDLVsQmEEp74t1Hrc
W3BOFP5VrcGbgGahxIME2vUrc4xCWTdavGXek5QtYb4aApOQ1fhcEXdA4tpory5E
ZuoCgfw9VQ7eI8wCsAb1htEIfjkzy8Ha7K1wvzDxceMEnEzFBHZt7TYsa584Yqyq
gw5licLJ8pDwv9ZF1GGUZ5hjfWe+6UecsG27prElBQpAsnksAK6E7T5VrmpRPWC/
vT6Pr6argAmssTj5o1BPxbM2PYff0SbfHGIfHAXxS/oIz+Wnlj99ul0vElbIArbd
YuB+xvnz+drTdWYJPsCv5iZvtjV/uzSwGs4eV5A3SreDTkG9mOdPPHzdrjBR36bN
0Nv/XCbPTTnCpykyAUJqCLKx895rTs84YEETO5HiU6HyuMQw0eI26yLg5UXrpgNb
TsGVC/9fYHzQEbJ/dvDidcRsnWhq45Nsp1E1qP0ym8767YQg9PPeYXnflF+mWOjd
o4HeoR7rFV6iSdDBmrDvPTVegUkkfEcD4Er8Pnm2MnE=
`protect END_PROTECTED
