`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c7v2dNuobjKsfP2LrlRp/CZCWfbNNlzJ8bnKcAVWhCKNaMNSX2u3Ryaeoz88Isy5
ajaeo3NtuY01mhdQlSkKuW8VFdq7TjLKwsqZkjamT4CF9sS9RV10LOQJ3SHliAwf
wYiTGM6yASHWbk3HyC6bl8pwqTEyDaTB4+X1ecpsNEPlhAQE6y2ZdWhO16LBsooS
Ii5oupqOCwK9gFEBEZiuoqeQqkL/Fvr5QA298mbJDaPmPdNBnyoWCFH7QSac9UEP
b+TRYqRzbS5/EL1ceLDBwkzidGWHWEpkoXGNNSyBkhe2TorBJ+7U5BBbqF4bvk6S
p0g1af0HfZrEZknnsqYV+o4t4K9roACbsbbDkU7ejJgAcNfKXtevwzxH+2yp7fgt
4iMTG6eO5jJx1dbTKkoZzxxTu/2FZApSDWPgCvKv0ZU5zUcKl9dFUwavUem6tuqz
QHrLUcRkPcTwjvygznnlDJdC62w75odD3Xu6kyOMm7b6jRJ69J2FRz48shQ1ditC
W98jEELRg7wzOlnIXbW+aXn1CJBlnXIvE/+F0ylyGRmK6J12beBXBOXi9NDwZj1f
/jsipnorVahL23LhndS6O+LIE/Z2Ioj2nuoHgAoL6QFVVCQcPwAy1oeFQDyB2IoK
fbYLOcNYXGg7d3DDI/4nlA==
`protect END_PROTECTED
