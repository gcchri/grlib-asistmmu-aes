`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7wKRS3mrEVz70wx/qq+tSBjEfXID89zNZbqcmX/7xwTOYi6jNvPkY382j14M18uu
ryAL9vi48fLMD+W9U6Q7yhKJ+CFhDgX1L3kvgLP6XVr9+Cc1BviIoSsJAkaq+sY0
54lsrcwB1YBQ2wcT5PGvxWlceIy98d4pa5Jo4Jc3iW/t1epZ/CPUE8WLTfzqlkNL
mtTId+fQXF4Hl8pg9bQeA9GUbs7mzKKiTkS+bGbgyj4DpQDROqnL6RuHYxRxVWA9
d5nFXGPCO/OcIk3kgtjcng==
`protect END_PROTECTED
