`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tl5agVipsF78T1CS0w9ElhcdvGkT1Md2m/1PHv8ELFbt4CSB23unHVNoR2EnAfse
lVMfBG856qgnNk7/DrabmtVL0sdzxWKIG10WB949psX8xSAYSv1oMeCA21rqdPle
radHFpVFwcaipjmOiEQIcimgG/+x13rSMXDj4H9P9jx8PLg18IQj03vnMUEBqa6z
gwHot9i1qQGuz2RCz9e6efVFm/oxAuNm2nA9pQtww5ANwRDtfMxygmLGf5x2OcYF
FsE1HOqbP8Cl0oE1mgO0IJT7ajF1N/zSFXpRKHjZqe/AmPyN4NklIeShxC6VLky/
K4QUSZ7PC8xnP8eWPKpbtg==
`protect END_PROTECTED
