`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
63Andb+dUFgv067+XEbfMkkvRVLSCcgVjo2Tl7rZkQfURtCWxgistpYqocrPzrrd
hO2gMm4toSYp/5G2AgyM4vbrCfo6xrLZRUYtZKhkMUp9DOvjosTCzjHHCtQd5OTq
ht1t2uLgtRsS9RU53LgM08q1wXypGyEyNWV8JyS6AuIp9CyQJpvNIbY4bTIXsM4q
sj0xKJ2aZ1417Hyy5TO7YdSxJL4lKGVJIubpr21zMYFW2R+DlxJlDWfuM5cmkSJ2
6hiTAwNRJ9kCEB6QCygDLTvx8tf3cN+99Qvi8ZE3Xm4+MiaeMo2rOFigyTHCjMWT
zJMvbLMAqZQCzaBJbVAL12ApeDPc/b05NVsK/eA424TrgaCyQMv1P0UO+SpIWTt+
`protect END_PROTECTED
