`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0We3e6qv9xCMXfNlQidiF2QCBQnMSq3RjRUpCJVWzlemT48Z18HXMqHcWDe67kOt
ol5uDcOekOAqie0eX8KUoflJD28PIAWbSPMquFW/Q+dmjEjaQpCFKd56lftHWX6E
06lzfyw4lriBWw4P0kaoRe0vLuBmsmrHJZzMT7xCxbcGNcAS69a/NTDOjd+a8U9I
fycYzhPYpOcqrSr6pbSwSmYggTQNEmlc2rmRnSmplRaW8O789L2tkhAObqDp9wFI
jPvQgci3oYBtgCGTN6mnqy9KH39Gp8rkyLH8X0zUMP0btGVPOgHDiu0yRpoYGB77
F8ylmvhH3bfMb9gd+DhiAwOaMFTIhXCBqRW0H2bEhHLEfCGWwHSqaT1mj8Q9+hZm
SrvvA7U9x8JGZQxPdZVHZAGpLNUSB12m++bASEm+Ie6beOcVr/M7MG6SPXjePE+P
Ce8VmjpIlb8kxjNAX/3QrqsWSQPa040V7d40P1ec4dznvI4ZsBFJJ2/Nnn9Qclxt
SejALQ13KpCR2f9lLpzoGNSxXDoqqwWHSI94XpbzFQx1nU0aV9wfUxmJAeQDwYTi
pGYytwn0koEFU00JKf2JVQxlolIXE3WO/NdXpJrGlCgNeSgLxgvXAe6IFcuCoAAX
oo3kfItFTXypzcpDxVxtRPaMgk6vu38Gh17UxDIGFuQU+xDQ5AcSkVVVJblR7ln7
e7k+Pz5K8yaOLA3pZYcgnIkQSYCtvMPsUxpOgE/EdtCgTaZzBUQJdvhFTnnVzULW
ewLw4Dc9vKQs3DsgDBXRyfD6HVaw/kUG+LMcm+R3q7iO8Nm1wjAzoXF+uy3sd8yb
OM14sP9Mvc0c2mxpuDb0hargqb1zACl/hf/LTVZRkUgYCOcedojpGId93b0W6Ety
Fdqkgwu1rIjvx3MfE8MsdEdv/XxDVbIDfEV7a9xgJxMR/abvOgkMWykspomBDnH9
DelC1EBBMjkyppWPJHsHbpk9xjW48P2qnexFrSSRR3pmSrUD+dOlfc+KQ7fOe0Iw
6RFAnbKUyunubBt6Wn90n6Xk+QurSFt4Yrw84EOXeeSfUYEixgGHuvLcGfrdP/CM
CnUx5CxFomMMmPKc7TxY2Da5gsEx7w2PcW4k89TBTE4LNbgqrFBgNADDns3v3+IH
bpa5BZJTdOkg2wjE9wHfDSjGJpyNmRpXhplANJnQwyxflU1MMaJ13ExTBchJTT5Q
HSsn/u/ISEPCsJny0BuWcrdMSdrYh5qDjxnJQn0PG/54lApdlGyfkcGNYAVOuCv5
I3UnDYbyR6H4W+5zOZ/1CQnvPsrG7/EIFHqgxI8g8yooYTXukArDwq7+IRY9LlFp
l47opqYTWQAJOStjPdvoR1h2ZRYh/IHoT3DAoRDaD5WkvUskvpcfwHYAiinmnQkt
R360rU2KzsE/q9GnCcBp0GZn37swMdfbR1weYcDfARSb9HlfgVmlcocEyiSMrB98
+JIzixmDQvz0zgnK23oL6/O6mDZj3GA0I4WFg2fNd+O7s+TF7+xtTYYWZeOui3O4
mJzJK38B75EGfqUNbzsdwhe+AX8/THxUrduPvPZ1m3ddWpXPfLBGG0Qg32/Zb9g4
9T6F7yjrxBBshN9cRJXc8K+GA5PIhJ2FdTGKZDiuZtfJpgYfvlLUHzAeXgKWLIg4
Nk7aNZqVWMafd0ETxg0bn1bnS05NHcy7L8BTHJfLGv7bvkTYmtiyxMNXZep/G6ye
0MftS19K9b+SUlV2MvhrHJpisVaFHfsIZ8LQMwrw2av8XqS6cUwNcgcTUF4klTsF
neTyd4SlTmTY3ZVp4tDzCO09sYTdgTFC514lnSe6cjvDce8IiYBSF0ECalSaTKVK
`protect END_PROTECTED
