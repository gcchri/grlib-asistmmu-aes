`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3a5CxM2VMWiYvzC3UXDgijemSmB1QoiL2HnpZRPFLVG8cu08/bjhvsUEuARrJAQQ
tVc/FnFUZbA7BlKgqqWI9ZP1fDn0VDl4TRGOM7k9iYZ6cU+f819h5rs9SPO2VCWh
nkQmxr4lqgIGoAQQd0sFA5KvXDFgIFiq8YzLY/lRKGWf4PDAjGBQr2xG4O7mVRRK
E8W00e9Nl/91kU13YbsV5P8AKmXRAsXiLMoBGXa16wusAuGebLuu1ram+8SgLyDy
KGfEjm5Ep2xpw8O1FuFE7819RoSXH70ZyBt5BGlg30XagTZHKILsVe5gtuKzDlGd
9TKWNx2TAAatpYamdy7ayYCEmM1xbJf/5MdT/vbSQ6zpm4MKo2uyM/T4Q/+ShZ1G
+6qm4wI1Ooxat9joKV/e/kswyOYSFlbz2TS4QcU89DisVDLM20TtlFo5MpUYSWNA
c0edvfOEw4LSpeDlTJ8JcZU7vN+kny2n/DKBfGYAaOrffVRpwv5vjTKZr1mauA6C
uztihvabMG9k26943X25tVx4HYGlyEzK1YKiuZhnZhwhxvSKelhQ3nek0KtTwPqW
xlc/8yPzBlcrgDVewEDU/N/0NyjRjPlomtfNL5BHV2Yx6cnKK7aKhUs/3ley7lXf
UtWYdt2F4mKEG1PmBbrEgRJx893ayLP3O/W9b0yLyKi5ysIAbLTgp72tNIZOTopZ
hRzLBTF+pearcnIuLUvif1ulwsyCl6oOxhkh6k5lyo1giLQsYJOmRENHgqFSXYPo
n7U0U/fUMx0+mFozFv6MdF0BP+MiZCZSBk8tuHz+x6gnxBPe5e5BFAb1mmwLf5OX
xK/4opHsMKENarP2A3Lnuan/b5vivb15BegRwp7mHF7GerGNlwGjVyNpqpX/vhUE
I560EsJaJ9KzUI/rnQyspJDOmUut6JNl4WMc2I0i+H06qI6oNxi0AvoqzVR6AsIG
du1r3WeM2PY8GDOO0gwWqHpmBWegoVOkQJr7T6gCqVbkmlsm3TnCUkIrXYcOvNHE
mixXJl8uY6J/dqTKJ/HH0qXImCnwEw5eriuKdZLVYIAdha1gdayuUn1z1IxoZQ8M
BcXay0j6IeafH1cddaLZvQZeviPBTuRJG9Kc2Kmrpa78AjTi358qcNuhIAAAqxgN
EHuW+CWqyA/XT38rMm70khWMxy6ChMemzdjgmz+vRIK9P1F8TfKckjh7QAVuawep
n8kib5cPUSc+gvi5GXD0C+JlC/xe55/2wfTs4kmCf/8YJmWw7jZuRxpE7hRfTgL3
LFIMV9KKAYQaOIqOD5wvivmlLugHSvkhxbnfMXVBCE2Rq2g9d6RoLYMLJkAWGZBO
egF4g8+LDQ1S463UN/+TCo5xyrpdruocRKON0FSEkpe90zdFoNU+H3jDda+SL7Jl
iJs8F+vuH4M2awoONEgQs3czzjbdQAuJ4DRkEfkOekYRkgJaywAQeWkvplaA7/mh
xy7evZz2EhHAyl3DiHESc7f32OcrbpI2FkSKJN/XmbKQd3XmMMN58LJAlIfDNO/N
gKDN+o1hulV86gDfRR+CAK6Ao2f5FwE1eC5puw7Pd9Hw4+ilkXAWx53jhfaAU4+R
wtnr1s7ZLmvBExn/PAG1s6UCEWmeiJPV1iVY+kF+VbzifHfGy7Rk3jLj9gOSMDsq
cpl3/CsaU+PdximwTVAz8nXsHYjIIkwnOoE5Wh9ysGjZ4ncqGwG+gPYXsc+y0NDh
SX544cd+BCAxzgGPdvjdXoS2MX6Lz1FGTPgoNR2NoeuP9V0j7aP9tusx3kB0zVNq
OfjmJrL0z7v/XtyBGz1P/zp1JwFpZ2vWT+5j3hEi+FCWCm9pP3uo3KNgvF06vACV
ZEkP9/EfoY+FApUNjczo+yMJv9UmkOZT24yxeChZrz9ZQ2mYG59OuoUV2hdo8twL
WBBPfrTBx646Xftsq5o5QwFpJcqdf2FbRw74AKcnZBLLob8WtPLpYFAbj2UWf2FQ
5oDS9Z6expBLtRb1RfW7BniA7CqFytfoTP1lcYvO7Y3oSPcZiah26Qbd8Bw8MErf
CYO2lo0qcI3BRhcLrY8ZCtOgMesbQXAtkoHI48/vufXF1Ew4SYj5k0qWAfdEjYP3
uBAyuTVmaHV2fWojFNJhyBmVpG2MwhYjf8mHjUbJUU5TCM6mnmcwthDkD6AK1JKt
fM2lTOweKqvPFSZtjXy7kDNFd1OItBUs0olO2hEAxMkYqNr+ve2dT/z30eY0h+pA
7knXdrtos9uz1yOxXP3XPSElCvZKNhslDlUsCeRPSQs1pOL/4b65pYQqdtM7SSHU
tUGbkN7PIe1drSDa8o1jZWwaU/acRTPbNRk5oy+EdrBmjxKJb+B71Wwpvlsgudm4
gOZU7E2811xhSxB5n+1u2s5f//yQ7Z3+w0Q7r6ejrjWQoTp5I0cegdeeG4d/gfDW
DW0vnvl+MxQ6tcf++KKnztUG/1sOpJLH34yrG8T6VPPMzDC9goyD59agDqbE+9cl
0khEZdaNcI3le9INPY3Sr3juryezjAQhCTgwG4hi9aVb0mdI2euhCkvpIkzRWbH0
b/j5Ee01gsJZFbnSpVF56KwvofXc6U1La8/Gz6rX3mrrJpwMbQcMTGLWTiAhZos1
5G0imGwA8CWtMjSnx+efhRdvrh2K8zv6DFAFR/52Hl8v2erZegT+FtnV0Ut7Jedm
xDx4xBi79QT1USxy0dFYqU8PFJRQyHkbKqOv5Gxh2SQxQ/rqia2xi15yGuaVSsVt
KxesWF6E0/efl5Vm9msJHMRJWPaVoobJpH7yGrb6lis/gpxlgH3kw/REY4QtqpK3
`protect END_PROTECTED
