`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LpTPFMOrzFnQHwRQ1QxOUHs1Jhbfy6wLHeLWIhkcRSo7c/ZMr9zDqqasHXd3YKX8
7ie3f4W5Y96COOMQBXKTLDH3HLHh/BViRNYv0d5nLnm0knZnCAIy1mOJ919GWUwg
JxE2d1Be30v3lZHNwhmrhKs9RYR9RUspwJwlCNPiFQejooSlaLyC1DFtfVwZUr/P
bHQx9bl8bfnXuY72fH588txpS3qcQvi91kD2N0gdWgfcTajFcyXcYUHabvofbPe8
OyvwVP+/ao5A1tFyrwBz0HUh7ORLaZEmNRsoss6gNMQq4ac97ShxWJF8u9N2Z6V4
lJ62lVTIICKmuHaKohj0PWqwb/kLCKnfOoXOeTlipEeshPL5tY/1589/R0HdTn8T
rT3LVGk3LT+TRVYevj3eVRSgLXWbITnTr8QpbkxOmrzQ9VfqDfA+oNoDDMT6JRBD
3XOEBgcdEZtd3i9in1zOVD7BjOJROiajY+Zt79aMb1I001KfCHdNYK81a2CRC/zV
3bXP0BSX+jgf47qqGHghJ7dec1dzruXbLKoHSMB2wtuPKkAqYyYjoMKr7u+iDbVV
g2TSV1WEMTImB1dahda1KxeXdh1jCq2gvmA5zeoMFYTjv403kShKKs5syg4VbrIH
lZLMhdzFiDLVyfX28ggDmvVxncWkvx3Q0tg6lhSCvrd1MynZr2IFPD2/WkkP5X/d
bNsSL+N+ngzGWNhyVErYf3g8ISJSjLenlG1hF1LxcFbwW8Wqun8HyRGDHUzIS8uY
dI+RZlifBfcNyXciQn4FoQ==
`protect END_PROTECTED
