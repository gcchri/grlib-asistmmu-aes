`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yyLhDTOnYLVfqZqmE32tTlqVwbtCirW7u6cGMBGg8lEJxyYYnaUeymEd0/d3vYbi
lu0RhwMsWfcUn6u2NJzRrC3Pxg5TmvTgVi+MFqzwUkGGmzssmTv+tkQPsm47fTnR
9Qn+D5/wUcPnwZhUpEWWNxS6Xu8GZqqhNhMak/3gPxNkfTcMWF8FGBrPmSmJvLzX
awouC3wjep1FPyB1u/dCcJplNesl8pHsK/cu1pWMNvAE9ejnOLStgYdzYsj+T7qj
5rOJ0hVl0elvxdxY7YhaIXhR+GbF+IuQY29hhcZxC0oiA7ydODR8GWUkIjwV6EWr
XAKafPGm8ltziuiGok68HFJCIHIZkvzspa+qMPnupKnes7ZIu+UkqMt2Ho7ZFNyh
L39GkNkRDGu0OMdiiIoBy+hnsVfkxSA8p2stFImuVihq0tgiUnUfQfTgahJzxDRn
/H/d+HO5b6xamUCnM2VUTQkn/JsvVRNyKuxDKkbB0Zhyb5otRl5bsFTo3zpATfq4
KGT2adzsPDpyYnHW305TlxeTCr4/omNZwU6ABEHq9+ALDFl/egxD6BAsEyvRBLqz
hQTqMQhIT/xwqni7/sRlg95ulyLQEZzwM7/VT8zeoTpVveAj/209q4Xu8/87Iv1J
p/Psql8BJWd14WVuAq7jQvP12XnHGIJ7z1OAIJsrJ5WClhqQTvDHB+rQLyRJn+bG
YZW/wHms4fFrqvZb26fFPT1kXbR/a8lwZWOsRU1GjcdRGHpW8vfh064iFpusKfsj
rKezUO1n2bZhd/4lkPS2nJkYCy0E2RT4UsVpP6cH0nOm8PBRgVrw5j/lVzMityGE
GUcnc/XHWsjI/wHHk/r1BHR6tsZOWhLWxX/a6uSKeqxhY1n13djsnlrcSdNp+WWr
1NxeVYlXTis87NzirwWnoqutPxdcg+gs4/Oy4aGhBrDDpCfH4PyqvGM8UGBlOZtA
sIYFBxTbHPlwRzt/Pgck2tFBwESJmioI4mDYwDrliIfFq3+sZmpOOFil9+DpGO1v
PvI7Kb0S8t2/jsIVn6nVGDkkvn3VZj8jUxxUAKUKiu8bQFjWcb+g9raG1VgOZlXx
TD8rpVlyYnKcf02cxi42k3Sjqs+Hq4JYZKsLLSUiOfxZQ67qqJC9TNMDh37Pt6gb
17KGheKWZs5cafqefz0tV/j5TtTxfzIVc9nYCsnwvSKVbZpTNOgD2iOuuPGduIZp
XIIjGfFJCgb6OxWqup9+oeXFHvNPokueO7I+m1/5duzMwgdMS/AK4bIOY9XYCees
ZUHgjG00jXbD15inpdZFyEIJyty68ZzJh0Y03dSGnft0/8S9aGDWjZm2PKYkVL17
4JKpNZyKo2cgla6KQ2hmz2ksd+q9CZmmYMuWAxeYZxuHeAHz4R4YRG0bWCEHulJs
LcA0jt2GBwjfGgYMtkvJqEhXQnP58sSlTJBrg9iBcU5ZAVKlqys7TWx2Dg4r3Ges
A5ffQesz47kkZwB84YEvbwihKTolrpXsDvnpQ/vaOl+QkqOKnXTM/PIOuZTilQdE
y4YmlQAhC6bZjIfoNWPVCjBPmoXZARQvs36zroTiHncGhLvdRZx1VnOy1veQgyx6
Blj49kBVE+rdmSkdzCunsDKljl9HwCz5gN+dwOr9c2M=
`protect END_PROTECTED
