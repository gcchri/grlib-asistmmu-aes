`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nlCeFq6GATa4A84mNCtPveDhSO7sHH/BQsDSseXhs3V6ZO/8318pEAOQ8xdXlL0p
Z3/RVdq1ok6Qlnr2h3m+dcQYVjIPYxRDZ2NZrj1LSYmnnqI6dHgWj42ArkabvR5S
7H3vg2+Q/9CDBSjByQvHq3q85vFLVPtd9HQ3XUw5e0VAR8+d7Q+Gx+U6VRymb9X/
o0kOK26njMvZDVv5rbqvLfVfF3iliAn2oHxFYSx57nu11uPyAEDESgSOYQEj8mY1
Mq28w8HeQuqRw7vLEjDLXB9MrTwfHp+IfhYbXKKATA7nPyoZ9PWlisHNx0OZQLCq
Cv/adSQ97RP3r/MnQxVWDtQkujReViHUtmyVM2g2k00nZKlpdOiyX07ZNjRclUx8
eurdb+4+XoPb/nPRJN7SioI09S8Q75hNTqDSTFqz2ym9s18fBBa8Vyyi4a3LapBj
w/MZAfDM4i/GtNoKfPD/ONYOf7o+6SoQ8t8Rj2h2GQ9XYG4s+/mEcjGxRkpe+8pk
fHwG678ygx1gELThTQGSde9s4SZi3wTkNBVupTTN3INuRT6sNk8aHUYr7Qnd4dCA
Ei9t908Vpb+cVB8tYQCbM/DLtKV+A6Jx+aiO1NutibHWtag6SSRyK9dkIeCgT04c
chmnnA5GNpx7+/FLurrMMbeA/hbDnqM3nD0I0eazVvnOmvHBF6AG5UJ1P7uVrHko
MhQ4b9SDhyNZuo1ULniWf9/MFcRaQnFuZ4rkud00ygzwGr8f4z1wvW+s6JiI9O2V
AJ+JW1vjtSJ3+tWNCOwkR6QmkYdqJfhHPanEK3lHqNejbijhm27w1IvsHy/I9BDV
`protect END_PROTECTED
