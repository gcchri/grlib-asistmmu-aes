`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
heYBSH/+LwxMXuWD52ZaKnFd70/FROi8Dzw4AB4AbKcElPErX8OYOzyvH6l+5jm5
b7RBorcdFFGE7rZrsgtLbWCk7b+6lwr64XTh8KypbXR9BNbHigdg3z/jeNlHRp9i
kq9E54tAy/orwFOkAQ/TCw067nKLNevMwzHjqaHpudJo3ijNuWG7n+mvUKWbnSxg
gRX2J7UdMw2lgAsWWWb5dYyysGtCr3D3Yyyfg/RFNSKPfpcOwn+S0VL/Pfovf8if
czNpwVUdE816Vr/oP96lhXPwGFZheCclTMTypgO89x5rVCF3pZRdvT7nwZtpzaSk
5xuCJ4pvDVvuJpyZcQRtuxQdSt0JkVy3PN4OCvEtfow6vsQFqvOvsW9CkfIy+/ii
NgE5nBkSnRgN3a2bCZ+ftdU62rMiOmP8QbOz+i6oWVK80yUd94ton/VALe16XPem
HRjvCTthMLVUgqwL3RufNmZPVfq7DunCvniiC5sMYKZat8YqjE3U6urWEwG4Yjfg
4FkCfiBvfO18x4xaJn5mbEmFth6Ywr+9FteKNW5G65py5vohmm0FIUKiYXM3OSkv
peOg++iSL6mqUIr2cY0HvKDmVT6ffK3eKeslC1HRD3isC7/N6jE4Z5TmDfSNnZ2R
o9q/Le3Lycy3V6zo/rMqN4XfWVAQ8Pmmvp9z828qjAAGczNYvBGGViyatexyRjSa
lBSA6Km9buZPwfBybX2nYUt29d1G4+Md3V8aKOOrEPrQxW8lLclj4RBYwPfwi/IK
0/5wvG0qkZEH0t3US+FpCw==
`protect END_PROTECTED
