`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FllxuoRc7DcQUE3hFgukEGo1IVVBIYjBK9lN0Z/kNiEIwDzmWSH9EdHH3BVtihbE
pT7PG5pH4sN+rnnFs20Hd6UqXMDOu5K1FybkSAG9DySYo0e00hiNzrqzUglJG6KI
Xikx/kI5vVAMk64AtXzNGtqQaM+WPBfEPfi540hO1hcDu1F5WxDulFIlq8RXpRIU
qLAWJwYQ4HAXAdrhQJ0Mlija2mrRvtnztK21ktOsfHhrobMEyy7tKnsYX6x+r8Ba
pbwWkvR2xn2kkX6nDnLDREMI6FlQ/nRd/0UjXWDd6OC7mJ58saY38ViC3x6d2Acs
HCfGo3lFS34jVO83uwzWPZgfhqN1hA7QB4yD33Z5aY1wwxUbL3IXeFvdEsZWaHAy
uDcUmQAYAZfJkP88LiTo+vsf4bFyBh1UV85Ett846Cs=
`protect END_PROTECTED
