`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
62qlLImcHy4XtcjcaOzLfO5MD4H7u+1GvOkBUa24eIq7gHP5XgN5ocaDq1LxiH6t
7t4rivYEafzTuICjLlJGvS+zILBERCQvNIoHochhxntph/BzNTyiMcCkflvPS8Rz
GzZ827dR/a7/0AHgW6FNO1uWlZ8RB1mfuKHlIaXZbPKkWKVkdH1wK8nchAZX+fdi
CggE0g2eZ5dygQJULxDD0l6dNOv/cE2+fLVmPMmAlZbm44/lXAKLM95kGotsOWJn
wm6ak0a38n2qt9yMJ8jurDy2Rxm40r1RQPF35GEO8LO0FpgNGq1y2mOA2JB5rCWp
p2+KT3AF97kv+seo9rkiJNCpq4rxYO2yBNVYYpuAuwtlxh0aU4CorHOPqJSdOk9z
`protect END_PROTECTED
