`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
53W4VdbekJVgWcrQEFWIJ77T2odynHhr/TODNODTQpLvufRkcgr2wCWOIIELcsjB
fnrXhum8GmeryuAHgXQ1Azafnhjm7AZ8a3BtJMQ1cWpMUx0RzcGiivlrGH6zOF+Q
uz7ASx3jHHBPYpr43Dy8fzwQJMn2jvaHJ4aocAvMazqtNRCjY+uWonbm2vhrxvWb
OEU+gm0/gcAWJIYYdZzEHBmUAyEbGZdxxUlLXabAaRCs1q1ygwxVp93DSSQlIQ2z
mdEf4AZgP89uLXFBVTrxVfzXCQ6iMJGVjA0PCJV60Q+WQmfPnSPNGRm65tjiaYyh
M6bcrJFbS3k9CtEXTLfMj6AKb99xQcpV1gm+G5pAp0Lu71sMk7kXUKATbd387/2p
3OJ92hnuAatpiEc1C1tPFh07oxjLANfi5POIcTyPQJfFYbjQxXxnEbjCXFn+AKzu
8xsNXyQR/vcuSZvFa/DIqTM5JlavNuGh5Frpy2Fp1gw4vyz6uzviQHNHQET4vaAS
HXvXacvGnOQb0GDNpYiJGHsAjJ6LOa64yYE+Mfv0VOTU8fcM8k5viYPi21t6YhLS
WrDmAxeIPX4Z1TTcYWaFNDkXWNMQGZh2cUmZS2gP77/75OzUGd/y270lm5IcKBI6
2k6ktYhzkJ7Lu5bPauFS3NBsFkybzhtYu45rlrs/wN2RDWUXw4MhOhzFYNRKcUwL
zcvgMTmTK/SNQc3KrrD1kKGdM0/8RBNo+eIsPnAUECTrNPU/B0ZwLfc8PDVSI5IO
RGJ9w8CQ0ox3qW1b0JLcHPnClkVOil2dO8NwCcc0Ryk9mgOfX4KG9GtVuBtMernZ
EPsXgOpLFaA2+dp9aqrsYKSBpNCr/owduPPzJfliw6+THxd0mbuRgPW2vTwoRed6
gP3Wdk0zjpdrVlEIYNNPlehhNznDC3uaI03HJ1TTEp4ie9U610O0/L0epMC8VQ5/
4/OkizHgPha7oZHsbWZPR0YcqZsu8zsx4xW2ZXG0shyrowOvw0x/ycNqjcxB1hii
vBuS+osGRQY3+YBPWzMFpi/3O6auoAQy2hZw92Y40swsXK/6MBZbitayIO10HXpx
J8KYuPeQRGXqY0D0PG3BnxOZq+A4gKeBQ8P1/5KSXd4WgnIOVoZ/klzDL4tyanp5
v1G6PXJmBdrKLBhA5tDttVuIu6W3h+nusSokYiD4bBPFD1QzAPlbvSfI5i+TVze+
050/DE4lTrDsESWrrnxjOpTcIf4fKlMu3oGZiGjCZlvoI0nct4iH0IIVpLOIOD9+
3QqbL13CZ3lOfv6NCUyMWhc4lGn7lbZweB9HHq1s4WJio5Cflmcr1s6OTG7CdF1N
uZVxnA0IghzqcPi7TDxcKyfLCXeT/bwq4yKCfY4qwBFkKqPGwEohU6PUl5xlfI8l
zsjG6aStXhRiqaDcaESi8zgXCAEwYgPr9XCmsmSs6qwLzjwnpWQ+raQiB/NMON12
0ECLO89V7c9hd6+XGDs3fW3rpb9XoF/QqvNNvAHiZdeAdWmRngswgB7Lz0fNwP5R
14NiKNTPS6rQ9P6OwlefPtErdbO3ZVnioK6BpRWmadg+2/5R3qjOw7yGv9sJHBR7
HDSzGGEG9GfLdyKrGwaGrRAlLSqrsed7gXBD5i0pdcFYbT2hoLEsZLhW8nfSPRjF
/hl3EIVT9MrYDDTFLBZUm/Ed3SadSwdXWM5AV17s1A8=
`protect END_PROTECTED
