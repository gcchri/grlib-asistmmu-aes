`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xeddku/ytJVbvhFXe8XUV9mFm7VjsvfLFrKR4EXV3jIli//B7y2nP4pFmy+xvHpW
ntl6mAzwP+2kL2pa7/5ho69E5z+U6gSO/y67t92kxWpL5Z8ignXIMaeKXWaYwz4D
WwTe32whPP/NV34MpeitFtUImojmaNwJIvjjolQgPAaeL5Uak6r7nEjsDY24oV20
iBTrwUYds8wY06J+VgeQ956i5Tv6iDSz32jc4Nrntbi7tudrsy5ZigSJWpwY8B7g
wv+vstrS52CCApd3n9RtEuIhaf8cDV1y3p4dx3YD3wrh6RmOl/XAMPU3HLw2p62H
Aqd+UPjC9rDNnW8OgYCzvX9i4etA9hwZfzNIFz98MgPia6t3vIAKQtUwqZqwA3+8
qwLILDC/CgHgfYsLuAGKpoVKvu2p9mmYHjyAfoPRTlE/2PXyg2ChjG3YdkiGJNow
64L/og3Eca+iTVQJ98GNnm6Q5fWB+nJWOlPQp3d0jD6iLM7cO216SIw3u67gB1hM
JTIk35blR0t3G38QpqlKs8/4sCG3tx9/gz0pCyPspAXMJxI8J2kpXo6bkyq0ueeY
QI3n1njngKMIol2TkDvKLs/ipL0WsSehakYvwHrNMKwDHGQw4y3tZzrzWaS8APbC
VO6JGsaUOZXnJY2e6U1QXQ==
`protect END_PROTECTED
