`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yrrYQP+7Vm4LW9IIUyp/+L/+vQAyAREWvLUlCQ3B+rxD1/pxKUiqJQdqwfIpb201
oktprn7XFZ1+DSAT+W6ZJlJa+wKWy6A7gzkj/Zf+u/YjozAuyNWR6tajaPz7kE+d
RiIgyUGRuzi+KTKIYeqRQfW39ZeL1GV6XtnwP9wZTXIIkVphMzlmraHPklAfrZON
Ec4GKZsOVHc2CZSKf4im7zYqUuwA2ukLoe+Ul+ftsE5CFvzfbhso9zgox941g+uO
0AIyJ0R6qba6WkmlUBqFcnUC3E/v4xlgui9ojNE0bNJbHtOdk46Fm7zAtG6fXRrn
0AOIkd2VjlBvNuCUwgylK8rsvSq+Sx+DRnJXgSQYN4zlzuJU2DoDWXDjyeQ7oqw/
Yh8fIyN+w7G4EueDMhCVtwyO6MLwhwZs70Z6c5h0kaM=
`protect END_PROTECTED
