`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sbr5uABqm/g8mzpeCAjMM//+3ZwRmeHVHn0GTCnwVOP0N6DTG18s0A7O/ZQKoZiT
7mB7xst2g0Z37xwDir592EE5cEC41Ia7PanGNkK/ovzs3ponEHl4HOt1UU75f/TB
UOo2zxWFOGBXsXIXbVoO7MFlIVVLk2HbP/yElbjTp/7VZVUgQuzRHkWJHTDNMpKY
o5g1BbHg1g7BZHVe2rqnVdezKUvNm9CYER/CgV/Pt5QaBJy8mamx2SUCrovdJPgQ
aQMl75QupoEqt5u0xlyvb5Xhbh9e6Ymjai4OeaHg9KrtUYB42MOitHTCT/gZ0Krv
`protect END_PROTECTED
