`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XZDgKUgT7rhtD9TrfhPVeFA5kXYPN3aBUV2NSINmAADk2XgASbP0uzKTVCNK6eBt
JH4nQScOCBySGle90upzX6tpfXdbdFMcWzckJjVSMeb1Ey6hcyrRFxGdyLbkqGzH
D0EEvt4cP2233dV9zjoBmfVLRDSGZS3l/Rg7+vipSXvkiLEPHfW6IxnvtPzqt8PM
a5ry8cE8acN+UiJL5M8mDcqG/X9iUmmDbLFadsIoLoikip1LbNHVoR5MUPFNdkHX
j18Qtso6IRar3GVesypmBWsyK0TVDOKeoYtQxgXcBtWkadIG/93VPONXQEdYXYvF
Kqp1crvDR3pjZJoW70SSM1dan6EcN93mNF8t/O71vMiVDUYT3BLdLNNtUiicRRrV
iovXzi23vU75/FRj42XxZ10Rt3WPq8dqUxQwDsB5oFwUy5oOnEiWkOZbzJvc3Qrl
amH5lkLq+xX8i/oW8RBEk3qoTqvhXt+p3qWVeufx9oOD45SrW/9Ak47bXLYcCTAd
`protect END_PROTECTED
