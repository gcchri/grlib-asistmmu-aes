`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
na/2eXYhEQlOoYQdeu9EAZ997Pt1FEfLlaKSFhdRmwsWkI/kpxlOoDQrQdkLg5DI
GL+0moQUrOCbJ5PrzQWTIWZDx5yDE4viYAD5h1POkBsEQ2NcQysFW5ldkeUYlkgf
K1ACc4wGty4q1Cdafp4kri0R+mf8alaGlCbDwTiDaUufnJDDahOjiDswWL07hnzG
sDSug7PMYabSiDirRoD6vMmjvBkvINDJSkknIuhezluFvfafXwy4WzCB8oE4NlYU
na3tZ+nfScfAwHEUSlrkwp1fP3+Sm1egPsPrHvbS4HodGJ7JWRXUeK0IDtCydMFG
3I5OOxLvxrbF9nvhMEVJjme0iwWia0X9Bj4T9lYts5qirdNdLe4/TECBLID69n6s
jZC4iwJtrXieyr+lg5XIiTccrYxbVvzy0k5VZVFI/Euq0PFoi8jPGAPS7BwseBUj
lu9IjCkru99Rxc2CqK+9K6LOO6Xg+W6YyuA1EpLlj4rex5wtQbbeVadFt1eVwKjb
RNxP5ghhOgFcPIpebuaVtbBens7kKX0GX/4bZyb8hp9IJfn1SXL6eFFfK9Sz0fvO
UXDuXIo9AfZ/kCCqSjAv6kKmOqadCxITgY1cwt5g3zar7upf/FvLmRWUurgswFaK
thmUAdkEY2wt39YMyzSPeglGpLsQyqtKm0rD1fbU7wOg67+4busXhe3cQ3mjiXgr
qukC1xyfvdpwZGAp+IWqGCaeXw73q6Uij9DEL5hd+qWDhGvg9Y6XFgRuxO9JDKqR
F8ioN4Vetw25CVXn09me8u5rcJMbU6X0XweREDkbfAc=
`protect END_PROTECTED
