`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gIZKez8vUcnjHOC3oHS3wgbwEBmkRFxlRhivXfWsPsnypp4reus7osz4n6Fq06BB
lVDeOULQB1GjRmDepTlKFaLEJthAWDGxrfehUgmlYpwJzigjmoJ7zIYdQuPnlXqH
O6+abBOPpTxMTshxsrGOsOmkoNyhq9bbkj1AvTlZE6xkM0dpUrcKkA3KQIdLT/xk
yfrjbB26XZzD/JtW4X3EyY+WdgRNZWSVNc9rC9grq4ogvIxVRjfZbcyHmUzh65xq
MD+i+G7Eh3uUAXXA7ITHw9uxPigLzAWoKChfUzHkOvVwR1PG0BMpIjt6yJPun2W+
KH25zG8UDC7vB9OG1Tp1JTPcWGBOqSSWYAgveCUeZSarCaxsb8IrykO8CINAnbLg
rVG/fcMdVJcA2f+MamTvNS/ttDAYPHy6mwSXdWdALhnL84Kj+fFkIrKs4RFxt5cs
`protect END_PROTECTED
