`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WNhKS40EjBWHyGqsIwWVo4TvvdQipTQUTkKlOsTavrQ5wsh+s1RKZg5TnMdYKgeE
YTYfIgGS5FOlB+TS9Lc6BlUr3yX9+8pbgP7Ppo2K3vf+Auj9QSSekxtdZeIJdzia
G13aYK+Jvt1Ly3fP1EKZwICijn5l++P9u+owZOg6TYkt0BLjK/R2S0/tnNpwY4rs
5LzXNpJODS2Oe3lYjcT/HMK3e3tKdYEIoYGgjHSZUWoDKEa00yGMEfVoY+TAsUOl
NDrkr0ggr326xlkr5PSgeeTSklBU8qWw9c851oDZgltXCXFlbJ7NDMkt+NRGDk4l
Ypntrdv2oFJf4fTwE8H06SJy5NneA2o8yN10hKbcnRb7YXscmZhxwLywuScUFmuV
/+xFMA+2zElhhIGuSOa35acStpPLw47jEwr7aopwwZL/vxXxjXPb277bFoTwT5/X
r4LB3X+gbyAs2JTyXeKv09bNf3Vhuk8+UlJDtMSyooylVvNk0T0yuQPRX3FyDEba
x/+dcIomPfVpRRUIs4CGttrn21J1Nq53ngRtt5A+TfBWtDig2YJTyOXNnBwk6N72
0MmpFUCRf3Ws0F+Ycd5fTHyBHyQ5NVyuZe8P3cTgvxxz8IQ7v4C7T3CAckaChODQ
GgZ9cpJgf9qJXNl8EtME9wq7Ea4JOw3OGaC1/4ibWJ4IHDxK9gKUGVyX+umgD8ID
izPQj+jdTsA7DafwwRi2NB0jY2r37jmC74DKlxAgMHCQbvdsQWXiAyavpkmquRhw
ocN2y3q/3BT4yw08zXJYNQ==
`protect END_PROTECTED
