`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vnqR5wtZS2tUDfP+jGhSFD8dizcC41ZacUDiCMYFEKSFe+ZTfUUW1pSZrqnDlKd8
7pkAILJZHr2hpQv8v9p4EOOGaojmg0FjnE9uVGpxJM3MARSw7Xn4iWd5tmTMPsNk
wFwrwMZR80xS6VjP/U11/wsG3aQcL3Wlp5LkrMlzF7ECFEeNWFcaE+Rbrt73Q+3S
wSbBU/4gEPS7flYl0gVDCvd4Y1G8ngeZ9wS38MeuVwsURqhkVnha2metXGjrpBmv
b0iAgYrylHbI+Vk3jV4ZyJMQrPSDI/MNtC8Frij4qxCrTZN3K8k2BHhUvVIWKyun
KK1phkqhNj6eV6oRZAVCpKaxRSaOwPnQDfCT5BSeTBOAcGH31T9d8k7bpnl6b3/k
PaCLx+RN+p+Cj7ZQQPRL1aVHkNKvykrqM5NZ33qWTjiWrAiiTWq4FwKvGnc7oo7a
LEbQiEzoskxb3DHDPU04mYQpWsKHALhdvIR8qMbPrFQw0ax5nTT8fMhTmIWb1TzW
Fl7qO3KQcN+v4Eai9K6W9lv22HD8vVJK3njWuVsdoJaFniBQ4Z5ivFaos1IaiZtZ
thx1EL1j/VMC/Gv4/5rrZw==
`protect END_PROTECTED
