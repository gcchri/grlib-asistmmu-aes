`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nLTOkbYj9hRNcgysbG5efmciGqiqQkjjSGHaj0XAxL48nGwgvZDAjp9uTU1ZxYBK
nERA7brql8v79FsaHVzpy2LqH/ePaEIjgYG4Fw4w+Ffo6xm1qY8G7YLinFezRp82
AgZV0xGR9q9UAtPvamkxZGFcGIQZLU08b627N8OWe+VwaH43yGEWZZU4WYpzPott
Le9jO+l0v92TzzDeU4eR53uOt/HcRXp1JXbLzyw9h5UU6F5oSekMfhtY+jmWJmeK
/7BfJmV72JXxBP+Y2z2kk5FEkPWQTi//UmV6idE7LYnrBV5UtieOGnJowcvno64/
Vt3bJEv08ETB/Jn2+1p08C2Rl2Lq5azHT5+3J2alQP1jz9p0EDRxPGQVBsAexG6O
ZE/i+maxOgFRqb6iJY9pHLDW8P0D7FYQl0aHOzvap+6ET/uk0Q6ZtFmStz4nOOIu
jOhf8xogqLVua3eqPNCaZdJFr9m2ZWem2VZIZuH4yuO53PO2hMHNxxDKqB4ABTsi
8mT0eFFSBw6VE16Z706t9Qx0i1EM4mNl/NAZ6GqZtQeGKMpscYLJ/S2UaPPqi/HT
gdGTLigsYfleFAeH7wpyKLn4e8Be6bHW84G9ZrBT4Be9T9iMdUSt0jw7dGxEHb+H
+4y+p0u/xlgAbHhlPKTYg5OBC6NXiFS3NNXKIbpZOH+DuKkCpj3MR79nE0OgDJf/
peon/Zc2auN7LLMYYPLj1OJE9jTD+9KhqfEK8BEVgsdLbNWIzZGtKgKaPV+krGjf
uMq3HmcOGYakML3sYwhcUM+lgTS01q+ogviSG/V0JC6IE7EFegtJ+NxHqOGFG2oW
+nwRT62voTXYmtEFvwtmaPw9FMS+J+Wgpeab5QctZqRppeOAWF4unABeQN8GuBqk
kB1pQzKZMZdUybbq7+VVRxAcy3Lt2dZXbF8b0n978xvLu/WXFNkFfC5AYyzBUPIC
T2LxYUheFinsfEH0otYVe//w1NFFAsnWfPcivsM9xuMZdk7wkcZk7t1afhWkupdq
jxgNtrfMMV057+TtlNaGq9pQAtqa1DEbeiedPPATGrAVe2gw0dMERC90RsoLM38K
9PcbyyFe6SdKhKoJniSBX9R5Q2Xs3VwAMarXBfLB3e5CBaXq8tKHgxX13FzD3B2Y
Si5tUilmQ9dQ6+juC2YQD4jyOtq+kqHWXi2VW0Qr02BGvXqGlgfdN8s7ppKVh2Ty
YncqeGR0uCVmMVM6E6xEN1emXNz9WvknUN/VTDrlAsa0YtekB00kXiNRHNThGzjn
N47cZz5ij2FjKwwMX5MAgeieG44KeyLgdST53PJUw0kO+wejEG9yDT3323ufoJb7
CJembC3hWp7K3utW2C3SjJCIMzRemt4JXTUUmbXBsxd056Hso82HyQ+Ik4E6baM8
ZFdglPsykasNRv7MVFCKa95hmCEraPb6djEATHS9LhOmFtj+Q7VHRC5qDllgEBKY
VcDU+2+BNppM6/Us06u0ZwHDoQ0v20t4aCcuREFS6LS04nBcPzSbxXudNIxEc0v3
R8jH7qzrihjx806CPLCDwC7/oFk4idbV5zQatV17FN8xRvShwJpxeINhs55wRt7l
W9306yHsfQYC3XYnRIIpmXEI4MK+lejBPH0IDUbrpIjZt2zIlZzo8QOXV/REsvHg
DNxuQ+4JvvJsm6MVOtL1yXUWNsscUI4lOxxiF/hJxXEtWQicTuN6Ci+URHuvKCgJ
EZLMumMHTYNdLLnz79yybdL8yBB08C2m9wh8Gq+/7iSg27x6NBnwHlmHmenYrtR4
k7EfaAo2sTlhSACfAYCrs64tBr+S9GTXEHfJrBNJQGEzpgsuJdR8q/zPWH6O7bOh
FI1Y3ZQ2As6dHvvk6g7g3E6GrHSg1F880hUaQELIyDPTMStiAdjpep2NjlMuHJ+M
o2muXKfwZ3vuCnYGMazxSgctYknBOvcNEraHfD+poylNHloDgE99NWGJNZFTwd3o
OnfHinOWW8GLAwZjutQoGsAO5E5MopDyiq/moVZwKdyDAw13soDTxsIvC/D/I0DQ
Ecf2u9XFAkNam/xp4NJ04GppuEStluB2xGaMM+DPbbSnyCBtloSslTXP21/sPeE1
lrnoq4YA/DqVyhHhoV8noiWZznvHENT8TGWMhoFFSn+P9YF+TWqCD8JxQUUKj7X2
1Cp2oHSXxpAlzOofE4i3eI2oRfR7ltVbY6+7FU86o+PQc0/g/FBTnFrf0ogWD4LQ
q3GTtvacwwCr2zyhCaGt0oaeWJlTlS8pq35QMeJa0rZFfzwTCoK5mfvGo2AcUWaC
OYR/w70FQh2WBJFWYCrR1ql0lGRtUB9BZoHaVMmOv7UWczMI6bUdHYYRYv/Gu02H
8z9K0Tybn1k/fTSa+SGGrUZi9Nct2PBBJqvb1G0RAvieSfNixGlanD+uPDyGrLUj
/JLsCh4Tn7wFnQT0fzmVhfaagPFOv47XktHrYrPU9Fc=
`protect END_PROTECTED
