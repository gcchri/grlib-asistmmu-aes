`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ji0G+G/EwYIPQbcaq+7wIIZk7Dkv0Y+9VyzGbyUNNnqPVfjgciNUjXN45hTN3F3A
H6Qe8ORPdvvoL/2UXuagLyBhW3AHvy3AHs2+AXOySAUJ67yxGAHz3VzbxSNTvpGX
Wk+2iqLweAX3N2GaTsY7bxKTdxfK3eE9W9mW/w61d254GS/xRsvglPYLreZKLGUw
wesGR9vkPMtSAuqSjk3Rmf5Q/YRe229qzVsqKSAYFcmBr37ZpLMui41vyP1xnwpN
PTA8d7+IHtJ7JRopOHx4RtxLsE+DpOFxuilRb1ecvKGHMe9wGnsAm5Jq2ruUBvGd
/beQBbZV4wupQZTS6i/9vA0JMFmT0pilMoD+IrCEfvi5QT2JAfyfgr45FfRc8WY2
9oFFjwiRa7t6mDdj3MkDGUvDKpRlUF8OjigSpGkuye8zEgC2PEaLQaDfyqZ0Z/m/
`protect END_PROTECTED
