`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6nqXREbezcxg/erp7Foxq1/7O9lXgnz6pfJbcjrob67DJDH7mO/CniDPnLXychvd
Zli0FMdbIAb/rzDAQHiCPMaxx48Q3erwepXq+MCwpPEHQkBHl4JX6nuIDP/t1ssf
gSYYpVzsnIs4TlmWunfTrHEv7rLOy9lfg+tOQ0kEDStOmvyp5o8XumiK5uRxjRHZ
+3H4nb2UFwMAA24SvoX3hlGoCypCb5c0XqNnysbZumoGzVGSB/IjnGnU9ZrBwyYC
LqsyZVZeSFn0aBL/FrPK1GJ/vKzKeM+BoLVcYtntACa0lPRvVifSOAwNUEIgqInW
N3P+qHBWkdXbfMFN9dulYnwqOhfPi2FwV6/6N7dA8JrilvfEHsscrupkdMxM5Bfo
DswvVCQajkPb6lxW3kksyd7Ri2Fldn39RLLpT6DpkryOb6DxTET//eZMEkUFpuqS
`protect END_PROTECTED
