`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SkMINfFioFc4OmpBFbKatciv9CsKmQ1loOOWgKYisRx3A382gjbn8+hgl5JLyQmU
Xc/WfwjjeaRGBH4N64S5MewAYx9YtVEO+YLrvwDpt/UJ+hb4gx5k91FqM3V0WGby
F6T9ITQSHIW/pUnHwZk7nVf1Ha3HbJW4P6knP43+4GHlse/NVLFZ9tAvKV8HmQb3
f0DauaZ4Q6sEhkwXwDBVHIEmLfgWeH8mki02LA44rDFZPVIRv3Vz8HOAZ0AHn3LZ
XAGznysMnOYuVrggLGjzhGIMFFSnpOVhkhWKx19f6FQsIjBOXwjwb+fpyXh7El9H
dWq2KobXNSRczzH14KySpsHr5QqTWGpR8S9OlujkDo6tWiOWejWrTtud95YGT84g
`protect END_PROTECTED
