`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eR2OYbzBiSLe41UmjjhwAaWMvbQvRfuzD6nTT/azG4PFMB4nNT5MmBKSuwg9y2PF
bj1pcMaqVrUuEUdUgCm2zg0ylFd5aEnN8QX7j3Vtz3U0PlskfB6lNLcXEssopAuV
A0pOlsOZi7/FqoJT+euot8zE9kT5vf5FapCUnkv+DSKSdETUgik8gFdCw2biL+ek
3STpOCHK2ySMHBn0QlKoecYYCNKg22mclj8NlW2WH07DXEJhD9avjwEGgpZSMeAf
habIGuupFROjrrRjSwRSiuT7qSEsxY4yrfftfY5ONsds2mNUAzdSJERdx3A8A0Ov
ZUo0c7NhJWc1U7UJgAWarffn81DEnF4hwEllKaz/gJMqMk7HVxfK+SVIsanIBmLo
KmHqLvnIpT13eRNC2Ag09q9xoQv19IsAnuCygo/LoJWuzT98a9X/sKrmylSQ1Hhf
qAqEGtJuSE5aXbNX5NQZAyUMGttsPg1YoqZxKFufHryWodMkmjpDMy+i7cUQiQtq
DR88XN2bTpe64Z0m4PIzQFiFFw526e7SO3Df/FkBJoB4g2xjOb96ZFFTqf++vQC5
Xj4dYbhpkPPkO/R8yAJWA0rlEdNqXk44MT4X8i+fQAwrNgyTx2hmiGwrLl46QTUU
3OmIyg1r4y/Jn2Jwe4w99aAoNNrUPSiqG01h9QiN/9PsRrN1KuoMb0OSyrutsMwt
KZXKnSUUNmLpT9tKrD7MxunEXyKzG+D7VZzwVEkjzcxSqhFYpP5vVEZ/HEN5ubp5
pIKV+TdNrjWHo1UjNepk9BhpDI6q9AXD/IUbVpZMcpEZ4w9E+2Pb5NyzQh7OfbWc
vttUqIXsUkLCdoXh0AegV9iCk106YzADR/WD2qkWGDvO16yYytdhtT1uUdcGnu4M
/vOh1qXyX2z+T1baw/sL/f9V9NuRLZASafn9zILtJdA=
`protect END_PROTECTED
