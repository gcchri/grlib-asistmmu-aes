`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j+lkZiKU84H0hTWRQTjQuJZ0ADtrqyPDs8w+11VbXuU+gCqsJl/XE8fSaedEEmP+
UPqr6dO/IHkldcxL0FSc8tvQ17USdIYoxK8/wsEj1Tnk8WSp1uSccsew5okj6UQ2
lgkLJ/Hq3fUJzT8npLS0Bq3D3gWND80BzMBBDse8n3NGmsynoi4nJC29Ash6/NKZ
KksygAHHUEH9YV9aE5/gjXigsbUBLFEaOMJ0nk2aAUcTcUGAIUPeOL6ETdTCUXdy
82uQrOhUbvSKhliTplI+tM/HKwQ2ZtaEvv/RS+RKHLnMn3ibpP/+spjkjqaQvZcd
RDhlFOm4WTa4o7oFoBlA/vWCYDy3haVS99/5m6HI/eluVpixzvSNILPNiu5akQbJ
L1hGAjQ5+nZLrIbvE4X+VL/TmH7HEZyVGS+/5jSlS2xrm7Wio43i0ja1BMNWWW+s
tpHU92xSd41XHjMT0LaiiRz1pXRTFFg09k5qNsk5kowSn9XKTgRNQAZ1PIhyhSzX
0FBrYMLVVDX71mBZEDK05adr0MDGJydwQTMYnkjihJgjN8C0Hpfgz/u6rMNzPFPT
z9uMvco2WSnbdt9+nj870+wJzrvXbjCppZzK8jQzsSFUBx13ccHdXdn4WUfpM4Ck
IRyE9KjaDgk9pSr69Mex0BlQJKx1HjFPd3iiKq1/NWMCf5qCie+Rejd2YuKsdhNS
14KzAfR7e2fPi3dZJq7GpXNsBtOGL+vWN+pVuPHMGD0wI5rUOaGB+oJb0vd15Kel
LaPQSVHfOsZoP7h46dvyXJBMKWeio2AOZs2luGKlTL9l8iFOkDCs6D8sZHss0N/Z
utol1vyts/E5X1xT3RtinGTDRUHZs7NrjO/aLc97rvwGQEBRmFBGmXgjy+hqKWSk
NjckN8adoC05FRFJOZo1YQ==
`protect END_PROTECTED
