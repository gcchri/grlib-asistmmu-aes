`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zfqAnmcNRen3RmRQC894HjwCxxfpyPhqlSJ/eJBz0NjE31zS2npvgKEQXJr36688
9ykgOWJFiWM88i3aTtdKt6wD6RBqgw0T3jtY7TTQkEwt9AXlvZJKumNlr9tNKUnS
NljAxkVz5Z6OfvHyOBwXVeW5sGpYy+rnaUOTLFDs/igwldTMytLKVALGmpDtj9R7
U967aJ6gRn86xUAoakXRzcT2iVmdmW4RQsJK5FuXKpIlwLdY/CEkSnfrws+UiMyx
m9YggRdAulFZZ2nfMdnvOnK2PEqOGYkxpRHGuSslSXYTxhVeZMQVETjIMF4Nh+mq
jYvD7oWubW8FR+YwpWYI1fP2zgLghOyuDVf3T9ePBGIE6F0NKzVtJcDNdgTwNge4
YUEOElFZ8VmLEVXH1WDgVC7ELrhf6dIJ4EVSYEyoE4R+DkqOKlVTSLAs2E3jz9Oi
JEz30lXb/ci99ynJmsPH6qNNVmNjlPo+4Xj/hGWfrbEE48sCf2n5wY6X6ifeFxW9
CnPtR9snujoL+lBIKw9Qh5wEpWwFQg0jnvZcxr6UVaEAVvslCIem+d+hK8Lyw3qE
KpSEVMioiQ+xb1DgEHmovDEc5xPj29uPdW+9HA03d5sU93YNmSu29Az+AYbWsgNn
Z5i+sXGHpJzBnhKSZ5u6FnT/ki/AJ4jrSI+HUsk5LrRcGQSkA+ovwAa6ev7byUmp
oUukC6A+kS3Kh0a+kWlppfCpei63g13qK4kT+ExRzB3lW2mIgRPJ8K8rDix+g3Tt
tfpMC2/X4EotDfZha7HoOWXmaShsIzdoxHQhZQbn1c/X/ANiDonjPC/CUL5DVXYb
XhscfTErrlPkObrqebrIwuDFmSoENQMnCI/LomStLICrXgei+mBRkOzgUuEW0Xt3
6yozfEZyDfxQ39jSa5joo3wr9rTJdYCCt29UOpiV9ZHpiah2yVr0quDrlNbp07pT
+6AM2lcTCAxQyasqGYc0P0dtoisJFHf2+wOnh4Rs9KGgeGlyXZTR4/IFzBRPUFdz
R6p/oHLxHxGufiRnllJ76zp4CLZ/7E+7Y370KF3rxmaEXOyOlzF/ZwxVLItkFGEA
rZnYRZJMY4mnQqXIPc5BFTj9tZMU1q2AyDULNqkMJlwZsordHfXhrYOT6TnzvZCW
lF2vq+iYS9FrIFpnaEvJlBoaGbIgqNvDy/QnnOOkg1CPy0ozK7UcXlqTIJM/Jwqy
JJwMHjL06Cxl6HXp+tnnVKkJwahR47KUfZvD1YBoiqtwJaQOHOEQt7+UcE3PrvPn
o+hbE+pW9QYfJUM22SSz8i8cxrvH4VFU8PjW+NFbM0OrstFFvt+uI7NnDPdG6h5g
z+MfsngQA6/rKm/sHy7uABPkz8kTX4Pafh3CyerejZKGvjdr5nyQDjN1e1FNCW/h
AG9v7O8g3LSnxxHyRo64qvq/oeaShkC83orQc/43hG5k76Ie0HWRky63WHHzeFA6
aZMDiUrGupmysNkRuG1X/C78pPy1/45puCMd4mR3y3wzAb44GPyiePrGAiIhnb6d
UZzAz7GRF/mcjoGP/UcLjNNq5zyuYygA0U0STxQJAHkqWbvvSZywbQxAEWO2VH0O
jTYrnhmZIbE9YyfxHUvM5Gy4GuwbJHwAAY/mp3YNmkrSraBHgWv4cAboYlrhx9Xr
48upMIYEhvQkKSxIVsXfYQB2xhUy4xxOuX3A1FiqFHglXj050Q4t6wLhDQ6OfFXB
y9wxsz1hW1YST4opHVIKf1uuUSSblb+J88MgARz9wH97GtdZIRodsfhhPX0rBxVW
tHtHSZDSq/yDOs/ua1Og/O2KwVHPVOvM8D1449j6fkmh1eqdx+5pr+RciGnHEPOI
Jc8PfFuQ/bIKW0XZA8QHVzeFuLhFQ+rRQ7GMIIUhPbZUPEs7RxLkK0puzc9U/ag9
TPo7m97Y/C9+IBanVS9ksqJDRzkaXZLYmRyguqKsOPPCaxqHrphgNKRGjKacrBOa
BsAsXg8PVvYGh0C8kZJz8flMDGl3sxkBmstTRBPBRDcmcSboqlh0SMb9dehOS9Rd
oUKn+TaUX2hIOpJK8NKeKQ2+hRpo0ihSIvZfO0jdrsXeYbVarrl2lPFW6b6XIkUm
HT2klBvpp/+5hCCzrI2Ybr5QnllazriHZnPfxn7iST2iB1UBY5hJ/Onw/ZPl7Y1G
1l6ddQX0O8SLgq0ItwTh/GDXFtleNXNuFtFkyZOZOkBTcpc/lcfMPJ1eawg/Sl3+
j4qFJDS+8t3Hhq/AmLg74NVuSfr6uQ42t22p0g5QQfjE4Px45Vw8EZ4fag0X3gun
xiKyyqE9jjfHkPqhNzkFAshpOD/IeCTNNLmnHYNqnBPDA8G7ilyloE07XzDC1Bjl
VXLJ0JRdNAd/jBw3I6InUcwd1dMWPKAMK8FvjPnj/x2q3qwRFMR3Z4jEKrWDIp68
2OiiBWCq36MYeUu6ZXegaDL/RBEJtE/eQaXQaccf+rcGtry4gBB9N4mOr6UlJSYP
nP+oZmZBE4/KDDqiGPx7KtzPMlaERlaYg3/VmWJQZeNq5uKFl02bnBrvcc5hF6+C
i0z2n7npIkSr5odYVYBkw/gGBVCHWbHLhRDkiPhY4x3Lk5cVqL/vTi3rK4PTmr+7
TsnL6MSmKk1S2SJtt6BOJKkcJKuHIUBkgcEE9UTJPFOYdk+NENFAUu0fTaK3r59z
cFy84Bl0nO+ITV+D0DP4lp5uqoqWFlDMuRw4R87XxlhyksDbVhW7JeijokAxgXn8
XAkmU30/bhfjRjl3Jlvr7b7PoelnFVvUtIHez1eFpfZTRmxLYba6ojCPyBToPoe0
SGHWrg4LaM52x3DEWY2OWTT2wx1J1nOauNr8TbC6kBF10phzGWjdCYc97lwk2TQt
TR/is3sOGE3J21dJrBwhRvD4vhGYesDkWyVeHziA9xJjzKdiShVhVNq6o3wA6Mus
rq96D5SjOwHUh7kKCwbOZ9eIyMYPRYuANDty5SPSJWG/H8Lpyaim7mvbGaIPGtJT
xW81EIImzyAQbOJoUdvJmrtPD/2tGXKeB7md3T4if6M2Dz3N8B+/EGkVsrGzgxH2
nwP9ZKOfuhPIO8AMHiTLa2quGutUuDU1WNvr03hRx96CzOK1qQFwH1CjOB6TLwBr
5gdMqgjTJjfJdzCxlY5LRIDSLmQSeKIAdtNgrLZQpaJwUf8XX1OAm8q+rg2CZFAq
cyS/KNwizPBFJ9lYIPbXGqsgnV5uKDD7ZmTRI+BOg+15Jvzowp22S0dKYsPVNNZg
DOtVKMtyEYjnCDYItLJSX6eDv2doKtV3NU4LTv0ltuu4wKctMg7xQlUE8A+YmxV2
05GgKtFRu0wOFomgb4huZPc4dlDBbC0yyXWq03BUs3QdRh4do3FUmPwa4sJ4Ssgf
68qAlRzRA7aPhB8LvZDX3DAEAqoRDBq8ZEbZ/Qs2pDYeltz12OJalVzl82EbR8PN
4Zdp4chdoPSNN1/Fx/ynW0UkHPjgYu0OGwVUOm9kJ3irakGrBufdjXnlsO4adcoJ
Bf37kXM7+UZPZdVEhPtS2mpAxmxI/jUFj4MN1WvW+/a7wXtOPkl47NmTMuLA+rjQ
5plaZzk7mILE75py0Nh8JGJJX+0LgKJBw9lOUomIfrsGaaED30ghURr8IEMNC+B6
ZstToO8aZuzYHVB1msDDGirz1lh8Wm+tIlrbIWi4Y2Bi938ydcYq0UmvcRO3dzoG
xsDvozQa4vzkmmfkiDrdnh8bqymixdFyPbCvtlzaVisCG9xCDjek2h962qfnP+Hu
RmHmA04+cCMbJ6LmeFlxBKjcPmKqmje3XZhRZeJi3wbTXkphmK9ICL/tvSyIqnyD
cVQSMF2L64GkjGe/6qG2vCcn1Scen9Jn42j8WpLRjQBgCkCrXqVvvf2LwM+SCTyf
GteG4R3mcWdPeVQUgFY5iqMw+CuXG6fA2ZwIhZL+ebQNKxajuxdQ6hJjcOG8ffOG
HwSAW1fWoN0+7yO4IJ+lCBSFDiT0PxYXnalBn0pSyR0p+GG19jlQde7cJIVOTyIF
d6p8rpM0B9EIxhWMQEqw0UNcPUfkwHWb8ZM3sesaMoFQR+R6dbiQYkGncuCAflwe
p/9yyu6CvYHU3KFn2bBLAn++PE57B3jK6U06X13sCmRtJFlPUc7FVzfTP43E8PVo
7lNO2HcPcvYqQG3iRDoDvxB3pK3+D02dhFSeRt0hgK1htN0uzF9NyemeqLPhWU+5
J0glOizKzOatKSbH2iZ4akTLYQ6uy6DzzQbEmiBPdnOrULSVdjt3/n5+qepIZTd0
ADBHL84RHDEpZaDMUpc2abRHt578WhbFFXYdIJb3yo7+ccVTQ19ebHBI7ajnuwLh
EX9M9OtJ+BJ+ntRA22DkEYAQ6JX7DHxb1kcokgKDSsksIcjQ+KKqAfRuljIOzKRm
TqAngv0P+TQIzx6aFZw/VNoKFi/XruLIcof1HWzcSCRjtT/kpsFrc4bWKlcMtSRG
RdbaBrfaXRrwYxVOy/B7Aa0wYMMKCTj4N/l1AZEs1l3myqmHA6XghB9+6g9PONMW
KVjYCtD75KnExFO/XCrAP4b4/6nGcgtaWMRme7KColrJUhtPFxgaDgyrpt1Zv1Wa
1ZidKyQtSnUiV7QVD4HBOZdiF0K7r/+m2myQKTR9trAtRrmwIQLyB0IxWxm5Nv/p
30Q0otKziwAp0CHkEQuphMYC3R18c6ep2xHb0OPZwFS2BaKwvu1NVqCt7JX+16RS
sxZ00ZBgQsjkPv9mpwihaGsCL7LNdYoBPccNxIxu+kRP4K3WZegzHxKq3VhzBUAf
K2eMmjCba3lE4FMmJRd2bw7igWAi/jMFgnMtcl8sq9nIXjegfTzEZN/OlwfW5pvT
zRJaIV938jqovcCCc3RXRHphSMHcQNCQUb5qWLleVW8/NVszf+DjPfrMnMXhURni
iPaQsOxhpOkjfeiOyFFjNL1ODMMMWWLSN3NhEa3ys0LRk4OygHf7Ng1PYpRV9gOn
ZmJYICoNdo7fM6nfxKy5I9P3dqC2xJ8ATh/UxWK+KO8Cq1qACz4Tys4xuTHGPKCu
c/WF9HaoDJrCHT7W6SQjDgvKK1jgtgvdDiK/cGDkwrbo78M11Epk4qyHhoLvuA+P
EMeirJlpUmm8Y0SMrOQMwRlAO5bPHGxN00gwN4AzByKUjV1jo191/zW9xLyMKFNT
fR3pEO3o9w+Jjl/SSRgam72zqSO2zgaqiG4Affcnj3d5Oj8xoaR9Ql2GdOIBr0Jw
5AKYbTE3GKqyJM8RRuqLx5Nen423K3Jah9zOnqNuQBgcummwoXWF2MIUyaiOHztR
KA8hLZQ4QLAfL/LYzOm6Zz4xJPNlLULSgyRwvWFRZ6xFjg0xzanh9zd9mT9eLy5E
VZB2P2DMTysIr1eOp3YVXtT2R12AJDRPXIlNpfAA/D9KDFR0vOFs+vVHPSQdWsn2
59yLDPFChHJLWVTp8EaJ57nppel8gT449uk2ljuvVttI92sVxMQzZ0rLJz3CSXFx
xDAzOSaDy7DOao2B0/9lWHSQxgVTXUmR1PbAjVO40+zbo3EaSZfev6mTafwxkROF
OX9+hlatE09i2p4HXRIOaJF/u77JzhR73p1KCDe+urW6ElDRUp/vuhSZmN6pEmTV
Od7rmmbWU0tv8nOMyHW0LtzzEnq0ZWsLlsmL5JeEenCwfIqWy6g5j0QjBkpHv098
jpcZNNoya991l9BzJY8C0CFEMGdEaJROTG4cIsd+Gt7apNHIie6hQLgXQ0JXa6U5
qXlzss8EZbI8youdeMoF2X1xJ/UOGL6/JRbWnoZB3hIWnKdumBm8nfN5HQqHlNI/
WFlsNG+f8eJONFcY05WaNypL1DhJ/kZEyN5hJuhRLAbmh3gEhDQJ2BTTCd80131/
QXE1JpOSWrIB4ZdU1Di1KxCKoEQCqT9fZxUq+4SEts3Kc2415hFGAg+ub1jK960u
+e4vK+DIZVuA/Io7sHw8k6D9kbqEzGRE+WmOwhxFgpKzf6i2VYKNz7BogM8Mxrkr
JB9XD9PrDBFdYqwJ3XBl+L0wEnDXmzgDtvxFFVFA3Bs+Vk+0p/6RAKCJwOevQNf3
7kYDl8+wW/nGdcP5LHbp3uoywoWwGbthoqoTBLxWTdTqVpqFnv5MePEbi9kpzIeM
o6S0uPkUcznhfZoX1T4t9Buq1v8CDpRQoA1zTkW3dNC4pzlO1dOMYH71vsNsaho8
OqB4V4CaO0GhWM3JXjP8FD98OjDA9jXlLyU5DuxYGWiHo6N9Ay7ATeqz3cowtWaB
EcK65uyPA+dw8beUgOHVfOipwYZG+9QWXVB+PLRlaacOg/SZWNohzt0ZUJMIdt9y
wWS+b+UJGObjUXsfuMUr21v2lXxVgkm0VoQLzi7pXN5munm2huHIIoGyTIU1s5gI
Z65f4qmSxaeFEtp8A0aC5hsbRhcNOQR3av81y9J0NYxsYcLlr4yfEMRXJBIXTQmv
K4zY2oEQPexCDJ5HcjROD9ZKz5LC8JNdLFaIxexShFmRgS5dkdqmYJgKYy27Yr+K
zNG79xpyUyxmd4VF4P8bEco9fWLWSUQ0InRChc7yU/pysU0HBm/dtNJ9edQD6ipL
UYEG2xFPo0eMkhp/W92s7a3dZuQsbd5wBqVjEij3gVWPWMjSTQ5O/T3W05m8JXE9
cMjkDFHnHttrwyWlslMJrCo4raWFoPgw3LA2ckuKJc36LLiKIAaojlg8ek/qTv4B
pn1pwerdg550jN1igkmFy88+Ey9FxPEKM93ix4zjKDKDfwXZwyxwVysaiaIqkSL1
5ZlL/oPz+1pzzDAE/e09dB7heyGrJ/5Sa2SFKytfz4xBgfca8howgmPT6UtWBZ4t
W4B5HWK85hKPGreDSBrxc57Giox5CAwW90b82eGGm6EPMTOggpKn0IfIXmJeOfCY
b+LGc+n+iaclLgvHPWrgMwoVK6hiARdjDfsvzv/1HR9W3emkXUPR9Y4vwoP/73PM
xHjlQsxGp0snH+E8boOzO6/LwKyBavGG17k1L9eRdfJG+vZfkHzMqN3LHtxrDJzC
OxSDltSNY1jVYEX0e9XhANWWYxm8sf18/sNLXXE9a8N056e6F1ANmFyzVxpqoq7e
4D54ArYZ6UhLJyEU02agiQM10Xy3WRzkEIjnFZu9z1muvZQdJWtU8+GpU0Hlf2HF
jtb6V2mVaUAVQAls8gcpiQK723QOyFt3HlMOYI25lAHb/8l2pi4psObAfMDIV5NH
IsJ2pv8FFp1kMC1eLiPrqRayR4fOpL4jNg306q8dAC71dNS4nFVA7Y13jAM1R62U
FejENE4agA4g8ghX98ZA7mtCh342ZqaKcGjbbLmWAGzOMBGHb+fbxyXWzrdMRhoR
qdHhQ4nVZ3Gu3GU2NTuVkuH8e4w56Y4TWdA2P8+15+vgos3SUV9SfowSIVc66Drw
uMmIEofwLaOnXPn2bGJjqybH4iHpFb7KubKkkQs3rSdGCldX8SNMfrYrs6TEVtiL
ubvpWchYnjhr9jVJbrPtEji0xOgaPrf+3A6o2BWysPGNO2R2fctp9WWNiCv9+dke
Dg/5rsAjG5R29ItpA6BHHMqLm+GgVYqT5MMkJEO1XuF5GinH41RIgZxbrAs7LFWj
KQM5iNzM8jIyCzxmva/Sd3Wz7QcirvuNp2ags3mJ2yMrZF00RB0HhpuwLh5ChNrW
gjfPZ3l2lYWq63nNuAlgwZ2Q338FzMiE2Ue7W1B0fSe8Oy4gWH6Pazi/LCrXMI2d
2PD64OMzsEiQBhcNEs3tzzWP0QeRWjdH4SrL8k/PqwfK8im3JPz0trxeGOQ9S77L
zF5dalXFds1v3PfhjNvmG5eUVSRCg0BNpvEdc9h0SR508gcJOdxqFRJZ8dQCRqd2
uWHClgttc78mGqyTGW/rNyVnWmsdDVrwHp+K01f3RhvRQYudiiJtfyEg9m7xTmvF
nUdq2gDZV9MLo9lUjl5FW3SrzR2pD0AwWWUlDpK6NahNbxFvhcCtG+WtmOZow/XH
urp0Z7Gy9F5/4wWhOpSk6hj1HRT2drm2QGBancZ/KIp3lJriSPZG6cINnjzMcVOK
4lJ/nLz0Gbvo3Am+BFBxiCNy+8BmBHHSdlEluuQcKNkfseFQ6nKPuXx7T/31m37W
KsBcXAo1qlO1ynier7BPdT0xNzvEyMibQ569sTlWJa/ulIKu8Yj5cfApjzmNjTMg
rxAU8HxI4G8QKlhEGDxUn5+fGExOExDXWPjdDiNlB9qy6ZINEITrM2QW9wSn9ioF
Ya0euI6pUSTLv8Z+q4yPQpqdyP0iyfzJR6yXsF4tJEJDnK6GBBEbRi7rlsrp+IUc
AsgDUwmvi8uuJq2+bj4vhmqnCmT2u0d/cfB9iOaYtxWRTKkmI2DeBBfwF70liGfv
RWL4M/vc1/6fj2Pp9o9cwU0E3HMA0fcpyxxLxcmR7as4GoOtf2gpoQfB6gdQtXIz
TTtlfY8tDEF8AK3f2o4WO8cdImIuwoiYcfvJPGfMi+4jJ1KablLdI2MwoNrtfbc0
8x2aEpkwgdjQg2Ir1reMx1JkLI2jAE6n22vG67tr61uFRHY0xP3KDirvOKnm62HE
jkAP8AO2Z9De9Gzd07CRhjAX+OKWXS6ljsdMJmObrTlnpFUj8Eby5KNohC5y56C/
3kS5AoWTC2wP/TzAZDM0fTimzvMZYsLc3WuxDIvyVLUKSS0P+4Z+qtqcNJktioOK
26BWMF7Tl0P4ck55bHl7scw4q4Ns5XGSKEFWh2PKQNm2+Th0KvvcldtGkNz5jl/p
a9c6D3vfC30GarplRBbRhnQC6Z1DLWc29upZ4Bz2iXjIgBdN9WKTtyNBWhUsNztb
tFrY3dvYdKdzxVwpV6qIF3NKFnmacjPcbu/FcXZQtRBZlXskj7uiwQykrrPFcCyQ
cSAwCz1kpCGUAOMccACgUBmcBfcckwTCv0FY5AuSHOrxgeCmGL7LzJByen7+3QiI
q93XEs108gIStBdbFQ1KN8OWvbh1EN67mRKF27UFDMcyupTEIBvn05ezyu0A7KdH
2OItktd66nehprlpBlpvlNw6sO2RH8GVIoXUl/jJ48PzdjzepAcKfkKK+8t/+EDy
DGqKE3pJ2cA+aGkfcVYOBcKOEPFxqbo0cv9Nn1RBSP4zVWgiHDZRd7AAF+rPJ+h5
WB9br921/d2iNFUYUBBEh/JEmhtN7yEu27PCfb7nBTHR5B2TlZqTbNZCY0co0lcL
01WVIFZlR0NB7qrD8mqogDW7AeWmbK/dNRybBCXaWAyJdUFiPOND5te7He6FLpQV
IqURSZ8vmL9XbILFI3moJ+MjHYliRRPu9KeFbY426Axv18i/5Xl2iw/qDQwqdf2i
BKszvv39KiEFwf5G2+nKUhY0BH4QnY2OxuPZyVKxBLD3ob3EqovlvMlzb4Qo5XdM
d9xIIDx7wyhj7hE2pT2cSKYu6K7PhYYLo39/WDAfIzSizRJBHbS/NoVD1XCk0l5H
cUvR7nyu6XUG0sDpvgeA/JihqzDOrB7qZqmuskkGHgX0pmlz8PPx2daLjVmkLU0N
pShF6t17vEl1RQC1ahlwW9CNJzmKbc12jBL/XbZrzlwW18GY3sqyZUUaTf6SyL33
0tL4J0RKgHNX3Wo558LnBSqcXseMdFHrgQw9nwOpG98rgxTuClK+pXEYsvEIW66j
QXYGR5+0LMU1jHjdDEB4co+Icz6TojAQYIhLSMJw6lTVOSLVdFKFi6p8UTOsgAVi
6QNQbBMWr9p3PdJ3Ihb37g6YZYcOZq4aicMTGGfd9x6n/jQC4+zXXHKGh9Vy59Li
w66aufWDdAw676vfvIUPfMNnZyEUWC5Bk2OaeVhb5RraB1RsRnofoNNXcl0+nffe
3yyI6Ad/ueD1BOlQuwy6O6kwFxCjch7cm/VUPJfxsdG94pPLNstX2Ax+Kmf6qMzz
GJSGloUTgYwGSOPFAEYe0NT0TMWNox3mvd+oOrPY2pKHtODG3GpLoL+EE2NP0JM4
yU7RQrIGRFYlGFraSz/zkcDKy/iKA4w9hHNDjP6hHy6sSvTHaViCu+A55pUIdwL2
2N70+C3V+8s5azLMxq4EaDeac3ztQGWd8eXYsIyCxXY8cgk83FdcKgaXyv+f1y0X
ubGnY16dX7TN94X1k8jsLJz6t1PRRptD912Zfvx09erDZcsTB9CKhXanrGEwdTnq
NIvecS5VreJlKxUePgciPln46fyrGjEuSashD+5iyY1tMey8o0SGXJxXWlO8BTcx
lyGGMrY5KFrSIh4LqY/VHrBsWX3IMe/cOE6AoqU+rLHnBcydipmQCie0+1kV0EJ1
MPCcuMjzcMZoqsmk7OzcUsKNCKw+FaPw0Qn3bjPYyjh4TdiHkJu1frS+Iy2jxhqj
rLs1FWgXflyrzOLNlgoqqOkIYof3ec1Xtqd53NLO7IZxykJfo1M8z6g6ICM3194r
3SKw99HOn91bJJ8wWR4LHy9HKkfz/76oTparP6em5hW8El8HYgGGmW+EjnNxJ5LN
V3l4gSY53SNjqq4S83UHwpW/u6KClKA9j/Ye4ZrLlPLOQzeFtryJcIdeHdOVdozm
8hXPrLZHB4bZHjQIp7F1o3wO9451Yv2KUvkNs5NYkj2A1omkHUVKvQZ+6nmC0ae+
q9qBz5hDVImM+nkRZ8JNlo9usvCycL3T3ljw7xC/RR5lkgkNhz+MWBpt7xFdjYcv
i4uHRLt+X7CMFWiqnPYBS1A1bcE0uO1xqqSEYsFmG7zDWILpqxp3dS02Gxmf4g3+
/RIocgXWTDarz7o2nuvS3vAyrXJBtw35JGUc1JQTbiOU9xkTh6hHu9T3LBasmeUC
ToNKjwGu2eg2LXXcYJTed6rDUVOsoU89CtVZSl/awut0lNG7NXqanoHebAVIufDO
W10P24GWqZbsMXTQQHwMLbKg/lxuYtUXilPfRxKn8c+Y9ctlAkZdoShZTf5gGOae
As7qGwjGOkXvE/e5MLD4xmRD/+ZJ8UJv0LWA6wsd8MXgjwhBkiYarF2o3Bm/rNKC
6aBcG63GxWfEH0CESXSK60ctisPDlZEPjSuwo2mqdV/ThutZXblyWiPv+MQjOWLF
fe70E1iZLQeQ/fBnY8+wypolYGkOV+yp3Fs7/IIbY5UCNvX8L1ZpSvo9E6D9HMa1
VBZAXbwIz9fKxSlmd6a501iPXehdCUQmr+WF7zX3D612jmVesoFuMMhfMd7DfvPv
QFBPq9qDjtIqefW214j9DTrSudOH0D+JMLS0i3B0At1IfECeeeYUoYK9Hl2N1I4T
WUYx+oeymHnNk3TAjzJN38KDr4grxTZDsQx0d8/OYD1vcZuxw6xYQz0wiR9+opkZ
TcW3HPvJkJAUPgHDeAknj5SZYbfCVB0J6zufZ4RL44qkcXfGpzJskW0drARf3VSk
zpZ41xjPfNiVqcW9bB6Nejg+DRH0U0tPWkMd4rBJDYCl+NJtng64w/rMNvu/CYro
+C9h3GNZBRxrQrpV2h2Q9XOTRuivpfEYwSFrjQNwNVvdhTyQLnAqNqjLIntnBGG9
tpxmLVaPV5MFU7HKXdya5GDRgl12tjX9fhm/aS9dzRoXFuvFzEAUx5q1mAieT8Vm
twGisXrsJk6/jHVoagxeb4xbXbHmdT4VkVbRVBnqP4q3ct9C08+YVAAWWcabYis/
nJdc8vNBRP/OmcRsAwbR/l7L4TLSXpPephjubEml7TYj9LIAftETAdF4iEDQlVYo
9W/LBJo6ap0qwAsh6AYpXoIQ62Q2fFsKbHfQJJzyaPxzAs9iY2hoQWLyuSx++3BE
QwF4XiXE1JGTPwHolPIV5fHnAqEohIVjhMj5v1lSLGwiPeBkdeYoPil84VnV8bJi
41lYRRrSZ6Nk/wNS+6J8MqCN6ZC3gviad9GHRxb/ALYscoBDG/s2ozU28HD0d9Cm
SJ4dZLnxJR9knIHW+WFKzMQdMCVttKQN8uwAttMcXaGuPVroqadttm97xWMdgFs7
FH0iCPqwG4AVM037ypjFDxt3BZBCWZIFDRP7rW6QeihvQ2Ms1omcIUlAsY2WdoDU
M3DrZmZegr22CCmMWUy+1XFnmDA4v/irwnihSdzpUWV9Ox3oR670F7mhbSporTCG
y5OEnjWspspDsoKDk91DY9VI+7Y1oXOmI1xbiIxK6qtKW34kzNyzjAD86EGKtCr2
kFqTKspjPoSze/5JfX7XtdA1A53ApotKH2Q3BNnfKxe1i7akTiK9Gcxkub7fkug0
V7ZOUUkw0pul6kqo5FdivHI9MEDjZy5fdImP81fjy9F3fdYcSGfee9HCxZJageIX
Li2MIVZFbu7kXRXzTeotQWwjFFZbEWIu5wrdfbj6/T9V1RkNrs8/SppiZ0m54GTS
J+XFhvEEzQ7mloFtgZB8MJerj8Hm5aOZW85XF63+qxIYVmPUQ018L8iAcWi6VnJ7
4Yfe/q/47ZoEjt9JezQePVMfJbc/eQ8khe4Yn/P/AFAqPBw9yeV3hNuBLIa/VuZJ
V/IFkQ1gNAKUsHt95v4QhzVd6yNmjOAJDI/0Q9tAtaPvMts2zvl1/iPY9LC7BM8X
YMRB+Q2E5c1nFSARfq8ACiOVs4jwbmDozvpUnU2QPuVaEmMxru53u8jGpYotrSSM
i1QuslgvjIowoPEdB2zsKA9s6EtZa1NkLa7+MHFQW9Zn/Zl+plopaIIS9rb67mZO
Mq3Bq3Ep/YfbcmGNb2p1LX/Z/DHKxVjuoJSuX19Hr01izxpM7jLO8JiV4jFVzr50
/PEbhtTmbWi3Ey4guweTwQ==
`protect END_PROTECTED
