`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xSKEJsD6leyqDsFcB5Qd8BZIJzaYL5R8r/DWiWaWIKEZ+WPkDf4U9FHSnbNmx0GC
RfD4AJ7TxcTklSTtbmUSIqkWsQSTVfdr0HbOxTq6R+3GxXkwnbjD9JTfrpFGJW8N
3s+cDBVCs27vu+2q+XE6zFWnYIVIcS35HdtjaemNPcnO3yGwtaXlDUYkeqPz5Hkj
Nl6fWkRR4eMIW+Twdu6zvYAVMwRPMgQCxAaRA/bQwo6rdCrurfY/EMPdtko5J0OF
dG+QiMcpG7aV3Hh+x4a5QHY/uQOvcmf0wborKSPAYvwBj/n/CbnpyGM8g3FaxLM8
iJFFMW+trKom9dygSearasxIaVCteRYLuXSNVMwnXeL6b7u9X+SNNx/Fvz2zJSjj
15ABigRuzVSmFqnjODKf8lE2tbaW/0eHB4ZqDyWXP4YOu8OGJRPhmizC0YXLEKsm
`protect END_PROTECTED
