`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C3RjK2SnSr4gjwvLgew+etbRQYEwlRIwyGlL3mbaoaNP5tCu/xIE7H2Gu47irc+G
caigHyQVjfiPTZ3oIHaAZJm5hGfnKMTtRQy4gEAa2k4M/BA4daItkoN4Pi7snlCp
2Qq/nw4stNrrHPJD4wY/dXJNlqrRBgp9NKiXWu2jxJCM0RvS46OoMkg6z7FVo3BB
x7fIFbjJ77QobDEm1ywZQXRcQ+j/q6B0+yjC3Pl0riEgU4QSyG4FaOk5+UBTMboM
sOuutRcS6QFiUzd0pbWR8M1Lp28iNx/YhiZVqk6hLi3GolwYSFpbRCQfr+h7ND7k
oN0HA9IDz1qXHmQUZ7zDf0hrE6DRL5sWWbSmHWdmFNr1q+Qx1c0oLdG/7jNbpEgP
Zw7hYJV9Q/icR+K61wr+cLhHDnUy/2OndS3uBcegrZg7ukgFK5PoE1bJPfw28H1t
Jo5ztWtl5SrabkS74Tp7haDtX65t03NLf3HpNSEGhPDozK/vWJp2W5b8OsqQCT6k
PUZEYXBaWekdfNrUILzc+kS0BQa2CNkX40p9bsKqZhUNT9WLeFFuCNCawetFdRso
z7xg971ow9Qz4h4/pXDnEBzZHh38DRG2nm/+C+ZYIUBubaiFMo/hjuIuyWg3MDi/
n48hE1GHYDkQEUC+zFQ4PMqiiCM31CmlVTgQofq/NVsBaHR17Y5mpXUqF4K7rNp3
4WBHgahyqbkrpais16omQFSplwObDDtTeiYdA5wNGTxFeGAY6vesmywUVd7se7gS
Mycj1Xh61zybSB9ibpuSnRCp3In9D/VLiMMHKsaXfdvM1zyYdP3xyAhdbSIgG8wP
efblNyKCqeF+wxux7iTMbBtbqc/vEf1DZqYyxG3Ewyr3BrCwAT9VKnJYJXLWgomd
3cCuHi82FV7kmUcqes2LNHCMAzYCjo9zx+uy8LULglptUcJHw5mI/+w62ODxwo0e
AtGDinXm8Kn5Ycq31cDI3OicQwxGT++LnL5Q3kbDh7cfjkrtprXQi0jZTgKgow1X
Nrgn1sAqhOOd6X4FAlVcn4NhaYIYECP5D8+8ZIUX1GWfV5/lK+mZvRHFjuKsGVaj
aQdAaLBOg1ZK88lz9X0CX0BrEbGYyP5vhiI8aFn+ZDrTPDZFWK6/AbtXi/fmnagq
N+qBrR3KjcgeKb6ihQEVTNewE/+9eHpAWFQjfZl4Y8cIKCvhIU4UKPWCb6AG6a7B
gCJX7h5KbiloVmajAMWVUm60LihZjA/Q6YJ848dAjHc=
`protect END_PROTECTED
