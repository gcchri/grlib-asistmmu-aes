`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
18qCF7IbORTVs/R6hpqw4swLld+/mfHs5rLzFFp1Jq5rWw1/JZlMXNV6Sc+VqZzo
eig9jzy9q7voHkWyuL6eRsWCqnWHRWkKRbKg0awjwV1vW1o4vUlrqBrkf7OZq41W
qKQfKYBi+kqmwh+NJxs/7rpj/5ulEwdVgJmIJ0Q8r21dhyGI/fsTjshZ7mLdv/KT
Cxk1yBlr0H9Olqk0qQnfeT983z1rflM7YRws5rqlJuGhbpHaeLFJkE6AHz1FnXhk
T0QWzcZtfXtVvp85Tu/3ejdof9l3go/VbDrbe2OObUDaESHdQSrylVnVfiJAoIvd
yVcvtexhp0lZO0pHy9SQL/gEqBMUISGQcdRobZJaZfj5bUpry+mF3vUKu9HBiKow
rE5ncXLZwcm7A8PMSkizBsoBVG3gzT/7u9pooqSHzB6MOopEpB395A5YFDfpKm49
`protect END_PROTECTED
