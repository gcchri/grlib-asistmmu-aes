`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dffFcGGpDS9zB2A5RwTvKLXdSvr7PRIWp8j+/RRxrmBG6QikoqRklyQUSzVipqIa
NDZikJQVoyTtosHjMmoVy17MdChbL+lIIYRtvsjoJSsNxWJ6TBQjJJmUKGsOz7yX
/IuOY+96oV/Jx2moJ+32uPlRUZUmeUhmRqJcq8JcZDHeRJDdmyvtskdZL6sgDxnx
aC1Nzl7RMFgestoirIymFPCwyJqYemkJpG5bkR/pBbrLl8Qw4xI+qlNN98D6Afz4
FhUVg7KcJle61NF24ORBGlBpmSgY8n6dw1wJv/SWRhp9dGzt/fiR7M4Q6DXgRnIj
3cAgqtEsZ/astFMBqoA1C+Xqf8BM1Tv26kbNipAPgUNet4xAU74yPdIhtFOHyLBG
jLv1XLNJvKF58sls28mwtiYpEsCPvqhMjFl/7HCWc5UVByOiyhyYWIlaIPq1L0vO
P4Kk0RVen9cQM6SDeKTLsbSZNJb4dL+Qb/koBy4TYigJRVz66omY4og/pkrsnj5E
`protect END_PROTECTED
