`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+YeVcDspx+5+vmjxBg+IS1C7X5d/00H9o3KCYqKFkBlkWuEuH4XStdFSFEiWbnK/
OMCiHAvYBEq7Iv2pAXZ7jj+TH7ljPqpD7lbl66bvMBoKrBzE/99djOLUad3trc1x
YZUOaTzZ6Tn1QRbE2Gu5ybHSc5/zfQICkaPDdFIy57ocN8fjDmJImuUYSHomz22R
6kciJ7nJN0wjSd/59yo0uL4we0eGmIhFIrSNmh7KqaWGZxyQvaq0BVSp4Ol2z9wQ
nVBtpJHJSF/bPREFty7XfsI+omDm94seS5l2VeSOr7gm/4fZ6ZtZkiUewo6l0hYa
zRYeXjLN7z/GEsZ3m8Iq3cKv25MqAiwIrfeIJodSLhhvGzFV5AU2AAk4tqVTWQKM
JbrZ4XYhYY3ycrBDqei3GC+R7VnM4vkOn6sxSQscGdEqn9xv7qeNXXjCuolVRbvq
JN3mix2oSijF+wYS0hLojPI07GUCFhbHc8KV+XfcqcaS6D/M+rchvO62JJO94VO1
bi8nlkgQ+FOXfW+eGZo9UxokK9xN3eMPqURZUcEJRWUsQjrgiKed/6wTfKTN/Wb2
GzddF6xuwOORIXajTloT1gmhp6oe1HaUZTYoR7R4XFd0EtpLxYJT1glEiDOTZQ+k
aDHbGvbtLESGKEN3j1Vq0PjKcxW9MPPrxiHeJWoFonQpMuWHxNNBmbOn3JMZc5Js
RqdzyESobYI+7W2lWjqu14pyiTC7bQ+TghSaZCI63yHorRGidGcftZGqj/3NvAGe
eOtLSM9Mh/uZfJ553w2+PoxnQ84eOUs0C3uNr4yYs0Q=
`protect END_PROTECTED
