`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eupIyFJZJXkqeoYkRCF7SuYQGbgofSnytKzpqtucanR9eUZiOHVrFsHjPIzj+pc2
THfz7Fl7PKe578uFjbk16w+XaFqvXWHRtu0NSozW99e1rbIrV7s5ZrnlwMtywBTm
DiASo6RsZRejLRF7oFaDiEMDF6BCGgI/1uXzWkhiZezT6v6ueA5PcYXIDMO8egtI
wCC6waEr1WOQ2+t3+q5d43hzK5BmPbxQKWiRcswudlKcpGH+21SvDMRZ+enx5lgC
Czql71FIFtKGdaO8Sa3a/nUwSoEeFXL7NRf4PEUTnoRjZRKZEYHF7AEUMbh3OrC9
L0p8JI4hMH2LARGmwUENWDh9WHoBy+3sFOYCEVLvBOYmursHl9z4cWuGBl3c/qy9
dYly48FFdxQSlR3uquEvvW7UwtimSo6wpU4Va6q3BX3oLfCY/x5K5Oqd0Qwm16dY
+rmTjJ6pM6VOfrDi17WyCkDiZO0yNN6RTyUKDri4P8S8WgeJWCzrUdq/0ZXvS9lh
LuU1WxFYe3fvjqMCBvpx4QRmJLlr7zyJNJJpJI5Xj5yonDQnQC8nXcYVz6FQPmy3
HjOV03nrf5drAt4nWwa/cFjfzUuOIaFy7jP4Ybm7SVp8gvvaUwVyos4GqDSvCfX+
f3SKkX9bo739DH9Strh2S8g31+xtkY9wI4jDHYBmb4lAEoBvsRLJ9UvQSUunpt2J
Nyv9xF9nywg1cjm0oxvbeK2MEciNBTNBmJ50oJsWDadx86LcRA2pQhoGNjredk5q
7HuGzA5yEFUnskBeiM55527kkrx7XVfkr+Axgzj0L1RX1RgwJkaLSfTKqsYMtIj/
6Ua5thsxvYpUr3rc3FxSCGLfeeUxdrmOQKz5OfX8hqF6LhdHa79dw++NpENaWp7m
ZjfEYEldsBHTw+DMThbh5iGbTc/WiLmBW5/uz+TVas9CHzvA2sFQCH6kQdemBVZb
1cfDaK2d/Wbm+f5MTti+w5hbulg/3glC0WqTYmCc5l+BA2W0TxgcRyudsX2TcCvW
kRqBXH+ZsAg4+W9i+igqLf9jZM6UzB06sYl5A6lDt09qebB5GTu3za4ZlR5Ph/S+
`protect END_PROTECTED
