`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YFcXQrfFXLtfF7MUiT13fabOMnKc6ZJCQYjKafCCm/7WcRxDl4mYHHX4XwIivD1D
/X0jWbTINhfVjC17SI2u3OB0jTHAM9m/TFU6M18GJQIDAlGSSU33i6p7PdDw1u5L
D5uKeFOZSPYAmswixOlNEglS7eyqTyYvdcvuJwuaxXYXCH4GAfGQAJYDsFlu1upI
QLgrYT4G3NyTWAo8OVCc2yMvRyuCUWP+HfU6PSsJJTQ/g38X3hMqWqJN+slEM6Js
tcg9PSjbj0RkI1NPXMhyaiRDLxEGa6tCnVLWGjOOqkMfnXe0sUhPShj8Af2V0KrK
cVxB82ylkgGbDcO27Vw/KSwACK9evZVCI11Rh736G8ovt+KQwpBdkaGqiD/IP9ft
/hzf2YmWIvchEd/Xuv8GWV4LMjsuRiCnrjfrKkI6bihEmLf8DFa2kvpzBWKeNtK/
`protect END_PROTECTED
