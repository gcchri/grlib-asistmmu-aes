`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LghNoZYoIpmRWFVzO3numcTfKZDjdcNmXHOEcqmQ/IQVYkOZACSBaFRCXcHePzgL
M8nZ5OVmEUDOq2F45UADsoptuZo5DKvd7qrjmZp9W6n6uj8PfCE+ilQIDtHIZ6/b
YR1UDmvO/bnVQ8GfY+81B10WQM0aaTe7+bbWwVdG/sv8EEfLG/4QUj1ipNv44tEP
6j77726xuQ07m39j8Vf8hMO8JG1xMnQWTNwm1/oWMAEVCLfAM48DhAg9Ful/PK7o
joDTSkRQ5IB9bFWK99/58TyGkUHbc5CTDqo2qreNaCialZboZjamvwaALtfgRu0J
ksQ/UJL/fDxVXuxg392w5jkU6jMkP72oHHwfxdS2WUAxtA1CsHaO8naHmdA/75Q5
9UuNTGymg8wLbiMf0WokokLovDbzL+/mS4iYMnORC4RIVa16GVp0iJnE3cLvqCRx
45SDJ2rTewLPiWnHwFCmH/BBJJLMq6Lvp+bDIv/EHtYeCyJwaKGjgwfJkbB/ufFq
u7LsXnnpjEQiZg4ehl+QH8QqR5dpJ7uRDZZfMFU2R6KtrwQdVSwJst+n4tP4a6i2
959s6NeTNFGA2SuXosegtaNEwQ8GKBhuvlDq/L9L1nuZBMo/J4LrUQnTT8+HGnZ4
hO+PuXT010unBTh4kvG9GjznRdJ9Mi0hQImmlt55W/XnT5mjsLJDn0y0hupwGw2Q
nUivEr3rtxooHcKU6LmAmiNJiiPz+viHEePsGFsE50cCFuKavSychxOX0KzsoIcd
74Z1i+2gm95BjrT5xUiilGwr101NQOXpgHBcjaRVNqo=
`protect END_PROTECTED
