`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sOF5D+qU/DnZWYzrPax/6e9NC7bsUtnnN3gqxyfaDDmFxkdwO/oJ/8JOPomE748A
JmJbFnxNTHVCqX70djsCaPDXGf8RbVw8qWXEaHW4/7yVvJxMkTCq162IqUx3A5eF
XY5vnPPXz5VeRHUAU6wCuxAOCyMo5pXlUzKf1pNq8yCCq/nPjoyd1DRK8DyxaRGS
trtwRvhgR2smvOPF0U9kFwkwStC1bHpjbzmMpG6Kr12NCQ5fKageo/pl97Xz4RHG
uZS65Tsqn5vfIurUzDKQbxg4xmlZyGFtWQWeH7RAweIEFcgeu6t+c5pwxOy8f6Ex
TYzrAg/q0B5uhfxfg6oXcXo8GAWbpbBKzEWo0q1x5IJr7ZlNVTM+nvL5jclj7VE1
skl6TNfXBFypQwouGByna4DcyWGQ2rtbhz0C+tpNbDRkZDbPIC80ku9oGlV39cEM
celQKZROeOUwV5pdhgrAtPeSEYu5hrscd6r9Bm+cQJCoZDEUXBRzs5YhB58iSK+I
vzQ65bcYHeFqAUhJP/JLNQ==
`protect END_PROTECTED
