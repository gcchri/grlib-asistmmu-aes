`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SboHiGL+gEhgEPYJn/Ba1ti6iYBDOKl6zaM90eb8yClIiBItvx7HTB41hag8/zzD
Uwg8Y+2QinR01u8QOItTQfNtru41xtDx2MI0J+hiYTdvF2QKqm7rDQ/rZUEvcn6M
1KXyNZLNBwJfFhH1tG5qwykViqVvVdxy+0LNNLKWuSjxhp/VrsPBce02qhjD5bC0
IfrsBK9JDp3wrs2hG0aRA5unHU1/Ns0QWIUJdbsbsEc2HhwG5DGYIEcR+dUvC5ce
YhNyqmSX/Ar/faEWVUMZgx1jpHw1kOXrMtRJqmaqRb8=
`protect END_PROTECTED
