`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CzWup+HaAs1JMrQFFBBqZXpMFWTtdHDTn95OPTIelQ0TYJMYdo9W2oqL/45Qa2jR
1faTDpqnRkTtIoSYEAyDzSS4rNwsgq6+UCx+2IZzqj3XIpKOVBQztpilO1/srZ7a
/iZWzjIcl4myyXAIwEey+Ejwe5yNApQn/F7sYeGdfnzntnxy3w0MYmDf/V4k66lq
nCF9fWioWsdQ84G6Jsrn+7gpv6MrN3fYBCYYW4+TF9KC0QT5IgYPVL9A5SXiYy44
KOJraPO8y9ZbNGrXIr7qyTACJko4P4zlDbwDCsZOp17zyCU8Q2JosoTCMSVVFTwZ
ACzFqIEAdrexAk5E7aCeITOkvB+oLPxeLrBt9hcLYeyrSFnuIqJJpKGM4uqXdjgg
8fvHJZ8py0gbE5lh/FFKPIW2NzZUsOG2qSCmGU4vJ/pbiZ7et3odAF1DIdbrbUEq
8iM1yyTB3BSb6eDTO9QS/oYoIR1WpG/IfeoXnZnQWrpBujgjmzXpi3C5wqb6Phs2
P4mRq6cANSmwG/Pa7x1cqLpnme0j2DWFxcz9fAi6gbP+0hhX7S8116yL2dgy5G6s
oa57Gx+tQFPqPZdX7477j2OhOzKe0t/Sh26dWEJGkC9OoNhEPsRXtw6Kz+kBNUjW
nvufKE9d8bOzhpuHuSocXAUDJmx9EQAR69s3qLrAuG4=
`protect END_PROTECTED
