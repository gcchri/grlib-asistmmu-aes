`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wdYs6GlqeMY/D3bcK0QRwLhDf3CTALg+4SX2t+srMycIEhryY1BgrhN9fQjJ1Pzx
2lt4zlFuoOAn6hB5V0/On0gsQJDq8yK5qVXJLB12oJfZrOvTj8mtp7yLjhJusN+m
OHF3SvYDrZQOvpmKUdCU7qlRc/ZCbWhAwsmcpcHTggft0NgzCdXAYuceccpVCpYr
r6IbVU4utiy6HaBtD+S3NuLq+ifBTXbonpvQXUMUnNImXyoagJdXQ+16liRcO/8/
Kr2mbvHhJ4pjz/mLxftkxWLsnEKmGgflpAfKUNfiBAXl/Z1Y74qZBUQV2+4SQGY9
nSVdnCQRx+157eGsj1WEjUPtZkf7iv/WYDtlOF1/svkPPyiOp+a6R0iEtSt7ZHC2
t+1n0Pwsso4gB/z75azRAEFbxBcCgxC39Tl0tSiyju3jfE11c2MYq0tzNdXcrjb1
79KWuFR9GJJqLUFYgC01wCF+nUms1ubTK0JOqPeeZDBO/SBJVdypr+LD+F9l3aap
W87WZHV1/dkVcnriowatvcZdL3oJzq3HA+7WlH4rhx4b+ano6ZN8+rrTeDZ4hTyx
9rOgMIC4BZIuYwv8Hi9vMcutpB8TgrfpxKrhwygQ/cYSfg/0pCGUCR/HGlfKYKK/
0tMAvfSXjUOnO144sMB4sSKdxD36e9yi3W97RvbjmqUefLcVU5cYZ+asehgk2FNq
mShLr57nFZ/rs6m0pwHsLSuOSH96V313fSpo1rbBHaVfg1dJWaugKBEi+Wbo2ubv
O1FjSWAlzWRxMVcCMbo2UsPShDyVLBXeZpl591xyRqIvV+oAKiIvhgZiPZ0oz3/H
s2T4z6NfLml9m7sfT7PdDXQ0iGh+FD63Lj/HNyb+TbPuosidV/3eCMmOwFDdeKbz
xGWFBNhLDlaW+OsximBHOvmZXxkaJudcGxOhIf2bxwnpNyaUEfOlgzhrGchT9Nu7
e3WlRpY4ZP14lbutUrkoI6y6EuRlZZOy809lZgPDnTrTgTbEgK4J6Mq10zUxMZNR
CIAvQm4QIMZir9NuzNQyDdVnI855MtyuIYV+XUK8tRQeIFG/auCgZ+5socxHwAgY
zwccW2uC9hgLsP1bPLQtlk5st7QEFTIpQxYSx2wUZMz+hYf/YjkewBD5yWGaRWXZ
mnhVwAAljWjXrSBfl6M64KMKXF6tAgAC8x887UD2T7DICOmQNWKXjxcnQpDoHGQS
tpXTRcYBkX2FKW/wprb6hIirKlfKjqb4RfKa4ic97CTO1prD7HL+NzGIRyPZKc4t
EzJAZdzzm7UTc3CFrt0ZgqueT+F85E+VFe1ZKYMJwDUqNsK9S/vOntnhWE5UbQCd
wwL6wvv5ZE61cjx2cZxE8e/tbnd4dJ+wZHz7IhSfHTiJmxefLudG0/VuJy9gq9PW
1sn5bUVy/SYT7SNI4ovB7eLvrk97VZpwlSJYRudnfMxumGCBICmCzPnXgL6j3vDl
XPOgFDV+qlY3p+BEAXrSv5y7rcQu/kEI6FQzS66nKbdWzeOf5uvAL3STYQ+Gbq+/
fLhGRkYo+Tr04LHb/f/Z9VmnB2hlubi4t9IvgDVE60Mko+9YHAVPkCt5sq6aUuh4
ZKIUVBbAO+3gDsbKVpPT7Mf7pt0VmsoaBPbpBGzNj7mrRWyvacGnUehfgIzrKxU7
KjystHEOjD+Zxa0HSVhQtGTJkZi9sWHkDNSBYv8Ev1At5b+yBFff1tLBnDaIaTPD
dZszRQlkqo4bgVdI1jV0NxQ6keno5yiG0NZT1UUq7IpM1TeDWuPrwVRGaItuSg2h
WyLu+5VJnTgF9/SmEGSxU+fme2mgW+snSVllsKXkLcxjoY11DkSnwsnykJ4lRLCt
UTDkwUb/NGqApFkCsnbHMCepRNFpOfNTiQdlTfG3VpZS5MOZUuyZb4wOxyEMCY2v
Ei+ULW4ur2wVku7zALBzct5t5yCYDW70lAa2F0XRmlxkUIVJWrliIpTvwCljJrum
W/iGLvjpPt9dxQ+qTNAXhJGz+w/xUToA4eDSlFCBcui/pLFjh5w7kWsrigCGoFOK
QLbgfsbu3dOF5GXc6spOnDJsDQQ7uwHid+d+xbmgYfTc5qpVm9xeDy2U4rbrZuBW
lfn00IyVXPL93EKBkHkEjwvp5iJjGUd7iLBinxB8FgDg6mo5VCy91iICgsRMWqxl
ryLeSIdZXn50H6+Xx6lq3RTw0eU6dX06jPfJPhgWhpu/1lySbWTDCMXGwLZ4P+uX
l0OLq86nmUH/K5XRcYux9QZLcCi6ZX2ZbNWjyzaRfY8AGfzt2f1uO0DQ3DBWw/Q3
gbgHZ1pDwgcL662EWdKwly3NncCEl8Lyu1vFp/SSThngdZ7PsvFlv3TLnRkbpjaD
dnt/VWwfao+U/6Ryk8GVmz9BO4oUbrv52YKT44aK9orwHSVjilvOGhGFDsBwIuF3
5wgKW/jS8qCt8YdsnA5qVHG1Ofu1nZ2jpaUEQ5qTmtUwEn5neTaanl8nMfFHzDTm
xkAetl6sOem5HOV5UiInnMp3N4dnfnG+7NOICAe6kpasFaEY635fuHMVIPjV94Uk
D70ppVXBI+Ms5QGSuXbb5pqmyY0UfSp7TtEwpdSpaCnzqUOBVbUNntNgS7/8VgXg
eralgSzpM92+52ZroTFS8onO1ljUPnDV7RkKagrbFkGDViTW7Ll/EzAkpqpDdGWi
qrwWDfwQ2TnS2DmDEJzoC3stUNI02vp14HRSIK2KvbagSC4lan253Z9uARRTFU34
mfeC4kduZxTa0XuPgKA6CRgfVlN6A7j+QdxYiif66bUTF2BMUcnxSKxSb28o3nXH
EylyQoG/gFSIvp8ePRvsde/gddfF0uf0q4GqnOCivnYZS6GBla4nytRRAE2H1m+O
/qaHJNCJvBVvXBuH473v3oawEvgbORkaQhHFRo01IjvozR06eOglEI3RiORbQuAy
AUPOR337v0v5LVKHil6IQjncXjiPdou6Gb78oX71kVO5bd9+EINYaio0sgZw6Sy6
wt98rTHW1UKAzxNMX5hpQqjmLGR9lkWPke+fAE68wJFCMXkg2PFVWyLSrgL3mL20
D9gbLrubXRGHeopaAhXNqbx6me1fSEup2nbXpLX1pogXPihRBPkQwXzAlekw40jH
WKuQx9m/rudaY7S4tulNpqeDDe0dIjj+32SgIxcq8DOc+/tRW5JeV26hTo/utYPT
NaJvsLLuIhSbuUtpaySQOT4+ZgXm7s1CgIks25d8CVQerp9u87HRztRvKppisrjg
HnEu4Ea8nwUVIz5x0zXs3jVScA7Tiz2SzgA8bw5DRPWA3VOOJBOx8CKFsDs9bcOI
JXq21Mw2Q3mk+FRiE9RWCU0RE95Q3oY3bJdGINyfGlCllug/3l7PonlXxCqHctiq
ozUM4DyodckDXAKG1ZjulHxUUGImOjEqDtgkqoVoaFX4yxOTnJW330KOwMbnG8Yj
hVaMljlm3JgTSiOXiemAOxi/pUS2jFuRh4+u3mVfCJXSq59s65FTE6Bm3RVeOcYl
K6OFosm9K3AHLH2JKxM6/6ShI1ZvEdKq88hH2E1PXKoyluRplqHiDO71eepWXa4q
`protect END_PROTECTED
