`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qfr4as5bsiJGet4j1ekA6E11EoqjuR61+vVkvUyRjLJwIQrGMDdJtgRFBmiZEPSL
kl/exh5B4q05jJ3Bx8ZM9mBtivFgkmnrOdbxPq90Ta5a6nHjxsYrlMSbeg6rQKpL
8cLVMQKnmyGVIl1/eOEkh1Wl+VCuMPrMPXEqxqMILFFmTmyoS05guHp3SRMzPw+X
EMFVnF6XDeNq3SSnR2UoxhRqEY3Y7gwkYy/pVjm+CnGvWvSiugDlO2zxuzdfSKhA
QMbIJQwxo0shcdBqtuG02ZB6vQhVOtUH5q6XrETcTSD29J218ZE4FgJnRHfMQ+i4
fOSyc8VWXDmsRIGMp9hUKQ==
`protect END_PROTECTED
