`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eqsD5XEji++XUg/WQQ+RjThFDJ0JJqAygkkGt0T7m6BtQ249t9xbqjeHC5NRN2PO
v9TaGGwqIS8KpP1OF1n8HPJf0PuCARIiRQ2m972IrhW6sJRan7CeHcDe46FK5EWN
jgG0Lr9r3bLJb20ypzMsqkULCRNwFruj7nbxDJ0YFE9qAGkL8+MeJMQvUDqFTyWU
HzgsLHuSNngySNirpPYMLGW2qqNqV0uGFGNtgpZP3+mvAgQHe/RoO/jpkGRey0mu
JBKu9eYRBdhxXnjfFyGSSE0Dn0TSiV3a6u7v2g7l2/uhE/EoFNvXjGqyYbG3S9UJ
ulKXmHTCIV7PintsCoPlR+/Dm6LEhIltD+NEsriGqM37AL1As+BpdXmPXdxykiy+
t5czlKoU0pJeIrDUVQE9dYA/fC8lkT5LGIk3nFD6fa9fbbZk4MPaFVFSQYtv1wDj
rTy7/2Dq4HJpLa7CxDqLg/mnzvRQNGSESVyR63b64HADYIkZ3LpHyazOBcYjVQRW
`protect END_PROTECTED
