`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ucNVvF0W7zAb8ql619wFHyAdm/7qpTdZr6FTutzWvbpfh7JgMxAgNe+ijiAYXcYx
LmdZQQ7ISOb2edwQbzdKQTsYf32MU61g4P6huwd/BVNFoiTApNACTCdYRWURFx8x
vezvDHUaGiYQHpAEiP5/IzYzlxjt9mgRBGY5d3YfDvv5gNre8G4ro1h71C96d2WZ
5DbfLZPRFaZEIpJ9mDtshPH80/eLuysScUMdhBZFoSh7OB4ED/sNoeLR/rt/XbCK
KZRsFDbpQXvRIw+DF6QkWB0gNSVx1QrgOFmbNFmQinsT2yIHutPNghQcYHQE6GXi
yk1nLl8hCtmtCFLPCZ9CoGJDCPhT74cxYvnudPTnI9/eHsirPWDy50uFRvmmWXbe
q6QnS5MfWQGTCQC5erZdifU0qBxanYvBM1Wwpkl+dro+TaJFqGzDkon6BItHEe4e
oIuS6aeVqRapMmmpnFqtB85Lm1jzsdD9TTrzQgIER1sCVvCjAtzQJvITXdhugaEJ
vNTlanB4uZMQajfizt32mm3dLe610p0JFZBLWc89aVhEgLhyZQLF+i0tUjpuIrEY
m1nNKIddOFQvf5sgTAl3RUCiDEtud4H09bgp65JXj9cI3LlyEjaHBdqFvY4g5urd
iKOO4Gvy7z5Ed1WBHs+eRLwTYOWMIBROJSe/uIxe0ztK/GYrDkaG8/a0X7X3xcBc
lVkUE38l+ifaDqEdOmUnIKLC+jQ9R+ywQcjSjHsP4WP5j2IKU4c6x/KxYWxSblLk
KPXZOG+sztV6NLYL/T/XHjZh1tZn8Couu/5QUQKqNcZjZ3tbzr5aQFIAAr6iCWv8
mTpYEoHRNu4T6LNvz6ea4qyVHHmYsfjUwlN3AkRTS91nWPah61M2EsDsw6UnNpZq
6mtZ2/lvUqntvXaMWv//3pQOLjWw7sDEmMJ4mjyOH41BL9GOkYmzXLGIX9LuZ9Bb
fOhYCOUkKUlTSd9TN1EWEJgijjDXEjC0w1yux7t4FsfnaaOy21MkaYqPWT+dtkdO
JyotUOqr9VMnEma/8qS06u44e7T5XUW+vX0DskXUYnDJ68fVmhchiVMby2os+lXg
GzpE8uo6hK0cZu6q5WstEtuqT5/RXj7h0DjlVVTwWr7JpJd+fUj3b3Z9d+MC4p6N
oE///FalDNjWDjng/4rctNLjyizfwmbpXfHkJzSZ5r+bJSBfjodre/4Jbr14UOnw
3Rerv/gDUm3UD66e4UwSG+PmkUu0/h8ZlieXxokPwGkGWyXC3xYwQ3cdd12l9w6T
eyghOZ7z7vmaho8EyGtrbkI/mFZCg41OWZJgvMKVAc7He0vKEIJ8m2YY+2fIe9UU
oXLoDKM5jNpSYFBuJM2U5qcuyH0xo/KULhUsN7916EpaxUE2TSE3xHw4WnAUcXLG
MOSWrdCB/yHbNOQjTucWfJ2PVu11aJzLS9Zy7f/A7QiOHXG0EapyAzacoC9qlt4L
ip8T1d649xmknAF+bcCkYRz1VOjvWakVPxFOTF85mf7/Uwuy2oCc1ZcOY0qvwsWj
UXsmBM0s+nfaIwnRemC3Ei2HbPTeP2p1oJU5IgmTI7U9fnM/hc7pTFF6TV1fpDjY
M/370ca7hsVYCeyusdYUkZrb4piJlk72AQzVr96cT432IPqpJ8ABV/P9INaPniGc
/4CasNF0sCCb0qT1Hzpt7/iSeutkeO5ZKgnDW5CheyO3UG9a5a1Nkyr9RbvzBPj6
iUZZpPtbS243KUS/jgzYCNi7azmM+OuoHMwg5MDOu3RdHlUMk+qun2VmwE3Y+dH4
nBGAFD8BfpI8FEx6Drx6rO/8KK/yoRFhGSRd8d3ELVvvFHNSbaKIcym1TgZRkEoo
`protect END_PROTECTED
