`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ds1tmc1EWozvqhZIHFqkRZdUedPW1ezr9pq13cofCzuI6j4PzxhcPJfQIUiGx1lT
25oUtUxBFB8nT0KPp0ddx0IkXf+87uR383pWQAJoaTBgRAyvx2U2YoAn2+Y6E4ur
Q0b60mCrMEfgymsH8Mr7jRDjBKVj3uRzgz/+0ZK0HGfUQyLFvC3OQkVBv9rS89cI
i6gadXVk+o+KuAbvFh5aKjHZzw9Xl+V56ROLm+bqLZngct68KfjYsZ3smOqxxDws
dOSKc23J82fxGw8dvayHWR0tU4Knl9pRtDc9ZvgW+O5ANNEfIlahFPWugTwjFD4B
v7OP2gWftl2lA3M4ImP0S//YXKWM08R90xy8IEfR7USZ8hzaNux0eHNQ925CtmS2
aC75/J02lzs+q8APdSsPMg==
`protect END_PROTECTED
