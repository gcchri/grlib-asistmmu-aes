`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1T7d4Qs2T7R/wCiiF3wMkslggLI1MI/BD9lxFiO3sr2a0HOKFFX/RTYnb2DrkKSw
KftU4pDpNY25BBT9Rk4UX+0ySS04fvu873eM7b+MQ8mHcIVikmNuHkHZ9O//zsdH
j2i350KwbJDXJ0K25PWRh+r/z7ngTMv1ds5kEpYeDVyYWszW3QCBIBHl3jgjfsL/
zsypxUl9ouUxy0RY430NBWwKYxMw1SPgSVJ13bLUcpgWYP4kcNEiYYEPn0zIYRbQ
XiNIYwibCenESG9JBrXl7zAl/FK9mRrqeJVpEirYRjRVrY9JP7fIz3bJnvMQ+YEe
ohUEGqyIYM8yPcJIyBUAdf/ezEauzoFg0gmGxau6oUoMfJwLIciBnKsi7GStitSC
51ylMwTuRzifebgMh787NUnHhlzUB/AIUhaBXsj+qg4nNamhxHewk5FXmD4YHlvx
zy356HTn+mRmAp56z/+ga4XQwZxDOl1sj2obFxThvq6Cc/U/hYcDdMJMeNIQ4rd3
WYiJYQrorB301KB2A3sXFzmRjHOdeDfCluobT6RGAuk2EEdqYBIVYZrc5YcKJlJb
4n4nmu1NYKKERzEI/Tza3RArLij0dkyn3EG12lSCRNF8gAqOdh4VWOfkwyfypTZv
ytB/wj1uZdlgOubU1kiFp8DWMNmbmO6Gks2QXQ8J11pY4Yu6+PRFo7eq/Wmn9V2N
99zEy5GwmtNLNVNqeA8BuE7IAji/+UYCbxmnWApmU1UJAzSpX6EGiu5ZFC4RFfpd
crjBRDzrMPRNyiayMp153lV31q4D4BYYhm/fYBwfTfARF/oEVxu4dYx9Khvctkv4
4q7UzJRBRr3gCR/1ktWFo+wReW1qye+QHtDYUOKo7VceIZQATvpp6KJsxWHXBW+B
d4uQcKdRFJkk0m0cF8Tg5ejSxcwpFdC/hH+FFq0ZgtpryLM0yw7obq+97lzYab0T
h2Yj9GyyNtERKk3CW+Ys7N4jmHk+QUcZhOtmLFk8ft0fVCdorB7mCrFzYVTlB+yS
`protect END_PROTECTED
