`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j1BqrdMg5uuqjdC+c9Eey+GzrEbtUTRFZueEBNeaJUIcJ7W9cwNV5xF5CqlHTsFN
hEnWlBuqcChgIYViUSZ0gcXmrFuB5UaJswzrxc7cYERf/4Qy3mBx2pj0l7LZxjaw
Zz8VfXHYEj31EUSTAYE25zA+9cV1xW1aJ53EultaSaDiqX4hnOTelG0jf0dO5eN/
V+xpUCcBZPnUXu2lIIREzJf/yRL4eny8Mi3ZEv6Co3cnsWfhzQZNGahc7p0BX6th
FBQVWw1nrphwByf/52R6qw3SaLERVWuLxsDi+bVqTT3Rnr+mgp5Z+XinZbn5JAIg
FPehdaqEA/Dzv36zHPY8NCV5LOznM+9JkKGuvfWQnaHeh12H+CTfFn56BSG0ezEr
sKtJC9yglcCLsC5fh72VVA==
`protect END_PROTECTED
