`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3hrWTZCfavgQpCFFMpFEno2k61utOEQNgnfBzxO8U0Q8gWVBXGrzQSBhSzLrJ9EN
fqLfP+c0mA1wTQuX/WIp1KHgNhpLRQjOUNLFhb+AUAcoTTuJnAFx4ll6sxpQhzYF
/SmCcJVVyvreaM9Y4LoXTWbI9DWeGmnEhBN6WpbTXL07qOgDVHjeLXdw5Z0BiATJ
vxzzAPf7iO8ZWQchBSvT/y29j0lRZBK8X8rLN12kPj2QEt70PN+4ejY0olGRjH5F
khcow8j3fOjS7R1Pc9EAYqvrPeWY+n8XRSwRt/Xcy3+HDiPxxZnrQWwKWGC9VSk2
fqBz3LoI2KslzXq4yWDHmtIIVjbeGu0y7GzOgmehc/eLvS9UMQCdlGOrkDPuz3+x
acHwgwa5dvNu86NN2rFpqcaoM9WuTqSy82ayMA9NbY0zIldN6gp0T0Oo3MSX5WD3
IE9guSlCXBFGg05pvn990wPbLHwp1X2kZeulYv/3UxHkoi4qo8W5lmZQCq+wmTMA
zhcKGUWKiY8vQHxen05RB21taAA8pMmERtC5u/A1n3xu4QfzRdlIGk4hQwC+QxrK
ZrJQ+7h2zhQz3JZcpzZ0LpvfA8fOIwuk+ETPTuKGK2ijAvxsbFZ8F6EVDIr6LWM7
6ukzEr0oBTf91tma6E1fs6kvv6XCdqZrMYULIipH7sbMj4wbrqim761uROE6srD5
QHTqqoGk7MzXkb8kXbzMimebf7QxUs9Y7U8l6iNxqUll7g5tv4VJwKDPGaH42bRQ
aX7KOleah0/WibDaitc+6F8vOUffD9L8uA7NmODZOlf51sOKZit8/KWM2RiK453d
XpB4YftQlUgr7YF2CSnh86i85PX2ugR12hE0KXIZz26DVz+M2F9YZek4gsSHYp5r
hfaU+ElBYJoMM0TDRY03HHW6XJkgn+kDKxeNoHkK6jB1f6JcJJCKTPkHt2JNNQd8
XK4ROvghqr81ZwxN6hvbHxswlo/KiMd7yqCS41RpNJLa0BJUW6hSmWyibaL8rVti
FTTwxvIbR+4qxGMNCVp6aRiR972TMrTxaN1cdui0mbXRz1XSkeZ45VhEwR1Ogi0d
SPPTR2EVef9Nckm4ib3qfjf3utMhRQrOk/p4v8Scz7E=
`protect END_PROTECTED
