`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tBBYzr+iRulUbxQtYju7sTYg7j/gOe4LrvobyGfngcQOm79dyUHEvAcCQmawzaTd
bqsO0J9pygDlY5NL5I9dNXiAkWkjUsThQFRWQAj7VrTN24LuznNRkoliSMy4LHF0
hPWg5TSBnWsVVPwVBjdLJ78m4NHZCb8mTpMe+B/MJvPL+mAohfDSOcukoBXwFl8V
Pgm2FDsRMTqOkoxsSNckawxdAnJRzWCq4k3Ed4Ql5g4ruzz3UJCGC0mvM5d/34Sc
mDSCqE9OtLG0+0nPDmEgu0gbJTCs4Byb0v0hXSgYlF3s8sJwfMzMkG3QEfEBeSUY
zoqO4g1M3cTKM3xYDiHElflM4e5wEK2DUA8HHOtgQqQ2VFy1/KHIDjCzF7w2yy54
`protect END_PROTECTED
