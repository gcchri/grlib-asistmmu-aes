`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TsmjU/+TodvYcPZcpVSoqWe8bFi66Wi3Qh2K38uhB3bhxbCkixuk35ep4zzTeXES
ExR2a8ea67ZFAAvSURMg47cNyzLfzenp9TzN/OOj7plKO1+EO/HGVn1rThiJrJSr
l9yJMmvg5V9gb552LUMySa5W5jNqZRs0Y0zG3Kx/FwcBTvhZ3JHQH8K0Hk6q0QEE
7GHuvYhvO+mjttis2R3oYikjN6776T2zjaCkZLh0/3GJZ4nbtYcV6uw97KQOlnRw
8rt9pA16QnQppe6P6lPT+XPohE2y1cAA6pbvPMxJZZv8RKoUZy/8kjousfRLme9s
BzXcF+85H7AMIn6F5avpDyyaezutjsra6YdvQ8dGOe02j1B/+2bGjdfVhSeAjEhh
`protect END_PROTECTED
