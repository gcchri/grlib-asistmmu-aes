`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NMpdANsYscSYPXU+asWmwlU9hUDiswIxQ6mYxnb4JYQdiGWYfterHmxhgVZxHgfK
VjKt+tN02IjC7aMOG28loreMan3FVU0jUKvX5kAp3D6yBlpNRa6P2uzxfUrMsA+w
U3Tr6x5RNNmva8zD60THpRHU3KCObnMASy8A9aabUNWrDr2i0IfoZ67tpJhjjYjD
MmoPxB14THgXPU65KtSL2gGpIi9P3niGBvxNItF4UWrXf/q8Qt6AkZ4yX6iOkmuA
TLIOKHoGfyv8PMBUU6K8EQZnWt36Rqe5JytGjFfOZra3EzcEe3KIXsUIbud9Vh+A
W4gJ9oQwOBCFkjzqdZW/rf+wLEKoKYeSRJJARWBqwnSzUbatnSe+qJ9SpqRlogyA
d+Hjl1xcy+JMeXvPDU2AqXUh2rFferVy6rDuf7Y4Pjchs6KpfX9/462ftrP+b42+
885N3YSRCkIky4WTv93skWceHYDYjcPAEiEEYfSGvBQXPOM9tNKcY0eeGB+rhjuR
3ukSHQr5EGBw8mIGboNq18znJwFfj0fnDMmZ+IBpNXcok70cSZTBsxD3d4ojMGeU
dcNid+0zWltLzajb9I1bGJUa84ernBaWIPpawXUeqF9aCY6itx+mhOppxB4uFjE4
N/+vADg+D2sw62m+kUs3N9GxvdmMIRrYazf7OZ0L/HKMhYfbt3nCjTqQRi3xOUrK
rL8r9lTTf6rFK9TShloBEhCwJ7PMpi6Ox/jfK8bCfujn4NM62Z+CLy4OiLh2ZZGu
FQsuTAY9dqCjH36CYDhq4eREHA+TaDPJgJl8h/6uokkboPicGo483XX3RWCBgAca
GZU8wKNiAMfPB4GXf/deN8QR1wOMltLF0v5h1rVW/yndte9nYJ2KNP3Ba3zXhakY
CQkxK2ZwyBOmwYwwUJOOG/dQCNdjafOljKo28raXAqPTi7v5Fap8F9HCTEbdeZZd
SY6zp5AU5aeipJwASmx3WHQ1YWepvPQN6rAw8YvKvIuWFpx+0qcu+dPqZlP+4Zcz
`protect END_PROTECTED
