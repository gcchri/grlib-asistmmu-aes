`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oEy6Dsox0He8q3fMQQ7W4s7P8tZCaTcl2sjvNY/t0DKRUqcPEW/QudroWK1lWXRX
Kd0m6Z2DhusHIzrwj0as3iwafbh7mhdeiyG9fheaZ2QdpBx8Y7djSvXPD/gI1AQe
0S4DaDH1/7DNOVNnE08GhKAd+VHHNeqwpYV0buGpDCgkjKyog7ps6J0UjI2OST+0
VS9dcKqGBoNERcMPmG/MTOa+pIRCLuaHRAJYNUvb4KE+vq/lQZxT3QDBJnYzzR//
I/q2DjVlekJkD6+WUzPT9PJY+WmRZkh66pLk4kWl0IkW8tHH8dZR8ouqW+uBCf3I
zowtHsMH1gGJDWDdCq5Ik8VKFX9qrjyLWqf5S0VyYVf4ebm3k9oiZ+QWr+UR5KF1
OMzZaKHrdhU907FHTLyNEZGWwQPh/oV7MqpFkRFc/fC+hn+gdFJJDzUU1+CvuaOL
N1kr0euD7VsfK4nWG2QF8MlWLkFXg7isKhAS0P3Zwnwpc0Hc6ulQSY/Ie9BaNQc7
FBXCjrkTVHQAIAno32YDuKKHPkW5Ml+PTZoyjfeYZ7wS2GGM2M4GQBfrPZMKAOnV
yk8vflV3ubn1MzE1Qo2yN5oU/H1G1m3dc0Ac309rzFIq1Q1brBUnkC3hXpnGFFKk
c/+QOGK5yCx6wjFA9lPv+h8aPYlkQEZRFqR+ZdHqzd6IfE2/T5LvkGP/hpR9i9BA
ORptbwjQw3ikALJ5h4BjQmzmQA7gHztAhLLks7YZ3E3S8Fj4iP4sIMOiOsSOIvnP
HWCSFDcWo64RYh1/29Sj3MHrp/95a1jnm6dYXtypM7yUr1HBxcjH3jMS5kDhUg8C
da4JrlMaQCr8u66h8HoXXO42NagSHZ7kegvikNC/snWEkcVDXgO9ymw8CdNjgeF6
RVC5fHYKs29jX9vwyeeKd/7QIxiMoUYZIzFEcLLeEg/VvBzhHM0bv03T8SkYNGwV
mNg99HBjHH7y4OezE/DU/suEdv+N4ksSGMUGV2ZwEtgV5wsDCC9VHHJsnIVwV4+6
x2Of5NfBqGNT2bgvIeUpVV1RNS93DskrObGEeat+2ZeHv//378T1ZYB4RLTwUcdA
5hqXeEXs7rUskClJpQF3+asscD7azhdpbIJ0oTQrw7zUyShxskY/sU4qYqOk5h3f
t5P/dFfdEeslphTfil4C2iUjCXVIJyywHwT35xg7H3VTKIpDia8IFuRkoDEsFsEn
1E0kM0ti9UANqCe5OZH/Tj5eUJTLYaXLuIysEjZtgc7KFGQzbASqylQeKBuRIt1a
KyiIWJeN9+4+RboLuKVK5Ep9KTXryy6Rx7Ddpn0xJq6w/LFuTOxTlAUmtsRbNJdu
MqfOwE7nXKfoln7HDBJqr3AqC0Cv7ohtoBqka/VEBS1Jrj/wY5sTedJGsXXbpBXQ
8adwloQmJFb+RNAjJxzuKu72l6sYhrqtiLmHjT9xe71uVDYbwX0P5j7xx4DiSPdo
Wash2iNsak3oaAppZGZJyQjbi1JFJgHydwxSoh8eUkYvCtZFzXfk8Vg6NAYKXpDl
cu8VjlwoLwCfI6eRuX8jqaUTIOzXOv+kQ7bPDdPEHN8ejRuEVDtOphDL8Idsl6pw
weg3LzDMh/UQAVmelIC72/eyyQKPNVkSHkixFqq8aQKXO9puoxWIjqo9YolYWKrb
5lK4OXolk36boyeCbIiAUQtwDI6oiob+XYRbTZVHmWf3Ng0J4sDgcChnc/Y+DjvU
UheGwRSw6FuhT/br7NsW5Hw+5bn7wQT3uUOJaRJ5UwNX/p8Cab9nQE/6IrH8pF1s
mPYNZRx84hLmJ74BvxnPceuptuN2M++X9NnSZsJq8XNx0pQAPpWrOFqkyDwc9BRJ
CvcXRHMwab6PDFvjUgDASQIk+18n6NT2wMqvZXpx4J8ROzMFR/xhSb8nfQwOJVLb
Z00fA85bm5nnOe4n5704CUNoUil52xLH/gMDl7pZygw2kaRamOuXrmSDg0EkDTls
Kj9MCoDddOUHS0S5qJaYIpMyQLogPSzxlp1rY0aM2CcDjkP0i/DDwF/nBp34iYN2
IVgN7bj07ZTSCypvqkZxclPOf8yag+LMk1o/QZjtafVHk54zBMX+vH/dkQrQ2j4F
NWeu8F2hQnB1OG2Ow6EabtIovZ4Ho3g9nh60CTFJmVrz59TcnLXkOoyTZ7M+T1w2
Im+u3h0z1MeuhE8TrahplG+zcJ6wNcFaHN4QpQsWc6/V2rhCk5IxNNTgZSBUQF88
OUDJ3gdjGzqs1W3Qljs6j3WuoCGt2JT+pGPhOOBZPnyQY2njf0Vouqs1iBnCvJHZ
jV6KSuxWm0VV1axyfeG48jsOlCvbYH48Ih6kZ/T3p47BCQ9t2XEFjWiKyNEXRB7/
CK880fDR3uV9TBd3osazJJVpXmuryojcgXwnPXO0Mq+LYkPChbi91QNLUO04VYNp
`protect END_PROTECTED
