`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mYmZSIMNvGh9UHaU0GRKpvMQwjjkyKIG6G4YJruVFK3m3i1eBIOKlywHAm2bhp7g
aEtes4baGWo5LuB7cvP+VsANHiv7DOVhepdJW2nIc7ctHk6f3BHobMUun1kHw/9a
bHsQVT0nhamGl3rXPhGWg2TR+k8yyGHwQUN/0VB+FMEajr2kpTB5r45PgWVQwife
ycqKcNAOgX3yVmT4XmJ4CROEtcTGi1t29iBkVOdrm+HGktAtmaoGzit07JOAA5A/
SJZ9D97eKsXEzvZXfYLSeM7vCUeiiBgI5J/0vldhtJQNtZRUkQ3tqidmgvjMFgsn
rmB0MaJxkl0qylyzyayFOpWg/xc0J6tyycFp5fzWE4C6AgR6boGtLv5Nl0WsmVhr
hAg3wmCDT8+gIr2MA2fexbLcj1JO1S6rcCU1VMq5sF6VYny/rlMG+Af4BBVL2X5G
b04sUADzv7d0S4k9KEGDhQ==
`protect END_PROTECTED
