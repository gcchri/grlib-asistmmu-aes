`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zQ5gSvEgtcT3E98XTf8WYsYi4JzgxQWctnLiaEK4rFRr1iPFcykFSAEaDJTWT+T5
09iLUDn+9LnOSebAf4qVr5D2HdUny/W5wvT5X7IfposbIEFVWZXHccwUJPmT/xum
Oy57R8p1s5NeCmCSqc2il88oI2UE7EcfNx5R38EC1z0jMTEHubgJ/cO6SGogj3sQ
2iuHC0gKu22P6GKIC++1IsNIJiwXTMaPqUcsEfjLeMTpXBCEes95SGVtBE/fUSm2
1E7AMmjBDfa7OtyofIJxzihjVz/anOUHmmSfUhDshE1glISQGPlhCHRg9F/u7gQF
WJZ5uT36wsRvK7rpovPNmi/U/k9vEK2wTSkWc6PSP7F+5cRNbzLl/FySszQ7R6LY
doi9htRMOBQqmpl5D1vT8+qPu0elmlAbLwzY0bpeTpS+9RaPRkipQJLmqWjhdUMs
3InOMYKmDVv4VAA0a2s4YgrICjfIAYIG6Clig2QTz3RCKEikXdYtwpXBSZzMSIbC
Y69nMxIVbbmJxWXYSDFA7fMfImHbXNLoo7B9eAmBSz5h2+c4C1qMc/zgGMCiC4+u
vJBKRfOEAgeJ+5DtEAmfj1FSlE59wZr1jwVfCBcv18O0NAcyIFhIpdE/nTjhJDbZ
p2QIci03L8g11dN+S52I/w==
`protect END_PROTECTED
