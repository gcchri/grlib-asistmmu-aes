`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zlnR3q9xdTatvb/2hDTqiOLbVKDIB4A7cMfV/I9ODaCzQ9iVelcuExsEv3K841tS
nayyK4E2ODiKSKF9boeIPGza1grrvE+KeqZMvhHECOyidSk8ghxZy9QEi0MkOCXo
onGP1Jk5tE4ODUSvyjOgLWAiAQjAj20423z6H5eis5XLMD9st6yEDGXlgpv2+JY5
hWolcCTHaIMAA7nkLmsApUxMAA7vlvlcO2cm1DuBkURwpvo9j2mae/LGfn6nZDAZ
4DFvsNrz9aGRtF4D06RILoTGCKyJArdcdNSJmu7FVydc7cSj/z7zbKus50BNTrLo
g8s8f6fAp4Lo5jmJZbn7zzh03e73YkH6Rh1ZjoAANtjeWqXroV3ChAtWv5gaoRXL
F0kfggbbiBNgqUfY24AoyNQ3lZ9Q0Vw6gtsnxtrUvuofhRCozbgszTUpThmZVZYl
6XLlCyY8H+F6TYrB9vqL10x1DmNBbZMfzWFNw4ST6jqu7dEJz15agjI+SDJJpxUt
mI4R5EazxciJoDvMwRWj/GojUdI6yByNDjCHgzu83hwtqOAgse5ml4scX2ELr59w
yn2nfC+sUSLt0o/R9qxTiQDaBAN3pyAVCRp9Qtv6rpL1fNVdEfWZGw0X+I1etR6y
RSpfR6VL6RzZNY0hp8fLVyJlWyboFn5XvNbPmEIEVtUjKiVn4myS5lV0rpAo6kDC
EZ8RSwfEVWpUtmpNLZBwAX0e4WRKSGMjrSqDE3E7KlePN72GQsnoC5WBpXWUy+wX
`protect END_PROTECTED
