`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cCnr/LixVftHP1P5Y9pMGrZvJHb+TyDzux8HYyWnRjFDpanou1m0s3czx6stJASg
CcNXk1ZYFSKKNsNtcM4GFaWrMi+zVQIZ/Apr9sX9rWMfJyR/k4sGmIZbBKq/kT0i
c2GDZEP5ODEBC5W/mwzLwH4p5we7uW5C7poY78Ezhep8/burlNGY+qvYax4RxFSA
UucnBrfDhdO5PVtig/xBJ6ovfMLRjHfOPmCSqO95OTdHnT7kXaPXzs5buDNCRGZB
7L0Nqd1y+xdY7VwPhDEhjsS4pPhiLeoppOQa+ahT8BnFkFnsAIHWLCms0EM5+XWb
FcUALgPwTU6Vr6xeSgPXq5MiUaABebMLeC9sPe1k2/++CITU/z8E28O2HbrCkztl
HcYZ/1Ys+tkFPCCamvWle0Qv29GayEXxMlYdsqWWEr/LA1+YbAknanBRt6SxJLUa
trciWNKbg5nx3MJDPhf0xVhIFpyqACvBAIyR8W6T20qpMNTNWkuw1al3s0acEE2C
pH7x0U11IjL0fuKhG3/l6BH1yZ0Olag8fWQD2buwTWBL+aihF0UjDU+t5RS5WVDx
yz8BeVLSKHn9O/JbELVmVOREc2a8cVb1mxXpigBR5KaCghWPihYAKedO5yDnuDJz
l+cIjPeAHC8plZUt9MR8nUXXDwSzOHV+jgQC4W7/ZuSRnObBATNrQW6aH9UzCeWF
Fmck3kt7xfbbZSF4rnRyvqihLZ9HArtZ8xdmvqAS34uPNs5vZ6UfoVlR0YXdOM4h
1kxHUaqNv6AN6IwLVCN1ZI0gHIedXRCHF4e8aoYU/pYjh6a/C2GcStdrm3qqDDVu
BT/m8sSEos6zhT1YzS/QP7WniEyT54uVimmkMA9g/cSNBaB3fw8slCEE7H/k/eNX
XoAuJphx5bOLVD7jxQfEZvyeJPNIh9i1scvJu11v1nw4KqfglFYhFHJiciezCuYd
/xJFSKUR32gZ+r2QdGBCVyK7NhdeYh1jIOMs/8aAD/FsldS5fBusGi3HeZx0lzKx
49qan7n/Y8iQWAhiMDiibxI5VshfswBtOUvE1c1urD1Ew6o96wXShCYbJmfp+R9g
ZPA0/DeCaFbhEa9XXxGIsCI4SZIb7jxLhA7Pjw2gBiDiwl6ozTsJdfvxE57/daZ/
5vGOPvBgEEbEdVReUPKsBHGKuxt7iuc/7NE8L5afq66xvYyqk5lFb2L9bjtfrwks
RnWLvCyOaQvnrj1CsOt110GaDZj0yA9eKzFm11vFeqIlcfTM1ah5qv0g1rCfE0rC
30yZHSIhw3N0K1DtN3PxEMSTf+zhlkArSYPcUBfkLsvgsRA7JLAL49TCoYPo+/kD
NEx0QQ4B1gu3l8D8BmI3CWdOZYbg8jD0jV3QjKwHkwPkNhtvpm93xVy3Hp6VWKwK
XFaTo8sCRg04MkQsoV+wfzlv1drWcRuQUS4YTR7J+O33q/hTQ5X3ooSbYmHksoU9
Pc9JLH6dzq9KWfrkkSJt6J0XQV+qoc+m/a3n4Ba9r/aPk9eGIGCBkgd4PfrtbPoL
HQzr3lSK0fisT71lBWIxRmm47G00LKCkj/JNQRonZPgbdakcY/48ljpAuQVcxWP8
l0PDIOxyMEl+26Y7YxMmkMZS4t5tRb2aTQlotkJhb3MY8Qg0O8VdYXfgXuPA9rl/
jh8qnEMsnroGWmqDXW+iAkXrSka5OjJ4a7KuXsCkckfdxg/wHewDWxub0Kj62JNl
Gs9gl6ks7w7Lmff3shQKPMBwXKt08PWoGiyiRLxFox//Nm5HldGFOnsomEE86tOM
cho7rSfV7F3fv4l+bQ17anT/FzGKTSS9BJJTTmLRuVbGrM3oS9k02S1Ix61xDC9K
pY/q+f1cVWK3pF5OrD/iMjYd+NAmUd3AONWX3QUImJEn0I3GAmWyU8JQswBvgWAm
TxZlcEaWpAFq1aFGsLEf6iHEaDrv0ERsc00SVC6S238dwD3so8PFK0gc5C2gEm+f
tWGdGinbXOjxG/jvbjOFWZalfWXFCl8kIiwMDFR/zF+IhxGon17cpIA3ks2Inf4v
M6//Js/PdN7+JET1IKcEJDt4tR5qVsWf4lmBGNIlJ9yXoDk8Y5yb91LwCN2epiWs
IdiBRxKF48lPa019UP0NTPFbw1PFS2HB7C0qnD2PoAnZi2H1BikxfeaenFnlC5wP
a5xArgPZ5HSLY6gmkp+p2McaG5gtOAhZlxyvp/bQ1MKDgOIkmK3UrXL54iLNTN2L
mMTnADrggDezTylYEauwX49pQAKTZOkL0LaY5svcsZJW5/reK8jHRfpuZQcQQkAU
a8qPSG7jPpzDsrZ2cFFphZrLBj7lNSh1sICE7wdoYwfh6YirBvYzfMpX9DaqfNWl
FfNSSyvwRXccboYHSfjpf32aZtKJAH1IzTPp4+5FGD0FzFJGJBBOuFxc9QNQQc8S
/Pjy+Tb5N2JmHnIJpMRrLNvUry6sAGL2rbzv8YxFpCIUocVf1taC3lx1Smkq9QUT
6neXvY0qkXxuPbwFCVQU8KxN7NvwaPCbiVqHCIrqHkMe0uGc1FZhaVXbATSTHqb/
W4bsOZuS5iMjpgexz1F0TKgzwVnmBm/OZ8QlzzzmI/nzabjVFRWuuJs+8Ex9mShV
8gsx/3njMsoZC4KRnZaLqJPnGx5XlxNl1YuSUXMEo/WSE3ly2WQjMzKhywmrseKg
8PdUhAt15FShvfg3QTnqsxcMZqFhsGUa/bkLzuyTsOVHtZGgO2bVjdgFOaR3W9jy
8BZhBkEJ7ibJb0WMPiC0YiHfLgVWRRz1RSCDhCja2lZz2iBzkmX13DHXbhwnDYAV
bxUyk4Y1eNfzQ56oXo8uMg9JZ12my79x3MLWrg2Pwv8U5r6d5I+V0hppzwbEqKA5
M5oa+u6HtbKgp0jajyDXM55zzjQn+S8h4mEdi1qLAo97xZiR5kTdAjKlYsJg/owE
3QLFb89gWg7zx10bb2/zof0Nec0sX+jlvi3e90QgxRc8IZwKjMOIg1J7zHcfXHT5
YZI+/0DKW2qn1QKDEWFlLWsSfSDyARH9sZvkV/4/O1lBb0w+ANfUIHMYIAx+ZVZA
NQ0S9jfvQ308Xi61S/bgDSXqhqvmV/3/dYgmUo/mTtntJxO8xUwzHy28LxzyrAQt
EbKl7YPbFpNjPf4Y9PkgUgAd0d0inDwklF9pTPkVbH6H/kBNoyrPEFUYv3MKS4D8
wMOqw8kDtLzWUdC1f8zuZ5Uq1m/GZ8gS2Iz2wzGqBuQRDlrEQxki4Kh4WIqJuWA1
RhduYXbO+Na/eMtrMYx0SRPW7dEsEQ2kVe7Ew4ssmXrxrJG3fOhYfnIdDtwGt9tU
k/t7sNoeY8c69VdSUmFeDQ==
`protect END_PROTECTED
