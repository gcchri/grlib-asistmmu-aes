`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oiPityNGTnGf25UWaISD8hxL3222BnWxkFqO0+BiljMoeBMwbqo+xK96RcwdUnEE
8SLWOROrHhWgMsvAAfdF56CvTaFfhY7tXlQAcS7w7oods2rJ2FYp6or4NM9ad/J0
uhqzz8jiBbL/gpz3mcVw1bXoCcYRBgOC7fkM0W27HquMzJCBi+FWmP8isalcklam
YWpWONhzOaVHnJk5kufY8zcT5cq6Of2pfuUtCQ0F8qNfUkd2aHvX9ORINsoPStcl
`protect END_PROTECTED
