`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
inRWGcxOf3XxuxSKoc7S+/KnDX9xyae7sZIBOVw41gx89HiUk4wmcgdtPqDB/xBy
VeZl07ZxiX+q4rlASmHtQtTtVp9ELBT9JCvQDZvzBi8tAEdb/kRGEuSCEHiKAVp2
JKWJh1XbXkdeUfDP2aNI9h76ugOps37CXbEaKye2kUbU05wHBKRnaqb4lDxlEcHT
CtZArn4GJOlD2mf1E8TigYG1TH+dRKCJ6oAhlDD6Q7b/5sZSleeG08vcQYKM4zGA
trPCi5w/a/Zyoyijp7TzverFN+46yoqzsOq9i9YxYGGocB+zaI/1yrOQh4BAQaiB
WedKRl4nbv5abIbrtHD6ATPxtFsHBdZJ9GeDw3k+NqBSI9mpNy9/5LTBffIhyFtg
mIHi7C2/Gz0BL8WVo0o/3ZkfBYDuwl/JAHGYS39qhcY=
`protect END_PROTECTED
