`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1RM4KShULgOCY8mGOwopB7emYfiLPr4h7urVT+yDzJrEj4n9PoLwsjk9pDihZo64
HB7r/Vz+x5+GbmbhCglss22caH/CMbSpn0vZZUZnJH01yeDX9s5pVKStX5PsNqzm
ST5DLwt0fGuQs5qO0ZkKJPhUlhmy53vWlrVY5z7uQdHOisU0lIfmsJjaHHe1dI1U
rypvTNX995knvgRtJLHOclPtWh8Icrms8d6O1ItNfIbv1RgcHBwcrVXp4jZ6IjhS
g9q8vePC5G+ZLAKNGmGluPFShBwIfnp4JE4T9wUhLonihM7Q1RCXE4W6BZjGVvmd
sA7RCLnD9nZKeqfa+z+CT3r2Oz7hFmphWi83sgDyw4m5pPJG11krCEr3kZEHG0LI
nSYix3omfNGybQWDkXwF+0ZkJ/f5Xe4x85LMh6YmbJ0=
`protect END_PROTECTED
