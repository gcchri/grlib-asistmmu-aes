`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KBgQ4RHmSwrmE8rVp5ADc2nEu5HFG+2ufM1NrjZVQmlWDYbxfqFAoENew6CWTewN
EkNr/vBiaVx7bDViT5bX7oTlD2r0hnr7RdLFcrRbgMv+i97LPALtm0vSmmK20pY/
QJHULphlEAwoZMat4f3OgGhVlnvljtHh4TSO6xS59FtnKb1S9Zm+VBpKuodFNArC
/rvS03i83PC85aRBHSRDnVxNiAjyQU74uusE3smgSI2FDgBwqft3QuuiYSQISTvF
zfJXijojG/gdv8ht2V3UWDpNzat39kUuIwpVOCkQUsAxWvakTH4V09GvwAblpf63
dPeKVHZcaY4wSLnJnUIeo75Bk7UbIBl/EpbJixBPLAo1+XDl9GZow7OXMxdlNAh8
0WnUHiky6H1sL1lYF6XGFgsjpFt5S6T6N/B9Rqot0WT90MHqY3OpC1nyDll27O1C
`protect END_PROTECTED
