`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iP10nueOdZge5UDQX/Md4qedktncxa2CLQ95TVeWQ5o+BMfkTROnLg2z/16wLm4L
R6AAy6WiNZaTJlFIDlp8m5+NcKM9xG/lk6wyJvDHAIbpBn01c9yYmVHUO9AYbE5m
SUUyW+megvZAQgKWvEX9s5BW7yp/zsY+FGgTsrmHZoIoBoI8A1VE0i1RGVUoaDsV
0mpftkh0D107hMCHYtGFs60QdEjKsbMCRCrJw+9xWR8zGCd/4mjjSMu7qDpMyyR3
34o4OubaO2Yb0GvcmANLCYXjiwcW6AZiqmSFd6/3JB1bsttTgBYnIrJQxftjXjeU
UF0A4raNfKjTWv4RAfi26jYx/Y4YaJ0REIawAp+kK1C/yJk0AgNkmCoBkV6f/5RH
bcPntwIewM6z/PxWbAUup4XXuPUjaRfFPp0Dwg83jULrBS+BppjkdjT/X9E5RZQJ
MWvLyxFb9ZPUkZzJ7gPrXbkN2hM8W8V+lI7yh2TauJlAieZpwZQE/vMV1cfrf8dF
2mpE7x/MXl+kUyLqrkX2G9h0t4ddDu69KJkxHpqIxONRPCdA63OfKX7i0gzmv61v
NbyLxoVQWt645sbMu4pDn+ywssqOaxgoZ/AAgHCc0r1jIOENT5+epKJs9qkxL93E
+no1EjH2aiULfvugHzT3PaqC2YuKyFkP9JC2uWhQgxxQy2dGG9haf5rrZuoAKQ0g
nq7mk0JNrTEAGOt2lzvAUTi9m/2QwsBzxZf2kr85pYWMxsOqT9SF2MFo1wZuxzTe
OlFylYLNaQAGDNA5apWKXc6WgSL41TdapBT0Jw7FgHQKdUOeUdCKeDUtrv2o/AIQ
2QZBhqXdNyLmNLLCxlHrsFCbnHV/t/yKMA1dU2En1h3cPp2v0p48wrh+Pk3ulHZa
5ZQM/hfPF/WWHjng7LJes5Dw6pFsOmY1JBxnzbjskTS6tvBUuEKHotvA+PNIurUS
JFlvrQGOYlg158G9TfGQXIRjCkDA4cYhu+yHuKub6kZnViwYw/yk82u+h/qDNafG
GbhPVMnbawhIcRWKCy97OxGFvUR171KRje8a+m7fLBwdJE7EYC4F3/uvP5pKd/r0
b0PTo/NNzJEX5PJcDX/sGSQHmQ64BOIXI32l7bItvjqgKe0JP++3WNDtm+0sPXB5
U7xaGp8/gkWHiVHmzr7IVxHgRo7oT+GE5ZuBb5KTS225quq1sMk590evc4oDwo01
xpgyIWMY83cijK/ghcGVHaJfBO/+ivnLCcFfX9Q30InPjB8DrdL+IV+G9MSLNEHa
2MGtJV1Ks7UpHC9keW2Ptk8cbK91eMYme5a1LsyMqvTrHrXwz609frAF/IqkG73P
9FAm3JEAIo3Vw8jbGdpT2a4yCf91sFuvdsjCfqJHIcCSMedceNI8cC6yGILq8NQz
Dl02ruZk63WYzEnlVBOuoKdY4NzvWfoFPXDBreKU9CvfWYkZUH77KNapAA/k7fwM
8YtaFpj4wUU5N3Ban8uht6Jx5WiOYR8ua5pjGE/nopL+Z3NSt3JkBvFEqK7OOTE7
8JexN/nQX1gQ2onP8C3X9K6V3dlwhmSbW5ypO1OoWr2UmthQIsjAQJtjhDtk/Nm5
2xmiXN6lQ1dklP353dgnW8jkkXZeKBJgRy3FH4zHyi6GSluWsn5PUvHBtbsmxVW5
wTY7ZfEQE77RTrNxjf5lKAmBnmNjs0VuIX7k3o8SN10mY3Md85WWJdjsaQxoDJlZ
H9d+pdK94XDed5WktZFtZZy3FDLRhOLj4aeUMw07mjI4TT320ylP8XuAeTUk6+xM
pAZQGN4SYMtmt0yVPqR6ixWUoqDziaOrsMyoBzQfUIh0Eppl9r3FGkNn5XS8xT/E
4ljsVyJBNxluHpOneZMHXuic0vvZhMafaLxido0qiUMENj7MGuDiOGiAGGyGtWet
ZVMU/yKJJAWjPcM5ys1Pkw0DoHIlUSfPaudiMWXfz7SbmTfTxLpeQ/YRmy8WCtrn
nUhRbJtsRTlivxcplgZIqkRPidv+GpbCuAy2+FjCev96S4ENg9UBdmHVqe9oHaMU
jjeVLwfxsnYXcVwHAiOfhIENq1SpTrt408Y3/QqpH7uxxLJGqx/3ztH4F6kDe0CG
vizHM+zBwhjP122WctaaDy6a4ihWFGD5FQX+Eg029MCJHH0HukC0xTvxXklxP6Kp
gdaII9TfRVl9C7qgvnnPJSuoZpuGnu/PuiIP1+oZlO8COpY75PL6j2OOPkWFbMlm
s1zTTNYiR0gXZzonQTN1JeQvNyoEmMsEWfQ3GgBhm12/6r9UXUt/DH9UELFYT4cf
Fow+gHSjcAGwqD0Dd08S21rZP7W8WXAjvTwYHF5yDnzARHPowjPC0PHlCuAl9Ll4
4REwwRJ1lqj2/B15QpPMfbT/oKSca7oagW6jnXWsrdVDAiofIPGZSV/QCB3sl8/0
bcCFd7kFvoH6sjtdLgeF5d63t2TDY1Gaqqg/DFD/KzL09MgSKKEGVEfYleTW1iRN
K51NWJw8mou09vcP2SfIJB/T3VGiq6mBmiQtwOp2CLXxmTO89brVn+Dv6fu4hKCf
Yw4OT2AGkp1eR7SlPvylYNPA0qhI71Z5Cvtv5r+/678EGvVHxTeyku6IxmgGFm8C
ZJe5igDoQQEy6sA5l1MoKtDxKv7EJNtxWmf6tjHmgUXFOHd0hjQ94vCBa/sGe/vD
XWpSdyvHDzLognZMC7wwaB1q77h0UW+n3exu13UOisYtSKZ6oNpIM+L7lbXFYbri
bIDkkAeYb2AWhPGw6kWIDKp+esATOcMIk08V4W0UyQcutHgKhD1xM/tmlbSTmkJf
bGbDbMlYJQ7K65VqUEnvXF6peNnImuYxhX4OmQSgvw7xqJcIzTc94rDK9tEaOWLP
4yLoa8VWF1RZVwXBvfgWMdJn89Eajfr5fgqZVFEaTXkWEjW+fZx2NM372yg04uz4
CLMbFQ1n2qj50FrNYzhlzGBuLhhMfjovd+Oo9kJgrbZOwrMf9NdIZ70qagbKKuUH
6BKftFNS8wJfZ0YCRXgR46cKlWY9xXrl3gSn11gumwC6kQoSXlAIBi4W3pQ6rwkL
FrLNq5IfE9snNJxoWVAYSbuRXoLhcPzhd5ao/y79D7gS9KFyp23usyBVN3aqh/3i
2PmLMP/Rlzi/PHVbO0f2137iT8+vdq65jik5aHS4jTEXzhv5aRiIck78paqZGFXs
1Qlnq75PH45+77D3AaHedvoErq0qN8nixSh+jC7eoz3jhF1ibMOyzz2z2xlV+nix
JDrjowMW0Fz3mNSZwUdBt52ahdDiNQgAw1M+7HzWvM0veyw52iIF7/6ENOny72fQ
yeLpy57ooQXTL9hnZmA1Cqp9GxcYI1n3GkhmbohILXDG/M1e2PSjuu8Bk37MDCV+
JGV7EfEGnhQcyxyZnZ0T2BwfZhJf/LFYvYfko9kJvRqUoIS5sx07uxcoXnf3YAZX
IiaOdiuXThClGTN7Fi/0zwWDE+AA40Zjqw7IGotah+bbFam9h6pbsj/dN79OYimO
sjZB9p+B90VBYNZ+pfyd13TjqsAOpnneBNP6zvuCt9FgZLtCgEOVmFlodpkyNCln
O9CeN8Y64YKYVtAlynAWCMMnWkC/KK2JsvuWYYxuarrkmz+kSM1zIFhOO1t9/GAw
NZ1Nz01UaORrSGrqyQOrkCb3seKxaHD4nYoBKQXUB7S0vRfK6R2AIrrP3eTfloLU
QMXKD4RIDBfy0MsLLF5E6Jd/CpGkqYeVvhYQMdMzXPWwgsBwVgbwRvQqh1uGIh7q
6tlG5uhuVjWfkEI/YQB65UadXCOf4oGx/8tKPQD7jzMIhbW67ftowKucqoFEaus7
YtDpal0f59fP+OmvhByi1By1kEhjDYXpCLN/+sr4nT/ioX3Kml9yOi128wr4mvsX
Xe1nXNtmtVstieQPpNWQ6eEW+wHVbpNVhpmKNQ/4lOY4gEWWlRkW730PEckXDgEi
RRZhjmUICADxjvuJ97POHHA4nYZXXh/r98rEES+zIjzzzYedvpqm7qjcZQLUwyIF
Oe4iLrLOWPskZwvcwk6cqjKNP07+Dcncwov0eTq7MQThxQYeQZ1fVGmPSSG0sgp8
6JP1y9sD6TDPamPVzKt02TSmQlwNr0IEAxTqEqZAWFD5blDxg3rBEv+XeIzkBgr8
j4tC5hHqfheEEifVo4ensYe+IZiWc9LjGR6K5dOuuLph/XAjpoiYCjJil0BRD804
GC+JyKqltHrA+c3U2/W4arVKNAE+luFj7g0p4cMRa3zK0RwoRykXexyPu1MJEazY
g2XIV6Lv+N7Yt//CYpaCOOwwZi8TPx5Ty6dRKxPiV4HjgUizxy6F/J4TTdtPaREy
Ygh96o5XG8HjXRIqNyYUELk/7wtGsmbCapHRuisZ1lIDFy4ZX04F4KKQesoCTkwN
fo1QdsDZt8mcXCmQR/qf/XOHK8pEGIVNxIbLr42GFmd4ce5n5gnMBDyKYQGwv+Z4
1srKhsdyjMrjp1vbEpECaEU3O8Y0L6CBNRnZJxFJ/7MEdECorVAjCdMOGZ2LAgpt
4ofkZcOpDpDnxPWdAOxnLK8z3BBLMfiDC9Y5/10qmA1pBI7LS6NUf3bPoaRK2Q4a
8voCk11h256utVK8i+vq9v+sXDYDCFRV6DcTZNagrOCV/RkLF8OHR8k/kzC9QQF6
a8yqA8eOFlwT7KVm7ZMYMoh5i2fQDPW/6VVi2XEYt+gfHL5zIB/LZgu58z+cnClk
gASGjTsaCloxzz7taDijfLQA1cbkRaxWrnJ0CW1JY7E/1e6QPjle6n9uvRfl3Cuh
jQDIhe/3VP5uXEqEDzuX74IboyAEcNDp/hdIgtsKGYJjgfjRUbvewzCBYZm4wsig
gPzciBMOSausMjS4WWi0AsqM4rpTDcW569nIvH6b5hzQUffGI/xgjwILhpwTN38d
bRAxpPMLUp8jeHP14tzd6v17Mxiol4DaFE12AqPPiqYKvw9UJJ0AkB7efElviVog
rLPXybM+P9z+FcgQY9QsND5dhOFjnKAiRe8X29XmaaGGA+8pWfdJH+oRLRafTzJN
Yw/P46r2lz2BnWeL7WFKlPs1bqOgTVfa12wvCtzon6LCp7qq3OhhwrBQQpMnrjsj
0pYNmtb6iFP3n0G4ZpTsUHqNbF8b7LPGuF7dV3N5WCsVIP7b4M5AN9NnF1eefsTk
OGN/isvrwZSOuA7Hx9XQt+oLJHllIMcpcqUkDYhn/KamaVvLv9bRxa0cMm42JIyN
N96gmsoK+IjtvOVB8SQZv2azgc8wjujyrhaAqbeU84hdasnH7lzehfU2gsMpmHZw
MDCUCsXMwdhKj7NBHA6aK39nxZakyMix9o07udLuScPZTAPuDN23BUPLKMXIRVem
IIAfYQN+BAA3YVS7a7VGfQ5wjcvcg4GcboRVQEYL5aBgaNV8pDr7L7udYLm120ey
Vwa7yIEmFaYMNbE22RJVe4KOk9WhcyQqhziZBZSuEqqTVpQiSnMogTuTihZiBrIm
yaFbptpMVNGJapqqYaRTnMQLimqS4hE9oKfgOnKmxykMYmJOBBEkAIrRIRq4ef46
kng0kH4EWV+BHUVE8yqPyWOTZucqsGEUUDDGuGrK5V2ZV+B/Pa0Uf0X6rgYcdSvQ
ZqlVgCaoYI6Qko3DtNgoETjfPcQzdhJA6clkJHn6ulyf8QWHgdYHz6YDSc3pD6Ut
XpQULA5muvubTymzaax1S0y6ZyQoKO6Yv5Bxhx8FkQUCEfK1jN9qPGxRkl9XiELa
EVQq86kenmVdsijJHpNX/Z4RSZ1Gxb4mH3Cm0GQnLavbGS0Z6qYrX9Q+Oy4CasCc
cj2d+UbRdi/W3nHFpvXeJG05/A6ufdhyBJ0eMsU5f+tREvGKsQNN9czCnDPk1G1Z
qrKKWmFkvAWcd/L0/ggLgHPwHInxhLPDFlqekMoR8HQVPgx/q1nrCy9POs+HO9Ko
Z/AxpaDooAp9PrrBlMJtVgfYTTWf6E5fd5ByhA1Q/S+naysX75w/yUgth7ba/fIj
2bviVf7brG9+ZUY1dAh1+qE1Qw2BXu9BWCpOgofuMhQ0X1eoRWX5zg9wbpXk9CoK
K2N8l2qe6osCF+OlbHAU/mwzt6yNYz2nbxciAOwZQ6mZftSM5hu7jvM/wkQx4D5C
BIy1kbPr2QFcmWJQd5pVB0BrGaCi21c8JVFBJU2jQ2WYKLRBcpJ0QTIOhKQh3YDk
0bO5e8crBHj2rL8uZk4fvVqCsvY+ftNk8hj1W5o3Yt8rIp+15IjuIvBGh3rdZT2C
my6XdALFgjLJrUFu2WWRshXGnPNeykqzz8GeB6FVQd5jrRQ8Sc3MQiFopZ8kW+GD
huDjH6akKC4fHryrtHVI5UDiV51qqGXyqHCdsBVBCEQHkAIxw2D53I692NhJB3BW
gw5PJNOmVVT7KPpIHHFrnPHxeNsgYCog+hlTO0pWvGp/lrXK9Dg/SjLsnZPqXSjL
JxmccjTXQbZzu9DDKEZ2Csj5zXbqEMZxKaWqlpG+qhFmNOOuXNrvEsicv4BXzoin
SsSY6VVdV/Z2GzdjX+z+FnAJ7uIHIS/lRTZdNBxRCYgOAVTkilDQVzLealm/l35w
dq1zPPBKhWGziECaEsH7vS/l1HUHgu9bjeZNjhp9MgPVZuSiqCID6IpbvgYIPivO
EtqzPHck4RypvjEG7jlrlA==
`protect END_PROTECTED
