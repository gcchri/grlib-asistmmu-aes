`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lmCCEPjpE+DApo4DsJeiRIaJwtPr5k0ZUkrYNbNEj83ETK/cVIF0cVLxwGb87kzn
E0RDsHdb3zvnYzFgcnSseqcNQryofgmz8j6rz1d7J8p8AVSK6vWpiGFBsaaZO2Go
snxBpsahsMIZ/u6CvngWBi2ubni26wU1RTwbYcODHM2CR5Akd9urcjSIMz5YRLPl
UdzWfGrbdChF7nvQ49312nQjbsaDAKiBHpdbeaVDA9D+lvzdndIBFX7ATlCSBmci
uVIMUB7oRXK9X2Ebu8NN2Dxyh9Ve+45fC4rhNllAkkmPaVXJ9C0ALUBGgcUDIP7C
h7mc3h+eCpIy2KBJcBotazMr0yU/QHMAilgV39kRrSll45Nf/0F1qVXztQxSsDOF
NTUxZ/TIJ13PqFWHa2B92WoOkjZ0RTge8FRncRuPa1j5qhnYP4uDsas2ZVqoSY3H
Dw4C5krIw9hBtFREYAdYZfDNXD9lzN5BrjZIiysJpCI5qAIvuU9UWJKwBP6t6uA4
KNb2WCHhErg5QE1a5Ewhfo5abIyeaYL6zsYe9d7kFS3FwKsd1DHUNE3bLLkQ0WzR
7CsPEq8KUAgx/QDOzoozukDkUmTCPu9rUtnRc78BUSQRMJgqL3bnDfcSon4gq1mX
P40uYb3FyMvyMcSlCfrvbmfiv24CqLMYygvBvFmwqzfHX/0WgmSXG5KiooJs1TsT
dlpEDLl6aycSYwVISOCC2AwymRi3I+4n0M04X2+NOY0AetoUpyClQF6CkfBfLHYV
5tOuzLs3Q1faNYdvhMOcrOpO7fooYgvqKnxlpfQyK7JntEvVuzfDom77qbNZlzF5
GpqgZWgoaaog9UJf9siJURp0pVPYkNMkww3clfRVCmDhovok8/Tffg7tAhcPXT0l
DTL60HWrNjZKcZspt40mZ/SFlxImSlqbBUj5lx6gZ2UlNLD237j0HR0njDuc0NLd
kLnh64Z9otYP7YdaQ1dcw/wJlRFwcK4rKC90kq0/bNwlGMMhbeBGgMqCP9qLMYsh
ZLBjIb3BOG8qRB0hUgUTkVjzj8meYLGVA5LeQphvjrE54sLVWTVZu86iGi5XxhxL
xUPrdWzroQCY21F/gHaLGfC9dEmn6WTWVOF1orkuwBFH9LxbYrYEAijVsdz7ECX2
xjWcwtcjXYBmGIClYGIzpnLvyay7lWZMYrdii2Oj3KP/EdeGsCI7lkOzL60HInQt
+tCQkqnJv1raghy5wOXiBznFW3VexIqqEetsg2zqOifuMtJRNfiB734DHeJNfcwm
BszQ9XCP0gOC35HMvyX0VQ932pi04dHAexTG/f2SS2CQ9qk1LQ2YAOOMlTXgdVOA
NM9R8HO8sA99vOIw6Zp247vgmJ2+8ReeMrrWGS+LEUOTJoKBODuF/PxVcV4UWPL4
LWFfq60PQdLNQSAOIUf7xmBAc2y8bBRby+y+mVn+bhU4WsImi12IgpQ9Edfqvtsp
`protect END_PROTECTED
