`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a4JvzKALJHBr533OL+64dCf1Wj5gp5atLHJ//Cij4GK1kjg7TtRWAjU14QPVOShv
uL6idQLgaOOd9SLdFq4PQennjA4+csYG4d0I50u9fjZ8Ezkb0MnfoaO4uDDm/Ard
6V0lj7oXYm3sRxj1rkNWdHjQ7ywe2XmdDVSoR5JdnV7+eFDvAHKnLlmpYwEXpStR
+0+NBltutVQzwdZrUvsywN+c19UD1roM26ZSmu7xCbcX3TVeaCpszTm8YcPiP4La
wcWOBXN/BD8mjyDrkWp7fXqbzmxo6eGMd888+N7zb6IYaefDwkTpGJCJ2UoYaJO4
bNzthIbWr4JGmcIaPTf9ojn9fS8KTAoW8FZ9lYFuA5USl6bQNNV8A3H5IYcvHgqa
4aFYANN0BcZ0+6Q4xfBWOxS6i8y/lstO/ctmAPRCpB0JoJw7SxTwaB8kVRJsoSq/
m38mtYYFUJtT9teiRVOAO5XRgVfsdWo+C0N2S4ezRqV2bNHDzbeT91e9hUsewaZQ
YeyQFGAbz89OUaDLGU5rJT/uzZaMBAy8R3gcOr60414b1fElv+q6TDBurwL5EUII
`protect END_PROTECTED
