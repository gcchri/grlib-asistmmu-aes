`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oA302A2MrSo33KraoxW+lac9fs7oTC2MM4lXDWWReVTPfkyyUo/JQTGPOwdcADy0
T2WNIbnrOEoOYpu4vY1ZfoGomWRVPktyF2319JESke7Dt+70S10/GbxwtKi2IbiU
B1FuiXn0hF3n/4iyei97GcjwzgHZaa0CwOo6WY1qq/C44RbRCJD9dDGKpEmMpmhI
W7cvgqk0/cM9nZBCHaK43qrC2NahN7PvIGiIq723HQ2aoykj71b6KD16QE6qnn2V
NKgeTBgjmRmGztMEZLoKDA==
`protect END_PROTECTED
