`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IAr2jBmH7XoOf4E3VkfCOPjmmW8/L4XhyONnOjbyV1Is+ZIO3oARaQKN/80/ud69
Qf0qr4ThPnp04JitvuNGEFra5TP9DGLxhpccPL6FaqEHZVY+xExv5NH1QME4go7d
5qj6iQJA8juT5/9pZvzn+xO+sX/9/pKF/WKZ4ZfI4+ogSwsVkNYZ3FoiJdYWU6ZC
w/kcCsEt/BQmQqLUodd4Fb5yVRcX6gLLgoPSieRmF1joJCrVdkSWleu6CR0oz0TB
2C7brLb9u0w9Io3JlgL7dwKeyFtd2gawJ3m30BQ11aTdT693x5CZbYEgmTylrjM+
EmlN/FF11mU/VR8aRX+0lr9yKCXbQbueukjRvrFKU+hACWWWjqO0PeuEhlfgX0Zf
MLQVJCnln3AgKwTNZ7e0+Eg53kVPXNarb9RPoTtxaqG7RiNabv57k54II6sY8Sdr
MQVzd2xOCZyFsOavSZLeZyJcygqn0D0Q5Ee0zEFBa20oAsRdd2NNpex+/1F0ELC+
crm+OvC4x4MnF0bzjp2fbrYmM4EqLq/8UJOP9inQ5E8sVNQw9VYzgFvaDUR/oLVg
ZiscqSxehX2eOkI/rUfgWDcBwaft1HwhPnkcckkoOGK61wxicAtM/3NqXPb9WhP0
nWIvbImgCrEXWfzHXGzd+bLdnMe0h+QFyyMMuF9lJ1UyZhq01m18Llalezd3o1/B
cln7W5AI27YLay6Kiyv9bZTIFGomRYxZ/ITWtbgsge2K37lXSh2YeOmUhr1FkScb
LDPzI09F6EIfwo9iFo1NZVltqIOQajmFj1XHdHBauvSsT70l5Ak1gAQS7JZoChpG
Sfvdj4db5OfXikLO+CjZTcCO3KBrsHm9MN0eD6ibw4S3KY3AMPgDTm5YuDVIb3k0
ptdVq9PkZeD3Xej7JMKiV1ZxYdIEKq57yzgwvYBMVgIJfdqAMl4BppngvoVn3RzT
0tC0LeoKdogdGtLwuU02PfpAMbSsRK2i5o/SiFAeNh7E+NIz11x5nL20ewAJDFyW
1jCDHWk7FWZt2tZrvZ1+njnAcuq+0PDYiu3/Dl7YmGexJVZso9Cg1TpexUeRUBGt
UVkZoglOLUqD19JLpDz8liJedgnVPes6wNVIBVSAk9rD4OFM3ODFtHZfDn+X7NNi
Ce0WWfH7OifyGfGS7Nt8zsOlrv5tD7BAMkRkKKSDEVciLN1te91hRUH9wW9Xn225
vfcVrVfFwkBEwcgQn7Jcmvz2jvvl+V/JjS5bK1lA52SHxu93YhudD3Lhk+SQIY/G
LrYklOmwKajbBdupKgMS3SpLjMCRBTgiDIMHILiLcVZ01OaPvxYpwKmaf/WjN0oz
htZK6/2YIiqu79WDB7ZVUNh4mvJO5RdOvarBkiYXj2fGPll2dxDc4cOknIDMeAJB
B0PiZhbAeVQhL6RXQJZJBT2NmxKwwB1pUAviQRqV+PpCnQva9pgx9E8H8w7glsYx
GolegFaYYmHnSCRhpm9nrUfTxoYZ/kd71G9i2/kHzAO/icqoNDlqhM7TUheXQ8sw
dMVI7Ak897irw2qsfKwp8v6PlzyL3DGqDrBnvFrJll+zHSwyslGO6dmInuTvuAXl
TSF7CEpWKZkYK6zDVvrHAoFyT7DqaM9VKUMtYhweR1TquwD9CTb8SxYgMrwlDSm/
iajc0tgjsZ04Soxz/jwZNmvXZ35+AZ+P9x//x9o2z+8crlaTlbZXuH5BZcJ83mYC
rs1bG/BdCPj704B/y68PH1TNbDY99ftkW5Kz4NxYxV6tsi8iw0+HDT3snHRxA+Dh
z3p/ujw3Ni6V8ex94KDl1jCpk6SMPkmWMvnNKd6+pFyUey/f4F3d+T/OFngAVSS0
e6xTzwIfHcXW5aT1NU5NxWoLPvmBhlqlgkjbH25KttetjMd6oB6lrOo3VYec2A0Q
YHrBcxcxdeq/1sXCPib4QgDG/lfPdL06Utc8c2CQ0wCLEp/BfGAR+o9ax5OivKY3
6wk13PIbhDLWDpjevO1c3G8B/gCFO0SMAEJ334hJf6dtYD4XmVVrXofcA5TGO0Xy
c3WTbnMUDyIWsqHse1rIA4zLPrja7PtBKEJ8Q6blnewn7SdeaACgNI9pt4uvUNLn
OYKtrx8bjzjyWUz45uUnHy66b7Me1zeVfd8ZSeu4241GMSqUT1ZGhm2bEJ+eNl2y
Lr97gE8G2+udLLZDr30p8d04HBxtXtOvJIcdBVbncJF3aYeR8CQGECuLc0JHtZmq
8xN6VZjckjiLa9ft4R/97s+8tEYNP0n0BVDqympw3gVZwC9bfXdib9F0gnqJpTnB
8/Dd9aUj1oW/7qTKV2LA9v5qKV213a0ez3FHO72+w6pixWOzdvwWkxlAvsUWtr2M
PQLFq0gYExRmGGShpddIpqTH0adBzWA8Glr71rxL9P8m8pR7e4KOcK7ekBhBm1b2
TjFZQ79Cc4m/RCPipAvu+/3I/83MWB1x99z97Bztx1li9hg8EbJ9rQii3HMePcIs
+IshBq20gY5ApTDpa5i/Qt9/Gr2a2Xdh4IW59cEI/Ei+6cvoM+EowVcYPCMSNerj
rbYGcd1NK+cRPfxhpOqFW1CuaSdVCii84xwE3nraTzEo+EXe6rVbufU3w7AvGOdK
Gy3wcof9W6nivxeRNlTRYxAsujkZRft6O6DBGrlli+7c6H6CQx/tXgpS4EUFMhCa
KS4dKuIeSP1sofg8FOp+wLR+SFLh3hX3Ul4IHqZSa4hA4QJO0c6xCD6SpMqFHqZK
YnTdV3hyRAyvsv87MFdEDensr8KdntI5vCP136ezoqUsdT+4e66ax+ZgHkLtObgk
voNUZ+DrY1FldwGLvoUZbS/aazZ6u6bNjgNPQoivOIVb41YdLxsiGTPkCxnjMS8P
D01rh3CRxTrlPxOB9+PPfwU7TJBcFgdZAkGN9fsUc3GY4Sp+csZoU5bo6SgfyrZ+
IJd0Ql8jsyEesOnyd/EmX4EsnJvcoYZ6+vxCbr7of8OLyWGD1f5mpKyYcxBvwQuT
Eb7qJ0W14GbYIMnw4ZnhqoGiqkrbhMGyetY2sOyMRtoH+6cS9sz3pZmC6M65FKay
TOX6tpP5yY0WE4jnT4jQb1sJ9nDp3Sr/haD7vIQU/8MCmKP+uIktq4VyBbU3wytF
nPEMoBsCOOQ4SP/2YvcZ70Ahl/BAeG5QFYBQIMg+oMb038CqvfETQFg+zxr9gzAT
uPmuOK28qpcuvZ4FrcFXCC5bc2P1FoNXdUnyZ5/Dp1XYn4n64O4Dsk4f/Plynjk+
17ohGBPC86P4CTLdYc/uKlrruE2B+P68AHg1IMqUZYxqOTXjBhNBEI44MXiT7pkI
Ui+06+PMWsyH3p9MhyZITjQh87YIARdyn+RdECvuTktuYzsA/7qmx6o+rHGPkQHv
3WWLiKkwLQvSol3ccz/cdW5647aerOJSzgHA7XHANspCSLCCN3JW0+pobpSsBC98
kb4ezhIjfhDfXAhOtgXkvtdpTZKUl/ZcwOC3DoCTMPUvH5CugYnl51vIR3dImnpF
J0ZkinuadkVyesKZsnNmjLMfJ3qnlNykRMUrseKDoZvAlP585wF417Ks+fdi1CO6
XovcqMq8L5cKcmcXzSQ09g+49Bm15dbJXTbiQeYlF8Kf6hZEoEADd0RKi/BcumXW
H/o0FjSwOUxh4NPHst3G8FFbiF1595xOSV0SGMCLpZcgbCCOZe1tEUZ7G/0BugXj
NU+4xd/NLQshv9z1XHuWHMQ0f6RgZxKZNx9e3/WSvJ2k4gwlCY2IVUxxl5m2U/hI
e0/aqydqeMP2aPROZESAhtoGETm/WvEqGn6BAgEbbUrZBhGlvkoi86/K54dcimSO
QhuPqw3LRjGUjU6aQ1zTZ9rCWCeKpP66xfZpiYvGfxT2TjzqglLcDThy/4YIyeKa
PJF2A004RTHEu7znQt6uC2DhWT8CfHc7uV42PJbTmSpSD0ok3icpu0Iq3aAwk7fP
q8pbqvsKcc/P4FvzxUOyy9wWf7LiZfvEXwxQLZvAj/ffUHd2cFnq/wOOjOTFEE3b
7xghbutWbVRvvMD3yyuLSIt30o9S2yt0vXBtcrcq2/0sNipA02zOEF7LbJsp7ES3
fce36lyaCDqgUv6W3HMt0YMDa3LddK5AdA2VmrDYDpnflUvO6PzYODHrX0W4WBZq
HvaGf4tCbK47W9Ds23C9TSX5RuQfC5yj/mbasuRlTmkbtZh86j+IG+ueGVOsm3Mv
lfK+IOkhTKOps8FBT1S/0VwQ/sKCn4RiLvqJZlrrYVO3FkUsloA4NPqws2Izd55z
EOYGPU4F4m1+vyuboja4GV6NnPRa123hXwsumXiIEmvhkFbJP+1iYWunIa2NPWwH
BEBA0ihxuznPY6uRZjH8fYDqA8gVNO6O3xAiLBzluFXWQ2Z26OySqPY/6AKJvppR
5jXBWh3jqQ/38xUVXp63EoC4gmO0x+47rAQhM9VONMxZ6wMC2YpkIIl7YQ4FdgLz
lYl0dPsTxO7jydINIUagpwEtYxjAKbc+3R62uxkS+F7nbN8KB60XADlTxRYGyVg/
vyY+eiWHZC9eCHpxVk3PZUdOlzvMwL2WF8NrOqVcbiI8SEw2CU4YEAY8nuTQ6ngO
8l+L7wOQXLn/a7XAQoOfdEznYtDTGCRWipjEcL6GKi6h3zYTDDAYH8T4j5q3uxQK
+OX2iCFTW8jjP6OhWtpHrKPegsV55AQ1nwqaQlSAza5BHWf5dPdosK7DB4KFZdHW
pUbXmB2Ko3tLCpZ9PJELbO/IqBhqGkOXPm+XO04KTX5F6BNrco8MhO3jFyYgVjcq
M/vfP9WbK60BlSnzbsNQler1gOVO0ldK/it+M6aiN64scLTXoMyfYL1lQvNhFe8B
lHLY5sxqiDGnAUiH1WiuqtCTdDvBydRmbJBWknAXXn61iHLgyENoQb3DY1VPaul1
oJOZnHpx5l09Rms41oXg7WrnX8pqkH74Arrsjrow71o2kVFdv7jicApLaoN0R/6e
O0cLTYnq9LGONpKixuESPeBW8MtSUB+M/u5hj3O6hnSVpKIMaPCOLLGWs++nzPj/
5q1g1Uz0tqXl2hDu/83T0aZUjIrtO9Ea2TTwYg8Iuca7asgb7LJhidVP8UYBVwvy
qls9EAGcabcoZAJTYsLmxVgqyQqJIp+ZobT1NsbxKGsyodBGUFFQVQhv0F+PxpSi
kUAcfGCguuUVq4KNi5kGksiAapeRr+QxlS4l91Ztob1WBjykje34MGKYsVkT+g+h
FFSEsf8Etl3KKLqNOTNuE/4KBCq4lqo0mA38r9JYZmYGKrba9FdKIrOjJ8X4xzP7
hyxzqotNml549T4dCDHpUNSKWapMlCSIBRe4AI5bq0wXa1WlqzNik07TV7I4BJEl
LiQG+9SR/huZa5PEzMhM5PYbMaA8jx6pJnCTcD9h1EX8YhwkLL+yQFmclZBZtI/c
zRzp8Ig2bfBDHyMTfi2fD53DV7Fdx5TNaE6ZNCIWzHZVxDmAG9EukO98DrFlxBoh
orA9IDYIGt6v5jTbUwuRw4nss1PEvfYli9u3MM8j/n9/lLIlXjQFD4kr3cttey7S
dy55FO8j/+40iODdrumxz7J/kUvOsIt5CuhCmYNdplV9jdVsPQ6Ya1jmayAHzOES
UxqV50ohLHgvoHSSRa7WSqM6xOYD/OAdiPAqocUNyTec/LQ8VNFDi1JW3b9X+z28
6FWJN4prEQqhDXhrD+s0pfvY6lK8sktDJm+5uNjHqUgl9N7NwYcanFz9IiNp4+q7
5h0NwIBrFwYn+eAZ8tM+w8dpXObx+E2CpX39PfvXrfmiAuMUvPftwDpoCfLc5vD3
H/4uXZ2CPh6fNxdxHeF21z8g5lQTyiSvdtauUaNWkGMFqrVIbe1DS41x3nxgCylW
pv6SSPSm0vn02m2zJooHQeqU0MaJDtsIYUtmxE5WmIx/jaLItRHkRyq6W4QFQmf3
wlEVqaKZ/cwjTtJVj2PnoPlud1qy4/E7N++mi4KnOw6TQmUn3x/C+aN/so2oCngk
U04C4WXHB4FrF1I3qcD2E0tX47klH4z8s/lwC7GiIjVn8gFR6J6+/iY8Gcf/9ehj
Zfac+BMBa8WDL+uV6bOCzgJlC5BCVx5gognC5f0RjmIvz9gcjjGNqe9gxTkFl2K3
SayNsk7zRelSe317iCdY4E58q6v/67lTyHp13US+WccsqPkp48f41dUppxTytzdt
dJ1YtRejoCNxVDwQnXH3RvziRkHsL8h4J5rf+bNFivktA5L0ynzjBrbOyrcuXUQJ
wSsPqKQJ+VELW/tU3FfVCO7YZ4g+N28/uBQa+18Ep6ikI+av6Fz01iuPw3fZA6E8
q9nfXjt/VPlx8eLCNIqjVF684RKZSNDpLTsGiqKERmNTPXHxZNflwFki92FW2fmp
jH6m8QtL9a1DEFkBolxpVLnuMaHatfe9VHx0O73UY+GrJkg+ay7fgNzTH/j0X6Jw
TSXxgaHHBodwV8JTxWNGVUricggx0g+EGJhETx6SRu8ALuFXcy1zQATBXOh/yYIJ
UucMuRvwlWoVVUau9vS9k1x50cE394MrNASPbt5U1HcRX6GP9tBWBYbPddAdoisD
TDeKehhAM9OzRp9G6xNKVsYjRqwlYpgSBB8DJYh0FKmIOKciNHe3bruKjQeY5GZR
pjbS+Ze4MMafgDdrnn+t0YdbuKOLdetdNJqQc/UKC1bW7RO2wiH440/2BiVQdiqH
6Mwru88mJM53QrrffqEB0JTJP52vbKbYmBIDMHycOtR9S/nPpKndjYHzDiCZQDvs
aHNx++0gU+4mh5gXAdknJ7IbcnASKYAg0N6ugFkMF0hbOxonG+WKwV4i1W4Pl4sT
AbVQ477I/D7lRk+Fov+sIvyzTaKD/sGX7LwOdUBn/qLE9To2LUeqKXjFJBL9LaSa
Eqbw+zkGqcYIvCp6UVxjbiiQUtb6m3o/fghMFoAM1DJQYJn1MWpk2jL4sY5A0L+y
HGQjdYG+m1wumT0npldVADT53GGI2ns0VSk7/H+C0yJ7m8ANT210hcOMH1pxn2nr
PrVFI+GD/e5oFrlgA9Z0ChpHs3rrK5wiOaCrFLFZU7xSX5O8zFVQ/q/r6Zfbong+
UGQMnd5d3alilD/ya3hYdgZ5P8g3KokxR36Ir7ISziCmA4j5m1uvRqSbvLWUFkP+
ImK7ulliUH19KBVVtFI4LrbC8FbKCnQwUGI/jNDfoDlxk2G7XDPj/qq+0qoKyvOl
s0dL8d1BvkjuKwuH26SoPQxR7lGdUHXm2K7Ts5ktC4RSWbBROTKDUZtES/3bdOoA
3FdKlqBKsQqVyY6HIOkraNGVK/Dm7wPzK2RpYCnlJP5I0Pww/WiEQLoS4CrvJV5r
1V+3xQw/qbqGSucdUEBZHUDDQgOi/o8Wg5ORVrwg53ArJJyacJNMsqxdjjb6fbbq
5WBkv59bOkvV5k6E94FvQLqEzJVzI7XdV7P8HFhJZAbHUYLaNNze/3IBKxfW02j/
vyQlcFnShLbMVt8FefOmfIyu4S+1QutR+cLcR0TJc05Iy7m9YDnVYCsCtY+oeNgV
JUigWfK61zQCa3BRNuwlKo2BM0G5mu5qcT1dhbNHMtN1Erbb7E2SiUuOawjq0BZj
Lorc7ljQ5uwGDHvzroWXUU/j/24hHPXXagWM6+ssyJ5r4/H+I9U8TWJLbO2nZUua
hVhPGRvOnEUIAtK2Em9pPUAyKiSn0jGsd5xFLjtetUCLrsfx3D1Xwncj5ppLYfeR
MDHoD/AneRKybiM80rK/svSxzAZZ+2oSdYk5u9sxLsNHrVUM5Uw1NE6tHGIPhnzV
K4YIXg1JlGOb78OcctrxWAd7mZSI+QNQ9BpiRbc0KXWjMpB6wmOwdse9+5GZ7QP2
mBaPkldOpnuC5QEXqIm6050DSJ7DkPBHZC5LTlxf9NQYH1RHgxCwC0VzUlH8PshA
4NF7ws9/fneb/aE1exxn1N8vGD0EvG8zyUQfhzWXOBS3KGvk4OUSOS5jS9+cSM+E
dqrJ6nLvQb2P3bvyukA1cLcObNEjYPVuEj2pw2UGBXHFpxy5Umjvr8uqABSVcqd6
tS/2qMNG5ZvJalZJsST1pAzvNP27NxUcs3p8WPES7F0v/4GQ9ZaZ92BRdFU1mAKf
BGMbZJwwVwpTFBwaDIGqwgqypd5XNcwIZQ6fSrCzArbGkcok0V1Oz44eK0IoM3gI
TB90YoWtjZBEQsJogm3jti1zUFXtL06bLkJILXBfoGu89SF2vrOg6vvfXYPjrIvs
h0ZlUkHgjJBpa+nYhr/adJo3oBaldhbqTMJk644S/Qct2MeYxifYFMPU5ACrbN78
jll3rqCIaPhepZISkWdK8+G3DcI4Ywt4ZyqCLR/UmW8tnzu6GkxR5NrIJJERr4Hl
9J9+4KWdhFoQJOAV8R1OGwgARbwq6eT/4ctf+jkhm5TYj9gY/P78Iteqfk6wfUpA
12slLSJVsoQ2e2Emx29N3qFQX9FCiIfcsTN38Omf28uZz07SLHfCzqLfxjpQPYlC
9jP4G5k0hDmoAwrfVfVqImdN/wFobOmKbTr2slssr0uyda+QUelYoX80xlnMpGlP
WvBOzFy1t2ewV/ylSbECRYv3yymYk2k/nXM7nrnOu70XbdQafPQDASuRKnwt43Fi
YvhvEeU2aviadiIDq2rofYzjlB/gCaPOVkr8nLqacsZebyFYtGT0OGYzwVSXCh6s
plU1/3uZKoEHZLXy+WdQrsl5Q1v/ZXz6KDyTk1g0L1+LKsBXbddALBINeMgArMr1
5NbdzvTdpMZabiVHQw6WZRNw3GF5iqwYLZGW3bB2NEfj3UDkkDK780/5L9341pUx
5DjpxF/xxZomYUfvX59xaWYSFBjYrr4LZ4SiWgtTH5dVkr7O/N47xfNg/d7dBuqR
iipEfPLZvcnEAUFUPZAmOggiSE/VU5EF6Mkg0GuTyqywzJfB0v4cvwgUXI5BTByL
Od7jORHtywaEvPbRHqBdcVxdNcph+TrffQRTGbm9iCxBKfI3BMeakSzUqocME2/S
SytFUR8fK6C7eIerHxo14bFHO9Pv/MkDOYnTAiUIOCqbyaGKUszB9lvcvubX5piA
er4AM4L5ebKAHMvs20nnHOfIyC04E456nWK9HEe76XiMR/8jT7u9FtWkhPgGS1ww
isGHtkE9E9IBp8XkgMO9vzn7xWo8+ZYEJl5L4vNzdwkJARDlXkUNLYKcTR4lNG8X
/nKVYW0JPM/fQoXg51zavuPL5ZVpHfgBFt1+aGJRhzAS9AEItJdf7re6ha3kU5o4
nii5m/CqbigHScD15bWbvPqP2lBXPtNPfMl+7V8FmbsE+NbUn4wCanPxFM4IKtTf
TWF+N/dRkVc8TAzZSsEavYFJ50Y20ZxYlFd2HC5h+LFXeUFxzl+V+B3cUp9CwOQp
F8aeq8pj3l+3RNG83l+8qkbONscrHrpAVH4RI6muSabsk85ggBgJ2wBLxIroL5Sx
h25lT640YjxWsHTc7YcZZxAJbr6uEOWHQ9cfFTFlSXLHfGsrW1nruZVoEHIyAOqB
N2eycBCTui628f4FOb6CFoi6gpZt2dRP0gUN0au23cOm0pRBJYOqHKwBYes7BNep
+n8NbGMc/BOx83zMC9NUxwOFBTd0TqQo5wD8w+mH22cA3UzDflFjgRx5JbDrw/aG
qUmN4b1cECUuucliZguR3lROKCyO1fcQL85yLm3C1q9PjIvjBFpEWXa3KWj76Rn6
fgjcNUmMKjMxpaeA+eSNhDGJ+GGawQc1RKSJaMx6GIncqW/+I5siOhOQ2Mbk8zIK
5rmpc6DSbmZLfiJGQP/mdnTBXWD8F2BLqPjOXcTQvl/2aEjAFlzIxUlPWLt4fr5z
39ohybPs6xVi0sYEB4aSz1iR119kqtB/PI8yZx7KMC9/CZ2CpsjvhWPpw2/4sLci
s5adMEbg/DWUct9/ewpP9XToe6pS3ifmNwkp62MSpGu7rhSrVaSJF6BW3Q4oohlh
MH+KfLDwrrAUR9Agch+IhoiIQWrMdOavpPiSRqybsDb8nvYJCizP0DZZI3dm537Z
a4IWpjVTO30bSVrWF8s4nymElX58+Td+BkSHOjfAg+cjbCX4iCwxnl2gNjV0y4iG
VbAAb7GSIsHzi9v843a35OvpFv6yKTI0bhUan8b9e4g=
`protect END_PROTECTED
