`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DjBU5Sekz6luvyI8fk0CTWSSAILQuEu2xACKPdRRv5vZSultUr3B7EP1o74W37BF
laXukws91FILZ5COYuLujHf11umS3ez2KptGbXIhz/oX2BEJJO+8Q7LdYZncIXla
YgLd6h+6x3TD+b8VfITysyzW+5HzdGjwsaEO+SdTvhnBYZNXOee7biPx0njuVuLY
1GKKQq30UZQf1hOI5PLB25xIHfdhymq7/OW8TULIc8u1D8KzHzOfj3K5NkV1jsgR
PqNWTTnnxa15IMA+aLMS9gjG3LfTdYsRhBNVwnt5KLV0OdDiIRG9H8u7QwafITbe
voANNIMiyOWx3KBg9dhRInslwN/g3TIrgPSMLB/YQ1SNliuMMHlVNjgVMEsUws7m
7jDPRbpGce8qTj+rmeONWmGpmY+NWf/ficFnhhNKnfiqimYO5eEjYwttKqkDeMaN
uEDWAfzWeTuNTbJvfv5SCvw3p8nSaNx1NTID54PGwHfoUqYTUyGCnlS3G1QMnxSJ
R8/qYobkoeC6TGzqctQ7frqi1PmXzmJ3Gfxmaks2o8jeVNz4IJKtNJQwsVf84643
ea4ttULPi/yszpGoFN4AdcGB2Zbo7Fg0Byrrygj2+fVcUbbFmmyhqZc2AYrXIFZ/
sD6Cv/vKA4HrLWHjJlFQW6fcoI70/jUn1YzSHRNBOVG/xbH8qjfZU4tflWktGTNG
P+/6TMU0OiAmz900eio6pCgNS+3piutkYW6ntHrnbifJO1lCzR6bNmyDAd1bNW6p
XSkt+TrjN6j9tWairp605KTqy03GEDJGWErCdi4knn4k0k0CuRJkzMtEFUxJCiwe
0vN3pMGJN3NU3CMEN/kBPS4ZZJ1jZ8Tj4P6vrQLmv5sE9ubZ+tMlQvmiI3w/6MNy
muMy9A8Cqs811cVPtyna2O8AL6gWVe9oEXrGSf8Fh4g1PJmlnMky3EPb2ArvLxDe
MJxwQZ257wpLgIMlWqlTuc+ppsyQvITVNR6mSuonG9os7rdRFzcDONdqO3CKrd04
XWPL9BacUqO5WY9xYckIfDCBBeI5RlFWr37oH3qoK624yG99mnthZWQKdnGL+sRa
vGQQa7oEKnIfP+TocBXONOBpUD+EZBULdCuwQ8SyY+s=
`protect END_PROTECTED
