`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vyPBwt0pvd9uiA/mZAkYhfZX+cfcsWxnH2PxInwWdnSAkt12gaiLmtl5Ed+Ev8RM
QGC6LAUWwysNyBDHOcnuFseu2WWpocTlv0VGZLCR6Tx+CY45jorUg8N+sr70GWhm
Sk0cNoz0Ry/dxyVy8zCkoDSbZBWwM0TaF235eOoDds1fK30qf0PHEs8qkxde/DdG
noeY8Rqpkm3qR4c5mNKfMIDzf8RmE/Tsyx0DWcBeil8mF4rP25+qXB5Os+zder1G
PC7kXPd2qn21fh727OxY2R61bBB6eGHLZd7H09veS64nIadBXsTmrn9+dak7y+iT
IKbsiURBMayXMUyyDU4oZZFIHu58H/FtTNFvgL+54yt6jgnhT7Y6d2airRu5mYld
vsKv7sOdd0ip5BTbmh2i4tGiMbYhuvvsm6pDjmFDz7OPAAPoYKXvcoK0CntvAvYu
`protect END_PROTECTED
