`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xdpRxhjCCa5KxKHEGr9icnCfxshZ9o+xlq7CLq1qwmnfa/23JQWwKSlk2Mf+VsbJ
oVbLQJ36FxMfzxJbEeXA/De1cGd3EQYxYOTUYngNdEN4hQQ9OtGNhyPeBQ1Qb9Ro
bI39nWbWC8KWJgVoFGqCee7W69TugrYUGvQS0FdSKOE7LoK/XJ4NeOCKpcWg/ctD
YxoMVywU3PFSo+Gli9h5gqlG4i9dy0TKVRlzlTx2nuCVO7y6TpXgEawHxWvQINFH
NVWpz/laKCQSaOLhLX3+zDky8HisE2ctXEWA0PH0/R4TY6A8CODIhYPxJvRRDWVa
ejjbAyNhtGb3WH1Obwthmg==
`protect END_PROTECTED
