`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uHUiP0QKgwQ5K/HnhsFymARU2NHNZasy6AtCESja1kVYhU2h0TId24JyCyN4NRjw
dcegZf0oPZUO71/+ceJKtiz91ISHnRvTMIEvmbhdExcaY6ron2WPc5ExUnyAXq2b
dJgwG+3kD4oaT0w2wxR9X1FUVSVCQBIECfUl7NAPsh8PrAs3PLoFqzm27EzbRwQQ
Jiw4N0z/vAjWMpr5egesDvCjSUjDsd3sbB20Igt+r2pYQq1Ic2E/AyhHJgLglQr6
zf1tW82jNfU2dvRmrqrnYYFZLPrXnMwXtxhiZg0Vp7TipJ4M5XkPCe8lvMom+DKs
z388GbZYAKFMUniKhw+wY+7QYuRPYJc80g0MsWKRkBXRf8/6af8CNRmQsSxnKY8d
l8j3mEaOWRFMjaNBjNwUcw==
`protect END_PROTECTED
