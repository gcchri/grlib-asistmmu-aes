`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Y/CEUWuXfGGmeYo/vLUIHMMiQIGlfIZJBlfUd0mXqZQ6M4BtnBCNpOSlyY5zMfi
BhbeAaFRZ/K6XpzxZq9migE0leTeJ3WYdGyh/E7ENSEQXbyvf0IspYp/Run1tMoS
v9KVcLFnURaSYAVl4VvMD8LIFIdbFxlcl5SeNOOBnuDG5yDqI12CoA7TS39/WpB3
FE1/kReqatgZLf3Oni84tZ5zV/5kTpsgT95keg0hrwr+qusUNxe9m9eYGyiSFv/L
mwg8dgig8rg6bs+c8W0CVJcn12fqueDvH+p3blhxmaA0uiYvnhYvZuakqprKb8EH
koax6kPohK2Qo/rp4cu/eBBAxxxeXpvL44GwJMFrO0gtyw/2NdJeAipxMx0896ge
0ptfmRP0Y/unhCCquNCjKBoGLXSBNNbvQRHB7r8SLxV5ziRF9a9dvSkqs2sb+ABm
hb8ZdTxuyj72imUjvV0FueZeiwjoUja5Tz9FOLyBe8CQOhzfZ5uUi0bBqOm5LuYh
h4pDJtcbRmjqHArXVb45sPnIqIDSFpguWv+kOCKpxspOy98HJ80dULNsBKv+f5RY
P8rfIfG42AnUIg5KCZok3KjA4qVb1nZmxZMr88zPMtUlJRIbVMayggk2sCXcE2cP
49+iLHgdElI5MjSSB4g8coS7ePMeZyYaIBLeCMl8C6KXvWvDU2U8Oxen0ZbTKz0B
oyE40IRFxpoU4A3cqBODVdmtANmnEe2PWCDYZeGpGnc7XFg5Byj4dPKmhAy0rP+X
V/8vGtKqiYWTkq9UocF2HxqJvqVtiQNFHzMfCgMELqbQBk9g0h2eVriUhbip9f31
DxpXV9dZIwM7y+92O12RW7N8pJqLtlwAat1xeJ7j8Ee1aYEWJAp35USp4P25cQV6
sKbNjXORVnjWmOvCDfs6BbqX39I5Vjh4baRXmV4ki9dQLk3INRcfyvyrlUgCAPox
+JYxjXN+7rWw7pfikpvQ6VefdoRpdCjxDQbJ2MVdTpDZ632WVxDAeT9M5TD9bFXs
i7up/DPQ7+OYcPa/0SeH4FAq+X0VHRU0U9tdz3cnvnHvECmFYvkWl3ibUYTkTc9M
EQg3oyEAivbnGVlhqhjtPPlnRQL1UXul2aHtT4Tvwj25FKWrRHdddG9RkUt9X0EL
9fxkv2h19kprdMG/+o576/wdelEl9Tu/Yr7KTQ7/x0D/6PYeB8RRyTgDLkz2YonX
i9oXJ2ziPGFw/TgyvOWxYizS7fNOXpv22qW6/V7DmG8rOq5U58yJah8v6gqVzQ8u
CnVLq9rV/8KQlf8O5P2GjZahpYTB/3NpIES+gMUucGkqXZLCEK1F0mD/J+G7Zmqo
m7KCh0rpTLYXGp8j4PTATqtHVksCenWdpKSDK3sR2Ni1FUVGfJvCqivRb7LWWKhZ
7CNGtcgVPzTCCy5AKKyaewzeYSFwGWOodlRnw6B2lGLIl/B2WvL13mTJ8BoqWmaz
Y8fNSEHb+SmzHFHeOe62GUcsRposrZFy7fXqcK49QQYx1YuYPtmhS1rI1TDre+q4
YX37TT9WxhiF1W2YyDWxPhaSqUZskWwusaV26nps14Jr8B6kweAh4F4eCEZz3DXk
biTz0/XpWSLaeLP5f2xsMsHEPmMf0UCT41cd2pkEhkRwdjPQHSlQceYvp8ad+Wc2
ItTEt80W2PbhfUqARy1lkdUkz5wWELY076yZQh67m7iT+xnTgs1omT/T5istvEKp
Q5rT+eLLgGtKBVNbfw40omCQdLvy9Ic8KdUAoMbvYv0ec5e2V9bYonJSFyxRI2II
CFAlcyw+qaOJU7yGrG88Ynt2z8lPLCGt4e9tkat6HmbssIgZtoiTxlcFIRMPJcAe
neM3GVUkPDKH28/xXBe30SGvZlHQds01ypZLJbrNCDfvorvAh24SZh+dYBAcpxQ7
WNG+OGIpKWAUUE/YPBCduHGMSPk9HaQkOUvz65yk8YzYy1H5Pj6deh2N4b37UQUL
xqfU7Fy1TRPGjjgiflhIBqt2yBkXbKqZnVY0qPmTwhq116sgnLuSw1eiJnF6jrin
pvfoO3sM9FHSdC3ysQT1Ycbz2VvRqPZ+lcsv5HR7aQqJJXg2IJgZbiImdPL3+D7H
nCAkmHpfjgKi2gRnJ4IFSasJf1I7MyDBj3uNQ0gzSeuLoi1AB2lwaWondIhxmBPd
GRfkFtSq+SONsKgsTNfSDFZTfRk/HA/mcoZLnmPy7Ijqv5I9Tp1oSS8HnzK7biAZ
NCrKtv1bOGpF0XydiovKSHEDNx6JsFDO90PYEWPI5VTgv8TtJQrzToH4ASxWWQF+
o/ITvhIRfG7btJfXIaNy0DEnIZRm5nnPVVz2hJ73Ay+w0qTW6JtRno5xDlXmxn8Y
vWEFBIUdirHLeQ3/Nm7TQX4C8FBoeLeGBCB3xXQyHVi+x4FR2XJbTkvj36KtPG8m
2vnlBf1KBpTt15wIbdwNx4pVc6AiNCdcw4FEep3UBGLFBKwgvrtHAlGLuu9EdWhB
QIVqy/C/c03ZE1MvYB3Br1rBu70VfQaXk2HdrMP/Uds1ANJIdoX2EpGOzklxVIY0
cByi7HeIZdLK6HGBCdcUwkip+XfEKJi7ROcZa90dxLv0mMjTbR7XhUPrwJGBdWDH
D0hKU8BK945es1qHPmPlZw/PwsEMrc1039t0C4F9ppGTqnRcEJ//uixyUs9lLijI
UaQSCzBAxKHEHXs503o+LLUNFPvdlOJP5Gaw9Hy5gbhNmtnekR4ppOjO13Eg/ZW9
MvGGf/E7XgJrT2MCvti0NLMCNVXLbfNkkuf8EZsL0xleNXBDEtSbGEajbmPCZ4v0
G8zoNgCVtc20oCJObPZfR4NbG3Keu7MssMmRqWWAvH6s7sSO7l565K2M4vzq8S7s
I4mxJM4VTt+KxdhpN7aPZIpu0X+ndohC+qEsYtdYWIIFW4Xio7iRGspYUQtJKaq3
zKEOvaQ9PWYjNcotAOwumsgBBMO0kGS8E2ozSoRoJVU+wP5srLNKuR+9L6/bDTO4
ixf1uR+fZa83K7F8MFLMvvKQFxtKWULDdD864Jyvvz7P3/rmM/Dbfnrwt9PQHskN
ileQAXBV2lt/q7Kvt1igd2AWAU9Q3UcIqIu8zVPmeNsni7VQTtcKHjSgqJgZMf+F
uw1e467fyF+Vy/MxYNVB+Ovb7LOHppLVDVOMFc+11kGnQLpNKYNLIyeEk1ZL0wZA
gV8aq2PC0h26lbm2LZXml9AoUfwqhnKA+umcww2Y/37SuSC+q/5miWXkyzXxcxuK
w0T+5ab97fwGLcyADlT3MqCBRVaPknbt+YcWNZrLFaxZkH+aLZt4zoO7BLCYvkbC
o970JnqdYx2CNb09sZtDKjMvuClKJ0FuL+CnRzy3X3MYaiS1w022gIqe0GlOQIBa
PfbHafBO5HEYiwejhtC5CqWtO1+JuaOIdWf3FLKSfzxrYVmCj42x92mg5tULicSP
UpFHBaxZm8Wn/l6ss6wki66UAqK22UTJJ83ZL/gqtJmrevjHdSq51+N+7gFdnJQQ
XwkCCNQ35zIxdjW48My9quuWamHtfDKSyWfhDbSmpM1JPbuJhOjC1KsMRS9fwsaK
bJHQAYUsP79dHw2wZtfth9Tn2EhuEi29ZUqYn9k0N46VDT3i8lmV2OVFsElPTDDl
kxM7PdGoAjHhD8CcQPN/DXTPp7i5EWxRJq5ThSC8SnjWodK5wExX0E0qG6gKjdo1
1YawDvxbJgTv+sVinEeYbQ4XI9/jNpI1YPmt+uI8QIx+rA47yGKOSC7432TLFwiK
YMzSbhUxxfl3jjS07Y3ZFuuErWFuy5K/GcUWIemz0bkK6XSOJ4QVbotD/Vw19Yy/
j+YVATOADroJxKBhmVEtvN6oZ53Qt4dEKPi56j7WoEMru/8xmIPTjNdh9CVA3Kej
JCy4IRV8WiwPebkQFN6XYNCyiWCmPkmFM+10LIprbnWFYIdoAE6/DGRmuBv9z2mr
2Y7IBHUFrNQVoOk5ncJUfxDUQiqU080wI2iNzmEvD/Hh923QgQI3S+SFPf+2qtYG
DHyeUX4NENom56B402mxa7KBr3YQ5KbffSw05gGRPKxsO/0K9YGBpAG2qkJbWEzH
d0tvNVevEc/WmMW+oHyB96pkuA2BWmh+MAczuHo4V8+6ywzzIK8i5M7j6MNrafLL
VWHjgZCYDxxqudKM5/A7UhHeYr6LT7jzLKIN08gvEn+AyICZeIROUBqK1A4XwUGx
7rYez76tqeAGleHFr9ybshFGdYLyaDUCvbCUAcMhmTcahLcug7SUZJyci4nyeiIn
kshk4fD6rcTQOXacGnU4cE6YAzOeLon3JEjjixjf30DiFW2L6mBOU74LylfXbV2o
iFWKP0g3CAlHPNP52yvHZ54kjEzSwIXYOpEZmrSu6flojE9xP0tWI07/BQXnMcbr
9KQ0FYeYOJsuj7wgnRAmriK5vnr/gs67Eo7drUVQwyGRk4Y7uQY6xex53fv5ID9I
nJ2y420QVufGuIjDLD3FhdR+5VP7ViUrpvRp5vrN3Cw7Q48l7WmrQJVWaYXJ7fTr
OJUPC69p6K+GgX2+gNezqcOZqAFNU53rzPguvaojnkCrAu21NbnbaqaKAM42ferw
aYKOdUlytkYbS5XEkMDNk03odkryeuXtmyKKj7Du5EM2J3ncl0i5CsIcmbS/5CZ7
XSr6KtacgzlmaPhzxNHjaH2vpetMzIGXtYnn4RBP38r3bhkLyjxAunljyhd7y58F
h58vPY0v4X5fFSesSN2bnaJ5B1fv3qmPbTdSXSUsjs1b5GzapG3yKgefuZv9+XcG
sLv15xn3QejJ9KasA9U21KooNb504us3p0jlfnyARHy9fQ0/ofFz/r4SOYpA3Vsq
su0mNCQWyJmkMpFhIcG4/Xp/PK7n25bsVivEY+vDqoLzaTtJowGZ8KNbjdtFdDqW
nPIH+EyXqHHzi61g+Id+KpjkIZk3gI0ND3UixEYUsCiFYRRJHQ+AFw80/4DJItV0
AbkWyt90oYjlPnjethpZlCBGblADlREAwHm8nELskOuca+q/gYadABVkIuvdKodl
zfnLvFCsHggIqi0Vy7eQurzICgzFStKON6t3oJiUrAHFjjrLnlk7XW3JnahZNW/X
86Ll1rUH+IUuIn6r2GhfdBr9+Mf3wXS1Llfa2WUY3VrCZy0Q1836IjaDBJs8Vk/Q
Nwz4jhA8Qy6aPLhEvxlLXSF+wlvAh4FfUgddMxSi1Z9MumHXxV3sp0n5sjwgATK2
hvy0I7luyE3BNDnYWAYIVRbSCK2uJtcC6jc8SJ3gKglS5jR36e+z8AhKPXhz/YcK
SngVA36HLJ+gkse/RqEB3j9Csw+iG5Ts/fOGpjBLSrXc5HNoHLPVD22LgeI0mAht
PBdMOGu/HbWnJlme/cwgHYb35HOckCRMqD4igHP0hcnFqGfFTxRZKZG2hgfMUABi
kOCrjWtIOcGFx0Sa3ldthxsqKPrCvjzqZpmKBtnk2VwmXJXC8iecmO4NRhNlCaa0
uWNsQf9alBid4ZqnJ2Hp7zUmU07dF/Di6o1j3UPWRECyRAkQSEerU1V+fw/WNX2M
S9to4GY6VclKWBZgsuCf96y9M1V/2Kh3FsQXfnZbPJzvNR6WB8aibPtyyld78brr
6jDCIH7Ic/jCFxVFKjDkNR/Uh7QHW81Yi3okHMp/3UAAniZfLfCBXldkdwZ9B73R
0/YbmKf20qMuyEp1878vKBDRKuvmoTWllkm0QZ4CN63PwP/sNco8fj3cS0ZKNAmq
yWTBbXDq3JUfqVrmdJ4ItMWE0DJ+gTIyfx/1ugGQSPXIOU31iY29IzCLWE8yWyEq
KkIwWPKkvsb0DlaD4ODL72p74DhIrTIkTSsNqXHVpcXzvsfTqtkxOa/II6PFNK9o
CanXkQa0PZyafO0dk3K3bPxktQGlN0SIw0/RPneiCT3FZVxiPCNmSqpi73N+XQrr
+mwU1u/BfzYDyeY2+IQC+eXnteHzOtB9bvtbGKkroHWwdjAJz4G6/bhNWrMR8e4z
VE6KWoMSXdfCT5glxpoXsBjYxP1+TSV/VQZQmWTmuRESqNEMm/YUUbRd+SIJ/+3A
cG8tE/idTDLfU4VbzgGVwZZSdXpenTizaHdvRObgKMib1onwG1VWA6emOUPFDRS5
A5sQcCgSFWJdOWMYHioKo/iZICSYqZwby5ey6kuS42OegKvtWnsRTabqqZFR2uQu
GMtcXuloKA3/i9PdmZmFz18DCvrEN3+oJxtQ83IPPmuoqgOr3Z127eqIHdYSI/NK
9elFX7kcOmFfkwzp0jxVoFGMClnGFSFJEuI4NrBGpuzxxJLiqmkcK6BIguH8or7s
ya8kma8OJ1LaJrHIafQybsVD9xLhJ/44J8KyK+uFH1/CXJmAL55P5cOP3kBSGyAT
UA1wIdAngRlBQWP9bxU5uyWhF0O7Wz1ppaFg2hikAaPkyrbgZptWCL7SwjY6ys8y
ffvohkdL5eY0z8w/pTvLW7JZRspSdFkr9WrM3ipPh/T9q6sFz33lIJd12dT3P7tK
dK/c1EkMJ6WzP3ME0RuTxAJ7kKtaK2teoIKE27nvGKRvQmGsPz+Hy1nJYwBquzft
P4xacbxvqPZk3jlVkhevH6H9ajRZ13ElcgD9DRQeiSxqHegjSPZW2XC/3/8sEoN2
DWNzqNYlA8bv8FjmmkmBikCDmcC491FB9TZPDenM2Cw5bhf7utmPurVYBNpRCyQq
KeZpqi2WUyHk8Jaal8indnOfc9sGJtfcK+0t8B08OesO0Mp2Zyc4yZu0uXVp6kL3
2pMCaxBIvczjvtFOWezR6V6YwMCEvApqkOVNJNgMCSmdsYb9BuJGAADP/OvBJBBe
kaVTLKpL47thrCH3EbIc3yha+byMioK+S6UuduBRg5jPkEhM9uK96yw5t3X21Ofy
vmQL3xu+CMNdQnKqW6RvI6Pxq4YsylTwsQPlEBUAABOC7UpqAgGdTemRrhRZhsWy
uF78eaZXJ1SzNUqAkmhkegwBTjVQdZ9w7tGaARNJbORRdyEUr58VPn7PqRPJsBCZ
WBgp1jEGIEy827smfU+WTQ67B/HO3nNjUaThC5ZIWxBsGn+nM1Q07xEH7MtWTpu7
yWRoOlxN51CF1xXHxQhWMNUbCCxcM/ugA4TzpSzmKboLkS9G88RGn2ZlC2rzXI1p
gI9hk37EoGdXJDtPW7Qljld0j/O5W8dU+f5dD03mVF6HQfmsZxuZyhxFxWRonjcf
VFRgOoThC6q77RFMDjGw3syXRtKVFHqPIkdeboPWSbBCxGmSK7aCe9WMGVj9M52F
`protect END_PROTECTED
