`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
38skf2eE6/nSUrjNVg8oXi6Acoco2bBI1h9PjOhf5rNNRsp9OgoS6C/zBW2pEwZR
dnbPhZIjiEtXWhO8k8AlBw59u4Ad3eAzQXoTOVkZCrbQL5TD9JKSSviRlAkzOHNQ
4HxGKqMcpC/nRfbMFPsOZo1L07BY3/ZcqPrOGHKq5+TcpWa/dEf8fKzLt8Ar+OE0
uwbgO+fGyMUCafbSKnfsVxh0gdnmswbkXN3xFPPH2uHKF1NQnr9bKzXK8bYD3WtB
79mXvRgKVTa9BQrEdeFUj67bbzPcdBasR/tx6cRcLxIr9jnNdwovI/bAJ1erxHee
GEnQgOSRX6u6vhCRkeOfULVyaBcR51C1FmKxC74mNEovv6K1Zg4+ehXG59nZruhC
X6fTzPrSUUV2frigkn1zBVFAAGc15UyHziZhv1gG/+ZRrwjqtH/HCQtVyS0eVMWD
cdTW22uCAq9yJvztVCv6/LWmpTCfMexJShMpNqGqukHO3HX0pDlzQ9kr/CRSxh48
ADrdCzm2AUMMYn68fpmVR1EeCRlqxfeNAMOstciTZfhM0DiQMX1YEk7XT078CxCH
fYlvm5lqmeVBva73pZ2csjW7j/04KZg+XwjwDVKgYf3ny0z7JCEwKHXnF4uwYoSp
bN4Rjtno2HO+T8jWeufqOly4SEkjSFJZoDqaRNQDYVz0C/W63s/zOGHeqjcXrF6z
R1wnkFheaPcU0lT00Zx74H3ydUOA8wEI6kYyNmW/XM/D7ZZFewzNczt3ma7sXD/4
`protect END_PROTECTED
