`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0vb5QVROCfJs84T5+BpAN/V19JzdL4RiDi0N4Jhmeow8SQjJW/r8VJPFoSMu/yI6
JkFSupaJmVG8GmSb0k7grHWRjvsQpflTY70hmK3MEXqYYunMSSQmi6r5ppabm4B+
tPjNINqAXnxQriU/p9cdMx/Vr1NdwtgcgLOs+opWUBIIf8ltPFMCkW1RoMkDY6yM
/PWGN87v5gLKSjaebf+mOybgjzqV+L1Y0iQAr8AINrhPbpkesZbHEnBip8NyNlXW
J922wURxa0gjl2kSt35vMw==
`protect END_PROTECTED
