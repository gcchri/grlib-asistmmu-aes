`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ni7KDuLCjdUdo1icLHt3gZyW9rGO/3/ptHh+WO93jnJo0ezTIMWOBmvJVw/DhTi0
u2fT9oGwf8q67Wj8bNH0rgyYo5POLqXLOWPFbXBJ0rJQP495w3hgl5j3NeKExcc9
6XMZ90frN/fh11pY4PiejjdaDaqx4EJFTAOqtCDasTQcV1AgLqK46bqgk55/L3lC
fHQO8xDtcV4QXsQ9rRhGxKsnNvQOWfaXTwGdhyF2PgwvKxTf+nUupUCBkAnrw7W/
59jshwVIj/170BS7VDXGFRHKw3RfvZCu2Jxv0EfLCRam1eBic6XyW960mp6iaEVT
6WW61n/3tPphwDpZkKFS6mD9iFUsgQlA4xJB0z6MDrCrNl6SYm9N71vb+fInRFg3
kRYET9aR/Ca5/uFC4+JMdWinN4MjtV+a0WiF0+QljYzqCTfiLt9DsIOtTAUsXzfQ
eSAKH792yN3aW9zztYn8ZGKj3AoEEXyq4+DGmC4LxxFqzvIXFVMCGxoFWU27o/p7
i+Xnr4sStqMqCOupYpfddI8N8c+P4eynhVDhg65wOdK7DMnd9gKKaLXq7yDvWQIC
obuM+d1xqpxA3/Ay9cXwKYOvFMMq/WxaS/otwiyOqZVBy1+4EQNFbmZXQWRnZHeF
sb8zE00rP9FOIFLKwm5yvAbqhfVvnj+mk+xDIZXBIn/JIY7HlJRVrhJbZve2iUzo
yOU3owC3deBKhKqQ9vgY0A==
`protect END_PROTECTED
