`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
doGWqsX+D4MhtBk2UwawBGgsnOKSpGVKQN+ianzfjDAJqjUN/74DWmCxK2VuoLZU
+rqXkdraHmnhgrx4KmEwhDA3z1QQVBgQWXYgO63yV50xiakUfOUGhkmWciguGcYy
xZftdBRfyfW+p8iJ46R5TqHFIrJVa1133krHrROi6aJElzdy96BfTnKEK9hN8Bek
NdvjtWHFUu+rrEJI72DyZG9li2Uf9qE5YlNqeaZqqE8MwcQhj+yreyMOaStI2H7I
HXyBdBJJUu362I96Ejb32gf28tI1AYU7alaqGyojcb33al5x8sguw7VXS3LyyqFp
uD/iGbOr3AXI7XtnVARqcGo8qEfncs5BIbF8DxvRJb6oBuCwVBd0dSXaSO15YE++
F2u5R7e3WdlQ3ZkkzJFYFAs+UvXiWYyVnb8vdfYc7yKKWoD1ex8nERg52iREdd5B
huAY+ZTTEzpEzSRZ8VXIlaTmCLUiMrHo5Jitif8C4Sg0II3+E9Z/QPffS8UCseWV
3OjZ/8g9Pu48Mat4KZSlGW5Wkd/FjmR4n2an4pbu67ZpPj1Fhifde+PapQcPGu2k
LyDuPKZrwdJMEjTUMhqh+sGmNzKnEpTgUKYvtjDJZAHm25s8wQDsOBGQ9xJLzsAa
mVk4GPu7ZfVtFzrDTXPjtMa0YbxpmTzlOCf5r6s/C4xyugFBLaXw6E8WF0MMJfC7
NsaSNEFTEw+oFpSvwlF755/+sC+7pfk40Q4cC4ZYEMiziTf2/XQeCoECmp2x4DaO
3ksV66fo+NaPVNAyYrCP7HJAesRXCZBYIagAcb69+KtXucg8NVkb5ouMnNE+EE2M
z6Wf32B3EiyJN3osrqtI6eeg1aT9fXHdk6qoGbcFo+tD1Tf5phLgy7iIowMhevHS
esZZg2oG07vQA9PQ1v3DmwN2PwppJPfUVDUm9PB5EMpFxs2vyFWH96YSL/2KjMUb
q4DnmbBaVKMb8BLbdI9r24yKa8EipqfKVL9HebSvcJQOhFlGnl7TK8GLD0sOh3F5
HxOIeMFsV9p/KKboUKgWZoRSylwKqZBTCogzvC3RRlcH2WKAuIVamQuidZCTUMLH
5UEsMXD1JII/ItLRatWKefm8niaZ7fgIk9ZFhsmAQjFeSMSujI6Fa9eyFzypQ+ho
B2SF0h/2bYAxFsIK8WTSZ0cDAlSbPNQU724y78oIoIFZ/aeEU2iLHogQqU7+P9kH
VDwqjdrfdecK+zBzyHv2G/TdfhP2Hen5zpFMKPe410s/RKLfkZ4/gc1g0GqLM1cg
IOkksB4zmapL8UeoIJKc/cEMQ7ubW6sUrTzEb+P99L2bmtLyKooIFMKJMFmkzWZC
QJoM0jzjvezsd7BFpqiv8OUM8g8PStZSXO028gU9MQigEVoUpSt0j7sjV6jzRHW+
4yvm+3nlW02qb5fAcX9hw5ALHiMaDg3eDXWQR6zn0F5UYECL9kbDK/gWmHVKPbas
Azel8/t6LvhsXTRcLqccLusJUrqG0cLNs7lk84vXWnH7uDvwp2NGYXMpKEgNyzIr
UggdN1ubISpgqF467Xc3PuDvkk2TUv6O1in2RhG0Wd7j2HrtGBrBGNvzb66a8pDU
MiYheJHAV0lMCpiCd2Qq0On3z3imkdTdojdB8x0aZ2hV5t9du5nEEiiVZXjefOe7
KCB8QKtvaydttyHh42bnYMPWaC2N8wR/H1v/W9A9IKLbwx04+vU146PlDgQvR3fT
cYKHvaVCmK5uogETI5m6cwaJ7fN7/VlRivECFK6netdUBGJW48wG/8hU7kaamVyX
SW2SxyWUn9yElnUnvlWRQEMXaK9pKaKAhLArpIjckrIh3Tb+ImhKPEMY2rle2UoG
z/DKKhIubjfMt/d7GinS2l5KXJoRPAEvamE90qeqlAVY9AixRc+o1hoynxIB06+y
S2153rTK9CEbAJ70n+D9XihsoXnd7Yg7wmDS78PQKb+2J/okjHu26o81uk2qp3ws
n+NTG6dTi+igTgGF4qHk99l3gM4/u04x6HG+itWQNQkcJ0BNdYW+IXyNm2u80cmI
eivoGG1oPEWuTGHyEQJmE75t2+2vUBn5eRJlCMfDMJAZsQ/m5o0MvDy+lZ8A5s/L
9AW0w+htCxgZlsWr/e8LzslwmxHtGuVl495qrf7FxAHBkevfd1JsVmM/YBMFATW7
aKisORDBTuteVorCspelZBNcHbASAeIZ3xirscesX2vkiNTRnURdganmqtqO4rxh
T9hS6ssMWE9Pd8BhtJFLeeHnjUVYIHmeQDiNIT1EBc9ey+aq3WIxyTFOepDBUJXY
eRhBtaOd1alI6aBlH0PkmBColG2VTo8YY+TyW+3I86yGi1SikXs9x32joraP+6G+
aymyAvSSTz7+aqOrWJTiZRimuEJIQ6C3oHkiHpu+DG70EnW0l3HwpNXi01V5WuD9
QBV5KjIOx60lu/uBepXMzRaszyETy8BSg/yY1rpgyhJCC1/lkbgg0UbqirZWu3kM
4ISxfuC8TqdOaLSHaLLTkXbYAxQrtioHTs3Nl1kFxrjZYXweF9Zr1/IIWKSwr08z
xe+/mam4Zn0SJW3NPjc+niCgwuPABhZ6/JQwvKC8CudMAri3TWqTCLs96lGldEYd
jleb+FzkUs+jCXCX6FUlcf0fIpgwSPL4l4ojziDmIKQY1BY3XGqj9ax3+sKehabS
mNlcBGUjvNfkMH7oGnm24KLWwZYPrA4FfWKirDpsIi2A3coZ88DZHuvFqQ2zaXZG
44Dn5jKlxjtIuU0H8pKtSQFt1Qdw5oxz6ZygImOU3YxzvBMueDpEz8LV0aUnhFF/
kSJlG72idT0p8whXPUqEK9J7np+vkj4LQKlu2KW42nni8vgGqL4zC9QlDvIzP60K
3f7Je3a+pjpEBv6B17dMhcLI8QtNyDCNofV1ct9Jsk8+J8i+pGayQP4yrD+X4j6g
QXYY+ZfD7H6y03HxRNDdSSr0Ubof1LM28iq3plTxskxemS08tpp22DwYI2Fui/xj
mbidYj/5l9XYxdD9mtyeFurIoVRjp3Q2kR+p2ALyb8P6EwZhSN3M614UNF47PsNh
ujtCu69/KfGl8XkzQw5SUoqbOl1dS9csEhPZnzF8aMj3J4aGPdkrPn8Up4Gm/Y54
uk5CptlOIbp0EZXAGqH28t5XCzuAYgls3Sbx2WPApyoSYgGS9u5LFzY3ciC7bL3k
4+yoAAXUkB4wYfMp5aiYE50Y7/qIZP45AVX9gAbnwuIrSHEQRowVw5tPRf+Rl5oG
hJBwbNJS5iF1CcQaJc2/x3MMLBMB6cGZPZHSgXMByLagIYvYHxoR/KtRSd3SViyG
1deArTWfba7gEYGfzeEVVlrNtB+J8dSN5v97/rwBaGXZAPWLGfYarjg7W6PUPYuY
PzqDCcBQUGgBhFizCYakgnO7zUxuILEh/sFT7Bh9ac//BBV4b+nzIehugJx/qdC8
Y8t70jCrWMPBhvesW283Vd35F4KFwIyQ4w+U+FAxvCLjE+vL3GcQJZb6S0gHfBmy
GyqQLszi1goJy4XZw4eQ8uELwZMGOM2A9VFU8iJIEe3QMCt77nzLZIYnoddduxhi
lHnVCMHPxthjjeSk6p/73Tirreg/ZgvHglvjH9K508oyaiuBmt8AY8kset2KtSv4
hQl+2X6RD0kjcSJVVd1uXk3uVezuPJXARcIrzmXU+lhOHn4Js5lI66HEjqzzjQ7R
jREldZVHV54nmempfWB3Vd6yzSBpuv4lLUymXeRt4pJQCo4pGt/x9zPwE8Xft7El
X6uw/NhDTJxVRNTFhw16Y1E3rDouJ13quqkGrUS31nT/+etSF1ntiFXmCtd7zSa0
BB94Uu+Dn9NjgyNOtBE7+fqBYg9dRES8RBmd011wzTpuoZq8z0I8I01082/tXtTf
JdkIbwOcEh3Na0OBQP41aDRxkGzUl1H9RmF2yYzGXNPDmxwJGwdU7eC2zz3IzX/y
ozAUhkMMkIrHWmLipIkp0Qc91pyRfX4WiBFX9vR01NzeF0KqmfNE6NgTDhumi7zp
MVHuo6QYpXogXrjB+ninVaCE759iZjb59ZMzSFAxNGvkDURWOfRnxg4VSC4oTe7W
gdpSFFfDDchTxTQnDK4qrJj4T5kUIRx4yq9ivHB1y/RlZ6OpRvRCxlhDv59krNx3
FpNJZymaz0eHk8vXrTZRPFA5oDzqYj7AhVr3xnpzG9l6FQ3wHIxQiAceTk14tsNg
lqXDm6tS2FT3CdVlDKpL1ac6yG6N+wOdubhz8qoHRl2aBoOpnUT47ZsKKscZQenv
Vss1qxfrVwX/W/qgru0QhhK+8rkFq+I6rnHILJvt0tmh0Ep9Yw1YVSPgA1C4myUl
QuQ9zJ1AoM5lfpH4BZR1+2Rivr+OFzMbcBxwLDg16rMlyfUPjbvYSlWvcyTu0y1b
Vrq/cC3POlacUHDHLckEm0lGRSNMNTQDvosQaCKcppGSLUeJVxu33Ld8L2uDguR+
EP57IKbPDre277UoW5Zi67YJwWiAphgvmv5LRlSNC4PoZnhdNXqITHmGuG/wKLo5
99Ok5YXlicS20rfUeDQ12+22vaOrNuu9nEfU7mou8vjKFvneCbXSKldbJn2ewr9D
r1P/scfXJXcgdC2YGd8vfy4EWVS354FDsGg+bBVvqYAAjJO4WgfBCy3T2rw1oYHc
xPpfCMpJHjSavwrxHMvte74rbk4NqnG0704CW/caWDVQZmmuuorMqtbCxrOP6vHj
LWb56PzpIFQXNZdnk0LsMzdtGsTAklokTcSrMmLd9wt/atLpt39jJ2CBzWjVteJh
T9opT40ODBlIh8JV79Xvhxx9gyUqrxxdxJ7V1pqmlZFLC9SonQlmVCeGwhqgYl+t
piokpOuhTThFES0ZszsQ+PPa6FmnWymVFbsBSwSO3sABXuuuVTQaBjfu+KknjuhH
WYQ+v5AbwWA6qW9ic2akL8tLt2UiO5xPclHwZ9j5W1vYQLEwtbT3WFM7r73pgjT/
CCSgWyOM02/uBf0TyG8+Td/CJOgWNSuMaTzfE59IV3vNMKIeNeAzwKM6ywxSv9Cc
mgNFMoaeEBmLTAxCrtIWla7n8yWLtIQgO2gDbPIUV7t278I1Z1sOq3d9G3qK0Mnt
I7BhzT7RC3wJEkQgJ6un1BvI2NtKkJ18ZVzk5IzYlRPJ1AeBwqEVHFQYerdjJs0Q
qlsaDiSZo9uOB+7SqOxHdstNV0aUOZb8du3iD141oZCI9jv3MVAbS31JaIt6tlPR
qGeJgIpB+B1Nz3g+saYPbLT8oRpjEKj7msS1+aGPzLeu3Gd0bNonSie8uM90jtey
JpH4n2PusVHsLM5en17oM6l7Sh5hvMqlevKbn1RpqBzjiMZWjxapxecMC7Ji8obG
YSjC4cpiUmJWsfx4nJqsP+j3/3CTmnTJT9piKw9eKWMd951oOZ2xuFd3Q8nC9rvI
hTT6tgLUvLZ0QzJ7xRqld7YU+r3/zgw7wJm1JkhdRN8o47kXDLf5jPBjBPWhf/td
ItUMDkkVy6vpAqWw44XPm/B8FvRuAdNlenyh/JRLgFnifc6ha6uduf8kvJa3nx27
lGvh3TPTGxCFKK+hd6WevBxRcVTcUXTSNzTbrYSYsfrtJRnyJFibR85H3+RtgHrh
vSdtUdgwIxvZeBG4pR16xJnlfHkkUUB6fJMvDEcJmE8gRnhh9V+3k/BLkJ+OMyGH
ypG1e36RhFYCfHJ2mUrmiHE534WDvzjI0kLOF8qHeT0a89ZEaQ2akWk/bS89YmPP
zjwsci6U9dFD68SklhKA25Q2Y/6xpBZZ/BSLg3afmckxfJlR6Iclwt5YiEf3aQCw
WuGe6OjrOwBu978X3IUJyrYqfhv5nE6lnsP4cvimrZMYJAO6sa43XnMtotm69R4y
ycMUujnCRIXQboP9mYdhNfFvQ++BQMsBnRPg0/DQ1C72DGD31Us6hjcYk/X9VF0e
Hjch5V8WuFnVpFZiebvHeYb+O+AYrC8jBnxptVzL9Nl2OhvfliDeltGglEDv7nHZ
JSSAKfFE0tbdCsUzw/eOYck09ZxyOrAD94LpKX3D1r6gG2/3XUiYJTkpaaqDVMVX
Ul/oyNYXR0nG61+vHWmCwEhxYQ5xer2LsIAX+8mh8NSyJ4LWjSyCWX8dARsqr6Gs
mrpBTPX+txZlxhRk3Who1hAUTN5oquYnzhjGRWN7fLZRk8qWDmvEKI3VZqW5BcIO
VFNhIQDC+Xx+jDbefmChTxVS/0U9+8xZ5k6NJ6HmOAuX8tnrd+cpH9Qov3I3ppq6
UAdRw6wtxdV/Mnm5CTTOfhOKQ6qJ4v+9GvKg80AZTEJK3coYNeeH2wMwXPoTZjmD
bZyn+tfdo0gkrv+IR04Bb6Ijyn3jkIT/2e/2Y3kGv1o9ShypIY/pQnfJ+FMe9f+r
iUPabFWKHMCeDLyrFGz/OHfoVcKj59+M4TUdJl82+vzx06Qmz4n1BFaMOEcSEh8i
znyKa/BXGvmvLUECsWFXE3g4dedb+4+Qo2LXLkUZ+BgVh1+SXKjjB2Xm30VRU2mW
2QRCeF5YRTdM+Dkickx18bv/zkeC5DWo5CnxgZAzCHikYkdhT0osk60Rshw1EIla
gQW7Q3+Zf5uJ2C5iy6L6k7RUNNC1HfAQ83az75nmq2SKOtNbBJkmvFo9MeS1W23T
RG4+h1KigCHZ/kQxwkNqHGSNwTO4WLGKwNU55coMFB6KdbL5IassS702arAeFHw0
yYBryjUY6Tc9RNfumJFqzar+0xLI6gaXK5vCs2/XkoVsazaJQK13jA8AkdLpZoSb
OU903vZy8SjMRNLaWjiKOKANDhL7QMWFauU8Rl9RcWdFtWYgDNin8QAnJ6IpHFOp
sc4mk7SBXySgonKJEZIzdEKIvH6wAliLotRbiP9faFyL5bG0S50PSIthvUvjb4vQ
5LdD+dN/TBvGYZscTtZQskT3kcgISn5T9VOoO6dSst8XEpqopus7vy5MHVpi4Sso
qCPzyH8nVwM+lgKpzfIGgzUaqk4pC9PyjaQ1IMglTc/hsUgc+8uUnGHobGgA7f2O
cK1BrwVVTUVGmuXnvIzJWmhuIyoyaTpwVnMkn3az9SkjREKF7/5ZPAq4YVYyqcc2
cOOgOkQfDCVYiPtLxWVfN4vOg3xc5T1nBBQf63NHbgh1ubEplT2Jw4FgA8HW4G0S
mqLkFnvZhQx/RTVixEDNDtuAzHDq11r4YdhWJZwtX4V9MBFxSwfcyg0sQl9Rgykx
08KUjhtROR6okqllFU74BGinCnnWTY5XpOWgh/HeD8Dp8utAQekvRvtN6A2XkH4N
GeagDdzM+RfR9axZ0MJxCJUTkYoNsCzuM/68szW6iuJng8FV+UOkaqiVIYuDiCgo
kkTJymhD6iohhZigkEsqDedBQoDP8MLpYewZBH3w3LIhzC8AL9sfGgfRjhyS4/oO
kBV2nDn00PWzJhlRquwGYmhMMTZ2WT2ECHGmRfUnWmWuF0NFIm+iF4S6hkS0IcFD
dOo2vtCEcFb6oYy6/O7Tx8MzIBxpN4VR4bkbQu6uG/OVENYvD5PT1k9tY07MFo1r
BoMrTEgR8Kn8iTvAqZO9Le/GNG/RjRMG4K2NDzAf2uWIhL0cWU3TRS+sFxIL8Gak
TH8BhAC7EnfYjudZylJwo9NejY/+ZHthqwdNwVQ77Oo7MDcdHNMguUo5nNzwV1iZ
u+4RWZ4S2ZafV7zbHuLzNbf01JFkvElySzl4ISip2Zsr4eBPW0kHL8Rsmz0y0twF
V6PbCeX6x7pArTLOG+/kqqmCqt/nMdokNf+ytssh8JiPqGM+Y7nJGijjgGiQaq8+
BNOAAHzPDuU7EvobJl6qjJoUw1CFXu02GEX8zy/zff+Sgtigj8lfKQG7ce/u8959
4hLiF4tYOwKKmqvzTj6fhFuB5VJuHf4dPzKN390VJDJoGFmAC2mz3PgoWGvqt85t
0OAM169Bk5wel1CN2iwMcjMje1KRs7QHCbJU4OulRHhQZ92Vm6f8oAcJg0PJ92tD
h/chCGYliXe2duYvuCVH4Ch9tiIH1ckNFwEVN+hlbPBG85rykxu4NWXqraypvEQK
uwwEyusXdxNnFkRsv/oUMQ5tJBndAcayuAJ2UC3iIvVBkmm18P9ssHCwvWDHsqnB
lCGmCNeBmmU7Pw6tRnAhxOaiWdCRbZUxrkWo/fwhmQiMD2e4gtCwtPKlBouNs0iY
subPzcvihlpjqcVqtd0YqlW1UhO2M+DOiwpohwrqL0GuY6n3biCKIkM5SZhQR0Dr
sDgXIOmqIHPf3ICqjDorVrS1ESOfvaQ0oof9dVyH8KinAro8g6JXpFuIqrgNCz5o
YojGmIv4w3+uvjvLZFEh6hWCPaXXun+4MdELrdnw3SRh44AkVr6htfJ63pibwWTH
LPlUrAARkaG0iZhVbJT2QiDbVUaqkYO5fYCBwBuC3KDsp7DIg3HeZhfO3XUxFHVl
m0XDJOFG4yXzKvy3EV6PNOTodajht9yFxbJTTPZyl1AlduVnu/hugqJysISVpZI0
CeJ7fG3/xcVhF1UZnjMoaPuIcUwv2ZzkxRt59T2GZcj97rZFLPVCgam/5R7CD2ed
lZZBm6ENN7kS4a9u1n8ipVYWJ6xTO9IfGBfRntPRU8Jsr5zp9C4Gpulfhd2Sncyf
sy8vvuRMxvDmo0+B3iogVXfEadBlEYWr7K9ber+WciWtZldIhuEa5U8TWpTKFJcV
kPK9domHJwvC2TfmTPbuT97t7CN0yzeg6QJRArZJ01AFB1L+lmhAtQnmpjUwBswH
31cakyVNwV6FPD79PtBZHA1Vd8/dIWbkX04ZjUSp7y0FzyZ0N+BoE1K3HLvsZk+T
4GnqVvs1D6lXjTi1ipNWC3m7pHIbd2V9ARNQ+wpuVHqVklDJomv8K5oyvUIGgs/9
ipyBA3rkBf/sTol14KTVJpMWULbDzcXKq40NLB+UsvvZLE2acxQn0uJ9a3Kg0Bub
9Ig0l4/4s3oBZbr07cJ4Ftohw59Qh8dtheF/6diVT7EBFuICXOsj1jUyLxayVDbi
KxHQ+050OBr2EhZwuPZJCosfnQwu18/FZOov6wxZpXcGybwIdSEceshtbaN4ymEU
Ki2dxc4LspqR2ppzIpDuCwwOrhkwGiRjmRFtYZItezmr4DJ7co9IEvEgyMtGTNf9
3By1wKtGtDgqNZGh6KI9sX9YRabY7g/TybVCcYLa0ldX9Wz8WF/QjiiMex1Tdd+j
9eur6ZF6Rcdc/WRzgiE/RBArUqyBv0LPbrdGKNkb2w6S3KObYj0fMGaY0PulYG8k
q9RT7acmDWmyIgoCw3UvEbFHzpCO3GXooevXLZWWyC2nj0U5rKc3IeV7rH7Oy0+3
JKdhiCuY7RGMJZkugkhdUuzopcyW916ZeAwhirsO0G2ACxLLZ/Fojo1OFSqI4+u7
jQUvQBX6yvYmKcpvGFWPIWZ4l9a1qkbQYv+v9ZklWDzx54DPmalEsZsMQNcrKynk
iczbxx2MWh5EoBFPEdBfo6pRZ+vvzx+uRJqyUUQ0EvLhUKzSaS5XFqJcnn5kojQ2
Ll1uLXr1DavQuWX4HYMOYnnYNIMcP0jZUbcwJ13wj7yzH+IhW9oUSEMqf2jqDUms
B7cvp4wECXrgyA92SppIAFJ8wBL3xivAiI1r1M/eXui20wHiBa55iqHpxndmwGVm
11Xr+necRhC+qxhVGZxoosDeR5ZVEDuawWuq6gHRcRFWC+o3Q1QX8M3pevNf3dd6
3NyNZOXdwHpOLhKgexbtmflfxYaOdXKlzq/R9EBprFCbgIrMLMnU4rUgEX83hQc5
+62s4/Z2POiYtpdPwxvmUf3q0/nPoJU+ROzXsPiCfSccE0/CC3Q1Tuj/8GnFaBJG
9P50SWaJmiL5xCIV7nffGyqqoIiCpZYV7/rK6t/JrKvqn/C1nDyQkDC/74l1UVen
1v9ShfD8sqnSpJRu7e3GKsCkLUYoD2PJerxzNzQuxqFF8xvl/+I2Cf7wBcHvAy7I
1S6BncijTlo/gRtT3+aE5Z/H8VVlHKhJ0vSLg0IlYYnQ1ticeAAidb8bwLR4p5iq
J9vH7/IKXuqayNNpF6UYKpdKryUR+ua7uuhqfu1PWlZKnNzfQvy+Jun7aUG7JkPC
NjBm7izlLpoS/JbsBm+dKMyg1ttB4rEc2jhRs/RHTNbGLXwt794ggQ8NzU4ANmnz
XXe47kAub+RQQCHyp8+tM4kXvoGGvEH8Q55IwNy/N3kBXkXySa+tBro7g51fdHee
0FZgVyHf/sProR2NSptJX2VAamLRq8vTzPX481XaF2QT6d419f2mRxJhJB6l4Ft3
fr/09MdUOMQ5Tag6MCB+RKItm1CVp3eOaPaIpa2q7nBaNEVm4rlk8/NrdN94asgy
NB1YLam3kLUhTBqelhT1ZIvvTdz1W9bRw1YuElX+aGJ88cCyiFEm+096FeA2nBHb
Bz+Ab2+9RqMTYoBaC0kyKaS2O7NsTJIFB7kibW/0FkOBAnK9w3UJZOBc0TTID3Xi
TQgmKXJd1XR5ADKoDuEbJeGTcs4BUjrLxg8FOEus8Mn0stCewK05APStLp6tJKoS
nb7pklcqNhgNAWQloqEnvg22ZuaaQyDb/voepOxU+HYLPh59CJ8nZ8ZaNrLsPE6G
GlJpzTUHegUXN5fkDpAns9W7fT+zxSXtQIEgCEhpxsxsiq+3vigC0TUyMdQjkakJ
Mtm+3SteIWmblaPhEOK8aqFc0F+6DCKi+MrInmPe4yqHlTfK2zu4EUONiZ97xrk1
wU0QlbRhINK8i7eY4CHX65YkGX1QR9HJYQJTWUI7C3GN70dDTsuEWz7MlzTtoEoG
beg7/tZEUqvtZDJ+pTqDJncThsWwUkWMHZTMOKmmFowV5gCqwDGBwNZLMVR+Hrtx
SqB3rCMsAEjwmC4n2PPuGbEYTzi6AeFBisMqfZeBra4k6RslRzNPwVvrf4vbGKMN
reaLjdOqzm/hPDnmGcAcuYgdcAmp7DHO3n4JHIv4pbdojmpD+22j7fmH8IJWzTQa
rTY6dK+wUhkeoMjsUQawDudNxpCkrc42ahnqRSssaPFqLEohMvQaoC+AAkIxdgM1
gO9wiQ2wIKkuWROWrCz5rXO4LfAmPx8Q5ICeA6lHshQ9FJEFh6g4C8itJAmdEG2u
kyO6NwZ9JsXHSiUug07WM+TM266twLDamYYrhkc6MYQ99AHkyEx9rvR3uq2zx/3W
Xn8EzSqVOptqVKGaQybXllf8gGENLfjJv6pCCqu+ESAsAyMLrEti7d+sOOifZDfS
o4EZ8lwziAtyjOR3Nd+wN7zdMlMlbauDRBKiZdmsMBM7LpP92qeifbrNfjZmW+jS
LL0sAMiDVcS41QQ7i/EYThC8LgKzaW0iCS1qtALH8Rnag4KrsDApuUuX+vsbcZwF
VP5FgT5OflUlx18AXQ4c7Y5U8M2MftZ/4PQM6ldPcW+ND7a86whglPwi2AfXrkRK
30NxXVxXgyMmNsRx4VVl/xmMEnsZIOmWWwVrHFqQFJjid5eAMFJhB+Q+oc/9iUAg
cS6AIHfHJB46FEnjKTyl6msfsvAEKFXlAzqlfvMUxovHiDcwh+eKu/muO9liGA95
2noMmvJWlHAuZUuZq9/eeKhdcXlnBNUxtg6cl978rfDltgn8rF78EjWWRqHrzv2O
5tIjcELArK9qSuuM/jXBwjbCqxhhRtrLVWdCEnmeRQMH+bGgBy29YB2J9YUNHIGR
hS2dW5U9C3lhZWcR134AZpmz4dKYd1iL0WAwg6tGeEzqEBDhnflN4g+P44at0J7s
hiL9sW21BsfchJSRISOYvyuDCD8kfr7GQcLzZ+8EwCJQPXxx7TFiDrtusaFDU4sI
3Jn07aO2iDL4aAN7E7Y11BtCRtsAtmT+6T0D3VnpbKRscz1tg6e0dZWBhXvi9ErR
CCBu8JWOzKipLZQsqgQ83w6CykC6wQ/lPXu02aUb99o1TcLheo8pOD9e14u6Ofol
h8pvVNRMsnp5Zo8BF4amO2EUW+9hYmUt7zdLcqAKMR/g09s3Xeg6XrPYHUUAfnw8
lIvNSczUxVIMnhnfLEU10wC8M/436RzJUTizztDGsBSFmr1c1a+JdkpuH82lY+8/
/8xYa4EwobM46H7Py2u/7O9vw/zEzSdSUT1hV/Py39ff7Mn5PFnz4gW4o7YfsCte
JtU2mrSvNOZ1wEULzEVRiOW2R5ALYontvA6cNHpZoBPJKVboRhgvmMoGBjivlf/9
XEo/nHOJd9jxpxEqB3/OWspizRvjniriUUpgB52OHT9XUPi9pqi5DxK6JWSpKQa/
pgx8OnSB4uSoZXGk3x2l7QjO9Qtm12N3a6EzL3JXqckqkWku/iaSNzkSlU9K5uIn
5ZpostQbTSqr2tFr78KrEWYliCYh8gicj6fqlmi7Jby+xoKgaSCjVv4rz+KaFS7v
eWpLbY7mfq/WHUF0Ez0lAWjgckavOYNXwDhcB4h91vyLFQZ7sATDH2FinF+7+UgI
rGmFuh7UpNHstHSfryArh2cMntqcUkRwA019lTN6h5jXmpUXg/2rzLEOhsE5uXq1
k2FU4wc44PINBfYSqE9OFa2Kp1mjnc48UqYjek2c0mg8yn48/j4HwDpuAHbXgU/V
YamB1LXP0DJpFfMPeOiiA3hzZGQ26awwdCVyqBq/D23ZA9+K4BwDRswNVA7YL10o
iBKtNTyKjKI0M6z//6GAwqeDlGfeivUPZ0xIMd+5eFAmkPKdKzLEIDixpzz98ujJ
SnsbuJfBSyMCUzntg43aP3hPN3nLjVCusf/bQjO2BkhI5Hro/fONRl3lW6hPf6T3
chEkFnh2JgT6SJQJeOiP2rgyO/mK+IjE1tRwUpp1KsIHTRXlshUpeMxIjKQvXSBz
2CkICCaswbk6PgrMiXoV7aRduYcCEhSw67MUiB7b5hzF/ZPradEdplbRd5XC+YCl
X9Nx25BBMsr9UgCAP+d+ikzzD0tfMMZ/nuWQQFfX9jn1cZN1XI2BflSWIWDoz6cY
RumfgUGq2Ak1Cvdp3thw+46xXOngp+cIib5O95RwerSa1t5IGuLogmRxp1p2Aet3
9Avx1F6HUPAk0/Cv1KRPqrVd1VUOFCOgeHJm3Tl7SsOZkTyLQklCQ4WXcpXoEXHX
Ptawnm3GFLRjCQ2/ZpZShJXaTFxpr9sT15lsoq2jS4uTQEEzoWfVCSNTllvRCQ01
PWBN06G0xnblFYmRjG38q6Iyf72C1Qn9iBLtXDybkt2GIfJFIKJuJe5xXgiPiJn7
nxX3eWxdx/0+/KZ/AJNsTOFReLvDl6U+eiuLJSg90qyojciifxqhdQYdyubW/PL8
pyGAnXy7Q2JZqgAQ5Vcple8+C0D7LMWAwt3MNUmr66uwkD/VnX+T+krbVNpXsKOy
4GxO+hvGZXbaC7MdrFf1gZNmRjbJu5t5h3Iio2CSv3358Di1QQMSDokAvVGrkP8z
B3M4diR0fNprGL/NH2vXQy/oxwuehAV6mTYgywAFYKH94fIJGkpeW5Gm9OVXypRM
aHtdtc1T9Mi78dtnxCuf4DAWZ2O2r6ZQldCfP1FRL8cG1ha1PjjDARuTUKFWYhhB
v25pD+N6Y0b4SOtwFIiZmzIH6C05/QXy+/MIEMkhygnQ904RCe4BIfzrYLinVLCw
OKv1/rQsauQHIvgwJ8xzJqHD9Hc3qWsXlD0xCKo++hD638pivS3E89HiMudJ9dPy
80LPSa58rSLckZ/3s9xHrhtQHu5Mv2wONx1V1TbGZ1XmXEN9JN+JxETs8l2D3H9V
9RGKaCczVKBW4KyQy7RKihK/6bSq5yJkQHoGTH9RTn+wXAxIOJSyZf6xlRV1ah13
nXmTemso/XedmbHfz5dDetaWv1QTm3pzcvUo/BMIPls=
`protect END_PROTECTED
