`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nefTbMG3o8I1r7reQFyWa82HS3M6zn4Y3LezLkeFfxnzUat7lQXj5JfHvdZC/ZlU
ByJPHA0ikgbx/BkhlTjsCTmLdpaL1Z7Ijy8mh3RrnCM/i82F++7XJMU7OS5lhwxP
I2V61MJmjZQvqIxVFmsvXyWNqgIijV00B+H9ZdgoVh/wFpoX1m00/HdUgdk++3vI
2Yv5U9J9xTSuM+K2l2W9FQ==
`protect END_PROTECTED
