`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SjvHEDM3lRSNxcqvKyNG90eWmUiLvnDXosq4nWuB0kkyAK+Ro5W69UsIotQgVxEw
/r8fHv6+TgEU8x40aZDTOYt81XW0vQHfNKsECiU+zhL0gCxuPgfNrpZ/LP0iKstv
Je7uD5NQglkXTdKxkr60QNY6kPEifHYN/mzJJfUVL/WCcFOfoy+zR2Tx9R3ulCET
SfRQ+bGgV9l0JtLrTxWHeQ==
`protect END_PROTECTED
