`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ZF+J+niOUTZv0Wblr42q/Z8+y31vVX8lu+zXlew+ezP9HVDADV+JSGMnkWj4N5S
AIARTYK9qCy4Hgy+MKnsiNNt7JfRdQnwoWW9Q31wjLP4yY3bdyl9cjGPQVbkFP6/
yvj6nAkm+zIFxlQb3TE5xAN1/Xgu1uaAxHenAhNTDgsUECsoRrppIL2AmgtJGm2K
Rb3OWYPaAv5qJiA3EpqrmKpbEyFEHo/5FN4HTbXbIKITSTp84e2JwOD1CBFW97/z
5n8GfSJbIUy3EtPhnS6ZPCoUv5HGvorulL6MQciftRWNwcqNwFAbZWMTSgx7nFS+
pz6l6d2+kIZesU9V+rnbnBwIYqgtpN55o3jkgJMf50SiywWVKoEYlxI+jZNpz81B
otgDygqci8K0t92LSY4rNLKZjGOI/cu6dddhwPK9IiJ+ou0EIBcdlpX/axjohxkk
`protect END_PROTECTED
