`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9QYTwe9Ty5MV1ZO/WItqt2FvHW/yNlUuUj+jQzXpEoxItFoSpCAgYcGSTPSmtcVa
gwOQMGYWMO5H27GKFbZfjx9j/01Svu+E6cSoTmzt3uCFh6EhQLH2mKheGBRjX3k/
Djh5P4kN/8OnIEX7/2fiklu5vql4t9yRgmisddRg2pCJZJ78dy+nJmDtUiRew/dz
BARxe9F913hAUKA8k4aI176LE1auWOrorHwJDuSECh3nnX8+SORA0qh4orZq4x/b
K4vfFDpuOBJgaZQzEayN2uEk5S596a70r6rW7gAs/W5awmFjUQYd52G0OTDEmmxN
fqhEuruwQShjepMMd/H3lCUJbd2rIJA+c1QAXqHqSvx28WtWJLFk2BBO3V6lSS3Z
Ds25duiJ5rGmkzaZ4XpD412tIFnce6uvqqvuGC9UrHa36IGAs988j7RuXHR97lpb
OdAJDXL49zlmYWvZEoNSeYL3B0azFglN6t6njqP6nn6vo3X6vXly48VIkszJq2cQ
NgFKBLU+z5yeVLaIFwiu7a5aHZEs4IiP5TpbeSeLhCT5g7V5uhN9xua30HD2rw1J
JiWbITi5wgpCAVWiXcmdEwpgOAGczo8Nc0ieeym0aFqvFy6AcmZOf5g5XwaRFuHV
S1TL9JV+pk1AHYrLGHnz6nyMRUDW4B0WjlzYmAaPNEWBH+cizO9ekVJppibx4Ij3
TNC+xGsnTfTqG4gm2VdZYG7s4mxSu4FZV2MQA2Zf5pF7Al53y3ebwNxKZ8bQcj8I
1kECZ7iS0Rmmk4ZGu+0+E2LtnEor+M1ff/nj0Ds+5x9HWTwV3xDb4vqrsPtCcfHv
1soC77esQztlSRgmCsiOTzXzu+EhxR7hS6RTE3ac2l4B/dCoRgHoQGdXhhUeyQj/
zQznDszHQrg1XBJIHjXdRVnhQqZj7531THvagUVFhTNEYU46MGpBpkqdxxntB2TF
VHobxdfLKJb8fKcmuJ6i9L9rxd5rZy9GfBK6P1iKyodYfpzoB8ssSPbOjnngKCow
MKkP3vzsvIkADEVZ+zQAjYPVn1pJhQ227H6cpqfp5RIgLbTWZ98PJY/co1Mv6gII
P05cJtd3jymrX4W+wXwOOHUZ4Zh460Deg2V1WcWnfvdUqBzOD3dqiQ82ndfBb0mg
qnjqLZVHDKd13BdXaT/yVuarZlE7pnGCYnTZ5XOXKTr/HfiVPP69vMcU7rT2xXlU
WrCIdoH4Qr1Pj/g97PqW8BkJVtYGQu4D6cxU68DaWz9ahrSVCMOo0ffvefb5/iu1
o6reXrQdIHn3AxAw59M34Gd1Rh75Q94JSRUwTH5xd9MtulXqleK3oehkA5RbtWn2
UU4LUBqqz/WhbTwSy+7cUflp+elrA1osGqKQM18VZfuw8YNAXwKHLPGy0nELznI3
7OjYV571skWl40B9pjFVWhFQjcU73RHa9j4lELuEqxrz3hUHTG4ytoYuQFQmXH3B
lrSJimpWyG0+agsyDtOaeldbdbk9HnrZbV8Vj01pX8bqV7KWU0FHCwVIZw7AtdUf
Av5yqyijpOgUdvsBLFam0wdtNI4SuPD966vva8QobEoc/5iF+S2KKu1gJ9BDJtrN
nu1nhQpb7eEz0C2p2vYmJ9LtD39x7uX3oPYvVAjgjNZQohHjmb0DtQFHkkFw8DHu
RctwTqYBdHknmsdSk/f09k0AKMRK4GekC2gnGEQiSZx0R6x16JaCUiIF6+mS1rfv
p2kDSF9vjaZYDmytT2uM2R1M7TY8jsW59nEBfeOQMhYM/ftdLyErneJQ1Zun5GY2
0Hd8OigvileyEN21oJ1jvJHQgBBm1cyvytMOdhcynnwROA9Kq7XaTcQbS3GXjc7N
0e3xW/4qIIK7iJV9bPXXq6Z+bifL3KVRsBHA7EHcp75xNaH4K7pldqxSk4e1kbk6
HgP1w6ktacOStHDNvqSTmJA59nfZD1/gUxN6uM0PGIQ+SFxN2/0G1z2vkunBcsPs
c0C2er06XSpZPw7O5MWDDPxZ3sthsF8ZkjdH3wIflkD9HP9sQJdDOcj/ZQQ6lpdc
+fn3tgRZ8h2wYc4F+T2s4j+BJtMas/fP1ImDmZ7WTLJqhvibuKb+UuOtPaENw+qJ
eWsFYeu/Svl2mlqp0ifhfhp6emykCkYOWzWscZDWHFHuuZWV5GnnsT3ryR9X4w9N
uJ13WUUTOPrl7r4I/bW2Dp93a1hvmgMJO//pgmWS/64wNbsXt3JU7Rdfi4HrpmvI
CPAvlXyMA9f+c7D/OWsW9DwHV4qVEG+JBuN3VhUOE13y0SEgP5zvLTgWyeG/DwJF
7mYzT1PkWn1prc0L8XFb9AkNtKr7sBZBh38iCa3WFZkTV1ZWb37LTFTYdZ0xejyu
Bx02HPNpzgEkuvr78dL/41oE23QNH17aXrTFiWk0ZglyRH88qXf2bYcXT/agW7gM
T1x7eDu2HXvhjQKl1LcADBgKdIf7XbG3SYp4QwLRLNUnvPU6p0CmmVGt2Rj8z697
+6wJPM+ycG4OApYD5iyp+Qgr4vtxlvt+Hln1lNEbzqFiNZp3JSTCj7U3z1CTKAOC
4jzIWCfrf4el+cF8ljfgnMMA0VOlWruHwG/faYiaJ6mjWOgESZ0ldggAIrYdjzpD
TYpz4gfBKukPy3qPjNUqP/j1yQB1HDmZFuHz4+lnW10NVSnQ+CSsGuQXfhssOOjG
wQrMu4LdTdJrqyK44k/yy4X1tW9gq6d2dd3trAXW/UBi2ysO76Q0IGpzBO7jB5Sb
vdbOjRvrVJaYIFq8imciTzc7cddEVgbisSvayVv7IquEVW2D/sQKVlvnuSr/9ata
rHSyPS9tReMuO51kE2/2DV8Sos7CF0lvZVCNu83by3+dUtBaXbM0Ay7Rn4r13BnG
xi6oiTRuvQGx0tMVwbJQlxD3EZhBHc0c8hAZM+xkW8bL9YEPBIlnT/L7TUcNY0PO
jy5HR1MMB/pJitI4ZpnUPvge0G8XT/YVoTDFI/iHE9M2FQFUo/uhaYvqesyCVRec
CFq2yYKVG9SxDGb4mXUN/oL9zSJEwD5slaxy5A/UDVz60emjdpjmPXPs/eDwSupq
3/nwmaoKdQ4dbLsHxtza5p78EPaiD9XaydHdZ3T9pFb0K6rT58GxGccMjMmHBHEx
Pvw9JbqAhLqNWLRjBcyJBZEyprmMOA340aY8Kox39gRDgVMToxGq3QxFxi8x2143
SEm181sw6qsrhHqyD+6rHSC9fuL4nidE5zEdWnjKyGuhTL5zBORZ0IhP4QfmXnVz
PZVLs8fsmUZjhSTnygJ3E4oPVNYCdJkLLHb26u2SfpxZgAESOap0gyZ4akpqlc7F
BF9aPTVNF8HwjRcGO0PO0wg/jHXiY1Nnq7S7tk4omFDDNNDEym1K8f/j92f9RYT8
8ZHdbGTUs0vUi+S9t/DQcy/7z+AVSXhT8YOZz/cyqJwRLHJ1G0+eAQbXsMxrkVXO
B3gnWlCkodxLQlzKJAdKkx6mlVjzD/FVO90XtSkaLSGVQLZwLK6qUKhgwShro81K
BGRgYZp3ltbK094mo9HS2iIfR7Abi7Ion6yiP3V6XkONw2E83zceoLV0ZmsGxjyH
IAqJ2xZj2K6L8PEwxp2hUg7WgIifKG9q94MlyInaL1ubRwLy6KGRUb6Fh6DruHtg
tBxXzOQVdT2lqWksDHhQSoXCOpGF0tVcOG3p59bA5LQ=
`protect END_PROTECTED
