`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mPXAY3VD0S/hmCtk0uAg5Szo1Ig9H2Qz8BJvsJEuI+YJ21n1G4mlVVp5/nm00Kfz
80w+AXwy+2clFbG771uaTuakTscamHzSTEQpUbE3S593GXllB6q6EKrTu6vO/jih
h+MAtupNvZttox2xlbMUzI1UQhGwjuhVr6DtD7SqUNBNcc7KNl7J2DZxMKMdfaz3
v/5idNSR57f1E7DSVGn53L2MNONLysOqm7daM+EGxB9Kzk6OBosa5IJ7M1nuJ/lJ
pnxoHwvn6ItMnn4UXfVKB6gj0F9Y0AXKj5u8mPVelTYQdlAby1tnreNzcrJBTaA2
yIwzlEzeo09GGkyE0DSRpg==
`protect END_PROTECTED
