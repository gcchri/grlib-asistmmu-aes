`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ww/lByKxXOtFKqczHrWqmFtS93d+Kr4hG4sbC0FKS1PxPlRMw4CpZkQzvo/rYl4G
mRxM2gl0bWGB37VGO6AYlv7xViRuVmGyQbG3b0TMosXWQUfEeah77jRCWYCJtCTU
/AwrD9ZZ8+PaH6IvGsiukowxA++rpMfC63FwuMN397pWuf6v47agRcxFbkAxGU32
DXVacArq5kL4IgyWj0QJdnqsA3YnhvrpC0V4mAJcWxpBeeuhy0QTb2Mpr4Q7SBbp
dJbgarlRi1RmDe/XocPNa7KVBBXxoHjHLGLgFfJxdtKyWdEjI0IZ8I18tcL0OFJU
DkZ6vJ1UaUY6Nn2pehBl6/vdblSi5kP8HYOqOGGmFUHN1GL/YOqFfr8d1Jj8HSEl
3WBfF6BuKOGBIUpLpJXqZFI9ycGvK4RZvLgFjORrTT9VPdqNAI12j2KahnCZibMn
OTec0bjVB+wJtyefazYJmQcBnNlpWwRYBtYU3pXCdTqD6fW9QCsHQFWvgbVpcDga
JQqxlowclaXkvgwWfCZP9dsF72bN87mQd4zXB2k0FMi41q+uN2GhU2HiculZAr4X
m7P5fx/+HA1ARKMz6leWh9RRwGf8vW15sD0p00K2JejZEDP6Jv8mqM56xs24C7vG
iqKXNhHMe5cIx5hDA7SjYch0+MZ3VSrBdYY3d7pWHVhAlm/pZyiiJL7b1QnuqOcF
BR/VEL25iGsYLJ4agbruwzRyhOv2PByWL4KAmeUVyzQ570rhCVqJBGWZlO/2NNsT
VVI7j7qCOBqWfoS9/kzabbxCfSH8kP7m2NfsvWqi1IkSgr2V9nmg2yuP9NIf+xe3
aBEOuWO/Y+EePDWhPnoR6b9F3QgyNZIzcp2VmZwx7L/QoRBcqP7KpNoiB+8CaP+k
FE3JyzBxvUiUUMlajw6F64Drboh3KO0QOIZ+MjuK4twQFieQPi/9SmF3iWzwOYG9
FzFJvvHnwyYTwKyVlP6sUedUs4LoizX/ohnV9p9tyLQKFOCt2otafNDAXsFpnHHz
tGm9OGDfg1oITUfJJ8bob/ISfxrnb0SNBSK7jVdmA9WQq5SRtmoHP/2xJEGrN5Hg
vaZqvXtjQgUE8BXZwl12Pj6RWrWjS6nFqkSuE2AmvCpEy/nETiD6qSTL2pgABgDU
3qhqDTdGBrGFyGMKR8CJs4LnuRKgIFuXmdrfybI1nWiHuqqtZGoiIPX3fUZAwQ9Y
l4PjnSj5Mv6fsFOed5/nZWG6hRPhNyBtDN65Rrr/Pbx2zhg3W11oRta4HSsPPFdP
ub5rb1o50XWl0DNJVVMHrMZMC5cv0fbT6VTYJHoxpK8jTfROAiNStj1EbHbBlDAu
W8RnBGFE0IwFSS6s6MWGRtjeB9jpR98hOEU9zFCRJqQs72fMAN+9FYjuuQnZ4MLq
5TBdWvhHiUbfSuGYwgql90tFlibfbW8BSdTJQurwv7Z8+SCjRQsyJ0qpt+4FxBn5
MgbDt50mJE0MstSeVRggHbYkmD6GgvVPmbtjP9QATqLXvI4E4B8R+V6uszTbBRII
zeO8oHYiaRfL6uimydeD6ksSfToVYio7USLF7541HWnMzsrAb3IurqatjP9673X5
8GFO6imPWd7zKdROVg6skMckKtVX4OKx1TDJR9jLkIckvRWjsBDC9GODpEHEK6yN
9lhu0GQWLTP9EwaUnodm+u78RkaENEX9WQWR+ULQ+l9kIML/KIvWa59ttNefW0rN
a8j51GjQT2H7uV+KYOzvCyNL4jcvZaDTdsvi1YQcAXpPKS9qojVUqWcLEe1Oorm2
pxb7pEMQtdK9okz9vZwHPYash8lHGzjRoutZLaLo16bYVGjlhA4RFe+J2Tt3CqcX
hujqgU+U6ukhrobyYEwXmHs0zxqlLx9ccfcBz56m2Fhe8/4LSPIbHBlRP++ZHmLh
`protect END_PROTECTED
