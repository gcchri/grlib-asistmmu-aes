`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NphjgvOyYkvWIlZng7e/28EJXfZt+ayMr70iUrZ5/ZQdfRuQlZ3sLEMXoPjiJHH/
Nk+0cEBARZKgRQRsJaRt3dMZJEo09KAUbSvRmXkdKNnPPtBd1Fyvg8K11fJleFTE
EwzrbIpef685AuRx1/JiLaqAwCYXFt0Ubwk+zqnPNjQUjbpIqchmpdtisRi6iEBj
LZKNzaG0wMiB1me1P/MUuf97HIWFRSnrNKux/Er9bvYjNagnSxTbv/NnSGUcecPI
WvHVJ+27raeonHlSHXlbiGm1evMx1c7mLf6glXwu7qZskn9axdKAxaKAG9vM4YyH
`protect END_PROTECTED
