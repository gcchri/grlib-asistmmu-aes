`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tyu+aFtB07bL4gY0yA3yjPWlEWQBNhbymchiRd8ySzvyq3hq95S9jyCe612VMAeI
j0kLRX4up0oVt641WL/6bUq4wIisoFxDB5o8VlM/e2PVtgedPQXIIIhfhTVd1EuV
W8NzLhmEo6MiTSvCa2wF563ppq2o1XPRwnIt2NbzpqdnpzbnjDmFbrET//4vfE6I
Ou80PlIKPNyFSlxTfICPHY5V90iozzZQ1p4bmmnrYGw0mywRzlz2UEj2doJEDRU2
1yD2qDBsw204oE80rdokvzAuhLqPy1nVUUEowsrjHPOPe4UGRO+i81JMdww7+Et+
zuHJ/VJ4g0s/u1VSEWeYj4VwJzK4W999kv3z5QjesK4JWtBxsPOuvl4lqjbedZTD
8wjAY5nWxPqsAYxJCMPSMExMYN2kcey8MKmWY/qNWkH2BbOup2f7f0dXzNh9gYYN
27Gq9MT1vWNqjkAAk3NVbxoHW5PpHqTkVUfTlJo+i8v0VBfrNcxwdVDd9xoLvMpE
`protect END_PROTECTED
