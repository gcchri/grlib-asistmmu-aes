`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1kgQegLOydVOl2fTrcGU2nc/c4dvSlzTGOoX9IZk7Zo5nwYRu0XpDrovEDFUOyzo
C2cdIMH8WYz/L500Bw5RcVLZ5pzSerwdrnZyMlI/YO3UtTcBFUdu+k+DhzcbzWzJ
Iab8KKy1KeVIQbCO3XlDbeQNGKjAK5ALsHbtG8+pcSfrxpZ8IoOeVlouGZDWBNCj
XiDGdmvlvuHQvFKI9Y0+hD4UZZXw/OmJOEt6syFJzWaQ8M8ad6v6Dtt47vX6x3b9
hDBgxfS6ZhIWf6PeHER6YPQo0YKoUnc+0D4/P7OPqfkGC7/6CbaepyTiogwv0B4t
gA5RmI3FiM/h3dpm4+ZzTKzp1Pik9GURNtq1XBlhd/Txe3A5dSAYofmX4fjNFTQ/
Djaz4671q1md0U8wp78j2I6bTeUAj3taLaEUQ51iVD84Ee2bec3C4QAf4oDiHRJX
20EokAzlyY3pL1+zZwiIAl6JXls8Rvw734yD+/mxDAeL5aCse5O/UuPuisrPkaOh
p0il9vwvDOW0ZVoCCArqp4QEVmUfUHqwUg28ozHbd0Tnd5/NeoDwIlTOlVOgmSxW
KOTA3uSZpRfHLyxSHVNzPQbkrulHvv4s/CHlJR5pSAwBcw0vckbD5mF5a3BhcVtP
sgAQiff/0dNaote9+hPC8qdAnKfMVE9fWk89Emtq0P7ulVhJx+pU0s5jsphHJjZT
uth4OgRj/LbeCtqnpdki9ypk7bgDNgg91x6tMkBnf9eyHZPHcbfAn5mDPNRjRLWF
h1O9CZGb9dXdehtycqgvjqwl05kzvvon41ln79p8gTTQNf1igVvEEMaCKoyXYayg
T40+KwPwnbaCdU45h5htpuOB9yuimWboTZZ/fOyMRhsxsKOkTpqvAxo8k4VEHCUA
GPXo+SiqaLFRCHuTCW1RsW38TcScD/2A/Cu0Tu9YlCLj/HHOZKgjALtp54+0NyhF
9kqtNjh+NLkEBcSEasozWeTiB18SsVN40v+NK81/FV9MnuvhKFHWOlSfNFYGxL0+
Xr8s5BfvSSgkJwaBftmzOJieWYTyUZrfMtMYIJIjjWqVz18rfdoMEQY3aJ97yp1D
hAKbsRZokhAnCUvBHbwyuj3hAzBTKa4Ktl3jb4A7fDKp9+JKfWtvCtNl81ULMwz1
YI9tkUCFMOCyur4VWhTO89Hqjo3ryMXCkrLhtTH4duEBaS2azhAyZxrvUxoW0oBG
ZdAMKY6oUYnem8eKFVdQbOUmSwZIWGx0S6hJeDq0eCzjgoiMNacRWKiqCbU4dOlb
S40fGHswn/U3Dtnfv+tL95Zwb4cVWzJp6nm2QgThgDmXCrWgaw9kOlCVK3HBqWt3
lhox7/Q3cB8KASsOEJktsK8ZBtl9YGGhxvDzyedlVz/B8ZoVH7WKEYNG+IVxrB0c
p8RsJ7jng3ie0YY5IYeeH+Wapo+m+b7YgIp8T7pBZP6yPhPaDHZ4QHnrw3HFwuyG
hMcSd2MjpdaJF3mq3E2pPxu77Al/kWWn+Uyy0CSI4lbIaIsxFOz7CTeeuaQV2VZU
zszij7HVbeqvywqDPLm2I1CuadJWnaFgeE9JE/DonrwyG6scJy0ADyDPboEvQBdj
Velbbg2vTh6LGEAgK5g+uTynVCUlQlw6hAc6xKUVdC6q1IHUXXuZGW+oBhX5iEek
0CtWwIdEOovurKOqGWoqFiyBLQTpreg0Z+pBux/36aKR6l5WybIttwDkhEwxiK+4
7Sqm5/GEaEf5dW1uJe56fCjHIfPxYTz3zf24sb4WFUSLxn1oyZeEHS0f7kdF4ojO
T3WvDSyl6O8v8EdqEe5wHI35EwdSxREueDyiH2Iy3ZMClw4ITYzT9xHeYqA0jcNP
YUSxd2GXAUVmKmdrANkCbdqUXfKbNKn+OIdC4GutCybrHstCDPRrLmQJ5Vnl/rXh
3tj3nGfS99wnv90/yTiWe/qai84sN1h8LhgpNqMJRRX8xVRj//0Bb1JTwWhuMl9E
n+49nGKJpdB6VWWS+Kf0O/wCqZFmsGp5L+kr3NkAeaQfdjvXkbMEt7z1c0CVUOc9
jf5LS46/oIyvKnifMXpUyuSPrKyXfQokPMyg1DxxIRdAVOBlyh+MY1eChOmC4JLi
vmHpOf3LTekWAcmyV9anUuQiIi8zvKyJd8bmj41enNK9/lU3yRSHRY/NktO5w2fb
domsn5s99n1HAjAJP2yq+jhiTrnOpBGW7dKrUOf/R3La3W/5mGnz+51SO2injBbz
+LsxNggJDlusu/dPIKVa+bp+VQ+ByvnWNEu0mVIhWQ/VO6ZFSnufFa+OMrpAwvWu
7w3IZwQnqaLddxEuC6hbtH6CaP3Z3bZkX0SQU85H6nHI3les/D0RAIw3kej7y69W
2NUFU9k8VkpXYUO2KM1lLdNW9j+lmfl4sQWtSwTxTaahReOLuxH+nmTrnOBgnYad
X2zNfSa5NTWtCuNWMDFslc8kU+6dEAw0ZisQqq+V1+ArcQREUpebjInflo3biAgO
pAuxWLVJwBjcrRH4HTqqralnE/7BLGe/HMv436+ekSHrVN4o1Thp4vlRGGYxPIxF
xZCJ4ekygtuoq3KB9JrKBm9qiCL39d4+A8if3JhzngkBomo0kHiUhlZKAC7EYO+c
WkeMMnincPX7wsUmK2s/N4S5bIRQdvxzN1+tv7Kj51U1nXEc7WsMFvgQQ9o2A20p
ZIyN4GqYMrvOTPYbsXzg8GVZAuzrf85io9MvpaC/pb4XyUMl1ByVp05LXq2Srq5r
tRVxglvgL3PYuPzdrDMLAEIZ2qsagVQtah52qFm1QDo61mmOzEUbLf/OLkHos4m8
bwPGuPzQjyEpYIxudBsLmSu5KqH9gXbTOt3m6h7u/bZbnpcQDoBJH1rf5cz9tMFm
b80Aa4jwQFpxW3ZWamilQiaconkuPSf1nxvT+TwncPQFc6LrLsEDF7gbOaD+ov6s
WKBQqaD8co7EMAihFOWZboHrwARkNTRzKDgmxjL16eWqUrUxlVfry7LgUWjPK/wv
BefhvXX8Jh22HTyndVUc/xeDaL9+jA3+43xKhsfVmoEERHYt1VjS/kpDMTlktJBa
rh57MX0iUH1SwZquWzVbk3RqQ70BYO+MuZ9Su1sW9oB7wYVjEQVuO6iKFKFVxHeN
LiYiuYlS7zYc3aQJrHias3tu0IH9ixR3bFMWKEvxuxI3R1MFobD6g05GXelyxmtj
Fdfqf3MDcQpBPff0q6jqpv31jbMrnWQ0VV9/yYtXoM69N0pURHRoGpgv3FhnGFZj
zd+RIruoWugnpI0rjh9+QNbfddPiYbptBdlzcDBNHxyVU8zckLr7r/hJT7LzgTJ1
rKt98yRFCB2qPRHn/aMXVJHu4iNU2QRW1aAp3LyFqkAFCYYxnhgJQ7fZ7eGtRQ6C
myDNAXoVz3eiFqt4EQiZ9YKSqFPOjk8KVi/d0SqJUBTYmOY3a+GcOMx5x2a26deu
tqlIUXra36XZArevlDvTBx/C9ODfTKzUcQ9yTyQMIyETdgZUSKXa37BuMOnxJuKb
hx0YtqVRV2lPjWayDXlevCl3G4oEDwoMJSfgHjrX15PmdI3MxhlgajtxRBC6r4c7
cbI1G84eTqQV5Iy8fSzHCk1lRqqoFD/m+Ac1tRLZfAXfY1Z3U2M1yUPxeWkUs964
DITpH69Lk8fdIG62FSlCmh0dqMK83cG9YAvF+Jw+D5TI6sj9dvm2D4oAVihzZ5Ut
ziy++MadxXgOVEY6PNwIt6Il5WDw0GvMn8S8BXz8o0x4LnH25h1BDMJoKVLmRSB8
Ese0xpbElGZBaOxM+EUlBRSQpTBvFOMqIikC+CdOU1RGVp6StUPmVogcJIen53Gv
vylKgZAdfizkVxEcbwi90cy2KLl9Qcl+9/Cfxf/5JoibIz4WsSiGKGG6XjXxJz4S
XH3XMr1yNlAUZB8RPfw78RI34PKmwR+dBXHTCoU8ixHbF5z5Z8+1scjRnMHlVH0a
4IMy/IrGaVa7ZlS4eJDI8XNnSTncoe+MxkTXfq5s4vkHgkqQ4krWljKHs+z97Djy
zVx735MIqHev7wLThlY7plPHhobZyUw/GN1QCRI0VUb6I1Ax6SDWQFX7i81gbAWK
CVfbkDXEqvdBa+5+59qK/Jbar6I2twu2HCm1rnMNvAIZk1UAb34xA39HDdXb8pKn
KK1wtaoWfNbyEKWA6cPT53p2Ji0RtL2uWQ3IYzd3an7fSJNhNQOuxzkVZhkBpaQr
sqkhQxcDzFv5n7zT6BbZQPzfoRy3FpFIS4zbR/fIFLccRwUvfTr9QuWPUmQd2J2P
SWKcszDoWssn90OoByjqL/+461oQfpQGOnt6zjGTvmpuXki+maGwdrW5s1aGx/Rb
C2Ddla+ZH6Vpby+oQpmzpQKIuh5KnsXLOn98EADTwY/j5XMeXT7m2dMDu6E7cs1D
lfuVnZGR5yNPscLoPky2HfTgLm81K05Bf85DhyXwoji/jvkyGaeEaHiR8q++5ZUI
ug1REvib7f4syBEKOQaFdgOgcm7c50iGqTYqiGFyapEsZjHASgMZCaLUTCiYdfA9
MnVRqcJxvnsTwMOxjrH70/k0al69XmXzdI0smXhuz1hF8kNqcoEOe5Rft6w8eJbr
lKpZxEgQCpA+sRA/BAc+nnA33Bw6EmLld7FKb0NWQZwLDfoJ4E/o84sIdXa83mfw
hoCpPSUWlHAjZNMds7PVCObRBuMIMgBJQvNwJGmUq7vOaBzYqn99wwrwRPXidIom
EBe7llgjTOCLz8xzvbNU6c9o6b6fNPAZ3dy72uCFvLBfWSEF69yXWaepSkTNgBC0
69DmXDq7GrFzYYobG1ynADP12Of1/ymWXq7JEO0T/wDV0U95UeD8F53vZ3d2U2BA
XV9IRYYFa0Ow7cwozMQdhxmCsj/putAB1j7q9S8Xon1XU+wH4Cke1nnHha4MKVj1
+iGiczsjzQGH6Dvu7x5CVel4UP8kwDALKiT9butjFozXWvQUBA+1eoAisWghaCOd
UjAbuniOzhQWSXV0x+UzJD9t4eLYDRxbT3+Jh11tK9QiRcbl4UYT8vcrPG9Q2g7V
0vD/8grFXLuz0c9rPEveKwpmTyf9CIIB48FkYBtCt4M44b6ZP6iR7yOocRNVG/LK
EBpweE/nJHRpvNhQx1U4QNirLoKjfM/h1iSvX2a5WYkssaJ8jh+VzO73DDEzfPls
a0ARHs75QGGeb/tysp0gKov+g83vfKRJuiaQAEf2MdRPDcgtDQHb/toDvfJo1qvI
9TCrv76176DlIL3p0UxPQulxrSA3s6BTQhhrmWtP/Nq/wztJjeCZsVexGjpqTYlI
3rTcRwDN99jloAwqA/F+PFVfblYsXJVVih6b9L5DeVl+djUL/ebCuhOlGNNIWK3L
N2G4a3KRYoBIsuFrF6rKPEPA4kVuSCrVE855ixfXs21Ve+1ndAhx/6NU7Dd26ib5
n1bAt8uMocsPhuqn2XHEM0b+pkUdFZ5SlXcgriLFaQ7GNTVgEOYNxF7NnLpeeoDd
UcCchbk0aMO+tg3XBD+qfvRBmns0ffZHembEQe0HcN++wyQeAmtCwm9JYvIJaB6t
JhVNs+Mf09NxRRnaI4zzlqU/MCSb1JANMlGcdy9A38p6lWuHJFirprekWbMzg+ky
eY+eyN3Iib8rme4ui3Vm7oPneGES8lFQu4UkKr0gT0ccEbguw6i80iXkg5uD7Xv5
wCnDl22ciFDxmjlHrCSQy2SR0xvACkjFf9e+fBL8QBeext8qp5NwZ7hPE/yixKOa
Tdadpv14sbXM6ZUlTy50W2HHloPW47uqsGBorevkto4OT/dRqDD0ABpsNzJX3zwb
pk8y+zHCOx3QlDjnN/lKfpY52Ngu6DVRzF/NAoUsfnA1FjcnojLOnUn+IxGg1Vt4
6qMnLrRo44l8uZAnNxiQjcGiNgIwHrJx+KKyxZlDmkJv97OeBGS5PooxM7xMYGST
1y+okU9neXow5SPY/DgEA45yDk9ZUT3lOy6SDavhiSZBnGRot+cLkc/cNlxIBvGM
5s3UIY/4+MRl4X8AJ8quRFnnQ86lPXRfKQz2WRJnBxHQMcK/wylI/w7fhrMSwgMc
GIkHwlG3ckyYL60eQ3qMVYr3sTBbFHs7S0an2Rr4u97MwyeNd/d2qM3eUMaHTZ8Y
FDhevsJGxzsQeQ3bAwPUIM7ug2THsCvycQxpiuWzZmuj/36QDzncMVPtmZLVal9R
uGDvcClQqSsXO/CqVp4Dt2MfaV3o1QsGxcOug1YzW92eys3BPxGanuuGDoAzsSnf
C4Vn1fTXVovND5L2pm7ADLbPKw8VUhykbdo0A4KVSeJ5TafeWq102NpIn3XPiIR4
flpCZFbXZbfS+UZ+enjNPiYpKoBgnz/sj1jYmlDwT1jHGWxmPcK93S0Ha7DAxmZ2
rU8GbZnojcp9pUdEi028S6q4UagzmGG9cQcM7XUH/EziXbXwGtPWHSQ2vq+RmZEL
EK/3kN0/f/yU6xsa7xKj+GOTfn6UkF+jm+3UOEyTgYDrDxCv0f+2P2Kyb4TsL8nY
FKu+UB9txHtA7XXmMNBYCUC3GwSNAb+/arQFI+AlsGU5QDhPj1YhjSHw0ct7UWkv
WkxxdEii5oE5XnPmGlv7XJ5M6ym3yr2G2vCUux6EAJQ5plGG07Ki9vYLLH9xBY+2
xmJ5S+s8AznkngNtAnH5Jed/IJhWWiCnNuqq6TVtYdCHDU+m0Nxq75O1FmCLeX0G
+3jh54+k//xfKwbN4xN1ZztjnrEVU8tZ8Vi/JnnmZrC8NYAlU3OPDbdqqimH9bYX
YISuj7U1QEkf72MgL+/PbsUVXQ/XaHCrNfATckXNge54KXBbFxbFO/X3oFH7FDIW
omd56xE/jTAEG0zXQOm8h5dQpWBRhAB+C19klorFHd162XvDf2/gKm+UH/EV5XRd
lf05pYq28KElwwshJ6eTsnbGSOgunwKqAOBvJn4dExF6jnvCuDLON1ZcVxyp3j5H
8+e981EQdf5CNm3znzMyA9txJxyyxgk0ulJFsHfl14PywTJxyJP/av6VyGYczfpb
NvsLuccqvoaVUbVQkiEtmUbdLJVN4/NzWww37SOiQ2qTqWS8qMD3Z4Ejt+fQsZs/
zyNgRdUM8hehkzHPFzhwuKkAezD7+mwZf4XDIUu279UxD6cgoIWwoPktpHPAR4iC
XqzRtNtVultmU2rWiZ4PN5go2yy/6gRreqmt+zODjFRtftzAydLCGsSOL5m3bncU
Ma4XQVqeqeC/aYTgOy65Rpac/DHhrVO/tDi+cKSqBi0V22CCF03dzPdnvINt9ykI
HeEMelZPQDmhkswjqZAGDGc7hHuiSGxVSg1H7VQIuxBIgouXC12dKx6iLU3XXq/k
LEezgVo9F22BeGn7MA5lItvYu8coC03GtPJJniJVGOHDTldTZt4vC0kscO2RVrrZ
aTvH72LGoyxJxbWzHWoUfByPHIGQ7bkOyzl+nzeYgg8t5npQJ0HHd6uPxlqYjvjy
mV2x5IGvg8Eg3XLjc5gxJCYOCW45cJeoqD/fvk7UaNuXzuAK51fJbpALqa7P9jml
25X2c2pxpJgoWOTqc34qNhrYHGaE9MXLyXGDqIV2MnLXQQhST2oz1MK25ULCDnQ1
f4u2ywQWs4ksfsV7CZF6jGby6+YxenuAspzHHt/hxwiHaKwEtZTGX4ZmOP1LVu7F
VfI7a5pZ6Bxai54bur5z5NxEAI4xHZGP7A/zKy+QFrW/AV50WhCndpbOE1FafSs5
rG0ROGy8md5Z3Aqmvndi3x0UY6SmEEY3fI5tioW2fO5+xHtUwEH7xz8/P//1ERU1
8ahnk4dRJUgF9URJf5HG+ujwwAoOKcsLTLyr3KYkVelMw6Fyd8AenNebZfGLVCNv
UA7TEPka11x+xqkNjbx7xm/214zzGAthE28/yW1jTxh+zhJd8/k9nU9OF50OJ5OB
TGdeOoY/7dtbJIJwgxYRtalNn61Ui/BD4wxHMMj/HTY7e0KAUgjb6pONS9idmTBo
myrQLf2OXm8T+5XysFvB9ms5uxEs+nXcr39ZwlFvKDVoR6yMEqiFtK1YJLcFF742
MeByniPZy8sBuszp6XBeEVaTb/lRaa8u9tLsanQmhR0ArVayiPI01w15Q/AENAYT
I3vvGMSf14Hu66ZWcU6niLJzzKMcjURqZjwSHKbCPVV2Uj5Z9+aojH1xB+8iqoZN
pfxtAJ8qyjxZZ9jfCrwDQOf2xI5SST4RdfmQ8S0hMMC8fhSQbh1o35kjKB55PYBl
+FM5g/YVb4z1AjeGrjFyaKsSFcwdmqgV/BJzFQXo6Q0tnBLT5ijYCpAZM2a6Lqe6
Mv8ntMaQrTjG/5bqwGlbSnCRyzdUwwJ7y3PPdW/h0GA6x4n2/m0DD8VEq70fHkOy
RGSu3uVIY3PKFMOR7fXWd6bbYC0mq8bHnoNmmFsdxqov1Asx2NPl50GeqdyiNGcg
bJAN5jOzm1U9k2sslCix2wWRlui3meRUTB2Y7cLdfNZk31lHrrWrmZCXaoffUcFE
IQ7YBvt+rXPBZeF/VkErChy46obMa+fIsKzVarx8S81RMf80mBmc9KzWbTkW3srW
ILPeEcS9uqspaC4r435s69ci9UgQHNt4RdargKEEY5Nzu5FITZEDXPwbSmxMpkgY
ZUlLLLsvo5ZFP3oMaR65wv6Wyi3q6ZwqN6YJN4aimzPQhHwLSXtDW7d/8/gOs1TD
TeelFSYckoKAQNbkqVUpfb+jI77YV14q7TcPirB1xkwIZtDpq3YNb5xFLD4Bhd3x
cRZyuSYZDixjuxhB00VhHzu6YD2jRvGM4zylq7T1bQ3rnNa8vnQtQB0GXr36nf+P
FcbQUVOjzheNUvt4kIL1amjtP3Zmcv0rNNT4IpwqHBtKGbi4YXIu2uENFlX9uKW+
s1nj4blIBf1gWmTdHj2WeuL5q234FcY+mTzfkqmfP7GB3akxuVaXqz7K3sDF4qDg
fcxGkfhBzzDEZhSd/R4EKVrR3sKfaGRMh9alBBxYCvSNN0Peal7gXF4O6fDq98rc
D0i6Zgo47YHlFUiLc7aFySLFzqrl1I4URrPvCtu9x2iX4hjTaPZSJ+KTQQ9TbhZp
kI5U+gwzoeotk/0GxwU2qGU6q5IT1gtqECKvLdhsymto2o5orFGsARXn24H6kY49
fyuGXcaBpOEdHJ4fshxwZ+zUBQWi87XH2/WU6RIw82dvuIbSy+f2lD5A9PIDRc+b
DsvGdO67ezWMxMQl3pE0ajc0deof85r2uf3zFReK/byrnZOrWlowJZQCVmnLrqmM
PbkeIafajklOkFsHuPSl9FmAWEWI8qD/GrUP0UGeHN7NCKscipSx0Tc7mZWEvKre
EU9RSlUFC9RCGCVqZc+5Qx8hhsZsh3zceqieALcg9rW9j7AoX+smVcUcmjXwPhSt
HUVIjQFBVL0YxnRvlS0rXKGklTpXVEpgusb12z7fQwfySV92xW1DK/jlEI3Vk2rd
7J6bLkeqcaYn1Q7t1D7oCTfcKQy9g53Ik8qpWrsselsqfiHoJpR6MM3dGMrbPBHs
S5xyREk9WyrEAaYz0iAKtIdSYZ6VdFrUDgiBEKjnquDXYscLjy9rpu/2W0cEs/Y/
Ay66UmtvUEihNCYsB44O/ylBkWhL1c7jbefr7NNAYCPMWhxmXYkLRQ0lwfV0PFP+
6yowmeL/1zYk2VsP+wTwvam2w4HNp9AJLO9Lt/P3CfSZV+a/ht+XEUgi6JeXqmhq
Keerp/AKzprHYw5M92q48v2nB2dA81Pm9ZyY/KaZIPLFyBPFNx4XNOvjglUNxboO
AQonNe1gChGXR5R6uJ7Ndig9CwnP4Rmy4CbdX8Y+Xk+3NSLyL5/ZOmO67EECOpGZ
+5UPkwyHiWL/rROLTkvvxppXxtYkCWeQQm0PAGtB1NqWOJHETO+jKp8p9l4OqGTm
92YozYOLh86UGOxb/iGO8GbaySJqfp+aTjOiElATkchEeS4Rfg8QHqOM3fHpCt9p
JLAMxllLyPQfGdTdG3CZ29N4hr/+tEYZ4qjd/a5sD7e5MN4ot8pNiBE2X6LLFvHY
jxxum11/X2yucPRuc9/6te6aLNC/fHqWjKn3Vmb53s7jqphIzk2zW+8tvlGyi4sG
T84dnCOrbnj5pYYhFrXwYLsKj6AVx9a9TmSqUElAUVu7m3+y3RFs6LzUVhhNoDof
VYfwAih/bV+IdsSban4bbWkLdW1PMVjqVVOOwJjZQKHPzkGIejTPUrJDdPPUAvq7
o3pYIQazw/gI2DlUJiAllz5hJwtvF3m33YfOTIKzc61c6pLf52l4AAg186ra+2bT
l4VmdY9R7X/7s4DZVG69ohiHDhMGXTV/kzFU73qNxRBGRKBbbDIL9kltlxTYVlKc
3oeQ8/nykYp2NMJ10YCkXwJZV8gmtePe6dZ0dz7rz6zCiaiptPU3MF7vwy3CJJNi
I5cNGsiqgYk/d6G+Gm61GHkDGpQRqQo6NbaqzNgvw1HdMk1e5p2gtA1sQ2l2c5wV
47Y7QowG34yNFAzTBGUjZeNSnRcZX5cOhMXPxcflEsL3ZN2FT1rB8mTGDd2QBDII
SXDoY1uzn40iKgStMN6fITDKRYpZAEUo5Anaw8eBPLP8r1ph+o3dlFZ5b5pmeYLy
5TI6lI+MmzxFlUBG8MuWE+NcldZ1nm8esuA5gAVmGMYzXtqC1MejW+aNmGkpNAkm
B5VBK8FZPzLun3G1dhPXOJFrBEBb2AIcLSmR5gW11AWo2fX0KIQ8UGqG5iG9WZtR
MS3uTJgYRd1+zXDFXkMFqxBfbLxj5FJbBnjhqU/IZCYf4VlmKfqN+Yq64Pz8HjFN
uyHPDXthsnQYIVopFFXoQw+Bu1p7VTAO2/drV7A+XO4nUt9AtB/LDH8ITAyNGlhd
hcBrDH172EWrCt+STnnOoWIIW3ywFCykcCRu7E55WnXEGIiH9IWwhGp64d1FWp+O
/3yMR2gmENlVTkb9QCn48xyJCod1vyMvpvcplIqx/Eqp2Y+T4MfhjudnadfQABFK
IdZNaYxa0ydoW7zSQPwhLklxw8nnTyVRIP6JO7FoEqSKemyoVcBp+RFcbunlhVtW
tJRIqIODOURC+7UwSjtTueTGZqAIhyplVMn6LriPTLd+KHAHFspzA706vzRGvoWK
tPMIMTTBi6k5CBVdzWQ4sDZhP/l7jxyde3Ee+LZrzrn8+noCR/3MI3ii27ZrTRJt
TF2tIJLnw/VPXAaxV/i0ZU7YRwElMEm/LKmklkO7TFC9FOG74DhUBYWla2qOdEtk
YjHh8ouFCv1T8tSxi7TTbaBScj2IqIqirgCohmt2EOSlWm1MLI+VoSefzedX+uDZ
BvO5ZCUHBeastORnRd5Q7sc0WeXk1Ly/QTkZW9ZPq/I7dDaXItU4NEPguSVFVmNQ
pSkQczPEgNVC3I+tvjcEyrJVRx4ELsKDubWzrTCU2TTlyZbQ8ZQqm/RBe3UVz4+y
KcDY1n6ihpyBhipdfBFuvLX465kxPdqjwdrcl4oZgkZwh/Gw0mU/CKAhgiOMN/Zn
QZZFmZT6+wmCKKj5zyyBzmSNdKkAauIceiaofvFGDQ+wmfGOk7mH2eILinKUvsGQ
xJ2N1vEH2mOI+JkHw984U11/UYmeMHb+2CiJMsl7iLWajjkNI59Ns5NRcR9Xc1XA
RjbL+PQFmN++2ejtJKIQrnQHPI3AD24i6q7NtpsRjE2mghf4agbwL7I5luJKDKob
vbh2Y72+6MI2OTYDdeJTq62FuSToL/oWF7V1phMo8xog2INFAGZceRPOUDCm1B+c
su5dxjy39H+7e3uOtTUKLAFrzrdoKhM56MvCoATkp+OU063vFl+zsKnFRnHQ621U
QFLY47A0WAcTVfUxmp7H0/lTxz6RwETA8ZfJ51gbF9QNGQUSqKsqHG0+QytyWctv
lQ/LMqz6wwZ52cLBe3ZYcDdIkSReJkD2wZc262dmzc3TkpGOje3OcgCyMjr8xpVm
mVYNFm3fP1JWtcJzrQSdIIMOJe4Blxj1dD2pqEJxlrFH/7Hh7jAG2GXrBceaRLaY
EBNqwFyQ0CHM054I788EJppOLojYCFPwMe3IPvurcdPwlPKUSsss1uWxGhMzr/8E
c6LkVrL863zeG6kRj7/mPnYwX95ee/XBxkexXLP49SBFuSNY26bPxEhhV3+ieH7D
CBJ2GNEWemJyesrtcr8xOq+PdeiLPU7zghaUKpKmKQN8bYaN6ggabkYjIpqKrjqE
8mqD8xyoVez/mCcKzpY0jxyK4l6eToHCQ1jyA8Eh4tQqhmoga2qKOOKMgfcJTn7q
Hkl6uhHfdu3hZ+ZD8BbW6uNy8lX4HrLSdridERMtA4XJBydpY9LfcjyH6qcFXj5q
ikqaKUI3cENKREoxd1Er4Gcyz/6YYvrujdtLYg2nlpqpD+xurFdjPuTLmgOMqQxW
tXYduVkE/50iIVBTazF4a1SgOTZPqUznkGwT4mDys1vYQIDS1ayzp9V4G/TtKHzz
9aRFxFi+7lFVNQwLKa1u6xpptlSSYZtVjlXeJnTDk+i/Wi71OtmuuWxoXK5WmVcX
KItx91l7I0TonStTewfiR1NX9m3mUPSym9twVL6ZqPFBIAJvq7M1SrdppgTHB+W/
e6724cXaGIDyknydWMZavg==
`protect END_PROTECTED
