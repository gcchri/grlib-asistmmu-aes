`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U/WjX8JAwIxOGRFWs8+j4wVFA5OkW+CZC9K14yAvzd7S0FRoF56xpugNlnvLObUf
GbeuS9GuIf/Q/OleZGfvbKXBwPGuWJWkvssxtFH02Yev88lXa/qdHWNzaay5sZ3Z
UgqLh0yts/ft+xoVp/LuJR/EesNyOKhJAN+XvfeA8iJkceVS/wNYaOlPBg7vFhX7
bvCPmhKyfayp+4sRXRjy4brNQzXtF9xC4P+2wAS1tQwFd9RSrbT/1niXhDMmg1Rs
3PjS0YHPR14TTrDeobuzbQhQbjkWpnoWO4fLD4cjFiTjv5cIEL0FgPZsMAy0G2CT
nxPvF4FhB9AES0rbY31z2/AONu9h/kuHmZYQcDjQIuUXLPjnsjMS5g0xLDJmlrN4
HO1wkWOQrUwb0+S5AxUV8xZ1rTSghZ+lS1V2FJUMTJV7IgtjEHhwDB1Rq2CJHo2+
A9F/lb5cuTMKHJVhVJpNqM4y1T1DcKV4UbVfhRwzXB9alnFBefP9n46IjidogrBV
jICXV9gtIug5kfpEC3ThGt+HhrBKp+wnY5hm38memeOvWebioY5+HlboMKPdcA3A
4WIGuwEYgddQcowuM4WZrkTefdoTNY5HXpDSMiDci3EBEzl+1I0lGj8OIQjzorKd
CiDFgyyibklFCy6vifNiBaWkXdwmR46D7wEuQ1kKi9AuR1PF8Rb3w5RY5pZYigCS
3M5yTyoG7h3IphrgGvleOtGbNeVHKxjf+S8Sv7r44jJpmTeN796vV2DEfpMYgAgK
cl18/EsFBxIp/HSLv54nQjj84JMcWpYhEV/esyFwuEQ+6xjdmqRfjogCeqmTsvw4
6QMN5eA2bB9khixIQLtB5zLf1IkwMT0ObgryymXk6Y3V+GOCy1qsbx1ZD6ZZrqbv
UeLT/klCy2XFVWrg96Q1G5xre1/dIX9YncEnmWuGAHEVZoTHTAKbNyJTFfHI4a8g
FfVr9FbXsrQ1z0oKxthcOweiJ4p+842Q/yMZE9VmTN4gfqdf0VBUZ9qROuQd+3p6
FLx8rUI1Dj17OlmBA+VfEI35mN4MMZPBH8tdLHtSQJ0VUyaVvilOEmKc697wwGFE
pr6KENDgqcXSd8Pc4Kopsip3jtacvwyssV0UIosRjGlB9P5IQ9RyR9MYNIIHssfa
7WxQpM7kD9AwqvFhBG+P6jywx3S9hxqcD6ftKvFT4kjVXcHwcfTDZ+m/8n0T+x6p
pC4WeaX9cmY1Na0fgq1a6Qo8UCgDX6o2JXtL7BI+8pF5zzoo+3Ix3SlY/K7NCXpU
r0VAMxFKF/E8oz+bsoAJzeuB5RhV8uVCz8unr4+8n/aIIvWz5RuSlxbWt25GK791
LeQtDAwBgD9ukZ905f3T5LwHAJnxWc3QdQxPlEt2dfC13GzmDnBJ56xyfTLwj4pg
+EjmWGDYvkN3r7iDinIKpJr2Etb8IH4fIA9Dw9n7CgDvQHnaGs8XwHsQzmk0mqGA
f52Q39cOr17P1MkU76OKNwQlN8wfqhUjc/hXFR3X2W6B8AXEsTppUsdTYogEvJEd
KoboZ9HfmDMzSvOziwTN4qQKS01OMlD29aN4ZmpgG9eS3uuv3vHz+ssM50YTXt7S
RoYHMxO3j7UruuAuGeDKzZVvTPEZT8fDpoPC1ylhPcLDUn/+o9ayzN52PBgge56X
4SLIJjxJtiVmx8IQugsQJRPAeHEjuYYU5zygPsfQOziaRBXj4Wc0uuwxyPXJl4Pj
LVWde6P3aEEFhaqUpIiAEJFIW6BV98+UIRQGBNIJb02HB8kTvlcCuWvHUTD6uVBq
3yKHmBbX/BQLy03HnesYP4UJI2WYDksZqIPgnyeCtyFev4mHwq+NS6sL2H0UYvDa
SJET0Rqo1kKFIl/a4BIbASpqYiwbkiiqjMC3nOhFJD48QIyoWFTesGRTFDfNwD9H
nBfF337E7epM0hkgmgLvf7SABQPmO8+h/Mqte23OFzrP7LbeBV+aCHcVFh3k5LN9
8ZgKlnWzcGP9JSAFQ0Oqu9BWELiCCMCtSj7pBGt7M/TKct6b3bxBCOrMwxeKl0+u
Bs4f6j7YcDOf7GDNCbi6Z/A7nTFyQFjK0C3WqRwmEwxnaF+UrHZ1P+q1cwd2WV7z
e4EGMFYtaOw6uZbLOD32gkY8dnZhLchwUJ2DXpaRmzr9xdGllsJ6vyJhWSBki71T
t5mnesjgrhDJ4qNc09rB/EHbfijEsMKN0FbjLaF/WTOCDINMh+v05D0mSdxGZWQf
Hd5aI9NDEca8OyzY2OPStXwJrDqYM9XIOyeLyaJX3SbpNCa6TGvpJ6AT/6q2RNOa
5u39rGsRti075olodhhUlQKKKl/8kOFJwLyLPYkcIFUKNmNffyTFIS3D5HkL8pBH
6lewcIML3yKbFg0OzhLAcNVrFErj4k2T+ElucgEFxEgA4HTSOvj+E9VH4IRYR0iY
PJ+1qTnS9ss6tSwPMVEPCPiwwf8YLEs4qkMa/8E8yooKmxEZDtrk17uc2wZpNuQ8
9s0A5EPGL5oAjzoN4dDWmPYKXGkeIRvcWxZi3TXy6SYy/vP8MrmlaFGC2BK9Dtf8
c4krLU88kdEq0HS4JVPEFw/OKi2LBwWXgBYgK7TxfHkYWh39tYyJCsLnONkhk2Iw
HrPf8xi1a97okodcl5O6ZKO9gCt96dFZ5bMecoVyVdfesJRQkNLx8EdqnU+dYJ/u
MCKyzc3Sjg5lTTJxxih8J/658DNvEtLFGEJiY5cD87t0qLSo4+Tv/7SlVlxUiYNQ
69s3/dVkQluojBuN/GmQtucKpRePSVS2NtC8KXeIzjRwRAIpeAZv+LUzVx2Yy7h5
GEfdZZVRe+UtOP7BpInZdTCaQ8qh8Y11Vb9MiqUL9WxeKDy2DYjhazrI/gaYPSuJ
VtAq6yQLWNbapbIcWqYd9+OBDVnwBJ40Xp+I9XLTyYD8pGcqLPwb86ztIxkWn59f
VjzDornpOeIOBMdVPf2Rc5P88nTnmJvVXXbPEDW1DaROnmaLguINt1NsW5dDphP9
TAnlewZnXw586aIdEsNuLqCkkST/Qz41xggQMISlgpCQCl+8H90L88O459/bv+du
d2B64zNE8N8SWF8MzaGUQiQMux0SR6DaSRXghSejL02ANwiCsLEfWseu615xf3px
JvtcNSaVTFh9Vyo7AP5+wG7vp1wxu63ZQanD8mFam0QmZTTXKt8HyY+GP2/UJLh/
M/pls17ldxTQ9cIF4Gq7iX3vZJUE7dFJRF2qka9M9Ul6n3QaiLije/3ZxEjdJD3m
GyAB7DeEP3w/3KD3Bm/xhvIAgtHmDRGDdiCTIOoHqb6/xpd9heKQrWhLLHbvhfVO
oVH3Iu8Era6DRA5lskN6+EwHRlokdC3xLU27tLRJz06HrN+AUbAl015drUAfa9N3
JsRo6uZYR9cfUWQmjL7D2f/brWgVHO1fzw3TKh8HrxqZ4t+L9TGojxnbKaEr6Qkj
MXM3a7LICn54xMXSxfezzjGDDxzOqRFguUrnFBFFko9qQ3YbbdnkkXJ0fmlG5piV
e10M3mJwNwLDn2KFn5K6G6gByAR/zhT4xKUG0IfjOM+TWx5Go0Lc/fZCwDfyLQk8
Y47Ndfhr/300DgEM/lHr5mFNg/DGA/RcZEPK0VTyTDN/GlPDXTTvDvEje2EEGMob
hQyQGkJiM+YeYhsApSYspWGzr+gqgkjAmNflQJFqZS9m8rI3OJpmUQc+K8A+ygn+
sPNlVZBLzZfch/XN29kIz+KxVPDGmuT+cD/lT+hqv+79pzVsdtiFieEl7CGh9DBV
qQ+oqCUTff5o4v4p2wBIOQ4XoH/dMlARObIoF3Ud916zTNmibay38joYl1DuoW9I
oRTU8vwVBxWUUKYPMT03o7GfGLlpRZdJi+uhrhXlBBu9++ubUzTajCRyeYr5MEh4
kaP+ZLZl10KFCJhRJhM59Xoo5iZPpQPW+bEuMxTG0jL7VLwqUeOigxmMVY/EHmI6
HL8FgZqK4OfsR4Wx2htdPQa4IwsyYUdUqMEKCrCcVaQzY0QtR/O0FGO3JySqr43A
0YXDHv0zgdR0uY79I/JFJGYkZwYFlGaFaNb48TMoBoK8onP/dwqcGwe3fQRS6mUV
FxuFs8XxDByB0s+Vq5VvJKqMMUfKpWYnrV7GIc4rsk7vKRm550GsUYcdbOYfpM0o
cZYXZoK1o6SiS8Djj/4sSO7Slq1Kg2Ic3wcelkKk0IPMD7WlQW4al/hi+F/E3tQM
uewqcDDVApFKvvKyvMpjpA==
`protect END_PROTECTED
