`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rQLSR8DzHhpzw7J5ey4318nFdU2gbINcu+Kpt2VRzfRmlekQ98AeJf4ZdZ/zdx5e
Dr+xiJN/T6dfavtdtAhFWilu1DjSH5uvon01H+5UDkRn637mUCKy8Ab0ipqcJ5Db
NTUQwqtU6XNWa4VyxdWc7r+u5/KNRr9h7Q7k7rFY7Hx6CcZeBBU2Eascn/uVBLD2
Sat89j/ayID2rY3/sayNIfjjI1U4Ur/qQrH9M03wvB0RKgfS3Z4Ehp+bVIK1yh34
ck5y1ecCalrORxA580CZt+wLzbY0QNZerMfyz1N78uRU6Vw1CVFVfbRI/ilFymzB
tIJcgu+TH7zCupFejrIIt5CA2v/TbqqFyM/TbR7qjRrEUfb+EavT46Yzcc5k9twz
bvHa/smjtRvXnR5zUzl/6LgVjVOGQaKGgZtfq1Jsfc0HKdAW8OIMeTK08R4B5QjP
Ub/YJK4xtv/5piTy7ecOIxZKpx8Ujadd1JOP7TfrNYg8ooR0dJw3fRjA+YvhErEF
+IVukoj14dfSZ2J42SLSVT1joVDQ9BnjSFFF1gXnTlfe0XzYfuIJ1LCQCkROxdr8
9kQ8SWNdwRacaWqaEIb7a1p+frwMtlMxllpmFRLqdk/RsLo/a8OZDA1YxJvnJJtd
5IQ8/4dX9r3UAVi5cTkcPxdscK7N0mE0BSlBaeZBiEmTtKiiQ/Gcq5fOxGmO/wnn
/8cjxXH66ObGIY/CM8UHXkD+9FaZWUJPz+KrmK8E+KI3FjSQV8CEFMdjJ6Cl/9On
G2Uo9QDWzDh2QwmJnsHxmRbpBxBDvcL4wiQy3ID5Dk6XiIBIdWnAXXAzephjMACR
uZhnlQLNORGFzFXzACMMzCUZu5hwq2wYJi/xVzD97GUwG7S2+L+WLv1GC6o3c4AP
qY6KvSJ9g44hAuFIclT5jmXLY7aP43OLE6K/MJN0XNaw4Hti3KFqDIreFjcFIqp6
Ph4keetZeooeR6Y7g4sAtMrCfHR4sj8sYYnb71xuApt40oJdRJehoSbIbw/7GTB+
Im/KrvI5oxWtGlPKRh/vGU8GKgWychPXTLE34XbJogmtDMKZ9xEvXREIzn1VLtqR
fuWFWxstbKER7/9t+gQFSy/gVXw3wsWAU8dU544yuWe6BGKXeLKKClCrBv/eiIPf
gWHvUIYrwsAGN/mN7huTeJH6RD0GrhocyMYVogtjpjOQ3s90iiAfPBoWHa18URqX
I+KSDykjShbmrl/hrtrvqkaDS00bNAEZK4s+XaFpyJfTXIxq1dv8GhWDKswaQNO/
4NVbJlAx1p3fZJMpn/SOslYvs7NmsNgyCAK7KdA9c75IZvC+xeuJTHRMLI+Cc4E0
NbArFQ7Sow4xfjS7zBbhmm6yoqTixitSuRO2r0Q8OIDV0UDxse41yN5CGgz+wqqb
IPDb732DC/ZpeP834IUd/Im45esBOLh7HcFV7e2rycA/hZzzlbhLEGkIHEsqSqW0
iJ092vmXjPvGw6T88ipjvuPc2lY0uKx04VFAQ/GYb1zUzOeEQ9DfuNT0H//PJS3f
BZHSsi64YBiIfuC1CQj8L3FxcF1KfKact87xiB7pxAdCXKbYCqi2KezTJEZpNQOZ
S0mBhTNg2t9kJnd9qN8Dz6lvX5J/0EW+hRsxcjG8I+eTy3OPaI+ykmHAD0DN9/Hp
jdfcP3Ba/7X818I/bgmvT2ZQYn1116XWjbabjSJsVaGTElzG83WZpQgPY8wcc3Xd
gkmyly0f9Saon2osMdjBStyTLdACcYzrkSZ580x7XW0jjiUcsfcQi8mov8DQZvs4
72derSxJhPqTuQCErkP1PrCJnt/b1JR2sthaEPOjdOG+3fNayHtsG/jDA1kP/rgN
2SwX5CpEYE0L1NWunkR8kEUEzc6jRjCkxDrKB7HVUQQw8ps84zOx+w10WMOqHYtR
VP4l814T/twIvxBLNgfHggAOCadADySSjs3qDY1DlCPIGJ17KY+J9dEuWNsFWT7p
afI4PNoYJRcl0E9oVt367qkKLJRH73YxQVCeYu9WN3WIgxwsG/mm9cy2ZXwhTaoK
HatV4EStJ2cdUcqw0vfT9EtapWqQA5BmA4tWyU9b1yz8xH2YOuo/CzwgsSigUB5E
mWi7TPGmY1WBR2mmTJvgbZMJxvkyFH/i2awqWaMLM9faDPplvyXatrkj2qRfhVpi
mujmgndUkPe7cJSNqKzrg+bkOLsiwvt3dW0J3v76DWV5a9JtzExHBUlsRT/BLNU3
m6kupOYBB5AC8+C4vHyj8CYkaaD2R/3l6lE/A7VBJ35AQZyStzmlBElUBepx9cYm
5wZgduHkUKwkYqyjmSYOaqHKfGjEzIBeE9HtfgPKtNmWVS3K2cSQIB/KfMxix4mA
JSZOfkoqFM5rOw5blTNjN1LA05qmrgsKsgiYXDPD4diQm3Jw9D5qzwyZxFnyR8Vz
7K3GS5npqtnlOr3wh76hAP7gowMh1qGd0mUFJ3X39S9wLaxWGttpNnGIpRYbxtDZ
15ZKhzLTvraUrwXjj2EU34qkFn0Ti/F8nya+DagvFeBZF82dfE8hcEjmy3CA9VGm
wk0BvapO7oiA5w8nNMeOt03DUs9RA3yMATrSDOraEyC3Ze3iCKyt2ZGketwxLUkk
324OpiLQC11YWbayMUqqEnNxL+fNnxA+TVn+7WplnZR9Iyj2fVRzHKR5B/3J+QQF
nNLCG26D/q+BGsB8NhfJAKczzqWKUyCT00LZIhaDYbohgxoZFnL1NuuPzjBzXwQV
UxyXvzjsZRmUTLDcIj6gyrChkoqIQHcWPIVKapvfP3gY2MDZMobaAzmMvd3JeVOq
8wr5lbTKZ/sWiirK8v42Kd6/znBmx3MYgCJ0iVomD0ogILTlACScKGsMcmibX0R7
0gAjm0TFIIKO+dHu3as69Il4NqvpBH0trCh9C2GleBpljbLdx4gEIhNy+zliMJyN
vOhTFu01tuLbwDjrJc7QNurV5wY10ccj+ydrGWCgh359yP5mpgnxpOLxgUrzNSuF
3GBLwLA4XyKH2a1BW17Jd/1h7jNShbP30sJzazB3pUmwAKEIWy+DgjU+1NkCKt9Z
LMan2UvGpGYQS5vWxWkkfP+/qQ9uefX5om83isU5ZzGDTwlJ6VVoeo/rQCIZqbe9
ywWhYUc2Y3NaxFfisfDKfbNa7CYrtUZDiNOfJIoJPpaD+CBYwUejz1TT+8BWO0a8
6JCv4GKaAkfSaBgu/O+CjdIKvrexSSJOQpA2FiPeiR9yapU4xVLflKnU4N5B8inv
13zMsQlDYGXtILS0bP3iAOTEmFU5mENsGdrYCNcie0FObfnEPxgm/6+zOze/YDMo
3bikK4SEdgRj5QAelGCkvob9IplXQzIorHs+7azWriHSoI6W3GkrtgXuh8hZvf32
uysbyDyxuBmfRblOoTwI5KLvGf4xYLTmWkckqBX64Wquh3fA/a+FH1Z/drMWVXgk
sFMh3cwYcI9/NK/oqtbA/QM7XvYJaIOwfnbIqnRPGTXwD8e5zz1MDW2H7TsYL1VF
2qSip4XZLuyqCPJnajvZB1osALadQ7cQ9Ff8UkuXDgdJSivjMvgNDCktvFOvIOFj
EeUDYVMEQXpf8/ChvMNwHwVx33zW0CGr4jyrTs6Y2W8GjdgSZCb7j4Kr6Wf5oauf
/N3p3dTdtgBN6zwBe6NxPBNA4rTYl0mGCqXlksGdvLV5Qfpgh7Vao8hsSU9Bd5fO
xB34KD7KZurZdyNVHTNwg0ukazN/t4vEUAkYanxYsJZ8RgSqRDdpHQlfgk92G9lI
z5YYEGva4m1Zd83LVrC+3ygW3tsmd62bcrcdbkWif3tuncjeRuEW3oTIevL2X09s
8eUhQnopCDGdX/g+iHk+QGDXXjqKFWqBTrN/e4tj5GdqO5/fBrHciulALt4quRnS
nWRXEEImLubkIUxM+90LEiYFJxswmSNNPb5IaDEjhdTYMaUwx6jQSnR07U5Uza78
KpZBzjOMYU9fqYwYS0il+MW5S8mfGH5k2n9bLHDkwhIy8lexyHacYenM/ZAtkGrC
Q7W9yPsCXrizNy22ln/UBymLScDyZk7+r0DYKX5oWvng01DXb1yM2ZrZbT+NhRwn
FTxA2mbcVZ7x4aodzcHyhqEXr4BxBqj47BW2Nyfm7vxu4Puo3IrksPvopzgGHm00
iyjuZ5lHjatHu7ROac7rvZUh4GIkHJboH09BnuEkegRyt2lcmIXhVDlYLBe0msFq
hAvJ4L2ycQYRK7O3TzHI1rd6VPd9clRc7F4wOGOlwF7idQ47As7/5vjaVR4GdcmV
/3dL+7oNnOEXl63A8NLcwEZxCJlkKfaAynVwMjMGXjXlFmersqkVFj61+HGB+3S7
Leaj3ofc0NZ6sdrJgk7usa3glxTjmtoaHJQLOmzmnDOi7etEqKMmU47Ge8yARxGr
pXUHv93rK9itv5weulDZK+nun2R20SyHS6W8D0RI40WZY0+kJuntrok90iYzGSik
1fXmkBejeufuYG3jiuybUNL8TE3CnXO3rN+MXY68BtI+J7IUJWgAsetuuxB8aYXQ
aSgOqo2uZmBTNV88yBQxqTAQjh56xNy6lJ6DPYt56wChq0ckGPLalXxDodtACZWk
xhSwceMjXrqXX0wz7VRLppcTqbqskubdjpwcO7y5NkoiHkZtb6geMvFiehRQjCBI
R0ZDMDtbxC2vSJktgi/xxJ2mUCpPST31uNUi0yWy1WcSsFywfDv820N8o18xbct9
EfzsGkfEfd/sBnL1BOYQeKi0DUMnC/etzQRLMkjNZirAgV6tSqL717i90nYyJVP0
G1WsTeT8EmTdq4grd9mc3lOvJkWi2NGuyV6wR2Ksg1VXp08HX/9PMRyJ8Atnm6a1
Kn/miRiI3iGHV/B4ejmUblnWTkJ5gzVbe9k6GObYePhjU4RGVpG7k9PBP2H9H7e4
QRD1GKYXYCdBLUrTF1y+9DwHna50g3YDCEvad4SvDYRqqsl8otBsT/J1yHk6oHcK
9IXPqR+GdggY/RQCHg9z5CbmRjGTl9JkqXJN/poiyL9zKzmhxK4Evz7Lr3/lKcH/
NhClbcMyK+wg3kMViwncS+UNbYCqChovVWQ+ZUjRBeOzJi+mMtuoIFm/jt5Bos/D
ppGhq/Dj44+J2awsWFUIuTj8XmCeQ8MxwDHi7/XbgYu2nYYsF6Pp8Rw+1Cb/nof9
EDwFG9GH5MzEbXIktdKppBxkHIF1BHLtoVmwEQoeIUaVVLxhcHk7Q/lmAEiBXTDj
BTzN8k4BiICPRE5eQsbng3K/1k0lBfni7yzQIT47Zf69M8rcj/ob0+AD5K4pO1Cf
fAduzTFMjtNkSO1whYINiAmatpUEhL6FXV4PiL9uQpG/06BJU08WYEmb+h9XnRfE
5Co0Gn4rroUiONiHG+VRhpuhEIhv2MDpinuZ7a8cx02E7PvO96YVQjfI+4Fp/Hd4
tnocTtEEISZEo8rU62bM+OR706Qa0PbCTt0kz0YsMoeYkJWrWSI9qodQFlleZfuQ
3gnRmMa1OtkgVIfPveWZYVpa2Ur2pXEbPDcDUlPR099EKwLyBBsWHuLJnmwVDEQa
bYn71MftGLCxPdOmG7FR2w3YEgHif67grXDfh3QoLNa0W3fQklp1zYjU6p9SAtGA
lMJIQ2Mn2bVKhQsVQBnCz6AZYIO/pfYp0WkoqkQXr+7DBnJq5cGiqG0H8Q1UswAn
K7pMYaB2o3WhsaO6OsJf5/QxFs3JvYQZIYw7SQt7g664dJWKIdSrLVH76NYT/IzH
16tjwGMHAVkEJHvm0gl4J0m0wL8KjYVjICOw4TUQ6iGrnom/58YQ/EbZhIKwZGZi
ikKxke29m3zUBAokRdRxHvlu26Iigv71BSrLmaNQvs4m4yi20e/XVksUWxJ3/Vj6
EyGjkHcIVBmenVlF1BoWYKMdAKGVaFgkGlkxwYTVl31cR2zKm6kUWq+qgIdCEn6w
B00wLwJGCobIRmm9dtw7kz/QRHwmJ8p9yENKXDLbIxY5rbzdV2whWk4+rFHPsxVP
yxg4yRfd6jvV+zKgk3r7fa1HBPej1aY9GwqD7QE7sCw2jm4k/Gwm/xXe1/rLvHhY
5H82n63kQEHsBCPAoSOroLx4EAy2qHJVRchzASRI6zW4VcLzqx6p0/1xun3tIecn
vK64QLiDI7gYXf1pX1HEK4qRXOW5M5/FQKAmSktSJ8njuh9XaCefgrZ/4iIU1ZJG
y4FiixLa/LuIdutFFwGlEN5lCyxb5jYH9CUd5SEz1X18fEUDFi8HKPNZj8cKRLfG
yAbcx9yyQLLZ6dR5DtrX7FE/oiJZ0OuvnpB3IbLU6+uW/5PVzqvFvqkRxGMtbNcx
jpSieb2vuEwcqglBq/+fTVFqzD0Ded1OlJtrD3vlL5qhWiPhWhyNPYCV2HOaipO7
yKj5rhUB65rRxpb2+XhHD0JeVP/1jyQqtOn3dNwGhwEvQy8erYCGLQIOf6HycC0Q
k7vG3zjh2TCWdBACONcB9x1LvtrDEEPw8xW+RXfETLunFpVD1gAV6rm1gRDW8sdD
Wkdjcb5oSk8wuLKSF++lm4NytQlPnf1jhNTC4+3ZCY0T0+m98QG0n5wP3Dg4DRyf
p7azA1Nf6xAfl0eZFpqO6dUJ9I/ubGpiU7rdwpTIYyl8zJ5NseRrDwvs7bypu3Ij
nr1wqqZWFzNeEuzFP2dBVN53R+1IKBYY+HbMrBopLkiFkFY21zwZvr44qQ4qtOAO
IEGjsf27ykeD6E9jBpjNjjojjL3MlcZPB3+JBYp1ViUpt5IsFINY3APgioYE3L9U
UDR+ymhOfctZwKoXR0fDXOVNT6SAMrlItmfRg1Fet3UVBiVR5MNOTczH7kInSU+D
bgaBfu6Ue0QFeCwfrgzMcw7kJvUBGZN8o97GE1+iGIIMQ2BtbLqKT3fghLaejFvL
V6GHy7b8zevWWKIf+33/ncXYjEvyiMwXgAt424LHjuYjkfP4IiQ+qNd7hzC/rsSS
fnJAMWwaO4FpZZYxtOyGWl2Z8xKj/Xfw37mn5eXwWa8lMB1kO/J79UmNJrHGSSCp
S3x4fqhaOIK9riFjS9vzf81go6jFi/hURIIDB0C8VQUqpkiVLiiFgDun6j51VwQJ
+PhmCu61fWLmhM1FmkibzLhqXUJDjJjS+HBsUTbvytcVELCvLoMgmgzswtcpdMDf
cfZ9Mybd9F2f4EXvIcDkaiQ0BJHWuhPvH/uIDOjB19vzcUuii29FQPWUJopVVIeO
c6H62t5Yc3YeaA+OmQ6Jqa8zZeCbHqYIfKVwyydcB73JSHTT+cgZxUHimI2JHBkf
pueJWik/gJnbW562256wcko/ujnBtaHp4ihSm5NhqGH2VfJTOBhBSpAnt8Y8WtH+
CxYmsKwmWPrxcdw3DOXKOlXOhUNL5A1PigW8oTObD73NBXvpNGBJ6zdQ8eFWim4S
SEFQQuFYCU4YhOTSRR2KlcAztg4tyfhw9P0jsW4rKcIMS2Q8a4whC7xoa2Z6ihIp
6+QhivsntUrL3jzOu+3j058r6qNs3rZ2EI+1lG3wmYHGmflZqjP20Kygfe/QSh6y
WQp4l4zY+85MWExGhL+AkTpSFjoCTIB9Yl/7WD/AQgkXf/mPNJvi74+tfL1FRyOh
7o/z8hdQyZ+yyIkVe/dD9mJCp6MXnkZ7l7nBlWST7k+vE8kdUplnLotEXmCrKPzK
7PsdATFlaBrcjtiZM2FEn/JusWSp4EuY4Zu36l5WH34aTgihOusq7hNkKAvwcbhl
M16NpDaTOPm76NQGw1XiuzQKCkWqJKK9JBMwnyoKQfU=
`protect END_PROTECTED
