`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tbGOm1ae68HFivYkC2q+ZHd7wLBvxzkrN84fTDUOtQMwdupbDDMY253AFZI9nqxo
kscxSNK9fkN6HXXSAEiXzCpX56YYtoW/ZvAiH9/tvLoNUrdTRHpWxjJnLeOOkz5s
DJ/BiHQ70enZ9v7rey27l8izwPGyLpuIPEkiFvospnxWGycUfY6PZyoc3pLkIwkP
u4p0yFE68itifSvKV2WwgXmtwrkD+lHrPUvW8bmrIGwlVjLNXCR2MVqbAt8/ukrJ
Hns6u2DInUEN7WWUai/O4sKAmvUj/gl4ZxAQU7rwqjTeYvK8QiBcXzgfNILZQ3oJ
sSRkBbxb4DmpScdMjGOPG1EcTA7cOjkndIrc4qCu5MYhwjWzJnTxM1YNP3sy53lK
rPCD6uz2m+cCYX63Les27GVdCxjyTGgPGiFF88h0XesbKPUclzPdAMVfriEG0N1+
NMSvGbkNVAS/3cmrjlg6WvmW3aT0wDHkwzSmYZ3U4b42+ms7ecA5eZNsWbngjdll
ftDrGBclOqQV0RHAkVuyyHJI7NQgU3Six7WhryNwxD+JkTCnh4ej1CKivNf2WHAU
bnO3Roluw/JB23hVxw7zds2+voQZx4bUux9knYym2t9B8dXUmhInBgZtXX1yvgaP
P8endNH+hiaaFlsBCfxm3spvCzHHg8aDuDEYoZkEYpm27bQBaZYQYQoxnX0XJDfv
s0LysU3bWdWLm8S/chmIWxPlxaeEuqcbetYq+Qw+tpN1Hyt0ZGW3VX/Kgn3QZx93
qspnrtveI+EI97GmqJjyQt4xCe45CdBOob+rSLv9X3ytaB6Sl2UAQh/6QSg/6F9a
xX6LOeexsDx1pZp9SBmNV1E3X3nC0fmDvJeSVg9UsHiB7eHgAElMQBXA9x4wqh42
WSGlJ6XrRC+Q5SS5fv9daSdDLyiRTcpe2u9YdRjNRMxqwqSp9EIs0jcRK/KQ/yRR
wVDXVfK5I8r7smc23mfYvDVE+1uHRVSKPx3F2r/WOq2RWb34hoY8O1eRLrhfTt/n
R6/nyKi1KAF/bvBpCCzkciJ5xrpoJ/lS2qp3KFTxgC4yBuPHMhuhauEhA2x8C79d
WpX15aoASzHOr4aN2NR+w4Xa3rT1avUgdznfzUU5xTyu8nkHD9CwOd1VjwbBPVoi
M+VB/hDebhVT2Oef4BJc0wAXb+pVrPJKGOyGaG8K+XcrfnP0Oe3s+rm+jpHUgarP
CccBQlfKzDo2YjT3M0V7j3XxwtTsz9aq6ge5AaTQkl/QZh8ZCon3Zup/ww79mTb5
QOCTqRMWIayL0bhtJG4UzfOGRDjKblRKLKkydQK/5n8kHOaRokzUi6N/Ag+QNmf3
cZoRz06tLxdwHlf/RYYVDiS6LDNHaW0uHSzMGVAcZb/DpK5oqq2sXlXOcDOK6HvP
TSTf5/08WpsW8NdyPp3fXhj60G15MA1B5wyQcd2RDJ2lNSZon/Ib1S1TPVGzqHkQ
dal42DLOFRFc6vldsLT+DQlfpFbQZi71/iMuAIXRJTJYFKjMP/Pk9iCsF5kJkCKk
`protect END_PROTECTED
