`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IJq9zPIq3iIqF/p0X3Fv8X9v1sIa3y3Gnhc1FBIzl/Dfi6/5QUfXATVppAY7CaR6
VsF2+MDNESIea+d3epjgnhFQoBQu2ROdT94caL2GAX77GamUgRH3Kw/eR51+Rbil
9VTaDqCIVTFlW2QBnkWEUzQ3SDAxThumXaApyd08EexdU/GnYXU++BESPldk6mEE
8jiLMM98BT3xyUFiaKpL2zbX4g3DRd9A3Ud9ZuG7Yv5R+GiYPUMvGmK6m5MB2iKW
kQCjCS89b45gphMiOXPfdg6t//ExzvIdvRPrqzWYx8YyJL4mmMLrr9OzW5wi6n+4
0H9kVtWGgtyo0Z2wvpyIY+w/CTDG9YGWo2SZ/MfyK9o7cBZpmG46oj0IUFIUj7T5
6BVeZZv8PBfewi2omcLABk8QBd9Pt4WAsvJO0+QVitePGr29Ubaa+sC25xmOuIT1
TTffOsqecFQewrgxfA1OF6pWCEk0hXrKh66DQH8XJbiA73qX7CXIbYM5u/LIZA95
FHRNJg7ADJxylYoBdRffltA0RSfKFM5JX2Nlv+NZYssvTx8d3lh2waiBIjC8nSVe
/HtjIniuzXeB7JK2cy9vc/ue1UeLAPwaL63a+ccmTCxnmGFtYzTUK9T77xVuq56K
26kDRCtQR7rzp8SsZkDvdThFUj4JzXS9xmNoas/lpVnYp/xiYdAMXSrWu0qV9UJe
k1Z6JzfeSVVW3TllGtROBAyrLLXu13FxyyZJuheT6EsGTqCBdbD9DOIrI0tYKX29
EGutNZmGnlJbiVWRWTLNpa3ieWbtzEWhCcktODt8oJ0SuwGeNH+W3bhxEYIHhqKG
i5NZtYCW+QScHnBlfUbRb+LFAStwdUDZEEZTQDprD/B8uzeUuNSLXWHesuW6e2Tg
6NkXiblEcaXphMcFTMHFac1Y3ufOMuV62/XO55tkWB2gKQrCHyGIZgnHxKkd2XrX
+l1jhnWfLzcalUqEWAdBLiI5LcN9iyKX9hmVIagQkom6+emZrMomDl94PuZb29d0
fO/IM+yIp5XPVbC0cOj9ZUbPJLhb34RNsSE11eQ6G5ve5W6DoOuHwemZ0dOTo0hg
rlQQETqVpIXokz2Yz6yaF58dzShX7MWlPcoa6+dkv5iu6QUaa3KX7Rdd50vWcpge
Jcipgn1+Ac30sQrW2fi+9POrbrQ/cov77315l9xrJvQRnwCf7dmvNxCrIH/DUUuU
bqBJEiD8G/Bw3s5NrPcugfsJq8/RNqbN0eJjvxkfa31Uj2sCsqssL/jbUrb47at9
5z5qvxCOWnQQKbQ7FB/BSjwFjQFPs+b/zc5tlE59yqOfBUN02Py8GaGU+CTrbPbS
V5VneOdJlLFYBtnbOWjRggFOnLWjf48pjTwU1CiLsHQbMRBiPVzGtfO6QOaRB4zD
ZwsjaGIujCV8Ek+DqhNuo2s90qAsLjJ3kpyCsVFbPYBBm04U9x97RBU9jzGBefZC
fsILyhCGSgf4EpjFNEFpCT4YmsVj96rm6An9vld4qAXfoHOlbe3LNWn9d/nVuw8+
A8CiGZNhMhopzOiko8dEFhb+cQQxXCS3/O0xlbjvKFh9judaqEbKvG18e53AFdW6
+SNoHQjT32qQRgZAvijDSUU3D8Rmqy6UsX9A7gFq1ilOaiyXDmgnjcRKmHq8HPnT
WSV4lh3z4FiGSpmRzzd6vABnBFxh9Q243yUG7IISh5UnUFY+JENnEH7CFJJft8tG
iCgu8zKaeG7xfDUPzq0JOb5trliamN/gV0LD0+5UKBRjOUxrGBmjsbHcfIZL0Jwk
J/5V52v6NIysl9nRtqbuqNXFBFsM0qnRGQzMVkfOE0CvjHE3e4e8ecR9hztzNenl
zkNdPqDBw9/RUPKUqT/ObUywQe/X5pRZL34hBYURx6lLVtmtON7gX8Rln+aUJAI5
BDlSlRLgBvhhISeaTgFPr/kCNjcvwFSU9xoerbkcf008OxwsBnRpsXgbd6JzA5/1
uhLTiBUnTqBW4mQYIBXwrEhoS2dDKSj5rc1wlfvH7uDo+NzyoidUOzv6cuagCYJf
jVK0QqTOPLhCVs/i2eF/+xxvfmHYo7r4HF494u1H3E4vRWRporoJ0+kUVLDjiuT2
ZJ2U5lLCl1M+4727wKDdXUS248GrudQ95RANfgLBtCJL2mR0DemNmu/eYUrRCfHT
eigMOQ+yZfd5A/2A8y/CS/N/vF1OEZn19NFHLPT/iSVfu3p8tuqEHpfR5/qpiY7F
A1S9dWnZ6+f8f/yg8OiM5jOxHQtsJPXhhYVdnaDuK2miEQ4UTGgrDWqN7qG+E2n6
t5q8uhjCC2pBMmWQrLVOn1U0I4/J1Eyvovi6w4R54U3EY/MisLG1SZaNI/D65022
Gr1YcyNyxp4CRuh642q54mrlHEm88UAiU4xxo/W78B/Ehx5/Z/wrH9uquXLCdZSo
+eEGm0a5dS5ksPbbuMdWKgPqtbcmWvgHiNHR9LcdfjqbNBjv3X7HJw1hEpy3/xJ2
GhXKPWzLJkVTU8aN2EIEETKWV+IiqkvNRNEB+zIJP0HvKrRXZDbQXxaxN0mYiHAl
f+LuSgyBRh/pJjGC8jL/W/C85ZsByV4SvExQEyxCREfRcvL1OM1rNA7+5eC+WGlN
+U3YPkwatkq0uq0FyhbqRMdST7cKo+6+pc7DNK2gjb41orss+IR6xVGGUf8h3nE2
JEww78m++7a50fGij/1WGuqd1z+SPZ8YbvBoH+FLv5msfnThE9dWYKKXktjBBgiS
B+qqVyYtauzVsoTxHp/xgAaqaXJrhIArvPdleYMg18gCoPEz+5yzsYs6bV9DRlWk
wOdJGyS6IQWVXfDEF+PdVQmDVNoFOMm73suYsG1nN779E4J9N3rtQkS510/HkaCb
+xAKUF+RQMqkNdEd8tYnTxK+UYNW0P50zdBcW8Ev/1bsP0Zdv3b69U9gfiGZv24d
5qcdjslhSf+gjKn6SGrcXc9EKFipRAXRkq2d89HKlKd57kJyIxiqijJpAzvK5LAY
/DyZVA4Wcyg5L2s7qu4ky56fGL3NfV3zNDTsvjYDkfgcDQ8dAHlw6BQayTIPEs0f
`protect END_PROTECTED
