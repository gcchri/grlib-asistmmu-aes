`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0RbkdAjbkDamxE+dt1vwjVy1eDZc4lvDWUwzpNBlEi0xJ76NFIsJv2Xm1vHCkhFh
vPft+e0luhOdfjHWwXAQSPcMYnrC2l+YVq2YYJzFL+r0Jvpu22cg6aeaBV390hdI
7trhg534YrIkh0KdrP+ZO6F/Ooqgrlz3YkpuZ6h+V6F/4zrzZZxAgqFBugjrzbE1
moADmwJUE6xONERkthft5T8sVGf2N7tyUJmC2WWdBwsUYschRQ+bHroUePpVsMso
huxASRaQnW84zqJI39kw42lr4Zf2GH8OJU4UY9Gs38qM1HjECDviI8CMYlviDjXp
ksJmJ5fMCs5VitPOqvfNd3vJ/H6L73+ufqd9b7divN5fwnxLtN+85+k5GfYffV1P
ZMOYwZQR0yOwCgDbqH1o9KJ3pFEGQkw7bzkux6WfJRdJ2Dn5udL8QTDLoDvDYFYU
oDG7d8/pq68UABjdQvDTqfzSppjEQvMgGOoFvOGJNejU0tuQW+G8R2mxDw3Sx+5b
EKXpAiWnv5086FwocU6kdpnT9C3KuX9UE1b2VNADblcYnDCW1fc0dL94BKG6qAEM
5snMAKkI82jgeSaBesEc9R/mkQsm3irj4cHJsG5VtmR3L/ILE8kliZmBIKqiB2u2
KxU8uy6gUIftZCidDBMPVLInHWHeolrH56D6YFnIOkVkA0aXfwTxvTd5rsyTH/f6
ei5Lrp9HY9OvtBqYuBYkGyCQoqSC8BfniWimjJXdziGZJNMroRqPbRndY3nfzwMK
t8UEZgRqZu1tdQabRK3wIhC53PUI1ks+K3bC5azalmWOb/cx52vZL/uVuBCjOXc+
6Sf+hexCBHAqzdC/mcfHGevXHDa1LmmnzCzPAsvmOF93GixupBMyN6TJa4TOeRFq
`protect END_PROTECTED
