`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FiDC2JPrP3NmCnE8OL471TiRq5bP3ys1O3xr0sXf4FZaCy0UPTxb3TVSpcmEDJYX
X2BpVIWCnm877mUd34orGjF/jr3G0EtgAYC3Y8tezpoLRx7Adq3+BxzNyDqAhgE/
NxxLsRTLERBDjzAelMUHyH/sfWajsYDZoO64th2JkOhk5C/K4Jd/uU59zUv9sUqu
ASpkUKURdg0uPqVRTCgLl06/tQlIuBcPID6Hwa7EtYbNwqR2LNvnzdLJfzwUnard
vKInlTSGczhTmG6KdHPsf4ikdysg4KITmP9NjR2rpFMFAe8C1yM/tVPBxlWtHOJy
qBP+iAiHJwQwNJ9zyGPpDBLiqDabzGDkcC7c467syjvQ7aW+tZrgnwsn27EPDCnX
NCTavavM4Cf7qiAkOH/nfo2CBxYSxSVT+8IgrUg15Z0=
`protect END_PROTECTED
