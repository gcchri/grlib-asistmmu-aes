`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FTh8RGOtgpIXOYaCymeg+vu7zuXVkxJDKKBhtD7eX1kFnleDDG77rDSb3ECL5Y/I
X2oImT/J1S5dj1hc9jJDETsyQCkD3jVcr6Y/MEEABvzj46GFXg0GF8y8Zh04HmuE
KJcwbcaH4z8Q61bx6m0BGuGb0WN8c0mMbj9I9VJB9AtrraEn6ch5fW6NX90r1iYx
2a8cXp8STvjkACNFGnjcUB7nk+4RDcS5X/FqKxmEpFFw172xKD7g7ohVpHhKRVES
5Uobww3ihObUvmiTXJXCrJEJxTKxX8XkNV6LvJ6QD9OcZZ4z2EfnNpaVHiQfZF7l
iZXzP/eWVVjCjBbRXGy8P9PYAn+6cmuOqDruU8NYEtAYOOG4hUVsijIMfABQPWql
hO88zt33bjZmJXKb0DhygmkSPslN5odfHavfTWlZ5dA=
`protect END_PROTECTED
