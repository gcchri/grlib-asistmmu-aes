`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zWJcRi2Wt7TfVlNi3zw0j6pPmqnOOSv/9XW6KHed9w9+Ahd4PlYC+fEupumaAZS4
zqChx0ePF7ktVC68b9wY6obtVlm5rfkHPDoAUvyZHOoQ1sPoYwz6ue1U7j/mWpal
ELMeCqRP962KDbYqguOvDUI+YJWnF/jNfUBiYOxjGvdMkdoEOxlyBkcJeEoF+APJ
ZEAb8R5059Hg158LoxW9MP/OkKmkrOuFxxl3HywmnhwPAn7sa8ttHrG9uhCAyhLf
CkYyrJjuik7aqNHbVvg6D6kTVBhY9xqHPrL8u+mzwJX1pQDwDsgE2pBQ0K9jH96e
Ql24MFRbR0Ivu1h5d9usXE7EgltaL6f6Rui0c/MW5ZaCdnkmo5RcS+jG+LElIQZI
vn9CasA/m7uZF4iQUKV0lQlhtkOfkwz9E7iAiWxVaKI5iZ1SDJJozjxh98NxNTl4
XALYkZTr9ezc30vaXC5LlNN5K9TmhYJWNqtqwwnPGql/aUW3ywUWc5REV6CcdHjl
RWybfQWgF35d9o6v0xftAa0iis37qYDRguBvbsEbb1rsRHjfcIG+IHd20fBcXiFw
wqGUIrn/sAVs5SXpD3GNPQYu66JBhp70UXbVroAWu5nxn0i7BtIgOMYRviYe0L0x
LVem+WAeq3ppQgyJyT7AwDOyhrn9S31m6JM6EuyCJsu7oQUoZ89vmBbrHbq29VRL
nax6rPGhcy2IobKq5Fm0jWIStH26FSjjwr334YiBbqZRQDHdvF+6FSaOqp9KOWKW
iff4JONDBQmza7hJBAtQD9Cs4EIaJFd2qlv7n+o/VwRwl7Oil8c2x90GF5n2KeOw
7qbAwGZFyWRq8sRz7WtKB99KfF2j77ea3GH/BXfU80V04IPNrwEfv41jkJlMF4dq
zTHR49Yhd/adycOdF9TTAp8V5z51x/QGMZTqW6Nv9A4uGPVi+wxBd8Z5Y2U0LJWs
15lhjth2nhtvPHBPpIaEXODYBbo1LmQVIP74RYQAxTk9i7/GNo9aFLKaRNK0ou9x
5Xoli7CvoGnF3RixYfFgVNIAfB5hZzEMRimQxSvaFuL5dKcLFGMieh5Tugj48Gqx
eBodAwBCWIJ9Nq+NjisL1GVBgEjgkFp6HlRLI2cr37T5hkRUCP0XhqgQgdd7r3db
CIctsSNiZ8AiE5x1PxM7KEHXbknjlu8iPI4Ybe3DVs7TgSLgllfdIX8Q/c1G3nbq
xEuZzypxg1aimMS6lzvAQWTX9/4ujyTE8YHdpsbd/D28b6unEvSMfX+syg/oBv7M
bthkKsRlWMkCQY6IzGvryIxDpgx8UvFmXfzWA78/CUzgD/oE0M80xkNd10Z5Z4WG
wiCZJzPIuLPQRsYC74yU0tsT+pYArSqCkUSa4mHCBlz2Qfw8I+/1b9Z15V/Of42L
`protect END_PROTECTED
