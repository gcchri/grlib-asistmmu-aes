`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jFkS2vxQCvuTsnX2NcBkfanl46jTaR/bl9XDL4o1Zv8oK36uQ6JgP0Dyi8K6XsA+
KkA5oouy+pWfK/w7rQz5tBmVi1hsJGt7CE17e2cBSdjc45LIS6SNN4d6Qq2VQdxO
axe7ni2uKjKEde/jCeHW17GOIulwZD7jCrhtkT4mW25ZpW7CRULxg/tXY2h7de3P
pUE/idK4cuqwa/5hwhsqcPITAmj/Cmov0Dmhkn+FcfAGCzpXaRG/z5zhKu/Soq17
rnRmbzRZeBH8hmAsIxTx8OkVQamoe4pVzgOV/jCgpxsl2kcUZo6kxUeMnNKpHdZN
nFu32b2jTBq1UZ4egpxUzvWuYgLzvanql4tWWuCUdZ7u9cIkop95cm2AH92hejoA
OkRKvcZiLhx31vIP8SsL07r3RTmOSy6Cq1kjcTRQCge59DfgLyZG3KYEmVti196P
FCNUK0sWpzyuQWlyVYjkDRwOgLr/8kFw0A1tFZUwoM4LLnToeMuFfAL4rlmVpyiV
+9htZ5op2ggleQa4x7nBUULiaR27cgLx8r2W1e5BHKlL/bsIk6hUUcFtil1re2y0
8pxZ+c4Yv6GSAf+fO2wk6+MKSl4lbRdqoxlqno4dLBCMZEwT5PGiT5fYT5JcrlbH
jcAPiu/Oc4b5H6Cj2B0PdH2YWIoowVyZNjfjdY2kSAq+Fbf2bs6SDDwjvoaeED3s
iuzFv0MV/8lfDQLAsUNDlLvyl5aCvZTWLGDSrod12UwwgzJ2t2Li6PQBxJs2LIdI
kX5ofu3/3xVOx+lJSqjGaPkGpzKYQEGNItFH+PgBZxDnplYkp+Cu3nXRg8VdF+sh
EQydI8guiRHn1WiTQrpYaSABv4ro8keyQVjow2WWZP12SQqOPb+e/yT1vMfsXC5w
W5n0+nTKCtkPnqA3NrjHkE9WaR+vpn8gG4pxP+ntwfGh1niimcZcPTbkT3oq/Wd/
ptO9txzZHrd4huISLM33b+FQB+5GMxcCx2QndPKnLqscmat5mJS3sRUbzq8zGRdo
nPvXUTByMMnUTEYqBJkX7RETO0ajZ3fQDjLPIZvwPcLPr6XQM9QbUzqABgQFCAzv
M5hkRcytJR53xnYQ9UBNhl1O3vLxOJQnR8AejfMct1nmQotFfMaBCQjvDcJ5sTfc
`protect END_PROTECTED
