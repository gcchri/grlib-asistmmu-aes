`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n5kdi2ObGBfRF8IKdYz2a5VRhwQoTWxu4oy0c1wBdtbR/Arfn3vY4QW02/vfFgDq
7kV+ppm3VcUr9MIT0C18TPfLH2Kh/s9KPJ0JqsXOESTAm8Ig81I7brX2Txwd1eTY
Mm+4K+65cViELhw2aQXPjyz39MjaEDfc2FW/YrIzWxKaR67T+OWyjgZcpa1BDQrf
GpsGRG+cynrvMsh0zrwhq3AeLATc3lQNSa+a2hdy6F2wAr4rTNcXOe26VvVEhxFL
R/eIPl97iWiSqK/o9EqW+wDSrEBmB7Ft4rkdA2Z7cNkAUo8ddHJ1unXAYSsoszR2
tc4DdUnrJxrfD2lcwLwTuXe0jD1etZMC/GzESZBuRmnP9XFYTlAxFvvJ8/CgqAIx
CCssM7SizKnlTD49CpELjzaLNH4VSPYfw3XQ+rH7+1/pMzTYTbbKtpwlemUY0V23
nl5GaAQzzNLGHCdjc3g1i5foqImY51eKeZBlAH4g/byqhlr6F9Ez+JI4LpJ+6ZQS
tweGTHHvxcUPDNapz+H65DJpn7zLdL/7UoYxA5EEJpeJO8S8QX+iLBZqniyStnAW
XAp/ZNRQsamZxUow0gQmiHutcaRApbmWF+bZyiOWOEESwJ0SNwiW3LzZ3rEwkeEu
YkU+CSsL3jZPNS4ehaQXDcFr7gM0KOzEnDBZsKKeI44=
`protect END_PROTECTED
