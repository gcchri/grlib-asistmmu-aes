`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B5F/6aZQMj6An0rYd7hHFVEOlrQqkeTPIxtzlpzzaem4++lmg44oArMNPyOl44Z9
EhEykMGOc6UbQobDxiUDeScHA3urOmejILPSc3TrN71D8UPQdpf3i1PGGn3QkbB5
NE2S1D+f6lXJztj7OpEQDgYHJbDB2Ua2pRLcDk3L+mbsA16yBaBar7WN3Su/9r5z
RBT+6ZUjT68WhwsYnFeFn4jWvgcM5K5pP7F9L2glL2Y+nnVAkhSCMKIAB2hqs9r7
ucauKV07aZASrS4S+tSaxWSWG/EhwNzajKTU0U1lLbzCidd4zPijxrDc3CKhDnGU
VcsXEUaegEE/joGY4zP6eVjrqWphRszebUQjcb/HzQNblxjqzqW6g7FTj2Q42jII
tnOxb7clECplNeAoscJDObWrWB1UF1NaOervMPKty1+2Yl7FHBFbvVugvQeeLc5t
VlNfPkHclzuLGFmoBEeyMvc7PJi/50oXYvvkZlUXZvT2r52C8VTcEvGT+zPKuCEq
heI4O6OLtsYpVkogS66tvduPqh5bi3xF6bDyx88Ge+j/Pva4+nkxAhQM2AJp0SPL
H5uHWbt1e7ue4+7SIlPlzWpyEsgNiLmRCewKPKIbzg3vpLE0vHteWKtTP9x3++tW
AEaNvZ+c2rnX91B1oWrSNvsfYZJdcWt1OfxQ7BSukDml0wm2uTDTKFSeZ6E1Fn3G
+sshNovGmRhi3dteCRJ7qvZnerqyid/s4y20a+tx81HLTk+zdH0OilJ0EkowJCLk
ThozZO8QwexJ96nuJLNo7+bKjUPp9rU6qdT3Kmw1vJmMKpUhVPmAJn8wWbVxr4Yp
+tZjaFhaCYAjgBi6xt/Q24xr7Ul2bTYTsFuGHD0VnN1/GFvw4CVtVr7xks1H5HCC
IZKRhJ5Ut158N4le88X0BKL9qQ9Fuw71bcCGBBVoGJqfsFJ7meUzlzLIcA8Dx8bU
h4qIYPk9lkDqg+xZHZ7w403T2V2LERApwrDj7t/1mUZ5d0ewD8OnATjGFva4ryDt
6d1hSARX6BpTvZ6roAhqqNmNd+DfkUZ2ec5y45PSQ+2er8bA7U9oI7d2ZQ9OqrJ2
QOAOxNIqaXsTV1EX8ZGhhcNr29C9EhWxTzQXeZUoSR9aH90efNTOb63qYZ1MYuC2
CWmnbJzPX6VG2Z7cITrvDPqHmxSDFyodT1glFuk2Mo1JJHTZTW1TnpjmoD4p0qXr
vYlyujrXe7XD5PEDEbIasFvNptnm+crtNHr/WBZ+EYSOAhgaIxok5TQ3zsXUywtp
O9DKjr6YJvAfhcpGIlnwcXqL8YX2sACZD1iVTwqzMDsa1M6RPpKxZE42DVGaHhHw
`protect END_PROTECTED
