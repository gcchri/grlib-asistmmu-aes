`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pWjofaeHqA5ygecItoCR+e1vMxAYS7CmIjSnKzEnL8wmRErwbJSq7Wvc+pw2srWn
IEL64bKqCHKoty4M5msrjN/taJKeDEtbaToLR2W4g0+PCO7XWbabO6m4W9u/8OFc
QXR6jrfwyp500O8mXfqlmTxJHXmOvcxEPBVRPlWjxj+8yT8vclETw36MLdZcPsjq
i/UWYCEFU38Cttppyr1w9jE47MMDZ4/T7ApfU2YajpaJMGM/oH3V69pKHH2H2huV
`protect END_PROTECTED
