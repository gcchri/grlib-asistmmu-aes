`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wYl+/FZaUEmweobI8wYMsZWuTWpv0lthypsVO3AdTDVmgZ+3U1oQUqWhph9ZrvOq
Ko3+EvmEBS6gUZCKWZkyMX7OmBghwV/FaCpykgmcHOPALS6sz+4jgPyNpsixfLEV
Y9HpkgYOpHRnd8X+f3jblIyOA1V/4/QfsPCfydXd73OeaHiDsIzNLbSTHYXAKPHv
Hu6sDHUM1z0q73045MFcxLtfSq6bPBXPPuN4MJZOeH4CWb84r4hiRHct7qIOdPyc
c7g45SNEK6rMwYmz961/fc+wfPSeJmk+dXawlpki0QHl3x2IfswokXzJFbGjHqVq
L4F/U8FaCMsam4iM0rPHe06QHSwJ+Bs9Nd5pCnBhBD3ygguz1JC6u6TthQ3bOEXa
HYNui+Er4mICtEr/EaTT9+65nIP1p0vqNiJ2nv/bXDbsSgf6LJ7QRrZ7/Ml91MmX
UJNiNKqpc5Ivc8N9qJ2jyUP73YwY0ZD31WjOIXrrbxxD4dWUw+bNNI9870eE0I2L
3O/OeMGUoxz/rKdXxQWpWACWQUCrBGclC3mkbjKtP5/RFJ7n4wEmg0rbVs5d6JgD
lB1l6AN/C5TAw6diPaT+jtJoVhyu+BH/7zViHsPJ76xSKSEkgzPbzJe8G9Ia+Ked
T254iMuGb3c3nC7K4Ur1VcZwCXZPvzMU86v+i0nV+k5Wl4ADXQQ1kuGEAylMdA7D
FxteZ40CN30QI3qIlwlX9by4Tod+koR1vJrmNdQLSyhJovtih2ZkMTZTjYlTh4IO
9EgNAQ7mhvE8EgdYi3KzbQ==
`protect END_PROTECTED
