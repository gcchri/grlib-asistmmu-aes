`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TYVUJFx1w8RaRf9MaFcCgkp74QqqGIAXU1I4hCO14IcdOw/h37Z5Wa50BCwUErpo
Z0j1UPaSccOUwc2shSJ+HtrClBCBv8LPQhGhaGCFjULcpDczdo8hCOjbLNYx6YkI
TPU8wjPoJhNiUH50edGDrgMoHEsM5BvihJFB/fop1KVQ3aRTGupV7D0Y9byL/u3A
jKjCTc8Le/remqY0daN+mAvBec2iEEVkgFhc7f30LtIKdWh5yEkuKuWEFMJHq2SL
qlNX2hi6wll6en0JtfP/uqwYkyx1y2BSVVsH2kfYvLLhZSIXWMeQtz517Xot2D3O
mlCjmvAnSJ1fnvDUUr3e12ruuZrhkN+mJWyp7A+OZsMFp3SBQcF/fgsk5JxuscJ4
hVXmXRjwfxGgEEsxq+ftvcZ5cm5vVeuRyoOMlsRxm8tgf4hHSIKoZ8TancLi3BMX
`protect END_PROTECTED
