`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hQYntjPOIcJkXGuarGDo/FsbSEtGDt/UoyEkjNnKSvaZSsSpziHnzOvZS1j7N9RJ
xf3o1wamHcwG6SgpVUIpiCwIv7+J1wAPFWTZaE/YcmqXiv2OyQVcDvAg07svMC+E
sc7sNP1CgitaSkHLJit21wRX+dps63G7IfW+7NcQDw0ooWffNHvGQ6AdS0MI/ktu
67icE/w0POmQIYR7Zo4nng+ofu63geecaHhtjY4GkKg9oYcTjMfZFzousaWsjnWq
AlL2MeH+Q5nwqwRRXdLeHZssgOMmK4e5Z/9rBKtvl39WHblAfY5LnCYfYEieQglP
p9FUul8szvI1oP68+CZ+/oqwiOcSHOEBLVhB+aZQfBC1HQrEWVbEeIwzn9gwAv9P
gJphGIQM33V2jgWP7SU1qBkGvH6NH7elXj/2PfxIYat6IiJagd6FqCABRJpyEbfs
JP0qDIY91O6IXhqdUu5trtxK+EwEYzlHkjaLFzdQzrZkmDJZnF2BbF+uwXtFDur0
nqrSmfqtkDAsnXYB+hf5OG8ChEwkl9d4hJy9nJJfjnI=
`protect END_PROTECTED
