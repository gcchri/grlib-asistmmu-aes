`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v3iOqpoydeu7xWNKwM2q2nXt008Tz7zG/lHQAiPc7GMz7EXS0A0iHIogvGPQH96M
q3R72+uNhbQaQU9bqFISAHWJ0ZFXTrOmmZiElov9Z4jL7kuqTn2+MJdCgCsp4nh5
CHGQyBQVX0x9JmVIONll134OC1cQSs2GNcJpsV7n4U/6jZWvbgYChrX0+36QYAsb
NWe4RruNzVtmK0Y8WsWka8rfNo4bf/1waxdypEK6H3ysRLBCGAtYGFvYg/U+AKsv
azM4DaKUOi7i0Nl7ap0/74o18+jEUE8NhhuzOhTo7QhB8Y0ZHZgxWPS29qNHP1zA
+pcX+mhn0/T3ZdTCexDtDQPFmcNN5NPjqnyjLvhbgcznoW0CxFakf4I/AT2kRhOS
i9wE2IlqKqaulqqD+Ynseeb8+M+94WI6WFd1UHSvCQaDiDY1rG68/cvOIruwX6du
NvEzEeIogcoT9T859Pzs2qxfe+sZJaAEQ4g+ygz2T+h95utJXQ3zUrcR45GQkT2W
lAVZEMZa43+c7PHGtqy9cBKGYakJFae1+Ynjj63WSwxnQ/GgsXDrEs5B3uaTonBm
l++0cmJvD+pL6YTXTOeJuRWSRc3fbozvHi/2DX9WIm2UyF2AyZHnM4jBj2r1LRL9
Tna+MlGJvLN4ppTHA6lnzW57aCTwthaP/+kirHctJXs=
`protect END_PROTECTED
