`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DgOxHeLjA72o1CiBpQSsPvlzIzKreRGR9yS1+C7ACYmx6ruR4mmymMkyDJn9CtAV
NlhYaV00bxNuT9adDXLFGClxNYEFIWYmnWGY6g4+/e97inj2dsf5I3sUULMCH16n
CoJRg/i8qdEEZR6km9ANguZcXkUZ8u/q3bA9Sdzwb/cAxO9BtS0/reu3JmPUeMvM
UpC8IL10jKIK/rjcLrVFq0WFtfmYnfseZcTOxpG9TzpJE5MqCq4bFVC+zkacQXu6
8kpOybKggizGXKkn/zQSnhlvUCpsEbfLGsrUZHc4LG1hQGD0uGoG4sHUFpOvY7mJ
khtEbrFg0HtYA9N4gszcdx4yO6kytlNjDZL2LXZzwnmWslb2hmQvWZEIGguDwuqg
BSGN/LQ59huQ1VNIvpaI70Wd9dJnUNWLGYtnzth1QmXoxyGQL4IbewOl/yC8mDh3
T9DE3M2mJZDWhf7U2phmOkOhDFoUCTFqApm2moWgaio8Euuhq7KTGSucTTi2X6tJ
7kfEY/JUK0Br0Kb//abL8f9lwaFxifcPaH6B8JbkEWL+MJdaULyy5WXBbfEqKj5P
njVGEKZ8GTuM9RJ9KUqq0d9Jwg9WDBvMD8q0dKY1sgA8Lm7TfRW2DA1Dzz9kbM+w
c+uTidkPFxzqi1U+XyzJqA==
`protect END_PROTECTED
