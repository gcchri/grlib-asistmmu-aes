`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lKkOuujP7cfwxmyshOSWJo9lO7s+O0V+7oJg0rggh5PMe3CsU8nYwrTMP/aIKQQh
kjVcrui/I9LAPuFnvhUcYNjihX2jbBV88Bc5KT05fVLFycaJaL2GzjclOZdrlUah
wSYZ302B9Bpn0S5NMELTIURMlTQsJgPe8n2hwrgm4tw3Glz9q87ZZCooTXya/nOS
oRQNVfMz72y395cTYVa4b3FoEgTQqBevcO4eoiwn/T0aN/hrAKK8Dq6/Co4LZXRu
/wJubUw+G7G56YMgG04znhTJ3dVgCqy4OY+ZOUSrwhrnyzipGHmMyDv3qFdqRDUk
XPYOHyKRAS9ewO7daiGH5Uo1ZL8JWclRzbhmTnc+0wWvXd2qFbAn9wfZjZmpC/f2
7tZh7M+YDlEOIdxEtTmP274R2GhjJynGMoU0ZvEbLBWwGSyW7XOPZa59ApfqSBlL
aAFNEGizie51OLsNkAoIIkOZGy/MWlJHGl8itVzMOTg=
`protect END_PROTECTED
