`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
neHxWdC+ddYj03HShs14ATHfE/Ur7HMC0y679jJiqccYk6wbtOyDM/pJdQiDCdlw
J1H2j8XeRAC+W0ngl7tF5cDToFFcQbc4+V0BibODhpUhwK6MbXY9uZqVh+8wtDqt
p+eCO3TS7FLBpQSbJ+OSEz7TXj160HXp2b0MrbNKnjNEGWf3xet7lPF8HTya9qOd
c6o/Z8ARRKca7G05QyRqKPfo4KMAdgPwF6ROJX5b93c=
`protect END_PROTECTED
