`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SwcOeCyP0IDHAYSZtSVZ/048KJXse+aCwEC0ctPLw2b8PYZmDFfQvpginIuC+aMI
QKNiNPLnzCzfhUEEm0Kd1Lnm6yZfsfSVz1LZdwCU8WvW8utAi+ERdvIVZZ0/7THS
kSqqsnKfTmaO8Z1TalAT3zfDfpnBdgcnvV6aNfsHt71Bt8Q7KWRcweFpRl2ebGLJ
OZsDezdehEco73n3Xfu9LsFq874Z+VTqimVyZD1+rDWkWQzDlXDrpXdEGPRpQCLu
rIzvQu9MGBmbyIxdOr/0y/7EoEmZCldme7hnOD8ANgY1uPYsWtj8MxK3fQiBgIKq
Cd1BqnnlGiXkbdDNujFWBzr+TjsqF0xw9F67vhgiv5GsinrRJ1gT9+pMzPcbOty1
bquwsAtGF9+crEOdVb+/JC6foW35f9izANh4AhFCzhr5mt72yw2FiPLGmS8wXv8g
vHyH6K5zbT/cJD13Zrec+wX+Vbq3f7Jdk8dLbIMP06tWzgP7jc5Ae9D6pz3/OkC4
5oNDM+/ujdtbWH4m3uLdqteftYn+8jzBTzu//RQbaF3w7aab3QeKAcZENUaFDksj
bsH07fhNU7E+kmmyjg95ka+Xz984nPhEk7PDIuzXX1up5RhTAvONO4z/Ob/lBY3j
mAnFFPxO/ZHqqzxUriTBMBNodVwhfXWUeHvfzio8wi99EniFUbUX+LnBt+IOEtun
R0o0gWDhv0sVjvZ+F5dB5zNUzrutGfHUwagfqMqJasg=
`protect END_PROTECTED
