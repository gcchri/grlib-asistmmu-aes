`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZcuYKmWB85InkUn88UFv3eeAmrk/SrgURbzeYhsrF+tXyTts+BbVKp95h2W7IsCu
XaK2DCNbT+SPWIRH5tHBrrvU/ixp0cu7Gent13BLxW3SQ4rXqP/M1ZYKdQFuJlmO
UsIqAxc+X4qXijoAMcKZ8LhzGlDqLjCiJHy7ZGdTTbarGoYNfLtXCe16ITVPyCgb
gnfearjYw2k0+WhBOelSWhRckHzllnM6t7UaLf9n6UgW/bBfO65/rtLMvKzSeV8X
TUlstKgiVyrDTysh9XtI4AzosRBnzBa0WskvBMhww6JHASwroM8bVe2rV8yW9FaO
dmCpMA6wV6Kssx3JgYtUOxkZh42DWErl/NqPwcXIT8Y3c50IOrnLtz9z+7PZq1P8
dCLIIz/QkOkgUaBW29Wby/QaOuW10PUqaswsVNmq5yyIs+F/WEEjPiQtfHR7e7NV
n9/2lSKha8qmsXWOZxEwnGmKqRXNVtBACoYuIprW5GxyAFwPDCfo9lfUJGRv3D15
08qC1+s53JKvnixkJxYatC2tu9zyacvpdq7nPamDXiS6tB2YC0i1QwPORQykpbsE
WV8amSwnHvssBwZKG1+N/7X2/734UImoIUJRAXDkneUZE4vZlPM8/ZXkRli65OyI
1XANJeQ/uS5ibZRxmf3iJQYEPTXsA+TsT6rpTFvimNfEgQ4ZuoW8IIsfTtdZiykq
FQt6CD8avwNVNFdaa0OXtfhkQJMHZJq7Ya62E11uLUo6eIT4r+ru3MJWpaZnvIRF
jtfHes1zBt+rleZXleoPUpRXxtqLq6lOI7W2D1YIMvzFu7QKuac9cs9DnG5RI+hP
FfAtHljFQzKQlzLCtz2T9Pf/2o3cT3bcL+6kLsvvYE2H+W8RztpykU90jTHY9/PV
tbqBCL7FC79lc/9/oaiSiwng7VaTPDlbigiZLci7r6q3TjFXiJHSyrxef7tmUMaF
0w5is18vPqchr1E/ketZTZdrT5yQ6UN5Xs+FRE1VMfEZtVWYjJc3sqD4O94+ODOm
2oAWDrqgJcjYy68BRsEBmG5qQSgG0Px7MQG3lISor7HnHVIkn21k0oFmfwchEBj1
Z2W2uq9nmp7AnJH1Bdommg8j5RNiHK3dwSjIrpyAXSUaMqxZBEgOSu35iyvGdPgk
aJH+zMMZiYZVvd3ERbq08ncp0mMSScdldJlHL+gYIksK1kQQ52jaoi1DUYtiRBbD
zKdHKhslhIpGImf6DgcwTTXlZ6zFoTLusrbpdditBkO3EeLLN4PYKgjXcV+0VIN/
gUtMakZvfh9ElntnWJMERmHWQMuWnIjrYXyT+lPG01/rHUcOPM0aj1QhVRQBuOEK
KcammA776rAPDP2edvNG86cf7V/Ilbd61q7lfZzj+TgDTS8xXLwv4R8/VtgdlrqG
bK55xt5u0rJ8/pKKEFay3MiRz5OT/vPZBGiCKaDx4XgMB6B92ZoQQgwllWNncttc
kTwWy+7+Axn7b0lHGZhfMJpTlapG0nSSa2SAsie/Ux11G1AsprXXJCDLPJe2Wdg5
cIGbP2iEVfv9Jtkz8rCxs9WUM+UGkcRv9hfeWQCPKUGNgFfyAdR4tWyn3QCrV1HT
d3aNL1yCeiGaSNiCxtNnYHrss36FiudVU8HEBQ8BxwUpANDbrwBsTdSExF352+mv
6cqqv5CXEvWvEFu0DNPnPbUByLJ3o5xv1NiklYMHrwrAa63Dyym/kQXCa6Bxmr6L
+XWBhPDAkH/dt4wKbBHjrLJBJbEviAq6j9XzRkS56yO9mXi5kr8IiH1tO/8fK090
h/AXhwRfJSmk1dKK9M5hl9Wb9eWjF6d1RN+spWW99CGX8WBnOvk/u0wvHXSTIiTH
SpRyqaA2etD8MqaVJLR7dGCWGaGXQOtKAg/LsMWyffAFZwmI0zmssHE+gaTejNfT
CnBn9HBJLimh4pY/Pm34ltFSZBtPaCQi3aKKu/D9JgFw8e8YdUYZ8Vyu71BgZ03p
ewOZz6Ck3NoHVV52UeT6tl8Rhi5+eaRl/pTzGeymA7vNfVhE3XnfcQu8WlAQ9g0Y
htCsy7ZkUAcS5s0BBv5B0kiZ9lF0+xe5dyDNNveBOE2LR3G28amfVEZNKri5RzKs
EvuLbDhdAU5KX0D+9toneOzDqZC0zXM0j86yAHnDc2w2S/fSqs5fhoVF7WvRKfou
RcD2CH43h8doGgV4XXye5nmHoUbdSbWgZw3yOL+UA+Ty2UiZBdeOeNbF0T9vHYig
rkKIUOPzs/qoVS1ChNvLHOpkLsSkD3BtCRa7st4U0Ekf6VyZ2cHYXL4NVBDczsvg
9ExJhwtQGoxPSfr228ZjAqQaq9TBAQxeNYJNBE5FtItBfjyqRX2gNA+arnM1a1ko
kvSsJoiHHrE5xEjuu4IeBHdqk0rn2QMDKimdpb0W6LeQ/7+t/mLGubXt2gp5egND
9imhCjkflUh9UELo1G3FUnplQsAJkQn7di03lwiBPDnUM7/o78cj3NeD1n6kU4Ef
29bbabIANzn5esU6yPlffC4dvMBKvI8YZDlOHI64Jiq8BUYZpmdgjgPeDq3R9Grx
UT7rsidO+Wrqhs1OeQG4bqbODtxQCkxl5ktN1XEkvusQrQurkwJ6Tjg5iqwrJdqQ
UyIK5VehbIN35Zyp2wgFtf3I7iUG2KQkxQjK8kbn7eCJrjMiU61yQynLDyM3mKSF
hh7DGOFWPNvzFzbAq6hVB1hrmFeXGYCPJxpX/4uo4ZvNiBsPOyjqUIeRwBDKBE6F
nVg9BaSSyvr5zc5f0se0NRkiu/l0/rQvrVG1B3iHibXatttv+txBmybHrGLHyCWG
IJJwLEMlq7N32PGg+7fmwK6tNmRtEyE/a4FIQ7j4GHDyOhbucL1nAZthsNFsiIlG
VUQJCMT9g0kOI8FrOldV1tqAbWKaYqzILhHEmHZ7xh10Zdy1MRiEeZZyPWNOtP9s
pvYoeOk52ZIWPdukAXujLBi2d16I3IOW87SLwyijKFhKH4XcMQFLbfzckDEaM4B9
/cfJQqJDZSz4YPXRDs3XL/T88DP5OvYBSZstIDLqqZ3FE3cTlLC5Efrq5g51rtUG
a1i81IiWrDO8P6POwusmDNE49uIC+ewgGGRs/PMoQlkQNOZ60q/V7tdYk2NhejXz
myX2LW2Mr8E9HYqxq5NM5M3Zdqbl52GVAGbfyNfUoyzzhdHYjRCRfi5DZ/uO/CAF
Dh0guNxzdsq0uyHvClP1eilyrquEnG8ud/NEEkPSHc9VCHdoH0JQ2dawUKdkvcD9
Vcn01uEjIKk68YHjYDMfcL4eAR8nOj+4grlFHK/ySnM=
`protect END_PROTECTED
