`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GmhloNGIRjs8d+li7HI/fYCD9HUTMmpylWmYB3+QYAAfpDtiaSE1Ri3fLlzV/5nR
N7W/YbGdu0+ThMBfpPhjC7VQDtn8hW82P4SQP4SKU5NsGX8jfXV3wxzFyBmnjPfd
UHCrTlAvhhtw76qQ/Kqka02vMC8YEkazPbxckgk/aCd5f+2OWdC3/PnVVzBVVMRX
eNnjbON5fUSV+CfWSsh1fcYCAbfPo/ZoWUJMGSvpciz5WEkdTRTfUEW6V2Q07YCv
RbKE0SkzFyuO7OvfUlrQlDzgC/ugtIXWslBwzxOijj3KKui7Te3kVcUMacZZX3wi
J39S1vDHwtfevMRm4ar1Kt47YIeCDD9mh/fN6u3JxYiaRR7pYHBdY1W+tco925mm
gSTyWRko0abNVCgkmYxE9Qn9s57CoQnDTqto5Aif+dDjVkOv6QJtWWmPT92IkSJ4
RJV1TWtNIHdSv6wT3NfvjieTh2IZSg4lMKiHTvaz1fFpSkAzCUbM34JDbCm76Rnt
/ROAegUsUb0vX84j/NFgXlaxlgT/C1gW6sXDsxmwvlyqs3WZ2pOoGpaBfg+WQrGS
7EyjkID6Fv4h+oFnVvvKp2wh6B5bPYCvkoGL3lCeVpk=
`protect END_PROTECTED
