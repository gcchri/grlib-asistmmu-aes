`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uf/EIEb8gJEvPvWAPEOGqtrBO8riTtUaEKhPE/25wDoGBtPXFU91OBsFnccp4qFC
2HQW+xKf+xtYkWK8ehyJmexUT/D0aPn0b+5YajfH+xmm/7bIRyK5ni48JtvpzfbP
XIE9EoilXRKXl7zLIyH+0t6X3AIXhqMcFw6y8RE1IFnrk5yCD7C9FwFo6RNiF0T+
ZqQv38PS1TnlG6RETaH888m7W/Vkmsm5xred92tNgdRrF1zKUE7r7hL0MJkfI23S
GwO3V5supTHZfhxm3kYIuqhY27HKTuvbkHdF0+mtqdyEA5b91iU22zcoZ/thhMBY
mb1blfKbYP2r58jUdopQLcnQXDkrfsfAfVl6P9Wa9q8Zl7b2tztKJVxVS/FBPiDI
vxgdH5Q+EZNexzF8FrFLa937pWESlqw4A70nS5YGQEnP5i1GaQwYeL+Rno5MvKzt
BjjoRXPWCQ69uMzlRnZiO+xnlLoNYZIEXx9EVxSCt20F3aDW2Daf85vpVdIOwnVl
`protect END_PROTECTED
