`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LpOt6OUvLkCZAfqIFZcUmYKaH88x1emznMSbI/umkTGbfzsWxgGSiAZ4NduplCU6
tu4V6/+GySyEQgb78/Ez+teNew0R++vO5mZMIH4qHT5ClDHCPKn9d3m2lEziGasM
5Sy4sbSfWQw2jvzuBFUQPIjI/D77PsnLySlGqHKORRzMg1ZXrlRTGDJ0oh5+iGgo
igHldJs65soZqPv4QLkai1relFOwPg9xnIRi5TNueZOXT4j8MQ7ZL1wgEj220KP+
Y+wA7Fygnyv8IDDdo16tCGJBKVZQAdUQfm1qvwB0c2YLEpP6uLqxo9datjEAl7mz
44qjQ3I8bsOIj+FTa4J+MtUJ/0olexUryEJs9p7yFJIwL6FUbuxW0WSPECjqWZnB
t9QYj9qoZuAXe7PT6aT9tNQ1bHDp6kO7uvyRWOZG8FkA8WoZIoua59ann99U1sli
1IAVXc6rOT88EAOZh/uwD6kVUDAo5+3fDow/Hp4NL7jN8iB7aAe5n0ooFDtV7byz
l97e/axoXxjoweDKESTwQuwcxyxXoVk3LdyYtjq7MWVVMZhcUFnwE2yV6+P+pPyx
`protect END_PROTECTED
