`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fA0GvUVk8NdapX5w80WYUTNxk9p43rE8xh3VOvjF/vME/AYJ6hWgkEOSNQEYMNYu
r1PCs+EiUfRINVILkzRo1A187vSRNuRw+IlPQgeM/lCdd2scaqsL/rb9DJI80mfU
dIVvDoC9p6bM/t5KsFHuXURPQ1pnTGhdOWnBG+pJL6C5cOeFTMKRjDr6gxd1h9Uo
t2kTW+kY0pXKqgDqGoPQD/woo/s/1KDXYf3q0d0T2uSfQvfgW1oMOQQnxpmzKdBQ
Tq2a4bNH38CTmvV8n0r6fNtZ0Lg9djXsLq5p0aBkpSPsKMnXTNK0eKrBi4ZhdgoZ
JMYmT1ZBNWbIoe77rF9/Hl6WtklR9Y0QezSUzg9TJN5ABKT59OZuRYY3wwWA7UnX
nMdaF+LpHTdxt6Et4YHHf2RLP4O2ScFMe5PAm0vtgmSyWveBZ2NEmAcPL2KtTTC4
TXDXqU8dtMNDiycafstcZ71i/bPiF0/pjhLKMNAs03Bfk8YGrkjTFXPjCZY/qfMg
TrzbL4CnXJOIwLJJGP8gh/zdvwoGgG+P1K84/fKWHfxvwaf/wsqb4IP9VQTEOvkN
5yGIC4MVy7Poji3wIqXvAQCpCUKQNOT0JaL5L2b286zl4wLpsY8Bzu8yR49iq0iy
tUmj4E5rXmVCrOlaGXOHq0nOHrtSS1DGdKje1kXq+3Pkf7wb0hlgycdxTo+6rFhq
Lxw1OEZOeMTHkdxmZzStQys0GlwqrWa8nEmBrN10l1BGT8VIAnHHxCyB7WgSHZvM
RJG1GHdxz68CPTNcG8EiwRdq2PeS5RGoY69OHxPWALeO5oolOiUdDCgSJRyX1Vw7
nNP4oI09C2ZMLww358NVTxVvZhPmXU+SMwOR34eRZzzHTQ/xcpfrQ2UjUwCE++PK
XVAVLXXSyYn6ZuTs05AT3qEdwQyt3QkpMNkiFz+pavR2RuRXOeenmftfihjU4PBl
ucacAgVCr3+euZ8zkJUQIyDPKCI6Zfo+Jmm6TgzmOHGg+SHovOE4y/udAD4OxJEr
6r0SzRCb1lh12w0glT2qcTidSqOIzGhL0ww9UQzLP1kh1fzfiZyW+V3DFCUZ9HDN
Xd2a2Uc1jvcaWv4LnBEoTWCtNQGCARi1T3HtBE5KE55Vos7vlhlcKySg8aT3cUEc
a51D1waOoTKoOBSPlphm3osYqb8vLrSl0c4TqUiHuVdtD2LxakMxPFkGrPWntxli
YYDC/mWUlaaOxd2ADg+y0D6HrjDiT9Zb/ztO0eR08yBbBP5WgrQi6l4FhSF9eWRY
40CCs5O3lhbn7gdzblfZytvgvlGEDWP+WS9ECrhg/L6Eq/TYC4XXNvYpPV33YCHY
54BBcneNohMioupzZcFbW0uuXXTB7qXQKc054OT+4pim6aOTqNLYxj8NIST4iEpS
5SOO3EB9z0Rnq5IOWN9/7z2lYmQryOL8AyTUVc/Hj5Wja99eVNn/wmLepg5tABS2
BVKJ9ZHXSEYQFg7hymDumQnxZuwogDS1zAW+Z8oBbqWxz4Z+w+LBEM6pl56KRs5Z
U2LKrgIlfRzEy/YzCnF+H+qZON+DELzedvvM0Eh2MdsAjA9AaGTQZD5QWPDXFbCE
EGY1Ub9375xHMcHkJFn97ZbSu+GFFfRn2qBvwyu4CWD0S3QRCW7XasSZ4z+6Gyt/
lduKG1F2vD8O7fcx02Lgm9RsL1E//M78/kCthKZEu705lv2bd3sEpPrf891rPSZJ
ZazPKRg5JdNxBRX4hHfMMNf2wwp/r90tuv8+qqkvErreVVAM5WunMGke1kWSry+h
NBm3Mq3JbaKck6iQ1CKByx722mffcxw62Wrh83pmtR8IzqjswOHQ7WpHxvEYN3FU
`protect END_PROTECTED
