`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vuiiSUi7x0dgzzR+QpPQKJqyaqPSdC7Oy4ef0Zxb4m4oxa/JIKDo8DeZGTB6WvOG
qkd9Fk1LycK4K1lu3AiT7gmU2jUmHMl0OuGwP2vEwpMXbQ/AE0CvuZxuHx0aV6sg
37/TIzHtDo+q3qRndkY228kbx+uHdE+EnORdWhk3CiLabypxk474W1G2qf35BowL
X8booq4AN2Ts8ccA4aHUVz4fG0Cf/62eeEvtK16UMD1EUlPQEf0d0JoLn6gJuDOH
/YEzO1O1zO4VK2mstLq5QykoQtcmuBhDSO44P3w189jCWxJbMlgBOfBtODr/VZ5c
qmaGgooG2yGFlqZt+2k8NmCN2Pw2eG8Hc4kbyVDuMjKIylmuvFqxmlx4rvj+TjBw
b5W3ZsA/uP5qmJHaTM1d/9tFW+bMEaaYke2j3wbrUpFbcSMM4sB35VyItxzdknJZ
pUq4pI1EsLV8Q4uCTTxyjPy63hEVJQDzCbQQNRM9FnXNUfkizec8sDYibq128pwz
WIkyp8ABM4t7OGpNcyYWHnGp/SNJGoKclDjRVQHtL0wLZ44YCMaGv3U3MHmBuqH+
`protect END_PROTECTED
