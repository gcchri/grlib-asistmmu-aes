`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HprggkWkJK3ipqguEUkzNGImMt2tPLRZS6Z1T8A/GyIy6MgVJMAZapGFDvtx89rF
SxnZrABQHwcnQVp4RK7FdP4m77FaORPH8pw2zUpf5LN/L7zvKEHQI1QVO6CgWqz3
wtsejiF9ZFU4jLjV0L32jgJSpOvTdYkU5DxB0vqtHGCeJRmpHsi8qJQ8pmjkYGpW
ZesCsuUce5/he0x1aGWzl6DQsxqQkZ0/D69J7OQ989zsyALuzOGyShB0wHv1DjNJ
PSNU7O2ZilbduxRX+7TN7/fP7/Mm75OYKvun73BN5rrtQ2mXmlMXTvCQ5ZZVvyeu
IqqEMP26WlEI97EdUvW05rcb70zZDouqbei1qwAKLJy2g2Y9tPRkafa7+D5mYI3V
kEmG8tsLX3N+LX7pGkt1N0Gs32VAMRnUMejAYbPBi2o=
`protect END_PROTECTED
