`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W866eVWooTSnPTWCPc8cuz4yVILFfaVQvSOwJKxEZz82TtXTz1pLhQ2nOBsSJmMF
GqkPnOglwJOhiuXnuoMukKjG9blj3BxxSAjo4u41l0daqNYmlQd+I6Q+72vTj1G3
09hI7tp8TaJh7Z6fYo3YnjrIHJ/fe7sZ9m1ZV3nM4nlvh71Grai1AW7e26uWC7tm
puwmYrxL0mBDKwmoy9Z/JMhv7pDJY1n1a9CittSdYr5FA9vPNKOH+9FAARmui1lA
OxknzKdATs4TVtt0JSdeA+yWkJJspBje5rg8xOyCQl9zrHhf92Xbo8aVi53aATI9
dTjLAKSSdSmaPCSqWriUjzHfaPXqHe05WcijAZpsIe8RnUSGl2INhBJQehqd6SFT
l1ASLJw/9Mk7UD25dh6fRd5rIxEyPXZjjnzvChwMj1/aVSaBYxaLsat/0xkI7F6l
yoWOoL9NAmxFWYYnt7kvftIUkqkDT9NPvEAkedUvj0AmfHZjL1BJuwK5Et5/np5N
N3EV84Hv0pbXJSHcTT4uzYRXYZFysx/DNumXxSIplGlij9stUnzZAn8sx74Pqr8e
NiaGac7cBvNV85P1uXjookZSQCiDJE4SNzlBNSqVCa2JtE5GO3rXsfeZTjI3L9JQ
OZhUqBFADYyL13abDU5eOBY65zgTIkBMoO7Eyg3iI9eajnhasxtyqdIZsGuvTxuh
6vBpmRzxZz7bi82Qu91yi0XMTEgJQTHkAmGZNYOIj20=
`protect END_PROTECTED
