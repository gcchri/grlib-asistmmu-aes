`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c1Fu06gdIe1YzP/dnJ2+bv/FwObZgmFnIaqTnHlijnWILeHSm1wJ6F6vxE6F2Lxn
Q89iF1WZTL/hquuoO8/p0QN5EKKvhFQqPnQh44Lt8OIxUqiTWFPs8akwlO9VaXnj
CsmsZNGw6FvBl3foRddyTPdR0Eq4jwsdi/165ZvvIVEsoT500BB7kQJ/Iftlj9Xf
NJVaqZcckxOeaZ2RourLmXTzVFHoAlaj6HfWynQ77OJqG7N/2J2ObyisNw2iADG9
4sKOXaaVzw3GxA31SBTFpExM5Tr0WBLETiQ3jBOXbzA=
`protect END_PROTECTED
