`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4gtNYDd93SvWfAvNrbjFr5IAID2MbVUZtyOs2NGDJbm2T0jyy5z5Nqn7WtqLk3EV
9ECrvx+d+K5dgCeStlH5OwE7hQ/zNPotUpfFxpIvbWXURvvWMzKLd2pKJNHVOse0
346GJELUpmio8J8MsBG4LiW+ZVDPM0EVhipnAatj0vADSlQyjeD7Z4juLsVoXx5g
2PBHibYsdCfEL+qraANuHeGTGLGv/GFPOc18xUvDN36S2df25B1AR/xcXBjWn9YX
3un+vN0xZJv43PHc/cKHaKwLN49DTAHbtl+bVfh/q4xz94Sj1feBJ88j9MzsJKSa
GNXeSijD+A/sAO3IxBSZcnu5WVTIRDF4qGCIAO+1bkU5J+VAcPb/0gjW8HFHuqf7
YzEIX4GIkCHrjv4euqcuniRorj8/Zas54eG/+UTcA4ZRz6gjTsxvn0BNTeM+tRPQ
DtKsN4hYWTDDrYmA0PzXy7Qdt4e2gZxvjIUXEUsbavQaZ7eRK/DRjM00svRE2MPX
`protect END_PROTECTED
