`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/jMW6jjJ5SkHaA140oF42SaAWYtp9TSeLJXONiXi7VbvaUKOfgI7iph9m0sMq9fP
NIzj8ddbfiwojTRmgaafjLQOG2CXJ8PpTZftnO2fgwR/BO2o5XmiZFORb1I6N0/f
zy8gmAD2HSDl/GOYGiTivfiNJiXn9VIqgaExoEipJ7K5jcYyiXs2PsHIvckWWznV
d5Tg1ScDFMlmrC6LDyx7yzFTo8IHLWKJ4LQfVzlA/A5gxr/ApKCbJIzVXYfB714t
WAsImJW3wJ5jv2l7ezhhC5JZgwPETjqmf3mvqZChbx2k0ONE3kr8bODBeg9JjRVY
uZ+0peOh/69EJt8eSExdfpOgWwJ5+gAPbVWQ8KMiSqNaZZNkcwvOJPs9t2AuBrBj
6u9zBOPZVbeK0VSoU2aeqJOBun03eR4vVRJV+HWhBCPvbBV81mmmBSdU0NoXdgkx
npyPWh6rp/c+5/+DzuoCmG45655MwRrXmXjg8cXegKtqpwE/q0dciPP0u5kxs2W1
3LcHYc007ZLmIxu2gOZTgeaWOkEoV8kt1QWULBLsmKtiLa/UGFNUWuorbianY9qA
cibuhFYz2DLBshF1sGnVEE5dzIJRDb1djYqW3KtmtmB7maCCIE2sX5tsT+v7EwnE
nuT2xeNuFmeXv1zbcQpBJrUwCfrWTOyajqef24HGDHM/KD/T6Cm/Fzb42VKRm1sv
Owv4PjhisK85gADaJl7g5Dbl0kkzwNuqlqwsRfDOfYJADM9G8ofoHrJyspEZJN6J
spjALfue3X1Xq5jzPMVjF2ynrLobcbhsIBnFHL/j8ASF9qEKFmaA0YH76GTlMicV
OXk5uRS50MqRs53j6xVi7GmWuI9GYC3x5CLtIdLBqLK2MGGt2Y1HjNrw/5tQmhYi
/bjI1bf4PIbjQawnvQRq6Knh2JTyDeO3cHOzU1I5XqYTELfPvh1az6kFhoPSeX+D
FoX5PXq7Y+X9MYxq2vrd6OfOV5mDyex5Ul8cHFba+vI2fHxJPF6fDkiVnCRZ4tM+
mFg7o/jBWhtKpLWUdGGv3wnKHwthrC+Im87OV0D27QpKXzkxD8N5Y2CiaLAdZ2cv
NgCOttcQ7fr79VSjBAnPczvlVPyeAUobnk68zOQA4dfDEAe24vdBXZljqkZXBhkN
6c09SeEsbNLej5WpQUI70hrE3OnL9yfrjX8HPK2JtMxjOvZs0bXW+gBHQAXCjOPQ
1LR4S/euU9Hxo9S1fm1XgiwCkA+hgr3EI7vC2kDC6H5AXDjolcx3bOedo9dbgfd5
rUGc7Qm9w65o+YFENO9nrNA2/b+QTd9QF0FulBcE2z3K7FSyNuPPMcL6zJnsBfd7
2pGX7z3CdlIXXit+jYGcK/UI/mI3c8BIjKj1mf0yQ4tG2MBvyDu4fbzrrGC2iq71
njD1OmztHLRAmHEHKS0SKlvKXmdM9uupSdyCWr8P5ezmVxUapJ/SYYrEpg4SPU6F
nJVd/YAQKBTbqH/Cd40X7Ra3Vfc92Awgzy4UXnjMqo6HVwZJA/KDpmyKQMiokZ2k
X8d4ISvYZbx5rmKOKaig2KJS7gPA0TUecaCmo0svpSVGlfwqE86ahTf5totYH8p5
sYed5kNgGZssRpmFFdfzJN2zbae3L+l1jhhgwQneQEGAPbHGy2fyvizKcu3ngxCo
N9tVl4tV/Kw1DxRHb9A4aAAROa6ecuCjBrOkC8zCwpyfW3dzZ4nRW7MgM8tkyyUJ
1ELA0LOJhYIKKbLI9EzCFUlZDEOsfgq96JXG/JvmGjjY2K1mCt0y2sBOjZksZZ9k
wgK8KZbEyVbtafV9sHdRdQ5MF3s8V9/Xi0li/n7BWIQzxCI2nflCNuqNYsc8Jzlf
lnujx5jBLbSi9Ha6sjXHeffMIBQw2dKiK5kHeGwoUiVV02vVQfu/K4x5fHzBf45F
vg/UKieI1cOAGlVKQIKZUjlDH9AUolbpYsfikcIucmbInEKYyiXPja4Iov0kQQDj
+NTZKUHA/+jNKoABNDlubL4eR1CqOtmVrA5ddu+pSWtzUS5Rj+rCBCMHuK/kpHHE
KGScOYeg/4pOn3h/LQmdLt6swZVbIpRaYP6WXnTmStfwTpoPgAGMVqhyaSHqx17N
gsA+QxP7XTwUGyHeUSYvY7c7Er1uIN/MlhWvC5BkF9REb2FqEn0m+ryMEm95kFDM
LRjuournGBOrD6wYpKPA+L2phhuX+9BF6jKonWhbnr8yzaRjRx3Z4NOvZ3rFyMH2
cZv00+dXxVZiGcCWbsejFq1ITmZZYZs87KRMMN6mTHWDosr9LqcTBoCkAZ+WzLLe
lJk68LDhj8yon2PT0aJNmzkMYEhBMiOSGZWzRUy8dbcw/EE1B33/oTASFV1Ps+Pu
fNY34GahNKg+tBaUsAiJrw==
`protect END_PROTECTED
