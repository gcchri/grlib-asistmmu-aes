`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7x/Caf+ujo4dV/8+sZonQ43+Gaa7uQeUK+Ulv5jr5sc3S1SaHtd/G7iI3RHnJGs9
iF3D7aMRkQrlRtqZ63Og3WwFIXlcfGWTu8G689p+X5Q/xsUTrTydcnVEe4rj1Kk4
NiyUIXkeuGU7GxI9KpS5vHVmabQmiIFuJ04GWcruv5b4tL0w9sSx/bEN6/z7W0nV
WMk8QgAhIV2VSUThMgJVzKKl+pcTfpA0fj2xPuphKIL3riN6f9PIU/UjHP4eZLQk
sdg/jQSQmWhJMX7+yFCAFOsTYMOQrFv3n8N2UB8ADAWDi4zrCYikyF4XJT6Uvy7J
EyRspaNx85BUEjXsKO+hVE+OC5i2BPLEZjxFGrj6pQ5uICBa+j/gsCiiLXYtrplb
h/4SVHVO2QO8EScdHl3SxcuHjqnzsAoZKzsb3kpWY9n34MoL7XqSWwe+dzNDmkDr
L5FuNuGa/Gr6x+OGF6tPDWP997Eqe6DbrEzrrcSoSLbhOaq2hyDaZtDZfMOrNRk4
F2NzgGjPXDsHii5FvUE4/5MolN4MpB5FxXu0tSCxlbh5ORisMZ0jBIXEJe4dypdZ
CME6uYv/4lvYFo2vniubJRD/eDyDCMUZx313FCR4Tu8B20zY/DpBMpKC24jQ+Q4P
J6gV0LbHGaI3WulTPviV0RCWgMB2+RKA8NTLxT/DOsC/vB3PxUjXtGEncrO3yuJ4
TZ3fWuo99ZZylG6y2W/Zu64KqEeqtw4G10bPdDenC0D4WvZ2/Vgr9vkkT987pr7/
rtNgyBuUJ1NgGhGFGUuKqwdjvOZuzAP1jyVuSBJiWhBzbnvv3BegGs6Kg6bU44zf
q30CMzpwassX7zuoj7MsTwz9gySD10w9Drwteuz4a7KIzqMvOSVSWYTJuehNHmkk
gAtnzwa1w2+qQVJJwlOx1nAzu5v8pNmlaK/UxgukROu1AM2P47hbaBBAuWc/BTtT
eUBg5hozN6F85dhrraFSCkb4Bg4xsCgSjw0fztC/h9jfHXSGQRYpYwX4ug5QqS5f
/u9w95JwqpYf6lirAyvQGrSMcs5A462i0P7fhXIut50uM67z7tYQbHd8iMtUf2kK
sdeGRQS2eet5RGqlkSII9q/w56EG+tVee+i6nHHU/5mMgBKFs3qjEaVmXkrHRjnt
x9MIgjHZiYl7Er2HRJx2LoTwALAzV+dJVKFrQTF9p6aMFOcoD4h+vzK31pG1LDXO
KkIx2rwTBHutj0M2jLH99iLdYhXYQZBfyzkBJObWR3sbC8N5pshXQeuNR1AGRCi/
EekJ9XUUd42ScUFPZYgnI4KlX7y0osMjMtkDqs1hkQtjFlGAPKIyh5IE+6ILqAdl
l60YJYqCUwr7zMWzrFscIL22dnv8WS9oVaP1CbnNCJDthDNXdULT6YSlXEYc4TLd
kag+9VJh3u6sAx+VS4XZ8EU2NKHPV/6OWaESTQsTNEaO624vWeoTl5X6JKlGNrOX
wLGv4xsgPMR424KFwnfMHSbQhVSJfn9chtXo/d8PcKP1//wyz+sf9QLvf5B9WUE7
RDzleeG/y1PXrbKgFIqaD7H2W2SNxC+jk8VMQbE6B5E1kNIekRYlWHg8bkKHo96I
yFuYVfOxiaS+vsb7qMzCmfXv/DcxLO3mlXNUXty3M7D5qsOuM17tUrvF/hFXeZzM
F2hbCLGnJb6BzEj9EZukvcFQSCtY9qeS4hWSqQRF2feUu4dC0Rb1d5MN0owGEM7S
ygW3nZldYCPianT/OjFf4xHQ0j48NhZRZ4RimeDNjORKWolO+SAni1C65aq5jpPg
9CjVF8nZruThbkocNEPSZw6AVzBujQi1DlG1bW5kXKOzXibkTlqNJHUJb1j74ExO
CdEd850iBLV7nXHk8JO1xxTRm/Z5GfU9CRNRoYFyKJJuItjgLfr+UyqRsm9RfPyU
udfRjCGDYTGS9hsdC3u5rvNAyVyJG2hsXFsQ/Jjv95KXskhaSg635HASgQJAi9ON
OF/St1BCz96p9V8npe4ilpu0ZeaDxzgJQYidOiFb+MZgTnUZTPyv2zfj/50t6daZ
pirnZJYAX0yoYRuv2POdkdLZFBeZVQzMgagWHlAZuyIu9FQ2/7xOK1FJW3VOxZaD
Sme/z1wdYn0gKJ0vQ9skxgP1advPrRv9EXLiDrkV3o0=
`protect END_PROTECTED
