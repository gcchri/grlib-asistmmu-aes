`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eWfIMDucxXzScw1Yu1abZdzU4BxLZ4ufj19AdgXOZpSFapy7elVEtA4Zp15+z9Jr
40yNeI05ZF3BZCe8JrLdMuffeky3xhF5CUEAbQ/dUrZp4PrLRttHP5MnmmLCyMEX
ojn/Guv+Pkn+iWuFHj2IzFU1L7QYiXVVuxFGL55WqIf7T/dRdyfv3+1FlcxsN+Zm
jzBTqZvynRz0hpB3ZDsCA2zZBZWJWCwiCzckPpIruO9zjkQGo0Et0P0vNjVEmPGD
WoT89eh0Z7QJdhLfnHFC/y2Bp4qIuVaTrJX+dLr0Tk0SsnPygUdtpupRqiO4HpxX
`protect END_PROTECTED
