`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HBCJJsz8aY6dT7FvJKEJ5iNwP6DY1O0kWRYFfKo7cTBZGO4k3qriFdzr1KjqtAYI
2l8A3yZAHBT5sprWaX0BUCLjmZKQOfsMJeDWfx43C1Y2fT/b1P0mg3+FfV6irTXv
jw8cWwbOSbHmwbo8yKc+SGXx+5x5yPwK0gBbpRDqy4UsXelxGvOR22U0PNAazblS
4EKC4sMB4Pow0D8ThLAQQkLD+nC0+dF3GUymgQEptnVjtrqoNNT5jO+Ty6BNCT3U
hk28pQ78JF34xQfJ766lj6l2Khdd1NrQT/9gDc+zn11/EL4fvXL9cG7BgLaTvHEx
LY48sAB9+j/g8Ej9PH7jNUj8lwKIT8nkVA2WSim+SsahIQus5qn+ZhR1qdZ2JUm5
sa8jL79jZQXxeuJ4eRzgXO7V16vA8885SIho7BOSQDUFPiwS69rAzpDlQ0i+f1cz
`protect END_PROTECTED
