`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lmiOBJ+04irBuC92fF8aun03kZRrV2sfpmMp59Wbv5bC5RnlNvQmTCgMf9ZH55ex
rzXI9QJcyEqmuC8g7bjctX1odpZuSxiEGS6cKMC7WZw5ZSfq4wg9elAPPYlVB9J8
YujrRd+M7DnZzDyBTQC/wgyVD2+H0DI6iMIisactGRUit3yUYt5WVawNNoNmfuEb
1azNR0xjdFyECgf75GsnpvGPV/nRP+sU5wu6uOXeaqrvyffnkjfFbM0hyvv6Ltwy
ZMfiano+RrExsuXRgixv5A==
`protect END_PROTECTED
