`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lJ8T9qQJOm5aGP0NE4iAO6KUk2nMh8RZ3OFeU7AsyLumrHL8zb0s8W2rY4es4HZz
9X5iiJ9e9UDAxYfMbbKKjMC2Aq41L2mfvJnAwwuQL4wQAj40fBACtS1vXJHmc4Vy
L30cisQrYtVPTk7W9+GfxelEcX6gV+jXEqJmNu2KaDFHndF7voymoNkExu1XRwG+
a6VzDJjsUS9OnhPBHrqrMxqG8SHyTy2D8a/yjVJHPzf2kfnj/97/kwxD+36+22lR
kjWlx+/i1acCGBtEPNv2tN2GZsGzHbLBMMm/GDIdKveIKIsjwQ30DUI3MBc5wMk/
o6SGW2IeddQ+Xzw98dtPYuKPHzZ9KLWOJkxhYF3UM7yrt+z9bEuySa9epMPfnnfR
0xFds7/2IKWMuXbKgfR4SfC3FsNlfL6KAk1d0EkIEzjiIvzaUXGdM9z8cfFgxjLd
KfgZBSqLZfpQWakBPoiV0g==
`protect END_PROTECTED
