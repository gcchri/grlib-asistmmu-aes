`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fx3xsBzlJsO5dmOC1C8fEI2fMBfVtyRoqK1g6xLxYJDOw4qvZgAWZmzzHUwCcUHX
THtguv/1SeVLqa/6hjKiAwWSPi4xINEMUd6sJ38flWyL/R6IUZAc6cLakCQIARmT
XEwX5fkrsyg8bGE1ezVsKAmiskBy3v6XjJ8DD1jc6FzOsv+4F+45uUzd9xjWRuCa
kdfa99zWnVtPf6reNg5IO9r6Chvci88nar2GvaZqMQqrolbe1ISjNHG8tbY0VU5J
7YEkEF4I+oEcqd0kZ//huqqMKj9rQu4qpLHU0OwseNF+6KRvf+/KzkrGuWy+ARSr
DmujgZIEiU02cfkvvypaIKT2auuOotqwvDHNC21Nd/dp5Sf2jnOA0eRB5TWqUGAm
HjJAMonDZD/8Bjy7bVqFr6HvDc1mKcm81ZoYg54l4r+lPsoYeP81nma5JS16Y2Je
5H6RW41YLEH/fqeNzqQumIRZBn+L4PpeD20etxey5PNAgFBR382gxe/P1bUJdsts
4CdjMypCg7sr7vJ5dQUv+8Jt2oSI3svn2pDToAG4cZ3AcnpCfZImfC6Oy9TmWSty
jb3epC+GROIfPG8kpu/xLQz1glN9QQfd/uxecyAXjpP5sfBHSdTu9UOtrphMvs4g
UtPMFT/eyNfVc3hTZuwWpn7CnnVGY8/wLYue9q+/v5lOkqLY44EL8y1KfjjtpwKm
zsLzDXzP/4Mzi5GRtZN2btgMpVMti/fwLZ97Rjnu5UJUvWfsButZ2wY6agVpFqAP
3hTAlmPo8mxkPk3VBSSF0hJFThBEMYWKdS1aZ3vUpDSkaAsoweZETvXfRT0rjWOF
9J+yIp8uT0NW0uVpsVmyJW1+XW/lbpfSsvX8nPhbPGAKeFR2Cp/8U8ZU4l7nY9E9
e3sBRxoyraqgvEapAkrEWsFOpn85qvZxYnGZynw05QFWss6IYswu6W5v+TdptbF7
hVYRINY/fv2XlEroDbM5swyhM9dTZ1NNiUw/mMVcuW1iH4xf1v1IVKfD+RW4hm6l
nXHZWZpLh6NJgGGR/3V5JCJ/6Tet16YygHgaRT0sekJPlwwaBTnV6u69Yj4+RFGs
EJ+dzWgzt0qwTHAz+IcEviumxkNeJ33q38xie8VGGHsDCl3MoSqgfzT5FH61YeaZ
vIpc3Z08G5BGPCAL6/sWUE1hkBAliesd2yRdOLeotARmt+V2VFuAeWd2xMydh289
9JSHaXMUBcT6x09ZiPZPJR0ONr1wifv2ZsTKmiX9vl3npZXC2J+BsdUNlUBDDEw3
htm6N0Ky7fYiAVXgDDcsp7ETqAiWlS5qFlQoXl3AnLTvi5YFVUgPKcbwCT7pJjfV
deAYg9fhmHJycHkTqV/Yv79idkGj4rVhpHsA2GfIH1tAhMDEw+uiMIdm/OyeqiNM
IhJR2d9tDP63Bt+MCDEeqsYFahr0Dq07SXjZs1J//NNf0ZBXpnAIClQ9xQaTUs/T
wV8nBZvXnlFSivYbrrk0ie51llEMeHg/eCuRUkGcZw36sceG4fFqMVsBI8Iaj4RP
saRhqrO30lZlaismHIHMpjCJJme2PK8YnjQiebv06fZnKO7XdO53sItIn+Bw4Y71
MSl+drSWcemXaP6LO2h55vvHmYJ+iVdPG1ILDWRzhqAeoP9mz8SAwNc6shtylURg
2viUFRawcofz2u2sHDSSybhmE+LnpwvFNiKj9sDwejaWdbb1sXz8LE06Bw44q9sL
r14Xys8vtCJsOG3XK92WDFQFFH6gMpkRdPWIPp9IOJ4VVbUEU/E1NMZGdrsrubTt
VwJXYmKYNr8gycIYGsxl+5erxjGZcGeER/GbSJaR8XkoKMQN3GQgue/liUNJBHTa
8dM9Fc9wxXWNpJI1Z489s6emQZCecO7Z5ULVJv1fxjJbdekGs/Ujt7hLBqiEBGmh
TORi3oW2TTKYi+1/dBCCP2KF+tiw002Xu+yJpWb/UqxZJ3Np5nSF2CJrJKdrzikF
KJUK7oOvVT7vTy1tl6sVww0ldrCSOnFHDCmOroNsjRAQdZL0uKzDYJW7NPbYhyQ/
jBoG3nzbhOmi/Oduk+yQlH5CdPrq8Y4U729fgKH6DaS2TeZ639Cvjdmjz5ZONpXu
FuV/EVEhpynMCmdfAVGXrDAWecxmh3ER+sQjzdr2TbzUAGHXj2nxPBJL62aELrIq
ZpS6a13IKi4VnOHPYkdgzo2BqM5LXy8BvSQ8oWpViHlR+aPBYdyboI2wHCYJcXE2
diBDkrVebwsRbcCq+9iTedOxqkpx1hZjXGqVRYJQxMQsGWJYQ8959J7QtNZDWFG3
VT8IXL51qSeKE5/W2bSZ+PsIaTaiweH7eWqydYGDyXbG6gdOaYQvHWy64lTWIjOn
`protect END_PROTECTED
