`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZbmMwKxolb7wbig1Md45Rw/K7b+aSZlb8zSMw7hmg4Ow00Lk+ds597Lgpst1SIsw
eS9+koOtoqR2cJNgKua7391ZTyVfslkEY4ul9rJ8EDNx2H+TInGFQ9/bT2XGbBY0
x9z8RBRKRZ0AkLWWeyhuAD3B7ILPj2Zdn5NhdiOVqDJxCAnQdhrQJI0UhqnTGshE
BfKM8/GHdLlS4BKKzeqJ7v5CQT8aI9TP4QGvFCJyGWBBUVM/DxkgPVLWBYDljxeD
J4sdB5rUEe/98U7MCs9GCifMHznAfJyMXNn7ihrlEFJzjqbT1JaKAyV/uZh7xgHs
k2rdeXRaTMrY30F0dSesPU1cICF2+NI9xt/7MvFt2um0OiuAsgKb8a/MlqKRaGGD
RMDOT/CXOWWS4W7BiTnR0FJuWe8ZrCcuoh5C3UK9dY6piDAMnqMwwRhneEnCDdSU
X1mCcjSAJp7K05V8u/a8CX//C87MN2r5EUQuZwwZIsM=
`protect END_PROTECTED
