`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W0w6oq0suUVUUY+fgtE9Jc9DtXnFrdnCD6jJIfMpRa2cCq5TR7anJKCNDAjBchok
D6GKbHZTUwxo0BEgbRWK/Ys1wZZTlvnICeVOZDwwvnSWqgxUs2hv4P44/IGzZGq2
9CgzCquJerFcJYaQmGO2eKTISWkrJRDLzyp6wegV/spFa4BcsCdItiwkoDf6XA3T
gU383TFO93SiO8aYiaN4dNaY2fqwJ1FK3cXk2F1HYCyDNuk901wuyLMCgWU9rz3h
7OS0EF7KDE29z9ykNcMiLbC4V7hJa1VlTyIc0IsBcphUEp8FNcPp0usyXO2FP3je
WnzLFrF142SAdta1OXpLR0WeI3JHNqvhT9Jy4tILQ5LTUqGREnXwg+jQPNWO12VL
lcaZ6YextjyBmp+Ny+CtC2/Jh+U0ZlocZfyYXxeOYPvxV3zEaKkBlv8KBTN7U1Jx
`protect END_PROTECTED
