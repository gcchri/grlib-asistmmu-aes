`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fyTH4ya8BiRlLZF60WiuyepPLb99YcRHds8nUh819GalIUIEUJWIFW4e6r1AzVqO
cq6qw2wwIXgKg77k9I9+L3/Rq7csfBJ73GHtFniHm885JJltqrCEw/tJh5lcT2sD
o72k3CcpnfRg8LHLDYwALIt6aT5O5PbLfzUsTS/7u5PZNXD0NZJ/U1O9nuSrde6y
QaJh7ZYFGFUm3y4jholqEcFk2vS01WrpoTC+WgpQvOpau4YLsoZNdpdZKHKKfnQV
irAkzMsOlyMV3U1nEiR5FDXg+jZSuA7OBwuxgo8RWuNyHKurYChkm8odeoxXOtX5
lZGTUippjariMVPCVFfFS1utyUQWq3wgf7eafY5ZanF0rD8sQM0CqhNHlZHD7BnZ
K18MkToOJpEAtE55tziXKG0kC+Uro2IfYiJvWB6K14JINRh58Qvku8USSmgKU+Pg
uzUQCYTqAfNSp8Tv6KRBryuUDbB1YHmnERUuXupYxLPSZJSmu8zajgyEXVvlzt2E
18mReZiVQl3bz5bD6pUF6jvBIhg5QlTkX3biVx34h3wakrAr/a+CZkItOBNk1Ktk
37tid/iLk4n31mBbgt1uD3j8KSScb6NYiNTrjBxwVcITFK5F59qgewhw5RN+R6wo
1pN0r/eNW86e4BOgIdbrIXtr1xjbaSdyGlc7hAUzfKJONd0ysWH4EbKEqI5fEncF
kGRtkx7rqlB4E1m4+kP6g3L7XwvjBzRFo5wt3GGppHAeBMvmbOgGKWBVw8rMA9KK
h0blCCRwt8rXzNy9OBe+6NnXh6P7Y9XiHLgMh3t13ouht709uETjOp4v7b/Vij8Q
2yUpTedBhqGvFULWpI/s9YOaEuXdU9UEXCdKUFCMFBRT8WehegSQsaqJpgmI7dZW
Nh0k5A8KsmG+hsbb/ToyfZBfbFvPepMlzNXt4pFNC7c8Xrp34QUuCFyH7R2vOfzY
ynY2qEzuvSwYgq9NwavmlvVvanbCqo4a6w61CzkM/CPEqFGsp0Z6wsEuEK7kfJIK
HHn10umiVo55HDhQo89iqrfQqW91nocCqcu0Nd+16dW1/b38G7KbJuiTjAkTdNec
`protect END_PROTECTED
