`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dY91hNLp0QOp/cW+bjF/kFmAV/EFHOZ7UwVqzZKHpshODwzoAL30cNAcOOnDzP+W
Lj7A3hkLlE/3YUIhAUSJAPpJO9IY3s9G2vvbuG0h6K706v1Hx9i1CiOxr4/FWxxo
onfjMZ90oTanuItEGHBLZct4Xns4OqkhUFXpGU1Wwe93AN+iItHTaGEdf/vYH9Mh
+RagQp8rIQPAdXhT2MuAXB7a8Wy3d84R/nIr/AOgOrVkziUl+ArOJUu1ik7tEXC9
dBFru6CqY3C+DUZyfy6X7xStmA1yexhl8GzIJTzY6IzcOMXngfWzAJV+jCAEd2tM
B4p3XPnYKT16jQT3qcIaORsOMIvdHDc7i/VfGz7GPqy+zPMgRfEvUOmOhSaG93cS
XimCQ7pUc5loQQ0hztYC7g==
`protect END_PROTECTED
