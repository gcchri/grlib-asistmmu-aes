`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gWReocxUttLxkKWIXdEuImic1U46g4ZwF0d4FEDjmFKU9krBnJgpd+kSTfNZnOvu
XzSUzhka/vWI+9btob6/ODPf+/2g7Bwers+K9kxn9JvXFbdZwbDRgvIJ4QaOx2ez
4CuXEgn+dMGbYeQWKqApH0Sd2+4YaV/n5DReqD8sjI0FTTMSgQyuAW1gTQ+0aBX0
3lWiTvU05r3fpSxgsuUu/9FzptJ8Oj3jr5H0mOMdVJ5n4M/eWKruoCPPRuiARheN
5qlcBiSnjhuFs9qS4kbPyn2W57Wu8b34u4WvxgsstNgfUz4iZmZ0AK8U2wHz+8Dg
Ln8LUAEqWRX9GuBwOJ0H7bcTlZ/RWWlj4Nt7HAZ43JZxgNwbdkJvwJ5tXgSkGMSV
`protect END_PROTECTED
