`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z7SMhMxFtjFc4mPxhDc+3x9ZMdU/pkxKDmu4t0ev38mclGVmuCWjzo+/BRgFJEid
bPPaWpUlWtVUeZufusYfl2uMBdLRj2lnwKkINB7LJ8I074qJDZpaw9CSGJhMUTfv
kirSpsfqT/dSMXTspb4KnFvbT0+WEqTbi+tXwe6fbrvSxS9J1Qdzq3xO8nMwwma9
w86+IKGK2Dl9X6dtn4LtmIfH73pg92uH6xHwVAECSUgjaMLvQ5wa7RyQwSjfkC/n
FcqrAdv3uRUohFB9irHCf6JnlAhesmLYv11q7Xx1R5eYguCnTjb9or2XehzJTOAp
ctVN+ZKoHBMCmoU3uoiHQPk6xtBhf7MNSSzylSREqZdNa5hYWMFmag5rwU2r9PaM
DK6XBCgVulWZFx1xh8JixocnGzrIRBsPpk5EGfWLx62EjE3x9Mgqb9LZNBoyh4nk
DglcSr9yS5UEf2Q1+/nTG//2gRjDyV3DNJL5wqa1fqkalKvD1zMkZYpgYyzton2w
9s1F9QdpbbWi0HTl60swBlpxZ6/PzujA9zT4E8WzyNQyC+abmLPh+9gwQV4eRAQt
Owmejq8cyKsUGolsfYtC7OCtbNaveftnoBpvCHSWPfCWpgeZ+9Fjj4KE2yrwsYHU
1CKE81hoF93hXbWEVp1f67D7DSxZbSqDvUJRiQCY9fehY3uzFZi9LG58fKxEPRet
nDBUQSXE9K3HB+X4s09C808J3XVR3ggClnJf824pZt3VJ9K0Q8HyI9D2N7a1prxf
tBVt7fH5+BNmWZpIwLK3W5IuPwQRJxhhmX+xwBgz0t0fabYgeS1tTTGGg3nLfotX
S8qWtdyXkTiaV5NPuO7MBiv07OGq1H6FcSfOEjwQzg+PrHGXm70GBZOK7Q+3M37/
QNuI3sdcePNSsEwG351PhB463Dff1lHehAdzJRyNXlsWB6DanxrZVqUO5HL+g9qy
wH3cLEHv3cRRDzlGcSwFfceDNRMqsfqWMV36a0SRM0sbmeewOs+y65RBmIPWb/EA
WwNLnVEIl9xQ23iQlHWxHUG7rAPTij7LAgwknriq+JNH/EfX9vhPncEqQBSiG7oL
EMF3JHa/HUDkHHQtZkLFeG7n8PREJjmWVNerP1R0GWz+aFqScCHMj+Bkc+JUMDoO
Y95rNj9N/F5Drbu7/+U16j04GTTpSjFvLhV+IOxmCKq3E3JUxutH6RSh/SMRotuI
NP6W4DlQB+ujpKrTbWLGwQ3b3GKiSAHACXA1NbFRNsuKz5xEmlyKuK3CY8aaMhiQ
TLige4xAkVsg0BOKXOIRg7923sko+/p45IngoXnFT2u+pkRZqT9fvzlrYSRjmu6T
PzxyeNVpUpWShRP+3Fed8mSJ7oZEqOVRkXPq0brRoLU=
`protect END_PROTECTED
