`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DUPwiD/dL7PVwsOkILTm7moc0qAri0f6wtTVADCckwHeQIV6YY46VHdbjEpmACpA
5DtmEi3JUFQVPDt8W1uhom2CCCEOWa2BsBjHN92Mpj7rHQURH96c/qo/RpErHAkB
/QNQgINkmaNZt0kVfNS2jjSJBU6D6pAoMMeEUF+YJQ5hXnT8mRZj/ED/GTpkz7dW
TqqOB1hR6zyGwtyXFqu0gAzZA8l2StS/w8PLl6S/8VRoBQZcivomAlKoTJf0hyrJ
wAlFdDN/S8AsSVAtzgiMu7uh+/XismK+FPB4J0HHZqpFm2CyhRh5/94MiJ/brlYh
9TMFL7jieK8+hAoaBl095iAjgpXcLEPD1n5EK+jr+me2yOKZwQnNNbbZcKrkfnrc
UeN1OrV8CxnTE4GRVejVdCOAo/ttiKYm+65LeXm2uVlhvSDq+EowaYxm+1oopS86
XExLSeKZ8+szY4ZwATSQf4U25ZFdwbd7I0VvCile9hf23AswSJI4touiwjjQlRG/
xnqvW6SKlXtg1h9UVZ9LXGPpfcg+sH1RgFrwGKnSWFVCAixfD183KXvqwoaHg5EC
e5WwD8rMIHlQBNB3TC6FsrvW6WD7/VhK5vIQ3c3Rbxi5TFPAGRsv5nVxJVPWq7h7
W8UmNPh9TDIBqNybeBeKL26LMvIAsW4hJN3WR2OGhQpCk8EZAs5GJ5MGn4Z8eZfV
t2u2pU2o97O7tVFIkbBqBK/3sRrLJg/P4lGO4FogNjKFcTqHBLZ7SyxWJsYDiKNv
E0K5woC9NNGQWy4mWXNEPNuvYe94sun2d+Wt+osCTWmGt1jSjqdIHVmlubFAKRPN
ofypxEvbVaKuo+ShJDFcoQco0bTquUNGBoxXZB1SoI5XVTn/BPV0w9whCRNL7GnG
mXK+QfXqesl6pLQ6VK7js7cnmB1vMd2kAWmNRh/pDrLC6OPMG+0aLabwutY9mZUS
hyQWVGj5ky9tugxdpvLnEJx7Eif4c5PXmjL29/QI4RieQGP02fUf582NyWnyoYXt
5YvSFucXjT4MSOvxapbGDbncqKQUZYxJFQ6NpEqbhVmtpFhyQuvm7crNm1TaiweS
IoPtayHNxjpN/OKxY6wFsD1C8JdSbSWNhSWzsmmPWzHaCnEdksfyOKMj5Dr36w8B
g29iC12E0sl8AT3hl//cTH4X2Rmqp6nyDO5f3OutmyCJihVY8GbLomlhcc/FuSKe
SeU04hPQy7dpIujIgIP5uk0c7BXM5VUUWOBvHggilEdWnrMonShRQ9Qek72VTWrW
5dEyfT1qiQpGb1K4Zvk5IEWlVeF0kkduCaYu6mdvgyw4LB0e2pcCJUDhZDUBHwtP
v3+3GShBObrkuHuyGAJvcIH+zPUaWVA33P32FjEhzSwnXM2qyKkLsVY2/KXaAEl3
BkuRhFT4BUgJbXHFXuDXI+t/yNVeEp/7IGAm5lbrCvjz/AE65oU23uwa6cRIFqfM
0WoN9SjQ9W1+tOcj9YFEO84Iq8LqoMizhYWjFVwkHuN2j1q0YFTcl2baQzrZ3kw+
ZJxc5dlX8lN9SU+BpnrCN79ULBR1EPYgq39M39gFZ64ZTQT5SoYZH6K4oM3+O/ym
U0f8laXAw7t/jLCYAj3rfGd8HGy3lA0IptO+PayOy68/sEo1wHQCnqy5OaPixoSn
0IkhApeLOYYZ2nBIXJn4D2UFEFYhysT7iBKW2Zks9BOY3DLSW2HsV8jmIFej55Dw
EX09jxlDsQlp8elQtxWeyUdAjMluGikgSOktJGfE7tO1eaapiOqWEpGTlhZzeBpE
bIKdRzfqijuPdRcBqc9E2zlDyv4YDj70UHd8yB0ru7BXDXFF57THyj3G0Csw10r2
u1MGrWkZQa58Sak/bfC6WvJoGF4DOG+Asb6pWNi46izU1QwacpTUl+enEQizNQ4C
Cw1trLxgMWH09YOlNoZqoE/9FyyBc0YoUfsvypnYpsR6ezUuXIGk06G9RoAwlj+z
us3lHydW6cEhSG8pPXsQZzlSPj5spkrrYq1fOG6EE0dU2z4qlkRZPxENugStNBab
5Ydkiwt429cp8eYTaIqVxCjKah49/DGlThwWVjfU66fZm4ap/K3Vj67aJ277QOCP
vuromsZ/NUhFW5prS2kqcjjMYxzSl5VkswKtJF2ItzIx0oQq0ktqU0thoocqjyhv
gmE2iz4xCqydiE0PXK9+Gvk7n6DHnt35+20UEm2WOnXkVghUBAy2KjN3K5mLggkG
LlVoyuMCobkU08Bv940N8gVcR7D3JLx+oHHmrdEFniFvlrzO4VRxLhccVASOg5QA
w5/ukkaFAZ0vZG0FtUjgHqY70IPeulwmOQXSbxnHneSXEm4qsimKT+t6wZJg6+Zf
64/e6YdX3vgGk6BRiZpKxkXlaoWZx9Ny8qCaUn7NBoUuWuuuUVYzz6x1k+mXMlj8
`protect END_PROTECTED
