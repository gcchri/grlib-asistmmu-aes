`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DW1P3FPoUWlIMjSjOKmp/Y+HUYaf/HBmdH4n1Pae5toIIU/uZ3Gtnqo4Voy3RPrZ
DPd3anH2Bmu4UA1TkTDBm1BXk1j7CI5lhTkiGzt4J32WYU8pbAPK53259dZ2gCs+
lHeqXtxojSvQbpAoUakJ073q2Qb7esc2tsF7Y5Ifbqw4Uh44WWQ8OCUqKKoBEBrJ
tGPkFtIcxXfbppoReutHgR1jUwmsMRGWiQJ1nWHbUjIUOJloiw6xdqXvcnd85vVw
NmdKlc+rqbmsNp/tzTv+8hJUyscOcP9Q2YPB0JwhnD4oUSvyCtV7GO7ILbwIeaA0
atsivQIguggK/+h9o3KgHFrWykqQm6LBlt6k0exD2kEdGGLEdNVWUg7Shc08gt5l
MxgSrNW287V1Iyn6blnGOA==
`protect END_PROTECTED
