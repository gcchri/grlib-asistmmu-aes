`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cx1XbvEMuevw5NXHyoDnvMFAqSG8kCQw7dP5/1UhiKdkJYPB8eAYItwMngfK2cXr
SS7xX1JozxnFeMHtP6z+sqLJaXo/h8ImTfLWstU8fReLITqu5x7Aku1XjHWC+uxY
3SrLOm0Mfep/KoNQ17NlD5ytuHAzJmyB9MFLgSaDuQENrP3kVVX284B1nc1gq1on
JMDyfp/oXvw2BMfkDpgKNpQVAj+tIEnOUkFaGHjWolHHGq14+AfFqPP0qHc0GSrK
NQlOnqXBCimVj3gzJeeAHI4CGFav3jMCGyYPWU4Z2PZlrdqiB5oGMXHxEFh08/tb
JWsF7xlduz49B+0rDLTLHA==
`protect END_PROTECTED
