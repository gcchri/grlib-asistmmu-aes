`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LOsh96LQEhaG6S8Z8+07biCkGo/1luVO71zZBbskHSwLlIrB6ZS/T4OJfAoYeQnr
515al5nRK71qomliqmVATZ6uiA9ve9w2bnA7sfl4+hJ4zVy6Y1qZg36PxQdoHihG
8JzFIBKjCY76z3AXfJSUCXmZZMvPyZdJ10bwEiK0y8HPV7mbY6zBbeaCfftS/1Zp
Lb8i0YjKWl4ppSe3NpgHhmUeFV1ppa/+OP6EjrUYQXsSx52TJtpQqzuhTix1Gwt9
VraoJPF9/84mAU2pAaKthQEI9YcOzqwycn3klMkZzYDwTESNLbHp69kSM4TPOUda
coFA5z+wFuJ09n5TjqzRlhM6Ltlq+xslgRzGusCRrPtusJhX5S8yYRzu5FHpHJn7
`protect END_PROTECTED
