`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fx6WTob9vfVGGIplxRBxEbxGHA08bWXPgHbllhXOOFJPKxqypfu5O2nWudQY+VDB
syo/Qhl/MP9hJHDKP1o5Q7FRg3Sbuh8JAoqSM00tC5J7DIQBke34jj7Sx2+++UWx
GO09aO664TUQNSfGI00WVyJPdrvwdNG2IU9VXn2+PByYIsH0cOfT+0OBPr+Re66V
qCHbJ4x19+Hl+FDhvez+YsLJYVXjOG2+FyeMfl23BgpKkD9fb8SXJ/4RvlxYNGBw
9GbPoLjYXn+D3/tpf8hCTUDJz5ZPmaKmLlPrh35Juu7hKrN4kh8IE77eyr/W3u5R
WD0GbrCgFOzCAXcqI6uDdA8zo5IS5QubQQkYSLdqBn5Vw1nY8/LWLKhqdkLjOrZo
LkrDiuniVhjep2WZgrAhbewo0XzonXxj2D4uG+tAFDpEebv6Pvi7cPRASa/VgZw3
nLHjpy2ckOhKXjC4g8Kgw5zGEEVM5BrX+TIba6A0vZtbQ4MmHFaoMGW45r1Bkp34
`protect END_PROTECTED
