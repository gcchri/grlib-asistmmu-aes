`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cq3WGBPukmj4r3aS5CznFrLovevnfwKKgguSe4Oaru7IArLWmmwbpbMPYXHu/4N0
T/RSWhxP3fozhF0HTcUc2853++0T9/nyfvmk2+l29kcLvsaPiTCeZ4aIBo1fNAYw
ZrAlX3DE+uDR41Qxnj0dvfNziz+PDMatr8cdeR0uCVAzCEeZtcLe+9bz5o5E4JD9
f8WlBPdH64Fdxtmiy43uNi+cMxsM1su1ZEHYheR9AXH6yeYOqbLGgkzEj7e8+sg9
`protect END_PROTECTED
