`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hHesiHwSiaDM5qHpk2rBXHiDbWH2h2XOYZx5NKFXa8LA/UBBbMk51sUe1LZ4tnUD
ayT+DBGe8++o3xP4ixwr8IY8llrXjabHWoBu3KY9pfnhvrh/7DoIfnWy3CkNeSex
G5UmrOyXuLQY9LYNCooMEr+76oRjXgdvoXG0oXNnHAdMscmX3AlJN1eXJEcb7hJc
6oFg20eXQE5qQ7zLh9/UDNJoc+x1SHf8BL3o7LiYeuttfVODCOXxEGBnnmAaWQ1y
tBgX+GjGDRYNjmp7Jb7LI56waCMQ0WsTOMwwPwpHvIvKqZMxFYsz/1AX4qQHw96W
o2OF0M+hQhp0riMEl5DMjmqRkE0BtVG7+QEZxwBTTSlrtAe7Kr8iQAFNxJBD0UJ1
e3LOO1nvbjQdBFQKNbXx1Mp7exU0hqG3b2ecXNkenBunwIhIEg27FaInD7+j6jz1
/SGdTO3LapQNx8EE4KINTDBWtQ2zMkr0GQb2QEsX8/B0oLLpEbzrUTct2RFAH0fj
+I7titRBIGlO8h2uTu7+AnMGJYJgCbeVuHh8aG9O79Ipshbpk2ILsXX3cCDiGRIG
S8irbM+aMuo8r7/+IlKH8/dUIO8gZnSLy2P/6tFNlvGQz1VTdeWZGOxEL0ZysBKK
uipv+OHG91/gMduU4LdElSCo/3JV/8whyOOBwasulDpsVtpvXTGBmtxTEvQKoQOo
+Avstj/tqPfYKlQ1rQ78IuVXwZsJPVN6XiW+iNjqm3HMQjSjfydCrcXKoGl8Pszw
wAmdNmUl9OSQOJpKiTfrYhvWHwuud9rcArgO5JkwXqhgyptvdPe8eR1Hy3u9mq0R
g4eR5NjlKpfwVQJziAtdm6HRToqh/Cf4AMiazZAuMoSQrLpRije+MwfQtfdj/SAB
Q30+KFSYDpUjI9BvtI7+W04NgcPHGThymRnIMq7pcmg/yk9sTKXxxiqcBPtCNZd4
MVabJLADUIljhG2R3FFn/RqhgmJbTLNHe8aC6yE5aSC7GPBj1w7K3YiKl7fNbSEr
HUEW/Gcljoes9hwcV17IbGm4e6WL/agE3vLbI4AjR6zxR7IGy+AEw1rLIaVEQeJa
QCqR+jPArtd6MMSZlIfNbdRJpDz3Q0BZySA/9kEdt7aMRtw+g1AWxadHTiyCmusO
3lZgdUDXk6ePSPbHjx/l2e3rhGu/ovijmt3LALg8kBp8jDP0XAHbfb3AmLZ1HC6P
2yyEKIUNU06n/4fsLgH2B7HYVk4s5I8Bvf+hZL9ml0FUQQhSwf1Psp0u+WE7WfwM
hMXRvFL5KPnTq0NAmvh1hJQ+VPEGqv4oXXIHXOX1jIn1jvb7/XB5RU+hZlgrqmId
ERd71UfysoDO0EinAnKjsqXs4yt+htlS92A151NcjqCm3SrGnDDLGhXg7oZZ7dpH
eOVKAZbiGnSSskE6FUGsRmwNVBz72eL85rE5oh3gpHOTZta0/1pzEkwzWG4L77q1
7nmjyPCQygbxyl4XHPLq/ZO5wo1OltIpnsUT0/rjaZ+a5wpnaaYAGXDW4uz5eQdo
+WFpw9lq6Z7cNo83U9p6bFCXC1MGp1h6WCvN1VevknZUTp76YbSQwHicxxGY/YXF
3REDcgpzBveisy60VeNISY5HQm7R9R54Bdj+sKK3I5+4MEcgibvEzbpQMBr7NSVd
BTunNFZPzw9DM8Fm/CnMNlyCPXBFsRNCryXdj4bEH5PbUV/kF0SVIpey2pNyeW+V
TRd/VnaoDUYielHWTge70o8vSxAOymIYWbzxcUbEhLnraRlagQJQeDAHBUoLBfck
mxfgC3tTeHyNwgybU+1opYGfEm9FDEtB7beXcW9qcdEsZrLC3/vbSvSj8Jko1LkR
83mEGBDc3PAB+sXjnU1TTmS/IL+VkTdhd9fzI/WiHHQc2n2ifRL7ttGfM+VgH78v
Z/RhS2OxO0o7VjXHiN7rfb23spS6/5nVpXHGT9dJqPGJ5zWirZMIgpU/EdQSfrrP
b5LJtSTXTK+Smg1rLOR/rKl+boCZgBY72bKclzJPYLnC/YEtEn/DgUJwmW0QIPoz
CTWTqxR3xnXC7PDFcDg4ONPeQ2GUXv2KJ4shSRJyE/hSqBJB4P81r9ijDpivZVRx
uiffJYXp206QTM3VvjL63ivcbMqdeC7QcfJLZ83L88y4j6dKcWumSbU6JU7KjKbU
SzDsnJS6Hv2umzEfCT//jRfh1i/glukhRMXAO97VWVsJZrgOZoKYdfruUGmatcmh
48lC3/5TPwElyd3axkwaLqbW43L1uNzZmMKgRRojLdMTQ+Ay++JsWYmhK5rIXoQl
CZqku3kec4MXUT5m4iwzy95w0JGYu8JwvGYaLlBcrcNxq05HNaYg7kWA14Eljn6f
2wsT7ePB5L+i8qVMeNgG2DYaqyHqFjK+AedZSJgwIqirtDukJBS85TzRpVXYlpYY
N1sS+QL4P5bn3DzHvSoWg7EbA4Gh25dNIGGIIwf4+YHS3OMRHRVEM5QbMs2EIX6L
efeBAnNj/UKMLq7Ia0QVOdfHHyNUW0RqtNXD2mMPzzlhklMcEwu8xvSu4wAiAeOb
WB9U06PkPexyo5wqdvYvMFKbETetUOCk7k/cfI315C3+oLnW4V/W0rOpYnJxPiUm
fz57fcwtBgvU1m5Woi/dko9zd53MmoZN2gZQuu3vDWl6BEOlwbTMRgwQ4xbr2g59
d16vwXrRcl4uDo/3oN8lP971G5cCvOJvbEL9qviGHq3O0FsFjxOb393bH/XjECN8
y+48HuGlnuwW+cktazLefSrWY4lE2NuXEyDKRviHs0DdS/18VzUbgX/TLddBYj0y
/9Z1Yl4uVojoohQnZYpAQB1jyyTcI20F97ovrMW4wOwx/bgZm2I7wghL/nmkVH7m
BL68nCW+1UlCpWEaF2UKu8y8LxJngq+nF/+o3pGhP5jYuN1Yy9C62oG8MOUuXa7x
w+Swv+/XNZyad3PMEPE8KyH7ETIBai95YM+g/LP8u3HJ8AU56HARxAo4YQI+kj7E
elMLtmjYRSvVJ+IMwzwqLXeqhyFzU/D87Xm68LMJaxjOOhLSwWU4fsCzVGrE7smL
PldNf0eZ5l4N0Npq4DbkOSbkZG02NK83E5CzvkRCJS3WVBjR3LBbNp6avqWtW5yD
FjUOL2sx8TRjtj7V6V4/nLh4aJx/lgEewZNVYsqAbu3H7b3sfjdcjc9KYABK1ljF
IfeCJt52E1B3rGVMN3KWb2tOWRU4nNXi0YPrvSPfuU94rZ6RuvtSQiK67NiBuB3s
DFFY7RG3A1HV/J/YkKLuSW5XRvcrhXWB9nIPwlCJIXDX24IRH8V8mV1kq1JJEEdK
YXva4v1pcA7jamIDdEG2bCPQIqzzDorBuGqe2DgDb9qhG/HeVH9sxfsmqsTQFruR
HQpe5hK9U3MV4LzAVTBNreTTnsXcdK8W0CbqTIhrqEwdeAROxPSfZdwH9JSH9Z2r
25Epx7x391dqKUKkzGL4fwcDRrIt0zfqTPbu+p1iqaEhvFjDp0eeGXJHvvZuTJA8
L7ylP2V2r3RujFVmc4t5IzKpYEIJZPCq2dIaJbQnQgriyfXCVnZ5/AIpskdUrwYp
sF9U+AApQ9xSNFKCuoRQwqtntYhZQfvRO1GvVmLxrf36QrQk50Y+2aIEKsIVqZZB
`protect END_PROTECTED
