`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y7NsJ7y5/qM6ESPZXgZ6ICQt28JNhIzmwNf/6uQTyG1ocLdlMNbsnYlv85BfxOIh
wvdpWRBnVY/sV9h4rUbDjqrmfZmOEkfdVNlr/vMyD0CQdf2tF65tuT/7uE0HdpIo
UVr/OS7NbiMWiqubaU1ew3ucXadDz6i2LUoF95Dm5CBTtPcmtHQLmsWtqu7qAjH7
eBykoP1N13+59dj0QnxgKka3+/uRsymPqRDIWdwiM/n6z/0XYJ6JEV7RI6HPkcLJ
IHwmwp4wCzJDxyLVcSD7BPp1Nh8rbcaZSYTrcgfv57EMeREG+YZBKr/51MUvuyE4
bDNppD+GkGTJZxYeDSv95jVD2bvngIJVBGYQXpmIukKNmKvanNdX0TcRPru3hDbn
UrQJwatA1kSGWXG82eP1t0uwhF8JBhmr5+Hr+h7Y9p0Q9XHEj6XzZI3WH0q4Opo/
zW2Q7mJRSRQoKEBiUbNk10gu+4RZvkEoBSb0EJvtWETFX14iJce9Z8MdbMNYP2hv
`protect END_PROTECTED
