`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ag1HkDFnKgbjVPA8yXcVj2zs0HJa2CLBF351N0d763FYKVcS0RNoJCrJmTbFm36y
auLIwnJlplcYkY3Kr8IoOp1Tfcr3bNctFdnDLXqo6PoM6s5aAhSgCeCtlfS9TO78
ciG8OAsjefn2SuwuY7ZoiGwjpmGF8BGnTHnosdcrYWvNHX32qS8ytNG5QDRzZp0J
V+ziUN+fROtVFCfcFvkps+p5SL8ABk8Y3SkImbZbEbSv4W1BNhl/8Db7bwqs88sk
Tu33S/G0ELNxutEkMq/l/bBVe9VJ0QIEOaHFlEbeFhogqmCCuEt0YaIG91b2WIxF
bits1KcnzTJjiJdGtToUPxM/KXQ4QhbO3SOAAInc7tzYA9gncuhWQUSgeYOBQmR+
y0Dr4bjOQhbyS5NaytHCEcmuAQY7pFh2Ozf0FL2JkNAxJ0yVvTwnH5Te+BcOme0o
pKHzMem7DfFWzIgUqStbVpYuaQ9ZEZqfDk37WnZBB0AOd8A7Y4r3ozm7ie/langd
abHkv6KUjTWlbzCxQxjPg0u6m++LixmqbVxQBtJ3axDhxn6ICcjlTpk2B8IR3+cw
h02yuD9rwYgRX8KVAUnRAcwYFr8v3Uh58v0dpV9rRCgKWiO0uPYphejsVSpO/RtU
YmEiNytEMYP1yZ1fSCFtyWBYI7BG/ETCP0hzu7NTgC7uA0bSuJP40V63rGPntPy7
`protect END_PROTECTED
