`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IssmZHeJa1aHoRWaXh5OZHSt7nXIQRPFbp2S4kbUSlKud3IYwalmr4Vv8wj8+TTT
YSGhi+N9ANPRBT4jcLI6c/HUKTRIwRHpeXmL+6xBe6ZATXkYBjX2qbb2J0S8GDxw
Yl+HuNZEnQjSdFCd549D6jziKuo4weOlDh7A44Wdzsul3mBNlA7qJHBSaWTPwUMY
TazWaxfjdYhs4XN6SXIcA3yKyBx/7WV2rs2eipx3vk3rqpaEcioWxkynDF6wFGBk
MxxR1Nrjtc2SIA/muodKm7mz+uC3cOutHiI7I/MoZQnGx/vQWKo5qTLBE1GDGAEe
wrV1l64dC7tEDjhiD8/4IoZqKIWjjLE6uZUDown/76a6vzcALzB87e9b2MJ3HLQt
k/pdAwMgzhuyNWfYR5JaSg==
`protect END_PROTECTED
