`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0pKRp6rxRdF8R0UmxJz+BR/JwouJCpGegXc2oHlB8XT4KyqO0U3suTTVXWiOs7hb
z9aaJgc3f26n04z+Rt0cWaQAeIy6GuIcBT/1apIaom+Eu+HDN4M9zwOZjCRDgJDD
N1hyDCuIB2j/XOdBUjiZurqWT0Ym3ioB9EQ4lo/3q3H9IKJHxj7SQVL0a6+239m1
GxCoVU4BiOYpa6192fzFzsAZpoFCJ5uUgfF2Atc8OutmPPBxIq/iYBh8alONEjDa
9iuJCNeOjVzYBnswn2x8JgbCcoumT4X3J0g5qgLcRiXoT0H+eh5NQAzV2Ug0KUEk
VoS89DzbB4OXu0J1N8088A==
`protect END_PROTECTED
