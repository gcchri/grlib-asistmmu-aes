`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mJwrCCp7/6xvqfrRgb8fTg4H1alOUAs2dw2KbS/AHReqzsj97VXcuHK1fK2au83l
SkD77tOCu03n3+/kUpxs9IfKUxJMgnMkARzetty7LpLxgDmS3pDpMbujdC8xBZWr
3XoNfBkH6EokwAedwrSaNVZm65FSuA//wNSp00nkF1U8xP6N6AkbWOk003qvnQbS
J8ATjq7yQ01zNzLQhuW3A/9KQe235K7WbmkvjuFyJ7vC9gP60HB2PkvIMt6giFEb
QXoa4AMVgDhVDbtsXMRNUuMupH/yPH1mLv3BueFX4Mulp34WutrmznPcC8FTA2Nl
uqINDWSIe3j1lPOZTrB8pYQ8UR2NTbAboVBkdqb+BPXSxFJL7EsMDFgdH1+zL8oi
RR1/3WlxuWnKiyGCHK4159nN2EHuH57vJ5yTCO8zZj5tWXeJmEwXHp9pe25K6034
5HreL2Vgcgqaxy/FSHcvwfP3E+KjSD5urf2+Wk/oyQkBNh9N6Lc9Hhrd4Vba0onX
8tb1NaI2Jo0vjQJTFb9oLJXtgh2qdeaj2n88rqLT8E6ih/rjrPldC5MHgxHQm6VW
98mZinL4fzrSvc7sbocUo/OR6WZ84butDNhxPOTcIxmDctAulm7rsoUC8rupDXpq
Fl4evn4NwCNETwA1RkfmBEk0kL3F9gz8osD4NlEhLbzCh31e6f/K3xJvLl2vjf6X
mzAOWhgy9MLzEnMFUmYdFakVvnhzPip6yxn2mxcBIOHp5RrA4YzDT9I1T4FqbySu
oT2kIj/l1ZLJ50f6RZULcqq/0yCWNphLDqScHOlX09Nj5okTlagC2nGh6W0gtr28
rMh0lvPBmBnxe7jwFUJjzOEcum+eFM5HS3Ams0Jgj8jt5Sq5tNhla82WZ0mnpQVR
YOU/phWMGgBn7XR2DBOm/CY/VsE8Wzdc64ukiQjo+87nyjtM4mqXedSPQ4bTTOPb
ELemByPHoGEU2IH/Qrn7GbJnpDa5Cfk5ijHvZjaodan3+RKycTC05YY9a7RHaZhK
zRoMEXP9hnAzKqH4JHu3YS3WJ+stbvJ+o4oOqXohcFGC9mmCvsrPYL/Yrx4F0O21
H7EwbtKXYhfDyQZ7wE/47NLo0CvNaDWoKe3GdxuFDu8as7f6kPkzk7HjkyLOkwmt
dE7K/7K7gi2DupSwQT/UOW81X4mMdW4A7agylUikcV6SdOehcDAucKjSRK0a2P3m
0riBAA6N1AhqlJhMsmBt1h7eph9W0sDf93VzW1QMD5Rk1RFRj02xNFe/U9KdBNKu
6yiAT2OVp3U/e1ZljX48chpf3YSunFy47Bi5jYbMWDJ+YdlyVRzDHLyIE86TpW3u
aqZQn87C1cQWz0eyswh9qda2bWs8pK3QAq+5c/t1JGe11X3YAvxGhbEgI1wgLEvm
FbyIWWF2sfirLCeu7A2ON5cDbGleCdtJxiTUJYQ3pJTnaRy30SSFL9FSiKTqYXmk
oy8k6EhpUjRNMV+TcFcs9IcfvpYFJLARMRQyydJKhlVMok/ZIUNOot8Ip0Qp3NqE
irI8E+lcOjmrNHngqJqdPFEI2YvUMootmKI6vw268eqRQiZNhS52TD2mmQ6Vcaqi
LmZ2uTkxUarEfCZopg6k77YuUlbveYGcvUnGpmc2DJixaMdSbFm9fXNKhi4gh2el
f6JAQtKlv5wUab9aExd63ddo7L0vHrr5fGTP20xv29nO0sRkfnh4mBfElBbD2/zf
NEU4jF2Cp7O/0MgU/3JSzA==
`protect END_PROTECTED
