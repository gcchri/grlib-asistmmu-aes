`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
56zVHMsRpio/Cmr1p+GO8sQJ58Qcnza3C5TeS3Sk59ZmCn5aQ0TXeVMFhVIuKhqh
Pw5ln20+PPJx23zHJbmPBMDhwzPh4J5BaSp8YhS2ZBVEFrJ7uwsiovAmykeYAzRf
VMPV+sGBtbaIjpGLetbRfZndEPhxkccLoxrz0PEJdk+9HMQSThnrdhIkgKvGe19z
1kI2jNmHUa0o02ATgxnf4izbIxnUt3XfoEaZTuRQ2KdrifjxjY/4CBGk9cHuodl4
R6BYmrbV9KqtnAEBhJYdhgScG3ul2gnawbuMv5Hg71+PIMMt4dqCCzmKM84KEZDc
pvi8v1zXq6exawCbfRmKaRoC3AwzcWAgBCvHPZbezjFzXmnpvUAYhHVVJV4/hiBD
pLZhE7BswllfD6ldDfNYytm/VSQrHYX5GoDTCyfKJ3SYh+14K0QBS2m+xnu5HkHy
Z8G5Pcitfc8Pq8t0FrhW+Q36dK/Nq0HJsJFCAzLNqDk=
`protect END_PROTECTED
