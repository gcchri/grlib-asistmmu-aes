`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EQdEOExtEffpStxVs/5zjfB7AY4YZxgV8dbHbdUhk2mJWMxLavYqJSLlSjgATMMQ
oLWhrayqmD7WevIHbVgqXvzWv2BjOoZMOEeRSvIUjBRSCr1w743r1xsvs8KuyjY4
P/v8ETl5zJk4f08TNgi+BxxTbilKfHe14BsOfb63Svy99JU+zb+B7WhdFQs2GHQk
hYtiv3e5vy8OuddeS8NogO9dmfDF6V5NWCTtWPCDYrohUlHC7V5aipCLkUfkX+YC
oW/t+fCpF4TSyc7mw8w0okQSQxP34uxXeteN4q0TUNs=
`protect END_PROTECTED
