`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wTWN5T8+zLKjbPPVGmeUxrq5S0YB307P1EgtH4y5LT9f5gA+OQxYOXRgM5dcbYxf
+Pzp5SpX/lcEAEuvBFp5gDaoEgzSkN7HS+n+3ypiAf4NEsP9l4kIUsIlMfhR9dae
PchqpuMiom3f1ae10SRHGdUDV7oHzYx+2kaBaTe7nuSQ7XLfviGeDS+0fbRuENN5
NMW/n/dKa93zutVxB/Gc40u2k4Ex+zE+DSRpTgilmRNzS7LuTzZm/TsgkrQuqw0j
5HSWL+K3UOKudYk1i/Qfkg0IWDgp5H1Z4qJxC1xVcFDcdIoAuoOCmnkSf8mjVY3Z
Bud5RZvCAMaW9pLZE4audg==
`protect END_PROTECTED
