`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mZ8nNgeVEH4L2t/79pDtQ4aTLRjLeFCRFPgW1iqLFxsh+f8cot9oxpicVeGLWOGT
Enitlc3T6SqX5vVaWCgeSy5FZJgKhpQEfuZopumf9/AtaMw0azhVtTn+crPqoeUA
geIKeEMlJozevPSTUnTFhnSSAbqf8Pzc7TSo6riSBdYKAqKSK/GSkOJds1MNVoUX
u3WRx5Dvbg9QfkjbyeJsQ3jkj1tmULIjezej+Nmw/OEV/jmxG05htKPe1IDyfP+G
PRn+1YWoqaaZbOKQUSWrllHkjcv6jdl6LjpmmlAZSXCaVMzJEiwcTPxJEXqhoQE/
FycuhKw7olY25tCb8KiKev61Ptah3ebEF63vCOrTll3WuqygIOo9hS7r9woARvIa
AUnGn8tWfl8w/81lc5EEDbcDF1XWoF/RfLq08GOYeOzSKUI8shm8sXdx4KZek730
w97k22rYjujGBC1OYqjRnYA061kuqbSfd35OQ3Uf4VM0+A1wGzSU53mjwwYu4ZKm
mErK4Uva+CbYGgcVEk+ZPXijsE0J96ka8gzQ6mllonrOBi7P9Mk3/IHRfVVrtPpY
yR1cqyzYG6iakV4s044/a7q/eESiv/AdFnlHoBNlXLo=
`protect END_PROTECTED
