`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E+1vl3/sEkcapfyEfjhbax1d6EWM4eiw2x/aQ5Qsoy1UR07DetVhAeOC8RBHWUg4
aPEGxdHarlmEvCBEmQ7ISTMrW7o9XSpfAOvtCudln8AE9u6u8UNApwPb8esjwTg3
wt9J834zejWaSJKc6UvqazpmhrABoxBKquexnINe54Ag6uqLFHuGVvUQcyASOcAN
J/v8O6+/zzTZeBslSsmpKB3nKvL3Jg2cbQLhEtS0jXFyTSsSXGGzeaM0MaxtToZ8
XCGl/8fw6b71mT42l6UY8g==
`protect END_PROTECTED
