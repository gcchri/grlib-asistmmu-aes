`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
463W2jES327DQsQiGOD7h5Acgiheia/GK7SgR4Oa7eg4WJJpY2LTJO+5sIC1HAcG
vruESmpD+lUa9+WBxE5Et0a+6l6SWh3jzpCJCHUR2/ZLYzyhHKlX0ws3NKf+NdCN
iXHl7IT4f9P2z/6WnLnyglRMRbl9h3u9SiRyHPDh5tabwUCL/id/j8L/7+DLDHUB
R4i595izKk+N20nCIkUx917+1YPLg2yojwGnBo7KmmLzErTET90nsFupf3EB8sDz
bUNWQVJDBRBpZFBBY8YoOOUQJ6B536zONyzszCMgXJDQ9iXDRsG0gKLxJXVFjF6J
1OG+Twbr9hxnz3NklNDtRUeK18p/Fb9AY7FnWqLvckzjsCzQ4A5UK0fs+ueIKpUs
69S/vUtzxACpRUIQiYnxRfdAU+vyDCFCMtGZdPcBLHs4rp39dmVQ7HfhCuc788OD
pDJaNvxoppYnn/ejYgghGR3QDrEKFR4pQUFE/fNLR33qv1pB3y59sWoM9LaKH13Z
HuJzSBASWLgcqM+xYvrMGrwOF6xdTVeuEUVdn2yzF+qruQcRPo9BJtcNKwUTFZ+X
iBH9OxBOo/IJG1UghiJiM29NEgx03XiygJ5lmuLzIYCvuN5u1LMUs4uJKgsA03Yg
9dP5O/YCW9a9NxGf7m2rCy2rqEnE2slYpzmBcKc7zKEgQIr15V1uff+GAm/dCli2
4SnwEMiXV7L7wbjND5+zFl8ubvWBLAyLQEuwy5z66Dk5mvO1IMwebniczn+Yhn87
a8n9q//xqfeOcdov73gdTNb+A+by+jrUv/15p6vnKHXv0ouLnq+v420YLByN5qV9
Fb3tOhEYuULprVF2g5DMS7Jsc/tMPhcn6Sj1uMc4Losz69nFI88mDauVPl1hRkc3
Vfx4u3NtjHJBlwjewrcWwUWkkuqUT8wPmPw3ItB5JuSKUGlKMeNQTcaRS5Pm2/9P
IntCIv3KRWvqercehM5KPp8GBHKLUO8NA0UqBvIjeXm4N3GWzN5flKN8km3U5t00
s9ZUsE3P/ebEAjaZobwYmbJik1JBGQfXtPATSh7cg/PrNWqZDVEQHKzIzT4F1WgN
NEg5ANhlMSdWEImDTdVfhj8IUKWhhJNqmBS9uULyakwnLNrvFDSSQKJakkEyQ36D
Xg5gjZrCqnNqjbwKbHSt6JX8zfczCZ5FgxWBo425kkr9OREjRhVdOyfqbMrtgiht
Dp0EXMQtsUB9mDPtw4J0dle2ccQ6soUErUcp/OUEfbLbpfhNiGQag94kwSs5OD7n
3nfAfPRzlZCd9Ci/YCnTT+otJq214YarSvmxR7GvT/qY3eBPjt3DUZGrWZFnvmqc
mo6/Uj80qM5e5J0jk7vPr1+eZ0DnYXPCuJHgUMNMrQu/YdLk9ai2nZ6YCcWXUjyG
uZhwyIMVWC8rdv8vq+dGviPpwVrPTAGRObAwJ1s/xF8Xm9JdXrVHTbuNFojE63+1
u6dkJPMRZggp5APLGbJ5tSGk33n5yp9TgvekfzxFS1JGA3LTpEzXVarrBOyh0CkM
GFyPpgruYiYBqZn46lfe+EFMk/Xsj5uTM5nPOI42tED0o9JwB6bAyfiiwpR0hNab
/lsnlsy/sIcxosRK8/SHQLxSf0mov2ioETc7qmlxsemv05VNGcX6bQu1ZweOtzI+
P8tItSoyzQeFPOYiA2siZ7N+3se0g4TyO+TN+vom38lJU0yaqgY1F3fPGYjytveA
TMWgnsaKvdUhqGzJAo1SW7w6chn+7cHTjrndirUoLFZ2sBmHUQ7CDKT0iEyvauLk
xt7BCHldIQAgMTDghAb6mRIk+2w++ibik/px6NOp+6PwAlARH0JD7z+xg4a7HtaT
2LnWZbtdgRrwljZivWW8wFs6HwI873GTVzqLsF6CEf+38n8Sxwz5R4S4CxSOrMym
5QstwugsvNJPKP9f1fBYqm63G89di8R4cq1RML1TOOOx9jorlQZ3nvDG9n2sUlQd
MyxC4SbLL7YqG9yVmQDnTerKSFU7YA6BGXU1EwHuekkg+6ApAtyR0+Wh8aftN804
U0fg7ywqGfVGu7qMl+Y8aE6g/SA+byi0sUCGGDDk/aoeLMG08EMDUZ5sJ2Ivh6Id
sFtKyXZzFoZzRgIsC4Tx5n86L1UdbOsI1r0M6Sog8gijWFVrHRbrMDnQqkJQVt/Q
OJ66NEOol0FqIkKSGNwErFqfvQKYLUHXB394afkoyW7NmgwfkGahFQbeAnr5naD7
RVv88Mt2+OOYSjiEmu29nf8vszArfGzBKxMeQlCzgqhq8v52HbyofY/Rfb+7O0BR
az8C/5X+khbSlwZHDyzRCmB2ONGOuXHOjsPdg99yixKPVC/J7f138F5G+jfbZ3nG
4CwCYydAtHdmcQxvmgYM0fViqcBdmQ5jqHLFTTU2OIa27SEAAhHAf06cY634viwv
koQv8o/m7CwLCnWVJLyVwceT/dy9dV+Ghb55nWDhk/qXMegDKaeJDuxMDYD6GN1y
2ug3INZKIs1EP7PUe9vK+C7noOCWzHep0znIo1oegdyzXNsqORURalsS8B1kDb+m
Hz9eDuS8xiTXMCk9EIdpZqSJ3mjONqnP16r1ETm0ruYFDRBC+MtgqJET2YLizkyJ
thHeuz5zEqzNwlLmTVCL9892av2JwAnLKs1iw38rwFG+1LwX63blSr/+sqT0kBeU
jlhVV+ANbR4b5vx2eySMLvXAERWiSxOYjzeK1UqHNz21LZEcgH088ylcm5GoYlNV
AM4uJMv5kxYFeLr8XeTII1a48IcTIjVIkFdBD3oV2SfTQ3ib7I23HdFuztC/i563
Q2O9OsaElg0To+xW7XybOsJRCoBxt/aAuccoJKZe8iTLOcKTQK8u6LgYI3Zz0BxL
Xd9o41giEVC520J40CU+9bGauwqAd7RUYMpAwUBazzoM1cwPxetf0QpTPxSEZ1Li
Q4LuKz3DpVhqienHXi/s4ViwWZYX3SttBfNQuxCoPU3D4ynnX20MfJxa8LKxClZN
qdwNhB2VN1h4Wq5qml5JaB13OazT5hxvPpe34riUfWh78+zNHdJl4ISsJcAIKNV/
bSdXC7LKofvx+tu6SOZSu8Mp7F/Q4OCUrcVm3zYpCFv/Bg3v1J/K0iLern5kqaxM
cfKRVKIrZ6ri+tbbEPKmg6S9GubGFQhWmgwkc35Qc689F00CgI9zBU0voDvpuPCt
MFAsPcXOL5SEM5wEm8Vq4omBY7WgZDmmpY6FX38syA76ZFQBzVh04EUTUad3W4hh
EQn0MRnGVbn+dFl09j0VjQHZwoGxbtJLXN6fAKnkQXo/U9YNqSlA+1l0tudUVQXX
9Q2G9EWGdbjHEGfXfEW6gNs/+hoK2dqiQfN2Wl80g3eLentxXm5DNjhZjxGn+oE0
+raUQMga/IQQybgKUUCeO9DRCdxZW/JrPJ/ZuCkFkGt/bbJSI5RHFCOngh564/1F
joXV9aU0AjqUeLDcJQJTV3bQLNZmuysg9MWkPwVzj7+h5WZIO6XqkuIjTzScowMA
THs4difj8Vbo5LFv/qmFn+ksnOhhZwUNL/X4DCcq1BOmmArcMhIBzIO/dDpt4kDr
LVgpoSRD48Loiaqn8o/UV+K+3wo2W6I9j24UrHjW4aOwq6UNc8RjBl+Cr0Mqpv40
23NJSDoCX87MU1g2gx3AJ6mEXHTuJwha3TCj/Ip6Y+I3eVWRVX/us4EqMs0ydH6U
9YG2IkrNIN3xUlkTUpSs4wj9HopHSNsTzgvooUigRRPAiym1HMgTSkfCBf5owoi6
fmuKffYGLV98wM9LeSiCxQ7QHffQbSPcYMm0S/cFs1CIDiEm2KuMSQbNhAQe6j5Q
GRDL0+MIkDDtoSPhjp556S3ON1tGcfw6z8nptgvIjFl3R70oGzuAKc88Fz85d78+
j6JPRVSl8nR7dLKztnr50A2yhRD+vGMZGPgac+eI4YD6kzdQZmumMcMHHYbB4o1H
Bjfkl5YEydKCAEnbKkQKRoJ4eXbLdeXZIj01PLB5g3nM76LD6iBHpsth+AZDm2Pq
ngN+uWPL195Ha8420MCXkqsNv2ZeKp0LVlFoyMutQUZffHaP93QAfYzBP6qq54bD
/G0fU/3pGVIudnjaWDMMs//5FK5ZfwmOR630dr0EdvOZ/XYc52hXvEqgQwwPeGiB
XKDPvGwBevueOKrEoQnMF1Zgz1o6kiWE+HAx0jj0nPTVNoX+FGsqEhWOAy+Pi6Ld
mWUunSCWeuBhAUQbYuYGFG5XDn0igo1WepUHuiyuNtftAIRHkJgG7g/fTZuVc6t6
iIecNT0JlfDuVOqOogSWiVUIzGP+ZYfzqIsOYVHOHkb8c9U/xHH0KMjZgqVI+p9d
wyVrdzjvihlxf+k+lJNJYQdJFj+Z7wuMVuOTrK5UNTDGitu2oGAqGdqVMKd5bOtm
YvT/RMqbM/cGG89KQKBewxIZ3zvZDnu7Lqd+UHixe33n3nyGUPOzhhke8M7uxGmH
/RQpDplV4plItU2UI3+P6+OnancWqXpgvN8mICItTlm+RNs5ThrAuP0O6q+1AzkQ
iKvJ+u9McErnpZNhiONXOP7ZefagqJJX+1NNwDWUErxeVXoigy/SWPeQMWeCWazy
SWUnw4R2Yu7g83+tybD9t7TeTZFmUhMcstG00vhrxQK3wQNyb02eGk+9EYqKQJ9r
ikwzjcr5vFXY989YW095LAAP5frWeEs+LLGVDKfkApPH3davTGYNYuWRRkpMfa8A
D7a07Crfy/iaJaSLe4Wmx4J1FRDKuwz75iedFB6Srx4VkEBG2r/jPoyPN4HxODOF
u7xc0TbJAZLT0vdEgEWnKmCRRystu3Qcwkn/tjIgNZuodPPjIXZOpDrlbs/5A6x0
zMcXC91MqF8dkCKb89NvePBDP0RQDqkslO6XYyuS0b4lB01+yT61uhpt/pL+5kHH
zLAYEYPKfuagVqPDPkaPbfaXt2/dHwN1p68ba5+IMfE=
`protect END_PROTECTED
