`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y2HsaSqE0IoSNQulfzhXZs2BPcr9uF1WBho0oZ/3ggvq26e57wcNfb3KlqsKHW77
On5SSlC1v1rudRwhl+AlM7yZdPoC0OAzj+2Hlbi7LX+qzp2VyiChG8OHJLzOJReY
MF8QuxSu+nceyjASonrDHSANs/jG59JYcP9zTc9RzoyiO6Ft3RLHbGujKhPJx71C
NHHmb/7nwYYrbZgJgHHM5qsCnoCu14KqQ8E5dMN+wkERkYolNpSwTc3cVMcY3UII
T/x3slKrcEabiAPRbX1Jx3sQFyHX+j428TFbpt60VTm4MWIe06OS0kM5d0Xeg/es
7YWNuMPI1qB54m9jrxSo3Y8fMdf5+2tSdsTTWA3GErcXIzb/9peKfycr9VRJ8y6K
QolYD9SputtdBelDvVNl9SXNDvvxI+uWN4kREZXfvVSSGk0cWsNnJ29VI/UZ+kbL
N7nJNnRnnTtYlEfq+lVY0HyMxHdVZzNfanCChKaMKrFrKtx2gRFSd41g5LDULdR1
tEtWD6EMB8KkYPNLybHE5r7okHqzOqmVAoIx+PhgFgFqqKHriZOfSf2HKPyoB1Wr
89ZoS2bLEDpvrZSU8T5jBNz9dhLHPnlRjknMf7/AKSsgma0CwIjSkOSJqHPC2031
GOBw4lAkyH2NCtu2lcxuzgzP5jsxisMtL/e1WCgBkz7nFkBVPl1PJB44xYk2V+lk
MMC0XN4sUf3RE7jhNOSbrrs/ERUNYq8nRg+YfLe4RS1mSNumCebp2Cb7fk7G/DMM
swkzaQ0wlhZeIZrqZllb7Y1WoJ6fl6XldtErqBgR+VKDe0UPseuUp34Avv576Lkb
u7mC6YDQaVOoI6DQvdvi1QE7C4GhwTPw3JxJ/YZzkNvmCJuZcRZJ/ghTNrig8+Fo
JVQWs9kfXnfcGboxQ06MywAJntylt8TcOOzQ22d/lWxKJV4JmRA/X/ndljNEXVXn
yw6IYghThO8qjKurWmQ7A2bTESKK4qW/3Ot1P0CWkRcjPfWctl7v+4D/5NA8GtMD
Fumgof94CmxQF6TAZnuqhlwgVseIENGBKTEOgcq894unwsSIGm3KSUp+P8rZFq3p
tM6MFedaunUoM+Kv5zCfR80xIjBy6Q33nxwcf1E+Y5lKI5H1FY2/IdXGI7tcUCSq
K5R4A5cqQQ1BrBaD+IRcg/ijdSBNncEIBogZrgNAjYxRsRYrZIEje3eMBkmXoken
QwBGw/j0o2jQT3DMULEysmyMSAmBuZyVau3uBg1Ke4vmpUC8deaksvtBcpWZjAxA
3feUJkrIFIiB7Qc8KgAximQ/Z7CGEvkQJj8CMzeHJZUofTzSpc6j/NiwTD8xjyet
ic2oqip1bY87cW0yB2+LaOVXK/PaaXsjXjR74IcNKED7nsZY+qNYm609mkfIPMcd
U3iE1i0b1N3I8w/hpZyXKW6jEhZXcqkdHbk85GmkvpK/Rn1HsyJCFYdzA4Q/opJC
3Opcs4wnIlTT8bnoOF2ktifwdrEo3139QZVxvn4tnw0=
`protect END_PROTECTED
