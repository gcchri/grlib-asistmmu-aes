`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1v1KwanHuRorMDnLLLMQ8ev/cX/57sYxZyk8VoAp4yRZkRvvD+IUPSYCCzXRdoZ1
kk1MWNTcDO0GsSQtv7JRAQT6KeBywKRVPRRKcAw6KQbptG0sycNiWM1wE5+XIDIy
K6V1c3qZ+x/tF3oT2kKUKuSLfhPvJSArHTx+Yc/JSI1TLyBwTEJZH8q1O+j5lfvw
L3xvzoWKwrCNL20xoiYJkMFTQNVnNvXpeXBKuKRL0BXodjLnrY1+X3Yzn5/TAu+Y
pViYgicaGYXzkRASLV28U+8raeBrnSsAVlOilubmxfwRaJib33KNh6BKZDAdVs1B
fceHlIEy6jgzsGFkoXPTCICQFTdZlOgSwonVLvUbJO7RIhxeJKpKIRlqT7RvyBzs
GJ51vg/R6UHuQtjpC3oqjxuuWzbSnTAcBUnX8zY8qKgADba6l41Kp9c6U8JNW3EF
DdoFmdDZNpH4ZXIzJgLfYqIFMEDZL0LMNYOdu4ii/wykDCjF8z1MI02EMvmQG1tT
EqVmU3gmnPSc7Vv7nCxSPmQ68Y2XnHcwL4E3649i99hAZWiYm5wK7mVJbb4j1GpJ
ZwHjnZC5y7+bgW41oqvbcA==
`protect END_PROTECTED
