`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4FfWeTndByIsIcsJAfx7hWVz0Tm6ECcd2QCfLsUedT3PoL1tZbjBnmrcl3ifhXDo
i2p21I+O4UfNP+nYiN+BVFHm5BE4Nk5cew5o/R8QJ4Wyp9GYTnmOFUNStqd0NP8+
9oDc0Yi47jp6tKhIYwKb9ymzqWQnCuVwo7KigHfOV28vm1JRdpDCDBqybXW4ME/F
JQ0NPdvfjX/6DTEJCPymSXAptTHG1i4gBRlcpEsotCUZ7IHyX5jLW9HbYReC6qKq
6hKFU0LrvpTSAeDOIZrpe6tVHwRFSVE0wi0xsYJeH3EonrW4s4HWSSxaE8DALx6C
C4Qnjhs5W64nFuLltYonyokIXuM8xUEKxKu7hBpHq68b8tGdnLIM9v7iH2CrUINy
46ljH2ZZVNUU26VMciHFHkp6RpvmpmU/YeQgsoCPmJTDP+OYDbRJ24j9PDDu/6a5
O5+/JE8zwbNTAsUYb6LvZJ2RURuUod0EEjMrUr4RMuPpOL6wPE7jSZQB6bATewo4
8XsmPvurowJEikrqil25w38AshkqY9KsXml011X9ZrwkxSDPzSse40ndE0uooo+m
Q3TAb/iZa5bkFm3f83HhoK52zX6RPKgsVufVGLE3CWuIAxsH1dEumtljQmi7ui83
GsZyQ4N039Gxykdc/5ByKGeEy07pmcAU5H5wyWTZO3a/DdRC1k86liMYuZ0y33g8
KfYjoxrX0nuZlxVX2zuw7pi3Xs5jR/xopj9Bb/KiEe8MjsqASfg8zvbAW85D0e/W
YLEBzc4nQiRYsJq550gWdjZgV439k3JZc/tGPPwZhtdUJxpWnRTjAaNDIvvjwUCG
XJZHeOL0s0zQ6JRpdW1SjnE2l9RgYExvV7p2GNiJXvqGlbzPkTcwADZWoSXDtny+
mzP4UzZ7zFxMfZoADvy9/QHkO52cyvAysQN8jSxyJHCN2rIp8bO0Q22W3JgIYNwJ
khydjx+ZzPqNHXamv5yT1xTtn4AlC3MHW2nleEgPc8IHwkvkFYGbfWkgSaJc9mTm
BhVrd69UmBc1i5tn08sHtOszjGYGGQGUUo2gtdpzMwc3O5OL5HEhavUOHxIJuiJB
5720PZoRRBV+Kc8yXE9cvF/jKyJrg+ljhMcwDt3lSecp+qLwdMv25B5MGQ4yPN6O
bYfXWi5h1mmYZUtA6Zb1nhSSWYRjQoQVLzRMPUkCE9n0rR5mDw6hU1rgEYFg8r7G
m6Uh5c9r+nsJqKBAAdMO/VIVff6It2LzEDjXP1IvXlgnVZp4C3kBqLUCD2vGrF9T
7wIQCVEUErZ/bc5MPE7XMktt4AEOLmjH8dzRn5G+YaVm3bqi81WXfbQagx4a/O7e
ObrctzrFO0Ra0Gx1YlP97DfzYtVqKuUVJS/MxYQr+pA988lZbX2eBu1CRwC5P/PR
EcMpkd2qyUQpTyyioezCgfv3ow5wUYA+rR0VsOBr11kkV81XgVVnV48jSxAsY3xp
z6x+rj13kEAM1xwNj4yV5yg/w2hL4qGTbMJmqlxVuCqzhj6LFpNLqTAaN/ofszo/
AXmTi4WE9ZdTMLfvltIQg5/to7v2GNUm9XdfZSHzEdwQoGxcpsRtlcQmJQtrZOAT
NeTfI0i8EsE/d8s3fMMvKnaQrgabqqHhzb+YCsBltg22lBh1GknV1EyoT/XqU6g7
ZfZBjkmxyIe/UnhONY4VfNQrE8nrkyD1MgTifOwz6Icp9ZGFVgUcMMTyLFe6dofg
nijaV1nIZXXXDFS+RI8gVSPAQ8bJX7w9WiZX2rDxVEIINM6D5dyrkSwruuiGeC8w
OTU7ERzNsMrUUDYgSp6eiC8mCVMIeq67lX5jQfyJFWxPqM2ietQ7Ze50PWT17yC9
BYyv1zi0NEl1fnciLhfn7fm90jGcaaZ8LXoTnP/OP/ykIAOKaWuYnB/v2eH9YbX/
eNQsvDi948/1MsIvrq1td0KgVrbOgUiB+fKkxvCDDQP1Ot1A0mbZeIoewLrAiZUt
CEenq0ZklZX5Ntvt3Ury+SxpTCFQGKwisJCV9+m0G2npiIgxdS5DFDqrI+dTVXcx
sZ4GIwhIhcwX8He6dZWTag==
`protect END_PROTECTED
