`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nHiGKfT6DKFBL3suV1oZ2e7lrzfCmT3YwTgTapawrmc05ICyNM0I/r44GIIDT/T4
nNsDIqW5rUwowWYMfxzmLIe1Bcu6XHCjn4Wyb9ztpnZg1HUIq23ZOC3eA0XV9k6r
uoijQV3ESqeVN/9nlGIeVSjAzENi71U3EL8jPeDz4QRowhNrE7EV1+wZkdEP37fV
fpz8uoRClfR40Bd5I+f5yNF3nkg7369Gu/PR5HSKpuoASb5K4Vva+qM/5DMg3rGB
wB8ko5+R8XiXb9scxZwBpBcVSIaLw9756bYiQNUwIDVpfuc4h9a7f6cmwI7Fnn0T
yY8gGPUx24ob0Ysd3b58OAu9CB06Ms2ONojt1nVyTEesbLfjKcKWPwWsIGybYNzA
LChmzoN4ERE7126kIrRzOjIX/gJ0ptAbShzyJOtiEGzI7pdMdhokGvLDTKArGOAC
V7Re3JD5oRCAixaEuQXspyyL0MCMfPWWcQmfkspsNkWGvSnMhUNkzxvPPXbVlkzr
pF2MCK+1OQMHHGDqtJz33rKEX1tovYACzF8+e55ljlkFEsoUrnSgJfJHrV43j951
MPDk+Esh4MYbkIioErd6hmN1We3K7iO4OBgA1/BtFAlPIcRpyUtBei2+jQt6KXBt
3cMRoPyPK5mkvw3l0yMgwGZUixPzHuN7FJRjBBNVKST6OkyJ9Ia3qjaBaekPdGDk
fpj+hTpzcGjQxoXsXlRyDw==
`protect END_PROTECTED
