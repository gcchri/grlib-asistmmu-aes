`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fZvSqLQwW+opjnH4AV9LC5dewV0NPbKC1mAjn6oeEBUxW7GdlGNpWzuMIchM+3t1
U55Vz5htZxdxwEvTQVZ71Yca7p8kLMeMPiB9rHpMk/jbbAsD67My6EsTR7p4c7Du
ssiLodTQfCLX1Atnp61WHbs9y9hLpaU+P/lAHVkk3Se0kLPZK/m02V6cxJXB7q8M
mHmGN69ARLojZKlq9bPWzbpvzT/kWv3SUL7AQhr7apQUlsorBQu5P8Kd2REwErte
i+I49ciIracmDlRiGFiQK6sjFUPXa+Xc+C9pgsS+bj3FBUTPA4dt6x36RDgbELwC
kzg4nhbPkomRLRzEZ0x8VZRiZctJSw14lO9UE9usWgCFIMdgQtMEvztUHB9byC3y
t+KzvGloyWG+Tt0wpDLwbnv7wof5bMLRPFhj5CK1u6tdQsVMhd258Q8Ng9pdFrOF
7/D3fxQjGsZkHhsjkdjOvuIvnUXPFYYIMByziYAwIU4qWNXu506yjPZskxFFWGNX
9PIYqZMbfjvRc18rW+AhFUhyKa/iRUCOqJKMB5rOxNQ=
`protect END_PROTECTED
