`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XSKQSRLNlvFoHOnIYUzev2ojjI4pHo6GzCvUoio+Oi4HvqlTX4gGHAhXGfT81d3p
wjHaZa42sdLTqWM5FpLP8xpxyJXIHH7I5yn5gzJOcmut8qIFlX2io73FdrfB9hfT
8rkFxtEJRLDw91e+E7GF1rneTt67VCOM2Y2lmn53e0fqzFw7pxY3lLHbU1LE+Ruc
KqL3XzfsnuKnGTdnv8LIj02Y+ShKhPXrvgrAGFfhfpO6vHJY0+kUUQjKiK2mxTU9
jDs0gm8kUUS78S7vpEV4sZkkeIRgJRm3AOgAVfwPKWyVxoODbf4gx45oLtcxscpS
FcWuVZkUzbmQRK5/vppLizCieCIo8ZeSizZc5tUHudwUsrlRrUnLlQvn+Y0aqjO1
J6ATDnA/v2knFJ184Uw/favKCo0/rhK1cmjLOdB9x/k4TwS6/9gUcZEo1KzQq/AH
hn2u+fQUQitJ4P7z2Z3R7MM73cxgM8J4pi5LcIR1hKl9C3K8Y9+Hk3cNL9T6LcNg
RU914TD/c7JO+tck/un/tmC2r4pDt7a8Na4tNAULvgRXSK67aZuD1bNrUDnT2hoX
ihoNkRMOEt7Bwko4yZyG5lTKKkU5/rSpxR2YYXb45MzZ+RDRrEDMvzDbbPb+SLJE
Bz4PvrtcJXXRgxdBn6jTvYewAs06atomU9YUvW2xZQHtv++1ccMLuWhxVGIEGMqY
MNAcA6fTbFZ33g7umGfB044/lejrPP0COXmxNmWuGoZiCoeOsh0U4+s6jFYTSFgR
nEdqDxkb7MhVgwQzluA6UqoAY9d0riOE2d6kZKina/oM3ne9zMBTHapuuGxFaYLV
+BkF5RC7RT9nbwXF9a3iJmPcuMAakNaRHQ+mXLew2L3M7axAL35759/tYvzsrWK1
uNQVWYnjnRlihWhuvOvpGAD9xkL5kwlC/u81g3GEJ9+NB1nO8qlGsNLsepJb9brv
sC4C+LPxRHpz1OBZdrfo4BIzwL5bjrBHLvNMnsoImCDO7pFYcMFd8B36hxkm6Tv1
iuxYxjcZW8UJPZQab5uTNQ6/xtm/ADM9jUYdl7Ch0DyZ+i1ja0zc5pnLQyp5niMi
YibjoWARXN7YzGZZop/iBzx50EwgWzMd8YAlaxYm3TyCF+xACLLyhgjb+ywwpxcf
Rm/sQr/uLsa/VGepmIgoRmjtE5RQIUpvooeF2t49r2jnoomajJEAqwfKvX1b7z0a
pjiuXA1OU4wuoKBqp/IwKYaiUSZETxj54aBQHCAU2sh852uxYFPA7Djl5VAPl8Jj
d7bgrZt7MqMXSbQImE+6/MomBiTnEcFImmwMi5fQQSrEQSWlF9YKatwos9DKr2RX
OPG1YH/DSXAatmCQ+Cg7od5Qyoq5sP32+ViPUjmFoTgFCTwLX6u+Y0Jd4S+rUWqz
Fzawq5hfHVAFCE9RhLtLQWclDu7yF3TL4v0lcppB6004Qom8a8zA5gAYgxwAv490
o4gBcR8fcOHqoa9XR7QOxQ7+emaL9icXWch/q4i3ZvcKbVv3hFZ6tMcUKMgtEVYY
KUXlyXYuIs2RjWfUncg3/yK+uiIhK4fHPp1DwI01PUlrRFpjWQR1VvZ2JidEGVvu
D05bg9y/hrQ6KDJ1M3TNAjpXAcmTPveU/xAuw9L9MDdGH+EOVVQUXjwpfsgER5Yc
+e3/81HQ48TC5j5StpAyXRwA6e8DsngtuHNQEHutZuRE9qbe/8eiHE2VDlqomumU
AEl6e+WxhNxCUHAi+MBF1Tl+kX0/KM+OJGNfO+p4vYNvnIYTqhVS2qwSaBjvUVkH
6vJCUOUGsbhOYRUbdiKqfIeIjzfbZtbV36qtXCunKQN/dPWsZb+aewf4LxpDp3tS
372NMyvykZEgMH7GJUn8+Uww/xouaA8sYkrFVXKngET4Z9JUwmIuBfORpPpVymG3
R1mRTy5LtU2pzudXiJeiNB5AnjXMMOml1PqhkIqlORgw97K0VdZgG7Bw2nYDSzkQ
8uQ3WjexHa5nvT25G7ziD6+kzOkG8e0xRgoa6ciYg1UUTNOAd2UPvuTUeVvUnyF2
0s1zSbvO/KvUS9l9lSUK6VZGBYodFk8DYVzX8tqo5H4S1lH9mePUHCJ4F497dJvd
DUqfi3U0fFJBD65BOoEp5NYuaGyM867ZYEGE7W2bRn5qnHyv3pxd2cmVa2/xT8g2
h7IRKy8jcAkpUoV8D/VLMCHiymFXk+Wqv7PBkh56MuSmHEix5Hv8s1dO3oIScLcf
Iuq3OplBCdsfysVD2rAAkRtDQ7ry7YPnM80dX/wWIVKDFcSm/eHd3aB2ZOxM2uO9
ACe2MNxAV2pHXHp6EKRCqhshVwQ8RQOdDYew4XQW5DwSCVbvPRENwAKLNTaBqgaa
W1/gqadXyKzBrHJx8rq8ihdfjdD28ElMv1RPioFPUfNj2CF5CEFGAB/Nfz/4lcck
+WeQj9MY35CvKg3nhSlnqw37G2IQS5AzswAwOS+QY2j/cOm3A3G0YpCEZrL5WHNe
wsQffIcW49HLwBQUwAcH4XXJKa9bpEabeDxXX1N7P5sXqSB70y/byyOwd966SK6q
BEzd4sePATqLRQsZawuGvKIgpx4qgJq+GHfJyUdd64Pb5fuy4X76XoAivKhJC4fj
P3vll607hO5QQ30M8KL9G/deWBRlpudbIMreVPHitGLCiAk/nfa8pquOOTqoHsvv
nyIwiebpip6pkV8bflYHx0AlGRgdKE5nTlpO7XEDS6R8Lq7nSK1eol3fIbA+SDoS
Oy2NiU0HQygNOtbL3qYPx1SjpBxGTmj4kYj6yTtk85mXOGNMMB5povbKby/krvut
D+y1j6YzSJApYa1K8RN9VTblSx+sLyuAKHxshpONh4d4n5zFt5fxyjw4lRJGTZAJ
JFz7KOiJqjjFYc/P5fH/Pdn7nEoOB+YobuuvvNofSrp+/pprlErpCW1PNX1hZpo3
ln98XNcHU8/NDZAbY01WeBWsccmYH+5daY5njg3Lo5SPtm/aHdiUoOpyU9Cm/Ekr
/9q29bsmymCgLVPWtngu1K2rZ1uqX4OnWG/JNaSypg5+Nr/utkzWlAFVsN07JGMb
rwCr8OI7Z3RLJoYVs7tg8NiXq1+p5j2Ph9hiIyss+GgErNEd3gAu1+Z5m/Z6SHPN
5AwDO/GnD6JThgbuiUidOsQ4nX8EQ9zCqInjgx4LyzDWGKDfAp6eeeHBGXiLCuPC
l56nfJgfULtF3dDWDrqdJeLctqC6Vs0ds5M9IkQyj9ZAhOFaACXfF3frIh/kpRs/
M01GjbBcnFT0CAUZ3yKjzIKjNKor4LdUYWwXWfDfLx9VUlspwtTY2FJ9u40s6P2W
+eSs3ORBfKCj6OkqnrKCRD6sK9TCbT0kittBIhDuktFkYwtoZ37S+tInt0veuwUV
XtyeUOmeJNOYfy9emmUDQ6nzbJFcS2pwGS46EuIMb6Hv+jhF7+RaSAJt0ela6zCV
QDcPBCVtwwtjFQfGrReddFu52tDmPQH7aJhb+ApWYxIdddIWUbH3BJYZpwSfeID5
O/NL8coNP3kzawDCBuhkD/FrMfL1ppGqe0YnzceJvz8Yl+nnkHZHczZUIyZ3jaBa
C4FMTEIFPJfM7cvRynDRM8i+N6bE9Ge/u0QhAPxXJuMSvs3TNgim5lZlaP45Tt9c
UG+SiVpF+/3dc165T7jK5opQwBDvM81lG2gOla9BsLxCZYKKUo/ypS47W6nCn86I
A02OVRt0oEuu3JMU/vAkQKPz1WEKEEzsNPndrDi3X1rqPBxibodi/T9XF8tPjirV
mxB2RgILi/3qQpIQob83dtftewirJIs/3pCK7hCd+jscesYleuHHTWZH+1wjTTuw
c+/UP92E3OrnHi+42qZav3OZUzD6Fy0VFosiQuS7U+eUXuhCOSBmIE41kGxqO2JA
SSP51rp2mW9/dFlH0WIiqa0Ya3RfLQRrMPaDwfivHVw57nf/dzcw6YrY3QLkQXua
Wo2LdQA2rtgHFU0tvgvGAsjoJ9BW9LhhTwvdeT3CZvw7bPpOjz62d/s2KOQet35x
Hn5xBrzw07eb7dNfi/YnyKW5BzGoUhUkJEQvMmJWfsxH9ymUNR4JAS1U5B9M70Uu
YEtM1OZOW6zRbBUCIHp8RNboSJnjRM/5Xe301vrl9xlP8r+b39GeeYvbxDMN7ab+
1d9ZuZ1L7Tj8djol3N6U4FtZ3f/5HB3T6vKSu8vARJpWiyxCQyeLvG+UiB4oaT3h
iN/JQMUyGw9ZguUroFCtn7faM3m8XPPoSVA2SyIXCUFS8j4K0yhMQMWzTLixf6eK
ZWV2Rx4lKugviyjB4TZkHj9FOKhcUlV8n3AouWpqSweyaZs94M0jYJCvb8Vl9Cm2
xmJTVeURETR9g5JVrHzA6zSTp5dpabp4ImNhpm2Ck4V7j6krCmrPNkwY6kcb3ADQ
Q6/Up3LhGKESgcqqJ20XQgXrziRLMM7sSdR9Nh8mWQ+ydrjDgChupFIHy7z3nKDO
663Va6G9SiVtwmxBfFniQ6pQ3LhYjgDKGmYnZol6s6RL89g6TlJIlrRnlDItMWIV
NdEjv+z5bZIFwPwnsbMxEDMb7iI4/8MR4lTBumSat4wr4AwNCtl62YvOUchC8fqZ
KGTefoWbsBYIhuYthVJNaXnmTIIeqsB5hzOr+kMNxpTn1K7YZptD2BduxKXRexU9
UaR2YgqNPVvYAfiH7ogy+lrDAHHIA6lBM9vb/avawsvYNC4vZk85HSfzGJdDaWRb
OoasZw4LD1uDu6pkYnCt56/t/x6z9GFwyAbMXoYhjB3ZIM+nQ6pBvzRUBX8pawhe
aA5alMOIe0jJzGPJTXoadCeILklTesZrXM1jBsFJh12vZr1PF71kqdQqMkqzeLfp
OrHTYFnvBdJfOio6trI6J9Bsmc7eUB2KtPIpyzHmin+A2lZ9mOHwMSo2TUefKSs4
Eqvox00BKEjcLhs+pqbJx6WBxAlHlSVxRqUGBE6ncR6+gL+be2aW4YSmlMcqQU8V
tVyOD8oQjyfZlkdO2A6Xrb1Jow6rsW9vnXSrLiuvUzmUvNNOAqrziXB+96Ys38vz
4w0IzJbJA08bDZMKcHdgAZfeyRA74fVuB1ZIPBRue9PtcuNFYrEAytjAzeSYyYaZ
tlfHQSNNuEc2xDyqMnSbDmZc9z0FrqG9IxWv/oM5Fz+ONGnzv4yJELLKx9cnq9yo
b7JnPvLPO9r5xxHES5n8UT38kq05RlpFTw1SXuTzWFeOynfHD3QbcAQAWkp0SQKn
zLrH3L1eXsJDEEsDAlgH03RMMOa7VbCsM42PDXbtkY7C0wEwHi4QkFlt2CykDryE
kYMRYdMJW0GvFWmY9/76mwmFaHXzM5heFAqFPsePxu/ESUFYc1cpYC+6K4SOJpBG
3NxKtRoC/Q36EnIQGW6zA8kzzRJuYqyTsJeC2r68XGXlxe+NrER6pbACZKIu7ylL
6OLgv2PFuRtWtjRDaxFOQZqCDs8EZeTjVll6ZS69TZoP/D2X2faKSsenQmkonG5X
LXvE28x1DnhrCrZ83e921XgpVmB1VpR0KzMRjK6gvjWpoW7x8PMBkadV0aon5ldG
y9245zx5UsWgBZugUG9ljMIWDQTPOR/zngbABO00M6wByzUVhpMk2rC47PyOItgV
UDHyQY1zK2b/ZCC0XLrTQJTzfkqgsAjxnQSJwFBAj1ov+r6P1N4mU/uDjU+lIscF
LerhndvjIOAWNphphQ1D695fG5txMFKuSRvdQ2Ciq0ZAyQS8xnNneOO4Fo5D35+y
mUGC0nb4xaJgTttXOzGfPl5RV5dUnBmuo5nXfSxvVxLtvyxz6xXPEPouaHH+2O76
rN7b2dRzmaV0HpBDOXFvLwCoyVO7gHc+87KKdNZs10666mgDZIPi+kU9AxQaaYnp
c7ovGj6IpU2dYFcBRoJdHB6TChHtZaXdT/YEHfUjk23qNc1NLnFB51/wxsSL2U76
yTFpqfOo8+7DUZf8X7FUAjux0YvmIB49QgeFpg0Z60p9aPm5ljio3e/SHVPpvkcz
Lj8sZipkzyOlqggnyjChAkrL9KRT+K+sP7V/DAVqSxQInwCYX/iacet17vIRPOES
C2qaYw6PQZISazTZ4li65tFKB8eAfxyC8cATLYq1UAR/u8kM22FRHaE6PudqQAkP
N6LaFL9owvZ2sV0arCVSyGybhe+CyEQ+9oYbBQHQs7+esFkyiJRspLU86jDoxhvd
tCokrayhXwOgCXl33mbBS+Hdl6mehaPKI5uR2BB/Ell/B7C5flSJc4KRe82Dtwtu
RjcNrV5pIYsLbZCoCsYTmkPptsaqnVUKvYpjgvTlpfbh2QF1AV/IQuBSSowN39wZ
12C6fCAtjLbX0j8tPa9IsSRuoheVY7hk6TKxeoQW3A836kEof6RNEt4HwaP1qzo3
HfXL0oVDthgo/ID8eYIkGGMa3r6xHKaBteW4Auunu3SEvsbnMnOlBybulfAtr76H
qbF7mcCBELMNSjgrsNwvQgqQksFEHMi++RtuM2SOVVNq7Xnf2bDNovp5LrsIi1QF
kbUsplgwGeQDc9wGk0DmKTvc1/fX0h5oNhCZbwJLv+iQgzenm8FYdtUFdaKg3MQz
CrVSQJ7xqeuUmCcI/DFivFF8qvo6FQFlpFw26cK+r4mOnUjFaYBYeV6looa2H9b1
ktIPbycYRh0X6CERm2Gnkf//x5iIu7lNsaP9tb78csmZVI98fid1y7LOdERp67al
IKGRFt4a7skWBmH5Vn6FUEj54ubRijgkVDhfZYuqquTcrjpQ2nTI4Zv2QA/ub07y
ho+QYPXnVC9G8rN92hOqIogcRlW1Z4CNSlJabM7Id67hA7WQ73J67DO1PBKEQgKL
gS5s3YcQ3v8TMjNv5wp5h52od4TRGrkWz9ELBknyI7aH0LBCZroVuSd0t1UsFpIz
fbaWfO+hioqXuTDWxLiJb4F5ZSr8WSvefJ44qQRsqlo1wFOjcdKh+taHclK8lkJG
oEEvhzgvJecNjianVyXpLgCGHYR8PqdNayTcpAbKdL9ZtLggGtEas8WnfguKF0Ur
zSaRv1ArgXpFH3UOWUVUtB4Fw3Uf358V0Kn/2IrRdHkzpfwFQHlYXEKuzlgCeELk
zk9xFV9Z2LpELMuNvjbC6cLb0xDIXAyDA3jgcFQDUkrF/sXMclPXF/KXa3jWk5TV
R1CglhPBHAZn3e7DrRyZFIjl7363uPJlYCjaPPPTSHa0oC0iC86OLjbDkFVyCMpV
qDN7600BhFJlBE/30g7FK4qquh6aETDLGYp9LUejMlm2VGf7Ccr4u3VnEIotK7Pn
jexmnS1tXQoxi6+6BcYcxr2zQcb86e/28IK9FJDIDfq7ZAw3O63flzc6FgO2FPcq
eev0JA2t/fGytEOB0EzKdWf/qzuFn1c5500nOzbxG/ByVqsFkpWogQ6WZk3PoJ3j
Z/Bzf6yxeu+OLtK4qvOqnqF2qiHRUh5fYjB8b/uF90oFF1pbw2KF89MV/IZYY7FU
ei/H+07UmuKPHu8JkFfZ/cnQFBUWEk6O6tCa0gM74ozMVSJrd+Yv8pbuBVAlpRPZ
dt8oNbBlbs+8rkZ6wXY8RhBPNiqB2sw6B8YtNBzIglyr7LUuof4ct5YRXsov906q
Co21DMjSKUc956GFUrXqBU+kqZVOJu8ALc478h2CBmxL6Bojl9cN/uOOzTuAtSu7
jSmanVQ/t8dkKaqmj0YcqgLujUeK9rnQxg6a3AfOZSxV3VGjFF04Ig2/YJHzxRsC
qkU/g12u4FKz09B+3K3kgUkuCYduU+d6eyEBQLQLgFOogMgOrMDLPD7fXa+aj8PN
YIw1kwMDnKRFIpxTXK8CetSSFWjRo1E+rgsJ0oY3rHtDUfu7k0bizcmzuHRMedsP
k38X5JFHRXcWBfBNKogUvuTzMBVV2D5XPtKvTjwQCg8xHaqCZ+ToDbbOQBZ0emQa
Z7L0e9dLOoRi+5OD4agsaDcbBh79FKCXnvp7Hurr9fiVLPy1b26qfByxdSDnHfc3
iMbYG6tbdtUtAOlkqjp82FLMVwu4KQ7tvVarKgVUWTX+rt4yqygqwyJOvsSRYXmQ
B6fgRBlvr4lUzZ8Lpy0B0a27vjRhV3zX9RKs+aPxJfY=
`protect END_PROTECTED
