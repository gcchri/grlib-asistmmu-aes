`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l+4kiG8kx/rUZkOmVM4sJ8SJwq1o+frjKfvxL77b9NVlQKBC6JUxtJYTR11TlVPu
X3k0NmCE3JzWIRpxvj1KxuEtEjXdH2TP2+WKx28GJTa/WPNRTK80VaLbAz/wPCvo
6nnwzIWaQiF77+1zzN52jXo0URB6Py7FhIEM/9peJhZTB+0Javmb+mQYwDJJ25KG
AMkgchmGrXv3PIOcLy4OJvqLl4eDY2oG5ippB5smL+NVNxEwn2auHTN1memWSaEI
bfMPtzByodzG0y9Acm65ziR5IdfB1bTYhKrM7FSUK/vmny2E/WSE/NJ8SaVu3Iq6
JjnqTPl4tnLj/6ilhbnyNrEhvNoMiT7Gqs3NRk0rEmcymu0M0PSOziXICsOYEEm8
34iwGq5hm1LqyBqWoKA36sVoZt0IQ/BPiuK5w0Fuvn93Qi2ANxan7hHUYHT0Mm7e
5dyAWi4aAJrC1sF2MlsrkbNjEMTrkAf4/3UcKhJy8ixAFc0/X9vOEkfE/GC88nno
oQ12ff3kxQGAD4gike/NXSdawuEUVwgk9pougntCo6LCs93NqAQiBLs3rozcQx0g
zLG6hhcTq8zjZLAMwIqXTPU2IlJ7TXNxBXV28Y00MI5Pk6zU6+6+kkYkR8HOHHv5
p82JdEdmEsWTkJRQUNi+M1vn2ayM2/jFnl24WKHr8tjLm6HHQnzKp6VV6eZDdVHG
ZMkyzij33GlZ77/0Ii9ddVVzYffrAYEcEFJV9zi8uW/TZFaoeNFPwrPT6o1XLecf
1/GRxCdIuAl17tH4offorUBVVBmlIR1Gwsdod4OFP1u7M2/XJnZvOqNdSgybgsdy
IavWgRKgPrCmD4UVuVewooeMWdG/OkDWkTsh62QELH21sL/qyfvcP4vlGJot/F44
Q5h2P1Yvf2wXP98jIQjhDdGGjSnEQIYz0XR6QeYwN4yDmJzZnaCgkayOhIhvp9rE
DeM1eU+I97cbOyDrykCKuw/wJTTzljl+WdXQ+sKGOWhN/IgH+2pkzI9F8U4HsifU
aQILbQ2YrCggtVW3HQ6wTu7aKQFYHp/U8kHduQ9RCeXXJ0VMRKwFCGMVJqqF5mvx
W56hse3QPvM2NwkcZ4pDwjMg7CGsXaiKX8ZozEoRe51Iad/k/CbBDDpIxAZmzSF/
H4CZaFcbSndDkl2JQDUMhDNMh/tB+zJMr28tfDt5enMigR93uqLfMsMAE/hPJcpn
iQnu05ytIi92MmqTDhpWWNzi3dESCw0hX9QuTzg+U/5DD85jRqWlEWvpYFvyUdRI
GUw3hLdPi5HQRfdTDqT4aKC5gmBaePtjiWiujCSPa183D4x2u81Ym6BHwyBnxvbo
xNDlG+G1bGeLApjBr93KDtFhSkDxumBDkU77uybKEbO7HezNm/tHypthAIS18ojq
CsFoalYiJEZeg/PZK4Fb6mv0ultypkWGndDesneEV1+DhTVQw6AvnDFf9W8ok1da
Ztw53kkwYBcAc5bXXqlRDQ==
`protect END_PROTECTED
