`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QqiAqW2hFr9WjkVA7yQuI7WrZsKWprFYT8KBeA5yThHKtkkMk3yoofz3H2ecztKc
JRSewhNEx98Wr1oeuw8iIEXWsBqW9ZZWEDWp/Jlv1YuvK/LfqB1O0L0XffG+pRtg
j5ltzvB0yUWr2u5hrD6pLfYKP0M8yMbAvEdCWukjnMrGREKEP1/2RLM+ZYaIKz0+
wSrMPxurX1XOKgcmdHIigzsulurA2AXwwKekXlkSE/FUJQIqYYQ6rd0MmpdV8eWV
D3kVbY7K52ClqnCR/tGyHvJRn+Gsc00TPmM0/4dwp67mznBgBczJweOkVoEM9mAq
mD/SIFPZGwV9Y+yZ1jWwAj8RwuCGMuJ9W/485dyr4M6bcUMUgErwznbhSPbzsL/x
PPkxzCm5eIB5kc1RsOUCzvpnFYqdmfNPGr6j3QEhY1M=
`protect END_PROTECTED
