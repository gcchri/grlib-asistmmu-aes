`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3m1wIgTkAAWDD65DaRLb5W5LnMkHPfvB4Dwyos/aBzYEyZzdyuljvaYAKsHh+paH
SpxawheP69AWrW2LsgXU9+VaHsnXkvivIrBAGj66ZMYqZCKZvK4ew6JTY4ekk1f8
aezQlYEr8LlPCVKhB2gz5bi80dRPUgmbDoENGSxgtUA4r7uiRWqBydlhn2DNY4d2
8UQ99G49rVfs2HVod4VDNLvwuUg7Ybnq9WnnLx2/vieLpELCw+TyrUFZsBbKaxLD
ParFYJ4KwNW5F4yz2HLXol8zhDHAheHBZlximwWS5I6TINaNvPX1hfm9X14qXmc7
fg9ESbH6t34Bwemonjw7X+9LhnZgc8xnh7BmHRRdxIsY/5ytTvWG4NhYXbIWoFeA
xf/5MlFsCGd9xwQ9S6kTNERh8EWRZQDnyqsAsqnoJ0/LvOqzNROhhnS2OGxuIYBK
/Yt4aTLYh9Kpo5GZzWqZ4EJx8igV3zj2m6MPAkefI38=
`protect END_PROTECTED
