`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UBoWpvQQ//Bf1hBbtb74+rRLR04PWf8SFhsztY4ZXADD/pya1PJ4oxbW9ZltP961
QPeDyXeLUQkYJ3FEYd8XlS+AXI/IRC6BQlQGThi7FCRMfYosum6XmwWhVgqI5PZ0
jNBUp8B20SrUe4Pe09dZ5cyclXteJ7L4YZJCJLtAqtvbyl0302r5UmO3cocn7sHR
ropH6Piz4ortyHYHzA8zBpCCMYEqaxD3U6Ol2ebT28mIOH+VEtcn6tPK5IyY9xM7
T6e+/NRL0BfxUBVJoubAEMt0vakqfvrz+el93kBSMeH/bnYMrWHEkcOWJ9vXSkZH
OR2GXERzwSADL2aMxNguJV9sFDWSsmMnDjmgUmAA9LyHc4pvEM4yEX9vLfmZMJFh
VKFqCfq+gdqcsO/8dVqkug==
`protect END_PROTECTED
