`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SnZdMHE2P/TEoeajffvtpzjOnPHXssSkq8t0uUzFCK06uQ983QRfcyOE+q8oSvrE
rP5mhBbcUboeEtr7sRt5P0Bl/DdFLCzA3t3rRFL3PuOXSYYgaD0bzO3RqxMZEDN2
GpXsekGQUtPROTaAA2+HjSnhYDoVAqCpo6bOcm46PXmwuH5tpM1txTWIZOvuxFNv
17tjef3KhqkagG5abpI0UECgaUFRKg9h4iDdF7FVZm1QG/A3aTXT68/LQYIS7kG9
UVxOkM3h8Fk4uUVAE4Yb2Q==
`protect END_PROTECTED
