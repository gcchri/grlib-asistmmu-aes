`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C6a5DbZMekft8yySkjTGVVaoW09ide8AxL+oPjDAInjOYniFFS9J5XMr5O5L+aEX
iZvObCggV/qXHdsDGFoYipgz9Zetm2bp/uBQjBqQou0p2i2chuV+BxO53c4I8gaU
FyVhQW315P28kXdh77x0gE/raVI1nKmtIuzkpQ1e0WP4Qljg06pi8WAt3J/dhYqk
VpMuIWeTqlxaYsyNELMwkbBMlfP7PyWLMDFNRbEer0NyoN/49WDzuKxue/t0ldxz
7mbbm9LL8oWk47LvVXvE09JZdTUfXHM3h/L33OxYXLrgGrYxBm3f10ZqOHLYwCJ3
udspO0YZOSu1bjunFdeyBG+SGCjHj0T1zMv2PjwVdU7P2tRSLC4HuelGo0GmUCyT
H4SFc01xGgTdLTvKkxQz6ReNfJFOxdaLS62qGWEI+v//0s5d2IjV09WA4HMOTHkY
IRyrNjsQh61j/G4AHnyLScKMmMYsF+MZI3q+oDUHAA0DePNmbvWVX87Iu/xhokwD
esn8oRiZ/RCSX8wcTvubL4mbkjX4J1XsR97eSAO64/GXiZ0SWvUtQei8UJH01J4V
pQCjFh7jKUPAj9oW/bhX63Un5myMIfHcvMaC1XjSxy9mlIE/v85r2M5+xwSeOVX4
7V0otYobdYZOHhzX2QdBmpuMLPId1crmn8vDZtkw+XU=
`protect END_PROTECTED
