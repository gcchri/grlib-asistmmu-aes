`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UmHP8eeTHJwT2VK0c984QY3wL/Ere9zrIB9s9LdoL4C2vuw+dF+J4mYpeN69A+tf
C4AyEdC27RlEjYnKSG692+wDRC2iMXWmqhdxChpvhxLgYaA+Rj+3iWamHB6cH9xy
OvgMXPUqmedYwtprq9lyzpEG6pZsMsyiUQxvf7JCIfhHESY6I/jKlmPnr5jumUs/
ZjSzhKedoCm71iWx7gMn2OYTGMzSVCexJ21ifaQa42zk/YMOfTx+v1adgHInvUWh
4uC+H95U+R5I0J2tRKGKOfBUcXERjpvabRp7WSq+CnQHvAQm3C1Qj6eq6uQWP+tO
zVhtLGpDMEZCuHSZ71Ck/51d1fG3jCIFTAwzp+WJf9fSZW8MT8V3FT24s4ACKMOb
aUa3zk/lnwFzTq0VGd+qXMLd9LEnVGNj+nz9AFxV92lqQdDut0+cdx1F1gkPPYx5
kzTquu9nma7Oj9WOLXyLy77v8iSYsFi3oNLDcMIz+p55mdb+39vvfjpVO6E3Mb+m
pWHgjzgtEXqF+5cbo11lZBU3Qz2+QQyxCER6Zr3c2IBBWPKz0TplJFZvXXDtN07X
4VX243CaBzZgf+yQnLSJwmnd5vCT7fS2mJh15ZiCWAAhyG9tcKzviXTyng3IVd0u
cD/77aQgnYdGx2tP0yPR4HOs62rgFCa4VFe3SkWidc5jw2zawwvNZwS3IjUu59RA
epI+VAbQVqLFnvKeOTSnjY4pt0Ul5Xy5AdGvxDeatO2JtH9bQhmfZDD4l0ekN1LS
nAWs2jLB/chfIVEujaDGKvC0LElZx93umuTuIeM+nStczKUWL4PRpFghq+o43MX4
g5mToVa33Dkzgst1G0LucgEOYvRHBYjqM+CBtoYp3W8=
`protect END_PROTECTED
