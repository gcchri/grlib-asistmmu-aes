`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IMf57WfdReX0l70KfqBhjartG5oHG7l8RfXQk50tpiBgK/5puPyAYB68V4nG0/bd
LIueGO2qzFQLhKrwOzdWlLo5kHr2YpunVYclefZiBTUnMYmPWu3MFo+fU5/IQvZn
/CVhZoczRXMDfuTwuV5eFj9phuKRYGiXArvWLrhWdtIzrlbB/5HxsIyUyDWSDr7W
f6gvY0dVs1x9Ki6yDDqVuRoJZbhKWrjHPbtEeonTslvLo28OggmsRWQcEc/y0M8L
GQNfS4eWJnVMcPPFpoSdSoR9maQil3HslZuKuTjjdYfBHG5PTdwwRouKGnGqbgh7
RZRT6s3iqhvObTqvZzix/k7bCPYG5FAhEaFILvzHpih24i72zrFYNY0cBWrHITHx
nlcvp3GykNU0aCpY3SFX2GnHtDv9o68FLIgD5agh/sRSmk2hjY3VLbZCMMgcriRU
W/02lx+Uqbks81n26DeFZWM1HvsFJMYtv+6Xebq16BVSvac4+aNFlC7lpc/aTzbK
`protect END_PROTECTED
