`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2UfmXhnvOIiruv78WdUacucPe453/Cl9ghjEcLdFETEtPnuS15bl2HGSDJdT7SAo
5hmyrzSE+5TAxAOKTP1+vc4d07bFldLlk3UY7n829Klawo2G+OmWe7hTvb2r9gLb
AZRngq1eeIYw5miAgoXJ5znt56JoDL6H0ZwWMykdNDIUYyeU5+kZ5jz+ZxefMYOO
pzbe8J1D/j6IcIiMFVRoNGmojnGQKj+z72JsWA13QlVVgwiLsoFuStcIA3FX1HY3
CBT2+6YPlKEZZjLtocGm5Jap9Q8780NrWqb5qX/1WrgwFo9Xkj9dCzQZ1zBMSqBF
84rpSWP1/XpwxDZr2xkS5T8JvsjWUPv8jHYrdsi6LZUAnNRoGjhPThqvdiaRv/OI
`protect END_PROTECTED
