`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2FuHFtrRKyUnxcKrlTCTl2ZeUnaWTcDWjiRzqBZzVcxUMeyTuxkMjnzhmdgtj62m
RJnlIZ6VD8S+kOXtmJIyxRQCbppjz/E6O47fowTIVEfrwrZ0Hg0AWvDL/UF7ZAbB
jc2X4qA9ww5brhIspnY7cOAlF37h26yAf/stx2HZ4WMIqr4jtthg16AtKIxZ6oCe
KPv6SKgbyeJii0KEuiWI5EBCcd+sQcbiAfUC9PmvhX8gMuf/X5sFwsuOwuTTdw+r
UUeye+C4QDWXhVyyIZA4M4NR9+Z+L0b3shqMKbEdEo0=
`protect END_PROTECTED
