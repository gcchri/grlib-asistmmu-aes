`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vB47RepMJJtO2DcEmgIV2R3YfYbHliEeK24ZvwYBGxsbbrXSqXa/hare858yiZCI
971Cce7zl8GrBBJWLVRt6t82Oe8QzNeFHRlNw/RKUnzJSGwau7HWowxTusx0Gk+Y
7c0KSHUJWvBUHNbYp5LdGf5+d2cJ1GHlLzoUGmfwo7tRx4C5hYJp12WwaJSD7oSU
8WHXpDU2skTRQ53kahpoAtjYNomx5gyrNGzdY1vtCdC2MXqce/hAy5NiyeCZAzZq
DhkkpAphh/0sogYnsUw7MllS+NZqQ2mgBlLgrZ8GAIt4ONP9qxUjLD6+nvBTOkfN
MPt92z0PYEirOCJBygGqLeOg8R4FZDphzaGpPclTEji0VRFVk3rW1gXQObBwp4na
d/oF5pCCIHOrb2cNknSNmHD1bMpBNhP2o1Efy2mwOV0tZ+wb3jdLW/CexmvXdZzg
aKhD+S8dp6JhcjhWw9nykJtaW3D253RNwFVXetFk0SauYPmUt9iB/bR6WfTx/jfn
YbTnUHDPXblBIasjX103dEWn5SVIIEMHOkDimyFvJNuxbYR/UGpKwqI65ERftdpk
uB1kfJjhxOFB3Mpfv6ObMBIJiyYWPpJB6HdsWySiNoUx+DFuF9Jb12qEoFSKg05g
v6PY6YR9hQm+rcGvRWU9BQJ5cYKQ27tdygQ0mSjkHhUVPB/mCDvn447H0OwTksHx
S3ABeODoKNjvAxE15TrTIjEB/ckmDutoQkml1zKkaARA1WbS6qRS5CZwUlW0/EpS
djKJb1lkKxRdDCxKmVYuPdkJIrfWhBK1JQNS0zAlXMshQF46Fq7kzANU5fhzKQcB
nZ4ocX2QbsshgK5+IIlk+MDUXh4qovVKLOYB4v1m2tM=
`protect END_PROTECTED
