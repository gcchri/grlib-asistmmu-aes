`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hJ4JGP9gDIqlNhrivXLNDDIvs9zH/OvXJrLnswKYqTuzKa3p9IUsnrVU0zUMaf4P
Q16yfiuGfziXSHBO1Dk/cP+eigE7DQPEJ79rRdi3ktyI48TedZpqhXF3CqR/3vPE
itE5uwJFa9LLvFFnRCsUbFcsfECOuoMsofHwAC4oi/qMCgqJUulg5mjVom38dP/F
NFPs+V+4wY9jFJWdZOhreesFG7G1SmNt2ZTe0M2K/YfTYGDgEMxiLtwaIKalh9FS
WeemJuQOvIBV2cY/JRP07VmnBUbjoHCINDrdKK7WCnmwKNtEV+kabu4wyqyeSFO+
28rfUHMeywNFsfb/FmvVix3yBmdNTnd0zj+qpyTLbj11ra+koQ5XkSkx2XCIJ+wg
0SScbQGlcfoiQwrioVYxzBc1lR9WTwn4pVcMJIZAyRznb1deh8ggXHhnAdwARfEq
o/M1uz9+UM5DSZVlc/GeGRp0fl9k3hPIwbWRZBERtnfosGFvrk8i78Tn+fhJaIOJ
9byBrj1bIOwU40RRlsAjfiBW7rsENur3OFzmH9r/N61lf10RwuDWLcAL9Iu8MjcJ
Rx+xUaWyFSgJiWq6EtJbEj84ckX0staqGidj7tXJyAVoktBsqo6q/zvQjo1KrF9p
FXv+bwNrS8yINprrvVDyJw8ZoLvs079rNbdViH7PrG8=
`protect END_PROTECTED
