`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
32MfMhradyKgcfF+jT/y0v0hZEwJ6c1r95w9iUEJCqfxcXiSLiIpAhE5qsO6XgLh
ZWvKUEs4Hdf5XbN9ZIgLWcAxWMzC+lyeasFt0mRVd/tdZPEbBPYWLNibmfT4b0q+
mVrQOVuk5Sem0dk3rk4AFpK1qaovWlrw2mdQBaDhzOCOzacGlfvzFNRnbZwCynyb
PQXPHWdnXI41ZAlhtp14OLBLQtSrwUDuviuk2oS7B9uHArvAz9PoIOedk+3aJ21Y
Tr3MQjpgtVJTapN/UK7oX0hjW3HDGfgDu4xNot7wrevNRhD6bZtI4gzRLBIraVxb
jV8n3O4kHHpRnaNoTQNDbMbC2GfIEbxiPTnxVYHDprIiTy1XbgZ/W1QzLQvJPTxH
iHBE4UnwsWIL+xd0cD85NEIbXKuKlyGVAXXvM7kWrWvQ2QSgAXvB7rX8N1juhzdm
x31a2kgF0s1ZMSFuEvPtFga9jy13pH3imTLcNbLkx9A=
`protect END_PROTECTED
