`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5bKZY2aDfFpoepevH1OjagB8/BVJ/DDkS2eQF0mvWJ1PlQ7DGSEqR4PTjd1wSUfC
ZqR6vLt1yEwtOd3l6/AVfKg401z1bwkvJ8QrEqwljNU+i/oa9eiLuHYLSbKdcGkk
xWP2lvUievY2h/+c7kg7kZcgu1GDTjrkfnlUBBw8N4uCZ6xW8jJnVjvKUq1a4/gP
3mxt20DXPLp72LYNvzC8N7Ega+w8E6+rVHNUGxpZOQwoAWnN9m0z2kj6/9AUuXmO
ftF7oPNx7183BN6ROEhTY7P2NiAdMmFLD8w5exhaCez7kW1L2sFW0SMen1Yj61LY
sJjICU2rw6znsojsW7J697H4yxh5bDyFVNfOinGTTaj5+UTYwjX3WWIHbIsEzZcd
S9JfmfX4RNcoJREUiyiqvkbFAfRa4wyfSRF9ratHmWA=
`protect END_PROTECTED
