`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hHfHPWmTHakyghotMNFXLJWh/xKcGCSMAuYQDwmrgNSEypEosCgfiZ4MzV5rscAt
bNiELWbwHOJV0057PADhmHiFr6Mk9HSvxSoynR7CdYG/+aT+egPLUetkb05kvy79
w41MwMYMUW0Nhck2fQuvqxtyqddySt3xhidIrd1Ms9bGmaePntmVtDZscvaCG+Xf
+fxfAWyn2KJcL1oufgZ6qHdy01w7fC90j24yKHfeBcgGJ9vCRi+tlSWZ1ggXRVBc
4TmnllrsgP+ldde6MQBGbvcvZWgpuAuDdutrd58H+NG4L+ddDQRutzO4dVrjI2ML
AxInnj/t+lIqNnSkp5YSCP7UieWXiCGUUeoQOt79188hZuK6OOA5wfm/m5WvcCyY
6lcWLMtyuq48tBHDsZ5hv8lf9lac7I06kJ9fpaax2Kgk0sw2V/c8AFKVK1cieghh
oeOBuqu9cIPpGrh1uK9HkWwEUWvmedB0bBvFoPw8UCkol0mc+Mbi//zO4dRz3C+x
`protect END_PROTECTED
