`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iEjpgNVp/C+EajH5+HydR8MTg8+THkCidbLJeEGaRmXXxgUJu/oBnUanD4rtfSgh
d9WIqAVrQQqG+ydH8gU52Phx9+PPjTbedSmqq1l/Qwh21B1DP+0K4e9n2uTDe0Ez
3ltcf9nYVmBKbfTYiZNIaKSESNRKu02Fyb/+1PAS9nrIbLLIsaZ6ok5NNkJRlxWL
5DHvR6lqZ8IAb3Vm5Zil85rFPPf2T3T+PJF0RVeE+v42SszRr7OKXKz7WQi7M+3m
smkT35H8ZyKvOMLRfiSSvhCElqCfHUxo2QbYMLpo5oMYkb9c+AF1xVcuZNogPyDb
D9VKKqO9NUkem071LPxEHPNwQyk3TxXgVyWVZcNiqHwClH+DrWbmvRkc6B7yLKEA
ultqk2Hly6LI0SZauXG48ZwbGh3BpY4yNG2bR0ObyCExvNGBLmeEXzbbH6So5/qQ
mM2ID6LrKye0ucN8DNxWkHJ2w23G4jR/oM9HvXymvDZeWybAZ7Vn4Yk42UUgFO7g
nnvY62hHNbEWGuoK8oPkQeI1WyLGLZp2MwtnIuwxGSeORIVWT/6nWAKH7133lGfR
RlFQtNFqIFT0NgYKZXlcSCa2HcUofbCxU2z4VV/gLrOdK4cy2LuZJCRQaK5g1V1A
qSNr+09Rwr+Z5QKLhJCTLnpXlLvIX0CzZAL+RrU1uunbVFRrk6/0ZaAHuHgDwcAy
s1k/Cr1XdKNxXyclg23HL81h7AX1tkrDbsmdG262N4BECCEXW3KIZMMCEd5/qGKf
gx7hhtmLbkgGgVnG5fUsAwD2GGmTxN/k/26Ye9hsKQ64RZtBvjr0yI/+E4lFVOSN
hvGMAeyBcLUroBmAH+7BQ/3LP9TI5H0eRR5VHmMym6ayLWbUkKfY+MDVswOW4PqP
yLRg85Y8AgGu3RelYM4BalWoGwW1DWmnsHsS7lM9FrSJgHEJlKq+ORUxNWTS5PGC
CCahyVTrPsSSyDq3vnMSkvKrPO+Je+ufFr+tTCbVNtMCroMFRYTm1bIEcAzhMVpp
NTbhhZ7UlSn0jRLbv5Ml1XgFhJ4S3jEGMS1cBOqElwOrKk+J+lXX+si9s84RDmjD
7iOni18VPvQMnMImMS19axO0o0wU4MX+7oSUwiTkSzTZahr6lw+aLwjJXdqLvoqF
Vx/YCHXo15iJsQcqE+phGPkHUdhRX1/I+YzSTTotJAzXL4pjJghT99LGLVF5xxRJ
goEPOec5VBkzSzpsB+6qIjWhrotEmqfo6vSQeXNdAVAOyesm2mkzbuNLhIs17qxj
jdHZRWBfBLsY2Zx64S2UbpWbpDzqRSJJuujxfAfYaQarvgnk7MgJbB4+9Eb3GpYG
O2s1+JHLdZhbCk6vi4oIChHAZSydEnIehuld7D8NCAmw8k0+qJMPv88dIu/EUSpD
zoyXoLOUIBwKNxYnKvRCf95Xp+rLbtQcCQ7O9085w7duH6y3XwTnq5nVSQwOzsjo
n63HbcwTVVoTr3PrS0nBLzBM71zZvNd/6/l0JNLx7+3oPilQG7FM+UthSOXrf5kX
hR0NvHNwXuRvWlBQX8ADJF/oEbqmm+5XTvV56Q2cHOq8mm3s6Fgc1whH3d1x3wC4
sZFYS9eFr1ebrep29s8ueJots//ZdVA41u+jGgA3yCezo8l391G6xe/5vUuTbnea
TqSoYHK5GMoC+zqxgNaHlehjRSm1xgL6cqLy36Wov8XWkddVcRM76eZ5/4YyY6zl
UNLmpnCqlFXuuDKvoAVGrExRk2Tk3CxJFb76/jSGr81ysicNRXKzovGuwczW/inb
4UmfpnbbSmIjbR8jzwCqm/qyViDq5iR8slqW4M1j3A3Fn7/NGUdZyCYmY2rQmFCM
OX57uprzKSTry43tjSyEo71OzEAAgDB+pqBOV7N6SBKYC6xJGhjmPZsdh6gE20Sz
jyh2QFZF+ZfRlJFgVJp610rabFXNSvRdGQ3S4lhU44h11ZGy0dTHoOQdwF/fcs9Z
9apbtPYjR4Mlk/8c/dotpIayeueIZozivcMoxKh6QT96RUdSBeHDGok3UE1FBrIY
4HpXB3XWROvU4eJh4CWvTWAktfPCmk1WH4WVBKPjlFMjYpdT0Vxr2BAL5hhE6qmU
eZqXX9pUgfIWP7kmOcoUt5zUdV7J6B2XLF6Hy6iKeDr3DpYZcN1ds+sIhl00gkxA
vIDtANtIyfP/P44I8HDkcl6k8PTkv0TqELZ4e+hcXEbKy6r6ffvi4z8dti4Ifwps
1VsAe7bwjleQvDLVuOkQxzvt3T3HC5sZ3S50K1v1MV6MUBhGHDjUcBRw7Sf1WC8K
XNkIw+BjbLd5p3IWXQGzQ05M10VT3gY4351vuBQurK6NQb/KHzAQNr7gDUY0XYQQ
sk3nmxUgsabhAIXWLW9MQstaJZng9Vcac+Cdxq6XvZmq99lbczsLG5v1+sForlxH
T8A8XeVpPi2Yy9ofyvkrZNiZCa4WogHduogKTe08GodLxitYGVAhj68icrw1vdcf
8U8GrZ2y+cD21BWESIUMC9tDgG7/oR5CwCZMZnaL4vtbEoW85mEYJnIToE5BOmKs
TBdGPC2RuWL3gLu97htqvyDNsYUJeS4IZ4zob5G4U0rhFqBYCca5S/u548IPnhVW
A/eNQj4FYQ73lZ6CAPjyks0EjQvVcmIMOb8Mx72CX5uVgeosrqXbNyVNMIsQVnNv
42WNGL7/CWlc4/220sN7LLwgvgEanyIn4Jl+9bK7s8xWU+f/Suu90IsNCX24JlhF
Kg98aj24Ik3/YE2pF/4ufbeu4z4wF6LOmRUBo+k2nnJmqDITmMtS9jZAwjJlqozV
J9PJMV64mrnDwuS0eUyANgOWzbT7/PrTV1/sG0kSchxDq+fJuPpren4ZmK8PhHoi
Lpk7TQEwwMKWZxGzSiLj02/mAiv0Qloe14aZVgVq3R6jG3mUi+ypXXPOGWR4cIQf
uNG36vEyMTZVnCaP1nTif+w0mPGs5joTMgEQtrJ4yiJAQQV5mm8CTG5PLIEwEu81
/0lseS459heMoHYBdU50nN2frk9eWkhUTmuuM0rqI1B2Tdi/1MlUZCskBSgo2+1P
2sc+0WmOEU3lvGjWC2JxS62Dj+cAOrn//yWjo5CvqAaI1oLIDDng2pNND5iOE+7m
AxQDi8qFV7HWgDbNjWooAK28QONT8fSF6quMygf8A8SmN5BmF/sEgvGTzSmDMqCY
GDuGsCynkuwUfVM4vWXHJCEel1X6hifjK0YNdkWc/VUI0q8QpfxGsXrroOqqvI6d
XTAEmr7jkarx/y/u5oA4ArhOkGR2NM9lIrbMvj9x1OQwTMP8HWaRnVOLgsVB/i7X
`protect END_PROTECTED
