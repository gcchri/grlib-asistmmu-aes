`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aa2ZXPzZk+/UQ59q91mv/Hfkp4NqQEqi2fK9Bks+KOjQLazQv/4xINvBF3Ri/72q
Rtbxqi3ypdMv+yxiW2CfWGMJ6HToj284uFtukrNsZ8/vh12L1XfIDEXqUQSNrDpl
858hxmyfyU6HvVIm6DXNfd4/4ANDpGiLgbbAgsxieUdl7q3bZHBvuL/Z7PbnwrS3
sVOL1mQBcJLMPj2W0H13LpecLaIrEItg7eu0FbbzxNyB/UNEF+4NOBGlDPbMI7NT
001nIeGBPAxxGmNocUgFSlUBl1EJ72eXFZUJkfUfvM71UNhhPej3ZLRlzALHKn41
2CykdxH4eFUpi9Z87DROsVuxwKnwNz6ytlXuybH8a24lAzwm9m8RVIko3I9nQFCk
K+wIRxtvOuWwjJJRwSK/19LGDiyxTPj1qV/kK//c6JY1uzmzUj64thhWiuqBw50w
+BtB8aDfYBGWQ/YgDa0Ywwf2LzROHw5NzfN7vx2gZebG5vY9IrNELZbnCarZxpU6
t4+uUTiWnkohlz37EOnyDWya2tFz0BZtQ/4MkKgdcfIwDanVw4KNYZdU4RhCEBJC
81NkhvSH+7J9MiQsGPDQfV3MvoVq7qsMfYsbXfe6NqFJKJq91Adj5vvaOavFsKJ/
tQihvxF7iT6CRvFQCDO4+SVrTkd2tJNQcobFjU7CF6Z6mFantSDZZG2UhGRSdKaV
DysRn9Uh5Z20lSO5JaVoVTV7wmigqokzmI0yZmXnAFNZDFoVEhDoDAku4LS1ypEZ
2+z6Pmwgx4dJtm4IVuZApdR1JdYKFadOIIlqFN/6wEvqdfQdswgoTZkpJTQjnwJ5
d0ELkUMg0Pe43bDpfCka7e1JPqBeBvDCzB1952dUSm9P+VlEj407JCVB0GHCJwVc
7wusKNWv7cOBHFs5lg9iP+b/15dXLPpuq+3JM9UvWBqVrDPnCIrvUngt/XYN0IBA
Px7dcJ4TX2zbjSV4sGcoEkWONhNT5E16pCJNCWcgwgC1q9uGNb9csiUErzZieVFr
PFzylWtzh+ELw/f8HTHdDAebKDdJoRC9vny0mXhiLLVyTumBOpoex4vK6hYiq4aP
q4oOp9ECDiX+jMFA/bBG8WZE5M+J5cfIHWCcj3eRqh1qGdWuYfNL5rNM6t1F/Ewl
z8LV/zT+uG1dzhxWthPt9R1vaMtvv6Bj2mShsJQjSvaPd0OlAOhmexHoWp6darR/
jF0Qku/mtKeAjKme5OZh6cpz3gMRPcUfQV2viJWL38+cbT8aMFFNxW5AF/c41eaj
`protect END_PROTECTED
