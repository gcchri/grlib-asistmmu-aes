`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NkuyW4F8cg38XA2dTMHgqgwKeebUQ6oSBRlvDncFGGa32cmqbUZlyZecA2yGN5pn
Yq8GizUQtroD3pr6caD96Ov36Qt5KVLTndLYS4hppKZkdQgL9UzxA4cD7cnlbJMj
g2+abUtm+JfbJFUs12wQceF/5HzB+E5jk29XuHz78mPvT+8/UZWp2ASBKcD5Iaph
taC4A5sjZN6fY/CMBTxG29aUD1XNH18tFk8+RqkT0M4GCSf1tAYJ+XiAYRmlucJs
2fYRFGN4grb0XWY/QJnBSA==
`protect END_PROTECTED
