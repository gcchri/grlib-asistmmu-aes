`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w8JGdswy3edsq4h884FD//wPdHaQFr4o5oHY7YoVs4AMqFpeiWW0P3vec5XYhL/D
RfpJItpdRqPLTET7ZBvXcpq5mOH21xhl/gurppafD+3Z9zIjXQUGl1L5PF2Z0IyF
nGI5CxZYCB3l5AtJ3mf/GE9/hMGtw78ZozL4PaWOvrxO8tEL9Rp5+VDg6KY/CVWy
zto/Q6WcoKXt7Tb3Rl7GIFltsKIuzW0E+0fPn2NJ9pU+kwSLy+7KHAgzLWCU+bK5
rTgxUrTcf8S44CoGfTcIw8dn/yzVQ1Zps7nF2+oreBfT5IrKSwTTqAevXB657Vns
vV82g623tE9jvhPnbULbZw==
`protect END_PROTECTED
