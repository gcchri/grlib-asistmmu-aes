`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GM/6f9r5KoXAOf+/t9Wedw3097VnL9/CVDtkRx/E7qMbgzVSfJhQW6Nl13+47LxS
36f8C6zozw0jPkW13BsKYTOM5icV1pdfZBEdb6FUKQ42JjplzpKSMk01gXrdiUct
PVieyQEtu4K+cBakaUZLDJqA1FjGXtuD5/FQuFQ1w2cy9mK4B6x37bOdLlX2DTyq
Owqxg/c3TG1WdONqNIXk0/199BxRUQ0n7Ytf04NJBrdTrYaVnIuKaeagR5WkJe+8
RAqsxJMKcOstT6Lh+BKef170XSR1fLNGZBD367MRvCVdsB2++ZylGXrviLiXpJXl
3pFGBuaD5Q1Tu3uhkOuhJj8RKt51I+72o3Gko/cFkbWE0hm3frqQlQ6j2YqgCd90
bH1BFB0ocoMWzPpEijlaLuXhXsyeEMiFsXirgf+c233pLEISpuEiKf11k7h057ep
dRezgb2vXzcTUmMQB977+TD9irjAzu0l7Q04acPDnF5F43uTvwlZiv+/6FOqQsPX
JtJr5j1s//gNwIAppeYjAPxqe3iBlOa6MsYS672b8VCiKKSrqIyFKGfox+3ToHEV
o7QIkfadIbxg7h2aNeDLS2NfCe6RpnzZ2zZidW4iqVK0a5pU9kqt8+M6OzUOnFz/
xW3Y/BEU448b8WWYw0UsYw==
`protect END_PROTECTED
