`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ATQM9+ACxjyxdMoMa0b5GHQyGaLokBleK+QqeiA+GzSSU/gGFtR0aBoKEbhGnWnF
J1I3XcI82zZ+7tzTAP3S5kD0FetCjOT2CaQhW+SlywFdF2fIMOkIxmc0wrJLROzN
Re5rZCDI7ySVDexJt9PVthnJT6g2xdCdpNdmSnrN2zgEsOzbRvmwST3/BNIX9rBN
8EIBAsonc60BQhjV2C1G0fVrNrW91/24ylN/r3+Kri3wgyZ/XH5y6h3C2smxSVTD
Qfnh2n30xvDJLOkGk4F/UsH4XkkN6iUNoSoKX/8XSleU3As6s5WbilpsdJJdVba3
rX+DwSMhPc3arluka+Ph5/tLJWuwMFZufP1pvA/tFA27tX/o+o3QySoQmfvV739y
v5xjdTK4OIv1E1fLzw8DeuLNO7uAPwL08trXyR7D+ZltOSbSC1mMAfgro2TfGDkY
gT392BEZlgHQ4vj3Hu2NjvTI4qUsU+xCQEnmA+grRYg=
`protect END_PROTECTED
