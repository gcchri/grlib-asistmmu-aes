`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C2FVLm/iuB554JSnDq1Xbc/JuNeMisC2hBm1cPk47pAo6P+41RNBQZXIGhrtTI7o
lDf4Nq1Y93Vf+4+ZAJBf60pef2b3YezADc756EgFuUW/5CcjmQPBmHo7/MGsiLVE
Bb13QBbGC0Xh26emshZCVNOwkXKsyjqytjJgd2+wk/fWaSAj6gyDDIT5mB4Lfsbk
/Ev7axjRKEKyjtbt57SWX8Sc5XcEVsd3ZaIRCtL/c2jY7eCTcJ9DJu3UZF1aS/dp
rlCxOVO+0eFV47Xr2mx3T2sIyzz1uF3JHhFkyTo+n5fILUV4MVrSR4PxVOaXiusZ
KOln2ZrKTBEQ7mBRr/sipGNc0Ql2OM3kC0V486ujBro=
`protect END_PROTECTED
