`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qdOB3XcvnpHGfUvRvh91S8oNa8p3fIlS2nO8Qd9HgHPjRl/UKWmgZlz4EtYxVHY9
XNPpeZADQJ/SPxLyNpvmfi/oyBjC6umfmogZRV2oRLh81q3/cMzj/RIfsm/UKsSs
27B4VdWkA80+sNpZ2exD8tqJuPrJptmmGlbbk3l6QlfcULW3T7ke8AUmvFoh7c84
Jhhmswtdlr7rhOYml0+C9Bi93pWDQbWUQM0REiIgHSMXduCR4WbiXzDxf896dywU
fosU6xrDoonr5ohNrPd4Ymh21HWk1TH6QmKMK/Opqko7ozPiGvBiQxvnq+IagPtp
srfNHbz2DgVMIRg/X0MqYSX2MNCyBmwwgUqvm05wyd0lMgrbCQD4A+CntTgADBqu
9vNg75lPFbgzEEKfh6H7Qm5H2uoGt1MuJytS20pXOeABsDq0Caw7AuQWA9InjDQF
v3EhaT1wjkUNJvWM0GwWK113YCX+xp83KyPPf5NOgrDfFt6ORdzh8zTOBY7Tr8Am
JjxgBR8moJZ/RZby61jDmWW3lRz+FQaG+vfEIcOGl88NFLeaC1K7lCUMZxfV+U8Y
zWA8qnOMTObKNlTFTKVR1QJziUvh/s1AXcz/VvxpodCYm8iTzLJlK8EbKJLqCLFs
LBFqrD7EZL1T4e734ex0C78jUbfIenkhBYWY0FD3V7QrgkwD7XciUgREZ4h5o+mb
aa3D9cp9d8xwnRfmhPkHnAIxAzXzp7rV/nqvscNPwFiwEGucTlzBkchQtX1m+Ru8
a1HXTWQ5CcI8V7ETP5e/E9oXv3+3KXoFY65FSMu3XxnYw1a1753eXqT11bWgFc0q
qs0Ikx9qjQe66QYQOn57VLwHh4TfZY19MBTjypI4KfdHRU8m/cphc62/gyL+J0NK
7O6B5tHgmrMiwh+Rrdnkkmida0cZWhpveBWeRrcyq8pNtQ9llUni3QfcX2rDMUKQ
Kc03bTDO1m/IljXoX12qlZGAuZ5wuRmqr/9PgNABUNpfrs2EGvc7Xleuel8HXRwg
1iKU+W7YA+2YLsIgi7NWHeZ3U484KI/VmG12puGf9DxkyvbMT7nlEA8QxFcdOon/
ZlomOZ/PrECKSRdMmvBk7iN8/57hwk6qz1ZXQLOVd+OB0bXpxM9refMfZt4wkT2c
ZdBBBlHqQ2yUKjSiu8mtXtQpOHEH6ixfadtqlh0tl3DpU4V2fUC1a1pA8G4uoEdz
MWOtZq/8glAWS4IHZq4TSlJR0YBlieTteWoKqktWB7mqJUwgteici/YxTHvMafPs
IXO+oj+/4WaUACiPUNran3Pm8qVSKL6ZZLA9xxxKoJWq0T+mEv/LJAM6ETw0nJyG
9KDiqX6PeolAicr13D5qSEy+Zxv8YBGbY49Rq/Zvm0OgmXmtPMt2ub5mF8yw/iaa
/B065Y2GzEWwWc0xDX6SiH2LoQg5iOvXCuLTnNmIZqoYBQy8LsA+vr9M7hiuFeqe
iHV1Jh5CYlUuN0z0qont8mp3ZZXp/xt5eVn/75smcCnVJO5vkURIJVAMSbE/p/+g
NnZp0s8hWY7nf9QToSlWP1gFJcCu5NasO04zDmEGoWnhHm9CMis8WVhucwy2Dk06
IiOTEfeRBjwkqpqSc3oBTqfcxtv69CnKXWNeotnij8fVMCfPcElj+CoAOHD65LHK
muoaZ7AFnaOYtqJA7GOt8XOY77IAFQHLzrBV/yg41fSsAoxSiN1tRGtE6OH4lr0E
8NyxpdSGr1ksas7B7/2iKiyJs2bPUJhKaLIQNMy2GhMtEhkT0aNS7Z/GP8OztJg2
vCmeK7NJ9oyv+5yhQMZBozftr3x7uI2maaJ7SdQIckiUItWy01Kiplnfj7BsPn5r
w2bdkl0pY9cCCoWjXKDxCTEWPt5S+rHCRXSSYSiT3DUWA1tpqUcca1s2owjmJZiS
YNe8MuVnJCJrAsAo8HzF/ITIeB02AnRQ8/gA50tvCIl9XErRDlKi7esMOsNwA6qk
G63/v5mzs0gS7pAt3VtecAmUH+DHbw+DDvSE3CrU/fV1DKmUYYho6f7RopllAuRe
iGp6MNEv/j9kYT+7R+ynpmyZZgaNk/Vkc/+4Az81B6JJrwDZHcNfFnSkCIwOvERN
qfx3QY/vP+bap8KDFWHgRctzFdfaCJqZ+aoB6KnrSlCKQjPARXJD5fNGzMMJQ4nk
SJl4/yrtF9dV2AhhenJL3kZQMfgjvlXiC7HACS4py1XHKtiAja5EPAaApWOboxCE
v8mVoo6f6l5rpUvCGtFstkdPCHyxc2+mUbLliV4SRaTeKtx6nC9A5QOihyo/VEtm
eWbe6ZgLgOIfAevavEpKX9afZ5tmtKlNPO+ya9Lq5ir0zD9CCAVCkc8kkYTvOIHM
fj3ynbst5bkmvGFnyl3joDKf+pu1n3kWkqnt2tM9+Xp+4aDlmuJAUxiUVtkErl0u
FyUbF7eXl3JOCdzjv9Vcf8iDB8tHqNX5ccJhNWlSQu6JDrrYr27393c7kmpanLS4
I3yA6swol6jPfrFVUmLKJwZbkwWfYKrKAq/jVYnj8U+Mrt7BeFDtIaLM1XH/sQSN
CTp7KGFtepKSpyakVfHhu+L9E6Y1DO2NMgM072mHsYXC347SIs0Gzbl3UU3T5vnR
RcXCKE4iYc03BLKDdWQ0OyxhLENRYrArjVRE00LqqZya+w4pHz933k83G01Kdibw
BdDv/c0RK2AwM6/9R4Yv6DUOPaEd0vc/pTK4pBm2wB/uthibV7pYm6yuR88NEm1C
YOPbPJmcz/1a3mObV4Vw6ydzfirRX5wurIjRw63uc5Rb6zQ1rVE/8P6voLohFqIq
r1wYOIGfUsWaRQOHVU6HUH+R5gngXQqEiYdBvgQVCDN7bJxjpCK/tHc6eR3Ui+zN
moIdEbvOrGH+kFLYCSxSIEgz7zdOfb9wtFiuJgfDv539thd1xj+/m6pBa3+hMiV2
aMCE8OXrQTm3CCC3zVG1nOcFFfZlFuxi1vfXxWNmLSYmxCQcy2f26URXJO/XuhXS
CaYKGs7kKGv+9W2ZgPt1Xx/ntLwXP5g3NJIcyurqL/wlVrJwCLxyi9BMlE0ctZqX
RFItdrAegfsr3ySfnKtQ9zkNII0lV/W6Lo/k4y5xnIQQP9wD+7Psn+9hRPC646d7
6G9fVEBIJybKCHaHbkje8kcFfB+eCJJunEcwyysREPoDV4bcaSHY+RqxzzMI377e
t7rfhBxITNLXyRVEHD634CVWJykHKWLtVam0lgeOLeZXlyAZqlhX00OqK96MXVqy
hyHryCGVtR24gJiq7lxKieibg9IV58BniXiCbwVG7+Rd2flib8zSq9B/X1IQYsU8
rC/ytgCF5DjIEMJ/WoBJzv1qeuvGCwNn4LaDspC5YtP0LH9OLwk484wrL0GVRbtQ
aK9uuhk/gf0bl0qOXgs9vqOs9+xKEpWx0czIr/QFoNU3jLMzH1RzoBs2jhgt3mjZ
zXhQgbso76L+/1D7bJ/jxES4J1YaPrZf5nGHiD+Yv91XV0/3wcTpmk6I0Igrg5DP
zbqyyPMWYuWtaaJp9hvgRRxK0sCDV0JEjNopKHPNZs8zPqWMEDR8Xl76prZGm/9k
OTk7U3s1u+LGUu0yJK6ECoxD0sC1HWCgsa3VdVhPMG95bGF+m6zVz1naeVBiiigq
+yqOtqj+MTDptUOpMsFz07YxyLEgKCVkipqGbGhVLjKp3zgOVUZrR2eAbPaLwb4f
DNRCsASL9L/DUZViVKdV0C/nyS79fM97MGr4CIbPwELihzKnnwmO8WVB4c6w2Q3d
lvuvscjVqZ+1dm94HNckQJyn5IWzc7YOMBJOGHDM2CmVXfjNibrc7sZVoRoQvlwl
D7S3LWm8OEbMj2QigEnCoqlFw2eNL47SvstSZDD8nZ19fAsRzEkkUs5oiCvyp2w/
FcSs1QgWK7Lxe2xYowRkJ+XoPX/KvkHN9UOjU7RCPboz26zm528TogMrz0KvF/qR
7RpszXdlzC5a7927W7oxDGTgVcvInDKNR2twnh3O6guegzvse0Wnwk1X7QkttSa0
cE3v/FzNR/8+EjGavetRGBE7sH6gCAqjJQLUi9dh7DLABR/8zwupUNoZiyRujVU3
PrOSJsNWhoI/c6ep/HkF/lRbvXox47Ac4FTB9J6aVMIUw6jNrov/q1Wj+erw61HT
srjLldoJ+srCL3C8XDw63zAv2BTNnvHb2hdx6kw2+8/PImH5bx4MYMy6/Lp2whsj
M2bcOyaHVvGGEPxIKt5XOiMG7+7KFgrTcrd8mb+SRZeFUnfj7Dzyl7ejZwp7bA4x
/gG06vhwketJYzFKoC6Gd1JO2dd9dUlptjsKQehlg4sQ5sLwASRxMpzT0MksVyN6
0S5Vq5i1VcCdog/dat5GpdMNiINQDysYYtl5zvEhNszceBPVTeE7t2nWc0po4k9e
DkQGXxWZn7w489UYS413qYrZ/oKjpRtKBGt2/I4tvIfDhYUy7xxM+XFGW9A/SQPM
ebGTPicZf3J1DMjCB1UqsJ7xTPT2GUNIbIZb0RSDarmuqnPjF3NRkfZCfHSZraTS
LKHSboH7s+IJfOFG6nyl5EezbrZ5eZvDiEVjQYZgx4TShlVO1OjhR7kP3RswNjER
AgxNzBxkyWzjfGyELjL+CIdwLb57Z1j2ozAhd2jxd/mrs67gLDfgJRpBwEeoRtxj
o15bC8eeCmC+qF/cdW6XSnucFj4qWkKmiCWSD0O6g6DNWYgX7VvP0aEopwlMaHWb
W2zJAshHz+1IgNeB6jASlJwi8gRlAHagXQd2YuZ7aCGDm8DtwBo1413z0bjZW2yv
Zp+NldnhwlXEFR0hHelXhQhOAYbrKiWDp3reRcdHcH62sSKOlRhgmYyKu0eBcstW
rQ0JPFRZNUmIbhOUtUZufw7l4TX3JgN29/VccObkripnYyhsAjjoL1+GT3vaoWGw
pzSF2PbPMGu112YDLiPs5ilwFyyJcYoTcvIZAM5/BxtMIMnABZOM8jTpVWq08jIk
8YiHDiGU+8f0QEIjGLTwMWSfNZF/0eg3BkQVDzhY792jvsCDgFOY2FzVQ/6G1Iok
6G4LwuPzRgNkB+wEpGJYnVaB+ysxtCeTzthkq/H8vYhG93dIyq3laz0/EAM5S1Lw
rjfkSPzKeh6m560OIe+q3uVVE8rTDl5mbGw2rs58R4kecsgPf/dSfP5Cf27NR8TO
1Ztp6t/KaV5F9gZdRSHKlSfR3PZ0VqwHo1mkZEp7/nrxS1qSK0w89vJTSAABMw66
h/QhelHtYjBBRsVzombb+dMNzP6gj5hOs+lCx62z5ozlGBIkXU+iFgoSqknpEz4+
bAyWN5oAAGaD85lkUwI2dFnjn9XnRJKznSftSqzlBldfkFAvzR20FSO0KD63sV9n
rx2RYZikmuyyvY/2h2aAsZGIF9Bo/nEEFAbd9VQiLiM2+Rholp80ugHH8tFCrxUB
Ci4TQB0IEsdADBDbvLsgAZFoJqn+QcOUSBYYenrpUmpiuaR2qIx2uRu41IXdjMpc
Ag3a3fe1iFjT3hcGeF6qI9GmcDlQKGrAgkT8ikceCcbdtMtZUd+YYjU9MEiax+SS
wmbwrbteMACKkgc3rngWwnynLru6T0DPXSIgZEEiWH7McN23KwsOY+7JELEHld9R
D6WPj0wUDTYzKaHLTLOpdLU34qeFvipY8+EMzoMH9Xz//et+t7h2AZ7mDLmWmS6q
usTi+v7c8Hx+hmqYhbiAmCMz04EfCm1qsXMSTjnQnhnBQfrNu4c7JywX7hG57QP5
pKZLYtyzJwARgw7C1DpBWYbhnDpgd4k/a2/j3S+572Y8Dx4Q6/aaB5FSLFsSlViX
tJPmCMWKqiWmVNu8Yxlx9oPs0LH8nkNyyZNCujKYkNWQmBlazn/SEx2/6vaMemOE
iwEyMtyh7ZzwCaGjjcankRx82h9WzLiRcDZK99bdx7ocftGPjXczlW1SCsOhRPuE
qYRg43uZHHX33DSaYGOYG3/pJA0KKqb42u8tu5Xy+a7Iy8JYCKtsDXsD3K0LTBKP
JK/cPs+NgECNP34XN7MZ60tb6E/keG3fs7CdI7jQ7Q2NOPXCCbdOof5evTveyzPc
GBDS0dvtp+tadkLhRu4dSD4TCwB+5PtV3sSlIAjUbhh0ZyofSkhDf5D7YLwculkj
hNJEXPWe+ucrv1vPl7gEir2M5vOAY5Ol3EIO529Ho9dH1xWrtXbiTkWQBlSCWZns
KN1oK3HsT1/S3mtiTg0WVby9ijQ9GMdRK3Woy+yn08f8RZPP7F9WE9yL6devIhHG
qmo69I4d313afE121CVy7WmXzvLCnrGl8U72dnQ/mfz7zgjf5k5oc4QHMAlyE90Z
8mImG6h/MaaN95on+b7DczHtzQMmBdqQLOW+g9bHX2/mgv0oG+jw0Ai+Qlx3MKdm
OXU5JXpM6ujD02eFopcHx/2FZx50gMKFigto0SFpTaw3GuPq2+tnSHN3w8k5uVNy
aBgaJWzBlwXIe36Y2EO/fQ7ugKvhH2Bu5siGfmPOQtlAwWLQdl+7QWcIOgQkplk1
1xRnxZ1Jxw+kOar2dfHc927oeOb8+b9TRKX6AWLFkA2JPTNHHDz/UTbXw9RMblI+
wOmjInJQpIZPv8EIk+W7Ri50di7Lz3nsCaRNRa0mGdFI4FBicpaxI70vX/UydcNL
T4wchaon6wDFpcnfTSmYOXWua8091p8odMNoB79byxO6DfbRr3lbEoxenBTDHjMI
YOZ5tMr7fOlrCu6YVca+Pq8Vl+oWLF0WPGk2Ansc9IRNi0oGjpSflsc+T2NiUB+q
RyiOAUx1ggVe+PHONafUs39SjZl3K7nX4HVaYSVMiYHqzBQ9msNUGREwG/62Clbd
ukGN/mr85Lf/ZCQBHth6KdKX5vptrmr8vs2cRWvJaA9lGJUpkQPMXGpiMrYxp6YF
zvFtUoBFbR1jqo5zB6tt3Sf657d9wblUbpyufGXktvibIt8k+sRTq+m2vR8dpHWL
Kri5rkTrV8pyEjDgQG8vFwL0fVOh7Omqv1mrrE9m+QRsEd0YXb9GjKfpbm/+Hbod
u4OFEoErhobq4zZPgiZ9p2sI30t5DdEghaz8B+um1P7JtZ2QJIftYwig3iMIs320
MikdnBnqsQC/T25Iubvytogz6V75W9O5fjzd+yu2QpzQR8zkUQcI01QEgG+RlqkK
Eziy82dbljyqRcgqeOQGB5QdnfoBMcJAZiicwmLytfI6CJROsSZl7ym8bjcsofyZ
0fLlEeNUUea7JhRas3kaEGDseL9RFPnJut1yyO3Wr1dqMnCLWVMU12XYPrHms8Li
SgNslPhqITLJTjgZKPZ1u3a/2VxDQf35EBwDConpQwXQBgIC15HRZslW5zI+V2ag
wNeMuAN2KJhTlnVI/bbAJjqH/3I3GgXmasfyXOLXoxwluyG3mzvTdXr0mLA0qp4k
/uqY5eY1I+dZXnr7TRiHRzogLdsAKw1b6LfDvaKYLylTnUvDxudhfT9OSfwN8CwB
XMqpgDlwr3JWTQfiLYrfqetM73IWf8hdiNnHkTJW5W5tYndKmAdzkAvqhBXCxDkV
R783C4zomQoR8mWz2BZO+IOTqyqyRjoNdm/PvYEd6QKZbdc/VYFXjoSF4MmEHgdt
cB+jQBj9yLymqIFULNB40ZVIuzjBMBVfdWt2d5pz0I0Srpa5X/hVmba1O0kKuf48
2iRgOUrsZvYCcNUIUVYaBJ/JJYTL5DxMmU9LPhzQ6CIocf48a5jYotJ8LoN/0lbq
yqOO2DTTZRhR3wDBd7Q1C1luJVjDtrxGXiW8hpW8FmnZc+7SlqVZU7iXKOEW4F+R
s+AfpiKl5almJ6wWt9J7gPQDakSzxwKAYYa+Vd5XclegVQngGSfsF/JOHqV09I/7
XhUqy2VbMiB9IFX5SAbxhN5h3Edjm1rbFwJpnVDX9yBiLsx3ooOUMv11XY0r5uf5
9RRMeikxw51H044moXjEKbFZ4M+8t7ezU/ufWRHldKeVsxkUIg/E9YlbpU35gBNT
/gDsqJRuUN8sytORsXe0GwLlKaqo0SbdbBkUSxyIAIhQehaM1Ii03HT6mTAWJROL
PAfLl6Khp3Q4TeY9rOcr0dHHXDyN/0H6mGISOYpjyip3bM3yZFroWdmXfQKH0bYc
XXTpGd7+ksJpF80LZiOVyGh9T+NzIMnbz2IPw6ya3RRiVJshqPeE3fFfvGAK0kLj
cwSbvxj/srWbKoKw55PxYhRvEb/meNrt7tCSdi6ibmexPH0pSHPzEBUfNpfdyYWz
CiZxDxW1R7Ssxf8ldjvYYGr1c1bDjXQMRwuOH/oGkWegr1t/O8VJoF7CIltFR2iG
z+hJnIK6AVD/EwcObC7CXXyM1JX3H8VsajDel4yTK1p7H11D2dyPTkPAIuRmG+h/
uVLk3jMGORvk8XSRNG9kp7zpUPzE7Cr938zn7NSgL/6fFGvJZk3PHU5M3K5wZQAP
DHkFwuevJKQDzuHP9HXLJo4AdblXIS1tuSMgtmOAigaMW3JcZ0QfBGOAy+LUioI7
PcFXSqgj9VtnohdSQwB27jc/cuqZbpV/VaOsmosG7SLAn4+Qp+xe9PGBF1ctRUzB
CwMo2zRPwFICJJaYo/VKz4x59WlJUnfARECxWA7ExjC7TXqLTPorkMWb/ijAg3eS
Ok2hluftJDP8W15Enkd1j0GMkcTIYfcv8fp9saA7IZTlgY75ODVst+07OnuPszzz
hcNMEy+OH3J4GLjkxbgxDKMwM7tTTC0n76YoqEnHysfkZleDzPbI53tuSpPr8G+S
BHmc02Feg/hiTCHprmzGlCuLzfLx0oU+9kVoceOe3jXHpVh4KoTAI1Lc79tNKhL7
xbAwqRAGgLFlxnUgGoRD0Q==
`protect END_PROTECTED
