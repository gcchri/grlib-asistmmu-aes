`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KZMQmzdByzWKOEDCdqXnrP5E3S+j6IqV0mMo1E7WCNv9mhaXUUnmWj5ExIrG67No
guoXMWTLlk2Nhlj/+Q6PV4HLeT0/nChdSvkgqzGiuda8Bsl9MJ2S0q2PMUiir5EJ
E4LfPOxtEslR7x3OAjb8/agq3zKdbok9+eASYwUa6c/H9PYqDvn7jGnLfvgpLIO9
uzlsJDRlIBDvPTAh8vBIAS44z4Myju5makPTPPjK55zBoTj4yX+ugSvxnp3pGfA/
oMlnnqAznBWrrY+XVPdVuXF/v9+11u+w3ArRaCCCai1EGyELUGM521/h7gRToGjp
aGXBfmqgfVZEbPKYLEwZ6p/1hR+h3dCGk1jL5jOVfJQ=
`protect END_PROTECTED
