`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cNPHF8UDTFehnVe/e4tOFJHt/lEzANr+KFKUn3GaUaVsllrRa7VvZFXIS00EDd/8
wUQGT7XKk0ctsSsJzBZ47HuB3fN4Y/CLFJcebGhwwd3bkHrb8+EeLsgmRgG00E2o
weJN7USixNsnl9WBMZ9CARZKciWMgKANDYcTSd3Oiux9teNNe7Kvp0rtA2X9V08I
7P8MVD51YCRoIUXsXn1rn1OUsliLklGw9gpwdQ8/Z6GOT6nVO/lgIBTpfGcvCts3
/rulLMPY6Q96MjWS9BBXe2o/5K23E1plX33A6lfwtA3fMLSTOCuajqmQhizuSZ7O
sFaDMFqwvj8XLSLLusztKpROPTRdZ8tKJk+UdhTP6sSCpxsQFLP7Er+4DUt42h9U
eHSiR5r9Z5/DwV9m/NM/ev9n+EO/wVfhsAgNMrLqVLCndBaEA2I3ckTD0Cu/EoYz
OqkShSKfy6m6BHGThXWyTOWcFSoXK5nDq2dC+9XwQ2M=
`protect END_PROTECTED
