`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VpXPSswntbxWjHzgkKgqKOmCLgbyQwU+uzkMHzeSpvFMHmcK6FnWqQrh/EZI7BXW
lyCihBPQabbZvz9JudYQh/McBNfMlIpnz7FCpFY8mdFALZEerrEINmdZXGkaCejM
6cfiaD9Fmy4rdMhkKzLI2jlT9gp/kUeXpwJjtmS+xHdRu0i1sH3FP66IWuW68xTj
Ud7upnUniwOXF97DXqzY9K3zXNh0j4zzwYepheTfy83ej2GyO3U0OMM96LyZ1r4g
Ltig41tjilJ8CpJewE9N4TVxXlG8z0Q+eTlEFQE/UiOYB9pEnnS/UE4ROOh5vul3
PzJEQxIuFk0d6WDi6jN24cYLYPd1/3Nxll1JHVXSX7o3cgVmHcEUVxbpm5htF9S+
u11CkmAHMgvWQAZPfjshsA==
`protect END_PROTECTED
