`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sXqJUqu0FRINlucc6OFfgSgBBC4Emc9eDHbdVE5pnCUbjbLZ13bf8qatjAwsdPm1
AkthqMkiAoqCkJvc3Oo8T2ELe/x7q1Liky7ug7lCEQfp9Hmyy7pkmFcptFJJ4tdP
GXxg2w9flNwq4NJiJyB8d86BZYP181bFUMnFzULdfVfZC6SRw6VPMj7cNjTFwNJS
SsPE8G4Pi9x0Ej9ghHwYqSmoZ9cD3p931JSzSkO4R3qi9SGeDnR5hfchWMVVh+ge
Tl85JATarEXwIfos3yIIuoc1bQDuqbC6Gx+mbIw5XqhsI2PO0PJ+gVx8C9IED+CQ
+TrYMjU2S3v9tCZRwjhY76NTVUmmPFnkH2a15athMiNMynhQmXXf69TX1J+oMa/V
q99kwdy9J94OgvS3Jrlk3avXknYYwIWcylS2kiKX3pOdep1KPIK/HviU+cNFNfc9
`protect END_PROTECTED
