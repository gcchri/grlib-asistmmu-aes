`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+nWMwv/ggZNEM8anmeIZExoiQ6vrEZ/2teO1wansofnGNAkJd/ly7Z2yItMiW58R
5dXVckysU88JZYItp8naYe6hLLKNnZqA4gheAdJwHkR38yXbNbAEfsGTaym05SqL
mQYpvqmWkvtKYjWnaAtWFQkMaVJD5VYSFHcHOmWLrBwhoweSVbCBaQMT4Rwm8ZSr
4CZSQiBMyLpRII/0quegSU43ekbv8G3f2ClH6M9kA0v78Jy2puWf093DKHFVSBrN
efbK6xyE6PtRZ/GNYDQL2LyZoX7ZhSgcfMtkXA9c5IUFfdyRAOsemSaapJcXJBFW
t89d7ZoH1o3oJqF6yxB3JIsK9rb0CX3SuIUqyi7J4Hp6OKNFeieahmUXBSRVuFBp
6LRJ2RnYi8HFvRzeq2L+eMpgYnh+dVxgjJP79x8wSig=
`protect END_PROTECTED
