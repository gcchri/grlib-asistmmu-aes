`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i04u+MlgGSYKHbDfPmU1u9Mr2HdOPUMoZAiE7rJy8hqu4SuB9qO6S4fNkjvu95am
Pg4BOo7tv1iVrYysNYxHwapx/gvb6liRF9WLBvjC8LapCw1hfoArO3o0ValkZ9vb
uoj7ZYXwLYwbFsP8iJFjlUTBpyoL24oq/i6pEHgY8RYJvCksjCHtv6b84thYBZo0
eotkMAgRxQWVq2WkkzAN7VYev8/4m3xUzA/8v2u0Tv+VDHgV/J9rfc3Zmu9pkkxD
W8S6gArgvD3SLOAncSb5+FNckuZH8V4Q2qfUEgAQeShzmGHNmSreBbD2kSGvf7pL
i28wO94T0OL+mr/7wZRuiUfFGIROwtY1idJaxt4rf94sJmxUrc2jGh24KipLBJHO
95FlyJYkl/FbLyr736uARA==
`protect END_PROTECTED
