`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FfmFb2c903LjEHRJWeggJgaoFBxnxOP9Xb5duVZfXkCkc/vl5GpT8zQp2/8Tsy8F
cM8rrrJ45NPi7ffZ1SbAr4UDwYEvXE6A8UcFRVUZ4st3MzZCNbbXbcxM8d1GJW5B
l3WKuJxuBlTr7C9YuyL4H6s4S40tNE+5FxI+7KdB2akg+Gj5SNT6OHAothb+tCOy
6SLkVeb5NaM2Xc2a5nWKuAbVDKkBZlKppklZjUizIIBpQDuYb3ictck//jbyyihg
DcMx7X/560SyNqFYf1sIx66iAA9DFivWzjpCuQMEXiwAdt0yPn1/SfiTS6m/w12z
u+P3jrKmTvsFaz9Jk4AMAGALEdLXGpKFrf39fr0FS49Cp38qKq2itcXr6OWiyGmU
4/xy98PcZRNZQYNmJ2pDjTZ7jm9sYCAMFxmw2hS6wBpATi8o0JJb+1nVbtgp1/O6
jiJ9pL0I8da8Vn+CKbKoX0TkzQ65KV30ovJYbRHq8TaOarsokg24KX4F3unCRb2W
gCUKpErs0jZr6rnGbN47PHOnd412HhqvpPcFN3LfHGcxorSo9ADo2NCOYYIOD1kD
yCtDTkeBBPJuYIWH0mebCWfqBaO9ZF5rqnAaGjYFHLOc70NP7DMD/LERq9MSuUfp
lVtL/ewkX/X2+ytMwzmma8OX27U4lR7CyBVBjRLSoTG4lH1VJtTC1oj2uIoAr+bU
3l2krOlkVDIowBaQa+QU2jmJYAObqLHlObreHt/1ZA0WReLgvdaYLIpvpvP2gyQJ
BX6ISUprV7lLJZCqiqPDr1hMo/sm4Aqo6r2Dv8AuEpDjzjMdpkNaiFzn5WjiGLf+
Sqg5oCMB67V+eO3kI2P9hio2ihCQHBWGPWCgpWDVkMta3Y3uz8cwuSunzJIZHf+j
FwW3fjiVvgnl++gYWu2RZvJBMBEI5Q9OS1/oe5tBXOjZFzna9uRonJidfhsO6ALk
B6mwlggC+ntG9k2/9YreaWIRyjMPf/B/Z0wb5l5Ku55DuaSamkGbI8DEiEHmn0OX
fFmt+XyF7M265h63Nuu1gqyZOTXN5tbEKELmEWzI8mf87xtFv33tUPays8bY01x0
+fcaUqK78PF/hz9tB/BiOFleZERYyIi+622udndnR9N2xEdt4NjWUttQG0qZVSCo
Y3Nzb5mexnHSvx4EhI7EGJnAqXgTysWNPAr15VqksubG85GaIWQr1BWnS+pR4aph
OlPvMWLsFiUqssUtWFXpl/Pl2Cxk+GPgluH4MM1j6Om5nbo3LBPISOgPAwGiiMki
0mHY1C4olN2BMGaSk+zCYtA8vgEKt4wkZJ9f0IdgqY04V6jSdXd0BVNPeYyqJQJD
hKaWx14r2cxGvZlkCexU7r1zMrzO6ydcBxXsJlE9C3Ss0oLL4EklTNOxKuh041ql
JLD7vljt+URiVz7pKoXLyHaSLUY2vBwmSzQSil/YWvcDaNvK+bieOnzz6Kfkv52I
PmZq6Jhhv8ZqNT3bkBp24XD4HPzb+pJBHMwQOiLhCVZIMMn4bxnqc1tL1snfybhx
HqMk5x7r307ShVamWTQp9jKYJXI/51cYOtxky6xU1roVL4QFi54yZVcVFuUMtN6F
Fgt74QxkkGRCPm2jkDLI1rDlcUUQiQ1q7px99nZgz7QjJmk5yW0J7a3S2hWA+eJC
6ecyrLSDFS8ziZuCxa8XA5GPVSiiyfrLeI95EAtEOs8LrfXre0CEG8NR4WAE9TVD
vjdy3+WB5BmW6HmgGOJKee73GxS5/vTdi4z6bPmeukd0+pIe288SI99cem50DOzY
LmiwKIaNNzcDkYGhP/jnSYOHOUM/L7kPt/OS8JWJlQxqa7csWGcBy9IF6RRhYhnL
EQZ98CsrYyN+BHjf6gwvkSsMJ6s9xLFTbTWLl65A/3O0sKRKJTrLTbeBHvPXThl3
`protect END_PROTECTED
