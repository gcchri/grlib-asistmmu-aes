`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w0LCtpVT7mNson3CdAkMQQfObuqcRuWQXJloXJUM5VWW3eKU8z2IaMri1aZhZfFR
cxouqQs1GbXAA93MINP9oIYDqw1hNe/Kk/wUI/IJdJce4Ci9c/TrOaa8WHjrANrv
ddxHlEtV2PIvpZXqiYKMHaUMsSH3npVT9myQGWo4is1n4cl0lskgI/tfK9yBfY3Z
aaD7wS2kRGcf1kvMofFaZsFkcQV7hA6OufyGuHFB0YnV1n3c2YY1jpMqJQy6AITc
eD4zEHsXFudl08pTDEK2uid3L2h3Yredb+M+NoswwuenEllAACPEowgZ3m2rN+yv
PVdtVDWZF81I4pIG6KvV5w==
`protect END_PROTECTED
