`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EK2vTAGtqAN2gU26U2C/VlYBoUL0huKteOEN94w5HPDLxw1/UkDVRqEB9xFh7XDh
utJkejHHk4ovwjKYWAnxtxJ47eYQcKn/pL1fJ2eKdtjpCVFe88RwY5rtNi2ne8l9
iNeUHYlafXpTZi0NAaAJbdXZwPag7q2IEJVxXWOnKdXyaOkI/dcW6iEDRi1mobna
C8bTfJwYiGmnINZDzsE6lmt+p5rw5ixR3qa//lyylPh2iBBEbf0X0D69FCfOUGKo
6PHFHTnI6+EmSFdJlvmoJ3Rfu/pEOZYBW97FPr3HCvSGmnbsRkL7XasQILFJB/kb
eOqeJnQbUubfkkuUWywToyO2H3frdwIELlfmvYVpyBIGh69AWXFGY98ze3cJi7wP
9Dta7u6rubZWoMp+uzpvQ78H+JL6vZIexzz39jFeEDKPS8N/FWmdu25fwqKiWkCk
`protect END_PROTECTED
