`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qnDsoQ4/iehVtzARcuSCr+Ohv82ovLAaA4yOL6OBAfKe4b8uqudpUGKLRuvlXhS+
luFH2fFae3wFZn7RYiqD1/E0iW9CIDnKIm5NbXrm2rOwJuasBB3PBnOiGLwogxxn
UUpns7t+lLmGzWlduZvstHZjFeJV7/tThyFnsFTGm7O+WUGe+b0sWe/xm/46HxuB
v4yL+MuPUd13E2GBxhq1roUUDXsKZ1gzVf4lkvvMRiNQGurj0XlBYUZnWWQbxo5w
+GJRliweYxqu55+ADWN5Sum5aP2fkwBocyHx3VvL76hgjDfyYa89A5YLdMrgmubD
dbA9SeaxlqlF4ui6Ee4X1CL2nMCP7ZrbROLRFlbiS5qobbikMi/G9Ll0iHnOMIMt
0CPRppxhNMO7AuyALd4P7TVn7izMWPl/pz41DcWbshCNK3JikT42KHZyv2fe1FnR
C4BXqZi9AyIXiKtHoBWRbkVTpEUEB+GEuSNzku/xZPGyuJJUK6GvxGDJtCsEahiT
snYOxynGnmkXfSRvedQgXgCu4iKUriRBOe5Fw+5hw5wfeAO6SE3kqtYhrk/zp5X/
3tbZVxFBsVJLfflnt5nav3EBoOgZd70CFNRT5F4ueKX7QzNd1A5uzmcpY0b4CWiR
UeaWKaOe5jvGScSzgfuLvYNkL8O8B48GoHujfP51FSofMSaTg4h4RYJgO5ue8tcq
QUZ1Wu0qCaaYBMVUb3QM8zTgWVueLjJjoWZ+YdtjTgyFbIDwqIBuJBhyn4AogLZ2
VCwP8QQHydItbXx6m4ypA7PdclqDoZkl7zs8E9xECpGF9+vMNcYDq3Fy98atPsf+
1itsMZcx+i3nhHwrtKqgVl1leZWkAQT2p54E98vFIdyQx+i2t7Qkt3kziBCSbwvs
3iu1nQ63ByO7wSQWHo8zeqocERg0QRFmghsdlG5S3DmM50SnlabLdkyjGHVSwgfC
NFoHgnrFrGJXEOsewzCS3bK4faWGbdRsZJVbS8+M0wftOeT3fhz8fVI6Y0crwf98
FNtgUuPA+e6AgDCs9M0unPAJ2iKsdx5GgXaAdsaoZhW3eaYRkX/3ct++mdjpydtE
uvK81/Mg/hxyzMT25qVnlkrcvSzazAOKKnY0Eywmig4rNMYrgxQ/tOsixylB/MSf
hGLiBbH1z6/GNE8K6hoDvHOakUY7jGRuQKvh/b9eHjGNs+k5uXuCfga4s4QxyAtr
qDSUPVspeXRVchYFo/9TMJlXpriUM/zLOB1MVwO3qaGrllF27PITgji/RqScrNc2
a4UtukCIgw+AxMoKd2he6nE5PPu1F3BYbycrA/dxjpC8PNGHhuJUNBYCu81M91kg
nrzW3GQ0JNeXuo+5LncHGIhoGR/BHXZqch+slEZKYv6h3hDHg/pCSiymqVSy3I/J
Ppctb300suasJFWI/UONcSwsSqauRn9QZSRsc7Skay2Qwt0dWz7/MNKpOP+mAaRe
vIAMA7El+RMFxcZ+5RBa/slE84EjIaRUh23O/5+Dbfzj+UtpHP4ww5E4xzQc8+2e
Yr+c/gjl4vdjmP/r+mnUq5u14KlaOt8e7sakY4gcbacLqtigK7O4wKspyrVpbt4J
GEhMeR3wQYE/zBItWzFqdj0ug9whGoUZJbTYZaqU4w96m6MlBuj3yqUYkLvXJVmv
x9JPNe04DQFRZnwxgEWAeDBK9uGOPD8EPProQug8Z+iRFpeoSRGzeDjgLz6vZwkk
6aOcDliJmjiziUwKR8VSj+WaRBd7bBKzlf/4B5qirY/2rbmJBHkuntp0p7nlwxSe
iEXACl5qZff4N6FtLWOrLw9/ZQvHmVT+VrnUQvP5VeSSUZr9Rzcf+ZCbFHZo0ckb
yp6q74vsb8syVzwbUERWtBdaHphXEIB1eJLU5qNI/IWbzTgWFXdNzShyxJgzDCd7
anFP6O567VbESuwDZvxvYX0nrdkB+HtPDoNsqkh3n1Nmh8dtapdltDzxOO2l8XHn
NxbHg3ZbM7Tjx254msngWf8lvaIMd9zpm+e0qcE1hpEfFUsyLF+ZQHcYST754nGC
b3v3kvr53PFqhAGm13ZXglWqSG24NHWTezR2b+d+/3B0rDMwWgSBBBF/iofx+hlO
4pN4WIe+DmGTkET10wzMcNTIseGDWPYi7OJDiuG3V9ekgIBVCppL6eyq69fTpmrN
RM/3Q7tEI5ANXwcEiDv7a7gU3PXo/eNVF58bDbZtOHz8af7juMRHJTXPMXMdFjt1
u5qawMDWVicLpXWPcmj9X5qZVDgvOhgghzQVMmujeae06EV+VZaJIxJeSBVA10dp
HbSv3OwQU0qFwWfmj7ghmFXUt7lpdRxkC7ULLgbuiCPIISk1hXO7xLLtaGUfv0sz
ew8Q9cXZaswvP/TP6QXMbhLPfGwAJURMqXOovTN31c0=
`protect END_PROTECTED
