`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u7QVPNriy/wC+9EO9hYBAMtMwMQduend11UquQdGpcpWpQPoPNOLh/g/qCbBx6C5
Qcg+mwarOkHjfLtrCZxEGkSk428ekAXr8p9h0S0sS5YozcUGQ9fsaPBC0JaZUHIp
nwc1LSYoIaq+ETMpsbYlzxWJWnAXC7OQlM6KoirMUOVC189duJiXTQSZgTQA+0q4
I+mnqTc62eMrSvm+nb3bTvf0ddLW6xTHfowpfWEnoz/t04nyicBxdpgePBKctcf/
evya4DCZuiQ5/LalKmTneA==
`protect END_PROTECTED
