`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
99t5lkiXSmBLtejYBDtjyppGbiyRbWQRcz6JogTLu7ru7Aj+Q0pOwQKJh5fIvDp8
6gSg2jQUVoKMyHHXz4t1eea/AsuZHecvL7hFVsPlw4GtUosMNTfQsaryCnlsxE9G
gXXCKLcmym9IK/8WZuZ/tNkZhVxSfboJdpxFAAbVAIL+Yd60AiNlBptKyXFAlVKj
PHWBV8lAOlqlU+fWOnLW+/HK/HX5uN/EIkKKkT5M2Cpy/hY3YfPTsUHfHEndweWg
QaOZ62AWmxB76vxFi24Muk9d5r2hMpU+x+/rLunfBAGa9X5KPfuPFUE1RXV093ql
QPwHr5y2kpT55lb3PgEg9P6fEz2mgccfXrAJKwUGs5cOZCAIjLN5Y9lT0XXwWfJT
79IIVxdLCp0Ifji1MYpL/ih8/mrV+jdjTBqmfzzAnwc1/EWyDxhmj7PbWTQZrVNK
NOiN82j3bqJLzFecfD6hZv8g8JczxzgzZ6oa77orOlAP2U51R1l6nYAAZhuOchpT
oKm6gpiwDw+kms0as6SRQImV6eIqeJd/hAjhq2keaABK7ARUEn1aUTl1qlzrBctI
R0E4Y8tbSYqAt82shP47MrUCsqn+Em8G1aH8uYMu5ubIHJMO27ivbLI4WsO5wX+z
Sb5XFySIJEhGVzftMazBAWEZh9SAANprCPgegja04RuhBYIWoxYTJMPHYaNe3dTY
pXE6nU3NGCHfpRPXLYmIydYuOFPvApfawDVRugV86DZWFddLWFJM9Css0EmmpEm5
8uf3u2BkDOExhVtNTXv2/JrXCZ/DHzWVuLFGHofp3KQppWPHt/HufzUP5pgvWZBe
Fpi9zaAmw8xj/s98391wVZ+wcxyB50TkeQaU3aIKIoUmHJlu5GtFxslkAN5/XYOF
ZU+qhFv6EkwHWi/49zuW/p/qu1EvBGc5I3YBH71sJIqDW26owKTV0dfPcqsqzEYn
T+KH2c+FU6thFxQcnupfM1yh9mvjx29/pJV83Y3/WTIAudUXDZ0GTHSM5IqE4eo3
5oJ+AsxsjievbLW/7Sys8ssW0U1UBS/bjF9qS70XVOckYJIBRgBshcqP8390OeeC
Y19UpuRejy3sP6NqCbvfH4/kgI/no0YoHW6Xrj9msJhcOx62S0QW8RR/VUIC1M6H
GcSG5/ZdOx6N4G9iU2iZ/+dtHfSRyigB40UYquAaZ7Zb2S94W9IRv+gWnDUPwfFt
8jHKV0964Ryh7i94/UTcuHFrXEVuiYFI5R4VF5n0amcTgHJ0K6AzYCIVHQftcaur
2hAgT140MheFMzvO9rVOQYba/oTYWsT51a8mV0S2HaxhumPXXxW0TVGWh3CNj3I7
hGlL02Ouwdq1nryYS7ERG1qzZ620Nd3SrIKZVG7OBp8HtCpbVZQyyLloYLrZBeWy
i5aiIlhdbF88ujcWjLu34ywNsBb70UEmvk7sDdf2+f1CqJzxD43p1Zmxn2nwzT6p
ERKK7pzKL0dRQixUXjFpy/e49nokkYGGNkkoEgRYiKPpTEWHzcCImabTIPC6nDAQ
/8pTw6vXx/8gBGme5/mGUVg1Oc77AhbmDv3FKYUobDcjHR5/Ttm2vPpS+NzQKRbg
qqJzA4XKCtaUaosFWVOZOQ/zkjbbbG9/Svjkx2LfQQHRhPrEqzNyhS8kXuFfnBVI
Z33uVNLBfrZ/KlhAcrftppCJF1HjOMPZLCN7dHBJdUvBFhjbaTnhDMs7aE2fewNS
Pxps1mxQdhHzYLrtsdBja3GrcDmkS7vuMgGXD41KiMkIrgI6Ny/9qHQ55hklE5jN
Y5WIAWDtGgkSjBR2b3APclvxzlmGohtrJem0VQg0rcq3o4ZhpEvb117m4JEafcMC
xoUItFKo0WZKx8RcRwTrB577YwOgRLwkKZRXqllTybCNx7K5bNBEvWIrpPCeXrLM
4flwJAEXESIP63114nLh8sksn8BBKkoGIVgq477QMJFup+fi7gBBCOkuxLp9xw71
lhH2gXJaEzZqUqqdTN+Xk/qpNRYqaszxMk8wKIKhhR6TCqVuCSLXdO6dioIuZ6cv
Equ+OnvBu1xO0fK1mt3M7NkFxtlL0gAwMowhP9TfOzkhVEV2udD1QBiPJLoHvfyM
iZ82SXGLX/8giLJzglSJNPkTFLQisM5xmtl8BjQivxpQEk7oJRLvRYW8BK7WTVnF
0zMB7wP6iHQgGIvrujaexHgtQkWH+OnbaHAeEKAl77ahm97fnF7dd3gd2vR3XBMu
P4JdCRIP0+9N/fjgo2/shSj4PCHuTS5O99YRfTMJrBoqbZSyQgoc6AVfle/+nxlO
pUQA8zdA8I+JGRrWx7QdGcKgJgl3N43xaUVlLHpjVOwZd+xfJWBMoGB8Fkh85Mm9
W9yJByHrpNJWFr4wRncnYaPIpntDV9D5L0JyNtZNgUZQKN3G74bZh0bmbSGMBpJq
pGWCpVa31z2u3P1HKxMyuttuQFpYeZwWgjt8dVTGSVge4NBihq+Xc1i3c5CbqM86
07tYgMHa2x+7lYXanwhf1HPCtpNLue9Teu5kE+kpEPi0S5VcOHnKolqkfJcqy7aU
0ezYvkMiLaHqOa9VzrUm8Vd1nTd+oDgW6DAyOuybLtlW1AwT8+a2jSLXNPEx2+Lh
H8u6LZaGa1G44+Rt1wzT9y4xtqjvMf8dBn4CUHHf1+KKe28tFCcR2OXC1hJhRX8t
yZkLVmcbqvUJUrWEsmOZyWdotpuN7by5dK5gWylsGAvDvSpLb8bYPdukbI6BYOnN
6WpJEqQHAz/5nldP0Nv8Ffg+rXc5imbwW+zIVd42gLImlpqujoPL7cTSoUg/Gexh
wE8VZIxTqdW8Um/lN0bAZT1ARD/SUSqSOUtyrQU3zE2oE6db6ylYs/jMQvCH2iwj
k5qrxSufeW4n9L27jnDKk1oboUMFGV+zJrYUApSJEcK+JqY6Kyi0C2+JZ+O+wb6+
gzmqQJ6HFBM1OjkcR8fYH1iBPrGNcpKejaAKsHmtBOtLd7+xls4U9CKUpxZ+hLAC
vl5qFfEx1JEe41ZGFYYKcTRZO3R/r/X41WHUoCBSiu+AJ9bz9d7i6fTjMaNJWeyc
EtbWEzCDOTeiy1ZRDDBdR2SxauBLpeJfvBufHrGLwUugMCpSqWyhm/s7vH+ONQ4T
oujlj9e1hz6bv8WUCR7jFAAjq0NTs93Qi8Zt12e0uARKi6z7JbKQTwEltQKCQla7
szpYAlF5M1pWNBU9TGoDkPn1PgpfPTr/VgZpGnsdPrCo55dbGFDW24g071NzPQNI
fjbtzIGg6pPaKRYxqTSsUPMmJSQOMgpPIsxB4ShXj7qovJ/4SNFdCRHtE2mieAVH
18vRIcN+P9J1EGAUxn38EC1zYDF5Taq2baT8gafK+jXEMITOiqTiDOaNuliWej9I
d04vQ4te8ykO3QDF2ezW0L+oJE1D2fAR121F+ZiWl6Q0oaKDdvJyA0W92TsT9uHb
Uj2lbTJM4RMIHX3KXaHYYCzDJhGl1cRqs41MLrxCJorYGCAJFdB7Byk3gby1jWK1
vfvttatigsg9MB8jQ75it6N5akv8azAjvUXoUNML+jHFiIYob9smFT6lwlx0X8mR
cmDDI/TNsMmcZJkanWHTUhzk3h2HQt4+DjRiWWbRZOTim9OP3cR8XuWNNLC7rM3N
EnTgNtTOs6MAPbTcUN2q+yVhvLPVMwOUjqgMXrr+8iofZ3eOLceigv7GlJiseD6Y
hY3t5fPZ/OJS97iYKCe91OG7+fXloJV1wLp64ApiuRD+MpEc5epcJue958T3lKL5
2suOW35beR/P+1+/mhA7c9Vp+AyWf1+2V1kl0/cihNg0A3IOsCL20km3y6IimZM1
Z6ovGXHVTrX4WzA0pOUmBoE7XNalvoFZEb9MWr/iHHnk2P4k+6qgD5x8uaFlPr4N
viMcf+X2RiMcrf/Jv2l645McrO/ZqJmKmexdlYi7L13q8xylRuqfus0l8DkRJHqB
urS+5JtfXShWmivN2sec5gg60KWRPkDpyxbO3P2hjHAVm5lF2aDpQoG5NPyyfOw4
9fok/9a1sOuFJqvvQ5HYGxNc39P4hrxhrZKgH8MuQFGz8Q0ktXcGtsM0y2X7sm3k
6eUbNdISmoUXPiQ5hyytbPQ3PzTmM1WOaooHi/Lu+5V1wYL2Tw3vgKFW0nGZZjQX
3k0CVX37GXD1pFPfWTVg7r3lv1IbICfhysbOOwvog2tWhtOJAojXUl8Om9xhDNi0
zbMT8tlDcSuclPj2tjAAEcZ2lstsAGk5JTt/bj7v+o/BC1BjRitZyCMAGuQMyQWO
um2a7ezNcgTEA/OrtB9r0AhQVC0O+E1+djdJNj09KpJ7cPmUj6J34LXEehazwwjb
2CTw4RLTGQ59ORRSmqb9tp4eJ+goSSMpgLK0HRUJ9Ms0+XmYX6xjuW4j3dU1KczD
kyreiObmzcCZXWwlVgiPBap55/hvESl/3Rf1/yWNBRsk26asMn80rBOV/gJZGVic
z5MlXLDIJm/y/IIqKX00m/TaBxzbOTv4ywmEX9AH7swju7IeO8G7yx2987QNJqQu
wwxuk1djZb4hyfHSpfsSVFuc4oII/d4TY91ndyOp2Eiokm8hH65rkDMgiqfLf/lm
CCNVWqVOALH4OubDHYBhqb9vLC9iyae/8X1RZX1KBEGZ7nYD2jYh1mdSjwG+vyIr
7y7JM70KmapVQi7LZxIzQEkHwdJFGpY6FDJcoVsxo7qe3I0FW+8nblIfRAofPBw/
q2r9uLwXGBc7bvvmHEIEqYdsJPNt9ZF+8CmTs/tk+AOpD6UIY2ON4C7VEHYvpqgz
nwlvCt+hXmSVDrAy+dl+7mpHoqOUtoSIyRmPhHn2CooYlKY0ROJMb7uju6hUoT8V
ASFx2F9B6u9lck1bCIK6/9MTE9drDvD2mgYIc0PH2mGpicZFqHjBbvTd4S4xHicX
TRiGc2NmNVxoQmCiPsMXDVs17/SSNAnaZ500gHevlSNKYrXBrmBPd63rKEKfFRnf
VWu30r4nH82HXvRu+ijz8lEYc8xZq5+jAIQzpP0yEcRjh2+C78wRjjSfn8GXzah1
jOIRIdIYqlx+GjUAOjpdFZNNewEw2UysaugAR3N9PCNMG1eFlp/1yhARgBUH6aib
2NfePA4XCZnZY10bJwAWpoikwfhDmJiPvlO9ZYddcVdSq865S5imNA+gWYEXDDNw
O/sft0Ffrbc9IccVZ3WPc0PLEbQorHPieQzusSRiwV16Q1uIjDUJvmZT6ARZzHI8
JNUhT9qBLyHS8S0PHka0PxQweqJsjwKcU1dmjcvSvWG2gkU4x03gLxxGOjSDN+8F
sxGDFlFdtQjOFRemRsQW6rv/hHKqXtRFpOZ9l5LHyy0XjovnnjAjZdwyqzYCDzpq
jAQsZ+ZHtvf7IZIxX7BJrYdSahGE9P0fZQok/Armh5SbTHS/Eucer8LBZ7XJXUzw
b5ayX2sXM+z150g50/OyFNfGl3qzlLmllJaV3QQsDvMuxhUq+ao41ZLV1PT9TRc7
TZOrf6Sb1MBb8PZu14VPv0omlIdLt+UR5m20j10RT22OnQBs8QUanYAcYIOdEpSA
zaahCpQcjkC+IaTN4MaZLiJOAHeUHt0pMGUUTLyYTRuq1N0cgkVT/iF1yVX/sEdF
6Hdm8tVQwNG2bzNEnl0LRu5jt0TzNHYMZxcfmHBntxFYD35R98+J5JHJWI443ZZ0
/asgh0jltCAbO+dwZkW7uK3OcRI9WRRy/wDy8Kzp/2jv7Ilv8xPIczRnqZpBmvFa
t3BuDNxaJzvDVs7i6n+EWHsJ5qR+AzKYtyuJPkvcPJ3pmSF4rQqsOFc7aUO2BEWq
3UiLeESGfFTzrDThURT3bw0d0GOLf8TXNrdkdvyibMf8wJQOgZXzPx/RRag4Da+s
4w43xbt8Y1BCiaIoRR0Ahs40S5A9vd4v2a21kR39cmFSNvziOSv5c2Fq8Wn5YzgF
1+3DgEcR0uo6Unb+/KpcnYEVlvM9ePGJhj7vAlOwamxsjg03D7ZWBypAPd4eLbSe
NpRj4zUGQd/DGbaBD0icPDZT4+aYB4nPBwYACOGKxKNYlbslC1NXsd/dwD3a8ruL
q6y4EtToG5+Ufxc4qB+MbXUM+BM+p7ikmQh1cUWZXwzp0fRXB6pzdp8rxpmn5wnw
I11jujjXNAYCvlWrKs7KB708DzEUEfHN2l3KuNmtEQbh3fVt1lPyeDo5H0LJYfKA
YB7Kh4q2Q9PmWsk9jP8nzrX/rrwce9VP/Hl+VaYnpG6cN15YRVYto8tr9xRRjLgp
01pA8m7y8W0O0AxrRuX4XAQNu11NrL5qB+6CbWT8hZb00sTCQs0k4CbHx4u3x9YD
G74AZYOqodbLcBqQ52LzHjxCbj1p9WfE/Ti57i81Z2MrdkBlrUVAvGKHUdC6GXeq
J0bW5nGnikfD7QQYaZf3P5TyByxqmKuwWdLtG4Yf8PiwvvkJQGO6onxk6koLh1CS
iwcarEVihpPihPq1m+hmfsHL9GEkI71mx+tFkyt4bX97oGw9e/YYPbKA4D/xUPv6
XGJCXCsC+FIu05qbNZR5d+YjOncYRzjEkaNGcbnYCHwAEeEnsxOX3b9D89lWYuRI
s8J/CLF6WEN9b/8VbT9vB1yyig+Sltr4Mj5KPvy3tLGVMbA/NZ5BRvR3URd2FyJz
e0ATKZJ9r5EqKJeyTzk2E21M7S51HrxS/4ivNgP/gw/c9UQO3YRJTJk8Uk5Lvl3H
tZ1aq0cfw1juZaoSLHwSvMcNrOQ9lBf+3m5f6LZ1qeukDGVBsuN5OLAFpqDwGfSV
VmcB3Ujzld0TAeKQpTg0YaX9xJquO+Kol9V7vB4WN4YkOqMDC8IbC51d7E3ebcnh
DntlmQfiDiN5fAEN7Kxl0BLwgRuJ+Fyc/llK7W5bPDGWBXtr5Z4hGMHmrc1zx1yT
7eTDMf4Oedhx562BWKAr2YgBvEz5TDFp8iSGZSF+UcZQAWQjTeyZH+FY560isPKu
ypGRHVGZrUckKP/pTn1zYaex7J3565aNTeuJTYG+pjEz2TggNTmvpCkoc/IRfyX9
f4AUI/qhovmkG3ljA4OogQKjigsGOsSX5v+/eLgo9f6qT51lea7fQUlHI6HE8KlR
CRd1MsPXUuh3oYJdcyTzenita3KhBFQcZRDDhCOWnVnIb8pAgNs/Qga480IbyOuu
zDJqWr/oDkCIWxtCuuRgy8HPtFoSiw5rHsHWst8/OgTxNdqRpkFsZBd8b3B/GzTu
IZ++rPzXdpt8kkSoZrGSC9UrKn3NR/SVPCrD0bXEKabLtM/SQlybgtonMe/Od2KE
NWOpXccK3XHbcU+2YxvyUDUqonpuQZBttcPm9m9OvCMYqlb78EjTm3a7PYcflgkD
o7kvLw6W6KAtQ27+KUZjA+huUZba9/ffgexW7s+NgHHq0Jl4Xnx1I5oqrmpoZmha
9IvKHniB0lXWplyYkY8XgZFY9j9NPuwaQFS6gj0ZlPOI2I5PRRr7Zd2nWSadzdSh
YEvybD0pPMqSkDgNqcGpHSxo8vjjuGjTmqNrp2TB8wA20EKs1KFfSjXmGdu7dlt+
nW7KZAC+oCr6t5HfJIHKg/e4sYv7LSkQuXnYYs7ZvKVYZCDEb6iiHTMOelY8v8G5
J0YZegcZbqcxsXz8NlmeyBVY1FD03TmF/0JRm8h22NWLaIKDRUaW1uaA7NfuH0Jp
a4VGFWLYxPsV+9rVs/oQ7DoLMAtF91TmMeuxh8fhXGf/Ed9brMw0MsZt1VPSd9iH
SjFrVKz6u3lc4Gyv0pcfNQwcETGshOYWclTwiv6YTSXkJFu0np19ryGL7GP/N2Rd
w/WCrtml9V2dOn9lIsztH0B9VabRu6o5/mIeOnv0xcRCIY1NFuK5tN2XPdTG2SKA
yfM6CmYFGXmvuxSc2ryyf9xJwqFRx/ZV14w48R018OkYTx/odNycdM/LYGVX2FBo
M/8cueKgG6G2YQsTbd1FUcZqVVS6A8ssyyZWuHMguupDtmlxqrBhXSdXi7xZUwFg
TW5OgpuwHBsZROU/w+mPAqzNk9tI/XLLpij3knfYdxdh1RoHWw95dQasCz5jvACA
ZyyhWA1Gap/nkY3luwqxfQiktPrvlbyTF6iyCdRWQ3AZwNyq5PV8mw82tsvzV16N
I8XYr4M2vvjAThJGs8mkbxorM1PDMeXhVELZkoMWfF0RGubpUBiSVqZvBkNhD+Xf
Slxe5xHmeRpot9ByoHSJBB80kQy0boFc+5XezNGYCp1Gfn7GGn2ySRWs2KpW7YZu
jzzNmiZQR0dX+OxNhLbnxzWl5+Zc1hXIrj339eAa+tq0knf4rx20UpBph2px7Vmt
JETiW4ity28jg3Oelc0FRKqbnDbVuyZ+lKTYQf1Ysrf9DpcPm9gI7sI5fHeL0Ahb
l6Dd+j84LX2rJkWEhCXWjydTP4H7jffIqizzsVYTX7sLmRKqZmNa84wfJX8A3olo
saDZ72+sawvqLDGrGJSoaBZyWmBvFJwgy/wshqXC7d7zS2NlPy5hw0uv/LlXpp00
Jc37bx3EUTGtgNqImt57JMbQ7hiBP8AzcflCDMaJonhEz44IDVh+hg1deYeItd13
+foViOlVHsUoDQZt53+QeNOfsZTtei85nVKBRO9waBPqdmkDyxKjOpg92ipD3Zfe
LtQD98B0/2NnWbaJt5XH3vq2RI3YZJaFMloNsOPh+SrcTTkUffbmzWOdvFN7ZfRt
+lJE+yH5D5HNkkq52tdSfDGFBUNDSN67NGH5I4Cbu8VX26jiisNbDSsdTRxa1Qv6
Odh0Yk6pTU+AUtrDo5HwiKUrlK3NM8e+SnFwmCTknURpOqIKjTCb0xpO0LrP2Fu6
JKASOOkd436xG2Dxn4VkzJ229drCuDur0x5XJGASYyrnPVepecS2WPjatynr5uc5
Ev6ZR1r65LfKLFgry76Ln140So7jZb8AyBBWPJ6xlhUGX8vrnG3eJIH/V0yFUsJw
ZU6q4bhTWNzl4+L8eH/NPypke/Y+Khx4NJ0HVv9DlqRQEg3DNzHzFRBF9b9vRGYA
oIvwLwWytf2PgxTU0zNko7qqJNNZiSb2Z4oXYqdYBfW/k00W6uXpOwfqAfc0SLrU
XsBzVYJN8ADaHojH6hKTmNFaP71UdNmqZZJ1G7cKJuHBYhMSBWJuTVe1xZgjRYpQ
h7dmy8S7MeOtcTGEjhnG6e6dEhPgwR/hW5Z59PhbVAMqctFbwXlqfKOcGhC7tz8i
cZgfCTW/wUdP5clyHhh4AN90kcU8PZBQBsBzOiSdCqhrydRy6lXFDj8B0dsdVMp/
JkTJ6ZnFk67zm28mL7pfKmFKDc+4xB5xXm6tJ/431D3J5i3sAfubsvyCpJBASPMj
6XE2pnZQdS56dSICRktKCTY5TMK0/w0Xx5lBwTGY5t6SEyx+C4aTrCuwUw8n+Iir
8X8oVbaXhaLZmnrNLFoHmUt3BlZUaWGCO/7K6Jr5xn2V/7YT6nap5EoYrmsxipWU
JRVaGhRVY0psl/vufXEQ0tM148cmaUE2dqg9Ak3Y9he2eftMjH/bCRfEZy/d5L24
QCOIZvpmA/IZI2NkSYdPqHaJL2iDcd/wiw5eY4BlvFxxvvF0o5XZv+OGSCD7Pe3K
+azmNeXWt9kUf4r/T46HI/FNmgWE9JcVNG9zpu1tjP2lTe5+lRcwNS2xKQlM8I96
XbNM8pv+3zuep5/Bz4Tc09EvhQwSF1V4tS5/5VHSGgsAzUyoSYa/J8oKIqn1ZBkZ
nRxlS0f28WbwKltamcIOoHrii/MDWhhMVhRqZdWWg+UewR7fofkIBXoVEvVVM0gO
MstuQqeyoJl3m0mv+QmIer77+b7hYvRWc/vhKqebbZMI1IhpmyHHzCLxfFiwm6lO
CgRhx1g8O9wNcRoKWATzPraw5cICeIt2eE+XD2Tg2uxK5uT+GKrLpExQ9LE1Txak
LSPM6q67d37khnc11d0/MJg0UFREs9a4mxYAkdcUJNYwn7jyfqwURXtMG/rI7Jt6
OfYFI3ayboY6dd4Yt7Q53h+Jx6T0EH52N1mPqNHSc+uz4wyw6d+/5VNbWITKO8PI
viDqs6aTa0zwfhGHCDFQ2KlwR/eTEz3oTZpoJQrQ7fZfjEvjfLt2gah+DveiLpdk
7jBp3Cn4MsYbgXlEs7OkJZ0nCF3Z70vhFZsFyvvYbsM9qN/N1yyO6RoT4fwH8ftS
nkb0V3ZeSUgRxzb7IzmRf7yBCA01qeOtzpeLdrBUobAgiYGa6VZW0H7574g6sdG9
nRnRkbC34/Hh7QiALdWdVa80vHenCpDzPpvhxMaq+XfR8a4NKl+4RdnjTRYlfNtB
/vPmlvCVor7xbjLPVEW9/G/AddEUB1EGvNFxOdegH86z8jaEfPuthpCbMoyxvag4
vGPMzkFLVKSj64j3yMXMfq+9cKoup0DRLtgQiWK7TWVMW4csllXiwpz/jHZ3zfZ1
O8IFBQKeyRN9dAP7xF0m58/8U+u1d4OImgSOK6LCBCi2rdciNEWODXG5tOLrqN8z
KuUMGCVXMAw0opRZZ86ZGTWahRqAzb5K9nThAlv6UvjmBI3pW4HKB3t8o+VVQIBX
cJ6/ofnBFDFNRkdmK/cU0xfzghvJQMnsKOr/iZChlKOtG+04dYzFN19nxdJsi+Fs
xh6FpjAlqAEvJaq/dnMfaiIrCZE0JfsoeCs+p8i0Ku0ZpKFPPH6tAPX7sQaYLtEZ
1Ju4RKC9YKKoQNiI5Tt+39lMFW4SyU9d13yDm4kUs3zKb4y/MWWRFVFPSTVgLMBs
55qtvt2fALhHd3tj8N4x5SPdUGEEhGqh6mwd7GX+bUK6Bf4duyToDTCzhGM/F7ZH
BfZ0kJaOOc4oCND+g548muok3HPlJ01WrTSLV0/VZbDlx5Av6koLhfu0Wf0TRxbI
qAJPIWJuGR7L3WmqBlBTMZxfjWEt2sbhe1X9cO+XwC7mQ0i8JtRf1lfDnVRtZ8qB
GavYxorqR/LHN06Y9qQmLlt06aCRhHuHijvsByyaQnBlxKNB6er/lDJFASpFt5Xx
N3ol/ZErv8tygl77b1mbXcSI02EItXUqqBDVxusZbO/O8DjzB/IdBHCHnOd3BDAD
mHRXLNA+wswX+FGEIrouwByWE5nzouMyFW8zJhwbHnw5oLrC/VggRAA/w22QjFy1
RqK80clQu7Lj/MoFKoRLMKb33Y48ZDT0UaaI9J+Pz5COqAco0rmrnCZDLheAiH0X
vhy4DVUqDOYuzUAWA/UtkOx2m50sQ5wCYJldrmnca6DY3lRwyJB7urlZm8piYb8e
NK0yz51b4Irm1pmafN4c5GjOl3+sYZ3oa4x3su7sbBb0wPaJiDvmUwSpVFDWo5pj
PWMIi5i3Y0ADIue2I1yMNhkq2a5O/CfC3RnO3bzZmp3BmWYuNYeuuJL0YX+gOMIV
TNHTv3+Si59FykvRmUtK/9SqfMkV6Hl+Hi9bhNFCHt8AtEpKk0gsA46Fus9NMilw
B39JlUyUahhDSKDTrTfDXfE/0kGHYAL7+2z3WqRiCvyBobMAGkt9P9dLTW2RcAmi
X//YS+n3rxue+i7Hh4wTcDdQrULArnzr5daZaNlvuXVrKIDbWcP6kc2Y6qI0r5wu
EyiQXKxLUP49LoKUDdElcD5y64LGITvgZFj5mjwTP7Ys3VRYJYpFiq8me+IeGtvd
h40OqM07PJtgbw2IW3vN3ZK+LIiYRfsf/8r34WA9Nn7Ifv8rzaThSViWYxRWeRf7
UxforpbHhwz0jP0WQfHZmXonDRBz9PMLaXkqwo+szEu3cPQghQrCU1dZIYlZt9ur
UEi/ZkmqxAl61U5RlJnqB1ucpUVEC3k9etEXfRj34FVrO8X/VRJGQrdrmZfzkOFP
8W11BicXtsTiDL3X4eG9l3F8IGcQrWVCj5pvBm8DqUehNIm6PhBAqO+6Lidb6UnZ
KftQ22Hl7+mV2MXH27/Vs341rZ6rBXf99kABUn7S0ZTqPDQZooezmdkviv2HarU4
rd0IytbLZCs/oRoYiNOHCFyJnqBV0/ToqwI0FtAzuvgDhZAjvG4O95enl46WmLJK
Gy9fn+Scs0lAi52XNsCGOSvbEJ+TYRw/0CxI97Hn8S3vEWnG/qaKsJo7lvnQqzv3
Vs+e7FcVe0jI4yCLDoo9vGUp2jYdtDJpMgL6Ip/WeivKBVG85ZebGu6nuEKKkX9j
8puuZDl4F/RC1A2h4ifU7FViMbtvSoJ5ijch9Za0C8Kqq/vGSlPTGMc9nFnP22Xd
rCSV2oFpy8qxX4tA5LcKc3+d4huwutLoQwqtIumpnmp72z0O1kuRz+PHu2OjhpFf
htHw+dL4NYh/uwlXViVsnu/eLk+vrHk7WdJYk55b+PJlWq4zzE1qgYFpdhwIdoWf
OYBxNlkMb4aGsq3aT5UIGaUOH2zSrPsDuHazFDxHja0HRf1I1AHunGL/wFFI6Dlf
3vtWUI2QDKTOWQFsJu11E0VuQzVMLIAn5BDk+orXBjcXHhJniOVMKqIaCpvrjDFW
4IvkUpVB0co1ZKv8kYbgBMm8S/ItWXCEfpLHOL98HS5DRkeObDHZCG6Z3X5FTD/U
TUif5mSNCf7GKcXWB+LFY1KOLB0ogL/LoIAfMjXa3cEOInrZkD747XbrxYVgop9D
9coYUmSEa9sW6xPjBKvB1+m0Lu3lJs5Op2TguhY/OD1rWg4vkELQ+ZcRVH8a0Is4
FU87oVOCN5zwP1knWu/kuQbVcPnS8vAVY6fliSGUZ9dxu5xabHjdV9FWZM2nd3bQ
tW9Yx/E9tjS0GPK3n1aCqkwlTgecdVQqZUeYar/TNwzZMAcGQqkPs2DopVo1TM2C
GeAX4lF8CrhNuPom3R38Mr/hGbvc8SeMWQdKG4N3Y+vUX9MR6EhxO4imzeQowk6H
rTER6P1QPe32whs081tW4dzBfaCLd00LYdxxAW0PXwHIbjujdZxFTH9EhctyLBGF
zxSlQ1pbgD9iG1aKc42VzJXK4OjmfT+35SMr55AV2C4kf7WWAFNIRlO04fOtvDKA
5eF82K/ZMAF0XyfSKTyzy9wf8ptqhzi0Vai3+4IZGW1uWBUeuzDb0lCv7WH0zxbl
/9nz4IHUkNMo3zVeI42paFZnpVJv8vi7eq4bQWa6LneCBX9tVOeij09h9FuvtnXq
Up9t+fZtWMHbTCTt0yGzpkefN7WP5J30cCmgYeHpxHinEJSSjrbT7b17qv6nyQ6A
fz9PuNQZnDwcQQlEvzJrYtGCHyNU6NgZWDfJ0FHEy+Ee0xmC0i6kUsjpi6jcekRM
r/NE30BP+sAawX4vxBe77alaxHrxoNaEGGrlYZKZS1OAezlI1w11oMvs3m8BRDw7
JcXlPyfS/2nF/T4g+7eWkJM8BDPW9qtLzfz9vn9F/3kKwP294PhFp6BCXChYUfBA
CoS20ClW2dJv1r5WrQgY5IAuQPFrtTRK1EseaeVtY3UtZbdaxGfatSSww/JlefBR
fZWaSprlhowCS+h1T/Cic1s3bA4kGj3xsCTUO4ls3oND/i0KjX1kmvVST0ljd6Dv
LlMA5DpRAOFoa8SWBsUZumWffYAjqH+WJpMzg8Ph2/Q5Td31aOIwqIiboC4WhBUF
IPo8ESfC2xjcd7GyGm3gFl359w+8E/tZIPZjCmMFJYEOevSGf+9MJkoKX9NA9E3q
GGOknU7z6dws+d/mUQGSm2drLMltkHHD79Hsj/PYNHIJQcJWJEbB4sfqqEkeA10K
Vsf2rw0MZuZMhYsxl530RXMwbuvpSyiRokw2B/8enUz5ql3E3Kp6sxFmkJrZYJB4
5NeJWA7X/pxhK/vi6K47IOB8TKtMBIySU5N8AkQlms7+56SVzMapF+FkgRdM20wH
8wfS0qo8rvMoOuk9T8GPaFpzb6M84uz6qqdwZogSJlsJYblejGXMdSEKs8Nhldmf
ONoTwyUAAw0A3BpbEEHjGqTM3ezxHYta3qa7D96t/KhCA/C3wfF/RAzAHYDMOj3V
uQNBxOf3rDCg4xy/ftyj1oo1ul0Gg6q8ab/md/MUsOrRxkIanxQSWpEFIR2jxt4J
xu1tqvvCfpie1A3XwPCS1myNqfwlr5FzQlUOyL63kkhtYwxPEShUNp55Bon6rgSP
JDFuitWSvtUIbVMJ9THdFYY3o2bY9txEDZ4adUpFMKlFyBpcCYunSt0gfLtMUyvQ
gdoUDBOYKQfLrIKiEtRs553RJfXr0g025KhoZrksvEli0wsrkjPCGxIJ0tNNQJkV
WMt37XeBXRbG6XmUj8gG93rAW6X20NbRg54L43xXBjIs7S28Y6v1PmSBP9MKYSHW
5fiNnPAbTX+aEniMDGl35PZER1ohhlQd4mJycAXOcR/uak4rzcipPGbQjpiFQSqw
cEZj9Rl8J96XQxGzJN3G+Ptn9gjuAtG75NvyViyoLur5+GBsChlnzSWr/t5VEtUb
VnlSxFF0L27/OptcLjimWdiXovVujAklMt44GgkMjkr/6VgM/r/J31fCJaSZhywC
IGCxtjSp8GOIBAyUXfrb/gWLEjMKB2ra6eqzCC5l6Z7p9YCsybWINEo5iao9YC5+
ZBl9Px/j6iBcDcZwk8yktHwRYunb9hoEthBwCqpYF4MGNfJAhPbdfo9fvdqXQXJ1
OXlJ7/Zx8UcULTYBdifHzYL8qxBFEEStBh/xetsPDtQ5yQN9FF6pi/xSgMHekgok
OckbmKfUW0iaZ/dsl4N/CZxom7Xr8Vs/f8fMZsk9RvXQHmV24vXlqySgwky3F6Ew
u8E4nJ0GgXOhvy4dqkFa3jBf2py7nr0MhunSOe1g7l+RuMjVJgBAAACMM8IpXZHb
WCY0mrB4Mu9uHQsSegOWGAdZIO6XIrXSzQr884oARs87Y5qVN6kzTfLI+SmN+Wo5
B4OuNTlP/ZboEFQUaV/UWqOW52yMOI7fU7ZxxrgLy1eEVSAK7crN62NsaRDlwDRv
8ostE9Jpq/zKLGvnFQY0KurOKMb2Ymmu1BUhj3eQn11CID0x+odEH9joseo83O/7
3TQbFEk067BwD+rwr+T1fwdBLtDvNt31ajfLXgUQ7c8NMIQwCdaEvEmUdEp1amue
EY8Lgl+lw8mR7bMK71dyA8BNWivD7hQ7UhB/Q9ESdjNlfZMZiVS3orlAU5TpCJGE
6LDt6NZw8x12xVeAmCDzcs3vbwdMC3AxuYoLvc6266i6dahIqifl7hIDqER+D5nq
gIuIzAw7mtYfIIfMTDvjms4UrnfxGNbRG2caTu/yo+AtQ6HtpYu8d1UwBbHp7JpN
ukcwUjZ2fmsuc/2lA1e3s9FhCa1EOvIYtZwAioeBt0VO0/F32mZEPt0iZn0St4X1
gtTSkwjYm9xCFh/ct7wQ6vQJBO/kNmrzQNc7776Dg8lQ8+fDtfaKpAvhj5qjYVqu
jMHw+nxjuqbwka1yHLMjXP20L1UkxZEZq3KuUtU3MyjYIvWGJNuGa1Q9P3Ir3Cyv
XQka/ib3MNId6lc/HRytm1DtgGQu9FTY8gUy2/xfGyQQ21fBU6/EGyPuuTXsEA2X
7p6ttCG3Tba1viI9CiWhyLRacRwAAtaB/o9Hf7Rnszszwnz/1lhmdcTIpztHJQuP
uuARIk51TjBCLU0XYtO9OkLfMya99IpOoCopvKfaJOgC0dhm5aQNijZNX/i+2UT0
NC3Iw4ODeNRyViwZXH9TDjq4Wbc2wuwbaS5elvwsMGM7cydQhRewvtoG3AbWGADK
m6hyxdqB0824kXn1B6dqIK+b42lGNsA6ysPx3T4iZbShHQIUPJwkLP3sqzm+hJ9X
RZHxvKUEHpEefjtEgKx57NTixyEahNl97PVKos+rQUtyDL0t2bz+2fNVRVAEHH7d
GDUYwnHKsEVnGhbeHzmMvLCvymY1zK/LxMdlLIAAISfjrYa62KoP82aQec42V5VU
Ux2+fCaCKV5vGdtetGywxQQ38zKXOn2Q+flQJKTfk+3wgov0VDbdPirVng5oWOR8
37TYLBZO2GUrFm4P7jrQNG8Qq/ytxcs49Xc/EXTKI6bHHF1hcCigNOJqTdVlc5po
foVKIYwoSYQ/zurMS+Etl5B4aB5EeL31rFJncW2YZg/fZAaFjmYNHl4K6Fl97VS9
uvcq5ZZFr8GUz2YjvZH6fOixSGUTrYHwrpsLmNyA4l+iQDnm/CvriYUIFPMo4Fry
1ZuXv21zbymVSzU3E52xeGVcoisY6Qs585cTxmCpT0YOpT8FHhokb2Qv5YMzPE3X
EN5q85sPZAcKfNUMmWSX/aX04nJ2tXnGVRPnOCoz4kGFm4z8jVmHM88cbLtTzs1G
vyCiMrN3oiB/0zqk8m031alHWsP5hHlufo0UfXNd1PEXm3c3Zlz6eiyDhIbPD8xq
PBh6lsKxuYoyZ+ervSDWZTrhoCAxDJj3SlRvyqeTPmczAzPE0/KRZfZ78+Zf4QLP
kfd+YBScV+GNQy/XuEXNYsWD9462T76IXUNXd7pa+HPm9FsZVcAzCHHW2VfGVekD
+mQ9sgh7OIG1tX0NvREyMYfMFD+rVAKrCvghiqLYjnlJ2Vq85a5IggPlqueO8hW2
CAEBKyB0i4ZmbkG0ihim9n0oQ5GxXYP4dTy8RyKWsJMk9bWbAvKkiaNvbLW0kPkR
taiXl2FMbb/eUx3PMf37PNQG/7YlcXa6838TdlXu1z+qMgtWuPnJgGsl1q+2f/hA
sUJFD8hltkfhlX8XgHQ7kpj0s5OE3wDDufngaJO3EJgCccEsvXgKF3umqACzrn5K
EIIhbfE9SmSm8aQbiRl6MdI5Jc7GnE1XJWmgwk7Vh0JZEejJnCKXWKDVu2bJHwe4
VDzslWgxyiCYDlKgMpTQMwIjpkL2yQHQN4NJ8XB6CZDk4PlAKuhnnMsUkLqi95l1
BfmAwDSNwvYiIZMu3Pct0dDzKJ+pCTnnAnYUIUD06Dx/qqCKFmhceDMsjpEfC5tv
xXWD4386Cy8JKWefqzxwwQ==
`protect END_PROTECTED
