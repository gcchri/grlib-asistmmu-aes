`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9HICJXlB4ERo8s+2q+bNZmgvNtpnOzvURuHBSIp9FwR46kwFmYFHdT4HR8cJNBaP
B0faVQ4sRta0WE8omJ/bP6KD6+pxUSIjliw6L/U0sVB9NdNldlD2qhjkWKL0v72Z
lIJCnpqOi9Zq513XyrpMD9lQ27Kjk53KhtKsOt+PkIE4iqd4a1FPEvVJf/XHGy5E
+gETCiL3JTxa0OuA8mVdSjSOq41pQdfBFFS6lyf8nOUHq3Lv6m0MM+Jxb0ug4/I3
RYdRw7ela4mQlgw6Oqe2fZflLhzn2jre2mJp/CW3BA4mYaUDStMDl1+33m6Sfgpp
GI+YHos7zHoYh/22NjUGI+Cn2NJS58qtNSV3V+3sLy/GMvxC/lirXCYBk9jv5ol7
HmIuF7Au8W0ZI/uL7tAx6ocKULTUb+c9A4MS9Pq+UIb5b+6Eaafdy9YQ/62gqduy
`protect END_PROTECTED
