`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C0r3S1bQieKu8FfKtvN8Tf+s84jQur8YVvNo6g2aiMjZNRR/pMgkE9jsO6rZdekb
8HNGBsWT0gXe0404YhOjx53QVbGkNd9GAx4cP1ZNS1QTBuGn4CX2NEA4/XI/Q+bq
cDXQokqOOvb2sDQ5FMgOWxd0DgOe3D1QV/R174sizfvlAcLnEwnLrFOFmopD9m/7
ebAXDWdVh43G1tVpJewPQjvCeRhcvdq7f/xWzRbX5wHnnD4xft2DJhxJXfDpeDSX
2t0qW6bfA04dI6hBequ6iMMFcUGvGX+NbBu1rsQDzMj4JXOHh0n6hPMLXLzwC1S/
sTSaPw6eVnp7DD7u7Pt6mzMK8O4XDXuoeLhG4a8kfkcVI8dEoSBhi7myi+Pg0k3r
D/ppW7jOS+T+ncPUQWXk0sb0Xnhn6MW+pKO2kOgQ+fg=
`protect END_PROTECTED
