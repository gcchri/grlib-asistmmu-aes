`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cuPooWqqq0/eOqzGBPfmxSqkmRcsYUWq8drswjwlUkEL06LuGiBIqPu/nymA3Mre
HToBxcOdaGLNZnBHbaP+5PT2b8bdxuEQw3ygXZPkh/3k0lWHd60UscLrjJCI+nwh
wVCooro/Gtq7T4bYPI2T7m/nMmjPYMzTvP9Z5iQkjFd3RtXo4HkxXbus0f2kiM8L
laixpMbwrCEkxbYAvtYx/lk5yiocenhMAx+KKoGLbJGVaYyiU8ZXBZCoqgbX9dkH
rtSZPF8LL+Qii5aOiFwVpRrRbXvkGS15GU7DgU/ARJ6/GvTKrqBe+VzHT78VVuD5
Igtvhf+sVqQnD+TMRF5ZEMbZUrFoywydAZBtZ2mDF3tXOB/gcSMe1EM5/eFRabfo
`protect END_PROTECTED
