`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lt7aaKBlqUeYzOvzVfASiNodaV/FBUdlNx+JHV92xQXHctt/LknEokxzei9h+XqL
9Kqwn0wjBiVGRAWL7Q9n/DAuB5TlhUtxUjGnFbFrpALyF2iYHR9Ju8uoja0I8Skm
m5xTfFZ3G++VNJRn4c+CT0NnhYWg9qN6IE8X0YOXlEWfETrTXgSFVU5aGC+TA8JC
nHs/QDwxCqBPfDLWt2nrK80kEP21arDZx+w5c1NqX1A5lJo+NJcxW1NbmTNH0QKj
wFpMbYNhqHiLWEH7MTPCFBstngbfehXk2AvHmrZXj/lGOpjrKjHE9lkwRKW5L01c
ptNNXshdg2dCQC1CAcEuvBINXU8ERHSPXZ3XvOYSYWqTaTmXd2dpgBYd8uub/x56
rMUYYiqdMkwhn4RACb5saigy8s8DgaZciVLee2EVPx2JAh2+iP3Geg1REhTHwGEL
jI45mJLfeZjp9vTG4ILB24qpkkURbcefiGjOTyWW3UY9J2omJfvu3VIDGtpvr5Da
kVas9eptporcvns/vPTIwcp/QOWeX4j67Efzo7wwfWQPz9AA10aEjLKhoriduev7
XrwGbi14XlYiT+DAkfzq+YMsNOPyZK/DxWJt/CIYSOF4IJbSFsg/GkjUo/4jIOKz
0y5KUrg8hBcrB7Sf8AjYPPgpBuiZrcWAZDWgGKqCJl54FLNAVzHxzrLG4jogQjcf
Tjx2P3+OYjxmbM+9qiW4hYCzYZGNf5xcqp6RVYkssYgVbbaUgsGX9Ag3B2ffB43r
Iz1bTILLPE/HvfEtCWkL2HkPtjhNI/izXUJo0CHIGDDumLqTrbxdJvg7Q5y9QUg2
Z+N7ZaWByKgIhJGBfumFyw==
`protect END_PROTECTED
