`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sRAQL6bmKb7QkR0mS2Eq/zyfmFDx+kLji4+9AJYt5HYXBfsBkB06IJEuwavT6mqJ
V3ERRwMIWEHZYGgRtAiHPHu6D8xMM4rMw/uZu2+M07PDr+a9DzO89Mdl5I7LBllz
m3x1W6cDNJiq3S261Rsrfarn79P12nu8tK2Gnc3p+97I6XxB8YfXgNzyoEAOefpV
WPwxJuENXystifl5L3v+rlGByF7/BFo/0tY1Gq+Cy8/326F8fVmb7Le7oAtdG2OM
vG0kddsmYhE68U3oA4vYSfzWg9MsJC8RH5kjqyJJwVddrB2IsWUn6ABBuxueGn69
i+mmJNjln9pYZEUWEZWfatYbtmbuC+rjqRFIjEOSdh3Wh+CskHhb1+t/RlJHKHX8
`protect END_PROTECTED
