`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mhzfS1nGfoZ13842+T3Qcx3/UL2KE36stV84zDv1rtFMdAnMQUOderItQcz8AbIE
IiGATLxfJzkovyqi1gulmiL5g2gzH+gyx8z/VU21XaVh12jCyANfkOaYhsi/tOxA
h9psA783hpHX88nKUTVCWn7EZkL5ofQm2lloxmTx35F9/Z/c8SM61g5T7adXxA8N
Voxa/SuWBOjVUD3wiSpkHlemhuNO0vw0yVPGzAegWfKN2vpoOELNFPNodBrDZ/7k
7DmBaVNCFrMvhYi9i8Lut/JmGENsfqP1VXimbIJfefQWzGMdTGghFhQqVLs/9AaO
C5X4dzKsHR4SOD/vjaS3IbyJBddJTSLkloYfaIEtLzbkEjBEOhi65Jrc+bxYBe1L
p/jaNVplsNfBVa40mXwWMOOwm3OIFNrEjICuV3feHYZVBBmbKUsoz8rW/QMvuAtp
PTFnw2YdNAw1ySH+fMPmaA==
`protect END_PROTECTED
