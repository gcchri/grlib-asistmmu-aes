`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WUHy/w7iRbhq5Lfh6+vaZHFzoJ5F/rJvaT6TEDJKbtP+g45QA8l+VMIVW8k24K6i
8jgEkdIkpRZQJMYELbQcDWJW9yq3Gs/pR904/px2zOlLsGVUrqVidVO2jW6s3VUO
7SvR3NuqnXwWcCGw92c3Lrm2+1nnVdaUJn78rySovwjkydiReqIA2LoYAqbf1v0N
sKpTzgsyJAXoBMtqft3B0yRZ5yOcWIKFNJ0TOoG6clo0laRXGhafQW4jIQvvVSh9
LpLl0oPnAKmtAJuLEQECM8TahJ61Qu7jhoc2PLUjuUS6L7rDvjoRHHkbPpm8oap6
Zhss9/E3AifFwrbA7B+kIlNpkNl67usSBM+yC3Tyux7wffrgIALHIUKaIZ2aUumY
QV5y0UaOKZZooyF2plyQcIpZqrWkiVg48h+vKGUap2E5OxumzKHHPD7Q2uoQfFkO
GW7DANe8OGC6bvIgHoX1E9nCLH7h2P4MfFqYEstVDaW7b5+KQJCauE221gAzzA+9
z5fhZnWRr9HXHiZyKObYkf3aSRLphO3rg2gYd2nFlLVMtMr7HZI6fXwZ0tr7IyRg
BSM2Au2AsASge7LOPuoF1Jq+NNhcqzICcbKYoT/yh5fPJhsvN+n8qIJxEPubWMFn
WNSFCg7AcsSzD3hKNb7fFWVhzhEmjOFFM+PZGuusKdCDtQSDk7K6WazNmfr1NftG
9RLcXDG0vlZjB76UkdPKOwI31hckrJdkJjZtIz61a9ZGDxKImZLQu0FapwTd/uT6
P7MGzpAKrstbbcISE1iaN6U+xGrzUfhpgbNkwNOdoyeGb0JR0LaFnK5qm9kOK5J8
2SJLh7SG5RfvAP/vgZH4dg==
`protect END_PROTECTED
