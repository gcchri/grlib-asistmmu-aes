`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qdKURgF8NwWpRHQz61yarqZinPg2ks/JVADmSVIVKPaKfecKQ/d7Io955BlUy77u
Cg6nSV87KLWLn4GtmCC1r4qkjbxmC7GQV2M4T4mB93Q4+GL2Wf6/E2U+dsgMTvXP
oKgU2KZlbu4qb3nuOaUvf82Z78ttxDeAX/g30EXfgP0fFbNKFS1fmpSn0ui+iVW1
9hX47pLukFu+9ZYC4DWQwuusJdh+F6CPp5SQt3/bIEQLtEhKSI8XZuIWsJPOPUS0
MLNkQlxv3DL97TrOaUdqnY/rCb0sYeUoYIB35YdtfIwnocodpMR/D2pTba2sSj32
XwfNeXB3JP3ApiISCdnZ/3ATkt7AKADACye1xMgWCgZ//Mm1Uw7UXPhD6FQx2nLM
LCFyKQp0Vo+XFa+GrcapnEZKYDLRv3Ks/UcCBc3ZOE3p5PAKZTD/sUhFRIT5e2hT
g5Tki0SdObvrAT+zaad416MmndTC9HHLPMHoQWmz4Wod3ai4hSYNirilzrTMx13/
7HIc0uXJt5Ip/sdqy7+93a2YHxwDUtYPBW0ra0GgWcoGmSQ0ffRKsgN6mgatg8co
PnDrphRpbToC/eEjd6/ZU3emB/RAY7LTVw9v0E7laKAxl6cDWhg/4asQl8I1dMGj
oJ3OcsPpGbBarHApfMHd+EDcXQZrkeB7EbgtPSHDF8lIoMB35lVXN3IoAy99N0FZ
FM8YpLFE1ZWrnjXslQfQ70cv3KChV1I5WjeFR6dir8hUrpER776IVwmpVredbPka
YwTRXiv+WmL5xzKsvc8dyE+y3eDjc93VHQLOaq5n3uCREDg59DhoPlJ5R7//bN9V
2nsUDQyKN/iNN+P2l87pXa/URtoIgt7En7qiTVHJEh8eYi4YRqd9HRz9iT7FbEV9
AjG0WiOZv7vIKgi+35Lf7Z80EzbyFHWzvUnp9NzWhd0SC082lHOMfe7kz00LfQPh
ZCU010Rf3p9rKuh6Y1O1P3jF7wHJ1IlWbD/VDmLnZ++/ig6UABBxtYwM/zNUDdR0
yTpSsoPJaYr5btS+AjZIe2Mwc1RSEjEoO3EUw5OFbqYTF1m69KPbmiwUDoBGOb5p
knRzstosBJTC+2d8gZAzlOnNzn2GtrRoG04MXYqqcTk=
`protect END_PROTECTED
