`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pPpX/ec3uHnPUV/vTOtOCAlIyXF5LBRhh1RKFmnnN11A79hrLa8+ngJc1H9P+IT0
QxmNd9kHJi3+EO0XM7pQWbVNERkIkrmcUWKrAN5JXPUL+C769D9XQGr1neFNgMWK
EwpZLelIod63Wezp6Dn4PubEVOFFRabh2Dh6vMM8WbhYN2Np/JGfGS5/9xtvamTk
8FrR9K5ylKb808uDAZWq75A8FF1RMrALuzulhNsF5pUJJTlVPbiEm1Zw2q4ecEMe
9zSbNgzYyBtnGjU2RE1JnOzEIc5+ocWpDBbXBQ742e2KqsytGAWofteWpXCSXert
csTyXfeIMqeOIWZ9TAswALPKOWhUTAPa6JUAa7YdL+YHXy8TBSaPSV2Zr75FkR1k
0InnM9pETPzNWpOrayV9sg==
`protect END_PROTECTED
