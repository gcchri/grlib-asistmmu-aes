`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CZg16BhVUjjSxSYDJBv3oeTMhfDVI7zAourIG0Kv5KPVDwH9k6q3kPKdvwwAGV68
PmIBS1sQ8F05X9rFz/LZkQqqIZQYXjhzCMiwLU3TkM6oWnK/BkFjRQ+ziU3aNSHJ
l74WtJ1yfsB/UH+2nhPzFBBrTZSTY1Z3hABV1oq7UwSz/CkiQmep23wTp3rsGUzm
7JphRLbvcLyAbwpahJg7RrRQnfRF/95FjGCh67xbia/fDW/IzhI/Jf9ZmcQj01lr
SJQnhROmsT01UeDZKvt2qwD1YWPVdgBqNZgwjiWIS6qoBe0MPrbx7nFdz1OT7rMd
edAOG1FnLofltF8YnjfraKWabtqxonupq0PKpXCUya0b5JOdsH9bibwBx9xSAZvO
Clq8z305MURO4iEv5uhvLvB3KN1Vb2xdRleeNRE9ZKo=
`protect END_PROTECTED
