`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GbW71ukgc3hVKKUziAIvSvm4gtQo5ieD0D9ZlWTpHbh/ez8icZIOTkuTHf9hmby1
kfQa87YumgYQi++DsHROAHswGnKmf9cjMJchKv5ZwsAuDHxmeekAWnk1Oftm6ZlG
eYDz04NI2ZfJckRTjC7GV3vBq7gri7Ej5QebLoDp5FbCQt+YlOeywcr+Sb7LP2Gu
pOIz0RGrmq7a+rCnIkkVJXWIMOL+sr1atyWJXq6DF4Oi2JWPx2hG5saiHAENDYYs
MLAf0G6J210UNxnz3e4JxLa7LcxxyvS70A2mujcsy0927oAHOx4l8M+fDfDGjv8x
bOI9AleMnc2PM3gFMsEOpWFQbZE32YkyNrYdV/xTKwwKhc0/W2W/sKiVcFNVJQvk
Po8zrDFVLj+Z9DnUGlA7ug==
`protect END_PROTECTED
