`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
88HHSiVM0owA4NtvbnurraM15Jj08jcmVOmORM3iggoMwBa0XYvhs0X2idW//hNG
ljJ0/wVXLRH/glP+eL9ohB0FSPa6vbdFrzhtWcGfA+nNesN5+7unWQqG1069bw47
ByI8daPswXqrkVf+HwhVpxnkzAIP1XvOtOj9XUPUciRxSHHDGh6x5+JYJixv3lYQ
Wn3DGi6Zc2TQIpvWd1rlINETr72WOG8/dMpIida8iiKlbHgg2O7OcdtOw8CqpoWA
8mEuI/JxhpKnpu5I8QsioaFYRFkVIf56EcW1Rx3FZc+gmAygOFMP3rgZ5lK6h65R
TNPbSQs0n+IDY/7i40vSQ4Dd8sKw1a/8t0YUreBt454e9/kM4HrExPZlvukitjft
Ae3R41x9gg4QV0wy0+TQTujU8jgpICKDHmtZCegCc+uxsikAQnAmiVvm0PbNYKOT
fXWYUzmGmfJ0ugsqV1hVXvV1Ax22ZOfVpDNOX9BN1s/LKFA8u5lBnPpRaDLGamil
zw/m4+QixLBlYEA2WWvPsIkv7z+AkKwkLELAbdocOcaB2avCEbtcDkwiOiKr3oOi
sS0loG+o38j7hAW9EhIW11Xwa/fpYRmSylZEAhX7rVOb32K793UFvUqAfEy22VIs
wSwJZkEZd8Ya5ZKQMElfVh4usj/V791SlKhU2un9KW/MqKtsv2JfFRSK44H89EfT
37p66kL08m9naYE6qVdMc4TG1elDjiDuZIS8sMiLGJ/TXr9fm41T+GxQQH83Vg/s
GKz2gdJZSqoAqs02WhDxmqepAzr2Ucl3YwaOHC5DN3EuISFZ2QLlC9f3lLUzGR/5
2HsPSVTqOB0Deuq5QNL28rO4LjnwdUQASwcV+CcSRCIn/6KWAMUZ/9QzbL+9O9sJ
DN22Oz9l69EXNsRmsddWZyGpnfSdNfAWU1GGIoPGOqAu8Vq/YJDKmc2HoHCDO0CQ
9gNYQQifnmbz7s06WlYEyXEeCmHnye6Y6LQba4siz7ryo4cJ7AucWj3igkRYMkox
OgnEeS0WuaJj72DsN/fy1Lg50aSrJ/ZzdRvX/OX+vPmv5fWp6qIDBIESjX+y7jTk
IM1oAY4DTPg2Jpn2sDfsfhVza9PDt4SBEQEs8bpudjdgBGMXFzh5h/jCbapYC8G7
988mGntQQAOSoGjyvWTVShLgU/db22FWiboi1PDHK1UGuCjOEhgB23aAqCxbtzq1
mkfMdMC2144ck3SDccanFMEz648pm0CUGIm9VjJz2hAoKeD1tZXWS157yTNyIII5
ZhkTdRTk0EKRcFUKf+kBlo+QwX06Ms2ZBifCx5Wk40aK9e4XnjsVrmPujvU4eg2R
+7uiwofhMtXXZleRaJGoKJSs3SG+nHJAnFhIhjYr5Axvo1y68zmIOe5bAJc2fyYl
XvhyTWM5+vW3eskXvTSSNLgComkgU+fgflUClAtvInVqb4+GCp08dZ+5V/VIx6fQ
JSHavGZesR5+3s5tbT/VcosJ/BGneTMeg1DzOXXuqWsPqSn3s3jLgQBTHo5RXPja
LJ5vy/vBr1ALz5H90X97sYpSTYLgcDRCec7dJnCA7UyExYlB4AOTL+TLtiX1LwOO
vUtzWkYgWVSb+Ma9x/A+6qGy1UosYBn1dlqX41ngXXODPQS/2hE4KSGxrldzyph8
DpOdoCThB9heqJwwjZc3ytj4/5W3nvXkEyZO6YluCCR8Kn/n7iBVoItVSZ8zfYkk
OTf3jXub3QCtKevgK/4aHq22HPM+pCZstVActFanSfnYJ16cjW527ubSHdBWgpbk
6XO7K0Z23GQqj5VKBbs39awdgDbSsOa5EmRyvhE0V4vOkXT9Q//pquyNZNhx5z90
RKuz+TrDZcOHpgDitbi941Y+nNB5mTwpHJk913Zw3mLXpW7vUYOQJSS0tAZ0tIXc
RDHj59pmCoVU7a0VZzodyN0+rEn1GoB7tLsZmxxlHWX8UDBoDuxINQDqfGfB5snY
X+Pt6J1pCK2lwJypcc9SR3b5U0p8vaVBYp5UZ6ukFaH2Q1b18WNj8FRxVrAInQnx
FQCzV80KVR3iXylp89O3BDlm7tAgIAYRm56TYqSQa448SPXtVWdKmZKjh4fxqDvK
pwkbooxCoVOL5rGPlMA7fKDC0h37AuhYHh9+HSZKDqTqEDHncsa4kNVYZPCRkPqL
H2X1Z2/fwMsoStTDr9Vl9drB+wSu6DTF6k49cvwakB2aCSjPq3fmvUDqKdqvaLnZ
UtNJRPXFTBVWaiUI5Q2hC720TBzajdRhs50v7AyYzaaGnl9ispDgwGjnwle2mS0g
30cShnz+CMvCuA0frd05VBa2GqLJrUXN8D+P2kmwybcCWqdK3vl8xiU5BU03tSei
DvHq8KhNG24epI3xCqHrX4xpVuESBiChQvtvpV9b3TYLXPnglZbYK+V/3zsYJzTK
YKlUPfVGDpUezBOiyNuRSCC5l/Glr9V2mDc8tz4zIls=
`protect END_PROTECTED
