`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1gMiKSRwlXQFh43FL1GagDenyATXBi1VnbeDud0AF0xQhorzEhcpz8s+iI//E38e
JkF3YdBGsCJhdp0h8JJiAtqqTiPL830+nCkIXvOYqKj8gED0396vA4ptdw+kB9IM
h6X6mUAZM7zdtWQw+XAJmSV7gPr4v16GDOuXXQYzuoLrM0fXI1d+TvLxBm2ZshSk
YQDLjUc6RfKDeqElfDVbV0T7rSll/4sVOsi3bj3D5PAgwXqzJDBn19uYndQCtoHF
ZV+CNrVIQO/4Us5IxkCIpTIhjj8qfVzA0ZCCRJhx9/CW5XlBljzoXijn5C41ghzV
NL1rG+97BWEz4C2rl15eV7R98o7awrlos6zLmGLWoWYoGnref25VN4tTYuv9SPVz
Ydz2KjYEf4sW5rlBoCxQA2FhJ7wH12FhntZ/jicV7ms=
`protect END_PROTECTED
