`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
upws1AoJ1tdcOrKs9tKKbQjwDmdfALAToaH9dOWeJmopH3y4bcHIw6f5Nx94O2/k
xvvDzo5GUM1wO2e+DEgXIqJbqGBgC8tjUwj9MIPUHgobaOktTHkWtMTefIyhPvNt
8lrNs4JdCuLHInWhYxgh7wX2z3idNgfL2V19NkOluEc1eM8piacbCOPiyLyE4EVM
VXDHFvIaLDMWnnNGtquW7+3w+Su9GRcG5THaAXoi51fV93FSTc3X8AAt2PmoW05+
J87/UxWjZqeDbwbKdE29oQ==
`protect END_PROTECTED
