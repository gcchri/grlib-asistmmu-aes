`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pdXuKdrJE3b2NX7AGBjvjWRCBpDYSJTpGUy5kL8jT3z69KE0gFnp/q4NSrsf6A0L
CvWbw5xcS3KM88QfX3/BRe6jBonTO1n2YPLKSOr0Pv1zbp6++EgdszYeesLQ9aUw
qL4co5fSACocmHW1SgsMAMZScgHWmpx9k4AlIvWEWaXo689R/lHg5iBHCN2m80vp
oPQbbcNSS8oaSf2RFOFaWcuUQSohgshC5T2UTyOmVogC8lzrBk5LVqqHX0PvYVWH
1JTA/MwzBKgZJMT01TQCLNW5vd/Nkr5CqgipmzD8Gue6JOX1Ke1ijMdd/81htAtk
kZXoLxCQQqbFVvB+HJLxbhOLoIUbV6MuMzCB35aBB5SE51f1diMSZMAV8zOhzwWN
5JHpB0yLSbNCGIzOYaqWQpXEjkJ3D4gu9EVTvp+aFMd69YG5Dc3vMiNvzGoH/YB8
mTgDf9U4ggDu4+T8ittoxfuEkJDUrN9BedBaLxWioz1nA4Lw55YLCeAp7HdNYQIz
PCk6XsXr07stGSrwcmfjwAz0VM9C7XOx7oR5nQpsbMG64fHOKWsfkAl4t6WrTDkB
BEFHW/xo0HUlZLNrSZ7d96Kg+GIamribjbAfiEvKrHBT8e+SRdz3X3YP7ppkzj+d
IWDdHbfLUlibZFFcm2C58d875rbA4UsjNqb0YqIX1iE=
`protect END_PROTECTED
