`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0yLkLp5lqg7AGg0Dd8d7pEkckxvwrDbRlpydrvTdo/mMnRcqRNkHyaQK1GblvbQu
lBqfADW4QKq3NZWozmBxecunAuJhc0ziqzWKEz0g4Zv6JdUiO0smN7rsXWQM70kk
Tr4wH181TMUgsTYokqzJqXpbyGD3dB5whmpoGAU4wHsOrLvsJkds6txm8p8OfNnQ
PJkTuae1rUPaJlt6TQUtiWMrradWnLAegYUWTRIm4hTe24/wvSuBATeTOR1wawYm
myNRYbuS00lNDJaDS4ULMDBtBudqR7gF6N7UribUVqcWcdri/XAB/A3FJE/D26Q5
Z+SKVfC70jEgQ+hM26YyQ6fhxGT17QROMyDj0i+fK9ER9uT5H1mnp0zvtWHYmSqm
xxNLzk0P+HdI0yIsEFpjj9VEBa09G+AMXxOA8ZN9/Qc/W6duVauQAauLYhNFfSER
iZS5J4K8GhxuXkloE/o2Pg==
`protect END_PROTECTED
