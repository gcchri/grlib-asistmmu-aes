`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k7a+BVFW2mZPPQfpyl4rA19/l9TVAzd3SefFJZkxyrhQXX+89PB6avrI50AJfYPf
XrBEC7OAuoX1UUd8baU3oqYEia/SwKmXnox0FpUo5LaLcaKJrtxIn0zQpZaGSheG
PfLCTwITYycmH5sgjuDkQVO5TGbRQv39s8D9/07r8FcJ3U24VNS4Di3CUU4x7B1K
YNJMxvLWy+9jalAKUvBZ2Ot4uCfnjoQsqyRNqZuuelVqmexZf8+riq5v6/4lz954
+1gW6Nqi9gKXa1GTtzRHGM4Of5y7RNZ3kuFiEpxaDmZ6orvk5NBYHFiZeFZKYQJ5
cAQNasAmFaA8zzERJUWutg==
`protect END_PROTECTED
