`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bfHttaQgvGb8LNtR3Vg+BoKpySEJvlhzFZ2s5348ZOfHJ+TJDPlkeR3KDZwHGTyH
t/vfjikvwyld/RkepcKuIuHyi2ERN+eEnbtT0eNvszarKuyyLEUDPOMJRXGtuZvO
f8ht96HO61Ot+DDXibXpMxviZIg5SQUDnVTDrCLXTwgdCqmKvVypqG8+Ai0YdmM/
hG7QV5ElEVp5nemX3IURUgA2+KqBJmUBx+4Tl26IC4gAct6cU2ENUwVWUO7t3YYR
GaL9j+S6UOX7YV/q8Q1jHJMCmvyQeQ8d8A0gux/XmKAemmNWWDb0i9R+sopYSmsu
Umo3iPTAeZsfbKwFUKUQwEfSLGnZgZp4OknHGByb9PLPN4JtMM7rLb4XBk2UkqbZ
L4jhRMejEDPG4gsbt9LF8JplP+rJimryft8K1RD7Pfe+PlKfgZkeuR+9WjjbT2z1
XtwhQ5FO01L3gfiP6GKvrQ==
`protect END_PROTECTED
