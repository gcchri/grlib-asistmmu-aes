`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TOI8J3wStWSb0+kzNZXLd7EqVXIipjBFFtm0PMsdyPubqIgLvCB+HzvB1WO6ixNQ
sWXMSeEKj3inYq3bYTjJRA5qYis8ud9DvzWVnfoxDlH1QT3Yo99q3//zGXvJcqil
TYE6JLOAqHXVlkzfAf8NgRjlfl+fKKUfXjylWAjatdYPXVvL9RagBQkAN+Y15Da5
jp7cd3f0vPd4OF/Afqdiyu/LNr5/5v3F1SkI3QloSDjIbwxVNrEgYd6htkxKwrgS
guWvUnVd+6a8rzX7GQF/x4QJC3oswDagyfrvfEcw5LvHkKfAmcdF12ufcpNyGHpw
3FDpY7PtvUqD0/du1yg5vZ3P/nHXCIAg785nanMhZVyiKYDDjUmB87PyKbysKFIT
FRej0uLuP3W1Jqs79HxnVqxKFoPEoKaT/jro5QXWUrI=
`protect END_PROTECTED
