`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qoae/OdBeSoYdMSqPaMbDgQ7mEvUoXjrsXn/HlRLyqyobRtUltqQY6wvUbvRDJ4c
pk0ZRajn77TghBPtKXVc7oVniYoYQHtEMHOTj+vttFqZ2kluafbgKlIsfa/yLTJI
NP8Mk/iruMkb+Z5hhLoitBuugD59ALCzyx24bS1MqPjGwcFEOAWMSgK4WTzOKo2W
JdryO3xBbD3vmrvM1UASVZSOgudcjvYoMr8XQZpDGX+9gMTVMGedC7XmGEYpwiXT
xtyuNBkeqWS8i+XVTynHFDz7evdOB9JFBBiADsVNqSC+1wL8ABDShy9ozCsfKRBs
uPrnO4PFzQWZkhXvvJLDf/flWCHaz2kfcbYW5Hl12k4Nu2nZONYK+28VTJF1i1AS
C0U0/qZyxNhWDceFjRRfaUD4xMM6Pn81+PS4vmP2Cjg9W1MOMtCoIjFZOKZd2oqx
9FAD9gw0PkC3KeekcChHi/AXtE4XWluoQIqhHVF40Y3W5LhSPZPpIeux/yXgH6ms
5+XX3r8cRdbvZkbezXgOOfJ3DP89qTOCpKuEdUBLQu3rtxXizENLdLrDtMLCOCOx
n8hbenqmJOA1874wBMyynycBwzOAAZB5II83Y9KVg62c/tTVYuCggwBlBTHGzdKo
aVp0Q6OUrBXqYIrNbd4/3k3rpVDw0zAenw5lX+J7/Xz2F4GSd/xsow8WEuiYs6Vd
6e/XaASnv0as3Kw+XLtYGjHqcCibS25KPFxp/n2qAtVcIZLU7hcWyH6Cg9T9P0x4
QvOOowDdRxvijZs71bHOixIK/o21ZjxvVkOVWYBxAbFGhtV3+0FUysDS2E625TLz
AkwZrrmax/6Q2ltKeWY43bJyPHHZFhREr6qD8lGnWeVYcocmsCl9B4PbAh9q13C7
Gi1aIZM6SlTxqy7I5SQZwnV8kJHD+M887/V48qy3fTbgdpALtaAGgvRZJN4Ajnau
kKV+Z+jSGEfI3YPe4r/9OjvEzfLTic2156o/pvjz2ULKtaPgjE4Bz4lZZOheF5Mb
aNb2oummzzIEuECvAgAL39RGMt85fo2OxWXHRqzT9QRanJWKERKK4sWbWU4DouCA
R5UnjeBZXAxdbpNoWtA6030x4+BCBaH7sMv/E6WyXCmQiLb0IkAIVYAKUoMAnTlN
s388sBxfj8Mv+erItoIAZ3oQOqfA1Vuz68bx9DMiig6XFambejMh8eeA8FwodEnn
aUSaqSIdbb4KWoYa8VPLGnWSm45TA0zUJjUlFsTQ8BGBkNDlIR1yrKuFauPLE6uP
jkWrFuqDssnRCIwQnyntK29VUzEPFNy+EsbQrxaA7LILKFCgC74HCsApvUhZFYCN
vBR4Ls+Wa2omt+rn8QA4tQ9wEBBYM8DqNSaJyeZtkHIz7Kg4VR80iqJKwTQD5PkL
TewoV+MmV8hfbVAJrF/Rk1xDlJebt8KJSEz+FEadkpYBE6B0z06KZ9VvYpcZ6XH7
IlqRYJ2tXRAdYMK1KQ2106OGpVSxvwEaju1DUiP4dN6jlD4TzEmhMqzpvJX1/k7f
0g+v9kzrMPVrOyA2eWBhT5TYf1c1uotw+McrecW3YLDeg71BU5yyAQvefQxzrh8e
yH5ta83NoBTzbdCBNoNs/FZdJ5gJ2yXuHaP7vkSkLiutOGqTqY6kdHFI1LMWuDfE
HsM6bbTv+MjTEWOSG4s2dh6XDUzf/crMvs98tPXpdjg0xxRxy/UQXEhUWWork3Ea
BDPYdPiiefNxq15Jb0bf+xwN9tC8Sz6vcibXhnEdTkOJLzRCD5n5JWXqxpRI8w3J
0PqdUBXlYAkfV+hD785fuWZ+sIl5UQAup08/hCUsNLHvilXbKGpcVLmdlx57xXDJ
E0q4LXIeVezkQx6dhoxidGi3ZLKzQAXTewnPghtdSr1O53gSe42hC7MZQFJmzd2/
BUXPtL9jdHDzQdbYPIoPUhQAUjTOENnCB6wyt5MDpayMH45cHF/yEWgXc4QC1F/9
Zmik78XOCMS8gZK0bde9MlPzqnUsa/X3bElYHZQWxdjy7HHnulUH5xlmbJRwXuVK
nqJfJI0IUxiEN4L3u5N4c44Ab3UxrvOvRhkiVmXL0s1+zCjnZ9oTnedzT0hEhmxi
BMdPJ1Sog2yMEWjUP7gj6KmwkvTX8gNiiJl6bTGG9IhhaMNshFBvG4gGXYgkPOHW
ow76mq4U5rWC0bkvXGURYZ2gtRXU6t+qY76NDLGeGok39GUBr7KDYAyx1aZVYuA+
XzWprWkC1BUG7iZ/0EhL9crNbLx6T0J4QS8lZFa/W8nRH69UkKonk025xA5lqvac
0myuUssolyIzAbc2AtWCoc3baTU+r0X6BfJ/Nctd6ki/aeydeplWQ8bRHXunWPXH
xsfvfkCd4sFHD9MZhCGRtj9dnKLD/TlmnytbOsKgAo8kdv5cB7akaJCCNsWvZqdH
D8OJhmzOXJ4logvkwXnOTER4hCeN1VUhyE1u032zTmL4RMVQzQ1q+LWGA98qxtiw
TvID4RYHvoXePt3S+0UPlWEm63vmuXm5QpdwT0L8mNIfl1H68FhOiqzYG0lZAari
38U0+VQExps/gFWnAoswH7+aMajrjwmEEN43G+myoMRwwOVMEtlk3NdyW9dMZSIN
CVoPaqTWOKGfn4b6sMC3F+5W1g93FbkjxCU4n4xKQhIScdNsz4MD9rmrxemHJDaW
oZPw2Vb0qR/KoBZAH9n7YuDsthhsrOIhmdtcOquFVc+j6Wj7UKs5g/kq3RK7Fwqu
AsFKysLnAT4LfdqhePeMSyUr4K6HTvicv0o1Ur7ONCsS/ae8yq6NDgxMhQyqCmZq
+tSycI8Lq49VGVtX2p1kUoHXFc1oYGV/Psfha+8A0PTMXzQo7BsD7r1qY9KpSBjw
LtS09IRg5ORr24cfgBeKsWC40zH6I0DblqrqEiCxhWI+408yvKPdIUUnx5E6P28X
7vNjda+G4TT4oeKrQY9vNdYx7QUpWxlFLYAcKzDsxzQrGVOSJriuD+LPtDlU9L4G
D5zLg1666+/kGZDE8QPZgi7ZmMf8aAfTGvSYx+7tg5GDSO83FNQSVRBq0gkHXQM3
9sE+aCuKnYoZjVzPJ6A0UZV6kGQ9NRTbOoac5KuAFQ/7y39ctbfC2jlYr/ZUkJWF
26+K7NhOCAF6jOT3/gWm3v9k+cEHnxhU5f34TB8f0R//CVj0ZR6iV6rxraG7KOI2
kWHtKA4rr6HEgz7UOs3BbVRbDYl29K8lbsDwFylahGEiMBZIsgaL1EcjUcV92GdW
TEmgZIlbhkGF9S8bi7gwxMby7jcA3ay7n0vQA2tDL81vHmMf9oZRTiwEigc33Tng
Dul2pD53pB2+c3FtywFngmigIBwl9hWnVduJ4bUmHADN4wnqQiZDqKqjUBMTKLhT
gFgbjNneSBJlY0J+jh2Sf2/XUTvT+8GlZeoHeR7ITOc5ib2OCEWf4YvPRG0vNPUf
Aix4IY8Lz1Z4LBk7RQtupGVJfvvGgch8hr/mDx5hENvy2zyh0yULWB9gDzOzEfmy
XgWUHUmpTtMLax1TkVS2UeEg9g0bUSyu/Gq9rm8gMx4C8yONAXjKwbUYXs9IwF4y
crMS+Jsxh6OGD2IKWxYpi198yjnKOxLIPYvHIaWaKy50vdZsFEoOguIJOC1ROa6B
lsLXWysiXAOflNXuqMQy9RQ6wdpnaRyFI8xAXg4gGVFYI6nqVDit1Xt8za1BwLX5
TeY59PSBsFlh5A4OBhn071iUP8SrJ4a+e7D+mlgBAQNsi8B4bObaUwnwphI+Bh8q
akoxhgFP1rOueh4yAP66s8KM4gM9l64UAbdL7sxYbfPNYxGU4TWADGCg0vHKtrrC
bafwuMMC9NhGEPJXDY6WT/ZNkURuwAmaVao/h4RX5kpBYxNQGshfrYVJ1iearO2E
z8UoYJcc9AVTk++tBw4ADLmHUcQVF14o0PuaQKBJIVMwUssa/JvCBbxdaVKWhAJt
Pcb6Xg5JuOFmmhv/s+iWvsG9HrImDO0uAvqbvj3nhqnVrq3881YR2hqPsRpul/wp
ySvingPiM4yoOIzHlOEiEAcdlrZ6p+xdInx3wW5SKze8xP8qndPfTgqC6pS3F6Uf
RoYeI4+q6KrPJtOxMH33m5Py8tFm4P7uZ+G5VpIHqeyjBAKvYOHXKxkRrdJQUGsU
WCcdxjDeAwn3kwxt4w2rMVwBmzl97XRg/H/bd9oL+kcd9SVdNF8flkqvtGcbrRAc
UOm9lKrhse1H3O7hqjlq9U8MIle43acs7YsYWULMPGjAnQRcXBA7SdimvHTsCgV3
fhqwL5A6AqqOrjUlCEd00V0tmel3Ywr1nx2U5QHT/zLwJ4CqbiMEjsGGZYOT8d3W
gj/tj/z+MgeKgjJJFcgDlcmtilPjQGLNPLX4V2ec6AqClnBTr/J7iyO3OTpv+/ed
zLNZjPXw5LNJ3L82Penby8101ZRf52TNp/igOGR1EL710vVu1DBbOMdcPcnFXgp0
Zbsig/vajp8LieX0S4ZiiMy8Rav9a6Zd5++Vp6PgN5KFq40DfVBYaDDxZ3olmyQH
N4orWmPIwhhqpVbRz9VabMk4AfJva5b9Db8WZIy2Zo45nn6/SENuLR3twboojOrK
n0bnmZ/9AOJC7IMHv/sHB8x50DivLoHhZnqBOi3DTjMkFOeGpOlMhi6n7sN9l611
MCwETeOc3RuSibXotkHSK9R3We1hVcHiuGVJFIXtDRc=
`protect END_PROTECTED
