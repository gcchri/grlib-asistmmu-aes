`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u8gQ60r5+m8g6ID03vVatImvR4+61vwa+EydER7vZ5SC8XZwJ89NrUz6n6gyy1nA
HpSYWxZEXK+A/BxIMZBR2mXrjuWJoG824rC978jbbJ2OoBTxT2ELpuOogDCXtkdm
MT2V5tRr2jztRgTZ7LPjXC30do6zioFrV4iDZ2SBboUes90jyLdXRiWcMAfg9ew0
F9l3SsJnMmcQE4n9UFEWQUMGPwj/CSzryDj+PXmeHWYXL9qpSjOo4GJ81OmKO1pM
YvsULN/wE8wGWhCQWCCvqCaC1BicXmdGTdzUzNydgpIRn1z762tK6/qpYSy6iJnS
Yo80rmxWcbJLQAYdP8N5zF4uxIyV/wahVC4tbWt9SGJH2R1qfc//J+j3BdgoMO+a
nrRkZe410aRgjBQQURFlE447p/RjNH+D7kRmHHfSNVKXVBTZeahfhrF+lfKgcnB/
lWe2AOA5OTa6WAO8x4DKiwPGrzWuq1OGqAL8fX86kckiEU0SIDKqez6LgAw6HlqN
D+QXh9cD9hZu4WBLttB0eH8Emfu/imd6UZ4D51PcS6wiO3wQ7uPLjlMyTSYcHtOU
ILWxbdnwpqZrAAJtEtrAhqZgYZW3CkoTDeWAxP8LzQbOEFp1VrIHeSvkbtzA4sZI
xl6ypUKUpY2AKhqf9cGpbfJKgBQMT1MOl4BFZs+NVkQsKVJYgEX8Ez+R7T2JpKfw
KaqDWj/w2QosKtJ4gEM+VRYT+CtvPLWPoiC27AGPWqcjqHENVYzhzdG1PI+aymlS
O4XdSF1uO6e/bnzH0k8DujoJGi+AzJfFb+tvfHxAfh1u7B3Z8MSRvGkeYQshuSK/
LUJH8Y6eo6KvEJPHb6p/w/aCwwwTerU0whKBBIEH0TBxlb0tgpZDVP9Zf60OO8Hp
vDTphxH2sUfUWADZvCKoLLyIj1wQh8rgxlQuDQKtGK9n4D///qGEcxcHkQn1rR9E
okciSnptFibQK8fnr5pP2JHLo6LF8zBGO4UPsoSgg/Ne9gFnwIY7bGJSjatZYUVz
2zLAQxyacpWxs0JK3+n1jMq4QW+GPMrUDNo7vMIzuWygdPzMMEr7p+eYgoLHAba4
ch+lkxxXu1r2OtZkLMSnue5VWKAg29NX6xJ9MRs6R6R5PST+ed0EeumjzNoWDpQD
S2Vr28dwrvgIGGAvCBC8OZAsiNRHpJEYzjTdu7lbww+Ad3IPTffAc6N+p40zWNN7
VgPp6lwmTg1UV8bobOn2VBo7yxUcAo9zj0zOIdOlrh4oILO83u1h0v5bSaooSzO5
mFc/EosNGPSWYkUfORZDSEv9o5TU0FMNZqFlstRmNgTh9T01uAoxGB4f6mEl67GB
hgnE3GlxZLl9kUMKHd8NIYOkUJvgMvupx/5AVj0JR2vghu4ehXSVpXUUIVvrcKD4
IbISWw1Fukeh0DuctsWE9+iDZN0BgFruw9wDUZtbwq3wNeV/+5nhaotZ+M6Cb+97
jUPgb7h1GMb4aEa47WVPRy36oUF8ZBdH9QUR8/A4HQ9kne10TW0brLOpnsiqKy6z
ltqPtPZQWlPkzCV/Z6s1w+RHsYYlq6nD15lVYKIDkrAlV9PLNAQ8rKb0yaNIFpue
swogVRjR/b7yXwvZFSy1ZOVqCIrVpWqeCLa/r4Eb/r+JfZfvyyuHbETF3ybS3g9w
Qax5EYkZhFpeMD5SBgFKNBFRVn9IewWSOlxJFNjT8CjW/pGSVIaaWrOqKex1BD6g
k6GmIz4onWGVT5W1gFSggwF+Hewz043aWRi/rMCPWZMZIa12RpWZOA/oZEOOwFJb
MNarhbJJ28+wZrv9b9LIyFlU0Y1BZrSV958BZgF2mLNXcl7b2JCfQKvHoYE1IcQW
iXtKfvJ/SDgtQh4+wN92ufwGKeMt8chK97RdO70ox44kwPNl+lpmlQOVQ1nWSX2C
DeoW/AqNUlCn8T8zNbx0klRqqFkhzvxWVdTLGJSjy0Oyk97RvW/8iO4ymxlGnNUm
e0JhbFGUPUA01PqfpkKzlrb3QSdT0OGWF3bV2pUxgzwdHN1IqIVS1SvusB5iiR53
6n32Z94xl9a8iGjSnj6m/EKfwn6xZ1QxO43g9mst1QFMFjZqPl9ovxEwP1TBoa9U
7r88AouUsZOCx1RVqNdwgsGWST2ymskMLuHzKweemQtKm7oOpXeRqpsLpWnotxNx
pYYM9jbcZiVFKAx+uVPcBOdYLsK/w9N84bWXsKBBAYfKU/YXvKrxzs/csi/lYqHM
ATflhLUnQUF9wNiUIHZbgvIoptPs2dlI5xIrYz+4wwogIPA5svbT2vWiiSKa5pmi
ybD7sNoMdDBaM2Qf/FX20Y9trekqgLM17oN6Xb11ahU9K45V7x9UdbwDIq/zRz9+
lHRnpzIpnBF3MClfId1oTI8S7ytlRm6hDnsWIBwelpf8zgqGuBBjYFOmurGW1Qtj
HB9GhRj3Gccjkr8bV6S09dbc4xWOz4ctOKy1XHSlyiNoxhlaW8PY+Srt0uSx4e1l
Wr9dfVw77ZjDU6TXnNqGp25v9xqmRw+4KIk4s4temyCYkMYjpU3LlekoYuBu3vTM
DHyWMf1J8HtuB6inVCx5r897oi8l42ZOqg6/+gDy/vRzC52RXWmJ8kYPRWh2qjwt
tl8Dn3nHkcFmjhXsniFeDxb+A1RkDexPSThmA436NXXvBCp3jQU9PKaD1ooyxX0F
Ilr4XrOUG3shGNO5FuogwYDGy6HDAoNBrsNVbBcAW4eUaXyNsU+l9Rk5mrLRq822
DtsypVVOyxq4Gx0tQ/9KghLR4Ps0vnAL5ja/RivCLJYFr6QK5fdt1yiSdV/4NIZt
QX8KXEMqQaPas3o4rvMMm8aolD3N8I5WZTVQ7t1EAHsi73pGozC5qISOLTJsvYe0
WnHb3yv+RAVsr22aYfrojH1dxYzzH1mZNDaUjdMa8hV8SNWIz6/NWMoVxgkNuP0g
DgWbcwfO38VxF9cOfJHFBKEqqyJKEoLcxFMiEST/FBjVqgKgZZ06C1P7cXvCbcDM
KVYzcBuk/FvyxEZK+CsYySO6j0YphCdOk6z46FyMObokXs4c3nmCL9s1Mc2w8SBL
udPISDQ8Wb/3U+3dzMvB6/o5JxqylQdHH7EpwEXW5i0Ltj3NhQw2digW3VLao7Bd
29YFzZ1JsA94ImbIqYOiUVwdxhY1oZdz6/YUQd8yqc6X7WC9xOn+GYayd8rPKufq
yFUc/KVzqeKFiED92XmxqJyJ8G6YhAyC7bquKfZJQurTZcqyz6Z8RNp5fD+pazFV
VIRH0/5fYPWtr9qY3Xn9cfwF73yxUMj0mWwrXb0wiFdDUq+y59R4yv06/4xgVFV/
zbsIuoweuNmMxx0ooPBajnoQ62GOY8i5h4DR8o4tZdEpDO3hCdUR3nfsd3jYlS4J
tmdTxUVrRiTW89vXiRGnXGGDcz9retBElty9YTb4zpJ/UHLOA2cCWGTPhYmQSuxq
8rnVinOTKCzIXes/+mAFNkdyoEJJ1htFvB/8RcfyPvnkfssstsI0MFSnmeNV5IFM
ryzQgAY9j8XIkU6mFzsSyGa91w65wqMykD8akLVmG1/SGdg8m1nbTtLmmg5yPGLS
NRq/yXVd6Y/1psc6mp4lrL96rDzrKb1UmpbbcDzqDZVRkeKQ+t+SDFwLQ7xRn7OY
QHzFjoagnru92/HzPkO3mou1vG+xRrvLgx0TWFwayqt3GThI+Rhb4ZuqThyz9UDU
+ycTJML6rvNJKcq+oJBAQIQH4lbQq6jCOemthKBY4TnWLiT2FosyoT3g+TCb0EC5
1MxAdS7IJ/8AfijvXb9LOG5BAsTisWSgxCHNZ3P2uQv6SKrrQmrTlq4h1cuxcrN0
O5Zd7w6JTdUbQpoRHWon8dFL+ytCzerSxRYsVwYGtQ4TutKLw9gyR72FlgESzWl3
wvKXhkibf2xPTQGSVp13BfaxT2rGbRSbp20HSKuKhlTPtb5w5v85rJ+gMGUHw96p
h6uXFYLC058B5hi2+AHIcpyHfFDfv4GYcM5BtCBHD/S3drsSf5QrCn9zPdO9/lMk
n7Qf2pZbwahi5x4nfzsy0fJaBokoQIaqKhlDtvxlBYVcmyN3peQzerq4/qdE55yV
hHkuZ9YDHKCRL3Fp9W6cJNL7DlkAbtbnfzE3kaR/5qwCUrm6aUT4ijGeZ6yB/ho5
0gJ+n1yVD26pDuEj2Jufm5sU5Chcy4A7o7QDPkYgP0Nd3R/w3/Ikx4FTO/goWUTq
8hyPChtIhO5RmBG7zNM9hB3lQuuvwNZ7jf9J7ulZpRyWgFROyWlMcRJ5dPaPnqhF
5ODiA0DDxJQutzzHY8g5u+6kEzv9wN6r6S8taEFtYKc7dmkjvh53QrthH58Qyp2e
LJe2u5U4CcS/YmBhoa/4s6qPU0OauzRqXmkfkfFeEmdZHqSfzHxW8evRJixvPkP5
r1c55qpE/jQNDLMVo26M6IGXnp4+kb0cU8swWrmmePsLP2RA88902JUh02TK/FgG
nWOqdxF19lW0myXkK9XrGKRq8GKwkveTyGLw9DyhdgFjZyQBOtuYNh9A7sod7IaI
BZpCLCkM84XlsxMneu2XzryoVPMyvHN6YOBtmkDVVTEc4L/QrTKdRsUCmZkiI1XM
c/5ioy3/Ie9Qp7vG3L9i+RbnbenhjxAQ5sJOzyjmT76YrlFt7zWfAuyfT3i+q8RI
154VewhpAcNKAIgMofKaf5BGIVuVITLTZFUPIelIh1MP6DbXWcwOnvUk/Es3op4X
ArPu2E4bo6YVT0OVcB0WKEDFZXb+Z6LUJbhJZlFLJZ2hDjXCkIWVjad8aqZPYD35
BSb8TNZjXBqCWtKLAJS+b/RtBvcZr8pqxgXArYyORJ2CxtGaErIBjmD784WCLRhK
9utPrEBqZGF3yDZpCr/gcCP9Wi8KNRaxOPwc5s5EIqA7QG2J06gMTSY2XjFp/HkO
lstDvKmSzBGXQO3zfPBBG2846ID3eJIfyOit1NOBuZ5KgkDamjxqrmaf2s08BVtU
NRDRboqN8Xt7ja1W5J/f38pWHQNhMXkCssZG5xA1Gwih4J2GC6zhXIFzfEzH9u0e
O5L+U0627/gtrCDNXucx8cvHHoxiJamOg4WSQe1x+9p7W6fVC6cqEvdrLQtFy0XT
vmlEDfBy/0iWNb/eWwk/sRruS31FePtNGp/A/OFVV28SlA8+OpFYJOvZdof4ywtZ
jaYJfZc8H4VkJVlP+3I2CNhoJkh0eaeNj3kcfiowhgq804tCTmBAioQZEzCSOiGk
mvITmrU2GoF9ya1unfr1FtU9ZQawlc6H0qKc+kGcYNa+CV/V2p6MQg0Eah2P84aZ
wMBm6qCXAIGvYeWonu174BP/4atzpkjc/+popDQZpT+u+5LwVotn/EvETR8AO5bo
shEetHW53GXwsAYRaOuQ2Bh4UVS72kDGUp5c1doenQ7182kS1w/N82QV8Uh4vVvB
WG3a73CGIWVNqHacI0nNYGm0Mooa3MoM4LDzCer/zToGJAJyAGYCaKYyVJiTo1Mf
njPcAivfuetIlo51eB9452FuToCkceNszZpvP3xA6Xozv6/e7HZ6Lr2dWL3G5soi
EYs/8Ko9zmLfXc78GaGbuxcc2ep/7GMs/aAQ3vPw4an944IRgghcB2kyxsJNmuda
ftD7LacOIWkSB+0/DvUIig1t7RVHK7G8BRe3a41ICDtrtSWoG/3o0+gdPVSKBaoq
qUoUoC3BD2BGUCLy7EDwCLmxHsYR9rDH3vdOUkczT6nf+Fe4mtpC10JACQoqbon8
PsQ4rWoeioAHxcBeeb3J88kVf5iR7LmojqiQlTzYCY/e/Qvju+4Av1S6Tqi1xNsN
Y1Mh/XMKg4w6HwxwrxD4O5KpCaN+DyAEsW1dpv8gXm6T07ebw2kLYrw7cAuNov0K
u44FFs0lLjezk1/RqKOCnFfYzldy/hfIi/ROdSOw1f4Jf/34U0O0anumZPgkQbX1
kCFkPaydnFQGA+bzy7yi/8H2e+S3F511QxuKnSPu323dpk6dTZT36/IrOGVyKJtM
tgL+8BTvtBOR4bVIZ607eJjImduFXqe2TkymiFV7Ni3gb6z9SnLvnu8ePV1pTy4J
vtVhwP+YecMhWfBDihvxt/pEHadWspj53xNqI8NjRMWSKuewHRDeA0J5MVCEsP2T
BaIi6Ch0oeU//3cfJ6HdQ0pQozFJb6FLGEuh5ajcnDcuJe1wqFbCa9ja04tAmrSI
wSx1dmdvnB2h9JFjEHzTLdW/NeKinXkHWE0AZE33ZUcREPoikX5WObd7XPupOMWJ
+OLQlyXNi06hcPODUIa6oi7jsfQI8KhaNgCXGQ+FN+PLJwoeNhInobBdX8OqiDUP
q1A5eXX3cqykUko1wwmNN6dy3ma6jQH3WRLSQRw0r2xVmVi1MazHIh3MzFpy31iq
nZ1fGt0S6pLzJh1Q+LgQS+6PEPJ2ZLJjvq6rJSreWkFWE+ehuZ6OOim0xjL0VPDM
iJzg6MMjc8Ojmru5f99ITwmPqqqVpyb9chx3Mc7k7qz0jvzKoQOHEUgywJJ/AQyk
fMzm0BOs9sAVZa1RwhpBakPScga/RlfzgY7zTVByhOTbf+uhjyt98eXJwzdUerSB
cwUnyk0Apga0X2Jq+s4BDN8jSMMfOFnLQ8wxS9zg3MA5lgPvz9obd/dlZhoLf1YZ
2YqZ6N62oqyeFceD/HI/sEN5pGIUjoZxQ5xw1NCo2jaRXEMS5h40YPH/CMkWjp78
Qrg5dDPxm5CG3D/54dwPQpB5uH91DLPbXdsVKvkH4ZMc1o3eUS283e+AeyAP6K0a
0twOfNzdEvE2m77OHUmoOY52D6gi6RCr4buQKzHoCb01bd2UugcZeQvJLAYG2rCQ
TIrHVDHpD465x4xkqiThgc5+lzs430e2TF7L/5WwS0fyUwk+39PcRhcxO6sTdyx1
BOxhWQUFPr3mrlxfP3OG2AkMWOJ2dx3YHchxP4bn2kONSgrp0pyu62CcKMCRhDuS
w4SdKmZBL5t0CwRSXLJwv7hAqjuB5bvPogS5Elbio6ET0uXem2K78Su7Yk1+1Ueo
C8hdQYkeQZtAzxzfSfGxLS1psqgLii6ZU2So/4P3XcTL4LVPLX18UHVNvqR0aM4I
bVE1Dedd9H3MthmYGDCLZkvTOUe3+v4uHn9rkz40pXU1OeXM6mRRmQj2qA0jiYfK
9n5bwXUzkfEKfcfAQ9tZvTeyoabO1pYWO7afBQmIyJsXaNIo+r2sp2aGgB9bjasK
LD+Ur80cZAR59O7SqMp9Sx1QPaSKCQFhqcOm7EjkZku7I7YNlzIGnFakCekvTx2U
ikj/jhOYg4PQS/PrxqCwW9StHV9hByn4hNJUcHiZSaOHm4GV+yo0W69IWmALJ2jx
zTGdGy98i+WFbHe80s56ZbHiaDs1JVIdAMdbq4TwaGbHPwcOje7zX59LVOowarta
56s7UI/9oVKpuM8jRutEaW6YZOOm8wL648S5SUGLFD+iApWh3rudtYeGKLKwd61u
3+rwxIF991G4w0btfLy5Aknk61OCIlHTPQ/Z8fwaNGVOhz0iy5gm5S8/ztzwYdky
cRjDo2Z6ifJc4uZaXLjkjqIhB1Jx4nT15la6bBZJpFsidbRlSPU1fES+29cNo+wA
8v8z8rv3OFKsYa0vnxgSJJO9iVy7c+7g95Ezsuql4iEvXF6yC1ozJfvCXMZ8kQ1x
hFwW9KtB/n/ZIjQFSfEx6qxW0hInLY41b2Z5NkY8jHJOC5sD0ZduoTgzKVD5Q7G0
7yObPwxy5bY8p6DCq0L0kvnnTlZbtMagNl/fShoyoSVfdUyh0r7NtsHEsAeC8our
uoeZ7asSqz3/kacalxP00CffKdYazPib/s0oM5ssSuTjfPEpwQDPq9YAoGOaEFHP
P8TNMKTrRt+iLuG+RTj/DZwvo6se+LoBtAXfzZ4Eg9ymz6fKdR19E3Fuvav6jU2q
NVhG/3DlxaODPHnL9txbSnb4FvqDJjhstOt3VaWaO/dg0Fu0ft2hJndoKzGd8ZfK
JsEgxMH/yZ8JvUFOTCNSs7qtHOG2j8hFBqXhVCFUd7k4mpV6ExqIrxjtXwwSTPKJ
ppfvMrzDpHxzXPq+JKyFYWSjOZgf7VsR9OJDpkH3mSmFidIy1EGgFSPYMoK5Fxqb
BxDGuHqhhsbzPxbQU1rLgtK4yKBk8mT3ZWq7MmqTEFaxaP2i81znnqj4UhNsbu5X
gMrCUnrqG9fcrUMNgZ1jjDmXS7mi0pRM0WR7rRu/s60+g2Jq3cNXFS2ElUvignWu
a7r2Q9tRKP49RAFa1rdjdiKqbG54+4o0xMdCNq30uQBjmqw6r6leHXKUry8YaDq7
I7b8CNs9cdimltJSmfP/FXsoTSMshCPkGMpmiMZNnohFlCyJBXq0zwoIAgENCpBb
jhAbzBjzkwYh6zjrfNqAS4NguFOUnEgu269VeQj8cYisauIdmFsA2F7qsEAS/XNx
796UyDYG4dYAKlKXy8DhLPmSBLDwF8DfGupAps6qOA335TRX3Tvr/Px/ricz6oa3
1YQM81yD9SiNkAS7b0Sp/znfJQuXlpB0W5xrCyxMASsSnc7KUbZuxGn4HkWRZ0HK
UgzkhRLH1sNuVVLE6UVzXaxPhKIFy4a9yXGpWMJNbs+kzqUndQ/I5ChanxT+xfNU
20bfbSiXaVJiE4f0fRf8yn+W1RNdoCRaJBK4lV2+CMCLSk6d3BU1oG4BZ3b87QEb
vvbA/ZhBe0e04FWkKm1MTlH547z2AUNOVP5Lymd9SX5SCVNZKCYwZd3pPNmV+KuI
K8yP+8yDzTPRHL9GMwhG+TinY5l0IQ4/uTpvJ7eiw62XtYeCZVtCBnyX+5jlvUwE
mAZI+GilWt2OShak/CsQaLQGei9/v1nm+LLqkUST9DYhYWp3xMCkBMrIOfmpYAnB
EVzHPdDEIjXRLU7/rBoI/BM17o+3oSogG6iC/eCfzBqLRMzx3ndcKUFAT2Ey8gkq
VdOUwrLmgIDjuThIqfykQhyn+av5YlKdzdwuZVa2GG53nTbonr5S2nwg1ckY5Amb
uVdpm1GEqMMjuWJ+XIr6p0IoYBgfZB+CbND6xTr8cfDNu8aE6tudQczvmzgrrMZ/
xXtXC+1lTdK1Heg0KWyCwHrPoyBI1dKpzLCTppUUsIE6MUozEHvMdxhay6FwvU71
LbvEJytG/eSVXo1Sk6Ed5lBIPtU7Q4KKBR+2ab3OPjs8NQpAmjm4CLXdoKs3AMlr
wRf8sfwUbt0fTwWneVxJ2tor6XfLhP7eJ/edRqZYMk4sVfc1B6zXNAd/CX47O40T
nSEEVqn+Ft7ClOuYe+zBsW6S+fD1EaLu+YSp7mFp5PiGagSQw8UwKGkArHboVHmP
BDtdjy//CPFuKTV0NdfwMQMhRlTdikbgTTFFAPVW3bCscz7stg+lCr2jVeTQX33E
2Ar5i3zUd695sHdsd2kG0dAh6KkQpV1yyDIQx/DZt7bx2v0gVx6HrxHkOHLwrxLd
R0QUE6VuIh2IuS44fn2VeNstP+6Cj6NTtmBxo2jIq7jCh11GFHQyLzZUgUweigyY
uXh+GUyKbDDiN4vYlKW40Iyf9Lc4dxTlCdKaKmsTcPg1xPbjK4OFAWUVsP8b6bwq
OocWkxhiUSmgpkt/K+NRpYwELi8BTteoY+Oh1OqKfWebblmeLEAWVYLkB0v8FvUZ
0hiktq5UWDdtWqn+3wz+TIGquvwrOxtQ/DAwDmiY6Ay+izv7yJ4Wf/Zkdt3DaVJA
C7NVef65p+61uqo/dZwVd9bTsDzNx58LyOXUKt4tXQgKtYdNkTdjGchOoKOmhGbm
tRp5MxuWLqLUlDIRpgffeAV02FTtUiK1Av1HWV3MC2asytSLHSiVb2NnTsIQCzQq
KpjNXIyMYlBQF3zZDPuFYgZbsn06xZeL7L/A5bZYSMau86xNwCs40eFwgKvIthLO
KgW/C48wrWJhY5GrPLcoq+aC+GKt7Q/rJILbJy6dt8K15U6JxUwbQHby5V4OKL0V
MzkHpZMtuviPKikY6hd/r/GCkiw78eqFkp2hIiunbbdJGl0ccpo3+BdYcLuUUlxF
1w7Rdpe9vXk5e1f9QGUtW9kJxgyubLFVZfqqaxqpP26tnAD+sDvXMHCfN4xiiU4y
yTnkv5VoE0NxbigOI71EQmDnZypz4/1APO7q9xBsy8hcnLRY7fRKi8UEZYJrGMsB
qna23BjaTCg3S6EnxvND42L2HW0ayhulJHuCH43h/FXSfawIBw0LSwrGxIrwFwu9
oipah6L/67W85LXiRVaZJFti6rSNeiIZEYTHVdwon6eMZQWaFlepfeDIVpNixeNq
fowlq9FZ5rrA+bVdo4aNUDnuah/+vNFatN5XUI+iISAPtubJdiRnvaDhlwO99/bs
AACoYJJ1JfX42Tk5EXFr2i0xBufcQo8Tqra1iR9byi4BW2It1SjbTNMZUKFy6u25
Q9Ho2QcKO0nvxDV9zJ4IqXpEPmia+mzUuxYF1Iu/IxJdqvlMiSbxfJtpsIL/Hwx8
+uPufeYBMnS7VF51AvrIZjb7cxLZpOmYSDcupA0OVXS8Cb5GhpsnqEsl/OE59FyW
/r8Q3hHz76ruP3BbV7lCAndJpjmSV+mAXOOvbwsgtVeuy1KyxEqhI6gtFuDh14rw
yp7+kDGRu+7i9RhbQlsCgWHUTwrR6ziSHo+6nslHEN6Y6xG3PVLSakShMAAThm7K
XSfmSGeKkv3cZyP4MQcVhaJFAdQncUFiJN893az20Pvl4G3ogajfDrg9UJZTUPXZ
ahf5olw3MWqSJhfadJ+uNaWbT66svW0y4NqWXLKlQXl80lXNKbBvesm0mp8jDyO5
sHL/8LzBLr+9NDPw8DXMipONcNZGp+e8k+ct3YImTt8FXMMISfHX0cueb/o44obj
jL4DVCFkYvoj4Xq27SGsdt6aljua8Ox2K/Dx+skWOoEupYE+nqcoQAFsi+khkPvH
9bihjgaHTrk13OywRLKIKHiNmx94MtNjKToCE9j7Cz6smcEIKUeMbiwO7kNUwvoJ
2qNtMEGt/FWEj/Fjh0O0VSLyTLFFFfSe+ZnSfoEk5n+9XtJqqBDqw/B+x21umhew
qbeJfK9UFb1uAM5R/+3T54uvfkzaGMz8X2apx1j4QBWrmXxqqLYzQ8PQyLFLcov+
8/NNQpy2vEjZb2tzpY1XfmJ0APMHmwOHFTmfX0D9ScZR13SWMhVMYo3SyP+y8LN2
6S6VhXR4+FEEnfcOBnNM7q7j/fzX0xfRPIjO7AxOgr00/IxSOY5FPDu4hN01XhLJ
FgqyaWWjPQ7iNW9KgAvFftaMQ3gAXwyWau0K5/ZZ9NcQu0EvqjutgL8Hicryacwu
9lQaN/lyIPER4spAuquhmVTNrflTQ8qklmG6Qd7R7oPoerZ9RZXSk2P96r+1T8za
AAqaoWhOH9+ccd8gyFSz+V9vzPELKBJhdT0/wTEhr6ig5Vha/f9eG0JojkuB6UEX
O8+k9hmH0bK1Tawdnnd+COefyfkO8qkHf2JbiN72sP7UDWtLzk5Y6qA72uhFTqF7
4de8TGJ5TTB0zRtuL/Lwn6bR7xuhieWqDo4gxdI4ptM+tVhR75G4ejBhVs1n7IKi
n976KeaPLyFtXeGXmHK4FH2qLEXRO/ZibOOFeZZA80cCEjBHIsU4yqQztpaS2ZKa
IVSbm+pftfUFc8fr4G9MX8zvqCA6ITtV4DdUyQLgN1t9JAYjGOvAm80ZrlCbLWhd
sYXvW68w9HdFK46v0PT/GmD00/QUANQlAjQf17VSQjNmqipi9wKB8xpLoErMmPi7
VrJxkUBKypO4fIttC9NiIL2mkL+vh8B61APcGYPxenu2qPc2xkbrzkQ4+S5XqO8N
aSBJe2whneiDxsB7CHACcPh3M6kQdLllZB8YuUk/kz1CXqTlRRRO7droxmsXGQ1s
jiUNu9c7VED5KMFyBt3SVGPyuo0yTpq0ldZaoQDkemiNRy5Bm24xGCXekEHxg1YW
UbH4wgujBEm1KnndaGOjSp3EcP05DUhgjr1P4O2isFQpxJpHrMF3j2SexqtsZ90J
6DRZcBsHvH/5w5KSoZrglGI9lN02dHLc+APRDTLKfPadIrordBKmhYe8ZMt2U35T
Phj9t7bBw8t82UeluQtS4v0vth0Ax+qNuGJw7d7pBQ8j6BVs/cdmmc7IodTNbjXA
Okj+I1T8Ox8fLDNQJ4CiVqwT0kkwsxrfLOMitjEw/ZlWX7zStXsmzJY04CzGOAWl
AYY18HJscwUARPqXeYIwnMpa8NF0oZU9bPnucrko9wCxIRIQhsPrY4wkuAkV5GyE
KMBgfjESn/5YPR4xYFVK0c93FBkkBxa5r3nZXILvd//1bSMvYcXfR1JONNTU6FqW
9T0ntHe2fRTmE7/JRu2Ovvbs6tnXPtH7hmano5uWeF9H3hKx/G4E07GmmyK+KDo1
UbA1MNTWVvRZHR8niw8TfP30uZxY99tE4V/qNeLR4YMiGf0O3FrkDmhU4vP9/NEv
oLnWWzYK0Pbcrw2lVaNrbKMhpbCKQ5wPp8wf60PQfJMON03M0ThHCuuSVIfPDxjJ
J+1bkohnyYk8V1/6GHVsA65uVllkhnSU3ONmhgaSL9j2tgS+veSkGd9yaa2M9v9j
FN21vMU44RcFkqfzxMCYA80qjGm2soEpeDcQJcps1wbDEY2naJhy9r9q3zF4OTMp
bYzhosZtnEX3T5PW+3qxhc3XY6J0Y+zsV9wkQidojPg0qXbS12cmPz3LSxhVnQ8I
V0Mu7M5R0Vn2a0xH19lJsl94lNlDf8QPELbW+h/21pw6legIpqryHMzzWX4PlZYe
oVtZhopTCNPduYw8FY28bvj2Fe6pxJPVslzCV/0jcPUiDvR1sIu9V7x0WJhj6r5d
v04Xgazy0A1vI+ZbBb8De983nI76yk14rIRbsv7SyzL39HYM1CtxzEsp1rak4EXo
qV6LSEK/+ORntcnZDOOPt0+ftLvREY7Fgw6VAaOr/uvGaTud5aSS8xu/oqntykSC
aT06OsRU+ocGyh6Gp+Z20xq8lkreG8m2CrJhtMY/5+bh7S4ydJ8cs67U45bdcYqH
fIAv9Be6O6/l5Vil7VE54f0VORf+9ih+v5jPrAxbsjxrML5JoIoERLr/mdznP9nA
bGKyXuH/4juiU5Tja7IlCapGOWJAThqNhQ8ok0ivb854Rl1803cEwmLc1Ocn/GM+
zNM1kw4snCj03Fd0/aSxnjXqoh7dUICdvu/Ggn5WvdML16T0ElBnufozAVNfIFhC
zbpHzBy5j3FpakLdmOcPdpV2S89xaohRhzP1ORKkULKp1mrrxLMQvXBK+Nopnd4e
jM0QgZsNLi2+crSkNwvZp/2mlMpA7IDOgaj+4GHsEOYDQtPWzMYShfZyWbhhYtcT
tAFw+ciJ1mSkMrOfc3YhfW8D6wngDucr3CK1EO9cL8B1Bjpjntn6vl6ifnkbMitl
q8zCQ68ywSbBv1eHlL6ambtoc/UHCc2dVNxBmnMZjvTvQXY0yx/flMQtExWdfYQA
gpvCpmUABr2PB/04iXazsyml3I9GK3vKDN8XqkaB238ErQiGS0D9m4ZcZZ2V2TMu
NfCvC3KnVH6rhQHgkZKY2EBYXjAfZ61u9ssCL5cDI9M39lvSP7ax1L2f0FwvU1tV
zVeIt6lpsMFha4NNz2vjD8f1ZhECad0zpVay69VqQn/bJXFYst9ZyJ8fpLmapbkJ
d5ALPm8aT49RjgSFlbIpWEFE4HUTutyXROvg3K+eQIi/dlNzQfznsf3pDD80Q2NX
mO4mKkLZugJrNHppGfWbMKxspcjbpHTNni/JEEWhuvHZYdHKrguoDocqGkGtZgqN
bke5u78tkQtWBL+YUSBAp3SIz6Gi7UK/M0/uulc33O9y5G6YpH091wAV0TPh5fuV
iyHQxXGQQwBP3oUAEGrPNugy1N1DABicnI+2mdnRHajOAFVD7mzCGZsCEWTvf4Ct
gGCvXYyNxUSsyzcNjQv4/bfTn9ADmlIHbufvjK4tkHFH0j12AF11KehrXCFMtYSL
YA5aT2hbGxy+zmnnM++N6QAzEVKZ38W2MB3+gY6UvJWQvs22PEba6j5r+jqqjFN/
nlHYJNpNj1SFma7rPBNQPKQlU0cUKrkDaoxXcawXOK3t2jCqcZI3kWx3ZLHETgZu
E/Kk0wapXXOgl/di2mvG5GPX4dkW6fSu2rx4YI2Z53hA1N0TcbcCPDZpF9UJN/P+
Lr4pX4wVXyWQulmZYZUa9bOVtiHONJu1HQoUiAxI509rtvQfGwrN+MBFaxPky/5T
qPEWnqUgdnrNNrMpCO3zK+KKOJ0ryey2/xsvDHjdZEhkwhy99L2j7kOm8l4/3Ied
3PRUakTCaGlxvrwYQZ/J53UiGaempW0y4Fs3RPNhRXlS0MX0R6mWfDOdtLEoE7Y5
YH6oyJpu3VFSY4MoiFa8ZaIJ9MyUpLnFX6vgmfg+jRj5tvnh4ytXBt0dUP25J7Lt
anYFija9nh1lEF3AEnvz9DYVpXaAZi42a70OCnJVsC7WKjF7zfr04b+oNvSJxpqN
RK5MA4hJkT3IQ8uAeiQEts1WjxlKhV+kWKlkFRd5rS8Zdk1V97La47dPVYgRh/+g
fYMUS/IoEL4tKzEnstBU3/EmejUoXhRGBoY3Xoqm+DvOKO7SCLgd0HnXupZQY2E1
wTfGG5KhyK4qeU6FBFSJ9SIzmMfOb56Y4PsKY6mWMFzfociFgMosHoncNt/3o9jE
fkaf7a15CEVXeNal6TsIFbjo4NrP4eyERN13qPKtXCDWRVnx1JpTFCwCYawGuwP0
CoZPD264J+3NR3D8dQ+FyzljwC+onCQTi9nfWnFDowpY93e/Lg9OR3AbxzBOX82G
xIwJtEGR1ISFyMIPvSljuSmW1enVI9FsZv35zBDpRBbhOGx3VdpMTQdYlUXSZnIU
rucrcK0iPaDlb/znNw9EhF0McR2izavTW5uLhL6bhLyOAAE9aNf3+MsMEue8CLH8
TT86cUAusfMTefBkoBnwbDZCkM82O8mJ38uRJXKKDMEAMnbmNo9AGwwCCALFe+n9
xJSptZCGIxJ0949XH0AHkFRSt1u/Zn2+qDyVDQtWRHAVzrNfXE71a+stJbc5ij4w
hble3pE6g3rGZLkYaSx9SvwKzNGDt/v4msz0e2lR5aMFqeM3JWM+Iua64nJqzJdz
P9nnj72S6e5psxtCrZMubrbp0HC8d03PUxW5FfbUaOcC6Tol5cQYip12KvtvC5jf
DedkPTFUwWbq8do5wVkVkFqF+CgPcInTmxoUveNaHXVqP1fy9B3TkQPeQuvGXWcB
iSAUafU8oGVXVJVnzAABPpy4MA8Qgwk/H5QEQyy9tXbAsc/eEBMbhl1df2e+Iq6S
YiySneeDV79UmyDAjMFJr1ors//tk/wQyg2fxgV+6/hRyFCxLD+y9uni4fbfEmC+
9K8f74uMSRmagYftMjAeTvQcT9u16oZJrK42Rd4lLTBmgjipW0LwPlCqCSWowU6v
hvrs8eq0im+zlw2k4q2Ul3uSKPEP/B6GVZkG0zB5XMwkkDpObhMc5I4Tx2cNYfFc
O3RYtPKhg21twrEbzFhUdqBJvUomtbCpGQfqKn70hXbwIx8K9htoTV/BnHWzsfgs
tfVLTPaEhDR8A+GIyTtnbGKu9wLd+0HMVv21N6RLoeYbai72HloEQhbL+tLrJuMY
7aKnD2lGGdQfCsyp2dklXFYedPtVAG3a9AJv3dVTTqrrrEdVwj8kNaWj/jQZdIBb
uVR/jYK965NdTOzwjgjVE+p5xHincYDO4gTr+1NinmIKN/DMqK34FUJ1jBG7vF0h
xt/0r+ZjGwJBFYh7cs8rDCRLctVvf0hTYu0ZWShNon4K9ut1srKYwYxwfnWTStPa
n30bqfJGs6r1ZOZnLKZuRF7enCwQpwq/N6r/PcoCJiMjY07qlCaz7l4hhfYscHza
LuFidvUCB+UoimSjowLML7Hn+g/8kOaFoiqB4xy/yDVt55vIHkJ7cCjmafYgdf7Q
GzpmX12hZBW4pMiinCcva785ti1D1HzEPf6ag8+kdDGm16B0fgoGpXdXJNY2SW5P
k3joshqB3rVowgGRWnf/r+/esb0gs1Pv1GIqQ6iHwr6bItxJn2TGzWbPRoKKEGoX
ULMeChqrtWb6tSe0vO3xpUkdmsPh75SZCfM4/TGQBFSnAStqOtPunVJZnSFH/5tu
wWH9T0hSVgRkLRCp4WNFwDExPZG3UdmrCSplGP98EtGCCk8NIpJ3BK8HKH9BYqtB
oET7c/rc9qz/qxJCxgitoN52NNzR8DKnkZhLa4JN5keYZz/J2YuE7YEPssf9ccFj
8l4tEBIhkLGumZwkehUCcpp7fLWmSVn8yTHRvds24C1bdWwjKY4Parwa4sxkEsHc
Ur9zxceFORrQ36Kku+8aPb38oS2OnBe/13vtSCdK/MG5T0fEelfh9nJodZMG8tY3
shU49xmgSqOqCqpj1ZkCg4LOl0yZljS6qujDHqgeU5BHhaKhL4xIKD3HRRu6oR3g
JUrovwfDtS6wwuXJi0k3VNud+hxeoUFUkkze/gEbgtWpIr/gzDvmNcS+kimG5Y68
GrHtLMc4ZhJjqAgV5TPNcNrZsAPAc3LOJBf1zhreBNYogbR9UvJQiiBLru0JfF2e
lq/+Ui2Q1W0/HM8VKuilnQ4zgDKlO9JxOq4XMi8EA2hSUbXHGmOJydG50EMOtzEK
5zQ9lJ2+A6qgHCkLt1ocT7HgHmBPRjkB9u0kyg7jCbjjvqghtJvzPu7BwzYBp9gb
peRJ9Vm24B2WVJYFfp/QgJajSB3DGkj5Eh+nY0V2Yd7PrS+haqgRGDJm5+nnya6Q
WCPvBVVQuUuqG9AiKFqEu3b4KQr98w6ydmbtK21QY6XRe9US01+5Gelc+D4j5QrJ
eXT29cx6aFSXVY5k/DngGxiP6/tqEiavdRG4xORtmorSRR0dM8HijURJ+xaGZRiQ
+PUNK5p1G2HoePiGnFJZnAGXFwXFmCAAxVtnRK6BTOfRulRfMq8g4b9bVV6z8zLm
3guxND3bRwVlC/zwufjCSPwTcVh1sfNGhTymbkeZTPOWiH/Ebx/DmNCz/6sXGZO6
BU5DfwOm0+Nb7wzC+S/olgRt5vJAHThuaPAfkKTHLldSKauWUySEba3k2WBajwFx
aYc2drbwHca4bf5CvxetEl2OmvHFsAwsluh3ite7isQfY+wlPKSAgvkAYUoYy8oh
lG13vanIaSS5qeflZtcMaM3jw8XCRaXF5IZFiHX3SSg+ncJ3JOSEUeeaSZUflNB+
frbX5MDBUnQZODks/UY44S0ZGmBHfEDKObAF+ZwKl5RiSyIeB6tVysZRAgxbl3qM
u+/4UU32Ruz+L8qQ67ja4AguhUdc1Lep+DsR2xwshKT+mQguFP2HNUIwzJUG7hfu
5pKKTmkWxT0uSvtgpt61uIWXCQnL6LpjoqXeSMil0vcNA9MmVkk9P5NbA4OiFSFw
HwjkWokCzXwrEXrWAsc0rKpqBk4jC/IHK/oGJ+T8QHOmxEkdfBQYkrx536nuThU7
2mxorjC33UGqSLDvq+kVtEsYWm0luQP7VEBn+uRiLDe/qkv8ZwMZ14rshtb8rTQS
Xsm+3judApC8XF+oakhDGvCMjgEcuDYDu7L105tZJTdhbUWp/Ag3c4SdOeCRZPba
zYIxk8LDJNIzNheMmloGO1bCAuZdSnP282+wStXivnMcxnGKZGc+pBojDwbKqSZY
+dpnKTw1bCBTRC7Y1uOu0N9qvx6/1XtF8HIQB1YcsY+FneaFb6aQ53l+vWxv6bgP
8mJPAdq5kKpKk+1tuMU8ALMUp9IIJD25sO1Ss7zMrlHL52dNUrhqrTk0pKxhFr2y
AA1HZr9xgs8BBfAW41awT2ZXLGCATlilA/60ywzZzIm5vbVLRTF3EAwB35gpnVbZ
ilg7pPAC6KwepE2zodxP644ipEKacOYUKDGuzZgBbpsBWUqsvGTVkREllU+6cDep
AYjq0psiwJjy1iqNWL9aYR8n09/Q83MSOnR9URTysM70E72Rzhggw1zN+2Au/r4B
eZDAmmoAsUnRZ156cUli95NTs7+ZdTszs4WLBTQvlXAvvtLYJACuM3AfMvDrEpxJ
EwfG1BBETZY4ghuDUcKnlgulEqId0ROupl5I1XVB1xAQRomN8rxNbn2tbQTdjHZj
v/GsQ/R8sawOsz59TTrNcU4sC5Oqg5a8t3ngTdDh+JhCE8eYt9iWzFBSa81jYMaS
Zm5AJ4o4RjotYD1AWZ5mY3GHLWz3YrMDallVsbOjdNUdrd/F2Q0TNtZoQb6RAS5T
ktAMOztW/Xz2hV7eVZ9azNTZmxyOC9vJLGL73y1DpQ9mLV3P7UV1+UcGahLdvYBY
9Kc9Ayu3GYGoNP+Y0ri/PsApPErNLPY3ePtUNJMpfteas5v+uFmX7DDb1kFmARLc
6kfoE9+Fp8tvpc53m/ydkx0kA48Py2VLtPltyN5y+MpEb6WpykarS96Ims/N/w9g
BVJ5NCicw88iVRZJdAgNgYZUSEltHpxBkUqNjN+FwSjQ3Ksy5FvSd4GLopVL/+KO
jkBET+cEa5XvlW923oWa55f8KxEhdta1LUa0QSVN/Ennz2VggAMzz0eBTBC05hwt
IQdZmA9YvimfglnqfEoD+Xqz7yhXoDeXHi/BKPI2Tid3bEcUwrqQr+xWmabyTt1x
6vb5eZ97VRG12KPQgV3fGNsanvlg4wlvjLM8bpEQJb4BGhu4iY6mimMlcWENmJ/t
I917sMP2aPhHdwLprCXgibnX/OtgGg/0usRoS5Q6MLzsyyFtVLCMzG5hOkGTNQEU
Hza3563KJ0vPqCfFGQ5ltngNlaHQffn9M5p04K+PkjxucHWehlm1NN1jf9FwPcA4
nrRrxOAfP3dOgZRHYfGIqI/nHXQ15xHKoSe2Dpvg9vVfYdpTlUSP7QtWcQkknSLK
imgToSkPy93lK6m33yN/smi1XjMG32h6oHGru5XycN+KovZ+xEvJjRS62bp6pGZP
F1FvnaFoJZEoaX5yCrH9eT4hu2f7NK9wfOh1a88hygBpzhboXvW/LeiFGXl5sn0A
PUf7VP0SQG/nnldTvLSxtz4fPJVaY9ZV/nw3EUJTfVWxn5umw6uoWL83oVmV5ts5
5LstLKadiGucjS4wukLp4QTjb1CJeyBhIW/dA4V8YXlv25DkiN+IAHZTRpr55O+u
bEyjdI6Hs4hE1HuJUbcBgIjc19JcPTLBTl1MJnB57a8ej2LYk9J5mXjv5HUYNNMa
dIUdOdkwsLrU4td1/FAu/sbB2s2nihBDJebw8uz1toh2tTaEoop7jvH8b6h2BcaW
p1y40flF7YIhz8zQYZXriXMQtLmQnpJXZ2CHlbq8g9oO7tbfWBWpsT1EmqRpeyGC
VfYxWoyNKOpnmQ+gWfRA7VUWtwSV13W9ToE9v3621aqSEZcB8vMPPCEJuSIIuZ4M
thUypC52kx0Wc3pjOz1erd7iBOof8+a8OR3+Jst9RlG5tYMYIeiunigol3XosIVc
6kBUIIWj02aamT/++kFvthYWJy7XghMySmvd5XICOUG1hSAfxgQnDFZZfn+/d+J+
SB8GOlFCiRVYGrQqszAnIXTT5qY59uLtUxkjKzIvulzW5rpKDWbTUe6Owc1Fl5im
OWRLhiJFeYGicqstR3KMocNgghl6tUNNuRIk/Rs1VfjVeqd+kFkR5dpb6hmCGptz
GeoXnT9nwlakvNabjfLI4HV69kTLh3Pg0gmFIaxevDg0JHQIKslxt9WquFHxbcXz
qsorFngNhqcIk4PG/rAhqG0Tko8kGcPOirixboJjG65tk+aYjLbc7uXteNSERIHU
5+7YCLPTJzyyqnEtgtZPFr+Oqe0mEZpQCsJnZDKzsy9CaWkQ6OV9Emr/GX5Gn1j4
b+T8CVKW3OMU/Y2QVhumkTckpffi0q6aEnPbHYc8ybBhwPee6za5/arWFencrGXP
ElnBfKXuCpi6GcMZM6VYNR1ZZbclYzLU2zqbQIaqzKZFIwELIdO4XFqpETDC6ITb
8pfdjQmZ6MAfyvf9WiFQgKVcycUpVPYfjA0T7T5uIilR4hqeUrEuzzHCT6Yuo4gj
jEBH9HGrt3YvDozvRftnr1PZWofNs2W84UtXxaP5gEDVNentD64WEEQ0Ruy2ATiq
1Tcncq1Y8qFBzFOKN2ELcJZwJIaqMdJlLPtjmj7WiPuNUIuBTqvRT0YlhaFTJYMf
lKzM6h5jzcDr6sJKlksaZsE0hRF+KGQ+MOWu4KV2vVJvenKTJoU/W9G+X56MWW2d
UJXg2X64zpA6wk3EFekK36L/cicS4U6UpwB86p/z2d1f8TypPswukKfwItBz6MZp
93ODxu19lePoLUebNtoE4T7sC/Ibeh6L8M8Q7/lWukQ8VP1iyQ1fmUU9vsuNTHcR
2jKIZhfCpUsQnAjNngpobo9mOvTsIbApOH9F0M6Xwmr2P3Ov8+RyWFpdSd0XaFsA
Tw9/p55OnE8Ty+HkrVF7ckmtdOrQMdBI+i312kNSfk8QIhea8YN4M6DTRV7ZQ+/J
YxNA7ertcCu3/uBA0bm+qOsbxXjE9b6uDpn6ll8GACGEVXVOi39sjNU2zQbkuuTc
c8/L/smleRWlQT5cJSeWyZnq5kPk0yJd4ubfhg/QW3iU+3gGIaS8xfp2ec4qO8lh
Eia8tOQJEKZ/7hxlTuthUw948Jd5DmkgpLh9hgbSvWMEHk5lQY2vCHSAey18p735
BNNz5Fu3cQk70kLEybuwZ2fFIZ9XBqMa1snPwyfGZy8bkT/QF7IQTPY+YfzwZQmT
02A2w0vhGdQWYZ+dm7gqNr8wP7XycZbFwn/Upn2F+Pa5ZUjM0Wg8gqvMaB5P1u1E
64zLnSybqkDEU+sE5ZJxkKmlihLhlWXFJME2XVpuUMOZoVP7kH5e0fPlgitQbVZl
3XbBGBE5c2MpCMSXJ1BPgqDld2wip/Kr3yP1teoL4ovcvOlKg5SPCNxX80Jirmh1
JS0BLXKqqse/aHxjAJU4vK1B8x3bP3GWV0ZzmCOp5rYudUxb97jdKXxMmiPBRgsM
YSye1FVr5Xd4JXJ48qmlb5z2Kd0Zagcs7Agq+ug+JpHVik7AK2UEKPFvp7VTfCeB
Zl1WKiH6+bzrjbjoCyuOm82i1jk4VSNLo4qJ1Tlzp7M9zoqifsUP0uIkhtwmBxSP
JMFZVwdhRFe0kAiXiIbchgCmaekNIQcu0in4Pd0EJABpiDcJVvtejLJayi3rY30b
mUUMelXF4Zz92NjR3MruuCIvB/Hh7xOR0u4p2OnK1qa5yEoC30nTugeLKurWfzZ4
Vlw7DxhGmtT8Som62O8ptSjZdf5LwJRNcr6oip2SM+jyJph3lwK6o0iPZtooijUw
NI7d67EI0ZmdUT9/ZqjsQcskOL6uvIBhyGbDXpJMDq8oW0+U8XAupnj5vTFEcSW7
tIXS6UbnkRvx44PMxbXqTsInc/KWvQKFs+qt6q7OCdWLJ1ncc/EatJJFjOM7tKkU
bKfndKpBB1R8HrzD7fBkeeUuR6Kb3N+8CtuejxLYugW6CSa2qGhEAdZ+taSx5+PN
BM0TPzGptj9BO9Vafx0FurHclPGfauFucNL0erZQqlwTIrEGpR21cSzznODT/iQR
7afJouKpf2G+PPPrgWloXiKL4fnBwiu4l1MNdRso9aa7SsjglHYxqEDObCn9NGUG
KWdaePAyx0UE1SBMOzVTazgd6xVE7Inu9Y45xdfw6JPZQy8B3tWz1YH5K4uF/d8o
nROpMD8vt6hb0NoKKmSC9fSYsW249VnpVH2sNCSNccVzImPoTZlqL85zyVQbO18j
mciMsaKtkPalXpu9Bz7VRVWN02k3ahLXgLayDJfHIfTKzwPR+7+4IBxjQ1F/XwOL
CSfOe3f0MOHd8D88kjWNXJkWbdCkvfJSmrlHiRCiC2/PifKaMvh5dKApyuBTn7EB
N1T3pWMqx4cBwxeSofRICsr9XHeq4Aeb5TDi5z9C5z7VlCAgwptszVQ+Vyu3JfWM
RPErICuzCC15cCatqdkxHI8hzbHGYfY/NqfjPEGhvVrzn6swPjKThG//XLdxDHNM
bPzeJLF6Qg9EAU2y3I4av3+F6K8jW/WQBSbEziTUZdfoaviPpaQXAbaLXaj950/v
yZlyy+TvqZxgwxwwmd7HPyxiinXHw0vmozg82lzqZJ0RnO4sAsLJeOzbqf9SXgNx
1souOS3mqj/Qgd55QP3glX78QFt2fOts8MMbtOdfaZwMWe2bwqtlBwBH2LZiZytK
H+IvGUJj6pShMqK4w0LlFIuJJ8LHIVnDZfNRCeg6LWF/9qZzopf3AuAfYCx77Vte
tepvlNFkjlh5bJELWm9TTYKWIaLRnM58T7jY9fIoQZS29qwEAfURWiQy3vYRMH54
QpCUtw8IqXpIqPXIP16tc/09z39CpX26wJCCcEI3Z5capA0nfPgMizo3nJ5mGchG
9wSY7uIqYjmoDacMFL9CKvgKYPlILKCQ7owmjBfuIw97bfreBkMy2YHUlwSAOVV0
EOpeuc62zUncFDhRxbsPx/2+tpIRscYiPIPYRCDPxTKLbAaO7nj4qeYFpsEgr215
Wkrn5aRzgGKxSCZclD4CyxNPPxQsUtQBi85w/pYID0y4o+bPR7J8s8Ck3/6NBw6W
5AxYE/3jVrDgyO+VzwiqO52M1vPLBH0tafa+RxrooJ4m426SSoYVhHBE9dLzUTqz
sGHIhdkanHUIohI5NEnxKjJIXBHPumZmT1FGFNKr5R0J1ZPIz4gbXu/65i4wXGcz
o42IufEq1jI7TYYOk0pDQefCEpY7yk4Y8Go/fRXPC43G5MW2g+8Bak16Lt8QcpjB
r3lw5EVd6KdR6Kv75yVppxpad2v/PwMUDaOQ2z7ESsVqeC7uYmCGDh8T1jIOgo1e
swfEhpHzUTkeTAJTk8CfyfjBtBI8NkbA6ML4mTHEe+Yrg4eyKPk4NCJNaD7ni3Z1
1rufmojFoPdqG/G5sZajJ3M2YSEsImqx/AZ8lYUJ5B9hzf6igIyApgFuY7hMs9pH
g/8NS3z+cTwt9v5m7BdHnI+9T+lzNTAdw7CxxCu/tAIS9zZJnlI/K5uf3ss8pjix
vpsbe9YOe/JZatjQd2f1PlPrzRh+OQXljSH47I4qzCbrRtx9yJl7D7wROMuOVZUR
QRu3J7or8CoAzl+sr+B2agvml5g0y85eVvuBpkRE/jfRP08MwmqtuBiVzeelpvuS
RC/TR+nylgzhyrFURENw/zyiUt/pJHcGvnqpSxJ322KMDI9pz+x1ZGVkv9zllaAy
welKyYNn3yrmnKDpBh91MmigmqYlyoG2uanJpmGVLkwWncJI3Qrv9iGBWtb9t9z5
jfpX+O2ibeFNUbEC/PKykwhKioKGOnQo1ySRoDrvC8B5HUGCM4ND2kd0/jxlyxy0
G3lgcoxXll4QOFakjrkPNdGT1dwp3/8+B/jFovTogNZM8UkN4bVfpCUUWqNs8Xty
Ls1dCohP9JPRIkgdQjcgYhYxcfz2Le+1facZ/YSz7Y+qzIkGyu6w+9OdjvahV16h
PSAOsqRcV2CeBUuBhJvzmLw69neSfdy57XImbPlVYCUG9m1DoceMl/G0AOpH9cTO
sbjY6b3FFbC5svPB2xRsxJZ3sDC9BB9ERz9uEWnT9uT7bQbubiqJ2wwB44ofYBYC
NBuMKqcJnzOnIIcLrpkui7HZyWvZxF8GHGfzM0FPfoU00sSsKUJXZmGv+2j67X6T
kA6+5FbY2gImFxkLTamVosJMRqcxBVpClt1E1TmQwlYAhBT4+2uRZeEX/Yj9f1V/
GQWE8m7HFW+qNmu+6SHGMtBSoV8VYBNcm4lD1pAO+AVaTo/222TktoMtRBYdUIFw
50u/La6EdBcR3QbLjFX6Tjfdv85/dXs4PfkrsHvsLaZfbhZ3neEd4miPxAK21WCL
cPlAt21ECQ5UnFbs4uXy0mJrtqLc+bWOF+9tebuH2WvMuAnanXaeM+BV1h4KJp5o
K+Gq93Q7+u8Q21UmU3aSNoWr9lUfMnQUcxJFFk8ngWUDr8+0+gl8x5a4UDtq42bO
SyHEOrW2w0Cg0bQW7vovpBrJBO8KEpMA+OG+ChsTx2k15cWCqZFRnNaxS5wqQrnY
iYsKCDH7OzgcWZftM5aQ/buPXr6gr4W6fpoVDTe9M97txu47PkI6X1gsBrHmo2uK
ovFLWd588YEo7lYPzVtFCt/kx7AYLu7rxaOywAyPzECwODo2N4Dv+H6BNinldpzw
plY8N9o3rQ0L0VAeRKkVhuwSU2rL+Ic8lu4PdsL9vshOmdoEE2pzr0jjbjm/fzw2
6rXmkibSBRUHU8Otxw5WzSKJa3nbyEGVplHxRXwm+gAZ5D3OGvzXXVele9GiQs93
+yUrGnEzfhyIUzuvBr0MrDFSv4fN5kRN0HalEgnUAOjwB6VwPOe4yxVOcx8v7dbS
Dc21urPTvOyFmnrt4HIiog/yJThmFNe4XAwvip6GR27tvL0GBqTluUC0Q45LcZ19
NXIIMG5V9WbDMwkgn5IPL5gOuQtIFRnvL6HlFaR/HAki5REYO54dar37RVse8E8N
uR9OPUoRkRfDrBbqBQ+mplN4A/SGCPzXL1tmF+BXzHF/OtwFsaFFWQgL9vgttchB
ff2eNQ+7YKd5WQ7AO4WiDRHc7uUZSImd1E1eYJGqs1XGJdWDmZyemp7mR9JMFOVf
jU/Ttfcq0hMmhSTS/+r/sHaQsgaS+h6fBSi09yep5f/bDavt2MBTeLwhGwGFU1xI
LFIDs9Ry4xgaJiWRHZeIvqDsOhd/SJwqbOKtTI6+vQhDoExqXtb4FBsTSy/w5EeB
AZ09XvEfYf1TEu9va8w4ccb7ewQ7iw7LOQ7ZPCqQ5VcLxXDkt5k+Q3M6D6+Rd3FU
YaBqWwBsUwLuXAWXhoYm3D50hZjJjxwfwVDA6eLvv3IxEY0Sv+aGp3oezqyEG8aW
6L21W4At7zF2lgarfjiXIB9JXtFzdubfTVU6rGOlKYiwKxnsJ4ehECn6LuPcRCwr
jP0h4JR3ldGTusSCgVgDgtHEJnVRYzACOCZGStUAK+bMvDMHyva9lAm/x7CuQ6y/
P4OY9GmAPWb0e+yMZklCYTO4RWXcbshTv+xIyzOFmuExgpug5S09mxe65Yv2eCSO
mBiyjf/q4A36IuAwe6b/WqO4qCV/tfJEHY6zCjSZOrbduCYGY7mLQRWhzo3Xxawk
JU8JDO1hmWCI8aJwDPEEw3jp5MKVr7AfCzTbIecbOWBtadlSDxnFcYtgKWO3Dpl2
Yy1PjW7Uv0s2+9HL4NfnSvmFLOr+ToMga43KGGvtJPEtGW4M5wzLqciksdr2qUuW
5zcZnvAfO4GoRON/oGu7mWxSSpOL4k1a0so/FqXcojTOJXqcahwtuln5voRXZ5Ru
4veDA/7x4RSQIxAiFdC0hce73XSaA2dExxk2EtzthwKHnE/PdgIgJYZccSD9Vbyq
udGVJ2Oftxhz1/qY2nbN/rQAsuMbyx+ayWLpuKFdGSWaEPrbj/Izeh4WmhTy32uL
PxVRj2lVYcXN5PXY4c/lDgBy3leN0DLc9VqN9HALLLyAvUlOUP60lynV672fxGf/
MflvYzOdOp78M3pOsuW6z2vOTzFvBRbFF/868w+OVm4AIYyFHsfIiny+Vpk6E4qa
qNy4GmDK9qIo2yrReNdWDCIGqzCLkR0ZL3o8TnyJHvlikGqVpqeG4+/eQFBXAsXQ
SLQVVdidV36IDBGwY16zxGNalT1VXj/BF8vdGG3/7HMscBBee9mqyeRI8tbi/Uia
dmkeCzAJLgl34UYYgkePv9SaHbrSl4/PHzmRpYOV+K3GUlGMY3KYlZ6qgeQLguW3
4h5tnw4U3LVFcMdf0R20whxHO9BpVZvhMEUqQK5rDwepVyf4pbQuzYNp8mjVyLPW
1DJ3N90E5LOdeyrqCfdW5gRpmyxbXcMoz/1WTnKzPjRKwuvzjk0J+faOj8Xaj20h
+g+yAu2xYdFCCEtTkoYM6FXVigzY1GAacyw/XPku6MTI5ANmh2ZNsF408KQhd1Go
rWuscFCU5J55j+BkoNzg73uZzp0IkoPBBmis3Wt0wx76oHKkIxlqCsrqpgDQDmES
iAT+haWFa3p6bzHJJ09BewQQY4FSFYdjVVCttqULPuIJxCm2IRNSKpm6vNUQ6Nl6
vemqfwbfbgkpopxKD+ZR7n4PMOQI+ewu7D5euNF4DmzATPu/3NgF2EdnU1xJ4cCx
t6ayAXWFQmNMHKuhRhCm/LL27N5WGIxS1JMzOghqFSx6I1ZP6NGp0J7DUfjeEuTk
Sv8T5kC3zU5fbap1Cb89+TgbcVhyDmRZ22yw+IIjOkn+TODtckBY9TJIrZjJXBed
zXFXgg8+Y1aCYSLWKmQAqmCyP/ofPCqU/jbm5zBwxWy10CKLW26Cv98YNPZFaoAK
Hz2vzWK+NUpmiFAdld9nVA7yhpzNHnLDqVTPuEnGtFYhC4NXloX04sPKF0Td3rLd
Kw3o8ThqIsB0kFny3qLoRbvl5khowkFWrAZdKf1Uq7GYeMhKspW8jiikGlu/H+1u
SsRHVnKvpOkR0FHQ5Y7q243OfBgzCRz+Ip9NgOLPAQ+Ra6Q+4KEdE3mb4oSN2eF8
wa1W3c+03rV3y34JAwDVKcHij0LRosOUem5O55EbHmms3e1+AMddIf+WqLdVCf1l
hC+yqtUgNK9rWwFzn/ZEBs2O+2zaor43u6FQOtXzfcZ5M03S5DB3ERYGdKDdHOME
UjjAiKoSSbnPEjoZC+eskQ8rCu/lqpGPOE3LMFD3wK/JxfbRwVnBwSFJG+SiU0hH
r+Yexirnv/ZoFZoDKGpQiW9B7z3YFDylSdlVbwy5wUABJciNAOoHplkhIJ17OjMi
KpueDUT6rXWz17RRKGsnOO3wT7MyjLdxYZcVNHuGSQJSnLWUkiZmdMnfKRE4qiyD
bWlHSNz1VFXLBKnAX29zWYHw8ewPobh7nII8ZMc2NIB47gW01gbz8qlGkdWxCZO9
sD/tqxcc2z0TUwUwgtNzLdeW5DAFQJoDumhWMsVQvX0UIGsmEWzXgWSQKpCKru6s
Db6sLwjvQXJBz7/iuTlIHSWURSiigbBL/MKfAbT+vYSskgChAXlgfcht89McKvw1
3aCQZGt70vAkw60jt9YW+ueCdcVDoFcaz+bZCTqh977PZnCpPFOfY7u2+SBmDAkk
7ni1Jm4lr+6AcaTa/q8LgDcLWTqHCpROi/60PyM4gUYstL9ImIWm3+Zp1GJROFHC
hmZj+StOrZHrf++2Dzd4Xh2bNDOCIwHwbsxh9HvdWF+7UR3Mz/qOmmLyEwb48qc9
clPeIi+kBCCiovuYj4NhLXfgudUNY18g7l0waVcxPYSJsU0rUGsCivJ82MplExGj
A5DrsZka2HMFHJz+9sXAenVPGZ5GKc5GKL1GPekpNAsP34NMcV31Axmk6FFt4CUg
V1Xgrvqi4mxXz1W7Xi/9BN2+2EXQp3le0vWRrqvrpIPfOgETjt/RKaimwYmcKqN7
GNAq0Sc51as+6V8hFyRalulMPU6vQfTmsxFvufoWhU8zu8gGMdWX2UFzKGBeKBs4
U0CgLxzO+uL/cjXoqiC70HKuWZuLUJ7XksZRkN5omMfd1tHS+NwjxM8nT/bwLgo0
rqrZsxF58+h4ToBrO5zmWCkrBniFwExVVvZkb4tjZOK0QhiyErqOUiECpaa4fMD0
/9kf2mmB0a2yMUswd/DQwxAsyi3x9IikgrOfeogKGnfw7KnVENMMUmEjWN/DT2p1
CFF3zUtVUycO8hbeVHWlqCi4DmmCC46wBeqsE9aSfV0ShFlv0NXXgODC/z/XzYzc
SyiLxV3rgaxFoyZv+3yqh9ttIPMhGYjCqtkJ+k7Aq4/2jw4Zb9BBA9bcTM+uzOLd
4CcjmTUQeU4/3fp9vTE3xwmtOcUkpo48kh00Me8L6U/LKTQVPpCV6VzF19JSFYU+
or013F3K0/mMsMazQAjgkIvKMBlkKI9XIwfDq7ApRO8H7qUVVmFprba5p1PxpsmO
PRaOjK6LQauNHU3E9GJitEf2zTFdMGtMGJ9Sop8NeYg0f+yEG2+DEs67ZgJ4kyJg
KXU1LdMyOOjGq9J898clOfVPeKaKduQWG/ZlrZlBHWn7vPse8OQu9oZgoibSrZbP
EfLbgiU/iAFhC5Dtm3a9aOVTpPQZnoTnAJnpdmCGZeA16LWbaG+4twoFt9WHpcBM
nyOdsh89XAAXWu3/aWbct5969C11HJZej67wtdg7FO5W0cR2H0itNVenF18oDE9T
G9pkTaAsb49gto5j1bOTv83UEs31ygymx6am1N9aXxxusjADq7K0q/+l+3BAvM8B
fJnJpAME/sc8KGbHv2yjEIExlYKlI8mUQrA9VEsC+xdwGprs65yiImPadxb3V3Jl
zuXYT72h+22Dp9I63lxSNHXibP+ldL7kullIu6OthrN+wcDrBHCkYtHOU4jLbfuZ
Ey6cRIkfvwTLijlYjfx7DymcPScknr9otQYjkaJPVhZYuvEzFedW88lTpDFKe5lT
xsJRgEr181mpammkXe6b8UDKKxytvk2/Ry3bEZZSxSJ0Yebe51JHHHtjua9gkt3Q
TZQCZA7Q7LJB/xxkhQwyCEzFLxWv/4nevF++4AkhcKWoyk42/OfNGZnATXoftWDN
UiPjvF0RhxrJDPjp5bv1mM6NJ7cEZxDgf7Uc8y7+KWnCmwhSmPQWq6KLtDB323WK
ULL++WCzV7W/ZDmjggmweD3DItAODVBMSuHokYakSBSyzISJicyGtn+3hFzZ3KHn
uOrPBZYwUDMVMGEWzx3yOc44+RACbyS6wyIupAn4yDOJt6KSJtbRrElVcWhjVh3g
mzTApQG5bi8J709Hwsh1zBHkWgEbkBYSStjRF+NFIlKWo6tmmZJB7oiSH8sxB4+1
nc72JcOxjWyq7Se+9q2cjkJ4ge31OqCRVBpyOlXpcT+erVt6ZdbPm159mwOOTSH1
+zLJ2BcEit1MRaAuIdjg8BaOE/Ohsm8Y8f/ZJcCgmJiYdOkzyXHba4CLmDVOfml/
nHspMkvnRnQDH34aQ76z1NDxXTUwNmNK1ppl2PAz+8L03D7JCTeuhYTc8ErFmd8w
HEmXTB899lxFXXdxoXxnnP4COCf2kUos5oPRMYbafZIp9c71yMhjsqCSgd0gi1P3
NRGfA5GHUUwWOsuSR6R/GuHmxBkNyBz/A/qOKAD8luj0XTjU/Ku1LUTgqMP3zvBQ
B9LJIUdOyj0eO3nEEpYJ57NLjiLBytGKIYZ7N7YPovvMYoAOeNtjvhLQR7sj/np5
UV0YLphjDXobmQH+V3Hy5Rxu9A5VFToIXq/pYIZiHu4W2NGuLCrBkS+NJGlfwlwn
0zn1fQSIimI+3zMYNcpT6aFP8uPYjQkKkUiSmIzMeDcJdUwagUvgmwrKUnLOQsb9
5wT7jgBAh/BhW3qUivyoar0wgry0f1S3GqsAwQDd5TfBAvE0wb2jKlhDHjL6DWHb
hEUvV2Fy0vIyG6hCrcUUtA0sci7rwLuJ8GtHqb81FHJnE4VzkQOhxD5ml4gg/ZjF
PVV82L3sdsqgX54XIzuqC9TO04jsAIBY6vWz+tIuk8TSJV4GOkgOAsMGqi4vkElB
JkCMpqEmjc4UqTIg7oNVLMp+J8O8KTtTirRHwUxCpt0QEvKTSlSbWPIRAT/x2TyX
24Zm/vJsXLwrPsDCa/fC7Qpr4flddzN3fmnHvPmwJ+qar6vw4M0BOz79yXBDs/M3
TKl7N7YZvTV/GuTL/0vS8nErQBJ5EKtqBBQu5Xofa75za8+7YBaC6Mq94Bd0pCcf
++jqbFcnc01iHL+yACUHfe8dGWrYIm4r4X+8m/8LRKK6DhdIZDb2BfBed1UUEFbA
WsZqwajAuAZ+Il1GkkE/zjoOMzOEbvL6gaFqfJA+AMAcxA6ErmZ4hhZjqhqtguHC
kwC7OF1Kv3rH3gYSD6grIC1wgLnwhZYZ/Q7OyQs8dZxtxeJstELsfyJAFTgo7SYu
XtEphy2v7dw+gzvv3BUUDAiNLlOhY/8YSbzy1eREE/wwmCs6pXxsdl87sXyLR46G
X2kbfi3paFoGkArN80r79zxyYQHw9FjtaN2SreN9Qe6vty5ypn0fvBQEpSQp6FE4
Mt5tLzW9sEI+LVWBZsV6Swk4rjFIs2mgTXrIgKqujJyfbLIBrt/kFz6iNL3q5GmY
0AoYNDlNl5Dx8CR1PNoePdYpQg+TpKx7eem6cKpKbUSws2UzTfwCvSbYb09FO6Ve
2/WMFDgSWQ36+CWqw0s57XobUjdqr3SqM4RU+1ZVlIHnKkU5f8dV3FWQbxsVx/RD
lcCiX98wRQ9a2JcggN5n5E1QX+got5mkrlk8qaTfjMfSbfznYHyXrZ2X48foWyei
dVd+VwCSZH2970eD4bvatBaI/4N1Tdc885mHo2xItNAsVQT7TnhKKOZkp5a67Qx3
gqIpOnu94iN6FZvzpmmq8Si4WL5m3hIiTcvVRl56bx8qgVGIN/LjhEfq5FAsogZZ
w3fqq1YunzChc53gSCCuxCcAXvDrXrTc51e5Od3cCIN4YTYuBPAKcKNV5ATwnjKa
C3seU6or9sc7/fbL0HsmnRwkZc0lVNMFZMIMSnq8YaVFm//w0hLuB1rlVDIhtUHf
w8x68Y8vFnFt4N9c77pR8b7F5LROcfVg46coGZkQGjUbiFTvOzA9r+6bzD8t8q8g
XRK/b4/NgdNR1QD30/9y+1hOZhSLBs09TPIjA0s7IaYQQD+V0gX/uYu0HcyBr4YW
+rGyedy4dAxHdH3OpwH4NgxzU7ixYIDJl9tS3MbExfMqBbcwedosE1tPlqu0gn5W
mhvf/wszB48am1TPiRM2TylXlRKsY5eQIH+xIKJyFmEPJGkAM/lkFpdi1BgaccXJ
x0lXiRiijRoQVy1/aru/cb3SwtbUgE6Zpfq+3eV0jBc7Oi/jyiyr08ZbyEC+fJUx
Fj90HwiNgSHy/LZEUo6rfY35KO/d8hq3dkDrO79DMwd576BMcXSTO0YyMdLHaGhT
FNe5zumly0muUB4+CrfsMsgU43GBR6KxKY8N75QJbbYdSXMNSIarZZY5htLZluNJ
1dEbTPObu3II9iO6sCpw6N9V17djXRnHmCAt3TA04w+J8V6a83OoINWVmf1QswXg
p+t7b6APc5SO5e8bY9rv94L2dh5/kU2rLNlg/w/h5nBgl2FWks/t5dpBOHZsV+GE
GZqtPvTuPeALWgXtaeV3Ofgsj5v4QZVejOR8tUugkIGgR31yRAeeSQKsfOsGBkHB
XfS7fN9/JQ4nlt1BNgpiWckeeucUrSgJiWMWNSxYdVzpYAAVP5FKZT4XNiRukKgh
Gn98KaFhu9VOw+IrAGaEG9o6SXR6opC7nAqT69qFDRRWwWbp5dCTk7BUf7cpA8H+
DoKR5rbFXzNP3jfvsx5iEKrN2p5ATSyGhJz75EMYW/nRcyyCGO7s44nJ0XFOSQ6z
6CVF2eNwe99oPPFn6iUwkfmWfKsGL3j0T51HxV/MEYiHHiwhlCWPmNLspjwtIitk
kXys32R4wN+bPx99gg9l6tF2TtEGEMObz1VCdf5h/EDZuBRyhKXH9OqrJy3pX47a
sN3N/RNVnPANqgjEYT7Zza1zhzxnd2C+/GGaueuXI5jeHSaJjuTZ/1bPKpJ+C24v
0iAbo5jkT1VIryOqwxFmz3h9Bkb2cI1EoLWfN0UjTCGM4hhd6how7PK+7sYx2Xzu
Gf02gkfqJObPrCuM5M6N50f2yoKwWGs8GMwTevWMdsWb7arkbztEQ6t3PGQTPHtm
CX5D+5atQga3jz9k4+wmbVqmDGxEGZChKx4PMgJRfE+oJeJSmKi47N7yQ2KQS/AW
NHnr2DN1h9XCqFq9DF97A5vePO1ru8wmQSu4ZK+rO7Ce8iGoohAdsz2OBNv+NDzO
KsXLCgZeupOJ8nbxDC8vey/SITKRdAXOvLTJN4XlCYfctdUsYXelXdPdNNV8XJX9
N9AzmFHsMrosFCINwH7Ed6mfBDrS6JC0xTLm91diqR4HUHJwUMi1/qqeO1nYQhx0
x9UrUeVrnlLyJ+hoZYd1EDSIGJKHuE0s4vlt2R5IhY4wFkUv7r8M9FsBxRJcQvje
JTY9tPitzwDfiEsc101LYl9GPqUGeXa3HW90Kgz0iLs0UJXm7ZUYIzFUw44KzTwi
RgJITcz5gqGBpDEhKnN7LhY+ULvhNweiaIwBtchV4MJv2QxQyeVpnEXSb6iQ5ZFF
eibvfXfMeiKysNEqjRLzgSPFZC9iHUSsZeGpCNg+Y6IoRqVBu+GKcuaAnbL5Ijtl
BeDd+A6N8QGjBhJmVrE4fKpau5UOaZWu+wWSNkO08wGdxQ7ctsfqFR5klHaLzFEx
HtP1+03dc/0AJKxXz5FbEXvKGgDcdP90Q07KLlipmTDA+6aUHWkAjfwe5eaE8rgT
Cu43GgrKlKwWv4oIcnlJypMQjMw8Md4R2vWvzQd58yjkqnI+P1PVHHh1MxIZxR0F
BgurQhrn7jcUpItwj6N6OwuAUBi6ecM/kR5bczfgXcK9/PeLgnXif2dAJzSF+ccP
yRSY5zPWarmbUsv2s3YK9zmqfB5EwZIwf8HcO5PiwHMAKWMyKe1M8DqaW6+uqIyR
74YfKcb0uVxdSkf+HNPamI/pTcMOPstwVzFG7AaoX1vl7vt976z4kt/wWubRnakl
Y63E5lWmch/4Aea/+Wd1Bcb4TU0m1fIP5T6rOSFqIZQGDV59Bl4sWD21hCf6cr3A
eLN8m4divZRo16bLdt7qdTvQ1z+gMotWqwfA+uqmF/lHZ5yymA39hPCJC2BRGB0A
JKCFlpkJ7c2SBRmApsUnWRyEKZo9/bhk8XxjX+bZHfByupdOxwAwpzYzk28X2hs/
c4vrn7tpMFAv0MYIBgkUbT5W3YaEgk/s1JGLYIH9og708NGaENtYW+apD8M+1lW3
AVADxVe9DlqMDjPfM0bMM7DOqEwoCaooiHmaAsb1EfMkAnwZFANNBg56C3MWqmRM
y4Lps2LERZ9Zzk+hDvFmrZ7vQxg7hkbiGKh6rHtNy7oqgo9wfJNT1lXtlOvpDb7R
8MSjrhoAnp8IvJTA6vGHab+NNEnxEBL5H81kt/f6vK4xTdxe/QwLO8HNYMQua31E
ENCGu9hbLEcWtke58uAWhmsESivvyC7eUDeZnrn+J2ESSMj+PcJn7YTefZK3WKun
c3pvIUvUrRJHCfkNu4zMzgYQdDh3SbVBAGOHGi+g67GB9NDV/jdfo2pIvD/Sysme
Iz08eZuTj4s7ezQt/HEDImyiIPjD9GuVjxqYW7ojmmbvoRhmkZ2Qr6W7dgy49z7k
pTgHj0DHdnU8vbr9x8zQyGPHVp783eBsquOnET78Zelo5QI8WJH2bWlmqdOkbBLK
HsxFQRkOKk60IN1SB+9AE1updHHbxdiVeU+RVqZNjA+O6vpnj0LyPCMGanAW0aeC
R/TvrJOKKdp5fxrbNVnER0BGEiwf4uJxmNurfQZ9I6N2tx3CjjrSmRpeUuHvgb7n
vOOh9NHDRoG9ZCnE6Ycdq6cAfYBFxDboplYw0fBHWHtxROh2SFJm8x0G6Ux+qn8B
m8/Cg82WtuN1YcteFcl1lETjB2EPn7GJPpTwrRSpxR9R8aZvcyb8kZ4WRhvHx2g6
7IQ+0XBrzdkpX8RcD5PAHE9DCGVgHtJfUdNqNpnyzbPSJbObgbvj0XJmPWiHSGr9
LLg+e8bksQx/GHtOVJUMz9sgGzDeoiz9NMpaYQhgK4yHjl9EEr3Yv6bFZjKQ5WrH
EZzMBefQBLejQkktX1cgpb9NEKqaiU1hh9YDT1nj8MLhYQ/e0I1VaI9QWtWJmA9D
y4/ZEND5wB3UMCGn3+zSrMl7PTx1h+9EkgiQj6kGBvxVnYASDwGOGL/pdWmQQmM0
p0KV8Y6dzJjaulvtPrVDAWoyIqrDGNl8VKCq3jaBCi32kbxlBgh9oB2NQy1D2iRX
0lGi4K/2ebNYZdki5myRfe+vhYZI0OnC7ZKSCtV3jj/3r+iir2vhdOt5RO715l2L
du3CaxA3erzB6vwqQdFJrCE0dcqxgOY8roLhnAtyWWzMLBGaUyREcGP7L7u/s2yW
dd6j7r/KtKmfj+zaWO7FbCr9KAd6CghaT2kBDks0Hw06zFVRH1IuucobtFdjlRYQ
SBIt9gXpF18Bph5cVLJRnguLQ+LC+0AVBe60IvsEX4tHNoMOTFiduqrqFCvzMUJM
hhK4IGGzjDi0WyzXlizY0iBuKMRua4T1AUzO3LIh2AXDS8I/d07yyfTfKYfL5Ipu
jP23UnBO4hh9RngjxiQdqgIuo1c1fF6l5+d51kFUHfcVSCsvZUpOSFRkZkKgHdpZ
c6TOp1pJVtAV7YHeiOGuY1JMVgs0ue6FJ/fNTX/iRxU2Lciqxk76cRqbxLiSzRhf
ylT194117lu2X47/7YrxhuWexn3xZk5W2NKuwhmjvrxDFBZjSzJf5a8fPsms8127
nXlCl4g78I2CVtDelrqO6A0Npl4Du64GreFeE2kDdJ01N2ofgVKzrPO+oC8piEs1
LzuDmt5uMMrZ4MfJp2DYvTRV9Knl33F4OFgzqpTeLZ7jA8vjb6/f3H1CoWbj8YQU
zjSJyO6yU0BFPXuN9g5BO6FZzS2lczw18GDIOxXWgQAe2qIlSjWICvd7ADT3/uM8
fI0O5dzOHTphgZOS9oB8KT3RDCyKRyq+xzNLtC/iQZ6D9/p2K6yC5OoeDI48WoP3
G1A2VYH7gBMDhawMrPY7ttLSeZln0NOEIIaSQv2Xi8LfOpg3WUbRQoP/sR6x+Zcz
eGunoeUdroUlVTK8OGJHZbxjjXZjw9BIuATb7H7uTXF6nbDd42fyn7RWA8t2GeYw
S2gPzuUC6HBoic0ySRRUOm8E67igMwN8pylZjtLkvcMiDbjxi99AFgBUU6m5AdTZ
yJbxm49e/nwlP7k3HP/V64SQocN+U9bdmLUl2ZEXFQo7Jp+5Esp33gwHekSNrIKP
oxEtTKRZ/lnSU8bP+bO87DkKxT3mPK5EmfPU94+WT7gjbbHbfLth+2cUey4s9lFW
jisnLCVQAmDVvxN99jcRJHOWI0Uhf110+CGP/0xJsWwH3JTE3HbUfEEw1Bg2LRfC
ALx6cKDIlPS5vbRK0ap/npsgAhlEuJcMQCrLae/F5RMZulN10ZQCH7gqwqZIsBwA
Xc9TQjnhDRoUSblze2zv7WQdrcZ49ERVVeGN43zzqC0jhOwHU/mdFDXFEAkMtp+y
1h+wbr/qOZQ5Hnav+w/hDizpevNiedvkOLgoE6NP7skcTeqX8A8Jix/+8it2C0CM
4YvMv/FnXSFQ9S9zWKcwDfdJ0aE15lNhLAurGpqbNMLAtvPjsMvze7au8+tW/1p/
7/lzBzyfFzGl/8ipaOI19p1qWfxH3s6iGu6oJuWrYnS4Ak0ZgOG7fIcv3JWA7Yq3
21uBGsBi5OXgWrl6S1Kk2r/J0WBp70qXB0KbTzU9xVyJOd7Qd3XKZySNu/QdLrzH
G8S9/BiYr4OqGoYwAgdEdRW+JyjO5urxeX1L5sUVhmfqzo6STgDz4QztXZdTGhfS
9t0l1FQ5iKv8KYd+aGicDzXfZdaZOXbc1kvrw+L0kMspHhl07eUViBsTF9zdBC6j
JirabUr85Sd0XrbodXVTQLOtAeqqj6q91q5DdOWhYQXem288OBIo9oAWpWsf+KJP
k/X1iMf9dEtniX/uwjAfAt5iw5WQryAA84tVFesDRhBJP5mxDUwdczHFMpWUR+t1
U/0n6T1QUJXilTD6gGo7nAlVMnJrf3Ct+1KJpq52UATadYq2JtYJqp7Clb+a1MKf
9mi3gelFAlP/X2rkzpAzt2GFZQu/U86hghh6hqMPUaswqGGWO5/Ln7b8gE+xfJUK
cjNdl60jI79hpgQyk4F6Trq6+1uvNBhm1/vPGCybJKVbKy8Ud/1EhRz3SUemXJMi
hIJ1D8l/iP1NHOXzw2rTzpVCHqvzM4YZyqXdeF4QWson5gndl02yNUtiqFjCFPIg
XH8fJ5iB30feEkc3kgslBSMf8iYm01Fa3BdVODGE1jnvIaxGP1aPFj2IVreOFsE6
mwcxbP5WwRESI18m5ZcWZoaw1md4ZN6J62H+bKE87UxhO6Yvm856TbvTuUc9zdSz
mHte4MJkPEDhnqXqLWEc+x0coGiP/ciSEC4hdR0Bom5RxITfXaPpliobPg79qm9/
D+w60P1k27lfVNUpc+FQDjPymGPXMqFrM3I1bwyGPTvCEURUD2cyQOp79VrTuEY3
rZTFYQTlWSzFU72Wi3WOELg/QGFVsl3VjFW6HH35Cr8bQTSTky2BgTFUVlj0Qsqx
pLUeU6NrHMNE/menPOMdVsbYwVkJAMUQnS8i73wVcbJ4hlmAgnqkIW1MjpCPAbde
ZRZujloQ3BDv1ZmYWc1pwL5FLK7UO8qyRc2YZ/rLU6HsWBIa3v+EC7HE2jKOXa8x
6lhLRdbsLnvkZWJNfqkr3XLanC/uv0wO4DVSMxOEfKjCQEfeYi11nYadkqHORsQs
jUmx2J4INoG5cEeDUJsa3Zd2lhMjSV7GEdZivj6BD8mG0zx8kDqAUfsatuiGOsaB
o1O6zP/q4EmEDhxJbl65wNBUQ420BQUrdBfkG1J46EotHCProMyvIBl6jqO0EsAd
vt2bIRVhD4Q7LBv4qJSsULz6sgRJ3Mk4Vq6fISM8gv0Aj7swxgQNZI65jmdZDmt9
gUmcxouL7/6yclyK1Dy3ZLXezQQV9wxKEfyPUroCOxjVOOa4xCr2TFNWC/rxI6e7
K5XAznADR+hTDeVm5MG8GJEuBttuACgGBh3lMvBOO4qb0WW9XM8QfakWbIJEBr71
RbFrv2ss9r8t5dk36+HRNnRncpffOusR9VA1re1mlAlGq54cLQCpxOdnp7/BG3bo
rBtO6EnhIR072CWLRu25J0s2IK72IFUVwCmNeiNV7CDkzJR26jawLyh3aZm6bKTc
0OKDHZ5W1b502yEj9pUTLRAGMqVB4G0sxx/2NsdtBbEvy9pDie0s90bM4F0Iz5sG
OZFCqUDtantIBSo0KPJDqqFsPAX5uI76IE8GvmH/4DR938dd8XCgrJc2dHgoz8x0
Zp8fFfv30Fe/Gpx0tnc1ObAUqLgyk2i6X9NZ+rvbjVPCMs5NhcrK6n/Bg+obCUAF
SjD3qaQB8NxDQ/GnXhVdAsnVevmfzf3jl7jYVY4yLJv8kT2yelkl0JxEappg1zjB
3oOtKKpDTLUO9J+XGgJ2DzTaysOob0VBI3UlePteQUrQTrpsjtIrEFgg+14fL9x2
pZS7HUsSYKEI/cURj/cN1Vm/KWRJfNXEXcso7A5KTOVYfT1kZXEZtqQdwEOHJ794
nj1M3LLvSbazl9KZGxvTg0AfyimXo2eCFv38ThP5gnyzFf6FGgNd+UgqH8xzYCow
QAFzqUbfi+qaW+yQjesp7CvUUzoa/WHVQxTrJSAf5xfFFPjOnCFrJcoqCM31ohrP
jjh1RNor6mpSbXH5Trbv/JVfdo694eoR06OMFRckwZfajPFEpxWCggrICHimYjrZ
RNGdNh3URSxM0GL0Hgba7VOh7PL1TOevE7WOMmiqelNtg1O1YZb0DMkHmqyOGTtd
z5Ni1fUfPGnTKxGA8nISy7BkmErqzktM/UAtiOsibqVhYQOW07gpMXotSDjmUlt5
5Tjm1tW0F/AHd4Bn2nuN+Ya5tkSKGiCApQFTXboTAjHQqCXC153xrFdbPywOtwa1
4xZEwhVcfQVcDlJcZHnhkNsi9wfu+2Xx5Xi8urjRYm4ZkbqO0MK0QUeSsSliOIdW
l+LZINp8Md38Z7I9CkcKSTz+1Vx/kRqVQbZ5sPvLowE0GOxNcBznoZoXJ0FnNTPO
jARdsYTBgN6CM0exCduczWjVRIwD6AITwE3vC+OntcljlN04FeVk1cqq22vgfgRV
xz0ICYM8CjI0JG/l4nR1bC24s2EzuNlylyy325oEQXMWJ6uiqSbh25RqV7/Tsbeo
5x7qrS4HMmPNYROTHLJ4ivTq58HWfZLiwAyOXdQIuHr7sNEhUfiX984NNv4o1jsp
fwg9Iw00CWLF0IDNDEUGxJa22VqbBMI4SPiV2qqBv17md3mrxBic5xFLlKUf/pu1
KO5ABOjsWUunKuDKC4MTRxltrlhkMttwD6CfCBiCB6+Pn5i3h1HAfmu274q3G3XT
pPwzqKiAcTZaGAxIbRUw2Me+MgRSxfmlEXRGQqb4+ycwknZ9i7GNPBiMyDL1TZIO
nQeiYwDvfh3B7gIx7NViUf3F41Ogl9As2PgIiTJaRjciJuibR8nPbSWl9mUNGxpD
x+Kpmh3HSrttFnfGkyM44srBP1UFAksZQZC1gkagHw+cyS6lFZAPdUI/mBC+gH4J
T1AcSJ6yo/o9LLBYM7tmaufh940Yazx4Np67ZKrTFyOVo6MWU2CIOnNdDMPvqPA7
h9qDT2GLFApnyGxT9h2XSC40PKFteUxn1h+4GyUjLrlJFCbozQMC7/rPMSrM9A0b
5a53Cz1oFm3nNmUosFe0aCn75uzyEJ6XeIJvZmZ2BsaM52OakwSQv00dw3NsE77w
7UuV+UejnKaYjTGd7CvKfse/WXAd1fpg9ddWwW8ap0y8EVjboKQY1XSIX+r8Ha1U
pNXVrmVK5+OXBQNg5VS7rviW7NAVsDtcPZhcF5mpdHB+n66tOFR8u1f5VLMm5V9+
6TyoYB1ZK3CmRQQh8E96EdvVHYTP4dmg9Mxl25uB8JC0kkxhCiW/R9WZ6DtHmdD1
OtyhV7fycopgLhbN2yeoolvN6nZY0I3NTti/n4EWqLvdCbWoEDKSf1EYE31E/Q8a
cBAtlUFdc5vDXXoW1FIU6K1RjS4Ox6A7Vvplmx8q9gWoK2u4X4eqXYQ+GiYj5sm4
SGd3ozoTyLhvLNIohQsE2RUm+h6gpjcNI8eI+mWGQ7ZtAt4fpgFhws9evJy1Xxbj
nDF6LmLlMngViwS8vo5ci3b2wLsPb594VmghHh0dDJw8mcQnjlhoaWy6gDxKiHJx
Hvi4ecZErrYkvKLpmFUV6w//iGeqApXhpJ1OImxflK6SoNOxpzNudO/8V618zgWa
ELvo8iGTs4lb2nbgZDsFriW6IHaCThetHsm9iLOvkQTfnrN9v4waI/8mTbkjjM/N
fhruldp/jnsInUDKOVa9aqE9cutzTvzEQF/sN6evyPsw0EYFaUJH3It0OoeGBEuS
cMTHXuTdaDfBit9lLNXnmMoH2ooHu4vz3XJITklz/o8AdxlCukYq/mr6PuGD/D2Y
o8rnAjIQI0v8yyDBywk/OFwRvx+/wGB7SKqV+BIXKDWHJLw5usPDRD6m2uWp8QDh
rnVYesymdtgQimWtaIP/iXfVcy9sOAGthB52PEXi8RSw9TlMFOW10ZFwOjPnGGhN
/woeYruEK4h+nNY8O73P1I/Eurzc47J/EDwksITMq1rPj9rJ3qtjK1AFmu8Ib1ei
FAA2u9aMQEgWvz6I8C1tXm8BPIBDVUqWm92QvxdTD02s46bk3hC3NizHYOCEVUQw
k7wVJs6QQdoBNzOcuHJlCITzDKynheKF7VVcQ8Bfdy6r4dq7dmI4NlobS+OlZVWO
X1x7wn+SG16TsKgHAPec8wlnkJjikGexCBMBz+ze2ukKOrBd4ncdLEstcjLYDfaU
GEjhb82kn+dlCMgk1BYBRKBn/RwBVc3FlxhimeuYIqpPwJeRgQJ80A0AKCuAkLIu
O0qYARINT07UFiV9K7mfOa6LONdG28pzGA9RVewP30Odmc7tF+6VeFDHR7jqN7FX
JN9rZ3hC27b3w/LMr1sOsAcsxsHhV+NIus4S8hkScJTojU7T3Et0Vm9DR8gd/KQj
E7a9vnWXL8ZA/os0C2gwwC4wfLJWVwQPhF53h7LdHMneh1huQDwZkiKN0f9Z/b5b
gaVzzotQCiE4SsJeMljv4o/xLytX1n9dt3kOcsAZNWo0TkO1sST7Og5BVIYBsCaM
xr3s+F6xEmeZjhPGHtBe+NbZnJMt7oJMPkN8cDO+NMRQFNO18x1HpXZQMxB0GrJH
VSgcOM5VqUMzlsYgOqjWCWXjGrHCcZNRBXpQHN3OnI5ysiMJOiKgPgOAD9mrjB0W
Pz+6J6I5lu2TtbQJdiJR0e/TK6+Jojx47NG44qNnMuNPCF/vj+aIRhOLZMSRWUWR
2No7ESmzL3s5X6y897t7n+TYFnRuPMraJ01pScpwRhsbA5tCZP6hWkaGEoF5ET2u
yx52KGh8Jlos1TyErqKd+y0sJS/bEsim1aWDJ/OYqDmS5UYQj45B9pibTBpy0fOY
IPG6VZJCSoJuMrk9//D2LfeSyUOxC+3qVVabMl6DF2HhCMDy6tMikK0TUgap7ste
A9ZV3JwVizE6qbmlL7karzxUlCZnZHIaAuWnXzZmsjl1duc694p8yuPx2W7SYZ+A
tXuU9KSiD3qqm9ndd1BY6BLHxuRHWl/XFRgvm68hUueR4as5lwYkNQJgsQ0QzitR
CdLwk1XB0BsdntbvIGPFcOwNmP9hluPsLPzYkDPH+y6BCXaRBEUZ78wnWl2+rXoI
kZziREEDUSBySmKgj9M1x8JIhL6rsgkKRG32HghkSBFjbkZUiXX6Xk3FGjOkEIv/
FnYckJXzVAPEk889Vh2a5O1AuZKd4xXVWiAyak7WD+nhPv102Tc5jp/r2u2RZCyU
mP1pgYhzoSvDUPxXnNSiAUvFsW1kC/Q8E5PqH6XPyYUi+sH7ZF27rDtgwxoXtqBf
kGVdVg0sijCdedF6fyUHxVPh6sQH9a3AunDRdRf2RKkx8L6eux4lwcCNBhyKtIMj
nlMF3zzEqbK7RLo14Ch3f/EVAlXBWVUYwNLxp1JXzprgo6bmLxZKQ3/2M0wQAmHe
NqWFMF5UhnOiJ3AAYs1RsD3stoUGNgb3cbNlrmrhVzwY8QY9/AMzsPgoO5V+dpGJ
O1QOlG7S8yZCAUdsF1lj0122vDiymgB7IIdVcOhXGQUPKG1tC3cEpYTTS4/jtYGh
f7QnDnqEep8X54/uB+Zkf9jkKga7u05kvywau0Ksfg1Bh+thIVhKxuMwza4NPVyA
GwoyiH4qaAf/80NFOyIT/LV+K4No2799ERonn+dDpTz3RnoesdW2bQU8FKIETamB
dfgeieQ4t3duCItF2S2WnGyp9TAzPCrK3c3NT0Vm5fbY9Ua+AlDeHnkwfK81lMSH
gt+b5z4oKMUrA/pIRgae1QYJpOU1nAosr4vCNlvpK4jqRpFvxEjSHHe9krH2/ppw
n3W4t7oWl6HwTAK40vGRhDp9asUZMcZ9462j2du9CMjmprm2NOSPOFo4+0n55LLU
SJkC8vGbA302lcx9tD7jcjcxTJkoYuaY6ZU+Vtyvodx2AYmOm2S3kU7beJeCwxkU
dJToHtbR3UIner0NyeqFVI/tuGY1SOvvE1tgdLZcAGTLdq2/AXyplSygkXmhC4t2
2+FqKa0LiRNFcYmU1kkTf6Nc7BPx6J1A2Ac13CZNppiZXlghR9zGlbz3YtTUSbiQ
IACvnKP7pDjEmRe3vNKrePihFR/O6HBnHxn2FRGdtj9uu+bjQ/g4fBqAM0SKNcK9
0b3YEPZnaqlJMNYYeaDUKrI1LpVpPp1EdmlPgjcJ5E+35k1CDzRxck7uzjA0vKMF
is+e+vuVqoMAkyXh9qL+MAkj6oqCMHy2v0fG7MYBVngHkvfVpFOkvvSqiRYMqiqn
VCgMYuwL+a2GzQMK1321stiOo68C/SAD7vGEK22Uj2DQB3AG9dyixC9dnrkhDYv+
zBmNIge1/UoYYCd/1DmH69Vb8bnR1WgxbX15sD17XGvDF9vXEPfFL/tK1nRQb/jT
jtCt6HaGFWgb89B5QF6weNZmP2yOMmgzIAQCs9kibyyh7ypwpcr0i9xGvJ1SvGTl
3Eemmx1RB7C+qz3PZccz99s9oV2fhiYh5hNFLChLjZvjOJEDzMb0Oyv3hSP/kgip
PTez1AK64m1T+S6rb6GtOMS0GWVuaJi59ZPt83FIqmWPXoud664xnGEi/COU0JS9
OPZwdho67N4e6KsrISq9RFGGm3gOZ1bv9sTXCJ9YwzWJA5tiyTPUVRkzDyfAIf4P
/kPvego/oeKrfW2jiFq2JcxCuHOfDsp/oT+1/APR6SBPeZX/WBySoOXF8NXeTXxT
DP2DQ2YpFuUlkRtxblTO1fMVbgwhtoT0Fp4AXd4AgijpUaAhRp8JHISbrRDN0rYY
aVfywwkBE74x5bMEX9Puv315B5sNo6V42GL7X+XnTRXA6qX4OtU6+/3HgaMgul73
qLbEmFj7W2Nbr9oQtyfyFr+6XSRY4YqwpfKrbG+S+I8R7kVAn98knwLLU3+n0KaK
YyybCKnx7hUl37QoRCf1MSyjMln0PHJretX/uLa1PG+RyFmPEedfVucEh9Qery+a
LiGluogJeYAxc5euopPMfIQ0mZOITcyXu4vuS3/o2njuq2H8MoE+24hfFt9uT/8b
6iQym9/bvLIAcn58bnWZzWH4CC/NPU7Us1PLcFBUDz75IqadXXuSDIg0D7BjDzP0
9286L/CM00vkI0AQRNagr+BMJEzDPUmywwaCQPCxYAjgo7IpA8R8wDirvKiry4lU
gt1L6Hi1cwoMol7wViqPV6k2mvuYrXSXdl7+zh44MtpH6qM6B4DJBJ5uHhO4lJUO
9dZPdCa2L9u6hwiw2tfvZGDJ9cNHv/OqtQNljraMFin7ofOxZNVbnceMAQzyFS+Q
yC6tbOFFvx0ImBZPj7O6t2bg/JKETgKErFmbGVmUbJUz2W5vIm9+yoyOHDM06NLy
YINfZkJSds6gcHWvcnBt7YMcH0bKAF5gfes6Yk88ML9D2RBwsZBEEbn1LktnrW1a
hT3FnvbTudSl3U0y0pBbSqkZjHPuHuqRNe08QVLl7QOnDcW9b4z49JGbuMV34x2I
5eZASq5zEMEhfndtzQwmUDNNfk0UuhsHmEIhMlHNjHKtwmqBNvFjD7km5DToZFGH
n9T97MXoimX2LP76LqiuUPrSdK8WG7PE06loXJcPKRGL0byEseePy6NpwMSKQJeX
Z1TGV6K6LUqO8aJMPE7JWNob9seLCu4hkH1ZFbrSEW5rhEX0g9YeEyg7sK3QYQuO
gQlpzknru9pZTOxB4ug32hh18+1Hyo1hB02wk/E4L+lez9KvJBEMnIWWWwgKZAj0
YDOVaO9PjdNYbKvu4qwLmvqIVjHh66L3uEWaa//BfPMooeqE1IiHHRzU9iWf/4tc
NRiwSIbDPxztOy8cwG63LFpQClKi9U90azAgubcZ2ZQRHMzqPu2KxMVwWPdEunBs
GGX9m4MAaEgiIUvhD7xxTlCZ1A6RxaY3KPRkqJH48+zdTembwxZ7NrtUycuGGfim
az+YIp5Yk87p5erbTnV4uSaYreHts6fH2V25xUtE4R/8zXQpk0xOJ6pZUGjL4ezp
RgSLDWQ9iE9H5UAAj5AxBGuAG+9xgIXHLre75DrCNCfzlfGwIcGqe5ev6IU5FNYl
aORhzm/fSlKwZi7XrP/XXWRH1ibFxL2GRopeSLAfSClWBB8ZEDr/Hi5bEViwMDxi
Zu16sgh1sD2UtN5ZufEp5lL6R8WuWYCkTsk2/yyUJh05k9gAhvKK1kdyMCy0Itr2
KqmTL1vdaHcpTIvsRmrUQoU3K382c+OVXtZJJqAiDFlkNcd/4j7Kj0YkNYrZxivP
NFZA7BDrD/2ohaxbpRpVhvU3zXxCofgB3sbZqpXNK4gywnmWRqOKrlnBed9JSFZO
EqfJFj4/6whzughVDp02FPaHuVu1rPPNJQ10Ekd6AJrCYHkb/riE75jQawDSp7La
Bah7VEq2WrP2lAcvhje94EF0fXyAdyb8HxWOsGJfTEptap/tHpXK4OwpEfs5Jqfd
HBeh2WCiahG0OgCAEZvQwNgVgX6NZCPU08saWFauU80PTCLrywXNi0tjrzdadaSh
Ficnzvrc2jjt2l+DSo99VWtAgFceijqiv5gcLNCpDBfU+5GoIt5tYRPROp04WBcZ
5N6NhM/1fhXY+qH60WjZXvAFz1WAFaohNwMpb62BS4kO7PpPNiuXs7nLvL60N2N4
GQSiV4o07dxiCuaFR5uvxW2DVyyZaI0ijZYaenucHejDDMc3jcyiF47hjcrXMeJn
X2LqcwBV1xgcCrPhmTHoK1PfFH5WQzTEQ6jPATfuITBNAPb0ShYKTlBQt8VoHzlw
Ev0oTR1zx9IzsiWAGPT0lkh8fRXKnH1Rvgu46rQt9S3jMXe5vbVPPJzotcvXgT7E
k1STqb1dhTFyyRn6+rmJGgG8YvZJVSc0J/zLv//1rnkXiOYxgoHLVtpPdatWVACf
IMYLnH1y2fF32oVu34Ju9/xlD1FAbQ2XMlXbaNKAI0vNfzH5Pw2rp04KvYKcH3pw
IbOjiVY8B2Vhz3xt0GBMUtQLGw7pgV0eQHNOVe+UzHw4Yd8tKozcv6YV72jubu3E
+RSRdmLKJ5rEhm4m6k2NI1ZLLGZ5I5ROO2vPunBv0E5xDGdcoyiiWlGNd7WVLFLZ
B88eeLcjLMgmfhMj6ZmjvwJS5U22UuLyBc5hsGEfOVmzHKJTVSK+Nzma5DaRxpDn
DVHJOQ1NLKx0xztUcYTlGUL+TGp9aWfabpFv/7NLRg4DmZLN79xzQatdGP25Kvap
Geco87DUoau5GSWuchXzLUCpBqq8ewi/kUvYdYOREjAronBrvAK7M4esbae1bjS+
LWHKt1+31QhsB6fPYq4Cy7A7MnNrae8+Lf3AnZxKwJ3dZbQzrzzmVVjECCtKTuvg
7Yj49KB/J2VJR1IHFgReAe4gbqV9Sq2lbGAcBsmQvc8Yg4B9OIpJA8MtI1VWstcL
il7RjTpmjvOSKHyrTCsIXxCd70YbcWySpBg52AOXtglLtmKRzC2WatOyoNNJCXYD
MApJuU8KLLU4imYwhxUqfkeuMKCgjtHZhD7/Ju9guRk6ZPvLunkS2VSzKYkiuhp+
BMLpEh4Ol/J3kqYST34gyHbB78Sg9SNCOyc4OtBI9l4RVtjauf+vxGJ67koG/CVO
pmtDg5/dwmmNybv2jMNQXpRAMFqYxz8g3li3tDTZciN7EyCkltUY6A2Tlb373tFF
9oAlRjOySK38ODN7IzIwHThGT8ZiqlZM3ffGHvVTuTASWG5/Poqa7Ue2GomgQy4A
KoxIB882OOKixzQ+svBEHr6PAn81s82p+oGPMzBLLBUBeMNi41/l5foDCcy6T5M6
P+65KGS1aKV557WC4Q8reooKV9z4/HInkkN/PJQZ5rTW19J6Op97sQnIMpbk3qP1
dUV2f2HGy7hZMA9ygcOV5BPk2snAg1tdCgvtljMg3ONmhOQsGjlm01bqA0g4Ddr9
XgcWfTGhmNGPpCYWJxXIpRwaBJ5rr3ocyoHM0OD5iznqexxEJJN1DE6Otm1gAewc
wWzhBcswSSXpIC/s53ViKMXKgQBjCndf954Mm/Mqp81Umxo/KPNqyfK7W++eKT3F
t3y4yOt2INW4rDtojxLzyQi2STmSpuE/WXvpZXBvuPPOLG0cXSN+Tj1A4XuEr7qk
PcOBmDPXWaxMGwTQtV5SpRvVlQY1sdVCs0zPsRAFWPrWUfUuRnerVk1Ewkz0kzBm
xsB0Ma8UKfZvWvZgUCiGM0wW5wDhwbZU8gG9Jhlpd4yIQotE7y+Ag1jsXe5JFzhE
FuVbuhHqlT2s4QbOyD6pfeM4c4cYdK9wAaGZIY2cQWwcUbRqEId6KkpSkjM6cTqq
gPAQY7aTxZIjGfB5GYg/91HuvU3+sa/+X9NQX5fJKyC49bHM6gO1f90gte1XCt6s
jOG9QhhLu4bGB72T7mqZVm/ILmujI6TXD4tjauG4jdiIMg1E1ez91uG3wps44O5u
QnUN6YdMWbi3eOG5YKpMaGMRP+8qcxth2AFpthRCt0i+dWdHBtQOSO8QAYo3ulFd
0+AO85bEOZzOp7bZg64Fp22PXV3/M0RcH44WFEOifbo473DLnl8VK+TKbIOxsi8s
KzQEgQdKHzvG1IAwA/hlH9LWiutVlZ14HMjKtr9REwVztw/FZlvbvM+AK6Tv77Ro
lHeCol4vagMTe0d+Wx5qMkxKkwGZ+hKhZw9zmmmXK1Vr3hnOgyBRfweUCQFp6/+1
QKs5RpxBdPxUMVjXXtfr6mrmEA6EFi1myx8ynHFr+0QH3QFm5uKeeIjfsIZBJuXG
9LT77kay2mepzANMtZ29kFDzQn6+7qk0sQuIetsG9M9CGtcM34sIMhKKl/pPRJO+
tMKqnTdx5v724v+P3Kn5/0yUdfk7LZh4hkZxjw+yYHH5EO0Dn9Kzzm95N8ILiLPA
BFROR2/x06/tRdUdKmrTP5KRTTAyEXoRDShs/CID80RiGNNtfMfFJtzf+mLnvJbO
21V3dYntI+1hz8Gvu6WZRUjk4wMlVKRyu24m87tDOCqPVB5hDeWYFZtC/vEO0YYn
gfldV0TL9GTWpy96es2hh2hiJ1QE2tDUtwPeK9NlqPXxsLPXwBHjjV1dIoOEGt7D
eHlRf2IWQPSGaUE8GL6vWhgCqUomXguj6ntSU7FKUGOUqOLB2hidT8x1jYdXJFeF
+SvjeL2hDnLYjz9Pv7L3OCyeaLd9YuGfCzogtdnaBdbaO39UW2uoJFpeIZZxo88w
m7WJ7O3YAbIbNCclqqvxCtCRcbg5OkX0KxAlKlKXoq7TruzkqaJpFziWNvQP/PQK
jpLyikPTkstvTAgEg0Y/jBeAmE3VDBB5M1HIqhH7uXqMsXIItqMEi1Y+YvCExGpN
gznhUqLaR6ggxTlObUJWORj668eJ6r9hXDusc3gVxvbwbr2XVo0VR9a5KDbpxcYE
/6FKqiCzl+G7GZ1seU922g15046benAUE3Jf/Eac8UPlwgZp8diZ9B7K9RW25d+D
lmeAJQYzs1MI4hcGg7TIR6QtTCkPuPDoLYkj4fSX8G/11bXx4JuqBsQaZkScJ4yv
DgTR7489+5vT+Rm9Fj7N5xzfgvXXsYVw59JwhWARUpBD4F5OYqYNRLFsfQQrk1m9
m6WUBtzfADoP0lHu1GvqONcD3CIwcbCaDalaeDHbZnF2Hq2iBePi59LSgandBMFM
+1o+/Xesve3BofjGiX0XW8fnA37uXe9XoIEhLY0r0oly7oXiDSPvWeYr3zgq5+ZN
VC3zpKGpCLgMNll03exRjfIv9RU3QRQX6OGev44gv8Y7igkxwIw+87yryPFss4qK
6U4Sv1wb3XfIfykqZ1yIQZ7CLryx4U5x8PBKJnNjgvJ0pooGBzRCn5BckjsNN9hZ
Kk4wxF5ee61QNwm0YxN6Vhrbh1TSCQFvIyd5tc9mZJgwfU+GDiHDXtPtHuuSh7al
XY5/YwjvEESRrrZPxhviV3zBKDysomRKSnvNwC3Paw9uIplMrTF+e0xExRktW5p9
lUJbi8ISojSNloF82ehQmCZFBt2Cg31qaE8QxIG3aya7Uq7m/TMJ1JS2509D5mqt
xVcT/9jfsSgjDnhMZ2VK3GgedZ+ssG1TLBzJ4f1pG0wumCIaQ6PO54xjLyLmLYRn
GwJmhy5xVG6YFZi5wV8O5jMH+VltxHUcuZ2fXSN/losZ2bClPH7YpGCNCUc40LU1
frxMe6kUot5dUc8MrmKsd44KdpUL1CZbhQ1a2C5UPkFcvCix98C+ylDLamwmq3RE
xa734llFZhm0YZclBgpGTWdluxVz2sj3pR22uXPijelTBfMk/nokZdGfhZp6Er1G
TyFJHLJL71RLlfhHylhhprkwGRKSzAS8zIiTUnd5dDQUuZmPnXM+6EJcHhdFdUI8
Kz0QZs4ZBoK042qSd6U9Nz5MYjfrgBAbiQljMMAojzsTJJuOK35xsIxt8H4+p3ta
0vL/PqzMPdan1aT5hXqAGrhpDUOKLK4PutKbOAvtZpVdgmCX5bB130zFEdvQ0Q2u
Dfhe8FXrjlBO5eOjQ6no3lZ37VGmZXslQ9dh6bNc+s8udpQNn839jBIrPIV1prqa
DVq++b53S2u+QJsunzbVhHYYUnfAOvbac5d1cpKyKK3WmyUDhAGuIWN48gHkPatN
S7m+/pCfH7kOOiHtnaiMwm1ZDeRqLQqk5+I3C5DVQVQbXErThxvJkPGzOM8vBdEx
em5+eP8qsgCkw/cMMIuDyBKF1/QuWK+mNJaqv+doNHSUClVEu9oJIyUn/KA82JJD
jM1VGBgTKSC3Fn5ukGsQAOU3Jb518cW/QeI2pF6CeQN9EsJZGPPQOPlrDx/p8mVo
IZKhE3nbGJQ6opAIHqjgIaRXrgT98yDOoOk0yqiJyyiemhRIKydn/E/ed4rG3s4U
0SnPJTfzHJjfpRWvGAiKcdXOpkOwtCufTVHQ/oInZLGVaAPOCz7M+ki4ipNA6hwA
PHIFZQeuRGNwN8V/4QaBKLiUwjY0rOqwU7YXNHDPosPZ3Htd2OiQVjjA7p8ZbhAp
ifjsFTdQdg1ukfpwLt+PzxQQDIrl1kqT58QRfr/nXgrzhsgCXQcXyxDVReeRf0ls
IGJznfztP3efe8It/nekvY2DSRYEyipA1sNp2B7Y6vFeskoWDZ754HbPBunCrppW
JI1f2OlfogYQQJCYis4utT9tmoQD5786MxflNsPSVgvLcLokQr7RNaK6JvspOSYr
ulkfpK+6GxPMpUQPBLZEo8r3Fm+VBCiNr2JXDdXhMRvxoc3At2+BQmHIt8Vh2bfa
RF9d9Az7STbj3OiWPiKgHeOjETcp/66JbWlNEd+rssCh06wG4g0qcjeCuSsSehnI
EJlRJYMN/CMdSLKhiobjI0xFB0YedR9bz+94XnF52GRmUIxEXJCNFYESsscjuwkS
k6HGgMRITaQDaYXmytpf5xVgpRhp2X5+9SKmyTxSitEiA+WgkW/BudtkUjmuJG3r
A37cvSWhtCKDaM7bzmxgbhFqG+O5cxJMUZus9zD4viUdTKNvlr7n0mTGU7Qb6xl6
zLncrE9i0+zspdzm1rdydJfKJcTdoaO4ENh4yJW6fIiXd7o4lImRaMyZ0prfyrsz
a0IJj3+hPoce+fW0nMZCMc1a4cc40BnUrw4TYZDjrdKks28j7kd62FXp0hp7i2dO
Ph7+An0h2suD4x/wnqvc0cIlQ834zeckTG8OB+WCUaAIdsVQ/rZdHrCFnhI57fIw
0I/7q9qWbmB/SvIxnmyvngnXKUzx8DzYQWAxABuBLUyynnsR1VdIJ70yTgNLEglP
WlMMxkqLkAg9biLD1gW2h1oWzddQkwgfUQx0VsXe7N8yuVNJnZ3TcqTsNtb8vNNi
JWHIk1/xVHwqMFbZv5AD6xtALg5BAYT5dCQVuY9lmSqsONtcNj1BzT+edKcY3rpK
QR5Fn7b9cUc10YD1G5AspLyTyirTFlDbX3VCA15d3K6zmQ+9bzJmm4DWv7HQg5TJ
vCbuEYA4RLMuT6CskHjay40ze8uSe25o9tM8gdvTVSOHEHdCAHATi/teNgTRuWor
VJ2Q1Eia5BWQBGa2d9I6AC9m5T2GmQWS9FmuYZ6Fyasbc5UXKKCAoU1K+gqxjpJy
CyUUsodYlom4NOThSS6B/kakNE+HEk357lElq73dhBZ+xMIMWIubk1jGoZZYYj+2
3AH5KyMNv3tvyc9/Nh4IQNafG7N7sbJXhfah/LB//xeIyw0T5YGLds+LZkXGizm6
ePOd+FBEPQF00XU5RWibE/ES9C/jSpI8r5tuw6VWd817u2Xkf1vtqDck+l6YX4PC
I7V1faw3ofzLoC0p0XkEPYzj5FnEF3ejidcaNBTJxT0F4jtWrdZf+T2ul8j7WE4k
ZQ52IkE2wwznnuKeRLWojNkBpll9FWhOEWJFyAH3kMzAI18vqNY2sGD+ZYx5rxq0
iE/CYCJi3HcTz5Zq58fr/4IVZimftvlDc2GMzV8DV3zLyUhnifbL2dzYxKU/hhgh
DB7ID+cbGT56xH1MNtlNr8dqJqcklvmMoKOHUGxNohZzXMoWMoGhQ2aE275NxEbk
yVUpiNPSS9ui5wOO8POatWhm12UwJPq+nPQ4lSPPcwya13lKGLCMEdZAVWQzrOXL
kbiN61SiQvt+VNYSUcdQW8dTSigPP99dK30Vlbh80lNUN9oxnjbxQd7Zcr478zYP
+d2UTDJqyrZtyaAER2ayM6z3mIx/SDwPVkB6Y/1pi/rR97IINIIFS6laiUrHg6CN
wuZvN/4F0UT5Qd4TWGQR3n//06GQrsKiRgscKoiCeF5U63XaPjBbdU/enoMP88DS
g1qR9lRXNewU9776LH+ab6kVAtVhW38D2BkFxjt/5278Ljt1xjX939En1CNKpZAf
EXxgrpTxU5iCjYIFzO0sbm5DoZOw66WfH46ocSluZ7fnF/yqxk5hrguELN2z4zls
CFXnzHFdmaYXpkKmMG2xwFj6c+KttxMJNUYsIeOMvDtYq7MN0nf5v7Ca48aNItFr
gdg2Eq4u6cvSb0ZKWeoIwxfwdFBlE7yDUsrt5VNT3XUR6xHpYFGODx016523md4G
G6foi9wld3mqj8qt1wu2dAazkQh+O5QOqc19mGxH/zASoYVTZ+zhJEhuSFsDtw0e
USMQYVmppI4dwb2tG4xOO7y/uZYMkpr8eMd+wLf6LVQbmVe5jtN0waOBBgoaprgl
P3Bw68S0HM3Yj3iIGjYX6stmIplsfXCHvsRgZvtFtFsw/lW0wG5VCbhEo3moVmN6
FGGDDEo/KGJV+nF96WT51TH1jNaLiHQqLxHE4DsVkyTxMipcqGRPjYEQTU0marJd
HeVGbSjSWqRhxTGiK4VZx4Kz0LUU2wrbhljpvpF/R/K0ELls/zdVaL2ohTfh11uf
7T3B3xQoHGpgDy6fjuYQjNg+0I42DA0suVVm+dPgSoKCgoj87QSl3j0kC7nA2Hr2
KLQlxEkAPtPGDscIgwRZXkZjLQAAxALSTGaFwLf2dwVbr4si0NMXpldED1xPbvDU
ohQJAlYMhGx9fcPqD7qCQd2TO1XPUkNbRMuTg084NKV5fecZWp6uqPCHmlB5ejaW
COdBSL9DFKjSToFobbajBuhs/9UQAd9PEX+gSCBKI0+myhKz5Rb4qKpnHt1nsdQF
UAv68ZmdYpkL9zr9f0tPAtrtvYKFbldfsVSHzY+Z9QpwaIKD6bU0ruLqtNRx0OD8
029LanV7yhwFo8LdTNeexC5xlGsn7S+PBhNGUI+5BYXM7JpH5W5ybcLJnlSYO0v2
B7XsCZmaJ6wfTABSkujU5uBtp+egZ6Wx+01B4ES7shKUDclPgKQkxVeyYCXAwnxm
eZqvO5q5FqdoV7q19R1PvIfe8n2NwXQemRcRZw75/+eeG7iL6/9szJAxDEQeo2xC
ExL54plt1sweMXfg5A4ITXRqpr5ahRlP+bfR6fEFOuN2WPdKeE5e0KPWMrCcZdef
9mfh1j+xLDICA8isMg5LmxRESYKf5KjXICaFfJER5S8JDpf0AwVH0Ab5qDdDu2nq
wM2FW1VFYiqsf+3ClBNV6w+KYWRIxC7/Tou88fEhBX/s6s9NnUPOl5h2xovmQ7Tg
vNXw8Bh2VnUaKGGWMfulKgrY+vzEiz+aOnAFTaOmVfiayHNsUBB/w0N63SMNpaji
mlpOp9NLqP+qyMdyK3rT9a9yRJ+0eSkiBj7K13ioU1G8X6ry09tn+vIghi7SUVkr
pSFrntk2aBPkXFadzrGvUzVG/d+yoHLfPpjH3UgmOMzZPoZYps2Ni8X0XTveG7QW
CFardy1O4aNYZ/G1udWOfw1+NjR6rn8Kuhpq8vhZEVi07ys+WmTehqp/a0Iwuk/Q
bja3sQ8oqOSv73eyQ5C6EQy13TNvIF3hMpWd+9n78hWK9H48X5zHoRyfPqADu3jj
QDGUp9IQT6wdjjbLdwyb2fv1zutzEy+tMkPVJ1esqKcgTemQ0UuXoe+SW2VXVsGm
gCwMkjhI/OFBVznDT89wZmsLWNLipN9HNC/FXJJW20Kne/E5cZZy65cAQil43GWJ
sSMkRkrElzDCaM/nJFeEmhg/fiNSLv+QERPF+nABGGJsovZxhti4TDk3vH2GJnj9
ajMGAfec2l94N0hfSBsjZtmKFFHyHwaBJacGQCgLBCnlKFebdKeeFagSIp+y0fS7
kDitoe4EBrhXdNy+CSbXh+Pr4wWCoH2ITTvgROMTI/aPXsY/7spJUe9TZtscLXiv
TziAeYPYdgD2TSRWKJEJE7E2X8+49RYbRtZgVeM9LtYj+lp8KejLQjKx2Ye24dfn
6GqYWbyjadonfuC9zGq4ligyiKy/hiJR9Ny75GxtVl987GF0m5W48fINJpfg07JY
yvgAdirUOn2P+ygNdKlfFw6keHARhyYvWsfSFsJplRKrAEn4N2qVILJJXmCqIwyL
DFQ+tq7wqa4bwq4v7WK8IChfrE4ln3UMVIbgO+Fka7ivwEfOwc9GynTK6Fy/l05o
/1GZWevSwd7AqcV+6o7uEHBqcs8hfZanzb2lDGlC98S/ab79rg2i89WwgVChT6He
zd8vnFwdwEBX/mNAZPEELLGMJdjrfX6w5EnlZRPhgIkGoenGO9gUl3iHX/lwJZrY
DtnNNNV5uL4MQ2GwDBCWuhlaRLBnNumYQf4upphD7GhZjPcSCGqcNRqvuyZwT+FT
u6NiqxS84hndQBw6S6xy6REE+If4EyjHPLP9sNtfjW1EjOEVpYOHWa/NpoJDMoMJ
dnEHAM1AtPZeHx4Zr4Mrf8adRK0Rr9iaEL7ysabaJkjvmuQJys0u3hd5nK3wjO9A
tNL0nsHhmpSEfrabXcyxeKyDgRumEiiIEme4tzTNLQOpZqXEs/nTdKAYQ+sa4s0S
3pvCNxgBfphttayvG+mkv89guwbIX3ArTKgynUUMXNge4XMv2eVFEU7sLPjc5qD+
OlGO8zTjjt6Xa8pAvjWrBjwgOWvEiwLLPrp8LPKh0qJnJ36uMji1g+VxEaiw6Yyf
x0P8dHDS9W6hbsqIUZB4ZmEC2hHPxjPuWZMEmDcoF4PPELBo+GLpx7sbJke7By2J
OJLTS1uti3lltOQFWDKMRcLG+pFhYuCjPtiPRH72PZ8F1KE9uNw4TCrXYIPbIXOC
KzS0BSUtZNno173B5BMXvVzA6FUWxlMyhbxIxv9CVgAXbgcDC5gt+/oDDt0+pxIn
adCXFroQ2Ynq4YdqWcEI8zP8Zw9qqj0h4FioCLC9tR/GEbegD/nuDGzfHg81Xgz1
ubulZ8GJQrKiaIQxdTmnq/hreUUYEvvdmSz7+J7hZD7KBWvdmdx6n+jHtGe8SP2e
9ZmErnUwpifcVCv4j5wt76gATEq7BCPXk0XBmggj8jdalSewtQWzs7c5NhHdXg7V
7xS1b6UBGrbZDtWCzm2yhtLyKSgYxpPo4uHEP5PpAtSbR+DUpCXzX3Ss4PD9H2HK
zto7cuB0KQh60TLtlnKNGu0iz1vg3dsiLnRrlEE7HoYUJlD5APJyXtQQX+dA3Xt0
8IeJua7taN+3S8fvoMNFVLjjumBrdJ8DG1ea/xfSiv8rM+CIq7dtwY4BjgSfZD5j
koiN8U1Mti3Mp73UN14ohFbA2uewmcmrRl9KWSf8QQL2fxmFjFN+xKkKhhjUFOUB
SOdt3nFhEFO4ik5Qd4qDmhjaxCjS+mZmFMi4F1QLoiDzI7M2NOmklT10xarlPRC8
wGCB2qWyOkTb8P9GUToHGXqy9pIRai4pPWJPnj79jieqZlxoqAU7SzuxK7fvuRRo
9SVmvvaezfdI19AB1MKGoJtWEhdZxWRNZkxDLSluvKKdZKeg0HqOPQwPegXgpgxi
6kHU7WzkMs4G23PY03C1sSzgOr0OqurBoDTvMnBBxxugsYSPsG8RXxmrmwFvPh7g
U4Ux36SQlsqCv0Xx2SKlD4cG2bDKPtR43XBoG6UPdBuqlFvoIgem2nsamBFfnMuJ
KuxFAfxa0+yZ4qJ9KpCksh9ycV5VKhmlSsQdmP1WYoInHEOC5oIcPL8Df9JcWwkq
2YiPklYUW8dK9nqVgFHJOMtgE1iKpp1OFl1Y6aUL0/effupFBNuNViC7lu867wo/
qa3vX1u0ilDNs+94m0T7DR4U+JZqEIVnD410VVjVQI46+vQUDdbeK5geqb1re4Jk
sGXNjzsp/zbkwy74U4/y+pXu2mtsL/F6Rfh1LfhT0qiVV4mbedSBqtz6mKVUhrkJ
LRU1vAG4codoYXvDISl/2XZwHAmd4Oc15Av/15Kbagu4TwWtDN//sS9L6tev3gbx
NlSAXl9qxg4HsyP3yqlz0g/t+2LFGasU683gnk2uJYtFcJ3Ej3jrhGsNefct+Meh
FqlkAvb861AeWJcNgKMPl0yKB1sGXmSAyY0HgsUkmq2n968VcFej/76UweyTCKXN
8DPR4bAhNYA6xIm2AiNwOc225FszukFk0sa1Z4Q9WQlGz06t3X/DtJDnEPFELgke
9MB1rVMHGsTWFjeJhhk7kG2KlpkDOc+HeUPQhcHTS6AphVD7Zn8sUMKvm5SWehMG
Bso4B6YQMkP8Gq5EgHtbDw7He8b9m4KZQ1OpvtWcO1xQoCoAUfHMp48jceEsDKXm
bRacbj0qLlZJrS+HL8a7mlL6cXsKb5Y0YJoVLChupyQHjd0zNPlRhAq8lcKFJ2qF
pFMfHffM6WNRVpVANnKNjQiwtsQivgJcliv2QvyS8M6e7gZA2ze90cdR3XPGo/4P
hYdBMsE6/5oRlYIVuQnr+MPDnI3k9w558Eus5hazMvzmtNMDm6VA7ORqc5OVb6Pw
C/BgkhpCz2iQTif8TUGOtAD60VRroHh8lhPRHXVJewXP4HhT/NKUCX/lVon9cMPz
L6v7MWYvS8bqR+BXfScBudmDVkj0eWZVhxmuKEr/r/Sizb7zfrNR9Hrnqgv7SXdk
eTK4EdZ9wi+IbtFM2u/SSWEb22SqBWdEM+4H+D0VdSlnsETm8l7ln0uH0F95a6I1
1ZM9u9d4gF4ovRfKzQ+AZFED3JiI4zrqZ5YhNy+uS9VWsjDMMY7oolPN1RfoVM/f
dzrSUgj9vDOqyhxXjWF/gDD4CKMazxCo0LVIMHlWrshah4c9EyEipNAYz45dtlof
neARZnHIW1PUkYvDsRS+ArRGoVi0lzpFBcsl2s6SXHIFMW+DN+P4wwI0wSJU1wvN
nz3Am923kDfnE94P7SKdxdC4rA6kpu6P8UZKgjq76NPmupKJyjgugELUq/xjwdtj
aCy9CXPNhiXZa4BZntDGjAH409nE7V8q05v6EANfcNZp5x7zM63jLrCx1YwHxEmw
TvVvYyzSGaFdYKliF/jWLF93XhqYKXJ9mQaa90pjWbDgbkb5g1O5up5hLgIhQCfH
+GR+J1YOXw9s35c9rMaDBaElRqZYA1R8SiOW3hoIVaSinQS+WWXBLoqLlM5T+kFW
JyvjFDYVrXGWQ3wTcudEh8vkv8gcDWbHqRZTq8fR4oawnDUHsrUI7AEQfsJxfNqR
K6TuT2DOxscQQPpV3xEwbt6IpMQO7T82xJcT51a8F9zHY7EKRO/DNaju+9KmSklL
aDuW0mV1/flSyb8SoO3HRI+nagvHnEtSbna0MQCmL6ND78MvktDiqyJNcmtwsuZi
RBmJ7DbdP6sONMrNaksldCBVZVd+rwQXfvdFOgBF63t7wRZrK9Ln+1FwqTvRL/5V
UIxcjO3ewZnquvrINM2FjQ1yPUKoE3+uhSFVQ7btMjxHkE21+4jf4cv/EVWbWZWv
DfBoSOvXnlP9krHxBhEGUvFetsAluFLEdCtpuaooiRVV2IezDVDhKwFDL1WEp811
4Z5STHW96WY3atm1ZHGQFxZb0U6vnV3ZscQGlq5IYvfkkMpCTbYzH9vTnSBGatpI
EexKcpLqZJYn2ApLvaZlZqhmJmXhX9Ncb7nyQ9pN5oB1n4S4HJFT/OJ/fN0RHKVn
zGae4ADNCKFIbRUPi7h+jwtGXuVZD44hTnnSLiORYHfWEVWTsFdeTTOO2Qw8x8JH
6Ru1UQTx5ZsZX91+Y0xSx47NV/HMRcHb1mZkIIcH+NOk7Sbr977n4wcwQ3GW9JOJ
qUA4NnjP/YTamJPrko5f8h5n7tgnwtc9svS4rEExlZYxFF3lww504wSTh6rEeROP
6/U7BchNSQvqsnmvL7/yWYpas7l/re8mZ/lYUEfwWRoUJWmY1lkvITWqqngGAaLA
8wgbXC2Zm+k9c+7/xNVo4novyhE8Gq2VeoEHLHw+LviORUV8LW45Fnw6me3MSEt6
wMzIvoIo4Io2FA4Xlx3teXvfTBiUaJLcTxOi2DRacVqRHcyvVujmm9J5Ietzwaeu
USGLPTxqtnw8e/8Buc6SMsdVX6RDc0AlEVa6Sv5y7aWzoEu949MNg0X1xuc8eE6n
86TfIVBcwdXEpZ+HiPUgOaUBqlgwIMrT9d1q7a3jngwhK63eLAMzTgVsBCMkIM49
gU6gMyfRkuyx49ahred1CLSUBkiMERMURLPRYTfrRqb6EzzT+iuqiajP9OOc7uEL
M1DlMueddzp7ID3QHcZzgv3cg/3IDe3/DJf3pygvRQ8qTSfeCg4JjlWYRHfszlQa
0qH/fVcvSIGlwKNCi0IVZwqAjIQe1PD6YV7WSMGxx35FlaHA20qhFxvLnHXayNzR
fd6t2jlLi7Ku0vj8zDFTYo1hKxHUFrQW1tjKu4dWdsp/huitfpilA8VRUlDx1Tc1
m7jfaPu3m+JnIiVttOkv6I9sFi5qiwTlycLM4dRigzqTBIFFjuMyVvqWKK1kbLh2
/QROFo7y7uJENDmFIhd0TN+dUaRxJ5Uug1cuINpgHh5j3krdj8N44OSjvaOP7VQy
RI98gL1sMpQbvJfwnN4OuKfXgFHiJal8WM1Wfz2PL1lI9dcr8mleKxDtc3ZxQGeP
0/fC5xPzjXQg2SKMW1w2jz6oHqiYjUU8N0hydWm+xLQk08hx3pyuwuVnEHqpHrYg
GNtzwFUQ/8lTrXuflrzqjD1MAoMj3W/FoTH3PyX0vRP8OVRUL0GMxgLnwj9ogQnZ
WT7n6xUU0YUu8CJB1MqjZXnfnF7AhHd/wHRNrBf5d+Sl7EGQUo7G2+s9BG7ow15a
sW89gJlR+xJ8N7VI+gnnEZMWn+V5XlRkQA2iJI9YB7ce/yILbOXUAGtlmZYl98aH
NKVelOaeuDz4HSboLQ8i3Fa+0Sc+XGq/cnGgwddkgscrLCmr+objR60Ua6F0offt
D6JDVS8v4Fu23iSJVvIV7NbeNqh6DK+cvAsdoysa/DJ7iKLpe7XYPeQ9JFvtaUII
GwBvcBOo+wGv3egrkOJnR//QuGq6tsz7Ypj0++7c5CTkLRfXHZV/zCGfmKxmuXqY
o7A3yXnd+cXX5LxBDKBkfrfNfLmUFb6d7aZ7Q0MDirW62JeQM4SHwxAmtv0xrr8U
GiQg7N3M6epwliQ0aOqYesm3GXpQhJLO2Y9KtD66C8fo0Dfw/pCWD74U8OyCcX7z
Nqh0sgW5GF9gMqhAZEHZfVhTWwf9pGAb03Hguw+BNiNJmijr1Bg0kxKCrIAQKLGr
/FScfqmEK8QJGZ7U8K/62yg6Du/6GbrYu4+iuU4PssMmptTsIi62cK2t0T9pn3UD
STYI/MKwVSWphm7fLqoQvSwWjuyMADmGX762ZCeUgtmR7Qx9I3YN70BaJj9FWU1q
o9ou7IbYAZh/T3+92qMXMeItVcbXSjdfiyjdNAcyGZ0JxsFWe2MsPPNxKTkSzg74
/NCQGyEXJEjQeufZ2HzL27S1V+ubvwY7LXwRNZ9jYIwE/UfNZ/8EHsl8QoAj7+Ih
TvFB4C3GC1PdcWM02vqg45RcoRbA3T4QteGbVd5m1pCkWLRfHLuZSb2JfCG92V8d
zO1nskaKwKVOeD3mxcVohiwOnmt8QDlfUvtXe7px6W5u1AfTK0E/THOiZcJCN//M
QogGtW1SVDfYPXoyGIUadnJGQmfHp4AePtcdv3svrxLXPJEclNBIqdViAhsNZusK
cnkEhRQBPJTsgP40dxAt1YOEG3hr7Xl+lfGZlLLztIZ++RTwEMbjqptHVLvcuui0
tR2n0RxPBoPxaEMwPB92ebKc9temUk5XtnlZlDPG79l3L7k4lwSmgmVQ8JpoiNuP
+VzTwX8ZkjTagOGDaCwyxgQroWR+6V+RgJTwM6QeUc2YsgwOvWsqKhuK9SikQf+r
MNscmSvVDVxms8ezoErnFsjJXr2Re0pT9SdjU4q0Biir5JpvXAOY7f/svI+cbGSn
nbB1NAKvcvb/rmzMTtnC8jdmZmsiqasVi3hJHByB17mPuGvTFkuApw4iQLUJ0s/k
g89LYmnseR1+cW19x1866BeY7yMtRx5V9jR/IDHg9XrWEmea0c3FP5EBiHsCX8eO
EnDiWYEf/flnbVjtkV1GMMn6hek4tFybF5cajOQV4RrohxogJ0XffXAGtVct6O06
wnvMuVLS7B27OvVd1btQ1ZFHhtE3p8UCzelzSfdtu+rhvc2/5sgCcB7cEjtPtp4d
FrI4V5U5v/x7zQ05H+WjiMwOFCSWj8RQttEmkf7K/prQbGFz6Wq9+7LrSqz+AI3u
cIQUeShw9S3gWCu0alBatqCMDJXKgL/c/6KwrvATSzPnoLod9m/Uy/hsYMMfd3+R
7KbA+TlzieF5uOHEkuwlq2T59QYQfdQmmGVRXBXb3XJAAYRma2w8klDSy1wGx8BR
c2jJxR62PQpd2CR4ygm/K+smSK3yhj9edaBDICdE5A5PTAc2Z4Ngs18+k0lkNuQP
iIyMYPRDtpf8rs26aeOuLOixDFovHUJKGb0VFzCmgUGa3H2l2H8aKrcsUyLZvCQH
48toSgc581TQOa9U7YPNL5ItpesLoYieNy7zf4YY5b8X0Zb0RSGDgkBoayvHs/ei
9ZjEyG4wlHfDNTwf6OIruz6OS7BOH1n6Wntefk1LdNdeM/ec8jHho7MALI/VWLud
R3NIp+i/Cv+TKSpodZzMUBoAri8eU117Nqi8FghEZHGtWHL8ogkRmkD8qciSwOl1
i37lSBsmOnKBMojgj6j3FPBWn/nGLiz7S3hewQ3RMiRCANEwUQI4ioWajkuIJKvn
hoiA7AOwAyFqxfWLpV6ULu0rMx8zutv4kMFXzA2Rgmd9Kyn9qoAoce2TMO9anii/
LfnyC1YIfVcF4p1QuXCfEF9qfN5QyDVCd3Xfr7RCiV4sPCIpEXmqEWWyLckuRjNq
NZUGM02tk7t4kJvfb5Xil6Y0E9N0OatR/zWmbjTYci4X7ZCteUL4wgjYDhaR1ZbV
DbadFLcrDXAEKEq2ROb7qTQoMjzfxoIhhgkB6CxGSQWGPRSoHdPuQuUWclJkNpVh
lxcrZBWYFGaoIvNaGAvkA9b+XvI4XBUq9vzVswHFh7+xM4oDYv4M4/f5wrk0eTNH
LPFWiT7p8cWFlmZlbrheQur2b52UjLiOTkUk4+rneDvYOqBhJydr1yG/YOWnOQEZ
Y8y0yIhD6tbHbu+Z0qveW7Z4PEJXQyfLQRkPf8oEFgsJKyG6WXIT9lzxnFarwWqL
qgrjGRuMS61yZP/xm/NgWEZazCWHnNyxxd0hUc13KcuVRQUqhPUYaW5b/wCYhMaW
9ygyVltWF6DCvjRngqlB07nLCjtAzt9jJQXAJnVNv1kKtcj6XEhMIpQNe7tKlLgN
4R449xz9kbnZKvG4ugQdd1DrLQH1Wb9uPeH3EfdDTe0d9Ij8LP1WwiSAKUuLTvT4
BAnL0VKSzAkRmMlfcgZH58/NP51sLbyPQ8OiAAjd4i2K75qlNS3kAsjwK6DxAOCg
l5IXt+64rgzPBwppAzCs7xz9hIV3O5f2gNB6YJinPnm752/INPkpA4ltZ63/exy9
YDG+C/xN9HzbEpFMXaClynQD4ZXYZJJOgJQM334dwfwLD2d1bB9JDajTL2DWm1qx
sy7iOBvkZulZ5onwrJE19d/svROvJVwd1wSW4F2RVdcMtFW3yW6zYQnAwr8h/0pe
v3Tvl6mC4F5AQepP/1s9J3vrFOAwTGfGYIqdbwMMcwnx1P2WlwrAnmU1kKtOlZJ5
Yd9x7yT+qXDrRR0tFGRf/OjMgov4gV7qMtD5DFhhzJNTvwV6Cqb2djYb+qL5S39S
yGvzYk+gatDi9ATjyLRkwfnvfTM0TtBoDF1PnkV08dZZcy2rAzOyTf2Y8mr4ZaDV
FRmHqJGpkG1N+Bs/pOr0saXGXDYCa6KrCpUwQkbUy7/hrvjuATa6nzABz6r7rGVy
mLxeoATA4LxozNQMa1AruepfZyFpDXbqU+Y4KHVOhc8rpbIrrekF6Rx9pl1WLs23
fLSnxKc2nFXbOZU2bO7Kr79Ug0VEA/ecDohilv6RsR1qCYZbG+czD+8nst2yI6qG
EIXe++/RMxJ6BJ1en2FJTFiQImylxH6TFoMD+ECV/rASUvG7zBLnUf059D2IEPYj
U0iF+lRNip7vBkOUFchRRuf/6sCR6RCu2g52nYGZWR/TGE746jp6+94E47t9c1hW
2kc3X98ngmWaQgV9miNtr/X8t+KoqUaj9Xc1AvjJR2/s6ivzXkTtbPaZCpIGdCMO
h7AOh+YBNa1G7JoBQukcjwl/oZY4gZZwn0VZWiAByzFHnPgHMWzq8N4tfj98i/3s
4Oo/mf0wTAKNluGbjMIjuiaQx2TI+VIqT3hj6dDYOrELqu/3ao7RNwbtcJ2eZuGR
ZsO2sPmYxu+AS7k7sSbCs5W6ciwKBOluzjzhh6K8SkGgtvwi1B+KhKJdT+Du2I2p
1SkSPiPH2Gr5URgbBbPU+UXgpkZ8f+VCoAHiNB6YaVG1KxFP95qSMVHMGeYnfCt0
iXn4RCPpKPKeA5WOJlbBzmCWV8cJ8htRQnRK0DLNlhagJR1NSv4clj7ZX2mS+44k
ESW94wCoEn6jPdmmZQSq7kjCd36GbCrZ+uhCqlqlyyA1G5CWTsPjILO8CDtbGE+S
CI66RN789P2fnYx0GHYipNyOUnXloQNU7uS2n987EmxtbqmPfs2iIJoFqoETiuW8
F7sSOOOtOMpY5PoyxfPcRh1Itg6EvLmh+sdUhC8Dr+Ba6bGV0uidWmOCiXt2UEAo
6qKitUwaR5taKXDQ9mo825sBo2D79LlRiyQbz0bZ5V85zLeh2G2Y33g8XWnwGNQM
9dcpC1rn3tq8PuBnUAlxeayoDezaO0QStrdpE+lxQ9txDWCQ+prxgwxbsqBk8iqk
wG/lh4tAsMq65s+6eQ1Rc2jS2iM7YPTawWgBkTouDD6aLGKgdx+n3xQ3siAzICto
F9hDcx/+e1h/aD003oGn22Gmvt+rLYo1TEQxzmDpAstXH/BVPA1DFpPoQd6Dbqfl
4xgknzjnIdpJFhap9zmIYKye3CXlYih9Cd6nP8UCtVSryNLiqaz14uqjJ5rVezi0
8sk6PPnGPqvGysK4/XstcJQj1ZeysfU8hxNHwALfxoJQCU2G8FhOk9AO+HvyfnKZ
Yx8z0RQMBUz1RysSyUtI0J6Lk//N6R3ra7PYxUXxKfN9o56XwThF0EZ+NxN2Gf2A
/+HYLuvCNVCew53O4nlBOkONnyorZ79R39FISwcRYQSwDMvVkd56D3WcYO6/vUCz
ZBdv/r/3am3SM6A1Gew+A5tePOiMxwqTNbPdf42XXRHcEkDNaUK6sjVsNWQEWdCz
yi2AFcwyXgZCTq4wefhQH8ebSJD2eWiNJpvL+qMBzAut+SZ3mUUzpM/jqu7tYYLN
KMLw/j10wYdtyCRJMVP0EgqoH64AWtKhc8wLHVzZ7S2KxX/shYjZSnYg0Zfk3xiX
JOZK+D/Ki3agyzVkNl+vSLuRMGGntpNHUHVmGjBHsz7Cs3ZGRuyTKRSN19cu09/U
Zp8PSA+xeEJyEvcAPOc10Jdk+n0KyTtodR2hXL2h3xbS64GK1sjEb+TK5nwJrWb4
lkkRbODR6jCqSsH+u1I9NaQ+aTJq08OFyJgLMj0IpcneHZYE7n7CtdGgDnHwF8ce
q2f6SqtV7nYhS42SJIniU56ibZMssm15L2M0DWasD2Wt2j79XiitOcdgk/D6ngau
57AqdENqqK11Zm43eTqglIUzwdakMSa9oLGUlZosJIduFp/wGAZtoqNrqdQkkbmc
eyiJnsouqjtvay9aBSEwM50W005wQRK+fehO5SeD/61VbzesaUL/u6X1CN0eMsG+
Y89Si4uaX61GyWHdAQlxhz6/uQXX+cnmcDYT3d8XTukQ052oKsuJnmZVDMbOkwdN
stYuf1Vr0V8JrDUhfFdGgqVFlcuw0ZoAMNDSywDQcT21y1CTGRjDjz9FS9IG/QMm
V5pYp5PhFUd7g1hJ63gfNouHUxGEWM1PPPh6uzYmYnBQRFZsEM8XdgQ1G5j0t3zm
q2GlDgiO3XsBlijYm9906pDMFL+N2BsdWOlNKp+aJrzJauWvP/iEwTru+HQI0Q8V
ZDsgPPc8ZiK445eX9O0PFeKpC8YRbRXeBHa5YKQyVV+yYH62wTromGmWXHmyDPwh
Cj9eSFu5cDND/FPyLeayz2N68Kw2uywUbMOoif+8J5d8biQgU4LP/78A2GKy2IY+
SKA7Y+/CGK/IL3lYSDrwqtaYNU/mh252WlW2FEt+1mmxVGvisDg/RuxFRHM8VUom
N4KMhlrUxyX3IaLpfufdh0wXYFs7J5McRUGhEzGh0E/sMf1Pzo0H4e8MZklUTZAG
rEInJgI2Gj+vGjxVyBz82gcDN4BYe4wvdJYfK0gbMXeDXgzs7MM7y1tuXYYzl0aE
W4NSOO7xfDIsPAer0LiGLAPCV3+/KB7jb6oZnpC2F1B4EDEGjKa8CADugFm7nzCF
R9P0uUL7gjW++a6ZCG+mNBGrFSzwv0/+2M1voTGqPSl23vLCAlo8wGX5GY4JKdKL
eS1+sokrxtWqoVJOnXyR0B3NW8db8/MeqShN7DqpRc72dGc+KwQQYVgzmE2huyyQ
c2DI2rjUOQpzyjvbLfXrbZjDkaxpHqFGIoClGcZ6Fm9kT90KSvtiKkVEU9/VP19b
4W8xt8OLjbu9HxH8RaKordqbnRejY2bjs6PT3vnqYQ+e2Tb0Ulm8iE7lp4OthLGG
tG7mk2T+RYkdT+VXw2DwvQNBhPTUMJK8lqtFskCvmAP+9EEOSRC8Az8e2vYAq3Fx
VnE7vjMviJGyimBGAjY+2rRvW+M26vIkBHvv4FigVtkCH5N9YV9lJ85UhclrMLyl
/SO4Dynh3F6bM5XCq3ToYZsrjmimN4BPm7aK7BiyPMHNE49jmXuluH43m0AB8f44
h+xhnUFx/GWh+Mnq9atFJt2MOwDxJpDme+QPczYINPE+BZZ88rylMprQYr0jA2W4
/F/dkB+EGB50Uc3lQR1hxHal6yuz6E4nUH80kUgAglFFRBSzoIoBQUiiEe28OGhP
75wqxinU6ql7XuUwaz+XRwfDJCOeCOEBghOThE3JFBMJLg4W/udCcWZ5iaBb5Y8h
Nja1ThdHK4Q5J7bZlsKoPFppQO4qPKzJXz2Y8YSbLJkfL5Z3lAw33tmZWVMkLRQz
QSM3ClB036dmap5FkL408V0HrlGAMwnxJbO+NZbc+b9Dp52kVi86m7JEaukJQds4
4Ew2TCdKVToGBGZEprfwTbJoY9xaXo+LXqw1S93Xqo5srDPWtkRVUkZQKhUEDsYB
X6fO7Q/6KOoGayv06GhS8N96HPy0o3zS9pQV9sHajS+plxYUGI+4+GgpzptMsIvi
iMtzQopVCuu9Ddj1/HdYvTuaaLPLfWnSL0+cAFlp4GrcP5EHx7MlhuOzx2p+qNdv
jAjNsSNeoIlA7OjUttFBJzf+Pft6hD+C0XkkmWo1J+/3XF+zsb5tAj5ZecBHIYOY
80bhsHODHiretzboG7lsmkvJB/62hhwfAPmFo7Tea5QWla3roXVGam+u5g6kFfO0
JW49cgqboMrWXK64F7NQ1fsmkuhBfT6eeqNgIrJu2rCxTUIJ76r0j5FzEeG/IznD
OgOgdCBrE0XwpaYOaGfPtRzZYEXSb1DyOm8j2X4WEyf6kxXXIV09jR5SD0+YX139
/dYiCvTbFgOE2khgM04mWCPDbmEtf7m38A93K/VgIAF1WIRpElNg09cEbBBYhuJ7
D5/mkAFBvvW9HLwW6w5SwdFkwu0Zv2P7fJkgOW47zZp6IYAgImQeonPp33PIncoa
SeOJPNfcu7KiI8rnhbPKxQ0yolidTcq0jOyxZaMBJywsNCACZEcWB3tJ2BxsWQny
yt1wjnKWJ6BnMZPzNqSsRdMb1teGKv6WXaYgmNa7opuI1J96sh9ApUIUTeiaQ969
rcpjPsaGhjwC3tzVecuaDmgvNc10XD37PeeHGj+sJ6Uxfi+ZNUhUt+cAYbqv/RZM
8gycgAagEesWuaqLSCz+HoS0Mdeyh1mDN0RNGktjhXlpDI8uXQWtJslt94j5HCsX
qLOsCFyBW0RrZiCEIycf2QJbkfW2wdsvJ9J1YZ8OA730FvtfUAbpoFBiiLTURzr0
amn+oFJiN31zpcvbVl9frXHBG1LsmQRF+wkEtuf0VlCkLAu2Meq8FUx2sAXk1QhF
RxzobHHyVid79TgUjs9OgG1WXm873EtDW/OSoFkXZWIYGTiGxT796UzhXtMNUVp6
qED2ghcuCGLquhRt0j9gBRLAbSwj/o40nuL91qBm/JFe6GXf/rO9kyRF61iGdyen
m5JrpzesAFRkWUUyzoI5Y0zcI6mIfBZgzhCuAYwpUEOq2eOObNW+ZQw+jbFsSbFJ
Oty7Uvf2K8NHva+K0SVZXtx3B7zA8JpntR/iW8TG1RzwIH/Jl0tKqOHdin8hEfDO
41ieS0lRie/IpRGks6mYZNOt+Eu6UE1FCzPrqe8XKB94NTqIdVh/B/GzQhdcFrB9
bbatSAX6L+574tykxH7mIkLGHfKiuEdtO1MazTSLqm7aX0PWDWyEHjyrtit6JQ5/
RnUOfOM3B+pNdxzWjH3/r2b3PE3Qg7ryDQXTo+4OX4BHXV5hvKsM5QR9+ZsiGtdW
HlUA85zXNvx4irvA6Ihcrwfea7idyhSzL1uh9iFWCvxMo7xE5ObgM40RT4U9OOkR
vBBotb+HSJEDewCfP8/9k630AgYXQTXt2msQGkg1t0LmQnsC+5F40Xu8CcqbLxmH
V16CK2upIqrPCCVLQuD/nPq/hu4fAckRKkJjFu3bpBoLsrHfZjOsB/uzDxxka5qf
wnNGcWNMNpNZuF+gOo1WJGpJD/fj65otd7RoHgpgbP9fYBuDe6T7xLEYlp5GtVZI
IwmAAa4kE+Nt0Yj1hyQMIK4Dxi7OG/6XyNKnBpFdSR36+e25kEmH5caMHLTZoFfi
i/IrY57IRBTCDFIUTW7ZigNrUL0/mkZOWWkR+ovsG2aylL1A282krv9XuGKo9QJU
fBNnzF3EbdPEAxXAh0mlpyCcKjdT1pW49Pu/n9jPwPZKieh4WkecUMUJYZqkwR7w
xQfSYIIYzxh8CLHg0+dtqAlLWkZMcauw/89Eiffx2+0xpXoeHv+q6NIJF3B9cKrE
dbIouBK1OAPXDxVQ90oG7XJyqwFhJRtMCuEcGlpmkksnEFl61Ikld93zeFrMUMUc
mrygi7gW6u/RWXk6N6U4RUbk/Nb6xvYQbHtRIb8o2zB7zkKc6g7kHM21PG93tsva
BdhmZ7qKtR5RL7GVO3ml3wY6Hq6nB/VxVlOsCfFWk3vuwRUSxoPWUm6t+6Mouph1
+/nedzhjBGxRBLCnUi62L88eTzBCp48FPkzCXLXGGmX8eHXjK/cnm5FFshmiHvWu
0XD2mxmG07QzSdrT9mkAx8+xVgDHQmKcysWOAZ2+AiQoHiclVWXJ80gH9lnmKbax
IU2bV/AlAhmXWbSpCBjS5PZdGD71y6ndp8eGEmCzck6TsTecvhVux0VSKrKSoYxq
fCPcfiulW0dg/5D2J7j+iW0u4kgo7EDOQ/HoQmEAkJ4+scdI7Od6Jj7z9KdqMZib
sAxor4zZG+TZPcHRB4bET1ZK46aI9h7V4ztmDHr3eTB7cPTilR4QREhcms+WvUpD
DjQJ3g/Tj7sugGrSwe6+9DVMjaSBw9VL2BTa9BW84NneMsghv56+PhhWgGstASMt
F/Or5XkGVtp24rgaGx2M+lhGvwicTQVo/InP+J/fNlKJvyUCfNZ3rj6q8lD7ngAV
L+pl4OhvBlJGKYMnjS96kricvN3v34VzyAkpFObk5e5Fbv1Phm8CLgpdGPrgTfgM
O8LkjMkFCIxwrXRlYX+V7Qz2KWw9MuhcQsocGwoHAR1Q3m83zRIrxRSOEcFrQWS9
T/EMUA34zLfA6uHiaihy6EexWjUC86ds4qbfZRH/nLdChpzZUFBCRH9P+ahL2a9b
1yyni+Ld4Od3rF9w48cPToGqL2SieIdKPOpieEtH40fLvyKis8N2l6+Mv0egEuFv
nXw5pEA3xb7EiDsP79327UiE4MV6KxQOgoZ+yCmr3QJKs51KkADbFyUsunRltYW6
LQAszavvEHi2VrPWxCvFpW+Afb3JTyBKXX6ZmFONw0LD6eAyZy/9HYVD3PKf/MOm
5N3xV25JHqM9sz7gmgmXQ1HREOhsbQPwzZtPrXZAOptEOnFc/damAQ3h3pI0NC5B
JeIBvIzpi9nzJeE8zhn8hJrJybRdQ3WHsW6TYqdFl9LV0MEiUTW2pzrnjTm/V3Wn
qKxMYHxDOi492l/Anh6tFZ2ctXb3IxR2cUUSoGdr6UpmQ1waFVnmDsvpceWvXDsq
iGBCIDyN53HX2KpAdClwLnycembpvj3AQm9E0g9bR+BH2Z4HJZWnbyb49+jDhO+q
TtttB3XWZ0hhe6RVlZ4OvJIOviVLFRKuARMxWlsmh6yF2N19ZLIVAJvd5ne1Lj8d
2aIhn7Gg+cilKIoxCerxp4h+WWn8Tl5Jm73K/qmPZ4Gct2/mCwj9fpZ/l3ZulGxY
qRUZkpZ3v0qosko4pucXlCz3ts905sw1rXvnUX4FnpsyYrldj9klrzBx6V5ruSxV
r+xZGrAIie0a/aCKAc6fnKBw4FjOPg2C3VgOOvMSoTfAUw9R8six7iiFJh7cIskY
Upg2R+EC0WpjAaOibRDJ45yx3ER9YPhzicfxu1bMk31VDOQkGj2WClM4EHXBH90E
o2lMRyIfVY3B/hL746+ZK2nlP3GKomStam27nTDjANeXViBcxABBhg1ofGFjQtjG
leWKOz4MDPNL5COwzAlLotve8NOD4nljNA59WJZnOcy689VUc8ZR8kDJ+8FMkDQ+
hASVcrQcUKnowyYKTZ08RP1NfVOLTGlk0R4CytzozNnF5QsOJqCF5vIBssJvfSPg
Zp/Pl+a0hG72oiu9fdp2vqtqulFpT1evUE9IqIKmjKln2l6+qoZXZ6HP3TxYQcaT
RFlPiuCuZkb922RGlRSEohsnUuvOie87m02DwCSrpq6k0CKDYCUsmXaQc7FC18oU
Li4Kap93J+8L44WAzP9NVBVffiNc+FMvY4aXEi5YE5SZOGuml/rJwQ4wdRZlsgtL
w88xcZa8TYB8Iskmtjw5rKq9l+KZXwCup5U0/P2br8d8id+dGDJ8yQ9ViOqmyD4r
2GOAFkETNfyfrVxNFavmlmhGDtyYNzXKInQt6+yiOKf+BaXhkjTtfD6lKbnGC/Sh
P0gZ2SHnfXca5Q34zaA1q6/L8fCTicHaT5wEvQNgDmOUzijvXO/KKoo3/cSPlZNH
uBP3js9V2Cu4V3NPxEhfQEVSIIGogAuck3sc6vpm0lmww2r/oBlOcpBKY6kM+Vlx
0Uvx0F/gGMCA93dYNHX9yOIpqw/8OpZ+jFcHzecWQigCrngvVB3OrR0JGs4sVnvh
W8EfKgK912eN3uCz4lQxD9yCGUngsKZY2nP09yO5cOctDcNXDkDsizlLBHDpoZdK
kdLSK+crFrcIuIELd8RGI6XUWb0wXlhTGxtb2ueOemj3sm+Rbbmg6gMuRdstRlWL
2KaoaUVHj8b2krybUTo8B+h2/vqHSB2/RR7uZtc6hYclAijMSJgWjO5OMRQAHEp4
l4YKl4+2rslHcHz0wO7ywJLvui8sq6iab1hIhncu41NXWRy5j9C3l2GS+OJm4vKk
oLU0OZU/iDlZnSuFKyhk40LYebXRqmd+cVAgYQlnfbFSpEklinqxROHzYsP16zlR
0NJGm5mz/Ls/H2hYHm8PD4ihmH28IxHyJgWJVcjhEOKsY7KmmSOHV4juOypVyg9w
IVW54C488ZA0skr7Ng3oqM/5nGDkzBUhzesGhd9ZVdv79wTgOoKnZhPAop3M4x/t
ikoFvBZrSLBJmCefSCn4rT/QTZ/O8qDrjeLFoIFAfs15kltMSAhQwCg5RneikRtm
EFzN7x7YQN3bbRc86iww6USHb5b6m1aLZX+Ln5eMJRx+r01vAm1nLKkvBbjTX9pG
KyTDu+Vhb3LlT6aZENn2CryPaTBwfMyh7ZrVxwZvZCBDuY1c5k5dVgMFH3C3h4LF
+HDN4+RRPx7E2onZDCgO6Jmg+tAh4/8HKZix6STc7Z7x0l+A1Xt2/P79Tu+D/7+w
2hDSLChNQIkyE1zJnYUXPnp046omPVhSYaycyya7r6R6mx4gZC0UE8p7ya7ICW9Y
+LEvdip+ArBG9EO8PqbgQlKtz3L715FCa1XNhgEyBNmN7FKsYcT2JBFVdnEjPtIX
eMQGyvmThOpVij5EboD/Y1Ty9xe2bnN2eGaPJlYP+3kGpaoICm9vizF+noptCuNq
CORJ6SSLx1tQdKiJiMQCMycqL3yejpKv2+1XJfjWbtx2LDS7Loq9K3SVEkD6tbvv
nrVlUk8SMw+XDJqlolL/2iT4tiBVaF1N0nDjet7HboGuMGWtoONx71SwndFY0fI1
9unsR/7locB/Y+i78XOU+ZErlU8gMOVYLuh+hF+BMGcsqANQRiunT7N0NPUEn9Gl
7wZu4Y9Hb9XE9FrgDiHKK/CSGSPNdb7LJQP3HbGirGY1lIk8FNHj1z3t1DNpK0b7
w0CPX5aA15sF3Y5E/Xmr5WDIJnxtffcwOBDqa7cLUiJeHWKA59Uwk7C/7K4NWjAo
yD8h12VRlywlZfzYLFZGvzDJoY96Urz+C/qHBralNzBI7reNJQbg8boJJuAEmAaL
cStsHjvgGGlzBUc2maKFnNkrOjugJ9ag3SXkFQgp0bEsoMxUx/fBUobDVGVax3yz
cJChbpcQHLpOjPsEx+or0DS+L0+JE1OnWEt3i+qnhYPBy/hPo3O2xvSF3Bgyp8V8
dowm5Hfq/uzAxwdGjAcHs/JOynhLttzadF/F4sJTADlL5YRpvmogntAmIlo/fJP3
J9CqT8H9f+u+MhD83CgEnFs19hxLl7HB63QTzQ8Z6KHybSiX6gwmVnu1KeBMbZVr
sMV39pQUUIgAiI7j32k/3NOsQwE1V8EBSGv0t2lOHI6BM50Z38hsRgWzsO2XUDpg
reCG09KihYmjrQ+P/xvtxMTKXt693YrqQPZHorpnNdDCcs04Vp2LSUdNfyK5Wfpm
U3H7zYhUOzoreJ/tt8lhR4hj191cN3hF/lRB9T7X4pCBEsUgIPb+Iqa64+rNA/7s
XWqPsWd9uW6+PmeEL2c16Es65Dd6xL1Q6pgGmP/YEhubUCg2tLMmOR0tZXwQKpB/
UokGe54/3OYGsDWGivM9NGwVmAYMBWqIxZtJhuJP4kfm+2+xoowCEdvvni3DA4ZT
ZgMNjj5eQn8DSFOC83sz+xOwmlZcpb/OUJ0YgFJzQDx3+kIEaYqMC2WBnAzbH1KJ
yWeqYd+SlETjFln0aivNqZxrnBQWs5dDdRbrSV/VpGIzc+mT0gDDU1Sv/+0mz/hG
Qn1vDbAGdjLVjTECaI2HkEv/r5Iju8fo8Z9EZdO90UHAJ591i9zic82jQL/dvwyz
6Kn47ymx6JB1M+iB9l2jE2hKkD42zgKL+Tv09vnm1cRz8/WiHa9C+u0ARpWXwNi4
IyqjLANKKO2O2K/VrmH5RpfvzDAGHWXObButGXWR9DGEzPtroQ3N+lj1zcrSWxFb
CxEkAGST2rePMbzA16I3XWSrJwQbQU5zvkW5R3u5kylA98UfXV+fIjv/abQG1vMQ
+OVu7h7mgRojthtjExdWMzzPl61cGGg6oaIymt4hXeJh98U/4RvYOr3VtNRwsB3z
SdpECIIQBeTeiIX8y3SNYk55IZrARv7yzfzhFMo25eURYrH6MSbkXjG441fzk6LW
ZIV6fYT5hiYUSNt7lvlJt6ChjvALscXfQL10pu+FAnnNvSxt+M32sTMyntKiDPIt
0QrSY9GUYj08qF74Z/aFWHKTFKFBA4t0xnindKb28cWGLNaJjlyedaG5mybk1CUU
59kTTM8no8ZarIAVEL8tsb5yCpPZgsGM6tCpnt63ej7eY9vaWUTzGqANREX78Bda
qzPPQEZPwg/uRc4xMSUCRD/5+72NwCg6WY1pdqXgPNYeJhMCcj3Z9mrop2/OdgWr
GX7ew9mmbwvxXPUxiz61OJAI2VyAhF7wKOjMH+OxoQWKohm0iCmZOlXvC6HfLkLP
6zt8pHqiSMHwB7aPYlDHRLU2TZDO8YiFtN9ETVMYmGQO1669Z9kukRojkCat/rld
P2tXdY8a+5A8osb11UMc8cx1IEPteYoS8O8XngMAI2YsebchbEQIlOAO2v5wTw7c
E74f82bF8deQ/SjV0kix04n/t81G5tTUGk3Nq9QcfVtZBWZPtTgtxPzFTwRhWlen
/qMIiYwNUKqUHATK+VB5i96lQwBFfVi/l1rI7t65ET8bJc6JX4cf+Rz6VK2mSokx
69+GQ4BFa1wXcuRWRmbpnnd/356AWA9SSSmXXvwEMg8nl+0LaRlKT8ziTugVW7dk
mtsJ/clb8hOKcLNQptY3qqf5+1TBXVZYp28wWD3AtI6/KmqA1xulC7vVaCV6x7s5
XS7gYz+1xMb20nxJE9hIi2I4NPF+DhvLHyUaoWtYDgIYMxLF1J815b1kIrUd6dc3
RtMtKe9UwzDp04QYFKc3lxUci1y3lN3c6TeIp1MsFaA/8z9N3PnvdWYzZmLoL2TZ
5HJoqLgg3AWNd3sGCCC4tyThlfZgSg519xs3bC1FEF5mFUtZ5+n7Irc3rGHWWFKR
1iIewifEpqOtYMoYa2coSH8fdECyZISaY+7nanuLhNQphUSTIknNXj/2RgtOVGiH
LscxHjetp2MUvsppafFdYSYVAV5kC8L0e777MwyHXN2cVhhhOskTxuDKHqplWZFZ
7p75jyKn1tOOZGA+fEj4eAXvP/qhIhKuEbzGv6SX6DSkYk3g26UYertvaP8sXK/4
vTjeBJtcLQh44LpN3d11OWh0e5Mqm1sxJdWN8Wua12fH9UOiMes15hT5mptGDYUD
1YwT60LmHePG4j6ME0+Rg/7eSF6iVg5wusvHIE3D0g94JKkKDz0sEEAsQo+XV9eT
byQdtG33VkmkrJDO34KPON1eJeSipxlZK0CVx5rQFI8jRsLi0bAyLCT5KF3ckM61
1KjrPSCPYpABpsSxDCP3mo/LmCpwM4UogjFrmGIGDg6ASkhCPvWoZvNC6gYxF6VJ
4hXsa5bYZTGWooNTP30QiBHFVPNNCSMgvChziDFHaJzxW8eTlkE4AjIVD2fXW31K
fAZBGG3+Tr76GPOYgwked/1Wa9VH7xv9SrHGhJ8OcYkX20TwjbTiFrq37e7L08zu
0K5FM93GhVIazzMX4sprY7DVm0iUX3ogfNntl4Tmi1CaSaNUEyVhLu1zFtXjuuj/
XgX3fvRcn/eie79D/ZoDJIIRJbp5SZsDYmOxuodtCAChxlOSciuXgvu4hwNtCjQp
xtnxEz0sGT100KcpthrmLo3QKRPg3X4y8OtqVMyzRfvhVaH8e9hJke5fT1DwXAv4
uQR1krjajxitysUZFwq6RzMfMO2X1YZW05aQVKjgOZnFUsrTYw/v2Ziv+zoS79Gu
/eqD3ngZO7xe24YXyS2o44U+QlZ03F6w4R5YY+/K5bQgCTY9L3Pn2NMKRyI2vFr5
05WGCL1zJrBbZI7N0HiUJzSbtMx2B2h3DxdgCc4sQ2VkWTtIp4TJTPU4shoDDuz9
jZuc6iL0X4hPXQpLbiq6uuOOuECAUNGRHaHjCc9DxTZU+YN7/HgPhoyNvYWmBi9O
tbNamp+L8npO7jRu4ofwBZ3rOSf9jyVVGUn+EMZHqWhvlUyMC4+/8pmqvkBNs3U7
kkFf8fWQi5962IbsGsFtOhP2R7HCP2YlWhPuuwHWTIDEBuyRs9tUkwJJaemBg02m
EjJdoByTQBm/dzxd0Ss55y85NOK4NVSTEIOEIgq+61kKDmqa2Pu6rlnMI8hCNoz9
PCr4UqC73I5iDwkeTdtCnxgrtiYSrDXQIa4RXePfZx8XCgKkz3Lj9V1nY3rwHHlL
LJd0j2I/Qj+cnzgRXwlMYtuo5/Sf/ayMtvNuta7FCqQvhJ2PIBFziINAAdEeQN6a
rtKT+l+EmNzRlKKJpDHXj2K32Z8Pck0DXCLGoWJ2JF1T0C0CIXknQMIxHoXH8/A9
9LX2LxmjRgJ/Ii2rH4eeip7s7dvSNfO9SPdStuSKjAj6Dg5H3ny0cEPSSEE+X4PU
bO0v2fkxJBfbUK/5TXWLvSchuClSV+XzzIp12NDCx+H0jCfrfpss+arloZYTJz0v
1A2tdF7YKyTP1AG0tdPCeH+GPd85tsLVYQ+rbUGUMZck9eVYGqQAzNT4bkY1oeO1
JrO2i6KUaC/wCgxTZDeC2+cRFMdYdUQMsQkEF7zYkziYIBxF4wQYbHjaQAClEbom
Ve1Fg3YZ89R1Ot2Yik3KlEAgrHjeD6koB9PWzLLHL/mKh1qxyUVE+RsBlYTPGLHu
jl3wN0m0eqeQW98sX7aaLw9y7Zg9IqaC7GvrsCMZlH6E972D+1vxFC+w8nQ4jJZq
6pYZA1+qyexJNGPeVHenmQEQzw3hw6Mn6pD2F6yfnjtJRFwMc3YFZ81/EtPzpIRF
vJiMbcS4wYPM461DSW8Ayvn+SPP019peh4int5kL1CpfObBxNIt5tNtJ9BFsF5wH
MsXLQVhTvoPPzqhRrKhd6R3bMK8y53wIzuAgC1jmK0T65v7KujhemFXy4aHdswyB
YPle3d2dspsQDsCAPP5vbkvLpwsQ//dPKelelfOKG+zlPHrszq5YTAPcxbMigqVu
EPlsmIdVJaoC8CBajkfTlw9PGSMZDmHhaktfkvfLo0vNrdRLBgebvnDKtvuJD6Dm
Sja+clMR74clEgWBehs4bF6o5c65LQsxJ2YPgZ9zTZT/fVWys4xeTZwFOb9wqB3Y
ZjgkDK9IuL3/CaoL1VfvYBFAZ7uXN/plouqLfPVrqmhjj6OQm7KDdKqgbF4HoDHs
uCOhdxJ98XZTJ+wDnNzPTdV5KbFIGFMkF/SqotfrvpGJw5ESuRxAAnEODVJu8L/a
UnYEQDMc0Q0UjDXHJPDrH4E0gA0Tbx09UsLe+tl9cSlRdlZjdTFeBvrXLyuR+1GR
TD1LkqJlFDu4j9zRMHTy/fRadWu4Kd7E6C9sAy4VJp6nbRI08wdG2NZpdc9cm8Rg
QEPxfxVyBhpBz7r4SycipRUemErDHpDL/sHtdGsBkSycFNOGc/Z99usQqLc3zgWc
kqfCwdpIgmAB46o2PZopp4mD1xlJnZh71KNdquu4cR1Mbl0B/OJZSKEIX0mG4+Ud
VQOmH2YDcRa7sDHrJoKBON8MSqlfmgxcZa5ERuYXuse81aR8Riisha4PT3sSpZTt
K1vYmDBH6fv0N6dDC61li67U4pW47+Wiovk4J7Y1gQSGi3nq3xlzN/xR4ap0OlXM
IQBzCYVyBb29uA732K9JX4nY5qQAQaaAmgSCzy+b3k17SsgTCV0WXgsDMMh2W1j1
sj/Olsq9JhsJaKmRWNaxJvFoAOXV34KiSy+u9N1b7y/uP8+xUakwLaQ/pDLzDd2X
aFiM7orjubjw/nMhLNgDY0bP9BBn7RaeZM2V9P8OOEa+ztVvZEEW1MXIPxEF0kmI
yxe+u5RGADsLK6XLCdFwy5K2PTHP8m5prnFslaIxyPakCXN52s2Cka4UEaECa9N0
L4GgXVrD99ME1I8XzQuormn/6b3+8Zv4FpXkN5ESRnSFT8RlV4gUUoCB7bchb304
9DjjS6/gcOidcFGamBW1hgEAGwJPUzymxtof7E27REAZt9zUNx5plutJsG2M6yCi
x1nxR6w0trVR30NrGuu/UNcBQdGrVg/5qBOoIFJ87IMZDnlbWzgBW9Dhqi+MCNI9
DFbP/j9xAeRkbgMXkHEznUdeV+lWacRFY8TB7cx8lflEx+vJ/TfSMo7e1jK28nH8
mfm/MVuSR89hbvf+SungtHmXlg0ECppi+Ad4J9Z4c1RoLkKHau9VzzQ97gX9Qut/
l2BOBndpJbdZr30KWHLk0VvZu1ngTvX8GCgTWowkBFgMoBTzT8UbdypixJCWPvuZ
u1e9mUnF4iO9mOjHwdMOMICLgH+9jWJyWfu+yx5oNq4saQtOrVQFGq3KSZ/bZT3n
dynIz3GHfEsAyex6Rjvo6EwFtocpZ9AQ6S3N5YKCzpa/crilPQ5sVCcvdkWdjaDQ
jQr7Syq20KUS0Yt6Nfyb7wUCUWucAXoMRysx/Y/edbS3BKggNOYXD8Hx3DAdpIwe
cuCxlKeeoPY08/CITbUd6WR/KoLuzsu+rPStEqwe8toYO3xl4LeORpJHGpt6YOsq
Zn5UzX6qwrm9wtW/rXTXAaJAN91AukqIcEC5vEseEsAOntLaTizDYmgAsB7MLa7Y
tR/pCffB6HwreF9D6RZ7cdJFx4BQ7iQ5fclljxDbleFvVKp8EPR3NOW6wbUvAU4B
/tRapwgUuEjQt8ZHWN3WLpZiNVnpwFqWxO42f6Afy4d5Pumsaol3sTGyq1tKJ0Td
u4sn8XQzA743ylZ1FYxRuRSHKOrnNmAe9Ubk0jNO212O1sBt4hC0O593ppAFaNu9
zvjPF618nkR/a7MnnuciaXxXZw5c6qaeSAZn/6oFjl2eshsx/yi/PxmHPqAINYr9
g6kA9EFuzvK8jNe1drJwfLP9o5nPIkNrPYpcKT34qgsOfyiOkOg5IUzmoZec0ndk
7S6SM5B+nmBSEjDcjmQNSC2un+6etZzQxz78IaaLMvCShitG0D+uwV5AAn4R76Wk
necZxxrCFuTrCRDRuo8pJ8ft7ATgo0Xb27OoZAUWcw+yMDKsoFtJCOo0z0ZhiqS/
HeNHVpBK0VKnmK1OTrLfjF7vLx5ykfndpt6sUdIWYkREE4Hj42r4pRiAk0/+VSs1
BQ/MRWbczv+KvJaOApUoK51VYr0uKk1/ny+pioTyq1RDWLD4uA7AdJM3vRqO6GT9
1XzVWP7ZqcXIf7AWczXhyHUXblLISLLDFjv22p2nsEvNa6OzA1a0Z2lFXbvBc2pa
lpa0+ODI5yDWu24qSGxyA2zcMU3nVfHnNOkRLfJUI0BwKH1/Dkp0hjQvxfRMWrI0
Xj8WklX4toih9QBoSCvhhokvUrQCdhMe9VKLtCbd+gSUEmZB6hjWI+sP38F8fLsi
PE0oF3O5K9++NJaAVTnG+BGChczHr3n/RYTvKXFkw3yIJdARU+N6/pVnOo+DjLTW
3T4rtuLRlSy1AZoGN55ih/OnX/PaoE7KkU5TJ0wBD1X0A12bo36wqpwf4BJ0CVYy
jByfTkM7tpUWAg4ElEA2IrlZZLblqT5orR+9wszSoVH6Qd1B1pR4y34+MCggfM1A
3VbfApbyQFvGgJZu7r3hx8xskmOwzAk3xCjJvJXhxu5HX1Ry79FJW9JV1m03dSKZ
t/PLUkWHmTlg2EDhAqg1XSWXN2oFGNHrrz4VT8HHhA1Jd1fYpu0Sry5u59XR8js0
kmH5eLm/vZnPBbu94sG5QgxoiPDXF15mxB9PC+F7ookWoisJ/XGjgCFPQEWHztp9
PGQGShDQWl1k+sIS87rgPvMpfi1xIWxXOzSLzHyVA26wnuYCStCvXV478r5dRhQo
NKlVxqeNe8WLeO138bUqL4CS8kiTdDW33bn1dREXYq97508ChZaJBZj1xs3+FFIF
wGk2ELqoNnZXVAy7K+o+06nakuh1Ze3c6kE8NITYYZITxFMey++2NTAu+UIHRznN
maRiMGyNFESeMHZV3na0mzaqe4PvuXVmrM2lxPyRKB286QBhoCYXzlrdc+l1ICn6
XmaFCBU9KCF45as8W9tXIl9A+hnhsFE4HEmN4IbDh10L9tqjIFlL3J34NmQZfB3T
5EzFAIRdF1732mtE/LgnwWgOHvuP/bMAHOEgbAUc8xySaWsH3A3Bl58Nnlz+3UgC
q5/DNZQrpLsLLu9uBMCYrkUHi0SKhwX91TLYaUrhAqaUnbYtoTYR5Wl6s0whiGGp
ta5wzYKC1zjkHjURWDigHwfSISnmirxcX5uc+UnaXIbchUPPFUrAdGbwIZpgEWjt
J89SeIIJmFc0puLlClLA18kEkwSbZc2VhMcZjKdvlP/sx6yoCW38aTgrBSkD9zLR
OFM4QXxSmQv/eIt8rfGH7qObX3di+bUEYiSbEkHscDAhrUPh2rtLZNwtzT66zma2
MCRtXHfxGAp4B48c0HPP8A35E6WzWoJiGc5RxWQ2YwfW42muTxeHzVXsBcYO95M1
AUm+zWPuNSAplgj1QJ4bK8PyfbgRX3Rgh2GO4JlIePdLRV4Hc4/daRHmfJicLg+O
mjGdyyL+eKXYU69Gsk3MnljgJ4Y7bo7BSKJav99/pxCxqjdWaQZ1UISzdtD4xjtO
1wXpNF2GEATI8aLCXETPncG8U+/Vol61ur3/EIp3F88Msrng1KFRUCb3hWDWdpXv
5VHZd5SzmNLVot6JghXl3UEWCY9m4iMiwjmtxMDRzliQiGATXz4755Yo/Dr4PhXu
3jFpwzLJJMe1QUeMH8+co7VVwjhX3y9MWiNZbIgKvD/SO3NNzhN9eMZiIhMAMmIS
6QkNy8i5XMySJyC0pprbhEJ9IwCG7fnIEZ9o5GtKaTuLDXKwp7AnsB95NtXAH5dH
k3x+MhZntyfKOXSInpGCleRKNdf7ahwR+m2VJppC8f7RdjLZSIHMTcPRf+9VC9cS
JLyVFxSdxSmw8Daop42Mws/wpfXO4ovqtA8P+5gtzpVbqrlymUR9+Aapr3j6iD3C
BL2l5asZVsUi15cCgalmGg/P5A0+f6OmJOaIgCqRof0EzwmOM21vXRWKarDL4QqB
JoZUI0PUslcPgInPl2OfHBqgyiXuq3v5g7KzAY/VI019dDgxOJuXF5Z0bL/2GvO9
ZAAxM2SSvND06ASNdArGsqfJB6WKcLiBdo1PUgcFLtF+Lr/4zBpgN68qLPekqaVo
+LrTnP3Ex27+g3NgrSfgwvJYjq3nDlfmUY6asckjdmnv/QUlJQK/DWoXkShZmzKX
HXj2Po7FVMZK26S1SNtLWgmoaYmwDOxR3W9AV2GENc0uvturfTyA7CEoa/QBrtAf
Zi7eVCmqEOoOvaMudEKjoOJkMH5lOJ3bwEpnH4ho79SyjLcJkKErXfYBqk/4jc2q
4KSc1lwUbPv3koiZoXi4E5w/unrzGjB39YYaSkX7nZINxZS5jwSuYQdAcFdLIc3M
QxhaUfkJ3Rw4IWjQvsxNX1BZDgNkOLBMqoMZql24sOnlh0cJLhVpShGXo3zfncgh
i0jvhCHW0vHHGQ2MFS90KBoTBdPKbjdZDnqDvn82ZKkoZnHFOWxFIvlcoY4MDh0E
OCfobJMAuEshqHKHjLbrd15uLU8eObQ47pgiyrsV6sTbqGEvFq/s7yZKssBPe3Zz
kPRt6sgo76GIE86+5HDoZRliEO91REF1AxLYdfJji8sS0NWckVqlzNhqAQWJ0AnJ
y6Dw4lO2+r+6vsn/lVuTPNuM/7snaPVqanJs6GX7q1A0CIB72jFI6WXywuOBkmrp
ISQDfhNW3wOHfqIa58ytBiL7FYQNmt3jkE82+7ODff7NqHOQ41cSrQEo4jPsYuTf
lNd5uzyIwZDXUqDPbf/HwyuIHV6D4HCBcflksDbuSNGg7MgO7UL/c7JtnIHNznoE
s9qH54VxZwBFAgC2HtU1PuESmGFYOnqPNVyL0kX7wmeirYRSGuqLzZl/7+lMgZv5
wHjqupK3ntAmcAnHNHZPH+K/1FyDTZkYvLX1fgn/DGEfqjq7Ay30EziTPsu+Lcce
NSqPtxnKOCCdAOzni7bqrUcuvm0Z/fknQoedYqI7kZZFZ5uIHtQs0f6L+8n3VfQ5
LJu/X9O1HjQRARYkJv3wORyfcbuRrljv3yenzzQwmhBtFh+gAyIBxgg6cbK1t301
/gZQVrA50PdwKKWslbDDovOtVO1yId7mqBR7GH4a4paY5lAIVnPqStJNSr0c+th+
Lenv+MM86dgCf4D5uxjGgN/AC0icUZLTylC9N6Rh6BMIQVxQkkaw0Cj+QuylqZRe
lrRx/QHgWseTLVaPX8CgFcStaUWK78RY4hctdj2pt7KRPemiPsfTrVs1iKYAzmj+
cETC5bnZgO3RUFbrRvT5o4/EVSnic3zaiJmoMOTpJ8RxU648T1clPkv1YFjl3OZW
/kejwMFbJ+Bqg23/mV6V4H3rGNKOiuKNzi7YSt6RiJ6TQ3Tb5aW7mdFb3hsnxRQE
2YiJCfmgICLN12hWF+2ov6E859TiRVGxXe5INiudnjE3/EJ5DriAzgMhBp2qw6x6
yzODB+Kg1M1sFBPI1GlOAoUvSn6hXpb69X8qNfRmOv3lYBGbkgWLfRkiJDB7YkTl
a/fjsTgJ/1zt8BEQr+bY/tohldcMIRgyr84LeFMmaatYSaHv9ubwXCOAWaC7jJlL
5HZWwRvOnzgbdCpejAX46fOwYo+Dgcqa2Yhgb9TGPuGNxfzb3zXf+5GZvh/xNa22
DlfQJZdV+dOJ65x8XmNS6Kdrf/psrNsFbQFqPrMSpeDf8DI3nCuwWWFBthKkFuMX
RFjlwmcailFffKysdBkaSgAGmHpNiPSvzGRrb30NgL3C+EqjSXx+EHvxtMiINFCO
yY7jQkj4pphD+b1wLxoK3dPhbpuj4Vz74MBo0055AY1z73Vor8E/WWQR02ST5pUm
7fEUmVav3vaB3YLumQW3rP94DUOHh0924Mlay5hmXoxpzRjQsisbH1upBTfn06nc
4BwSg81rEPr7OwAMfpDVBY5xU0BI90Qv7YZWhNiuSFKa8sCnOkGfwEntDS7eV8rp
eUHVdvzq+Nhgw9kcpR+UrvWsCzdGtqIcJwyTNXbVu7jz6lOJTHbqto8XjZiDgMhq
kXWU+Yhlj+d76NFkjp/yFvPT87NSi2GcLGflmNi0v2HtLb2FvcNxf90ax2h1nsh2
SMCnAwHg0h+TUOnKRop/krRV8se5E8b3Dlc/6WBm1V9fcMoJ7ZP9XUxfAPr6LKUg
gL2+BuVJrV2gOJnzDzGWO/ftUXLrHw5EJy3FAzpBC5wRgkGnegwVedCukQsPiiup
MLScm+1LR4tMdYV4P4tbTvlr1N0wg0RcFI3SnXaSIqIXymflUWF5fVxk5jbJX3hY
MI9/E5hq8b8L0MjQ3mt6F40zZNfhYwd5xFeCQ+YWyk7bumZipTO/w0vsMWxgpkuw
2MvvfZQdQSVjGImBk7cUkMZB3MaBVPMKxCslbmkmWTy31oehAHr2uHT3bxv/pWmS
IlkgCCDt7pnflqpeHEt3wv/yBOtjJnRg5rrYTkZN4hRrQl1H60brryH+4UX1E3EE
H7LdgqirqGDFGPu85QicygpddPaV8t8WMdEwdMP/1WlXDZsf2wcij5I3ca+9f9ep
uAyjVWgxq5hUTWxGRKPnTvWsV3rKpc56VYNlO4nLJZlX3ePUGOQd1S+2FQHuPT8m
oVN0B9pgJz/3Oz5PuK9LJUnh8nXM5HvB7IYSxpSqEnlfdj0QbQLLDZ0pzR4Wh7BT
fyi9SK15xdlDOYIc9xBAFL/l/gvE5RKNObgQ2f5cep7OWtggwBKQQNpNHJn7c2ag
t3S3ggkWtXuBFE9mZ7gmS+X4YXiqiBtSRDgqlxa0Y/Eow6mL7AHy5laceTxhEjg6
GF2+5QtHnayWVBd+VlzNj7D5abwfS4CJGw3nzEq5DBOQTRZw3Tlb0SD51LPB4cKu
gmbiqfAPZRVWr80b2qCvy9QAu87Q/Vu0rnZQaOKVPABzq852YErMauRSmy6GOUeW
gMmL8upM4FEmUOmqlZ24WogAvEvfDig7/5iddD6prAjfCbfmxYWnmROCBIEDm89g
FdiqLgU41AAH6bclIZSxUWfPozTwOsKadyJxcjsIQuNY40vO7BxIU4+xOfTH2zB4
8zWSrlzKlC46LIIhx4dIoDXCJbFaY9UaUIhLiUoinvJgTESla1gQV+tQd6miqNJP
+LhX76Yskvk5Vr63gYlg6w/xAlHpUUmokixkD4xJ5bc0u8jeuvFaIOxAC3H4ideC
MUGTFzY6MzFFQ55RxN9goKu75YD3i2UdJkzLbdHxqLCOgXiQjrzwUISGQ/gbsPKv
0hM450DS6s99lCXEIHOO3uKFGguuUAbAzW+4tPyK9xWihkA9EzG4sCgw1ONEWHmd
82vmOnHjHDH86BrkADe0HGOD4uvUVGwbYGytuM4Nr2O1QC7fPABVgVibbgN04pTG
CT8TK94ouOjc6J2ruc6MjpmD0nyxZkRuGpX3dyyLvmZHGqTPPU9uLfqvbUS4p5Bx
BVlKl4GqjUzKqTAFEOFTQX9h4k2GeglF5noVr8wP7HQ9Nb2Q3Fcbtq3/Tq6EAYRE
k0LsNGU5ZMGRWbOW1mM+T914AxlGjzZPwkTjT2HWY3Qoq+QJBw8PGnuW4OLODz2i
/6UWItK0oY6t40BVn+3nJ5Ht6qvE/c4GT3dL++RDAnd8StegCymJE4Y4g+zKl05Q
rFrLSIEJAw638wX2tyDWzqS2JCRCuRqhlNSA8esEFGrX8nfkCfNGGKdHPVIPC3ri
JI28YgavFxfCKhTn59kAeKQvxbtNcdSfaTCOeJXZ2QcoJGKOiXd+nOiyjyhFkIA5
qUKlLACC6vyDG/He5qqN5TM7No8hQ/NAkHpxHVkRYHsJoujHkSAAQGtRWQo9d4Ov
bF0jCJAgJQTXS+ZYsXHDEa99hsPM12OBlmy8uR2T+S7DI+bSMF5xxyYaqkUrP/Jv
8VTghIb7z4YVWuq/Qr5fqDqFjBdOHx8PZ/AhhXr7GVjWG7Pjz4EEFBRpz9LVsoql
xDcIz/8md3dcbGnRQWeeBlML+R32PMmInA96jCKlBcN1t5R+TFDaXcRy4iUXTXwJ
9uGR6jZZvWRjgjF27KDTKqjENV1KAi26W3lElMCTKtUTqgg7dzXiP3H8uyANKn1u
xLh8GDxzsj/YaubgcqDWCb0cKf/9AODBYGnAKlIhY4CtJRUkXdr8pbGouEqrhbxk
w5owELS6SiRxCmOFUJ8mO5hGOKQ9BPhXqL7kmp46wOG6HBYpITELfXpYlFpJY/6h
fdCaRj1QCADjD3lcS3ArgyDbAp6P5pjC307fWJykc25cH/jc5H9MKiG2efsheFOT
ad0BIlvbNDeh20wyddt7Xc3oqa0mOAH+MQ/U2jXEcFvkGxlPKcrtnKfH2bS+Enl4
cMJo6tQ7G90q14Dei8RSX3/kHdJuAg7ZcQj0WRCDDi0ElSssUgZY7IRnkojoZoqY
Uy8Wot7rikX0AljLOAYe2/0AeRJuRCD2xgkG3EIlbJXkbpE9xAHvIq5C+YcxwT3l
eYLG+dVtnsyWC5pq245QgwwUT4yaC0iU1mXy66xgkURzwauWyTpudTqtTAgRNFH+
mTD6W5j00TpTiAyhrUQ0sBqH2QCJwehytTzMMwd3MSi9bNXwThx4qaUuXCdvsa1Z
hJfGFJqV9EpQhVOPzgmQCFBRquz5ulRM4e3s4zXXUOlnRTxOfLTwL092rhjmysw7
JedtC/FSI+rKIVdCSwfEnpKrGlDVikTR3KcBO8vR/PTmIjRLC/Yq1CggJT4kVqwL
WDdfFbAJ2WRzlJ6jdR51bwHYddiz/I4OPlVvgPuL1AeV9sk7QU5XTT20IRsY2jrd
Gckk2qBQmPSiClNAQPgb+XFXWuCwjsSkTene5g/WP9WFtLp6/glzrRe1jV8vpCsL
Z0EbSdiSP3t9ce6htHgoOa8TXgoKvZKbkP+0U/cniGBIW5aQ8nTMrwNGkCGCI3Y4
ph9Z07wDIFrOgcRH13bKAvp/g9LGQVZhgGq4gGSIzCJ5kAlZ40HHjQUNI2Zt9ICU
O5IHFCbMOfFtmU4h9acs5TM5TA1ddPGlmNU03G45ctegkBSKExhLxM5+1XPKqBfH
OVtfE2qYxRZXjYbl8VuKWlD6An3tT6M9EVUesIde6eiezP9FKCSzDeurEvYW4mhX
aXEYR8UPhp+Y30mz9qG+xsca1wVFum1b0k62CF13tJnfSsFKaJM9CAXWz25eQSN1
Bm3lpfuLgjuT65ShnSJ3WK5OoSFjuTUxKRmOdQhT347mJJ1EzUzk2mFCJQRqeHhO
kfVgt8FcKAxY9cLntKaYS7rsU1I2MrGJ1BFaluyRVba6YWNDEba/Ow+P/Q3qdMJa
6Dy8d+k+z2ipy5fIk1P2CJk5WH7u+uJOe9sneAyg5aFgQ4+hzv45fOG+0/KDC0Ut
x9foEPvH2AGK49IWYY/UCwDcpl9w5jXyssqzMLK5n4+5PheyU8ybD+tsAHlKChdi
ZKfgR1RWUGVr9QX9s1a+SNLWRH6ClsblyRpbn7vx4axS5MMVlKCLWAlkCG3Zgkfi
trm3uh9d3H/iwWso54/IIZNaZfT9/5PtwqIWznLfebY2vV9u+xVn/HT14j5SWZ4o
rO94Tw1ifTzo8xVdbHjffUe+wyhcjTk+v4ta9d5sTpUVXQHNexej/ltTc6SJy/h8
R103g5SfjgcCiXldInupjPnnb3tpyIOicmpJfzEo9+gA3X6R/kirM6BxBMGkQUei
36qAxb0xyLMDLtSLxSz97AHThBmcUy19jkRXLbHt+976PIyBepQBXp0RXXEGhJXi
P9ThXC3wVtjhDa+xRnf7YhseWRV6x8U718vlJ4/FdRVMul+qegJWxY7T9SCJrEi0
QGPALD8dETzFp8nUi3FF3kOpMxp9aQ8P/q1M6YVRPy498p9q1rRQM/1v77xkErlA
ntyW1D4nqOpJ0KOXkOQEFd01ptgn7tDQfPxmeW19PHrBY/5rWvMbC8IKdYdcUJOB
dlGD/8ISPqjFuYBrvYWTFshRbi+z3Vpq7k9hnsowoSAmKtAHSdu8hZsffdArfUVx
A8MDGlBdnuJGh21ZFwFIUXMgAQP/i48VLvR6b/0Nt6J4Yc92HjIIfXgM7/HC5nzd
RWDEIZWG53eGLiEaNYOtEi+p2rnSOvod9hlAqtB5Go1R+xIgT8+Pr/9h394rqeGd
HznkTVYTLV/Ac+O7qcw83Xy6s7VkuIp05GNlQhn2n8QV+IMb/CXVxXADGLUs0v6R
baOlHS7e4LHADcwSFQDAzjeeGwNzkYmDitln7u3OW8h7No9KJzdjStN8K3i2Y2eZ
kbK9vKi3sLzTvfOcG+Zn78lfs+EBb2Q7o1M5xeJ/1SsanZKZgqRSsHvE2boeOzZy
DlDsGSjA66Agi+iHanSGqn2dBszLrDa5pu+IoYpwVOaJOyzGDtpAgOzNUyyJ4QEJ
ROYv1uz/5bWxzFtdMQVFosgSo7Q8xSNjvjwx3HofmAl00bKKD+GiG6Nf0/sF07bQ
4F04Ix1rcbynjwalfep4XP3QxFSgS17k7MfE6y4eGIb+tlrXBJwWDpRUYuGv30kL
JSNVH20A55tbtc3cSTmwpQKyDzbfXVxKY12yKjs3Qc85mHvID08p0TXxADg871Jk
3wKjQs3lvEHZqZUn/Bf61+bCxOeaqLB3juXRyNvtWNiwQVH/xnEzX4PWNJXqY7aR
sTEMjFNEaoIoybbq52o+Spe27cwuVfzPxA53EaRn2jMrxC/6LvYJCE/9HIAI4l/G
Sf4cXK8fmZfiWonKwy6YaQiu3h/6EAUF5EiAIEZx1oMBnt7Jyos62Vqg/T0nABIr
tVp4Hd3ME206mwmnbycFDpWSPjmJ946zMS+QtcJ2I5W/M4+qWY5pei6nPMGM698n
4GPb8efCBkWUURngOlmXVi78uVqPY1cXzFOs+N5fvsR8ubBietJOe6DZp3UroXDJ
y7PC7jcR1daTCzecsrSTg3TVLIGWnjld5Z4mFqIUM4KFOISNkH9mtzEORMTFWDC4
GiYZ0jxeigdTlhPdYhdF4AB7B96F+5F72zLp3DePokY/NcPkNQk4LWPIqyuOKa+t
GlOefhkT/pHmMIZmLy+EHs3mzRmd7Tc2iXPlN2xkDLTNWyOp6fJcPBJK8DL9zo67
aL+Gi6z8aoSlO2ONR4ri2TbFcS+cSMYPJxr4ZYXewtNl/xI06xn5dNWyRGIWiVMa
Bx7G6e8Hu++AYdK62qteeXxzWLyR7DS0oGpthQ0oMLUNKGtE4kaNuidP5GZTlh3j
1StZx+MF+NPe62FYUnn+zGKekAajE/8RWzKhy4rv8yDxuvj3XnzqZoRHTkaX7Sq8
FoxDmAxVgZB3GIloW5bdrH3qPaPZkPnIoLfHs0LPtZXmPHXH4HPB6VMgBGvlWXmS
9Hl2qXzjgNihLhLHxXM+Pd6VAMWJJfjWEcG8kF9rxlWsoEEzvuZzaE7/cCDU8xtP
riJ5Qgvg+ap4o37CVuBu0hROKvorgQQaFvLtqDkiVrL+PYqKnQq2736WpIelnSND
6CZBmbCJhM6XxLKH2KhUm+mM6OUCfPakRgNA7MGRR1mjL/peixpQ4D/BhPN3dkGh
8CWWruPvcB13K/f0FPiGWDSjrq1BN54ChyyQFg8WX9rF/mJH6zA/SV+bqLp/j92G
2f9fi237bUKMnAm9bviXT8i+VaEmPXid7ldiflxz8ZuywGDxoFzlSteey0P4c1yq
o1nP5vOtI7uk/Cl4ACPDSsjSzRi09eqVd9XN6jhhOK+RZExN+M49lzkZQqeQGILu
mPWWkCOAu+dd8UB4fDwo9JwOf7yqKZaU0n2WrYZqF0S9tDLYtjU4FtN5C3uP/PZW
hAR5mO4eBHpptnG9o1LiTKvAjM8PbuHmbz76suKBht5HdTfOnh9h06FYpWTxOnpB
BwjjASq4+LV2/95C5rC3K6wnoOT+Bo/FN8ltGJD1XDIBtkKjz/mgVTD9ByQs2POJ
AY1uYesyjQi/tdWbgqEzN8vGqfwHBnfXnKzh5zljgCiEs3qX/N64ZQfHjIFOTyBB
iSTIepAa3pNc+taCaK1USQaFcpy8AQTJQHZgYfgZQUoao4qNc/vLzhsPl8JD/czS
3tDd09AN3WFJMsMngaYqKi1lbhkx8LUcRFcKiwBNs42uJJ8Ctma25dLeAdkgGx1z
wJsEPy/LzpZRwHwQuJ72vMvdPtewcXd7EmYlgKnyMG6cxalTp/9ygI04n4PttqMO
5Z4N4qkKW7KJP5SUTlYpWTcDqq/O+TYhgrPUp55SVo6z1xeRD/o5ae8ZPTBoOWc4
sWgGFWvSaTcbRxzdqRs7LErnYCFPtvV8/iFKrOUybYdsVoDD3h3ujQ+6st1UOgR2
jtJYs6C2lZoYas+LyF0AtvYFosgrWib2v7dXi2WKOeIlwQAgwSKlEOkgSz2djryL
qhAhYmIgL6dBZmF1Qs6sUxpPjx7PEmxdCH9OqDJPi7nJ1jKWnsVmAJtBmeU7okz1
AitYPwW3EyFUn1iUQM8/xjuiYkRLlAP02x30OOvLfjnur0XfS1c6Icawr+GX+TvP
BG24qz+BAQjBsZr78IPsTM1MEp181fqDUcbWox0lmV2WYJz7MmsdC8E57GapG1Cc
BKkfQQY3mwp2WT0UFHG3XCzC2TkDlziz3XxnJs4qMOub0t43J7unhpwbpShOufHi
MWoATYoHPqbODDN5nRn9w4AfRHrfQ3Y0kLIWAGv6np6nTfWJnQzYx4VqEN5LUlbI
AKWIW6jXYObQyblY04ROhlgXcDYJp3IhYiTTr7QYsaJJHkRk359FS56lvK+7DrnC
rKV2tcbmH0oxLKUkeXTE6HDasJald3gOhp/WupuDROwhJHKJ+3tJyLkPvTcilsGo
7wQvVvt1JZlO+46JjwcYyFWMRxYL2QtMYxivqOWl9xg0s+zWPRa9vHIAfayeJB4E
OEibjBAcJEnNBjIZTMQyujiDgKBbOkl2WerS3OR6cIjFDhVzHzRukQPPXprtoYRK
fuAYpAmbo4PrWoQtvOfftNlfDZ1cNppK2PdjwsXaDb1YMub+wO8TUBcKeL0GMhs4
XhrhNi3LoGHFCbYNch9mIqw9HnPFqLoST316IaNbH871ZGdbSRdxx6snjHMNCdrU
wFac06KOHpmOwD8KRisk3kVtMt98o1e3iHNjS8iTb/Fw845r6MBggdGqA0bOng4b
1JXX5DtHk555NurNlONvZtNWUQh+0j36//Xk2RTNgTgZyoFKzxqhx0d1KI/7tgw+
S2oC0lBMLYtY6H/8Ds5fdnUabHHglKzC+orjUphXNV95rQ2eS5qP2R5bEpmB6OWB
NBPyr8MB5Zy2E2FwyAQgxs1PC2fWcl9jCNoC6k/yQvnzG2x9Wk/BDs/+wrQze/Te
y57ArIaTbNx8s1Tu+QYEX31UhkvnSudogqk3M5EJauBC2cOr9bZCGZN9NbI7RgL6
wQG0nn9Lv/NTxi5RH6+tlu1zlETSCO60NLA0XyD30iFQvTkqDrCmV3KA4ZnGN34e
FQZ23GiHZ6ELMn/y7p4Y5ZcpPbizizhiJ6rmPPAzPKwsXCeH/KcV4PiqTeml6qaB
xLLKPV+rAUvrA0/4xo4yCWPmpqzpIAsNUuxqd4c/ZX13P4GdnhQ/UFI4ViDW5NZF
A7dG29vmjXERYXA6vdV5yNhPzl50oDnJHtQ+ESZaB262vG2s/riO9lNeZGXap2Yb
m5mgP0lvQgKUDiUfvcnEq/lmL/kHxj3pcDHJMQN5Gl+YkxRnOY8lMigKJjphaHiY
rBFm49KC9O+cOIFOmoQXsRA/8kOTDHQEHRRu+sv9p9WeEIZcE129fhPQCpIYlw3r
xIVkKvg3/lVBw0wrqjFc+HRtf1TAdLIO3OiyQHhpqxLjgOukx+ogSnYiv6KXAk38
6bd3nbIF2Z8len8t2eNb/X5vKZmaKHQRRFhnh4oa/zRMrB4RdvgLBSBRVUbV32uI
7Ck3P+CVvV0qqtWejWDbHg==
`protect END_PROTECTED
