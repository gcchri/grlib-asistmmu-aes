`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Eg0WcN0NoyyzEx8WslxtMasWGJSe9ZOSJjko18d3HFyItJ1YIW5MuTIVIo5sk7AY
ZbSe2dygtc+PJ8CUX8e77f7a7JP9aup930L+aX13KddDD6GCdnX9lWenwMOSPUCR
8uvHzXbv8v9aZwa058uHAXJBZrr2pf7YGdcURTqFjxuF++4ahjZb+Inbmb+j5+6T
IRXXGzuCIcZGldPR58cqpcMmKBZVd0A0+bVU4oWAkwvu8JXckq6IWov0m7kWjfIB
xcN0vVnkIpI3uCidCTUtZgzoB7+qoQIoJ9M8zqJEdilrUgmbkRvVvTIyB3uKYEw4
n+aaXJ2Fmu4dXLc3mjDs4RGKjWWQl6GPZdaVMgsWApJrRtxgeHMmaRx83TyU70KZ
F0rSvv+CRjiodDq5kAFGBWtbGWcltRly4+c0UuInVt4iL6dEqmqM7bxSwqK/1KSU
`protect END_PROTECTED
