`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z7/sF65/REwvOAKg2aT/H8G5UVvYtv+5e8zOSG3OxmvSQ33pPpmFk9VJGa/6w92s
Zhl7EPpnoyOoeztnYSy9YRAxPbkHcczAnTQUkumbv9cByEKoAPFw3xYUMaDN/svI
VCinScbhEcPtdb+HThSM7n7rbh19NNo45iLAKVw8pZUTuqNmJO9RZLIZ55843s9f
BpopsXfLbbCfczjzjJgKGimKpYjzqJXkXBA3FneUuk95T1Hfotzu0MJYdPM3SIXS
E2GpNysP3IWL60bWWhWJN7K1Q14/Obz1Z6tLVmZjXv+WdcxS6D2Db9pFHk4AGH/H
AQgiwZcvG1vvSml3qJw3qQ==
`protect END_PROTECTED
