`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V8SDl3AdUSkz2dMcVdN60sOfok+o/LgeoIMo39Isl2/jCUV4TIqSH7/O/nvW/QHR
DC2k3Rf7zScG75cggSOBgsel+wderjYOlf+72MfJiV+3yejKoINsQMpuMcZN9FK9
AyAQm1+UZp4PetiF5DRjDOWZTDVIlv9D2997PvbDnBni0ooy/DO7Jo1A00Z4vTib
eFvhdq5Tsqz157Uc2HODTrpAgeU0dRd0JC0szEIXO2K1y6Ch3cm8TDgNeSGtXwr9
hMr0lvVTeBGtFnBK/HM+Pg==
`protect END_PROTECTED
