`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y+mK9tEC9oyKv7sFEH2d4DgzI5Sycr7pDMMedg6u7NnG4c19Re9f2MAJmEykRlN6
6jURT1uxljlDaeFgzF6JdKLS6IG7AUhBMjxhlkHuClj/Bn28juAEuM8kYruSlGk5
Tfx1g7Vd3IA7wwHs9sYrsjP1tGvseUcarjc1OehAxa13PK7g2jVwbnTcVTBPXo/x
RD7d+JS8oxb6Xk4dCmGYhVFiuLJB+rOdqJAIq6/UW1vJohlfcCdu4PsZFVte3cQV
w0crLnCox/ibsykljxAC2/8L6kSUnsmhuDt4odYIGvzpRDBfSTwLoW5c82ycBnYO
bGsKOWL1NGu/oYwTdN8txd/K5vGTJKZx11tEUZ7ZQ9EgIh8POdJmlyFdxok0bA2S
24RdkT6lzk01481eJusIo8T7SeUYVil2UpcrqtlaMc3WVTcApIUAlzosRSDzVmz+
cUaeILalwc0nTMzOTGF0vMJNOoQXmIK9/r9VKsvBRfbDr7176csV+yXgGu3Sdg6O
O7VwHcNshN5B6xh1pYlFLEhorK/T0svAhqoNcVYobK/BZmQCoHjd3W9kc7Y2Ctju
OdY2Umkmd6dIh9IGBop4HGXE0U57PGbVh1BOWrN9tVb+JG5AIN0DMMGocpzWJFOO
xT5IQPAeRefLwU5W+SyWPbT8zwj+6K6ctWdS6apmwJjZvfiomwL0IOdF29LI42mo
gf+78A4LYjgerOIZpAnxkrJND8XN+x/Ch2BF6MGsiG75sVqdOcjjeMF4x/ZkVbEQ
2Rlu0W9p7+wk1tZKIgLbUOvwxVFQnu7xFH+UV2isiAawKRrQ/7kSjdcDK0wr2V5M
GC1wBYiE7T4zOojlrfK8TNAh9uk1rbGjy6gPSU5asZiKhTpE4NVRUm4Tb95X5MWD
mk5Y+pJbcnZDvZX92rT3H2tC+d3z4ukUCmp5WV2fpl8hUnosd/xA1+fZUY+4iWFf
JCoy17u09fjfOxgLfWisf+BWA58ks//ibWuMNnBd5lu0g4VXz60CpOwq9uqXc2sC
OSXyrwDn2aJ2veiZB8m4JsqAB3MiBpp7httVdcdawnGo0KyZs3nOEz/LqKJg8oI/
ShqZ5n6M1NQxTY9m/ON7aYtipDAMQdNoIgVLoZWtwbdYLJ3wUCUvlhpzhu8zSQPL
`protect END_PROTECTED
