`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wfuz4Z4eIW9ITl3tOYlBy225aCahGO6P0K80JyXpPBV8eB0qtDjz3eBR2dCoZkj4
UVoOx5zhrgoT0iQ/W0exCXO7+vOHby+WyYRd49fXfE7NmNQVvl7jYOwerzBOJxQx
XbmqodSvm+rAqoF3bXCLt20d/6XLqecKIwLlQ37UimWJ20OFmLNUnqEHi0rPW37x
Yadoc6zXWZHyd3Dyq1akurS8ygpLTbbgZiOMgm2HkVfDXNaYxwb9y4HOR2t0lt7e
17X7Nk6v0j9AXJoAnydYv10P7rgkFFu2ftvTV33pPyevm2VPNVCYSQFwP5uNxcda
bj58pnaz1CW2EEYN2bRzRKU1zdYi4WC4rFVVHdDZiccBc2VN6NZwnAw4UEhzafnx
ola5euQ8nWsL6Ui1+Eqyk7fNXRguG7Yv4SHOgVzOZHef6oKxPS1daCJ5hPRtga7B
3ImqEvZPYaQ6GVn6DJF+BjZOtePn866NUIa5ZeRYSjR2uACkNiZpAk+2UNhrIyBk
v5eddEjLD+IvDIvM4/Y77t0BkjzsmgUJA2THk/reaCZGMV3yG19k1G9jrX8Mk8Rw
WVvb/Ad6SIO/P7bdJLZ8P78E3+o4LoGyycA+AZAy90acXeKQTZXkk3fJYxk7a7dL
5jpvvhofy1QnvMEsZPefjD54WHrf+LWawL8bkQ5Z9h/sxTHe7VjmuZ4OUYK+RhvM
Bc1aC06suioI902BwtzCJoZg/2o6ruNG+6VDqh5CHSFFqr7Vda2sJ/rASKd5X5oy
7/GjvdKnqU9oKAUAFtZ6pjTZAzgFCTAYA0UZ63XdnMkLXwNNjcmg8+RlDylHy5JL
4cl8hF75sczeAz8qVLhV3jYIxOzkjWPN1BIY5+7OhUHjV3PKjq3mpIMHC1a40Cn9
yEOB7b3q50dPWle5PI/hG3v9T5iIlcHtaGJ+0eV6+UJP3omCO8mAQdhXizYO8t1N
iVVYyXEozVO62yzHNl68zwzHjP7AEjz4nrFRXgm2ZxyBI0I3QyBnkKU6LXGvNUJN
zKh23Sc6wa5ViuGCdbRLAmKcwpRIha9cYKTcd5nNND6c66lkPMqBhAj09q3GS64H
sV9JlrgN76xXomlgsSnWKQEllIaMDnKaTUHBQ2NkyoEW/QNqmwxZbyX9FiDUjg9j
7fOrIZDj9b3EyhagQfsaSb6wQ06CoCmRl653hBPpSovPMgK1kgFDXuxR72vPl2Sc
cp6/Ifyb8jmNtYvYAJCo+ud4r07DXspDPebsicLHdRlMLYizFEjeJKN1YWgP+Urs
sfnB0lFauT1BzVzjFsI75FaRQqoM8qP8r/TYrZzlEm9YvNNvTq0k9Hpv0uooVa+K
kh78pDufAP/boFfdcPP7D6Pocab2lW+OQDt9cIINDOtoS1X12z/z1SLtBO3/qx5t
lHc8rGiYeRwccRkze1HFAALr57lltkVFgfajvJVfJFR0zBD+vk6UUN0HCduYwx9A
2bcklsJGnPWf/fnBVjBJj8GidxGZpVXXPP5XYkVUSH8/6EFIVbL0wbuJf/NxLub5
cC5EbEuaLAzC4JOEhJJ2T3sHTVVUzr71+B7V1EYd1c+u50kAyieHRseCPyfv4neE
Suvwa2tKfGFn1MBVciM7EleYoEzuYxLgOTE60+HIG6tZYCeYpnoq4BCpBTHaLSws
yf2s/NQtuHLktT4ITvK05m8dSs/V2yZdAbizm2oYd6rVCKQVZaKd4BhhLxasJAvu
Rojmm4X7TRkFHhp5A4X25ZSyqjuRCA5KVYixjWBKcw3O2rZjsMGyt5HFjqWVQYsr
Toyf3goLCb7YqogtU+V/et+/qwuwxNP6iDVkuVrdA/x3lI94lhYUrygDI9fsaU/M
xFYLoQ6lveGH2ilM0mG8zBxq1PEgsWn+Qs+vhaH7vNza1ttG2Ri5IvlO2lK/1H9b
EOm77534/bpNFnJP9R4DTudRUyGgQ5xlcqxXoPyCRXlDB4ot6sxfjnb4J8MU8Ipp
VqUtfRxQovZc7uySPa1JCcz6x4yXklmWt0/kRo0w2ejSd1BtFk6mQGBOzF/wEcFH
1DAZrNO/NGChAdFmOoK50Nqmt8Q6ciAr6R4xnkjpmpMmv7zmcMiT/Aj5jFG0n2oh
ynpOfSfMl3Nom6q1QrJ0LsQG/XFwcfA87thBunIzwSNFDnPaxRssPXKgZcoVFNvp
Ufk8EcykyKAL5/IFt3Vf9prYY+sa0WtB/0ueanp3dD/GdGT/1TgFQNTpLkcMw/Rl
/0MDlW0vDZIF64bhFfAC5XLy7jZ8M58x7w350AfKK+g25u7XFfEjyFPCJLe0NH/q
g/QziBkIJetzkaOTqr4hxz+R7/E4/sSz5xA9QAXPVRLVg7qYI3HLichVUB9mLm3X
rDDZ71Xk+ORJqEu5q17CW64LJJqRo84QdykdVqBAy4fByBr35KINHRILdzz146h/
MA/EVw3vlhiSB1W3C++HWEVlR+KH0uhsS+xwGzcS8FOEcMWQ+7mR40ntnJ2Jwa7m
0UGGOTC7IaOrPEG4/sTYwOHYdKGp2CfAdhn3m3TI0OeeUGyKDezsYT1IG6qj2RAV
FP7Q3kSgMrpFPlFsbP0lU/qmR39fjOtBKx29LAkX5JIOy30oSfTGcpDUjFcbQrd8
CJRbIHO+IqVl5HMvY6tMTVROKS5D7Wk2uh/wYkqGXWzMFL2XCVpqxUlzMn888Evw
/9F6cAXi/xWZ4N9+Uyv3rHJg/XR8hm+BAHsfpNAPnqH3F7yEmOYQ81rHO3oWonRt
BNk0GE5UtS+JYx3atlTDbyPi/MEWaybKZe+cSMA7N1eSK2eJgCwKqnZ8fEgs1n0C
HTQLbHLOn8SUAXx3VrSAPnO/kwhZu0CrFY5NYAatmyXm6bATgXFZWut5ZNA5jKnV
2u9CQZJy3Rmg1Vkd755QXvo6cEpp857qBPS2nLhUvCGmiX5qCsnj056Ru9GzH0RI
Nnz8a3+in8+WIncfoaxwLARb226fBCkpDXRmvEGOz8YsMVhkyrs0N404NEYN4+V0
fmS9Aokw+WDPyZ4AuG90mdgVmXjKLV6U7QDvGNIUbmBVgsVA/Gi/XkUmD0dDew16
P8bSfwcj3CBF/sS3R0UQjZiyBBQ5c3w8lRJd8J3Cj442hfqQrGHeBJeuxPPlcEVU
W7Imb2ozCnpgOJD0Vk0uxUBHp8T9MGYs/pMmM5EbnyzgnXjXdsORFebw8vfqF7KP
dQVdKcXpeI/s6TNSkSQEHn57FqxTDTaFfd17i7MqKslvTmxPrxCnwE6I9sVIfhq6
x/M3jnF2cJZ4dhKakUDUb8Z+23e9OTEvqBXqJGqq7dB/PzrzDOnFIYRuU/+aKtrm
badlgqpWhFzbgU3d4ouPtlU7oqBxRstn5W0Z2Sv8D5JvhmK2zV+eOlhc5N4j8p+J
LYm8v0cGWCOHOvhumHb0aoEUq6ipE3fkj8jxKYsPkkydQ0j7tLaB5uM9SUppHirn
85j68l3fyrPBF8Hcq7rpptScJ97lB3SHEDMR4AKE1vDSagkrQJuNBLcZl8Z1ifm3
Ybj6SWBJfWHnXZTpr4+Kle2oLjqON6vfiVZ76ap5IzR+WuGi+FLNDsdburJLxmKL
cnTxnIaz2Jrv0VnhOr1ksrYKva1Ik8zQQtc7Y6Zadj7l2dGstuGqVQHvb3FqBuZZ
7IGuDiJ6hTEsssAyVabLaA3iRO75pZUBSf0GrK+sBKGt1DlFsRXAXQh6bFhcf8u8
OMMtuWgnxqBh9+Z++cGW8Mn1/Lc977V8kCSSlIYtyOO5FBVAu4hgGUp1Wu3qwjry
MnVvqRNLTi008L62R3JDCIiVmKEExrx3ArkYGYWa089F+K4JSOKez8QkDAFLNoPC
cakgH139OZI+WCOpZZbTeFExfryR6bgVVUY0T8C/ipit2fNnYm4CI7sB6t8EX6j7
p9f0g21ZCxhCPlpAPkMwX92prVBTYdL4oMS5JGRLgmHY+o5KBsqAfCQvGDVq7gXL
IrGky9EgiEDcH6l7s9CQgjjsmt/0CYbfSZM7fTaiyuwCzuuxdCX3rZ8a6y54yove
Bd/5j8fok1YodAVfYoSONlTTuw8hovT+hRczXDUj8hLxqygjtXPaMlXr3dw50Tbg
Tc9FHF5jNDz+I9Fb/42/7wWJYfShCqYSOyDXk1RehV+zNMj6YNc0W7MMjqQAg6xQ
cDqSZvhnuGFX6Ho7gATTMB0ulVTnUrBqEsnsxMyWq987/KQGFX1ruKNwqkHpgQNS
MhAOQEh7g3VV9HnBa5bbOjghPY5y4dhgigwOTb3nnA9JtdhjzIZhACojVjkOj0S7
QBtRKEYCMwgIGKq2E+9I3l6GAgIK4mvwn0aXkFEYwZ3kTXALEOhtcslXJyG766Yc
tdC4vzT6sdHHLO2kXf9cZ8kB/iohMR0bTM4s1uUtOJPi7T6Kacu5rSSJDWq1Ggh6
ysv8Pe/C8x7d5AajybnkP9GQud2rdOr62Qab39dLT0fJ6utv6FQsqXQus8G7X7rs
Z0RFnjyHV71UJ1vMbs43aQfwduNSg5k6j23dXQCHY3Cf3p8MWGLyAMH55QZ1FaMw
by5MBw4uj7kFkgko6+UCAwX3ZH5PKAfs6DeCcBHwIX9TFTIBMWkd4Sxkr2oTaZZz
EdpGl5yH1/RW2dQ0+viTXFP24TbhxxqjB+JpG11b6bsjYbGSfDg/fsK4c8ZtvtYh
GYnEqY1Zu9a8Cf4SvDXwo489NutHqsucDAu2zDWAR7qASQijqPq9uIPI7UITnwoh
ezmbEttjsW08SnAiKvjNDAxDVUDbsAEdEDzorkmmcK7NB3PW+WQZ11raspjBaKA1
52Hl4dqMj+UiqMYZxrSHED8a2vopBmH22wiJXqIfNkttJqCY8GW9k8VjZtPkWE7N
kz1k7y5wQdi86jtzPcOk2UNNpk2F+bb413/2WHsZ8FhNsy8WXTaWsWPcyyCKaH1z
/WnqCuXLl8rINK2T2ZCezRCfCQb66YI/UjLNC9agJXNRPmx0ZLYTqiQUfdFCYRxj
ef8cXtpRG6h5uv265GBtxooFpt6YckT4Eq/jXxw82u7ohz17W2H2ILVkH9kyb5V3
8rqxJ2120WsXo4H6NETJsenk2jgf7qef0zZGpN4nhbJ3heqbS+i7gBOH1KMRV47g
0GhbJhpiMRuXzRNeJit8MuO2QiVghQEZtddJyF1y7SYXiPiCpb6lNoz3z5AHV5Nb
Nq0lMOTLulE2NDCfYU3LV01qbxwqq5DBrJn+KyHC56sMkNoHUUzMLtph9fP2/Sfi
tvGrYD+zNHS8Aqt0r9sfgw/ykTUmurhuUC0VCVrw9cOARXWFirIylVL05ESETxjN
ylMFUef/wjEcjjIYYsaGjvPjtbgeWSXy4DifPlpAFHrQpd0fD80ujIcaYEWcV90T
MMA1WspvX6Toc9vK8mF91GIJ/pILLcCQsuwgVa3Rxd52ics6V7znYojCuN045hxg
4Esc3WNKTk+KXUkcKZsZtbF0DIicSajLuddpfDtinhs1fiKnj68Tpy4UozJffkU5
A8Q+nLxMlSLDRQxwzy+Ta+6ghOOTPR9+0X4t7bIeRu7YEs/gGTCCGn8PDc0pqNlQ
d16MgQPY4HUwUFlqI54SruekzHwApEq/yaHdxnyiLsaVHJ2+J3Eawik/yAZ+tBwo
NqOS2RFBqyn39KLEW6fWwZWAdqzdZ1i2uA5bNXvbguw/vqLQmKUYHdkyy+vrFs+b
Tkx7sv7lDH/lponmcmUcikK1lTkKGKR5U7L/uFrZERbWt6/BiakxZm8O6pwVRIAw
7a3O/dnmF8eyfmdOnqjcb8OCGoVVPpgxEx498p31veMLFd0WxScFAmKBp0i/+Y7y
PDcCusefHyhQu9VLvqF7FtCefX3oFIf2aMQ8v/U3baG6N3z0yARZrqwAWeBTX3E+
KuBYNz30O59mxwih7W871Uo1MakBu7dBPl+v7bus6RmgfonCgmkrzGOR8cYByjIR
fei/+jUjX43FjCe65DmKhxsAS5WbfdFkMCN8Cio62FAJ9UF9E0GNtxXhP7KOauab
ZHuCmN9tf1C5m3vz7/yjV+fRLQaN5rBIZohCFDZcw6vYcApiwAL4e4GsyDH0Jn+l
pmXVTyRajjsXrDaEam1XS/k9LxCuhvvUd6CZ/tb8tANHTRJuzzCKhHhiYiwelwOU
IJyLVROYYGS1jQV/CI5TAujFDju5Cn6/R3klZvoMeUDHhWPQ4MdtZjJXwXpt8f/j
+z9JlOacg/QrwYUIiANe9g4UuSH34S7WfZWMAoRAnanSeeG/ircl6u1d5THT+9a3
zKPZjJ7ZnCXMtIcjXq5skMlKf6HGW6M5647OWR1RkpOA7RGDLZu55pR/QwRFa/gT
8NglG04GnhSyXP9AU1+42dIrMEpSX9A4d1o36h6YrQbH4YzhS0T4gPOmAfvkp/IA
+zq3mItru4H9XcppZJllB5BdD2+omIxsEHqa+HHtHuVsK8ETcohBIY+aSODa1W1W
JFGOCI3L8DCtM40nSfhY+cPXC1xZC1kp18hCDwqnCSnGUv69kv6c2yQsGqaVSSZw
ZaQdOx3HeLf9ekda7J6KLzyNbW1lulg4a5i74p7I+7CENecSPKZeiu4JqkkEWpQv
vYS8zmDgRRWmE1X8snN8LmVB8epw99GrUAMijM+xE0BRCkBklgGwmcuvUZ2pcbcC
KRbk7mw3azCtFgZjl40f4Yz9G0gjSZLBo1ur54TWPiUupY1sRC466s34/HTkJPKd
wvjuNguz5qiY+PWv7uDOvwX60ENndk+dTkM0+HL6hWcUYdcYurB4wPFtkY2HFBF1
zmvWRkdk1vgSzn0OIKnggqfR+i9m5CAACT+mKeamdSSmrDSE/GPJMbTPNhV6ZQjs
NU50XF6yt86nyXu3R9jZ/DF3bO2XnsDLMJNcbBbi+s9v9y90fhL8VLe2SqGgN98k
KoWYn2Cxk0iEvo6/vsuu0ZEB6KDL/wJTxU+RrGfsimF7gmD+IrgBvStGt2O7XBaJ
XZp3gAuPoV+IdhzwIo/FDSrD1URw3zdZcn60yjiKNt1FY53x/SdVLdgdPRqIK0jt
+o5dBp9d6QoLn+2o30l82Aqt6VLi0Sft/nitDodFt73hNDzuKtXaC7Pl++qLDJ6D
ypQkGbAtQJc6UXFnh12cDHf4gWdlO2NN1/J2p6XsfYlhFe44jJbtZLBaz6+AZcLZ
0ZrUEtei3RhIq77bMEAKhC0TgrqPY6bxOjgteVyo9xre49ZaKzCgfM/DlY29UFOk
pyDz6OsBrnR7wszxens0LbEf0qWQx9yBRizZmWiFfX90LKQLUH2WxBQEquzYFA9O
jGIXlQBc8mdYoH+6DcYsPdNulModLAfgkGdyijkkYD19tz9zP6LEsBv52S0eqyYJ
qA9hso7GAQ7VAj/WpvbFHNq22klYhcqsGGpyBJ7ALFjLu1+Te05Lob4ewai9NQFh
AiFoWeU20UH6i8kD2gRm1digv921X9C5CZP7HSm/RhjnIh8xHDku4wBPmq+QfDAP
erSdfrrAls0m/7w7E4+O4KUCYPu//hluGhgIWB8r0nnvuY32SBRB4wrPVCcDjHTw
oGt7CyQccGADp/cZjuJ7gFF4XIkvxb3sGoKMc+E+mQJWpPyKjuHZMO9/AIh8+rOU
YTJv1UENoZ2/Wq5fCG9Uehu7rgbtHnEwvB9t2S2cMPl9MsvBv09vNoTqFVzuYV3K
W8XhVDC+seC5ZaWQ8d5FXAfVTk7bcG/WpGujGajKda2aimiKRkuMzYO5tUz3Ph9k
9hGcO/iJuBKL+H9vHc+vCB8hJQEJ5N++A+ubtSYL1UvItZJA807fNEWdxcY3mL3H
JiaOvZKD4wA7CkoSJc/G8POTZUwLQ1Br+nlK7xjYQvnxkJpI1umD+aZk1Gg2mhvl
6SIemiR7TD1kTGxz7aM8mnTMVy6cOVxmhzGFYc9zjsmhqz3WrY6fljfJmjgAR2Qc
h4U3yhqwF9a64QtQFf6Lcy21Njyfq32iZf4L0imzLqa2grGxMcc+yrJLYBbm7/l/
nq3CNMT+xbYwhug9pdtABxVDs3eb0kT58goxNPB3F1HO2Wab5EkN62tScdSvbaXI
e3MnvT/9o/cc5tCxV6DC5NdPgJLqcEBnwcFYf2K0Wli7gRkbm/0MXcQq1O5howd1
fBZqK9IKp0FXOxjA576uCOVnLm56cYATvl97Wpn92eU6oncBxgV5Dgo3Wil3onIS
XfaPW8TPOO7ojPyGwVoAkSN/w3vQkj5l/w6nd3PtC3uKj4McdgSR6UofR5YPuxIg
bCgCJsi9Rn4f0xGVJ9NSUvysAl1+Kc7ub7bwSCkaBYuxxKEbIvqhqrUr5EAddvWX
PzmpB4U7TPSQR5jVTvu9x2jLuSROdFjW0Qmlmg+jJqhZlRRdTcMU4G6tnJFsviBJ
PFmcvxGJCpPte1S0KdIl+iDtqr5KG6Jobu9FRRKzjUm9BvVvur1ZUn0sdovLs3+o
/HAwuw7PbtLZ4PbwKduNjo5BExnJluSGp/bzZ4gO8fE4UWJ3PiS5eRFJr9KyB0iI
O3PqW2vXV8jEwVaeMbbcooENUuY3YS6IQfx0LFUfDPBwcXwVI+tIUlMluqbxkHAC
+NL6xWIFu4LFsIfIXpP+DSABfgIwGmqQXfDC6iGeYdCSiLzYfEbMhY73/C4YFrD6
bsj7HZH/aXx4B/Q8H4SyP9aiaAQjXtBXGzdo1plYW1apHcSqFdc2252RyLMHdAwM
B/5y9nt4jRUJDaDn6DNiPZlVudBDguzVq12RgOtxgp5YXDaj1KTJLEOpVIA7ap9F
cZ0JkGKGvc3YvHu+faGmBQo0AXFA6+tZQL2lOdzW+IFJY/NZ+GBh+geA45GJ20Xd
Qga3gaTbJM3DO+qWflb+xfy3tFKGVbUUEVPm9NYWQ8NAJzjIy2BgLy9hYhuhNuu2
kw1E66iCf/zve5Y8ye26cWmU8jPPOf649Cz+dX65TfOtjcNiFWrmO3z8zhxlHiIv
dPM1o1ZMcQhMziZX0N1GPnRKy0AupuP5KR1+iDjKgLWM8DhM5MeVcWVBfqAkd3Mm
h29zxeqEfKtQxxZJIb/8ypKoto3bIA7X9N9ln9+cw37/d5sM1RHvyZlif096LAyo
ufuW6CluSh1+7A5mzD+ymN+5GBWjjg/B2MNapm9EljJ04XqwUiD2SluEcFCaEu+j
w/kzxU6fuCD1YNkO7Sd1yoQSRDSa9pgwwrnbnSmw4Tnbu/R4pg6CoUpZ9AHsHcmk
iHrP4qwJIqYe0ihYFoMoQhBj68nXMpi80hi9vPamD6tOJBmG8NeIZHHmYfRsPhae
+YbNH5oBdZF6nYbb4uP8PfVZY9k+mcxQXQUe6AQ9ABD2k1dXcLcmSgSN02QXFPNB
g/+CYbz0+iPcOg/xpkh2ei7M4jn4Gm1JC2gZZkPyzx2WzGlpZJH7o4e60wFw6/OT
m3BJztjbtrG79mp7cLJCQA5Tq5yFq03KVqwqQnN+Q/40t6WvPKzaBBbROFfh6dds
OiSU2TcG31xpybeqMfJ6LQridUfHYnmqVxLuQbYG/2xmRWOb0+lD2cQK4ZbRXKa1
Hn7AovToThrHbdGP4DV+yuT57/THQ3nzJyD9uuEMd2990m+vUbEvEkIla/Beihqv
KytD0/4XfJW/kUXKt89gaazlCkvJe526Tz+zYLS5rcD+AhpWzaSnksnW4FPrSyXv
skofXN4BChYLQpzyQH8LUmoN+LyfM5RttqemDt3w8iRqbsoYNmrEPq89IgZAEOJS
exSN3+VsjpWDYVw1NdOPE12/ZKzZZdcWQKmXkdPM+OJ+OCWM/TY2YIlB5RY67C+U
VuoxId+PC82zSz2FhaljPPjLYQmatHHXq7Cc97RmCZ6iEwX8Pwdk1ztble3H5kdn
EkTrtcEgnbkYoe+wh10D1UfTxv6DGXdQ5j5mKNVx727AQC69o2qt+YUMR391hftB
H02QUIKjaMO5f3ImjEHF32DRB8TqxJsZwlHYX69eAlvnNc3L4bXhizktQCXSiTyv
1dpEIoH863VGHdWBwbKgFju5TgfSTMV+fGbgpiqCH9W8d0DLL5i1SxYw8uhuif8I
d/Yo1dZA63EGYAAVYdRHvurPupL56AzW89ud2e2c7Pg/q4MWGi035v/JV0j+UOHt
wZagxzgHcLS9gIjvLFCzfWQfoauwxTqed2Z8y+ri4fl3aJ2RRynNWsdVGSbvGEYB
BMI30WWdpL3W2FIQuNBrDGPZNNAxV+m9DG+IxLqbmeXG77iB8J0sHgdywS9L9Fh0
D6wmzDiHtR8C/XOodw5qzHkStPxBXRH/X/K0UJ83ic6Wyq+00H+H21MSuzmHW7HX
lfM1cetp0+dCt77SZ6RD6uCnH4SXQXPzIVgwzLAZARFHH+M27O9jGhmuQQk7IGSF
PQfJ6h3tkBd2vF8XVBoW1Cz/pthLumzx8U6nup/QDN2o2Q9Hc+3kMAvKcuMkOML2
Z2qxbHjKgUVzsD2PGXdw/V6SQOYa6ae2dtmintLsi6i1YvKC23NFF7jT3+kvDtZF
sL9Vovc2bWQ5JtMlnsEN8NCMHUHkV/jcx/CFIP+ndMcRsAPs4Fd1stPAsTqIcMmt
sAsJD1zToY/XPdNICbUg57xRxvbyq1oEL4uQPAWGesulCceow2vcX9rEMuGVebZE
FYjMXaqWgqgwEJoAdPzHuNWpcYQI3EdeJdazVf1x24uI5R6BRK/fyXQSR172CQ3M
UpESxPeMRhIXMgKoYhk7Mpe136RbfwIEmDaRdPeVKwn/euLMeWgxPWXbgzZLSGQD
raW0uSEyZr3dvBHqaO3SJoBax2D8rR8TEvlfBuRM990G/cux+srWH+/r6MB+Ycyw
wI2/BG939aUu8/Q4zRI+Sg4GRY69LMKjLa9IUKfhN5bIWvf34ZLuW5os0nZt0zD+
u409PQJtn2gos5Td/PFM7sY7zeA0USKw9ZUAzCcC7k9p0BjBYnin3aeY4UioqADc
Y4evrQjc5vYDYeYIzdLmI6kCO4M6bz0kPPMr3dBtj9qYem2S+5UV/Z/gN4oCgwft
faCvJlvQuDhdMO0aS9KGa5rdYo/LWhV+a+WDAmQj70Fg11e9ofCcIvjAVuX8VmLb
BI/X3dYQiNEAhSUQysNf/PO86IQvqUiOU1nxObtRPPhuenA31EqLzMgxa5gjjZ7e
2xnXw46wvEoO/wWkow6iYLH1oJ/Jm2Vt/DqN6O6L5mAVYa5FguOQXTW7RsL/LTgW
eBpwjP7xKyUflVACreH1Z5+E3HlEagfdbee9UHP2c8r86qrbfeMA3xb+zNCZ/7Dt
+En9WW6bCS8jSpAZIM8q1bXaK442yWhbUbwAr/QnEVcaFXZemlMIrhal8gg5SNTt
DQaVMPFBSSW9TGa0dVXN2n0XfSBoN/BNHX6XFoTwvlKJLPrXMo21jxa/5GfM4RJs
uVg/UroBEHpcTfo8qqySvqySzvz7morOAznjYBGAmB26HGqSVssCDZGI5jqnvx4/
iKzl4LvSr2BhMHAv5gI2RhH9HXDiOG5gH2nZc1XzqBiKb1+bcizB7k09YIF28hGQ
Hzph2Wrnm2xTlP5O/DGucTjCUDa3s4tZZMPUHazB9ynj+ln2uNdGPE6u/TpPKnGX
ugQLbCVb2+9T2sGNoBAwQESBjcepZC/2+dcfk3VBHnJT/gsbPS8IO5C75Ji1g0MF
kqXq2fOy7ctOEnov0YauSllx6ZbuzWirlqJAr+O+w4B9g2eVQDulWQC3JIqQSgmT
ZWZ/Yz8apbUxJVRwksgamyzo2PBAIlhhWYOGZtOsybsSR/tIPtJkK/gQLZD1U1FT
KACin08L2SLn4qeeEYtyR6c5gNNClxp6kFOzfZg4fMGSgA6fEHVyXzp7I5XeQZql
vDr4f6GR6ECkvH/2zzQpR4FwmrtDw9Nf9xor6mZUYxuMMjaUik4qhZ2UeTARzIZ7
oOL9uvZPKy1fNqkrqV9Ya2s6LDrAT06AN8DbFAMArgsFW+Wjdr4kmptxabOHDAf3
yuLk/x2sEiWOE8FdSH4eWlTluH36h/Awhtp1a8LEiYX8utf2UpB+dK4WDY2fwnTX
br9f3JZ6CCWvC8YEcisYQiMdLRhjSUKVlCxCF0HAcGz8u7oTPCo/F1R2QMxHIaIb
P41YVBWsTA2bRcJOp2aW3grOPzL4/6OzEL7kuuMZkvvTES9/0ifUvqOPddmdzhXm
rbnPB6w3fhQBYd8spqo23dbLjiZ9PAUpPUwRz41coxz278Sqr1c8TyyT4HibE2ye
QtlCZ9pGAYVSZnVnyisY5QUZ5v563yjlQ9PIPviX6yJyscKPkZRciKgmltq1Kabl
NFm62fDRSR0mrw+XbGSrdebkmwsREfusHKRfSzA9Trlqf/1IUribQnceTiznIwaH
5DmCe9QypBc8VZ3Kr39k6aiD8t2Bk4s2iDQRuOhjp4Nk+CzoB7BsvLQayQMKU8lm
kW6ZYYfcbkN9X7wbjrdq+Dcq7hPfDGSqPQ1y5tPbkZyeKlXAqpfFnC75hH54E8kG
O8NgjIkRPw6LpMz9h+9U4ky2f1YEs1ewCt8WJhklFwZV7JkR4yeTgTFVkJVk0Ux+
E0pSym0YxEQo1QmRysmY2/nmO7ifLAP6sVJqFEPRhmTDA7llXO0xEtuUNIIvl852
cCnIEpkxjkijrfk7KmqiQ7DiYxEr4JJ+SlBfL/s9SO4y7L6EyPQQtn7+UXaCXZaz
QLSIKc4mAE5oVJ6wW3t6fAq/ePbh+Nd9/Ot+fFL12P0KOmHer+gCi+ZK0ZB0hRma
GoLZwWrTxxBqSL2WWag/Bz4VqLEAJFsInC0reiRuFfvMGKYUW04Es5eBDIvdE/ha
im3fMRaS+0U5Vv2nN0cHIJ5Zd7TGs3WOOQKGuh1BQqbVbQbaGx1xj5JEkTeLrmNe
16e11JjBSAJXxZZqOo4+J+nkZvoEY6HP9hfMGTh5wkNoUTvIbGZ1GALrXUS3NcZS
FftWBGOKMgu4RSzyFgE1LWG/EGcx6RYwCo8njk1b7OxrrK6ly6kgsxuQYP86yndV
0EotBrG1V7Y3OHloGu5CODLOdPBBTELnZ61Y++s0pr7CzQ+C7fxgryODnDKpTrct
odGpYumiY4vuPJbZa6dyQZOCMlyiwSmTwOzSXWxJLzZuklehs8PWyhs7EDvMC+FZ
iNLas3RyrOz4tw7HYfChO7+szuSNWFU7elUkH9tCmpVyDx2K+OZWDsBsVb4LVYJR
2eHaX1ovV50sRiWiH8lYywI38dN0HU5aW0wr7yAr7it1EfL8BEREp3sy2IVrEiT7
jWrSxVY5TqaHon+Amd1Wyn5ML+C7PQAuMyXetjJ4jNdoUSx4zQzT2gUttGD1gtw2
ULv31BhMaaIBLXmz4DGNjZxo7ocUdt2liBlF7E7b49M=
`protect END_PROTECTED
