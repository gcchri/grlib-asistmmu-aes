`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e85pBJS44VGuOEhhULcdkhsxaif+5KRiVuRnAI2drkyDyfC441XpWh4I79RCD2Zu
lwBlwKtFeJa1kxlBQHySKKJv15HlhkL1pUbt/iV4eaZ2N7FEf3cLtWGODwOIM+uL
f1B6jg6nSNk34FUnz5uR2xqLUTmjXLPUJQEcsW9At93ccQtb/YWx2BzEnS6PbtUb
FuOSFKl00yZhD3KNLBYfwNBAymGjESUJmwbCzhPcLI00gFx0IVp1Ig1xj6ZxHy55
H2+pxx4RQ7B+0D2ur9qIvwVniKc1A+Uf4xzXKsrNXkfi604yaRxGiwZBYzFiPRtb
uH/wmzmK9NsjJhGjGNksb8cb5ijQtzPNpQSD8gFtw0kH2yy9batald9ZADLRTrqs
g4pNIhYd5mRYlVAW+OixXmYNOU78ZxXW9Hs+L+QDti8T7PL13aSfzaudaKBE+fNm
sNaIAF5QgsbgHx4XN1gbPVTvAWRYxVhheu9JnBiz+8s=
`protect END_PROTECTED
