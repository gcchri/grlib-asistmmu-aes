`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lQzyR/WFIr0Ep5pJSu5zaOIysS4jepHCGgT9KtbJ48UbXiHG5cg5+84Ui+FJ2SXc
lTWzTwe26kHHQ54n53mt8X6BvI4XIQJoN5a6hEg4p57lI5nyHliCREFbLnU8mlLw
lsG+ueMHyqGdAvpt13hbyi6Xe4aVUWKDVmTIcdzuKk91s+DO1Iiaez3dWkI8+yTn
QItG/QSAW1UOBiktzkMpOY62Z1xzyqJKcGTJonLo/9egC6KScnfolkXi2Je/bhCt
qUjaezKFUZDQlIkmYrpq+tp5hB4s4DHjbeC6Yh3VVgPEFRW7F7YQZOvL08vvjKb1
vX0GPsy16cc9ADzPG7/+uKD4irB8KUbdFbA6U8lgdeyX8TtgCKDRx5jVbsqTwh0k
0GKpRtOWlamsBE/+8l275becQ2U59TkW55L/zZoJoqz3J2kAkY9gVuYxDEzkVrxo
2h5l3FHF3+YuBJVOkEGwe47TvZ6ZZdYApZIeeKZ12mMSiUMW/ArFtSNVaIT5yvJI
aiwCGD5am9qkHbsah591d1nTQxTjUx3YHUhL6Czo/3zrQC00ehnMq+2DFgKJGGu7
nxpml3mZPGpu0HhnZH3cYs8MmSNJ9EdVhtEE3JOGm/8yJ38tTbR1GhPkQ/4x996Z
Cgl7cM9nJaZrnW5kUNxsyZ3LczeUw7pP8fyX4pUimrUa7tg8TIlurhzmnq6daQZS
eK9G/OP3IPFASKnfbtwUIwlnbvbwtO50GgteOTjZl6GISyr7ep9kLvgvMJ2HMRhz
ggiEzo65FxyDPhdkKQE5VBrOZPwByd1LvVQLQJEHb/gCjzOvvVV0CR5x8h1tpf2c
s/JmN689mvFcQADGdqpfxM5qIZYwFOvr+/cxde9VJmHpBU4zJ64Q4BCAOECkdx2X
yX3+sNVHiuNb6wour2bFB2jysjWqu4jB1FDgkYpyg2ObuwymwXkNJOxJYm4gHDyQ
+FW00BzkT524w+8s9Y4SBqjgvvN0XkyMH3pRZGx9V7fpcBDjnAM0lWdBMqNx21+L
byssgfNIk+EnKsF2jxqRQwptvnpAZbN61MMk5pTgMuC/wmLpymaZBGVfT3pLSQoQ
aQE3yGgCdGt3mVM/q6Qj8QiUmmDbMjqsywBlMoAZXLTXj6Vp8/sKQXJ7OMkI3bpB
Ki4Iv8kGLncZtdlmuUNSHrJZXKjuEPaD+hTQTVT5yBd3Ik4UFYjpLS4XoNjrUGS1
xsyLEh0R9FtBGtFUTRadFKVDIh8eGf/iic6etBU2GhC2f/fjYnUGQG64TC2K3lyN
+v1N/5kQ5Qd5amQzFMglJ8I/PLTua8XLp+Tok4voUtkZkRJUCGmL1ZY3GMzaWccF
zHxVmwK+6pW/INq42QT9ruWdOHdTBOUs6os6QPme2aUP3u6ZYFXAwY7JsbhNsniI
QXb9OWV5lDQrSt2yymow3MfcUb5LOxQNNW3uQpWjjbP68S2MLGpuRfBveBnzgVqK
MlG0DZA+czaOqzRW+5bkaIEiSQ24MdPl1U8JmlbsViT/0XRHMyFiXuSp9mFyCyoH
/JYFksjf2KHFIxkLKkuNz76cin/Gy/zmy9RHQa3OJQ653PqvlA0sjEuKE5KLONOP
OvUxYJCU+deLNIZbNY18VX3cHUXHg0TCv1dYANJ3vGV5gYfZIfaBflyLglpnP5Ye
94IaQL60+8/EESVsoR+2Zw==
`protect END_PROTECTED
