`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0BH2PEUt8tUT6EQ1WnZcYogVudrdae2GX7dD9Zqn+hpMrqxA/NM//lGwP9+8O2UU
UaFY4rCt7TNIzjAT/hz2UY6KC04oKILfXC4bTExOXooIbujKc7wU/4cW7mXyXxWD
Wm/aBzMsLjvni8qFTZaYWTcsUFdiUw01xISu4WLsONQ6HHAFANlakdAAnUHYFiLU
NlUqY5sRl6EoViCrF/vy9kIbPjCUdAf+TKoRiFaTaIxGxcbbajXl4VU7fPkQjged
tfcHkl8she2lZE0Q8vYb7gRD0MfKW96Q2rgqbMmVMgI27Jqcj8ed+Qj7MbWxWCWj
U5wDpLNi8sSPuEsB/FggL3DYz67KeQlgQtTr1ZfWriyxq9kh/sJ7qNiyAyNfyx//
`protect END_PROTECTED
