`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DAU1Q5zmbXLk/yViJrRV9jPB9G2yBynaD7tu25wyC4lNkllSuLhZVCLsHyIQKzP3
0tZfy+MV4jBQWMu5/bvY6ELNV7XF0a7MHGvhz9SoUm8ZF+nCoJlG8LTIpWnrX6Hp
6uh3sy0Pg4iTWTMRTJszeeOGkrpfBuMORqCtylhHnZTmI0Tm1mLMkCPmihyGswjL
LeMW5W+8ZZDBWl3jxIWkb+d7uDsGh3TQD/a19WB6Jbc72zrJWFwACoQ83JGjheFP
CwXTDpfRI6YNQJpXCaDn06oryug10w+t4in5KRD4cGnLVAImY6r74xrfE+xNFLmi
+VkVKcq8OAg78CX83SLIVg==
`protect END_PROTECTED
