`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Oko/dig6nyBKkAzzW10DTGChDt7JAqTYvIrwyeWH4uLj+s9Dqs2A0GXon6DUwwP
M+yMylkvoqlYY3rzqJDU9WlMeErvj1z+iBJplCVT0rfpFPBB7I151sigBYZmBl3l
JNVhKZECuLdZQ8QpAQwrCGzS7SKE0YA9GDKguoo10lKzHWbv3ny7n9OiaVXLt8ug
hLpIbNGygarYu5Um7YwIaM7yCgzTei+EsLyRXLtXt1Omn4EXx5shFogIQq9sEeBX
MDazqzRHHZp9DPI73sg93A==
`protect END_PROTECTED
