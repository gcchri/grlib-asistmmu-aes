`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hUsuCGZxpNnuiRBN8PTJyVF2pDdo9DgpnT5Zb9iaFnMXM9nW77t+VoKK+TVdxJ34
pu9G9kxroOnGMVvW/lCeiMYi/U8hmGnNXg0jPfCM6GEdAv7G0O6pZ/mAzckJXDXI
Pv7XSQgFtN6dLqRUBilL9GNqFYoz2/A1UlDb21WW6EHdtyRI1eUBZ2tAKaBMijJR
dMBLGLyBTei/w0Cm+eJgABfA0Hyr0stYtfGGoxiiCGOypHB40Swe4Mu8i0DRgEr4
xcWgeAdGSCbPyxeOTkNRPrBpDv1F+R4IJPfh5Fd8OqRm1iIqwU8pTreVXARdrwT9
c1QW/X+4rAXh8WHOmNQXkcGVJeWY6qJ0fvpHeuuu+Z6jCn7xxopdjR5R23mVe0+U
hbTo5sIdI7i3/uEb5m8+PdEDkJZYvjv8djgKLmy5N/dBPYIPEQMaJW3eDCJK9xEn
fe4wru1ND00foif7U6D4Zlqp/1wosG096VBrVd4yn1+2nvzRkfted+Na4PHtUXQ1
ac6svZu/6a7iFRZwCKJdltLSkm/SHDma90R9HRNcniCkvTdCmJ52KMRl2x6GJDpp
geVFqtodhKOOdHAnzbjGfEB428HqpoM/L1YjqQxsqJrJ4hG/hAfbBH3ryKRDjTI2
KcNlfGE8qup1TpLbd7TuZta9V5FUChqOHj75wlafutci5Y7dRGHwgXHMQ1DgbrCA
F8RQEO5JqqxOdxrIFTuXiDqaZHTfbPslODiZGuwnvRDg+isAYjV4Vo5q1JFj74wr
LA7W0EH8hP/8eUs3nxg8DSeqGhG0w9T1A6cx2/krDfbay1u9ZoXAXCyrXa96Iicp
tmLcMAfMaITkjzJM+4U+f0R3l8GOKUhvOJ6GjQK8SdzqDBF/cxI75GuUlfvclGKz
cvIfbQb5Yw3ttwvWRJYDvw==
`protect END_PROTECTED
