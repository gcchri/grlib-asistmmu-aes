`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6I6B0vSnsaZlnK4XW4mWqw8uHJEV52emmnR3l1oB3jx54RuY1UKgbuea7apYaKom
rVHgs62zIBdzQeJ6uK8edPH1ujX9nlIQ5X6aISXkNjMsIL6J4xaf0ny0GJCXIiHa
wlNnNblxwzx9zJlu3VA1haeSSYlj2RzK/ZM1IajOPz4uLmH83zyZJuvtfkMcIvlr
4lq1Oj1XGXqI+Zv9Q7HCA4M2J37sLc3gieqxHIOxZlhImSHalIWTQyhAwaEHdstn
DoB7egLy2xCHQYZpkbHAjvR9NbewBDbhm4vaPt7ZaGRm2qO9g0DifT6kmCvnNYN0
2H4NBXwHD9eQx5TEfAYvbXGP5Izaynr/IiOAKvCOHKmvFYoLNwNNqzIsSQp2TFY2
eee+cPgS8VuuLpjQdWP5sVH2Oq8LmMb7bPuC8Zdvhf3UzIbGwMZHE+cXCI6q0lAa
mYLSYvqoQHuO2PZXT/UsXg==
`protect END_PROTECTED
