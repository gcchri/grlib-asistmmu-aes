`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XupZcUfFTCfYJTusSJUBFOCMGl8JwmBfcgLGvpbggZiTyrXX+E49irBgkkp9yyks
EOSQlefXK7EC78BJ8bPHcHnYI4t/Ck5nYEbt9/Zq8wtusux1m+wPX7ej9PIAvgbn
9p1fFmD+AVUQrkklu/RIwr2M0k/p3RAtE9UyDhuA4uquZJwsGnfNmkS0ZfSNC/Eg
tgP8eT3s0jBWLDjdUrcJSrqky8x3SVWdNakdp7aeRuVLQbv5yjQvd/99cgKajVZv
5cPEGUU/2Lu3xqA0xJcpVzeySyYqdAtNzq2MNQCpE1YsviIgl3Mb4OnZnYsWWOpY
WXiwij+BqZ7Dn+wiclfnWBnLnYUe7+onrZn4YKeexD6XC+eRckk5EbXNwYtygeTt
nqteWdenWGh5JY/JcX7qy38CUiN95enmqQ0Sad+kJX4WdK9NTYFQiYQPMhxv8ZCu
`protect END_PROTECTED
