`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3S6ab/MV4kXsiNzuTFY6oeOA1mh+hGyXagcYw0mPOBafbW6TxyQ13Vz4d9sQ7RON
V/QF+TG8g+auuchvPYTMX0VVti0NX6lu+2uHj8FYXfgZWOBu+XDhNL0iD1I1hOs9
6ENSPRAfWW+xUNjQLvEeBhVnGgGdgj2dtjstCAa3UAGNNHMZGvrHo6Kg3H2I4t+0
Po31MfDljYkio93zIItLttLq5wotEVQF9uSy6UdWFbfiYhvX3AlEOZJiUqB8ZwBW
nVhSnCwKPQuWG8SUdpcUVf2deM6WkZZS7SYryOnQcEcPssqf354Ob1FQiRs0imof
Fo1FPP1+1ZskgfXAo8VWCA==
`protect END_PROTECTED
