`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EiDrvy/wD2FCgYfAVhQHIHSp997XOaNzhcxmbowAeBX9iCsYKXfJTpQTNMQDw2vS
xw5cvA95V6/Ez2o0VRwf5XOx5AgJTueHHBT/ZQo2eWQxnqflg3rtJEcrvO6bUY3F
SICOpOUpsKmy9in1rFb/ETacItIaShnTDX0MUqDFAc7w4PnEdkd1ZvyD9+4YLf4n
mZ0yVM3JoQKnoIES5LSH8CXPgvZExZRSEgrj2JHHREbcvs3bBUTgGMMigf1aI8lJ
6+/ArCT3NOOUQVA//ffiRg==
`protect END_PROTECTED
