`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hkrP9fXtZm59AABhcbE+sKXlmqTlE80qcx+rvJbIvPx4I7RGa02ZVBVKVt+1gona
zqC58tmr5shnjJEQ5mNyBEBM8DC2ioW821Z+BAvfOaYNLLSwjTNHhs+hWVWSt32H
wGuFwmSKE/SUqnyz+Bpr9wi92oNZIZGnZdN6BOAvYPxrmBUk4Cd0k9X3VLEHUG2j
0jkDLYnnI2kLy4oQ+S2dAM6+S1bkZBsqwMRox3R5hkNd2mxrx9GeohFAYqBB2lmV
zyqqE/SuTcrJqn6bryj7V66GaEwgi9rA0gblvtqqfW3oQj8OrA9ANePT3gtJISLS
ASZilpFGs5Be8XUOBvRXMA==
`protect END_PROTECTED
