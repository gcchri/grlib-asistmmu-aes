`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s2EOPInmiBeh3xYic7DaQ+wDssrzHLq1H9ad96UBN8x2mMTS9r5S4nfil0uWU28C
s3pXWm28KNpyCVZvnW8KPE4Lqp2wN9uEIVtQSXNYVN0pYzBMQiWVf8NkZp5go7IN
rSKRY1NzRewXLEGxDuTGxd38Ur1UshcVMRxYIpTl2J1ovA1S9zMID1WoBDY01QIR
txG8BU9k002Pt5PUsYYuaiqeOC8S3pkct4YVjOr89xX3lBuEarNvl/M2lczWpzzb
/b8g6lMpn1OOu944UsZyLlhoYg2m0A7ndy7zdTJ1UFWZq2tTpULmfrNrLTCI68+L
cjLMe2Si04ihNXtgEwn5motq21V6QlL9V4dB4ONbdyaRxq4BLE12mlXdtjoBxq9w
xkAMca702JtXzJZ0pCgzJw==
`protect END_PROTECTED
