`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IR4sZkYNyS6K8kqd+sZi7LLMu/tzyCeB12jp9jIQu3lJaVbmTc1f2UXgP7CQjO1e
rAFuLGOXnjd+f4qQ98k2ei6N4RM/gkFURsBIaC8x8QpyIcPa0n0WUvu5A24s0uNN
VyDPxREc8H4PSKickF3/m0cLb7AfXyfW1TGGNCarNkIYDZlldkBvDKaeM0CvuuM+
KwcmaYqsLf9gG9xyfcod050oi+vbn+BTW7LL61U47ZqiRUpEv/Rxy3jWXVAxQ4hO
TKQlxe+zu892nu90iKBTR5mLWCbPFx7NiNRttpa1HcjtI6DqffudGR2LnPhm7L/J
MssqHYgpxSggOs23LlXLeeZMyp489G1gOFI/aSHa7XKBGwA4S6j4LGQ/B66hGbxV
kAbXchHrv4VSrZr88R4Lt2nY2gP0J9QCrwT+KhJQVnnvcQaii2yUJqSwXBL3tk/N
1ye5g5rm7zEQulNqZ0jyN775ASsXbEDO77zCuMs0QS0eUtbFmqSdbx2gmDjsWgOK
CkSkv1dKx8zC+sMi3See/z4Aus+5nsPK7oz5/diLdf1cfPr4udD8zgUQiDDCzQop
HuqwN9Gx/05in7rl1JK2h8t+pKkiVP1ojAd1wfva8nwQ0GhtNubqRwo5ylFEJjpD
iKautsYh3FYJ2/QgvLQPE3K+n4f+7jLEMPhvVD/mJ+6K58GVGK6+7MNetiVt8tJY
cvcDcxaZwNwo/YrWv4/d3R5fa5ZtwnoyDgY71hg9zD94R1PFm9k0/SenQdLFkFA0
KmTv6h9gMiuUHmMsiGgsqTNef2esepqvhCC3i5Y3/Fx2x3C4+Op7SwUb1b6Y/iPH
/Kx31oTLD2uQbXLkF2VwgQZmRVnSwdEm78Lk7Bp2jj51gi6Fj1eZa7grNPLIYg3r
nvSJGfnxV1rZoeZ3HtPHT1La37jtGlHL1mFlqrDC1HNu0qYjZQp/o2267LTuWrX0
kFyCtHDySWulDjM2T1iXjA6RaXEY31cayxeL4eJKr3jbChN1Z+ueMPLYW6g+Kxs9
4lcNnjWT/BrRLaZWOBH2HNgipxB4DHUdZW34T3cPgnXhuTETCSnZ5x3ME0TXTuMf
6PoHqNHGUqNlnX2arbnClDdQbArTbRBYT80mE2Oa8hSzv5vXUvPoZVIKKSU2HFgt
4JASpNKPDjz1nn8ueRkqDvopsMdXYtgeNle++LZ9Qu40cUPnkxL/EWO2CzkEK9cf
Ojo4noMoL7eE+3bCmM7O4nNymCOhbDtzfBAaeUwhuzKTz1cDJTIkRFa/wjMvuOLB
89HZPbuAlM4j4v5lZdyi5L8TZLsjj/ywdmfZ0CUrfLH6Shsz+4yYwgKynx6NrYrm
2gFxNK6N+e4rEu5vCrSfmWWTtFFpWOiyWXVZlsYVistRcAok4+X6XkRkpmKj2I0X
YKQuPiPeKA90Z02XL2cCM5qcnJPU32ySJefgQmfmWMSWj4bWum3T4zP//YTPhvuh
0BPxO8w1+ITeme5D7d1NsXlpsItmSItaUQiItRj2vOqiMMOP+t3coheYkS9Hn4OC
BVWIExFZuU8qhaVTFX4chJA2KknIV+X61yYl7OSzBgO7uGNFFVHCvZ+EbafeuaQp
4yFpV9MTZPu2mCKqglcGdGXfFF689/1aWaQf1+kcXvtlgV/D7nSyh+eSqcQ9TK2+
R3D/Mu1cb+06iWBekdKIrGktk1AP5ThS9ZBSdJDF5oXlaD2tzAZw+gf2dbO+MR77
jrallB/NXFtv1/4kYc1/iSUDlvNyxvosF41npfU+j6+p6HglC3RVJrcalm9bDUX6
/ulo+7YSPXV1f3JiediEOiNpkb11/xKoIcmV/QFUMzeZgd6ybbNUe1wDhTeAm18q
jOtft1kzktSBG8fE2ZE1UNXCzct3GgCWa86EHnIN1RqCdPOgQ0/JxMfPxBHdw79R
50i1UiZl2Uk98LRNjw4dLn3xwhn6FB+vGzR3BHAkqJXyqSuZVoEMzlc9Ugw8uJKK
ISJsjru7C+2mzP78MGEDbu488OQ8RmS/bDoLU6jXoI9YJwr6z/Z9wUXN5EWD1btl
KgZ+wVFkFE79PW4+TfD3XouiEwiQ+2V5zkKg9iIQ1xfK6iKU8bdbF5oSpdyNMAVd
vZgLOM4bsyRV+6H7gY5M9POGHqk1i/6ygv1r7iSV6zPxrGmMRNFrMOFSpb2H4ZIF
swfIESUQFyJHa71ngBbqTr0XMGOZbjQBnGf8uq/iyzeohC4u3mnP+gaexIz6mvgZ
9C7MO0XwoGGcdOjgC0Uvy0BBEbzozvu6SfbnVRHvxkunFSXA3t1iT5zLLgX4piJF
6QyBcoBhCIi/uKuNd/RmaYEsP08FxmzVcV3d4p5oy5XS7wB4hXDRkKH2h8GOIMnT
Os0CmqTOPhJp45zaJ6Tgm+YL69M85p8BvNnkOu0m5DKWiHqqgK/zxbJWWh1ThzNq
lDSaURCTVqJXSM3qdlkrFarqix9wEcppSeh1nI61U4cGZC/o1mnt0NLwUjLxLjiu
AWYghVJVO88A1uKk9TNqR5/wwpelCqgU1nMONpsy5K7PZxpGIwQcudAU5UTKhBQy
4m4eOc9UjwjD5qAnob4krG417wUYXA3uJHhu68ghvH1M8pYyw1JHyxV1lDqtaclN
p/WzhU0mkfZPetUbxnj872tuR0lvbtT1jhv/gxkqswQo+qLWDk3XHHktw3Iu1FCq
14+WLmV8fyTAenLVSw04n1/BzFWstph7za69LCmNIutQOOXx1Tg2Kmvcn0hv2y0B
t3ccAEWd462AbXjCYxbwmZ+0fuunYjTjjE3zO6kw+EG3LYJb7NloSQ9NVoZIBTb8
/ooQYOWAsLridm6J11SZqq932E8CJiMoNJM+b7JMJxp6er1dTFg75peO7jPo4hw8
If1uvV0uUp2cSNkYvpmG6eV4ErPTEMBSj4qCDDdgK6srdWSBAs4cXjytUoZ7hDtf
PyOnEstBUhcaqMRF2iAz2ByKcKmAh9dfvC5QE75UuUWKss0MACBqjs03f2o7vcM0
/yyDFMM5Rq/lxqUM1ulq/AO2rU2o/YftwqRgzxCRQNlYjf+tSscv/36ZWUb3Nl/i
FdBPihXyKopXYCEJsTI00AGXHhraM+e2DGpYSuYljMF4p7igG2Qh3B4OkhJEewrq
88TXtNxVdtK3jnvi8g4tCPHujswrRBNUQkH9hUzpQHKlgtYeAh85mVNSWkkxS+yT
Qle/E6tPqMjQvvqS/J3r4Aqiz5C6pAvGYBVv0gx6Xan9Vvz50qwzQ3Yn3RXT49QX
PtmD2dUFRe4Kqb4UJbimSsAnbPagV0dO2JBpkGfHfBEsNqG4Xup+f5QwinzKtmMM
D03DcDkhgJg66PkuoKWReQMppQwh1Jz8BojsuaBIMOfwBNEsb4a1Tc8SJpE/i2Ki
ghqqVpQlmxtb+ZLvZAgCGQ+PAqmqtbiYVSxbNtC6X4KsPQRjVSrUAuXqKzJMcQmD
ymHKay3xM6PFTJ+i/H+0fnhqqavFmBPAK4ezgMXhpXCjGNiD/MalrF4F1NPorT+n
ohpjzQHKKMBr652eQ0c5/Bd6jPr+705UlGIeL4HFEU6YOGzOaOseN5f4TaT/I1gc
1gb14qtO62qOuTfiC1Ud003knZ3JGHCxqwNbJG9W6ofsxCINfBVzzguf6w0+XJ2C
e45EYA+Vitx5O7jqUQDEbKeHL/tv6sw9V4pO8YWmO367tndFgnDpAwWjR0OiaIbx
yDRSbhdiw7v/sSScyDc9649TkVRCW9C7X7z7T9JQBXHxoUcaUd3EUyQOULF10AGo
yX4QyxSPZPjv37ZzavkoE+R6PWokTXDGSWkHo1kUHa4AaGRTiRZAJR8+M9pdElvT
7x1ZWuFdPex1yaa5BVAza2/bMMEuVhy/TiuU1hiWVKJuhSr15wHbG+2jBM99R7go
BZAKjVWP51WOuvO6TbSzB/UlXMpllWB69HjqDkGNTQkue2eCCr0Z7wKfX4g+GSfi
5hXshnPUBQcp3wnsyHPM1TE2Clsmqb15V6wdTHh00/2Ipc9cKoghaI6HyX2OxQQ1
2zVl7j4fT9TcjrjNGmpU8QGi1XMllgc/BMj0uQAKOLBCmsGe8RZ6dk5e68YFu3oi
0WQ8n04umxSdczrYQhtg2AEGrWOjZYuvHwnFFeB6fvQsNYfR25NnaYFTJ/b6dJXW
ZtOK+i5LEfYkBCp5G1+8g4hrA9DY2EZ2+dsa0LZcYEuHbzaWYwx6mBlfwSpwfk+Y
+CyEt+ty2e8nQcqWFoiRbnhcCgvdrdMWlcIo5WivEapTNE6ektw6YLHVlac+iv6P
kK5WfdTAMRv45c7u+YrAlMUdYEbJFbk8dPp//sE2yuoLFnEfPUSbfMI1f3Rvm6Jo
/YsTcewUBIY9jE87x9XnoTDM4vkZC4fBIh7faXxc9JKVNQ12DbwLNz9NN1GiAd3n
JqgvzK4CEGMH7QdzC3XeBTmY+x4/q7WYQyQGAxOStIxWIq692Uh5msookjpOJ6bY
OOY9+SXzi5eubOzsuS10myRzKzri2pvMxcky/+SjuHnlosuVUO2Q/cB5xIm9KSKw
8yaVxO6c3Y/qH4L2sF4ky8LAYX+Wbv/ZnGGAz3xoDyyJVPNH5ZerHNWFkCmtI1V8
sunc26PAMYJYcpc1Rw3MDo0xHcq6p90ZCtUkuwOP0MNY/wlq/yUpFOyC7GzFPi29
yXqyYmqZyJeEE+hnUF5NzWG17lmZGxubhdU7m1dmwwM47P3GEjU/fgeGh/37YNit
/Orr+nyOD31GmUcHUzYg8UKuI6+vYVsmfhIRExUla9rnpTJWN5UBwhehCBtX/fJr
/9yk5nt7WRJJk3cN9zAwJtP+bVgnIBcNLCbwobQYeTj5SF1slPMtKRsX5cnhatM9
3Ibt+VY4vVDGByypDrQ5Fk/TSg3hNT+NyL/D/wb2bLdkHldJKqFvmXy04kx1sXAz
TwkBPF0vMlFmfnS8XYcZbrrmQ7AFT6M8dFTG8rl/96VtX1IwRTbBKzg7/Y+u0FFp
8lqkDmQ7Zq/s3pB+aFyfaCjh9fuWs8zsR4JW5QnEFDmf1QrG6k8+DPzq3PeI9W+T
fNriLaON4/4LovGOmN3mB5WEs8W6oTP+ZiWtUK7z9VSyuRJH0W0jr9aUs1SxNE3D
YxcI1FmLa1vZq/LMeAe0PhyMyHqGzF+sCvPaEB+6tTeHi25IHaN5N62fY9AnQhwA
sxKH/3buvfzyFeccLggfdVzVluz+8PeBz9KzhQXQHs9qpez3svUZxfa7i9AMPGOx
Q1BLmTlz2nrevp1Suc3YbqG0WI8JUL1G+pctpHtEQ8FTg4yMMVcaovlhd/fg1NNO
3VXIfVuNQVjUHXyfEmDG7ngtBnhWOggiazemq0dZft9LwbsXfGPbPKwSaePr4MQQ
ixOVcktLMPLAkaAunN+XqpLTB8KgFddg/mVjb4U6Xij7jA0TYVcRQ6ZmzlbVGfsW
iH32prAJXjxyPxGLwCo7SfknVZhonCxUuWoZwpu3q6rXWdtOPYtK3/WOO6Q0zV0J
tysCPJ9Hgs0eAevETWtdxvW/zuAkz5JcFwXs38Eu/W96Gx449jQin2YvZS44Dk5l
gLlo2cdmxhQek09i3eIIZfjqrFx+Lsh5lqll/ySQZWz49lLnv2SKwEuAfWgqKnj0
SMEvhQYWlMGo0DBjJ3et6XHA1PdWknodwkWzUN6pnSCs3j0tfFxkhsgZnzqNTj8S
RXij55ismWOL54LGgaL7Quoi8lAMlY53BPpp+IlV6P5cVhYl6lqa7NVInbeRzJbb
KFMdspDfZ9kv6rmCSYL4St/TzKZ99enuHpcShqykQoYU0c0sHojMeOUKHdOv1Bu3
drRvipdHeOg/xSCHgtlvtw/n1hKcpXPqiUjVFsjBEDBQf81xoQ8/YLibaH3NHMWk
IikoOyDqB4nojws+bDDJ+kD2QnpAFDujanVVuTPXcj9Gv+TxEzdmgmhZGQJ2Fsyh
u8vwnKqbS9LUXw2+b5J+68/t0Njf2djYcKRrgx3WQLCXPBp6Q6j/cYWwPmo/jPap
scVyqOt/LEJCShZyZbAHvve1A7nv/n/K1pbii0H+TL2SmAvSs8ZLKH7S6cqKC3Ri
+6xsKwny+WssZghbpeuahg4sS/XzVvitxGanT/TxwT4BSf9JAVpnc3bFlJML+01U
xZMex03lnEPi8AKflloBal+o5/Ex5ScvcmDs5qxbeLw1zw/n/q3CtAL44gbIApFp
SahMrLtpkPAtqQF/fa7Ms3f+bgAaVboJL9WumBXPuD/8Kz0eozxGasSYxA61czUa
3oEURTey63WcRfX2AKzmoPR3gfDp2nol+G/hg4GLAl6kcQGpWsOZcY/c5b91pnmj
+7JFek4romNqd9b4tpaHEP63QqDKB//dpzFoPKYA/1ZdTs7ob7fda1A9sorWROHf
IM50BRw7JuK8myAIQKiSbIjgm9e20wSoMClR/jon42OiskVRPEw6vLynowW+ME/V
EuzeeJVpqPZ4nL9sk0CcxD+bjVJsbtkugwrxVaSNs+WK6p1i5pCDOQf6XcsIxPCi
DfrJnwrmXCzDnWrurSoqtfsnLh20p2uLDtaWYKwQHgT/DQLKIU8t/KO3InxZ1NtP
dx+7OfUeNdkj0o3H0ZyQYhf6x0HvODTcbYsoU7L4arCpew1FjNfT7CYgGIyX094+
Pic1D+ECwe3F2VSIq0qgiJhoyVkiTlxN31yU7WM1Ut2wJTEvDzktMtvJmeRSGOok
61SW6s00dpRha+ev2LzMQsH8EgXIPDypS4u5V1Q24qkfIR0nSY7DsU83nMEDc1LO
uiGW+ghpgv/5lA5IqjO3/BpmXRHPHTzrpIbbE5O/3Sy7VnEu+UppSjgvAi74Q2Jw
8cqw+RU/J/ZOTBCDFwX5mXMn4qdkjdk61baJoLY/rLVSKHY+04xdQjLKI4T+5gmE
C3yPcX9lnYx6EfoHimwpwHRKZ0Epr+OmHZjfBOu10+W0nuIjc/GDvvGVxINE9M5u
I+B4O/0/56H3Dnayqp191cOuDCtk1Mqqm06GVtbFudquqeb8Xl+Ta5AZMOPEV72F
cFUAhfIv1Y72fralGVc7rB4jOl/0FGTNZ2LJPoDyf6lqBeuQ0UllGEVimAJ5MzNu
WR3H5I04BGt6trXUcK6nj3Kd2OCryQjFVEZ4E7UjW5W3TsSiXtVjdTZ2hEdAKAi0
Wc8W5x0Foh6LOVAc6WZvbLmN8uRzNqgJyfukkKRzpI9xD6bqibQGnAmPM6sTLAqB
XaXaZxuWpkVILqiiakd1uwjsRcibCbWRC+mra3ni6x+J6S/VPBve+4FNRNaISNbK
6bXPJjcyWfQjmWF9U95QHJiu31xX/YR1OxgRRe8g11Arry0LOkHmNW34GpVTv13B
VlQaO2Z2rGwFK0xr2ImmNapUyVlrsMNWjVV+aWT5kLwPXtXfpkmuSgRnicLsJ8o8
EqMDAP001an3ADpfjaZOJ9wesrgla6fmJwHKd4KETXsZwaTww2qXsy9PT33wr5b6
69Fw348ilBkDVtDFXzrsDMCfp57QmSnlNlEuzQmB3aPHcsYvJM3kwKgVNMrDOqNt
UAqJhn3Rr1D2Plv0NRXmwoH8yZHTruJNRCmLUegn4cvJxMNdhOc6RSS6sfcKXqS8
ouAsWXI1rE2kOI63JC1rv2Z/abM3GrWCZvGbfny+PGXrcwK3btTm1E+elkWldCTi
bSHh5VZzOLPWd0mIHCGCn9SOnk7JwwYUcERjSytj0JSajFf8f04RckQiiZOGcCrN
MI7Wi899AzqQpJoHko/uQZ9sZn2JtrSWCN8uMYkT2eBxxMk96CwQt3sgfnvTui/J
1TdQan6WY5DP6S6HMqswU2QDHf6kDKsH7naNWMJFzjyyDsHpU1TuhRx72EToPvEF
pXS43MUK5A+0nAV2ZKNGTscTCKCmS77/YAyMBVlVPyog/Aq2oRQuJoP7vMxrfXhp
asTlyW8z5qZcggkgtqO2gFaEioRBHdydynXYx+64l74PebDomEDbbj3JW0yQSO0y
ccYSdRdcqk7RKgbm+ABhwGOUfu+/su/CHflOQ1AjJhxDw514PmBm1NLPuj2zIYmm
8o8V1OmUtsgY5BbSpxOkqzmKNOBYsT1w36Wjhkh1wCvDSfQ+/w/oPiYYshLq8GFB
LMF6TwLwyQVYpmyYpt2NSS510o3ksbG/RXgS+YwrXNc0Z2q0yJ53bEsWn1waR7OY
lAPO2s916i61SNbK9z75CQjBcI6rlXKZF3/iM+Nohe1oRNNTYKCvInCZzhMf13cH
mx6zUd6q/W57UJmZk7EHhAIEi0zyYssvEWpp4zIswAQ=
`protect END_PROTECTED
