`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XDHx5ExhYpZfbrMzbevQIfqUod8XvkmsICPZTnGXhO/ZsLhv5AoUXKLXD4q9p+u4
jT46C4AhTCsbk3oJQr/9nltfz+W3i0rmQUzVjRIFnAe2mMCHzj+iS1WN++ue02YZ
oIKLfNM35heuQSD4hRysnGyaMd618GSFWfq5EPT15BJWrH78SGUSmxUWlNdM1Oth
iRFeIUS3IfOIsT/b3VubK4MGoakKtzUXKTAtsRvLSgR9ms1RAghZZWEBmEiB+0rB
FeE5Rzn7jm4g4tXWtEDwYJQLtpoDSIg7sioUREFMbMC5h0YmQmphIXcaUCiNqTKR
XlZo71Y8/QMSgsyu+xMSTpsJlxKlEUV74Jq5tgkWOmxKeru8jqBDbeuvsmnwHLmE
YR+7hgT/64ogMOFZydvXagLLQyrOPmPx1FIywjObuBDxzuohWT+v7t2pbusKgj7c
K9lK2m6sfqj7cFB5lgLzyOuoMpn8B8ydPANf9OGb7/cbYhYjUD1QflaKlVSt5U5U
`protect END_PROTECTED
