`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oMSVOSZW7MUUPyRcgopJO3VjnX4D0KjBacipeBiPtKhKV5Ewp8F4dBagyJKnpJns
Z1ojYC/b9wACeErNj2BMZ2+8ppwn1NUevqlziRl6pN6MLYLyoYFYf/mV+ccDet88
Gp+7yLKqKYmJjhAAkRrekGJDWhsF3B8XDliDbBUtrCw7eYDFWc3kc9CSRWS/YAHZ
n0faEu6Bhfk5X231Xpm+xrUOe836LAtuNX3SQpHMsNdduuWiZwpXCjp/DdKQeUVO
80bIAfJ7+xosrYisaTqI70osy2/dWCQkBxuugqWCLPFN7HfaOcHaZh2STm0na3Qk
rceptWlgTVE8I0QdA6EUNA==
`protect END_PROTECTED
