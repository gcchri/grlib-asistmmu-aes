`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HMxUNZsMlsztt2WC5OQATA/2CUEgMbkBlTMu47AlXD60wtslCiIcG3J2F3YLjQQU
XWL6zXvLyKi/b4n/6VxfpMa7kQtqSXkF/1ckeF/gw107YiJed0Z7VVeWdcJoMxUV
FUZzFgqZXRVpLvRtFQjyNL7NV7xZKwaa2N4yQZU8b+zkIdPwDMlFTIfE5uhtatvF
dzIyr3qjK/uaExPvh/Utr25NPtc6YMPbjUkfDKRTBFm1cFO6vD+VJ9aCva7iRZiL
DLQgZsYB1oms9Fuq6Zv3dXz3S4mFS5V7AVnR6zIbyJ5inTTjORO525V38tsTEpb2
uBBg5FVWsT9HYOfECGLeirbug1+M0dzky2ctlsG9jpV0vobNE062li2df4ugv1F5
EdyvVkjXvYwPnvaGCj8Y71pP9lzjOPS8fcPpwwcK4z2uSxAB5gaRJtshzxosVzSz
CBkAjw0EgXkWE+pdmXmkx9SXit3ixl8rdHN+sT1x38V4FXQMKt9ZktqG0JtVM0zf
78onXIp5n4xgpsYhygrRXj8hWP6WMVB5kTunpBg7QPEOScfn401DA8Y7eE/EOJ/o
16C/EBrAVcfwywS7aVdU/53+oDjzj1AQdN9Pn+QAmI2VmAvJZRmDKqaQGc2cgQTJ
l2ZSA1Tfsoq2QBDcWHgftQsxsx3CN82a0gETe3lENB3tbsekX4lUFTPauJhwCs7y
TbOB68bcoxN+RDKM3tOQ+cP0PccOXo86LFVoY/DL5wHD6tI9DZ3a16Pj1HhZ/Fyn
yGe1F3KPvLxMd3z1W5RmLo8n4ueAFBFBoPNZ7r6CpQIdpdcsKWIklrdx85JqrPuz
wp42OFo1g3GWBeDRLsSVM9v4q7+tQNQsFXmoQiOM1O080xyTd1viuvVxgeAIgW0D
eYj0B5Tr3UEkE886qh4jbP9MP/5ZRnXkzqC7cKPGPz32pw/rEY8qKLuSem6cnnqK
`protect END_PROTECTED
