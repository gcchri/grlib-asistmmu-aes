`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BVpODM0RRBjkHYpE7l4o4wqAPhg78SD6YZLb1TNeBYsWiE1te/oJKkAZAjdR1ijp
zfcIJ726X4DKVEBuUg4Pn98xrEXtkcHOjwz7N1wGg5hheDpdrAIpZqw8/g/xtGA6
xoTO7s/dLqWVwOyZQaDXBPjqa6iwCcP/sVLlLmfphOarmK9t15v+Ark7XdmsmE6o
n1iTv0MsC07h1bGmu1K5EQT1dNV8jOLJwDetkLYtHtRRBOc+xHLxSDYmUKMfOWkC
oxBKSrI0ftOcmf2lgwHjyn1TIwRDp7osOx3CFcJhrXH67VHlAWu958rsp7DG25ai
r+Y+ygK8hDLRWA6+fJoFCj2myZJUrPOaQky/0mfxP04n1JAesEHntt0iREmmfeC0
nKgGrPGBxOCw0EJ3X//AFvjjqdGti7pgsge4uE5T1UBCQ4krxbX/0px6vZmBKK+i
+k6AEsx5EUvOsd46IzNriYFQCh2gRFKgdw+1A2CaZXI=
`protect END_PROTECTED
