`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9AnbiJsSZwR38nACvosb4DU9c8zEmrYuhBKc1UGu92go/o2VL3XsTN9Ip2d23eK3
etxCY/v+106L0n9B1mF59JomdrBHJwDCqK2viV2icVsPHoiNECRO5baBqIz1gwDh
YhmztgAgzWYl/Bjx6IqlioDflGg4xEK2163vWhwEPLdPUrvdlGqnmO0H3fP/35Fu
Ya+qLrH4bZ5n9Mbd4f51oHCkfEFqDcgE8tGxkXQRhUlb3ILv22BbyFwD0+Eiz3nH
IMh+VqZnobnkry80NUPRBAhuNCPwxau/+nX7xu1BkuKfio9vpHIXvdPD21cGoxZZ
XWD9DCoTsC+BpMrardqZtA0yLWWFlB+vT2CnuUygNbZqZlDO/FwPzu1SpYzVqDdQ
ikHupdTD77b5KodNTJhNlHhmyAKYJoVgD/woLhSQ9RMEZ7gHBh+N/2dKIWwzXsug
3wEj1rxQyd0j44GXJE/TZFpsX+ajgRFTMs3V/S7fQtGU5lFsO66TcON0h78aCJLT
5CO3sG3CRlTsIwhPBdX768LLoaarcCRVw5f7xeE9T8Dexcf3Gz2RvHl7Qe+sQ/UV
jPBtpJ0vP2k9uQrQgLEQMxZ2DJ5ELboXvN9k97Lo+2jvzYbY56dgkJUYAeQgxazg
ByxDA3KA/N0C6YyTNRwzwFRwz0Yihf0+vKy93DHfF3fsYC4QbLBQN2sPpMu8DSLu
`protect END_PROTECTED
