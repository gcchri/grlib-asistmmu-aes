`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
olBiWjWfEj1RU5cmugq/Yr6LfzHgfl4edo7/6BtcOuDA6rIeMQDplYsPY4FlsDro
bOiePPrEVoeHjG2qgh08aaH3+hVzjwZBWH+gUcs0v0WLnA4qr7H4eMhE+qSkDlQw
9srbUh2WLka4nLoe5GI0nGYcHPbgXZwS7eJA/Ua3F+YG3NJaOKC5DuKPzwQMGAd5
rYzVk+ScTDw4+JW03nn+tAzGRvihX4yaTMjV4ewT75GyLoFs9URig1csKTY7cZNf
mEeuEl60hSpmAlZrevpWMIYlbWKEokVa7X9n1qv8eM4HYvSBoDA0qjsQ3kmYrA61
SlwbIeeHIiI4n1O7ghSuXLfwyF6mZnUuH8sIFsaREXg=
`protect END_PROTECTED
