`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dQ2lqYEX2Q7g1vJ50QI4k7it1murZkJHNF9v3sAy/qFlPx1ZfSwbbdL0GgXIWet1
te208MWCFcohvKDeVdgaw0h4W0y+olif/bjLLQVeppuRbFiXouEPTcUhWd3clwP+
b1RVPqbCPoauKJhn8lGzBfalknUavGX96mPAIDkFNJ/B4vHJyxNsHRqPWl4SYrPu
AySk0UuK2f4j05u6p3Zszf61ErvxlHWWl7qkLR7axv1L56mBd9gnz6WJifwyaVhW
DSV2HZuLlXPSp9/qmPbJlsl+ifcn0DSqk3w8yzQBMxZt2D39+fnQ2MFEAeI6+4Hs
x1OcOTROqcp77BX30YpB3Vk4tvstaHAP04NiM9raKQVl9jhEmBIZSlT4X8UjOCWi
7wrb82D65xaM8j0nPcmRQ3CUmqwOjOtti3OXsWMykr50w7aV8gRf1gKyGJ5nqBnA
IwhuGplHZtR6du/xpklu+kWz5QAeKJzsMDhBfTZzahLc/fbUH1tsFPWqh6GFsakB
T8b0z1niazPAsQ93hQozKNSFxK32pkMsyyQYY0j0I8gRA5UYXiuLhZPmn41jg1H5
AHG59LPfh0Ry9uNqMs4hCcxdvvth1wxZFOe5xNhoZn3bMZIoRufVi/ztC/moZEyA
WEfsFCoMVgzzGIBnk4crwJaN+KRGuiO8YNmZ7sIBCgmuJ12/cphqTXNTkZXaAwM6
33hmeIbsOW2w8mssiNQSpsjDGR3/2VpCOZ6adg5deYbN1U2Hm5uXIzAyEJKrbESi
`protect END_PROTECTED
