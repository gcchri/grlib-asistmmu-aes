`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LyveffRgHGEz9TB+1p8txLx+VwXNjT8rSd/geIEyTlyhVTFlTg2yrsDd1aP6rQsK
AhM6NDm+gSHfouJ8LZcQt2zCTnKoEb53OCtFjJ2zdvUFbXuc6/ZcSL9SmzL2Cbt0
i9hjM9WMnIXQ7M9p0S64ETXvLIpVzXRbS7Ty7upW4mthEf0ew/fTqTZIBMuE0mN+
Q9sYOvtrge+KR0acZlEXJ2nxivoBZIGXrks1uPevgyecGd0ndh+eJveoxDbA9b8A
Im0CsmG4gBjvw6s4KVBUZRJRJyaAZ3k18p6xT8ukpRIH69f4mgDbb3VTMNISA17X
0mFKFQdYkv4vamxyPkEJHoJbGdDouENG0njdz8ngyLhLrapac9DqP/xCPPPUKf3j
pGZo4kLMyrVWW65FmmUasNgWP90sEFSwqx7GEa1YMHm32omfvLalmu/3XerVlX6L
2qDKk88o6xFDqapfmUVBv2vL4pgz6/gCNQyTo/N8FX8pcSpIpsZM7viOaI0NYZJ2
E53hFkWYLykT3NPJfRx35oNoiljHx9RWmq1V0nwNenr0IZpMC9Thyde1qK+hZGYL
ZrHCh7eHtv3HlKC808DMtg==
`protect END_PROTECTED
