`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e7WZTAb3AnWYqYks4+0e3u5Et7lABMJl2RUsIqjstHreoAEjRfESWlCeHbmNw9Ua
vXze/xPeZ4X3qBJnsctFtoZNz96VE2OSvilYDciMH9v67Ps/3Tko/xiFoSCbuZWf
Xve4//NdxAfiD6iaCofbQ3um52AvuugyyeGpnOejvc14XYy65YIdiHB563kOYGW4
76d8tuHE2eR31YEWY1wFxchR3yHJsVIlTYZHrPPCRlm7irBe300bjALrK+E4dRMO
eYUgArT0mDViCZvG9dLV7xds3nH61qnnO+Px2w8wcyTW6oZn1q18NCYbwRYxf136
TfkDuYGNkqPvBOixcWjTLnpOMAGjybJqI5bCbKxNbJGQzR7YvCL/TTTCszColmYh
qs+5k2OhMkwmJEV4RVRMMBvc6nHxQUezBC13BkkVbcf778SDwutTTcZIOdjNmFPT
Z3tkjAvsVPaImQN9RDE6yZzLgfo75PGAZIJ37otp8JY=
`protect END_PROTECTED
