`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BnYF2PhGT4Rg1yV+2nAfpbt2OjOO9K56ICth8CxE/JRCE0JZxNX6zix3DANdsbX5
U+3iE5phBcV+8C3613C1/8YrTBB5WsPA+exy//0KuPwywVLhHAvl5r56VTp7HWOw
UjzpoPT/mOXxIpF0ipRu2sYFU16iPQ6hkzwge0gElwKWH9UFvGkUAuC7ki7O3+Sw
syNAw3gNYwfL5MmlH8DJPSdPc9XrPU4BFiLkQSXBCiPE4ZvA+oc0hT+7Iljz+rNR
wXcEjno2+rfjqs0THLspMzKhQVhzWplTyQBWshL24jyKo/XtWJ6tBoXDe5FZvvPW
6RvkJQxoyU1tTvVxQBTqpIkRBDeqHF9+HfHdlpvdmhK0EEAxSy9ZghcPdjdl4ozm
/YVxlV7fmgVMDE/qQNEch7FpJSFzKUyFXqov43muNPMwELaeQ+E22hHRqayWNlSF
vl6q6oCAmlfEt8lHy9FWPe8JN1zyZaA0rR7775uh4R9TCtVG/85OIw/JzG0Eil3T
NFHDTmJ8bBkXfDS3URTl5cN9xGRlzw50J4t4FFuDJpiujRGtMqYiNqDGygj1esQM
DrlQFXi9O9HizGgeeZjvrrBXSnrO7Kgqfikbcr0C6WThtIzaP+w4F2EZkt9GTtNQ
bRWsIT71dokwEicyliJvdNO3Wh0yAY/QPkctGZSSV7A5ODujTd6piuB4YRnrUNUo
O1v5TSjeg7ZDFIIj9SxN1OuscaOxDAy+40x8IkRhBrd2PlDjBHZvNynRmg3ClQEc
g9sApMIlrXRRnuwRPk1hhTlEJ6aAbySlhA3ZChEWOcMtx0qqt8oMKHOKIk1lbGpN
BjJLtFsSOUBrTVcGg+dBTMAD/ycRVz9eGwMqbh4dXpwL0ab2FkAwWHKLVtlLkyGr
SP4CbWJctxhkflFlk8cDbE68qg6VJPIZGZkg3mXnPSNwfBPSVb7zHVf4yJ8ccy57
HiOVC+Vv5+6aT2qpynFE/YiQyhkEq+BBjuDzAJfU6bsxOnrw+ARpWVz4bicakSeA
0Fknnh+HiDurgqThlBjuX29XCQK047hAeqYVfEdAmvC1Q7A+csjsWyuHkiIBTjO2
5YqFutXDkLvO7nDonTjCUMY7SdxQq47shibK6UOInS6BI0e29zgajDGZXbdLAgna
1Me4FvBnCr6JNmwcQdK0PU+bIUVSNCnWlYZgLthqq29Gz3TEZBEwJEHQ40leg3+K
/6rOaIsI5Cg1EXBebeub+Qxsx3srAkL4VXrng9YXMrsag68lEHRA+jCQXfAmSznI
ytMFSBfOObnQQ69MTbCnhyh7svmmXd33TAsdwkOApe3sHSCu2HjPWKnxDt5yNdwf
pwrs/2l9cPMoA6AurALWubPzdW5BmeVfY5GoM2dyzONXX6Pk/L5/NP36UmIpKBUd
2zGEEnCLQ7/0Y9y9DK/1UUsLXxM37xMLZF0103ckttdsx8r788/ftB2fE4Wh2EUP
45kqHSyP5PwfLwmXvJEzhSjC7Z74wdVvv/74AS6zk11cdzsojz/JQafhVznp1SW0
Ed9H91ohQY0MbHPhKBT0bKfPQcqg6EMVq5/LbQ4EgKaBN3xMVlcSlP0t0D23Udjr
zV47r9tTi2Onk+VxPnv4AWeQDwiEwJoSzwaGICBLBmAl+6MOG5G+WlzXDPhWWXjM
U0gbUZPeKg62nz6v6LsxerBcdE1ECpzcMxcqCRSmkJHDzYRqkPWO56siqdLi/EUb
MjHI++epyF/ThVh4EL383M1dsGgL0ylD3HjQBxFBg7cg9TVPQOGPKqYSzI2RhwsC
nZeIy+cz/Xl4ExVuu9P3hzJm/21EJVGlVOPdvPVqqQ5P8dPg3TZUFcfst44Mrzty
GvTue9q5wWx/AglkWvkGop4BjkpYKKdEp0XtCxxRDbboAGlLQUel7k0lopMXBl2/
R+FyB7hGhFPOTg3loRDF7KgSad/xaxerIe/n7KjzvjNuqWyEoxyP3VKEC6plGFkv
gBoqHFo7Zb94A497JyrJ2WfPAO9m/qXdYkUKqYZwTEu7GA4fVLMtiRnMyWAjCReZ
mB+oyU6mhQ0AQL4BchM0A58g4mKof346nKUOKOxT75J/YefrpiZQ8bNbSpCAg1Rq
wBY7tm5w8oF8tS/Ncr1UMRbs1NkodczT9gzxVEtEpx6jYkx3ZzIjB3sryxXod+Bo
voKSD076YALSYZ6Rw6CH36sEuEqoPAbFdAqwE8guNQ6gmfMu7hANG85BKIGbXOyo
eoMPWI6qbonPs9gPz5ZRD5BJXYujYz0jxl6mLobRNOmetwd64gKUADwbqULbxL37
vCsfDWHAF+nPQGykB0/6fC28Ev3jSwvXZhQSrcgs/TzTg69XhOlbh75uEERNi480
EnN6Ing4pDDjEm7Ijzx4xMQ4EW44YiBr/FB9rzO4XTz7XzFqknBdrs0chpaEmot4
GgR1Y1IL7u1GnpzsOJ0irf5EvLNXzt+lxKQT+GMiKEEslYKFFK5o9Qv2HGX0KJC8
6RPvLAc9bHh/ZiqhFt3SZB+SJVQYkoPHW5TGU71LbfNfx+GVmAnMrLGdgsyyu6bi
/BCuI0e9v0ykKeHe6OmYSeDwniseMGDLBDrZheZ/dHxx7qkf6eB7WNZdtrYAq7g0
b7MUjFceqeqEOELxL5jX7IfabjIWj+fAt/pasK5ZU5hmr9hKpLaIdmLP12SNnq9q
ZN4sdqey51RUgKajgqgvu6Fg1NvcD4NoUu+NjTezxrM8FHniPtg8HqjclDWnDecZ
HELOfPcmKoz4x4WEyIk8t26R0TkfP06W4k+FD0iIj1QWSa0o9GGMDXIur3tvNDqq
crlqX7N9wwzxQCQlg2zdqb3iLSBloZ2ToxHGDJ3oa96YJ6rbM6VgvM+mdFTtnU3i
4XFa4ex3jcIUB5Aj2f7otkIkQ9sSS/QsUHQhN942/6q+Uf+s6ICqiuxN5RO9gUnQ
5mPB3pJD7p5iNHcmOquf7IHx8+dV4Um9P+qp2diOrFlBomu7xjZUPstm2Vdi0D4k
DctvGEdbGjQxZz/QMUfrowVckQyP2rkrfKcN3hZPpegGhbcuIXEyOUoEgVd2amtT
CTAWou1hWXmAoe1ndFm/abAs6J6Ntl0qwjlAvGp/WpPIuSa2CYiFLtbCRg5kEWI/
JXzgO9k3cvda86znoa4ZmsyzLRh1Mgk14v2icS67UlIVJK5kb+1EiudAtyC2zCWE
hDyo+7ef1FQ3T8Gt8rQL0wshMw1QAKXWxwvEFcsuU8gQ1ADJROT8ZIzSNTyEcxL3
92B/vX0lp5bLBszG77uhB5OQEMp4GYi6prqfTOvUX3SbEFEvyJj8ImZmOzby+mdi
/3CU/lTmrLai3JbXlN57xapL7NhMvTNiwalBwRk40v4sUyzBkAhR/MRqrLGBlNAE
9HQaM/1CWt6H2l8CcYMGfoe6ObpZNJZC1ayk0j/1UtqucqRGDsNPMtobY46A22vQ
AuS8hi+COJqtr+HI9Mt33m+HD+Bgcoy7PDsjlbjvYrDudKwZOW3Vmn8xBbmcshkt
PV3dRrKOE3R/XKReszg6YSQSgrYcwVYsHDVV0VtHrU29i4O+C8XnTsf8M6tMAVVb
KrxalaufpINCUjwwFtjQEd4ukJGa2+yqQpMKILOEi0S4beOrUgWkODOQwAEinWNk
pXFzHDKu35buZknbZ+p9+cnAAEjHzPR6wyxZU+/jt5nGvI/SauM31W8/2Tx2twAp
NY3tL2svc6g48GtUz/zP54vTXicDJlVVv/IxLCMxdi8LPlrWjJRBm2TePabAONDo
82TIzymVVVeY4UdgrIP/oTC7zJlKVbcCycuJj7c0fZcm6wdwXQ8u3FiC9EZyCgTo
tTLrVMciVw6eu3VfR1UjQMxJDrFHdwLk1JfdiayosECwXEiNR5YZAw0JPgVOa3QC
43vEU7t9ubGMHfKeala5GI7yH9ZBEbNpUjRvwPrq+cGHKbG4aSoZ/TTlpkqVmBwf
Vz8QqHIR3jxDV5UUOdhukMoq28t+VVxpoEGMf57ZWvT0FDOn4FLjMB9xgpO10JRZ
BsOQhkObAyaVskWNyKIyIchr4g+uuSjrIUIu+tdX2Av23ht3X5xcgXqsSfeH0+xp
4bkE9b3XM179Yzxjp1qQWBcUz0ViP+rbm88fSOBPT8QfscZrIEu5dDJMjtrHVAJg
g3mjojSzF2POZXyRb8Qh+chZB32dUE312l2k7rJMZGl4CTg6oyOJwBA6uPKeULIe
YQQ816sXwvU58z47mfgzWHFioUJ8WHiPbNi0k4jgFbdJ/jgUA6YeeApdZmtRIqSA
CMR9zsyAd664/RShZTW31WQu1srkgNfzBIVBoBK08PCTaXnV1dKC45dvm2WysYRx
g5Ldd/+Gq8yEQaRSiJQ1q8MgSuwNPw3vaPmeysV4dS7OGBFO55BmHpcK+MZ4loS6
c65V2Kh8XKaRln5OmiMzZvNCiRl1mRkxkf3BDh4KHxhx+lWCmJyNXeRfj1OI89vU
PbO7nqJUVVLv4Tpev7wIcW957ZCfiU/WWjFusb0HmjUlpKLWEHFef/pTFHwq7tFh
YlqWUBLZ30oxv0SDbSdVR238SnMcO/kVv0OF+7O0mIbnCaKbiYACU2uRuv9om5g5
ntKAzTHFJQ6VLABrBiw+T+cF3W6nUZZW/InBx0MLAPcarIsr3n9GwJGIhXH0hzbA
0cb48n2JXUEcrDuqbis/yxO8dtj0PcAL+euWkQDjRkPnaD6D7SLDo93TVIEVoac5
0oE/eeSrJDKy8d19rWOKOvZ7/0C6oo7chB3P+4WYKCUU0EKDWziDBuazWuoOG4Yv
5eXEYi7KbyUcgrlE0uwR60jWE1XbdIZabkrf5fE55BpYrRKoczh3c7TZJ1r71zUX
yxusBBEt1NqpLsFE1emx+WXRuAczLjqhk2HdSochbMivHqF2qYSFU23QPBT9z5nT
yxcVGDMUvr5i7+9aGX0tkFOzkS42QsLhTv/6DniDLwZRcWesIXhcrfArj39j4/rn
mlmQKuZL9/wOHAgEnekgG7PTD7psXQ3d/6E03Lpd5G6XIL3MK6rckvvecRFF8O+C
HHvGxKJsPdsNfT/HX0z1dG/lqt40bW0dql5IHa3cRqdbXfL5rqQi/XtuVqqatYgb
me0X4VbcMzWyeMoDFZp1R+/B2y7pl0tnU8POD6kPMSx3L83NSuf+fSZ7pH9LxxMd
9dDO3kkYVcQ4ot+AlLCb6M9NgkhVff4RprRFkp8vLCQ5iM63R0UFOEjUU7gu2oKZ
rplpCuZ/D6XdKbobdM6bPs3X6ggAKU6nwz+BTfeeY3RXJlWaaWxghVmtSMAUr0wU
Ov8mauz7odg164DQBA91VvCv42hBPWbG9uaOEC2kUkEicwEnoifDzTyyBUJynQt5
rWISDTjRTUwXuLZxojvwtmAe4Rd/atAXF054+F7Y9mSAeAHjDrBsAykTIDXFHkwi
lyz2BfKD29fqwVrUiRuXMBBX/pmT+i1qltwGwkoR/zF1STX1O14WvpD5RDle+QXz
gR4viG2/S5Q11pzWugstKO9h10QGlCjpec+TB1bPzUqpE7BAalMCIdKzCITM3v6+
wgdfeYoobDpOUS7VTm39BjUYULC9xbWvDBpuREyh/AwP0kPcanuwh1Z3L1crDqyS
3JsOd7CRmvzOjsj5qVptG9RrhdMSH0iCnSkg+s2lsh3qinNeoruCcrdBuTDstPzH
38EdYVM4QdO2itOG+JSIfPet/RfwGjNpHTsd74011T9BpdAfVWAfor1Ua7ptvpp8
3wDyjglsXLhy1G/WP29JB+MKlc/QyCw8GE02/CwjNsBf+1rzWMJDiyriv5gFpjTA
cEMgeNd4SF70PZD5+21pBFbr5PDHCJJYIATERYJoFeG+S4nP/6XW+Oi5YyUhkH4D
EvmWVb1rmKw/Nfa1+0ab2583Xnsi6pSWw2WpmfHYirW4THV4TVrwjWEZAVSFrHyR
VW1Ei7kC8X80fGUX1mNNfFUbulgBRQnSe+VVp3ynqxX7zokp+0kFEnGB3wQuMrh1
RnkgRGQr/we9vpuF2mQJy5BqzweBXXHqURGXPaJiV8r0y2P0Pt0tPXfaus/Kg6Z8
iN+iuIyKK2VTur/zOSbXEvSm52dNc1yhAd92X95d+9URJdIjLuV4ZfzviklOGWSF
6+I+1u5zmUHIamSb5ZOV7XAaw6QvY6f63cMyMkjb+oHSYaOkbgVjAo0o09gtHx+S
eCN00GEqn6/xU3ZVKUBENziFP4adoAUq2DWOgiQJJQZf4Lf0w0ATjKsXBc7G0rum
DwmhisQTM8tULsDWz9IbA1H23AkVaC45dOPND6VlEOhq+NAXK30TjFqtJky8iPC5
uZLm4f7bI420rrSsrJgx1ey2saNcGLC7TL6YOs0+EcFoCw/UVkxTquhu7fz+c1G0
WIOKr08O4slh9caiAFtGyx+OkzeLf6qXghKJ6MVGfXWgts3q5Zv8tk8NLMiZfx6d
jcbvRaTxeK+JvDFpAHy081NByYTjgkxTPUnuj4qrHo81K3HDyn7+kh0wQoUuCtrP
h+XIKs7WVWPP/aGnYtOdRnGn3BaVckySHqIHhfLPRxrlh3Yljsy145ojcGNTN1L5
l74qOJARtyiGprSkSXUZOZWTebhke7qun8VzB9J6SWAc9/z7YrFL117BeASjbs5a
jnZ8Ee1BOd5p3IIbP4bGd0x+6Xe5AdCSkzbL4QvVGamtc4iOjNgvGGoUGXS/czMk
yBvzJz9r0DFxsgk+TzoDY4JXWiaQj+H652WhX3nxeDP5slxDOHJ9Z0e4NcF7Gv0r
8z7wvPwVOKO9YdDwEb758oL+/DWIhOP4nx/LZ1AblT0oGaaTCPe/6FQhXY+V+bYm
WP/1u5l0VbVWIcGRFJYnnzausbh+VrFtcfHgyZINhZVkD+z55nNCt3Fn/T+DQLYn
vyxyYu3oDzs6Tw+8dO+Dd19ZMD7a384lwWoB0qgrBIyXyaFVyQhj0sDamYbunOfn
G8GIOMrp/R3orjP9x6gTPvy9r778VACJEoP1NBHkd2A0PwK+XHDdZHFZa1SiEd5F
N2ikLc+3r12ZQPxXIIbXrcCoWWJvI0g9EjJ4z1Xdh9im3SkjUXUdtWH/fXZMMW34
/6ZsDYWqpJ3vhqWjENvt7nJ90PPlDPeE4DJUGro3/TkpP/JA/rDX1d+0qaV98jMv
xj7aUV0m8hpbQDy5n2BcXkGHYQkqO18siQsWFeJLa6BNn7/+zzt6dcL8w3m3EXPW
iloR0XxAjcN700Y3KNDhlDqbGI//Cv1ZK4uCGGUnEoCC1F/mOoOcJHjHDULrUWvx
3rlzY56QpGE+hxybUPTzC4a0VPbP2iGe3TkdEO0DqAs5aLUpgPyG5SxqxFj7VUGt
Y2SMnlL3YpwjwBT6bJflv59IEdkEeXtGagsMnQAl4iRK0nSc8wr7U5hiArG3xUdE
8VPrdM28i2Bw9v2ZmgUGjrdR+Dg8N7EqE8SfM7FI/lsblThaXgBmm7ImpoZk0hgH
0PB/yuDIJoTtgMXi8cylmgYUC04990H1MlTyFs5Cu1tml4FsE3KMoY9km63qp8+n
uEalBQmSboTXaZUSlsceHghtauKxzc53n6LqaT+a0SQv9g/BmWshJ9W51NTn7/lY
nsWnBWfY+ScjOv13F+2Wmq05CjDDclgys3ZA3ozyz/gdL3H8XayEs4dh3cmuVKMi
fqHDAno+CIwLfJ80QoxMiuYTqv+OznmTDuRUiG+fEgiqe/vKY/4365SJ10q1KxNQ
wdIzRmjYAdyIpPMXo4eCQBMpTEU7MDSIFsfNR3kFdB0WLn6h+p/mdvmnDXiJsuMN
tNUiXAGccOq7gAhiXP0/8muqKf1o9ISADDkiGq002gtdb5pU4pswqUIJj1ShKd+7
VAGsFFCxDSfQBIQGIWeai9l7KL7K1G5h/w2ZBYy23qINhDzbOCG51ulyjP8BvteT
vRuWgMB7ZgIwZgrZttBKjHJS4kJbv0vqDHWYsyClm007NfBBPFOj5TmGa//S78Nw
RxC8sgbz8wIjJu0QexDpzKfIza/fPtUWx3HE9Yq2Mszvz0BhzpzDU0bmXej0k4fQ
12bnRzi/ABsMf47XMD1Z+qMdVVQtafCq08Xh/0nU7hvrih+TRuabExSAphBsIRYx
5aMshI6VAsYA+/HYWi1cNdhhHoveM4LBBYA2M1KOwfhiOo6bw76GYpsdOO8DCPKH
8lQHgTYp/+XhPcaxg2AlPhulRF7FN89tUpT3//FOj0pX5bSyrrKOuckLFZShBdmU
IKw/oW+/Q1vrHlSTHaGDplaoHolFWIuYNQcl84khi9/AbSVfWNKd7kXfrVCrfkd1
kLKasnHvz60TjV4/uEV7Pc2CkPXOAVprMr63IfccTG9aSndox6u9OhwRvEfTTJ4n
f59NC5JelwqT1v8EY4QB5icVSxB+V3h/2prqUbzseUv6IzjKvVoJ4ODLr26nY48R
SnjnkzNJQSBrdn7KhkBj+n5VrR+PbayvZUYaPimsUqst9qFld2Rh2f96w/5cWj0u
L5TITZCExTYPWQQm4VXtlUk+JVRtxdQxqTWlV34T/FlW2KcFxvinVT+VUwLWxbuK
dPAezjaqT16wVZxY3/nqL5eA8hu6dqlwEUUbGyRWByg0r3x4Z84AloYxLuo6pHhj
29ZWrwQZ2DUj4BnBPWU9d30V5WI0f4d5PqEjkInV0jAl4NfE0rsz377cZQdutA4t
u9a14yB+fMbamA8gJgWybd0Cc7+KGb7ipXMnRmaJXQO8sAV0hberEGbOqG5GuAZm
V65bLJZmYK66gKArboGtOw==
`protect END_PROTECTED
