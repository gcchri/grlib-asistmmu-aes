`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qs0OFToyBDshcmw2Pkxyf1PZQyV+KO6EALtFNKOwmqPlHhWuDmF2IAwjkj30nj/A
wtX79oLM8e73XZaFH44v9R0wBEip+Ot6YNQRdhPNV6CWYbq0hJy6EiM8ZQo2crsz
vjge2rG1NvvCwngq6opo/NPGzS0Sa8f3yEpNTI+iZNXJJdZGIoAD0S/+uQQBqHT0
ED4DYJnUN8ovy8T6qB2NrSCK4EETqBLkUpSy4ww52lIwSREAdEZgZZhPIdqq9HF7
nGVn+S/eQr1tuTIRLPRGlL82VLNHjOW1o34QyKtSAW8Qnh6ZMPZ9HSSeoc4rHkfD
6LgHlWy7uN38mJjHi183qbhGUFPxK9RuokOfP1vr1LAUisJG6xLUS3P68rJnM12k
+alkQ+UPwqvuFYk9XcTGgkMIIm4T87enW6r3L8NlzHT3MjXp1yV2IeaHeJHk9CpK
YhVAyi8ecHfGHfTrLGgKinfjMiTbS/t6uFBeA+iy/QP8+HQ+UTOM0l/Qf+KS/A/7
EZPMTVLXiA/Wq7n4x26lQPvI/mYc6iHBfLJEitutLL7Z/M5sy43OuMcYGooPB3Tb
oHySqhgFy7H2/Z7IR1iIGvX5PDG8kmmBeaEMnxipSW5q9SST65D5lee05VVoF2Xl
oDS++yP4P4a56S7WiwQi5vw8RXIhxMAzxcxjmEL/0Zq+S9/sNHeGr06uxv7ZKlLv
6Y5FkVD1dHXrGYYaT7KdNBbgechmdjSAVXmqqS5LA86znHmjDNnLcI6hI9TqgUOo
nDdmCG6pLGWbwRGmz7WTLbI5nVKo9D1+ZsVQcIGqDcHrvNc4OkEPxELFEetZspW8
5zoIDcSts+06KJp+YoNPKn85yQypeR2ZHy5CUbsXgvISWAdc6vaPCUkzGmwHZRQq
cGwBBPovUGvGWUmK6rb6oKw5dwkAPHFmKprbZAGBBpCMXPi9dU1OK7UUJF+UbTXK
MUJLXi0MN/XpqT6wfU6bV8zie/0Fo3aIj6ducR+bLhlbSKqmTXlAogVV3DPfbX2Z
6i09anwff/iq4WYF/MfTcGxR5xPSu1E2ogERHn2d0GHxM043rpDcovvC+8wGymAf
vN0/e9KaE0raZAXSD6RA1sytHsYFSy1uwCUXc4Vbao7SmMQNUDhIFt06/Yi6p0S6
ENBK2iP6Hj1CWQvIS4kt4rkqjOqWgNW4uK5VuTkglAhn6rwudP8YVBVkjwph153z
wlQZeGQQaC8xBI2svEkIBq4Umzus4ZFLr0caqi7Dx+mb9w9GGXmT7Koa+SuOZdBw
qnM7cXQ+aptpD5nOaiHK1BFqwc43Zsj+6/0CamA9ZHczCnHIh0rQHY8lQmYOhcYB
aGqF9CPrcd6owK8WmD2HNxeP40sXJeDo0NWbmGB78/U+lm6yYVdGMqDPfNePDs4u
ItICkMzc1UTDmob4DdiLFWzEbFZqhvsIIyQKlRXYgMrywVps5UIUyq+7fto/WZsZ
MM0t2mvvAX28FH9JS++Wl8f3BtDbgbzYZXa/jlmGMTTQ+G3URyrk7fVWGdNtwaGL
5Kh054Hn5Syg1dJ9/WHVpR7o10kpI+NijqwY29JplFIHNnJeoSNx/+GCEq7sIXLZ
0EactAcsKdgV9rHn5MnVgUn/S52rGGlc4D18y2xnxWRNWgEsWPfMB3g7ThIZRlNJ
yRir22RwF+m5/RNI5FB3cABUbCiooWOzsyfKK6ZfqX/BwWtJDhOnpqv6fXroGzLz
4IhRMMBivcPbi/7Oicu/DT9Md+liBGoKnKoIfegdvi9AaYQijFQWAsh7vQGwDmC7
zWyEISJptmmfxpL8tk2f66kLbrp6wJlR3stDVDkDwARWoc6FpIHhrXL+ex3upEsc
X//l5X9xT+cjMuMUtZ01SF9aAauoovsQc+SLVAslIRqBQnKZGu8WNkleHXdfft/l
`protect END_PROTECTED
