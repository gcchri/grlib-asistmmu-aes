`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i4eDMooZKNItKlnVU6VciffBQZlxbWIix3thzIj6DMy11S+zuxIblbYS7rwRHWeU
qCnU7wS/U0Q/L35gYPUHIsxusJbf5DshIgNa909FIL/7cO0jj2FVIeIpzW7qE5f3
RGxSck5Ie4QmNQ6kHEnD0GWSMxQcpOM7KDmCNAB7yfbxW3wqiLcqLwJMNCw/4yFX
FEl46YyVS29xdeISSExtB5/LvkLdXpaqB9y8wSEJUj6IxYIkrIlHS93qrFFSinxG
UWYcMAkeSytOiJiPVuLyyHVIOOXDaGpxavxWq1ElmhI9KvTYGYaXOWK4WMPa1DQ1
`protect END_PROTECTED
