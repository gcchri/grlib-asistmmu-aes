`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vHAHnmrKTbGfni/Wbx/ydnLfhrY2PNOqZtC+6nPtUngiGFCiRTcwpCMbhlEtICbW
oGULpZf6981QLgqtTNHWtM8IguSVq/41VsIHd+WJCyEvtZdq268/IEn/WIFqkzn/
gpGp6okwAgdwrgTBpVOFwnsTaRqD0R3SzExhrYF9KWdhEWawjs9DoiVcQnh5DWHS
C9omhhMMbxkZpj8moLp0gCuNdRip8PGI5JL+OJWVNmvm//luRaP+FPLzY4jU+ofU
wIPcPqxitVKTWdaXOpHQkQUUd8eSceuMkgdX1vQOfyKW88mmqrlV5kNOk6SF4jy0
iyVyEITp4ZHFfqxVVWV5t9UYslWxD6VoRoc5r/Lr9QM=
`protect END_PROTECTED
