`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8+YC/GqFlQ0rq3LXkjpyB+KaZ+EkRA3WTM6xNUJaMHwrA9AAbEBECKW2boTmxU1e
BAnWx5vkUHgvuyhNc4cOwQchCKVAfYVdlg0tI2qp7nPevOAm5qKHvy2xDd3mYU08
Gdz1YE+5q0w5ap1u2CmhAeu5nEBPkrFUoi81Zzm5sRs1/maAfzNdl1lJtaMDgpnu
YoRasDXYuSXIUBMrR8yuHPi+VHkv1wlS+zUmaz9VLAHf3pW6hgxuTQA7LZJhKapL
L6WcB3rNmR1Fq2sMTxYQpP04XQmfNHNHxR/E5la3dONOcoronEU9ov4Ryo+6PGSk
wWKhIlXE6p6raoKXOxCvWA==
`protect END_PROTECTED
