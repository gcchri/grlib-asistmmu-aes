`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VYb+wJtgVvBI8FnfkzDu4OfFo07t9ID724aI/aIdjDoFYcZVy4RtLYfGgKYw3JbY
gOfGjPZrWSF+XjGQ10puSToUnouOTtxLMHZZV5IuVcXmja7jWHx8llpUnDxAOcjv
ZYaDgfzy+NATREq6e5Ymmviy6Z+qIU5vW/tA1mEteCch99XXjJuN03Z2lTvXJU+Z
UElcLMXuj6NUo/rhxjAPRs4eN5fFpNcBjERT2ewxTFM8n951j/UyjUtRAg9q1bS3
1h5B1IVcooWitmiI2EN1eGoloBsPYVkI3LzmUCAQ8ufTFATomCxLhhAr6FpQk1JZ
WvA+rtkVLO1jb2VXs+fPo0PSBKaR0XQmiT8FZ4xsngI+VBn9gjfS+a5WQoAzI9iD
S44LeCsPwU1lN/z4z3RhrKchNvGvrqYqsfOUnMz2TVPit8DOibBHFuWNfZAN5soD
/AXmccHBAgI40j8YYWJTLfJ9j23s4xM7FhEFpFgSsaxcLpbtU/hhHPJbCPeC38A1
aRfDNIrnEe+I5KhWOB6FuGbciOBmXB6UqFb25rzArp/WksaN2VD0fYDBPnViqWn3
WCkVKfzUJpxJgkiowsqSP5YClAzQn3B1bZMkd41tf1/H3io2xuXbsfvro6p1YPJs
n4HU3XBDvrGI8X2LbopbQxc146NnoOIpU+KIvWD7gtVbV08W4jJ8/DTpZE92saHl
nXYpo48FunKAe9OatsSqOqw9cytiDlqtQd77HEnq539JDvA8/5Vnn9j23cT88urA
MJPQASltHPko4IjV6H4RCElskMCrTqIx5ZDnNVg2/C2f72vmYsk9VzZWVhUiTu3C
PKgQ1x509pgGbogn2PbHMvDurkt8iJZ0JQ/dnJ2VutX3t4b0y8yd+zSYCV77FREq
/SCm//t3CftF6dkgng/4b4fKHyiTdbJFxdHZyhoVxVcRlm8Wf5t/OaSLl2q0Tks8
AKWZUYelRBwnXEegiRBv9w==
`protect END_PROTECTED
