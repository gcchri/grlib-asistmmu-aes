`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hL262MQF1SMarVTklkQDCp6+MMKeRmAvg7w1x6pAKuWj1SF+FDQxiqpCHghbbhbG
vLEEKZ0wjdKAl9dkbDhnP55cHRgPt1hFqsgzlbDitKcKwpUfMiYU3VFDisQau2Ce
HDJiU787EQhC1rfKn0ZwHXyMFmjMOiqekQESvUTGHRRvUeSL95ZT2niL+vHl6pJo
Teq4m8QBHE5wTUTfTjAS9JT/RNducvyI5QVuNs6inW19o+BRXzQeaM+YyUXL116n
Nzs0aJJZRqfjvi4TrxTzNOexwUUvTQ7mHXZr84qW/Yr8CWAic1SHJN2JMNS5T6rS
gd0Z+9wzNw6XgjuVzurSzZjXtAMFBBU5yVQUNvlf1gyeASiUMKKp8cdhhWjjM0Zd
svzRvK6Me/a0pxmUA0GoRJi83UFDrhYOgP+SbXWoVxswn9hcgl05e5yd09Y6ATmM
1j8V/tMAOsA59zlZYRGgKKGJkzwlHnCDqojFbDzvh9hCPE73tPUHbwhf21A0Q41O
j9l9i3RqotdcInYg7SjJAJmbcdspK60NehjISL3J+IpsiVBE01jr2J7k9NpqV+1A
bu382sBTqv+XcXAnEa4eDDMXMYWH7/2MltP6b57a8gZA7jEFcsqjQBG7BxvWrNRT
EXM7UAp+5hoI05eYBsf67x1K/55Z0BrVqzile/x8nPt0UT/GH1g5i1RtNGycfUKn
ROd/zjR/5L8BRWedW2auSpQscjdypvH5ChNIEA5EtGlP9+bmje1XNUdgE3FguFfF
NP8r9qx+3K3fNGYNrZl4uKsDgHz6LxM/TtiSUK1pAiKdW0Z06SqJRxysK0pT4H7G
gj5JpRuu47wYlZO7hrWhhdjBs2n9/uC14YdTUTwZNvFTXx/Vkfw7WLkaM7A3xTcj
FE28a/zFuem0Idscn1H4iX14utmBZzCWtxtSKu3KVJhdGo7UaGwj9Uuhd5ENd56d
hUfMzQL443CDAgMhCUmwhA==
`protect END_PROTECTED
