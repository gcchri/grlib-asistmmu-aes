`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tNAEubMVPKsyXmJu5x+5x/9L4c4K+kr6fPuEdiQ8JDhQsoeREBxqrsm6egDnvxR4
ffFSQI07dM58I+VSbvns4Su2OxAX0xClZ6qf6JesAko9a021rUOAnvO/IaYDUv1A
e//Llb42u9WG0HoNRBuaKhUpNF2s9lcN23jDV5Uhc/b1znf3CboDHAoOmOu4zowQ
PSNnDNeDaODeGxoKgP8TLVKueW0GzLyss8u/J+CDjm9PkZPEg8qh/aFYcdgzGsdS
T6v5jz+FwqgyFB/QLe7xR+rGuozmZ95KsoQcMhUSwauBUihFrkH1Rgcr+/tIe4UT
5sEYEYjiXG8OyClydJJggIGYOcY6fDUXdVvaHMea0x0B6VpTIOwekHJCAgqq5P6n
kEC5foe8I40l8m7+AncMY8sPhuyo+UsP5JTzV4UtEUpWe9YYsBW5Ej8IBzsQz8VI
6svv/TprlT0cXgVNxWeTVX+AJD6rn41QFJ1C/C+hpc7qzMLEkQPEIVlSTgU6XzGC
ph+sNszLMYbHEvsLic4PYqkDr08Fuk84HGopQF+I78F1joYs1OElo0LIv+dYkzXn
AzgfLOpjrg0rApgtYZuzbCz2NWO7THS3GocPltj+ys8=
`protect END_PROTECTED
