`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IOoHLGPr+aWoTwK8/KCZkXz+JRsmUfVCqcDCYitTDL4/ZCjAX2fvX7fNRrNGs6Ms
camRW0p/dZJ5KJU0v/aGTEhwyiP4x2qrrMOfS0kxpX0WR6C7q+0BpH1hmtZ8VnwE
B3mA+1kdxExvXuhxCqB52R5FtZWiLcTxFEZk5mEoZFi6WZ15as9/RHHnLCVDREi5
WFtHhERk9sRDHqbwajODEZP1p+sAvFI6S3IC/nxi+84A6ispvExXLFS0sqo3cF9x
ezDjOli3njB+et8x9TYeFVK47TparBeOZRaWn+yIfMFQYgim0VFaU09xNuAlrLwm
TuyPwzrw8BZ3iddhJ55/qb9+1QNe22DOqZkRvYEtQle8kS6n5P1BkVbTs6x/Oq0J
FNfNABTr4Mi7FxXBGFE+QtsKkRswAUElouPnIXIQTkPmbTT/RirQXlXQbFU8wgal
lbiysTneX32ougQJQ2hHvg1LWBRXr+b7izR2cNva0jU=
`protect END_PROTECTED
