`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SPY5OKF+GU0Eqmsz63VCYfJ3e+mB+WA+zfQ7yuUeUd/vB7IwCk+SMmW5fuf9T6wN
+3g98dmtb2pfoVB3L3rk4FgQW7MeOKbsNfP7Ngizh6gOWNkwk/Pj86U4O/cHRxeT
zCe8msJNUl3XHx3J2c2FWZMPovN6resTPmMRAEsm17jYifoRaLiJEzhbc+ATjeYK
0KaH0W/CDYQ6yHZdZyEyqLzs/YkZx+EXOBjnLf3684CeGMZJCv6hmBcIj0TqKQiR
EuKhJ/v6gcwk1M0YD0vmHT8o46yFpAMemDpX2LRbHgeJQ2JeLWiosVJ2vlG14aDg
O6F9cSCojQg1/hLzb8HuTA==
`protect END_PROTECTED
