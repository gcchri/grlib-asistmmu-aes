`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4v3ayW8FiZjza9DNva+NmfeLeBfJSSX6L2uLgijsWH2GJKHeocRrsOjjZXAPI8ys
z31JzoKaybU4pfWJ2uR4Kt8TSOWFyQZBPAAqniPUNdhbMOTYYsDylCLfjsp4Hu/7
KaCO5M+tBzsr6tU0Xl8+zn2rqtshiHe7Bv9njCQvXOFaquOUvnBYP/Zbcso8Yrdv
1HOJHA9DBxQ51rbLqI1y4qX8NPH+BBlUIM9NnqjVrTis3fqf5Ip+3H/cuJEGHYpt
4T0MVZXal0+/FVvV6+aroh1rYGUgVFV5KpsLimm9BEFzEgJKBV0ybU93eb95CYGD
Q5U8lnL/TvVHvopd2yMw+DBjxu0AcVl3U724c9vTLKETxoyYFMXDaf3PuA1FHMEG
mCJRywapHkJO6kcVfEYchl1+QmwGdfdFsWv3ZUvYIfjiScslw7HXeIAF1hbOs1RB
`protect END_PROTECTED
