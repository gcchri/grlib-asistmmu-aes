`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VbSLOtQKS3tmpGnoFQ70dMIHAHyhMXWwtwF9aCjQ9+Z6kqQRemRQdgFgscxvtBPX
6KUPQ8bhSSR325/uNNWOGqqMaoLXv+lv3Bp2JPyg/whDcqk2bd4mwnIenFsQkJC1
50i3KTW2CBHjEZW5sXdRCRE+CL2PoOiZC1dvOSyUga9YgRHdC21jkHtxlzCgCnwR
5Pa6stxeKD7B1eo5ncjdntfAVyvvTPsgrH7PM61ylEVGPWwzDNY5pfBi9MRMPS+V
CB/Bfx76EGHeB60hQ84FxZhDHUuJumVaUj/U6EfkQsiU1517l+CK7XBGFyCBbsMh
JEragfEhLx6Id6N8tL0jVTO995CRK6EYQDA5CfV1zY00vanwJ4KYsdi9pI615xy+
OtkXgEEMMoGx+5cIxxnd1csCt4vofyBhGxfm/ZC3ABUR08qSJVXe04IpDUtICWt2
0Nf0aYR0l3findclJ9aahZEghSSVkHrLvkHFBC6j2cHIBQxKd+I0ZULhPr3VgoR5
cvzJaBxPwfCyA4oflP/eYJbS2Egv4BHTbYE1esfCNapNfsoUYml93MjdW5cFPKUa
WQDJ5zq4xeRaEXps2e0G77tsyYlVgD1A/GPJw9thB0jyp3CNRGXOgU5VGo8g6OHM
7zgS4QZFinF2dSLDQ9OkxbfkI2gFucK1mG+nkZAe5dccWWRPbpCaKWwG8bcMoyhO
+m4FzOzY9WxentgdAJC2u4EcIJa5R9tQ1WeedQz9B4KyxFkhA34kJdIAaBQkK2bP
1VFiHBxODa1Td4AP6iu1E4fZLJFmaLT5MsXd4Td4fMeiMWyaZVc12d+zViOG3c3X
`protect END_PROTECTED
