`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h5MZBKYUFgSIQXCgrWV2PfePzwvkviNhj+SHhOsRNN8oAfH/KBYQq2NcNN6OCAyj
vd4c9zjj3w7HlKStlSjzGzTrBQ5gM/6BybJidgeAi3nTjo1HxNCDXkDA5QSaW/KR
0ca/1YbkQk/QIqNekgSDYeKK3O1vXjYXCwyONQAFCZLhQXRR1D9pH77sg80rn60K
gztEINPBhLv7td4PZqv1//Na0CpD/SBt3yMZmEe0hmqf4zjDQcQFcRicAo8UB6pD
I7de40sJsRWvbaGqWbx7Q39V5TjJNEQHlzsC90YDlC9iYGAsGtWSXBEnZy7bjOcI
ClyahibpGFX8GvG+AFpTo77Mr6mUckafqVNcX8H7IcuSuaoo+5lIFsloLBc7WG8t
MfVmNfrTFF/6W3/Z56OzenHUW7HXgQKA1+sruSZk1a03yxJxFTq6TyavAlnQFV1L
R2yQaNi0+djLZNOQh3M/ocSZXMU+BMJEUYmGlgQ/dyPyDMzX+8MG9afPxO6/Zb7D
xTZq1seW7mBKCXP8xRu0kRTu10QKEyf83LBom3bqCCnbs/Nxxzv/vs2/dDeSA+jM
gfIOG9CFZo/4Kt5FDc0DEP2ff9cY53TihLaf9EwuesouRFvF7BoNi9hRItJM1Aq4
EpZrrc6HTm0JxeWNnIMfkw==
`protect END_PROTECTED
