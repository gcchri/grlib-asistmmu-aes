`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mNSxFg6TnJgDT/dlXYq2dLq0Ml4JZ2W9vK60Cxrl1tlPA3sZSeCYTDcoBLTKzLfV
IGEGmOBsYyzq96g7QE+hvgKPx6OuWYvnoaOTrv1mAJ7FPFOkDTiRBDtbTRzpcDs5
jrZvxvCPvhR16EX5m9PFE4s1ta0u2rJYZgZkhnNLBYAfxDnHcXbeCtTAI3vvceA1
Nv/C2CNPdn5O6FOGc6bEvMJDk0K18pgTubIvvkksL5jDaScPjh9e3vo9CnV3eaJc
7xNNQbjEXjduqp/aM91sS4AOXv3/IhF3O00WrTDpeiFA39mD+pHlQ8qoPez8gRcS
F/kpaELH4OaR6Wv52kuc4sN97ZFHeSOjOGOcWA25yfT9q14vtDNldRjCb69APTqL
VyQ7r0Rpzt99pBjeqVZyb1FIjViiGORds6IrxC31TF9G1uxE0TvzrzcVzVeElIli
eq+Hda+/wJbcYdlB4nPPpY6Renyjtbngl60VaczqxYCC1txgOhurzJ05Q04LPv/w
C5yJhMRTntVLFUmBz9YQOzg5O1XloXzU+HcYQ8Fb/9ArKTT07jGlt/ZQSQ4iQmhM
k1hHY1YjIWHyQ3NhOHryC4WbEZzpek7ve3MkdSauztIGLweKP5FampEuS9blqmy8
LGKe7fZXoGg/TWC4f3beVSZZNVYzL2lE4sEOxLNT9EczO3SA63iR/AhZiedJ35Ly
`protect END_PROTECTED
