`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0bzeKb3XvE9pV2rdCJhVZyxXWuJVAsZdoR+GANPca2PbiHAC2mZp2wcYJ5ixNMig
/bb/X0lCiSi/NeEV4P25WPt8APp15sECs8UvI5HYfW5wwtEDD6dCQoCg42uAfpT3
6vFQUv3/DK9Nv+187hq11Hq+TOd8pEUn9k+SUj92doRAsvFXXo4Hh3MAOFvSMjWm
w3V/dk1PfOQcmsNXOE6U9pAJtX0lB6WYDHpMZH7q7WkOopT9xYQz1RUsioZYTLfU
I7+WDhCAYFwiUOkW+HiUtYv87nYy4ugx7aZm2JG97pWLZN3q+u6AT+/LD8GxloD1
RWHnU5yOVIXB97iiSpOKSUAEOEJsUXn2gAR4e3KOIuiGVVtZ1ElCBJ9I4Ih27QXE
UjH7XIOH9zhTR35NyDJ/gS+Iz4tIapMSyESd5xipwFdpZ+gviKYt38Q2fdtUkD5n
oa4fXKj+znzsckKhl6vZbr+zDRZ8smPQlbEhs/Fqq9JhDFiGgVM0XJexaw/ZHWYX
CwirOW8aCJ5x8jpxWDOTNub+70o17bqPHc8M4uidBmWBS/qTohrUIflMQHl2qZDA
/Q34r2iXVoKikch6fCElRytuxW5tVnQadO/j3ftKu1EX4iENNkt+acLNYwQ3Gkwt
efxTd5Gcs6wklbhZ9zD1XmMEgzRX+lYD0h/p5AxbSkRy152lQEit0qKRcGuLR47e
M7RnrHieO7HF15mbHcdBG6C3q5cozxUq1qHmMXg5Q/b7wD8UUpkcgE9Udz1BIrRn
yT4mvNjOp2ELghCkAh2k+ZeKkp2Wrd/F5faCJ2YrYf9gycdeaiD1PwvzXg53Hbz4
Bfd6TsFxp5Y20ThvgY0WEHfpEvvWpO8ahRL/mN/dxChJhX/+wlBUzjgChyTxzIng
ljTtTPVleTguV1ICkb3jMju/aXINSxu2KxUAckbxk+g=
`protect END_PROTECTED
