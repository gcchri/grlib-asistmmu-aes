`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xqoSFvjSZxBImAism3Fu2tNNAMIyGse1aYLxsMrqAWbO3cewW+xRVaFqUSlojP9p
/51FcB+wD2RlwvGFoyB8gM6c0UrWfJJ4UDKVz+i+xbeC4njKF9u9RMoqBtrJIXbH
5zKPgPwjsKQruWANK0jrFAulGNnsOKqiTPxwzc8aELdl4VxXjCdiv5e6gX6CleVV
K9vZrB87VuOenCMXmBR6oEpzNW2aAHUT8QT7689iAyP6YETnReb+jQ03fyIwn61P
4eX5cOJTU4FPlpGg1VwfwA==
`protect END_PROTECTED
