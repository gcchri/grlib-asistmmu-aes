`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4aFTzxE4aEDsSza0HjlXfsAMxlORBEZ39YcfSjj0z2viIAZSEr0cMEbcmWZ7sLHI
j0DcDnTCDiOOfksnpa6w4P4+W0tZk58vybyKRw4GDKRUXMGdTMTL9HpUGNVNRQtm
u/eUEIYaetYjoF4L5llPgSqft1+OfnEVXvmKyA2GfHhX1dyscWQ+ZGvJzcbXqIm7
Pttz01DF7whwTxO/SMZFiwzW16zZBc0FTDsVM6V8plnAe8PEJ988oRcje4SjQj4N
WAIYFvR8RX4zqMGuVnlxT043OkuTXd3vdKEe2+x+VMzd873mkzbqcOkEtydp7x04
WZAAdoFbtNuqDwHaZ+hORXJT7BDQShR5M5e5ic6jNnkX1WeP6ajTuzVpWOpiy0Ek
8wwLloSbxMihNSWYildhGbJtkX03CDpdr1sm4OkmY8o7Xc1bEQcNlhNTKTqv7ZBl
aplbs79+24D3cmccGHGmHe2j3u/yL4cEdaMRe47tmE+cbgTdvOjfYyszthcyvaWu
`protect END_PROTECTED
