`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gGzKE4L5PBd4wZavdyNHcX+wBxLII/cEdsqXedbE2H/p8F690yJHIasBQhZON7ii
QZi8qiHihV5wLJgRUy+gn4cmV8lYrIW7vC/QcW4JDP72v6R9p3q1lGmV33XAiWSR
6Q9CtwH8Dql8qmVodCO6x+VKkri/6eruq6aoipK6aFrfGy0pS7aKxLgf3ZpsP4Fa
lxZ1GYKfpFjeO0jgb4vGpPAn7KaEcIOHcVmlR2o/q8icURBnGdUhgBAgg96iAS3c
C8xc4vJPfmA43x+Os0RTXBartf6VWxa4+YA2XMD8ZQmIXWM9+ZMOa4qX/T0dfOQf
57AZlr0BHEy00hGhRegHuu3EbB3xgyeJqV7UxHv14W2JDxI3D4Ujy7sQ2KeuKKeE
o+WS0WwrsRI7DsQLuVjV0psHL50BEJ2Vxpsas0wjzPJHw4d2oL/RzqiPpeSKn2mv
96tOhCrninpwWtzvpbBq1cM8X2aYXy29M9dK2TLaYXDIr4CyL8qWtXa1BDRjzwhF
i3LEtK3dM0Az9cGUO3gqWI8OczTlJaRc0vo1WCH5kgtR0yGNx7g9OUt9QiXBYIfz
Zw5Qp/ShLUyEP5Yv25ftGZzlgm00UTvpDd6I9XUWdHAlzZBW1e1Oy+EcojWXU0aq
qjuMSCwyTSKZJzXZIVfiq6DYMiU0GI8BafjP5ccNb1DnuHoSLqishdu4NMfVLAKI
kWGfLhLv1X+6lZtGTGRsCXTjkYvlqDrsm7hC4ymEnphwQ/mneMx3z0PQvXnLWNrN
ZAssdzJWpyDpowv1kUY9Ax1u7HDR7QTmMGCqN5UcO/5Z7R22aly7874ToG4VkMja
qu/1oSruOSWLXyKjS/PbGgXpdomPLtu3YMeFE3J324SnZGZAu4Lodi51C+ZlmueZ
`protect END_PROTECTED
