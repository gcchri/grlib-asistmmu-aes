`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yWfsVyOF+VU87M1xHymYzeoTo0siAmqIGG5SqqMtGKxBIJVb5XhyXm4/RrgrJEh1
jgOMiY8EyjABvHihFDTKLnR5eGS/AGUo3+ZVuRSPndOAj/P6kk3czMGhzXGBRqLc
Cd6mjF+UoNK5vTGM+jPqrX1k2qIVNauA0gGFH2AmCKdxq8FKxkKYRxVzVJIV74og
gwqyjIoUrRAtDw7CugmnR0B4uzhbFkxiWWUdIaLVAmCEqtof5W643NXQoipC3Uk1
4g/IcjtgPhRhNbhSN4uarAieaShxpDbXG9ugaRydT5sBxKZYe9uyPu5JFySkwhco
KkaiAJ6UOKCJaxBn3mICa3EkcvbCXdGLq7a/jz+ep1YRKGYbPruyQFegRS8k0poT
Eesw4JAP1adHWczLZEt+fXdoFuG1S8I7hh8yAoWTH5xrCM1+OheSNDEXwBOP35le
`protect END_PROTECTED
