`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b4m2xmTJhLOIP/k4JKJasfSkE7VFB2hqadoWoItwrLkams1m2lrQHDH8MTGWoAwp
gav2HKpduBm0OO3p8ADxWCZWTMRuwWQIxmDlret6TtyTeDekqvCpwkuYOFZC8DVW
4QkIyliHc6DSSDaTbsBcLvwy+MHra2YWu4Ou7NXEDv1O/FTjqgyaygCqUn0JRkam
/skycbUqrH26Kr1OVV5NWTwZQt7hhXVY9m5NKYu/PTedw2609XIpzyq+qPFRDlN8
bLLmPKGHLVoT+At9T0EjdkewdYJ2wRSFpjD3la1LEnPcQrD6byNJIaOArOw0eCBP
ap/VVu/cNdykD+E7sQL9J9BynYTLPC82bnr4Qznb/jjFQOWGOSCWnC1GattVPu+s
LDVHF5nR9qAEdkB+U5A6uAm1UnrulhPomWmitwvokfhH/M18SetBwnaibxLFtqLn
ZJMbzoph2cq1NBmhwU4Jx2SgJDgs755e4H0q2VLbwoxz2qoBaDq908ybgf/+Crgi
nbgGX43dSXSVVQRAhnL8NFW9Wt5Kr3jZa7H+pFjpOJ/rhpsXUoIluLNgalADkiIK
VulIMpYdwCFBEttbVYFqlwwLKu4WGeNySOR7bodZIcRzxEpTYjtlJRdiVdbPc7mF
`protect END_PROTECTED
