`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ze97xRH/da0jhMjoee9Ea5brvTlP5LIuT/lvUf3XB2P0wbFkJs1i248uOnnzNyPW
7ekyEk17vjgKg21j9erp9HvfXDkK5UEPynX15PW02iIIX6Dg++heb5L4Tw0RMN4T
E8B74YORl3ptoC1RM9SvLaYaqe/TV1a2N92etruP2pKCeaEpA5Yc7B0Zp8Wlsr9o
Y6+iA5T0NBpneF0ostdRkzu4NA/pKHgVzSseEHsDrmnTC3KN+b7IYe6J6bTYF7f8
+T5LVjrdMi6q4ay1qCjbgUyqA+IQZPapprRcusDyR8iQ99gqYJPfNvxfAPwCgI4s
EOfP7Psxn4FVCeI8V+zyaC8iNn/bbYTUkdfEEpVWKS7oeFbNt6XzNonfJs4f7WL3
iryQZtjMSXvJ5FbKP0lgi9UPy3f9cmapYiSXEDiN8MDOrK/sCaDJUyUg1o4kPiXv
G/5+N8a0blagDxvfkSMNlP4fhMaJuunIWuqTQqHmT+KWzzeXM7RGh3Bp755L8qAQ
PCKVY//vcAYxboKxsz2vCrIKWvJzzMznrL46Q09dqydwN/kQXHaXDp3HCE4p0pEb
eA1YlTQNHwBbvg+OvzCdqyGANDUTLz3ZQRV85ZbrUv3a35UFlw1tAmjYo8Th9uI3
YigYkR8ABwy/TTUi1pDPCvtNFRsPgeBOqSurMzv6a3m9qBZNMxq93dHD1jMfWG2y
PElR/Xcs86tBtZYoDPDlNZN7FqCXoEi1SQnRl63uJYjVdAyIryh6H3S6TJvjKXvx
3wMrLGUto6/RsWb0uz7dug==
`protect END_PROTECTED
