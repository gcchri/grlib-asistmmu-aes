`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FouunvWwb7eJi+zFuWPr3W+I2O5a9niQOTrzWr4wDWrVbVRpbADQ5Z3tLJQb0/gY
pJ1SG8mDrK+2PbX9E4xGNDpdM63AWpY6wrMevMwtEI/3dLVZi7Oi5dTzYICs/Vyd
EsIQisvyZW4ugxYOlsY0dPmRIgZ3sWvrGC08t05t/IYtjsnyLPYxHRjwTyK8j8sZ
EWNoAgO4cg1Mo++iHcVpQCnJJhd4AxvXmmSHKLWZSGRM0XQVMIta/Syv9dF2usls
vmTL3R7vLQfcGaGYMvqi5G0+iFe4MB5cY6gudisgIlKd2yfvmgSsyZpq3RohJVHJ
HnI8aZkfIIQFXnBiPF2uC2gkkoFplQOre89I/OV3N3OXxpbDD2HgHZW3gVPZ/J7+
lGCwLBa7Ox0fpLOGohyB/1Z/mD+cX/1SwKeVuIIKb0SeATeKLtYn6dCuyucdiV5/
gTC5cTi4UlOBghKNYFjJgFRNGAh8e83UKtn/TM23npiaQamUnUQ4s9lsxgZCi26B
OsWEh2F4YxafvonCAcnxIUmVhLUnKJw/MxhJhxTaDR0jdXrfiG06RIT/PXa99LKb
N3VhL3aSaON4ZOr8dKo/BUc3iAb2aSb/QpxdXbFiumrrhn5CyxegtNePpiAtjK4r
7GjpdUiE6Qa1k1qGMsWhiWo2t61pi1s/I2lRzpSEdMrfwBOuTfTu+7vx8Wm08CPB
hqIKZkAoagzrIinGb8i783b7hiti3ZqMjBWWWHDRNilR+NyrPE3kNbGAtLxdwyXd
dFQhrDG3SbKUrOh2OuadA+lN+qhnkeSuZNOs4KfxcS2/bNLUjaMpEnVOlt/9nkmA
X2iEhxC30cwI9jytU+R0HVnBPU8do28w3Cp5X81gFfPvrfvSTWOjJOcXIlftiXWy
G7N/A5vgU9NbsxafX3Kngr8zJTNa+dzLPsN+M7tDJ22qrNwVncpGy3CReCFcW/GR
dSEpqml0eq1OkgQd20vEkGVZaD3aVYqtorgwShfwdinPwPnwzNUyn/q6XbPvclAW
oBHQO+2euQMscbg8ZVJPedOxAimmpGQGjj7/QxhTjvFn8SEGSlWseRIAKxUu85VU
0SkiJi3rfECQmJSaQoqPCCELEWFAKiQvtcRP+I6n/nmU68Q/An1sKYpRg6sF6KQt
e0JlnBnr07jgF/hCP7x8anVy4PINAgZTZORiR5pKgilBtuOL6Sb4CDZwFJ+hHoab
5HGlJQSRYC40oroGKRPiqy36EjZF8flVM2C2GXiw7cdVcOBd6Uxoq11tl8w1ZjtK
7li/nzFYdI1z1G/YtCTTfSoRG0OU0W2lzd/JrjY2dOXRqcYqlOAoAY1D5kFSKzdi
FIT9BUAYXm80KZGVnhtKFA8Oqv7lEEqSsfSz3nAKn5iUYJMg9/0a9R1u72IARauh
lziVufcOy2AklIyqyXuBif4peh/T0YabIGk4ew+lb+FkumlcdAt2o27CqMv2Fpl0
uRK00EnleCenWOuD2C4/M7TIAjGQj8HOHOL9hxf2TiRkvwGOiw2XmzqhDaR85DAZ
4cEQy902qFDIiwDn2x6lYY/vUXSDUXWyj9MizxlNGqMgviQH6S/zcvaBmv122QoB
6mUNu8Lzc3fkxHCMR9oFV40Fz+4XRAjlUCgXBVR3RempuFa8+yjcs4um+ZUakug3
Z0qGSDmS8I6WxRryZo/I/4T+VX8J/wWUMJOlI1Yf7MNye+muzefSlGRPKoK/6BZg
HCqnQHPmzyftz0iG6kSOntEDUrVN4G4s+AebfWzt5o6LGI/QnzUEO1sjWZz46qcx
giUEhkJugUjAyY13naGX1QwIn+6w1jyQlTue4UMvEed7RUnbxNwAQHbOQkZ8wlfp
i62gYU2FFjAWtunVl6ENWixS6oThLXaIkyz5lPUX4s+SxHGUwTOouF1T5HJ3tQjx
qUWm1PUFg0q1P2dWmTCtj8rAQGbpAxm3DYVmzQW7EAiJdGh3q3ZnNjU4/CwHt4rl
tlwLo/Ql28IqwvTU2SRP2HXcS56hybpES2S0UWy0u0CdCnUW6WTJ/VnCkAviBD1q
sz3/YaNUjcSlHHoEfsOfPoL0RSqVkH/cLo2ADPBoOQEmcLZofpuywHykqdOjZrJZ
WCyzelUmloWym2y37YMcLIcg/U0DDISEXH5wqEBKU/6BYPW+oaet8M+gLFjovA1Q
mH8/UpxaBNVG60lqnor7gjG8D+x1cFNroAmwdSfhtdWiR8/cCAXuDX7T/uKe2ndS
+zpAuL2R/1Y6ESdov292+rqo5cE7NLDcGTd5hi4IOczCHQPXlE/GUuWP6iB7EiNl
mRyXJojTEX1C8iSXLObOcI4jNRghY0KQmQO5GfLlbLZfUsAeZmlpkiPIhsr9qwzX
sUMDCO3v7soQMZxEV5VgctvhAewrLAJNQ572frZEvuB1jAZDr6KUTrpoT0gJLLA/
jVNN8O4nkhlJJ10M7fbWSH5fuRdl+H2QQneCl4fwPNgRLSECymHl4MK+69tTb5IM
9jDJxsFX/Fwa0zrJnGNjdQk+2eooE9VcFV7PphEcg7ZiUyFkS9uLYZZeFCHcGboJ
bT4ot7yrgDaAeWUJMclaG6RjpBOkoiCfrhfzjT9fKH057AiMHLHmwU6Hxi3tbWhh
bwhMWJsnKhpVPzR0FJkgG3p2XrGZZ8o8YxB/t7td96xCSRKsXRAf4jul128RArip
5R3M0hSB5sQyDn1xnDWh91LMFCuzEG2Yq8UPyo6YrfTo1mbJ3kARdR+4rDbzSVgt
yfOt5vnwC58IMeTNWC1yf16SFHSDSLCbtwuoxrcOX8/QBLkDlt6G3pslHtw66nz8
fDg1pP1G0s6br8MUMJbvjUwwfz3iyHtfJCKhnlfkI0OJEWT5nMcyCHrYzF15FcDC
foMzimMsNzgGq+5TFBll04NVEQkUVrbG7gY32HjStUTbLGmapWz/EbhPt+jENVEi
4WtjGC/DqUKNTAZx/+FPiayST8/fgPnNIyvDbPKwjS/qAC8Im+Yquc6T2rvBV3KL
LV4vBaedLrXuhnsm82uvaoyC/UkDpPMndVgZellkxuzIQ0IvVInZZfSuEevZeXTa
ItNZ421WmgjbKkdLpbC1j+77u69KSXinvSD8p4BVxap2Sge+g2M6Do253tRAFfQ7
59Zbx7JfgH9cyuh62+VzEZ8cQ+ktUNXjl5ifw/UF9ZWZDcAHlzPaJeiKOKHowhSa
h9nqDEjaqUtfaKSOSOvvUFlEVnVs6EWnw/J+tR0UOfLuEarCYO58PeAEaDN8XkWj
2HpG6r5ng55+q+nH5FIPpFG4gZT6TJ75HYr6+fslOYXYhi6mZdp9DbCc064dCOr9
dNagLXfOmbWJHF8tvryDWCii9raZu34GIZ6B+3RBzRBT0s3BQ1y+1fxVFTBpw2g2
7PJv29nt7ao+XupzxehobyOh7lVu4cKDJO4OPJ20tusSMDFUzUUjEc8oopPNnG1w
vj4k0ReM4iCq8IQnOHPnfqIzIfETIkp/AWPt0DnS2TWDAfJiqmFZ1anWgdR4X03F
OD1jZUq02iKNq8MrEX2IFWqfgf5fGk2YLPoVnIoPOAahOKqylQqwoCDe7T45vuc8
d1/q/woSebD/ORXGLObI1Cnmz3u64CLztMJWjXNlZP7qCYLDZwFhq6PyjvV5Oo2a
+hOuZ43XDMKTEu1qmwW2pa9wOf45NfuNKZpbpTi/h0gJJkD/UITxcjg6D+lUy7jQ
3JREoA2wbkXIBmUqBiyOz5fBOLK/OyGdYVeszhkNL12c5bzT8/1eAH6K7tAdHjcu
RWZx7h301lMumNsIOi61Qu7jhqhr16+j32uHLzERJadL9UM4yQzdvy3GDlCmuSf7
N0ir7LhM0v/L5VMZmMiJtxb7PB+9d3+B0CPThsCqodzo8j0JIIOtqNYtc7w1o/zh
Tx+6yehKWRclzNYsYcPsq4uCSPJ97fLKj4kepRV88bAeei4yaeEIWPSv9kBkayqF
X43tI7JVR8eS20GSt+iW1ELQBXcSNh92VIWhk5MKa15U/m67BdGy5fePrBVWeRnc
t/9nT+2I3senN37qceh4rwe023AvgZP1Ilb/ThJs8kzlhFTgw/0mG9wrfcWR4Kfi
`protect END_PROTECTED
