`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sXCtzRNvnZ8aw+oAo1PU5NNazPwvsWdC1m+188VbtYfK1ze2yPpJ/aqouc7tSQ/k
fcCCRCZ/r4dRmXDtjsJ7dNcu/4gA+6eeMOR38Dw1BGgEJVDM83YWAGUncAlP4Jkz
SEk2UVjcrAcYODRFGVeTaC4HZF6PEd5uJd5ZDraWNzyCles8wHciIcuSSq8xOkA+
fAbNRVq6Pju5PuaxVbJLxRTiSpuJMfN4KUqp/dV6sKFuuYWgxC4OsPVIp8zGTPVK
lusaKNZjSVgSWGpGEAOJJ61mUByOotRc/k8f91xrK65l2YbLIr4nUjy8E+bBbd9u
+/P+p0hoBazfGhNNDXxdfCn9g5slI/ntqx4aKOrtTG1/rjsg0IwD2F1DSsxH6e/U
l7e54KdaJtMqb9H3hMCM9Nkox1pGQ/ytORMPJocU4LvmhFGsq7iU4bt15q60EAR8
5xkNRrBiCOxapbmIwxrJQrXtlo6Xa4kfx9ie8h4GZC/Mms52Tz/rdvuLVqb5FAgu
8Qe1Ztu2mw17+E9uIbTk4/QdgtVOplZwRwbyBkN5l2D2EjJdO9GKFrvoJ8TFR45q
BJscfj+mIPy1ikGiDEvkAruBQ1JEqQO8UcqQvpOyww9RjI2trEmb9ydzkSeirteF
1sdJmwTOCIBD3s3dXudmbUwfupca8sFTlFzoCeDIU2VMyF2MTCDrkzN/89KYgaBu
J9p5KMRVsZLITk9cRp5AVuJNMkgwwQKrlhI31fCeSksz+h3UaYErLZMYdj8GfmUr
JZDJx76pFn4tPDF/uLFR4oJo30OXUSrU3R+TkBBiHdWNh7YqNgeTTDsnXqrnz3Cc
1TFI8aXAO/MNxPDuGVzuEI67FMA2u1oBCg06FTQ9wsKAOTj8gcZK1wnvixZAYbgN
Jt+3vCTkkTNOc+CAIg7mdTeajYwLSVWfWRJMM2Z+SV3n6E0Kx4EToelPjbQtpsVP
uGvsv2AO3aKjnyDz3Ul7JSyfTLr//74gxgnmHAEXBWi2X1Fk7TdqoGaabzOOdgJX
nP5vIRz9hHjKOVLqN302ZyseKoprWtRB53m1R2PoDMsAYjnCbkJUpamviAVyZF5d
0xYwy/56+eaXSWvycaijeSCzLM/3Wq0uykVYKe5pE77+lqv54GxQAV/veVRLTmth
Db++eZ7BXmspL/SUdmB7kMF2XieLjHEUeKbH9eP68+2scBbYrP8MS3bFlZH7Y9No
dtO34Leju2N2rk8Gi9xNF4rLgCjGNGvKldNmBjWjfHu43/h49zLFofi18aqgBebB
xFdAN3iH8U4sgt15fB7JxYpf/5lDEIuJrSe5H0FztzQLTMFmwhFWP4WAN687sTsR
Q0kdY5bohjQX67vNQAbBId2R++7Kea1VjabXq7dL51pwsM3ifOlWJ1DMtA6MuW9A
BZZ0w22i1zhnOv9nE2qlW4ZLuPuJDPbdvqYbkpXJACA=
`protect END_PROTECTED
