`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
caljOKiye3DwBJOhXrASe3NANJVOOnZvbn3PTveCz499XwudDmsiBFD0bk0zqNOe
0ODn2gmTkLJ8jKdZajJhTpd91KQJE26vwVf1w4QrqsXvDqgJpOnxjHR/RPiR/FqT
QekynVhHX8N2Xj2j4hEiF+t4/vE58P4P09omQGduvBSOAzbmBhrPA4XnIKDFeYOt
6eKDEK8qedzS9WwfhFMrd/IusVtGYWeRHKPLbs3dp03Lo/ujtTk7aTsmcyr/M6Zg
DwpMjYKMaw8LougWhWlC83kBMpxd58IlmSr5FjNNIxGx8v18q7dQ8SmVxClOvFmB
VNz+kZrT+wRAt/D19gn3wA==
`protect END_PROTECTED
