`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SmRVAmAUVz0+7unt7WH+Qo02w57z6SoT3a939uK5bBGaX1tOjEsUX7UDnYtlDBfx
E/x16VUbWqmrgKFqe1QfnB9S0qu7kL2o2FOiHg5YiBt2slOGUYULmgq1cvfRQIRe
RKJ5UD/bUqEP36GsF1D8tp9K1RTAgmI64gcqtKrr1taD2BkJRMmhji6Mk1kNMXpi
MIb9zQ3ktWmi1+rKBBkdsnKiUOE4omexuSOXlJj4/sEeo1PEgNjjF6HQ8AgT0A0X
+B8MrOWCLN3zzXiwy+N2ezdaTO0y5zs9x6fiSJNY1ukddL5nP7KrEsgw8ikpRUnU
Z2iAJLl6rpPx9WyE399nVHSD9xUyR+bL3HsU0wfi5vJuqzqY0bzKGSQgdTsyLB9x
g9Y7tJYgoGSIWeRKV7VEbBo/dmw38VfyeUgibY/7OxdfmDrO4OadDA/MyxT309Q3
bkySDVcxPlL32nG55WZTNlGjzZF3n4Ge26XDGHR1DN+qDUnlqYwtzNOOYZQT3VTt
zpGTgOYzoRj/rhRSsyXhisMX7D2F4amwX1/n+rKEh9QL1npYyAfL7zrq7zn9CmVx
wjxSNCL+rzI1uY+ZWxHC+SvT8AmUm+scMynmiA5h+cjlqWSW7wV8YhHmDjs+q3fI
FRNDLZ2lB6IMfMRSUCuVasznV0/r791ogarq+ovmPBHsC3E3fYKjcmwUEhi/rN8q
2hnFli4tnLG+dkLGwLpp7H1eN+7G2fADIqaPRt7awr5LeXMmPI7adIxtZuuR9eZX
J9NVfSqIZbHcmxqPPrG5Vhy6w2cPY6pMEUJRqo/nGl7ZT9dmT8HZrSjVFfGdNGZJ
2dXCQ7deaVQECyBNALI8uzFeedXf4HCMJVNDUEeFedMa25lrIAi+S2HzHBI7TQlq
kTiDSKo+UU5zoT15NqfaqTXnhzpCQ8xsd5/TN8kZyMJqbcQwli1Gc/fnqBCXJ9Bo
awrPMgzwGkFrOBgMN4tvguhLP4QnwGQJkZprbCiqyBxgHSN//PdLe09zcQW367yQ
U+my1DhDOAg00I4fJiN+prcbxGFSGdDSd+d4xGMZLLM/KkNcEVal1OJLYIVMNqnb
jMFvn2fPQCD3l421qm5IyhlvlgfUuWqT3e0xH7KUKU90UV4cOoDTfQ6+V+ZuESMw
Bo/1zkx2tdvDIdENJ1+Oti7g/Q7kimyDRIEJXclnF+IedADKIKukT36b8FETRwzT
gIeHoyytUc5ZE2fUXT79uC06ixZbnqiD7utXf3Eq9iujlEpp8J5ENi7xTWxEnXBU
lIAUeYF3Sx6D9mTJvZdT0Pd6v3k2LD23WxqBJXXiYN/Z/4jqgF2guxEgeQ6If6eI
HMKWsxlwltQytSNg5OT2QwMf3G1i5rXdIdn+0APiOQs=
`protect END_PROTECTED
