`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EYAuLI6PIu1OmsEs/5//K02oL152m5DQeFYCwTDmuXo5YABqtCmTUSFwMxgZ9Uj2
S60QXVEBgVkWrR+1cqW57kYvOmgmPhoHhZwDH1ntdnLFiL0YejgQBufZSAqGo3su
gz7g0avxZgQABvAp/yBsA+pn2Oj0Fo4Qc7rvgQl6ZjRplTKsxa8H5K+TSj1jyvSJ
YzcQBIr2qTq4wPIB7/d1gal1L+cXar/xolJRDhvYw8BlT/I3+0A0I4TofP2Jxi+r
nrtWQu1dEJgZajZJd40VUURKuvgzGRLMhBOLsntry9/wLNZORVuHI7rkJpnkScXJ
yqn9mk3YLlM/Xtok3HOrYmKqmrr1ypeEbfOJMeUikBg=
`protect END_PROTECTED
