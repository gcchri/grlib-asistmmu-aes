`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rM7eO8d4W3ZAn3DqJ/V45Bg8OvA2SNGpGhJOhMCVlyK4xt/zS55GfUB3Nj62rcxq
XIxwMJmFnWc+KVQw3Uox/CBfhV6Q/ematryxO441N9lpCt3ORxbPs+IkvHBWOwnw
ohRNSZuRzKbfclJR6t0xkYJMY838rGAhbWsq8LSEXShaKKlP/FsGb0dtk03HLJwk
EVhBLa0KxbhIiumK0+/ptI8i5lZx1EN2SVZZ6jrQAUMmrfM0myQ5W30hzlCAtIae
x0DFJ9cbxcIe5OotSEifabroABLmfTErDiP209CU7Qw24VShwAbWKv9IO7luVMsX
j8wgAlotLXY/BwtgSSg536Y9z4GhBhNuQ7wAX4CdWIi0MRIQ9qPJDGbBVJ1tFt0c
`protect END_PROTECTED
