`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9IfNL5JXKPrlBR6EQt3wo2eN5nHlgWyAJHiG84QUEypDG9zG0+Rt4uZ0qJUo2KMa
GK8UQ159LJDWSnBKvNo/yaOyEFWMaInU7dVlb6aGMh2e9buL+dWZVOOD5oaCUgMV
KHjIKVOyA725hrhtaTz2MjSt0HK/QwO/vkPSFDHpTp3YyPR/Pql6CLzwoD4HHbzG
v4ENjh3DqEgefJL8xjcdugWkuBLIdNCQpKRplYcXBC89I1BFt6XPJJpwEiQnm3Vb
ly5HDwjNshaqrcnDkjVvNjYEnsvh5+Tedw4BW5BrhimBtruqz8XNa7g0vB+kIn3I
KQ5xqoDwaVpMV2iDvnmq3c9c2ogke4FUOVV6XNIhAhUB05ZrljZt2IzQ4D/MX7pe
Hq/xP4P6zeNWTJhCjTkQnjyu/vzjFuIDFsQQ41G96at2C8xwbaoF8untKTeMn1XD
S+gFMMQHaKXK/V+ms55Je4vhRXktucTNWrvf2/U+YWVprAr4n27XxQMgPtHrUKx0
xk2YeVZkObyNHrzZ8AwcZKLiiLbvke4kUtvmao09Ap75n/hLsEbBbr0Og+9b/f98
iZ87ZXx4De2z7rlMuNF2uBRgm2CXtoQ/1qJKld5H3amXJnDxE0HCXH0oXiY71k3k
xzir+vyF7v2bBf6Z4SqJUan7FtuBz/GT2EfuoJIe7dSLjFBpXkmuyfIl6oY75jGH
SCXrjO/6pQs4ahnZMGc4OowF4lmBIZjvv9JyCFtmVVOUdSmt30rKWOFPuJw23pdb
rbuqkqXrfg+lt+3v1b2boHdC3OA7gL1i5rhOu1mBlu6miLlNo6mhW9M+exHP7nIu
2Ldyjw4YfRkg0O+ddM1rsxXQAVXsrKiGkb7EfR0eAVcMoGSNRU1qTZK9sNZy1KYC
3VWbkHviZ73wL/MuzSlEBV1ekCXR9HAiFBgR0JrJgsf29X/tPVZ+9x0I95/fwuDS
NNQ3U4jjV9/1KR+freoQDc2mNOeLsKrkenDtUPf8bDoglgoEt9Hm//Gap80cWGO4
ebXwdge38x+wjt3nc4FFC+gEkd0KGYgCjjP2nJZdrXZ4wmXv2sx1MoQMD468cNtM
xBeDFp32CC/Dp4zbEUP+LBvDCj3N682QiwxM7msl3ynTYMdr2fUHBcaGr845iHzv
vLTEtqB+WMTbvJi763n37JREJgE7dScTmr9VceMoJmRTbAtjQzrN/H2pbEkpPtc7
n6IjFmvacOnerkFGvMfQrSPVe1iuOdbCHngUBMJcO8W3a80g8++HE4si06TL8+bU
sTMkkdxqMxbaB7Sfn8nQnJlkFTPanBTB0hkTkzzf7heY1O4Zi4Fn3XdvmAy2F8c7
A2MLiVI8e63jQZs+z1jXwg8xt3AXnTyo9rX1XApdvE7/ttVvJzvBUIWnPlkNUzIN
+pEN5j21rm5m43MJlLKsOzBqk0Lh1Ke5jpN5Xwh4k3rw8X8eOKsz2cxruC0EqH8Q
QyoSvMz4mgYyI9c001bOkP1db+on6GHevqpO+rg2wshIBY2MRLUR/qmwvR2luPNF
3kw+rE8OBOR8q519V2M9uOONhqkEXcE+PsbVQ4waKO3u2EqxLlSOJ6PRhwDreaZE
T/0EDm4CeLFhNY5J+juM55q4WvInxf26BrkZq+WsVKIjPQpUskmpyllQtN40UXWU
R2tx8jTTPVvgMRbJ0qjHtgDtQ8jRQQf7mxLuitgIHsdggcze0QY1n86def0dBwrq
LmvxPLIxnlPF1SvR9ZJDZg==
`protect END_PROTECTED
