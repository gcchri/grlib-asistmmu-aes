`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oIucfL1uWqWt4Y/k79XEcv+uJxKdQ6h+ZGxovSesXH44EjCbLK1VsoFq06b0q/4D
jy5xJdlAY93TUKr+71db/VSKMmlT1zSe/spV3P+nHMdv/JqeZ4ZX5meJcAGSdhlZ
S/Dk5ORPv6dfDt+Gq4uZuS0/v1XTFrXW3vDENYJdDeG1uCppRikp6zS5nQm8alFM
bu/P6M0P1tjh0PC9HETiIR7jI18tW7QR1cyud6jPRIJzKuEVyrseED9O4tilQugl
CmPEQOyFYI2hmrK+Bb+IAYzvUtLJc7Tw/FsuEg6wlvvwcSoZSjZJzbURu311qXR5
jHpJlZaL8tvzyXXj5q8xsDAkj7AS+9doNUKgDLBDxOtNS0sVjd6++oAw5p+r7dPC
gBAmpFU/Hn7p5hKQRNMef2lxZzmw1S8FjpsB6LKsnCr5vz6GFeq0T1yx+5tuVtsV
WuzTSjpmYXOJkilaWpk7QGtBKEMsLFvEvbFWgRdF2Jb3SqioxdzZxjG1ICe3Xut6
ckoVaXNCyNdGx6ha4Y9cFrL+d7xt/pVFCfKIkEAEiO/rHi0Neb4+dOgEJkWGjyPN
hhSh7U4X+gxJY0ApnHBrd9zCr0ruiuaG5CrIgLm+zRt+0xCd5Ay85qzHYO/61vlD
MKGnzdlEqvfMRbx+pW6JO/LTFC7SQW14kp8vvMnI1PvVBgnU9L4aknQaIplPs+af
YjuFWT4d4TbB9p24G2kyyQVvAU++njFCh6DSXajNPQYfVm/mtQRRhcxhZeevJSMe
xolAbNRcswO3AjMGB4JXEDVTSb3n74rk43smjo+PhaViVm4oYRB44bOK3D3y0Mjc
ZRnuEjpIYKiIxd3o2LpgoY83iw3t2J8g33y/VeJzKfm8Ci9OZHjzrHQ/JyEPKp6b
M2CHV3+QWyHqNI1kjAeXLgB1kZtsCiti5Fo3D72sfYJ5qAhPqQF7DejoeFidMsoY
EVbIiJ14rTIGuynwL9mglQ==
`protect END_PROTECTED
