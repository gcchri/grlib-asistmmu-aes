`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XGQij/QWC4JMuzmf2lQ1NteT5PdE5tM+lq6B2ZBKzgkRoVp1aAR5FaW6woaZVYJF
iV3DN+ZuucguEnuYI6FagrQKJl/+FOu2+76qdrKMCfUZaunfCCyCJfqVbWp4toBH
JK3i59fIsfijvrUFbn4mnkSAX2mniA1MzRzhXiZgxVBSi15tnKC3ey8mr+uNetJX
pLK6glzYasWAVRC1HXRpZ36gRmVCXDZ8SSw2DWfKflKBS1Fdjjm0ggv/33UeUys2
wpUiL6G00UiiXTzRa0PLTo/uPeFla8Bamid4syOXjMh7u1Rmc0fEnS3voMRRX58d
3gS49AiPtUmU+l1V7CszDpJft1Ma6iqrT3622/DJiWWB4spW57o+UoYO4xy4e2Pd
AmF8hJC9/d8uioUsu/KTqABXsfPxYHSxSahIrVdhEFU=
`protect END_PROTECTED
