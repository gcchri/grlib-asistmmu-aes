`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kZooRIkKmB0lvfrmoJLcq5Iq5KccNCNNLekM4GMik9+7pUx58aAhnxObjmaf2VBW
Wckls7QVbvmvRaVl7qUTEQn4+6YOjAjPtojYXs6DfehUTp2S3ZeAA+Wrl2eXoWmE
Hgp7dA9NTnbyof2jS6BHdIq/kL4bjemOvCcFreW0M6YZLESS+FpGIm52YfGukJz/
QnXSXbl4zqIbt7BCq0IdgAjHOnk60gGk33PShVbcLDJsZG8PSCciewlGaKROkUDj
VFAC63b7DmtpzedkgEZENhYfMJgVc3ESvIx8hf9xOF6jPBvDGpqrTftk2uFXbRhj
gU29vXXJ9Esc84yrSY7AKcJPHGTxiiVOynE/1PH/OfOf2BVLuRC+8YicTiLxL6dz
qB9DU2VtUqvSsz8EoH76eGf5bEIfAH8VZmK9DpzVmsPlx8OvHhuxq2cklGgHCm5W
VerpYUS3mPE19iHjrUoXXzIIsyMNVXUzdPCsuaiT4BVhhyhU+nYytLvH3KmLbpOI
rYqpjMnvCtau+iPRMhl2mEmfPtwnTLJQLRAiELpm/jRdCBTrju9zJzAMB9Xa89Dh
j946oBZHMJDzIUiq6ajiOHDxUu58S/+mv4Ta7CY1XPRMw2hZC+7MQk6R58uzdXkU
CH8wPg4TZfXsaEz2230rEeLL9TObqXs2X43VbxhqQO9VvDAZZW0Hm86iOpf96zEC
ocz7KOQi5UHLeGhU+Q55+dTkjEY+tpscfPvTyLjIt1MbuJx2DAkaqDozqrGKYqXy
`protect END_PROTECTED
