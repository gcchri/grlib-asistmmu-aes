`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sbEISOhe5na5DcgGO4tB6vCKfUE+bYE3UflfwhS549gdNBIqqW3nF+hj7KsmRN7x
T7bWHUulVftJxNsgTL1LW+BzB7mfH9SOX7WQsf5w1QFweTHN3juR0FsfzxQMPEXD
MVNJsi9aTetJXwaws2EKeVDBPF9QxvIzEX7ue47DCZ7tqrIZrUIfsnQW6964Z7FO
rwmLXcqWABbf70l23XsX6ToIUIxnmp9uzbsRMTcydYjWgIp1dsNhHYxElwxymIie
bTSAnOQxciM38wwWs6N6U6IVEqgb93gVgzibS6xYL20X0d8tLxLF1Kug91BHKF72
hGZPNJJj5VO0wmC2NQGwNbtYCczM4MK9095PVLaOkGGaFFCaIGTmXZvtEgc5KQBI
iyxaq2V3E0a08sbsBB0/MerSRLoMhcebiDGtOwA4qWnChdJHVvEwVF7n+L21Jwlw
`protect END_PROTECTED
