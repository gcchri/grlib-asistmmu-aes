`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iEsYaeYdsom1pkDBvpnjjXik9l4o6fwniN3w+ZRTYLU3m7leGnez5SDRgdR0g/O0
SGB3MmaS96MHFJOOo92Y5HNB+1ytH5q/GY7AF6GD24xEKt/YIWMXHmMTiFSCu5Oy
ZM5Lrp5/iPgI532Re8fI7jpuSlIbu9hflI6pUJSVS/lhWirK2vDuUN6JrxldaMPf
mCDTOVsPO2PGn0Gwy92GAnZ5gKBxDsP4sIBWMoi22VrcT1B0FKcGwK913Ekb1x+m
jz92oW1hO04oUuwKj4sHnIDypNQMx6t7f4vIjj6lt6EBRE3eeGBp3OD3alWCBIU8
sLfmRxRZir1ndu4vZLXRFu5qozdRLkXcZRuCWIV/coGK9HluPQFmum14aNl1asbC
oWyYaB5uhKfY6akMA2aVMnhuXDagDCu3dQu6BRox6kWanHBk6ELm3GH7DwJZTyjy
jMZvuDZYMOOOPu4I5KJ4ewcmVrHIToKtTblYZBGg0T3WFXFfzoCvAP8Bh+LhUMQj
d+4F9z0r/YM7bsYDSKfPugOTro3hfohIE9qr8PyeDAUIqfomD7hM9qC9NPII3wj4
mVP0tyXZuuzRs/Ine7tE7K6xfzmR/3/DUMHjaXqMrNiK/4pKANw4M0rQa5s2QRnT
PPSeR2ePgH/BkGPWCPjzpCdVvLYLZF2peNzeTXsyMIU=
`protect END_PROTECTED
