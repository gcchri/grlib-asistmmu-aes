`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ZlRH0h7YnusoCkale99JaE3s7g4JSrRRci0QqPGNEPW49jkK3w53WXWcIpYcAUy
xFx5Hn6UTSRSWC25/NtMhJS6hNHIzZBqQFJGsqyLNwy9wyLv8NJx6RoB7vhfRpBK
2ZnZZti/od15wSiFy3PQmPoiMgIssAfECuCOw72tQaniVQITczacNnoYgvQN6Dkg
YdnxbMAI5mGcDLGUqDXez4++Afnop8KTSirO7FLgGjDHD91ahP7hRgirViQWpSaG
g/wi/ojxp6QF74J5vIqdI7y1TAQZK9i543XbVhYEPCIOjYb+Ju323Q8vrsKWTt9R
xo1gPFNW508/dgjY+ZKWG59sgqhig4n4GsARtLeEjYNOMpqL3QWjqqQmdyBpi/wA
jRRN0AgXIZ1DSTqlVgR7fxoIX5ECNm6iAuK0VB9SwnM=
`protect END_PROTECTED
