`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HFPcjxlBpI0/NN4tSxOEYDm8XplKMPjGgZ08cxirtojhAgfQkFvSTtWGYphs1leD
vgy+COMVVLv67lWysRB1mx+KJyuEiRV3X8ejahO+aEeNLIZck2sHuk0dOVC4iLU+
G+UfPbG0Lvm17c+KtQsZfTRCRrgFpt8PTnVwmEWOvOdayaLAqOhjXLvT0Mcifwgf
9krNQXXJL8wEXpwH55f2es4pmIHQvqQivGIzu7dEJDYWGm0OFolYOre6jZRpsN1a
Yy8iABq24CbsxqRuIYWc/YIdetRFr/VjKSTn8ljCu1QCCjZjwdZuYuEEKR9hMXd+
EpnXh97aQ8QzLyb0osSWKg==
`protect END_PROTECTED
