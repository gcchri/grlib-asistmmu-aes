`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ekMUURYBAwvKGIps9o7ezbQYOxMZFdhLYracTfLCRUNYaVxaDxSW3OCwFj36uivP
RIGQIEJAk5KUL0QmqWYZml5xuMokMh4hcBxARhWRJhm3iQGEyf/mwWGrtA7Y3LXp
isuAuPLDNGW8ndr1JbTV2E+QADvqwd9mEHQpa2hJ4+zDhQBuSJ3AZONDgtwg6a1q
iZSB4ZeMCKQXqfgO3Og4G8or/CPrt9Bu/za1EOmstwDnTo3SIJDqRRjG1GggSdyF
26+prwm8P0EECl8V3CAlnyD9OhYUvzUq75UtBV/SocdnAGodkRdZsynlUbj4uPJF
K9Yz1yVSMO8Xuu+79GzWmkL5LUl5NwrCx4WsOEyYbbJcuYV9FPljZamDzqTtcGoA
b4yOxd66TrCBF64VlCnhhB0Yq/pnk7/J98rFVbdRLf0hAoiBoS4UT67p0SU7Co9d
cYBdCX0PeZNMWHvAABXVg9d1l3nK2PVivFPGMDjkCX1Ny0qh5CVJB8fQhJ0qMs7V
m1pcxDUzIgp7O5HqN6C3R3JIz0E1bCQnh0nIIKXal6vpxIXfWg8aHEXJlxTPr7s3
PD+dzlBHf3HPbxvDjthLJEz0khiWJGOJL0QG9y+YcGfZ5BAPHwuk6M2Go5AH1JRd
SZmMpA711ZQWD3lWb9sNf+3Lmjbg+knyielw8LbSVRp8z2NHmWMuU5WgPjcxdBj3
lh+qVrNMSHn4N7FAWCEOStwtTYX2gCn852jfz4lSwB5+UnPMPmSdTQ/i0nuK/x36
2Jjf3aUyP9/IUw6QznC2ugzRkm3VC6C9SuDEpYv/LkojhqhdpEh8sTOGXLxQMEOL
GezyIcHN9Ij6GU9CPAwj1OmLqMxJZxJ8Y0b2cRAASOS/BASNINDGDsz2mC4E2juD
Xdpn30F20gSVv2MokbrUFLQ5cBSJUc52Y1Opg5L4dV/bmqNE6yDHNdE0lEPqljIl
PQVignlEcESCXT+8BYDUizL4Pr0M4dHaAa8nBw36STJK/bHb/zhU+j2utExRMU3v
qGf4A5Y/qtvAX+Gn4zljL8oVgOST4TZFHTh/j2S5tFafstHbgvuGEBNZzihtAUxR
3FJLqb78F8Ss4apHaWg8AuMg7FY7gX3YID4Xg4O3wcID5m8Vv3tUFIyIjWs9oJbg
R86v+pSfmvcEclwHDBII9asrFuU53oYHdusOq9w0iHm2/gHACBez717dlMNa/ruk
9dUkwxmkpukUgw+5OF2gt+cV5PN5kQkIt9VIJ8/w1SPyABYtG/vaOnBm7bZsH7Gm
LYgZvvJsunoxgd6k2uWNoQ9E2ItR0TvvVshZtkpneK9NJ8EPmKZ+Ve6cT3NRnR2E
PbTuotBDV82p/6NR+ij5S9Af1WxN5S7Z6I8WwUJKPnQLy9/GNh40Xn3UUEtwfGcf
bfFuAP/m4VQQfZHrgRd4MpmjDD/krtcgABUXqGBPkrEowkHgSwceA+FhB21MPEt2
CasnjKXPs79jns+egCFV8CeuhDBJ8BxFsPKcqELdkjGAt6szO0/a3w0paAa1yJeu
JDG0L3/eFOwqfZR/Q7ks+aJPBeDwW2PHOI1L6gzVsYddo4FJ4akAFX/adZDVjcos
855KP2e6xAmKm8WMojdgeomTrwsdBd5+bWgUJvTfS7SLjEEnusqPdNBIizK3Tt4Y
RAQ/Od2e3ZSy/jP4KCKr3B/iXKmGTYCcyRivggXCiMexLS0Cz7i4UEnKVW5HKkSQ
uDNlgYh0qnmv+h8imf63og==
`protect END_PROTECTED
