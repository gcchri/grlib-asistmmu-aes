`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VkfvNLZTpCXqhSNYN6quNSw6ceyTgUYebnAdnLhXIRCaB+Qb9wXyGP7aPQa9f0Uh
ZFyO3drQNO4mgyH0nqKcfUw7aumLUCWPhWl7ae3TrUVkbVfYdX90twgcLYW+VXUV
LMbimrk37NpmUVNdaYHQUFMcSGyQx3YvIz76T6Mtlk6nJmjJmVhrgk0B89XFyX4V
LYA75d4bGLDfn6FMKNmCiEr+D5MEbBlw/cpc+73oMhPPOKjwt7pYsI4HlP8cNhWi
PE7aDg35zAxngp63W6F/D3seK9IGo7psW80UkuLfs5uYQX4Yd7+ITR4AHuB8ugqA
lkaIWzcy441T3VGRg2at/kTe1RUgpeUdr1pllit6mlQshzzBsyPPUTxYbPLLmimh
7/W6K3/AFb0KVxG7qKEzzdLSn1U0xfeNzURkrqqMyq9xAd501lNpOpXqWvnJaDVM
nBFVu6ofyrYWxh7ZMLEqOAbKThZy/CuraHZQJZijP5J5U52wGjnahX/g6+QwK805
u7Sk0jfQ+2/xNIPIDl19wgqIGZHspO0MpoRsXE9l06ZW6rWTrVSxTXytGwYzE5y2
62igDwsDYoiQ+lJriQCMS120CaC0ezO42vydbM5VRcA=
`protect END_PROTECTED
