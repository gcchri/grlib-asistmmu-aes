`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KqH5T3amXNTIc280p0LYRh0ZgWXQQIGtskwlgpyok8ra0vKOWCXehGXEfl5aF0UJ
1eQDTboaSIgGNUgZ37MNSCwxbXCKzunvrvDeFOZ9qtMdMQYjLHF9X25w/jWFhIdZ
Fk4REKcfp1ClwtKhDIMszmd9wh6/LK3UYNIMl+fnIooaF8W90vtOwsTILzI2safR
7ZZtOVx4jP3/M0xX2xUslFjP1lWCyGILZDvryxDr2+hg1RlS7P+xKzQxBLU2kQoj
Ol/bYAdcC2JpbuPfuR6abtbrkMTI0pwkfD2y1G40VEtlRCXq8nqAex+hU3IIoPLZ
YZ04Ru0RGFzLFJOHz3T2nnLA3+XTLUaSSgRjcIkhgd4Lq5T8oaiV8GgN/ijv613Q
U1BGLw+Jx17a3BRhY8rUtZSHq4AxEgvwsLtja96Zvzmoyrs6Nkqzj9NLZaFv0uER
BoskLdKRIwPh8mFFSQ4DVptrsfkXnqWac3HSZLSLTzMCytJcCHDMXileoHS7HR52
QFL30sxBtBRglgxPinidnA==
`protect END_PROTECTED
