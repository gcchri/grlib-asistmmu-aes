`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xmYDAugzhLPWDSfp/SZ0kOLOvq0OmYvXPnlKQQs45HR+JZeXg8gUpc6qZmix1yi+
H433Rpb2Fhcqg2TezXpbF+RhqV1gcM4nDfUUfoJWFgCy2SjW+WXCnZHpM5910rBA
6gEvWyyTSNb6wR7pit9XesT/0cc6WvpbsH2dtRp0iAOsc7eQg9c5DFx4N0/Qy63U
ysb+1OVjqK5j8biDQ4sB7OKgZ4GxipvKusnfB61jBo7trs85rbyJD0BphzELm1dF
HDPd/bOLWJ6T7bEZO6Epb7dG/j7T2+MStmxdghJf1FgvWJOzrkY3TWDqCVFOORtj
rjdTCzQPiIlUidByQAZIeKQxWhoDA/1InGLY7Epm30qxW51m9PMSPHp7j5hvq2MM
gDczb/xo3liJNSQ+/1H7Q0Ecedi2p0Zi1/tJjPq40A73q0lc4KcqlpfrzVO95+Fo
Jn0MwCeTfiEAUsSFPsiNs0fvzvoRh+CXJ/xskU5c6wVp1b8JHHk5JuURaOxCDdO+
rFBw8qO0CrCTU1XtiJ/pgHrq6suPV/yhgdNmiJOMEhuuC9Jn3DRm1XNTFHslPCYE
dyoHWaNIrEAgCkyCZlxEm0WI8yB/YxZv1KFkQWHZH54=
`protect END_PROTECTED
