`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OaU25EGktNfTojbJnxcitlhz5cVfyMlGQfnNuDRuKq6D7Ym/UkugWdWyNyl3Qh/A
bQbsjo6O1IGDbo+ytSgyP7/jAMM5wonrk6Vb3vqWL+dxQ9A4amAc9f5m4Ius8uER
9d+wvnQgeW7rqtVw5YkCcRYgUzrdRi7EN5WQ7rVXOvcrdzNphFfaeQqPDzPHd545
3wHY1Et7wIpNn2UrrT27dMWT88nmHjSbTODuuA0Xr3lDsE5wbSLyLMGrmdQku1to
8ImLXzTml/dMOOVp1zh2cX1rr18U0qBHzgL4h99A1j8EAGIEn1VbUK3SIrqwG+Gj
CcOxeVrN23mg/xVgxqsE17ynF+vdcs9UmJ/V/i2blYvUreVQcoT3ljGgYTsejIk4
URftePW3UTNhuTp4MJRcJAXRxWSIzcyvi6jhoufzDAMv4tXoobC4ysXSnCPQXjWE
2pm8d72fOS7y7YftIFyTWEAsRiIk5wFTXwfTMJG+d+yF5dcBLcehqg+VJOBwBN4/
GnkNii61JPyh1xpfbG9c3Gln/YjnXPpldm9fyOozuPljMERLSVFyTYfjZZ8h52nk
1phNV6FqbId1BpyuuWYOloQbUZX0+P+dEZyXEQxtWhRoAokKXm7uplyTkJvVURlU
keakloRlDmMySghzueC5Pjz2X06bFnE9SSnOfS3E1frWttuimhx70f5UP5ovqRrk
INZbyt6xSQ6ISE4x+nyLsLqknFX6uFZQ3pfGDUj+QIyl+yBti1N7QD1/ojqzfX/F
B+5HpB0P4X4P8g1KawoupA==
`protect END_PROTECTED
