`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bmwlNVhPfrP7TLBsE8dSu94IuWJ/qvJOqeTyioI8U3HjuB2fR60wYIHsw1WScXk/
cGD+KmlCM1Y3lGiaoiAHius9da8Jdt/DMiIVIh85JIq1vzS+QAG8ekyDHQ1iRfjt
DLkQMMe7nC9hnlZlCtmxOp9yEbRLoqpidPbUutRav8bdUExJt/43YD+0NvfGqOCU
7bXPnjy9ZYsVTXnRg6BMZRmBhPB7XZj6dySFIvNNNEByj9nui52j2qOt6CJYo9Ml
5VuHyoICJfrMzw9sGvUi5FQhRv0xGh7HX1ipZNZ+xy0=
`protect END_PROTECTED
