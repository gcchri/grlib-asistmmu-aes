`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v5fHaq5lBTreGsq7Hi86QZA8ex/8eIwYtaXHj3VG6VUSN1g8Hk9++s+gUeTgt1Wh
8lZSG81Yd62C7OeLwHc7dNY8i9f/jUnyrrG403OhSm401Bj71oLCBcDonmcXsNMU
xf3UvlKlqyjg9OCxJMzC5OQbBqMN3BAzs1maHXBTzpCe3agU92PW1t4cI/DVVDAw
uBQqQiarr20z+c0DYwkNSv08qdRXYkyHp/RZXaNdYwJ2t4OT4obejD+2RmwPa95J
uHTf9Q82K0zTO020Srf2ycFwnXLCaxA4YkUZbi3Q+oKZnK7rG33ypPlEctwhS+MG
YH+nk84+XDjkHxRnTZsZsiZX7xGZltaraKT9VHc7riZuWpqOFb4bFosLlQOk73Er
V0bByXNP6mIfyJd8e1eNHyMVu2eXEO88S1i51ZwKD/g=
`protect END_PROTECTED
