`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t+8nGK8e0aUFvK3I5YN5vR18XuNdgFf99ZzEtxvmH4y5k/bAKLJSSA4pOBSbFj+N
moRg2A8fJU9Esrom+9uAAFkbvCOrysTCzOxt11QgNzMVLVzlfCy0YAt0hnS/bSbW
PlDPI0F8/OhOjooOEizXMgffGPSQM+zBS72ZTF7lUvMYjpjr0M1dySM5F1tu/oBi
zWK/8siZQi+7s/Ga+UHOwXalObufOLkPJclO4ksu8LO1hwtbwBCZ01+ePiNKJBwc
79g5qTo4ECb8eZzzgLBjWgT2kxtCRPyCXvmHJ/5UhVYPDtyxyc8+WkW6rnPZ/yLn
WI9EMlONAs6maqgoo5dq9AK1Qm4+sy42flnjh45iCsvEN/58qDDYo1KRtroxLFBB
Vf0AFl/IfQ28Yix47bHo7AZ+2ZnFs6CER7lwGVFE/E+o0/ZCsg1MmnKw6sNwBknI
ZR2mfoZdP0nrnZd96vnq73KZCSjlFopk9Ql2qhKKMPFUjDmeFdG0yKbnYrV6CWYy
/NB9t3k6Oz/vtorJBBl4XDkzQjWaOlo4BCqgXdr5K8kzSQUbuGPLFNlAWR2mrp4C
kxKjNyeZpFRtkdQR/rN5R+JScrvTC2F/3ZLdgCwja3JGp69WZJ8p+DpRjfK/bPv2
p0RAaUkXbkO/fXC/d2GtBcoTFm08BjDl3y26PeIXD4GrAEvcgsyBqXZYjLplra5U
0T3vsvrtFAVDPpMST9pCLtWJbKCa2uAHbprRC/2QIbQymenOUVbnedfG5hct2ldk
T+WWC9Dbzh3lHDBwyEodBDLF4gji/76jKsH+SC9qrTQGhqPZ0hh7/UblAe8WqeT4
gRBT3ceI0wRyiRuz7Vv6liEtEBiwz9NttsZyFgJPiX3jrLDdRjRKSvjoxuP8GjdR
HAcI50Nc1+HhEzHa3vXMlZ+752R0GhB1f8Aj8cT73lsDHUpXOVNGAK6n8JGMMzYn
+MkltQi1Nw61uzon9TBWmi5ULEpFKzJtmfd1d6KtQdgiSAwgs+JH2RcuqCaaSA+q
3MD3f5AKvgI6eKR/HYY4HkKLMgbiGJYIfXGsURBbo51GpMyyzqnshuAOfNrNJEgx
wteakSd4FggZcM7yjtasIYFk/qjP1hNOFcrlunigDVO7RlK2ehOxL/YHq44AnVvh
tqCFB2YornK6/KDKUz2CqhsqjSPR3/BNloIV9fRGgGXww7KKJ/BpUl99iZuBhGS0
UAGLeJQR4iKIXUQ2DHpkc915QjPvwxrQZ74QLSq5KOWsffNWVWH6rFIX85DmOr+Z
IFrFnle6pKgkhcJrcGM7n5zy+xExyKiovF04vv7SK8eWB9TY8fYKtotatJpPOaSi
MRdl6CswqGUi7ZopIZLppzfVZsyRJj0zErvv8lsSragd9RCrwFrzW64AELCLfXax
sHFllpqTE93v5EUyIRXe4Q1SOihOth7R6TePYMhkhwFVxtiU/NkruCdxiM/AjZlo
htCSAlLGYFMcK7vnnBlFb19KkB724gsXmHoipW/KL1dgMOBnP9XYFmA3zpgHpsAw
jfxbsvlhTd35Mo0ZWsUAoKBFZkdU6VdLST8gf7i47dKUpFrJvyoaSeBfMSmiK6wU
n0NQgfdTQxrjZAES5s/E7FUwibSGsie2pYRcBTl8raKu6Y2vTAwTz0bvQUoWwtVO
nrPiVWOfspLjkg0QHv3bm/54Dt5p6Xz1PcqsPFXgapowEunpLuLlhFxElqdwGhuN
Ybs6p7LbRS6hjMbT/eLqufYeV6e9VjqLqkOMN2sLNKB3gjuUxdgv+xrrzFQSDhw6
`protect END_PROTECTED
