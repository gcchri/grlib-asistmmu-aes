`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jaYH6cROkssDX3RO28BT+UV4qJOLo8w3FY0VfqY/ss9xKDDUm0Gm0IYYBe/fufqD
qyJdpSMeMLfpdRVz1B4PyyLVboKsNv8VFLEkD0iYchj1lPl3L/DeRbHc1NNTttET
H+wj06XXSplA+CoVs3salbjLWns9o6XyQc+vCVd2/8KHrRADSez0SopX4USiM0eO
Jb8VTP4cOymrcsxmlSX02MrKIOG4BdkEhs/QR/e3S/p7CSJXKyBUMPntq8ybSDZy
CfX+GAOALO1nvbP+ETBsgLx+WVKx2mPSOGiAzFJYdnYOamqjKKyZt+ZMDGNsGCjB
B2x2SekYZ+cH5Mo+9fnSTQ==
`protect END_PROTECTED
