`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i3G/ZuRMzk1KwK+Hu2yp+4z4xh2ZU4AAncSkB9Kx6YzDiJ87wcOcljjfrWBgOMs6
w1dqT5i8IS1wWZ4N5sIVZyTSayXS+wyHnKhB+CTgyfAnsVyIUlwe/ZSs+OdiyQ/L
XDJTY4a/KQzVlGYKnO9pn5wtUyHkEGa+d2CBSVjtd0gLhbardeBqanvupKQY2uiM
hFph5J5Gl4dhE7j9tf8OegDIW65H/W4AfUwZRHl6sENfTR/LbHQc/gcbrdY6xCpM
8wcAZNbPpvGM1GF40LmlRMxE6fODG786+9u1OpKID/9lTMEEmEIuxSApLqgvzvwD
I/+RLlLFOdR5naRhL1dYgW/sOfKlhLKbz9PnKDpkHV2LB2+mKz36B0ZBIzNvpia3
aRBTw+UezLzj6RumFBNZ1hpc24hwV+j4gzxybvLYIiLQ7sbekuR2gIe+u62h6Jy8
KIDkF2MfrVKq34n8bDhKYXta6C2Pb6JOo9ArgM+Sxe3ALM7G0+oZNV3iJoTrcNzF
6g4+ktPJ3b1YCDau8g9HaRGde/64H+LAJ1GhuzqnwCczrLZnXtysvtc6ZSNTxTDM
uoIrFZ2pdUExO7XWO3kVdgxpdicRFRtouvCYrCb8gfTGtqU3FiGInuZCHyRLy4FD
4frXetTPKBeQp5M+C4f7vRFyZ+uZQ/ymF+BDKWXF1F9JSgYRILN0FBP61R8ekM4y
JRzx2+rJuNMagMxRiDBBCdZiYPYrDTyIpVgX+Qxfsxd8xl3btaUh9lqSnbdROh3B
AXms2T8NflgZLt39AdJLfbyWM/kSbJgtDgTAGAiPiUwKq96OKW9qCNeNkNmZewPu
sViAlfpDjZB3WDtyOI/xxUySJ+60wTAPQUKlTGlEJxWJx9iIdV1OUd98DtBFLhPy
B9eg7OEEEw/1zAmNuWElNWzbWU8AnDkk+q3x7f3+WIPdaPR4i8et5TxPwwPSu/Jv
axORAihgZ0jviviK8oBoiXOSFe2qLS0McOFn59IUvmGRLArbjk5/5evdP96JOsHp
IkFLKDYexZ7O66Q7kHPe8Jw49ao7r5u/TDG39sQzrVfPgCbfyNJGzXmM4ErzrCc/
hIWSYSNEhFeQIalTPzyWryWamI1FZVgab/Dh9gnWAMTTT2mDvZOhcTXzE5C6UTN+
6EnjxwVD+3Op+918yGPghUj8K2AA7/UBgyq/1xnnNVC5QQNFc/GCpQiaaVwzOUcq
cqJkkLDq3rqtwlwjxO+cQRoe0TjRDe1YU/ukaVUtjYrt5M3PXt6H9a2gsOqdg3LB
eUTx9NA7cEdjmHzMA+8ttjVjqJZx8zef0CWKdFmYYlho5yGGf4cvD8xrCoYWKiL7
AewvsFtxsZx8NoXI2yQ9blozS5LZXiwOsP1Tuxvulk8nDIVYD8kQJLqrsD0CLyLT
4UQn86p37383N9NlhC9GQuhiKKaXcY/PZPUf+B0XYP/D6g4kkwxe2oGLMUitjXaX
UvWtgYKHKWODn64u11IXnpIaTig1Nl//sO1vvFAuzMAIQbWkQcEwJ6GTNLi77HUw
PB6JcD2meyf75uHOljCeStg1qPkf3kbgCxTfgYgXY/WA0bZLcnf6NZL1LD87/ZmA
BM3s3sfwQe43LhEmZ2liRjyc3cN86DVcpJAKrFdRz4MsSqCsHlr2lUAhGyTw6O3k
c4UwVLaSntfatRqOSt7mlTFrTt7aHiJAsDfqbT076EvDgX02mwW/c/4Y5+l/XbJj
ALyexZfxKVS3j0ezavAUwm7tYHnqOVWNkHTghoF1dlCxZEPqcLWRIgObWdCbAKNs
p5XVZLK6ggqnavu6YKCunfvOV7qsUYCNPgLpkik9gEsagwKrVXTrCmhqOblOUj4J
xWz0p+fo0CIm0gzm72TL92Y4bE/FjWJrkQzrbckOGzkXAQtITQYjRkF5iHC6tG9F
lgAy9MJg3IeYobYjwfplJm0U+D9hTK+2mrnNIBwWPfvAGWVj76KbHPf5+xQIT9rF
`protect END_PROTECTED
