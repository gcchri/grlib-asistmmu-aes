`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P2e5qagTsX2zS6EZoPQO1tW/f+P0RJgHRcBb5oSH588/lGYOtbmqWyYoixVmF0cW
EDhF8wnz55lzAIHZUgkCTz1Xghs4ERwhz005VHzUpy9s+YqU10Asjq8hhaAItIiX
Gwi7zmLiKGNeqhpIwEGLucK9UQu9fzmpwEzr/VXCKiaGvZHzKZ/OFACC3q4iKUYc
zllimUWjC/baWRdYaLVYU7CeDXc/mUG1ZSbvdK+hw/+IKsObESb+X1Rkw27Wx4J+
TAMx+zuse/wTJo3YCG2rmJqr/pum4+stiYL0r9rVrIE7m3U7YYILOW9PclfN63EF
o1pHtllCkQrH8aMWh+ru+v39iHEbOsSmiMx6oD3FeBXXBPpy0UNJguzJ+NvTGkiI
49BM5Whsn0Hy3mmIUu+gE+3a6wtjoFKz3YnetyWNzRS1r/LKL2AxTDsQWxMeLw9E
XCOe+QA1Roqby6X3Q+lFQ9Bgx2DTX+ZuxoXV/CYHRzOeCH3uM3S6wGfMS3JM4kb+
dmUyhuLm+oZbpohYMNE1m4m+5BEROkXy2bCqoV7vOMTDzroFs4k/xK0Vk+1cszpL
sLxmyQ3uCp1hYnWB757il7TYEAfwzRzTN7WlPKrMUV7WZWOsSlAT/kl4uk9PyZ4e
/rsNQCzOqpJewyw4WWmSJg27sry1sbCNKoO5f/A7giHeOUsjRuxhSElvWLLlFZJX
cwGCTgUGxbN23TY7sKKsfSu9dPeKVpD50/0+yExrzlZV1IDwLD0kToe3syJaBAlK
pgSZEEb6+9ZsSOjPbsNR1KOeZytv/Ksp3N+L8KEVobhf23IgxceAZcMHZNdle8Gg
BkcDEDUEwg0YQk6qNkEUyLFSTRdqVoV9L3VlN7uzRukna27oFri6N8xZPAHSdXmw
AF6FJCW2iBM5+3B1Vc5iMnThCZb9cKbevd5gjR9wgzMIAnVALQTpiX9JeRm5Tioa
91vmZETkyeMtwXOdXbtnZOM3h7jpq4DwSVe6EFGNk0KjUqad7WEUoOH3kGb7hDXr
ud0nhuDGHMUL2tvxZ/ju/3zuwFYGHxLwd1LAVLeeyZIWRlax27f89C+gWRYINdpA
yiRSWs3UjEgwl3YXFkNmA719SYAuRUy/XmQZ1QneWkssCNP+vdNq5R50g1Q5OAym
cHO01s+KypC0EjL6couJWLtEWHPSmN1AZhf4NyQTempMXtXVN8C8z+5YXLSZgth2
3iINa4e+WM09Gq8juGgqoS7DgfiAjCIrD0PrwvE1iOoe+RuUaaIUzEaDzNtUgpQ/
vNbWO+dBRigsrYuq3RwvS0bG/u/oyO2kotxBQtdCNNDHxzNJpCsxy2L+yL4ffBgM
bp5Fa1DWuCQxN1a6ly13ePIDb3EpMxVrNAf/b6n5zrXqSRrlXoZUfKYJoZjshPqO
CVO29zg5sHU223294AV6loXY5G6eq9K7O4sZv0p1NJxmssOF2DOOcuo12aXNN3ie
Mi1JveeM7AQFNCvI1JbNHMd6bjA/lOiMBc69JABS0PBi8DFEL5ix/syyMNsBNG4j
/6xFvNEi+RTo1QLyAGUuoHHPeli5dHiD2YOQxLopwePpMmSy1GllzDG/XAS4Hm6P
qUGtOtkI0V+nTyOvMAakgqdKFxD9SEQt1EMeFC8NiQatK1bfJBocTpOUw9oUxQp1
81U55dFibKWPAG9bP0TUPAY6+O7EdRa8Vf+MFZPCI6n2hKuOonp/NLAL2fflfK0S
SUDtPiAAzPk+nNuSiIJ0m4ZCfcweurnQPQn2faru2yOc6o9in1pssefl5kO2vfrO
WfoDMRw4Hy9tFQlMb3cA1U9U4OanIGnuEzqAOHNZrbOgUSarPBVKZ+J6z3EV8B4o
ezxYMNCpqB8tyZo4axi+YjdSV1WlIr2Lbpu6nRiG0bUGho/NNXul05YvzWPw8G0p
iY+BKUHkpkAE8E4a5b03+4VCiWdp61CX2ZJWy0P0nmWhTkY533T/WPbbequbz29B
Na6XWIUJnwQzrvxh4D3U/xxszzxX3TyD/boZvUoHeH+Z5W4QOy9FVsjrMDfTDVkC
HBfWOU1Q88TtHG1hMOrpJJMMJE4i4C85BrGFq3tZguSqZINGiOfIpm8N3zgtM6Md
moH2jws/HS+qtOL2zWO0XkFGkHQ7eCs6iA8K06Sd3uVXlXIaM3uG16TiYosf7J4n
ET3Z+B0UlFdH34WY+ooFwuJDnjH7Vjv7X1gu4LibLAZiEWsRVCFJmXoIOsfIhmJn
5Elr313plaaLLb3vLe5EzME/nO+Fm3DOdUbJGDMqQPneWWgNyTctwX3fHNWUmYaj
T9cycqUtLGhKCFvfqk5XKGB+FcAo7O5DJW63KCaqTxHsSJxFxqjIjqz3Hb3v/Kxy
D+/8eBa97AyOIFh0e/nmbtY3vuU9ck6MmJf6Vz1giu/5tlzI5HEouaxcCsbu+EZS
9kAHDpFOvc6q42uzH7brqwOjUhLHQFTK8EQn3Knm8GLouXB8Kr7SjqMaXCTpwl5L
4hCDDkz14akzDJgPxjgHlWjEM5hh7q+XHk54vXK2Usmi6U7pRs5WcenOSVLyLkfm
aZJ6VjAjk2ssYx6RngOsELtl8F2BnLxsnI5bwrxI5j4I4FyatG9ZUlEBGHv3Ry5u
AZpt5URWYvvB1tTuLyqmQinZLTfk/StL4JBfE3RQcu2ETZqWg/DhWp0nOmAjlA/S
M16lUUWCM89TrutX2RoIH430KcVfINOubB2AOY70BKM3SN3dBXLYZ3yXxZT/7y1y
RZ5cHVOPB14ABa9BHJ1MWPrmEItOJ4suGg/T6unZQbmbMXW9YQDPO7qBmiAQR0CK
OLT+OMpnsEeLoBSTzLLMCZ2uxEFkjxwIA4Ystf45cooBdgQ0dEWs3QcH4HBTO+VB
EQmxnptx5cTMUpR9cl/5+R0yGpzqrRAT1om64cKMwzZdRTDMyNXXJPhquNG619qG
i1+sCLXhHwND9w/VQnRx3Wtprw66jXRfrlVwGbBXxkOQ37obBbwuBBbqJ/dfdk2j
PiWF7qwcsCfQ7OPGPGxsegxUWmnEvvVf8yaFw6ZUv73Qkn8r6J0cSc7UT1ws+nzz
8eRQ/+vtn1ccAM6LKDN6Yqjm5yG2LOdJBjx5r+k8rG7cZ+SGnqRA/o3dWrHyxqI9
aIENQSpUMbzdhmuvVbqKY24KIsxEizb1mv6Ziw2zZTfLfzP/QdckFZ4pCn/1u/Xo
bZkVv1wA6e9h/P1CMky4Ebo/uTlSGdDF2DtJmvgJt9KoPat5UDVzoW0MDyO1TDPN
+TqX+To8l7p9dyCkN/ByrQooMToDnGaZcnPrUfSbwWo=
`protect END_PROTECTED
