`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xJRtzlINjxT0zAgujdxPkskW3Fo8If6VR0HGOp7iPXOo+xinm2/A0sQv49FDwRsX
OdnCW0OT6O9dPPy1adqtFVFd5ZQaDFkx/cspNEufoFjlvBE6lpcC61CY0nJEZD+9
OD7eFFOENhTHHk2aoQGncfBCFDashAcq2IIaY1phHytNwl4u5Ewbg6+dx+PdfUJf
/P77I8xekZJKWoElam4//wQnWRTZx47aMXK0QGK9gCTbyzDSERFdXXVSGw42JZ2p
X+TfwpSDPndBoaCqIFnGtTK8JH0cLa4/4uKJGXwhhXjMRH+jI2+i6OqJ+4tHs3VO
KHAV5yOJXR+gaorGrtwTJu54lmI55+f0uFaqSOKtf03vOeez+6AGQHsxI/O/iL0u
hDn6Jc1Pw8MbbMNjQjVBRA/pY7/dMZif5Xfp/+nkjsUIZW+sBY/qsuY165PpK3SH
TxsvLHBV+lzdiEmDD/2DzPP2NYc2yTyLHt94TLmJajfnqVne9XQs/aPqUixsV4KL
yFo3DSNalMiizf8Hi0Gnhg==
`protect END_PROTECTED
