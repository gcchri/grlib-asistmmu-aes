`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nGJlXsOxgl2yFN0uPWZgJAcUvF0Jvr2AgwYgRo1jYhEU472beDFohKnwnllLDKWA
hulnj9Bl6fnYf7E83KrLMECBJdrOvY2M4HJ+aHUFz0todIeem3FD47YvCxM0RFm6
Xj2e/Vch2mU9xtQsiwpcJLTXCQ45ltlT7UMSsE9h2ocpp+Gzw0fQDVoVFlvGk24k
nIDzNmPRQyQ097CsGnCqTcczJLZkebhZAgJoHcGmx91X2CQOhaSW/dGsjPHK5HDE
azHKdUF8y2hff6e/aAGQhTtUx96h1PRqB0iGAEnTMI8/K35wQCUX/TZdbQHEQsVA
hiVwv3kpAEZcRgbDP/KZwRYmdb78LQK3j6ta6Mb/iVhBW2cbHNOYj11Qj0Fhjz2B
jJ4hgQT2jitoUdlgMbe6LfmZ8kwqa6Hu9d1MaASTSBdXXSEVTmDsTM+4kYy3nGoB
zxudVteMc0iUiGZuwX13i3uT4iVSbFGb/w+WiDXcLs2JCkPU3Bet1tiAL+mCiGqJ
HlV0nP/p/wo1bJuS34aa7svryW4AhnLpcAyT7iFgoPU731MRHDcF4b04e26G/sMw
XpZD7XZ/rILLsbob87YeqdqPDhpEh9YkJ4AmntoiCFSyT+W5cBdta0cJI8vPws2f
0oPP25vQBVQD1QPejApIn1dfR5YGMOz+AMI0GSp3lFWVmus05wNQe9KcU4kz6nQN
ws8Or1arWHQ8rDuEY3Dg3/f271VOedhJ2lQW1J4LE10tvUp+sdr8FZ5WxhuKwiyr
U+7HBnbevZv1aCawyvQMFFmfpjb0ZH2ooPpoy7OPsSq7pkfvVG/0tf1s4J5ZSqyz
R0TJY/cDsO7vUEtxb1vWJvBHV1drWjB4gPU56ul2p2xQppLspx14renstJ1GIvGh
S9m4Q6pB7gziEzAtQWFWbw==
`protect END_PROTECTED
