`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wr9kbseFYaW+zUXsMMQgwHKaHY0x/BHoWmhEby0h8cuKIO3xwXquETzjuwjqLJ1U
AkNnsAbvvDFPU5Yhln0sv5ub3vhCmZnD+aQXfWZjp/YjTp5PIiEGU27RsjpqXXWY
CDhqPbMyc9VEYeuL1LyXGIugMSBKFJLoOPLCEYKYbUVAh8t7PoVNHKs86Gkdrgyg
tddAW1jcnGPunl9uHQ6sAdy1QOM0dEdO48CAebP9I78ABz7G0E0JtBVac7T7zG+d
TnI95RUgwtEEzjzXJwSI6r6StqAyk+KDKnCcFgnzpY5AaZelq/S4PcuxuIzDjXd7
M9TZqZTf28R5fPQSd/6aHJ8pYp/Gtw8Pf3veCBBMrcuKmK6UnHSKbE9tCvkxQP3I
IjCXKCEOTdb03N2lWsslqv5gXW8MMeZsyDlGFEWzXKE3htftxs0cs+vNDvhq7Lox
kauBxjajH8stTvvWB1Us23LvquKlYBybdJoidoIVuCP0yK0yRUMxiDUQ493sgF4C
nVA3VnU8zV+rQHN+VaMon8X5AlcVmkaOEBOvilhzqZqcOF9sU2MYjA/lPoulIyOv
zsbwUAFDDrzf8g+R0h+K8PljOui4kjBv1UafRkTJ/F0u+Q18/4pIfRVXPSuYkVre
op74jG6BlnPocpgmYr6UoA==
`protect END_PROTECTED
