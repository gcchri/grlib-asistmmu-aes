`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vZOvV246oPAgTKVvF6v1vakd/abM1YQQHNlzV1Hs/YIGR4Vqg+Wvn4n8t2FCrip1
+yBIENKfH10UBBGoiIsswRjmUPHay4JknjCZdERpxmIMVoH7gSHUMmdlHU1PvftB
evhYxrvQg/pfxPcObw8XTj28o1rk8dSMi/pKFLoL/VnySefMf7juVFF4cushuAEL
m4c6ba+2VJHlczSKrQFlV8hF/Uw4WT+IsvUdAfDkFjXKbNeiOQA/wt9jRSdUur6+
MdQf8Jp8HDEYrY8q8+nF5iGgD9xmKKQx+zjdrRVnlpQLzpLman/WmZv2Um+cqtRB
fhVUs5je5YAsed/4j8MrWw==
`protect END_PROTECTED
