`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qt5EldVVkyMYkngLVDNP6HYdKOvUi386wx/e8jCE9DEeZMJqsXLLMySTmsWmjxTF
IS1gwlMNyqAcXCnN7+Vrn3JYaOOUNvcEdKMeQsu0bJyFLbpSyviMAmZ5MKGh762I
lh5iUY8TBBKwWMCeTQ68g/WGcNR75S7FtpjnG2lHa98ficKwEae3GNWJp65BNQTY
J7MH3hrJaH/fKJuJzUrG/YrRN5rnKlyTzFAjUqEHD29TfN0bQ1Xt/EZr2VQOqBoB
jpQeYPN8u7d8izHsKC0GZ5xkjdtGkoKOLi9+xZ3Cas764z/RJac5E6OMg8YAoK9s
xWXq3sJWgifxe6xJivQsX7wfn3pAO64M/lRi2lYSC2ISiFnkzIzVGGFPa5JnzRF6
qRcp66G05XuGKUQaP4JkSSRxZUoYSaCmyrgWinYBQAiQ+pqr15qK9j3j8Wgkg9PZ
yMcZeOeIUhbbrBo5d9KnGKcKLcATeueVefpfWRyITMH+cZb48bnPcTMN4KNFFH8B
zJz/XWTtTaZqi8ypHJJqcJ7OzYSRlPId5YmBMazzRpj7VXghi5naR6tRoKLJaIvn
XILTPrewaUJ6AHztgkb6JHnZH59DngKioH3NX27zP2/qmlP+grtwP6mXqZWPQ9hD
+teXCJwOYPQP+thViywHnEbkKRsRWD95AWqvDtTf+D8dCTk+TtvyN9mHCO8K/sAx
NUFGep4TQ2q0gRRcLUkbPYkYNd6jDZ/FCnetkjkNabtcTlz9Km9d+uP43dlCi8ay
ruxqXDiplyDEMp3cju1+iYCX0uGPcXe28pEKNqFpTpq9fDTWu5a+V3CAhOq8GOMV
ulSK9DGcvy+p+DHY+vJPS7o5T5W77pCP5htrQK4+BoORU1zWXJy3n0yGrRpSlHPA
njk9LfMkihC+xLF0fOT6r7Cc8SYVbYmsyo4NaxPUY50ysaK999FHyw09xjxhGSLc
Xz4r0KMHu8zoINGbk6Uj5QejBVhPd+bwmrjaEeILPQz/h5XXIr3bU9QJxHOu+Mr0
K7zb3EY9H4J4jaiAlIHhOgRxNy5ASOGmzTmQoJYnll9Nt1z7qYUvEFQSayug81nP
nIZlNg2SQdLuznxLSUQv/bj0kQ2YK1qOUXPOBg7Zu2gE0keYM8x7ehHbrj9Uy4co
H+WPhGoQ8wt8mwbwDrFG1ISYgwULARUPFQeotSUD2+y6TaNW7zsnWM9Os7GXYO8l
09uA7SIfaLL1GPH4znT5PhsW5hCgP8J1iNOiDAwxqDrnwOEp9Voe1lcY9bmd45wT
YFum2xgayyjalt+JOZSG6ooiklPldWhbegb5CTpKa8nx9ZvFyEBb6gLMxuQExoPL
1Yfg179eJ6Tf2RWrd3YxvhXi1FR+DqpK/QJOZllW4YhIljMuHOa1JTKd7Am6jIfX
Nj4/1FvDUhIqcynNAavpQTueTodVMyTJxuY2trqBp2ruBPMliqFc3+GvU729DiFo
2KX7G9b8ok4Xoj7CBTNbbVw/gp4s4FwZExFV+l1OhsE=
`protect END_PROTECTED
