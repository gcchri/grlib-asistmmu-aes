`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xYu2m4Wt70F0cfY/ZEyVA5jKG1DdupyETHMR66lCsyYR+fW2QUB7dqK+BE/XVrOq
6Sdhu9fFHBQfJEL+4ry60dJTm5aKsR8HhT4LL7fryKlamgQnLw5tBIEHdWGOO/nj
nXfBNWPrDtmN6c1uGcKBieZHen3tmsqttdtrZl09H8egW9nPwng2Q62elIDHAlSI
PUZOca9S422cLzlsyon3+FRGTPB0eT0fvwgyEHz9XwiPnjCkuIMMQOwqAwRv7osz
TwZ/5bssxSnmsddTZiGd5YsBr5w8pgpi+kKXKTDgpq58DnTRe6KRely9ci/RiK0a
1kzQl+EeRHj+WaF2f2rNj1ZSvPUPR2d22U+wPqwciATINWN0GcUFbZX2xBU0h4fN
1bgsbSeIjq/FiZ23JLJfF+tDB1kCIVuxYiZQjTAW2ddgdsZQjiJSq4oQS0doQvIi
EqdDAoBFYJJMpmEXeajlLtUGOQsrmCrBrAKRM3qWCs+IuoqOz/S8gMYoHHcwVqDm
a185d41ODC243aCSKbI0bgAECKKBYywHmtyrgjPLKOQZTJVEPuJ3+VQlRj//tnmE
Aga0y1+7PxOa/C/sXtg3j+e691dIqjSvxLlrgT4nE8yC7BMYj6IM2zYiEibsRgLv
S46z3i9UKE5THy6R3BUi6+ARqxv/g4bOBzq5iUZ/qvFEGq5MTGs3BiTBkMqCgNLT
3vmFJfBhAwJHzqPfMFETVOF1HCkH7XIlysdxfj0eYY5YPT560KomnA+J+evx/4Ug
zKXvtCcU5izNs2PFMiDRw1X15jYqLb3ccPZnHH5GyhzPKeIvmuDuWXK1MZ2+jThK
+F6ZTG/5sTcLTkytTVVQ8m+LeYuKsQfe6SgIeQWOkEAv99i0UxegQLl5/8XtgBHx
1nZzo32T+aTDUUPgXRfAUY2p+r3y2exj77MRVSfPRCfNR4qRfUlWrU4v5IJq1g5B
vLWwVzNbbWKPOFjmvkMFFZpKWeY8d9h16Ka+CYAC4p1Fne1UP9Fv5X8LKWsdz0gF
qwtgS4kFErqJ0TJifN0HK1k3D5m+MshoKV0oGHn7Kp6zjzDONwX0zxvaEt+MlqAa
UqdfP42TAyPdc4yBVeBwGg+3Xzjd42frKJMlwUWu826QIvMdhlFv+yhtwUuJazQX
zKXacz97w/60nNRG6/xpxjGmwbl+TOO0xPsnEUyhuvwHmiSqm7dAwhdEDfbPL0cq
ninUr0sfgct1Ij+oqByE36mfUdJ65JltmqfRjmjEXEc7xzuGGiksrRXRsTRyfnYb
mAO9o4ZcA2vFElQNYZuGYw==
`protect END_PROTECTED
