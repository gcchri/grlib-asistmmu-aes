`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uzpmKVRhpNarll9xxW+1B8JGdF5LALxyIDnrnge2Cr1bG/d2iIL8z5b8z7y5bmxQ
1KW/I1aOHB86e55x5rhqbMx5Grbe0iVR9ZSxIPjxiSyM/wun2RJCAn0JBh9AUMA/
ZxlxxPWij99VLidybtV0jCIz9clEjjqs//5UmxJ/5TVCGY8NMbIviQgNiUUZybL5
9rqvvLd0tz7tIQadSA2OOZMT0v/0H7/TMFuDQPzwMzeygFFpXqY6IhLBZXi7OOHI
KJn2xm9xqEL4riYu48XjhNl+srBAJ04BwG0hONj9YrpcXHOuT+VEwUGpibMDF2k5
Znvwj+/FqNSPWtdJK/xub7bwFiIjSHDB0ylUBAZJQFPyWv3tgmiOTRgjWNW98bXo
hjXYP3pAbfVMiIi7o7ToUOwuKSe7b5/DcX/2m3UxFgGCdW0+Hn3q9oPOr/MsxIGV
lFWVUr5Ak5oTTrOW1VqR70IYVS4D3q441z8t7LypptE19U8zJE4YRd/d1dQ0w1Qe
uBbmAGZK5Y9P3ufW/oBxf9+ovYmOo3LMdgEySqt7u0q9SSeaMFLmkyqUNM7rXzU8
c9t5qaT/MwTrRzdyc4h02Q4sYFM6M+TczB9RBDmI50tLrxOYb67clQKJdy/bfVZs
pPid2xFIaFG6OL8Be7j78oprwwSJwdGdY7a1vPH3brlfNJixflI3lm0/nL2cDeL9
eNWH/nIsJFRJtFpJWOWgyMiBJ5tNUuMMvL31krH/VZ2U/dDB82eqNDNfzN+gKx2E
K6N/TXk1C0B01KkDnrpVXKrZ5b0TwBxV/VkqHk6kU3yKWhskxcE40CMHvnqgvpQX
RGQzhmQ0x/9lgtmHogM48IP+Tsk0OMMmJPWpb1pubLewuZX6/JUKUb6IKv+QOY7r
LXs9McZ/RXWdFGneuWSRGssMgHqNzGSRKqTJALHLMI1C98bvegDvccPLTaRGW9gK
pj8Xmtfma0dMIv4anzJz557ojyg8+FJoGH9gtBfD+3iH254PbxqY44MLv99m8VY5
zLig/0dAqNdHBGWFB0O2T8acB7pDuNV8wIBMTpoVfZfVN6qmz2ra+pSBF1DvmCq3
NIwjTuOB3H8kvVtIGeUbecOxBdBhYD6tUZi7vZ/j0TnT9AUm+OBkrFVaKTaC41BN
FfKr9d+AKdnr/TExDjj0CwfGZkJlDIhXIWi6WQUxlUb2VArij9Ijke3pKQ+ww9Pb
9/9RR/bA9HKVUl5Wis4lpXYrRrcfX700rt8To6Z+sAjQpRDFVyxTUGAJxCnd3tFD
gWGGENzmBk238pHwonHdVRLsan2YSCHSr6KgiNJwUjitQiWdsk3gvTOMfwNAOFl4
tq2R7Cg81CiA1Tj9f3P7WgvZwYps5cbfoKGJ/Loktak1SlGgyAApDbkPpUp/1h7L
FF24jVGdb273hnSlOMBTpKEKiLIlQFztkdNx2QblgACa2ieKRI6jhqB/M7bQmf32
JJEN6EAWGb06J/mPD8wzkuxLH0v4OVtQBDzlIYjzRz0R7FgcUaiq8K/FxgE7ZFNn
ElbFl0zwbxg2ne9UeFNyDDKhuoCqYyAtmnKUZQ4/876rNB7jyKIHzudGWpIYxo9h
dH9B5VcuWyCS5Yz98gqLkf4ksrGdsLAqUde2fY/g8R837xoAT63V8mYONndJI9RD
npIft4oZDsqKlc4M4q0XwxdLleVkB10Z6J3kF51WaE1GT6ey9wtErDNhvDkYr6Zn
mrNrZDdwvfO11d0V8UnPsu1EH/3msXzFzC+k38R+QZODbYnDk9giQ874s2cwrtM0
YSh4hzb7mA4SGBQXoUigVjt5ZIOGlaqTbynrks104t81eDTQRqjpJAoLZuoOqMYg
BEEKl0fLM+6iO0ye3bdRziZQSfC1co1ddH9OWY2rdryN9j4YT9mt8rl0W75VxP+c
kTTh0pa8nK6cISMwh86iZ2EofbtHXmgCnsxGvb6IjJEzWBKV/0tNFSf9sXBt3nzW
4F34QeIb0Pc/UjKJzVjUSJcjUGDcXAJ7QPfrLH0hi3D8bhU/YzeRijLc/WHyUoI8
wEyMbenW64ZtX0GLwdlHn2moR9lSUm3/Zj1ADKmZvGEFJxEL194/x1J60W1Me7fv
OAjc7tfo89GISZBrtQ16qdLROQXHgxFS/gl+GEyvf1irnUidGzWqyAKC9c7rfger
pP/Wc/rHst4/+IIEyHGnETbfRGdddCM1V/3rj4cTw3BzKjaFmEKKgMDvkGk4nHFL
8C7gNi4YXi0oy7RMvO7/kZ0dekWEtNP+lfBPqJ+VBk4OHswXRv//KGjKjVCTUFXU
NN+jOnriLVWgg2oxDzmVhHxilmfRFnbvIOJuAzNpPzNPGS3ZzNtag7fnzPi7JbZo
WE+LEIMpqPxUK4fkcGAziXvSl17ed9Tn939DzWn+Hp04VkD1fi8vu7rjDVUzjQOU
dvChITBT4NnKL6ylBJuNqJugkW8G3nsaiXJDOQk0J5JKX0dTN61MeXYOjUyYEoI5
xRi/wyLIDZFhwO8PHLv+5mKNN9XALSuXxP5cjJvlTuJ2147amstnzVYH7r1JweRe
2laonsQzxwrPkpXzAR+nT4SHhyipy8ELxv1/EsZ0gQKIjKQRizn0PyoYycGUfzFA
1/8tWscziRTRiGEQ4R5DARKX9MN17DSy6bZEoJBEHST6S2SASst2aBwvNbH3jfdN
5Zfjkt5EMe6/VTQKsItmGcWciAmDg3kThMuIxa9a4bjGlVR+LLumvFdhF2clWTxp
q+OnWK8a2V9M8i8WSLXNCRY47DxSm1mbatdPQ4zEalFpTai0Er5dVrSMxoYzCmRU
a16clUc/coBkza6pcOE565QWgEX7T7HEpyFK3Mw16Z2VjSRceHYtDGmrYsbVN7FP
U/RxK94fKS/bnFnewm9S/aWtqOtq8NF305JVnO5ua9+OZTfMYlHiWu4BQiExyr0B
1/F1q0li0ueMPv0JdEVMyVmsf+buyBpEOV/32ATvUO3AfRTYr9dODxs86tFEnxlW
IOuwqVP3jmCwRHq7cer29BlKVA/jlvnPdTi41kFJfxWqdd5iGiAP1tliwseYFe3H
8IjHYRlU/53HxL6QDDtN4CKqik6Fwnye6bNQl4dL6/sykmf6yUofQKTmZEQHYqX0
4OO+xOxxJu0U+y6pIIXMYhKwD+G9SBkFFuw2Jn6D59gTVZPXcvht1jrnMadwrqrU
LyLVbWWrPl0CtGXKVl88AVTcWpzJT+kYvAWE/MKftLzUSD7qg89R0d50z4hx0M7J
3kUUKXcqphnIWLw/Y6UEHO71+laM8sXJjRkVqEOSIOVj512CyKjE9q3vEhyFk0vu
XSAH8ZRn0n4nhZbUGfthTkPlDW++TICPm/BF6B3V+mUY9lE65fLM+ouiFR5lt4JH
2sVQzbQF1AC6/vK3NwBmuEZOoQ/gWoNFhVZRw/VKMOVfG13kncmdsnmqbv1vpK/G
jYAGt93eqhReaHYZ2YrPvdjxVc+/KPRKq736OOl53HozqlgVQIeIpjB3dUq0GOG0
+52XPTdvavXpL1gnffdXrA==
`protect END_PROTECTED
