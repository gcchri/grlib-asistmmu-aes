`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3RwPutOLwvC2mKBG1rFaPTiEzq7JCgguZYowHL9p69AidRghpPbtYUHOUYwmQgPX
EdLTTFBwuhucsIX1pr/mXKnI1rRC3Cz77Ejt850AM+KiwN+QKybJ/nECl3Wp4u68
Vw1oA8yUMPrTmYkshY47WqZFcMG2A6ldqpBOhy84K6UBzGpieHIadXwjCCss59mE
863Bh5VDaQETxDCetQe+zulbqddZ4VWxy6JtI54IHpBbFWkmqPTjXeGdp0o2KKM5
ixQEjD6qy7/CVU3ZY0POIHUfRXE1ggnIp+VdvuNnqIJxfIZlFs1CnPhR7PY4yBaz
`protect END_PROTECTED
