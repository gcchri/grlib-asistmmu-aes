`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xHYI2wu9SuUIxpATIdQj5Kph9bAC+YJS+/goIvBcPPQxfEL8BPxUK6s9OjrByTio
k9RkyVG6pEygo0FIy3if8oxbGbTUBfZonpkFPFoLoow1UwZ/IiMYieXLUXMtFBmV
VJX2f/I7VxNeq+rx/aa3BgZqT5ECunc59DTYT5W8I3wA0ebSalRCLn6bKxCh0/yh
9HFMIFMdqM6nKMc9zE9JMDg8VJJ8DT1Cm+vHZNthHnpTPGhz7HYWsBootUvhvm9K
jVRjTey5QFWvz95eEdxdQmUZ579tPR/h0TSBaaXibXKrIt1QHMEJkWNvhCaaHdOq
FDunCOE9iUZdRw5NjbQPGSaiZsGCUqMmvMtFPtDoTtGsWZuTtwy+G5c/EQK1PLcU
DBGnQvSKo7Mqa7Q+MXVP00Zkgd51SgTTCetWBcCDa/ySLKCQljydPSfigdAag1vX
a/8s3ggEY1km662EI1n8XjVAHyiMldgubzRlNp8joYK6TErMZ5/tGibBrK54Dp12
MbrelTQIVvwLnxeXF5fZN8ZEZd9EnG09WlL+7aU86b9WJlca9c2n+lY+Va2VK0wD
EO9Bmrab7OmeLyN7icp/ZByfjbX3hYOwR6p7VOLsBaqKy3vjVMPnBcpGdjJF5Zo8
Fmpw83aHcr9WQZKJaYHql3Zn8/LJ0tm6U0IEDya6HXTjtHBFm2JQ4mPlvteSNkJ2
fV8Js3okB6lUfzPumOnFEU5FRQeJ/W9r5C3GzuaZzEpLcFJkhFp4j9o4CVcJbAoW
4XNTrSAWBRre1PHapyYgKY2APMtSwqfFjVUupuLB18v2BrsFiZFoWOewfozU5goI
JXJPmK1Z38OzRI9GHDxUWw==
`protect END_PROTECTED
