`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zt14KlB8Opx9leFzzvPZZ4GjB/Ejg62iGg7cWAnPBmAkpmTe2m7vOnZLAuDisInM
po0lZvu+MFOT9xhghp8S/o4lf53S+0LV/pq0tb2W+x/dvHFwJ7nh+LgOqlWaXS4A
GAGdKa3h5QzCeWndoM1h4iE8iqaowHCnE1sc9mFpqCRMGHjcZWR/YgfGOBeZBp7X
F/2SP+EH0kZNYhWBDo1Me0FKcXLUFjBnoXVb/wO1DSvxIFwWHqwA50EJ0pvmMH+b
3gWrehW54dFE13q7fVlYu5it7qmqMufMimOyrlV7otgZ1kIXKICnu+fZYH5fBd5C
c32/Ujr81PgOMT3cFe3IMXXw/ysPiWNBCe72zr+re+fjHcA6hsVnbWDBM31Ns7G1
BMVW919u+76bWQf8JKklAWRF2zVa26ugarJu0sqYK/MAgTyX9SEIJdNxMLOW5UAL
G4Vp+3JheGIqhpzOJDJSFlKYQRYFVJp0RENzx1d0ViBwhR9+CsJTZFaU+3Qwwsuy
UMKqrwDibO1IE8+1zJVkGH1k7ihN/5g5NcuqwYR8oPIqwe5Txs5BEcczHxofztyI
Ny+LFfRS53nq9h5OEAMpabe2eWKzXi5YjsfTT6a7uMXroZT0tg5s6eDg5m+3NtS/
KsU7AA69zF7O+Ln3gY5mEMFB57M/QXnC12uSSKt1CKW4Kl4SDAhQmgYPhrOMeUzv
j8+DweNQtC36X2a86uL0x85Er6KKSEkNjJGSva7pKW7TpWGjOSt2BewYDW5nLRdY
5LpDNx0hKYFUWnZzbPFaqrK1K+rpjXRt5x3UAMrRGH0=
`protect END_PROTECTED
