`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4LqOlsGFQgsW4NLrkZhe1xtxEG4BaHSmGphQ2FscKjZgX5hC6ajPTQTlt/SOww6l
akSVoA4ohNZrUfkT/r4FQOlopRI1o5siZd89eo5UeA4nIk9OyQnLMCtXdhESEB/B
HoW1VPhKCPvMtBAocp99/02k/zLsLnJX54WvyYQft/d3Mps/y8R8vHvkgD4Z+klT
FAKQn0WjRHuCKmDxwnb7aG6n22vsLcPHz47AXC+Rb5AsbGae2TFkQJetNz7CmoAR
GbojYj9muvSp8HcRVxeugjd8srkjRTcVhH+rNzOipIVe40hyLioSwM95dMO2FVsL
vwfJNuN5+4TQLC4qHvm/rrGDOweD5n8IXlqZg8UV203sDA2bl+kWuth5nCGLKM+k
7RvpDY9PqCCniXGOi3hxp/Tf8KsrQp9VuM6G9VwvgURUUMD0OJHJe8TLCUn0nndK
1HY+SZ9sgf7na9RkMzZtUyave8uQXPijhxZZDYo6KMA5HQn3DPfJ4ipiWLkpxc7T
LDRzhc0BATa0MpbLjXl84DQNSLq4e6Yle48Wz+2dUhGs1bQruwES4ETqu0vLumB0
vNZOw7q921nU5ipKzZTqiSB2gsV+IBULqB4ZaUoqkusOv0Lq30+JsU+mdFZYc4Sz
u0oVFK65hdi0WjL/oP/3Mx4Hi4pNmXgLTZS2AU7oJUdftP5Yf5jr0bbml/2hOE5R
B+658sq8BCL6JeH2tQ/s2Q==
`protect END_PROTECTED
