`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p0YN2XFyBmMIh6fDfxxa6Rl96sfi8m8Cc4f/R9AXl558K+dazppC6yTBIC9ZZSj+
wx71PKlpJI1f5D1IydCS0T5w78N+IVmJqpqpBnjv8oXsrTtLSTeFV3+1jXw1LQta
oNyOyrquSmDYuuB/zVJSQASQCxack1oq7OIl0CTsB8jYRtiVKtoWekgHto8efD+x
dgAsnq4ADhzf4NLD0Ei+vL/PH43Ndna04mpzeChT8wwzQbYcvn25kwQlvTH7/2mX
ybk7RohxNk66BbFE2QOVxdOs0EG6w53Win4Vc9l1kBmF12cK5PnPwy35FZ9ipHYU
eIrT4wFdsRzdYQL4kx/PDwXuqWHPNHvUaehy5w7bk+/b2kne05wi/GQoprHEoBtz
mK/9LM4Vc1S89NT0Kf3N6hXCoOqTH7GV3cixyueCNz27DjhzZSjM77mUsb10jQ5Z
gbP4JlASQJ0YaLZo3LXMLSuR1R7y+wrTpLIgp1ct5pwCFZlzkn8uUaPMdOBpacPV
3fxJ57DeJvI0fsAdRlJILf5OlUhy90phA8B5IbTfe1RjsQdHUxtAJIh1KZnIpZar
ARFXmut+0H5O2G9nDDTr2x6O5Pe1xrtxK3mz/C9oGf8Lb4DCz7hlXHlHhDQtGwzO
jmCnksT/c/u6lSOlWodcdw==
`protect END_PROTECTED
