`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kqeaN2gZH0DUy/QeHHuWpkydrKYBUUvsWReHN+j1x8ZgAtqkA5/ewcuILJj45TI/
WmeFwXRstUU72tKwg8YjSL2z68A1n3Mmp3mgDXDwP+loJ0o/pJHtGKmzlwNGsALh
jMfWHF5krhQG/StAZ7m9tK9vNlKQoM7YsKPij4Y+294hUxNemeiXv6MNEyo3CVPa
yWOhhN4/zXJKCBA1Pv7r4KCsJ3TyfvtRyO8UEkp+sMZGIQqxFvlBvfjNNCFlCh/t
VvtF9Rkit3CLpcSFTVWWFXoqTX+Y13FN0ucHvqnBaz4/TURf/m4jhZiYJVUDm8lg
J4OSOUXsEHV9OFDzaOiz8BV+9DEDLgRDlfWm1l4NGMj9oYb8QBeCoAZzf4mZ5hBp
E1ZXaf8mluqlesWhI9MT6/DvUbA9fJUztfxAbRvftsQ/vNDwy0m8wViPzW7QHfTO
IbPdbuoZGU32uQ/jGrJ2zyvYsuDZsVMZdY92DdDXrcb4h5D0b4aqaBjFWM/OPTau
I5swSAt/VG1Cc0fqwgkWSWHrm+P0721d9ohtvwlsrIZ1TYThYn7bBdHq0O5Kd5so
RS9/6BTWSlsWZvNptwMpq8PqLF/mIzFhE3LFnnElS1k=
`protect END_PROTECTED
