`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lm8/PQSOb9NE/LsOfcCqwY9KCgS1AUjUNOv4BOd6pnVubtqz+GafWwlu3v4XpPnb
hCrieA9zobn+mv2b4aBL9RGKSXL8gp7UdQYxL8F2tWE19Zwqii1sd0UGW1/6hDYV
KLkiGew2kTsE+ZKs0NIYZV7LM5ht6y/qInpxaQNNfDvkvIlvfL/Gl+JzlNj8Ip8T
3KWPxMJPixLMkybFMQIvqMEal32bei9TatoQRCp8O/87xVloF/wIQkunhGrLBne9
b19FMTMDZnqO1KQH5bmmV7O7A2uimxqKphgRLsY4PDQPeZHGNasW/p2dO3nUYB7q
SQGz68bMCqgeXGRuS3VNqxp/Gu3OFd46qMiDpWTQcJZIc8azcV4Wus1x10vxdSB/
vLSwhavxcUwN7Yli+S4u1+FBWTRntsIbQgU3Jhge2kfKd21eAt0dB/0QTX9+PBLV
Cgpc/uP37FDA/HaRBz21woBQ/PgqAprROHksIM60mvWzxuCRCcWqyAnbtsGv1pS4
KAhNHiCuVvVkGO3TcBtPAfs7KDJahtDti+pirUPsgpobV228QjKOyBkPJqhIkE/s
oybV4rdhvu+UrIgVxrxu1Vy1gfajA7YzYErh9g08pG7rheBmXUyC81KvaWTIRE8x
C/AbvnqzwcUUwSlVC7EZACzo0tEKO4Bsdk+kzT52U/kyAv1ndPxOk21+3jyZiSZk
t9sM2r/vwVN7q9eGJRUxauzcmmvETEDAYZcFTIHnwm/NB2aeTTQ9pTAcMxFdwR37
sDh6Z0VSKZda5MdfVZ0Hb8DHErvCOhc6Sj2shPhW51dKBwajJTSoJE/3BnQSEuQP
DwB0p8lJBhCaYW/hTZIcKZmY7IAmuSwd8lEZGXA3u3MIYMLu0WP/igCANZq+RSTx
RV4tnhf/J2QCvkaKiuaRAbWTRAmgurHEVbCq8IDYqGpOJcBmIfg+4a0SHO5zIdnD
ZXIQO42p5crAldKve9L7GF0ewv0Cl3cmWwTZrK0ch0oxjaZyAoQBIWFbeWNwO1Sq
aR+B34Ffc8ewfS/AJKWPHyxkF/unwsRb0tvOgqAnS/5cTlqOV0nIkvrkDywmY+9z
`protect END_PROTECTED
