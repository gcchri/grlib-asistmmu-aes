`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BzHuO+o+DDPBykPe+q1IghRn16eNr/nzfkdqhzPBJKPXFSGKhdmPfhBM9fvVkcOE
Gr0DlUlo+4okl8Ej+FTEiqDppKMxfof3yn0gH10qmchajZ0xiDf8mgea6bCxruQ4
2ai15MTAjox3b0kODoi+oLF8TjRNjGUNStC4ahn8fuObUa6Rh1hHKsaitFF7pf6p
DS7fywSo0FcDnN4iew0me8DqiR4vqVKSppKuzr3Ng3473/wXWuYDsBAgHpmxzeqj
20Q+PEi6BAWhF6bW1fth4z/vqsdZpbS077XQI7IYT4zqo6LkLzaJwy7vJX4WxbzT
H2g6uqFxZ96HnaYdvzfvB14LmJl7ShMiQR8TqzFEejokfSsxXFfIuahoMfbIwpJS
v/5ntyVj3zsd1vHVtExFoZX+St4Mnorvb7/VuNRUEnMTuHgboF28vvqgl8Rkpgru
gV6wd6ZzOza25NhVPwK3Q0GbPAcV0IbLW8qAtOnMApRalsyXqP9i//GGY4rStYv/
VXdAF4qoc467HPnV9X1ZF38UTqFjGrKDCuhrnC2BzB8zDcKfIVidrAW2jbaXoS1Y
RBvoycz+m2G8bq2MlxlMzEfMmuvImPCMVlrKYxBgGz6MezWsaqNJiHTp+zARdtiv
t0DwQlttEExawhqn654rHr2j4YB36KEuz58qScczlOiv2r4Fp/aeMzhggdlYTFwv
HxtkprKc4f5k3SNyLXw+5Kn4FDwEokDnc5/G7Pq/W09yseCJG3AZctw3VbrU2AMb
fRLtcQ4wo3bth28drFr0w5ZphjX4ie+BNbod2nqgAJcANSeNVVC43qshosvUpqzU
K2rpfrLefeaaaiLy6GHIiMqO7n/8WTXRr3YxnuCRtW3gIN4KWwQnWtsnAIz77mvi
ovxbQn4jYav6bNwp/YWdhkKEHdJz9pzPhsqTFutL9O6xirbBI+7hOr6AhacyqZfZ
7EiSBqOKPHrub4ywNfBqjeElo1JMhrc8kx05szNcjxFSq93o8LPrdBw/rWdNzzq4
S+nIcp3+7+hc3WaZQbmf7iZCgzjRmtOLY+Na+QmPAKnWFkZX2PABj4VL5vWsY2vn
aaVl8viwxUT+QmipH9f++OQisfi+gcN745mk48ZOj9xXYVUBmWB9FjKJ1MjI3Fi2
nZtFCNWfwg0xLsnJ1VYVlvgs5wpPj0JOE2ZnqpEeT4xR38KXNXMUK4RfOd+vklxa
IhKcSYJe0fy5yLAg1rBfZlgBDMRlu01Wusc9NK7RrJDbK+Az518GGAD7zsbjUbeT
1keerfDvtrXqVpi5/R0dnkx3cKTdTjKFH33xTJMHxweDLMG8+Lk0K7x1MO2EBiyr
083hUIvUSQyX3fUBYeM0XkBvkFWi6yGI32wbiiH/4hMlGm6k+259+83ORY5ZOLKi
7KP+tZS2/GNWnixdG8Omz7QO+2l30i2lOH5A6IlZOWp43Zrcr4hAXbkScmIBxEgy
IRfoDC43bEW9JzGrRWX3wxogiDnae6eCHbyR8ZL6deISnBkIrgntHBetOPHFRbmn
jr5eTttfz2CPYD1kZ2O8ehLW8Q3whXResCPNC/iFyfEUzwgFmfrBdcQU67pMZahh
R4ZuMpt8uge7+I5tS2VXl9J9iC4fH2cqEGe8x9GEyFJHzMaVUdO8hdkV3/yiGE+x
riZwi2GnSvZHJ12rmR4z7KwqUY2/kpkYEt00ywZpIbMar2GXa7Ap2L2oyNTkFtQc
UvPq1aCFUCUiZ4sRjiHLxFpLFIgZ9gEnuR5IWqgczXfjELSLCpMZVz9rP+0Qrra2
hR8rhsY+I42WZGua50RpGRS0BU3nDptxMidr8fZJTUDAOlJBprtY0XlBbdgAjpst
ous4fBBI1FwZrzVz51LbbI1XIBvKV9vaXC3P4WeFC3DT80TOpo2k0xO7ELM6V0lZ
+wwQGEFzholkG/n7DItpIr4uHNvt2EfubzopPbqXwd/ezYsahpNoLxN9WuzT3EeB
D0R2/Z5ufabZtNJn4h1n/zDyM0VsysFyT5t1LR9GQthBygQ/AZunKIK0bjBNlIxt
bgctZ0eggLgXDhjYLSzdHvXwTdlrvimikDHz2BMu552qnjhNXFkYEVr1tvQpLKDg
q8KdJQasBbJTv+zbpL8QH06eRHUMXgR/ccaSNk8o8yRNfra5owlARhylZ+K04XFq
lZWvhlHVP7ddE0NgIZDPBzp4vw71yhA4NS6wuHguFVDUPxpWFq7PltH5p5Gc0iBI
MPBJM3G0QnkZjfSYrHOMSosXeeMq/SM4Ty3tZ2Jly8iplYUH8J9jvA5qNOVB1PYN
GsTKcufn4RqHqgycSxfJ8UJM/d/owXtSwSnI9p/G67gPFxSQhiOnbsCejM4Z/r13
5U7JkvGKq34r4kQ8sxtJ56jR/S6hfzorgqTotagujWvoBt8UvC06hM/nCbSkZgw/
VDAbYtfVzgjjLLZyHowHNK4sOInmpvYcofjRMrP2+hwDeAb0md15QXPi5gaieaOV
SkfSvafqZPEvpvzybNeH3088o82/jt1cMZnMoScCPn0E4iomMbuhG46srAZWm2In
c7hGVp1B86cAFX647yo4dHQ214UsH2Bi9MegPksG3u0jKGc3RCQnzPlxVaa5e247
Fgi5XNDF7R83TnrxIXY95eI/RUiFpwpECuT2N4B4hpn1Ax+SpmYzu492MZIgyCwr
qxou8A373zXHWLlKHCmxeb33uHdjHI7gMmGeutZ3h+AzAVlPRvlOQBdIlcQk8Zx/
XK03S4w4afgtBJHnHzwqI6glGI8dXgNjolhLA6TQCVTHmaH8V1eJ+kawLYxxB0iR
jGncLizm6LohuCSTFHYo228Bv9M3AMNdWo4AYkDD2zFzlsqhg0bcPbEjCb7mLYwY
krOIHm9jmt2AQyXpJQM6w7vLljBoog2FPWJvaMdIy2FBdQ+L4gV2FO/UCiZ5Z5FT
LJhR/JptFuiVa0NDvoOCsZrEFAdRMYqm0BTm81JPzZ5T0YwSr55JF/9J7Q0MZCuK
LXJM+vq9E2goYmcJSNOXEah+YZbQgpvOBoqVG708f7Kj/q3DKxwQnjrX/oGRbVNF
3Q4poa9ZaovpvtTSYGwkW34q+dsrI9Phx92433i/NP2NbHAihYDFV1YodMvn1XLq
3DaMZSl6n8u9aqtc8sCQQ8/pmKUkhY4D9ZX9fcEntSNUrlwn38fWhky6CKmQaudd
5xXo3I1LM6AqWWbTpUgC4gvQlV3J0gwxxhDkFM/Wx5T21PDcR3jee4dxNjNLzLqT
g4zNhBP+KaMvQ446ZYly0HE4by+XC+wvdJJ0V83Fw3Qtoluu8stEDutMLr1s4+HH
tMJJy2HM8QYXiexfvwIr5StBkrKO2UsAacruUnb6SqwMSWKmg2BYVLU/5eNQWEuD
P4klJ/23tmUwiWXUpu5MS3aLfGhUsOuJgVtRvrtQdEW2r3kUjE+Ukraqoe3rng1c
KBZPRNR7UFV2vHIkvYJ38n079jWgG/yHBLaKTM8FhrTHyHsPaTvRyHNWA4lErQrD
OODxc5ntVGOoIb4SnN9ILFPtjeO3qhQ8PXIzOgqRSxiCnKUjUsg4bD/o3w/pzL61
DI/9opUDzw/xGuNg+uxwNGxSKYbxhZYht9Zxul5jhZpiNUlrxZwQdY+Z+x4YCTpi
BgL2wcgtH7r0ETVtUtHqNMA+v4TyGWwkX2K5gcnaBhznNHKcdMquZn0pLovODSeg
FcfkhFgjqDBYg5M0KEgTugKJd4VoSLJo3tMxrq0pg1+1h1W3aNype8WLFuvUyQy9
NYE4ZHxQicPjQZzO7fxuqxpJjf878a0yWAkuJrSi7+kqOBq190vIjOYUd9c3XLMV
Dov6XTB5FfOxM9lP3nb1eP9OmlpR/6k4rxa9lNmuBXZ6Gs6rP3Qkts0YvmREvnlI
TCbYymDhqawguQ6jDtDXL1a89zU+JsQ4ZGoMyqX42mYZtkeq33eqKnpZP0rRHBv6
T8G1w/XRLEM/b/11K/Tu/+PTIRUR4VQlETepKXFXP21cDrPzWnKHrT592x27KOTa
Hsw9V/RseDDi1QNn8QOH1m2Ue48PLPZ74d8WNtis3uYPKdUKd+nAkiaF1vEs/Nbe
zNI2XshzH0F5ZgciwfSfVVTG9u4ahrWKA2rakUWE6LcRM+lIe3+zA4mvcY7L1E+O
FXBr5Kpari/vBXYLQB3IdI0BsecA1XwAGcFQ3BmlB8qCYcCGCQYQ2It4ugr/X17I
SL5kTpVS8/vrnoMbo9UI/w58PKidq064sHxOHYo5SoqLnKaLDvY8isIFBgo477Wc
zedphVA5rKtukpQzR6F4XfZ1OTM/ldCJ7u0W6E8bT9eJFUjYQtjHHZpuxTqyG0Pz
8O9LTb2fWpNM1hDsA2+KQTLIl/9rfxbsepvD7+k1mqK5cuH5zMgMP6q2P4KjYxdJ
Z5x9QaUoPhGlKYcsap7B7WFfbDb+6etWtA+qHoKr1LspefBZyCdBtt8OB2ZT/rx2
4KkHuF+YsldyweVUHjvMHM3LZK8oSU6jpp1I3D2vzDctae2GLSUCG6njQ/XqFTCw
Vr9PQ4YpuRXwcjZYoDmTNoTx6a40j+8JJhCNK/CK+ItwJ4GMYq7P4kHQDJ38mYV6
nvnpbsHTs99SJEzbS8fdFe3ytBF3NTxuPrDCDdWMN2lIlZgfUwMuTLozV29ROE98
miDG4KLozVIoxib6nnTvgN2xhHtBNjkg9FyRAyHQ66JYFD/hcOjMhUOVXsUroUUw
sR2XACfW87VimlsmFqNL9szRd8MKtsNt3KZv1rZvZtxe54Oj7nDc2pDyhbw0zppa
XWJUfkkOvIrV4m2I2apxARtYOeJuHLTEXXi/L37TGGbFnrcZip3Q7ZZCx6OdHPWZ
V6XE7ecPE7E/hvZGlrZ6FfAfm1FH21/llmKMRc4eXxqiAckV1/KX3mDJBxSxVKwa
elng0A/C4DqcVCKtOvif/lmF+njdCOUFZyb/UktegzsLPNQQJz7yfAjuoqXCuL9p
MFkkFMtvgVLiYyRa6wX5hXnhG1j+yw6qdBuicvbH9bjz35uNE3mgEJ6SCVPg8a7G
sXEGBqocal3vAJKMEbeCoZV3EQHd79uFeYR/oYRHrosH6kd71FPWRE9PsfRdtVJb
V2Q4kRIh4KiEM8976BpFNQE4votuQFYGGDrwwqkex3w+kl/YAf4e0ogQ9X7FegMV
mmJbhCmtpdfLyoNfHcAcxlBsiyKzHxCZ9410Ys+8+YsCuI1BU/nyBO8xslejMx+V
s60aFr+D1FYczsqX+sLqsMwRnZ+vGudRP9ug/JLyORMfNFcLg9YVNdEiOqzx08Ln
j19hU5dC3Y5ABl31Tg25XL2yk2f/D3nAk7ozcJSelTgjpa5O0fkEiG232v3I8Ft4
UGylNcZAtIa/cNb9GIzoXeMlJCPh3BrxZVUg11p0GgcA6z0jBBxUyVdz9hMZcG+m
kOtFDtvS7iAlDjdvD1nR8fCBrzm3fQkgi73+cqng6mTpnJvN+UOdxbsbyXJbwm/g
vFYhweehUxaxYTPIx+hCa4SRDaKv17PYcaJgapay7pjGqKZU22UQSG7Azg50WaIN
jk9Nsa8Cua4lqmKX21LyML3rQkMYi61cgyCZMF7bF70oz4P0wI2WL0nfFJuZMkFY
Kg84hxH5WbL1KC1cMwfz2CfVAZICptGsIHRIaQmIQjmqvneurRxhBsBKJFLT6EXA
4CGuex0H8r3Cyi0ABcQS0J2/46NiBLhBBGOHBL4zo2zw7NoLKzLZH9ryRWEee/KQ
pSiTWMxOvHB0gvXtGAco+g==
`protect END_PROTECTED
