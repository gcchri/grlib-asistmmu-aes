`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/bFuVUkbGKKH4/iaT8RYjl0EgJr8iQp7CCYGVA/m8pmSVB/aBJ7wJaQptDUEbc3q
jTHBdMFDv0OwqLTpjGPXUOiUp7b6EhL3Av8JjT1oct6ENV6StKtr34z376Z6Erw2
1wd8azAC+2yqCEZokdKap1nd6tDbf8Y4LD9JdBZsVkJ3rO1EDGtdgTP9tTR3VEDE
xE7L5I7aEQiZ5WGRBL8ashrlilnt+ffpo/wt2gT8ib4nPL3MlzZ7/1GVKWO5mwux
9sDJbhI/RBQwFeknCRBHNn6/9wPmSk1IZvH7PPFnwewsl3eK8TUfMXwFgRTitrpA
pv2cLKya2OQ1EmbKva69bnaMIJ2btVJLNrpa69kIthLEfBvO7PJcJibIMUD1YtJU
QOdfW1/kQapoRdSxNsn/wQ/azyH8nLq9lwTyrfBxR6M=
`protect END_PROTECTED
