`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HLYNBxjDE2nZplXiHa3qj+ksMFsaEFAzrSrKc4RRdESM5N67/jY4/QnBc3HFE46K
bgPJE5aSoRuvHQprulj44ElbI+Hizd9aBS1i51hH2ax2krjsWDfkPyrHFXs9ucFK
QBKappY4geZ1NzUWDalzur/qKS/j0UEK7eiWogdtuwP+9H8d4121FDLDrM5ImPvz
FymMmOyK7OxB5I8D77jULfH4ae9FFpIKfiZN72+G0XWr5Jv/+/Ptq4AkBMsdsIO5
0eO17IlFDyie7KppUt0lMYsqzgw/I4Ck/Su9ZetYEGxVog8rwudIz8NRNtsBGyw+
mMngLSgKmwfDgOjkgzvMbg==
`protect END_PROTECTED
