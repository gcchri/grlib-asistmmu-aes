`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NbdPBiH+O6jxWJk3JrWLP87x6azha04cvfEz6NkBSNK5sDsPkfDBOcqGq9hSm2wt
b2kxlpQ6nQUdwUwW2ha/Sp+unwOGQRvq3ATE4g7VEQ89PsHLgQMOwEhQ4DM9+JGv
mgkGVtNPX6ftFCy0DtpGU39Ioo/aJG6aAw+V990KEpEw+gxLZrxTUEw4TlnvwPs3
Lj475LBHh6+JYcRZkXaFOqoMF2/mJoxEoX2HqR5rIiDcPcJC0GA/LOSn0X4QdmEj
+3QWhH9Y4dO6zMcMr974QHpEBQ/p83FoX4nopQDPaKPRroCc1NIbRBwEWBij5af8
aa5qA4fI7U3ght6aPxkmsYpzg+rVGl5CHMAsM9S+FRRrc4nAXDGx9AHvXbmChUow
3mMyNXXrl3D6J3WogLU7FMFJYRP6Csys8QXmcXy/Y3j9e4LdfJVKVF6OdrVSUjIX
gbAS9Mdq0kMF49nWaFg5vRqJ6wNdz0LGWwJT2KeDebMg6yH/lUHeZhx3vTeAYphw
nnC2x5LkskEfrvBAAH6YVwSWYaGSduwTwxZ4Z2hx4bx3yWhGcbH0Ni793pBh6RWA
ANqhy8fJZebtVWiJuInb3pQN4Ha8g0ywLeAA53WcddLEMxUKngcEKHHO8WiR9Dwm
Lprw7LUUb4Y+oZX4ZGIT0PesCA56WrIeIPkxrzBP311wbkmWqeSDp6byzN87bhPt
t+idUkhws/Bk6ROe1AwD9rcdhpNa3/AIhFNZf3yclk4/st2NEhYXU3kWYZPXuKKg
alhKUd9Uvvl/xmVO1ANRmPRigu6xu0XcXKIFcCR3dxnvDi3AK1VPcHYOsthhOPa5
ZVvIIuAwzYFni4HX5c/2/58r2T0JdC1rGrOz2gHmBdI=
`protect END_PROTECTED
