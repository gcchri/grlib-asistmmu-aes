`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jgql1G76BqfYA1z1QPwGGuCs5FV7edIGs6rH/8AmI3gQa3AbDHzt4I5L6zkVGgRj
fJ6xRgWdOpWRNq/q4ZYItaAMnP/NqZvnqcoC9VRA90Q9H+dRnNKWA0Aa8nRf+jaa
5LuWq7mTEuEA97vzgLxKcd7NNNajuRH3JnBCI+pWM9lgzuYO3gTuZU+444qhhCv1
lFxjIozssSp6w8q29/yhDgdoEL46eeGWUnpnyse3N0drW1T4In0w3eA7G14JdgCP
aJvW4aFqIlXizJTgMbVRTI3YVyKPpSDLPK/b3J1gBQ1UYF7KqUGebGS0QzOUhPWc
10g9NDS3BgHlekHxRGIgRQhfaX4zn5kXIXbXDiHDEav6l+cViqdAVYu6VO42MW/v
UOvpMH0MBkpxdAjafIGRCiArPAeAeGL6qpNPIf/FK/qMrl2dJ5eDv7jH5QfPUYfC
shH/ahiT27pj/JrVwq7WuAEQnMeoqCX0nlzPUOBEQsqF95FmD51u+gxe0dhIEZvk
tZeApPFJlqieGs2AQbB8MJMYNQTL1kj//4wC2xT+YPv+l9SykiJlPf4+/Skg4Dsq
eMWARh3LfDO8HvaGceMNFJ+vZt3OcuO70vYeUJmqEPBaZINQCS+oyZtN7dIZuSwB
sqxQoZsm/Lrxi9VMV92xlp77b8DTXvNc4d3/IIrbWjW5n1WJm1DvT368R8JpKXRJ
F1434ZoKu9jnmUtI1vJCuUqjxuLx3p1tbAwhuyT1gse5UKIUgFxAf1cCRZEHUC4o
8cDfAr5FBCgbe9rZEbPXcrONJuniL+2iswH6s9uPDMXOfrN78ZTVI6x1atwoZTXr
NDht1nn0uf9m4EWSBQd/sIGjD/CglIld1m/ojcx8q4XDtLG7cIj+RcvtpSiBVe93
2ZUm7mKg5XhtOIrlHryyhdTa59kWIp0lh58YVhYq1mA6O2370NDFUGQVHZ8cJqk7
iUDPpMZkeaZ/nB6LKRvZlQnjSQZNq5ZHp8BI06BAsAFFpgtI6Bpxez/fXCrT4WsP
6W/vNDZFIBcWcmALtlsF3wCQvjywS3lt+fVplJQhISj6Yw1BmzMqoYEFqB+ceVeQ
53QFeO+qYUM9dGz8Uq4MQMUlEqwhVaevoC6XvsBYLrKnK/KfxI2BEdFeDixbfMuR
icOP06+kfpiyrh1Ny+JVrpAJ/JAXKXPJJRZqOMH1U2Ywe+7qMaTzFHyCMo2wc0B5
iqqae5tHOPk++wmqt7hyRmVmN7BS/SRPC90PwZfFlsKBW/fdcW0AGWlfBkr5J+bd
SoP0bjWZDKZEKK7Vv+d2JtfVUCK9xlDTV38TywMJolfancjRT/NiJ5gcWe0BNXu6
W/4tljy5OeoRetlbaLrU9gFpG+HnP36mmlvdRf79OF3HPDtRWM2KqJTbWvgSj21s
kOlWytrAQrTHL72j7rnWoO4yJ3mwRrhPFs1A+hmuE3fmmc+EVTUWjiDpLtA05hjk
KR/TXfVaPxXjVsnUDyEIE6Jjks9jDQs0i2cmJxvpBUJaJKksQYSNjhxn4f2WkyTI
8ovOu+fBtIFVhhfJYsIoqC9Mv6ZNZT/RHYQlGEARDl/Qk7tSsR+hQpfOv8gCiqRJ
Uf9dWnA0NP/6bGfRelu7paELx2XcF2xjjp9EPc2avpwDpexhVU76wBE0pgxXun5D
m7p6yfq3oRQxmXplPVIVgb2Xx6vI5JlulPUYCjXCAPHyV3osY4ER1bkQ5RMvPKC/
xiBMECW+Y3JHaAnCcyYh+A4Lm+znO/Bo/4a8Qq2Qjz7wp+S+hvyW0kxV3UB5zko1
pf3azVDY6N+L/0S7TvHqQal+sZ4y50LFXR8EC/DDGYcWMV/uajgJUDsE5bmUlr3x
3lWME2fWZLtCTr4ILJwb/smQk/Emij4eN5RCRQrW74zCxuODAFXK/Oh4zEgZPSwJ
a9mpTVcWJYiBWdV0zSlf0YCndOqlhYyVJh9c2d8XOrod/ZP8rPgclFGL0R/3tXhJ
B5z4ofexQhZHiiqrVP/+tf6fPrFajr4dY8SnSivfErkf2VHmgtqRKj+uwSQLu98s
l1Ponwa8Jh03NgAYkljWhIAXsP8esopApGNP9kgQBvNbGDnTvI2dp3P7GQ34sEad
VtkNUUx9cYZme8lzaB2myH4BeenH8Qe+u+kx27ueO2w=
`protect END_PROTECTED
