`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L/Ti/VXzZ5DPCVjE0bQlz5SwWr50thy1RReWO1NPEZOqtdB1zK84NFCRzuVxsw9i
LFhh8FSyyUi9i5wrivJLO/vqoCDKXnkhjg5HWKsbPFWiLEDBmIWgFvYvfzrNxSSP
Cm1I8VqOjvJxZhWHYddvKM10gqDEYypCFwoxkhCbg790V9kYptoMjSJY8laKi+dG
lVohyCF45eciklhwiWYC/j4xYwzQteiUv4zdHl7ctzUs9Tn/feqVRJrHavTHfMZ/
8IBx6zNdz1GpXHNU+NjjUY6qrXvKM0ByIB96Ov80D34pClrPFczMNPINzUVC9XS5
msd505rIza+721jDJL/yjgbM1zEkb8FiD5sNRv+FwiRNS1cr7Dfk5+fmzm5Ypaxp
`protect END_PROTECTED
