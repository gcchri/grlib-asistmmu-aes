`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NfcYckLGz0Nx13LbqEgdTVAVbdNgcg/yZqJtwD+JVl/jSwhSApcoC0XJ7OXsUM6U
0EI0GYdn7qWSHd7QBhD1cz4pNt7MKeEWAXwnZvz/cxSWjSQyGMDA6Kr8MtSxwZYB
+Ay0wqv9A9DSOt3URsUvSw9quJA/+0RnKubVpt5NdtH1yCyf4/3idfuURqXWrahW
pt+NVv+RRWrO1qUJU7XvZWoIzHX7jf3b+W4O7U/z+k6LTAB/V7AmngOK2EUq0/Rb
ZLL6VXZmqBv2U454iLrFdipRTOIrkOCgeH+fMZB9BSLZMyN9fquKUniXBPTYmomh
ytantLm+k12Ng1hEgbfyyulYagDQi3jCGiokSXmWb9u3/XCwdoRkkEUlMHA8RC3+
51enCf2w1lyIBUx530n4JkE1ep8D8BCd3iBlezDl0HRicPb6Z9J/Xp8ptDkmNc0P
JNziny+3FQgVCD+F8N4kjP3ArobmMJ7FRVVZra92bIq8OHrjh6vasNf/7JqyNXWP
`protect END_PROTECTED
