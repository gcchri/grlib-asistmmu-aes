`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iJ/aHtyjTCvNutznEdECJDCkKNLShiC3qGFJ3Uw3F6C7eS0DiNcUw+3GZ31H1s6x
Dfz8RHTMT6nMl8ZgY2Oe8hAiimEEyGmOXERDOxUBkYkzVquaCZovNmMS7F8N0M71
Zbf+ZaXYfDpoyh1pbnUP9Vo+m7Asmw2YpCzHlSaVXk6OBcNyQ4Jj9DQDPmqB3RIf
I7rfDKhDlWigZxAmgDk/UEng55N5RzMab0UvXi04xtAmGH/z/SG1OmP8i6o2pai4
zXTRstdT4/ujycf0zFOVJ5/4pi92cSUnhWEPXs8+HsPWBIKGY0oLklH49E/PvCUw
xaAbiVZ1tp8hGlZxZvXa5JGTHtH8hHTr+diEDuYP2OUzeuW4OGanZrpdhH6Ijelp
bSyHJMXINKYuZo2SsIUuRbWU2awhUtVZBs4p/FN/vy0=
`protect END_PROTECTED
