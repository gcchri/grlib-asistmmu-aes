`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XPBOwAAzJeuWx1h8/49Q1dagx6iZ5PX/iyM+CsoF2k9D1kg7HiSsTcTEUg3aS3ir
aAMi0v241MNcHvo2RIp/q2i6n8hqlBVPZXl/fj7tafW2IJTtK58KkCeF5IVAKvjL
8hrs3SrYEf3Q95Kn2U2LfsOnqyTzHbPolKc6sUnotSQ4FB7xTO2l9FoMd25Ydrc6
fth/3DKxJBxBN0HxHJe4v3V2vw86aSVh8ctP1hWEfHe1M2bR1yNjuTFiGC2RoK8K
UXyeTrGSClq5nWFdPuHAMC1hUZcvYPgAqq0y0+9/4axfBqhU3+LWQ2G8GpIRPPmi
4VXi0C/9a1ELpVC/pKa8Lh1xbZ1+yAa5gBFsisGtRh+L1HLUcM7K3eWcsQ5Sfslk
k2kWJgfgoJPoYr59hE9PZ3d8OyARf3tf1CuVpLsYSSqKvCfuZrFHwQpAvpkDQ8Oa
`protect END_PROTECTED
