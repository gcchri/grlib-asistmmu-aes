`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tl6Rs5Y9xtaxrlYJPRDOuDWwMZ3lNdr6vVXKzidMR2fdzGQKT5yJxNXw8DWCUjNw
F6y49P8SVzP8Aju79QQxWXVU3R9py94MmdvQsNZ3V8+xUu+SFjeljMLyxFGcKXs0
l3J2oMEaBr0q7vQpWYV1jkQCKpXcT6DqmiTaOV3b7ie1tCOD3Ez6gXtdllE1xB4+
raPK6WRmvaLv7ASikLFrgQbq7RcKLODQWpzbZb6PNxMSZEOtCPN3bOBSV1B2324Y
idvO3EcH3YnpnHWpue0Hbdus35hJemRozTaEklui8OalG+vnu7o10QhJjCc77BR9
rgJ/XbbFd5PUGZGzv84/gw==
`protect END_PROTECTED
