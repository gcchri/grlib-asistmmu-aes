`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fPvhBi6WCwZkkDXANkjFkk+gB370BA9yFc7HVxiQQENHTIGpSp2TTmWBcH/jYOWE
j4pwPlXHuUiXIxrouRAnxK6WrxrvYXeNTc1Y87wbwKMrJjPRCxurli+WECoSoK13
mNxy0+WCNNvLlJIbb7AdX/E/cPh5Kdv3Nyz0n6gdV5dfs4xAlMyBl3FKIr/GqEiK
Ggl8SgZfVkaPQH8I0a7f+G8sz0hAmfFjVTFNZkAkHsN3NcwmonLUcthYXmXjcLiI
f+nsf3ZbQHJajBeYKD1dQw==
`protect END_PROTECTED
