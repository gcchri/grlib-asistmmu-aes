`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vKu0eAb+IsIN88aydVNwODCvl6yGWTekj9nGbqJnkUiVhj6pBCjhtUW+vcJTdP4e
qKVEojoQ5f+evLDPRoWlfilkMXCEBm+eNUqF1eZgwvpHEJryaVftEDsiXVLFLQIK
iYSRfYt+BRx9nImM6Hr3xch9QQIkrWMdKBdsPyvUk+SbFZqJIyrf9wIsY15I5amR
OmodlSpHkqLCTwgQAsCqaK7SFkyq4IfhUT6YaffIyWxY4HXkroVkHSIo8mxDTDJ+
DSDuiFMom+71EAcvFJI9M6hQfGOQ//kQJqjB8wFqG38uDbMRKkQQdvNo75EWdeB6
7vQAnIHCnsz/kmXDWVdBh1MPf4FGf5icUtCYHCvxz5oMJFg1kW5ngSPNI3eSsK38
c2qZK/4QCfHqEQ3dCcWQK9x8Nc1Ox37dbuZZ3Y7mH/WhDB48OsSefZePCJ+N7vXm
kwXTLgm6+qrgAIwocu/DvFv3ufQ6/U6uSPxixbG2S8MNtkaGcggdZ/CBwk+ucuuG
S2S5itRYvOmKjSHc3vqENA+vUWVGTFLhH7+RfOr1rGfMI+7SMeUo54bOujvu8T+u
jM9tSdfyOBlunEgy03j3UTk/CCa5TF7KoF1nBU2kKWmDTa8DVOS+t67sv1aQJleU
VlpY8UX9QI34adIj4FzOPy+g6TGGSJuJI+PYlnPvK4fGHKuabfLpijBpfGmNBXhS
WKtwgq6REYuTjWI9ItCOc9ZUSlgl/jXE7F/96ljdrpCS+dAO8F9g9A99KduD2qWx
ODeW2lcWfrZi/k4fV1qTc6YRoCRqN0lBgzB+FSj/Lutvj46wfefqLRHpQnjObxkO
3LxFbxRo2wFCueIHvXilM69kcFM18VB6ag1LhGfEU7oNAkxPU7KZkISKMOgXM0v0
i0eCc2RLb8yhrxi44Fvu/xScaQbrkPhHdfxmPLVmhBIPG7jWRhZ8XtEkfQcVDFn0
5e0Gtr5OYHLZoNaeOWL09FXpiC1Qags+99+nVpKVcqDuhBUUeA3njtcaIX7pWrBQ
`protect END_PROTECTED
