`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ptzd+WR0vlJGYReDSkl5iyKQ1zA5PTOwoPyCzm0q3NdS+4d+SMHPC61vyKjRQLDn
abBcAq2sEktyml3BV16yF9cEHZfwETwl1VqP3TlbugWsN22lYYTWVY3Er5USHaD3
lBZd0XnxBeey40rs33AMTB6RHaS6NRQkYkeYA/FXhxGxUydcD/lXuF2x6Mw2tATp
21+ZfHpH9SzenR7AIl5cK2cdbCWqJHJSK8rg+8s/Z8VoZNyjs+0Tuh+V7tiOdeVE
O6dPwoGm3+oMMryY57nBFHQx+ubB9PvgHiidg5kcY2bKLdual+PDcB1mIommZwcJ
2T0skQ+Tje9F9DMO8wlXW7ScFOz3cUHKImgAedfcLPq1jEh6/Y2jcyOhJksorMHr
FptycExC/4hbf6HJbN9j/BXKYEUDcJTW0YKJaBq7dhAAEk7q17qHslzx6h4zieUG
mL+g85B4LnqCdw+OnPduI0oG1gB08yFnJnM9CHb+JHoCuzbKJrduQzuAwIfzqWnD
KPrq2UTDvSCzOvw9vQ5ualMXPn2AejX/VZTeyEAcXqoDo4bUumDqXq0ORc3ORCel
V2emXNsRMutzJfbGgQ5xwrJL62xesR+mpYHG1tRYlUeZ7g/qWM96D/32ssYYVnzm
use1Rx5i++LTtQ0Q1C05vohu2XGB9clMQBPOIFPV0WcL47xHcfiGSpGPHuomO/Z3
H+ZB8U3dKK9aaJPD3c3OBL8yc7+ouhhHjdxw+YrUw8BdyDB6hogDvnOqcFTGL2mM
acKRCXiOfnkExqVv0Nmw2dDZzzlj+A//NgRelqaM2iAKz2YJDh2dZp4Rv7REXgpX
YUiO4Yl+OC7vL6OjYFijP+mxcY+q/wGnLhRXormKyMoGdU1pPWg1WZBdq0Vj3lIi
lwbk/mbCUtabKQ4MiOA9p3+E5zBP+EbntC7FPLw6ol5NwvDLXO5PmKOsM6ve8h9A
cfeANiEp6WYbHv8SXSpQ94uHNgCGxXJch/W27qDNXrLkPFEULGDMEDLgHZTdeSuE
ELvwoYZWL2qEWIsv2gV1NnS26PUoNz3eHS5vYUiI7MeSptmf+PMGD7lfxTh803eW
YIhVpPLun0QlcTBNiz2gIiy5WDARGkthnUQ3pOD2lCt8aMrhgNq8hzsCz+O9JJJ9
KYbdozp4GFaxlmwXBsfFf14d8rsl0TDiggAYPswnBf0xPj0q7iCBJych+9/cRKVq
wNo9/nhfLzZWMcKlmAhKu83Jt6GhVFWA4h1ZDtGDv3E=
`protect END_PROTECTED
