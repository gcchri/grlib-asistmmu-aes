`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DACyRKZplWwmXC0u/g7Mu3R1Wwp7TTYevEn5fkHC8uwdPhp7jVW9z6+sGxLjjBZy
kDCjS1qYZHSRDBwK6a9NjUly845teqBsax1L2nZgR/6AFK+86ubMoe7cN3vkA81I
bAo6yX8QQT7o1hxRo3pmigO+97JDKAxoyBN3L/EiCN3EnKpepBxPnx9my2vVDwS8
9Y16h7cn3w7MLlY5NXlQuUvaYYCcWmZu8YH8wjiVxcHCBJHqFO2jGMmU2xVKhkQC
XvVPD7F8bdK4DpzEUJpB9xgmntENMw+HqLlekaUQguQ=
`protect END_PROTECTED
