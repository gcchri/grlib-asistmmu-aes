`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kD41vw+STjZK5s8ci1AB+qF4QO8UXHVzpmOHZkykavnKG5Dsf+BQRE8KfdPV3BRk
3TdIRNM1mFTGQAjA4K0g7dzUy1pLjJQeUjVG6kPEtc8UqZDYqsVp60vAWiZFaTrO
6A426n3eyCodHMMDJhw+PxgkFaaAIbClhe8mZYMgH7Gnn8iT+xM8YjH2Uz6FTBw3
9G/ez7F9Pn7cqDvrUrr0G8MVlc/l2N6XUnmP9UzUTEcL6+O3h+iTHIXY5BQ+IG44
wf7B0KcZDyPOP5SWwUCt4VJTZxDgz8JN16nuz0+I3GRbCH47ytN6RuBSH0WHnLIe
6O9ujm0uucNKoNYSWqoitYBoLWOcyq4oPFRMMp6e9I60Mi4jJXgHV+mKRBfqGz2X
ZL99o6aod6RIkmGV0jBKXjXBhjhMtsXGvutQ+Sry1Ho=
`protect END_PROTECTED
