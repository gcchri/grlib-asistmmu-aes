`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x0lIo+4UzB+jDwpeJNPm2yr/cs6YxzOJiWeGKYscEQYvrS52oB1kdMZyotjGg58q
72/xwCltNZcaRUO+idYAec5eezezyeEqPOywOgHIgdJp/Q3abviiCformEOnY2NQ
PlkoMcmXK0+dHAkyqygEtxnpApT81wUVxASFFhkczTSRYxJM6oitdtwhblwZSBM9
SuQz0hMxh0gjJtNFGL6L6vmarYZKt4dG6LCJ5rMMREQcbO8f46RAOf1oUMs4/Kxq
owOtuuGiy8jg25am5z3eTvKw5TNniKXeTZYJb/fa8GDtuxnr9mBFHv76tw27IzL1
qNSYkcUexuJAc2M10+W9+YjpHu9wVVvrE9xRrpAim+7EznOfxhkTzDAcQORmzrQ/
WGwt19Mwv01b4eIv3vkYBjP9UbNMv3+ZkuSfd059Xeu+e7EzDX7BAwFvWEMRCHJo
`protect END_PROTECTED
