`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3k6GGaaIwbV+/zv7EvT+BPFGTuzQVEV9YQWYCzbP0WWmbzi9YLrwfgIupZF5Lbro
shvMG1qpFgHCOTY43+Tf/uN/91mpiaj3ThE0o3abpy+HYZhAnBAf6ItHvmH9oP+P
11XjBAFMtOdweDEFz4vBkN6ooiG14JkowmGIxPsD/TOv5PRNNHLulkrwPqLG7OmC
j0G6AI6YoDNu1w/ooPl/I2q1zesHRIacbeef3hrAshfFEchi0t/fvQSqAAW6hWbq
1fsFN/ShapEiak8+dmHgbcgFjLqQGtM59LAbwsY9e/Z7RbGNnj3uxd9pZWRlF1NF
GU8xj3jD+LsQCHlsFDKeSPXUeRVaY4tS9TI6Iv3h/ymc4g0w9DLXyGE60asOSS1V
UGSlngjF6DxgCc9OXVKyNY7JgoEn8ZMRokCkoQuVKZw=
`protect END_PROTECTED
