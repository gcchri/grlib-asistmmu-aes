`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ND4lVMzUMrjJPmflYlpUi6APKhe81RGNRhxpZBql/shXieaIOUhM8F5mWQXnkiz6
d1SLOT1vv3+emozyjEkUY4yJ779yjnbVET83Jk5jNqeyD93otq3ZH4ax56HfGBvF
FTPuXRYMky1yqOQDYia4F4VAY/GjnrJwE15rR4R/HpO8PrAUdOA60e3hMnH4g7K0
qlf/bFjo87XhYE6piV4ixScJiDXhkuCIhQNu1YNjJWECzSMq/0CkAnyt+bDK48O6
r+z8P0qgpbHUKo8JKJbkEB2xiI0B0r0THL00FuOkvMa4+UYC+ORG5Bd9UJDRroUj
Ye50BkYk95OiQz9PFA5KBpuW7QPKTJE3S0XqWkNllVeyTQLUu3wvYTYgfcyiCkB0
dsN985ax4/fcp21FJ2FM//1maAJYNlYukvDmb2RHqWaDKkWxFelwTX0dAeY9vPkg
zyXie7TOAX9nNNBzpnrZnlm4Va4IgUshiK7Zmxd4X5t7BVd6qxKNJ7FRHulScrTg
gSm68E2oisFzwno8fml7Y+KHWbQCXFy4wV2iU3PQnEErXx3F2RAcF1bQJTlY9xDx
OxcAMZXJDvP+RFVdOzWpA1I0R+V4Xjk6XZhUpUrVw3Z3FDMPVJ5h2sjfE6vh60Mq
C4J0rBpNE4t07QB46Yp0s61+zeYknU3/dwnHTB7bVhJqja82AmSvopb/S+2tjIOQ
`protect END_PROTECTED
