`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Dfa//dMnmrWhyNYQlsCcMJlKRsYVMHh/7r5yax/imWBMwkXldiwJmbzdMGQcBC5
ye73df7bMyxk69qjmr6hLafV9b7Didwba89VXItkEMCsHRCzdEo2nvtDBigi7Jzc
qilHqZckKjjD0pIJoVwMHK2VE2h4sTkJejzCs4e2oMWA0eU5lW2EDBl+F4mDMc8V
kCeuN/yqufpgq2maN6e9Pa9XRtH9ZLPMKv1NDpfRb98XoGWPqVAHL2jgjxHG2wFY
3bXmz8s/AmOyy1Nw4SF1x1+0UgA1gxfL+8q9fv8w37gQWmPBDa4P3e0yvP7AU5Tx
14SH5kRX1BlNHg4RMl02/9Yh9yJwwz4YhTOfEF7smldTeqgcNRBt9sZ6zfC0Wuy8
wR9uAMZuErsVhgBp6XBYU25a6F++z55MylEU+ji4qXxSSAj72vHomLbfDmbH6HdL
xV5Ulv5yfKRwYxdldhW3pZL2i/csHNIflINHxgR/ahEh5NunbEd0/LLbYnU5t5Yw
p1zkqCovIQ0DU7Zbc0NtRAXCNARMkjOEp5BMbp9d8QQ40dC9Bgvn2BAXst9u43Zf
zhQFNaU8kMf9ovNir6x93Wf5XOtWjp3VxWFkAXT5Xjc/yLne9apVxVqtQL9pdsjp
w4xK3lunhy8Hmnlvqobu+3Qxm0IYNxNj0GdWoUbT0v4RoTDmx/P351JQLmW3gFTd
RJD/1v60qiPx69FV4kujWA==
`protect END_PROTECTED
