`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iabDzuAEkL4VQT7QgM8JGtpT2g3qfJmzOPqtQyGmZFhxTWpeV6qa+ekD9/t+ow3l
sIZ7v4pRib4TintFWDEjN6oh32H9ORjwX/GI/E5rXVboHzSUibtPoOx+E6W7ZOOX
wVV6qONHTe5r1h1LGDs1v2fa6yAtTqIqmou5D+F8r6zEjIkfzHGsEP8q3wh/GWew
SfkSDBeMi379Z1bor/x/BwKH52zsgRwR+scqeuLg0asKFxChcNLKj+59X80+o4lA
E5mc8LwTnfkf8JaBdXCjQYkkmjgxuYRudCXOVBM9hDA=
`protect END_PROTECTED
