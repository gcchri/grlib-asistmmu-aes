`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z/mjdrr+xSdJHWIMOT0eIWXtWFnoq+9aZM4LrFv8ey4JLYKavjVPCN1HaiDIUrcc
YinQxeveF/m4wUF49WN5rpQrxAc/LT9hxTXs6O1zy8bJbsZ+wpY1PHALPhUzARBQ
JG57VuYgMMbutXDLjkh/qHrGz78g9a+e1yh1Y1Vzpc83s1gLj+14L5TEeaC38rzP
no28SOJnkK8dRRMTpagiDodxAgAuGaWEF2jpBAuzrrO01QgyII/DEB88XLpTCTxL
WbLJ8lqoEJb6mw4xS2/ZwklLHZPzefw+99kH0D+GQ6B8zw+TN/4uzRhbRCkzYiyR
zS+GOS8B3VZSReJXUKXUVLVkVJgd73GQsrtg59BzDXrh143nNarTxaqGwXMA3gd8
OsXa0NKOky94jV6WD/fWv5Y9ibB4Olohl5oMTUF8lWYmSHcyqZ8ksKLzRMscUBXf
AKRxFlxCUm9RgImyKnvvGQilc78t65mq62CrR8gGe35HzAhsSM0Qf3HTB3Q9eddr
XjpVswQfDd1qNfpRXAvLgIE9DzN0Ye7Xl+Jt7RHUWi3FX/joU+fD32dRBE0QYxle
Bx8tQQk+HddIZm6S5eLqsvHfkPq+aPnkDW1sN2aQJ06CFq4U4/pxLLYbu8opLENW
aPnQ/tbOCsshwKlfoxOpWsrXLGfQL4uByWfB/S1AizcPj1qHKD/cO7RADW+4QsVX
XqMkBfpkAbVa+JJXoXya5+2pWvXwrfpShlCTN4yrNjPphKBJzKygugehXM0AYnZZ
M6uOBevuWQbq1zOtZVktu4j22ZCYtSr7rHpjIA25+8PcIKzIJzQzVuaJUkDFQm76
Lfg/H6d8hnH76NbIXpou16+6GgZF421Mdtcd/CLliM//Y4keHd787qVFJxms5+J6
42g/9C7t6Y3DV7XiRk0GkjFJ1bYVFINOfnB9X98a6rVQcmctLvx7Ti8jwBw78wNL
+UXONF56QUK4dMwfwik1yFoQk4tYg6kQuYlfte/1G7tCvmlAxV7XDmakNFTeikOc
5/EDtxqnaOFkfu0a+uvaxSW74V5A5J/1jKW+xzCdxJHs7UvEB5fqyU27iFBaQxla
`protect END_PROTECTED
