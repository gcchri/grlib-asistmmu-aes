`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rmPXcbPYRPtTRqejN1uU0eJ4xcuuUZGeLJP3rbciPBe4N6BbOsyI8guMbxSZa/yO
nK4dt0wcq7oXs1aOplhdhQ2iO//p7pK5bd7NGhN1lei21+/Um7DBae3X0a+aT9kv
hMAff6JQilYAiWhnIjqEEStXWehf6oh4iPoCUfgLxt2UFEApOKxhE1qFrbIBSt/Q
pk/6YTAEQcwnakDDkQzB8Rp9poWqxaV3Wus322n3ZDRVi0AFyO35LpCTAynsz6VB
pbmTMS6XGsMtDAud/T8r4Q==
`protect END_PROTECTED
