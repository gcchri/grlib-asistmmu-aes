`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vpGWXP2+DlcKD3chOeEsX6gvNTHl+EgIhym4p34NuhPk9F1WK8s7CpDJ5XlwfN1Z
mdsB9NneifHw6HAx7o4gd/JyEc8njfRUNdhYbcwjEetrezBG4zTuXo5lEIdkqjvx
VUea3Xa+5Ruluw/JEkuaD9Up5KVZLXJyfGW84Pix2V8GNTT5iysKHeF+p2iZ4651
aiAYRQw5hjELHc0hzhu9dk09+WC3sk4q4d+zs8YMLNEEm82XAQF1fZwfHdS41R8t
Nm2zZDxBrwhpt8pkDnXDKRg2lGem2EsvmjsHBUNvUCs=
`protect END_PROTECTED
