`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CjUx3ngWrMN3RupIgKfZQEQpAQZXQu1BaadjC1yVF5g7zWjCQmv1Yp36baCVlk93
YRCFR6vzXWWuI5qDwxxJjUzcG+FKoFjK0pmVBOJcq7plqPQwf1r1wgQ+g6O/z7LA
nkiRkbbY2kSd7pVreyj1tOhtVQzvDFtmMlm5b3v0wcAQonI00PpwMcW6dKYyBJj8
gEVAMT0kq9KfbK4nwcqQHHbZVc+Acc5DNfvip5Mai+OrkQxlZw1MjAEwH+2/La9B
mMLlQWT+E2ZMt1hnImi6wofBnCEiYLLQyTemtn7IsLc/q84X5zs2cdhQVnGVhNXo
rOHDJ7PKCYCaeeA3ap+oIaZvtfLXjThzsV2eCM22kOW1Clb0M0yp/eFu74KAxp3c
SgaDfJI6s1q30FzA6K2PA2zUUTWI50QhsRO/AtAge7URu9ly01RyfWkpMBovF6a8
aSK7p/HTZPF21MEC9+zx4rHkMoF+OYXrfuYM6CemnXwvYx4tuOJ+B/Y+tpkom1r4
`protect END_PROTECTED
