`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jM6XiHaT/xM4dWgX2uSR6k3DioCdAft4bN1YiR+e1bT0/JWCf0cYGh0/YETLYOjx
cX4/xBaqQ3JmMDgTXRR1dfZXiIm8pxavIHggqSkniT0Xxvl/f37w2FLLX+yPtZxw
3EOeDumGOEI6GkNcy1yWlzqSzHMp7VC4pB6pupBa7+ZIQ9w+YHSfel3Z0WzhmnJ1
m6BWaIXJZF57E6XCA6IUgG54ebdfE6Ubj63OnXknPLZGMM1UwaTTDsZ+Wc7TrVZp
0SuK+5pQQvrsO9HJjtBBD2Z53VQo5OY8KKiX+XUWBl9siyLkXjuw8MFozNgoEOXI
eczmsOHZ6M5S1vIkMx2W806rwPyc5/w+SysGAgofr5votZ0S/2UPszBDaPRof3K9
Jj7Hr/0oYdzADRhKsqwNQPCJXEkefxh7hJDXlB9iARCxcBVk+Fu4f4IGKaHkQqj0
mKv9vlAhYioTIZQQx/Oznw==
`protect END_PROTECTED
