`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ch8OVVpuk4W6VefjDXaFZkuLjpoZ10hpG3iYG0V5wkr+h223PfEGWGQ4O6GzzB+K
p7KoYgX4m0POVohfenmIfWMLLgNSCKrfhnfMqlQGzk2Jyo5b7+9fZrCTibghyBZx
RrCZEr6kVtNym2sVGAtFJJ96xQh+lP27+4fYXHaz7UyMHIW5WXmveYjLGVqFEvBJ
A18vcj8Un0R6ZhAoRdw75d5emDQXbXlfg9hFEdPBk0KP1/N4WvG+oF+vfWRoPRDQ
i48Jf1tbjgHSkgf3tY5aDe2g1AG5EDAs/db7apFqGYTSQnVJbJLRNl7YVOT/ABHr
TL+AxMkmvFfb6aM2ZM+yaM7o3j1iuCqh3JwN6WmT8sqB4NRjZgo2LiXl1cHT6GC1
nPezMO4b+IwwcDGUEEoPqCkwcV50PqCp55CyY9owNmnfRNDuTjuK96+hou6SIMVk
jYYceXGVTkil1dwY2NXxpZqbjh/ceRLsHL50zAiVbC6N4vy9gcp/mgSR2Sf67J7Z
h+iTWFVnrHkkaEvheYF9PtNxMUucbelc0gaKBifQRBZG1uL1wqKerwY/yrOHvdMd
gpH8h56S5OUyNVFgcme4hxmYw+ZRrXUX1ib6U9oCwp0lLte6+7lv58QSrOP71B3o
g+TRvg/NeAafwIiomTR2YA==
`protect END_PROTECTED
