`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CcnVrQEGu2iUYtBOoxeN17BbLMKOI+rUvZbcozn51CtnJXL0uZ0Hr0tZBsYPnk7e
RRYUmwkG6LHobq2NjaEiJ0Fu6YWczfdQdXNhsoWOC+MyNxxq49IYCfOOpAZJ+62f
FpANaHH581UuC6qjHIHOXgn7tKnORUuj1v69SF8Z4X2AdtYJ/hFg9bjnxJKGrGBq
295ouM9rL7T6hG9cId40hNm5YG3UymlLebHJ+KTPVzlCOS6RNBB5X197qql1zvRM
tFIBRkM8oxb3cf97TN+XpBhXrJghJ8tcg083oQ7f37E=
`protect END_PROTECTED
