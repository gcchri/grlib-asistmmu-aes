`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IxoAX5YaO3osFTH/Wa+t3Fy4bMsZFVJHZRV6aihEC70MQjkcyj+FCTUxNCV9rl+f
pBbM8bLn6ESSYOl5Kdz9VqgIsi6kCCvJVcvEnFEuVDmZdAVgywb50on+9vWsPLIB
yOpdl3HwGEcnbxXJjCDpe+0NOGwd0I8LOcN9w+4ecdoRWQTNj3d2amB21q8CTskl
ZKO4NfC7US+AFitMs5XnGk7l7OHUgPhwtmbDVund7I1awk4Sze72p0QZxHCjRRbh
WYnYCR2r/wRLrNoO5ww9o36q+Lk+Aaq83hocw0TGRIYU78+JNC2jG/KlVdMj/jpm
EtGUcMvG0gz3VcGUlPnqLttHkV/N/0DyKuqJhjFcqiwTt4CCOUNktjJunpR3hHIM
nRf7jMVgFE38TTXiz0mdxjEIFl36eRNJzjYJy4kKaVNRW/Xq++pp5hgxfjiOxfm8
uK7pi2RqqHVxGkYezP/XTDK32tLSMYUGQtJADAeF/Tg84QrwBHxz5hJQUiBsym2n
az+7nmKa2CV8bPkzMd2FMgqFR+tqFtpOUE7TTo7bVXXnw3p7OblvR3SLyyEYiObX
CdnfdC9nHmzS2nF2h3Sqd3zvQPyEfomfZRi5YbzMtERUDcO1nnERFz9zu9nnH0vk
mTWY2me+OHO/LpOj6xOeQKj1N9y1MpnB+vO9pKMSFpMcLmfMQ1JuX4W7OoKhPwVe
z3gceG07R/Cos5vUmxp3nh1WnaYHWqPCmCnhdEYlw3es5HNHwldW+NZH8npqEouV
ERCMJQWOE4RNWm+7vlH+n5Z8MyI8rXd8nzMeNEOuDKfXRA+WC0hrZx2mP2Uwiiyy
7U0JRX2kH6rufk731R3amXW2uBFWQIHzDQRPf8bbPbJ5Y4dpuUBi4HgXLTUGTHNx
xNupf/aBlBSXfbKjQ5a+BQgd/rca/vLuB1BGm8gDCHfJrKXOBai+wpQshloG0EBz
DSrTHIBKwhFNmUQaLDPkM+z9otJSRLNvP7Awo6vFYp67Q58LHGzmN0ucPR0XNIfv
0HKkyvkpeatt5wv/Fhf5pkHpCotjDX9WpJQvYgy3RfD1EtykvSfbJ8cZtfDKkK6M
QGOTIf+ahoB/CtBhjFCxOKIKGgFguR9M3cRQQsHgB4aaRqAdOPIDhGx/l/CBQEq5
O/IqOET3Ta+ykrHK9VCkmojFcCCNiklBN38Run0PiunBSXCFZlO2c0R+IfuJoTaX
IkxHFK0S4K25EU9Z0ZFjQ1GLLaeHNIpgu6SfeejYnS0vj8xiIgpP0w29KoLSDMHT
skdssB1m1y9m8688psKBT6LKsGLK+52UpCNf3NyLkNWlFOFbHtfdbPGO6AWKs6pV
Rikbg4bhBaE9oO8uWIhKYEcVMaI/6g6M63wXJEajN2Q7eCI0bBXnr82QVzIoLcBC
Fl0Fj+vJJ/c7bfrNuHHWfYPfnjkt0pJb/Tx7PfSKrHCVv6lfowsi3iTCdxYtZjYf
ga2AVCqGCTob/RqGx36DTJxZ9vmQv+sQHl3Rx0NpVxzEjvbHoFmuGrDTDLmASp/Y
cBE+Ueez3/GHu4fOmHha9Cs6c2Jxyl1hN6k2PMkDEDnHp24bnZOSJiSsss8Se1Br
W/iCpQpWcevfEknuK5BnUPz6iul83uDeEwYNzkHHKgWjmIyLz6t8d47YrUYBXpvo
aawr00sXDnztz+9F4yYUb84SXvhrYLRu5gPcI3rY1WR/CT085LaC/qhQ7kam8LIJ
LjjZGdSqC+jHvjZBS8tiz5ZwTBEVhpnoQWdGU6jwHv0mmfHE0OZ4H9kpbtuQzoVK
cySVSaTT+smmAStMX8aT1kS/XTn3dimn9XjMsFHpURh16MbhwNHB5cI7YIh/eT6y
vUXwPW7GgBzTBXcKFoDRfJ/QIBFtIYekaa9lhRjDOmBFzrq3PTlJNuyJoZvDZpF+
XTPMoN3yy1uGzcguJrkzPhpvQHlm1GtF/Xe39rmCskz3JKp6x1kjSec54o7VQnaC
vAp9dfpZsKouOuzcl+LzmoE7kjramhYeByYXUh+rztF7yU1U8bFYbhfjG2aEFhRT
biznnzYA5jWxNHnYl6h8SfPWuG9QoWMCrrGgfddHWWmx53oU9C2eXlEv87MOPmVt
lJjPGoZjOJemlNLSXsyW/gGiMKYTFM8lEhDUvTmB4gTmTFPlN4Jv1AIuOQQtjNlM
ah3f0eSBxso91mTi5YzHPSFy+Eyvy+ntbRniB93QcRkmu1c2O6Uap1/dgeqVuFCF
Z83AbDLogZtx1SRrZlJXdPYgyFz9xky/elC6skgTbutDUOO754oVjSfSqrbtpKzw
UbODvxFhpcDHZKgYG5bkOX4FzNMZBrrGwF8n3htrMX4y3IpRoLpWSpyNDeXxTbxH
swA4yNePFZU6hSjlbPMm4hNQ9YWRUUNhnhJZY4+jxmO2yiqy19xihh5AH4auXC3L
ieQLC8qtU/VozjJGOQBLdY8w9IqBlyWr+AXCrPKC9JLVjXd5PmeiwoV/JIcFBeYL
3Fm8+y3Osdm89qRaHWH8hIjNJUVq1TucLLE8YzG9D7O+DKzb2rUDwb8dcpkds7Nt
ETRb5ZASIWiZBkoeXpfJ0MaMKMS1QKGRiDYs25ZoKu7ZjAHz+tS7FBF11DAIAwcQ
Ob+t8Kst6OLkP6gBYgOCZahK2XA7Z6TjjYZBzQ8/65c4pY3CjeIbP6kOAHTnTnrV
hxVshb/DB53VWNSUtggv9VOvofaTYeEq0ZLD3WeEGGzJGqVSOUXBM1tViH3qd6Xi
846CV6NlichI3v4vA7Rf9NBKklMfwSlEckEq15KuR3bWEptkbc3Gd4rSuK7xfJA3
NsD2S02nibxvmxpsGidQ140KP+AtyK2vO+8Nug9/TdWPVrVDAllzMWl+IBen5vKl
EDG7ZETQabw9HYL8nemDgPabfKTnuvIBlX2CgzknmTKJ6HFvKwi3lXUVdImKWohl
Hg/fjnpNq7l5d+SQFZYCYHNkUHjljuX7U/HcYucgkTp9u0+PUjQy1POBaID184LY
5DNzTFLosxNJEeN0acR19iSm7evj3loPxEzmAKfuNkg978FwpO7ak5aXjvMZDzm4
Rn8+RNn+bTLUQb5JRyFZiJkJv2jAAzEgFVkDE+GIwUxxVLQW8XkHvzU5azXlTfmL
fAWvPM0kbKHUH54WM7lmmQ==
`protect END_PROTECTED
