`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vYeBO3fPlgGR938HdFacwwvBFp/MTYid/dynx8LZqdYLdfi8+K2M0FdoAl/TZ687
5MGtwiN9M819wgu51PM0fXksaLKC//ZtPk1fxJJfzWCVxhKcAwjC748NIQx/OnmH
uc5ugaqhIjfbWi7mOJ2K0fo5GCC93MAGPLoAd6YreRLdL7pPi23puAv6sQ7E/ou9
z698RtzCBHiF6iXJIr0/vPM1UPYNkRT+taNuJ+DsNRbZEEkcWIEHWTvR+dYMGtGx
BdphQQWXZtTTDo/cXjKlDZyh/LjWyfGIrdOv3zr/xfEl9Hr54N+P+EdT6ddUo50x
2FBYQX4RIz7U73jjnlOqyNkpNwAxUcU94vKB2ZuT187zqicjbm20Ist8fPwXWqLN
`protect END_PROTECTED
