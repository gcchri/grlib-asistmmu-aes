`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YP7LSHNCt2w6/zLis7UGeqpd4KMbeaX70QV8V5Y4CNYVXOFB+4BMgT5YUSbSXlou
rmRnUv5KQRxMt3gv9ozsfx/kq/YA8rUxRjaqZVpTOOMXG7G0tlZnt2i4Q+U2yPHB
C8C2EkRsDK09QZr3qdR1j57ZDo9B3ugg1rIEy0WhTPI/zmqBk6NF+EhqgaIOAyzK
XBEBbgN9CIlN/eJ2g1i1wo1QJIsdWXKdwgq8YjhR2Xp76L53khUTX2tIzoVAAWvN
ufnO63HFuIFs5l+TYpLk+hAeQSNlldyJN09Lci6h/DscX74LSXj/q6nJ9d4bmoLU
sZgrbkG04UaojmF56dXXSP1p2QKDkorDHX8n7ShkDt6CX1vCsqzwiKHJmwazLuVO
mjG0kYbalF2OMrsoJUS38uVMcO6WqsP285iaLlcCvAU=
`protect END_PROTECTED
