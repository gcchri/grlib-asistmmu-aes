`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c5Id9kRlK3I1ERii8y0CiCsZ2VEuZo4NEAMilpya7k1q+XUSaKOBolFBr5fRzbws
5vq58aGShpsfNTxXmKu2LP2SmCXYHURlXGcK62otBLzQyt/9kj0M8lewvZv4iYQr
OB5Ba/peqXOiVOwmbTwLEgqBDTl84pikNMAeq/ZEZ8tuSZFKnyMV9u1v4RWkW/ra
lHIO/bkxOBcI0RJGfFvNSZ+wj+zVZx8bu9cjNl2eWFvw0++LO7x1g5xUZxqD7SNn
d9Ytfo2sYcRmhs4KYZy0EQ==
`protect END_PROTECTED
