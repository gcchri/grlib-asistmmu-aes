`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X+zro3uXzZkJT0hpjWtdypBYItjq+SBygeFGVAY0sE9H7Klu/M8HD5zk6kl7pUh0
g7eebh5cH3fQUZQa2AxUp+81UExUE3mek9xBmg6KH34GEplpkeCyF4tWHA3c8Ai4
89Lo24XhP2/OUzMeRfDUAvVHDjH8S/yqK32v356mieTdeXg1l5daXT6ZswyQPx+B
S13pHSCYSDvpWcqhxCPdqHJWrQYtDX18dUWcwqcOfnPzNypqsSU/BSnEFiAnv577
aecVQzBf3Gxam+c/0rxrRLt3MfbQsMCCUEz7MdLltmvnPl5pKCxfOey/FEeHgil4
c6Al1JW5qtZe+ivFWzsyZWfTG20w33b/qvTNhb8auNjtwp4lNu85KyQTNnhCZDP+
caRS6QQWNq+d6KbIl9NJwEspVTSAUwRYTZ3Ruwos47mHWYYo3GMDtg4gGZ6IxIc0
Mz0Ze+Cx83BVriUH2ZnZyilx+1U8eDNEgySATuVj3ZL8WLa8IcB1TFglHbGFfJtH
Sy2CxLg0siPQ7OnAg8/WsEIy1IN5ySamxfdAtdT7Hwo=
`protect END_PROTECTED
