`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dzYB6mu03kBFjEZMyRhzQLlG3orqgIgz5VxMxoS5NpxeYEMsMPmlUddPOPhtKB8/
iW4Gy5li2983zfoL50qX30kn+N/LJ7HexR7UWcODDRHfnVNsqN5dWYjG+HP5BW9/
PqfIlXi5mWFG1/epBrpCPU3BqQxQyWWI5VeD268A9JAGcl0DKJo/9QZKMB4dLXjX
U+5nwuCRZZHkxhv9VBhv7JY45LL0cB9mJvlKtpWLmzFiYNkzyBpbQjz9DCIYDHvd
+8LhWtC3V3jFrcqaK7H9SplXWlKwFc3W7YsFV90GTm1GZ9Lb+ofYHqp9imYKQjcy
TYIEaoKWW+hYXX4eFBp0rKvb6NNLgbIHmjncLlp5sitR/Agn42ugjwMGcs9Zk46+
`protect END_PROTECTED
