`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HUM9BH63cUUpSkehRSDIviJCrOU/HzYsBxr3DqhSV5lzaPke81hctFNOncg3C1M6
/j+KVkeUYQC80zFY27gn14MOttADLUQ1u/1ysCllMp1aV3U+8ZbfOKnRD7VDIiYM
3xkytLScUi7RalUUgLiUFA4TW/kK2x4OgwJnQ5/fHmJ0RZeIBXBxGeGo29SuiVSQ
vWqJKgy54nsOxY/gB3Kqbuje+/weYAGfsBe1cEgP7GPS/TdPkoHr05Cvi1zGlN9p
ms2mBt1DPYBSCIlgzWvEeU7tag/bLH7jqLJGqgJ5Isd4Vt3C1LUFzcFb2T2+rT8d
Imh/tHoHiJcySFV6ZJ5bhy7EhA/fr9GSzWQcbADq9dgu3xF1ZB43ghJiUU49bDE9
146T+J+MrUEnixVmZzf1SYUKW3CCJmWJhHwV/DTbp1tN2eLIBVEri5UqgtTcx2Tn
IPmUDF68YrKO6gPPPPf8uPrZsEx4HnWQIVgwNDUnkQgld6ksx3kkJAFtmnZ2jNmc
2q9n21S5xAguvSwX5RZdJ/JZTkhi/6UVwXCCLspDkk1n9VUn0KeqcvGrA9U+zTjn
sZXJO0i9bLQs877e9bAX9Vt+jXlisrf0GMU2SMfF75kmBCt1IG3M65ONYvSDJcmR
u9tEst7wk54LcSw7bb7MaxAjXKp8BOpPfv8mXPo+e/xlmwaSGjnOkRRIWHx8BTsg
4HNNY+iD1RCkmkXV/DxuQdGrkx11s9UmvHgwJtC03HfyRQP0LDzCN1ak5QtcjGAy
GFWGpwJUwumeDY20uGVFVw8neHtJXHfTR8+ZeF6lqT2Ex/s1fFWGVm1tFHPUPb0P
anVwalFHNmO1hr6q9ssGk36BbUbj+IwQGLm8iEk5pbaODiyLvi+7fAqUFKuGDnli
rjDy28rCwsadnBIlO8SJC+cYP68tQ5infvzYMDzp2E1ImrPbwzuO7GkOeRDvkD2p
ndxNrR22vctRwTc8C+G7gTg+u/3B62+hl/tJY5AZZjVDhIHJOrvRdl1lFoa0LeR2
R4I7Bmv2Cvh2f1g7IDcnTKZUJhQvMElzOfei0w44Zg/mtQ/0y7BJ2/c1y6nNgJxb
2ZwLXoUcbTDr/o84vjz9VEQvMfxZdoxmLFA6fCrrDfl78jvnf0oF2Xz++NeYpb9p
`protect END_PROTECTED
