`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Wx19rayAbXDllSI/GvqaZKRZAStKmG/5QKhXWpyLwXqTu+5UQ4UMglo20QN1jFy
OKQ2LeUzTAPD4UG4SHFu8gw6Y74b/5X2bS3KYTscm84OpQFXAYbMRgfuqvyk3+nP
76WVcNbS0EZDw+cOL+i8BUkDDM3vEcDT+MAAICIy9DD/Gw7P/UFK6F9cLxHULJOl
6J4aEbaJgO9fdaSfvVO9S+Z+7AINe5NjHU32FaPsi7UXrB+E4vKSGRDNQ4d8D1UJ
`protect END_PROTECTED
