`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i8theiB8DtU87EpFGlae0/5eM0HhuD6zOZtGb6iV3Bu3Nndb+eo6UvhVJ4+GbEpc
pv17L5QikBRrhcLlzZ/TTXFSi7Yw7qvSrgqgeapPqIxuMiQ0NaJfefSYvp3C7m5S
Os+4YLb9yr+uOnCRQz3zy8sc2HVC6mlEC3EYCk4SRGodlm4Tmbak14WPLFfVJVf/
EDspMEdRGz0AshuWdjAPHGibpq4a0XbEO0TDHERXFu+gTGP4qQu7fLTwr3SjKQr2
gYJo+6vPJgSR3UmGq9Qr4uWl9HnlfLdpiQpWbamRJAzWVbq7f+McRXjj0O61klYR
UNiw501TsIZtf6FukxtkzQFV65CEeafH/w9kQh6si1um8ffOdx5p03e5ONaaATCG
LVpdWGX4s9/aXRvQIxWcTgojj7MrmHGifet+iwHgN8ka2Zd+rmlTFVMJPS3p7NkH
RHHFwPr7IUdsuVMbYnL0ao5IZgpSuwdqmDVVWRewij5PEGJif18m1CB/JlTds8hg
nzdrVj9V01EkYQpw4nCE0scH6YeWWgQMI4iMKwsaMoNMlDHgim9sDvZCEEjLoG6J
zz6E7D2rMnm9sAL83FrqBYSGCSqGI8k32YhQI8fzsWYoKtYCFTPvpX5mE6Ri0Y2z
EzPRgGgr6pRBgAO7Seasp5+Q12sRsd+lhu1PFPH+1yYgnAYld7/stZCxUXUbqwKA
vsVHiWfV3v011k+CLMIaEizG2N5OPunJ9SqmfXJByUtqrTGvrfxB3ObeH7cFvyYg
+Mo+RLRwdwJ9G5z8XPrl4A==
`protect END_PROTECTED
