`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4yKYzfZkyeM6cWeIO5rcZWNkkLPDukmHSo078Aufe1U09DqZDZstOEXUyydgqpUX
8KogdumaEaWxOjO9JHFoQR/ZCCI2UGj9118imGiX1S1BLBtpb4aYLi1sGL/QHe6M
imZ6dUp434E2UA1ehQtE8uRQTPYXqJvT3e2jTltpnr/wKexjxASRO6hnJS6wquV7
o6tT8hZK5SkZ8kPSY/hYOLvrvSBGyjge9hM3zzJyt/zSSOzkWMUzxsb0RKNt9AM4
cpupHKhSjH628wNaDaAEriWTyuLuOKwGK8K7BqBz8IGBUlGCNhCzMD6NBjnQvIBN
xhRRGLYqxtkQMnKgFFLwa+hizJQVdG/TfBbrHqH3mmapgJoDNLagOjmaUhmj86x0
gvcUWkoeUz3SIaOB9jeQpyDQX6PXGeH9Fnp6XqZP48hZMp+eXeg/Lq0PkkXE82Pk
X+KfEYTsKVXVEns4yu0zv+xJLO+T9eKZlJiRPz23taQ+rZoIspRov07cV0xxX2Am
f9bv4jAGMUGE9Mo58gvohqJF+LPZuVBqsqJ0SW1rKU8KJSu3G/xHOCqumCcEDZtL
TA4E3y08eP0x6+mZj61AuY2v8351yuxHVbA7IOAHxwobiVeRTWYWHXnQh/1JVE9E
CrzXBW+jRSY6baf8UzCSxilh4zWsNYgkZ2B1fW0K94jQxlaWWQke5w67yaQ19Du7
`protect END_PROTECTED
