`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kn0Kon4pleqmKlXKuHgDiE3XTsz//viEd94R3PVtvPjL1ezTXhmn9zM2DYvBVMs1
bHD7e6oqE1adnGbYI1sMSKa4dHKtMct8o7I0WWBJUtoWLvYyjKQTVwW2DI9/GpoF
aAx3mBiJM+iHWAqJ5MMiOphVDh4ghEnrgN2lH0zrT72N9Cb/WtzBRx2S8DLyutYv
wukVeQ2HoaGAVpN/YhpKqQhLY24C0wQ5HsWMxIVDc0VHv6dFz5Mzo6+08ey5HB9A
pLzAYGOw/a9Nk9S2PI+uZfLSbWkuydqWSFPUbNGKF175clSVBtRENOSQ43xYtJrS
Un56CKaWBpNxdmHaxPBuFN3mrtMk9I483R03bb1OdPvIrqmANqcMwL3+ah8aybCy
tC4cVGCI6M+ffrUzw89ugymtHjnb9IUBJzmP8qjGD9u/mh35h47nzV/fu983xreP
mRU/j6r30UhZ0+5YbfiGp+BRIP2n1B3qGKte+uOKBdH0vvma3M/RH+6ewEqSLlIz
qSQ4Nw1y24T9sBepBEnLuK6pbI6UBDBCe5vM/X4xS2Pv34LUAUqfnMCVy6y3UD+G
8/S3PcLT2pgYgYw42suTAIfBT2n71ttdfSJ5ijR3AkHsTbYb5uwNcxYMJKwCT3bE
PNjHprPS7jV88G9hjJS/zShsGXiUm9z4Dm+Zoy9z/mlGBXbIltUTQTK4pcgKzkh8
vVkx+aPTtMZu+McHFf0N5ZfzOOJwH6aErCQj/PY2PRuJdLHkjfm++K4Vbvi5HuAH
FVc/JlDjrhzaHnILxVX7rj77UzFgfyg9a5O4lTyHdXKtKhUmRD7wo1kzfTGmtwu/
s54YYj6iTt2RwWIcQr7D0sA+MI4BQy+XKxYfNHE3iWs5yC5Go3YsBJJdwsVf900d
E3DW8WyqwiMpuQS5etCofuhhnmTVBnoLDJ+PRBJ7xfS7JIaD0spDxzM1hNx7Sp8W
JQx2Sjty0i0/3nQB7ufTi/YLhpIvwDdGZWTFUFQBCcdRrXzNAEaOu24bk9oMnzuL
iU2DcTFHuMD36qAKzrxSsT1x9ALa1NnoRZjoutdWYSzjGBZVJ6gslJil3FDQ0Dk/
ir9qQv0KOpQ9Ohql6yn5nsJGM6TbSLDHn+4F1jh2vYwbXoBAJD6O671+S8i/zZR3
vBuO/1PanfGY8DLV4LjM8t2HxQ/gSZw3TFxGL6gEiPvCYElTQjSgCBEVyET2LUel
ur8jl2leEv/KZODE3PdXkexdKLPVyP5w7qmjGXXlhPk/2Gy0ceHwhZeD+sdXaGs+
zaHilsosS1KtoUAiGQCRjAQOjygi7sR+prMIGUpbJCuB9fczbYo7M17uP69Nhc25
CYhIy5VTlxtrIAi1Xtlel+iJUwxbcHwD4dsEk6I86bZz0tCY4YNJ5Zu3Ro2n8kyK
swxgd8qb5MdgaCE1gfoeKxsedT9gPtGNQ5OZH8lS9cilshJUqFYTVntshljNjQ4f
Qg5NhCH4Hob1HtHOctwvSRW4LouX4L+jWxypEOziWrzWfX99BNOWLxM+XoYMkRGN
xAi6XVi500EvvtylV9Gcl1/KnCdIknnLzb4ZXhL/usIkpFZr9zCdU3/AQPpOhPrd
dnyzE3IHTyecOvZAICx4Myvp3oBnFeuSX9vsZOQbflXl8UD8gDJc4AOdTt6k1kx2
MgVtS5d1vjdRdF0aqxwFkO+8Nhw/yIEyZNguB/e5NcMhTyx6rO1V9aY5UTaUtBV/
3OuOeqddCDOg6ZHyvntmLb1ZppE4F23SGewNejPF2+PyaaGKNOkd7VmtOmLgjy3l
KWIoGtOCTFi5zlyHoglKpEo2mzBJ8ZknysClOgl0OmpZ7KCKu1twzuucbLvUSaUO
VVH49+SKfny3qIIaGs+YKVr2Z2DgLg6bn3irHyR8SfBT961vG3xLMQ3ltMJT5QUf
enfo4a4o80Gdbw0ATeO/A4Qxv1EfwqZ7clVYFMlTGIfx8FT8Avs9MyF5o+NosMwf
4ZFTo+3E1YUbMsYDeLVMtqunWS1najWRP26e9LoS3ZbkpQgq0WB5PnI+TkYYrOzl
8xfodg/tHrzV+xB91oc8QsuaEvo9pP19ojLX/WGgp53yh2iQxWMNfeS59qKA7OZy
3MC9ZHndl0XyMFkU3nDSi8fe9vu0hw8vvYxZ4fIEmcy5//iGtYzVjnI6gYwU4T9l
XrHvgdsr2ka9mD6j/ZTY1vn55LT7trEI1UeulwWoJ+GvKSvVhdu/yENLnyHDF6t7
KHD28kFek5LcyWDmQw/jpCXS3OQjXoXNffVl5EGdinajN00bUMgwHUZJFVjzu4Xh
ykG6WQZRhz6vr0058Zd2xedNjN2ZHJ+szhZrSFow9vajeNayrq6EFmG/oCk/4Ijy
DDVh5uUiD5secxBZQSy5tFnz/ITV7y1Y1QGsX+SRzTmBliykgj4tpvzuMgORAIV8
0Tcm+yHbK28bU2oyr91spJWIpWDkNzNXo4BCvupRQs/fxZP5DInSxUfCpYAYSq1P
Kucp/MOlzGdoQi5U+5XxD3Zl2gRyqrXPy2PjUFxKtuKPGSDGYUUOzkz4RZR7LLPX
L0TkV/EvuyJJeWPLshaLOjXgzTzgK0kaKQlO5xiMnAd9MWFPRtB7qZZDfkd3TVV0
dEL2KrOg6nbmf6jAjMz44fnPQ1GVqU2jzY8ZYtEw1a3bKsmY+dYfi4lm0q/jARyP
bLfjw0ijwSTcLTrlrVxc+G82eeZnooK947HxYUP21jrvW9u9IxzDlDnhH/0U9Ghg
THxuDKw8Og7B0JHoLj4Qp8D3jb6qEtMuQx4qiPlx7EjdawCTAVI9htJHwMpg3zjL
cN7+m4CKVirqDOOWzy+Bbsje1z6IR1eOEPCF//h273T0UAIeCef0S1j6nnSy8/Ud
PAzLv0nA2MT10gAHvCujArgQbTIgQUzCGQgta7hWNTNxAtC2BHehcqci0kIYzCJV
WQUkpPhjgxshNHlY9dzYQNHv6utxL2Eil8hPwsMOBL9O0113kKIyGdtJTtB7dsOr
0bMoDIif6GsmuxGDQAHADXr6RXRvX6xQlZs+fJZzHmnpJa24YFRGGGZMOkVroOvD
mvajNeLp1K9y8t/Xg1JR2S9cgXBZhV6gpaRO5z3AvfUQiFkx7EV/ima/2RDVUQaL
t9hN9QA02GyyzLRwvqaYRwZ18/BnvfrZJMaElclElZGFYmLZ7OrSoM5mx2UvuM8d
4ZUqsNF5FWj5S5i74IllBwpWsaSbU4Lmhf42ziwTaFcypz2csSe4K74nc+WYPuKY
w9jLNoPVSwijhG6zaAVvQ+8jC2jR6gAbkWuhI5W7umhG8lqlwtsUg36X/yRewT9d
v9yzqjJ6GRCGKhG8XVAhfKh9ntkLSOAYlQzBafABLfveAX+KtyqHctiX+nFizEOB
TFvcC/gI/NJSzGIahnkLkRN+MRhskHA16EpYKy1INDj5jwSrBP1xMiska4MT9pW8
AfLqbvSC8CS5tDz1qSZkIGLnlz/P7oiEI/r1C+yavCIvGSfZrYYIbpC9+qLG2e6u
5gQh/7XKucF6fBYe5P990iW0eifj/yPi/CkKvCr9AdF1WEJrukVsCk/UY9UdmJYd
J/O1xIIFcx1aYzpmmOq9p1HI3gjd8qwH3kJN29WBUNuCvGUsgUOmz+p+RiZsDCN9
xTkAMqJ2+5OV4/RVTAVe5GB2MrTZmfucOABJQDmXPK7os9E/BTEKrzE3CXTI6GJa
dqfNtoGk9gy6ETfvYfpYQIoQZ308Eh7ga0grm8QyQFcgGP7wLv6fTQ7zfJeyP3JL
YoNO8HntO1cedLrgvGcMYfN6Me2fwtn2KmNxlgtIvzkkF0WfgB2n1XJDSAN5rWq5
FyjYi5uqMOudkTzG8ZnfEa8qhO23uYIkGn7szYdVi8XKMnyvZ69WlNDNp2p9MmTT
ppMP5QtRHkJsb08NtTo808DXWDDfTBgkaZK0VKBwb3q9tq9R0xZ8Mk7QEcq7mbXT
Mj32L83aAb2hLEbAyBp+vcbFRQXCHvg2cTxm4jOhVE70lCWlwpNjbLqy+AWi6h++
ogflMd0XEGaGNAnqs5VcO0Ry1nvCF0M2dPWd+ou2k/96CPDr5M7I/1vKy+ntTNss
idAgvyMHCmrEH566BKvOyg==
`protect END_PROTECTED
