`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
shapow5WqJo0VhB4ORNXpAOijJc+ODFTqYGRTQE7M5xJIaIecEX88YifaoG7HlOV
9pdFRSEfvEdS/0c+VJXlMFfZfN59iN3oToDSbvO4RxaerFNjHz2SBX1fzd8/0aBK
5e5YbC0PXpYqSBt6t0KZ9c1oXHXTghLMKX3ttBc9hO5UUgk4fAwYTSn4z/nIx3Vv
rHp09JdGspecbdQoe1CzN8Kyn1WC5Lxgd5X8E/ShMxvl6RUF8npt1NfeXlYPdZMI
ItaQqG4VXxyN53gXnBT5tHPa8q4JnvjyzRZHM+xC+n+Qj1fif5vrwWYbUPK/Lawm
vIeJ4lDGGdlCgEkzqnhdbmWHfXYo4w0XxHEnQaLxMS2sBqR2HsyaTFPKBgHtclcV
i1XJMBI5qoXGwpIA9KJsSts3OsqKoafn6U/WWrX/+HH1IWnvjAUIlWVfezOP3imX
oFUGmH6DwuCNKNcJbB8tUvIYaaXFtqfUTIr/pzEkPlsx68zOyBoBF6oZc4QNvsJs
my7ferc2tTDVuWlqfmT8f8InJOKq9tJPizh1ytFf6uN40AqQkuwaaNqixyhJoupo
r7vrrN3WNC/ipnYg7Zw5+joiVJRxDSxMU0ohvtioLDPW65x2/21G/larey22Chwe
XrMjeDZsNkL2+ZgT5sweVg==
`protect END_PROTECTED
