`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CM9s/9Au5xjiGGzwshDJkwxITM84HQcKxYLgyudIn/TqnrZ3HyCYRRUeI5pc8S7s
MyHq9mF5JWogfPWEd0jD2q/M+QnCjOwwjVXRR3dwiwGB0mkBzX0n/m0o0WfYnR1C
xbqxxIzQgEnFFugNX8y2WtvT93e+TcvpV8iHHWC+vVBh4Qx8khyw+sWTfUTJ9r+j
mh/A/mdQd5VXlmcSURuNs6itFPeDETEpst0Q0o7rgFhOjV4QVLMiygfJBJY9fIJT
YmH3nzUxmPZAzsnGipc5y/nLqweA3DcAMA0JEJs4EV1euq9UhSYEgULFYcHgR4hV
1zHFDRMirgfwWFHX+jkdNWYDrmRdbEilaQQGBUtdblRrShipnk8FXn0D4Q63SBcw
Z/GbtIbEhxCwUFBkFIMXMDrCNdtv8+OwdbdMoA+MqfVOoSLS9zfGWjIXEd7yDBRr
9uD5f5A+bR2vMEBE6AGA80C0AUdjyszVzzMc99U2jU+H5jXqbc3SoOsxHxPoDSdm
CGcPa+7jqtKeojoqQF1ZPOcuAPILNpHuhhaz22onQNMzbKq5EeUIgBRoWhaydCiV
+Hx5wc6wVef/Aws/wIr+4S4hv/CwJjvSkabL4NGo2BY=
`protect END_PROTECTED
