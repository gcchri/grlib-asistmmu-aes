`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4JSo0p04z12W/o/IMtcyCYXKQdnJqUYMpSJukoIwmj7TDoAFMpsWlAIl16xRlUrk
kdXIXurx2jPmAVT7D46TcgJizVJv34wKu1zFw1WVRsm8w/g13R1M4Xodq5fm2PE8
1v74vonAiDf/Ga6yuXij5KGqhQb+q+M1hrvLbwBRVJgVPtHa9N36Oq7GUcp9VcYs
Ebdet1+oMY1VRoPKzB2pWH2a2JAWlq0xJv3fUDDv7F+saWXQplvp2POJgMjsoHJX
/L5fIzmM4zrz7wXqdbKb4ee3wqKYRzKfh0IjGqDI/Izn0M4MMyF5eckqgQjQ5qhl
UhLRFrzJAualEmAXzmNGdZm4j2d9pN+AFxnz2N5PDcR/iB/f51N8NRGdTnWokhm6
u+PF/t2t5S9soywyKSWgQneT3yXdSkiU1a0nOXnR3LhQBLRG/nOArewgiUfFy609
4O9NLVtw6CH6Wdws5fafDEqaRNCLPtZ7dxN+BDpRKNE3EI8cp/25t1Y2dTFhho5q
`protect END_PROTECTED
