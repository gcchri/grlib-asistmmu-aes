`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TPpKVLvcbeZ+eafbIdJrJk8zNteZpbOsk6wKPa5S1ayKlZEESBPHjI1ta6bY8V/j
hRwJjbee1oRncGZYp1NdilSUZbK1MKRdSrOC3A37isIKqSGwCowHjV2mSZOiN6Ay
CQi80beQmpHRD1fvVCUk377oV//7sEnjBeZorR1GPHjlXw65qwVQnYHCXSAbjC2R
vwBQQZS4WUOXb5gq/c3n4SAJlHNHnobzODM6hV5lv2LeBQVwp6Lq0/EbB990WJmE
U7tTwuA2VxiB9ZdohZ4+fT7nFHyKDI4KN5e1OggDMVDelnnW6aZHuxVTS3Eo3k+o
U1gBvPWtNlONwzI3PK4b1MLbKGBb90Nc4c+1qHK4yhHlMflvqXsGbYHTCvxuAgig
fNa1UQ+xJ15GBAG164BTBUBOI/BO3kQwRXt3ZT3Pcq4=
`protect END_PROTECTED
