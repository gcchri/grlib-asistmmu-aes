`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6uo7f6yij7fTr+VPUA1I26A/EYHRhYo4S1TSFbttfiLcsNU4DkMefGkbRDRWu1K0
YhDk1YlFbIA2T31ygJgO+pw/loJUazCCP2s2+vmB7rin/fSqnZS3bE0KFwRKoPDu
EU4HaICdIW612Oxil/4uaprqHckBRN9ecwAijOVaK+mhsfjdLQY8xDDLinG4EiiJ
LbGToUylcbkJPTZ+qiqLWovVo8w4VZ1rLhK2rs/0mbALO8HsXaFr5z2vsThMJrsv
X21NSByEP9iqy2K7K8PQvYdxVIrFsRJiQfmOWRcNWJ9rMmvwRxjeJnM4TTGm/oLh
okQXxtxIV1rlwRFD5U+c368wSmNfKyn0AaMtNI+iGqopbv89rGKgjxA93Rxc22OU
Q1omm7JydZWEPKgdepl3OFTc8TIN1kMFKYDVJJNbAxy9DJqA4CZ0HnSw6+0h6cC+
vbFlES0Qo6PCMAx/9dgtnsU1L1tJefeTZZNUn501x9bP7hi4F4f/fef8LgcbBrjI
jbrQv6yke+ZVNOLISOwlYkLRZ7og9ot3GQKEcqVsBRA9FPutpVUeBPXV9/hyKJkA
C86/0FgZmXtoX66i6yQlpWw06HyQ/1fG3PIBPvmAKquGPqCLvtBzQgEdX2CLTW+5
tnXtlxJb3frZAHGQ7oA5UchFZjS79zE86IyctR+1ZOM=
`protect END_PROTECTED
