`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S/r8AlYGQw2HFp8UvH/edgWOYK6qqYe4DhGNHcoL3U2L3QgfPgzIvJy9hsphtTTz
NSbkJ0TTlMnWYnxNpHbyrcr/rpjBgpLKK87D3CDv6glvZTLsnRGt6qJ1SxMIez8h
DiwzS8phEa5/cUjZZCKeUVtei9t3zAxfHGk14+W7tMCRunTVHYX0nLy80OcN/qmT
yJfIDqlxv6LruBuTr2k3+aDKFPXww1lpbw1ZYKyCGPiJpN2ct3Nt/RYE7oTd19Bj
PMneLaEpBZ5gsEccsvXvuoLWreCQ816x1mhQ3MiYuwcA/mxgQ2CxK8fTn3EbMbfr
mkagGzeTbw/DgszROIOwWmKonyGlICU84WFhKVHiPMAEFYnGf7rUSmMffyIFO3AA
d1u6CjBPkEDDiQuJ2dj6eHUVarLolfddpvxRu6KLPHO9FGX8HO9CMCNffT1KM+s5
ts1Nq9PseYGIxbtlpUM5Gt9V+iRBc9+u93dulN7MKyXbduWZyizHa/csAFffH9zd
ydGNuh226RY9KnE7jR4wFyHqCgxo2dDKDvTYarCwYx+qA/BtyrKa6gMfoscJfUDV
m8HsEvDNSF43+5swV7EadGef2E71aqtxZDiCpiAysFQSGNX3uJezSqUKV/qous2N
JcAHOW1hqi0sJgjNEpF2pIKjOgx2Ggbg+xqEtQA/trgqfhHs1POZ9NbFGUQGWD1T
VmL6KRrsSj6HrFMtWjsiTOA3kX6D4J91QD3uI/zaYBp9yDKPd9cCU4b5kRjvp67f
zCgg2U+8dEbu/dmGvaKZSjOVgTB8R5OJmRebF8tzCAkwius93U+BPARdpmTayhHk
x8AvxqAIOM6xgebqDICRwl4+CJCQWp7knYYvbOtZVxz1cLtslkU/5X70DZFRg76b
QyhAemTIfdL3zZgR291+CLyxDLCswk1e7DDmXdcdObDLxVwaupeyXqgY7HwJwC96
07hpSKh29o0hwpag2UTBTow81zK8PcAqc/PafZ5HwhMTQofb2DBCNPKYrdnQr9Y7
gPaIDAxwfXe//rmXVOfDC3cM+rlEzlnRUcblRFoGr/v21j5MBkIDpBshzdpHIAJQ
c2jS5iTsfxYaeO6iSTIJrQ==
`protect END_PROTECTED
