`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DoC/cbpLo4yBxFLaXryoHZ9QB2bg2tRkF6PvmcOOh0d8hp0cnjt2cMXwet7j0XEn
7S3hUWapWIJq+GiO3T+nF2JnnjgSc4tKQfNiBCXmT9ou1IpYKqpKbhQsCcHtQcel
HuSbsdYYPm6o0ks1u5siCx8Lo18Tw7pj0vHxAokcXKp5Q7LlhGZiWSJe2aWEnIfw
U+mL5tE6vPSVSLBSFpPMdxLMaylsh7u6+rKTFCqUg3gPEthRWk7scOMs9u2T+IbY
ZGd3tuGv2SE2wOr7XD0YBAk7qNj1mprw3rygMgVQ4OIheiOoHDI9HkDc7KSdE30G
Bj/nmjXulbwfN3gutdQZJL19NlyzNUy+lcF7y4vDN0YqvsQ4r+5JGQi+jPV26SgC
C/9pMc7aIO/i7KKGOqriigwplfXniBANRfOIrPrWlioIb9gpr0WROq077ecJgx0U
NMcvyuORrxQKP0YmCtyQ0/zi78zJbi4Ck6kBcGl+m5MC9x5TfRQmKGtFOO6pNLdd
QKMN1Azmpzt/8AUiXqj8h5Asf1RO8dy1VJMUaFMVVwA6+OjEhOzyHFwLlv12P09X
wrwS6TBKjrmhPd+NQkfCQRoa3x5C40itFiB6+Gw9vdh2KIDgYj+bbWJoC1LyISa0
qaiEe7xXvmEOeGNasDAturmxdIBaIsN14gRK8ddc8SCYY6wXmQZNJYEPhS6ygVaS
m5QzW5tm9RwhdZcLMneehqTOGAO0N2vxp8u6LYa4pSGiRNvbMmE0MqQ7awcsy+Kg
St8fIrkJeaHSJVcAW/g1rch9b31ZbDqrlSdV2sIX75uG6GBQGbd2GwAb3J1n2ITY
idlC5uhTmYYwyWBVImuV83Ja4UbedLzN9cWHaO73h+Mxh3kBoVQ+ad5LEyV3TXzQ
mJShAG7CJ/IHbXbB78RI7GtHsL/ZCZftQLIC5pFuZRl69h82FZkTkYZSDNqOjsv9
+qMiaScJYKMprCXNgoxM8J/Lr7Bzh5FOfyczCrzxaxIKYBhSOzvWH/QWOG1aQML5
WXcTNWAa6yyA7KZyL04Cu1PPtZ8QUPy3g3xy8fQWMoh3meRTZDEqU4X2oU5/PBJc
GKq05wOwIimRL5DBMxqKJUPph4oKAw+BoPbhz4lpgYv0eN2WtBbVaprAm19ffRtc
8bjKI9MjaJuB8UFHY+uD7KcDA49GXfKlhcsbV25gK/4BgopL9zSOXgGTBvDbyATd
u2HbVn8rDemLxEcYKqQcBm2kWnfa1IPNnLw6RgdPShJJFC1h1hwbnJdICH6KRKn7
LUyy6G2vTnPqtE//j0LWETZaBBVA/V29X3L69WEGmdXcWB+xxH7fTZx3aa4G57uh
IiZcNaIPrfNgcu5MnCPbbaVj1pH/qfM0chXC7NUYl4m7ABDQ0Ehdtvc6V2geKo9a
g/Zli5EGrq6LO5DUbGr+RHWvPtUGPvpZxH5hS/2kbdUvfp3cfIpSe7yvKvBOAw4P
WCEmg7jloNNZlWjj7/r0uCyS6prOADDulyFp8QaTk98ZAENpQLqgjyXYgaZLSpEY
HKN8WqA5yX8b1HXNChavDwhyynwdpdLg09xMuHhgurytI0rVeGMNg1tZc3v+eJup
83/qByF5CFa+c1myCosp5A==
`protect END_PROTECTED
