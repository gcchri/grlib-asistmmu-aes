`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H16pHrTpQnXT7KrL+9AwTalh7suDmLVBmXzM/e9bR45WcnOFKbyVH4dlG8HKzrMQ
LNhJCu1I+SlXmWf1xJbJ73wdQRcQLgAGZ/Gv+qUxGC+NWnm7qyWw6JrOBKR/vla9
wOlKThZURpF60qG5LU+Yh25K67mx1MlRyCb1SD5t8OCCHSVotN92nVPWQAGbUohx
/ra5nHwOSTwpBNz2zEUZJQd7C/fUXlwqXCsoqJsOkYrqWqxPIyMgJ8JvY2BKhOSL
skOs3SxNRG6BjKddtZdliP+VsxW2ptip/zLoOwQ3O6kW3kRtgeTCWuEqaAetzYlG
aaawTz03fNzDrW0SAB0Scz8G8SDMO7HKm5U6bzvdaUPnVXvR33nkVvLFnROWppw8
G4Poo6dMIQEoFKsVZvGzhOnm+e+gu0dz+IhA4Yqq7q8F9jMmQ0QXJd2XKfuIf3rc
CNzXq4Eb4uIUIWg6cemVsdS/jhVkFJNKFvAGiWgh+TjihBp+LaxF1WBbRZE5ayhV
dF6okZlMWj4FHsAN6NjRgkRg8tvObgfzb66rkXNYeULg3eboMRIvAWgmJ0zggeRf
y3cL8vI4cdWXAyohMrlpGQ==
`protect END_PROTECTED
