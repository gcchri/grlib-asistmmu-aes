`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rhkm4lKy2L4CDBZSVfipXnYphfVzlc7cofAWqi9ErRsWdGj3wVbkFeclbv54rNfM
s+AJ5Xnc/qw/WNw905UShgBiVmg9jT6n5es9wm8ZNAQudraYsmaJPmtX7zEAQAol
oVT7AzVvymjk33ho3f0+mQqI7QK8KlHyJdWORLDVu+4Yvr/y1yJImRP1CSh1N1FD
CA9Yp+syAGYmn3lnAyxNjcQGC7oxMSCW4pOa+c/x+wXBsGhdzbc6MHHjYodkrvU2
ox3zXBkh5b+iD5aqKRi0akSNg+93ypzgHbCn0WvF6yZQEJTXKW/F5A2wo99SZ8as
Fi1OFN3CJ4WngEiM9NdV1bro8egf4bfeCmLmyw8soW/pn2PWuFLQz5gS3Ua0hpmu
p2Wt+rBp+/X8Ew14xyvF+z7vxjsskAQH4vNup8YPwgioI2eTgWm9C3DiZWjdNdhF
G+hkhiYEUiyzAR6Afs0vtcJ8ZO4aL1TncIad13Yu8k+ZSeJK5RJIR4o8X5ctoLIV
ImVEK2GhHnDrQ8JLYrRgXJ+iF1zHMPXKagzF1hRm3QWRoAhL9hKfr8yXNfAluNZm
UQ/qcfIG/rxZENplUb6WTJfawDKRrFr2uyTN/ouPzkxCoAso5xV8IRDWdoBqCJoI
8NpHudZGfLS3iftt8R9A/A==
`protect END_PROTECTED
