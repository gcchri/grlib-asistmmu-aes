`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ROliv3YyLVyRZDUaa6Qvl7mFA76C7ZUBx0uPndc1IvgC0QO0IdPXqv6uwPlmohtK
/ka7jZXabLktPoMBN5k6iaC77m92Cn+x4s2CJKDocAZ46wVRTQkXulpD3RFa7S5S
7osTGkv43s++1hO72Gdx7xG3mTFEJMH6osT9MznxmFxkfavSYXV3ovWvJqnaTzWe
wGgyNimxe1thXBgPScxMeRk5DDRqvadotueO72tRhzm0FF3t98ehWt9GvZxfw9n4
EtwSf5JOfn8ghjmnyluViXZDTcJoppMqDANmrKCx2XNxsXcGqbcSk3fE5aKe1fuT
Gwkib3UJkbvFCXtY5ZOzEY8cbzehEeeBSJGYO2Z16l7RLv4qPprY0E4jvm1ITcZW
8Ws4vyTBVqjKwuOWEp6nSBsGzZqzs4Ac4pk+/RU80c7iGJp7q1/dyNuZIncj4rOX
y/cKPdm6jjGvcz+NFFk1kihl4iReQd+x5efBYNsJjdotft+diuk5OTbXhTYAe8pq
mgIOHIM80kLpSW+4Sw4BBNlVfIpnTL7sn+1JjhriEJrT0GKoNm2UKGP7mpw48end
SkJzEB0xnDiM9aPqqnWB1c7gzo6+1u3njcW10O6ajrKJXpQO2XTN7rFQVAR89Jhw
N3xQE+ZGYvqNdcT+wAgS6VDDpCdxxcforcAQWYFTvlB8gNabFh7369DnEe0GKsgu
wpm7CdTeoE0o2+pebn9jhQK8eM0DfhokhLVfhT1GSSOTavQCfdGH8BVQ9BHLNdLO
0BPHG79IgVhNj35yK632Y0Ws98+IKscxUQBIPJdNoxihNgA06C9PIQm8Msu9pcS5
nxCeruoMuKYRD2wDS52tGlvddAs44Gx6Nx8rTgFGTB+e+EIJC5ChNLejUhu8ClSn
Cte9Io4hajjCJ3aCgMAZrQ==
`protect END_PROTECTED
