`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lquT68lZR/YjCV6Q8ja/Ig+IB3eyfBmPraaydjeMYTukYb1Q2eOcJZ1FF1Wazye9
r/abSykBfm5lGGbKq3eq2IW71FVe/Yi3z7BfVsqCGXtikmHtcBLl/apnyCGUHS3Q
1orR1Id+PdUxPBnAKisCIW9Gq54KNRZaH66aIJuMHk346873TxYATXGkKqxgCtA0
NxwPvBHx36NdPxOe5Sn7baA3tPaDvuV33/XvrLJBiFXhI3hR3YlrlF0HSBZmozwf
T+tkP4bmWbfku69QUp2zZ1tePK6syHXo2aHD/SFzrP6BmX6+X4KBQAkEq8Yyhlby
1C7FOV38pwtW5GsabA8xHchLtEcoehy6L4FinqU7fCqokwaKRa7ChpBKyx6CgM7z
IFIV0rgExXPwIszXNuSNQw==
`protect END_PROTECTED
