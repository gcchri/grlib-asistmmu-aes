`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eoQc1JPVDV1yLPlExlUUp0bIsUpEkqCAgBYe8luGiI76GxxMbT9Uxg8lQ9F6mPOk
d/r62LERUnoWxvUjGPX4cnrSU24v0BDmL9KbjPNNPMGiQDlFfpj5mK1mTSB0ZwZB
Kv+orxldjnnEbo4kTmKiU0NuHsjy4zXxjuyGt7erAPDNCPToWH44fDI+eu1aUVQi
IXp4ecVxPROHVSPeIs03+04cSbFzIEGct2QHvVGfLfFEynG7H1F0NMAYZ2KmclET
MZzkwtt5zJ/weT+ZKpDhW6SKOsDMcUstbShi0W24ytJuRu9VR7T6npzoGUKGcXCJ
FDnShidFcABKgo0D4cxTzgppaamU5MpuFQKT/PpsV031CU9Z90imwJ9+4rSbAlMV
I1Ql9niSzh7ErMeUZWBBKHbUeMGYZUb77vNxHBXW9GPVDDi7LyxjsCdNV4gv70/f
ZlSdxjOHt43kKBpCvB/EJ+8VC9gEZJ3hLevxrYdB00kWQTgsPJcAna8pXJiIUDO2
XZt6Tt6kItiF+dC0Vj4Wo6FrdhKPmSQ9RdAfI7TI9Lo6G/l6UgwkGvCVNrh9+V0U
kO4ptEoU4FuEZ1f/XTPh4um3b6ZbrS9OXWKr4dKYq+yO1Kqe/VlFshR/shBn8Tsf
+uaO9o5pt/Hm357R7ExsPdYmDxpnZh8xNUQgm0lpwuua1OU2v84JwO7GY4Q5tMBC
vVqDzral46A7IG2rlQNSpMQEtQDZ+MUvsktviYuW98ywpmRywTcRQA8sjTKxH8ry
ghKFBQK7LNIkeMCLuNz/YlPHpMbIR0iy3eQ/WpUKJr63blom64LY5YYWHi7/Dt2v
L24BgDbAaI/zvRUzdUSrR6MfjWlniTvXPtjILlPOdHOl1sDLnidtFMyXmkQd5oyV
srBlHIMCTpmfmlpqntNkDSoC9yXKhe7mUrQpu7PMqyowpWcV5bw5HKE96GgzcfjN
mkGHEij41O8eHFj9RPmBucirU1QKcvjEVkOTdMR/DBcY+NqR2gN3AqW5FCbKWRsK
aEDwB06BFbiE9WmihfW7gJndng0ksNO4P4WiO+qFxOVlrPQCzut18jFowkE56MNp
HHLxesKvgrCqL+DieF/bYIKU4gvjDXHS349Jn5OGfQDfINwJtr7FaTupj/+kGcqC
fpTZVgDd8hQX9wcSSKB/1B8uzYFKbvQ4ZHnUY/es+5eXFzyBk8OWkE/Ajd2Hped9
Pohosp6w/ALRDUHVTwXyk1EbsIpG9hCXUvKd0l7HgC3il6coOszFCtrM+bCHrm5c
TjAih2uDNHQcEvLW2k2lLZtY/rO+TBnmqfA//k3tD6YDhq8CFadctMFza2JkO2sp
71jes0kBPpUVFaKF/g8JQEmPhJA6YI2nckFo4eCONh5IYmAfwzkZxOzNb2VdWgl2
RYCSFeReWHBPS14xSMOqJup/9gWNms+YLfKO72Gtxjh8h5Bgt1seEjYeeeqH5Ais
WSDS0V1KYsmd1zalkIdqjR1n7Eaa9vkgfxDj1P/mNiMLlTGeNvqIw7xa9YJFo3d3
gr+AOEtVaJNhL/EctriteXLQEe5KiwQ1msXgry8YgQA/ganxLmL6zrEtJq3ZdZ2i
yfhoXWabb2Vi+NiDGqBQt/9p/qbIdlFS6f2UJbeEAJd0eImz7Mnb075T4FI4FLIG
OKDoShKBD17/FdMTJhCJQ0FjI9gEnciRWqXYRCLYP2UJi35JHii3DKOOS7q/fTCg
/5HWTt24ph+gHluFh/reGeV2yZqvmRfRNpINRDbA7Z0c+MiqWXC3P8yM7Uu8GNK8
fArRG6NQnNuDH4VT3KiVMamNZMHwpnA4NWMZdlLJpjP9ZiTm2iG8DoL3tA4By3Lg
P0hd/74BTe3Csowv1gsnTSrK5ZJ4jQBe8RR3HI9F09vBHmnNcxEd9VBI+1SwQhTi
CmtYpSzTqeIu+Q3/xN9eSbaL5/sKqJlxTjQ4XfSJc5VjX8gD2gk+GiVuXro1R77T
f9OUCYgWzeMYYAWeqNs2n+NUwRi7cmI94elkhiyMZ/BcrVKAI193dlsy7oc42g5E
aa9lF+O8QvAVuXwqPGE9RLuHRB6Lmq771dT+eN3R39z4tZ6IB143TKe0RZHEUG5w
M3zkV8dBCYUpqyw/YyLvn8olfQGfOgeMo/1i68P7hVvu1LsCxNVAdRhFbADDvvEZ
IJBKU2OR3pXZLcW5It4TM34Fe8NIqEA1lzIwVrDO6apmM/NLtwjTWrrAM/87/nRH
ba+Y9H0GO5lM2XmNvh9AsvZZkQIvzvAAKYxmegPqtj2RdVDJdt29y4F2btm51wb8
6wG1VjpGbltb0Q1GtEBr3V7TLe8M/o4TGqBCJpmqlSdVRySBZcgupG99fYGF2c0d
LnIlqB2ysIikFSQaczlzw7qaFvfAlmj5WwCl7K5R2Q6Z5+0Dqpjn1QerAWaovHIN
ywjeGCP0tFyCTM82TY6TnFy4wHd+ZNUVSHv24fmuqGAv5N0ixZ3brcuENGWEvMKB
BD2/52ko9BeESUztaw0i+9tH8inYgFkFyBXjPqNmzUESkOQmPmIoUtCFEp0raG4D
JJNzqZJ2eiChts4jF8rTg9JBsWntSk9ryKtWxPmQHbA5CUhw4B2Al2f0mBpgrWvh
5Vncy1Miz+AYK0psNfEbJkFvF9acbg7x4u1GZVAg6IuE/kryEgK/ulI11Mldv6bA
HIn0oOTCiLG9jlGq/CjUsIn3dejXuXtMutGmK04CaJyfpOmMYf9zlqdSGghNvCkt
VUA6hs45bNlTTnhgXD3Sy/y6StgydzQR6xqrO7iscbyOGpxvWz3fcJfTYEa0eFnH
TBXYxeLVFah/gUFW5Y63e3/NHwiJ1/g3FB24iLpHH+2XZW6VxqBXutg521JmCyms
RqpC72FZ4qaqu0J/zEOcIQ==
`protect END_PROTECTED
