`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/x/KBt11mnWyYJaMOC8ycQ0f27FBwBUiV+HUyeCtm6Pg3zQ94Mx4kbjMcnnkIx27
XoPjMaN1mSeNyLD8Az5arZYaCQVRDNTSYVjlCkEOHlj3rnHcuinrPxKsw6GuJzVv
WD7hVSQhOhNX0BRysdtXPmbOdH+ftwKTK0b7T3cPaJEUjF0uXI1kOYKseYL7heeb
m9POnrfL8MLsdGa9ROBbGFZdean4KkNg4PL8IZGqyCC2ra6CW48GwqpOV+3kYPVv
18Y9gHlMV1NBKCWlS4sLrol1kkGe4hkiDidxVHEE208YeMieEY2zYW9MAvtegcDk
ftfz/OP3tCl4jABHqohofsy5qCJ+sOkyZ4ALBymxF9/DZdhlrSp5lC+xkwEQ1Wzj
lSVD9xRN9sM7Icpk22NZ3usIW+ncq/d6Qy3w1+XmHRCIG96ZYQlfQGl2UdtPyW2R
VBufy/1sV6gfgmV29kK9NdJB1kWVbHWJnN7ipR+7qoKMaBnMahHUZfYgHBYh17gQ
4UiTv8kvGFhe/PlcPQH0kxXz+OdZK+1CAow+VaEHgJrKCrBHcnZaNo6gDXW/GkKb
HCG+d14kwBPude5HbgiuaQGpEOhSxMdCNOUFow2kvSDpjza2kweUbL5Bxy6yNc5L
hJIm5wrVibngEXCIIUsPFhV+38HIyJA8d/Uc60AN+8AdXDkpAqi10MAuHshhMdWR
4bs+Q6nWjXHvaAoFN0YAqHoOrO9hXZKE6k6c6CIuDF7DxCDyzBhsngEFZ/tT+cRE
sh39oGlh1ewrQvnb7QTzEtuwFyA/k0/ybUENCE+TRUQdMxClvJT2wUCTeqZhVVrX
1WpUL8+cs/WLKTTqFPXB17IGNuSrqbzVT+URtRahsi0YkJCQ1Gegsqccx9L2KM+R
PMlepqsHHEdGKGnTOerdtb5KbQixiPf7FdX/zZUw/sJ/Nw7UQVL6BbH/cMgYxG5V
V5hpUJEiiH4IV5RwafvfV2+avz5pSqw0/VhFQWh8bDEXi5RT1Vq7Zsje+25BlSib
+xw/KbzV4sHCcYES+ScXLF0PoJ4DcAWekctMzAZPH8QywxgCk5gxPW2Y4tYo3rZ7
PRccmk9cq4Wv8YI790ZUBCwS9eeq0LZe7VzOihI/e7BFClw913ro1YifPKZ+viTn
unPYvJOVyxucGEifZu8PeimfODrY3gARMlAFVHhhNi9vPYqEKdrD2dNgSEhLkOnM
s0VEvLrBguk5j2o1FnuInQj3nPh+PK9K7AKI8fOymfJhxkkzaSIam/FNjQDHAVpI
vT+XmDu43dLvZM17NDYTFb8LRxC65+pWQ2MXgCuTLBBEeqe2xQY6Wjmf6+S6GgBb
v14HJWLaT0HGod9EXav7j+MPMSCnaC31lFw+KbcUoK1fwdlxvsujpxhC/KcSKu31
3wNTR15+5ptnqNRwkyE8yvdh7s43vpo2GHiMCFN19gHcqQvqIId7djCswZszMt6G
4Cw/lzokTigkYKsygAa9Dy0zX0gsh6F9B29qwld4a2bOymgIKFE/3LjVzawR7cRs
oYQwb+an4FdeGNfwX4ihJQepCuwPRewoJjkO66nfHtDkzMFSPhfi8FmBtPwXdpwa
9DQhWFlnQWooR1o8uqhAli8buKt8CTIv7yMQed4VcC7Cq5DUqgiMJkha9673BF7H
+OZG5sToI0dwtW9M1oyXWZOkg0KTy6fDxkfUqmpUB2NnRkM5Zc7c/49GHjEDGV5B
KxO1Gu8XJT/f889CpKp6v0P84tYjWyhs4GbG//l2+1QQqVVkCHecJQWem8mIOoey
z2G86lptdYyBBDh8OuJb1d+/wjnwRdWlgzAKC3ceHFbZNEHcM/G2xYlv96YRasOC
eei9mR4YbJZXBTfRMKoO3Fe/DQd/W8sALyOrxEBXuQ4sLvaqok7udkQWTsZTUtuH
PqxhLaskNp8DGcNJyMy30jH7UOVMYJUy6gqO5XrYW7YeGAgLsR8cWCASLxAgHNZj
uNgOeOl9flJ5LL1oEf7wVPrx+NGbhZqvbipnqW+8cnab8hZ1KgGxSRlylDQk52Y2
GFP19iBCV+HD4ixCXP5HLM80J8If+N8h1F1i0yIJ16Jga1ejLkIISXMcEnWr1UBu
JkGUwDTWDl5I0bdKWhRc495BU9iB0eqwdW7hZ2e46TFqyFPejGT3a9KsVsDpWsgT
8d2CbGQ87kNnYLSndTyYFvgZcevNOVjGuUpHASoLYXeJVKp2RZWdNPbQSYrIdfSq
L0Blg9rEWGkqONk43XSJqU1RKBwqddSR/KhGvRcSahNIKKLigo6bb3NC0Y9ESfWc
QcCnTvD/eN/bIMg9U17iGPhVeAyI2ugSwvZi8dfgiMTiVj32ka3+HUVeLH57oftF
SycrmCueKbibamCqjF54ny41KwiwN8aOfJ5IjtIzVUwnxVFi/DXHmcuojJPLslnM
5/15rtuE1WjLxEsdj/cOwfrRkmYcTK1Ub5p7aA3T3bXfsrQws/MlL/Nh2AxGjpu8
7xGiGz6kUslRrXoe/WwFOVOb3RFFKKB6f/udnClRBsJ1ljwmhCL4qIAuS4JC3fIW
17MUeFsFBkJzMj8cUgfQHoPAApRenOlade4vGOnvrbDhlCQwljrOjRBtFoOz6qFk
rFrRZByPo0WuRAkaRXjZsrPcXXLZkCgmq7oEg3UqJoFbnueGFTn+l2+7tXQjQi0b
+w2cF9Somklg5jhdILjF5Iiop5uircV9+P4gstaqKl7RPaBEDl+n35M4mZG6GGea
oh0HHV6Z4BHeg6A/b3Yf3pu8FH+XTr4FsO86X3udbkt4KhNK1BaN2F+wafaAiPnU
WoFZM1m3INXra6u9H8Fqb/EuRj/hWHSpo10NjxrJk/Pjt7433RA+DQoz5eViJAwg
Y60mCs2iXIda3iF8c2q6vhk21rFYOSRtaDtW9xUEFUgBSS4Ykw+aVcnjl3tDWA3s
An2heYSxvHxJNSCc/dntcGSos/feTCRcvOtD3oJv4JNU1rJLej3geTtirv+aqGFI
hYrnoaJ4xkvJgBHi072Qtru+BbUS5k+YrhVOzj9cWYxx8uaFMFnCt554RKiRbyxw
rsUlOjUl5Org5jUrj0zF63FU8lqoOnYO13P7p1vF+W1v/na4J2oAYeajMPDd3RSW
`protect END_PROTECTED
