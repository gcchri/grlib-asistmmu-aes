`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iJ2TS12ggn1/QqJSL7EvvE+6H5peSeyFi5fQ5/8dfoDUMZPJyToa5UPz+Mzejr/v
xYVZ8vqQ6P96FvAiQ2lSdL8CitUnvgaqdeIA6Dk42o4pgG1a2DLhbMpjWesmCVna
x9C2nZfHNkaoPFM2SPsr8t5pHCFVrC1446m9/mdPxKyky7Q8EoPP8E4tLwCFuF7E
3ALLS1FISrvwkFMpvg8wzzHaxR09UR3+omPFy6z5pDT0T5OhuGrG/Eh0ibWUMmlU
kUis+SYS+pYBtCzilESx3RIGFtZx1dPKBk6g6P65bXIDX+OSujRVYwI4p5jh1fcP
57TsnKJKoZuytn31ooN9kH6x1O47vezxk7sfd8v6R/YnJR7vEQF/QHBMZCz3g7Ci
fJo94mLH9WkY65WLpd2id1J2VN+v5UuBQeuIA9S4/v7D1SOVfNtKObz7Xa2hdE+j
4c+4oQuyTOXrB8j5SohzAtsyy6HihJbH7VzA8cpvjKxFZAunoCrtAuJK0/uDdynt
VYer8hFQVtU8/ZXRiAYlPqZtc47T6y21V+wZyuA0CowIQxihlTSAmY1qJC/XqfJV
GoW9v0KSugkDkmlcvk9AE1n1nwbF4FaNgD6eIO/ONWmkQDeNRTtneMN3vCHdEPKz
BXqskOQNpkYTg4t3tnxZHieo1VGVVl7wvvdvpXhLFLRmkMJyUQllUNzgDqSpJCYi
+BKGxzWsBhsmqv7p1FdfJ6nLrBVXbAl5L/WLqELC5J0JvS+p2FdYLNih02ZpbBKK
9mQRdUwzhpay5/G8E9ArSlvMHxhKdl8HQyGCZn87Hg0AsKIODCc5Jr5lcMTvLPGp
MZtxeA1iBor5PnaCy3SjiJkZMRBO0zcvjorYTAlKUquthmqLGl+JMplN2eVGfBip
lwLzX27i3Np4EB6vwsldwp58+Pc33nE7fHlQqJwjA91qqpb4DKJMFNFbJRRAda8w
I1m+0GYVablvX4oZyYTJ4gEWpY8X1yIsVO2LaZkbLt/ZwbA2tvcA8bITEcX5lw0P
AZI0vWNm2Pq4bXAnI5NL+bzx9F1InQdjLhMtT8BxE4/5zK8B0aPkXACTiD94uBvJ
UVK2NMrWbICz7cikV9hATDh9m6jB/rvhwVPGaUVuC+OPTgn9bjJgcmD5awRqi8lr
c9eXUROj8f5H/hhjXaDEFUFoA2zE/2G6pZlmS8oOKPoCqv2SDuohKZ9LCgQyrY6D
iLeiD6775FcSpupGJb48CpF3gcrrhpbzuATXVu14Mphw/EXveu7NH02gRqVD0f7m
DkyO69ofT99e1aDZnyIYQsHgNLLln3kJAagi7dDhKsY/NagCQIWApy4I9H8ECqu/
wnjKgbLhpCKa/JLO94kj17U05GODca4nVWEa7SU9bNvjYigj0gnTJaX5d1bWQfsA
tkgYUto+dLlsBEELHjC2C32kW/5mqKPwMFRpnXixFODS7YgunHdYjXbkoyHbPmTT
CiSCTPfbTegKPRSTTQ2b3kx9c7V+Rrk5uP5VL+TYtYZpzYtX32BcmAmf8vv1lXfu
oA5oAIInwc14fhSYwBHD515i0yvUI/5KiSvx3lpEu6V6FlXGHfJMmbobtiSGraR5
jkhrm0sMOhy/mOA+J+79jBjEMlGOen0ypjeFO3+tSm19cketGKEP6zJhoC9IjcRa
idq4tfmQtKJY5XmZSDl7GxiLJd+JC61mKckCC7x6tGNWmcBDKoLCGdHCiOTO+6Xk
3Ye2O/4DbNoAOwCmStayBIqZl/Jh7WMZv1KUEQnNxinv33QFuNdFOv3RcFAYebSC
1axlRo2K6E6hXQvQ3Hr4Ke0GFIwjzI42+EwmNQuLhtgH+d+xwYJX4GaUs3RC3XaE
qOURhaOUkocR0fAUcTc6BdfO17xyxZz3aExopQ22OVRYdrCNbXsCPO9VLvQWv5T+
ewAtIm1J3vZqOrwG8n/UyZT2nhPTXErlCynfBsGyEAePRlBURvGqsHUB5WvuheLy
oLEuxrnenJm3EmgQrH0cZxaE+qCz8nggvkShUFF/FdaJ70dIEf/tACsQPQ6H/k4N
KmLwMtPTABa6V3buG5qqO7WiqTM0BlzsBema2hJAc8NAMU3MrL5zeRgKJHWqXwgA
FRhxXKdjye/WyGxzTnNmcLa4fdBkZC7wufQEZ3Tlo4LcK77Ne3CkJKwKS9CW7YVv
s/9v6J/ulRVXmZkJkt8Y9d5jKvEVi0/qLJzFOGD/BJx5gPZC+u37sKEoUyECDhTp
ShQgpOv8vK2EFzLkDQXldCaFxpE0lfV7VqC30QjyGcHdePJxCNCH752Utv2zrXEx
EITeRhlf3ERt3kYM5TNrKt408xBFkplyQgrDi8c6ebo8qm0fvfoNxXmu3Z2Y6T9g
i218WdhgMBIuDiRbU3i+jvHNQICUWzExNi759/P+XySbHCV2sOtVXigjxe6rqD5x
6k92z8vGP1JDessO20posRV2HVCP8hpsBFeG5PYELrpIjKBymkDDxANoxJaDiRAu
C/NzAX/XROWjcy1HfFJ03EgoNydQMj3lzAw+5ouipILC13FqnbGoBMpNGRGmTnFc
RJdC2cYmD+Uy57u1XU+dJ+Q7bpLkIRONUFFOgKjXZhfri1q223slgNlJR1SULcUq
HOTJP0M4QHzNx1XP52j9AivAnjDW42SPOGrxknJhhTD9Z19ZvJ3QKMP92axPQhce
V2gr3OMlBCH7wXhvoAPlwZd1QftSYWHQqaVlsw0SAQnkFbN1wG+AZVpem8FUiqRm
UG3eO7gOYwLaFP2l1hyAIw==
`protect END_PROTECTED
