`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HytAGKNbuED34T/lOSM63CQwbeM18McUNbXRKoreH9eK0raDQAK6N1whiD7d2Sy9
2oQNChAt1OSFdiKuGb/tAAf+kR2fk57laFeuHEL1v+wJz16NgGvY+NHnCVivVl3L
IU8LMXYPwR4HmmcjS/i8gEK2qlqkzX0jazD5/B2LLAm5bGloqSXeVYvX27NI6Agv
0mmr4D0gQJFSD4xOXIbC/0otaiDJUwkX6ZeFuL3L9XbfYsUMj+4OMmPaU3n+QJs7
KMcjg6qiAXw8I6YFmpwAy29+aOipRhdIUPK1WxBhpZlkAcvw+POsnd2EpYvFyc2b
wLMjqL/WvjGXH+KyW/j3jZckxW+/i2DBeSn6HZu7dJooLMoVnkucWWehWl4dwqbO
NhXr97itJJAgmPbPqxFSqtR4BGgYJ+wEydl5WL6+KlHun8qFRpkBanZwWw3L0Sq7
/zvGnJn47zTFzeq6Qpig9603MlCQ+xRSPvRZtIC24DM=
`protect END_PROTECTED
