`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bOmctSSZLFEA26gCjUVFLgn6oye3VPnmbYbCFROgwBk9dzS5HQTjgujBnXti0iFJ
ewGbP+vw2OInxgFlNJgjH84lImqVoGux/3Gv4FwyEXAZI9y0GRMH7BJYEc+yNZpl
Y8rONpujXnfIs8Y4SthckYaM2mgb/eJYS19UGro7ZsdeOQZFpKnQvn4StcPpEdwo
WWcUAmDTnUjYca6dI56I+FQWMMkqOdTQhyL/T2/lbyhr9IHePsmQynzsRXm/rOBA
4k0xL0LmBW/U4R3v4M94dpoVWegg0p6Z5tzTeLMGh7wdddDFw9+GfIwdMElQw5BC
4BneyfDM0F0HrlIyeRGcxPtSutlOdJbxm9w4jS/fxy9E5pu/twZ0Imf/c2/7sA1i
Ld8ZlUgnYg6TROYlp/oMGCg6pquQfWTLKWmaJcDsTW4=
`protect END_PROTECTED
