`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TkaJYLrCSS/I3eAw03Qrv1j+UBz1pzF045t5oE/u0PzivdbLnRhaBal2PnzHktUJ
QOY2f6BVtWdPrxvoJgyYF2AkHmlNHBkppvp/lLli3w5ZwLp+efS0cMfhTgYr6LAx
hTtpfgC9KhaGHWUxlSEtaCMTeHJHCBBSvYYvNFkJNeVkc2iX9NpjvRCoAnHzbDBe
K7GPjyVSkk+HUlZZqZlnVpQpDvlJMb379kwk0dc3jvl2sXkErcpiKzNHN8PMxdmZ
NO9CGT8Q7K7ntjZ56QISV3Ym+ptmguhjx7dmFsV3c4t7mQQjCHzK5WSewjusiYPj
1vBxWukyMw6X4YDxzPCkGUDxf92CBPOy9ORIt6ubNI4FeQTJyTnuiqyLSnEIcEqn
EWCG0HytSDbSduCvlvi3LLfYLMj0YVKJUM0OIeap4iB6FA+N251IMIN45kxIygxU
`protect END_PROTECTED
