`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IGPE4Jee4DXbI9NQRRoGnPdnexIfxkkprSKWcmJWRYPCZNGgkkNCGfjYEepYPwVb
i7fS7AFW2dVtZwONXPC4ZCxK7cTueGbXoUvwnMZZ9t29l+gTL/k7bFjerrE34tOl
Zq+m4r2ZuonmPejQ1605W90NLjkML0XHFMOhAUkqSPeNQxBs0GSnMeWsTmFFvjBm
yJem3cqviH6YxKh9MRoR6uFX29TKb8FgkaqaX/lXQqdF8chttCBfDpkruvCtGlzS
Y+B8D+1j6MDkSrBWb41FSMWIfxSl3XUuxGaL7djft8LR8WeNjGaQci7u/xdD2+Cz
YW/jAk5uO48eUtxrnpL19+WNZDgQ9zOVedNwXyCX18YejFfRAIUgP2NmiSj5dL4v
51xNKsms6mOxGxtGNnUTGswtG6k9nfG10OqvKcNey0SnKH4FrewPoz2kv6SeWm9a
jsHS1WvehweopVbxN/OM7RaoZQFQuMWRz9+ApJmvCQez3AJw3vxAU+NGkiVX8uGK
`protect END_PROTECTED
