`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0y+U/Qt4PX5fd4YVBiaYpdy53XxShpPSuw76fM9USeoSJ1NoUCJRm9fN6IQUCzIU
uIHKz8hxtaP/fRcGBl5dtkDJjL8qPFAH/vGNmT1w5CAzw/ALlmEbgzsAAKVrgow4
sudTrJBUzzyPo8/qZmv7ZvzDqM1YyDsQG4Rfh8mIx+P6rkM7KJLz5IL3Tps2NdDp
t9w1PGhsHoIPc26XyvUKbtvSs0MlRP6Dk8O+26o1eWNwZXJT8VfOPZmJfTaq4IvH
ELm47NxsnNxpaTUNkte/sSQXQ36QHm0be2Kvuh8c8swivqjNqBO4zTjzMLuIT9+y
IuSULOw/dT/lVHKj+GMfaJ2rNL+1vS9Lop4FlwiVnWn9eeGYga3BlBm98z/bD88f
dbkVi4JYnWMulThfBUTVdnh1PaXeci3CU1SFMYBgAuwyXv/YjB9fveUpPLIGDT6q
ssN+w0OhzROavJB45y8W24AS2nKC/Uth5gr2kPqOdqygvA7MVlze1be+sUo0bDe+
MPtLH6PzpI2f0nPZfzwEW2WDJ+ilfj3BIu6mIqQbXr0Z8IdCtqqnOgztXqEZwhE6
W0Wt5yPswCVbYn2h9T01jMXuQ1BW1kZAuV2yv+tDXDQSqj2UHigy7yfV5tVY8RqH
zKp8PKW5Thj9yEJrGtNHz5kYCc1OF/FyQ5IVG374f4DJuIwCAGWFECz6RM/7mFnz
C89jC1h8ksDAVlCTZ0oacTOqeXkKz8YxdHE0NynkFJgyaT7evOKlByOoY1YuMbBd
aISuf6txNIhEn6G29uATOVBaKqudvMb5EIlu/ahyeG7NM7VwTp9HwkUfP/94yhBN
KWyb2rDTBSLddOIKIp0/g9t1oPgRHDyAs9OgY8mzcYcLklS4bXHAA/hJ4QrSLCqx
UMGSlhzroZDZtLf4smCySMCLZwewNzTBU/C9mQ31a1eaKmM0PlJBmXT+LOkMklve
+zIkxnF30OHo3+MhNqpymwcgRUxmwq3hHBenvaRPgvPvK9ijnprINBovXKF4yBfg
sJ9ObLMhN8hMWW3vGLbLvbqTfRSOsvCNX0TWss0Tkf7ueye+AyX7rbvIGS7htoh3
TeCy8cbWdsZHxdT2qaaAdk1l9Bd5BaCg8jbXZx/ZRzyE+PVDZr9EjnkrhK1rHGZR
xRcI4mmcyPNhxDs8CxMyB4s7qjKH6Q3VcKwtApoORSbo8CFxUHnDKAmmCF40mgdr
OEGcxajWLOX8OvIi5e55yDvZKxjlSL7hTxbMSjrH4Bvt7VKNAZHiAhz9T8h0H+CR
XiR+ZunGmeX6UogGB90dThcwOXRAKmRlx2vi74fbBdp7AIzGQEOPhmKRlN5SCaWC
aSrLDJ89zmKXTRCgvwErcy8ziZ4MhOUKQSzrG7ABG3npOSjxZFeuIelrdlVuObHz
c8LXn4vPRh1az3fSkX/2xI/FZ9eSqfTnpKUUmvvfYHv6tGPoc69HL2XGc/sSLRK8
cMgheYx+MoXOqY2k5stTaZZe7s5O9jvgrn0gYdyh7lfDR6AdruWRFmbur4c3vdiu
VluAv9BMcjApM4WVMKRIzVCJBgOMFDSYDIpdxEkPAcE4ropeZvmiv+9T+L0prMWC
6Dq5PTNzQLI/l65dbqBW7G8bnj9AE/EKlZHchTLOiVx4at3154L2gpaWMxgPVSi6
r5Gp/cGVZsNPpIn8PxN4C6haDja7050kMdeQln4XcrI+fRq3eFl+okT5jeswFwi5
J/ixNuN/+bSTliHQ2GmDNMN1zFwKx8sv5psV/iYoarmpVlEY/4oiy1OKGnwqoPSN
w304zRzH5l1dC0BKQm88tC2aPMBvfhJaRERD5J+Qpu8ZBNHMdid+XoeHIKEKXrtl
wfhH+KZj3PAVsbUNW5PTI12g2g4yn3hyauhNc8c0jQUfQ6lcNIxtO8MHt62jlJuC
djTLSWPHv7D8v6V05dlxDd1sNTcbTLzt+Ny9tQjQJsy8ZebgyhO17WRCN+LnUe3w
i5q4+TIs2KThHAP4Q9PXB8+dVNHT1oI+fWuo1jWzaBlXtDfP/O+lRfSS3RE+ApSZ
aKxafCM4KTQmaaXnHUvU3A==
`protect END_PROTECTED
