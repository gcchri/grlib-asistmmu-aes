`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W7DQpMK1zbQv4B2lTMOSmsj4HPTituXjlq3YOfgzG+lrq3/cziHGOXaEsJyv7/GW
PyZkqx3NKw7LF7KbNwnEkjIVtb9+DPBrDEIj/Xmw8ZIbyDAbbKQq2JwyYsm0wU10
+6j5QwNKVAKFKO4aWxUvzBL7cQuO7lu5CBx8j2ZeY6ZbHrm1ZwgU54agMIAT2Mde
6OXf8YSwhMs/97LJmz3i7lmDgoDJrsZJftQlCaHP1pklBk7/tyxNQL2B77778HCQ
tcD0Iiu11GKrff3sOHmZDRc2HjDD6JZVp6aObgLjVWCLGCPwkFtRA27Z+O7X4Mr9
5j7Ql5ecLwRXzkY6MqkUbfufevFjhCQb6dI+mWozP7DjFW6z6V+iUGpSlG+nvwTN
ewGnXRE3Ht5cEPFJrRPTwvCTwjwBdF9CpKEHzAn6uFR2Z6ml0rb01viWJ/ZWwCfc
qki03iXkt3tyFRWBhb3+xnPC0WjxrPOyApVyfxAjMixpg+NYRWnjS1Sjtipw3HCO
Q4Id3K8C3LSLYt0lRyQryNL5DUFRzwkYcX0iPTYW3nlLLoXtr1wI2X5QAa/HCOOb
Kp8Y5jK80JlNezS2KPD9VP4rponJVT592lN+aRc2OIAuUfkurA2Fw+yD65ajVEx3
AJYgDM3KGGhtyT0OY0r9KXa4XXkMotffbnKz/OqW7NfgcOOlaz4HwgmKjtfqURCP
/WIo7BtDnQwwZSqvdimvNwgoscsrmHAkKa3HzqCmaeRSvZy6pJ5yMxwAIwBpbWKV
01wMMhRGK/JbZ2E0LDmoeHpBYvAskrLcpZo25m8Pv34JYrah+FIQW6BUcby9khDq
fe/wHmjzGYGZURQ2u/MSz68TBvIb0M4+JO50CnnI3G8pBF+G9aLNUCUmMnJXfcc1
mLpGSpkVsg2fh7F9Zqgb7fM0NsWgX1t7ivIy3pPG9TEMWzewhDLoAoE5jw3closT
C+SE6q4z+4b4ksuOGw0uU0m9/7Itg4xrxFEY0ABCVJpKE2Kz22q6Lxuic1zXdyNt
5gUWBcDnF4wCeK68x10FJWruIC3FLrKQ29V8cKbLHAvmPaYHde4zCY658pSC3Y+r
SnQPQqwdeETcjiUrD6bGonqTk1nF5m0lHcola09x+W8DIgeSDzilmlkE6iLyKv/w
`protect END_PROTECTED
