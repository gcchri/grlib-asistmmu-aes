`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HF2WUXAv6GPg1wExLdJ8foT6iWslymK4aJm25jK54kFffPSXCJYkVfp/2GHZtPy+
EQvngqlgEZXeJdVnMFxkRJz3eHL/GF/0/wB8p9hch0t0I0PwFwxdMsifW4Yg3fWJ
MvYLLQt7uP+8cUXKGJc+rVkT9GGVewcU3Y0LcZseYd7q3OA8qbGc1ZBc1T2dGSsz
2GOA8eJWoANHsKm0Jv71q3ORjMmR3DKs9leGpEgzLnq4B4gA15zGuXndkcRC4oak
AsuG/KYyGeVdUqCEpFvfQFQOnMmAn7oMOsY051cdtx+tohSRi4MrhKXqlWTBNkT6
sl+6nAS1df3DOLKKDkahCQ==
`protect END_PROTECTED
