`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fEWSQW8tXitm0eGOgaxyzxuKnqjbgzwfvhWmJiKCKOXqrcVJtQS9ZBs0FZKdtDis
KTSAYTyIFkw3M4VPaziEZdTyPyAwtGHX+mNMCLm+bS8GAvKbVd98KHZkhWUaovUB
NuzC21BHre5LtG+/QxYyQLEIHNgzelHwr+AzgMRgsrgnAH34C6cK6l3yDnzgScjy
k/auuFpfBWjCOXgNMS6zqbowC7Btne74Zafh1aUP9Cnlig6jeOW2B9SWoHOCT+3m
zyECQMndWumJRD9UUmDNnTJpjUrojzXFyVGbnpTbsaXdHHSj0+tMsWsZuQqjozWb
LoERo9s1ct6NeD7qeutf+JWIdgcYTRKRzIl1i0Fp+zSUgWUVV05u/yEXLW5HCXaT
fMiIUmJv3tFPGQkDW6wG23OUl0gZOoci1NVBwOgGIOo/NQoPlm2lgSgyVsO9Kgqb
/fEL1bSPCbB9G1eRJqpfbQIgQBQ+TfqVgmt5VXtDj4De6OlwfxOzfqIjgE1mZmo/
p/hVxnN2yGJVRreGAQw+TmhKBjQEqczgNkXbU3aGXl20oX82rRXZx1q7b3ufUHry
Q2erVadmJlmfGFBH2WUV3Owe/gTy5ItXKgZvROg9GlcR7KScQIC9Ah+J+OH+r15e
+lYonTcSdug1XZG4p4ayewE3RLtqI6qVzKbWOfDBEQ4REqhxM2p9JeJDYG0l8u11
ysH6HTaTEs37vCYujgKIZSA5Ce6fZGP4h5T5RXQXQw38E99TDXum2fSpsIVK8DVO
I7qwtOVIFENiWxuqY57lc3Q4gF1vemp9k1WLVkA61/IOcGVMd5kWHm1LqYD2QU0F
+fAATdtfKJM0CTvOLqIVKg5dgtyuehAUxKhqY23tyrWCF3RptFJhgpt/XWXNbwag
V/t7qkRu/u4Qg0myaMa19A==
`protect END_PROTECTED
