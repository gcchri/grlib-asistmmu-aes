`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WKj2k6MrjqdpWnnWdI7rAVcQIVNOxcRGsPjQNc2GHONhwsPy0IYkloQ8wjdqhMRP
8Ta5nY8IjbBP2UpLeZBS/ht3eVjV1hyUMd5GeZM5rE+ntNXEw1o2fZsO1uTN5sm6
OkRvecwdz1XXcHu07BBM16Z5NRy7VBTC7Y12plKSKY1uS8Jn0xqEJy2KeqWFr9qI
FJVqFdsIIs/yLCDmoQBlGHbLPeW6mD6nSWgn9POMhnP498rFqZ4jmdYEEwTGnNPA
yDiKGOd9/AU/2e9mwPaTbdepBv3KrwN4NEibhKx+Va1bEC+ZbM0zlrL2N1JNW0ql
huJEJ8v+mAax3+JD4ynnccb1+UCPNPQ1iMVn62KrWNoMAq94yO81MNgFVV6XEu+8
DX6d/OJcvJyq4FTPJ01fwwhXlBOgMzis3inip6NNYgKPN3qUNXxafmTgihwFz4LU
TXIpqLA7qdYulYuwQXeMV32OUAwJPS1RVSFYwmSfCTIF6o+3xdsDrfJ0CJS+qrCZ
sJfWgc8PdktLek+AFvYilFcQBZPuWmcr63appv/QZ1ekNalQ2RBVQj0nKyyl1BWT
TqwWZ0LmvMyMjHJ6LIiCwpRmzUZ2HaU2cpZNkI/GtPqeVEHqRM0dfxwiH8V5oztA
PctSozid9BkaloL/xW2IeJi4J1GjLwFAFHne0or18a4=
`protect END_PROTECTED
