`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BWfMPul/0d6Wm8eLvOtgadqblbJmtObRiaPojRg/YYZwn5J4pNrenqHvYxeT0m6i
L/FbBIUJ9fl2E297YXk/hOsab0mTIXwpL4/613hAMyg3WwjJG4TcSopiRlCHWsQx
bn+5qQEcT/7rHDGR2TymxQIoxwyQXhLY5Gq/wjIKbZ4SDyOxC5e9kLsUeCbww0+D
YlXXZr1IHqdXeEJtZ9fGCQGfFiFNuqEVY3WqtMQsTRY1WFfQ2EERM9dondtPiMlX
mkg4ZmTdXNiRk+f6rjU45FVwFiVJtT0FtziphPMdOPjX2+fKgJt0Rmz4tIIpv20V
C+hhY5zhihc2k6jQIcwjhPlaHsztebogY+8OHHhNWc/EHh2tXPM00fkQ+byt/Z2/
ewMEcJO++SPYeRqNuLLjTfp1rrzn/Kk3e6lkf7TB/mbjJyifWJ47iCWl8rf3q1ih
8ki/QgfkMiIRAi6V9zpTeH+HW51NYfDHNYPd0frIcyNDFOrSwdCLd//VthM6H1y3
yIbd7zMGmm7SY44csPtQgXh4587Ed+DiINDiKc5bcSNPZMSth07eMawC0Xut4OPH
4IZihTsBzOw8hRR9gxibChnqyhuS0IaQf8cS0qwvUOwcjnohajMtbroTZDF/cvSM
pbj9blYgSJN3C0Dwkd7yLUwa+wQEEjX8dCFnpvZ7NzneIlAoag+wEuNwTTyF3WDV
u7+0FI/KV806ve3w2OiapoV8ZfribqqaYV1aIM8+wJRlTPnoCIcRKZJSA4zIAQKh
TeebCcBxVHTzfLW0zsYLnNorEJZCSMylpgy0icxOS1r9Ugy6ttQY32fhSIlzzHLS
dCeoDPJYXFgvxPDRbm/8q1oaeB8B7M41LZbXzhyNSpt4CDqjfQ73EwwzKq0kRGWe
U6tfaR8NaMo19nYrYmf/kAud/Vgr08zGg0wN5YhZ9LAhAo1m9zk00GWndIhkjdC+
28Wasvuv4PDlyzX21MyaUDGwt305W3ltctiUEC5nN6TGSnIuGEba42iZDFIxxAcV
VzyP1348v1hUgTSN/DClybUYTbwzBTVSXKnyxjdBHwPwx3SGgYatieZ9kTJcJz5g
h6lVM02bMIUGEHWFMGlgkVAD0Tp95ixk4XBtXPgR8kRSjGlwO/QKQsylCDsn2kmM
zoZ/dVLXOezThGd/1HUkXebyKjozIMy5qahheU8RCcTvc2Atu1ovpmStsndY8q1n
ts7W1elO9n75PRdz1pX0DVckPAXK22nRR3jGm1IsLreeCpwmAdeGOJ0MEvpZjAp9
ffLRWmR9lzVVZf4mS/JG8Ox39Qp5Bupsnv7F5P+FgBeGoYg5fR8oxLiQpXq82oe3
DFYmyooswviciYNcBuNYlIM/+BYoi1NtHAmEY7iB+JDQNHw0DFlTqTUUy80/dfZD
L6yU53YYk1/SEbj7ybBHe9HvfuodzAdQ9v8PcPa1LQR4l/U0z2uV/O+6q5V9YOJX
AlsfwtNkaYkFAn8mlllmSvrJ3yCL5PyJnNSo7QkeXi+sZPlxy7Uhp4Sd23ygr7sk
JUAZzmrLCagk+tgVhjA3FKTPEQtokbY4F/MPr5Wx9+A41fju1noG4yfSAG5ceYrm
5q/gFRnsBXd6PXXiJNHP17kbUYNB017IuoMTXacilezgH/5t7jFwfKdVp/Uawfju
I1//I5qac5sLqDzXVe6ZowWtqBLkJvS/VUSbEldaZZooToGrbRdYoco42uAwCMKt
jNOicpfmhQPPAQkTp+NckrPfqoHv8x2ejBixO44rZICNb3Sz8y+e8cBQRaYFe5Eh
tfkeJt0G/eEfvkbuAI7zkIIXG1SYe45jjdE+D3sxXf4mDeJ9HhiW4NUlE3W6yYHs
WKum8LQokPpRhvQnH1j0Az/l0+62slw1XiJWJFYU+OFi8WCgEVAwyg+4uSKV8JhL
emSM9IoQ2UClA7m6q67JeesGr0hoQTROrGdRVdjWZ35FL7OJjCfOM2iZUvh5wRlo
BlapN/N/UgmMfLXTE5KhJTDrfO2Ye7F5VzbfEfkC4BDT+3+nb4TDG7/VdZDeEzvZ
0PIdr1me/4975fs5xPETioisRlDYNzry2X5y2XiL6HxCbYMjqxZFsyjNgysLMCF8
9HUyRWUkT8cWypvqbFuq5wNsQuVPYuUCrJ8Wf1cZjUpA9DEfWoFVBl0U89VuaA2U
zzgzTLg2OU/oH+R4RiZxER5sSxjwdgLJ/dL2nryQN+Dk+odv/AbQxr9v5tgAqOPe
8Va7W4f5dEFqvqqp4rZHp2UhdwzGCBYy5dxEjHlT7EA7YYYFHdgbVnLzMTSWpf1g
eTM+ouWPytbLNJu26X7HPnQwHCTTkrOstj7pMVVWp39SbP75UPK4bMSZSPGx2IBE
T6vTPuFOcrNMbw7kxVBChQx3iGhMEiAk4iKn5ojRFXA508mH1MpUzeIsp2Urfeir
hYN/ffcL4waJCeQVhRz4eiZbA2UGpsTr9oVAIwHUrWoJdCeXCUSYhTsTPzzR6Ko4
O1uRDDFTGf89Zl6cMmckVvgfEjs9kF9gQOfsGyeREwCxSub+63WY38Huyf/xnRf5
TpZNR4mc25sBvOxI1onr9XIBZHwsVZcXSbrubgX+xpqk29ghHc0O3tJrQVCOMP4m
HB1wrZrmU1AHzOBp0iW6Bo3quNmCyykPogetTjOlkqm7Ff5/ZwNfwiZ1qpkETLCg
r4R8wdUnfrF+v3A6P05GvqSK5CtFgcbe0St603WMTnhkHU3xq58Ftz0tWSf/fdxi
jN66n7fy1rH2Y97kEJM6OA2meDLVVEH1uY3nR7tUIFPz+G3SMEC7iJt642jollAz
rFlThApBhjhzbTLg/g5rOEvjSO/M90nsps2oGRDSArpNV8xa3NM0h5ObeCQWITuJ
yLC3NceeSQaLTLzeWJllFhS9FYXgK30R6UF5v0DjbzNgoJqxTgYNUPO2uy23fY/0
QW4JX5Tct1cSPOQlrTP7Ftv0BmLbLSq5QHg6wr21IZ6j9wLvJniL8ibfhOzImM/J
w/Zoj0qxf9ai/9b6aU+4dptPVNQpBeCWQswnzQEo4I8=
`protect END_PROTECTED
