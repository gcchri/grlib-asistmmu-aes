`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aEUPRVcvCObLKZqgH3jRiHuSX3A64m/eYyPppH8OPhJz3lO14EAWpu9YXhlbJBw0
Az41YRq8PH2Wx3UZe+9rzO0ifYlb8F19MnaaeHQT2USf2LO/ZgdvtUuKzzpNVOE6
oCuLgDFYO2RC/hzCIJG9pD2qWUVtTlsZZl091Uvnz1zyq/nnp6yaAGCjP1HVkrZU
9xF1Y48fw/lH3K52gFEfHySBpGFXxFPKcNhUS0a+LMvLupvsUgr2Pi2ArbEY95F1
cySHOiPmpMa7qJQLcJYj1jUiJyDGHE0c8LVeTuiQYvxHc3VAbi5QXDotver/Mo+J
t3v6Ij0iNZ9Cby0nn2RYlQ==
`protect END_PROTECTED
