`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r2FdCX7Np6VAHZY3IvqRxxpiDZLDKsC/8jrgmjAC0ArrAQpGWIC48IqOAXTIc93W
UVggEl/NOR7+xINuqNrICX0czCXoOX87gjFwAZG0qeL1N/W/w+Y5cW1ZcwYrjCUy
VXzs/JolX4eN2q30kC9tX53lNBbHkDnYS5ytXNfqWMblIcbDgmRC50DzswRpnRgR
La6ZAqd4/hmyLvF/NcA49ZeWbOVcZtfdmFbb8yGfec0SGFyOpVTRVQw+B/R2SK1e
`protect END_PROTECTED
