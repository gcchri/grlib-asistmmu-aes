`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yupy824u4wmTWuTHddIO4szALjnTcGWQq69yqt7exNaNpxW48UvYZs0fOUAnIAAD
LDh/u9EsqODgfrnFvhGP3XRrMQZ201BzyUbQ83/rArz6MYeEuZOgPPQuYENXghdP
J6PCjzW9bkJYLB6hQz9m9ENBiKhB5oAgDRtyvKfF+/b/CEKYfOiHY1DsYr/bz2BW
SC+Y4mJxYxj9aGyn12WmYzRXrNeTEyKnTBgpKC/+Zb8TIW1KakKKeicPZ2zTKOGe
tGFDANZJDHqC+/cjxBSvVW0QIDpyIfN+HyzZgiGwqIxlgReuTvD7QJJKvALz/rls
Bf4fFduFYw1VwBmHtyoDKGaMx8AAvGxCpuF/bjOKmNVx32l3aFy/c884vVBMAjUx
0IXGRltzBnoyITS8KF51XToltPJtmQge+r31ZPeuCyPJFZACjYdkyYMxqg0Zh3Wm
TmQEfCY4fZkaoYRQkOiLFERc08nE2r/mWY3p1fxOZp4HBVTUYsEqfhHwRkF9jSSm
uDJbkdk1PbVe+MdcnqcRiTWX/uUc4A1Rhg4Bu9Onh6ZdoGfdHerrM06QdZmPQvIy
zqiu1HRpoyQY/FKA3MBIzlqxWRMbMXv4QS5+x/VD2lQ0zO3ctSWPAdzbbQ1Ysb4V
OayUbZ10B+g0slTCCv5Z0HEk5zlgAc+RhFm89oDkceUMJRv+XK73VrxPXLVGpZkw
RwRHym1PHOhQGANiYpylsuSJU0tYMLlSxqQcuf9I7B8=
`protect END_PROTECTED
