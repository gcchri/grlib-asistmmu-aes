`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M9naoCcUSGiSwSe4+aeYN6qY3LCZcLCw/YpUb7ozCfvTXQIq0MwqtaEhiPQxbNOi
gAdhrwOCUpJTCfvOMDnYbaC+wOkmgQZ2P3B8JE1NvLH5mIXPOZYyc2sEnbIPiCS2
VfOaVSG1P2DVXJl5shTb1EnntRrA+L+eF6RAl4tAmlPhWySuFQ13BkWZ/k1QH9OX
sbQy/wTkT0X7eBWhZ1pmI/kNg26dH7e5KiBaD7en1n/aglL75hCyejJJYl8VzkFf
2NIlQJ1+/OQ5+vVeYaAYIAmfjtd0dSfaKw6b8Ul1xUMMo1JpoS2SpHI7FtS7IjWP
EkFktp+6OJFDSw+uXcPIQPh5GtVbyeJRp/FA3QIMw66gX1U2AWDh1pdipWIwHCpC
+pdJLkQp+iNELB79j2OP9w44P1C31gGSCEBLkIqU/amfwCSkJ/bOJSECMzlL1Gff
iXksMTjZb1M6x364VP8zaHpXjdV4TZDW1yB0LWDG+UPjUtrtp3okGk0s9BVrvSQb
MUmThaokUxd0qlXRpgFa21X+ow3uh64gw7gwB2nYBVSS1HewnYW27A17FR88VnnO
8yLpQBfsyfOF4RfhbHdfm2JOEWMu7j4Kl9TgMZ5j19J2mJ79qhL+Nj/6n7Akb27m
OnOd+L7CkTKdXkj+Bph6EqEVGISey1MMWOG2uP0bkXhjwuPGtTU2ZwYi60rj47j7
/ysXZlo8zFdxntYcYn0V2Oa67IpGIsDVvSg90OO9XWrtxfECOwtaRMfqQAPxFlGI
vk7DxNjov+AB1vG3XAlwSFWj7YFUNpXWQO7l5fhG6Qfg/1ikVo0NVOMPXOBsvWAX
N8CbSNR+jPQ4HJj0wUO+ZGIcWcv0Y8tU0hphACy7Azi6WhiGyTBxgXs60x4MIFI8
a3SeParegsKAIKWx2cGcrQECCltZNoa0bNthB/qyI2ucSLgQRdbtj4hAroe1vYiP
h68sOCnDhO68KBZvukdPt51yB2KlExejwlqYKqH2k2zag5ayhm3vShba9Z7hCyxK
nn+ulMrbS14jZozK3F6jX82vkoI5lgm0lcRlufehfNbr7xzcH+IvYGmEkIJZYIO+
ygYQBHR78HNtCHrbHapXY0UUljTfcLMtFz5Kf6UJYoDKKC9/j/xR/I047mmxxkLk
cfnJiZ3UZqKzRj9HH58nmspX9XVKg3WEByOtrtkNLOEK26mj3iXIg4E1v5nPpGo+
r6MEcUwI6t8LgctlKX9SuO+KF5VbQO6jC3ebmmL2i86nIIQOnH4Umnw0siKjqtR9
/CD5C2YYrBx7A6IX8bTKUBXceuFqto9922DU1X929nFJe07uN9Y9KIn0JNioUb9C
tR41qZOx5JdJGEEGctzSznftiyUAT3VDdEplngtGRnZqcs57rNQNlplbMGT7bU/T
ZESb2tzArnW55dlk+izOsLBUaMJFtHI3Vz5nKe5whB/ayA76Nxrqjc+zdG/BXb9+
O22hiv9UjMtVLbSnwWS7uKov27ehYPvW+mBtHCkYBb3r18WXS1Sponq8jlrvsJwN
kiNIoK5ow3is8OZxkxbJtzKz3mkOHTWEL7HmtpfbUq2yNWsq+Zs5AH7/12st8thk
KGR0wQBrIf+EwpQ/jCQyur2e7AqX+EDR/9k7GqMQ7IVm6p5SPBzQyK+WvbyZBI+g
AlvCtXRRwT8L+UDlaCMlNd3ls6b+rXhgvRPR/3qycYG/Z1T6oLntJJBRCKqfL7VO
xefYyaaqAchHyS9xxhxM/d8n2zADjz9sLCn+LnG4jk6Iwo2ySgm97DgMvK0OBdg5
1479hZHvaat38R8xqE4YNphL0/AovkfHY2jIbadyZvQBEtjD4duNRpbObU/Pqaya
qWFtu3pLs7n92BjMVQvIa3s8BPsk4UY+YR07K1GXa11hcPB2WzvZ91cIL2kFtewd
ldlYg+VhuTT7cXnKjw+0jFj+4HnC7qESMa+ysSIl5SDF5KcYbgdEf+0OlKlEnnNQ
RbxlIaZViLcZJrP2xjOkP5oxxyH/02XAJzP5QUAEHw9xTLXEWVOaaPcI5WlBFuaf
g0vI6cYzr68FE+wPEB6hMDxNSJeciear9oCwCXPDJUXXhVDKQgNpz1Q6Ecy0911u
X1FewjANB6+biNeIqeMz2ZGQPwfEIrjcaVW1SKyXBlGIyZIdiDrW5B3jEoivnHYM
+q2oYdmMWTcVmk5zZeRp3/EVCrsAaNyVsn/mkoElZ9VDOVxQbIQ/kQt6MTmoKR4j
cZRmGouU6MdYknfWZEecxJNSC5qCm3SuZtUZbSMjYRHF5eTHc01bRnXrwXChCGi8
zoMwFxtNCwQdH9szXmGfR/Ac7XQHodYrD8o984Jvjwev4oY36kXRnDIHGUumJe5a
1Tb9gKlH/MzVOF4AN1DWLNXb3JUvqlI8XyyCCTSVVbQ=
`protect END_PROTECTED
