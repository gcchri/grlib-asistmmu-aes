`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yrKjbHuQziTie+AllYFyRH9WxVnUMYx6kpVFYVjBHnAQzA8GmM9w7clqhMh+3QPB
LkiBZsPtZkoI8BVTdUmfSKzBuB8ay03BUgi74KolzY5oWHenoG7L3wGomOl5V3rt
ZXttlV9OlnUmN+OPyP0ouvgdc4wYksXtdB2KLzgkZcOq2EeDoIk/dnPMO8z3F14+
2Na2yTKvqHivwlxds75KJViUnWgO8u/02PFdAwm+5n5l39C+8ieXHeqy1RymOKpC
qZ5TLRePRyCfT/PIR1Dtomlh5WdG1v161KdB4pIXvQE=
`protect END_PROTECTED
