`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q80uIJNI9yE4YA7A2TzfpXmiHzpZTULeMBgzIhp3AsEeX9/LCnzfiWwrNTJ2JM3S
hOqWH4epnbygA/HvehySweUpNopnC7fGFCdoePaiKc3ZYIErBlGF7QrBiQL5RfnN
Q4DNCdRPl6GqAMNaZFa30slSFwJEZO1tnhwCGjiXspwB3rTdMjZOuzKbf2HRs+SA
i/ja2OwEBi/jtaPuMXHKhLi/choww6J46LATBRza9ooEKvNlrBCPwctrIOpoiBNf
XvP8xFQ6I17SBlxj0QeiYMXzhAgUU4iFBdtH9sCqVp7zz5fHwlfvlW7J8+V1xAsa
fFYdIWRhGLUrSfrUwW36MDf+C0/5/mey9/4uE89fiqk=
`protect END_PROTECTED
