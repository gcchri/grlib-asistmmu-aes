`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
72OKI4DAXBrMUhcnXtT/u2NK5P0IgFWgqib3E3f2ZCsJItmwdcoaoJnh5AlU/nK1
95Q1czGAIH2Ccy6dk1LR+MYXSNKgCggeHOIalk9ZFV92EARIyquY0ZRPpi4u2zHq
CpRldAh63EN4AKqL7XGW8PMKwFNfQ0DqhJEIV7GRqOQARb2jVc3AdN8HjTayh66G
LO2t4g9iGphKKWb55Wnwud3cDaE/SGU48Wu/My0DliN7/jSD1ZbRcba884piD/8R
gJDGq0LYpK++BiYFUbXtFX2oC5APcv8Ti55fwqI9cf73s44idrwi2STN1u7ZMNMS
vT0tpkc92+SH977oriwE3JkYkfI+M8goIvaVbyDpt8pNxv2v71qH/Ud1K7ptRgln
4fV2BmQ2fz4zLQBttyS89W+zgkWGGGYuNbPqFzUERI1H9chjASU15wMFGRDMHtuG
Qm6iqCeDKHWizoCiHoNWaHQWf0NZ/bbWHjXVz97mKX3gLJB7P9bZGdw1XqVPwSx7
kYnuDCcslwSVL7Fsr3Q5siVvECWO+kdW+mn3I1GPenWh3sqUOKNt0aWmbO5OLboe
9TBTya77LOhkrXqt3ij26c1D4foYaQqOr+Etje6ZeOFShPr54svWXjf+vbz+vzKD
cVg5SlJSoOC3OWgJCKVuF4TpI6Aeme/koXwsKMNqmDnN8RRQ69/6VerjqpKq/Dmt
76vvJdijLiQDd9p3nPB/8j/gFQ+THeZbVj+fJKkh7ZMGp3A3m2F4X76dFwe7CsMg
bgU4V5hKaSCOTxGhlSf4i00gHalKTCdWEn/zgC2y067lAsMtnhcB2o3DQfxRpjam
SQhLZ1JRQSKOmDrPNpuYKyI/2/mEKXITSh+bvN//e8987EM/ZS9/Hq+cvpsFm3yq
zoj4hCH2LCBmbebRmj0JNZo4Gma5w4CPYxW7NwL8TzPb6hHfxWBxzozf/8E6t0lA
jLk77mmQQxLcgfBLqy4vzcRWa8DefmQOc3cL7rnlHbC9bNsIIoDTp0m0/ju+gAR/
ovmnVtCQWe+v7iVcbe9+0q+TXY/BOUKZw8taFPeW4LHRHeRI1yMGnkjwnOvg+rNZ
vbs+TW15JqMD9llcviQUCSYMUDEhkH064n1YsFqBcVWibTOtXUY6iBXc7G0YsdiQ
tS//PT8GabL4n+mR4YaOy72MVMK4Cx6EeYc20dHOQ+VG2NkG8fryQdsyhkuVcHqm
j36sa8Vz4wt8dWFRY8prTTsZL3/d/64gnckB73azIMh7Ar6Vw67LYo2/gj1JGIGr
4is9mgbcC4hcv5qIDit5NNuR1aU5fFlYfW2aXFOX9FK7XtNCoRACzr9QGcWsT0kL
V97cP9f1kboT5kMP+tPDQRH402RJM/EDM5NO44M3K0PKY2K1yv+cPkHJ0sjsYdid
ajWno2kDIhxq1LqEmSMaYAnVKcaSV8/6f3N9JQ2vbrh5A2ByS5vPVmUcJUVwbT88
zp4/9sQQvOIdrl006u1W4aFiXOeOb60rvEdAl3IDcjHhLD/qS0I5vlWO7SVJtBlI
LoA/My4ShmkY8xWzAyy/pnCnEBKf0TZRi14T/43cQiyQK5mpKB+iZ84ft08r7Ej8
5TruwHMNZOZzGcl9SvOxEgESINCM2k6mFhm1/sP5ApTH7fCxZHdhGjXy8SBvIylk
nD/60b3Un56dYazyAIo99wt9N7A2yjkImoshRju89rO2CCsTiKuMkMTEdtdSZtn7
lPALI0gam9xvNl99NIht1IkHWJ7OUrqhURiezGeb+XQsaT2HpCeL9FIYvmtmgVwm
LlzpmW91ZyVcoKJEgz5LI4gH7E4vIexImnWkJcMOChwmz4je3aQBGjAIuJDkRYZU
LFkU5tanxXTHHvRzkZgN6sMUqJZmNCQ3HuAK5bd5ERK+7BZGP0pQTdRD0Hwpg+Ua
r8M5hZhSFQl11tikItRMHPmnf2gOZsblvLnJsY0c8IPynOaxx7Dq1vaPbU5yowSH
YPp7SwrvDALNWnRx70DXKObHIWZlO3SsDYMKmPwaA+RKcsy3OnW/kAG2SVu3Xvyf
F55yATntWuFUG8iVc74MM9dQwzqdnuw8PqI2/8/OH6TPHxBzHSNNx2zIGSQiPqbK
bomFosT9XUss+X3PiQXjZMSunzGDgn0x4EZjEQQm48MsWCxNlmPzVoDRS9orhcV9
7eN8Mnv2dmvzc5H0lRgMty1B5p+45YGHsDpi2HgNghkw3A+rrhw//hEn/x+BO1Wn
o6kZCnToigqNyKMf+rhsxMItglM5xOdVfpcHyIr1UJh4CRNj/syPq6LuWe6b22on
QUqiFY14cPqFZ09TYH7IHH9PiP6Ra11fKrBB3kqBI28TnnzPN5hFu8zJZ0sS3Qfg
Qke1UFzWwiEFgXpI+wkGyNoREF2VzZ4pOTWRuetSx5L9zwP9UI32ESbXCO5RjCLy
DucubyendkSimc0oZzfCWwRNnkR6eZ6g0NAzRHL6cdDQj+EsEioV4D+v7vG2+qey
mdNH4tOKpaGtZg4NLWap+0VsjmBLs7THADvUwfazesJnvqdnGv0BNvW95r4/1IOB
6gCpBEC41Xxs1MRKkYp70k7b1TeHbARKnRDOPasvxgGyR+wC47xDsEOn1zpnpK8g
oCyRJsfP4VSAOMwk82sMxN0ZujwxhhQ/65ZsTwauvvc3fI3905wDrkAYC/6qaPIJ
LK5+imrOluAyDHV8NqjoJvFCxXEOkwiQ8C01e8LAUZ9tNnnprG6+iZfGJ4EWIxRg
cb0W6+K1hTDmu/SAy3Bg1cPumahUuv1jvSyYRWsCyDiXwNpcHZxTxzz6KDfDR2CR
XgVsXL77sFP7w4e4v5WRYEk7kA7TFTRRHloNmKSnCp6w6ixQvOdusBbdFlGIEQkG
XCTegqo0GGlSEgQN3AWEsmU/fY3my6vkJPS4MpK48qsjXMHHjYkHnToo1HIh7Bvv
SAnZCzD9n359BxhV0WvJzA+xNA1Z/eH6KCQ5KfZnVGJHoaV/u3Xz0J6PE3mLJimn
zz5gNhPq3IR88BYlDGP3Z1XoLXzc61Ks/pzab8V0YmaB86vNrAvnJO/18N9g7Ix6
i2q+8LmM0gWZh08dV4jGRQBBJq2ucv5EAguaPTdVARumj09CpMXVVv4vaOcB1MgL
fFT+NDq1XejpD602YGRFFH64Wh/M1PRE13glvQIb02UKFQ8qvmER3G8INukdHKVd
9W4xID8hbB1Ve6/jo5rNxpMUlRGVxCL13RMYkkrwTxMe5iiHPd4ZdyMBO0P55hXy
ddk4jTJC+39h0x7qUe/jabhtQOxsQEj89D7SZibcJBUyjmfGRdeJkdmdGo0ybyB0
JiPerAlio7XgSj/eRFedY+hkp+Lsi41f765D6WdEr7S3VI5mfz8yxaOLBK3yAH1o
9vCAyWFrKs39Wcg/gpJF/ZvVZ8XoZkwR0OMLpEE2MlOKfMCHEBrBZ9tNvCc/I/AS
rtqjWZ2ezjbF8xwTvk9HMTg4Ipdg34N8WuIdhDlOGH0bQ4JRyDm3kMk89ETjnTBp
pN07p3hmdZb/12E9Tvd3Zd5rOrF+6fU11nFsmAHj4SRBBrNozAhJlJVS4YLOkfHr
JRycAPF8zpgQFKUrAU+Rm5aH5JiDkXXG05vHh+ZwMdyhKT/I+rC9D0fcSYb8is0K
480Ab//Q12Pn7Y4z4YmbwGffuUyg6f1sSBewpaF6XqHbpUMPI5ICHhzXEeLmlsAy
yhDg61ht6NXw4HVONi6PvzwM187vdRUAFGE5Qb740/c6NCjo5xBwPAr4tt4VH5uR
j2++WlQaFM7OKQKB9Ho3b2fnt7HXX9fTooZCuZjtqabDTQjnpIKekVT7UsraEzGE
zCMyi0GM956FKLm/9CW9uabwwmccReCUpJhr/8e1U1amaRWDvej+4T7C+wqCeDEa
22D5xkK35mBl/5YnmvsvLmFjSB+R8ZgSdyA85Cid6V8GYbA6iLTkLTYEYlbMTmuY
F08Q7+4yoI3o9WMZp9wXzG4uc92RYBi3gRf6hSfRKx/Gv2mRTsclx/CPb9Kafl0/
cdLZ6BIdgRfwDbK8OdmVck6WViJj4q31zT2bx2sRjbNN3vbW40TSbupXEDKA/O3C
YuJWDhzN9M8gAttQthx6zuz6OSZvofghpGO3wJomai9Yfk72DCT4KICtbtxGYoYF
Sz864hJbwXxNuZBLYGHEk/5hLZ6FH/MDacqbQqw9T+WVjpbSxvdMvre2bFWw+6XG
dlrdgFlvc+WCcDMeX0VgrO26aHvyMvgKz0pXTsNe0qkRC6YfCMWVI3nw51rwnKzW
`protect END_PROTECTED
