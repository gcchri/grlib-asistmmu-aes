`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QIPcHYsNywWg/WTYiZOXqr4Z4vuu2OyIESpI98Wp7wZ9fM3P6Qfmjsc8WRZhN3ym
5U5uL3jGMj5Aau0kDjMnjguGITmbZXrPnul83bydS7s7Q4cCcypq2OU/o2zmH5DN
KV5uIG+V516t0r9WT2e90g07Xdp66zQXQthCn87smaLJkT4v8mjlgp/qCOoZlIyg
26em1wrbnhzSnHoagMgp3Xgigx3wVKoZ7A+Q4uKZR5zhf9ySdHOUNMZWvcwqT4uN
CfmX1UOrrFonsDAzsdxJwcQoCnKUq8TsvEBi9prTU2eckeY3686BbbHPk8l//4Gb
LxTc+Sc4sV9aWl/838RDvgef/F46wJov3CbHXNUrk5SyWMCi1YGRmL88Erdn+iOw
PEBk+uAX08PJB4oRf1+lU4VjBPvU7GfIyZchud+PJvRWtEvjI0sZlAaLsOP5PspH
H8J17NmptBMRjIqu69ZsmZNEJPg7Wl4mslQn2wVBIvtWA1ZZ3xy0zEEkNcKCSGHa
OdE/gTTG9IXEGogE+469MnhcvrfV0IEH3N9ZvhHX2gn60wKt5wCcR8cTwaR5VlIp
JknteWcSW/5BikJogTlYOl/UFY0qsgaX42oP6+2F0e/oAp9yLxbOQY+ND+qyPQsE
EBwAuLvblRIJVso2/Qg9J30sm91yR9SxhxsKJOWF7h3jnbGYwBX+mHc6/1GIXW6D
cxHfEjQiB+RJ7U4Px07yRFjrwnJGFVMUBgqhG3NlADeTiZziX89HdyH5EGWwSibA
vZ37hU1P7OgxcNC4PQYLF16gQfrTrivWb00QQcemDoHW3pIzjIUlMEpgyg4lq8P3
2MQ7z7qqIEQpAjjs/yP9DCVn5xv5PyVYFBZ1g+TTw0Tap4PZR3FzHZmkIKKt8irw
Rhww1BRFn72OWj8stRg91O5WuDE8ZwZCZPDg5YtuusdFJUT4yF8NuBm/mXjmEbdH
7k13mVszJZLJ28A5Q+vyE7J//5Zp94Xtp1YCsHgsb8r5RgLdZwvqWvHsLqrdvCia
xkEzeRIKvGYjdeMRQ26JDt6On/yWfx6XfGjB+LmQ8CNVkiY6FQeuNwn+51r5pX3J
W2ErqI7K1O4mBtHkwEpdmg==
`protect END_PROTECTED
