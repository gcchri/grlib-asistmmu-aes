`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/qOqIeRclHNssJxDb6dGeQcyHU9as1Vi66xS60DFXEnNeTLQzl0FraVzth9NvYU/
XH6QYJq3YYzg4XBasJd+78sp01pHuovSN0vt8t7V7lOGuAcxLUpOQMpMOhUyZPsK
tftZJk9/n0PBH3JSA0YXLH2RAJr/ipl1+e0AozKdYsir5WJgDZJ+SQzb5WfbGQ2K
PnMUuzk+MRR1MR4iTKZp5XujqfSYoiPVDHEaQo9XP6IEK5sWJs5hcgLHiFTWifw0
SXc4wfBDQnErnN8ESd/1WYX+DXdOhrj4dnawow76urs=
`protect END_PROTECTED
