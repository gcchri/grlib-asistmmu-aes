`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qNOkP60QYgFWD+BrEf/4J4tNKGU1DDwCCoecL2dMXgHqNZeT38aUrlt0iOjV2koM
a6dEYYcUXvZcLy+M6fYXenDWUJ+QmHNIvs8nCaLc2qMYrxSo+29K+/DKnZTPpKAC
uNCvBoohWcJJxLkyScnXjYwyR3k0zy1xnTkaWXYFiRYY5oWA8mRIkTC15Ik2/XCu
9DO0G92/GQTtTI8aw7tXNv9SIWrWgELWwEJ5goexsPa5GS/XiIoB3G7KjHM2LYhx
6hADttVqjHD7tjXBLADBN9SDS+ZDSZTo6Od7QkczM/N2iJRGVkSUWBcOzdy4ykyD
xCrHfq0Zwy71ZItz6nNoGA==
`protect END_PROTECTED
