`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FFX4RFgHHgVS9h/kx+2c3zqmmSRD1s38omcPuteSsiyLJqMl3V4r4GOP5UOcleXw
k6fnSQG3aMr1RLBBaOObbv1iXTtmZl3X9vPyNMoyKf+3uhUgdofVug3YJlP/x3SM
GKpeqyIgaJaSMWGzC0vR6klaLsL8Q2NsTyRxhFLYJ3Dz9sUq3fdUHulz0+RbcZZx
ElpgN47SpIUiekD/OQN0VTlY6w12xQbjCZxChm5LurUt3rRJipoDiGf5rGnVG2zA
o6vZwD7Qn+cM88+k+8Zyh9SpDHHP+gH24Wq+jW8F+/RRy0OrULfSR3o05b64bEyG
d5jOLEXB/hJx8VB/KAEmET7lZ21tieAPsy2jx+p1MP5hDOEhQrk2R5xvcTmBHZMC
nevgbIJupczF7M5Eo6Z+43U+hxuafmrdwbMUFChjemk=
`protect END_PROTECTED
