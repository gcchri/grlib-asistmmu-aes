`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o15NbB5fetzDY64b+NxlYfU+1BLgXqQKxSsRiZki6xE57Sl5sNxh0DTct4rpyvwU
n46LcBcPsY1LcMfsRhPp17Aj4gT9BKbUQiMx3trACmQsotitu9nEilTD7p3fYp/t
DPsk0EZrEtCgjRroyk611GLpIV5KjHOHylXHMqM8EIHC3nafrB31NbCVujxHx5iE
CotLDL+GTAiY0baZ2sA53EdW2JAJYqyZeL0+KjvgmaFiprBj6P+AKmIkjO224zcR
FZbGQmgztgWrl2K4LnBAlvvDXl3Qvpcm19He31fjwRT19IE8f89qChWfhRumJ0nl
gmqvd763NLrWaSeu1QpreuuakF3ClmW7CR4mqA4tCefpkHyU2NyMIBIDhWdTns8T
FewNfJdLfoK+OCKrWXF+YE88yTWjcxagD/Ql0jNVZw9P9PJheZP0c/Lt2xLES8fP
897zNdv/wcjHru/jrARdVoZNxZaGx3lVLMkW2QA4ub5bETy0rYQ1PWWBe5lUIQbl
wD9yLa/vGWYUCA4hlQv05/XaNZLeJv0lt28GK/0vC0GQoLsej/4HyPtyfrHtNC/x
vaoIzkVEQrEvvyyb3dt2LxQ31GVtlXjJzLFnnOEMRKR2ya5Piq6kCQEGOJ+XHQ0l
KuoeeM1KcE7CaUusS+mSOBO1W0qpFzRYPDzYuIHAkCWZ7i5ir0EWjj+NG0E5TAqf
TVKVGgTnl4z0xAxZ095nANT/8YzrKOSmzZJw/6aL/b8PeuQM6eCCv4krizi7PlSo
EjIOjvX2fw/Usb4XNRr+XmN83CC8WqVzCVDE48DGGjRjqR89bRCBZkAVi1TO5Zzp
/DbCkzbsgFiPHNkptFkNmnUREkOXiTjnRUYul4Z2iyo=
`protect END_PROTECTED
