`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0y7AMJNA/gM/UXC+nEEOc1Q2SUBL/Jnxki9gbliuvXlf57WqGr87F4wuDBfhZ/Dk
evsVRLLU3q3Rso2cALtsybBJmh7Q2pjpazCLUxmYI5PBdl9B3LakUqkgAkS4ZBNr
hNyUy8/sbJmVcSNrmmRz7ZNGeM0cW8Rlr7HWCKpqBHKn5QjmVUa3avFotpumst61
6ZmTPqPthjbhwasvx6AJkI+F3UQbqSExyc/RbujeTg0PvTBZp67d0Kz1bpsWiJ+8
e76WcB8Gj0dSyHpXwcLcdhOFIAOT84sYBqxDB4p25rUzh2arWBSQInkujzTPDNsm
a+qYyGWz2J3P4NVAP0E/2ys0MdYZY1mRyxgSV7+JRFymG2T8XJYFSDTnBk1A85L4
x/92Sv8pK3jt7EQzJZLq5bemb5HUnKJa4BFUv17JrUB8CEFS/B5YFTF/XQ9fapR2
zXCwDOZG76jrOB73kTPR/YlAF0gZSNawTJGcGrQ1duROH2n3EVn3gW6FDRKKcodM
wzjB2f0UzNjhCkAVch61ohgEGXsj892sz/Sh2oGdiAvVYSIHR1VpnToL7OcsIRoL
l8gtwaqctnYKWBYLtNmz5drHFB+JLYraAOsjIPnS0nsqPOvXnRBCtv7smCiA01LZ
`protect END_PROTECTED
