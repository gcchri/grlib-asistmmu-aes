`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PKwVQDCVEe6eOli3QvSNf4kJWlzpK0hNgeKLEUzeEf78qgq3tAxgMmcV8AZxhrAN
5wc169Z1wbfXibEVPRZhr1aMKFERzh3uNxILUp7NlSa2vwpC61SlOQHlj/6Aeb3/
j8YQJYGPj+GK+NsSkXPNIqKhKOnPILqLpzM4Y0CV3NFqICSROnRhRIi3kr8D1ShO
z4Ba/KlJbnsDcwzgonjfKywy3qkPw/ScyylJeNz3I0Z72HdiH5S9bXwsOMelG00D
4V/cIwo9ddle37+q5M9kfy5ktTT7V+U1tKmBhNq8FVqI3RHvuDGGY8GGtjZSZsQi
oyxUlHARAa4eIHsmEueEVwz9tcsihpLg2Y/xlpQ35AEJ2t5Bj2eID7xMH36rWbce
JpvwrfMq11UqqHuFZS5OggVaeVQWAmHPxEV+fqJ8Ji8xyRRtLANcKXeHui7oy/iO
Alug3YM2lNEkBNbudMGeXFHw4hf//YLhD3ZAlThK9V47h+7+s/45T65znrcnGdci
eBc6MntgJhBusMgrbIXkPo2X/xI8wZmNH+QSyI8Sr88HR8TZM9bU76GhUV1HzYEE
gS3+fNzvCHXu83H+/WXPzso/7jvC99kp1QtUs/Q/Q1VzW+JNnsWRZlKwhNHU++pN
MV3P4UDzqYGnthmM1X2Och3IUqKa+TztG1n/FzI+DX66UeFrxz3hF9I06RZ9EAZL
IXPSivpm/rkg2daiJAbBWT6jI+1jLPj5VNL1Sn0W1w+fBSqhtFdIvsT6+DJ64Xou
N4exSBqmc2oEZi7P4VTp2mtVP65un1C1q3wQEYbO/GZuby6PNW4JA7pS0V6SPhzd
0SHTPEiALWwa6fVuvRX6SXql+5xeMB3EwJgdHfkRFF2mCe0vsLbnBkfvHm7e/tpg
eWG5dfRnME7zadaCOYLQObq9hEqYx1cnd+chfIgQ5oiRFzhbUrLETE0Q9yyjNUo+
GSlg/cRBMYP89DYq34HdMsRzL8tzol/YjpeQUD6ctm3JO8gYfqW+xBDW1lFkXDTX
OSOR8EvUAhfNFMpqh0sPDQ==
`protect END_PROTECTED
