`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+nEZii9/rALJPXycSFdPfRxpZbrTsfRBoqRN85nDenHnSPuSglodI23Urj4lmuyh
EjSgPGHSiZ8LnUPskPjJtAczF3M/pJMkeWcouJwkkEGr0XohJVE1Iltwsct6JC01
iBKXR9X0nVoLFocgkFZct/cqN37QgX5r2Tn16PkDbhYKtrN1QmLWmPTIgGYthy+p
0jtf2m159o7/77NjcYsrO1Rw65lrDC3SeOyDkj6SP/W9qb2F6EUnkGf23oPWw8kF
8DtAvxOWEZ28LqDqwT4MK4QBrgWhbUK0R1Q/v+IJXHEkt4SRYt89vN9tEyy9kplW
xLNSd7O1cKCjNjZ0rU2o7W3y+J2bdYWHejCbJnMhDJ0mSQS9bJ2NFtBVCLMaNPoS
6/N5HANGWHjyZjpcUrd671y48P52uiGUx/KiRU0ne1YLG3dIJjDQSRlgR/U/O3TO
HOFQ5NHqbpqzDfyu/fBp6QI6jgncxCQZywhN1ZSh65XKxVRqgFvpvNpscjK1Zt2/
3eZS+uOBvId8PQ5yR2mLVALWYo26ODyuxAkvlf11vCzP1rxOGf108QxFUZvgOACR
jj/9bZm+FFyVwBnQ2/KRCKVjzhWoPksmIsvG2xH2qfOCsQdcIXj3KSajXntKLlpg
kiv57uhECwS4iwwTPvvx7kFgH8gjG4Cfblxi6RI7gWgPJc1HKt/x9R+zSaS5xpjl
umjU7Iy7F0rd2TX3Hk9w0ej20Qk0n2yqZhEyDzZwbk//oAMZ2dBHcW8cyClbEE49
CVNDSfUgpg9NH87c3Uu9eP03hylq9bAP5xYhaLtW4pd4y7EpXCzfmk5GAbk2+Wbk
/rG/+oSHetMgs/pNL+VWZ9OpLH373fbP6YtAgsIqQ1BG7u8GgXfW8COTR0prxPHN
NeXfF6gxXhi9c+TIy/2B3fm+kJRV12BkCYOPrr97FfCYvy1egdwvNPsxQ2XpMCGt
j1MIe2KG/pXL1NdhlWmrZ15gXQuTIn6XAXpoiluD8HD7rw4ysIbhOkQD64HXAD4k
NnBufG6DmZNoQ1ncEO2ZaOneO2ZApeH6Ie4PqiVNkqplqrF44bqigJgIHHBCR0c7
s0xWnvAbQ8mkAjg75bJFG1QR6yokGCLSKfTWhhIxB+ombTaAyOhWfvXSxfWIIL/x
TOtJvYIXdcVqqW+0B8KtWBbGLlLVpnc6Lp+vMG9//9Gv89IyT5snnd6jMGEO//UO
4EEsu6dNFA2C58ySaoLTQbIlMut8fabGZCk+6ap7g0fMYxH7EN9zegJ+JHRA7y2L
dYMY0TjEnBRcrQhObbDn4wBDt+sQItUmz0gxUXjY/+V+Hmj+ajgIk+9zmRhxIeSb
kD4LAR6G+GKWXyZl+KyByQMfiPOD6u0RTKDCDJSJvvyVM17b9Wdg5wrn5OwKLrL7
NdG7d5lLEjW5tb8wNqY8o4xttNFXXnCFSHQV4qrsmSH1RTcxHbmBPV4bSeU/468f
04TdM000VzsmZFL+sDT2N8qB4pdwWP4Tp6W2IvAFUd8+t8hp8cwXZKnkPH0lQ1pW
gdGXf6U+JGqzVXsod/9QqLK+sLUweZ3Um9I7qd9edqwI8ewcCeLz1KXe4D9R/Y6P
5JVODRurawIAK38C9zKaLfQ60maAQlO0pZuhmhQVf1NO9kVvKkDKcxmFJ0AM/uYd
Ot3gVC9JFjP+yAZBPs18kNngOeo9jFiZBx8Wq137SHufpetS1EagPSWYu7t5bqlJ
A/yXkimYHnImFfkSNpNMI27RiWAc0jL/wWOPQqO+i5ih5mrNhbijnpJIH+j2llUL
Nl2/xXwDSTs+xrOSX6c5oweCWZYnb5BdZ/pIIZ7MwHaF3N7qgG3WP0BQ749J6iPv
i5I9961Krxm6RJ3lWXhj+w==
`protect END_PROTECTED
