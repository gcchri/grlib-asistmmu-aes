`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3mJUNq5Q1bC0UCJAiewtvpjWWDCVxuJGF1VZk23gUE5plxewMLtNXeg/o13BK9Su
w7pCZtLhjZmQ96PYk4NwsLen90GGQoELDBFE2KQK7HuEsNrxsYg5Z4Tum2QnC3su
4cR17yqJNLpCxKZmB5kiogDEWHM/P6Ark69hwzRCSCIUxtW3JWM/HwjtiwNGGx/8
L1BG2eQqw+L1QYXYUnr8tNwVOgEgmfbIZ+9csCx0/BAribXbrICdz1qESBXKXmXK
+ZkPUSfzmTXTHk3loh5GD3WxIgd4nG3cg/d1VULebV+E9ht0Hrf0P9/FtaWGJl5T
vnMs3xgyS7OwR9Salf7Pw1bVvlisuSh7GVE13tzmSUo0CrWHuIsYnHUpVEEYwKqo
`protect END_PROTECTED
