`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZpMWReLS8M45D3E4SN6UhlNSqJw/JE2CA/5U8Ajh6N8n2Pb/iclsHxY4lEFhiM7p
vPfVdbrX9IkxdTZ1Jq0tIxvjDoHv+R3/9A2nwp9o9MlfDFQCSMaZEELFvg3akM0o
uyZseruBxPVHC0UkyZif0yO2DjBAcAxHKV2e8mtxo3FZUlFQrY3fwM8ekqH92WKg
uD6DcT0mqRkpZSBN16JHrIeb/w4OmPiC1JWaes8dFRtL3xk24pkxs/4twi6RUxMQ
OeEfOfkCnr9gipmtC1Te7x20sVk/XOV7I9Vx0fr6mortMSxXCKeE2s2o+XmDK46e
lH3OnvRheatXy1WiK5gdz/cd2gqIZdy+GvroOdAAR3EmPjD7C2as4udhkkXO9mOJ
9+pZ82UBTiglI73A9oEDr9dr5vRZG45XURLych9TTmbyWXWByXYMVBRy3QvkECyh
jiNfm5eCz7NXp7VIOypqxPIJK5aaicg4wq/nR+nQqcrjFNV1Hj0hn8ITWqc633LG
BbK2WGq1cAxLsIqFl1kbiAUbc6VnCPYvkicYJCd0G6IP1QJVelByCsoeYa/PMQE3
QtEZNOraXrFi9fuMxs3SX0T73PXX+32lxFil3ngI2pS2xSE5vVZ8baKWfk5YLYU9
QQfoLaVIU2IHBkkYjKLNO8Ugscllp5iryfbkpH3J3dptQtwkcFw1tuarzlFCQl5a
HwuixQGMiVUiLWXxAMMp/q4oRhUrgrNYnyp63FLQi6ymHGw6LOV/0GMXsKFFMqJK
R47LILEBSWRDZjefCjD8uXLRbcSR/E8vXauwY7Qv9fHtDT4TmgPfK6UG8+gvDCaC
P5FxHQma434yaQsdlu+O4PTvUPiPvp5Kiu+msXF2IpG6yazTwQrByu8iDLzd1lLq
705pz8novd7jpJeWIuDHfqThU7C2WFD5If66Y/dRiYo7oFACdXlou6C789I/UpAJ
gMktBVBOPLNnJwRq/wyQek9fnpAQw4iXS+HIHLz1+KjRaOdGP0S2k4BGbH87p6jE
bq9zJaJJMilvz1Fr60bqIxIP3bHQkTTB13ngqEpk+MLBzfoPSu5ZF3OBvQt4l/yW
ilMYVBkIe6Cj1bMGGamzbx7WFkVu12h6FnZFLZFXYOGO9U1zs8QbporNlrf+bG75
uOsAKTHaUDuENOtoi2iZ7cpGtJssiLHCfHUJ/emO2ddewu1uFXOmMyE98u7Dz+aE
aTvo1Co/0/vOpc3arWALsz3U1VX5fdjyRuZ2RFCYG3O5LRQMzfCj6tuxG4HoSPln
7gaOJ49NDWqGwAyHoOOpkylxoifChh7nn6iMuUPo+Q1hk0RW0BDFkEQEkXiR9QRN
tMunj8e3cvv7LWOG7UVlprxj/NbPHOcbwdhN60En4QjC6dwxSbOF6hsUcOthAhIB
J818h/+ivxEAbPpn3tW6LGsjjhvoYaqMgl1nCU+jOjzi9LxRWlenxw1B7G8mnk1g
PUg7FqWd/fUCo77UNEBB5ju8PVkd2htaHmmspqCMN7Nbekw9uS2QNTkFn0waryET
tOgHtmqZepC3Zru6ex7rccRGo1UIeVzO+DepBs1adGq+WH5l6Z7ioUERoGmSrQZ7
ibo1CCodxsQfUJQnPHmUrUS7vg1hK+nlNkHNW+KnjphrVi30kEwOXINqPahiGzV9
5eLvf7AfyHs2C0osBUFOIo54vtL/vlYiR66KJbawFU0Trac91k6BNh94GFOKHdth
Tnp2gXGDqVlUMZEYM2AWsHECAFkkGePxluWJMw3BqPF0KkML1DDDx2WJV7OLM2FQ
k9IKU8ob1U6AhxIVf52yRTvCOUXnYxJrI2l1ASQYmd8l90U2IXEIOMQgKmlG30Mh
4Y1+IAChL/qG1sI8tvOx09eCmKRjMCOdrb8zmGbtWwXeEFFxAPwyBjHQZSDnhEVJ
1fJ4wXsbHx2jfe781963t71omfOQZIKg4LbW8XsfdU18/OQEIOPtbqaNBLfZZue2
SWfJwUhCnvZ5XlokytjhrwFVO4m41jv1QVAyJiYf9G8ifb0Y4Mm7PfrZThLJujx+
/2Ji3mw7GJV2hzKXn3Qe+fSC8//vckRHQKZX4EdKKtG6mUWvbKY11rQJ859edQZ8
r6flLyTGsPGrxXUE78Bm1Ns0u2nd9zcH02X7d4qFYvuYU+jzglfdl3xUteL3lpCd
aOlwL2T6k4D2ydR26H0HddHtBMpKqu3oGEgAWNrKHgG/B1BposjQdn05DqtCpEXO
wBU+7iAGgd/SFYTQZf4R8JEexm7RpZ/v0BwTiHxwQql8wsJfbPbhhpWQT+JYYcnZ
bgVXqGY6ytT3R7LZMRk+K25gS09hgQit2h6Jeauw/aO0PEbh1eViQJEvJqhJz7rp
rDBndcE3wMLO+3xZ2GLW4HRRgWnJbZruGJA8GB0c0oT6fXiKOznET//NyRwhvobM
1yAIxjLvkpUefPMMIw17T9hmMDhecqoVsJ5vw3YBtZzJQILpi/G0i5aj8xh8s2vZ
+Sq77fzneCvtNTbhr3UQkIdXAFaUKxBqaRg9SXW7YAsrQKJhONQadFdgOt/zAdnq
sIwz/UIgRXZ8KBO48F00OX+Ufnq+HxgvZ4xkD6kibMB/6gFRCIfupZhW7ORVQPlu
wDlpkFNQrfoDPG6OXJDunpB7ElRd+XN2zZaethKrJW33ZvMuaa9KsKxgGENa19Iz
aI/FtLw+klLzk0Jzfws9zUQU/97jJfnjjgKWbHQVS473wHnWn86zC3ys6VhwQcP8
3kYveeCgVhg2aPq3o1sZJm2oF2OYvDlPGv3WmCu4btJGrAF0Rr3X9XqSSRzPdVSf
fTk0n/2ymzLKhgL75b/HNdY7e94hFx4PNBOKiWiSbl2CKzY18IEYI07pAFL+k7LV
ndqH/zcp3O+RIcwYKL9DvM+x+HPhtAYn8r4mXxE5zdX8cCWmxV8TiLPYilx/SftG
q43iGb6Hd3mQkmbYFPN7OuGFoUnQF6Zwjw0O9m80idpTLiQWcTSb54yQQdH6/gOh
oTEU7CJW8p8wvnjzy86BuC1HPtOR1lm6Brl9d4vD2QPFEpNxYxmVObAeC9Ync1x7
s3FyMs4Xlw1C+cL+aikAc2FS09pPDaeXTIP+z1vPCKYCWXGO/rm0rnifjcC/D9R4
zVG1NBeAqva4ojm2YiS5tqElFd7ztIPMS0NaRnQ+xgg49TBlHM4qUJRijK5bxxGP
FVsCdEjI+FNnu1XLmt03WIBhszReDuT5mS2E3LQEMO0zzWAK2K+oH2jWR3RYqA9O
8mDMXWzw5X6J6oXHWAuDO3wnt5hwe49K3gguYg4/Weggxq4GQTHwC0LIUvq8g0EI
mmgyYR1JgSPrYdWL3hf+EZbEwszIvPgxzkoCDpWiSskl/3c2eD7YUlKr8Y++J++L
bNFo7wW4QaRkAReuyFCYKdaFjiLslFx5I+FlApAEA5fi7CARWn5J7X1xspq7jSMz
IrpkKa7++gOsXFZzFlW8rayZ1bj0/feSOWxX4wod3hw+2aLsZL66aY625XMjC6C+
7dXvTtTY33Eyk1tNxp/0ZdkZN5LoRZG348mPK2+WUVNSRVMujkEAX3KUbjcCADNz
BvqmXa8bySa2eLYmh7ht0wjVJCfW6WqiE5/nDKqcWUtIZEh/+Rf5VmwbhVlw9IA0
Ea0yn4PBWE5BjT3iaScybQ==
`protect END_PROTECTED
