`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rUGtcQNIqFl9e1Bd49u1VIAGZgRp/Pzv5lV1a1q3jeLpwnN7x5iEBMPTFhv66mZV
RKA0N97O6HKC8wB+nfMx2RvkI61yCUt0jNe7Xhdg2degYlKvtXB03ZY6tRSuAKM1
sMuHef/8qcXlU27cdywKJf0jwVHXUcfrHWrwvIvsipTMkzE6e+PUdXaX3u1AozTn
aaiJrWoIH5uw1i3XuAkE8Wjm2CMcQa++l/jWrliXwWpEYYA5bGJ1sAKoh0FJbGHY
N0etL/vlPoMxhGo32G9KnbNPFeEYV7j/R6odKzee8eimLFIufZ+uUeAzjDQNs+jH
qKPaHQovaory2TWfD/Ks6pkuGjAVoVpVgHW/tQ1tdHFK3oaKFnMpsTjhyOCF0T26
5qkbzbqXA8qthTHDGOA6YbA7nYbUJyl3OHNpfsRu6W5zjNetnhceXYZQXUc5jwTl
LfYqVNomPFaYmUDBaNx7on0Kk50pLiYIIGNw5UyL8I8=
`protect END_PROTECTED
