`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hrvjG+YW+IWeYwiZYCAhpUYeyBqzWEOrTdjyFmUv8P/W/D/ksJ06zVfjczJN96yq
eg5S8O+wrBDXIpoKSnabVK5qwVQL6QT0djNJh/8fAGh4IUIToTI0Ls15oCYrN0UQ
nfZ8jUOY6cwLdLOK9WjgoJWeQ229e42z8vhKevZOifHY01YOKnf/IiSJ5fwSBvKv
PutcAPj/mAmTK9KbeqMz+i1Hv8p4MPZb2uALQDBkd8hyQ3zviBLp5929Hpt0YqG3
N5jKKxwjbyj2UXo9Nil8I5ivVhxAu4Es6PW+fjT/5Vq3IcsEWWhbsbjjFcuwvE9p
1aq6+Ck60UNhg6dWmKLppXWQhFjS60kretGkbMWetMYomrmciE0WJP/8yR5bGlHm
PFY6qCha2T3p2X6qP5qlgwqBHTmoHhbSvOcQa2l60BM=
`protect END_PROTECTED
