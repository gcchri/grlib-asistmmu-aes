`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jn5vX6WahBKBhl59MktuL0huMflsWIkfoqbg4AcrEcDboUrNYmq9uPkaV+02iFwK
2S7CE7QVhP1aPUSVfDMIJCzfXRBiWVwMU1haIrXS1Dr5ejqhgilTGbX+G0xdrlaz
iK31Q7/OeAhAB+OgaeUdhV/WTM32KEoeeTVVL3gidjLHL/qJwnIl8Sxy+IqsLppj
JQiHfsPaC1XscYiS4Q30Vwqw5vYRSa8M9bgmwNhUifgF4pZ2e6V6UrSCvECpvHJq
Ct23qSiKs3EONvG8fZD1ickBz+9LJO8qJ6i1zhpvjfz9mctegyhzyjAuMbEPouDf
O+fq9tTQSNS1OpWGO6H2t9xuUK21QKf9O11ud5Xl/hpYxFYgScqiuPZSjxzOvG3v
PgRm+2nQrhd0xpd9CyDNxuf0nItecAg+54wosrretO8=
`protect END_PROTECTED
