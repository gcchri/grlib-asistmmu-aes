`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LD4PSIfjDEpJkJe/fg8MNTE5W2tIzQJsI96ne+RKlrMNzJp4HjyNjBML8qRxBZ1z
qhBYvJ2LAb9bs+Eb7d67gZ6OWSnrX117b6RpBQrBgh03aiwSUTtXOcnDTnImHNiC
Ob+I4YstQrHOqZRbElc95t2BqMv9+p7UEX3PJ5g6JeoI+THoJdUC7HlbKkRQSjoW
EVFtAIn02GZPTk85EzRax9d7y4VjUdO6yHNW3qOeGer9XoNutsuexdNlVxX/opuY
LnAg7Hzct+9MmKCBJlGqEqJ+T8RHTQV9v+qONJaYuV/WPPQHvaEogWJ0Ygchv156
LdVb7bwZyrnkPrWpe3Clo0XPirlOCADqrCG3HuQhekT7QSgUMndjjJnRn1mgYWuQ
/9UUovM+k+y9SKV2u6yVpUoCO1JogPa5latLGP7mZ+ir0AW/VfokJvOTLve0DgO8
VuCYiDVrKLCE4qDLt93DSGk/adHgTztvWCpgeB7bbyepqQ+z9QW5eQb03EvCduu1
`protect END_PROTECTED
