`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W02mu85YjQC2303ANfa4GHYyJMf7XzMcB5OlzP187fCtaANhler0cuJGFnsdUnof
AAJfEexEiZ7Z+l+9dxvYXKYOf5a8brtLGrZYkFOwc4OdxwMvNgAnFUm0XhJTazMz
+XH4qVKabdM1r+iK2KkT3hlIB+PCeCM24T+zcEEO4lA+r75ONOyQVSbQ9D3TdfdU
JO80YEw2nPK+o8C6fXHVf/Ep0KsJENLZt8WjMKSLt1XN4VefLkEjDYUf0b1d+mey
Gf4btssr1bST8UgxkTBvtW87nU8l3iF2tp+vSkZxU8VNNXrtyIpVlbEParosPmX9
V5rzfdKcjpZ/q8MOYoLNeIE+TUiMDypbn4dOF9O47+je5fNob65k2C+m6w+CD8xP
Ves5oE6wyJY1ZaV8CWqaW2wsptLl9aG7MpAfi9eguQ3KE4F26T+/y0j7Myx3/8/F
`protect END_PROTECTED
