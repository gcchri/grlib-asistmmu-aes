`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C8ee/9P92AdtAKqG9wCjtm+G/Ag8RjLCwaFRxgGIeFdBpzN7t3PeevYWtfR+36kP
l5CppGDRitIKORk1YXs8LnKlSWjKIooBQXnZKiFpDQUaN279ilHM14N+VfV/trkQ
zGNcd1+ZR+cNmgeMYIGR5jRddrEOi/0gu+O6MlH+JL7cFr1kf0Lfwngz6aC/aD/Z
7Al600lyhJGgprYlkKkIB5C809vOmWlsv5HBB0WQcthiKPg1y6x3lFNiTe4HA7r2
8w38kuWN1A6Hft0sFe+maLMYFdRspMPWLYi9KIi9eUdHE5HK+1mdHWHxCBhwonl1
qyhddK4dHyhU/otrXteoru9HGwgXVe9g/KukHNCpD1msQjxWW8ERBvmSr8wzeRuP
1zLrH7EuKTCo+RsyL0YRFN+5R+TywVFZQzUQWLRko2T7e2AJPRthKAgtQ85FTeFt
v0nuUFehcLQ2yVBW2Kf6P9i4D69xk05AMwo4X1sLFlomekBX0uTb4JPDR1x0+Bfk
qcEPaAQTEwUaerfOHZRTmRjop2W6ZoNJvQasP3aLSqkz5xtFWjwKMwkscOarg7Uc
9SLo/x5cQZOcYIcZz5hjhF+LCvRtoB3p7mFvAt6JLjYrs+P42eNQauCrU+zMbYOA
1zujJ+XaiUDE+GhRLJa1Rpj9Ya4lqmnJRu7xXiHZ1rXFMiLVBE1jlcy2DErjActJ
4nUITzIxKYP2dob5DH+txg4jW2CQszMGPDMnQt89ezJM90/rZ4jQBLc7b9mD0k8q
`protect END_PROTECTED
