`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QMWW7DOgvQp54pBfQkt54DX++ld3FR6KGusuA06NhaxENJpw9C6UfCb789XK97Qx
524KmgiITvUXTGL2jKl/w6hKaISRZM15fN/uOUspDEVkRkh7x8ejh9Xp6iV6zAp8
mY/6sNwnMBDu/Tpqfh5ZhNEXnBV+iHv84ubkwhJwwtsig0tXROTXXAnfnIz8MpQq
kUyIWgDh95MfRiH8wLEaWFZpjV4/eVYmjbKhbeA+g7lrJl2NDyAj13/vHiIcmqee
kWW/05Z1shdkaJ8ud9swrdBjcaz32nsQQ9AtPI6balIv5N7HUHjJ0Z2FvbjD4uk/
A6NGGh6Eh0eRwChQF5d8RcEb6DRxkpQ5+OFyysThLakavkKGQidfa/F1C2HolQVo
uFX34a/KhyjEnLUjWYKApg0q200A0sBJWZNcNpOkb/j4Xq3WZTdQ6Yf6wtdEU1Ey
+i9Rf3ypYaL2w4l+GLUuyXV3ckhCygvl+PFBXueelHy16IRQm3gMYK0t69LJqwQU
wtZOThnNIdXReP18SEmcFDP+UQT8ukxUCgZ5LNzixEmIK95skqmogSezrPcIJMqW
VopNdmlrHq7hlKd0DtKcDCYN2UF65RNiKoLANvyemKv04HgSTsjCvKW5EEupfQsD
ipZe1OyialGSExf0ltzHQazP36yog4vUyzoEb4aopkMg/9l0+FlhkAwjUbxwl2uE
lOWy/wf0Mg678+COcxqXjRxyxynFtTQsWBFFnGNoTury7hkWawQV3Sa3JRIdOtAF
8AvYSy00OQLomtt3PeISRQ==
`protect END_PROTECTED
