`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oi5s2qy3n8htbvcEviap9gpyxH3zEvPLWLNguySl/jZEBqJv+aNJjocPdu9Njii4
AVjm5rnGDUTdWF3kgzUrwcGSnbWG7z41nTHAz20J/+W4+kSyNOgmJSAdhPkEcy8Q
lcDGX3KhpyxQuSLEC6M4hKyPsNvtfYNOuQ0YNaKug1/sl0wGUk79OEaIblfiZM4s
MPaVW+xEGYleXEgt95ctbMLtxF448TvmlgnHDQHyF4IwxJ2gXuMRPCsjAkJp80HI
WYrRZzZjOmMzF8F91pa19w==
`protect END_PROTECTED
