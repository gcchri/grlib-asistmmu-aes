`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IQ/UQYzJ5erag5IDzvBwYrEUktRfsElvfUJxFPnMHrUXCiONXXEsLeWcdglNWNxK
XXK4/B/lNqtn7Mzoua6B7mpJS21rPwBgSMcNEX/qdJx/XBf4eQY1Fy59a1h5n/K1
be01ckgwXSdxgH1sDCQSNPCPZdA4WtAcERSp147sTOY+RJJcPLDgVt/9Ruhc7Qnp
QHT5TKlxwGUs40u/54XfGBkyqS8Lkhm5l9MeZgc7RzhNO3xADzIyzQjLgwfPhgN6
nkmsDW/I0ASs+utcZQozCUANKzxXtbbkfUeaCoxFWyqJt7H6WE+4pM1piKwa/62r
ScGPC79Du4pMNq4YXG60OIo3WWLcbvuf6lW5B4vDvn6xQwIa4i9aDtInSR3odOe1
HqER7UGtMGP8lPm2PbrMb8JwKPD3b7VZFWvBwniqjVgjiRF4Jj7bAqeRv8QYuI6H
V4uapfa2HvEQKn59+LaCLxXQEx3BZv7pyyA5PlfF6nQ=
`protect END_PROTECTED
