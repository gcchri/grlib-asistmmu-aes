`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OsbwYR4tCN2vgHWaculh8Gr3dodrIweGeld+TrBxVC6QcT8vsF/EcQLS1yOVPsAo
pa3zbFaS7AB7gQzsBEjv30AWp/BZn7AdAku1G6zlkU9oJZL8LuApvBEVByORL100
wMVekZEZl3Uo0YHrDDTI6iuxOfmM3fCyJIzUR/Y7Ptf0MsrHN8KtSPP91gYZnkX4
fYjx6KZZnBy7iVjlPHbYlxpwyIGImFQqdtMd4GfuWzT0ukIaZ3ZtjdNcMdbguvb0
QQdxKphL17SbcEU69EpMdAbpZ1Wq2yOjrYxsqmGo71/VhTV3SLqxkvKFKi5XScH3
0stQLeO+H8fV0ZV2S2VkM/GXujtshkJjiCAEfoStOLzDmDbd9/XcEYGqEt9eIma8
Y56bcKfJcPFcFfW6ELO+YYLuiFsMA7RHPCZmma4CtILDMm5luYpzNLBy66UbImFX
wqvUUXCViEe5Vd9YThcyiikhxqhnrmC9V+FLPVpFhml0YW3zV0f6EQznoL52Kann
W6wiqntDwFbTwlicEYx6eRtm+JaTWQVEAFF062XEos47/uBSQWoK6LNH8nMPrewt
Ftuep+MxVADERqVTQU5fal2bj9BN1dVe2ghpQfqTmUVWJ/MmpZn/ksTMVu871kX/
zZWgTOosRVi32V9YXOvFcf2CWvYfGKa8f9yJ7nxMNhANYGepA4EXpKcyY3yTVi3a
AQeOGI+90zNzm0O1WiF3Gc78Ps+gGa5RN3FRw24TMOb8sJCAt+wSf/EBcodzBdtc
Kd0XE4NmytsCVOLMl44LQS4fNyALJgdQ2aZnRw8qpzgFAXL6yTHK2VPcoQ3aeATz
TO1F+dNmVnHVZIVX/HoAonlK2KQPoP7njNctkYGCQXcre5Vc5n80H0p6hEBc+I2O
RVwXjFzEUcsnnnS0xt6IKEN1REPpHZwpUwvDj1MGeMu2WJ1o39onWxwkx/jVHODK
BMIZs2hujIVIe8LlvI7kNAGoNi3khaaqbfMoVIvLu5Zs+cRyWX6RaElM89ptE8Xy
ZU3j85lK65/7TWm3TsXRmgzPgq7Vbl1apU2pNFDgiQbOWVIpQzQQMBvfMUP1pfWG
snPmdbIqhdRlxATOLQkB0CPmjBI+FFoSHla+cfZc1j/26fXZHsXxoeZXi8VNOTzR
i+oWnq4+dQqAhI819dAn/7oQNGrERLTF1rP43o4jUno1xade4rIC+2VZ1/yUhXc0
jEXKxghb0GtWPlenILCmZSlEQdLaZ1MJFNrRl0zwYq9Tf9cXesn9brKcEuIIJaO6
xeB/yMwNZSEp5G5AJuZbS9Kl1IHhhyAd6/n6j4Bvo/wKMz/5qIFz+rrtkTS4wiCS
KjmVHTQIlD53MUckUpoQSoKuBtFaHQ/pJDUoaBQKY1/a28XRsatLYGIIEKJYi/cy
sm3UMin2NlGA71zDhz+sLKtory7PTYyDA5wld68maJ2zI8gi51v/O7/QynTHoT4o
MidLtXwalQ0h59xRLGjaXW0gl0xD//5I+n4l5tRrL2wID0Kj1aIAusm3EN/dEVmY
6XqNFc9xWOkzerPk8rmUGvxzJQJTHJyd9XLsK6KHrVteDE6bwbEqNG2cuPuCCbMr
RYF1/7aO0yxzOHTdz38ZHXPL9LKJxL24cMxoQe+ggDudPCso3MtVA6h9yBxiDSGI
j45gqIsdHK6SGhu/yPAGYa3cI3CNpkCtztB9br1bQQUSBtofnPvXrvBjU+z6e7lb
7bYCHR4da7l3vL7O54vGbHxI7xUZLnTENc0PAuTWG8jLuGJ1lNuVKxVu4RTognIq
dd3Tv1EC8CHoj4k6xIvbbUShHyYbfcvIooz82OCzF4B8w89F7kyxOxjDVPIXbelP
jf5a3qMLCd0tMPG/wOPXL4c9zWGKjylt9yM/WyROcl6rl1jd4VUAgW87Z077YBq5
YZdepGRgOPupb/hwwN03FDX8EJ0+5sgjhAuc9ivZDdhp9XJRgx66am+tRgAEg8L+
LEr65xNS9RE+nIqi2grqqDGQRD6Dn66D40ppKH8Gawty+hN3pBiH7wR8uv+mVQoW
qYJL4REyhl5VKaSwlU4pJWzoPRulShZx1O6L+EL0la+tiAwuALhUA412pjv1g5ZO
PwNnENsDp0M+qghdu0Trb/dwf6YajnwRTt1Z2b5T8p1sJ7hm6aF3lrVV+Mdh0UTj
fwnYQ3nqarG+V1xKCtD9642OTSaHO0P5fePa9UzbRMCU3gK5MhEHbHrJfooLNjit
Cb8JBXjHapiXFMabJTcJPDLbQ5QXX9nPHzrs3gFty/PEuag+6rAGRhwQqz+6jtjc
LyUFdG0BinEiWel35TF1Xpe7gaKZ/XgHXGtB8xOs34WMDiDLejFRRm9EjGDUaXo2
RAFK9ONlx2kJqyFnYg3bYE6xFOkxdEctrJJXXdjGbq0esrX0GLZuJ1EFpgV9gc8d
5LkyAQMhTejEi7o2RQCejX8Tyk8dkrzHMUPyprlOVPEeFSDz9gWDzB+4onVd6Stj
7YDIWCK6IXp3NmF7aGHyjix6OfTP82G7sbKkqI5l50FuHFIQh30RUDyBv046mosq
yXRqS+0EMM9b9zS5Kizma9p7EWlc82uzNYBZP6sUyFszS3ZB8NRQg5sL20y5TujU
ws4j05Tz2aI1AMvtmu/F2niBggx+QHaMxeJIzLV8/yu8IfZ8DU7HxZ1TdldWeot1
CV2WiU7yjHv10ilnJulI5tHevCa4vpT/rM7ZyXBxcRNiJxDolMLIQh7Z0OFN9N0b
BTv3TO/8nNqgi1Zl5B1sHajWP9ne1RVtbqylObKBmQPQC/G9r7oV4qny25T566d9
abIiYnvYCpRH5OdHvRSC7GmQOXF9K6i76pih9BNPqLpq4xv5cmGFdxbam040aLT0
H+NxzNBezm897T5kytpL5ofproJBmXCuik4aUSJquCRk2w63BRL2v30Pz4ZCuwJh
+QMvZWGp/F3UZQvzSW9I1FZKOU1kH5asJNXIDmurpYlDju92UnyO69l6cIbjI2Am
fHKFl4yhNO4eOPgQP+oxS8ZgM6GFIqRtnnP9IPjax5xn9QGuna0YPY/n3vMDLpGB
d34WTZr6BV5nsKkaEdWl0jah48lbVeWQFQUSU8fqgjUeqZMiKWTdC0FdAkA14ld5
3A4/SdEvc1KJcXFpuGxCTELzrz0rcKDjaCCUjjiLlY7ZJ9GVQQX4qxjbgn4YtLxY
jMB20Q/XWmg+gH6AkZkShItlfZEAJ8pu8x0Uua41gV5ANzf3mZ9J2miJEZrj0ncs
46XMVnJeqfkDZZWVPfxWyUpKR8U0mWgswL5b+RGncFFzNR0irHOnEKXb/9+30w7n
l6wrUfArykYbs+w4GvkuQhj5ytCyC7JrrefNQ0TLmR91O9EnqRXSQVnx2H4ioxLu
eqqFeN9tAcyb4Yah82E05+vH7cmppkm5o2Y6KxgepOcbG1Z0E8M+XKzyba/UvudM
s+fswS/p8HkEr+eM/dHq9a0MymNNmfkwLRZ0qeUNNGfqG/jY9FJjg8rcx3AuCIyw
bLKxmoVzm5AYui9orDdvrg==
`protect END_PROTECTED
