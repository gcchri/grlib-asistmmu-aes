`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sb43Q8mq5REwC2LEsfB7wTku/29ZxqllmllKW/VPMLknB0A1nyLxj3LD/59RSYto
fRV571H/m9ewq0abSXKwvj7J5f+Ki/NaVZT0Y9UTguXggjWZupRtCfQaYRBpUibm
P8HdWHUO7OAJszlb4solNNWC/7kDz5OcIbYzA0plV7uli/fL6AIg4vB7xvfnbOs7
U4zFs7nQ0Fuw/h106GFIoI2VfFs5ROvAVeQEtdSDGC86+C5QvUqoOVNNcbhOTq0a
KTPCs4g/0XdiHovi9hwhj9pPS9issd9l+QLxk18hzZ5ESPS3uEw7NA/1RwcPO+WO
kSQjYGFa8EQAdC47yvQWbimXhSNwPo9z7suidOEJgw6bUGuB/QgUu/S3Bnm2ppjA
2gMAJGy8lkHHf25VSHLimKYg7wTrriqg5hZZGsLNe6EzX1cK9uIXTPpwZm8vlhGZ
swaC7ITVAVLZ49f4hI7ViQV8ioZoLktOxVpvW+C0jTPsuxgF8JF5bclHA30mzGBc
xGeOnSvsmUbASC+lAoDhag==
`protect END_PROTECTED
