`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6IjAKLXYpMJShq3ngHgyIkZosUiTmuM/GPu3DoRy6vrifp6kbdwGER+stDcQ7Cx3
1qw4rKxXu12pRiZxkNLu6bDudOcfya7miA+D3TGnuaWwgHTnrV6HFT++3GsecPGN
k+HdEWa/3Ia7d1a24d2qqM2YEiJ4qrgK146rVSmCYXTd02D4qT2NIuRP3LreI+ur
0Nmif5zlfrHFRp/RjmZuAToAHQCVPylb0kkfrjMjeG8a764o2kcQu0clOyTGRoIj
+h054CWIgmTP3qMTBT8XhQu7I81z5oCOU5YKJYQOeKRYi9t9dQ50v8eywfb2xRo0
AqUQiHiW5UjdJI+O/e+BbpuwFRPSjwttr8kxBaXhGpgBgqq/8Z6rpguuWjd8ZVB4
Uxx0VWR3C84C1HeUyNpQEcVSeXwHL+mEbX+klbjRPp4+6uLsNKHmIRf14O442fbV
tJnLtVSO4ZsrBWf8/+dR8D2hP3d140m/G+g8nE8fENHREXe75o99UOELUNVi5L1H
7QYGRzo0hZ04rbx4Vq1SVyOoDm1KJULyniSB28eVVi81GRjxnZbreYqBH+6HSmrM
5QoXnsc9qhhH0NN87trXNA==
`protect END_PROTECTED
