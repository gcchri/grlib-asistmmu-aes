`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kbd/FlOKcxAqO5L85I1zxT84/wQPT3oHul62m9OH1Gg+Y6p0YOKFLaMaoxmhAh8w
IRJVVX5vBKWE/tZ5QyKZDmaxznynww5zul6k/YK/WwAUn8ubFbPzls/ofY2ROigy
uIASjxoFArwZYy9Lj9hKrzi+/OuugYm+Oe6wZWTl/bqoL1dCANT3gskwrBOQig30
l8wKVtFPkP2LAx7HsVtGHBFyPEgUWeIaliok2dOk8rWZ0jEgXkPFcu1RCrZCtKhm
ymQoGAAmMJBQpBSryhcMsbJuImBxmZL1S74Y2k8V4hAX8QbRXP27MifKn8uMKD7h
0Bb5iid/w1/Vad2ITlsSYr0QyY6bFAQGnTzNzK8XyfoXgiDYbCatKt5evJtANcaA
mkcZ0vwExZzVXU6+SsUvpmIT1jjqy4Uvcx7/zU58rBbSSsoiM9k0Qpj/5SnfgEGR
kb/qPfxZFCMTm+qd5F1uXc++NJTAERGauJeh3/93AcTsWTRl/tuP6ohEahPb5iqU
P+MerlsefNVydicRWf2MYch7MzcKla1mbdC56sk9QL+tOfLFHTE/EzNxrAjVBIgQ
DAETz7fac1JM+PP/4nKVa8CUbx6FQB7yTa/uRJRVC26pTc/SUHu3epHrmBDH1C0F
N0MxUdR/NAhkVSnaRnsjBHV6NTgt4N+q3aVmWe3Saqe/t84QIIc9jEgVTYeOOB16
Z0V6BFYUQ1kw5KEXVVH3+X53B0SPRQvzi2gZmXF1ygF8uyGchrfcW5YJ9LaJegn1
5r/lq1eejPYwdeY+6R0mBPNYgNaq7BmcujKG6NUBlKxtLNCsQYQU5wc2Y9XojE7C
CpHIbUgP17u9ZtdoImX9v1MqM1wYJoATWu6YPMIwP6ZYzYvVpDRCHqENL7BHbRgk
NJDTs5A3UuY7Py33j1etW9mTWluRYI3vr4jjgV1/6ae1ZNK12IasWnLEayXEmFaJ
yoPiTZGZ2JsDJGd+0TD+6xYkNDVRy2lgfc7tHb+JKLyrpiTN9NwiyDqLPwrHqgAg
wz3O9Xp7CA5KnNilBBBfg/NY3k6SS+y6/PQ9BUhf9CCnBEG37ZQTHvoZ2qHVV0+j
ebABiAYGocfV8tiWfXQNlp1DLKG5ZBbiEp6UvLO7vQnJ4vbE5IEQC+ojAlnCOWpo
qGQdbK0hltqa5ORqt0Qcw0n+MaVj63vmV04ReBreSaRhqXMuzJ0wnMgej9ueBoq0
FAe31EwzrY7mSQBUIyW5tu8qiNQ5VjVg74TO67rrIyLt0TMlXLqHEKNrs1XDTaim
XlReQmktm06VZx7CBJAoUegSe30jCy7er/ujSHKUOruta0lM8jJawfmX0/zefCYr
sqbSW8l+Q+mHNQ0UuTf+RzK91PbmO2XxdXrlnmClfBcL6pmTLOdnI8wdb5LRBFns
+aF979UvDeQ0waRF+SPiEv3vOs854WrPFzfHNovCTCkFYPHLihJOOf2G0xuBLhPw
ETQJLrdJSp36agLBUnfv/vq5QBwUU76k8kyC9mq/GMYr1sSSuJ63nGaTYxabOMbG
ER8hBeXU/p6tfZVVduhJ8bMtIxqHr+AcEp4zbbVO8TbMNRQJBV2j7JNHI2NYOaRs
y0LticmFDydl32OFmn+8Bk47GTByU+QVZ1R3Xf+Tb/euWyl0dUJkQd/67PLXRV4Z
S2NP/Hxxy0XIGMPRCEmRT9pmRqdWX1F3ep+4A39paUr2UzLYvUDZz/6W8QhvBh/K
CJ1c6ht/9oSh1HFfUcC+HJ1TkAV4Q38VT2R49Dw96unTL3/IA00O+jrGIH6EoHWq
6Ib/dJ8F7a/n11gUBHbJVJ27enCDWF0Abe56HvlP9p7iT4LQk3pLrY/jsiIzWZAW
dvMoH5HBxfGhe7wBGZLDX72bC2VFAgg/1U9gD/CVTvCDJv5gFZAFYnSJaVYhv5i6
9aU6ADOWF/5Ny5Ad6FONAc1QNtG/dhndbptf9mU4WRcoTUHvuzNp5HRmBjvmDT3l
`protect END_PROTECTED
