`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jpP8wmTLMlzJuhc1FZMTNfDa6g+HmUEAMRS0ZEgoa3vdBaKt7HqlXnGB29bjrvL0
eQmJtIwhL8d/Q83V3Pr5+aa1DSRHt9ttyAN8H19UFgl23suyKBz16UJpTNBAONMo
W5z8ZLKjBfCYGQSwJLMKfCvvpUOCjUYvyaoKrymGVkSj+4sRWHOnLlkbk06sEyLU
g2BmW+lgvnGQ2j8Sr4bYJAaJ+4AR+npKhWJW/+9MfyqBU/sg5jyOOU6+K2Lynt1a
gfWnI4aQefAZigpzFvHg3PTmZA9rtBEJTF7aURWxpfSZWtByOEOnZi+2xFwE/fjd
l44l20f65SzFxzOuAuYxgxDADmwz7TeHDQu/ywjo8SSyxOPh/PcTRx3ypVFv7u3b
ww7rbpF1obIVLr2niMsPoShGkI4SGMp2q7GWemGpidroAkOtzq7AGyqSJf4KRsf9
`protect END_PROTECTED
