`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4ZhQR63xsCRAfiBeOXApsRIwuJTEaiivXJO3UkWaLfPy1h8/4+Ra/oGMXemX7Mwa
okc/RLI5mRKnsDXMb1D2abQziQFikUI5AS3USieyNfLL0UPJMYJY3mBoceHEGNeV
M/StdeiECWS7dEwE3RxePFa9PE3A5M2x9dfQxMwATrqWs01q9OwOy1d+2gXWmOfQ
1M4PLTVJK7o9IbAbH8cS/Pp9VuegXCiVPrG/xi0Vn3jQkxv+W3YK/agxsSxNZphL
e71kH3sfm1zf66awRZfklGqb8SGIqO257qHSXGrh5FCDarYF9ng3vKwMA9ZHGNPG
ifxb0ykrs6wtxGVID5B7tAJQc6b31esLjnSy657tblZcPTeamtzx4scv5vVAu9Nl
NU78RC1Pg25XH0rBVmViOloQ2cpRy8zppszHByYKh/ao26hTTl66fpKjLDhC2RQY
29DtD7VNF042I/TMaPbRVrn0BkCH1NDbNJIdhqPAAgnewMAFHjH0cgebQCXHV1D/
TKKvts5a0ASNaJ19nhmUSdiRXSicHstAlA5YXXCZwTCHj28C9Fa9LHgAwPce2y6w
VkIJZkMeb8NCWsF2Gp2VF4qrRfIdz3/6fAU5B1aUm47Dn9Eqroolz3mBTgZfKoVg
mlC/0C/l9mMKF+wJrXbMUhG+o8z6KbRM4LzuKuVh7Gvv4CALOMQ12zmLHCnWCHY7
ssoTM1A3Xr4qQM9s4l1dx7498fIZF5WQ3VNmnsDYl7W4cNr+eQStQend4oniPkvj
sLurOvypoYkKkGW+DlUTtyemsrovk56H1EZyuiDiPm+GNNHHe2i0LM/2y1K0pgqt
avrif4WL7El6SPWlzB33CrTKvrRLM+HEiAdgYZHDjwLOkFn+cY3oDYggQ/7qy2Hc
`protect END_PROTECTED
