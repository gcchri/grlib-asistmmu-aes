`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GOgui2RYyXz8tZW2Q3oBxwW3LOjZ6QkDUhErd/YQASyT7nPYb48HZxfe9CKsdJyw
Klz0aQVl3UTw1n+ja4RVjCSQqojEq7W/FxrSP7natH5jg2qaagv+YidgEkOxZY9A
DHW0y83GoLuysIYclgQh6IakhlLY6QL9sG8HuXbBkqmTS1OhbkEZIsI2uIN3duHu
MspVQiE+we8JUIuE7tscR1Ktioo7nIhYlvWTtdgIlKHh2jZStSbKPBOk/w9zAIhD
TQJPWO/XRWqgaYBCOszgfhPNcYoX/8JNDxaHhKnNzKbPiG5/4SPMunQmKhYVyeRs
9MXNWzky2QsyjhFK7raLj8mEdaLYRljr6djEfymd0y/ehuqNeiI6mYiLRdjGblx6
w5NOj2zBxmxqoquAgk1LgD90J7zEIxPiNDjKFfa+2XBuU12y4D1sdQ/1PEmruCBl
n6e8XfKYb+S0dh2uunFhQZGudt30iqHsstxaEU86sQIPCrLZgt3XO60xFSu0GXNx
v/LjGls8yzskaJDMVkkwo4rmB6cNLUvgat2HRlLbnLRsIHcdHBd2gmyDpLbgbhZG
eXlp0U04QrqmoV2J+nRqjPgq8qnnBYC35SM108TbhHmGzIDoDrfAK7GFiD0YG4g9
m4gmUraZ2I9hAHtf7vd6W1RgSN7jJSqW6o4nby6l4bBUnRJMnRi4x4jggbUOgWFt
NS/IW0bYoUWv5s6xVmyUgx3IF3AUO5eH524NAylmccR+Dqow439F1/vBkcvJ2N2P
XpzdVwsMubtWuhooOaMNAKyGxtKBl2cURGNJpsnBaCSyjNIzxRJtfTVHv8e4z079
8NaEHSnG0bs6/UGcvVsj8D5Gu3lFmCFG/9TypzNQfhh0B2Q3xDSzHPrBVyWYN1ud
aZB1pV06M/54Beibq324R4APJCb2eujyhiSnyY6OoIQ3mpMFo+f1AyOLrJL+82C4
bjVq35VgkWraBuPFWpyJes+nd/vBYQY6Ob0Gb3eHdpXGg7Ig7GgQY1LGUJ8tp0AU
nlT79Sl7DMii+78SauyKq+lhJsrERkIzvh3WkkezaEUeXhjByyeoVdtDQNcr22Nu
RdHJAeXP26UIoAFZLy1NRUTq+wjNbdcWpZkWt2PQO11TY4CFtxKmX8U+gDnagggE
qgRDYnYJHiuDlPTHUfYvzMLRsBJBw21EArFV0lfJjoRNSR1XsmizilQJgyfzItUg
jIN5NRFRb2IsXrauzk7cuiP5dWtIBhhbu3peS1STj8kDPtEhC+2gueU6tmuTOEGk
hb4q7OO6MDyS2CB8SAUvOxrZjdMe64EcA8tgTnsyd4jRekYBqivMC7YNRFrkMoWA
V7CLG4Z7kW9Z5ZUqtIxNP8zggArodcdEaZNXtv807vSsdyqh8lshX1UkiOWm2ULl
aYwjxw2WTBooHnm7bOpVPF8tdJVx5C5YJvbF3fb1zGqORfiXLhTG2ohcRjINRke4
B8cksGSsKSe//3IhZUMUVrRV/46mHs3D3xSvDzmuOTTFInK01ljIcZOyM52ZkBqr
SK8xA5OeI1xH2KH8xH1s4pjcRQsgvinz2syHBCgp1C4yErFMWab3c9137tjgJL5r
V2FqMTdw17IoeQ5izPifTxz8AcmLs/7F9KoPefKlwgF+lKcg4bgJXA9KWwsoEQ2y
q8nOCgof9lB3AWBEwZiN3O1oCYPgRxmGUPb2s1TFC6oLUlWQQIQYXrHTnK6sAv2j
UmKDqp4dXEACP5uOnZi7qw5miDDd9s7QJALvgoz61Xb0AEDoHSlzGe/Lt0Wu9Ws9
gBhQya/jzDmtRm03QP7mHxqmqiOkGAL+wLARW+QaVKp+b5+E/qSyei4VptPdxxZi
1gOy4YYwGaAaifFeOeHugKlq8bN6fqi/EjywS+PZwbHuseNoNws0eSI/rzhkV7ED
9BRWELvSmgraSmjXV2or/9J2HkntZ8lJUYaaMp1icC+h9C4lWCkUG6nkBhTIDG41
fn9KaGgUvw06qk+sKbQ15OLAa5M9hU3yErMOHi8NdUJlsD9SdhGU8msPVB6axNLh
CwB/GhLRjaRDo4F5qB9SYjcE28NFLhJKWHaLB5gRyyfxg5tKAl47eDVM+x/w4ZAE
69ctqPjBIyqgAipLWsTzqXh7SncU3qC0TFmul2uuDKsmW+eAL4f/lQDGoG+CbpmW
CmpQFBXwhPpf14HprUxGb3zj0VR35crhEUxurOi0ucSF5oKtUp19FVoSdoOsntzr
L1uxEC+tquqil704mnBjNk7afZ5SXHkyaHz1651JKcUPwrs9FxzRa6ec5EDd6XTS
Wxgbd2P1wb2MVg27F7L2p5bacff1OJb/ExQIydmHvUQ0sh4U4WXoCrLi78GtRZeH
qk3lQLWXL9HCHoJ7YSlYezldDJJeND9Xe/cObMWMtptD1y2yaxTPCCvJfPbI0ygk
kwx3uK2PGF46Lr7jukSyqJKynKPSk5DvqpYwQ/+kv5rgZHRgrMUtOJhi72A7kAwQ
PXRKN19ek1zQCnMEXwLq3C9ycd6h9G3UMm2G3aoaxVRNqWP7uN5JtQJT4u0cAmtK
KaBzU7jd1IzkGMPhYXYUqpV54mvxehl0eVAON+3Q01yBMqgYTF5zfvLYFvgIABmm
6EqHVDBLBWWz4WuvmOSuBY/MESNP/VeY/qM91NoB2NpX9wYY4xWbBiYh618YGOsG
6KUX1YP9nivpth48kEZ5fIH+gH1ObETFeDJPnXqBZuxPk4GXV39jDSlx8wFVLlYV
PHOTQEjFmUX0BdS4oORKU3RlifDxwyBP+zLTQT1Xl4vKA9xF8lGclIfEYOs0KUwS
mqtYrsJxtbA9IXphb9RGafdIjq734B3CBn/RxyL3T+OXatOqTdsGEFv4p5P8ulU6
xtv+aHxfML+NKZ9w6wj3gwW24LzoDC4IlpoGzQLppySbPfXfZxyhev9YoRWpuQG5
L4ml1XH6yllKog0FQHjwuvmRfZYWo91IoyXpZnKpiEAYGe59zNqoVWi1YCZAJyN8
B/FYy2jSTlGxYQsI5ThYdaARkNOXj+ugk6ZMe9K8Rbi0P2O7cuS5XQXzmrmwgzsV
1nG94FvsqJO4rCYo2phNi+2UQeEVsEEwS9BvLDuVv4hfKqrm7VbqQIzCPE2FlYbA
OiBshPMnH0TuU6ao5wpwCJ1ihGyWrewb/Ng9CFGBuDM3yha+UHLPDrCTh3h2L8M4
1VYUURByGqeDGw52BR8Zg31vnbR9d7bnQH8linXlk8LxljySpJrCz1nHnNtZ45sR
R0MiDoTPvba8YfpFDN7HW72zAfaQW82USFNYPzVLR0jpcGCpxgT18gtdDAx7pQs3
IXAqHBE5RdjMQqNI6CvEjG5cpV3wlRpBjbWGDTxJj0+IChKZiCLoIQoiHR9JzSzF
C3YeiXGyQF7Q5NonyrypLv9r3dlH6BjpZ/yk3oF5sZYnd3BH0b9D0FbO8G8vnqE6
6rPnX0i7Rv0RWOlwQB6wKD6TzioyQ5r4IAB2KH/EkrT5K9LZPv/Jo8+JUJqlFwKM
ItLTZ/RolAo9DwYsyJuWQAuQ2EUgJQGsYZlktPS0QWnCG6mwF9RR6Oa/EcWScymo
QogI7FhQ2iOCPypEL0vmUQq15IbgElnuDDSTXCYn9rTW9Gmpf0xDymipGxUmT0yt
Kk+m8Gc0sFnCQTA2tTg+G6NctuykGEdOSZK+so9qEGsurUYgLCfLrEKq+V9Zbug8
WIvcMh/zsskBwSfK5fTmZ+Wb2Pg+BrjbgIjGXhwN38lKA3sIPeahSzJryQXZDViI
frrmKnTkVKMEzm0/E02sgD+N+4jxTZRO8S3sNTfvDpxbe7BTPsdLYB+gVfmQs5Jf
9gKac5frJiCY5zP4lcWeuW1Dv4TTl2ZK63EOKkrlooX7fNYbMUZ6lAtflPxoEkCe
R0FYBLqDNHS+xqhtkC2vDE8lU0jDLynGPrr60j1DBTvNmx2iBF1wVzVyQXsLYIPM
bJUMlMpN/KpedlphfXSU3EwArUbvnW3DK0nmsPx66BFIB+hXXDz9ft8XF2as844k
nIuYKdflCqsAqIguDl2VNyA1QQdFQc11AFmexE5FUdEwhy2Bzdd3hD36tF8UuEEf
8AbT/P2M0x1qQNXbIgbEpvn/KSvEcioDQoaZmNB2KDjFNZyZSlnN/wOuCP3SJdW7
5F/6DlQH1g170a+2S50YWfUfX0TOCLcPYBAiet0OCXChsnhuLWOvCRsrd/iV+gwF
OexTD38v5iYDKkBiZdXV/LkyW7NJKp24v0SNjwNU8VaCz/cMDBF/oVHVJaG94X3M
+cLUHMVol9X7sMbpmCZ3iNqFb3/8y1FHcPg5cH8nG1WSWCZNwkPV7dl5fG8dxo4G
uIH3pmKRW93NX+HZK+wo+0wJEFIgYAfR9i0KOsTWLHaOvoaafnLcXp2pH2ur9AUI
4scjfCtQh1uoIxXvUQO78lcNwD4FtEN24rzc5/oyBMJ37rbtc0kxFlPgtKeFYRRF
ZAB/oigmp5QAHuySj3K3YT7+hWnY/JXmxlRqumEb/vmrvpq9uHAm0T72N3i2ZcDD
cGcec1Wuo6LtPA+IOspv1JR0yP71q3v8q6mGSOkby/To1Ap+N6WpLcrUJERr/yjt
GGbzSfSUcuQ2waNXKi5Sy2OhWf+qsJWzurYH7MDmBMhQQAqEHM1tjdGJPCZdOGMw
esDQ9vBtGOCQZNKqqwR74fj30dsQwOPBI4BklK/GwX8aG0w4ZuKFpCwFbaD1k0ru
mL0IavEwbjiTbnue9G+BbiHTq81PKd8yNhrMtdGY3zerCpKAiQeUc3v2OVwZ1Lmy
Zg0VRsMHcYW4Y8lmsf0j4t/iz4HCKII59t+KwMz84slRzU33rGntzzYm4/MfXfDY
6DzECxhZS9tiiDmViqXPAsO0KTZ16+4xQO/a70nciAB+R62jmeXMpr7SpRG89uuz
oQtB9Feh6d3M+3s9ULKPXM9HUSaf6UywS/T00hnNaoucFtLYWsKoXkWBf3mGrv+2
UlWL1Y6a4vXYhfP5VG9lgtwiJPHviFO27ADfhE7Ui/e16dX6gO5AC7Zo9Ckj68GG
3/teTta4AcnLLVPmfDVGw7IE4Q2z7ObpkJxtQHiJdZZr+P0qRD93E8hfHz2zrJEL
9nBDCS86JqPgaq+3GOx9K34ZD05p+P+gBK5RuxKJ9fbeRP1auEd+apbEsZ8Kvx11
28gAjMkBUireHAaa2eEka4FsACP39MQfFbHFamp6zCCd22VIyiTbuUN+i2x3xGs7
S1zTO13ooCdY978z2ONNIlBsEssmk7a0wanHUNbyagI+Ay4+BHzQyISbQ0Zg7bcc
vBIUwfzas2Wd4OdFByssJXAoHMbA6jpljkuQ/AMVwU7NdIakNo/AqufOE0w2Ewhc
MWTmIa4ytK/e6MX0Vj703UKr5a71MAaCRLN9CiMjYaAFoDpei38LxflyfmKGi1JA
WShmY5SH+3HdChrUqByCHUITQgAW2cnl/p92yNRpuue0iRabZE1+hJQeR8Q3lcUG
NU+Guh9/W4tR3NeLXBHssi3r8ky/O1aZzCG1UeAIC50=
`protect END_PROTECTED
