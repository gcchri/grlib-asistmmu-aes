`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5y1qWVyhJpdGZVwR1naQYBtNPtmfD8JGUL1D05q/e8FJFRmdXFNNF8ksY90tYP1y
uDExAVpc7fSDiOmmB19AJ8NDiBtvmg7nERz6NSvGvTQof1JDDHTe24YWU8RogTRJ
WsJVCF6GW50MkjJWsKy3c4zGJ/eR4WJ4GhfFflLOExTbm4yn/eS2fvoIY0ZkOkMl
lS7FiqNGm2yOwqHbf6IFWCEvxxmO35pBVJNFuIVfvANbGtPLu6ensncMlgK/5fkh
JydKk5eEnd2OGRRq0UuEo9I51LipV7cdLqd1kIh7qBTqHM38J+nOSqwf4LPbj7Lh
iVaW/t7BgUeqG1VTYsUSub7yMcz3qvysvKnFOonAuv5QGjw+vZBIdVhbEIF96loQ
exgSfjZYuVXk67BrckYyb4frb2o/xNL3hVLTr7Smj0g=
`protect END_PROTECTED
