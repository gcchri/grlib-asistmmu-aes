`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qPEZ/IspSkjUGNjhXgYoPT8me4QUYo6Of6H0HNNtcDmyNsRc0Mxj2VTbhmQgHofn
cBKijn4K2d2FCtrPkuwVXgkA/X2ovzjhX5lWQXv1Zl892g4H+cClCrWoO6qmrpOl
DM2ZHqBMP0aUMDZ9h6/Zc/EBNvDLYze02mBi9D8dFQhwnse0vd9B66mBiw3IrRyA
Zubgp4Zp0lezkS0yeBQxqZX/HDi3hIIVvDmEy+huqO0A9OGmDmks8rAbkCi5ImtT
ee9ru55j1gUkwV+OYt2r3BWKjRqS6sLJbDLgoIXB4U4NVP5d42nvXlSb0qDtvlwW
lrD00GxXE0BDn9e+F6Q3uOLOOkWRHV+K1Agp0WkpAVqGRBrKrl0LV8Ej6FRc4mnH
nfwzKqu17YMzSH5x+59/BWCTbqIoWxtoXIXjKwmUPDRYpTMjmH74sPtJ3VloyW7m
3UQAU/DLhZ8nPiSZvnVLdC6SEz8mLc+ox1ILqdTKlmnqN6vLTEVyspq8WD1FZDDw
kHxd3rHnFoaOs8UO1H5Cls56+oRBzEqpxjufNhNu8Isde3XngGMTRUPBgEwx16uO
GtQgc5Bs3O/VwTU+jGJizw==
`protect END_PROTECTED
