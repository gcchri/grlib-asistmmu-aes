`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WN3VqNai6oN2SyjNfmuEk//o08OfwWEKH86hSFXQHsEXFm7ylPKn9zcsq1oiOfzC
x+5+wan1vS8sQjiE2kzeDJgTdKl65APcL+FLj5DzxjrkuNCepDF/Xs69NYQDNgaj
6I3GfJYl6GYzJ0GMS4LBRDEhCGpSm5HHe6zpQz3frFqBesuTKd9v8p3eBPWdb2gt
R9nZAFvLeulP4RIdrVZkyTFL6qlv834NGHA4LwDSTxr48JbW09hpRJyn47kwCWMP
A6IGL5UWjiK3MFaoiJV4jDzPzCGmlPpOg0a4i41nuADFjPYdgiVnHQ9VeP+95hiX
TTCcVEHcsCSZ62pZhT/LNbUCIDZQV767ihpdvGj3hwdLQv495w2WgrT1koJHPhv6
w/X1fbLgpbNQrEEIeYZfwoPBvikSumfTXjUnHbiqHbhKgFKxBCssfdNYx/7yGJGB
Vz0hesygQwOZQoXrhob8zQafh41lN+IPF9R/p8MFUryOdI8v1yi1bWujwfOztBCE
lt6P7gB9Ed9nQEYbATBB49JZWrmQCVSAwQoveEeIEzIb+EQ9CwSXpJ1u6bsA/w7H
H5oyD850EuUEUSPXNWYKvOyiKrIdg7Ngm4aeFsxkUJROetEBCEVYxKA8V8CIcBC1
rExLkf3x/1NEQZiQ6XagZLFGS0j819yCjOmkG+U0k7RQGYBxNLvnWu29urj9SnpP
cWT3+7sUcYJIowBWZz3VSDkPiM0XjV4q9jFhKYcsYUlTqq/anzmorZEaMlXxMoil
krH5qx3Auuxr+BwpSKf1PmLpF9zhRS2iD12lGYaLgyFzkoK3RUZ6uAeUfXWUEeE+
hMaJsOEYyydtt06kgu1/npM0tbnZx0USxM7eEjcWXYM6FhtXev8ex1TDGUSh0edl
71VhOOzrFD5fMPo1plQi0Ir0VX+jkT4o9rrUE1YEWF19+9wPH/TxCuoHwiLSCCjZ
A/Cqgy6ATThtf+Fndvw+7AAsOLsIXqlSJkV2+HAJ4jpyj42vbgPbUZDjXsNDQchg
4R3vLZfBQMj2AG+akSBQwvQ1Yum9IhiSdHopJNsmR27qCjOJoXyT/o2Dybpv09QS
VluRLRq1mj4Tp6SWIQPkjvGUN97zgzoPv+AgUsPUgqtx8By/BNMnHZ0VjG6dZZj4
Pz2u1o7E6sEP5MIwGLbmcMSQAiEm9RM+hX0fv4y09d06CPb2yOfYXaolkV2ysam4
1w8ztDtBxvX2Js25GkQmgFD4yBPr0cCw09cFV1Td1umki++2mMp+g/JOUEWIBMLn
U5vXbusTgC1scuLeIcgxPY6konjyMOTaVH4c+QFDgXnmOl9AaQwaF6u9XRsFSPEQ
nYA4H7VraBJNOCrn1VpQMct0d/2I2X3++tQUj3/ijQVG4N2oyJJAPUL/EY4jZqsZ
tV/WDnOFLjQngJhn20n5vTl6BkQYUlO97PlUzurddLQ=
`protect END_PROTECTED
