`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4cmlTgAaqTLKi2A4HuoAomCTngsvhj3jncxhrze/YhN40CN66d7TUEA2FCv0KYLA
v1A+oSJzDj7bqavfOCeHz+0ImLmiHgkd2yFcHqlNk1CG7BjWNZiVG4JIy/4ufeCO
R4sdDsZvMwcwpiTDs2jlrsbvqQQJfbfTzPJ8E2qZFuCrXAfs41AQYTIjsgImgvCY
5UR4SrmCFgVx6EzGqtIYXQQGowjDIPiZrbVOLiR37ljr28PsNHbx+nQjMCMdtrkt
IaDJRFh9kUJIKbi4aHVPCM5iBITPPUjHvOQxr/J6fwQFYnbTbuitLdi0o1Ml6b1W
H1LKZ2IxgGLAaF2K/oNrNSoQxd7d1IR5A9KQUaIXxnafqJXyHn0OjG0WUFLkfDWu
z44fw24d4wnbupaNVMdW48Em4tW21Uwbqo110XVnLe+Ib8aL/26teYzb9iOgtEBL
uQDLc6Y1Xr2nPna32xtn61xCZbRahYd2+hEPrk9fe4yzSjwW6KSsMk/VWxeLuPej
ZaivUR/Hr7QVYRvi6QvfQV+8BHdbdO+CmDDxRprEwS6J+44D4Q3WPYrZoI1oYqBJ
JB8x336cln2+8sNr+rUb+iQOGteRHuKz/ukfYyQhihGXtvLABFpFdGqKLthrT3L5
F5sUfQC68v1ysIAe/NP0ualsk6IFIHIG9Yy9ukhvvdwlMaXknf5t4xXWKZINbfQd
bv5vJaqy1mSaXAjoeJkUUA2n81ItVeyOq79p5DIejNDFJDL8PuIpSJ5PGVKDgFn1
8s6RjaOoXXONGlsStC9b4Cbu69ozSaKU0+XhQzi92r/r35XezVnMVNRXolCE1mOk
23rFh+CNHwrgRswMD8XS0OcGPiKTVEnQVF8nwdT/wJTXihe0v11reyPAw9ymOHRz
y5yX9XQsbrIRJRpEAAqkl6CIGLMK7z0eal75ZUzeSUYpgCRpN4x6t6H0Musns4HU
jT3r6C7lxkC79ckDF3+aA16xZ5p7W7wek2Y4s5jNRAytaHMBpCT1tDpo5RaL+kIq
MzXo/kHjxFli0svJrgFxYZffsHobKEPdiRwj9kjswuz+10vkDVdviYfoBo0iPF1G
OIMy17q8z35Am6IjvxKyWRsZ6v89wjpYzcM5mLrxWNmJvOnY4HNdJemY/h/+n1pR
Xzm3EudI+Q20LiTByV5ixhn6scf2MLrYa1nj4hWxSA8P+24KOA6ohDxAavKMuih2
WnW2NM/yiG+G6olBQNyZlvDap+9NPUlJCZVw1yK0A9NPr5oScymOyHNivN6b25JY
7t1w0Ze33GMCkIzJyi9HQ/C8n+159GpF3ImEgAj7ePBkhPWmRwCYi4DrABIF1yXP
vtn0OgQllYseloOEpmgx7dLW/5JPELqNvshRo1Iqr3FTnjRMJvzZj0yhsNwhpy3S
aV7DCuQQitMVHfvcda4q2bXNRdtgG++BtsNJkN4CDIEmHv+EJ11JOkM1s3zXbJpM
lOrNsXxDqeWwmvK41/jRrvGNiobgbbvA76XhMAlezmMDJW5tvZo4ywpZCisVKvct
ehy8qMjZcoB66ngun5Nm9xwnMhRWrHzarpE3QepE4lOqLUOsKV62f1DYOmqHgdZ0
h836y9Yew8VxJMFrj7aHYPYI4R9jFLnH9FzheSEoXHavUMUQ/6Iwph/Uderz2qbG
iAGaOSBTAzi54d5HuB/Zr1gaqw1MVxiXcTFcAdfvheenkeyDe5F3jVXQo1ZG/6VC
JIyK7J/kk9rKEk9Jt9xmXqOtcvlDX20OCiEZF3gbWsQmn3fd0w38N6iFyC0SUfmL
/RARJuviRofQn040/23FZ3TDzAa4tl3GCa62jto4dVp7PJKYH4NEdzf/ttRP3cLD
OEkm4//9KXVjC8lp/J1hXRPMdnqBdfhY3SckL90dZF5AJQCuRGJcC3UTs7ZEthKR
R0fUp1v7hbRoMSpccP/B89b0KEeMSY8fSV+aWayTAlF172mH95nheNnrjk7LCr8U
S80eXc6Mf7JkzWaztUGZqPMynFV71lREmqgNZkffob69tL2mL5Yp8aj9i6mE/UQB
IavUEOrcl29bQVrVdGCziw6ai0TDYVyL/NLm5huvsnCasKcuvAsltwEVq+Nl/+1L
XcPdLf78pGhBWZtVRCLsYn8XUgMHCwYhw0GvnAY1Tp9Vzg2wLeJZaNiOp1N6Ys3b
YCgTQ6JQbBzBqDfWUZhinVNNl7l0cPr4aRTxbgZPv9jtSuRMSjS+MldbCHT8Li/i
iyGq3yaPEDMZgAJcj2YxkUDCRcLvpUrvKGMxNPHISPqoFv3Duqkw1BnOXC0S7vMK
SN+k/oE1J+mFZqSIv5vdfunDN/q+vBOylDIfKTToBP5bin6TANrGMrKXjMKzgJQt
LfuNgX0S64GzWvmzg+SUkmY2phtuaty69lXIqB84gmbfz4C/+XTvQYVpJigdh6wX
aaTQ8UVoOucl6fSrIUAJmmeENwr8MgWwerdFBoX7jXzNNUoDPpsknYYu0XcGR/ss
NNTpiWcf+K3RD4R+0zmgE7xtpQnrJvuBQA9G2+VtsyN8NamuzUkG2M+JsTMqzzJP
JkgQCuAmt+jv8rSPEMsciYqjQijR+lkB+InTOw9AKspaLjKql1J4QNstPQtrxo2w
qh7zQER1qcSkNmEt4Hfqzo5RnmG4fexHPMIoKHn4AQwdDEk67ZlCNI/Jxe3B7Qvl
EDxXMpbf/tBPIKeoLIeupPJ1MymMTxt4SqqPEhdLmZUt6N85SHGXOWlV/Dz7aEAi
Hm1pAITYa/7+mIubhIPrsPrjuEhy/XLJ8HjW13wfno6e2RJ6At5bwJikOcwYZ7wN
pnc6YlzVzwssoau3mWn2lAqeXp7gQIf9i1xaNlYidECHgrl36tDnn+O4dEUqy8oG
1zo+qMOZZGqzHgxdnbGLVMk1e+jXQAETrFxoIRCDihTzPuixqix3jdT+s+d/yEvG
XpNMzO0b1liBtWvGk3AMpfvx+I2jnNSN+UL76Sn/wjHle0B+pchtz/yruIlBvsWL
DS9nYHsnaCNlJt5HbY9tHMf/8ewf02GDqLseSgFXNkelur5L+iTa0M64VBKWMJsF
KXiIANuia0PNUmaouODjBMirg9QFNLlelzQd9v9FwDjauDol+dwiy9B+fcfkcPzW
Zv1q8i+hsvB6z2nGHjMIRHbTwWs31l/A+XqTuEw/DAazN0Odd1wX5hvTgSYtigLl
pVhxYPZxYY8zHuytzW1ZZHwY2ufUyX9cKR9vbdhtPA01coKLB3YXDW9wjoBuco7W
7YCk6YAlmEswfez5gM92BMMHPK1KNeMitGe788yVE/7JPi400jKR9aP8JFbpjZiQ
Tg45uRRMGF6i4COBtHlwfWkxGAvOyrQDbo/vr6eRTpGI/nwJR0qqTA4w+PQJZUaB
UuaW5qf+TF+zqiI7kX5wWZcGPv4HQFroHEBpUdkgWdwhzbWGEetvGE/1qmOGKmnc
U+6nrYsNjziA0ToNozV14HlpYycrMPlH6BUHh9waqfysdaLA2g8LizIkwfXB80I/
RKogXRVCLCwaqV+TKVYOV4nUvLz4TAiokk+BTIMfsgKlEPdgR8CNeW2eHT4rnKrN
ZEaFE2v0L13nHDkoHPqNpBetAqWDFEoB4Z8vPfGzbxMgNACA0EDcqX4zgJwK8Jiq
H2XqGCvk/fLUi/5Dvruzhg==
`protect END_PROTECTED
