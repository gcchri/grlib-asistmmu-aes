`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q/U/+CnGfXk6BpkDD27LltBMs5WHRXEz4ZSGCeYQnMIid4KL/Ttx+8UW1uCizlbk
olmgU02zFin4Z/b8m9xoQbUt2veb9qMUtqcfdA6LWUSyF4GScfHh1empoyDvqKO2
V3Rg21/RVr6WBHyXF54uz8sN382jR2RSfJfMc8n6vC4XvVdjm9EChOf0Bxk8HI8Z
yXZ+GcUP6pFA4WGWcswf0kpBleyIFXFg1afyxLxuunZCEeZj6xrt4rw3lG7GyIUZ
J2chO0NME5sol7WNyi9hAhZVyKXcviY4aP7teuy3DJtrVAVCIRjniUijLyTsya4h
Ic1L6zpAl/iml5AkEnTZahzR4I9Oxx8x1gCR5tX9XQSq1+tsYzTrKKPZsVLksQZB
gJ73vcp1hPNbO9YVANtq3wSXU+PTOgz0eRKYpLNDmBTAr20MeWjZukcaf3rfrRNu
9qtKfbRTeasTS8NDQKq+ppKfsYOUhjdNrwCxbsflocODrdJz5kG7LW/Fv2kP+mbi
6IB8F/Q2wFRmzzLoEZvp/N2p+HO+wb9qiL5aKP8f/9ewy3G1X6Q3408lprZYdg6C
rveHl9TUly4yAfnprW9aCBLnCuKf+qL4FjtXewzlb+XJVx4i1LI56205l2MzNz8g
HYqQtvKM6IgrjE96cmw9VhH2BCgGTso5TLOw/B2UnUk7QFXr+qCK848Ok6l/RVzJ
is88O9FAasnlwaH3FkG7lrL/v8o76mDPa/cG2qgbY3SmqAxwX0eAIXkmJwrfthce
60QryNcaPT18Lw8NK2uaOA/JGqaxoR8/58BwHQhDJsUHXwJK+Z3fS2uq6hZGGW8X
8SpKAcP4Fp4UIx161DoygfCi9i2RKIXnC0LtO/b5Yxr6EUYE0I/sFKPKdyR4vUYE
e3+VeFDEAK9bAgV7f4I+9kkgc1A5q2jOIEtjSWsynsLKYXXJuhYEkUi9HVVGNWhD
loR8k9i9HUOclASuP4uj7zlvJCaV19pik0wvnbeGQ9q196iv+t7f4BHau/zOa2gw
veWR8sehAPkDeQk7Px3kAqBY9XFcpoZlfJBlj1+kCNHkY3jm3pQM5CxDZPm/ygnh
uXz/2DEgXUsLkEQ/DAILbfamfu2ob0IZQysamTH71jrxl2o7spqDiSxRAED0DW4P
9h6GJXcTj2iy0YQarx7jQR7OkKcrg60/f5baUEOWVl5BMcWAkuNcze3HcVUuRAnp
1EOSYRZQeWkGhBjcfj/nC1LShWfZf/e2rcmeawMT24Ybw3J/TyKUYeMGVCT+8kGB
+67/XQkixqv0u3EpAsW+xNrZayiG0znHJhbBOHRQUmwCqFdnhFMP5KG2k6OLylB6
mDzEvULHocVlNKDqTEzN8AdY5HPn6pRffmBsqDFDRJ58vwvhC+iwyqli2iRFKtG2
iU8Rf4bA6x0olf0Qpb8KsIm5fCKkXptBB/qeWMTOoTZiNhcuN5otS6PZ5HYJqGJY
k0phheS3/kZHyBxxE0fXeRlagu9eDuatbdlipgDApyczRlOOrvNJWLJYERDTc4t+
xFtQVufBxLpQgTfaxj5DNVHD9hIzBQUlGXMkWuTHIH+dU3N1Lq42rk1XeHUVVock
VbgbLy3oNlYkC5tt47bB5vP1/vw0mOjj/PPUZ6h2L35zxV6znJS+M8dfGuRSW7g2
XYPuqxTQwRCYqXQLVS5E7nrXNydU4CJDYdV61nZEfssVsfcO0X5QG9akwirZfkN7
hjqfr8Z5VoKiGpJFOVTRO7e+DuZOxoJ423HetF6lczCzE5+FS1g4/xQLBOeXR9Ap
NbLS+FCSpfTIFcFxVAT7Uk4oJH0s4QsgOfqDGJvkFNTaJnl3gXKMhX8sWsr3DZ51
eGRPylmskr17/9U90PXK5hzNa5kxRufCsxEnANgTgPRrrjQZ9keyvLZH0e3nLBxb
B5txChDr0W8J3RYgrymX5bBwUYK0qbZWa1KdEMVMoKYV6IEsbiG2BqAnY6ion4VW
R7L1GTtxXVmniJb3JIP8BAPu8yf7TQRJepg8/PBMl1HT5pGHKpdIUxWyXfgVOULQ
Q9Hfl3XGRmAcH1y+20CUIuJ40ZUY6f6JWbn2LK8bGdCBhjjHNJhPLk+tq0VSlljG
uDOKk64NQGGsXqWCkbsnJTFyAFOljg6rRwldMlzg4eziMBqNUgY9pvpoZsx82PeT
x9kWxzlDZCN+PC5o3Ts1HRb6Lg3u244tio6rm17d2ipDdvsf2G7yysjEmDmF4tpX
tQyKLcKnWhrFvKcRdGtIAIu7NRvLP7gkFR7oST4xgySdUu3D7E7TxQLer6LIxLu0
ZqibOWOyEXo4fpaR1TYIskWYoYJRgJnUyTnyT+CwnspiyDHSz+ZH2Xld+/dg52J3
4/kyn0EaYh+O13EVDUlQLxjzG1vBh7Y0g4CXiIQRHrwkodpd19pqIfwWG04ndLH6
4mO/5NZQTHrvPyDWIJ7mk/vDOyis0rKSOeogHNE9/D5au3jL6IFaiF2NCQVM3rKT
BcRmJtKnniU5cmnMRBEVLawxQl37uAQFPZSLrTVEVyO5NmS/Wi9gfY2y8UHRbkYR
HFYYtgyVWAusYgwLY/vDYKTRRhxChGgV85NFzgeNvNByxt0ICAehRlRV1p5Iqkgl
M7eC5Ms8JcoRWm8d12SXX/3TsESrnR2hi0ck/fHQR0mvAG9UMye8pGI85xyHTYgn
Pp5r+8ej/tYVMSSb2L6kRrXjO9W2uaojUsjqDg/AS3sB8WkdLqSq8jxiLKRbs7PM
0CsdtZyYTIa26P0z44dAQhDgC6U1Emaw+idvgBH1QtI83WvNYDEGugR1eKqJGpjU
fUwkT8vUS5fXvazWP1YoQ/4UcuEougBqt7MqxWNXV/WsktBpwtx2n9iTjB8245Kr
Q6eanlzkFYJWJTmIwBz0TW1l7+dFTbPtadCwNmGYwbgDKodM1PbPtOuZW2Znu9is
S9sYYiy0vcQtDY+RtUGDNiqKJjTd7Q2a5EdimUw8W0Im+/8Yro+rse7hb5AYratT
5/+koBLox/Gf66Mf2wb7lpBx8QOZdx/WkbAGLlIbqMyhJcBxx/ZiuzKECnXtXDMO
eyR0tuqzxQsqhsyoDaTK7BXqTMTJMXPmKb28561e0mZ4NLHssvmhsGSjhkBVbMm2
3dJ1oRMR/qhvkqUshv0XzwCHMX2iNT3JrDOAxiqMHOdW2DAOAv0dM9LkZjXNcWSQ
0hDeEYoxpw8RTLA9WPHDIByYMyqnDQfAd5TbAWwQ84xS1W6dJNlLmeFCXbJyCWVs
C2XFtq6B1sS26z22xHNuBPsPlRquORF4wTVNc4ReJO5h6MEFb5S+QVWtWQCIi+Ez
ChlDWkgu/NbVpwzbVJcYly3meHtuDR9WTiel20TsT6kQPGrycBWRuGX2ZLPdElxr
BiCgDnxSgfZGfMCWwLEDGAfzTh2RMQeEYiaFGKliNfagTwtmvn5EAvdQqLrracyJ
nP3fQSrqh/3fYwBa3uAOi0inPqSkT4TJnQIuINYMwNaoVjd2V2X9XsCKh+UoyRRs
s1fhmMh+kFUkHX96OMEYu7SyY/IXbSCfFoKTxVZuHQ4Q8v+xDKopoGXialOTFwWi
WYnOK2tM6g9J328zwr9ynpyrEyzAFfutSXOX4ZwS2WeKQfI01vtH0WpejQ9YTb4N
mcXShaKZbhvqz1HgbicIyBJ4ZC8jZBIimKKVTt2IEUMMPisDHN/LT3PPLYu/lDf1
iMZ6TTNwn645F+NIyn2eoq5Cn6oSnwKAqdrdym7sdUlXX3znc07sKDXM8eiBFHiG
f4xASkOYMPzxa3gkAVRSSI/v90hRmYyXWUPkaJEfrv1quhZbhch2YQ8tpvmQ2his
9wTfSAH1jVkspuSqbZ6it/ulHsypPB4nurZrbVFV+Nw/KzBvoptp3HTsceL6mmqg
OsfByOXTaGm+eUJ/+edl+9ftbwj198AWqZNUwMYrFudT4ElJHwWW6zi0HOExy4JB
hfnSuaNXALt+oO2hKDSr04UKPkPoN2h3LoIz9fwGA85jvLfq/6xL85KQVc3xpwd2
0B/Zz6C3SbtvDICptWZgxh2+Ytr42Fzw7wVojdip65IHgevPDMX5apMhHTrUmEve
Bbn4TKIEY+S3YGaI/zmspPYXybQpCRs/VzbExxJBZ78dOF6bdBBE1n9B85VKzcxp
rvGcp2hFyF6tICBWQrvr/r3maJQ2xtTqhXmaf2kOAGoiUpEre+q/LAMvupeT5hNT
OBeX9SONGP/ZxS6z4xo35g==
`protect END_PROTECTED
