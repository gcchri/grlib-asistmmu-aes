`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ij1gI/Le4lMSfm7SuxarUOs3iT8VqdtPCwWsyf4paTpr2A42EG/ly2k+hEnWPg8R
aI8SV6fxS/kcUOEtNQHrHbQJnPi6koVi50flcGUqV84jrJi3IoebsY59nsMcDFNb
xcgwMQXUzUkq6w1E9ooEft8nU+fU5vi1nGyEeuw2MX0hMo3hORVrDOAbiyEa/0R/
SJdh51zHviP68GrBVu+P4GhWv9pB6uSyqV7ovUNDi/wWVx4609/vGmAw4x7oBpoc
pTIrSficiKX6qtZ1X3ERA9t9skvS//8OOJJ9VbCBxr3JCpYvsLn8YaTFyxcn+E2g
og0WTx8YeXDsiJJvMdeUum2yaGOM1x0cBoFaM6eqg5lQJus867QYr3b6sYESaJzY
d823Tp2bRTySoMjcF5LNNnuaacs3k6eflt7xMekhR45ruIDMiubzH53jHxnO+aPA
5lVm3/Dw19AbxNbpb/B9FR89MdaXVo50O9ffNbxJcF6+D1MVH648gZC8BjcXmezD
SF93jZT6WDKL/HlPcj9p4g==
`protect END_PROTECTED
