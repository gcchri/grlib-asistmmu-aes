`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xd4ccFU5Cu8AKBQ+XqHwn0/9LFISxCYbG1vOK4sXs4ucfpfH2x+L2JEF9lZbwJfI
fg/UCMnyCIAKHyroUkjDq115myTM790H/arooLGK3DoYEa5i2qaYkpvjStNfjaRD
VXStLJrC8qTnkO477KcqdhzEH13uyXy9O/8fU+GD+S9ivPky6YvLUheFeIgL29T9
oOpb62VCGrmk8fZGMboUmTdZPMMANbz9t+nLkM1GdWcp9g/Y+fQh4Vt035EWcXIp
WO9uTLBuyY8kHgXanRsCLbCqV2+0tKCHDYLU7o3NcUWRe5aNSTUMpTe6mNAGay7x
JJVBXcWsQoJ9faQT1mizivoXJSr3LxHV0FMdV8zRM7ERbV2fJHqSBbYnRS3H8PEE
dAX9ZiN1P2eLeGDCq6/DFLRUybGAMuzscPVIQoci1ZCU1jyB5nxRsEkUbVtY4ur/
`protect END_PROTECTED
