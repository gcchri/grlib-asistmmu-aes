`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cyjJky+FuAzJIuBKOpxmY94OZM0miQIvtDaOS78EK58tIEKgKkYQ7NsqpG44Jdta
jKBlSqsMzy0CBealbs1hHSznCVpbQWTi1lO44E4Rx258efTTRQ6k+fcxuyh49zxt
nuJ2agpoUQWpPtCT0OFjyX7bqqeEz93ho4uB4RrYcYFl9LGmnXnmrKjBle5bvXjG
KUh97h578DtiGCKOoy8edojQgDBoC+YA0UrYKlTvSaD2pUujqQtOY5qF27AYnLnf
3ux9UN/3FyBG5wa6LVPe6ZtRmoXaA+IjGCJVRwO5tAd5DeSrA0UCbWmbzNMG95+u
BJ2HxnB09ja2WsYUs+ePiZHunpJkXrDBxW7ck/QsYdNJAnBoQbwTTzL+igBYJ8Zv
`protect END_PROTECTED
