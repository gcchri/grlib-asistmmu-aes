`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pluxqxQzzFdiXnw7ULCTkA0HQDjsAEzJvysGWjStcE66UIUvfYuFt4uT+Rrnp0WM
XUIbE8PrgdH8cJdT8vPDKvMPVbcQhJybnxSrSgcP4RsWKzO6vt9eTHYRv/2a4Dg1
6InZKRqxOvxupCFitguitGZSXllJFskshml0Vn+AgXTOAOM54nJODbPRDVS+J9DO
uomTMHe2KqEpmRtHybGi3D2Y9fmKh0rTWOVecmFnR8VbMExg9zM8++wasmYUwE4s
qW4ELb94b9GSZX02QNYrkOOf0CUX6PEZKYvbYdBbYA4HSsDjqpYN61KU+HbLeilh
1+Fcp4+xO9hIDjX/6D4RmKt1/QE1pLljrgUqDrQV8SacLbhsaz4ONQlC5IZiCOeq
1fAh4xaOQWSkC7yfdHYUgFDl3hCvbUDoqAvSf6bapuHIOa9I16Lby/H5oKGaKNvf
HF7LJBVCBGpPQ9s0bMwhLmJBmYfiC0aLQoSUP3QcytF8eIgobZ6s6pCDwCcbVrQI
L4wXGjA+/zOXE7eZTIUSmrykO8rHR6zpohmscG2NSwQ+Kth6rdbor3XOcwpmpyyn
j1OPJ9dMFjMEg71L76rAkLuK80iDWMe1ltak2CaGppo5JtppeYjsaoqpVKlxclS/
VwJFIPryCLhDk0od157Ug0y4pn//bVwv0V+42U6m6cNpIdM2OlCAljz0B/p9Nmli
lnHBXBZyJNSbtHCBQPtdZja7rUZoCFOFr6+PvnpJazD1KtyPIIaUuOW7GzJN/9iT
NnsQsM3ZZ2MLc2JxK/4kG08AcAhqGqH98YYyL2L4Wts7CpowRKewVnLebou+5PPn
swlNVnXckigF8eDXWxQ8IporR3SPlf/TTzZEVPsY0/mvlBvEb81bhegnAPE9nQVc
BGkQgaliApWj57fEPYrr9gJhr/8XaRG9J/k6o2aGuOLgTXinTaj4xnU69yrZb0rb
+e6mHyHNJqNMqZIBDMOK0s/8bbO80mWUMuUPMDR/6W7QqjsJAqfsOPCdK/5cVACs
TmA7ZTWP51qqWX+PY2IH4eTbe7in/P8sQ+uH37d78VyN47ma3QNAC3LXzuO2vpC7
QafMAY+sn9rqhFYDTNGGfG9tgYriQJdHm7JszN0IIg9k3+rISDK2xjNzP1B8yobo
tFZhHqPeu1Hx7nonS8ETdNtzGH5tb1pUgjkz3wKTuQOfFQuWXmwiWPWWNK8kWD+k
3iAmXpBTvvu3Ek5Y9gNk/mZ9rjHFKNb9yRlyHLmauJZzvJGt30XKrLero9mD9fHl
Kl47/FyIAy0w7IqVBm+46imVxNw02dDqK2S4ziqYdI27+4WSUy/ENzXa3g9UoHJB
XFS3FP0IzcUVFqCI1do5gbGljtMdrgTsTkJxZgMEGLSZN2hrMTKYSkAV1n7r8GqE
NSna2TUnnQzAucZOXdXUkhidU5PItt0057qGncmll136NfgbeCkNVQ0Qgaap4uYM
HlBjo+1HwffNZF5rQ6P3JHY9x3YPA8ZXbV49KhBWWEH1b95yzLC4vsvn6e3O6iaf
59rn40u8P/dTTYNqQnGWrdUkClkuJohiBcJPUb/0I0AI1FRscHtwo1VLL22lOTEl
5y54um7spdxnVZCEC/9yBI2Mb9hkE7l5HnFkXneHBJOO0g++4s/ozT9tuJReG9mc
LpbllhH3Jp4l8RUKfNL4JaQSO76okd9xSLURQBx4rF11QFXKDmF2od91+taHwrjQ
juOQLSqRdB2cOGmoaYd5d0jBFQfgoBZEzj70ne88+JfDTWVJhZ4Jms2sheLPEy1X
dttKyKWgD8zTKhApx3iZacXD7SnlKbFyLK+lGgB2KAJy6zSYsTCQJQofY3d8mJ1M
dP4LAjqTNYmftXmgV0jz09cQUVLRttJAhUK8Q2J2raxdxdi2FX6L81zvuzLfpcdk
oT6vrr151PRvDxQ8ZzLrsPdbvWmdpoxM/V+olfQxeJijJlv2X6ObQQfTYPAyI/Ea
aMuDJ3AA21CUlDcjcME+frD7B17twexO14qIJuNMjb9hxD1+SnCmGCeNn0Wm4vTU
939g16YGbv9B3+hW8EELZg==
`protect END_PROTECTED
