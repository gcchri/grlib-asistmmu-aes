`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lkuGX06zMh/Gi5x1bdiwfIzVFX3/0T9QZvnUqntIVsPgi6yW45k2syszRaMcr9Sj
4wokg61b2p90U74JI+CCKVzk7ov+VWsExg8WgY8D+9ujwGiLeP47ublsoo/7pV8+
hvYh5d6TWWghudGfv7/NcMT0tLu7LfY1PHDtefONI+fahZD/HsVJ1VUiktx+RAz3
bwD/lBoSeWqczfa5bKtgEpjr7m9bQnn7opSOLYH2gtEKFYoDXVGld2STTcMiNDKm
lfS0/1HHAaC8qAP6aMJ86+GeTKCXzyFeoMVB0L4fNjnE8bfpR8xLlHsluH5DlJ+V
oaS72tQVYA6/16BmkYLM9A==
`protect END_PROTECTED
