`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7NDdTSFwWGQV0gmLZiXP5xOuCUjblasahJbCjoPKHFXBRh7jMgYAoxZoKYzaflYs
HYKtGg65QOjvjgtyoZvh+0Lf41yrRwvaI/AaiNtl7Y8qJKHoekn9fILUZghAzyXc
lSsL85imPjTZNg94n/biR/nmUmSF5T5Bg9jarAkSMuI6KYZjf6fY3NaqA6Ne5spc
Le9CQ3auFuqPUbSonxA0/v1G7bHrij7mSLZJYq1lqPhntjkSHhkcOi0lz7bdRd6q
+NuR1oEcdQDx6FH07eUGa21MgiBFV+z3ku3jFALMp1NcSo/bi1C63kecE1wDtISL
ky+1ZenloIxqF725VSUVGx9lTeAomYwUzJIge/FyA01JLx6tfih/k/AgSIQ4ELaT
X5ccfrm4ArDaDi48XHutcdD/ypOdQEdJnEORXx82z22UY7x8HWVFuLjtnVkxz8nV
AOQrLi/NLI0JwQ8mkT+Q7PpGyz8t4+eJ7Zp0pVJQ4wrt6CorvyDJObw2O+/NxkZV
9Zn2TOuZTU30BhsqJMkmkXLGoO33PRmE+TwsJc3dp/qiNWA9ZBnKUm+twyi7+TG5
QPApHKXVPOcxZrmGVCfZE3agaQ9q3tYBx00HLZ3irT5d5exq8mPa9ZzbDpDzAsux
ODD7ca0+jvHQMfFDfh+HchzrbYSp5j3gYzaZGdFyYl5Cg2l29e3/NPI3HZAG8/S1
Ng5U6wrpg2KOGSc2ZpI5qyNKkWWYqDH/WfqIYrzBrNW4gz9IoWYVgh5hcoYitpiQ
Yf1waXWYW7uejjmPqBGmmuYSetnXtTps9ep34zKPSQ1VneNG9FMtOSt5F3pyCDR2
pJV99DIuFMcbK97W0UG+MkCgOE9tuBYidpiFFCLV1VZFuxDOM5koeEUPA0EDaIjf
yKlendnekCs8X711jqfU46cD42V0VyZ8yZE+/D0xFELkoin7lOv3/UkvQON9wXsB
xpyWkbDSSkDHPVd8G+f1KyRQ+e4BKwpxrkfmS//4/jHHuOecIcKAWyFqw5sU97Sl
ITOA2XCMTzvXFAFfT+Elh/9IC0Jhj8djcREuOETvlBnuqPbJfh+zAh5pfhIlNoGN
r9mwdP1uF+P+PdHy0feAqQOwPE6B/2lN2FlZi/OwufcjQyNYvJtwozPrAhtHlo0H
xEFP2gu4Iq3Rbq01yWJx3J7r7WvMI27o4vdHRupNkDIUTLMAnA5jzyKAaphwPCXR
OnAc6gYUVfTtoLHh3s16enFvn9f8mINy3AuS/+ig6wzn3KlL4KAIRnDHZCx7QBR6
sFt7OLsfqgQL/89If3SmD3y55JvfsWgX2cZIa5+NhUU7Mh9INTZNonm3uswxfFWs
Jhoh8ez9U51+h7tJvX5mMFMX4XICKQAdMOLBd+eHXgTJzy5vwrp9UQOVokFxqP9f
sT+Zmdl9qBO18NmV0E8+P9Ory3/KSWrzaRjei8GXfq3rxUuJokxsZpHm/Iq44P+X
SDWFucAGbidL8I3Y1hXBd4Lenh9LfoJHsl0c2gEOKQeiI8k3Y0pb4AzkbyX6eHBu
w1otdGIQeSLkfdVPaCtPaLTY8vKD4S9tpvbDfJZARDpx2R6OESVdjhG5uahU0MEv
TZXnfDwA6ZDY0lARfVcoGRT0R5zz8R8K0Xx0KmVngFKTT4KFUDLayBlxj5FInLJM
lKyd04a9eoCQ5NeN+mJKn5aqx+kqbHcLqfFK7w5CJdQQv+dtHrSa46CgyGt050hr
wdN1olJS3AF0GgmdRbhJP/haBw57ZZsCvpw9TwFqhr/v74QTSiKWHwNEt20Xm095
FGxDTQZXnoCLj8AZR79CkNn5hQdmQCvFKU52CVUkcudLba2DFAD6L+6/TCKPG+N+
NILqVAkgNmEuRu7ngGk7y+keUlBnkl9fl/8vltmn19CJNR2xHMYhah0gVNK932mx
2bxmrfNcaakjEVkSifIc5iHGBAX6/Lm0NJh7e17w2fBsfA1AL/FriGeKPXtIq/5X
w54TkXDW8FWfpzpFoCTv36OlhFqRHXOKLJ8FXxN1cdGUtXJ6+qpNeBCQ351Q6fJF
KynwbO32xLB0Zq6VfrRvQbw5E+Pu2NbnNpc68Bp8c6Q1IAqQLjsRchuSzVOg32kn
HNVgyrHRn7lsJ+GK5AXl5cS1SbZUbGHHrhOYqn1tpXz8ne/39X9CB/LjPMCkXoSX
oVGxwPoBhL4trFzz606HpBJ7c1GRFdZCFQe6fyeCgoXFgSvWg3o7v1Xd2bkCiscL
euUNdeHbu+5UkirjN/hetEnLolYE2rqXqk0+I1GwAqkd/Q3136vMRRUbisLT3eIS
B7rPAyzZA/bB0ZLsukUtY+myhAR/EF8IL2w1qVMjqUToiY3xSxcBXch2KqFgWpk5
5woMEf9K2t8ufEUHmbTsKy9BMfB6qQlq/CVARk6+mtGdkNz0jAN1oY+TIvRO+9Iz
VGu24Va0zNdMUKALgCh7rZyZ2BEG8UhHZ+qes1NWfZnmcdH6hgpEBDUnxlNzl/N6
lS8pfP6D9JbW4kI+Oq2A41jB8XkPxeIf798W03czofNalNJ72CsGNFxCXTFMLmZP
hwUpOQTEsoLqG6J4aZ4kyhFB/T6Gi1azgGK5LmbIj7lnJYaFhbZW5y5Pxz3QNnE2
mPH79IKtd1lOSH4LLF0ss1VOLsf6rLzHUPd/aZB3BFRGaWe8m61R2lgPnuWhNjDI
23rkBWpZVa6tTS0kS5YfY/5fTIGVoV5xE6gQWgnghLbJjZUkTWmrrnnr73JBqc4b
49/YHW9w5JOzA3rIXbxBSLviKF/jGQeZkGqMUGd7jyGQN5JmtGWEpRHfCD02PJh5
oekl1Q5iueDOz+24iNQQFr9Y3NOw1So9yYQuiPdCQu2J63tiPiqdf9l9byrouwVR
qKwg+b8YRSzv4uMxobjPl8q2g0d+taHxeC5OGAVQwn8jVFD3Bw1b1SsnB/x6Awhr
YrIcgOXRn7ISc5MAFlMlTZsHEEwMDGyMUG61Waoh5zj2EttNgr62dpJAitD6lP0k
eTgrRNx6gTdrYGnSCNsv5eC/eV5dJt5hv54ZSalOX0XsCDfofeySwjP4gGteo8U4
b/V2uAEChVkFPnjXxCmPrS28lrW/lzLmi+STZ+nXL+i7DuoTa3ZSM+VRx7UMYKcZ
w5EvqkKaR0BJvNUSjnqQI5mSByjPtwxn9NAIrIYHgj1QZCaaSjQhq2yCaDqxG0LR
CxWiqnQr9elXK7YtKHLkAS7Lo37oqOES10MdoWixz8qeOu6lvmNLywtCoqv9ARhN
HWw8ZDivVHlFfWbnzpn6a3Ul2tNj0dIJvbg05A3LhJpFkutJ43q/DoDEW88IoyoC
C+0JY7yWObumXHHvP1sDIy6e1LibNrVMVep0HUAr5dFtnYzvmMbv+mUuWZL29TRM
v6AJ3Fl3EuWYD0z4xmBEDVlPZ41Tu/EJkglwErp3563pjt+04ewQTQ7JV/EjpleL
R2U+fRL+JWM/Qz3n/cQJVnUBqsyobF1IQipHwA9gy0VJ+wkWir7cvfeu8ebFXy9R
lCEhJCccsAOJckpAfxquQg69cRlGNSpT5MluAOkQTopuKngKIL7LimrF3m0cqD0I
hoZ5zCYi2LTNGn2wSvQHSvOryA60viPPQJv5GtBaSiU4m3rmp7dtz2+MZuqWzPYj
/LWNc7vFvdMu0DVvcsUpqdhfA96eIWqHvMIECHFwstS3lSRfwMkONAWM7hx94WoN
6j01/KPOSjX2Xdh6qgKIrnOKHyWUuktZsQEe0ru2NLYr5ZdYyQq/GyuI8ZJ3cac4
qVQVUWcjY4lGjuXY7ozEJayNDhoP1q7Cs7ch2Ai7/kHpqQdH7GIPTt9QqIQREa28
vt1N/PX/oJKUZg9cg+Pc4xZ0exdpgzIsOaPal4axTpeq/1V9FMDimBDDOh0jDFX0
3v4XGTC6HskuwzK50DLiEIw+hKGg9erbgkLkCFpwUTQsGuC1u0IB93rr5/tbg5/d
SrkJwofIEzCXtKqYbw2gQvquQNORuDWqCsTPXCMfQfC6pmHwpT9FYOX/Ms/9e7K6
HfqNLiVUtfypiiL/7F86jq3/smktNZVd21QR3P3vBei3kWDp+1Wa1VMZmGq8wl5G
MHytZRtWnQdWc2UcJ2/9Du2oS1zxv2++KXkrV7sPh+xVErbbiep8DCSUUbeJ4MXE
l2pZgAQ1onLlilyQou5g7o0PuA4alTIHA8VvvBQ14nvFcD0mAgtvOqF4UuWDgZT2
l3mSlNF+CIxhayjfydyO8cqgfOB4kuNL+xtwNbGsDiDM7ZVXC+ab7MG1rVkM/2yE
moKaCvEeO+zt1zi5c4ntldQjWzjYzKJmcCIzR1HG1T5eyZK9FJqfW7xFu3sV9DM1
`protect END_PROTECTED
