`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rxur+KClNKUm+lMbY18u/eV5rE+qrDVWuWPx34clG7XGDFnNO4o0OdcOpoBtGKIZ
81f6mD0evSqJabsX+oLRHUNbLfE+HeSLe7ZPfwilMHEuvSqzJ0aRYP7cicXHPRcC
C4JhQLC5xYJa7shYGpJf6MZb6tECjHIgCJUeIzhZYStihEryu3mtSJU0FDRVLSHI
86tx4wDgAL/1xd0+VrVWQtR0+dViR19dmCuScqu7nwGO+8QprCajcDJCFeF71LSp
J/06x2Fewetex1ZH0W0J2VoldwUuxeVFWPZwNASsZEZU851tefqZX3PS+eMuU3XG
hMgMPRkW0KIxV3+jDsojdp5E3xNSEExmtgt0+JOfCNH6sw4Wb+wGsVkBdSNyUe0v
/Sg4GCRCfVIa9jztfWhTHgxKdoGBiBi2PzQYz+gQL/UH2Su51q73obomxZm1rQoV
D6gR38yNOwrLX8HQKJvBdPVWTTMYJBHynm9w8Dlgidw=
`protect END_PROTECTED
