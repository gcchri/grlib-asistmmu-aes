`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G5UX1rfGGDOSQqtaAgCLMgPbPGIF1of1JEz4xQdL+d4XidJBDPe2P+50Lzb47fnE
pFcvc/2PgX9QClrdCqdMC7I8WB5o+za0SW46lGwlyugPkmCt2H1iI1j5qUxW7zEG
y4DLof5JEKB9L4bKHDWMGEc/7UVG3dK7DsTN+I318Y0h3jkW9BLKdTs28uwPH7nE
mJodUB6FzbdfDIhOk9HPbLg6R0EHOAhgGRFeKjET4zkbqRgT1ROotDSOzwtka5XX
BGP0iFNGLF2nQzxEx06MxIZYvMS/+2xECa9zGD6iCrI=
`protect END_PROTECTED
