`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H+ebZLq51A0tOBnjET7AJQEgfXe3m4ccI96RYGsZYZT+RP1WoS7BkaBPYswqzcY/
m2hr3FDyOxN9ZbkHtmCOKBRDZEdq/biI4GZT5DrR2PgKQR1hPidNu1MeTPZUfL94
besVzw7OHl+NcbSALH+H2YdFclRv+5ENsr2BJq+IO8k+PaYwnP4RMkLePaU+8FSg
W9NgEpPTQoVuSTh8lBEPNUKkz0YpqKHNfE0kaJTMuVa9rla4KldNTCrX4wLCGJ7v
6E1GlgXlnTXN6VaXD7SXLy2a1S6y70zdxkwEhcIGBmlCUfyOW8fJW+tEKS3joSOq
FDY4YtqEBvjP1oo7lE1wDg==
`protect END_PROTECTED
