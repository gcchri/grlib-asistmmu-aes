`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GjooN89IM2eWi9uu3fo7CdqRKSiOYARtpg48Rp6OjFboxZivTBxj9/FlDDrmrjZb
6WcAnlhuf2hUSVwkb4zw6+CaFq3V6gWA/RSQrRALryPgcPc0Hzzt6dUvN6UhhPNw
dxXVjn2/l+UrvsipHNPN2wBY3/+t/mI8LzCa6N+7ZJfNYhgKr/aIH3wNd19Vdg32
K11cetwjFE3Hu3H5kBE+ymyY8UKhxuo9vuTt8Tf347KGSSOc91wCUXTGE2teVXWR
kHOxUs4NVtPgoPxNj8gWX7rYhcbFZClnCxYOdEwjdN4SfZqvclQ69DuY9aGl1cJC
j/VJdSUXMvO53PHfu4M1Iak/3u+8KuOSxxRMZJ9cbO2EyLC3D6fDfa/7+FUYUYCe
tmcSOcvJia0Hi+XMezD8ikQ6qPQIBK4tyA/cEqfl3P8=
`protect END_PROTECTED
