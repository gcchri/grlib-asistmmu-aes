`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y+Kb4gTX7Yi//oXrMZat9SEXRO2frNmS7136KuscGhKNRTnzYm2+n2vzp5+Gnknt
aNQ5hB0TK8EBUxfYjj1Ma4+COsqJSoTIeZgRZW+X/AacML9dumavBTmNzDTWR5SR
zm3MdueP+eP0Fcg/A744GWTFKwQP9rSvIxRTFt+WIYHX5LdBkMz6YXRddpPWmVLO
P6cv5/toZlwwmazTnovWP8JvSEd+Ibwybl1o/5hCWPguDS7B9gpOCkGKaOYG47gg
Lws52Q6QCoyw68ECWyBm3tX7PfsAXlPrdr8CTKJAFNjvntD1eqgeHZkU4emCkckN
pMT6pGcguAaabxIWz8baJ3Z4lqKpfTkT1glwFCILGTGovXpuyaGAjO65EEnZufZO
8e1ZjGvsA84qaYIs+a8N/3dcwi5vpTJ79lgv/dMPptnMV6//LzZpqpYJzzbHSnfH
z9eyILVwF68+eM3GesDshPlxTJAgWFCJf0fOUCrC8GLG9omI9Wm40F0tE/YKcVIC
2xzicXLqxc3+DSEVmMCWeni58nBIOIvp6TGpnULI0XV8NTDgzL1LhgkRa/YTdAFV
pxr38hnrP06KkMlA7RNymcOlpuBSXg1B0XzGiU6YEC1/XmVk3jI7eugFDmatRFx4
FLBAiGd3wJZ/9JRYZIyIoFLwoN7hLRDcteI3ZkuY+Yu+8wMn2mZ8YEkytAXPGFXp
qbJ2Dwdvx6mir5cfcYExybygmk5MKh0h2daFAkyBpuYl/38F+lUF1rmBUr2A3cDI
FO1S3NPWaPT1opNWiN5YmNKwSoZdq/Bc5l0dNcGKj/WNhzS1htdmwqZCEq5jywGb
oiE6oobLqXZsxgisyiEQ+gc5Ax3cLd5KYt/N+fRJZb5JxPmEYegw8wPj9sqAMH77
W09XaaPK8J0oZARSVyr2FeKed+eQg0A6AIigMVaoKK8rfWUk3d/4HnOHaOljd7Cs
GQxRvfKfbm9pbpD5i6hjpbvorBoNYOGHTgyFrA64Dm9FL0iDxbAQ01OXuJKIBvBx
bKQ5R8+dDWzKndDtKR/CYgsXgmFGMt/uHYwkuMyfylc=
`protect END_PROTECTED
