`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6sFlxrmda3Nt23rNxM/4Be7uPNZTvCC5pvGjQSebYtXxPHwc13lN7vaYThyGKs/M
bGrxWG7faWgo8Z4Nj48ExAy/yo10jKk2Wfu1zKWemuT8KPn8zSM+av465I1pN4bB
jU/XLNgI8RzOyNOfU92kbTwOX997r0cwuYRrU8w8wkNmB3BQ66xTuqAMBsoSXdT6
SI7RRmy+wdrGlMKpmNYf2JpsxWYEYIOLMYtdYpOF4ka4mSltkrSBz/RF9UQfyJq3
hIGeqEeJmvzD5Pi3BKhqupaQAC4VdiX2IzEtm2F2GY8eOvd/2RcU7RWSGyokVshU
pTUnka7rnW9il/eIY2V1vjoM83XKoGn28/PQJW/SFna9V1rbu4mbF8fiVE8t6inf
abfvDUsbhmg8L2TR5xiuf6R1s6QHy6AYm+7bbSx6KKI=
`protect END_PROTECTED
