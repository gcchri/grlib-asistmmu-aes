`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IBrr79K/J1zjpgDD5KozRTZqKw1a1x8zrUnQMtxx84md943aPuFhFscBqYSeUac3
ri9qx8TLvfFUXhwn+IyK3McbL+nma2+SUA9ia/9xjvOGL2oRB5QxOVsbsVSzpYj8
mOcoVxNk4gPaSHL5R84G99TnJDKRNNdcOtT5y7DEmKUyQ2L9OX/UIvPtpft9dMxk
kHiUp7xLVj+d4jRo3RexIx4sFjM/gpBCbMeR60v9aQUSsWx47lzvV8Elal7DHFzg
hIOPbt02FH1PC3R9bkviLbzWnh68GXvRklxX2IxP0zS11x9IKPynkuDtxHBnPOLV
dSUtcUcl0rkYw33LwZdY9+kx1eO9V6MtGDZl0JpqyIrYjXB0N34GsL10+dvIFTpS
t/EC9XlXMjrE7git7tU0P/yzeCdGqqC/y09mM366N+EAInOp6Vu+DKyUqX5L0r4L
jZRhkiJA3boFkYuWvSrugtIje8mlZO9nUkpfUpHeWpxMBTF7R00ZY6AQkPwM6V5Q
ELuBYU7hNUIJomCSscVCgnfpERFRpr4S+vOxawL+Ows=
`protect END_PROTECTED
