`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xp7glcMNNX4bOQw2SjeV0nUfAs0+b0FmZoEcjZfMyHXtJn1ZI7V1qE0K72Oo43h8
vfn/4Tm+RE5VE7iHiJv0WgQz3CYTdouUIyMYinEQvWErg85J/aZS0K2PdVEdtWBP
oPZA5wRuEywE+lOw5SjFZuLbdXahOaEEytmCQNhxGW/ZG6RzACfgasEnPELTH/aI
Y2zaKN3uIB1opwt6xQjsBPcwB5Zt+G6v1vDrlp73rFvMjyBkcUC334p8CShShML4
eJf1A8/acjaeEKXVOAk1wn8Oov9TRkWCOxXn5lFSbmOUghboqlnTwrJPoIp3ATpg
C1dKa+IIvKH16vR3eaBtBTVDjWzDGDq9gZzdqx2DpL/1hbMTCuecAE3MwvjureGs
7PzHwNf659/8uE5v4BxZsDgIsnT3hWrGpTfAxywl7xMIyXhvi3kK7e0SSIx4WsY3
iyg4DNPfUfntV614EGr0TcopDUTEwjstZ906UkNQM6vaWWY8YwEPbYoXm4I+wHG6
8U4ZsWVEJssgxT32haW8bFJxW10P1nlKE0uaY8Ojk4/0YMVdaVHIGvZayf/KNnkD
LtF8RRNaFl5GbYdiVE7fUA==
`protect END_PROTECTED
