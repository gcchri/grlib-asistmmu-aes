`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9U4W9b0PNB7g2/bC0DbuW4yvSlej2xg5Ewk6rGG7tV8XH6ldLy7dwh/sNTTu3WNt
bKOvhNk3Xbt/Hry7oEicWQ+jWD+AwvuFFj/jvKSqDAF52aO5xHbLPNEpEOOCK2uQ
lLOly2vSMMSvSwqHGzY7ylRV1j1essWb7ax/EfQaMKpIKXEqDceh3c0UnH4lDzrx
JVsec8MNnphmNu5D8gHAXHwRYQpubj880ydE/Vpiy2vj9gQSi7/Al4TpEFRa511L
WAKvvMGrejzmLXUKupJ3I/4P062BWj6w0j2iAMpQmNCPDpCQ8Ik9SgkcnidBGu5f
NzvBz0MD5wO2z3tmUjnNJbZyP375WN73uzCN66/j8kbNH8nvnDhBfSlC+J4MqTh3
itFx4R5hkap7ILuBaz1FXI5EJwZb6t6YNsp8pzYML+el1J+1psgLZcahsGwEJzhO
`protect END_PROTECTED
