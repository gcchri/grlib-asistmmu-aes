`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UJp7xw0iYjPA6HneXgtTdG82F1LmgBxDciP3Z2jMVH4jpDqCrb3qbv5B7bwAaHWv
ZlIR1mKrONReayUEVuagSN9p5KzUeCqLLiN2beV8OZiSEwvKHAYnevZmJfzbCuRA
TPIO/xZgh/fdpyJTrbLEDRxnS1NMl26/9krNUUt/aUKoaLx0C4VhSVPaeersRRug
Bo7wXr13xev3o0/YQpJAB/6BKsFTL+xg8rvFUdvaI57Ado83DVTEJwdlrr9THmK6
H8cYFhSp5jVX5TZDGO8HbcYYEn+xz4BiTNNJDcDVG6IOp8A6Foj9AiEfoiH381MQ
MStlZYhYOKFFKedLtQXyS7mwdJkl+uTBvFPE4nVSCn+ToxbsZRkkj4fKn3C1ETIx
sa9l8FwtHY4KTxh4gViW33Pil5KHaVkfi4rZJJ9g99s=
`protect END_PROTECTED
