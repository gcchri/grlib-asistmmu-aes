`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bcvJpS+4HiRPgwokYZzyp/Lzxe8B8G+qywbuwZ+hSzuDIF93YxNZOyKBk6Ru+y9l
fxlsWRp55rqTkNXE9YL6AGe7imo298u9uLUht2ClrrhkRqZFEIvJCoz0CFO/jmqR
zaqqZdoq8k3rjxHocBd3m37hb0zKDT3Pb3Gq43kpFdxsZPTdoNBBBQ0URgSni4nX
UqJlNsXO7XqlNgjSpaIVDomeydB44WPZsTq4Hsfng7HXED7FhPryqNpfsR89TEgV
CTL8GT3oRNeWFuimmuF2mb4cNJ/K5qxuNr4Q+vQEGfuE9VAVAdFaqw5LiTuEUiju
ZgAMqjhwbSi2eonRfRAD0EN1v8aeZlmi+Gl/Wp8uIimaKtINvUmbUoYWf8v5+0Sk
eD4nR3eFTSPM99UgV022fhgfD+G4lBXEhpFFK4B1iND32aI+dxP33TnRBzr0uUPl
batrZwy+oRKeYpz4C3FV8KiSssnttgbfMLrai6SdvUIkWmivTM+Mo++70qm3HMDc
tD+wZZeiVDYD6z4mV58Kqij19KWFlP90bDQp3T9QKNKR3vMPIV5yM/4kU/GC8FgN
qqHWRL7YyF91pACQ0WoN9IGgOpDEC+Rq5x8k4pwpOgT8Ok4siir6rHi7NCjgvrzA
EVvrFi06m3poJ6lqfupFw3oGO9KAAmtjvsP/vmbdwlo=
`protect END_PROTECTED
