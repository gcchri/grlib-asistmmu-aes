`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BwVeMLTCzdv9Nw7vBjCUK7nxPpRlWR+Z3BWPg35IF3Gm4qMZ81pOMNGdnGloH+rJ
PzaO1/LIvOh9jBNdDtb+9I7nQhc/PUG5Pt2n4Sf4t2f8aoo3KAafwaUPIWwGUXNl
qI09uFCj9bht61rAhS/619QoZHK/v9WWYGWUVr7nCMve8wG8IecvNaDCw4LDsSnK
7g6NEi4bsqf78CBRX+PRR2MGJKTz3O9HqG2+esc46SYrZsWDChippU/DyPXqLQ01
0baI0QeHRtSerrPNc7ac9GgpuNcwRPI0iaT9gs8T2IyxKrC67FYODVA+1aHmfW3i
ACaldH4c5rR0vJS5AG8fx1gf238CKWZr3rm6yI6KWhyJZiUQGZ/8ax2fNvR+N20i
UixuThgwUaoLvjEmYaUFJElSI/daaS/GQxRosLcNCFLH2r9/8AVsTqrArC8mLjuS
`protect END_PROTECTED
