`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K/QNw19YRqOrBbYxxnC63fhPuaatl4Ql6XYsf/nqkzk40VWtNtCocd5bqdlh/DHa
QI5TlyXkp7qKI//pONAj/Qjm1eI9ZrM6WCUkhiMHSABLeAB4HDHwnitLe8sVrhV8
pwa06b0J43Xdr8I7W/H5Q82Us/CTB2KFxIQl4H9WEX788rcHOqaF2WRh0DM5HXin
zrp4ZdKK/KMV/pXMcoTLCk6Y5YOobW/+o7flF3RZtSH6rl5a35d8dU+iilRn3C9j
/wZRD5RGVFm6AE9Lv0zxLw==
`protect END_PROTECTED
