`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E49Riz/LBTJdFPhdlNMUMfGKnRTMyaZIxiZFs2IoapfprsstKBMNkz97c1d0E+WZ
fgSqi2xuSxMkwMKwuYMrvGtCC09s9QzRfVqdGLLtZIlR8QDGEdlrSqfnYLYZ/H5J
VYrTIw6syrOfPpRN0JOGQvy+rSBZpQOwWiFO2CM5TJnPrepM90QW65DpEnCucJJ8
4voB8qCCPBDZcFVTLqVRYu1JlOsmzwClrc3PBS+qEnVEryiuUdYQ6oCVkJjV894P
2qGLt538vGTuZzxGjknIR2tOLImQR5tjCBhdKBLiu0gmIVEBeW6I6clFAq+QGTMk
tKtek66qG94P5ajy8P981r50NJlbPbheSk30VywQfnwaQT/7ABxEq7pHnuMolMMJ
MX96Yzu5CK0ojeesakXAFp2Jye0MlXylNTDg0okSAjeLVt/cS5h2Z6ea/77HaPYn
x3Y9Z6DSMaY5EjsLzbaGxKOBbMWhoAjiPWBcdb9VDKZetssJCCqEdIWvT59EfV3/
0HfDeNwiDLqr4ynJChc/MlBYsRf8O42iIGbMScxTFR3PikCu+KC68WW7ma3n7H4y
0o0uC23aaR9J3lJrXd+Xn5hEqnGsGtzqXvbq5FVSqAvvwabINNRuv6UDUDYigPvJ
YtMdkZWKyp4NRX3ECNjAwCR5J8/718YYXbl//IvNUXF9JQLDzLa90TKyW4/SyshR
5Q8cZSN1TTa+cjlixDx1GA45IMZZNeG5/Zfls7zxCqVp0jt5Pa7j3GjmPHQASSgo
Bdc9bsHqm8C+VQmZryJYYic6qfl/fEUeLPPPaPpiyQW55K9jh8h510Db6uWjY47o
OylQs7/dm33ykK8ZnFXdN4I4hKCbwgpml7WtT5CcCK1DEGTlAvMblSFBNf8Qzg0M
IuFoE2+dJK2EcB3I3QPYC6aauQhNsmYHe+YFNHSHewwou8pB+zv+S9IHT49fliBQ
Mpr6Mue+dTj3t4aUHEIGbQJ352+U05czkabgD/iZfvScJ7AwZ7J8KgTqdS6gDMRl
fwwCRfpJ0sNP9LMPGepOBIjNfNuL/BEkQv5qW7B2sc/ocP9vW5i0H/ShkJepqxfT
hEFWAaDkWPhdy2S3NYnf2UbHVRRv+N/gp0PUkB/YFmAgiNMVr29t1XNZgfoXxvUP
x2wWKvqS8lVO1cAof8dJ5WGL+KQrfaDZju+j/x4K3QczCBVqpWsPQ1cqiN5EpRn1
I9QNZr3bCdd6h/Bez1DzEHaXRWpRsBps7HNsUbKiVue/MDjpp0ndXmoOMHCapfJd
EknmoZ5JsHuf+kguzC3WoxiSDV9Jxs0+S7/ei1Op96ZbPKx+4PnL46pgGwsuwkgD
bsF32vUz8NKgR9ODsD+Tzuh1ty0S/6/Rk5jGCAjRtYQEllLA0PPpta3pYqVMn2gU
ookmJrgCpM7R/1wJxgcKEnm2vvi+un4QbUJ6aF/TGiH0p5lrKUeUMFewwXcUPvx7
KleW38lOkp/8fYWwVFgjzVJycqAD9qdCVSlLGgY8hAJ3DkDik6lkZC1NrYsSLIki
2iMf+CsM9GRIaSZhwsz9TAGTEOOC1tdWDWXExc8UNhZPGFLKOL0BsfRfHH18WBWe
8OyQCLUn7NAj/VvqMf52MXuYWE0vvyTQzINLySYp0twuv5uQPQ5IKEGImLJSWDW8
/Ni8mZc199uqZyimrDBBpJGrLlgbiInnTf5LewPHzaKC/jRn3V2YfONIWw+pcMbV
3kc8CDtlpGcvP9xSjNXR92magkRrXYH0viWOyUx9XXBbN2RQRPq3iD/4LpTcuF8/
2vlhRVSym/+J4MfEuVi9612pBwZToJsyvxANTknfVi8tkbUWIkg4KCzBGT2yMaoR
LST5EC5AVQ6EuTljawleO0UksOn26R1YC8CQE/KeNDNs4t+L39vIrn3q3pvlLvX+
R2z9td2vsF9A0AOB4FO7ZmMrvUREywuAKnKoGw+pvnR4eaJVAxiATMMD0RbrNJvR
ozNEjURzgehrNVbTBb2jZUU4eSkUmsPYbZ/VBtXN/B8Uo3+RAiqEoVh0IE/jCJV3
EjTEHkeRTpDKe/qb664ZU433bEo9kvQvQ1hSzIeQSVy7b4XtH9nI+2flWryoqWqG
hmrthN++CScvMAt+jB89Rl+ueujNRjikeaZ4wSkxpPR7rA703fjUI/ClMDGVnEtQ
5USZzq0feM21lYQ9WFZ82B0lysXFOEQ8QeotJfSjLPkz47Z9x13g0xR2LlX3rZFX
sV1D4vIhdzocoSF/u8K4QLa3+UJAq61OIln/2IsF24QruNtlGk6f4XUhfc4Qc9RR
vV1XGETx8dVbUfPFkop3tbsTsTJGGzRGVylbnxJJ8jhw1+SNsFHBbGt/9en7KIoJ
`protect END_PROTECTED
