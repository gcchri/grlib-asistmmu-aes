`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lCYjYY2bAHI84K73Vo4SdqqYmC5QGeYzyVT9pkNCkwlp1mwMmddRD+ytUj8DPBhu
YqoCtpx13uuZ8NB8FuTNtAh/Bzc9lpeuOfJBG8kgWhbQRjjrygZSRdpof4qJoe8I
rXzrSwMivDkVdQSJNxP7GjWOTxEcizuqHdxbNdjZgrzM/P5klLZGfpylF0iHLpzH
h544LLkXYSmYir/pKTnNz0NdsSiTPNW2JoAfcvZz/ttDhX/G4ZhWcf1D7+6YqNH8
tRG1GVMH5BIh8s+4gxPoqmt78/qdBMsdPob7kCB7DhvdEOI/TeSHimZ9lBHjB6Bv
c10lUJCSVR8q559gWTi9b3PQL0aXeeuHP2SS63I7SEVKrhEIIGX3YkmL1Ec/gT+W
pL4iDkXBEiX1lUDv/PovlEZoD8ENGXDLXVL628DlU5Od/MOyv1jw4+LxE5kdc/r9
zolOPS7cjYghvlX0Oetzh6c2a4DSgeDCEWjs1He7/voXTSYOkByrvrJv67njpi3j
S4hytArt6awwxJylwIC3P1O7G/1n1OE/XbxHLUB/UTVTVXatt2GOQssPCIjK+0fP
drlvMUWVrXOYy2EaoaVdPL5GAcQWjuO6nDwQAv0i9DAMdvqy21YTa1fMhZFLSxKF
D/JYSI25RyliiKbRiVOuAbcY9tADpiMTAYvfHf/VFJSAC2XWwD0sjRvTL1nF7Aaf
SsBaFOUJ2c53aMDA2fQ48SY6lik3ImprV5Q396MiXo/KCSwn6HaBRDeltCkRmpxx
6raG2RQZ3bz6g1jFt5Um+jwixFNPuj/CkZI1HTFJcxKPfWtwQZbUNF2RMGz/Rflx
mfvS65P8bAIwbd50+TJgSxqY9Vp1jCfjXCoFJ7O0o9FxppmeKOTqhs/2JiegE1HY
17WXKRJp/G9wvrAtJIGf7ciPp3FCVPLCwS5nfODydM93pKIeSnKWi37o1+8o/MMC
zoKWnk28gSFFOShfF32YT83FvdHdyuvwlt1Q7XTy9mM4d44cGvqlBP1B/gjj1zmy
g7EIOywfnDaqV/sg4iqtly63L+xBJHg1BpggiUPfbTs=
`protect END_PROTECTED
