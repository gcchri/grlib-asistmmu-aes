`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bMqNIGYh9dPqn7JlEoV4ZFIGQQ/zlcKejC1QJCMx/lpvJF6lOPFuPSyDwSJXbcdG
DLH5+Ivu6ihYFtngwMUBPcwhOgQrqpLwUMz1hBWJeqhV1sHf8fZGLsmT6nVQ9Vnz
4MG6HcgBZY6uHsa3VwU33MdnYwj1uXXqed/XW7WDtiOTWVGZV+Rspi4IVL4xrxQM
P555T0Dyu0gIH0mg+pBDARidyFy3Fc9yI70ZC0H7kwyadxpxFCAkhLK9hoq4FnYg
jsxegKa2K8gU9MnmaCAFa/na/7xhX7HMQ6QbOv7yr4E1wVLAOqyUV1xA9a9B4zFb
XTkl3BuPN+QNJAeIdKtmE8qAsqm5s6sKCeGScny/XEMqan28lqR+3pg6IKisrAnu
svTSW8RtFIGT2s7Mt6EQRqJ0BgL29dPDiVKJKQMYOq0vyyd0O2K57Iq26EQ1HYLC
JZ5nCpmPQGeE6jRqKpZ5gQ==
`protect END_PROTECTED
