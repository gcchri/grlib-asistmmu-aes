`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wn36AQLLdQeAOqWVaGhzedkA2Xvt7kUJG5wfiOO2zIILRHE0wY+LpSbvWjYWn9NF
QkR4vBfHAcZCRcLkSeFR4pa4vGU1ts8q8egHXXlzsacrtmOHy6D2iofAqev48ioM
RT87p8MCLFGo4kZhJjUGfqcZUpx8gG3jJ94RBxuBru4/Z4nDK1zWPzPRvB/bk1iv
E/ea1l5mfOluawEoLYqahAtAl7EFwC5ptU9uKl7bSPdtmLbqlGMqG/aJ0NmSr473
HCADgrqcG/d98NLck5KW9r+eAklG4MFBc7AAzVnwldhFRhLbJB3xui/tCmNSxf8V
v5Y0fyeo2WFW6/LDIkGxGE8FlxGOqhP0UK0tIJ/H99iqZsm2NQUJIgigsqwUw55c
TOCMTp6e9TymaDPOmr0AHfgbc78WvWm6hmsgvurcfBo2q8xhcvz5kVVC6RWBE4g/
xPv93i7mCW3M5zRZSYehnvRXXvA3s9JtD8L0p9SFiROTFXlozQTeZNZLe83eQ5mA
YSjKe+KGN/Y1+3+wGDX24fJJc/J5TVRvPuXSz27Vyl/3PFVHUMWiUqmqApa4Secn
Z9MBlhGxWjmOGx41rdM54rsOu04PID1lGWb9DCoXE8av5FmRPkkFWEtN34vuS8dr
U5QRsBL01SV+JkB3QdNzilsSLuE/MNBKmq/aH4w0r8VFnmaBpUJiRu+0+r6IiPPo
xyYoWicFPutP0CqhsmtyeTYLEFoBdDKB8ujefHRGTXA=
`protect END_PROTECTED
