`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aXO3VmxOlT4JKV4zgM2gnXDA5VXg+LYWtJUP9hbJL35PMGUIHFmHkv6J7VM9OXue
nglJ4lq9LTwxlmaRur68s7ZxR2HN08C1r5ON8MHkWMSCWH5UWsXk4JhwG22zNCko
M+Pe0N2PovgeYn9fGwQtgYta5CcCdiJuFsQHl/+4IwjmQdfpALwTnNNwKDpWinZT
Z7GkGZAkFIL+J/SEmlW19uIlb+hZlWKp2mnPOOW24l6W+Cpz2UDT9lin7NQ8kvpY
R35nLlyZTVz3FvZ69iUART7ERXJ5UO545D9XUgB0O9Pb/Tx4mIAsdE9JQ2HNhKNS
JHhN8ndjYfhmY0QpGG9qy1Z3JGSdAxX084oDqFz/PaPTEl94yR5doXGANANcnRsE
nYAkayeFdq6YeC9oMH5XPxCsJzTPRqGP4+1hNChkZQY=
`protect END_PROTECTED
