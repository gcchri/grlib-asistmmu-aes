`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JJhMQJ/f7o4Z4CnKGB428BIjGKUqo8Hl66jEo71t7z1iUlkiOCGqZ/9kehspdH4L
W1c+wn1q2vGQf2N7jzQVWM0zNk2NwRTbgF+eYJNcbxSiQ5zu2ZWGmLxcgqcoJHOd
tGHVDOr6kF6Op1nXpNi2Y1pRU9rSHhVhcyIqowBVca4XWdPjqdUmqI2Hfvo+cYFt
EstH/JEc+uMjwpYG54cGXzp0KGmRVeZg1X62mwDHHfaM9UZ3q4YBFsqcUE6jGs5r
LT3X0S2++w4v+MlTvj4Bli3WiVdarJd8JEq1VaFf2an7lHCOzzUKIrQ2LWcEI42o
dGVMTPcQTbMHkdkB7D1QcQ==
`protect END_PROTECTED
