`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ssejgHiUAGxMdWb2j2IBiovwhrFujWJVih8laHBZq3Fa1X1ZGnjlcblJmvYbs5au
LDsC0Fn76nnZpqquI7zYuiYqc/EJx7XMyZmdyeJjKM/kSDbKMR0DVfLKKRIlwX7T
L7Hd3zp334aGcffXM8Q2Wpuk/HgagpLjvC+IZniZOJjOTE2ESP75qIcszh784AHT
v9WsSxIbhQ18DXzCioKGGivntFksuGjHm+Gvnq/Hl0csekjXDe/NNKEGTw117LLi
foVM49Zu9jsQTlrxfOHrX9rDYpUzZj53EBWlYRFlEzvp3qZ4QPylgysvZzoisltI
++qcL3nqM9zmR+Cm6sYgF1P66icwznEK13pn4GqR6li4nFPcJlvfoUyeqZMlfywb
TiPYkrg7lDF0u7QVaW5u1o88cxCgINArlt2sjzfT9V4H863OIlBQN+l4TMs3mPHM
xmVuVt+zeczRCrGh2QNvt0nD/HwW3mzuSuY3dbKBfaU=
`protect END_PROTECTED
