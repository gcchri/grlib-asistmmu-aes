`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LUPCFgIV2l4Amyt5arMRquV02liw0fzXj5N3fq/aCQJ3Lgl5VUtbZQwDuPYoFFA9
O22QNqBGHUXeXPjwUFRxqTIFEYsVvYp+6TARr7R1SFP3hZF5Yc0HrzkvQggmaT3a
WSaWwDWylwKlDC+h8SOth+7hAh9RD5Q2n+MqA1Qmxey5k9bsM20eQ+ZvQClN1VeH
lHuacCwEoBpJL27AqXqGP96nFSvV/hMhhsfINzKyQgkU/2tWwo3WU9+2GAwTWgMt
xT4d28wXIgM2vtn3pd6Snw8/BWC7/5g6BZr5zHxwgcE+7tqPjf5VOyEgRdx8s7/C
Bx42uds5z/uhLVu3uVBKtqw9Uw4HuALE/rk2ppmboDq1BnHjyIJw1H50Rk5Jrj+r
Itig28esGuLQw3g5G/L7tIer6RVRkvLQmTwaFStUVQe8pcnBH/ZQ/XYA4PF/GsXl
Fld4mQ2fgk7WdPtdNfFElkFO8Gv4RC63Kxk+bESeB5SBw6Gu38GMtCEHM91Mocrx
n51OSpODN3SOZC53/hHvoO635Sh+Ll82AS9etOR/C9MTp3RTkF95d6nYcwEBxzBG
f9by1GDMVAzCKdFuNUhcITaRua6c1qaKPsSEsvW9lRdn/pDsTD0gJzVstbMIDgbq
XYDQW9oP/a2KFqW6QD53H8WSHrO5I9Rc9PcyRddYcl6RkGoJY9e6W1BUZJVtlUKb
LeqXpQN9mlzL1tO73PjH/oYO0YkQzXJ1yae4/EppYvlfwPU2MT5srZ3l4mSGWiBY
/wfqg1wP60cQtu1OX1drClKaE9LOqw6+lS2s8b1hROc=
`protect END_PROTECTED
