`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CCaoIFCG2b1NLra2/aPKULxSH56M3Eck0WXKH7N8qjgf/XEbzkRMFlnrNr7aHauh
RohS7OATf761rpZTWja33JRjK1A02AGvxB7+jINzCscdsGxrX2u+QOgwLWAYUwWL
L5DVJuIwcROzVh4Szm8CQr2LNVtK8C1lG9y5fORB1bcQZf2JarIQig/0GpFU1I5L
VJel2YZ+4SFnRpI8lRWS1PVM6tYqG5B46XvFW+3T9qyGyUy+fcfSzxqadbPXTzhS
P0fgxWoEvw9o2LC+SSEn8L74q9RZQNlm4K03F4VB6Oxg5rfJ5ogFO1HQtJ5WdNEb
3JFNuwU0gAMCZDzbsNtrXpk5pzZS/SJqbZ82sXTD0f/0e/ndMcNNTZ2/KW43NkSj
rj4/UgrrYp4CQgwVfOD6evZLLJVzev3BI6RXHRTIya6d2MX3WO3mmu5OALh+FYPG
qnNWNabcby0CO6/W3l3MwhXmPiZuMFuvfy5WZ9kuPZHyEXHLNJgtoii7c0qopcr3
q+q3eIOBGErzKGnDxsapr8jitydTwhHgYi8C+aWmK7l8cgGeRNwlKpjzzcxbsN42
7yUzggKI7mfu3zfvtSjEk1Ampb8gjo83Y3d0Tk0VoK01kmREHCQXi/fXY5ZENMT1
rmugshfBq5Hx2pFTLMuWnEEiELE6Y29sFDbqKweDFcPndX4pr7BsFaoL6tOmfl7S
ySk7iYGp4pwjbUeAEpNgb6Gx9IYL2ReDNWdFYFtxnuDzsos78s+CzpC8BqeHPfjo
K1MN9TqNtHfkaCXCoUgr9b3eTe5pIBDYzE7gp9tvF2ixHoZ+a37KZ7swx+QrpjXi
9dl9SpKiLp6+MAOlcCZ1HFZIPWw5UEpk4cbEriL9Er+WGcyu47ysDTGdm7t/O0+Q
PadwfeirxYams5XrdYDxjQ==
`protect END_PROTECTED
