`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f9rJGqL/OYuFogVHhSzWLp5JWsz8maFe5G5RlD+oEeTIkZq2tOhdLK1mxoblmaOf
3imnnBZyYrePKyrUiIgr2FNVq1gCBNWoGZl/BY3BCGjEJfuHAotJu5gZr6b+mUgu
QBkiDrSsna5+UbAPVEhf08HJb1H7yW5cE0Ixo4nroDo13QV6P8b6s9SGbz8inRGr
sGi3Ma/GIIkogIvhLkZUQFh/g63jo24EnpHg3sBdVpkGcVkhiavEC206s1kz+nSs
//4Y5SyzwD3q6wtX0dV8pV/LufpGmvWTl1DFPMUKYFBR7UARZ3g55ZBr8YxxXx3Y
ZOu7NyhMqhQpU93tSvA3ETW5yoj5UxzyeweXDXM48GlqMrCLv0yYeqhlSR2nU9D1
zlWgDQ/s9lfRbr3SVkskbfcjJgYQ/qHL2ucAD8lilLlhh8Jby1JLAAprxvtyObiZ
3O72p4WZjwUkZhBGM9G3zZ4R4+7wA0MNujnnXpsNXnuSLvp6Yg7HNoX6ixRvEHVe
lLCktzoBfz0X6h+cf3E0ZTUeVynfSam+FxvIsjGKpy6DtgFiX65ob/hNb38QeTAE
nNuSWVYO+5lg7KgcHQGQrSuoaCrHxmrXtqzR3PZFQWyqSEn90g6UzRfjpIgblAty
O+HJO9erzaP1WYsPeAVTOmCKMDRzVtG86S6IhGSww/YXLX8xg4ql0MF8oMpu40ro
U7YrHha0OCXh1PAWP2rcROFfUox1snj2PxZEBrOF5uZuemXul382li31AfwyZHcL
h7CB/nbTq8ocOTZOpKgo42fnWiMuyHUMdm2zXxACCUgsRhKh9DNa4CWRNYUYuegw
4WEIgO0PVplaSpfo/fjDK6/lqUblLOVvGK/jfM/S1giOREiyW9FS8bn1heU3wSnv
+fzCzd9Mx+n0Hx6+XLNiYOJ2ch7/4cIivSUaQVuuLkkV/Sgpc4qW4/GXAb3sxouR
`protect END_PROTECTED
