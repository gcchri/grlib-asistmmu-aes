`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v1+AS2yTOo95gwF9gkhzM7zHscpdh53UPvKeXF5W83432bygdHGrmVuoFegnPVOh
X0KguwBKxUD9YER59vxEXvj05qC4Ac+DW+ndf/+JjA1ysxYA5Q+gI5w06pyVY/wI
wUTSpGORL0ccV1+gUJNFPkmfzYb5LZ14PL/8W5ntFVZlDT8+4SEJodE4Zu3FM7ql
aNY/dFjkGbb5JPOhKltrqMubF8NHUWjEwzMlN22QL3xLwx/EAXuzeirXu9KONmT1
`protect END_PROTECTED
