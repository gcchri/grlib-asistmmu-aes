`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sfexTXhjIiJfUD0uXeeAefZI07htkacmxg5CHJeiAUSa5E+lowoU6ExkT1kteV3C
kuWfjdqLF3E+JulrKNa71CGCmONIQTIAwOYIustsHzzVSLtRAKZKn25fBaqWUAAh
zaHfqbE/OyIYrulAz7SzWNZ9hM2HJ8gc1zUtXL7fxbbrZvTaGMjl8L/rRTaHrMAg
mt74HEoEixP/RJ0AuTvppQb0HuL2zZW5NEuESnc8rHWWmf3syiAbmWTL/PjuyAmf
pmPh9v7kL6Pu0hrPKNKOBhXW5BCWIyCUXCmxpN9GZzNPpHndwb1gNwQL7kKi7eD0
sz//HIdabyzbUA3uiEXUmXi+x6Jxw2H/cWdrQ/3+qnaDFgnvfcElMzjoCXqJBesU
3AIg0G7l3n2CEMA36eEiwYv2NL5o6QF9PYeBe4CjvhVXJzcBv7YC9wviTlCqb9zz
h+LlAyAn3Hf6t7Adh6q/bFFC8MwI1ddzawz9UZkG5MjLCdc37vYOxjIFLVH4I0+J
Nmj0zWWkSjz2iOKkC0sIh4+coIhGCFGNXZvAifOrJh5zz5WBYN4ar8x54MkYv3Zn
Wt0XiDkaLrrpWG0r1/faf6gN+XMIcRRFRnBsLsGY3TlNJa3XQRuSRToNyYHEd2wt
9GwxWeTKCjzys6yhhaFzo4mBvUDRHyMMcg5p7PckGpVMHPArjhz4bUrY0854bx4d
28Bdrg0C+1r6fbcpxNvyYjXJXjqJ0/HswgssKj4/bplmyelBwgltDQJJMIOqCIHD
MCAIxwlxf4bpEvl3xg2oCoWuJKf1Aj23wWbyr6qSCk4/eSbO3cDsF+OSBldsJvPf
T2x3GuokhxZV3SHM91EXDbNMjQbujMMozWdPYGV1g7U4KOCzx2g1eZ9FdVxclyYf
H0xChoYZQ+Z2ssfPlmc365INU6+jxqs3/pwGrU+3Nv6QK6BY2ikymuQoQXKwnqMu
v4ER60IHGazhXPwAuFeZgZlrky8wEuu09gGu9OkkjPJczNLG/Dsz1SCqQLo32Jjo
MxnWi4a4WkSxYJxUqSQLbZ3eGK7/cHPPaOoEzY3QaxN428ilIRi6H/thfx5quNLy
zELOQY/GwhzhW147AhXCO7/+m3n4vMtINXT3YEMhAcJmaBpRRTjwyJ/F7dnM0rYX
DeKCrWCyBsj2XaSM4zGAX3X6SnqmRu87ACwBW3AvxWEUhluq1FBOxcnna9vp67/H
2GogTlpp5bsEto5cUhaqGruXPdFR7Ul0b59lDI9HlW5vRe530lzW1TLwT1er5XRO
JT67eTXQgGyljY8oDEQhGa6JHB1NTxUspq1IhSYIKB/2r0vfKDjaLN44/U0OQmzZ
IoO29J/lxSCaBTkbf6l06dqzX5uitDulTVEwTegyrBRtzjQQv4jCnweigmtAWIbu
3kIoYcZ88ijO6T+QW6fIze2KmcYpUvzwdFH4Xj2zFNFFLs5nj6qALwKi9NyN2EX/
7blbuOh0enHMGBdaItV8apx6iavtLtEV7C15rZ1zJAwls7KeKVkzFpo/PnArUonc
2jOO584QPmndFC/Lv2mGsmr1aSfCtOMcsv/knvkt4ZXfTjdP/V602mdZOz5liyKS
TsdBc8Cm8pqr/tjGgfIwn4u50aYO6OYw/ErLNAqyzSemzSlmECuyGxvqtbKzGV4b
lG9CSEyRZXXPSqDc0F7Pt+VanD330ZrYxaESrQLEPUKce6G4lfLlMo1hp9FuMgpB
hS3OJOaTSfJBfxs11IEVyAGIbveplKQlgAaKU9seEO64kLSRnDfLjR8EkDOPVwZj
J3Aqdv2bdjYG5O9NwwVkwHTpOVTDtzsGs2dxECHk8Ehu4l1V7r92mbV7OuAbeHzl
77Wt3IKKiphOBkNbNDpPfgmCUJJz0VKMW5BsEobtzelBCuhMxSyeOUOtw08l3YRc
JpkcNh/nb8GDppztbTwcc66sx9SRwnyK3wxuz/w2EPo1IDHc6S2FIaCkLhxw0NOm
1yQ3BqaVEFPBm/Jzj5m5YsbMCv50W+U9cIktVBuljr2iEoJigBAUAPOINYRgrjUX
awDp9GURtFe0EutSkLjFJArsOKpU4voqaxAhDuw2kWh+wAmkTm2ne+YxMfL1cSHv
tWRQBXHM/7aK5ukIU74dqUZnO8/JfOGBDhI7VOWSaNEuJjmpxCzTnl5sWMd7t8k3
/nvS/YHKKTsSgzyN8rRYKYeiQTEmu7xkfkzLAZPVQ0cEtfbnc92zBPf383gmOtpt
LcvLMa32WxnUJrp21bkqYa10+/dO9XzaxpKK/FDAhCM+nxnyvoaU6aDCpt3EQS9+
RSEesDHDK9Ktuoh7o7EpQnFG1hbrxITueajsFQ/OhTQm4j/ntpV1jkzA4W69e0XX
nu5Yi8wjse/MCDMmV4RwgBYl+4XMTuUy0gfFCSIXCaNZzrysXV+WCGPRt5ciWZt9
FQcMuiqZjHCeDLNRjksxNizDGx930KJxAoRTXfCvCDxVJiSkPSf00gFTDdSD+rUf
4LG3LwsEEeNh1pcx0caJOWVMmGo7RMOTp1ohXZXQmuMBXkzEF1kKiSFos5UXwaXJ
hc6+v73nC9KpLzjvtV74fOXJaRWwD7CgdzcwbL5yCGcHHWgW+F1a+u9ZF5+wPezy
ZD2Xc+nDXtUPqBRGTANpK7DIWtOH5XK8VW87I8NiudOXjABx42zhRZtJX1TGln9Z
iPIM98YBA3fqvtgGr3XYZKHB7sjSqmaiXr1zKV4R3jTRmRFmI7NCm/SsRTCgH/HV
usrQSEshrk3d+93xQay1LFufUqaZAPoBNLewQc0FZ6xSUbC7edQehHhLfweiqt8C
iQVAnbThVIJ6J5oz6dPKs/mHx1YZmOvf9kBXEWeRvsm/4sHb8XP/uSsGC6Dqyfht
gaHYqzVqtoZHnGNv3u9GUqiiofDO349xbKljtilkflflOSSjIfeDetp0AJ8BdtAw
MvPt+S+4aYdfuRGuoMPI72D1CQc2t6qps44UnQ+7Nv6tw5doMsOwwCJVwRlkEb+8
nQloUNP0g1YqudG4V0yjloKHht1jlHZ3WSG3KAussCC4/cPeQHg23ZfrFZL9XalI
o9LEkGJ27c99fhYBbWt6vFgoSCb8RfwXvKcrk/MTkG/moNMuBu4JmAYPbQJCyXxG
QzL6dLk4YrxUJ9x1KM/P8uftORog6zoYuLfQqjCDoe6Zggt9NcewFqqexJk0Yzxq
bdm6s4ERI6pvtst01xpyx+UwcmHjoplvH3GlCdU1nGVm7CKdBdBcQzIkbsrXbnnS
PJ9FzBc+A61BG9fdeGTd8VvI7x5RnuGGutqRlEFxHtDkHan1yMubrpKmnCtYjoo/
nnFWr6pUwPb9jHH6cLs7FHBA925QYtwofzoLB1JJZkjJ6kYi4sWOra/nna5IcNg5
PO0zfjrO6dBhlSg6KJlNDmxODLBANn/1QBRiXjjfjYkcVaSBAiI8SC0hNpWWZPV4
GX2ZGOPUhAfKQ963Ng2vfJ4wkGNbG1DfJHhr1qh8FU5cYC/OfGhBSKoCAdUwP+19
sQe6ouz2WfTfMU+UTIeLxSr6mIm1tLCXcN1tHkFgxgyHlg5zmg+J/ShVr8DPXUe5
GRjkKfhQLgaZMgS1a+HzeyE4T6HvkATOu5xZTVqDdJBLg9IglpPmMWXWwdNvZ3BG
sMKbynfET+Ra5N0VSOqh5ZDTIgMsUfdPnMmyWlrsgll4atninf0GOMQj83RmMlkX
drF6e50eS/mCMYNLMwlbyPbFmQrjU1/sFGVcieQCpxHXegJnEzP5LpeIMEq0J1cS
VyfLhFNPbJNq6zBO96RJyFLEWstC+E/rEn8zOuuksz4Gh62pD4D70djpaTvobMm7
1RuH/Q0L6jgU0cAW/uaOCRfb+T6jDJLfswzGaDc4473WYVRgX0heAmYYo9VENjmL
PDNusnoZAU8rh9ZpR7gaQNtGA3Jwx6FH7U9+kXlcBaKHSMkznNWSZkFYeZoNGfgj
yQ0nyghlJ5acgcj4JremuRSrdyWGYbNXbbOEqjgezRBN5fpaYdyRPEiNwV9/2GBi
l6/Sn9Cn3RsPeJX4c2kQZ1czNoc3N0iRAXlnn5tCpCpQR4JiASjQdY+sLsM48dNh
hcTlKlEtfouuYq8jkBzqQeuXA3ZK69Wt1g1ndWuiX8y0RZ2njjUkWU+JE1/Uyo09
VyKqmAtxzm1mDOwJxUOWdyMgLJjNyQAC3PqAbYQbfr69SpVekDe3kdaQ2/S2uklI
didErg9X/wgTItQR3Jdr1zxiEtxc7muNve4ByuE0pvGUpfmE9Vw2U1Us57wxhU/C
S6HwBRfaSbqs8AmcmynSDKWks8tBmKRjzm6+lni3IJOwQzv+DkNc3wHPQEufqQTz
RNSUabNcpUonwJd8N12lIhGWtUaA06MrTmt8d+muFetwPKNlTv3nOWkNe6kVLC1i
IUJY9RK1kVDHZ8CarCol82ourKPux6t21tuMs/9wfsQ=
`protect END_PROTECTED
