`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gB/qavyE45elyXQJB+NqQohedoc4WhPljIDVN94lX2Z9CGEeBI1LQ7kRtzcaF9+j
hPr/oVp6U195YZmVT/q2RhVMXsMZAjBs6Z6JZw1K74vXRvd+zK55FgYXfn09ZN4h
IgXjfH7mUqeeR3b4ihq7XivLRspADuV0le9ge/h53hQndoT3LVNQl6r2+iIHzqbL
qZIewHlkr86hzxC7NqnBSJu+Si4QClbQcNd8R7LwlUr/9icBLSyFCovTRUiwG+R7
qpvhHNElQf5W7c91JHyHexQxDDtlgw9FDJCp1eTupfSPDzrYG0oaVtHk5vK/P8dC
QfobVXa4kbyJbV7rabTMNE5skJnRUR9VQIVP7WDpBmzUMoWPSTpUh6IgZhPoqYp8
zaRxvLGC11kZHxDNHdwHYXF78xUlsqQmcOYQCVZy79YiGhkzAMMLeKZ+yUBqFXcB
8T9j72FKhPfMDiYQ0xZc+qUvFfEHWZ2653a47KOy6lJ1u136NEmJzmo7kN8tK4wP
xnFSnWBeubCmZXJN+QfiTaKj4oZr1Hbifab/2Go+yyUmCjtVWg2nZXPDaDFufDsI
i3/0Xmv74cVEsn8/01maMWBbIgFx6oSpiD9ryeFcNzo=
`protect END_PROTECTED
