`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zjBFiHH3PCi5qD9u+Nphrt7obw2ORAynu9Iyt/oY2OQ92IcDjpslh4u/sRnx6r1n
72WsQUjgR6N65zksXXT4A/gUgTcUQQFaeGMsu5eRtnGxhDTk6dAXUs9ahELYYVQ5
+Pvf6wRzBVOQ7Dttm8m7v7tXNgr7mkghTHTG8l7vuOQcwl5wypCrL6zjhBNPOocZ
wNq5zjnbtZD8wOAqrvDrvu05hyBgf5qM7Rns3TEKmSNVD1ZN8wCdIDkV91QbrPHL
32BdqgzBJn4Iwev/9dzQc1q10dFb43ovvF8MtwrJJ6RyRxgX8mYLhfQdj3EvPth6
LEQ6onle11O96f8TXmOAYKfmVCvBdK0gm6DJkUQ7CuTpKFcyvWx6IqSY9JfGnIKt
mV7SSq/W823vYD0zem0ke6cM+zFK0riYHtvYhW+Ph/xrCKA2pYWVOoaB+rJIJxAt
fhTdb/ITVATTv20ZSRVyAlZpnt9OpnnM+y1JGpe0hbwrFKSuqzfMzGNEmqt1xLQT
56UXrFC1af/jhRkaSsB0j7JQnFOZbG3oe8BMn2kT2Llb0rae336HIWAayL3Zo6O8
uXNrZdG0xwxGfOvs6h8pjZhB/xONAyIPICIeKYW4etcw8gTvaLEFSIJescK9hfId
VChCE6NZKI9hqdVArFChVyApudm5x5NLh2ezAUNmnDiTe8/TvPMGSBdpXhPJY6Ul
Zi1M7tmvxNMXZorf/JY5AEaX47Sta/3paK5ggYLG3GqmqxQkpnhiv/GTEQAPKwzH
B92wSb1/2RjBSCCOWTP7Y0RViuJN3BJ7KKBLDARcxqLhmePNQIwaPCmF7xUUFEqA
aoeGzwZqIpde3XDrmEXkodpJK1yXPqCMSOEHK9H/cBE8K++tAPKOm5nLeC81H4Vh
EARnlXe4tn0i8lBkTVD6XVpVGQpdLokGHy5Yr0PGBQXm9GlmSJ9hlIcvGuYuGUj8
`protect END_PROTECTED
