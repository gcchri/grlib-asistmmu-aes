`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2VZMY/nD9e0EjWMr1tZzAXkObmXKqRAxnznqr9iNQmxCXTnvuDYelCXkYCO4flwo
PCA6oQ+SE7zPRLHW4teQkYyDVJOnj/JlRA1QOURxDUF6rqZjsRtQDWq5vC7JwO0b
vSZ8GFJQsK/57GUjjMZdZqb6MmELiHDcRrNL9thsomaV+kZs7pUankdTIz+1CqrV
7iv/1JbvcFBrPIZuDvkcXwRszm4BETXRP1NjBPnh5wWXFdcGtYvb13rCTUtrqLHx
RnUYFqIkVbnv4xW6AuY7whQ4s5t8qR0L/66Lf+ErzLuKJ/oZfAiYwhN9NvESiU74
UezhK1yqR/87U1UUSTnlIQ==
`protect END_PROTECTED
