`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gEkYAQ4LC3XcP6ZxnE6IWi7g+2/o+7fSUwvTlbtlBxsJu70fLSyBJK+5dSisgLtZ
26cW4MuG2PpdEbnMG8+BhH/6QJBOiiI5GS98JdM2KLsl5AwtgLYGc/2UConu1ppg
dMfLCFIzSxBCUkgzB2JTl+GdR7KJsyOUBDyrKlCUvP721HVCfF9jmElcJm2ejxLg
oZLU3UU7k9ruTuNozfZ3bJA2bvGH2+gksTC4bxt2swq6nXdTE5DnxE2ptUa+DwiW
rl8goqNctnM4tMtfkS/ifVJbCrE3Bly874aWjkRSf8XAW2Lluh9Y3dRt0wlgb84N
88XbXfvPwkZ4d3akyxD36O3TIv3EZQpILG4Cxe47tFfyUfDOdEnABjXLwiid/Flp
FURLtzB/6Y2SY1Jr201DMy4WF4ueXNreZ2R+0TG8aI83RwYVHUbk7LrDhDm9RUe2
V6qZoROBrPEB0GkM9EyGh2KrOxtgnqHMDuhNvXjdLoKaOAlLvZrDzvyUJDzS5wP6
P+QLhtML0wNPrQip/6tq5sfoG8nOaYpnUHQHA046a5HaTcklg0ArJb0QUeqlDGti
u+CoFM8SeY/7416ns5p3Nr1SWHWBvmnO6m9Kvmq7CVpOUD39YFinT0e1zrmvEwVx
yUOzzHtyak9Vgr2p2EoKEw==
`protect END_PROTECTED
