`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u35t20sikSl1FkdJwCknI3CHhpA+32NexeflWXt/Iqfy+YQVRoMfELXBq5+TZ8Lz
+7KReZ9+qtTt/q3TXetEcmR/D2IHY+9CHMGCjjSALtxelQTul/UL3ITqKGDi5Zs1
lr/5lFKiFqoDeRyzV/tQcnlrEPAXCsnf7jIVnmvENBvG5LhuPb4fwWiETJ2PpaGI
MSdrj9YXSDyy/721Vun1BVwaGHJpMmx0HEA0+w+FBAimvUwsPHBBtgh2vJxZadJy
GKyKrnIjsMmPwHDNejgqrO6+nxFKyu0OA6FE0fUwpGAyiMmiCfiMkHcS5ooh3FbX
4re2QiWNOIu5T5rtFyHzhhdwC77Y5Qc9AUYP5FcRvCWmBkYG+Y6wy66TaYfBkmo8
zrQTJyZV9H38729SAg3+7srksjAw0QNxAxcTetUd8rVYsi/odBnYG7WDC0gJX736
HquOVwFnqqUWJ7yKrd9oatIoC0/kBUBUNW5tS14C7OKKOoM82mny9znfxm9MSsiI
ZDeSa+KXhaFAp39PCC1yGeu8OBSpIsY8uzK1YObty03VnFi9uC6JWHfsoiyr05Pc
LenlW/rkwZph0qaAl9cqrR5m7G/yLl9VEpVro3WCkTZ8aDg9f9Pdey5p+TPGXjtz
maNJVebSqxoCFOrS69XFP+ZU1rOnAGBwJXgElDS+JO5RB8CtEeiZLQItqrIHXeAm
6y48dgZ4SCeA/cBf1K67WpB42sxvaAJmbIXBXE0u8U2T4e0PTWyYuPs8kJTvwZSb
6V48D4+bC98wRwg6n0ih2GO/3RH/AQuyUafL18JadLL7ZAR76J3BgKTV17ZdF81z
Rd33de9rFbv2kbLhdxXtK/8Wl12aqGyx7t093+qriyYx+9ZwppXmLvgPuDncXfFG
o7SOcQeK2hJ6wjcFlM7/u0T9UrqZWrwQNlxG4/Bwqtt+Ud2rLqtdit25NMGlzZdG
VtgQojA3ZojjyHLYovLmE3+xezeIDMGFtezi3S/VrjYg/R7LEaY7iZE4Ru5vO9Xy
lg/A/0U1+LLEOxJUTLfQnBXkkYDYb27E0HrbTtQxKu+tHy0OQOnaXLxL8turPh5K
MMq+kKbHry91yW2Y0PrxOKqQRuQXFShGF0VsoqYziEpw+uDBJj/zpdzcudVPGadu
o4J2qolGZgIOAKMY5KFJJatQtEiFwNg4QTxskZW7Wc68pqEM2VABXSgodbSI+5CZ
6N01cewKEoOuBhIIxQzDqmtzuQAcxAMLJjnoSSS/aGYcmbwsZDMy67gj6eTjjpqJ
IeRPaNp/Zkg6RWMhRBn97DkRnbpqPdkdjmFfScTH7El8VlZEn0WAzS8TL9MchvwE
L6ngiY6DVlL55MnA8k2lXKFrbB91qfo3Ko6yB7GVtn55U5HJNgKZZuHjjKLqLMHT
UDz35tP0rMfugVIsCwgtv1s7adjDYlU+JpN4QOuZXCea1YfgUMZYaeTj94sJ7xvg
tIaXi65KcNL7hB9ovqOwWM8aerNb/EDU0xHgio32aSXMCKB8uO/VZMTwT6oRu5t1
wwOAJO5Vc4jipJhjdkQqBHG2DkLMwzCuCkUWjL+fcfMs0ARZ7vCzmzxEo2gGS4f5
L22Fvy1XfWVwp+r351KsKEGFD0vd/9UT0hCRzemHZUfCzw1ntRIxY7sult+dMAxN
HB4khq+RhxsYdOrDvkKiFTNMAWUbkGg9JhH/VpXpYQjFZw/HFLQD2Jp3leUNY6wj
VtiN74A6CbvrFvnlFH4hUj1NzIN2ZRkr5si0XhtnhILfxbDvKOF3Mv4kKUm7oXsy
AyOIZhoEtD41ajUbChiQ3828qmS+bNMtIdmrtAf6Wfhq0IOCEYnjfqRrMOGBmgeq
X6VLeUEUZo1Ef7AjA7WI0lNnw/4kvFOLjPR4UA73pdbCW0SnUrSxii7UtxXYZZwX
9t503CjzuhG0NIwS3lGtnW1JJt2HJHUeUmLr0wcXmREggp89KUPuR/dq8Xwr3BhQ
/hk0jVBasUjLoMukKskAVA+LygTXaPCshiDyko3rtNSm0wquZ+1aGSQcV/A1Xjqx
mBn1W9VjOs1GpkWhJ01GiCmADG/6aIOgWkkOjoFeokpKAUj7os5YHSIsSz7k7j22
rCYgsQWepsNUmuQoxrGGXMp0sgnlbRfYueecR6/ZNm5p0ikrS8a1EtxVe0gmZjJ5
e9S61WuBkjRdHPf8EbfU+c6/Vtux0Qjuvur4xTM3l9yVzY7K3sHsSyh8L1TnTozx
pRozFSB47moWSRkoN4pXb3jVATfdPB909almjNw65MsI/x63lQmVM43QPwRTPu/l
1vKCnL3mlSSorkbVBCwXbCo/gWJic9HNMfbEKcvexvXJIttN5hPNJry4kw4g4S8W
DSLzFVTomwF+kYhGVukyldhPmVT3ReMPkWCcROs6MA+flS0Dauef+FdPO++QNxah
YR+dsSMlNe+V70oz+LU0JqZvBnfcKerYMJjELgcAJRHd59nCQsbG8G8RATZWv7w3
QpDiBeD5LpG9On7wX2Po3dCRF7YPAchLVnJCUdCsK7MCppm4JU/uGdSixFnFly6B
/0CQRzn0JQ1ztjU5/SfHW6xcBa0OmIUKRVGRCUWxdoxcVejqywCH4c9JNuI3iiwv
wSolnY9zHG+FbBmexnfgJ5VE//5d1yP0HJyM9aHjibT5qtdE0J0VMCEzMWgvdD78
sZb1rQPWQyK8lyUs5vWjJeiv7vUOyieqBCXq0Y3FOX7AjVE8DbmQC04GrBnHYTKJ
IM4S25Fgw68lsRlRHwWJToyt0/hR9U0MnC583DQT3gS+9Fg2+sOxzRqb0N5g8E4n
c36pt5jiA/g1wLa/UJkaBQ94McxERWcW6sZ877ii45ZAbEVsQXg9Ce3La4OrLb1K
8RP8aP4j4TYLixuSBjsIi1ksSHYSYtNesALk6jm6URAd+zYe/S5BYTA5lbfBnA4t
xp4uEDSbnOw8wDvqu2LAKe7TX7wRhsAcgV6IjRztxlDrhc5DBCQHSekeOGkX/mbh
GisPSAFwlDhtF0ovPJkcoU/Ns1jU0ZjnC7iF8Nc8f4execAL8p/LLffTwqKa61Lg
jBKKC4uND6c1IVy05ECXL5ULVpKwKWVBw90RZVdmA0wvBxKmbpWPuIuUpC1p2x4H
wUx7uno8eu6DDdLoWHZWnN13isidKAc3Moli3R3cnwykUVZry2WyYaXMg8oRq5z9
5YVPkPFophnyfJDFf9a4wVF7TBq8iCyROfxm6u0Z7x9pYuRSVG48VoJENZl/fI1X
5PE3CdLOE4sXBuzoeYyZDbvLSWjWfEjBAsne0Gjb5g5djWlJeS5i5WLUMBxDDYTs
cPxZKtxqcs5y6GhgURmTU41vWPbkEq2/axueBpiWR4jC+X1ThN8IAMQ7B6L4FEMh
htYh8HFH1RDJDUKFArR9FKoPLDQ26u3euMkVuuwh2Z+fOkRz4gMcM18Oe3l1wzdC
BAqwdu2ShHrGxWcxxyJX7DebjXxB4PXQyEm/2HSzSW0q/NXCaXugT/NT23eV3obw
rHb4IyAol7lHvKQEiM7YFkbfudDpBh8S3RNqRoHCX8dhrSIZ3U6FjnvkQCJMU+Us
e94/TBIA+Cy//WIb8JGtYrJCBNzEYGzTgIJ54SI1eWAf9qFageM1VtOrjVoqgeDD
ZLwaTMxGQnjwpUdfDuetJ6omYKirh+KqZVliFfyKRQaUALWJ6iWcdFOlEQspcrjQ
zfHcSsSUVJHKMYxgi+bGlwjEl+ulh27lMWFbjpubGknGE8NDDA4L9u4rcFEv3DS4
fIRMQz4zfy6OVPYSuuUCrfcU2n0NsmMwWaFtSXDzZTndy5nhzl8js3p683D3SPjR
76TuPJrFQAID04rEXHbTdpD87QIy691ZgEFtpSGdcyBItz9czewPvpAN9NXq/ci5
qBxds/xMDS42gyF6ggZjQRdCXbXdvxcA9YWWQvu/Eul8/nyCH9ro1fwUhzGfVLqs
h5CRXCI5ftSu4YMokGRANZ7EQnPLEUyedfn3NJHW99YiVT4yAIiOKZYBQdu1phQj
RWdvu94U+hRjIJQrt8QsSQUwBH+Fks7DMmudjXfOfYdKBO1l9Ogb8n7z02Z9H1U7
KnEte4tCzwZzW/7kG0fC8HSicNBMTzmuLcGqwxnLGJ3dUPinKn8ZPrhsBofyjgws
NiwBSKS+6hPytSnTXBVQxMlWemfeliyAsIi9MkHVh+8ROSjGDYDB+HiEai1C+f6Y
K3GK+osR2yvufxWftfhOqaPdbbLmHd1d+yvSOgbUKX9q52pvvA3KsRqwkl8ecZKA
+U84GYOHctNaLDxXRozii+25kWuCEu9A7TXu9KmBouLCHnuG+DL4ujqyynsOpLxB
FKobcTNuZClZw2SJA8fzad4MRplcwSrHn3MLTUIjzUZKBhG2UUT3KLQLDbJPTLdb
ByhL7+Jo9nduKOGqI8dYsnVzKoXZkC728Y9FglnC+2I/bQ2YgtrD2bq+x6jUSbKH
f6RMWnwfJ/6qxxHrvlK7Ac8osKXX7sO71Gj6NWKZ4GHAbxgHNkl5K82VxKq9cefz
q+G0hRmXxN8VX+haZrp/rEtFDQ4L7EN3dOTywy3+oUoeQtxJysbUZxjxzODuhyom
Y+TzdI6w7kStl/W/N1MaIJynXY98YH6b37LRVOquoA8LyNWVUyN34MGHjwhaaoQ0
G1Vnj0VbyaxBjvzLWXEXfn68as4o2ND/Yhpf670JlztPLJArngnenMpRDpqyMq1q
9yIzhxEqHOm71x70PdGhmvMbuSvqLRvSiEWlRyJjP+W8rTo0zohAucZp/hgl4Ywt
DGJbVdmoDLOjCTvb7e2EanRXA1tgTy1QGYhKQAAPwV+QNesv2aA6OKlnAIgTowNM
3BemfPdAaeMzo9a++soTW1B1MMo+TrHRf10DaiVCuShj/24CQyOdb68uhRzihFkF
vlZnsFWZ3M5Nr4moLX8U46NnKhYNzd9qda1Sx/VTlmGMnt72JTHKyExMjfaao541
jPf9SAt1lLwv+JAMvLoOJUkKpY5LyHSu2C3EQ7llJExwuWKikaZKI1vmHz8P3lfR
+DOI0Szoc/S+RVLxWtU75WTXXsSEEVa3+Ii9eniiSjAsYuMJwplPVfafx0GmnrjY
kOxdkXaakJdHxyEpc3skv9B3CX1qiRxYBgKr5C6Zll3qQaATKydh3k0ESjOO8vs6
XdDC6BvQAoKx3dvNLG6fXKwrfr7D3Aht1sK4K86O8Oq5e0S3UH1iSkMCd4yE1C1Y
7Cd6oCEzcnp1qA2LzkzcbypK41KghL0FpOyAetD/uOXv4QS1p6b7dE+iaKkrlgAF
zDYlWwkRNbmNCfUEtybnV9cSOzWv8vJG1NnBErNBMvbi3l43/yuT/rhe7o3PL7DM
VCfU/PkxBj/bNR2UGsqSv8v8h1yzU32eh7T8x3eZFBMJIayW6dZpvpdfvQgYaNyh
ca9/cXDUFCg+3CiwEQvrb/YRFWkQswYF0AqcORNBH0DWYw066dx3xBAyGs1ijsCq
BGP5wdoLUrukjim3Ia1EJMKYr6wbV5ae8RaqO94BaJB3+ErW4z1ngOIFPgA3AKTf
orXemkDbZKqpjvQv9z/OD+kUi5PeETh96jcPHNtLFp8RjybnzPtjHqOp9FfjIT3R
4/utiBTpzSvS064mKyClmohTXsDOz2m77yrDdT5nTkETurxyUd7nM63mYIhlkrXt
ESfES+vRMU1jdQF6k6Kn82F2Xjphv7iBYYGwlVDTnQgqvzOVUF9cKe4kbLHfbLZ7
rBEZJW//rIiOxoRTybY68c+6VXxCaGqJB9wq+KnmG8HVsoGuBh8QdNmIi9ZRfaRL
ZajFfdkdOpRcPrBNtguqa6/7Wqepyu93A6ZUeaZPZBoDOygxaoqP/BhrQ8IE4hbK
1fa7eNihKyVAsTMhzJWkALlp+L8qz2hCf8GhpHjK8IrCWkf4WYsNvAwdHG8Enc92
dLk8/NquSVCProDgpM+hjTAVrHAxwjaITrPzLY5YX0JRRUpzaVsDFv6LhxHyXsTj
foz3whqlQEbhM65WFvBfkAY+b4eHBXd0JRsqXCaYT8kbjTnrXl4mnWDxxiWN6MLo
uLrBQDL3vWjrrnNELvvYpMOxusAC3uuvIpc4oDdSfmnrvFUnPFnXxvLKDnr1lMxc
4PC3STiFyFR65GaXso8GYX376DoUfA9/poxs++Yp905lukzMGxV/XQBxfSL09u0H
mwsfvQzQkaDjyOXqPKbKkRQIA5TNpUVVi4mAoLCGdon37T+HEPdq5vtCtqHHJzAF
WVaOpBQANK76OamWsw6TIIXdgmPZcYdLQ3Mw+ZJ/AZ2C9IrZq1pRoGgja3cgYtnL
mYSkojueu1u+ncfc1Rl5E5bcVVYynPg8Cjb2DBJgYJsW6xFxnML1X8Tv+jlS0OdB
MAohiy9PIEsiboLlRY0Obyff14I94Dx2kSLBBxDKmgN1eqJCykxnlhJNiMeO+KZt
E8gsq3ULK4NX/T2GZhA0EZ57LHMrApqbTHtuwuoE6+qOQYJ6lylBPN4anDzEzg+u
BLutTtIFM5xrnJuMNZ4E9gKFiOKTuuyI/qvLWcHWhvrLC4Ckk4dwG7DN0hvYoSZO
l6ESraP60uJvSUcoPwTh77+1WzXAVOm3P+a9I9r26GXzWYo7XypVHZ4xDorukCqd
WEJnF1s1O/hS4ztd3G5QNr6Xzc2CJsYNsEd3PCJgacFhiAr79DLnGMEFJasM6yR7
G+oOFslG+cS13VCRVIGJbgtP2Jb/FuV/waP9oU7blYiowFGsNlBaqzbvIga8EihX
hfgJYsslAMWqu0XcEwuMMEVRv9oTmDa6gpMsyKvMrk1g+2DcIdbElq5VjShqSHv8
x7BU/9xUk0Ule8VNdfAmz8u8SiJw0OLKLUF/Eh9usmjcDdUmrmZE9Q5gj0ELDi5B
BQf5F5lAhLzOmevJCETzQINwL7RbV3OCcnxTOk5t9+xGPahvvcdb4X5qpjA4ogMM
AcXNeYS+OyIRfRF3mNMI4s9oSZwyf/fhuPeXh7WlFgc+fW8SaA4tOJoY7SyhzHDX
axoRmqMGRiQm0JMM8WMuNejLyB1JMUikwyO8tHtLHcold0EdiwycySKogjS5LpPG
QR2o0snxaEJLcMozVYElIg==
`protect END_PROTECTED
