`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R/yXfCLAS18xQqDmWu/D/Ke0LKUPbaHndco5ESRiMbyTcU+FQObLbCT5NL7XpoOb
NQNzT//CIS62f48ndgmXtD71pG8H48QyWTcSw++soYn1uL0cL9+peY5HLIsdpw0w
1HfVsGIQf06S9PZMn+vPAKczC5ZCZy0STb34Tq3zzaEiy936uV5KqKXdhlPHlhw2
DpxZK2rj0RI4XH2WGTWCX6kyVpPSt3woHwaxYDZbv7MZMdXMNGNhzWTsjjyZehK5
SXz/HkreNHQ3o2PXPpsq/10He2cpynMRQsxcTtGmMSW9S2X0i1WET986hTFopCh2
ob4QPDhcVKoHaRUUWSB4EAq2Jq5YNJFfr5+RKw7/WJseeSa+ndNyrWmes3qHEGpx
0r78wso3mVhk75w92GQnpt1q341Mx/pG1k5KZvHLAr0vqjGjX+kNM6NqOcTMgYXr
frv12xC1IFD9fHlQIpWLrA0YsMO0a90oF3jObndPUvKfS2pisxJCeI9fMqieazna
+WeuRDuxNnlVF2+NaWk2xcjOaY65uQCX2SHKmCsAva0c+X0d131UPVOIGEudigxh
QW2P5k+BSf1emOxfBsAPuYmYRlMk0CVmYR1jEAdmtGMtCbZB4ctfS0YYqvAAGiZ3
+TU9KDGWhIlhtsnsi2P0i+3+dd2Xmfy0kuknT7FXYI0dmkClcI3Yo+YT/x/fyOk5
`protect END_PROTECTED
