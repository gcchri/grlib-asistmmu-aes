`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KJ03ufBE6k0MHiTpmkAqK4IbvPlUkQR9uicrEpbYtenDIizcUNs14Ao+gzGyxcwo
iggXztLwZ3JxknZFgN9U1wcFjIQbf9OhizHCaKd8pLG+6ofDIBqnX/OwQPaKHbNR
DXzIpoj7X+tZqAu4oyuEOIIW0bit2ZaHByQqRY3oNdrXEFxqGDPZ7HB62rkG+ujx
ctpvNywhN1MJEHxi4RLuP7BOqwioRcjpIIH6Ndlev5FL1psMTAlzg+K39mM+ESXa
UIviNfSERBnZBxm62FQFdN54xQyAvKc3gYx5kl8WhdcvMK3YRqyCF7urxpakumIv
vdLxVJm47fZ6y5RQ7mGqwn9rcrXQ7PsDXgbhJPqRLVKSpwzaxUvVwkyVAtrc1oa6
Act11z1KxPYtwtAAVSdhd5KruWhUr/fIRBprCAr7lRorUoRcCovNQg4U8usBuY/f
FiydQ3f5VinS+UrBkA8M0zqaDSu/wtCy9tCxLRFcG1TgbEHmLEh8T67OuZ74OJOY
VzIgciu6usWZTVhAhk39AJgwop4LNP4R/gMfVL2INiw5iVa8Y/GqfshLfu0T3jcl
6/ewgqhUf6PIwOexQvmPcd2Ljj8A0kSRlSbOKRrCwliuU1e+U1RYN1F2eJvUAm9X
+a85VWhRFwckj/RDH7lrESdw7dFKK1/NKnoPLuUZhdk=
`protect END_PROTECTED
