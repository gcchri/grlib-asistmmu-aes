`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wV+9ZCayRfZVjkXDcRRse6MVfUS4exVA+kRW2qrPFYVHc62zLiNPUwKPwpT5U9rB
3/J7rD5bpW9L30OkNCZWxmjZxzPkGRZF+4xBEH/AmbCbDlIoyZSdIhU+H0XFQyYl
qRtIGeIfPDdhz6royODZkRjKaoNnh8m/mrQ0YxI29rQggm1dwf4DKXC2+52E3RsV
fzE43ZjgmNb/2EeTCPrJQNDWxbNHlqV9JykSIhCFYO42jNZsGAZnid2frbQdMjzZ
ZjPbFEio4migI8Cyx8KDtLLeafWzzscwe++x6ummrCFSKx08uUlD3N8jAcyH1jOe
yMQ5HCHFZDQMTZBOmsPRa8z1D1rVZnQTybWAxhEZXZEi1Q4x8/as2nachyxdK9D7
i3z4HmpVe/W67qKe8QZSY3vw8ZLiNs9INmB0FSYmWwnVrqL6ghFMCfTYZoGN2F+2
F5QsyOt0LrLQiseOnvo8x9OmXDmFBwdn66d6pKxJDg1aJCHaKajRnW7a9H6lIMNg
dcYg/XhMCOqeEVpB8V9PHKjcfydU9yhnMJ5Lj3ULmtX8TclwCLqOFUdIsfDbIYI6
DN1Sxmq0ekHhg3cFbEYGGwqEhfgb557o1q30irIu3MO03IfifjGgm/rKsQvFDZc+
v+h2s/NScLfBXQzR+X9GEAXfLadBFgZuOMAJtgg4s5dFI5SHMgcFmYGI4wKs3xGh
u7/olr+70GPjOaSelj0wbVpb9s/HB0CD51N/2vgdHoKH0dWx/UKXysvDF03Xk/G1
J0+YSuM6qNLOThbdC6bBdsc941p2Zdvhz3Zws4lmCzbSauMOsAO8GfHZF4312kO+
9K+ZpfrDSzF+fG9qWq4iesnzkezYEvpIiAk58AgCy7/UN/Qq5zdLbqPMv4VkjXGx
S+OV8FbEhL/0sQuyJcQI1+gCiJEv3GWypwT8NfBm+4lWqsfgbyZ0r/dkSmQfNITR
gNtHMXtDlzoEKXJVMk30GVY+rBzxS4JltUnJagLkuZvUMcKQO46gmV+xyFeRSXUd
`protect END_PROTECTED
