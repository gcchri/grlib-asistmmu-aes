`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
62tm6s+BwLUyTTwwsksxbK3qqBu6mr4g+DcUft/nlEZo/H/GTle+gP2yo6zvkqFm
/jYdR5ZEwjeKWhhVMNaoa75TahXKWFOJd9MaCvKjnsbpDR0DX19+/d6FEz9HYgyS
Qq6Ky9z8upybdTbSoyivhXPeOQ/9yzLD5foBzfYSUctZaCo7avFVZz80A6W1tkk8
Y1N60imyQJEPYgLUd6auqyUrn3lA5QtOHiUd7WR5JvghEttt7yVUiNe1F29uG5uo
GjTD0f9F3s+N+NP932/2S8fUAL4gTPO1hLEtIRoLGytAd65WMZYYfhOSWfCMcRdf
36aeGyhbelbb/iNwZqLtNw8OKPP8qGWxQvSFJFD80pO+3NzG3dE9EDFdy1cFw9vp
UObhHkMJXuUqIoHKMRjUNJ+wHQCqroH4Pus6+EYcX7LXHgeX1k1/Mucnb3qamb2p
z/lpN3UA4j4yy8Gf2Bqm2gAFUvrhDzk61xpj2mJ0/2PQH/T5O+So7XQp12Pu8Yz3
Aazc3pE/WZoGMN/Z2gxTXH+gXn7JxwkFYR96nar4hDGxZvYD0GyhjkGssrc8yQIh
fT1m4r4R44hzg7F5ooQbgNpvuWbCcy6jymP8/ukyGK/Y/Hw+zrC2wqhp5BV4L71T
4697GhrRl+r0fcXkPplo7Upmed9w9R3cgwH4YgkCPOtOZsR6AyhMZGg864aZiEUR
8kYPsjKnUWPCRVHkntcllSWelMnxovaLBLPidKQxY6vJ1fIFN7RE3qpaXnrzEsXd
gvzYb8PdY1rPnyZT3Gzz5goEOGuBKgjQ2XuRBXrRiUCuXxvJWKbJH1/L0pGuWx2D
/MRIYSuU5G3v4AJeyyq2c7KNXzLJkmnyFb6yS7lvdssIH8HuzCJAgOLZqAILkTiU
DU3mmhKYgGlihQfCPRwiHxJVC7G9QZdf9heb/ws8vHNYRMi8wC6Mt4R/gJDMSLCL
68tfKveoR8uKjsKZXqvqIY1hYcaNBPdVes+QDTaE5bZ6JnRa8+D6Lnlz5xdLP+sl
F4ZhLd6Hz6eDcSNrC2oG4O0MgZco/CY0mUEOsoA0KEmD4dyW6RXp4FvHkzEKNpiU
KkVjaIjOuTFMaYRKyEKT2hsEf+mFQE43sClboFS2pF0Ay7UdcF5vl0I4h9diABzk
KsJdmDE0RJfcFDuVeOR+ziPfK4iFMv8Cbn5BVpXbziFTQ/iFZEHP+rOj9e//icmQ
WZXrbYezvnAV3eWt7HaysZFxO6IpeQIBe4evvcgiuMTBe5RW1fwtufFdCXBwDnsa
IhjEWYBptF8f3m+Aj38SB/Ri494oRuFQvIQAZem6wfHPcttIeWwFkTrSiLzX9HtB
91QFfSehkRjTElo++3qN9Qik/HwSTJLS5NlwO376CQewsfhhg50wAwVppHIyHXbc
ic0DtefjevuS9ArHDG0gg5ZdLnBn1ZSXS4IDBgvhwiGANhXeJdtFNIg1MyWOB/nv
7oTZWfZfPLWozbuYQUaAVQ2WG9guiho5lpy7YdfsuTOAymWnHEKeBc9Ts16zW/X9
vpB0SZN+plyphgck9zHDPaKynVpTLNjEksKaQrONXjHWWxhvMe65Kwnlt9/A/YJY
`protect END_PROTECTED
