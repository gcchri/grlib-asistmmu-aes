`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pPusq0x/ekdC2Kx6oZJPgRp6BgA4GmsR/R2qcX3OChZZ3sxZ1xxcJNxPu8yFsu72
Z3JC+4g4vj8fHW6wTVjAkzlxczTz9D1CXbJ6uwHTe9bXs0Ah1vXn56EHZ9FhPw7I
40z3RmMUVgav1YsZkqcILgaIiSssdOE7AHlByL07NakLkfQKACb+AAhYTVwkkz1e
sMb/RIRxgmIlaoR9WINMtLUV+XvqyFGfvZufme60cI1cd4NyOP42AL0Wxr3BMb9R
D6gmwAObBYNxxbXtfmw0djjECmvDuF0zeg80bNk6UbWkOZdL1VhoCicIEzOExsAE
a+jy+fgVy/3zB4IZSBbxqZhzAZP8ilSSTiwCW7UnJ1Sw1WcOFxL4iEnGOgwYCc/m
Iv0okvNmJUHgPvJiVXhZowhMe7ttYxLeBqP6ZoaKSgpGLxvuX1FU7meDXa1anKJa
/ukegZ1s0yETzx9U3IpA2FGnDiCkXLrAtoJcfIK/kZNbBWkDOyniglxCvIP7orA1
2HYTgW2uNLvZzSQ8GcbsGuEcuxMqer3NjCmt5F7VEjdft0oGIuDoogGtmWyXMyP/
HeiY76Do+T8FPYG3fq/M4f7Ccz9dby+PbDypP6ZverjOusHXFbECEa7Z8DlD1szF
61qExiVZiSwdv+N2XQ1ASawzrH1XHSrzr+h71aagpJ6qCgB3u2vFyo4TPU2U92QJ
`protect END_PROTECTED
