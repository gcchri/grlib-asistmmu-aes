`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IsXVgKq5utrnugtV+dGB26TRZClQ4IBA2mJbZquFodnz0KTowVAuBV546e691fcm
hJ9vfSdEcBPy7g7E8ke3aa43N3dGvjcxyRDXjipGhl5GLjNGusytbhP/10kolpyn
bjgtzSvoHQ1rQPloP9+kZT8STFleHkgI5k+UIcSmuXuD7m8jsNtT6w2vAhkHX4nA
FVVhSsSkW3rjb6bb2MJ3RUWTpzFnACbni5oVZ0eiQunI9xTfL5otIcGigRMOJ6Z2
r5DDsxSKAUP60AqRRNv12Zkf8cNeCyxz730Wh7hszhZM3uwpgOxIYfdducPm1HDH
I1izU6dhNSjLR7YXZJN+9JUYndLj4Fwhn1vHw91dg3102eaq1WUEuaiaRrAr+3JF
QvC7Z0OvHzNtMKkgM/oBD1utriFCUMTFp/GI+C+hlC91uzglZN17nJclN7o+ggG6
1b5nog/X4Hve8DvM0bBGx2uZw+SozHVaJawqBs/L+v6LnusoYUpDkO4IvzdcD+jM
9+y5Hocdx2zT3zVNW4+mcT5KeBF9VVkDrd0KCD4Q29m/c8gtftowzWo5Krk10f0y
Z0A9XudFLtu8AvL+xDVBPprJt0soEm02hvakvQgzwSSah50YzWOQ9U2flORVR8ms
ZZt6UzjvjLXgMXUVUDTvZqb0uh1helXkxlhn1u42Hd4bJgGotkuV2qPkq0RpG3Ol
LbE9sLzhFXnvqDuptrGc55dydDKf1IJVYsmktJcb6lIaFYizJBO8jiCKaFxHEek0
qD+AO4UlWRQ4Axyr3leBws3BYnkEEGHT8ofcQe/YAL7dyUFPvSz5S4wd/IXYFagr
au63Y6UWCh+VtiLhuGseAZL39HiFVG9d2bseT0Os3mfU5A0zBXBO31FeOmd0N2vi
McqdfL7R+WAn2AP4gr2XPe3lgyza3b5XJcADvEqeMkZ8XAlm5NZrcdkNS10X0bWd
I564yhIRtRa5VdXxO/BL2Gbza1vHrwzGIIHgz02ugwjmL9FdgTfkZ+jvEPRkYJ+g
dIlFvDfsrFMyiyWQQPSNi9kkeBo9N3DUd34neJcmrl24Mv72EYWIAZX1R3Jk+h88
eSx/wns+sM3qtRUPxk9lo9rp21oCk1efCIZLpB7BUL5JPbDJExY/it5Of0dMd5zM
ihvQfqUdCXHO1lt1y4cazu8AXWz7+EHGlTDZsEO30aI8YV9GTF21QxfcTKqm13wO
wGQrh9V5o01lSoGLoSUghdQyGdXXncR4EZTB52XGf6Cinm0unTSA5qkgu07H1QZ9
JIRBrcEwbMgnOj9uvTxyQfXKK0WKK6AGTeeLdg12jRhuYZDiffUJuK4n/UoO4olX
vWgigAJ6YTKHcDV+UTs/q4J5aZh7GXwQyjhAyEFJKJkScBw9is5dFwSGNmaarHOY
yxTzOhkTL3aL5P8TbLE11ucKBRKoGevPGIQfgstsZjsel/ZxVz4xIus6Me9g7LWl
UYh3XmhuXO/62xDfN4//HkFJXFoHkBlhZ7tummErTLs6E4wsr1BqLoKMrvEy6+Dq
FSl2izr6Fps+ldpxCOIeVXlCuEdo1tl7CGs3j34yXgJ+E6buT0Kvfa8s+kSNqb7I
fO6oHclCYpPbk3xQVurCqI6hbptbnUDUQQmjJPHrzB59hxjWdzNSE82WID2dSd/N
lAQ1dMCQKFAREA9Qhao3dQUsXXpXewOGtBvvHK6xXxmRXKZzdvpywYfqQaeclIE0
wY+ik6dv9xqhTdmdH/4DM5dx75/qEkgNnl2kL/172cZor/KLuoMdmQRw+3WWWcVv
fsiVfpdwADpq7jQ7j/GrUnDEuUjOrXd26hs806CuiTmwbVQTnGnb9KOhw7pTXm1j
j5OfRU4fdUJmU8hM111EKnNRJwz51rRzyH4g5SF1NiCRjgf/fJSAW+2mn4h97h9/
435Tw8kOtaojPunDqqshvKnmedfig7Kq44WwEKm4LiaK0zvW837B16rSVxXDuubO
Hi4I2v5ZrfuSszigNSHKF+0rOBoA5dQgxk8oWIp7KwICbXU1jYqi1zQDU4yXRRRc
ByO721GINE4l0nPg5qGFqqP6e2pmRMc6HD0BrsPoKhjmrN0xAKgd12nmxpnV6TWA
2ouHhockAH8XfcAq0VdDNtxbCVG1ktv3zE/bsOV1ATE4ndiCWbhxckOZfWad4Q9a
J2XZD1kX5b30h0na3mvo7gqVgkypBMq9oEJQ6VRnDgEyVQKAgbAxVXL/iaa6BKqy
ZxUiDtUSDdishY3RxTzIJ7h52dd3FTvo2fGzQQi9aJp0XKVZq22aBtXsngl0n40n
Eykp4XnTOrJiwVHKZptWuexltWBLQSgc18NnROq2xsJ0G/sMV3hWcphtmOmn9l5o
3ubcbYuifvYM8TJz+EYNKEXnBADdB6/qQPA/KJ8aOd3e0ruG85WnJUSzW62g2bB1
V6jvSMZGO/hiUk1/VEOzGE097drJ+pC9bjTXX6oV51TZYSEE0SBGvnOZbo/GgcDp
NN4hx+IzDRuJX6NIQWZbAbCH17OF4KpCFYd9CwJsYvqbel0QNm2A9r/Y+7VHASAu
Uku8Vt2HW77Mhz08HpAd0WHs/siAZXcSAlbXTdUxnjaZeuN/bPt7K1I46BRhSpD8
XptAaGuu9c8Qmb+z46WEUdatsqjDo8nzCkD8JWRNeiEIjXtMYXxN5/JfJtfBSjS9
35cbf4f/M1aIqrYWCrJRMDhpKxYj3ibl3Y+TZxOwXAvSjrH4JqPNh8OQds+39XMG
7iNDV5fibgXa4nKKSjqIlD+bwA4wHKdPxReAcp/E0w/7RnBuPHSX8Ay8AhfXrdEc
fV4qqXZp2LMnKW1XVe+3+jcUYNk3Lt0Iwy28ysldke8r+gFZNpJPe3MAw9aYOcX3
qYXUMmnyvjf6iZ4TWYNgnCN8k/KDcU30tcXLmkx4cg2DUujxRezi4eodRIrqL2nc
B/0RVU7iglSkH/E7a+HqMtS1Tuiir07NvJApBizjeOHg1uKewdset4FZapGA4WPa
kvksuZwFThXIYz5A4zVKxXWQayCqYQlgMYTnqSefcx0g6Rtywc/oAR7zUKTIoB/7
q2rAcRIa8JC7wu403kyS0t3Vrg38Bu/DXBNrdzFYnM2+G6tD1+erXcpWFMcE9msH
HmnGN4eixLVUITkq/pJhE9uChmWF/f3mPq4kkUUkZ8yVqm19T015BcsJitOSLJd0
AgxdDQw5gRb0LH0xD+NugTAupUcJISldpvivF2HN6GGkwvCFP2kAM3Oc3HtUO73g
MVG0kmS+s6G2AGf6+ApTHwxQQ1Lno2zu6jNxacHERW6OWZsz3c7o+cPL3/GNZB2u
J+i4E5DAjHkbTNBrsm1eEO44ntZttUucczi7Eh4ootUGMKKrL0dIGUM4KfMNWIk+
C8R8xZbyIdh6fkkGz2a6pto9A5e1cNxTLbnsjEij5fs8oRo9T21D/FD/7LIPNRhU
6Vi1L0xrWY5GLABrdrxVPeTfk4DABIglt6J8aGo+AkgAvFFDVlb845uBHFFWAgmc
kg6pd+zzT5KYsfwl/XbIM8bXkKDD5ZGImDeX8yl86hrmbEATdnhsK6ATh4l8tlAO
m+6Gsb04Ve4/rBj9YeF7xaJaGJRKEHDxE7zS7+R7vccNV4L4jqax+8nWNWT2RHsH
8sptKWo5W2smsTi495qCkmwYjdwq3OXBhFs1jTDHdWRP5w4f4wZGEOBG9H2uixwQ
p/66W7Li0D0bq37Ay3KLykN+iwkOVzSYyCPfWtjeyOqutLqRxalZPHrvQUlzLEyJ
IxGiIiN+MPbGDArX68HcpMWotjjCvKGRtgN0WM2EnibBrJsIMYmQDpFRpX2sQJwV
v+IgOuoYgGs66ZNGyUw2c+QPQm7mv/y/3ZTjJS1WFj3pUUnnVp4es5a73VgAd4hB
c/jI+Fb8usMzX5EgJjASilCNeLXiRcUHTzVVq7Q4Cu//e7+VtQcWyCaMb3PKY8nD
vxYJnAVba4OONzTqaqKIF8jDB3m30QulaXU+3nl+t/jxmtkHN49ZgrMlw4TQqc+i
/xrrSC1wBHuALJOJ/fU5usOx581a37it7HZn0VQcwqzkoQDuIJonOa9fRZmf6G9h
dpd25qeKguMjxwErEreUje9Klj5vTSuSYFztMyuYKu7Xl18eX+uO3BehHHWH5T2Y
Uql/AXXiPO49q3++6gPjzjZ69l5MQ059EHe17rbBo140fJRUQUeo5C+cjS2Yh/c9
w0PAZJuUwIIgCaDfOmaCc+e8URhb0VeABNP7hCFYpeBy21W3S9yP+vmnOwXyxlli
2fZx/fhZezSwYm93fO302bSIW3QFOCSZfdGje9PYEAtiaIe115pkd4sv9UTtS9hl
DO2H7CgN4zTFhbJD2VxVEgQ+t28KMDeH074zZ+CNkoufNA4tZ5Xe1yn/S+pJAd4j
i+G8BfT+H6vcX354qbgmfLHmXLg/PIUYRpSizO2eZ6yZ/G4C4fZ84xS+vs9gnWX2
6Dj31DzBnDkAU2ks2lSubCv59Nmq7CZUEUHcuHYgVvZKrKWnkHb64EEGoD2BM//M
neAmblTv2cBNU8TOBfFo43B+hdNTAPkV7W7VyNICN2z10Id5MVwj7uaD6Cb8LT0Y
6ficRtmoy8kTvLA+aJw/+uTHTbfmuqz6Ka3/m9AACr54X/g9PrIvgHs++NxOh9qS
elkXiWy14HGI5PkwkQMPRVo5LPkKACZ4wbXr9DPLAw3lc5X+KFG9o27tBbbnpeND
2LOF11hRaCjT7qC7TL8q2kb6l2fs8n/FxKeAJGHwhvbEiSbAqwWFaJMLWNgCpoVz
B4A5jAwDH5kCk9sHkBslEpSS4wIlC6srA8g1Ck234arevHUSNKmCWQRdtr+nY8iM
gvdeek9WhL1J0I0yXXuXxP/K1dJ04E9R4dvPTa3buOKViElAEqnJ4X1xVtoJgGXH
L2UyDhy5nRiPSkn81Jee79nr+CXkBHYIoYzI72HolccZ1X0F15XU37MYGj045JkQ
ya3rwKsSdjxpyrvvGNJf7kCZFHXSxOfY4X5Hju7aiJWQ2sFyph4bD3yVeQU1rGbs
FK+xqtRaRwV6z7GbiExOU+C45TBKU1YIGIuWpqGoSp6mwH4/O1lBPtSSgXn2y1+A
pX13N1Wg2AjVdN+ybLCxIxNryhT8WUNU13F8ZPUt9/ulVCVXjbrnxpd8yT+OZPm5
HhWdICMETKvbHpNk8vzL++B8MMcwIFybvciz8hR25YTaA1ind3QA7DrHcRoxKh9+
aME9fhzoJ78SgtGTE427SbKL3H3WdXpTPXgMrCjpviA+32JFAs7Q6E0O6Ia6J/x9
k075zdRqJONCJD6njeePqMtVW4Iu3oLjXU+FqhaZxVuJ9b7ytOUDEcjJ0B7rKXNi
NIqUZw899HjkXU6FNNn0FVmhNotWzLLBqvtyORNhMv8Sk13VbQAdpmXzGpSBYZqw
sbiuWN5vfm9CbArM+NttC1IUHgQ212bW7miaa/1EdX8s5dUzw8FIr8tWwA4v5AlH
aLRiJ9XPa80xE4VYCwkLzCYeQ4Ml/NEwACwIFm1N1lyV60HJDM5xh2JnlLHsDqzY
3ulW3M1w4005oZt6v1s8xHBOt4qTC/Cd3tNMmStB03J8ThJYLOpTHSJe9Ad4qbQE
UrKO1auYFMdbm4FaNvtgejJkH/r2bKQ1I+cqq2NrQHZOCOg21BalwmQkOE5e+av+
RE2qBTyl+PDqY/UYbrGqA69Tc7SOKozwD2uEAk5RinRaKzu+0G+6HtMzpIJZ1jXE
kEKP0XaAoZC6PpRKUWemJ5UZJvq56jQUU2qHQJHPYnx4pIcLhhQ7yz85/Jb39m4L
EcoH1hMo7WTCRArK9Q1ITAiumTprPAheATuJds3lOtl65SmfoLKDLZq60Xhys0+O
FJK0wOukxcVoRfQbP7Kx3KWP0z79M5HrIU7aiceAyVSCfpr/qKITfNIL2H8FhZ30
pZOefEXIlJ3IYlGJPLzE2lV4FgxgMv48uQzt0qy1swOGJmPrd6yg2Jt0/DQfSovE
1gfzUC56t3XWxKNdbeOvRA3NT8dk3yajZfuhxbuo9OjjUxcky6LapJf6+wRJNGTv
AhfyMhueWGNOnKtIntk0myexu+sEw5imFXVH8cnzJ5VUh4bV+vi/bqeEFsuld1yd
1VEHNfEVWp3o+jZAFuNKN5i8VT3abZwpWCLTq3nq86zVRnuInwqfrlHsY+cGplVZ
RZat4kdxv7rSzUpRCIeqS7EljwSEpV+7Cx3aENniS9OZnS4qgV933CWt7tKKtFr5
+BKoSg6g5z3Ayun+uYuNWo733UCZKwsmEJRMW6qkPYsOS3TpCVi0nH7Hb2jUSvOi
jzOSxpjz+v/rDOT4zmqlRPwnbY24bzMJ8JKzSKHHboywYj1i/e/cgfml+iuQ28Ll
u5D0AUagxvgLXKPfgsYpoZ72t+wXYaktRhzsC1AdVgcDJ/6kLsWUwEOuyOftjdIE
rCCa40yKFejJTl45QqMCyDTPRMAxVH/ImZkQIrTJi4+RLlgoq8KweazETbVVFw1l
ppx+6flfJk6a1pOD2k/Yy9R9pQi/49waCEgldvm9q+9pFNJXs0gncau4qq0v5hZZ
uKMVBKiM321jge8Fe2xXbeRm18K2MAstAmHpBotu0WqK6ITg2erViBQdZx76d0EB
lZLbCz0RtNxTq5cyeHhk26zOXpodqm28yf6rtCKmPPa3w4l2JgQ7eMWLhQZ869q/
elF4iiCvl5PpyHZTW9JR6P4Qf+HaTq66z+fN1JJ1Nf5TP+Jdzsi+50t6Iht3c/mb
7sEXDVa7Lb0TLwGnCUCyGZ9Eo/1dO9L0wO2FzadDTvlzggY3/1myPDwKmR1BAeAn
BMQ4e4Eh2XlGLnhSWRx2Kec0QU+vccNPhTGv2fHsHfs7A4Hq4EFhRpgVWBF1xf0M
vUTKVEC8BGmnm5XRQvlVKo3TsJsLOUJIyJ3fPPZlRaKzT6DVJwPEJeIczKcp1VlR
/xlnfz4Oiok04WJpbcDaZURzFUQ9gofO50+lwaqlIJfLM7fzb7vkH5cWaZLJLw4r
QMjJDbNfF0+dDPgtRfErjCBV0yWU7nuEsB7BwQEakrUgiCwvKeKBecpV1QxnitQP
2vDH+I34tRHCx/zimCuMj4bqx2gj57krPb3QZqaNibRYiKi0CWQoJv2PRrlRc0/K
varRwezw8uWk97kMKkDLBgYy8eKmGgrziT+oRkYWrP9rA1M7UdwjfZEwQC0cq+is
66uQpKWFglifxixuE+AnHaiAdEUuRixTyqtCR+iDx4cd5ptXALwQtbKS+PIN3c/d
TSqUDWzaUSLkETP5kKeRQOiGTBLyXEklivXglGEn/vv4Q6yqVaap+Fhp0xFUvUb9
YFKFErbUIdw0ZggO+0+OFPGVLHKAMc3YDGcsIFzW96OWxgSHveJdcuP4CuFcILr/
NvAYB5fvWKMwdv4LVdsHDw3eH6VeYlWC+GHd4xFulbYtoWQMzYoDrS5WY4aKL5ss
UTMvEXCQfIVQI3nbpdlSRdAamQYcnxmzAaaggMfmu8e5jElr7AYPCaRUsPjgxDpH
h+7MoQFl+9/xk3SocqFazEKy/VeWbKZg2hkeWkmtePMI/joLYXohdabzV8ZKmg4m
t0NHK1PN1AE0YwSR5XcffunueIzDgDRphtonzgLBzGSxOA3DC85xkCWDyubnP7k7
VGrrGl1UEoVOTtu8XoqSe57WGP9csRPdkg4B2/Yr0mRq07/vV1dncq7ywde4soCT
CDIZEM9q7imlfTkaLGfJn+zbCvHAGXSN3xQ4eQIbOXcaD4PCI0zxgbSUtdt4Ri9i
4wGqkM64us7NUkuJe+cKDNMP37E59UV33WpO0K2GNg1WRMKz1wF60Dj2eFO12eHd
bCYmyOVLBgdYmrGFhmlwTdAULdWwCD3oaxCN4UFPOU+vXQGAKOD/y1Q1iowMJl2H
g+VKoaeM1LnJOHwyJ9UusICm787CL1eCUgLGZdGi7H3CVWePQ00tOnJSITxTdJSs
JqWR00SGAUW0GQfXc6QhJjWwN/NQLfZA0SjZciJnOBfUlM4O/E3Q7X2rCDA2TT+K
Pn9PmRMmG4pvsiXGS11XN68ZiHZQLDY3tpTyLVPEpSQXTKlTUNOiTjS3fqXXfkfr
cBs33f6V7nDATS7FcuoQ2RrKYG+QUlrPhOBwfQMa1RQHgvO/QP5t4xXxWCbY6Gn8
Lj7w44LpxnJqPOjj14X+U2slhqQt7R78r17JHZfsshDE5jUXqb5/bTtZJtTSD4dw
y3tmwvFDqB66DLdVswBguNycoJ0364caDkbD9RSkV9Od3BJBB7/QcvZMZdEiZZNz
6JQ/HAYQ6UTB5vLcmXSZoVWpWeoBxwg2DIyuIDvOZiAPpr2OdVaxGYOxO404xb/y
nLbgdjdMD1i3g8YoaTn4Ge1bWDOq0Rh6Q1Y9RqRiydpcc3CuVDEsCORXue7JJ9Jy
72WBNhV5pgMCtymRfc9Ys5C3HQhe20h3D5WhQ/Tsi6XGLpHGF8PTvmSRLbNioL31
KwaXignzZDYihkLQ3tTD0XP+yA8HI1E3X+58EwPrDP26nTEHh8oVvMUvgR9hXTa8
PiiVFh4ZT9k3sODrBMlAImutrpJzKX5MbTCscBWBoR6pP+mdeeH6UjBKuFcaSyH0
xduC0ygZATyDXjjEIT3ZU2NysiZVsEC1gSvbxzughrXVPT9uFJz6n+fGaUx5H0q2
QczkveJj8B8a45VJf+inrVImbJ5UfsgffPlPe4dZyKPP+buw8zL3baH+bfUJ1S3h
7+sjgGyOn1K8IA1wug8x44sWViiwLJCdUuTNEPuT3Ph4kTpJxbdud0pQEtvyzw3Z
J92NliO0R3+lbA6ZMTp3M6s3ARfQ5Q8UNnIwZxHEeS1RPVGjSYFzJyoYDOEb2pd4
1qWCRJR5uFU+YblmPWy5odOBZb+C4+bA4q2BQ0gyXVyZH6XiTu0PG2COH9EYzupL
gvI4sRR6f4A1S8LkFWjUkzJ42jioiM2dgjr8jkNFsYJMXXMZDlGZ81FYfxt3Qi+O
NjqTrnKpR+6czkjcuF9EC3pGJD8XkyOYtx/P+IDzfoK70eGfGK2V8MV0rf9AoqzW
TU7v19F+rGniG3NpHR+yS5xT3BfwAirfFf/96yYxUk5NNVzwtmbRm2vzRa/ctvJM
kPFuJWS4sfKGtyOFVsdn1lL4FJejmddxtkUZpGewgAAmzgnV22+Yh4EmTCQNm6X5
3mgnVIWnJzVdY+AM4W0V6mRsQirz4wS5paDfBGtXR3XSpylkecIDa+d1dJOs3Ur/
gS2DpdAEZvq3kR/VS6FsiSH76CJRd7LVU6WyBttMqdeHXMvb9eFUG1LZcnqbxYug
MP4mCT7Mwq7QV+yyns7CbetDJ0G8h9Zbsjj+5FT1FYxau44E+kPlnCmE8U+OVWZ+
U+yBoUaEUjBAVGEtZjPgpExDBpQXeR3pnVF+fmLOSiUh2EDCGQlWMuCj8u9BFIzK
qEX16Ltd7InFNcmr/GYmdakM7mCrfKNNqEj4HIb/iBLv7Ki+6q3qaLDE+EQb0rzi
0Tj43Vuep8v2S4aEq4f+2HuUOYOdyeWSpiw+vXsws45asqk6U/6PDOAHsX1gsDrF
MNW6pmiylcPUh9j+O6Hz2M7a2gPH3LC0ey+0WRAynXQ+V5kiFG7EnJB9etWaVNKa
EV2Px2K5Wk/iQZanJGo+cM+uyd1V4/taG+N100c8d/kqcieuPC9dT1SWjF03P4xN
/xG2fveuSVkfYeCigpHOqbbbrRyejCI1a8HcI05k0L8I+dpDvJBFsnaL5DzzHUEv
0Ar3iFuEOh6IYFu/mqxYCDCnJdJ6ivUqxz98WWf051txG7YQKlr7wHVjCtfkEvAi
oMfjdfMkmyENnTdsM3TQzw2qAhZnbnWQ+sY3m8btqbGwv9n8jeHtYW57FDfE6q4X
iUr+QFf8qA58yynGpXVz51VG4PSKmk9EBkBT+0dZV1EB6IxnL2obehSdVB7tkh4u
Txpu0DRSSr3NZJKOatfXVMHS5Hu2K7PF3n+0XrD2/WodFyUjY7L8IXwoo/QFn9Ed
N7SOLe9VaSmY5ZLdlV6+4ckPDUaf3dmcFbp530PVuhsofHshzYx130fVC39gI5nc
IB7z8kHJyJs3YOjp/IdcurnSwUid1xoP2iTXhgjkwj3zNzokPJtovG5ymKmT0n+2
1OjYU+DxEfFjpDFhSmRiGNfYCXx91vgTji4XcRm+NE3u0cJlIOLA3wMXNes6KY2Q
ZdgzF/swzRF3iirmOCY6Ikqn6N+kLjA9u1XAaRcKYqkEN1+r4ujkRenAHAI8B89r
7kdZ7s0k+GhGAVeNiFStBr2wRhoknEbZmAEnLsDVnx39sCo9NTx5EAxCrF3rq7+V
8HqymnwQwWaHInpbQGbJ7lQNgwgrg3XvRNAPmeg/d/Tar/WWuv0n8WZXPWyCTTBY
aZteOHYYfA8niMNiocgk5ICHQTo2jlt8P4aPEjqXFZc1sJOARjmiex1WA/q1OS3E
dpEJ2FIdnsUlOnMJ80aBIjHQ4XNZ/D/w7X4raQ6tHlKZn9Fw6Yq2Kf8M3iyaDxAh
xy1effca2vosDEJ0w9+wImccGWC95HgdY3wyjn77pSryZklzLf5ZdLnvNNbhF82Z
WMeWodggErSbmiO1ISQKeIXvuGgOXZeLsV7RPOPvjbs/nBpAZ1pDKGd3hZKAyAfx
IsUrZc98i5ZTTchwWZTTDLTegVpfHttuto4D2C8AI3+lMMKISQRBQYQCKdpbuxDw
pEhrytzH8R9R8/a5J1Wn03QoL+kZZ16ykDgRsuc1cdSc3RMZQyj1QPk3pnhy0qds
7rynolFsqM6LjJ8lpGQ1O82/zSlVSXjnYkJEJjokcq0Eh/FRUgnPRb19c6x4jIQK
AF17uBs7dfk9LpGi8Awl7n0yOESbQjWl+QbMnOKg847wBeadKp04wINeii6DnlOU
6bkhXVbMLPrDIUfSK8SjLLCpnR2cs2k5OAT5dG+l7gPQ1ZEb7dejka5c9umyyEhp
LA21NixbD55QYly0mGGa0WtCLUaB4gYCGj/VjmVn4G9t2nPKjkgzigct2hN1G4XM
cJ9R5LI5LjynA6lz0Ia17RWNCZqdtQDcS25eT7YNr/S1ZvBEzmElO4KHs6jQAVK2
yNGSke9brHJLldN0fUI2ucrK2C/zrXPGxUOQ4rV/Dl7f2uMhr7SarrGAhurm1ZLY
FjM5BXwuzURg1/HTSyOcfLIbm5nO1yEbNor7NF3Ap2Mwfh4Fimj/sHlf3v8v7g9O
KO5k3YJlahAyuYVlv1x7kqU1NQ+cxtdFAcCQN5y+WeTFh+SkDjQVpMaTAqvSI7gi
DZ6Eetqmv9E3x5YFj+AMxSCeZvrOE0kG+a9+jZZN1Z+MZQEJvadKaQktQHgAt7oj
MhNC53Y+yqSDXJqgXuRNmwqYsNAvbhvvw2oNpKus4K09jGiuwQB6VgR+vdcukoOf
1ekr8IwiDZT0XCZcygX5vkpXN2SWThR7Ip7wO5E1yogp6tmEcI6RwdoMv0ecWDTQ
nlgqiCwOzdfW8gdAcrqjeLF7C5EAStk1MeP99QkQXIbdzv6WaPmSirUKfgsKjOLK
KtP0+6NRYgRCXWRUeGFtPVuK73rR+JAiC01fAcbc9Df42xwqp5hc6ziDnE9R/255
2rr22+XGfWNkoNRyidNYb+s5tWUFiiaKVSWE6O2eMnSgL3GvhocbUzK4jwsbNENN
NzFDKo+946KYbwggak901Qsk79YRyFxTeZmKIL9D61auRLYAM6rDfUuBjgCutved
35xRIK07OvJ/At7kzlLwcfIRnso5Qx/ox0Z9b+0TH+Btql3IdZDdnFJD3oBsGCpR
pte9J7aqsQIa4pBSJnqfoW/LGuU9ti9glbw5sp9oc5CKmCM/ZGhe1ncV9FwQCO7v
C1wMZaQ8p0NOTuYPJvTJXEHzgiP+1Cd3LuVfSbZUEeSxwPucIJVgssBSNr8aOs7R
r7LZ9i6Nu6c9AQnzmkFIKAHGBb1ByL77aO6HHTS2UW5pNHNywB6oj+0c9hr28G7P
FzUys735j5p83CbXGXGrav031v4FISgN/eCbbomqM7OJQF6EXN6QnBu3pm5ZS8mm
cZv3hviaSNDD7FPOBaI2/TCfLb7gViIf6OwO0T9MyQwnxee/Inh7g7oNQBGmxBsU
WRqCOednVWRFOT5bW4vtj7zZJiWueLuTcyrjq/t4wXpnrYwiIZOtqY4nN3B2wBV1
5b+nNJgvXv+q04sj4PNhFBXJWBiop4lA66a5qAZ8nXocbJKzYwgpynWFvLM0HfiI
/xrMFKLcu+xPEKTtDV+XE3UUBkI3YKe+zJhVTNjc78zdsEWv8snEwrkT9s0d8pli
l/3TZZirpsXX41vPcCrTPxDc92NkpXa5w6W1GWE5CztAsDUPawSNSswBfCPnfCo4
4pXlyCTW9NZDu5g3El9PWmgfWdGw5aQ8OIefSsCP+p+M0F2Ccu9S2/DJPZFcNOyM
RS+ejJZMViRhxkpzelJfPKNrjHjShiWdbayLJOpKjzTzqYWWT6TGvyNVJs7xq1pT
cuxw4yjj5noa9hKDh9FbHE9Le4cMHjKVwKBlGytA1IQdhONP+jpdTUzrkg4Z5L4V
5cvVsc96XUKlcBmA0CjpSYZFf2l9QPq86a/MeqAakjJO21p65/wFrVNL5MoYA1Gw
SkpYuTkm2bEQzB/NK188xOhUOzyt6lbCJ8R1ExIIwQymRmQxAXptESX5buTVjU4U
m3MflN+XYlnJnUMLRJOQkPM8F6lyFXK28Bpthf9ppwFk2ptBj2PwGgm98S4MzQWB
ci+rp+yVsTnJxFYLZVqsADalXX3KnFnAi+NW+cBTTEEKwxPsi54DV7ka1/6Pl2Pc
4G00hws5dYwEpyPGCMKzjzf4BMwS98/kJYCU5TUVwnCjyEryEYJVherUWqB+dHbi
DxA2cD8SPqfppBRb8dtYiJb0bFJWHXipyvOoEDkia1IN1BD9HZ1Nky7IyfBl7xfE
h4WSguiqNiRwzsm2W58b33Vg4sJJeC58b5M4extdYGqCgbN+mZ+dpE6EiaXDy+1C
VP5ma91JRBN6v+HQYvUDe5xJDTlhFsR8et/jzNKygznDKw4mX7zoJIH0jiWyaAhB
3uJq3X4S+gjutJB+pOjw2Th96I1CK5NmVJj6sT9+gnBqQLfP/+BAzKXDsIG6JoYl
FGgRI7PRWIqqH5ftwyMeA23vlFxFr1WfLaQl4Sq8K+Nkiy0hG4r+gifA38jLJZWI
Xqowofl0P1Fuhx6uZWTfZkeT4t+Tzhf3kYjGwjk7yLEYek8K1Ow/ELsvUbFVNVfU
Ht1FEWgOYNGhLcTKRuvRCLzQKT3D/5iKf3xHhSyiCBpPmItYBMeJWd/WK+4lcyqR
qB/I8rcxqX8+puMYUUZl47hQiQeShCuNf4dmu5YZaS/hoJMyGGtQSjDzs8W7fHaq
qKFO0Ursv6oCd81SmwQ30nKB4fiJzXcmw7iI1Aoe5K/wccpaZh1v28Wb7YfydWZn
/VEl23Uf3Yhr3AsznWPQDOL8w0bn5+H7qaOKy6rccm/ZawPlYkMBl7e9NoY9UMGc
8mMiUjt8pCeYOhsL0iIKyT7IMTT9dumunONenu5/N6jntPtc9t+tQ3WObwpCzTtO
ibg43T/LcUHHBaaVdZI6UGCwu4jqt2UIC1BiV4jkEqiJlh498UcNM7AT3dj4wZh4
1CS3WGIfFZRkDh2ZKWkh+9tTrrwaLVC3XQA94xC6VrKa+GLUrUK4YtZ60gBahban
PQPi3qtzSlLWkMUNAgaRhZw/QNjzKPVxYSaIprwhZ9s2RPOzioI8VM608j4FWocu
YEcL3njB2PVP3p+FjHLsQltKpka5yKL9iuyMaY8r7IYS5r6rRGYgmGQCRIXAdv6i
Hb1eXhhls1yaHnBhtVLAKSszI4PfiJ6qU2njhfrDN5peaWPFanSYPSGjMYscAwHE
3tpUQhQj/aY4WHDPcMpmQLd6N9KWgHDDH9Fm8P0LiB1nG7Ro7SJhNCxGDE4JqaYQ
+N45ylZ3/JwfT3nxR20tHLIQwVacaozCF4+Sl2FpIoG2RMC4zfOB+adn2nm8s3Ki
H/OkfnR1cExKdp9k1qhBjiZjEFW1jbidSg793468tBlHrJuigz+/hEzAINmIZC3X
gc1eIS2WBAkQlMPSnwDyCGeT+AjrHQ7sMqKR7wkka/blFiOxWfq/AYMaWTDYsw3j
DHDLmjio0iJ9zwWdQ201SgUh2H7Fkvs436LpvJGuLnflR92vKF5MlXFMZUsV/dUC
Zc7/ShA7rBxz2kzKS/DUuEWbIfAlHX57xtFXuSTcVilpD7lbuB+xKb0hVQgK+fGZ
U1Zma0PQxkmZ0FkgnS3jPVvYm8EzFwjXcJ9bCDoSYYoVAguWZtKnDAe3u5a6DSKe
hlZA6TxS4ulGisV+LvhZd2T7zKihqF7BHla/kuSSBN993Rc6YNWuBJGAutkJvpVB
WV3t0G2IoIpcBIWA4LRNMdqg4o/kjCWRcgY8RuW+cmyu/s5Q6QTx1svLr8ESe8rb
75nr3xL8V8I0NAqqezTpmRKV7jXVAZafTro2xxLMWgLXUSJZPlYOWNKpv6+wdKiO
lvPGFZpLU5nRbMOERnR2NfuFPNuWFnJ94BGhsxJcru1Dnfl0EpnTZZ9o6CDQ1f6R
ur7poxsAhzBW7DYSTbGG4NwPt8dUrvqVSVecvcEhCQ85BDwJy6jalyktBlOhElXJ
I1iBCXE0CRXJX9scNW1MjIi40ytK/Pp5tRaK3c3P3YHpVGQ/+yaJTMugxZtoi5lb
qt8IAclAcAcuPLdJa9Xl8w9uLQfmsQxmN3IsqeETAD5HEaWIKo24vriyiKIgJUw2
Znd6DRmM8eE8BHwwVlMScJonIj1mNaR8PLoEYPX4fmaYuYLIuGiPujdouO+6Ipn+
32I2peFfcQzcDwmbGLgG0F0G+0NfaQIED1QX6Ir12YpWDMnu5Auvv18aarM6xzNv
Umg2Z34cEZTYRP/2oGAjauOyk16WK9bRSrU2xMfVQniyCQ2e2Md/w8HmqV9jgEBQ
c0JTw1gt67uO7LiI+O/wQ7MJdtEGNU5PZBzo9tGNPy81pm0p9aTwxCNYTOuAMlJV
HISHxDbW7zQt65Otuniq4tOzY1jDqAsCDDx6KrmeSKPfaCqlPnNgOMmCIvoqFdog
t3woSM5OPFUAw+k6mfsspr9rs80DRSK8yfC6Ed7AFL5pcyxV/IFxwEBrhWgOm83k
vOchefdcqMwBnTUb0uyhqzEfZ8oC2vI0IyJ65kU42+WNCldZ6N/6lwEiH5Kv0z9j
N0Sq1UkcGiHlkhtSUi3y0qiQuyPWY8M72pOHXvP2lq8Zey98Yj4Gl/C6D0+bguPx
PXiphmx5YEIwz13f6RloChU/gO7cGohLbu77C0wlYM8slaytpcTPu2keUIDktdsz
JghZDmii6JafiLL1jA5FlNSJ/b5J1LOZBGK2RCmvkhN26feI+tv2RE/dpUoHklDW
KXm5VvMrFDIrMAHOyc4qtO0MzGMrWEXw0QKCQoKdyf3bgMiE04Saxq7VBbVITDNt
i5wColUtfoNWbJiHsj2rTb9ee98R6L9Vbb2CEbxh4HDs2M1njDXb8i28HhjiOpYB
RgzI4m+oKtvGOxzNkiGLRsIEqwgQKPVoxhUBXdfot1DpE0EfHoRs86nPdntqV8W3
PB6EomEpunUrZ+Pvh4w0E7truE7g4xlvWZMNyPXYviEsOYSugJSrR/JBLp+RuFfX
6yQ+Xzt9pArqfOYFGR2R15csAcFKKasMqLisgPpl2TTRAU7+oeHZ/zBunvkYW+en
t8Fsy5/kJlQJ1LP9ACF4RsesWseS8LOsothNPKS7x4cys+2cKG9yGo0oQN21W2bQ
NKD94OJ2AbpklK25oXRyOrGPCx01NREeAN7jyZRGjYLe7R8AUh20q70w7ia1eApv
s/OBuPb8wRXc12aUQ9fBTH+5pVRAPJyhjeY/zQ75Hu664K/w7OhKOgK5BPnUJElD
/6ifMEjekjZwsuwpOHm8Kuwk4YGf5EFhDyYLACnoSI+p3XN7rIYbrzvDWRFH+Mk5
8qDyQS5LHWOK4FcA9fSXr796xLGWZRx0hs+S3QYSBtoiEuif+fW08gmPOHxKxWXQ
lRQdAE4gFsB/QE1b0G44gDwpQnuKNKuP0WfFccsZUYMAWNMesDiPzPgRy/kQyMPm
5gRIF0+6dPEbYk3in5pfV3SToVcFsgVPIUnINoT2zrplhEtAR4FKvOhiPC2hkVyS
ikzfPPW+skGLQ/8woYLM82c2ifx9MN4ban/M3UfS2JvKfdR1UJUMz2/r6q0sEanz
VZZ8bQoKsp47VTcJHazX1AWfknWhKShwX9AxLERLGoJydV/jFx6z1CtrCLuscCkj
asw10zo9VLnTTHA9iv7ITF9lj8fFDnPi/5MUJw799WcEQRq02U8Sf7Xjy3f0dRUb
wHgX9UCVDzYMy0CniHq0nmS+LUusl0OGS4u9UaVwZWq/kQdd5YPWeHSJeuhXxYdg
4s/cutmoRZ++cEyi/ko3T3NY0+ToINsawkSVA8HB8fX3WqzXNfXzsvaqCE2HKbCr
9WvcSgGeGgPO3xh7q2p6RBa8YZSeVl08FyNTlGSuem0QRtVtZ+AhqNUoKJ5I6Je5
iBpVcRd4ZcRHqTxMoFav0reMSYM6J2VxWbSKlDfN5i6Pe0Tf8ZY7vhVaJBy7QDpY
ozDijj9Idv1/ga8YuBqx79axNb2/hENV37uouivNgqG7kcjIuKgWM9IrMk8FtkCn
7yxTb1f+zQxImV6ykI8mToLoGeJ3K2Z+Tegxuc/s4t3Sact+OzcJ19fZbd93mw6p
jBQ9x7AP8Mglmqu3cXfq823nAqn7ElRtB1qUpa0TLqSuniNvB6i2aArrmuEVC80s
L5XpTzoDHlP6PAP42L1NNBl2LEKuc2uDZJW8CgTytn/nta1glo7nmNC3hz4ULMXu
8fgGkb9gcE6updARpQZty4kTngSxp0nR2RKAUq6GJ0b6La6DG7O3z3I67vOogyUe
bNLTW+QEAKThG188LcfWzkZF2P5SK97z2znCObFgAbN0VjPuSRsAUx4A4PDlbili
dc15UGVAzyXV/f43OiXBSnHKBXZns1X6MtvUini6fj6eeVPG9XX9dJJi2wk9qrdf
GFQoU9ULB0ucowheQUoYEiRz34xVrkZubwKNIBA2aCNNcVy8r7iKTFpjujouZ1Fu
9SUzYgAhfYEqB4h/kRk6QNM+SCPFDtK3+uljxNUHEDC274U4dFlhrnE9znkFZ/ut
f9HRoRzZUu9PaB5rLsCtWubmVOPNCRaqxAfCoFivTWPObAuPXr1KebuDLLvo/qFK
2kmdv1SARxwcCtSWtYyt+vdKlcbyactS9zw6dgLRqZGy0c4BOUOvwvyVBsIoi0aQ
JqC9ZCqeJ5Qy689w3TD58qQNtwxif9W9BN6QRc2IFumNV5WovbJOChPcs8lhYPgq
a2qp7rNYMj8vnzvhcqp9iSjR+pQRn9q07FFx89aAjvWjghYVPSvsqh+s6dWVPiLW
5LnbEqpjG1O1aTns6c90SHoPqGfKYpK3iMbu/wu+ThpU2HfroA8iGsiZ0uwLfAfy
kPHEURsV/Xoi/G6+Jl3FhJuie+slUPOkOU6Um12ZsY3vzTZAVntXE9j7iVye7emn
5FYx/KUjtyAR45pk22Msm4Y5P9TWcwIRUspY80VlLe/VLY2Ll+apiOIMs3ZHlSl/
GgPWqyRADHYAxIxa1dW7oqG7k98SA4dsoeLoUIPN51Vu4AJwzxFX6Aljm4hy0VtA
oulMC4vAYKlvDugTGSnQ8Y7z4SGG32YACU2iM88AfHKfARWHIM2pYt1eKXSP5jdf
fT7DTdGl4LNiDd8zPYKMuuvpFbhqebFyyKv7GgA7ZuUs66uYEhbSGx/6YlA2oYiY
xeVrMPFBIj5SYxe3w6OG3dK76Bp8IutxPRhoo8f03+ElROImreIlXqA7jS3TEN3r
1OyC9E7L8lznbM4bPow/HVbm6wjL2hmkLHxT5yGsPPsHNI2fnO2jtXbXvcEnC92h
4Bmg5MCRUaijPtBRYDfE8YPnJoREcGfcqRx7cTc+Pnhr6Gm23vLG0fw1VzyNuRBf
c+tgxKIBNnh0Vj4BsnuURGLe1Y5QdPZZ5EnYPfQUnVFSs/65p+4qmTw5V+x9HZd/
SwpXKHVRsRhY5hYVshgoCBRCiw/hqXcdTQ1PenU5AgNArJQTAY9nrL84EHZbR/lp
JUzQq9J21s5lrImMHa+00Z40MdY8Zr8/SdMy2uVrq+mcq/w0FA8koraSgi9uWZgB
XjhR+iFZujubU/f/U8N2UIHWhDzQbkhgqUuEWeCph91KgP9Nx+KXjUdiqpP0d1Ha
Evkm37ia085FD8rLb9KPlLZdtt0psK9Vtg4gi+1BZ4I+skOxk4Wo7DZo7woYOdrW
oA3nIYiuzQzH/9UBtJChcdDYwYa7fXO+Gv3XKhFVOsaT31y5Q14Ub4ZmZ0ym70ql
OjreyawOxwkD+k98rJlViYTX8x4kbDPcKZK+FZyJ299UB/FjdwVVowmliKANZpbo
q8WswFXUA4Kj6LBnmDi1prFMwpwODsAy5RULzv6oqKLBIkZoX2toFeStTDFoM4yu
uJPvT9ECv6ti/HhZOmPl1F8w/m19khuR9sa4d20z94AruDaB+aXxux/9cYfKwfy2
XACqBHODf+3BjUU9V4JdDyyLAKIMLNodQmiHhQRjykJLA35CiwrJ1yRH7+a1v4sd
ZjUor7c30kMhD5LvXnKn2dDGyH+Q395Bzim9LK44hI/4BHqUxY6H49/NXzjYzzWN
yb1xv0ZFX6VQRe2TMxB02ZpTyE/gNR/3+vpHIU4Wx11o+2B9rStDBf7rxBPmYAaZ
LzmMGmvM1aJS3tfSpGByGjDglqrCHvM+UPAXLvH7uvC4nWY4uLYUMy3J9Q6QSP6X
2Uq2qdtqr6Fxqqku0rPpnyvc0HATQTpNjiqPw2488hWeAkR2oyXdPSCgNS61qZtm
YtxXtLbAuLxrzUu277Shbau+GAc4mMI+7GMV5S2U/ReZqJANqZn/YYtdgifr5A4V
by9GSfdKNaB2RVFv1UGWVZPU6vWlCf5YO4unmYsXpWAxIOB/ir49x2H+3HSWWWJC
5vM2tTdNX7B84YqWqoFxjtvAEIaFT73Wynm6j07CDPh+lwIQVB/F0TjNQ8hHy1Vc
ZHHMCJK380yewIw1U+4p9/QDS/ImcVL80lM3jZX7K2phwvg9eD3tvOWqSwl4Lk6b
IbBHc06/I73Let6rCTWhvRL5/vl3mPV7t1MA8eSe5TIXqn6+AMWJNtdQfi7MpkUB
6PnCzW6ZH/JvNwmZkB6ELbmTVI0L7iNBkO+dzzhPwjK0tbVeLYeZIeutQiIhfeB0
DkEOHAUePwpto7d7/e1rFqRXsviyf0LBaBhDkyiCAFauPs4sGskhrBWi3rSqasNz
IfpsIn4sOBtJrQE0fYdyixT5cQT9QIdxieOnGOeg7L39T38Ugb2APs+CTeF1h44U
UOi1JnOZMFdO8g6dsGyyIfSpw55K4IrNisZZoyP7YThlF2J/zZgrEfJmx9tU1/40
hJfSc4eQA7XYzeV1d7LHqfHCCq9RH27KBoUXP3DgXspQGkw6FaERnWFKZjBi9S7W
Q9HHaDx5u54KQFHw49Yg2mVnYXrPncaGc5PyjFVe5j95xZak0Is4k8nyjv+EW8ie
wgmmuP2awUXCitW5BRAQ7aiGavJ1rEoYnGXGYvavszP++ojs0TRzKXGv+JWLXBPc
Z3T0juxihxP0FlB49J+8mVjjbLsxj3jZ6kOGxNO7OprTG6yAow8f0dtzq6q+Oj57
u+ASwfPJlQURn1wG87tf8WNbXzGAAb/ENOpho8xc5Hs2syKsMosKskMzUpK1FhHi
3xXdy5qq/wzxzHjiLvqabqsdNU9EU6D4o+4+5bgUsDf+seWGFA3FJYOyDG4kX5HW
/N+N6uFneilrE7amCwh3fyHN55uRBdR+fabNCxLGfVzr4+H/nHHcVFOB023emula
UmVqxpTsrB+sRtg0laqrIWKGrQWNLg+nQjRl5gUcqRPc3JIAYPXQgA/Rnh+U1qVO
wpt0V33GlVJvQ+vXJIIXk44KCSSBc1qZZpv/TJE1hH0k1zMfQeAMr4MWcsh596Ir
yUQG7qTRygTHgVND+8qbpIUN8n83eDZQiSYui2EsxkSkJuYxj4Y9TVSzK586ha7X
nK/TREg4cIjkHLRwzqpfbs62QG7DcXISSUGYmV8o2/ohUNwGyjYTP7stSJnWosib
wkpgFLaVjkODnD5S+/QXQA6dNCylqxHwc0y5xzqJSbtpJNr+yW/3t5Jcc+NINEAx
Y7OweeoC73wi1MK3thh0iZxM3bg77dCxcjZ6DHsumvy4on+5VHsj2nl9iZVMAC0a
ONxjrWLeimF2a6Pw0jf1ulLqdVVizc+Fu9rIpYzRfmpTtrlj+eT/QXs9nNdHNDo8
7UUPVJRSoHA2oE+yoTbH3RMZrrd/RzFdZbmKEkiGvi7cGBUcOEHhdn8N7s5sNbBY
PsCABDOdciTRkLPfpkYQFJUmQsdRKY0ZdCgHSdrtX6tcGcVCzigE+5AS75L2eKD9
tnhxNlbkVUrq4/ItSOEqoUSEPB7tX5VCDfeYw96wzRoY18JvBCj/cXd3kyLsheRd
78ScHuA4I3nehoRATNmFU0bRyn+sdzAqTjoxEjoZU14tsowlqYHos0Ja0VsgcWcO
Rd5zMI1WOy6Z8mVuqXKizgN41zC0c3/1M93zukH6TtVALhOJpwmJ3a5JmzXjUecI
iOVrM4TKpS60r1oEOzCW52xRYb+q6xL7cHtvp0CaGNOCB1JC8+7OCbXeCu1ntiuc
PsM4Pu0RjhVaOhbwJmob7rnzFzjufXoyPM1bYf2Q3SWbcuKOTxYYwT+uxaYtXUui
0EfIEY8XSxsF1ew/a/AmKv+/rUXaiwqeaV+oErTTXSoWu7lhn/TPUZGowhP6r5mX
MLWePw441qPB3Eoj8htsQy8pF5J4SQW04pIhlttv+dklN/OF/s5+KCoEimUWX2v0
wejs8jMReIPsHLm2rJLvQMIvDYNQeZ6tyeTWI01SOaimJeOIomEYVvB5xnEzEEQy
KkVmUilewPp0V5daGCfpBNR5gK2H+cK9Wf26FtDTX10vdUVLIGHWttkK0RCy96PY
jaB5m9v+9SjgmX/34poggzs9EzIH1pkYm43kIuwhA3ccpTW8avkabEM3RODngHn8
7viNzWcG+5ORTfZzrId7Z5FQSTxeG/AqGBHaILLVLQBJUuOeFJ5JrjM0BuY91Xm7
AWlXRRT3So+CWC/aBp+J3CY5fvSoBDCjuVUYwOBWlItnFaSg5P+/YecrJi/5VwCD
xTNrV0/8VAn5DmLbTMzGWo1iiImBcnFfKduBXMmhqnWGfIVyDqG6Cvx7NPf9nkTS
DuQxFItEL9A+/yvAipW8tBlAxQyyEuL19dbzYFZn1MnLTODM0O0wK04daEAQ3etK
opTnN3YyCBNPJvvcEgbnAj60c7qX2w+agf6GpLimUB1/9WAQOSh/nIfuY7yMRl2t
EQ0M1Ow8he0RdWKFhwom320UywC6tG5dqGwUlj6CCqdFwd+FUGczN1uimSJVfk/U
cYJSNcvItkIGqzauWNQztlE/D9Kgo+v0gk7vnhHkHqAjPwfCT+m0AcKpUVWvabqO
AM+TQ/ZVC9Rdir/6Ktw91960uz8GbQ1PbMK33Uv1hyf0VoCy4XDPZ7H04fO8tO/2
bCevbp+Q8cIvHaUgaJTjeRU+KhkfrfzgnyK3YTEq3LB7NCsoHwnuwbWmwbqnyj8D
enl4Nyh7/QpuXzey+uxLaPgCF/Wrr342qK8oAdaeHWLcmU2sCTc17B2Uvvw5RRfg
ST5ne/6cq0czef7O3x61Twi40ZHxiV6SUHSGhcVHJWkCn5BPrRcvvWz/6g8fjLIt
1hjwu+mjo+pv5VwXc6uy6XjoySgHvLL528ia4H+zlX2pD1HhBkZbt9nJQr0AaKsU
2twjsZJd455Y15O5ZxcmY0MoBgBwbA842PdeSfdyhfEXRi5CTbkrkH99c0IxPvv3
Op9IdpWVJ2eGPLzFA6Z8qx/HLQLxMwK/uuX0OC4pE8Sv1g8FBHWs1keKD2SWfmPM
9j7VVTIHOugjQD8Yh5c0sybDsf2dr20hw9EIkMlzItBzaTo/vQhCTHlFkdOIeg9r
D281o+Eyr2fNf3Ax7oWDXVnTOz62aaydCY7P79v7ChXT1tJ34HD1cAUyAamtl/yw
70Zz/IeKCfaEkTlOgmXjKGjI8oXvFod12A7sYZy8bAZZVZ1NJYbh4hedws28/Z+A
2HkBwNMS5XfJQyYUNxkqF7rg+h5HQVHbJ0BzJEYW3OyxM7d5hT8TnplutCWFycHx
zHgvrg+U/OjGcEOHFhX+MjiVnKzII5tSe7jUFEcI2+dbKwgND9zKEMVLru8ikCZP
DovouP5FepW3bZvHU1c0YEFHxhigAUtWm3nQbkYiH5Qvd+L3ptsGEChbMKOBzgJb
z7ulYOlyNhnRTU6iV3wzeleOLWJhJ/HqbaBRPG2xzCxZGFsih6uYDh3y6hYbWg/y
4YXmpUv3j0PqI8yIE1QnFQgpnGxCqQm7Aa3vuOzEwTAa2AlxtkpynuE1OVYDpl8y
5VHKIXNz8/kIytHVcFb5zYleMZZl7qt+eCfSdE0N+DQhZ8UWFy5Jitb2FJv3FCVC
2+jL7lJ6+LqVwpEht4TYSdXyH/l6OKjvurXTIXZUx3ROJZptDhgqDJeQeHyd2IPW
M2zV2tpQnR6NihtsR3/woTFnP8DreGjiKDFwhRWknrXf7VTnykuGMeg8/9HAKtTR
1PLoK6iRLTfUQuLLvCWbyjX42aqUveQtAMjczm2TtgsD2g5RnbyN6s6k1vE1CFWq
KVymHFSovpVwgcdYeF5FIXemX3RZPJlbbLJdTkJjeoN+9qTDSw5iITF8OLN5eC/M
oYcQrx+Go9dhvmZcUfXxQq1PN5+aFSn4VDlFUSZjizMiQe1xdSwoA8uf3Ctc/wSZ
cG9RCPb7VS0W6mkhd+G3s8DNzlILtML96jCNJJsJEPgYJ5Nei34/JRaYF5TYf+Ik
k8MIwsWPH0GiCzlZEbfi0N7b7ehY/IJo6fdfxr0wvFOfN5IwrNEq0DMhhzNstImg
tizWiRR0YK19ZlDBIWXCQGDD/z6zA8gqwNVGFRyTvlxpbLuftl104tVwbvslRQzY
jho56fnBb4R1OPVwdZnLj1P2LqmfTO03odmv68FPUJy1/uui+0DzM9Zy5JLZwapY
4it4kRa7EcHnEGTjySyMzbiQAQhcFAC4XJKaimo8kZDBgjoz8DV6dgAfpqfFHSuF
ze22GyFC0as1KsNzrhZKS/nYCrIOYXoPxjo6pgUUE0VBR3VUu99qD6ZNTikwXq3q
KWkr+/CESdJ5NzN9xNgdFMoHhMfOZEKnsccPfbrKk7aWZBM0jSHeswu80qFEFxFg
ITCFBL4Y10lqv8XeyS62EcHfHa8ZYh6M74bbt8Pgd2WMB8TQ3Hftjg2NQrPMsl84
OKOUGae6GVOMHlM4PnfWTuP/ReQsg2KrL0UeI02Ddzi6xAfgIwbqVuEMfQ80ag4M
gOsT0j4tgBIXg0nRpRYN6AwZDvmz13xEEe4HQFBZAjEyEWqLZFa/mC87PxMgjKjj
18H+ZjI+SAwLG+X79pjHmCXaoL6yZt0Qb7fdc+cElviHc0o/jW3YvDIUnu3jL0n3
EGI9E/uS//0tZoIOYeydluVPKB+z6m6+89qnnW58sqwKVxkuS3fUppg5bHacm4dX
sT5uUmMU9zAC6i5E0W0/X4+H0CdqB+Jual2T8X+GcgcvumYe3JMBUXnDQ1TKJ1JV
ZEEkelW0qdgq797dwF3A7wOLlERD3OkgJ4s//3/6l6R4Kh13UaqwD/F9P917aLaq
biD/3eOGZv109LXhY/mXU7OsoOh4RR3/ogNxfMfYbdH0AyXf6J7/kIxjh0P4btVt
sYh75yGgkzFy6yocoY5pnF8FNwweZidLkYhMMd96h75fstJbOa1JfdeV0o1JLpAV
O/tXB5s8iH6xBnWDxNLirw5RGKT0w+fAZgJv5CPe8USDaTFCj35Fbi88ok554WzY
L49muW7qO1LGR46lv6Mp0bHKThCwQ9pgjx8jqZ6sgUZmqci5OJrqv5OSBz/eunwk
YcLEmfPjq081pmF5Bhmrwd+NtZomAp7qhnV3NQVsyFt4khPswsKBoWpakGZvtT9Z
AcPYRX7PftWpLXu/6KzMMWkgXy+BDj18lpr+RV+IR2msXGCUZTDlR4fy/uYxXHu3
U0/Fv+bmtmyPYgakTrvSDVxUzng7OUeIJ/X/A6JjejZAF5PD/Nf0R3E+5tfaHRQG
bNUxZSw0KsvvFhdjm2rruOwDTIZ63GAtloTOAAC/A9gHBTtO5hUY2hMD8LwuQD3j
JATjTGgoZOGw6bWKNp+fP6wCr72ng5gFWZF4YrMPjRTX1qlCpabp2T7c9c+/r1NJ
yPCJeUrKE1WS/9pqcozXaG6s7vLgPTiCfcPAc2BD0/4D5SbQHOKsUTfRWbhkAguV
IyvoxreMsP6Jsiq/VLuxOMUrvs8PDbBAVUYzMOJ5m2aQipMyMlecjXNYzxqzJnHK
7V0iyIDrjW6hU5yYAVxtG8ubSolFhUr+bQCuUhXenyuu4oVuFXmcNrjCKVvpXXyf
os5dRPQ0Wz3ErggUKFCbxC1+Pf6EVW2L9R/ijUcqhs19f30YVEtyQiAfPHaaVaiR
pnZkeiZV1vFBDDnccxLxrECcMaZlnja4+6giGDT5+hHY7NizLx+LS/tvroj8+YeJ
mmMTgnmaUipItrAwpsCkWEUNOjHy5rT8c95hmECkBo+gq0ArSP24NgH+vRkkXwDp
jASFEZ8DEugKxuaQVZdH9gk7EAUIBBOX/iVTHmTW4VUYE9PBudI95MYhfVymdKXJ
adVZJbrSWDftNUqKTLs9Ji1n/0nONDmBNdXx9dwSnkhb7LVRwXFJTdNVtM6u7M6E
LjcKp58YrXC7Cza+Thrk1QxoAcOS2Ekw6Lfl27MsqV3FPlvvMClHO2Hfy9C2+uPE
rSGR7Eq8sKMH9jTGxYD3ouL9qqYt3ceD7WcBZHh/MOcpVJUIOC91WxN44ep1FFrG
I+qrgzEWdCBWhRoAj3l9evC2bz/xF2913E+aYYpn/l6qD1MAsIgfUtAU0pBoC/oA
4j+gr8kwH+Sg2Lz0FpZBWkErktaOoBk11xrSmvAi7P1KCT5U4XJ5UPcXLfLjDoGy
JPBwPI7vLDmkK2b5Nj7JadCkmZ9mtlsboNc9j7BueuEGAFdWvdxB34tlnNCt//xO
RBzR/6wfs0cp6JHEfbpwzXClr9v+Fhk61qm0gTUE21dPp3TQcwGEmyacQZIBaV+z
DxfAnyJUJFVfmYALjMy9lQXdZarBHj3PXheplWnl0fUxtirQxe7InSECBS4S6Sea
9iOQAyZ98EPiHcixV4AU4Whh8SI+VX1fJnAxO/jjzi7yB1QmDVl+PZEBDxCI7/4W
dq/px71Lu1Dk/R5pqWNGzeo7kG1Y9+4GxUqqRVir9MaE7jeYrO9eApzQu8tpLJGo
f+XykHnUquqzc4ePsQtzyFQTW6fICXbMA3RmK8Pu5DwDydi0YuoGDsoH27dM/Q3F
2MnvvzNlW9B6sbKgmtgleTbcuqNh5PisgtOFOjNJBLVFczz6h3eXRBenWz9+HjK8
voiac7kxJZaN2RznRpsEWcKozlULbsWt+iuYo9fJTjfah6LoqnAjSEMtrt2IRRJO
GQRDwyZ/581id1fm1ciOxSGxaThte+79Liu9q8sHNBzjZ8TFGois54C7TxeBSkxQ
NctjOYNX/yM9cPE8U4Ot9U6pZZFd+Zcx2hKzVUcFzi5YCodlzv7S4erAFdsNKEMk
JK7dmFfsCpxxNRa+ZmJKe1rpt3PvFv7ECRJ2koURsdn9dYs7si/EiM9/pTf1vpPQ
Ay2Fd+nhrJChY8MMS9CUD2VijrgenhLiR33hbT5CJe5RjHmoxnY+lOuKwAP5jg3F
G2g7Jwv8E34lkJcsB/ms+jftPIm9wqCjdea87xKgK2NUwJ6McYguit3wD5uEbDY7
Ok5t8qWD79MVksbRE0FIIKXrWuDKrNBlfdvRmdUK5hC/tAUw1PKR5y+SxK5vcZIQ
gNbIbgQUEnbaq6kfgJO6pA1TPZXrF460sNFiolMa6gG18Vy0oowrjouGypJxgEia
ombn5sEMOHpqqXcnKXjkhOeCqiTJOzlxsye2f4UKw+qMDCPNCisP8o47Z5oUxD4U
zjlUgle0+JwLrg35kMQn0ApnXSOYEiBNuaAx1uaMs1sjLcLSZQ4Rqt449GrmSUDK
b48wy1vwj8UcknpXu7/WbAt09hmb6FIa/LBUssp69QfFIyMZ+kEZwLj+JpuL3Pud
9v3zkKfEkc2Uopz5y7bag3ktOukUQCYIe2H3hkrP+m+JHUl+MT/JEPhKYQqCn9yH
aczDS/cP6KnpWpXz+tK0yJTz9mKHkyG7HfjMjWEMNJXtzBUJ2RwqZCaWbL9s2B7i
Q+6+Jj6evkvUiZEd7OxiLd4GULb1Yv6hqVyGgZwLmjlsOV6p1AKou2XAeIuKyTlN
oyWMYYfks5h8gWdFgPDIL+pbnOMF0gz0yZPtXftiA73hKIU0QcY4LTkdBBEfVugB
neVIf0HMeyyObsDlaHBO3fw5ouLpmbyX3No/W2eWnFzourZmcvfC7oZkWQbbD0bx
fHWjhQlHybNRpdOH4xSuBHSCxA8JBpgbTrkv83X32N3IcJG4pgJflxp6o6l4ICDk
AyiKnO5+4u4L4RtjLFMZsUfrxdVSfnQOS80L2tk0uPbh1D6R/9dp/FqMkdIkRRFk
C+PuzsEu/i8wlQYZml7VYUlFRVrnUpDKWVhtj5IxXRdjR4v2mxGWuONGjvKND0j1
w5QCmjKYS/QWFJXaC3SOCd25BA6nb6WyxFj+FtVp4gV8SrAxLkP4DUVcIZoMBLiS
b9AqpuVVo8M01drYIiqnaeoapuC3/jxsFr+XwfRTDxsQ0Sl2beznxw2fkwQ48HcT
E0/8UtCXYHMEbvbBfKNhxCbdo3arubU2wz5nnNBGrcxWAx78egBmhZtdN+gVkx3f
+IAj1zHvLA9pEHVJQS7R/KXzTfJlRkvO27Qi2rc+pDOWvxe8QC74N5KsoADAg/mL
UKRsnl/mI0aATGPi0MUXrR/WLA4i29EDlKpSEXsgzqkmNfmsZzXT6PhW2sB46VnK
gG0logNKQhkVPrz5aqoZCsSMg166y1UmHk9JgFMjuNfxDej9iM2Jp0SkzRiuXay4
flJfE2FLSyyTD3qErRFVViWMZXXWroe3wAIVmXrXDdhMHJkh3wvZxTfjrDtH1hVK
j2PwSxCKL+US6ra+H/rCUxCBFOmknRWqSRL/yqj6MJu4QLmsDuCEjB8nsntfwjdn
Rgw2K2iPJTbzdShE1Ap2BFLZRnpUEEytcXZu3CFyAc+LNotxgpyFOKnLWd2nrKHr
ukIyBCyV3wTn/keGt/oIY0QqOSu2srVr6+eszk2mvQ/tCDN3hpbGBNX3fTTLJS2k
HtKRq7J7X7A32vSdTiTVyv1TF1+/P+/aV8YA3Z5M+CiTcwRtSTaM4sHQp0w5xq7e
50tbK6gE3rA2FlY8Fn0KlF5OaJnaB2bFQXG723z9oILr6IpbodS4qSwRVIkto7XM
CmZp5ex7GnWvjbZAlS8FwZib2QeFjhtr8zgFtYazv6tZckc++z8Q1Uh5nuIjRK2s
L40pBz6q3pMT4QZv246iwrngXFEI/0smYZlhUkRIZ29rZo6q7wusx5CBADApqxhH
/FV9JLbI3vdV2niUuVLkGcqyK6RUcqcAvuxWUevXvCZyGG9hGFxJRmVEzinr1GJR
d3kuvi4S5jb9z4aHjXk0KE27nduCtxrYD7ucDbLUJfwuBAbcDEfhTmJmrNU9EZz8
i3UQSMCnJ4Tcdd/MIqvMow==
`protect END_PROTECTED
