`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Snsj+nxaro7Ggd1CCpMedzLtmZxyjpE+fRN9XvyzoqHzJB7rSDHFHhDyPe6OPN4E
ICGsDdOv73hdA+F3zI4Y8iktePpA1v63lpsEkjoEJscZtomnDljZh64eVN17XlJv
QerDX4yFVDnGWpqjEu5GFVHOdOS03SzIjqZeMrg+Va61wbBs9Ljz6G/efx3p/LLU
qdWTi8HbovbUgRorurFOT/b+UOuOJKQkZy/F9RyO4quE0V+7Z4xb5dn0gcmYCEwu
rTBTgVcxFE3GB9rAWEjTkHUggXWLzfIf+E3QhJnWLpTo+SY+hrlcSKMWThHCallN
d/nOAddXr7atQOeqIElhpTtVpMtzFmXIUW1RDIGJTpPIzgYI5W8CUk4w3D6ouS1/
+aR8LxU6GjdA2xeQLPzGB8HFmhGnhNwymQfVfxJKJ22zScFXP7Hg7SEzy4Ut7+Hd
IIb/1pGTJMZiaWmjVIzDAeElW8UCOk168FUrb/KjBWMBioqlF75YqpU6tPk4+6Pp
AtzTyGP/SmcQRCFUdh9KacPmytvxk6wP5frzw+KVnRNaF7xUwaBwCqaV8zhL1iWW
Dm5DsfFQ+FnHWUcYHrdHi3WYAnh0gaKnb3+MlVS42guKyoem7xhMr+HV79cNop00
Oi/HE4kWM5sUV3jmSLmQ/hJGFUZSXILzA8R/7r74LQgxXCyQLkhp1qRYjVMGKq0i
5oGXXVa3sEifxfgsvSzG6Jt85LbLLBiYSDUb991t0ee1qk091Xl4cgt+kTIqTCOI
`protect END_PROTECTED
