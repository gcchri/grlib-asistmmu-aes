`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lF6UznJI6DViNQXlwUgzckQ6MktaiXmoUIXUwTkCVPv5dRbBXSLUdlWAR03/tomB
bkqtAkkcJZI8h5YPhdGlWS/1qZBi1nIRPsbsfalOuQvU1pNL/csC+7V2l1MphR+w
rPx1EeEt8+7R3e+dvuVA5x/PZ6wBTzd70EgmXmpuF5y8MuX7Vm2AhNLHYBusTiRH
FHdJi11oRJbYZpO210oyiaVFZR/uPpdJXGfjFfOjiDVa0+i6GX5wnSBJIMIiZMFA
CqfUC8ImJw74g3sgFhlwqenknePe7PYm2b83/HYdGhPIg4IGFLQkV06Bvit7cSNN
ksoLZGX53QwYsjgUwd/m9rMpC9Rm8lEOzxj0F9SU1JfYP9tGbc4ysYEBMvMyQ1iW
w/HMLxe0FAp6zrK4vCEapymPE0XMIeg1rk+JcJzRvMdzPyKWG3Ico0kt6ts+2dhP
xx+K9y8V3Cvl8ys/lIiOb8cjp66f9bjIRsJl/U9t7oBNdE9iy2+sLi1bbD0SlC/D
oZRq1Yq6d0ksVri7azme0N5JEDB2C9yrUlor4R8qxDh2N1dq59SYVfFpvKSLcU5t
`protect END_PROTECTED
