`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TDImxLJIASS/Azy8kt9l1g+ITuL/q4y6mT1U5yX3NxW40G/0dRB8OGv+0IBkl2ac
JQ2sCQTSEfT2CXNVsVVrwAyZQVxLBwJA9gF23uOUyQ/tly5dUUau1K7M8guduBge
MCPWi4fRG7+r+UvhOG7VXaCwjwqvIoWF7ytCNPJ9aL+0rwwswCReDzZHuVwY+D/O
XdZdbMzJzLHx02szto7H1xUlHSNRBkbCEHb13/jfHaRkoAPl/R9RTdmkGoVxLtlt
IXWMRR0putRMLKH69WHdkyKZmziQsjiejP3teGtzAOmdyQL35bL6UXZxNE0hory7
o8VX87eyQt+ET+yeb2LNXw==
`protect END_PROTECTED
