`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
woj1+2mEwi7/UUBlUZ3GO6hmwy73uRUFqvpMZUTPM6uW/i5/3SLgkTzuL8jfAKvt
fC1U9GB3Sx1+LhUG8jlMy3t1eN++Zs+qPfihF8FI5X0iTj/pz4DDMyVlXIIbN0lT
0c1q3VH1ep34+9gNSjJxXmIHUUWLTkkJkSNGBisPKZPRO/U+8VDiYFiI1f+sFcfd
uAaYdu/U4wxYuvaRSaKZz+4Ig2C+WflgXR4BxpF4rcnKJdqfIJ85E6z2vGNK3/mS
uWjBsTL8ozA/zpkGwUhBUmdbbzT1c2B4anmXRg4Bld8=
`protect END_PROTECTED
