`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pBrNthHsSa+X8In3uKz7nVTmNZAviFKN0pUXHeuy6ub6FtSSgy2JVXHpvpz7YmBr
EWm9Lh92BtQ3NuO8SRfGsfcNOtgjssmcIe70M37HaT1ZTTbDj2ZFK7TeS/qzNtSv
c16S2dv23hH8mHdJUt4Xr2aK+fLHD4kZ56sGT2ukWLHORA02IBSbu8SmJt3trjPn
Se9Cr92yt+Pqmz+3hTP770Y6mCcjymoAeHqOpl0Jv+e9BMZJ3WU57MjT9nmOhJiY
TFXiM0uqkXP/cCsZz/xkQZZ80HdoqSrLTn0nT0mxVtvs0XotTxt0Zc+pKdxk40HS
nIUIel2QcRKyxnsfIh+x4lm2dAft5xV9zjAMdTic0w+lkxqkU2p682GwgQbqZYEG
jstpoBEDZGzLwNOD087y9BsCsaumUgG6IyoesRSNAUP/oZ8CQSbRr3mVsrtaqXEQ
kQBSMysKvsfdbn84CFWb+o1Mdt9PDmZ/GyxwGUjqIzPT7LfcLDCPB3n4crmvJR1L
C8Hf1D5nbzMYsHjjxxyZvbHzdPjHsngVoReZZ58v2/J4yreyLhpkfgSeRUNQZT8e
Y7prpDwBXYkdHJzSWETW4QZ/+xCAbTL+ryPLTJfzRUVKpngpDdum5iT9Bkm6HB3h
3Ymw4rjLkXvm3y1k3M7Oh2pLy+wLd3lPFPWXDlMtoxRfH9OrAr0LltQGF/L1Y58N
fT87gUdKrtWtmNwHrzQCtX7CKEt1i2VJ6QPgvoYSy60mxuEDeiSBHXd1MNUoCtA2
coSuVj7XoMg3pWFZebOmj5ogH2gojvgY1BU5wsrYFENywFYRZglOPvgzYyLcmfDb
9vBBhCFV3BSh3rM2HHel6+Mr4OB2FX49+U0LKhOD/uvfTK8RhlKylJSDx+OKFP7v
eRwds+TQ/EQhziq0vm3C2SYg2fUF0Gan4zskxw1uY6HoWxISan4/waDde0985mmC
9oG0efjFOCFYgGCVEnT0yNabuPTww8Exsz5D1bxdbk1ef7UipBOLZkHTOvqi+iRL
9qMJ966/Ps4utKrQGDD0dglKwNH1Inp8TdreR5OrIumLLb3/0rztLID61onSIjHN
NDOgMbw9A2tdp6zjKO2FKd0atACaDfTnMyq5POmUj7qa6wiB4EcJhcZjvpgHRfni
hxkd1/9IBeL8Ltqwf61Fz4mz4NcRH6+FckUI921/Mb5O12aBGZMcF0WxBe62wrfu
MLaPS+zJBxOjIfwdDDyU8jOPUExQDCmvUWd1Jrkz4IZHJ3pIHw42oLsGraZxE5gy
fGTRv/Gfvmvxcc8llsnl0h1NxglmeiQ+s/zDeY4lmUvTpMFxGpjesSCq4PnmwgHD
FswhSMlxQdUB5uiYWijOBNdel21zuJTT8Upcf5LOZtjcsvzIZBTzJ+JA8GIwk76/
7eR4vekKAx7DP/YeoRL5xeQ/LID9BnNh8j42/Zn89dTmglh5c1oFU6NbKS4Swk+Z
WP4/2bZJ8GkOYJWKIVDBPrpUzfI9oT9L2sUwDWkK4gxbJCLuAdvrTqugG4TFeFf2
1ZhTQ890wd6XNr5V0mSd+VS5v6WCtjCo5ZkEUzc+pw2uNyiZ2NL8Qrvd5Ff8C2lb
zQWVfZDGPMxUxAKn+R4GE8Grjg0r9wqE7ZwiVF+ixGR8JyPzYMabAEWnKirXUBiX
oYyM0ojaoYialta7xSwdAZG8bd0xWNitsivDH1kJKa4CrleHmV9DzkAmx7vFqh0v
vwsTWTcfIas0auKzl1aXYXwAnHYycI2NTJwWSFqTyf0X6s7p1+8sBEyPtPkfWfOw
zQIn8xYeMIm/u7fv8Fv2Wd75Sd5NFkE2Nhpcjyi5bPsEqPBEtUyT2s9kWfTVZ+Sy
40fTeO2TGwmNbb+iEHFQS7TR7TBm9E2zMA9r863C7yHjAMCAAFntuXB17SJJXncq
qTIyWuPmBvO5Q1xqYIVRxI1SFbCWSzws8/8mFm4ct8ygjiyzP0zlsJYfgv/vxM4K
/oA6KXsXkeeT6VDFnTO/jdlBjpSp4ngXoOWz6fy9v+6a9mWG/5hpddOZ+2xX8U6i
8fvP/+F+6UVj/6BuhT5LZKLqXeg/IB0dY2hUZVQYDyy3aNxxEG5qcLgPRE8gyaZ2
EFUanUSY6qZPCGsc8yXtWYuY5NV1bnue1XEaSBAE8vZ21c6U74MPoCZ+4ii2tavw
N8iKCaRnc7YmqIGgxa92rQrrZd+LOZBaStFRo4/k9cU9KMbGqeWqQFxRSQT71Nwe
dhdyWYI4qmZqjIG0iC5WDv47tWIGYBcMLjCXHDP0p6WMyHenXI36CBsEZ+vlzFDF
kTg8KhM/PujEU8VE0lPzPWQZ51GOWD8Z7VQsvGinAl92B6iFaf1GazDfLWKsv1wi
TGgd4seHiW7GnhM4PDCN1KYOF0aIbqFWyPEGIbciHiC+XH/wo5J+B/Ru7fEHEuqC
As7t7xHz4Ju0OVEFTOKrH646VYKyhSARFh8PsrY0cRHMYwuG84J8+CnBORRrvurq
Xsrzq4Jsh6uYMWp9ki7nc/aMy5ReF5JKYuASBhLrw1RKX0bVwQnzNtKnxxK+s89V
uVp3lULfQgpkG6NFA6QmqMDts5B2/PcGr7rEsQnkbadgzPj5jF5I6Ii39cVz6lhb
N4KL9UC1HktWLtPMml1C+CM3iLrNExkO//6FlourZaZQ+jAY/ws3EbJCeOdhqnng
Dl9PiXjKA5JHhOlXpVP+qc+YB/5n+Yze0aV4O3BhkkXoHMufekNdaIUjhYnxusjd
rFkEepi2i6eI3fudobJYGljMhjjN+HftYltT5urxhVBP7jp7uvZDWnw0VZXxFnYV
Jfw6/mc2UhBDKaS/AN+Z5qu3Wlirr5tipqmHKlJCaooOK3+D+iu7UfpRgCaGDNZ1
4nQEnwbaEv9ttl/KljPtN4UV1M9+K1MEwX6QTr2UTF/Kyp/pznLrCL+czitrDPBh
YlDCpUvYbLTZ5bTiICU7Wk6d+gJWQoGKXtsx6jP0vG6QOmkTDiF/s6025dMZQfjr
Fc4x+qZA9pndiY2zmIukHrQz7ELeHZKfa/BXyRomSDcAmbHc6d0+WDXg1LUEAtRW
5eephGrjtNPYcyQcCVdUyj2jhSZIOQ+6+JkZgEY5K9koJJNVfclaF/eI0o6NtlF7
mvRAWC+9vtkcuCi8ANfhSHyReLF3soz3cCmPE1Ne+MeCiRjsG+ehDhBVLVoSPQYn
tl4QvbdkPZYnEvdhTOPhoEv3ISV84I9Om4/JF/lPwCYZxtJBd8gz2WnpLAlL/l8e
eh/eZG8lUJgyZDWMqDnHcx+g0h5UHBTDLw9oqVmmFD0WEi07wGTvMrn0p2IUHzK8
5d3WQasrv7RDDTh8hSNr/Jh9MP247nmuI4F9KfDEPDNMX7ajslru0kxGt7H9dmyv
SOm/h+fIrBTSuo8Ou4Jjgq8XdFI2qT6rQ1iis8PT6GeiJy4sbtMdK42kMvALn1rb
TGSt7rf6OE0giAzACsQow+XqkfhPXSfra3XzFuzrDDWHDvg55NZhecgncsVt6SV/
7jUXl6oBwayToNdodFaBuu8Go/+J2eBgLzAhG7+QekEWQK6n9InsZvaMI9Tzf7s+
+OT48f0yBk0+2fyJti4V4+UWwD3a1wtbatgOf/8I0TGiDdR0uVwrA2/AhMC9NpuL
`protect END_PROTECTED
