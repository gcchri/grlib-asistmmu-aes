`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tCi7UqRNP56pgZm0KP6kNceBrPoD2FQPiTDfQvd40UjoMG8dhC+CgKv7SZjnyig5
RpEt79KiGHzURJOEh5LqqJcI+dwYqkqejGtRy28lpRhw2337blvM9DmGBEUSfuHg
dLThEq1fjibZl/+J8iOANzQm/zzpvMAB0JoXHiU0N98KNTaVrCS73skAKpiEYD84
J6ec3cN+CX8AYfJj6wfh9R2bFMh1EGR6vRGMQgNI1ra/GSpBgh83SfSwaOZQYmFN
Rra53D4siE+/QvMWZK+thzKXyhdMD5iSUAc5fypjyaqLs2ysPDjM3iK8k3WjaOWM
41IWeG3xvvx5IfVyvX9+AA==
`protect END_PROTECTED
