`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AJgVHb3thwthl6spIknTATuLFPGHu1Ssz3UUi+eGg4kuBe4c+zbxOkkEHIxMgxV2
7PYDtOdvCPY9LCMvYJj6fQdc3iLSxd/vsq+mIuT3osJk1om0RIHYmR8DSEPqAY7r
HAf9n7rv2Qu5T58fYqwCrC5Sln+5RJQ/OI4b+rnaH5eSRJkmx4L9pUCjXWzQglu3
ZVkK9Z6beL8KKH1hnBNLZaVw+N+Ke5U9tNp2bFitdbZgXUrAizrxEcJjI4IkYmjB
vD9VX8WrXtXWfNRgZoH/1JOL3DHOojooDIMAgyPi1QIS6+XrsskTgk/SsfagT8/t
PB1yvnent5BgCBGMuKnLDdYWQ4T5reeGJZF6vpI2erums5Q/WqzkFHNPg9DuD8HL
UCZLJ7v2xDDH2Fhqg+55lYGUd5M0v60Hr3YPUpK9RP0HuVHF586aNJ8K1MGWZMjO
xAdt+rUqorNBiTCJxOwgTNO/OziELICCzQcIBJxW8pM=
`protect END_PROTECTED
