`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W9vRYO6nikjCyHxrR1wnjp+tnxLH57IAeG3e/xbLdHv3rm5pKB2AJoAqhiVTog5G
SJEmaxU0UI5NuI6bnFbrdl8Xa4vmlaFLcds46n5GPPJ/WyeBN8AkjRyv7bBMTYVt
znMXQsl0ghS145F6lWsTaqFn86rBFjqLe41P6vz3BBceFjMdJN8NnTSEvs03zT6v
HDcs3UlhIp5z8K1TZgU9R1b0tm+XUQa+nf2Fs2jQLl177ecdld/D/KNCxtS+Ze9w
lHskDIC9woO4pOPhs9Kfp/jM+KURCj2e2qRaqiffAlm+kq1LCkqnN2fxuJ+Ng6xc
UdLY89ln/3wt0Nz29XHrn6YbrKEtrnxDh1Zqjd5CK5cqNUGuHLCoCibGDJe19Ous
DMLfkE3o07rmed0/cKCVIY61gs7G0jxi5T2hFkSJkTFI7yy2Zd94Ts/8z8hbvwnd
daP4OSKnpLX7LlOjRNSDEc4Hf/nRll+M3scPNgiuFKygy6Ii/1PooqBogt+IeARL
o+iF10uyiFy0o5mvMXQYwxjFn/Y/NjU+KrB1UleGXcXn9hmxkF2cqkrm2BZdCZIx
`protect END_PROTECTED
