`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
srilpMAIWS4pIlYY9iNghJwOTuI4sKIprT9ciCujAnGJ6YIgzAT3rQhJLQsAhOnG
TOn8iFpGAaQPB6BSbjA5DK3/eycRIxmiIS5yGrUFhB8vmDRrc1Dpi0b1Znyrpmmg
+OFRTXVSx6zTCoPLPRKbz8JM6Pu7OyRc7gOZjQkxfYuBqSUPioDul2ID9BIPvGWa
UANw0vGUvPxhT7Im7/l+O1dM/IESnj0nJ9Y0B3Gq2IpphJQgwJw25ws5H43w2QRE
TalHMk/iel2MX6/VXYPq9shJoV01oM9bWJ79Su0MUI92bMTsHgw8e4WQmWEjVaZm
kWNaqGKyNU43o1HfqQZLtjA9Bo7bgWKOGu2cZbpW8olTvcsxUrpnQklOn51CVXDH
Ss9V2fOyONFNbM1CV4s1UwwxyEgM2pB+x1PCfsQshEZEaTUsWu66NNtEp3Bb6gX1
Ki2p57IBr7VcOrF5IHDMuaIZLUeNG6ejWws50aKxBIIHY/r1ZdZ2JRM4NpWlePOa
2WYOqFi4vxoVmbWGRgl6241UAsfyDgyFQZurk3JGGj/1AlsUStaE4CrqYJzBXUCd
`protect END_PROTECTED
