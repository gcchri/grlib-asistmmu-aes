`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zIdsYs+MwRGKQBspo8jexWiml8n+gaVKmIhcVTfZ9zL96GKBG5ZpAQt7VKHXP3vJ
EneQFjcATXX7p+qGT/HmbYSGOURJOFm2/ynP60KiOJ+xg/zyP25qGATED5WB3/5R
C0ttfA2uJipatU81nM1IJ1yIkLsQKmPlsWtuh9/tAaAhMFqB/Dks74z16AE6ktJt
984c1urLSL4AUAIdSe/EeI4lhsMDG2Atw5zxm5DGX/acCprajsMRPLoqoN+6pbT8
BOA/hK1iXM4L3sr2Q+aGOHKTDcI/jZQg6H+2Tqsl+rE=
`protect END_PROTECTED
