`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/+XSkxIyy5UZjJEyUpbBjsz8O/ELmMcX0j+jpwGLcPVkhL0LXNNsGYi5HIYhIzid
Vf0lVbQrGPHQWMAtL7rdwLeiX/5whjZOFY5bKiYIUKR8SLOK6Pf7ZZOP6mpZVLTl
r8duh1skIRWoAfI4x4DVKVCh556jJ4UXA+bNE1/Mq9TQ6p4bq3HWUtKVbSm/EM0B
+HW2hqCVW0OOX7TOKCMxUFFOv0wWtar0subBAksSOYl31grLt9CqZZwOrogDlhRj
IBwlK+9+yqLoNGf1dK6oshTviNLFslZbUZAWSVpNqUT2wemw8eESpgQi/Uj8DfSY
vhyV7aYKd7JBe/PLpM10dzD+tjG/gN8yabCHQMmMiHOh/UQ8CW8NlaMCuLLAISIQ
2FxO4YWQwlwWgMVdas98kw==
`protect END_PROTECTED
