`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QxCj3BmAaobqzpeVHvSQ/DKgodCX3HzNTz57nTtZn3jJLPdVQYrjtyHOztcwIC6R
J/fcP+0fNf/uk5k30UWtIn3ReAikgZxw2qRdTppfsQ/Jn5j3/9fzxPaN1XfbACT4
nwf20RycblOtNEujCYhONMHczmLus6E2pDw0BKJR8eulTV6x6JYXT0+wv0lM28QW
7Wp9NrLrgXMt1kH88T8DserSdosvXmPS2ZDP1Yd6qgQf47Jdm8TGlcn8gF1inhAA
GbgeIW54cF4xvRN66jE6gUf5U5VEW0IwgDg129FQONVLHffwygzO/8L+UQIys10d
xkRXfG6B0Ly884VB5DUIX9uED7AgD/aXut+XPGlmAphBhzMjRsIjNtX1w/VG0ma5
L22e/YGu6UYol8kOEFyDxWAfF5oJCxvIQdKvjVbxsRonhhQ7IRb4mjUYqVY6it8I
eIkb66L6ZzJ8mLMfv2FrTziKUwE8DJfuh6/HqoG/A3Q=
`protect END_PROTECTED
