`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a2EZG3zJ6o3DWZYoSrQEB4lVw+0PbKKhhx7ZjK5ga6clkHI4JcXpHsqYqGaNDAOo
PYL7extdfTAgBjlfNWHhvYFPvCAC7SdHVzz8oBRX8eXPadHTclDqKfNg/sCKD1MS
ObDwPl6T5ASD/InXjdH7tnIxTGoJ4T+KNjfe1Lh2m1+ue+FqCjdTImusZHucwIYu
1Lmp+5kxzVrUfZQT4P6MWCmwvAs3LbUhUELBp8UBoMb8FpeuDCy2xvQOK5tsNNwh
WxIWVmQz/LDAcQbAw32BfJXDafbulu4DkH6FZH1aaPGQCS2BgJEJ8i1YKi/VzC0H
W8zjH5qAm96PBSOa0NGfDhtEB/JthM6g6Cs5j8UEvmawt4mtCM4jrTbCzpyNl/hK
MHvBNDFZTRR0yB2N8VnpysIbmZzW4D523MQMG9kzXyuJ7TXw5URBfyNnEZFqUIGh
7n9I5FuI6zD3gK3iEQg/B084l4rGd0hv36237KxtGTxUAVVzal4Egyo0kmf5Zmc9
aKw9jBEt0dSu4zz0GOnPX0FmnQP4dYvJqRRT0R3d7i74beCJasJWVIwA2ZM2aFVN
ab4RGIGGs/O0UkMXj8gneP4o7vivCmUPlXicMJwFqt+DIMjnson8P6qjoQmUr9Bc
`protect END_PROTECTED
