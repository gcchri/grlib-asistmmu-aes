`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Foee96Z8r4+rtAev40gPiiYNePEdhJA+hXkYf3MJLNGAfN0xrlrYb7xd4qGbB5A3
X/UL+v9OGtYlNgAwQ9IzG4NEywRC3g9WANCpq26Az/uuH4ZxKYZvSmjxuycz6h7I
7c3DY84w/H1ZaauZdRUpESpsOhiYcYC9lt9jwK5jKGhV+lADHoudQwgIVux/n2bp
+AgwjM2YZnowdm1Wm5h/R/pq47HmZNbsHJTwViXhN0R2i4rQxuGRAcXGdDxoJiqq
37YkQpdg5pjoJml+KBmS0KftJAnNLEB631pTAMTZONzcE3sEoOqBRpqa3B8kYK1s
lM4S2Z9XBL26Pz3JR/LXtiiOjRjhcC2oC8/Ybjz3YfxIBfpUb7nQAQ24iKnloOGp
+Yfv6ar9XlDI12u7vLbFc0nDNAU0xGz4/1IxLQ2hPZsdxQ6XUkP6mEfn3Phdx8Oo
6KREmyPw0QBM4iNu29MJSC6SwSoZ4E+qaCcNkYhwT8v9qqv3IxD2Q9ZbxZ3FXkYJ
aRMAtSrCmcTr1lRV1iP5Nrxu8mTqXZLk2pav5FxhQ1FB3cq2PkAL9FKTnJv3VIdY
9WpVq4mVll0fc2DdmFTfYi6ZePs9U4tRwf6yTClm0p7TMQho/ded3qrB2UUdBvZI
63bLC+6JFhkKPLta03BmHYfkZ5+64l8keb1d4WbdxxAWI/E+Ngv7V9Aw7C4zr0rG
x1hNnRW/tBfyS8bLkivyqKFxTwiMAniAJalRQxozB0ju81LQKxsiipQR8uwK6uwN
5qQYgxGHI+RKiVvEtTq7R8EeWETslXvWoWqVgmmL1+EYIN2eMuhvyEQJUtcLb8EC
FfLHc3UK/KfgsbJq5HhjwH+kp6IYncFiI2IzWUWKUgaiq5/4GvdeXTrSzHpLOT+7
Xbx5VYRs5utxDdCgZvm+VFcSojfQg9DMbIhdjRmhlR5Yuj59Ja/9HBOPi32X3GRD
B6NrtPLk1JsqIzEsQfTN7hN+Cozvx9OGzvztq64lUV2XXPaggTiEcBRPzuUfWK6f
8ZDQL5QcoVywnBJzX8mDluf9O5qI2Sp/S7ToOVvj7JPtC5BI+BnpK8G36ofhwGL0
`protect END_PROTECTED
