`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MIs5MCbDXcEIp7oFP3M8gMyyYvHYMOBBSmHiuXVlHSu4moF3LQkQF/hwZMbhGXC4
4IsBqMmQa+IjzIfTZA0y5q6RMrfHmImYxEoZsvRkAvrQiGuUJRcjhzrI0BGE17kY
kyxmjEY11qAaCrDh/YCtZk+w4H/1iswG1B5mul6HsonTX9dNY5sKbQ3qK35qsV8d
UT1in0/7upe27225jxZaoJdoxESqQ14v0exONR4w+cgwSM4AJr9+pTAJfm/CpWnl
/v/wEqtv/GEBU16+04LHg4v8Squ54CpCweEnnP2fq9/TpT3riLXOGJLKlsyEtuYL
iKc4vBdL/gbyTXhdUeUMPi5UmUpHw30jHiaCURN/axBc1DvckdXSsFe4CMTXK2U2
f/e/rE6oLYg//irnX2Pcxi/00xC6WvvxyWxLSEtWhvTVHmUF7MR/o9zNQD2svQ96
cAam7Nx6Q7+XpuIOz3tS31a6/Es98BkH7GlTDmlPk78aFd1iXuaTzNsL3EWHIcoq
`protect END_PROTECTED
