`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HMpnnkO8kjrqPMvwAqggu3rpQzYOFS7J6318PBorQdOkF3WGoV/LO1GRLpe3ZHPB
A6iDhfkJhx71qCWdrdc73zrffTrHHoVRWDfDjm6GsGV791Fn80vV1nkKAe+2F21/
8/Rc6uFsx09VvLIdkxDRZ4zmqD3PddVj9IQWYvvlunNFQf/+qJ/wy22+dfF7SRTo
aqfHkvtOhxc+t8yqqiILqp/dOSDta4iO5RQ5/atetUBjVOTCE3ybcoCJ7AEE8bhw
OaoDKsJgWIqFUEp3ezRBVr0IbiCvz8fMYLfvwi7Lmn8Cqdev12ic/xAXYEPPNT4T
m/u7Qe1uIuBjbfO3o7/V31OkDxra00srFQ5syHooOlglb4dbOo/boIkoXp5AvTZy
GDV9l73WrVc/SKIdJxwLEE7sr9AfMEto0hwx1B0UokvfGPqM2TlBZJUyrEysVXlP
2xzA1L7XZ0TL1+UXz77OBccizlQuMKEGqhd60SouvkoQqq/Oiy76Fgh/8nUJmGkd
PFhNsDO7Uwkt2Mv9fKwolVMdX2JgIm/CEjOKz+GyXwd7y6CES8di4bLCZ4+fmgQy
80RivqLjJJmntqyQ5F4J92FXx0bb3qs59vbulK9gbZ4Y08bXUW2epj0/0AzK1iyC
C8daB526thxeiJKfhZynQw==
`protect END_PROTECTED
