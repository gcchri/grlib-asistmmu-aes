`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oPyOHBpaeo6XNwofM62Ty0pCL9qzUND4WUh2VRKBvgrcXjXE+Y7SGW+2WDH4Vvaf
ZAySoXrAWYNnBsdSDCeN2scj7uWoO0vUJ7VZGEJJawgSdfL9x3V4q9NbMkeYtrK4
l19Rehr9iwPgWNVKmZ7P58V1Tw+udF0TYVrEK2ULBxmQnaHAOauAU7YWAjFciaIR
VBUy1rC/2YfRE4y46wc1A70tKzMDtBlua/lHOiDOM+mp9XXDPixbUWB6jWBKGuRy
16ukdvfxigtdRtem7WNMw6O1o/e6YzXAKY3xoKpTUd7azNZM1Pm8f8FImrNaBXLe
ov9ZklMGwRPzU0zMta6BzJlrz9U0E/eN4nXqTlVpybDhgukIJ5vGDMFkRJXK7wXc
WShVui8/buCONmNT8TnoF+Cx7WfJoLiFCYLlwkCpK6VAvypvXUGpEOr678ohITe5
`protect END_PROTECTED
