`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sv5evJO8Q4UVSVkB3ep38ziw2qGRyVnc4M5wE/ORvgoO+CvjdxqHMJ64cBe9hnFE
OPPKwprQk6HfJDAlp2qL4CSRGjiqCwN8A/jVx584Es6kuPcRnFj5foL3bUbqJxSa
U7JBtQ+2llzMu3rUQ2gggyfNX6HZdvrfiFDNd/3OoX2w1eKtF4flrtMGVjlnTPqw
RBaBbbWypteRocHyHc3CmBvIKf48XwmWU5UEDP9i/ALhyp9GH40ajCE9Xy0YN8Ax
MTDafTxtMh3Y4TfmNy7L7X4y9g7sfGXO9xBkq1mKQvggP+umjCa0Fl03BWL9/9dq
I2WSFEmEYut32UHiqwDynCkyqwKgLw7t7F+2hfKjyt5Idy3YIypoORi/UzHa+6X9
MDF9/tCq3ZUw1cFU01zVgt6HY5EC+83/DBGjT7IbXVXAZ73H6W4NEQaj6dtBhiPK
iGeibMtdCeW5suEP4zxCgHTFlQybf+UuqnE0DMF9XLg00wPAnkO1qkMIcbDfitlA
UgcUeZBUerXWbi2wzVNXlpw9nP0rqMiWZ81W+mXKG0FB/G9ZV0U7It+h88hDdnWQ
EmI9KyuadG4JwrqpByMTGwTdCkhCSfcLVEJTJ755oLgSc0l1kVigbuX6yjeg5num
OPpoOSq4fseOeGrgn/30caaZR8h3nlIjuhZmfXi3e6Ul3aZ4qguzBtEE9JgYpjtQ
csA9dJp2moRosp/YWTsTmOICRV79lffr7NQg+aYbsC/8pJ8YV1tceX1cek0n5H9U
W1B/KCGH4s97909rlAWq8rB8vjwezhBUPhpf2f4odjSpW7tCE/yfk4itQxNumvv6
uhH0t5rqPMWXAzhU/83gzAN2cC/KxdVyNwRMBxjg28VKkTo8/u1752xxdB1s/D2X
murNuCqvhf1uh/iWAJHBop90DEmi5c+QYsiGInbxgd3ufWmLXUFtA3LXHZ7i3hTa
`protect END_PROTECTED
