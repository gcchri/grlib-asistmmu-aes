`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
64YeVet+tzY1bgkZ+KOq7/wBN167ZuIT4Nuu1jsepCkIt3En45VKh7ndyM4+sodu
fmYS1iGZUXMgSkXOQAQFu9HuEmE4GesJL8TbFR+sQlHzxT9KGtrWZOCf1Wg67vmZ
o9gijv8aw7R1TtYnmazAfbK7dRw99z9sMOk2hXs51buL9fPQX+WIZfSnKYsYUezc
Lr9LVpbPcFUNJa1YHfXH+zInWLGM2oU4s+kOoF9JZckx3Ggbvi8GOGRIrL/8RLMJ
33Tpbe+PPPbBt7A420ThnW/8yBn/I+rS7/+hAh8Y7fVVXt4xJA08q84LvyCfnrWQ
FHyDf8nDUiSId9WTWFkEKmcPX9QpzZgdPvwAc/Xr1+MP3/18c/HgYQ7RUIZr+2h0
h3DW5aU2FAZEp8OY5GBnFg==
`protect END_PROTECTED
