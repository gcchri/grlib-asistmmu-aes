`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YmSUbLodrFgWUYORpSAP+tdrQ0/zZC5Bzx7v/iWchPbpUoki8ZkB3DQO5FwXyLXw
gE0/05OZ9r4xCkg3n358iPO4OXY3SDAea2v6bZyoBJRaoQeOLzi4Xr5jn6YLiQG3
mAeX++ZZg2JRdcPKPiND3IiURwBUvkTzhf/4Fb8fB4sQH7jdGeEu4UnYm14SSV5E
d9vqAWnpXi5GyURIhcvcEMXdeVsqbVmFNXRLTWDBs0NqKRy0FpLHiJssmmN1rIcT
w4hd1amTWjt+aVG4n+2cRDAanYImNGQpaQgZaAcTdh35pSHgf/dMe5JOs7iJBXLq
V+NakM+j6LLP+q1Hr1GAl/DRn6muvfJI8oqdj5aLtvOShseP0uPo5dKEIIwNkqeC
TaLaUMSfNn4BQ7XNyyrDJI8KFci+XH7EoSbYAj6mt8C/inDWgGx+uhOGpB++Ijbb
9kjiK4/tufmB0UFewOWzyzHHfBtBR8ElrWHHPvdUw9cgIY1Ror7tiFaoZdF5OWvE
zrcBt/jaBO/+6pEMwV6oSl6bFKJOzJ+ehjMPoTLV7WrJ1ZHBrta4utTWQ01PHXjM
DxGmRyR5CzYAklXxzPsK9oDXGC9uD4NE6+ARBQBdn0T3PFAlHqLy6uySw5cdZYTW
PSnJVU/6XqSEUQjzUkg5dnn6XiZoGPNgPMnxWt7FVFQZ8UHq59LPWbr5L8V7G6RD
IyzQz85lQAdLGCVv7ibxRQt7CEFu/VhCyVm2+jNbCcMKreksB1CME9KLUgD+UzxJ
8OCf9c87O0uVRO/ATD/tO/SPBd0zv/JAd+6Ey/Svj1KdeT7ciWzJ8xQZLxeYlJpm
HCHo6GmWK6BQn/FLBc3kfHK/fxqEhFV2V9Jui2sEQ9jcMMEjhC6P55Lz2k0KTXlP
BX4SkSJ9Sc8QWbbwFztU5ZAUSD3zG+1AnvZxNpvZMmiFRowbWMQsCCLJhSYHwCPG
TflC17zFE9Hil4NrEyPeWrGXSUz5t//NJ8rH+b9JL4UBm9HZnL1Wfdmz71KrhSbH
OFFvrP5ztPwUdETABBsx9RngUZmf2xjEw+BYTNaaRhykeRaJtps8/wLU77eZBn9f
`protect END_PROTECTED
