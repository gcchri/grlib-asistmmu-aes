`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2BRDfB+FNxxUe1xDZmhT31h9MXiT9GGBuavBAAWsKQKVxX15tgNh8ioxHSSeP8Tj
ibbdx7DnvKWcK1ootZeNeESvryTSoKBSz4lnpW06grR5Fac/BwStW55E5JbzpOQq
S/VNg2DcBEvchF9s2hUt3b0U4BC8xbwN7fU4V2Cpwdr8TWosml3pv5xcb9GiMV3M
XsGomiJbQP6lkMpWDlg/VqMdMPgBinqXDpYUfLVzqnBHoP271oD+J1NrC6m7jfgt
m5So8/Bbah03hzV7Huv8DDFhDKYw3Q43J7Z+BUL6T5KLG6C0IaddNW+5H4s4QRQF
BGcTPadYzloLgxLuta9QAokMctGpn/n5+NNz09LIoygFPvHSRuSth634Up4K36rD
DQWuEWOthznVNqfzQ0oYVZN2ULrbT6Htx/23J0x84vrfGHq/sFwFv5ECz9OwNMES
j94Y2pnA+TYLh8npq31PppghUNC1K8UGi72QB4X/hD8=
`protect END_PROTECTED
