`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ofHnH3CYg8DUlIOFhwlrC3wCWpVq/7v45w63s7zl0APaLakpD1RGKiWaQ1heUYXf
uWNIcyOjPAlu648z1RLJdIfjmFLMDLQZbGOf4h3wyAZjEug6mVMrLZUbwFUYCESG
6e2YT0j1VIVYVO/zKj9uALnTEtE+Og4oYPKwPd2dxSHPmB3QCJD/u6ZW1IWnWkTL
hOvOsdFUwfBj+7jyEOe3Yva7Fe+Cr7VWhavfTcwanx0bgsBRCaM78kWRxqGfc6hC
Cr7fsXJ6E6ic1Dj9DHupcmkTXcA7Ka9R7/3AV4LghF/QSofrFBcFBChS5cJHJsiv
LeIGvTjYF4Z5cBSO/LTr0wDREKo/70KDE5bFdYWlOfEhkarUTsSncIzXqvI2WUwP
vfHAq6CvGgyUyRs1lBd/c3DIm6CMirFieC3glUQKIB4ckup1R8/CY6IcbmNst5rd
eQCxrXTEg9vZaldfQBAoSB6gbMW+6g6HX1rBYnXrwPo=
`protect END_PROTECTED
