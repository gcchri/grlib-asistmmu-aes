`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hjv5sIEDP99/+kpZuT7oaADRMqSBim2Cq9WvzGx+m+jo9uwjC7O/8OfZ0eVGu+iM
cm+byhqyqZI4VMq3sJ3cldzxT32i3cOnJJZPtAZSOrCSmrEzBfO1iYSkwTP9mZqV
spgThKU2NxjlyaDxe6SU0H/7gvsCm/lH22PLirY/6R8UN4XbsrZjIMiWpPptsctD
g9UPm/MKYG2yBoh+qqSXfrKXRm7WWAqN2nF3w71xwwOgxknHRTTmiL2I4TIh2laZ
NbmHtufdzRgDspn0ZaGKHdN9j6LURAOebo0dvcmYqpF3VgUPk8TgOkuYQq0TihFn
NH180VSLvbpK1peSqK3MTHd6h1jgofhNf5cKtNPJclZr5fxbse46PVBQmXINbdLC
N3Cz1ZpGM1iikfNnqUXFX78E6aDNywEv+3Ghov9bYaGgwH5WoYAGWMhxaxQdERe5
6YwMyXF3+RPOc6qZgTcd+L2A/brw/XA9m1qBb9GatK8FKTYQojTlmSTxpzSwiYId
ge5e6pSa17bL/vnE4dqzdWVSbca06WCUB+cBPv+Y61GGIFAvsmxA3jjh0xJ6b2k4
0rC225U73oZ3zXTKUISOSu1I73O7EsRMn/EX/DeHtLBcw6LG6bs11xokLflZR3Du
apQoTCyYSsFVtLk10v0rCcILHXeBw+Zk4yvdKtZ3Z3VOWr6VkZIa7QyS9tYwoLTg
OXZLgLcK8M6kwBMFgv+fG2DRIcU6wNGXoTfQKgczBA+zKaS/c2gE6TXTJTpdZ08z
m79GRIqtGmeUF3DYnBbxp4PhceYFYpB584Ts0J5qZPT9LWevlXLjXs0oG+hUBVlp
7cwb8WksmAeMCJO/camH0bVm/H3ds5BSXUiFR6NuAqs+7bIl7WTajA3X1Vo8FcHt
fJMUb/rWXImqpmspGrTeELxrg4HTMoJtSi4PNBGLyCH+MgoyAliOLFlCJOLfvLJG
NzOhHCqlKkHlkPgl1t3hiPqaX96UwXhIHVXFOhMTbUB4Y23iWocNWT9qHObVIToY
vQVy6QFHOEoP8dgK10oeOzAhj4kCD5zZXGKWmhb3vU6Qc8HLf7r2QSxNg6UH6QFK
AEse8DBcbuL/jeKfwJ9RalQBp6deWbSBmOEwe0gcm2rJuLAcHQRIHL3KdVDRwiPv
oqHBtWNtS5OR3JxitUq7Q+iaKfB136+5GnU8tK9qrB029+ps0QLNti3jcved37qd
T4Z7BFGFGCuPyDoGu/p5z1dASnskzaHlihCKo6WmGvpoe5YKQxHkthTwcZEzGDSO
P3jYfgTHkSxoUizvK14MZA6XH45ux7t6HHOngg8d8CKULlxrRgCS3cFhsRszU7Wj
XXUeZDqwyo5/BxHfAMeBTQNRJDSkrPpPttqtSzF/Bda4aw9CtXjn6EIYeD1dwtbW
GbXZnKcLGxPM8l+u2nTrLzToPwb/BpMyZ1nUGAU+mLZZYbkPlxCLtHOuawHn3fAv
gaYoTSLpsKZ0chnC075KKhsS5ldJZLOK2xbrNafeAEMSHQ4lfe3szBrMsOu/W4+Z
gggq6R5YJ3ZQ82B+0luD6KSwhmq2lqhYLMI6RHyY/vNlCxM218L1RK4/03LEVlTs
tVBIsXvVRGCGOft6fXkkIl8NwDM4azZdhJKJKhfeaBJAHIYxjPxKrqWkg/IQMIPh
H/7xZeOWmUO3uNx1cfw9dVixjJ2d3C07VP04Pv3LKf5DMdI+RTKT1Bj5yWrzhN/J
06wcY98nOeHC9nDz8yJO3q/Km+OwWo5/1zbS+Uf70G64Hmg+fXvmL1F1zqXgOuXZ
YimwBR9bI4eawnOMffRo83lSf7p9A496+NjrqK8Tyi4Lc0ePmgmbq1Io4HZgi/Pm
wllCIGWtDjzUxjFwxOzrE23yE2EmXg+RArC8BKlUwl40G2UnKvyb6v2WPQlsbWr3
5tANZdMBEke2Zu0PDFKmLPv2ymzPQSHz0g179MRcyHDSZWM2FbdiQ3K7Ir1VSZUm
l1UuaZt0PME/PyHKA7qUPd75tju4BW82gNuch/9GvWmb+xyX/WVZb6wZ61o7+8DU
j1yBvNE9PBpv+ZYiCKZDolU55r+NH67libyejIeUvBeI10YIQR9S0DUC61VWwOj6
EhMgqpQWMk+GJn1ihoCGSgn/KMt50wQkoMTZl0Ap9ypNz4fg+mJNTq/1KsafeLx1
ssC2kV7Q/IjnaNNZ/D9tAsgzGXdfAZZ45ybzLTZOVNnh+Lslm/aoydJu+0nW04Ov
gxpfd1OzhOolvGCfftf3RdnD/SrveCq0sCr9arJoti/caKZ8ydkZ0Fpqv26nYvL8
j6X9naiGGrlwwTfPKW5pIJmSSkyPJgAg+Vs8pJEJPkz+DEVJkuZ7CaAuB9erVqxc
8KylgGm6UyuTiuiH3hRxQgmKeunevi5ENGK0FCWHKVxbMDYnBlhxSXwKMbcyMoNq
WS7GvXDQwd2dCXSW/8ZTr4Hq52WvbatE9AdflDeV9T3Y7VzCR2VHnqTVe162JQ6r
Cxog0cVKwjQHcOPzj1YQM6lGAITXFxAfZqRxfDzovPF/ZSextJiXNNg6ayn3JyxQ
0/neSzTBoAueJz6nxMJOvck6A6UKGUoKci8nnf+HoYH8RAWznAREjy+L87svHtf+
WHZtH4l/gDv0wkpG3g7ehbrQXvvRs0awudjNEHjqegIf4rMdFCmxwchI+eNL3ioR
OQMA7xYaLYnmEz4Mm3Xw/khAbC7aTC10XEQlaR/zrTUtinzLV7uYNI2/rvDOpDKz
a8yqnrWiDBhtDTR5SEaSaDUhk1HQw9sRSp5UF3xLiQDQDE/GxyacYYYy02/oI8Bw
SAZQlGqGIETIm+OB/PaUbsiqAMqvSZ1mommlX4xiVcs=
`protect END_PROTECTED
