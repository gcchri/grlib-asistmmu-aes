`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5//zXZt2yzJ1cRpdY8nE0A8fsM9S6PiIQHg/cyzaoaDkurAdcv6mSK6VT4t2NEVU
Gk4DxUKFBrdLMPbLMo+1NykQmd9NXXkDu97nbE3WNZOe+TtRD+sQi+qgs1xVCpPB
6AfujgwggGXhMAvWDPOHwIwapC5OF3sULOyH4GJtCq2m4RpSSwiiWOtFM6bIliAe
ClgPpQLfl4fJHGKSFuf49VZEFFhgXrrdpliJAig7xtS8zyS2vIOqshp2zKVprayD
61jE1xPuTFT2EuPh09LIUnSaMibRLcE9mBHshXCqCQ0X/D0pG9sgFRC93fQZdAXJ
CbfZygLAUDjLLeqCqMGHRNaS0LOjqxoozXUpPVmgYncHqSoSuzOd30gxVE/aAJhH
KWN4IKYYbCJjZt4SgCGeAirvUQveD9YE1tfCt70+2N3C3ziV9VKJl31aLYtxTX2h
QJtNO4nOQq2QPMW4fYXfFQ==
`protect END_PROTECTED
