`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WZOLAlqmfnXh4bdjVBguoengvFpbmmurpdfRvY/XYQtRVM6JnKnzJvFzrVviWaRO
e544tWBO4bjUzQqfu9dW4hnb50gFe5gMwOLJYW/qXc+gggx7kl4fiSOryKXkH3LD
aWUYieu98XvHfrS9GsIglKyTT3wkLiOKYvUH7lIx4krth6D/LNAGZCqV8V2FPx6e
J+snbMme4sPW7+I1lVDxdLLP//B/DqR/YJXMT9KM0nGaRuAIqbax1enAyB82blXb
OO8gOmzg5Rya3cf44OTzA+ylaK6uYgU57sddyP3cGhrIAgwKPVnmARUg5uKrBIsu
/K4tQFWngsw9b5QxqLXGcq4lx7Z8iUpDEiRip7VrUVjRCpziNRE3vPVhpRqFvp3H
`protect END_PROTECTED
