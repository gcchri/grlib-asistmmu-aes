`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bsbrKeztmmFSr9Ay9tO6vwboWL4fIDc4zDCZh5eErVfxFBSpR2NCU42fbXwg8r/7
EVEH1KVXj84/LlDNXqu834aw6vVXDVIEsERMtct3weH+fBAZZ+s4rYbAY8XzJff+
TZtCMBMsiItHb/NCLyeU4tHgBJqgj8OEEWUyxc+aqpga4HDSojfqK3XM7bcBsG/6
Nl+9BHPR122JbALL+Gr9d2rto6FWI9MKw2ZRI8NnKw5Os1mxxC1lLoznJSnrZ65X
vruUHEmQI908d+9l5y7SYh1rlzHf2bTARzBc8jKsXBJMVR/bPhJK7EMyA5IYt9l9
J/VDQPUXCwRjU4oPlTppafjJR69hL2w4XFIGJ3YtZNBX8XwC95cMJMKM70N1EDC0
AqFuZPxbsyD35lz9U2oaPniYt4yg10dHQnRYCX3FeIL5Uds5fA+HGNu030z+knN0
kwtDpQCWixP5xF1+l448OTeRlgL6ezEOjKSWxJa34pE1Dor+nfZG5FXo7ERnbeCd
L4LdMSKzWB7/MQF4RSOLPgGon1kRurDQhSogD7XunA2sqHK1Sp52OAfcXdzWRYOx
9LsZTOnfVWAK/L0fsw8ONKcoPZGg2/ZOYvAiIux9feMTrJofnmcy15W9yQzPpBxc
jJQsIK65DGWVD6BzqsY8L+Cw1qdzXZZmAlqqZvEDCuLpYQ4YaLorG32nRPVYR7OB
8LMnNrL8CPFU1eLEwtub6g==
`protect END_PROTECTED
