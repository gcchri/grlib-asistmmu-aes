`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OxXP/z9LcaO8s6aBmrSPMj/mCwjYFFrhhUdgl62n6tjwbKflcLR5hDN4937xFTlm
htXcm3hLlI/nRfDEMpkhmqYgTqqPy0vyt5TKI8c4HmB0dvqIobioYgd+n/bNwl+Q
Nh/oxSHE+eJd6E/Jy2FJLNPgX8nDUf5joEKIlz0PF1L5n0XxqyPt0c9VwzvqMJW7
03Uy/fCKFAXy4jcmtdJpNUhdeIiVy4WHCJAgRGFwVc3kuyM1BrGp4XR0/1gCuurq
GmC0NJ9R7to8wA3BPRiJlBqMJPU2/NJKimH8gteBEwDPtc2ZR1mGXyjsY9gXkk5g
AIZMZWSLkt4C18y5eGw34CcgdyLE6WNb6Ep0QQkoE5vL4VkBj77b1NZqHKMEJ+ol
foX1f9QMYXg1XVufkmEdfomHfo3G4/79eOGwhYz3eMfd4YIjKSOSVvLGJ28QETdp
R8tpQmYqVP/nZy2y8LqttmFtAO/JrNBGiT4rQj8Qxc/xrzyLLsE8UvwE+eJCrPLs
3swAEFUD3hwoWA/89GpAXRWxQ+1u352GzONHxlGPUMe8qY+c0HsPwFmQy9WaOcyh
RW/dDJpW1Cikqh4OrpEJnil4O4+5NTHiD96MU8vp0KAGUNvKJwQoUdplw9OC32ng
qpWrLV1DdDbCyW41YTvgq1VGh+s7/NxA9ynVgUfwUQ0=
`protect END_PROTECTED
