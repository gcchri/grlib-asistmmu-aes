`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
66ZG2x6Q5T3GiUaWwOifRywuD0zVTZRQCXuwSJ8CysHGNyhunrw06lnWLiuspkit
miCgaawIjoseX7h2bGy6PRFEYxXuDc+EHgp8elqbnPYRJCzEu5WKsdxGEo0hIwow
Ru6sZimEMIxEaIsQEJOs9CU6XVPd8FIAK1nA7Occh06fiar2f8Y1VD7eFEI6UmFW
vhBsLZZ6K9VfHswt1IugI+zAZ5l7Owh15FqEzJl6dZMb/m4cULyO73Ew2uIr+FgR
mXchznL9Gv1c5aMXseLZc+DzqtP1WqWoNjnp+GgcHCxT/cG4pGDffUUuPa/sNvhW
slvkux/WLxZRsSsuOi9Ij8EbspTq46SiuIYe13ILOo/lsLYO+gN2IMDMuIbE8Cc9
Sx52r6qA23ldjq0hb145Ladg+N0KYh7IhpOLQ67XacHcY05cPLD+NL5qUgEMAdv3
zrQkCHv6Vuf82bc1j3eAwWX1Fzs2hrLjs6o89WHF5EHpUkTnVHdJ0OsKzczsgiyx
PtdCPoCFQidKZyMuYx21cVOrFT19RPPFbrMuZNvxW+Sm4YEHBsQ4hW8SgQOBigOP
eiOq+65dlIfUfUGSRZtHqJYHhd3Ocb2Pj2oUdiS1Zqscy/bVWGKx4oTR3Bxz7biD
PWMQOdiGtr3zT0TV8phGODQmfxj53DVPyn23U6180HrfP+avc6JoA5WuekgrBypN
ruO7OZHAr8BzwlwVbwUhRkSGc96xafXOcEGsV+fD+oeYB7KrVDTqimZAOsHh7RE5
NHmvT0h1neh3Kvi/wkaD3KzkKGRUAlvD5sB/i61Zf/m/cXlWOuV5DZmR8eTdqFUl
8dnmGyaj2gN1h9Of4oB6phSjVOB50k+4kTM43xl5n1s4dpFolw99FCUXCKJj6PCi
4yRB2mvqL0M0Nhs68XhLNptTdH44dY2C8p62focmPKVzqtGrKBhGeeM3fPkmy3Fa
BwY4AVgCqhIZbfd76a52K/9VNpTfeyRTp7/wfcm9c1LRakR0O2+k0/XJgIbwO475
CZ8tO8EEIr3QuNwfOAybbS960g2dohJOgjLmvb2XqlAkLl7dQ3XRBNmzG+xMxp5Q
2zCvHnYdCxIJxK7ha48vrlP0heNn4lUTNba5bKJ+J6h3+ZXIJA50jPpPypK1/eJX
hdkOJjYl41EfZwHHjJs8zGvClwZ3TmToHRNkOYs+mg/JnBz7QSkcBgoIKtGK+q37
lcSHeu2jz0CCQEL1UlD4SOWtNDgTcvYlXR5MidfGYvnDLdqptI5RFxfVt31mp09t
sepMLTmdhSakqf17IftZIanFCEPyaM4y9FzAvf35QQ4oL1vS4o+h4vg/xIgqzitW
aTaMNjTd6tGF37MaoB9YlfgkMN2wlLzhwNGWLwna/nDV/iqAkuqgdaFrGpadmh5z
mvDw92pR8slQODlSSFSh0wqopuyiWER4BaZvdufWGVFhG8f5VHoyoTXIdcLj6AUp
1lq4W2gXeRZW14QZWQojwEtbp8w/77NZpsgDO3AbPTNO67+UdoV3bZXXV44ev4HO
OftuHABaA37m95CiVN76EUi+9CuJkvffN7XOwmCpfMO8gMngClIgCjikYWjPo2Fu
uCfSbn11evQXsNA8Qe6dhX/g8xUUay8UYuOuGDRjxA0ILBOXLLTnLfD4xEJ37P+M
bIVs5CGI3Br2+y3RrU7XSXH7nOSP1bYMftOUGG1xNFBXJ/rvfeuB/DhZj6gIoAeE
7iJxHaTLANZzcNX/lrKCwd8dYSBCqIVOb64qtoCVW8+cBGhgem+zl6wgeo5Cmb1Y
QIrQqwyA1t7ACcafjvZaXvSXGkEnQsj0Xvkvq4yqRSEiiw2WXMcUN5ZOtLf8doHD
qRFKO4xMRwF64FokSBAkcyb0JFNwrmletnk9t0LrbKGlef1k/cKL3mnpIjRXrQWC
wsKkk2u/YGv96qhOMqCkP+KpRWCtvJlLdtTmH6toSuMuGFLfe/9iat0JiwNRfOzE
SLAZZWLiTWYipxvJnjzEk2rBDc36Qwy7TJe0ndmrRQnnb/hRjTQMxgy5rN8bhGIv
GJcsCiguKeKCSbwLcNfMetVp7VmG1fHJT/ZGOgNV1Vj3cNiAuJy+RQsVtikkQY06
9LUYqLzwyj/4xQ3jZPiUQMfP2+nwxtXL4Lj8FSI6xeEXDOcG+Ex/DVrfWd+CKaVq
MYrZwlPTMjWOpSY2AkYuEpgDedTBMvUuepOlgMluj9gOcVAAvf597B0H2ZhlAZMG
+Bbusg4gNFlJVAHx1FI3KrArF3E4hpykcLQYvTu5DNBTTlMtazozPkSPvlSW94Af
N689SS9Pwb/Buy+iXkQWbb8TvtW62lEfrFTGSZlq74/Gj6Nfio7NVqfn596naJj6
AB8e5qhyn4akvoIudleBIfAxxzuG0gtObsPOqjgWyOQiQD1gmR3KmCnQ1EcxLw0r
UL7rOPQp19DKQ4IOTiSeVA5t+cmFw3WYhlpEhqZf5URHT5rT8grHvlxQJHQposbN
P6fW4RGBn9gz7h2Q97BdZAqMhhQ3r3j04ELq/49WRyFtqCXuppxhoLxkx//ls9kZ
ijp49UYEqZPbaiK0z37xUl83S7gaJBorWeQ8KyxZSRoKJ+SQdlIQ3bR+6AOj0CQH
MUYce9DfqSBDPYzqTZ0leKPPeQKgsq3jzp5+WmfKhf6R87PeUhfOwOJuXvafSXvf
bPgaFSwgczv3pNjfIfOrDmOlqSWSYh86UTWEJ1cFyKCN4T4HXD81+TNdtMtEQ5u6
rqTOacdjSKSB8oI6CwEVKbf3+t8ctWd6Qqu4PpstUGJBo24TrfRszN6/UJRvwjhx
3MIGgcVF9kgztz1/GlxG7KX1HWW2O8v6/eLZdV4QYfiJ5SoB80Yu541ST7qYBp4J
cc02YYAg4ol1N3W8PLeB1K4fXkCUjlWQuRcN1Xf9fJ73W7Mus5Ivdwyh7UXqoLye
F8dk3gJL/tare1mGtp0CoUQg87kQEtgsgBhBfKaqaPClFsb+p+qBxR4yf8NSyHGy
FUoX90+GLh7o+BsSs5NK3aU50vdy3Wnb8UdXFC0gDypPdfHzXd4nMc/1DVRVIfeb
E2KFSSTVQu2wqsDcdD87H5KkIo1T820ek9wwbsFsq2UiMsCOJxIgKMF5VP7sJvxz
grohTZGwG/dkmYYLjZdWg0IW4YBQakxfPkGQwi+SlDshQq36zcqnNdKsxAOWatFy
U3qyc8hbD2RZZTzk4AroCLtztzKUHnwQkESt3JHwXnuWks448k4gLvc/eBxbw2Ve
0SzmdSTvePYPN3JkCife1Xv+w7QE7VaTdQYIVwibLbymQLmDvIMAszcMkZCLKlUd
DxKK6PcALbRq3L+O0SDlg+IIiTLUiH1cUBbhv7cP4PXM5Q0ZPZqrWXkmrLqpSolQ
rtSCilGWfmYKUtW7MC+d3QAB2HXKgl36c8PwtvQQzbdfInQLgCcTcqIeT56lqnVq
On6Fvg1LMtlyNG6UmYcRub65bY9zclF0SwmXwKh6IDzH3dz7RtWsNxVR1nBF7LQf
45UFoQgMoHP1gjtjF2TqvoT4QNE5mwPFXgMQZ9N754y+A1cFvXgnyehtH+5io2GN
9g7OpijZtrnHoWRlmhLM9C4KSEEphL3K/0ApBcrnBi4KSsJELP5HDgPkGMq97+qV
g/zYxbf6EpWuvJ3ZYULFtobVUwqOyf8PekKPsTAFPaZ6SrNSiiMZMEoI15fXjvbq
4xy3Cx9n4jQUIKFczsUCGHZm7OV2N0oIpExSyH0lJE+pwS99bULzDfvwjE/cc1hV
1FnbPZh1CLFX6Uyw/+iRN9NJV8WNK82aGVV6GEIIOMCnfEMIjJKt6pqAtsu/1a1j
MpQWw6QzcSHZd8+k/B5tno+wIlY9RIYBzPCzRym011EDtYNJUvT5RzR74RpW3rub
IEpt26HJQDvvTydv/vHkRDF9yLukix8KEqp6RpSeKhhNuo8Q3UMaKJpoY5nJlckE
EuJ/UnL3ywSSm/japozuVKE7J+L7+f8foPyKPZY9elpFzUmGbt4tCQzmXDSH9jwc
TAgyQzy6Em43/5JkqMHvtV26/UUEfGgC4B9Bo5iZrWyQFaysrTgzwPOzX0brNlS1
CxMlGD6ll4AV0gx9IQB7JJEGBULvyc4jr3TiE4iade1IiBAA71Rwsd3jkN1veo/e
fMzNcVZLLeWzVI/gQfG2AAsJadXzUgPzDjcH7FK6anhHNAw0CS/fY3/d7rcMoBWf
CB+YAil/5oWCy59KWu+Y+S/xr4igqHdJxCeV3DWh1ipF7MIe9aERVjpHUfmtx8ok
lx+GwidFfWM1lNm6kObMee7HmR+s62jq3lMVmUK5p+U3ppvyhc75gi9ho50yCzzp
MEdFaOWg9k3TXBu/j/Z5vPOed37ua+RYqQV0kSaxpJEroJftiz/NXyJM8pioUh79
V9LZXF7MHXj0slWBAj9HSg+oDS6axvUj3NffYS6uiAEtRq+844UR8iIfupTEbDTz
HstxjmqdCjD2ZOh85MjWsAJYaUSMXRYiOjGL9ozBAGEta+g/qCOJGRc5vTcD0C1V
DidWz35XEXwPKI5fGaXA7Z1cKbmynBsSS5a+3n/xBe/mYSP7B78jhBW9vmQWrfVe
uJWwbeoqh0twVmO5/TVQH3UXuwL3m1o12lwXYHGHN4hXfd+ZR/wK4uSbv5rsl+Gd
rBRrTFK2K8+XIQ1/5hHIZwPrqQCcmfBTQWd7o5cuMI9rF0U24u15lun4CnSXWCtU
QvFAnAiozN2Dw/loGNCCVRBf9pI0YhJuBGWVKVBdinVcEusUMhqxzQ6V+OMJ8ZaJ
FzdbCXoGWYxPOecyKcJLOJDLMo4WRz4t57pVBIHuEDpBcoRPHPuaFCOhoMwvxcqd
dkDzA3Y1Ipc2c7/DxM1bPAxXKJ33CtY7RGZ1wRSoc2Kxvc6Jrvu52GGxN/nHTMtS
WuosmlxPd8TwE0BqOSw/Q8DxZAzNuXIVqTpY+R76K96DN0TROWQuNCZpZ2tWkZRQ
tlNPv7V6BJILBsh9SBrGNLuzgcCLfCiBTP/L+MT78xkB4xv2Uf9QNZsmPObXp1tr
5pjRg+r+8msL6RalXRwb9zsfdfhlzh6YMTLexuoxFejMYfT0ZopEyGj+SkgsRfXi
fT0rcV37ooC5c/ZfFwaPvbaYAwM49M+cSXcFPYSQtD9Bplhr9aF8U1J/1GJdPJtO
Ys1yTKuP36BKkRum98Gf/3DrxJroAZf+uPlGrQIexKahy7X0pLTmv5GUfJVsWhxW
BXjOtDywWQjtb5cSVIR99+wfdFatZU7hP9sXQWsaHfYRR7kx9JVOwTM7h3bMVz4a
96U0Qg82gGytTMSTmCXVXQVtlPtkyYGH0Oxq3j+7Is9AFw1SS7YV9A+x2wWtlN7i
GSgQt1poTPsS6AzuuFxL2P4yxe176LSsDLfeu7aGuqNcne8BEs9ep8yCedgfbFzX
8dsn3lnipZPiiYnGVxcCRIEgxHp1GoLX9KvUJIJD9EBFnk/V5OXiidBtJPQ055FC
tz3PScuiV+vPkyjr/hA6Vbr++kj9pbSVgGXOn/HdWHLhDOv1HHzvGCRTkjCyCl0N
zzaBHKBKvaZ56Z66d6K+ZVtEhggf3Wy3sun/aK6FzigBxNOMrbMYmBpOaSLya3uk
daJUCkRSsevcFf/tFc2md6V5VLQ9KcwyuugYhRTm9vsM1HGVGcRjWAwzkEJBa2CN
0ka4+EgG7vBoFoBvhHwOY+3iD4MNqZajOsV3Sli+/sl1RkijFX7HFbnDkwViUwwu
JT2KmqtXR1YyQ+tsyL86jPJlcIEisYSB64K6tv3qK2w3vfyphbeOEc1Ba8uL0bex
rat2hV2EWg9PDPy3+CfQ/WWs70fRFoB68j0iBiSTmvCKLgfqX2TgVKO1NK5+MpUb
1ybUkvk6+X+ld7mgxQKWwusT+q0V4AdkdwCkb0pzUC8edhOE5d8kRfLGhky9gMqF
BXRIJmP5FMQbN4wjipxOHGQ+n9mLTDgxqqKytTW5Mzxp2XzpisKrHpq3uuaHOXVH
3QX0BRfWQYNB/ab2SNyqWWhN8d0DyiHF2oQoKm9BtjF9a1xgfWBcz9GUqyck6pod
cf74yks7OqK2PvCDKO1NiunBPliD1pip0DcTyhcw3axqKTjLChAqxY0FqHipIXdb
Kua6WdoYTQkPXs/m84II3ZsbMu+xfo1+SzYa8uQkaw1YrN0BeBgp50mE1sKMu9OE
KlOw2sWVNZc3Az42zJyRVfev8HDu2IQQmaSG/KQK1r114NlSZXhjn8lpTR8ktYPs
xZV8TQ+XRwJM+qOv2IL/OB1cy06dKEYB0ZKin0iLKoH1bN61zjnEUDYn4ZXNC7zb
iD9oIsU//L5g45KMkggGAFfT220VcWeimgUByMVilnMclwRToHAIvHDghiPsiuNo
PJP07YuafZKuJhqfeO354Pr5gJXxJpIU/Ew6yEl4hMN5PCXbJsmmF2bPOHIUBxzY
0xcDFijwDpFn3U1VnvdMQPJNqUfI1ysMSFKfdGLbegCMp8AfwpVf/H42od80q78/
wbDpzFNCbaxBzyBlXIMomQPKvZxIDbqt1gu9F9z6VUOxt2IOQdECVfLjzN+PUJj1
D5+TkMBrYO7/cEB8PoDx5FCo7mm/a1EbwANkzPCuDeXtAA8XYz2JTM24cHhmXYAL
EtOITjwqQG1EAnxeJuKFMqYqZNtFEOKttV6N3EDXNClOVSO2fLhRwqOQm48/um57
/+9GpZg7fkOF34mUNT5A7GC2tfT2NqkAm2BoZP5uJXe5iqm0K8Q3FgrLmguHLXmV
V8oAfdwIyjTkf5PxM9A3ad0We5v5Iz+XKOdvji6n9lua4C2P1LeVgCkv9JjhHYCF
PDe8u1KqVT3GbC8hSDX2ks8+HgibAhi95cbPDRHRrN6157J4NixTu5mhqHW/A+wv
8Xd/LkK/s+tW0Kpq1d8eeZwW3IaaZCu9ZYNxIVkwHm84yQeoSB59VYUhvSsFDz8u
P213WjSEPsn1PDmU+FtDga5nLmtOcnf1w7Bffs3zFG7DcJ0hANHvH/omC9yCy53M
J8YMEwz7fShhZCX5qt081rlTf/fMEZcLLnaIFKRy5FAskhjjSlYc3bRst/AqeiI/
1C8d0tGkLxVI3GyGttn4xKkHF8phj+cClTfdms/XOwkco3eFgiwiNAMtj0+xLJhm
BzD+8ER2i/BHOP5QfKKNrYXLQAnOGTdM3mZGAk2WvQUCGjoxjiFJHnvqDzvkZqnG
XTkeQsLw7XmDLpYMPFwOUbriiwIsmTvuLcDumnTFTN7e/snE+XTgYhRy4Zo4mLI5
aoq5IeXFta5Av7lmD6HN6t97MuPh8t1ppx/2vyn6neL5cWMrJBv5YFANmsj3AM9A
nscH67GMjyrcrcPdjGawm7cBaV5n7EtwYQdiPXCTJlWEsC6n+P5ysjGFaElIsebj
/QT3mrl+JLiOijqk/uGMJ4s2W8qids3WO+cCpso1zPzh13Z8bTUHGj8sOoqjbsjr
BY/lJjbaQiO4KnNt/b0CUFhMTwxlnVZeZssv0heS3lymhpW6U8OJHgyd4XkVYvuL
EEBukJDP2LX+MTLPbtpueq/XM0PAcyI1T1QauEMIgM/irDyKjqowxXZUodK6t5u9
3djd93INUfScFPLzCIKm+HTtB0d4J+fwNAhT/i0M51U5GmxE7GdsIemeO2sffZG8
Xsa2X4C/JCGEDzNpLrqSaRbBgcUVcPByashutq4C+Hpi6+Ksk+yu0txejDD7HMRp
fJ6dRdlEkiyk3gBGf7Uo/DG5EdzPv9oBGOuM/PH7czRZrjZ/eKGBEmodhAPR3U+t
XJKKvHpZSdrah8pu42JHR5f/UEhTOE6PEzxEQO35An25HHDpXU+J1ssOpHsNl8wD
/JL5t3p3RarDPFaPBP4eylMhdTkeleiIXvcThhynu78HWdwt2N1QHn4mSZiTpqLX
jGLp3eleCE0eWCCgPINPDazCXHP3oa2gnwhCwU+P+bWlKn1Unlka06n1Rf2hU7+p
GfKx9CvfsdOXcSHLPKm6lUQhCRjEajpD0R1++H7sQKrVwG2Q4FLB3UB/ElAZgrje
Yy1RV9CJrOM5LbJo7JDqzMkUNTeZdh9w1R0BclEwnbRrvnUoa/t2ydnBh5HBQLtn
a4erFCH1jjkTbnq5n0prQYPyZ3YmNcN/xp1DyMLQJeUVsVCp8cFrtYqA9GT2WvxH
86R+8UE9MCrCTRGdHgzGnIAijUWUpKjxvxAIC9W/VTKLtYAlADcFIK7w53uRp5zn
eqrhwMkyFrKPH8HbuII1+Nb4PN1bVJDDWWHltH8yDd45r6kdMbtojGzs5jxJ8HBO
+C6kOo8VUKef/KVJpMNpnAA81RzAhKzKIBj+rFIxBFkuQP4SakKlhmvgDtsjLwcg
uHjXCacZqJgdXjBc2mW4/ZOOh8MId6F5HqfZ/M/0rsCeJ0pgpskC+Hp5Myucee+K
3sORSGCHuWjPEe5VrnUzbQ/wdNC/BEf4oOvNIy/EsZVu8GQNMHUfh2Bru7T2FH+s
y2i/xqbHGj07OsaUNrj0O/caV3ZeK1xosN24bwly1UrdKxo4NAaSUCGfGdJfboB0
k5pR6VGnbNups2F0oo2yvntYDQjRmp7rq1cCNbpxDiKddIE9U/uuiXTkj4OnhT4J
EDfps8oSjLO3/70BUXjEOHX9KoWV0S1kmDMtZJIRnrNXf6bs4prQPZ2tcoO6FETB
oSubM0ZfsZ1d6cf+y8CJ/v9dqBOz72x/9dV0EkC4G1H5w29Qp+5osBn9qllia7Uo
HNluNyR6/hHLx+rRZpTSeqMP6tLSswz7WYYNVG60EhFB3Yj7hoRhrPiBvI/hXAck
1XffYXSR4D7MLs9Pe4sHAu6D6gGs6KiIu6pqEg8YAN9684JfZTMe/yrDp1uqx/Up
+1vCfgbz8m9duh7ALWAZiOH2NsqjSRtqz6G1a+myr8+n9MoScuD/fqwYVyw2T6eP
pO4R8lWh4nuPPVppnX9xw1A3U8d5Dk4qU4trV+Hp9x+ambF23a0mBYW0AZYkWrOY
Qt/ntVWNkeXgpu7MalbWYT4AIN6hRDXWU4l3s6W20Lnp8MZn8pAw/cPnxRw4UUKN
9xNp0x69vNqDA9ESoA1rPProfCyncYqz8MUk8zjWyXGw6H3e/R1VHfQX/lKoosO0
UVtecPCeE7U8C8kTFSZsc8z8if0FSsvJwYQbxz/coJK5cJncFMD7ODaDmgr/dMUc
uvNc0Zt1X0Li1scYLS9JJAxnyNDc8x//ZqOVJvmv4Zu3XzeRONnDHUTJAH2hOQ30
F8vQjq0WtlYJdXuro7ndi51wBrlIbD+LBCZUOPk4Mubu6VOCh/PpIAGmsPYq0tse
TFfErlbTkLs27FbwR/FKB+mJsyi070lTt3hr++BWnug25YLujKFghVyGdPumyDRE
XWR0jA1qV2n2h/ZnOPmvFon4N7zkfAIQRDEddVGKLlnFIJTIoj/63wNy4moeL45H
hoM/3gLIIB0rjfg/ylF8IZAvxD6hi1AaIIlLFvKk6Z/71bqIE8skWfXgkLbvwjkP
qhNAgeGl4zKNEGaC5VwlGsneDwUOKVe8qhp3SY7x+M7TF8DPDQ66E9GONj/bj1BX
xSQkgHBzmZuinx0/khO405ICEmg/ZHwiF8EIiyEQ+voTCiLwObQgz58bdPF5+5Nz
DZ81RCpxs79s9RsP6KPUoadq/X1weuABNHHnLfv6NUHK1sLCJP9QwcbFr4QaA7Y/
2K6u9kitdcDLNN+m3gCGqVpjNTmhGZZX5lh3+uZA1/NZnd/T8xnKT562y9TzdoZv
sI+Kot60PGot+ttrDwIeou1qnqrUw7C05WA1//8h62VzPEs6AbdPy8+LocHAn1Hz
uG5FXtW/a6Zx60X5vOBJvzFC7duq9xLsKRM4XAKlIK/8KFraOTGnerZQGDvCsmCU
JSui3aQGpGM30j48wUk7gqaFAxKGScXpYY8poOqaz1jFjPOljfAds0lAyLR2EZwg
t862hxUCe40XRO4jD2+t+7GtrLpZlrMDSf9BqF8yTi/JmVoAvNuvSKwp9sdisnIe
c8jn+DtTAnWGDbAhbEFXKUekqmvTueZJlqbDgTd0LU8/bs1NsKDfRkoec/2C8hyz
NULh3r+N/ofVT0UTBBWPhYUe5Vaemp7ichPPl4KitYP5PP4QoZUPE9fscVxpF/Js
hAGFvV6icliJY4H6Z4k9Myk8dyj7w/IVyt3ceMZr0KAVlqqZG9xNltAI3CvtaBPV
6LxObpaVuul+w2KyB9VAPhJwyv4y0Lf+qwLrRzFCV4XJNX/w3XHQrTo48eJo1Tjm
oXpnSiaKLbFu7GKstHZ14bydxHEmbg+jjit2+8p1I+pyVbaWedRpnoHkR4FzprBR
2Om338v2yB1PQilGVEiu4QW5UOu4VTlI9uTqPSMtF22ubmAgWE0X6MjfQlAghE1r
lvPzOBsqos9fgtMUaZcYQohT0pfP6LykTozz+bP931EEi4b4p6AbvCTmyxbMr6Bv
uOV1HvbIpCRnWYx0Wa3ZBvWrCd0dFnZVdbgjkPOjpxXMPl+rKx1zM2G+CzWXiZuj
Uz0zsNSEpNUgydCnCXyFVOyL/qlCoeRO2L4M7A/IH9wZoqIWFv6y6n4qKeenq5GT
5+T8n0llp43vHXXxR7ze5XrdG88zuyiK1xPuKSeNh3LxGRN+yFizC0GkErVC8XJd
+Wv9/PfP8yC+LE1HFqrlo8Hu6EZkG2FO9xygBgE9rrNdcQdJe7s+rjY/rGLhNVKm
q5jIHa8UCMwlKY1I2pZ61NPZ9RzqDVRrAjynnL9LF7sISKPKSzIh0p2NUORcewQ0
r1nhuf6F+EUXnRUWpM/m3Gc8A6KQQP5qHV/wxgweHKOTy0vX/xuzM9C0DlCP/6cH
nELNIZ/OhzhReI9fuew2umEgE/lKJieUpYH7xV5cwTW6ktC12gvkZdQu/NenkcMr
ePukEFLd0FlRUDusMpjh2clOLwlRlqlXyyz5DQUgRIy1XuhzmRigX491WXT2Rhw8
x77fRT5L8dFwk4k45/se+ZXUK64Vz7ahaaqMkjMj5dlxuse5dxDHikYSdzCDaEUy
cHIbMLXRDNnPvPZk67nFTUvI0DEUzMtQx5GYjiDXUYMYZb8RjTdf20Rq8UbyPlHb
VXp9lXuBDxIacL2uv93Y6jhc/YM9/aZl8fZXA1evcirYPg3Dum9vX3h3ryJa+Qnw
vHeBkixhFLUc1dDpofq22c2TT4hzBMT5IjkG3qE79+BSvJozKuYK9eYLQUuVr63b
R4UXtKrEz4yQ6j4SUghS2g0G1ctrFeNdRJamVjY0LheX6+sUE1GsB3iklGpWe98E
Hj7jBXscVLAVJN/x2EGfvBkv/Q31AnSmPLnlEKogQVvn9dVeWo91ZayguyZHFd0r
FZpx2mE6WWniKewW/YiyTc99H4CdsSboAPD/h8rTpGC//8bJzM2jHQng3CeoGEbc
AT6+LgKo/i8vubIr15MffGyy7fRJWgVynfUe+daiO5qLZCcIKcq3M2ESnCdCCwSb
DucYc5JEhdb8wnz9uqooxy2a/N+sQPIQ+UsQaiJqL1CxiBSMMgmHH47ew3TB9T95
9TAd4iL511iqagOgYrL8eccBwAumyobUpyf25WQJS5thACGw2WIpRaGpZYQCNIQ7
CNYx2PhdjtC5zbO1kBOZQrcij84GBpeCKE9SWYEqKoaW/rs1B77SBSCMPvelHqJY
2tv4mT/1gxQFhiyeIVWYv4Du9upsmHscpQti4bI6zWWaioE02CKRniQTwVtkM5YV
4EKVUHZKNCQwwTI6Hc6tMYrA2EhtrWVEEjmeUOb76KyLq3b7bzt1wZ53MwlFXsht
aFhtcGuOorOFy3bGeLf3vOU+2s2sxG0sMHmFf/hwKiApdVILbHjkpaG+ECjCvm9Q
O85J/l5J62kBV7/nOkUF3QaZyWVsSHAmF9LciwfmlEdH5hdEtn7UG6ISBWRP5GD/
SY37Td+i7vwZuz2Ft9ydjyIL1l3ycT4q5BHVA0aizxn215U0YF0gFvrQCMxiWNcC
vAqBzLS2LfWQlEYp2FMCgc2VFwN+gARSDX5fPbTXxw52sngAGpKHTZWUNSCMJxu+
4OVEP1hy00Ti7cn8H3MuMYEsx1AdgBIOS302h1Uxrs221xEaLHx+D/HGRJZMnMoK
yFmxy/vD/BrSEEMRVtAkSwlgzMhUNvEBLOm28qWFKPON3cZtm598RaxmuPWKjOXF
vl2C6S35+VeKfzJGHDdv108nT3IPQGQ08iWgm9pzC+vlMDO+xgTIrIe3yjn54IUa
6u5Y1a2eo33NR2EsVhn1R/LmSuRbfAUJDujtUyu4HaDHDmgin9dFENqDGeoEywEg
w0qtcPsXaq6mMkdtAYZ3AugfDScSL/Llw4IJtktQ+WNUKembRtZa95meBFtnS2xJ
FyE97MNzE6BYQ7tcjoVYQukUtRvmRhHKvsBPBC5acErSgarSyox/uEjJTIb7MCpN
6R/XK1N625hBlgY0zbej2rk2zqGY7siiHA+PmsaBImcHsXXj9OpL6XcH5gv+Yik2
Kln/c6J7rPtUSr8RBiSbhMi9jvLjQ39IZXVJ64hODUW+HOyT02ORZjHjp3Z+a9OM
fzelqXG6/6+h0unZ5K51XCs2NEKEK+3C5lg56TpG24tmVy2AaiyZhlo/IzeyjWD/
hmgbiX+Ori3NThxq/jQh6qSaEoxeBN1yg2EP8/1ldCtrgwDohUlQg4nWElcbVhR0
KaxfODQzE81rXd7zAplsPfy0oIR9v0mcGxEs14nyNRlZUAt64Jv5OXljZkZMM0XN
oTpTIuOLILKTiWCm4z/AJV2DJutwm8H+yiCKb5M287Y44cLiZnUId+WQ6mcyhDwJ
5fUMg2OF09pNl4rmhx6wmOl1EAiYoL/Hv3CeeHllGaUGOIVjWtMcgvLmAaVQkwR0
9A5d0dH3EEFQtceBXXNDc/YFNCOBoMGHjeMxhQX/hGCbjaGug+JJ0qf6s/iPpCdN
/2zUZTwBxOmXssqqDVYCiTV8f7wYuCf7nz/RN8COSeSdn7U4L0qO5VXkN+XBtTlV
fy0qedSYXYl1ZRahC+wncho73oQkqLZNgg3Yoh/9RoSckbwidgixbZBazMqEdccB
vYs/OKnW77mITiIfYPRz+KSGexsgtHphiKw/FWf82zgsrHf0iuzc+Ts1XOIwHbcP
GLFDT2p/q/pOj+TLHfsqn6dxrpFE6eFBR8QAQurz2SJUKxJ0/jvpZ6cxyu2fTRnr
C8GOETbkel7CFHVkOm0H7incITVz3b+nZCD3oguVpIcrRu3uzesltMTrSZ1Wqi/2
yrtYmzAIdjHZJgL37UBdUOFg8+Jgz8pgVlI4zkcdZhKAYcgdUB2q2el/AVvws7f3
Mh4OmEjzOWsBp5qso354gcX8KH08JN6cvlbcP/wx4xDle9CfBph0F+hxwGEkh+zk
hzWI9l57JJcGkjgSenHYLI4FW9gC7YeNoiyqF6T5zNKn4m1gpfEzTKavFx3Frbrz
QJqsQ8hBvBDQ76Q4lacwn574sGowK5czgRAyfXJ5mvjesnJgEcSvC9bjmMU4IOis
1ddHX+4N6jN7SoSICtPyOooIp4xUgFos5MMwiS5feph86EEy9xVAiyLIXVjGyyfz
tq2hImNYMxGKciDK6n8RvJEm99Q4t9FbZKvAGOyo+kKsOfYZY+67MwYMCEBd0skU
iR+ejicndrrCnq9p867ylUz8Hau/NVTSHmZ0qYsHvYxltFSGtWM5lmHiU1So+4aD
ZTMYuE8UnzSzh0XPQLUJrLH2TA75wd4LwYXc8V19eD7QKBXGypMP9peBtYblip3x
AiCZ08YstD14tgVVOt57TnNr5IbFSEGoFkdVRw4NaVZu8SzK9WTiUgAJ7kOEmH3y
SNqsBxkmi1Kl5KiavdNJG8UckW0N0RkoxITDno1gX2RWy0VkTG/63WlH5JOq5yN1
TpiAj2mI3FKsgC2QAnhH9LWfO2reFNi4gRnSjWLGpcAhgDs6UQqYMP8yXelGJhWm
jYUvizErVAVmwvqRCtWaYmvj9QnoYHVDb34YneS7AbqoqW8jSiysZJkjiF+1iKpc
0xdJ8H5/2Cx2n2AxgCAjOrzkPhea1yCG8Jzx9JF+0SODZ/zH6IG+vQUXDIBFKVNl
2UO+BFC8r8LTvp2qpti6PkG9AqBHG4s6TRjpWwZwp0DexVkbFBU70BlaF85ykZIQ
Bcm/0RxBbuFeSQoEVJXhQ8libCTygYgZbTaV0So3J63t9TzgHL3MX+j55C8mwM69
a2FJ7+6vbV9doUCwZEO6lCMhuXuE97TQA1wt6cOOAJnZz9Wuf3mFIk7vYpix/o2R
M7xVxVoKrYeigC4I+vUF9BuZCIn/9u0HAyhnZ6CzY1cSQx+0psEjKxrlGAI4pyQ+
2fcCpN57Q12gp8UsfP1gskrdWd3j2zMOvOd3rz6WJKTnLDtUlcZHqh5//9Crdysr
PFR34VrfiONzyfXW9DnTGqM+LSf3TI6vvVboOFj5sVcD1gXw2qh8F/0z4Mptl1/c
A/YmjzABHOXctxYP8C+o8ddT5tWoea3BhIo4FyRYnG+RWySkkDsf3hHptpvfVSyo
sZ5v9YgmkUwIX+zmu45KMsodFpOodenbBygDhB9R1ecpsQsKTs8GOjO3UZqi/d9S
k2zSYVpPd9ZbV/OZwed7+laGIxcpo0iAxl+05inhY+zaSeDXjLG5pKZvVvDCxqmh
8wnLSDNFS6S++r0Eykuq1Pi3+93N/2AyCzzv91p441+sA6O4lILRtqxWW2nqlh5S
k+ezcoreTVKbEiXq0y1sFwU6V0LEY2vzXJRWTWzq68oeCX1LFQiajMMuEeldbbbZ
ZEkzEdGBzHjpwJ6rCJ1Cyj13DT09hBiKIzh+qZMQ5TCb+T1kUQz6ZAR2uGmavaGw
CLmCNawYNymCx+HfjWbxriAN8yHvGnjOCUdGiVGlZrBG3ICDSuI0TZbPqD22AZEJ
9tqD+w8GzfVd36HKRtv+w69gX2dKhs4JDJkPhQcstxT8XxXcdpG7hJSfhxcRennk
LcoVrGrTQxyTGADbHpWVEZMxSY8B7lv8pdm8CSVsL/5r5MtpORgRFJdzS5N0lNt2
4qNv/DDUBIbS+T3w44XBA931sIa6iV8zDw/L4KcKq9q/v5nd0xtDLP6VCkLRQqsk
HexUYAMxN6gpdI61rwCbkhvIyeAvc46EUqku6SBNqBbkmNO5ZIDbSpvsHSSX4yVN
DIxUo3TBICZm9dfgvHfWL+dMXYAOICuSFCGYF3LUJJp6EnveuNbqr02r2qMHmjto
V58QuSAd02kLx+ds4hLDZpwPAIFJgDGMII05LGOzys+FmAWj/b+jpZeUVRWUvZxb
j3jYSoFP3F0cTuourYg4L1oesdBT+gBSqRtaOXAx3MugtdKgA0+UT0rSd3A0xMyD
WZ0N1xIcFrHshMiOaQVk4VTHiV/191/Aul3kWnxIT/VAiCxnsTpnR6S+IEtoP8ii
EthDDrjIs/uc6bfffU7f33txBYXujpOJpFPrcrjtqGQPuBVZj1+03x3klY0xqOrI
PM7y2YvWurDvnVR3jdNCmR2iscX2mq6lKcuqHFncdtD5LA0bdXZXsgWEoMcVtHdz
wVSrVtVz1Etgj+pdppgsujS2f0cSaP333ehCitYa8UxAX+buXQQ9QPE8RaJkuZBL
2+lB2xk20EmIFbreQkMlhxjCfRezwPJ95gdFC8FcbcIh2lGBQ81SDlCATB9lsR9f
/Y20uKc7/OAJDuo3uz4D6JLdXHT+OqCZCbqanxB9wSP9LgrM2CvHdGdkQu/wq7hr
/WG4iC9qJlHvWpqtvf8f5YWe5/rvGCtOavfSKcHjJj+zizdbiabXXe6IXEZPkXb3
HjJopdZCfFcOvxBIscZh2EkKshRwMyEUIbeZOUGfk/d1KyZKOIGs0ZU5bFjtryd0
hJIx++R1lwU6OAk+a5WS6ZMZuUNdLw9uVmaF9W8xU3z2QF61UFMa+mYfFOFGSUFQ
EGUGS1LN2iJlQWDKMvz6cLALJ7fgEYOXOY6Q+7ZIL7Swr1srWeC5DVpl6PpRPRYM
QCdY/+s0mI/PrZl+aiYTgoKastxMmYlx6wUUOza8AibIN2s+kRsIF4woYYHy58Jo
LH2F8EtWLALsJwlYeKqTHAeG2N8yaJdeqrrIVvTecSZhlXwBQCl/pP8Z4q+hvpEQ
qbDkBPFH3sjBtRE9XNzbFrTZAMPbc/qSXTO2UHvzGxVVDLS5jmRN8IbSDIfDmWEl
BBL+c/gnL0k/X8nGS4t/cR3nJn5OEFKPqXadQD9zexw74eJOVy38mTfJy6WFwazi
TaPWqdg9HY23fWWeqPuReQa0eXCVAQwO1gc6DbWzubPqerXy6kzm+BWp8PQOoGo3
tyssOFI8XyIJ9EgiHTEafyakqFDHH0l3VeUneVuvKWS6D83zRQrxcEBOG5bQoDk6
CnO6FNM6rirrME8RO9MtER/boB/Enc7Dm/3201zrsUAEU1AFfvyMpib1mDH2E+ZF
yyoy/C7dm5j774Z6ljWA50XNmP3GMHbeQLRu4FIqZfu5zPvJ6qdhSx40NaNJs68/
8xIdveKjFZskgbo1PrETjNJMNQZEK6NOrHV2H8RLWGxCwEK9+Cs4rnr/zl1KQs7y
5w7N7qYfkGb3cbYIJcdHzRmN/z4gwGICHK8gh4tnhaA1MRm/dmk4XsF9iO+9DTmu
+JGbfvVG4ido8EVfZLLovLmghgF4+/uAZH1QdmHPYvmG3b2ZcSYwCYzD+XSxr7Cz
gM2kNZn/qk6jQPAA3fYWfF3Vd01zEqI4yhxGsk9BXIZSBvSs4jPWOw9kJ6Bpykzy
z3lTVgMtGcdsCY0XFe67xHGhiqS8rKoTWNOmlc87Z2vH7VOG1OG4fmwR5Wj/IIRX
dWuL6IX+UAOgRRTD6aHrgl83FXbgwY4Z5xeVPK4uwXvlWhfgjsGG8x6nziH5Wxhp
6eLaSiTvpmwHNnoHTUWBl71Ul+KkIM1rLhFoJN8YDIj9exdWZdw5kDZ1qDYwLghr
daxM5MWglkz3+AICYtgLRx+oxRuZFDl5RrzlAosroNTOJdCPzMcHpE4O56VuJRxa
eixYEg/Rmj2KMDTjQjo+RB0KbkEDXVH0B80Hmga+nxJaB2qhMIJEQufefMr0RYME
xkGSlbhWTee1G16IAT/1Bq0EP8woqpClHmsYh3nCUF5RC3vR7MxILyJtNnbUdEfq
9E0Tz/HtP15ZHy0Bd0fXi7EGkDOcSCbjyz+ONKxZX43VOJCFNu5FIsxhZXS8hbxj
gByPBMt6z1l3CeTVf/e6zbC8OOv3Pvf8A0z7qjR4Mo4bQcOtOFxxrOKyJj+dBD+0
+d/+Iz7sDxzbuFo/JG5NB/FoqfHJBhfF5xwY4aucqVZ7TaeAFD/T62L6tS4nXnFS
+iWfIylbETc9CKP/AYt+v6KHWW4P/yLpIomygO0kKX7bF6s8jOxNb/pk6njJxeg6
u3W8CRtvGYFFnbWooVMZa18lyrHaZXBEvOiYVx8Ee9ZcEwceGmjp3s+VATpI9M6J
yBNhYmxpK62Fu78QvVnLo6jPl/bDMqxssYJWIq1R6x7zdzZfc793mpI+geDPWHHl
FjipzvDJMFLY/h80gsHfuRvxPOlU1BktfRRrIJI/08Ai1Qc0I7k88W/uG5+zgqbr
uIw8QaGrF+RqREPWkbr/sBLXLXbWs4rh3ZcK0p5B+CtLEWeQg5cTNa4uMHtBVycS
tDOhD2no9Y4cxayXcO9cMH9cz5NeByb55JVE+DRx+ityyL3hNvgqfpk4rczUfZNV
s5ZfXreMdmzeCtwchKSTTdsMX+mJNpCLBBcLbLDH4hfHgfMTEdUhFIdK5SlniZrr
92MUVFAtGr9WLDSgST9lyOIdFjEsOcfAhVSasBhsrYPZk7UA3GNqQvlagLdtscRc
zW3KeK8wLdi3Ho+Qcy28Ro1H18LcKq8g02Do6605oJzqZM9cmfoGEt0/QuLrMi7r
7tA6K7LvEvDlQPyIHPiKNqv/PE5ixfwDHyo/l5i5Ev2SedYcql5Sbz2PzKlBw0tk
zu/PcNMG/2vjstHjgv6gAIGRHMLruzPw2LHKUKJD8fITbd59Lcu3HYPkWnXAM/eu
pmwJgG4sgr9zL5OfiQ5R5CiIY/1rVX2UAt8IQOQf2XVbnHLHohFI6Dw/3Zsk9X4C
tcAf7O2EX+7+5TRDjLzsyKSDjs+s/0DXvDequTT+gS/PktOCnCXMbYyjq8KCeUrZ
jofv1jqLyUSPRzejQdZxxnHZ2qVrkKRWDvqnfu9BdSKZjrYDA9XH0dOqoP7Z9qL4
biPKW84OsXqnPIfhK1qrLXGB6nZYircEbl+v9dr7eZRk2B6/tKtAsJ1gnUZC52Y8
LbXRT2y8285qG2vdlzLN/5NOO8QIBb5LBKVnqsE+FgCaMS5R8YzfWKnuz1bQU5ra
CoCP/w7i86cQxpnOj73CE3qFfeG2DrU89eD06bHLDHwjeYZCnB7pk5YiOi0gm8pA
XB90km9BnDr6FALhrtN50qSu1PndpboVKyDO1oj8Ee19HKrRm1cBUPEd1JxBsG60
2t96R9N0CDxG+UB9U8DJzsiXQUe/3el5M8WS8RtZPBUQVLbEyWlatsK5a23xjVQg
hcliRjS5sIHvED1A+DgV1SgUN8p1bV3QUC/3JZuTPdvoGUk5aATffjOsXB6pOzIt
tjf/NoSzBm2uaEWBSmizYDNdV4tJNf+BQenY0VIVdPRm/wYXxGpO5/sseO733nMx
Uyqf1hfRs+As0kc+p/9P49EyCCL9iFZRen7S84mA8ydOlOlDNPfal/UEY1rbMixn
yVk34IxW9DHdUBZk1MxGn068qSEVPYF1iJ1v6l1NkwCCwRIajZpLAJxBOL4TZlTA
Ogr18BuftjCNEKJXU0Q7hV+eBo+hPr2/6HShlp6oR6YBKmiuDb+MC/ulKtT85a4W
CcVbQFRjON8V5mWrEzKTtR3yYU1DBkbDkNdsioub35KT6X4QaenPHTvY77kx+3EB
3y93pp0uJQtXKTZQ7tDOhOGIA3mXVYc6zpPZFxKbAwiYfhzDb2fO0gleXA7OvfTM
JWjd4JjEyOKSPErRzDvrvJQhhXUvjWU6qrJupgHpTLm4tusBmvH9nSqEW5fCYHwj
96Jvm046lbyshqGE+nD+PwrX3hN7keVnIQ5p3nm1ZAfHYQFSwePyWJhTf/e1GR1z
yKFEASuzSoSr+wT/QJzUIqQ7nxQwZxyAaiMXEjOB4wshwGN5CPBIgvd11NhX1Hjk
OatYmjB4eBGhBRICO059RyORv3E8ltHhXjQwqUEvUg3tfynrmtqIYuy4uyarJlhC
QskmQRtxUG897BzWjDoqO/pZR2ZDvPvzjNwJU55foivVLjrVZTxpVt3+hhqTXywT
SiZwkXGGSCi4mb3HSmLmiV9b0wA834BkuPVCbMSmBlYzIn+LBYY059n1U4i3GNIk
18U/bwF3MkqPgxQ5VrILTdxiR8NVl9vMnp55rwXqWNSVmpkuO8ywJB6mI0QjF9se
Clqz47fMjrF8FbODCnNkOtOb+s8uECBU5dKRmNRIdLmYgFp/KG81zt9aW6tIna5q
2Xo2ZxkuQF58gumf7UTowwkut0EsJ9KCvqJ8WbWfqNMxMMlYVbnoZydaASKYSP44
+TjxQuW9EyB4IlZqn6HYIKgbC2qolDokMGt6kvdZnAVoxEA4FbfeTyme23eDJaT6
cGHg/NvwgE/2caPGz91rmFVRygmiWjNu+8C6HWFBNKAmpY+l8ZiINgWU3Lbgdhag
dJt8fa9slJeUUwTlNoVxbHtdWYQRBMug5LVkRslID/slpYvkdMuqx6fY1ZWvelAz
M9b4JkYlYiexLzTMo6LLjI2vJTie6222MHDvZP2FFOKobpIihUxWNEUrwd5vuHrr
xYLWVO7yeBpw/kbKbHlVMQh76vfa68ttz4U79v7pS/OK4zwY+U8gkJrLr8HO21QM
qlMtZD9GFWz5OLVQ0kolhIQ6lCIFqAK8PJgzCGUKuAqJX55MyWFQdFD1eM1KxJT5
g1cduPUIdG61LSknUMsIm3dKMYy9ubhyDYh7PW9DmCpTtAhKwKq2qyYHQikuHJ0Y
r+GogzV3qK6iWgCfS/bwN06xE6ZHdNhQLAYD17J6A/fMDmYoms8iXvRFeXrOpvsz
tLIEJRLxEeColRpGYLm7s19B39PwW0nlZmTHwqZdxaxzSScfKuTl2qm/0c5AXPVM
GtN4WO7JJGpu1Rb3dTebpsJxzf5XT/n17Q5klCsOBW42kOlS4OlB8chCy33CTAwa
hPGhpvWzRhz2WQWPKPXi58BrkGB/a54eLAUunx/HlTmvHDIXilS9FeDrgODhs5wc
52gYR0d5V1zD7E/e/ifAxawGyVI/qJgni1Ou22vJ09BUA2OvBPLhqZs7nJHUSLn6
XQ2sbBmQ3NzjI0nEG4XLo2tboInHQb1dIYIavLK9C8iGVvCWXE4NhS1LEyRxKJ4C
tFgy+TmIaI60UO6tWINi0JabUbTndxC5kKxoMowWvVqYx6vbvkp7El+CZVWkfs/Y
nmbmCCajJEU63pOq1OWq+5H0gPX/ST/Fji+zl3qSPRg92VJ8UD/t4jHeGr6CHHGS
DUuTGSt1lHmtfy1GjkjrYqhZdgNxkHeDZgj5Flx8OgbB2JT1LmWeKChMXsMuMWMz
w9dLSNSLJ9FCs7w5r8p6e2JGaP3olMpTizNeOVipPhyKEvx3hHTT+q0C7M5WQiNR
AmWjiaQHy9o2DRslTAnU86Xdn+W6ockMw7x43fJWKIsA2N8BLDN2xUEbUM0Dzkyz
+9c9XGP0/KqU/BiYxR43OwYGrMw/U5Mzn/y+33suvqNkV/ubYCuLjMFW9m2U+j1C
HYbEHmdli27DGmjx45b5z/kB0tMEBeWpN3GCTsZF49XYrskY83/Vp8xs+glBRfyY
6cElzozB9959JGbA8sCOL+Cy+dGampeIFd+U1YVDgsZUU/4DiujJFyFPZAja+l9+
iMYk9uiOpxMxdb4JMDpLoQ0ca61YR5+J2gibvsmpO34kZx/YrTuP/g5LQod6CDo1
l4zofkHnCsWpGyDOY/SzlOH/UgLRq3Mo/1fqElymo93Bj1P7WUtEnoNs6/czM705
64bOVZEJxX+oQ9jek2at65GivKuw2J2A0LL7r3/I9k7j8MZJ1X61CIfFQT5T3LkV
LWYlaRsVMtaK6dM8NgeR+qkNP9q2tt/ogjKVJMdLzoJYzak+jXeoMDC6gwuGJNSx
1RrY2l0x4rLHU1k8CQM01t8l9Ur9k8xeA2q1besJfEaXbTZGKKOwr4L1o/DFBeYn
JcXDrOkX4X7zMeOF5w8Jpnq3eE3DTa4j4n+RUH4shprU3aOURcJsoXogoNc7dDPc
kE6TcTiuVCVcBYghpc0vBbAC2O/alBf1sjHFjLCb6sry7jsyWhox7dmeWFqHd4Fs
HzkFIEdG1Tx8WU4Rl6q3P9ENbYROHQ2oIrkJb6azx46MnmzZXg8Da6FpiBTj3kAT
ApDlbx0LjBq/soc7sYHnRovZ9oSsROTf4PuCTe8EA9AFP0BR1glrsxXiWXym5o6H
jQTmfE83iZ66s8j9+82PkwHG8/yl+Ih263tfkTH9C8VRa/00NRLzAxkl4uv8E52b
UsUCBTKnto48bHPU83nIZeBOiZnCc2HqNt9mEykc4lZil9+RZ1a/7kOKciGB1wXt
qr37oX4Tc2sBrQ4aCjq5Yy8K8gyg3W5WLedLH607l2mDSsoha6TUefLAgxc4akjP
Im86toE7doreRpbqvAzMN7F4RbVO2ahyLqROD+e0gqqnSAQQzbG5sHevlavDkfWK
uAjNs9smDn+/8KW1xXHhFwnsRbSBL0C9X+xt43ycjSUAGcHr2AZ5KVhRokuPoleM
UUeRDBMNQ4DS/EO4+BA3T4CDfK16sd+8DCnGqJPRhiwWWCB4iKmlSGmQqdvUz+cl
IIomEpiVljnaUAkYv7WU7MGG9GQX2lBx3pu+dzu4leTfBDSKxq/lKFoDz7GuM3cz
g/xcN8GETuXI8C9GFcI73+fShAs8nJKD5lS3m6tJBUNVXtd0TQQkdDdUVVBcAJz8
UmbXUqUbQ1wwzFubGkyG+70aL4PrxdgM5pIBYxRMftNKGGyNE+/HZRV0RGkpqIly
kl3YDGqNt2M/QliQmRjBkJRbidizZgV9T/j7xrreUKDTG6TXD84YP0+XGc0wx6aZ
MuF3Tx6+ZyGhkpm/SplMmTKfEpGnS6OQNFC59Uh7Ax6MbvaEFz0nO604BHV41wZk
ijDV2ra/L2nRHkPuybzv4C27XfMYWG/0P3S3hS/8GKirNycZtYllD2hQs050egaC
rUVWiUEXPXVs7W8EgvM4wKgWf7HVH1NijpyzgAN6ChQiY8GRbkZ4usCu6pHs6YA1
OmKwNkuVA1XpUdG52rsm1LIMzCTRm6Y9dG3qMMPF5PVgQUGONzsGy8GbYa9XVuEm
cNCk0Ldhhk+gq9HNWxixagFyBt5VBwLmNj86UzLJN5R4YzWg/+UZRVHbCAgpXyEb
j7ttlOVxYptmXZLVkHfhDHq8dfpZMyIPz597XCszFeC8qRd4o1/0kSpGHt24LI4C
sK8Xpm+m4QyzGoiu2RMaUmesR9oUMMypeyMfHv8VF2z1yURFMzUMnOFJi5megrZv
1yIUkkDLu1xky5yh+sH46eGzHopir8hS7ckeFKwkgGVf6xzgAlHpy95XCdz5ZiW1
B4sF7j8xqVgX94ik+knxBXfsxKLn9UV5e93/dMENmltEQrHgsQn+ad9ar6yeq4J2
V2Rp00pOJH2PJuAZMXVOVEbtWZq6uLVB6TNjYDZ3cFR1/XQuX/WGfOzCYopfVBsZ
bG5ZKiszs88qly0CPP42V0J9Q/kKM4818fhXwXm0Ikqnh2ye2Igxc6wvwJgomZUA
sW8tM2pxQzyqXYw8sXBBK9Oc+wRQDtZyrBq7dZ8WzIrQ+4mCIDppD81BG0srDU8B
Tp3FTTt6sZNy0psml4kbJqtf5enb46cg9XciPzvGnPyf+PfONTpamewvA5MK9pBf
qWLKVOHsmS7rU7HVPTMAOg+PqQKvRM5oS/QwyUTzu0YMn+6zfKpHbEDMo/4PBdAM
BR7ORhHIxNKkrjZQqBvfUIHMRmOKQ15Hp8ZWZDd23MOEitO/NL0CXfXz659yabxF
gmfjGSTjsFA26Yhp9jkXeqL+5yWlLC9nv1Dn4goQwFn1ozyV2E29C+JDE3v4/rMH
h/pi34OnRFyDYUhdJEJBTpOPYHc4CmFYGcfiz3X93w6YP82TaaLTW44XvNeZ7jEi
4BvC44rnxXY/J5ULE7RNw1Y4l3Z6XPbLFe4vOM5Lb9jnwdZ1WW+EE2XoPHIeBhAz
D7rZ83Kv7wFZ9mncVvCftP/Q0p00TvN2g5CopEH3G7jQs7+I6THtLuOhJgpXjIry
g17mqWV5PyDaY5aP4VE9WHaIHELjJJRpf41iXXG9fv1RBS6/RSe6FSYvr8ko4W/Y
9qxd7pOyzJ395ggW7dXWVagIPSf6QxRFh1S7B1vTjicjl9ePdAqdp53LJRkO+2PM
HZhZeKRjIRlB+OSc+ealfTrYNEDlix4yc36jebeW1uoo4KgHhwSMhk7oDPCjsg94
6P834hmBpwNhcBfWh1ZemgU94giYbSW7PEozX5ERyGkAvJXCURhidrcMnb9k+dCm
YYxz1aqpRhBQdpUC5+NpO6cNT3SMhhhdjTfkSNkT3pJFuJt2OVYhZZzFaxWGnJ1A
RluozmLx3R0nT7JxYnSElB9C34Btyt0Dn+A82GPTQtvUgfnHOcBv0V6wmL416wwh
7geiG4+lJZJ9cggesTwyOkde755/qWQ17ZhDygsJYcVt9mjoCZAonzV6mmzD05Ws
OAQbcldG1bmmSeizQHh7G8TURiIoN4rD4qaEYmjYqR/NCvJjtO3kqHPQ7/9r79W+
C9MPZ7Ubp6qCcQl9WWDCFK6edlaQ7FLOt3UZmCbR9P1KUDhwVGWCU3m2CPJvHNJ9
yrHddtJW4tNRG1bIB+cF5LDlohm5c5nOyPYmTGDN6u9E9XBVMDPeGtPkW6BoAl4R
Dygb3vdoe6KDoQmyG9tjIlTxnVLZUG4rReNf3Rqua1HB7mfCPaBnIStlkqncs5P2
dKUEpKdfAFP6FaZiBuyNOfzE1YiLdK++dnqCcTl2Vo7HNC9qEfurvF01+sunDDhZ
JHxOArlVaaRJgGxJ39+ejE4FamsIV2RE53usNYft+XFVrRHUdVirJqUYCHfQ8FDd
UlWQoMcqpxOyWc8qHIoxPNk1R6QZRRY/BIzzoHifZ7S4RwMobzC9h1sEbZFVa+OY
PlGCuL7kd7tuzjji5yslQatxVxbqJY7XpYi84QszSXXk4+iFFLCYxjxcbQh1df+p
TlGOtJlg0V3ZbrO8PtEKvc9deh1WUi8QrqICT98Y77a1cC0HwqxJ/WmczO+JQQ+9
9ryLUxjKJklFhYpTvIl0U3tiqRN/1ioK0BQ/xc3vroi+OuTkqLwa0UDBsoEK8IRd
dH1QN9FzJLllP1HfCNGsQ4z/Lnijmj7K3xFNbDkdNXWAUuvsNbLM7k2o+5GBHKfK
XCclJASKmqEC6jJt7M6I0m/eVf8uTpI8MEbUjgF7/J9TKPyloldHjHSax+pwnvn/
PCTA97Dror6rJCF8GOwvTMHJbu1ud8+5b76yCGxqjRmjGrUu1pK2OCJshextPYL3
O1FX8YVMdqsFRA98M7U5kZ3JFfJYyvM4U7iAQYjLBibhl0z5BCfA/6W40SiGjd0N
sH0pqJCZdy9BXw4TellrGCsw/PtXlIzh7z1mg6fdmtOqMbG52M5ciJxoI2hYLh8T
gCjps18WTTd0KdrzLSEFj/RoJ8qbuNppEcMKAk/FpNdWGgjY/NIE7aRG0JRSis54
ugTz7TJ4Y3Ppm+WmgSqm6z8jkRfDp9KomcksrdW7p5U8+P4qZ9BlPIj22QD6AZWn
5T0uxKij9Nklod4NxWqS4LlGZf2sDDIvwKS0tFFPBiEPM5EnWbEyRc7uwIQTNUsO
4GFo8ZMjshsnpldsP/ooxyAQIGh9Shoizi0Q5yJo7/pjlREhCLd9pCPjd20elOoL
dmktuJTnolRoCkXwVIaHjQkv3F8ODfnUSQXqdGlDs+9e0hOIvAGTVpWJeNtfO1LD
YE4GupVG4kU/kRXqRJTuG7t8Mp4b8lB2CJDMdv9u5GTAVJuWyxzG4P68ANGWHyQy
K2l6YH+LrSwFXzVJuU0+lzlkSwgBdjreG3OFRLZmL7urCpm+VMu9mYT0PMLMCZeN
wUugkMK1KCgmauukkypeImKLsWskF1z3LI+sJXupZ56fDi5IwG9b5PN49bW0Jd8n
Wm3KlfTxNGt8Wy6QIYkhTCIEAY8rq0HkbyDKmc+QidExEJHFgmpEVZ5Z4HWhZBSy
PLAENN6H4deqScG9qlt/JxeumadjQaY4Qoy9bkgKXV7cDoCXkvQCuzF3KqomJ0yq
JOaUbeLh9Lp6cpU3hOtbMzCDZEDsuBGWvvX4vRiAB2vSs8WSJaBAAOdNprK9pvOQ
KBXT5nYLb/MrJDOco4RD9nfrgCcTlfZe/Z05omdwq6+9hnw7xKQzJB/qbUmEG2Q/
KSPPvfDCbZRFYuhiMkgXGRatibV6aejkHWn0OMr8VPYQSwNP4iua1f3HXlQA64IX
FV6kP/OMFZ7Pvp831jobEw7/WmBOxWeaQ1jc1eeWpPEhaAJ0YZzGwgkLTDAMBZLr
VX9Eipgay28JZt3BJg2VB39JyGx7WMo6m2L5e86szd58GtQD/V+SR7Elr5t8t3rl
2xYDnjpKVh8u8Jxo/SVnfLyWzHc1r1SDUD4ge1Zs0jF4iO2nJ9iuF1a5d+fbf19o
A/EK3eHUpxRd1vdUIw2Q9usLZ+WRsapWuxakRY4UNPxEvCTevP27Sdogj7GDZYwl
i3iPwvj4G21suWM303oU0ayRIBGP6f4+fGOU312UNKwJTNtbvGwNYwZNf0XF4+Bv
JvZmQBlvMkkzAeIy8pFzUTvbBV5iDBUkz0wpafya7vHb8LFRMUOFuk+O4qiPQwko
77rr8+7t+WxVUS9KTaXSGb7uPSM/dYotfPEP9frjdXMcWj6pi2QtcQIKoRdaeIe5
XM60M422ldQvCeErQWf5tcyD9kdzBgZTHclkG06TlHUWnOISdL3kYcW40FaHYxrc
pU2tQeQoEGF0HFMmKuJDSG3ZZW8fa80mFAbxwBUYYX0tLS6XyNMiZ3tN+dOvxpau
SPNEetXE76tl96c/6jK9Vl0tzirM979NcOewHVwHYshjdUzntVjswQyOafB4bdZv
9eFH6A3S/Hs2C6McT5FWRXY4gnccXTw8mCjivFm7fViXri/4EgCjNosrt6YtGuME
dDxcP6u4H3eviCSPCFkmPHPZD2Wtd2ISUgiUOdLJmafPKNb3XOQRyo1mwsul7s+N
xaKcsvC5jWGbnkxv0uOeoPwp+D+qe3nknomv8kmHfsPvByII/6h7Pue1KjvDNb8u
MmJ57+4PMIKgVY2zAh1L9qi7kaScmyDlmLUaUEWGAaQzrCMYlrNevwV6extbvbCz
yUmnfLMSIDy4Jv62pyFHLnw+JisbL5c5Jo1mneaZDPjCSKTRacu8bj8fw6KCXGX1
z0K6CRe2/gYm2eYPVRh6Q6qwQiL5uNFkc7HOrn2L/LtQJLLdpzyOBsrhhpMGfnqE
JXvfWgcpRHP99pr76bQbadVFBDos1oS2IOJegggciksX8EwKNqK2CZXrOB2Hd9VN
4RMFOpr33CMOB4c8llfw7zMqIDqLe+YRRlHMtxwuUSKUUotYVnSOzCKz3AkEU6Hd
39ZcjvtG+BcfHLktwwr+XUQOe9cnzlYBeWy3kab/vvVPfVtC60Mdh3eflvdFW1YJ
erWJnkm2DTMEmH0KqeVD4dviGgxxf0Air8fXFBFgnfuyZoas+4IDRCmRWbbELWOf
xPeBWPV6xKk5fJZGDHiF2USQjFn09//N/1KvVq9cVuHQHyscj7yYz7aazyieuT41
FIImcp/SuMHqoFJp928GjFM5S1hzInzTJqwYEPUY5xtR/wKEQRtXQynymFVHSqjy
b4yZYOqtycFBmdSqNceArr4SM+E/wNdI+IOe5Q3VU85yJ/TIbRHM1ZQ65lyWpI4k
rj/4i6FsHL3KrsqlsAxmHjpqkGlpRxlu/nSiOMxeLsDOKShzhEZ+DERWpec5T6ge
d+RTTEvPf0k5Ue3u4ZxmE5nu9chdZRULo2Bu95T+mZ0ZHcgKP8dGffnajqE95fOf
P83oFpsRahvgQI+Hs5eMCJdir302dW5UDTvDiGO9V2YZIm1gOtWlIkSzlFe50Iwl
IQQqbJQ3b4h3YBdx4yl4JJEtdkRT+RVMxexFHUXysym5FrvQFS1XBwccbDMg3RQa
UNwesfhWBaDFf8h3+ICPcwIwcJeT5lLoQFoPG4TtNlC3t9vzaQ5oaVjGb3wqBgec
UxFLvAbgmh5bgHxLQ0d/vquxDMx7O6xonm5qc1yCQ05WTLp0+KgxOZoRBSM1a53c
wsMwsqiAFXauoc1QvXNxxCiuRoTC25ljf//8iN7EUHc25byEQJOZ5FxZUTHuSnJ1
JLhg+jFWgdipcY8f63dxclSOxS+KyFeZs2wv8iCn1KE9fBbNcFL6m6Rqxm3jngxX
/B41+5xzUAuVTkW0oeRwfi1bCCTbJBPNroTxwF0xjqeA805mx00L8sF5sIqb6tLa
cU4KYaS8KD/G1gJKefkZsmVYkzt+owS2L/eDOX4NRQ4Lc7HAxI7GPEjQH5h/0xPz
Re3BdbL92rsGLXHjzDQd3QY+yIM+pO0LSAfErYmLpd0NhNZZupvpIszJ1PpdVAiv
LSfiibYTd9mdv9PpEx+kRMBuvALQjFA2kXPLLX1WyHIDpl/Y7/BNt3lK5uqQ3QrL
KVcymvRi3Pp/Wiml2cdzQOAFhgTdFQHSNvYQXrdkmTwlSt3n3FofWXqxSe/zBXQ3
jQsPemufdkIQZOmPGdn69yz6yfvZVJ1OWrVI+IsD5HNcHxiU8Qzq8Q1NytSA1wKu
WA6XIhd2fAHkY7V3wJbrVQlft8MIMuuxtThmCWP7/DofkYpjnFKcUiY0Rt8Kljgz
sPVzEteh+QbKx+b7z0PNveiDD0Ucye81Fj0lngVMx/AQdOQLbjuHVERcANnmfaHE
wb8u1wD46IlbfrmE9caKcqdKQCaxWjg4msQsOcVB+4r5lczBw3/wOouHJSqcdwtn
shteP3b78Kwr5m+EK8NNmpGs71Mfatu9ONh+Edfu0lScwpheRHJMOPnkhEwlpV5Y
FHWNQcZToQDViJVJw4bbUjXsGA9b8DTvfsdaQIct4kY4TKivutUkqRqCchEvI/FV
Yt4Tgg6RQILvAPhR+4jpiNISEdYbNdioVop5wgWyJCLDxD6jtGTE9timqgwGKq0B
LEg6mAzFNN44VZ3nAAIZ0R9skl6+6oPEN+I1dl1qE5k4oSZ7sEEn9LxRrd2H/8lf
k2HKkz7BZh8zClYRcH6ENzzJZjURrdRle02YtwCu0jjKmqpZd27IMIfTaEocLFSK
HdNhSyRVjRlGIb0bIg9WVe0pJKDS4AnuS9VF1BXpz/UilnbZ7yZOLNx56J5LxbeW
HQMY9KeaJkjHLlO3/+HeWhD8G91jjkXrSKY92yYs0EvhVaKNFLucsb1Ypj1DLVkX
5y2nHfyrzA5mtjXPeKFmN/63sGTuTGBvleIOf0e3wqFYG2XFQVKiclIneVWXbIhT
5SBFMa/aDCcT3NNGecssDbmxAE6YnUAMb5ugsx3EW32h2lN0iX01x/IwMkdnEZtU
0jI5m5xBHOX0wBHxJN/38JKePAYagrj91L/tWJIqngDpyYDIs82y7aRuzimGdZ8I
rkIlOFtpgMyGmtkfF2M6iJLiVDcAhlo5E2FPKwtIczDpDG4lEIi4BULaM7d+lHxG
/RVbK8XRdmCUy4i5iWaEuEAnw0/qmrCM60mrCiZIqgtbe1O30pveRlmApDtr2XsF
xfHB+lm58VTUiUap6xzmJzAEwIEYKR4m2g/AmGfsho5d5UpHRrYfCddEcYAaOKSO
nt2u312ji8gjcnHchlFpVaOGJqPe/psMS+2ukwIr4DFbnncL7RHaUfi9hN1FO5Il
eRPL9QlG3Yh8sSrWnLa6sE4GQ8PrwAcYZN5n0DMLooNz87acom2Uwjqi2KV2wSbT
c0Xw+rxCsLpvLVjx1TQ9MgPWg7YQrMpa7fl3aZNbmcCyH3UtP4/826jMm1am0doj
qO/VS+O/VdsbISkXvICaTtxLwtRITEPY8c7jgMW3S9vqal6vJCuZcEaVDxyvol0s
kRUCVR561KShpOHYI34juJaeEYqkqPJ0CV9N2kQiIwcInclOcajDA+iaCBTcWBX2
INylgR8bY0Ucy09wrno+W6jz7uHqTOb1rMZO5odK4/vH/NujjazvsMfoqe0yEMrf
72f7Cppyn5DN2L15NpPjLkbadMFqBBE9hARfWbDFz6cCj+QgVC7PIA5O1Td2NHr1
2oorZWNjj3oRiqLBWoATw/mLpWKobKpTEltCMDZjVHVTbOWseL4Dwj9BYQWCJRlj
fk9Iz1VwCTIz26O1gcIZ80sDapQbHMib2GV4oYeuFDg7zvM9pUM2bO7BVtmqmSoh
baTAdjSMtBUYsqOCBXPZHI8u+yllPRaC8crvGYpvyh14G3m12PwGC5xXUIAFMDw7
24Nqej1gZiJWpdQsu0+ckOcTVcHLUEgjvAXpisg2SDzLW1hGGK+FWG6u82jsLRcQ
c494OGpRIdwaByG6cLis2sAYIDwdT5fuVklF6wYxnQbgOFIVkDxf1k0MqMeDPstq
6P5NdCQHWNSWingwKnN7zv7Nzb0wnm8mLvmDd+LC1z50QRo/NrufsyBTIOi8Fl4J
GoBraWYY02e3v5MwqUtYjaUcN2W92uihGBgGSz7rK02Bt4MDqMx2ZeRWmoHa+uVL
0+V/dnCpkeM4hYS6J1aF59Rid+ly6PH0AH7p/aXVZKbXoQwv2ae8m70cTbWG8wMu
dCWPc4UGcdAM3guBecXL0xTQuwdAo+fMRpxrffT5TC9brHRx1tGmqUb957ZFIwmN
oVdUwxQIswwgIMWgxh/T09JmXj+gh/q3AdZ0hJ1nPNmqs94V3OPzcRwNB4W8j2au
FUzXV2fF8ImRshUNXlHRw+ViQKweciglh/LybxDdDymwD9OYMvVR7Z1cKZ+626uD
cO+5oPQ2uzBLAMX29UOVUfy8YKNiwR6YGG2su9EljKTQxMtptNpAA38so/QP1CGl
SY+oRCZeO55uDRcHajyBCdYlmnUZbZ+uhdzM2U2eFKCsPNHTBmgYPltzo1SiFvt7
BfXwbCNqdxW9R9zAXMVFN4+biiKUvNxWExJ9tvOOSJzPDPT36Joxa98hb++LEYD5
gIX2MJzYVCW0lKO19INbiA4MvBUsNcsSb8WsWEmSEmwvETq0hUxSulWEj4Jw+ZLA
FQqPGuudzumpYJTHFCgJax0LlI2ZSwqGuSGWTXavwL9/FUx9p/09zuHx+EZZPYN7
/Yh1U6fr4rQSuJbRikZfEDCiM3TsR6HC6flD6clpBhtpGTMkrR9sk7p6J0tH9aaT
aSMUaZ1WUl+kLnRkGPiYHlg3WAFG54++w6wuA3cf7UmRbgwCRVLQjMk2rdaC4kBk
qOuGzjzhHi/ujc2rJ+vO/7af8FP++FbI52xHqvDhmRUPkYKg+ewnld2aissEQViR
/1LhqnzXkj27L94z2QOz/bnYivTqP2GwVb6APPkj55xkQ+T431ccL/ifbNKNnHcw
B2a0nSB/7mMfptxCGEZ2b9hsXgwgN/0wgOF7AAMYW8Y3VCtZvwbR3Ee3+KhKn5i1
rJPsC5l8xe5YtPvhRDpxT2BCcTI4Glf6cqD+wzwSjV9ZN3fqsN7/EevQNNm1wggG
s2lmZykfKsZrzQuL9e7VbH7EUOoSFBNboyZSZcRYbL/mTCwXoO5S0LKN7aMsWnSI
6Q8QR07x6FWS9EkGxgHOFLxZ1wUEEzC0lo+q8HQQLY+7r9KkW03l2a3RzOlGnL1T
NUtbFROURGSCOroUIlm852ZaBluHGxKHkBVyHZ/anKsjU/Vk/PpStUmbTcPEKRx1
hDxDwIwi+P4Mj+ejHYcb0tSnr9cU1LHqSYLecmEKREAYrSXtO2tGrgdI5K0VQy0P
9tqK4IhiJzbSuJd9RV3/LHrpUWfecLrVIoSNblHyuh6ofj4ialsImPc0cUgAchPg
cciNgMKzHyFOXQIqNERNgLgH/to1Z1P02/PQjr/hl7EMSnW5tNHJLnt/O0HqqrL3
6DCLfKJCga/k+q4cdaKBE3b+8qkCzU0rCikw4NV83dMRyfS9HmE9QGWLFbdtmlCV
lPAlM0IkvV3Iq+c7qYC7lDjvDSnLgLTc+vA3E+Z6L6IFdD/+C+90FQ6s7X/desIa
KRWErepjRu+TBV82FGXlRdCh4IEMkwvpZEGVqtMwLSBNG3y4zDITexEcAVA3roDt
IpmEUICSrE9L3ukjYJM3N7F7mJIEOTq1Aev88FUtCvxRNsTFfpUM93Xmzzd4rOs0
IkerjicUj/yTzatOWodYBRSwbih7CfdgFG8em87/ugu1IwfwPKUDKuoHoD3VTvAN
38KzQdOyV6XHDwiWA66lvRcpSyd/xE0veJ/cgN+dp4vt2bknNolnOpscMku1NX5z
n58YEVDstqvwDhATLr7MdWNPnfA/wv+JbveB/jT0etnV/kpaYGLJK485oco8BC2I
l64rImjTOMkwxsELTEY5bpuJRhB71p/fZlWL3PAw2V0YHX4rfHcjp8vYIIoPYQ8J
+4T7Wpr5e1E9mWCf5FeDgStGxt4XmoTF/wkEo6vlr00yvzrSMNrDGGk+m1n7s5kk
yxAAJpsljXZ51bpKckiX/3C16/JsSehjnUwFf3AhDjhactbFm8niJiCBEUKZz+jT
g3eAYOvFcx5Cz63niIrkmFwJ0sABUbSyz/mogktGuv6k/zw07grrKkAkZrPdql4b
kBFfleSFaf3J68U1q6aoXGytWXMKuqje4JyAGnbYZR/2rOiK613if8Qhe9OBkVlr
4bP2GuK6I0P1mlLVOTq1PAT677I0BUMI/GbuFRjiyz0gcjZ5Op+N+XhoTEz95aFm
89SJYISz6he6BcnEGMSH0XMZy5IM9LOVU7F+Fnl2KjUdSu69t9O7Ro0cEpvhEGvC
z9PkwGaaw9N0lOdnJQ7kjJ8o9hnj4q+/MJLs5zvApySO9sQajdhWApu4rDugadfD
r1RSLcO/9u79XV2JhmCH261v3n39AeCGf81GoXHtjDKcMFESRYQgs4Ni+8Dzclr4
456BhB4tAJz2o24uu3rVTB5BKEofejA2WE/r2KgldIKqvOgvHmKpOgyAx9ukcFDA
4nlnIzQpypuaw1MayJn7NSsR67XZScNSBxsZ6975JdZbQIqP2SoNiwHDJeVaxstV
XoMhJgUeKG5TjdKIkBo6aQq1Zl4GbDSNmiwhtOhTpF9ZT+1cjMEPDDRAO8WzMMFq
6kykeNtK5nNbTEb4Tg8e94zSxui7rpThj2OJwDr49+UbrA0sqsJcj9WKZpEnOpCj
QYR9bCgzhUtUBMbRmRE0I9kR5cZ+hzNHCvmlSyauQgTSdB74D9e1BVh9asUGru7C
Wh8h8dfhlHctN2ZbsnyJGVZY+nU41kdf/P+34IP5V7T8HT50mX+Ek0Kcet1yYTjw
FThQOOalmchh/nj2IzBe9rf2z5PZ0kaLr656eP5wvciQvhkw2aeyl8GMDSI7zrFa
/+M6aYcMvyot8krgLljZB7Jx9Ojy95xCbht8pgmyps/qHfeSaejpqXzRLZQB+O+1
6UVT66z3eo8RL/WbokcJe0f/r5DCT11YJfbwYvqILrk0wWAYiGK1k8icO18lgUnv
DKOBYHn4Z8Y1u6NFgi/2eWuq1ekgt4DGHE3zH5O/6WD3iVEdViCzOLHPCTM4dWTx
xk/A8Znp99qz2oI6g07v1JfpUNDrMQ6srnrMqlWav4EFlrvtLLlwMKjcYAt5m5NH
L2gVMPyemrc03UQFkrSDGa2cky2tflghXR/9c7/6H/BD5wFXvHTCZxSashPmDTn+
ROZ0lR3u6r6BMaKFCCbe4QfDEqGOSFS1BYwFf/pNxzwehh1pSqsLvrsCiulNJ+kZ
CGvx+xcpfpAEVnyOkovYzYZ/L3zpS1lWFXpewNbtJX1sU5lGfo/5y9oktT9VhsZx
MbUal1UjqKyqup6KxfsWGq5eyvShZf71HTYkRFsUQaXFSKltosRC+nQUqojDBtLm
cHVzSeinbEyN8SrfXpLF/JTGePJA/EJZRZDOoVY3v8w8GpQfoDmsljjy6oxgUEi0
CSuYIo4oNgSKi4Vi1FN7x9MQ1ctLm1WVVAmVoOx8rgWTVAgw4M1y/qBv/73GoUiQ
TWSpIceZ280MZa/vvrFycxvBKNJwhT2aclE1Wr3bdMt7NET0kwMxgZqSVQpJnlZM
n8z8jiBOtRt4j8SdlA3x7Z9B51efZx/t6BW5f39RL87pqfk7ceV+K/6PDffA+S+o
it7EkBxcGRe7EzsbRWPKwEL/qr0/P5j5ShmDUEoH5moDD9OGhuWZ6gbtadlAr/fH
C7ch/mD9UUrRnkIu/fFnZEVePLB1jLp0Oi1iJfBNWaURH4pg5kAryIUlsgWYSa1L
PVBLhjg8GxdXjRSZIfKrs3GZoZeSmuUmKxP8YG51+MJMRpKBq34l8vWJeRWWKbGY
7BGmoTwBVa/CXbKU/ettDfGJYS7WEZVPGn4TVIfJzWRfNybotxEMQkA3HTUHvwL9
0M0P3i+wWXkXt7pm7Bs4IjcJVOTuYILJTHjW/PJXutoOoilWeH64/d9TYvKIdUAF
lZ5rxSqhfgMjxOm7xYx8b86lkgx51u8XYpq1Gy3OyXq6sYME4mFdUzVQRgrPYMGN
LJa7rRVsMTcNL2isnqGh0JN6jYlAPOL1qnjwqlLcldIwLb5AMc7wMzHtBwcqIydR
CTUZV0s9SjoaDXT4c7+woRcO5gzB6VNIX2FSSuHUYKJpiEbmUJX+kI7Pg4WSFttl
J+K39tOrKVAwATYngxlipNi7tCQQy0bOQ2R7nZBF1VtfPCSEhLJFS/xry17r5Oim
8n90HV0CjIS8LLUIbs291BGYA8YiZ2zRrobuuhgn9MQx534oXlGDDGlG4Fmgxb/t
EqhB1X484WeNOH1PTSmjYMdx9NgrdfvlUzIceAcEAU9+cbgIUAszNnGgWEvKHDZi
6nHXbqgvPnW6uU5XVPk1c5OHLoxMCo6adMa+ttvKjYQsW6Tmums+e2eV1TgKYGhn
Lx+ccEgTB1ehAf2wCW/bzTUQKbu8QDcG5QQdwklqf9jmV34/WgkVdWj3kCX5V4yu
fkazc60BFjNCH3NmJ4GU/t55dP03Q9FYHiCtZDlW64unFFOvU0NDYhsqWOX9qb74
Qop8qGOR85BrCPBOnesgq5x5g8OmveKwVR6+/0zIkxQ59xZNAUftqkdoUP8cHpfC
5ELHW9wvgEYtf4IRLeHhn1vIMPsGRV5kU7C3ULDOOqsF2tGd74VwnFHU9JNOK0Nm
rozia0R4KtA9nUyLAzWw4AhqKUh83W6vRJpwcstRul3EuaFAxuFJ+yYEyXmR+vtm
tKwZf1PL1hRPXDmKP4ygFAWXQtk55Qr47BD/ckdpz9R0sBO5jzMK3d1sbhdh2UxE
wMVGp3qE8y9u8Tk2QPOwSv3TTxYdKQO7drxkTSwyIFM9OTtgQWanfvV4ayoBuPOV
EVs54koZWi1uLbfaWZRuDQV23VHR2qe3siNug93A8gZU13aFNGGhzYjPKxYaBsbZ
OdcCvWOJrGUvYzCd4oBK/QO1zezwcl3+d0WkbBnVUwfHKR1/YqZ23dBt/GvfIv4G
v9JHXRTHUy6sWM2Gsh255d309OzFJcbJ859YmC7ly9Xmo0uJazJ2pMXjFced04Ab
54ryOMyBgOTMjaNeNUZdpecy3zzeE6ARwuuRkySKk+7cdxQAgXS66hJlrFHvG+HJ
xBkQZLYP0vV3Kd62+ZSLWEd3SBLm9Iwu42+9g+knJXWlj4/sr6idtdxuNEYTL4f/
ZNg2QS8i6e3lKvkvDWxYkL4ofHpKwu03wUjESRJUTTBYqNz9gkVX/bAEkg9eqzkM
0HRbsyXm6QSzlf1PyIGOpR2Sf9TSzwy96gjsZRe1ksdjDNC0c3F6yQxWT8hqUhs+
YteKCo5OJB9Mzc3/PrlLw7ly6lgCAT3B9kQcJYe8tLzJiHkmqhyHPOYcB82LHByi
9c/iuDsSrr05oTQct1D6vBsnOSwkTjSwplFtHR6Q6bYyGR8mVv9vt0RiTFnqBtA4
TeugPQ6tVBLNN2aT+wWEkiNgFoyahgMUiNtPcfx92pVdI5jlDDfsC6IttrSiEAj+
WmCZXMjKPjTsZ7tKq9SKKLBv/B8gPIWbLYzne86F1WMxudQtJleUyQZlEqFMeqns
ECPbsUhXRX7iasW5k5iEuEMd8am1qoB1lvqbUf+PipY+L68GeRaBUPXs82tIPd4D
DMrRLBaUyN4+e1VU2lhcQvyHx+QbSo91pFIIGUqepwtgq07t4gDDplALY+HH4lOO
9C7ynC//2ydyede66yIl1QPE/oVHipk+DVnF7Pe33zy5tNnIShMZBUT/2+pgz7vO
JvYTyZnIHFeb9lMSSam/cY2GES6DnTa1Wh/tLigGLr7NtntWlh0RHLW8ONP9dbc1
oqtp8PxeFvPtIm9hhDkEqyOT5vLukRwke3G8+slA0xGXOFhyUXu6cMWg4UUlSGIC
6LLxNXVLRN+ZqvPQDPV2/4+P1QWFVKspJeNQvfQtr8iGXkQwqrL5SjMjBpSHmGbR
+tbrfsM4v0ELyzjjMP9LSNBjYqL0QQIvN1zzGlo5BekFeAzAJOEubJ9mWdZzXoL4
o2miP020myChKrQG04m8c5+o6I8FwTD2WWc22m4DUlMnlca/BYof9ROYo8Pr5qAJ
gHTDvT31yiwWfAH4B3JUFUsFhn+II+l/fzwH119kP4S6GpBFvcBKMXSi5WVRhWVs
KW4XUcy/NKQyrEu9KU99TAMqH86dH9rb7x/N3V0hjzcNKyG4YpX3eeLkkYEX8pgB
BRDHt6EH+qqAo0LcbyyG5KRfzXi6Vx9YYmdF7i2moAy8PzN88hu8pfzgFC0pB8FB
+GcrkEDYCzwG0TjnJSKYH7rqFTCkXZr7w2A19BFLacnnRT38g/CRTi3SDrScNJtR
kGyNPqTKN72RQmOif1HWofbKS5DyYgqu6b0yJNcOXFrpnT1Wlgisj6eHPuIgO4iE
OziwHxrUkWISSE/H4HkfnzdA85FcufhqK30x7Dcjj9itW3daFInz49mvjYWsO4AZ
PmT4Y2gNPbkR2xpD73tDDwr9z+rE0sPUNdHnX1VnDeVbcD4GalgF9K/Oj2/X3kzi
1AUXhX/aBopndIWBe1M0S0eQR0BqVDawZDyCugD5dcNsuTT6uEUtAyPH+9OdRSM6
UySGfxzMaXvJgRBI9Sh2GDvBA29pkrDT0KCSrSxAwHtUYjAirn74vvxri7EiwdUq
9WN6xhzkzXjFF4kYESjxVIVNv1o7FD2zFT4HO6vUUeHN7eckZn2zEr+elC6wF6Cg
sHqb9k0ZnqQAmr9VpV4phoHVj+TFeJ7H/T/K8Ip3F9Qv05sJXkVZSs58aWrSRE3w
kePrLxDOZxM9vrugfH2P8NNf+QB83Yaqf8h+jYF524BVbUhqbz/vTE4jt+m+f6lh
9M98P2GKtoBISlO8DNYyCNN+Oz6xSk9NBMVbbQW8EnylRFRB43Svh4Hq442wvr1C
EYoBXLn0/eGEG2Y9Rq6cYZ5kvNfMynTuWeANrBD425529PEroMKsrXf1KBcmGPaK
6Nn6IuJ/pVpdy81wksdqkhuWrCKpUqXBXmn8B6hXQbNfItMecwF4AcYmxpjPEUIr
wVLbSJ16b+TFhQ1xiquBAj7Lugy1WWRMqvX6iQIBryWTxUiWw81v1xmhKGkcOV/f
2h7Z0EDdaxRkHOFvUJSMGMKia5jpFD9TqQShWzNhOP2YJNUxRIIKOEmOZlZTaQVZ
uD70eX7gHD2U9z2pBL3LNTQbYVi5PsUS53deS0SBhe056CeWqMz9GP8ebM5oIB99
KjTTRNFeqDjnV+PWrjUmLI0tBTqInbjAAlKO1QC6qXund0nIu5nBhYI50bQ7sAC4
oFbNpcPFZTyiiomix8/ypMp1P83BE7NDYYkS28FwjF6458UDiThwjr7gg04Nbk0T
pjVXSRV4dS8wkG+m8RpZOVaN9R9YgWN27wll3FDFHjcO7FBj8A1x9XK0cBiJYAjm
5PJkHtH0g2bry+xnAzSXZ7gGoxa1RVwLZ5Gp3Rhjh623wgmWMMSFfL9OIg0NMgr6
WJ9n2fOtk8b+h75l6DkUbFG/Lr3Fi9Ni8tzpWEQuQpGWltlRDb184fjqjaifkPUO
eSh1IupWvx8KmqulvZndJF3ppvSwIqPDePKv+59C6EwkWQuot/YQrVaxsZyV6tjZ
RCXIEFkK2A9eK5wue4eJUI3o18NMo0PoAKM5NcudWaIPWpwh8YWCPbHMro8fSEsq
U32MIJzkNyr5MMkSpxygK/1Ay0Ixa0hY6046cixTE25gzeyZmYvS1oiOYZX9lAbf
SJCJWqISU1kVfbcCMtu9gtGdqnpufV8k29aAIQjTQ00gQgXjpUERW4KHVP5KfI+V
CbmHfflUUZ1zqDMoIKuobgvAlwYXiW9vKZ726MttD3uTe6iGGwRXByljUowdIPfS
8aoJSUQ5n07Vi1jVVnIUSSkwbxWdxrZZRPEEDV/02xkGrp2j5fURfxpZ94xapEjc
+2OEblpms649dHohZaQs6cvBzxc73ckiAdrdkF7UnVIGI1q+VGBoBGsLqieRDMD7
yDPDCxJrkayQ2inODB6QNqvrLZ7pyZh3FNNCPyj154kBViXinq+Bjt/6aMO1ibkE
9v8kn631JfnhU+qFRx05D+SQSSLYVBqC+rqgiAssHMycVXh+AcMURwi1O6XmXw/W
KLK0XpsW2R5L7oA7DlSyxQYlDXFnbw9keMMbvRJIg8P42V5khER84E21NJAgYg84
Hz5LCv05gnU18ysDNuN09y/zTCJzjUbWUNlpPwkIPnsUvx4o+8apgPQ/1QDJkjBj
nqpx8bjpO7Uhptbc+/OpD5pV4g4I9NxHolXxvS5are7KGb6duolbYw5RwVDSBUqp
qytnObovtEQuPwGcloUemGYkdHYfXx/YTQVIeK9dfBRe5Aav5Cthq1QhzrHTU8yN
XSfueVswDd/yJneayC9SyydMszgLHC1Ee3NpKJq5VWvEhC9J4jo4e6kzmwPM01rM
B/xMqm//tpcyn/CoLFxSuIAJQ1zpiNmLJLChaU+cG71OjFMYoDWaJBrpXrJPbVbB
yzSyYtJyrnnqXB39LfMUV4tGUDnJS0rieDl6+2zCqwLOQN4k0Jy0TuhK30neMYKJ
kbkTDWsIbtgAnR2rNduIkHwKTAoF0hikw4DETLagqDkomQoMBm1jdPNKC2AjMTt2
7M7cJV6hCRDVAtitfhdoABJ9LdN2PoGLscDH2fUTjaBQL4JC244iB5FsQq7MEMx7
wtpRiF09EJC4rMy8+EmqQ3J2K53SLYFwftcUH1E6jPBBs/NdJeocdNGOUuM5g4kW
HOOv+lMWjIMupayfogAypXX4uM+mQnpyJVhAjobJ8R2lChHN4Dulyk2cDi1Ko76J
ueCRa54BYybPTCndT8hsRWNLS8z2p5KsC2T7eeNlzmC3ngqD+v5dUE6CXRXFF9/a
oXJlaBmpw/qLW+ER2BlKop5BZwls2kM1yfFj2s6H8Y5ldqBgYukw3jYEqz3+KhB5
98c9c9ePttOaz7OcV76c64X2YLfyRJa5+DCUgRAg0lYIxYkeFCmWHXQ/UEEIJfdW
YIZ82QTwi+7I2MZ2w59aY78PBwCdZve3Rbi/rmbzhKzi/5gQXV4n+yyMH2Zcw8iM
d+2efaE0Vt3LQ74ZTezSZrrsrxoICEbuJIt7fp4qD+cFD4hPm/A7Cs7pg+XHogYO
vURqyIB8W5omH48g1dkAY70LwS/YjoYBkcjMO+Vjcw2Zw6i6Yccq9mpqXOBel8QF
oBnGzeRnNvQhlce+we4kj/zBpdZf9p1BCzwZq/Fv+DVN2DdO+jqXqbH6stWP01qd
9jcrfqJ7eVl8SP5+w0u8vpEzLTENT4L9FxJWd5ZwNR1Ap32uO8KXyFwwpuU5F4AL
xWPZzhwcsrFpzHuyZ0bhyIzmrOHzsBboMMxAGLuw11xqgysF4gFDxKHPYqsAHCB7
6Q2izULUroUocEkTcsR5Onzj2E7qfZYwb9G3nYqJM6LYAHX1HJzp4qiRzpE8RUSM
Qb/IBXOaMXRQC8+9G9qcFV90eizoaUEcgiavPwhTmbUYYiVCIU0gHLBxHd5RzMGt
J7twMjES+l9hlYGUsH5eF5+6tzccXTPKsKw+w0XB8cn0+x5E+BI4ikawvsR6KfbB
et8whlu1WZK359cWlzZ8GxdGw3AmjGknvHLF6g4Z0Z/O/JQiK43QSRZgZWIASYNT
WBHc8kPdqGB5aoEPRViDSYcjjziL/MpjNuyJ854GpzP4XZnX0vXFhrjl1FpV5VgB
olRbayakFfCpl4gTnLI176hB/Jv++6ig28gDMSd5aW788Uv/2KkUpphz3TYNy9HJ
PIkMe4Vv/iBSLH1sk0LXyrPao85RZjh8hcVYPwyy+3AXjnI/QucF5oNTvMJrKOPD
azzpB6prOyU5k56WQXFuRSWkGpXfT9LyVr6Tisr460ozcGIPFZrBilfg4ON6J30u
DHIoOM8cb+mc2GjTbmlVv5SWRAYc0Cc2d9DwTXfOspCbd1MEZHI5JyNnQlBFOrhd
vG0vDLLhykz02EZEzCbiH1QUzK4Wkjwhb2GGAJ1mRJtTYTglm0bHgyuppTakAMv+
6D8QlfdsC1wlOEawVySZ2It4Y4tGbLTQ/FwfcrS1Qs+7oxL+ZMYkMvyrdG7f583d
0TYfvIH7CTyGqEfZYnYIFutV+Zneb8dN6EZp9uGQdVaYTYlG/gpevxNG2xcWlYd0
xyy5FlXQ/Q6V2m35OEPLXBfdKvcdd3fxdyXh/Oa9apUuf2TjdbHABrcPtAf8NJon
zT8X+CkrEnK8Ccn1viWtUaZvinCBwGjNbM/o3lRTlkCFMHyJIfnwnIVU40zHkB6y
Uxc98WBlY0AlwrgEV/cGdjzSGWDNYPWpcBrOTnMs9BxrtWmc2b4i0LrGaKtE3zt8
C1RZQGWzqf92nLKDiCXUIT/wVIkVG4C2I8dx8s9nWfUM5IOuFtyfpP8zy+21joVb
WF4pImI/CcJRKStRY6glPOsOSFLUzVpDDFOiGVC4mjGXuCuHRWboDmAflqjE9Wv/
/TSVmHi8wG3uq++8Tv/VGmwhbgTc0ynYKWueN74gn+CdgyUwkZPzJl7b57YzO3BD
YO5tkcJ2MDkYUPjPWQVJ960+ubrTZmLzmdYCD10ElZ36twKPwrAvyqSW/Cvhg4jX
A0LoLPQfoumNVy30FW7hYauEhC+QplQ3Vtbq6XL66OAu37WfgopvnoIvNr6hKRUc
L491xvfyIL680uBBk449wM18rz7zA3LMG6ywML19wzDSCWqfsk88qV7zJ9wLoh2b
nWmHlWCbBea+lyC+zRo2Ikf9871+70M0ZHyAFWirWp8LHcGA8bMwiXCqa2auE9f9
McKU8X6R+zhUkho00WDt3zy4viuHuoOyjtDjYrN5/5LPoJKdLdTqKh+NQl0x/Y42
JRZFj3PnmkOaJdeWAaF+bMRC3FqYWvnyKkghM80Ie436BXm/19VAY8YsPZ/zuPQw
/dmAndirhmtpV/yNyaZ61uDHbGBP9Uf3Ngr69S8t3dqTTXVLoiY8KS3KfAW/fWRW
Y2beeQCTU9IIBUcPa03sfHV4mLOQjHYfxjzKdxHEqZqWEQt/OV/N8m1ZqndrnDNc
95y8J6t5OC7vfetvOqjl/AQFAHYdAi+hmJZyGWtvLPGvqHWPQz6nX7GlwEqZs65k
dtiraWGsefLu5gCQY3iSvATQ5bfcUiMfbrVwiE61kujFGhrmRwENM/5KMC95v/Iy
m8h8LtHyQBp38swHPL0tq7C7ykNqGty+P8sSkvNdf4W06KW0ZzJ5vLxIynOD0R2q
1CdIbYOjQGhdRs9+qo9mmufN2t5jrgnSwrtK0gskE4StroGqbEIjmQobZRfg8k3x
6RVyOTpTOwzIVoFc1keNmgef62w96zb3ueQ4+7v82tSLPtWQoZU34giPjZ9qF4bM
a4B1+N3AQ650CijDwO2Sub3tsN30OLMx0UeBdmqu9gsSkFG29qKzFa+YYuhbXmB6
f2emTXJkzVfTFyMgGckeC1d+LhEWI4js9vV2ndEvABmkmWGrHVLWQNcb0+0YbB6d
3zv/Mt/Sc4nBjORJ1n+CVtFwL9YFDdhz4HOA1qoyDr8sx/fNjo08sOjr4q2sMXvy
+g6XKXTdGpxmIC/FYcNjMuRbgxvg5sRTdVzU5xwBu9kdlqeT8Y1W3SrxThTUPOyb
kIeOgEElAndEdnpVGqdlMjxNx29Li0Tr4Sr+2HtJ8/T4ZZjNWfJGgUS7Uw7zMwfa
i069byzpVLXls8RHdrnFt+8c5kN62QQ0kEmWsnOS+dzoxcZnQk09yNaGxY7iW9Wv
SLrqAIuYFqOTiksDh6OYEVtpBec9+iN/wzlIL1zg7n9vOO7G9usrJmViRv9/C6+a
hFCUiXYdQmZwx4XPYmsTpil3f0sCjjGnVfuLS/1RJQJRxRodYhmWWXQ2sOkUDDLk
/9TEbxpJfI+7lNYcSXZWzANvJK8iAYWIkL4QPKA7dZyrt42cp5yk+j6qL44WPdrY
DtNbOwj0totMlunhMolVu5fH3ZBFZ2aX57U2LBucymyJ/gu4ATb/2ULJsylV4f6S
jwO5AyERKlv043/D4UlIf7e9ZcQbs4+3m3CBHOkiJDzAJfbF1DPf9CtcAhOsxVuC
TqCElZdoA9+AfM9MX5l0c2AoQZeF1WpMAWUZaQmH4M27CDxHuEozP4a9hpvkIjU1
I+/XO5aUMTqByAWbMoqgMpG9wL04d4wbz6706yDK9/RQzqmEfYkq/AgIiYKAs4y+
ucctAZ1Rb2pH1Mw/RXUvywCnqcLb6HrYtQHLwHSLK1xqMUWIejHH6/s2ZVQZUAgw
JS6l6u5bMZ4kukReDIAcyuFjUcug5lB42TCKp5i2cDESYOSGCmm7vViZUnU9Uj1u
wm/cKerlQojpld0YNSAbLsxe8jmxa6/t6VUsrqsp5tMhzF4eew4foxhNVKtGOM5o
de4VUukqMTew8po/m5aEeKxbNAChIpjYP7LcKqemrRR/c2d48X0D7Px5GBfRsfpf
/GXQizf1i07Rpxk5chy4/OrydoayeWdkF7znHgtvgnpRS5+CPrqMWO18JQBw5ecv
BwSc9tPe3tiYYY511+B7RWYVq/cPHYOdVqzuY2SeKwQI4fil1nzXYhssICd7B6tb
698iYTZNJEzy6t8M2pqJgZywswJ88BmK6o5V0ta+ZTbySE6/F9kVui56Xo4+oUce
K3/fekcf5tAP9XWBTK74FFX8ieZou0Veod+1hZCWrr9FsjfNMxOBlPhMqpo3GhOq
MOlRAjRJfgzUlMlyYMYELjvzeK/EpW16hisvj6Uwv1cdzRNd2WU84CliARe/2tTl
TOpeSxaiuB87wIljseogE9/oZdWm1gFZbq9tw+hx6pOlcmQjzypI6vmtcmk1X8Zo
6ECxy2J3VBCfs9hU3VYPGHdNMbvcgCh45Vv1wXAt2HsOFfHSFHUbkDfi9Px+AjzB
hZae5VBZk1oXnQfY/42bKb2G98BJQmuaiNdxBJR+jyn9do1g8nFx5eOUYeoqUVGh
yj8a04b+WcoeRH+V2VodEJh1h406MQ3cPnrSTDx+RhWbSOxZhPNUjb2G3dS6+bCT
rtd3Bly9WuTJbha0DI2fmAkRE10/Bt1NXNb22mj9/98gpKuwYyXOA8qIXlBV02n6
mb3f+/Ynup9EgJwg081rh2DO3b7ks8dIfLFEkyDKv5fj6gzaXD4/2P13V0TlckLK
uWgKLeMs6O0j5VfwyA0NrNO4zc/eTpFqNjpMEiw5DDGiOJNTpOto6SVq7trfdtJX
cWZHanLgvFZ0aQ8UhIWM+p2eN+rk8ThDmZSykVReSFfVAEh9m1c9T3ftDvC2fiM5
Ot/sZ2nhblyxjR+Kd0dPQp6V6GqbzN4qALkfJAAZ4QYHeKLXp8ZisQJxy4rATgw0
iNNbDrHjrUwJ+xaVThcQeCyRjZ+3Nz/8n9gU+UEmL85+6sX6/5Y4u4b/swii6VqU
V8zfGvrr4zkolk9f1xPn0fF7GiM9+JlWsX4KfIlF2LsSNQaeHHemahmyRUHWXW5p
yuyuFEKjDIztBTeKiRK2pbjyLRyUe3EX1R/pQwPH6caJKz7MZL6n00SMc0P5YvLi
9Vt1uUuwCRQbrLVYdoCcmjYZ4VM0laQi1cDy14zeM6Ea97LKPYz90iGGROISpHM8
r2liVomghVjmh746N46AFNg8pHBN72Xtk1/8TBQFoJprv/Tbv/Y6eZjB2ZPNbOea
Fh6yqr672qAKUZ7MtR3ygETUJ4rwejC9ZUd+u0o4RS1bid6tCkZhGxeScmPxndll
yWR0sc//kxMY8Dr/g/ejWisDSOUjmugQneH3iNARvmVsb8WU806caygFq1Y7g9Zx
pgveMQHXSQd4g9/3yMJnFIPczyxphp9NUYqtWW8OCC9rNC519RBNt2QbrAvjeCHh
1yyunhBcgx0iuzM4CEzafovNkPnCacbm1lAViVxWs/eH6+FPlzavjOsCgTtAW8+4
4PI8B4nZsINFMTW1RuYgofFo3d9SDXrzLHm/I7Fwm8GoMi3exfPLVRNirKBAVg4O
G79DJKYY63Iv3BUesIpwoOO9hmkRwoXXTZHsyOm4WcsteOhs4EnKL3a8186Jnz/A
A4LtSQi7CyNG000ye6s8yjaOyU9mPxATlinxBKTyyt2GZf00lBkNlbh73Q65M95i
KiYsksUx98Is6SyLCP0nsAWQ5/JlaIBAFt8abl61cskVG/+E4Xng2Xz+2KL4VkJW
6A8EPX3VoHwdbGoY0sIKiF/ZqlGlwBt3NX+sGVWAq7nsz3YgU8jCiNdk5s5Gr1op
mPraD/dV1LIKe9mqORitOg8XuSktwesUWUxEG947YppBljUroAgs3UJ7R2CBxB+K
RY6O6iU4C86HTVRrAOdoNG4gIYmYx1H2wH1zpiULv7XIm5k61SC5wrh8jjnSh/6L
fd8CHx/RqsUfLbT1m/PyhQ9cKdbcL986O1wH04bt/DGNIcq8n7koyi45J+F9geNt
PhQIESK3wrr3e8YUyKpjDtUt3wi+gCryumu/vLxAzdw7xSzgDLaSTcx6+xq0/6jf
EvPEWnB1SegfXdGRBZs9N7D49J9dyf7iN9TFR2KFyptv03Y8AcK40nKglNPQZsb5
Q3NLAm7qb4dDgQMHMksc6gFSTChQBr6wIo3+PhGOB0LnNZ9J5u4VPFjYiM1UXYGy
QeYlG6vHfaZmiDqKtY0X0bAxM+T77C8tYT4RqPYbbBpYgs3BV1N5+c3Fv/QVT9cS
uekYLn8LkbHTFHJh72yRfrK4OtC4b6xPAQjMqhnnjS9k33WTIvNW5UPXaQuU8GYk
TWoyKCRxb9o62sw+AFN3rp2eGhEeU9u07Y4qIuRPY1QM0jAOddmGy52R/tQWdYqY
zY/k7daEvfwjj2PJZ+J7AF6D/MBSDtdFSX5hbuUwIaVX4MOPfca7nbdwAxitccb4
On2STAVTaNO6iqYepD1wefy4QFKa7K0NW7AiN0ug80bJYN8/tU3QoTRHGiU4JDtm
9a3x4/OvZh8/vOwgPMSD1bHuQTowYPisHiV5dr/z5m5RYcbIqEr9DtHkj/9GJr6L
Y8fCc8ky7KtlYnZEplY6UEW9by4nzXSz948sNXktz5VfRuXhw7NFcCS1TVNHdAcX
PW4J7KDET7hZC8SxKm7bn3Jaw+SlikGMsV4lR9RvM0ZjnfAmZNpOWUMtEEXCkIIh
TSpZKklQXsYrbkW1x4oxsYNMuqLKUASqkkayvyQOsDLIdpiC9o/EKHu72PCrkYAb
j5rQZWKn5rcbQLY1ApNm9Q2rIitCPw/fOvfSFF5xuQjh9FY1LU7vlDZPdtcwhsCG
g16AT4XGgy2cwpx9rMrLcd0DQcjHT7gdSKNZjmh51+dmefc6hxsuINTTZXPPSX/o
fZhptemO7uSqqnd0mgkcjcmZsVfkMGjeBoqyVMgwT0/zh9umhhkHA7g3zozkZwu8
eP2LqtZLnwbFXj8fwtKcU3hvxxbBU39iW2R3PSbCYdfxqDUd4tnWWnbakjZD71aw
ToP11Uc6LC+dkHF/G7VGQ5+IwkbNxxqls1+XenaSBTaI72cpENSWHCnY71kPkoIH
xcxl+SRbNKgaiuDA1x+0nz3WpIqXrdBZFAhfqHBUXkOTNX93bpu4AfXv5Rf9XwXc
7VpfpVGx+dcosKoVoP78M/XTP1UUh0G913O4Egea8IBHEyTuFEdaD++h9bdDrlXx
p5d7m305bRXW6JdR1PEzJ75bNyJ5RqeK1tamKMR+WqDzkUT6Mmip0k9xN1igLlzc
3KHzjtXImzJlpDAY0ROTmo6uRJarvvHo229sdJCHh2y2FvUyCcRVK4qhl5Mju9n3
pLl+Hyps7LkyzdEVQ4lLEJUZNQcIslqpMaFS1I90sC4paizojbs571qIEr1w2WYR
H+YuurGg21qfC4WB8aaWVTr1LFXv5Xrdi8fSiCdNjsXVDOnsNqCmCstxt6hkgx3o
vrvie0S5b3DiyHsM0/iuxWFSIUtqYWBVdZdUBPCfjA5NopmW0gzj1EAatgMhIIEN
Ub857GH0ysdY5IxN+9dTucH9KczI0deMbQWNLbrx8ea/UmeqV7urd4JNRkwO1h96
j/wzSgfganrhnkMr+dRzquf7KbJwA0kJw8PvkPM47giL73P7odVHQ+q7DOkqfuD6
MHhSyzfZf6Du8Vs1Aa5kAYiYSK1dDiHANzn80hcgzChjvdC4PbITTFD7HXT3McW+
K7+o5cgMqDgKSkqVtuSP8cdu6SnbcYKN5PPBAFj2riIi+fvtm2bfLqzupl4wbhPY
rN33szf3zei/rRU18PWIrRBEEFfl9cZi9+EH/cwdfPqxMa6Hqk3d+Dres72E4R67
668SMO2RgK72/XvxgxlLuT3lVyqRzgZuwWIuNN3I0RuQveRxAvioGE6SMvbjBVAp
Sozzz2ux/USoT4dLTjAvrd97yl/jgWP887fO7wBuCjpOBPHw1SxUjREcKbPQaHaa
oEF+MZwXpmM+iDb8GA2z4oB8ui+djsLGxi4qswR8VHKrLS5iqx+VMNCcc2MkGl4k
kOJbp9DM20urO1I4eoJsjb5UUUGbAgfDersrW5AEg+RTeSy9U6OPihsS+PmQQpDp
GANy1VDPYA7kiyS6qrJ+NzSJt7FY8SlNDJBehVQdV58e3MUjyUsabnC6Z2tZ5Ynj
AJWBs1eWwC4XneNNYaUAm4xxKjcrMYTM6w/70IAV9UJsTMwJuv1HeKlXHoNLWQAi
ZisU0U/cNvAoS8rKYZZ+EDfXmvrmkfOuIc88VNkw0DJLdr/E9kN2XZNhuML8WfKc
SHTFi06d6fswUayMOxe23DMgAeYlhRUzAXMsQQfN6qgOzVcRSHoZQwYuDtV2PMVq
VXxXmppgcVBWlr4shPK3uS9k7vfBjhDCSKafqsrypErjzcN55Yo1lqnRQ297ESZR
kK8JfU05QLlMH7GhEloOqtsA531xbipFoMTwPY8lYcbwOb9TJ1jGiqjmJNVhp8ad
hUX9lzEc6oDbP/ZxVNrD6n/mnqWXD+qqPgugspJ7xE+BzIE0L/1YZvWRXDM4sIyg
HdlgP2ebxQk9Bsr+zVlShXRdljoMEKFYWa1yCAygQjZkeb5Y+ThgnQDfyQIJTFlT
wxOsJkkuf6qSMSgd/OWh1Wejv01j81cPPILzWHOQBK6GYVumFdGmBX8SnBNAH6FF
lNWywIc7JRfy055/qtKLIeUYknG0BkstyY+eMSFcqTnzIwNGVb/CuV1M45Gu33at
ReNC9veTPN/mI43sZvlR1vp/NkHUkVBeK74m7nHcdoFOmxoiy7Q096EUJi+Vs/VR
YviPOgaObyYoK4PaRrveLMxBDNGwFzqwJk4v9FTkN/ipCp1W5q8G6JagnS4uzIyl
ASKC9Dy3TgxVYCH25rzE3ASV3PHLRSdT2jS0hTVrvVK+ehHywAsrThUUdzPIyi9b
muDp4Q1B6aaXGY8F6OUsOJ0doYoAlcAMmNcIVhe9Unc/Wg9LJP3LWfZNdmt6EImD
8p1MwcUi2RIZ2Au3WHaCT8yDucOf+ySPkb+L/zhFGAInpZw7ebc9xpfOr3pACGqY
ncfg438qD6CUXZQNh7RzMKbE9fqK8JBBdtrxyNrEXwuRL5/cu9+al84kT/w68qLi
Wvum48tVCbmcY0j4b/gkAisR7iikhZ6lwVS/KWvxOHeteMQcuKRTzxBZ0JNRJeSA
Y3WkN/mnIxEewG3IH7WxS0K4WU3NcizDp4aawkI9PItiAeDpZ44nvCu8p7wrNoKL
FDke+Bx1+BvlkIWe0pyyuIKFpMTwK6jdlC2M57oMiiU/qbg/PgEClnylOl8BSTzF
rYgV0mopwj8vhsLbZHJYfibO2QQYc95Y8j7usSXPOqGqA38zWoHduH3xoqMEIFoe
rM1nt9RaaymXqYzkljNnWxdQOvC1cMh/+hWiPdZngjUk2K5x6typwWggGIYOYcVT
NAdljNzgrasgxTp0kPCfa/gHASY6JwSH4Etw38UgLmThqxVscAOklFWdbRx2X3zS
QmCanQAlK7zWuk7VfVIpwFP69kvk9oTLC5MBHSiBHw8Pz2XqCJbbjfxvLTRc9BS3
S4XK/NJ+mtZWZOKgVrHNJ7nEFW6p6BOyU7Nor94YMsiEHwatZ7fpkhi7l3wmIrkz
p74L1v9OTJQuZ127Dpko3G59tG/i0ZVk4NnhZQBI3ldIv+OfwS6YXrH73B3wYRg7
1Vp+IFFjwmoSugh9iFS3ECaFCigRcAbvsOPxdIHL3DV3dmVqkSVP/auhfjjmdQDY
W+5eA5y1KVSwqDn2cUFDod4TMOHdkwSwXvedl51SzCohO3+susOUuHlYWHj6ixfN
gQz0RV3zFZe5KXOYonTMi5Rb//OMi7D/Gba2Nvk02XwYZ2OJOCmFz7I/2u4bimzl
HQ2MoVz/vWb8Vbv1NyA63IN0HgRZGIDkqMH8C7UtqYfU3moqIYcKpxBs8tHCy2ty
OGDNz9HeBj5iaeievdRjrAHv7+px7pnvU6htolML8d9Wvj4ey7HRbrE2W8zWsKLd
x2OpMc98x+VaFkot92KZZH+NdbsGJZWerxUXSS21Fc78h8H7yrnAsbZS+iMURVMD
0upY7WGDAwAhGT4F+iZikuNThkPPcZYUH+HIT4W+ENjbx2knYPVMLRvI5kr94Lz2
78nzZnwavnVVqEdH5PXzJsFPQ2PN7TBpNiKrVCv/3XP6DGg9LDxWmG0X8Y0ZiQsd
SNpFalH6F3pXeXKwbBn7QmeEkierPfCCZBX2DtC6ZLq79s2uggjtow56FwxqABAF
y2AcM9veMi6FFthxUWiTk9UUlJBLET7ApOhrZF8D/DCsqaX/sqYa6aZXA38XGeiM
g+pK5VhfxGDoGUKIS3pcBA6rcSjYU7sKQ0zfS8HtM1FEaWVWQ2O3QogS6yHUTb9x
bztn3gBLkFMkydAep/41Omp096puvfUm7TS+6TgxBUMq02kkXuS4zWeqvmmyEpuO
tmT04zbeYdbvhoZ3XKuA9X0m8A7/uWv0OoDEF3lRcuBaMj1HgVBsJFLhMTXnThGT
Xszx9h++dzsGn/RuzsOqZ/kszdXYpPoZprtp88AuXRsAJuH++bs24d/J7tByByjU
Wo1UrtYkRnk4QdRlHFSv5ypR2V1yzTGIMIMMpAYCVXEbViRmjSxWR6i/f9V6BZwQ
pXdAvFVoa+l1Mw5FIny5d2ygnO5ecm46MgSw20ZOk7L8YFxO9JqcEQdomy+6AMYG
tIirxsI7WlofNNOwEebL4xQeC0SoeXR5QfP26Ic/MEXwTRLZTayg28BSKmx7CgC/
x5DymXTP7vu06ZXj4FYcwL3kAAtWQbiPUHKRVeENhPcR/yYBcGfbF0CxxQa4sZpn
ve5LRBR21t4E3a36BFwk4aSjraNPxZC/BKoLymxSJc+mb022P9QrS/uqmq8OyTNT
oMe49Ezu3mRpd6Lx+unhi8x4H5ATQmxqCe5ulBDfAU01N6NMb3YuRg8NQ/XNRoAg
9UnREEa0MnW97UAcjHiFldUpNTx4knQCVEE6GRmKc19QAuXY93Qbv5udShAsRE/w
k4t/iV+HJrQuxkrvrqZ/BBFsHb6k3qeJmCflel27Djlsu3Ie412Kt/Rnkc19PBuB
IOrOEN3/R8BOEA369jWRhtmeirYx/gPN40HZMoc2f/NFXqn0dMSWKNDe62BoQmET
a+ai4PVDXUh/VlFXzj+dhCzqWnH5rOCdHzqPxksufcwjzhzTfYBhCV1WM8fmm9qq
/3Mycp/e8IFLdBXkrtG7e63SWrR4BfU36nSQukQNKpWn52H1MsYMcAWgvOgUXb29
aqrBhYFs20/638+wRYO9RFbA1BT/YL7bNb0/8OcxrJ4fkpoOem8pLwR8Vcyzjj9g
0WRM/XFNSX0Zn4AJkc3kf2YKwkAPzKKZ6/j5TRAR1jDxCCB5q2MW6dxeiblwn2Sh
tVdT+4ljrCw13POrtA4vygUlHp/VLMXGE9AacWZe7m0VTTJaIikX9JjlRe+GaOaZ
l7uG9jV3ctL2Pnx4nLkt4IOi9xOv/OycDndqgQv03sAq1Pqe/1TsAXmiFUxdoVY9
fwtu0rMWt15fubrhLRfI5xTgyriu52hGITcXvwqx43P/RUS2sv2jh7KPy+zjJjFt
vZiFaHqq9qaR4llg289q6Obe5aAn7XXmiI8L9AxElA3C2YlFIXn61ubCxJNUIgWu
ytoqcwlj6Tk7k6XLkSoiykO+CdbREl7qZ3oS5NFFhA4CSP4GNHxadHXvcR0fs5xD
bqugL+QhBkOaFr+LQ9v3JxW5o04EejxRKIT6gunEY+WH3eoIbM6IHYU+lWnj/ziG
4UItaBttxt/hdz6FKn+M516rvI5xIjtZd0J8dJwqd7EcLlMFMDfh+RKav7JKqXPA
Uey/UJHgCIkSyrRJDv5dbZSWGiGm7meBmnijE5v24JQUCCbZK137nPPTuyquruye
zFeEgFW7W9H8J14auWJU3+7qRC8wJbHzEd34NMjEHw/kmCnH7gY7tjhs/ZMX3ZfF
RT1N88O4szEcu56zN2t8eIHjqMLv8RbiOoPtI1Qk36f7z9C2hjgPQLudxkVxlb9t
evlpQFLEjcqB8iL5Rz6F1X6RoR9ytntJqUQtOvETBgqrEk6JosvpJsxN2biY445J
FYdddEDIojMgyyfV7vDTlM4hrcJ9dQEM+XSzZITWC8v+1Zjx8w7eMNgNk8aa4f/I
CUIIHbY2J57pRryd2p0oUdPsbRyBWsJiBjArAVJODjJ9lq+W66Ju0IDs7dKzl4Oe
m1RMKI0MQiyY7sXOvTsbYv2Rd1YjI08w6plSV0kjDNWMxpkM0jq2Bu1hG93XPVpG
HBM3ETRFXVyLOYGuAZZFuL0NAlRoQz+ELJr1SAjQ+PkFgT2nc/TyVx01a3k9vUps
mBUdQp/dxDqnT6mIKadiniNWpNgAndX4VlVl3WSlWCipbi2wId0tiuVo/TpTQ8uJ
YmTkGh4TCcDhU9tLCQutjl9BMaH0grNbQquKDiVaxURmt+iB57NSyLvH0k1lxvUW
cxxuZ7Hqh4H2BUsd6cGrcMRLc7qMXn+/Ir3wdWFOz6K7MoOLu/KsKP1cncaNNLWh
yTqARg3uz8cDP0odPFsirSZw2gjrJWsachihddSepXRLAlBo1ikvd5mKrhw5rtyu
EOLn5i2MazkLv7YlYecAX/ljLlzsnWgmVi5s3P7OZ2AhLwecaf729WzDmfHd6Xcm
ex1jkP7UY3/gsZ8BH2mq2459CHhc9RPfE5zAXUBNcZk1Hl+05cogPSdu1/01oXSz
uZ5DrzlUpNPa3SNkwGiDg3cebYSyMcVR5RvFKSltT4wHYbSL3i2L6CgNOrdZ5JX6
EDwhp4kV80YyZ3bug7EYtD2s8/pD7+gr/3xfYUBGiINi0T1tiNead/m8oNDVYWRh
7U8Wu8DQrNaTrZOwNjkevmaRBtmtGC9IaKjnaJMZLOnQwe710ssBRbL3AN7fpt+C
jauPi1r6xJ69xmH0jfRLmCWBD3phTkyECrE800DkKzY4XYwhAUxS71/jOk7z8Vx7
rKEnlddwEt3UirZCnHyjqKcUeOf1WjkogtJkz1cjr6da7XstfZAkknJy19Clyrof
ajC5ZszqttriThHjL8X2BmKb6bRssqFH3FS8FU1fc1dUsHar5ksDEFAbkC+ofjlz
3VAO+q23t0ttCmuBchQGLHg7bj5jNWyyX1vOIjmvjGZ5wD37V0H0SI7ubjpbDyjB
wLdo0v4NUZRwTowntv/UE2ZkYHvqH6CSR3ey12pUp9niNE/TBZzSmnO/sc1qghhp
1pXWzYlwbkLuOL111v2FARiYBOPuZqHiFPmM3IsNQgHPad02R2qTauvstwr9zi3W
n4unG2Uj5ZhmI1c9X4krA/4PCFal0IHdgEPoLXYpIF0MpnhSijMbmR/t4iIzu9xn
JP+Htl7SE3NYt7aIONC2qE4ZSVLIfgfNna/TW7yoiDMTyouflyZ8FhDcpK3Zfr1J
VEJYKFpP9GaR4MWEoRbBQcfiWb++IZhNH7txtZPAfMW1VjBqKOU/QpoLmQaJhNCr
PLGhD87TKBT4LPH8Dze0jrCVsrzatMWcPGD0k1FojFU3fEVys9+qua9/ULqDMeO0
WdQOO/6X/mxA3RiUdcZrL/PhsWBjAcCxDdyWjZcpFNW9a3xn2L2HXRlr80RqLcz3
CYQvbqDtKiz0xfsB/AjXzDefyJvaIIjpgCij5yIzGmMPMG0DU3feB5Ag48a0QQwF
6MWz35Xv4JUyQmgVWIwiypzTb0xb9C6Q3pnNmyIfCPosPdy827Nmfjwr0bgCbM+o
jA9TiCJb2ypaz2UYwY0SAh/eD0hmNIlwrgnej/Ex/jfe4I4GRHN07lMzPS5v2Had
n2ynO2eMILqMXfk6JtI4pFwgNZI93YdQUsQtD2PyvWZ/XhsyusI3JSDBB0xebzJb
M5+f7jNOv8OV9O24LIJvQ5JBH2RyFVviLGR9pw+hkhy1CugB7Thf8ELQ3vS5AxTw
/m/RTlaX/DP+zFLbCFobUqTz+28WrITV9ymEAS3yn47axWo2jZSPLJQ9qQW5LeDN
T5eB5KZuMdJfwdIH8oGKzP+Q7g+gELVg2Pjfz27yeKUQ/b2uX1m2eBcy4wh/Q8uv
OI1UeY5Wx8yKK3OS6sfBqTrToA18zFW+5rnWWGJSgBcpiAMXzDL6p6wio2BZiJkT
aERNQ5zoqZMvrOCXfxPeR5nH3V/fvNM8iBzwaZ1Jwbo1bOuwwa9MDje1Gd4LAcop
l8ARCCBoFuo1xwACSfC5ge6HO4MDRhZLqz2T4RNI0F14hXhi4V5/cf5y5QK2cfZf
rKKQnigyDVCRDycuMCkotdzbrhdgULvqAuSliBBh1Qnnbo88RCx1AWAexiYk4QFT
L7axW9QpPl35mkwgkLesehDmJeZyzQrPpFODqR85SR1cgynj9Xz0yKgaOcwdh94l
G0Q0TDJzE9clR7YL/9PUpkgaxbuAgJpudCO+Ba8/8V9DagQ5BkTHDAnrH6DBZQGQ
ps2yM7rjSXlJF9Ne/tfuAvFWAVCatmW/y3ZJib50fd1RQxQrQABKlZdbn9rffcVZ
++5W8XPFAhK6WuSRTKDBYs6EQox01XXCkaK9D9CXagtomM/q8sfOr3pJSJcY8Gjd
4CszWJ2JIyHFsWyWTT+MGFbONX27+FrCp3IZybZXrQxl12upjfBclmLV+xYrVEDp
1DEXmYlv53XpR7ybA3RAjfF+iEIVITXgMdupU3gUVUQDhivoCc+9pc+1gjIw3Gga
JBBWJLJbYPMSw219WCTHP3szYK1r4lOZNDqgKaCwSANAf8N+RPDncPhKZBhL0wAA
ZlEAI+P4/TumwoZcl0G1DiBL7DsNEjKBOKx0LZSCA+vZds2WECth5Z6QNIea0v16
XUTzobwn3riO/a0K3xdE+BnPfl+61udsS/IVRsFSluYU6R1C9NbaeZd7UZ0aA0aL
SjjEG9Uwh0Tj8NqrVFMp/gLO1RUcOA/Xsr2HF3ZpkS9AbkaWzXriXVkNtUKR2YRA
LX56oaO4zXzyHLzaG+KVhQ5Hhw75dlqe3hwXPE40n15RX6qObi+xoEkL3T3ycwvt
KKfq7VkwO2Q/VSzaffWR9+ah7joDdVmJHWcvQkv2r7NbNXr2+vLn/VaTO4vJoFEG
zpr4y58LHO0egdSASMhL+Hnb0EvuJKGoKc6rnt+/0MYoo/F7QBeFihXQIveRC/lT
OK26toblOkK/Dnw/IpnsHYEcTrVcNkWCH9DOepTUY28QlTPD0oUmo0v7j0phwsAc
K59JR4WcBdlF3lhbWNm9r60I4IGfS0lCQLidPYgIg3FRBAelvW+juGi/T7nZKE1I
KrhDqACW1MbrhfbQhfrxthY9AmlFSRJtSGkm5ToXRhnlS69SqoElhjo+E06sczAR
v4qjvPwU1rz9hmc4+lb0IprryT6mRG7GS3cgyYloaNOdGM+cyAsLXG0Nh2SCSnSR
cBtbdkrZJwdu0lew53aYcdORwQNOEfS91/8MxM9NILzLQjwYnqQ01Nfzf7iHeBIN
IBGVmbmSvg49SeaMNYBNX4ixhfrqebFpEAbug828itKCK0fR5W93PfKVk1Mz2XH0
zYRYb1wW5CQ/f7BdcxI4QaSPuituPjv61b1X8p2DMlIbA9xULqNRlwovZKPvBFQK
k0BSq2/nb7Fqx9bZKPI1mZlP0jhh4XcgiuLf+rYeP63MORJ58o0Abc4lahKXEaNj
tc+4gyJdJ6UEM8OVIfxsy7bLdyLF3U9M5nS/3AZ3hrTDKmtIhmOA0/XScXtj5nXQ
79ldzU8QNrLwDLXsSNQl+3WWr2ZPBNncJAAx2pnY4cD3zfDK3C9cjn0klSrAF0Pq
19na4EBqzstI71LcZZ4rZTS3gRiqSekZvbE97qzj+ukUHDCOPtDEgaVgmeDXZE+c
t1S0vDfTqivLiYb8W0+aGgdEnWBLZu/QzJvl5Iirfcy55KPBZO0M1GAU9AFkDsJU
Nvp/7S94sl4q1CTiP6ydUV077J0LZnIH3tUleVTiPWJox9oUHFvISXD9p3SevV1Y
szlKhDIgX8rJSaYgCNOWFtwS7gVQFnl8UxxjHUj6PsLC7wXfrL1d/9jZU9uXVEMP
/oxlHtAGcJsB9peEAg2Tmk9FtpQ9qDffurFKTsEs8SWvlXeZ3j/th4nZgD+SE4u3
zkSB4qL1Ud12bOs42AbKaxe1k1rq+na6yZjIxHIUJNCa34borxdsGyJDkBM80FmM
l47/V1MJDpMcxdQePaOjs9hCAPzU6sr/H77XlSnlw+zXCJGBW2CwOCoJYSD5bTR4
i9iDyRvI+M+hpEGqXiUiWjF3Fyc2eNbVjO+PCztMzm/bJwrinhKFGhpVQVDwDcK0
qiunC2iAVAs94bQWtiAwLnHESxuyjOFazlbwuBHfwqSmaf2YY+Y/Kn00H1o8VqDl
NgRRyfcJ/1O0MdlQsmgpzPLhlw15yxjX+qri3PSYQ6ebwuF1LvNaCp5H31ThhV9Z
i3/MGjBYJ6TU8AWJmZjiMwcv1bwo/x3GGBEWm9vwz0N3TKGpfBY5cjGUVHZPdTz7
0UHcYiO78bKzzMjVIGGqSURWq/ZMuLxexSBeNgvOPz0L163LfcOp6K0eAHzpE7b5
hv+9LpJn+95m9Ovt8aLzbVhpxshm0A0guNHheQtbQ/YmL0xJoMM6ZeWWznGIrL3Q
h+Umld/LpldXTk9qBhnbClV3LdEeX2UUK8wS3ZWyVzMgzCF/VPIfJmVPp+ukVyz8
tg5qUz/tN61HT8SS61IEI88roSMzziwckB1dFbVAPY7OrNBtfJyV8jI/189NYanY
mBQ/zU9BGbEdvCPk53oRvaFRCdwbTqaJv9bJ5r4epeHheZ28DieO+dPD7o80T2Sb
oWUiSdHlJaKwO1fwbBfAxsiOjm7dHeNi/RIf//H9XNCHJ8dAWDngvwq7qy2fghaq
m95GP0Sss7SMC782LPKuyL/hBjH3xlRnPlrczeJqxjZ4SlQ1XsCtKlBA5KSX/Hwa
bIKoeF9tGgtHp3nvLUTvteRN0Jarb1Q76uCw6MGQVUIhy12tFfnUPzal3qMc9em/
hywoxUvwtxZnWzqtnD2mVXb/H/YMDIdq5Hc1FNWZFSZCfL8aew0neMCfNjMGebae
0y+S9Ue5XxdsJkAegK2yx8ZBAJGKXb1pyglu4f/Oo9OTu6qepkkopWF2o9HxcUyM
QYZq8KhrEcqRdTC4l6yyD5p2/cLrMbw0v3gViRgeBZDjCxhtqnrjC3z57oGatZSM
dxhekq3+Cxsu7aJxi6t+HaPqNvv8sA5uLgzbMdaGu4Df1GFYyFvUjDN9BLiKSz3q
aBu4N5FFg4QHM/sY6/61BQ06T8CAnohFbCeXOqvlMKxvLrkwmMFDR46WWv9lqQrH
PcfRCBUUDau0F253XEVyIqtouIFxLr7Ccwy+4xMA7eK8+hddLPFzq2tMt7tD5Ru+
9ijLqGA0qKU+xTd6T8IIo3um+A+zArsUYwhWguPsZ10OK58bNx9FXNTWJqXdeiF9
FSXKwfFQvaTZpQoQoD8ecvHEBDIore3EVPoDKFNlSNLr5dbhPUPFJ86DFQan+9hx
j5IbuEjRbBxe/se8+sQBUhjW1mw9+BCB7w1QBdlCWOdYFhLzGeQ6qEGcOrgXDUYx
r1Db4BzBahuZE531plRVo+VDHuCRESvANwR+5YlMWW1hCXoCVEa/aROyUUayy7/h
TaQnCTmp2VygxuSH1KVpnuxu8V9XOS4wfKgWAFiHJJIRKNUe9czv2w+pd3YuxeSb
kp3EkwIRJEbRKtD/0ZwDPcvicF4sAQp+M1kmJnIAVCBoty2mV/T+lPamZiGwcv54
pHemVQMLFSmKcuZOSbnACHnCHAUPchYU/gsmcH4KrZmTJHggqcQnwbfN1wrhyYLD
ML2p+QOxoAb4a83Ue6E1k0WuhNkr5iF6qaXowuQOzE4TsNiM1k0/acEOC+/aV9ef
DtXwRczOUicgXqi3hMfXvF3wuTw++OnjWWO7wcsYJfWx3mZVPs832tb1d84NV57C
OF1B4EthGxelYBEfgqXX7HHQiH0k8N3bfjHfqbMSPCpQUmbNe2IE+EVq39PlFMYH
4UA2bJwchABOZwbPeH0MER2UmT22SG6UpKUQuOJezoTI/rydQOVsWWhcEnOt7Qnp
w5m+6sXjsqNuiB4EDdSZPHwYpZkz76U4ttkyy3HCV8jdtelWMThjEuUpQFnTtsIT
OLmVulvL7nuipmGP9rOd4RgrQRmHqGVARIabO/s/rs4TG+p/YlcD+Eujl8/HCm2s
YiBWYUlPYsvCKU/JPBeq0twXUFMx1cUNDMwSmnfwaAK/2utBtPaoFGqMPOOq+6Ay
8Pb53zW3cfRBhpuUE6f4jG3Yr4MKkFuskPWNLqBaxjT+54Fs4IzNABgfe0Rx7Ox1
BBkaabRG7BKULU7XDAvf2MpIuZmTU6etcl1+T354aHg0+4YDCwmDYrBZvPKUtgYv
aSgENRHP1jVGLB9N8u8PHN2k1ND6WbvdbeWqI7JD5mnbCTC14M1GU+7QMOtza/Fn
lk2JqCVFGY8oy8Z+Jl3+dIB08Lmh2jL0E2LvdxyjyaxXVon6zkO71lifsCLJx52Z
r0QcDp3ujJSXs9llkNLTmvHxQTL1Nz0IYwszYqaTQ/dUS+6XiN5/yB/h+WR+5+sX
eErVLAj/OwFQlOCfVIm9OK2V0hD29QPoK4DsbeNcHFMvsQyhQsYsJTtXNJQVVF2g
bK7AcUPGMKqdczU+O+hQkw969y4XzvBoLMO/HkgaEQ8spAKH8toqXWriRdLu4ppQ
KCH9sFdxOlk3jLn6vfzYdUML7M5M2DgnZn/cwhmWWJYK5oI+TTbLdgkY9DIXLPuB
U+iPAscD3kdPdpyYOWxGn0Ox6p08th++B889IQex3madTiHalhNA7XMsrYmvmAWC
OSxvtyDiiWOdwm9FIwmJ53qqB/e+3D/GHa42/OEFNY3k3LSiGqWCtVHhTkgHavrW
z8VqenKBZ2UQTf5iwUNmuwPV3qJlyavP6WCojoqssf9wFiA/i5p4R6lriynpzgOd
PMKZeQlJinT+UH5bKw3JNwFEkLFOqfJj4XRVmBP/oAUw8F5GkMYqPWofGIV41FTJ
/RSbfFyHJx9yfkDG30SIBQJpst3OcGDu3FtcRg6mbryV13UgdZ6e4kPSLPyJHUls
Cz+NfsTubm7JWNPVjyGcQI2LIxiuKQALP5wYVhi0DzBa5WUFdiG4JbaRsxwzdz15
9WW2Q0z681rRouYsDPjmFXFloD0sYIkYQx0E5dr4ZYYlD2sy52Vw19g6gseEEEpV
FGYNxFxRLGwmxHW6ZyQkzpz3lzY3YgCe37zTOj4c9RnF1YTA2lM4Ll79wjY5fzxT
xV5khqC1FynjnPpxriHMZPVSrD44vX1m3cgvDmkDJSYMksBBzKZXGelD5VS7PIpv
FXaRS9BM+AmwOMDUQmJJ+Crtrqe0twPd2iCfWuVbvE0gkjX/UTfCXyAPDtd1rZ04
JD68FVVbEObTHXbd0STF/hu8VkBA4RnXVgBSDTzZgRYcXyGfBxmTcfr9HVbC3SmP
x9GyerOyAjkA1Pa1rq1E9s3j0ONoIrKddvRWIPpzw/bvOEYAhOC8h+Y79DbM2XS+
SLqQeYmNJ9K2Et+Hzbcox8KsLXqlDb4V2IHrTViFEqEAUgfLTOWfxGKChjRBopAl
Rn9EWNHCWIYwFZ4rPCyo0zRlp1t/v+kVTo5rCwd0olZ/W02v0hirXTGk1p3FM+KB
l2LHMWHiz7XysgY9QeehwjY+3IWlXlj/6dwQvpERDDtZnkRxwRb2hhETOo+3kehR
IRg8/ddWseoYLMgnPy236R2fsRFFGGOzk6L2RggfzcUoLUWB2F0e4Jb+MNmdCmXC
x8vpG1NWr0znlZK0rRFATawsHcVC4DHRNvOwEYkvdNoBlJ2DKnaWG6y+Ite3dlgg
qv8FNpVZPYheSjoaVQmLkav5EtiHIwwiy3KOEb/2hmPTceQCCjr8UhNHabKVzN8v
WcghLOB6YNj9EO8ncYwYb6jLGWG5iQkkp8B3x6kpi255OwrCd6zmKk4B4n6YTVJw
Ywl9pkfQ1/Y3Vy6GV+OgobpjQVlPjsMHbOeDSNYjXpJbwWqfMPpGDZ2UPo4q5U17
e3Y7rgeV1ghNT2eSiPHspBt2JaT4Jq8HE2ovJ576t3Qj5Oycm5yZCJLD23R06281
dIIEByawZfNfRnWoTwrA0el39k+JGb+4+YgHwaynYkl+cbrRjBTjKe3PuvwM7qgq
kzgteh1fxIGKO+V873aoWQfn++1cOGsTu+qitjcNm1GK2kFiVsu4jqAZWHRvim+Y
TFSBmhwzkVHD/UBxWfgW06Q2Hgg9UxuWQ4n50NE4UIr+/oJu37lTpDpWhnOGo66N
sSBYl1FFDlgFoduOAxtjP5Gfdc9azRY71xejuP4CyRCl07eBhrHrYqKHJ35sg86u
Cf+RAWBCaMFFJyqVyRsagta7FTtnpvM8WkULnxg2jxTSt3NMAwu+OKge/AEqmHxY
uZ68///vx90PicUiEVMk2V7AtNjETgH6R18Q3kVy2IkjEdvjqwRU540zTkIYUWJU
VopXHEvx/pSs0NdMo0IIiJZEFC2sbNQ9Yxo9vNaAcPkcn3JyS0s+/sEcvhGO9LRA
gsx6RAlZdUEkM1tW3E76DnvamTytb6u4iZe4CluQjTcl3FOkY0R+BfYtOqf3dSAX
I/IuL9W/OQJWh2F+xf7D3svCJajakp/J3YZPnZIX1Mr2Szf5NKJwDu+49mYHKC4o
74zcuD1q3fkZa42HprOKaPGFVlLXuZQ+Z68obZTj9yYVaRr7belU4KRVY0apgSJY
5pEYp+XsL45ZLD5ruc50h2JnOQpeeaWAD2oqbgqEjmzhbQlNBC7vKlJ71DLHHBrI
SiJaROfAYA3RCq/54t2foiIhs5BXQh7vmk24mbHBBSek0UlxRXfZP0NYnkQRxWjE
YyvmoVvXLKXl2OLsIR9csY8T3QODJ916HXkjaqaA5r/MBLdo40TiyKFduTPgqhq7
Ptc9a6YFAFlTX7SXb7DbxX4mhmjmy4DWLvqSXqL2iK0VfZHXZYFvXWBJ28/P5hbo
XY6EE60Shm7D0koCp2JrDWTVPwTrw1KOad9Mg+dtIyI4HO2jE2pVjr6y6mi9HJ1D
WLO/1iW2+nwYvKcBh3iGsAKujOIsxVBFe7UHKdE7ISxrV86RQGRyJsTyu7J7aiCA
AhA7jfrTJ2RYiakmkNu2ZUDPRd+YL0b3oqsFtX3VG9hfpZY6qlxZynY7CspcpoIF
rTLVHFPbKpviep/Avd0B5E0afYQTgGJhIg1s1wTDUiqEyqP7ldNHubaJTwToh5pR
X/FlKBML7ao1ay+V2jOXHSdJeHHq+urEukY5Sve1qlhJ1apYo34U/4DQ6J8aN4gy
hz+ldidPe+ymsvKtPpKCDwkRr/wv+oVTUWnB6VCWwT2JxMAiKz7nOwM9hEuoX9LE
By1rg5UHbK3NZ/LKtWKOxACDWopDyGRC9b3xH8sMw3ox5JY8ZwYnhnE+MVyZkRWB
oriH27XJtn48ltWk8ZubdKpjzSwHbI9w2zeiGaOraaaSmCVcVhecEGPTBNeCXEjf
+BUG24a3P9oFfp5mu1hci4hzEhSDFoslTfOW+eQpxA5IoHUMN4MdTdST9HkAx1Xm
Scil07o6PMv54HmaFshWxQSCp5CjvyTmIqJ04CDjz3R/geasbdTt2o8FVPV7VxEP
JX5NmmtbZljyforLt5CHunDtrnBh95mm1eLO3gzKybI5XFUQVCKp6XK+Yf3ByLvJ
yXVlBUPkQP+5SwjKtfUJVebkignrlRSOtSQCfl28ApkMZicPbQU5CJ5hXQEiMEAY
otjCDu8nmDjqHYanz6VRsWgMHe1E94W2k4zwObIw3ktLzWqgdvQY+wDvuAWcrsim
3+dUvZE48EXWBqZYMXlHAmK6tlHBlR+wRq+MlN/KINN+nV67TVkH5kBDLwmxdrKJ
5JbtVJ9BUuuu4jCsKup//YZkpGTp+TNrJlg/AhgPSaf/Zn63G+O6P7bSC/ajNgPC
nwMcYRSQJnJWiHIEIsMuswL2ftcla8rcbamo2EqeinwQO1kQIyuhtpmv6isOT/oN
B5yPd+G6ssaPiQ1yYI/Hbid72mgeP9Hw5PEazmlJZxhHA75wsvLgadfnrVyoxPst
CElp09Jomp0Ardmbt7KY8JO+clF8rU3zXSIjj4Gw+diJ4N+uCVV8NtcYn1EX/aEZ
zBGJjGPUU0IlxYHC0x3h01YAyxUA8PuGhxnC1WYGsaF7lXiTSjftb6NfKTA8M04c
Mkt4yofvmCQcewyj9v+3fMHbrKv8hWbLlS5B1c8XdpwyjsEkRQS3Gh/dC/gCN2Qo
3NlJ/u1d7KR1wEeilLfXNbUp7wblYiKUIvLeiF6SwAkJKFRnRiM5oREDHoTGF4C0
t54bBAVAs3Ogrbz7v9HJR7dns3l0nl2lFhbUa1WgM7IWoKljElzz72zKss4/B55v
JucaMYf/usEYrcNGPZQ61HCK/UlpFBSulNI2KneYi8nsyGj78nJ6wmTaCmVjufw/
m7cnJTYyLx59eL/viZN9A8hfiHsNuKMp9809pqx7Gzz87XXydRkJj6HAdZNZuE/f
li5+qht/6/wuHboYgsOf+hqRmKVDVeAjZB5LFFLFZ2A+5Pxb0k/BTmuwFPulnMlf
XNr4ly4RQvz/fWHokKkoLCMtW7H9KgM1LUepkq23+W/vlKvBnQiSE/ImB9ZWAaJ+
sg13Ti1mDl1ZukXvBxl3YwB8IwHzH8ruz1n7wtRNVLPgUfkHnaOLPFLENxhh7Ta4
BOqSzNRj4QiLgKb8oLnODcB5Xm23akOYMR1ebjk1RMwQ3Te+xG8FuTX6barFejWu
1XW6ic0bvVvGEgWaOOrCem0yerULgY6D7kxpewD/+fF/nvnYGUEGIK4WhsvC1vhy
BFwe+fUsWyWKaifAwYR4tiqkyB5ToynPz8UIFsFT5MweBX1OJTutIysvDp5Zzgsc
g8bIH0TU0Kdkalp0oyF6l7A8sztORGqn2YxjkgQTqV/jVsJteAfxpthx5cqeI8OU
rfmaIT5tgBrEGiy+5pYUiNAQJXw4RIgFq/mHqU1Kz+h6RkibWZ4GX7TfReX8meaI
JtBISo8FfYp3NYXGUvDRjp5wWg57TVmrSQUmApuh3Acgf4uKa4PU+nKwwHLG2e1u
lyN85UjgReKAQus8utUATFDUe0BI+DD92ejcua9wgF12/0L/8j/idvt1n6w9nfLn
vavpraFabPPl3QL5u6/5urPlAIx030bFQSEEOQwDbRU8CssKAZwumv2pfHQIBBB4
3pDoyEQfQY8UsNY+wVfr5uggLpTJgGm4t+z+k2SKiHhX7QzYXk8d4FAc29FZD7pv
JCPdwoQq2tS2FOV7AU0e1mqMDSSQBBBGnhSMPjgNCiaKRzFMHQLfJblSqjvF1r7m
SvVJlPV4xBwda6b2iDgnu+M5W0myLn6B2iyVjhcsqqPQ31A4HXeayQmjmjlRcDgZ
HlK4QdW5jiQWLvXCSHLio2oUZFAoJyolX2pQ21sduKV3nXwa+avzaXI6D/Vpwhrg
kasFV+Iystqf8te3dFHqzJ57xTvfallXV/LLYXRYU5Hql6yhsA4lPAvWtDEXCPHm
oTai1ek8a3LYolmhPBFOZp7yboqpYFRiF2kkLdLqC+jlym3NGZqabsaVc5+WKLgD
AJXaP4POdh7cX1gLm7B4VgWC05E8KDNgV0OL1ntWfRQPnK5hwINnfdb2yJdpPx8o
VbqwlTFqU3IeT3eZTqfl1Ad2xoyhKHA4I02XitzEAHwCwGvB+JTiyKZkjmNrByj8
YRPlRI3EXij7sz9o3TcxbcVpxYb5xnzyKB2CCZB+0NAhUVeiQGZYp59XvFAkrLvp
WuUGOG3wEIrbq2vSIBGVfGYc5/KQeVYY8TNGYy8v/4kljVqTbApggGk3q7ZvUkHw
7OSV/gSvRIOWDzmc4BYkpEp82iDOqYPJezwhwjcd5Yo9xSFtzowkrojjfiJNaPp9
LQMl8fkApU9MjvFVBJDCOE9fUHDoT8C9tvD/DvzixtPpkFp2s/jBhf7Go5o6ozal
+VStAmAFLeManu80alVm+D7ezMyDpQYHNQjVNxX0UlIUhaTDX00u4wMbmhR2Rl14
AiWPOBfqd/1gE0jww0tJ6+jymqcx5Xyd88GkLgUJfHSXocA1e3WrUuPl+GzTOd8w
y+g+4yKZm6n5O2KZslMLNvB++wNScpqL+PnJ7cvVHWSLR/Q0s3lxLladL5vqLOu6
mSbNWYsBuhXg/BF72wJ7n5v4VniRGQdCzbDRz81mqVufCUucgd/tO8b3PS21/ESg
YHECaAHbwiKkF++kyApr2Op0PmwDrJDhgxeDY31awKzulnCQWB+qLWvs0AovW27g
cIOhXdcEpojeJnYOlnSkuYOdBOVn3UwgrswIcF0w/K8Zr8Awcj8WCEjvRLjtJtah
XUoh/hxXcuNIDG9ozcUQNcACfrZ3Ol8MdyaeTcD/bQ3WHDdkj+avvITAyGpBWBD3
BNMi1y95CrGv3wPF3fID0CpArZTQhRl2shj30sIcMhgfwowHLNej4ZW/AiDKyv9a
c6ssmqyLuy5m6CePalmaNCnZMrLoN45tDrqqpDfcakZOEazi1B2r9mVgdSNMq93U
sXLyB3NNeYk5XNzevIB5tUp2X7Sask5m3AzrDlckCqQU/srRfPF0yFGfoiiQUWl5
RN8b71eLnA8EjxhhEC3msecPDzMOkRZh5V+NwJttr1N0fQwiYOvj5FhDb9aHZBsT
89uEE6Q1K6h8Nvx3LFrAp/Rm/biU2zxrAgIBXecavVgkDhNkQQkadOKbhNZdnRd8
WoEqEKZ8t91qOU1WGAbsZXvw1fofIETuiw+JAua6STs8627OQG3dRn/8AKF8wGSB
d6nfzpB+CRNMNsepoZL3e5hVC3BGhQbgzWR5xi2AgSZkxwMgKz0rZMvm/jzzvDHe
bPDYiBCXJyiotptz86qd58BvYvcZwVbXMD8UvC54sf7Qtyh8YNnzZFQk/zkgF8va
YfPII46cc/fERjRFt3suZib/bAmRmmHZtN+Ab0b0tkVSaoogFepvlYtVsyzatNNB
0N7DxrsVXOUAfID6WZ8Ll6NQmsjNF3FCffkPhVD8Xn8CjHnva3bozQphTzOMD8GX
BCTJOBRSAcRb/VSBvgSTvClWaXXFIHrmMNLgr1+mnXM5mKphv9DTman8JpQSF/hj
+tuD7hNKdb/gmY44bsMDCPyuZDtFbsNz/R5bhkU7P2U9wMQhf/oTAJ8nuKH0iqld
1PcNxxiA0W0NDVwly+wZUKcXX6yu/gnlcuPWhruVGckLGfoJJs1O7a5Jsv65RHeQ
5rMHh2N5A3aUIi7PqLYkOSyLS3K05I4OAoVbBqVd1wGZUcps8eQL8ZzY6um9sKel
IzqAoV/KWCMGYvvGdEHmgAz0X2OAj4YwkGaIc/9iILI6zf+g9+z5TA/B/roWRN8h
30BlAjy8mcOAkE6OSlXQxWWxqJoIwFE0My5ybVperetraR1EmjrqOfTm39d0p0mM
oFzWsP/7lnRFXBpD2lH3UfCkhiyhkwujOgZRv2vSMg2nyCkgEPuMoMrF9LLbaVuw
/c2KLx+RQscQvI3g/24vR3epCOS4EgfmjKyO+sGfdCh3CuawOSgP+OdJv9CYl4eD
Fcvqixh+nG2vVsJxbvHHF8jhkWXC8VZiwpBl1GdgM20ONGOKey9YKBzbrSNkGia5
H0aCHATJeh2wB9mr2VYheCrdlMmzX6ajy8OvQIa1gf5iO8cSstp+mZ2HO5P27jKm
818Oo7/LNkYkk9uwn0e49+nIsMjNVGbh0wufw/4XJIdUKhxdMEyaDNcv+U/IPOzN
PHdAzupKkr1mS5/UoY3Tbaw2fBenOfZHUcsHYUQFGqK4+Xv4vNiQEptEWM6BKHMr
njZWYj8Xw/ekS1u7fY1ilA/b6JOh4AOTv0+elV8+pjER8M9kB15Xxvd4uv8Cv6HE
LvVXPu+Ed0QKflQ0cdvBdNgbtULR6OdKOaCCjjVeJ0HuW+VJdPeJZV6soBWkqmAv
UC15Q+7w6+91xO/h9wqDpvfv07jF5elHgLys+AK892a4ZdHTweZFTx6FpQA8rJW/
Rji6lMcGhKEkYHoz8PbzBMkXJl2FvOshahepLmCAYl9k/QTWB9fOw+2eZJjapvCj
dz47jsXLrHtoYYmj0kWvABb8/thulZ+m+yu3WecYjXoH4b1Ge/O8p9uqZEEGU44y
Bi52j92icP1OqBBlcEC7rVNU6FHU86Sv7dGSFbEw12K1IwQ25NxIAOoP5NE9IpXU
QS3Axsy3CszRgfqSd+XvI9gxttry3fcWWEjtly0sQQav3PX7hzwLBpOkYdo0zBR1
+QVOJEumF+yryJsLrb8ajBofZZK7RwQWT2zIB/XVUu6p/Lox96cPzjEv6G7TRC1g
fiafB6z1DOqT/njwGjqsp7lVnSPsGSj1XLf2bq/e5DJENOWAz6bmtozta/s0SfAM
yZDcyFXAbLx0rUtS6j7Qagpu50OXbfALmh+rDR9RQioCYFIDa37iZQbbwg7chpAM
Y/rDam4pHuPa/p/cRmg5wC+H2dXTb6dQxk+5qP7syhsXzX0hDC9jSi5+nhxg3gwy
CIMBO2sJrioRj3hXtoMBhy5/C06m6JnxiD1/FlsRihLqzP3p9lotxpZ1xuGeGlv8
HQxeoB0mdyznYSFmW+1Pw4ggZOBRWVPgFmdn/zV//wddXeEyjgOl6KR7kDw0nntO
jfJhVTukqaG8unA+75OsaEZsZiwjZcr2mjHKMQAWZVCSqfOerw2fxPNF88vi5u8x
JNc2wyRwhVT9L2EIbUTHAkjGHuJVaNbKre8vWRzCfS+Tq1UO7qcseDzjSU0qNzvK
b4qmEcp8ry3b7YYbKyyH51+HoOGYIc+DZ+wupJH442/KojsqFPWwS71ukWk+5iUW
axkb2vY4jFXH8HRGdmY0TW0CZKnf/fJMSDEI57NJ4DynkOpG1nqaFb791dX0/T7s
bvW4NRtnXha88VDMiDzDf1ZBlH8A3wQv4bwIWbW3j3uC2P6pdqoBFkIenwxvi+1j
u8usB6Q/39MBLp10hQKQom+TNMdldYszJ0b+PzlffQYulQkAzmQPSP7Yczys4Cep
Q5Q6te9wFjrDCcRKBmEdZlJRrVi5k2/C1fS9g39uCdS2ynMp2fnl0QBFxFpWfoxC
Sj0dpzRzeZ+IMviFiXXSw9dm1DUXRc5di+TyulDc3bbpNOwmb6EMQR/OHvStnfjX
jmVWIpYvffmnmScmkU9iAjA0Lb7lpvE87tbmumBNaC4Pj8YXRFOUF96QFIIvBZOq
YxShea9cPDcB2oTYlxUBg+mTZTg5Hj4Fc5UwkZ7wWckTFnsFiscHm3WkmoyaQMRR
pwZQZhON6WwgoHpqNuAyHPWTMOBq9AtP+445WLsDlBmZVXe6xRbDK3qK2VvKg4Qw
0z1E58CaJXLX6Ev4eemlsi18n+dLIFyK+EXYMDJX7OSMVUKfl5PpbxPhMW5YPBCN
ONxN2kLl7CXRAqcq5ElzIT45qO2VRQm1VDAeI7x7hLcpIjENQjNlW1xM2tWmWMy+
z2eS/O28dnzSweeC29n8xxB/jce80OQfEn1SJeSoW02F0O7+MjfZMZAvbhhgrEtB
2fbX8uf5r5TnfdHVUycxIVy1udx16Ssx/kIL0Ud7U+gdK/ZDD0F575s5h/ew8PBQ
uZydK16xk0AOH3F8nuU4j5s5zbGDHeE3smiuOhQRJdZ9/CTdQAdRxxYP77YzAxnC
8+vYfskpCBBHyyOCNJ8fDwMggs+yUPvHMx+X8jt0Fgxlb5gB07EQnuxrBmKmD/rj
k4cOuiDpe5UQ9Z1wAn4sDxps1CedSKuN/B66aojnj4cMfPhe9TvU0BQGw54OFnpJ
4LjGo6QES9dcbl8v45/M3So5mINLWF19MZyVNg9Nf16MXAlN0toPE4DGfAn6mEqE
RRuB2hjFZXoctjG6AtyQSGr3rVd1jKbh40QgGh1T7QLLzaIzo7oP3WO71njlbxnp
YwVVEcj6pXc/zY4z3GBt6Sm6O1CXoCQmhvHBiK7TpJcs/xcQq9Nqx2qvWm7aLmPF
Cyw5oniT68y5R+TRBOHFsTC5gD3mRTRqDa5EYI++6DIvG5brmUeR5p6epBxHderk
NeoyyLuWGF2gJmTZ/PPNNqgsBFT/EhgKQTF/Gj9SQKfoQ5USP/ukhB7UrGqtbP5Z
nc13t104CF/osXCCXEPQRr0QY7fBre51AhPD3UBsFfcXAoijOnxY8OWIiK/goQdI
LTryfRipylr4HWr53veXWKXswCHRySCfcwkU1Cy6P/fQEuEWJY2gChX7qjqWbkOR
FnwiVoGML45BUpI+9CXWp0Vy4mtHmoo0kgdlvwfMcJy5sxZxrb8KZCV6a9Yxj1h4
+i/i9MczpyV18/rRed5XyM7ih0e9p975wgUVkZFjvor9I1jMrGrZWtu9++Wy5GQz
O4LNJ9mlXi0A/c0XvTOEn78NKTYsm3zxcgCHH4TviCyr+Nz+s2Vqd68rs2QIIgbp
RsQuaDFoH82J7Et/4mqEST2yMlhv6OODj+Cy4KQfd/zFq+eL57Qz8BzjmyDqhThV
3dhIE6qumVBmX3htGUuNpTMu3EJUZZt/HKZznc7XLOnaETH25lAsp6PHmXZj2QHI
lc0+rBYqNx6EsQn1Sbl9+Ouft6ND/XwBIUoHe7tUz6bLz3RCYLIAYUzPgTKIv/W+
hZVBMdHCtZllDQgr0KFIR74e3AFAwxZGlNTcXzkZSlsTyBm4ypyWNW6KR3yae/kv
htAsk5sG547XkOhRUTDCbEHjeLbE2Y0wbClMR33RwhwQG3TdLr1RKai9vLBW0yA/
qkRzJO2m9F17C3cuodYlvjaok4PFX2F7BmxfYPmwKychiMMXpHqMu3m2ETL+vb8H
MnjyLLz+WYud1Cp8rymj1FE7d1usuzmfjE6mGEUL3zTxuj3sRJ7rv0TANpNay+hS
w6dXESkGI39TsfWDY1SUc8Zut9qsNS822BhtPDvPJclMexkn8M4J1j1BpIeOg02z
WbOYuP8bAqCcG3F/J0J1FNmeM6lN4ijtn1xjhXl/KrMZGNnIYiHmY+P09s3yMSjN
eeSrJ8m5gm6AMZiLUjqv67tXfxJK/ut3VGVIvr3oWphT1SMBVUMDJGAXTO2j3yAW
PFhJoCmALkKGt99JIRx9zbQVrhe+5t3mya9NFJasySiSXTx8FhHW5sEg0cS1cdE5
4p87ifQI5aR0BPd8723Jq9bLj8Wncth33sBmXXFVi5NFpXIrofhER0LW8yu9sLrL
6TyNFAHT026at1IXC6A+VfeA5pMUSAhaaVFjcJ2GI+pzQ2WuQpAnXcrDU5DpU/fr
URiH7w4sgX+Mu1yzsdrDrcHea0H5AAlWJ15asMXeI01AmIxGvQ5PxPcrd0EcASpd
c7DDlX9k50csEFSzlSEhRCQyFbuzd54CYltUAicW2qF6i2SmjfwTV7zKx519HdWe
oFJw0WpXoGkUZSYlc8GJfxcKqa480iK91Uv1r1ALx2fWKrGe5sVd8q68YUmqooZH
xZUE8G5+uY692m40S9d91RclOcKmYd7BpRqSzKV4u2FMaret9VNYL2iyPFpXHKNt
L3ONF7dPZIqgkyKUdGv7rj5Gg4OG0AJ+OIVGsd8qYNurH2/4ubQ2bdWc63ZATLFt
FvGdClD5oAJwpI8Iu0bN3hcwryaMxoxUwlhBN9B8H6zwJ0u0MhqejE/oLLg0rxm+
rjNQ6y/4eeaVnLI371cpg5w0MnaK9zWoK0kfJJ1Eiw+ne1F4V/3USlwOQEmaqVGi
Gm+cu6BRUgR7wpWHpACoLmu2JByjbGHeOs3okRsd3gLvDRVzR0umlamKlsZUTxTB
hetYVZgsFOO0IIl3dBJyai3LvIthnPAU4eUvpq3YkSBJYsppDbo5zYjgz1/aMjFb
y4LEL+2lAllHghzwGz7K1Z0D2/uoaxGAvuC0WLWGEAd/SH2VPXYu4ABHUkxaRbTP
KVKQhPo1cS1DGs8B95OaH2gPDWnzJ/IDeTqClbgVtx34jRUHbWYN1iTdFgi4Jg9f
QvLiTejXiUD5skTotqxCF3rKTjZF2HDgVW2+WuzdR0mNN7w18CMD5VffufvSoKvs
9rysswnLAfh5ZDZOlfLD9UQL79mMOLG8H7D+kJKOkXUszAagud05MnH1VBoy2h2R
Ozpw7yv1Z0v5mmdkoIfS+x0MZh87f0ljz2pgwB6RPMB3ENohmz1HNn65kULf5h9f
Y2Lw9JVbI27DxaZDUvv4DNBl34ApmU2cASvG08YH3HIndGTXDPR890mmZY97VIcd
FbweHc9eLL2lBJcsOeRbsD+YRqm+m3WHOWTWCIYbPKsS5rpuP4S8X6ySzQqv7fVN
XikfpGkS5bhoMQcoaEgeho/XvNf0Jbn6lHEbPOvYiUuYGFp8OpLrpfAtu++ad8UX
vRqdSSpAmZ65ZJ1KiEOP1d9JVrSA2YsnzQ6NyjNbU8cWHtJXd6UDDFX97TFkhznB
pVUcb3XP4MWaBrc9+Po+KJYOJqXnVT6YmnKZ9QLFw/1dmp8tGQ/jhWd+S7k3RNVs
iz4Icp4dg7fzb7lpvCUsxvXuIMHElaT9zw6fJUExz/GHKZnS1AG15IlodKLJi5R1
TGo5fNurmLTYMM/iA1b0Cyea0YE3mYqEk0E506pBKdJFanMO0oy00aWEPn84iirR
7vPEyG2/mKnOzDGwDmIndeS2ypfegfmnDMVxuNy9leUsMe2VVsBrD0EiMdcyvowX
t6lxYIYhynrc1xIcoidpIajhAZ2XtPyD/KsO2wkN7tMjTpU6tE8fKiu3Pa6rJ52H
MoVhppl4oMwtLcYlo+cW1F55MxRKsOsDMFBJTCyO/LfjPXfeO7y4/t1kH3SzUWnM
Jr4B+FHz9SHKGjV72wIQWItFxYDCqXxTqfxNvuT9LJPy+KqdFxcz6S2QKvXv37Hr
1Ktpk3DedoxE71gJIEV/wFmyxeFkWkQ4JvMYk3NnoE5m76Q/9OfCv+THSnY+Yhza
6S0rX92q06aT0fpTTNrW7Wmv8HM9qmVZiwgf5rYuAXmWv+xZuTxOM0sP3FzUJlbo
XkbI6jPWgrNZ1HaRoF7Cy8XHbwz+mlvXKkTj4AG1rOWvZnycDOJ3EDDGBEvxbM9s
DBZG2kmM4xLkwm4Z3VWce5x+YNy5AOzBBCjXGl3Et2biYsd1z/T3e+CFplrfJ0CW
NoxcUsictSKsFvc5xilreJFAFKx7EwTD8hVf4V0SKiGQr2HyzYksmxyOldvoa1dA
xK3u/tYbFywjRb/FX04MZ6mJvv/7sd7mcbgvTzD8Ah68KKvNLSE1Hnw91HsHuE2E
OYwx++fhLMnB8Fc+kucyBBTI93ZsKwP03BPeiOw/YOnTSpCpoOBB3nbfOOAQzsA9
OE7SuIpMyl9b3FzV74cVIqq+bFAl+4GkpHtgMqIs0GCSCGHbnXf77eRvS3iVAfxa
7D/CBWpfHecZQydgCuB8SL0BY6T1osTxxjhjXGT3CbRL85yeWg+HljaaGXQGcw3U
TrQEr80Qa8a74iwRVan1If1gcazqs6aetX9FID31vRLfTxHJce4jDHRt1lCP0D4F
5eKE13qoxJ2tAmpQmLGx0DiTIHybXubz1H/VprUHkgCrBBm4VmqDSmolsOPg0ydf
xDFAFfGQyt/GQZOTKmmB64Rr2kL+29K4wGnV+qd149IgMus/qdIQpDCJZXbN+cMG
p13x50O6fRjnhsWwmmZ5CqJvGXpg5wsTRrP7fngeB114L+EjZ2VJRvlzh/5FnjvK
WbFQXoBsKqg0XUis5FjsDuxbCxbI2QTaMgXFk2cgJl8OzAX/nmucEdiJ1xPF671O
1u5ky0m227Qhv2S1NVnJR3UtOZepYT+d9LW82FvvEfWIPcSMDrZyXyVvM9fX2wfw
3eMxR/d7jCWRXFfiZ4CigE0Km+mMPvFV9Be6W3UTUq40pyz3Ss1z0qskX8Nfx9vn
NGefzPqajB43N1dJTHznolkg2opX1dAgqmqHNZWInbUtGyUWnN55gAjhYQOt0zRi
QG3/Khhq3V6kzRKdYcdyfdd2rmN6RYsKfBNR3pjQFqXM8XJ0VzDtuIvmLELL/hpK
rEJknByXvaQ+6wSo9L//HpbxGxTTpgFoGdWO1JyHW2TtXeYog2FeJcvLpA+tewmz
Jtj56TRzWA+v1eVk724t7WONr1Yf6/ZuBkuocLFJzaG9p11E3XCZkJpcDBOqTGm6
lkewl+ClpduDCH3KxTUCvGZVxKAVJJQwoGFY17cYwF/B49ay6h0KHjg8TI+x1KUu
kTVuaojFQq1LaCLymmEVz1PeOV02/k5Te1rTn2naJD7aiVubg775YoXodWqF4dpJ
zx2X5vutCQnQV1UPlMtmzL63JPh3sMy0SWHoackrXSL3pitlnd73bjQCgeeVMSCz
X/TVa3NZ4+u8pGxzQ+ozJAdaSY/ELcvcZjuvXt6bLg/Gd23ce+Uuzk/UavWHXmP0
gsEvDOVJE8IqDdyPiLv4Cofb+BbMq+BazAfKHLnDkaBVe7/jDFILrgAqzE9Aq+S8
XBUlVmEaa52plV9tNIA9muiZdos6Tx1avkfhBNjcMeQzv7UKO1vZyLCqSKk9cAMR
41qAMIdwFt8rgsL5K/JEJaT3MOx18JsGmIxUKwxK7rlVofur4tvAKqbPMKI4HFc3
bRDCubtEjuMw0Wg6xQgI9uRW7CNkDIdwqQQzfvzWCrvTvSPTfyX+LoJrNzwwIK8V
S9Jqmt25HdWWj5qQbUUCRYr/h7J+cvhSYYXQwE5kW9TsRdFg0fGv8vY+n76lhN5b
M4ZmoMJx060hLfe/zNksv6etd0//wwcOYx7sxdQlnaooo8D2nysoVjjMqdSblTAO
8tZN+P/dewKi2DdrG2q9/TIh1XPcOiUtr53DEV331VjOHzWDTsBgRJDKybAUBtYE
el0jKOAIEIfJHC1uAhr+ifot1Ugog0Fee9MqXgetGFI7Qywrb0lcH2AD52hUqTfh
icBO6YSREca7DHHERsw+yxkCmLVZpeCc0YYsrJm7dl+w7w5aHCzM1TyCbOWTLvk9
CzvrSYxOLLfPW0qa9jcHqpmLvb8pH3sC9uRYBm/QVTC9ZQZpoGomxuH+kj5NWCeX
W4bNf064VbPBOSR+/dShs/Hb/2tcOyQY/1JjAXzf4Z3uRmbaN+mWveJYgIKXkOJt
Qlu6CNBRE8ozeTwHgl6VRqCV3wW9mKzet/a3yBrNTBKXC63W+nW7KclHdTZP8sXq
JTd/+ekCbEaGFi5dXL2RUr92EUWpDdEkZMw6qf/aNZOAGFUCu3ZFQ/a9h8wOtw7q
t7J2mNbZioLeyvib0hmc2ItaaNOdiVeiD/op2AZMOA8p86wOXuz34bfglOyBevE0
/n4IhuVISsV6hxkQjyGAIxF6SaaP4GPHIE4lF6j6rBtb3QQN6Zjo8Lqywact/bMV
FyzP8PEbaUfLG3M2M+dUNfWzrr+0qaW7AdbQOM0V2BN4hyXQ2/bHmtEfGj5874bl
DfvrStoKunhG09ZY1SWYtHj9nI7eiMVj3++ToEIsPNajEMLq5HCT+Zzpgh2zJcRR
pSZ0hol5j9oKxanjICgRCQUTz0zTCnauFKCC2B1jjohrTGrs7KCaRfzD2UTqtYM1
+POWxj3ZwOOYr8z8QiCsZG4JLDm2mFMp8N0l4a93mbxGje+mFpim7VeXqpZgzlwo
sXjGThNV+0VFZqpHELANl3boJBCdwb+7WxF3OD0kHMryAxo/biVNVxRsNqH4vDuf
6k2K6upf+gymQqP6CbBKG73d6IYZZjZ8gPr2je6i1zhNTXmhUw3f/AYLEUo70Lb2
uHeMEU02VXTDPjr9iRCAan0U/dz5bIWSGQmbqXS5nCw6ojTo3EoLBTBpcrwPMbCh
6L10nqkg/p1P5U5j6Zy7mxbUSJYLz2sIN5cmA74QIq+uYWBn0a4W87oLh2eaVO+h
NeaEZXjWsFgX2rkYZepI6hwI33uSmzDRGby5YCHZUhrWIAKFxcpywgSaUYbkwtNh
Hh5L57ttsc6BxS8MVf/xDV/z75UX6anHj981Oiz6v2Xq49MZVAI4jod+aail3lT9
uzPJSKOGY3v3qF+V/i6rLcm9V4Rhvr+2ZLYCnuBh0zhUZlY+rDGRhuy5IKMetGXy
ceFiIAevypSOSkH72iH+wdB6aVUTU/R6PelMul6dbqeqtJkFtFMrNFAEknRg/SDA
ZBlg4oxSyqV80pGjtf7g2xja28AYpCUrrRz3IudDXx8h+PFBo4HPvifNknO+8Fqj
W9mXLyV8b1Lku3CpWDNL+NlNk9jvQv5slM6beOUJb++RyKfau188rteQ0Lm21Zop
zTydp3TjUNwAPQEjWVdk636JVtr2c8k60lM22ZK+0JU6qmqPMFjTplI3dEKoBC2k
W1ZTbXiN4UebIxUoKESGjz/0NKiJqNPeteBKJbFcN29JH4GADDvbCMwZj1mxUhWo
1e6erqwjzgK2QhfRfYC9MqvQjTV3hMUg/HmA3wLfG0C4fkfGTpCJML316ydYz7yX
4gaAp/iuUExk8JxrJjYy218wvprSJALTgMNtcNOL5UyBuIp7IV3WzDOmgU5xGe9W
1+pXza8xDT5nlcN67XVsy9ezLUBGP0w839FQhhyei20BJydBb5vYRZewl4lgeWuC
SRGSAqnQvDJHIftPKqL82Ap9RPHgm1qR307+7wdMMaLSgPULA8BuMp3DQrqZBzQU
L+9XtO93KsnzXtqTD5pLhbxXcxEE0/rBGhrITV/75ftn6PL1Q4RCxF8mQ2aPlYsd
vjLQpyW3JTGQSaZjmlK7pg9SIdGbg4OEwsUJwtC7s9vb9pqOC4gxztT2ERb/3ilr
pdy2/AQPFT6uvo0tJcNSiMWGiMALDXVR5NjBw+KTjlXexG3QytB5jgJMGlAJSLJy
7V3mHdrYr0D14txsEDfkqOE1vIP65xj6pHTwIqPw75pVTsGnAVmrfkzlTAUG14ud
Rb6sh87omSXVSsbK6sWEutyzWTsH36ZB7An3NHoeSlZGV9fC9RUBhxmQ1OXKcrql
pvEwdDCBlM99ta56oxKpcLkMF5b79yYYHBgDFJ7cgk2M5ttRVPoVEbNSHtksRq4a
TycJlfQBIE5IdX3TuvXMvGOooloUnh11TxCCyJtwyrIQDq2MDL118a7WVWiUI/SN
mR/EdITPxW5PDmLDABAYz1+N65eFX/rvSTYqi1eb9GlaRPaYYP+5yJvLbHO7XwKN
9gSXKFY3keuLsM+yjF5niZLAydIpKAOtHsXEnnmVTYgS3xq2s5upumei1cStZjMr
Kw2TBgKkD3Qttt3Am6vXYvBVwodD3RvOr98SDIPxSHhOki0WSob8Wntp7FCpTh0z
Y2lM/Ui/0oEoyMrFN/pGW2ITrJiTPHry+sfaRrqJn7e2CPDUNv2LahGBm8CZeRdk
sySJ1+F30aAEGGOLIpo26UuRtHn/onBZDUTR65oTSd31ZmNKgAYuECUDMyKybQuc
mhljpdauIP/wc+CU0kQ97rWrqXZ/FnDSfwiUBj1H01mBlNcOJAsDBjYDuFJUEHk3
F8TXUUij2bEgtCnStYjZVj1clynsAcL3EDPl/CYmlWT64sTEdPbMhQC3Ws/nQbNR
DBRGpT93/u1hJpzirL/0jz3uDQYx0lgh4N/5mQIkASVJi9rx7l3zBhCmvpfa0ky6
zG3Rnk2Jeo91LnJHceRVQPXXzc3t6eHMxqU6wV/muVsl1WOH5VOoTJLuVlmI3lWj
OJuzfTvuYPu5PqaRbqOmwkVKMvva5U426AAfKUwoTL3N7VY6BZOB+tbEuNHCIu8X
D2gi+Aq1ujEiWoUkim7m1LSLKef2fLXp0xoi3NLikFu5cZeBKOoUnGlclJl71B6R
uQz+nrWWrVIep5oh6AVJlO80alcf65I+ZTaZOpcnDYL+NI0LE780TpUtMr8jr2+/
vbaDrOAdRQsjCFtr8jJdg13Qw2s6sTcp337KE9u2IWVJHHP5WJgtV7vXO+PQFyRC
0ixd0ozLMwHW6QIMzzJoeXBV4slmr1/gtYrZgNMP4s95nx7rIWlPkbwesposBgFi
mxFdCFbjCaUqylnSVIkq9ZStLSy6JHKR7Z7slzCZP0LIpu0NHIhLEVDmA1HCEFqS
nEMIgXlMuvcDz4XlZJAteW2Ewdm36dHm7AAJzx6UXwQvVrNvThfS0EcoQ/LqTd4/
3lg/GXLvlsfnxxkjfD0dJ7erOqjCjfN0JhCqpkgkyW7B2LdeG3Y5soBKgTIzN4X2
eR5Sypk0Bf2Zx1XEkN9PBJUBXe+jvFIExT1g7US0Gtdlaobt1znbaxwxZWwCrIl2
J4NlPMdCN3NehIfM/1RcBV1ngWqEFa/EfULpPmfSM43l1jupai7/a2GqqWaiI/tm
82O7jxzanooKpay3c80oEi0LG4OpH+eOe0O4XQZJDWJiBOpaW91ha5Yd/bk2enGo
xAQ4I/71m2Te5zvrueoFLc+GMLOE17GBzEnpFcdY0VTYeTnyDWDkhGVkcRCpxJEd
/qWbiE54wfaxaP9527h28led306jdF7KNs4s5uyKk7gG9Umpv4RTKYJHJ8qxUeDs
ZRxd5APrhROKNmSTuQJDIEFCcRUbourfxCwuoIGUWpRCCWmfys/6eHD5M9PZ9BG6
46/0aGoRa5xBhDRDUPYDH2QyzepAfTW83bM7t3jhdfJyGsB/el/4W8dROpQKvLyc
Igyat44T9IhkK4UJ3oVp4/KEoJEdX2UT17UCTgRa5H7kFLzGO9mVKaGfFCieyn1s
g2XmEyQ+xUCJqUO5HM4dTa+BCCN2Vdr0AjS/c+UD9Fi/Jj+AyXvfHUUv0r1mI5ZZ
yFOAmbQcmFbN73yvBoBHZj8ab0CUQieMu2wQBbGCy3R4O9lJ56cF2J+jsXqsJ/uc
WGCMMdT7O9nD0h5VvaeUu1Qj406AnQpgr6j2cyHwehyKV4xNUX5wD+M2Jlsylc4+
1k4Ng2Y9Nx135yDxgDfg/CyCn4CUScpG903aq4kfReKHLXPxSZvMCu7TNdTbVyW6
/a1feGSff4ypQxfM+TvFKPttRGWFpE47EaBgxZIVW18qKB+cm1W8cjwcc+kaDUlq
G6WkGQ3zCpBlE4k4VWjmC+NPqvnZCMPfrbPeLonuRIZnCBKZi1sky/1gIH0ldcp3
ww7S508Iv6q1Umr1OXqy9L+ZS7YNiUiAdXWC//KNWyrdjK2TM+QISdWR9tYKaZ3B
kRRkYuSbcT+g5AzBqsXBGNR75Zg2HmZkEfgvUSxgPB4UuoRH79FUpPbM1P4LfpN4
z5USaoEgxIL8QGY2DBJb8dBS5KqsG8LXlUdfoEbhePei1fK0N9Gokt1Jz6IwOh74
aK58Y7hM2QOMlcw6OqM6oEsZrSLMSJKzZ9ZFd+7z22wxA7JB6pV3uMY4ZOEeGCHR
/dOQ4L8Ite+CcBsgurmNKqC5Wh9146RD3KH8yGu0Sy+ZSvss1jqbMjbUZCsyLrWj
6u78kZWs/JPe0eAA1vLXUuDG26sHlfYfQX5K8B6aGcwwetjQfKgjeg3UZ0W+PkIv
f9Yc9gDAkEnJdct//popbwrVScq7VkdXQSAlvUcDqNz5DCmVONuII6h5kyAfXocx
OupCm2O9yXQSYkTKU1UNhKekd45yvaXVp+x5qGY+lrfzgFvbmBLl321XsqUbYOvu
5OeruHOlCCOWvHF0GmJ3TQNl6b/ZTOqw0IC8VJWG3vVYvKkUQcnwuoBSuzJNMg6N
RKuL9sTBOMJdrY+6ZPzexT7EIh4CiV2NOKJ0lkfiuUnOn1IMxQfPYv20vl2+oYez
XeiBHEoVnQ9mq4d7KgSUvIgD/SDHDquEGY3Wznef2SJlZPSnRZ2okkeciPFFmG4U
AbLG1aFQDbH+bGf42unOw48FhS9QEtX09mVNbW9nctkGo4QsyBFaeFYglJ19ahm/
Ony6sYI2KvdVvXzdZTVcT6pMUdiB5k1laaRxTqVhi3EKc1A/qdIGeoOezPrgYSu2
vLvH9j4yZ4NiSXPHPoVHd5v7BDWBMOEkVh9vmWnpcz2PLzPFgWBC8fDMpS3mxyB+
uhRsDohjqmUu2igzfa4b5NAAX/iHQPoeXf462XmK1K4uM9wWt91sDgMjQWXmLokg
cnQewkyT9b+8DFP+MhfQGCq0p6RfkWZDO9l5qO4BC61Ns0dJIuFfQ7U55zKe/auW
rZQ8zBPOtFfepW7bnscRDspFtGUkDRvDOUwUOfh7N+gAM6AXMe3aFKD2/+cgmBjl
NnebDOTW0fG69ducksW9KoWRtrKs5UoG0wbfVYQ+RNu3CNgIGTaYJl9JqM+pI9u7
tYATq4QmtSPuYQsnCM/o+8dMH82v3yBYuXpslPZnqRPPwJAAIFSSXynsOi5cjMmy
O+PK2Z4wfcGWyBGgesjp5XpXKojBP16jxIAqi9OxrDzFT6oKHYndqdUKLriqpopz
HXOINHM8jxJclsMTZ9OFA3IQvlx9A4Kfu4AyvqDADZ5WeHUj1THwHK5zG/e8SKpT
7IhNmp/RmiunW4+E0n+4fN0hCu/ZRvnTzNeXFhsl3LUUHBMiZWUJFhK2qy5gScJh
doDyf+XQdt3oLRWL5qRqsQ9js3DXbV0Kv5khMo4PCpQduYG9ra+VjBOfs3SoZi4q
WAXRksvpbVhf6mXdfvGXqcyiCPsiiOfr6DnQULq273pjhbmbNNi9mSfXNas2H4tv
3myg0NpZHOCqdxGqih9Vpn/TvISEuPpuR+5Kyzcls6hXsyxdqlFeOt3VRaAhrnq/
9hAap00gGrMfPKGLGM+Ja9vDzaOip68HC1yzaz1cHkEtj2SOWZiFMw0b4hZ6WKel
xXQ0UgcIYWQ242+GCzzBz2PXGA2q7PZz7FRiCjUyXPYdH3zKwVImZlpcOSv8v+45
dTeh2ub+bXdTomt2A0RvuE8wuLOhFV5EIds1mO90vWkAvMEOaFsc89orrCA1QHJS
6RH9EnxB9soJb/g07uT1VHwvBA0jYNSAD1whg/lwIC+Dizda3IqTqwvgpe0qvpvs
jdJTk0TtPXwS9TedYDbrHkW5hvdn812M/DWUMFBWSM92tIM9w0DL8PxQ8BxTrpEb
9b9H7oZi60YfA6ibNhuULw0nZbYqHYkMWAnCE0MvjxZDhjvC1rU39e5GCXjf1Dt/
whustSQp+p775qsY6wR+HISVNw5ZyWj5L6IdjUOxrFRQfgeo0/PQTYufZVKjdvY1
MmEJztLzzae55lU8jhlNJpPgu7jzLjZpK+8xp/XCW99H7gynJyqrsS6gkZhdR8NQ
EhUNAWtio3rHtU3X/hgVuzo64hyGOBLXik0w3TpuKUoRThijxEHbI6KU9LslPDOL
Sd+0Z8iiZGlLQn9yPudnOFC24OLCN+Jh8Xqge6dzClJ8UZKjNcTNFvXCF/h7wbDC
W1mwHoNVuxAmciqm8N+aoCMGj+nt9e14mkOOQIqtVueoDIvzPU+A2Dd/XbvwD75x
tgGTKjjsLVPYxh674D+ha45zS2mq0jAK/SafrjuzLY0QMoNjehqTFbaBSqUE8AuY
ycqoAqHnBzBxzCx//eaIXSPEu1tahClkU1ANMRV4RRdpXAa7d/UuvfhQl69qs3Tz
clsxUxEeV4IALi+wOdOTLvZ2ZlCbCaJwg+OUV8ISmv5jkI+dpUC+G4cnSiVr1Bxg
f5IulfWOBRBPAs8gBYcHwa9QCFbbKtfH8tATkSKBuxaOr68t6AXkaly41qu/L7CN
b/fCYg3tZa+XaIHiLZNbJKE+8Ygn2W3ZVbdkt0znIqX3B63q27n6rbbaXG8h79Z+
SuqvftU+BSGJ7kIgg/2lJWScM7wmxsen/2CBNF7+tsB7O5QTdjx1fiHK0Mm8Q9DW
xSdnvxtQ4SA5ubqhCSPsCzGehw1PO67KXJtWFwc3w25jMxrsZnXXAbN//6J75yoT
XDR9ApE+NqnkmPbyxwgHf90yLeQAu6IvUw5kz+b0AQo1ovE4yz9IMuiwlG+Ctda3
LByvqk9bAXn6LVrJ4MDlTuZ62kLu/xEiz4T3MerBJcCuVOXaaaJNlxudrJiIcIhb
dxqIpdQPRcaGlypJD3egdvpuiAz0q61jaFTuGWACPXhNNEn62w1Re7LDlmSYNp1f
cDtNt2spJrAOSSFSeJwQrKOsHE05D/miRncRbRGUUwME/5ehyhd8aatippH2KKiX
VwOKXazYMoCHZVgbYMlS5g3fErU2JFmOQzeMZzdt4EloV6UuPXkdTP0hJAdqiuC5
v8cBOd52MATTGS2VrtJVlsgHTMYoqE5DTBdo9c85M6XG8iF7JPnJSohz3hQRFvwO
zWiGEhbE4pB5JhcnbbXQv6LmFl0UfA99pg3/zaBDLmCK45QlSiXsjNf/rGjEU6oV
yzrT2b8BN2nUg0AxrsfEFP4l/NmDAOzXfHAKwiHPiXrCIPUeFZ6C8idxAmAoXACD
SQoRnltOOzvoLcMVyqZMGVoqetJHtYQ1yOnE+WAh5mQu5Zd3w7RQ6D71FgzyrWEN
dClyZ2YFiP/cUB0Mt+q90+1o96/c1qoy4Jsp5QsFtXUdlyjA1eR6tdTRXjbe15gJ
NhXoh5PDkmrL44QrEgGy6BM3Ca7L/Jw+IFd5bXjsskJDMlUguQroY1XCnLDxfk6M
pol+q1elfKS9pL/+9DGh9339R3mLitqH0S/++wwTyXBw1UYQiUJO4pGDs8l/d4bf
CAN1YdpqqbLDszSIcUHgYWcmwV1ZP2aoE/0KsAHhEiN8E/tSHwbGhfU/hfV5P4lF
mksAmVK0+yjplUnSdAZVhjbhmBmmAGD/WMGsn7/F0tLE47HqUCCg2jdtIkU3vfMi
KjXWhkZ0zaGxNqdAWqa+nkp91rX/o0I9zmmeCH9qvBGS0mC8EfezcSdknfVVLY4J
lc9qw6h2K3AHfrL66RbRB4H9vdDoMrtWunfB2MHukwkaF9LjdYSGQ8AGXc1P1zEk
62SUqzfNAH5MPd2okCSC/Vf5BVv4Ryo94wzNFIhGB+syjIDGayOy1eQF6L3USSa8
RNYl7YLoSWvjAb/MjqwZqTwqZ9LIC0agz3aMizjXY18oaJ6Sn3H8RM53jT8v7kRK
QvFj0smj5BzoSm8a9cyyvpyoi/eb/J7E/ZhAvGSXprQx22KnHH4+5SprLgd0BQ4C
Bo9hTny8KCYX4LJHraPKuugSx/mN+VkGMZFatCY+sYteV78ORbjrWwJqGtVvd6rn
McJz7t1VskhD6u62FW1DK5PRR7zj7GhV9X9NuiqscWTy1cCTeoWsdOoefRNZKQ7M
VOWck4ThMiMSVzDzK7yfnuMPyatLI2KpomvNQ8GE+kMKZcPLGgY2IA5gtM4ASp3M
9Ubtn2t1fcdzsOxGNHY/CYLnQe3hVSTJLREDYqOMINhmkl0otlG1lL5aAG6VR0eI
dMNPJduRStFg/Dr52gXoQaJPRX8EsCSQKWV5caqo17jpDn0+SQf+QWOuZp13WeG6
ydpqIAbakrHJx7lCWxEco+jrJfS1smVJiYthknBCxJymJzesTKAaT5Hu07+t2IY7
+9GHnq/0mvuGkMt8gEdF5RrwCgEUfipc0D3oqAyobFPoSfFI+WRO4QtPKpRWOC1i
gXIeIhwZbQKmynIcqif8VI+Bmob23AMOW2uQh8ZOqnNCyP+9UEUT8dGXP9oYIx8W
L7wedtxAWaEBpZUkCrzYtoYIYiLgMr1F35hlrUIgbP9+uWjAimLKS9cESLZS8agS
XmBIyrcxAVXoK37pDKACgzMdxoHSYIRu1TNM988bznVWV1BwYsnQFiU4LyEwLfu3
En82sMc9f0yGjJZVqhg8gSgvefRWV1f97iMTcaBJEvV2rMFZ47LFiybdq8lIDAux
6bjxS/2wwkhY1yIl1rFXn/EnrgMb8MpdnjBqI1oBZ8vioUNP2wGaIEXnhysHmeVn
DQXN9lIhpcKPF039BCzYhYDcxOtQJ2KySNaQOO9dZPsf8uBISwQALIxzzjiOeRI2
3vKdBQhUukmn8LQq4gxALZa5VksknqKyzzyURDm1CngCqoWCXbJy29E314DKZVMJ
HG8SzgxCB0MwPDzss0Z2AtTS1HmJMSMEXsmZi7njDhLAgaHauAqdyhs39ju5h1o7
EgnQHGQsHMcTSbh7PFuFWSzgq4hRAJKROYW5D4Mp2Zs3VAY2/kN7GcG36TGGwH6k
HvrAsUp2jsp6MKgt6P75DCRXh/ZughPhrqarQOUjvg/DtVbIIrXSXzn8pkDoJjMQ
ibHG7JcZ0miaRLvvb5nzHoEtpFtPubGpdYjj7br6UFHlQBquzmyQhGD4V4+8JTq4
c3nvnzjiLXXMknCcfWgotvEO8XkxiYV/sj6d9tiJwUz5aWFGtrdRYD+YD8Pud4Ey
Y2oznBWXhuKhjqcov2vimKemNrXCOBmxDXsCAx9hOF/RTHmbSe6jnOr8gSd2JTv3
58dXKCM7lRtwQ1mjz8NfdaMstn5uBBaV20y8RsZN6Knxb3PoiIm4qCVqbbb6X8V2
gr4RIH4eTeRKOKvPkXYSdVEMDlk2bC19R26I5wgJ/XVa0uu1npQLEgIvbrEUmdP1
j1RQu/a5C/VpZB6f95RbDZBVojYpzVkhdu1tgLl1maFojtg9+Fr+r6ls9S8Dfqyy
JQaKr1knXuzGQmQ0CdBuq1uos2fbLtQyLKhsyjJAM3PSAcIuMlRRJu2cNQM6e5yY
5vW0e4SWHhtdzTouC9j5M08n+twrdSTKkdT+0xwZUPDWNVUhpy43cDM0svxLbMv3
uT2kxWtcBmlj+FRurJU3fGhh4JC3kfoosunTHdfY82lgkj6BTm4fS1HvY6McCw0F
RJau/isgBlDRHvcjbVxopX9mWExkYSiiZ0GahqX8jTuveFrK/SNBxsRvTrFu1b/b
+6nCC445znzIX/Vbri32zODii8SKBqNyDlyiIzi8lbcW3p0LoHmUyaa7fi3coHhp
+NThZV70tf+LoMKJPiKqlcp3be4RbaOe3gftFvNVeWmKvmjA/+q9U7pRYled0OUF
KMZTDlLXLX14fLl8jA0Iq6C8gqrCyt15P1EGJXVNBUjx67E/D5NlMyHpgR5NwyQ5
LpurOzU+fZv7SG1SlTzvzk0fUxkUep0JDMmsSKGAEjvVft3eQya4uKUga8wPx1Cd
WAeCi5X89L+9ICkPhfqDNOYLM6bVVou8ont9c6NGSLadQK6pmFtAsAJJ7DC8cvnp
LEmBRiHHC6qk+iP+3lufXjKzgc0/lbm9NObda6yMs6E8amHhgvzXinUKu3Ubm2hE
qmtm4NItbnWOKJ7foK6u/ySxj05G5psoo0cJN/t7e35CnJSFxiAMxue/lHZIYRAN
4lUpPWFlJm29oJMGzUCNPYZxmZF9pIkpEWh7cSp+gxAkGRn2Zk8C6BL9HWz/IpRx
pUSms3kyggBZ6aJ5XV2wEtACNNxfo4SOCekm9QZeX/cg9wmjtyTaNTHZ8pQEC+7P
aakkXn8gyAex208WhEvv7KlwWhNy2Vco98PUAau4xBcpYit+PdvuBdXNJ93UxGfY
3m3hByq0m3eXqfR2us2EFX5Z+VrGhwkkUnXdK4pEz3FlQnu9QhU49YUTwYAsFUVy
D/hByztf3Vh3Cra9hafAxpTBjtZDbJvrUFxEyON0OHO4ejfBDSJ9L6Ee2/4R3v8Y
23OB2TG1osrCFSW8odJKT8dRNMv9SkEQoXOC1ZGX+5GNlt82rsUOaQhZMpmzgyuK
qugHZtpTB5E8ucdTnhdSKnlFECOEZf3y2/nZGJ8b9RidQ1UphpbPwYjXj6YRYht/
ApeEUBZP6tAS+0uYRPcNsFUqRSyRaUqRKCtsBTuP2MP2BjLEYgOpkYl/VmBONUO6
AZNjhUV8n4fISY5alS1HXXHhTkOyKjIvVIcpwaE8G7zBk/o8KP5jrCMvhs+7Kxwd
XkrssIj60n/kjpnPEFFnGgq3eSWyTMeKaXXiIv0IHXOYmKWWeIH+hZeg8NjBwq2f
guN4qnCX14xGCCwMdQu47dp1lI9SYsaHd2l2TwHvC8GYjH/LOEl+ZXG4x9RECTL8
0h9KYBe4BD0Mku66WOw0Wj1t6xT9bxG1xwplExuC7Y808KzRlAh6qSAGWGiZJRZo
rdM1lW64KL4HoL+itp1ZYjw6jcCG03FndScrI7GBMHMXosfnplOCGSEbVRTABO9J
GZxJ5fSImc0HE6T9YaAkXA+yLqQgibApBnrSgFdPxCNmIwJ85eU64xLrJ2Iwbpm1
bv8o3cAiCl5mT6RAgDyT8wG/aYA9U9l1ZOHzH5oHoqHNcbm5tmeBzOOPu5fKRNmZ
CV/wuSVN4TSorYuM2Hih2IgAlZvNemkVF5IANLpaQUkhWzBY9ip1O6asikIPbW1q
WeK1hY38Y6iycv4TynhTcduaVUsJcSA0Dna+0gYoWjSGEIFWopITFgH1nfGoZwnA
zcviTc4/tLJjqkY8f1nAohDJW7twUd4sAFW+5fZGUqK4o+5eybXejlQBDqsKhlwR
zO5BlxGCViJsUjURvn658lay9KOv3A+aJIVlJP9T7Teji8/kcm/7t3JKgA1k6D4v
kqhwYYRoPD1YYGmvkS66J1c/Z/R7XPbJLb6NgqgVT4cM2ZMKRFQMRNVSo4AJ9rBj
g37UiPe2irhYqX/fKxVX30lYLeDp+FVduCBHSvXogIlEOCK3kPTrptkIBU2M/inS
IGI9aX0rzIZfq7s5mTpmnCu/NhtwLoYJylkxnbNQAjs3Exkl0RQVSfMTYsNpyk+c
o3IZh2AmvUbXvIUKix/2lQSLIfZFnYBAho+z3wgTfzYEDEyVZrAQogVG8skRb2Sp
gKpnhvUUe/jIKrEodnXovxu1J0nDCzT+nJayNN1101tiWdUxI6BU2zuK6uv8tNK9
Ge4itbMkbml7w+48Q4PFTvMMXaLPuBBIeCmFAfEFKVT5pTnKSwHlGnDAOZBVpwjw
LGRuEk/rM0LdY7XUbrfqUgADzQ028rMePOhQ8Pu6YxbkoSePTsuQ6z/fF4s2Lq/w
6Hyl4g4wG5rUpNV+v7ExwtOo4uMZutqZE4L77hlqWGhSlqiFhoDRnEWM2YhFDKNc
PWBkBA13o9zIwKpve/tSIG6K5E5o/KaYAdnjVZ82mDOVJNUUovsxKfkQlemXVD9S
jWmsmn11MzI3Bp4AB1RR7wwKJ/YTCcQv9sQxCqu6uCPf1qdo0l5Uaum5UL9IOSrP
8x1DrEhfVVsFVJ9kVQDLpt91DokUUCr8XHNGkdUWzqsomRXPl5NGrPKobs5qhiV4
pJ4sIeHqDURov3o0AAU7u+xiPjXRPbFucXvVOfLhpH0bzI4ucPKmEHYWuG0NybU2
cYVtjUzu9xbIkEH7Eut+GvmASfn7el9a9YmUDuvWDbXirFSdAmqvpBVYzxRd1jau
fnxASa7aS9ZtwAk1Bp0htcG8vgPUK1b2xP6rZ4xgXK42E3eEM3ghZOJgbiIFbA0s
9PxKgzSQcPj9kKsjXTvqEB5HYKApsSIbPdsXBmKug+daSQlkiCm5qmIJba78pNKz
nAvAL/X7g+T+A+qMtYaqK1d2c8Zc+akfguo6dnzz4GWSFy0hJQdd0xnVxgRH0xub
fjODq7NO0hHZwlj7fbMm7V329zWGZF5UTt0BELPtmC7HwJnhBn9QT8ThDJTt9bab
nAU6tnaDaETKaxtdm/Vl7NpzeT1oacPc0cr4cYLKnzPkteaZMfHavHuOrQ6LZTvz
jyB0lCfD8jHatYyozFol86mSIRT73glnumswJ0mFYZVz+uw3zZRbTIsLlYvs0Cuv
v5RQ8AlAjYrZyjzn0Y9K9EGMzk1/c9fKNwv/4Z3GPMDLDIpsRVXmjTtp10M9pU1S
XFPZ7b7/Vmr/B6qvMABM/c6FRoIvnJDiDNu4xPQPbzkAxQWhOdlTpN3oG9n4a1kz
x8upifE8OuAD0tPOdAnn20ccVHR/duIz03vGSCuGrHbEeQb0O6V8XHG22rEwDQHu
ojwWD1wpiF7WLXhJ3DS9Gq3H+7AvrJK8f0Qro8wGoq0WWckVXfOcd3kg17IHZpTR
Z6XPMHfGyCEkdXJuGhYOCK2NnXlhbVBHJqCDS4EJ3cvh+t9LeSmmIHgejNhepIS3
kU/pLanQkLqbX3fcP95VK7J2gU810xHMnCueAJmSt9ZMUqxyVMdQ9czZD99qZv1M
OAqwkpvYZW5pmEJND8qyvti5mTz/eS/n04voZH7ce194guBTKNF5V8twMiXHlVlG
tR33BVzEFI3jjUq0+KnxVvFF5/hIK4X4661hSK+279ngg6dNgIKZje9wh3wynPSw
M5bsigh56QiwLCsvh2j3L1/43R29/ZhZ6tw1pBHEDDVspvaQrI1JOWFK60Bc9hqY
LhtCFMVJ7Pt6UGoPVsk6htfD5i1WxJTBJIbjW1t6L8owIrGJX2UoJoTS9tmkef1t
5A3CEiRqHg4AFNN3e4Y+AWNdch/JkzAZsE/NSPHU3DogJzYGNXt3z7hVUwggn08c
qrt71Dwk99N+3p7vx8NU+r/GWpDQrM0XJdOK9LGr/AhL7VND6SuVSCeWTFaDZzN1
9rd+gRsPAliI4orO+5TQ4yVUurOWO2WSy5x2qa5w4vkCRWJ4yF9uoyBKimWpeJrh
71xFyVM8c1mjbHgGJif73LXszUi+y7Axe4ijA7cw5qYEhdfJ5Qr7kZ4L8D5okLf/
UZI0RnePYmKFlB/gJk5AZNSFHpsybMF7Mvo3F5KajNpmkgPdELCJIU9HmXCRoUl5
DGB0edms1yU0RTp5e/3n499Zw5aVfh0gsWSd5W0jBRpmCjug7hwOv174tA5L1Qzv
vmzQ7joO+cF4fTg81ULDMgCn38GMGUpvZ3twe1/hTFlvXcF9rAynm7oHoangXaMa
dtfSRrIxDrvDJIXOCCnfY5OWSY/UWHUWpy8fu1B173qT74kFET8mYi/gUonFmEw4
0ounvILXZQyfH4dPxRMMDQDja4HiYim2FJ8GdAPsDeeLs/y5jvNqQBMLRnwA9rtx
2f2tPcmrHDmx/4lDaG3CiaDPqTBqnDHDB12pk95BszybUQSuJ/S6/fDaJ1jO0/2l
WHu3lYc2teSx3VQqg9Lc4S5CwWhFAfBMiZC7CHoBlqypBrQ01KDMY0Ds26rMUt8y
ObUJWilwDrtHhX9Zqo0rNBT5eiZWJioz/L6RjzA04Y3Isqsd3DidtAL6ZafTM+c/
HZtPf+OAoqIWXoL1adjTRN1g4VJLpplrkfc/xMai/sY3eqH+aXOACIGED7UxZ/Gm
pJ2jzGEsyw39B5OT3jUDa1gFtxUfaLUxX6edG6Q1V81xaenzKcTtIClXF3KoKRzX
I0KkS0QvrkkvDevUlnrV7uXCKR+ZqGGacLKh5t+NRHcrT9FLHnmFGygs3BlArl2m
0dCszI6UGb+LC378BjxQPI/uO1MGEjm8CJrLxMD3+MAcmqjT2GA25BH19Td3L2Ez
FUI/OnA0LbJSxYLN8a4Gd+JKXjovo+WZMoz3I2rmDndjeebHxYJkzmevvrvp3J9m
VEHYt/k5KPzhNhcfiyVSUtfbLWrk0ey7uqJX2WlpvTKpm3w+W7s1ar4JpyVaaKnp
HQyaiPqI1Z/R3FKCCZU6ySdQgm/wt4+d1vB1KR58TNxwQnUaFpKVgG6j3xWLudF4
jeSogoeo25h5ZPiPgKFHzcr32PXqQBEvZbFY32P6VkRF6sjO+m8l9S5FED2pqR+g
4b1/purUt/V/J4ve6PBOb8BUCBcToin8FGNulZ1K4ZmE1f/wyvKa+sdjPIWzWgxq
44ZPUjlrMhOsKlFSKSZ2ckGKMz2fOKzjSrA4qy03zM21tghtO08oUVkCPSFXnMlu
kzPCAuxc0zRuHRyyhnAVkkw7FsY4JMKxUTUmJKRvHqq+FdOTQBOE/7hagsve96u9
ld91zx/sAR3Tk3XZ2X/f3lhLj9KrczcqGb5itXQpiayMAxvzmlywLY5c7YRFXpAq
27mrZD0kPFb/uAmaTGvpbVCr7Zeh/nTV8Jg19rvkvMlM5XnJQ/9QK4gHvyDnVE7B
vg2hHMrlM8nL1XTGxLyGCjfJdcfmvuOmq5f5QRk+StsothfkzxCLjqqxN6x2lHOu
RSifJFxijLIcBZ7hN4wHPu8UUAJOAwtYw5Nz0VxG1TSpv4eIJy4xNXvdAA+jyCe4
g23gDwwOX/17y6ohxc8pG/EZYtNQHONrlC4CaLgDHe3w3NKW3Z2D1Yu1rV0pi5yM
jdp4tS1WadFENJ2iIs1GKJWkhBg2YBaCsw3HZj0KFQnUFGjwELOtP80rLMMgnC2q
rJjYBcbXc/vfeJLFkqGjZAhVFJmAvaa8gEDwRn2/Lnh1ojHVfVjYGXcanDK96zn0
ofKe6+WVsdvED4K8coUL1GRUhw+9xGadD7UJgsjOLjGz7I3F41nTuKLyzd2qEGeh
b9xFcI13vssygM7YEHDZQap9mPnKzHOFbop63TqSX8a5arhBAEflHXm+869YxE14
uNLbWY9L+pUXOg9egLRPKYrSDzvcUFn/ObOtK2vwJ8Yb7S+oxZhpVkf0YU97op10
OOpVyIV7YKUHOFUVrJq0BUxT84Hm3NbKwFxhcAPRy5nU3tSSHTzutW4u1cJjXSTY
VzwucAZk/g3q3w9nwjlFh9KO8W2FUU3Xw/pS37/95nCHiWj6tAcw/5SZrKYiD6U7
q/lvaFWbcHDo34Ah37r6TKgQDHe5KBMh5vDZpCOG6e5zzOwNK8Cz5khJgunf873j
HgCXUTfrZy4sqb0JIfloVtl3ywxQFPAQfQ+Px3ZKCyIP7LZ1q/D8imfun5FycQze
SaLtMnu+ANsoZfCJhWKHW7JScYxqTN575DYlbumF0x0/DkfMmUo8TJ+H9iAyYKuH
XwMpizCo+PCG/xv+UdX3euVvyg0jzqjRdQmn30HX2sc1t+aV2SQMO+Yfw1nkCOao
ShuekC/Dujti8EI2hiwkcpGElK9vQNu/ioRiY6WAbc2RsJQp9vQ+b5ZbeO1YlqKx
ojoEwjvpxPsFzLqBndSEvaghOclg+Tg+fa1KDmxxNNmHmt2hnQRfi4wdUTR5fW1y
HY5/oQezNIgObOTrIAopQxwA9U5rUurBdrlHxgmYtJQJk74sKhA585AlnNy6eqnx
/gW23LEAKW+zHh/QkYjvNjHaykEiQHIqE5yYvRVSFTgh0B7g80D+4i1dbLfSKa1P
CLEhHm2tRQd+HeOH0abgiVz3fRLHXR6yiu/CzDvp1fgDb3eu5EHq9JzVL6Tesqsj
4+0yJF2TbdDbRXFsF19gvbm9ko7cTnHIaBO42MH4YCbEVya6ccWwTnNAz0msCUB8
RmPouNhsoXVTflwA6n9p4fcqK5bTpUUkumis2CSdYEbZHCsNXRj/Pe5mo5TafL7N
8N6ZxSe6I5V6vlZJogOX+1SOq+kXKgC428yX8l3avCFJPcbZZV46UiwciOTEfBWh
AJ9sSopJwTnneUVGxk4qnWxJ81CxSkxhYJD1xR09cb/agJDbp1dgHfTQpDK4MVcV
H1SDj1ezrnZm+GpTotr/3mTgU8wfpKagHhFtF1aY5rF+ZgasgRuPe5Xhlkaw8KIE
xKOl5GSaKJDU9ukXAlChHUCoJXlN2yM+blpCw0eVSwE9MI8pDLE72F5nNOkAu18P
Z4B3NT/iTzLdLc6lHYc9p/D+NMYZ4SKWy2+vFdkFG4ld4fJHdnNKlaY+5aYW2Zpr
gfFObaSjXLcR0+GtBnQ3CQJkGncPhfVhPB7kSSldvP1ROjOM5kLgU/MxK9Lr4mL/
5mHnFOQIsqV3ClMsBHE8cJZkzvPL16s0FIHkCQX4k/cMdMMmBz4jpOtIwbHYTtbT
0rdVMF75LrDF6jbaw0HdqcFSeqZJ4G89Rmu5b9IZioU5Kp8VotRm7h3cR/CqM3Um
rTv7xqBcmyTlH2BBlMelIG2DVrEXDe63VUZ8GVhYQiegLMPws+ELwWXBTX57O+As
rgjFgZdm55IZ4pLrCxg8cnxnJkIPlt4o1njFPyPJMrR6zd2HoXLyUuCGX0V6WzXP
wiWeuG6X1DYk1akjWugfYCnlw5U7RWrHJQ0fMh/76i/0rOrmXEEYf1pYleLE/goK
FqlGVNV5/j/SdDx9Ot8xEcax7yT6JieP4Nlk7NLKq6cpS/pw4xrqgu8x3P/WHBWw
auGQcseAUSHP1TFiIxcR6KoYP3/hjqjkl585h4d0NZ/dDHL0+8BIhbjkdIpdspz2
LWcXdF3/utK3vwTOEaLQvpERPp5UmwVLUedlIh32OsHnxbGdGHpEL9iyVAcDGxsn
ml/AhdBNph/7pFfndG559Ko4VXJLpZ8jyFgZb7NUsph1Jra34XaptIR2kBeJmFIw
RKlsSMH4exh7KwvV7wPV35/gjpkXCzyTO1lgu5vyMrjsn19cKapf6gHUv8JbFus/
hNBTJfoMjzlyNB82ttA7Tf0n96H21VWVsURhbpiACD6ArqDPfTFt9f9/9HUTdmZo
HxK3fHA88G+fkN8ezQlCMBp5+EZ4bV9BiepSTjqJoXOxY7CL4ieRL7YWheOOEmuH
Nv541XxLTFN4xSeVPtYu242j+lG9M6HjRdFglgv1zS2h5hqVwmnXFwXNLCPGo2YW
necvj6mYynt5hvWcOOLOgo0xmMRtVXXn9Y9wCWVRYHQiQW3npFjiIt6tdo6PewQo
3QM28gN1eSMLmNC5TJ45L1C7i/pf9c73WgT50ro1Kml6iYM1osDLEn6W+2LBfJiy
5Y1yAxINpevKqNRL6u2bHFBJlXf+I0b3Icb+N/VIoxBgLtsfQUqbBICFIfJi4H5j
kVxfZr/H6JJR8bfsxnj8Bu9VT528V5zLil7SXlIVaTHNocVzNiNH5QBovGTEEppD
TfrvXcNNeuX31/oo8AqKbi4RNRmMK1W9A7txfQv2vdI9KUlAab4Q4vhxPRoXmLIV
YQ2tzYpFdkV3rQqqmKi7yFKHAPtX8lK8bnflWoc23RNUaVmwW42QP8zi2UNaV4f8
kKH8yBx0vksvW5BVS7G+sKUEjSceNW++sWFNshZFZQusJqFYa+/nC0EIQu+/iy8W
1B9rxVkDlRPQOsbmPRMHMiuHa0sdpa9ii9hMuiuNVehbGjKCtYwPykHEqGA9RhyH
sHI/81bz4WQAheRsrCwS2aJ3I3Syg8YP/1GJiczGAZ4Fqjd3MhzLDldwYNukJqZB
W79dvewtzs/1jQaxTVOMOpHQ28vG33HyXp8am+0e0XoKfO/beMXBuPU2TDm6YKLA
vU5KiJiu6z54TY2V6t8Wgyh8THcLurU/WJgwaAEr0Ejp8I1kfgir7mCIkn6PoUO6
YKhn5YKTGrSe0qhzmGH6kOYaCVHAsE0ySktyIeZa6DarRljGyid7NBZae9TivYUS
7cEp53kQN9mEf2WwBVEZ5O+SYjdlrc34oeDziB2naNzTvTXRJH70tTukDBeG74Ba
F/47YXtTB/KmgWRYaCTZ45Sp3P/GJm0rFhttkZY9ri9UbN1e7aeTcVObhWyyXudA
mOJW71ITr2MCqZ94OqoPzuiC4uGGHY9+Sybieph6psXLAu+nbAdidYuJfqPg0DpM
itBQMBLBwj/32SFkFYm83mtV9a2A6qULFlS5adwBvGpXHBG+kRKNEXeFcXqsdL65
K1RB5XItW8nELcvMMb0+CsTWKGyyek57MqVzZNjYrECTtB3Lrd+s/uryetXiaxDV
3emz6PHBafACRO+vLk5Lj5HTE/MQ1zKWp1BJ5HnjZEOANNSFGRCG2JNsfHALbU3x
IM7w4okIR0r9amErz7gw6zqILpqay3R2ri2utqUCJLeKB3a2nQnXDUbOcFo+CbQx
cSNnx5O5uWxbAkLUQEsQIi77tHedKJhOVrnHorbHPVh1nfgcwAdiZBGzU2iPF1gO
fN1TAOGGti+RFnXBez/TKzo4heQgVrYghtM8wXWEM2F/C5MVmkTtZ+N/hLJfg8C3
NdMgPDSNbeYsKtowbOY7558lbcuGn5GbLBBjUVHoGEFZJlKZ3+U6Jfba/ZBAsThS
5lR41oFmLgztSp5dEx92hwA80J92R5IMEIdYDGrSfio8fLt63U1sgPIijJc7jady
i+brOhKGiS09a+fmmAxxroJoquwnGipsVxbeVgkkxYntZOpJF4sbJeTR2inVVt55
Ap5MAURrXUcXZXDL9RbnQjOSNYt58KZm0GJAUIwV4ktBtTl1HJsSn2DryKkKTe1R
Tgy/70fkXztiM3RK3w5RM8vExxC3O7ZmJORmzNd3h/nvrOqnDR7tcYJ64Ib71U9G
BbK4joYQTonx1hBYj5qsM0lBnCNnG+dAV0ZJMxDXY6i2hK2M7paPt3eOCgaD4SPG
fH/yE5Q/B1wcGCj50bsJmOnwvmSZEZx5SOzmzYOB9omXDZPTmMvrypQoTGk1bxc7
K9HFnLpvzgGSwCbteeMqCGLcUQuV4Ov+6hLg5GlsVYFXnp+zC5kt67+hl9nN13pL
h4DwVe/QZnTTA2cwGm74oFc1CTFrxGPzOzzj30HBmo7q6CODkzcV6OkWWHXXvWJM
CtlnQ1FeOQCtp6ZqNDO+dCOTepg+KwlGaIXBlAQNKH3tgJxYUfhg32JJxFIaacBx
OkB1FMblr/Qap7rkPLADba4GPdRxbD8po15RQrnQ0C0PCUfq2PBtM8oV86x3aljH
0fUqNjyiOKJjtMwWnJvklVPn8gfCtc4lABhbgNstsFLA43eqdK3VpInXF5QEtaMS
CLhRWYlwMnncDRt5Pj1Z5S+aH6OIe87MUYuqj/t8bbHlUg7PsMJlDKaJB2yLjD4u
QHD7zJXIsgxWToEgc87MBhYtVPltMFiCyj2wLIYWrzqO2/qrXyIxgPHYbyeSjxlj
PUXIIRm+E7WiUz+LURGl6L3npX+bSS0apRS6tcKBZEGxsOCH709aJOK/zkQr9ORh
PiVU2bM3nccMuiHf3BzjGApqa5inV655+1Wn8IuGcpq4MDeN9tfyX86T0e1J1737
6NEkVO4l2vmuua9gA4Zg1FNbbT/9nYjizef4KoNpvRZeP7bk4SgEiB2ZZ3uZnw4N
IKiZcnxXQZQzNe9mN2SG+/+2L68ZkINHUAUmxHqD2DxiGu3z/t/1rWjqfPAbTPx/
sDN4vcy7Ufvq/IKD3F6yT1sHBL84mrhmJCnhl/1biPktkHMDRDw146Ac2gYbe/g2
2XZe2BUgrrgMM6F64CBa756W2aQsBeJ45sdZPOhD1NtyQ83lvz96J+k+vdeZejMR
HgeQx7LeE7kRMDjYYNWNBrXe6NskJLIrIXf4R76bZ5Q+ZvQWBlKYyGsaVQOEeQ1E
tB18wRhlV7B7sbYyIakqu4VYBc6TfJkiVLcnZ53oi+ZyCaUAnmj+bZHyugH82TsP
Z0soxzrRb4/CPo/R9Udo4oww9f4/wSPleLT7CRqN0bDcuj/sIDtTvV4HX/lu7naz
1YGo6BVeUmz9UcVn8buOB9FKkzFB3Z5pEIelwcRG9fyCevfJ1NQYFi9PdEzrbwyy
XnOKZNf5k1AGIPYOXwUtLCqwkuDOB+Rnpv866JjV0U6KM+AvmmIekXlODGkySElW
5+AkoJgss2I3bEZIYSM1jhl6JMrNIauVqw0VUFq8QCWgnVeRVt7sz4p87mFUhJ0Y
qYIvVTcgS5Of4X7AIs++PTJVfRJ0Lj21n/pVgIaOHmjdBi5K1hGvE6KBorqfDZlo
xQsFM1CGXjaMVxo7l47m6GsoaKBVHuYMh9I6tb5lOdtZJ9571mGYIp4d04DpKPLP
FabxavqRNt133OC/JC0LipwQ29qq2KhUvPEaYK/QxBuKL1zXcS1pHjdfRIoxnD6R
qcqZCJLaXMoQUjJnDlvlETd9M+BU59bGgOe+6lkw8zigXs7DIUdg1gCmB8ZzJYQF
a64xDgc775GCxS/UgsPgLHX1p9l6acR13fB0ZxdTcAg5D0DUMEhNH6q2IkLQQpjz
bgmHGXL3Y3AVhf1hq1k+dDg9Y3cidZstzXn8yXz1YZK3ZBjajXpOwtcdYcVHMSa1
T63F8hNo9TnphwOz+EnUl0gxFjCWKQfVCN+woJJnN1xt3m9JdEre6UQ0nAZRkxrU
AbXXlwTEM5qnBEd1P8BQizkyv/wm4yIQofyEIgZYjPqn4AuQyJplQ4NU5vhpdVYp
0lrRauvf8ek3VMNefhWOhchnoTTorYipyvbwbLs+S3ezLyg6iIOw08ybjvceZwPb
Z4/ox+lDWRo5zBENuU0AU8XnOuj10Ci6nwB2O7c+WODGhbKIloKRWs+A6qP+sryo
WYe7C9osJ+i4hAaTVCt0+JPvzJWqLEjdtjx+xUy9//8axEhyoTVksRXVy/0dGmdB
GF6cfYb5YMMWqSx69Ycaprcr1iqsKxV0EdcA85HsL+/koC10g15onHZ1ZC+pRz7j
058mt6yLbo6f0LC9h1xV36s5pw2/ObCH3SGcrvpz78ptI+pVEtRhaGXRDKZcNkdm
fu1G5DyvxpAVLSEkZUOcrUkAUFY/LoBB5TP/rcec42v7KWmfgYyRxQEe2ZwIqEfK
xIWk8Mff7lVVgqLxAmw1rQ8KwMK+cx97RCKgoRRuNfc0Ok7EPtpm7jv127WVwmA/
rGUueZLymtbQSaYwOT5uIq1I6qe8CG88uotwLStx9xh41TUvG61UKApUDYGWAd4x
FG9IvqZSSVop1ep32CLSwlCNawgMtSnDBreSQuXuljfxjXEa6Ro6jHw4RUkvYUWg
TFjzZ/xjvX4zG/D8p7/lyiwlzM/GGPCaXhmxa2nNrTZZn6K551BHOFyxqeNy6sJZ
PSTxfqXzL6bUoh5KSabwk2oLsaMV+HuSrxSYwSc+vzTP0Z7oa8XGSG5jCFuJHPRr
e4QQRlxi+IwnrRQSekcZtWy42YEpO6OxoXIXrgpbI607lmHWdk7nY8uM9sh6CPfK
7nUi0FU4yDRK0RVx/FZiueqvQCudiGi2a7/QN54c2dfzwzqhl+UWC85zazhTQbE5
uMCyuDmgu43tN2bzL+VASBctkx1zh3OgmQvGbEInen0ACdUf7wMU6Xm96PwL1pzP
JifeVzXEnSFOf47qA2YYSzR5RGTc082naggpdroYzqAfcnF2uk67Io4eHVl3y9sx
RcbPO0bU833YtIfxPtU87/Zs2P6HIenauQ2V+UPo8+vUim3xgIrI7E3qA7yybf1f
n1JXNmmCGhVWHIesXhv1xMCkUyh+hnb3tnOZbJamE4JbYDhVxk9JhLY1dbAvRXo9
GZe+A/60tq8NY83EQNgpY1tUz5Odi9rjP3wFMAk/o9J1j6UVHOxGQCasfOYuCcVu
pGWDbcPh9tcZMp/3Mp7Zqk8764fAoHAH7MqfdYUKucDslUVXIzY1ScFke69uIW+G
ePF01dtlrBgWq0SkSQNBLcEBZd9b7ISyLxT13C6TZaQJ2onT2v38KjJtVlj/m5RS
mTiZxOEaLfdlRP9vPQuTw+Br+w0+1vBnRh+NalD5c/WU2rI8mv2He0qZOBJ0JJzY
yjXmE9zHN2vCpBjXoaG4EXWFE5LBzMS2fljMl1kjcenQsYxG7j4PN4IKqw1n8Jja
2P3dDvWEM9o5sKCovUYNLnWIkyqoAcTS/Gamu9/ujY5ILFjswpim0uOb6BhwBpkw
PdBaGWuVffh7/eFDH+x2mtKttXTb6aZ4eZ+O8G8TPWj/4t7UBF4E8+AywN+GyiVC
+sxLzHEF4oP+KNez+tHPHWdJFJ+9byrklWAK4QrxwHR2cPOCQp23kIna/lRJdC+4
Tk80sP7fxIj/nyyE8Qs8+yeMrAz5gz64soM2R34MwsGcU3nEYkKEPnzxxSCNNXz3
tn+NTeBkXclJ54D85DbPJ4N+fl0/1RNsq2HzdNuvt6yNlSC+IOs1OKObQQQempV9
g8g39/giboDo4LgnoXzGurQVNdPrNAQvFCp34ohTglHgB7RYLpqqX1ajeBP3rP6d
OLq7WON535Gz6fGKgEO9RxQnALWHUHQ1ZbooiEyBvX73TH6JjBi9ZHoE3Ch3nf5R
NRVOaCBZiOrkxqmx437K3Mn+KHz0ohmOx2MBoUYYlxaqzTjQFIgd4ZrJtTbpWrWv
MLGT64ZXimms4jmqCD9ZtYKob5C2hsux8o4Ro3Q/PEhoqmdFNobC8wShFfmgNlA2
LiSilQQ7nb/evGi4te4LwaruQ0jrHdQ739xdfMIhgEB2OiaXeJ0ZtcVahvwmpaKq
Q5P+hACJr3xgKHcrGditeBhUtm7z6D+wG8Y8+jbSPPbdkKQXFZLq2dSIWRXtHaTq
ym7oeiMs2rJYeooU1CSwyXW4dCOLtyU/XuowrM9MbMOOZYDfexFiBG9S5lY1t1pj
KdILs6QWVN56rilcNEA7K79xrApLuEwuUC0KRkGqfgq4jnA2OC8QhwcBcSptJaP1
D8OpmIWUkxGuBCnu+7LknUPcmrrA+aj1JDL3koRonnT6G/Qga2br+j7E5psg8kTz
bnX/3Z/JSvoiGsLCa8eRC33j2VJavtaHXfTZj1CXidsWImqxuPyTActYyj8+Ey2Z
Bl0HKYd7Bvx9DtCmwtk0dTA3+mAJQpwVmAV4WizPuSx5s4NAE8l366GRsS8pShjf
tne7M6+6ibrRQ4lo5cmyPQPzKDan6ffdtR7DUZINs3cdrEGQ9mbwQMZr3Lfn89h4
4iPSrteUPxNChpvrIQxANHH4iV02I97IW6QZ7YUyOKFhceIHbvYA3/IpLWzEZ6sO
jIfhEC3bnD/zjvE3XJTpAlr7C2ywjK/UXJwuaVcyaHxGLC+95ZB3UFqkV5hnlFjC
Ls43+k0FkTrDH3r0ih8Wp/ZCfpaBgp8KFR9cTfoIs+G/io35fvO4jLBu4NrThx9H
PCAJoq7ToDa5/LCJCExGio7FxBsuU0+jgWBSXpEkBn8qsr0xuwsUWInZdcoE7sjf
SDgKgh6nY0P+xV2TcpN1NOwTl8f2KIGIBw4HY1QNKdZBrr/ApNbn7eN45VRzKwqN
cPeJqKSNcWeEWoig/zl4YnwsTmzl/h92j5grIYAoJfbX0R+/2mt878t8Oav5ltBc
nqFtYMD+FuErmSlDXJcHpzbiMh2+kvcXwhQ1UECJJwwme9kEPqjr5jNwuGgxRgX2
bc3VBpUCt/as3I8oPRtUSGy1v8wGm78B5phrlJpd5RoB5F+f+jQFBD6mTwG7V1ck
e6T08nJqoorV7GAl0zzT+75dwWWcoeOXrUQqzE/W3qaRYda28tX4MN/04x471Fmw
h1T40ydqZ0peuaaY7CmvjLwAcaxUzFBSELQ2hpsuGof+a7TL5N1tiwfSr1r4gOUN
kFPmRrxI6h2O1OKVXibdTaOxfDVKCPDH9qUhoDEmOSUaVMXc+ChEmhq68tDtm1Zv
anjvUp4hgAkZDanZRzTGZNwYoA+K2Mo8RFxrTp45X5Go2kfLpvUqN7oiG8aW26qo
yPJPqlvHzCDW/D8dCAIczJ8UnLaHwB9DJ+Dv4AiYLtllTYeI2E0MXrZR/APzcjNP
4qJ99X5VZiaRkIVrkVCzT6jfL6mkG79eOGeAcSNNgNCpq0jUT2Z9xnTtTV/Gp6QT
35H8q+CmUEkKPiTMXoYAuPIe1CMwgfd7CbNLrOYyBT+GgIrdqkPmH7M9Vrc+KfTx
ZPtagWfm5srFiwT/q4X6hPMlal5/eM4ulPu3V7aTuBjORCnQ95+RBWJzssHj3+Ky
czEYNvn7XzjCdfIv8yQ8in804hLQKFaJ/Ds2sx1841/cFMinZ5f9hZUie8zb81io
WGvvUURqYeA6W51SEbwchMUje0DZcsw/bMjMI7U8Hd5BQC++9wVEjj+DEZ3bTpGo
lUWKPpYqY/85b79/HxY/bN7HfUxLv+ahGHN9sM7Ro1rjzuPEdxgH3p6dkETnE9FJ
si9WAM/J6bGoXkv335dRuibJOkiHRH3czA6zVzhviLZr7flrJZUHLPPLB2rAkKQA
S10BcqewR8OQUIfTyYmh8cbuYbG4SsvXPWCPwK2PntDknVg2IQ2QNCJu+9VkDXEG
S/d8T0An8CeGtGQwcA1Y/niqcEGrikCuYyox9bleY6I0KqyPBpwpUDuOiC6Rc5xO
0mgCJ8hfy06GcNmV51PeqhO03sImnebPFn0qtcoB9MSrQsh/z6BBXXwKXYHy5OMZ
Nn8k/hQoGOM1KoQQQSHqvmANL24NpQNIZFhjds9Vt1fe7OVaRqtsQjn7tmPLtZPY
pTV8nOnSd+IQOFuqsWin95mwrosJy+pLqOq6qROWcgMcjxSEqUswOdIKgekESn6D
hZSDH6EgXJU8EVbAH1QAb4Tolq4lk32TvqftPqwMI9LOr6a5N9ff7mp8SwkMQ+9F
FMplYNtx6tJqaSHHhYwrW1EPoiMeXBDSVCxCc+AMsL4W0KyhClDay2Exu7qA4Yo4
rWlb3p++ZwfyklnvG83Mapm9n4nV75K0y6NwVcSW6PKzRUxTwSSnEdkJB6vZRHDb
NfGLbx0LiGbq8GEgpDR9itZa5zj7fa5WlT0diiY1CYbfxYgV85WWvn9Mc/JnqFqy
HhG9iONiQW1FIlThWLW0N5w+qHdAZNaOfl1NRWwgU18p0kb/UkeRbG+USo0AzQRx
OgwJdexhpfJFpfVeta6pOazTNN5ivehMsnq9fiIyeTY0JBuN3viVoF77PrDsaGDl
aVFC06U3PkN+P+2uBcKQJIKDTLzzyxPEJYjgEKTrS1v4G1UOFFuXQ6izaStWK6T4
jdqSroiTWgAUUu0cr/NMdfgTsdG/DqUa2n1yyUNYu2j+mO/mStG4E+xcHGb/p1mC
wfOE6f78ptBNpvUEucpLQ60bfxUPhkbMQf+GyXiM4u4WGXTTxg4UY70ZmmYDwUeE
68FQsLqQ3Q4NlVEciT3+/6/TW7eFtFbhPzCX31i290PyeFWhe2zh3/jkQf+fVh5G
WPIeuFxa7MKy8qZCy5iuq3/mnjDbm9cG+05T4U6ZZKU0eC7Vo/1C3eaPUghBkvNw
ydGWHmCYD99piv/wuTQqUuku/CPKFxhNRlqg2L5twxnd0pBGRkWJgWxpQxyTSnJB
tZuvo0ANUPavXd3Z3kJfWL9jt4VKYYgBweXrPNWUzQskit1Qdw+EN6x7bNVQr1Re
EebdNLppiDmmoWVmorSgnZk/vtiw9wikExMYXZB70jYcK3KXlSeiUH4lcUKPbJJy
6CebBL23U06GxOSIFjBpHESDelLMjyFJzqcw8rNWWZOtz2pWbzC/YEi4TXFXnvYR
AWGdu3rNeQzHWMgDUYFQ9eZtGgzi+mGvooKREKPOIgCZ5P7aqrotuNzR4a3V3HpN
272ZUxZkTGD+y3qWADRUt0yMlZyOfgCtZAoaBFHWZmhGqS6ztmlDuQ4TYcduH4Zb
xAMYLHSpAVpJ/alBijErfiSvMSdfrkejdAiVJEVgJmn4exPBSWenozInCkn7Yhqf
A/lhc6W01KPZQ68g/NaNIzvUDC+oEhDLYp5tTuWokkLu7plR5+2R0KQfWHU5tI2D
FHcyR+n4Q+qRW0OG4N309rD1/uQQIi4O+cZFk6x1ydnTzZEngjW1HrCs1Sytilm3
VADELk7JHtaFNk5li4uY3wBU8PiZ/qUWxyMbUHuQ2y+4fzJjNuZ78M8anwplzj+g
00XC6mOfR/+yUiIBp2/hXMvbvOuktkj0umwiXRjQaaQTxmP4JyoR5F5l17NEFhn8
5v200D9zddkJi5JXt5zPI5+Ux4Eq5RKZewARt76wqP6uYXNpPBRih5yWMocPH+C2
iRWvDNKq1CljMfbxuyQGyi3leRPi52BHmCwimijS2YJO3XfETwyOwSJmnUGtpBdD
GcGL1pH1cFzBxXPI4lYd8g6nRMJSyGA1j9oIX+DU++apYY/+tn4+GrEWRq53WrDi
xpfXAL7vG2YqS3/irtCXRsiAputqonBTiCILFbwBxADGZfdRADRl88xrw7dVV9x4
hKnvcTeHZwhz0SRmtxLse/a539Cy0RdnB+Lkdn7e19upp7nID4Hhx72UirvEes20
LVLXzS04Z2QpotzbmTno5iMbJcVTIHOK6HxyXgDHbwjagVGoX+THloghb4Nv7R6P
BbHGQNL8OdBZZG5OjfYzhIRYKb3XnI2hVMhWDZxa1x0ZkHBwgcJpGAhNCvxBG+4z
wXqRRLNK7vvqR9iDEt+oM3000ud+o3a4q89vZ5wNTgIkIXfr3o6KZI0PPpWYRyp3
QFhjpFsvCfz36dcHlG0C1IV6s32zetnLjTeU9WM7NTKzc6Rh5TxV21L9XQe6kp7g
w0L6donQGVpo8uKo/NnCsljwDWgt3MleEFmycIaso1Bt7UlPDQT5oEWC64PU+BH8
O+9wiqA1p4ZVjHm+nsOK1W3hMyYO58z12vsZlLDaurrFEzi4U+b6k/Q714xijtnS
i0Msm6g6mtfY7SH6KMJ9zpaLHO7NBveQbY5VUFetdTDZK/sXvnYyMfQMcMhmSUgU
g+zig1yOmN6qD0HpmkBKFHh2BEVnYfl+PlyUriGHxkQfZeNizs7ppIzptCQk+goN
TxIIZSkACGeaOpg/eCC9OqPs3KUIYXOF4ohfyHjRPpbihFYP941j1pYK8oJ+xywg
qI3S0KGOtHkt6kCHOTY0ZtgqCM98k7siB73/87KSWVYe/jt8PO6UVPnWRBSL07P7
t8jOp54UlxRTUMaZLec7sb9cTIXe0Gpe9PKJt8wv709ki3+Q2O5KM9AHmH74D1vv
zNTAJvfHOuwZA7YgY5JxkKbb/JKEjMuXfKtkgfY3QOT8M4MwQ1Wi5/ybSblYe1km
Hj6aix5pKquW3pY72PvEbgPLUBjINA4JLEk5TMHfW4DdjpUVglKjroqKHu2ZFxQR
AtDzCwHcsjsYxSP9z3pFRRwqIFtyZqZ8MeBbyWlhsl7HA5fNR1Rli0lm/QnEnMQ+
SlxCvpdziTfMCg2XHEBc84dcbPGYNPPH/cGorMa9fuxL3j9SFGfE5TzU5R4yDsox
/ZA/+7ne3+om7njPnvcpccDMWt5HaIbnSiu1E0QQUEaeq/dBbH+QXhm6c3I5VuG4
LKNHN5+CBsQl0SUCmGj671IeTLKPfLnQQjgGMN4MAXMuEoCb/hr1R3pJ22RPWlwB
uhDKqlXE7o96i9eff3bB+SrSeLalkfUMiRMsUQR4pef6OYPDeokHnuDiDOsdrkMw
1defF77TP28m0ZBSoVaI1RPpLlakkLlYkDGfv6QznxYEL4jlwR/ZZZXmF6Y2onoh
cCDG8mcRVjWAT+AHstRqr+thLfTqbFSIBm4tyAOFz1Rq1+SogK3JrtrMYLfw2b+P
T5yhePqcfQzq1DPO5D6H+zkM4dxcHmrY+Ya9voGSx4Wt5msAKYznUuzSdXjyVxLI
4UC8LQLdDXaPtCMM2T8Zj0MurQPpkOIgalZdUOf13gokM+7Hc06/IxrbrGT2X3uq
SvgDTrdpgyEEpTCypae1Euu+tvxk29R+M80q1MOOr4v5wGzvxEOSUSSB2PHwb1vk
wJp+qa+POjtoOPEzvNpUYxi40Cc1MROdRJTe0SgKUA2ZEsLYgfUwVXLHbAti4m+i
yzQuQCsyKydqZpL7IivaTUsl7933E1EZ9uR/zfRXpIQVcUBR7iT7gWrJxRsNEgHQ
+4LZ12cdKA7V1OZF7IBt9jnUXLx8TIfxPseFBi8tECa8ffJPRmLWG79GHaYlunVO
Ro2PAVqGeEiDZCfNDGcBL/nF4XMA3abEtOms1R278OA0N9AfV4eJmU5Bic91BPtX
Ae6iY+MzuVzj7UFYeHB/PaD46C5UcUTcAISH2T8AzZ7OKeM+QEc8gQBOW/wuZDje
p/CDRaldbQa3u+5sZI1d1rwMfBp5vs9ILzOabli5mzw4e03dqH25Oa40WGhMQWRb
NIJoQva9FxKhjMLf0YJpWTo8ETbKl1bD52oJgQQsWxS4yUYX0tPFKg1BNEoGBWSX
oIPTTY9zNEGKSNQtqY9TEqoi3+KiB6aVEBU3yRmf7q9tPiI4zJkTXsIU1n0O5vQw
xXeLCzPtCJ/k14tSTFWnEBNhFdeLyUCgMZMONCx33CAWBqHlot236wPzOmOYkAlU
QxAO56JudFAt47oz/W/Riyrhkz7GsshySbi5NVagr8mFTm54A8S7rhoWizfggTS0
cZcOzZyIZwUUmr07G1NpfOackGFzjhihm0xzPgte/23UqrJZMolfJMydSSYJGXSZ
b6AF6us5RBt0jWSuqpCn+H4lWnXW4PsVlOV6Fb+3X61z4Sm2k1IJbPqMC3jJBifd
6hlrXrODyWba/ogsWbNdcNjAYg4WY4rRI+DuL+O26YbU4OgDJMGIjl0FePPVq66a
JyIeQhPfI0u82ukHQM2JraLi6dHhuXtecIewypaj9k1nfL+kxwTodnCCNO+Hz7a2
+QhYY7nVPaaTMm20DOT3VNgu5JFBCWlmXnVve3juZmoem3lGVFVpI8xRmNYC0yQM
VFBbB67c9Qupw03N3Sbn029INvl47cgThgzcb3tdwgX8GJzWUhCKRMEQkT1jNHUW
KSnvWfC2riRJZC26VWPayBCxvTjCk/YjIwUeSQ8OAqelMIXsxDHDAcS2toI8wlAc
A2/y4MA7M5V1a0HwASPtsNTJwit2s5WhBl7sXdm+QTiZ7Oa+wwRLtNNLuP5qAlDG
ae+lVnq7tPO49JbyeVX3IUcjLf9eaNtQVHEk3IiVtXzR/YBWwBPUOm3XNbABL+pf
ZjRutQ1ui7is/A7rTUM4IpIbTWpohglx9uMKJ94ic2IjJBLs5GhQ7MI903AO+jqM
oYSUt7jQ6V4/+DdUMdJ8t9Hf77AyVt8HJX2ZN8bYQtuKHOGYOollcQxHiK+7enku
iInKXQ1MtJ9KehKCxEyjAbaFnyfyEUBDNrnBjUrpWDoP2gOki8sTe1IairN+YLCV
wONeu/3V+Df9gntcidGy4bAolNc2gO0qpKgtkKzqfbACFsuixDoAmvsZ1e8F08d3
DxxYDsufrEUbmORfX6npt2p9SEmxuVJcLMx/BsxmPdmgSEYAuuKTVctzdZXmJoYN
zRkc1TJDTsJBLQj42H+X7mSm9+gh7b0IUX2O+SLguXaVESGRv15opS3keHBr59ky
ptBzpD6goXJuAgzP1v7xoXkj/iyFFpkf9U4gqwKF+cqh1zg2+gFMLUk+6HN2LDM8
rrm3cl+CwGOf5M04ANHil8vD1Uam5U5ZcLA+SZOa7N5M9JDIwvWhhk4/bmsaKeJd
HdgJp/BYQLxjD/qnXgyJxNZNRs52zUed7t8/nnTojwZor/LgOo9p3cyrfn1vZ5Oq
iCWf3XSaKddPz/XbJdl3zzUTsvkcDnP+G2VeVUfvW0qvR9sOtm4X1+Xely7y3Fc8
rTWc80Qmu1p7oc1FBsfx5q3MoZgrYW8Jk7vRyrBU1l3NcimFGc4rKgMzY9X13pD3
maE1toW/dN2xp0RoRlLPYO17zGkgVoCtDZC5jFIJSwhEp51m3riNoS3mooN8A02U
SA/Ql+plIlB58UH8tN0tn8KhogbHAaCpSPzY84+aCMSPNfBqVK7RiM5oC8Qf6YSH
bH54dLVLeervCOCTFppjspclETISlxHkTslt0GmdhCj+AzXmTOOGz2aw1+rLm0Ii
qEdG9EVdU3XMofoBLa7ZVm7aTzoSzy8v5bIvmyK9ydwSWrXqsdpBsfGFlD0kYyOA
Z4JsRsKs1dwCmiT784/mKiMOdJDsmvgBG+uDExSaizKYxzEzpYYl/nK9k0yhrB6w
i6oQZuTlK9Ze7O3ZixKEGYJPbpybNK83osINrBvKFoIHw4+QlVsc9atVG8Lzvg+9
g+zFf9Ai4GDGhZKYlI9DTJaRw0IzVWDKzgXsW0AURlzBGsj6Y8yPmy0CkKSEC5Nl
h92CmdYPCuygW/m5wj3a/ulb98rrP7fbHNUTZEwI/pVh/bF3D9pKlDs89Et7eJnT
I+2xd3cHqMsjS5MIowVQQzymRvhy6CB48uf08D6Wl55Nx43+nGurs1hiEI8VSF/t
ncNthHEAJFTD4i6d14pJL9bXL3YvbuCo76tSWJA4lnOVbRZGzhl+kdfNbUR6/quV
CrWvAK70KlbvbXucqPbD2Z+yXo9YRj/P6MV74WjhM72YA58wqnyI1EgHupaFv9jN
/4DUBF0skgqxqhepHL7MZWcGvKwrK+u+t3Q7TfoSxcwhJDZEFPjZAUMXblVPN5pH
88fppaIXDA1elXLBfR1Kubs0t+DpGLFOf+rZyK9/LW/d7cu/M0dyGVFhrvBp3BNM
l2IsDlUrTE8hRH5SDV7eJyWFC9FHHdj+CS3/6rHMjqaHpiYsbxaoq1ezvfCesoTw
98pMUq4vogVK5Wgy9TChbe2ACb1FMcRNL8z/bhU9hKAknsjOAOhSFmQ8ab7v4l1O
OCeo6vd8HkCjYs/PjDDz9hlVES1lBcElrphEt3j8FMBPfd/v1IfnjWs0bizqImVn
Bd/tDhWpIQgEDSImR1v2CQURz0MvOE/7xrxiOswbvrMPqbtHMSfa6TEO442usk+K
5x4yAQYxzb3nPDrxRXnTIUX5Zrmo5kY7Fe1un978Pfb/Aq/kghF/RwOiaJ+oODcI
+mb0K4We38cJZxgavOU+OnBo4wQIbb0FzvtpD1DvQ/bR33A+kZbK6tWGlH4Iu1oV
QEiG4/kl8zxTxb7jDZ5eRFv/cR4ksF/Z0jywnxBcazBZGGUfV/4tNYT3NTt3XLJn
vq10o9wOsfLlIuGrSecw0QpFmNFVsrLu2OVKc3Vqr4eIZEqKwocSY/TzvYH9RzlD
VfMgbPj8Inv1TqF3URAwKbDE8Uebo6ecg+R3vOPTkuGud/6sB5qDjD4MS3zGYRIC
EVS8jhUErUSBwUFZtruscazSwZM1rmI+4ZoUz2+p2In8zCNKCMFhprIumOlaE3oY
h7ADFts1RxRgdcpaA/m4jTgcroloDjQpJOh3LKA8qprAO0Iwkj3fD39Gk0II4mtZ
7E7HFNDc6PntPZIOexqjJ3MNlV+94kd1i80ayBeOWodhpFOmMGWUleUwr/Vr3wGn
wDOO7EmS01q/faNEOl2qasewyalG6PcE9QHve7gwRqquWhXIwGcMR73Cve+c73b0
SYhienHnRlYfle0rGIWuhkP8890F+kCvCHwjmyySOScM9y9A+FPpa/M68A9tfeen
/aXVtxqMkKexJyizCWjlZAlO1oT6xVQC2xCHEtEuyJvm9bV6xvbFe/Vgtuhe9Ia3
zpl1pT6Ld98KVEhrVyxUhB3fri4+5JFVJa2OLiBtUyhUSCGJ2oyVGvVt0TjACYxx
UWFOpSp2EfPqYXrdOQFb6JUmoj6Zn2Ct9fIE/Tv05yWJtQiqCsAx5Zk0LCc72QaQ
dnPSFVeRajpWJUjOQhfYxzkrbD5XSBEfjPXhgqB0hkDyBy2uWnXNldangWyH0Jv3
twbGRAnVY7h4aUpDr4DQM685lULXskMkynG3/intFeMmegCpfzrMx8j6UfP10HuE
6/TVNOT8csERdG46S4BBAfst++pmPWEcc4bdxo2yTn6Ik6gQOghNbkGZXkkZKQzr
uhz2lIrKe6Fttw9BSmYIOsjIRPjPb/Cad+HS7aYJmhKcVaD2KshOxr6kg7rpejrC
lvP/MuZpnEPPvG86Kk3Le8sjXOGHwDavJo6FMhFtm/8P/TzY9vJrse13vmHzyJYU
WpppA3ofLG4TwYd5VbOQA32sCMtyTl8Cz6DWqhblCw4mACa+q5kZymt3wWq6Ly0x
xsDqjKPRZG9l7knP9pClO2/LifjLm32uy0qYNY5dBA/YEQZoiI2ntW+3fdLKrMyD
zpXOfBgehgnwu2NGYhdi3TuHV621yN1qi5uhMCjpOI19TgDUUEifojblZpGMsS6z
pf7oPz6p8HolbrUzCk43Q3bBo+3qYo/b7BcMzy8XXcsGiSm/9Y52HgGmMiP0z4mj
dCeacEAqu78LaGIbcEonIhZoR755gB2IG/4Qj2liHcISgHINfiyzVG8ENGfsEPCz
/mvepnIGgTseys/eroa3IgsVHolT6EOjC109Q/pU12NDlHI9qUNL6oGhWec5Wrd2
/y1wcRdJHeuA/WTN2ku2jqOfd0OJKnq+sAFxsIxVcVgC3ohs3QGRO2z2hc3ckD56
W66+50pyP6j1DjAnHi3SWtGoVUSpm5KB2kZFb06DkfolSWMgfVg4bDIYof3mPqFO
G9bGW3ujDbsst2CfowoQ0Oex635B+X/wmRl7GLCB7VhoAgdR82xUUhEBxoryjFX2
8U5/FE17cyO9OP5c1WACPQPZ9mIl3TXLtue8khJQpz+G08dcnVyF7b3vBZlvcoFa
1Uwid+COe1ks1tX13bW5+OrsUIPHAWWlARlcC7d+tKQvZYP73rw0EExET0KOI7yW
+p23XqBOXu140h9Jptlh97q/zC0Funh8jA0Bipak0owbCqc3Y/nAcRFhqq4W3xhL
TPPGo2vnPMIPGWXbnfRQ+8XRCBk3rKL5Zr00NDI/BH9dn1EILz8vVsSb3G/bX1T6
GXx6u3WCl9EXzVnmSkAu85wIJ42kXgbLUYtf/bjjndD0k0KJ16Nss7G/ljJi4M2N
H1J6j1PYGUCbpECnJtJLSaYqCh+Lhx15i243IGUSWRxXNRSN8XKxM6p2rLAzmd12
dL3Tv81yWOnwy5nt6XoYcefiQW9pBhz4XU6IOPLjAbobU4MIikr32R5W7uKY7HNp
Zx3bRueIj6k0vHS7ccc5DPhmuglZNLBV2SdVUxFXE8OuEteyG7a6LzlUW253+8Yr
h5K3pGfruv8rpGYFCSTkmgqePzLgch4TyptiLxk/TZbGPhuE352VNTj1DoVN5F2A
yoJFhmE7yMCJZQjE24N1ouLLyhNid5i7g1utVnGfOA+pdgFt4xCF9vELo3I3TPGZ
xDVUu4H4BNblH1SgprlawVPdOLgNA55R2u26EGhbE9SeUT2YF3xGBpAbSGTFiBCu
85iKPF24tFH9foF//ZPMvlQ8dbxpegK9FZRbMNbvHxAYXc0l/4mgbgrKtP2wBmZ/
R0EztOuzN7ZRe0XfJ9Lx6P7Ho29p9jRxJ4ZL1tOs0nsSG/0oysaUyxcklQgcQ2vJ
fVbSqV2icHukM/Wn6MSCxT8A5uX0/k9DSdWHumHmHQGYtSxUnd4mlEzFGiRPBJ++
NOqcEOVKdNtYWj2CrmEg15//785gCNuNF3uU9VBpdPQ3KNCGkhKH6GpzkUuMWIEN
SKtlKZPr6+9lmsKoZFhix5V6IqaYFbHDGZRVcQw1fAMyxvwiEbL3OWOK1/9g8wST
lJo4JMmZPp8ji2fnU5Ek2xf4wLzDeVeyPvaF2VKEt3nY70SazC+GgNZiK2IyBWWj
4Y7cGd7qnqz8s6Vmkz2BeZjaGPV0lHQTCk/TQ6E8uW1X0xdSMJH7EXkQuqsVXm4d
1DHFtrcnZEzebxl+niBNtiJpj6gIsqn78BtXmV40s6cp7DNxKyDaKQopcTus3yH5
FQJ7DTLEHt9lcHIeWJJMyzT7jAYDpTy0NtQ6sksUrQV/ALOnMvPTJkgDw83qZrWa
0XVhTXKU+BI4SgM9xeaGLIE2BZdTDk7jZgWC1PVdMFCD28al+77gJddujnC59Op7
DB67fz4l8R6wY1+gBpubIOQNXYVZSNiqi/8TcFFjUvBkuF9OhutWrRFxCHx7ljUL
nzbAlTu2B9qn0kkdHrM3tAb//jPPhr8fAW16zRnpVH7TLrkiR+k6Hi+pbY9Ztyeg
tiI4Fzq6mluQdTM23c8tX+MeBVrMOD1zP3xKMrEeT3R969u5lDV7mg1RbsHjadnr
tKVVwloMpm9keHNzdpFqDbqGOrRwgg4P4tTiM+cuJRXt9zCqmj9yyftNY0d6wuwK
AsEjrD1F0Tqo7EQpXOAlv6H8/GkqD3ycpT2ZrFzDAhgTQZNLwuWkQ+fjAxQGfVWO
UapTiq1e8yv+gvWB8KNjGuBltQVEmFB3XtoDzfN5SdHZvnaN/BwgnB1TA8n8IvBc
TeFryaV9PVNV2T29ciR8aykh9VKQJKoAnqpERIydthX2nuab/jdQYpIqyJaMUV/f
voRLHwDlQE6xDXpxS7K0Hip6BeMTL2g8BY+yySA3aah7roAYQIAsIHbMnPgRLYUG
VPvktMnuoz3dE6mxl4npjNiJ6yWIh3IVBE9hJRPkWrz1WjoLO+GepB1ftGYUwvX3
FXL8/JzHJcN4fR8TPBRhyE4jQr4W0FgDeztdEk4sgVravtpmxKloG8M0xlgoZZ1u
H2pMInhyvqaEEaBJMTEJEp2YwBFXVMm8It75M/Id9zYa2LUaQeIT7B8LmNptepVB
mfyoqbASVABS1wfLM+f3vFKmebt6JrNQkpaqbG+z1cFp3PyUCPN4C3zFkimPHwXo
muXYlQzZKLigx9DnLc2PLG7FaIJvHfm1Rlq8J0UAYeJDTwKgE7Kcj7aGI7URtFav
ftqhfW6E29M2pxHLsnFxZJLHVqQSUmtwqSINuS5//aISF7p9n1Ko44ujqtGEK6eH
su4kADEYnD3kCB9uD+XzKxPWuLg58aYi5DZJrtq1OwOD0E/2A2QCpfZnigy/MAg9
hrb0c6g/L6PuSxtt4CzsNBXHS5C6nxfCKiD05QTWfWyhC7RLNQtwe7UGQ4QE5SV4
97BX1fNGGbEz0QJYOMspMMDuGYLCNWXWpM/GyuJXJfEKFzfheUfQpACGPGZSGiti
7HgWnO3AvXx+DjK/igwj9gPZdCsti/tdAk5OdK0YikBQhrZfznOvYboA70gCOIb4
pSlqAVgO4BFWgSOpwW8PVN7071PXARfad0TokaZIN5kCKcKS2D5pSPG7YbijL+xv
s1k0VgWbdDYhPMf7rGuGCfFXRTyDnzmmDijSc2MSNUdLcjxuNRSXdEd88eYAy32G
ArdGuu0WUX0QhUwkvz2tT9kAVR/ThzlOuCHHdcoDQe6pT0W2fnsJS3qpWmqoXvZO
l6HRuNYmOOuNTSyf4pgC0f+MFH0cumcJTwUaBJAuW1UUVBMqdTau5X8VtW8J5DAZ
FOOslFQ8ApgnzCyjCLANg+2O39LCyohJgoa/qQWl9JxTPUADQXrgYcVj0E84loSr
BYAMAj8jVnsyOHeB3WFlgVYxL0tsxW4oZSa+18Bk/PJJiQKi7lF4i512c2XuN6qO
F5+lfVjZGLI2v/3Z3Fpt6kboaxD7pny26gGmF1Bc2bvbCSEhOFcnrnRhvhe1uCOW
3sHosHoLfxNYeuTpV5b0gejhKpusZcJmya2KeeeKg7Sbeow2a+oQ4ji+kvgvFYgO
ySnP6oRg6HxtNUr3Wc7e/5bA71fmDrUrSPZFJbxF9T2qQqYmzqx37V24C2NGYgNC
87v+/7KAwN6NSvTPrh68AfzJCeH5phEMMdWSEu2K09+gGctBpaKqZNdn+H4BZHN9
CK3ZLhNW/fceYtAFhDMyIxZgdfaFY43rfjqOA8bkGHC373m1j4bAJQhpMK4GuBuJ
rGvF9uJAcIbpaQ2K2F567jcWaJWRgr4LOqGs2pTHUtaQkcusszajuXuzya21fMNK
CxzSN9uk/brr3pue4Tyso2rPCcMelfLCGMwJUF4LVuO/7z89gc3j+MOkHe+6P4KW
uaCrKDvYQo8RgjYIAd1vazjsVH5WVC30TyFfIpLFdgOkuC0EVE94dTffZYSTHIrv
fvDIcyL5MKLN3MnxkwUlEWt9973R8Gs6n31IsCAenwJobbJRkXZdqAp/rdp1w83M
cGLC/t6umYvvxs6m5ooExKgy7uba0l+rCYLRhUjLv55ySrAsEjdYxkIhTr2fFjdj
6iif2Jls/3VsuBinXAbGYaJDtuaoJExYtHdlua3dpIAbnpwX0i7VxyLRnknOV3HY
FWJkjTD3Qz3jrHLrynCD48ig1TdRlPVrYEL8Hb2YNgFDKZugdB048jcP2QHAON89
0sLLi16eR/WLVTg7uk621xZ+gYUZTndAD0CAHZ95G0lqnosL8dy7wUtSavwf8CZG
pSRn5iVipVsTbifPmLwKjhgPk8QKcRswmvC+zKnKNa+2a3ZCQNgq+70i/vx61PJJ
qTGBivqV1VJ61yb13SRlUzh2tAxlpMqmZmejngDTzFMS6OfMuLLIMC+UjraSwCBL
OtadckjY9KOrs+oq1ej8WXQAUpjbt0C0aARd997aX8XJQBaeFUVVFsUl1ovH4rGl
sKB5Bd4nK9ndzi5vh1jdSo+kd9OoNvvMUCzXip65CU1GWtQ7JSVJnvwcFFlAJ9gH
iC2rLq5HCdn1xxm7z2jHqNefFQRJzlAEMSOEVRxbGWw2QKoFlJZpG8R+mTDyPRtr
2PeleSYZlJZ/bowUZufdXYwrPpu/Qj1E7RgE6LXrXJwZpRHNgHwotqRXINkWRfBx
Ls3iiordkBvmnTWNWiG4i/dVz1/7QDhn7lPUUM3/kcgsYlo0V5Ta2CNwiB6wEu/m
Px7lvYWpJIKz8WeEnLROffv+BGfDSLltRVZv4QZxlMnXXTeCN/GnEaXkO6p00vSM
BXy7CncYCkaUw77Ul2h0gSHnexah6QyYuSGHvThs5WHn24LhHBXI2qeTlEsidriy
X0IWvuOK6URfA0cVRWz3FaS7raZvDfUJkFkSw87BtZlZx1cBXelUv1vknDDPQAoC
ESLlJFAeDsxkQ+ePW/50driKSCA4zq4DIko/pSwz9WWiqewW7PpaCRi2AuSf4DzG
f1oYBbJFu8vQ4Tcu9ls3Vg9q2UvMgwTRJuXjnrTEeDhvGaeh4XaoTrsGwYfGD9Iu
QxUpYKU/hE4COT1CxlybAXJvWUjt4OdIdqAhgVQ9RDuKtrDNH/wlY/SlakO3i8Ui
D3FFgp2Qea5AAJbQ3I0MJ2MbD5IoI7/7pfcVGQAebBQuhkcONqrjrQensi6IMRe+
NFpLaMOk/mIMq7gRHXPdGGlyooXkYn2mAEK1IWFGcbYyb+V7pjfqMt/ss745YXY6
5DixiuH8h47/UIDI75QZrdrB1sioWBnnd8MYZziJYPjEoCLFNc+F5nmxK/Kr32Jd
TGCE8uhWO5gbd81uBElDBefiD2gOCKCXevfr9wz9mSSbYoS1GfQftqjB00X4tPUW
0v1MW4wrJ/MXIxG84jsu5BHyFHfJ00HXHhIrjnEdgy7If71AtdSRWz+ts2KjXmeO
fM+N/WMeWSaKXGOZNleVNdrUf2T6COEfGKT++PtkRueZwC0BOjKsm8tUBNrWMWdi
+ode2N4yfKATz4ucj/1uLpqaG4JJ4e/7t3bbdolEdSLafsPMuKDDb3fmbK48U4l9
RVIagtto+A73E9U6uFRVavhmUR5/VNIQODUEioGFqXKFH1hr3JwRBrBhBrnZftK1
fT4enFos/zxa+HlOQToeBiu5Snz1qh7qLUxyYrmS+RxNS/l0hGBLBbGU79FwnMnY
cO72GQV7qF0UsM6oI+jSbLpQ3Ch1bPNB7W0vUsfRLGpogjZBspGgL7OK1IfqjFA1
wV0xfwUiy/1FfHoKgsdhW/gYCgQWzPNvaqrEJxa+srkU7Ui0u1hXFU2HC35hhUWT
p5dHP3L1/TvaqPXp1VN8rjLl0gEUm/tDIJ0JZXtCE6RGJtaiUPjSxQPee6PuSFgD
X27cEU5JIV0Zw1BwRRktBtmFr2IN6KHeBN0l374o6CHhLXVEbBzx3Q3/nzqRVd6w
STlEEeRNZbVDchIKvHVXhZISYD1kq9VX/vdFYiV1fldsWlNY4Tps/QOQWfgm0saN
CuNFFU9hMZtjEduR2xfvo8x4DpCTzCMSACMpTvYPxqUDlSe7Qe7pLZ//ZiPkEH3/
K2xFBsLovjzKsUUov+BkNd8Ij9KN/4nC0HdQV+/3rhvPI2hU/cUMpWbOiVgS8zPl
nDiqyTSGf27PT2wUdUGhdHSBl0KnAMHOconX6uTdzEZHWSrnTsVDr9Udt1gzVoRW
vvD0p61kHbNdep5MWpUdbNf9Civma9BD4JtDw5irNdQlskKRKHoeXRvBwPBERkuA
2/7UFOZp2YLIcS/FPLAm2REHJI7irx3gqaLkrt2lCg6K/nU2yse2l1k/5KPrVa9a
t2B9kuVrOeJ9+SPU4yJeN6UWHgNofbcKlTyJfSXuZXDgBEV3G0WVdIH/9aya+xAe
Lc8Qh5DT8xpZV4icUasZ859I0RfMZrabdoXa2FexvUsy+N9aXJbGr+iL8W7Z7PqI
TXBDJRtgGyvXAoW+oRtL8GdrPr9YRcOuQPGDc3eDVVPcl90z2xNj04ae5fG6Vali
dfG18UjF+HRQBzaD7iaA4EE/Q7ndb6C9G2DPGe0FNxqy2Lx8V016ornWyYXC//ji
vXVPOHBz9g2QqtPtioO/sNIjl46DIv1EZVrIgamA2/9jVhBxz/NszhGQudM7dq0C
PYY4qN4iorHnnKgOqIil3QIFdrwbQHiBUfelwEO3D+fv8kSJTkuP9pBAdUy57qyC
6P5gMqDUN1INntqys9l3g2WgOimlBh6a3kpJNfuCIkgBW5SDPbb/2kJmo7eenKqv
unk6Q7rx+7QgdxLs/Q0ym/opYvSfMzAZRcQ7KZj0RBCy91JfZTR9Rob3YQ9bBwEq
qLOSxNWDbhrsLVdNxbZ0bmvBJUFvL/ubiG6qGC4E7Ssu+TePMhFlX9if6gg9T8l/
38ltiVN4wrFNl9b+b94HwafZbM1CqkfpDzY3fhlO33bRmcivEM+zKyq+A5ybv9Cr
eTIBTSqvMDKWpxBYqbKzJPeQc1qgWF0tvzX4Xh/nu1rWl/8irtFEhGwlHrlSpyM9
dFLcKyPM4hBCvPLOs3/y05DI1C0aYdPwdq+zTAxwnOL+vaEEo6cennejg0gDU2D1
mWHM1Gxff035VPPvczjPBWuM+2aazJtuAHphdvjDnLA0NPARDMe27MKGZF9Bl9hq
z5AzoIpNGiA4fj/sHKSXYMiBIelKdj6P637N3m2upoaQCiM9h8xdCGsTjQFb+MRq
/bFGy/IbQ/Y2cA7AFTTDcksZvtraR8YQx/RhpGR55JPyN77M+x2VMn1jkH/YyqBB
4ZUDWj+krY0AGenwfi7sOgsbGaWyDKgLT1UYia885jcmZR6sEhlp7NFGfybdwBES
O4PdT4sRwPqW7bL/CC+CrXoy1SYth5kV9KL6zxhtQ5bzNO+omUB184cUhMKUfu3s
34RjuorIbCZOxBeWeOHDJ00129Aw3p99+Ld8RvkeACZqLYtYtbZH1FX8dF1JK6yD
iU+BqbdSNjFMBxHhCD7MJY/ic2fWqlbCZPNxc8fwRO/wBmTbvw9A+SnETwOu+YIv
3QYqKlG7bAd92jtNxRYlJteHglNpRO01Vxk56CTo8FugR+A1bC6+VHlBTqnmoZTQ
l4ob1nRwaGRkkWRiMgJLdNLIWIzdC1pWVu7jm/43J8iCBrKAvC8DZtXIBaC7WfBO
hY2QMv86efo9ZLtEAIZXR8RO2tENYlVpofXECFkVv42I4tOMgAFmGvRb8OarNBqM
DTR4t2MEpBHcyWRLnBzd2W3l/z1LAwn8CIG8Ua8VkCfqT0FcjheBP22qUcCn+XzU
4gYcFCwpQ2M3BwaPcT/DDYzt470eMjK3RbYTfO/3wTLuN7f+1IGxkc1bgSeGLdCL
2iTJl8cmqCds0GuLq2Sgg3jJa9ocPqUdb0DcEk2Qqsj4IV/Qd7L9e2WUEuwiyC+m
WlA0bbtiLJjcxVLrGogF8S4S2ew9helHnckJJQklSehwHyTDytCHZa+YGlve2FZ/
Yr0KmV9deH8jwJxikZEMlVVqYH5k0qStv1dixM4abKfyoPzb7KGKV9SKYFNBhGWh
jnVqiF2cVuWvDpbbZ+meagdifHrla28KG7iNcbU9jXe3Uc0eMTSLkK+6+2cAOHuV
J2Ch4O3nK3gQ2tm5yTjJGtJz2vSbm4BW6HsYFfC0avA8Vbn5lm/VUZujzxgtd6Dx
Mq/lEHOCU7ALPqHEKl4Sta0QD6xZLZg8z0zzd/qFerRfiM0lTKffe+ZNlqwidYIh
YKskY6TFM71hGawNXtQohPB2jDIojqHOO9mI4bXs0irvH6x/f39QQwxah0hVPm2D
iYDyI0r7T5mI0ExkdKf9ANB3ncOFi3VOMCqbzBI2KCiBvN+6f3EcqfogwYJqbIXg
IDGT4IlDG3PHFUVisZHcOeyAQ1RV+huJmbZI54Ed7a89u6yEHA35CHFQA/PJ4a/z
CKpzAVOE52kck1LokrnMiCwL0uActm6Jm9h/oaqyouTSxurN+dpGAn1AZXvUycgx
JUSHvzWFRrM0FwJ7lK8CKeJ4nrfXabq2p6y28xPaA4+QsZqrNNXCMjkw/RN96YPU
o2V7iYpZ4ZSZeFkBh9iRfTxxjOSrvcCTx+eeJfkKBkg+OFm1lFK1EQqp+EoRonb1
s4EfP7cVZxaDrW8U12Hxolj75c9X0rI26qbpCAxke+odmAqPBayRYmzUKn1KQBdh
4UPph2io5mdGNm9MSWdJUlqKhrQiFqJDDOKdeGAOhorAyEhEkbfdge+NEeU+O7LE
2L8NpMeUdHActtkBhXMgZ9PFRRBe9e/KW/k6VpOuUreq2Dm195wx+e9ky3so9Qt2
UzJfSf2ijH75JrbhJMTMDCZSGXrLy9QDWYbBcKMKq7EGSjKqGLxJq41G0Pz1q6CE
rJJR3tkezpFXPyoFUAcoJaC5+DbQg0LWvzdPLqAtlV1bziy+TznQitLn72YHVW2R
6ro5dMRCP29yofKPCggvbEsxU9hVGvNaegnNiFTmpGtKtDhQym05jf/E7SCeySVY
w/P3pkmQFXAhaF0BhEftXQ0ewnKYgeguZpfQkwSJyteRURLarKWNDgSiUnwNrKIS
COWbe24D56lj/GO5UVg7eOy5erxi+sYonhYk94eGtMEJ94nFLWNTIup6lJ3Dq9Ps
yR3Lz3VG90QzEStWgQ1+hwTY2t8CinwdqzZFcp/BDkudrGOuhuJ6uoRYv33gnqgR
0LgwRcjf65iRogsizySSd7oidwJgX3p3IzxzO2TVcMVrQsvwlLCqlfel6O+TyYLc
Q+WIjUTHmM7FW2iT0TO3j8PgVGkotGTBqdXde835WdTv2DSBu2sOJ2Dz36J/Qpjx
QdgaSSaND5JRCfZHXT01DFBIQHHgPIpJDNt0JrJENFlpitglWB2uP8OoqRCKNvah
sjNS1/8DrrnWiGkCHoA6cJDLjlSW0lQd8O9lH2uDSe08BA1TBiNKV/YpvdxEfygZ
x9gF3lCwI/x30zr3yol4WdiqNyXtxVs64TOlQbFHLQGw8NLOVB8ZwcyEEwhxgjtE
tEntzT4szH+qvBSIIXUvSUNGeToDHdEH4j96kopuYKRtLAY3TqKG6cVPG2c+pXA5
JAaC6DZofs0u7EzxFcqo90VzN6mmarkQ7Es3OvEYjwPBhRN0YTyuF9lWNvRFQmmT
3lZYxl1qYboCDLgiyl2AYWcYs6w/lqhmbx1SDG5m4+2y+nQRRXZCkcFKuw+sQ+kJ
AyvDpJeaWjooSpm9QFNvS4gZr4ALKAtAtYnG25rLHaAh0cmW4bT1/WKxUxD6d4RJ
gAKCuB0AFfHBCeR+GE9gznHpqtk5PIZ05K9M7jyslFDykILW0HvGkYpgn2zux7r8
BBkSAWgUNK1zwDXZ1peNF1qbI9OR98GmjllDKHBeMgSF6TGT/okrrgoHw9DnfZG2
NdAbzM0jT0sN4roE2SVm/P08LjvaZIumFg9UweGZzuUYLCBEzW2YraqeiimqO3p6
Kqg2wzLQI2DWbgpFoI5OB1rUwYOdNRQ8mLUuBxof2Va0oczzo7GHcpDn+Z+Qf0Ai
/F0OroJ0wHu0hjLdqUGfe273SDUixIMfpa+eBEJ0TZHWRN3n8jWZAVwpcE5KrmGq
RT0nxWGg3nTIhzdMFZBHhZMbsVF7VwGzs4ChSYgK5SugsqT1V4ZP5D+/sBlonEoH
BCWtw8EnvS13nB+FJcXjWSsaD57EPT9RZur/EOfe9kJM0w3flw2XQFe5xhdydUJK
d0vNwJf0YDUJqQRatVl6P7SvUyYIfql887T3+AomXmj2pDyfoF5akrECHrfxuqSz
xiypETUdemIDUyyKUVHFl0vHXQk4sQEWIlFh05tuNK/7w5B+PpCreRvQRHoL9S6f
HhebQPzJegj6IC+2xHSfYjatYj7EfWHYsw/O8Wn0e+7VyYW8/oDB1dLgOXP3dd7P
59BTVJ1j+2CT13xlvw+C4TFxm9YIPFukn6EweBHjEXicSXb/nNYiBXldIEa5an0c
DzerbvS6sk3ctg7WRHgdafg9H6Y+POiffcbQpxvjqyYAEQQSrWksf3rG6KCf6nEC
Tx91JY2csgT5Xd1p9WG5WzN8VMOADuys9ejTAokylG/UC4yniogei8WLDa5zC12t
DJk+PBT6o85l8tYZ3PFrclN33uVU0d4AlV/TN2MZ4XB2NsqvOFgA2By36Oqf/x9c
W26m3ttHOAlkAjtqEvXcaJjeSUIipJ5HYcQ3lp3/ZnAr+odzLqDlytP8tGXzXAUS
y2qN1aSZjpTOviRfmT4Kv+yBCcPCSDpYISW3TUxKFbOCpFGqHoHppAaGjXm0pPvZ
RieKUu/THW7i9A85kM7SxFPx2N4qslM+/TWX4d87MWH7+vtI4Bp8qDd2iBt9agKI
QOCfhZ036tDvDODSrgCHXYHrIfiD4kp31Y+gPwWMKC4or56aEkECLSR7wngygYll
W+1jqepzIKubSGXKYbDJyvQyPLigFByusWJv1v5txn72gelJL8rv/XbuZy5LeJdg
VHDmh4e2Poy5BPjknyKOYSVPqqHL5yX0IDRtudpjqgkaCDj4l7z48hb1JPIe059+
4HCzdVAZONErQgioI8ZpHxrc2C9tOHW+ZGaZzQwNY7u4pgI52RtKlm0DT6S5mvL6
qOgq96tdrcsq9xMpr2JDFdDctuXyyyMxsETfrNF72Q8fl+BE5OyulGPdle98b1Sl
Nz+d/shpIUezZozEw/8/lFJM4ZtsTVP7fcgoTMPSCaoVom9nuUp7H8JINRbeetoI
+7j/9LiQhErMDxppSP/OQhA9tCU8HslU7OzzD3UBVstdFyxUooVGpvglb0Tj5uGO
0cpktRG/jnFLRM+U6wZnqHuzQhJ+jfLa3xH/zNcf/T3lZisqeb59XOcDoTF0zBGn
ChBIhkmhn9OHHvbqFxrBLkTLoQd6YxssU/F7dbBGDoZ+g4jbVxVIIEmsvpG31owF
Fj9zi9cyM1uU5c17JaH4WGHKWsVYPCOPktoHOhta2t7ZMk2x9P09A4DOYdGFBjOW
E4PuPH8Lc4bDY+GmaKTxgRLDWl23kMlaQWNrBj3fbzB9yQWSeGLy23lRdQYse2kJ
vjegZQIuCdx96gpAeQ/pBY72A7f6nRw2ir/bsytnIOsiXUscKMZsv9KwW3htwWKe
M41Ym28sBAulj1fYIZcI+UOJUxGNzMoWg6Mg6Y+2WRGSDPNOVc6HLMv+7sreHJd/
UWu3zIea4nGXmYpGYSF2Ulo+gRugInusiPvOAvtW+DjfmJ9GmLAp/pNrQSW0+3/z
UjQ3Yr+Vb9Hk1qHjPnPMjwHYqJ8NUN39g1jQQ/v3HrwHBoZR+9d43uAVrQzw4625
nWSsA98gSr2R5agP1CjFnaia403Qs6SD6yW4qFBgAqCHQtLTlTkTD1vFS8jHvwDr
XV3LGpCoLdrdvxEcKXS0KRUzLym0oOQuiJGsl0wwZY+E7dCMtzquc7d7ZMwFA/Ul
zOf/PxhscrQRLAkw/vIpTOP/PoT73/Q7ZbGjd2asGHVe4ymZwQSgcLAISu8h5+6R
uE6DHpDrsP6Der0sqJA19JKJNSqh8BWI6zRxWBMK6PLyEKtPXNOz++DupnwisaD+
3OEyl2gbYPvPiAxVYgw0EdES76RGi/t0eHsA8aQp49JXw2YI6BcqU7FtSTLhDWNU
T2/st82su9OX4HHMVKcnX804tHUZY3FQu9Xs/sYX9lghfHSE5+PD5FFrhYqHYRwc
1UMI3Rlw70tSdWgKR3Jkko+VzoHQCXrttRaWgZRatCLIUy36lnciCnVXC94wV2FH
DTjVhiwxoxPK/NqT1aigu1uzxH8j4bVYWqM0aHLr2W0ICv+ypdxtQ1pypE/9XrQG
qT8olcz0ixUSWhVQD0EAz1sq7kW70fDJPUNALlZHpZSNDaZqrDtnX1NlipUwrBpW
jA1MM5KyK0QKRH4TKgfFMyOoqpSypylnzkcw7uFV8kI0OSEZtgOxvZqaTtfSUv98
xptrS4oBvLwPcbK5dl4jzWpibLl/x2igPsmTz4uvzFdP4PbQuKPnYzeJTaKEEWlU
F0B5P8RpdZqSOAcfdzwLdgYZBH73R0ug2JRAcU49FvlqHV+hhSDdwL65Gr0xDLux
2oyGNoA36UDBFQ3ceFqtVtStGp6CZhVnF49xaTCmy9rbHXV4swVir8ZYrJNGjDkH
1NwLxfxEoSqdWf2oIDbyykS8Nf2QQrBCi+vQFRAKyGccvqENnBHMSvPyTZYzmuQS
eSV/JXJcNvpcUiwcMEHOVYIzM4WqfkZ5mX8hMVKRL5rlvztef4QTxrRvUUzkgFc9
wd+JV7V7g+Pdk0WXMUOSpdawyyLqAknLwMfrpCZUjO4oDHmHE9MFjs+RUvPkRscI
5LuOTunDhAJLJUToHkBdfd0qWQE4KvLZiD9YjTURTZVqWLh3lZV/Me6l78TcXJL4
+EXxrWAWlm3k+sESPS/EuzfJh8s0VDk6dBvrE54RBNJwO3nuWigAoBan8GLRIgYc
epTihVbWPBt4BBEQojm8XzgydKkAj6LwyxYA2g4qVWeUdjDG9khpZIcj2xz6g7dn
0GrNs3+3SFQhHR631XNZOZuN6e61i4/4Y7kpXovKMwXwmCN9oGZjA81TCsIhLpnP
UR9KB+DZjE+s+qsXyTjenHVt0H0nHgSy9y9QD2LmpoyHrhgp8IXMclwNr9Lfsyqp
BGT6OYVzFB13h8kWsJPv0baFbOJzUBEQtdPZ79smOLJbFS/ruRPSGzcX7nCCcpbb
378VMq//IzQ9CPQnonBJtkRknei7b8N+3ZPyiOctq340Tw2k7M3Q7wW2V8EEky2k
rFiZddrvYJWY8jKllfohX3jzajuClR11AhBYVszkcZ3fm6/qyzZ9bei4X2V/YNvc
B50WrvgMJCr9iksCLOoJ+uQksXA6WNj8heqqQbJWNIWmac+fiS/im8/xiGGaRHIN
AF6p/W24KxOeEqb/bCujGCSt3sItwrlb9tEXLTqef3IAo0ds7T+aj0HvjYFiPomy
gBdiFg1X9dv4jTG0b0vDJcT6aASDN2EgtXR4xpwIh40xqssHJ204KLKoysPwsSy/
Zxpqb78lobr1xG8vQe7/7gO7hpamLCmkeveng6SwX9GWr+/7kZvvqVUi38GfAG87
Yp3nhZlAh9hg9EvLn80OntAfOIcDC+1PcRjsUe9vVs3jY8aXuvUFdBMASKLH+EKH
4gATI7NwRtCNUmwc87i9/+BpUb5SCJlC5WojVHBJ79XlNrB+S5fKxVVARM9xZGbZ
V79W5gioYS8cwf4g6BjDvFY7iMKjfX/tEboVtu7dtqfXnGAdm+F9mQnizgiMbFPe
rHf1DCeNnRCPHYGElMNKeX1zykSpd1MTtTatpVzsM8XIDna4S09D1AfM2J6KAvCm
Gt+idD7M/buL+STqztrgGIT8XtbPFKUETpOSBsRhPa6fda6dHBRS/Rw4LT5Z/whB
IDMsILAkJB1U3R1syZk5GVSFMGoEE236gUBO3Q8DlT/JCMM8tymfNd9lgtCZVuqf
ieDN2xa766S9SRv34l4Z1FQiWVAU/lWW3mymSZSe+4Dkkq68AqCtaEEzNRit36lD
rJRCOR1GZsFSLSFULhtpSDXEPuuN9TbySi54eGYr3l6iP5spQCRcXWm3TqVgOCju
LY793aIuWQC99ivL6VuA2uxJtMXdNVxXoVLQWUAVc0AiXXVg5A3QAosDvwvoSEvw
i/0wtkLYdXfgwEnuTZ5OrDd1gJtSvCAiJgD56AcwXNyhqcvB79EJYeMUFHTUE7fO
WIjCQTDRa/WwdFYXwwQbrWgfK8i1CUbokJtT45jludtNKQLpnOVj130uLBw1T24V
SBUfGc2XNWyRV4kN60LqgHkVQ1oH1EZqrD6ZnswFOB4KF5mIKEPVhcCRiiqZQ9kb
KEQZZ6yXCfZla/M7Uc0YScVtWwWdc7Oc/4z3/WR2e/kQtjQSNTg2OqpK9kRplLjM
/J8Z72pxpJcr3qNq6wOP3mu5dCsG1dRje7/Xsy9piFNXPBc7ovyQjAgAHpkJcIxk
pu4LZucKCTghhKUEyznfitcU6VNFqgiuvZFHoSfmHyij5tpXD9BMv3mHwefLR5kC
4EnTxDJja0XLIj7wBcD18Ah46mwHCJEp5V8NJYsDpP0X3raoZxyqyoLLHUBZ7isR
mvqf/y+7Uf2wzWne+6kjLsh+fZv8fw9N0lrF4ovePz5VjVznO1h022JxFJ0hClWg
XEXeb4scnrx4cNumB+QDqQ326flEu+yLz4gCl9lyWv+fVSO8fHmTrh/87Bt0SMnx
UcR510UG34Gxf4w5FPzK9dXbA55g4nKrOnsE5khmi8KHzgDRmdo+F68sXYSphend
Dhq8IUNQLO/GXWZ6T7pxprxuwnDQhIHE9tm14SQ/khTvjpIFsvikkZskXh8E8+EI
3JxOdWl9ZoUctQzMwLLe4C0cxtagidxNmpFG28nD1aVRqfcagOTheMFicAN7t8Ov
0DNHarOPivcKerDogTJzDIBbIe8TklxHj6/wd65posWqQ4z8PbJTeoT+TeuAE4e5
5zRi1IZAT2xb4fIgDHhZa1YS+9oHHK3WotliZ3AHwXT0rwetgdYl5+pzRawQHjk6
V9cziqpW2fxhqkXUR6Kk0XMTu+arefRmXCXe/Wvgbn1ksdzW6QxDnMZGr2bx6TQK
enfkRKNIJzL7dp0d5aGMD7p7Q00R1DFOqKANvJ4xrRLCKn8w61Iqc+8oZOPRoDHA
NgBRyTGF3KeL4epte8aB82CIFZp5d/Mw0QbW8exClkJV/o5pt4Xwt1kKr8O//M9u
09LxysEaqU85uAQqaSS+zLpep9Dtl6J2FdNxf2/Os9P7rrZB7IY5XLGMj0FW6Wk0
agJmpmypGG89fENREyYF/+67YurFWGPwBGJ9CwSsiH8VxgxdMyCPKCUD0O9NbjBC
2pQ/qaRZURx4oKSHlblM/Gm8ZJOAhJgXhDdBY+pa2iUUh8mmFDF6UYJcNn9fEA5T
lMI+A6wAU3jFXMArF4N93ggnME1j1D0QTHBsA+1tMGPrEblXGR3MRa/r4Mfcg5AX
wQn30vx+2AUiq7ia5+JWYTJXWqTEljtq1lprSthLVeSLmbx/WqvkFLGRK+2FIn9t
33xnbd6HjEUrpF007TKXN8PE8VcO1Xb02PynbwwPKJw9Dqr9CT4lOt15kZDIcLvI
qa6RDrYY+2qLWkG5Sd0NrM3Yp8DpFM7vSh6cWoJHjpFvN0xfjmalZvwzVDW6Uoth
5Sgzg5WggW0akw+zcWC9rgO1vBiIpOZtlyiA3y88xry1fQNN8An3fiJ3TpaoGHOH
9rFcEwyxhOcDpYCO0Q7mJ0HWD0rr7vR9nZ9Odr+4IPkBzjOk4KTkFg8DAcLAPPvv
Hfcl63kv2l9eFbg2WYwWbavkBjJjQAz8a+C+BLMfiO8kaoRWe3gzVjTX/ID23Efw
sRRRWCkSZvf8tPYFLftXWK4jbYMSqAmzQPhFtrkhrQrABbAA2L8nBzA3unVEdqiS
pEuOZTP9Rwd5oUmo+8UeLkSC5UQcPHnKr7P7PH+u6vkf1gAL8GndV5qx1FQ3Y1Tm
kuIFTYQy0VN/5+f54Cev3PThse0jY94mI3EhlwJy3YeryhZaiG4V28MiiNbEX8ew
kJ6rsAo0SARK3FEJrS/YqWGFpb+2VJQ4IfWchwYL+10Gk+rmUsmS5NHfccEHOZTy
Ja2EgmxtN93LKeKOtPOqMptK5g8FUAAIA+63ZFzsF6URkJ24qFzB4Tfsoo7XpB7a
VHTvIXIFFrCvZPAoQ989ReGRbTXM7cZS65ZfO2zLVmMAdVsiP0Ol1ZkmOaoa352a
mboqhYIzd76wH16XvqL6Alf7Golj3/tmaOCtzDL4o6FP0D2Yk7Yn8FYkcVrLKrik
vIElWjJ6f2AUriohz4CkEOvdaGNvzqyDATuFVrfPVEA6erZK9kH1vlTDwP+cMGN5
qV1qaAzavAuWSmXQ72hs8p/gPhz2XUaUIRiW+nPUAIY5him9dCY/RwJp7L9gzz9J
ws3lhcmTGyFYUC3EGGO/BEKx/G2wLubJvyuves248cncttWC4xPvJTakN9Z7vo6g
lukC+i4m3D3pJC86+XiVOCp/hHvR8jf3D2c4B3KqhP0vsjwSXQ4IIxyDh1P/fyTb
ig8YXtXzX4PcPcjF+Q46wFYPrBJyZxTezGysXuGZa01N/mi2B3vPjhXhWbG1xrf6
FqcygcBCTcvZ5MhpyLL8tiUDbg7QpaucNCIqCSfROxLW6pOV5eUTk0KqlGs0lSjP
KJOqZiBxKsndQtJQ7dsUgnva4kNqnYxmtMxc4ZAIaJ8E8YPxlsFY+aTUBUl9MgEJ
nnKYKFMJtQgaF2am8xFFVmqCf8WM8xe0Df3f2despI1OmQ0A1J+pYBJrtIUKH+iR
XAU3tPmiEmdcitDFXcwbTBAGLUW1nX0BW4ZEbcaQWbvaQHUAakoSu3pQRIA3//SZ
r+sAkPdtTVMTz4WN6pne9ZtJfA4L9+v5HLfTJagav/by61ZSAUHNhkeJhDOjxPWA
vXBgboa/3XDzU0YQvft50eem0a3eqMBs04FPH1fl6Ol+sS9/Y0JoiUBWqKO76d0l
nx1JUF7mE2HxNJM+XNwf/47EzQE49p1pkW3xbclP1OTg5Uv3+DJE1WTQkN9kGwwD
My95rq8OS9MTtYjzrhdQM/Nv0S99H7nWlRDa/ELYxS6M2hLmIeO2pSP5SWJFMzDG
HQx8SdbN5uNuTIxEfMQj6PhrjDCGz4Ty12vGjH57Aa35IjGDUSeeiTaIF6+FsQ0c
MwnK8qAnl2tcjCr4PRYg83+aFVlT+VRBbflvXplLq714zv1eiFswPQdEbockdP8r
UYHrBGFqH0cZElMjgJ/2CjN/Aaj+dawKmbC05Ek9uO/uRGoWtOVB4HDu9iR/0xmo
FV6Ulec8CRSzX4/NoLJLvL31la75pAkZKG/lhxrNHBSSDMaWbmfKZPoppcAiCGjP
6lKSZtjj0otN1694ds4SSOB5uRuVzr6ZKaOUSN9li9ET1DMUkuONWbzI9egvw4nU
4aEPgBUtllQ/G449J9FuCZTB0UVfMfTXKZAK6iq7szSqUZj1d3MfYoM9eJWRviKQ
zRxUSYl7ucDPlC9dT1l+iuCMK669TzkM4+o0B1gcTxrViGBfEIydZQiFcShVZ2wL
91UcMqORq5+0GUadGuK9hzVv6vSilYg0ewIRFXLGq/oRBkg9Hc1BvRvec6IhiyCE
Dqyk6p8aF02Tca5OTxBVC1cFckwn30M0Jr1PUCQgNtRvPcJAUhT2nOlXEP2AXpdm
GCJmLK0Dmlqarfd7g5yKnhk82jqe0IeAywM6KrzO0P9qkAkBvalC3qZmw6F+gZxY
F4qCBP+tE2iovSvJkpCGed9UK50aMSMPXAvTeUMCIXztKDKwb2colDfANVbEOwI/
Tw2qiw7GBrn9iYNpXfhehXpU8X+htobdTm3W+iY6DfsnsHpPGJzmVXsjNCSo1yTv
AhkWhbLzXG5u8wWEX4w82GAcFsVdqtIRYuSHr0g+TR83WPxbWYB+BnhlpUBqYeGk
ETm3vLf4f4gwR8t5QkX1A2f9uq2I0l6y39323Hm6PghMZgqbDNj8ZeCok8RzKIh8
WFVQnP0KCuiYGDVhHO9ItZh3Y4fi59v5pJzcUOrMkBxKqJKZtXDQUOrcBu1Zu5hT
B2M3e9tg1miwgyKKd5FRYT9xfxh2xK0so16xJkYbsV4kszxC+RV5KI34uR3vobAS
iS5D2pjP2Nz496PzJX3jQ4kBYh6Yzz3E1XlrKOF9tBGiz37SIiiBCSeC5Kl27GO7
TyU/EfcCgFesqfN8xY8j3adDb9cmk9AfnSnve9PX8QthFrHjWBLF39VwDXIX1p/a
1lYg0hZ97NmbK1dmh3Fm5fbOvfdYabt2LauyfNjlDU3+ktNI3QkVrnnWLGeUt5CL
QGvfO/6Hc2HpSS8ug/h/2T1XItKw2nROoHOswRuRhxM4x6WEFtKc3PYp2AQ2czLI
EB1A+q50k77QTxYpR701u8NY9wuCTgRwhEr7b1rjb0/UtmVlTnAg9tgD0XftVQzC
oZDcAoNcH5HV06SE9B8J9eE94oJSfg3O7oyY6mv65UEqcaCUnV8cwwAylMRUCqUJ
fAORG44VPwwWMX7Tl5p8Do//eY2RzeY/QQp0tYetAUEyhzmCi7AAGxzWj3MqLJl1
WHTmytPmqn/cqUlhjPiDh3ipgPjBDOVMnDxJZkXsGswKWVOL4JMnpFDc9Szr/zEZ
mCcR3+JlnIS1bUUhqJb2ojltWI9lolbTLyrFb8AsFAg3Zh2pDKD4f0XEa4I+QrCv
2r9gQbwqYSP6gdVsPy0J26suJZTlHZtiBzN6ylpqk+q7si+6Ie9NFgjndl9cv7m0
Rex6oCm5HFW5nuZtSdEreSPRJnMEXKX6M3xiAm3cQqtvBJSUcpRrrrD+Q9zPV9bG
SamlQkIOWrh0IrF+hgu69TTA0AwKr12ujcA5EXhV6y6WQE81qUfdZjJ6PoByh03m
UbveNIy3noLG6BKbRjN+Zzy/yX15QDQu9LfNUc8sZuXzK2QAhTW6inQ8D6z8UA7X
PMb0BOUcGhxi5qDLiuTlrw/PpzpXaQOeyMuSwb4YV4vWt/iLUjUe4//2j2WteUOB
DM1jCxVc+zT+vwyfQYBtuJ5p85DOLxyZKK1qznlTJoCYzwtCdVcnF45F73OYpFHo
+GHJkeVy9rELSNREIniZMFZbFSRpBHdBHx56nJyHp2VbqIQPO4pkrkT5hviffVSU
Y2UNH2XS5RtHfnR4x6VV3v0SZbuNNDbnm/cU8DXwY+tzZkxwWoz4fSWaIr0NFg8U
W/L7JU7Xt2Urx+yokBV0Dru6ZxM/dc4+pY0IFVWm0AIknD/13PHCoHxfxcnI24+U
eJJrcDXYkfdNk5FgqtHOTskQ/oMH5ITGGVstdujUliKAxOYzSwOnnbxZzGxAf0wq
iIote8e9//oaStBlTuiLS3Uj96OxHXn44rLwM3KQluAk7rFZNyl8p8097njkf+MZ
3JY4f7u3OEAnbOoPxy2IwgEMV3smzlwITR4iGkpA0yUlKHyU6xP/F+ul/E0I16QK
jUvzR6NYvS2cyMxr9RWtNvh4CIMixLqZMxmwtzj6JiY7BM0RXD5mn4eWYZfMRRa4
grl8n3f1h4VzEdvqOAP1jUmlDyTR3zIraAoaA1F3u7s1xM3bgjmzyHU/nj6BPt5J
vb6cN2aeaN5fsfQoEoKisBlDzzbgJdrifEOGtncVjScBw4/QspzIn7eR9S2OuZzv
tCAljIKE0eTZ524wl6RpXyzq2XLq+4ciHMKkeDH9JrmyS7HKAM7C1X8hS03/lZgC
iY/2lm9rgyZwYeRLrVvshtr93J08X1lmxk4+UZhfeJunVd2MCbZwOQszi0BR+7K7
waf+QhLP+WkSLqKcvFNYCFGHoZhHw7BYLHnGY/Jk7kUUHrZXIoGSpM6IKQKSJv/J
5owBPYcYoUt9uKc0UbihhRrydXwSKrDOFHYo5PHUghfcssa5tlXsrZxZ1GMV3s/4
G+xgzThZMx9xruQx/w56LmHKn3G9Yqjjpr56ve0nqd7QEBruRgPbcIS8f+ow/xuJ
p/Wder7eCuu9JyyhJRN9IEMnDIArLdYoxFua714k04wrxz8TtZr5po8M2gbNm+Aa
Q6uhTqh/+7ORRGpCFIYtnk+dAkieh9geSNw8NKJIigcfA2Rni/k7tX4KIKWns2Rq
yzE8Y15/Ix9/YQJ5Dy/6GqHYwLD4H/ImkDte/erVVGSJ418eq62uSV4Y5h6TB2ZE
QRmUxay5QdpCSXnfbVjW20RDj0N2w9G6Adch/UCka/wxPDwsKfsxXUIhTV6I2rYb
IGHu2AUEnyuD2DfEBO4w/FLfk1dx5vY0SvROu10ppBMLXLSETLliybjabQFg7+5Q
I72ztGDlg2clHKGzAL2Uy/GM3grZkLutOjzZHAvnNUXE0bY0mqLcEAY0p+Y1c08/
GG31uaq9Uvb1yqUH+kX/yoZMH0yzfcLj8Yxk6zqD10qvpDjZUFoDGJec61nufBW/
woTPlcITr8usnt6TuBkxKtbVCKlqu8ST6baMySCTfpOHKCeAGDRxn7CKMynNp4F3
qkFCJHNoJAURb5tZ4wf6OE+JVrkq4AONzjMmzimsTOx7XryJCaJRCcqE9SAnTrRo
SnGtz5w5xvIrn41j3oV93KRHuv9YZdJXyLULHE1Ro8ybBKsgMkSAvnuu0XZLf7Jj
gpeIRvMwkuyxXnjbnvIGNo1PKE23CkVa1km1Yx6r3ETwfGH+2DTvlnj8DUFYKMHn
3bjiqqQ3CAULlqrnP+dpIYu91CcrsoUGyE8GkuEJe4Q09gjn42ntH1pIeYMTq3ip
0cg0pjPaSD/VTAW7HUaDvnm4VYSQXl0CUZ+3ikonFDuu0Wmx8ZiolNndI1sPn0lw
jlf7Tw1qkjYfTJIiQgTBqQ+QmjiYuKjxOHEinOgbfb8921a6imNApt9J1rXfCO69
0mxM5447+GDAvOq7p4iopfIy4k8KAQZ9fGxjO2bokC/+9lgrpksNsQ7913Uzhie9
0WmYQuQgrq+WAt6M4pwKycpoVqXEgtFqPjxUrOlHTafRXsbQDyemFghVYyIOzJ/g
8kCzO/gBTsGBxfgiyMV2wwOacjd+dY7ZkbplLqOLtXz9bRWtI1Fx1q5Ts+maN5PB
LJYUc2GGxrSVORtJq4CZ0EUuzhhgxCu4KPlYAZLcZJa6Kf6Ge0osy4GMAcIyAaqw
ih+DKZlbrUi0r9XiiHZ+kTr76J6ijSV3tvad5ntn+hfZ+Tnnf8cTb5zusylB2OD/
/Bj5zaJ+yBz+LbrOiVTRBNMLrzGBXxM4hb33WCu7dXcvfhCSSvmLhaeijTP1La0K
Ppdal9S8xXq6rB/fhr0HWMsRSVgOxAHMg+9ft9vLS3J2j29DoF3THdmeypLOGhbY
E47ZeCoQQMPELiG7d96tvQGmgub7LgWEMkqfolwltXXN8DcNr/P1X2B0eSjNQHfc
jOewlvkOgki+7cV98yJekN3TUh64BUN9hfYZCgBaIQE8v6+QBMwTQwtirDEOxHIy
ooEiI56XXjzpy11xavsgGjuoR046mgzQ1C/NJdrIWhFW7ZY84PtKJr64oNvdgMdh
U0JImKImDyFxPtcsMeBViZIYmLxVp8LMTlqIW5AXT8T1jENUJ+NsmV7BQCIUKn+F
iWl6rEVNPrdmM23DGyHiUMlQQaV/rIGqOf7OVjeuIY0rCJCcQ3cVIVC/jn0KwdM2
tp5BRj3P4GN1MPb/lFmH/G14NCvzE01a3k+CRqvrse20izBmHj2amWBFzoOyaT12
RNU2ntpXSPYf1LxAzX/Vv87So87k2Yw8kaAqnOIXGKIWNzXX43YNF+Uw84npxouo
xgiw6JjeRvzbaOnzfUX9KWQVCsdZK0ZEDpbtmMc5zTzztOZmW3mdRxexxomO+sVc
fPcj6dspAClkO0X38PV7Kkt85FJVvvDc6XkuoJMK+xenvkE7ZOxIfmhwLLB5Hmjx
vgkFytt6juBs0fj5Cmu6gmkCHikZi41ConNJvXpF6jIICH4BbfdnDSAicjTcwizQ
a4ga7SQ3/XBXa983pPNqSIhnGN+Q5jMVDe7TFEgDehCXtvwVLKy1ne7G/rlxFeni
7kip0uUo/w9VVPzwZQVfoS93xyuVF+p8JoP+38H/G97pf8t3sC+jmbZlStsgtWHu
GPIb5NNTUZ17iObJffGqSgNEdHLPo7cX05Py9wVr3hFAEGHedZ9/WtCf69m1A2Mk
P6H2HppADHjKaKW4a+jpWDF28DV9wtTJydstsgXGzbm7IIQ+t9rrM5RTDUXJ9tMh
euVUg05LTcddOqlPFyMfDiIKdnVZ1Zyob5Dz+XF811W0x62KHVfaCx+zVdVQz/GV
nTYZHRA+PuVxbmruay6BFgLg6oif/jbsp9XzEq8gdhFxraW/mW8f84FJC1D9BbcT
jBg//DUS0KRqS9SWJq4WfnKU8XzuXjhVLshaaIci/NVcNAvAqsJSKbHtdw+BOJsm
hO5d/lKpECXIvuc8ElQpiQx92T8UoP4nuzET0nSNb6Ffz4UdkyiQOF+6+hVy/E8B
+cJFgjEmYNyAyPo6XcGztRJmGf/9vTMj5RtG/XhLFwTdDiDNVXzDZJjXwWU3kfjZ
C3wOoKx9ibcl5D/GkDljPkbQIs/5Huutsc/3utAxeZ51WWjyt4flF4K99/o+sdbS
FSxiCA+Lqb5UNSI5XYc/wKDVSBAkliLJOhTVHm5F23Kh063zF7Dt5EDS+umdiMBF
UGHVcQ9L5B7CAopvnUlwJUUudacbK6IlpjSCjraXibr1MgRlxSPGTNBIe7imFl8Z
lEX0802C3giSW6v0wRkzrXNukrSDputpRe5S4H4/i6ILQGf10GXICVONE7ENVckp
S87njPFlixvZKJW/JzzI/DhRKK+rz+vI9XB3zhaBKNl+71rgleB7U1B9ZNQOvddi
XKOZCNyrKV/Y7jHwu10A1vjE2su+hYAZ3bt+Hf4beKC8ezqdqyzSv7QjeJuS94mM
bO5nNIPZEC5lfX9n9PyD7A0DXUlN2hZpsJ9UNqeQAhuprE+ue1mBmTsPxX09Af6t
JFCafgceWOk/+wedqlQYPaGBWmS0odt+lbueUbkayJOjDBBjlFj/lY39HqLaKvai
rOvHKwELyz/jBFRfjhWG6PwXGwgrXNtZOWbkjxoC3Fxnx/ShG0EENfpMbucat2/L
wI30ZJn5q47pxyj+PJwLHWKdV48rUBsY7I7uB488IO2nG3Who+v+x9mmvDqT8s20
+KX/1yhA2gd0hY7nVVevyTvpfMEf8d+8CjMR53jhfm1kppiwmcXfG7mvbltqP5nj
Sg2xuydIIf0GZkFZ5u0djTslTSj4Mks+FWKORwarIem4ZVSflrbJYRbgyVcy7SlS
3FQy1nruB0RniN7SYDq0pEkaKJu9lCXLSYNXNNUekhLeBnKM85SFpUv++rhCR0HA
yIIALumiMseJXy7hQvpTyBN0h4b8iymazrDO4+pTo64hRO8FKNZu6mp0R9okpvJJ
YuqN4X8m5FX7QEiELa32eZ9CMaTmDHGrPpeokfyuOKZtmFPBHBh5VZSB1VRmzcwW
VNoi+hrxYuh0B1cMMkB1+xDAyTHOusX6Joi7Tfe05ca8bQrBUmBVwapil4BnrsmH
j0P1eDwnGYbE58yxGLv+4nnSZSyRFiDSiNkKrOwZG2kDSNd+x8C6AMLyWsT/iDxz
7/jzF3cpC2Q8BoGYuPhFUhhm7TsYZ4PZ/nEId7h2jrcUqCc2IQbkFxIrErNs7SzD
GkmJsrQ18cxqtg8yLnyz5W3NJRQf/S3fo7s9tywD34hzE0ObCGpmQLjRJ+y7+Csm
jglxnpzNms82IZT45cxMRUooXniq8jcj43OnXRS/F+3cJhc2W9yMhJeEbs0iv8kx
GEPp2CJalljhO8fnZbad1CpNtLTyY49jAtsUIe5tw3ho17thw/BnQaLAqi8o539N
0UlMDP0zYE4g8+amQYIYwpOdwiuP95bpJQ4ZxkfpXth44e6ApIiCV5zZfl/9vd+9
VbxKb6g6km8HlbSAe/chIK+RwAloeRoGSAvQ0wcj97QzcCrbbDGHdR6a93rbiwo8
uzI5oF49a3k2x7C64hO8oHT8lnamdvBcLt4x4X+LCvnrlWlJkbEd455xsQ/+rVYF
NnZEyZaXxHAYgtIRIYyXr4dRqpm8H2yket8pvYdvBnI7GKWoE6WOdlXJMsnfebmV
tOVKJxfEhUkGXjYi8EJVZMKHPIez/yR/ZTk8Cu3l78JApG9RIboyavZlbsOnqPWj
Y2UJZUaSiRIoy6inE7MBG52wTTHoiVd90anDgQ0glgumOBy9IHtJ4kg7Q1uaQFlD
XrKUsDOZQ84JF+lHctLCJMVZJnzrtbGWs/+SknhsqWjqK2fJLh2K8j2yLlkj0Few
9XSHXd5EEHsqPoulFHqB8HOmFKhpj1dQmkzRGlczRV90ulMT06+MuL1t7Xwz+68c
1tXzpoK0lKjjiDpN0fu8piJ46kE10A1EV33uLdQwET1rHzVJf9NTOx3CFvTMcpOJ
rL04YfntjHYF8fOa0oakPTF0g6xIOUkZWiiWHHMWg6EmOQno3Nw32fq1jfb2IggZ
L58YBQoxqkpUheL6yp9ACSHDvw/VyDa8FSO5rm2m6px6x+/3lYHE+LkR/iekErSW
F9xOU9JrBHs0pYFxELiEXMVfX3DzF5hf0qM9LZXGvQPITze4wkeLijhe12xXxVCI
mTE30FlglbwMUyg0JLtlwEcp719GLOa4233J5F71R64aiAvxpPCveAUCSFileic4
QnBdplnGoQwZ3I22cfowUtMTXictsfTrNml5Y+7DBTavdm33Lf1U6bJ4Q3kwbb8J
m5hJo3uI0DzB2O8T8q+jYNDze+icMdvf0kqLQgaZwOUqj5pM7TcT8qaVID3dR6OS
KTSKGQh3GHx/xVsyavDHQMy0d/mEL11OXttT18b9mFbpTn+jPDeGET9KmV5BGKRl
HYcfT6qTemgwIhBgnZ41bh0Mvw9t31nzgi5VhIr4e7vQItlZwTcnhESRnhr8nE30
feDFU/ADJuKIdtCb0WkydE1IHB4ZjIQRWnwxyhuljBinzUEtB8+T+IIOBjeFt72m
Y0piZWko6Y5q1mx6F/B2qfk47HAdLU7wnwC9URHXkeJym2IPUtD11OZEVPKjnrsP
N3i8K76+O4sZibSaMp1NVSgqPBgqTP38Bik9FpwLHHXKvnVFrGoebxI3cp7bjK/T
BBoXi134NwR+zeQMvxplPlWRt2k+6ob4nKdqgPoN6u3mtekE9+rN26mQ5VwwxANM
cpvHqqpQS6EBX/BvyxvSCl6UlwCgiN/yTPcdOXLI76hJ+1HPXc9nAlZKnC+J2q/4
sc60dU4sznkXrjiQsujoSt2hYSfxoAvHMblggHRikSqKzvYOioTABTfk08y8Rsz5
XOYKZeyJMUGqPVPYYrM7hUzv6jJnIzwk2zuJpXYsnvGBN92g/a7zx5IbSN7DcoTV
2WFRZ897V9TXQum9qgPtr1zLh/lTn7DB4NK+kt2r0jv9bQmTP/KcrwYn6VGPJ9cJ
Qpt2NrOR+cjZ/iXguJkNBImqQgmqQ609Ct7oqXXnI+IDWgiLYEjT54B+YS5Fp4M/
l0nUyTwawYSblqUZ3C7LOqVFa1WWmUEGxBYUBgH6sfCdSWKN9wI2ivDoB11ShN2B
b6N7xdaHPdzZhTtUKlM6j8V5yWnTzv+7betyRNEllGgs3ENubt/8j2/assJreUFq
sacsEz8zW+k9kt6uB59vT/l+GxfrRFVUXvYwGbOmdT5QnUut8m24W34l6PGKyl6L
BrdUJTa5fzVHPFbKz+7dsbV4Uy7JrJ7auAxrjJC9mGvLR+/Q7pUO8qEsj0Bv21Tc
6wd1Eky3xBjNAn43HmCgs4koJH61IDvB9vmLk0EqstazL6ZIz3kCyM5q2RILVobB
DmPARFj1KsAmerGZXF75hZUBfpZ6vwl6n9z9A9dEEffJTO/qGZqmI5DDoQZiZFeM
HrM40UWLsOG2x/+v1+PAe5VbDsqetyHsec/9/CPuMAou6MHprkHHEahA2qsLc/fG
oeic4lt8Gw+BFshL10/0ZB0zYVSLAIg7zIabJIgqAiPa7GnGk1q5cKTQ1Bon8jla
2CtRqxciyrriONsNsJ4P/vxEwOEh/ZU77sMLOcnMunwZYRP0z1yoDWh9oA/sCOxa
8Eeox1UlY5KQiQ8Zr28/vm/Il86cMNKie5TbRR6zyd8ulfowxGuzUAhk720ECqFr
Q3f7L419FmEBxTOaEV55VnqEQvJR0mHvujcfGPbbZlMoVn1x2sPRRQYwhTBKW3eW
lKONfB4FaTuaT1gmWpJnUE9u15p5J1+2vEXUzVq9mP0IneR3P8ypinijaeTH2cUD
ylHatJrLvdtM6dTinD3icRGtwMkO3/XXcd8ArvAL7nsiZ97i5M3YIv3waZ/VCnOA
SpsncJ62XEXAIWvKjG7UPVanV3QnxdsXekUWmfDcexMR2w4RD6ezSYsCEeXyklII
bx+bTAFXZrIxHwOccPntXBtF1Rbd6tYyuiTwGXVwl9mt+eTAvktmtY2+v6dovnde
OesbPj400QJiFT7cwpkcrFwI7gQFl5WctSSJapshg9mekLYOBb5A2FfrE+G0GKG1
F7+1jL0qavRjdzxjHUUFw/PSBmf/EoMZt7MrO5piBftDWn1jOvm/U8dfiXBZk9Qc
O+nc8s5sYG8VebaqLBznYad9fttoJjf3UWp1RRyJ8hDmrF5WmMU8U6We/q4psKst
SvPY9nExoS0UcwLuT77w4wsuJDuckSwaLBYWU5IHroDJ1FkOza8cO2+igC5ZtS8f
F+uAf8ZaSkFmE/BKtC0Gp3vK7gLcrzNAuaDaJ/FgKsph1vZqIZpVjuzncCrdI62F
5rrS77iB7dDXrOBz5ArB62ryweLXDetlBC8asyzi5fB6Ce2VALunNmxAobPC81sU
9B2OdCKqrvSpyTciOkOQq3x+5Kq+GoP61C3lSbLGF75vSSWUFC0V31B73OZnDHlh
L92bBtKKTLFZYaBAd8vHiMATvBrWNNTlFXRxvV/lOFQ5LbWmCOJx1uB4HX65eKGm
fgkQDTs5SjkL1dzdkhMzLonIvtRYsAJKTfT7DsUPFDjlr1CY6jsNYvv8iMm3NqXQ
3aPio9vBWRVWwANQl1xQhTiU0sf84NHl9sAmC2wrq1R4FxNoYa02pnm1DbBLSQhG
zFDqWr9sIBMs/Zu2ILTy4retOigaDDORyi8thSOp10HyfrLrxGQ4DS/9F2tIZmuc
6lM5sEuHSeWf0ehsavdHSCQqkAlBJN/ul7rO5wEGZ19TFly0dn23zSgarr3EXjH2
mAp4Ijo1au6fonasnKoP/7kuaiDuvRdwZWbEq9Dxrx93HlkvBj2eNrdV2L8E2/6b
UqiQa+fCgz+2j6xs4PjXsHXruBT04OZl8QYmphXyTr3TsEW0hDpX8R5z2nn7Sdci
lIhZco4wEPVdxsNT5YLG/bWV1H9+s41TuOfgZ4GyOqpYtoaI6/TIEbnNw8LKq6rM
3uhLWkqtNKE/dVCT4Ufc6HaihQCz7zcsUGyr3CY+Y3HUoDDwmJdlOI7S/Z1I1yh0
5xa3StzHTZGRfLuYNbad3ajeV+xdiGnux27npwGMCzWWjuOGLl99uqUKbpti65rr
CgqkafTcQ0pEMW0m3RmzxqPU9eTvhTSN+gDI0JE3ze4DllbOSk1bHt2kS6HpBYIT
ycNsWw/3zVJWnUvC9vLdimdcmVuB23OFJrWBKxcdI7tRPL4cYFE4vSeOISuVSGNc
vAN9lOsk2tI3gOC69y4po+SwhHA41rHQFWLsYEFRShgGKPrsjwdEuXql/XmDE4KW
EAaILDKGzg4lPlKiEOB6IaUPsPC0wH/awBlZsJpRb03m42x3LTekJoSp6viuV5nn
DsLi1lSafZp3dzjB91oiwRvkrBtd7MwxsDQuS7YWP4UipZJs5KTo/9ONZ/0uR/c7
mbsxGtUApzC+pZHVuqvrc52z7AfQyimX+/hyZUoyhjb92fDdla8WTC1p954FkV/f
bXm2aRpUnLPSUKn37r+wcrMgqr+deqD1Qi+mh2GrEXd1zLVK3QzlBcWmRgnHr0iO
gm3YdSdQOG1b9sXqmxPX9Nnu6rt499RtKmpEtpHXYV9ub8PTf8ljTDlmxbvwIbiJ
rq+uV9JDtrtNacHHUwHeNzVHwvmgmNROYs3YPNCvUhcFSGf7TSGGk5NuzaWas+jh
Lmh+oAsjiLx3rT+MsF5sV8uLqYl9RWaRAZyhvRrw4Wtra10i4FhelD3JacPj1zOa
3h2W6Diyz7qzpRWVH4OeMIskBPajtgv+3KCYCQH96VAP0cx5mugynhIkohPPEjpO
odOU43jwXJUnN64I0vLT8XN4OsiEs/NTwkj/2qEevaYjbu0XnFWpa2yLoGN+Ecvu
tI118vgjjE2GMVMu5ESqk0OeRbaBqt3k0ERxxpljFeinS4pY1SgMBApGsJICuevj
tazYHvBT3KQGR1/JhIXXoEKXZnXedFvW6932E9KVtGKsld/A8jjt7XtmGcUMP0L4
o2dZ/IoWi3VMxCGyj4E6+7KBcFkTSDRkP4wpW/4tW99I79606SgpUjTblttDCsvA
rIugDjUTmdeLnfDq1GkDOU2x/i6nyYut0ANXpyENVzHkLTGPu45mT7VThICntNfk
wTlOjETjb4F16/ggvTQs+fi5JTrHOng9XokEz9Y8yoWrknFpRR6QgzTNJsqPzWhk
5e6vYCy4IhaX65mmq2NMBVd7U776KfgKZDHjNrQ1M5wTR6iCQnZtRAawhxe6JZWc
+Tf0jn07Cw+ttH5kH8gxrQQ/RH2CUuW6KmmMWyM8Lgj/Yp5HWjwyjGaNGBvkofdF
fU9broHSJ0vF6+ixk7Nk84kiaA8Ebeg45+LBxvsgQFaJEwTWCq9us+QrEr7WB8bL
F9wMQAia3u7fFVQz1TxgJed2MlVKd5KmMY4myG0ECIIgsZzYMHzke0B+UtQSoXDB
zD1RkymLQlwdAdvUy/73ux+mn7pQWcW4MppCN8kPqiCLVwL8k/V8j/mgZPY7v8ks
MHo43LTgQh47ErqZIgf1+Dly4y8MrE/scXrzQfARcIBqv1rreEJu0GSBkrGmkF5W
/MWHTDsn8hq72I3NzBxO+7p49ryOy9W9yOvvf5pBwWLX6dhsxS/E6juJXb7UK4gb
/9mOMRDJHybtjVPF+ELkESB9+Lf+IxwfmnvB0dAj3rNdojtJS0W2JYEP5px7/PQ7
Oys2aL4OrHYwrF3D+ZL7uOpVXNo8mkWl603M0yGjI3s9r+XsArepx6qAOTzYtjeS
s4FKMLg+hdaaTUIn9SjdlBVYkKacIWYJ959y+Xpcw2afBxUH0ywb3cqUCOhQ9RO5
m6SNvgDmMG2P//UiNgND4vl4DydJK6e9aVRDk5IoVz15UVSKHDgKNHRbVfJL+O6d
MUhEgy7Z6OX04XhaE0mq2JyS/WqCKjHY15DV+YF38l50xRW+uEI0HNnNHUfC15uP
JPCDEGRJ3DX76fLrJfyvmd4UE+JCzZnXx5i5S0F7aZ8hNsWsN0Loc028CAEYwPIp
yij5xo+PTN1bXYUOlT19siuy4LoW5zSHsTp/10Bvr9fuYK0YL10RDIO6Rx0CbHPP
gxPA5bXGw2RzKtbxkwiZmB/2Lj0hJCsoYe8L+9o5wAkE7x+N6YJDomaHIkOr5U4S
n+TfFVQUI1XMhq3XFiq0QU5qLaXNhsYTIrMt/vKhMjEe36ilB2W+0mFBhGCUUBqo
mdydU3+6M5rclgnJmkPJCFt+GolenedMm2cVQ5EHcK+B9ajzlW/Trr+fewdB4qph
ZwnbBYQ32kPWvqnHFvEuk9hbpMrES1Ga6gXUVPKzD+qQlGKIvicPEpep8BxUixKK
bRZUPqE/wzfDkGGe6xYtaPEvhrl/AF9iLPYUbUqrEJi91b9PuwUOkonryjbGf11Q
EELPRKKNDjeXvAkYPfqhd9TiaiMsOLqchb/U/NfQ/uwfinj0oOrdeDu9evdoHi2w
fPRfJZdHCcL/KQ4HcGPoPrfRby++4Sb111R/lYf1afYFn5sZ8fMpD0lq4halzJie
z7p/7EtZe6H6TMeF/oZdA33qsaRdoe7yim2XxeeBXyr8Q186S0StmsHPB1Sb8TGF
WXqb8ysTrqsfS+qC0/RdwGkM3IMTze6lQE7Oinl9n0V/J87Bofh+FTy/1aKh2Rbe
8ZrCcut8KlkRt1+N4ENwZ9yLM4zcChAViz9KnyRwuFFWMP6oMJftutKYBquhi3uU
pQ+8pXtF8CiGUydiTGtA8/3Nw4/ij7ngxe+3tZF66KjAHHEake+x2R61rKazWMl8
MuKfPZbQv0mslADJYpeS8muoToK2bmC/caHhyJsJVFqyKz1f5JTyYeOtXKAdl449
bx3TXaTR1QxSulqVIy12jIS34ozzk+yAyjF9k28qwD0qAv6Q8hFIgNUzZ63CI3We
1xo67xTXvBEB6tPBPBqIv0q5YosLXHqScBkNQonZT/uN5kmBqWfcJej13UCi6Emc
BiX7NkOHNLQ0mVV2zAzIrIi9YPTJquWhV9hM1bg7IunkJ+ilXYrjthLqDGCJ1TEB
3QmUk6HTN+oEH30ywr0Opb08/DvR8aVA3QmX0AxAbq6vrogCdUHP5ECJ13lL2pj7
zkdega8HysVfEMyLKPNSU6aULTbB4VKgEKmoJ/+pvyFFY+1dzr2MpfxuaYp/hCaO
9xJMlXmWznNbIBvJOvP/8dOG6PL+D6VcTNfZyhGjwUdHoRZI+8aTjrGGVzCqlVWj
LMDxwSpCTNPxlfYX5aCjgKM6OCrSRZbwzS30F5XpqN8CZ1Dfss5ZLkj+wia9s1+3
bEan7OC0bBXFgE4lcRm9b5x98xQ4F3RmxGI/gDK1tzWlmUgMZZGIprHyK2GeyFmp
YTRTSd61kAnq22xhku06GHJTtsNDLvsnKNm5cOBKZw60mWxmikK62bVtO9YYCOyG
ovsNq3DQXmGtenXTweeE2BMTQsDrIk74WvQeIGl/JpfB9cfoWjAoLCjLbn/uXFOS
NAjJqA3ucRDBtgxaOshgy2U7KmQDQJAWGPMUUg6Dfl4H89yIK41IafpEGX0mx9Ud
eRWIWOxcW/2J83IcM2CYLtRlPK2bUGQViu987CEcPJ5jkrkrf+j1m2IT0dyputUw
jb/rBmeVPCt5MT0XkjYSI7PDG/8km3rDI8bIT4Rjxw5sV29zW3PaI9Js8OjCRTiz
hYwtmj9m+ier26GjVsmACWp5/VzF0TZaWleriBfyI3e1wnSJDY/hcD5zsjBR3m3H
P6dcPy02wKqcOd2itxnIELhAc85bhUfuJcHLNzYmEV8BQBiAq7flO0TJk11O3VCI
WPlvZV7O6M0V3oEPoU6SkAgeiJPcf5Oy2NHgPXGhhujB6G0Kpkt3zbZ5vHnWzf2/
38OId6FaGAsOayUKB9ZGB5zF5GulLDPVrFnVPVgJFKT6oHR0blEBDBus/9hL1UcD
MBox18Fuzp1ZirQJQjhKwQBeUhJxF0yqdF2BcFv5Hn7UWMFO96kvOdHga0X4h932
+xXkNMvAG0AKgOOX38pCQr7Bvl3Kh1Tks8S7oXm5bgnFbvEDOSjk5EKT3gI++MAA
JgTpEQsma7VCzJgybaz7bohH+StpANqJvL2ZMPuTYOYoBhZdkL59qMapRToJFG8u
orKkLXbPeFwD+euVBLsZM8pKi0NnB1KejUQksfIwWn3rQqQJxZXVrWDI12EUXz2W
`protect END_PROTECTED
