`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ccC6DXkYi4y0h9NXwX+YJv3S4MNfZXmM8oz3D2vC3GMej2uElLGnBX/ySUFJ2kzM
RW+TFwILyg2O0wZxf07qqFUkedNO0HH6AkJULvWcMd/6j8f3rAJqhA7XbgmoVLbD
hsgJ3kzmgZDR5BeQ0zCrS7BPWInYwawbtsYbc+sKYsoiji8tRfJThish3LzBQujA
NZAd/O3pj8lO3U+d7fysuAOTirB7M080wdGobyyRUGpeNrjWkwWuvwKiFGVf0hAZ
IzCdmjaZ0cZZurpEa/u5WUPqelxxl5vswGy+7i6gF35CzmImCN6t0jmL+2Jp+MV2
BoKuhWqgj96qSo9JPB1kTLw0iqkxZhIDfUeUimCSqgSlwb9FJs8tCFyYk7AA1X3o
N/sI/XvHVuJAPCctPIplh7avdvZlLeWxSyf3nhxif23w/kz1qhuTzLoezV9Cp82H
jniX0KcUQQRDR9OUvXbkbMJQVoHK/NY/BwxqMcp3yzkTpurlC3l/JoT+lgQFD0AP
81120Ime5NX0WBc3nXZgiWDWfYEHa7UfraJyUKxWOsz7PqH8RSBrpCcRNkNh+tK0
a5EQ1bOEtyXxdTW51iP5B+ERBn6Cr7FMHEqryPLJpXvcf6PNKAR5PveI+AkfwnmI
Ez3Q7SXBhxbxQQT3B/sD1FLVKMF7K+g5TR5RbckKZnVQT+wMApKs0Lla9WCkGtTG
FxWgtWHUhFd1kZdsScEI0c2B+TcxAyTNnNvBhCpJ9CHAz7+FGJacujVo8/cPMWtZ
dv2ndwg8XF4jLT5KpD/1frWxmcdIqFH18CvZyeKdX/c=
`protect END_PROTECTED
