`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OCTNL9pdFj4znknDFIDfpuULjSXTefWC3r6LaoIl92LEP7DuPO476P1mxidLJtpa
C0BkZkqpWH6YFIbihKJgyUuA1vjfLqIcsKgrHB8dXkDdbckEDQDIxDUo6M04OC7l
iAhDo2vULmHqIWu1qZFUSLehCQxYMZM89V+f1WkvLSdOmVfd7yUia2/lzHQ2xZ5j
9QZz8SgZY7L8qFDkeLTt4tLtfSuWIwp0HBiRBT51aBChhEYpZSY3GpdF2aYm+d9D
bpV+TS02oMX4GKzWHSMtrncj+fhNPeswf0Mb0GbH9Cfb2OWaAhZCvor/ZZdTj/VX
cSHXEmp9osOUMr+WFIdySD+GO/TTpvXT8p1DQj1TgmkU9a9wWtRHNqNgGS/ByXWU
axfeV76iqQOlMaEaY9K3goE/Wy69OwIbtxHzmASvxE91ryC3EgYNLMZmxo9DekW5
4zfva9zNw32JkfduXm80kWOOt2pGqNwJeL8Bk9osEUEQkqokqTUJKcziQit9Hkvy
`protect END_PROTECTED
