`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IxTZgUe8USVXbr5IdWIKiqXXz/LSfc4f/BUCuXKblB8j+omINOJEXwjhta9fwCLr
P/AqP6yGOVj9cwfPcSkifO45yMCvcoQgsjm0JuL4xZxdaaet6czw6r4wrdU+BFNh
GZD9eLfjpzmkeUam9xekocxgk4g7zYBEBrpNAZfk0JZVtFgq8NgTUFt4n3RUXpd3
u5UaXQGQAAsaWVW+gX+XImGaUaunf/pdUn6DK9QfkhQGEul7QoXk1Ca8qcGy300I
HJ7ybaa50f3FbBfCHGngd+SJjUpn7evAyoecXNJ0PF88uIJBvhy4M27EJ+YjGpLb
TpCQPRL1dkbVVWqALNvQd/fjLAoTW74sgsmuZOhmVyOxcSvowpiJCroF/u5LhCPp
90EPQAK/XVO27uqCsIKKWNojH77uyxVuj92+4KHCzS5svzOih+ctcpgewMVtntCf
`protect END_PROTECTED
