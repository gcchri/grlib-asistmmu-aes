`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FjvPPjtYNigr2/8qebkNLGC8nIv6jin9+MyULG0PoGGOz/W50tbrAu0/aVi2xjZz
Aa15olSVSqN0ggWyXEEe/GQI2SdDETC7u53659TBFT21y/Bm+oZKUxQTrpGnNtv7
dM5uhiYdyTQcjGnf4L8umSZrliGSBY3TDoEQ42BoHei2i7CQOJNmWGtgOi0xUyBa
iHdi87iENRzlWBT5ECiArTtfWcC2gBnEeekqLAPRfO0LMzhxlNbrEZ1ubpTsGCkW
mndttIybGRdl3VofJmk/6EQ0T8cxHuOkTLXVHXpU4mTQLBwaJWt9lAewsaaQNE5o
c46gAUZM6e52uw54OhLNxQ==
`protect END_PROTECTED
