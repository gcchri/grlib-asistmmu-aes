`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3r+5o+PX0NB8znx+8I8cooRF5W0OJH3R5GyFnH3j4Os2u0QEq94Wy1Tx5kRwoX3W
ZyMXtTzRmbvHSX4f+hnAsXzXbrNMAHZAdtrzhpgtbZFyLEANOqqA/CacMXZqy51W
rNNfuftx5gxjP+XAyLCRoABDI7X4nr3xzSROWHprpkrRuEDcjYozyp4tDqnZHoBG
o14tbP+XXRy6yl6k9ie08ZYPfiBrxtiWDNTcEiGzor8rxsrGe9Qj1YNoupNf26FH
mYYwrMwJKhW5HB6FyQEM6i2HNYN0vDXp4ovSfLSHTEC1srwnO17+HJMZYIcalhYI
6Ye4kgZnC/eMDzJwoQn3a754SshWYapuf1HPLvPaKnHVx3/5JGCKDfWZBybhg2LH
KdVFNK6dP9zHzOtIzZphU3mlUB66nCgoyuf2ecHKz1g=
`protect END_PROTECTED
