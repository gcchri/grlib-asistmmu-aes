`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m3LW43sYCXFFRYiBjWR4n8LA9P1v5bO8+k+LA4VKulqd9Pqv6uwSdenkik0U/hkQ
rar+HDzCHGq2Mcihcm1yPFFpo9n9p+0vmayqKXhb6A9ee3CzAJSVmAUR7uDNloua
xXp3iTPQ5CDiSCSmFf3jeCdq+MjWKwpDD/YnRZ+BuPa4Cddg6oFtxLfvKvpL+YjW
XcPR/0XyS4NZlD3lkaP+TAaQm2ffKIuiT5ofZhxbGhja2mvecjzUPLQOMgsSNUTY
CJWhzPn6fpY7wvD9rPhq6hzVwEVHSuloe85tK0kdHl5ao1vx8dSNL7eheuR54Hbj
G0RU08axbGVywHbNHpHGwjFcprXREubIPgZGV5mkgUZSWmPCC+onFErQjwIgyeDR
1Mj8s8DTIG5kI9W5Dm4tduAxP9ySTgm3b6RanT26O20Sel4Y14U40CQwKNmjxkYQ
Jmqc9jGkSfTQ9E6ldF0fC42o7WT3qG7qfPfCl/Z6WHM=
`protect END_PROTECTED
