`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/tUFdCSb44WL5xdhqZfz50Gs9NBoPtIUxNuvb4MvMg6JlMFJ4sLb1NQ05P8npvXa
s1dk0ZAnCXC8sYSTu22T7bZpB0CMIYgwEBJ6Ei0qb8JjugIito3OkJba2Abaut9T
xdEvp1/HrJ45hi4uAJzM2xNZ6cjhsZ4VOwdoVO2ec18vrvXHE+M6gPViZWDLIfwj
PNa6cb2Y2PO9enTLcfwwabRKbqmkdXl0OnvKztSdq2fYvAutnU2gZG/LegvF1ps3
28QKQQedOa+/56X978Op+uZPATLvLbjrsallMab7Qcm99NWq651z1hG1AMML0fsV
9zoQBoJdLDKFS0K5zZ4mQHnkLnnp38VY4h6h/ThkLtfg0bp8m6yUPcA/mNM0y9Ix
HndktUVjVZG93AzvNByysGRs0S9P6fFTzOFL0zzVwsRhC0E2bJfJ0EqhD8Z0xpq3
qW+jMKt4MiBVidT3xPwfqlIcL2RQ8d2/SPklWaYWVAKy7b+hMJ4Nzvi1T7PoZtm2
dCrqYxHmOC7udb5cIfG7s7tS7hHDKIeKB6QUi7Y2OB0=
`protect END_PROTECTED
