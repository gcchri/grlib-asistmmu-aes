`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MQ5T5v2/1J0GlrcUN8j3Bnj7QhT3Brxe6jizaCm3XBCy/70G56aPelq24H3lGD5J
di/uUnWLL8XdbVlK8NLxrfNelapM8MrvMkTzz1rIwBc9fSdhopB/o7xrJbHz1s2p
CkOucyokWXjXelDO0R3Yb8RadHD1k0fh6tKl2jT6kqCDDQ8Y7SKgCmJLyId7n9k/
whwcXVlZV5L+r3CjpEIsO7AP/ITYf2n7bzjtuYEey8ALIPsMeHWm0MPJm75A91xJ
hZeoZmu10tB1a+mMbcF6UK1BK9qqQg6BEOnlWwtzLVCvVR+X7+DuVcKS297nyg04
mA+9OUrqpHvz28SqPiQMBGGV0WhdlaBkiDxwVY9JM9LMrm0aZADXXFhqWMP45/WZ
VA8c1OOFbe2NjBpg2/vDEV5QPbMFQ8mwxjW5Zw0AQZCBYPGcVx0kyRrihUjQwVWA
ez9T6GAUkB16C02SoivM1OfDCN4jYAdHtrZk0AygEQieJpyelx88ZaM7lKCXGedu
NFgekQXOV0aPYzgMdsTKTx4R3Df+Ns9r7lZ1SYK9qFACy2m4JbJNsO76feOnL8kP
s7hdcAPCYn/xDQ0CXck3sRGiWHvKtfzlzIp5Hmh0P48OB+z3IJq1iDBJWlACZN+j
vMbyV/Gix9stFVsOUA2RgDpTJlDGVIDoF81xAaabK7Hqgl0PjXdez8TENs4JyJot
S1H/sILwEMyWq9rEwBtbLP1ecTwQ7q9BhF/VK/O2kdMCWYcL763qCnzWNOekzNDb
lT+VnGWlOUa05HqugTD/o6x+/sijsN43BV43oPtd76DGPBazhEQZGrSX64ckvUIQ
bvpilUIzH7JjWSxEJzXbFILKQqm9GylZeyl+16vUwLE+PdbDQBqnUKCbREHccFkz
r/DXfq6SApRVbBfunspQodEb3CQkf7PY9gwjZxl6+KCqOBIux/qME8bdOwEP9mcl
GtWr0nSJnaGNKG2vYjFEs89Z5cwCKIkQsc1MuL/fwZcHBdpOKT2i9TUZgkR8iim1
Ju582boXHjEGDUuMLM2+d9wdU+0mj6bSrZwumlsdBQ5Sn4feUF7hGtRgehu57vve
vYABLm/reXud96xXoY5OUoJR7Wap+yTiug7pArqc4VDUk9CvALxLV+NJOY+u86VP
3U5xi0aKHS5JVvjZscrnp/rdwiiuMMBihR1AyUV/37ZNJ3ygu8YGPz6SNQ2CFSdG
`protect END_PROTECTED
