`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RP/1Dkj0sXOpRLvkFWop+EQNHLwaOriViqIbk0OT3FYZYBxpDt+qkkDycRqTkH2F
g6nGCftW+I3OzFKh2LiEInHn82JPkzUeMtY3PI8DXRmUaGWAG8M35xx/rBx7mW7C
tEH9xLJeLBOt6ie+9R99+CHh7CL8HY+ny0guLpYoHbWYUr0zlVtPYDnsvx4MH1Tn
Set6dV2xfSR/YzaRt/PzGkw3Du8hktSfSOOqkAHtuoqS1h76Fc1Bu0isdXFsyVTY
oyjdqiNczd7i8IRU3gwH+PR6bE5PcyaZ9TvPngApZpp4hhEtn7nCmZpeofSekIx4
u4Ylbms7HDmMr4dRelHRgQ==
`protect END_PROTECTED
