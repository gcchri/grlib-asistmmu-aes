`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ES3GgbjRyTT3CWY/GtWTwh/Lg24f58yOt7RLYfN+JkhvLMG4Tfd6iEWRMMbVb+P4
Qzu+4xgZ9SLdwO8wJP6/0tFwqYGDziLzqlXzYymu7b5OED8U/OdBAtfUTehZBQNh
ueuvFsIzzYgsbBAroqvKVUUBFnh6eP/h7PBVCXB4FcAftzXFyv/nXI3LolKTINzV
zP6w4FBD+apyrmjLtCLJrGrGvX3lA787iLdDEAgrIGj3l4HaoKyvR/B6V/9A/2W8
Xj8xGZvGPuPxFLc1xCiLMekGRvR5Cwmzup7pEK9Zn84=
`protect END_PROTECTED
