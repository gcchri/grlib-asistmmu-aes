`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lUo+oRnKoGR5CFkq++cdgzbWzC31ndBMllJZeUe//x3ykgaxBS14lJOTMz2nNIDO
UyMYb0HQKG4QoHC0AGfnFdXcG0uJBZXc5OW2EB+NcAYrPyj8oC9N0u1ccV2wn4Ee
kEdwmkpUr+6GiaeJst/bDjOhpifl0gfhaAwMz2mwIvFyKDlXBjN8I/u0DfHYIFlS
y0PfSeXnH1EY6mdhDOLHM4bNXHtxiULif4XvuUCIRc+BMTHIUknlvhUWlF5AdfCy
f611SZ/Ih6tiXIRF2k9olxOA6ztt+Tyrw3Li8kQV2vOzEyanojZFfIUQ1XpRPyKY
3Z77RTcSFncoZ0bm/ZzBPHwLEJWRXqn2wJh2NgGjOIdHsgzQWCWm7FpL44SdNlgz
3FOg11LEdy/t3pScbRtPS/2vuRP0e8MSDqam7tNtSqQleejVl0ME/CcBGlFposCT
nq3mx5opCUyg2dwQmEMjuSQapZlRSIW6sYJKxGrjzl7cQTsUiPKV2E1nUsDrH2X5
Wt/zR9xRlzA+u7ulhDop0w==
`protect END_PROTECTED
