`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sIUHdSOE1tuOV7DvOhr/VT+0DBuzU2V8ZUwp4zzIzLouO1yPg9PrlUBx56Ddwhly
ocHEBqExmZUCZj3wv5QNq0YjK2H0LERVbCPwwMvxYYY/3GVCRDEaPOYt2VigEZKs
OL74r7JKgwZGnJ2pn795XvIg9kx3WixEcWkWEMlKYw670oJDV9fo/6vm5kWjbUcw
i4JwT3ea7lRXMwLuKH1IDV8MKfNp0C3cJX0LLoZJ+5k/VnkU3GuKddt5TgU73gr7
kmRz5XYuCX8Mczsj0KiGrA==
`protect END_PROTECTED
