`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gu6lbCL/hzNGK0WzgMIygg5ki4YUwcEMF59amvLG4iBI3gfxhigTHvaaeifvQavm
BkPchMwmwSxd6BqJSqJQf4Eg74rTPXalwpR8AYFqlnpTbhADQBsvg8ZuJoxpIncD
puKtRb4TtpGLqmT3y6mN8lwf0mIqcj1G8ixTB859fDQYmYTvfOrM3cwq7V1Tt5Ta
PjyHSXTBRBQNfOvu44eofE+bCgHEnktnVwISMjGgEXM/eju4azPvdP2qp9o9GTcU
GDy0J2/amuNVVMf3um53P6J0508X1X7xJwOtyK4Eqe5bWHKK8pvvRDaIwJ0QoRI4
AdCeqyE1vjWGHMwWUEutEa0ly//3ArbEDpqdl5OJcBDU0ba8t2YNk+2yzg1GgtLj
Iur54zr7QEHGvdpHZ/skNPnM6pfacPMIwFwYr/XFc7vuBUWbFNkUw7h/AleY6vx0
T2b2LUyMi5WcvwkOpLJH0lGrIeABGLXhbWbYdeYkcN/PNjh19L4YLaX9yjDSQBPy
dcZyrb91GjqQkS5+ztxNmAAKcUe2re3X18rSF40wS4qEA8OANCfngJLNECKvca4W
2fLpITkz463FXzY7ND8KzA==
`protect END_PROTECTED
