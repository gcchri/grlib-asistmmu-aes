`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yr68NStjZc4VqyxTWL1rC7IbujJF1MiVzRVXH+LlXzakfWTlhMD96Tkb0GO8aIlz
rtBuMk8OIHL32hBm3UcRwxkNwNH1PKFhfa9no+1G6uIlPnBVewbCZIDRGvcKj/ss
jQjMNkn80MeOFTTiP4/GmVuMGksvZN5N89bs+LHf5AGngNl8kIkZ4XGo1Kl5V/cC
FHnjTiHdsBIQn3/V0qYdt4KN2+W268QL5RxR5l3mw0JHWW16LadezU/HXhX8n3rd
iWQ3LefkRmuZ9lh0IDnJ5Q==
`protect END_PROTECTED
