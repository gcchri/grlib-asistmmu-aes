`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tb0KOjJkNshsgljE+DvETuEM3Ys8u5YlToI6g3wHNYvfO/DtaF7gukjB/Bp78ZSV
khA2ViTcu3shdfHH2LsiVKtZEI4NsunD9aBqHb1BWtxTVZcxg4YXa+y+SSTOxtE2
8YhZuJ+yATuBAnlNfM8jw9/DZ7d1NAtTwxdcsElFtLY8v9/VhZQQuiwySIDQJ20h
u4hO5VgRyrFILt1wU/4mYXI1CvfcpZEhAHSKYiYr/oy/C3jpq6+qF2oVjhteDwAM
gWcO5omf4ykR5OWSz4Fvq6dGXwfIFTZNcduWmVg5bPS4ZcoEBdIneuOJFzsbF27u
NDlDibf2mTQtGxAot4MhNxmMMRhj8K7vP6+DLYjK1c9tDSAHVg/aBlOG6/ulhv6Q
/8NB8W9jKJR8FuQ7MC7Yw4GGCOyck1rNK9OY5eXItvD2uKJXvb4U7brIdW5XL9p7
7Kdz9oxShEpKDnQK7aeBsCL5c/HdlF71Gm80t3Rq97tXVT8yEgKekjsHpCHrA1uc
+YExaoX2jH+Ev76Wcoy6G8TfhPDnwfxFrxFo43XbZBabHveUDiVG9LTpEhJHiicd
mzpeBKoKB1d0hHoc6OAS4oZjOMHlGMStwVh36XqLbmCtEBxYMxuX93liqVHL2jpr
R7Vk2zD/mFMrW/uELyaxzJh6fEAagStycb3vWd4cbkxitcO3O6WnSn6bbux7RLUx
/F58N9YfSBi36kHSfKy5gHYDtFV2aYv1AHJJ0frmFJsiqmjSirY/dGYEnwITbHOJ
vnJ49EFa/RXp0ai2LPb5HDHdCE9ZJWdFhAfjz0gS17NTX9BUXFFW6jrOc9KWTmRI
OwOdhc7neNTP17Zgx1tGq2WZUgf6BWqpT0C7M13CgjE7sQal8BJnU226qLFnXTFj
4FKbXsNNPPRvdudkKR+LhW1w5waqR7BAM6iKi0pbp87/vmLeHiwneuzOEXk3k4SS
6aruafsZ4/momDVAsmWWYkhOSa5kl+pgYCGm8oRmA9A1m6PFJBw/Rk9dZQwTGIOl
1g8gA0nt9mwSVKx4cjsbewyTOAsSgi40IBbiutEOGF5BkBjBNPzeyPqLPIKwitbE
gGWiGy734FjFYbrttVO8gzCTVM55EEWllzCW4tXdiMbPks7AZCEd7agP4Lg9Fjkh
cT1UwkLi/Py5PG8A8c0xycoqg14wjajboflqsdgH4yvKjEfKHlObc6gPwKqIgI4k
klwhq4eMW4kSEU4NFW0SicNLXFZUfdaoEDLSDQMm+XPuKNL7xtHfu0M5FFFhLfZx
FMNBCAq/5ZksX76cPXTVXQfAoiN1PGKHDMfg5R5Ah00KMAh1I/AkcfD4ZuKJDi7E
vYw07Wj8lBs9VvOREmIYPP2ZM/+FTj0mdIUr5p7SWTydFNHC0DKz3LWgAX3cCqwO
Zusnmm7+A8LqiHnIp3LlZA==
`protect END_PROTECTED
