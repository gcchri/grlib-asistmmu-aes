`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r3WVZyrQ2fIelTL3zNyPNen1DldagUoCua/B8uDlxS5HecKbsSyiX54tnF0OW8CK
4sP/xj0WyzOfai08NLfzQxSWkF3JxsiwrNcGePpAQHWnBwwZM5ZvKcvRbcaBKNc0
F3V8xwqtWOALx5Rm89QHfqRvyJ+knb69siYsWUSGUIFYS5uqJPsqMT6TUsEgtmWg
Sjs7egbGmFvK82/0wEEysoZqqTxK0VMBYXKr215hptQpL60LWKdZnQ48XRGcvtKh
3BVZBN8JF+qD/qFcvWf/DUEX2u9VP4/5FFbu9zqLiPlfRTmSvxnzLXP66vZcYfBE
rz6T445V4Pqd955Uy06P1KJn7NVanE7M/HRNHftRvejiwg5UjjRK3jLAM6lxC/2U
kNLUUfhH7i4v+wpIVBtyMl8pwnsJJzq7J7/ypiT5xARmiubeWXG5MfzJoiZXe5UX
MU5sgtUqOL/hofb3hVUKVRRYJOF9A33IcDsZsrc05fznNcaKQjN0gMgsar9wH4so
e/wys/m8KsdckMYS+6GWe1YeYqOPuoRqxszXmGNhuERJ9dtzW7C31JamN4ODCdKc
Rug9Uh6t8svf7NjlpNai1EWlWj3qS2FPxRmc4p8QK3hdjl96mczbYcujCwlBA1Bj
JqHDtMf3YSNAdOURCYaJcpo+7Xwt0sFp4RfxUakHVftnSrwC67caP/BYmNFZQPJc
i/9BBLGVTW9h57L9Jj6eR9ClmInWNy1/33KDbj7HxUpR4ljxaxA1U+t1OxjLgJuV
ySdif6CoXKXm3/bjQ9MWgcSlyVuUuUjtqK0HhOKf5eoUdSPu1HgAXWMZrGnU7wWV
uxr03luvgZAGffjXxqmdJg==
`protect END_PROTECTED
