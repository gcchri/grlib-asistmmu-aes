`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w+cfoTp12hj9K1P/JcdWcu/0t/SB9jud8pRpOQ/DGVnL8lwIF8Ei8VzLAGzEzB7z
vule/+meIP0DU9FxfQ2zQYrdfwHDxuSy62aHjNtIxPGHwNAOTBQg5g8Sah2EPeaf
ILHyAKRs8gGuJKum/N+maM70CcHLg/t+MCIwwup8l0IUM97IAre7Hd2S2jZ5ojwH
SzWyXUgcdcqjE1kMqK5rhEDiScHJURSdHzD35lF/RtgJOWMR1MhwgGdTg4UCTjGR
9SAvYAbJeaEY326oX5YtMvBdTUcO+enZ/EtEKLfr1uLowZt0FXCXJE5NaoIunj44
n8c2WYtacvjkZ4kCRU7Fs+fYjDSVJcCH98VP16gCmqLjjc2/stROSij2tzyxayjN
`protect END_PROTECTED
