`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dR/QTI9yPo70SyTEswaZ1fVmbEqBHffXo4ehNbBdNAzKPUbyy0/kRzBHe6cu1VrZ
gsEu8q3LhVQ1ZHn6dDyF59cM6CGo5oeoWDfnvDzNnJsLAnFeaBH6zd+G/0nfsaZy
J62YpDu0TkgJvlm8aHT/oXFTxDQMqxz12bLsd9DHgDlwRoGenRDog5MCqi9ywtkI
nsJyKr2imvR/gupNw8+pL9zEFNxk5o3iJoQco46O4ZKkdRyVmXV+Scv14TXhdOsP
qze6aXgR5D5/5V8u7zj99HhmhdnkuGtezkbPBnKr6UDvotNvlAeZthQNo84Idx8Q
5mLXkXvE7W1xGatw0+gzGwr8Mh+0wskwfR5ribo663CRoOsjAaWz+8O90zZXWMI/
WhqRGBg0ObN3Nh9SvJCzFuh/eAmFrKi0Ur3YQDqPfxoJ5BC1+JYVKU8iLy4KKJXt
eQXFNGa9DBocWwMEE8qeHI7u4WFI5vzqOfqZK0J4gSAaWCz2moTnzeJ8hy59s1vF
sfHxOp6bAYu/S0TJBX/AOviQXCTqk4igeFTzJmJa+X2TMQqmmQXqoKCxySDrm2OK
f+8FQOFhf8gPdy0PWT4y005RIjvAfwskLsN80HBJxfYXXpN42mtCI3BOeJI25aet
R0lx90R/s+dfynTZJ66pfDGWc8ERn3gSYW6Xa2GhDmNBOnp2F4tJyp+SbukuEl4K
9Lt4qfZTsQP7+kNQjrIQCryExRdH332MDeeX/YbrkoKxIdVOzn+0OUsvAPR6tKFu
QaPNCJF5Ygm+u+dLsRcu91GPGtYvAujnLZqJQ8gNj3mi/LmeGaXYBFhbEYOq/EYr
T6CxlOAjBzvoLg43SJ9hw09nzxDtNalfm4TCR+6XalB97/ao+1+vGORTds/P/EH4
oz4gYrVcnrgcQdNOcb5/CX2qc65Qb004h7BJI4ojY0ediCDLyMNu39eibUb41m7S
ufAzsM4YE+m9YEw8eUetjd81BKpxYvICapD6dJVfHqgJ2KGaQrOOpyKL5EXad6WX
WZECKGEzYsDy8B4DEbqTxbZyscAJy/sBSiAV9zMYBylf1uimdhTvgm+HW+6TtvNZ
iUvJRwJfgKg0s/H9vnmcrR3As8j+nY+tvxORPK1Ttd6dTiOFbw4ZaiLbVBX/wHks
wUITzvnz5VATF4QOgHnOKmXijedS+cISB28wOK9nqRjKrmQTqoEtaVFMQdIECge6
VQdYwAkTokDaNCdcBmn/8/dikQhNCt66Chkd60rxqEBBAxCLdIgwBVzMnWm5VVEP
POyHAl8vCmAPFW69eRYHUT6UYthGiQjv/E+qOuHWm5jUvqvW3VBLEwkLRs6beo6P
yXx9OylFJeHpV0/7y6yHN+AT+qEbxRXIpPq3Gz7afNRBro5nAjuN88KMOBOgXe58
ZgzAzfQtnMDLRibmtIxDJBsu6k9ByJt/ByF+02FdPpXuVLKE8RuYhDYzhuQfH56Q
04xvkeNxzTfFGWNRapO6uesACzgNmgMDVyRraaOCMuGYkTpjfbeS0hvRe8ENnoaI
pg27cwro+7xJmVDls7QPrZ/ghc16E8Ra+caL+vsOPjyKn6AmbAbjDOshGcmy5DAI
B6pGHG1D3rIaOYGY7u2G7KMrrMgs+4nL89gPjZvaV+qC3bR+qwTCiQl8jYWMXi+O
gwSVup+eqvRxtLSvnlZDjCWcEJaMAEtqtEjitL1NYzCZfdn+icNxAFc/YNeDenAr
wsABQ/CJI51m4KPo5iXUydp8T9N4NUCUsfOFqQwLUHdJsTn0RCK7Vo93LABctcOT
xSTp7WWXGFwEJdbeCRLxbmWoBFMn/rlftDGiNpMTTq27BBFKftQvKHELT9JRa7Zt
BqxnxJgj2+pCcd9WAG3YZuZe3Ud/3Y64qNwzM22vGCYH4+0Uqe732NbyXpUXFylP
hV+08T+TTeU0cdHcPjoR8APNWOu3O4MX12LcyAfNAehlYyWzw41e1uxMdrJ8FjHX
5FJZpwUrhqnRwJ2CB/F9JKzYitsV2m78Tlc1DsmfN+t45AaOQf7kV9kCOEogxsSg
C7zTY9sCLjbHru26NpWoURv7P5UvjELkTOSUGvdzG+E5MYWYSl53BFcfSEFk/+H8
PGNA5ATU+49DBwMoNW7oJxNulGEk9xyEwEFb6R9OqQqy7+oP+WoMfe/P4q+bnDVF
epS3e7GhuzWRCO7I1XLFDuP1XW4V2ylEY8Uk41JlBEB5fIKL2uVHjB4VbqEVWeZ9
EQyQ+KJs0MMacErXgMUmibJWY6y+6j7649i/YQy1eYZYBKhfiN+pExRJlNd1DXjR
H93YIAifS8yMf/6hIt5hE2v+MiFBeez9lAnQkmTSZonkG9Kqqh5Bs42TQrFz9z07
lgwQPfqKymNn79mp+zskk4ePLlnqppi/v4Zga/J6ShCL05ZtOZ4x15HZVsusZlSu
vVyLJ96gqyK2PFhHzPsRt4u9gUOZpSi0xhy67jSq4NPwzQzmSTz8VH0UG8a3/7OQ
g4nC+EigOKnwnaHGMKkrCWUqCldAYoZLVRqkccnFZKfciaNBlTVzXDXyg1rUKBHN
uBxXcZiVfE2/wGt7iMtxeOByKT1SBWyh6qh6ixWGBT0AWuGlMi2NUxHUBv2dYlq3
LkvIqHRMg+9DuGMANTRhPg8RcD1se+NQhyXzhjZM8L6i66EDX4ORWEsubSveQHe3
yUldG6anh4lsPZl7oUjb5YSgcCjd6ROLQ9bFSDYJWieV7EL62q4ANg1p1kYsowBY
bCSbzqu5P4CetcEOYs8Myb/OZ4YFo8oMCydmSa1xhZcIhBCcrhfsKpWRp6E6ff/a
VRd/WfTHWpPIwTocCt4NlQvz22+JJYnN1BtwSWyYT+DU+F4HV6VKuf72pkFvAPve
xTvkIrtfnMN0QTwIlvg+Wr0TRMSVqCeIHgdEhPqDdS+oUefYYnD5Ko2xlo1TrKqF
1Q7t165W36ok3xNJKyDWeNew/M2+euS3kqAP74373ovkbgLELVFrfO4s8OTlECqT
qX6m+Wp+SyiKvDvzUzhL4FJb31xCVV4TZVdgCLApyYlEwMq175jNDG2PYs/FJSNw
7/sakh9M0i024Fx3WumbYz8Txs40ZlrTHFT+tYKVA9WGpw0xkAKHzCOPaAu9XAka
FDlkkPFgnTu3dPBPJhxfyUxW/tCXXwksRIHhoEJUxmCcj5IQHWnitvjYlnS9G7GE
GSG0i1yt1g97bwSjaDCYjQN4PMqCOP/gCp1R97hbi4mH/qiBQGO7DT+K0cg37iVX
k7jMi2WPF+jdjj0TnEudDJDo8HivIH63DqsIEP+2H05aFb0sKqxnux7b97mC1UTG
1SPczMHXz8FFmhasw6yPteisLA7RqLivpf6JT6RFLkE/sEzRw3G+AY9NL5sBfvS0
XkSU5lgE6z+48znliQ218t/OvvJyfh9b9IadVLLU5tvTevIfam6JkmyUKQEWOgVA
h8xAZo8ZB4KVp221+nuMgrrsvYF4sS0HEsTpDWKJbrm5EEEi6s4LYQwH1Lgu97kU
Zuh+ypt41mqYo1fPjEVIVI+74dEbftmXrGx2UoWqpcgJVMqAqdEEone4VpNoPkX1
iUuJKlzH8lLTLxa5W4yaySbwGcrTwQsBhutsr3+S/4+oh3SLGjmFkeGZbQUCtLt+
aMarzqjJMBzi1REkuwBIu/kHbJxF2Rnpl912lJ+em6bsT5ZeOv1ETMlfU3SsYa5w
ATutioM9ty1GxP6FszGH6kTsUv7ohda3folkhVWrrC2BuV4ed1F/mUqVhbBPgEYt
dRam6T1RVcDv0irIeV/ljHRVsvaMzb0gy0a0/ZmV+Bu8lZWVVJeS1w6Y1x8fJtE9
OEuOacXB5ebzCg0+DxNcSYiwxg8c/b5s6vUVoiJF5OwjeogRmYk+h9+7vG6o0z8f
jkJsoTmqGg/1s8m3PD0X5S2gXPzbrQbZ4FWsCy6czGB0nECcljemlpf0Cxx6ux14
27Pj1K8sH7fHn9GkPZXZoS0PScXhwAGZVowRy7AU9tZ0Xzip416RCZ1KBkYB8Ytl
Z3O5UT7ogbeMsUmXikWI0L9WcOv9n8aWbc1h8W70+ze+cPM3gxIRag6Z/z2mJtPj
PXCM9lsNmWWoHaqd1LaTz0eaWSQ6qEFdk9RpL0R4hxQy1RzmydOa/5C8OxYB8JFU
3qkGl9XBWLiuuISZ/utrVf1Xg0l58+UganoLVn+4ZJzUTtdrgsS+XsF77JjdRmdd
cOCaDOhz5MqJ23Fbt1p9OhF1EvBdCJZMgWclWNtCsb2tApfxEac2RAqns72NAxVE
iP/tj1OZKgbSlmtKEPjiUCvWjXqcU0DvOdNfm5aIrWNX5vy4yLg8C/2J9/T2Agg9
b8/HYi8B8GqmR33rB1r4JpH3iRcAVQHadPsaVTgZQ3jCieKUIEwY4o1m6mVztNgX
Ga0evT3U70U7aMiixrV2teU0NuerZX7/wkaSvJRhm2d68fu0KdQKt/gzEe6iht7+
gkESy8WVBTZcGYQ0h8TfXjoy4KIJMNJsbyJa7R4ayJ3NJg2517FoyxwtVH5XFSxd
ATSVLvslPS0KygHF67AnRfFdVV265HsQfA+g4xNtMno81m2qXmvWjlp2rhNWV3Vn
ZqJM8w0Efj7BqwEeNLz7U/lCPOgjxQaA0rlP1j2xZjfQXHTmA1rcDeP04ajlxyNY
kOGaxHBNBK3L9vQ/7JCHmPOjlTqgu35XIs7Yk36STBZy25FYiIuEBRr29od6pPtv
oPqXpjC/Pt76U1yCTTbli/9YKSbJBY74fnj2GZBGyM6ZbHR9C7pUrTT5DOLPppC1
Ab6qKTm30TLLbuBJUxp5SzJJeTKxma93Q543zZkNs+sk1rNcIsbfr/OVV4sbL/XI
qxRrj1GCPcVwdADmXmPaYZ8eAKydJMbf5bdTZJE3Pb7vsR2rKD4KAtnpdrO6IGcv
mZ9QU2zHuLF42dybNaRw2HnmO+8OLq33Y4iGSjtZPxad5iMER/obnnB+KGndxcJ1
Ohb6uja48R5yW124rVQp+kze4XRf2gc3yiEgbvmeM3hHDivp62a3lnyyrhYvzdvh
0bsZqkT3BJwfhYc+YlWRo06cTc40fkMauRfU/AMn48KeebD1xMlrWLEWIFMckMM9
PnGlf1FuiRBwFjNZ+n0wLO9PA0hqTAXuWTiuUxmg9n7vSvzZNawKfVA+dUGrhtvW
u1XZmQtgEJSvYJwBu2OxxrP0DKMq5xgeY9xhlUi5e0ID4EFmghjKHVcQeDk0R74O
kxyja/RWficJzs4+ysYJn1L//N9ABDVu7UrULNIBPZdr9ojpuxSBkcXz+Rx+HqzV
g+FNGiRHcPah5J5Pc/gtD8bN6EDcn0Ecb21nbF+IwEpLle8E2vO+3bC2jtb6cy84
z9JUunbpqUvjo3mWkwIgzOjH1chd4MLL+iM15dqDvW2rB2q/w3nwcbz0i6e4g9Dn
LWyOvoQQhm3kxPHIKB6fWbsl2vvPBaqflyNGri8L+7m06DcqeqM9/eF5qxIKBz2w
2j83+SDK2JScaKWKmXIuVEKvrTfJYLF3ApNqi+ppEPhGtJYyzfaVY/7HSMgqzEOD
QfOwS51+UjRhKmK/9pfJJ+DKYqzm5t9sodf+3+cUT4KxejslYOsE1rSYvmyEKV3z
C29QhWscvHwqBwSPoOg9NjPV7ERC/jHBVgRvCTu4ZEF9pmYGq6JgJb7w/2zClEBG
6achOu8LK5F6JRfao8OGtoyMsH64P0r+uiY8/8x4khUGuwDvQ6MrjMYoY/UIqnAX
INaF6vBDkAEzYGeDtxDUN7m2Zeyty8n8Cb1X4/MG4qnhka7fe3xFcO60dFnSy0qP
4OwsiIDHvY/dvZj5Z/WHdwPw6/CkQRgR5z8o4Bh7G0nYgN7pv+N/KgdUk+iBq+Ek
HLhJGjKUp+TQkSlao28WvmFWVIuGMRDXLnaJ8JjOc9N7wZotlUngD1xgImRkUAkj
zQ5mi8Ing9Yuj+sLZT1yHsJbZmfbkeXS269GfrVzFdXN5a4209xduQ4/MaZKpxNy
wEl2OogLKj+HlCVryQpJwzmzPx3iHRkbQxGBgobWBzk2uvX4AVysH9UnDdg2Arta
TgXD35fj4bMyar1J9qQgzAelMI9Zd2avx/ABkB0qZMjLmusm3lPLlCgLdIMQxkcS
8FITzgBXcoyXenst8SZoVaJN7uo5Mh4uctbdW/pNqTRXe5+CHhcQ/TzXhEP8na4u
1I/OQyQ0nlt6/Eo+x5URuak4PONx+h5wg5OEmqnx7xHx52swwPxeZZfn47lXbTV5
cFU+Oqcfk5D25ZDM1FxpoWX8SgfAj4fZQcAb7fDORxYW4f2lk2ZT+hnRGMC2dppB
Kf55Nydaxl7kxOX2NGrJ8n3ajJSngAU9NntJLKHcHB94Z0r/DdnBNZSXk3n4D/Ya
u5Z3rhnrfGqcnE8PZIotug1Uw64Rb6eV1vjPqVUj344lginzIyw5djK8FXWr00xN
1ACYOFPpxp5iTE8/jsLGrSTeoDY9IiPw2i4x9+HUx91ZnzMs+tpr2prUoLZcxpgE
vl9BMNX7mzaiOGYd89qOUi2VFeiorThc28WMOJdcqjK2M0Oz/Lrq40LSqsEjVh7J
97t3Yw/x39H7pdcgV3+Qs6Wum1MJZa8UNALdHBrPoCorv4cZoYFyPEV4oqWNPvqb
pq+pAfgq+4yt8/F/14YAvBtfpvTK4pcu/poitSbRjt9aRzSzSiDHCeY83KizUOas
gUOqOssUPLzFn634+zKTeodVf/9FM7d5Xdmhw0xupr11cXgdK9ZikdkaPYe4e74H
MEhN9lsu/XK5B6p7uuBnWc0f3+E32skjJmG3EcgtomAS4gAYKoi5ksG5aEzqq5KS
RAeLDFpC6OZhrYUwCjHNAQGgEyHH3IlAti+776UrX61RbasS//fXHaVk5YYX4gwG
1sWaDVi5LSN29gZqRzOyQEPeSdaebkUa2D97oRGLUpM06e6TRHGKIrMGhoEQc+sK
cNHXTZJ8yICpiBhUP857TLe9X6+55d0flTSkxA+JbeXO0xkugPayL4RNOv9qsiCm
YRP2lXBWJiu4hB/rBLABX2y/KLNEUbcKJiVhPmegDINjDJgqXOQPnQvsOMYYQSke
V1bMX4Wd63Sq+SXxQYzJvycTl+KeB0U23WcYYPWML83Kc7XsUeRiZFyE+la7yUJG
sUC9/3D/xxodHXQHYyf95nt5OOHV9Dx8vqmBA6XdEuzoDCY1abY8HZUG/bfKx/Tk
5CE/VQzGUIQn0O10Ehu3D+Rqto5PFQwTSvK7IXLZV/DQth/+u1fWrhOV6nH6Xnxy
4XXpJBaay7wHVbgF+J8iLgVzv1CrEbp7hhW1d3zxJGkYbUkYv+FNXBOvYSz2JYBf
S5P4Qy7OkiHd6IxsAztv3kvZq4VEDVIPxL/KHjgSAH+BL5SMEEBBjWFgBwQ/9Ovv
nCo7jCVLISZOLLINntMyrGJyG2AP6sq9ZzEXl3ENI2DlEbGfPaxjADshg6zNTWcz
4v6F2h9PPVOGtiH1zPCo7wGTW80BeIWCx/yoFGMBS6SG6gbnAJ43hcs/zXJFs2Ir
0zc/VLyzUC2IpTL4kxCGnd+cI/ox4rMFAdtGQcKpbn/6DMlWvkkcI7If44ojo4oE
VVBP9f2dK8ENzQ9H+ZCAdhFrV2rAn1EIVrhstunXta0ppfYu9JK9h2u4v5eiQmlc
fHo67YwdPbhNfLTMjBJmwGjP7xaEhEPq+zRN1MCX447KdBb9YNXJ6Zx2uobazr42
5Sn/5UvEfLccYJFZOAPTAX7XvZbmN7nRR5NYb3l6so/xINhSaxsZcAg6U44Co/G9
aKWg0y+9djAHrv/LWgWsxCSXAfMNp+OlrxDcs9YXCUbJz8KClG/81ryFfQmoBIKQ
4ClTFIG9dm/jPlffJVseGH/oTNOok6va/GoNTrVPQTOAsSDNThHbqYMeGmyWlCHP
lheIy6zo+Omuc9Oy880kPg==
`protect END_PROTECTED
