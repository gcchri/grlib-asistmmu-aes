`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tEBaj6UaeEpkTk6MjvyDxyqGmG1ZGlCl6MN4r6TjXplZyFskeJ+zGGnV4mLrMPFE
pNPkkISMOUAdN92GA8PY3t5SVnPYvLmU3AOBeUwOs+mxefhBu+MmFmeVjcg+M+lH
j2NfcAS754ba7eeLZjBbG318NGxi2T3ziZ/jCxlucYlJtntqoO9QrfyUSL3urWDy
SgFmB5ZVNuyn1J/IdV+KE3O7UIus42isLl4OKjwpQVHFM931OFYQ0cqvquz7Q8r4
K7g3ytOoh/D1RQ2gXR1YoRkzGf5SARsq40d0sDBASCmA9fmN05GlBeBW0+57XfLq
`protect END_PROTECTED
