`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hv7N+eH0CdjtI3kt/QORpp7ecnKxfhhUjyVAY8Iln3rHbATPeclU/3PoVezOJgqy
x5iVqchmmOiTBiFzZOtae2vXlKCfCkBsNhgi0try089kxdjrVErRZfynVU0P2bQm
5NenPPoRedAsXZzsUR9eKlwRs+IP9ElXQ9DEVhfZ9d+nVc12hzdWBEaUWvv3zEv7
boFcyEgkjaCW+Ch8wDoaG9RZoY4l6vJt5QOqM2ZjsJQi7klQ1+ze1kMCPmX9lJol
iXDvxgorOLUoAMja1ewHZA==
`protect END_PROTECTED
