`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4EJkInv0ZrLhafbqCsfBgS70omuour0b8sr9EpK1+hV8G0XykOCDiI/TL3B5u4Ux
ddloVATNm2TGrH/hDK99iPyqVbD4douDUNfdUtBB3Jhh9moUa6gjwCvRRaeqGCoa
pcIFhBgDY0ZL2y74sN9lOh8yeHA7Zuks0sguGH8QEzngGYW9SFRZLh5Gn7KWwN6X
5Bokv8Mr/Z9ea+eaLsKCCgr3kua21Bs2sIlxT4n1Hd0ZxcUjMW1ADmf/qAd7xa6N
9FCjjrExdgGhQlzvFHD8ms7X44pI4e1XyZK4+aPxIwP9rTurn3cgyJ1eaLbrkUwG
rK0n3A7Dxehak5hlKv7Z8Dq+E6SeaO6s8YOfaiWvHEJxLvHjdpVtuB0LsDKbLlBw
Hqx/w1J5H85CyttOJDTG3tXTqNTgX+AuyPbqEgMJWvw=
`protect END_PROTECTED
