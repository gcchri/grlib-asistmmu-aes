`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A1ZORWpcm+wFU8Gv5eVIkWTwtJrVnqqgMKY2b2Wi6EMUFPuV1Z/+zjSbJd9wcIZP
nGC8GJdebzw3NLAe1MOHNtpUi4V9iS5YiWcrwXhA9EHgEMbjrwqzVcLpHExD9H3I
NItAyiiiI5dPwDkAjgQLkYuAFBXt5Wn576V7u5TGQoRE16lUli/ZOfUKaVVYA/Le
aIJMdR0PAZjpWxxjltgHF+f0isuAYcnTwCsHNMs1HtiU5RGhpFVVG0FsifLHsMTu
vjWsKZJe8FJ+0m+lAT7G54nesQx/Jo8ObVbCvPVKSCy+LdzsH3a3H5HMOpWoSwct
yHi0spjcFZyUdQgW08zis3A+I/8gFWm3UaEPzMmONokcwrYujfO34W3IoY3Yv2Kc
2HV9wsBU7aA+TDCfsJcHn2myd1jXe1HJZygyO4wIizPvrNhlYkk2oIZLrWTu53b5
bueu3Y9nyLDZA6LrCddBNydBi0ZOKVyQlmoJkMYJv63S+M65hp5zcv+Af7YM6vq+
CUpg7aVAaPP+63cLKe3Qqq6X2WJW0zgdafQMaS2jb0bG+sF53fKaDBmBfL6glct8
lIBRRIpTSwmU7Uko5VHfUe3zas1Zg1xNKU5ahZm5RrsXs4eOPzmBenWl3pLiETbC
vb64qvBmnkfXZaosHen9A1nA2YxoF6QbcRWAYv5YhEy5ZHsBcRiYQyQKab0ET7gB
VVwsSrqAK7ILYKkCzATUPqo+RjiWOdMFr4sbU3N2YjQ3U+pgXpI9TyjplB2+/xXS
pdhkgH2CsmF3eP3Fap1jnJhQ3/WsjqbMMXRLC5zlHzwQ7rHvJ9QRsggOakm6Rix/
vBDh0gTNp8PJSL4s4IvxyMQwErinpRlV65sylFTcBKtjVG1fAIIAS6swrOT1zXNd
95ol3jo3eGw4IIQZGRFP5u8/YOS4WnkmIKgI23eqZXvtioxasN/V+wOW2Kq5950c
L94IZfwhZ4t2RqGrk+lpKbXw23MD6JwiWvhI5xyQ9eM4h1MLHXZ04msD69XalC0X
lfHzK76giMYlAYyw5vIuK638wC+aPRoa7BOBPKb1WBjkRo9Uj5XG2Vu1XmNi5H8v
Wc9+RHZqoK780pJpDQm/7GY1uCHpPK9n5VIhsdK7dkCb5JuE7OoLCHDxy4q07P/d
UH94q3AI+WsZIVQ0/IR2QCf/W8dflU/1UzphIR9/RQtCxefupfizBDSO+e5M6XCH
Rh9m8reGVEXEsBTC1kKfTQUvA4sudNMwPr07Njxqec5YF+v97HTEfdrkjNdhnIte
zEgx9onOxBQ9ADd5TOe3anUVJkO9A/q8LAaUhdoQHOdBPkF8vIAlxLH2G/+Bs5lv
L77AoCe/bkSw3Qd6fI0Z3tGA6WHop0Mp1WWTZ91xl8B4NNYBFHzagtlElyOI+Fqe
yWwG+lOQ9zxcNcMSaTBql9D0BB/QXk+Ut7gKvSvnZSROT+QLD8UAur/84m3kZP6S
fFRnQmm0qFWMam7ekjgYsr6XQbD8QGZqjsGyBfl8aP6giJNTVt02JbEOaVn2yjsb
e2sc9mDGS6eNxof5Uouo9NJbj//l/0xxet8TDxKWV3iQSvXu/RbZbRjeRBpQ3IwC
ZNAdU26kIObC+CFEMkCrUS8Etw2VexvvPbdPCAvF4Lc=
`protect END_PROTECTED
