`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ja316AecA5sUIbGzkQebzmCLB4U7ASndADTT3UDPsRAywq/YBUhAf9O61WepTwE+
oAsXgho3iLuxErh5eDJAjDhECYXO+tBrhYrOTkDXMPHK44R6wfI9Y9REmPoucoLI
oXeTzthOyjBoYDMKlwrMwAqxBOluR5xosBr/dRF+oCupnT0VFT/GOEn7FTrye0bE
+KE3ujJR29mVzxsaeaTDG63rqsuWg0WYim0GtrGzukdBa0yCE96mURqv2faIH0AD
48dcnzFD7+jhrzZT2X8omUgwCz9OJZUpBy2nIBq0eKWeGfblU6TDn/g+bxnm4Cmd
aTtW/fBeemswLGhuXF0Otg==
`protect END_PROTECTED
