`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ip28V75BRerq8kvXgpPAJ6TqKUlYGHZDwEoDYfMv6XYoENo55SEHh69WA4fveSHc
q8X16eboebcVSX0MkE7NPEnIPE/heePJ4JImTpGr3l0EgqlrTTZrsJ4VZ5+8edv9
YvDV7/QAcmp/9jkaGCexlxJzN1FtENv9cqcWwQIkw4RYxThu87POvBThjMlg6gYm
o/TMW21+gZmibSpWEI/agUap7rTVfrWygJTrKaTSSYa9hZZR5NNj2VhwjiFPLj87
TYVketKuoigAzbTE6sLHt21Y7HGh/rTOX/ry4yDmEbFeetjFAb5yZMb3/qOFmXG6
ghbbrYA9pSUtN1ZjZS77rCeRKEhsfAO2r/KpjDSL8KqqIwglEXCpvC8+nkIrcg/h
eL7Ofc5tgsHj3AStU46NQuTVpsd8v4letWTcO7M2OefvdDeP8EN6vw9axNW8+UfR
hKoBlt4OU01pN3EmbftUvH7HIdF088DJAR/FRyLW/0TRWaa6aVN1c7FHX+Zti7Ds
M5akUEYZz/fd5Ndy+vZBvob+ygBR3gFgd2U8+R3uSRx559dtwrDy9dkq7nV38rvf
0ZEiSVB1HUWj+MeHNGXQMdzoX45r/XILixU4CXLJNNAa+D7eF0WOMbXcgRAJIu+c
Tu2h8929huArx3bl4sZmZsWUtRQkv4qZAd1tXu9Q1AoFrhQE0tNhMFL33LuoysuG
Yz+ILQva6nRoXfd/zdDVyEVmmwyqS8mAVKdrqauS9Os=
`protect END_PROTECTED
