`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RBwCxioza0Ir0hGEkNje4fyEZPVbxro4d+wJtorfhASDsI9V72SbD9tdEclK0FUG
g4WRaD7zdVvikUMsE+DqUf6cYMC2mO6Ve/KtGWskS9lh7+q4CV05zgwqpNd02U0G
dN8NcqFdIhe5Lglo+XM5tQeC69VE5McaHAl1rKiqgwRBwNt/wY5XtCQpa9DC8EN+
fgfFZzfKv/vqEBmXA6JmHxa3FvwahGuLQ6GSWVQHhW660SrgrMUpJeqpoznUNRBF
mFdaoKOoWCLFmKDorsPGpdPwN+rKi/xjyL9T4rOEX8mYdfzc9nO/T8NS08nf4wHU
gGsfQfjGE7xEM10oqBTFnf3u5ph8/DbPhiu6QMv1bISxb167CgLyOT2rrHyxT9ih
ssA8gD6PyBxNEfk4So6OCg==
`protect END_PROTECTED
