`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lAVllCGhNlkfA6C09t7PIPprHRpBWceVCVProgFKs0RjXIwHbzJjwo8/FM/Yywbv
/efubVvrJv5RFCcO0kjWfrqGj94zqnxBO4b4kKOjQFtwqFQglHdpSxWiRQwO1aqE
NiFNDLxDdKnGIgAN9vDSs7Y+6yljWaZXaRMcwzjWgFQk44qVF6XnGYQRDxXDg/S7
IWTK5jEbEd4mGfg9sPv1PFKZaosVPrhMjah2dekbGg6x4jjzntJChooyDB1+2ysu
rY/ARAggOv7kUPeBzIK/OnS+xL2P4p5ZA+Z56WIoKHs0ZfVdsj0PGt+yIH/0qP8G
/I9XC/DGRdmjuVYiGPzInc/CAHu8EclkuKn/KtT1gt7vNpXpN10u1WA1T1Z2hRlb
pTVjtmD/VbRGanwY6GLf6IoExBbun2Z9OSweWkX4ejpF39nM1h2sdqlQoBYrkUCt
c+TVz9f2IERKoKFeCgzibmI7LkvlRz9878I8X89ZYxsKhf+QWwMQOPwNX9D3wZZv
Q80wbxDWU2xKUfgOJVRh2LGrx8TZ85Mo46QDAw6Akh18bTTGrzLHkshBfeWWpggF
QW3YVZHE96sjJuuNCHa7lEZ6aF7zGxOJ1d5/dyH7TEEd28wobFjTi6rPmk21B84A
t+Ab9z/DMLHRX6WsJtuSYnhgr8UdCRz03x5mVwaZZCeOAORY5odp356uyxHxJw2x
9ZoWKStHxgrPO53Fer865uUANaL+U1VpO1eRXWZkOOfIcAfdCt620u4ykg2LKq4B
Xex+paRxAHPKFoattUZfi2X+vq/+vr9M8+AumkZXWdlACdBKLr8jCQEUo8S4tx9S
by+ny/vmEY6lSsKiqqLAi8+i7qDCoNV8oMu+PjJVgFnIcRXU75Bx9o3UWODg7ekR
Pykmvy/EokiebT2h/cE33Rq6wS9LrJ1EQGyR49CMmnWm8PbEqkyUCcpV/F/ugTwu
8oaXyat7fSIDEbjZQ6C1mPISdgBapqZGwqLE/bh57YNtPNgedahcaYazvd6TOqKo
adnaRgk6NNlb2j3CgPDyYTiYCrjZBXkhEBpuwClzozeOkjCqRpml/nVUiB6Olu9N
3IduzX03kGN5VSLNcln54za+JwQdn1NYkD0RfVmvbafCVlOkLuLjEPcRasjLNVFW
uH7ITThbVsulxxT9qh3RVHl/m4sNSHZSukvQLhXFuk3+L9EoXFFlVnJJkCko6HqB
sIC8aIsGhkNFipDYaOc7qrhIcbNzvk6L/7Pw29SufSRFzGTVpJAbPF9rsg4UhKsE
AIiQDFtqOTGyCGc/QjWoBCOqMtukQduRdsEm1/xUdYjvryNhTZisWTIaKY0vfxSu
p1MnZdZZHlYV5HbAlXWUYDrzVau4+MKPIMxFzUEDeoC+SzOmpZrqpQ0RgrQlCtq/
bK7MJxHgZQ8JCm4HwbUT1J3f8eyw7VaMZsIUReaUXFuU9Nyr+F8K9F6aPrupkPWQ
wvj8W9TXDey1dW3CgmPF6q4dCv8cwbmggZOXIxEaat70Oz6PZoG8qpLEoBfZhKoK
RXfeD2XEQP2hbnPqq4e+5kvsx4k92ujIc5eL7gf/FxJje5PMyEVh2Qty6pbMhcm4
DTW7SzKDqGSjipANdPvhXV/8pl+1MLRfUDxyvHPSUhhzOVpAvW5sTu6+Tg8vBb9v
jd+qJitItCro7+46Ijsz/EsDeKna3s2PprgnesoMCvfafj4rFgZO7H9Lo2nxNNa8
MWhiq0rCfeS9CLJACCVpqSUV3vcGOsRr5mSlZB/z/occhHR6oDyU1g7d1nCdaMTC
bnFuwmdRX8Td50B0nyabiyGCYd922klovDchmT3utDsXXEY6tCw7tifRwYVj6ZGs
NZSZdUhhwRkdjXQEJYcB+CuglOmaVRUxCbDI03PtLxSXr2Lv0e0Y+1RM6ByGX7ps
0EbItai3chtp3F2MjiZAa2HzC/XAuiMhJZS0UdfKEYwnxfSpULOA/bfyHLGKoQwG
ng+x7oKdcCqFqTsC5FaeLNyxT3W7qlYEgbPa3x39saVzrqnpKGf8Ito9WJsSuF9A
SEAqFXAGK0x6LcG0pTH3kJhfopwsW6GY1TSaEsfkMN7QfzMnhNsfLSh4Mzku1eUM
aqig8/jxwSqBLXvrTIBJNRe3c/slS27GpQOdQOUadV5flNqXwEAuq/azWsxcx1It
8rIx6kND4GtyDlNVpEF6DI+pclA1Txpu/w5VjXzhB0z3s08g1F5u2kAEcDgpDIJs
dls1Ld9qkrClM/mmD1K22ggBl+MKdktzlreSn1QKJlKDqajNGX+FSiaTtbNo0/h/
EKqgZOXReBgEFd+zUhSNQjW78Q43paRD26/CqialwNYh5tTBC/QLCNfarMnSgyid
dP5R1r+P8YlWkSxnZFgU8rs8YVivCqfe9s20xkrvYqiIB3GrGgIklK4c6GwIpGZe
pNj2NFoUhy6SiN8yCEUOdvoTQh5iko83HersJwS+ZncjUGsd0KI3M2r55F00XwXr
Ox/gMosb1kE6W9dYRK3yerW3kr8jpJM7VDktkaQ9wvrmVt9a/jqUWgM6IPkv2fWK
LCKus4n7VT8CPKJJVa5MB+T8qQTILF+uAARp1RtUxc2G23frfNbSX3aH2Ax8VQNZ
5dABEihoIlpiiEoGkiT+wmiOQVmYFFh1P+d3sgkleSxrg+uKN77aZwTcxcNedtN1
hi57Dlnc3jM5S4puaqdzlJVuiNICmR2xWphc9d10NOto1u7fz4k+C2tXkQARKNxC
P5HXuTXL/SVVZgusZDb+lw2+c3pukUJPwA074t5AN74CN2/PCdYkWr+aB1MQwirc
MHNbDDc/TseIgZDsb4lgWGceZeWmXSdR6gAxUZvtNbZ2Ar7tYq0Iu773undxkEoO
+icngONfWMEXlWWybO+N8iNGNOdVRnM6tIrxIHX4bCXR8AVZo0byC5lwd2IAQ4zm
fNE6M/xXD/SCOPyiJWyz4PAZUUxRdplLvV5dfrfYWUXt1qJ7SMq2g46v3YaK11T3
XNxorlFET7R4x2WweuuRscaRj29BGCLJ/zfzs7dvRz/WCBoxtGS5U1XwN0r46Rc4
yplkWeqWo+IeB+kTMJAS7ooudbrBvhiP/NR3peq4+oDmLKUqcr83xUoaYPzwxEgf
ogzu0/WX+oFZfAOov5h0O18AKHKt0NKK56rIFH4u18JN5ZD9un/T5RuI1vAcB8fG
uQj7KfJe2MAEsHx1qfuHFEECmN1rwCCmubxyEwI8NiwNHFqHkOV1ZbZEu/N7Jstu
GUKN0vv/hyyWCKFm6RrGM4+eV7JIFm1rkqEijJKIeA67V5+gouG8R3EYFTvUwF/5
wqs+HGK5gP7T7dg/HyDGh6J0ncIGR9JoExLMJhKC8muNMgQJvilR7vLEe84xXHmu
DI9s6DYJuePfLTM0yA4FcqsJdSbiuwuLTxjvbRUX1MM5u5GP5LhsOJentgtnAEkI
MGyZETXI7JqruEKeQHSWpYwPOF7lEGBlJUhgiMZcDc0U1hPBFiabrKgfzT5BOCDt
yiEYsUlLmNM2w0oK4tih5JzOW2a6wSsNvwyFcC5pEIG9xlofF7FfJrdJwzWHX5Yy
1wyreXiOCKa6JjPXZ8L1mkKYCze+9cqmt0LFgCmLPvSfOheYZTuzkm0RpQey+kkD
DhvrNQ+FGDBzmbfleMycjNw6gO7YSS+ewfiNqQrtz74iWP6Gsi2XnDuxhyEzULj7
`protect END_PROTECTED
