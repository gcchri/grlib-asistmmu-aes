`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mYYFEoRPcGgbs/tY3jGOkHQc8s9JdbkR/bPBP5IpJ+vZQHLLv0zFC1+fC+MiJ2zr
RHIwIMo12DkQV5fp3l+CvtDJGoDtColBVbFPmkCyNhsLnlj9J1MdUIV1Wwkp19gY
ZwBUPgn20At+sbvkVZTnhkzSGqs5jFalcq3UmBh+NtoyZF6ztC+PJZ2UoeQzvjOt
3EGaTo+LkTgf2YYcKswZkSMV7cnbUs9Xryn+/FtcmcFoYoOMIBKqNBwVnqEqmLVn
kIESS3N0FX3jA4AtWgIb8YkAe/4E62S21T55wvlMf+7az4yKLprr8h/yoDE4tPXF
4cxCH9C3BgIjkA0PdZ26iSYJbU8OoLNxQnvPKavYERLwrvVAJmvzfpxan5TDPp9/
NdaDskHbJ8XjtcvDSlVOIq18NzyPiDV6SnyLnHU77gAeWUpbTtWZ2K4f6SrMCW8H
uJOZCLf6l+uJpuGoKQyMuMOJggxllg5vaNadgaB70eoHWY+whNCUvqbiHMfPOHrJ
79rRdiw/lqFrP+Q8pzNlfLUCexqJSY5QUum8QGhm7g6VfdwQSK4dUgysVYjUtkd3
Hb/q1BgRVd8I4/g+qqJJeEwbMNMZxldp6duFkeRRJN34Gg1HUTR3dUZSCnq0WRxz
RgRWR+Q/CL/HRum5fUcOMGeM1tmI7aLrOiABsmFL0EGrK5lMebq+5nI8wkB0lV5i
dFZwSxDbs4b42GBiMwSuB2anwJCxVVvtxx4oQLonRICy00KpdpKSw3pafrXGKFDk
AYxAdL7HFqpOQMWewT6PG3cRKonn/BVVtx12pe8+kYXO6801o+c7dvljGRHUjHCV
xYiV2n/2pIrkQp/+FYEd254NcDhndPTFyb7+giDw6RBm+btbxUvwmeESjBxNfKFS
DxOllFkMh6x9zDizLEOYMq4jyyDPlt0qOZAF2M8eOjFw8M1WLy8ZURQ7GV478s8O
m+qeMZKI/yv+fqgPLnjT4FaSveRbU6oBLclnHWbovdMqf4wC3A3aV9jCrLd0hnG8
UOilBFpeMUv6DvC+J0aZtJvAFqLwz5+TdbpUdp0YnyGKMqtmsX4D9TzRWavWE+2Z
85pdFt/YNzaBvCNxemsb/iHShfxkErYr85JRmO02AbnfB859gKDne+Q0tO545V5q
BrJMIAMngV1tMf3QJhCfjzrYQPDiNLTik5zWK1aVkQO/L2miU1dS9HYaTQNAnSpC
b9hwNb+Um2KGF9H+CEW1FaJIg2sEHLhYN+87OHLYm1w=
`protect END_PROTECTED
