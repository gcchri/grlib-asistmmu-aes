`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xOIbeGy7NRuKNfSg46TRpJC/XkWJJ+Yri1R/ABIGc4KyHA2sItJsodoy+x7umPXQ
X3UpoLT3ArGcMXpjyrj0rLfaikiDYoXF8rwAEKOwSOfr7EuEUTcOi8SzBVZQU6N8
tL48273D4zGCvL//IUe88MBqGn8oOqa9fJbRZqX1Af8kamfbdskFXgPmr2nQ3SQi
CX9P95UXWTDKA0CAPzStCK322gzUIZStT1Y71ZvBJIWCAlpIT+suK07ouyRX3wic
HcuFm5awSY5XDqzEjjMPgBUtyjARb7o0W5116DUpHwnxZh0V8KiTDd6ji6PMndtg
alhsLDQ95+7S2jbIFerXgTMbGBhNO7h+WFNw3Q/Ic+v531KX8Ly0wQ4bKzMkFQ7+
K1V7E+/1Dxigod69HNWoBWxRVCxS8UwYI1id2PsfVC3VDZO3gYJiWIm4bDmPvGL5
6YytqJjS34QgN126kBhydrHpnutbixMN5Nti6l469xr3BaXsglRG8iOXT/1sy32N
LZoO90THIOh05pRiWfrNvGfDGRFrNKiVOrZM3wArCdA6FVIxg0wo1Db+a6SzHtsp
imLoNRkU6NtuAUmwLwju4w==
`protect END_PROTECTED
