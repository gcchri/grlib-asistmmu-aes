`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ge+mJZxRn/nLUs+ezQwQ0w7F6X4kpwi4DDzAncCryH4Z0AopMdPb2KRrsijGMdgH
LW/OQ3OjpOBWowwm23yyIx4qg3Y7juxXe84eZJl5YS65AuhRvIlqIJdCXe4sHouj
jEU44z3i7fx7YFfEHvliod5V07FbuJLFG4QNNkuUeInE/+lOz21XjFago2PB/FcV
Y/zIOklUubtEmJC4H2jEY4IYEJcrEhBMRhTGucTyrFuWADXneVy8IhXZBSKHckW8
OM1P9q9dEn5Du05v8L/SzbY+AjH11OnRP8m/aFtCaxSnwvyCIURVqku+w8O5kqrZ
LppJsQOxIdvlHaHB3nmJ/OW9seKCM70f7RZ/eC6fwawdztI6ktgRl+p6QBxYuWqi
h3pMjGtyZJmScLeXhS54NfX2+sags9AUKuTL+AY3Yedv60bwPmTXehef36QIbBhl
5ZZwwIQCyggzyYgePX5uzsBCUyhJhxTTRqY/2JICtzVXPHlrahL2dycf4K1z9vNA
krPrHHklzGqH/1vOl0EfDjniMb5m38N95C6aJWfCCi1qdnpWOBUCVhN/tD2aAcpj
cKbw01fg6H45MFjFgmIxh1sjHDhB5GDBQd+CvO+TEFh6YIIzJon3YrD6wA85Aho8
9+BbvarcoCrqUVTCJ+8h7L1FihOcfT0LQXLQSfofwmFsIJgLLuqHbSHShLLLKiVc
j5GL5GHqfXwL3PkhqgN+ddNmcDebmUJYTfXUhrVZz1V+gh0Ppuv9KL4gf1hvmbjN
hUklRxu/x3JYGS2/9vKRJxHBq2Kh7EcuIvpKRP3P/FtSJMjg9LXE0ec8yMPNJQg9
obyWEG8UtZzowFCZXLf8rA==
`protect END_PROTECTED
