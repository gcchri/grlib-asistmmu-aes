`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YH8dDFgdbbNckAg1YUSzUmwMjZ6GWx8YKXHlxHp/Lxo09jpx1iIHlgpDTsSeAc4B
zgDycHfMz8ZSfSsmJeGmh6KQnqSWlFrGBd3usa90MEH4TClMYaSHRHeXpOmXaRie
f4LOZTExL1QQz71rxLulxUMMENXjbvKKL0JWTVemEbNA4wr6W5fJ6yJ2FXh45tV4
j8erWAusZg64NbV9mx5wwdS4app2hUE8wIwVUAv8EwG2Cilaz86V6v3W0ygPejR0
2DjJDQF+K1ysQcWgGVAf8zlCPTyELqIXqiNeTyC3ilHVXZZrhU+h8LDsWzMDuGpo
ydzlRi2pLzSjEagj/7Qoehuyl9RyvQQucy7GilqA2bmK6wasYZi1e42F7HtYgVH4
`protect END_PROTECTED
