`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aY0EdsWPxI7U8iBWeCiwXTG9DxuDi2zyihldyGEwCFJ/gnYDHW3uJF85dlb6ZKBn
ma3dNRD6vqozssCH+3YFuTraFHet2dg8WfLLg+Rig/U3q9k8pCNsZadYa8zO87BI
hj2oGhl9DeozYP+IdEgTuWdEwULTh12AsuC9ZnCMncIdQNb0qUYS56gCMedSVu6E
rZ0JRwxGYHtKFozWN9028ogc5/eaadhT8crimtphRTdQAN2HZ3vVuWUuBwXY3ZBQ
g5MBVfexNbicbpzKOYSXli2jp3cjry0jkWF0CRcDfKad4JulZSxv8UymR5PNXWP9
G00OZW9Zt77z7FWktdBdAt9Ww2PPQRtGba0SAKxsnrhIIzQ2u2WZwm8a0lZ7qzoF
jTLSbkfSXp3kJq/bPQaARVbGz5DJQVD5XB+bdS91r3dKB6ee+ALSgYYU0eXu4r2E
6q+WS9rL63tVftw6Hk+daXwyZXaCcuNdeUw6tCF8TsPAG95Nl2h1cxFmaHRiVMy7
nb1BYgK3CQEn55NchafCmUTtc9X8aVGgRlAemKe4uFIhloG57ObSZ5pmG8XxwATd
6ijxAzRd6HnRCp282QFOVLV6xv3wLb9jVHV26x2RwHlWH0x75GIHTLy1fKHETxsB
VNJjyDGVY9YpbefWT49km2eaQDcTxRCwe7imgkibNrlZyIpqUtsXxFa3NTyvRQLB
Q7dSmuiWgsZQ82i++WLO/Oxaco6pp0WgYxmV5lLZA/RNKvPwu76kL7vLq4mpkhCg
0brWQYc+22jHpxPfniygK1sT3rYEpTW6702o5g9Kt7EviuFz9L93N2D4DWEHsbor
7wMK5Ek0OgWnxYL5sKMtpw0MrHcAsxjDqiLKDYR8iJhOsS/5uHeOpC3d150eoSXW
yAvAXbvqLNFaGR+RgncgPCw6zH4cgNxz8dN8wxzJNpDVggIsa9kYqGj+WyjasRXd
z+ZeitW1qU3NAMKPPoKzOaT0w5tSkslbqm7jYm160UgYc+Bp5zWdQaZv7H0e/6qI
ghF80r02bpf7k7h6DDTaLQp541YuQN4f/Gq887kQovhHZTgZB1uJWepJWI/xqQ2E
w8AzN9dE+1RUAmonbLEz0LVliCzY/KsBao5Eaw6nGrYb64PmkSbJ225szCAA4/5l
BXalwTA9CstSgU0y6fHsmVw+KB1KqSAf0b4UNddvJGT3iguMXvb+gSi9NGJMoc8f
KL5hsRE5Hok1yY1A8zPq5zdgbiXin6uEM7DtHf6xAJiECQkgPEMzvYrtxZYUnadH
T+htLZU7v2qavBR/G6LE2NZu6hEK77zz6gRCnFVNQWqlRgW//bAvf1hnrEczV3l+
BgbENHN8tY8/mJgTAKaEtp0IsA4JsdR1IIUCm9dK1wWjOvLaTsj2B/hTJe5+6xOx
iiASpp2zt4QMsRbJ3jxlO7vdJ4sOBekEVp2NsaSVdYgjYgiUTksydmiw47eS8bo4
1IJ9XCt+Wb6ACp3VC3jT4sLr0xQLfmg5pCdNQ3G0EG+0v7TK++kIZjxsYiyzRfUv
yDsfzq8jLDEyj3sVfFn0PunafaQLkBbwV935lekz2TXwDzwVi6qNKG+DI07YWPYw
Fm1j6EiQ4H1trRA3/NUWJKB13UEEj9LygmRVNeQDV/2+3NKdjvMMgAkwr9q0rP5O
OEwyt7gHKaji7h5mO7YJANkXsZqLyzaiqNLbu+Epzst9nogeI37e7gzWIu9MKIvG
gZA1bUxBHZAEeT/Gu3tB6CkS1ljRTZqBzELS10Gez9CJx/KvtFau+okxdgJNEn2d
aBFHbzBAAQNrrcWPkyvHpTOzMil0Gjb5OScpN93O66VYkD9TL6FcgXrciEdrGX47
Kg5GE7+qm/UpGOlzyFM+vZMrLH5isddfkFEJ27/3mw9nnkam6xHosdVz4lbGOcYB
ICawNXDyvc1Hb9gcOHtiVyztEClMEzooEVnzV2yezWVHEnk5FGLDhHW2LVxwxUj2
eUxuRV59Ii278juqveoe1NABXNCtDVxmepPfxRdtxpBxyY1ZzjaBXwGY69mXU3w+
bk76utwBUABYLC1N8zug7Cw9gE1n2VLAP+z5KRtfmgZ//zMZSqRjPedsbOg3V48C
cJLuL0BUwl1lD/1jiwOBfa2Dm7gs/TVMug0iA5SMiR3yBBu3iKNX2HnaOYajN8t9
gcQRH2BbWSV/sEIgDdtr0NQN61E+jYDLsUpYd/4PxqVulsyomP7NypCF8J24C3zO
P45e/99Kl848JeI9s+riWn16gzUKTNqW1gSIxvza7R9Kc1aYlXLq2Hx7KT/forhZ
iyaGd05Of29PcydRlLq7WDvbOVjQwV3XY3sO/sgRkuaDucObwbK/L+0sKjNw6viL
yRaJCN1ph4E+OCk3vMPtAZIqs6+e+tyHiezqJmG5gT22kai2LwRKAkV7+GzFmE6b
Rhlxuw6QmROTJau+KCTJl1/mDsi7crJQzzgxN2KuUsvbuvCzCmlAl4EuuHmHC+LP
PCiOL8f2KWc38X50TT3iYFmsyQi/PbBHTpySLAC5lHrk6uIe+U5E6ikSDsdnIIPz
JPBvQBQIRDIaIQ5VI1n4a2GhMHAVWVMtCx50f2/Ma1qSObXrg3HxOaAvgvOSR/HX
Blmy/ewt+YLIE1S7+iyWzT1xG85gpyGOfy2oyErmk3Tbbe0rDfd3MKDBBrRc7bze
L53yyB2pSl9Sk6zr+jWy/dwozFRQ5z4Lh0gVzdSAqT6ieSr9eZdyEz3XIKrgOY16
PSxRzSMJOT6hsmsYqGF4UiZD9YqN6RjOWwwAN8kdQZhv/z+hewg4NGPl/JgB5n8n
E0N9u9hjN6ufKM25yh62RpY4C0bAEt8G1r8I0Uj6X7ZZMu+Plwv8ksyDvqFtsYUt
IJEBqzJM1moZ59NJ22m93MJzymN22lPnrEzBWO3m96M9E1cvTNILq3RZC3WYFN4t
SjfbrtYaRlzu6CyFlRcEJ5yXw31AShlqS7HMciJ6wmK3RrlWcD9Q7ZDV3BYiEbxi
y7fcRlYCjLrxnzETlBsJNVDpvoGh0lQ7z4ZdvCnPnlJAgG3Uk61xW/sUwNCCqr0n
+dvqooQpkPfZkrcU2Pv+1vIY/GDtwObB8/RXwnQz8Lh4LCvfTiOO7/GiJStchLXF
aQfDDJIvG0Qd0J5aZjvlQGxWMOTm2vX/Ox97F352edbUVtYT7/vcXcX5pOK7vLZY
UB5axOPdQdUGTCQirbBn4BhpC9jRC8x0vKaXRwEOGU6R76u9SgiqazkERiFlqJ9R
6IeZXPyhNf40uExf7xsjMQw/9OQ+FNdJKLdtxBDiNlnMCRIYfWQrX0XByhPs3dwR
GCDgSV4nEH81xkY0dWBvGJZvbMXjn5CFfTU2iXWXFkv6Qv3VqeODYJhXWEdYFTnb
Nyz6/LcJB2e0hOAn7VlLmHuVnR9/E93wRmGGp/+Iod4PReTfHGYfp5LCuELZVGxZ
tkb7r/PZ3eH/5TxGPcuiEvbCRJCNqNuu5ReFOnwGAzG70ZpN1y1qWFLrzZrFY5Gs
lLQIPXjmpIcr41KMwX11yUO2SwBrqG2HjhRJ8k3KPI18tHWlaOOA8/e+h4qIoue2
uKwkKyd6m8UX4k+sQlFsacstP6pokAMVT+AaVBxLz5g=
`protect END_PROTECTED
