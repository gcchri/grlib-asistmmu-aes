`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+GO2Jy9ksr8rVdxyYToJPnbYWcJvwfLfpT65kMeVBRQGLRHbBOYh1/jpsfrdXOg3
tLO7LeqKFkj10DS+TjkgCjaRtmesAayZh+TRK6KZoBi/EVY0GIklYFevenT+XwMY
cEEJP9M7NpPmJVDqckOAaCeNMeELOlDgUiQ0m2B4wQhY/xXsHPvaT5jbN4PCG77A
g3rTdVLe24J73FveUExsrCFETXD2nUou+AvhjvqBQwwAOpWwvERT8xvKHJVfqrVu
DrDVnFU9EChE2Mpx89ODQWncMaxzcyDzgWshM4XGXq181yVGDr173h7NfJLpBDSI
tTOHvPJwYNqVN/sCnDAfy91SuIR8CwvA2eQD7b+r3xG+gCXSb49E5GnxOUGitrhJ
T6gjpXJfWdstjao4pZoUSeLggEfSuRX/c18kr66C+XrvQd7JOd+73bR+jVWooXW5
0GRnoZPxjIsP2a4pl6++kEZLPUI1SPv5xF8fgt+fTdogYfykPuLBffKVW2OFXGht
BAuvKUFKqvUQ2vbWBJndwBQhRfeavx2kaQO2aY5jv9ajLQi3vLsVqdGZRoVC/L0O
jwk1/Ruht3P00NMnKz0HD/Ypw9LRNzrWQmaVVDmspqQdyoH+/ptosYZiWmgWSg7f
XIWUcJsYpePLkTYb8D8Z4g2nL4SReSOk1rvPVnelAjFAGrD/FC3qnrHdb/waJEE0
z/KEJtOhMpcWbqMjS5+G1pB3QobIfXg31Gk6Y9WGtEmX3Hn3OzzwE7h0iWDWyQzj
laxixLrpzailhLl/KAIt5NVpsiFpX3+76S28wG1fF9CNPj1qwN9tRrLtAP9/ZxEZ
r0UM73b6EhpNUJePyAEngvZwzXZfsziLqYKhLBTIf3Gg+N6p/y28t/DgLQ/b8lor
ClydB0Fl8wHWG+rnkCw8NQMDQRQEHLLbXd4EGiqUlnnaVDqaF4Idxy+zeMRBk4cj
gq2ILh7LdhdqbiP1pMjCTTDwq8u4/HUjPM4BfQJkRmM/csY8Vxti/N1CIpSwfdkF
qpuaFlvQmgHEUyVoe1Qm/EnSp8n7f9sEUEw6XoLXzg5PVh/EX0z6joVvEmV9Dv4n
8sytKSRDh1YTflBXC18IBRt9XuIu7pbcL0Wz4vTw8VRcV6CjN3NNMS05pazegT4I
Eg00JEaKvdaYxIUjj23FkXILoVp09OYfuJYYdVChSRS/Dku2wLwxoA4SOciQ/oYo
zcVElqYAxoW29BVYu0nsQmct8Yo2AvKi2FRg4q6BQwT56gAZD4LJJaKTtNxk4BCz
`protect END_PROTECTED
