`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nEd8/W6LjFvaiPvRnYw9TEXGH4WJ4rNESvRTbcA3FDnt+L5tbrW+Peszr7P6T5Lb
5jujVfvq1HSGqqlE/+0mZEldAIpEtHHxjqvrnVnbrRmXJ/Xtt6OYXfiHYXRj/ZUH
fGfmNB0a73roZaTdHUzi59gTYaUXs+6twEq/dIeE+AyOXdO6FqjmxlKw+oXj5LGC
jWzVqHfDYt0g93jvXu55BMNXhDdqIB1m6weffgNd/A7pR58u6iBN5utmNrmPp8Oc
Y+SC53qlD5EFgYZmDaCaMQ==
`protect END_PROTECTED
