`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JZWXk46U90dIC3LpSqoUaVgq5toUcj9bqdVHJEXz5cbak5wuep2Zp03n8b1HESM9
B/qIKejIJcSqMTkENYJYYrJXtu577Z0GHXaXER8YCdG2bsvvAvIVlXytoJxQcYdp
YBh2/nYx8InJvFIz48I/hvYhMbOcrm/wayvSBWtHQ554d0OioeSim/h7Ru/+x4Px
YDQM3vSb7Vol9guT3H9HjiH4Afxb2xq1KYixEnVqxD897cFVsIU8AaWxhrWmo241
YaBPf7RnStkvA6DfF1rFCGqD29U5TLsOoJ8fbb0HuqGM54Y3iX0Mwcxj0NbGbybL
rNIylHftgPtVakRNeYSggqUyomKnzZKVy+obXRpnBcjZ9qy9fybzXPWU3bEz8Rlh
Z6C6PlYXEqqZrepdTpA3kEK6ru3VtCz6VjuYTuIJnX2ljGFnJN8IGClXvAgh+kgl
BFxGDGnL6lElWXx4gwzmOgJoYcT/EClcBc3rZNJeM8nBP7KXsCIY0NzNpaRqGhJo
hLnvpndIMfGyZSak+5oFBeKr7TyUHsL8GM3wjbqsboYtOUZrRBSohfwOVB7MvfQp
9+aoGJsTiPzYXAf9mq0e2T9gm26TBB+tb24yvGs6REQiRmmBvfDksMbp3OAGZPVq
qZlLtzk2CVomey9E/rtMNA==
`protect END_PROTECTED
