`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PZXLmdKy3Mmf4ShFyDin42ssPoKehJxIVEjDaqDOIa7vq05QDOSn9mZ5CY7W470Y
3cUWeCMqtNiKzVT+fAaeT6CipM8s7Nz9mkWlw5ezGFjNV8c4w8gzkSHMyg70N2gD
KG3zEXNfIwPhq5yRyF4WCSoDas8B/prG0RWYA6YmZ1dwEieG8GPpmTKyXHmecVCu
d6uvRFLePCI4USFdctf52rSGONbS5rwLxELm9yZbvZF/OkjzPNTYDUhXxuvIMGKN
SjDzgBuG2zPtCeI6IEgO2bna8IVnCjHo6n39s9Zw2w73a5zww4fvmoz4pX03P5OW
1b9eZDfAWJCtFdlacVfLMKwS1YbeRoIyDk37RAzy/+zT2V02yyQHNvhibLc8fhl/
M4Ny7jW2zDuEt7fJjjLwtRIMoyQXXFSLvPYLdnSA4yw+Br+QEvl99U0yY3mVLQjk
bwF7ydU8ZCe+xSfy1nwT3nnFXhfPKzQWA5/QMTR+Do9CrZxWsfMuHeyOarOqOG6r
WivTUJcRxstuZVUOqnYbPe99HB4EYQDTzJrU5GrQn5EM7fjQWQuhMCWOexEPK2T3
/vwV16NtxJBLOgSlg9BOQRNONoSEWpXX42rukkK1UegbzIRmkwhAoQ+x1rjnzhjb
656AuGa3B3U7pzuJ7qjkk6bd/gF+hEKV1ehoBvcY5kPpA0wGQjB7BTdHybEnRT9F
ltgX0lX1cpQSVzE1T2xorcOInnS1nwpooQEMLVc1yI+euCaPgJhhU2FJkIgFDXTH
IZzi5uQ339R5gNZexMjre/pOlBBSnx1Yx9kbrOQGkjkVT0MPhINUkPuJ9NzjoZHX
yGF70nX5mBV794+8wICmeM9tRh2HDTyxj1v+Vy9rS0Ndz23crqwCOla995XgTrwZ
W3oaOIQk1XEluM3xk7CUqu1NG9AZ89TEpvjJypag+khnxIEHJBrxY8QrCVfRw/Zm
e0Gij2OhfTT+398Bbx5Nog3jcyR3iObUu7O4jlYlN90371ikljcPsZpGrNeBviBY
LSQaMYXnnjqTqYYzs8wWuQ==
`protect END_PROTECTED
