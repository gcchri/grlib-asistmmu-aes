`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZazhP+1MJ/LDRvuU4XlYzvCdNzYutcvuzeOWdFB7ya+YiWulMjrp9f19fg3n3W3T
uxqK52/WdBnpj1K7JFlHzOzZQKFSeU9S/7QbEfQykUkhW19Kob4lHvnQ/MafiS0A
xzVuXLhQRWKVrNfr19NdxPJw8yATc5WVtCHmSOR5NFJtw+msFTKQ5jK5W+Wl0M+x
LJFh1I2ktS3iJGzyT0h+siRQKnfLdFym9bq/HMSgjGLrZR449JQruECluREhRpuX
XjOGleYZTHEj32HZP7dg8FWuQd8tx4U85Ft2alKy+3iA7QoR6iIrhmo3DOLGqMbc
IRVR2d+rhzfE97hjtW1g+tCEXSK/HZrf3nOOhrOrvhC7eH4W/9qRbNN5QbH71ZVE
sgGZT5s8dBDYz5Bwt9k0SNJ2TVfXbgViqd5HgNThlKcdgT3IlRBARYKNzXauOwxr
`protect END_PROTECTED
