`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2xubSx9DxNKAgKB5w/boG/ABlkJg16hbZ9awhKNpv1VlF0JVK3WmzTUw4i0nq4gX
s2ZsO2NJ9BpKxU11LCLssQ/F3nqA+I9U8TJOaJS9WlIrYbumq90CbVs9ZemfUtmB
jtgYtAy+ULbhISlp81PNjpr68XjkIgHrepbH2eEl/8bkjHJpYCJrHVz5ic/SmD6W
lbmyH63b5C+BQLfa1+EGIf/TpQUxKgJeWzWFdeqKKqrTz5RgOMaMF+AXQzpoaJ6V
JC/qSErMECjY/+JZ7V3oVqorulqA7Foeyaa4KP12AL7hFiQUKM1fG6Lj4/Q3WQqD
wCL2ZO8YoH2T2hyBcHRDCrvT3o+Ecf8/BnLzTjOMexW6LV6vj2+vrYtEvtvdZIrJ
9rc5Tg5w5bZoJ6hRKxJh/jn8ljlbkTy1oWXcIY2qbc3DVkE0P9HXB1d2f5gW2gT1
ssnj/mFxOMtcY+ekAzyxYjxCchlZp4ws0xpVElzJ4URYeDNmPZi0I3mTbyHTayDf
PgvHvUYKWGSZCBk492vSfLctpHLV3HBvtEcv+8GT+RWg0yUqVtS3B4frqhVHFIWF
AIJD31G3FUCYdxHwlHm64VDYN+NxJRwS85QtUqh+IQAi3wdVRhNC7vOWSlhlTvke
NW2yBWuDStbDxZ58be1+e9BLh2ve6YRMso8AEm58fWW9YK6P+f/FmyaejyucMlh4
uYFkv2P3x6W8oRQW205RSveFvYxWPuTRllz4aC2qhyv9t/EQq6Q2uf3aseJJUVAE
jEa0yEn4xKudhCPj1fymn+7n9x5jZnh4VxU+C4w7c3Z6Uwkv6uJ3Gz5UHqLfa7aZ
ImWYTLXdE1/lijPmh7ejL28JawlnQ5Dw31DSfw4m7A0=
`protect END_PROTECTED
