`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Aj2ryCqSuLggUXqgjJMSmZuUWQwZ/x8I/wFxYb2YSsku2itg19S1OddzHbx6FAw
d44ebCeoQdHx3vcWu77khev97d+C9/en72JC+Bq1l1mtAcV2/VhKhm7ygrcCNiXn
kCQ9ObhgWRly4vzFP5CQjo6KqarIhFdHFinO6y8BCJ1jnvQl4WhxbSx3KxFb8o0W
4fDvW9kvo/ixPva1mHAfJwGRFrPWIghQcM8JYC3SLCl59Ezdkt/4rhL3VA9kBHUu
Jvk/Kf5BdEaBPaqMYeeWlxReoYtTyHLOwXCKkE4Co8m5o6zU/xR8thN2QjyDQ9Zo
ca2HSYftmbr7q7o6/vSjs5hjas1D50KRfu6kPRUU4RGKj5YqsNJ0sfxviud2eOeH
q34q/EgHY2zbUjYXGPReTUW0qcEoZLPP7io8zpneqNsQNPpLNIDLXj9Pi38E9Kqn
`protect END_PROTECTED
