`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fTJoQuSGpvB0493/nZ8nN+ijUADby3LIITUVGB8N2FKTNBhzMtoDENGfwYw0ZtQn
fVq//Ss5JRL3uoCj9acrXlpFAmdIixagNoxZ8Xig4UtNwbainNrht/FwBsHjMUd+
JrMWaWJCfvh4jy6zrIOvY4LF6JEsOkevDhkkcjQf1Rjyhakhmz+ty8q/T+qafiSU
alt0F+WwI4MGpN3VIpPcGFsxc3YFloh1Us+e3JYAw/J5lrvthpSCwwMn5148Zr0M
zeGYzIkzmj2JjrB5Pn6J1CfeAMTxvS2X1o81wnaKKuKDUweHvde5o4SQ9BWIvHRX
sVEtk18U25yR9Sd0rh5Wow==
`protect END_PROTECTED
