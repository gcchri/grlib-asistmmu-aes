`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ai2wVc5HcVgSloCwL8PqVEuzgcqtLGa4FoSxmshVgG4TKTdfRHVcbkAhv8UqrsWi
ls4jtFr/+94rp0v6HN7YCXcOY0Hfd6+ne3K6WRwm6VZ9KdvXZ2aSrHJkyzXh13/x
/b6vSQ+sw1SRfvspAMcVErR0LkFdizQZNpzMCuU4JFx6uFAZtgcdiu3oArMqSNdT
sQMYgD6Fmtjo615fSO98CK3ZrCPCTojFbFSyohXKC/RwZ01Ua6KSVjwg0DrU8Oic
jegye8yGRV2IKt3tt7zSrt59nPgmnZRqYMaJZCvtpilamM0Fv6HxzKwmJtlnVqEI
ZRI5eBmpDdxeoCZi1rDLLnI5yY1vAvO/FHLY4yRwv2IvdqTS64vxMvqnpVJvns0m
zCG1Lcu5dWwJ6MTeCO4NUQ==
`protect END_PROTECTED
