`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AWrbKBon0dT3qD8JYHDlEMUcp0AAr4gfxQdQ4FwawqJefv0PpeuRQI+7MBFfoX9H
iVKNpsPnOuMw5b1hwHmuwb9RjXH3xNExkTiVt9a7Qacrfsty/ryaiRvr1P/+Zqu2
/Bh/cr550jNP4wBvt+iYrsoX63QFeT6IzunQ3Qxaf8+OVabSRsrIXL8+vEN1iBXT
S08osWDmjZaVuTR/EspwEdMgwqF3hCUzwNWEJ8ocL3gOQHG9/T4RaDADj8gcwxHr
7ZWf98VG8dgAWwkZ2AOqhtSlsGETCANFWgoHDb9vzD4ldN39oWKAg0TafzyDAwbK
5RBgJAPvD57voCyW2U83nAlWqpwc9+m35YAj3YBTcrMWcgtWNG1DrX/Z7SHohKiD
RURdRnchz6XKjRIMsSFUY7dkcMiZM/l+E9SNN0PzQBjnb4ToK2CQP12lvWNrPesT
g5Og707joohoSgxiEbVj6Y9LHKCqDBTDMrc5MkKTXMxMWFp1Xr4a1TXXiYEd9NYo
gBYNy/HzTH3BZc3CKKs39KsNK1e7l/ZXdbkHNtCEZYLn7XoBsf05GrlL3bnp1a2w
Yc2w0YF/ruqyZwXtxREV2mOvIAfMCj5FG5aqzsy0yroEHeV1p50RadTCbXYJvBI4
T4YUB3+o+FVcdVD0ks02DEdiSQjZgsnU4QRe0viNb6AoWn9eshgCvOQmxE3ZpzQ0
zbvVhyuCXZ/gP0sIX5rjofo+OlVjq8rzwxBB2hQ3pyVPZCuNxgX2bfQbzXE5tLCU
3gbiJIz+z/1nQcQjEjZKrOx+35MdPcniVufeStbVQ4zQPP1zp7AbtIEbITEPKgO3
9aMlXNHK2Sj0BpCllEUBZ74gwyHMgX+WLvQz8iLE3aIptkwqAUIMtT3jc6SW6vUJ
dtwahm8VZN/nvt6lfNoy+no1P6Gw5N2d79P3hpVSrDWgqYlqJaAxezV3GBabFea0
Q7cHNey2XM5iU5wj7YzL87+62sOW1T8rTOXZWH+INcdu74QON+3p+tKmOdttAJsQ
ZXiDWX+zAkBpI+VATQXdzwhw5SUsaAn2xFWieTJjEidqEl9Nu8Nk6IR84yl+O29y
phzmvfluoxtIbhZX6ifPhEWHkLbFd+29hxrWQG7GymlYp/B9TuGNrfrSXkebnCfU
WG20Pyf4KK38CcpgXcInwycLDGFhTwSaVaL/ZGmcOMqt/hX3H0iIRs+TnIeDp87B
soHrfcSYsPWfqmHRgRG9hB9Yv7LC2vAu0E/r4Q5E/X4M62S+NhlNZEaWAZLbuduo
4bS4m0nMoC7TbT9FvdzOuffrmZ/0s/Uk3zS6fDWHTFxfMzlXW3XQi36PbRW1VWEI
7gKoMVHeuP5SqTp5Hy9Y4bklgvXSAi71ge+D9vXuQ2GUduX8YKJ1b8wVeX4b2dHT
hqprLvqugNtrv1lO+g8qEffHAza7NzFrSjX1w0dtRA80yxW7UF/sXLKbe6pwuAtN
STwz7E4T4nz6UJAMq0H3KI/y088M51udELuHL375Al0MTtU5rc6QQmoj/ave4zgy
NMCtAwIuGKtQI7bQS1sBGBX6CHvIRNUr/lT3d+OVw1/CtMjI1Ll4bcMWoOFer+K8
YWPvIxEAKcwOLqIY39NuGvuiWzEJRQMUvCQUTwHrGnNFp70hUWXHHlEd78LeOdBG
wclnO+UTr3nluNpV1riAU6U47F+vOFA76cbQIcLZ//T1PytrO55/hhmU5Y1+4/7y
hi+/Zh2P9ST8g1SvYjzm4Z/L7AZ+53pAeJHW0NB2Kt8SNgksfCg0mVnh0Axo1FOL
cffJ0Qy6EGCflWw8uvwxYLUWummKFoA5S0nQuAH+EbOazF+Kt7d1b9hnHkRdPJe8
2lF8gXtUE4VewFFhREqU7jg52jX2kaAl+BqzBYAfHm5vXxvacrjHf5MOAgVjnKU3
lUkX73g/NCXMUaWLhVm4nSh+bVCfXccZ1RXNI+IuFa7g6uCUyyuALN/WhpGYZAA0
355hMI9U9vuv2fwbTg6cfYhMC0vHtiRc/y6ltFkhhf+0RuHxX6SrIGicuPNFob3w
2n5NTtRLHhSnEi6CyysiW1D/zIs9nmoXqnqagk+swnSnPioPVP6cyK41vDypq98c
afYSM5GLUP9fYnmv2QoQwY01Vg4CJYx3CWjkGaJC7ZN3y71+zXTLxD9HRUVSgm/M
S+V1Yn4X6LO5EPQJjUaYNOuLUV+F/psajatzTgYxAUU4rZr5oW+k05PST7wkgyu7
IERmzTGoHXWRAwYnaS5gA7SnesyKRmPz3P4zrIv4TiPDhYos6T45CyG9kApu2IEW
yca1RDIxiEAnUhUwl0zeUDuTiFTnfDcp/vnN+wCu6UzBQKt6fadtDdClJ1b7DZcm
SXylXTkIqdHaPgUXhIZUhcme9zCg71+RXDxC53ur+m9NRBGIYE7j5WZXsRgz19bW
dZI1fFVJD3Cd/QjqPOMTMhEAXpAtHOmFXNmwn44jSs/M8nhCyhS7tn+nbRocAacW
2bRvKcb/w1DqWzvu1ZvLsJJOwLHoppHUSchFaG/2OZ2LtzU4zB4Jj0ZeQfAQRiYU
S1gRAdzCjdITAgi5Fd1iRsk3WyfMeRvKVcEI8oSdFAlx5gBMHhoErLEnK3Qm6aD2
jZdhPoQS+UR0BiWERtAR4wh85mA7t57YI9JMpfSsC6tW7Yhv4eoUT4av3VMrrZC5
zrBy1yS59HWM3DoBxYX+7Rr2BnO1AnhzQm9sI67D4DT1QH1KAuXmQYS6vLzS6Or0
X55YGG0uWpQ1MB+AxFeySwMmB6uE/Jwqs5Z3a5S5PGY+OT/CiS9NLjnL13atJMIt
8aQZ381X2gMA+YVNsxVJqLOQZ11y8iWi4og2kkTLopeS7boHhrbvIKGF15719uBT
LJpBDhEWdmlm1A/+Mk8GMVNBMzoIA2ZtYTb0/CoFFXv1p4o8T+5iGk524epHEE0I
QoXTb3Wo+WLluEuRFEblPRdMPncd2rUsmaTUIIDokNbcszyUvIjQl8OlkEM0SWda
3PE4ISNYpfOz/rwdyeqB5Ywemw81CtLI2VU4LCtFq9GvuqVEFsElX3Ryqw1rP7T/
oFqwf5cr3LuBF9wBQ1kyNvwig4XKC+xjYptsWwYXQGiLtv3YDXjBLt5V5QQG7+IL
W/q6P6JHmGy1pBa/7oIKK04j7PolgdFyLR4CHEHT2DEI05u3lQdSaLGwA5DyKEiJ
6YA8IcanipI/sZ0A8xQeU4glJpdqlom2yyjJ8/i0k7pnQ7YFxwkof+NXAszu6rc6
rQpAd27S4dakmIiYZ6t8yZr4dXsaT99YXm1OFQywWiqRHIPQ2ZseIWC873AfNJBy
Ol8uDwVE32kMZbKKQU4BTgAtNbpSDBLSlKCHn2I9Rcph9TuRXlFa9iyJ3qmSbpgi
+UqXAngJ/xY3m/4YFSgVsEHUHuFjM0xEI641pB+Qe8Y60e262iv+oUy3cvwYqcHq
5fS2d2XcFm12yHHVgpHp87I36RdqpI0SfL+QgE29cKU3ia8DVyMFInPQuuP2AYow
t56eckCvsXup9PbMHr016YE46Jl09CzpEOcZH+Bg4sY9+pQtG6KZ/sVcEAxtZlNE
HUrr/lRRgidMdq4Xl2E2BrkOMYPSLjfTPoGuVxUecGjioIYSCszjXXYd3NemFOjf
II5uehfkbBVLnnaFph4sclaIP9MCVpVeBsrqy04u7z4HJOOBUA12gibV3pYnLT4r
7P7u/jDJQS5TBmfpPblpDtyZEAW0Xfo8wf3fohe8ikoIG8jAYvJ1ptqRc2/ybqEQ
bA3tea905Vak0UbRFR1rB4GniloW5qfIKAW49JKX5+pgNZ3eSg1XplTsViuxxEcs
ux6U9STh4jcknAu3W91VSbP0PyIob4Es9YTZDmKgTdELpFgNc876ceMHMPXYtFbN
KFkWs9ItSJ/Fxaxx9yYHnlm2MGUbPsd9aPX1TCuDOOSepIUbValAh4SvhEEFiYJl
aiMkWD15KR4m4FOwxzynr3GiT2Ll5Yo1C9UJJgS6jn1cYIynu1QtOvSmLSQSJdBv
cJhOdQojHtaVHdRRn+S7x1SPRllzA1dpIi9GeOdF1KIR1yfcLsA1m6rBKAn+7Oxy
tGUCXv7hIizkIEneDqiycTk/Y/sYV/aceXfMVEsePm8vEgG08cLgqYxBzLGiHZbN
ymFgQ8NwLC4PLd+hzWmSDApNFEK7K2yr4y0o/kkCBItjqUQGvA3NxDmdzTqLZi5G
ZoWPYK0RCyUjKnMTdnbHuexcboOVaoabp9IR7yP/+JI42+F9xvEpXhd+V6O/r8KO
570nQgX53yQ6QIXGD7FTzJnpdPOADm289J0GckYip29P1zEGPNSlhqV+Z7BtmlTE
sA8hiuLo42su35gWK1BsOLejZ2SsgmYEHDTG9PzTPLrYKCwXLSbp7IuGqIH0PKVP
eY4tPSougTjTi6Qk24BZQ1j4Xdi4qC0bLHzdMp4k5IqTNd4dDfnr3eJpqDJHDVzW
8yb2gNwJN1feOHqB4ySI/sDya9pyY3Tkl/vbYp8tbhtN+6OhBpHbJJ0Jkn7NyKZg
wItDSC3CO74xpFPth/wJz2H1fgKdNKt5a2/N+MFKwIr/pQCFghPEv9uAFilsMWHw
G96AKMiipNlUhv5TS65xJMLoqDNL51ldmAKUgnvgAmHkyptOwTTv8RAsYQnnnUpT
Hmhv0AiZUVTVgpwmv5cW0j/dcU8jbc2bnP4d6KPQYCoUzXFrk3HlvATI1OPXhEsK
TrAdpL7eNwiNwty6VhJ22P3PGzeAr69iCQTH/gEIeYExsa6+mXPwyVZWFS1g66ZW
MqVyzM4ps51C8EM7b5DootRn4mQN5hohn2V13khQQ0FIbv8zRQUMzD0HUJcD4ks6
PQgac7HGwMqgCcVmVtdLOk6DJ/lUIAhK2Ht7I5OKdhqS7+G2vfClzhf2Qw1BQOMv
6Y7qP8yQl1HXeiOzlwVfgVph6xggLEMsuT1xI1II1zm8aNJwekiXrS7ZkQc9/rvQ
HsKL3jCERomNue5Obj+nzOBzgZhKvRZftDVDsR5VqOQbMPiaT+XOFbNypjimu3sv
VsT/RT5UgXRi5+CeCcoucLi5SwRSZiIN7PNqxFmkjdLie9eICawa8ihcuIgbO8Cx
vcYq7iDQJMLiWYa5DIgoIG8lbOydFWj42UIyXL+G++2xQuXyZOIGiYBziY5il5ky
8sVaEDIHUhiTFP5kkIOjOoZTnr/8wT6iNAtuj/q9pN7SOTJ+44cozsDNqT2PnZa3
ga8KaBh7I9EfEsGgkTr4EaLL46kHertU1f2qJz6hMERwF9htBeDtri5XAks/3ff6
8ypj9x/HsH8rzPA8vUH09x9M0giQjqGKGQc7aEL+EQgfVtsRPqn0BGSpdZYwaQR1
RUytQ6YV97yz9uEBwP7zzsVjGPJNPeUNubnFcBDR3hRolRnsOKi7CXqbfJd6GK0Z
hRQ1z3nci7yoZM4xT9JhphUcWUx8kXvnTmMmwZecThGOZEwfeYXPS+hEG9fG1KOR
rQC5wzp4a0odFOHnbZnA7BZ0rxdLiZ396ujecF6ACwwC730hiDb9R6SusCDUO9B6
1GQNQFubF3misBctfQRb513AsGDw2iVQpH856JLSpNJKWtB1BtpdIvHL8A4fRypy
hSiL1kXcags6LEAEBClHSRVeN5LcpUJxPCkSyr1ezYMT6olNWYX8Ax6q6jMKcJyt
JyEZhwK9WsdxAnjd7ygncEk/9LRl+b4KMMd9soGU+kRNqCqSqZq1YMiykfDM4Pgh
Guve4OIbDobwACI3uaKI1e3cAdPbG51y/PvFF4Vy/XDfJnFf+hc6gdshpSf+Fhco
UG1AqUiZDMTtTGo+PXQcNqpLl48tU9mFR73d1kP/xYDppqTrszto6h6P27XLa5lY
DZ0OuHFh6wZpK8FdjDNoKvLqXJ+RQ8LzVjnfrvW4f08pSJ+y0rIIRnuGSXuwz9hp
Avh+kWUmZezYmc8eX99KfBUFEkrGbLG257qjDPjUvqw2XR8uT+g5J7sQBRIDlekc
DrInxdQnAojPCsACRo3Qwn4PAyJnNJqWw13ThReSXYvbAJzJAz6ec5BX9Tz+orkq
b2o5JOXXP2t4e0QUs5KT8NVF8bAj0EuPqHm3nBOUX9Ngl/EjikhyRczZ5o4lqPCY
OSdOdZ3KYjeCieH1HMzaOI3Lg19JC09zluLMf+92fNZPpRvrMwZs6YsG/uJumlvC
ZxlcQm5rYPKuCqZMnBD4TjAVXX364qnu4U3lnCwpBkYdsY44vHrKwvz2Tk4qJrbd
+mGJy1aKdA5JSnnv/mSknW9KU9dSnzXZjn5oJ2sEAlBdT8emXrtyGpdbLaLJvT/s
skQOo1yl1mxFSPLJh9MzybkGzgWmRSsDhi7Hs/lY0fNk9LsxRs9tJncCou2f+0yJ
CYtZgjpD/CH86X3ZQCaZXFw6+Y5OVXfPYy3T6dD/Z6+9wjzzTXHhK4D7kh6GOH/m
HFskIkCuOHuVXzE1+wYRccmfGM6wdxn08C48cHeU1ec1mhMFzjXvD8Ds/P1mflua
TvXsqy96tYnPUpjplWLEmSADXYfiX2EkWbk/XAbX+O8k2h8Q3f/AIfb/Kc+ELR/v
ZAhW0ymDkBayCXoXSvWi/FLEbJM8+grpYZSgs4ZQI4JMBsuwCF8rEsPstMBPICXa
fJGltTyMPUkAGCmMym68Bikjc41I4//EfPZcS7tDRx5ed4vyFSGcEeX0NxpPkNwY
tvynKT19lG7BFx3wRQ1IZn5odz5sjUk351lnsR3IFa7a85qfxlY9M9++ESFSic1v
LCHAB4y+T8a58RiujTGiZ5dY3WHx+cXUzG/4/LE+19itc0T5X3EptJ1VJMED9dlS
gq9jeudwRVWCyv3nwVe+YP4hMxtepZ7GIbqQyrQTP1iPMr5wfTVkJa1a1U6j+XbN
wPEBnelmKwa7e4/ovkBRdu110qcuww3sXTHQxLKmYqThiZggHyZ0MgxlSiztDClj
qTBBudM9H8J1ORaSu4KzKriRM0vc/bfQFmay6Ppg1eCDXkyWpXgIq38FvjYEjG92
u5BVvNTGpO8ILuhHv9II3CZUjab8y1iwVdltOiF24yj4gmuRMvW0KJkGsdrlUvCg
mG3OH5eN1KOWvFY1vb3HOSHouP8QT3f0rFW+yrSu32y8WwirntXsKGObC1OaOHpk
Aob7I0jpQSFmdgjNe+ZpJbo8BZREeWxhJOthiMSESS+jMNiffjxj+XoiZsEK2CLW
0zwSt8lpfU7V/iGWukdRjIzADKKh9PN7drr6wOb+GkRc2ucPFfVQn1FVj1DrkB2q
Njjzs36UTaC3D/eD43ycG+WxN6puprqb9WbqWDYrh9PvdwVZPmI70UmzWPPscSxT
F3p0SUKzntnoeJYd4WFe/PBq2IGnince7qxQaU4/6zJxqjOXRy3YMjl2AGMmH8IH
cQ4vsZn5dXMeRzJaIlTGiTxTwagVGL0AlAEqf2SES6wyc8Lz61OdMfL9gCF/2TrF
dzUW7lWSfVLDUCPTlGyY8OD5jfZicYxF8Qw0AalAZ+EGETadbbhXiwjG+hBOgkbR
AkDKF3ZSmJGQ4O1ClZHe51lb/jqZOtwx+Ib63Li35X/EzlUZItOHg+Ty264Xmu+E
sjM2EtwJRlsbxYXpQwJz+IPrHip5WlFVlFj5t/kD5ONjiAdgkiHET0yk+jldgvOx
MKo8JH8JVLxlpCvlVr/fic8q8KtE80WW8RwBHdxbprAwF4XMcuvlFIGPrOj1sSEf
czq3kY/idLtWyQC8PTofyJtYS6G/dhZwVVGXxwBhPzLLOqyaGoFvZSiOIAycmqFu
yrbZWEEtBGIfDrVtJyyb+T+Fhxp1KxjWKJZX/I621jSOgO/ZiLlofL+svlJMKeGM
u1XbVWirdU/jreQbBu40NjtuUaDYPVANXQkLG67ZbGS10pFNsLGaJZMVn6im3/L8
7DGmvigwPMldW/kkLy3COOVHpStKvczUhPOVDVzldNB3Ghr6ddgrOpHl+pb827jl
Ly0Wm+xZEonK5SU5y/FkduSGeMFFLG/pHbOrV/aQqe+9cx7oNp8IOrmUNP+okf+P
bQbu9o5wNEWkyP/h0XaDinJqsh3tjxMpO6z5L66EhwNAiFuu0pDhRbbFSyqwrSvL
vxPGbTnoDoIoAyRg7AESroKk0EAHAJakVNqZu4F0SD0V4rCH3xryo5K99IBPdx3W
ADC/+lfF/DSVJxxH9Hj4DnYdYbhhrww3fslP4eeEfL+e/xVGRg7qkSoFnap3SjW6
LWAHUlo32A+BFCmIL/g8blTi+X3hnbcUVBq1dNE3SdnVxJyqf2QQ2x3qV8TfK+lH
fAUnzBx1m+g+qER4x8xHwVVI4VIbggwSBPsFD/MKL0cqSooQyUOIHpefAOJJFGVN
y6fLfWj+vGb49ckpHxcVe4X7yC2x8doqoWNijr3bvT5pWVI62P4hns3iClyUSp+C
9Uf4AYcwZvmjJeJfSa8oGvZOpVzfzZkDVwMr/HntDCnakBRdpUHK2k8MkoLDLGoS
mV+rWKlQuUXKJzlhEsUnJubI7aTXXiKujFAEgvzHsUlZ+mIXfN8qVJsHHtIJ+7wP
JYbIVsqVO8FYIuE03avZlGAXRRSk5l/d/Djo3u4NdlwscSnJ824udxk2lgUkv2nr
OmOa9gH46/fWsELGG/3A+W6pNIp0q2DSmLrWzCWPB/CvSEqWqSa91UQ6ioEZI8ea
YaC3ExIBiiFmJnv8jertexOHjASKXtMKE9gB2Whkj7wcHzicOkfNGWida0yuivOi
ltLPloDKGRswZIPar8/bQJ247+QfwUxIJ5OExb+6AoweRha+OL0Xg2zMM5PIecRY
lMpeh6fmIWoMBYAsN623rQSu/3clIB3214/Ndwo6hVgSWUoNvkNUPq8pqGwz4ZNI
9SAn946owXz86vWpmP7LDLCtXEq5X5SsUETVDo3eVLss2/4pIVP1bD3hN66qYsnx
SYEq5zb8cmddx/id5nzcWLdUu4DY+e3msp8vYEnHTdwtPLnsmVWAAEqNjtWlSWgp
mm+P12c+DAQKC+MfmOaJP0uX7qWQhJmH/5iMwnV8TL6/kEimzMxyT7zDTxzr8Boi
MiZPnDw/a4x7sP89h6ajwjtuUMj1DnB3HXD8q3CwhtAu62QkiaZVr/UybQJgEKNs
Ze6NVENOe2GGxJGTKEPRDq//c8qVeyDtgJdjGruL2lzXy5bF9laEP+ehvf1f26iC
UDQP4udcPBr55A8MaPrvUSs7iA3QATGe3LhZMEiZprg++SfZixIDI+IKmnHCABHk
xQd0L1h2Y7whnwAEXF4pmKZJ/5iiAbx53+osd/YP1vroHMIDr8xKtrdOx5llZxba
NB47xPY2dYSSyTXnZ9XdKfGsWyQjcdFtm1Esvxkd1jEc447m1F3Ln69lKSu43zrQ
v1GREi5RTrO0YsDcbxx27hX6N6SS2z1motS41tL3sbIAD9n1Yoc8cnnW0g2mvGrO
NjI8wlgYj59GgMbMG1UwFsOVhgh1k3FneacyDdClu4e5U+598N7wsVT5sX7bj9Nk
YOghBK7JfyjgorGLiSqy5xHn1ieACl6r06TEpBi5shoZF1e88j+Ilx/zgeUVcVNE
lZpTqJQsSSNpNi0OCgDopCJrzpxukP285eJ8veLkONH6WSRQJ4kspJvKpSb5wItr
RGh7rUXs6+1olsOY+mB8AheXkTom3Q4jU6PFkHLh01FyCNTTJcv3b8MJWJN/9rP5
mjGVN2nnyHGL8CyH7ojHUgCdrBVfIha8Ewwxga0spIglF9dyucK7buhv9sZik/z8
kN2OU3FMGrb1CBG64gA5VIOBFFK3LZurX+F5cfaR3CUt+UDLFcbHaFfrpzR4BNaL
Z1o4obMA/I79jaqDDcH/B+ICMNqKCwwnup9ljB4S7cOLJ1/HbAk1lMY+IWkQMb3N
JQgZzlPNX31jntWKVajBb7PmnCNSk5aX9XHKc5iT7QVUztmtqYaqFEKlZIqyBIpt
I+ASMxsd2TGvgIfQtS3ot9UubWbKUX3XuWHrQBCmrUuAyfGdd1K0CfbUVBihZtFT
wLJFoFB5Sckc8dy7LkAqIcZcgoA3AAWYvhQRHvV8uJvgI2+7DC0GHk9WX6yv52rF
EI0xd1FHlbNmMP8gX2iNf7TAl71gDtmviehQK6hEzCARHI7TRATC01ydtryjyxzO
6uv1LkJgzJ6MiLA8KjUKVL7nDJ790cJg5drq0xwVcBdJbt4x8/WUMovKzVfTSOM4
/NKNefmC3Kb0G3FQnmOj6NVb7AACao9PzYSRVzNPnMbUWz+125iTkr4LYaxPGy81
DpM4ZwsaoapLa1F32y09Gtx8OGW/NBHxTWMn6DyY269yfN7adkNXARqM7YzLBLNj
LXOaDqs8IIy6I1GxsFcJJPAblfcS1ANJff45coIZ3Ai/+g3ZJ3Egbx3Txsl3WU+q
w8PRfZOizruJrCKfTeZdXKqkvXZn0id8clpogVsy9E7wZlvp3v0gDh5nkiyQPu0M
qwEFaMOT5WgQJtewit5pBrPwjsnauXEHP+64gZJlYZ6zm9MWe7QRqBF3Yo9HwoXI
znWKmcqjqWqQiK9YuUL0swsnsvEvfcN0jva1HFzWDnaYVkzOM1BbZkcN1Gad80fk
Vuw7kZ1cFbB0MnVs7UR/a0RTAUJLvs2Nl/Z6khak7f+mZqC/+YWiLDTuVMHygeMF
ChBx7y7k3duUp3YjMVdIUeIC9s5wm02wL0gTgui/iPLJ7iXyzwIFWaTNWj9G3UwV
7E3VpDSw4GTtknwywBpsLCn5Ytf9uigQkEjlc6MyvhRWui7RgJRqb4Krb9oMirzB
wipclYbbYCX7GsEAeZ99ILpCwSU58p2Og3cBpkR3LiniSP9oftUqgaDzSBgBUM3p
0q1qhidOQpnjoUttGA0OzgQhDqffvN1OkQ5gipxp9oaImPgWADUtZ+bRZ41d43MF
MQZClUF4YIfGmRG1kvPO+7DuNo3ecV2UQDfYx7DxxoIuAfzOy+7361GbtMz8KJft
BHoSm8pPBmiu0YMdUCstQkD5bHl0Lv0sUZDsDFUTQ/3JTP5QxVIUKmuhPP1RYg8A
7DP9fsRMdsp8ybZ72sQQvM2ieDDjVbNYKQJ8Qh7ZZF7iIs7wHqtY90w11ZxePOpC
slEk1w5TLVyfqP811HaP5RsWWcwdBnDxVy6SsVvKoQaj0sS5s2IvvIWkcF9FgXIA
3XDpB/z/jkE3nJ/gmPk5VvWzKeYfj0m6+Jg5v3dVS677NnlMZ4jhDAsQdn2r8Vjp
LL9B9rY8BdcWk4hZNSLoQGlirGrZniqjgiWQRyta+/mJ0DKDlk+1WylD7uYiFqrf
VML1kGhME5iFSrrSXl05AxBT8/k/MUi6LT01jFk1cc7HNdeK2kwoF1BNngEDvSnR
e7YFrho0HV0+yUqMmcY/96ZfDfBqai2G3TDvudX0AAMbMjIFS7lG6kVGJ+AD4Azm
mER8X41xBln6AkFrFhYNegioZTnp/Ni01/C2gNjnTf8+WlB/zCwkQtS2Q0K/eFFK
1cw8Guc/7xw6SwRcKvmN70tQy5KLq0///BgYEPZ5MHs1AjuGFsbwU6IwsHzhB4Xo
jdTSSSOwl+sjqNAhJcExAZG4H38GkFwi5fB+61HRSymK+IkPquyg9FD7vBecG+lm
lEBvbZDYu7BW5AFJbmRpn2tOcGwCKugo59JSUU58Leb+L4zqn3xK3JCc1vw9snhL
6oGE6NOcxtF9KqbdOwPf0repTRCAwpcNhBrzlpY1+6W/HBKhEmT2uiY3GZ/cMhF3
7sttRPx+XLPPVZK79yVincePXETRE8PN8Tb0jchLprYF4BUXRs0DqVWlJTc7x3F1
0hyVBadDCfkXBPQYTYtwZHIj8QWGYHTxp5xz5xDiw0vgQBSadwwWnNKnTwR2l3pM
FnYDHbdO7r+PMlWGetNj1fwGf+jBFuQI0YpPia0MY9pLmHD/0GI9kJKTpEab1CS2
7dj0q3x9hMrRdrKciNdbLUqdl0/HII1+oseqemVcUadIExR0giia9kmdSRbb8qRr
PoJZvicIVxvGql7bksVm02MuHS7qfPTKNz91W14QIUCg8Df5GWS2Y5LNNiQKln39
BpRS5CM6vYMwGCqrThUiNbJI3XV5SCV83HeWhng0FXI0BAgtDGSpTo2ZmbDr+0n9
No8leqy6usTMIkR9VBwsYs+KjrKSRO8vE2h70+zQmF9O5PW2z5dcRb9gcAkBUDJv
vHb07tuLWZnud2C8Dlslyc80T/ppJTYXDD/z3lOdeEAyDGxUEHmzei++KCeI3rkf
Mr0Jd8cirTnVikS5rZa/KSiSEI93sv/P5o5EFyHrahVJvvpLRY211yW6Ob4Rn5Ky
FYd3sh52lTDuWUixtZCw83nvKfz9+0jmfN2jThzP1hAHgkVO1TwSnao0nCu0k7vX
D0DCVXA6KsB1u2iSWZF/+C2AdTHwj5aN70b5HsCRQYLKCjfDmfAMDv2jll5NhdHk
uNawun+qOA9uce6x9RSlRhGwsGXi68oCO8b+OwuQUFGn8NmoR3VRV+kyP159naif
/4tUo1kvNY2oyzvfkEjomXwdrFHmOCuc0IVUP2hkqRByn2cICoMl1odMxyJ1NOO8
/+L81jG1XbBj3UQSUKMBubV3o/eIZhfuVpCN/PKAKyt04sxmRXMgUmCWPqfjhzrN
T/6pROYoG044PqM21lWsNPy3aIjA8RMa+9Bh3CtqfMkLkDD1JedyvS4dk9YsuAuJ
UIiBevi4b0ebOcmTaTpzfVBFDwz469qa4YAxDhukHU7K1CjknYqNeX7U2SudWAqI
zuRK/y6H3C5Fce7EguJOc7wq7ZhXJgcWUR+htTsZkMoVKLqI5eaYgzpc9QkHsW4z
T0CLV2l54XgNPq2dc2XvCpcqgCNKB8o6viLt2fg6RZl38mtpbXQd4kS8B+dtgb2W
ESVi9ccZvHE+yRWMePCPiPtXJ4v65aKRFe748cju5QPF3inn05ISAkc9BpIb5Qvt
zAG98QrddDOmbY3BD2vbEWVJgr4h/Yilw25mpJW9lvH9U2qYwf7ZAI6LH+MCntg5
YErHcsC7fSVeMDO6N4aIXwQ5qCH3DSymkiYstMjcVWNz+B6x148nozbtyt54ugVH
iBpuYP6GOqGgG6U1dlC8tmr3vfzWoXK/tSqGWR25N9NDTn3e0dbIZ7ew2LjlkG55
7pt9q2vJ4Nwk/08pxK4xXZxXvvpeWwS4+scF74C4/ELWARCuSVhIlV92t6LYs8y8
ikvSJ+UGQ6bBiLXFeRkj8BfqsDC0e+nJ5mhmA4aUoMni2xPHObsk443p3bi8OcMw
Ar/Ls0T7OtGAH4BKlnWfpSlfdKIJHo7WbW2yaSOLmeiSauWN0Vo4o2wey2g3txY8
MAvdVBZlqOUth7qRrwQYHhlZRzl9SkNDtTIQ4ZwVo6hWhPZvRYj7LcanBkpjS0L2
4+qP1yfmkgwGQTCsKkehsxgOCxe56vgONYlUgF34tV0647D8N9+FV/ZJkvNTk3xP
BmQDpePsEMAuWIK/IJtq6+gclukbpeGrP5gPToP8kZNJ8LACCpjFeTLTvrvbg43G
rmyyt1GtfYCmPe3F588ZIlULHxOzKOQ0wpK8P1hdGvmoMgq5Rl2HYTAdarw8aM1w
RwwCUU29BzcwG/1EJckL57wFWAmHF+77x1DUSsY146PS3S9UAcmKEbRYjRLo7adb
IY1zRZ/rQjWADyOoCcu/q+/fyrGzucnlfZDvU1yOjAKMVr+CjPGH0rco3n+RhfPB
gHBWYnefJW6CuIIaj4DKSbE9D1QrT+UbCoHW6zogKQqWuZY71C9ifdPfpOMB9EAT
Oif/LhNrcvwOF8ETlrNGUkgvRTE0x2iDBxsNe1mfjJkv1SMxQXEYqfu/qgcoxj6V
+eYpH/XUVmfJ5u6d+eIGfcQ8MdKvsqxEh14CYF1trnKcs3pQJT/HOM6ilQ4lmVPz
fto+5NUjddG1vr5eM5IztxiEZh7eul/FEr7Ez43pA3KlvVdHMIo2eim3HZ+72K7Z
ceQHlTrHUux/7Fg8IX0ucITF9nw67EnFBNgNKY9v6RzIN5h/i6g4vZXTST3QAJRC
9ioY9KY4V/01bhQjTjzPe6h8DSF/OLnzK0aAJoHZxRMchKNqT4SgEVoSO54ViuEe
eWath8LT4mG7d8G0sqQOuB3y2CNNx7wptUIQ2UoI4mXHrcOtDCR3eJagPWN2VBZD
5szc7WXvni+RCfbdvgop0qr7DF16S9lQrUq47Y7NdqhkJQaPYdXZAuYBt9SDbbEG
IEK3iDHGPOBeN/nRxi/slaXymHpWV38J43fpGwb4F54KiSrOml1wPtJMS4lFbXTT
X8m7v8oNm0BUToGmxOxFE2ErB9ktOvcgtjc5varoRWyKaGd4r9GiRks8Kxv5W6jg
k1qRLoUHAZK1VAb3/PWJUUAVM+cdJQXgZZkoC+mMjmrMthTqhpQBHZX7n7oeKbM1
9/YypueC9ZTgEugPjuAGJHquSIKVgPbZF+b/4SCAF5FmH5Qap1KAedoQSXhvqtJm
IIgXBpxc5k+qZq76c6zOrU2ER1sCYbL6R662vPnIRDlgSVkU2iSqo4XW4C/ygRNy
51Qa1Hy7x6ukTSpKxT1y8aSVI4QVBIhmemRnd5SPgoVtufyPxZNhM6UpR3zMe2mA
frf1wo934uz3FELf9XHP8+nQ5YYOvQnPqwVWeqKkB+vKLN9mxGHjOWKSOWWQo3VM
MR4SdlSWbWbYXeWm1pjrHHpm9jGSwSEWnV8y2AXcGMwp+aT4vqbsHBPyNDobJLfn
PiQlRYcpHgUi+JLt8t81EgmvDQQ0wijAV5uZhVaDAMC4OI/gPVKaFGaOuxCz43Hm
fSXMd+XlsFJswIJ1GcOue8H7MsnLbCOOIgFJAaR28/B1EywpyMYV2M4BH+H9kSzY
XYA784cZ8nb0Jr2Ky9bPUz44dMzE9xgyrPlFl1rm306OTJRgHniIo+R4ZVNBINg9
1eXQsOJzXtug39s9DJjdac2mM9z5+1ci1yKvL1BaEETIQPQLZqXZsmBsiuNuGrDS
fcIkQa9Z9ZaP9vu+VX5+Eo9BDjf89mYkQkVO6AZEWlvrKBo4e8CnOUXy0U2RhVty
mxFNH9hLRp66wMxsnfLq05oxQz/z7ycjGzc+Q/7Q7Q8MtUrbOPo9FuvTKHUOJOMs
/0KXBHKIBsM5S2MTFcUdwXS6xhfnRIIoncbpIbt+tc1936uVA3n2yufJwQ4LLeOL
LJT0xRw9wc6RvK+I0QvJtueU83wq0kTa2hNVQYiIX3RDedhuAbEeSCHbv+0yc77F
y816ahLhk7NDXbyqPqgaUUdgYB2VvZQG4rOjQJ5qisv/pnEDxoWxi3c296vVvKtk
zYPjGcUkmxQFgwXK3Sm1AgFFTq3VBdpzyNqeK4tNlJHUQ6LAm2sSJ2KlH/5g84pC
3LhY1QOp5Ywhlw0Z9VRC2tK9uhU28gT1sL/sWRQkhg6ff5pnsQpi1Gd93dcGIT88
fqKV8G8/jAb2PIquiBn5dc5gJbtSrKFkSxgHASPc2aR/d3UJrlmzMgyv2RXyBYEO
nWYJT50VH9W/2zvs98sDDFXyA4FXSKa8Iy4Z4wa9WCccdL0GSbqvcgLNHA3sSYHq
rHHQmpGZX3LHZ68I0UvQpgRYnCqXmnx8Yoes41D18hgSLzG9Aq+T5S2rMdTS9UJA
88j9utWvDiTDs8HiOJzgpOo2iwqmflRd9rkvZa4+5PX9oGZspYdXkNY7Ay+U/0wo
tNo5rhfacXD53SrVE3NYDwrGJ3fFcdrNIoudrVXJP5IAc5vBlN17w8jVxkSazhDV
a0oPzGo8cduAlNeX/WKvORPuW2+2P6ieNshViy3Z0DNC0qu5nKHj/7xdoCrY4MwI
PkRJbbxRPdtiWN08qJCs8ng28bUc+qy73yqf0lg1O5abrKfHWWaBTqKHrG8nET0r
MSAYl7qP4DYeLeBo7N51csyrvOG4bu7a2mBLodBIs4PN8CZBWi5TIZCL9SuYrm9R
rEA5W54GwxF+wJkKGFhuRtKPiWFjDAAuMEwvAxeS7z6H/Kaud9oCpWs1ajEpAdb6
RZG9UAeg85MTNpcM9+cGdStsH5DvitcHE5EcQiDgPQqTzjHyySSY20c9ETodt+C9
3KmCb9XMC7KcxEGNBdLG6WVmoyDxTd0eT/MS4YMacEwPpaxwEEeYI785hJRgu1yW
fHc/5IEIuOnM+UfrsCbs2NxoYAWXKu736HXg9grkCC6b+J5zpP/3mQ+3MtfMsDj+
19Kbe1ppDmjDUVjrTk7YwQuJVZ3xJbTv++PslZDqoOIgElhFVXtfp0PoBIUWrSMl
xzMFrTPzgcIIEpJLuzqWIlqDzoifEZvSLkjZyxyXC1Fz0wuPgFZ6jGPmInpauYbu
fpdQe8yEPW9m8WM9dNPH4OzWUfMhtCXcOzVUiup/Ccm40VheeGUeVgt9lfqfYTIX
fr7OORvVYEQRqlMvkYVqxObQyUrLD9IfuwTy4kqnfGQQkmkwwXcY4crN66KhJJes
zLUdDair8m0sijehddENy6JT9RA/tLltxYAzKQOwdwIMF7eRtxqW8sqRRY3HRCLY
FHZQ6TYjl3O+uwax3LFG0MGYOA/sjRYz2Z4mQ/m+f1cjmiPW/cy6Xv+ljY/gY7b9
f/s7Gzg+T+Le9VtHdpjZcEavUPbOxrbv6mPxPnmPHsT6wqtaXaw4dz8tlrh4tZF1
jO3KjqBP1FtpOgCPU/y1mEOTiJ3mNI3nYBIfMq9eCmka5BLhcSEsfgbUVMZDRVpZ
sVAWPzFcjntopmbtg7oGcoq3Oj0jBDaznF/lstjOkyr9S24p+4hr+ZCRC0exJe33
NrKQzRiwNrMleugRF7kzAVdUBznrIFKyLUuBVcCgRjxhwG89Cz0tujZ9hAFj+8og
LO+ho2bNEh3uiTAJowJ8X7VG9zauzDWgO1KhuWhtz4Bpt2b69zVRdQiwnRaIok4D
LTf53U8WghpLv8E0//nERGOFtRHzBLVGBjX5Dip37GvL3UzL3YIm9gOHcfNFWdwl
dxIzYehgHa0k4JZDl7XiwZaQ3dhjH7fpfw02jkGs4XMPEEepbvnRYcSF3cNIbCkk
0SDcPgi591phhvOrLfVPwA+yWNxdDubxFwE6E8Tju4m1XwO9CSl6RRUDsdVwWUlj
G0UwHyy+ReBzrnV2Gvw2JQ+eUZtyCEM6DlWdIDOK7Jga6hVkb0bRFiNoT7nr+rNF
tfHHcDzDyYxT+tcE6LW8s4aQ0Rd+fPnpoH2F1EZCThJdTpZ/70Fe5SZ4uvK9Uu5V
jhpKni6yrk6Vxv3TBNr0fkrj2duvUTSIC7itHaeUHmtW7MuJ7WpNVRPwv4X0n6ph
woVGqGx63WCfF7YEBdUXvqrL+WzwBHLx9LKAIaz3GhUvblHKA8gGB8YXNsYwqpmS
A/qkshcxROAcnbbGr4EEoFgYzThONSQYWkbaE3IJ7kHLy0HQF93PnDrV+3UKxoUG
7poctwbUvdIhx7lK24plivYxYoyNh1G+TtXgICUTcLnWzY6B0xFoEVeXj+f4t4uv
6HJ3pxkdevHlWCae8gDyOqPrQ4sb66Aw0JoNByG+IptGi5cMfa7Nd9PJSEQ5dZ2d
po2GKYisDE4qWovSEQg4quwQstvxujFiXupVx4e4OKMtMAP9PTcjCAc8H7TvFwPE
La9iKYMs67yQmuiwvEnQu2KRrwAvkTNhLtiFc3PY6dd2rz44P+KsPVxY+O6OE9dP
iiydNIp6pp89J1MusHan5u5QYIXzaUJ+jVmwhyQfQm+cE942Lb0DqHqQYdBj/naA
yIWgWPFWJyZlCZNqiz4cZesRFIwCYZ9IOtsxo36C/l8T+qCU3CkPq4v8z7RBiL2I
euwqfb6gYFmGZLBblEhGyg+ntG6xG18cTa8vEDcxb1GEO9FpnhhNfPOpSgXPW92H
a17LZJbyZGOOK2UoiTtEOgS5f1Pbh5oWWhfxxCI2yBNuOdALtE5wIfUdLmgGEybz
ZumF2mjX7UkddRs/4AwxekMAboyWRCYpeOWDZVi77+zUmfgB2narwoEQdGg5G1ag
usKAjLbs2j/95mKoJOLBH9+v+g/Z4xwwEa6wYfw/etoP3lRbGfoO7FOb+3rkqiGT
a/oYgmMtakWx4jo++VV51srF/UPuLDLXsVsa5nhffzCPMYFMVqZMsOAb/TrhPnvn
+wfMpiNqpiRRh7OedXba5gCAMmY88W+9cBz6ZqdgxFvLNhmgQ8qO8AwzzgyPxWsZ
1iWHwsGHWvuNVTIcATepgrnTqg6cVufu8cN5B3Yr0OW9EzmFehFnWjXS6tI/PC6U
9fpgr4s9dC2FWNL25CJ1rIRF6VzXnOyrtplYRdz/aIasHwO2WQXCLRbc5yUN0Kw5
SMsw5MuFG2TZcX/PfCPItpFEeZORqld1xGxLbIW/Z+FPaqTfUuMOd+Dmln4lutQQ
r05tc0oRxTNW//RA75bBnJYYTO2scRf2SuZgn7O3nCkUrLx4Gc5N95dtozG+b9ju
rhNy92FFa7rssrspBCH8RR8Rs8/8KFmqEA7Vr8zo1LSDyF12Xx1Yw+kGnf0d0nBN
1oxjfO+04yBu64hrU5DoHPpdGISDbBeKfpvPwBZLcQB2oseb41TelamrnpCDiwLN
oA10EV6hmbrM+qMdQSAZdf/gLPiZNuH4ROKOrB2GoArzcQ3N04z1KW8nSXTrCVso
6JwBzI2upkVSxfiHcf0rPymotW22OYb0U4MPuyNpOfbSIVvzbG4RVq5S7LhE1mwI
5gsw8QVPDSUSo/7AT42QlhOJcXpIwW6qncen3W+0d9EAPRvtwwoRekGzK2fMk7NT
LMkYLlcJGz6yZA6+zH3qClzGMO+uu83u9VmNGFNE1FiTY42QeIGSNjT/xa6qF3oh
f/D0WfDeEZ3U9pkK1YUhmmn/8/FltdQtSVppvoyCkTjb3JXHmgD9oRLowswCVRKd
9o0qy4B/GuPY/AjJPbkSvOsGLyXIKs24mGw7xCGdta/OEzgs3wzTEXLBKxXz7lxU
pjEcm0dZ8+0pbeYd5Vx8QMZFgQLWJAu1zytTq6o+Kp+GRsXYJEaclOnwthePnk/I
LoZdoFs0JxEfMm4Y6CIrCjFf8r2DcybgO81DTpIKdxPZvxV24eZk1TE+bAhDL/px
xnrFg6dKs6XG6ZDWgWnfClWGm9e2N84b9vUHePCOc3/vtY2ZVhP2Fips9kEN9j5b
/WfRyOh2PdSjkX6uuA3j/w2vlhJ5sVHtW4SW/ip070M0hvu0u0/MLenwNciQJUfw
G2z/ItuNfDN3wh8uzz8ikPXshERMdkEke8hd3oxgRVWviqKyEXe21fNhM5hDYBZj
+47/aSGEVMiYs5T+cEaWhlCrc80y18mDUoUG/fdBclVU+aJ72jFyPI0qsawU4BSE
P/PqTtCVa/OEltUS5nsJ0daNYnbgiqWiI6iHVn4Y6fKibTv0YwGcmdmybW/uGCFJ
pavejH8bbcWjYRStyGh0p9j10f7+gOSuGSFdKM9ptifcP5kzxQV9eT0IFXd6CYrb
idHhlqj519IhSXRoUwSjyeR0i5QCxZXVQ/utpvvq1XWWQigma6AuvJHA+ht8NMNk
34Rwh2FhFtWSGU2dXiuCUbzVyv0bndA9z4wzmcMPAHwIfo1MBuF/bV4d4xeFhvZ3
dMiHby8QcqXF0D8IVTp2o1EpKmAmIRkitBR9viPJNvnkxlg6yqrmTZ8d+NBnhz8R
GuYO331e/TBscdbGyon5xYkW3123CATLxG76TgdkY8zFERSUtk/N6tKE0d1o9euX
RJVXuXSC/udXg8EjdKNIcKDhhyZ7UXnodE/c2DcKdFB35TMUf4FzFj+Y2GN2yTpz
04LJTSW7RI9vX7F8Ut02LXPvHXbz1ek0+v7YOV6NhLSIf9IT1dG8QWvNS9omej9C
eEMGOm7MFPkwi7bbKsVyPE2zv/vp1xCtZaGBy1RUMJzoCjFpE53PxS4Euxh656nX
n1/jWJOdeD/m3w14L7FxkqA5AMj2Gu7iedNyT/U3J2SIHw+RUPwl4lU/RBFvahLB
YI3+27ejsotdFIWxDgm4LLrwY5ayGc6DLIg37w5UrpzeRLVe3puAk/A4fu57o1v3
GPjxIvwJaGnXIhKnoQIjAaQsFX9+SFfjZ+tuHnlpAQk3ID3o015ZkiAta33XTsr+
jPcT91d/mtOdrSiXdzfVFowdENVl05kAaSaAoOUuNkqyYZ0ttDL1+YcQfzifK0Uk
6YWsxaA6Uxq/QCnks3ccf/uqwUlruqykIiEG0I9op5NdxSFzoZjIgmEgZ5oB9GVt
DK8b/ivfIWg6yyuMt2BIc3t3bSW0+D3tyeggqVuSdmB1TKzP53gp/WX7dQtuHhDt
1PnBAPrraREaAgaWHJySlH03IRzyiErItGnMnNjXoIA=
`protect END_PROTECTED
