`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CENah249tv9hoo88UmU4z1WFAqF6wzurg1ThIrJBQhGBvhKEpIXYOKoPMQADUtV/
ojDIZOZlom7x8XGe5thm9keg5CjHoNkgQnMefKJOiH3whe8MeoGVTBme1Greg9qv
VqHRalzSYYEtYyVLwiCe/L6zCHpnWjLE3E12fk3xLK3JyQLFFB0BbUDp556QGqWB
m/8vfwm8s/C9udqvZuPVfPEQ2s+WadEKHNp2H7XpPnfAyHCgpmSdw0U1TZNR438M
xDXdZp+EorudMDiJ47mQz4J8A//qDN+abGE0TkiVZY18yulo1YTKOhy0OdvjxnFB
5j1l1tipOPA7IbHF+VCI4gfgeYjZOBqPHX5sevJl5Yw=
`protect END_PROTECTED
