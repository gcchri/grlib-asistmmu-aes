`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yAyHGucrOVDarcZ2YxIPMd/n0vvcr02NA6zKUm+3pxWAsSWA0IxHAk+F8eyfEp64
ZzOTaEoJSh9m326g4aNhzVX66jF0ZOtl/nQqjuZY5+70d9Q9ycdvpLWmuPVQ7XQj
XwlNSv4Yv1FoD8hTl4rlFV6y+26AZL46GKqkphzDDjyc2MO3LOiUgvagGNnq2j7g
Saoq2uAZ+7MSBXFsT2HlUbkgtRlZ5eW06WpeGIyq9b10VHnS5LoSC9fg8p9/cbY5
qLApbgWkUkWql4V4yUMIqpCDc0ilHfFyb7ctGnfgnfGa1duL6MajKpeQzrFcqd7D
OPud5j2elb+CmwZmdmd1xoAgQR7JpiUFa0HLxO9w/oC7fWtO+91q0dOfZLxVhvqy
8N5a8QFiDs3J/qyiy/Mw1pnlcwpc/maMVId2EVmEDFAToJjLRN1hmDtzqzXcpVCF
uVEtz7VDm2wDApFReL6Jvd0VbnXDXNAwBFgD2appVh9Ih9Rs9BH2Ya+sLMhoVjGB
VbQK9SYnp2jzgLoAuUgBQqg/xMkBVR84Emu5+FWEExnOZOLNXLZPgvlQi9SdHQLV
oJutrC7g7LwztoiDDmBz9bkKEKQT8B2O9Al4pk772/7rQRXwvqVg4615UFniV61C
IDazef3MEbpljPYZ9oACU3kwRrm6qdnw0rH8XlDckjDwi8akvuMe1fMJOBjDj+ju
a3dcKeFfctFboaGwG3Oi78Q/5OpcyhN7IOxM/DqQdThPOY8p0xT8PgnA9gOomC+N
15sr/5Incddwh2E2uv8g66VI8PuT325P9fJQw6xDzpofznAK211uKptpndIxR4Ot
uvWFRC5gQV+1LgkROONJBbT98qRZHaqXpfpDhp37BxRcm7sh26uGGM4dFjiJIjXm
ujtNp073D4pdN80NVGSw7CdaOrSgBYI2s2di/kBCJz0=
`protect END_PROTECTED
