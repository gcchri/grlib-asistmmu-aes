`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1K/wRoD25KMoN+Lm1o7djddQXW8aKp6s6vKj4mJBQ/kqBY6iUY5Xg63vSl9k2qld
GLHOkbMdgrGtItjpuRfjWQs9RgerPHE+PftAftmYmBzatoHtzmXY+P98Mszgk+y5
LmoTlf9JBgjnW2fOutMB2tKNg6NhCFHSjr149BTRWMbxlnKVQm1uf5cAp7GbmPI6
nw4Rh3YhocrqARaxm2Tzf9gSfjoL2nOh0Pq7/NPq195POHt2GZapSguwJNh7CHi9
NFPeKCDj3Ky8VnclEPzeuURvZcPj4SV5RdaGpy2oJH+CwAbivkcTwELnx3CfqBqI
812iVYBO6uBZ9I3y1iKrng==
`protect END_PROTECTED
