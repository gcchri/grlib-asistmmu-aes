`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BHykZ1GqbflOs6n1uSzPoLNvvKP3Y/8fi4HRhPJWYa91kuS3AFd0+vl7Mn3P3AcQ
Jbl0KnYZ5alMDhV7pbdtd5tx5DZaJocv65+jHbztWBAb1rwWsLB4nxe+iO/02rHg
geLUvXcFHc3pgtKrRLdjuzJptewt3HZwpoFfuWMdBX/3IBC1m2AGHvbaNmW392Wx
mKiMByKKfIJbfGTW4vjF0/XMJfsOsApJIgSKtIhmvmigjQcIVzr6ENvLCy0bOfQ+
yi5MQMzchn1oSnw/M6kmEoRydlMV4FUCngMvmI0FdZnknPYLG4GXdDZ2dGmuG7Ju
qltLiX2Y7XeqPEVFEB0dm3W9IDK01eiLKWLqR/HNf1MGFFPtFD7pl8PRJfak2F4G
Xd924YHGaqB8AGYNzvssOyAG/eP7iHgIxP802pqy5hvhOtl7+MHmiDUpOArNFJmF
sws0+JguLB1c4f7IzMkeZ7Kqcmzu52uiiUga7L26+kmdxVuftwVxmXm1HPDvpOE1
eMkjc+F5r5oMqwmLCVAzH8ak4shOCgHner9I+v5gxReVwtrfpDSWAYcog3T4dTOK
2d9COP3eE2LFYZ0yiv0RzaE7uIm9kSeNOMhLneHPidiNNiRK/8ihXzNap0/Pjw6h
rfXUCX3mTmkP1zWM8nQWWamYr1a9KKqfi/9ZDRB0zoqB9gV/JqtE/uOoRfWciwwq
vLNzs1BhpoQM0mKn/xKoUVE65rpZZVQ7ZbxTPVTf6RtnS4csnu0y47jE1PA96jZY
0PaQlwKZYLLmTNTql94fKCKk+jOHDsUfWKxzgqFprNLrC/i8/o2vz7PMuJ3IC4y7
3ewZZQBYarUIv7CZC7tdXD9xIwr+wOLwV0SsVGDYfkSJalpsgb76HWlr6i3/NyZD
Ivi2v4ectSYUjj26GWVVPxsVl0aZCcmP8GcsWGMwzB0ivdZpKXgcoP9X2O+BbWwj
wi2KDR4SkavM4x+/d/r8wP/xv1XbEMjr2fY6q6u2bHifa2Wo756q4Vf3PF0CnKPh
0JEzWKvUtn71XciILN9mnfd/zDmBpX2uejeZyCMutkol5LLjSFw1VnPpuGlmWNli
W+KPWtGYwjOq9iLgigF6tmWOyl4QvrlDeSwB0v6sbpqadQgNkCQVZWUY+C70ypui
RBxSfWYH4GtsDhw9RBd1kgpGAqorEhqCGk+PUk8iXLA1Ccq9hWf2KM20pq/MioRu
AqsKTzWQ378QMfptLKsYQFDGOdDAlyWVMw0RxK74GWPunk4s4szhT1KpBK+c5szt
naFxegsvQ6NnVYPUiI4BAkXsRphcRJmd3kyVpRNdZQJEBS9UpvdZscoeUWVwK/Fq
qMY9zArYvebijwNLcdH5Zr7qk56h6sLi4uR8AxTi6s48vLrR+VxAxOTNX7axbsDY
`protect END_PROTECTED
