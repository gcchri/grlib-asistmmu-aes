`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gw27uI6EMfTYcy9UycmechFn8JEW8WMld+D7R40JnVAHKMkE6jfQ1m8NMwODxLEe
YyGv/l1H4kTRQrPGmZTXhHvwKYQz7SemWhwepFP3yrYFG6CQTziphWna5Ga2f0wN
ZJqaUp42Wla6O378EPVUYGa3Hlie8vI7JkfHRg7cl96YFEKw1Pg5CE9dUHdRzVjb
THqGg2kV20I952fZqVkjyZZJ0utQo6uA6zOqZbpy/dkEIl7EobTs2jsQqD1+HzF9
s8Y9HbGbn0ooHqdOBCQt5DtNIQOltcMG2V2BpZvrpsTxdgeAk0qHC6WyrSzns/9o
TbnwprWwomdjwQvrXIEwOglJ6SpROu6HCi+Q9oIUBn0abW3U+vrFWkR/qsxh2+3Z
qxpNMCdrtgB+ltxq/VPyPsNkRfNnonS187aiTX8YMzM=
`protect END_PROTECTED
