`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
egcYaf01T1tiuUhe8DrZjgbUm+a5c3b1X5O0eRLwTMQvKiX/w6rjVL23y4JApGFO
uXXN6kkf7cM97PrlQ7x5JGI5hbOh4IEs+YfcSOzOpcX9v4yW5chpvdRoFGR28uk9
zn5a259rZFFWEGo6b7V6688OBJe9Dlf+umckhfMvZTiHFGeMRpfUW8HjsC+z8o19
YmcCg6R4Ze4/bFeZ82bgXw+g9bXdmYqVwdqU7HoP0ZPETeEDdocogM8TMOKchdk0
FRJi11z1lWgTbcwMB980cEPuTNBjfUXcVxFefaflk4Smf9agPcbDUr6vzj4s46mV
qqyZjTN5ZbiAfZ14MPWdVpAszkmszC9yH2Nfp9WiSn6eZjX2Mj7N7nYycbMbY8Ri
Oz3jtfBVWQH2jF2m3VHib7dRXUgE7yc4q8Xuh9aZmEagm2wFMM2EIm0WDbKcTeGZ
`protect END_PROTECTED
