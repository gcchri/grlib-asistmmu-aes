`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
meChi43ehuSbpaYTgiibEWgsIkg9YaJDr74E4xDP4Rq/JafnVzG9t6NQ+EIL/syE
INHhpwL9eDKb6QIvBIpE24mJyGLOp33+im+x2p9R7GiHJ4v3X0dcCZL2WmPitSVk
qVgBgv8ULQhoawDNfPnkNDoPFjG+91NBzacck7gDC3IvihYg7TpSJu2YGKkYPWom
Ikkaw1es45j/nT5xbb+Es/pyM3TdresgoP/VEgsO7g7r0xMPiusICSFuY6mttgan
IC1pTGf8X3TAx5SwE4D0Oydb+9zUxGWunPzpfwoAcwRIk/bf6/XF/HF06kBVozE4
GIV9gIUZ71olA/mV/62878plXxUxm3foyJSPAt8OSSSG19vo4RqrG2yNX0MXXPHY
sLMIWiVEEWIqwB0L331hBR9D0Kw6FAvct/ubOwrcYnswKU3oWlXFgCbD3Oz080Yg
BA3VIHH4wF5HNLFNmQa3fuvFUh34QZJdU3P4nRPznP1G49rqhC4RkahWwCWLvkKh
Fm8pY1V3GXTPYUjbwzqJu6k/X1mSGc2/ixDt0d1G+xhCJOAEDvMEj+R1lMrPpgIk
G0ReNwAMulVjH3dG+fqPSgwgKbkCcTGwu8YzTkg7Q4d1cQQxaWaFtWrImFUE+RJA
H+jUkDvMZWN5z/N0uxeKoBvQSewiXYg0JHDurIgV/dSTizyYnIW5IJrAJ8RdI4tT
wg7vF3OKROHolsOxmY4qeQlmpwYJXNb85jIH2T3t1a+69GduwhsERqQqKN0qfbhh
vAABycFO9NJInfjx/hfSve2hThZc+GIEeHJ570/DVx5qNmcu90OTW9f3G3a2Siw1
RZgUosxF6Z6zk3asyQdRoy/dd91HHUo8ky+Aq6KKc0Q3gr/aQe82ht+iTsulr+6W
kEv0/Iy1z9bgZvzSy2PTfmRQLNchqee9AEPo1WFnHZKFkMBgS3SikzAv83sOrixk
eAszSL+M+0tMdoF9SdVCWAjCVXlTzgcGmjmVz8NGHscuYxf1PzTavoVQDZmTa9PQ
yRpT4VHnNTthwx/ed2KSj28I2GvTRr04yrLxq5vHjajePm7SCrQgkA0H1jjvJ8+R
7yYn8ipvQnwNHFxCdnXRfK+aif+MfyfIciyOZ5JlvELTr7M6OuGualxZZ7zheEbR
SWVIu4h7zycvHPbX063Vsa4WXIORs9GMWyT+TwLWDMyqLlZrotc9XbWSjxyYaxdr
liG6GqxP6hZrrWI8fc4Q5M+o+ZMM9ag/jf4/+Hl8HYJ6jjR3jaZ7NpfJhDN/z3bY
e5S5GnsJ13Trd7Nm3xO3isO9WOqSIMsBXXf7b8TWiPcnTEdy4xQ03JCZSsuVdRQ7
+/HuNAhrsDVbvkHP8fONIP3Ewb+2r3AE68u+TxKlLDr5PR/4aDaBXdoxYQfMpIeM
4gREae4DYD3U0CqzJS0lpq8Bh8+xH66q6MoFXmKKEGB8SLg0qInByzSY79MnGHY8
NCGlrZfZyM7+u7/CJ+3zk5JMsieqP6M3pLpo3DM5HzVguQeJjytH/c0l0c5o0ksB
yWP4O7j5nj/slAHuFSYrE9zm8GOM+nl+pDtPHweLym7eiLpym+BTGLfZ+bks5+59
JHcReB5dXiHtJlkH2lNuc50k7INfs7x0ZUlnm1KyinsHCc+EL8x3YRG/TRHmqsEH
Cgmno9nPNko4/hii2RSsScnLCMYjV7C0EqneQa8SyBjuw2iOwENW2r0wu/y/v2pD
wSzoHT6ZgYhLdsrpfYJmHQO+m3MxdwlOYYzVi/4DhL5kN0LoZqiai8/1qXMBqtg3
naoPO3VO3vGNWK6FWUfXw6/BWiFSylldHS/GzsfBx4v8LuWKmLJr2zYQQZbi/jJd
zKqyZJ8zK0MReYabPCf0eM7mmlU6G9gFidXsNm/NMGEqx4WkRdOBq4vTrv2qRiHA
ALZ+MP3i5P9QIBF0J+XpdiA0DzcjMpQCPaggwpceREEuECiY8vysG6bb5xF1CPyk
ffIkFIbsb02bFMyx1Xs/klPuV1V/vIW/FeayVVbdsYUamMgIJ6pkziv5ls3F/G4u
zobLBaQl77rhJ+j7OEVTKvWRKWqepi94dAG1oCl/hmjM6rtl8DbLd1UmCz6DFnx2
pq3jq2AbpEWWQf0LicEc+PmQ1CAINWbgPRx6amMh8njYlk+3zhGFSc9uyUT1bcI/
pqgbTQk7HzG041NaijGWFRkRZ/QyeAmjyuKO45J/zufFk8NoIl+N+36dg7lULofp
JNj8RHga6aa+o9B7olZs9S986BfHpXXRDbkcvERhTdITfRGg/GVjK7E/C99py71b
JQg7zCyealqXZIRNYUiJ5bh789qFQcDONZ5h+30lz08GyGAxEPBGlVgPhUrpdA9O
cH4FbyzKr7RTVYz2a0oho+Ljdr/pwJcGTGxlLlhZVvnu6g9/nsvAqjCGIpOcm+XE
5ZYutVYYHOp6fUisbyXeREPH9oEVvNT3jyVQJhdjkLtvAneVMUcEvCuIoJ1Qg0mj
fxFmQyQA8yANfdqKqcltWfD89kqpbulekR5Qo8j1L2ON7jL0uaYt86pnvfBCK6Na
vL4t5QjDvxkA8CyzBmMIaiOmrtN8Acd0tzVwsti987LCFVA+KC7fCWz+upkjiPee
jN84bELpR8n1WmCo8ntQ20q41MrZu3wU56cI2yFtMkIOePCtPvyJy3PqYMp9Ea4m
hJiFrYasv7QMj72fhOTTiqyhdRdyfCWt0Ww8Dw/hYnr9mvBHmBkqzGHfFy1Fne40
mKcv8YyQ61+fJDJqdCkvBZPU2E2afZUc44AQFZ4isqgS6fNlylS0j6zCtD04QTVO
YTXT6ZLNNXGG8Z1TuL1Hfp5rqfonRTxCf9yFS/3w1s3oSw6OAUpNYk/rtl90lAfm
vpb/vovBctOPu8lnF0gZYA10yI8VBN7ddw4nY1fwisnvj8HabAurHFnC6DHIIPJF
rrRYdB5UTFr3uHFuibshN9pMQ6F8y4lDMiQawsmpTWekXaSevxPnYdVCR0S8rt0r
VSoRV0uh1je/6Zv43UaI41VFASEMaXS8YskEiKnNF3XDnPfVl0o7FyGcR80tQoOP
GzXxU39eUiFQ0TsD949VaD/RgppAzHJErC5jYgW+MPST9OGXS5Gsb/NNiZqqFcI4
su2zwVPKrPxMWshBnFfrmXXf7zqWIzeqfIhCk8xx7HU26pSweix+xNCkR9sBq+3O
QhMykhopZY+XMrZE7F4XwwcRzjLYrDJk6UeoHEBNfwUlLBpvPFbg4/qLJNXhPmXs
BIIaPkGB+aYmqi7xvUeA5KYxEvBMJF/jSpHwWQxuObFgzogKTbfLqZGuA+d43Var
6STk6xImbUVl64QRWyog7ySWcjT/vHDok4T9MdeVB2d/cRbgaOpMI/nCMvcjQsBv
+5KRFUr6p2qRrYDRCpnz/sZzEAcWTUb0lVo1XgNLRLYtMRAysIFRE7xBj8/Tbnff
Z20NJtW74qgG08sANqhXTm2yBBUOYngAL7lh5+TRhB7uykqetyXIZxVqznYM5K5r
xAl85NXjYz7D4F9MT8XnurDNc+47AVrxJAZ6+ieAGyTzZoVW3RwvCj1T67A8XDSp
wzKwStk53T4ma7qZzzI0LGMxnx/poZs+IPDw8KPkY4zVGWLEElFnwV2pahtaXDUC
0EZM74sqsGoDlbOVDhRgsRnca+qspb0JbhUqTwVWZ9dwLzcWnfiG/Qftakfvwbce
BTB9S7C2upWvRxoswN6rTagZAjLm5OcpuD6vpT4G+6jAL8OTTs6AIQ5Rtn8WHzGy
WUbQmH+J2dqlQUeXfLHpSIyzatWAgzg5mC6V91SvuBkI4OCXATxlpVPz2J0HRiZ5
8LdyNaAMLbozwNs1fzVvDi/rAVsdh67kcYRji9hqyZeJBjXauG580jCNAz7HQAfG
PKLw1lEzGYZUcLvPuhN+LxUUigKzYKVU8xG23qpPBLhBB4gTwPKH/fnUpvPcdLl+
SUQKPT5RNNlxtEPPVhERcZV0yp+dRIXWOpZcCWKevXnuZSymHclvh9AOAwsvfv+/
lT3s5+RUi5qCeBr40xu5ftI8KFMwELeVMUEd5xIDY1vC2XTG1jSKem1vQaYBqxlS
9/3jiCywx7lN/LEy4PJxuTu4r93SSkaItBg6SAKvFqc4TLK3I+4rhBGSsaNbs5Iq
11r5RSse5RgmTA/D8kg7erlvEJa0SaIcZ79/TMDBxvL6lISLhhU49wlnMG1eOkAo
lG+JFCfl57xOqK7XJlT9xEf8SWV3v9/awvqe5SfOxz77dqDTm82qKEILnXVYhHQw
Qt614cw/rYpiibfmvTpw/kjxNPmY+KCCsnNZfV1UCbkjBKF4VBBXkP5Pf2NGJr58
wyHcsGn7sbic3VeY431QxklTVRM/l95sWsGoTi3+AivJMAPVklkmYPFCwVbltYK7
2DAl8luEB81NHV3xpTOBEidi3Zy6a473JtsP6VrieR0gb+M8Dwjc9j+t1FA4xj9Y
cNmkRsQOJ6N3Oq5cv7bmGrXEIAOhA2Sj/s3t/MlYeNFhTuc/Qspxu2tdfy9o53TT
HorjGSPHMsFzxUnvae2oioOcE9XLlJDEy8jZ+6Z4S0t0ZZxSs8BPCpxwHy9zCM61
NOZn3T/DJP3vKhMDMFDKDTeQyRXWz18oqpVdBnJLAlMBhZTPhGTVk+3a2+JIxrG3
Z7vI9X5p5Rei0U6+JNBrwIevmJDlPP1kQHp8XZh2OVAwmR7N9xwE+QXix+9I0oGk
emGsfeUr3adIBFyVVcn6hr0VQL8dhI4eoqdEFO7+1gSoqQtcu2UN8U2/Yq3PeUSn
j/K58ZoyZGvOhNFN8xfNdf/ujuTV26TF+8RkANVGFRcXShtpQ4ylkNV2w/1o0F25
RipZjalbqlkPl5WFd4Y1AXvLXo4DgyIRO2nGC3LtnRt/0AUvBOuNjU+2F2UMe0D1
q62Q4O9frWTmZcUqYxARu0gICPbf956wy7P4bTye1MGWDSQ955HHPcQYasDMBBQT
0Ii9Ra6rZ4TYJope2MPa5e7ieQP4DPwTMINJq8Chkbwe98w9utYMsN/oylKJbiNY
asTC8lMNdHlleUO7WWyz1f0ZxSr5udvtS9WS/lVuRLy9TKHQOf0Xno76Nlw/p0O7
0Nsg1M5BaKX/gklDy+llU68BvVHewPeDhcRIBjdqQTHJE/s3V0nZTNmU8vmT7NGc
6UB5//PU6/lprWHXl7CxFD+OMb9p7F7xB2TfuuSyhV3fqgxZv2EitSwhPjuWfRqQ
Ta4q7LbCKppIuuIuW1yhYBNK7PeZ74AWvBEMoQoBI2Wxh9JvXWXk4SPyiCGZd6BI
WUCSb0vhcXCzK8zfqm2mcoRRzZBdMXRh3iEWOs7YLkLJId3OYScXbkgATobFFNig
KoLG5prjsDlxPf2Oq52lCtxBGclvSutEVKMBHD0vl6nS13eAgz4W3sB/yXgzhe1/
BpmUmmJSpYdcCDHnFNayNM+mOADvHGIdtku0BFsk3/fb2QvFzvTVXnQE6PM68utP
KxXKdlYnvMy4ppIB25FsgwJ9trHn/52ucC3R3A6Hpl9Ko+VJDMBPh7rFUnjaswHq
DY7JvqZOOzn8Y/EFbDeYGbd3eLBmUhx8KXM9EFtzIvX/3qFQ7xZBNDeprbAb4Kjx
ph+Ny8YREOY0uc60tV4UqTWiMLjMZwtmm8ZuT2xTPDZRwiNlzN3TKhjYXg8T2mNP
AnFSFyzVTng4Hq5KlmUApOoKQg4MEFIhAq9iG103J15lS/rW6KTFCdbeN5c7IjeQ
+ibct1Chb+l5t1BFHPUVHb3gad2IK9cfbC8e9cDbyT7M2C7RGCAVo4eOwe5YXmgs
cpdbR8OciIcrDLVnkRLAPrUWAkx69/OO++q+RV3sgaGgTNsc5xwHja2A9QIyGv9c
5lVbUU5hxMYg9q91k/vvdH4p91xdjATYFNfiLM84THJmoxh/72cxO06f6oLGGL4Y
6tS1rI49xf6TJ2EjKYdMVM02xo/pB9hSdpYZeftwVO8Mk1qD4k3G3CWj8YZ6hRqB
uZD4zYgZuD0qLSUAtRclvZbeWsPiu5dIhIDL5L3Lh2tqTLwT2EbAVme1WFBAKxuB
QQR0EVY4N4Q4qQRyekLjnV48cqKBoGpEfnFsTPwg9xEYB++lLYiuwDhNixGodPck
g8CoYHJapeTu491Xz3JJJt5YKZ2Xy7liHnjoh+5TsIPA+YbqcZe4DvvH9Ev14nh4
LsEgL6wLt8WxgzqpK1R07jpG9i3nGzXCPmnffWwlTtKdl2CFRPdhVbGi4xdPJ4RG
3iNemKa0uGmSE49fMNdxVZT5Lm/lW/wqBqsnW+usqHplyrkcHj+AXbnhp277fH4P
us53LQ35XSFJsPdr9t4nuPfl0mERGUlIh4ZvXeSJffdXK3ntcjaIPaDWbA3BC5+8
d7dOr/U9M8DyYspFglRoZSlRhMLwvoqYW148Ykoh1lbKwJHKKSBoQuXeVhSo73fP
du79L5HB3cx8tjF4YuBr0VIr+i2SXsF4AeCMn+rngvdk10Bqg2LVZOpB047Z1k9Y
GT88QhrKIdBWeUJT5oJ+oOtHq/tqtUFf3ikpsScbzzg1/3Rrr+Dv9FgQXzSGFpk2
HU/coUSuz7SOLE7HIMWYKscogminYLk8MDX7rZsRCuEoNGXWCU+SmTU1hK5nzIO0
bnUI0ZzebDCqUkdHP5QcHwsSty0pr3Fs1TF3ZWrFuM3h6JuohBgIAsdnRfmzjBtI
MM37IfeZOyY2yYR4OvirXH+5dMth7X+UiMAHO/At/WbcQ7LRXdP40l+6cM/FDpB2
ffyuGPdZ3XaPoGQ/hZbJbBiA9510OI5HyepNJ/H3+m1IEmOep+w009wL5LlcXtYH
I+DTz2OoIMGGWkAMAQMjvFBwutIRqOOJfXK+1Q9UHCYQ2KOZC6bNUPN8eQWrRqw8
dOTZEyqJq94t2un8G+1mAod5tUTkqLBaL88lXhFqNFmL1AA2YLOlX4aodPv41Y6u
quqzqNK9u+Mjc6K3wAHBelhVWmYUU6QEizIFVjpm+4lVXDZKX4bfz1jocUdlhWCN
S0r4+CzGCBvAeNXMvRarJYixeSC+gtW7D6vfoM6QkcRlKNpVyUt0iAF9KAGANKll
Ts0sIxKZKFGonLP2w+CJ6+cSujWtlAh5PMFXSxJ/zVWfmqC/zEQcoFo37qruPeac
hEa04pw0vH78zDFeCf1Q9ikECOl7Cy+aG7mMxLSrKQe7kCuOi+I1TRZuHGZz8UCs
GVK32N1OXFVoPB7LIf6MWYeX1Xu6Kl22v2GjNmLOrcwU1zt0GPKC+Y5RiG70KE2N
f7e1gPXFWljYy8uiPg2oap/fP5vhU5N+G7QZ+J+xkcv7yd1nL+Y0Z1sNHJ1KAZL9
YzSBEoCxQxk9aWWcRv6FpnB2Jw9LtDrw05RECSmN9FfQqIWhi5XRnwgJIdcnsWe5
GMrQ0b5Tbpdgmr++4MPjZoxkmMPxxyZ5tAbSPPAxnItzzCvgJ6g+XjN/N9wJy/X6
iBuP8BLT9v+ZFDwsSerMxtLh3Y0OBWTyWHVVbREuwkkJKiI9LBswC6978JXxVjPG
oZ1KchMIIoNuOKPhttRsmv8bwCzCPeUiTnWObi9zx2c6fndRS8kb4YrzG6RSnilU
wOpyt96KcEL0fSWHg3kmIxK/nK1qY0l7KNBPlWMbpfW3KYuyPLH2F4WUmKi3pRvr
T1lraECSsZrXksu4V7DtJH1ngnHMS3Njl73u1+ViZB2lX+fIUj9AzvHyFYhKoCO3
uRERkP21eommz+O7AmL5t4Wtk9Kz8hOR7pc+DKDrRr6mJhEC0wUpUMQVJ92Vqz0P
CCTvyNvphbCpbTmzoRHk734TJcAs8VuQvhQKkxUaHKB02zJBBAxmX2muvwE+i4Ik
2zbFCjpa4ySi6eOSneFI63cRs4tNXWPHkOR7VNvipcuwnwZt5VoJUpdZvDj3Q0bo
6nN0MNmgf1dYk5Q4dQyHXUZYl0uQf4UDVw+haLAwtG96oFld0gJNoQ307bwTPMfO
CxNp7aZTJC4CCHM0pqKByG7bI1cf80whoiBXIEAtLJuh1SC3i9Vtkyit13ipGYwP
lEMsnzN/OdRr8gdJCJqVAnThHyi5QAfi9SgubHdZql6OqqYwYV6VSkbch0Ovey+f
lz8KFbVIMuUya9iYNTv5mdFxeIyhjRRGaz+/Ja+e5uvyly+6ITirUR5LvbdV0PCc
iZv6TnYIk9xshbYc1G8dB3S6Jg6/DXhFJsfrN3BUmcV0Fs88bN0+1IYXtDjtMcO2
0MPrYc5uXJtf46aroGlOURwaXPA2cPtM17/cUnYOqMnLWGdv3WNsBRlkLE5A67Dx
HbmHHWBfcguhiXCzZTSwMH1TZ9mHrshPZJvthTMAdhond4ZMaScT4kwU8QiIPg1p
o5lqX/mFiby9WORkO3XFUqXreq7wa3xxtQcFePLSu+dyIWFDPgvm1eOglNlJbRyB
md8tbPoSLBGyso1pQNuaPrid4XgWmwNYCoA1wKZhV5g2soQmoinPYdmqhgqKliD8
5LvqWaHGB/mwxqQuFsJwQzu7WiS3aSnBOzjy9XZtYZMYgiQQmtXgySVS+JGY0o1E
14n1X9p01GCXIoE1W78GzKfMteYXajlrXlV/UNv662pqOTZZkluqtVqSB4iUrI7z
Ikrp0sPSPJZMoPTx1e0wYQefYeKbGqjvY9BLhRNsjJ8oLpCtjWOF0zj/53roGjH7
EIPw+OyrjM+Dzaj6uJtjdlmXSB01FSDEQilNXrPMHUvQZoNQROybuNa94CYHqpYJ
BKWRPeeHPI/J2NnRcTxWtQRGbxRI69FJkG+OAIICNEHlZtR7+X8ZIaZB0A5if94n
5O0PV5u6T0PXhZgzK61pEIxlH4sYTvlE6XS3mt26GpT5wZqR1mcdmalI9CMJVTtS
1bW64Yimi6d+ha+n3hbch3YpcV1jVJaQXLV5co9VRk/70NkP0M7Gz6+YrrKr4aml
t9nV38Qx4yix4KFEx6SM4uvIBDe+K5ztQTeGVj7IgAiaDjt19Go/Dw+cD7tCaYMh
/BdwsBRT4XuAN+ax52L4/Z0e0HgVCwVd4uN99VA7S55KcMTU0ii/0CRAmJnDwGg9
9BYGTTBPOp9z+HeQlKQUlCSuv/BBOOoUt+bkJyc9zpMSTi3ENx4OgnylTJydVh04
gLqr4VBdQWYCtCwhCWCwB5LfX7cTgIwVikjykwg0Oeh6/6/T6/LfJ+cqkR+Dx3El
A+KAM/GsBRUfMnpq1Ut57lfiHUncEC/MapmnqTwObpdcN5WIDgJ0jpLJa3wwSVWi
UJ0epd4wPfLM79wV5F7CNzmYviDfqXHi8g28sVvcTgznydFSbczkBAbAEgN2wHU+
DytWAQDggAV1qPk8ZR1jKpePeOWFt1lHRiGiKbfKcLDPNxX8oR1MPbf81Qw9AhiD
Hw0Y9qxgKzXakS4FIzBiBgFtHeD8MCZwJPBlddMbFo9iUG3+KWNb8E6/5O8ybF/s
i1rTnE9HPtLYw62LEQX1/KuwihI5d6KXu2adIsfsPwTKIEseI9hhPTSGdpeW7woI
cpSvud9YJrqJHvZWaT15MLnYJmherl5mVPQjSykPNsMnxw+FC0hEnc87Pp66KWGR
pp6ihoSRVXLK2ngfRjtbN+g+RJqHW6XfxTUPXV3WLSSdjqLcmE6v0j80L4C/7ipn
B5L11asFxiywRXH53FmSzpxKzYODDGjFrPFAcb7V5k+u6LIx+rSrT4G2NnB1KHSi
bfiAPCp1SnMY+JqwqRACwGhCmovzMFvE5CV/bZy2VQwrTvMvN8K7REGVZvLZQOe5
8n+FhcZirgbc+iwizV5FherV7IeVMZTaGFLo0UTRCSQ0O1YabvvjCi72D784gnwf
zXQO+BcjmymzBYdF+5jvbJ7TiWS0xw6zduB4wGiVI84W6Cv4XjEld/oCvPWjX3V2
1VrL4FfDbdc83TpVrh6PsfLTWl5rRVzC6bELOq5VggfBi8S64+5IHLTjUjbUXMIj
rm88iDxmfAUAVwGvKE8ED+hwWl4geWvNtBLArec4F1fdjzEQggv7AL2kxWFe9ZW1
oKGKYMsNYOXSyTYMLyIMpivxy3RT/l1Utr2Y2ODdhFXrxYaxdlABpyPfty5r3OAv
o3ZnBSgZMzFETzQJJKhH6KCeWdagBIvIYDhpKLn1fbZqbjT0fOxnnO6Ocudaz9uN
A3EX832daOyf0BzvFSYS9G0p9t3naeHnThvZ1mi4HGtkJFX7IB3qybfAV9dpYwIh
2Dv3IMs61Zd2ZhiNUNp6CpKQhhfwmjkRWLHVEaiHt4JjEGZZU8sGnWAe/zwlAKRY
yYD+7RZNd+pl4az8+KLxJU0Ch/MewPIUaeuIPnl3c4pLAcwsOxr4LCBwQ+VtmB5X
ISWIymouBYRP6J7sWp4vS6Jw8+IZTCOL1BK5WPH9Oucuixhv5f33pMOF/0qQEPd4
r0olsiQzeE6ygWsgmTP0gdICg89GAbswVNqTa0FOEsRzUlHyZXqiYj68KfO6Dh+3
LVjUUv16UX6F68F9bCs6xUYySMuInDr3WahzdrKNxmsLJ17Saw2OWFEaiMnUoQGB
tACFSD6Z9m1FwIa81qrlIbnrC2yRt3cC2cWFfz66dBOv3PvTtTsKUR4leYJo8c4D
AcwTb/RgpQG4IkdVPtSeKA2F+7a6d0BOrDpO61gMpcTVpr9mQamZsuf63YRVDPK2
3P3aB2nGyDkE7ddAV9peUsGRz9Vn2OlsNKHqfAeCPIKYfOmTda9errGk5zqgHntR
KPvWgjfAZKjCNt7AOeExM0emCyMzVpiB0Oes+4yJfJdguVajdGzOurj+qTOVIp1m
sU9xE/M/mPHafqcFxX1wK4Ef+osu3SBNlgVcy21A3ZetUN7no6QNxNBgapbHcjSF
r0MK4+1PcaOIOZ+zvrU+2hrE4BC3ABMsr6otj9mFzqRka5htyalTehptqou2ebHg
YHE9Lt/yPx1QTIo0ueMOx4whknH+s4PV3dwMZeghBkGxT9OUM84jLbzaIpLG2hm8
cUUaXs8cv4JQm62CfJmWdCMORD7h49xJNooAq2yIT34EkI8NKN9Q+qFrhP/1db5y
UMdsvAH7FfjWaDyae2lXvLoU3AhK9kQi8p/BVe2j5o+GqtCAiM+lT+2h3yE8O3rS
C57ks05wt5PWI99+fAQP9ItjkbsNvdv8Z7b/4q95GPsKmnZagYXvnzjRl2SN08bR
vQZAyw5eLa4w1xeP2FOtqwgwKkwr7vMAlKF9LJbUdC2AWP9Q5gT8VfEQWLyfczhr
A6GwNkZsELhHcgtSb3qhyF3MBcITbrZWK14TaJJIREgt3WTXzEQMijtZv8sbY+q4
k/cP+5xhYFVjchx0ZDezuXGnSp33Ry1n+ZgbK7IFRv2/1ybyAJyolLXt02487FFr
2yUgEs/hJqFsH6TKCY5G8V3fqU+fwrrMmz35dY6KoafLVmgfJ/tc6MaxywNCZ8+y
ne4tXPfm5WrhYDS9l4FQwWs/5QjcV0M1vv/0FQ+Mx/Wmug740WZhGglpSPsbtwwY
+hpc9bBX2eGii2pLeg8bUZm8EtxDYUihjAX0wYcR5ZCdkCqpPiINZ9EL5Dy0ZhcH
uxodDL0BFpYmW/na5Ye+BrzvSUxBRZOeSVjg0k+6qbWrY6XKBK4CTDevdEpFCHAN
t/yR4jEir20Pr30stBvGBJhb94iNysEceLGEOpt0aaU4pBrNAvyMcrgGLHPMBE4s
VhkNqPD7XIan4af1F7KH5WhzHIYr5vat1+y1JEx1rLKcvJZQeQsK/Bw0jnGKt+RB
YHmQL3L4NkMbyEymKgAddylTX3vKpG9s3cfrfDmXZZuL6lEkESeOdQev67Mc2Wn6
ekZ/uT18YniDj9NBgfEZflj3LBjFOita10qxjRb3EUadtHZWtfBbCXYZK5FHTr+y
zGqbBDsWRPquwpayPJeDcQkn294MafoEVGr3QL7DjgJWiqiEd+ThFISP9h0VNIKy
6YNc4kgL5NLZx7RPpnbUDEEsri9iydIH2e+VODzkS/0hsYJmTV7kF/dhaNEJAl9n
BqUO9GXO0yH2RP5SzNO5ocI1dYsg5E1bXZXtZfXrx9Jl4DFtdS4jvPJDAzhY4FJu
TtcM7qS2znczpNslh/8xRJo2s4KJDW4SujglxQyF80tYj+Na7Cf9Crq/SciCnZaW
QBcQj3c0eqXUbgwLzja3F5gmyrIUuMwYfhlfUwCkguNo9NpRLlCQ2UZpeAKCndOb
L0V052pU4Q8rVaMAMkwVaS75zevgTRcWqMxOZn9J9udgveu0ySwZZxD21K3WgXXB
RDyP13QDdNULA7mWfjxiqfFjFImCiP7RKwy4Vj6Qjl2vv0jvGXi9rDSXSECcRbGA
68tqS7G4kpr7oT0WE/3Cr6nrfFHiSaNjZwiiRdWxv+wavQ3F5Co+bdDZESw+UEGb
aTuQjWgCUJMWV7ildAJKMNWEnsBmRmZoaMw6nZGo0LD/Fr1IfKVc/Z1wFZ5e5iOE
nFvlveL2NKD2S3Yf6LwsNsXHV0K4ieFLFNIVnm2rZ/4ZrPxT0js7uFIUIzO2VCJU
6oJQFC3Vnjgs/OS6tNQqkf0BTOh0yE8SPPXh0RmaqwacU9Oe0NA1YMPnG02OIinR
wERaMXHoIuXwt6JvQrHhRWZPwrbiPPB7CMrOKcxaOWK5y4AbNcA+E4MbRyYAgvux
jviWlxbWVbVaVe+BGbDpGG3OYdtl7Zdo/Cne5v6FNazy8xLfDcS6iys2A4fyGcyJ
XFtOpE8TPAXw5+qq2cCkHSWz8s/US+jvuINfEFlFrcknl8mAIdD19f2Hu97vVSH8
/CAoMwBwn7P4X1QcmUFGAIqae8qJ9QPR/hU+aGSl62K68/K1G/tuN+LSKIW1Fq69
XgzF3aHjrGVnwTz6WGrv0rEg3PepjaYuv6J8FGdB5K1D9S6WMEqKGR7u/2oX4hb9
66ZXrrkG5b7rngo0xBR/loy+m6WwIUcwIYeZj1FxLU8Jp9w7BJm/o82M3HoOg200
2RcjwQevyu7mY+5A9l+z6Yp8HZv8fOBfyZKa3aPZuOcL5PKrMSlQNxxDg71V+YSU
oj6dxKutlki4OYKfTbBfjVd+d/Afh2wz0YgD84BUC4fATPL5AzjbliCHcSoH7pMk
iIu2C/DbhFrzJKrOfg04+Qs7opfe9cmmtOksXx5sQfboadK0uhBTcFb8kHVU8Fnp
sjEEJYdYXpiXMEPGTIZjd86JAsNDbki1wR5qODLO+CISFcDu8ztVNbiKKJtk1Njx
JASjXTRoy9ID8nI9SyGBsscic6Bqbul4AKKKxp715MS9JaNJzqViKn2rIYpapJmm
C3YwZEVT6iE4JVmpATswD3t5ta7C7JqRMZdGGdZwsli5gurWzWoxp2hI556wCVH9
uwjXTE1C+iLC6LtuLu9/VsXhrvNX6st0qZSXed3g2ZPC7yt5G1fPIblad6mPa2QS
mR6Zx1DmQAK0LcplTKT/+dM/3HozQqTbxBksCiunwbi2yY83nerZqEgE6c/JNz4+
wa7SYzGc36n2tKDHKy6aI0y4MW5leZjvKfM1EpDKualqVtiRMU2yDMd36iysTtPo
kERPY3UP29oJG3RbYDwodFzY0+C+jswFGzyC/CxsTLredWvFnFpF+Ps4tL2NoUqk
g4IVU8hNa1oA0xZhIatxDMAMIaXeRGFtCvJ4QWSBvolfj/NA0U7AySkAJwJ/DjW3
CMQWzXGYzhkmIfKIF8voJfhIhBk+mJOnN3NLl0aqlQ6ExEojlZDyyCJ4aslTlZuw
SLRneURL3cAa9LyhpRVVe8J4scAjn6Wj2LpTQbhql/3IGJXprxIRA+pQS/10A15G
yFuQEbVNSX3zx6F4qJhfNkoNEOjRoS3CwVWcoWrgd9qj8NXsSMlEFcPvmzs+FfV1
wwrFHXOfeA4cEC0xkZWa28K5ZKwU1stbj6EMQ21UfUl3jdLKg26uZiRP2tALkEu3
pLgt/dLFtNQE014igYQo4QnoZhZT7NKkNg01GCh6MOSbnXJXIX+EMD1JBGt567Lg
uwTl1+fR8hYbR5+e88pWxto9S+4mJssi1HLrC5lfRNPQT9Qrb/eu8aFj1KEchPz+
vYQpzVl5LicBydqB5TV3p5MwxNEr5IhZLgL54iqvEhOxBTSaIgcHscZRl+muzH8m
04FINSs4nrtIT+27I3lYvDvyszRfqvnrRxg3grBU0jTCkj7KzOu4ZPWkkl3F9LcV
G6x9XdJul4RgwUxO9rUykQ4F+wZLH0jBcIagZOh2dIt69N+1iDE2VD5h5M2gbzd9
1h9MOP5SkA9sLL3bsq9xaEqzCf24xVqzKIq03CqJ8zEiq4CYtbjoQuzOq1csjCAV
Wv/Wvwua0nvEj+0R3/SXwF5YAMQxhD5fWDHSUGPJqWhVApT+DFzD8q/QoJgt0DTK
2JCGTAdUd4L+tdKSPYjuLx+HUl0uyty8H0L470m+eh9+k4kllJyuoE4r3Re+omx9
9f290HXhpRS93SEEaJnznRaYDfhXOmjdIcXXWEC+j1ykH4A0jPE88ioBCHZyrjJP
B6cOdKsBuIoL/O1+XQip1YDMhMJa+tY5j5iFLleul78/Z1zUSy0oYueq96yRI0D/
9qBnsgoI72UmH/RmIt+p5YMEFJ6TwwAzBQENTEQNwcHBfUbqP6pA6420cJzVQO0d
e6nARDEQBBIU3Qewz1LDZTGebMtdXz0KSq3k0jvSFOuzXGrMBHSmuwDdrAer8PZ+
MNWkawse3mjeTektipx6X4oAFSbWVTZkPm6ao5C3RqViGtVGW9kAn3EV22Ydf7/4
UDQhJzPmvRtKYuxJ0T1huCIrnNHEkLOE208mh/lU3zEjeALAeGxUjfvwA9+mNg4Q
ic1p9dMCiy7NTQSrPDvtRCr7qJ8LXjeecpw7VhtQ4AJxx9Q7if19uRPjxyiWWmbs
NiuRqxgwFdTmnH/d6VCYgKL2X8W9tm/j9EcJ1Rfk3JZgF3xQQCuKnC/C4VqNfCJG
hrv+PtD9nUojLtpIM4E08ggP0FbW/+pYB2JK9LZUstfehXiMgjrVEyqd0g8zhohU
bXaiSstN/g00VwELjS1FYoR7lnsiTPvBawTVMzAOnL14DQf2MhdZda+McYgn/ZwM
o9BiA2REv3DHaKZxrV39h5sPeJKG+MeWKGY2z0xVkhArtTf7Z+V98NLn6+OYOYHj
DE357KLrCvwLlmMZCR1QwR70UlbGPT1GvedW6xfE7o4ashN78bikEfVvfkGs/50J
JccqyrNQyYnq066OnDafGuHdtesQR13ijk65ZmPFoKTjiEpnm6XLg4bYm/DtpopP
gJIRr/qbLDZBRT0mTSq2NIKTsj0rKINHzDopR9XYdYINl7ArmwZmWy1mh4OifMCv
ZpQO97BYTXetC7cf4sYg8jxOk4lonLEsCPpAcBDDMITdLkYG4HKayVqZ63EGOwyc
ZYU6AKAuitKBBvhmPA/QB01w1GxYK5Vm2OotkgzNwglf8jobAz6wE8MSPbLO9+m1
o3U876Lwer/GuxZcVZyYXL9H3aDqPqD0xuLELINUBUWjWcVVxCjkaJv7UU3gPMMg
mlOPrBg0BJVXXwqFHAJ/RkOjCkvNkGWw0tRIN8mR/0becGCaJAqb/4eSrSNvu5Ek
l1Xye9xK60Gwd99KSuU+UfP8Z3VpKxv6l2KtLyCj+yndP3wt10HF36JNu8jk+ZRo
5CigUhb4W8fxwuhX/ncvi13nCSP+3VjaMgcq2+Z4DYJzABsd+vYGmXXcp/2DjgIY
JrVcjzU3jm0KVZkoz3iJm5pd07efjqvooiC1ghEI8k1jS73ZQNOpR6c9525AXssF
2zoBv376zUY5/M6gcbceOj+B6uuMFy4p5M9z2FEu3HRadc9UnIkx1nsVNCnagjJy
I6lntoUQDfUpcS5iRdv2RXfQT6RZ87TDer+YHYUu/nVrqpHqyson6o6+PUINQO3T
gq0fRcCwDHiVn/L409Ch0XjXvS/Mf9jzrbuMZwcgshdpHwLxogVv+ZYp7exIX7OL
MZ1BWNuMbyc7CzDXXpkDzo5nEYL5qPZbHiIHyk++hMQXXdnbTCtkYgeMECVfWFDl
KHiYc8KAkcAhwh+e/DHB0nbZUchpvE7mYZGJFlEsNxIUVomLN0bSBH2F0jqSyvg/
sVQwNxC4BN+J44ZnpsjQ00QdyfJhdWVlaZkfJuXkPABxyI3QhUUp/aOeJo8QFXvh
aEje/ss8SbCafUZjTqaXf4cbXx8EkbfaV7S6Ynnskwr4Agqiggyij1aUeBFFtlri
TlgsxY6Uhpk85zvzExEwpItN3ummwg0zcYJbUS+k09MzYMtWVq4sNNJYKJriQItD
UfW/ZRRJKxEWgkiCZ7dBtnl2qLjjcCNRerhb1WlULHyoaRVLQu3B1oWvlfd3rNtv
hP6QHqZj2YWAkBXA7OA7EwrQTd9XR9NGkJCfzc1pg68LmkcioSuZWxGpPlBr+KBl
MWpJAB/s6dzFhGcp9y4KWhQJMnOoxk500hHaUyLSQ4bb3SqOBc+T3ka6/BqokflP
QwudwFdURsypeqzu6F3LqxKSfF2nBzzSXpy2Gaju1NRAFQWslw+cF4YANuceNAi9
NCYxmBCioNoDxDkuzU9pTLhALcqifu6Pp0TKpXd6sHVbbERLDK25Mx08QU/p2b7s
avek90vmKRH+6tiIQWoOjeYJi55jDrDz1UtLc5KQAgzzUObxWaB5ZoiXiPJLiZyX
2s9wWFFzT8ti8tFdAZDiCEv1bVE4nLUvTDboBjpYih7QwT5s+/mh1+VTd/wyr1e8
t1mrUUEEKgx87RDQ2ibvqdKjpFQVRQbvhc/tYa+rSH1E5YP55C47gHf3No16wJB8
AinTuI86dT8VkqGDQA0JMjp7TCEt2a+lXYmDtkSkPWWxoB1Wu/oerb6P+44wCtMD
`protect END_PROTECTED
