`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t/Fgeit6hVTmUbLVPrftxDrts5PtquMrQUX9yiKMPEnYFlJ5oxRTo0qk5DHo5bBu
+2LyezJgDTX1nn3ECGvw56T3ueYdilyWctDd6q6LKf6g/a8bn2lUE97BJG27gGVj
Ha/5jT0Wk11RL1whw2qZVrG228IhI1qkNVahaksPlT61Eww0y9cGpJBhZKcCrYmQ
zZhI4TKaklVG3Y9zccicbh6YB1JsgaffvAFUro8xIZCMCCNPdFCgJUFPnFGskYX4
EN0PrIRjyNzI9fmXfAMGitIXGiPqAURS41kpR4Ezr4o18gTjYw8T7hCBPc2yuWk8
z5kUsPZ/yxEkJHogSalXHYSQwFvOdP8wx6qpYZV3O8Gqr4JEusml5BJjQ2b9AfLr
GD6qQCey05STIU9qbTuPZgISPJlAebK+QivRmyDtvwnBcIaKwHpWwES6Ij27vADF
`protect END_PROTECTED
