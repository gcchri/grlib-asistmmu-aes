`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Wzh51M0et+vpkKcgcCoT6+QdI5AEcPEwVul9s8PcLL8Qu6cidFZ4H1I0KJ2u0yD
QmVa0gnVxl0PlCHNpri9YXGfLSCy/gfhFa4OdhIIlvqbLgnuszXk37aaIGuBKG1u
Kv804fsR9LQTK7NTKJgWKP0TDB26Ppc7H6jaW2rzjYx4scrO37jJt8eyL3md+uoZ
CkzzL3bA7hdLbRlpD6P6eJYHXewYoN47nn9680+XxXPoVbn4nbsUMnqR3JVpWMeY
Uczj1bsqGORbeoTRmKdU0If+bjYiwzat4NtThs/dvc3iUglKgTqoBDeNax1M3s2J
KRjV5PSxC8dHrHg+/Olfy+2jZ+7NLkPjjXEanYr3zUvGa32I50Is0ypN/h0aZXmi
CYZAYuamUT7OQrgcE/brVQFho59eQnEjWby5Xtk6NOvZe7GKqoYcwcMHc3oWNjAi
JvPRsgbN0ciClsK+FxzNGjLc+Sbl8XO1UwjgkgcADsdN/vJ7Ak2tNyNepBD90kTu
WitusoXT7faQEDTsYslRwyBuSXOwQ36Vxsoc/njNUVu2ItrJ9W89+BoOR+UKezMk
rnKPJeiA+8+SNI80IOATzH+fABlJX7ToIhqTX960MHjMXPA4huJ/SWpZ5cvXfMLO
ieF8Es34xJEjyLCFtIztFAg91Jds9GKp1738PNKwrj0L2hHYITPzWFo8cX+98Ie/
14xgilhwDHS8hyVcw1QLoXllFrflcRrN/doUtALj0jTlsDLkYpGFNE7QKToFfXKI
Rjk+ec6vSPVhlpVl/c5DzZLlrNhae4xEmJKR+rlQqDM7OUQp5UFgFHsdEOhhva4R
3vNqtRuCE/qBt3S0YoFMVg==
`protect END_PROTECTED
