`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PLjMAzHUYxKp8DDRka/f14vvaAMAopUK2F1ZxAI8WNuvFkO/++yIrFuBO5ri8bP2
tqN4rCAbCE4qG2vUcGA/cGFgw3U0A4Hw4sF75gsu2/WAheq05YAVJNV7llqzOmtR
V1FfcC3C2XkG5Sp7WjJ0OPYnXeV1NgcBRna2LIyQcc16acpbMkGdw4dmi0CyixUh
Hj408nwyofCWlj6m74PIRlbdB6uUpdOwwCm8N0cqQb0/SzLCUH9TWLMHmnEmSJcS
ci21B4/YIUPG0Sc+1fsVWcHHDZAqD7dVgjEXRzR8ckPmIb8kkjsu/k42rRQId1xl
Qrw0pH5lmG5NnMqG/ECevmXor1o2SGsWCv0PwNSGW73aVcCITdWdtFvxE6L+pV3H
+ITYh/zT0aXdscKFxgr7neBAnVBsOyX8pd739LevzvqmixDz8XX2KbvpSlRhFza9
bLpcoOATlLVzuihHchriGalDeSEtU66weF93B/u78KC/zH6h8vHlD8Luq7UMtF0h
87FGi4EfU+nD8izXSCALxYAqiU1d++h/8XR7WlqjtINUi6F14oePlLGyTW6sng1S
ji/5RC0xNAqmogmL/W9dWG6J4qYSsURw9Bh3FjymAhu/jRDQIecmBEP5sHVVPq+J
mrl9RzIXmmumcylxBo/tASX822FMT7TVS6Zwi41WkuHVE52IT+ShP8/9GupEfNkJ
7T0gfkR5iMTN5z6/c7+9Aw==
`protect END_PROTECTED
