`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oj3/9LfqieWeNrHqQXTeFquTpJ7rUZhHtrvNJiFMxPKxvfKCI3zN34hH54bUdJUV
gtqUd0BKllWi/ZXcTo4eiY8p5vmHWCPbtWnbk2FE4kH7VkROp+FsviWIuZkI6e/k
a5BgBOM83hNpxtY+2uWC7jJWviI0gDbvn5wSs18BNYtQq1fNyjSc/R4o7BMo36Fe
0SWHEUOy37JEFu3exTZEpB/sQ8prpFwy2W53Ovhlm6T4FnBwz1P4XSv9WJjKOWxq
efK4vN0VKb7LeSZsbp7Rc19tNiQebrcUPX/LxMh5NKOxC2RyRfiSLbZnYjT+2sC3
T9CtRQhXIfiOhy/z0QhYdjxb+OrV9hza+LQKFOsMqIGzNd5wW8D6ne8ZJaym+urx
J2aaKXS5RzQtlj3uMD3dew==
`protect END_PROTECTED
