`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iuC6DnAUcP4dbKWcN7BQZr4634GkRsjLJChF6HMVkC7uCJufKNtsOMtQH/nJViAS
N3Pg7NeSfSzyw4R5cNCci/B/Jlxz2vbmzopXmpk6NZErmTX5oihJs6mWGXFbFrEi
OdMmbRtq9LU9EkMySf76PUwtrBZjt6MiSpB/aLan5FGgLGQ1SgCbuq1bJ/0Rfo99
2cy7ejOGr2qD/8mnVEHgIUKgzWGoWucscZhxVHkwBi/aEuUCsEpcuv+n7XUW6iF6
4aktfLzed4h2HvEsMT2lwMLRETnTUt99lxhWfwtOMvwbxjn/Ao04FwG+XuMue/OB
520W+RsWS8C1UbtMa1Bhjf5mbtLpLbUHtlcHNYx5/0gPYdwa+pgGf7Y2W1VTp4TT
vWqXE9WZeiaog1QeRLjyrIMqkqvznMcz4B2wU3/S7g8=
`protect END_PROTECTED
