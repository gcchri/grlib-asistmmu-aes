`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZWXrv4gPJ93FHkDbDGiYd6STpYrvi2Qd99HD5d2i9nskHkEAv34Horp660wTd1NH
1uHpNRGhwvUnaCOHoNGF3j2V6xsCnIq1ad0HNoG1HbbL06au1XsfUWn7e4p+JlFh
KQ98K7xEqahzq2T1/8siwJs5MHsu2gdnyzz7TgQhgS8B+Veu887YhMhUL8KoD0s+
t05QpdiE6ziKw2NgsB+7BHkx3bxGMoctNdWw6zPpPn8zScumgQKUVO9Eu8aAn6TM
cWyLGrrzXVKn02q/Z5pKgLNoJoOXyE2Ba/XWXpLzg5CO3uAx2sDHmm63T+44+md0
YLH++SrTiWCW9vkMezNb/brsv3zlah3UKl7tQziu2iedL6Q/dFAuV5+4OuruR3cu
M9nvZItY1dNFqxu/nSTOuEWtbUqYpy+vcd6/X+8gs9FACMSvW4O0WrRe6EPlYh8S
bofFqRiAZvFYgKbjGNTM9aPrZunntu1tetRcRFhFG6ORq13FvC52+iXx+XMfx7Pn
AUx2zOUehUnF66778LIUd26n/mS+DzVS43o4MA7jiJZzYwbTETGnJ03UDuvqhEUc
bGdWnGRx/0EmYP47Uq87eMesWw7znM51St+/ckTussa0bLzboPRslCp9fHyF0rZ/
oSoWtw8Yua2O80ShBaUvmXi2Wc61T127t54m3i6zxuUj9lzxwIJgQgI4o0+tP3jb
JODONkn8EGmAkiKzL8UocukXQ12JcXuZtNuitK4PXUz3DhK9pkMBCY457k8yznKD
HdwHdvD2MJxuf7dZdUzmQnqq68ZS6BPmT6LEsYeSasfLXhLUm+m1ta006H2NidnL
utsBbmYEl/YJ1hFSCE68liqSnZ1NZq9CIG8LLSAd8vFXwePvyJn7SC6jnwHy93xF
egr8ztRN0jnXUApPNLClrA1I8WZJFf6dZGMiBXTGiAbKThG63DJgfL8AA3dK1fOY
VvkMY4THqn86lDoYJe2NeiJRUJK8UBPfupuu5a01xFil9gfSWOGm1lL0Ja8qPnoa
zdTU3tmJflhq62jc1YEBZb+zm4b9BKa41G9z885gSzmdeNeM8ltSZz8zLSh7921F
LxsCj5NGn+PUbKnfPU709BRv+y5dSILrNNq/4ZqokuLCzb+EyPCqMVuluAUQK8PJ
ucus7P6oDHvYTV5bELBZgGjpzILLSlwHRyMEseyKimDne2DcPrgKXQy+rwKnb9T1
E/DzWhfDM06zvrI7kYJF8pKZQZ2RrYW1zu7oSz3X90UsFIL8jZO9+3f82jQuAS5W
EcvwngnVZPDw0qF3o0Mpm19z3NBLQyx7REyKl7AmRlUU7UNw+o8z9A/YCL2TLNdu
4tifb2hIr3/aWFvk4b95iCMbkj51bDmvqBLj739EcGKNDGxZ0Qwd5XWxA4GQYuus
fMMegm33qHI2Cu17CxrK6MW3zs7PtdL4ybEZAfNPJJudXLcC5vP1RTQAlQilzx4k
lgEY6b3rq/F9uqCo1V9vlidVa0ibji19MRpqs6MPj5SB3pJ2bjuZneuARzv2ToNG
vZeSfkiu4qGOrbe31pXaJaYqqmkyd5ZMrsuSohUDwQON3owavlHlMHtlvy4NyPl+
+cnnZ9IIOW3K0EerffYDJdzzcLAq++aD90T4kubK1I1RInuZz4cdJ7AyCp2y4oQR
GP5h+zjsqqXj3vhR0eFkQ4IdTgiCPZOy7HxRUMf5RGtFlA3enQ6ejb1uc5uTotEr
GihnJMRwltJz5OyfelNEoQV0ygUt02dzWmhKKOtm6YPV40PxgWnvmaP2nUARVgOY
zjk/77VieG9mMZr4+KXdFhSmJk2zrXIgmB/E8ILLyXf52VmGa3tU1d9G0zgSJyma
HsIA+iW7LocSrrV43n3/1xZV9GFoyV9Dxn0qYfdm0Y1fkIZG90PxW5YEEVvY31fr
kheMIw4LbPZtha5rL+6c+OTnkdeqlgK7sdoSwaDjlThnduySIej3viU6hSUBtJ4K
6T0PoUbVtfZ1pDVbzy/3Zx+pH7Ds1BS400eiBsEh08qUZeWNi0ja8TU6gh+up/6s
goi7d8ZAGpAJx+aBbJ9aPLA6TCw88iiivu4xp8++FVNObnogIvJFN23YrM+r/onQ
mczdI8ITVOoh0wrr3fqZv1hezzzq9oPDLTTI30c2mibdiR2sKTkkL1FyFjX+qU7f
KXy9KVV16BPiXvpZH2KHVEI4GzhtL/xlzCM2eRzhV3sjjEG1ydJRceLRujL+yeZa
PTn9Mca2VdRSbPunYfb2kXIpViHmzCSwxgBUIa4gXubK7Y69ZsUQG1HOouvt4wSS
n3DHAwQqGOpq8QRvycwSQT+8RqntMynnmtBgY51YLleoyyUJOyIqtxGgHUnyT6ea
SxwQ0I551DRs7wRQA6eSkzQGoDCWlqDvl98X4c5xew+KupDPATcCYQ8hM8k+f9Tw
Oj336C5sXOYR3sSW9R9LHEQLRxEEgAHGa5oMjCx6Z9m9FvE2E7rU3TomfT8mDTOZ
WDhG4JDo9qa4zuN47+U3UhqwJhjHy33tWNZmTv7zVKtrsmpFkmxboIQl4gO6x6ym
PJoY4mCynLIp97xJQ5iLv9qJvhY/MrHF8Tglyxp6RiK+5toEFBaGNaxLuV+N8bPB
LVYyp9RNfoC2xIRA6CmSnNsFcXmRqm7p0g70SbqDZaGQfhqRqb37KbQTREkio1A7
axiTvbrr+tywrIOR+uG93AiN4aIkDfxA+h6Yk73UrxcZ8ep3MmvU978d3Mpk/BCN
/DQdGnE6OTWvWZlgJa/FMOqlzGlywGvhILKs3a3p4NyIbKHzcujvS9n2Yk2Lf9aZ
8LnGp3ZkS4c5aaOsOdT8gV1I3ZanMAe5YeQsuJ+xs38cNuii290C4s5G6hMRqtJL
K88dI1yLiISIkl5WH5pCNlaOEAI+M6B2nAZ6/82OOlQ0ePz7VdOWfyPMbYRtx59N
ACW3W/4nu8pUxrd+d4NzoNKZkq9lduezlp1kc9Z8drpqjTpFANkyxssF5cOX5hay
SuJ0EcMnlx69uT0BazzDGFnNz9xH1RfmUBki4+/QuALPbcOdx2W+GPz6UVoZWNQ2
dk8PSF0Ah/RWS9MAEFKIu1t5DJ6j8dMMtaDfgM11b0QsN6WO02TS1owuP3TXdRBI
zI2Cj8/wV8t4UO8ChEMGjjFhP+Z3Tm0w1HnblucLn8oVXUNS7Hrh4m2/ttcFuade
sgHsg3/hvV72z4IVJmxjnVWFqr/l8zLxZHbS9MzlF4beIWHHky0McAgkxCR7T4uD
t16xGHORK2I+k8StbLlmdMpc0HLQaEy7AfXlp783R0nZSBSNQ08q8s/2CGUBM127
SuicrVCpVt/fpM0RIr1jQZff9T/SdsxsEDANVLXIHsYP4m4M99Tb90yq7LzovbF+
60kpCg/rFoHuj13Pjt9RKvieuPlFLwZsA9JG38mNuhGmnJ5+Q+EvMgxCMeiPGs3u
bpkwbME4P2F4o8wC1nrboTkGMi+FIkjEBOGTmBCzpBj7n0DPHUvwGn6LsJNo47bI
Pl8so5FUxGek3pdjJRvmplMXB1J6oxyQJZqKRL63zDuhC8NYJ5h0J2oHf8+2Wf/a
kRehCAuep0ddEKUxbFEzB4AscFnZ2dTPyu3kHwD0MDcOjTT9NVe1CHoalMptFvRJ
9gm+3NcLvplFqyeaPBAPgFRgojC3GCJvMwqY+xWAfBrIlKwyBumqgsU5RhFWOo7F
KsyRpj1asDvf/wMZa58h9N/8Q0/EqH36EG1scwBpp83ob5wfcvdslZ4fi+K9HlXT
T4+CAt4VnK+9rGznofZtCFe4fykIJl79WxcQ7DLz9zrZ2KTkYldDCpJwEbLUddU1
RaNPed/pVgRxxOLrhDnKOg3pw5YC00TTv4EKac8VHKIAMXFKa9ovICCrUAp9Ru2w
h4sbLd2YPJc1DPIQAPVAFldMtELZUvQ7HDpUPVvSmm2qugcTVbt+Bsy0/38wpmmq
7qjeOO1ELI7ZjzF0S7C0vkWHQqrSan2BZcVjTwJADS9aH3UTzx4ogBgZevs5blE9
MJreuarbq4oqSZKo1pDC8I5jIYlGF9trzoJfccl0hhYMnR9X9e6TlppFpLyYZgVX
IMXt9uiGftKAPCma1DiBjOXLW6GPqykBdJbdXLfBuMaN0sav6zjqyyq3jiC/AOT8
5lLx9Q8J9iLranhpfH+fvlKQApJ084WNErfYkOvCHuhJ7PHKXKCpntDBF7waEjKP
p85ohSNEVYvDdhyDC4pInwowh6QSFh17+af3f3tqejChlcKKEUmSg4J1En9+jWUE
ZFZac2sCScYNgOJ1WGg61MGLdrWHlV3CQilt018dx40xX+JYvu5AcTelunbEqDtW
i64qJZqU6KI2fKXnU0IaFpBOqPWAd0amnfJOxeKRZRfSXiN1rjoXWFy/n8G1Vj+d
bkrscdRqNzzZX5zLYn+uVkaaOwQrIDOzA6qSVOiuE/WCRknki9XAa9csHkF91McX
FgpKNQgO9LFyaZYTma5IeXFAZnF4tp3iBq1J3xei4oiWF62ptzRULLAY5sc6zzae
o21wyQlZWuX9+YB/1osfCFvPIa0DXuQjillDAMxvEqpnUXuZXvXpTWhOEZXco5Gi
i9k8GJK5XdmEcS1e8lCJLVsz6GzKVE4Ak5dk33hmojU4AHuWEnbYJBJ4Yykp9vGH
ZKo2imsuNfcVnLwdLzpL/BfwpSUa0vYz50127qLH/Y4jFAEFa02NtBPmHihC8nGj
OlT2hYY2M3M43LZIpVqUpV8NNIpPQYt6o0vXpnBQV3FeCPZivkiHSVMvOrrGT6X2
tRbbOoMxozwmEdgM4ylNDvaRwolOfnfUcEqAuuYKgQSeR6npJYKbsv5BPo80gyLy
WvJtV3esjFQ9qv5aReCUB8lSByPjfVLOcNjlTWxuFamfN8Zi47WBNEbRYwPYM9uy
v9fLhjXJ/ap9+oYTWq0cKopyx7ncUavYd8NnBq2Ev0FJ5BAEzh8DDW0JH9XP2pQV
vBd+dl+a0LB26XBnmU8D6FgFlpm8SP7+noYtv2vSYlSRfOKk0jyuigAZLTZQk62L
28MWUGrXrHneMxnc41glsKQSm95mHd7PAaNue5ECZSNmPZaq9lBKCcIVBnZwxObl
fC6vj6hr6Gm30E9fm4FtYu/3c1zNOuqH/6/7YVbW1LevhjvX6Ki2PDCeECInS9QP
+raysF9ltvS3/D+O76GGtuDZit3XN8GZFDocbImJCLp9KZyjKo0WM1rDuKGtFTN9
bVKAF0vCW9obE+FD2AQw3XyOskjgEUxmHr92ZMUh7cRw+sW4oPDcoUQlLB4QF+vU
Ww54y5kUSl73jW/RGbzvTaNX8fG8Zto/laRd5nPYtOAw8Wpa82jw2t/U2ZOIICCb
G3TQ+PDRPJOk955ypOOzFKaAkkda2KNe5eM44AL6wKQvWxhggwyT+J/1Qfsw+8Vw
zwmvP6ApXnnrrrxvAFi8VYF1UtOConY+6c01QOOFTmHdYTOvpSWzxBRihVwTMBqg
0yMv4V2r1oAPWfcs9xzU1DwVUbcICUpoI3hNFz3v0PUxCZRI6L5PyncrVRkfd3lu
Zk+Jps2w0dG9S+jliHo9euJQo2bXe9J5KZSFn3kgfAZHPRv1BmdGdNB8dqsTf8Au
wGKZuEwPjpvet1wnXUEdgVDZjBRO9W2CiS/huX2m5KHkoyFqWpZXjQa6oRYXHj27
lmeMNRDYqGGSgDCvPYFZX5+AI0DBlH/XI7G0zRu8r5iuUnt6I4jGrIFsi1lvVuUF
H2vOun7JAx2Rip9COYNM2bDF32xar2aZUOwzonzYe7WKD5CE3rgJN0osi6dZpJcc
DO6TZOsWL9meJVfoGnTVY84p5MzlHzdqDjDcFySPUinZ+Wf4CIxOpf7kdJ6lahzJ
XnKkgEa+t3bRL9Io73geb07nW0LWJZzw6fSWq/BRQgn9nkUTNRsW0mn+q/Pi78tr
ulWMfSLSLEs0Bwo4EaLhihtDXyiH3m7cgesmCvciQIZhP+mT+XAd7TeFLB3NIMgx
2F3Mmfsl3qvg682slLpz5i0UWu/11cLV8WP9aP18j1zB1iZoCE/sp9eLgunQiMe0
TPioal9QQ4BTHZvrUi6/G21vH0nJH1CJFifLG3pXnsYc5JAWijfUTZ/YjWLxa2pP
oFhiv7jSsiYHHGup5utJISECv7+hHlTOXgyoMaQMhHZowWs8QElqxVOHX1Jsc5z8
a3gArQXtYFL7ouF7n75Gy86ROiJpSm6zWfJ3HtlOh8SygDo3OFWVZY0PKHDkSo6g
ow8nuphDBQoEBs8quVppMXQdlhqAJHpui11LKNN6P63OHjOLjsKIwlRhs+yr3+JK
LJtK0MoxD7qXYXtMro0g/yzIywE+bBfaKnWjvwEYMNT7eiTd02VMLXdD0wAU1FB2
KxyubJoFH6ZYte5SyQZIsfU0+Wsdi1YQQG+eXpLh01G1UJv3UPINaaloQ3qXj295
Zlf7kxpEGjyWQWafD7MNZsoRdEdWxN7FdNurBcmD72Z6x0zRGz+O0UUT+/44Qqxp
pmfcU9zn6iorAx9BM2T87WzLVtRFU8bv04iLI7Dg3doup7k9R75RizXMgzZoWSW6
hkX8nsky2mAe/V+ayb95nJrhPb3UHUU4C++AiA83NdsY1v0DsiRCJMX2UByHqscl
tgYssH+JEw5BWXQ+eZdgBk7DJ5Gmygv4bl0+iDlp0xoEXcNnb/EJS9vnd0AFcpYN
26vrm8xF1Y38otPTumX3V4pfnemSCT6bXQZ0Zxt/EVZNsvt2VO2xs/1IaUmXtF3V
VV0pObC1cwTiRutyM2u9itt8d1+F012s236xCPIDHWaBff8lPS+Z0owBdSd7MkPe
RUHQajG1juUJXK7OPXKaCTvgYWmFnpIOt3ZOWGSz5ZJMIZn9lm6meUfnU3BcO6bu
qZszUMv3HhNeLbE+kF2yghooJ+i8raVDzqSlSKPNAyRy4CP5pDuZlj+YnfUcQUqM
G4zs9/cLVbdypspw4+j57BOr+RyYZzJ2YwAO+qwNMiNqUp8RJ1bTQWQsbfkwsYvu
ES3d/kn+hYc0Dzmj1btiNrMwjjYOVNTtE3oUIrA+YYUBAg7+n4NktSXeYFvJq0/i
npbtnuzwffNNVp5GVIb+UNsQlG969/LeG/0ZBKh1o/pZ3oN73hVdzKc/20p3CeuR
ZeeHZdteILi0WXjPdcv2+NJqcV2BSZv5hlZNrhdBhpz/SSDF9d8RaiOhlR0E2GCC
vyDfxesxgjtMNvOT19XxJDJsMJ9Z2lc5lZsVB+jfxq0T2Wtlen0CVGnyGjl/pu4E
G//0N/N7+FK23YzgtILaP91RBrj9uVj9xvgc90vErBcg02mKBgRIHOiiTVWK+iyl
Hh92jxEFmy885qF1jBXcl2ynXwGrJ3QKeUpAHoZzOcYdNqROybop9OHgxTQzMHOe
dsYfYV8vavRycQH6ZOmQWEWXH/YHmFMYhiKyEFI7p3mH/NaPnqF0gwnb6Zc6BfVo
S0ek2pc5JqQuGXI7SjfSYPxHccBxdSqB9/DaiFPNiHjFzeTBUejjNRKRv/O3wbA+
nNREzGmrQzGaHHTZJXQ8Vi0YgX1Dtvmy3mqrmIniWp3BKbVcvUGXt8D0it5wmS5t
MH+qN7pWlyOD/yxFKiEzu8SI2NKBnn0X3jjdGOO+VEYrO5yboWCIxKW5R96BIUKH
9X7CGw6UmlGhZmUAMMFBGxWaYMcrz3WLdnWoXHV4ftRDduuZ6PfDHTJbcLMkYRiv
sRjpn12BhAnWr9PFTlRb+loVHHZ+mPFk5SahLi2FWKR4P/dSmVubhr+lJ2jlBJ9H
LMqOfVlPukO3vKoy0T3UemSPdBV6NEfLF4mzf5ELt1O8d/kg42hV8sT9Y2mVguI5
NsUxIGTzOMSop4u69Ev3CA+6hagwiXVAAg+xBMChfUxOuJCsHM20IyLJ+u1ezwXo
aGG1gQMhlWtZoVCQaFpdbWmQPgZYc22lcffgafxpsUFJFVrpcuyvwbUC/UqtAfr2
tq03HrJqBs19qBN1iB7d1o8aAnS5blili2FcN7RGb4DrC3SyDIfL/7UK2/yHalwI
hLozOmuO4fJvQy9trZ6sni+xkuyog2b8NRd2kDmgeQsSyLK6yy+r91VBMD35iXoy
HF1mBbVFI7Za/uFOByNoKdYo/YRr+tRXU1bpdrJ3fN6yR+f1mI4Twk595nWTH9J8
hqq+xzzCH/1dQH83PegFqa8zaiMWrc71cgBlgLWFUSFCzQBE83UoiBIDHZYhTgFC
GiDSifPpiV+L9vVGQTAkwQmXjZTLHuH5Z7moEYvM2CDd1xYPQMYLoJufRKqvaOdE
EXou2SsKTB4W97nuvamU4kqaH/xheWA4wpzTq2h67UkSNLY+MKb2v9n0Rkc7YL2O
f0idBzoPednsbINz9teM5+RL2hYPhgXjioYVcm+hErZmibHBdyu1r+d14oR9eqg5
golQ4W+aRJFVrbfsBWvgJd0PEbIfL/hIZWH33iakXA3gTdgA5KhW5gobyNfqrVOz
yzvAC86bMuIAp+ow0fEmb6kOh2iDdX/i++arOXXZIw4Cgiwyk65yYP3oj/GNOjd+
Ljej3lYayLD9/mJpVfT7zLKUXhzte+MvWlo/CEtmsWPBloJsRr7h7co2mXLhF/oG
+DJh1FCX2oF/ok2/KibY8bn8qdXYanfFuqBa6mfsnIem/1+zVqVanhF6e+gaPClc
gZhHtcSeZv9fe+Xn7H80OQAXoOqFrBcjxXBQWIZ4bXpbSIioyi0hcdNXF3VX9JSA
gL3mTBmVKqgVIjUi+2Ws+9YLw7mXzJWULUBmSlcJtTeWVdhfzfh+uAr7ZyYSUNOF
dL6AN2kKvfBif23kj1BFpoDp9cbIjX+A0iZFdqymnpggpT70GPA+0Fw/5s9Dp5FB
+4tC7h14KdiFk7ydZz2XYGOOGMjUivYPVFoTyIR9Li2vfP6QBYxX9eoqBF4C6szv
RuJar2+nHakO4RyHX6NIL9cllQoUuFnX/VqjpJrIybui0zAifG3Kb23c14y7Ktc9
DFQ0NqtC/IGMi43I6A6k5yvZYPKL34D9i/blq09BgZBuM5gjIsJHCGh8KQw6TnvV
vxOXfV6F/z1SCeOulABEheo5UwK2++GccMihcJnLZM2NmY23QRz5svKsB5bAkLq+
I8Iq2qnBw14pSdcTDw685dXRCx9c4msIuqyT7OS2Yr3eFrzl1j430nIjzmmq5dji
3i9s2AEeESH7qbJIRW2xHLATu5GU00Pjn+80LyFAuMdB/zZuOlsi7bPLERtFZ29k
lSWyY2kFL2/siAVwiZZleCVJuPpkrvVEKvCbuVuLtIt27ZA8+a6MQbInqnmVXcHk
LwmgxSKwWU3PrS6lttK/pA9qiaPEU0nYRfQxfUy5McuroOqb96lXkkcXWY1cisIz
OWs0/19QRmPWj3gWoi9GMTkMVpv+yeLFRqiu0PtaGNmcszkg/9ZjUcyu1IJkVcp5
WXoYPPO6V+2zl6XF+cc5MG36DM3ndkAHyR8I69Mlh44sXj+Kw12HsPx2XBuIoLjp
Qb3j3PtCUdty3YWsf+xLmy2v+6rVVUqewsEIpqhUwLUKFuCEYbthJR9bMqnI9R/O
OCoLm+yzheBt6CUv4QT5CC1Yf5fJjB44CibSSTnDowcFI5kbFgS0dtY7libY7WOx
wSw76DGTVnDuK42PzEp7iknFyyvR/2ybqdXxLFodQ3C4xS8dhxmHjBEFTnWpDqLo
dd9IXgV2o4BJWjwSfCT7F/s6irbTeJMJbBqtZ30kQ7Jct5pRUg61pKj59TEVzRFx
kgsX3UiSOFcos0WD49axhgLfLdGWT6r62hj682r7z+W6OJOUfgFSelDY+L4Leeec
hFlu/oeNKLXgUiMKw5CV/fCMV+g+ln/rSeOCuYvtixJHGRa0tn8FTlwa/TZ6aHPU
wkRq8uB6qC6UTHmyEpW0crLUiO4tmwddP83Vq69igzjdntqNiZwRk4+imuT1zjiN
FOtNeXiNz/+wBa8eJJG//lQtsQnj+keKcQg4LVL41gVoeKb0Vca4/gPmtKcuKUu4
9d9QeoJsLyeh8WELhnYq+RPUUEnm9m5n0nZCxCifrk1A4k3hf2Qskoc0Fac8KDd3
pOo+aotuied9uvrG9YODiQO6HsJlGgwKLaZiW2383D3WdbiddZiAg/qBRNVbSmDo
/YMWRo/We1mOWrHQjdamWUZLjXsjHeOYUndmDXEHKgbkvHslOWsY9SfkZELhoRS5
3/88ms8U+d8h921rTkEGqSZBmuXYXYfqHGSgyTXwXEPxuoFlAYQs5xcCGYklUcXa
isDSaYvDJ3HZSOpa8KOQnUemreznd0Jm9d3cVdF3s7qk0M+/jkDGleEqFKtw2phG
96nX0e9NIS8jpGoPd6yIF+4I/VwoRgKWerVDtIFkJV6RaZRx7HFbKzU39vLYdTmF
FjZZGPNHK9IZcR1WUGRQ80md4MT+icUMaUsJ5xJhYJfz4dZ0OYdd0o7Mrma8OhPa
oGR38pQpa18voGgtppQm6WMA6F1AxDADHi0EfPYXQelz6r5gpsLgbH1Xfkl9kAjK
glMEuWu68uajbcSvx6N/02DEiPZvgNg0SoTmDSkPPl3vlybCwvjsFrgQO/6H7SYS
SgYf+4A996DeCigMwd+sc4ErYX6VwC2JmXkghAuNEzI2U1/5HYJpbq9AkKaNtg5v
63//458wI9WOKTvfyk1vsgqn0PGpg329dufQlgVLsMZx1FOYvJdwNE/1GqH6pW/V
nhbl6bMDZ3Ihu2iX36D906CugWXwip9bn4GK5H8DNNxGpcs4+ZKqHP7dIbX/v5Tf
d4kzKL46B4Alv872VAOQlau9l2uQnlYiRH0XAPDDnbiB0WnQP2nVa352ddq6VfiU
JxofiIktatkoppaoRbngFoHAQ0ewee2O76neHXXowE0gxHXTx1y6oEkVTERC5bGI
2/BSo5gQELOEe+XOPiFDgud/NAfeMa3kzVn9pMpn3/RBScgalG+ICT8OiGwWH/PA
3GF9zkC9VF0TbW4WRgW2UnlnB8/03YEre2cTl52rEDshUpWVpjHweDMXYiG5OTsG
W2s3BDfXHBtW4EBm3lQdRjOOOy46xReruNUGU1XMzQ6MmQfRBCSkxSwQjB4jn1Vx
gX4uUzzeIvMSVpuZ8g/6Hb6+zsAsLLMmJirgQocCSGY6DJjM9RM/vTwfpSb3KIqF
5f0ItMeEptJOY2Khfms6yGDywDiNgv13UT7y/nGmFNxJ803e3WXC0NSSDA9DzsTo
wVvdrIspyPfroyXMmRErw9Ss2vNA+p2C5zZrz+wEYaJF8WWnIzEtZDny7VKwSgFJ
5AELXVHhOwQJe+bxEUkXne3tneziWvPgnYZUMX1ESKPJkoLLCRfqf+1wz9RL8mib
1HICyHv3f0w+2KHS4T7g3RiFJZsLNW6z7Wf3WD2mMCeDKM4J14Qe+87BHbdpxw+x
E7SyvHziLKLcJJC/6gXVEny2Fp2N4PmTTgvYvxr8mv929Gl3ClbZ2Dl6k0Jh3dfn
qxU1l5auOQz0i3i99Qtpr7v/2+J+pY9qG2QHsF/FvyqCHiRBwegu4I0O0gSgN2xw
6EUTbQ05ctKh21WkqB5A6F7qypKwB8a/HWea8kn500F7y8+xtC1HIFnDOAQYlxeP
51VHPtH67QdA9tiYRzNYyHXtJmxmH/d/OwfstMqbq+PB7mgKg5erDhUTqX8EgzGV
+oo2zHxCcZw0zURuy2sdOKGca2XP7lWuQShTvrozEMxD+xsXWUK3e76VwhFmpMlR
ZXEkZK3VwsQ7XHPS+HRfCqJXGjGs1RerexoVLMatbGRbRKaJtIdCvtiITS0ZDmq0
rs2PncA0dNrYfE33EsJelnPrLrXc4sGfnEIO4y8fEWWmMtg2sqmKarddg5+V7WWT
QmJ4TSSXv0KjBQguja4OwqASqVGKyNQxXWYfRMUsqvt+pDXAcMWy5uOKBeGAmwp+
Irov9zvCCRlIvPxRltuyndbocYD75U24Jx7VHzLZdF3aZokBwPpkJpSly4lOJE9S
DgqCyQQG7XXl/JKf8TtSNo7Ydt1OS90Afa1f77j+GRD4lXRuEbpV8KXwbjzEY4dO
sairMMhCG6VH0i15V4MKNXnJQS5aZasJjq9UAqtATy8yy8UukcJYG3Mg1n0noUHT
Yoj5lCKEoMW8r6cG+OpokejKH/y3Twm+CGxc9tSJNMVaTeWld+UmgrrkRCnR+Oij
3u6csC3X6hcgV0lnziPXvPy3Ltv5ZYQ2yHfTV++irDdbhvBsn87B1W1rWbEI48w2
SRIQxKrETz+9wZbGx3FUNVbx3xXR4BoUgxtdMfDDPwUflg+NkHFOPjsyJNj6A4z1
HuuXauqdCa+yz/sVK6NrPVmeFxG2QTMZGpWRoutotLdFi3LAiUu19X7wsfJ76U28
97Q0AihsguGOdB49k9CpVPSD49gydOYDubepJsx+0xADxt1z4GbLp6bUtjx+N6ST
l5QZIzicYgHTLXmF1B1N2Sq7B++Zjzz3ZG1zK2mJznlHHz7ASlS1nqSc4hU2DxT/
+hWZ5Fyap44E7rqJmK0XcJtVP04fcpQNX+YLXZAncMPz0UqEyUpU7IenuRaMufdq
cPh6nq9naeBcXMSinepyBkRfxh04fstt+dcxd+USw2a773uMBwdXW3AzVCc0Du5k
xxSqShgPx16Ha9lJctTU1TGR/q46w5p+aYLgeTdFHSP3LQ5MjOWDTs6wmgWU4UH/
qdjc+ZHBuGK397PnI+z93yRU148Id+ZvOWekVuqHfv4tuqg7LecLqmYBgJIKXCQi
HOSOu0L0l480X5EHyniyqELiMYkMNYi0CJlnKR1JNL0rVdVqZ1oLj50Etnzo2lPD
1hltkA1U3xMt4rrsOQ4NYPaCYZ081iYQGFcQFwuHZsy/2wZ0Xy/4lBcuppsH0wgX
te74WT7zaVqdDyVrXSU4J+yIycIa6D5+vk8lkLw6OIvv8ECqg7KHsFKOhHDS9eBV
NuS+NE0kiynr5aHJI3zuCXG79NepQEIAIWjmrx6jxUDc5ZLLpjsbB/ooOlWjLfM/
YBlQ1RxekPssRAZUNxXqFJZK+m2I1Nexe9eqneRNwFHsVrh+QDGLH//D1GDhe7rK
pkbzAKLPWm+iLhz40YJl4DWcMG1Y+HnUDe9w3H0jMEyH2TD7TCROQE+bkau+BLHe
PdBuv4kkqKI6VuqPwcz6xXzuShv4oMKEj/ndx63f0onY4SpGc2wVVRAdm5RnbNnb
iQ0uQE3doUngBsTlhStUEKBTkX2ODVx6usmRgEanYcSxGZ1gcHXeJnGidlX2CV9A
mdsCc0DEDyxoYD9YMBWLBc7jcvf0azoA6h1GmuWGQTEBs3Q/w4UvxZ/jYTsiyLQG
sUxkvXn92XluwCly06nnz7CUiBgQrf8wa4M0K6BAojUSLaAKPWTZ173g7UaWD6Y9
opuCnTvs4XpE39cNIgQ+BgThPHhqV1vwjJe7ZjgzJ2V561S5LlU5JRn2hFciNNfY
/Bu+QiBZRUzMi7N5qJnqdpU31gMc3+pv5WxyUmJRtOI6EbmC7gl8HQGZnb0t+7Mq
Z8qduheYPhPb6YFcC55leyospHaiwaUqI8mfxMgXPqJ2iV/BnfnXkAn+daUjjFCA
CTzTzwXs4ukuzrffS8YHupqCxrSVajJhBRpdPo4kn3toDsxUWjZsvb9VdkyanZS3
EeYug0GC6HQWA+Ktiw0rQtGPJyIXXfZS1L7Zf9WmrqZFckmna7aWHfbn+w58WVNn
wbkOrmKmvfHqVngi8THPDsxaZWpcX8tmaD5d+x+J697rkmQqoKCMxy+0F9Mj52hc
TGp4+tUcpMgcUktqEkyC5sZW7L7hIzhXP6mNUnQchaouHA3CJ5C5s9l2zfDfUS2S
WZsxa7mpyvVfyx2yIxQwmH7dJV9Kq2ZEpFotBBEXc5fSW9tpsylsi491YhEZxzJp
wHcV9iVEg79Eijdf7YHYhf7/RgO6y8qu5XPpy58oHbW8a78Zekrq1kPbhL3Qr+Ds
lAVqo2ufhTZcMC9ZlLyzLJkhQGWQRSH9+hl/jODbx06BDbNYhNzw8VRnmTgItENp
pmy/+HyHqKW6nlrGHl/NXfEsASMvfVRs5g3f4kAQiy7JIVO3mpQw0097hVxsLQ6i
szmfJe8DG/PTeEb2lQxhbjeZJsGXdj4ciL2wXScROS6nZpMWnbPQf5ZlgA9ShSVf
LYFq7t5Kr+GuyMYdRhmgpP5ydjzHvrp+LGfOKyOTQu3/l2HM8ncuDzRrlxs2PFZ4
V7lZjq4XmJzuGFdzzOZJQBRCc/toIn7oh5o24hOu6fS13EA3GCffKhOLuMzfB7eX
BvWcZGSNq8eLbHXsMnMWNAUG6RexUVBpGq3kbyJH7keUohQnFE7uCDri7YyzvkLr
GdbLj3OFIdfzUDR60JndnCUKn9vz41oRTh5QGHMfIRg3gVQfMaaRVQvqt1pPITqw
KQXLOQ5nwBEpxfi4D6SHMeBqtmpKBbWLaLMZZgvHxpvPYgCviIGibVkhrWa6FBc6
5n+0+NhhRDpaUGJMvLSn6k2g4BCfLQNEuiw4FvnSDgqnTnSI2GgKgD0O8UEQiuuz
uZrtSKb8AbamncXJf5G9YOWpglFPqxtuWBWGdiYI2J4Rd9E9SFrL9eJHjZveMssZ
FgvfgIX+6+YJosaxeF7bQTp4HVlfD1Rr941uN8aTsdG2xh88XcoM0LHpmOu/RUEj
sY/diX+Ca6HSqV/NfXXjMHTAQJTB1nwV30mnTbw/HuxEljNsckuAraHmajAWTFNp
bb8SSxKwg0rYqVnuMgFQji4L0V9E3uUz3J3XV6FsZU3qPX0C0Lhi6uJh+nBUkJaE
GpaJIEmQTv1269Vr0A8rKfQHf0XNNsntk1eT3TjKt3SofJxlcmrPKGgokIzMzMOb
IKSHmFKExKotGEOFOXV0RxctkIqqDktef7A6oj1+6Zre1muGz59DCZV+yujvDxHK
cPsUrLwgF7QzUbkHMpvnqGW34lB7Vwh3Del7nzVi4gLibTOZtnoAmMWL6KiNWdH2
/xqngBF23lbgRRreDQOHGNRsBcxJNjrvSvJp3y2QSJVPxUMVHV3CQO4dd6KqM7Rt
zJvGOff+YgiXiy9bbklDfY5TDIJBYG/XIpGW7hlr+Y3c7aPltk1C7tU3S3ZIIOtu
boRhhAboszlUna9hfDcfcv8XHd2BzBQ6fcHJGVpkVe4IA4rKB6s8SJCrisM10W1i
bsPURtyoCa4HzVzr9gZjVxJ9LwQYUi/S3gotAVa+W+xPRTAzo5PtesSi7ttZPM81
0ZPjwh6Z1QQx8yw2rMOZ0HMqwhCQy8nXuWzxaA1WXLFMSZUSXSU0WjPoNd0rDxLw
ZnIdKGcC/LB1d4/llS742KLI8U9PFlL/4nNsFwzGic8WOXIeCc2H2AVyInpoiVDi
a6+7ianOZ27BKCFxtwF+AOEo+dlV3wyMBvdl8BrTPZwOyw1bbzPgQWjWe4VA4moH
sQbZtPvvmKptBM3qAyv9FPPurwgeOuUrzp44/S6IZejN+enkTo16iBW3GKk+p418
9O0KjY5OS174lGVnsx/lND5GU0hpy/QZovu8piEQhVrk3Biw0VZhv29Ce8xz6dNK
KJRhNJPFJlp0DUhGPTSdEupFYo0kO+YElpih2sJZIPbChORr0BcMOGT0wleLckyy
eGDYfM9wRaySa3n9+dDRsr/0wwau1e8k0/HyykkULWea/MAzFAKDaz497dNiqNUU
TxzDPWMuTgikwEd6vBfTZqgXyWuucSPMkE1CGA96WED1h453RTUfZHvLzVpAdYe5
GNMkLGhU/rBKQguAepmJeCWzyf7ue2PbI9D2OvHTgGAAAbQC6iL7eA8rDQ7g1WOp
hEDlZ6Bu0GazKXPoGgi2lh8+7LkFBNPChXbcJ01aowHZRg8XIb3T6FGBCL2EU8Er
/eM3XVMvPn/B1/VlpJ8rMEY8gCyGImqCrfs+q28Db62jNWWNwENjZ4nOmZErzLFT
n1YqRQTdJn3DL3tBPzGR628W7XBha2UEok2OekrN0cyxY7g78ex+H5kBllONQbbW
y++/WTO0f3xrixI3bx4358wB03OlqfjQgPxLbv3gcOJY6O+w3ZuXZvWMglWnoSkr
oIkwkkxDG59hfcCyM3jvGCrqYG0a9ARoKGoZCBnJVp/ozcMUORn3DBhtlHQ81eQ0
cb8uutcnam/qOnIhym1K3EQY08557DPhpxYFX+M+JCh1xHNzMZEcRfh+NBJCmpSX
lS4mloMhI2uqC4JpzKQfWiSM+45rLwAzR3MGtDqgjjy1Jx9sqLj2s/HEJenQLg6z
mItt2yvolkfn+99fHx/GzbRUxgYtJWh5MqQdIj/rrb2S4Vfs4BNe1z9/mDgisLvA
NGZwE6dnbrymLkF4DupvzIuAn2r7/yjA30v+FJXfh+kQs4PVtokVETrf+d+ZNUtH
ZI6/Th3WDDhH7iN4XRX4KoAYsbnlzNkngXEhwW9VL/wfMa/y08Ym3JaDJaFBBe8s
IM1s4vMItIZhSoOHj69HhTWMjHCDK4AIVzEN/vGAUvddP4JHPKnMdJvz3J9y/04G
U1JTwjk6ds+YydAsjs0enEP3/mIFN9GHIG8IN1WgcW33/ZiatLEM4fLOe8RLip4Z
lrIErLdut66risB0cxJRoO/Vft1dXBjWD5wEyH9bBlL84x/C5IsxVN9cruGkPpiB
yLBfLn3U33xf1nSqDCEMOdp/HTidVdoQXq0v1xKtkncut6w/QEI+Yfwsg4kuSZxT
aDU0HobLgInIrz67ZpqtcGNyYPvnqjJpl8VEld0vdDtZ7O3yhe+N0/NIsiFXpOiD
zDh33/th8cIEpf7NZO77DSUKDKY2xxA0ZmaJ98XCJV95vwXml85QltNSsStjt4B9
uorJOFiuTaUVpJpbAnrhctuYh4kXCgxofzvXnd64sjNd8ONnEcNI0i2OvOOZyyCV
KCYvWo4uZ1+xLhQcc1FaXC8IDHn0Ud1ovx3+QfB5YcMmb5fORISw930EHwvw36ed
8/XKxKruiKAbfgV8aiK3Zp2lOn8qqExrQtgWrWfXk5k9CtYFr3/ENlf/yNQ+azKL
ZEUYM25lNApVS3hPgxfOB1OTQOE1lbjjG735Jsoa+hBQNInV1Y/qCautnI5fmcNi
j42DS3AMMjIqDI8wt+voNfJtea497bHW3j4jZcYo1ZxZQExgYW0fiCQQkOcMQl2Y
VgaXcD5/kxnFEhKHRNTm4yBxWS1Isy1xVECp+ihp2gucYpNBJkZS/47thoCEAWRg
bLTetVCrJa3dEu1H4cWhBofNjBSw+fN+yVf6TQWUulM5+0rOYOXnNi4KunVBHPrG
4Xz2G0IiZmsi6m4OXc26FIb9hUQmB9L5zOEl0DkHvaeGIc9D0nOIaX+/IShd4fBR
RDmozAZI02kHwLlx8H3C6Q+mEO24d9zhaVowQWYiiHEoFIOl17o5cLxK0hgq9jDr
8n9IfWQjQ+68+Vk7LkWN7Je6Bqgo7r0sBo9sWQ2xOsB6Q5tZaQOAKJ6nfdG+vSKa
UdeGJ0XqvVlNRrxpa7amKNKSYE2aA+7FJd+eEY6YcA+VcN2Q1Xl7rT+wMD/wpsgg
RpYAFFywvBLzWn1fQ3Xo+nnWHTgScZGomsxT6x7da1s/mtE5WJuSx5bCXSfbHW+g
9wEPzINcyLHUYr0yOQcNxdvakAsx0FNwIkdGYZg79EHA3OjAU2P1PqXkry+OLB21
ls6bSoEodW3axeTDQHuUGuVUCedJVfVvY8h6fEly6lZh2cp70z1XPRJ794CUu+NU
bS7KwewGMhpHDHHkaZSBczpOjtkhG/gcNDkvK/l94wMBktgiT4KZS0FUw/E6zFgq
sWXmwZXMwgGVVoDyzGkbtAUh2q0MsDMkeslcSvhRMgPmEg8hpfULPAufrgY5iO34
XPkg+Ih9fIoBb+akUQB5UyGgvM2u5MeOy5NkR06iBraiKssAAZsrbnWTQdmvjWkN
CWWjN2zux12aqPUEJhnlW1hB9vus+cFd4C1G3Wug+v0gOL7tqEEG3KgQgIlRrPNX
OA8sMvTQayL4YG8lTIIl/jYD8Hl5BDnHr/SU2SVqnqsKNmX6roj2yfX8BQk/NAp0
cMEGgZBVpJdPzPhEGbOUjv5rRYu9ouYSKomOmQJesBFd0iK60bvQeOLLzrSeHlh4
M7mOaCX6TjcAzzvbTM8QdtQmrx2TAnvYL64/UY94qFu6aDBrWZ+YdTi+AVD8Vgpn
sqhGto/FBej7O+kWZLzqkCiZegB7/cbDw41fWy6tL6MRjRacFwQXrPjDPhFosJrv
LarJOqGE5wZi6VJMO//gwzHEsDwgkhjRI17muz4EEERzcigHauZ3FlmDXikwq9Ry
P5zwfuA6MDE6380vlbreXkA+Q2cDe6H+gUC+aH3GAY8Y9LR/AP3LZtbZ8FT6VGNK
PtmnB/PGSKV8e+M2W5avEUeTLNoeeVB7Qb1o4NPfr3Z5i3bQka2gP5JrtjH6h/s6
95lpxjXGl8gRkn7ranscrbflcOij51QhH2mH5m2KTZRRtRSD5r7HElfJkM/hl54I
2Lsy8CD0c98NrTsRUwks0pC4/5mvnit2FIdSvtEb0PMWY82/v2mG/fYVBqZXXPLk
BonfZ6CSqXEOtFhOXb5PnlVYP8crC1GIjCV8IK4fClH+mDBmfMM+X6qL/oydr7Ck
sV60F9FGAei3nb4fRov2fGGbk2j62ozat3V2pZh+CUY7lEqOV9BXOG0EoJg5gVgh
VKD2LmVvBAdUyAwSugfprH8pyJJ/okTlOXFTj1x0E3H6BZuwGp0JNmfiwI8pOqgv
vI5xF2kcB8mPjQYj1GoXpDKSGSxjpgINlz/SlUlcXEKU+tJyTaP2Jm+SU9OlTcpc
iH7Zdcku8hXGZKcR5xcuRmoK3XwirwIRTSvT+9+E63t5CaY6JJPtXRA9+MywxYT+
Lm/emfr6T6HYmBeQPi7EUlAWelqhrxYfpWFaE/BXyj1SU4IJFvvsvRu5X2k5q+2P
0iq6ihZOPkgKKNR6omUZ2VA4HPTzFPItfy8g08d/wkSsslZo59yXPhmK+u0XYfx1
RlemyaKa3lfRL4Zuyx7DxBQ6f79WiJJgYEjhFZqLdwfYFqlur5/pRGKhe19tO0tO
pkmrHlUtU+DrSdV29LyXVMRK5HuKfczwfn88azukJ51Gx+Sf21foFICS+7c/UCPU
DLHDraA0qv8JMgB70mOay0Vy9A4z2GOFxQPa98KkeKRfWnpkoyk07qTSiwo1/VFg
m/DCHiuWwH59NjpB3kv2CiBRbqOaazDBsTbOw/Um7KwfhXS3NFs/HeX/Y/XUJNeh
UC/gwsemwF4VxC6lWjei+NPGBC3VcQpolXOhquJ/q0WCQzdpeZk2DUyoAN7RH2l1
pTMg4TfRgKg7vMAV5SFFyUXOPCl0bFVfAuvgPbtyHIOf3Dqcw+OdKNQTnoiT03wl
amtxyK8XAfKiDaarzeaXY8PrtU2HKZra86IpyaDSJNQ2Ub0hgUnIomaVmHv5H1xK
ONqgOWNNK4PHhSPyNkpxtOWpmw8ukeTi5pwM6XzxFssXJUDdzdPdkRAFr7GFMyGD
rJ6ojaRGakN2g/MrKvlrlJesvdtqr/MK2q7d7cp0JgYtjc4w1rD3XofgTHBvyJqo
ff6C4JJIBsUjlsN3A8onsJ/CNsyaK3PqVdu4Jseo/zFC0wz6Kor3Msq7+s+YiSBB
VxQSREZgw/b5f3ZWTCw9kkwOKqCgdaTK3q3U4fikCyGgq8Dv3tJcOTfIbZLZR54+
T9h6uUQyEcRRBc4dG1PwJTQuXlno8z/aABZBLvej9wKbmCRzC985LNeIeeNMPpdt
t7vQoaEbtKfvUdKPuTeSUw235lc1tYidspMvmlEj4+7DmhSLm2a926RFA+64Fjo4
BqJ8vhrN1Z4nCq1ggmhPkKTQRWpkz0Hu9ifY+CIHUVtvRjicIvfCKoTlNiGj38j/
3x/2ZrZFCKA8dHOA9qCHhtG71hLmDZqJHKdrzd5wJGf9+xDwBTsIrhXFDk1dviJV
4Rq5YAWIYYGJsG5KGFjX3i/koAKZv5K/4AaC1ldtIaxi8l8QHziOaWVbd399jG/d
VKD4e68nQ4NCUa14MWdOigK8mvSz6g/rEL+oHpN38JFioZWbvnFucyl8yTIBYbie
9mTqFZ4bO1PJsAAIQ6/+SSZFKCrLHXkwzyhTPxiHCQEEobVS7yY2lnx7X8m1eBd7
n9QFxy3t4KSTELSTW5daRrLrEu3Q618n57tCO0jnYf7ndYiHTXcV6W46CnL1S/J0
g89QtSGjOhbrk8JtI4ddahfpzTeEH27M/dkarAxuoQyGHyIEanPNSKrL0G7LlHS0
17JL4ieq+H4sC3w9mxwEzdrs3NmU7zHeUAv5c1ST0cX4YmHhmUZB20hvr1d9bckQ
KtT2VCj74ixAJh6Zx9mSA0mj6X4TTNG4yqhYFCRskskEmZzp6Q/Fk1TWSVWyRIif
oXtUXFk+MAQ18IeXhW64wxGWb7MSynT31gEf/kJ1pPC15sPVGCxnoTa/kGcfa/um
fFwXTv9yEqqvx3Py16YZF+sGpIrZ99USe0JnAP9cg5uKLzDGPTSSgr33E+Qtt9Hi
wqkMfOW0KRxHu5rs5Ju5vZwwkC9/Gt0PRO92lc066No//FJJ1iKNPftaZ8z1CjuB
o3qKnt178y9Vy8uTpa6O7291iKw5dtrm+54cWEkwKquycQSn9ZuEYzLkxN8kFF1C
1JTXOPZ9nPM8AHfU+hyXokmwxPeACnpTYQuOSfU/DOWvKaU3Pdp8KMPxsOyIXukR
4PgW3hcQQmG6fENY/p5vEEbzTBXRaj0kzZTofiCWU5QGrpijauQjnHftXTEzU+mz
vB7V0TBHs1Nx6XGCsYQupKrsbMdlonUZ04No5RNRpByiJYoWOg5KhsbNinJb3eBL
V7g7D0ssE0bKvmVH/UondTOU+xqS1vYcbbyz3gvNYCVbk0KH+ZC0kyioMMjCtQqg
NUulFHKCAZLMpY/CrMjmzOeSxzyaOMPeyd7okK73QVXSuEnpbBE37GRflYdDEWak
SF0K7wi4v+lHAog9bw9knRJ28+1JU5aV5F9uRpcwcnpCypGhZVtejQs9Z7uyYvvs
80G3vYIT1nmUrj07Dvm/B+51/zWRF6/FjNJuvkVSLcFt9gsPgva6Xw+09VBBubB4
en93r4mh0GVks1OZUW6oScKkq7s66a7IG9vJnkAdszvi+dxIuikw6+sy8UBVK6+q
3WNETn5FPUnAy7IaLncc13oMjvgwolj/zl1PviBOFurgxd8O3SYbRQA7Iian1ZVD
cNxSlSkvadB80E5NTDOCDz8RJP0i4SPeqJcIzsw/JEYS2AqB0bIxRjCkxV0Mm2wQ
IS4rofwvrMAMl67BxGSccOZt7PHNvJYbXGiCL4UzcQqhz7PZxpEzAL+e3eCh9nd2
7fW6obA+P0CbF25HgxFAjz8UFYGyfAfpoJRNzipZ1fmKsvsqx7gYiANRMBGOfn9Z
e5GiKPnNdm571ejkHwa3RvNWvK8rBIGkgq9TIHzcBPgiZikAjz1e9dPTFBmjtUtu
c9mOilYHddfF3PW9Dv7iUu+4+TYjIkIu+Dw2ZiB6NlkcSFmTs1Iq/nlMcDdRiGFW
rW6PJkwZqRYKvdneA7u+gIh7baWhx+MLNA+OJ/FHVLewJe0e3JjNvHSXiEZwgnvs
Ye1YQBrJ2TqB31lVWygisi9A/IJY83x2e2h4Ub75Twi9iWao6k+ErhHERbOg0IBE
apD+W70WSkPadzDMyMNJsp4ec+/FDVUJ8pacS7CCdoOBVkzdkaKfK42CUfyrRQFB
zsWZWzi2md8U/54gwf8j3SBlGnQE4MKXUPATXrPvnAAJicje7iHrAJSa/O3FT15W
bVCtGSHdWem2oBodm5mWr0gYcBU+/gesj955CI04keqHHdrE8FHenHFMZocOMgw3
LyMRlNm8mGzqz1u7AJ3jwJj/7zXYu2AbJMRZ5pzlvKAQGo7oUd8u3wgZ3IkWz+d+
50wmHCDUzYwaOKTwSqJJiMZK4woFaaxEqLiZLpYubqRlM/B/Tkg0eksXWAg2OZps
EYX2BU4cQQu6W4aI/2zN+3TDh2AUwaZIxuulWarqUbBUU023RwXQSVvQXjeqHDf6
qPMdNBEUN0c/rWqUa7BjykDjTHOg7IAOHZ/uhnK0cx5dZEiuAc9X/SVdKo1j5WX9
glKoz4ATtVWBNmfoVHtBelLIMO9QPmFp4SHsScgG8nUYVgATyArM8iZdWQCDyznF
/leuzzCyNsTBsTV7pZPNgmY8XnYvZVgsiTDUu8mOh7WT94sevAwF9ti1uLyjTI3r
mL7YpavUJ4I4vcwmYmVbW16RGph2FTWkun9poVdNkybLaoF0113j/2hnqcqLCnys
AnTSvE6iU1PJEsMbARlTYtHRGXJF8OgZ8e/QPR2qt2aY4uo2HP32KBQQMxoHwIzY
BY1ZJBDQ8wUgV1k5H4hATUpDgIKQ5SrFv7QV+Uzh4VuLFRhx7lRyZKEIAAG+rSxA
Yr9GNELe9C4/X8y+cExlARaZ8Np+mACnXZ1yzlpum4SqsYtKJdivio1GMK4ouNpP
n7h7D1dQmsZH1CJDBKmd3WxZ0KYpcRBwOEl57M8n1FzpDqeSQ6yCzT7+IB2fglnB
Rsfizl7ejFB/xa6+2jZPsXwq/+rtqQEvrN2/r92GpNXItpZJCUAijKcmmK9DXiOo
5MF4ffhn/PB03j/VDDCNayyfn94xhX/wBYnunwvhM8T0aTuSBHnCkaqPSh0nySJE
uyn+4YCT3kloAcbSvjfZC+bxQbZA85m3wHFX7nWNqE7X51hNEHObV2MqS9rG08wc
RoBXtHabCXmnFCV0L5Hh0OsDcjtwQQcEmSZvL4iSd5ygOgfN+o75p+F+uuGhBa8t
Tv/C+aPf2bXAWBgOyfPQsBLnodGwEIzI4DQ0oJWFV3aCpz0sXwtu9FIPsUkB3lrp
6TvJnwKz/Rpb9SNM2iW4c4fzS3pU/oOEnlhR26egHGWG0dikvLTSjLYBryS62plG
bH/Udi7UdAG06PgUZLBBI1afIMak//dZzUoua2ezz0481VC1p6DWGGEr65n7FhVw
pk13Cz5VO6xTfrh96fcW/mCPgurB8F8PmsP5ZpM+Rknr/OnsIuJ0l3paXBM33I58
a/IS0o7i+Z0YGtO/xiMIvs2xQeeKrgwEwLO2bEnnzTk2hPCLLoSxN2vm9R+7lwZB
Tu0EEcvCZsMpt4kg3L/AxCJ6+YR1GnkgIu4w9R7yBZtrwnd5hI39uBi7LBvuUVpt
LMJZYnLakIoK6XXZihaHLCdon0ODR2u3LERt3dHxUWwRlYX/qiVG87hKq/KMFvJL
MVZpNsm62XBrVzjQ0CbVPbSsDgJrsGU1cjQRgGX1X/tp9f/v+PL0kCu+3rnmnWhm
1cA9QTiuGUgjkB0TKfTtcSaJXoGOeuOffSFOJ4Y9oK/Svz/RgMKmePZ+XhmLzliL
imFofgWFbMOG3dH+iy2V+iyQwE7wdxZxTWOGz2VHoH6Le1me/glFF8v2MZqVeFVy
B9OlPnjAsqWhzRL13SOSxb5GSoMhwvtBl+OWssPsyl6FnKDh6cCS1sfHbK6sbg64
hi2QrZCpNzky93fdet1gOfMghNbiPFLM6NdR28P2GRVWaW9Dmg+OsRktf+e2gFRo
nhTDQs044KaYw3RBuJBQatmHUT1oK1uG/Dm2+PgxD02QYI0b2miDH9peFGsYRp0g
bkDZZg/Asrww1rOFxVLzUNWDZ9bQiysQfZcHyx0StWMyWu5ymFK5PVRcoixkkJKl
1JmqIz090/bkKWU68oUS0tbwYGfWiFVCMZ/aKPZVEhcqdaaAiWbjatszBirT298t
HtHzcK69m7aUhhTV0WFdqxCoFSRTzKeBbij7HDsl0AOEbHfsBQYOY+0dyi0EAcO9
3ETRWb2FClSFnKuJbPZlDrtkvCTRCjToo31RrHU4i2BSjH7VccDHJM30FCYWK9ol
nR0F1uL6yfQrfX5H4e1ySawBwcfHgqlQfrhjIDmOuIFJb93Lpqz8sgt2rck+CQyq
ucmxTuMX4f42nfmRTli01Hb9JtDYGruS2Jj6fbud/WJCS1N7t+Sp0SoLNkK0kahL
siO0ysbkQCQDo7MvXRbRpKA7zNhQyFMZ+nQWQLSpNUsXNo5Gau0B8g5+z0s6EeGf
whZdu334+5KpxAaAbyV1y+DeWjmeOfkW97zfwAr79IMMgzTGAg4ipZMeKXzxuU1m
f/fPH0Yb4TOaTozGM8b11Uy3r+izV5SFmly51Ei3f+5+qiPY+QIypwtWRNBSOUxo
SjPJRzOleSdsja1uYeKmjDH1pST+ABA3h6zZIOT+Pyzh+dpF7OgU7iHBEf/I9EDE
jnLHCm7Zr5wAGiImJTRRiech4wtbwIPtC267SLEJBQvvFiwrPN3UsO41/4x/yrJc
JvCQ/kbsObwlAHu2bvDBqmHLX3ErQI+TWbSJbjmksZGvoQRq7iXlhRIIvj/OkUcU
BNQr2DvBw8rQkCQe4gZCPRQy7IolX0CNjRkMCqeXBWLo+PRUd5uguHa40jaXCsnL
GZmoNs6EhMQpArOcMkv9u8ImRw5vWFQPTuNdpHJuxHCvztw/ZV6ZQ30RFvr847D6
+VVHx/GCBW8HwBAt8IKMKIDe14g+eQIeq7WbAKEVe8urZBaGKBSjPl0W6049IcFR
0FQxgvKoPGR3YgLrtCk5xTQhwwM4oM1K5q/AqTxSzlWXqyxhe9M+moC8H/VzlMvq
ywr1cb24dzars98EZAibVnc7n0Reqz0aIUcTy20g6/4328rwJh4cgv8xt9rpOUVC
64m1inrn/5YlG1RT8XFngt5x7heKpW0M69+BcVJYvaL81Qf5Nxm6NiApbiSI+GB2
Fp+cZuYjSx41bbGD24Qhf6f4JI0JukeCIUNGCOO6DPyZBJ6/Sd60E73qk1el8+g8
dm7CMrzNecKthjWeKG73J/E0uLXhdS8ERXK4hxgEjoWIeez+d4DaYaEdwGudmsgd
G0yAOQKqXejO856XymkVHegYiQ9Iuw+z6rGNoTlAX39n3dc4UTqhiJkPBXrIou8X
jM3/iNcPl3QcPhG1QvF6hm5cWSjSfR9SG62Dbw4rXnIEMOPKkivoeDU8en9Y5flm
o3Vqr9voQNQLo6AGcIeKQph7WanAabmrVge9cv71RTRhk9HSg3bxbUJD0Q/m+9WX
5gniTO+KWAtV6APAR58p3wXQscfVfkpkU9sBP+aw8lGD6tqTXAylQ1qZYg0hDwLK
0YV5WaA0xDbhv86wHkm6q+AJoK90pt6OIVYQJ++wcIcBANzMNTCpnQ8YubnUqar/
pYgDHu/FOIpBWvErVXTXInHMdXKpzPRweR7gEgrz129xrHiWYBLXJ2B02uGoojkC
7XB0aihv2bitRq1UzCyqcJde+v5QKmUOaycSy8jZYfAp9U0OTzL8ChCPwIkh7y24
jhWj4TIDkPwQKOsoK8nZEIOPv2V1hmq7NOZOctpfYoCyG2H4Ey8rKT4p6klUb3QL
dTaUfxnpporSrjCNSgPwjNJI18jgkxqaWtjcXpoaE3d7j8HyVlSiIeYxiPE58Jh/
0sxwYzZTH9AD623FOPPG7z49nDf05qWyEiA696w1N7FuIwSRcgTl2hZkbRZQDUsK
tT08nUD18ythUvWwCp/rVeHzYQKR7XFyFox9gWztOb37at/R6rNJJtrpi7yMp5IS
PFDQgerKRp63MyzTNKgoI16oTHbT3CoLdWopARO6em/LIdX4+hJgmLqE1XtJtQ/n
SuqaH5HSFSOhyDKQH4n3AQeBOFnqrWjAutRy3oNOlScDcpF1qYVn8u1XEG3KHQem
rwjEGtq/Askqh0icr6T3Qtb4MaNV6G1Iul0KIFeQGMGxVvjnR9ECzQCteQIxrBfH
HG4Ia/h3bcBwDNqQncTOZQBoN8qbMNPIuuneYgwOPH7WJV7AeKW8N9sgprUZOvOJ
AmRa5D87MTgT+wDdd/436FZkxhs1VOu4yuh+aKr5fMGqptLnjIGSszoAbpHA8VaR
iOtKEDQ9EtoJia9CyQ7f8HNj1qxGSlnirv6PnrmsUHWwyV+6lb+D2G9y+hv8XH32
IrneVzDByGIVxB1wQB/AR+6dEhfOpXs7Zd+o45yXa6Mr+a/M6Ey0jwnutRClvuGK
Y58NA80BlVRrr2Sx9y79rj5utsnifzyAncTObUQsdldV7+6SnK9qEPU9hPbrvhr9
xfC9Zqg8n8XEyvJ/SAKpx8Yt+VkCUvfzsqGe/WaIW6E2LXlwSED7l6rAfpQiFWR/
Gp7UKezoiCvrzriT0KML5nEl14gKat2BfuPPgDXj07+wRIKMcKI9Mp171JH+2EB/
7DpLDe6bdz8E6jMlM1N3c5mK4LIdln//id3UDoOAPCIk8fhK9nTczmTIwuv45+yU
MxfZUelqli53SpWYgN3XV15+uPX0sT64zFaatq7aCvWr0UYBsmj2Emhjcl3zSiV0
Lg1+vJqqhluX+39VZC5cn6sYQy5hiumZI8JHaXIlSR/J0HzEajHZfInF9jA5xsyZ
McGU3F4axhRoEraMxKP2aP3fpvODFlFolzeIfyel/a7q4ap9iiUTMkiYjkNZ1O1K
1dJn1pNxxAEeWuwtnnNLRIIKYODmwTbf74r+f0RMJYtw2k8cpyFQ9s1x+AWr1Wr2
mCbkWDrasXERJsFP6ZvN+sPoTl3lIntadwEBdTuZ7QRbGXz9eb4AZHNhBiLt4XmP
7oxwdEULEnjM0IkN0JO/XAY3dxNjJzZqSbc4sAwJvfzNlgxhskA1Sdfuk4VCAbMO
09tY3aYdVOkSpQZmpDQ8Fc1k47Bgv0B2JwTthMABTK4hVhBB8iZnt6C9Tug2fZMs
FqHyqnZXjg7KGAoomgOfoJrSEZm7ihjSUYZd2UpBBaGFdhROQesWF/oXLxHnOjni
x988Ns/7P8R5edSIFSm4ggBv0AUaAGGdKp2SEEDJ5KDuj5+N1RXZmEXiQQY3E4J/
4FYs7JxQzyawXTWziyihodFxH3maIGwPrwSZCm3+Uon7so3W3HGKtHf9peeifArg
ZcOy50mIZnzYT/cswFP97Gf681vY5PvLypJdQCgyhv6D7sKNK+W1ABy4vNnHn2z3
VUeDq5e0PwEBqPJNQTh/jM/Z2sHKYaZQs8Ery3XaHWxxk411YX6E2bZaJkt39iTT
DbKdIManLOClB+mJVpfsgmLLWltLotWar0j5BsjgfqiAFIqz7z8t9UqandX23+db
N5LmQXdbkubX4+TEy4tbaj0zKVFajmPT08Xb0QKHRUB4fylZ/XHvqQz79FmgedRo
mlgMNYjXZLj9fckqDLBWjNr3h8Hxk3cGWucyHKYkAW4lFzepIL+QtpK5ekfEEBE9
xt+UiDuDUCW7XvzhA7raPEf6IZ/Aqp5cJcStuFFBm/JZgUc45vQsG1ZkJ+HwrrhY
UllhYvMIT2cMsIS7F4HxOR/qxuNVjXBVDgGaUcj0P883QfIusS3T1DnFzYxiCAoh
ebHwjrMJtwIOZOPtHMl/Efc6akCtBFhUCMcBOdgQJ4mJuCBZBOB97Q9HCuh+s78P
IGykQMkgklpydai1pyd6+vZ6L7xw+BjAa+5gkX/dwtBDnVSlR16cC3e+xtAfZqHJ
HixjpQQ0/yg5fwyJ+bfLVdkrDJZcjEf+PJtrhun+GFCOTlOg0vnAd79oy+/mtJkD
Gba/lbrPXwcI03o2/X1/MaYXZr9yFzBOdixNFV0PeQhbhfXIpYU8eNSWSK0ACUtG
EcWDE/Olg/uayhI+GRF5fNKCYnhgnqHkTXOjPdtFAqSz21W1P/8TbsxB/xeDRPAZ
Y7yOXfQ6usgpUiO1U0DUms1H60eKntZYR+vheCCr3cZXsUmlVboUhojZYknvUIIW
RqfZuGow393+FbVr7JezAaESUWTKPq1jNC6w9fGizIy3YsSx1VmTRo3Hmok9iS6a
ToP45OmjGVE+23I4gRIC2etuKZTS9PDmvaHxZMDYVqaIz0+MmsYtaChBy1J8NlJK
GrjaAdzZ1J6FkoQuAokbHO8CiUFXeffEGUgYiwCapuXIh/Bk4v/IvJnoLhL3+N2G
TEXa6sZtBevZgoY0vklmMMrrg0hZjK4rEopxJK1Qsbg8uaxVe/koP1uUh40QaYFk
FOBfTkWhlA479zMDlpOKnIArIXPyt0jeeULirMFZLtekUsCcugUQ1OPBrx/Fp657
LQC4LjkRy41hK4wgPlSayh0Dw5/lDG8zbDG8+kLzU5Ae5xk/0MC/QrAWxTo+g2g6
bsBe0V+zvS+lyu6wPxoacX4EcYPXbBbzy9BHuYIB1r7XUyZyKqz8x2Bx3FO0gRs+
wBxmRpMjLdquy21I8Jr8HYiyeCfL+9iazSf5eiinb+rLQEN8FNGhm3/o8nx9rFzO
xdcYT19TGDAysSTg/VV8HChrRUxfO+S4U9wI3U2Ce+5xf9hT5HEkC5yj0u7Nb/jR
8ijkqW/hpW5nr/NENx93HIhwLwUfs/rEc84dxCo1NhPyRVeHFARUPd2E0/XR6RQN
lZRgOzamvlO0IVcLBVhGyE/VzbwM+2OCfenwCYhmySIn021gUGUX7MMuJ0P/sKsT
28alCSDPva+2Ef+Lu7JI5aQZlijELA02mnK48TcEX4+dyyZx0MnstvcTaPO6M0Mu
HFkID7fKIMExEpwi3XYW/PXGbC2y3+dg+VFU0nYiUNxCvEv9sr5RK+UmleMxIIqH
d7A1RmvbIMGBzOWskD8mR/b1CnET+56F4gJxM8/zIhWoQ5Eh4f/e9rF7wo7anRwj
xcFIvHQdse79cGgnKP0QqiAIhG59YTzcHax/8N3d7U/dwjXXz65gKgTJHTuahwdh
toLR71RZ/7Ctrf0BbKrSleyXdUMgeFdufTFWqfegOUS1gfwItFGJ3MWI52c8gS16
jol529AFW4vSDCHU82yPttNIiZnaoVIkg5OTCdR+ycYpYjdksKrz/T4KpTXk0W67
dFcEEX4bBYqU+XMJzYPARBs13mXI1DfijGd5h0Md6VX5CFRxIBWFD58mXRsc2rKR
fItLDYGuWKT63B63Dnd7iwvHV+wVUaQIyS/TtOv3BQaiP8F6SXvZYpGviwcwk6BB
+tLqU2La9mhX6m53dqeFChyfVHhNvUFeTYJON0X0H2qUC5OvdVaI5/9lvMI5Zbt3
WpRDHqDd3y8q3p2/yVGFTW/8auQXGdfmolQr0ezwRXVdjLu2ao1OpSSy36MCZJUo
LtKP30YSMKJiHDgFLtyqMfMCtTdXw9sDRPVv2KG+MwOTCaBSwL7sjq4pYs0orcHc
UW2qYG/Rppu/6qswy7dwixl1uc/7Z8MI7HiRZ4lgYNvbOsMHnglIw3Zrt+r8wXdy
gNmaj2AzPSfjjbx2zTVaUqnLQJq4tuSfqmdzb0f4113adqhbYsxO7i0rMcA0TSp7
Vz7C098S8wLILzJ/68FMmtf0AQK6wJCsPqR+MdXQVg5B1LrGiwRYsBUmvyj7btmC
+LC/EArG0Ot/4IW9DGnGr6TZeIkvCJ1QLhn1jRpK/DZKHDG8WtNbKsiW32X8Ik7k
5tbpGnOmJePcLq7nlpjeXkzjSLE/aYqBIhAEUXThSpAGWnt/XqVF9fH20svUQMTz
ZzxKJkTdS9H0uk6dS8RgpboknPMvS4Sux+QdYfh/nsUu3C5FOHgUXdNS5n0BRWdP
qEVnzJNdBpk8lBHOQS5c3Xl91JrZwXPxPcP1uWYy4jjv7Vd2PoX8Z8ez4+p0ggcE
IjhBugPi24oPJmSn2e1Yl7YiTf+dzSJ2eI2MD4CL5KRULDCWvFUt5WwfJJ6ys9Nh
v6pclrnHoCfEAnxlCJnyqYh1vER8kAph9JM3pRcNDh5aNEX6Br6Cfeawl0hgbAoU
7PRUVbqHKKSByjFKysbCjfpm5PecTPlDJwPc+L4vwiInk0x+ob6WCMjQ3JqbsAnv
aFFoWbkW70jvhlhumol0uo0yUotCK9HYrFwbHNyZJo2aa0YovdfKW60nhU7QgB7v
OrtJExJS52MTvEmAbIJ8LgsJGRrj6ORSfnGmhtjQYJgZT8z9wj3rCBhhWrbXaVBR
gyDGq0/m0JPMThacDn53Xy6eZuNcz/ffkGGlxJ0ZzXWhyHaihoakwSvrZQN9099e
bzubznI9fD+DDJsp5J+FThZ1+Pko3+8Deq6njJZStFKfZTbjPDEWa+U95oVtsY8L
y+GZ45u3Y2UU3UPeWhI6Lxc5OKfrTqMKbRswQTTF+DFqF/2vSzq9uhiwUOwQ/xFQ
bKjKhwFZpLEA7vLEHIc5jOOXMKDSQ2rypmblbrTllRV7Z5j2KxdNb3Th6nX6LFDq
r2ukNpqZn5+zoWRLoThQmZXstKasOs+9IpXqn3Ac1XhTmx2IL8Elwb2vfV5X1kOo
hjuOr/8ed6eJGdZ1/nbyhm5gmKAPPZ0s+6qlCI8mP4hqCN6sgMt1CB7jqNMq17as
SZXF2XDyD35n0z6GPaIynhWhs9jWiikY6k6gj26NHtbt/ad2eIedR2jTvR5nIUjY
mLrpogycHaciiOlTAemkW243VwTx13aHzfj3mQ1Umlrx6mlXknrcVP/N2DBsOm/L
1H+8CHudh/2CGZ6TdeBxzs+5rth3vaqCYjwLpT/hiLsAtTma+iL/OiMpxojytqXH
NUX2c55H21BfJWoQ+owk7HrlIdrLIpSxY1oFLl5RY52KoX9PIeVy94BOKA9pOEDy
0qUjIfDIU1Ma1hxLeG6av2t8PwAGNlO5zy5HZ48+YNQ7R1ttEQhigZd9CWdegnhS
wx9S/cl1Q+ZD6QCGPNHu5Z6MGQJEJpa6B2Kgphr06BgqMjkw337e98J7FVhr35US
zzUuYf21E2MM7H4ptdatYMuPsBF4HBqS4/VnHFzjvo0yeyeX0rgK5wb9egN4fral
ZAqNnLX6B/9dLTd4dYutyMg1vnafE5Q/oZBOPdwL36yAZs9tDsimfBbMZAZmA9BE
BJrmbpPExLBx1cX6Tp2h1vHd1hHBqJVW3Not7hA/jBkWCqw0cBgtu+Cj1G40OMWB
vS7JIcmHvI/WddQkrQfpOyc7d7lNXvFJgZl8FZcBEJQPi572wczeoFfjOOLa80n3
i3DwWZbseqK5xKRe2FI2QLLl3WkZaYaSf1y8IFPC7BRcxR3eCDXWjq4b44tKUiVo
8SmaTfZbKjuymF6N9ZriEHJcu9u0sHoeyoXOJrV+HIJvDjIEfHmF7E7K9UxBx8Tg
IBdFsqALE2z0vtmFF0rmkrhvM1sab/RPD9YfZXkvneoNdJaF6I+jMEPW+cW2syv2
6QxUvwBV9en6LBgNizOvVs56hwL4vWoGSUoAbL8xNLgqsjbuc/UWm1cyTQ8wGAEx
RyQ7xxdL+5A9SwS0eFABFWAkXMZvGaAnGpudcbrWsBMo/QH3j+LLjqwdsrbzxCxT
MRGT+FI7QXdwLR9H2Fdesf9XkcaxykbO4BmYDcO3F96wwyJdLLAm6lOEviFy66Ju
F1vPWIU9TOD7yGP0cKJo9gIaZMEY1ImnHl4cncdU2g6BKLDsI+39oPr+Ttkt2Mh/
MTBX/RrB+Rl4zG7zL4qQ4DOphCmEHAMRYWou1IZFa9vEPeubMvor8EpupMGRH4kC
ZgTWDNyzkeTcPRibZOD9N2ykbacBti1M4v2qAjqTezLaTAUB1U0NGIppvL7G+XL5
2xegAe6t8q8+0w/2BKBmfYT9CcUSjRrPqPYBUrKkceq0LlQlqPWTZOl9ye6BEFPI
BKj9GIZ5dILSzDldE2LDkJqrcetWoOGJ1EoLHl+w5HQ2hKEvRJ+Uv15s5Ql2VIju
ZBNVimU8513xMw2q6PVeT0AmY/u55sEJuEcuaYcGne59z/Dq0eCvZ5+TV6SC5Y7x
UAaRkcSUY3D8gvAXCxkB8ICUIiB7fOMRu8BzMSIMSSCLW3EVYcUYoIs2NSfS0GHV
ZWyQcVrH0+mRWsLAh+v3IE4viFi5HVKrDvYdurIJ+FDE9dQG2JpvKzIUxWvjVVko
sbxxVJL27BpOQNfuWkSokMjaJpm+INhI5d2vVSKJVo5JIo8EP6Bb01h8PAru0ZRV
hPlfJjUZL2zj3Tw7ba1TQdbHoEwIGtoiNM9BcU7/PrCeytyPJ1sgdZHRF0SDnfii
5GYe7eUPQHxk4lfgMRr1aAZgqp/80m67UHyaY1Xmtv+NO4W0RM0qv/Boakh+qxpq
hy5rL8eRNlvUIwCxZmYlLe0uCMdwji1b1V6Fmoi/qEMbNpencr/9pzl4RaDkGu2+
WRATWyoB9rT8AP3P919RsDo3CQXo2UU29E5XdaRkKLWyEh01HxWsI5IrMwetzVV4
MS3jdlDSnfbmYUqsnTh8FEG0gPyBF9cZC1qRrZxaMglgzK9AblCsaQJrulTTD0NN
ppjbfhwakLpFN60LNqt6+op28uHCOITPtSe4FnrM9DK0A0s3rI28B9eRGYgRU7TO
7Mv7uPsCj9+IpAS4T6CFBhcgtQgUrI/1wqCztwvIaEwl8q+J710ZZN8lw4duCsE/
+0hGSs+oi3HXdqjfQwSNR7k287NZjq8TXlJ3F3wD5Nl70uI571jMc/KpF8T5OQpJ
SM6KI5MY9OZVGbfAsOyknFSlBFabYM5hvJHZ2HCH6D932sJlzgfQPy8phOuiHno1
bkD4TyQpGZ8PkThPIDDOipWiuqusTgbsNDYLBZeNjMMxoQPILaGtDhKaBK2mkJZh
R8ZuDr9SMK4AbwPNhp0kb5fRIf8Giv+mWgnMEjGIxmIfo29PAvRo/jBrDxigG5YG
R2vBDxGiKrvcG37IrCYmnDi7vniR8/R391YWVFMstqE=
`protect END_PROTECTED
