`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6kWhZywA7xFHCmpEDi4J528uOHIVYgjGa0CL3HQQU8+3ryFKHldpiu+FFGlntpgL
Yb57SQmL3b3ax7RxpMaoPG19ZY7z6cxkk4LYQcD6cCY9K/+Ea/t20TP3Kk9ZBBVc
zDQhQ1fLa4F959J7QrBMTBnuMnMmKXJ5hrEwMqFQElAFJ0MNeuWUUXRth2Hq4bMN
/aJ/cqf+TFoNjaNlzh3l8iScnlMbs2vS84MnP9A7jik2IPkibKuIPIPOQGlABYTX
VJreFe+A+cAi6dVrEkrOMFF3lTFAc1fEcI+tqdn9/eOXfdbgaO3bMRtVl1DFGE1N
pofv3zXYq5dmZXHhH+Yci/fMROIGJdz2pCUkihe72yS7AHPiWYE6OODauo39MSGu
nbEO0DCRJdtSuG8bG0Nf9ayWf5J6ErdOGBQbO3rOzWul4U6plcikZ/1ay/fpdUsl
iZFYLB0IAUck9mpWdbxF3ZHpwUahoicgxgam9KVOIXQ=
`protect END_PROTECTED
