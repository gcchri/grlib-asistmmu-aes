`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BY1OuqGys83skVf5XURTvdoXa7NaBKddhI2Eqel8FIFuzAFuf/PlVQxTb0K0Q9Tp
+BpV93JzMtK3EhCXl5KMYG3giN/2LtRhTxU96hyc8mndh9R0kC1uo9hUD+LsqWUB
lg+2tpcZ89MnXfWsJiu5PX15ellFpr3asMYABSwBiekz7rPZE8Q/LFecnlniHAaw
h6gFjLdYwPeB/P5u/mpdsl0TQb3pggOE7B/6r3WoKYSXihvEWOPeaaS/q37AqeUD
qFNzkC5Vu4a479HAq3q0KZ3sXwDfDWKDLLDmvaKDIpv7njXE1vE2F1EVVusmmpWo
zm028aM+/kDRgheyS5kp6h9CqvinDVIOv1njk5fp5ZXdwTyAZIlOVzzd5L9LDHHs
H91QyGOOucvzeOROvrZhneZgX9jFYU8zQUQbOfjIA10=
`protect END_PROTECTED
