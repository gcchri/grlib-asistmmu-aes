`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n01o6eYbLEgAN6OuMEzrO08Ea2I9eD3sSGMTKWSBIFtEoeczoZFXIQBGHyxyQKZd
wz5bPl/fbK0oTThev9i5RVl2eYHdZ09Pczm+FgcXd7vaz5fqe6+qQiG1rzRs5+wT
u/NnTf6/CRUcVz15xr/jSOw7FYfeVMXH3C33t+e8iaSt12xGvygrQb3gNTUd4HcN
WoXyhKTIQWtQWKUdjaKzVv9eoXQTpTodfos1iSBXNPXxu3p7JFJrtufWcBbUGz4a
pId6tOdMPD+eXGavOxL+dvgcx2/W3YJCzPDWSxfk2RhT0WH1t3c18JJqFvARpdaT
Cd7kcBYN+crTFIl7QQECeNSi3/tlU7iVimYvIuTH8TkvG0sgJlwoEhawwV8cDelv
X9keHvvl3rhhT8Ji0V+6GA==
`protect END_PROTECTED
