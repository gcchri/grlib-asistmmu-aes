`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6eFCsaRQKc1e8DzgIxuwWoB7no9IZol2sQv9irMIaGLVfkMYlyriU9OGF00h1Zeg
EUq4IOnu7S8Y5q4aFJgogqRUYSHO304/FJFcryGP5ebuvVlR+a4fMAc1LCXAq6dN
iAVXZqieIMz1tty6P+lFAlXb1ZcVsIu69+qNyUXGrzX+5U+0YUDxoo280fFOkG0o
8TYSz27xeEqktJ/IQfanU3OFUuDOuswiCEU4K6qDUH+nvBfS7NqclehojwX5AHU3
osCjrwcg0hzhJNtKaohBMEgaMyqJNdYwEZL6neQPgf8GX3cMsaKiO9frzNWsqh0f
plmC9dmkByoAK4PtAgpMESS683Z7p59IsLmaRJUgBpZ3YN4qJe2LaVKVe26/sjsB
hzyMNi/RdjtFnCraFWavaeyDbii0h7IOTSSa1K9BpwulrAYsiZdvUrEOw3LeQq5z
HhNz0VSfBIUGcyxBeMRfyN0HTVoeh3tgI1SwlqBLU758MK3uYrTGq5r7Ul7nBtbO
KlTUdRv5X28bMpcYwRYIv0giNYJ/cOajJRAQNAUljtAj5INgVWuf1+9WYrXGT7qE
D4AVJWrMiiqE+yoHz37PBIfzJ6PJ5Ni1CB7BS3Vp4W6dCDDUHY7irrJ/8+s+T/RW
/XZT0yb8+5B17FRcy2uYBrDK766+NJkkQIOAmbDhgcHFB/NUwv35fczO6J75CCWc
7ChXfqBk4pNcSAudlLmtcs9dHr56pUt5uR69jM+9QeJsPA8qqO8uWrc8ns4QphDb
zT1eDmZhK21/NtsvWiwdwrbV67qBrdO6DHVeT0Q4pr+ygne0oU6tiszgO1IxFdr/
HlqZjF6XfLmYiL1fO0j6AyYygFvFWmdd23i9ufObAK17BSkVxkmmmNNkFMFDbK6c
UQWA5o0mdHUhVY/En475F3k++Vtc9eE50jAGrei0MtjaYz5hXGgFB17WJmymCcLJ
`protect END_PROTECTED
