`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OlosIZwGxF6YcJT0tYLIazVJrMK7pDAbkWhpFTJFpgfQpO89ZajkkKJRCM/Cn3Vl
7oyrDKcMeQFeUd+qO7ytlzTGnk1ufDrmK9dR0y4C+6XedmEIg0E3tB2GGsr14Wm3
i7n+PEem3q/h1thlc09+cXL91RAG+dgNm8JpSsqJi5O+CrYqq1jh6Qw2g+pwQUfB
qBSQquRTvr4HVTYjVyRdrMgOSnRpOBgwFMDEwFbpBxaduCRW81FkRHswH+CMjJuU
7oy1edyDqFkjHTagakmr/u7uH1NOshUb4278NX3bWqH44mSJqkiaYJ2J2x+Ybbuw
gTB/5fYypsX9/5kMDuO/oz5OQTtiMDytIPkE5q/341b17cAdgiNJBRCKiEfGiAG6
u6qh4cmzxUCN191h0/FNJfTxJJIO+8CTtPTtcXW2KltNvM8mbz2XkEhiTrPRPEXz
lS9jiWf5CmQHfrsJu7fTg6OPBN9N4FY0VsoPX47OTNC8nqg2TFWHsvuo9nt87YuK
+9+DHUE4IFd6FNp0N2QWvIsqbHKQmAklK1PP+keK/OyXuRupfPy1ZvT6RqxzmZc5
izldBHqjCLc944ZLieSdos317zZaK0xMytKUKG6/X7ljx2dmdnkBLheSah7WTnsn
ZXPSyTBtvVsG0ve75FeU4DVUsBwt1FfVM+7ahl6/q3acwofIjDog10GRPFayUnE2
Q1PM20soM6bkZeumXaUQKmNs4tC5EfKBLfy/iwPmugKUGQRZHUJatkkGggpJlXUm
2EeVLRiXWuheKjPgnD3oXishIpU7dbO1LHvIEMQ0ZynVogmLMzeccV7qQTptGOeJ
f2PwPCtB1OUfc/6QrO3OXw==
`protect END_PROTECTED
