`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tWFAPPl9w55Du9b/QUF49ypXwNlREURpZDiw1+JvbZHk+9CxAE+7ZSFSpOUi9KuB
EPruNchOoDsKRQy/vy51PJGKnB51rkFpiLYLyDeinpDr2uk2JccvHlB3JGWFFsCf
vTJJx6GFBNR7raTbtAe808ckrY8Aj5C3vTPWFgApA985xtiw6+y/JVcfI1VCUxzb
I9tZFkcEXKRnoPyx06A+7KTgj15CGVF/7DvPwii6AdtqWtx9tPLx1RJQYGNyjfeA
AhmsJM4YmXcMoBqcZtKvCR4Ka45Gy7a9tcUMzn6fH+ygm2VsZVR1Lv4Qq3KCSFjO
3OTAhYd/ZO7Rbg+3VqhosiSHHzDdHuDrQlkfdnGOrJQNyARGFcaKs6Au2UWkHzcc
i/Tpm/u7E+QRBI7rV5oI0O13Zz/QmjPNF4DuGzPnVTFOrlNGUQc4TAfOv3Vfmud8
Jw11YdUshxREInPRVV6bXqGKcOTJhSfC2DgamG1Vh2kPsdYZ2G2nod5o7CUA51Qx
`protect END_PROTECTED
