`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vNpQfOwuc+oF7jrZdSft6MluDKyWaT/qLVPL9chFeefU9EVRO3jYigkOi9Z7rR0i
Rm7pWRc8wt+mwoXqYAtO1hkf7yXu+91rsnBDS8bS4A/iAZKjbrBKgkwa5nPgCGu/
y9S4bRX/hxh4QKNwSMM4a9bc4fx6UyAZ4jIOFxXeT24qzgpcsaa0sIfLGZo2b9dq
X0dnDmkVS5j7VTsodZNmODz6lYHJXYlbRaigTJaH7w2fKx//ErREHaFE5XZEvtNh
aEp3yKE/0nKnxLTMN3fOif2damW6y+8ek92xCyjsB960eRGcX5NBnam1zRpCfjkc
IRwgJHAo1L+lgJVzRenMdIoapgGsTI9piXO3CFq/Kh7CHWePsZRpuzCfiK74KzMP
`protect END_PROTECTED
