`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
430bk41uP29NO0ip5mbzejxOEsXrf2rQIud+vz5vOj/sBcGBM3VeA3a663fZS58l
idQAwJtmFeY+UnNBdRAxBwbwhMs9oNEXOrzdNwoUxw9WiUkfitr6DYXrMQzwozzk
SVp1FIErs5/LOzs6lp/kownh9l3xuxvA9r+3e9JU4X4peI4/D6QG7QAZL3ZCBGNy
VhEI0GZg0UCWw9GQVCqj57mwiE6sj1FhVzn5S0QDms1NrWu6R+16KNG+pcI+iy9j
IWPj0Y4tvjpoNAhirASqON9pD+XXIVOrQ90pbprp8k0=
`protect END_PROTECTED
