`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6M5FfAORAJiKMTCgyC2grw00U7P8frMMF4wmxZjnAU7u5qB1oeX7vIOH0RoCEn3N
vUxIyF5Wrniwk3ijfiqULE71EbWlpqdMO6w2whmpDGGi7qI9Mk7BsrcgUjoP1AJR
39GtVrCIGRKyvKtvHa54PMwLE2Cl+ENBygRRNEdHA1H+DIvWj6sNMdYqB+j9aJOj
keoloL1UxlMgAatAxNB/13Vz5EO4ZzRBg2CsLuVtJaoC4McNL13Eq9gR41oNxe3/
41vnToDBN+J4oWNng1SdC4E3mSXgNo4ZwbeyfJJIbsKSlB/GmsxYpmc1O7Lp4BZv
drCLgwiKaRFbxzay0KvV4LjTk43uYIg1Xr7eNyZaUC+cS3gjiPbfqB0DUWoNLJr8
TloR0u1GDSNW7Yb1Yau8eMOSh7ypeaZo3sfDW7YEqrIkYkcyIHngb3a5O/vvy1Hk
XkSvfHUDCqfGqpcuNfcsYZA8dqdvX/A97TuS36vYoJs=
`protect END_PROTECTED
