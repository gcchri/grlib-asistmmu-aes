`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HvMO24e5g2dJhmQZ8Gzfp8cQxT73WwdMjma0Cd+vQNuVLSXLRYsVW0tPv4opxj4i
Vxv17vWSjeayL+XekBKBlHSiiN2ryr7yAlIuKd4B/GC3mrolhNw8HMMyAk77D77f
9hhDz64sfWWlgRJWjhUaT1jx3PeQ1EF3BBLcrlyVmF2QZv3qhN6nAlXFX9CSU6h4
BHdL7Nmj7T8URpkhpEBXDQj+N9/+MknUtg8aWH1VLWXPP9wOEj8j3p0OSBJmnaVj
9avTfhUGnrPe+Kpw7r6UM5TBQTJ3hW6soqt4/NDFVnDDlfKSPOUq3zZrnMGojICh
N5DngznHpB/27Qzvg1WKZi6sCgMvMYr6Pga+TDUt0ndijayL1yZNjl/lQBGzgcxx
erwA5HmLlBC/V6WHvAKmd2Ccqn/2v9x9UXYAearDX2r7kthPbwR5EGzId7SVmvXW
ZKP9ebmpXBQA0SDLpzY39LjWHbA3bXBZGiHePp06xIj15WbWmosyKWIguvwxN+5o
OFpxzaHyjUu3SgL6Y+j8gH5foW/cN7pWApGdEFyxPGUEyvrGIvqC1VbC0GnJSzoS
HVZgWgnxFXxTPHrk2GhEEGhlItB03oeA5FrN1LuCsTzkvdbo6OOMDrsa95U+YjUC
HqDw/k0338Qgu9F+OhBH2A==
`protect END_PROTECTED
