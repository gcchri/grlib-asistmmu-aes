`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gtJoVsSynVSy/LfABXevPhJE8HUP6hmB4mB9LGTQnXvanjI6AxDtCG5eCS21ljfk
cyFw0Btwrwt3EL0KhbPmd9e/Rq5K8xDIs3XkYl118Yb9y0wIlPkOzryTnada0JM5
go78XCY2wjktS2Q9R9f8O4hJuAvSb6Ky/osSTF25NzFmrT14ADAAy0kEqIwD1CNn
B8S1TcdEq2yPnZJW26vjyMzao2zPuYK3wMlni0swvSG76mY38K/YxS2q4IlMQq5v
WxOvQB1H6ZKlddE9Ccw/K0wCUnG/1aiLCS/mKGxkK+iKsSzDgL83sSODZRG5Wkjq
`protect END_PROTECTED
