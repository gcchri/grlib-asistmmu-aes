`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2MIsAxCDT3FWW2k0gXjyKj9csyXg072WNLgT0huLsKM+rjipmldfRt5h8S4o8iGF
e1vFWXQKhde+4FT11rteI1UdYY/if3S+i8HB0A0tflky2ceFtmPb4Two8v21Jn7T
zdAqpUgk+WN0ujcR4tvwOtFeOiwDSpcgsRSistt8L/3N2qOT5b0jgUPgmfDgdlkk
0cz6zmT+tVWkKlE1cJk/VCwn4/uI/hK0N3sXsg8ZxC0mIfKFZcnSFgW8f75l4jSH
gegDktYvWI5nInYB6PFwrBmaAmO9XC2Y0B8A+zrIfefXPNQU/bxDetcx7XspbCrL
YRTxHS2ZBnLpJNAx4OKQMcOxZ0u257fm1Lp/sN/b2V89UegZTiNeBRSLPW4Bkt9U
b2QdVowUEmiZIcDOikV7KB60YvDy8wotBKCsxHohLr0tEcUjmjGTjQWtoTlFckGw
ej5J7ebRnL/US1adKCv8xfzWPj/nytX0bSP8yNEaOHRVRly1J5/jJNZy1NXpdT+8
V88ThPHpdszuVxE55wnClzX0FR6YHrbtQ/APEYixoFU7pFm/ESfVkJydR4l/ji+x
3OOnq/IzhrDe4rL+d8rMJmR3MD89EQ5Gy9C0gdWbiAAxiLt/CVpcuryIAAqibZl0
W7O7hEvrgaJH4hFYXBs0P2OQ8VplhvLrjjtUjJSlkF4/jPfRAoqRUCFCrjjObCUV
cA1u/nHtMLU93gxcQx6xSa+LjOmINf2UJNlOgTc2pxzbqyrqKB69k408jSchzTsu
UZbVB1Fcjg3mZimNl9smrKjhekwVGxC9/bNTFE7T0Js6YbgdqvzAAAKwlVuSm2GB
YmPoVDPufBuOpcAFKVFSF1hogBT+z/QbruIZhDLhR5VwIuyT8+CZWAxXXcIL8Ryk
q5dHK2dkQVTLMfm+VVJwYbRb7pMm15EfnbL0+5kYJCLyhckDNO8Rpaz/BzjMp2J5
5OKDAoXqSCQ1zPNDCHe6O5JgIC+3YcqVf4DtnZOVVVEuCTNpOmVuJatgDHot+dIm
YzLY035DpLXViF0poFNedUXAeQF8OJ/227PYmDhXyK9EttdMsPy20dGUn5x+HDJa
`protect END_PROTECTED
