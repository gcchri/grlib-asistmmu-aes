`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FCS7PEBDNRX1E5f0pCD3AjPILhKwQOISq5Cj8E0kd5dZEwrkxc5T/k1pijLKPffb
Kk3RcH2M7jEoABUucptJ6Xb/KRpFTgUXP9/OYF7fNi6C4hkNsh0G+aYQFZjqiAS5
Y2wxzsThpPkgm9P85QJtd4qkK2a6OwfhY51GsTtc+EYmIPolEGMytiK69o3rO4K0
uj11VA60BinRDMDhEriKnmZgOkRgO7Bc47qn99gPZcxl+nsWqxxyG+TaKmj9R+KE
sKbzifBVBf0h7nwwodjbIMnwrqsIYqzyGBIzucIlTsHl835pSHiihMdcCsFthaph
WkdjIDy7i3xGOHQk2sfCQQ==
`protect END_PROTECTED
