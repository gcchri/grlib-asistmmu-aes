`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QC+bUvndAIv+WEgxH7U4rfBNP6Xd+6N8CahID5J8ICb7I95SQ1I8WKiEoqTRHGO4
BwyqXiYlOpgzK61OWbHSgmq6WroP/X8cVg/HFYJ519RYytKlPszpCPdy27LKg6tE
uANkEfb+sdNFWxUhx6+jKL39aJZWz4BMZsjCjznGr6kNLir/0h6zsqWhxJc/KywL
uaIMUL51XATtMKMdFAT0usSxYhufCVbsP2P4VQcclcwVlamTVWbjn/cy2Y9J09t8
vbZJ+f6ZlI236PF1jHvSzg==
`protect END_PROTECTED
