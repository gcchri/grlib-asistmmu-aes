`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bsP9PxtYZsPXwtR2hrOF1iFdM/qIcoUaYluZaBfV00fW4x65SSyB2/FkZXNJUlaD
To5ycY5zDWHp9FXMt+HidHZUjSBgSYq2tXq9SlMwiN5dWpySK0Y9TRY6Ak8qWUBR
2DRTf/5ezZSPV8T22l/3VPHwOOqoW3JxwWzYGzfr5KuxFYoeE/sgyoMWmmxWKRPd
D6dkAnw1+IUi5T0FAsXBpeOzpWWh+hGanAsCd+gLqXWJ+dzAuDJctlHJ5+k+grF4
lXbGhdzEsgOdGNHAFbJn2qG8E+8EZUHuzeucEnrQIgg=
`protect END_PROTECTED
