`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R2oHObVucHxcmlw56QsLwA5FYxH46FvjgxUPWcGYbFKcjgXyJgNwvdz9YrhcyZm+
G9ATIpbX72S5fKXXqzCnyOEaBcLftxgKK0grW/9DtXvDoMNnLz1XGAKMj3XEEiFs
J6fOgYS/WGB7Tn35GglAdHVSu0zCM+VRAxcrIxsblxGK06HanZiSjjEdoNwYm/Bq
DtAOoFAGmNv3EHhtOZ2yQFWjw+dwxgKC3qfTiORyDm36ND7PoPFG227/JyqbFUBT
ULgGEmuMij0R/kpb82hTUAe6mlc0wzWvGw4pJ5YOz3TRrbS+K4Buz+OM8bSaZag6
hMHPnyy6SYEmg6qws7LXfChbxL7RFVmmkJOevoskDQX09ofl9Izz2pX2kZ6/MyN6
Neah+sSaQojtsNH/zpG5BHT+xQPhGhligecZGBEVmXLLnQPTpFrhZFP5FWtZ8u0o
MVmGxX+0n9rJtUA8X7GFc0plL53b85ecIeRHIAyJHcEBGc+jWBZUku1z/K4INZug
zJohTZisPikgWnndWrgy+/8NSczDiUeI7wtKPiiaJPpjpgyOVDDqCQIckxOxcrvp
lfXSDL6RDHyFfkR3zZIPSmh9UaxZrvcyz8U9eHEpTvet0sh6dNhfvL7rytVVx1aS
e3Y4rUsPsgX3+XsetdGt9GsxCMx0RsjWzC0BecyogJWJ82h6rxEzLqqQcitBscz2
+EoSkY2pkB0N2+w8o2ek4J3AU83oFZVu8fKqk8w7QAqwYGuBOnZ5jWrBVVZDc7Oh
oymoc/2Q7UbhLDSlXenGlBvgZZh7ut6FMgZwwxTFEo6FkziSEAWUsG9rbA0sdYhV
FVGXfzSONCaYI+UCS4UaG4/UQvG3K+AjYDbQmKFc84Zuu9OGzJX8KzF73dhZFuYU
Hd6239IKfh2j7+L21CkBS+bq2OMWhE8wQK4E851UpKeV0/fENT519T8vzSrxIomi
TIb/XIZlWiCGhRUY5wdHA/F5fGvO47Ms6XTIqA2zdp69w0A0NWkOwZ2GY4ucWSOV
fIC019yXol/nY5O48Xsm20jbG2i4II2hCb4iT59+vFJEy7gvaoxjGjN2I5RU0B1t
Zqw8qXV+r3ht+IN4rsK0hOO15vy8ms2OpMK+r9swhBa4kLyzMjTCEk/HIukuUrb2
5G5Lrw/FlmlasDhzAK0YKygievlrXeFP1HNKSkAyClOgfN2TMe2vxJZflEISFajq
aGMkbJka+YiOA7miGJ/vXqk6yRHUxLCq+wSHVH+SohuYWpdW9yrjeZQNBjCx9RcL
Jkys41I4bhM0KCet3Ah78m8s7mreeZMMCW0zVqLZcAOKIosh8moQgu4StyzXv/Gg
kYkmmckjxaWy8YK1Qa26E5bMWs0BLgl0LhnZ4Ip7DsUHDViHYpfN/5c04HZxHoLe
Z9bNe5Gx4zE3VOGAwf3nlrqk62r0Cr7E93Z+Nuk6jap1pXIz9Lv/JdL5io0lebsF
oIgYCUanbirhHlHW9hTt5RQkrwgDLi3T3kjW2PK4xZPmaj7s4d3OXoo5o/NDyEsR
fB2gBHcdO2BuxSLbX4qSxUWLV1X2pxkOF4dAu7cQH/XrhXE42NBbO8Ymd9r3tWye
6f/LohIAbuvJamMDfFB9W3EekJivwbq6YLAyMsUb31zCTjl/gHsWkJUd7y9rJ8XK
Y0Xq4CJTXnMLWD2jSDdOMIC2KpX1gOgRjJsnNPyd6F/cukQ2ajQ64TIO/1S8/4m6
AuahzUECWHai0VnkHac52BGGTRciSfsu1QMi9U9KNXkKGPddDHWeVMU0LnUFm9ss
PKAKRqJ/IaKj8pvLukKmtRZ4GDhQcBEKxilxFbC8KN7BOB5yxJ3PA34MqMxOdbSh
SGe5m6H2C58U5B4JooDFdXNZGFNtIvU5eekr5ff7rI0hCXQDsVSnCUytI3m65pg6
xQA6d2TIrtbTubnYZu2S6X//Vx3W6P8dyyid6eRzMA51AR8S5mBRrFgnWT8RrgbY
mv0+tLAdOJZGEsfhHMi+q9k6PYh27oTiUkKcAjxvdlrrwg8IwkN2LFRAjHaOXqwq
rardxcE06zrTiK5UVLTRV7teXyfso1q9Ml08oz6khHIQ0F44tiKUoEt1JF5WhHZV
Zk11KZB1pgydJj6bBT8CY68EXVl8gCP7DRi+x2MmLvFRs/3FpltVBGztVEkluNss
lpDFEyMRKwjvgEpGn5t7MTexweLn0qCGM9we4bn2Tb+8bLwp3/IAzSBTTD00AMrF
S79aZ9GQjJQBCVMiWDw4fzdSGH/yC/rqT2vgG0GjjrGqAB3pxNU2Gjpj6L9HxUvD
DYmE9pPMrKCdk2smai8JpXdA9Zqo5IzDhMXhN6pQX+Whrkxyaoay3Z+I2pv+4Nnx
iQWh4uUbMFr4+kglJ71ZTRnyUdlKc4Wj4ryAEZC8amsjQcC9VWcHZ8uyvOmXTc7O
RNwwO6wBEKuTyuYsvtT3/rYN4gvORxN3TOMy7Wy0rn/tTbhi7AvANqBXMQAVq6ws
Wds1cXI0jQTc27kTr0349EpHlImcUyv9mUMKYyrH2a7icddfATH/zcAVTD8kmhWP
0QNwVfCmTto3r42qcoMXn4fs8bbDD2Ja9zY37oojgur8abeef/jS/pUPHNa8Zq1E
XjHJfpTEX4IBk1trwKPmFdkh+2s5JYwc1XJQybg2L1XKNBmOY/+Xw5uitvrJRkND
86G0rMzfcwSzhwQxY8iMRHuDH1Zho3lHDq9BAVWV+BHVOfySqQAMHsPa3QynYkXJ
Hn4aYDt2eKAy+fhsBNuNHtdOE9RMLLOYCQWgRHk20SK27Ztw+fZTnd+ivgmGiG8G
u0T44ypf73lzf6KAEi8mGVluE3HLziXbhWFmXu9wvOYFo7JTj5DfaztiV91o8d7Q
66BqBcvTcCAotMuReMwwOt8/sHG7obYflWvC/bYpstQt0ltuqll+so6dqT1GW/bo
NlAntduOfouQLGY5k67jivxlFJ3Ir+ep8iswWjO6OSm/EOOWPXo7UhQEm0syJ5TE
vXCwLrTuHhw5ZiEWcRraHRznlTvl//r24Ut8ANgWiIT3lLRG1t/i7lMI4d144s+k
SrTk1RTyUgf+eC/HoREkoh7wo7VFfDvKXlg2+8QuW0dZgo/OBQBqMzi3H+79Sxvi
K4oVyHIk5qIRfDefZrDNMTecJWEX6vXiYvRmYjTgw0hoBpPIE02HKRruGwCqYTTu
xmW99RXxjqIn/OfW+j7JaOJlIg8vkp2IkpxKOz77LCyyOE7R3uZeUyHAI8IGnoJc
Ic6paU2+RBO0gwt1IIigtFU9R2ZuPTUkm/NKNkpn7myIyECVlTwqB9yFGV/hhNb3
RdH22MzCujf8vhVsifCl9Y2vBw5NsI+GOdSpgWXyYgGgpb4LWypkBsbj4oJv/RPe
oGwn2//SVX7kt+Jf5NaNWBXFlDQwx60Xu9AdbLJh+i8ICp2N/pnvAghiUgPYLYic
C3vErod1zjy04cDrNNqO9TW2AG19XtabkwzFxQsDkDI5Vi3Fh9/q6Fgapc8l4gtb
/2hLU4L50avTCBldBHXYLLc0lz/MzbRy/KQJf5pzV/t8CYKp2kUGsBOmr5Kvzk2q
xtOqox7w4SFdPte082s/fuFfLSbD+p2Sdqqlg01JKFwGgbhI+BRI3HLpBR9wsNMi
WcOY6CPWqT35Yqe2agnjBplU0A0kVvEQP8rbNnshBEI76oOKCY3NtKXB7iPKYgGg
OgKkB/3rB0YpASBhsqkdPwN9XIXW8CMAqZ9sEoz2sUkPQd/quzHb/e0udLW1capU
0VmmKwL5T6YynakjZajTDfiF/Dt+xEQu50zgsG9Zv06xJub6A7J8UcawsCu7zmLA
Q1EU9HaGJvKDXBwaVDdJeR1vpBLE/Cc3Mx+rg73vP8+q7eT+DBCoJDF3Qaxnmtn+
/iz2pvWxfmrHz5z08mC3u4hix3DuyMTH1lkgTfj2LHOue8gTnIDB7HtreUzUb8MY
wkTVuqDo14yaSvnl3DmAWdnonfDnkt5IiqQOBcyY3Nzm7rMyH5S8Va4BFP3h+Hom
8Uci6uCqhiEO2jEygIjt17psxu0OOLZLNuKmN2UXupu8SXqOSRJc93+UJBwEH1FF
zQCNLCLbCz7itnxxSSY8Ev9yVIJAG4pVzvFF+snFq6WdmzqYhEG9U32XnWenlfVw
6xHDdcOen+WE26zBe36gWv0Eb24qfZkcQkm44onlb5VFMlQb2lfhwqTmVsh1v6W7
vt5dBqzxQhoweHC00MU1csicQNL5rho19Zv9JJupTKro2LEc4kXr1xrfWS1q1TTW
nVnLWhoDtxJ/XLOIxoBbqJqU2Rtv1ZoohvpWIlri7Mb3gCjtZdB1AU+xWIzuK2wm
brsMUQVRzSHywvznilJDfQJEWB68ZOU0hGnNAcO78t2uHNeOf3OH8AHuafUjqQDx
PwY6KqUpo4Wq3gJOK1KLtTc7l5xM41bf4bud2bN5ADX2fWoF4OVM/GXzJIFml4bE
wpjpY/BpWEkiAD6957w4SlMEtdhFaynv4w8A870Whq1b/LqthtLGd+NZFBW+xbZb
QHVmYTr9m+mWfV1c8Y+HVGqV/eD97zGhMJzf6z+wsQ1QbAqxpM44svZYbAPnR2NA
TAxEy85sXa1ifFGObcpUGNwsmMDx1UzOwpcTlRj1muVCxMyKCpGNsbsKIvcRjK7+
HmhCsob9rdWvsbLSrVetRr0kz6rcFhUGhQjcZmIsmiDgvOVlKX5vHQ6cL1NkBGhn
6KuhGZslFfAs9MYnrwim0vWVUyQuovsNuLaKb1cjWYAcsPoWLKusIuffqaf8GqUT
qFF7tZAXhl4VYfQryrCTXD7NW7ANhp4yenrlLVZbRpbBL9m2GQmGGOui9rphavtp
eicmosG0/zXbliRe6PRpGL0qSijmwE841ABDFavloJu7d3PjA7o1g/VNZETMFda1
dddwdEZRJo6XgA6pBNM5ruFS5z+Csg4+oWZPcJ4pN0Issabc3QR6BUDKDUjFVKPj
Kd6WTc4pbE7G8dz6akVrt6IpUFeiH1C/LE47QJKX0Zk1PG63iMDxXPG/KQghvD5e
fbf0RJUrGy23MfiEYg76Hsn9F+IXDra7IIlDH6ioAMQShT9ty+TBqdlF3IsBFWzo
RqzB2PufYsryNqDY30FVPTNx+bFudvCloS/N3RpOKzgaoMdolYzXxP5AgGcshtNo
fX5meR2WmjB428Kq5fdszWQceief2UmeWwsMC/VTFuwlyHzhESzy2k10u1ADqOU3
MR5X7iMvtCZF6lyzZS93BckFgRww9CKWLrX0d3JiXdS+qGKe+JB0fadbXQ0Xer+R
PdDB41RGJBsOqKyvdhmwehc48FCghVrJ5ldI9Hq3QUKUiWr9QPsJn1Wcr16yUqWN
9v83rU/0dqneKvsatzm8BVDdFSkOIIjMmrQW/okJDPcKRbUmIIJ3xonuiq44wgJw
Kq7+LhOjjPYSv3LkYAyfvpUwlVlq5vm4xKOBxoiv/RcavDHO1gAHU6+SRYRSFG7p
/5n5vbePweaPx6/xq8swuOM5hsdGQy40cFahIWoyHxA0j2wAoyNBBVBVhnhoTDWk
Zw6z3yJxrMTSdyaB5IwNjM76tGs5NGZ+xL1+bUDH9+xhAYg0PIcMVcH78D+COPdQ
U2HaC07dQBwZ8v45OanwbtnuePg0wlIe62aH7dcn1m7zZllcC8+rB09hht+BJBny
OJjiOReAoTLWWzkFSHmxP7bxBNTb5ph7N7mnG67v5cdHryA9QtVf9a4+Bwrs1YEJ
zyKO+Y07h0obPJAA7SzTJeMIRntjo1aha+8g2Brcs0D6HrWEuGLZMl3QzPxoj+Fn
gD5G4KlZN4NbmWnJI+zt7ZiXl3ImoIIv4GCPfGxQdJF0zbMeV0McXisbNg0h9fUn
vLG0poCXQRkJQX9TafaTQpDjRgI2YJLWn65pBFvqoCBXSYbS39ArJVZwtyfmJ7ec
HOnWw8Zr/vLDuvuCCgxaRnuterBTzLFTNLyEfQHpEENT8AIHcpjoGGmY9SNrbpho
hC2zpLpgl/rw3gihzeogp76U27vYDf26ShGeeM6nUri5HkQZl2gOQd7lz5H6yXDl
m9ccdCEqDU0GXEgoGkPdM+PbPX9iF896513YUClUiGmyvMEmZJDVInD/VAciUMTe
9g6lQiEQEhP7n/qa4f+EIRt3mvna1PLQSUHda5Pi1S6HPN6izQxsjVfmUXD+w6fl
u7cMmAmTbOAeBZl0IMewJNk6nJIdv5X30fm56aYNvYKD6eQobie/E84iVmJyhmM+
IviEBNKBGXSRx/E1VxFLdVWNMa4uTkL7noCtT/Qv+/fUb/V4+fJW803Ps5B6C6bP
INiDtKo/9JEwsdkKICOgeONS7lVRsxNh9hhmvxJUOPBvNXwjf1KZZarjA7qBL9NA
sLz0v8HFPG8jUd5OMcN7NurXyswD1x4+UGIpNLTKyY0RpYNkl4zYj677zSa3B0aH
PQzJnDToNuXEtpU5C+00pxIFNcR9mjKh9pq8LK07EOjOgfmLpT+7MiC4XQXjI3nc
8uHgnanxVCokhV7f4U8tfWO9J23xtiCjx/RaOgsIajYB/w43rXBLO30lTqTuxzQ8
m7o7Hy0LXQs6jbcEOWKTsyPpnLMoQKMIcTJ/kE5oObSV9gY+AQPECqv32LqO5x/K
pTWCvwiddgbQHeiY1ReT0IL7X/E5a/eR0lFz0UJXwEpv3/TRPBlOLVx0vRuJWgC0
bgYmtjXBc9ebde042VuxsrprJOCmVKWt+O4eJVyHTfYZ/Xg/QG6FBa+jigxY3PR6
7jl9dpx/bR2QpcylJKWDsJldD8bd/dm6VoMsR3aauugPBLqtBZ/4bTTl0taQQz+E
yynpOrFBbhJaKkhsx8sYbi2yoxA1RG5Q619FeCadhnjkb7ynikGBRKISSL/4jf4u
dBs1LiGo9uGeau3xJHnuoIrLSORCxs+AajHcWxLtuHGqeaRqGuQlIV0Z29xoyBE6
bdsjLNuG7lW0Mxf9OIuKescVDtbClR1UJoDs29vE+beBZW0tkILwMU9HSOSYsOAi
nG0vMdVr7MWSstRYs/Y1aFaXqDvAfn3bDb2ZVE5gOSRk3QTM91O6BrO7mRjKpF0C
Giyq+DH+RXbgSujCWirQYF2Y2bLyy4juFhAsXD3Q/Ytz/p2ZSufJW0pPSh7Y3Qs2
/ZVJpclsR14h4zqa/sMs/ltum04Yjkwua14vPDtIft+9JugpKftnJkzj9W542qDZ
DI5pv0zofjlYh3+MIS567esR/Bl3j7LX5dQZu+gEFRBkn1Ay+TiHKwTK9Vfa00Rn
xCRTdB/ZnOVw1B6TgWhMljUqYFhgcAQZjWX4hcGkqomQdMTAwutBINtWusYH94zr
KxW5CoRbM4XyL3zlAhsZ9y9aJt96FMuN7M1cCio4AtEVpwkNdCc9PT2dyVSGXL1O
FsxGn7nSZPImawpuCxcjQxDSEjlW4aNOak0Ya3ZTkZNUbp7z+ZHs+mTYtY+ZZVYP
a+4BFfI/55XaczilRZ/cG26HUB/swBYPr0f8B/jHIiTcvAzy4hFAlQrDM9mJfNfz
cWQGBUUuzqwGCFmLd8yvODKE+nkyqi5vTWDaKVQ+w8OnjjpGIZ7w8S7w4mkJetLP
BTa2V/0TSxIl6gHiU4KkX00xx7UbKtrePYNJCIINul2+Bobm37P1PXNWsyRdxn3m
ieXYQsCAQliSU8ojel3VaYhN3ijaP5RIcFSgXF8MgsLk8TZJkLJhh04oZJMupLXl
ggJ69LRsVVpzTggJ3w6OU3OnKQiQ+IRSScGVMGeRoe2Rzr4hx2v9eGGvMWdiDydh
sAcHVl5O1qaR2mrrfHHLfoI6HRbYjoHF20os0eWiiNt9i4Jou+BoWhDB17ioDXaA
JYn1V/h0vKWD1R84jKtsJgEIdRkMR4oSxHKuqqIuTmwEgCiu/ubMx1uS7GCg0uqv
w3Bg6p/TI+tMr1bKudViNsUDLIy18djkwlkaQ4RyCjrvQMfUKAV96gtJp8fuAjIl
KZ5zT2MkMRYatDPSYyXZ7BpoA80g49K5cbhdQ9YJNxUzKpjYa7zAquJjD9PfTYUl
6NW5dHKK35pxejxau4AuFWuxkutb3m70JsIfwsHux4b58hk4PfyDkRnb+ZsIPBG8
fFLNrBy0A5xd2xBtTABQKRF4FzUMxMCAeSFjFB7xvLe1Tm69iDN2UvIriwJjuSBn
lRLUZ5mFjbjyQw66VWOXNpVvv5OmteM/oVTJ6U+tskCCJY6evEo5fq85YUj0RMxh
f45NLRSgVdZliCE25uxGP8SsbXP9UGt1J7WZDgyxakmFp5+geTegHu62V5n252b9
wgC3RaZVxxkH+JKoAD+cZqaFPZr5bMORnI3lojXfFtus48+x/FK1EUgPaAjEYANW
H66JKTBEYM4tnlfGie2jLj9fMUlndfkHSPqt8cMcJ/1UMHYgEXV9Z+DHB2UOMdk0
9QIiKtBRLkvETqr4yePCTSttxhkW/gtQ9Mq3L8IPZGm8UlbOcnafRqUQBhh140rC
TjZCYpW6RUG78YdmHsgUGLbsbNSprVG0Slxllm9XyKHmWGsnudUIDbcwOyUpdFjs
+0CHlKl0p2E6RFkH8buShjWDYHAx7nbOBD5sccWSx/rApsVaZoctDXmEu1djRReU
WgPWebiChRAeN5xaICey65Gag7bVnFGq66H8uyKBP4A2//0KgKf9rqFhylwhVFPO
Sk4PVX5L8/kNSmQa9IVQBG6tyjqBsJiRHxK0m5H5SYZ2tD7slV5rKhOEL8MgUyqJ
rkOYbDq7m+KY9eOaI1vvN1ZPG2exh3yXAgxr5+RoLwi4vbtkWPeNXofJOiXIL+qe
36PLfis3O6R47X5Tbt/n9aZA63vL4Hqp2NkVjYmdQPJ0V1iQ4Oywvvo81xnXGb2i
98T7vbmEoXpWsaOi+vaUqLaRzMG7Vxmd01+sFllqjh9mN6R9obIJwR4pSQHXdbyn
q2v9ov9xbJTC5O6zIpwYQgi5R6KG+2NtpFr4q86ADE9vPPORSdmMg3R1s6qnogwO
KNGGMp16U0iWgvMj0svznpcFUs5KFl60dnVIT6uH7tmK25juh6/ifW6R3gq1ryNU
MyImXXNTLsNwGSCuzN4n3TiyBcTZqrhsuiDqXgKC9OlAkGviuMD16C2vh42rGzwX
pO3Dk1fp/9Qxi/cY1F92k+wOU5gJcuvKMbZbc0WcLiNswz0uPKjSq8yJ/6/kBzTM
c+DJJB7vQj82WpHV25P1+aFgTHDtKKImKtNjINuQSnkT5LykDVprbi5GsSkjkIel
w9VMEW2tuGx5S26a7nIQLLUObNkElLQNAo2qxjg17Wk+CKdRDwyMItKNDk26IAgp
ivqElZiWWVSrcIqDbHCdCVTVJBI/K8KTkSlbVopDXN2lpisTtmIju2qA5qAYl/GD
p+QBxhuAaHPGbxpZqJSaGjqT3BFiYwT4YgiXMnwY2Z8ISO42k/kBSaTA4T0FTIBK
1wBOHdGK7KuaYm12/AOdjhTAKkkU/ehOHPuZePXZwEhD4TFvGE508FRwg3gZlpbR
fzcoCC2BpOug5wFdjD2awRbAMurwO7JWeQnPijNWK/BYzGyjWB5UC7SXUHwnrI94
80V20uwy9kCbzuL/eAJxTbdzJ89DNpy3ITtpaLPDMKlDtTnjUBQf+KIiZcKJhgCS
+Q5mqaN2oGBheYPE0nQgdVdbkS7wgKY24Rs9+n5QACsLMwTeeY7Hmy642nUJ03A1
nFFucf79D1hQ6kOWSaAlTOHM+uvDvQusWjahvWS58GLB3KZ2m8APOtoGcxe+fmcq
UUMRQWlp+9gwNDpdIkS09DFW8tUJj2Q/wsCH1KDaB+H7wD0+jx2dSvzwD/bUowTs
KfBjVNNu36A5RrCZ9gSfNan3Bcvfgg5uBglqz9aZpDIbF5TaNUIDO2uIewt2YVy0
uIJAWDE6SAvAT090nvw/K2tcwwfnpjiqgN7glmnwv2u8wAAsep4BPh0UjvwFrCZl
VV0VSChW5q/3PIu7Sf2mLPMM/GK3TvRsBPwDVOX2UUzFaL1qV7QgRTpYSgjyqEq8
vVTo6XbqG4Nk7vm6wg2ABEBsogxBVleEGTOVDGIQKA71wXPI4UlkG5UAVDaK5xpz
snOReSOc38gzsm7HATWzw8gQpeSX/V2BwXXYnLMMr3dpicavxE8ad+7CyRlgMeT8
npt68jX7MBAgTA57C3Yz5WdjqUh4WASS3OFNf+vfuAA/XfToHPvgXAoUduAiC/XL
uiiaqIlC1/S8kmGPCOVXfzVWS+EMrkM4NI8aqX/zVqO7b1q8Ju1rYSXjok52fPgl
QZEJvN3gZc8mMocuaGCrt79f6TyXHWDCT8GBaJgFebHVKil0VpfvuK5HftPpeqlL
yYK6ukhX2LECBeX3fEr+1vRmWoIqaVjsyQNzmQWMg9SdN8iggvuUsTVqBVCW6tKi
mdjeeQGkGUM6wcETr/mVaf3lf8ClPAyj6i9xtRCbZ0MZocHkv2mLAz3koGHYeWGJ
x7UnL5GVXWJQcfBSFB1fzssPGExmsDuky63p/j/vQlLVWovhNCwtyIA9YHsuIEAk
w8oO6929p1wGEJ+3Vb13BlRRSXJWKn+I0LfArT755JRs/JazgH0Wt77Cz5ISWYs0
r680SeXpJKC6NOkRn95DEtOCtEbiTP1shooR1vkt/gY3Cl9xOSZtnZWcBjulhGTJ
8ISq22n5xVFg3K0vCWu3bO2/BtZ+/DRYd6giHeZF22WJTRyFdBMLXpsgb2gjvVBU
6rKQTj1b5D1kEd7qLDkvKYbU2zidbNl+SC8BMGhR8SnL/Jq20TSpNG2oARWeY81l
bhUFNL5gvFbb6dC/dk3OoDRKRkx8PBkRn/9MPLc75jVLjQITo7MG/imbNZlIeLp6
4vvpddUqFF0CooKdazM98kAU6xMT79bMIaXwwpAp9NsfEP2+YDa5H8qCTR8ZsGcw
xq6g8QyPp2UHetAiuyqDOgwyKBHcc9tWlV+1YOmP9g7R/VBn65bBlX/jfd+BCzVp
i/ar7p8/3kwO2hvda73JLI0wZULUA6VtHb7SH4tpliosfthZDQcEG0MV80aZ6RQV
8xbBt+c5PaNVWh1SzuB85HLWh2VIDHYLgrSgf+qTWqHNz83uNtgffA0S6YVbKUu6
E+AY1tRg7DUEGSvF6ujeeZvWt4MTl1Q5iFBnaJQRin/Rqy0dQMYBX3KBSDQa4qyB
1py1mKAhfpkopCHuik03+VXdOOHc4IiE7+oMMzX9fNxXRrmhZe9Nus4M6THU1Sbr
yqIJJQ1O0ujvjYLfrR9PMYaVoozzJaOO8NQhqW/bgM4yZc7KapKBZUPECZs75DgM
Nyuj2bRep8tnlXtF8XEetbTfTSILwWyfYrUS8DCTpU4+BABJgjPViWuoNuCdwK3B
KMu0wSwtNqf+WOaPPUUKCvUqQb7DhZK6l034zYxumi9UtRnDym3R4XbRtYtKAy64
Ae2AsFjU0dCcf0Gxv4swhM4OyrrgaNgzGyXxiv+wJmAkUcoM9yK3DO6ZgReTd1nw
gZ04LiHgzevZDWN6ZPcfkz+ZyuhvPpY+7ss5ptonjSfBrU+JMXa6kOFXt4L9TTys
T847PUoYtP8kRO1+YAtbqkL6Vw3Mfos+xM5sh6O144Ppm8I+sd8r7YrglMO15Qlz
NxdSrqzoSJRVTXYp7Hu4q31ETL53hNP9lA9TWSrRkNOX1/8aAM3Jv6T3GWuFsxv7
/f0arnMmfK2ZnfOtpxZ685BITw+31bo1tpLgYwy2XbZLcIRI2+LStL0xr6witLb4
FnClOELdExREweEMUKkCAGH9fuvpjJwsUVgjAHUGEiRvLBKlGJYD9mCewfzusrrf
aO7EojfFwyamK4oIOhyVgoJMeDhQL2HW32n6CrXJ5A+VEAcpmsQlK8ttrV5T55oT
TJTdJrWJaGCcJP3YUcUJ65BmPk1Hv7zQ/tcLeYwruezK1iSojk25no4K4dZ97177
wNiSq4gk0jrHfpEvvn2bkD+ss+wZg1WTJ5/WhoAlIoxUDU3kMYzIy6vB86RICsHz
5JnLv3uwvmrc1wr+S1wnxwzdc4IEnm6Si5P7+XmjJ8LtQro0ST1NOQBr/g5Y81Fw
7wTVqAeAtTtSzhgc4tDO/PNChOw8SrSY5IdcCKcpDTyiDYaiCWkqh1Y4XsnENaHV
32PJJjQ/03vhFwoDti6WyCJ7rg1Ip7YFwYjhuudw15XzsVUIVe6DENIiPnSHgHrS
BKORvik2foj3/zSYEuoQGCklgJF7GjSVYkRxpDs/xDUYryIIT7Biq/wtd/Vuaqlf
K+4S1bE0pqdT0HSj0D6HSgr51zzGJJ83zKFhfKn5ZVy04w4IN4jEDSwhLtu3xCa9
EZXzlDOEgI5zq7Yvk6CRGVzKng20AdhSlZzl+SeRw2b6BTT8lMVi1vJ4J0zK6Vgo
bvNm8Sp+xsOv3ATfd0EXEeV4djLKhIUhZDWhJc4ddbYGCV8cCyFMzWlLGJ4l153o
3A62AevIGVaw/fvd5eWOCC4RTNo049IsrrvcY6GU7oPduman14doNWV4Ec8Wf8z7
YNg88q2Nl1wYC5I56T2uF0WXOfhOmBM504hqI2cKo8yZCsScjOjTPEzN5s74LEbd
fxa88MwORAn8WTbjoP2Hqc0XLBEfa6QBr4z+5U48Xn5yBIPvzGJRbR3czBhfy4pa
7lnjfvutQTSiWZAAo+syWThq+jxPHQz+myHPbInH+alzeY8VGwBroqy6mDhrZi5l
IrmXEg4OvlDH4nZdHqmy+N7k1IsXoNslPDvOQ64+tey//kNHltICu5DVghWD1hg8
esCVT2GUdVPc+4FH9r09Zn92wR9EtrKG1drMB1l4IUNIBYXoIHQHDTuxzC58R4W1
TwtG3WU7OMn4fnwCW7qznGtNFJrS5qwKd7HkdSMMNOqPcSEI0eqoYCzkFkv4ncoU
podv1HqH9X0LYD0o25jmxLJJDDwwh/bBBcY+AXBsB7MhjWtQ879U1cwuR0KYfWY9
/skvMXmr0LJrWByToKtTDF3NFcEzOhM52/M1S03hnxTIm/nBKzo6KR1thU/MpFco
w3reJ3UOxlHNWJ30NkkhGwXC1VVou5UumYUXGjb51aWT2Gvc0Kxyqbhiclm26p5m
o83CBvErWvAjmHuCEGAOaeIIUJEK6kky0MgmIBn2U7jKVyd2+ugMfsDEhROnNiLf
dUeiIhT1DZRW/KAG9/jkQDPbpA23UFNkAN+OdSokbA8xZoxUNzgfzWhP6POts5cR
3Xnbbl0NdoszyUoLvY2OEMDl4QKk4i0dnZwytTADTQrEzoUSaKLKt8/FBCdlLCle
hNw/VRhbBweUbPwTNULp5unEPNoU9T4SJ6brvOwa25MzweBZ/v00wVNFUfQIsLuu
+bjrJLzKoiNJ1cRnjLpSZB30CxaTfxNrV60hGmMS9JbtRooPMtb9nIxCUAue0Zfu
vxm+nBnMV7p5SFqvodVepvKKFtdPOeMeFyT4Bdat4RWfPV9vNwIxzT5JiyhSiHM9
xy5skiIjXaqomYD8A1/12H0v1bomFq4RfoQUwaxv7Kam/2wgr4uO4/bPz77L45F9
4EDyWzHIlylN9OCvweOBf08AtiDcI5388+jyi5P/lZiCZDY8hCktvS3RsONNDX7l
CMPws8ABS8uOpUkrENm/5o0EuzNKeM4vhJDy8ooOW6aTir80cLHSLbK06ugHFD4o
wQZF2BXFmFgKk/dl7VDBmgtfnHYYzRsKL1r9ylm84i3DB6IApyjDh1xOzIhYctOC
WLjFZtaHiERDQT1EkUx1MItMUcSvOqZJgwCVlb34TPUI8CPiAsGJ/yug5kR3Dnbi
BuhngxneZRRbTRl2xei7Qai/DBelETWqCSVrWl5xogCh6gGQRpF72DIlhxLG/Y+4
QmWfmVB5aJ0wshNgpVoI4//L/qmJNWvmtB7ekxmKyqidxFwIoE0A1Oyx+ayVRZYF
1KTk0R4U2NeHMDVBCLZ53I2YJUabDCWxxHqoWB9NP8FESQGXQcEZJbB/MtdDoUuM
q5UgU2je8ORvCeaycUgZ6gkXPc60utdmm+hvIJe/xhhvSIC1OLMWibsDkeM88K4R
cZsqyRUDDLAjaYgb/fOqQwqdSt6s1+WQz+TjfpwnrXQdMNpR9uukoF/efkkVuUY0
kvwlJH6pZqe9oUpSTbD9zEVopdkFfVm7F+lrz2L8usntvRN0wZpb+PNdTyIZ6hAd
IbFZAJZ2y8EREYDaO07JWiO4mTawH9NtJSrBrlYt9ZeTIVs35VK+6Z1yMGyIHKOC
FMJ1d4XliQx8B+0Xe3vdGdhdfnCZP6Uy+79qzm3loDp3OUX89v3B9TSWPKfpEmuY
RUOv12fzgqH9RY7IQAmOWe3mXhbetdrUmhdxTOluWvAw2920mtXInB9nGURcdeJD
VHGZ75ZIj5uRTqxh4FwON23m6hPjJynqjF+JZnf1OBV6uIQbR9EXLok2M5AIY7mI
uh1lY/SReWN5yfRLMdmbXYJof4p36fYmY5XfckHK60bHlvNBC85v1tEZMXL3+9Fb
GtzyCgp4KnxlKOP0c862AjzxWkNmDQbD7GoFBkC0SQbr3itlC8iVCbuzYfSTJrqU
9VMgNIqdUVzTM3FDCa6qGOQeNvQy/OKncFKuM4WOI3IL2MST2YbTeIupxfKO6eQC
OeJMF11I/CJ0FZTgkm7q9S+1xXLC5mo7uxlJPS9Ccw+XhVMHFbEuP6tlGP29+YXH
HRlis90Ax06T6CSzfVzNqcXHQTSGvrKqIUL/rnsbdvM3qu/Zzh9Gdi3stdYGFpbq
sfrgLjhCFx03ZVIbcx5k+qzN6KBs+gRvgYfC2S9vtIRmkq3eCN6R/FMIjZ41pS/I
c21pO3oSegppt8gP1Pb56pyglj4v5mhk3fg9d5rLu3e5NXJ4uG101iEJ0T5I4rdW
s8W9qk8WGNrRr0/eUeVEW1mPgmyzSMy8XZ4czJTMz4rFKtS9vgIx1kuaPqM8edRR
wgoZeIshqwmzQErusVKtgrZg7RV/B9TkY+kwsFf43t9YYc8iD18oAyZG6YiQ5YbW
2ruLfX5S5cqso8dVK8S1yc2T88oyPvgwa6chyD8stwdWvXp9bG3nSAbtjsbRYqP7
`protect END_PROTECTED
