`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V/xiIiB/BSrwy1zc+v6PGkONfoVxqk+JBx+7SV6j//jkVjXHkZSz52IuM85mgB+W
M1+RJp4J2XIkOGnFBXcRKiugEWNSh6NSHIPC+i7VL6Qc6TH8Bl1sZsdkrx5OqZRj
ybhFo2MWM+zvq2lyMifVMrI9rbN3TIVwzSDn5xjZIQtmdx1PfAZDzPeutIKvikFa
O3MP/M7a39RclEO0exiNdOVNrBgMY49jS4qzNanVihLTSGNhrFrfgGN2S9TyVnCe
mbjbjWyk8gXTdgo3ZGQAlG5fE1VH7YmYphiOJchYVJrSWEnjnFNqZgT0Ow73M5PP
bIz1Jai8ASbwqz71ejZwRw==
`protect END_PROTECTED
