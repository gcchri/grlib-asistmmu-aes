`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qXDC17dxSODbIXuJebF/irSvk7MSjU4hfDpvG023OTDC1RnAKSpS7v9SAHGC1J9H
nkhFfVDT9bFgfdNuY0ad4Z1AfT8XFWgBsz72GViIOBvbt1PgJu8Wrewk/E6fRrac
Se28jmZnZX4KRgYXk4zSEZ9I72Up9kFCCEocrYmAjS74y47t4w8f6nRmN4fzjFCv
8hHFVyXvE+CaD+Ict0aar2JFoFtStzZUxUvBUR1NdEkJ7oQEE0odAuPParChmEL9
AaN62MRRcP7PYXzt0/zGNEDce+WOTVXhNwEuNiu90VZCLq2on7aXNHguX/yRhJsT
IsihPcFAeswA0ZaJDjo4DIkiN7BXtIPR6o6Vxmp/81/CCAMlrG4gMZ5dYiCW9pD1
7swltMAXg07dE0/AJBhU3VDoq/dg+60dbb81c0Z3qE+34FUqyd7ezYayG2dbvxqG
kFvjwMQy2i1ZZhaPA34eALdVH/u2zzmpTwcLF53n2onV/SDj7RzjvGSlg/7PB4yn
`protect END_PROTECTED
