`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mG9nfYbAbsn3HD35KccukI4F8BU7fAFjqL0xiA/xkz6ZFdqonGyH10u8+f4RfSI1
N8Y4BEpcCZ9JYL9AlZGk7pmMfuhEY73kEu/efv6h3rpGxfZI5vjZaJqpMyE4HHdf
wvM9RJDHUnmnccrb1QGvQAzbuyJBzFs7XXk5aHlvm3l8lM3890LVetJQlTQ219AF
F2ez4U0/W1bCikbq2U6Gud65+L9Kr3RNExwXKnnGk11uN466gyPStH+gxY/YjYWA
QBS847zYC4rLBjdkE6aD8xgVxIY/k2plX6JM/FVu8uPgX/rXQOB9HWXJxMxsRSIT
bv8oiCxJMpX8cRuzwBUURU61Q/pHDTNi22Nqgfumk51A2nP4tJdIBd8kUvD47l5t
chdLjFD02a58spm3liAVSnJmIyZaks0cGtRhftCGNDk=
`protect END_PROTECTED
