`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hTcpdZqhryoJjEKsp3ySWYCdzy4ZVgDjzds54XtHd35oS5tk3L4mq4Cry108CBDF
y9yDhkTX0Jg4qfm8sJPPM0t1PRPP0p2RMMv4ng92p00goj4WfUIMXtVW/9JlQH1P
aI/Wx573Y5j4eBSLcX0wnzSieg0AjbTO+nxaCjEW3w1Auccc23ttpn8kUoqkEfb+
03K+EcT6q6KIzhEwH2S19qaWym9A/M9VEdzcr6i3441Z0R+QCqcnaGBLDJVOX0/M
0HVDdTOv5xy8rlpXOrJlSYrSYsGYxNQRXbz+S8jyh6+rQOVAwUICfPY9y/YAYYKK
+Q/iu0NBUnrEOt78e6lRjYykzfUPQdTKDpf6vsfbhluHIMZObNDO6ZaWUl4Fs3eH
`protect END_PROTECTED
