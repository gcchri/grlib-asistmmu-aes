`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x1i3LqT84jLT6qR09+18b+daEpOcaisUpdJPUd4Srn06UT91l5esZm2YXXFAsECI
fDhC7NOmQkVOJBES+XmxoonixqHhxEMEm24Fc3TUh70LLRgR63a8369gcAp6cpPI
5fXq1EP8muIvC0IKD20un06w4XQ8eUoooFqSwIpINdxw+UQPIrZN+JiZM12AGs0+
h8fUY/NfOZUKehZiUGDk1QWbks38Zi2gqriH9VbqZ4tHTpQWU+XBatH1nLrxDBSX
r2UlD38JTeMeuu3BTf/tNggfIemx9vQgIIF1LzhPvit7eoGcyBYzSKzXY0y2+ItS
JWbzSx9n7xbNZ+h3E8LYIIhkEgEo8C5lpKskHTk6kSIYdd5aOQ55A0x9fy5XqmPP
Khy2LtkumK3+B4FbjgKlO+IlY7xmPMx+KNU0J5i+r/wq8Ai+xPFwSDTRmQkx4562
9hTHYADJ0JEURqpCdMEgVfGCnXDJmgod13jHbg85MLqiBlRKhA/SJWOqCiYZYeA/
kNruHTQRO/sbKFMMiZzBYRPdC6BTK1FWR3Nx4P+j18K0U2A99HXwwhwpwGAL1e4r
9nY8zqh6ewOzEIIgDQnjbGsDyN+gTu3VWo3rGKGF9vUXTmUW9k2BrYz/kQ3GlDha
R+qOo+WQ8s36H4jwlHcX77ttXrjX6wff8TIvn7Jb8VZhZHptTdm4Jf3jsm/Klh9M
fHszTQMjJOvtvasSrr1i36RcFj+NsQ5vVI+oWBx3Wmelz2b5eNGMyjW9O/ZjhgA/
Dz5fbo8PN+VUNckz5a291Zucrwy7yNnPDtb01j5JrI125lPCqFiV8/WuzDfuSR4z
zQFd1/V0x+ZEF97OcOWAXzg2FGEEn0hwnjm36RWMEbeu+r+rNbQQYkomGdHf6HkQ
kF26Ifsvee3ybsjry/b9WbyGfeGTjT58CpydZ3mnvxaLN/SsEQrikPfg3upejQsq
EQGp57sisTHPs8b7LSXyXVCIXc3udUHWbw4FPR6z8Ozd8NYCL8sbZFZptexQr/H6
hvZxKp87b8MQSEkPbhiL1oRHyfdVYz4W2fXLc2ujgpIPB2ZhCnJryfCuqix69wR9
rlxGCxbUKNU7g6hGAvqF8D2J3qawQVt5H2ylwu7VofaCjLeBytGj7DY32Ae5J9of
eusphS358iZ+Q/yQRTVpOuRoojrNvsaNv9YDrlDS50wqkWo7QSvtCK9OLAA46rfY
toUWRuAni1wFFqz64y8OZv8xE6U6OK2PRLRdanqYt0E+brIYnlgvHRcuwGZrY0gW
rz3P7C1k0RkWhuKFc7jUHSkMBaYJqY+1uqLKp/Q2Wi68j6kHCSCOU1Fdeqf6getn
8/1I4g4QtiSAb+K64rJ1IIkF1ihuylGJPJLGZRWbh0/WkpeaYYMz9NYgOGcaKpBq
W18sWkzyDmZFzcbndcO44np4K4YGK1NFnq/fRLRmD9KKlnj3BM0qD/4IAxRGFp6r
plgABT2BMrLhd092BMvxsUEa3ds7ilfzhoPtMETuN2wbZpyGJHTvOPu1pS/JMOPE
Qm80ptxeHFGXM0V+23NZ0nb776PC0PQRW4k69ZJtGcAigUggA4aL7nYDpC267+no
UM2ZFu79ucBaF49i98qf+1HNzsx7T1EBc6raTN3GN2LdlzUoF/HDTrdAdzK3TOvS
SAjBEptvdCfZFT0Lo+WBGIt7E+1WTqtDHN+qKamye1sdK98qRy3SlbKfQYkx9Vq4
2qp0jNVxWSr3CQF3qF5qcADlZlXAVNGGaE9xB7ridLmIqhopa/pIOkXQlfMqNNGD
+xuX/17UaoqIXn0YcUQmO4oq9qVykp178s9K/Zm9VA7SXwdDmkFZ4LIoL5U1L1O9
AFQEPqiRemoo1L4jrQhKhNXYWde0mfs7lce+uunTfiuDsrIfPA4BIgSKOXUwlaok
L0vJd7ZlKxxJ7MQSuXMyEiKqPVnbgpZgeW5Kh56mdk5xCw1F/U1HOZBd0dfTkpJu
06UOUgp0hERfMrfp17EgWYGOzJ9OTZyUfVLqyFJFe5f/n71156KtJBX9D+/MMLng
iQcZKj/oa9yvqGywceAb1HNZOR5RlmktihP75tpinYV9H0VGg0WrET+dfLqPAOu2
ZXbiu1D9HxSq+hVQIFko2d2bDDcYEeM00oXSU7siFxUq/Azf+/s58pWJ8sF/mXlR
DrJxgDWCWpxAMtElKbimnNLVtXAX0Lsgs4Mk6BQ902020N2MpN0XR9BaGzRr/o8b
DfvmkDQtD/iDTf3Ed6Urso9urYghP3m3ounmzZcmnR2kMoR/AN/rFspvNEVICDhr
eo/gzmHV79HBPPXVcGeTCDip4LSUK3gixMSrs8Gt+t9Eupx9uJ8cwQWEZsS18bsN
M9XZtf4ZVlYQG5L9zbr9cDh0FpLa86F6+FnPoM6VIhW/bWvbGAarlq1piPyJZnpy
tMNQvxBynqfyEpYoHYSqAYlJsAaLqJJOquh98tZFnBcvLPz8KHQOyVOrDRb3Qcnm
oIqhii2QXmZPlu4Wxu3HvUZG2bgQoIVnWZLuT3MnneudgqQ6t0VPrZW+NvnklQws
wG4MTzOKXSlG/TgQjp0zX1dVjjNOwd4J4eDT5nMf4uW3HsNI6XZj2BnGh6FiUGxN
LB135136MLDlCwP/pDNpyQGt7ic2BMbYknUrKkdZJm69tA1AV7gnTsIRYydWBOWW
`protect END_PROTECTED
