`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qx8WCnIdbcjrlUlAmLLkqD+rcijRPbQ+Jfj85/EifdlatWLO+iEhLl1XboiBzpPJ
RPomdzf4mQjGdi1DwEu2GEIT81xdg8e32SmYkBYO+vU/Jxl/+knnLIz3skAUfnMD
0NDL1y3EhfUaTTCZwdzb9QyWadtSv/uf+LQLOOA5iiZvr8NyR8BT+3AU7clzLyAK
RN37GU2rb7+9gCEZvdTbaifTNShxyrlam+QfozoYi8ob0IeinlHVeLegdvw+yqVC
VGt5xqFsh0St5+rPEIWmGTmACFJuqlwd+F0S0/0GpvAKRa8IWm4caBSZ4WvKJreo
JVnIvflZXLQQFtD2PEr9lHr9BZxrZ8rFjr78nN2fwIRUJhGMeshJO4NBDh7XLsei
4PXPHy1T6Hqzd6KyYy0hVceGor0cxLJ7ozWj3eM8PmkC1E9/CzmtiqMLbVOMfo2/
rtPl/Dd+nJxD1gAEG+RtuMP4ehblEVml49csHN2zguq0lT4w/HMxOgwDhFAI3Bt4
eWUGFc9LThH7NAR7n0KKtYmsaKjty0mYWrNXHvdyHfHweJcIFkHDmrRmDvFBwaZ/
6wCAUsCUl7AT4ZZYunU2Q/VKO+7l2t6r05FchCSU8a8UQItLirzEZh3DP5oyGV/H
dBtXPtUEX3y2trgibccA3/eyNwSNr7YHxqQHl87Cp2DXMiqBigtWUOXjflty53qm
BRkCBO3b7ODf/Rs95mtWSw==
`protect END_PROTECTED
