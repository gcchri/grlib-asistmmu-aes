`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mSPfK13cVrmhEr1yQcusbbDYsDdwVbWKamOSrAR5U0ocvpVvkbtfLqQtjzZX/afe
nzJeoGJUI5A4UFGH16v0GvJwBBRTcRZfRLYHu9i5AIL5+Ij9GbMuao+T2K4dY76f
FJe1THrj0PSdBPVsCGhD8infyn7zSvXg7CvJzJ/UF+D6s43BahpM9VyecsS8HAtz
WicVXqlRMsVDsxdJReDuojRvKXp+T0Wq/vF8Rn9vD4zeM5yg9uqL7pjM0Oj/lR37
c4oPKG+j4Nur6c4D5ZJD6aUrhr5xsOS+9rmV5e9FMUK9csw0bLFurobPUXuHgokT
bZev8TEywmf2Wwuf7s30/A==
`protect END_PROTECTED
