`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aGOOCvXiidoGOQwf/s14L7yMjPryNW8WHnS+1XOp0Q+hVLDTBv8psrNtlU6Mj8zn
sPUt2GChw4eS2OSn0p6teda+1j6dRxYx2tiTFaZFFwMJ3llhbeWMlcWfkeOCkkgr
2eQhn+iqC547yRCf7q29Gvdtrhu1V/gCvkJVNboky1ZdUp1u8YP9QQkTzHXe/XnY
5eqB6uFILZlaz6Mu9EzqgAgiH0VD27JGkQZp9KObm6lnlPpSFb4qdJeTDzIOqIgD
j5OdfqJrfv8c7nj0Jdeslr+cU+Mkllqss7xlYmDDO7CbTNL7HlshNw4T5Y0JMjCf
Rrr2NjkruhGuTJnGS/9Z6mokMu7ZJX6oTYMYjNa+aCmalNXID3Zgfc9FSWRP0H0t
3JWpVx+SYCmlfDevs/FNJRMrKoJfSO9YV3W02IftZvYK+JOVDQFxqAkbIORC00h4
PKHEnLs6WogJDC0Qa2DhDosI2OD9A30kOKgLcN0G2gik7bs9L/JGS+HUtURaT3tM
AN/rCOooa2QNTgpfA2U3/OOWf3lS93aBH/EB6TMotC7TTFR2VN9XIFSM2RNZXINF
8jp8D7BRNx4mqmcmeicNvOXZxMwWAE9nkRE8+HBzJjU5xyu2NyXT1p+yyTJI8cwB
FSEnyzkszucB2AeTfJMtl/fT9/1Z4MSDDLw0fQzvKB/3lWM8kLu2pthaCD95wBd0
X5F25Fb15118P+nf6S5qZkCHbYNn1W8e3g9M2zqw2+I=
`protect END_PROTECTED
