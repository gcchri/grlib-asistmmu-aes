`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Paj0gTYVtXMRpus7vra87mkQKSQVjOa+dVOG4S12B2DA6lybedEUZahfRbXAntU4
bOhQ1ZelYZhScuG1P+27hpGUsoUq3zIOgSYiJzrOC0dyJS46V0hMvQ/mGLyTxd5y
jTUnJRKKQKBeYAKE1dO8VydvmB6EjdnEu7hqQd0yDKxAV6V/hq+VIblq0t+f9rEH
CwJMfJ+ZsT7bpSL81sWwbTD5+5yJcUOVwb5IK9OkR5qleqqA8dqPz6IUwqZ5ov5G
pIzNx3YcNQNDV9iFfEPWTaIBYS5D6h4UqC+wJevWsFnHTOUeX8nUdsmN6Gn5MvgH
5wBwG0c3+wbFqMYXEH9otYQs+PArq2ZgtElAbNoV02/hlSCXy/QpVmn5y0g5FaCO
5UqHlTKngCTyRvyH/dVUAeM89PssZcVPm+3EBtKWEMDKzS8fmyOZ7Mk4GvT6liZ8
PyeSVYQMZKuv5JOX2e86KGfBhz8z4zFCmX60FCa9xCL5mfW5Te2w9pngIqmaqDKH
Ta4/6xhmCnmf2UZRG9ld5yzOMkuoQ7gXDyJp7iV3z+rVEXA/VoJx45DXT81TqvRm
REcxMuxNUH0earhyCyEmdXLL9IVLTPUB6Jd926Kw73kiBuV/XXV8dHY5QpHBysrl
ETd3NFdFPp7xxstpWFS+ojxGANNWJlj4tn3T8et4CS9DC9Rz7/JAhGOWJ4J2wnkd
4cCfjpwqriHq0HM4AYnGcugpiHdSWEwidWm8vyvyhkaKQv2YLkqv2bj+Z8Tv/Umb
UE1TIOe/LIMnjaakHECkJ6eCqrjHnHV/GL/XyzS5O9teiFbMSumv749PEsyiHAyn
b3ZFl8+DnaIyy4LnrTHaMrUYOd7pGNX9gIqoPrprrTu3xKGF559qZt6FnSlPbICh
pud3/eU8SPdv/ogT2bFO/T1CJQ4PY3RaTb+WqYriMXR4VH0gc05YMyiSpcqWvYYh
0P4iGD1IrLue0EsWeFe9xOVJuvXZJhzUV+NewLb4pb9/XBumr8vTpbqdYJEk0WS0
VrWmWesUprqkNa1KW9sCddcq1sFST/gCAJVUNzx30faDfQy+XLIBQ/rPe9fyV3iD
7h6wfgNiBMN3bAHWWejwB8G34ZpZYIdGsnL58OGXZc8xok1WGLmEKFfsbXlOHGgk
nU8wW5Emy5d4YqtZPE28Yn4eeTdCNaMs3VEdtIgGJwpSWleq6C93T+v2BZMH6Xyo
`protect END_PROTECTED
