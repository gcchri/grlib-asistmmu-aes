`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tUJa7d9JOdlozLNPnu/ibCsQyrf681uAxSs2CrVdzTrEtnoLLrz3+I5RcX/LPdAb
s9P8JIh+6e4Jt7/efC9mpBuwciba8gLD3GQh4g4aHPJvjS9oKYuFkpz2A/S7ygjk
XpDYHgBobUOxpZHsTxHmeZdIWziICATQ05yMWNySwhtfM2OCJw5t/nmMtUuAcSYJ
RIZeWOrBm5XmiMNe/hXQR8TIwb/c75goEMNu30ThvRL62lGid7QCTU0JCeApTXbC
diHjOF5jmQyMXoJZ3Csz7j8DJdZfUsdpgwuut6sVv87vzp+mRPsHxYyhTfImO/TV
`protect END_PROTECTED
