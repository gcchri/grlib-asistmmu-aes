`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FmTBOJpPY7Uoz9nXKum8LIZ9rEvCxtSVTXSAD2zgMR+6j2Zy6GH9pKTwcCoAXK60
ChsI698cQppzn+0b/NvT4NZLA8WUrijbC0xR0kYyLSnBnvtuuRM6MeAEy1nWuhIa
yGsjoZiTzxALLBMLBr8fBExC5TSBsiq+YehLnBCiNowjegAHc6nkX76QShDxZRiJ
t1HkC1SsH2tXJkaH7WT7KfcA04ZZ+27ipwU3+DMojVuLY3BtG1ssPJUDzBDp7j1x
cIrSwDWvZS0Tgm0gu7X6Y7AfcIg5V9mFvSPVl0PK0X+NihXn5vtLMeO5Bcb4TOl8
5aZlZPuBAlCVxVxI1zFg3/CXjCij+ptg5wmxJ7iu0D7KrnW0zgmvxOQBXARybreX
K0VgUL3LzDVDjn5ECg7UBpCjpYkI3ohOvgEMZ21OzgPjjGiQzV/Bz5V9QkelIgIo
qtbVqz41/kYH8zCzTg5H/1svCU16vpVHIq/n3YPOK/Xv3qL60DXABAMPdzW+Y3j9
3d02f1TUtqj3Y7jPm+4d3KSWKXiq88bv2lUKzuHT2e4FBQ8tEHOiPHlNPctpbk+i
LSgB6kQO8nAYl4ZY4PwGam3onhrDLNlnMTurJDBtEY1qW7D+yJhRMGfN5M8ILFJn
Mlmtlpma+8S0pJKLMi5FnJzHTBeyMBFCuhL783OUIvQ4vD4hwGIGt5W8s8gXk8X+
XzPa9Oub+timIDDB7ffW29I1uhzgYRI52QCq9cGjzXEwBAe67zmsppyR/bzXA7yZ
VhozWTi8K60A/s1Cvi7grkKcdfEEty3qkbglBn6zpkS1FfwcFxA8Vg4mclZBspgj
uZihNyDQsncGU2ZoqVcp/RXPCPZ8PvE9JBZ/46VOUhFXoA4YI1avfZBJ+4AoFkRl
D7ERZxoVpcIJLP7KuJBmM13WZw2T/y+KKc2sAlcWmhlWGbO+UmGfYZH4ChjUZuHI
WCyzt/kpYts+NY+LTltL9/Lm7dNCMbAFmK1RXnRGfvln5N7gQDV9YdTFRN3wUvcJ
HCT8WrAVWU+2jKpqnS1bKjDBqeq1Pz9/qu95TAH2wU5Czju9jkzwteG9yand5ewj
Gy9riio++tF5+DzrvHtgY9hfi+G9nvhsIS4Eon7t2LLYar7lw2yonXyZzCCYPvgB
Eo1uA2XoHvF5xzhbpeb8LWI6GgCmKkhkwpvmZh4EZhhGHgtqmBDAyHyyQ5J2MfYg
wDi4CqkzhCLvt9+wvzvma+wvzDCekG6+aNxJtmkrFL6aG1s08VNow5EMkNM0krfI
0/iB9CvCIpbrGNhsFAKbjLLbGhpy4fCNil6pK36+XXK2xmYNhK1Rr7qulfOXxzs4
ob9eblJqFn59sL1x/75G+tnxR5Th9nojlowQqAK/cKjEejRhluQ9QiALCQGM6pA2
CB3fsmzlYa4BwNXKngdUItZE6DRH0M9o4j063S1h0Bp9zWD7OroI6xXYYVENJhka
7LrmbmJlfM85JO7SPvpzisZYWJa+trqpFIVdsYMJlVVyS6jJutsoiDS9J0D2Klv5
oZCfuOe9zg4XJ+Be/91Q9QarH0Ng9me5axzFmO5jI7PF5/85ohmxgMCE8YXS74C2
+j0XwrphD5XuxO2MsHLASSelwI4dNBma3784XQHniT8cCImNWehosSm+33SenfTr
NiyLsUSa8rpgonyTH+Xh3shg75sNlrJnau2s4pdulR///pPWwRok3cxnQf/BNhp5
Cck5LY2F4Np9XXwQqOJ4XHltjDyUyQFAxDQknT1LU3AzkzJ+Bw6Xv5WrvHMci/3p
kjsB6fz+HsI4+WG6VSfZ5w87HLAk6C0f3ujzaKVvFnRYhKOZ/Vjxwl5EPZKcDcZi
cuSap/bM0WLOHiPTXZN0Ltjn6v2uCn5Ih7u4maEasxAxupglT0Izpla7f7nluwyR
pl7ZgGT5vhn/cv/QXTbFgB/mXQ837ydeWllK0G73gK6IpCIPYOWLnUl9ZrLJiB2R
2i+S5HqDTLo8L+T7XkCwyB3AJNLDsuMnOaZAhh8j55bIXAvtv28qO0obfQeneDPr
WfQbpt/vjQ/Ax5zwwt/XnQzsyU6WtSqz15isi3oAhEAOvJZRiXge2A29bA496Ph8
kt5hc34+t1HZa0SUPMSBAuXP/nWVpicXKeGQ2NHYaq9yo2iEFbx3jrY+IRo8H5WC
dBazSEaWsODWcPGnmZSuqqDn3wg4IQv6G8jtGNA6zVAWRYfAYzaKiMzsTzaKXZ1N
1bpJAo0Tx2d1Lf0b4JVX+lXwfLc3C0+zf2JCA14ZD1k19qkyJlnKyblUkBRcgIYb
Ru5Aa+y48y7BBHYsvc+yY6xI+FkXkWvGa1wWh8XeR+n3DYlozUSWsqi7JYMemruQ
MghXEN+Z8fn9SUwCvUE4UxIdik1+nvHHL5Qg/HOxRl0K+6+d0RXA3Ycp8UM8+4d6
4XagBh3gGtf/4J8LyiiHdpsHSuEfLrZnMeWjS2ceW2Dgb83+vfXTGNZmpuJRPeVT
uCpQNYJ+Jn0UySUzc08weoCC9uPGYJ5gu/B3ZtwbSiR4Ida8LdEgURB5T1P4qA9T
Aaq6BtsiMt2CIgNiBMN/091Dr7qcBCw76QSA4KAVuFTA/NeXYhFsm4surtHby1lK
uFOL2CagLIAH5xDR1qBeY8bSxFpnpEkGgGSoyRs5MUrpGq4A/pzQyONnb9L8ktLh
BjJQsRJLp/zj4KJKxAF8JlC7ICR07pU1LLQH5GjZ6+Wfh91ChPtLR5qY9DjhGp8c
VKSvbQmI3H9aDM76ktX5c9wlIwNyu6E7cLrpMssGM5MjrJLE0sqVaPjc+1p9ibFi
UUSPVvgrbsWwmHFpfqmUuw5bxfHhhB19J9vu7WUiSny9PGAT52Dpwvanf8XF7v/V
YGjDVfv3pK4/fM4/IO2qJxuL1iQQzlfjz8EWH2AJbQdEzMR9RgPgwwlfi6XGIk/H
QWXsYXDL+eOg1Y/kefkejjDysMbE4h4Y/H4OrfLeCw+8bLVxUXMJ6AYgKAsxDGgR
Ls6W7pbkSXy8SUvXkfrN/8L6vhqvf/ya10dGuGLGn/5b93IvjA/ynbn7FsVQUo5M
rSDwML9EXh3l6fo4cF8UN5Gm4lwCwpwifxqcEb/m/Dag0ca+UakvD3JqETimvYEY
IMB5ZCuphjYMD5n6XQiip7FwZBK0tbAw1LPaZuEq7+M=
`protect END_PROTECTED
