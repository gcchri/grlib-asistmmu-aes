`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0J386T+0GWy3l7CMTOlx568A6Nz27vX/sN0nMRwLjW2MT5gUQdfu29oQRWZnm8ul
OWMVbLBE2nGFEpzKMzO8CRR5kOGBpWcXchPymoMiYIPBiERLZPe0SZXVxeavs0nF
1qDcTe3azTj+6aQt+iOczyAwJEx3RadJhRNirHZ0duV44mzdHnXDGQS+XXuB0EXO
aJLe2iDYnkojGBEgKJ8dPgnvIVruHZkl8/dSzSb9DIzj8UsX4Jjq8Z5hGVz/izI5
aLbQm222YLav/LTho1W50MXTyE7shh0s0FIgL0TnP8GREynY/buiK3O2LRhyg8om
5dwNfVwzyTiE0nma0PNg545O6elrcAn7NfPRGMpz5YyR3oYPTF6NaXKKY7B4IYsM
KedRDwKohSCorK7xMZhsr3B0e8xMr6ZBRK7qEcds7KjDOSUoPXF71Q+4fZROqM3f
NGM2T/5Enn2Eg+d6JUyeI/ld09Ls4uvWsGIPtLHhvCTwpHTFnZzaXUNOH/aiuyp0
89oubgxaaIgo/Zw4lJpaSteH5fYs8JbzwfWsufgPX8bCbWOreiBWQOz4EHor+xDq
OtURIFnrwPvOcBoHaJLCvmzT4KhoFvU9nruXQIvlDUXmhR8szsvCrV87a9NZHsob
0/AElEwX6TceOtNy0pIca7FkFwnE7kgcjn5lbQf79ZTum/6Ed0V3gHR2ydf6R5YA
RL3FVR7kL4b237c2e98pwKpUwCHc7rBZRcS09zz/9srPemT0ihehsowAJ0BtUd0X
jMZldwTClXGFluhvd6i9scWoEcpwvO5JarGYRjEtJF3eel5tITs9XkKr1G9xmuOK
0dL9xwXivB0Jo6ZemL4xJztuKOkm63mB+t57+kyIdugKFM8KWmMk3GeKcnOE/BcX
e57KCDYTJnmsfu5ebDVOhqw0DxwJEq6FISiYC2vwC9W2W9FrYaq1d/oF3oBehTKz
An5nlOs+A++cUCRevEr7wSac82kxF4Gm7PkiMG+n2CfGL/hWniqOdUWhAxaSDNgw
0gWqZFf608LRAdGV5cAut4JlmXrkgsv3dmDicmWedy4MEj0f2hG6vNqglijUOJC0
lQ16SdObB3LDxFeukeJfQtRenLLJM2AD8RGOZOw88zk=
`protect END_PROTECTED
