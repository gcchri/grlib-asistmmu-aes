`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CKbRSFe1uUUpVHXkEzUUPIANgyi97/EviJP1OKsADs8W6u5/zLMQDjwGi9XOpEEh
1y4U8ko91mrfmrxCQX1K9I2PFnZHHRSPofTD3MX5TSKzfiheM/9n86ZFRsJTNNIT
1c8ZkWMlCKScSQVZ2lG7D+B6U7sqJShAHsgGKx/AX1rB1lRaguzpRs1LGqShEyxD
BjFO5KzPNBuji9Ttw3zq81Pdgqtc1YWF2BDtUNyjPPfi8F03BtNqxZPsI0VP3fdr
dnapXpiJeLjNRtzjtbThyRs8uVM3QkvzZ0L5rgHSTjitnQqwhVaLECmIzuumffSb
HnxZkfGm9x9yUp7X7pm2+d+EjWZdoq6ryPRgA003PKmy6rYbXuF2Ba3nW18UiTgw
IcNGcJgkEaH/UA3uJWAfKGOrY1LYD74E3j2cnrJ8nz0nnBBXurXSPlrh4apxycDO
iIk5XHwZ+VN9tkTXvZxH+vUl2/AUicFEGBGYd8XAkez1xneDisa8dcJHtEhHTrIu
OGEoR6IvwlKGdSuzQxgAEyZRZxez0A4k5Ct4vFFIagVeNzRQnLc2bk+oyoaJveGi
+0HC3vvHpCGmXjHGHOQh/53eF0fWjOW3Hf3X0NKVvC4Wu8CCMP4gTtH74HKtc449
jr5Bh4rVtsNC8MotJ17BvAtvhK0n0OZ3IKyXSGHF1bQ+j7g/kx/teKMvysLTqnFD
I1RjGf9Izi9Pblr+5sPi4AkAoRJgBgKLvIaFwtyPQo0Cr9UEGyng9jUkGRZbiB4E
PMRs8MhISDmSZ/8QJMAde/MafrHhaNuo5SKNjNS8pcdRVJbPFaD9LR+fE48CQxim
6OBsQhDRlKbAfxoxF/K33j8eY9929I5iNpeUx7u/zW6otC8+c0xuzhXkarcJHSme
WwzcZFN8GR8ldBJrCUmJ07ZwWV6sI8o1yYMcJHHqtPgtKUE+HuPrmi0p46YWxYU2
IYWSqjLx3761kYRv649wmDNtusgoHiwi8o2sjywdTs9XQ5l2uT0XXt3fUMtbAdj7
`protect END_PROTECTED
