`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eFWRjBsef2AeooUEX13lgos+ztmSYWRBomow4BYiqv4tpu3xokH4HhTT41mDEsHR
vRbCp07dj8UZfV5pPf2UexxgLIXo+7yA91dz3J9CwlDmPgdgyvFy4RQR1+HrdxHl
2LFuXBW4ttm0elc5r0VvnygwgZJ5dq8i/t9mtna4HjQrXXseciwK8HI19ETHzmDI
IzLYTi+299RS45BR5s2k/Yd6GjYFKfLkEADJe7mMAEsnVFQFPPXad9KSeod8GtZo
DbbOzFiGx/Ep4N5eTU79qebCDnnkt3e08cKKLaEeCuQZLb9ezorgx2RulpPnewT5
NGpVTHdbSsb6wRN7riRhxKakan0Z/qNJ40N+Y9WGDBw467e8wji8iJuYdTEB96kY
AzTmhsKHFlZ6I7GgUTAylVsx0EySd7mLsLIJhKNof81FHSFggKc6i2WQrsECZkaB
LuKSpB9Z83/tzZcWj5HaseJLwIACze9ZtnBePS6iwnd9hkRxaXbrZDlXKB93J8TT
`protect END_PROTECTED
