`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6NbEdaTly2UeYCsf1iV9FmJRe/Gz+laz+gjuSUZrzsZZh4HgBMKRuZAAq07tOCzR
vzXlnWrD4/Kkr4gV6QYR1pJQEAW3bcHkcoNzE03bSoYiE1O2RxB6gMepTJ8XEaeo
20Nk/OXeDz0dtjkUETJbOrtbbz++uytakysqJ9Pc3NPrXCZ6dWptcpjDZGTY+/38
CQ4RMmWgbPws4Ye7Lfzfg3tUzLuYUYiIYMSFXMJNePvKRXUzukmuyGDPVNVRR83l
YspbncKniDZLKr+XUQqOqPkBv1pWa5hD4c4xutV86ZmPhoukZzolhiJg66wXdRUA
xP+yGNAAtMZnPQcKHOOhA6IN/pYy4GW6U4au05NospaZ6UIXA5DSz/ERPk+ME8xp
HAUdWudOg6zQfpXSUP2GLx3nKNGibPZqQtn268Cm94+W1eM7L2Hb6mL0LQMZnG4z
I3LW78X975FAFW38D5pCFzhGVyI9S7ihk0GLG/2HcCnUE4z1mJfXB82eUKxGYq/Z
UPk2JHyvNxhZaVT/TGy1G4f+FardVNKwtpdhsu5ghGvfJBBMeN6k+7AlUnVyXeW5
GyMYI6/0OlnQL1YjcIM3ZfHvO9IgVCrCxz509hzGBSEPB47oCuY4ByeughgNFo22
pPj9rUZtp80fFkwodTC1o8p3RqBMt43IH/JHFNM9AYx6cSV3cFjMgkhTmDGbKIEZ
3TJdQU5yO6GP5YqabKwlqQ==
`protect END_PROTECTED
