`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JajsNrE3QA+6WXI9pEal2lEnOg3Oqr2Ym0sQ3Mlc0EVMcvRoGrXAc7TqyhlPz0Kg
ar5sTSuuYe0iqSs95r0adcmt6kudAj3Oxfl/GjIlfbD8OAVSXsXfggKexHfU/zpo
ZUlogc75NcBZVfKscEqms2C7OhA+BRwXDGTbSxnxCGOA8BZUH+szQZIlZChKdH6M
g8Zqzb0AxZ6jzayu4FXtxhySI39/HerlNDkqyH79mTok6psm/om1v2VpkCZsuGqi
Vc0et4cZPMt6zl+NdWecBgU1rbVU4pV/6Wn6avTolKH24KWpSXV3kRBNspLlFZSu
KeyYOC9Dox1BjtHZtygEUnFGhgvP9/KIn87aBdhiapqrVxcRG9tMmrbif9ag/Dux
`protect END_PROTECTED
