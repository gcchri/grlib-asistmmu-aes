`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JsQJjYclpDx5AEMV5+vVxERXonOT+coCgodOfCdqyaZecIxekd5P/w88kzohB4AZ
xo6pxtoxZDpqr6AhzHQE0kuirCCya7ulH4ATVx1gCVWa4WmDjzJ1YXpYBZPGkCpG
OUmj5TuN7xqSAoMhJwwQbJYuE6gN+8fWkdfM8ox2LGkx5ZVnY3paKa/yoyAxBGF6
JSl70o7b79iG89q76oTdNhhy7dt6rCltMIlaiAVuZ93FWPDi3bDkbIcPvWBJIgaR
2DwKpXjx1oiWVILVU8jRs4JnuZaw2dVfHWn00QuLTalDBMZGGyR2AEpjSvECw3o7
q2ivxxrssqMBIN+mVVIZq/vs8I1NSC0I9F077mF/GkoYvj6HGN7JMHuogVUYJtOR
mJXz7DTeuaJlaaNla+7UssjBGW8J7CKwc37Es0fu6Wfu2kW3WkIH2fqGIFPPmn2N
`protect END_PROTECTED
