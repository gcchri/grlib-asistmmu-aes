`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0BAAUn7O2GFx4dT0R1ZHz6Ts4F8sMe9Cf+yRBJEtW7CwUIioToJZzy5dsFBorfCZ
Lh3D5hWz2muN8tmOBOsG8P6eiSEzJxiYSA3ThJl+eg1A7E4BCxfyV9YI56jbUTzS
yDHQBqcJnY136FmjIiJ5FlyH/I52AqZC3bI2m70KZO3rHBWblvSsBA5HlQLrOow7
KKPXtioQX+yIPo/5KbrAMYuKGeNfUPkhBbV9oivb+AeDW4NN21rAL/3OnNkQ5VJW
CDGJkKCSJur9w+Is3pHIecm3Lt21jx53uYwjYmYf63Jkwn5JdVLNQS06H8HKN47S
o5H3oM7MW+J9u/HVaAd42zdsFkRTjQ7Ha9Usv/0YU7wJyzmFumTEyCAHprSzOfqF
oLpehcfyCWbZQWbxwIrlFIh3T3qWY4bMYzhZ50KIdfU5wwxbKO5NMgrtltVVhOec
poawE0YDLDYZx3sT+2KsHJEDQBZdqoU0caGYGOOpgfqXHueME4+vvjimElI8dC0H
GphS39Bk26Ts4spbu5TAJX5apofOt8ms7mqhe1Zp8MNbvqgr4VzTuI06N2+FvopN
wXUVYTq0w358a2QCVo7MUW7qDKaYG5h/HOu8G1peB6mvEIFbjbn++uzN1LpTWtYY
`protect END_PROTECTED
