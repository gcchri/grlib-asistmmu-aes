`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Suv5Z1sWVih15Klh/RjR1So++s+Pl//i9bKUxU70hpHK6wAMhbtejH7zeDQZthj/
b7gegqTdyRXyKhXUtdud2nozDQtZZ9M3TaPlPg2iPqW96PkG3qZehp2BVbA3enGj
FR7YLEKEUtH6PsxO7jHl113Pfg+q/Q0uzHzRAR1vrTVXjni0qbbgAQ3zHRBi+ziz
pFl1KxVbRvY4upfxfDHl1Wc2Nd9GDWmzHiNIpAROnMA7maY+J4R4Vh8EIsiLpaa0
tZeLzKqoeHBcSYAfxHiPCM9fCXWRE1TVSh3aCitj9PIouNHIWeQFC6HC8BPke4b5
FyeBsEZaNkWf7nkBEK1CSfH0+bSMKAERuQ4PR1g1zIdg9KHkc5vMrMrWSOAfw3NZ
NePafUjruucHcWHwcQ3sRGXbpwRfhwRBom1qvRC8Z4/LYxhkYqxdi5gaYMEuvuPD
QJ6u271DawopoE8ZE5cT7qkfSQgj34/1Ca+6XjOW/NHLj/a1OfeIfKjiGzmJhcZN
gxoq8InyeENFQZVJq9Udxqq9h4I7wRRu1uRahWN2Fh3vuW58iKdt/r+sWlbC7Xiv
Ng/gayBv7LF23i06w+IdHcWeh6q9HzntwzXabYeQn6FafUebEzeraHRU1VKilbG7
n04Ljwkz3O8fvofvgdDjdspPOrtNZAvy0KudiCvAs0SssNrob79r4f8DvwrNmB6K
5NtwQOwWPt0CmRFw4Vu2Yu2GbrBbZBDqdeLBBEUeeWliN5FbbIQBxN98VZmgkjGf
3DBr1DSCfkkMa7YyRUP2O4K95vsSlgiteLg/5YHi7o+sHRyXhUk8BTz5eqw4mWtJ
bhICgnhDaNi7Lcel90f6qpTN9hE8NeNp9i1jCK8cU7WHparcwYpiIZDTTS6d2JY7
MJqg8zDSrHLZ9BHQ1XrM5Q+q/bHyRNpTQHfHcZyl67z9+aXHhwndjx3lF50Uon/Z
joKaE7D1gZxPZ/qtixE45xZ2P09fn8qbYiBGm5Y8ehikV+I2OBYbt+57svNy0/OE
`protect END_PROTECTED
