`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GsZpDaSqE6nrkX1P2xMLG8BlfAngJSdkIdH7g25h5BpaLQnu2hfTYmcr0kIeCSsX
wISaxAjTdzZks16XbDMBMnkUBN7aXwDzuvsKmcSf3q8f4cr+lnr7RUKZ2RQWI8gJ
WDBCLwgLJjtd84Z4CMeI0cmhv2bLjeAobrouTtU6gpzP3zyV7U+oGke/ya7r2WTi
khCTD1vVGklz1OMKkNBMlNZmhbCmLitWJMldVcWwWOTZMS8Ru7PTa2E0jWxKWz/R
1I+fMk6IzTi0yBjFubeeL3GtQDOCdgJct4iMagoINf7e9rGhClNayy5Yqvt+VDLg
rtHmfe/kDH8xBp8+eAeWVfxVfg1Co2kPzJQpYZviK6oQTdwZjDwQsyr98m7gUjdS
hiwRUNhNV3tai4YiftLKijXuRuRMVD8SAioCvjXHxZ0TEmQYBbS9upgc5piZyzCr
lRu4G6apJrSeEtv8EH6+EOWA7Sy3Fwv+Tf5yRy3c6fy7Omb+bY4kwdeu3hh73o+4
gP3+PVgx/UgKi3VHc2zwJ5gUGY7dMszIo78brWXq+AxIld0wRP9EOXmf6L1CCD1r
tyv5lYmcLlMgcYeTDrvhGKYA/xxiZTck24yDoa04z0oFj8CIX8vEhN9VXO7sNt+3
4MDp9L1F4u3YtaqjxTXsqc47KUYdcz99kxCmDDTYYdyJWdEjCD2fy42pyNQ17ahX
nk8qlDHdQcyptVgPWSolaje8RXgLetlsJlODWup5yZo=
`protect END_PROTECTED
