`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nvO2sO8z2UV74kXgFgPg8nO7DutG0hO5jTha1Fu5VdD+nTbmAwmi37tn1xjIc+7j
+koJOZeHbcoaJIv62cG4tLWUKtSVv62KdG63k+ACXZGlU4UoNG0UqjVtTUpMsVnP
wNjnPIdHLFdbFpr51VhpHiWRX8pPRJEvwCbz79Nyf3PWU3Nx1n1kbXAfAKB8QlK/
5fseyWNeXEE38Gwh1DLKNH10nHgy8czyaK4TAZGG7BcIAkU5Vms8fmWg6Uc7Zzug
jJkWdxllw07c59MoTxZUTR8yasLzSajMmknWFTl0qxTZ12tdUmES+ujoELowj9kL
WBh8IrXrR2cdPRcKc9BPVz+hso8cJC3OFiDbGVUnUeWJKAFwCr/BLIo4Zi+Uupfn
6EpAkV3fJfvqsljsf+4jFyzkd2goCnuGZeMgugx1qUJ4B6qO8JBqJVodGYhgWLqE
v62GlTNE1Y7l9fYUJqqYbtWNGhmTRk6PlD7Yvu9PbjapVHtSCYRjLlZttJBoKqu5
7ibJ6MBlLl36739QTWWfi3/NsGWgdkFY0GYsK23P/z6Up+v1FG2OncWcKHu0hAnn
DTavA/rdyb5SF+U5lxpnLTzDW+KkAx5uanj4tRopsNcVL0nuAux3AX6EGJs/zHgj
qGfgriHwgY/eoVoDDnMV7LJ/Pnren2iGevJ971fwPSymg793l4t6Va/FvVta8tko
CoTpJyUvrISbL8jWgFTvBF2IsQyNUwg5bRfTC6H+bjOKXzN38hcSC7zDn1U0rvV9
zntFztMa6by9O1GusUG8+wY09gSFB0cLfVV/jsHsUgcmwHkj87GSo9J8C2H3CNqR
C3d0nEc/pTSqWK3Z7X6pnsPOnf8Nnp0Yl7tWkr7Uzt/f3tnHH1szdwelEa0gic0V
N9xuPMaiSEbR8RzDtOXp+R9HhE1qg6C8lCF3XZhMMIM5nxxQdITDWMW9ZYBt9630
aexCZ2f1tuQ3YjLbLd4PUtds0I7PZmpJcWiM9LXkqrravThjLjl7BO1hyCWeAmV3
IFiD6SL9AKX/2T4M7zWE2FmbXQWu9TgofDGgrcW5G3N6tfMMB+lsVNhYj9yZCH1M
i58T6EaugEuLs4OoIa7usbn46fgxHX2G3T9wR5vEG1GSQGrwhVnKo1vnvwJz+wQz
XdWqzYjZlRLL6HAukEyxUevJNncLD891NZLZvHb28s9F8ZWsjYYF30X5qcVPQWQW
L3xRENHpDR6HIyWy+oCP5XVmrg6hqW0HhOQdI3+fuAJxGvXyySGUia186XkfHEg2
QESsBJY0ley3amo03c6aeU76bMkPtkWBfhfISmHIAnpl7gZ451NcVKyi3CkFW8Ri
bkIZKFkEJc6YBVH6jw96Z62c97mDr8DI5aYIn7WdPYP4t6OG2GLJqfKBIRR0rwTU
2Z23rQ/BAtOTukNFCcaweBbUoJpx0q5bDt1QwjdvSA1LjyGYWKrTrQp74t8IM4jZ
m4al/+O5d9h17k8diaHtRw==
`protect END_PROTECTED
