`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hA2KAuQTTTAWGrojnv4DXbkcjvm0bu44OEC2y2kJuMy6R0d4J6r6oRYqxqf3ghp9
W/I9k4A0coyTqmAQGJRfv2mfcs9FLOU0Na6TOcEcLZVr4ciLO8yZcgSrH6rhvhoJ
WXldiSJL39wxJTwl+z29FKlL4guSSJVpSLVMyEd22pXxputNnhrg4YxY5bgnrQvI
TGBPssxaFoHLRy1r7h8MHtDVxypHBVBoUOvYRxeMSccfXk3Jnc20N8/9Rm6bGc0N
1r9uIgFq06dGUF2Re78nAlBzLxwt+UGNpFnV+xxzgHHDTbzjG2RwDtmMc7Pv7yCu
uhH6lQULZwZLVJ2tvT1rllEEac8m8Cn5Y8QttiFSympAd5OR5IAZrP7VHP5kgAxZ
a96boG40PdnjWILEZ4m/XIe4NPNQs8nDG4eepT8K0n/LFNrmHk8ge/xAqLhlniBr
oKk+YoPMeyMVkQFPhFV1W5yfItlv4JUKKlOMRSLyZfklsmNmwVU0JsaXnYSIwy+P
OC4eDqUKQo1dAuAXAcANLdZD8er3CGU81GR2gCvuQgJ1SaskKN/o4Fe/TSvyHASl
27iWnJxi+CeVooXXkg6yvZDzJPzNuTO/lHF/VadqUiuPBhlSNT7VMjk/3umiB0cV
gJcDqdqYgxVfuLOe5pXU/nJz1+8rsp2bLdESXeJ0K32/q8qtv6/kIRTZQARUIOZF
/0Px5R5Y/mThBcdJwy4ZbENc0ye5XEMHdJMnIaHAIodxv5J7auPKAB3o9ka9FCSs
956SMJJ7UzALzON226xYMw==
`protect END_PROTECTED
