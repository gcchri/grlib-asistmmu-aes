`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bxLLbyZque/owCiDnpJ6IQAfFoooRnrRwu/5Sg5nPjPoMD4G+j7lC8PLnzVc8883
zJHvasZF5LQliJghkB1mhlxl69rkxczpu+oLBX3o2e0m7tak6TEgaNe3ASmcAHDg
n/8lDL/S2Q8e9WRSVINhZuVJ4go198keYmkuEUmnUCA86ILgzaTLo3Ovdcf4e4Yy
25itKeBWTzPWFdgja9IzE4aLZqkfiGBeZyhdPZeYiNS4D+r4q8/wD4Z8JqICmYwP
MljrKq8YogM/UCNXUs2ylhLRkYrbPu5+zL4NiO/GAxARDzg8vnuuAc+4gOyHoLix
lFVgYHM/TLLEYp/lD8Dsv3ysT0qsgo0otdNqZQFouY/tES6RjC8+9N19SCSdm3J9
H2PEZkUePNjc1vPOF49Rrlbqf/3g2XJ0ohUT+l118enkc8ZKSQmagD+p+WbkilOa
b8d/BJzVtAdzELtqe2FTC3JuyH9O3dWjAPGs3xmsULrAd5t2jpcIfjkE9IK3qV3M
626IWf7CAVGFtkcADfMlyeu67oDt/IXNVd6g3hLJHNwXTtFMn3MCfXq2Z7q+jOwa
eNOSDtGsISixk17Tzi8BKaBgS3wW/Yyfue5D5pykVfhQl5/oSRkHximN16ZMv5qT
6nGG9Woy07GzJNoKAgogA2uYNnn/t9ojIEeVwbpylATvSAXcC4U9Y738ngupo87k
Nb7xSkZJGeWS/A49KLYH4A==
`protect END_PROTECTED
