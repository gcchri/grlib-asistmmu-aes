`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VsgG13fF2az7572V+L/YWR7nD5o93w0NaG2250gX+dOZZcslgNpmnizB1yLfmSuU
Zzrkt4ZdR6vEWftw1UDq4TTL24zKDGdR4LmTOwwb1TyQ2lqckL2wYMzxBvTbOJkR
Sui0I4jmFbMQPp0LY7FEtVmoCYFJLynk6Wx1DEBqNKpdEtJ5enrcY9yXsRH04NVU
05VeeZUHtMmKM8RiJwgZaJMAW0m0qe97KDTuwncBhP6AFXP450z5iketRKmV2UyC
yeZEJXcLKFqYKjpfW+eeUWinpwZTTc8+6sojVQlauuRPZp7ABMH+2Qtzo3Rb07Qh
I8i1LBl5OM00yEOtvufBa6EnN5/2djnkSqH0SBOyiXmI56gC6u1Y3IVW4NPd3ukv
6/tsXq5ZCc/hqqPRvojtvGocr7INC8CNnRWPRxCxWXQhqMmhcm2XxRD/enjLOccx
3MWhzYyRB7TQtMOv7uqGB2zd6RHBtHQw7tpRq3vjDQA=
`protect END_PROTECTED
