`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KuXn8vamV5pl2aBl43wB2utPWU0QvrLC0KSXzzrxAehVAiIeFKTg9o3G7vIWLLgk
xYhMeBej3eEiYWirhysAh7VCQpfabkABovtpfOE5oZxc6BDpRbqtNNWsjpAExXhu
/qwzb0AFwBS131JrFmy1fFk0/jDnoe+E/R49EHWJBawvcCti8WMsYBE+eERbHY6f
2ibQsU6F4WXq8PMbgdULdadX8BBrXMienP7E5/K7DlqrigR3/zc2pMG8SsOe2Y8t
xrml9Gw/ycmS6beSdGXrfBTcA5xGVjT/BhkqBYsQGMqk4D1pqMQY/ZIAQ0zfTAhd
gix7XbRJSxfMnx3fRo44YGLUm83creD9RtiCs8iUbOHzobRn/T4V++yaZIQbTZup
0RwtUjqy5u2vBW+JGddvrl/W4c01jfd/kiTYSa8GafdZN5Dshj6asspIAxGF3ase
cbKS1r4NR8FMqjMNGNZRDthihFDQPiLrcvVfBjJbrFj1WGacFY9zRJETLMiKiQXh
jw71HylwCnokETCesTiYJyayo/Epmol+nczuGOEGvG7EOiSupXB1rfkWR0CGWreL
BBpCOc7alS75sYF7aR1n4EYHielRrpBRuM15YmWA3CmZxbeOD2eu7RCpVZ59NnZQ
YKOxPL8UhTI0Cke1SOp04xZOxs2RQA2w2GObRB/sELaJlcXS04xe/saGf51E/Nak
8KEHcBUR8LaoHtaLXS0NjWr9kZFYJ7zz4wsJnSutAYl76fco4qZURj3Nuk8wG2Tt
do9277VvfeAvE4d8TtYHiAvdVC9n47r4HD2lJif/M4wy/HswZFlCYCfzZMqkHVdm
srrYO5AI1hpcsC6DmUNPGkXcYw1fCVHHNhOI9izY3Ybgjyodf3cLMbkaFdq5xl3G
BdRF++O4hbQ/w30M3eYoJPwA9plYhYeSMR1m2ep9nwu3B2MpJvKdZwwqv3ZPhgpE
wn8yedtuJqwTZzN2HJOfv880235deTKmuwNWQezngvZz1DVvoap/1fkZ/JEKDVSI
LqIjGANd8wsMNU6zwxLLNAt3+EeK/vBvyvZ1UAaNfxQQd143gHMaSPSXcMJGiNss
ZsmKXCeRoEbK98PE+vGMY5L8U5wMtUcqswO0aqb94Kj3uY+0qG34wzqLeAF3dzJ3
dRfv675cGlqpMQEIH/XEAfTmxKAR5SHpZuKJuE/0e9JECdXL7WZ1hIpe8sTieYKW
bYbJPhmqGF2bsefzg+igz22iD+3c/S71ClRHeDFEynck+XZqM+v/VPNAIdcRe2qN
GP8wkOanq6R6+AA++nVYIi4AZ808QfxLoeAbzUj81MTlM6WVpyMO8we6ZgxUSBup
1HQ6BbIyulBlgXlRjmw8bhHFMMN3JqhpLnPqsran2hVbXrHD38p/bxa29H7xuvQ0
GXiWmzrvfSkCkTpI3YuBFZif5bHOCA303GCAnOVZUF75AswjTcc2ZKMeF3684o7X
5TppS+QlRal5kyoNL1a42dDQIEEHTVFvs4ecI7LtW+NJaVcPM3agJ5hCOHp9Zg+G
4EyvLT4AKrvIMRbgRCzGd8CKPEOH21lVuAzGKdVTFZSVdlhiEhx3sX0yfynjltb1
qjal8fHa3zO841X6q5qGaAJFxEBNLGQCqlHfscSO0yEW8KhwCNBtHmsouWOJyqpB
8ugq34BM/gHaTeuTEKSrsGupuI8XXcZMxaOPBcsJ/jt0c0BScIwEwiSU7Q409O7x
c0NIUNBqqDn2j1bvN403S7zMCN36Hta9004YUyyOqKYqqFK74h7SxhiOwkDQHOUY
Rmo24o2qpFQnF16DcT5XzVktf6Lv8t9s0kXBZG0N8hSwIAfhb2yxnT3xegjkWrr4
4F2ca3eJ3MlL5qdrcoOXeFxBHamu/UhrnMXybPURdQKv1o0MlfYqy/sF2iHy0frt
i9Z+bGXHMCI0basl+BTRRxP5ZhDLw8aJ0swuzSDlD5FMcgpQk8Eqtle0tggZ5BqF
iPM9Yjr+KUffgYCuJfI7fdMWF6Qm6TyMSbYBzGtjaWHomIeB7XXklPG57jOJgh1z
keyu5iFrIX9Ol1Yu/qS7n9t9Bt2spCp2wYh2Ye2GpNKxpGFcnWdCHsn9YnS59xc+
KYXS6u3oC/0MN148y+yz9/biEYoDBIEIL6Dh01nhejhKYtMakIr3QfEqKn3CYohh
q7CYxMGM0H4ZQzOkw5I7bXEuDap2SY45b5keCWsGXxNp4lIKgjBVGhrSN9E+uih5
sLEFmsW9bQRFofkKsjWleBRPaQYPu0F2ehZyW8A+myn8yKHb0L5uVWG4MhddyjEQ
aqQHefmTfk2r/Gm10oYCx6xdESPLExD0bHhq7UEGf3/n6roJkIGvG2Cz22bTd/mk
6zkLqB7aT+rNXc2uIdehlEPtv1VOoOS9CFGvPtlb9Q5BP/tcyBQiGR0AyMuzm5KH
oXjtlOH7rVs3wejqaPITcPbadpws0EPSRl/BT0azkFAPZ8jJ3yrkwP05/azjaXMh
7mmo+xCGlBkZZ86gYZDHpivDNkDDGPn9Q9Qb9NVTlukH3zjy1Yrznb89aq32R//c
ITAVtYL1g/i2CEuH8LRBCeeaAm6Jn1voD9Cw2XssmpLBHzTJ8yZlV3IFgJ0jnyGs
MQbk/4u6bfpvaQW49DhboeUOfxl/0wK6tmh76+EJHS8JklgQ4F8NF4QcOTK+KTV0
Gmpq22CogOSEo7g8dGynS2T9h/Pm6wKGoeL0j/GXnM1A1tZ2MY8Woix1xn3lj8e0
tGkY062Xxlp5JBs2k4m1ssnMNlE5ArOsRr6U8I6tHJjXMyNsZPtQGtSM7plQClFq
6/ltZM7fZS3M5lAXbFYG47TVkBYdmYgKJCu4Tl6txUPj3HHjVSF2RXfGvP6KwxOn
AIYo8gSYj+TLGKJMYVc4IkOsKC0bbqr2gxwywW40aaw5dtjtn7UHFihrkb0MhtCo
v7UbPK0cz/8XaMLCEgcv2RGfqcDoZm1IZrtjedtvF0+GdZevtSO5EzYbgMfOP3RX
ZGYcrhUVv1kRuof24qW4x3UcxOuHE0ZehwmW5BI+7L/eYPitfA4QUm9xG4ik2kAO
Kf00Ucs6zP9C7ptguvBHE8vUSjfJHEQndxgnVVrOqjYtUs3Vrf9jaI8uFQaF19BM
SKN4RHo5zs3cLnTKlh1OWtA5a2U9kQboWR9ig74fN/Iilw2MidZiGRohWUrf0H7F
EFJJ5iaGKDabNRoQTdDkdJX3aeFwdq2VMVgeEr48tFERkCFqPgUU1xh1+2DslQrJ
9sHS24zPApDKwUne+3hiAgvxcwAccibVRP7iVfDU3ikpiIpReooS5XkIGdAYofCg
LTWsviNNlLaBacsK7D/f5uKyMe/H8h5ChOrTH4Hd8A48hSURF4bZ3t3rpHcemTD7
NySXAnDEdxxctPoOW86rk1R7ZYdu9dbYzH4VBxnctZ9MRhpLX0Uw0ouPIi9f35hz
ERowky0rQAAjFM+gnqr0cQLTB1AAMBeqfHiwhe+426njtpBULVAzjhxkuZQQNglh
Bvg3FWscz/Gv/uUs67pj5pGp7cwSuOHcQ+MyjVqv2Kdb8cW+Xl5/WHuUvWdr7MdX
MUNmmDPEilpxC8rEUfUekAewVKiE0Co+LR9E2AHqZ0oAOo7wv3Gi1+t2ABrunuDL
N1Nx4cHONNGzA4EiJXC1ucIHpqBgNEOp4Z95mt6STFakBs4tjxFLqTyCplqf6wor
abl2sJEB+AauMXujT+spPTETrksetQYatpGYBQJDP6uTczVrbR/K4+f/EpjyECRF
iK0W0uuwEVocAts6Y1x/ok8aRCQgPgbha2KqewMa5yHPX+27ZwAayC1yHr/7d2NL
tK74Qp9eQN5ko5YUTeydaDxWyY0TqqF3J7awwLpULNoslWvme//ji3jNZFWMhlgX
XmzxB/cFRxkEMzOxI1Y6Sn0ouvupGgA1/nWnwekEuhGFW+DZnhesQ0hprsrj6hIL
xGUvjqA6d0ppFLgdZEkZgMx4Sqq6G2gwN3+Lt/MYXYv6UENmouH+tTG6O35tftTJ
TihIQQu470H4H6j9R+/1+8CuQkXRR/g8IRP3g65KlL7VW+afdSjwfcVdZg92CGB2
qdvWeJVvOkhexu4tEu9HqHK6JAg0FzUqsyGdnawFObdlSon8DIemKByhHd7/XpU3
Iu1luWCNqfXeG2wXfEWte4Iu9Hsv7G9Gu86nSAYULt9SmZcubJMKvg+2syWdiNwv
GwMYNc1oIDCm8E3XN2PmlJOo5ewD0DG0hMVfNgCAwz8U/H9S5g4Z2MLBA2cAXDdz
CAmy/hFGPwzHbanvCgS6CxGxy1g0zcc1JFCuKqhQOzJN240q3V/+Vo9LiThf0Pic
OJqjBh9HVH5SBCm7HmVQNpAYkszWWhgWxBfUUJLxZyE3xbrNfc5bVWFDjtb2i7QC
zcTuybIUzHTL1bYfFspibC9aJHmNwR980Jf75B+CmWyak9jhrLTQkbVSXYXzVOu1
ZB3gM+f62n1zt2egatarifaC4B0QI/ez+j8EKl3T1L88b4fAk88vVceoXx7RZfmZ
6m/gBG7D+dDxsmY/32Gxa4aJymSPlvo9DxEkiz08m2xV3ytSgHcAJVkZcZcYNTWZ
pPK0YLjSTps776iBJCWmW0k+fLQv/NM462aE6GI4iluWrPnH9wfjaE/eE7z4aMp/
voEMVk73EoJuGE9ZrEjRqLaEBLQnyWCkYsR/CLwIzv6fTLJDcTCVaBBQOqIIjg/e
ZQOhOYnTIEVYKqzza0RYROfrQfMxaTy7gYGOaaEdqcohl1wqNpBUU/hXbidkR4v4
83JR2T63SgQfRvoQiTfWsS6Y7ooZpFxJPeQiTwxcIQI13tnl4XrDVE1b29RXOoOf
5zvcGZ+hwAke7zfd3X6hXvcWR7MNOKxGqF545pumYuY+s0XRRiTeTBgHqelLMH4a
c84oI/MkeQCL0NvcKiOcNQtT+ZYsQ9abKmOUuoGFYXZMS9+8oohRnLCNyKxHU+PQ
hlpa7XQONtIb2/rgDGonHOoDWXZJEGNslx6gEkop9471hpLoHONkumJTwHB+OrKF
JHJizO1z+juWgK5l/tk72abcwTW7KVo6EFuoupotWfXMzwbjHpCbPnRviZnexGs2
C5wOyIWbyf7RO3tsM5QtrjYJusgVQbcnhQWF+UdFFTy0+whMkHOL/z7HvYXIGhi9
u2ynmgh6p0LDl7lXpYuPX1iEBx01UtL6HOFTPPFsCOXXJ5LZTOC8NjTCeNsS1vhS
hA0ciaeBEaRCz62vgYyagTD74yx/D7Q4lEn4rPWIRCjwDl+WhG2wdbv40ObSAjQy
P/oIscB9HLp32lH8Lg8u2yahCOyLbU8n2B8Zt4r7s5rHq/sX7IfNkBwV06FMBHyk
efFDPm7xyjM6oGZl7xTFMg184oVIBnt+Ym41/Mh7AzsDzwRbxSfHO34bbZ568HaH
gAMRJdPde+qiFNET23luH81Wf2Yc+1Jt1Vm0bEY0fqMnK44IozvntcaT/jZ7n3X3
sNM3i0vKndesrLx5G1Xp5JsdVjm7KATgH1JpsX+0roYd5HdCYBkN6ucfF7Nw3dco
rLMIjFmMyxAh/InOBul9Hcw36nznVYkc6UMmUPZMcZxixh1mf75+fZyQbQZDKaSD
ZIy3aiN8kCbrSo1CgsT0L8ZMMotVUNxl2dd1O8RJJFMDRsa2unMJEzXLwqj4qSJO
xhNn3Nzn2705mAJHFnnOzs3b9Fy0iW/Mzm7nya87iozA210/vnZCNjnyDdGB0HVC
hckflwNuuQGwMmuCJ5HGtjorPm+9eIHwC3AcHPmi0j/yu4daQuUxwN1XUq0j7VRE
M6VQ76qauu5Ir+1olH9cJlKdFFOK+ZdCSpD6UGeMyY4/tXBkJb1QoofTybnJ43aO
7YOddWMjFrbMcePSNIEEWxt55p+GI42Xq7YQiHC7CL2SeT/8i3dkpaGBS63wUMsr
uz7BUD2IyleCLIioUDcwtB3id/nG10Ftqxfhagt6XR2PBcKBQWO+SjxUHqplBRWo
h29fgULVTz7piBmLFMgUkTGcQTPfxvBTkSs3aaPGWFbe/bDGZmDsomXdzlnrssj3
RPkoJ4X8vQRisaJibKMo4VopDtg3g69SMggp76m8onVvyJFV53dxWdC/AgJ+e8vN
RfYshcAzrr9Lmn+yQMJojyslE2+leXT994FCFyVZgsNXheMoozGG98vDra0wjUwY
9e1a/VCrHpyfY6/PnXuQ36Gn8P8r+v4o3wxRlIxm25jCmLIc67WZIgcTO+eib3cX
c6vI0AeqtnskeDwsrQ/5p6ApwTqL1/iW3vj/I/kqLRWWJh66XhGMAZ8wFIsHLhap
7i2fFQdIjoqBADsFfnGOsLExL+Mj+GBHJx4+HsaYB4UysFiySKgItk+hvaEDrigW
97eJab5wYAOMECgu3cjjRHibCexgYOirZEd8BYfX0sMfIUtqoZbQkgsJGNbeq2TZ
66oTV/nZA9Gl+q4BunONIjTgvqNaw49s1yoRPPx8QszCmWWSQ5JcFZheLraIKiDz
SYgwTQNPKVatGFkSMALglxUXxrJjOdj5WwvVbe/op9gOaTc8uMc9HYV1CfYcHDvP
53VALbAll7ekUHI2YCnMTte0rFCjcid11VSsqkVsteU8ecjK3Sg8biy/Ebdivqyk
O01WmYKgCqS1giIIq4v5DlqIeKeQ5PAGySxwnRsl6pt3AVjZyEUggi2091KutJc8
gAi3LOCwfLEVOwfG17J6RxYZbPPheTs/hzj2YtF8T1hXphHvTweVJ+LK7Qg+ND3d
HfmmrWg3ji7Lqggjjcul22BxYMr8hNQAMKPyuGNZZM4Yb2QvVUlHKx3O31/hpFmb
XqEEvTgVzY6fiInPAf7FSmso6TbVwFH6o5PjipS3XFdjuqN3NrqdPFIhCuXz0V9E
ggjTpo6HsjARN+5HWxel1bexd9xLjfvU9Sbf/eFtSAo7xoduOm91FcZ19BNgLTeA
nBRP1FgS6mY9cveSZFGRWx9hEb9B0v9cIGSch8kPTZAkIQEAXfMjgh+mdxCmYJUp
r0KWTv2C1M2U+2caBMtAyRUj0UFMrkN/t5ODmTNn2fPquxKnHLTofRAL3QkYGpOS
PA2LFZgAbz6eiLiK8L/iAb19yGBdxWWHNUSNzeYAe3vKlQayb1lXlvpXC5hRt+3a
XyXOJ6lzLV4t+4QSbSb3di5mHk7ljK8H82TgRejjMqUvUEfzoAy/HC6LiPm5MbA/
/YsYx1Q/j89OVhJOIkmD9nlP2PRgRkfi9pATUnn4wvXUFbaXrZAyxF7KrEokX1hq
rTktkID6w4c96JGl5GjWvh51mdlruHyKVFENgyh/w4StW5UkLAPhWhoML5DRW/Sw
wuZFZYGzFXd5yUM+xhNB7WASlKPQF6NkU0OF+O3PkJG7Exa0k3taZMTC6CDuJQCD
UkDTQrjS31v6s0uazaVkfJFuTWV0BBTsW9BnqlTP9ky0sZS5vFJpuBRlwnWXupph
hynl4xMUThaUq3L2sNibI9YlnuxJ/kIBntFmR9Jcho/JWJ/X65CG6FtVy6WgVNf3
0B91suaPNa1UYh5Ii/d0AfJNfuSPk1liITHrMprCiVitv4CKWoqN6kurHR9Loq32
E1m4IJqH0W/jgBejfU5ny9Dc9e40XoUwqbfams20/DXNmh4ikHltb331Xh11hXgz
U1AQ4qZqt2PuxQTu85kmbI6YMZn9Z+TPdDTj6MTQBAwpWmYbxlO2qzHk8jCBroO2
+MSkkPLbGzYKdBddRXeODeLRIeEa+1Gs5QnFR85GZYYFLuEKE8DZy7dFu7TvQlZG
6Gob3PumCvuuHZzA1tA/bRoGMlnBP34gCSpjYT6x7dhkQtsNDb94vnRXL06/Zeoh
bTTy7KGeZdXzc6+LyHIDV3CT0pfs6tV+WqTi0XBxikcrOqVQyV7sNFDvXkFc1+ug
2x9h//t5v+G9o2AG//4f4+DskbL316cY1PCPlUfQz2q3ymfhaN9ZBszpfdKWAUgN
A5ZHOei+CHmo4KQmOrUuCyUtfcCjSFcY7pbQPdfDhgFmFKblzwySy+eBmhzErx1z
gnEkLRhP7BOtyQ/YT6/HFD652pmo2n63oFjqUEnD8uzht0Rlm0URTDQ0c/orNJCJ
rbMhAOlAxieIiynO5n07MTQjysjcjn2Xd4K1sEXU9wPdx4NolE7y58+PhCijI/I7
UGpaRa6GzgExwFe6tQPHq0EJNq60ATvx5JVl3RDLEhbsGIJCiY+76gXIjRkCyH76
ljyzDP26Txo2MVwu/dJyIc+sPo9pItyQmJ5+o3TIEEXXUHd1qYcsMMROUVzovEDA
6wIQNncp3dim+qcpg3pCmqKQb/+KEi6KlNAvASbX9zvDUNstWgu2lS0/jH/NvCGE
IMW922ejVod7981VB12MrD7uxd/JWN8fN6epd73uRKHFDld2kjamU8OPUo1K/7Jz
YoENk3eZ4i6Dl9rAwkI5K9xAKn/LTKPrQrdL879zCCo53cz2Bu4/ksN3wom2b+F1
asy0uol/TPboCOf9JfxV8nl+wntOv3knjZp4FyoJNa4GBZ3i+5VO1/DcMjzzuq8J
qU1Ng+8w+/K4QYDxF+hD0Qbv/pF74R7J8lyZ2d1I68mTju6PNNU2/wZ1By3EJ3JW
uKqTEegn09mc9cOy25aQyJ5U0nvz0XtltWxj3DTaE1OEEALXGNM/RkcCJZgioR8B
xu3alF0ZvxScfvBJ+wOMq+WZYh/1qTMz4As5bekEzDaFwyOAmZCQsfNKPZqYYf7u
nzzCeI7BmnwaXrcrS7+ZcbjxIZSNCOYol7kid7dvWIuhsmRu/quYae7Xr+4nMWno
MFXHeKO16n5SYXyNpmehkxv8VwdiJ9rdIQg6perpt2eDg0wAqoCHTomqPGROaq55
j5ZklF8JG9W51o3/rhBwxnVUVBGufxuJuBZmrxEYqcPkNgan28c8aUuH1QfdVgI/
7TXcTxh29dB2uFOwk+r8GqcocEbRlUkn8zpxmp8MU+UuJrK1iXF/Sg99cm48MThS
5lRE7vH2JAXuyDJ1JGgMMjaxxElLLGSZZTMbYs+yhwB43yWGJEvt1V1FNXEgcLf2
6sCnjCRMUFYuFyiCLZH+gTY6iWWF+O6wE8IElLhn+Xf3hHG/hFfPv/ZVFCEYqqLc
pSyfyxy3VMrZfl/hTsVdBvMUC4Qqf6lSDrGdhRESLQALzS3ntrq/kHPFu9l6VV5m
p7DOEqGRdyzsHwigh3L87cCRxTWPvH0JvTF+AbHKZlEFzGLsGZNL/GnpW3GbfbIy
GVXdMykrPMICfsjKEFS0TXU78j3IRYnhbbADluOUQjWnFCPN5aHDS/3lvqU3pjva
PVUjRVvoSNUTZv65YyoujlqLPE1w1jhKmDE2x3WHcWlDOJWVXp1YG8CuEcIL31dV
ULEJT7ZBoFrQeknl/Lb492BR0LXPo40zbqbjmg8LJ7c6bdxi8YO4CjQmIT+Odjee
YSUHeqMbwsJYnjG+tBMQRwk8y6okm/OjZmDGf195ijUhIAlQwIUzXvWz/P5HMCnH
Z12xnvSUxoYCfoVJUE3mJ05AbB9ZWIMNwDjlMHfHqdGthuzEMeegbzjMvOXU3bKx
fBNM0q68g2jENfHhcFKeLqe1a6/ht8v0vipA02DSWMHwW0BLa29BgiYszhvdKSJo
hMCDuz/IWy8yWfTDOL1UAqug5HKKBQ0VryyPZIDh1CTMtWJryrVsFKVjILVTFQLO
qBhkGS/KZtrT5Gi3GOeT4ap5KtibbBqNpIdAf/GHqxrXLeByHWCTvSnWefwHvEQd
ZtVz6IKhq4paF7h80Hq7E3TDebImW3VyX85GUzkKWckqMXRK+14tUyNHvABDVubb
OU18GnCx2D12XV9P9AmQEAVWiCuTH6QERx4VW65VrBCAJSEbAmKECHwp5j14BJi6
3ew4cvKPnezedUomyEsS7I9jGAYIFGw0g7vzI+YGgACrHhjbTtnOLCjGqyAlhTLc
Tod56ddmp6prJRv62SRkJ3gkuCLOkZ1heW0nYRk+hpwSyzQdNH5L0cSc0tKGHkJq
jBO0ULWkrOjLtlJQ+XE5MmNAotD9aa5288PVwxjTp6JDPOYIbARjrC3EEGl6527x
YKxRTTirlvXWz3VOZWQ5ybIyFy5AJdgyyhhPMzqf7WIbGVFY0LAhP3gzQFDHKsZU
8QSs24D/Q5HlrY+k5hREXNSwG9PbnJzMz9riIzrAPgU5DXZkrA8/ZoUvhJuLd9F0
lgm7XwW3GdUe7yUnzfV0Mwvz/MNnC0mMuCbraitZQvAU//G9XWabpP23Qto9iwme
ln01893keTqDhNVXYuI0pciaWVUhuU8e6/7CCeWeM5eIkrVdw3PO7SUfc/FGFJkI
gT2qw5X63mgXwkakr4v9qinbsZfadJsR4lxgNtW7lfddbt1NrtldRPNI4NKnT+5E
hKyHnwmwdsbBz7UBzH+jxx04CCoLqugHABw4RytcTQ1YEvDVbY8ejTSqYAb3e5sE
cAXGFa1FEULQxoigt50UrXJe2E36wTsz1emoFZUNr7SIbVTNg/66QCnpaY6RgqNr
nFk9Po3X9gspBA6Uw2iGx7kLQg6B5zNCtKQGm9FbexmyoMOy6/cTvj0uepD8kt+Z
SemkHko8yjFGRjVyhhTsABmdH945IL/FbmLZtDRInk0rPB1+lJ/gEMcXU5/5G8va
00H2hEtTNv+Uw2XNKBJLPfafVIKonPAZ+qWXLkiuoiHrwI6ZRH52b0azSVNs5D0M
4XHR+Ld6b0dYUOuvFK0zUtDhwTQM8hdZQE7I9N1+yVxYCMvyZ7sFFIvwqhDzCahA
q5gPyHKpG6weSThfAC8YCPz1m1j6wnSrc30WM10bv4d/6IRMsbah8wp0glr9mObP
sTYwbgMJwR/VEv7tkyOAWb68cQ0RrV2ORqCrDmC1pzPxvwZc8Y0m9QZ4mNy0x6FR
9mA6lN8RgUV7R/YRslWVgSPx2LAd9+nzuE/4svMAojTB0jRtRmxzziUWfNpB3Jpp
ZFlCI4TMnlW2InrlVAUcJeJyhjc5hHGWbIOtAJ/wqs16zS0NVvl0WIu/aPmG7oK5
XdNNifrlEQwYo27hoxbsVd+EeeSPfrGbPqtALVywARGlfVFE8IepDf4hOyUCh63Y
154gOWqPCs0GGiw0j1mnXm9O9LUo1hmkKtpCsle30EEMtTGkNhnrh3/ylUpzw7wr
wTAhbN1biDJ/oEwSbG79E7V0L7xOYSnA8flkteZSsWHK/1OQP1QgCzwfUh7kCPwv
U6Ar8o7s9SQ9XYsVmI3BtisFixQS+OSRP3/CoYoox0JijaK5Uy6OW0WdxwaVigot
MQadB99xGnIaTMkuCVFXe9HCi8hmcD1Hinu+TpYb0KO0oQx6Ip4HC7yOvXF3o/XQ
5CpMuIRE+EROfZ/AH7b5e9SYa7FTnjewUT479ko57l10FeuHnpXqrzuf2RMazTf6
J0nA2E8MAUuD6hGs2VDq5y+PP4FO62EYykv4HiZ32msB0dAMgIRD20OB1gb1029q
QKdddUMqodddbE3bzO7qsgURON2aBdbzRezRH97VmDpVYj1Y1WIXz/oG3Df2/PcJ
GBr1BFrRyA8Mx4EQAG7W9ATeM5uU2PX6eSUq2c03K+d6XZu12UYzZwJBSDIK0bfR
exSwHwGzNWRuXOPAbW3fw7zfCL+hCrK9VczaNoF/5pjOY2C/f/3lP1sRuerHvRAD
ZTwB6L+E2XYJdUO0hWDjj7z8N4kT2ld6v4p+4QYqFFsuR2xsqyIdl5yAB6t5Bcka
kFx7GqVpvcGG8G6f75Z+xCZBz/aoiokuZb5L+KxBac3Hdjqre33b6FDyHWAeubxQ
pZqyqokK6A31A7m57YrYRBFV/CT+y7zX5jeku/tXy9R3DxOFTPIP7l91bs09XgWQ
tGPMojEZcHKQhTRx+/YypjufieYYd/fw37Q0Y+g+Nh7apig1wob+sLC42uC3PoKL
ob+EdCzWicJUL9s6yCCCvZWp7fWAo9i/4oq5/PDuyy4AXAtfGTOA0y9feGvLKuj3
FY95o97Yl+ED76drtSdlFQ9AAMaryrewmlZO0KMyTNTZIsGvUbzv0O6uxlEJjgU7
5XJMrzPrfNgMgSaxdpWNCHb6G7+qTvEaQ46WK10fTZEoDMBG4ErzMwm9WMY499Vx
1ov+eRCFStRr+dXHgTALr5bGPgS7sO2FZKm+beMkzN2laxfPfsaOGO/9GMgXDlNl
KiRs4ato9vXdCfOkxJKizvZgnXu/904e6lqGwqzWg+6g845dJR7iQHwjc3pGqU41
Cry4xaAPcxVFlGqqXoECFQB5zLLObdZIkC7uEyswvVppGoa0Au689Mgo9GKg0r/k
48UIbOg8lXmIwx+MnRsyZinN8E4dWQJ2s/DViqrvyUwckZhEFo2JsOM4yPMzVvxH
8qNM0jr6OnEPQzkZuLQJ0oDm1o19y3+YtTwcM4rUXV1slL0a+pMUqogfw9Rxa/R8
ygAujyrl0oVKjRwQeZPtORhJ9zW1uMbyNG4bQxA2MXsbBwrRltLMTG7kdABi/gqs
mUVVBdXRf576u4X6FAGSolMvO7C5Vbm9mjz8CjuizKKbfTM3K3DAUowKj/C4nuOJ
yKaCA34jCmxodu58uuQ2FsZ6CDGRW3cZz+PIKr6oO4M20B/OD4dvtp/GyAImv3Pc
9sdlOMgSsyYqwe3CbL5jF2XWXxu8bI+26lVYLORMJPGaJTLjfrQi2F6N8Kf7dJxt
8cM135NrPv4p+67j5rvs0R/XcKwbZORfdqYKzzwmGDjxV18LT/bhrywEiHmNQ/FT
WXfFgzdZoSat+XbXd/QwRr0iNZ7pix+XEyGZuKDpOnKrAdCuJ6B6B0btBnZTrdVS
XKDYrclzVTA64hyKNhvk9k33FkcVX0m4ZOrke9FHoTPP9Kwh+xulNgO0dl4lrPcD
cgVTCr8BbBYdzjrOjwUfZ3cjLaQNORhwF+HRhSvriAHId0yoxNFmvWhRF89/U0hw
ra45D9NoNh/vmH4ZyYkT0rGcVsiMsUfaO72FwbvNTMMBbBq/FQeh4P8KX4UyoZzb
fXP7eKTOiHKr6nn1UuWMLHK6AEIBX/PndcxdPOarbCOS5l0GOKWn1M+mQ4DKwz+k
w9k6fvPYKTXDdh1yuuNdbL2zIc6AVmiVuKm7Csvv3RgXjNJXBdtWTQNIl/EGTdnI
Pvs0+b+JFSoePYT/7qByynkTCOTFofNHupsskEUPqwuUBUI9bwJybMNeZ2owrCW0
O6uIExX8O+ehTfp0/QvuWnrQyOrJXSZ4Uk56XKxsZpKhmTF8uP6/pF3WvY90aNoY
j8E/Wah9CI5qJX/6AP0s79Kg3hB+IH5gMVOrPCcB7cWLBmqV4d4WOlsMNLkbjwaD
qZtRjVG/6Jlxq5poRhAwsg+5qysHMLXfPZsOkZ9gwl7YyTF2useah/ZtyjX9MfIf
ttHPYk/R1yEhsULPJhKDmRN4rtXXm0zorSj3ryk74qAj95maI70Xoa3gm7L0JAlE
/iRm/Ya64ONSdljJHdygU/N202a2Z4HitKKUiOnUqu61YLZ1FS5yXw4ffkvCy9H+
owJ3GfvVYmKOtYqwOKxqnCYgROm3k++GRE9GqeBpur7xv+CceATGQI/fxHYPLqyq
t3EiZVGIZr/SzPCvasZQqALZfm3qZIyqK0YrxcyQzsjC/OAIYSVgzXugJYh+zXrx
KfcXOGgBRvBHbtzX8AycvNJ5QDS1+GE33fPy01X7rGJHgWfEztnH1IlooTxkZmbi
f7vgsfot7cGyKarXuwXaIoYsMNP709h/Z7g2IwlVJr4rPFesLv7vIzhKyAlFWXmx
z5n0Arwp/m13pLHgrK75LXL2QES/ZTwUtHSLtBtK6TdCd6r9gqhClEOO2iEYEgdL
ZkjkRNW5R4b5gR0uhD0tAm2RH8wAgJMAa9opRexulnQi8SmvlaRLQYT2niW4Zu37
A/3XyUZFcnTEOOPvCtuRE+JSK5/204unigGf+SNBRWIod+ZptTy68TQ0p27nuNAN
Vk+Kw4vcUj+gHazw1NnFk8H3c+z/pWLUZ2MLtiXvLnuHSQfHXpPL/Zm078BzH7ou
1NUr5yoBK0YrZeQvcXjrXWtDWryShZXwiLUDT0wq14VoPv8zOgg8Ior9+RHmufIj
lLkLuZG8BM9r+LO7Y8KlZwfrr62N97krbCm9mOeRU1bMv+AuSzUQqFu9JAEYL5YW
Ck4/HaaRjvR10D/p6RvYtHRrE2C9u2U1b0Z9QxjYyIZ2u9B7qJw3bTjlnK7UPjCS
TuAKUptkB4ivIPEUGyZSXcmsXyh+d0w1+W0qSezgZxCyMxnMGLVWPzIoVAGt3Yun
llt0ve2yApxcvPXA340gLS++41FxSzohNnVZSQ7IK5VQCJfI/9moGK//3Rt6+VNq
jiCF3IpE0XVdnsfKYYVzoTsXcZ0ojKaJbm1ZXjOAoBhLTdFYYHyQVWUZENKZ9SZD
sAAIzI67DvTfwDLB91YGSy08AuhNMh+A4PgGRuWZ4VuEvJNcSdyj6GM+2nxgXs+W
leMVR9qyaGd7DHVn55F8K1152j0BRLUJobnplfycJywb7zA+vcdZqW2VLwya+7qf
emoi8tvsCvT/9RiGkcpbFAN+JuCXSQakJFx9rTqAdeZyyBu0vpq2xfuX8NWv6bIe
Nj+ydyDtoyqsWRASc2DXJqQEvROINWdXqxGUqiERepalntA5qsAt2oGzPDU9wmjC
nPMm49eyLMR9cuaJ6TU43WIvpJd3s4Fwlx6+gA7RBzQNnsv74oCP/olgjk5NxlHI
6Bo/sbYFFIgci0TinsddqC6Ocu/hHjIQC0o41Ewd3+0dR4go0hShIeBjzqJARXOl
7E7pwrM+tfR+j59DMhm0H3mD8XgUrFfjFqi8BvoMuK9G2sjBN0L/8pFgwfhnclKp
Vt5GiaZpRdnIyIp2Hce/jFHfm3WjRmF/wqw5/w1jrZqoJo8r8IdCA8OB6bKhVzZu
oWhgSGVKuWKW99olEPDC6hLGC/aG7fjCdPGicQSNPA6UM4bTdg8f8/0T++MweBb/
mAAclkeDbNxYKqjimUnD7xc3quNgCXgZ9as0PyqcYXQjkKTzhUAq/u0pq1vbQYMl
XZ4uoWhJS8Q4C6RzP2xz7HDJ8SCiauOt461J6jm1arWVdUx5VBKnGjBsyVDaeOwi
uR+dTHOhU/Ynct5OPZ0sEQxcd1miN9UunKmcPJFHex7OyGN1v1+vyMFVr5C9Mk6Z
/9t2rbg6vbllAZFMsng8lp5lz5REmTNKYNq+M3pAjtRy8B0fkrL9y87jiFDGLt9f
fpRtB4KFV62nvBvPmEYKpyxd1D7My2o1YFTUaVnFYqgtzhngq7UOpez0n3e5lu/y
AHkL1jF2OWdgADjLrKn6XGUZpJdEOo+2ZtCvb0L6qVZv+sxdo8/ACF2lO8IOMcpb
fMy2cGm4XqKzL847v8A2DbH6cX7N/d/3v0GnXl2es9wB6yMaAcAfjOPXu0l4HO4c
BzpmfJJaHKS2BwlCRWpqONfnoElBS8Zekir3y+qbSWjZK64TX8XgkJn7RyABkEdv
T2TkeQNNC62GCaQ0zcFGnVeHo//rVgg9/jqJTJUCbfdfRh6RnpHM9391Z1QyDztv
yBMUh+qMUQwSV60k+MXP8FTwEkonfkNNJNT+sI2qK73ZcPoqT5OthFqPTSmuA61g
awerP8jGlfyXz1hFwo6lBMiSSLsW5M3WxrU8x8XigOzH+SwQy7LDKKHFJ8bS5GO5
EF46SbBS0uX/awjDxixUj4fY5RsAOby6Jgd6DYC6u84td4EQvEG1QWv+jSSRF24b
p4hrNUxcOaziYIFekmPaA8BX3eORtuTbaBrRnpnWYdh2NxpAdcRynVYIPtiESC4I
//wRsumIIJ/5YMQlZcuTLzkFRhBaFNwHjb0qqhPFzh3X+3AKr0ivHP7n3tqnrMt/
ZeqO3uGGe7SwKtnNtT11Bdl/6bdfpl8JTcobxqTLHKZERuijbd62JuHNtrtulj7j
QiosW/Cy6f5Z7cjbFozfh2C85qFwuDeKJZmu4aAesH7d/mYes+tyLXb2kNcpP4ow
wFSmvRRavDdrzUToqIRZF7mlut7vJTamawjhN5q3FwVoKeTdBbJkGAktRlVGrhZD
SpXeOeTSl/MHDkYnsramLrbmVApQz/WynRowEdLNPT5kcMNPv+Nl1KdkhSdCxo4f
RuS92lYSw8zyqFlhtKkHjsnHVfTeoSAhrKdUl0SzS0XeKkftxHOC1iBZohU1UpeV
9pQq5nimroK9z99bZyPys2i9Q9gxusfOawkIwiM9YFeBUGUWOmsbyHiBFb6OfW0a
lU2Pfhx1u/m0ZWcDolyihxkeErDms3wUaKJH4X7g9X74lgKUYDl8sYJfRKYEPuPt
+k+1SfMkM8eKPHHyRwgu5x8DLBQoLPWux6BUyPmRTVjp3TfRWBtmhSKAYxOOYv6A
Kp08l/mLhlI0v1P4Aw94gaEOR0j+qmfcw9Xpj1PpUeaElVuqxIiXHKmtU+DYediX
DW5m+130OiauFKlkz9cjsMT6oe6R2DR2CEPVhL6RNbZR857QZxwYHXRRGSKRmGbJ
h1zfspsjsKowmqytNMIc1HYxWpCzZoC3l1iTKdAp4/wPxWrNoaXxU5AzADU5PxVl
Jzrh1xv+zsUDql3IU2VMowCmp/ml6BgZlNRElRW86pb/EwRSS0r/8GWcdDBQ0FCZ
/Ml6nbX2E46KFewha2DIM5FeLDf7f5G+oeW1BaBqrwe8MvDBruq9XfXByld79TEK
XQL7WGxfkYdaev7p8lZIXAfGmzHl0uucNxp5MGOYwO7NvxurjE8P4SiCZZt3e7W/
0e6RVZUFlz2609ejy97QrB6BLr7CumMLlBhngkTInGhdM4GAB9iXOqOsLMNGI3xf
HxPIyUdbGC2GaDUZ6+lVvCe8vRqCF7H9M1OBAPiKmzXU+a/zZVsIIvUa+dHg8pfE
JjUcFZuiJOjI3722rO6+ahgUXUNZv/pD8g25EUC2+Pk4XC0kKzqIdfSs+Q3Wfk6N
p5jdxPOSwLMmQvHDSC0b4yPclexS6PoshJX3iqeK+JMAS34Ua3A+Lji/HpiEPYqj
qoVeFIaRS7iibWNrP7yEjYwkF4hB/VCS9H68vD4E5iV7mhTcU1z17SQF50xzr1fu
LcWdsvJnVbX0BFxTY/sag6uIUbxFtrKryZUHGlvcDaaXHulVDDTJbsysODylh8o1
UOOfEUIJjONLVD6ohjN+WuhF1TGGeQwN/4zKS1dRbiSxTfBlqR5emal722XPhxVV
ORRrYz1gFQSUn0inDRA54MhBEbqieZMSUbJTd2puiqHlJ3u9pd3hS6orhSnmapRn
MgsGujccsEFQwBxH5E7N/dfLiYVCbynfswvrZAL6zeXkLla8Rpe1kq+Gbpfv/2L6
229yGc7CY9wJkAUiKkSx49kdtbQtO72tXx14Y9v3TvDjzSDDYCqy38mzouieyNWg
B85+Hn2HPisOJGQ8N/S3l/TCzSSfIFDRePEapqLZcLUZ6MLQBzenJwgFuhFJhw3G
h2v1jQM5hVq3NFbpgioobPvJAUJd1QjEEF9mLRxHQvVn820wwZ+nnJc+03mSTFsR
fEUOGbyhjxkSxpDLs3Mle/BM8WwmvlIe12bceKilRkRISKxB7YFTe6KeA3pdPMst
YvyNX3nvvMOmmkU87GS21iw3oPpPXouiAaMYzpMFFqnjeP4xUsuVEFCRc3YGVe3P
n9q1g1DfZnFA11byIWFtA9lf9NYACUYedqWqwRDEGPNdsNhyVVs6fu2JxttsZUJo
K/Syh/eVQElYWeqdnWjzgGhjaq8iwjs4UOwzWYrTy6CIFw+dN92pDefhPCys3Dt9
KX4fwqfiBeRkKtsaipUFVXX44RhYivoTt6MxkGVyohPL1Y0qvnuZCpy1A1/sjStP
Dn/gwH6+Rzc6R0vfc/HhAi/LyHPLGoojF0DkclZ2m2IG21a1qvZtJpBDrLEyUlsd
hHNRI5K/szLzKVVN8hoIPSGKX/EV3r8yaz5qAOv5mIm9E/NhptVZnILg+fhgs9vE
GU51YF5Ev2O2yE+q9KyFRmRD0X5lMXJprbfxJQG1O74LiyaSYeOxmLiqUnIkuZYb
8r1UI4O3bzh1/cS6eh40/N2qz/ohieNaz/RovISW/nA9c4+2wI2vunH3o5ohar2c
FNcUpp1Szzchj1MvBn7c/TVUrafGo81kfLFoqeWT/OuCYyhBEKh1GVGmrfKGVV7P
Sv+QCKZogtPgnNTEvwEclgbRYF6y4X8+eXdDS9dIOTXroQztyZlq7Sg+dMQRT/lg
50inwSvdV4U80S8G7ekBdUSMHgiG+mWaBx7yGeDeAdOrdaUN0jdciunMC20vJPmW
EBpVXxmZ+/TSHkaKJlsM8oxY0we+wRTpIPHVeT4WVJSKMj0Q/Gfatz9Ra6tH35Gp
uktPIxs6G1W4ZIK7VPm905dcrXtSMhZje7y7PxqLvPiQQiefsZVDS6PGSxVaIERo
XVhHnbJ1Whn5WbnfpxYuQp42ptnhgtkJyUeGF8Ye/Y+aBcOpla4E5CWiOVpjhUTC
bI7qKjSgACFnvmGySXfQY0aOQEnE3WHkQ1opRhfnXk7n3qHTT3hpiwvWalwLF7Iu
uSUXt6vr7M7sorRFyP4I28bAZBkY5MQmNY6aSlZ1WmV7HHgW228eMrZHG1d+szkH
uUU1nBCe3ng3R7VvNmva9kB+Eyaoc9Qy7BVJMJTZftr67BbLMG9/VPTm804gBJaU
D83qmKYd69ggxtyZZ0e0awcP9XEZINeW85/QPLBW+X+jSCvPsj+xG8rXtixvjx3a
jcDlz7vOQ5gaykBUXUofDSnlRWkQ+IvaI8pgrVbls4BjqicbOlUiJArfpo43Gxk6
/dyU7n+B9we8ojCBv3iMrFHU0DQjIXovE/RMd905z09HXUvm0GWIRkhBcVEEaOj+
8Ol6NaUdaABJfcBatnuj/H2LPinOfvqYuypgl0+OAZBEURcyOM2jCu3eE7ce5ceg
BmmXKrYYLkpxPcSoLGzSeMhfzCJgxhoU6gXM69MPjjed6UBXg5MmZ96j25goEJjz
4/JZPIONUJcGSOKvkrrIE0ummWdEUZcXj2pw6MYXE7l58vOAyz8x3GmRO76qRT7y
pNRmPmsiPvAPei3dgnIRlHbjFaQgwTWQ3hucZMCIh+oAACJebo7v+GlsRQdHgRVw
KCr9nOwxOxI/8NIwhVA3+ivaNhghhL/LynSSaabv4KGDiT79pMIe5byukqrA8V/C
LDU/XKvOlkikZozJAzaBjONKKrbaE2y2Ft/rxtGyleKGDwRUoIC8QcdoC8eMN/IY
ZDD8l/vIyIWIPPKwkYtyQpMz3z+4Czmac8JJbvGLv+Y1hQYY5LFvUzODZFnhja2n
p2KvsU/EUYCKrcKdSoIbDIL3VVexjlg60PWqjPHdM9bM8N+Q+qpO7bNrEcXE7Ti+
hMNDWNtfPfsaemPUHHWFKnufuEkHhstAudCCf1Z/kMRx36MZTe7Oc/05lZ5oFrEX
uFVy+YGRUs+MLfxzVSXx4YxvdGIT/KTqtH8QKgSbdZ+Xy9Dm8s7xRY49TETonyx3
9ZJRKVeGk+XC8hecyJkewQzbqRL+HxtxaJbV2IHLv1/ueYe5ozsO0pDKPE9uzuYf
F2NZ4uYRbEwH1pkCxexUEMBJd6ofVcWciKmsQc/RoUmsaD+Lp/yt1anPxCe+8jSI
e3jLDkk4Rf7rH0XL7hlLdSJNDdXN4AttAqytoXqjGBAr96hgszr48hbv0zyJgmYq
Abh8Qj7MkcJEmbZ7sZpJWysGp+JvvIPhxzg3AIIItOCQxvcv82wTHRkwbxQ3fPWN
Mvl4RY9TWmJOwYc99SR7QXOWZ7PgvSqBRX2i70jXWiUJoyeLhV3JmFJQDrvEQLml
atXgHeOE7iodhYLyimkXGbWIE8g4dNnejOV0/d1EW6dBmJ32yUVzcqQVcplf6AnU
oycLxvrrF7z0EvcPGc2UJ8Jc3oc9oPmrpYlY+22EycMfzzIyOQil75qFWpOXxKf/
GXlWeh23CJjJo2BQfcZllG2NVSxNT+wabuLsEHnIP5rNnGEnOKzloygWdci84na9
pfP4OxxKlPUR+u1jIJ9LVD66kvc/Tzn+Xs+Wivly2BKCSPiHDsw6Eu5WceWj7mCO
l81gMsBsOd7g6h+8xO44fg/BTdIoVDkKvRKZcgkjFKpcU0cJ8CDbJhnNaeOv30+F
8dviO59T740yXbK/ucredBh3bQZWrhwo/8QRYLXTqWwYbSv6YNNOpQ4VLnzrTBz5
8mCf0tHzPxhY+pfkS+9mYLHRo3mjQJEs8X1F3HDJ3Li7T4LIqN7t2PDaAQ0HSts4
YAfyIOW0RbEFcp+Lv6NrJzqs0CDqMUBoyW5ePDVHah7kRrhPqM7WyAbS/grHIFoj
owXSWJMGuPZNLUdcdZeVtoSqZ0kxqqZWpOAwBz9BsRF3fH5Sr6zw8mbov5ufKXwA
A/89lo+GAbQAyzwKgsZBttqxEtaI9PqHnBXDmmkYCeyhfc2yW2DeRnVk4h4YP/E0
qgtr1+HuB1je4YQ0uko9fFiRQNWWSH1acC2awHKrKt0/mIpUG419rHoYsGpP0LQ7
rLUi5iNWOA3Mtuw+yWQUGCMLxC2KyS20SgSmkSyigKjJIq3zQvQI2+/Fhe0GrVjq
2YQSZcptshgbijQgvjHuG9fpk+/8FNHromgccuJtz0onWaKrvci5YunXjTy0dFay
JTAMoz3jMJLHU2la/QQWnu39bFABJqQIMgeBf7g9gwOsuszP7tqcCUAA6UeHqIOG
2K/xkZITWs30lYTgKOVZuce4aL3xk0iHenfA7sAOIxqx3C7iYOGp/6Okbh866Jre
Reasplv9vFB0/RuGZzJKsUaZlfY24CWjIBhLrkQRFlg=
`protect END_PROTECTED
