`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Aq+YLRKLhAkImvhxipmod1ntFv2rPrWxOo/Nn6QWRj5xbOZMzqAidjUEzHa1jo7o
r32qZfaG1R6EPXhsKQAwlv82Cv1VhN7y/CpfdrwVGqhWcseGDN4FNDu4yP3iLwxn
pFus7uwkiRNsaw5doKPmGFKydHTWCocC5p5cNxdJAR8Z6iJzWcDdetzgqkBKTdUh
rV0q0kVof6LTAmK+5AAjIwRGpTuDI82AWxfxloXjcfwPKrKRowKehjiL4YiWkr+H
W4bu4oGYHFI21rHCu8/BCumyxDWQ+k3y495KuoE/PsF/TlUt0WX9HwtutQSVLLbn
KUnhgKwb6OAeYWQ7ZEB9Q/n700T6aV/ldTRLo6DWhkYYLPCiYsaqdC2jZ7tF9zTX
QWP1NE1A9q0AzlbIlaKC1wihkQVGdpSfS9dZHmFwWqmUzFOs8TLfl4FjHvBIlYdA
h0bdO0dZzdhelksTa6RSppP+6VpRxOl793wIExjTY6lEXy6OFp2YZHxj9RWkZ89K
CfcIl5NUwpi3mjKISrKc2nMmm8dMaDgF57v5BOm/FFAh9grEmABkfg5aDDFwiQaG
zjsri1gFn0fcXqv01VUwIg==
`protect END_PROTECTED
