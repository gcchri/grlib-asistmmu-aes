`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Lcb0iwJ2Llhb//5+zJielUDSUZWoeYQWAEwc6V/UcabG1IcNHZtuqA/QHav1hm4
QjqNtBQjELNzhVUB7nu7q1nSXN3c+3qa3GwjKM/rqP8c2z9CobukPN5PoK6O5E2l
3XHs1BwWlNCNw+jUlyEj4V9i+gmAGj1IUpxnZgswh+TAnWxtRPfrW7pSQBEhfoGr
tc3JHfPYCPMemnfLGvc1y3YsUg/5rMXMokap5fDIpn9/tgdL/B+X2Tm4AqXCR8mq
ZRwxbdiVp/X/C48OOLLQInyg4Q1Z7Id4nCmtEW6y4Fp20HDn1YI0cKAUtkocDtqN
b63qRu7y6eGKxzWqNtZrTfTw2+1Dvk5JSqh5+hU0a0dSjY33y19G+OzjBarmCY5b
5Awr/KHRqQMvqnj55W80/PKQo1yj8fOE/yITDEmgQbep8D2akf3+zQ1nD2488qsh
YMHamM2xBRywUgdY53iJnKjM+jtjQhPynGW1OaoikC60wzrxozLVBQOW8/aMLSEo
Pn0EAVfGwPbkY4y3PmGCcSE8+JBUN7YIOsoiKqxxwRlmFexyfXVa3MGHTV9kyRyZ
Ih2oS+8+h80Y7XqCbuWCC1PgPq9xYssGTjRHxFLTRdEPAfvzeLrL/Q/ncDjuMb9n
uz4PHjSKu7mtCh+fnq3ZFBhR5dGrXGB873qrE80EUrqoGFxizXhEG6i82jPCvIu+
7eU9AGOiA3rUBb4BU/Z9I8M6D6DE9fNGAEzuM+bt6J1Cf4s7DEx3nkFPeZC9BwsR
5pckysxIo+jGbO0qdqLXsBXFAXxwRkczl1bEam8w13HtGiUlCpvDO72mygdv+0Vp
Jd2dVKX6G0feJP41evvd8PXlCquXlR98g9LbFRu8r+jU73SId20vddSHKktiZGET
JGJlJVqhijMjdeAlTsCrvP6nTDSPC3kvrB7w91lKlXuqZw6muN+Xx+lvdB0XUxNR
4JK1hgLn4J1AmQGAUnvfVu+InOQfmjzrR6czBkNYG9YdmMA1EhCniowiIJZE9DPg
vKRSR1ZpiuvXLW+N5GqvAZnhZHWks5rKEnENKPqyfT3umFMuEnV6RC0yrIt1sX7D
9RbckMO3cF8fpkySQOOLp8oMB98nNQojcOqB83PKUcMth4cCIjEzmXZn3dwGLZFG
oSQtZx7IwhbO2ytnJLmvg3oG/KClHrdTqLDVmBnemtCxgrJ81nTgLInKnCOXwgZa
PKTDyTAmA1F7qqMz+Bp7Tw+HmumZsda7eN+cGgbjmzfTPcdtZpTBODlu5BkBjXnu
3k06nZpzxhfgKfSACPmKEoSNB50E3SSVOrEuK/z108LUwaFpf0YaVMelAR9+Vlhj
LdUcGJFB+bay7HJPpc7e3EzO3kvk86JiZh3KRAU5G/Gsy9tmqw7sb6tnqC2LgwEg
YFSE4nTI0X2nM/z45dEQa2ycyRZ+/01ZYY9JBeUn6/J1xyhKnvSMPq3k/2nPmXY/
qberDxgNvsnp6s3GN2ludm7J3o6M2n1reCS4vTwenn29wfCwi7hOT0OdCQiftNkZ
Fbp4eLNW4zegslbupam1eOuyQn0T2hFA9Hvoj2qLVLX8GLkirMrhQp441IjuFTBS
BOxBn8+4TMy+cEm6YRFb+vEKf/2jwPxPf+l0CPgecdyzKPEXZE+5RyEKqxQ4mv0t
3rATiMZLUTVA/S4MuYL8UqPifexD5OSdLlo9jDsqVR3yBw3usGSM1Qzpxmu/88zx
/bYXWWXpdT6q4Ot6saWqgD011Dn31c/bfMS9ZfjmLW0FeYWVJ+R0htyrtN36BdTt
nRrb1Eoz/bTqpphNGLsf/0WNL+sHk2OUaKFITDnzrwYKWaB+W6gidzwRfplJOlnj
CuP8/olhsLMsGqxcdH0/MOTkcyzSTDzEvADr6sktbSj0dvIh+V+7+Y9vtA9d5pWb
6ih7cQ6EEbLykULuvTBVmLEAESZdRRdf/xk/+e5w5OSNNP4yagjajRDgOYtbr1xs
/yfUtq5kg4jgN0lZ8zQbkUe1zjQYrpOFujbzpNZsqxJSSx+FmHCBBPffeLANEkCl
XeTq48L5xFUcf2Aqh/yNxZx+byb21qTgCr1OcDx7UtWXypO1UIDq+w0H0nmwtX4H
aXwHQnYgbl1rkFSMiPDF7QUetUwpktIo4ZakzWdmBZC11jNYL39J2jqom3KXLpPH
BJ66rH8UIbRAIPYmxwrKIK4JrvYlwg91yNR5M8pe61t5qXIWf+gqSWTMloQ70Ekm
4WD8ofBf6+FMlSVeB7E1O0uhpIk9dH58TK5uLsn/O+hTGlXxu4breEqMmD50gZjE
ZuwEj04OIL6Ht6fXPjHK6txSxsuX7jdPO+5y4KFDqMYK5RJpYesadisC09DyOyuf
Wl8Wteu0fDCykPzmoG+QSDCac7mPawgwht3zqk7K2XnGvjZC7Ua9qarmomA6+651
xNECIpNpHNna9qDT82cEFuoPEjaPDlLH1cMKfi1UAgSsIF/o3JEI4JEKxt9JBZ2d
F9RkDZp81AoCZpuhUcApH57IZHUnTgaLvMT1LOOOCdJtBx8kIJiMaHhtpfYzOF2F
Xonulzo4GISeCMAX23rxYa2CpMpN0oW3jabWpX7ANs/SBLES2r4UtDOGhBFMmsRm
qxCO+FGP+RwWYk61WgMoMzFW5Cmw1WgqNqLBg78bZF9Vqxkyh+gtJxa5NLA6KP8m
CiqgLD/5rMrZUCQyMlcQ6nACWtfzKSmxeFhsacgrJausWp3/dRBdkp+wsThMYsLG
Y5P2xo8+SKn0Kb58+Ax6bUkgP1b5ZfmCNxrWkahSKEgpXJJupvLR6+kPW/42WQ9T
z5W0h1UtiFHB3f+/2zLu+2dnZyyO1bN83b2+AO2giKdqcuaK31t6NMZtPunylph1
t8Nd1X4HLbuuoYskM6dhqRJEP17aBmN7Xf9dEiCNP86drxd2CkunsnGJnMdfgJiL
GqwuN3vhR6G179JlRXedQhKwmYktu0m6SA+oId1ni2kHxMDr4CO38eb4ykPcuoCr
quP+8XyydCZX7rsZbE2GF62Q2QjC35d2Y/xdDpv0auZKoOtfbBFHDTsv87k529IT
BERJgoJFMk/RA2/ekps318OHh45xwPY6fmlnG0WkRk0fR5ylOmO+7RUK6ULCuBeY
hnc08HjI0A0jduQcUQxiz+htXjNjOwGPHFZeI27aMKEQX27arEl5v1r0XXSfwhhO
8tDYuqxrScdq/WokcQmAbbCP8hq4hG+p8HX3XuxnmujNgR96MdAI4/fkJDZ3cHlV
nswmu0yZ5VaSt1oylUmMrQmPcZlV1yT5iIeOsYYFaMEYT/JXRxy+TFncS1gGnazB
0yeg/6F/IYGcHjfuW/NrOU3U2AajvboEWMaTzyLG5Fa9nrFv+P+uVnxAkMG3xECs
1eEIUFWx3ebTNWNXeecga/b1KPXZnIL3ROekBXkNtfiqmiL3o3FDNckklM+Qea3T
SBTh/iqKaDoCybObTGreSVlRfIZcQp3xN16w9Zny+nrrjuRTVVGFYA4dBIJwyWsY
oHg+mhIqEApESAeMi7raS1l7Y+/U9E9ttjItK772rSTLEaY3LwpYqRYFF7OaUfHX
0q/vY5+mgqGmUTyI3jlAZpXnBGXjnn0+EGy2u3MVRti3zWvqPmtcHC48xxeKZiyH
W2Z2wybedMSxf+VOBnX51IJkiAAQmMPqeMsyrIzBx5n7jHTPjCfelq85Oh6ojCic
tFRk6yd1F/CicqNwwFPBRe01OgmpHLrQqQdQjaM06FGQSkuycb7ZktY7LzhtvD2V
ZtpeiXWpLxTnTk/p4KIpVTeZQoWWgAOVQUxKqPTCswMbXXsG9vURYIEVWrmJlnvH
kIL1OPNWpB0xdL4dcQk3HjP0n9KnNoTSdBNnn9VLP3Vz9FgqCJ8B9fRATb/u/9gT
kkiHbn48iD1gTznjW3MA3dJ2cdu0uG3pTuq9f7pwlLQHuc2rkT7vjroqwXTmd1uU
6Sc7D11o4hiWIoa/+9RqUgyhTE51kkIh5K9czXhPOMt8kCLsAE+k6Ra+XqEG6/Va
k8dZsFjttX7Jwkmp+mNwjJo9IV95f52CfTV2oPGEChIdHf0LByxk+tk3HHvNOynT
uaf70CHK+baUiqGs+zrRWnHYyNddQQx3npsvq+vPZCs/8vCGP9Gez8VsRRUHr/Ze
qcOW51KFUmG3J9G/W8F+sEXc29a3Q8rttsv7QT67WTiMSrkQ8K1pkCC0R53WJYIT
qZNf95HLViJ64xK7sNwAB0g7b6mLsUynerYXErv+j/mb12EG5/86QyEAaBlN0fhh
V7287Un6CfQPPxpic8Ip774JGhUjDj5Fj5l60jPqQJsAoyIhRAEdtojnm087FjA4
Nf3qAWVX8VPHAA32qiRt4ckgKIGH7XyGXCUp3h1dDTTlYtrvJzeKqLtXSglpMwa+
0Vmz36Ap7Oge7fB2oLmNeaEqtotEohZbQ61I6EpazbvjOF1j3v0H2/isgSCIKV8w
on/Wb+gcD/oxeJS1L1/Dm/6jcgvVQOsTn1oL3/ZJXvbLZAIOJjfIGZpap+0BA15r
+xc24jTMSDtUxYvJ5IFBrf/pZuJVpQa1+Xeb/mOkIknq4S2TsjGmJMKvfifo5NtP
wbRwduU5Rs3NFg7uvmjmDWt466ln1lPsDTzweXXSXz2yjpAHGnJx8uyTLlVFibfA
Wky7853hdYC+dVrb6OXFhHSySnvB0aiUddhiQnB1RbbzzTFtvdtXgfG8d21Caipf
czd5KHmdnONYKymDeyoDDVkxb94aFoXgkV8t+BKMrbzbHuVBKVMQWf7WjNt+sCcK
DWhBj6A3L3k5v2UqaJEv+536UUFZ9eZJNA+1hltlUSJ+wdPuv5RYWgu1NoW6LcAt
sKlb9PTQccqKbyEJ8A6o9bLkJYxYiwq4920NJ/0lml4kLVvtC6A5cgyXIQHrhWWp
LAeJuuihca0WNldeRbcA81KRH/lxDq2LEcgaq7Rtc6kbLFQuwAUB2hwZtYuO8Frc
a8tTa7MZNo3iiDf6UKU7Q9pg6fybM/+nFpc6th3D4uujt5AwBdrK+/B1lJQvCJw2
WKpdkpP1kGtXyfST1tzWbNC3q89KLkJnFUwVZCUrjQ8Fxy6Xaxc8xMmU7qpj/zZ1
u5u21DANoQXVY/8p7PyTloYWCdtOC+zIudGeATv5vu7GvfZLs6sIfAPuRPNiOiTs
Z6ZyYiPlILZdWpfWHZvbYy483MaNlGhDAILHmt7CiESgzBixY/s3m1ZB/dSon0G/
t5ef8ojcpvDGvruVHLjvm7s38IynLeBG9v8NdC+mMFV451YM9q+upFG/peITEe5q
W5Z7bJaEmA6c9rhTQ0iZJnAyF6g2d/YINzzrr2S4Bl6oODYPhHwdmcYFzdAVqC7y
AG4XjzS9h0grzuvviS4EHT6Ofp18NOSr0HVazPbtnylIGQmyQHQDV7QqswKtYXJs
lcnPrSJj7Tbm2k5dUSUvBMn2d8CzM+djeTdLdX63r4x08qbeU6E/O+XA8p5YrDDg
GvEqijtgkPfjZNb0oueKktmra63VDbGBfbBVz8uy15/gO3MYNM54k+0RrWBzpul5
GLPSGqrVUIGiqb2Hz/mvDVR9FqK7wXdEMPnbd9SSbISGdG+Fcg7WkUpKAQhZIWBz
0t+Ie8uc1jJj0mUT43Oi3OCAsCMDxbS1K74vFVOy1ZGbY8/w6Q2GPMc3njbAy+lm
Y/gzXq05+FfSFszW387K3Apg1LBNnPCwf46Xq3lZsz5WV9B5xGFWzbSHPZLsSOTb
ioBF0Zr0N3mBCKOURZNSCrzebKQX5eN/4f4IHFm4aWhu5x60MUTVq6t8931CcaLB
JJNqrTmHObt46HT5cwtJWX6YcKa1qneDe6rDpZCwKBprZM/kK6/d5hTF/CJg7s1a
t87Yy1VEaVyvcU4rUKoaFoR7pqiQ8+iMPX4zcvbgeaeS7Tc3ykP2m++Za4pHeP/r
aFo8tVvUi5YFl161CjWSc+uTaatnLOXvgi0Rw1oHw5zlp/N8ANXHh9jMIJJH8NHS
OD2NnWDPhK4SjlXYgQenuYBJchAFi/Dr36SsmzTHtNGHbYddQ03V0qLFifC1W3/0
PfWf31ersmNfkyVF4CoWAgFbtrRPIYLgHNKvVOVox2zZwKb1c+oE86/PTvkIgYJ9
T2j2m4p8v4m9+q8FXAW8tbJj2LtYMDhrGCVE+en9NLJtR6IiVVJLcZ4DiEoBFufV
ZOvlrOglPLaQE9OXN7+7pzSNfrJEdBvVFbxdsdXhkxOGUZpKXNnAEsnswLKPDVCc
BAEexKa9x3hwjl+cPbTkCiPrBpkh+YrnqT21n9q49LO+YjREupbF1v7mz4/uzC0R
+BDaPNi355UK6n+7TJ87hUkjpO7X9ogf1Te30GdngtFOzfzrI6vhHbUlZ4WsiE1z
CNpy9Izl+3bE2xTdiQ3FuzLrTbq80c33zq/5q5PRojhw6ZGROL+OANTaT3vBH2tx
Fkjdu0RJ4hGDNvTQKPJwNm8aJTwZOf9iinGRhyYOCJRY8mxHzbSSBDiXM2aGcvIU
eCm8+fIB0Dt8iSEnROwG7VZrU6LbOmTYHrQzgrCtSK4B3ZuxBvjM223GQmf9hBWA
/RJex6LCDDA+yEbTxBcdfiF54aHHlEx5yryOfGliHE1hbXlbQ9yAQHJTcr1jubGu
A74EOBWXoxXq+6paQDWykEE5RgbZKJrCVtLqtRW4PcuecdL6IbCDujZqrrZSuPBs
dhv8jrsBWLUW1dmyjBtxh9Psb3JHrDGIy91qnKbb7HDgvJyofDgVg79gNeL8Gxhp
CeX9drv3ZLq3ImWhUOoeQJjwdMVjCM494ebr4IVYoPv7cazULnlPMF86QwnVUz59
zKHPUaO4NpYdg2y/eaQWgiiAbXzt9RXn30dehCiY8tEz1bLpNvsBDL7U/iwboU4R
kAwW5y3TChpjBkbAEvCpC3lwo4rcUTMHScpQmgxLTfbcGt4mjYcGNpLesOeUG5J1
W5E90Zb1bPVWd7T9f5kcNL+DOMGOgkeGE+XgzVY+SgMXO016NFbvL9V05N2N4Sin
9lMIP8H1kEnQOB5G3SWLwfvCmeLGAiWSXgYzQ+j3yIvO8ultQKiZ/H2DUaITPfor
POB9fjuLW9xTwHTTNyfqUMGeYbXyMzyGuiV3cC8Y4phej3L1dbvsFfO497kRpVZf
7KjnFRavzJUljelaLIoAMQBz7q/zKwUkrwpNVNkUDazyJwIcrEVrBEIkkOc2PGsF
ucZtXLDtMXemt2diT4HvjfpIBENm6FoL799RUEnfvOdQlAmgjSlxXe7MkRGw1fs1
7LR6mJn6ZThRKxJBftMVjaCIPvgKT+533mHDrtjjDLY/+IC2qOnmlQJvnImcyJ21
e5JV5YEdQcv94SaLO6O8Ou2cm3fzDwggRxyeheHiu2zOqCAYUHOUj/o2fMcmZKqQ
8eWUWgKEQr8rijTjdkXXX3iTNE/kHU2tX5qMRHHKtd6APBa8QwKBgrpDm00NGpNR
IvVCiIxDBeU7prW/dyokqjJoStgEsLzF3o5O1NwI+egpSlPNpCo1QE8Z3g1ImOHx
0YnK5EYYt5I6FENmwUXPOHFvDP7lJ9rXNufu19nP95TUM5M8OmcCzf289eCa3zRW
jYFiMV1QcTfooco8NFNY3SEkRNeQ9xx6Rs/KDrnRT97VYk5XD7EQELILtgDslHaz
FtKwYgblQPuJhXuk7hzb3xRMpCKeBJv8sPJfEO4RGpj/SOHdFvCceLM6cFk5TG3t
KpaiFU8wL7hBMA/7hbKhqpr+URvNuAl9SMyrEHV8COMoxCtsmqRowN458BU3SbzN
Lnoc0pdRYaEX15UfL03mQndiPu0xbsl6QZEOBlCXiE5sYikbPBlVvQngG1qld3hA
khupblFN51X+iw3k+q/30FrFlZErl7l+ss6pLkh9jt4t5oPCq4a4oVv+Vmxrr4y+
H/5Uz8P1j4Swt/ASUg0RyIn6YVI5mlU5oZVHScRFY2kYRFUFrN3kX+lPelV9sbkP
IwdbBwYvsDAitRFcsgxwJ3t86JlHDxP+O2+yYNMGqpg81QSdlCu1/K60Oh+J0/Z5
G704L0rB57AFyqGHbkVJIcBBOpFxXqr8HPeOeFAvXA8ZuLZuMcaJYYc7E+7kIBxh
iFljY5YUWRYjUfKfuSbxU5NUNmvXbWhQTrEC/Am+Hk6jL1KhBGJwIswjPxcRfPXj
Eed+mDiKNgv1HjHGBVA02xCX0/R4vOUarP2ko/CNkp6wNf2FA2vhmRKGhdrEaU3Z
NEsf6SOSBo8TIBDin4kwX9mjAeiu2doxcoUTNh0p7/87RUM5kpg2gIzbhUwvvZpm
H8lNThWRuVk9w2lHX0YoTqLupwVzmzHij94eG/XT6gEd3Om/blg+3F6QpkNjbUBI
2wklhYT+6EYdrC8obrYqPfulzOBbBYSr+9Ah7O5DNQd7nAwYY8YSpUfa86+3AQMF
6hRuuaXjc0hGSjVBPdQ8D0VXhqmMmRFcyngdCWvAK1NY675quz8G4+XVoJSakC7I
PeXeTWMaPMumZM2dCxI3kOx1wfrW8s8VQrqC6jjXwry44o6IrILQOX7R3VfP6nhY
igz1lvOwIbutQIZrvj+e1LclbWV6eHl53r7x9kpr4WtrcJF4JRBGgO9UvGF4Yo6S
owieg44cLYZ0/wV/tJ807+Z650jhmNYDV4ie/NjsNkWxXZgc0Kb/9em28zWyDWpt
tqXKEJIXl/Gg3ai/FTY68IKFI3HkkscKAt+D3skPBx/miAOQY5snzqtCOsV+gORa
ARWvmlBArHbliBRkEfXixjQoNATn8P0NgoWp8gsye9dXOo/qa6ACJtzhTd5IppfH
k0/jvlM6x+JyvltKikNaATiH1xUimsco8iUmb31I41rqJLwmtPztmh8P8iNmdKc7
foRwRPScMBIDQV3pAsTn/+uLMCoWQfvtoo2LmeIf61uHh/ye/9twrdFu1a7dhxXX
10qVzuRfO1T5sqi+jLDgoPNuTMeKy0Jj7ybY3IhJkM+/OZxSxhaSe3VzlUA6Vde9
oygRPYSGO893TGMfFyrOXQ4h/4WsTjfE0uyZGrLYP5ipN7eOsSJNeVOjnw9/fjEA
44b8MiiFDlSIqzDU0OIMEk30l8rFQKBZhKlbVO6a1scytpkKn9sLTYAcbYNCPUZt
uK1XSHYaUOahaSTcy15hVtuKthTSPC0QET6WdvRnLtlnTwwqnOhL50z10k3GjucP
6/lTs42L9UtK5zYCTUbZ5iF5wBfEb8bTQix4xlV11hsJCMCwMRAnOT2bZh/44bNu
B8rGvcDOp/2in2G4+9tkPD/nuc8lFAxxNQ9ee2KZWiYavw7UG33E4627iRuACmcI
rvmKUYsrwpok7RyT0pppGczXLpshcStR+LquMfFObI8bidK1/lrNswMPRziG2dJm
o0phGoXgD2nUVKjmmeata/gNOXiWEQ5aVWUeXbaTjjU//Edn3NdPMT9Pf7kWMgDB
nWEw8eAmx2Us2y2zUBAKJM/KW5PcSrKK4flIp3GXRrCyaTPY4zizsQVTq06OEv6H
fIZC4dYDSdkZScXoP2nFQ1y9Q/v8LqZ4lFMQLDb50Z2+4Qdy0CVfSw9uaTiaFLDM
I6I1SelBwt1gTwXwshZsselzMV5Safj8XxsYYP6kZ1JFbn3qWEIDArPA27F+WOPD
DCRCjr035by3Q5oi7RTXJlwqTmTa8L2H8Jn7On2U6vuRr/sQqcg1UZTqt/HC/NET
mYO6dk+0hs1ytd4tvAGnCy0bghKZ+onAzk3rU2Ke9Dvu+lDrLFK3SzOmQnLSRem4
elNcHX/PP6+7a32ElBNNv02h6IUNwbNZdqw9gjg7405aIeKb176lkwbtN2wbp0js
LcYi8hpNNu2PdjYiorJLhT4Vsy71162wiJOb50APPGoIxktYx0RQJG3dDBYmDQE4
7kql+O8RmepPKVAeDIM4wdwMvgfo+HiKjrniwp2Nhzi9C0teNsTDbUiPEYog3cjN
2+5nmOGq7opKzCty1h5uKk4ewF/E1221BKEXNMPtzD7ByExEPCUyYG2aUrpfkUL3
a8fk8dDbwyfcmwVwF9U5FtSEAgSvvWJh850foCl58ANpHO1N3WCLBvDNe5AdaxvK
JW+72467rcvcM/kFdA9lrgkw1UblUxoftrORiVi25UlQrLSIrJ9UnBFM2dXo97K+
y9YjN1vE62N8Ve42ZbIhciusiO06ptlVbB+invwyju+EbzwQP/IeAXYG3Mi0qDmz
bUDmsRpxqgrtwJ30X9uNLawV8VE8/hYtbP1wYIKRoK6vJQXpH4HoCoTbM6vgaQ0+
g8XsCPfdT5kuQdvwmF+yowNedGwdihOD2ADX1Xy6ZyjQJn71/FxSTXLM1hsmZCes
2O8bk3lPR/6VcpW7pRrmsAh+EwubDNN9pLWeMwgEEHzbFqwV2Mql2Sxgm2vvmT0m
xokdoh6iWOtQD276NcMQg2Rz525pkLbUaUQMbOtepYNbzqxfJneTH3fF/twajbbm
GPFpBndEk2JiKIskaIa+1ZLTWAWl8+TjPkvSdx1GBko1L0CEnyIBroADiVGUeKFL
59e9uh3A2bggmvQlUmdzwyOib6689XU8KNlLkX0qkHphfIrJXYGJwnR67rnRZ0o5
MlIdlveO1gnRihCKjXy48POngaJ1zxA5MELIVsTS+p3Wj8k+coj6DnmkMlPel5R2
2QL0EM9s0Ka7HamTKoBhq2mM4gXhxU2hTaMIr9heBy4AfE61oMxSwOmCsBCnIGt3
UnIxbvmD76PtcubdsO9kuXv2Y3uozI28EMjntE1Bk+67mVdOEsuxeUubw7k2kWWl
wLOOmxWMs5m4P41FeP6zrKNTMglakcgUZahg0uBLOjxMSBC8zeZq02bh1i/QtSS9
a3oU/3Lw7kNatmy9d7qW3M3yeRDCSWPg9LoBYp09ChiUnkPJ1fMvybcNlW13W9Qj
2JwupHJ5Ik1CeaX8NaHxnwBT7Lat1zVJAsekkJohI8yQVpTuBS4MSR08FOsWLo2/
d5C80ovmmEV/PtJff6mvRF6s/Ec9Xy2uaCOJgnA85YbASVq5x5OUDvkGcpJMPC+y
XJg8/Ls7ljDMxU1WX1qyqElN0b6uKsM1GL6tV87r8JZhx/CSnKXg4l/ZLuNz2Bf5
Ei2OuJi2xmyqoZyIVqpYFJ4ijQoBB0iJQtt8HICRnRH9uhqZ3WUytzbQAQw3a1Zx
4aZV/bBsttQzWQ2isl+8aOQVTr1k4PlZBmLsxFIsv7ah0G4lU8fFHqeTriByvBmP
`protect END_PROTECTED
