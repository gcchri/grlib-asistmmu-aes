`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ov46CDG//zdGyFQsskjBmvOFKae8CAHpnwnJr1j7xTCKnwlNi1kGve1nPpJsksLW
5MkkOT+ATTbOg2V9cx5WLH9AlPWiKYwIKQj65EGiH6RkPtU2rv8QBECE2VkG4pBU
T5fltErJ+6WgOe48eqziPkQmLqUWWC6IjLCFcSmcZ9zKRINT1kB5OXh08gII6+DB
BnAgpB+F790m4bxiiwVxGAvQtxbItJWp8m7Lz1i3OiKOIJxggvbXygUrAUEnEo2y
PdnJxI/TuGv4flivtc6lC4yur0fpCGGmYFMvdn1hE5cwYSiaFD6d5JOQva+zZFCu
QzMfjOfZP3qvN0+tXviXUY2OcjviRq48lUi+8xvx0W8vrUOmR4xb94DMrL8NF/5o
CXNynp5m4LF/szqCnCIc1H34e4zUGm6kRA2Cl8Z5+PDTlKYoi49X5F+G8H895F51
xvNF+04QGfNRyKyL5wPMcBmpy12CRndSbkE9HxmgKJO+AHeIyFR9rgaAkyg6OCz5
rqVh7mUtJgTyE71/TWQ33c5uvhTzyRu3ZaQe0i2b+WUeTdQBkPCK/mxXeMgKXbM2
dfOm0lt6ko4oOCEGgJSgfu1QRk6YizT08BXQ96brQEcUXoxuGG7JNfnQIQN1O0sK
w5kF5dBvgxwAX1WWcVNr31Ju4eVrQkbwKLtWfs0E4wQodyajdTUgUDQReJJDmmMg
lELuBTyFT/myByNHGvNCRSNDUTVm1jKd1lUmEPOz8oiHhtWrlxlrMXuHhcFvYEO+
7oFMH8+qj9tHtc+WdjcgNqgO7Okw5HhBCUHxRQraixRhlDznxKYaU30g4fKzG3zC
Iq2NWQbfVVrxpR8gbTH13kwPn4P77RX02Dg2G9oKsQq4bWBAiiSii6EsoPt9yede
jJcbnCMaGWxJpOqoCAuvUei6bgPT1L7zRpef+OAWU0w+LFJ4jQTYYziA/awhnglM
3sXsxlI8ZqoY6/aQb7VO6vKDcgmAzwFqHKGKBFTDOf7trAgkPpfaOzeI6NxjeQJ8
tI5pn+hCuptBeEuVZj+uMBqHqCNlwlS47IlXURHVUIOmNKkWu6uZT/CzDZuLm7ln
ernrHk0EoWY3Xs6vVecMlXmpw5FhsbtD7gMPfMHBxl6Y/m3hnx+3Suxe9maUzdSZ
y8vUCsWwuLiSCuvJnmesBki8SzvVBoxS210EPMtoHrDSqxP4K77aa7wIPX5a6R7o
UC8ej/7S4y/6TRgcjxWIlqdVpbHZZzu5VZI/hQAOyTYe3ljfKjNL/Kqbi287ZjjL
uvgC0RRepU0J6/C+iDpCcLJSGayaHl+DmEC2KaF1WFfb1GGCJWyv0kMBehieA1Oi
FF+YQFIE25vK+t8kJ4FUbpBBZARbsVDbT8jNQ7DyyowAidbeQ5I346G7NXp1nkTX
vTI+tHMh76/63m0g8O0qk1GkWUVGiF4lj9Nj2xtjfD4foyOlrmGbjgYE9TcjUqQL
Nm+0vtJK/pzamP2lhAElqiooye+jfSX+E+deNvw3ltt31QzUzV4ektsopsqOzw/p
W0+qG+jf6xEO8ehAOsmYuCo5Zds462CShzdhR3Yw4myGLFpdO/W+ispwrf+lCvlm
pK5sz9xB7JbbKXlvPF3j1vnOA/yoFmOHqCqdXmuk5kZrygicKz2asV76iJ3tdO5V
HdW7SFzTHA3McWNGtA3x48sThdYGEmV/pu2rT3RW9rWqQimk/ix6P/SuPSLws0w1
lGP/+d24nsoBMcZOBs1QXPkwJ9i15+mcRvkQGwi0q1IGgcChzenNeAEMU7Me0TY/
OpV7JO9Q0tq8X+J5Lv+/tRWxCf496SH5RT6m0skYugTm+OH7UvCnz9LYyXnq1gUd
2rGPkdwBsow+90VgPNh+qmzOn/18BJ84ZX2SHMw2NhpUD6o+tYkvTDITMlXf6qPx
gDlR4FdNBfhN7/1v29qy/TDv2+dbYfhjBa9XD5Dc/OHWgIZFxP+8lZtPk2Z0Ydp6
mhyRjZb95O2q43f9jFEwLMnN1vRsJom+dyJ1790j7GRWIeqJlE6Pqz/yHtissK1v
EH5TIs3R83kQ9Bjy/wV4h/qgMTLHwnU5wls96Fj5fd/aaJAVMWO8YOs+oK1ROF0H
jkc7yfNCqnWnZAKFb2kTQa9Dcw61c8MZAx22U7PLs0uaJiHwzvx3gHGoJ9OcVeG5
zNFZTcOkWElV94CJ0tSYZmiEIXHKYBb7eW1gxSjAjzg4U4tv27kEu6Kgx9hX1zgv
gfAeLR64yYR5luIVpHuYr6+L/kZ9veBbXkFETQvyVdF9lWDmQfmRHZy9hvwfcFt7
Hh5tGIs/yDr3JcCuSo2E8p/iIVYmDLbK/wkyK8s4qqnxtBxQdifFuyB7W3gvxYZS
V7UY7j+gSxMa7Q93sh1YdmPlt6OZxClKIDIPKgLHhOO2m0DJO7AaGeiR1nmq7UtR
Uqd9edMPQnO4siXINqjnAEWOH2c4BvV+9jYzG0vSQzpep082UJkP64zTpM7wzpeP
Z2teYx1dalt6tMKkBRsVjHWr4QTrsC+w1AqHTc9/czbgy0MH+cPsCFl5dK5Vw7uL
CsjQAx4PhdIZ9RfpJ2Wx5dy6Av0PHGsvZRGlGFsvp2n/8hiKMINTTiA/Df+QD82s
0RD04vsvkMYemK4KqsK50cPvNenZZp5/izbuWIjLmzxUPjrYddQyfPNWsHUp7Sro
vnCJyCNMLlfX5BWd6TW3jLPVsXdILDlUvvTrk311LQLt5OdJb97MiVyGB2P+m8hm
JhUUp7YLYflYxJzXmRmNxCo7vtFEHGsXOFr1G7RdxQO95hBaZucsctBj1+XpJ0hG
6yQZ94tuW+OpZr1uWgfiwlIBo/Qx55UYkoZo0JkCf2sDj1Hd3qfqot/3EODiwV/O
BFG3jg6URAQnbeWAdm+jsmDe62sk26i3QHNQi39OInyuLB8XeU14t8mEdpFiGhLM
bVYKfMih/+STYlQAf46R0E88qMLa/I9VO4BUWkscazvlwetuiBCTUAxj/vBH5dWo
L9qH4IQIdYzq8sKPIYn1R2FVqdx8TY7+baBZUMzL+Qn4txTdEy2IuvArp1ZAdydI
TlT/BaHAZWDBj64heYQXUyMrXICL9hAoBC/r1cZWaklkz1VoOgXJ39a1XyTSEip8
L01Yd5qYCnQ94/OMFb9Z9+exlrldRmHvDf8mOBxhrXPV9PdpiRB2eXALKEYoJ6U7
X5SnaaYFJcb21FerpGFiHmSk7WMaY5vcuQxlipUVtx7HW0w4GkwQjRyW6jSwMCrP
RrtTSEkeUrI/3CSbrSPWHDQgoo0rvopvhJtY1BrFFRfumOK/34W+riGVrjRY/oQQ
vddt+C7+7mHeWy2l9/vdD4s3LS38K2cbuajW45D4nVxM//m7yo1Q/vicQsFou8LG
JoTFQoydOgw9yzzqLHVQP5RCGB287sfu2uXfhl858vWaKxkFiH4xfGbMLlHV1wWi
Ahhwnw3vN2ynbpBRdNW5WCBExw/7JhP3KJ+ZxPCaW8Srd4FW8ZIghKrI2wxMy9Dv
Gx6Z5dDSa/65s0DNV8e6K9W57kZ64nyGU88qzKWCmCbNBeDExo7hqhLuYqYHQyJh
l9PL+s93I+L1GLd46vAiIFlRb7Q3i66l+QfhqxdlR1LrQ72RBbwMckffACbDv8d6
yK/Vh+c9tE67kJAHq9sNDPCGFldauBc1/ZYvIrORepxNJswjkm54cMv52Bi2rCUj
ptPj5Tt3g1RJnp2t21MVN3zxt8m6U68hLCAWryzynAULNTL6IWKmIteI6/4eCzsp
aSIP1qeW7gfQ7/jReAKDZX26GY5yYgWUz5fGA65D5UNjYLhr86lFcXw69V/1yQI5
orIRXlnRshgy7OFIYTrIS7r7lP6vEiXQyYRljUUxG3eT4e6MRpGeItXYGv3uikt+
QpJhy/qc25nkbpOhlHzW7sEW1RYT5pDC8ByKjrzGBIhSqqI6zdhT33KMWRhORRm0
Y6tmf+DzFyjiz8/cwUUQjFv+eg6B2KAGcb9C00JDIDc7EsLhIKacCQV77NTg/lLK
sPSCYY1DGnGGC5OEqCaSNkHylBKwf6BGw/2F8Ae2taIgcvjVOnau/IKWpzZ/Y9R1
wF3NI32cVy72ANM9BRtMhJLO+M8wokDL95y1LMJpFc2OSurnJt/P2gGhI2JNxtrU
6PGvaVkH+DHvTx1zhLRIV3TmeqSNG7bvUKyHfjJtu8O0TkCziiCKlXw2azMQcwpH
oWkP+ZYHB3PpEu8NECsiyXUwwO/SEo8ImRBQivlOMkJg+qFjq3WFduLeLYIwOk3g
h9NxiFpxAVosLXjC2V3SW2GVLANcfYonYvBUxVZrLs5yplATuMdgm8r9z/jjKc21
T+M9JlY2x+MWMrRuubvJ+Ma17Q0QNcSjIWtqEKsXPy+FGjaKYClMMIEV2zA2pFmw
OC9OJyaFL6LxTk9qL8+OPMVavj7QeADS0uOAAGN+1FdH/qsyYozlqzIeNPLKQuWd
DHXU7OGA9HH45r8IQBe4TloLUzeAE+sYgypn6Xq5mQrTvWiRrXTxqetdiOR1MMTU
rQXb4A9lMLCl7Y2T2lXLpWUQ+oOrHl25yvylGFeTtIgAJUs9mb7I+lZYbQKFFDhj
hCCy6fyS08By/EHe8Lg+WxAXmRZhathhCVIhj1kiZdhlZph2NCSu8fwebvZd6a54
CgWTc+oj4ursFDbGYZKmSZLhuJJnkpu3D3Yq+KjUCvCCGiueUsNQtY7lHALa+tUC
Rqgr1c2VwDzxNCB+Ti7NMfwxr6w7NGewzCeyznSrVSalpn9V6FBP9s7WYYruKFUv
b3UYWOkDBW9c3yQw1SbUGWDdH1qa0A1brUI6RuXpTchWi15zcCabh+5YY19ugWje
C82u+7tx8A8yvYhj5BiigsJOaKo2GGJLmy499zngvZVv0NHntX2AP4lag9TY6N+b
My5jNopQFM+b/IFunC1dnSGZUy5oCf8ymUOFIIc2KJTfHFANTzg0fZ27NPWZJabO
1H3NdqqxRAXRa1vmJtt5Z93lGVQ/uQWk4+C0Rfh8xc3qicH99HmDgUiWNm3VxYa2
j+KBPq6ZEQOk1qw8fJXuKf/MD6OFV/6Qs9gC/G/JzPg1iaKP6npfIip1VYYBQagj
kYBA6M62vYlD3hVcBpHxyRQadAsxgQ5YylHK2GVAQRzHomY5ZfZo8BAQr/YVgggg
dqGXj36sCnVe6pT5EnZoRJhGKVfSnq8H+yw8mT27V4//AcH/Jb6IombgntToLcta
hP4e0D/rGpVUS3GyiBT51R3w+eWqs8ddEDHqmzX2Xt3lfsqAM7aTjA8lhbmtHYeg
AKiTEbmAs54f8rCJCKqEYvjl/l7KES4W0f/IUK76YUMD6aLMc/ThbMDShuwGzk7N
ja38R+sK2BIzVbg3v0w2qivka+54Ub0g4HP5D739Yevy+25izozAcQlOwIRiusMk
o9hU4TvZXMM57xKuh3pnC9oFq+6IUr/4tlUHahIDKGpV8FiAR+nZgpLQBnGSgn2c
4t2YMocT0HarRcn4I+GGg8Tu10hVQ0GRZ1ay0cJgKuzPKJaMZfy+MQR5fPVrzzBN
IGLqexTI9HqqvHJXQ5Uq3xvCYnK5NJO5D006bZ91pzMLp34q/1CHT0DZK9n5qyV4
hOv415oLZBQ0OIxdvqQclSU2jfRKuRsJPgsR0yIKXYFHXxF/yjUv/3Jqr1scPl5N
BdjVxYarfHsP4BzFHjh57hp/LA7MHacWQQzZkKBwxnsmRWUk7L0CbtnHNy3U/a0g
w7V3OLzsK0jGPz1SkVclFRAb++ZGpxgYNAtlk5c0aXFPACyylO1DpQT7JjP+jDv/
n/3KKPvqtDSc31TTqHVxRBCNqxLgLLg0yp5PQQ6bVHq3MoZQQNw5k00TYEUhLI/R
JZ3jpROpvdXTltOxYbvXMEW8AoJgqQSZXJJaiapdc0ocPDj10grTUV4ToHQdKvlp
3LqGGGEpQZK3ea4BRAFGGlCfh36wlTueqNt4nvvR0f4uRsz+bHD9KKnzR8fODwSZ
TyyVWNq8FimbDM/SyksRMi7an3PZSLvTEZvfbGcSkCoC+lGH99WxvNfiorZ8I4Is
nJJjunxAnBmF06PT3WY5g/SBvBhevqrbi1PNHRaN6WCuC0PjjDBa9sljj9OBN7QB
d5MrtfoJ6rpE5Bvy0NTQfczKwWKiwXrtIv84Rg7r1/rGnL/a3uz+MuN6yZRSUJcl
RK4WHmxFNjUXScEgiEbf+UP3fzETWRbWUIMIDnnE+QL2kca3+9gpNF+cfbCkQBj7
UQqp4/L2/k7GBBmNCPmN+Bnx0aeQCzUPVriTZARRbt7j3sHK+LeyF1LjD/Q/Zn6N
LgBpRsZo8QRhBb/PX9/k/f2aA9TZZiFN8oi8gynsxLuTKzokgTApTZprsHhr3IcR
1ggGp2G50WOOTQAKIx85tupFQqjbFAwSrA2vAfnb7mmFTy8Qhopfptb6qevG3RoO
1CCrO1zkGIqhd7OzvtHmftnF/JaYyEVv+8my3vMd9wy5Vj9HaknEPo1wmJApkpCu
ULoHKNE6VyZp3nyQAmegdxTBMpb+TvYxRU48zPF0xFnXyF2QSVzcoJeLuzeGT2Mc
mlRbRCrHO092AV2hUsqy67TparbXUIA1vyP2/xVc4J693F4t5eSI7ShP/S3UzNKo
VYI6cXKg6Ub4gCuxbwWr8+cfrwT5iTqYswmK/uedak+s5B3ErcKf/kkqzCUUznuL
Abc3c1XbpeIZkol3m5T6LqZY7mZZKEutrnNtNHIrDM9LInyKelwKOgU235Ln8WWM
WvM6WENuoD6Lty7udJx2SLZiv4wjlOCiXZl6fLC6PdoRqkExAJ+1q0UwMOdQN+em
+hYU0NpUYuT2Y2oNNrzsq3wYXf3SYgesddMkWojbdyV24zeyUW0AfD4b5JAu1Uli
Z8WuHbxyHIvb/UN6U3UNnf8cRF+oNGU3KtNJWoE8KuFB+5dhe9S2PIW7sDqoMhI9
ZU5cU/C3jO7BhIDZXl3iGc8n4VIrF0cUDKkTr/qiMBimYYaLwSMqz4DJrgTu0qaS
Uh7uoXXLlxp03UH4jAmCYp3bt6c2PctSNjFqdiA3XMGJntgm9bZtQDd0MFBmuDWH
vtwfYJwfuk2JlBcuTWYnKfNvuM9MpjoW50tTyAxHXbtyAv6zUKDkfGU4+/2y0hiK
JzBOqiyd70OhfFcDuMwUP4W67z3tEc2WHJaXeKm4xXjVUYXZSpGBtmp2rV4zaByE
YdJrTKmGSyRzC5uLXu8B02DOhqxlDshYXz+c/KXBiIyWsbS6KbAZ4jxic4GTp5vw
ZB+1n4BKVTFB7zESP/ltCY5bXy4WJRKtjaHygNqIMV7bfeDCQtminvm2Bw6q3lbO
0svwv9a/LwJ2NhOGJ6svt3GMMMptTA1SCP9hosSP5VVESywpt2R9w/km4ztiAzjK
vEz2vfuCOnudaXLWp8ehJuMjF1DBuzRQ2cwDdvR07BOQhRsic71vO/gEzlu+lXJN
dhEaXx/rl8cE2miMoXscIAQ+g7k5T2cRIaT+I/W4IcUEO4jIlpwmnximierumjgT
Ry+9sBe74QXd8gylYVubzjSOaUdcAqwWYB4HnGK4AZzmNjQscfLFxdaim50AgE5G
prINQVFcJVJ+gfZ5YCm5JCyBV/CVQu80Mv0Yzx9RQp4NkZl7tu0SSSN3LQAKv8Oj
UnTrIxffKWdUlMwwkUn4JvjyzV7m9wm1gnD4NhAvCIgBD22oENeJqSMGR1RKH1CC
EI+sZB5fSd/1oaexSzue+JqPh/L6Il7ZRqdqAb0344q8XqkrerQ6E2w9DhEOp80V
DjC4xQE+MVCK4NqODDuY5W079DxMfX0yjxb29Q1CwKlw5d+jeD2BXk8d6Vl4eiZT
m1kaNLjUEsR5zqYu1I3WSOfynAiTV9x+KRcSQWpnJVsNqY8doA+QtTezW98JbBAV
oozYGhbKYsbtqTb+MiBzMuXmloyAZhEY6HY/UPGz19SMf07w9jY45GKzreuCiY7N
0dzDk9D2ImnJXcKPKHEGmwfAFC4LEdKamSgpED/hInKjAW9DUzhzWeYvpqH1zmk3
rI67C/+POupMjs6JUfjEgdZjyACzv90Nfi/VWbBfOLaLmEKQnLavMJ6RgMAMRElK
MCHPN0JCnBdpfP8c1na265rCaFsRBF6XFvt0eMhShXGDK/GhjsrHn2lIYQ4bGPru
1XjKZa1NXqUqv6rwYegsz424G7i5/ftJ+90mGqeHZ1EuWFDFtfLufEM1eN2nRCG8
Q0l89fZsCHmsmgfYbS93gAfxCKNt05a4IZYudAr9nHEsWuCF4ME+dI5Y4CSCfpiG
kbIWDuiXnTpMfd3aa3D0wFj76bfVEDq0qevXAL+xn4A7bC6KLFSZc9QPi70fkLvJ
dOsmFYglOyyIcHhYLcDA+jVSPZ8IaDxxYjIoidkwDU3eSttd5eoR+SW+MwVIl7Lr
BCLnSn/t8O0uXPMES0VK2htZldgd4PyzAkCMh6NMYSxy3csnuhU/ts4fOcil58e+
2tRD2w1qFuEounkVH3z6PIZzyO5P9eRFuB2HCtyzpD0yHaG4bEcqt3R46Ak4XDs/
A2HNqH2yliaJTJvbf6GPv0kXywxS2LIjXIZSj0rPfkeRTpZDE8sh714aEG9rH4YL
1J6zu0PXVMJcjVqiY7220zD5WQ1yEtOJkMoq9SCBWOEBB/bOHrwqrbxjdE8ER9bU
AyewW7LDmxh3QLipaW5wb3bGgQMy97syZ0fJhZnWVsamuJOc54l43/Gl10ZVWcdf
2rbQrSjSk7Htd2xtR/8PL1cgpC+GtEUxGqEAa5lAXEYyXqWa7qULuh+l4HwThoxP
svCaPuictO9140+lifA0cSdde35WdnLH1ORDMAiQTm8ghuzR1cPSDmaTlxu08XnC
eCH1qoSxHRPTvZPGV9bm19wppbdwVwLTPOo4HnQOwxa48nN6jPVOpk13FalunlC7
Q7D1ZRxAGtFTO1x5jh1VcANDbh6hOzCPWgnXo1BTdwcPateg4j00+mmc7u7gm0c3
Enpm91IR2xzTu/6sxUhw9WypAJYpim6tISS8vBJ96jGC7Ieup72g+hgjnohizfKp
FIhFG5aAIGpQFQcQdkGo9crZycrbnP3IJbyjpKGntMXVoRyNVAgGBnfLvyNNpXXM
lvmlvmqX7PVxsbIMPB2yCRn00BwOYr4ZrI1APEvC1GtacaUNXFMANgmJFy5F4484
nhiHVXJ+K9eKuPR/mS95gkC6zAV1Q6z6xM6C9hllGOz0LPYNVhl9LaNdw40bavFR
aA5m16JH1bVLOCDheKVwr/cs/gXCXEJuU614UdSc47T3NEQYEC7THbCU0ytwhe+w
3qC36ftUsd7WpseDKZXtWZmF4VdPyHaC7W2XFAnh//bGBcbDkvGstIIIgb3Rhec0
KpxhoRpH7Ac6v0JF09zBjBUsYx2nFAV0DSmnZiJp5mQxn3IbSMbEb0AOYwwrSY2w
4U9B51gCSCYMGpLmDAKTuLoSMwIObj8zkWL8VahJlXuygFvuGc1sPvdXoooG47RM
vi5YZj4sgIKCXz0VtF+tzRN1EH5v1Oprbuj3c7ntCDJsw7M5mgXUglAOhuLlEbj0
euCaiWmGfXKichP71AkHcRjef0j/RIuRTZRE/Zt69DBqDSbQSuHep46a4217IH3/
cZTf0i1xDxUMhMnDWZrezkXeC2dl1hOupkJUggXofTuCVf+lAelJ9rWK2ZmQyO8j
x0AQA5xdCyvvl0QxVdfu9MUPKNXviUSSPsYNeTOXbwM2RrT3SYnzakERUaX1RKf6
488ezHxHxE2g0Y/pAsrk5ZWtRlT2/U5lEFD8evETY4nGgwMAqU1gUfrsNOhcthwg
0k5rUuU/zOxmw8vU8g9rgsV2QmWjfTj8Qs8iuBfr4WE6zinyzyaVZPw4I4pVV1G4
TPifkm/0r+gOruFOvH0LB5WkLxMncJMMrF3mwgZruztYz8+ZHvRHPDlkHuBnZo6v
gzEq0bjt6UtRBkN3V6VAfA==
`protect END_PROTECTED
