`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
llv85qXrmoxtuvZtBbw0zY3DGAdGO59frBZtMFuKHT7Yf3rKPcIVchbS7TuLaNMl
DqqTHnSOyvyE4/rDAtR3shxKaVc6BywrLPJ2E7yIxpSX9ycOhYzBQxkow90sCdHK
ojwUpuVtmMFTTILjjK1FxjbABfjdt3DO8lncrycKBRgxDMSqFH322LOBssN5Cw4x
niZ2sEcqUUvuk4GUrCmhvNHCbOcAgxM5FkUNdRFjBjbz3h1GuazBLPsuse3vAs0z
fHO9NIXXasB+blNzOcx4DP+5tIFJ9ej7qtriY9FuERYiLsirIDkWAgQGu3BDeVJz
NogKrYRE0MjNRuTXD8PKy11EnkzfDD1yx9aGFvCVNqrpuLMNdMtfz+3hnO3Wwtqr
yYwrUQt0n7riL2znEdQXKSE494pFwPHvoMFpHVwI1zjkPwmtOAlCo4igv5jzsmm+
MNggtYah1smn3JFdu4uCy3OyyikEVu6TvtPI9mE+PHUdNGkQ74aV1XQuYX5b/iKr
`protect END_PROTECTED
