`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rf0N+6iThSGmNa7cKkXmn6bS/Enwkpt6cbkygiN/LmhuFCxmn9o+WkvYiJYLniNQ
4Om7VUoZdA+4RfuwdV25LSs2zu/gg/8h+RY5k9BCgmz60UVR5AOEjUT2DFiUq9mS
bCHYRIg9BqkB7KNU9N/HdKO2RP4O3Vp8BJbrNwc3EYGZh/IOmrn4GXv6HFoPvsdL
ek7Of1NuYXRgkGy0TPudKUtrbsv0Qtzb4VpXhkzHYy7hBXzw66KH3KTxIXX55j7s
TXj1iZRPxdI8e+RW4xXFfc4BtwT/jGB7tdTKt8naWBuYXe5WR+eF+E6tD4RKk32F
9kGmVJTKRTYlQaurbo2YFlJK4S/HNgMLoNq/gDFzJGEG/cALCdEP+DJrQ7d3rvsu
3gy5lsffW2mo6u9PcxTd+/TidB6FkOegA49QIvtc6dUH2bcKyiOP7IJNY2fd3tqm
5IF4Yzek4S7P1ikxOl4fYoLmcBGSo80luuO7X61LXvg=
`protect END_PROTECTED
