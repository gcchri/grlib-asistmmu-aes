`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WxZ8WsljX5MNAdGiEVlqScsj9QYMzocnr2bm8ZpeOeTwNM+odKF44/rBfVdL6Psu
V1Vhlh8Jg7/eUvFVga0CAfTjxZ6FupE22IuYq+XcV81352XueavRbf7mJg+FW+8f
UU6rPiRFKa1MyKgWRseEoFOKCaQizKDXyJMY9U2Yu11wj17bcZl8D0atbFHZNFOq
c4dvTDHA1ZuVrKRoHK+7pc/vJUHtd5w0hBfDQp66KXb6h32CCTx1UbxGJcb2eTYW
0EvQEC6ppkDjRMwcJMAKkQ==
`protect END_PROTECTED
