`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JJTUJMYBVrMuPDHq6q3G/Gwrf1wjZzYPNIetzwoMocXEsHe4GdWeWRTFIJ8IIuu4
x5Pzgo1rozi9WWLl2jJNcMxpBjRtQmN0GQwADlLu2tWFLp2H2zTHhTfFmRusj2+Z
INLA/5w5w+6fiNZrLVWmHfnReF0W4vhYxi0CJcnNIp8jQpEFy93ycSa/yAiZrYRG
e6/Sw1Jrm+TBBrF1K8uCs2jbVU4fAn0At3d4B0pH7lELHGQOW7xl7sssM5H76EkF
YZmqfNTWnITpBTNuF/oNdpkf7vFk4MLNvFIsv8hHqShfvMP88Imd2zQLy8blh3+l
G2lDG7CrEPLuJ0f7Y8Z4bUZaPM0lsi5qsBkd4iTlIFB8NDB89ZkZ1wtcwuX7PHTu
7wC8CS1jQdAWfLCoIbBaB6NA6q7xrLl88Vr3ofYc5LkTQyUD2WK0NfCYXg97NBRE
ct6U4REE9ru8AtTXe7K22RGTbTlOrpy7TIyqJ/m4lMqDJiq/jW9dWHGtO8Y0QOen
L3z8QvE7nv6eB96oOeWt4HgL1r5QV3JNl6FaIcE5OhIYe6YJuKV0Eb2jakFTULxb
hGrK3iBdSHuoB4ZJ8hDwFS0ChSp7VGnmjiNq9zJ5IxLHFmNYXe/51r3sfb/+HbFr
3sAxQsylcwBegaiZB7Ji0F+mtgF+TxVZE+VjIUZg+zY601xCp8NV6NkyOT789WbO
QU+p4qAOO/INwfST3jpziExkvqN+N02gDukkOkm7/LyzbayNjQbnLUp8u1IEh97J
aZEyM1x6g2kk4EvMH2mJWMAMVY+dhd1nyN7q1Ufrgiqr/pqq5k86f+Oezin8CK/W
DoocxPLLRUsFrtDhOwZXATNgTl/GDav1t/yGliCT8pPT3T22o/ndk3dVxXL7buEU
rWbt1asESmlZ6fChJaxKyRGkTqQ8qGeZlvU9AznlylorkWP56ioGu+WptW22I5O6
A1g8yxLy0a1g0yrRmNy6ordiaTVnNfRkJGyVbPj9kQBg0HQfY8T/9pjW/3n3xjz1
WQcnBcoK6mFqljh4kvkgawS4UDlEU55P9vmPj4c2ny4r7WoLfzvFva7bTnWSIT22
G3SeSeqw5LHbx3plq0CbQruy2LqyQqJCGFCJNjoOnZKtol9UK9UThMWn58tNBnfq
nv88eI377pEmqg0MAuzT4n9fUQxR+/4bE4ohnnj8cUDCPjTEyziGEFmqIjfOq1+0
jfMb8889jR7XAeUCzmPzNJDJeucXmlEhyhESL3e6SquzLy/CHo1CxfdtSEcX0Tqh
iTRGhgdb+pHZ9lNUhEASuZMdnAfm15koHfDw+sei8T1BnhXSzm9VdJGea5Kc9gQp
uNlmnPgiZcFg3NZFCEYgpi1d6u7KYZu2UaEU43W9rOnrB05vNlkL6P5M+I9C1kHv
SrLrM9XQY7iSvi98SfS2hwG6z0W+CY+C5zz4hdmuIvqoHJk8Qt4yTzP7KYcQ4iBH
CzLn5kTlrUijIfWtjOcz2HnyRuKIsTsCEnLnyHx62kU53/kgy5wIjaKMzRWhMZq0
Z74cn7N2gopMs+YfS2GWHdgAkH6zM5Ubdw1yL7A8c65m/yNa738a4S/bWZwa49QD
DhmWBc3nzKrfmN0TlLISF3meZjQonb/x5Mxit2Hezh5o7azAD4XA0k0bVZUKBnxv
8QNmRUBqwNtJMMqxwBTEXciuhHhL6FNioi70DNGWC+61GBO34P+QHf1pnE8uR2WX
d19axZD1Or8SWQ4Ql/4Sf/xMlCBYNBYyL7uAMuEI/84Gxl94cw/scyWXQyJfBvEY
9Y4A1jslMfFEUYcFuX055XXZoWaAC0bmxJQpW17sdt9t7+bYiW7COHYHYN2wTKbM
dnRdgkTIZ9Z0njMCnEA9qqZBwyKEAMRBl+m8a9EsxB/22w05ReOFO8Rfr6bK1/ya
IeUfUsJBG0RmDxUBA4oziUHH+Sxaq6SnogXDc+9DJmypLUd4QKcp9Dr+Uu6WaSWv
9vy4vs7ELNV7GGF9CLE9DQtusbCnQwYucxwfXcxl5uQhqFCSq9dJM9bDKHnLWa34
yywSFSh0i9tUk+5/WDOZVp3BfpvttKt9QWjhhXmBmJOXIYqSpfrXDaTVHOh1A1zn
IFYDNpicsf9RiYkjopPhH20/+qgNrWPSS4TxGnFkcKTcXpOeF+Sa5mVwAqcADdpJ
0V5JADgmGmTZHa7hojORrVkyS/K2GLzjv/gRdRhw0tufEz9vhFzIecmum0Kk9xs0
DZKJVdrifC+ryBvVIz0DnYHnobQW7QcDgnsrxZXK1i7lqaASD6Jv0vwGwGquYGR3
clcWzd2+NNU1xFIQt+NmA6rsSdjZgW2+LGixVhzvYBAXw5av78VGK5o8gWW5XKwy
//3+oVivoKew6nUS5g/mrCdvGKOstHmTtPQds904mN9En1w2f4AAdq0rAbjQRm/+
flUPN0L76l3fGGrkof0YBWG2DUm6pE9cRI7Q6XUfW97GXyA5kufejf96Qu7kfdBO
Ek2OCjYbrDq+ssCysFi6tAp+i9/YxX7iIncqHvB9H8mMlZ8R/2KvYkPsj7nay3DB
IfGeGeW6xMIcjcqPXiTJonNNDl3W4HrZa+MmwACQbK/y6NG+Sx+gZdwtbfmzfXPa
8WosrqQbZbxvj2S2ZutLXwtjjOSG/2mOS24PVbZc8ZK5OsWWJnQLMEor/JesTAh6
3QbuFinRqZNIEgqurFu+f0sc1VFs3I/aHEbAGYi4rEpC4ra92P5BU1E6ZOWhx0Xh
NIDascR7zGatrr3XPDOJUWfsPOefK2BaObjx1086Z7QrQQdgv1MfTo4FDemF1es9
xezEueJbI8aIMNdm/KqFL6cjmWQ/FjPZlPauPfzNtTmh8gzZT00k4xwedPKZcGFi
KnvFzqtY6x7rc/RDshw8Ky4af8k2XrccwVnkInjcZJ4bvnD1fAbay6Vr59pDBS/c
B+he27DlzV6LcYSbvtm9Tx+G91/52WJtSQV+c1OZwR1S5N3KqXGxccNjwSvSmPM9
Z9R8kNh0xDlZndI4tJmBlqrEJuOqHLb54IOGDyRn4TbCbLDAKg3YZh+2hyiWszc1
4+tZRPmprjIMltqOuB8KHZ4JFWQBTTLsUvV1wrMTY3TZsiJ1lAcAZSrMN3VtplBA
we+YBOE2e61KW9S0w6KmIaKIWQKOnl405bxwvasHfYJMghoeDtdmjC2lJeXuDR1/
faf04uRQL/keu4jfS062re7EvWcpCvir62N6Vo/r4V4OLZl/4xrDsW48ekCgCyfZ
jjnL26omVYAuFiOjXBZ+ncN/iA+JNVM3QudO976FmM3YZpwD4aVcwY9hSIChdh6f
WmEDOTREVMzVuwUIuhBKoK7yFiHlSxKag0Vb7c+zkSHJpDdspHfkcUp1Saq5tJHr
C2tTJcO9SyY9O1RLjCiJsr4dxMwDkk2+ltWouZmAuQVQplk+deBEgqcTUheiCspz
gEzAj1PrrXVGKH1LMzdN3IHP2xwULlYiPMYNoEua5AhY7iaagMVdbaS4UCpmZvbR
ykgt9sMcPdFVZjHoc4rTjhg8ZEBUpt2wdSDiaqqO5hos4kItlxgw/lqK7WvSg55N
NhbtDbXTm16jxf3Cg75EwQzRd48OYRkcO0V5P+hColxvnlXu3eXDktuuUzKsW0Md
45BmLePjPs404hKTwb391JNHoSfevjx2wgQlUoAoYut226PjIciKD8k4daf0G2DJ
DBRfrHbkfCJLDmgwoDgVyt3H+hYNWn8mgv/e26hSQ76CFul1/LTiPlctEmxm9cK+
5jaYx8seldo7OvNqSt47zD/iucRNSnYLP6/Vlkig5qXM2NVAfdi0bUSVijbk1UdN
CUai31DXvU21d3WR4Q8ILSwgfAwYOt0Yw0HVDI21WFxSl+z8w3B6ebNPaEO02zLT
swsDjIQqzqHqHUTuP3vdIu0UXUVg6YcouZy1Rly63IAv4aKhloGE8gKkysmnjmuQ
2YL7QpUb9Sl5e3O+62n980fII/0XKvamIiepuNxRVDaVxLj7/KRCw4YPl48RYZdb
R3ohqLMUWbq9Ao7nQn7dlDrDIxPLqOnTH8TmsUf2zdkG2ACgRd8cpB0u0tHtIJdb
kErQCmZp7iGRzIwIDgykAk/sU9ENK4fvw7KsPkdPK6yxjsGkFZmFb4eHM6Y/eF3l
uK3urp3H915ZTDohoYsOU3IMs8V4/jgug1mXatb0ZH7rqsEHhy4XrMNTFPkUHrge
blSvkRNCFchGYRXkrSNg3ps6Op73KvCOMTIPomR00rjuiS/UrgCYQluo2F/dkymF
3aGkW/sMrXLVwOeyOSOwCdQToYT447q3p/ZhXppviNYJsPq0eDrwxrRK8CW4gPyP
TrOvJ5RQpvL92DBtNb/aiZBI3x+WQGgCqcHz/Q8TDtbpC0tNenTlU4hCXzkohPUz
zo/QzAQuLiOhQiJbare41kUTygAkcA1ek2GZpjIekNvjbg9A6fZy3XQlwaR5xY1u
q0QHGG/VJ8alFol80J5YyWpPRN/6w7KZM9XckGOL9mwen45Q6Kk8vp5AQTsIAVkQ
Ym/Qado4YSamIENGQ6Y4O6mrEWbJ3Pt4TSlxCjeJu5U1h1LzBdw/if7ei6R6dK3H
bcrFMdT49JUpSXATdWpxjBGeUxD9ClbBUalHeg8OszpRyNoYmdr7Q73h525y9JkO
GGeD87kuv3WQwhgHHcS0VZp628sNkihLKDNRVpOVxDpxLMdDs/dYklD1Mv3sJ8yu
L70iKVR7wUAVeBpmUHlxCM1IQy+ij/TV6BsGjbKvA62pyPKWXfaOjFacA7oYkGcm
ohxJNLJvY7dsATAaAKARkWN57c4IDvUnRxxJcR721fd/heO4mfZXpZuAXRhUjS+e
0Sd5I6Mp1k7mXIAjpfgP32G6ZAjJwFcGgBiqvI369D7Yp3JkUhgQ89rEyv0SDv8b
sU6RjRq2pEQe46yApEFB/okltSfGygX7NjSUIbutUR2POAmvWSrX+SFxa4AOdRkY
JNhxBxJ4uELnrqiBYI02IkxE9wOK/4GTygAskm71nDUS79X30NlqrVKLfkmkydw1
OTCKm0SmdNnp/BeQ3/vW3atoLNMozZRBMLROFROOkR5sbVq6DRRvajWTGHJ5Gven
qwoBz9hTT58qY9AqR205ymOrcORbrGFAgoFhHkpHs7Spt24eYj28kDrP94BnImIG
a5vDkQUaVG0bFc3GzLW9zl4sCubo4scU9lMUsuAeTAhO2tRoprzYm2ShUcBdwK1v
dSTD/fF1mLlSiKTq7D7PU8JrqVBtZpMJM0W2Av23sqU2I0zDcn8Rm/QxMR8KTWxy
K5WHX41DrDS8OmF/MSYE6dpi/wN4pbXiFLE9BYC0S+KUXFXg71zexgwib1k2G+th
INIxechICMpXOWF60Ctjt0gB1+YQY/eUwq/wG829I+WReVz0Jg2WjBUkKKVQaJRg
SxaBeHOw8HYXgAATqgiCmyheJSHAzjO2bMwceKUrD43X2YdJiS6bLa40qBMp5Cqt
2Qj1ZLI9MtIRYbpA1xX3mG+b9AbKXjvFwNfbE6cJ5wzPD7neNO3Tdsg75pCFbZ7b
X2BGbL7oDOhnaSH+x/nhXWTggpy2hHUReeKEULqqbOzhFIdsgpBQHiTPfHT+TJuY
Wfbs0BVOG1jbO0kXmuA4bXqLozjbk7Q/rmjVCBlH5ucOG2oiFSr692Y/19ro0WD6
8rmBOxHnODw0y0aBC8dTPlqeHT1gGnC9wa50hxdii/GAblSi+RorYKy00ChO3a6+
q3+POMWw+XgvlM/VfY4IukClisYY/cc9hvJ+0kpomYavTf4+4h9YlZzK/AJPcN7Z
W45KSEkdGKpnBnIfSg3zhw1FW/ibWJ6sFfFklNx/Kv/KBu7uDaV6MtcEc+6/a56i
NyMYY0fuxRejeFEezwqyvRACv+Bx7W5vuhvC8myP5a6REj4xL3ah5TCAaG/MK/+y
7DjYt9SLK1kIi41CC5HpsR02x+iRJftujB9g2T5o6aVL96pj7alf395ap31sXK9X
a0YLe3BQWQu/54+q3ECBp3Si+lrvqpvKCUZmsSHeJS9QNUsiDD8FV+MZr3H72qP5
usoNZmS9F99RynmnUvUyk7c4dMcf4gIjw1vUYmNXRFyu9zJWG1wrk1H5g+LO8rVP
ewDLsGlq61ZtsNGEZItZc71PyJkwl0fx3ILn0AboB+pAfszSI3XQkUrLArUvHZXW
tmo3KdMqN9mkBBikj5G2/BMF7IyprzCp8WytpnExF7ufI7B79X2luyTJ7f0qPkDr
N79Vln2sfDIU6CIR4zblR5GjxhTFA8wj5OkaLc6viphAnNw/8H8GKXwz8Vbms90z
63YtHJtFcP2iBxVLahpiy/YMvnu/+XU9wrckL3jx1agt/SCo0ezMePX1UOq2Fl4V
xb29lDe8NZk59qbmArYujWtL1FO++1w0H/5RlKMe2dtvZdfwianZ9wDCl8DZ69W2
zx+VraqbLlU8zYz7EF1qHoRxrr9CIqEkrgOy6qB2epWyCzwRvFJNdWwQSvRttp+4
gAks0+QmiafhtOYNHP7oYBVOfiKWnkvt5cVcxlNaV55vdaaDfuuiuuO0Wj9SBZZH
3kslHCHBvCyjhoziPJxRitrwbVh32dAzpw1DaOcFzOI9ehENGumTn7rDRxDtMwLg
SlAP3YuHhTFWIIEgGMZNUGcFLZsgEDK9cReLoicvEzGhs+jfxCcKrhrcNItmkiMr
4ceDofAlAFBm0bksWx8T9rzg2A3KirSBLFB3QFEncTj9acctFtUTpatOSRRSMqFT
zMM08QoxgHnVL9Eg3PfMcVIKnjLzn8yMYDUAFfVc2kILiRh0qdqmcMnfxoQ9DRTf
qx9REYnsDmv7Q/NHZ1SEw74vqZhR5Q05YgYqQcYzy4oltQEJP56dtsc8pW4LSTwd
Z1oPXFhg1xiB0L9YYCKuYXvPBptV/CxvMhyxhnj1x8E=
`protect END_PROTECTED
