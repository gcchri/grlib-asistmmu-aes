`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P/q2sNh+RBVmUg5aXIDcdbhjF+IT9So2b92wYJLJ2+WLzd7h4hGeepGTlllwyhpN
Roq23oPCxOiypk+VI7SE/+hZfOexM5EhUEOUb37fd7Z4wSiX6F6E8NMzJFURgtsR
90DtIbcxbDqizFYkpGJ5dPqKxjUD9MgK/RSeC0TqYf025fkMGL7ESHDF2TjJ0XOO
nysp1MtGTOgp5/FiZ34/jJa78M5Bom0Gte1aarC1DVcR77nBL0qfcjYT82TuQ48o
X1meoV+mQ3hXaW2REu9SrCeMSLxMzdNKEokkNFbjzN/J8BeMX/Z2R77Y6oibC+t5
bSRraQ877T7dg9eepAum1rTktPfFdl/FzYJp2dntgKfZtXZGttxli/gKxS67eYDa
Lg+LxsRhs0URzQMMaCrOKhoHieE7aySEJEwPfsBXpD1oHBhFrh4gpCXvSJVC6i3D
mrwgwoeooAa/P9KYmmmCRIsA1ollnUCM1fLCKGB6qQEZTbYVq3GMgJRXbTlFz9+V
EEX0JgWKWxBegekuCOZu/sjwR2KFwl/5fuVDGBFGhOCO71eZKSjhNm9F9/AE74r+
u4zUELkrZ1DjLuXrKfb/AmbBboyQe9lnuvmUn2mgE8HgoORj8ZCOlvTD0HOMBCZ8
fyqU+yt5OgngVxvMWf7KyvuWZqgnJrSvPJSXGaRLHBQZcVwFdd1sOgf1/HWv3uan
ZhnGxND5pw7B94qpj6icR38tFN62/xPgQ12/npAmFQqfJ9aVnP6i9kJ84wcXr+1P
SR2mJdMl850I/47Mt0OjvgUWatQJgiQtixTgPMQzCxlHfUDWiLYqLrHyqjR0XN7/
9I42qwEG9NZ7eMFB04ap0S6bSJr+2tR0eiulVM3VrJoJdUHpFSi+C0e1GWAR3Ip+
ePkjTsJxbFzCpys2f9uzA1b/ONfjXm+qhnOfW2sJIeAoG96OZyNqLjw+Q9mKNrKg
6zuNkwFLTDsXDkfF5bhp7IvZB7NihvEpnmi3BvSxpQg1R0Q2KvGSPkRlhvhy9GtQ
`protect END_PROTECTED
