`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4rFAYjQivTpBoN4aT/vUQaK7Q4RljA9u4b4pTIuDXnwd9jaexwopEYnR5IDwhSY8
gpTRZINBDoWU7jFiFi1f9hHwd6tNOd8k/y9Vn6dFXFJCdrO1G4m7DXX8plSLHyFU
AmN8FO1Wpp1EayccTM3xpcgS3pOsoQiIMGy9t1HXXUke1LAIagAMTpJvcYNM4vHc
qlAb5r62mhfhXywxjWcWG7aZwksCVJCyuAfR3C4i/V32yQ6bS2iQiaD+mtr5oBsd
u4cqhW9ayUNfIGk8C+wUtcWlpbQHTsEsMMBzkwE9E9IJ3nz5NerlgEbLXAfke2Rc
uCzljY5EU3NlT0f/RUYg1N70neCO88pQQV0gRbCpjV5S4jFQtcBksSVQygiFavNv
lQFGtZRSwHa3N2DFHgNVVGvY1t4ppoz4yoBTEKs7bfJ1EkPlXTNHb2PnhdT6xt8S
dbODvuEb8gmxbfeOAEt4XihXMYUKntS9DGgpFY7vMwGeGf/BJvYzDc4CrCiodv7E
cbDH9d5qOWvhDWrw0P48V/OE7RkeYyMZiV/sdpe/BGHHTcZ8kw7jCMXIKaP8XXtw
KjMiaxkcqILmlxF8svGxZuZmeD2LZ4Hy0PBKYKPbt20jWbIB0zV22D+/53aTuJmJ
oa2UCs7Cq1ZUlZOPEAST/OFX378tYEYwt1/hmAMpyFI=
`protect END_PROTECTED
