`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XNGEI7dAOMhagfjLKXREefX4EBXxA+EaBfPGko/1qcx3LqacTgw8STu02ht5mLey
t/xRzzxFs7Xd7QFAJVX/vmZNavDl3tPxV31ypn2eY/fZ+NXHV6pj5ypFKpSPq/jj
0uX7sE76lTrxc2+MfZSEHbB4FKZRb5OqtkNN9iSqmE3j//db7d2NWHRsQzRlPjDj
nyk73QjTBDSFxO34J0A9WlozgIXmXT1WS4QUdZHSBS2n4F3aGqGn8JIDEmpyM3uB
G+XqaBo3qyGop7qCcLMviu3NThxVoJgH0yUwau10+Gr4C7kFYfTuBxodKXgRJ0Ii
A3EPv9ZLN7Sqs8m2dw5fHRluwevGYzBO0m1IVAPNk6Qdwo+NzrWtqFIVgfII7f6y
Un7wNvsxVV7tjzoGJ2Cr6IGQoE3zwETK11AkP4upsba3uYOftEQMH0Fm9gzubtkq
MjDJpySmyLTC51O2N4qaCKqnlg4l0uaccYP5oW6Xcu0La2B9hmY69a9Acpuz68Uk
kn1qyf5CovIyL2LS23ablER3cJmVHwHxw4Pw2G//qP948PnkRrcAalkwEW+YTQgJ
MHaIe/Chc+KwnZ/Dcx9BYQtaZwblRAodumlmgdAHxN0=
`protect END_PROTECTED
