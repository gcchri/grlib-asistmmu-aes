`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IjBTzQogigJsM90YO1afMb3OJ1Bq6I4OZzcEpvB++nRspMnl7AjdHt7uczv8v7jK
gAM2CdFIWDo2Rs4tVTVkxLIVUA8ALj3Gjy5KgoYpkig7UdVzx1uLsx3kBw+UC/Xi
fLw2slqJLBvdX4Jv+Y5YuubGlmF/8+VrwRU3TRO9DzkmMyK1vEsOFBmpyeiIf8Gj
txPknPvnOvWPT50yNFizay43T5tfkPsZrvyFfZQvImzFTuV8GW88gAKgV9EgPHJx
5v18zWLF5xG40cJNbHxxI5X2eWkrY0PphqmXrZGTS8Q6KVp3AUO2VVsJtMk7DBQK
CF0DR9efanFA6LQcpUQmQTLjD/O/mkRYNFe2mAhV8SxnhMFBVkgm2aDE/M7p+OUM
C6ZP84VCXg8T2msTDfKihSKHF+U30E6BEnRh+VzIp3KZflqqDRVwRzam4TUX38hP
JcJSReu7/a55tDgqtc+fyWGdGTb9I0CeTcXFFltlv6eF3iRZUNEeYWBlBJ1/bBEM
MGdcsGk9a/Nb10h5Jfp5tzCtsOuhiHgfgtFh93X77qEe05XOABPK2Q1+w8ZjFj+2
R1zswm5DAn2OlfQekzWsKRp28sAQMX87ql+nUG/gjPWqCJa4zpZFgW/sBwwHJ9yw
7HRZzF6DzwV3diLKJKkMMwVE4hqV7pwzCKJpkVO+I0dlfjC5FbJR/9v54430vmjU
+KK8ltvOG/GHAHWEjxaBKfxi7eX+/TOBijcpJSGQ2/5c6j721x4NNSFdGsGyXcZr
RmPrkGn+vJB2oyAYsUFVs4bOAERJ3KbXw+HvB5CmrPrkX5/Mqyu8SgtVNKidY27s
ABigWdj99sz2kmdT+tpYJhtf1Nh2bbu3sfeFMvJQefVZuu/iFg7vQfSHI4pvM0kZ
mXQs0s9avtUTw0vM9z1YOdXovejGgqpPih8NyOU6IerVd9V2LJ2FpAvoUb052yul
xor3OrszQbUxbEfoKZaxf2qbmRxDcJkptF8rtuywiEbhtlysjdKcNNDHqlQUOAIc
/VVKjr5DncZL2hC5uKHhRtw1oXSxCDsBp1Ts08Hrmz4zMZLwXffF1BoI6FdwH1OW
+0oNOjRRVxH0GFtYSWjBTm+qa4/Fm18vfl4CiPu5Dsu3o8hfZco090QuGbATAvpb
Dc4KI4HNh9wwig4YbBLdBA==
`protect END_PROTECTED
