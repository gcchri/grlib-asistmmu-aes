`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CvBf920cO7cNDfbaFHDIz/Kup0IoQK75ysAR8+7BcLBKBcvEnyZE4k4YA8HKMxme
NGtoG8aCZ9KyE9ZQyzdITpKzrZsWinQF79WnLFhamacoztiWqNg+20xfa6sAsQ/q
42kluDxl04a07m1C8tG0xGYjxwGB3SGF+LmXqBfuTlLZSLPLfiL7T2q9NbaQRPgj
uoDuDD306jDr+5vIkSTICxLfSRnd3ep5+VXIc8Smxe0TWlsWCW0gdbp2uPUh7NR2
Tc3WEQ/5BlCM7mkxkHiAsNbK/HzRcEmV5IRDxzSwQrs=
`protect END_PROTECTED
