`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i3rBbU6oz+PuwNA+dkworR99CSMnxYYnHlk5MxrFQQY49FZRudvdH1azsYuopaP4
IK+1k5/K178+hzOsQGeUBQUP39BAI3RiRpSYFycgDUJ7rjFAyPTr4Ls6yxY6l8P7
W8QSS/jgoswjt9R+E6CqhRaVL3apgH5n95OKp2ORy1v511CE/WHmMQelHMcTvkQh
I1/qEgKCC+8dBreC2mSCr+PvTS1bAi53Ddsj5wgcDPGIlujsCrow872ZvdPE6IAm
bVt6rGdfOlNjvyiFnWvtrNTmqSHOJj86pxfLk/GvR4xG8dL/LVQv00l+luNiR49o
Me6H3rcWL4hyH7btC1ANX+Qu1AvqpqPcQJzGSeAeHO+t/jZQaZ3RIfpmHrUDeyd0
lQop987T3O3a9Ai6A1Hjvw==
`protect END_PROTECTED
