`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gQC8061rGZss74rCYqcO8/TDECX/KuzcedLuu11LGU8AFzfz51IoYY7JtotcYLM6
bKp8xUM3ybfDjAwN35XofUBnS7F4yW0vvoIw8aa1ritVz1sX/8WtXzoYIohZMiAq
jwMH/XgoDyoRtxFxhzmzC0TDbAJwizEA/X3ck39cpprF2r7PK6eu+659vZ6nafCF
K6CE2rmXlP268Zb6H0ryLH1w5I3IIoSb/JxEtWg9JPaicdTHIdVUBFiP73uhfZEd
dFDRMie78LM8B+gaB8OfHMWc7ffuNZ2P3GjD2gmiyUhb+5q1d++dvF4vI0yB4cYn
kx9erktJOD9BrHunCr676Hl3+XENoFoA/Nj3Z0umOL/1An9Fcy0g49v7jcnLpZMn
D5AYzr+vI0KgX9Bruh7z3JkpULhMmV1xXBKrpmL2mM6cJB8QURDXHiB2vss6edaX
UJWWPTiwow/9tQF/GzCAPhtOJptkVEyDZ2gUqeSBXgZfNQqLichGC1tXlZnPp2Hw
xOEZEQ5zgiWvhyI05oMoU9EEUoVAwsh5cVzIMJl7/D2p87Q+lfUsohD1c6sPo70J
ZTkkSjYqQGizTFlR8L8hf3g5wx/Xfy1gBkr6P2bk5mwWnZ0xeQrAw2WD4yOYKXWb
nH6khLG0q+WjVylWlCe6BxaLLL8t1ikaD+tk225+q1G0xoho6avb4u4+BOed2Dqv
ZIyKabYBXQnh+pe9Cpv+Kb5arDPyhzHrFtRGtbONXdRMlt7SeYCXmQ1iVynLiQOz
1taWuyKBZ+0MfRSjE2ZCt1LD2uDvGKLPOmKnvzKUDsxwBoo+AffcfIR06cpOuiyp
86LmHb541q7FFxh05SRywN+kwo3/x6fN+Pj5TLtaNyKE8MQZDoifN1bO83vO8bo2
Krqcl8Sej4SBdDHEkfzXZ1T5iuyfC6zf7Cva5huw8r4=
`protect END_PROTECTED
