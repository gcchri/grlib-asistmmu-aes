`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/ix97yswJ5ipmVrKBFAoXkSBYpDMNLsfl9mcY2P8KXjMjBUcbUJGZRY8Ssi+vPqi
0dVtLgbqcw77BbsmSTLZX8NEW1EJ0aO1TCOvkK7ZJICLC5afmtnulbO6oP7YHEY1
PlZ44o8S8yqF6a9NuleleaGDKFaCWGuiqB90s7RSTsszxjcZ2pb03F1UsSQ+l0Uc
Pkk4MANYF72SAbuWxul8AL4NPw/wjid6Ll4wUfKUqKu1GALUFgkg3A6o58cp1RPu
4rvFz78IVao6NM9VSJxqbI4bKBhp8C4YYO+dYhP7tlHytd7KoB3WHxbIaG1ef4n+
TGjSi37qm0IEbkZcuF2Wsb828+lcmcI57X75amm1lWCoItHOFs4TZeIcqcFI3nJx
Ygn5uuCXkLPXD2nDMea6O9gqfi24/ZBmz3tPkwSur0RqGe7o1xTQMEMqCtFMIv8J
8USM5v/avPaAEMfl4pLhU9K/tjhBeBXXERwRpeMNhhR4ipl+gTp41bkeKobgPRav
9AzaIdZNdbhdQ91+em0VMncglVjE+mSsRid5ryBOByxf7T5RNykL1NS4yS4dhaFq
vTylt0xfPPmgAdswSsJBnfCjFZazq18FsslhfR5/zaUlC9kAyPvBSWf5UsX017vP
WKXVLLflq1MPKcH02JzaRzfD5kBKo+s8e0/Vum78W/V9irLA3bR2zjVjdIuILM7W
f0o3Q3vTz6SCu457TXtSZ/Ip25xJ5D8YtXNSYU9pe45VAK9PzpuDkea0O1Quze9I
qhoQoU/z8nbQFOoYxcHgJB1sAN+0BnQYpOhyeJe5blrM4hKb7oJ07znTwrH4OJXa
kq35pf1e96xkjBp1hS9NIGleL8HkK+/rQU1k3QFGbzRdgGs8FXNQ/9Vl3clMPCRG
cNSGsmOlaGe8lz/jG/S6GB2yIOjaXIHTqer8ZSxPtyiOgi4/cBQ+SRoU5s5Dg1vl
`protect END_PROTECTED
