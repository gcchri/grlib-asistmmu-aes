`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KBmXnR2bMGkHmDKhpwVg3j6DHHykuezfMK6SLzdnaA1K9Qh8eQ9rCtwiU7nCxEH2
pmJnqWMT1GR5JzGFZEHLZkybYDLpbxSX/NZxjnImsxARGk7c00Pn7ZNwhQhcyBPp
SI7cYO+P5yd8gEMxZN71MoPOhRa2XRckfCssBOjEI8ETztGodvjiL2JJF8I4LSEW
hDDLy1DNiZ1NlLRYBG1WcsyXrBcSxzRVwxImWj/mM+VYC36GxVqMyQFQ2N1Fk/LK
UlnXjY7cy/aWnN9VcrOQ7dgZirX51HYZOvD+XRPK+nEL7jFWZ7nW44HF7TYxlr7C
ULocfscnydrnCzgL6SU9fddxD9NdFAYnEHQHHoxe7opR/c8PNF3ho7LrR82Hv8NQ
TPmGcM1i/dFg84U9sibINSaa0sWiciUtg4U37ejQjlww1cpRRkRcXHoOBKCBHROG
`protect END_PROTECTED
