`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YNH2nRoX6pMqWHO1oYo3HHqyGFUsw8bshzWsmXzorqgE9ypSQDbIJMAGnfsJRFmi
lMytRWTVOpaS+d8kttsQJsb1Y+O4WbbW4MFQ3VDI1TJulsHPjBxiVy06JXuCuTBY
FTdKJpeM2Sla+8oBB1k+6tr95o/qJOikpGJYUyJwzL7Wwx407e4Q1gx2H1drm8pk
9ZBYYgGX6MWubM5r1LFd3ZE59hl4J8vDl3i6dIRkOEjbGdxXACCEmCHLzKFGnCet
ASAS2rjRs+Hvke9zCq1PU6/A8veJKg/+PHm08numqZAekWMNXbJ0yiDbdL+VgtpA
`protect END_PROTECTED
