`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rmt4TyUSVyaY6pzWzuN/eG3bpAUgQ62YcY/+VKauSwkPox41j5FufnzDsFFiYQcq
aTP2tcEnefXVoNDr90lD5PnqNh3lvAiJapLW94YzEk0K3sCN049nl/HXilTS7U+N
q+4C3MbX+fcDhxZBcPBAR0H2UQtV8FmcwAXNbJf7TmiATQQ/khqRPfIq7CoV2UXN
cp6455/2SBeOJiuDGxRxiv8bMnuCJyPJwpXSsXdSrnM2hTXxzLtfDBVZYDQi7zB6
ugYkaPpjhTmqOcNE/QZcelb3q32Hm5MJ7/I3GXCui8WOGD0LFPBTHiS0xRZLWHs4
mZltQLM0JQwHAOO39ms83bf6slkFmMQhzR78p6DPxpqCDhlkzsPMX94ZfSU/TVHs
`protect END_PROTECTED
