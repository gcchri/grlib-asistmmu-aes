`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vpbVZpXTU0A6I6348sUD+vd/SYEyvNncC0pNf3UDL5/bFasaFYuhhkqyp+hZX5o8
MpJ+u43MLGi0Hkh/E823LI32+YkTG5lI5tcVgsd7bKjsT/HlHcHs7BFWCTws8cio
xKOtpEBbrTjxU3ZawvzPBecH4Op2WRV6ffeNhx8RJ/6Vb7gNWjs4nVtiV24M+PR2
FVLHHrujGw1j3ElhpoFwzMvA9OWAFrq141Yi6uUQHnJN/OZtisI5CmuzA6ZrG5vm
I3S9CMmVIa8BXGSCXzV2WeysMXzHQkpU2CvnTfEV5IONRCqQU5RZQPeArNRzyT6H
cQH0fGdta+a9PNR9H24EWv7Xa2/p8nO8+YeW3A5aRBJvW7jddQaj+OiT9Opoc0Iq
m1itJ2kHX/fLP4QMkY/8GuxNLzaxr9hxkY5Ynz8c3qJzrpkTWNSU34T9FnQG18WT
6BsKBI/f6axC/MSoXHS1oh1zVSzMO1l6sWYFdCipelZmabqyl0Vn+GC+R1i9JPIx
8G58e3RVzRDIrYiMQQHxiTOknoJCglz2AvNh7gRo3C1+qqajwlPWAigojrWFZDyv
`protect END_PROTECTED
