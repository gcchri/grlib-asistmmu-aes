`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eMnML9QCtP2tiYUUhCz5yHFmbzqSovNbcwzT9biZDiiL2YOKWaDsnz4obsOFFx1s
chmIgWJYEYQscY8LH4DHQrDUZ2sXy6pYzpwgotCORQukBoDeqIzw9xhFqrETfMIp
Z9N2BGY9mieNuHPOWDegROFhqFpHAVxKKX789HAaLpqVE/K7l/0FRKT3SE84nwP/
TKdQNd26oNdj5jA+s9VzBgHr8HblM3M875g7dPNJ1PUMp8rCW9yxJblTI7VDIpJE
H7svH/dcSqcRApWfFRuMfga4UUXBfJrpQSUkZ57CCeW3OPFdiEP+OuTj51SWRe+V
GDY+hbdVsvvj4XCtlY07bnRZYLZGNRRLdhg8exNHeMnjTDVO2m1OUOKUgmtO00H3
6b1WXGqEby6CHgHaGtqde/T2KrQDtvNoEt5xoyGsVVySD9gVQnZLsjftQ99Jm/Dt
cJcD1Uv5Adn2JY6XwgTp6yJyqEQv/TM0anXiNbFes3DbWZ8Hic7Y8eaegCjlB4GS
2fsh0vTK3iF7ChRy5TNog5DY+KD95bY0C+zJEFuNXrSW47ijsrKEjqOO8smxy7vX
2W5C1BBkJthtQPwTgzlmZA==
`protect END_PROTECTED
