`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R76qIc66Ni+P+jWDcvi410vvKhNSYdtlmflCmrYfr+5t170efWEp618J/TgkdPBB
we4EaXfvmN1J3Nbebz3IGeX5m1MpsASXaaUSzXl+G9+MPTI3eoWUJEgBOYSGiWhr
S45wthWRynVu0j/anbJZrNsC8jHCiVbe+AVloe8ovwlO6F+9ijtcoE+A0znwRqaJ
QKDl3GNdJ+rRWvgke7/OmNVtWaE/E/GgdXIRGEGM5RHhg31zg+ZjRDmV6BHluk4S
49TsC9pWL7MbtGh84uMbIsx60FyvWWlj26SLqu9NFdvOFzQMqkzLzdD35siI6QE7
bOACWC4rAZFo+J9MbTst6CjYGx5anLRGHjM2LBZl3njXLkNYcT2JPaaSQhBurxM4
1Sf3LjDakDRZFL1yWh6w8A==
`protect END_PROTECTED
