`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BPBzQw9HrSVkECs2SJy0o/ohpgoSjwDPFVGdZw2ma7XXFf8qwhk7m4Q8BHZYvE+a
aMRciOaCDUwbOSLqiz3Lqa7hzlCmZYxUUxZBfeizBSAgiJi9QKmS4qbC68PHcOwC
WEInCn8DbJkBRGb3HQP9rfG5xZmBtWNip7HL1LwhsEQ1RVE3/5v5bMeib1WLf/Gj
bluDjSkj8a0/JfHoqYUm8Kyy0YPPMRWCn9UgkzD+GOQbFeYIDbc5nYkPuRCqWP1W
dnTdHrJQlu5IQdZcpqWWYZetwUe3YMc8pbbSw8ZWh2OMcOiu1KVss8Eze4UR2zV4
PlgBdQ6mS5xL8mPsD2+YMOgGdwYgXgp1S8On+sGcLnm/QNMTZ45IyEcXZbWm6AAJ
ozUKx5RAygoDNQedVT3srks7+GfqKelLMu4IN5c9etex5GjEwizl2F0FsxqUA0jA
fj8+fl72f1gdFEloieh4fTN8WJc1OGsfneJZbMJaR35fzpeg6TXpMSGDwL8Zoicv
l1enNMhcJ63TI4KgpZ8z9X4+6F3gn/sBVFwyKjCtjE6SdiA9+ByCf+kw2GZn9p/S
nSFVHktVH0PNeXwWsrx1ci1FfhXQr/oJcvRC5wDdFnzm0BcKK7j6r9l+cNh28LN9
THkslovpVVtayO9Mgcjc7vxD8qRNEQjgAeW7ekDUhBV/JSbBkzZdG13un2NVAETr
6RlXciLA7tBag0PruirOoPNROpKLY75Viz5ElTJfJSuvGNxR9yCqEhPpBi7Tqdor
4xInbYn7E41zMvlDkVsOZE2+R084JiLwa/tn/J10FvYxk1tNlhgDgFvcYCKxFifD
ZikULbX4MqlR9wnNq+zelJqiFiCGCmbSAuODiZa98+dkKTib3bVvo1EIGDQZK6Tg
fgwCB8N1hA8J2thsB5+SmXOHAon1nFdSjv3Ny63t9LkjMneZi0Pc6Go5fuOnDQtV
l269foPf2B2MR//WqdynhevKGEPcM4yk6Ka9jbwR6iDZsURuZJYdbLNezK8EPXxB
oI7JatyXhtvh9aDFcguLh+TG7y0Uchg2Su5Q+k5/czc9Qe/99bZUZ3rx5II/n0F+
tIfcRy/jp99JdVKDn1Cb5ykR35z5oFXjMJfMf2/L+mrd+AgF1mdPA4DDkkHc/PIv
2CErqmYsxsNRf0WriINO4PjzmtdtPYaOWFXZwqVmqmS+PJ5vx872/eiyXYFlCaD6
CAMqXGE1lyo3pmh25yO3epCrsaYcARgadq0ron1bKf7KRyP4gCZGWwIP3jLZvpDf
yBKyJLqJo2NCse8RlcobCMpv8HDBrzmwkqIyKR3m+yEmwJ3NBp4smR2fDxoAlYWx
kaMfWVJbYSRJ84YDkYS1HCKHPqLqo29gIUFkrydmGgyq/giUBx5CPPwNIsHzJcww
L3UvJkt7Fv1bJBO229WfO/wg30tcRzYbHMKSaODxfZs6f/GB/UwTMwvgBtsNZIsp
PV+8tZw/kx3JAv5IQ+SZdA==
`protect END_PROTECTED
