`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W5+8QudD/n6gZXPh2lDfLz9F8ymK0LX0V3SAw8hEVe36AlPPPJgFN/O+CUQmBWr6
56U5cWK+AI4sR+8N1bWaBC9oAbYhURBoaFPr5t2dk6nXmt4s/mbCQ1grV122qIQt
W4pDJx+LQ+8h9wLmIQyIwBWfz2sxfGpe9dx6cnFBUGb49IVjswOB4LIMPQkJqMxG
DziNwUZmqz/NmiX0+7lAAZFB8jMyOkFPH4xM2UJoeJADY4r2LvB9Vd6psWsjR3Lp
b6j8YwAbbpwixllmb1T0rqbB4t+DVN2gzE5GHbK5Ip/vhRh5ZtrEt1sF2IixV4Nh
CEObrggMH4kYV4BwE5tI13zxMDNKWcq83POovELgS7+OWCfOe0hL4JtjQtR02Pl3
a41A7H8SHSK30+4Xo63eG9eqcxU983WkjhtZXOdsnaJm7p2E2tm3IzCH+b6SudPi
YEsPBRQ+8F3ei6RaQIiS1gZpJPAt8HFQZtTWj82G5PZlGrM2P5GcD/ZysWLCctFW
Bp7W+sf/Ijjsyl/EZ1jGunk85Sva0VOn5aMpLWGSP0piTtAktjH8OqEh+Aoo+3QE
EuOKxAvlpWii8tDgZN+3dQ==
`protect END_PROTECTED
