`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1s/YUm14twK4Sdxc/BS8f11Gbsn/KbLCVpPqKx/m0pALbZCm4PJv1aqT/cuklqNA
PCkF3JA8jCPrTbgXY5oYY3L/nO9t88Tts0jbgGbszIuZauNS1Iz/k8xVtDf9slnk
bkttby+6/u+9y8p1Mq4zIY3+0hanFRT/n+91YW9WC8wPiApMxwB9h2Au+0mlCQ6Y
poHdVqJ+T065KyDop0nmmhldyhMBdBFvUm2JV4tZwz7Dec9zg+NEO1HYUG9xduaz
WUBSCFtCesvi3A+THEvQkMrkKuemAxe0cIHI146dJu5rvRacGFkqa30zgXTpZ8bA
hVpvB1EtTpwm/EyGdnHoP+eH5yoLQJzzhDcCTQArGVwlHnbzZBX8X28ZQdrReu3q
g9zChrRHPjBbk8l3LwezsO7bVnV78KqivHXWiSQt+vH95IpKNxn7tf+Qhb0jE5SR
ECwXzmnVazv/rb60ZXjV9+e2743qT2CdXX9GSZ88KsUG4fbakROwCHFRGAoFQwk7
qQlvqaEZ5R5yAhrFFMLnl53aQ1+p8HhYSXZYG51jiYmKZanm4b+m2CbIUWJFAXEn
a1nCwhhOb+cEsugofua+Yap66rySrE35yLNvOK+eXmqQUx7oY1NrGeCfcYEcRJ0A
40J4MKDxYoubUJ3ITz+g8IsUKPPSjp4E95cSABI/l5IvG8/Cln4feHrDmP/1eDzt
LjMKzI1EOd/bmPBGA/i8WcB6kHFVL5xgUARLUWSX2xd7m+Au5VTQ4Ny4hBVJUfaG
fogrK9vkP89wDzl7vcf0jcoVxAeZweKKoaf4SuQii+OYX0DLnzaajSwSW5gH7eY8
kWuDH9eouHyZFJHq5rGNuDhbF7o/52/lOMq9v1D6c8tPld8eP9uhJQZNmJKGP8Ty
UjHozLpRP4YTYOgPHehl+j10Rbg6pKHu1PzHRbl87VT1LNNwcmQrh+SVIFbfzhTg
bH1t7oSylhftkmAgrVQba8tsshvQkyq7F2Yfp5T+eAHqaThR3Sen1S+hotJ7KA89
FrNGEV71Vfp9CpSlJ5+cSs3TGA+opjjDdce1f7+lnDItBwvD4vQBLUKrvOdPXBcL
DY3P2FUf3gwkNmR6DYv4Hvkd43cqaQpW+U5Gmqz1P03mIUDB2+E1PjSCy+148aQr
h/nsaqpiObbkYaZfSac1wrJg9vblvK8kz3LWn4LzK6GL9yM/g+Z+r9FIubXtRoTk
lfTnn9PZtm68y7lucJAEjSdr6xr/oh9KAyos97u15mG5g9VQHQfBYzjxnZPxnojV
Xl+EVpqlLFzuC0MQB4a38Qu8iR0K2220pWTD76OjaN/b9Ay5yPIioxir/GTPiZB+
RSe/iRHx954wghMeCW2xWsvnfdtwq5jxJ35JROOb9ym6JDGuqgCMWI/DqKrmn64D
KdaMLXxCL2eN0/QIexM5Q6/NE8fARZIXZxVfLYdz21SN91xvgrSDOxSqsqpFt3c0
fTk2Rwyg5pW7RLghYrRi3g2z9YXsFprzr+PeLqvQf869m96RltHZXfp4mXVZ0r5g
1B1BlGw6JXlSM8UPeSZvyXaFcQtr4g+KP4YtF8VtojIC5iuPaUAXt01sfI2B9rnL
ALEchGwdonQCWccPbwvAyh86g155mfQ6gH1hckAyQiLRaAYbOhOhOfo/+oXolmGP
g52KfjHmfOQGiu9G1oBD3zlvhEg68ZsSyheQ9ATj9LuAh0uKv6KsaP+B0OjBOyPj
LxnqnKhcHSpdDyZbO/d2NYEMAs1AcAwUc65W4M0zPbeXi4wuwDNE8dXxdV3EPJtw
vu5Ya1saMzVDOchUygCXg0W+uPHG+p7DM8eOZ/FflEmWOdk3iM8FUeku+HCDreDM
vC40TS8f/tjkW48IijRKvQGordNfHmJDm/9d+FEtC/ZXX4HakQjr4jpvdI4vwVbe
RLDWMRaJinQ3sEDbe+Hfzj/ALQBGhmoqNLajzhHoETn61YlsyaOYeRszgCyvWaDM
SgtM5vyrbet90HeYaxPknv/zlYkajP88Y7CQphVSAZXXb0coZ+FEe/3cUq/744bJ
kgFaFcSIBU6owZrx1HFebr4yG6g4DlK/wq7dW6xukZEaarPj4H0weoEa8oy+ZJvZ
V6IQ7bIv2OjOrAwXIkmPDA0PrtSjAdxn6UzTAhonA8dV5oYUhbK+AeRRBwApcqAD
unrvb8Nfe8pxh4Hbapre/CUkIrfi+bFzDJSsvW8EyJrI3flAMjR+EFvK6+lr3duu
3l7eBLetSOtWOdo6HTLZbfFNP3tjtVqUh4Gv6GqLS7z5Yu3Sv1rNewv4r8M9Povc
DRmy59OPcYyp8Fzq1c3n592+xCprhXhapo5bHf6CYqSOe3u6NqH9cQxm8Wb+VTXB
v3nBbCcT3Ai4P5taTDJTyX0QcRtETyYZ6gInoSjPtAGB4mrQBuaCvYm5upisiok3
C0NTkS43oZvq55V9x4/WqejsuRKv2DsE7lYfbm/ZqQxG1I1fH7AIxKcGzbTbSJmh
IRADUksfdVX+kTon8XtrT+FVDRzxmWB3+7rM3lR4QCR1Qo2uNbijNmZhGilplWKn
cwC2u88aZA4jW0GMqZ6YvZviVUuSMU3gjJGXCyp6/XXCdAjtjqNj35hcqnJDPfwr
CX1Ez2zZGtgquE/4Q89z6fI6UmxjpyXSMYBwq6Gm6UtjObPpnnnRh28rDZazPwip
CJtVLOWoFYrECd7DZNktd3k3RxriBU+YNZMMabq4sSeFPCRItK6GlieU2gGAWTDR
ePBBlM61KBJ9j+XsRkwmeWOFrWgLs10kjLPyWxhpE9+A3c+RxtybmXsG5Jmsqcop
IEpX9zLLYqHjGkUNBKfkwfV/mDCpUiGRrsJpcscrkrJlsLUEvSvzN3Lq5H0ou/2A
+yRbfEQUOWY42rO0hKSB0uG+Cbcn6pfEl8+0CS0M3sMud7thJ8kx9+iClgnCwyUP
QepdHpcmV1SI3XZ4xkAaVvGF8HjD4uHmiUUWGPakFR86BK7wOseqfmSYLMk0QOBO
HtfLLlzFu21/gT+13sLDH7Nne1RBml+FtWkbIEGAyOqH9jbuWUlik/Q4OY3CWLxn
fqFaNPzCnXNdSS52wtCGKSXGLNVyRqee+bJYY1JOBeqkIbZeVIKisHWx1996EJvp
PI7j1cuazuEhwyZLhDxFUST+IjkbrrL1hB5IX4pu5qRCcY65sjVsvdaZaO8Hgir2
H/MoUy6O8mc2//DM/QuEgPwQWRY8eudcI6/DFD5dLF9OOjofY2/jXKdvTcbM3xa9
+mJBOc8sRbNfKQ7lNnW88Cbl7UOSFxOcF5/jVQ6rCEbecSDcQ+WzCKQv8HDWOAEi
yoq1lkLUyqjHC2FMK8SJB5J+b/ako1CPDglArMr9XR42EynYo9DpWNp2IAspCPjJ
WYiaXekLfDRWqsVhH2XCrWuz8MSgBTt0/28pr8ObWyr98fV4naLvyj7RUBbtmz39
S1VpvkKkV1P+QwlhSRD6rVbQ9r9iWU7eP8UOzVeeQzRzfAfpefizNShog/etqV+S
Fx7mTPZSPzvw9ikc9TsfcMklrqJgRTH5qsrKUInWrYf9ckbG1WgyLMVwUMiwLi1Z
OI7ct/mxNwAO6MdRVkH8SPM1pMnP76dxzMNgg+Fv/wkAamb9jwfkYliOpRGFVw9V
dczhCN0qOaYTOtEFyybVAxsUJcH8AuGmKkb1rMOv5F3SqpQCszss7zA7gTZ69nCx
icy+VI61zxbSxDnGT22EmVzNyTVZHj10+dngbxKAZhyP6Nc8P6knG/TBUH46wEg1
peu93D6s8Qxpln0DuiozTlLm9pvgo8QPnzQEPn7qkc4FegFcZ6lC42rOQ/bI9EzU
7yl6hV6ZgQj+CG423YR48Q2dScyzD1G7WJre58XonnX/zAvBJgh0wju5BR5C8VDv
motFyz4gqWiM9+jjK5CHOheEdy7zjgYktJwgrMWT/uUPNOzPFCz+6XjPDRzjfiib
JSU35e3lznFOjQTG1UNoF2hJqkKWPzCF9ItolYQ3v3A58M6xboaJsez+1OGonynX
KChZoOQ9jYH6uQmDWe+NjnwdZVPQBPrIIsLQ9gpkNbVujOD+YnT3lqVvARP5JdxB
oKJsmMTik82cbZ+scvO3o3nDqjEC+IM8ZgDRudEsaQXEgH4GcDo/x379ayq74ZIZ
ItI3QvpsdulafnveyE+bp2FkhK+muC4JECvTJGmbtzVzHCGRdJEIQ/c+AzO0iyUA
6LKrourDIYxhVpuxBsEStiCgbzE65y4hyDdOKBylEjSfwNhbd9dG7WgN2LFjaYNE
CpftDgkfg+orxyPpSupRGRAw8QcDV64NlBT0gjlEOeCsrkaZ3fhEDN5BEWOOwCef
YnO5zs1bKmlMKrsGuJKbfzEcmMOPuor6Nue2csoKEA/lUnIXDzt6H9lSbntLVfk3
6jF19T+4E/NN92my7YHB/g9qwZ9XtJzvWBLbKzzlKhncxVS0G+/MznRsmil1B8/X
/6C9Dl5LjCzu/ePbE6ZW9pgLwcsGlBbqqTTL8qGEbIG0+DC6FaxtvyCccF5iyS3c
i0KXHDzqmDytMJDJ3aL9JUcP8YB6OjvOr+Yx0uBRcFRu7wJUcESaJrWlLCV1WVF2
bg9yjjIVP7IRHvMdIXldFN0VxwouSam3k98RQpdzXpfdG3OiBKkLeszVpznjrHVU
zljCu2nLLXUVI6Ikj3lOCXD6AmM8sBzIYhqGQhPD8kGZC2zZSn1HLcaPq59gErhb
AVyYyk3IiU8kw59ijHZemKSnuOiNvcdT5gyPp9Nk8Nypd5MprMeyr7lLjekWBikA
P0fBvyUsgkriIQLpv2DXWVYizFtoDfbaBsU4ATHZZYLclZ5ghAjHOHI78wLyIyXH
pdzfCgo8UBLhJUjIRMY9HeE9X00gRtBXV1JpfdOTw2JEUai8peiI5GZOvhv6hSjf
uNqare99IGRg4UXWa2dkqJlUMPEykW9btR+ThsZUJxAz8jQP60k8g8aBEyLtfwiq
GEedQxXpbWPnPM9UPhqn/WKoJL5Ly39AdZjR4fN5mgXT4EsClQxB/PehzBUjJS9u
LK+rblM7pg+OaMza/cDNlNviFSuw5eSKJHbnJz3jDv8IakrwN1KLGkinEusNhKyF
IZpfV3qrA9rgL67VpKRVrizMGu6gZFHfDxXA9V+NWG2ETyoSJpZwIFpi0o0dQdAU
L1tno5v7M+ztqoOB4yXhbrgG8U4oFFPYZApk0LOU11R1v7YFF73vkEtHBZVzaw7E
U08ULGcApkRDcqC04nIkPzLeti70eF6ZoecKNP5XybpUvumW7UABPDU0zaCOMk6V
4jquNoGNrcs7ahjCNpbEsDxQCJ3YDKSvHWDSoGvwsv0iEPMddfbRoSk/vwOcUclN
qerT98B5ymGKZRTLCXVhUdb9po8vH3jPzmyB6l3YBa2lVqcuXaMcvPtHrsFgAMp8
//wPeQhgmBD/mrUdtXv38g7QWA+HQF5n+41dWA6tbIF3t73DTVY4qRHlG+mtXVgx
Qz7n6sMi4SJupP4QQ7bN666/W0q4FfFSt9mdGadWFib7gDm3VqBLVCbDIJsGR0IR
3J2mgSMLTvf23K54T7NwB8L/m7VqTBuAXhrbKJLXYOj9eaSkNHELTEF2pIHwbGQ9
Ee9wcOaYtkYf2WaM7emd9W/HNCeFINHD2eA0+TuLlFXnNI8oiq8vM2GhRxmpSqHN
5wOjAzf3peI92b3qqTpL7H7GHLR0ZaYZFJMlmEWZxjkOivxawBSs4A18gAwbOicN
VpkKAycJEa3C382qWkx1S8oUYRz9jpDwDgbw/seqVlJ6eWmlDeOVoxs6zNhtclBo
QMOwI+EzBYqwQHbGPerw1UNRiyHGULKW32CBrpYpPhbGkE5XWeDg7YrNtMP4LFXC
ewyb/V0ayD++89v4g6YsoQWrkShQAUHpXmQOXMJ7yZVLzcys0UH8a29qBTAHthvF
cU2rgA+D5BtO8rrUiFctp+dY8G+fvrn+9mf8UEdlqoHEs2UjiS5jEKyO8NbHt4cD
WGElYTbJt58ad37EtRiG9JlHuDlaPyJRRpLSawaDLAdy3qpsXEinhU6msg4f1liM
FR4nRShGAi+jGgJSnlwat0ZMNqwN1MLT1Qp1qoYePMd5DJgXyR5KQKbIjeNS6Z//
VvhXg+LWIsGVH05dq0/o5++hxjpPsDMkDBqm+fp912IoGOmaGs5d3Mz05sxwx05k
FLMdueb6n+cdw/YxHhs12RNdMYplB18SOSK0n+RWBB0lTB6sRs/ZjEbxhcV+WWYU
qZHfgN+Y8LhJjJYi8Z53In+zp7zXcUCFM3XjRSr5zGPd3z//XlOG5hNImpDyLlB8
mlu2/5Y5Bt+D6w5eio2Lx15uPblLGqeACFI05MLJyvk7Yh3wMFV9yfK9+vsYUo4D
6gBVDpjVJ+YZ3addmMpLgOZ7WLxVmAu3IJ9JnTqMOkpczebdStWvqaMo/uMwOCCu
lqOP+uXUP72OnHDblZcNntzg/lwO9jlEzus8g3kjVan0NTC1g/584cn6uvAuWW66
fq4eDJcL0ncbPE3XWcr7Di9jfhKmz1cUlvFg5jeOmE01i7jRX12E8XL+uYQOrKue
fitbv4jziMPvC3Z7Qqgua9FlYitaEX/GjxJRBmbzClnagI9YXxJbg4tlsWEQrJyN
7B7nCdFM+PWKRSY1fOVyHkRGakdflUroJk2YO25V1ozA//vU66xrOUozYmNDLKs7
STm0pNZoj7cs0iNUtQ/stXjvXdWg2tAz0n6uUKy5s2FT2oKIVEAfYl1oVBsW4QaN
lzFg6YNFizXchfKCYaS5B8ogmksyWMGkwRECzevxxlKSMCAFDG0zy6bByVHQWTZY
SEPLnsLv7YQnRsxabkYcpVaOmI4+n7URWbqpm9OoI9CUzWgCcbuQjWcxnDroyD67
WOg2PxXuU/niH/Iq1A/94RdLa678rIsNdt1BaGlqOnBo6R5od6/dgHj9XZFiQ68b
HuWtJAPQl1YrPNR8DdFHell+z+SloaAvkfDmcv8Cu33setOPHYIo9ulOiaWDhO7/
nKiFP6LPCTy5FRPFvgyZZlv28p5JGFxGg6PcvMDM1xYH5duvDRy8PBYT+cQGl5CU
Hip7DBJqmYINveMFibou50FCMYJd7/zaQLYSvFmMkubBqSQq4z9bIkZ2DrNkPh2l
sSMEfhpEiZWY6/Tn3M5+rjaJ5DazzcUcZuBhXPIE/BpjQYDnx99B70RdYGdkGism
5VqAxj94n6V28mKGB42jy02/2wUuLfw+arF0f1lUs2ghpy8okbfTBwBkV72fDVP6
64TOda0tJWx1fWcHCuhl+Jy9GrXrJ0giq7RFmsfLvRBELSRuLpMti/a5qCClHjst
5QiIOkl8m8k6XNIlv1mVTByl7FHfJlNbvBqosqdXmsi9iWtQ0OLtIhBcW0ld5Xtf
br6baggpAU0e7NiwboqqnFNhvG8o070oMIYKdgnTdgfA7s7hIm/tSCIKBo5XVZrr
DasSQZMDTpEysNZwZi7ktomenO74+ro7D5Fgh5hUiSqPfqdYZgQRLcd1krh2bFbX
E3LCPACdMiJuKJPXywN4gH9g4gNsW7KAdnKsUeOQnod9DUZZ1rSwNMoPRBAv0xox
elFWy2zudKnL9JIyGiwA7kkrPO1GNGmxaXKoeOvJ0OpMf4gbthRIBZyhCkchhZnj
7yHx/lQGBljoZp7tibFdDLiwRp9xYR6YsCHuQY4ssSQ5K2UDKGWyYYkXXWoDPA8N
j0qLKK9vC4ppWdVf/VWSr1OYb4qzM1stHVkL/sqUKoiVDnkI9ykH6xO2DKt57sHi
Y1fSZXgbzRKBYVeMojZTCYt911peRzFQQE4yDWIt+aQh1+YyrBYQvKYjMutncRCU
os8Y5O/p4hMopcks+wXrA0slLyTwvgXIMb+umUAy0ZX+FP5FxTlvsZNG9GbRmi08
wZJ/QsgNRGL1m1fCNyihVzHWQ9ks3J2w5T6h7PJo/LN3A/GLloW0HgbtoXdGY+zF
7CalIf3bGcTA0DRSvub7dY5A4labdIjUo44I0oL1MuUXmszFubnkyGCKpJI2K13N
2B73oRsnIQT4JCQtDkBvR2irz1Wp0+noN2mApx0amaWXsnAZjBueBAobhtXNeYF3
wfDQMjUKxJVr4FaV6xJej8eoetHlKr5Bm7BOBzxZ3VTQS3KILPkZgONfGe2HTp0y
4MdfKI8bVEeQIapqjmbHXsIkZIGTDcUOubN1O5gQxhzrSTukR3EHzYJMdGOgknv5
DLeJmIyz1o76cCGEP/k2DHvbnd1iuM4QSOb2OGyCmdOZCe+Aka438caestR37ich
MNRw4MLIoY/Bk9Va064O8esXL70nIbCZNJqOt0r7Sd1Rzy7k5EItXZJb9abm9OP2
f5HObC4jKOHw3kG+iUvkLIfPjCXV4BHFOTxqFiXgQWW8Zy5TXY7CqjEWbLY98w3j
o/pVBuwktcmdzxCVBdhehBu1eiRx7pDLEYpRmvsspqLNbA+MuPahMvFdbO+Tel6X
JLf6I4N1OfcNNwYATk6s81/21GNFdJ3VPTgOzgjDR/TEkvlNfvgaNkh9LkOHKx1Y
1nA+BM54eWlKs3bxvUUY3cRVEBm1YGDnDIodulCPxuSXcs/6BmK/qiLhp5id1Hw6
olUZgUdXHc05cowC9cYLSjYZfthPb00lwaPsqTFgykhBMGp4AbwthsuikA8pGfIB
8Xu9M6DjoftEbjYcDfQnXgDUNANfvcSNwIsh7i8KQ1ino/IoXeFSLdE371874tis
iaUN2oOmPUbT0jJPKm3Sg/qOp6alsFOG10ql3wwcgaWeba7KfENy8vSEmESPOJ8F
pMM8pOgD8yG841Sja8Gphlv26E5v2PQhHmYOHAvP2GQiUqjp6rb+ZZ4vGy8d2/ig
YZtPwiuN5rc7sqFfNFZ/ZTKMFN2cfBRyCRMtG4moud1aykFC+tNEFEFTZ7m0VxSO
r/lf6NwzNVxZde5D+RVGeab60Hx9GWqLh02yKYC5Z203S6qogPx2Kzi286mwoKCh
GffYX25A+sQRztkMCE3tNJ5TsF3sDvf08MqkH2Th7oCLrU4DxTbIc//idY7WApfV
KGFWLv9YZzAO371w64xZOAmEBLqFlDsgY+65DxRD7GuputpIHJCgrWfKDAJlZEjZ
KAPaWQ5+I9oRHbhRCKbpAAiSMcAeOpyzBNR1iX5cYEaD5f9IY7KYjufmhHBREp5h
2PRT+elEww2sJrAL2UtIIM9Py9DRQ9j46I55P8C/NUIkV+sBznB+VxCEBl/aG/9b
xXp831mc2bmWn6DHsFF2/qU8vayPwuCTvCIckBGAr50Q+Uzsim+QvjgXq/wgpEPR
Se3Xr3TCBzoEKXPSCheCWPw5OUC+LcG0hVMgB9GbDamm2uRpu8xqMjWBpoI4g4hH
RlEdAwYbWnfnehK0pToFViEtBAxPemveQgO8B6oYezjDF3YswZruSrxIga5ZoJov
Ekm799YLemTJZ1zu86YDwePlmMnGr80VISEg/C3fbPeoZ4pL32Fjtzj/v5Sufq85
T/RaTClgNI907Ai0Wmb96dko9zKRSv8AIcVDM5TOCEb9G1mZttBedPyVLUFfZ2hc
kjlb7iLrtM7gRITOG1Lg4MqXG3DuBkp8rhRGlCi0nF7TOJCdwVIAM1Kfmf92tAvQ
TMTvcjMY+ltmGWYLlsPq2aq55C0B/H50nU7zX+DLKg2hU8eRp2zGtN9n77T1ixR1
iM6zBG5j7YStZ9k14cQ9DAKnQ9BXVWLJfDBcUOHGr1w8sRwQR/0TeK8xnz7JgZee
rQGqlIvqHvvVZD8olpQ5VlTsY20sErI43F/iR2e3p/O+2zlJgabAed/JsPw4VRaN
CXz32rbDbGhf/CeJLNEr5VWmsu2AsUbaVqEJo2ShwbxN2vmbHtpNb11jrWE15Wyc
0wUDc73EJ0hy/R+uOXH7P21doemy2SZGLNill8saDAeDg2L/aNBD5zc73BtL2XmR
3MaRswcvkFcDgHTGz+0pKatwpq9ireCxWXAx5s7LMGJIYKOiA+lL4rGqCt63aqh1
lP8LZ34+K953GOlxGvotRAEKg5hzOB6LNGYqWgrYz0DZNIJxBIp666ArJqKRtdtq
uGClctNNNmO0ApMufnsgdY3z5I57HOjU/bsvUBWE9dzHYVDbk0HiQ4iRHg6Glt0V
K/UZoYzLjamb7syo9cieOkQx8ueaTQPfy09TWL66vG4j3KF3SwgV/WqcmmhtEgFa
0cJrWsTUciYQE16jenueXeDPBKqqbmA4k7M2KijMmGUMMFK5u+GVyPt0OSLBxy6C
5i0MZxP6oqsh3FYQXAXWCuMIWichd2O7iPivhNri7UmQYoSPr1YmM3bo4xLt4YVn
I8Gzw4/Bd+yRByS5K/8FrwAOfvZkwmDqBvQXkopEXQMXZ2eVh4TQsb1sxkbncKuA
2m6IlCEXGy4vduEiujOFfdY0LRy6yK1/v/gBntlmmiPR1YFwbLrFLlKtGlBRDYFV
E4jDEDAA7uD0fscVM1bA/mnI9gxnuud//GTiIySevpcx8oQ3iLcy9Sp8y4y/UbXU
b2pFH/RoThvi8Ep7iKmoj0ra9m4oBbZ3rC/A4wthofeC5z/FYr4s7apVHMP3KODT
iHBTj0yE6oH27LXL3LEaRzknTajnNClHmIfMOKGxSnQ6EcgwEWwdrUcgjsFaYLpt
1kHUrgOlap9oa8RQEQgt+BJQ9oJz0DeA5EkgH7eNED6I4ELHqPgpjxfTucQi78Mi
tEPI9Ual0iCI7rdVe+qo5+KPXetNqCanSCVQaenFoQ9Pi4ZMqT2GsvoJHnsHnJ8h
BgnCy5ov5bVxcdCLQnWlvP4JM0faIJlQqFewQJU5o+l5J3eRpHIW349ZOrmrBbSU
J2OHkdZkXa1uu/j8iCQPZKndJsYY3a4np/Ebrt08iTdU4ois8ycwMzEUeHJnorOw
tItdzPcSPr1v3UZSx6OjTY1leVyZ2ZTClciDOFZQ5XzutTaJVSXB7cgU1YcgZvkn
IX44Org9biREhMw5aGE9jiwcVY5q7OFRfaccFEQQKIPr2MOchCzC9mewh7iuI+LH
/nxUW295m9qIFyfbpgs8aXWn4Oosazgylmo7oyQCUCScdm+qEADeSdm3h6cum6Xf
IpLNNWKjEAg+kYH/pqMznshdtu9nzfdlSS80YKXsYB7vGpLxBfYmcEPMppC7NP7Z
paV+v7092lj3qXK8lY8HKeIngGRKNjxnLNFvtWws+yDZdcDcv5IeTMvqW7hlMJGQ
52Nf2GlG60HLB0e3W33uI9HP4zHTX1RKuuW+VVctOlcGgCEc2MRwqJELw3Ke9EKD
uVkbfFI3zaH/EDgH+oIpDDQiYBeoHWVrH5cyStFHpglOXca6qZPJ6ptoJ6aB9m3K
fnf/fnI1MI097jIF0vr2f2Am0VR6FBlLF9GVdXbJijnkOrgMGrt4mJ2Cv0B0Dwjs
bavj22tfjGtlfpi23Stq7fRJ0ClSOJ7tE1Xe88lxOF6uf+InDyfBE3rNEbBKIBmX
mENB5iq2I2klH6pxIsoKQD4Ck5Xpa4gmCicoOt7zoc77hp7ZMxp92j318079Zm5a
wZJJYUeE+LstY24ycFIRvhAhmqElYzd7tpMNiCH7C0yw6O3Jr5kkn1F4FO0U4J0W
0SMpJqbwY9icyJor0F1CZGECZbiSA03ViT1OQ5Tsp3inGa0UGVH4ecubWrLSxb1J
GqG4CY2vXiljGlvbPkAdUywYGXiSs0SWnWQAeDHsdr6GKMJHRSfJpBn7VosQMrbV
J+dVoDfVHUs6bOofql9rfXetzjZ7vftIYQUqTRT7qX0x6zKr5nlEs77t+K5yRLl+
z5znb9Hm2wjc5l/Yhv2Sx7FiGUY6xureI3XIWZi0mVN2LCabUaIVO9pX6tWsVT0s
BO6kXxprsvhB9/dTKnpHv6ptGBGBMX1OVr4adD6aCOJT/qQOvfrdb8XnicKjF6IK
5fVQ1OO1GkcVsMG+0vH9tF6+gmZHjbxqhEYtX9JEKVzJveF8uyomtPQwJG9W21Zf
xaLrqVS5k0DPawnABqVamGZodvUzPlgzuN774N4zYDePEfSPGwXkIVuGBQDHuNlG
CB28kFcAKUoSm/jfQDx2si7dqAK/Tp3BRgBz22kfSjNyf77BJ1+KrBg3MB/ic5ZO
mko2kGl4Xcl0dhzSlGLvIyZEA/LAUQObTtksdmjP15Qnlc1LZfKP2Xw4UtPn05NN
qVu5Y1ADUJLPaQSt1y9uo7npKV3V01wIE+U/tTzbPQtu6ntif3kT8Eyp8SxXJbQK
x9w3lbL7li4l3YuQZJOb2ijJL4Z9FARzH9F3S1EsCreBEKYUsYyAszjUppwNe/3t
OFUjEieCrk1bbI2aziYb1u6FSUNOJsz6As8agMQKmY89LmWEC07zTmM9SK6Bg5yX
6n563yluA7sCYgXC19faucbb4rnLolwpCpf5hKWregQRgXWY1nc/PZffASoLdWVm
tE8FXtMMmIGP7eysoSsf5/B14OQAHPX7o0hgmhiRcZLQ1n1ERSGFvGvTP4kbI1Ds
SJDEJg9/33XWYWjaK9S33+Vrl/ynZxMnBp1Y0FUkT2jRlMJqIQcoW8tFDVlooqne
H84qHvS3deXhbFJe/I0oXss0/q+IlrVTEux4MyWr1euzWBn865oHwp1YpXFsijng
VfxetzilEHwFuQO0xhHMIEc90YZ/BRGKCtr0Jf2lo+y0/Uchf0GodKkwDJwRTcHR
Cb4nfbzv7cFnTzo8PqBxFgtdM315a54//2jMEQ6163k2jzS97ty3RZQmV89/s8B9
J2ZxYZpemSNr3BhQLXKG3nrkAW588JWLEm7ZJqDzE1KNhZAT+BTUGAU9HnJkQUB+
WXMKNA6UaEnV3/IyAErbknK55q68RAoZbJHONMttQPWi3t5aD0aOdYVLdbTtiENE
i7J0J34R7S+LX4B49YF5K3SnnJTmb9ERFDAkkMlLH9IWXBE3WzAzICpsGddwpXIk
FAeZRQsNWSKFtVXXOl4BjB+qWyQ8D0J5q69flY+LWW6dsY4X62OHaFLNnurRwGE2
zBaz+jLUsZSawxqXIHEyaj1OHRcIDIXvamrjTrUQWQygpY1icuJhQ+6e2zculfvD
j8aXLbSpgND32nZUu+9Z6lOQvBk48tkO4eI2MqroZ8KHDDr1eX+YWEoCrK4jo6rB
IKKmCVEGajS984z8TjcgRzox7AVounF+1pweRrw4G1Ga4WF4+bp/2d5spkrwrzhO
6IxcY9OF9QgcIiLvMDJBccgLz1DqJY3xeBKa1adKt1biWwz9W595E8HmoSReDLw1
5vPKJiAm8jBdK4GvVtq8Dprfjj0f4qcw/5PdkcBZ0dJtrVlyzSD9o3F17zJkCQtj
JINK7UQlJw7E6q2z8r5f0jl53gdhXwWkWbFFgLio6fhtHukTqoLiec5vZqDdhdWF
OlCCK02/u5StoZGEsk1gXsKecHUJ/6E5miueUwyBi9AhSkTGlzXTTbhyibYX9Cld
3M94+edQzOXw/nS+lSaqVkLGzfhsVDCgY2h3gkVEezaOn2OBgqDIWN3rzJ24WyMM
W61qGXMgyHBT+ghiiDEtkwaRmCd57+jgdMVAdNoQVjLkK4h3iEFos7S+6dTkNw3m
wo+NwvA7lNo9ZbWtGenavGvMCukGms93kaSbxTYJIAf+S9DUinpf+jGZWmJn5hsu
KlIdWdCa0T3ArCi8ni4bryGGcCngiAVaNSRRrLa3JJhnDx2hFffNxrigCWqhyUvW
hPv7zIrS2Pxq0F3OamsgMEXr+9fWILVEI2nb3Uwe41xAPtW2Z2o7dS3tGB3Iobdi
12JNnYRxR5bBIXskHPEHx++u/YMpW4SZ3cSub/u+YSw9u0C22ZPyqjcmVGto15tb
QbG+EOdz/d2lrTft6bHFPU1z+H8K2cXTqforeCSI117N6+MpgyYxhX+vMcIMCv3H
crqA/a/NLGGE/zBOWCt2g38etMVMxxcz4NL9kzbFmXYe15CsAi5KwbQsmx9vtvXO
sNVKYy8VaGmFwKFCvIEI5sjbXoxA2bZ4Y5dXRBBkGHqWMW4q7+SKwucgzzdciDjx
FSfEJmqrIG2A/jMqqiKIssai8DzDV2uhIvk7YjX+5y+wTtXeloJ1B1Gxq3Gssb0h
KG0neqnzK6p4CZmPsiDZckyWyn3lX5vOX6qGqjLsi8lHW98vcnnkfc/dZxZYVBAg
BPbg4Lbuu7RQCn3QLGm34RTXapgEiyfvpMbbOLlOSBEH/eYc5PrT3982g7aEbY/r
h9k56vn45OPQKILA5iZG3J8dSDK1URWt6qQGOs/G8H8FfrODeuXY8OKDqB4SSQeG
Dz8qa85DCpHKPi7K/P5v6vfQeC59G6VbTZuYJmbiWkJhiDr03616r4DZOdbjfbls
NhYBWyoNV+PP0RnMFMQqpMIjHSLei4ibFICkrCGI/BqcLhJKHCW+K3ASlIt54SjD
fY5jWQp7tmEDymzmE32kc/hTbVci1f4uvuM7GMyV9jQhUqJJXKuZer9sSxE4zzk0
FWKmZeHW2WHQNyNB69l9eU0YRYxbSeCFcWY23dA8Xkcn7C2Q/2KSTxYRwy4oKOrx
2pmblUlphtmCkJsJHwBDAJgg6s9L9PwwzR16FHF5hEgERAlMMgY2NpUbXZFPr9nD
R1Z41+GUxD4Is9Lbh0I9N2C9WL6mpJq3NoHEtYq4nibPCEpjq1ZedTJUFOqdFPYf
C3hAJRuce+k9vWj55GuScgc2ULYXDbZgRrVLm7t1xz32B6wqI0/ty5vFvgYuk/xG
g4JphJIX2vnIIRUtlrBpG5maqkxrDT3gelLIxMe0Seb9QOVAkggur0tiOEeZRitP
rB9SMYI9cNZyZGRbRTRI/dRjm5wqZk/I4hRhZL+X/qrqt6v11FLzr2ZBknLD5GZ+
nzrPWSi7vw9V+8E3UtitEl7nAq2PjXMtDPhNWcwGa2y7F5MTKoJcX7ws7tLAqyBb
dF/DifmC9jgu8OoGxM6jVUyi7MIan5r5Q33DOfRZT57v+fW1bFamvs7q2quHxce7
lE/FU1Qsg9Ft0oIdVFUgHn+4AAnVmwNlFVzWMKjDmb8mL+X97t/HmX6S3mKg9MoB
/Mcu8T6qMA6C949pIfmKNhKy5QDzlTVF5RTXrnfKdfkTr4rZECNscyIAmYkDcHVJ
TP0bUA7uo/JMjhCZ/YIpBajG518dEnSx6FYxhaLZGxSBhXpP5eQZPbmRj4KWF8et
VNXGKNTrq+WlOETls4YjpiwPyj4jMT1uac16UQUQX/mqav0TNpt+Xz64S9/9nlzb
NjemzONPbzxSz2gSKkrxRayyMzfE1OubHKs7HIPWXHvSafkDSgP4UuUcVWPTaine
LXt12JWlCrwpI9RtEBhUCHttZ1WqB54Lg1HwSvfM+sB628O0gZW+zn+PSs+6blB6
VA0IEUC+l8P5V7ai5CXj3bJmglplPtl4xUGQfKBfr90mqD1CI3SwRlmETpbl12J3
glbW14Kkb+Qr7riUc4uzyRJAnzdwAi4RD585HWj43Uht+T8ztgxWaKMlUxLJ5V+r
RIulvWPTc/2/Ved0W7/7C8m9PZ6ucKMFIwUoJPDErNfRH8l+izy1hyzDq7zXlZTP
6IfhS/Ga4gnCpFGgxhFq2rljF7qWToZ0vqgmynhJ9NoMaGo6aR4K8E8hdIqlzhwW
WMa7N1MrVWSLXi94w/uCzrdUQDCEuaWeAJdhZfBDeNDNg7zW0um0c7TkhXqN9TCG
As8UPvfP6U3vlg/Z7KafO6PhDMy3ZQBwbc75kBIHuAbDEK+BDWSefOFNYe2e7KsT
+H6dQtMj8Knees4dxL27eEFDnOnmRonk4EXbccYiRa1hOBkTzZJNVeh7XfANZbBf
wGGcES4Lf1EQGsP6FVm0pgCy0Ztd/K2t+As7/eBXrQMZx5D+x5MsinD2FWb//dwk
pZMYYy949c0AC7dhYl1U7ElSyzCMFs4zoulOrEvhx4wwYEKzB7DV9rxb7krUbLAB
sGn4R+FMZqo6KwSUlZcLsLHP3LFI+usNLkMKrq60Bum6TGr86dVh/Pl7pHKU1cSi
Ku9FtTJbeM4cM1PErAa/08NaORklXRS8NboxkUCbS/kyJx4QE8+frLHIpHL1ibo4
VOZOt9pUgJIQx70ZMpgw9TvvwQ54Z11nZjZPSvQcZ3In+a+rRpHlsOkvpNnsOoDL
gwgsZ5/iJhGSooxsd+zuZXqsziYRxjSqxhLxEbT74YLhgyXI2khNdBddPWqPTBSy
SoSwwRhjRToblZDmosNA1PTvd0EayetHnL6JraUy+xrBCgNP87CaW07rJJW8l8Zh
WLes7RMkWalLVQ4yCM99GuWJZcRCS1wBEb1usRMmXU8oSSQ13uPoX4YsLM/iWdSh
hIYjju/uzi78Ml7x5MC3wn2AsEmp0+9QyQfSdHKQCeQrGNXBdg/M9TkTo4HVF4IT
yx3uwK54O8wUSQGqa6/deRX/xumRc8hS70aV5wV2OSGYYzQI9YvzkkTQvT3xaJas
CXT/Sqkmr7ys2Ftq6+LtLgyzXy5HWeHs4m2w0gmPBEi3Egot2sYgoefFBGaBgNBu
67YUL7FFp1NzxyxPUunjLxwkkXuTmQHLA7pXaRJj5qi7G1yFduQn9IrKtyVLN6y9
5Ap4/0146KKAbgCiDPpNFE1accednyIT7HsnNqCSBPq6pn8qn+l9m3l8GHaLnhnU
vznf3PCdH6zO5bpKIJ3uYqdSBBHTZqG5loyvRPOQU1ExfpVId6sXPVSojUOqdesw
xDpklCxkE1+7XkYI1o4ZCRk+kJuByIPrXy94cRpOGfzlnhPwemcl+qdC9aLAVF4n
5r1tfEPkcMscb00D3QA7ZGEDpwJFkNzJw4NBU7fMHzWNdSO8Sp+8X9gsR6CRaMGW
jeqVD9FuAK9dHCuDh3G72is9+4wacoraEo7qTio/ULMpDkv5aDGMBfse7auoMBr1
2FaWyaCyfsuml2DG/EMyJ7IzPpkWDvgKYSlo8D7f/h5ahG5dKj+g3dG4mp8JRqua
ItBMh+FhO7FImzOWy7t6jcZGqM9hAo5GEE9FCmO8pS7W0ndqk4tPYxQ0cUtMmtEk
VJ/+O7qvXRVE1Unn36Pzf9RrlgggrHg6LYs4jES2JxNwYwTQDIdCttaFZ8J5yO4r
iirxXPhK8WNp+Rco0+YAj2xMa9nbLqulJL7uWae2qz9B3anojWqr3WljomMv/MwP
RQ/RhZyZN4oYRi6pC9IjXthg8RM7rH4QRjDW1xT06ILOXi94xQQy5prjg40T9U6t
PKm8GvyN5LyACymGteFRH4JLFw9WOYsHSq9Qs4q6DoGpjNRHokb0ndWNtgR34R0H
DHcEe9eOgZNpFCi8gyHwxfkjc6OUKdOFt8mJZ52yLktVB6DEln11XCtV1uftbGT3
komlAidYTzc/Iu/ykY05FDsBUtXX4ga60KVd/PViRKp8PDjs/cf1soiH0IigIGHm
MqOzHqYHYgbimswgYMAU6QRwuIIpDGuxSB7Qm6fDJwXFj/cenXEaJ6ppsVUCeJBo
CDcquI7DM33ug3Uc3jhl6zC9UlxpY1/cLbODpX6JnvLaEzggNBOR5Uawm9mwv/8s
8kqgYbtk/LgORFgbYGfuhIS6yPzlnPlRp6BEJuPmFSHXN4d/6oq+EGV1yPjGuqc8
GTs31XU4tf9zNw8TD7JAE2EuPx1qDu0xay94agKvVYUBRUJLaXW6JjcP8p8MxcOU
9tSexaz/9MlmJ9VgjmDqYpwwuk0ZQbdbS4xF0HILXE/L/P20/05kDyYDc89Zq4Uu
+/s6ZFVGWJo7NnOGhb+az0Y19Z8EZUnYXAGYmJYtv+z1LvuDARpiQ0qh7w40XEDk
9DZNydXolY8XJc0KIYxkUMuWHIZq2IGC0oVKsTxSmBQIwnJXJGqDlZTUts5jHDtX
AlUixqnIr4WnrZY71lRySpXjEqxTJSxJGDb6z/zOe6nHmN6pTZhLYy9yaIT/cQ6k
yfaXXR7dqsXe1ecYrJGbPBiuPJ0Fu3gZJBnB2b1hSZBszIXQLUk11wQkte97cYrC
kT9k6ZbNZSDjsdPGTFzC5caI/cm0qvDTm1WHsmEosjGtx63jvlNcei301NIrnQw4
kSCHhCkjnpiKYDTa449vEQcIRzXSiIaPin/y6eEvbT/bKn1qN3FvDpVwI16zfJnq
7fynQDVNQZTJvuyzg8RkRTPP+VNt7xB42s5sn3AvotAVxKlJ9Xb3LGSG0z26c9Pi
8/j6ag9inAmdfIS0g1TAiiTkvyLG7qWq42hvBIqfB3wSqFVrFp1yJphFmUOjH7jt
dnhfs4CAeaZv1tyapRJVYDYMdFZzJo6dQxvHQGhcp5tqXIyjC+J792Jr3GBqCNT4
De29VYaWv6Y2wlUbALBKzPvrwtu9d47qyipf3TAjCRyU47ty+0WkiMoICpCkkRL5
OCbw5a48/vjzBVdxTmd2U7TW8HsXXGc8KZDo5ZU7xCPNlz6S9Xa0BNJvbIRiVS+J
4VgscSNebyU4+QuVfq0alKs4xnJaueJMpTK48WHw0H7aYnNRRyHR5k3LcbWXN1dH
F4z/yjq/SFMZ168U+PXCmccXs4u4lY17+ExmiR8sPt94H6/sgtjr/qdNfr/+Wd6b
rUZ773ZgQBnWpTtLblt7MBq/VvRetO7xd9/bkyrJeWJpeclc72pcYLb2giGiKMUe
BODbk5Z5Na2/9d6YbMjZp8X8xr7M0KqWG2MGFz4G+CoauzHSBqJJQVl8Sw3qC73B
0HmmnoWgAIpF4lTY+lt+0kK7ajNAFsXdIiIpZRrtKoNwDXkUPmFcep6yR0ufvtoM
qCkKWW+wITH6UesKTfW2QBGhNBi/JiVsaXBMyanfeRwWLZeUa3Wt1MR14WbjoXz3
S3X8bEU2RuHES2MaWLDiUbpxbNYlmdpZXoFGAH0NGIyXLC7q/Jp1Z79SVR2hTzOa
k01J6rEtpBnzQnYiRbrwufNed6gyIbi1UzNozvXYFsauFuyhER9Bk4DqANg4l3EB
KH+nOxpnUdRAt/s03F157n5eVS+AFXbhV/hkgB6VyPo/3hrAM9grfyOjfgqjGQs9
iMdEB7KvzoTWQezd9M175IpJBm11rWmK8RiOANeBgb6iU2UQb6wOQKLZtdyMHL/r
BENK5keSM9GO9ipoe3K8kTa2afOdDmHK9e9VLf0axmzJW9Tdd+ehDYiMTcVXbqJS
AhW82oKdD0mh9/ADgh/iOyLA7JSQBQeazVtQUGj1O+0XagqSEl/jmLa9Uk8HF/bz
6pquBUeiFxqJ8rFoco60MwWP1RvfR99zwD9WAOeqWOB+MfXQiOP1TNg5IvkqV/u6
b/yfRoZ7TcijgaJrdgz53h3XImPnJfduWpttmlmwus51JIeg0Q+6oKrEOi8na3ln
q+4jznaRz68HWTeNpzCe8tjawpkAr4sV3j0vq+MEwhOs72yCq4mcJX95H3iXzTJW
TV4TfW5NKK9TVKCrnxlq+v/1xyypmNq+izTjUBelUG2hf0vqDCL2m5GZ+HWgYWEW
acRoaNLq05p2SskZ+9qTo4Wx+00uEugBSG8wwLhvhNiLR/HjmpTcuc4yrxgmuLyS
LPEARfXqVDMImY/JL1evRQin29LKruju7eFXsGktTZ0SiEFt/26FMSp4LLfFAeZ1
nG1SE67D5LtRhcZkaKCKR5q2OLl2K0hM0lx9zPzimC4qMf7kJanWH0YMZMr9WH8A
/Nt15bzM1Tg/Aj+1bm1uvP5mgXuitNpDh6uwL0razBRdKyJQkdU5fHnNZbXUW+m2
w9dzsH3GtGeH+I2e5u9OBA+1CZUUEj11cunxf93MQZ4VtG271N8vSFDLkuRDt8fJ
3wg44pkvp7iP2/hTDGJapZ3i8JlgK/Sbcngu4T+5bRgPDyP7oejFexisroKjuo7g
96EDjL48fwTD2ta/OwRDUdkMW8IfNtQ8aKLQPbtFfD2bSNA9slGlNNK+netywzat
6oSjMD55NA9TgiL7PtNFqCZ7XBOHHPdy3SmZi0AQrR0lf1cZfVAjiTWqMvIci+tq
KQr5dB5g4VEPiynEsuZQHzTqC67uK4NzmSm7PuftykYKuga1ryFpjwduRSZtIlC5
EJzh/UnGu3w0mPYKbWZzqxWldrfAgjcZmgPrT7bcEOIqDpMOSFcWruDn4I4TPa0v
0SQl9mrCyISzrC3Yw66Bk4SdqXBlvxZcC8SgawWQW1et8Pvq7I7Y6NO7bMpFJbs0
NcP9F39R1ybICCRxTcERx9TBr8SVRiHy9Sjzgn7nti2dFVfSVpNDgPpoKwD6FAKT
t6RjnhgDEfSe237n+khF+Yi8CCok+JckBZ4/Ylw1uYYCXgB2u/7SJK7s/W12ElLm
oMCHYS9aQGK3BCKckCwcI1vRbFayhVSUMWFsaezF7RTG3DHiDFBdJHc+6NdpEaJe
SMU43rSuy7K2pLDIhA4AMlHd09uaDBTPSalw59mXtfvRAr4ExT5q7G5Ukg4Qubqi
i0X1aQKtznjwOc0UU/vFfaLUkwftqrv/b8N2rX79ZOkCmnuvl8OhKOqQ5nY4j/wA
EiiOHPS5WSfNVYXkH09PpTwPzU5uyaNu8vslvJzsdNByHi2lcdWdbOiRIVEqpQ+p
yaJ3d9koq+eyIKG8PTqodtjKpCvSMRy2gNNwvTIsvMNuWErdELvfyLCMPJEnLZUO
y5c0AsFqzScXEtWnqYaxF8ORLeuUUiICJxIuqvtzSps0LsDhITnPcSoFidOcpk2p
B9V6JSc9OVGktEpieJ5o8ouhD1E+tnvuK7DTqZV/XgIR/xoVYC8qpbSlO47RFfgI
dOMpSbJgBcnt64xEzYUFe+8zT9FBv+8srUMpn5ms+sSETSx1diXSLVfMh39EYPNI
BI12fZ1IrdJ1yzZkuuEbxER0qEakrACfbpohKd2OyIofBMcniO/I+0F1djHPi8o3
ew2JcBsXb8dGSWdYCMT1SY0fXPgwsDwx+KWnM10SBrYTkGIDdpTyGhhvPihiRPbB
wF8qHreH4DNq+b/Nwc5mtTGAamUWG4EiMn38tOc2pV2wX4JvaHUHh05lI1woNJa3
QAk7WZgwIPNAs9zza6I/tGDuOjp4R0ke1B+UvLVnTuz+ExB/f/giVAaXczkAayas
yxvxqDeRmvZayLoorcJMXS2Vkb3BObjj5djmgzwCIDnDUeDb8MtRaeh2eLpWBao8
EQONHnOxlpnUkiqasxfIwb13sIREtoeNxkbt+PyfrWt+ZWTwSMBu81hSPqSlh9pT
EpMT/4brHXOS2D01ptrlJg3SnBrH9ILDWM4n44C7s0pr29zqnOdwUZeWCxcCZuwD
IJokNbE5BRAXlTOQuw9Yfzp2qbLtGkAXd83L3F6EI4ZDu56aju1cj6BNqbLBkLBY
5WMjJK8DVEmFP7ToIqqya5ab4cQWuoVof7heFS4qjBmfnX+5DDiwOhNGXcq4oY7s
jMcITN5I1xzcGDZxiBLis4a0NOBI2Z2JvxOI5u+7A7nwDPoCm/EYffHSTYDwk99i
AbiAdLLpM4ufA87int+ujG2vlE+RCH5FD1Id/UkSBo9gz9Xu6mTjpuxC0caArWRv
wbkQRJIiS/3K+7jIGGLP8cZ22kB6zWCOQNbdQRwUpeLqeWYLJQ1a6A/Sz5fo5XxK
v7hwC+cziXE1Yvx3E6zBeFegBk+X1/nuiIhUjf438hNPLdGjHmUAB/gLWdyKVY5J
r1UI65w0VwFvnksKuvqTUyAs+Tqr3ubSKu254HquoAmZemmHfetC2k4k6q4ipqvg
LvfTlA04204yjEfNCohxQQ9TlQLNGC8ZfjduB1kTVT31hUzlGrhO6xVC4hQAM5W9
Y7136865GbElYn3qkdvmD5+xIjvSrNdIMD9IIl6hoYI8Pg8f4q7TVDIdqhc+ya1r
Zoizu7laLJ4KW8lhJAWDKJY32Uu8hI/5cksqQJj8eo6w/kERsY84MRuR6OK3s1X/
AYtkmHuVjo2RoX70f3koA8oADxdd/XiPIsuJdLfuFlF/jPbuwlKhlDYhnM5ACcwY
fKeu28KNejLNXM4xM1p0FeSxYUvfGYfC6cK2Dxr2rSo42kxfcJAaNWQhx2c+pSpU
mRydR2O5C4dkMJHwm83FMP3+loZxwU0eDAIIXqsnXvWa069l242y1NKjuoXbK+TF
xpdsURw4IE7iDLtQPjZQxCrJgJolgS2opDUlmAGdopfsCz1K6N9eFeybIiUUYHYP
BWqXluCCxQpH3rOC3qrNaKEmPNTCMBhHOTI4LF5B3ag3zE9Wrs7HCJ2KcZSy8z9k
xfjluZpQw+wIlj18DYu81Z71cuExjwasxkYYoKn6gnbhjMRpSXE9KupUcKrQbByR
94tlbtjIdYNFs1GQS9QqwoIcXonSw4k77sjmsllWZYtQU48M28DwkruUy1gIXOI1
gd4+J9Svn0jsg9gnFC8f5LGqcpPFCEI6ZumV+7vrCY5Q6UUiG+IR1NA5ymah2pFB
myuqjod5JaB0mMf3Kn3gj3QTnI4JWdSeARAEIavPb1cayo7oz5yGMJn92+Zd6ftZ
P+LIkfq3Bc1ZqUsoKCkSgiVJ7ROQl3Ig+5DTHsSNFS6On/qrn5zAj4B2kv4c1pN9
ShA7B+cLtHzF9fx45350eP8A9gv75UjVaGm3aMnKnSgn6VjUnG9iMigWsObaFEeq
myAcPn7hok7DgelJRf9i1YbNgt2k9i2Lt3kmjl0a6Cw7rIwffQtJb8IeXWCOB25e
DgD3lFxpky8mnHPmEEU0QynVGVJQIP8DSZJGNfofbWtJf2/iX8kYCohk7jxLaDe6
zIrePhocnyEwUu98ycao+lLBmFpYWivNDbsR3jiy2dHvOvnI/yyeFi0ezj+G2nQI
QVN45wjFyKLxqZs+xFQzVYI8cK0MMDrSLL9dkyF06AjIuD9Zp1SgD6IDxP2ZUYdr
Og23yPcf0rNuPA2LFCZPkbvQCVkLvErIj+yeq6RoTIMONHZNRK/UCZrmclROFhsm
UxW8Y/dIkmts9KIOAR9E7LAD9Q5ZVKZ+KjukeZN6dN4wHpGsp+6galjbftU5PXok
hQLg0+Zmihu9LhtzmpitKE0glSgYxulyfTHNo+0kNWu1aXYy5L5HN2KXu997XzFe
6OKkaxcJ3wxUZcuLMARIY0FZrDxaV6oShpel1b2dJZa2011vL5AtXaAo56f11DOD
P58WvfbS5r3u+T5U7q+htYbEvHRRRdxDB0+5c9X+tvScE7bBTvhIGFS+XvjZBuS0
Mcso16TlPLZ95oSKdeiFZIeWWq0/d9YuzknUlXdUGbsocyXCU2DSgJr2dssEbajs
qoxxg422WBh/9owqet2bM4+USYq5hoHdqs2VztBL5Uf3HmsjEzHaZH0B8fM0Ywk4
8e09zdf83URM72BMWbRQnbE5RPvDAEPE5SMlfPARhOXSifLvncQ5UdJmTumUFqip
HOSMuEktFLUmE4lOWiutuEatAKS+KTWS678yX42IjNNf4D8Iv2JO53bx8eyo2bJi
IaKJyUJ7mp43jjEMKEG+vQZBqDYhLq2ikCDNCJh3WS+99WDUd3U3ntsgkZ5vsQeQ
vFxtRspqE0Oa3fVqANzF3jpz3kfTIo0Bv7Eu5y842HjT/qZKwPVI2e+HDKQQmiQB
Z617Ou3w3sCHPbtmwdsaWXW6YykYjwrCUtnd7vBb6nIvq27JvcOCsyyoGNYszA/l
xs2m6I61TcatcJ1kafTS5iTa/kGJXQPqHlW/ob7yQ/b0G4xDETonJ+lmWzPDMbS8
4Vnr1zIpfElZ4KCX1uxrucdBY8+yjn13Dp1pEV6jzpYpEjrYOT9neAZz6qwCJAMk
iU/EqFD3SMJ8XlK8TKZ3XhvETy7TItzdB//RcVCzW1oRO3ujW2cacKL9aNN0hsm6
xkfGJKXiK6pmwwpK1diDNq4as+aVSTpDVmQMy38CR/CluNxAPbV+VWroEbo2AI86
3qbFu8nydo6oxwPZTIda4Qp0Tenu/YsRalnh4r0yCaywF6Nd95fxb64J3/Ko+sj5
MxEUHThShYZOzygLSB7HNVaVLym47eyf7aPi1MYbq6uyzJrGVpRUxKuXKiqi98MH
tLXV6BPKCwgyhcXYs7pQQLF06KFLrmG0Ukf/9vaZMPvUpqskKULcJ3w0uZvK48cS
MeaCvfXiOYXggKDJBWQwOJR8Gn5byWwOgLKS2yWtsCHxr7pkG6/7t9B9+q8fYmIy
VtWfQaAS15aoVeTWEzdXSl+uYnzfEOYG0tpLVU1nq0oW+q4XK4zRoC5hX72YHFbd
4PfPDCYgBJBveIM/oXlf2owUc2WoACxLaanj3WSF1W2nhcQiOFfXhTWjZWY/Cq06
bgqN/Ykxrx6HyCTD7rZSTso0pactZjfDuyYiw6BZddR+XDVbxavGlY4ax3y6VvuL
jZcvyiXVPBMWYNgran8ABJ+ljaGaNdEtGS0aUVbVWWEC5Qg72EZ4QuLY3eXh8GgK
c0DsEMj/6tFXwGmgKxwswM09c7k2h+Q6vCYThg5d7yT56E7LNx1xmi2bHcY+ky40
SGcX/23K+ECl1f9QsCIbPGvepVMu+c1chZ8YxN8J4QDaLgKE18HgBCn8gAFyTvJL
8j16LEOS406beh4dPb5RuyosLjYO8T5PFW6l3HViZ7OXUbVjNlH9zLe3BBsOLnwJ
MXIMvWQkVVj/Ay6qweYDqbkWcwHS98/gu5iLokIvMhU4j9AamXEWVk7jNF8/Yn9/
3Gp1SAjyI4c0dO6zVGpVPrUcTqwN0lkQkEfFlaE8A8q9P7jJS6wnUZYPtdyqa6v/
BxeA/wpcHPVyzqoz80+ys/PPjYVRnyWo0eBkI/ILszx0k5L86YciTRuN48t3/Tl5
SMZMvWkYd8ByKW2zEr63KzSqgOkNiFvGDwbeRtxuzgfpyP2plabLxaZjtuTv9rUz
gkp9sJsVW1b88mb+y99BLrJ4ctegnrKUmgSFX62XP1xorAdQ7ntKJqbDg7U0vr+E
ibsIJhPbMuxjDWqFY31OaiD3Pf1JlpFdZq9V9epYcLX6LIzZUElBYvJVQHdfZi+c
cF/Uo8tJ+es5ova64byKkd/1b2PO5Ia2Ye09mAEG1vH8x/8ywQRzE5FTuUJ0iHx3
RQMcoqUk+JO5wpHrDnxmn48/p/L6blp37lQh93dRdWP6aqOBPdAkwMkgOqTbgn3e
gD18j45AgbiFBa7tDo4hb7GZkgSIa39lW6bfPB8RhgUxj+39hfv3Kl+syjWGZRw6
pQ9wEZYdElP7Y+QiWatRtgK+YSKaTlWWvnOWqWZgg/p+uWHip2lfATV/zRhjHGlM
mS+Ni7uWYdq9LWYHjBXo2ShMwmZ5/m9iQjQOhn7ocEqLmA7889MTqMUdzwyeD0xo
laeL1sfb2EKz8n02vAR/BJ3jI5bHXFZrcSB+8/46aXRlQDLDCzxoUsLL1uvGkeuC
v1nDTnlrovgLGvi9t2q4x6tW6q2sx5WNDwzskdmMy/Opw5LMaJARWeYsPpePi+ku
4ylgMMt4ZjNPtvR6or8YBjJSOf/lugdGEGBkwSOJbwM87YLxRoI0BbszuHbVc3Oq
YEj9bCmXkPUf8WD8k92mnriRp00AYOzvCUoehQetIAe/ddWFwvGs+g6FrcOtnMoB
i+6nUyTOB5glZbsMMmRYm4soi5tw7ni34V8sW6AArhmwjkq6YhSqpIbDb71gYFBR
Op9OiuifGPd5Ubh4BFL6xDxXh47kxsXsC/NFwu2lJQ6ubGAwBnfVpkUfjS0OgyCO
JlwYBOZqvbDNqXP4jHS85bpm7ACXDLVfs0Jw4Brj1vy8o6um+A7MsqCN8MqepgRc
eoZTHkeD+9+jssLMEkPGOJQg4GQrY7wdRJpfpvVklv0yHlJkcWEaEns5pCeHvUY1
8M8HUmthbomxKZUl3MT+8X6LS5GDZK1gP9+jtCyF3Ul9zHvh2uTbTYGuCCwuXPrT
T1ufPcCZQpsfmC41mLXygAL2qgNtlPfNezgE/GjObVu3ZzAnSA6F2vZOU/fQpnq/
AoUa9oMblUNn0FHNES5bs4xN/dFyD33Ec1BSfM3TkNp5MW9z5raJpvUsarKsYLoy
7rMSpKMvO+WcDCmYkNPmMdNd4QqRH3GYjLX1tb0pFzbKtWFiQfXwOv2N4d+9+I9V
J7Wi59kmAVy+ZKDlwDYXQ+A2KzUy0kYToepkmTkpln/+SI19PJbhf+ZfNyxqyvVg
NaZjhfT8PAGRvuml4JgF4+xFjQ1S57n+56IkkqypPeuFU0Myno0ZHRlMtFk9BaPj
fGJyHLDoz7adK6xJ/LCudyj683Z63hjd0h3dl1d+JPFg4NZDDnhVlHmCD9Z7o7i9
qaN3Q6IWkSE8QTFNo3yoISQ7brzNXEPnBaKgD4xeyYH2Bn+UXVgFvP2a/ohrjS9Z
EaGKbefP7R6+Oza43TkfkUubbXV5q5pOEjN8SDS7dqTEo5DsD8+PBCujM/q9Dzf7
nvH7iDEjjn5SaTwcflw+xO9QUqa1vmMLBHxC/oSY3Qd4PWYrhS/C/VctysfRQnXh
k8nclonL35l/ToXIzC7TqX+UXfaZ4za/Jb/gAaUYp105lWlVvpi1kvqXoti2QuDt
BG8XvlP3o/81u9CJWSvWBRZsCPWXBbS4NDrs5gTVJSC38A/6G7d34k7xPxIychIc
QKluOYje5qcaBGXgSvba0AsABJ6MezOeHCVLWe51bPha6DhS16Bzsc0mkCHZ0bBd
j2Scfg4vv3kmo83YfTVB4RM53HXhw64ubuu7YCJc4sHF0Z1IEb00gV0S6PTYPVCi
xAWw6Z1GQ6oszqEoOE7tKS8bwBXI1plywSlizcqJjbgjfHYy+Inkjwnmfy8hM/oX
/IgOwPpw5d5C19ILMrefUsWtaX7NcUQQL9ZsltgBQ400huTiNUF+cCpPfq1XiRef
QsnOTp131pUPtWOKcyBOn0DYc84ykZwKRxLhPVwzhffjW4HIDgWkiKGzREeGrk1Q
cFOfgXNB+Y0+1hF3UpUOU7w+cPrGhDahUzIQy7GgHCO0LXvkTHaBbag1uJmMlZU1
JE32Ih1rmSrfeVLlc6BNETjgmfFhrAM4EsOK8ynsccnG3WXta2TJ8h42CIOxwSbq
ltqBVSQxbh6GGdIjvgXpq+fS9cNr2Eab+hgCs54BlgMoM3huOOUJ5YfBV8EndZkY
IIy4lC/uLCM/fEWzJz4py6Cwe4/xZHIXXRoB63t8n7rL2WIv0d8b+kFOmTfjg/6D
D9BxYLT87ArEtBsbyF68FzN1fEOAs2yvpgX+IZiZzi1O8I5IxQURdS0UKZebsLvZ
qZXywVMmCIYV605/zRtenfeRO/Ha68KmJ0dvtWPTXL7Bal78+ZPnAARVQRpQhgoD
jEHwXQxicGxqWIpEkeXmz1ZQ9ROQhYO9Maq7drMnRO1cVW+82uaPR/IjmgOaEPnX
/22JhZsd19NEJtAazA3BtukKkoNpqh4OsC9bxDLCI5hCPtH1bZDkSVvcbC5BAbja
LLEMjFIN+GuBkYhsNhG74phrsAFmj2n0RvPva6z4UEwbU4HsWiLkUtwoHBKXIW4g
pmtVyFfvN+XfRWWaMG27KvBNblBjs2hKpcV83BF539rIQCxxdRfkmSJOQT3qdYWp
ISLIw5mMZ72YbmtsYJ+tZcv0KySUXHOO8Ei5lWALcJcr4ZK+/kx20IjY9EcXs5qd
U3hBqsmpXH69IQ95fuYEvPWWIwaBcy0nNNwD3XirJnwclT8meD83Ps1Ayj90ZyMy
NAEKzzqj5U3Os5iVAKgHWo3JvIAWqnlrP031D3ue+apBb7zsBvMraTePRbLDfMuv
TkHjyhX8da7+8on+aZ/OsW+SK7hBAmHwSdO5qRyItH2+q+YlqEif/TnSJbk7vPkg
cSbfskenBCmwOCDbFpZ5/hiKeN3VWHmz1BBX5gDFXnyUt8RlBkylm8Be9LTXTeml
ANAaQD0SMccKe8kEtX8E5PEVS5HTFoCSWH0rLldc51E=
`protect END_PROTECTED
