`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z3HN/J3Lu0ArIYIBkirwoCo0pgM2etiNfDvWX8sLQdyssTwxK9yMeI4p0vOpcM+w
dNeF42TOWFcqkhJLACHZFOS94HMNaWn1MOmfpf5eMl194KHoo5tXUtuVYsBV3uIR
ImpJOmTWZHP9c+lahS7BFqqRiKfJ30wUZU6sebuVIUhaX4+g9u4pgBczQp7l5gUJ
5w3tQh70MUQ12ZlekyQ933dv+lqZJeLoJldRdea9CQLnJc4Jh5MEuDmTJrhh5rwr
wOMmHA7wDS8TuGMYaVNIWuE6IFHWXuAv3KfeKh9M3RcKJHtcKG/3hhV+q7PbvBQS
YWANn+eB2I8a5/xFqgcaneg8h75ezhkDXDpok9nuMzjBA+mtcPmKoCi2rNkI0OSe
PAnCLaPVm7mTC8AN6853Sm21p6dBuuEHlZiVwETLEIdco6M8yff8hd87BCiqmYfr
zrI2/u8iNQ8BjpcjImiK8HiujsMpKUcd+HM4ZWvQ3JDiwSel8nVq0oGddtYS7Rp4
JUD9wseC2j4AH8vypcPXaGWemoLmfDt9E7pqBmKPDE6dZJV8YgfoolQSHQDMYhiR
cBuuBEVjaMJNPcTXjOX+ZYyNL2WYpOErysPti7T8IAS6CFYLr06AjouknYDUIfCo
cSR3qM5Sw+AsTI0sV43f5xT8gBGlw49VLoraDtaGFtrBB/oDIippSQ0Sd8jO8ILt
bMg4rE9KtqyBUjJuJtL2cbuzF0woaJx27JzxFXzSXrYJ1VV+VaoDB/a1m0nPy/DD
bUREfbd81UzKJmK5esU7rsheck7bkJM4Ld7o0GQQTsUtzfHcSeCu33ob6xRbCTaG
vioAThc0A2UCBgz88O94k5WYH1/yuTONrEha/FOiEiNFmVHosIskQNMyhCeVtAWM
EVlUPVJouFyBW2zmm1itS1iw0+FUtFoyZctRbbHlRo9XbzAGN+oXNX2CBUy/HVwI
ljz7Ai3hI9TQa4ZQlOJ3v/cdgKp3QA3ZZUBraFc7cxOWSEFgUoR5H11EIdIiTa+G
BUhVjfj742Aj0iLJxO8ZyjTNdr+Cx6xKZ4GWa63YRjNYtyiB63U5ZsM6Qij4gfa8
BnLmpcqXQSpsrCWu1SvpD/6v2wZrokHabKFzAbd159GpcC7Dsfk/4rbfZU6Oxokc
LsM4ujVh1+PL0xuAqUvd6zXZywgoV5AuOMe4cQuWJwM=
`protect END_PROTECTED
