`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oVNiFJSikP7olgonVUkAF03q9y/yPBGGoHuy89FCsRVa3kCIawlFbyPrZt5IEkA9
XsaGGVHjjrOdWSUFw7OkqzB62hDP3hlPyQW4mnS+3hDmTA/oJAaV137GGPgxjFvj
fOz5f7tKglSCrrJVkjwp1/ulVNRUqm9TCma2BkHzsAKRUMY6sieOwYzJGMqfv1qP
i0+mdKze784bixUbfuyf+uMYFs4eBZiN8WEN0pFS9JOToe5bElgsL4w3FjTV9ANp
jzo94KCZLnEVB75wvWHkDTCKu9HuXfZQ0fHW1z82tqpL85CBPH0+oN/7oF73OsZY
11THchLhAM6YvyyozGhqe0kvujOnUy7krGKW5JIaFJ84kyLeoUsv27z7EmjZrl4B
W9Whc5d5VAvTw0eG/AaC9OSdcJje1tfgNo/wsTLhpBySkWAXRKEDS47rlEwonzos
Nla7ee3oF27KzXmGShMre/5sk8X2hDdYGO1XTHP5UPp8jkqGdZcg04hMrZFpzC1a
ARzoo5EPRANBPHvUCS588cUbisSXf4fGnNwjUyXh9MtiT1dcQCzaA9ysWfQqJ0q2
Gyh2Eg+gh7/wPRCSBEE45o64VocYJ3N70Yj3FiPc2XjjMcS4/wKQxrFPlP2wYCTM
`protect END_PROTECTED
