`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EkWZawGYnv3xs3LlmITOxYAitC1Z70dgesKmSxOVDDb9RLqjtPKlXyrnkP5XnCs/
z4hgvs1bqwlKHGAEIVg+ng67t+AITl1hhDSkhG+j8VZt8wJZq5TTYKMt/AuGpPah
Pp3u33LTLYojOUGy2gwauAXSqU+98twU/KTBN+1M8DUCtZnhdiDyoF4XUW07/nIc
Bfb9oafXE/k13t4e23q6VccLTWDa1dWxWpYqJvdoHAuOoEm/kkxh2o9rh0W+gbzq
Ot2lxxYVgxvl7v6dfGw3SbjkiGsklNBLF63Ua9/jqla1tnFI5TEheFvh09XxO9UL
OV6Sfwk9XCfJ8eYywhmJ5X4gboF1vwkFGFADKB/AgNc+HOD5POfRZBpABVvgpy/N
aIOja/2+kU0HqXNk8PlWAwvdi2yKTzmTmoHCNnRr+ptdC9jhBNZh9nTPsRjbEcJE
QD+ZMdyKeyd/0TlPkHKsTzyzmQHmJ4m5eyG/faCjEgWYqxqjnZjV6su4XAWB176G
by2fczRki6VVy7wlnJ7cbvRFK9hOY/b2nNJhF33GpAbo5kOBKS0JRaRoO41HmPYB
nAbqCh1C2rJGUrA9DBN0C7jNfjJraOvLl/HckqJX6jVBpTMk96ZqPC8h5N+NrDLJ
/JECUOk4Izlq7IMlA1KWIg==
`protect END_PROTECTED
