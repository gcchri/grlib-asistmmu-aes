`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xjO+bx8CuolndfRcFwByNY/fIj1AtftqtBaW3oYM8jBrJa1lIo3R/rer4jrZb6FO
zKM7GjzSk+arVoO2GdRyq/Y6fVNPgGuLhMXtiRZrxCeW1RjzjaZHJH3vfnzGI8H8
FejuJ69bY3He0JilxPUwPY3M2lu13YqIzpy+pzH3Zxc+/ayY2/lH4sTukOivqyZz
bcxB5DVlHJtiGsxGcSRYzrQPPAPISZfekB/6pCIaA+FIaNQXfo3ya34GdPjDSAYG
oNCkxWgEXCCtMVbyySEmz0OQ0fmb2PP7JfisXsp38mVYCTlaHbaBdg4hMnl6i7Ji
6roNotKsxZY87QEbI9ogPuSCFl8F7RxA/dUtrMv4+dKI8nowcOvuFV4I8K/nLIWk
rdbUS88PkSqrdZe8azjOdNXNX1XlQJJBtAFjHZeO1yL6hBefp+vTaD8THr+mlz51
hg4Qexcza4GglbHoGS0DgBrmJBwdBFU7FQe4TD5jiSl9h2kQNIE2LIBJ3u6ZhDp4
ddbT8Qd3ZJmUJs4RpRIPF1DUO1gvbMYEN+HwpikqSRgZzLS3pe5Mu7zPsDFsHmrG
S7B09bDRzcCUGlmjpXThbX80J2LyXr7wVyOmrBKtVwtTm22sYq0i1n5jHGnyyKYF
xF+ZGpaSmR/NdNIGzGzViw==
`protect END_PROTECTED
