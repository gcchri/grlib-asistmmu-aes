`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h2OgKS0Fz1IL2eMRU8R4G/I0yP79N/oUc+kKR2GxnRwWlz4/bx/NoM8At6lm5D45
0XYw1lx6dTUsxGdsa7cZtlpDaDaoEXvMsl4hANzdk4BZWHP/I38/drOim5OAXj9O
jmB7l7lYyygZzYqssJt4wVsz8UVVmhfKIDlezoQsPke0wWQDuMKXFCod/UwEwpMV
KfFXGyqf1LZoGatuZ3/Rbc8oUlWmxOofPwDJrdKD/BjKSP8yDsjAtiQReZAR/vpD
8+ybD9plecIcfAN8yNQJn0p8WTmyyTapLR8Oz4Fd5o3byNYWHcFpoQjDehmML/C6
fecm34aFHZHjHYsP5Vd2uclJQYrhpjeNwsvwwj0S3/FzNKxd4fhkeuVcfCJF0tD+
ELHrTeC9CejL2EN0Du+Tlxb7lR6nV+gQAePgQUGBKnuHCZj1ixqDtgMmgKAEesdY
qMT/5Jl2lJVtYl6V7f65yUZk3CE1PfVtGWXaJj8tQxaiFAQUkpuDhZMv5F+eJqk2
U9D2I9odnGI8R0qA3H2pRr/LOxCY5+b6TjMQmttv6LUvEd9D+3dLTKWHcpW3iAuc
3ftyw+lXBtr1D/Nogg9Nr3sI7fQ0jFCaHcHBUsAvwZUkBgiQSCQ6fa9J1r33r/dN
Y3Jt8g1T9oTQcqImZwGcipCjyApnwV94c6/1IXAhvHA6TQr8rHX8TNPE9Cn3XtgR
iR131TUusklm7VNxGfpVVYKpNjOWx9NsaXAqBWTnGfSKQGoKqu1GNZ3DymOizkw3
gAIdyGa8wic3S1z2Bomxgq1jrFxdV9darMIfiA2hhq2PV6GTbaDrb73LGCbulXMT
GsACVKvYBfOGbjyb3I2fFudoylgg1tmCwwVnG3yXf3WfRv26qfCHmMebLOItEkDl
JhXTcV2+OsRqKXoKCigbmWAreMfbdBGe6d/eF1p6bMrL6CWGTeUQAp8/LGWuiiPY
yqu/AWl5jkVgA84res0lSEWLAF9Sjpz8vWzsQ1ocj47UKiCrgYbChhJlmC5EcefM
9f21TCeHurUja5TBLgCxCm8ZuYgEhv9fmizBGY2BtTsS3cBJpIvcL6fSUoRokhmh
cgJFCR8l3fIU6wcFH9Agx+vICGM7GeYU4WfQ5dfRfp45bDQtQ3XiET/4o9u+evl9
qyGmi1J4q7I62vNVkD4GiTo3a2X5vNbTAwkl7ZbjRQmlDu+KQNPO/0lTp1O8W+3p
9OdGjHMabeDmpytZNfoBafADkY52OSgWG61USwFQDs3ZkWGliFt9x28z8xcO8TXE
8VcEn05mrtGMqYghSGEF0VJqD7jdbhODN38wAgCezO933y400t1BA3MQFlwd/17m
`protect END_PROTECTED
