`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o9FZZtOytjoIURJe5pNFe3m5NS8xMv+OZS2LAF9cvLETt5Vp7NbhHGnTDwnZmLxr
yMxJJh70jhypkfmK0ez2fGncIa1eB900PdyNmLg0as8awGy7L/+FlkrN8zJEbsFy
Fnj0iCRmFViqDFfv06uuhuq7C4OXybWNbe+xQVBT3ztZgAX8v6kVXvA9pRS7NZSS
igHopVrDukAJfMcF9255Ij9e9HxJ4C7UV0l0CBhE9Hhs4yw4X2XtM+Epm1ATN9yi
c6Sz2mjciKx0iMY3saFpVUA9uhF0G0yxnYYfvWkNDO2xvLBrdB5pm+zwErzmYrFB
6326O1T4QDkQ+ou7DPUCcyrXtPlaWgSxfH3AsJfG7wNIEpkMKf8PmghzLwbXMEC1
SRRSwh1YwUn1VQh3eTWBvg==
`protect END_PROTECTED
