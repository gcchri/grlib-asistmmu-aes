`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fj8R4Y7tFqIaY2PPlbNLYIPtNQWZWQxoZ8klhSnirJThpwZ8HfE3mfY6In/+nb3v
9cMlZZjef6DVmf+Tmtm3+4quFg5GAlyON1seFX2D6XFSyo72sWydl8wBzEo2qI1N
06JAkkGNokuAgn1UCdo4rpbPz/ETF1pKgTB1FWRrz4MFzu+XPjd6mGBBXrnmawh5
48DDPNZJMWMnSuTe1UxtwX9MUchbqN9nRUGBIlJK2AAeGZbuWghTxtc+43upGt4w
GEHtcI6s9mQi6AHXCSfbixP6b3npRXKWl8OukCpBZ69Jvfa3xzeXJnRAPtikrSdz
v5Upx+6oAeixFqxkdX/AHJKxGWhI3J3RBjwYAtdjKI1RP4f9U00pEmEtF0xzDeJE
mfXXz0doIMlh/SHwvKuyQM+5RFurT5l8qZ3k0uhzHzuLNKckLxTp+iQCvleNzZwJ
tqnY/D4zCXb8qwbV1cF5h0a5WPlZ9Y0wIbMscyp3PgnY9qN7F69iA/emgcuyXfoi
Wu2I1pZZ7FAORqEEba3MKk0iRlAGTWFFsbjFFdvVmzgSp76pzgX4JG/2lk4fQXnu
8jlEgn4zUh6Jj66FXevYw1Y8RSgvi+HXe1SIYtEBhBLYu17tS4OPPIqdd3Ik1XxU
jggeiWoD9rPskaKTfVY0ZhtFd/rCSJc1esq9s/xCToz9HqRe2kHq6lIFr5SWo6rx
ftntRV+n3fg7YD/y+cleQIgTT04Q/hwPUPgVKKWUY09EWduFRro/rTX19NPTVtCc
V/27m0Mtc8TJk5TPnm57ugDY0mpsnweB1qTyXH3F+aE3mareELyD0lhFpyTh3VI1
STGc5xZhgYE6KLq54E8dY2hX0AID2Xf5n9xBpZWhqE/YYbMLUg8K82Qu5fZRI20P
VIqMZip0RPI8JaKQ0g6wgzPNLjc6ED37VY37qCuwaCcs0+lb0D6E9UI24H/MDQee
mzl/9/HkiW8GTFMMi3UF8Gl/Phh+uuqQJcwcG4tmLjQ0vg3GyTQZs6Riu3XKlP6Z
7swIS7CP64X9Ayyahd7VOLaA0wcj+4G14SxGrL5MUJbSzyLZSA2hSB5uKU+jGQHY
e19JZNDfJyCozT+DkedsH2jtnx7JPJSARNp7r6CRWTqeuPw+95D6iHdtYckQK4lD
+K5gJj07yXTWetNjXBmt5IH3Swl/tCHHphl7ys7++EPe1czpzoQ5+iCFdvh0Kws6
Y89Ro0MD/zrB50KKsVVRxMUdYRtHie3gTapAsOeQtJq4KJ70aVc1kKJ/3JdFMsth
a+il32JEYY4KANf9x7BWRQvlM/G/P75Kfw5ptVDzGCxG6TCZDueEbgZdeHtzpg1V
fLB0FfzJ31P73WOA1axLbEegPFr6bG10KeMJWY+GAid4HeXFvRfP3lpnC7X1yD3r
HsXcRsZ5oO4ZcxScNFoiI6DRgSrY4Pe6qtGHSWizT9a/JPqEWQB/6J35kV/5SkhQ
CRhrnrWDUBs6wLV93LfCll83G5kZD4uJzyH/KIdLs6Q1Pjz03NDuCCDcJhdufBBE
EP+F2S3W4yDnu1j/uIZ+3mkKoE6sZZVDHWR6OcLrqMqHRDwnCHTOT0Rzh13BCOyB
0qX1byLTaMh+PJYOx35/V/dwFxGidMWzxYm8vz1UlPQYwGf94VgQVz53yFfi00Dr
pELdjByPN5Qs4ieUtGtCmwEehg4poOZddNEwzc5Q7BHo4TPb+m3EfoekRv5TQDR1
9orFfPVNmgy3kRTnVWSSmmZdY/BGU9xR0AnL043jUw0HWg7QTbgG/ghGV+3yLi2a
d7PHZPF62vNLettYV1uQ1v5RmV+8YUlM4fWLCSsxUWUqXLQo0oLfu+7HbU1IoIiO
bZ4ToJm5+Oe8YnoAvv6e5N6vSc8j7A6LOr455OElKnIEbkkhMOKp3BHIZQAcii7l
UwkiBMuyYXVwgsUE/LIcQPFgbjmJNBDWMrsQH1btz+b8CsWFEXscr5lpxny1nX4g
NqOtvCOMs9OlZERSNQ0M4OzMynCEHtE9YACt3bnwFuPaVLKsLA4fzaSKSmo7lII9
0o0J8+Ps57pmsXqCSAZgK6R985vFeYcUJLn8VXo/+qYsq6mek7ZjYgOk9x6a9otW
WDz90Heu+Sa8PdGo25NLDXkSHEh5FBK0y+co5saYA52+0MRwr1ELw0sNd90od8rF
HVTN84JhRH0nwNxAdjJ1NNn4IQm2A60bM9W1lbB45OHANF1hUVK1WI1kXbsduwOm
uZy9bZybaV80k49nIYG2HuD08diRflGBqnZEXi/H/cyqO2s51RCTuh/v2YEXlriH
Bg5sadMGiT9knDLHeuFkQo3Jnz2WV9yjt8pINT4DR9u3cQoA62yYTvah4alcu0oZ
mrWJWDVYFm7K2Kb+Jzm1p4HfbW6cxnYcwFfE9zjeF+z2YiSWV6085vXyHvPI1R2p
ht1xqNHmGonnlLpo2UgScNzJLyIeRTag7vITwNZkESS9mWblrXo5rO5+FiIOsRUW
rksRR3HZ4jbBx1DezQku/i/RoQSZ2Y9jWJmC4FOH1cPL3FFFzFnH4Z7lw5vMtful
oRO2B+gGkPzzENHWd3Jq8MDY1EYu08VwZecnRuQUhXRgeSdHtGrwLLnTKmKJ2yvn
bT+N8hbqDbkvwa/LNZ9Bj0M86jbV2lYc+ojbt4c3Rho7IWF6hNA55LCr2rysBULe
sM65sJsqUZBx2tymkZHw7cNBzDpD24IkrL98VkvbNsU2RhBOcxmYjWM6gJFrTXtM
rXMOQTZ3WAkwj8vLj9KHp1A2MoPzden5NuXSqcAqWJZ4hZDR+N4ipGxaWxgOkCoq
h/ynAZg++7qWoXnQJ2u2s16opfgbFaMNDWgcwQqznuOUqA5ylA6Tb6SvDwsWlsXs
UMXv/jHzt5CD1I+u2yW1xSyo75T2TRtjnj+Ha+g1VP+UXJTr+J1an4V87uV22NWN
GASPEN++HHx++l6aIzE3ZZle32LHq7VkMYf/0rGq7S9fI/WJ1lDI61xMlkutHYKr
6hnVUpT3OKFhQfIorNBgazWtcWJa6lJHJ1pEGEbjADtX7qNGefpfvpey/Pdh8pAk
X4tCwXiI7f+INdNsT7us9ksK9ZyS/bNWGFPBBoJ10tQpORqR3nlihInTL0ObYOnx
OWXIvI+gOu7O2uFLB1qOoVzV5RKs6AObPmIWXkutJ/EQ+hXp9a6EKIs8RTtQSUPW
DsKd9ay8aSCAOzTQ+kBAOxCA9vK7a1qqS0qidoUV/8oIFIQ1tVX9nJz1JNxNx4Kr
0q5PB+gWA6TkrpQynuQcYl0dbn4rRa7pwPm2w/CA9Oipw3Gc3PuupXWM2PwU6Gds
W1gnaCiTEY3DbJJB3Z7BHannmHP/EBDaMQ/ZnTxA19vqVoNUdrlMChxjilkQiJf3
RjOnGq1gAKOLOgUnVJcWuZLgf4l1JmW9oUWQaOZQ01Fq8dVMfoGSsxCFpf4TldjE
KhCM9uZzx866x1Gc/VRNAy54urCmLC/D2rjWLVOgRwXzJm1S/4LEqaYoUoxEZKO+
dTn94Qch11x8LJHhgxHX/xTSJkb/NT08lU82iqbGzhEYFOkFMw2gy7sb5HO+wCS2
pZ8lNVJuRVQLoT3WZoU9JClEfg/uxGO9WwFr8n3YPH+eB9jDq63WMWwMCmnqHY31
jCu41GOQAoQ5IiHvPKtemvku2b+iOiwAVYPAVknQqAfDvT0b135i3FjIUS2oiDud
wS8cQay9M0ygskps7rHqw0FXDfDQsC4tgLmX5GSNxNwsk1pSUdCmumZgcYp/RP6q
PK3TbnTlKNjXajUCiYdN/bPzLhpf5VArnLcMF4DDJTxEUzoRGCSz94Ch6dkvlB7C
RBKOMG9pC4QVcUgZJEQGK1Ggy7pkTujNGCNoDR+bEA1eh/xQmsmID+9TH+nDnwcZ
JTvdTw0quUNXKJPQmi3ycxjH8AB1D6k/7vK2UjGm+nOx6WPGC4l7ynU+GXKE4mS6
Qb675tedo1TWm73LK9tugyTA2Zp104AlHGxU7Wk5+yYIlBlKf/KJrFUyWHyQj66P
J1g8npRuhqxwY5Qfva4rfe5bvKQrkf6weWPh2uz80mWN3I3VxtN03d8P6D/4dKjE
IrwQxpiEgbmOqj+2WpqDybK6nvaUmdqI9xrYUOa+KNAQp5i+T9Znno7IsuK0HUfk
GYpJM31kA7hmeJaaOaaOQwTpiqm7IuhgxGztzp83PSzfI8QwVHBOAY1LcFhE9EUW
FboA61EQO1bbkqeHZjMQf0sUW/8++SA2K4Vsiq81APK03dN7Kt/F9Yksvp+RK6s4
NwNLGBMyZpt6bnO5BeU845t+z8U/+fMP3TESfY8endGcZkqwVHjEJeSTHL+hK7Ux
EWoqt0Jhef72KpP8OI/DIo36uqt3Qf3PVgIGY4+rN9nH5qTd9XqrDcX4I+1ie4od
CPOcPji04/QQVR0qdiwip7g4BI6oSc+p3KC+ghAH8Pf9FMf949zMMImM+CZA/t8I
r8RHsXdEFeVUkD2+qhm31c/B5f6kHuxZ8A0kPut0x5YPgTAj+cBK15UHM3Ih/uZ9
uqzY212HQV6EgO9XH8GL4iK1rKuCmjY1YvvxksUeNyxRsvd8J6UCTP2ftow/oqz/
SEWb23jLAeOWrh+G2oXwXPscwTKyeRgjkkiJLdLJE0ssAiiuHmf57ZTy3BL1bvCr
nPzu+KisWm4U5CNnz1htg3cpeJHR64MaJ2rJUS9vxVJsSDYlh5ULF9HKFTAi7sfm
Aiw+I0nmyYqsvlUO9696/T9U0A0r6LjnCPq55wlri7b1iAil4fizc/MW47yLA/j9
kzKqb23ltnV4e81ITczpmj4LajWbVWQVfHbhu5gYErw+bnfpfNN4KDBdgdu1M1Aw
7zEtnMCPA/7l+nanqK+SspGXFcrsuS80ryv+yG1vftSezL/liqQ8ZlWgQt6iiVS5
PHSlGULJp6VpclWqHd8Uo+zwCZYL/RZNHzREMEL2OoodMMMRQ+xY2P1Py/XyHJEj
TJO+G3w/93/o9UB6pmYLfJXbYzZnYccpWTNkXB8ne2+1SdbdKj2jGv0MbE2HbeXZ
3lvLoYoT4hTt6souZ2MElXXsRB/MuKV4FKTnyx1M0sj6CRH4eBBxEWBtwjyzbUZe
LnpxIStRdOgShgS1eHsnCgOzNAiPI2J0LFrOcjO9sgOJpRkfo67a1bleqk5sG4Ao
av1+BPmjRkt11qMdA9JRfTDPHWV/MWI0YdObLgVINS0u7Ns8ocgvRjJ42q75j1cf
TdIRmBHi0pIaVESki2NibuwrK1wEOKruqmkX/VjZaKoiuDAE/kJuGgGAzL+Cwjl0
wyNOWGBI1IOJkCGnrUGLBV2AC3VZdEx4PoSFOWZHLwnGXvIclHba6qlhFrTerCAe
Y80+ZbpuSemekwLYQMkb/HzPoP/+GyaHtJqL0Ywx3C49ID/C3dwk9yDO3Rwnyv3T
24ZqvP7C0jvmIQ6F+LkRy0JEE3hwPgh9mTql7OYjmhU0tt6Q0VDF8u20NAp5ycx/
LsZEkFiaNBiBOnCEE59sg5nu1d5ngCWEVHozHWuBE266xKsq1mqRS2FYJLr221PT
aA79NXZyhl0mnJH8dES2VqvNG9bFfOo+9FanmWSWWsBIruCy4rQLdXU4jpwxZECP
/iVrZwixgPaqnag551OvIj5vseCrPC2VDqXwekGA+H3SrV2DzdyHAal9MVtLZS9q
bNPX5yFN+mTtdD0+uzzfwCUric7FP7w1rV6yVmsdz5gyWT30eh0f19iIh/eVzdBe
yaDZUVuBE5gPDj7R80U2QeHTCoAEisVdu3+BSST3e/58dBvKsXqNvqfFDxZWw3Qs
+MgRvb46dKk1UwSnEeqa5+oirT9ZWcFzECKVOAysYL/JLklCjrpOXIoC3iDxBDJ7
6+OPHORakLIOTGx4huHNthnJqXv+ZfxFwyhI+wPtVh9sZTi6ttW0SiQW/W4DIvnV
VnChl9F9pxPBNa8E/9WEJcmyf/7o9V2R410Z0tvlEFQHjdlljz3umqsWXIbF8xiY
sNfE0k2mlcm+SUUhv0Tf/0d75aKuyWdIMRM6mnwfP5czQBV4PBksQ2wVsRl/cL03
WZfahlAnVStmuLDFEypumj0GaYIXoKRi08c8Ehc2rYPhRUU4STnd+n0yVsuehN85
YrMNekuoE/Zw/y+lH6/1OjdDQgL1TRUcAm0NqyaGIMcxoi3syfcBQ/qbKhj+fhUR
lZ5KvCOMLia4D7UEGUZLfO26Nhf/rvzg1RGnB3OF5zGm8X+vNbpxESMPBS4gpcWu
25b1LwpXqW0zzjzLjohACKmAhuTPcUMfLAFuypPg4B/MQKU08VXM6qUquuCFzYQX
9ah06yXe5gmyEtw8dznW6N9ANCmbT6Lu5fafnNrWLFbn2soChfO3n+hRhWALta5Y
+Mz1s/jIiCaQnFghfYdUwGmw5/EHTtcxm35qYYPVail4c7K1Zen0AzHeNKtn6vWP
CQz6hPFIvgAHWMMmtqSg0UWjdMf/7/BTpBMY8EZ6VPGp35qBRxbZQNLibqaeqbLq
QslhCW39zeq64lDgOJFM3dsrn9MCb5733cR5DCxrEkV3Ge1O3r/EaP4QkPw42cPD
MqQMkbG4HGxlZawA47WxaH+eqecj0AA1ZJ2j01BW0czRQfpMoxV/Z5Pp3CpDw1Xi
Rz0NGfqexxUJ3tH3gwj2CaTklJE4y/QY3WCngn2wa5eztp7gzlOov295sXbnRlZp
6JgHZr2u9SilTKweNROzu4g5PoYC4P0cw1JrfKfRSg4wa5lYBxcgGmgcY8nqXPoB
nR23MzEQARcErzOB9XgpTgKquT63Ssfhp+HtUf3BzzaWHUjNrdJySKLxbw/j4Dgs
ofyP7ym5UWFL4PqgJCKXPBBbeJP18YCXMLk++YE4O7nbsPMfZswcpnvCksDgXIFK
a1aGgd6hzsIZnvgJzUc8RAuwu9Q4AZ9ccQoe7qXYSTMP+fjX+HyCX6rc7bc0H8+e
wZMf6H9tDwWK8oqf9lv76gXmyC2YQFoZdChBqU9QaPqO53/VQ45idiQO4YIkZ+Ex
ilstq9iJBVA3iVgOR3fTxXGVk7/cnOb7O52Sh/L1MfYAi+NultAd1pIx6xX6TylL
PsnVUfRmpNFEwtzl/ttPWi4q7KrFuGOzZaNCRl0gcxEbLP9PzCVvJC0Nz5gARl6j
2NF0fAsPSkx9uc8A1BqLXsPZW9Y1nfQpJQcKZg0ojpD6B/CzbciOXM9Z8kPj1uSv
HUOvV1/rF7ucmugGRJIrUgCM07VRjwusjThW+NVRx3abwxzhMrd3HnMAf1BuZRNB
kNJuQYcSl/8hba9zcywqONP+43qAa5JDKxP9Y8GLpTUXx8HQbBABPgWHK+66T/PX
BxdkY+AdgtHKOCtEnVSixwjEFPeZL0hWTk30VvTkoU5ARHgwUwptIual89drSeUD
X+dAo5vPUkxej1dS/p1VqHHD8XTA/t2/n2oa0xlrKXAYaw/CQx4d21VHwg7C/2Bv
xvLYiJd1E/X9JjADjOnQ+oqjO68X0MZq0IYGELuKSnGD9T51l64sj3RX18E5rOBK
tvt85ocqK0mXv7Az2ocqy6QozepaqJpZ5EASYDu7mv46rfQWRoCrQn07FHIofL2z
kQpf12mLbwo/HD6ojIyGgXGjLwwyRAZ7EgoQnOw/YsYc+owVJ08J7yJuPgkEx9hr
r9BJUZyMFLvh/PI9EpjcfgVWCkstjURMAYfjyvycw+iHa+NiiCk+R9qEtklOONQM
4Hpv/mgXq5xIBfbGt2Me1gzPxivDkrgrrEj8QAxyKIdHMGyVtCt2RLeTVHw3WBRE
FNnVqEdpCcXzqsPULbpVrKngABVwhzwdeZHhcrfmOZ8k1cEI+N9yy3UIlbqnyEcv
oMJHW5uDWQIVZaOIO7YPO3ED7KnfyA7KLPE90VRy7cwfRFr2P1mj/F7iMvzqXlcM
1nBrYQ4/q9KjUCFR2jfm+/1AUAaI40Qb5bhGaP2lwKnQicMzviJObdcnepK9lrlJ
PVUzLEwcMdQY+d1DIJ3ArHmf/+q1BdvWPlKPt2Co03Tp/wduL3nzt+nX/L1FKYuw
/VGZ9iAyyEWLaAm420F4r4royetdEoyQquYrh9yTwG6wl1qHatliVnvuuTnJZYla
LDMT0+IMEzXYRP9cqD0AO3KgBX6kHP426IpoabY30+H93iPzFr7vYPkkYOud8MVm
mUKjrHGRHIGIDLv0vtumXrzOKU5t2SYxaGD2a4eytl17arwun5NsSaT/VWm18qqV
h7e4K8tkilCXJ0mu79hi3MC6rXJrMPy8sDVsAySIiWljcialvPMYwLsDrCEQOReG
14Dih7yftjb8SvHq1SQviW6ZUi3B6CfTsrrTrg/NXMdNEXThgsXTctPmf+UFp8NV
lJMwclcmLwNfQNHz4gWdqsVXYZguFg7OAZSfn7B2pymKsf3OnMyR3gYKjh9WkkUl
SLlZGxvgLbBpFp1zFEJ4HN5SePR2mNsiZQjv73NNJwvj56kubwkzNhVVPMkaBYu0
0Am5yFm5o7wyQGdl/3ARvxZRSIoE2aahVYiBxUAaNR3bZhP1YaZoidTCcAYhmh5w
GkjFUvZ6vEeyhbRF+HA6WqS0r80lZmCn+TzpEtNsG7EcR6o35yxqGHJDBJilr2EU
G7JaHe0/upAKPYwrEIJh6rop679W6hQE/8BH+8wipfSXdVKnhipngBkreNB6GIZG
KNHBjVCydMU+7zRcrfxXKGyun49Ub2bh6HbynjhKd+2q3dBOPzwypY2+KP9BfNFV
oFSIw3T9Dj1txfkynp5CjPIkZ3Hj7NGhJvD37qr2FdryMYx9ijDBTk/0Gc9rqkQ9
dfG+NaydLJ/DOuvoQUA2msLoldS6JUgqeK5vIZpO+Ypaz8569GIo2I1JsM21uKLZ
KvyQccXj5rLgxyXT7qzzz3W0H9LEgwuOnaJDFclx4IPq4udxLMCbRPPymo9zGr+4
rzeiwdzdzGRXsSS+umVSiuwoPRaU5DGa+bSan3niRkJ6omgFES1j+BBzBnLHE8xN
q61WnCeYfMAAzKfYKXNMleCsi88RkQWQIO0464Tqp92UD8S34XS62PwCUCJPPxYg
uvLAHBEtS7gvT9HIJe0Yt0xcIKLoVm7Mer6FoBH74u+rXyxDRVv4ie1rLWPItk+f
b5zaNGjyymQabz+A2lseo0x39jljze0M4N03OMtAAUEnoT8RJaszW63X0l+mAi62
OCIhXcEEi+kyE2BZ8lKCYGQ7QT2ZJwJCEKthK9YW0SPX4U5kpSq6S0+A8d4Slo4V
JX1T2MvR1H8GyHyxXmYPIXXxkrgyxSOVUYWau0Swu/DXCUDoNLbQ93aUoNEIKWMz
Av4gt02sI4FQrKwkULzsuQho/U8t7+R9bDnhA7tqOoc2MEyqZbwxHO74PJMESTqr
nYEOQTaHK3Iyg2YG0kvEXXNQA5bbjrCiBhk1d6bl4raTHEaM0Zlia1CGh6hsYdck
EvHij1CZDgzwBzGByBCHpzTEYgYLnO7JRs9rrW3hGccLVeJvxT8aZYOG6A7f9t+H
cx+cow7PnQeu7llO92y7R7lz3wihQ4ptuy+FvAEKrJv9tDfA/yixt2VnTOBAozkV
CD2OGRrx+0qRrhwBiJw10hleV7b+dxtq/GDHEdnOd0e+h5PUUVMRSr/vlnHu9rKi
yeSgN29qvhMlXE5sXvHuWZGzeN6j+8Wkc2setK2zKXyi+2cHy9aspRYG5Dl7qkD3
xh31bSAUaR9aCYV5Yr3Ph9ruWSjkBWyBesKMzdiVYnSbbLiJH10312il/ZvmeTg9
V4ubLPNht0I7VLIYtq6jGrJKtXZ9KIBhw51rjTNLzJtR2XEG3TmOJLRWSPfCa8PT
ytviZF/KVuWIGR5INoXa9wzC4hqz3XOgO/EWlYJEEeOSFgfZ1ND+ZmtIoE5PIrW8
TiykfutvdvnTm5HX7hXqdMwI5xfyTknT+VYyaUEKBZmoOtpgDyfZfhpyr7vU+jHJ
Oe6Dy1rM14ohbnL5bUj/qh9+f11UFLXSGk7kmKHPl+68UVynIrYZWZiBV/DYxEYt
IULXdz8wo22froCC4US18XkmI7wLdZZxxEtJFvex05p22cF1s20rIhp6bpOtSEou
mBp9J73CpUxyIpPRRFHn8O2keBZnM9aoJbUDa1HGV2xM6xiNP5HJyG6jp7oiN23H
Ebqa5GZwarRPHVb/e2CQe/iwePt3EcSUBeglXypiEIFX6k7FmrdjEqeagEg9sJQ7
aXxoE5z2iVLZZDdCOtQ57DrLiKzrq8ZRASW4s9RkTUZOLkgYIUzj0Lr4gAuTPIDO
0iEXlWnmY6JEVY+zPky8eTGvzj5TuvcChfjLkny8Y32ocKWszpERmyveehXdvch4
dNjiC6dx5+twH7/qOZ9wazTdjbOfhUdF9yUpts/Ho5vZ3EF3kIZZBLLZgI9D48I7
m94YLMApsu560s2kZJIvtwE2o1jjFe5s9XPZjVjPnaki5mw6ZNJm55Iidg/uY8G3
XvPPTxiKCKUc3KPyZ+BPBhX2/x43EyaxNgruR0HX9eeYWS9/+WyhthzszN7cetbd
zRU4JlK+4w9ZpwL8K3oS7lslbpJqgQwxq8tHpaG8twX8ZttwHv5NDjGUS35KdDfT
zDHK7sKppUbjGs8Ff/IzdfHeYnC/99QnpPw/amlA1A/oAlawWoLlLHlJ83mrZOMs
Ykclb4BDPSLx+h1ogU7XocNMvy1/ykFi6hvw6DW7t7DCiJZVljepFzxi4Fdud469
Dj6Ih3i/E/26udQMggWfYLV7VQ5B0A/GVaFCKGrGnvkyk5JU0/31BSqw/Vaf02Kl
PVP0dtqjVNkxDYNjZAGu3eA8od9YpB/lbzBykw3pqXlPDc3DMIZtNSWOWhJzewSn
M08TdyFKbCJDwWPXHjcGzdFx6D2HJflP1Sb5/IVgYzWsZ8jTk0cGTVtqsRoOGTe/
ToFt0xiVGpfEEiZX0J+Jzynwc0ZsTaeDn2GLbid4E94m3aQ8QrnKh4D2RIbk0yP7
E1AeGj1GAxQ/Y43tZPIUFBdwgj/4pxZBwoHMfQ5MnENiAsz9eikgjaY+a+WQgYfs
XxG76LwtEDZeoS4xYtmR2//6DCyVADmOngk/5MkSnqqAmzO3sYfCRIdK/MSNIIYF
lD8ej0aS0iaFvmLlnZtLhcaOA/kt/jc3VjnLuFEGybPcR/5BcobVZFbmcjmH2tBH
Va1Wm42Q5d89CrOAWVB2oToacJnY7RfQfpOzmZlR2CYzFmnvuF3JoT5fpwLdBQ/7
hSQC9gEAfuBvrwoAQiaAT0LGfgOAZOCAy0MgD2UlmGpaRbi4eYDNKdKfy6Y7AJm+
2ndIU6qu6Qbf3Flz5ZpaIsVOH07gn+yBBJy5cHFFv3Igooxoe4AUa0eAgOyaQN3b
98C9l+CSK9K8L4mDKwjnSdAmADyfjN0KC1OFKP37A94bAF+nvB+UWlOzFMejI3EA
EWS87a7YAUEcwnqp3FFdo5iiW08jeQ6UiEVfsxwlu5GrKu8LwF4HgX38ubHOjRXc
lG1322C9ieu6UF13q9r8NIT+0nUHA+ANS7VqifJOpliPzlKliRZDDy0usEjon47C
7N/sc76h3wpSvkO14KvzIeU8jiLdm/I4iZ0VBdqt+6PaOFTU4XVAgfPSlid7VfoU
nsggzrxJ1k4iKS2KS/o8rVMTVE14tt6UxkdGZqaX1kkLOBE0Ev6pCq0pDLAmOJff
5f6Kk+3e3cPLD4w+vFO5e6wDxXIS7ZAu1MUXtRuaoOEtp2YmO5sbxhP53DGUaTkB
98+F9qWgJ8TrLhr9TRmYLtTcL13RtD0VFiK3sSKyhSt/jrhFArQ1+laGsa2vLBF9
tSSV2gq1o1Nrd17u3EjEYPyz9t1NtkbrPep4SEilfCuXbNqq46iPSbElxg2fyCPB
aPl+ItDtg3/l34v4wpYUuUCz3JToJAMqmbrtqQIkTXz4K2QKp49C660p5cqsGvnd
JpXsR1NWE9DO28s8tFi7n/3nVFF8QEaeZImNbmPDJwaEpUtU6JKcNx6xYrNVW2zk
215hgbUVeIt22dOgEzpHZ2E4u0wfvs2eY0hU5FiOd0iCX0TthIYsO2Dnqq2NYjRu
EPfXvyIsbzf4AjPMrnEqtNZVL1JH61lbz3EiYfxd00jFpIMz3cqqG7I6TNDyv8PX
TvMQjIjWD1UsD15HUI78xfWtC+Xa6+Zx2UBtDLy5V6jDvQGQmfF21t3SSJUIF0O4
YXVvOLvNC+n2nXnJ2K0fLs5IuY5dhR0oK0N3D/ebFF3xIcCXXN2TLNPMq9rH4Lbs
sIgIAbgW0RjPFbzq2Dg5S3Oj7CI1v+KRosCRA6qNfCXkXUms4TugQpbvSZTEYOL7
AA6ioFQXq2POvoMhjK62rqAwU7ZvujqDxFjGzwpAHCHE0aURlbkdAtRPuqV8lNZk
79uRKWL0KAhUlVrp8kcePEbD0yqv5YgirgvbiRrXRkhBAwd8mPiojKbNc4Kq7B6+
rAaPeQJwqPm+CcT+aojXD+ICBsCko7QFYY6jQAE/ZZORW2CkRLDQfX7hnkbs1OLJ
irIpgdl9Jru3ZlHVb1sARJDCe0fUxeaNQW6fPggFbveVQiULRMPNTMZSQY+8Yq5O
eqrJGReAH5zYkYdeHjWltaHJSjYm4JTE5PdALmao7kAhI4PU6P7yU+FYfJX7kN7+
MJQ8TEczHXkgiVtBHZai2QQSKyFguDobWIYoB94c8kqBCv7E6/wNf7iRhhGKon50
5TFLcUB9FpzExJC1Uq6KUBnx8c/CmRExmRS/e8oNs2qTtRHX5wSoinl+cC4BcTOP
76i1jKHUG0nWWtpAMAqCcJ14zLXqa1ystGGAXm9UH+NH0O3ivwu5Tb8m8BWjIHY2
iLTC4FnbL8/CYqOPVkG4GQXaBL1QqWJoQvm9zdNfazOrh1U0ljW8FPy9hrs15KAh
j31rPV+52Dg8syi5OROa4bmQLwfgmnrmHoBGJAZjBZRprWMLNUyMt8TGlFsOwuW6
gpvF/EHCaHUeRv0cdCT7yaRiCjQVEMKOUX9za48kNjQPYKJwEWRC6U0Ko6G6Hf2l
p6GLFdgq+vwOH5c1Yhf3LRdwz3U9iMZryndFwKv6FyjoHQBZwXRnHWAb+8BkDkCJ
i78BZ79+mODbMU7/n2tQsK3OqjOHOS7WahZU1qXKZtx3Zt0iYiD79sdkiH17VgeL
1jZy1/W2DijxH9YfUtY2v+/WCK7oc48tmFZ2wRQUaRyGhGZBqeSHkOJ+/uuXrUtl
9NL39DQF/LhHnGlVm4xnQpL/LbW4woXj6mPng4ENeloPXU3WLGzwrVWZzJL4n1bB
Ym0VwAz+V1ATCn9sJoF02/i5I+HjfwGAxOMTDrTYRxO0hbOcmqDevMlpMEEIXZHZ
DSYIsFRA9jaxr44tbNWCR+lSpgHAIezDcApqHAVLT2vlPgA0zp7QZ5sYoQo5Ycnl
h9eIMdSRuWsbN+zcxwJ+Gr90Kn4AQWLKuYBBV9s8MI813tYtocnmt7OxrAGt9Dwf
Aq2aGzz4sKHI4pRvBLWZZ6xpnPCNdR4kttdY6r9S9DvYZBnLbAlnCMgbMYB08fNq
+FxL6JJsoq//CVFbxitTa9SWGTYUC9PV+hO4qjljDXvRCabH+09n6iGj8/Fq4UiX
IbhixKG30IXR+fUVi9vv022JyVn2IizmewbOI30Uj7ijFdjOTxWql6EiFpLEJW+y
jgwzGGB0ddKgUjXLBCPNV6sQUwzirimxX8KZ/qf1sgyTRwV7j59w0slrCGvmMLQG
cwRuLLgF9vEtMwo+Kg1BnHb827mPMlTja82BNNow383TtcuqgTMLMdM+wcvc/Ohj
9AHR63PVK07JGb2+r2HQoUXmikBKVDjhtELDB+HYsRd1ZQTRrb830PaHPT1GBYKU
vBtuonD6l3wUUq0Se7ua3uE/KUGWtUHsD/PHN1zMbTDdgUBUTTjS9kZyH76o2/QJ
kuBu3vITCFPr6SvYBCPvgYvKZD3llhukQRknbpa69ZiagVNuR7Hp6Wa/JfIeMMcK
mQ1OGrFPNxAbASMuu+iEPaDIrTAnmVScvE+u/iG7igb4NO/Ctisw9BTgLUlCd5NM
f4miL1I/LXNr3qmigvT0XHAmv66bFo5z/2XA/hr/V0KL+5+DM1J5X+1MaDLldgBp
F7GkD7bNIs3I2LBEEtIuSoOzJlP3Z2UE5wSC359u7dGAeCiMQQw0JtUfAN5b69rb
HE/QizR1TS9J2NIfw+2Sd6V/6UNESeHBXCo2ggyAQZfh3ppGZYUcmpoGU9Vslhxd
JojXUUypXbaSaOQ2jBRtq59fsAXVWK1wpDMFNdzSZqIgBDGg0QiFvwYqxHkz4F3X
EF7z/HDvF+xaM7RNuQmz4U0D8QVD2Njd4FuM03n5QhdmQFVBOExqs6HhnPZxs4xT
kzoAOoT1XbnLyN1hlGojK7m6DLMDASdS+Z4LUIohnxw+9v0kapDS8ppHEANhGGVb
sCOvctwW7K0U4uKp5lcj4MeWDrVfMRkg/83ZGxIVP6u97nCQa/lPoFoSt7Tjc+kB
IluwSzQzo2LUJ+l7HUbGe542BvGMmInNPvmJlqLzCjRrjUglyIp7jFImz8jzknfF
tqyuKZepFhvrqVCLrjPnkc4606sdc+T9827GCEu5pM5N7F3Zemd+6YT9Ol6CGwxx
dtBbjuBpAcfHAgeZPy8Uv0ADiuPmlVKkxlyagQGbiC4tk2nMO7Ls69+Ssr9Qzisb
vhYUqL+FcMXGzqZ1fsCGr3rER55pZrhqoJ0ZFl5qL8yPcB56qMKXz4zpk7mGWCZb
6Oz5cdwQeGg86sFPNaI7rzoZ285yRze8pLZDzT74gjIvCOo5LW2mf4tuF53wumNe
KJQTN0FHLlV0wi/b0KKjBxXzJgdSDJfAb4p8Pu69TGXbtdZI/orAjztwVTkyJCAv
P56B/LY458HlbAu+JKY1eW4KRuEghcuHEzipHFlaTTh+kPdY+onhjDp+GbSecj8v
odnbVcP6wsHrOntDuQO5okyvDj5bNqzb9K6r7EPjis2Hn3OhlDs3A2kD5kW59edO
VLEKT5AxZT8YdbqvKHTQMKNDeHqqQE19vqtAk3XnQ61xss70+zH+oqdKrbHMeP+G
WreBi8IY5m5Xnymn2bE8s1QXj8w7ahWtIk2nEBPIytyN0uzYfbfeHmniTJUgVXun
Mm2o/WAMvPsqM0M0MgeAJ5SoK/OxSYGF/zIzZeXAOvxrU/4plP7geUWsVKulCxI0
OEAcUS4gZhLWId4VhozR07MWTWOdAlm5txazgJzHmVQnkFvoBqeskXImboJ9hyKK
q1CkUzNiIvgyaX3BnwhL76mEagU05nY2OchUAxuH8PGJ3olsGtGYbwyby/Rj/thA
9LMA/2fE47W3qR9n5UddSYzYCivSZgYbcfVFCZnl0nWEwdnJbMWUjCHRRGMSOnMP
WCZNE3hpXfsIZrg+UyG5aLT4z7zMEi5kmyAOSBLg3GesACuKzOvAcasUtOaTs2ht
8J21oQhiQ02C+gGyq4PFWXPaHBckffOC3nDuhLfcUGzFWoeksXgkYPtalmlKCtqu
BgPf3oT6ZThErIktvaoBP7NTnLuvJ5lk/X4AWMt7WXYSOO0OQRKv3W1oMZyU0Py9
0JoR8RfStFgz/RukR+CwOqqVEwIR2L+lYM4tUATO6WWzZ6yUGUP+lrRZFIOfKMJj
5GgkmMjwDuN50RsOyjYOTRNjHRSmhn/maX8l57arM5NpDtjFDLUuTIcUQEukXBS6
ThLf8mRohGkxoZ684sUogtm5aBTG/z+iDD/9aIqWudgQX16RcsjFF8jsdy6lXawj
IyqQxP9ZB8EaqnrPzx51NRSXWTWoWu/JLa2mzTrA0Xb+oUKBpnQx4SJ3lvWJsXRm
xymH5ME7MUWVF4ZDfkfma7Srn9JXEWfQnhhNKXL+fpYWD52GZkP2PA5uzsVbxbH/
SkvKuBEItT6wAJCIri2NSeab+tuV38yZBixhjrI77imONkDDaSoA127O6g1txvmz
xnocaR6b/zLcaEAgyYUq7Gvvu02OwCa0qXgE2oPCeBrdjOh/SzPkeBnYGw/bG266
vLoVX8vctEfbjpJpDVDr8hrPS9GbMtTRL5AzFP8peH0UOq+8haTq67UxpXB+nrPb
MH8yt9EFnft6KQ1chXlXTnez8HsPDxyugGSSqSRnpnZxtX+k00A1ngtGD5i963RO
SZXMoJDl8nbjZqZHa+HfnuXCfaqq0F6+KOz7GpF2p24RgCP+ukSdu/5R5OoeEZQB
koKFBQgcnYVt9sRGixL8LwGS+qM0mfxAn/BJUxzbKnbvtYAyDuEwqHE7mpatD4h8
v6U6kX/WSrswjNXog8jVm2k/+swLojSuL/uhM2btsZTNwpVgZPYMtoW5b7uyIWrT
AyczkZwBxp7tfXxLQp0k3iEB9XnUMEWvwBUh8zFASIE94jIpf4x2nWWUAwYMOQ7t
NheoWwdDrHNOHisM4ExP/QxS5Cm+33sof2rWVhlsI4+lSrLaVJUYjwADWLldkc1r
cpdtKlss478grrXp/aIgQCLzK55LQpxUoP5ndXzOWtELkDA0DluR1UA+wEY+dXm6
huAy+Ox9G8wy6OxqkQ7e8qP0a2uiUz3x34QaocJE8sqmn6PR117ErBxdHxoKMd4O
qyrCdfExjsxvBVfmdg96eAJZVMsEkzIWDYh5t77B5QFQfNnk/yx88rq/zcfGv/Xt
gcuAL+H9dJbsjengMtB7IAjGWT6pizncoDEy2nUqGFMfS+SAy/ccWh2xu39JoDDN
KpAxb9onNWkbz01rhvVv4QmWPhBFz282b4WGRxd69LZmTjpaXJ72OBwUFr0/sd6c
W2oj1Z2Cxpp5KUBbgO3dLH2idM3+YueZTspNOVwJKvSj8om5+JjT2DhAv9BSzTbp
g6Y6mRAwbCetVRL4xu2yHDZ+i4B4tIE17IaQm4nyky429GoTMBOzigr13B9vWSNf
j4+3bd/tE7roek0bYUhEYI1Kxc790e4X/+3Ft9R4M3V3R5POFqDy+cIpE1Z2hLDd
aa5+iA++51hgzrZIJVyggWhEn5EFoivC4h8CXc6x6s2LSAcy/WxJJH2Zbz4yttdi
DIncH463k48zehOvlBs1VzP3+ZPzQrg+xS2MCIKtW8jgoL61DsZFEQT0v6ysb46F
CEv4MPTXBfx51hsVUiOQ3J4UiMi1eRbVzw1T5hwUfzoDgQHTXDYPmy2E4+g5JT5C
ALFn7M8oFGcmMfH6GITaZ+ATf003rwS+FbIt1fzmcCNmaVchUeuDGkmUFGpj9jX5
0o1h6JGWjyb5m+trHfQdEPaAY6+Z5XZlS+hhZFXeFz3ZvcUtUQHwvQhBP2EYaJ/v
2FFC3Mj5JINL5Nj3vlsJJ60vRvZbZyrIfdI813eMSl8=
`protect END_PROTECTED
