`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
umlIBaEmZP9eXB/gp8pIQOyYY9VPRW8YUyZOdEefAK3KslF61mcyACKDTvM6JOLV
VJzUisF45t5qPVyeuDvP5dRjEiIw7nEh0puKjFYMcobMUpLhgnPl2OqKt7rKXAJo
m+hxhQF0A87KQmxsM3LAeHOsx3r+/7TtyMbPqzNQdRH6dWEdOPlgmWu3mqbjdRgD
NkGIUVl/dUxtRLij6a7/I8P0wehwGgq6oBw2hG6KVBdQJAADCPgHatILO2qqWE6r
0MyM2NBsgmS4zakG4Wj8gLnyui5PXxYRAwLg8HRoj+gDC9ERqs5zH81QElS0Qbod
nBeKmtDlWFGpV2/hY5vN9RDZlCuUOQnqdXC1bt6+CAkB/pZ6fVBIeNnt+/QH9I7f
0hNl9hsspjD5zCDBoE0wiw==
`protect END_PROTECTED
