`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QvuJhrw8xTFEJPL8kuSi0fkPKI/v+kAgVGFucQlB6seaKbW9GxnzFPaEFbpu5Ia4
7K9goqdE/EP9hEirp0od+olw9fxYu2blRnB+HCMCXOrVrZrRi79lPZIX92XVu6re
qXrPct1D2KhkVPn3W3/w2wq0GWljjkz0zHVqJcuntGD0vAYtqdJHIbQ1eskGfql+
+CGbFt4BzBB9p6ghw6RDbLJWxQ1MKlM84li2dFzB8hhYtPz7j8pxTGT7jx28PNsx
ae04J54AwvYLKrgbi2CLJXT65PJUCGS/aLzM9kYMOc3uB0kdZXPiuV+4oeUc1maD
iKtSpt8IqhFQQPySL3+lnupc0KdywiL1CrzzEzcbftgziCwio80XHqb4pp2BrrXA
`protect END_PROTECTED
