`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c97sQXwNvHzyk1W0PH3xDD7QjNJOlo8k4zX2J/XfY7HkLI9oD8ItScdG6PdmTu4l
pa84gbuMIoZ+H4LOC/N8yHOBYFNnlSDqEomEff4Hw3LOcSkPYpuA2bUWw7djDDpF
cZNG0glgqfWlMBmKOKYKg+I6BWqQPuefkeiKCmdDrqoM/WqmaMMOFfaiU2v6fXsn
UImI5wlJcFY0QxHuIcRHadOrb9Gm1py6GESR+oQx6ohEW7VnKnKOiRT9DnjZ9cVk
QnOQs+wbV2j6h0LBkak+KFB5BvSuZ8mAquNas5PGG6vAZOTEIq/J276ngcghSCTZ
BTy3nG9GrGVonxZi8+UvvqUkhCUV7k9N4kM7cZOEuNfDSWKWntoKFaR33T27wF+L
Dm7P7Aw3o2b0Gfxrt0Bi26Gj+ggGHkiY1S4UlKnWMr7H1YtmjjuYlizqafmf4gEP
5I0eE1fY5XR9hlE+gEptS+HTNkWNw7Yf/vKoc2ipzfv92RJWEuq0htKzCY9lRzrO
9o5Vw1Q+KE9dWrZQ2vujjm1oV6vJjIuIln1fVApgDPiuzKNMbOXaWE0xJlCe74Qo
CkTBKp9fDcLrEjp06iFt2+lqbiaA6fyZ8pBDLvF37pq2/EuYhqPkePHXltDphhFx
T2AWkcEY+60fUAjARKFnzKLb/1Fuih3qGcI8wBZHqQn4Njy8n/fb6VjYS4zmctp8
0S+BMOzVh+RSS0CAQVEC02WqpOcnhtSDmZTxWbHIxTL5eWZ/eiH0qxLRzH5nClCe
5nhMwmTKCgVWhluPBCQRvmGv289cI8j87DXKw1UFH1cv9SgSzsafmBumiGuwPAEW
Q2w67cE7ZUd1gOSlVDIqtxwpjQxyCmGi0XSZjyOkZB4Cwe0RPX5iCFIJtm8DOaCm
RQUUUap0OPNyhmDlo1fRo2ugKADOmF5HwD9XwJ1Co4wqnHE+Jvm8k/MqLTyGG9T8
cbNF1YuGT5QLlKDoxrPIh438HeNxIo7wvg7iZs8cU4NuFjgMfyXP8ls221s7tFaD
ghfMksEo3AqQgC2w9xAdMInTxohohLjWGrV+y2M1Ww0naZKi1ahiIW35wmaFSJVc
NNpz52ed6LFwxcT4vEkyHJvwywN9L0NoTpqxc75e7nTfK65GeZCYRyQi/bOI0aYp
ECr7YFegjYZ/2wsBg0Fs4xulfBs+oA+ajLdo+69hCcQ1azWn7Xdsp8taIA9eSIYx
gIOOCar8d58EBjia8Kzqmuwf7tqeSzAfdY1UWrzL/EdZxlj9JrvP3Yxo3Oo7meQP
zNEbIpy+yt5lwWfFTVo1AHkqq4Z+D+cqODWN7xVazyh9rprqPUQ3PX7i+h9iUsGA
OFyNTssq0Gf3WIjRzjKbvxnjzagqZmGqkxDC8+qwZG5bmoaUXY1XMsvtnrRnAOBQ
GfAo0yh+ru4oi/akNlTF2MJyfcapPVlioNLMQh6ewfy+eKxFElhKhNs4qfuXUAdc
uyyfkdhaxedjplZKcVanBoD+TbfEG1SHsd0SyUFATjybu9ZTUgfg9V5VpEYCKKUU
AYvA6IhrlUXdeBvqOhOLd3gkUmbtHmxxwZFI48SxRB2A4rA3h2DKp6i3WMtaSXK/
hPw1VpTOz0JXI6VoRDz+2D9FvO2LziKo9ZMjhdvTYF4YoE58J1wjzi8I2QVtK8T/
u7jnWbujF7QyLA9KWiBDedqaz5v6vwJV4jUxggwJbAkimTD0eVei7zD3wC/NZQ/Y
NBO/xuEjuMGv1K3+EKvGeaBY5SHGfB5dfxhx81K02Lh6k4wyp1rGTfr903ycOfr8
81+DyFMQWy+8ZfzmIWyxu4ewt1oqipCAQIRKpCBu/hJkkOSUhZr+fIBeY+x9Z19W
pttIgGbriuZffDPdQ8qzx48TropLwTGNt7vqMXwplyWB6AVq9Qt3PXaTYG1rfsDK
oczv/8fsr2WrCbGq1WwoaFG4pryQ8T9o6MgZqQYCWCJkvWSSGUY2pZUUq1LnUcMB
`protect END_PROTECTED
