`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UmVtdiixqgEQkWmP82cJ6Eg7Sr7GiehmAuX2xLipu4zASeV6rLt8IEtKbGO/UUkY
b3pozhz1Emc72+BUDYMXA7JM0AWLFtjq7M+3J2zv/P/fsZX48my4aDToDJKDExGO
UvErGYojr/TJ5qqTW1eP/4AfGwF5aR44IihzXhn7RCBL0dMZOwOt2Z2VfTjddHeU
1XoPAFOpC4uZziuHdaDBkiT0ZsxpLojY82sNx6BgNNCDxyvsN2RqKkhFnYtOKq6T
14llk2v/G61VpOTY0l2HKNg4hYiMcgxhljebg5iveO8dFujVpT64L79njw5FREDN
ayBhIJUo/VXkmvbuZ1vElpphAtXLCavhJ0fH+goyKn9APjH0x4sY7dF14UKWF9P4
C4evRzbwZvLEiiAyaLiVDBRXhwz7xWKmCqbxHkTB5SPwW4OryeCkzCM/Nq1A8Jnm
MgvtGTj1s4Tk0lhQavLksIf/7KGmhQTsUIIGaGwtwtzl0ms71wdry+4tbpVJoWDe
p6GOlFXqlPW0M1xHGp7EDF0YwbE6L9GFwhmjNlQ9Tql8hQJWjZ1cfy99fHswD3FK
NcOe23SMRXdUjBsXOvtERpBfxpdc7Tpt4jd5a9sW1Qui065oIz0SEpUtSPp/2swo
GomaeIBFUl0SP40stoCO4BMJYhG/v42cECBK67CNzqqIm3ykuLdsFKW8oG8Z6FE2
paI79H8fgkv3o8cDZ9GhFnqFpDVMiaaBeQ326pU6BA3fhwm2cR1ZlA8vlCyvLqUP
JcOKtShsnSkj4ro/X9vt6aEpMdKpVkGVi3RinzlxgJ2yje84EZW8H7Vay9d3oq3C
`protect END_PROTECTED
