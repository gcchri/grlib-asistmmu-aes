`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wqaVmGE0pvpKEJKrq7hI1sqNDDwJ/hAzUmVFMVuwhXMKrYPZ/oF4BefCxN8yfsvl
mfr7C6/mPoXzgD46xh8DvI1iH6l9wOdI0DEoy+3bpy/bSrFYZD/7vUvF1ENJA99Z
cb1tulqMjdJdlFz3MClD9Mgv8aDYcb4M/hNttmedORiIB5gei0AWJx6HImJUtGOO
sFP+t5S/bP15hR99zp/6EbJsB5EzYC/5T6FhhKf5zsvEDLUXrzw4GIroBRytG8e6
3DlV/z0OopRheIjwlOpwD+I08gvuLcKsf2pimiVTapJWdxjgVm8H1MOkiUgJYQOV
9QX61Q40s9a1ztiTan+PeQiYP3WSi+grlO9oUz8TquhpIaL6KFYTbHxRSS0ur0KG
UUMKnLn4AUmXjRqcvLQU/QLNNo50SxKjjGAnb2urmoGcEgz7dbomypptuy7OKFUs
`protect END_PROTECTED
