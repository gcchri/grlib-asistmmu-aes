`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lIoKcbG/39kQidbNo/FGWLF4uZjAecV9R2OYuOYU+7kSs2yRaCQ1l3XM7HtEl3Ng
SEOnRF3+yqu5rmQg8Z9pcwEs//fd0vwO6Cd6YXIA4F2o5njVYx/gG0YPxzEnBqIm
gqrenZ+aHkWKklK2TUO58DNQbtsmzVJFTAuPRUhjTz1p5iQJaojWnzcuxMTkssEx
cGxVt+GKPvAjG05TC1cGmXjF17T5ZW3lWdaqn39uF7x44hdWoIGQq7HFD9a1rOwt
TtpeC2R+BVZ+bP9B/iGUAg==
`protect END_PROTECTED
