`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jwlbkMvQREJm0lVDlyv2Yhhnv+zON1mWdOPMtJ8YpDHWHQ7m8TcBgUjDWnauR77N
UNnYVfDEsveFZyoASD1c7iEnmvurOP4raeNtcDhx8Z0GQMvMuBquq13mG+g/YDs2
IzZrXLx65fBMzIGxN80j8bbVkqqE7P68USSvYCkSgkog2O6s4LNOgKM8NSkpM24V
iFPLC4zyGleey6JQ5wSSD3T3nMV104dfNGPvYkEdSVhQ4AaZ3r+AAKR7Eknzy+uO
LJgQdaSEdz0MZnJewRM/VDiIr9CSvIH33/x701LH/PtBnbChQ035iA4yBdvvTalM
MO52FBYrkHV6T3wz8/lnSCQIpyEPIVRCUWUeI1AcpfI/GzvrCTX/5b0kbceVg6PK
v6PNYA2gct22I3SH9kuDiGSdnTTyLXFajIG1QgYELOwe9Kly9Z7GvryBUs2CdK7f
7tcOzPE8vVMjqeMxi3az6vGMihyonkmlk7hC4YkMydb210FPatA1yl04v3lQh5dS
`protect END_PROTECTED
