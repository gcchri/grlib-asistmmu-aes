`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BGlq90ggl4/1DcZD8M2wHDpSM9EeQ4K1hUHsxKpmzJmekoGURG++rLbMgBpz3kse
dA5oO+W5OdCUSyMQe7xHGfjY5ZVqY7oVF6HfDmSH4i1Z2LO8l3Xz4jxFITiMfev7
U3prxP1vTBGUrgIEdjJ7V+BAAqaX/i2qklbQ+W/h3F76+LSiHgNRL6PUXEBrbhAU
XQqOikNlRMeyVgvG52zWZz0LLoBQDEFyEnppAdcXuyuCX614abpnVCow1CT07Dvx
`protect END_PROTECTED
