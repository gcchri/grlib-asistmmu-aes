`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q96x678MjrmwajQK2oVY/8dRv/KKSuVWdXEdPuyin+qi3cJ3SQoBt8o0bXRV99Jm
+TNPoDEN5PX9WT7sdkVMsKB6b0BiV8Jl7aUGgexzr3kJjzPsy+o3RT1l/OGylGIX
QYzZFTrz2EHD4Db490xawY4LfpuXuiY1Z7rmEMtd6zS/mVpvYuiozqS2TiZDS/Xu
TmnVFgCzQ2C9IYzhDqYFRDo/bfxTMbODFEZGNuuxchXiw750wO/P1jb3sBmvGJcm
9gTuE/z5QugLgy/P2bjFVAyif1IaA0rnNiaBN22lejMWxq9K8uKd0UJCMyPwjKjj
`protect END_PROTECTED
