`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZML1C2EystlvR7pcmXgViZB55s5ipIy/7eyAnr4WSmLFborQWvdzKRwkYFgQajdM
y3oII82EMnpsWqf+5c+DuH8aLppImu6zSdA0QZyNPUlbHdRIA1TzGZWZGSThotu7
jxen0yIgChG4ODkf0Jct1WNRfpDXTpevcnlehjXeN5DlVFbH9rhV8hMKKwf+3APD
oBCe0+kGs8hfa1vkc68dFTl4Ar746WTfC/fbDYkKFEk5vh6iBFuRawu9BURdB8M6
qLqbFNvc5A1hNuc7nwu9UKsbSsDorJgJ3CqJ6yNCajuumzBCbYLzHuwjLadk2SWz
oGKY8ORpszBoQsrseyYoQNbdF1wQ5Nkd0ZxfSXA2guD/+gkprivxlcgpIH1NQ9ZV
kbGv39mPrx7PVzN6NEoDbZJnTTdv/PCYk6/liSORbOoT2uJq2cofpetwuvPurlWN
RwZuECLUWG4dX1woDlsXnqOcwGXQ0M4DxYsF/Rejq9r7NnoSRx3jpC2q0XDE/Z+r
XZc55cmcJ/WtfBjkTDZzWE2FTCA81wY6bo+EXtJhT9I/i2o2OprbJdng89oIfgWr
NreILve5iZSpJuaDaPCOLc9BVxNknYSXzmKR+aW/dLnm/ff468gKvrQwcEEAg48I
fy/Mw8CI7ipY0UoY4L87z11pLDSmILpco3Q82DhCGfYZGxiM9hRkk8niAkrFxFIB
Yt8RpHLcaqTFVjax2o+izv90hXwezg77g97C2w5dZVXVVGKSdF3zYGOYZsnB8MwZ
KZ+rBK1jgpcOc54UKIZtpyKC5nJEaitxHCJk/ogiWzem/wmevVeLHRIjty1f6Xvb
XU3ZH/y/TrJDu5xvNtKCp2I+5jPErG1KV+Z/k0fKLj0sktHU0E3OuxedglM5J6WG
U/4+QyOEFLh9G+cKRSYelNCDFhGPKtSprwFbU6K1jFc5h2m+r15gTDcX067PMM6C
kT1PK/K1AIuqfA4cjtd5S+shARkY2yQZj4eS35l9BBHZv3fHPOQL2jQhOgHU+gcS
MsxVAb2Ww3sXaIBro2q+sw==
`protect END_PROTECTED
