`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rNM/vCiJLb5TH/vuI2nPHbpvb/pnmEL1dirFqmcGJVPKQVTv6RZHP7rTya4wWbtL
eZz6AnMXrTrsJK5S81FKWOqXRdk6S5mu7yDjoa/lC9SN1ulcwo9UU5RctWRbQXxx
MUaPRLIc87ZDwsKM1H4L9Ln11GL/MaO8MFMi0Jj5FHz9nkNG3dH6VndlPMEB4WXe
b3KCZhNH1qMdkDHmfYvSViNRwYAxnyAZTPjBIUSrT08MiVDb55CPh9PQ37EvT2g8
EA5RVwi2vW/8sCY6goWnXBDqAt12jZVz3XXPrPI5eMGsw6l8i/YBNKqEXa0/mByZ
q7eYote4bGjHSiqcXebnzA==
`protect END_PROTECTED
