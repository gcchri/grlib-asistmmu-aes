`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
buNRbd3W5GDaBjB9WReDDSutMbSBiH1vvmxL9Ls687r9iFFJba0KbOyexiVlUlAq
0MNNCMR2nsi+osQJpiXFxDkonEBzXrSH549ez1P/zKlwljOAyVLpdtGTg48v32Y2
4z47KUFoG3A1DoHOL9/lYvi4wx5rkRotfebOlohCPzOVZxZFiZBDeeze0gXyAqxj
oa9z+eVqczmpc7c8XLpjZtHVVww6BV5zBJubew9P8i2+xO2pDoBvidsJvf75uY4J
e+raog+5pCcb9GlONbCyAXiMDB73C9WipTyWM4qSA8PFG5DQ6febESSp/OLJb2X3
gMU9J+g3q0WnEGLDfNavog==
`protect END_PROTECTED
