`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IyTd80KZ7X0ju7cALQcsF6QLjKy5NJUWgILKz07BVIuKdlOI1T2HOyvqRy74sO6Q
5C8GSZkAawZ6Vw97fjtFn1v16egCyskelJDSrIzJnXF10YmUgm0LReyK2mezqN2t
nTHy2J89f2Yk54ykcvZFG8h80lzrTYKiyhqMziqGsRJ1SGIfwdgBwFSSfxOfTREV
7wHDn1Q6PcsCo5qJTDDokuNfDJoZhxeJJUzaIqZhYYmIhtG8YGKMTR6JikUZEFXV
8xPbF3CCtzxI7T4nsT+T06kNq27CDaNYLmOCh6nzfk+Fa7Ofhyv0cK5E2a4XdL18
iPBlSXbYp1KX2USikZ7xuB/2NymxggZdxATAqLgWN46rn1qVLjBC3vJb7Gtj6K1S
GYlWtUwzdlCBnb5NJh4FkJTvLg9t6XQAQGpkPWYQXh+4svpx+Whj8yOZ7sIpZK+A
GCXah9/N8YwkWsvV2r9gd70x0zwxSpu2BkfNA92lNDSfMVMuh5/+Xvx5HHuI5B1i
NVQyECWP2NFeBY6OuzSAwZ/g+taNJA/ZVP8c9XsglTyEdupEBklZW3FQWx7VE2Td
5V5TMq5WOq8N0Yyp5eBEcso5NHz5dywA6yGJ++51yAoz6R5NqR69b4lDeznMcKLp
ohTseU3F2kBz7Gkzj6J0MUsNUEViVBqYPHOWm9JqtaYtU3xi1ksdaabrODYErqtW
rhCI5+CP+Qp1fTgT3kX8WBjMm6AJZ/t4149tVvMuAlLmE+es0/0Jy37giH3qIzhg
616fR67JwnlhkAO+jBKFgSxnmYhgfe3JWBDypg3bB5iQ7nobC+pADAeEVBvKvM/b
mMP38jheYBQTQOXdBviqJZgpwZ3ByCXVGMEIgMqblpgfyltoUZdMqGiEUeYDO1og
I8GJA5+tmXN+jkVm43nRFvK9ztoO1FObXcTBN0pQ5I4WVfSSAj8c8012fB3W/RKj
wTzvRlN6R+MIcTuJ6nstjFA00h+129rYnk461YbGVgoydCKrOx9WIYeeFZWzRvq5
`protect END_PROTECTED
