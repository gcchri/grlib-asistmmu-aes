`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ETGF3xKnss43R3v9VC5qKXYqvNyaUL4UleXXTKHfJ2j2dBCye6ZWeNg/O2IDPB8m
tqBDeDey2vn8lHrgVPVbjqYCh+iptQvA5kU6Evy+7gr65uMKjVZ85o/cPotq4pZY
POgDnTnFyrdlTAVzL7QTOEeV1XaLQPvat+XUScehUi6jEJmR7Dbs92+i3m7dVkeD
1SMSIUsTwTP7gBdA0l2IrGGelsn4AFAfNrOeG1ljD7RTG9sLXg9qOeo+b/OSii+Y
67q049NJWNaZgcfJSGaZC5Gd61HC+ZFUcIMQitt1/Zq6j03mmrd3QBWkBDRhq6J4
p5LbiVniS4cpaxhPRPkdyVirXuvwPGJeK3sMFi+zJd2PQROAo08aVCueLjdCDuMj
j3Apjf26bFKFb9JeeKBHZFQP6wp+NMYWUfuinFHhI8X7xDX1g2BQYOIQVo1J9Vci
`protect END_PROTECTED
