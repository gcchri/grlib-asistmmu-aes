`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QBX8uhS2tBa7hptPeZFwrIl3VYEHkPTAZuJDeDh3sFbe34NOcu91E+XEGig9r42F
py9ExOXgi2NgICEhQXNVmFbBEy/OJnqfsHiyWelE9KBIb0+LVDRV6kCBXCe5/z2v
i8lsv3dOXjivjlM7mK/VqhTPX13HiS37x7m1eA7W02PX/C78h6gMp+vHML+0PlNA
Oa+s5LqPnUepCMHfpHqWTStd/jb75Wb+hHBP68VCWzWhq8bTeIZgBi/aCt2UPMfO
xdPnlAVJht4xALZAehqXtbxxosfP7ZkjXNFNnXUiRHy4EBTb26UXf4ToJXgmSfnL
BsmT1OI34E4eZQRhSIq5a+m5izBreu8/3ZSHjT7qXpHLm3NbyK9q0hy/VxFP9yXQ
9cfc67xWcmW3WvxXSUnYwZsHFMylzXTQgDhcC9IHqQJUGCkphhU0tG8MGf1uLFg7
P+dDo6t1fxXrAdf4l1jaIhcw/X/qYodM9DszK/vVbGR/zjbpvoBrIT3sgyEQ3NED
`protect END_PROTECTED
