`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OLvFtCcIxlSmKUcVrDa2V0Rhx6MB0p2gXGHAL5ulRZEtin5USwpOU7lzuV/kYlzM
c0O6hgwT8wXW/UR851aH50F/f/zOWJ+zyHBE0YNB//lmp/z6KET9M8jWdm6lqyNe
8HYbWbCn5t4gvT37rHzHQ/UVhFyB+/48CmSdlVfikPfPDyqVwR3XWSH221mZ+FrD
/lmgt4zgMZKO2MJTi3c/lrtlGD8mJ5migKs3mv/dTsaUayQJxTuTAtux6VKPJEXC
P+cgCRa8D7LEPpBmawZK4EijL4XqdHA6DCTecbDQeoGph2PsDBggBOJSFCc5w4+T
e4vaekXZGOtY0bYeYSjETjVB+uclpHQVJa42iP/wsZKM7+J1cmF8+jv+MZdqAiHF
fGWVP49cUzs9ozyfCa0QDSQefzcFE33hhWjbTb3QQTuoUmYiRmvbleBx+OsrVzGd
4QuE4HpVZP5OoUb27s4wm1HPymDNkyWYa+VASoW0DTUMRw6qhFisfSgYPqTAhV9y
G41SpD/dDTPzBKOzFEMzEnMqYzbXBFXHZPbaxpOzo7VCzLc26Coy7JFh9ZaZbJfk
TVpgP3TO6q28ktpQsORU+RwK/N1lbn6uCAdZxp77YLFDBdiE8lpRMpl/NJ2R46H+
vSPluWFY+WcqfwXdyHOxzingoSvvTPzNJtPEXJtPxKrU4TRNHuKdKfv7o7Jdq/Cc
9W/F4lWF3VDI2l9krffNmp0F1rwxhFWOAB8BMG3wynDlrwjjV8nlmFj1yX27n1x/
vXzfuqXwnoAG4rgW0VfwRRXDjWRri0ne8vDG9Bs16/SM7it6ZkjYriWO3l5VJ+Kb
HskE5AjXNyRVOh6nTvhekjsCoOwJuKuqd0IM2CHBNpcQTtn8FOPMmiOKK6TppG7b
eKh6ZnUVx5z2KOpedV9ZmJgEFKsgMvLW1kW/dFqiRHlbkhB9TSnFDs8PK9+VLqaU
ditdmEigKIf+40AazRtHTIpm2KY6DvoQSR/6p0DfEaUnHO2BVZeTmAbEMEPPIF2N
uORCueZRUqzF8FZziL/iEl4zw8oAgXHYC0hAlCtLYDbwVqZIkFPNVmqpcvQCODrW
fS8TS5LCLwOUw8Nxzj+MnM56+Iamu0/kEB7N73FTO5VbfeGkAqnwudWnVJulp9QM
UHANgs9biCJ/Kl6uxe4cbFWuWjrsZLdRThtOZGfvx9csroP0Vs/QGoFJJWNzlPms
YHwp6qH9+b/heXlxMNelrujASkCu+0nKcFQY+YlKpTPuTtyLDgj4dxyC9hXYj4Xs
qW3GGHl0nC8bMrFbKiB9xQMarJDRcrp7l5mrfqXUK/WUBvE+ImTwqlIsPUTUTlUX
KCfuLqchHbwBAajG2bI3PgYnG9eBKDa+tC49Pwg+HjylMydyVfEu6/+LaL5YfmBl
WExMevsqXnH5CYAuOY9g+iOV6rB9O3CnV8THtJ/6516vM9dSdldFaagYXFSztJov
PTUMcN6KNQXRDD9JsPOxzejsjNETcgAaYX22v6cIbAZj1S7p2hMyjPv1dOoiI0DM
qkGBQN47F52opYPmZKsZLEllqiHYyfeHIo1i8fmt4eYT0jU1/bidCzucpifC6zkD
Njz+xhLz5bsqFLNPC+/XcbdhvXzBLexLVH1rmtpf/MCyoHcn8nRqyt2rIWhVYE1s
yyXDbxhb5mGroEzOSYi/IUq7bJJ45+DZdT7ukO5ohYBe820bSTAQG+5YwW5sFL/g
6Bnh77YkHY55O+rmxC+S0417hzoR5j0Kf6oNnk8qw0l+dnyqvppOOEHjQ2R28i9a
znILDv751X6/o/e7w3v3xnBpxKTSS+BKJvN7FecPuWba0AKsIrRkOwohgGAW/RAD
jTeE00r0y6BTjX2xtcc8f9DZVQ/pHLDm5lSzA9770g1uU+z1oyc0zPE5AO2DiOrk
Ckbh7p5BoCDYcRMMN0qz4ZD8aanwfMvfKcjglGf5F9ftPuH8bcLVgLPh7XhwSTzo
P1cBLOruYTu3f/ZQEzNOQjM/N5HuNE2NmKgY9nMJ1fPMT7rpFndFcZT0a1sMQY96
R+wCoeDaZt493aRNdt1uIpVpTJMH49lx3MJQ++evfyngao+jOKs8fzznQXG5WYUN
OVa1RqBapsU1Bs4mdM006/zqCeTJOmiPO19evhCiW9KuxBOzwuTj8tMoV1FsBlGr
VZ3sST03OsSSw38MwomRUOu/pQmeE36xM3zS1VJeZq3f7zOBJxJoURU7buecudP8
567UKz3HKdTanm6gd6DksbQzxl3DFDamzLmg30sWgDQQ8tGKIRyKvuMxrJPil4Sp
hJ6bjfOZF5DP3jACirKB/5mnfwjHD5nBnbFXy2LN2mVm6HsCrGAvDDoICo5W0zDC
8Q3vhDPlWfjcDXab4lPa2eCDnIWGm0V15fb3qEWabuoG6w63MQSZHh6LxWOyEAaA
kn/vm/QCut4eT2/7gT7F2ZdzkPyDc8ytYIT9TXc6TwancfO1YwSiOv++fPQQcNWR
iO+vtKvGpxHUExv9yoPVRTcJMRSRP35XrpaHtThNRkCNru0wMbQgQBpHltkCeqOx
E+OgIvYEz/vy0aglMAKrSTq8nIuinJIpYTmiju8jjYmWaHVpfGqKcVQO33Tebytp
zgR4MCftCudXsXN2rGOnmkHtdlsIu34kbOkShZ+554cYNg4oZCyY2wFGKz4xa0N4
b4aOlO2kwpw4H5i/09HyOml9NSBEKUfSEK1aBREHtjQlViHHmOXDIndUGPNXu4gQ
2wnNhodOX/Fkq5m8YGE3kZlAUG5sFHwDi/w/IWZPqucnYDYo1FjtHUCKhWnZtifw
yVAjZqCDVLoSr3RL8FL+NJXEbJW9vybsnooGqeUF4+Ir//+vwk3EHfeVldydWTIQ
4Nup6e2PGN96txYkJDhfV3yu21dtLB7ZS7230K+UzZFhJk6cIhatH8rZ+afiHEGD
Z5Fi4JKX4llJS+1vW06n8tox01baCxhlfAj4DqwGUjY/bErOQNLN88SXkUdUCdYZ
rG462P5Wq/sVaIWsiewfYmIyWlu56CBlT+S/4v3AgOa7/riEakrJaBQ1+yb9W/QF
Xij7QsAUskJJ87hOETV7AVdnlrlt7w6eN09sFBDgv4vdBSEmP+Eg81h/l+T340BT
ZDdnhNw5cxWqFwIM9Xi+BNphkayjxTRAU0qugYl/E1oD96+O/BH/OX6oaHqHvQag
HoL0GHNnZlrfeAA+zBstQmrIM9NBYFtVelr86VQiMOV4kaCQKxLW8ajWGOSVSzxS
UIwsdUBDgzqhqEr1d1JbkLT9yPn0LDjOUT5wK0PpGoUCV9d2FZ7DQiHQBX6dxdyp
0oKWaX9F8eFOvjycR1XfXYTcrQsaYT6bCHnqdQG70ynvH/1fN0nXlqKQt3MgDll5
PylWQxjxz9VyQiZwPeguf5yWuuvdYNIDjcLXxBcglYyUBqfE3kNI2XblmQvl0mym
N2K5CdYZoJZasxY3RqrYxVzU4aYdvEma99T6OUkKz4sWciLBrVELovpZxzukZJXM
oZZZS8lJCSWi1fNg/gnTuzxvriDwxXLg/ipkewrpBgoD+uNwzx28uauOEvSJ9thD
vPi5mTu4mZr1eqrfsKpkIBijhA5KSAxW4Quu2RwoTqolc3k1IpZAWSoYI5+mEJVV
yO7GhzCL/XhEqTPv1ZbkXVocmKJ7N5q18idN5qTPiocxilJiDgSsSWlUWQMPlv2M
QQs/q1CKlyPkyTPCybvxn4fKwYVmzGpzjN8X0dza8ey7XpCQ1d7d2ZKlyzzgjy5P
g7iUTA/A2L+3lsbDTQL7HZ81NNw/M5l2TRBNVhFNseyGBNI22ghxkQnJxihNgqEA
fktsE4Sjv+FqSYe0F0cLRP7rOqJxJ1r2EmCuneuIzgwzWEQVpiRKWPG/6useIax4
JgJ5dvUsNKXrmUDod6UG1s3ERP8RDnDA6fzg3UhjoHXauI09M865M+j339AcJg5u
Nolq6u0o+DP5VPznp0rhRV2AfGRDy3ewGvTFuPTF4PrRBxhFlpYqRjxJ9OwrOEhp
vE0tYiBkhhMXmDWSFrY/xMVYC3HBy1vxfxJrrAzbyxrLZ4Oxeyx+UvoxWZNr21sm
8hb8csVDPxD2OCvUH52myJjxjWrg1cNBikSjxpQn7xW60926SYxlXcnICNnJQCm/
3DJepyKMn5Eynk//1QcEI57UXFV2fLc5AdLo+/n/e28aHzXBM4e6E97G/FpksPRv
tkkCY2rzB6xoNbU2fFWXYqzDMA8+28AG7iJtrvmMGbjQK3WASp4y+w9H8zxSykL0
RukXBhZG+/EmMFVL7uFYEshQ6WM7n+dgOsrq2HP9/sWKNGJYgVncBM50XFFiqf44
RtlKNbkvgwGYnggJ3hYVrUywLl1XCxdjK6PjNr9muxtgvNkFVAuSyDn0CcZG9OPc
mkNN9LmyqPvOEppPdL+gSCBG0XADQDemCOGK0fbceSpPgVe2+I5aAs2fupmKWGac
4Z+EjnPUL7vwE91rmJXBJKuC3Q0dE8NafoKf4MsetMVzHxKSzSw9yjub28mvL3FI
NFgrfRtjMFlmMghLybb8GKRmlR29nqAwjGwwMIPcPsbZqwHnZtGlceCpK7hyZeqP
BVUrfJFcpSFMNrJhL27LPm+/R0T79BTnsayhyr6fLKw/uOWq3ISDtsV9NPdzM+gu
55y3bKlX5t3eFBnRq7ZZRs2YOPqWbkJWgXDWLTP7Xn0Qk9CAMOYUNHTZdfi/X7zk
aynaytiGRsD8SAsc1fDlSctx3uP5056Djfb2Xtvi34DO2PuKoFbyXaPDG3SJHfu+
qI5U9aeRugtoLBK0xXvolZNHKLH56ydAxVLVSBOejcUWQhvt75hoXoz4d3gaaSCx
4zJNV0wIEoh+0cX16aXpiH+CD5kwhuIbGzcNHOJt7LqIJoxMZGz+UjNKE/kOz0Zo
eehqeh2epTHRfrkOF98IrcpvL/wMmB4IHKWvK88qO6f9m/ceunSzkKf7YTq7VXBa
6bL4WFEVrPEvajy2Jz4j7wbWoH54zRWusiI7U/a+qHtgjW5XENc/w1hUSDtj+8hq
v3vK7wGqhMdtf03lusuVIZ2FMtp8cAvF2IVdiTXM9+sk21MJK2zK2huFCSt/g7It
hIT/pbReyVCXFHcSDWly1LwN9F/PRHVsXKH9Z4oLMMZXPWd4XF1WpHpWlICzEwNO
20r0qSqQWhOUmm2rVst5jsLpd7OncH1tAt+upJW6n0nvSEoEcFmHMX0kxm+cF1AL
OYonSfFg8nV5HudSRHdEbEwT76g7ScM6VawEZLrtWLdb/XYjLu/y8Nh1jcTaJbPl
cfn5NZB2WKQcEbZUOrxhdQGNslDRkxxsCgqnyXZnDkoDXxNoKj1VE5sxKIgDrXC2
KmXcl9lzNfRpNgFGo4xsSXVXdV9HM6QuQzIB0NHPGN/Dfm6WU5rzDe4UujFqUGmt
zbl8xfu+EPHu8y1gwU5PPVwhqC6N6u/zNnDV8zG52FJ0sjbZVcIGSEu6QZ0vZ8uu
rFw3lJHxyHzKJ+oDUm6vI8FFXpUr2V3h5hWaJ69Jmc2kMN++WYPCiV8RjJc/sbjN
/f1sP/mC8SITk2AuQ6V8ABvPE4zCkFN8cTTa+p0UWY75V9JxLiO9znwWuuVRVOHJ
MiQvYHvdvne1KtQgA9JgocAcZM7iSXH65HmlafhiA9lZ+xv1T4O9vSPyqz5jV+dt
+ZOWNBtbxw0/IduScTLnxNcNvjp3FIf79d2+a+RIShKfcgSkSmw8Dv3CFRI5AlJC
5kWPVdSGjIKAeE+slIJFchm+QyQglOH4EjoXUIAvUSV8C/ZFthDnY+O/tiZh/2Ms
AY9YTYEHg8i3kLD4DcWYNWl8PCpwRAguQzu7txRXCfkwAaDcBy32rZaUT1x562oG
qT3JolUfgPPADNlvN7ZzXgHqRYSNh3Q399WGf8W0ieQbCUxZM43qn4AAGY+tuoi3
t/Ax6VFYcZhxKq0vKfcGOSvsSbrIokdtsgpwH8Ibg0jdoTlQBTmhZkfdYpxhvrGm
WUVkkfiQIHtJcdWPmEkpbzA+0spBcOY2YxnQMCaPPBvjIrtmkxVoUHgslWqBXAy7
NTcG7LKBk74Z0e86TJyXQlWQ32yTKT/gsZxStiRtomKGUR4lqAXnqzUwFoasHB/v
S4iGwCBB/a1uJddaC7c2IsCw3BtEnTky7iTM9PmAdfytMlpEANH+GHKz6J6quc5y
gw+17vYqlRadG6S5OqcZOGpDQTeK7s0U621VyS4/4vyianMppsBVPkCIsZO8pFnV
bP+zRdEVVmsookMc9+lwDO38ZpcUHw2xEQuULB/iLXD51r/wlJFWRMGe3hYLYOXR
8hTkWcRQ7ImXPNmHugOYaKEIrtl57hmiJQVag+DLbLK6GLn46gOJPaAz4lPdlLUW
/viKYTNo7kdFcBSuYcL3M3IDWbgrvulSuIY6464zBFyWQfjolFeDyXvTPl1oZpDQ
jvJ2QPfQyc8TgfWAngANzZx6tc8eCfGQkeRVvD+VAtk9nt89kDvjtugmMZYwuQUB
LkpFxSvrlihNtz30PvK317sf1eBUyAG9KQ4VnTEjBNmQ3805il6wCHP7YIk+5GyR
aumGE8QpoP0+RRkk+VV+4+1ZNlV+I/gdvb85zCoYUidzNFwpnT8DMdfpaUyHyEa0
QMo2VxI9Z0nQug/1sLOwu8XxpBQxV3DJntf1Ld+MAQUCEqoRI3lL3Kr6GkJ6GUiE
6tGPlfotHlpRv47lgwSFqYZdog91ORcvo6sqMbid2Jzl4oBGmjCLHK2GIHm4HHSq
AJ0P5Ql0WIybtKpHclw0VSGUyktnxob/5nwRQrg6o3u0Xw/dtW8f5qFSbuqmAVEk
FiOI4nRT0XJYB39FiXmWfFg4KoN8Y9BcGVRwpgUOaW6IoVV/KkQvKmakvsnBiqbU
sUIByhW9B6fdVDQIjduzo7SQNkBXmCdhbou28e23EXqOp3d7ya6QHHmLTb14fLj3
PZHMAWTTAsCrhA2AJx+a9bvkQMyhuEFbvdloCxhbZzjAPksT0kbFq9cNf3494qAs
ygixRogwnSF0DvmgsNcauDPEzJB6zbnnNdZoJZ0xxQvv1d1owV7sYK7PtouFAZiq
ktGtb1S2hvPOJxJS8hmh5DXWpUV6y6EwhKRm/N8o1l7075l379NiPXGn8demTbNG
qlQwgTOBS6d/S3XCJKFhRhAGvtNHEYXVgoX8F6XOyYs71R7iXiJnDf936hqe/gPy
XyvoYBzXcdKRux+VcSAcFk9eZ6vLljEJ71eL/ABOJCeW1u/9Y9XMDMKr5mMNwTm+
9B2JBv5tecv03rNt6QsfjoUtG06FQSUCbA/TdlVMqoWmtGCgBqjOg6MABVI/WDra
EPSFsle7M6zE5OyunFTiN8SSE3md4/KcuWVb2t6wewbJSrCK5oCkk7HaJ0UTjF7a
0qRpjL29SHjTRcRIFkD64D+oJ0x47bPcpMGqNjseiThq4OlI06P+/oIbrq72XQs1
B/Q38xIw4v/B+qIFAYaeikLJilVC5dSTxO4/uGkm/9bgVzgATXAnHCuDPUV8HYQX
RhLm9n1ECzvz1IDuzGHv8X4ieCGYfncJYd8DR+iyNfuAjEWLG02dfVkXaOY9xciD
tV4vw5LtjExBEtdfiWGfeZFo43BPjurIId/I7Y/jb32uK2IWS+n89VX8xC6Loe2o
/2I0JzOQrzoQdO1dsk4qyvXLHpstsXtDqPj6Y4e40H709nsIe4wpONg5AIzkkurz
OQib4uY1wwrUcIdEOy2pOTu19IMYJNRrEbA0Ey7VpBJSgNDW2SeIwcOooLe70FQk
JmXfhI1/70kYAJVI9Vzy/WHZBUgFqq1DD9FmpTMUN5WXX5xv5jugqEFsk2hg+uvf
eZiPruFfqygu2nY9l/1ti6Zth+2EO/LXC+tkW9akFEkY+HEI7cGvC+cQQtujtOMt
iADpR8wPQLxBT5vVm2CpZpASaJ8iwCmHDzyavUCx831KlStNTCsMjiQkbaPAn0M5
vQJ3dBPGlP5DxFM0TnG0sIJmO96GG7zT5qcNjqWxasBNXr6wd5yH18EGRuWk7k1T
1HArPBGKky7U5J48dj+FntnQbhSlsEHmZHJrzsfRpTW4ypA+xeqSTe7zCXqb/BM/
5k86EOnAdjvDVlZiLoEPFwSi8ueSXL5wEvYtAfQd12HboT9yWnBK9ZNsPJdaH22g
QDW6IRepsX/l+ItOWuhsNYrqOnbV5YJu8ZoNWem0m+sP/Gxt6cHdEVbITftuhZ5Z
u7Sv+A2BtkUbkjF8KZB15HVbQpjpKJjqmf2I03ORWMtgCG46f5IicyCvYSLU/eze
0fClJEnLqq9on1Lrug+9k2aUrP2KXohnt+HE0DKuR1qrBTAXUuTB2D8xWZ93BOdd
qFHBpEbYFDTXoeqRFJ/b55i61cf9c5yoBHKCm5n195+ld2cn2kgyCntYhMT3B0mG
vU1WEoJcbh6Eo0+hsyJawJU6QcijKMqTCpUVZW0QpeyiM16tPq+SCny++u5BJpgR
o3jeXEka/QF2KkZ16YckIUKhcl2qQbpSMHf8XxHnhlraMXAsmiuBYfoxKA6ZSwLR
fbPzylMciPbHKRJ4Elm1wX4Hc2ukkk88CHD1MaWofXFmG3gpadX4W9WMjBLmEK6g
A6ZFaqSoc/g3Fbp57mSkO5Q/zSAQ7BE3IK5OqIJcNFw5abbJQjo8LqSNQFI6qyay
ZhRVmDfZ0weu1BwvT0lWRY7MCspMkMM/LxyA26HgtUNp9DZ28cQ05ngTRLo1ycTK
sJQEKDOptQFF4N6goqk3flARVXRCUZGwZjcR1WP2xdnR7YJafbxGJvREuAEJy2uh
mju0EWfnIMMqPlEREf9vkwax4T0mLljQ2xQtC8F45xZpTGcDrINnYdpeRIaUMASD
6MQTKbQ8eBPiWrsdp+zjODg4nEm0KB6Y/3tPL/4Y5jagVnhgkwHh0HPb7YHZAxLP
uVzK4rk4rCdPpKIrU9dELwm0MA7POBGHodk5qHwTS0u9x0o+Q0/7qZ5fjKZkdr2o
yAGChM/aFNYO/P8KNZ2nsXFl4XooZWhQV6ss/Tul1Su4KzPZAkA/q2MLFoGo7uTH
69aJt2j2jfgoEKN7LPs1SxMCDfhuOxBs1zdjasvEDD7K2HByY8IaNZcCGnyMR5gu
c9m1YviSKti6qlxTCng/3rmgiGMp9FKEOv1zoc+7wBfYRnM1hCMfo8RAA7eMWRMv
3rJHWVOsNd1TJMYGJQweOzp4fCaDEKn//BtkOJgB0QY1TxUKayvd54RqFbkGJnEE
U6TPRXNSBxmjPISq4xIqyFA4nUXGZEZ7o5d33PcDd1mz/cgW9r1vhvwQzMk/kmmz
GAtfsEyeiNAIPIHcVXf57b0Q0R7dhlSkHgF1BoH74+XLf2mB9Xz+xYquc6Z1tbf1
wh966eacAbKD3j5TNlU1C7cMTmkDrU4sYTXjIL/SnPJU5w50AivTyZ755bTYv+Bj
yBxjOm930b7rl3cK8kOM63SDuaAjWGR0LghvhNgPLVojMRKwhU6YYc2hu3w+gI6F
kvlxNXJGxrpsG1szeWspdB4BxN8+gJkVdxNNQ3oRZWFE4tGRD4W+L1H3bim7fOLO
laxiIoHbWS4YW+2RVJaHgzb+ASK5lcpTHh5B+6GMuTt+Q9F9subhqrF7/2He1tPF
+8WcO1RlyN4oBJmC2ADx9DcE76fZAg5FkcHsDPqlMDjPAUVjovz4ON4//WQ5pxBR
cwWpE6HOG1+vkNxHpqdPV6QVR/yZ/WHSEEQxLh3ER4ZFU7+SQ5DqiUg/yRkpuRJJ
iHkELzS0C/ebUCDmsu2763XKiMkI6wYXx1Ww1D2UC/FTGoKTu0QeZHLF/5QUqNwC
Gqb/vFmKvwUMHN/O+t/a+HM5PU6LcrZ9n8BhhxyPSsvhdQRVRfMIxRpmsQhkOU5g
NsfxKBYdSKVSFhaFkcKftTADIWfnij314IFX8zs7AE341rb6mC9hx8BcsoCYApYd
f1jutRqcRZs7irU1ytnJGOEsrz+5OywoSDZLqN4kl9epveiCtbJai5KZZHTI9cu+
coeKppe0qNmq7e1xszqL+87NYkRr++hpuTn4h+MamI57NWTUBAb1gPbe1E/PJqaU
tvjqv5cKYmC3/hWAIiNHw8JNgJd6eSjsZJ/OEnx7meOuzttYNGO+kKfWOvKXROlj
b2nRsbDatbQL2gqoahYajI8Ud1QAme3PSuwRAYQyJnKsMyYsuRqjMLoDXbstF+/N
l0gIXST/zmynNxkhouUWh35XH0CayuvdZdROcsaRSupfbW+6DvRyTOJ1GIsD1eb+
TSg11W4+jf+69I0oZIsRpMpdpyxVVWdcBjyWb6+CalEd9nxD+mitLqTd0bwBrahr
qCAtj18fd9SXuY28Lb0BrCzkeohsBVStuU2MTAhgQA/d5jTeVSD0ljnTO0b67nL7
erHOA8maSr07+ziup2FoJCzkpd7qBwCKcqUBe2aWyCuPO9/9RSzT3OAq4Oa4rzUK
djtCPa14mS0XmnbrbDy5QQwWRW71HJWL5WDHSdLZ2cm6PE/zpB+rIJ4JJEC47St7
IwjTUt8HabaaYYOEXQKUR+h9JPbPwkpm9A5yWxX9gVHmlhEjjOOj3u71IyK1IZr2
MVe8ZNCGPjiu2D7IMPWicHrkSMTmOoB+1MqF/F15TDIqCB9gz68f+onxMEqiWFnq
sKP7tE/ah9LNd8Uny7TIofXGHP1VP4XotNVN+ull5B/jjoaBmjIml/RJqTMS7hIv
OssnK19NJ2PLyw1Yv/fBCyb3ed7uejfW7iw3Jls03AFZn6YlOG3YJs1IyjPjqsFL
H8NH69RprDMUUavSuiPbaYfa6b/BszqFaxu3Af6wTee0/IwfiIvNaNlcfGraz+Df
qd+eIU+3ezad1GXPYjFr49llFaYikEz9U3j3zLSgjHOpjUU1q3PyT6BxmijxIA2F
pAHqvK02hI/NJneS3o4DbpjTG5rJlwmiMqiKTRz7TKaDnASe1pTSCymfpflRGjaj
ZJ9Vzw3xYFYYhC/6HnvBgd1dJZG6XXU926MARVCrF5l+LjBahOnOEw37ztgiF1Ar
vSbBcgHbbDd0P4QOr1R4QF6LGWiNcEaS5lv+KqywFuVRKiVrBbE1/+OXBS53vWKb
N9sHiS9U0c8GUf6719wARKaP1hiXCuNiGeNBNhN1wZDq4nUSuNdZhh14Bo7nePea
dtEkA3MJH4AQThqnE34d4Md19xYYNso5+oaG2OJqdQSbyIQlEoCLgesoDUYrjWA0
ml5cOZAInJ0EEvK1X0+EWIYCGkb8KGfwzvNALFmDI3oBSSNBdyR8x8bMyiKIZQIM
lqmuc1AB8n8Zss7pfF24fdMiqyEJ/jOcpUBUgOS+zPYkvHtnORFA2mo1tqWvNDur
c+8W0VKN16vThXw/xHn7IwtGhGsi1mdWLUHLf4HBjZDb0VDzPYi8njJMQUM7v5Ep
Yaqys1X6wA8fs5Rp2yrra2rrMkeiQP8QXn/mVvnAB17HmbUaFJdt40CYHU0rVziW
l/9k5u8jfUjvl3QgA8IVVN49/Xn74d+4BllgYZpxxji/2b8OXdM+/G2bS8vBbDVd
+I9VuoUAM+mxszY61xRN4vznokfsVcmriGTzBqjo+lyfmpy5YLOeXeRo9YQ24uXA
WDx0MlAEBjnTYPhdfO6l/ZStYxV5w06L4sR5TZuiMR7IYYJm07JXeqz9ZOsJrHRW
YrBRENfJTc1xKIyM8OsDXNxxnol9Okl4diMUcfuBbtiZhQV3QKP2mF+N97p46qog
`protect END_PROTECTED
