`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JCn38vG8YzqMW2ooSnpAB/tNdCeav3GKY99RxQBwJVpMSd9QIt4xbPPb7ahnOYVE
nPAwwU+3TKaPEs5omV7UCxRUwlphqA4kvZFNd7WDjy6uiuksqxPMUKXOVKqY1kzz
XHeP/nG3g0Hx4oW7WS8r7/72EjoSBtadY97lFovGS7Lmv6Xg2stIov8gd0s6XyCW
tYJm7QbbQZzIaKxur72H15y6ZRT9dse6ik70UAJJH40OPZVe5k2MNu3vyvb8ZRur
znT7t8OecNI4kI+W590VE1fSDG8S4M+vgGMY7XDKD7UVzC9g9dqBK3Oj0efAibUC
/yfH4sLNVo2bXF69JwTkCCF83fGme+jeJ7ZFU3pRapEBmRl+mZN+xLg5168z6BJG
uzJuEN1A+U67caStVfxifOvqgBSJYVqmj++PimHHUsSbMwQo1dE0kAYYIl2s7ig6
IR25wt/4/mg+ijK3fN9XR+41lLltZOnUchOAI8o4/okdCcAjorQiopCeoyylKHD9
rcO1lor1Xlan7Tscflqg/GUZ2YQmJksLd11Y7PWQaluUGEKifXHyMc9ZKsqs5Va9
nz5HuoRUacBtyEEPbRV+ww==
`protect END_PROTECTED
