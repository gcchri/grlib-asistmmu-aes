`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1RE0ggIcKUWt2U794zJQc/VV4BPMevpUyygYujrMtY3QfXYhWxK6phVG7du8Muoq
dGarSzKUD5x6KzEIpbkKhJvDiZv0Qi3n6FjF4ZPTAysxMYeY+dsP2pSYDihS+tDP
kZm1jO9oCgQDbt+Mr+TESTt9rs6/+JhT+lPC6k3zG+aii1Nj1vZwPpm0O7aJjFEt
wHA5cpeqA0tUoxOmZNcnkd4BTtsZ9BSPdCWgVcl/UyM5b6EVXareKT9rnswjZfNr
2GIik9HhpVAVuKy00P7PEsrusupMlXxfSFZP5bK30nUzlLMMvk8+SYhBoUJiaJ/K
6gv1G1dUGpIXPDM/MHWYLIitm8r1cA1ADi+AmSokXDh7hTcGy/1dyAAoIWj/p7u9
JD0W6cXlEdnNEcv4e9J4qdDRp1hr+UWh6h7c9AfzftABeGvfDCBGk2dQqxum92u4
voXqCXBZ4c77XEVvTXGDmDAQDGbqQYX3EJrtV0jCaavdkiSlZzOmz7OVnDjKVmMN
k1Kp2QfH662bt6aqsk+9k+/A4v9aVNOnmUlKjikohFBy2SwCjAtCFUVsb5Fg2O/D
cfWQ9LmKkxoTHRke65kfuhNt+60YVZ0N6G9b4bDa/NHwJlYmVLJwA6+YiwUc+8bI
BUKtyqE2+0ZGnqWvAjnvC8k3xr0aoatdnFiOelSXUYxJL0LLDzXoGBpTIZr1WTAf
O/8pWKC+BXKOgXsKxBEUxfHQFU2kJK69obm7EDES/4gWcK+8ISkWoJFWGpNSigam
4OoU5GnFJo7MSxPpTCL92SN/L69PcHBpmpMqz2gUcWh2yfqqX1qXv2+w+/Z6wt7I
un7Ubhh8tW9RBvXcCghX3EumKZxjS3qgsqK/G7DrPDjSqwivHvtqEMjYi6tWZC0B
S5PWsLVAmHNBQhN1sETGGmmyos3aK5ifz+538CTmmUI=
`protect END_PROTECTED
