`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rowD4geqxCCiejrZoMLZJ1/+nCjUwSQrxq6YrttVWFgA8G06xSIRwpIJZ+IBiTVO
wxJNvs9eHamouLvf+pOOQdZBBllE/hO+SKua2AFMcTra/uo8j0iqA/KCSwrU6s2t
9paCUiu6FF6cy8Eq6jb/y5loLuxlZPYQSXCEjLp+IbysYej8wkbMxTQeLf10L5Rw
NBIQqeqvj0kEIadykVlSsNU/GQx64xPwQci7A8CXAmf47XgDAeSAGFmuQb658nra
qqo18oNRYpptD5dCK0NdqaFodkVyfXnJQBFXeUvJXifEAx9+8EfMF8oNzP3j0a4H
Zn4ODThRISGYAWBZFka+d2NfXpha3psBET5ty4KQtbkuaAjRnkvSqCTD7Ojsi6n9
y/IPdqyxUnKoQiMK0r0s9w==
`protect END_PROTECTED
