`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PAPkkVz/nj6LCnxDAmPu+wk8nyaegy+8AIIRkqZemZsYQftoK9g2jQ9zlImoEZLh
cf+hSDvsnfSUH/QDYj1TLwQa1B0nJMbKrXG7Pq+94IM3iCVnCa1IpCEb1V/osjT6
9Es8jPekAcE1v5SrTUhQIhqDtpkSmFq/ziGJfYIWLlX6nmDdrAecPFqFc539J/MQ
05CQ63aykiQIAa/eDz1jyl5DleJ8U+jMA/WjOMnzOjwhinSNCn8BWnQZB+I/XWmX
MVSTHCj7NPLIxI8Uyl7b5qCBf7fob0pCY0KLvvAoKsmLL3IxhTnZT6oL3lNePe41
lTwlQYO+YwNmUcGvNT/iaw==
`protect END_PROTECTED
