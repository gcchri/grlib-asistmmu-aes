`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cZfDQKsl7P+zP3WpuFVZz+quvsMH6SffvM0TGgM86k/IK73+hsJmByHlOpqMBJlb
B0a6SB5LpfN53EnZKA7btLx91v+DP8Yir8JIWhlK+Z2Z7+tUPB+X8JLHDGhNvJYg
2eifaIyR0L1llyewpQ0jxDpBh+s8QyqplVmjT3Bz49VpM+CgjrgO7hV8svBXaEnY
UzgYtBsFdr9IkUJ6W5Ek9HxmKeJV1YsMspMEF85dQvaXmFNE3HyLJUUMkggMTz9N
shWtcUGjYSV3wUTcnOPykTdeu3IJO00ziwt/z0kON44vOxNkwd5qHRk7jaT8d0eG
0ok/EdoU+olYNWTY+//vgSwbS25LMts6a54AYIj8K0PjETAmoCQ4t2W+TsSPpqKX
OTs/QU7BWBNWixkOjLJC2G+EAmA0Lg9yAO/ZKOGrv7Q=
`protect END_PROTECTED
