`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/n99pV4XbF4VAwNQI8uqm+ocjyN60XpkjtYwJkcIqX2fdjXArTQYs/Z+oQj/xIrY
PgO47dGgHBPiC7vP2/RFovhDTtt8N/PBVw5t7OCp2Fse4NDCtZRKko+dgO1gYPbU
QVyPREhAXSgbv5eBz0OD8b5a2Mj0Ul1QDQniz7tplkCdtkudBlg9TJV6mx50vThC
cTFzPw71ZvdqSYAkKvV/gj6ulRD2qCBkWV/dJGZxoYyrLIKeQMtSwUK94mgbVsfU
w9nGkiwHs7LrHAPocCBTDNMc8tOt1UpYTx0mjorhj/QnrGsRDoXRLqyzqnOA5gSq
OM0ygUVfa17y7gFKvZIkIN/sVayPEIqfKzMDaH9V04Oe3N99yU/9HivyHNEMpOfA
lP4G8r5sJCr11Uvxe918TZB48dofVpXZd6UrXLITNcRFAaUGGU6VBlbRjxw7G40x
`protect END_PROTECTED
