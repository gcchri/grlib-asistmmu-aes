`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p4rTuCa/vF+Ej1gsXeApKlA3+iHcx+P9v0gmDPvGSAkTjSx1yLLKHRWVS1bzKpKq
CIdhWAjtmhZj9xEmhAQ8Q8E/XjTID20b5EDmZ0VZ8Zq5M2GgIQp/ygWgKA8XqLzm
xVfoEVCJ2oCDLShCrhA0KllMNBVcfVJMAeHYJ4rJzIdzFPmRy49G5XmGzMpMaBEJ
Z7PB+6aiYKg6DZ6Nt7mb4DXBLlQ1uXAqL1pUM5SzCK70GciYZjUlf3Rr3Yd8ehgK
H3+ON8AKop6MX13Yjj7Oihb1HNeDB1lGiS5/PtQ6DPM=
`protect END_PROTECTED
