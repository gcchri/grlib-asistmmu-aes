`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
20Z6SHM6gvTN5gF/LQFnvoRsoGLUr/tDeVWpgQqDLaQEeYmRsF35r8YtE0z0uJgP
Wp4FkAMh4ccwtrOpeHP3HNqSgXnGMpMBvY00zNvjSNebXrRCVCcQxfbQqiIx2yqM
pRpjJX0lDVW2eMF+wKhnTtt6QCrY7cDJUhZB0iyVtJiNMEALelTKdpNqOoMPUXRJ
TucWLm2j+bUKMZDzy/0fnS84MuFZTJc9dvWMKhU56flOqlUuZiYFEA8b2o5eXYz9
e6HSnFelzbXMEuAt99n4Irgobdo8UkGWMTJE/SzNonc60StdgjIsqdlcks6NV3D5
8JBlBV/NSasNTIT3fIv+i3fmuAGszHEnx8HMj/hLfs1aoOs6UDy3tD4briEhwUOb
wLD/SfH7OJpgXUD2rGE+bt1c6ORoLsQZtIv4Onms2xYMKGNukM/sMEqgNodJTXWi
6d9XdmAFyj1R9o4x4wWbej28WdwNM6gqYS3FDzjbcdBpgI4ZMdSHiVjlx/3QExB0
nYspSOfTB0XkZMAseDSBh6Y30G83LuQTB78zmqDwnz+vmz8jphY8tt4MUZPeBgTU
Q6OJ8fjPA4IuGSShIMZBqAXbzjxL0fcZ6O3wZhraUr8dur6J+jXcx8PmNF4LH5zY
i1wUHaeNSy4Ssdtvw4FPkA==
`protect END_PROTECTED
