`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p+tPugICVpMHf9QK/s1BFvYEuf6DcMnSfDjYY0YIbtqP4+80gb7o/Rp+gUwv1paC
XsutNdXej33ZRb7khgjijbFfk0dp5CifSnA4tdiNrY8a9ZKYc57p52GR46+xI+FO
ns74cMs/Wp9p5BPyIv/BYCGbIyijrhlKPBkNHQH/pzqNw6M3X/XwqEF0mZTmxLVt
xP7+h1C+8wNkqZJZnSiDZuvOCqoQeifba/jqQI8Za6axbI5/M2QjNgRm2PS+FwxM
l+gH5TBORv9EIUdvx6tH1e5Pj89P+LH0i35Q4jCr6LQ=
`protect END_PROTECTED
