`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qyj9mZHio1QQn7w4YshG0XRdEijO0dm943LBjGaontporJ+AjxTxxAHvH9WdEh/t
gzt2u2jQlGNhreFYwpIg8/hCWSTZ1HBSClMq6+njuP2zl5QlzsDZ8ulkG1xrjirN
EwmKDD7YLCgTc9h+dJG7SwoHr9nJh+Du7t+2hbUqV3IC/WRSO7HwFx4duEfpk1Ed
texbwubPhanFtQAaV6Cw+RoHZ3AxAJuprhaDrUc+ygKwaOk/YZ9VDUKJhnwtBGQn
p5eowOeUJAWOZXvo5voOQOgz6+LshAasiMd5DUO60PHLFu1H9ajDS7PYhhlFJvIr
V43UauDI8kC6x8EgNu/uKD+pGp7X5W03QcgymtjX4xgPpOVjBeEo/xfD2qlfuRyw
N6Xr0aHh/ZIqkgF74VXdwftdE///k10XieMpENmWYkyZXVW7bMzwQx7gnD7FjbTe
WHY47FbUO6m/y2J4+M057axY7EJlmoc84LoUFZuyWjaVzSwpqA37y6/FaIYTG+33
csf7HyjjHe35mDnZomk0F/9S14o7AQTirFyj7qRoqs3uxgc9Me4BATQCICbP+kmL
rMb4LKJGUaUtFoGm3crYex8mruU9hPMAkuSG6cFIDLjLLZXjv87tCYwMd4sN+SZa
Rgg1uomh8kPperid4I9A54S5FgVc+U3bAOCr3EB3tHtfLWm43MV8sv8uwfixgyND
gdaMuQDHJF67LlYXWKph7IGpuxTXB9H79kAXwLjGx/ef+VXfCCRLs5TxEfBlyNv3
oyFHCy3QTtn6VGZM11TjPS1PEyu48ZJ4p4vcQyDwNwDxuygKWsr7KNphyDLq74pg
RNljNY/aXf/Q6aUAwoTegoet7Q1FdI93SGAbsULzt1+T/2QX1RNbBxISLPYYwPZS
9MXwMn2uEaiu3JC5Tye7nakc6WKqM0/3XHzomFtgbxydEEQ0UkeVMCaNX/oCZQ63
yCipgfovrvvwfLxb37CWPUpGUwLft+M6tOFY+xGZKks=
`protect END_PROTECTED
