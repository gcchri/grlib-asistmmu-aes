`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VFWYZsaaXcnRVlw/qkYZ03om8ESwZC+WD8EqAqbE55rPcm52zi9nEbx4rFgHAmeu
QJ9v8hcLjVT8EJTkkJfuNnLqbd7+Dx/aAvkWxDLNA5ZbLpXs8oTEOlcZ3EglwIjp
dNibswTPFIR25zTGRu1BUxlHkDcw0314mh4+tEn9esB7FiQ8oymR73UjSzLJQxey
cmQleq1Uw5tdIPuMyhCdIwkxr3HdoH4RTgLNm7ipmpKga5J2w58ODrn6dXobGioV
2U16dvp4vhsm/6V2F6vPCIsPhwqqCLsTWfI6c7k7jAyK9fzZf6Ctu+reo/3MG6jC
IfcufmjPQbh+uR6erfEiXy+cUhhFebvS2ZuuKFR9BYkDw3Rodnx30YiYzy3UL5yk
OfdcJjcX4fzj5z1Kuk9Lsw==
`protect END_PROTECTED
