`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YBoLq+eCmuP6prQ5rKe8LKFXr+cBwo52EqC4M6hHF5XBOzRq31CZl34yugFSJOLN
Gi8eB4O/OSTxZttVQZtj/ihnmTc8XzgqOnJ6y4WlggPtkia7BLbzzzxJ3tBLRjDp
rQEux1CiwGTVYZX0BCHc+uxkWGoxNHCQ7dv3PjeLq+AC0twUWUPmSxXN1cKtDxEA
KqR3TxHxE2onu5DjnvhYTmA9twA8cRbOyVuaY/uFLMRnS5UFMmwxpxyKnkTdb++u
KGZ/zk9kxjqdLk0KFXDBF89jbjLnYOV327oSuej1SRC4JBNJXjxb0uRiUzI7sGk9
pnMQBjMfmKKlkPkNPsDOTVO6Uxdwgo+ducDtu7kOE2YZFp8eaSIUxilM5Iu93nqR
aXOcUlOJ3k7RuErHUi9yfr37NyA/UaWYdG3VmhrEzN5P5zFi1LcFoNOre3RrVoie
o4o+kl4Mpi2id6Q00C4814bO3hjAcpwS6hhljxmaNpk=
`protect END_PROTECTED
