`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lrJAdeYwcy5FcLW6VRl6EHXQW+svMZ99vjfdWF9NAYkAu7Hp1GMOXWVaNtFvn0iA
2MtvqWwv7RNOM5ouGpoMeTycZdQP+hcgWbtrCE9VDacqROSsvfYfvmTZAYGO271X
fKUB82YB+cXQry2olrOoPgNScgoy3j2IB1xC4BlDeAFATFu3hZLaFvvjQgWevM7I
M5/A1ToGum8wDRL7SEeocuVkRpBGlEO65d+oIuLkZDbLP9o7XiEPZLio8g3KPMhY
OSf5UPIecdmx56Ey9uRmjD3cnPtMQTvjRaZlXXJEy+sglaoxf+1IJOErlAChpK5L
JvKpub+dUL1MbaFYO4ADMzuSez2Oa4ZDCunHKNw+sadxkVoxvJwcRjL8dVpLbAU0
3yjDRbPYRcvaDadZIf4jTA==
`protect END_PROTECTED
