`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ogmEQ7jDQGG2AZsYZKSMcxrAc8GPW2OT3C3LoZLH5tEL5HEEZpli8u4w9MFxb5xa
SAUNUeVkOJtkv2nkW8lEalOfGfn+wXZkKD6CM7MsRQIfRAwb7Qa8cJ5l7aMpAh+D
B3VkZ+OJSnEsVnmeaYmUdnTUX2p2JWvCq3QdHEMcXo3Yu1W1aqw2Wy8y8NQaWQRO
1Sm6Kz2gFm5gauafx8WEVGX4XwV9BLW3egD25R8ZKKAfz9c3mn1W/nPOGdxEDkvh
1Uek6CgaoM7bnJE77FZN6n226/sX9uIVhM6esJoz2BFDjwTsbGv6HrfN4PA20B9/
D+ZPgTm6rwzQCD4GBa4IMnZaykt/B3UwWgPFmP2FAS3zkbgH9JUW1ChH5f9UScMf
SWwaZCC3vNSMFP36B0QdDdmSGytFkHOkwvWKB7vmdUCW2+4BydnWGtaGwG+2IfWV
mJa8HhQr6FvJs5/5FpfF5kOHVtfG0GwwJbI6VfptxO/ni2Snfeo7wKZdp2+xuKgc
L3JdeTohPrcaLjdkyEnzeO8Xp2FBSiC+ufIZX/nhcLh9TTOlkpsW9/iP4PlXTSNP
tJrY25gAeGg2QxYojD1g+xo2gvWKRXn+QNtshwtjAk15IbAPQ/ly0PUhvi8SczHL
RTGL8/rJyxCcC0sOPMVaYH3Qf8po4jLpZyT9Yi3rdQJSY0CyMr9lNw0Q+iSPj9RF
Y5liqUc109jGfINR2gEFUu4Mqeu2zOoHYGIBciE0oFHSOvFPGomBAOJ4ey8CXX8Y
71nmZTfCSLneWTNioUOhX7jc075koYZCb6/JOkYug6M=
`protect END_PROTECTED
