`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LT6/7hvIChBkzSQc47kLu6SSvqsSwimPMYu5UKjj0VfVDCy1RWHEpgVlq+19Cp2S
ji0P+ha4r9xoFR+d27zdsILRIyL/sYoOg8F2LvBOUdgqhKCaGznnyc71zzJi7fjz
3HjVqzP6IOSpA3F7hERwQ8Fub576JzCq+JRhLfA/b/XvXiqJjWgf0tz8ULGcb11N
0ZDc7z4E2Nc0VyDuf9HCCtKqRaEpXIdkf5xNZ21YczJ3lDT5yJhcoF6q+11SMYKF
P8wOjAsNgrSFsFkoUErkLpOWOtWAyutwWrnFQy+QWfo=
`protect END_PROTECTED
