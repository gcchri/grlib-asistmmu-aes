`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DJtSCDYHcjagt9r/CnzBJ2BwDxtEJmO6p97rrbaBbijTjRi5f/DpTR063tmzqAkK
DBMD6AEQznm4riXScjtctsBqdQMyDAPCGJNC8r9M7We2YAu0n76THIJ+UQzv4G+8
6Ro4D4Pz5yy+faAfKclf5T8WwyzfmeB+sLFTE70t/fGkeA9lApjOz0nBFUZqRsyi
TsDl68JlV8Qf3jgLwbwlG15wwjdWLrhrU8ZJZ91pIPMiJsmh6zTb4F1QcxzwfjwE
nopgAWmvSPFoyafIzWktmnHcr6R/qeWQWgyTvQ26/ZhY9D4VxhvcQbU1npT9SW4s
6xam1Km4pxsxJBz8pIB8KA==
`protect END_PROTECTED
