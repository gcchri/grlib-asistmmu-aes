`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QVPz5tlRRoBDDDI6+jrfWYmmoCeDbr+ehsSyZUVtI4wu1h90MFRZimrwaw8yPRLV
XkC7qAaheirk6VFyB5tktUUWRIcj3532WsNLqocGabtjzoB+rPn0Qk4Bq6qUNJ+v
QMp51zRuVr/wh+KqZT/i0Hh6HAOPlauir0mM492TlQL+u12wKELjhXy9ufZwjRBn
UWUYPlAydfHyp+B7KaOYs1Y+0dO/IU3xvVmmdK4u/lVcLwcTJR7khN1tUWzI8I24
2US8/7vLXQxlP2ctomS4FOczbDW7I67uKw6rMoSwOiASdVf9jFmFTxzY+2izfZc+
7Ud+GRhT0LScmdoJioYZOITMfUmu65RHLKdYpM7EUgsnQAE4Tgliizv+bYuK8OAS
sVmKukhngdYzAduMEU/lVi2ybBayFhiHA82vsubn5Vzfi1NwPEcf5sBkW2VB0oSP
KuGQb1OUDHCFmo66cMZBUqv/XX2lmtDKvM1WyRQsHemA9GrqcCuTlS8d4w6nL1wy
qiE4LT9eglwea/J4d9ml3ESG1wiqvj/JTHwfilqwG0r0rMG7wJpGIETOACHc9kz3
jP6maX4YBToRttePQsTjEUqZH11e0Jez9s6l7uWAz58D0kaeXBd89I3H6AzyNzcQ
S3JuN3HNGmwejzNTj1ko3LLUPQgUknXprxR4twaHQ8A=
`protect END_PROTECTED
