`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QogpYOtQcGO5ncupq4uqcZ8XvgiFToymJInv71GyB6N4sOMkrw8lotVvYDXroqQm
yFQCv3hfygxKbfOheguKQ1CzJPEKC2hKE3IXrIEUY3d5zEi/xwtmHcTYXfXOFQC+
2op+Y7dYHbBkx0GU6JVVrrxda9drO/wYEAvm7/eZNrtVacLj85CgGrhDLghUxV1w
mkjBkOXWDGvuMIkLkwbKOiQYN6e9oqIyiaRDYlJo9VPfGfidq3tUptlp1dL3PbMa
L0gnTmq2esvy3cuptEXjiuIUhic+gfnrbOS4RxmwNt/W7LslBRCfLpjD2HqNb4zu
1L4PoRBfnnAKE7tV2/Xs79kFoBzBkwjWfje4HW5+IvSMndwObX+eHSFc/GKNakTv
ntIGzI0pgjanAejOzvSf2w6QOBst254B9HyHIqC+87fVrr4Okxx4jxt/PxpSX47u
9kBxWh2PICqQ3uyv5eY5hg==
`protect END_PROTECTED
