`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X7BXAR5RAvrSsWObqOpEoDWWR0rZIpgcWG+aWAQehcw2MNJ8994ER9HnysF4xORs
NJckTApbE6PfCXUAainAE5YNWqXer08eiLa9KqyxHFVG2aGchWv55Ehk4rtqaiy0
EaoJkDOwyqniankLIEpoa4XxwJL9kF7Rr7BvdQTfxqEobQUtzDBH5AqzrwlILBKO
S28wk06PalJgELGvah4q5LCb21lajN1g7UdWpUY6HIxPmEA/HJ7PXj/nlicTiyLh
NIVt8rs5CwDrxCMpdqzAeEa06fYC3RbMY9b+0guYQ8LOkoKvZawvIXk/0dXO8Mwy
JxwRaSeKjBfcoJc/lAKVnnh1oxGNEng2at5IAl49rIZajbv+RNCuyIoIzVmxBsNC
E/gJh6yeNoflEoAAgo8gh9Y2qhxjDrn4/QzqDJ8i674=
`protect END_PROTECTED
