`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Np1U/qsStwkqn3m19ffa+UQPwgo8fevR8L8qg805N5oaCiKeBDok8pr7oXt4Efj5
cODmTnHTuIMwyUAfAK9dltTJcu0z1t6cWoqrVw+gXQvtfLeNSZ7vGcWwPZcI2e3F
joxe+2FQXK2k2zSX39ipKQfyS4Yrm859F6DkRDtMYRqaUx1JmoYsTnDMIb9QiKTD
D8T1MnWNnG4/mDT+e80UZcPyNKI/hwXsmsfrrTbyN7AVrSUgfmG/ItlIroMPCnaQ
14o8FlrJQyBYAoW3wbFDwBQ2bta49No0x5oT92uLgepSawHEaaxqYcVRYJ89Lepw
A6jVwTNWsMJ2imXxvr1eHGLSyzs1hOLYaXrZlug5tD3R+uKyJswx742WauBsXkmx
pcKcL/7xdtuEXXYKBt3PqMk2oU0t95A3sFP3QjOVorEXfna39u2AZx9O9VwJZ9n4
6L90Wp1QZ9s8RZMuRW9PiXemLTJkTcTWTU/X8FagtCj857rq1m3IJbAF2QVFzqpQ
Akr4dv4nBPMKYU192CNJ1/xw1EJcDdVg5Ce7lUqqS/quHNsNlU10wuHRNTsdufd8
oxTmJPkRpyGyGk4ULVpZVaGPzFkKuwDuMK5sJcY821plyVcasa0kH9QFSRdavINe
ahFIXTHADqgGX/ZP4m5gHTMlAOFkPtgRknHhx3/uFigMbrxDygnaghibPopl1pwD
ZWVLw/JLGOCTOM/L4WPFRvai0mwVFha7rCgvN9vrAxEubBxZD4ucgwYtP8T1mOqV
4/FmOjr7fPDhZJ9Ww1lDolLdNjynFVxm3z+VVUHK6MWLYk4zom7fpZ5HeuwlCcqj
AjfPZrFnIGdV9V1XpbIWq94l6SWGxuSXtlqldgjW0EJsfWwOU7htWGPaKCgIPui3
v9LvFL86PB3dchW9leOxLsilezB8nI5EWOeki3WRVeax8g8nErDp3ot84l51EQbS
2MAguJ6BOlf7cY3bLznFM4KjsoK+qorIioaTbH4tYXWrZ/fgTp8ONeDfshVIVp6K
HvNcxcE/AnR74w3emVK8N+23PDPiaXibkQVfK7TYgYh6ZtT6oRleibtsOMHexwC4
akiK15Nqno8DSkDBHW6nH3Vg1z+wJwVd0XQJgz5vRf3HyQieMsqQVz4f6hmAcy9x
WZ4wm4gJ3/mtvL9W9Umunqvz1cXg2mNN9yEhMUJ/RiknGt6fnX3eUCiAjWJBRj78
GUCoPR0NA8WpHDeNpMUbHFHcoNbnjQ8pkNMBo9C6fvY=
`protect END_PROTECTED
