`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZGGZBfPlD0iF/awGaPZaDXOBg/sFsUs2EuJPs9slJyASE36y2c42QlDjXFEvXyWa
Dter1aY43CCV0E3tZIWqZKvGrUZeS8TDUgE1LD5FwiGjzvQOPA4yaP8k4tIX7HJS
sVdtpmI1FUp66JlpuOYm1PibFr8f5UeJNystl9tzwcYM6r7LQW3Ot2O0GUBdYLoh
gfhQlBfbd6c1+2AaAQZPeaYJZtBCVxZC33ewcupFWLq7i2tpJIH3i96v4H7mj37W
cQeOVZL1ZW5ztyxGV+Bxd/xcy/8fqCzIsbk6EqvMFF6iQgAm/4ESW6aL0SJoIrlH
hBVC3j32mnXch3VN+4mptgE25VpeHBnfeIqVgvbPth0Rvcnt4xnyHs8/AZo1KYAG
Vu/O4kAuBMGybRU/MJs17G6SLaVYMLEXXnp6qva28oMWKo8SbJDh0O8qRGXSYnlK
FksdMcqq5Jjp4RGnlsy1vyVYGM4J04wK/Tp4Ir02OQaDDbt3D7SXOIIbKciRlWej
RT9M1PX199DkirCrPwu5/BlABNRcq5MMcd2KSziotAwjGClN12G7F8A5d9n5Gw3O
Kcfzzv2P/mW57BGvPnixlOlqfxJFFuzQxXm9pKSJxO9KL4+VEnWE61E58CsrEKD5
Pu5/6N0QN7bmdfguBFhtS+ZYPc+aHwoMxqLU32p8Qn62X9kU1HX3QAC5qclZx1/f
EbN5u80M/RuK9+faO1cr+SPBY2Agbj862Y2QitgCFg6r0cpFM9svnyJOPWusD4zf
4el08oyfD1Ofqm49ZrCmt1pzTe/NoplSj6UZl147TCI00UpQd7x1WU21aitzADSR
arouj/dC73/c1sc/vCDWdVr0CVyboMccEhqO+tg7y9iydZBasqCgBJI+csdEwlEw
UwDaSrmD2QWJ+SOye4WLHYyF7gDuwKSsl2588fI2uucWQLiyO3ip2j6vuKoNRVjd
4YnjnjWvMKcDaAni/fHbyt1RHXK2g4Pv7Vdtt1yvAfCWSgPHkxxZS3vD6sU88aiH
vsbqMmvn51YYw/+zWHgXllCzzFAWim6xIdjJs6hAMbvDkCRqXy/zKKjpSdKvZZcr
ZnbkiNz7kv0cXRvQPlL9U4lhscp2RHKUZZRElndVmhc=
`protect END_PROTECTED
