`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3KMwhZjv3FcVV4g9hcBkTOcgt5a2MZQb9ncIT2jL5sSnZYsu523mbtF/fWmKWwp4
kQ10zTqBhfkbBFrUkX4+2hJhApPau0o6i4Wz+BC5lVz+ndo0/HRdQCd6XykJIL4v
5pn7IYzN7dcRXeMar3Wiozv2cqq2Ro9rB2DVeDSwinCgKCNeJ025CR9KPURUnOsk
TsAqEZyJiZ+GbJ/cLul5K/DDu5EgFnHRCT8cV893uLqZD6zTWd0p7j04N54BWR+h
TR7a4yThtwEiVhsG90KdtlWrZQkhYhkpRqxbKZ+zx/NJ379TmrN+gxY5RHwd+uxu
9XVDiifFgwQ9qEjHavYvWyG5DMAiQJlaPJBZljGIdJFsW0ZpRaFYesMzXajm3oJx
NGWasrV0I4ArMVaOvuaLB7kazZVaZrpa5ak29TY9Ei7YnNUP8MmQyIFLvD+q4EZb
`protect END_PROTECTED
