`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O7XS5fZazhHPcVtnFPzEGSeGsyzrzq8MwcGtV1TPePka6/WOcA9VHsrLGZgWiBT1
hsEe2neajM0xcSAM1wn6tedkA1PcA1NEm8yLZKncfCBHhLCuaddnHZDFe6ESfKC9
jKJuwoBIgik68VjXWw4rvPGLonOubLzwCUpPnFTrm34Sz8O7OvnVRr80aTTbYp2w
WmvPutc9scWANLq3EuvdwTz6Dk7dnOogqI/utcARzCujWahw6DN9UA1uPLofIw+K
pw1CG0DOilMxiXcg+Z5ZGaxT/y8bQ2aluLiXMbV8BXPYDaLDcntaOKRk0ip8hikj
QzVpQxwaT7+OYWusty+iEF3sP2zXhvPCuEV0tL6PQHVp2HwR8MVIPGPWhBods4Pn
1Xs8bnOFzAZH36UDDVR34w==
`protect END_PROTECTED
