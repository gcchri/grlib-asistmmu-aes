`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yoZuVk0Rigubh+p+2xlabS1IGBsY7YschelmIp3cs823COXEDeg2tc9HTW/qkrTl
kjvwq72Etc10HfMMPAfo5V2z5qk9meUsxYn1dqKNgwHBr1WCnvedI2MhgV/XLOkK
NBGMh78vJHuCvpBr0SLqueFzXZhcBTwntYxLZcWjYXo38BJGrznQhCW7r4tblhIM
3lmLMI52ds2wMOyFd7ai89TMeUzKyuoHz2/mxwnCx9q56LbRGUMmr8cJaFUQeVmi
r2/vMEFYBAtWlLl0sc6xeBnURxPk8RPuR3VLSH/3ocGVabh/FMlFSRfymeWHwvKb
CE9IWdyVHury+0CW1SP7cA==
`protect END_PROTECTED
