`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JKgsSBlQXHFsX4YMEeK5M3V9VvYAleHt/ZGytzr8Ul599HxaPLMw/NXXcue5UCks
i0P/VA58xV9VLmkGjg/xaY0C35PvWfcYND/3rWZ0JzklxglbfpiYc1tHm0GMTaFz
tGs68J0klvUPFGDrucLuyO3Pn/9ma8JbRoavyK0tFu4Fo9M+JdsA3QblpItzGitx
jQF/zVsqDFUAvY/dRzcPief3D1+OekU5Y8QCZmYFvhy3AVqS4DMRmnlAWLev8WLo
xrFOJ1YU8qN6Y3a1TJ/+EhLIiAJdZBqcu1u7ZddKyt5ffBin8E/beRsIb95lAnc8
S46nTr1Sdh+n2hVyH3QfDG4OOg1UDK2wQBRm65Y54XtM4rkOffpWdtnIR7/RaRJB
uyvZniY5GX9085HBWJXCLcBkiT6btoOE4W9Liix/xHYfHkax94NfFnbFRyX9DltN
lmhSt5DlaqGOdYsVBdtYuBGmkqClYNtwsmhTkuOnMBB/Z35SbEgOkBj4HbgVuYT7
nR82kvAbXrYjwnhghme4nkPNym6IEuNGVj7Pzo5yA0pOSBrqpucW6vYCg3mArBb/
cBaTZWILJ3epu52HSLRmY6vjgeeM+xGVEqnJCoMjaovvN2AnKVbxLl9Pw6gTQmj1
u+mre+BqBuooJcYtEerVP5mwDgNbh4AkC7uvCBXd5kRh1jkSSO1P0DMmuo6r6Yq4
lLD5iiUZYuqPIqxcKFIxRh04+gXZx4jYdMFMq4TSu5cY9/WXFQPimRmUm2SuRxz7
oacAO56hcIHZt6eA6+ZR+icYj98FdG5am6Q82agwOXXXkb1nLa0y6GFDeHeIELWO
2zgkLmKyUKhgDxmtIg/BcIQyqvKKsNUxx0McEOZeukrxlQT9SFpRHd/ApmnVzpGP
ZdX2/0U7Foo854g9M156zS60hPlZxVH+7EhM9q7FqSV4GC53jY7QuF2RGs3+imB5
lL7dFLZLlMLiSpvq6mQgeoxv30gLd+HFa3EAcXesRIXxkH/XvvIt4awPVQs4Spf2
kA4eElAYxsanw6tUpFRQ1jDVeksXSGKzY5kXDwPeHM1IJChdldth/sljOsXaiyST
NwSMweJOtHz6YPd10jPVvGp3G6yww/0ws8iGZX1YVrToXIOa5EGXA+HcAj/WPyXn
7dvUYJfLL6JEhjLXZbJ+L5ACo++wFImcfw1Ep1FhKuarDrEVnS1dvuiom+X3CQyj
ceYJpUnx2akor3PSSxw1Rwj2foWhQnYn4GaqQKdkJQdipMoNT4pWG7khpkZo4HhM
O4hxkAA++h1fgBusAZpkRZEeYcr5SdxJLW5sWlczvGdiZZUf/72hVXsoB4XxBUx8
JKwyGbItJQ+ayDIUhe1l6xuaAe/QbVzjUA480X4n3putTUX4AhIkobZciUYdVcMN
sVrpcBNPE72luUdF0FSrifyJi/XcTQ7o9/pcgalRi1mLMForKVbw/6nxAaPXed4f
He5uFpZvUHvUR2xlwWkKCJHLWLPznBNPIqIR3WxxADbbHoWvgT4rcYQ1P+I9Hl4S
RuiuNydyaLww75csHnCWd6oyAYE1v6eMdpGZvoMclrZZP+HzOKUgEK0JlRroVz/G
g6H6SC0NvmmEWw5Mo40QsJwgnSex12n/anDcpLugpSbDmx4pIwjgVWBtI1HR2Lme
C2nF15QfnF6HKW0tdSBSsLgGH6kmqVZRrctwy7vrnLbgXKu/H4aEsahlG9NQoUDl
rXxlXpPef7acmIWMi023Df+/beZb8FuHyiYzAWpM1M4zyOjxKTQaCmahvjBM0i2y
M3PdIcafEj5V4tUdy0KI+QAQrIjv/kIC8T8rHG2LBLQaKSUT11O1PIxWnPB3hVzu
6cNSwIH+N+Sc6e3BnZ7fvVpvmnsSaFeOLDQLZNSrtWMHZITC8ZME42CmMkGBApQU
7M010GutqGpJUN5Hqo+AwFLuxrbo37XMRr5n5q3tzHckRd8F3OnYltXChJ/k9/pA
plTf/kdtaGHsRlpgoNwN0VzYIHr24vzTEn2eWH8JHWuQaq/L59KD+Adh+tjmmuwA
jfPqDPaDKF0TfohCJLsQkMf23GprCAONaoc+eQhQwczemi1QmBP352OsiNXP1i7X
ylRiTssq5uziugJsxnaA7fkUYDx3eP0HNJ9ziJvQvwio6IdAz57qnJZJE6ZwPIO+
kENuZ89f52QlqT577vuHz2tWTlm9G4nQ3KDLWVF8fbIITl0LY8zyqq1EUL9WCsqD
6WvWxZToyMX6GvH1tNshU2PfV7N+/0dDFRp5MyvtXInOKWlcWmwUCLUz+lxa6a3c
FhHYpfSDdjMUj4AO0HBKrAuAzMqJHLtycWryJpsPQb32YwEK5TXd7AXI36VWXmmu
RBiWDi36gAXITjApUGGQ3nW4egc2ndDq92wBhTMYKFzvzOYBkFRFRe3gTs2kROOb
7zacOS9n4fhkWk24ZAO/ito+ymRwe+ifwnGVA8OV6avXBYgJ8xRRiA9KQqpPRP34
A0QBp//ji/FUtmItCyv1g/a/bWdZL9g+qouqgEOqOT4ImgBiwmjNzIojLD5ZJnif
V2tEW/kz4fRbso+wl139SkFD6bPRWgVthBT9Tc/5dYA7s/PydG84dAM9+tiA2Zxq
2ljKQkeG/nFJFeuqPaVPqmyqc/x0/rIN/0mnpW2iwBpE5TT1Wmwdzp/y8O7faM7v
TGrX1D/2j9YiH+hw3BEMAbQqKGcyj0fDGlFfscwdSIV41GthmasJNTvxRqzg8oAd
H4fXqcG/+4cHf23ReGBlnjwTreJVSpyUWlDYj5fu4+gt2/c5OV4dZif+zKbJj6Mw
g2Y9djDll5vJYVQ/+kwCr15xwGvWOWecviQwk1v8OJ4eIN6qoUrULLDkqhpCOdLg
czBAdQOogimMNWPrEBPlcg81h6vL/Hpreyr4POOFSNcXzZUXHmlUMc8/nuTc/wh0
ZrY3HT1QsGSEl6Su1NgozZh+9CYGWW9yLGSRY+AmzsVox5+kZ7wD5bwQVEtOPuIK
Knjv7Kc+IwWdbB81vodJpj6X4CH9Zk9xIobLp9IN5eVhEQkezC8IOOfPj2h5UP9o
PBj6sanyibPoCAP5691haxVN/rys99OF7r5ADtXgiUrj3otFsmYdecv5Oiy20/Rz
X+PanNg4RO4qDX+eJKQdFnW0GEb70eqK9cy1hR5ZrM4bw4sYw4iYpTAtkiQx68HE
dId6evnf8Zlb02sJfyLbLUVjHSwc5PWwsmLcy7FfG5pn5yaIITAGZUPOFbe8sk4i
cgXRuUPvoGFtTnNOaAnV+TRW8sFEdoEuFxjjCfM1bqHRkY/o4D1kD7cNdee+pQJ6
6yBXmc95zCLrBtJZaExdQ2Ahm2eR+Us7XzCpYin3aViAEd7s5MnbcBrXSY0Xa7Z8
WX0Ijnypu/z5fG/Y8NacgS1YEXNKJdql4PKZVWP0IKosetgKlorhMvn7tS5uMOLg
Dp3lN3+otB1Jtnc6sMsLo6sSrjNNLlRBwl6g/x6SeDonRpgdorwmz/GbyTtuY4Yp
z2jXvhPDf8N5Bd2hzjoTIg2wvGyiEPdIq/mMpewsyqn2PwBX5ma04jQcE4ak+guL
deikgpkWFqxkji2l5NRStm4WYnSA7Rgog8LJUCwxWQxoUshc4qujkZ+UiVoUD35R
+STUXfZaa4DAvTI9MqOTuJlfs03d1v2y4EHB8UWnEjbMOLK29X+DMHS5iDyMpGyT
caBndjnIFGhky2UWi5W/lw7WpFdr+FWSRfCAkmPUIbSbGRQlMoAVI8FUv0oddcZG
hx6n2gOnT2ntgixCpuWf0DEl8yIw0t7jeq187CbPVkxdCNuo3rZonFHv8/AxtL+m
YkJ1Mj6hOIxNTTX/IhF6NnSjebku0Vu6VhtMp8pINEXK1RQP120jTIsN68ThZppY
aLD6rFMX/A4rzT9vpCOyEIdFDCP4rGc8Fvwcq9+jvrj7Ei2VgmuZnf8K2uyBnUdq
l8BexMJTY8N1PBmYppzcRlBTWb38eeJVIobYafvpRuI1FtpsScqDqCFsOGsIEZDj
HzvUhaWc+q41AqFDJ7m4IKVQPhm8mjVCIfOqVsk2Qu0pfZUI+9QqRxYy2lMIJvDF
1wnkg7jcMXgtsIHD6eyHKeGlxaabEaFcBnmF4UeLqLZ4ZHVpuK/m8uW6eLnQtpzU
qfArwdBRuUtoqhkTPEy0kc62+c0G6wWpJogTS5zdNZYS+Gw6aNFlI0njEymt9w/d
WPBORX93dfTLJliT3RRqkWGTN1miqt7hd6OZYw+9wMdB/U4z4XEAZXwiV4xRx7KO
Q34Xy0fZx8DaDtVSG7PH4AAFyBtFiX4OzQTbCqliFR2fexNXU8FaVgIx2VCBLCbx
6Vua0VrZV+ryWd41dClkqr6ODyb5+hIVmdRHmAHKjiw2LD8giV/f1M78DZS3mZxg
vST1UAZvhuTtZbQfYWb40bJ+B7MBjIkc6Y4Xcg/Qi+mVA7nPl8df5fh0ghC91ThV
HSIbegpwyWX0Q16ibqUipPIhWcNT+CIrK7lzh/J9pD7JSAWCnu1qFLN5eUkutOGC
MUMI433I21tfZY/Q27ZkOdwSiax08+1yD22BykgdqHSCyNvI/4NgKXTv4SBvURL7
GsKizvqr8Yhl/ua6vTH1CsljQdodCPfmWvzzrTgyP3pO9KE+kN9fJ8M67bs0R9lA
vukNhwaKhAocp7iIJ6PKLYJP/na7qAF/zZ1acyF4A6uJaykR3d5TiiG0qpllfuVL
JTjVpoZh4SFkRvEpCDm5fKND5A5SH1zOFkhsUBMtYN8nq6aoK6a06l5PnFgjz916
vH0Rw341kykHzh0bWKb4f9zTmTbhDvXhv4D9oQxrWEkCcgDOmH+67vdoa05fZroN
xLf1+/EkhusGj6vCajJJu+Z4kTuGCsJ9tlIoS4yVaaw1HT88y2CyC9CTW7xBFUFn
VtwCdJ4NeeEg4P1VdfAEfWlexdGZ2I/dxEunDgjdXtT134HoEXWlFF+2Pm1D7ZQl
fxwoE2dqSaJxPy4PCfwLxl22nwHw1ks0W69NmqLsi1QXOywoq03GZUbw78LVm2xa
IIatmVo2nbGiLAk0fS2A7OscfLq4XvX2Wp8CyaPGP3BpAdLO1Hk1xE55McgBC1gf
SABwXn96msJvzMM1rb6eW6cFCU73CcABOElmG5a60MvyBn7NtH22RTECqOTsuz50
V1fZC4+pJVqG0W+Txfzpb7HNEglhgyls8LSLglYvHF3zXW9zTvQaj39H85a3JAwP
ClTkOPT+XTt8zfUlLnRxFrogED49awOuPLMSwCkFpiVO/lcC1yKSJ0JF6+FsJzDd
CrnZN/wTFhz59KREEn0SR4WNr/mDYhlmShN+kLY2eE9W2BK81sxgDx497zjf4frx
KEuVZmkLhxs0QBR0wr54aAK110aCP+lMbV6VjCVY0DtbuO5fJe8KvJKyILjmEXmR
/aWrpFO4fT3UBb27HpnHYpG3vAAmshaeeoa8hJLFyrM+vy4BgZIB05MWTNa9/Ct5
VrKzEV05KJzjUQGmxbxTmfv8q+oBSnXG4bnPifnoD8NeXfaGZqtcaInW0yLeq34k
7qTt9o2Nxnd/txKp/A2CfuYqhRZC984j1E6SQJUZOjl6YbGMCcPX28svOP0akw8A
LJJs/hE5/RK6T7HwBGXiPjElNJLq/5Y3rosgA6MROWW5HxaxgLp5Pc9ILp5bdGOS
94fnFNPaiyeDs5s/KmkSKQ5QK/z2zBu0M2mgp0dGSf8wqPCovvlOB82Y+QXCL/7a
FUn3Ws8OPKJw/a/kkoOGvlPc5tRITglRCPqoY21VWS4faYmTolfLSVAOK8QVgukO
ukRbDyXRMCd+DqzSnnOkvQK6+Go9RjnVlzPdnCtJDb/DEMR5zgYCfQyVbz/4yDzq
3bgjb95sg+cLvcTKMlBqDfpNY3rFOCzP1uc7vhZT9MHHQTneSsBnuwih5I217IJi
fek/txy5R3DutyS68BnVDzMPJPEd/iZHqiz8HvPTBbBIOzHv/cUDhpcFtirdgeRY
MNe/tfZWmfuD9feoe48VXSV6QPEM7sTzpZaC/U9OcxI7Q7Ne14NFAlGalQr2EPti
AwMfBSWrEmAuZvYyVtKu4V3VXwNUKBLJ+rhoEdfSnnI9ARc3qAl3Lfi3V3ZVP9mA
VWEjZe8LgER/0k40M1pSa6gvp+Mm2j+82Wuzta9Sx3LbmGzRilkSY+ttYM0S8qNH
ZsQj3LqBcw/Zr490Qx6lrSkKuJ47tjUQ+oIi9gAgkolg2lAPp5lthQyehNFM3XjF
N9reyMFaXcStvGltQFgjO9q/qsSQyhpGA+XXfg5dT7W2XrMN5Y0kw3lNUq8JWjKH
DSkvunFVevl5aB6HP0GSXHZSD60tzXPZQ6+v+RjEMRd2SKhJrYAfnqvxpHOZ+ldq
k5e//CWljqOafto9ifiF6Zv9E+7RKPtNRFJu764ZksEnLjomfJVqvjB7s+GNiwHE
Avbb/Vnd9Eti+PJPDCYkz8OMqQ1pJsT0IjFCNDEP35ebcgzhl5OAx5fKU+HJLdtd
A21k7cnbvMTIclVfjBsVNe20e1Ddf73JVGSVUhXVZGqj2HKPY3JWT+rImahUoK5I
wQq4JIgzGFSVeCGs3iLYHwNNtLO2ENTkJbHEfS7CTPYGxSAraS9L1l3fI5OKnYtS
S6wHzmo729W8AZ8gioenTPNFxTcTwg3JjlQWJfOBfxBG9yEvZYaEYSxiq5KHu+UW
arBTTriimG2d6nOF2Eu3g5civ+c2XGAFM6hJy9lNEUjBst3LMS2BljRo9BNFct3R
46Z8LAYrTgQnK+ilhiJ+/Y669gLschqugirJDSt8kIJY98wFBgU9yrUW/kHDqwN8
yLOjTMmo7MtvFf6eRmf61htDzsXwFoBd9PWeTYDyn3E+Gi/QEM8mTMgw4dgeD5sW
u2aStIqbQiIuklLgA4agprnYoHxSovPKScBry6IE9FJ74LAVR1l00rdC1LpVr+uw
TcdlISRpY1ZyBD9lMiZBw77qob0IsinEkP5M0HmBsZIhFEJIdrLmXNxcFLX1mhFG
x3amVYnSr1/QTJF5KMZN6KawUz7padsn6fY2k9SRQjsjFpEIHEC2k6wb4tuHsWNr
5ybNrDuMsaXPIag9Z6UAeeY0FFflWSI8cTWaGZod5g7MFiGH251/eanqLQnGT6KH
V5jXrBPp0aWAWwDfx4cBkte2y2UfP1gVWaNMdw3KxgajT4TzO/KF/4ruR6u9WuKe
7RZUMtNmJ93SCN6c4HSVVHHX6NtiFj4Ro1wvTK0bXudL68MMWJS8/yYWxrGm4GdY
sPKQoWnHfi+9kaGaqIFZ7+lAy0RMTsYtG6ZwPYohAmxFxAiEY0dqBgztphsjUmhN
qMqCogcDDU75xFJ4Yq7dK7LvMZIVVwZ+KQLkkSNfgBfwkBy73k50vZEY2YDchIRI
6MviJG05LQPzWMvfcGkZ0JRoI3Lf3LyuFmME8Kt6kkD0wtb9VEYrgme7ZmTsZy3B
cmZND3uZ9vc21LySHEl53ezR6xEmq1JNbPK1wOASLxsD3/6C8MLM4U0LTP7vdoOo
zod8NxvUPxCMmsGaTtB0H6NTXWoGgkEzWDl9IBMDjw0wdghKq9Mwg58YbgUpqfrR
bemS3hhfQPTGphyhVFTh/SKcN/HsCEXZE6aC0pM0LG845SD1GwLbn5srS7ExoBzz
b7JmWWs+uOkX5h8SzEDEQ+3HJfli541/GZuoYQp0z/Q7DdDgube4XVZevIrnhWzf
FFG1ldEj9nCSkuMcOloWQneoy+ykX7EneOi57d0FuhUulLV02nskPWMj6GIER8I8
LsItNEONe/8fIrgUL/OJ6JMuSlodPcswXsJNZoas0KpAUTheq0HX765lkfqlfK3X
5C1uCe7KBr78pAtgHdRgvPFrloaoxvEQ1X8TUjNcC7D5zliGcM3V1BIGIn1WM/U5
LjgqntYK7EVEZqUTDR1UaopTucRGDFQffn1iqZvFivRAuIKidxSP1fTpIKEuwn2+
QC77jAFczkw+OsYwBPYuKUExZMN1SefjgWZQVOhjuhVyWWsb3c0/pO96YugbHpPI
aDxDNdmifnbpBkZS0o7it7BZLXswruYrrCSdZly+lu5a+tEO788XGFcbh5/62nKC
xgoj7h/amY0EzNZ/4ZjvssgsCnv9+RqZN39LJogQSXXDNz4A9XlobvZdk/14aPkA
ip1s4Og7VV+GvUdQlMTEAw5thYrJsuzOk+s/peBDqYsXlSGAZRolsstohe1//ISm
Pj+TVIYXDKdtz29rHM5oVTYITAZe3XM8nH0ecRVTzi7+ybYj6i+tuzSZZEfAbcRI
JJarTi7+mWz0/9PNCL4yigFCswboiPYDtTWdW12qrUqmPU8HBpJhwCexlFy/fQRm
22N8CPBGVt+VMOxG6CaJeDTrB4gNBJD5fZF/7bvsLVNbLoo/qBG64L0rD5jIG49l
pvifRFTZnpXtPN1rAXdO8ERlY4pjipTeAXgMChkOwVlbGv9WVUX6OIy+Im4ydgqA
XzEB8eCsU2nmbzkC3osNo9+8d1/qYEoxkkKIXfspyk/R8Wx6R1Adxo/6mGSnmbSm
9rFs5KBaclAEWiufKF+C0Nk9owbWoH+5Vn+IhmJAI03/wwLCEgNArrV+LeW8Hyxa
CxF5hLMOt3SP+UQeCQqgi9ZOz/ujC9u+tL5TvZUSRMgE0sh0pv31DQHDH49UI5tQ
oYvVC0gjhCowGBJ9nyhzPvW/2XxQo0ncc8SJdHo7zcVZM01TpYuZT4BCjhJVejLU
MQSnL/+OCSxCzkxdmmt6xc84icxOb01wWhRiM7bQR2hvKx858dCa5zM+DWxp0Cmj
mhTAkrxPuQt5MzgNeYviGQ4+HGo/dUGmCP95BinRroLvjTYqyui36QDtzzy7XTwZ
VPyobePW1zA6LKXtuwVRVs9v3lWEHB9SrSFPb+FOm5TKgBA5umQ+TFjk0bsd/Lrg
V0ewgX5qvLhFP7xhGHUz0D04aNmlnpjmBrN9HkAwb2RNuOF7bkhSdpiCLD+VFWV4
gm6zc9Lph5v2sjDDuenxWi1jwyU+UGwqc4PM4gWTYAY4nOvXjGUYqDDH/5JJrGRt
8PyZgSH4LfBGSFjGS/1SXscIlRTqefWpnTxb5iXQ44g6rnYIKt2JID5Pb8+brTdb
5J9LiR7ugSna7AVyXgYoS8KWDjzBuJVcPyZVTmgJ8nU/eksxD385C9IQuKfw2LyE
dLNsS9p+SkkcMbyf6FAOorjDmTv+53bEXUW5OoIKGhuf/Cnlzd/DjH67pO6+vGXw
+DlIk8EvnNhiZX9x2O5LtbSjzWuVEyriU8XULQQ/TZ+1QcxReJBUGBhbLcjtw4oz
rYS8o+DF7PA2S74l+2pm+LRcggYky+gliWLefCVvagrpn9bktmOSe8XcTkXQGi7O
KXcJpvJ1nzZntY5DiH9oZkWO3Zyl6JvQGVH66fNBqlCiU83Iw5vpjbXdIQG+z/MZ
4YHnvlivkTgiVAQJo1y99/BcLHsVuZgfyjfBf7KLC2JXweUSKMVGxueNuGoWDq4h
2CurnJrmPA9uEIiHeVj/aAulSAx0ZWa+hOJAcp7piB192QVcWzC0Vs6Tia2H88v4
6WnoU8JmijLew+h6q7o4sF0BVxI5gZpSjmiOWONRqfc6ls/Hesuul3q26KcIQf1G
g4qUVOmMpSBhjN/P2xzPLhk2gEsBesvtBayj+DftIt9m/s/HgiFdJxCi1iz2lAdu
TE0imaOJn7JgeF7ZHIZBmQ==
`protect END_PROTECTED
