`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lQtBOvevWQA1GBbP0rwcFwSMixDmdVb2+KaKX7EP1JL4ySHKmovDlSZVJhPLCkjl
7vVqJMAuzhuFn/ukVQVFoW/uh8L+ynmKRijcnTt+hgY9RrLLU/tTeC8QXc4TfVw2
gQMw9u/PrcMvHft5ZsWTZ1QzbifEur2whnYUhxwqwiqtQUiPJA8hDSJbS+ZaM1PL
3P4SNEhcFOyJIUO1T854KggtiMQtmH2jUBwWevnOdiN6ad/8Vk1SwWgdMiUojB+M
IM1sWRxf/6mcPrAJUZ5mJt3cKcJRz1/fXQUI56uXw83wB4nADrRbZBINsxBKmUXu
Jeiux5xk3TI0Z702d/kWByPInytaizazeO4FAJo1Go9Ni3oI0T3Oyygz+KuJ77UZ
l1Jupwn/zY7oxXIUfSf07ptEz/3eMnSz/Hdptd8aJuww1+Ad3wJl1rzXsdoyMkyd
qnlnAE0fLNlEVsDxydLY7VeMhZFHISO+PUs6RzZ1Q5nj0sE0wAgN0U+47xTa46X6
pami2G3FiRgtyQ2O69C96xbnnm8+nrWrkPtA3KzKNJkEc0YEsgx0dfixAYkk3Rpb
40/SJV4iU+3AfHp5NkfnfzSGmlaZmtFA+GvI+RsEVPIRFIerimQodkw7h9Nn/T+s
khy0QBk5E8Z5kNVw0mBS1wr16gXR8nh6/y5Mg7lfttUu91C8IucN1AI84C5AjqgQ
F1BZPR/fxuTPU1kiFR3sL3ABGvRWSFXbajBL4FoRJXfT370bzLjR7A+462u15om/
nImLDsdUATuVnitueT1OArzfR1ddQu8JzXGkl89Trv0C6N4+fV4igdr91O7XZpkP
alxctGhm8lu1y1JPuzeW5WrzTwkKrlkHxbJnp4RsPDIGasMKOQn4pFZ+9GHRsJ6d
QxLhDJ4JpoUqH30okibY6D1LbUFZb3s47Ja2IfQ7xfI9UWz3VggGEzk4A+EuD1yf
TjHP7qvCfAvup7VEl1k1fOkeyZHWv5hpHfebX3Yby53BXSHgsSBJJbmYdNS3s/6F
FR7F/ouovL2kGcBSvU4uOOygygg33n8S5yRIT8X5wGINf5r2CK2LnB/U3f6s6b3v
8MK5OiA9nSIuowS0YsZn7wKmAeYQ+mgqSSxgibm7GwD7tSaIMvNmlO1Kb4LOZwR9
yTa0RKqXpTE4tWTcCM4uwJ51wNO7S53qCcSQc+4SO5cYfH/PC1eo38Wkz6uBh8Hq
xh/80qYUEvqDuzwjOFKtWMzaxyXgYNq5ZiRTcEnImY6+6a3Tx93tA/vyp+9nfrrj
LM3HNcAlcmsqGvxt5CxtU3YTc7Vp6FYeOt5+Iq7RsfoIr7cFBJ6/D4umr2LIOvhA
ihowd5aE7A//SRJykC1/BFhHieJQoep3KK2f9RyUtDGlCRRSbJqMhIUm1afqeBZx
KkfaMRPF3n1i7Kyp6ni1hgjbMeYyKFFEc1inkQNkqIdMn5lPjVKg33ogsuN4g4A0
jzlX1USX4B8d2jxNKfnrKQow+V965d3QcP7X939raOQ+OpHAIEJXYTLXrpenBUOY
cmLi8D36NUk2RwS7coPh+dhbf6ZCpW7UEYbZHV26YeRS2eFIfilcVHRw1il0H4tQ
lnQ50QL01emSmBMLttmsLNadSnmeYng2U2KqGpbdTkuVHxP9nLy31qVYSGvWGAi6
5+PWJg6K/DrPYvQ/ejJQMOmN/9qe51yv0m+HG4G2Q4OurwGUUciukcM3pBSIoXxT
icyqRXe040tfha1itLF/dL+4xn8f49Bf5l3mKdq4jWvn3IUOiTlEIaLsf8voik/e
VCxGtSIVMkcFgV9sHM8Qlr6h8DnKFwDwFqPoAheAxgGexAQnoD82PVJtctND/FlS
YrA7A0hNPVd+748RBK38JnjF78acul7my0TiSRcses3m1erlWBfEcL7KBhyDJjQN
2nlCUCd6ekhpv/18rKvq+m6v2/1umobHUg584PngO2j3VTp+JQQ8n9CJcFMXvc10
wk/btH8XPqyt/4Z21U7p5Md/pg2jFPYaCb8N4r5bXJrnlzCJXp8VS5jrTxQeOAKe
Pn6D4npYGfNstOw+hAYXcbps1BPGLmps2KwTqyjK3gNvUP0QGJE6zwPVVENyj03g
p49P3Ax3Jw8zWjUTW/HpDD60Gl9VVj2ULlPN4VIABp732IWmuOsuqtKVZBbWQ6Dh
XseVvPXpKlB5ouq/2vh24jiB4a4QAdZ3nsGcHy/2ryrwOumCcvwiKucedKW2OFrR
CYvtVf3UnsWqoHYe5+6bHjnyAQQvKbEVGtmDx/D69O/dv04vU2xZiOdOriGZpoU8
BU8Jn57G+HUH2QP2tcgFVrtPuDoRjipZjGdZBBjKxvF+i3A+grH1gWhUMVw5/mMK
GT/GDB+wyN/TQDNX8iCG4t/WR/L7OjdNFJNMv6XO1DcoDKQCBg/IdPQQIso5/lNR
47HslaWdh1Wbd7vN4uCgh04TFXFxcZSZPDJ/dM02bRvi4Q3XVl2/xnTtO5PNEy8d
UrdXlurbM6Ke9iEXB2OH+qfYZjJdqcwlyJOxTlq+7MOOstdqkXpAqX1b0Lnj7h5C
uHP0Q4P23lm5CO6Qx1WcN39dM1Agd0mA1AWTuunjvXkDIxCfkdnTtGqS6HHE4ySS
lzB7JoLFphB1t0tieUqNZs3a1iWFj2q7GhqqnIb0dilS6oe5BvBOHwSljASDujWf
HCDgfnPwkCDP2lEt/jUyT7i3WYwxTU3lwd7fdSF6Qjp/YKVFHFqwIWkUVhTVVjXI
y7ZxGmOOgKv0GUt09zMjqqZXfYPNbo8UmcrAgVVb4Lbu7rjdQ0xi3l02vT8CFJxT
t9VrekLuAqO+GVWphKr5rgXpyRT1wQwFIRSn7ji8wkcgz5SwlARDfJUX3bSHIhHH
Dn95+A+W/Ympu58p558NsLD2WwD4RDLKRTB2tpJM8cJezpWxKroEOOHNmpL/UjuW
cr1oEjeRkqw5CLAfIfznnTAihyVFfLbHd+xQ04Qz8H5yEZof3AnK9plhQNXRMg38
pLPKczOh7H8d+rLCL+a4vNKiIuxoUM+Bp4dU8lLQKowfwomiDTx+xZcyCumhKi53
8qHKE6ME/sR3xUQQC1ZCddNDrH9uFaznSDFGYHd8QSwWzC2jHjFFlRndVsfNJ7GM
J+95sKJ8Abn08hj2UlTfvw7Q2Up95wWOWRgfdzrFvRm7wL7cZncq/RrGivvpdo25
kAGpMVY+OZhetkweDOxRVWjnRZyxIjNYGvMf7YD6rjlrLHPbGMBFEVY5XZHU7ONJ
6cFmYzVsvdhALaDDKiAGA3/FpyWo7wzNcjonMSCXL7FYlg5yQUU59zJTZzBeEHft
XBockJL4aOJ6SzUOe5yATSBrAEhnUT+1DvrI38LzhcPxZcy22wCDYw3hyEiNnuc+
yM/Y/+bQF+KmYHz6/zciz+7YqC2jqmxlCKyjAdRzojDxWYLzk4N3gvIlCr/eOyWS
sSimdUuxkgY3w2z7P9ZfkTOhkuHMgIRjkTuy79ukFkJUSTyR/UqRUVpHbirjYaDa
0xAlQCvinAejGoEMHdMR5QQQg/n7qA8sF+P2QZ0ZGrbMguwbu12BBKPjYVLZG3EH
4OMGppnRAmflcMCQG0giCGcqzcG/uYcVqEvB/Wz3E7HhalQ+my1GgDnSsA8/AJ0c
CusRpG35kMKJQEFefLY5j/o0QZmtxN0IYBeo9NXiht6snNCrx8lOCnQR5OzyYHdN
Ze38sJDkKsvg2uBvwCAHAfSJN6fGzRbMmzQQgAOIMSwQjHa0VKSnqWFDQRVCItXX
viB66NSzeyQtuvj38cQARkw37fcXjWCM0ozYANIyDeH6lXbMwthzOHTFg6PH+buS
nWduG6auDAB6O++LUladZbAjMT29vVuDhUpdTeMBNB/LO8xuKXaEo7xcl/WYLF6x
t84iy46uF0w1wkOI3qIAOAvvQHfZWTocZlkr2+2jzlX/jOe2/S7U6jzakwfanU/H
65z7+LKxOMPpMONAwlnKY4+8Z+FNiK6lzHY69vK+6jHPZ/Ssm8tZAbuamk0Rgm3m
45KS4IWsdkAjNCwVwziKwCSGspGOGl3ehft2lc/n/ISP0U8p7eN/lMGLpaSEhVWX
2xV94I4Jx2YU02TkLw08T5huYeuDlmyCpntWxSuUvNF/X+xTHO/toy0SKv4nsZNQ
LxHZK06NT/jnOM00YFV0WDqe0Q/i1yL0scEu4dTYusk4arrEodcpkyyYWYTXx+6h
402yGCiapUVFX8Dpvco5Jz58The3WMqwUvHWLUeuJg08f9xtRUek0Q/iX6U75DTQ
/uGHEAx94mp6GcyRB8rLFxm+qHCz9+Q5rWxxq1upOAK2Wqe1lMT/lMgegwBBQSY5
A4aEb3CUcbBFjzjevQg/1WvTDW94VCASQgWtI9r3oAO1nd97Cwu543hKJWOktkgF
bNncDyQ2CV0UnngkgfGBycD+recnqUqwzB6zT1xyX079vTrvaTzfcEl76MS2TmRK
/lC7M2GTEnDoHORt4t4cblrp7GIbhia9/ZA3yjVs9Zgf8RPjSkfjV3ASVZDeWBjO
9TkWuSYcHIluGqsCQUOMfa1IVDF0mT5d+ZUN8SHPiPJEg4kPwF7XbURibl2zxx/v
VFjop6cA4y8XZjfsFPwBNBrGvM9gXqWbRAFJzNBpCQZN8+OhMvMnMn9phLEVlG9q
DLo7DLQfkTpbKj7f79eEujh7tKFHyBb2PsV/f9O3R6qFYWEOhCSX00rwaOCBVhWT
F57YPvB/Mi7QtmI3T9iWKMOGMGvQ8vNABV4NFQQXG84inNzR+F9c16xzM+qIU9Gh
fEDROwkRGGngmxNHoBAYp53o7dcwXF9i0G0wwWCdACNUyh96MosUn0PJWwPjXewX
fxszdV6dtFVEQGelpfh8fNc+lVkZOLUrDNEsi9tW7ZYMTqSjQvCcAqYG8qTA8oku
IInY7eXq6qHLgAUbJBa5J8T+6fQtBA66HgSkK9SG5VCVNscRgAAf3MuLUBudAC7Q
vUhLwNGDabEdC2UhBa2tf8e2/LYwXNk0AsfzZn/ZyvYm0zsBRLkDoLz07UwRIsxp
GVl2X3LApFAtl565cq2a8nUWTSxPnVX63gjQfJeQLslGzhosE2dSiO9pmcfguxYm
zryUQmKdLiU3qw0un3m5B/w4RDvGBZ5H3YQNSBLKbbfMUnNXshrRvVcNgU3Mi4sA
5cjfyLeE/tvmdwZEdmXYnUkHWNGCvhNTKuKaJNOjT9GYAEAt9nUF9ki17DA/VrI7
rTRQplAk0nMH0e+ziHGoMRzmdHZSaTJBY/ExXKJTFptSGyci7KohXnx82RkZ/uJT
THWmGJ3oQAPaA2RX4JJhFztYpMd2tvwPdu/xbIt+GO2LOOI0ML2mMsYBQUPE0Gq+
zUmSm9443pnNZE6qWhIg+AViqdCzGVmocNr+48OdJwllsZAIOn9WznedYlocwjQS
z+c/KmZ1iwjZizv2RXbm9CgSM1qGy7eTSppx0p3xg/pQ8ZLelmwh/DH7wAmMcvHf
jQ2OaEI1p3kwVXiuw7Y3kkypunRZRf9nWn68AZMMgGLzc5vAlQaqbelmxP/jdmFn
dlCDpPCeZGfWKGoW0MdXud6yUlFMgZUAlzIa46+lqgLg/H0xnDtTjbz7HNlKcV4K
sOK1SC1AIGnBLxaaZW9f3leZvLBAFnxev2ximpIXgSZZrZGUDmiGA9Nw9/nWdGsm
IdpmrO2t5tVRto6bcwrk0skVT8eA9Z3ZwaZZGpm6KMQyzuvrt1/sgVItPut/36S+
x6lFG5qDMg1j93Y8q1XvA0TMy+rKME/ktHMeacpY/GS/OK2Nzs4EW42JM6F+2gFO
MnjE8MP1TiDEnt6UW/0sCUzCjUmEU/fEnbt6NoBOn1EUx9DFkLBfoMYznSrkYihR
nqi9IGRviApbFRYhi6Uoec7k2hg3IylNWK0ItRrGL+uusFz3ZEkRcCffmJkux2nb
2kQ8IwzEgW4yJBcLs6x8jUbii6zZpBc7LQacFnFhx8aQYb0v7/LZdtuhuiioKCmD
fuAWdCimemYtoE1ULKxiYQ2Bv6uCs8AtcmAb4SCH+lylcfMuBEGG9n0y+trdCjPg
TeEt13hwqi8TTVCJq/DD2BGKaVykwyCXLaV1N7WdhWq4so612gyKfH6Eg3hHVLTj
cih94wJ7a6EeEXRfZy9mk3DZrx9gt8h4qCyTE2IBY/fglyso0eIO3N3r5wA1ynuD
jn0kKijtdu6A2YNHbVdyvgoEwLtdbLgPxXC8jDDUcMt6otQHhFgwq45iI/o53b/1
0mFeYwEjjltfr2a0m0IVGcFzvGjF1d94zeP0/+R4UsCTIjDKFOin3vsuWqpTd2lr
z9tqiQ/IQwRhnNqdyvAfU7dZoeZxD1PWHt2cj6uzu8uKfSiWt4YNR11espyRxgey
uro6rbHOJ0VavnVT5gT2h+ZRH91E9HCMX+UF3CzcmsnUTN9qB9vhOEyQtCWBvGbk
R53oS7YL5/4D4JrMFG8HN0UgJOU2nuIqCVmLJthUZNGZPn74lhwwAZHJkM3zoiWN
cy3uBBjI6TUqoyjRJKWl7e+hYNU2ErDsedXnCAdNbkzcRcYqKWkb6sWYutMJVvt4
A+G+QQUjeCdTL43C377ORfytmaxYLfXujU7rzUPMWUBDbYi2hTJjOj6wCSHIJHs7
4Q57+lODQcN9c9BnSl3Tv+1ATSHgnvn4nVqRXrkgSJO8THg55ulMqlHwVOHISJqj
RvyIpaddA8XjDCuMNnaWDl3rT017HnzivVCAtahO0P1oiiAQ2SwFbCSKGc5axSBI
suTW3uCM6CjFvko62KfSGPznJTzatb6Cd1xHJs+4DBolxRyK9FzwCTDzxQIfdy4W
zU0qVlHAdEyRkfggpQ+v8Vrs4h8mCwQfA32ONmqmSI8uCTf/MKA1iFTkzbiH7IF/
o3Epv0zYGtwUrEM7VxOVFiSL9aw1RvF/Df+XKZhWzX4ueVpFa+mSC/SaJ94meF3A
bqYwqrBgVQE5GQsPT/Q0whi68koeuE8pTjYiPugmRl0e2KBfQH2+FS+iS3RBWEhA
RuHe2ejhZsGoUqDBUrzCi40iFGo4itgFd6VH55B42NbVqUerfkObN0QKRW+S3Y13
70TFMSaU3ETlOg3CRsPjerdu1GFbmOXpWY2abw2kqVAzz+SGvqC+rKuADyBnSqVR
lamaB8sVM8vreKgYXen2coTollOgjWf0QfRUYVRYqrjmSm5og5Y7LEF5WPTJ0NsE
8N2389gfGCYEG712q1bQjAC7TPddxpryYjca+x5nYhmdbN27a22b1tAoiqaAOI2z
O7YsETb0Co364R7gN8f0ebnFHnfa/a2f2M4u2f+M0t4lFXWgqtrPtjdKU5T38vTC
64v6C85sIoGe1RzmFPSyjQhGY+XV2dGonzJpRFbaq6x9VImfc06aRi6Qsuh18IB0
S9GORGzt1Ku/fVAEwK5NIJ39f/sg5YphP/Re/Bh4+b6ZJdfLFPoujLJ6S0Jw0kGc
/AmuG5X/qCBOUGszVpxlz4EAsUeKsoCwk+OwLTLhoZRrFs5FFxYAOykNzUzyyoRD
8m2UQbQnuf3+b+PdMuKa3+jZBmTqueMzIb2H6BSX70Z8zhLc2gYVcx8VBEDgfuXa
9gUej9gT9+B51oq1lZK52ngR8/1jeE30AAGDsE0GoM1ABzKXVnPzrq+Mn3S/ERc1
K6w0fBX72nWB5sJyC4encQWIxlQB+axABNxWuPzNnv8YpaMWYpnD7YD1TtMKRgi7
DPgt6oV+zJfbnrdqEZp22e02q9UQ8CimP5azFU/B9HZIt9he6gxIg/pJJK4qQm44
W2XKvsdhl46sRQoXg7k8acz4P69TsqV4mMcT1fW765i1UqX+ZJ0HwbgMKEhX9rel
yQeprdt7LomXWbah+rFBUcdtPj2m3lu0olpR3bOMcflDMobgngLESm671OKQuNJU
sJqKRLe8K6K8GcJBGx6K7immCt2NyXANhUhSacRbw3fGUVSPKePaip+dxvXt1hF8
XASYBM3N9BDK3twrpiZMHaaktlVQ2estsokkr0fn4aTH8O5Yfrc13Cd9/jFUBDWz
GlJUE7IXBpYhw9C+gYV/H0YGA30MQXy7betdSD5LYQj2A2L7tUzxthVlxhTOHhbd
/D3ZAYVf4TRXI6SR//yRMKd1IdgyVcQcm7eC6Ls/tMpvnv2Y34Pyd3KbjNzaEVWr
qM4ibHU5PgbTXMrEp/eeKuwfHmAwOupDPyFIiEtwX/evJmJYZxqVe/JudXR7bOau
xVxXuE5ZyOeqNv3rmpkSFnuk758q5SofT72ALu/knsTfk1p++rmTSKc8epF5HCfo
EP4TLMPoIvaBEsD3cOqMTPl3eJkkhF0gUagnoqWK9lXC+9GnlwyXZZuen7HJ1GXZ
1NXqXdmcCfmWwnETaYpBdJqE6oP6IKNTSqBmbY3pQEXVlMGaccqyqSb+lra9XVJb
g3XpVlf6DOrrYimvRC4yMkoX8rB6ksnz0/dNo/VdM9cLxpxa+aPw6SfTo4iwwd3/
3hthuyQZB28iDF1wwtL7FF1C+YWHsCK6whov6xDyVO2BVIM2T7j2/zyGsAR713Qb
gFO8+pFyB8Ch6287wtnwp6dao8y16s6WiMKvX2NzyyCTCkFwTlHpxQjPCucKL5+g
0revWI3S8AQSa2+6vz7r55Z2McXNrqQltuGpUM4KSxUYnfH1ydAUBrKoq9+skdZh
3ICtaF2zT0vPC/mqy0qTX7ZlR9XJkTY+Dh/sNaHI2J2edXootAV98/T5vsdfLeNa
2DO6A+sOW7AAzb3eqD+eGkwBAwIu5ZVvg2uNYhIi139Suxgez4V3Rgz/abcuC67t
xLxcaszmuE9fklS5bvC6WyaYtN5fm7IysnjlQULEUD5o7JrLzMJ7UsCzrce3OX68
`protect END_PROTECTED
