`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rpz9oOfB3y8q/iQ2Quz220mj+v9vcGv0h7tLdn+laUD/0TdL8u9xPEEI5VKIWKB/
ciqpOxpfKiJq7/ZGRq41Ss3qD0BU5zK/g5X0IuGoG9N3uhb/uV4Lx4VSqq7zQhBS
s5VCb0o/61D19V6ldowCR9S8nccqbfzgzwL3bkTWH7c9WSOkKUs31v2hcMf062Xa
+sO3HIHqPdxW+2bQTtaf/OpCn9KHKHkAWLAWs2hzlaDwNXL8ufprLkkos0pWBazK
RLXWvxMhxnJsorJCOBILKZ8ExfdONo8aS6UNVXax3weIunUwQxHb1vzy9rh2tY0R
9Kge6CDBW45+o0DPWNlNsKEmcfNC8OTuKl+7Hd45Il5IAYs04DXWn+Gf8kRYuCl1
IzMqT04BibSjgxAMeYppQ8IBuX6DpRsqh1wKiC3vqUFJLSG0cOztayDs575i2Let
HTYjAalfUAEgIubECJVgkJov/8WItR880Ma2wDM8BKy3vP3FvHgNVP9WPYPtJXqZ
fYoQhuPI0keAiBzNkJh1sy154glU2c4bPD4UpVTEkhhODIyzWAvgtkm3XbcTsgEc
m4EcSNC6FDfDW9r84QsUI8A1kJD9K8TSzA3P5iTQiscUBlxAC8bUV8mdWJSWAihv
`protect END_PROTECTED
