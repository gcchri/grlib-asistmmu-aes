`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/vUOWEP4+xOsJCzr/titbMG6UAGEHn6e/tSm5mmabFBykMh9PwfGaYcf5EIHA93Z
KDVXrvwPKFJ/DxHtfPoWMTsDZnkXCiqKuPYYvmTiTYu7eJIylDV8VbNuLV6UgaPJ
API37NjoQ5hlznlxkqyMeX4IOEANMFnGsM3kG9Qu6eJXyKfHjTO2c50FzP17vnN1
Y8vA/WuH4PqOAhROpV/k4xD7spqDcKIOOimpuhuaPEixMpHrOEx9835g5NIw8rXW
RHCGQ0NIRlmGdzowefqRzjZ30yTP9wWtFoEXLp8z91dQCiDWI1bWCU5Vu542Rxns
hXTtTBnWFrTu9Ve3ful/wMSOk+qzZAhtX/K3E2/oUv+yZGsxe3+lQ7fI+2s2ED1L
LlyHQwtLujESi/zuLoxvqpg/axUfaZn4kBIknyhfmR5ly26IdXEoLGCUMZKOfRO7
`protect END_PROTECTED
