`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GVZr9rcLCHIzPm6FpzmBRGhO+kxTeHa50q7wLb+qx6CXHMPrlGxZK8OgD1Mw6xYW
DDrFo4sYdG1Gk8oi3rvEfA5betHxxBgsHQ9VlvQLYgjsy/eKr1SfDZFPoQv1ChlA
lX0jWM0jF+c1PRUAXqv5y8Po2XGcg4qXj2RZ6vw/9OCW7OO4qvrnAKTRMNNDIVKZ
PXvATsoq1anCcBkROs9BFYhEnJQgZ6pvWJK2ALhjomDaRz+c7Ju2CxB9EokBGEPf
Lu+nfYbLD18ON0h+qLNZwT6a7xyVvVrIGgCo/aQQ8psgfPCrLQMVvlL0dJsToesO
VZd+raopk/g1x2Ir1vt/EPp+fUM9aMt8K9vL0ZR6MZBVvbknUJlxSvGG3a+3pteJ
kYsko1S5LWCuiSQXAUHqI0O9Cd5dVzRm4BAkokw8H/qb1prEnOEiZsqzELVzHqvf
ckPj9DQ88MO/p//l49oUAklbtI/1PW7t+74GMb1kzijEelaoWvjm2o50LGvXZmyP
xwYaX/YXETnVGvqctS0Cmm6bl6E9pB1m/NJw4QUZQ9i9uYDwrI1Vd4Gy7rfMUdIn
QqmErdBzlpGnptRKlgnpoYc2HsXlL9H/cCn8O25lSzg=
`protect END_PROTECTED
