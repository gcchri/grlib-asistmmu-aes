`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CEtSyB1nj++o9V+opFFA3bdwgxsNBqMCt5W9ki10qHxdLdmm/7lSd7t0GYqNAWgh
oXGFM0WtRG5amxOek88AaC6NIiWyh5j/nOOPsaBori5xgRQbbOmx9Eei3yoCZqbu
naCegi+RFRYQzfkK7zn3n3YtqAR1hH8yNKVgKpug2g83fP9XWUiTMz1/nCNQm3Qz
m3q5JDSYHKZyBlrIDw8C+mhkSl/8i9/sq4IcPe7CRrkbSxT93zCvY1AmZNNXk/UG
ppXmv1l7aoqB6w85ETjq8lDXxfryaXMCjtitydby8/c=
`protect END_PROTECTED
