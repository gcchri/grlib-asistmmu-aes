`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tVLVhnTa75QDhoChFnI3PDFjvXsRWoVPPwDss/ly+6zOevlYrc1TwfQIoPSRAzAx
x2QJT0zE++77nXpcx1xA6Q3f9s9soeO7XwcLE/WDYHkmJWZ5okN3mst4Ar2ESzcD
wFQHh5p7BQ+lrT6CodQXZSavf5GyWvKU6cQOXDFPOCGJH6/p4TntgkePOQc85FNW
8uvnHYjH3J/JRnuWGoh04xyZEw8b/KYVKZ0JCb9yJpxOX1pD39rCJPRGjuQGqScf
fUeq6730JnDqky5GRLtGTZ1omLp3ipYbEgFd9xsBBXeDrdd2TpkMH+Fd0RgsypQl
`protect END_PROTECTED
