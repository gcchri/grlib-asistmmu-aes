`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KQKUjmXjJQ44jdDwV6TyIqV/f6qoh2zqAsSvDVLGAMLCJgZoyRqgLXded9zzConT
RldzoeR8W7MoJ51HITvqfuKoVUCD6WRNjZ/GQfboUUCaYDOdL9NBGF6iwC6W9GXQ
+9BvAqdxVcBRuUz/jwbtZuHqPfWupIQrMFrsmkN8WE7dY+wuJyCS3zQiXp6GwZi1
iZJ791RSdWvoW3HKtHUZyPSPfAI2ZMBfoFK+GFN4M8mBQ3Vz9F22O/3SWhthGbPa
PX738hGPCdzfEQb91q+XehXrTQp5H2gxuPKWEKbWuvHxIQv7oYmACkZY0MUQjz8P
IDKXvO4kBoKxzmy/JIj+UizpzTx/S5Kd4LnwcOSJeds=
`protect END_PROTECTED
