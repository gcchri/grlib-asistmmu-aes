`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QPZ9gNJkex5HcPYkbUNTvSZV9xZetImUvJDB5hYGtcpVF0d2LRcNmJWoRBxYU52l
59yy0aiaMRQ95s/D92QFRs3smG190nj9mcSVVmNy65Ki12Oc88w+LO5xTGtlINsl
1BJdzAsmOeY1idTk4u+095oESEICmtHWrDWWFM4jG/RO55PYNVl1grJgNMdxp43P
5wC+Py/ZyTycm4ac/o234tyeDXNy9Vw5ma+BwImokaIG1evXnuMcUsf48Zrr+3hV
0B7LxmV0QlLYq/acB4Vo57BytUr/VKfBfJuXlZ1VR/7EO2ywwvhMdtkg8/KBV0qo
bzn+a/3oQSLHAFQbieI113BvG+Jhc00sJoQiiT/8AIJbwH44MxFdy/0Zn6r/rQQD
SD5sHp0ei3rLFCwaN1LdBsbzVpaAWgiOg9gkEtIpebATQ5BdySz4ka9rR7NtclL6
cwMoqqOmX6s/4cZ3veXZppNbFg7PNAyJsf2ZO8uVF/8lrqwgtOiW/xOsw7yZSVHn
1ESLL0YsIurCunYOEBgdAFO76GpyCzuTkjSyNO+pZRplwzaqY2rqxV4wGo2DKeFD
ldhBPFEiX+LPX65TyJtHYqxHP2QTnRpU3gagDfMkP4WOZkdzOtC4HCbb/h9AntPh
S9ggXu/8mKQZ2j00mVuewA5tS0qHXDCC+vb7nNTbROGAynXppJDrGBMkYO+Z8oFB
rm8yCpLtPZyJYrMSzwH9Gcc6WRm8uLEsqhuuvkbtP923PqEwKTvzTIBCdoA0yTFy
uMXLCx8EiO/E3/GjqD+NzLokpyD4iUDChx1m8Lzoy2InxA2Em9xDF4UxOLIZUYb9
sBABKfFg67cuzg17LxjuvteKkdZxQK3zmOb1IttgPxLsoTTcCHuPOFcQ8a6sDcf0
JvrulD1ucGWoWrsXK8tk4YOTfGraSIvwp+oCqSij+23nJ3YD9atLP3BpX8gNKJup
TfpkHKgIUQGm6ygZjWLBdfjFtUyPGC4F1kylxZsNZxGu2SdjjRtAFxk6rFBbdJw2
Kl+l00TGhjtA5Jas1LpgCV8YQSC/Y1EgdcTpr+BL2c9N938EAXZ++o1WDaJTnAVW
V65fZJ54MNNFgNZ+x+CnPSO/MH8ku/He9mOiLjdtT1N/n2x04d5Cc7YJSNGSPvjh
95uwQSr5Al0/lUUpNqf6X+SqH2774Kfjd5KN6PMI+PAO2Sbw4RWq8SrNKJbzv34t
1JebKxNc4UDzNxmIub30wrCskX2OY+CPzzgQcs/kTe1Uhy3rfv0x0b4XjnRwEooL
rGacieGpyHy3wzK9lHbLbcX8gSDgAw1oubo5g+WiRnDWqt46g5i1ugieeoJ2SMt/
/pD8cM5C4ckvZYh7a1qF20roKsrwzyp2GxqwgGXhztOxGT7II7fY9Fu3vAMFfrhm
6x1y8fe32A7J2gczi2ml9uV6EON9NQQCh+ouGeHdKNiglSZul9nPEhCowXy+bhlD
mDRGorCTm/f452Qyx13yzKeI6CVVWlKzPOvBy6gvWn9reNN1mzBAjMS7NCc1qzf5
K8g6h2SISWnAPnMzTNKC58RdDkLQGZDyyxc0d4EslpSddnFEvg/qSWFNyc2Huxfo
bRKTv9Zf5DYLj2Bqwh8wW9cP3C7QzP0KimpB1KrHCzyQNtocSAvOfflm8dWeFNqn
xB+Gs3Wl+P18SmtTGDZ6lupy+dZ512nZU64+5JUKyEbXxdBU9R1XCeDHlxG2Ehdv
pqQQ6/WTiREick/E47VV3rTyM7WAzhfVU7v8JQROv+EvLtO7dNl/HpTJ+3SRW2lu
QnsJ6cEspTcQ42Odz+dz03UQ+YaQm+Sw+j6xC9iSpZqgOJaix8rZtY92MlALHWCH
SWT3vIedUwUjZ5r3rnzI27E/4yp5iEYHBQ8P8tkQNfHoGeyveOjDHbbFGo1pA5o/
o/N8WV1HLgsJP6ffjQV1uG6aGbGk9u+hWhfOQjvBTCnGx+gRsS76quPlyX38+lvE
mrmC8PcJuWKwPzI296bXc7dScbp69eo2HRKCW5ZBVpEPz90nXYUuR72urAcTqq5B
pQFYIdhV8DGjTYAZd460ne0fDQOwtEVFNxtP/Dz9xQXo6+4tZeoNdR5t4loCwtRa
sYYHezK/uIolR8pPhinoLU7gGAqFoOk8KUW3hRrNy0uFqNqADKI51Z7JU2xq5XAC
CTpaRDNrfLPNgjzr8u+luUjUhYgWpxb9GX5oluC49v6NGtjWERPKCG+vl76rhHkO
qaySaluo7Gfk8cQgcyalMrEIvVgT3ux+TIGvH8FInvrwiMLOHXg9EUprBiySLGJS
iv9pOkwVU9vnRTmR+BD+/ael/0GGBm4ZCcURfIZ/irkbkIw0RzmavmeFMPi4UCov
0v5C27edj4Bo7+a5BvcUNYo6g+GmlQOLrFqwhnXk4vS4Vt9cbX1x/nesi2TJqIWa
v+A5J+SHq0+Q2Gom61TNwJAzqtuWDDJ8UFD9eYnl5ktvgm/35SwubIB/AUITwEsC
ucMzsCsny8mMuVNtBpmmkTX9YNcmf9oqeT66ySM1t7WgnolzyczCJbFTXvzxtfbJ
121ev5zPikExSEUokSbwzsA02CLgiEQcpx2/Dwv8D1HKPQW4vgREhk0hBYp3JKq1
4GpjGQucTM5B4AKIXgwfF65/Q70+DzeZmUa3wTCWI3JHWmnAqXDgUw/UgVMZRKpB
Q88OIWZxmpALHIOORQhyyoVZWNqLl2bWEJl+jUzn80ejP6N2ImHA5cY5jAZYY4/M
okAb73VifRo9BQE8UmmjCbd2TSEvJcn7hCc/7yrT46+D5p31omsg5xlbnRQbdXR8
5c+xyZicBUL80IxzMO8TecnY0HoCGm64nu/tWIy/dbDo5fKrYV+lNMrBdQZiZ7rR
SOAZf7iQwF3aPvnV4S9YFpg+XmzVKuwfs1QHv2MUHS778LBn9oHGg8Suc4YoEc7u
k9+w31THKFiAA4PXSqOruPNwcQa+sYWtknBJKoZbmn7s2GDXfoMI2WsDBq3oAmSz
VOfVoTA8idcmSp/h22ea9WPJMn0IoXDu9y+7/AmkjHJ2Iyw1nlhexZTdCZCc9ygJ
kOGLRfPT0mRpkP1M8Cf2TDwSVCV8az8M4HQHdRzp3lW3VCpfkzRlgmB80t8883Gk
ZRjBWauXefVgC2yxGlDPNELVZng0vr/FJ+a7XHXAdSPit8h+LlzNwCItjEYvz/Rh
Nm50czTgmqgC3e4LW27XqEtdAcfaAIcIfE1f1e6EPN+KZHdMsHGMgyVHv9tjaUDB
Jt10lb3ccsjeVo8hobGivP+LKGHEE0i9/yLKiGByuM6FDAbF0x4P9FNOqBsyp3dN
DyDTYblXsSI8VK8yuQoCA3jJCfT/a+iKRO6366DFOJr9NC2WHaGsxfAD2KhuGpwW
3L7tE21uxxcYLVqXWBDB7+zUzOmYNuyzYUBJ4AiGJ6z2JRUlURyvLnV+hbxQc2zd
9e8TK2HqmFMmo9U/2MdIdz+TGYD0nNN2La0ml6PQlXGNB9+50Rb2S21DaMcFmxF3
vaiRDpGSUgiBAFfjBlErI3520p1Oxis5T6potzKECwIAvgBJC194GMlbRMNNXFLn
0N8H60DvzEAMLlNsGyI6WUpU2+7tZg55aVrsWBh80xxawf6PH45CpAyLjv4jpGzz
GS/geueJmZuA32CA7fU6E1xVH+8z9oY5WdfL4amBUhS8WrpMmYKYmcKnnruSgFM1
CITcSrNOJqPWdzrgtW+aMoDNQnazdQU0WRGEBrWrbFgMIc6Uau0XgKk+g7ekR59Q
u22v6aXrsoBKG2B81hwqkQ==
`protect END_PROTECTED
