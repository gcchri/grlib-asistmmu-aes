`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1U3d2rQEd2CWflmAVdsOhCd+z+KN9QB5hFv+YLejj5xgNaZ821TvgC2Zrxa+Frsr
KLLnlznmWpCMbLznOvOOZDzmXTTkz6dL4UiIz1bPpNL1ZsoH5w92UpXUubko2iiA
jd4Ro1jJPED6LAgUCNiyywyiS1R654bPnh3FSZg6Y2sGqIXMH6p/orwwVXGuFp4n
fKtfmpOsBNxPE+V+Xdnm5XKl3rUGrlh7kEJkMJ+8D/JNLjmBRnNO/qvg5HKUjmI2
xTESC/aso8rDIQyd+rJGtkVdcZfMy/ErQ8sag9vWuEoUUVmAC4cCqv+Zwwhxuyij
caxx8/YJpDZL67EHxKYz+IfFiwYGyuZltGEj+8K0bcDGs1uBpvPRg1EJ3MbHHgjY
K/ousHxh4dE5UaKq/+f2IzPqgCGC1SCmg6hzLSz5W3acTF18X8s0ht5z7tK+fbg8
aYhMMwb4w1QgYZbPqLGlI9xWc/gEHtF8XSn6jZrEqvcKx12CY6W4p9Q1baxoKxPZ
VBPeqDx0zefuChm5T0WFxN72vNf3UVcyNabDZ8VTeGnFGRO/L1mTEmn6fPxf3cmj
BInnY9KCEvOC2jWUkP8qNNCV6js5zVI5iUqepQ/NUw/o7o8A/3+E4O3V3N5AOeFq
Fj66hRu0CrqJdbOHV8X8cH0avoTWz1ECBTrDM6C27WWKdPfNca23gFTN7j7CEDZ5
ZBRdvYOc7xKJ6rHq+SvO60t+JmLibGHTKXfJyitqpIJWJrpP7dNEXhnKBGhicgC7
fxwqIGfrngeDo9YiHA0squ8AZAArICxaNiPxFs2/v2RaggK+8g8tbCfli+ePv4WD
4xOcaIFHT1u2aHtOI3Vv/gqzS7I1AIAlpsj4JDLX5IeNljf3tSMTuve58SW7VAN7
21wuJhe6kZskTrcp+AZy+A==
`protect END_PROTECTED
