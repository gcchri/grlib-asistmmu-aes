`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NE9H7Jh+59Kwd/XwG+V0gATeBrt6iQrbGHrId0RzDcZ8aYxHNcxymIoA6xUyXAo8
xzWmdEmLN2xT/tYLnKNSeh7hznt5F9OcRg7Agv58k6JTQn9m+MuF8ZNzddfF4pFj
qpbwuocL0oT8jgZb7zsNUvVgO6N/UaKCWl2BuHgzke6a8VBAggCMbkOynOMTTJrx
8xfl02mBnE6tQRGgtosEn+s6U5ZVoObhD+DmtTD9ZgSoQBEET5wtF3W9AhWDIFfk
5e2hN/pZYrdHxrKH3hMHUodl8QuQkdntniRWNrTCYbRl8Ylz/BQwCjA6CoS5gg14
MMHf6k2N/Uo23XIL+qSE1c8WkRk8t43rrgYo6TUmiL/dxTJPm6bLC5uV3b70C0yk
p/aCidwp3IFLc2ED2JJxZO1qpWzvE1TsntAfvBytB7/IgbZp7NqbHScJG1mvSDK/
4Lb41gzSGz1ARaAtYdhzXnj0auUVasV8ryJNSAQtpsn/Pq1/wvD4ZcKLOIjoFx+d
qF51j2+kxH65FkK47v0x1mw0ZkP66zCoH08XbsVZq/WkN/GPlqhoZszIGlasvoc9
i9GiikRpvNV+qvtsV4G9Hg==
`protect END_PROTECTED
