`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lhpx1rUmi1AYbygKDer1EM0jfOlMHJMrhNGAHr31FCkSkxWSvC0w67Ycb4DSY2/G
dU6HYObgYiwEp4ikZEoDNGIbKzigWtEo3vpvZcwzNPFsXCt6Igu4M8xDdP3w1kr+
jf9ycIm9ZwAu8LSzSPbmwYV9oeSDKu1w+FbUygkhnbDibEKOX4pFkd0pARasA5sA
ZbAxJ4eknNiiLytwG2XuOVSb97ZmG1CpGUiCzX+zjgCv+O9cAg3fEfI1uHVrtTBj
VhURlgdq+sgXEYmGU4qKNShbpMv7tIg6oV2eZ0vdSc1TxjGfVvu4eiii6FlnyJvu
HxO7vW6PHP6M0U53uf0dFY+tjZzO9/PTlpSBmvyzEHTwWWxhEpSrs2nZyRTUAtY4
E1TjtlqQdDKvsklksVZw8lgM8eIALjyrVS4YOmDfhOE=
`protect END_PROTECTED
