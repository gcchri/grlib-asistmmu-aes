`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ubUMS4vMISme6hlbj7K8UpYjkUXbyEzlirsa+GcCn3CJ2qxr4XfS3qAgbkX6hMrz
F8r2ORj5Zwhx5cU7EmKsljYE/gy9Bx9m4SLL5dzatA4JIyv2JY7SO4+ThrwGU3zF
i+HtV0ztHhF8F/jZUU78R6z+AW0+evGR17CJPOFAhoNgTm2XUONTQDeYr7/oZx5q
Umz714oDrjOUxHO+RDRxh0pqRA26e5WpXL9nr6CU5xJnveKGc9u6tIdVpE/RyWXL
Z2eSIGsJ0uFgnPCBQCFWvQ6CRNkd7WxSM0Lxt1W8I7SSPrhmtC2qlDvjYEqCO7dJ
T8mzGLSVHT0VqnrXzZyHbXKMX4ziWgfPuDDj6FCItbfmmzHBCZaL63saVddy4qRh
n9gZ9oDtoyE9SIe7nrU8hQ==
`protect END_PROTECTED
