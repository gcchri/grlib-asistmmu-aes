`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vtt4UgCvY5srFHGyQAW1oR1CPOdP+R03da9tbbNcFbQx9rLneGhwpUFIqMvW43A9
P82zgRH+Hh/m95a4dqJjKOTVX4p+IELnnEMxqlmaK6xBBSDwyzEcEbNK9CVkR7+I
0X7/fWGX8z6iubVSrwlN3A4/JsTyD9cn5MAT5Qipp/qk1EOxmFKp+ZJAhigvC6a0
Fs+Vni7UzJbGY6LDuDO55qeybmtm5qGbCGXtNUEIudISWNnj1C+faKxGJtMx/HJ8
wIdHiw55QeAcOiv2Jg50IcZMZFBJ3aJfcJpmzfEj7pJHOKSmva/5qmL4l7unVEh7
JB7L1xrogbnSGOtg77O1ZCSRu0ov3e9/TdWwZUVpOpMIjIrORPZSlhwqJweTTlHQ
`protect END_PROTECTED
