`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tbt3HPh9HecyCXzCn3yvk0nZfV3HLPGRZRWeaBKG+ADfMFO6AUUDfxGYRImPjBoq
G+45bkWN5UgSJo6KP1Ft28SJ+kFrlo2KNcOZSkReBGiHNGDliz2LJfL+eD8PZVus
u3JXpak3/EzGdWTlGg0cEmmIPvbWtelUrjV8xMcT5ZKSYvl5/w4LpSLBNkdoHtJD
QINV6Q45X6J8lgsIi0xXPmy41YXJtxfdy5BBESVUK2dZjOERFLKOJLN13Ipbb016
faa1FwLFQ7PFDVsTvJ1unYa9Xdpn8RofL2ynw4bQ36Wmwr1hdz1H/T58cOhmyICj
dxMyTlsLVs0FAowDnQHVHKv5D4JrqIxB/+XctsskjGLOoGDIZskjzIpMmVxcytkW
RwnWX0/1MhwroTe/S+dgyEW4z7sZ/v2aTM6Ib1K5oN6d+nDMqGdNLolktrPDnyB+
uwHZr9TTt6YG2NceK1kVvP5yE3c4N0xtmWWQjNWK+Ou1XNXrVwFyXKVRHcD1zfrF
VN6Tj3zC9EHufRwCBGL3T+LebIBQ44dJGkvqt7WmskuwVeU9kqxBmDg0XV1owW6+
QoIiW1pdrgMqiRMYn407pQMJtBY0VzjoxTCi3sYU/KwJ2d2ayg0QVb2hijmC8FNs
d7jzAHCpOrrK4f1/kSyDFG12XXnN9Nj874fLterlCIg=
`protect END_PROTECTED
