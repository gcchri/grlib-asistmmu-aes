`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hioZEAeHvmrjwV564+g0jZES7NLo1iTp8mSPU5AVft+gavPgAC4TxdLP6pI0NfPN
VQKW2ZX1DLzSmk/WIWiTqcybBs+d2xrvIuTmqJmOBILWdHh7/uBakIiXKlR3xFGe
sxG5tWGk9HgcjnHb40Mz4jgTXhz0VZtNBR+RX1N4qrWiVEEmuOgGCaQL+pGy4H9I
Imtib1HsAOxlEtYpbRUJeyZ5QyXPmH9TxH3bM2p7O+sOLaX8sd6gTBjtxv6NNh+1
gNdCaZpBYi28wuqB+/k/vBaedbW0asAoB7qfQ/9KAlnhX8iz1NymKSyH0rlhxKe4
7otqcKesced+zOazsp79IKQt5sFXF10jSDenHJmh6JuaoL0ZBHPlggihswHe0ihI
dz327gYJDBumrCK/SsoymOqjF9PrwmqW/Lomz+JT73A0viFR2v22Hfay1yukIB2H
pUqclBzETSy6BzeUwj979NAx0m6pZep+GSVQcX8DfD56vBEX0c+ZNP5+R7C0r2TD
JtuxcIu6YpPJs6ZKLap6o8l5Ngu9aJbNlnPxLNNYjdRw08wVlUfljFAqWalr4FCV
YKWpjbMogckaCSadWHovhckLlBFWhDxAUtVKLB7e+nFtS/+T7xTomJ1zR8WPCqNd
Rjz4fY2Hf38rQGsMN8TMAjGgUuMRrj+23H5KcYLOGsH19OXqyReJkSykfkYdkTqU
0JkwZWs7xazTfizu1T7k9Mghf8CtX54s+c1ycuG41TGHrc1Q1JgTpBgZzzJCznlA
U997HEYga1XdUQLyxD4I+A==
`protect END_PROTECTED
