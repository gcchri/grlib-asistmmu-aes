`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bOcUAKfQ54f/wUykzopJEDIH63fitvhzDwmlksK2yL9MS6SFM9Xca/uxMII+ZgSZ
c1fD77P4tuy1vDNbTdb3G9idiWEXmE7gHGUmg3yk8xvGtz7+4Bs6ASkghlL/q2FP
MbYyjxAYNpt4Bv9HZs9ecmORLHy/S83uuGEzaW1+UznC3B4qR+e79kuxXwHdLafZ
eGj/p+/ymavd6x1N/e7c6xIecDnciLP8+G3MwV1zvtOGD7uni/GYdc1DlCzDgcDC
BBd8nWiyUAoCDmKSFMM+QYz2ev81Q1EKcoBI21XlDtpKMqUdo0BN5tYpFq2RIHzA
QX+2Qt6yPeKUGSE5/Ut2aT6LWzLxfhnXSNEbotyuZs5txjHlqiJd3EUR6JrGPOkp
cnaAp1Effaakm7Xpl6AaXQpDtBdj2H9SJubxZYr9+pHex8BxdFAcYt9bmrbrFB5c
xFsHj+D6ZUhlMZxSu2EoNrEHXmnUWV9WdfvYl8yJWYBHcUuGF7Ii7ddLcgDbG859
OOagcyrdAS0B5d2ztu06Ziiykkhy9yzeZhf1AdbTFgo0b7ATpu4J5iyJ6PmMZnpx
`protect END_PROTECTED
