`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oPZRtqGw2oXMAiDCgoFYWh6BpBfFn3/dfmMKKaQDMwW9DM5EsnxUZP/P+uDoOg5+
AiT0eQNNWmioQIpl0hAYdrL2IGrdG0d9dVZsfbXdvXJ+ipZVdnoMuca+0wzNSkqM
FPmVAfeY1bjZFxmIjOjTR41TIgk6nXwtzw7OkOqdJujU1SHuKKoGu7WPH7MLGpbY
pij9NRGtDoOJRhKIWVcXFEJLKB8ceiUZ4081PdLHqlOJVdIalzLgKke1QwGK3pm2
n6LdzM2df3VeR68hdOKg3tYND3GDXNCZ4eyerP+ECUFaiq5TJz2NAc1EB2YdkiYW
3eDjJ+vzOPRHK44SOxxq8Kbq8azEiUa/BbSjgYzaqulb8hCJU12lJXJjLTPfJ5EA
rj4LecgM6gS9mc5vACvZlBYkKUMI1ii4ACjnh2cVouc2AIWcrN2pdLWRmwf/yv4m
JqkT2Qy+oYFLvjbaBq678Hv722r/qFr+Oc9TGdaFgCapw6crlBpdESiS+um+U9qK
f0DG13YiLgheTCmHOT3pUQG+YbxqSQsZB/JxokykHQkgPmucL71jrK51k2tJDRmu
hLUIy3YEpDD/nVSBi4XJSWgDG7Mz4wspwYxNxrMYVai7PRQBC0S5yy6uGDJ8/Dja
lwoDKx6QL3njUNx13EHwt6DAmi6M5qjOsGJ+9rMo1dNodZOJHUkSHmDl0QmWEdfy
m/l9IlpahMnwFUfpbIj8Z2yHCL4b+2ti5ljmWXK2kwW8ZF48Ky/6uUaLLbwqa51q
fB+LHPEVS/RfJrvv36POOgx7GrRD1pm5l+EshkiD0G8SnBjCyfBkrR1ZrUpkyvBs
LY8rXDdxIfhI6OqCfX6dIK2J0Tj2NQ+qV7MTFvakK79wbFrxfXcy1wbpNRRivCnF
2punqPECp5vO1J22dK8zE4sPJARS7ld16AdrRt89IAC7cYRNiRJ96/eeXFK1Lq8C
`protect END_PROTECTED
