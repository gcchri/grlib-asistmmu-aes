`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jip6bKLvno2Q76Ssz0QSpetncBDtD1q9/QYjLjblZ5Zc13tbeloSbJu/50IaaUdn
4X49YyNACWYKpf/N989BrdbVUGfmuiJwA0zpeMyb04PScFCaDMJ+GwgIpV29xuxG
MuP03qvOfI6YCe6ojY7iLDExtC/43KOMzrIE2OM6fA8zwROfLoz7dbZ4eHXjFbNK
10Jg4qmkmC6B0er21a8SgtMu0QxeEdbX7r9GgFF7xKL/YMP269bnFpeVYkqUT6hZ
Mk4ymIIvaYD3yr0ePj9VGnn9rFWtvGCXOtGNf/8jbJ+Nzt9mqcRQchYDlrTk8soy
n3Aibk4wN4TLuG0sVvWskiR3gTipm2EAZ3ATQHsviMpbAA7mDuGl3COqzmwOJDE2
y6jj1znsrjTcdmW64dozwnPE0+dl1Q+Uct4t0eNY5a3ZM2bDNqwlsxaObF4lfHtB
jUflJOEfr59yL/Sq/APl7HU3Xp8tKb2n49wY79iaRQEJR8thlJNeSFMJMY41zAdd
lFKkoGIVkQrJEztBFE+VaaitCBW0KNGbLrhkFuV83X8Q8pCy7hf4yrpFH/lJ4wRd
p5zRPi0v7cyu23dpgAFoGPX1EqaxDzzrybkbvJdmCGe9dK4lotDhpLIAPvUuVuu9
bcerdQOm11PISwy79n7evJ/4AJNOpDS9OOX5BxrYAx5Po4qOUVBa58wCSy3Y1EcK
NN7eudNGqAdGJpdT81zKKYJL2ZU8JtSDBfNw3VbqkdyHm2JsnK+MoqK6hCRfnSy7
HMd3Xdk60JQMULnObHH+bcGPN2EMx5rmMpl3ur0wmheH4Ru59bXygZhZki7BuQ31
LkpHy3F0Opw4V3Wq3tTQ9LsyvYgBatlbN4N/atowUixQlRZ82qidiuwjsrT1MD/3
C6+gFyNjOPeRWH3CsMKtxc/4tmOTLZzWLOi3F6oVY2v7HkEuh5dFEWq5DHJHE21I
HgumZhlONw/2HyT+J0ieHslfxi9CwcPLiGbkXuWV7M39hxwPqSLfKzCATojSBxqr
TNZFnDBHr1P5g3P1Qply8jFfuzLr82amR6XnDpU842wJQxzdgRnDQA0w39BPYZQu
V0NcpaNY+H9hK+eg7kMMusXNW5cSXJhSIjuPHwuElYemjX8bduMq7c/2DKcJAzlT
Oy6UcnK1mLbSs5gqkegJzJaPcklO0GrS+LF7Ro27cr9AIXh8te8kczGLEhEiZbpH
zOOvGGQDo8HiYm6QmAhavEoROL1jWCloCzji+PhT8oQTWzEpbNgg90GG/9KVrwwC
Dg0PNRtpmX5V//NmzaFXa3EeGYgRhfJCEGEXhmz1YCArHpjchjsJR1dP416vp6RC
kZXVCIfOV9v1yRWTiCuxNsMwKmGgTGHC4BvtKGB1+4cQfCCobk98nEGc8Peb55sX
RatsjnZ/iR1fdVDiXYWWgak6Oa1W/lrfMC3kIxLtE6nUpktvLXjHtBv6pAyDm4SR
D9jtdo86jbYM1AlmgRAqemrhcVjZ0iPmiyhfngPmgN77TULqefSfiwKhQRMorPhd
rMfjlPKpu+CKD3kHNwV6UIFl6+Yj9jmwhV3Bd0TaI5OeWigAdbxwF2t+WlqlAKid
1ydNOEIhzu0WDvlYp8u0rn7KFcdg0plmu5GZz95x7yoCIG2rLLW1YPL4/pvy5DTn
G+96PyqXoQk7CAxfeoowlFdisomD9T3HkdoAzkc56E9LIsy2wyuXJjz9M7WYGC4D
Roz2tUQjCHNMZDBNiOamK6S+ePbdB5Zz4Yboxg6yp0+cXp2LHBDumwtswn5Igz2h
3xiCT0j8fqfyV9JeowCYUdokXG4+9imDGUdVaEeOfv3BuiUAdASOQzi3RsymKyAc
XkTraTXwqDoZAuU/Q3Wyu7rBw7vFfDu3bE3xOTBa6A809buN/exA8eC4H4e2GioD
MJCFo64ehVQ3XyM8mLGEjWatZEAec7vCa6inl/HZk4ss3xkwISHWWHKKMcOyQ/RA
XSgaEsZPXRblND30a3/Wq+xz9ZqHQ5zUSRnEz68O0ltGHw7InZh0MQu+d/wbEfqH
oiNMHbHeoYi76nxA5BSW3m+taTTpaTwTxHs/YDelfZfK1Uoboy8CUWzgpo1O4htX
PHo5Cv9ih5xXRTWCQbzR/6XOO79vz8El+NCuKHrs8er3hSffP9gTvfy2LmuyvlTp
XAc5PR58j+Q7pNgOwNlwhJoxRd1GL6luYLLtCnHMtFybhGK9vEWUeJdNIWw/Xv7i
m7gdEipKGLVIHo5dtUVNKq/T8IQGi9DMWOExIK2Q6pw=
`protect END_PROTECTED
