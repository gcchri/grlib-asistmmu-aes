`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MkngpafOitspBy+lXHJkt8TSBG9rZ4iEJWtEq/j2wACFRS+/NFL+W/Me2ZmAOFSi
IYOAnqy/FpvcOh68FlRgP6luOjTb4dLXcwuEt/Sp4B9GhbaIfZpU9lFJ1SfDbjve
HU1FerCeqvJ12uZPpyJ7hLP1DMtFTB6cVMTHuCIA+hiLODOrtdwAZySOp+Yji4op
v4nYTjZ67NegEWprc6yuzEkFhtoHPYY4VL2hPmDzHVIajVrtc6erLfJncPnZG6Mu
4ocE22+i8Fg7F8HmEdnZdjQYXCxTdPFoDHgMEVjSMY3yItkbCG5uyL3/NGmMUA4T
1b2GqZBNHNQXLv1PHN33lt+d/yOopA53D9Nqd1GzLYeIbBb/XLLGkduslR8LiRac
AXOyOYjIgv6UgrDJCu7zyKIcf6b8lnD2inoY1Fl5Me387U63Fh27qBW12DOrAD0Y
xZEDMu0YAb1LVqe/J4qmmMD7ORE9nmv+LrZw6aFIpfrWWoqQg+986TsnKyco8/Dx
ylCV3OzupCM4FNwiEChThyzs4C6EXMnq8VKcecOdTmetpgLnNCz+HBQDJgF5RWKf
Ef9LWrzplTLZzgrYZMKsXeIfHiCpH6QocizSJtjfqvPIDEgZIfmbZKR/lKAnvplx
Ypn+uztoK6u0gDqoOuyKjJtSzGjgXV42mmwEKFGonQRdo4iB0hIR37i3eD529xXi
g7TlKOeuh1E4HZBepZAvdCewTFD7ea6rooLBRO9MQtTheLXnbjB222ChpSjCYAIl
IlQD5GXmTsQ4UNhdUOcJlt7R78ytxT5E3tjt9Y69DvoeFdgscIvTed2eTYG6Kf12
zl1XFT5ag07aFlidzE4rievydJF3k3NIg1qGFzkwIwQal5HWA42nNl05cVFRo5KD
ZvVj8nQn3u+JwkfhtR4a0On3+ckS1K8+YNV2JI7aio2SvBLHEzIf4DnTaJnT2T0m
wAjdrKjse+IUUJwcQGoEb6Lzdr0fExIBdTc+p6vvF5tlfe9v6dZGNMCxOm2GZ9Hg
TnZS2H2Kzmrpv35gBn5nZOxoU1XMCuLFglKttHI62nmnyOD+NAdGe4ydAJcfnWAn
O4K5MihRmzYsOvsUFNO2Ii9TysG6HsPLyCbune3OotJvT9DQXyvMJK03SnXutp/m
ki51j3xCxPNlOwi7DKw2v6z/JimU0R2BQBq1PyqOulhHEITV+MBjOk3KR4C9CvPN
8pUZRjzu55sHm70I8vFPwQ==
`protect END_PROTECTED
