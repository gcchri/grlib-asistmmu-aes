`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ixn5DrPfMPonoaXlBonqtfkOVZJzdBvhI3wenRGum5xBNvGY2ItO52CY9kbTaF+C
1yWpHJ/tHSS5CVMiEg8nABPpLlrPy2hlfLuliS5w8GcY7YLmnDAjUJa1I6C5jeIC
/vJLpBx6FsrUasbAJtG0TP2LTvGHGP3nPcP1bECitzepIy78YZnbHPa/tAC+ZXu0
PyjNgdE2cwmV0IWYegL4DEALMBGPqMte4pub93l5WxjvqUW6kwhY6++jr2fiC8Ok
TeRE2kcRLXx8jGtCZ02Sr4megZ2Tc5/OAzNQWxTQFORS9sTb5eA7AAmxqBLx0GAG
XqfDSyUaAQW4cBV88EgZP5aEtvVbiFVcRgkNFfyjxZSTnYQnJZXYTmwqmzwiBCDZ
ydrxDnlt7S7GFHt9Hp8M/h7DazuwkOb4ZxjPRwkZxrVCcZbROlvLMQv+JJnZVUEJ
gjDi2kGafaUxprYyWqxyUi9ldxXACmqut6Ci+siYqpVh0YE5KcuUpqSFhL8Muuji
Jv0E9/7t8y+2fl/tGBnDRylfazbvrt/IczFK878L8AbMCaKIDqbbshuJWCuCJ9OX
s88IH2FEOpepcCnbghjkPpD5lBU+2U4pRzzB/Qa4UgOpWiFnTrkQR6ivD9jxxccd
CjpyZtzsC9Jr1hnSQXyduHHT2ZHx48RbH7HAwEVLHl4TUhIhI6O0REKOAYx0spaf
RW7sxPEm3ODBWYyeyUOerJ/mq8nwRnmk0o+qvEJYEVtHRm36OrCx0v0QjysfxTmx
tILmqZ+SiU04Ej2XJR1bYQTtBZpMG7uVm7h0v0wqB7x8SCcnHKNBHPlXcWuyE4Yl
qOc5iinilGJru6szvHSOWwy7fhNHQFB7/w0Ek1qihHyDn08RZw3gNUv51MXtGdu2
6dUti00O1K3qEOPHBdRCF5rELMWgZncyYxWPeEXEHYTkHk3BJxTrlJQE2QAMLbo7
`protect END_PROTECTED
