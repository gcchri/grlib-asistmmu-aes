`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bWkqn17p+6SEvytktX1H7vVuH3qIlhgthdb2aX0FPdTBrxVUMESyS6PnTtmDQZtg
0CMjuBm2hJqzkjeojaLPz7mOsVNfgsSEx0ZKIlYwKQQ8FTh45cSFLHsf02dKZO2f
8WzDWmCmH6FTCcwVksT5KEC/0rvXwrgEY0JRJogP8tgN4k3uybLV7nd8vphIadYx
QLuPTcrQjYmPf3k+FK2g7AQ7j2pUmOW16xUjNFqs+bxPy20ZL6ds7J7mehxbAxuI
NsSPnhxe4M56wIenO4JNaZC+FSuiXi94Sn453sps0OndCDkMMw4LGCXUblQXmZqo
JegX8P9oOdEubgpYOs5fUewUpaIJjrayI4kijW2Dno9QpcbptoIbYFlMqKeV0oMr
ER3dzEuvjQ1n5nzQivLMAk+RqhlhZR7nfUWtcVx85SA=
`protect END_PROTECTED
