`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oh3MJtu63oizwdJ7V1Qqp6PsPZZHIVXOvhvGfU2NWMNElTF6A5bpe1pet2xH1qsW
QTxXaAREdBzYY/FRMHralUUYIIacNUjQcOdQv8xqfMMfBQbhnN0lXt+uDoYeLFcz
PIPc/X/WvM+shY4MIebxi5wXXslKsVpzq//S8NYRgGL4JN+yWUduDX0B8y8K9zxJ
yCuWig+sXH2LNVW4Iw/HsEixWckc3IC5EUqf5vTyFbk5xreFFiPFjsvaDcfiJhmp
Ye20tFmNDm42zHeMUZR/8bFvCOeMr/XWJCyJ+U4yA2bCJcDgUXr+JLrrXGZScmxs
oywBWn8UeiRWmJmIzEha5uA7mk0HytZv1p2uqGuB93FfE0akDCvcZVwlbee3KRBG
`protect END_PROTECTED
