`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B2m/ovDvH8gTn52HhTbKrIm9KfMHdCzIDaPb3Zzjdbz3yiD1207ErzYWvOxCokDg
Iv3TvH+pRQqhJ/vxIi1pWN+KhnP0OALPlxjO73+otWg+Lj4odcqcXswaNFrSoF6S
94ibjiFFQXC2p3IDZc4u9QZmlWzMPRi6PBQ1Zx9JAr36FhNzRPZXaJZ0WNyEnPte
qQo2M5Cwh8BsGUI/VNFED50XSw9vFYFQdEiUUEgHztqBYsKD6sABT28hDopsnDki
VxYqPMApWxz7t4jB1reySz1wgrtE2GerD0RlgjahqesNArCR6Dstbhq282+7stRM
kExqPGYH5arKqPZcsmNpn1EpSpdaSHvVLyHYJxP1eztQNJ8lN1e0+in4agFUcvXB
aDBuI9x1lmLzTN8cWBtm8A==
`protect END_PROTECTED
