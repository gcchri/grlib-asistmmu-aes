`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uOFy3BXLB6pf0V146GxWuEg/yTsoDfC3gHEOsPp505q8lXJ2fIyAi/MgINAv3nKO
Oaiyhd2DlgUoiB1Iy44Dhvkg4G8oRZWUdZAB/fYRkDfUc2KJ3N3NnIndqoNBOJSN
OlqL9D/6XfLgpruzWs3dux4iaefslX7gZ9h/i8Sh0S2l+4aoqZhaPACQt4UmcHBi
Y7EfZJJlH5hkVAyi8dWzLXfIzGmqR7mwDJDkZ5sr4QjbU/YXCXAm1Wj0CEa909px
LE9j6efrult+z1fQf2NRFgly2qD/mzuxyXB7zL4d3+jXIpIjMDZzI3iqbMP77UeR
Cgy07AaVXZsO8s6RXHB/RSOi+fQACbg2lX0kib7SvC8=
`protect END_PROTECTED
