`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SkgExes+TmiDMSWXAs8Zbtbe2LaofpRoK1Lvbb05R5Ek+/gjdZws9FD9ZR7umbPK
5WUIchmcczZxQ9sAKauXV5fuRzF5gzddmh1YaldYWIr5PBF+Odk0FDMew0oCZ5dw
87omjACQ3Zit6l1umfBlheA0x1n4K9Rn/g2RksNNZh6CNheWeoDCoRS+uspNb7o1
unTxnxw0oZxx8ibG5SbT7HQS+xd2BYR8MxVbvCy0xuP2C5MEEiJS12pg8TqFRi6j
cyC9jUUZ0B70sTOCPtPQ9UhjJN6q4Pf4S1RwxTMk07BsnRYXePN7kwl3IVLuBvjH
VYh4qgwO/j3DzmFPvKgwNgZnEq+aMTels9UUvrB6Skql/8jczVaUANqvsQ0rPS9S
iYe1o3P7uT7unmP8yp2hkO3PyAjpADYUowfB+o2C6crx5N83AB7BKw9UNz3Blx+j
LIwdF7GO19/r2ANmEgue4sqBMhjCJ81bjeOkNtdFu3xbYDZcpx1DZPHH79J9JJmH
sTE8sNVYN2mTJY8YyGzMDTwgFDDQGk2JhEKQWiNaCaPUIzBimsWyqorW0lXC8L5L
FDMYlkicU4ON4nZ/B1dPykpu95EjCzF9AbiHgr+fJDc1OU5zJ0MRwo02/P4Y/Lk2
Trx0W2wAjcsrekH/HLDE+Q==
`protect END_PROTECTED
