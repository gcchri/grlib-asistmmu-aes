`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cGY11ETG9Nky/0KbPHhdtxjp2jCR6tuiuW9gd0fabjrekIyoBD8iS6IjDz9QyoHD
KQgyopv3bRYax7UWqI7MF3VMJRfcRgYP+XSuGZ1nb9mDSQAzScrhOAVreW3oLi+9
M5XX+1QeL7oPXkKABZLabxDqcRsYk9CENEoDSXz8PDH+Ku2MBTttcO1ClUJF3NJQ
fwLFbmTglp6TpBN9xWm+PVYM4r+vzRveI9HImmWnuv/KPgQKbeTUxIt0Rwu4yiB3
aX+pWBNfxTgrKyoIA4qCbtUwuuRKZOPVD6ZrNKVDbSRiAWETc4RlD4gcJFam768z
oe94Y2qobB0haE7T3POrwUxohnkFPQf2danw0f8mwi0fgJ8AvMavMx33008EyU50
3IgJHenNhptjjQf241KfglQ4O4HXgVyUu249nuKVZXtKn9O9ltzfsDrPJE7JnGlQ
u1JYog3+pYgchAZS3VDdc4o4dcfyzG6Zyg7zaqzMP65OKw/helFFVYNw4GfslrW+
`protect END_PROTECTED
