`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oDLbrnYLPUnVhZXf008fqPmGLjMuOkVaFuFtbbhvNGPz1RmRVw/NSaN+P1k1U8l0
9nLTSBUPEWP0KBtJPI8K4e0ksL0VR7QDKUqsu+dvCsyunUaBHAAEKfKHyJKjrg5Q
8O96q4yaUOuJL3g7HixOe7YrbpIgoPoL3z+0r9eg3iC8BI8hISxxQjfW6U4zMPfD
cmXGhXgygviaZILlW/zMZz+m1WgMDfcOeyiqH9wBFCTIy6SxiixpQCwmIObVHmUS
5mR/Sf0vptKhZAVILL01FI+lk5XDdSOlscgBL7gHkVgZ/4bkE9H5Qs+yxnaQEoTT
/8BpE5vEo94KJtZuz61FUmFBPsgOo44SNzat+BwJtqt9yFy8Vojw5jMHa1hHA98O
y+6IJw9NguFzssCYQT0petTpvhAh8j1R/5f3jmGjwPs=
`protect END_PROTECTED
