`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BFzse30piOQ3WtQZ7RVrFr82jAEHMMt4n3z+Vd8HSLN81Vuh+75m7h2Zbpcoq2z1
qm9bsA1iNnbY7qhGyq0O7wVi7jIyFD3kLZygzhVEtYtRfyo8j8UCt960joi1MI78
f9r/RZwKgu+Ue1Ru6OpDCv8ykrmGJEGIIySro5eukHwZ2ZO3jB385o41lFvoGnKS
9dJ7f4NYEjCwGVW7Y/0Cqxuqpc5tCF0Y6x6UO5MO/EUEpjqwwc6RDlYTN+4LDFqm
`protect END_PROTECTED
