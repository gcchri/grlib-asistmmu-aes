`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xHU1Xaf5QSDvLI7OHqv4GEqlj6ZOI2D59kZMVMsdMEUrqMdWxqykh9XIq0XZMsYK
WOR77enP2OkiU3SG3ZGXOCmZWDUsGO01+V6xLYLO1isaunk+VGj7w38A+Wqo2p6e
nxWFAeokqceO5+ksoZNAS1nB76Y3Am0vYjLuV7mZXTiNT8nC+7L1pTRIb9xmlZ3x
lKSTpsdwmVcKe0w2lozGLswqhaSCfIwxadQjxwQ8l1ET5DixigkKyz9Xt3lJzu5c
sY+hNcgtH17d72TgwHWXAogUSiiHyIqbvTgqY6MY7uBzjcP6RsV2AAcNafFnG9tN
OSLsAmntcfwCqgCp6q134AEMaRR6NJ04cadAi87eDU+IX4E470MyQEAI0kuZB7xQ
ni//YFo2FQitnTC/5CobOyYZpCfU9Lj3+mQ2qIfq1zhTB9cWEnvi0jkT8mV0bgVI
`protect END_PROTECTED
