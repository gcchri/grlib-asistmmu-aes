`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WiaRJOor2FV4CbQLxYtg4iw5UsQ5MYtWkAvTQh15bnon13+v5uvPu0Pbl4JunJ0Q
XfzMWbxmL7hHfgOLDiK0hFjyfndo5vJF6XgA4FFVmjCyBDYrTGH+bjNhybQoa6RD
W/NyC3wa6N1zwKJTebFd868CI5MoiEA4cZxbdCtfCiMofTb76U0yliDmIR0U66Z3
+a/vkW3gBpNOVpLKO0JEJzz1B/LZ3KEWmyBg7YNTuX73GWrd5JnRXVegN3DeElJN
pFFzK4Lf2Sd4F5iGupb0CspKLjmsgGRMzgPyEj0UpnXNZXhp96DPfsP4ykbtXoG0
be1VUUWSf/a1mwBWao43j+QdNM9mJGWVbB7oTp/CrC/q50H5/uOoGb9r5g+p/fcN
1ACTMRJlMuj+sKFDBfr8hOXN2/yGMwtPikTuIpi7F3npmd/HABgDVBMZOkq1bmyd
NjO5W0t8cx3G0kJTYhUTPVsfpmpEBRcYjEKevM3DRIxmB8LbII0it26GbO6rzW1Q
obA0K5uliivJq81M/lc+CRj6eeG2pI0TgMiQxLoDWAfowauzGCLHAXCsBaKoBslz
a5qZugOw/dCwroZNfddP2Hakg8HWtP8fPr/8mJX/TUw=
`protect END_PROTECTED
