`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6M2LPr2rDh9dahckvQ+AJri/IeXySAHhEPXoeohHoHr+YL1wYuYg5NIc2wWunIBS
4UT1p1TnmDuD0OcEbsbhnO6UkiH76w3Lzwgmg1gwzOT5L4BRAQd1HeUVXl8vS+w5
uUrVUQ71WZ9Ym5z9Lxp2L9F2PPj/TSVS1YC02o5lUQ3vh8umXazqE0lj9b/+1l7I
ep9/Cxd0raD367BEg2sz8yyc79E6AfdP5umM/jSMZWcd57zhuGMfuKIoQyk0G2OX
pGc2Ec4+PTnHdfUAoLOvzu+K7NQkopLAb+cAJW2e9rvhyfmbAoc60zKEjq0+BT/L
DJwL42jZ9wnpSyF1a3wnJ1rNJLGWLUPVt+Fwcm62R9BuFo6ioJIQDVziPv16rgrY
GMhVlguqGSziYpQQvusrYHYHFLGgm+a6vIB089DCkIQqAi5L0wqCof8auw5497QG
dwf0mM6oTF27bQX3LZqtaEYg63jQ9/iAA1EKKt4MnAySuNPYHBdkysbHsMFu+p7V
`protect END_PROTECTED
