`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hFM6IQH4pkySOTz8dO0PPaICMSnxzzaxWmUjFphbu8ifLmmxu7qcYu+u5BMV5kgR
LPcYy+ZI84uHcA1X74ztxsldepR6u2opFLINk1+7obn9dG/S14oRceDYeb39fVct
z/rsaaw8DnkUu4aeRrB+A7bbvgLujdvZcwV3+HIsxVuEZZkBX69lGRzQ5moGFK6m
IgxR45McfDUM7NPBd+ksgNXW4aBuHEIA0RKxqreGDzli5cJ1Ntguj1tISmGp/7FC
9hhpCDcs1ZFWq56jp4u9E6W1ycjbGadmEN3kUboOLblBqWTeU62TSwE58XCWnbNg
W5ZK0rcCge3G2PCCvLxp090mSfWBYvN0mql9mQsHwzuQcECPOgU2NXW/GYP6b17x
0c3r5mr2sXDqVKkQbWAfmf3chkn7vCbIVxmCLKdArE2kXh2ymHTBOd6S2DoWbtkn
FosTKcIilg0chMYteaUTQZ0TGP1T1U2ELeP7hoXQtz1jOaMxzZM5XTjPrlDg6dJO
wNim/gbe0ebczULBakC++3JmmqWCggdE5Dm7c59O1t6aVgq8nDfOH6VxRvM5qMFr
Eh3uWTPmZdXGmc+DPP5mibzQld8MyGoxgI7pBH+aI0usLOjCFfowZ21M7aPegZfU
cjOzBW8jLOEJdbo1kDkLr+otQEbxlCJbTl84uRc6ewY8UOr+ISZ+xg9gs2ziJpuy
T392agO22nsDJlhxuy4AIgxfk+iqw75Kq17SmFwVVYiXy54Db3nkPK2sSS/QygC7
5aMUphdUUOYwdhEfodtwmRBAK9AFl1G9oa5iEnHBJrgZ3E7/UnFpM0cXhAQ4zXkZ
Wyk35jgnG2iSwHoBOl0ijV+vhE9/0fGxLxNsbmvgN5ui7+/caC3ausOB+7qXEiYd
KE+j6YgUz0P/3n1AT58IRKSES0I9cWqgxs2eY1NwWT1sgqJe2i1D9JjWrAO2JRqs
n3HkdyOpMhYVaUM80u31wqRTF6A6sjhXCGdLbmCKDJCJ2LnCmiba+SlU+wicxrUx
t//x66ChtWv+r3g9gvDU37P7j40jAbCHmWhXsoGIq2v/IiRRbyG2z10Vh9U8HE6R
u5NbHSQCDteiWinl11FTGWS9TW1I03DQtjeq9CPZMnxSS97z2TUwXRNb4JMhwrE4
mINMEjQcUzcdUuPhuddpSbUOIblbWSXXIjICT/HSzGhcsWCrTT5DpTKsVH0SH5cL
2wYFo+6XOj05gW8BEewt4mzpoufX/xv7KhfiKrl4Ec8yLnSZyxem4Sln6o4FBhMj
9XctUO40LaajwGb9jPC489DgeXA0c0gIUqzoZpd+r5ZS3It9IFYgqrd1fOW1AuDd
6B+kcYggqb1CU/dHESwX2khWute2wd20+SQXqhwqhJQTRIPh+Y/dKxuXhncWMv0i
LBO7wNLRYCZgofJ8vjS/jcLrOLiCB7+N+pZoHBcPDDKMmZ2xijcmeQzwT1f/5WKh
ry2oRWBOQUMMuVwvwiZdFr3bZhvOM43AQuCFp3D1AGe5XbxvUxt7fye5H3F6HZX8
9yaOM+GEPq/sBXJFnz2sy4pDpjJWINSzKYtHXf+YIpRK0rnXncsqIMMiwRrcqp59
/M6e4JN5/C0+MIAavty8frkvSRx0frS1/NZ737tzSK3JW+efYYgWrwTpAnfSdEWU
8JbJYSxl0Id1V3IVVvoEBMS1ovHckL3FXqKOHRHJHE7+o2lKKTOKx/qgyRvbcEIK
zGNR93L51TMuPDeLs7YGtAXep8iV5Rha24G72feFVOY3IFWRNH8i7C25Lzi/jl4f
LaZqoanNuB4viPcz0HeNXAd6t40mtD5UjRvmqwM4oyd6YxO75Le0sxNzoS6By65V
XgrXOjQelO68JYMADYfGi26OmP/vgSyztA6TFfs/WrJlV1CQAUNG/+m7i4gIHN6h
SJcetT6KStQ7AJKkJvOgML122L6NtehlkD1Dk/a0rXl90tT5hqUU5kfsX2+RDT8u
HdTo3n/RFS8lB413SpA8GTxDkVAe6iowm+z2DVlWGeXCUF8hYkqu3/USi9scQWR2
c2l8uzCv1LSP7tly6CYllw/W2zbCQ9mdJobFv1+kP/c=
`protect END_PROTECTED
