`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S5igvXsmtzRNY3B/M0n7IVBQhxJHDGGLy+cljxMjQyhi6tBXx4bwD7DAO5r49mVc
bDz9M1DJUKIOa5A8KjUq3nXT0EfduNWK5ncQmKF9WUJZnU/j4aa6jFoCl5mTXq+4
kfAbI/grL6jMVpiRLskGvIjLLikqjmGQVTRfET/3wydVo+mPMsiQFETMkBRopOfI
O55zG1Qn/7Hk6G1DPu4aWGaWx278hwfu1g4dOUAC1Us6wYGg8h0Az6SH8cZlVJEO
1r4fwmLWYGo32lLPuFsiFIjKYS7zKffEGuZjwePkZNvqUnr9YADsJau/QfXG5umR
Zxjo1QjYbaBamLYzY0pZJ3F5P07lg2vBc+9Wrla3mwMVpDOmmN55AXYw2WvWaQSM
`protect END_PROTECTED
