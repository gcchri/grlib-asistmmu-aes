`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8iDiH8N+T9ugOV5WpVI5H8qk1Nj8OkOn0rnLOPmsw9QApJEdwg9/lkwI/p7vk0vU
t1HiwqxftuFrFotrmmJTJsmAVlV4upe20afHyXpbKDqiVnHnbyIqSBl3srSNmdc3
EWGu9NZ5sGPM/iYAVEUPrRf9VOfnNjT/WrMWhI9fFzvgLgmRhoVMikRI+qK4l/8a
VDqM6bIZvutCvOo4Rp2vpcbeRlAotTF93QjGCIl2kYB0WvD7/oac/+kwRwycQ2Ti
s0slixvtNaXzCchtH63kiB/AR0+zwiVnrgVOS+k/iGiRl+qE65Q7pgESJrIyXvZq
WFRVlSBFRDY36Q0wzdzUKM4Y2NiPiyci3ARq6bR0QyCgN6McWj6zoQNNjfPIfWrZ
ecTvcHR587vA8q6YtCZfXIsB+//H18h0Lbw5V7ix4VBXdYoTi9mYr722D5cPVoIX
30NfzncdaI9XC5X57xbshc0BMTWSlura2Ss9kojUgTV5gCm2qP1eTbPFYrl5quwh
M4sDHiUsSF/vRf1AVGdr4X1idBGaHf8UCIUHejyNmOmNVl+Nk+MSyVAE4XamCkj/
FJOi4tKe5IN8CPaYNntHahDkO4y7no8EjgmU5slpluHNlQezHcT4PDZXsseDVj2g
k6c9v8j0AP9qmP0Q68Zc7KeI2BgHIGLZb9pEjSB2RMyseSmu/ezcgAR8mwK/x6jT
PgrqCJnfhj0Pp9YZvf7aET88+9yloJM1dJw/kNDiXyWaVMWq9MPMUNscKWAZrbz7
X5dZF0mN6f9g+ODYeAgMem/97bY+Z0iE/CVLWNBXc7hcPmtUWtJH26U0DQPLd+Th
WyJWq6D8w5I6kyXFeTltolyR8Q92fD1wxudfZpohptqXVizWyFvQx9/TABG0uehs
c5W9dB6lqt2dSlcCRWTL8dxvZbGdX68w+Ki+HngzFuftzTbWDPz4weNrwWTRmML6
ChGYVtxcJvzq/40Yho46Oq8rzQPvYuxRt+lpakelvbGVPHevczvkg+5RwUAp4Ytl
A/ru+s2KW1Eb/pmE7Crb6E1iupGvPnGFBaLQXZ+Fqu8z9Ky1h9oyBSq+eopmLCWg
GONjdF/0PK5n8126MKR4l3b+kdFQbGrNMuzdGyHYA4LF2qxLRk7C2S49Q6OyD8Pp
fo41ZdCIug7Q/6XEXUzXMeOi4otmqYu8KKZuWPMwXUz/Y5U/P7NMf/XB4eeUAEcE
dEKRAd2B0DXNCcDU/l1oasR6NzIeO7c0Bbl8K73n409k6fo2BTG2WS7lM971xvua
bTr0W/ZU7bzwZqgVIegkijpoLsLXfr7uSQ9isp4lTJxJLW/qy/2TCiuyIOr1zsQq
NEBf77dHeLGqk/xx+hgnYbKX4xSXlcKVUGgcaANkS6DscA9bU729QVPfxsGGxAo1
77narSpe0qY0NN5oQPvtXAHQyZ2JdeaoXrXFR3P2rcMlJCYwwRijaZoP3o5WVrFJ
+7Yo9Kzjf3p2nPJ2iRiY2x0RfxDwAceyASoiICW8VIBI59XaALGnib2VZE9amvWG
s9hOsLl4yVkCb/xKB7e4ozePrObTzUdWhRJs+dtftBtLQarTZWbgo4LCf0dshI9I
8SnAM3B2d0bP9D7npDdaTUhvulUFVjjP73wpA5XdIZtsHVFEhkbB/5PcwngcV9Km
bwnAAqgBIAyNFxJV7YU30Gtx9TY5K0seElv9FbWakunGfZVoyfwSdE5OxkKlHHJW
+PJuXhTs0mu05eou5Baf0IX2rOlIuDLcfoiToav67a/PZv4lUV+nBcFxA2PXOSus
neqYFrV9dLqFyr/rQM5jEco1tWsUcfQYOxG0PPntVmzAiB/xDSc4sTWzmh+q1KaZ
VjG5RYzGVPVI+ZpAjBYgzrMggN11yQk4a/hlF/Ia0AkEMDPLs2dngndBk7fC4Yj9
P08Rd1u7EkOtjwD2HWDcGnvg88gTXOlLB3zYNTg6PqdqjVXapATz2GJOVZASDUhO
l/Lbab2bWE9nNkifRNdexTm40tWaC0ZK4YCXsnAz2dLqUkNppe2a9NGi/Gt1jBhK
on9zSZOdN0Kw3VY9iHByQAP7SIoAf1Eemt2k6iJD5uS+Xkh7tOKeylQH6UZz79SC
ldVEeZuJqE5VoJxGxOOXtLoOzZ/JHimTasqHgyawbAvQRGRc3zQCPTMVWmnr9lKz
h9kLoMeFaRcInT5S147Z786Gq6+MbM/03yN+gDVba/P8C4ehuWIVTgP3NIPvSlLU
EXwvGzrwmT5lV719n7vDtyYAf06eSLFfnETkSrebHdSnOtXFsqjFAX3jXpVxcrS+
i8dOq5OGmDYQGQ8Zf85IaRDg4SrmfdYXXyfGaRU7Fv3OczTNd3PDQNb6FsjnOw/n
a88azIbGzvzSJSUJqqtCfpb+Ih+CbSXJ7MZbOafW4xOAYyeJtKPEsBMAe2z7YJr6
4QUP9VABo7ueMEXcamreDdK/eSIp2G3yxlqVrwAXySJGgJA3uEzF8BROSUbP1X4S
tr+kLooEP6OAHJFhXUPHkiHgeOfOaJVSa+8VHro5EyTxwI1F272wDpDyjDJulu6W
EqlXd/VIIO2vSfbRTZ6rt+CMmdKtdbrDoUfK+CjFZHwZam0j+XqA4oy43kCYTjJC
3ezkSXuRssZR8nyGGQa2jzqXLwlV0Q+RhIEhzdrd9Hdcl5OeAbUUMwDoNNx8b5dv
+xTlG+ws/Q2VGle1U+9Eu9CrtSD8u85h74xDfrEWOWgSb9S21VE5PynpWc6mtpCs
MX0J8Qihodi7ZlXeeDR4Ghc4wy73kDk8NhEHmcKioyyJx2Eyz2TJSAkIcAVlz9pb
d8lp8YUjtiSPbbMmPIj2RlLkKPkv0+P7uBc6tkImGCWT2PYDstUj7RH98P6KFxCS
wW+sXuZLAOUigYSgVEcZEWy39fU6TzVI6B6cw7hjX9eF23ke7oDoCVtLqzGCovjI
PyZhGFTbse2Cb1Q1V39xIvEwsyc7xHY7JfnoMzRVtJdxanWG9H9606P8BxA4Vbb9
Pgf/UHdjP27/E1+1mxnlpSzypII9wYHcAZp+rAVoM88ZVzXTR8GGDoeFZNYmwEI8
E4bRCFEv7IGWAnR3jGdGI4sFW/mhIWMPb87iX0MgUPn5KYt3iTPycfzRHIJoJAxy
aG9ugO85qcAmVw0IEUBGJJqSUrz4et3FhzweCSTOiEn1MP3gVP8ECR7ICUm1e8NL
yybvdm/1S8rtupS3sZwiY6al9U4zP9kJhnLSiOVUkm+He+N7EsGUQDf+yY5XPfbK
SzPg+RTj6KKorkb7N272Pn361/iptQpmm6wZm6+tP448pwSRvgDyc7OKRh2wpi8N
/7UhNw+eLR4DCfbvRKod2kc0FZGbBaz1G81yGSqX7puzES7dDZsFjKcii5wyjjeh
SRqb+pAaivst8Ea9uETeTAJ2EvW17Zb2bzUkSWw1GKJx+AU9NRRIjultOTR+uLFh
FJHWG02Ulisa5JOO6hjJDXfMU4kowQO/5KoU+fSVisn8TiVM6GMyrNMSR4/WK4bd
gpVwngLWgrs1rgs/TI+fRaWHqYgRvbHriKuYBF1irihW2X9Occ66Wksf7fSwzAAB
AQ0e3EU0fKF2q7ZMHZ3g3ngmj4rQw0kTo9tzYLDdGuZw0eYf+Z7zK5NnmIz3x5rV
FLkLytTTFK6kjGtatHXIiA7y8kau53PRby6SFhizuEgZ3EnJX1Mbvp7PwWyBM10T
E8BYERXhpR+BJqF92rHQCrj/cf4jCh5ljxurkfJVQT5JLFdlcS2gd2u4Uz5WWdVF
5BklC61ReuoV3M2v7srw9hQX69jnYpZpG5YA6sVeyJZc2vlxvz+ZPOHOuWE9UaJM
lGnC+X5S15sBbRXEC9Oly0aPHvBVE4lVG88Pm2Jj+YwceiRbGWqN3dttkTjTGB4I
Jwku1QuPuG5uSBNGzleHzpfQoNQTsgP90h8mE7kuMDE5r/udEasL71w+NDRwdyEM
B1OUCQOhjSiX9RUZrEyr8RPQH1Dv1LS2wfZLLZaNx3Fl+LgV4PpbddyPmyygGb1k
gdXvC+cfpCary7eytfEwx8odld+tFLr+8QufdXjhMD+QZtOGBIGTRPTvbk9iSP7y
px8UGWVqgYQXu1ROTfy+RXcinGi++B09DWYxZ/4kKFsDQOJUeie6vRl/klZ+7D6f
vAm+OBAFpZ99kNTCQ/rq0E2HOOTkS/K9Rd6uNpHOtsLFwOYHmREJBe4bQjNNaK0J
nMqSeLasKvTc92Kcyp8SFygrnPw+N85YFCJq+6+5v7TyprY6NQH5GvUdPPCxCmCN
ssserJ8u4KaEZ5hHFN8nURMtDmbdGS0nS1dWNEy2542RZD+ZL/hX6LgquMkn8+/d
LBmbEGZIrBsFQ3Jy1ySJhwlzuK5lU+TvRNlcHy8KqDws5XOcY7Ab8XZ0DuGLDXbD
TZU+lnyWEoe82cZsvTNbctQ/wlX6GB92YruNEOV7In8aT4JTSfvezbbHgKQgR5ZH
ktWhZgG1D1Ru/TEvn1e68ci3TInimNZRq8rHEzXtoS28uaT7D5OXKJLYFtEUjxVF
8Ckth4EZ44dSBP2a2mTztiyfMyOpI0zzq9SmAa6/DnIysgYmy24v1JDKq7NmZBFo
sy8qRz1dFOxw6HM94ylF4PAm/ehHszzFOI6V8kzI43TsEAKyLfiSxCJwPyXMEoGP
1FEkadzxc9lNoA5C6eNwbJd5kP3EEwMNPuYIiZSt6sV00Kxbf6ONGYtqh0Y6MNEC
CE9Lh3jOA5SPiR0myCtWOx5bue0AiU+lCs1XXZfvGDFiHVl4jAFq6OPL879mlxnZ
NPBuS71vZMzghR7L5irJdVFDMGJHCTyfTsQrFOK4gkH4m7Uz6x3/UDKg4LzJUeR1
QmWK4tnQF79pEVtSPB5U9FMHIwlnZCD686aDnAnbNLUqpzlMpv+k/RweNB7vnPtG
/Y+MMfGmy0E2creXn/NcY+MS+nHyF97xj0wn8ZsKCLNUn61SYLQupNFVvOijnQNM
tg9O+2WoAnMTQzOJByaWTz4cQzFWPxc7Rb46Ql0btvYvfdRrxBCXJr5UzJ2fBNKi
Gk15BW7H4zZNhVwSfac5nL7ezqkXPZ2Ci8CBrPJeCFCW/j8dqYTxLN7xqVboOuF3
LLicTrNStlaEUyRFpufG6gbgK+HSFNGM0I/1MTVmN9AqE0ETg/FMhrf0kYhkK5Jz
QrbI+n9aIepCM8T0Ki3Pu2TSvLs4hkJvfaGrSEzUe3px5R3ou3Otx44U+EgJ4UEq
AUTY3fY1VHXarGMmkjtbrOy11SBbE0gaiYRKgDcYcZuqy1DyMkyG+ZzyoW0DOPHy
fypVACzviiFgnaXKTCW04kfPuyRMYy4d2T7JOeED29TRALpYlzevC8JGtcoLaY73
SbYTDdZI+bKCjs11w1Dvym3HD/bw/WGPQwZMcsuux/AiSimuEVebA4K/7nDvKs85
`protect END_PROTECTED
