`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t/Y8e3Brlf4mGHQ/rjhF6RSP/yAcfS+b832Ltkp9ywDHEDGi4xM/oB38ywQENTyD
TrhNxvNwsfkWJ3eXkHCefGR78KazOZoCDFXj9iOAYGN8xmiI1us+CjtJQ0P8CIES
P8UrQaJA0zbIjmxBSgH4e1VAFa+0oUPyBlnK7CvA/MUsHEToCDfp4JGcwI6s9d6A
DzSh+yS3XjrJjsA30HrraznLTreXN/l/qISUcyMWJK8dMZ0djjpn52arhK/BQyzI
2V1TpKIPeva+c/RWfrbPxho3PzGQQ/+q+8xGnEnj4OhJcZSlYtMTl7yYRGCmubut
LrfkRPWMFWibspmSQ3q3TWpe+NQXv8ppV+Y9mOcbEeGK0AuQKDJpgJRjWxmXF4M+
juWzdYKpAWND6OOFOjQbYi7dWK/EkQiia/qTMuDMk1iljGgO6VixItYYaD7iKjnh
bisezllRU+brX1oqiu9I/Gqj/zIH41MGbJkB90Aq0NRZgilVRSYoaCtnHRlgODCM
UWrnKg86vxOS5GmOSvTEZkLY9YD0dWZXd1V6iHbiT2vWvsnF05Mkm0HquDgSHqvV
ppIh7tuoIGiJ0jftgyn0GzqlyowfE5JBjnj901EwIqz/7GK961Qef+0tRLXuJZzd
PDZVFwpmoYUA2ut4+JNtHxPMWcvke3ni0+svUC9BjJ022nIa5AgZcOhJR4dj81IE
in4N6BT9Ja1V29Nd5CMhrdeR1jd7ab8l9+gkptIRUOALGiHuv/KXIwtxX6xShTvQ
xiDtzmy2ay/N4u1GE4VLZELGVRTZrDt9Z3Z6aFH7yJk0XHuUE1WUkreYHL0ILDOq
j7cd1YHB7XlGzCSRLA4JDdq0N4ZbvgIP7IHiis74jyr4VvTsZLzhCSCcgQJwAp4q
UfTmZiaiV9/v7v15kWP8Fo5sG1kMLXNS+6+2nXxgBVDNLeVQfIX5cXS9CHrfohDy
2TEr5EMt5Fz8PB6PIQLxvUZmRvUJLE3hn+lnhhUooVg=
`protect END_PROTECTED
