`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E48+ZPXrULumDMl4Doq6Riw6hiAArev9fPZvH7VZJZ5WP25CzwBu32GVxAAbyQq7
Dnh8vrpTLcABeqGCpbTDSDzWrgz2V8waED6wimjU27F/tT+ikQyNpTjZvkhT21ry
BXfjRPYo+vYlIhwdBnkRCLK0YZFdGEp3Hz3hwvomGkhWduTCV/86VTGAXbIa0oqQ
XzALzvcaOfsaFDHxozL8YaRtlGCab0EtqPXlsnbZN3/sEukWiHH9AldkS9yhuJ5l
G9QIXbs39PUFsqGjRGGh7D3VvwywlIYkOSfgY181uv6b/4QS3vC74bEc+AdFIa9M
P+mixgTFsS1joYn/OZLtkA==
`protect END_PROTECTED
