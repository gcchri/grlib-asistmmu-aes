`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G2hohVZE8bjsParZvK4pYanf5urP6CHCtj/LHe6sSobWep+35XgDM/Q2/48BZSVH
O4G0MM/fLP3JE4Qg2Vxe4U9n6+ozoXbg1gOZtVB9BoAdvGDJYgBV1XRUb+Sw4WDy
A5IkAWbpO30n95DIgBac0ZoYfHh7e0W7kzEr/3Q0uj8u4MfgGMx4Qi3QDpi4qdJN
JOdrVUnNtZBXmRoeWdjgzwwKSixc/Whz9XRKvOoG2TMph+GV+aGHPBN07pOcUAMp
xYf/H8cZCmbW6cNNjz6udh2xpaZ1unAQ6+9stm0aMnJebLccoo7XHB90HdZNu9gg
u/Luf1b6rk+mKwr8cOCX84REv+8KLOSiuZJ8xUep+CoEDzm72JKHwt4Dzlz2IfzV
2y1ul1QkJehlzLHJ41G+LqqEF8rnALG/Wjawn5ChxRImq3cdw3QApk93eOPxvHU2
mIzEzFLCyTezNLG57TXQskW+7+nafYnUS6zai39JgkdRFlPMMGNjgbjsL0tz/c35
JRirjrkU3oUBItWYqxZWlAG/Rt5oOuohRsKrqIdCpltljhuI3ORffUqukRSHiL59
M0daMWEIV+5nEfkZmXJpNQUI7RsxpwOLq3NiT83S1Z0tBWKTfI4LpfxMLdknv89o
xbf6wnuYrkiURaNKAK26Ig==
`protect END_PROTECTED
