`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cawngrha8uwaPolku1vqs4M31bB7lF/MktiCiaQb9PJCrFwrmY18ao7DTWghdlqd
AUc4WH/d5G3AhOLmxRTO3tYCzL4hLDLgm6qxecavj4lanKn1iq4oFvPRpbWJ2X/X
UhC/PInnhPVyRko4sJi6Oa7YMBB37ZW1hmaX5r7vAYFXAAGOuCDRJvWU86k+1xAw
3h/yLL21g495EynbAXNPi57RyMl8VNmldD5gDUPJ0wJaQwo/DXu1HP5XeMlftVVT
KlgkXCdLXlzmRPdYIFjRT627v/7NvavAmVM7q3t26dYgu4Uq/rG/i7f03nJs3Aa+
lRI34TzoxBuON0hyRvHGV/G8gnpukGP+lU2YV2EBktUTY14irkq8LzQI+MuU3im6
rvVZtAGbqoHNpc/fXPtBiMDEMwKbhW0aLhkLXur0NJSGF7AsxMrXumzHukoD90/d
vmV0EDkLzscwBOc+kJUSRinM25CpCk6WY9ZAWw4tZyU=
`protect END_PROTECTED
