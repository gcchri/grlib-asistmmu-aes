`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RRjc4g3NzkO+4bmmFArg3iV/MtMTCsz4h14QKB9Ust2cBiMBNiqUIfnKQagnf9x3
FVjiIthKY1wooKClfFNSUsWIn+DfVfdWHuZypojYjcyjS/Zg36TOBNDjW+NLjF9K
difezgjObtFh7vV/Gqybzpc7h60bt0HTGjb34t6IGDjwMtNataryttMW6fCuvydt
5FtsvkJmQ9LSv94rrxalT5XgTI9iixcABDPBWN8WwvzMVXWZfbijJpFRITeP8oEP
SC2P+iL3CYVggMl8teFN8s1VT7ePDXKgXDj1Zh3uBUxOQJoMNASDiV9U5OclvyG9
XxAvz6YR3iWBbSmLkteSC5iaUN3u0wgUy0l4kDVEzrnkwcnFnwltdNr0LaTtkBz1
Cit9sxDhwKy/f3lPUD9wZRPZLrV4Ruk5k26cD6/o4a1kEzCwoT7Sn5n3jUJzgoaG
V9ifW+4BZZcbvHX3BjD0JI7ojf6G8IFu3nHhHarJEN4Qs+cICVY5RmgJx+xb8wIs
nVu0yBYNRMGLSXqjKZx7H+w3EnNABBhA7yxKLKblmZkUa9Jfvynh4aOvVJsrNERC
8noxFlSDSw84NA8rwinjuYrigk4BsWUM4ZlMg+6KD5Nz0fi7FMZu9g0RLkjX/SLJ
mUMC+hrhtryQ6OL7AziJjnAHU0j8RdGjKeZE1ntOcsRYzPmfCitzQ2zlK0dBUR2H
`protect END_PROTECTED
