`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AkFregn4mw9BZfCwtA+p2nTZbGQSvbBuKFDkdBh9uPfGBBsy7DTJA5FmiulRq3kA
SFUps6b3hF5n4yz8v6h2LF2iOTm1c6TwUek0VXzgnocgTeRnzZ4qPuQZHw6QYRBM
ESls2KEukSxFOJEhBv1MeTePCfj062J1+L8dxk97/QMtSM1HiXmgrAWnpZH6fkh3
XuZA1eM9XKQoWC/FhnprhG7+iypxvCTXGbhAaL6jOq12tmkTwoS2KFh2SCvpwqpr
uBW2pv1oIdecExanEwug6ZZl0KfnqfXMOx0ARpK8kqomqqP7ugtPbsaG3H0Vd4Yd
tWtCbZ6FRanJ+pWe7PAlfsWkpqPoUJay6+jedukooQ24Ec4xzY/UeBYo3e3PjY2Z
zPcYbFpYdj9EF2T9GnXu71HLUoDruECxSDdlS5WSyATSTR5W0FehfbK8VY9N5C7I
WXtrNQBSaUJRGuSViNjJg6jnskrVFWpGroBk6PJruM+0H+Z0nSFV0MVBkIAnF1tQ
`protect END_PROTECTED
