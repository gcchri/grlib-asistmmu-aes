`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EMGk91H37R0P3t3kGBGlZSev821ssKTs6ZzcoTXy9/TCDJLbeR4vZx1FjCUurEVP
IJw8l/lxdWPP+7UROxrdH9j89Xt7JAhCnqtuGCrIWgWJ5Lh5BJQ7BOIDSHRmtAlY
Ef9BZtBMqPIXpp9yjjcJHowPSq4rntiYRvy7RQ3K7LJWiMHDFafoPuVb/H2iBbKs
UahXCn3yeZH/+251cuPUZ/QjvynUD8mltTn4hoEv7j8vHIgRv+zz0RBqShzRxh3P
bat+c2rrOZzYWwt9OZM2bWubNjvsz10N+DOc1wAvyghkkMYbPonYkuOLPkXlIW2n
NlR4S+BXMxRpZTXv3oriko5c73IuhhCSQnbv5dIe4/Iiynp41QCNy9QgBXYlTLDY
`protect END_PROTECTED
