`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OIbRPpWtJatPpwNm7FqShGKkdd5EAa3l28YLfF75drq5F79etT8AQrtxztyNAa17
Q9rVAJbSfMAcSPsNhj+Gu+d0SA5Anm0yAsut+1J94EKUrrsgGPjugogt31gdVYng
E4CX2gmW8/+NoLBrrH4ttQ2StMgGigaJ8oDN2+8g9IgHBLf8Qk4UhE3rpaViRgcW
3a2eVJp4rpHNuO1m8Psczkbgv+4zlAdP4NLl7fekk3wt8Mirq/qqh133A4QPh+5g
Kn3CeLC8LP/h5VAAi5zYcM2ksjY/Zwojz4TXPmS4ZaZsID77OKCztZTd6OIclPf0
EuIT62hRE3G3fohZ/TMQ+r/F8JwLVvHgSKExNcy0xhRhsOGOQ6u0PQORAZhCmhGA
hADi2r5F6tzVLQeig1KV8nfvX98iQNCDXn4l2fRUkrVwidV5U+BT0cDAL0zhOWOs
5k15gBE0HwgF1A9ALHjW+vmTZLh3UyngejSxQ33cEV1Qj7I8WQnmEyw+dpbL/tv7
3+MF8cUNHk0/dzKdlGY0mJljfMLJSohYieD/h5seYCs+jRrv44hqQ+hbAksmgyxa
SbuK7jzB54kfoBtOPAdeT4Q0FuvILhov/53fVUHXRlG25ah2mbYcOUnYbLNoWE1o
eYyF9EWEIcyiNc1OH+i8xsc2heRyTUJPSIxewP/BGBJca5/Dav17XgE+RfmBXP79
`protect END_PROTECTED
