`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mRkV+9dmxbysoFalmLrG4K3jjvfUFnkE8rk8o5Np4nksnlo1BarwPuRN7J9mGOmk
/mh4gcIWgneHfjmD5V4992sVgzdBtBDdIk//FRWDfKJjQCrJTDaObHp0XJHataFQ
rbMAobH0ziODzJC+q41YI5WGSdnJOds9+SuZvSlFodS5y0oJu1n4vXOU2GzXW9QE
QDDv/b0AB43gwO1DQsGFrpvGNuaoXYYBNVj1slAlg9AQe5J3sYEDgpXzjyW8OKPY
4L1kZ1ulxhgXyAkKTYqQ0qvsoxmbDJbwg4yfrO3CpsC44Ctl4sNA2hXOqrOyPyAj
zZGDeGrbkdyrGage2oQQXk+KhsNHpiLouzyiXJRtrNk6aGMMJfwVqSpyaSM6Vs1V
67RV1j8HxVcaR1CCwVnKSCstG+hjCExJgz4MWc1LhR1YQRG0MyeZlP/XCGjqiynu
`protect END_PROTECTED
