`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mU5v3JWiKb3KgV7Tzz6BGVCRN+xmbcq0Cr5O2F779j5whzZxRUjMrdjmKezO+FJV
ftbRo+tOe7jt6tj0BQhx/HMjD5cIFthTNcrGsvNXzj4GuT2yiSY5g8lhf1CgKS4A
dUI5pwmnAk5He6A4FoVAEkJwFAuU3e3HwNITQWwd7eAUfHBPkwWdc+3pYvnTpqM0
YX5mkPEalxRV5TB9fsZc78dFeft1EjCm20PC9uUOHAQ5iOz4JKZn0YW6lpLfkc3U
qpxtxW23xQKfSV5IMNsa8mvl2UuCP2s8tKFoMCmieJZISzCUh1hZ8/53q2bByxpN
AbO0Ca+LKhNd2R24iJq1osiHT9x9hfkyjCGxB7ybflkMIzibrDdXMwypNQ6i88j8
47f0IiQ30nS+/ES5PaXRuKi7wNUSgR8No/+fnPGv5+web96OrtGuo4GiXRw6XHjR
DXDlXNAFTI1FJbACA6trYJQBCfYvGCTB9io+2rhufBY+zSsGHt0I3cPlefWKYwfI
dgBWoysrqqQNIUTdNapCqvgCAT8UsbIi07T+lqi+w0YhbNln2rUHFhWy26hsW3NG
Djml+9li8JjTfj/IQw6akKjvSBFJ6CFD0LhNzYALD0cl42MnLLqk1SdrzzAys22B
ghL+F/OdgwXvRz6qF4OdgzqV66Qw0CE6tFnb0P088Pb2OwyA+6hARf1cxXLGB01d
Q1qH9K1f+yrle4uWkxNVCEHuE19QnDMFgvqPEf/vBL8xUXLeKY8t9IeUI58LhcoU
0USVycILTUWrMheC0sb/ODFcUIAVuLeUWZPavQeMYIwgTbDIO+KNZ7AOv/yNIBvJ
Pu9pySipqfxU4kVqcfyRgaBj8XWfr+0v8TQd63FPw0vmkZ4Bwc1Y6GRvHHj7SvLA
zVwz4TP1Nz6gP0v+aH14PUhRuxB/Z8OEELNd4oPmK2TQoJXlIFNIQ07N2qMAx0G8
OlwThQmwzq5YkS8N15PuzRbJLgVl+meLh7Bl8WVQUpnJfdaSVMThUX/t8d6IoxN7
j5t2Z6/BvKUGrYsmXrY18HDWYqAIW6TqlT6zP6+KItYWtgAtebqCu6eiM9yKWI1k
n9MuFXbkZIPNLoLwWLZ3gwcARRfBXwP929GmiS+jJS7JXhqbaAxBzl7tgPOSwhTt
Nn8UahC7+SPjkbDkEusiHiERcgiFUyZfieGGlABDizhE9vHIyv6kmA/xRHXvCx3P
aCK6QSdp8R2Ff/Gr2jRoTeGgowihCJ7BvE7D5ioSAL5J778M5Pc694ipAdE3E05n
e5BYaWoFLb8khlmC0QjC/4c5uVBdHasK1mM/Ffqv8hHuzJYioE6hOq2i62UBIOkd
nr9pEM+Y56SMtor64Hhz51GY2nPFT0/J/SVrRnBThw1cPCqzqY5wz9Sd/sbu1dJP
NAnAE7E8NeSSc4dE95DG6EHW3SSepcR/sNfZXA+BggM2UNIsa2QrkZBGc1YivAVl
euQXSubn/hPzFt59l8x0xmF2k1aK9a+RWrStnRh9X4fQsfgRZ5frJoV9jJoftWHd
B+41j6pHz3pyYKYxVeCX5g4NnGmV6jiBirYZXrgiPSEHLGkhOYuBjxyoE6xFZfMV
tNBeLFVA2Ot1B96aYfC61j9pqkDxWs74ISJYvIhPlTYrntQTzWqDVwuVtCp3MwpR
rAVsTGjDNYFMGC19xNGQ2nSQnycHH+g32jcuFj3qTYj6lhPj5hLDBXGIZk6ArYya
O5q09EEIxP2aQhhNl/ClGO0K+yxMoT6ZSVn1WrnBUs83qpLjGOpvU0ZqOSPH3tGU
vZq4bdauuoFx+gh3ZdAwOxbrRysV9jEfygpAlRI52hKpRHXHHlfHH2fWTOlJ8/ff
YAcQ0pYeXnxDzpEjkLkYLiHhgfTQRnNfb3tbcgHSwgjkCDq3ehnsahQ5HhEbggCo
8vMHzCfAYbB/ernZ088nGYRZvn7O5hRhAqH8zG3ELEngseotkTJGXVi7R4K6ZTCG
9v69mctzdz9Yd/f16hljMKYKV8eAzhJPd0wk6YEiJcAiCKzU/xOQVweZBTy3bxLT
UFusCddD6XiKGtLPUIKRpfkVA/XmVsVY2Ml6YtyOASrJB/xA7GRUPPxnRrNBK6BE
NEQtpFJIr0MQQpTWbHn/Z4Z8d39znn4eAcxqVVBNBnnAZwC+YIfGJ9ooe1c16yJt
KYv8J1loqmaAu9hL6BJZznZo8Lpv1buioODXgUWB2IiDUNwrzEvFM4q154BcpfMn
kntgWkjK23iBNmECuOGWJ1flfRncl1+o3buIwZqfiR8cEgxkYcZjENQZO2LZcp6M
j8RlAAzblfIn9svoEbjDPU08IOe/wwzeP5JDfjHGJGfwnvbM2tcvP7unxB4CCsXf
9D+ZncdfD+qlvGFJQCXsEjqBkJ2tMsZc8irwVbeRUPFtXbMsGblNIMmfLBtJMZEn
0nyzEGNP65S5L503BaMyrIMgS09xoEe9haJgB08sTXLZ3aT5CrlLBxZDz5uX3GTE
515fMDO0i+oNJrTQiOjbtpdsZqSob42YBVgylFi1bxO93OCGYp5IUxUQvuMJe4rk
/eAERKynwh0hEM/43F9AllodFrCxHUAxV1snqXaKl0IWiu4HYI6Qtib/30Lv8Si0
tkJbej7wsYZ/i6GmFwgR+w++/fjTbC1GWCZnGIa1qOabuI8vDgA+8K24hfr7Zb0d
TXJCMxVHZxOSnDOxD9+tW8BlNX3gQTZX4pQN2iz4XFG8xVcOOG3hsLf4mbaJR+Tk
WZnmMlXoLaCAYBHvTTNbje3rqVkxwX7aEqXHcx00dDTqNTL1k10u2nxq1PmgZdWa
Ye/iL1K2qTsO0oGet4lKRvTHHk8aDh26PupgghkwOfWuiVezi+DTfgdk7dLa2hyE
lFZJwJKZ8hF/B/jqSqiMKT+bUlnj7tuGp/jF8No8PdZGpNlu8murKJ4rX48Q2dqA
s+2TwqWxzhPLBNwCapRjllJbf4Cd1OZrVCfreWUHnJi8Nz4ihPhYdNhTr0M32dDQ
tiklkIKemwlRMsDL9u68vcI+hhVQKN09A6Ko63VWS66+Kq4+2lRRokCNm0k0O6Ns
KQOZDuR0byoYobM/jD2g+U+oVB0P5dY8y+c7F4taASsOHQVDBm+upvEpIjKFCgHw
b6aIVaVKN46AkV+BKN3opofMBjuiHXR6udkQswRWzl8NzyRzDeNDsIJFRDcBtlkH
rneCZmyglmx9B8ILg6XXwWbTCVRoUnhVUSQdThf3VEmoJgmPAovItjdhMPvBKCLU
7yOCzEirJrgzNLnlFYOjXvIxY0Vxk72oVVMERp01v/w3Mi3XiSZisOrpaoB+VdKP
wVKDddpEZ05pjj7OHufrxrIZ60/9tUEXTVZx3+ffLuygI0IOje+IdL5OyPDwHxJi
VOitrygWY392ook17sZicSfkY55KcW0F8ZjreTtBmfKxnt2bnWsNoCxjaTm76M1d
s+RRfijwQ/j0+EOwxCHVBy5SvoEROJHDkENgN3c5rSJ8PbeHSR9I+1EUbrvtAg2n
BT2tud2zotmj0w98UJE4KCxvqyig1JlhZY/maAOU8h17jvX1e+CjK1BEleD555MZ
UejL3BEAihrmzlWj3NB5HkBG3a+onRMYyu2yHA6BVvWT/jicEN2azXdB/hkAGwgJ
xzsRQiGuG+RGkIv4/75wqw==
`protect END_PROTECTED
