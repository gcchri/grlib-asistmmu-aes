`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wofJWllochbGCxcDwmn6Ar3v/wn2Fg9Ap7J7Vj7OchNHcwDB0Ll9d2r6JEEuqor7
3XSuTX+VIXXUaE/nHd4DWQDmUVrBLwXqMqxsqfQbaw0/2kEIZlUTqqSXGSxDucjM
+xDlQXPL7WWErqR+6BHqsFesFlxeQBtfyoNrjtQCiCDoyyKi2S/Nq7lNtNRUVQep
HqHM97w8OmNwHSQ3F/m0xfFmdnqzX/5E2KL9LsMXqvWL94ztnVcR1kNwjPdZ+DLw
jtSH8nbT8EEKO//5vojNgnxI6P1Ox0MxQlE2NOVFAjVze7vDgzGXXDL9pZlaLCxT
zrAK9UOpruIwV+G607hq4l/BSCz8bjnAN47FL+qG0WEuaqKnN7oh1NSmamS4hobd
X31HifnT4ljgbozX2ggqOA==
`protect END_PROTECTED
