`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O6t/bxB7NRaWKxto9Aymzl7qvA/SqVANh5NaMBLq/XY8+clxTl7MLQrG02J/rWe4
MEPRhKSe3B0ht7zosi4/WflCCY3wkG54qrI/8mGPcYPXg+lPNFcArFFd+jiRVqgv
446FuTGmG+ezkdKzyfz+M3BTzkxTg155nUmpkZ+dBXAjuhsS3AQbOhvxwODwvVXG
xIzlZh3NB6aF5GycTzuKl0QoXr4FgQ+NrOwLXyBWP++o0FNrd0hSlbCu36hYERzr
+/2M0me390h4/cmxoQW4I+LmS3Ez2iI5BIWkgiOEyyYi0STXGhnBgi3Z0c12wIdd
ttt2YMBgUHiV8LHp11EjLh0uLbKWnSomcpGQ6a/bij88rf+aODYvlrdMaQPi2tA+
jk3jwz1ccGuT8+izuapzMT1OPIoly3Hiy0ubglYUYbTIl+73oCRtV6GDV8qj/JRb
1qxKaZFRTAdX1UwlwyFXLENjuvyNTyMXmURSDzs0iW3qSGs3U4671keTOqcsbCfY
`protect END_PROTECTED
