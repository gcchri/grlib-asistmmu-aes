`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Sjt8Q2N+sZnUuK2teYH5WEGJu7dHqtZO5cfkckqlSKQ0BbRuHfw7I5PteBFaAOn
7PdgiYkmWbhj/yrS4yGUbhrn0B+WOORAM77zUjVDxspeCJdA3k5eJ2da8a0Th9Dg
GtodvlC8yqWuXloVg4to3I3VgQdOCABifyujTEkfPHEarjSWq1kA1dklkohXPVmK
W4KiUc2xIILI84Cky9afoP/4YtS871e9fjBE9HOQ+Uq1EOJbRbjrdm+91s8zc7Fj
PcydTBgKA07kZtBX/9Xj0H3Vg59rOqoK+x4huQvBOajyLPyVxzoUOIu2IxKUxvVT
w63a/dahaMFvHmp8DUp8EoK+k+iSQ+G6mqfnNF1+YzgRLw/AeiZnshvoq7lnxd8T
dWJVnnXqEGlfdWhw//inGoU3++VQyfh0GQYS+WIiHiZDVJiuQK72qZXd7y56XX0R
R5JPDQy5FhmLswRxv7RVqteVO6C1WU7fq+zYZpsmG87VrWp6uhByF6wOx7p4FV4c
tv1v+I+lMTDLh4SLlNai45e5Ew0qldeNeRRh4ZxgRVvVTtDXTJ/23JakxFEYI1Mx
0I3r3EtWmlfJ4Ho3Y6m53qx3wViqPcVwuXyHBnqBeqZFjfnKck9VIbrwFJNNpixU
ph9/RniULhreEzqzXVpIMsqGZNIqkpAVOlz2lgpOK/M=
`protect END_PROTECTED
