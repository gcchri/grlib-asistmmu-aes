`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zu+XmcbC06yWEOm9CIiFkU9sFfYrVBmOkmwWs01BLlEtVkDnvtsytgLMYZnycbjT
WzSy3AfqFDY6jiJQKlIhQteQHANCInzxGTS6I9ggHEBUkYx3TmjbjzsddxQkf2xU
+1adeJxgjA7pOBBZct72L1bI6aJAS5jVm1AXH0o/WjpSsQk/ADs2odkzL6UUUv1W
o/hFS+RSkPfsdKwJF6z2iF/OQL2svh/FfKsaLkhNQsJxVMYqZkMivztpOtHihB5m
cbePxVQVAnYmXmMpJybmAFl4ZG2ogOQmhG5VO7McLXLRj/4UxMYEy5ZqXaxSpDPh
pQh+SV4Xlqn9jOuS1fwvhGNxd6ubUbuk6gK92AjbhIhmLv+Vf9Dqp28U0DCzKqrF
A5IXPf+oeDncD3mIp67YkovHxmK+hiDR/6Zu5yRL4ZSnnEZNzW0MWliSeM3cSGVu
ArUBvT7Jb9yjGgcSYW96PQLZsICo1ZckkkyZRCYuW+J/DmnPDMBMZ7mMVaYLLVE9
EbJvNefavZtQY/eoFkwwkCDtoeny4jyYpbFpHqHcXd/rYoMn7mujrcZz2Cz8/bH9
Egx/Q1Dw8+x5P5U9bXfYnf0Lvk9AVWRdKbRSUiyC+W2VoO2NpVJmHor0N5Lkxmdf
rHfgwN0eDur/1NhXTyzcPbVg33Y5zh8A+9+P1Gp9YebimsGBleINjTqaAKgyzN2Z
8LSClEgOoT3Kq3Fb448kB/3aEQLhVgt2WCeapS5ydONf6UvlXJ3bbo7CtHl0pVaF
4w8yWIt3Oz9yZXh6WwdshkDR/Q/YTixKALq7NbvnB5yBy20zClbXsmTX9F+lJsnT
1YafUPerLZXM2PM2xSMaanjEgz5Fzl38H8JhhT9+Ww9VjFWBjJhTdWc8Xhc7FG5A
nSfHOrtSEKfe6RSUqGyu0konEMUcGALITBWfYhSeEC2u2TAfmnsZVFLQCQDa1qk/
kJXAapwqQPoJqFTjRBWnmVLmqZNg7mnO+PpXymjm6CEg/K9tssDSTHRJlJx8nN3A
3YXxJGCiQ2pn45v3nobnv7F8d7XLv5LTe/Qy2kJqCOGrydlyY2u+gqD0ak3LwleQ
wTONiMYKlPAzQRFtWSHNF9VQe82MxA5YO1Qt7dcDBA8C9Yo0+DPEkHonjVErrVY+
0uOjK6n8Nmf789bylzSSleXor5srDFJO+CRY1F3uK4KjSUptURXlSQkQ2fLaI+Dm
2WaeS6imU8hXWfq9OsQL/RJOTtXttxpz3bayTmUNGeyQ2JJ777r3lO8Wg755WEaq
Jgy/9vOQgDKkqv7ofSNJ9GjjDcysDou0LoWd8e91J0xuYHX1nz7dwzAo8oT+4xD7
dfzGI2xqf2+04huCjDggYLINZZkpTdbiTSj90rY0Erq0lYfATNAj99CpKc7UMMwN
bXM4pflZKB8lHtPSLR5/f3n4vzXD9/z4csQCZwqBiK3BqbS1Zhfk+yfTM2sRflG2
roPrcEJI9E4cp2aJRUHWkUeP4TV+O0ATzWucnZQCPYc7fObzg9lMmezkctxuDhA8
U6Sbmk0rHgywGJKjEEQfzNcOHMHQZSnh1lV1IEMhW0t8WgSrckDOhRT6dSXohhCC
SS/ifv64LCZjr0Y25OixpdLTDPNYnetbXePkFXslZv+55ojamN2xY7fWD02MTU4E
4bkZqO4LBHyAeDt5Cvgzm6Do53ut91XCE9WSzepKOwa/dolobsLwTAgW2ugxbXLY
BdnLi5fXo3/KYlaNzLTNTUoSTyOu7OBsWFVtK7+urJxCc4jKRJWPHVEKQJkjFAtE
x13ZIc1ni0erh2CqKWvVcO2M2X3wdrvBnVSbrKOP9QO+KxJuOGn8LzcPT4IG+mJl
VnjoEbTY9GzAUNRvuDQJOBxuQeEz08Ank3ymkfE4O9DimAOlVPqpKdbBXnOfK409
8KMUMFNjK0C/KfDHe699NB78j/NKFI4QZ7rYeUE3eBfmZU7SqN20V8DEZN7YTO9e
S5OLVAd56wwVjWcMJzKQXWoOJZaxrAlRe9cG1rnFIDUxdN/Ds56bPoto5Yafptm7
LwBhX1hiGxDFJNIGL9BTAcuvdHQM4VHHvG7h2gEt4QKwtmt0nrv+bdu45kIn7yVI
+ECf9bUkRKPI5knGCyThv6a/SJFsOKvh9+8PL1bIOVX4G0TBFxgOM4FdrTBtk0Bu
sKY6Shc761wLeoI8QZuEAFunN4hcnScbQD4U2i1DM5GnyfGVXiY930o+LHLiGOlQ
fh1mWkGdx8Fq7z3e5180BiSZsZqZOOemOnA5b+wQEi8jImG9yBRfR4xEhMWKPttV
omJlfeJ3UaIT76uhIXcfssR7LxTPwhrgoZQQCR9C/6Ug6Nsn19yhEqk2vDrhBqht
40PmSXwu7EPZHAYC/9I8qj7o6cYblnGqcQnUIRydLTsvhfae1o1jr1OCOZ9nsBST
jhNmxewFbYoM40WUdyTrfNZqEBP9aA/ZJDwbSGIYKwXwO0w205Q28EXCctZDUAk3
SI9xyrQR3rOYmUoVvPAfkZBg0V+y5kpe1OrP4L4Y0KKN5iW6eYYNRMh9KLv41Uba
A1yC8hIY+yMVrmLi+XsjV21TiSJajVuV84rni/NCKocn6t1cACL6q1l4X7vBYp1D
6yLgFmYVjOVrRdk7uRBxYwQzjD98ta2EpoTW4+42ql2IA/wKeZdqYhE5x4bGWzUt
E/+asjkjMG7l/5sxABu1mlT1vvBlht7UpnirvDWRSSZHVLseAe7mXyzLMch4nr2o
ztUPrKhUXC9Ll9COahiaEbs0xTHywIvF8BCol+Ylt3mKF+VtKcuasBPoe861AWNk
jCGK3v224Tuj6fIIxwhFUsG3/nkpfWhF0pr4Xbb/WWNbHy0AMPm8ZwpN+qXHMMeo
VXl+NPp9O19CxNUBxDjupPzRDafKkchR+OBBSZ5YeSCD1IkEt3dEBfOlXNeWiwox
PyoabxQSqyYTuu/6dY9G8N9CHo8ZhrmFbAA0hZs+E5dwq/QMLjwNOiVlxG9gq4/6
vVPSr7L3xsYfQfsTuPayBaHOEK2HegWGOBbFhHTfLfKB2LsyRMN8gaMjYb2JvHqQ
QTASp02z7lH/w4ig3dyykRga5jk7fpx/5U5PnCAesY7CkEFCTs1k9nOFnEBZbGNY
RmHZ/r2JQ7JOoC/mRRaSRXSbyU0QpRogZMwbGa0vMFoszN9wxz5A2xyGSZ4A8NWG
xqi3k9CpGV6PWjIUEsjsO0/7v/BLlIzI9KfDrwIDqPUXakXEyYreojghlQxU+kr+
4OML+jXKsLPC/Hk20DaXsvxM4fCwv92x2v3YvYzgbg6gC6w6x32L4vyQnGpM79/5
l9AQ6Ow3AoytnSQZJSe8wbkdjON5IAkoPPxPH2xr+UvMg/mu4GwZvCwXbrXz3xDk
QwVdM8fA0jfqCKS8wD//NiRPxy0E6FpJvKzaaL8802bs8HHu5ghqLIuJ4EM34TJ+
KfxusuS/EPmr/x9zCzHXF/upHbc42nFG7ZlB7Umgbbv8fwm52ss4FDybVp+kxnXw
Jz42WFi4V5d6ZVVf2xNzOKCQccBSsFTjW+vMmKhhmxl2o9vheExDa0r9eXX2B5R5
xfGgzPThdstguCPe5FKCetoGrv8HzCHlVW9Ws5sjDnAFiKLRTZ6TQmzQffQjzTTJ
HWtk03I5QgHsAc8M65QbzD8xYU5cS+nLwnfh1auGgmbghhDNE3wAjG+3vSxGvOaH
jbYxUp8SuSpn/V2/atvM2JsADBEMU4vX+t7VVtnVc1t657o8MyXX4rOQHHSvktz8
2woaJ1l2CHDoRrNqYjNyS1dwny1gG0Eg8unxH464YsXtl9TPP6VuAr4lZJhFL5PO
nVIF+X4/us/ue97n8rBATy4kM6KitcL1QyRDuGtV2y+V3uElgaejCqYgPsE57Orb
eT4GWsHwuBGP6bMULf/NzUnG6WmTa7hUo78TlVvtOAWB/CS6+YvtMkrV5RKSRuZu
iuqh2P0Q1vdzU9Kps3n4les1fHxYusQvzqFWva7JvvCGscKp0Qpm2Q/XBjV37c8X
fL4uBpsuIEmvPO2U8f9sUsH2Gj/gpxrDbKD4Y8N0CpIqn4OMtACnHWy8N/Y2k56g
G6gG+u6Mz+kdFIhxZAkQhZkcIRgv52TPYiD7HceBC5COs0xfRd/6lBU41Muhvsur
pIBt6zvMY4PAQRLl2Iw8DXmVmkupcvUQOUIOk9iqxtbf6LmqV5JPOPMkeX0/v9qq
H+YUk+iJxdmT/DgguN54oEifcXIMz9zRTHqNsbtmsXHbAZf+gBP2j6Fg0huVKltN
CbGNPbmYBvp79RnuYXtmYEsQi/icH0WhcWzdF7o3jQaU4uYwqlWLxPNHVL0f8SGB
hL79ByFaaQ68q3CKmBtlPxKcVKA62P9AOTYwOEow3iaNiYX/4PbRrNmXAQdM9230
VSVQhUnW3XpXLio2QZSuCDOrHR0+wALZeUrkOHMeGd8tQ6Aiew5mLVw2lCuTd9a2
/GizXoJNfpDmgVtRO21WuIiBJPmjYyC24NR+l67uuMZPWn3Xu9ReV8O+LZIMAjkU
e2tlfki+MVu9cVjspZANsA==
`protect END_PROTECTED
