`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Aw5g7S/UTtKiHr+tbqsObAlTk2sJC31wU6U+TmhgP9lup+6Std4Vmzt3UcHMCpM6
MgWGXU6T/2itBQ/Ah6iibpcZLVqvs/Z+0CBpKg18X3YjcYxgeQrXdHVhW2/5eifD
Q9CmB4S49BWW0xR9MWgAmbk2kMZ8sjMYbE7AfVLRipu8/Xtd+OX6cNfN+svd8Lmq
UGiKuTaEDJkjBdXglLuOLvGf/hsSr5+ae6NqwTfZQZKQ+j0I0ZqLC6lf8P1eL5vs
LhJd0RyqzyQY6uZWEY9EbFbgf6/tEXhRLJXRp5LcNOd4rS9go2gkcMfNZXS6GxEv
UTlcE4+nYznyjuQ5LLbvPc7W2KRDrDzLrrhOu7REjzsK9GNA0KW6meq2ojWFZhCk
59/QNeHAUvjM9Fh/gjypKQ==
`protect END_PROTECTED
