`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5rn4hhReI+2iRV2SrHkzyDVM7HR5Yw+P/cMdUC79aSREOCnkZQeVSu+dcNfso8H9
ONDiNCf2yeoCHu75wxuajGS5zB0QisgBHHQ5Dgr1u1UnKqplC05t6yDzMdp0rdEB
rWUPjTUQfnCDVbcz8zBAmGliiHFcreUego7hfE3+Zpj1tEXeGC78djx/L/23JlUb
uZjo5bo5XTgvpjS4TAe7iw8TQfzq4YkFc0MZn0K9SnKFsT/PpQYhAwok0Y2/WF3v
Hvrkh42ct8C1HgsW4b1GNHEYifq3OQZ+NB4zT/VjB/4vbxgBU3I/HOJNulg0NYqF
r3XGY5ofvlecuuZSF9HH8ikHpFQwRjX9vrZziLgXZ6SdTOsRhFsaSOqd0Ho8blbJ
eQRgED5kjt35RbbkkpxpuHwo7E9deVHCV5uee9tM+p6RF9LS9152e3P/4iCOHJj+
dvzA68PMk+a8I6nNiC6Pc61LQ5a1dZzrcMUA9uvbL7gM976i+Ok4jAiROwe7emF0
`protect END_PROTECTED
