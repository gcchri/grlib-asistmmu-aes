`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SR2sixaTu3EOvBFV/4X0ax5m5N/+88fGisvQIMCTZdDGIhVwF0F8KcrOQyUo6AJw
KJiEwZeiqud0mO+3+5XFWkNNbEARGplaO5w9nuRsuyRy/MqQc8xNkkIsVGbvm/va
lyK2NOFU1+QGRNwmQICLVXUJ2OqGFa47N7YZ+PkM0nZs33GpAUcGkt/hYUjtJSON
rQYJNiuckU38hNrfIrITvPAkNLgasF25iVwR1c6TApznDkxOlFm72kyYBx39hvVx
bYoZbg4YvnVXy4qxY9gvNKMN6BGpAXcxcHnKLn2o2Ne3B4mEq7ol0BwFVU/nW76U
1YbSkl7ZS+3tIZ9KAgm3sznCq6qsBCDq9/rjfpKHHacRiE0ZQ5mmbJDglOWDpixG
U27zSYBp3bC2uccviqN946TYSAu0fd3vjEwvxXqfSjDkI/wc5MCGey/2MzdDit5G
GkCU3+NXcbdQzMN6/bS2aXg+EMH2TpxWPhWBfIN3lzJX+vLpb9hg2Sg82nQny533
6h0W6xamWPPhm1kNk+3z0VPXctDAQfd+uKBbOFEI1s69tOWVGHjn/ZoH6xOpdFec
jGVIafIBG6xBeRk3X+HE3fAWgg7LdxU8Ri5E/+twxDM4uQxOjq+uIkbpqwDFAU7P
YM+2lnnFXceNRHHi3ee9n78rfy2FDq2JSIM2ziqc0GyoLcwLRSos4Z9jWg97bqaQ
`protect END_PROTECTED
