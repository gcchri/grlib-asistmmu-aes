`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v8Uk1/NRLCGZW9b4/bKqcdmTBmiQe6oBGbEiDy2k+oS7+tGus8WyErxNfZFNNBmK
cbTRC0w/Wf7gqjlmpw808cb3cAjmJIkj4pYyTs0AbeSkE4mZUd2WAcmORniunbyA
qWQSZiA0V4eAyWb36qpcEJP+flLqGzBTqoSczo+DezuZ0OteUssLxHy8UhaBe9UR
FHKLXa8yj9Z6bK08lQCWisK+I+hgwKMKWV0LN/YYvm77tEzREZDMo1jTCuQFbRGb
/APm7yrJ5IEKZF/sCRUXN5CUBGGjCOxeDN08xC4a8Sn0o3uVETEWzcOMaaLbV7Zp
2xyqv0LlXVL1958F72Rw9Pt3+UbEYDny1POr++X58a4ToiRoLSSPETeSWWf05B9D
BCfjlpTuUA2tXoZrZoMkOa7fPAI7oof/Qtmfu3pwBRVntOST1eoM73u0BcpzLu+6
01aEo7m9Mgi/QEiK8q3SafwbQeD7VoQBnvRx/FbCFkcxiNvz2YXtsLWvnRYdtQfn
i8wZsOKSRLHs1M422H0K53NAgvyVp1dmpU/Yn+qKf1cUeDJLtKMKQNe/QPfLli2z
Olz6iaEtjuMjpRfBzIf0zugkMvwiQn9iSQLto/fMhD4BuG1ClpgVtHAIisZzmaWW
e/rZw9eak/H+Pc6zwvb+KwYy27CR2Sap8KmGYyRYfZzZTg2lZqtfZl+oxQoeqsJK
ni67EJmM4X4NCM50Qr1u8kiD13lqypBIdg+Tn4ynbLdN+GWJA0BZpgwGIdNwc/27
26vzk4IG1E+1rGnNg+RgGw==
`protect END_PROTECTED
