`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hfky44N6goI97PIoUwdhq0GaLrEMrnJ0Emudi1MnpTZszbjrK+qcOsEjtFjCby5j
1Vdl+3tTiFh6IuymNMqjEL9QAumrQ3/W1PdCm5sg23waS3AbGfffXNl+srp2lJQk
koiyC6NDlOdjrMy5x3jIS8TwQdO0OIEBwrCMhunxJ/LHY8TCOU64NiiI3fRmJxz1
9EsEhbiWNqP7t579U9ciJ6N7TP5P3qKrUhLQt/tQBuQDDM6YOMZXVsm/YxvCmru9
XI2+Dz5VIsfsjMFxaXFmYPOYm8tHXeEbtM2jewgAQFORniiWAj7r3D/fxmJejQeh
nj/cQMu1etFlrUGBZSvwx5ep9IXzrHl2JmDTkGZFlPqg051qP4KHFciERoK0B0/6
h/j0Kx1LLC1i9dH93OG2wPm40HONHE59mtt1ca9r/pZyiychltm9uDJCWXTGXNUX
yH58HK6T1+8928l1+UZCY8+HNEEXBI6Q2wTBB2zLM34=
`protect END_PROTECTED
