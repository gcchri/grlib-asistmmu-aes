`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q5HJbH9f2eovJmNsuJbKValLznevbNhu8b4B6p6d3/pi5ODhEnx72jK1LBe/KEpg
ae0d3YorcozALSSyDGMdrHtKL+ITmjNdnGdpECcnJ8XQuFfgC9jSIBvc2dClHwy9
6gdVZS2xz/EfzrLcnKzhlexWlXiAohaRULb8E+F+5wok29cIkPBpUTAHuYngRYiA
cwI9r7jPyciVAi/TV9U2K/CTN2BqkgBeLtpYvEDcMWveKOKNzZXF/A/CDCBvSZQd
RphbZVma36ZPJ58x2oJmd0JNimgigNre3I/Q2yI4iiOBMg2ZxU3DAgZ20k0I2RMT
4tjfGvJtlTPtdIre4t1AplH2cDtgx7/PT6t49VhxrZvTrjigAZ6rrunOR2pOLWhS
2M7mLdAUjc5GU2Leho2aFnWxrJ4eeEBxvGrypM2//EpZOjinjpZKeZPfNeTtRz6z
amkr1b1i0Z2Jcuv6LW3mJSwhui4pIrpepMEjjjgslvCN8NMtqvpZs7I63+lfFtxv
4mPpf8+V5blPIPcYdCUWyVuIj8/QYazzwqpc5vcYvNmFhR0G4Ge6oxqu+Ywrd6iq
IE2cRQclBQ9mM0R1Pd3tGQ1E3L0qZNhAczktxkThJely1uVdJFzDhoaPpt8a8Xj7
PHu0H7Cr9FHuvdCqzIzTSWH+MV2Yeg/4sIu+gHsWlrcTs7SEbDGPi4Yct9CoUbfw
AVeXdOk/qtJXY3vGn5sdk/7SMjt9DgCfk6FWrIMxiZVAnK46HuDt4J2hvWMvYo9t
KbMRudkzieN1S0fd9dQbsbVDKFcg83Sh/I/7P2eUH3EgxjcHC2Evtwpzl+ayEAwB
EXk9hM0NcxhA8fZe/T6fEWAB0U2q3Xv5hVesIt4VURWimMBNB0fpn8i23B9JrRop
I5qxx0MrLNX6vFjIod2ElO9EIfrtcTzy7/ATYgsI/B2GlKRbVlrgvwxvecHdWBQL
7y7IHPuMpJJG9BT6JuJDhvPjJ0KUAiHS7aoM5qHtcoBzc7y4+WCeF1jbwWFN+PhM
FUWoM5E7q9ezii1Kpt6k896uAXEDuQIoelLyjBZjbpLicmvJUOCz8mMo6yrt5KnL
e1fKUIenCkTwx3dS1KDR7FUV/070mwGfIvtXtMqFDsAhApLKmI6xCY2hgPY/5lmb
nEPsyqs1+4zIMknImpF028aHtkoRKEZPc8n33PQCGM0U2D/PkPC2+7qKzwaAKGw6
7gWzN3aBUU9Vk1m39JxYuCgIw4pGRUJ2u+sxwnip0dHEmLNSrTmQ/Jdzwrp9WSSr
iYM/tXoKtQ6CZJuCHyySTRHxlo5pummb4weZGhT1Mf5F0YshCPvI2QFL9RW1L5Wc
1ZapDBEFtAIK4/dLtWGTxGiRAk7vWgdeSfzOghqK7dHGuFc+H6VZ4Px+X20Deyzp
sgzbUUC6lHCm1QL697YfROG4v2YTbWGGL1Ay5fBoGDKZDx9aJmFOy3hCbhyT1JRp
lJfpaN4kNC1gEEsIr5UY/tNGV/QtRl0ZHJVGMHTml3j3pS36Km+g2S5QgDJkZWV5
j+XMER8mdZac1DZEQnSW2FaQPwkaRIt0qkQFJhOKcHnjBlY2e4u2iVm1ehXKo7VV
Ky7TbhVi42mjoeuhTp/HwB/B/jdijOUjBitDk8v4j+SKcfDXtkhLm0TytMtQZns/
0IEgXopSPL6CqO/016MYflneQeWQeWnK5nDmHTF37cy0VAQvro+WUCC+8UUUMvo5
sgpTmA64v3Z41d1H6sEuuy9xzirq4fp4FUicwQuiaJoO/4/zXSVA2a+u8W/S9fO4
DV2u8GA3uXWRgAbkGainuKlTvxc78Rj3WsnuJEOXj4xWa9HOpIP01S2I8GH5NU8o
hotO6P8bnqwz5sDDvJ6NK1p+YGJetOoWVKZLYnJAcdwrNVZLOBvHDOS0Lc9ZIqec
omvu+VLHxkVPUo3QsWotRgJwgIwbaLnellhmPUbZosXlBNFA1DlBDi6Y6PCrD7OP
rJBZY+2UExm/YhySRmF/kinz3hR/ScOizoPUqaZgxvGNIYHYNXXTi/g7zHN7Df2v
Wpu6lpZWVMA2QiL1yBvCV3P23Bt63bqjQU1l9txHX3XxDf/n8nkA1GHzQS/IfiL4
f+VU1SEzjnj2alvFDdL4dODlp0nnYzL0CMIT8pM5xIlYPBTgg4yaovuwimg1FbIp
H4ZyXV5yi+Fvej4fzqxzAbb4IgQzfwVi1NyNATqIycM/P9aT/AJ36+gCFdWrx/aj
aqPlXACvPRg/vjQc4SWxH5Dw3iUcMHgUbv57PQzNMCr/9LoRXMxz1s0hItIA7qyu
g1V176gchKsU2H0Tk7QWKLcpw+U+hGl1SsbMempmosgilZdv3so+lnp6pEKrUlCc
blFpyYWVrsnMjWF0+FeORlHjpaJLEn/gZMGX1Yzt2lQoZ39zdhB8g9peLQsrcuqu
zGYgJCVIvu7NSrECwwXNGqbpdPkhFPamH6kZNzpwWfIQaV1LRvjFAIj7heIjQ2RT
Seh4xejbsyXEgEyxCYyRFVpTtog8cOj2IP81WAaK7/YsK85e5QKdQVUX44NFPO+Q
4/TxxTbXjJzlUbtdzTifr7tQMQyLT0JWq6NUjTH5mPSoEUYXvsq7JsbRof008elj
5jtPKpghJPhxMQPNNbZdQTrVLEDmBHPRQNwfil9BnLH09ACw5aqMoO4r1WzcR+K4
CaYieDx4FLFwh77VAjcfjId3FD2ZOrisjD6lnxl7XtJyzBP0ym4dKOZx0h6MEbar
6JhPg34I8/JBZdKJpRI9SawqEzeoHR2WKfdL7T4RtBBSF/czclqqtfZKW6OrKwgC
qJeK4P5W9QK8aPfHH7ldoyGSrXMfSx0T/N3qVqJDSqcvS1DqUwrE9kn4fFUl+kkv
SWdXpWr+7mYZSy8z9CqD8O0WySGTrie+Jn3fuvqodNXv4+gcY6x4Pe4Fdec30A0B
gV33wUJwhPeqOHegFaFV78SSMIihYVcXxLKf+bJKULZM3p1CrZFvDj6tmtmpM1+w
hUtBruIGNGy4tKPpmQ5V7TXyIj7GGEZIETZmVuls06Twi/7CM2rY8lEBilev99At
lC9M+L40WoCkcxA/ZT452hdkxwdQ/hJvNCIOltoGQQabKlJJGOI7hCGSAYJTolVA
tGoT2Mc82UW1sD8atjnV2aW1dJi+QrMF4YcVLcDSirBX2iMFeJpdmQRw2T0FNSwU
tWAff/AUPWcXF1FzFle7kwZtZpRq9Ln4JGsFbMiyAliAWSxH95OrXqDTlk57OFF9
rjW38kN1kDZiaZ4WVT0IuG0Qmk1V36HgMQOakMpW8SBH4jz/0RIYEhjKHPoN5lup
nGT55tgXv4+WwAxLEb3vrCMceD3ibCYY1Kt4LrzSbYtEhWEx/6fQzMffHLKQCQJV
DJxUctzHtYxBwITXQu8PFYP0d77IwOb2bdU4HjsKOoDDd5RR4XvrxXTMyLlVVZ1P
AvdqqsWvguY2SThD+S8ouOr10beJgT4fFJBZlbQr9RJKhVjlLIHTjKQKJiBd+PHQ
2zs8C42LHIcwSdtYU5LLbl5Vv8vzSE4VMiStZFtnc3RoHINY5U6KplAON5oNcvVy
yiIH4kmH5AvT/Zf5DXQPjs9hhJ9D+uqZjARiQyY9Qula9rIlJUpes28pXXUQL8hS
PnJvDTpYIiuU8mxt0NhdZRuYD56Y4kzD/6jWzVcU1ZGYfa7b88HVcz/W+EZwmS6E
ky+gGKA1QHStceXPyNUUlee1AGX9xgCAIFdw63x5q37lHx/0kIh3loezFsYTj8oV
iLRAwzum8onUirN1tF58jSnSi5AAc3P8HEp169pohhmxkI5h4+yeWjlp5M8A/P4g
O9FUshPnYwTvbcKRjVeDsw01yaw8Lb5GKxgOfT2uk7YM81om6A4slSXDfCP7Ynwx
2scbw9/HJx5DGIx+Phz5dvEYRMoLNMYXgWwQm1YiCcaLrX7JndkH7I+9pwhI5jDM
fdoaSmJwFCcxEQDGqBP47p5XU+3YV4XKsVwBOTWQ1W+VxLaJXwYadVmLTVLgKeu9
h72AWts0p95ajvcl0faSdzA1tz+B1bsbShH7ppla116nna6mhTaEb0/YI/j4At9r
cfUcfpbqSNTtpfERzUDFJgkuHQpkErCUXVEaj5i4s5jM6DkTC67+/ko0OR76GxCu
MwvQy5fFFWLNBU5wqEHksma6ErBEFg0lBqQ24m3R4AucSfYl1p1LHe76JsRLn+Ye
HmCIyoPAZZVQIYdx29a9Z+TbdY33S0SkGY8cqq2WLzWQbX/+sXIlAgKSex4ffqm9
bsRaVEHH0zz9E+J/BcRQj9opg34ErTqJbtq7IitsZWfoAj7928ipIIA0uyObNR78
t+pPs72yTkFGBE9GbiwqkpfRkc8ASzCSRX9BoIeQGCDM5XM4GdTVBHU5v7xSuhwM
jBN1Yxxxk9Qa+NC/hlaGQuspSuo8vxhTexVC8EHx6mcKUfAtEtFncA4Ku8MxehN9
vx8ZiXbPiTm3+OSCyP18RypWdItrVLeHZyEKjR1Ui5PPTZnXCwulTmjCzevIqT+f
Dz7XKTPj05gul4AfuvgJi/UL9LzxsFGxRCYWHa5UIY51XjxQS1FRUstbbTe9kNnx
i7Cjl2nxUbtrTZFBLWhXHAA1u1njtKquzGKOskEIogc1BPALIVCJg2EpKzfxZ8kV
pIvJMfyIZ/hesBB9HA5DgnW4g6psszbI2Na2Aihc5P4vhP/u8R1a6vhnT3qjM24O
awW+5ZgahVuQcdMM/Z6HTCnFyEnt77o0XNnYOmdGnjwWG2fQEqlAIQy2GNoJIjQc
GOOQXhec3G2PRp0LO9ywJe3KP7X7ZSf0Kr1NfbpfyVfcMTXgjrszSAFtWoXM5VCK
IhRRi9nWbN9sclHv42ord8vXRW5itjwzDJhXi5VUzCVNpXTPY+Hm04j0F1abm5Bg
PIcoP/TuzkQUK7+aBNBeWfR7QIV3zpmEnG3u/Ks57gs6pwUWJ7ujErFkEA4P/VL5
lr0DLeFcNGoEDNXLqUOoumyaNZqh/sCcVwlPBiZAphws1wEXcGXay1zmGBO8vB3/
XM/Pu/je1kkG8mLPb7ybSOh3g2zbN7xZ8Zec+B6yzp5ykYckpA5ptQBTtlv6d6O4
3ljWdNnGQb6DVPYXk1HoQv3dqDfTeocSYLmQOOxCR+oxuSxl3BDI4Jx9h3cH5Hej
Keutn8CiFkun0td4vwpBslPEMZGqky6Qz2EQ2noR7GjNEApBXGbCfyVFHugu+ogt
iQnhrmKMmHrerKjU8TWi7m7y2XROF6A59kuLk/6CuuPMuxvwFUSeqmmppLedh5S9
RGia8bn3bLSLEBS/LN08TWvfsEU0Yrlbzte5hC4ywMmXFLj4UtQArlKHrmKHxim3
UW9WuSfXXJfQHfWNG9YvSwesANI07mGOflNCx9oqgsyr199T0cU9Fu3ZsO5PlSz3
kHKkMLfhHu6/jp1/ADS/ooqRL/O/ibJfWkQg6o8QEJuEmOYBZAg9nQCnxWesn/hr
/BD/ldh3Xd3xeXUF59S3mvg7noHJjbTu4Ol2tbGCpkLdXOKc7rBBrA7dCmDgVGaj
EqIoJKCI6QlVjouanKenNrBqI5C7OSzmLOlJRVyyo3KF/Ukt0M7KsTiegWojBwMa
egEFkEaV4T4VIqzF/ognAwvmzek7fW4pA3q915ZkYiVKjjqrqsEO+vj6M/YJE2sf
c8F0TxVgFUPNpBgYMbcYtpJNHbdTwbyCdd8AAGu2biSFyhzP8SIByQs26/+SrkoT
j/GECS1WMW9MMzogqjtqeEiSII1OWKYewSAa2K95CJEHF00ZyB41q98DeCmpJIGO
xEK17ikCDVG0ffusZqRKF32pEmZjkch5uDCE0qEditsKFibbQTLOOS2yh0vMBBB1
srDQZrxn0gdhMx3gNfWNKBiQbZXyWKL+X65feONtKtqrGWYFbwwH7x6WJQccv8w4
JZ5lOW9U7YF8xiffl+Aze2NBQe9jriH3ATkKs6hcXRmUJEpQQo+acPDTmJsaDkZq
kZP6pW8ExFlsCMM1qqFKClsnKXu7poNRoWDhSms+oZENq4jhBrslDjc0fN5vwUdG
UQssnGq9+yAhzNMezdhb5GMX6g+8HkxEc2t6itz+FfDz6lcFBxHoYhm8u3Fy7sxe
xB0X9qtpHe9U+ZiPHUZoS3zOXvm62M8DbWEsjtgqzn1jf4UCrYZEQ3jgNgEqyWCH
8c2RHOeRPnlNIdjfDBJOFjlw2qzgNDNyJXr5GfKixB11pk6cop3UBjUo908thEUq
Kd6I05F3rEKI6pePfpYLqHRz6qtlkFn3Ka8D2ablYR6GyB7qn2yffOjX8rgmX4bv
K8d+vXYQhgu3Cd4U9erxxwNUxYr6rnzTfa25xHAminVaC8xoMXqYOq2/JnH3+vf2
/O6aR+EMbykgHZ7HwuKq+89eearynwcI3sqY6hy9umYrp7h9T9T815jXfr3XfSvs
UH1ELFk4oRBesunMMiLt07WFcKcKZX7IAtGDLchhrENmACvXFjoXqKRoaQrXEx/x
QzaOwbxEUxvN4IYyQTumpOdDHNJ0Wq5HC3Cs4O5tILnboEhpASnD++tn832RNbbz
hMchK47aGPHMJ+KnwVQoRfSBuC+HwOgcBQ0vi/KTnhczStx9htzNU/3ZYks92mEN
pNpeEjTX28QZBRaF6NvqzqLTnWU0abbtNPxIwJk112ObnV3epqee2+dwzjj/1XqX
BvZrS126mmHOQbzbvXhgkIvfgIePNi9t6LGEkQpYlsS/3B9JiNieuK92u1lFiMq1
DZPlCiNr3VQtcmaffE6B2RdmLo98/JtMaxUqNk9Ti3zb0EK8Qh3W/v5/51lci1HX
EFk5pmEPrDC5+2QKe+3h/VFjf2gLlgcJu2WrLoteGdoM2kk/URfqtCdPrCWQV9xm
XYVvQMjUV/f31T3+vqRovKRAVp2DXz5pXxW9p+np8PTf9WOxD8USbGaHfNr4H/76
zHsZwIzz+oXWRw+BNRHY/ksNXsk0syYV/StTa7Giqj7WKhMlLyRoNsobSjMGaMxU
7yzQkQPbHY9LBT8KDUbzgSny4qJ7aAqHxv8X21IAZ6hi/OFgNRwBfzueCXQTWwID
9m43aWG+khiV/sTIoW0nB4Ach+J0mfLBK5TbbiILrtDR4GA9Hh1iu7PG5j5/X8ds
sbdl+Cmu4BRlIHdGV5Dw13zKQNFLQKqfMgCKlzYcoqLxmFrvI1jsOfynEuC6pC3q
ivuR1CkhxPjd5ot8CDJKMGgwElSnybip5ajpQwVZ9qFiSqAln81743dHaaQqNbMf
/sBa5p+N6hB0Fwi7Guac/puQeH1QP5BOS9H+JhK2SFhKUfIK7e1t+ypq4jp1mqq4
crfHT6rC7uhK4yXVOIrSu7ruJHvOnbY8kAV3VTuYGDJAuBNdSakWWTu0pGmuO2WB
78PaoyQs6y5hWkGMhxHdsyAbBDjLrH60E7YUQ58JdrExZoDHggseAnZecPdqc60n
/Ej6o4LMJy9Fi9Zn/dNzkIPIBUPADBTeLJafZZZBF2/wVK7MGLcsrAjBuIsG6+tt
5aez0rwzptPn1UqzL80UZItM28Hk8m45H3rBd/of+/iwnQBPRSvBXyVs7SOcjqrE
ygM101xKw5Ozu3MAyUVvu1EV4WsaomTszEUkvQyfVXCc/cwzYCqK/jYPcArAjwUL
MSsgmhmT8SdkW4H86NxwJhr3MFNRSMMQJSrOu2pGo4wliIqxgdKpZOPuE/qY0QeQ
agkU8thZawaNJBDb1gzOqzx0eLchNfp6K5hHk+3FkjB7aUoJ4wTZ/CUMjB1dvwGW
5JfqFFwQiJZ8kOR7Im1zDPbxKBIlCKutLCi1O9h0rjlC8rSrVbAYW3Wpv0gWFHdw
YiM+PQoptailhWW9Dfq67pGU6hMCEM1R65mLCHiM+Wpbw3kSeSFWt4asFwnmTWuc
UBKLRrZSYCm40eba+Owyj2KO2w8FDA7ArR38VxxtYZGLXROlCo7WvrubWSlmZajS
iDnkMdc7d9XO8GcRdniT7qw2V6hQaf38xjKOx8i1PjmWGUSQwSmRR/xJqZqhx4l1
2MQq/5YEPZrcKBF2CFDJPzAKXV59cVy50hAvRKnU0wuXwVFsRgQLciNdxqlFktXj
yoIZ0pddvavFwKcEX6rJf/a8Uy9rqaK6yLo0SajlubQZlNR2syv9TGx4jlfhTzhk
5ztHR/JnQHUsspAeU/U6sfavLBf//fGSBJVVlDHFzruuxSw1PNydQgDHJaWD9p9N
Awy0bDkn4HAZ9ccEBl1VzyBsT8C5CZOznrmrdcaKOs3HWBpD5fpkUiR2C8sGcEFD
uow9EqbwfaKsnHXNUzdbuBXqAeeL6EY7mbVBdLcU+u4tRIeBUy7E7I3vK9Y218V1
RroMD1G0yBWMPScFB43OUpZRhWwWMrXba9WhAsVQBmq8uP9VEUckFJzwFchbAKgq
If3KZYm4h7FtEpvvM460YwEF5hVGOyy47VGPcsh6lNV3X6wK3lr89iTxBnTWUZlF
p8EDaGt6hzjaFMAygEAgy7M9uUQQH7FK7DMvGCZmSFmPCfsyeit/9hPv6LiVvGsm
WZTJJ0u/3gVYyTGN4vPfgFcXgyU2lla+uygzEDdiBug1vkgvPVx3lUg/4hPIiVIm
Uwk8QwuSRmUYAepn7h/CSCN0le0wtPbAQfKpEQUTpTCUR0UlIMfbAxaeM71m+O1Q
XpDWgEy8aR8eQ3fECLjVhgNgo46+Up4bMxY1VVW/LeBIRTyL653LIWBpSq5q1QNX
HxgZgSL0ozW/h08KzRxgLgjFU94HHshJLGo7s8lAAHLF9JhmhwE90E69kBt1hHPM
ZOgJkUhiFrgmgq80105jnOhttAwou06N61YXnWocN0UHRrdeiPIpopm/GH0XSkRz
HqpBveR600tUfWTNDRIdpA3/IuiDXTLyRdoJIXs816/saGbhF3O6ErnvdoepyYy+
jg9/G7/MQjbq5/L/FVuClrGxZFpQlmG6NglFpOXlx/XovftxF4tClrSuPxUrr+ou
DmQlceVFpORD4FY3iRufhvBmwqekwTn+lMxuxL1QKvsg3xVwkfBnaXESzFII6JmQ
5EzLSf6eym8IhibSyaWeDYZMdffteDWXyI/01JfmxIIu6d389j0Xwp1bmvamj8z/
fOvwqEjLVjNQ93SdxfH/DJEhYlTMfuqCEXxhWN63KEBRsERdMfpG4m25SUGaEapz
nh1MApj+nEGCc87w3eTfK5CrhJPBI0FFXKzdsDHyDOIeKsrE4qPU91UcSYw6HekI
Mk2AesWBvuzY+PrzuijDSD1olRKwC8OoIWfeAYuw/oDgd3EdCNqwdHiBJALLGR8M
b8qWYEjkfX82ajrgfwmoP1z8ilR+PkKGvPNj+8lYTfX0na8ZXzJqksaYsrJwQUNN
1kK9D6l0LM30zUMtOaLiLZ5vF7bndIlgqMgyo4mt/CxEgS9kcT+vndRVvOlJjYFC
/cgcJg/4BaSCvFkd/dYaMw2L5rNZh5igl/2qG2oOqH/6wUSxwdU5ed7+f0VYbJBm
TRUnfprkJe8rbsJBqIBwCobZmSvDRYvynCN8TbUW2KC1J1FzVpEjAjQRPPrQ0yy+
chqZ2lJkPDnFCaTUk3hoUaa6u0wVSgKaf6u3XMGNmju9DrpZjX+7eBRIPn4wvqax
VYXeT+dptr8r4cKFYHEQtRsS8VcS/CbaXHuQ7meQPJDcMCbQCVjNBOGjpQfrFJT3
l0qwIRihX1BxoweM6P2PHEhvZZlLclCnn0015O/wcwuJybbi89KP0EenxIB4cYyC
xicOPoQC3FFvrukRhE4aI8Hi0g249qn9CBduNq2v3Jx04yexMsGTmn6DBjNCQWLi
4c8tH0mORO0cSK5v9ukFJu7Syr7hFm3/n+vn7n7uI+xnAGGXvE/zWYXqGNu5tRag
ZETSOFu+hUmdVcxYkIql/2T7Lz1afucuvlxDV2ri2V7I1D8ip7BMk0Sh/8H9gcqf
i27nOrpBsttE4u8dJpxSatuf4DK0o4gPv07PIeSpArSRCYv867s0E3ZjMLkMSF+/
SQYPndJn0jZ8A5uJgtQveas9rStTb188o+FWBZr1nD42Ld9r+A34E87N6iga2wHX
5xblh1SdWaSq3x6KsOFqMA==
`protect END_PROTECTED
