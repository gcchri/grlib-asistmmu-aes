`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c5jMWz2snIjmmecZlIzEOSPIimzwd6obQzy+LZxY9IGa65uW1+9pzJ9VOqvawO/s
/JkAkGwntuHG378qYLsT6ba8WvVaJo8pASXJQsMmyjlY/RZ1zIIx97+q8D6j7mgM
nZ81znOEikS7MiX8FCAt0/1bDykHOTdl6rDHCTlEGdY17ZYM9quuzfbU9aHxopXc
hbFsT186fSzuJDO+HLggdxGjCFeHA5lUTZaqTe1lP+UqkgTti+CPfMWu7hR1w5pI
1zzy4NTo1VIJ74ahtQ3BH3+OOcqO2x9/X8P+DPajk5+T+sOU5Hd5SgE4ca4FC6yA
V81tqG6rtzcsWPfXTOlTXA==
`protect END_PROTECTED
