`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RLVf9N8aGGHlIff7BAm5Eih2E1XQTfvuhJ9aYH6U1WAlRRR2GFEjzqu8JT0K0XVU
eyEbD5bNVhmgqYzpt644RIAsdzFay8k6MyC5krM5wwYTofNIx2sD3fQ0cKZZoVEZ
jSdoZhx19Kjaq4E+q3JmJfx+RDZo5juEEXT4Ld0pIPcy34Nf6zPssM4iu7pav2Wu
6FB4Kyt5J1f9LQK9rxawEGmC3UE0NwUpfEO+EyjGEsSRCtGtaSSUHnsEbMTN9mWL
XDi0/WN78GO9O4CzN9YpexnJyB2FJzcUA+QepgpoDOdB653xGhGHMW8BZiyxwB9b
XcaC7WhHcv54huRGS57mcVzvvTYhkrZiV4pW/XtF95PhpDeMz1iSvppg0hEHDRe8
d2YARWx3K/rioBJcjvr7ATzGemE2ggmvr568pBDH33kXaB9olcxCSMQGYGxAd78P
Sg1PIn7kFUFc0EQ3S8FWUjJA37ozcww5xPsOrWgMf7HRP4Yu6kfpEEglrLF/A+UR
o8eRXxTe9hT4FZyNaSQIyfTkI1qygknAJiaLWW25VyY=
`protect END_PROTECTED
