`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j+NZ6elSVJF99sCscNSWlO+QDjSjUT9ENTD3bCxpXygMc4gmZBaINjVqTZ1Vlqgp
MQk/ZAzjB8N0GF1/AaRYraI7PY4WWGlqR61WP6q9io1VwKzf577ez7l1DxY8ib4P
JjSmrsn41fXxxppfrqJbwVy4y1lsAxsUAnfRFLeA0rl/VelhBZVUlJXgHgY9YCdU
hKE08iU7h0nsXrA8cTQFHYEPoFrnMNK9ExDDW5JtK2WmWgO3G2lcE9+zMCzlKd18
ertntPM5iUTbIACA5Eo02QtLeQUC+f7jKeD/DGeh1pMGkg0c5QRDmRn4A333iHEB
c3xuCRcNaxF7ROznJZ8QCAB1VIFlEghnLuG0Fqcx4am05f2SerkVXuc+z2W7ulKA
x3LhK5Z4OQA0S96R7tXkVPGETjFCC17dU7N+eW/VSs0jEwjHpBEPvsI4SrAKV91f
NpVnJ8tvdBvErhAwDmSxK4et68ILieiY0zlqPgRL0dpcmLVCAnRNfs/FFu09++Lq
oV9NAvtIqL6yFhGBLg51SQNTHoIv46PjElcCMhSzRKTsftMkdinzhuRavfBt1ChM
DfBG5m+QSCz1eQRtJm2GH6fNUtuJLA4kLOkEF67ZrK7Wlkdjsu4vdbciESG7OWhi
aw2ztLloLFfH1hIG/FKcFXzJ3RN9zYun7Di3t746vrGhYNvxsYMTyjzPX5xJOG96
f0m+zWrPLPS3iPi5cUjVlZ1fJcZgiBkvzUY4LDAeevWuxUNzGU4cjpWWCYMkuMK+
C0kMaYTh6t0NXJhb2kjyjcILt+PaUBn9cR4duNmmtLpmCmMgurCseibLCc+Ban+e
bsgxG5+c+ixeQsGk2x6VRkqKd1C60u3n8RgD7QwpOZLoLZDr/KEPk9ziLbBx1AkO
8AfqUwZqgnqUQ8R4DYYTEIiSNBI8hxuqNo9hKSgqlSJXHlLHtZS8oLPalj3fS2Mo
SNONS3PdMAMd4Qlgxa3tzZSHCf0AZi7vGurK9G+4jR66xiDMeg2p4JvU8E+KfYMj
716+AzMawNp5Zmx7K5D7xpd8pBr1rwJ3hSo4Q3KmRPucZ4rvnWu8MJTYrCnRw0iy
LFt04BOBTG7JGtqUePfhNMSES04pA22r61jfwHVG+ihvZP70mLwy0FUGAkuj+8iI
J/oyjFCLOJ/sKotaXSyXmambgLpjUUwlknOVL7NCGcYx4PIDAfSoZnLWcAX/Gk0v
rMN7XfWcqSooupBdPrb5O+S6Li5H9XIM0ecWAEz6v++lyMXeCbCc0cKRixmx4YxE
cAOjPP5162pzqdmxqFuihHMDzHTK49o1d1HjPBKiqDHudrKS+5N4clqahbdPRKF9
Np0hZ01XXhaW6ZQuOlLEW3dlq5E4nDLU9ktI6VvOuzfKePct848HxZ+rmLRXN1NQ
Sx19EsNKx0Z5OXlfUQA6GkKTpb+aaZpSF+hPWlP+C+YKpX3npUVg8WzmTZBzdHBT
FhW+IPE56Th3j8yz6cO6gUavu3JsFX96IPvuMZjPr+KTV+IacUyonA/BSMAyzi55
N/igG3jcrJQ/LaUrSGvC1WYrIbxgw8acWNxB6cK+6gDWOJMuItBdXo7Jf65yIq26
5Eo5UuY8SffQdy1OSa3wSdiEWP9ZV/0StmzbA3Yg4b4CKg8/9XVPoovMayvyXyDf
V582pb9Cl977amr4Ol/w6yXaVPltLHo4sEpCcbCgqjAFCTRx3B+0VjhLQVt50Ijy
+N5iMWoZxWpEnPMNc86ah+pGW/tRGXjXyFbnMAg/YdVV24qd4b38FSMdzk/XVZUc
2DsxP0qdrfk4EI5iKx4AfojVgBXLVBibBQURVMCiUqPvz1d1RmQcKmdXS5SHpFwM
/ukLNUg7TadgjaHS3CMy1t/E1s07pRM2GrLWkJ+TyPamgMFrQ0ckcaN9GSCEaEC5
cx4+k8KTBX4w1+Lh+s0Mxak8StYU7i7xfZXpGcGrABumfkapXCJ8yvjI1xnRIYWK
Cp0J40hUYOzOHr/Ll9BLChDWp0HaSU+QhUJT5TAQaBugm0VDZCk9fka7qBfiIQiC
PGaoFVuR9YmDYoBiGEl2jAP3FZ+lKPqON75XRHIV6Wzi5W3lndQRuVZjMhXScl7H
REtYxVtEnzHyR6wcibmCWJ6VLj+QCnyIQ5zlvJFONKk=
`protect END_PROTECTED
