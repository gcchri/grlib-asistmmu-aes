`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+2cCCud+04aJUM6iDggnK6JqFVCL3M5Cm5nn0mGVcyH9qVhTyj7multglj+QpvJ4
ZakIyy4mLsSW4amiB2EAbaPVUr7ApdenB6njgsMu2VHnyRzQDfAqocg12c3Ss3im
f4k/wU/IFPARPZxsA+9Mjm9ZyxaWtwZifPxjD6LStSgt8Do0xn7X4omSCb2c7PBZ
QvPkwgOk/HRw1JqxVGFpLW8dSeFreHpvFG7nY/iayaG+MwWWLrnNGIy7KHLLdUcP
IqpSRXaVZybRDY5SYL+Lcs8jiLkFdVOvKbJMsMo63KjjJsJaE53UOXYsb4h0YiY8
GbjMxUTliKFs5PnXC5Ch73Ktb5g6YqlcAgKH6vLtfLfDfPvz9pD7djCn4EYEoU63
x7apt1VPSofQQ50t4IkJ8g==
`protect END_PROTECTED
