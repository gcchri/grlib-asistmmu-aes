`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i5ZuR3fp/i9I7RQvyux8pycRagdnp/NbqqS1fezQl/QpPNzITya68KfkYi/2qsdh
iNDpS4S2pGGXXWBvEmRqHNO0wQFWdkFX+TwvX9J3x0u70Ro96ktWfqOeioJO0Uda
NrfiZl1szHvOopYeTe7UjWAGWECORVkciCC75mq8+GFbnVfWYuf3hyvc3g+XHxxx
A4qg0I5p8yr8Znf/kI36PPyf01Yka89i3U6ddDIeY9wPAaPrFIT9DAAdvvzWfXtV
jqx4jB5kJgVkJYWh7zS2OG1BvzGd+OKt+1T1a6H4p7/f3aF32s/zOJG5iR2zTAbM
BsmXFVHXJh9SnlmOl1pIE08JGycJmfi/RypG+fCB7dbXLZr99B2tw0wkKkY29lOk
9bJ2qjubdCTn9/ql2ZDvxjsxvreNxUbHrB2mPbGdFjVF1Lql78uu/dZe0yGSVnAh
Np3/NGGdh7wjgUmamQ1aHw==
`protect END_PROTECTED
