`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Devh+XjyWFxD/lVqzh8MV4mA4Nz8t68lsJ7/dtkld/IxCIYiqE/tOY901UpjdEfR
V9cCcrsNFWm7innE3xbX7dIE7SN/65XitForA6+bPP+VQAw4RhihU9D1wGsUSLLB
XysScrTgwYej83zjBTWYkl1puHB6uPZS3xvxIzl6FiGUFoiO3IQNOe8pa1B8gWZy
GgklEv3e5vhyokxKDs22Sc1PdML5KEr1D4uXMyOCTDhMtSoytDlB29dXVto79UNz
6N5uqI7Z0/sVaNf/lQ3TliTprkLUbeIxQxi8eKtDveNOHPuZwaEA0JzS7BoklcQD
7jJdk06lKB3MFiSw8RCIQ67k+hBgzUegIMhCKjuyOj8U6xJMbEBkf4ao/Qtod9zF
Pfg2xKjQdAm2BQQmmJsHetNHBXffjwz6B1pxyVVWaiztXdXhhz0tFDi8RvOZgCXl
vBoLTM3PUXHeAhJfUsSKuuCspBzTyhbxwuLBFv55Ov0UJCARgtHLwLl2D6p9/zYW
oTOdRF6LZAsUwLQ3ChvYoFMWXA+S7FXCeFwi/AmFmOFYEns94pdZJBA0ZFvGQGRe
23JQ3VuLH33Xdq4m5G7oP+lLrTTUg0i3gNjCvnlp1jWI4L1h2icYWTFYgHsXi1l6
1wJ2VSw3OB6Ga96zlM6KwOsPGHeltGkpXtUupGbu5vMEbjGr7B/9UFkgYCWl8H08
XBu1zRIhKBirci1OuBqOL68ZkLhVIq7SwYyg9kEki0pahP0yLD8TfVGvO/X/KVfW
AeFrVwoOSBsNkLgD25724R/dVQdk6FXCTbpTCBKEnTEPBwSl3+sTyKGGM5uIKGc+
BlX0gAKjf5iPxkupAayLnbNMujIgyOhHzPzwMYbOnSHSnUXmzqtlxOiakZi8BVij
DZ4F+NhfACwxA6AzyOGYlAoJMblqyDyGDlokIFxjK35U0WZTj1cdc3S+ZeL6RE4T
crYK0OEtdiMNQES8zDGBS9uYKTVvtS3iHt1VUMe7gME=
`protect END_PROTECTED
