`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s7xhwrDaCP3pbro05uD8OTumk6vp5aZP/HeWgIcNEyasdz7ieTNQubYHEZAiqWLK
+kZrZwGgq0yOWbNGVCRx1XxqCnpexGTUmyFzXyiRJxxKfa5tZkbTT5+1T3d/ia5s
2iSlCCY03yINpsZCPHgGSLtAggM/ZqEMOi1Fk8c4vafi80bxWpo8EQ1HSg1Wro2b
/AAIqNTAHNxs74pDz0CCVVJ34YhF7inlyk1KQ5BfrPObsHaU3XNi5QoU0yQAh8Ve
r2cZCUKHbtqXhAlFZ7SNH/HIleyky5auXmtdwadQROgJSk7yCvXWzTf91cLQn2hH
YvUdwKti0xoKCQmd3f2YUDOWRHjkquGPbQAN5EdpmFxFJbFLxF3xiktLzeTkALAr
YUqOk6zOVis5O4YLPZIS/fVc7GMbNPNPoyPkgnheAOKrzolRXgw4HjvFTd/VOZl1
NWvUpVfYtkwNHHyU7P6/UQcB90igY0tfO4vBjCUobXrshq1kGArK9dJOFUUDnfLr
8/lSOtiVVELOUFyXgwNDmbnCoGv+PST3fRX+IXOBJBbJuRp1J7uLBc2rU6LwwN0W
hNBWNbh1V9fuE4frAZAuNEa473riDAvJ4IphIHVEt3ScaBppEOzMFBsTLs6c3eGn
U+5IyJ7gqOHw7eSKN65ArxdtPDwUUtCpTKlbyHEKNRDU1RoMLTOonTwzY/X9H6or
0IlNZVjwMtbr1RWBp/qxebRXeq8zysCPMMfFoo3pAztg5YfQvwRflREVI0Hn51MK
GYhmzVSUxgkVZu5xI2voHxzGInk1xtB8pWPRZ4eSZ8xEJtFJvUlQh7C66PfSh5cK
CGZRNTm/OwfB7UiPu56GuEJaf2yXVY5v5DR0+/x87Zo2GTZfh0LZFYjq5sh16cyJ
v7AmlOyfjVFXp4Mco71XdQ==
`protect END_PROTECTED
