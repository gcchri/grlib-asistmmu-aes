`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CSFfEbt1NlC5IfDeSvXvFSXV1hsPvW+fTzD1bBunMfElhP/rYPICbrEwC7SlkZQ1
Bc4mG0OipQiItoPy76JtynLFNOsIxA67xoTvSbUwuRqUUBiWlFT9s5o4pNLOoUTS
zPGvQb362wgTtqtBY711X2/dbjE57PBGrBwHNnYb9chAbedzwT+APiSo84UODDil
T3XAPPHmRRye+Eye1dLKowE21DzRfka/ECq0IVapjl7YOvvtFDwkYq3Mw1hEcIbz
ZuXrlloJx3xgYgM9qqATZWNneWT3dvlCOhMW5vQwlNg+BB7cL3/dAFX+AJFI5q9m
yOkox/9Hm21ne42geFdhsmVZkDrU4ZHQO62VDypTE5uxN55jP9WrXuMnET0+HMf2
1ISbAzOmiSP8X3810LsnNcs9Wdo+5glJZ2FrjdSXvAOdxSHKWd3fJAXzTOE/481w
Lwwl4i8Qb3VR1geU/Fqwk3FZCtXHLCIo20+3EwUw4b12Y84CM0qw3mc/ic7a8Bza
BmBZD90s/Y0j+iLOT/Hs2UkQUijIJyHm3KFPq9sYg490A3oyP3/eTyVC1tjIqMiW
qo4/pxwXWObqOSm4jgUEfNvGMJfS10X7Zar3a6hVJmCVESWXvLD5EwO4Ewwi6qL3
`protect END_PROTECTED
