`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h5s0cgEomTxLrE7+PUHW3kTNU0FeWybMAuHxYJIaCGgiifYJhiwk7qsJUOSMCt9a
x8gY4koV0FRIf2SKapdZuhTKZ4P0AtE2Gk+5ksYW9qMJfE5aDqx3xQKthC+pc1+/
MhsZ7yKO5JV3jaVeX3QlXosjlJscVdMSgygWvFbVRcCKqn6+c5qTs4sXQN9ZI0YA
4GScslTdIysaZYLwce/5odSB3el28m4lhcyw6A5/bUOEzA/Dq0iCNo3wiYvPXZzX
D7sfUHGp70I8qOcobSCb0jnbcerdKVO3Z7weKFJM7ay0HJzrOuhTd1QwNlA54X7R
hfpSb7/9CCXVwdzB3RKis9+YOhqX88r81CQCc3NoazPWsxtEtJTAJXh+sZSCuHu7
0cROzbkRZckn6SCKmbxg8XdVO6ATpuPwwX7KYFGZWL/k1PYF7z/rqg7a6UyDogw8
sa/Qnvjh2gh1uKIEQlL8sB7BXII325d32q2xNSxMzCSjnEirvt2YTzpiuuUUW4id
cIav5QxLxNpQGn2idSliG0dvKt2/lKa1R6ZJFjWe8Gf740IcXSBJdfdKs4WEoqiU
vLPoNQQPMwLNpSHdKj6N2ApYn/EahFXXo8pwamf9ozEXDIL/Su03N4OgrjXO4Kzl
MOibRvAGcl18bb0sKKUWcRNHg/X3vSUZNsk+TCkJcwDqDASPVE31Uy2WUbOxFILr
Y+HptyVpwyclhF4vUMYCMKiljRINqFimy54xfq/d9Nh7Zg/d9DSVL0wb0nII6icA
Zkzr1SsOWqBlnqVfr0+gL5ZyrJh7OB4k4T0mnqaZNWm+f1scsFzoKw6SUHtX9sfq
NxgzqxHk1HEmdhVTvCs+/hfoDz0jDQagYfS+qujv7pPe8r55lwD+6OH8/d4KnUuY
Ye8Ytb0nroifbT5KxZhG72eIJOrpjttJexYRrH1SnUiuPKaA8vBCdS9EG8iYsGoJ
yrXPXa3Q6THiMBPFehERYrRe1GfyBWKCn6tQvhmWsK7DHtklNCh5L+pgxZ2X/8ZJ
LEsAm/lM47ELPJTGwBQ6uLybDpia8ibOemSl5mQ85X5TE+Rl+UitmNPa3IA35SvU
rgKlwgSXmnvkeAXDBlWowTLwl1FEuq4ZMbWcxWTN09EBb1Jyj6I9+wxNJFOWf7/Y
/KibTd6lK8ZN9VFl+2ZtM+s5uivwaEOs8pTUYd8xdg1uTBg2r/KVNrN9Tiy7DIx7
ft+mRLCgdMKyfi6rp76rAjaryWKKGTxwMp9j8W7lKdaFsvbA/6xiELdc3aL47dK1
`protect END_PROTECTED
