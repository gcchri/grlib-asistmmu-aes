`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PKtexK1LUzql9hjYuk2qOwxjaX+xQtpWj5+CVvGlL4N2+SFklB8TiXDTvTxfsJ/t
sR0RP2mFr3Ll2ETFMVrfE+pZVLKcOybYr93KfkZOq1CetW/YMxe3nM0iNdDPPxe5
azpM71PDfFqIphkmSrw1LHzZ5VH2DGaC0XlAnXXBQipodv3pvGyGapsu+U09zQRJ
hWRaDf0ENg0xSKjLp9uV80KvyJMih1wlKywNQr+FIMry38ZqzZiv+JNGFHs9BkN4
tnKsOhRmSrLjLtxy4Pn3c7rqemVlNCYsBT73DxERmtAQRsGjGOKSwTWGNVZI9twd
FPoJmuyv/mmNvrBbTb8wq98pT97DAs77Dlil/TCfX0d39+yujAFcCd6fka9SNKkh
vNjcdb5sTYDUhkHyMWpNEHGsi8ZQYb8dkvSBCSd6QqtbZ5lrxT+as5VSEBJd5Bip
fSL7ZXtqhxIn5GZVSVP/F86pUqtdDXGpZ3Pgz/3Op709aBYgrLLraND2r4kyCsvN
TZQF/F2MQ+QTs6hCQDVJhcerfv9RR43cM/uB2fF2g9K9c9KdV9G1gL/6l0aYuete
gM0uIkQTPRDygWX3Fu054O646iVeXLbax/hzZK44X/kLzFtBl86AwAeNnyXEKNI7
0WsWgOJ50fLrBL0uZoC75g==
`protect END_PROTECTED
