`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
knJ5Vg2v6iqer0pUjuQnY/NKfFDooOgC/02G9P4Y1OxAQcpqyWWptgCyLaQJ/MuL
53wjCstYvNmwSGfz3SPS8AchaqdfnHMDlNbyH8ANkWIeb3v4XSwXw/VaNXdJXnhM
M2N4kkCgcwkGsVKNN476C/1TAhcy+GQWFcZOMxlt8hM58TDqa9+/WT32/UYMfVRe
mYUiT2nS4TvwzfDj7e+ioL9rGjAavghfOVhSladuQV2Vm3yBbb+zwnupbqlGGpwJ
PLqsnrse17y1LJx4AHe0rEcsFWp8Is9LNryo6W2Zb/s=
`protect END_PROTECTED
