`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SE7+iuISsQI9iZSkWUgvEcweXTlwl+XEmJxQuRzSmHVPJgXlv02UxKEgiMF/Z4Y8
90sej5O7k/vAnOE5q/cFsfj6unLGTwdi3t694E7xQEsiqHY8WAL4SfN9riYfw13Z
6RJ/b+3wMM8eQS7ou8LseI42ts9qykvBF5zkC5eTRuuZ63uOfSXLhbOguPFYmsjj
XFT0+mf5gKM+FfThjG70taLx5pUV8rCDvIn+/NWXiaFV6dSCW/sykSs3JoybIOd8
zaAnj3fgW+ykRdHIelQjSAgHeafY+KswH9Q1xZnST9IewDF3/TEVO2v1ZgDjd1t4
GMRM9LVC3u1dTFcjKrtDnq0/+5leDdVsek5HX8AIOoBP2knxeVzRBg59k4pjGpC8
AydQeDJPBhyjL7RkjmUx1w==
`protect END_PROTECTED
