`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6pBVQ9TMVWBVZOq0A8K7Nr5VKfNxY5k5L4igdi/Y2VR1tKkOXLNUEmV3iIieRWv8
znCBenTXacV0iVLaKlWc8D6vHlOi7RdEZnwSZkhN8uI4pG4jnIWSf7EzLH9OQLj8
bStm9N1kGT8ugxT4muUBhxdtV+mNyPiVHR0TMzn/3RQhLoTMWS2spTQStOhExttT
9Itln+qf5oDAjmQSohfTEnODkbJI3umlLZKUJcez+GlAVLPpK29q08LLSwfwfpjn
TCSeWyajxGtXJBdHp6ZQww==
`protect END_PROTECTED
