`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pnNuwLN/rJRpDlLV+7eWZc9WwOAlLQRdCutSOMI5aXCXIIK3gKebMMNBmNsC2iy7
XI70dK2vM76zrdtnXh/SAV90b/fEwPREUE05Z+GdygjVUSJ8LmS6lfVzIz89l5GN
7rigOUKmvKXNh0bTSI2ydFK64VNM7f41oiT05BypUPGkrAxUN9Gwp8TxVYlMEvng
wigyBwnz8ihZId1sdH83jpYKh7biP/o40f9cEglzib9OS+bzTfeEyp6GhqXHjP+d
1gYN2hJv17bkLQCUcxgGfGpj27EHavJzORPIj9az/0kDkdjTsyZUqm29JpyYIqsv
ozQy1t4BE3C3rdIlSBJgKvXxRqdWnIL96ETvHTYcZ3+QaW/9mzUUzt1nB6z3jNUI
EAu86QmW/Zan4Y9M9UFoSv8qiC1YW15VPXGC4OAgs0fzaH5uA+ZcEhoyRcKg7ulH
Ns0u0D2rICq4UKvsU3G/P8qM7xSnnBDxP73bTSCeueK16kmmU2lkun+j/CmeKfdP
M3RwqPOhObEJy96eXLjzdiT4B/w3t9V3dsfPW0kvlMHJlBERhe482Pt1PUocyhQl
WidGv73dwQTfBtw7oVW315s/zwyaDOMQGIK/QM14jOjypeKEHukMf1TTcZlYFQya
r0JK8A8GwffdBgb0d6mPpsmNxt8njS2udtgG70KAUjrGJvqA9vGttGfPpQjO0HaQ
lU1QDqH1yYwNrUnwXz6KkInffQVm448qqyjDIZh6GzE=
`protect END_PROTECTED
