`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KvhXTWJccJDS+xfzpv6gp3Uid0D0Cnm3mVDa7dkCWi5FxyuHhqN86Uqm6n5rGTlb
pkXKYetsEGJUcmMfZMoEcAxREDUkoKmSGmp/DjINJVW2C7gfOYfQohKF9bywHloT
grS+jMq0RprrKlJ6vjOUbfbl91/eLeqOdlMdFuxpHT6uohOaCMCwhcRmCMXqqOQD
7Y/XLFXe7KL6+IM7ezp5mux7XfYnrsWOjCkKBkFmZcNfJBJmblvEXqz6xQsG1AsO
7UvjIlh4WnipMyWh1GpMxaQMdYfkstOBXR3WeADAdGTrWxqUOD+qybohG+F1yk+T
YDdAaXl7oG1CKfXj4uFcmfUtzL3dd5dHEh1jSnEsN7ImcI8AfwcA3opZZ+pxA4+0
QO5DJSjOwAAwudfgZaliTOgm38M96VjB9ARmREbEuK14mDHQ9wfg+fgS6KcH0j45
1RU4h6WYo/SbUIxR9TmcRKXvzPKzCx5RGJwK+JvLkeb1GLWs9l2QLGactM+ixjsh
eXEcmCCHkP42lmX3L1BGJMwasLHxSXOEKJETByReLV/9doKR/MeqDuG0//VJ9Hhe
vOjNG0DX8ua/nPGPU3K8X7rqgAtxDbF1tXElC/Gpt3+ThIrZd0dm02mCT6fB0aLS
yI1e2D17HamOCfTkrLUw1mJCBj41sIuJNHH/zUsDb8q4DpT2jZ+7ZCJOqeUJvDzE
oSJ4O/yb7sg6SlVtde8MhXdgVOOT3adUe79cKFZP00bNXU5slapurDN042y7iErz
s2K5fzKv3ajp7Y+EgxaT0JjpXqGsqz/6MYRzWKL93jZpnm82kvq4v7v6LUPgkg9G
l2QHJpVR4wZvr7jhLYbmGbnSQe7UUAKHBl8OOUPdU6N+AMr7Zaknl5RocX3tpVkK
KpxiHC442C78+4xLdnF+4qc5b7KEz1iD1UZGUIJI9Jd2GiURvmaDogv2yH+1Vrmx
ZLSqMBMLjluHy4Hfe/Re0DQ4pbdygmPj7nFegcs0pL5aX1VpSH/XjzY7oZKRIN3X
vHX0SPPajBHaN2miBT9KuLGa1Szeu/CshKLptxJ/RKsibuoBC/k5B8Ae18hxVli9
5rI49iBGKaYBA7uUNpcPUOmr5AurFAXsR9pdPVmvcsU+BmpsGOT0/mAKG8/gDedR
DDtq2dV75fsFi5KEFsbaiZhLC3zmXz5AHdhE16h2ZxTJuiL9i92eL5WtO04jWOhb
G57yBLcM+t3SRhu6jv7nSvVWtBQ/56fg/SlS8arsZ5r1TVL17x07aXAlZ20gvYm3
024E7Alou6r+thHlO13degfp5w4aThbohfhE9V8SOruC22DPYEse8PJPceRM0MX1
qIQOf45u3crtfuc6nGe0odJOdOeep6b3M88/88XssXUJzmnB/Ic/R1jLPYl+O7sc
cWM2IlKbKNS01Uh6P9awa/Q9pm2WbTJgbkZAsGY28yB8rjhKVd0YxLwUVl8iZANN
8AQNvTWpkRF7xGSiCEJS2jLoij8yZctACx4UdNDDoalSH3jQniOEoSatXO5luvB1
MNDKv5SSR4q5CV7o9gKta8ajhHA5i+abFGEmwe4n85xKQiQyV0p6yN7enN3t5OUh
M7FqPXdmbAMjus77On7he65lpi+owXl4nrlDJlkL/29TSRfL2QjFzF2S/2KdzjzR
O2os7OJJWxwRMIOTEIgdcdaI0JEOdixXaENE7jITN67it19EduzD2YMQeA5guBxf
Alftq9D11wQ5LL/9WKX5ztzbzi5I5LQTJmdtLltCbWe1+bW5Sg5GjlDsPub2Wjj0
6v420Rl6tieEQlgCErYyp34vE2PNpunBJyPrbVLdzP/vniuSpWE7JN25CTmLp+6H
ESVa0Zcmsl6NCLnWPjLbR2bSzzNX7D+fHrvjgCyFbVQ1z+cC4Rw3POBJk/OFf8C2
76+EG4lfc//L3tYTBH5JGjWu8kTCdEaDDQJzXAcfi3za8jmwSyyriGycXPc2MNd1
WHv9w8BoJZhJYgsT8ZWt1StAbvHGYgJNo0kZgHfbPR8aMckWDrjiITNzSdxr7g18
ExZP6N6YVTdqNmA3FRYBWf7d0z073opgGg7ieNaANN1iIGE/DbrfNEml/iQOZpWL
6bAYL7A5leM85X0JqUdkCnk0VvhVG9iyJQjvGr7djws6nyoSq/6bxQ8PWSobEll7
Bvmxr7BBtWzBxVCUvbh0YqCiL8ZPDtSkWVAPsaUB8+iXJdaOxukoHV/uA1FX8rT3
qArljDxiprCR0iJ82NOQRbuVMJrNCGysKfAtwLRpG5J66KeZjVvdl8o45DJupAdL
228yGoS+iEK/Jr1PbVedAY7vklrdRjMZi2K6eZczJSgtYP6SFzHm6c2juSxgnSID
aZp0SSpaJM/+rXPd1llr+HQ+8BZuN0dugPm9v9BRUEIRuyb90zUpAKAR15+MTl4z
wVHjuo8mYwUuybFDqUF75Cw9p5tfAx3cRgNqTHssqB1cqy5q9eYDaDX2cU+bLWcM
ZBbTg3ISsTo1uX8HqnRMH1/i0P3Q9XyZQraYgtRFK6C2Sxf0zqb0a86u5477rZxX
tmnnqDcNQVoMy0niySN24Uno4z7B+LAgodye70j8th9ERMgO87yZfhLxTjOYBnd0
Rrt7pruMjB3psxU44/0teGdg7l/MwkYK1EyHR0Sv/9SPnBk3k7/afnF2WGBSKu34
2mju5Ruwg/C7+vRnUb9JSMS37oYg4y00DG22KhQoXtCthpsL2vfZUSqXzlqRQjbg
DrdF25c5QuwvSiXx6k+L+xUAwitUDnM/53fYV4rJc9uWiBFqRrcS8puqLE9JAws5
LPE+L8O+7nGh/H6omW6+hl/8qBBeXfr0N22PAWmYyGOLdvkgYDOQu7ttXZpD9xwc
JrNdbihbrubLK1YgvLTlTAqZ4nF/nWrvTwXRlw1aeIzrTm4nN7MF1wecxo4oSPeI
Ke834z6bO0l+CJg55MRQoW7Qh3bWx7osA+Pu9UNdTfdo8xUjkTE4Y0eq5K8cjZlM
Hu/Fbou2fnqyq1XVqghc9EAfnah7UqhuytlTAKGAYsCYBWDUUiGH8UxGkPFECsYG
idGWMSJkLhP4SV04D6prTm0gG8t6B2hneXPQPWrGMeFMxYZWH5X7tz81Jm+/YyA4
FUB1fsu+QBSkkTNDOHsKKWEVXtx3dCtkEf++5161YQKjFBsHBsWtloiV74d5NOow
OipWRjykdGOW89TRBgynpQlWOCTCoHkODESofCCs1fwXTCgQVRNJZS62TsPPQ7EA
PdJkbqFLExr3f0EBVKnO17ScA3+eJvCoZ+U1UFf8iO5Ur/OELYyyKjty1+I7zzs1
sQdxLbFWmPwWUptXdzPC+82Vf59APPs5fRoW63nldF2sWHO9Pos8WE+5wDWWS5LJ
H77bKCS5J9lYmVJV9Wyu/QIPqL4SWYBEEP+51uzd79fyolVTNB9scC9KwUsyiKUP
+TTPeGr3pwjpPmn8kMSf00K7W26ZNJ+4o6cKZ7OKYCH+OPk2uAUoQ/i/uG+1kbyK
Vt1Ry/bBdO0aJZmoNb5vDW6FPwL0a7f8wHxxnPVLf/J0q8ab5w/8o5xAb1YOjZCY
Fc6xnVl7iVeQFy8cTKyn3QHv5e+YFZgxSLxLLMva86DU40qQSpQOORPPWzSCNDRn
4CprhlBn3LYgNRLLUQFje5zw0Xc5kO8qbqEZS9oO/v869RBqtozM8RD6GW1EoCC6
8Fu9nyqU+cJOnynKDkiT3Y6x2dU3bdl8Ky/Aoi3/e7S3re/Nql+/SoWOYAUsqbc5
9ignbzvK5WXYhmhn+PmjS/G8HhR8JWWtpReEuZvwXW23vYER6L+MzGzFs4fUbMZ/
utRoNY3wHkMi3xzWHI+bJ9RQfPUn9UlD0t0rTCM3FL33P1+wzAVoUcmLPhlw9uBh
nYIXZoGb2tf6RmArzXtwDUrOEfgbpdFPhWnyyaiOkKpVwvWTjfuWN7EmQEOS6Y6z
yH21pxAo24yKj3mOg/yqmvGMeG6fO7OgYHnAYx9IRneWeIC+v00u4SQ4vXACYiuX
rehpu5v/cocFZbUzCm2gSw5wFLd6jJE3o+JUmtlkdl9YY+xSGR/HrEuWxpuIfqK/
nuIZjTIbfpqgiuTrKzB5a35EQ60bIiPrPNMIwJiSW9nZDCPk9UzAXxyMaFbzG+DP
mK43j5beTdt8uFALoWN+zA7kRN952kvYZTVPu1/Wghb0hP0C6UHwBQO3+baLh/Sf
oQ0zA8xXLTABHYzWTB5qtnQLJIBtyyC3WfKIxutxF9oNQDh+okkHc2ne+/ckWi0P
VpVWEbaDwj1i3hyQ4tYTFYCx+WAuO0/xGyDcZDv0duCBkCzXHPhA3GcGopfF2s3x
4R1smDmcFje4TDL55XGNqV4ZjTPoqVYk8XDKQgRQOmw91PsaB9wfS2z7GsO0k1LC
kfYRI3vsd1aU0sWeJ731tQrRDfis+QAPDNrh3FppKim6nfXN5UV8OwtGteB9HWzp
MCNTxk9HQHFYwUiOAcbO3Su4TB+EgGvxuyeED+hugzk5vRqC6nkQmQYF0dR9/4pt
aXbYMfFwo54MqK3UJRMbqqwxwzVshOmoCJ1hhsPd/O7rTcRL9YjWJE7AE7v4Y3wb
esIkkxVKz9SJEeNOHDua2p8m0w4oU65c3AZpTmPxlK88Jd7d0LI+7YLq8Xc8gwVl
2I9eZAYpe7JCM46sh6pDZwtXRzohurHzQ+nFx/YU+s2EFnJmk0ye1e6pyQ9ZhICC
3GvEho7y5ZOScFsbWIzPLE/6hYMD4ryJTHQJEnEXkdemfloA9ZDkO9CX/etfKau4
7Ni7yRCOr14KhORDsbg9xtC4VpNWWkJuBadN23dc4ev/DRV2A475qscXj55R6ksZ
4aLSt5Xpc6hWygAqVEKi3ow6NCNI1cbddBYlSpWGyuDcBZJIdH0sfQ+ndzGzNXJQ
lU7aCD/eusGUBLF2MMq7RkiWhO0WPuJfyg7RltdWIvfKKC5DThoFNnnTkLH+M4FX
S1qWLeGtQTKFbt2o08E9d827ALLH/ch7OTAAc02nw2/8474pbNKRXSq3MshfAgBe
NG87p/OIq2dqcCHeeI/upVU4eW6BGZ6PcgzZR/67VsCxzCpvhBCT8tUtJxKDLheO
ydBH97jiEU5a0CK2Tz+zc1ECOgmWJi5C72ntJJsAkPSsL925lSbaXpZJcRLPVXwg
Wz1PwLd4SiW9M4wXZDJSk5MdZVMkF3z3HFJcjeWXGJT5PHjD5unVV1UE7kjqNd/m
/zC+Gz0TimaNMa4Kj9jAeDqoyoDZj9qdzBljxgLc2FgIallLi+AZOVR4aa34Vb8G
6tXFRiYt6RO9yb943ukU58gqit51csmopGLhuFP39AkaMmH8X+3RTPM1uZk3463k
271vIqiUx30bkQ/RgUrMGRp6Is1M7+vX3yhzwy259os3naGmCrxLKve1/TRNTsWL
S0ECelPETVsliIudbFJ4v85i/KdFo+ARUpuHIDVmTVR2K0RUQqG4PEj0uXEXvW1o
n7fTkirM0nDx6FPNMIePcQsxlY2elFWrwdj6A44AMF2wu6ftIFaLbwEsoZPny/s8
ObQjj5+Mp0freM+36od7Wk/kMR4xfGPyCpIdhsOxa5CUTJ04oxohmOehoDf+2qr7
zmuXoabEu1Be7Egz8Z3/EyiSrSCVT/eFaSvmr8XUkGwIEQGhmdOilnHNxC89QYqP
z57nCps50x6z0hYn6NZqyUAhCjpHr2vExh6Yv3ZdkUSkvJ6/mJLGRiha0AdLPX8R
4nB19XIKsfTm1AU6K7aw3/2bDKGHo0YqGIpKiPmX6+qRt/qjrlJ3gjYR5zBahwlC
iLyTeL2OVvmSMtpizyot+n3qAzBpO9RaYa3pkhAQSIx+tQTilhtJxS7feAsxuCaI
89SnTq2pJzT/obxf/M+BJnhIgr0lspjZtASXgrPMclH0fWY2tqGlUePRVcKuTkM9
p64pqPXsq7GsGxHM12ix/HHjdqzKrw5KS+A9/WV9+ui64YMauOqCkA9dR0N108Oo
cxnPc1BwljQ00KON2hLMGUfLRX5BaiCBKF8n6A3EAiLDvfP0fybPrMo9NJ09RK71
6dcYRjSRrlI078A9hD/b3Y455qH6AtayouysHaBfahPsZ/IodW/R1eFcuzM3SoHk
eIrzn2lWwIsVy9uIMjvS20xEekcFL2SE0Hw9T1RNGxnjs+NkpiPa2Y+5QgrbPtUR
AeMnhB5JmRt5lw+5DUtK+kTe7RVutGYep0XqFccP28W5wTqYC1vEgLjfDzisqlMN
rm2sIT8OnPDnRypPPzhjseCr0T1+sRvCa/nRZ7V8gVrukTui/d62mvMJ/UoufoeD
Mkfy1JFB2mvWL8PCtqgVLyWf0gk1cb642wd5r2l7rCH1LjPBBT0auKHr2KB2miDy
9sbriEuMiYUkw08mADjC0O0A+YPflbOdZAM7WPYLpQSB51T4Uf6vTWHG+s01m07X
u4UekZyQI5mpjZ3G1+Q/VRNYm8oW1n70baK9KD7Ww4t7/OXbhI+OXJPkj2nep+cp
EjHvheZ8CFKp8Hd2tgM8O8ceP6A9LjySdPfAV1ukl/DMk0ow77vNpcUigry7dPBL
Uz6AsIi+Ob+dZlenMlMWEwgkwauVCFNkxzwGNL6NJXj5vV0WgZeeqltxLPbEbDv3
prvv3RTUENQ0xBkd3OAh+f2aNlJv9XE99DBOCx0gWGt8tIM6ot2DszM34dD9OEOF
xsx6VTUf+AvrqtGqP9T4GYK54ShqVciUqaVC9z13WR4R4XxnBL22SVDwavxlnjhH
F87iQ9r2ZX3lpLGksdzBEltdATA9siPUPHGT77qWYrChjwcIqQAlz7ONPQDjhy/V
4sZogpn5y0ZjEFRNH82HY3rXwSKhjFk32i71QBwUHJShD53UUPVhbRpLM8/+lSn9
bm1QL+XkDwvuk7maXlvMqFLo5lJypRoPh40Y97YhD3xKOwR+cg7EnwiPUyL8WAGV
AnVVKWfKYbEaAjuYS0IKRZJ5nApWJMLYh2sV6Uun1mvhQI7QAEDd290k2MsBhQnr
02mGU7FF5UttPoYZQbFwtDiqKWT/9O1mpO8E2myiDl1OBT2JkUkuFoZNrnfP5Wp2
4qUueVIbUQoYpjg0lwXYkBLwXkJAXQzBSdG+VJ7zK44BFbFeNPDjsLL8XE4kNh36
qZjz2tnvbio8TZP1nBVps/0j3gZYTKs6OzkKmThs4RDx9ASON8qT55sMXy80Euza
vB4eHqNZR21hOAERfF5HEloZWqE0rWZ77TW+Wq67afWbvDEOpOZ5iBLLIWGOhsp+
J07ijisuz2ESJjv8PfW/ZtOg6/fXnOCAsxqWfLRwcBCl2jrIeoHzvgNGzkuwNWf/
IBEOgmyqIfiIJXvP6BMGXeZVgNEU7E9ukikM7isNhT8d894Eont3c5kp4/yshuY4
z6LaKTQ/kfcXNs+X3I0S3OBh5VNGQBtBf6VuSZPDI1H/dvxW23Da3KtDZXVPbEHp
7RU8suZIEqX0hfYqFhnxhIgl9HKVLSFC3hB9i5qBG/Bfk1ZYfVaW5V/wVbMbCPLr
KoHGrrmmF9lgaAwi1agWeN7tib/Vgqfm9SxAHc4QK+akRn7h4zxMVlfGg+p7MZU2
gc4Ps3Ka0OvEdKrFJiq/yirrNA1zlKI98CCXHrY6iwW2TXdNFB5eXFPPz8floq6M
9/VTqkrpQFd4bafdMXkXtdho7Y593EGDvzcrxQkTw6RUYVKD+R/f1q+ydNInpZEs
Tz/QNn+QJ7vLNdzhSaYTaF0xmvlM9qOXdJrExK5l/8IP6H8kOnMAKPEdt7Xjps40
VQgYGH4fmxPDEs5j/oau0KtdkAXtmLNwx+pFC/BDxeetytGcPIJSwkZy5yvJV6g+
5Qou1HqASVZeTT9sEuFa6n/Hd2OwTExCE2XO9XpDmnvnVGvne1ck09MY4K4cnjse
l6Fqw7eYa8/NPucpkSb/GB7M6Zpe2Chql/fO4w1oYPFzraHioIGvRMg1IYLwxtBB
IvkRVrwdlWA7FqxvtlfYstlNdTtkW+HEJo8fXM3trhcaG0DbyNrfftGdZNk7ZilD
P5bsyKoyMXFEGuBLRv5vIQNCfx2gq8PfgQusrfvwodNn/AyWGJ+LNmOj+KhSPeqz
MxjvfzEbgUV7WkO3twpvb6zTLF/D9D/6H2KJqqw9QAxDhmrvP/lgy/pflIxCKWML
k1BdD08l+IIF37k7nAieGbSmFt7vAuBAtnSMdMLeTaT6EdknC9z1NUi9jpNYksNp
fMuqvQlp5GmFEqQfhrFLUTuokAOYCowajizJZXekHflvQsBT5zZfvyC5i7RxRGIG
CexWqVS8AfDQWND/xhkEE5sU7y6gEgO07uMam/srf3i2RYB+xdBkqunRtQ2sA8jY
+5OwJsAB0KvbqHNmmzi//gzX2V1dHy6ouT3yz0iH76Fqcd47cwHoaIYRXXqq4FAr
dOQls7XyTnDGOOMbpdOuNqpE89pL3aDqFXQFdG4qmyz77lBpBPjnlDXR4Wmzm1mS
CafgePi+rDDy3qfiEZ0wLyGIaoh28TCdTadTYLP0czQuEYVH+qZ51RsJuiYFxRQK
vTGCq+Fs/uCxNDWIB3W2JxdVXLoTuiU/fqig4EsoUoZjEQPeP8nwDMxV5JepqbIo
BVUWV5XQBIzOpFJBh0Quvmx2fbV0jWyWYOfypQoQ0+/L7e5a9v/xI0R3DMqPW2xI
r5nEubltpK8yzvb66rGp8d1u55m7gXuLoM4Q9Xc6tyaKwbPGS38LQwMNKrGPL024
AUEZM99IkQUgCU3MrME0JVmLKaK2nvcA+di1rtxHJUaAGr0dohOjvIkyBrUugxv5
IG318d0Rb2QSai5C2Vn/iN5MdcTZMHgCgjKzrpe/hiWG8GuccrFdC+0h/VflNtaS
bRszyYzcprQVNj7zi1oo4FdG4D2AzbcaGuDlVwB1gyxdUvAScvCbt97iNfHedcqx
ZrgeNcgGRsnpMDUhmxH1YfTVoSQyrF5vaOHB4Gb+j/Jox8ndDt12Ih5zGxJrouj4
xJkqzsgnxKLEQJKlD43IjpVGd9U1LLDhdJhxkCBDzUGEjKd//rJrB3NFQX6hOQUF
ext2Y/Fkvx1HyAugjqf8NOPEFsapgchG546yLx40ZTpFyJwDiV3/Qxftyd6DcULv
36ARdphKIklIcH7E4GZKesvdK7vX05LSMLdai+FJnU/EEH/Ae594ESAmZ/BgdeBz
KdO23WPJEDCXoXEBMMiT/SC1EOcLxUKvmmP+tyY1ZRskgTBdq/rN/C1DeXPYTAes
Y6YGOHtYKuuACoyAvROiSZO1N76+vFvwoCJT5NpUIRRhnvHBrUvIqZAURs8XDijc
ctr8d9Ba/OsUZd+BdIUSHwq14FkHr0hMPCS4agWDBRrDlr2TeEoBp3jegDTBySfk
qpuoFqs+wyL82KMp6V0ZARWn5Dk7VHzl1Gtqrk8n7Q22qoJaWUd5yM7MZgvklhQT
Yf7alEaJ6af5xQ+5QnX+V45zGqLV6dnZ588v5mPM6Sg1cbZ9KUQM5NQf2wwRspE6
LfHme/MCjUmOS5w33fRHAZpWux36GluCxFE4nxWZ+Of8T0EQs934lHnZEu7pNdiK
ZH52qRCRwnG+sHSYkD0m+ePsmYCLEp7OKGdiFEg3gZEa/xPERa+5IB3rfQpjn9ZF
5ALXZvuu/SbapTuqy4SPnkYiW33Hcx+19BktJQaL0zTa6+fSOPJiaZgQwqjUkLqr
s89G8M5FKjdvP2PbPIBRKMcZZcxtHSqtqav6aFEVHbCaUhYUSPjy3zSf8/9n3DGd
ATfMmzoz/bXTmDXhgh7ZoKXpPWeLSdGk8BqBlX1dKzrTx9zeQiUBhi2Bk99Y6h7D
QVjTI8LwI4GfcduBXlt0y1kIEKkys3CRRYifm46ZPAI6u4x+hDeLKarhGkecV/Zi
pkBPn21FedEGAL6ggx+bQCsy+3AQ6fLmKQXjcXdNzb3zX1coBfayOGdkoEbaPvU4
4bwA/6jiF8gu9On7gqzUjUOp3N2Y3o8GoUhVP6Qrvjs1KeV0P/0xI/hzFwnagleV
5jFwTr0QpBVbp5z7wnl+xK1vmIW00B/KxBkiSyXnT4036GQkz3C5klTsMkPd+XxY
IEEteyyiU3trMzKxso45tR2BoCfY0l8iRyU4CwHElre6d0FMrtOQ0M9j2ObS+O0v
enJ/8MIi2SgPP6vGBFTnyEujUeFo6z+hBuIXcqdacgDLgyswaMYlKd/d11eZkJ6b
3BDw6a+K+5LfW5MNNUmuvYPAOMDDMrMeeUYRYUZdZZDZY06uemV1gOkz4nWpitLB
vYHqEgFvhEpxwmQoyLsnOtzaFKcnUISrA/CDhH0R/5iRFMPB5lv5s5+tchIgwGTQ
m8yR23ercsbl5Afmd0p776XqxwfcIktMTJqc4KFLYWP3p5cx3ENIUPfrmi2xjvbR
LK7XYB4ZbWTqZSSkHXSReEXWUakTgv6/qXk5lygJwEeab82akZwsOyPy0Fysx+jH
IkJjV0onSBLSpqyXuDdW+A9JPpW1CVSDyrkkzfwPoJlMbDbeDEfgTkVDleWTde4V
QFqCjABqpkv5hWFDCsL8oVgI1cPWcp5Ji32lfECGC0dNYff6YWi7v0Nx9s6mnoBk
eJ3cgzdTh+vLOnQLXKLbkk7rDCNbNoVK6Oy7frNdYuNDXmDnAG8sJ7t/qg1eYvUn
FTSKJbg38Es9xHDDoFYI2yrr0Ylzth/OUIK6xNuRS5O84xubjTVZVE7s4rJEbn7u
A0yMy1ZIUBpxs7nrXaj8UxcRrNCrvMBZW3JUizoNouKOKrcC0I4mO6PyOpJYgJVC
UqWe2nTDFlKdfGHU//FO51X7u1tOowo60b081sBxDrvnKTj1RxUJ4bNMUiGJqwkJ
w/Ns0Uda2uTvC+PapjGleZDtl27Feub47/IcYBPX0nxwZFD94cckpKmSUgIfWw0O
MGeVmGJo2bGIgSY1B5JR0fb7s+AaC32XX9x2q1CPBKBRZcimKqizihDZcYVsYF4d
Uus7J6dZXraAGwZDgIZn4GQ/KmSXwT0ijcv/ZdiwxpjBUDP7JlHG/xxLBBPUMY7R
eQ4cZTyLviOAjBeQkoPLp9vNUoRrVaZ69kIcm/C5N4YJBmv3GH8XpCNfUmqKSMoz
qEFMzbcpBCu2OCS9RPRhngwx7eMqrG5AEBlHjC71fEhcG9rTHv9brfRTLlFAFmbS
qijgcuvl+Fsict4Pu1I7v665vHFAPQX4N7OTwfsmIfQsSbiXlHNVYsfNzRJqqaB9
9Z4kDZ0pU3WIF0G0cQGm/DJvTPiNvWbTp8VBNzflG5rKLatku9pnkaSaLY652zhv
ReE7qRdiPeazjoEqEUgkz57Q9i78Tszk+Z+B8vx1nj9Id8zG2jeWEqCChhpmKWtq
TfY2Y6fqg1+FAOVb/eT/+1HeUdWB58ti2lut7gcyGxp1rdcLlS5SdnlsQfHrSvu7
vmGf8E1fFOdgs35jiokNTZxHKygArzYwRqvlIhrlncBcSW1tdNUIXAPxb5TKgzTe
m12xJ9qaaAFKzZK2gCs/HED4c6geQsZmO4EPiIvnjC5Wxb+nKURpjfxIUYZ0EI3P
bFPTY2ogVN9B3wLw+VqpYapHuWT+EUPzxu8fx7giOgjUe0s/DtayTrlUHhbB7bM3
+dvi2bplBaAmYcHvah2BIf/pjBe8byNNRAP/Vfl2+8NSbu6WEXRKpMG2PAM7QPdG
cuwte7cawma7TGEHb+TqVRc4DT8QKxDFlaq4oI2xYvjmsur2pbEyy2iotpS+c4m3
o2JmilOBXu8Y1Voobw6TKYHB+eJ85eQe6YMpUXrss9GqmApc/Lh80VE2oRJlYwQ0
Cj6WQlhpPgLrlu5+sg+lctldKA+/s4svzAAInkh9gYMKQIEWx2iko2Ng+JsEHHyq
K3RJq9CffcvVzyoQMKFW3CmOKsVHY9roUbok32AKhMaV7vFk/FLDx1OFApDbUvw/
TsGrp1iPnLNOZhm3k/lZgtPb6lXhSn4ppyGXFj7QVF0vxwYJxesRZVQ0y3Gl3fU5
IKK/H9Bvki1jVuhNGJkGD7n+56xjJNi02JU7Lt8ahoE5QrVBQFF/NN6G9wfH3y41
MBtfxNXclc/1Ya88OvQvUjdlCX5fJUdHJ18JPIBXQPwkHrmPW7ahgarw8IIJ9Otr
xXaiOjdjXZ5tEynGcwe0qYsK9lhFBR7IBI+9W2MeZC7Ggu8c++vqhX1mg1HdWGA8
JVdHqImPKg3mzQlvfSWD1moJkl05BjVCvwdoGylLpO2eE8yZZo2p/OxI6noBofaz
uKrk1wVSdTbDvdpNulCv8wRyhOBih4SJvJUBaWAfSydJYgPHcb6847/i+T81TSgM
Aca7KIE9mjY+WypRP+RcRZSm3oRcQJTlaQDKGgEJ60H6PTev5VFLj1BEwAQ3WfJj
1yi5zN/fHqvLy5HJGYJ/M/4RSPkfgKLW9bkriubOOM790X55H3vu7foKDa9Esdei
mEOOWGTozHA0s/W/4e+ypto4DF6rB3A/XzVkf2oAhOfQQ6QzUBuxUKei70B9zB9t
iCBUqzh2rPLenWGZxvStdPgHxWszurvsfX1q9kfBHj/4tPHlHV9BPdGqA0m/GXoQ
C2PEBSqdKxjMktQkyjr2dgyZbyZvzCp46JcXylVfHWnUkBo4+6qzhQpHMfrM7eqQ
0ilnCF6LHxCFyg1TCGKaxOHXGyrecfJNXWIuWVaZ8Kv+yvLwOo8f4sn0PPLfeAoN
T0FoZwsndiGNi4RkWsS+3VxJjaPORYfFfcnXKSbyWmzG3Mo8jt9F0Evt3oIPT6ur
vI88AgyJzSwIxdaBADdpNxR7sawUSNgjuK5T5HH4WGgEVy4ME4iplh+kfkYjVSFw
/+DFjwVugMK1h1dSETlcu5gANOuT33klkYKuWUluxXkrodLh5r8CkPFkykl7amCi
4vc0hyXoHoJlA6dxHcdgSiZxC7llaF3KPULKv4tG8LYhe5Lw+/LdWcqbPJYhNBo+
S2RYv39WwMmjvh4QUwGDfYXCMamejl6yG6tgYT6ollYgS81/sMKMfniAQqizXPjr
V5KGcPCSAHpJFSs8oxGPwg2PBCuoP3xkWgiWLRT24GlXpbMKhCXRCocePx5QZFvF
4g0tBBpjqqDhgzj3IMVWyodLPF07/QDrCzobMMzKtWmd+BmYTBKIMNpUFTBSHffh
d+2li3TDDbzkDHj4TM4v0adwNy8ErNGO0VCJXqNzDSDIcDdWz8kZlCO/4vaj9IB/
UKHZ9/hcR0NhhcQxg845n/90JQGdOIaDrjWLHdvbEDFS0R//yayTt//4mSu9FzBD
rf23FCmIVkrW9zkDai/Z1v3mtGpzcaDzxT1CTdmQnGUsz9Jn0xw1aGy0jSHJEQX8
J1zcViOoZTBvCwiKb+F8oB2PbkbAlsBZHWtL2+B8QwuS+jj+tZY4r1or45tIQZIp
wC4OMUl3fZRO5vyy2lYCop7voAjkuucIJRZSqWI/MDKjLOQd1j45SSa7qckG+lG3
00CCsAWvkKu8LcVtiPPiKzz85KNE6q1j+dMnWH84OoYjJ6pzFOQG/bRAIYzRPqXh
K72uRc9hBOkcLdzpFiFW1Qc+JmqiCpLQuSU66rqUzUvElICNkLE5iQhQKTIB3JtX
Eio+usyLr+ddAMmYflo7uDXuNAQdEH+GKXDLfWYW7F0NtEcQN+pQ9Ugxt4iLTvoa
pOTxuKjcvAkFRbOAVp2VnOMWLxHXc8hzNG34VEtuQL1IozVMwP+2SFRv75LFScyX
Ht1I3h+BLAmOeNAvJI1aCg5ui/7nGHZEFQophZqzGMWV+Egs1IGj9j2KK3Ack1HA
jHB9/DZx9Hxg1fvrhG+qfsFZu0a4eD7v0g8jI3frFQ+AzNlW1GyOxz9YlMz/VPVT
kLlQMbcP5SZn4e4VcNq0UiVWZ/eHFZQzEAMFmB/q05gSbUTx1gxzh1AF6LMp4+fT
TN4BjyTmEVeK1YA2p7S6V82GYTClNXr4waMtWxLC70mUip/YiNO0bpSihIqxOCUc
WJJmhjJAEiFzV7A9vOxHD4DCBy2ejsUqnPmGnc31E+KDgQYtAXgFekLyV3fXk2+i
QgSWUdK+SNB20V3uta/lxoO//mf3NV578m1NFIWRTUnp8L3I3nWCcTgcjrD6kqGs
UKQ7TW67SS6/qe3zlr4IOjaPHMKE3XmWjSgYB/ZOIwli0Ftmej7EYVD5W2Q/mEGp
CxDdivbTL+4vRRqLTmZ0gShwbsf6NY0pLeNmV8zU1pqtYlz1ciCVrsyw6ipek9lE
+TgyhnC1zDff1lfHRF81lOa3oMqlmicpCZk4gLrRhd/775dbcdODbqln+hDodK01
h4Gd7LI4bNZxVNpsxCFxR18dH3imU68N4yxXH+HgPQqNLdHV8jQX+hdGg1zq/cHM
2cAdyd28KyaKniZWf9oXJlUx+ZHbwKM6odBLjcKjOLyPbjQcxcp9Sf+rHXkDqN/o
YsZkrEd4wwtRomENaVCN8+MsvYAjYpSUem03g+fr98Tuo/nH0t4Vv5AotARozK77
1cIdsp86izRUbQJiZVRwP8GmLnlxCRnV9mON4G9CEt78mHeH/N0QQRmSc3Mj3MAA
nQUMZOJ3GFEravSKme2Y/8zoOuEPhL800tlBG5ZFn/LnL1nXJBZ72AJDhjm/P4LV
Mmu0aZMiB2sTf+2NYcdMePgJ/o+vvpIziBCjUR5AF4xS/Eh9rtr9vhok8zTopMzj
6BqHx9e5Hm3aApveV830YD9G1sA/BLBcBXc0EJPEnSvd8Fsl/2lh5PotxESV3268
O0m/Whjarj/MaVAaS8vG0mnC3Ok7rFHg5Ga3IsetEyB7cmcGFsCejvfpUNt0bHwt
nR13svXq3ejBsr/LZgM/nN5wiiJ7B3AVySB4pZl4n7rUFK6QvOnK5/FsR5iYjRlR
Mul08AHNiruBtqqF5vpfWn8pF4J8KTxjtpgAj1YGG9CO+PVsIozvLZ67QDI2gU0W
MIR7vibyk+5vMkhjwDSvzwfoQNDDo+bW1FrKdX8WkLcLfTlr6wQTZKP1oaaLJ39I
ErUTdXSfftJ/6tPyYHh7OMZPXV4Xvk5PaLh2+edHxjEiZ3bbQdexxo6SChoj+Fb9
NUnQ+7w11cNm7jpt3iBxtrtrA6ZxHGbsUvY5Q8peXEPO3S5RCWZ3WsNHgMTcbtGZ
qNlNIboRd4zwwGvMfp/6ZEmipHMPc9t8t9rsxYWlDVXisG9L+gCksyT4vpjLSpN6
g0V8tX5P5V2W/dyOdd16JYsEbHSh8lDeGAr1rPy1euFh5D/EtqgbtYsnF1vrVd+j
x/jPFICWNmxd4fS6tkD96GksvKLxHNWGMh7AJjyySIJ9TWlXN4sdouKl4QFZCPKH
EmLNRYRhDxZuBrD8cV7mwvkna8s7tf/WV2efTgIZoSznG7cEMoH3mm9eEmfmjmlh
4f/TT9XG33uIvFJpT+Rfyu/VdTe2Wf1ncPYketgVa1TRHY2FLOAFuD/GSbZw4nGS
yNzmNdGZbnXXhIqxgkDPU/7gMtsw38c1dOZy3RyCm7u63EGvNWAQmyrLyHQwjSuV
tllJovuVKHA04NO2krUoE3TnUUgjMNoNh6NQVXdeHBrOh16oVCTn9BGqdKTuQg1K
N4JGcNdGn9UpOYiDNTJUPjwPUuEeJJUPzKGDZY/dUn6ihpcMDZ7UKZZbDwNbwfOi
AA5u+qbmTRcSBVo3wE/bTHmbvoOnpAMi0+TR78PErj7NTHqTC4tEzlceLFY4rsF6
ec+fvm1aU9sJX50xdaqHITRcY9xA65sdRnS0p51MR30LkA9hhM9ZYbWlQnjjr4+C
jM/UkX3Ld3iRDUua3LGTiH0OTEEjwVcLWjcM9+t9h4+VbQenonahfmP5iJ29+dqR
RnYjKXWW3A9FnIL0pVI5SA0KDjCSk1AWnRt+xP/PyR7Zau2YQwI0HEkzkVwt9Xso
hFE0buJDiQc2Bb6jCAX9uH1sDtOzdgXcTm3QmipD88gBdqts9u+hmlTrDryMt+zU
0XE74L5OZSXfCLKbbE0CP0XSjx0p4IqxaXm0OYD1N9niobD30IZbJeAi6tWNWLmo
v/Z4kvYgoV1AHtBDGCsZYeJh6ezjKwHl9zjMPbcW9ZXaCMPQcJJdCzOC/xdvcOU7
Mg4WsWg/rYtN8lT+2rT3xbXPZCIsjQYgTezA6jCrOLAajTLKP058+SzVhrJZHCKL
KQ4x/5Ng/MYMfbcS1jTgyFwxSya+LSdR3gAaZRjwdZOBwrsASI7ckJw74E/bjWa0
FyRM1Ez4ulPtrN7fIuuOQyjMBTf/VugaRyqTEWCKI+Atu+2dFO9zGZqtcqtg3CNn
rFrms7WyqLJI1DJZsnPIj2h0vJi25LmHzLHwevB9d+cssCv4zriq5Dnh1pyXhwLU
eJeiC6AStrD2I+7tmKCO172bLdTC6UJYNnHsPT7pKukHOMoFKFtLQJ/gbaWeTNTI
yz/ChtNnVYr/x8ifrQOGQOWNsePhBZPtDsc0HwvDeIGGoNt1F3t1dQUbkKhAxoAJ
ODqYVy+UoSfjbSoBY31fuimCMv4OptYtsaXaryrWS0j6ZNmyrUUv6OohG2f8fflT
7RSCYsnQNhlM0p9h5SUwHUeEuzs0RNmVBiD+Ubq3lnz7nLltEg4VvnN2znZReKAQ
75RfykAzxW6sjuRj2pyoqpNs8p9Hg+eY+P7UukSQkRLj/ae5GtipCWeUUmMfWA6G
VKaC4Ry2okjVpSOQjc9n4sYe9MheAMJR9JV++4Dk/omXkx+0OOWEq1Rck0OI96Ir
XhW0/66V7Sr2erhM0CC3zHjJmnfXLiYxY0KRT8znI2cXA2Q2HjoTozlankqkUKU9
xibkgP7n+HZCg3idksX8zEP9CK/HRwTGV6ZqdUVLvHMSwbbkURd4vfO60/dxSvFF
HEvkRG+ISi7Fv2Ki4/Nkf/FNfZdMFJJHR0qa0aLkFYjK29/EJBWjlbjwGR5UTUel
ifmpRYj4LnEtLDY7IUBTvisroRaRveFnG3FviDQmzF4t3bIcXIRsJhdJg0dNiw4I
GWVcTO+yoIQ49rBwx148Ex43pLA7Vs5b0ow1dWVajn222FSbamR/vMbBpxrREy5n
mwz2STkG63myWKBKB6m339QViCS979kx4PhpX2+zKgUnKk7jksFJxFXVEiaMHAKP
byDCWkQWykX1j/K2f6wXpbBWdlYCpyjiS2MuR48SVJ0UzbAlqgvsf/YQwLuEzgCo
4QCiXXTxwtPW0Ra+iEMQ2Re7JZHwR/gL5C4hgZPLDm/zr1J7wCUiUYgs/dhadBPu
cVdOm3Frm59gN1j4iWqvvv98HzSCwE96j2gkButvVLPASmerB4fFb/JWasj59CqR
Y5ZGhdL0MmDzxxNWBbFUCPUAACxsNMjGwxiRFwJMvyOHM8YJN/a8AvCxm5l51OX4
qM954q5XluwPwsQ2UOnZygAH2jDOrkBDUx3f0LDFjFmH4CihmYZg0+hPFSmj9a33
L7VnNpmAW5UDzUON2XUY5/tzjattA+GI3q8lc2OIyFox0YDmzG3oQo9MkaqBsLp3
Jur84yA60sEWb2/6ua7i7aNsBRIM5T+IovTmDP6BKfzAwD6dnkLRMtX0K2TdcKBr
VtpBmUKP5QtRi7V9sMvnJqIhctds099GBMnwzk48+bRfNQrwY8xkHV+iD1EcTZAB
3zQ6zA4UZvVmHqIEjXUNpqDiDM2RINxF/lhdCdEU+tEAufVwWnOaVbuTdS74QkdN
ZzE2eOPd1qKfY+XeB0u5LY5EpDGc7PMdLszAoXZT9qd+PhUgb7j4AQeLaC7efnot
y2hDeY5BrcS+xRkM4ZaDTJr6LjycI6pS3xvJBffIuMtmRtrzanNUae8PfNytuct/
uGMk6ViW6WCPaMKsXjxZBkaAaTK4g5YPWG78paSzQsoc+lISnfehjpL1Q2FFUS/o
DBlFlq4au6X95f+XmnXT76ZarmkHG/92fJA47N8q54i2LlepyRAzJmC6JMgPEJmz
Tm0VdLEqx1M2oQrT3Ja6L/8cJ3i9jtqHbq0J31sWE1V0ho8gbZ2oNmfJtT73jU4L
DBtEKZT40Li/dJ2arVOKzVznEyBpX1REUUi7ZWmZeIFEnaC7WJc6VXikY5g3g/dx
hWTnmiUVn3as6zhtpGySQ1+BS7+cdhQBdJxjb4KzGnFa1hBgXyLSIrLpri0bFH2m
VclMrL4pMP2EAJ6O0LGnHNepHqEh48FRahyIPMM/vBdTWKBApbWSk2TuOfdUrmkj
SGzCL5Esai1GcgeskT5ov7gxhmn4Jy1Mhho5wjr0K9+rT+mbxkGv5jofPGg5busk
IonUJaIsDUlJxZSBbsGrJfddLQxlYqfZXW5Dg1WspvpySkQmP/ichj9wDBIZaKVa
wWmorYtisStt+YG3T+tWBep18ZZ1X9q73MT7/WMGdjksPVYF8lrr/6cFmWB8iSM9
qS+i1Lx1hiFKne88EQJiBNT5sgkTOTr9Jawv/FhngyTtqNAqYVeinHKZJo9TCW3x
C7BHsUQ3+iBWu29ES23KwJMWfd2/ro7/UMWeJEDRswJDuIFiIQH7vEaaEG5AxEyG
hkfG4tyQGqetTD9IYTByGfWUJL1s52EmO90dZLLiMcBz/TUYtboF2KPhZWfuFAq3
2cYMq7omvhk/O3pysuhRZCwhRQLiMqs2OYEWp1GQnz12CMuhTmRrTLvES1ztp/Dh
tpflA9qzsrcTgkNvH+vMIZVojMpOSYvFjpPkwZgJcK/xZEBYZTjS96KRnwRc80HJ
Q/JYYESPmYGVOQSpJ4xV+hrmCOObPP3XOj6VfCHeXIB+rt0obZBrdRtjgB4hKErW
D8eNA1pr1bUEShoOxZtnqsa6WYOptvgshQNVYo1OeLSydGy3LY8xTSsJF/RIy23Z
ub4saBJYuRwv3l6sazWYUB+DuQ7JGSqPNXqWtZe51YgJd18PnY1T5wPSmDCWx6fi
8HqRacLVZXE5Yrn9YPoUcbKhIhEKrqg7tsit3E1NeHiiNmZJXflcC5PMxhGGvYjQ
8V+aBwaMgKjIb3uWETYrRoOdPX8t80BckD9P/r37w0AhVoW54UxHBKk8Xkv+tglq
vrETPe12/YBfxyZFYDt1rIO+ppQ50RcErN4pa6dOq7Yw6A+B20126LEoaY9kJj9b
ZtVBqYtxnQ81qrn08SqxQ0yLxL3JLkLw+ISupyBNh2PvIzRiR3/R6vGXz5cWk8Lb
z6I/PKbg6Z96I/p8KirhKZJl5OxL4INT7T+6DiIDdBNlxhXAGxf8+ZlVEZ1fuBTS
EatDvtMgmnVSteVhcmDtcvVHsERxJfCCt4PFuRH6FXIipvIvh0oZM0Fx8WGNYUEM
8iMqS6CqoD49FMGA+mk9uEwyOoq/hf9wgDM6exPxxrivuJojyssLH0a6W7+pgYGR
FOvRrVjp1uwZKr2PoA4e+J/TPCyVWokHxojAe64rXTOPaz/fYpwsP/8LAJUupWik
6InCMUeizBL1Lpp8jCRwXDE94EzMxgwpVhORzSrYZRjMzlF1HpJVeU65nrJV8c2M
c0IowPSdsbqu1g7rVypXn36W4TM5oKb6eQibr1fYdVbTU9I2rdyEo2/SHxyUTv4U
3e9rc597T6Uitgtf5MiJZchxazlDY3SEyG8BpAjLYrOcSuWLjpd5gH2O9Ng89pB+
pgzmQ4KveUPSqaWSM+taLx+xWKeTEe/kzrHguZoZwoaNESMKSB8wYC/tgoaMcIKJ
4Crbxf8QNiBbgo8o5X6gwmjCAzyBefaBtEiAv24qO4z7mtBNCrqJfJjF26YT0gG7
FA+6SghDPoidcEzHna8gSZGGuz8gFLE4GiwHrilTZKW1rCu+vy5nk81ZaZeDsOkO
VxDxgCV6h1xPD9CTDtChVUzfxNhCmvlfuMsIKuVlSvL8s1J7mGljBaZQJKqsrPzC
o1Sp5olyvOz34tKT+ZVds/pn5bmWx5/LdXTxFJZrtQd/ZS/MzHOJ+GDzeGHZZN8j
+tQFpaOI0W7n9uzttkm7EWAQemlid4JqO8SL9Ntma6ScBC1bcCZDi2RKBwsFYdqe
sG+G9rTmyxsLxcuPdQoZm9xlIREMDoozlObeNWI9Px0=
`protect END_PROTECTED
