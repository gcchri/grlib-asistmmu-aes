`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zzff9PhPkVhdoo2cxb+niL3/iDibnO6ZSdOOZDA8yy/fcahiXGICVWxrpA8BuQeH
owjgjqr50oNzc7xjcMKdRupa0+UCkMpv40X2Z5xqMGC7UlwelOhgOP0SGvOJM4wA
NoY9qBkMH6SJUI/Wt0SjGnIaSzTwtOqE+E8PjPYOO1i4gws+nY+wZylv2QuzzZbR
LltnLRnhd0zomaeSJUnJZ8C4nw291IwEZtYKMu7dLq3dXeH1X679nbGH49nXJc/U
9lrczMFOZjogSZW319XmNN/5JS4zOW+nMByiWYDx9u6vboXFSyVB77Kmuwf8J9Yl
FlFBvllztJ49NHUg/gTcJqUtir+JdrzT619i6hQDl2US/HnHhN0O5UQu7BrQ8gtn
YEk4BHnWNl4cCgmUp2dfP9GPNi6wfScNtFeq3pzHYZWrISVpztH4feqRKLToqePN
xrjoCLBABa5+2cUHDl5T1BxU9quNNbzSJj3SplwdTGnSsgihDU5UlqA5I3UMgMO8
/K58t1+5G93t/4FyLvFkW5rFrAihEdvK6kheOna1qLw3/jRE9UemYGHKvkyYggjs
6kzoHuoS+klQ1lJiUmpsgADtysX/+iCB9IsIJQ7mzkwH088PpELYmkiok9Kh/c5G
6wQn79E+jPBVOAs3JZtF/ItLONjZfIo0IUBWEpbcksdUvCCPEA0Nk5C6hMhsRc2J
1JT4VxAj3VDbwYRICW2ei8FbBVcn025IdjvammBgQo5W3lY4FmxKcjvN0DFtlBLI
/rgdnGuk3fZ0FH6XtTcD8QvUhGcPhfhjq9HanvrnKr0tyV723O9IKnR+N00tgbLH
3VpJNGjoidyItLC4gKMjpN/uCMj0acnJQ7eWBC7xeGfcYJicJYMYQ90L7tDHQAR5
uoXwo9DLczPwjYFwWERwXyUcVNqRNNq7CX6d3Fk4HxSTJ+jkkGFAh7NMdKoRlzEw
YhNAk0J6LWXQ/wkyhmoAD0babOxS4oJF9WG0YlJJYppkMrVHyDJ3ZHmFGaHvCyRC
CGidlvY+EHDtSLwDXo1D+EaDetw0tXHb7czVqcQfWD5gZhMwYP/FrctpVG2vXUeX
t7CCiTuvvcuAaK6agqqRWMNN/UsnRJZD6dc+UZZ4m01yCspFz6Gl8M7T6SBVpvFP
0nYUrwOzUNRfb66YH23m63tajpkOpsg3RzILL3/yhkLqzdNV2S72fNr0edneH9UA
q1nc7N8iQMfuIsOpKen1ntxUxg8nm8v7Wa9RuOYfA9SdXIIx1R0m29t269jlpxv3
aM+qX4HTXF9C1mouUMhRj5oXIGEKeaT5wK6VLdFOSkAX6egUEtli28u0B05l4+jV
gLRXyd8u6muUb5IrJfPmJYEoOHVeUNdsmM55LOD9z7vR03w3qLr0S0n3NKNaYY3y
UUOCJoVLkGvpTgiV9XTkXCSK+Mvy40/+z0IAvzXsN5un3pd2qrEMDf1Kl7DieXgq
FRDo8eL4PyeoLgCFqCW3JLD99zpFVTr+OhwG3flTkA9cGaAOE8n8InIjPLzChKZI
CtG0sQWtdcfoUWswkIP6q0hn/TPSqr9sgGKRCegRXsF/0Ac3cYB9BICd26uqOzpu
45zOCsBbhD13bWcjldxUWON59lWbBMvrgE3FdiQIImQJ9DBIy1UeADs+Gw5t6MEr
9TIHQJrJDSBcu9J3SiDRJ4+TH7xJEiulGyJnB9SO01AwBX/IhNGV5jjzs5Xu/Af8
tIZnjPCQiop9UBVR/HCRAEUo2IuGVB6LmHTHOqJZC78=
`protect END_PROTECTED
