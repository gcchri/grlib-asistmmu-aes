`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DarPAkxywezg0uw5/F/yZgma8sxaZ/hv/AwA96Xov7I34oj9mFcK53HptSEjizy1
fni8Yf6Nv1hhyVd9JcdXGS/kNYCbCuzerZjUfpN2e/I+IUa/ZsKkdXP+ol4T//L+
pzFGcYA2MIr8NkkGWN2KY/LbT5sOti1uyRgh/CA9JhcmYqNOAbZh5HIh/+G+64x1
ivdnmD6C7mFyRAgW//3SMUxdTlLnu6qYB/kceRJfmSWKzAUqngGzH54xAnhGwheZ
i14PZtoDEwhjrKaIFpNQoJw22NdrWGJ97KoAk9wwGw32WlJl/wVb59S95e9YKEmW
j+o07dS4TqEdBgCYpPBh1bP2dOi9lPVBeLbEtp40pDI7TieXaAuBBhdF2KJZg9/i
0axVtDwmSxiTERkzVQBpchwYXAaaYO37356Hv/bznSsjOBBUnk9jB68+LVCVXUMd
C6fh9T4UsGWS02JmJotuXIfGWc/pdPq2AIiLwQQRrrkCDRPiI2b4KKll18HI+PWB
68zkWN8oObRxIUheZt2SEfgS1asMszOmm7wYCK7olec8CyGxoZ12Xpyl2OJar00D
gvQBiyoEHvwI21JmcKqCzw==
`protect END_PROTECTED
