`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BlZC7hTPkF2ECXCCmAv3WX+tam2jTCUoBIu6811fqKaStBD8+DSwoi5TFWZni4WJ
8KuvBIV5BEZJUthHiDhdTUdtY5GO6vO9IduLk5k+8D2UUysHUXZG45f9KmdWCFsR
AHldz8MVRMzE6V4cX1ybLFY2/UN4tQAhBa9ixfbM7aDo1lMlw4U9yWcuS1zTlev8
1oBWDE1+Z4wycNGoMXGMUQ8GmX0Kpr/4m5vkCUXP+GLv+E7H80yJylhRiyyycK/Y
zvpDIjb2e/IqsXBlfnIXrVumPRRSjAvVYVjlhtMZFk29e1N4QgLnUtsEYWVYfn13
aL5jsK+EAkDQJOwbaWvVnW5MDfeeL3nsHkr6FuGJpBmgknb996om7vqQzz3ljP+N
7YlpoMArAmCjj9r4xzbCNONj9RzPWE7+Qo24yFLjawqs9qqwlEGK60YqDgOsHl9f
WpHLBP9kU+tbBvNctwHQVlPnjlV0J5OMUhUrNe/DkWWHcd9Ynmc8zXG1GnAY/vYV
+RnPe9+UZH1uWSkAIICzRw==
`protect END_PROTECTED
