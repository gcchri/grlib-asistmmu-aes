`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eBAswfeC/VkYzauhwAsnuD4I5tQ0EhvxtRdQGvEAq9HSH5SYBtGUQb9ZVF6tdUx9
s2oGlirA4jUhVe2vHrEfJuOIu3LPMQ/HH/EMmlVeuiqKd9s4P2Ix6LnCL/KQU1mL
zzKaC31k1sCTCZJOrbH03qMh7C8fpnILF7sYJ4V7jlKZ9R/pWkK8+SpNoIKf+B3z
poPkTLl3eZYK+gxosV/9yJfS9+OskPyQYhMSVTs8NvP9yGOBzyrTgODqYymCymU0
vi7fqjYOoByYHWNmaK+D0DRJF47DASrgUXh4nf2G+JaNZiqZde5S2WRONTQ4q9i7
mdCKm3SMBoQ4mnMQHWloOFG42nZ0pIcFA7V1Ja8jM9Wwy0dxMw3n9azKIf7sA6Xi
54MnJiFxyKkI8AlqwBbQ07/3JLsOmm/jFj+NFtuJflNhxnDlV5aAcfCEyF2jBlzu
zMHho/1xsuyT5jJhOI/bMz1LcbzMWx+1zCDhT5rYvEUIVG+DzdflOjUuyw6hfa2m
n39rK+v65RvbyZzNmy8qkRZfOrY1lXtwJRdjqkV0Luw=
`protect END_PROTECTED
