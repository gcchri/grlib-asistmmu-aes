`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jTJtbyCDK5k9ZHwblUKLP1Iu0YoODTnhXKtlelqw+S/A63ixZeOjkczvGh4WDsao
mvYq2pYhR2Fl9C+Eq5sgAEsnZ8lcgg3PVPXJM59+iz8yKkw1IZ2Z14e742IsO0Bt
MUMB+zVSWUh+1Td5LzHddK/6fQtknuAqdsGVmie0OqKejjsgVYxWANVrL80YIYOB
P/GhhrKP4ndNB/OcymxB5oY/Wj3Hz2SocDQ2G2zeXqE6e7jmrORpfU/tLoq3ih5x
g64NPcuifhlsyiLFWL+Dhg==
`protect END_PROTECTED
