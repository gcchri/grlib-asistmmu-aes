`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qNqofilRdapsVNK+4bfP7zFJqDFTP5J1C6GqBmfFOujK5iJvhDIw+XMbWuu/2j17
LwWpIylXGJJIPcAtDvwR1SDSEFtjxJuI8BqaWDu5/Yo2eDUF8nU1QJ+ojQK+M9ED
vU9Y+4TQFYlVxSizM57p0jfdM1IJtssliYoAwKlloXT63uHrD+YyafBEnuZDmHzw
t3ES1Mj3PwAc+v4d0yI77BSKSOeW9+ZW9SZPDkerPSb99OlBbQ/pPuMY4oVQM1fw
WTGbyVUD8ZNBsrZZ8cngRx66Glg9n510esPdT0D6tbwgueSddqesSfl2PJjilYV3
mpn1umb5jPCr5s+raG0suRumvBmTK8Db//pLkxVbQwyrAhW4nVB8i7UWMWlAQ3P0
irLJ++fklhfyPhYW+N6usuqdiCTvTlYGQQK8fMXQKUvj7shZ1g0eDcnDPDVUJ50W
qfRGHwkPj/G/NhVGd2ZTssojMpa/4T78gEk67355XFQb166DUBkTohI2hqQzZCTm
kGuAYelW4fwPXICIlo0rXJUj6eQAQS2ilHTV5bcyBFgN1m4U+5lYPeBR+VB9P5Is
6DPlI+Fq6+lI2d0D8wWNpmMKM7XA1Biqqp1mkvRlx4cM4pehSHBjEDDHMG9bulpz
8KdgA6/4jryQ5Rk7+84JIePMT6mR/TTPYsC/U3HA58HbEcKflMUHftn9sRglqikQ
Pvy79cGYdDHlwiabcl+dIZm8DKkbhyMUnZIBJVrxeIhfAjxrxXqVeb50/zSl+Q8I
s96tH7wgiCnZUilcKrqgzrRocHP5zpSLzeornI28K8yplAr9PAKbin+PNDYrKrwb
0OX2F2j5TyphlgpyrHnnNisXqK9H1nYL6vbezI9dWtbg+Y4DACLU2fcrtChdJVw8
z4zOxaEpW9TLxawMQMs0/KWhrRaOHG1duOyYvVSnz9iyOMskG9OnkoKjYvVtSb95
TJXydrXiqlxF33OR1w7VSFhj/QR6hZE6X4SAmf2Z5mDewH06jR9WdYateKi9P0iq
Ac/q1Vp9MHa5mbJvUWGNZ1UyT1tO1C2wQvNgS8CSUnslFwhchSJLzu2j6nhpw95v
CVxmTKsxzlhLTA4pskvQGM4LfRu0P+QVwtw5EnO2c7TDhg0GEXyqbKQAW7nwduhe
lX3k9W6YUJwCA0Se4mYRWs5KExUArTyi11MELgEkMBwgqpwM1t08u5pFlZyYK6j3
0F5C5NB424jbgHcTHwqR5q6qlC0xBzg9VbUo9A5oatMkOXuiy4RznhMII0KLDmmA
y9vnHFQaDamvXmEISd0muppWafIlRZNx8TXFZDVlfircEb9FG0fPqTkAYtYVf+PR
WaJW23X6OIW5O1X8KMHw7JVlzsZ9N8dgbjNADefn22lmRYugJVLuhDjsaPyQiaHF
f5dG7WGDvyE1eEhXiT39k4ux36pc/lzq8IJ/nfFhtHMHEndveLebkWyKB5ubqhkf
iWb2eSjiXEB+6ULNXR8MR9gGZv0egodI0jGoTM6SIQBhCyN0JYjIYOocRuyZE8RN
p21XLjqXASSehssuckwrAlN7HqCJ3KSqOrecegi1uI0BC476E2OPvAKsruZ2YsUL
pzFnCGslkw1n572CV5pYnOngsm47tL3Ep1Lv37qOcWC7/pNJOQKh1CwQF8mmY8/N
arFHlq7KC8dWep2qN6AYGKMpfBYI4ixxISaJ3grN8QyXUJcSTgSy5TZrZYFPpSOk
pGkf/saNdxtB+JU0zw4nWnrO2LvTiUFfKl9v1OPdWshSZIg+nPO0j0/f/Sz7RRSO
5O5+h3AAzjolRzcb7M+UhsXNa0xry43r26TzIvKekuiP0/96gQo70WRCBIrUzjiP
tPT3PZ4gpfJrj1YSR8LZHVRxUeQg4hZa6n3OhP8PXQBG6OqxiWLIpMq6PCv//NYc
tYcV+2SVpk2zI8SR5xWUgHAvGN8YQmyp389tGAiph3GgX9jEv0Rj1qyKQmviPedd
aF4ui16+2owbBErYy1zQwaikbog5zVv9HKh/8fyt9Hml7QvfSwgymXfSxWGrFsav
hIkKYv+aag//GTEJXyUVEU2WEiDQxEFJmgvm2k+XnL07ygZIhpCioRCSKGWLDgwS
2T/+lZE9PTMinpMf7B1slaP6iPvQv4IaE4PzkgdHObCnHUOrtx3bWgB7WieVR1g7
3VLw4p73t1aQReqqdtQL/InzQDDBiP6cuy4YeLTkDbCVtwc40iApuwBEY5hcVFEI
DA9hdGvfNGj4YiCh2V2q+g2nhyYm8No46FAPrfo4WUGIfUutuN4JxcPLidlKujSi
mqY/jkJEfglxt4QqAbyjTj/zhbxLVFNgnDZwDaDWdiZuWdI0aAmb7gS7hJ8DlhyA
NhiCsmmFTLhPViyGKLvQxLJNVy5c21COEdHaU66f4u4dRQ+872UDQDb8hUYQVDhE
GNjHx9m4ByLi1Ifufm9HiM0QjpeLsmozahk+55f6JL1cSFuHyctB5UC184lQnpXd
AKPv66iuQ4X2uTB/ZvNSkDbju0sMtLh4jsGhcRGOF7S9P/ky9rKtSZL6IRFnCBxe
rWO2653ONWEGDPy1oJ5YwrPqAI7WXDXpthWuDJ4hfVc+2mOcmA4ryBtxlaVBHLpK
Taeg8bcjT9F/P/GlB0U3rQ3tnKqBmx00h7o5/n8KXR7rz24cubW1+CjCOGElMcoH
vgX6+KfK91Q1NeM0mjX+DQOiWVmLwwSw2Fgr+G/svmaJbGw3/S9ergFMpmRFtC3M
ibAb5fv32lnyreFGYPA/RaMDb1eD6cTdr7TPdo8UYiGVxlL+3i+Zoo+qLy7Hw3Zw
u2E3BQj/CbECZDMHdbqH4f6L9XoKkfylJMwpdREcF8iDGkPesfiVWHmnA/1DdLcU
c3zxUS3ft3ofVXoDP6MBcH/A0QDQOm712rBDXuoIf33c8pBQsVZORSWESHKgOqqj
qWFB6uGLPaeJunUq1oIXi2/n7oXQXgHyheLLrKx8QbtbXaPuGWqNFwyYL8EcmKvz
gq2MNbrb1zlPDD2kf9WkhjZap57Uak7Aiis5jbg846KECbsdDbtCRVN/tiJ7aRpq
mSlQ7wzgRfs3jv053Ft/pgKl1mgaYDBFonfWfmqDiFkxr/bvjSSq0/EqE1cAifcW
I11BIW8w5iZ58nW3Io2LNquzwE9aXyav5/QBjaHy/limxaA/RovXSokxjg0bXZz6
CEVrfaZQCcyCLA9f2OPzQXslWEKWk+9BbIMk88xoSHRx34nOMm8FV6QsS5Fc2PHv
`protect END_PROTECTED
