`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UwaetmN6aTq96dfYPz4HZgDOsK0cnaGs8N71kPeVVxOsaIFG2Eu3OggoBkN/imKe
Je1LdQs5QqKmZlHzVqeJg6rQ9lIkZhgMkxsw0t9ShMcKlGG259sHbPcVgbIKClMK
lSIcrKb2ovWkAHdEZ7TwrHme9tpGaTPgAqMLe9k4/ZZRrue6bIjAijlSZz8nhI3b
ZdyU/SqqSLf+EGBsT493wpXxkgppZW6bn+UzZc6NfvGVhWHILI9uSvB84upcFHOk
U3gn8984Ul2o2gQ+9WtN/ueM7YzXExqVWFkFSPzycLuR5Z95DeZ6dwKir4M2vZ5q
MVkw0rKqNOvDBgGNCdxqA3MQifQTO0T9gzAdcOrn4s3xYJsdC3kBxWoCaj36YKwY
mqSYIWryzkkoc3nfHSc4ma/md1nOmSyrh7oSFzYi28WWdUYuFl4f12kbpYT4TZxm
5UqTa8lz56Fy+s0fS7QPBeASLvObIPDkYYij7lQPwZO3mi4lzR5CrizYGrhc0iD9
LmxlxLJmY1ZFMeCJ/gzobWdbbqXI2mGevGesdG2YoRIWjiZK21pe79I3D9oYMYpy
Scltvj2j7rZR/TrPItYKxknCZ5r2ULuscXeDs6hFuG4xmH3sMmZ91w9fIk2t33dz
JkFvnZf96LStUrKXuelOEbkl/S9b4w66NBemTGogL0I0c2DFyp2N3bTPrHLhs9cD
7XlKk+1zpyaQ2NBHsasfBnlBTl68YbhPKE4jAUx2A7+JckqMDhiCHTqNJ7mOgXIw
6oDz+2xLTDTPb4v+Qn6Mu8p448Qu7ReN3roKzDYZ8MFHWhAzuv9dNb+OCF3G43N5
/UIwqs8mOEESGgzBxp/XnPRSWNhaXvwKQoLqCEBA6VFBjQvhbIGkWeUNTk8mrDnh
mV6SihfUC0BUcwUYdoXP8pl7i2KNxcv93uoP/5GMP+saxo0ThlY5naFZv52Q134Z
/keLxLzHcnzebNCngcu1iX2XNcR552YteQzcGiZ5IE+EqZYI+/vKc/nNfk/SBDsc
VDO8Sv+3BY5pdPYDEwwQ92HLP3SQ6WE8FSUBNiVDjxTVNeiMM6w9XzcugbDU76G4
m1bCk1KOLys/kJy8TfOC4N27xAIw6PzqhQbEbuJu126I7hULgf2nRZGOsv/BcKL0
L7ksvlOtz6T52pRVdi2h5WWSfjvvOYVmlNpIhX2mfn0D6MBFaa2VV5kVBniYTexB
bZ+4Jjk5ji96PSn1M+Yqt3XDy2ZlCVvKm1PuuAzlO4fdOW/oB2mRSk0mWCQXB4s+
`protect END_PROTECTED
