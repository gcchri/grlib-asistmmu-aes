`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y/isVB8izhhJ9qofVYbtwxRZYLRE1ie4yuJcD2HzgFl1ZPJdzVSfYvw9wKbN40zw
csj6eX/qdB4A1MYrHJkzgGGPyL8U+GsUu+vEDuhpjBhueIdIwqvEFwfHQAjVrZQo
nqGFkGdxAWQWRIKuMSi5aWx9Wc82rbwAXKA1FBlV1GQnIDeM6eKsW0lwiJ2Ja/sO
1KEdX64kxT3De7omyjeF57fvxqUkMZG2xcoy7qYG6RdZtBwRVKtHWhuLU0YD/3SF
GgTIY/oZsm1Xanmg8aUKKX2wV5Asy3FQU6bPHOvwUDICF2dmmMQ/pZxyV5XGF3VQ
gmtaVdjKbtYkCDjeP6tOL74JATL65ERZJZClBlXfnfqbTvlyaiX8/sLMVX81K/RN
/eUzjbbtLTLlu+rkw38giTQE9lwyG6movNd96dwcUUqC7d1JC4S+xoIFSEZMMbdC
uYn2VB97MUWY992WOX5agv8My193P9mgeHjjzFsmvk4bzSzjaUCWZYJNliNAc60r
BSF3w8nobR6o+8A/afj9lZwd4xkE+Nieij4Gmlr+PPN+cw+Vq7VBifQcMqGkvVb3
bpFd4lpOZMvLxBk2josvlF4yWbiYhSZQtG7mfvPHvlw=
`protect END_PROTECTED
