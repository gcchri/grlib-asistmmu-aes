`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Bu9EkHxeiCICuaPrwMBKjCa2gxCk8da0xjU9cFy+z1+TcnCV/cj8DxB/gfDccpk
9Rxynxyj+6i8wL3QeBS5x4BV1nNGU1SDxwhc8qmnBemHzMZj6A4XGMYXOemSbAtG
7LwWT4q9Lq6vOXRWuZqVMN9cjD1AJxAAlC3rCBJQ3D6SYplww1xkBdmoSgHIHRJf
hZ1lepTJggPHr1Ti3XDpt3ukNCoQ1cCGfIOwBeQENHqVwWC0mIdmWNQSuYdZh/FN
`protect END_PROTECTED
