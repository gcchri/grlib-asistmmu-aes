`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nRDZ+XMXJiXP+e3BIoP/p0MzfJTttlisNktNaY5ZW/HXoardBXqHRonZ8HGssxAB
HdxLklSYVjOdZblCkCen1jIewGa/o3cH7vy0A1rZxy5KXu1E1r3XgjnRp9PJxhHq
BGJj5XGvkCsWSIYLm5Vj4hwYSoDYiB0GGfB9CO509TtwTLbK6ygPd9vMNcO8bsQy
HYECLXQPma+H+QDunRvPn2BQE0q2pXl3TYDhKwa7GJLYG9/IQfMBb76cZDJLHCmh
ilTdBPS1kY1u499MJ1L5OwzV+gXsW6RgMjTcpCs22MGo/OyOgRZOVufJX9UZflzx
u1giKiJ7UK/rQz3aLYGEW/4Zir58k26Q7AVXwuVYhKs=
`protect END_PROTECTED
