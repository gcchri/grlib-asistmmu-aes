`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vIXnEzJVI1OrRRlNS56OjLniLCzNy8Xrp/qjYejHwc7xLvSZM3k8U/3ZE8I/CaUV
vHfb71YfHIwD8urJssiUsxmAXNyqqhUQa1l9Z2dXuN0g5/rMqIBT5OFgGbkFMPa9
19410QtmZaMRje0p4lAMtGb4+SUKeMS+mtT15pgLtoUl3PE7wRH99jz07ww6cxck
3P/dn79MRjToRvHsDY+1803Bf2T2NCCIGq6Bu+f8oGEBTXtCQI3r1so8wDuPzoq/
SFnlEus41qbYD4lyjukxmQP+yElQEynC0qaxHV1LuPh9R3dlFEA2EHGildBzzvWK
4mlxp+Wri2PAGRM3heiF7OjR1ujjJ4T7jJxlHlAloG6hKp4Y8Q5Hz9fn9EkyxRsq
kBiiBM+Z3gex1Gx9/V3FRQ==
`protect END_PROTECTED
