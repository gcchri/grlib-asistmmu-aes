`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I6qpXI/ScmLLnib3UqnaHzQgpFViSZRaskKm1HAKbo1b3u5UTYZEwX/mlLecU3ma
YOReQM+nwMgFwgUakAM1zYmxU8qbYvzr+4C9+GrzkZ5yP/2jUDFsyGrtXlMAzDn2
nzoX9PlLsHfB0Wudcc3FFS/mslUHl6otFgGajtXGm7FwO0fauscljKqFcGiGVyOm
biEOu8gHXdGa8BeNkLqSAzogDrvjM3Yk6/Mi2R8ZC53dDUA//xAOD4hDuY228Jxv
szH0N+gQpxgYTHn4I60G5saQnKvgbSeMh6dNlK5I/JM2WDDFwWwZQDNlShRaKwh+
sajABxCt5DXNBLwwHtZnzY8ZZaw0h3ACUO9z+l4x/LzE2+MiHs0gORFkHs7NIwAN
z3XOkBGowihKW+CIhJmApaH6V97Tp3Y9Q/7pUqHPi3jBnuSGx/C+yl6F1663ODBr
/kbL5m32397AfCLmBeLhIOGtV+/gBNR2VIHOdyZkPyOavaFbUIrdAkjJWjbsOThA
RCT5WHsyRzy6We2uIi59b22C8Qz8qOiwnhkADDt/nRy0CTdNTCov+oqH93smsSRY
bGftsEMeW3cxWxbAv9+D5skiJGpUIfX2Mkk3klRFOiQyuxTrrb80tihszYwv+QcG
rvLf4oyuWC3sQq9Xn8J743DNKG67IhTqrfl2yk+tSRrUvxTyp9t6TOoe+dyddAk5
YVrl86V/sxvWjTV0lPhHhrXWWwQB1ZyiDY6jCdpO4sG4QkjuqrwZvSGWRhkeU+tj
hI5aet4W3zHZ16DhX3iw4uaq/YGVVIGpiiNHWFBMfbiIV+gCKCW9X3X8t4UMwzYC
uOS6bW1h/d8YLoNfV8kKJKGZl56MBc6a7ZFC18xQ13G7Zd6pTaoETLVmoGiif1Lv
m3cXj/L7b0+e7aRfX8MlTtQDvwVq7p6V+DSbiu92cG6iLmRX0xHlkPk9g6yueUQC
VlNz5zjIyE+e0HwXZlxVjF+fpg51lbTFiMEkFL28tZyGnFgy4Pew/fXHC752xFek
W0un9lzSCllpX0AZ3A1anTZt9khtnd8oK5uVFL0DL+Wl5QTiqkNB5ni+O7PB33c5
ZfMS+v9BmfwDIm2d+wsUfY1CSSZCdP+tBS+JfbVP8NmWNYhkfKHPj/1GJrRfPI3Z
sWXGiPyQxK0FIMPf5ZCjXPcNEOah6QrsONUmPPvhvVThdpfDFJWp2hkrv8iA1/cG
uxRAdZY9cqUZYMNbZb9+S7qKQ/5jHlRzxYj6FubWsSRCrhs780X27ToINSzXr1nd
hDeNzcyC5a0Gl/2g/ERoR6v5gspt/W7uNw0pkrRH8/iW5d/s4P8UpAy87qsuwMie
/4a//Q1CLje+PZw3EFCzaQ==
`protect END_PROTECTED
