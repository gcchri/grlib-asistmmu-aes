`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3TW8m+ldoGlJi2xEfLiV460pGiPY5/MbYTZcbiiOJeXqkkOgxd6F4Z6hc3Vu7MPZ
BR0YkHLYsMfrv/S8W8lRz6s5979+DPuJ07ed0FdbIhGX3zK4pHlTwc1JrFcANp9D
ZBPxuao0bx47b0/rjPRlaXJ7lca/SZENBqrvTntOogl9diz1RL+Wg2EE9OkvjEFR
cbO08rCPhZgvFzJ1i6eeiqbVphuSq6mU7aongZ7vVf6XCbK0F0qy9gUCgmMrI0wD
xCZHVtluxqNes/7p8ph419ELZi8AQphnWEUOe6c02ihUpKQ9zAte6Iat7+NitCee
SjFq+s2WGKACwrGBN52DjSAytwKLse2roerfSWpt5SiiM68E/tUfVlhSpchE3jPj
ZojcLOs4EQu5Uy6OMA4pUSaKMBJ59tk8EmbLJLCkM4LVNYUvYV/yYS0wVLYocnot
YCfAxyXAxvqD/zmjYhx/eFXrwZ+3IpCrrLy5oL9JzAq9rA5P89tRrnnxyBKFbeLm
u0JkW9X5t/aSBrw7SXzU0LenPI1Q0uI1ZcrlHxlDdwax2odKGP6yoQQCA4ZrLawV
d6O87aYp98YCDLqs6UJHFwlAunE7f3Ccn6mKfKYn/hHhoMfFQt4RhuDnH/V2wFkz
2ZiW6/sKTOqP82UKfsx/1YlUIGupvFRByC62q+mFVzUGz1/7EA7JaP8jHEskAjhD
TF81qxfAG0DQbC4rYDDCCzpoP7CT77XZW6709xrT5h25YqWZrQyqlsQN+p2r/gcx
65/QjiM31ZWS4qsR0C9R7bGPM/e605CnDIlA71e2wPgEZXa0g6EzGhZo7G8paDT+
4SG7lqTfBDA87gCCHAuOm2PLxsBt2OE/bEJNK3XIRlXGAw0+/8pKxXsomylTp4jW
et95B6Q5QhuL+MZOUNaR1YtwzI+ZFmzj9tUL1oHjyyABgrWM/rjGDm7SGLV+3HBP
x2TQ8NPqQdpu6ka5OUy1sUifQdd5YZAcJCSp1lW+u0EMHFs9ClJjziqRlI0Oto0z
wAZj9XLy7OrkMByHS3Wc/GUNVZFVclIVkR6xxbstZ61amSJfj4L6QFTaE2WmvpJX
LRipcPjVRPXLto/I+laR6ixZ5M3eigwAlQym4L/pawvmlw2GjDAF/xLE2k5PFDby
YSOU7sUK7obJv4wf6Pc+st9B9D70L84GCM3TWr8lqpZ97WHam8u6X1rSD2ABjWrk
HNo4K+Xg1Pq5L8gAgRg8rYE9/WG+zPxkZrsxAvJZ86CXXfs4bVz9WNb83ui0npNY
`protect END_PROTECTED
