`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Db7XMSXjIriqGnZm+QO8INFjFwafAz2iVRqUYpb6WL564JKtTwADHh+sSLFdTWhN
L6lRPT+V6x02m1B1EleAqPK2HnyvlSN38cMTO7p2MBnZHqGVDBVBNLQFWBi+RNaH
EiMDMuhjQipDvDK9oFst3gP5aQgdXUZ25mpz4q786l2p4qLjfrFggDO3P/3Tw+z4
CVchW64l7D+KUXJUiTWh0GIpVsTCozBz8riPPX+lrJK+rzBosr2qfMvddvJMwwew
+sGrgsE1iMmeDaUJGwLejrNRKDT7jjBybCcGNKIEc0+4O4oZKuTW4BEodMQIj9cx
eWDLfy+QohTsBdtOOZjHqSbAiUFaav1GuuoB7H/LRVC6qnzpBzN04oWqBdht0VR0
`protect END_PROTECTED
