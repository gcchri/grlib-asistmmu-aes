`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
thTM4tIUGxciveNzwrUhkJPt0gNOZ0Ix8pzH5P8vyGJTlIOwqQaw8KPuFSv6KHGW
Pk8XiDmNd6hjreTDJ1ZdhK1KcdaIVTiO4USWrmgy7JcNJhPUUKh+/NvBgxRJYIgF
FdBfojyO8AClfZi1FB+U5/gmgzMDDq0JB9mKpiIQ+TzjN4SVz0EZio/QPeCQYfgh
dizE54JezYhN0dOIIoCeBJ93d+eVAu/KFzkzW+QD22gSkO1+XUQ9EwYwc1HRmnGL
cUTDRIV3gTKskpO3Eq7+NGw+8EQU2pZH32MISFmp5oqPXRdioayrjRpqaGwlumQR
A1ot915A9P3jzFyFHCkuNZrJBx5fqAmZdUUonDW2N/UXoDRqHKhk0IPMQ7aAzCWI
T9m3O9Ynu3QnrLuS88GdiOM+OVTuNXQUShn3y0m/8Jpp76wT3KF0sybSQLy1sAxK
oZBbbd7cXsufJdSyXMy9fH2+RWAQ4IsSuwih6BcDJd5+9RPLFcYSQLqJ5BDc+cg/
504yx+QxS7JlHydOt8AsGmsp84WeK2ujv4YJ+KJY0TsEq+STHalj9tlPTkRgtenL
`protect END_PROTECTED
