`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4jW4FPQgBW6VXZGubIladH/SauNgq09ul8Wt56lYEz5JAg6K3kjLop11BwxYeMqe
PC74/J1WBdNyOHV5iV5X6XlljU86CDnXIueHRrBmNbvwWVBrfw5mc1+5sBXpfAav
B6XwTN1UBCRt3IQQMx1LfDulmslEtPdeZRswrdgu8PyD8eoJlerP+J+mquPT+hwI
+zLphUVq1nQOLlPDakWQf8GwbBWDmfLHomX69iJmQ539u25dPCSQ3S8OmYny20V9
FwE8nUnBXuBELXKmkIThKJzkbVWo6Sbvvc85KBKKcowcNzm35OiWKtI6ta0zxzoQ
/Dhj2VkCOubHtn1BGJcQjodeg3ftE8pNo9uCehviS/1l4gElclbCIGhIs0V11sMK
`protect END_PROTECTED
