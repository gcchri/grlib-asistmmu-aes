`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ORLzGrjB57CJLSUKtSKXmk+o15QW2U+HsguAvo6XRyjfNdJ22aUVSrCAY7/mfaml
60D0MGuMDxXd9BMPJLGDk0jnEALppXIQN0sXHkVEsuvkrygbGBQ+NnXdizXjEUMr
p7U+Tc1T937mhN8hnb0d5ZdFq2hdLu9da8D2wof3zc3umT1j+gxOadUfeBtmlfH6
ecIaZf4NYt7I1+TydozP9lcqpw0sjYuKItoejlLX0Hexp1YeCocPSaPDG8PitfPi
CIRuung8q6nteBG3JoB3odIPJW9AGrx56NKH99RwJ3nrdztacsDr8zCqc3hJSj9d
FSxMU7Ph+UaE67I1AkMO0ydgsqsfw3SB8XwJodYIJpIBrDEoelhIPv/GuMcjTZ0b
AiLyWvpmLY5K9GkJa1dCkEt82vZVdDDxmx4SnLjnxAhxd+t5LgYYJDT/g3mltlR3
mGLyCAN3ykxNJ3tD6y/fCQyGA6JcFG+PLTw+O2kSsR/FqcdQayCDYHRFJefFaJ3h
ZHgCcuE0uQEKH5wAsY0aqlQeeRpr8ISYmjADDj84hg++cshuxe0M53BqrpkCxxaM
kmxeveMBSL4eP8C3gJiXTRgUlPS0rDGKd6rqeXnEacEAwKDXYGs3XqI1w1DP/5nM
oQ+TGFE6NWxUvov8TBtfXMM66EPZ6wwlEexIEH7ajjXq0agHFUKhnp3Osjnoyi5f
ltcAoVD3azPbwdSk/KQou/7TTfVwwrXKuXtBj50byNT3JGO+Y237j3pwsy00ktRe
hoDvEZXHovQHqG60rHtv+W4hokBe0VPaH4lfVWbBPfIHoOPARZSrVYIa4oKtDrMb
EuPruVbXWhtidmCxtqMWkFmtR4usnNMbgYGDXzm9Fme7NGDFW/HcBAKyvJ+t4Y2O
MTjykiGW/RSWA2X+cZFhckAfk5IZrvgbJm5IZeVjrDCFleqpTDGqszpt+aM6bvUL
9sGun7W6/fjgiy478jGaDiJQHf1+pGNhi+k7EXCA3D8nGMpgaT5EuGkzUgJB0OP7
qV9ka0YhFsvdeQpD513JJOJlk+KLzUUZeLsgj/aZkrod9P6LtQgp71DlpgnFQNNg
+6G8GhG7XuTpU56AYA5FtWDxbn8weUr98JnQcZ9m5988qyjcHUeAgciAXaIaOiVS
QAAtEi/lBg3959l7zyp8vfEdMPhKPlFKrlBlHRny04jugQas0JjucJj6QhnPzbvH
64t9qY5nQw7tcNl3zLWvmHzWWqM0dESbP0XDa8dp6Ddu9nGQJZwA5Njv5jneqT1M
tO5rv2dDUM/gXRRhn7TjVpUxBzu8SN3W1AYJci97oLWmwtcq1cwEWnFtGNhicnLa
QXX+wN3m3CF51zrZK82gi3XF2F7FMbaxH57D3siSbMB7dDMN9rtpdkxxnvWxx82U
PVj6yuvMVyM3u9eES89DZVTX0NY32GoNn68X6LcuezG2irzuqqySFuIR1+cVQEWA
QLzh8PBFDWC6m/z0cm6eCisv2wU+wJP2yjRbA2ARH5+jc29CvbKbjmC1NV7g9brP
DbltMgdOryQmU+pOIfkDIGbd3IXmMZKEL1JP2b5DadtPLXcavr+Sd0IROlO67yrm
SdBmsLqqLJFPcvbxysYazPzpR4zPtky250ZrXYflMKvkBIqyxg+SQp86JLKPH9l5
PlqAZGMU7S7eH5Pr1wf6geX0Kqf4j77o1Wod4/h6BFZG9ZBujRQ2SNCOWVDonqN3
yYMg1vzuIVGYKPkIGRQxjhxRZOG71SEg/PEA7j6nFOw=
`protect END_PROTECTED
