`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CBHCeDQwpPKAy07Uk3LDRhTToEDhjBvhwzrpdvFKvTtteApeHOHxs9Pz1eJRSmiC
KvMpxXYCuKJIwJYvyUvygh0iuaGmISnv4QuXjfQA7/cFW5k5jUSPjtuVJEmFhJhJ
SPH/nvNTZm+6VlkuyHXmGieubPD9CBI7NP7P880BVUceEz1Vk771WJEG2/r9YMpx
86/4xvF+jdKn7r7UMbqrUwrRrQcyyehc1yoJvvSmlWbQYYdcSjeFkSJXWRpeJySD
554biSQHby7BLOif1aVHmSpWhosQushDUPSfkjXDdZqDGby9ydIs1K6X4GNIW9+Y
WU1kI+YKRHlBIF/OOSn1lupiz/E2GezfKqr6BJoC+EAOvVgJ3tOxMdDCmnH1Nh6V
4bOUp+kX6llzHf8qUILnKLEqNJkoPNS19WDChZpAQW0=
`protect END_PROTECTED
