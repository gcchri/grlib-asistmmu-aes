`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ltAoJ9Xjbz9qf3++JWknXQSfaCUbf6PawoOMcdgMbJZjjNv/c2yckVSzL6WIObkB
KM877hQlYPhq8v0SQJxyS2dl2+IUu89LoJJtegI2UxrYRg4/XXuPvMo1jHaN3RNN
fMJkx+BWl5gtnbIPzYEwoHuT6Kek91eZLjADIkK6VKLBxN6tah4hr3vVGVd2OZcW
2/sWc6a/PeKB6YJnU9za0gsstpa0mAaI5z0/hb7fg3wcQoV/AuK12Ki+VEANvD7U
gJ8bL13kxEH6fR4y7k1kWRj180SfkgLcnmnaONrZp8WSHIdDrRZ51S1Xh1uxcPdu
3Md1ifBn7UPOoM+dIXvPjUj4cHseTBL1OAbiviQzal/D/CVi4xqCJOOVjhthPmmR
0VepWC/96br6/I6rQp5U/boKshXuWM7Q2KWt8oJpCDuevukc3IC8JCjFheeY71zA
Q4c/PbicmfKbNxmeMkMYMetz6jAViIuecmT9mYIGngrRGikSys86PuJ365u/kN4F
Y15SEBXEhNuRi+6wLlQvRIaWX8sSmxjUvzw7TB5jHB19h33Z0ZWWycPv6wV+PGX7
3pDeHIIvHhKG0gehpSVjkrNgwbxNXZNyBS5CSJ3BaGI3ynB4CP4bH6GFEJtjDbPG
dfWQnkpXM0totGK6ugmLDeDw13IQhJHt7FMiZIs9Tl0SsoqU6uCuvieonyNqfyxC
EK+Q/2JMU67A5Kn5THdWpryM3ZKe/EWJNOX0/O5KZL6CtIoZuDbLZfLA0PZ691FY
D4ZNRjX6Gf37BhX7Hl9m7JEo0VbZrNlZD4gp7SJfSCf8AaJCPN0rv03bOstIMFDW
3tibe0oVjz2LlHKxN5hj1yl2NVHR3lncFfLkxknQCWvLxXRAMY+USGSKPqdOLVak
sBVcRmQkRjylIgkvjt/NKpUw495mUOeRnBniB41L0MEo6vvwwLlY8/xud7uDvnH2
Q+ea0Phs422rERGK6gbL2IHa081dfRWbFgeeCuUcJXL6WK2Nn/tHd6BuR4Wn4f+W
E7g+GzOm0vSU0mZFkGF+yj07k3WHKheP+q7bMuOCrB8QLRvhs3jraj6rNMAlJhMz
1zxzqmzQjKTkjGUqT8qLOrFDNuk948vjf/GpIqmRliMQdN6Wtlau2qfa3YgweCgk
I9R1Q5dFBIrwqahcdbi3F46yFkrguUen+0/UpSAv6I0eJglRcEQYFmCfrZUUdpyc
jJ/fS3WzfsAtcY0Nx5iBsmKdx7B9FMtrUWZiR8gadspTqi9Jg4+EN6We0KeG/oEM
1rplxDn/GVgAEc9XrR22HlBEqBdIxqOPjBw3EbLXvXbVi/z94+A6g2VMOCGv11/s
Z0QbbIMTn7zXFuqEDk8J0C8YZ+rF0nw1YDHTKGKgcUpcRLenEgfSoCbj3l1ENVqk
sfvd/B+kM9dh963dx7HIORQVtTT1PGLwbAkYoyx46bFiEE5PuGoYFH09z0Imf8n1
Ow+eiPv1Nuteip5MhYyl3nTi/TY7/FgUpYYnqfiPhzEEXT09JrT+7u1CCgQhsFNj
xd/2JntsuMpewMbYaDb27JGRFf5FJ4vwNrOCx5ky2XPvuXEDG1juIkWOwEmSXj8m
STESalSlVdjcGtWFsWq3eV5qPtzPuh1BKmOmDLKtrHSw0Y993oOZ8ukSm71L16xp
utbpudWT2JKw4c06nTUzXzZfwFErNWchTVoWjn3XHiVug6qyYOjLEefGuMbiOiiz
WRBz3S3NBQnAaYK8+rOwk5hXQGaRxoUG6w4bArNvMJB67FDwnIxKCQ+osRcsoswi
PFAWOdtFgDPiZQa6Wae/i3Z58E2yGXXt/r/gWFiZ1YLL9bZto7XmL0nJE6JrCXsA
I9iSYqlFN7qTZ61YvHj6zx5ya1FaTZ1vyeOv83EIEKsfpTNri6wbfVn3CNvmzeJh
jbOqgaYaQUVd83vJedzLinwJa4ZeWSYGZBUFo3Nq0r1xLMzUTw+HjDlvKvwSAPpU
wpTeYkonP1ZrRWj4WjCyqCJKX+qkQLF6CnAfEugSrIXhfYNI8KE/HuTeEtyh2THE
Ep/rkunvHidPB6sNaV0mO+0lQ+22HPnhAfWJnRxFS0FSSw6a9FBOf2haCr3Wl+zy
TrhrF8KevFZodEOsCnBNoihYNPjLUmdzsJQy5SZpQkABxOvHyEaeXnE/jzBdSwWB
vtIE6DWNTvXXs7750wzpBQ3w+CFcITaNw2Nw1JJbN7gNU+OlcMNMsW35/Li7NvYt
JoWfb1UJwkIW84jV6jeyJjFPyMevabGZQT+ndhTGGApMIGw8RiEA8Vl8kr18vOmg
ykCfqmigICxCPPJBhR/N8eu3QnQuBJuZKTA73QF4TiO0w0IvAD7/Nzkax9brUXfh
3Ypitgen936DqbzPl3BSWbdMCrTtFMZir++OI85y9Vv0zlk5XqJsBluL9oULaf2J
/D1NMp+IilQf38JWtk0Yc5k9kfZfLNVmrqSH6ddnpqMDeikV1nYxQuM6Nfba2BBU
4tqdajtESS7DYUDA+5XskyEj7RYg7urm6c/K+uEc/AnUQBQef1rbPjpKzeRz2Za6
yz0Hb4Ujzr92Qw59El+KVGFD93e3srCYzuaB8DejFxmX3YIVELmV9xUgTrxTxduJ
3/gASypjeyGUJGF4zPMrCgVmzU8NeMJaBJ3giGeXrg9G7w6big85+FK3vnJZD6zS
d7Rae92xdSy11vYxBrpTFSI40Bh49VaLQpI5PV0Y7cJ1JfqbEz+vgK3vbguWhdTB
ie2eTj+mew8bye+NSYFoL2GGzLCZiHS1HEPYE9AJDz56fNO17mqN5LtqdoMzN3pz
pWWjJBFf8zSmnwQW+WNfZ05w0OfbfwK1Ex6kiCdZfg9YPJxBJ8wsnL6QMRE0rgOv
/SeNUPOo8ntrcPuErfDeuYYCcMjc9drHhxZpou+HpNzalIbcmEfW8OKaFhil7CF3
Chv55HbDGLIVix7V2AoXRLJ/setl2bSGIOJEKZqP1Up0y5X57jbFNXMGdlk3qBsS
IFKLKQ/9KzSsdmUU/UNL5aSnH6yieDd3fcZDIPC4Ovxvv83zaL3WlCLhwPcaPrIA
0eWSBFMFVl5zMHAyk3mrDV+/lYoq7Vbuf6GuzvedhaxYgYJk+xcOtrPLNHqbQGe1
HxU5lD0EGJGwhKmmedQZo9seRHoSrA2ykMuKEtnArBC7jWl1Mhr6ngvccL5u6js5
kkzOU9+b9n0Z/jv5rcHRxxPaRpV0F6c6uGunhWvTDZlAYmoFW2FH+9nlVu8YGQhb
RTp29Tj5ZxyDcPSUmWGkpuly6D9Dj5nB+RuI8+9OVFCup5TST6YVnTFtn5fvUyPz
QPdwcBTycR9AwEDmzrBAHCQiU4TwygcB8hmRymEDcX0wgqFJUjdHD8WYE2CcCOaQ
LlitgpDj23sotLW/o8RiotWGpWDKZ7AfEjzKUGY5I7Gyv3wIdJ+9Qwl9kvlT0iHp
jw/DMi9YjC65p6ZVAvNSPFgA19ycIpJ0Hk+vu0vaInlhTWlmq+jJIS8Bb+2dps4K
n57Q8N5h6RUyHYli52iPjVA2l7lIZL82eqGS1p5ma53McwVQkaXVONwXM3R0Giz8
EBLR5UQILvPG5DACtKkCEI7WZEOgxDqGar8CdHX9xdRIn33cXXtsdiP2nOQC8OXt
lx1d8/bhoioksWDqOsdm7ln2O1lq2fvLb9gyn4zjITe57y+6U7BQQAifGzxhh+0n
kbuKZt1I68DbUWBlTWoJbvtaSiyBuLB7gmH3RhHz4c42xMjpxkZGwA3JBUES2fVy
emxvL4eLbUMemoh6F+2IfjW2Lg3fI2XbsYgGUsOm0XyVi9+OURwih0eh6lL/ZxIV
SpXhJ7nhfnjEvBSTo9R+Rp0sBgIEnZsi/onbV1ho8H952wwZAhHG0uFgnUhj6TRG
f1jvNRiEkm0Yh+dQcK9awT++ZzyYWPGubN0RY+mKRIGbd7aqcVieKmy7GXHLSwOk
`protect END_PROTECTED
