`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aft9MO1us0PP8TwM5ofjSeIuXUkpslIS/qdgZnws3veFQLTCA12zgbt232pZKrI7
sBDemx6W1jDBlCUjYq+vjZUZ+XbTR6gLzwxU8Vj6vId9n/ZUnSgwpcu6iC9niVYJ
MmQu4Ujkwr8bOkv0bS7ydd0CcOJxDZ1/Yr2181EmElMFpTtU1Cg0dRBiY4vKXoIX
7+ZpGqFke/NrLFX0bSber4ZoEZxM3edxlYZL3nvJS69dm6GylifDhoW7ubNeRvUe
4NnWq5nLL5EABwc3o3BQuXHWIqUyg6i+YIVLx9lmP1GkHFYv0CEvm1IU/Lg58yW2
1HjeKnGyJFh5dFUcWBxIoKkAlun7eX6Fl1NM9+zhZtkqT3smt31t1fTMl8wTl2xK
GPvWKLuOgUA/WNIaHvw/QJx2sNaEvfPItHEOLDaJV3kO10nfEPZyyLeeK+xUYDH0
9sYTr1F7AFbwOck9kELanIVh0+0v7Fz44oYE/qNLBcqEVGaCcR0YECbxeAOyM9lm
Vm4dwfIaTTVOjfyZZcwBNQqqd1z1jZAUD9seHcu+hdxscA0uvARtIIytRQhL5fw1
VSIMU1N4OYHM9F1VOmzZQmHwamHfEMubU9z7Kl8MLq6DZmbYjRU9plt9K4WtfTa/
TtFHwy6dGZR6AqN9tL/1KsUXYRaU582N0pjC41V8bMsFCSDJzH6mJYSZibrnD+gi
YLtlWGRCUxFRUunJG2ywM/pgID3uCiOsM1RqJlUzikHeeAmwWXm2UCdWAxMlC9ax
PwPuA9cqahXccTlyONVpIfBdCHIhN0N5Fk9V+rwmKavVyrh03U0wsBbxxxcLSNCC
ZgHnCCW6u78uUp7iBsYqOlaE5KNfFbWCJMUIkFAXM7U7b+cerG2q0Wdc0GxDEB1g
6UZ8iLdjx2l9kC/zLqILPWprgWAM14w6mA8CqnOpx0RML1SoV6qmUgN0sLBpzDn4
dLfdXDGhXk/GXDHIrHRXe7tzOvXSrq3SBpw2HXjxPdF3Ih6NC+kbwWmgAy+xkyc0
mLksEcJhf2Cx8mQHeZV5knUcvGH576tpf4XrB/+ZtvEeTjyxhh0pT59l/xLGAPab
JHIW10aCcYSlT1ng1rMuKCXBkqj42RsQO50VLvp1WJOrnGSA2tdXrAUgLCDvhWXi
HoZSOUO0NLuUZ0sVeVR/YIICvdOXVSEmXG5d4Ar/CmbmRAhFhxrrdmUk6aQPRlYv
6uYRBP+bXl2njYXk6AljIiYbNCgVRLYO/rKVBNRC7ZrgdXnNSUFmVlVm7kSeD0Ws
`protect END_PROTECTED
