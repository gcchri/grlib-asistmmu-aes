`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QFIX3DozXanct3o5c5EYC8VglS6EjqVkwnb/t+DOUjOxj05Zgb3D78+3xRQfe0jk
fY8yXskQIt2MrZPuFeOtvC7IEDZw15W/btm6AbwBDA2zoLkpTvk3UQW+SoqPLDOf
4ZaTWnC3aWZcPwPir0hpQhpLBRxrXVEei7kAE3Bm5gxY7Nylo7PI2oktVEUjVF3f
p5Go1Gnr6ND84jjncrgd4UjEGZ7hkTGZtTH6ZNiy+CSZ0w6y+LaQtpxKb9+OKQb6
nxY0ShyUAcQbmB0keGssCQ==
`protect END_PROTECTED
