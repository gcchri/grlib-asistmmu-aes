`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pQgmAVxeMeN4OitFpvae0+3fMA69F4sjAbwioxSXhFkZV7eqDrt/eMi7XoCGaGGF
P5xURVfZiYaDVAIcyKsPqpycvMAyZ+0+9t7D+Ok2Or7o7b/eKf23OjzK1Xc3EyxC
kHsSvEHnN6WH7DiFHgyBNmAkqAlDC2LzDCSY0zfPeQPA8sm5aBKT7/mbRk814mno
21efm3K1hNA1P8Uq0DjFCwzqhdf4edDXIJ30yxRfKCf2nnDDLKhIvw8oynOo+8gz
14YWgDa7iF3Gq0jjWiBjfphfyLUN+aNnCE//FpItJTQ5vmNEyOmepxFptlMhCQe3
oziz3Q2onFTse5K9p2KpBDaFIs5ojfbtJbyIM9rsVFAgbKF19hZc3FQ2wncnahSI
vBraLzqFJs/oUxTkBX+tsLKewX05ubzRQeLLFyJiImZ0xJRATeHngompKaVOlYoC
zmTBb5LoimVTeygbpKauYW1epoksLcz3tAswEJjI0JVm3/iy6MXBGEdqh5CquLug
J/Uo3MzQF4qma1gQq/cLVU7kJT7yPn1XG1AEVdy+ms6pZxSfZgJhgecsxsICXAQk
j8PEqTJNUSQcdkCJh2l7wNIkmsQIk9pAhy5pCXKLnL5rJexbr6AIZnj2lI9YTCXa
2RByS/GnK9mEwwFHqwq3I0kJpChJvc813wzEIBj+DahALpWuAGWYkL4v6Ye4YfhI
gLRS+aPvsh1JWNEJTfLk/oO1jy20b7+C1CaEOqUnUlWP9CkR6BZdrJOC8EH4VEoW
nisKQanaHYB97xd+l6bhriiT5KiuGgIvIpnY3uEskRXJqg+cbk1hB0G+vrbP5woQ
Y9i0e673nTiEg6RzDOW0R0BfMHo3Hr5nvpQQ5zpz2M8XetmssQYnZb8BxcszgvED
ql9SAQBNg7kGsY3D7mdMwkSR08obDUsHSzgfrW30AeIeOYe1jHxF909+03dtxLq2
3qnBoMDZKJmun4DwY3vDt5AP3h1QftZqrYggCB2Aiadn/4G+UpQRPxFUS90n5EPm
ZAw4Sd4fHab00kfjgY07A3Spw/VwzPP+S6c0by+IAcuNFuDy2F5U6ueOXdVfWfZu
N/zGo97zJ6nmnLYwo3DGEpAryXd8clTUxA+I7tPlC/YW3heq7N4nu0x5JvVd5T7n
v6q+LspUHIYoRjJ+u92oVQvXR9nZG87BROGVrh1/3qjGR75kQpsjhD9cpSHTO2Qd
O7BmPr5nouihs9ePiG5kjJntnHIHKgE9qqdlJJd2FWVrGGJDfpzoaqyZiZO3PUBN
`protect END_PROTECTED
