`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NOJuE8kwpCOpXd6GcztswAHwZs0D5VvnMZAQH8a/PGeL+mh1Xbi7V0Q2GkZ+0VbZ
dGzD9fbIg1FfR+slXhYHEwNX+8ARDGi8RUmfrEOXqzBgmOEMezSgzrVhkQ1fJbDI
0rBMf8qGsLRgTElE+v4T70W/ye2QzSygM+RYUg985t58tU7bjT+V+FsZotsHp7hc
qyGyHsMPzDMDeO9//O6E0vuS92lmreUl0gSZ17Dis0Nfv0k5GGCNo1GXHhXA2eJT
OI83U1qHFqUJqaHoGGGePKba2Ly94bBmNI+GRbjuX+HkPKTaS6/2pHRCp/TxoLAO
`protect END_PROTECTED
