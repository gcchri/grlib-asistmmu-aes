`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AmH1O8UVGt/Hzc4y8W48PM1gU4runZBzYPvMeRYIeO/xDchYRGEx4JMOK4Ku/zfu
CWDBjzSrRBA0hHqUUvuQkcpGdeQNewO3AXXnqRcm9GUO3wktW+CuTc0aRDzj5qPS
l7obPQyz14b7aKKI9iRd8uJNoVxH6CHc+ha8KmXO/EUJ2OqHrkGPzQAw3gRWD31t
+VfBfGYuNlYkX0pu0tSxENfKFbYdGmbkzt+QIEubtqul/9b08fYmU4uc59ogfuWo
1ay5KpJqQZyasKL6ymVU4awIIb34+ABcvaRTmYRpR+3tFlgDlJpJ9ofCCfr4XE3y
tqfzrozi/ap9FEXEJPxlsbsbYSVcVPVgfv+ogo5X1lz+BoBGpHQjYZwx8l9+YyQc
6bhwsXjFa2WT6sZpA8nzcHDs0orqa3ky5e/ZYpGNA7T5gCQdOCBQnNBatG7E11wp
UH81PllHNoP88mUEBlNx8f3MZhf9ursC2psim4kP5gMdcpSy2gvs+wt+TmpNICjV
uga03Zwb+aeZ7dBhV5LVGA==
`protect END_PROTECTED
