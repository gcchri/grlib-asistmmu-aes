`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HdJmKgz+gMQG5od2RmpKUoOX0jm7nhvkF2KsIkVsL/cA7VYTaC07k9f1McpG6Rso
HmbhmTcXB4B5FNJkhcRmNtuu/w1Ir0XBb79JbQxS5/E1mR8TWTG4whqUo/W3ZH9P
16NEUNGtYLVUG7DpzCmIO3+PxCYmJy5p5SKRONgxhrpxKy+vtzwE4RqAzt/3odlz
bM8F6gf98tka5Gi2KwwX3lV6C/6X/l8VfEi8R13Ah7mA2F5NY0BV1/cln0BvY98Q
HEKh5YzxtOg2s0+t9TVRAXl8/p27r5s8N0E0W4hPJlQAi1qdi9lmeiAi4pRiPdGS
Z9rjf1DgWPl+ZFtNui23yPwKwKIPzpGlpPSmd+4eOeVDsFwP0o5ytq7fp9iz6bao
+MmMhGzqDIjr0Ue9ewzbChi/IF4ROu9e7CGIGY+Qe2gZW2K5sEI9FpY9WH3aal9h
BVkI6x7fqkEIWBdLwurJ9AWWM3okqimiwu8AoTOd8TrJjSMzzNhQMA5FJj2zuTV0
Q9BO3g1qVcm+33+SkmxcYZlSUCcxg3tFDktu8qi2qDo+Ap26yUG3ZBYvzDh2YnPl
edUtENMNX+hawK52X8fc9w==
`protect END_PROTECTED
