`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1J1BailyCBUd5l2Yb+PX5cG8p4SY6PESruoKHBw17G8TTRoKvesqVUpMqVNPujSZ
SD3NWqNNVs7g3LgeT/T/vkB42D8Ne14LisfKBvT/4H4XG8qBJgEuuMPjje1AYBV/
gmMRTdgbEK+HCDtlpTGhkNOYgAz2Trfv5/+sG4fFT85Y9TjRVzZKmEh9xoszrKJZ
7zlpPd7SuqDn/3aSHQAykOud8VGyBEZqUIyocVr4xWupLlWfxgzLAf6e44sMNIfj
oz3Od1Yiuc/yn1vB5U4Uv8jc94u8gOhcA+G+HbqHKbI9qD7A9cJ9lm+C0ZFbaIvz
+o+TAIImgi4KFDUsxSmm2A6OvnOUC+Bz+NYJIlT7eJz5C+iJqpiFruAr6BCafELZ
bpRBZxij7OGYimGdn9ijl7rwE5V/NUaU0Kae4wHBl9w3TuMlSOO+atMxsX2LLKrK
mEJQlXzHfVCv9mFKMXq0fY0iWXB0mxsSEN/Ikt1b6rk=
`protect END_PROTECTED
