`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cgn3ISnDupFxAej06BREJeqpitzjvjuGwlY05yfJ5+hrgO3Ha+A0QHNxCTIJLEsu
5/+BfAO3cvdplNq4sYrRkw+W6VhHu6MpZXyMuJ60EbXwNew4txprskSVpgyDA5Rh
Vzx75iKuUqcg8O+j0GpDaPjPZIDWDnGUHNPpRfqSzx7CeYIBQF9JJL/ImvFiYbps
JnJ8iBvJY9YF6T3DLF56egy7Dx/7VdYzNKpACRCV1BNemrf8AEybTNUzrWb7U0SD
tb9ymg2ZR9BVz7AkV6l/w/AI7my/Js6iMtQJHHzVzdUuBTFxd93I/ZrcBMlXz1+x
yzuAyzRkTcNWKOyjpJatUYpNVrlSBMLE2yLPaHTjk5zWElOlBzgx8N/8+oUkZVnp
2iS5BoPwyJBvVXD7o1StbME+gRuHKpubfnU3IRCyKvlJJ0aUa5PkY1EoLKrhMPiM
RNaP6TYSNPXQaLFXEF5aY7/w5LAZWBgRQIEtzfZim9xfXxHvXhpOwZUOSw2U5diR
SFnIsROHgMlk55t+S0HzSZTpVtc/Fo11CSFnrkKoi6OTrnKBX8hGl70R/O2spP8e
ZLsKKPJLvsysYpPp3oEoJEbBL/S7nu3LDtSdueszC8skpIgrg05thVQTdeiFFeBe
UoYGzmaF+/ggYlxl9ASoH8gDZMppPzmTE8McnUwwKSb+3MMziDmL6WlkHeBEVNsg
WSZYCUMWS9VfCTQpBXJYZBmjcMh9A2e2mnhKMFP5Ga8JFOqfbNWvaG54TBt54R4o
HN+FCXbX0ZuVQbcEVxLUTxh7o2PXBiQdpe2gaozbLOIzXEtct0bBBLUKaBQ7Dh4o
X5VGEUy4S32FusY30ZaYcDw5GQSSjlEnQVe+6bbRip+YKnEEgxo3+ot2whHOD0vD
liy5KkzV4AnEQUxybSLQEU+lVAVkV3Dh/Tjy01Azeoq/rM1F08GwbGGi/gG6tiun
pSbCqZfbFmcmSTOsgo2dQAoKY6qYyVwtJXeVcQ3Ts3apg1FCkAEgFNSUvy8OdvzG
fLzsA0MTehY7R5Nl+oPjuRDsj/NzeF8hiY04SH+DGHdrKDDS1JaGk/nyKuQSYA5l
gYPFYxVHnVQb3kKIQpvLpA==
`protect END_PROTECTED
