`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WbMHcFIVhCO5mXOffItWRIDAxtc2nG72Lp2OJidX0FEU0IXtnU3QMy3MkVoqSBIY
wGYSFarQjIZFEOOciBEaVbUMf6aHc9N9KdKVX9A2GxlOUsvruUi/kaCSXd1DalfY
DklWVhu1EssQti7JxoBlB15iRhQDp22kciV+bHBeuy4vMKJ0TYlUv2BhjQQ2z7Ol
uvF8kRiv6RqMLqWqRrAiVX4XrCg3FsAV5dPD8BGtHviu0v3d+fZboZydtl/9z9ko
me1yOC7V/2RABCtcSIe6T5fLzg8sBKCZWbhm7ms7fed9jXDJHylAo4LcihQT09/H
jHlMcFE96qzwyxe2QbnLgIDCFuAHK8VoJfZt7m53rhGyPesiuvVf1CZsPPPz3yAl
UzdqLgTNPWZq9xH2804rId3w1J3yZZVpcZJwX3COB/8=
`protect END_PROTECTED
