`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rorVFquXOlWV3ZYOX7t6f11LsunFmvSNJdLv7wQJIvdXSOJocJn8gcIkmrtDubyH
4WhCf8mJ4hD4rTguhOO+TtEpWeLmVBkSXlKekaYtf2mHcTa0wASwjGq7bcp5h5FC
HAEkwPhmOrMGNJ6iB7JYKoXjBkgwP5Z73N8588j0We2U3e7jfZrEE1rSKS51p5vU
y4RHUShok2kLkuTHiaiQQKZ6mvVKYjihHsOARVZMwCiRktrZZ/CvupG5BEnEB1W5
/A3L0eQ20KkoziueeuF1dJUkVM4vTU8cnZCxQ5RoSiD5P4wG77gjCv4PX5q37XTJ
rTPza6tYYf0Q4jclHvfinLE44fiZ0W9K3+70pgfFwgpro6XMBxFij86MTqRvIl3A
QCsZLmMr/4fy25E6Dm14CJvryn1gaU/Msm0/S3nGj1GlxwunT/AgFNAU5XvqAxe4
HFwITqbSXhEwuHAZ0dxv7cEBDzaYhLEB5gixvyLUUUIGWbzpR/ZU+jGMOmhM4r6W
s/dNmqwDAmD3xoNmct1rgQS9kWKODTMQkJLGVW5jexuqIYMqKoAy/EWyUXVQEnkN
il7bqSo2qltd3ODAsdTnJnGAiV6GRDQFS6gb/2f+eq9VAgWZWLw/PmWwNdf+UIai
NMbyxhmsJKvlHfJYoQGFKsgoqeLUsCH5OLtVNVL1dXPeibxGujy63VeXeWzAdHr8
EUHUWnpYsKQ4qAjByQ671cutB1s1h1w6wrTU0Drd8Qm2xo4Nyr0H3dgCiO2x1umG
sp4fe9dTxylks0Vop5EiyWVE3fn2QCD4i8iSOsCKJiw=
`protect END_PROTECTED
