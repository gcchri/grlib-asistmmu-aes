`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WxDTPOJWwV2snnIlPaT6E02nTDRmsP151mkJgtTjFFEyV1SId0EszU1RIUaXZ8JE
cHnH/NKXMW1Ue246NdZ4wyu9e5QS78TeUNnKGkvmNvGiU+oc5Bn4Z2t6WoXo2pMH
RdcV2qejRpfBAXmgemwRwnkbtnpOFSTFExP5ma7cFI42LCfCu9kLpXKYNsXPFSnw
bFrR/VrIh+PtXZAGcrb3GdeYakI1YgM/eeNMJy+oanIjMpqJsGkAZwhnkDtQiwBr
dZUl8sKrCnG06V8ZkUra9FgbKd1fh1WSpSMlPIOAvoeAoT5G+gAJhwQ7TIZeSjU4
XemAyNY+aGnOmSmsvjZervQYAF3KJ5Jmamb/fNyL+sCtJlPSCW7o/mGD4Y8cNKeP
krnflhI+qEU0lIu0kPOkEhDLy28Pbmwh8n/yKbmmIlFFkt5JB3sXrVTsrxNAe9k8
TylaIWf8vCddHKpOnxfADU2kZ1WAveELSO3lRtg5SGDlA+8l00CvA6s4foz5Oo/G
girraMXTTxUBFICzdFaePJtD7nEmlc7C/diK9LixWXpgFUKyV8D6XL4Ats4+MyFT
x/ilOqn/EvjXhfx+xzEcI+igj4M27DnGVOH9yOgaGjlhbcW/EkcBdHmGy0znQV58
OUxivRhsq5mnieL9yEArNsXhA7THncr33nrx7x6Qu0y0UL4rhto9abOyIWkHfrpZ
ZTQzLuW9GCmdrbWB4Cp7i/XBemcgQQi0E+yJbhAQsRMAH9hLOZFzJFPNYkFne9Ns
TQ16wzouGechiNVV60rnsDYQM/XhZ2FbT6xVpTxos4RMLGP7ySY/IWgMa1Lhj2kd
FsS5c7Om3Y7hrxxxUfoxsNQGs8GrXozfQrWesA/h7HFJeaEIFYqHIjKgEOa5SYF7
tO7S6Q8R2agPx65Y82M/qrFGjUFR2NL8J52tf+FTTWAJLbPD1TuVBpp/Gmpf7Byo
lXQdDoaupCQPHX7e0oQKjnJASunYLEcZl5qp2RDrvC8wUB0ow5W4c8Yly5+KQJRm
asDG6KREomKVz7NIZxe8HInnpXiZ+nqxLeDquKEOW4iS96U6A1bJN5DonazpVmaA
G8azDVOstO7ANdICqFTC9YqGQXh8GU+fOPOnHpRqJIcn88J6lejFVLo4KAzqBEzG
k/rmqi09GS5/gIovMbqApo/zIA3tfCrEPOjgcOMa4cfkUZlbF0Wh0hkPZpvO2LV9
iMQj/cEjs4veStITdcRxzIbB/Ps8JUm+g4LK93NzKWZU04sSB/RtxR5ndOaplvQS
yBGW6tFjheqYAqblTXmx8tKJhrAvmdzMc+XbrxKwjBO9maj8ZUjfsX8B4GfLWoqq
Mxe7YRgSInURaHegOgFzsS5bpAPYOotO4VmDpz0yQGqiKfcqLFYmX6cd4iazKcKd
5yHic8pOx8R+hU81ggWIP2xfQ/vnz3nfzhjK252iNiZ0hqja8ZufFldNL3UHK1Va
Bb/l/6+MS2FksV6G6TabDr5UzTq0k6G6njw+Mgh7QFvrN6RVJjFigqOmc749DS5G
s2IrzLyQ5vv73GrR3xpu+03AUstBCw10U0TMbanbJYInDKotjhW2duUzUh/nHiiF
S2tHCCgBZ7XaG5p5wwmQU2ARDo1oP0KO8enygkS6IDmz9y+AaNCCaqJ6Ut7Va44+
c43zGMS9wgUSl5GJ4IVk2QDgC0pC1Yoe0/o0Fc7+LjZOA4oMhq2+6NHmhXcyqPk2
hATwLp0ZFxQggUAtu1fxfAlTQU3BQWUNlvSYkHYOgAaly4wwRv2aEkPNJmVE6F6v
we2mMLBC58l4io1eroZC+3flmVe2d6hP9N+kDws82xRifRb3NTmuoKu8ta5Yji6a
Pc+Plje1H74uVI7btwjtf4jge+wlNbVDeNUD81Q7df4kDCla5jvbi26n0/L4NNp5
uatZB39yxnlUf19or0SO6hXsPlXny7UoOKaviY7X5vf2wwXKY/MCm0r0IAMzwzNw
UDyW/hJO4sbVNVEczqgmyCX8lsACac2HSJeNGXbsY6pjD5c4ktPgsurueVb3mKcl
pT5NB4o2rfzo0JEdLluGabpGgP0yWm0OkPIoZVgYHkiMt2jBkPyGGNfxTcEUGV0G
sNsQoYf/1tsaDAoFOvEc02B3sXs0v5lRVGifQJHKIPy9lgYfdJfaS25H80xaqX0j
bqNXWJ+Cpmnc1rcPf+v7N3Su0VtS36AdRN75SsUaOmyvNtbApq7z4R4U3R5zH0j/
niD978D3kxNfRrwwB65PAIexZOQm/lRGANb/xOUkrfbQZbWqcFL4jNRyCclqA/l/
SGULM0qw7lmxg7p++3aPR9kk5NSisQUxF9cMAlhaVmEnovmjBzzC4Nrnk9EIJc1r
Jts9ADxQaTQtm8qg84qlLJgB8bN4TF2seB8HM1bGW+B0MXsEUE4SEgLgo8ik/UAi
ClL6r78MpJ4bAbDXfkay85kNzSbf4a/mCuG3l10O8JmWKancRXlPkQjF9tnKy/wk
6w0LSSWJNbynI68FxUb97Nov7JJ832UxyqjOuulJmkxoDWU35ZOs7yOfS+JHPKmt
iBlCLRhjz7uy2F8XnJvCLaOijx3BVYtnMwh9We8m+8G5HcV4px5sT/8T8TQEDRwI
oZWfsjuU6zZGSNREIiVYXKseIs+3JqmDsc56vi63Ut0tiZrXPwQGp5vG5ZKQDhDA
Q79oCcpq3bRuvgFzhdsIZ43i1sDJ3V+YsPvLBZurL6AJnWUgrpNBA0f/g/QUPUKl
eTpymh2FqIsD2rbSP2sgwOgwVqDhHn7dbLit/e7QrjuhJO3kRsBAlhr9ndHJlve2
Q1HTNN7tJ2NF8uXo9AyFhJCeka7DnIt8KCjNfY5V7ivUf+SviJI1zoj+CPFYEBtS
bPnADKftUXn9n+97afALhH+WmipFV7hJLB3aU5gSzRZRNbtyXf6JNBvxEpvXhl9T
Su8+L0xjRHkJ7+4kqBA7T+T/xDyvONVZnQrkanas3RA/vRkSj6ooimZsOPteMd1f
epBcTZ4c+Z6QniN4hUou3Yp7TVgn4U4UmeGoGfIU5ZyXIPp58phuskgIgxvqWJOs
R3XT0IWN91QezXB6RTPH6hoAssMKvgVAcqNKseOAiHyBqkHdxxCjuGQn14ccMapG
c9Yp81KzuSC8UTYkNBUbM+vslAZflGgufpoIhFKE3VafablVkdWtcHfgEfkuIDB/
xLpqb19Tm6gHQHnDYHoGhf6OZUr94nOBsNPWYL1KQaYdDxr+vPWRxar3g+2k/1SB
gR8i6NshizpceCTgP7OZtgGJf2TszK5gpLvMi1Sazks0o67BUMc3abADa/CHqz0W
XOuOIN6YA/Y6c9f/fCeon4/8Fq29rBOlRZadovTHs2sRIRV1FN5hWVYzwcuYqph0
kzA6T8IkpuMUfHHIY3RtudAdlV5bxgTS8LRKxV1KE6sOZuIZHuMQkAZLnX9uHZPa
73RYQTbiYgMEErX7Eq7KGCZwrppB1kC5nwQ/giwqoPUFGOImJf52Y9UnWb+hwJz/
WBN5b5+oCv9n0fp2bwuXzDjPboa+b/MqQuJT58/T0mxNhFk0F+0ajeS/nVqbcvCk
qtIW+cD0l/4f7jI56CagWN/oHhvCilRisJkdiTtZqsap7+RMDSmxb81Pm+8j91Nq
qHblcnBOqXrNdWIdQz5yY5t5VKEYQrdKElTlyEY7R+oY0SYl01TcGLHsJFEZdDEA
d+A8BghFeHskX7ijIwLePq/GZdzNRwFDVHbg6A667TsORMUAnOuPNxAP+uI7USC9
QFmSBFT+B1ck3+hlajn9N0+NH/n9qijVBS+UdQsbO3G5v6nZKJm1BGR/q8RGRUTD
rmuZW7xzwvneyJBWJ92K7hZAsAHKLB78xonV8w/5xtqAX3JmInRrZ8od8PD4A7oc
7yhqCZNih2wsO5XSdk2qJlzjXsqfsPbew75koBWrD526xJP/qoeUqZ5vs0lxtiBz
NFGhxUmWfzgCo5VJ4pBeZBvNwny2L7qxiGR0gOFLgxFkqFfAoKpngNdqATOxPmbJ
naZumAw5Bhp+/45KDqugD4jfotS79Q1u+RluQO1wKF8LxbqQ0+wKxQdatjyhmFyE
Xffi8eA9+NDYdj9GZMZlCybZdq4C7C5JNNcntKgZ/EPlyhn0yBEfjS1A/Dzp4/ro
79wm0qk/IW1tCubovI6729rUXWjYbU5zHXj9Gf6NTaK/ZUdudOyXKM7fM7BdNM1R
TOkoCk28grq1ITudBqqY/OGayvNBsjg+cjt01SSiDtf7Ki0I/9/7vIzokNHqS8Wa
rR7nCfdLeCKWjnvCUB5VwyuNlF2PXxJ4nVHQWkfQLSA/leVtRyF4R5Ny0lGksPbM
wUMhRnDFt6VDTovb3Izko9OHwHARRMOQCQGUMV4WxpC1dkB73jFCubZO3Od4zF0+
LDHKq8IUcwCopR4lD4kySxwGV1xc6VnV7EG1oN6UyedBI2iMT/LIID9ZWQm3QMm2
n/HbgaOYyIuujtYanLxzRTZEl1qyrgz9xwknLc/55e/z6gXUH/ZWjPn5ywTKoGuF
CWdYcGcCrUS+bWJ9RlDA/dEqdpjXSbRYnKSvzA/QrgZ6Iup76QdMQ7Q6QbNT7PeW
2Qn8A3FfQtQ9b0ZxShNqVqx9z6KxekW5/0lmoAOykeGiDOvEZfGEFc1K/3ufE1ST
TRd7B5cKTdeb9iQ9eb6VpaYfgpNKvCFTz1J6eo0h7o3lSZzKRX+RSYFnQLP35d79
MxyLCtfCENSZtknxrQSioSIV9g6FVE8NB4scolUsOTJSAqcyAroXhjlxzmJTqraU
Dnbwc+U4VTwX4ZerO16oNgw+qrfc1jSdlKWPsM3Pi0DXGlnMvK/9g2TOM7QNF2Cw
bluTyBfBLSZFFc40X+5qLxIDKP4oFXe5aDrZFCd0YcVO+AfZXAkQffpUzBswPwp6
B1TgtslKRRtmogM7y0qXFrcj0Q56Gzmp6tBuTX/UdyJuphl6uzn60c+7Z1TeKyHn
2OSOmnqJ6rd36a6p6dZyNkfeYESi4lIWx4cNlYA6RKpiWa7xB2dCjF+ZgZhj0iWD
7+yjQASqQdBI6kPGfzH8zbT6CcciB/5FOgal7BMBK+7bIaPX4c4fiR4zpH4jjWKG
Bm7KbHa6kiauO4uMCs9xFLfoizTmym88BUQ388qstTatQdEGq/wvuEM77H+BCkKY
3b9AdFMMiQlx3C6CLLlEWACvM25/RbXczH6O6uvHRjuS3w9GP2+GXVkI+xixkTFg
sCWYmQzb2RyR1Qws6hQr+mr6FPZYopPZPgxnzWIsd8oNFWmQT/IEjUha8k257KMF
0r7EKiWEyhaRFgmj4Ahs/R/+YP/lLG8+XVsvqGSGZMoa3nNOPQsJLu+Mf01D8nRu
aJhrI4DzXcwu8CothO746EAwrcqrfdvxaJBo8eag0E4g9RUmmqZ0anRZ5Y0DQtZd
Ud4T6WmprBGxkDeuDJmOK/EdS5TjvSc0T7zEsAdZyybM9wP7u1JaCXiB66IGxZBr
obpo/6AU2VGrB+lgbu5YWreP0vG6g4L5VR0LL5wWZm7irAeqcnSXmQuKpxK5dSIL
pC3FXIBTLMdmdpxgt2g/+ntxpvu/JUrmXq/o1fkOoYxZ9SNN7Rx/qx9jTW0boKaB
nWseJuLaogMYVagR4yixuSikgklmc4t2Dh58fVW0c9iLlRazt5BE382QfjMHr8DB
`protect END_PROTECTED
