`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m7efhTkZHw9AyyGbP+7CYMzXFeROkyPlmdL81q2TlZ53AUGTXwAVzRFDwPMC7+R3
rNFalGAAZsu7iPiXx3S2Pauv3GVA/5cFLGvfKyLPgCxKjTs2WdoWaGzFfZTrormK
dIX07+R82Cj0OW0TCsqBRhYCOBO3l4SB0TPqaP/cwzt+1C24Qr9tzDXLB4Y4dt7h
w6Yr8V/KIeO/aTSSOo0jtK01nxiXQVWNrlWRY5HXrOsTCeGPOkGsexipAiLzwuqF
URZ+rDeszXk8ou960xLKC9nw1QyljE09Xiy4SoYRUG22Wy9KHSSpDu4Z/EcC8aZD
lHKWMyow1x2yk7fERxlD48kShJjlDpQUiOkwlNgYwlZbmQBGBxZnEL8Smidh3e+s
PRO3NHSJCf2zM57M3YGuSQ==
`protect END_PROTECTED
