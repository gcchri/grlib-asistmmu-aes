`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ukarfFybijVNfl3MPUl4G11I9E5UgDhlJuVaYqFD26SasFD1DDmrOWn3qfRHtghQ
kr0xQFRNHkV2rZOxDGVbqkIX984MKtS28pQBjqps02bFVGTNCDxMbgyNPWPSA1jQ
A/wXNmCBWNiD3So2byRvESc/ASK7GnlM2DXZOnWiZCngcMf9TtyPgLwuE1cQezS2
uYQ1IWR4rmufPSBRSEc0N2BzFNC2WShgnUpZ+9fk3V5yesn8tryda07rrg0lENPl
UvWo6TQM+AcN31T1C1L3KxegVd4x8zR7TQobU0AmGH6L50E7VTm0bWo8VEeV0tZN
bS8USfVMj+aRdQj+3s1jbbZ7eg6Q192j9wn8iWqWYus+H7PPUruUfII9Iu7wMfrr
3sgWCQ1K91c9z62eWVDeKyItzcfG1N0ZaC5mxwOUEkS61tTvd3J2HGq8MGXFjJPC
czDY7j92TLrp40GEzCGyFHlAQ7W12XeZmohMMbKcx++aHNvXHv3e5KRWQPDs8Dk0
80MslL+mg7upcexciMiNqz9ZedqXHYomJOq6ktB50M+TAMWUg2nP8ITIf9+b18/4
pu+vekNukTXHiwtuDD+HS+nyk+qGBKc93QESikCuZulq4wd/4mp8PY4gM4Bjn6D3
TuPDoLaA4wgIANpDohUul9K9EPKmgnmgtHpnz47hkMyYtSOdrHSFwwQBmgR5kI3k
T3yZYsWZd+1yhepBO+7tZO6fh3IJ4bR8GimapnDUihQ=
`protect END_PROTECTED
