`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JsdshmgagyyvnKBG1Y4MArCgyqngKUvfAZqyjMDq7XnRQDNGEN3Nk3l1hpZaLYrx
wxDAHyfVvhbhs6vpxOo0mjVfiWmaPSsZ3eVuGB3AYb9xP8yjGmiGVWU0AJsdPSey
qezeo1au2nPTZjdgcdxlI20o/jzw18sMvehMafN54AoKh7PLuOn30vwOMcyEoLrz
4y49jeHJzeDVIViTPNdWguwpphhuM5Luc84L5jIODiziLqlIzPiNAHkMRIfkTZBm
HHwR4QKO7z8deTm2f5vldZTPltUGYj6HhGWZPDz/sw2nfPap7LIS7vNE2VTROfS2
HSfnCV5DfZXzaQffkNasD68TfEmBoaqvKmEdjFHw88raAZQLNTHfoA2Uzb9ETvHN
C59ppMpvidwQkyCjBFKcoaEzpY2tmsqSxMMglaRc8bPR55Tv/RUYEJsr2UUO0hCM
g6z5mDC0dFDRKcdyPXnijkp060AAo9Ov49j6H3eDySVlLiitLS2JtD7Llvsc/sSR
5/IP43eQ1t5rmcgi1Nz0hxAEQSTWZxgNAv/JtbN3nIwcMWCH/jDMWeLg293HjDoN
xVUslBd35H/bhvt54s8ikfofeIVQoFLbJIjOoEDFq7DoEawf9DGXmNhijVCGFj+h
XSACuLNvGglZ5gWeMSJOee/6rzhBRtagj7Mmg9ETtSPOmsgTr8hDcgjDfOQykNh/
vpY0B0THJx17IOpy1N3rVMnxQFv1tWWMrzC7HQ0XaEr1xE0RcQLOc/UMm5uw5gnO
KlKfVbpNu1NRubRNpXBqyS99ftvD/TQFLC3El2Wm093LWcLgt31zBDVknLR5zPxG
c6Vn6DuHosVPjcxPTt5bPNHx0FbwBkxkDYHjzx4eN985AN6Qr4/hFns+8uBk+QA0
wtPAICcVGXoSD4NoRV7VYsq87NeYc8e8MJ44GPcJNKeLDF93J5kGBKclr48+nB3o
l9PAf3x2/wXvHJMOOlS3CVDzKsLpwGKzoUF35AGozGqEcnFgSsMJFvaMnmyTR3uO
N41K+cG7mlG1IhoLRW85Vlk6Tyxf7xR4ENs63CMBkEpRGu+fk3ebzS6dn+97pnsG
Mlgihrq7qbOhV/c4WMO8B43JjVtynXiH3X1isCbTqTL9ooNnLvfc32i2RfH9jg8x
XNT1WXydFsav5RC64sVeN18CArxI5+1WoNwbIf4XZDmPkXM/xBu6kxj30t7JDJ+f
u5WLXdpTbREJz1czLXgRtynsgrIWgPwZNezWDNHvhWyaPpjL+WywYfZmP6cB/Fe0
wYda0VBzQP0m3KAWZN6HVBSwBJHloxNwf9GZbPsWjinMBI5hNSj3FdhEyroa4MQK
+jgEnxUmRBifvR5Jxk/r5FqpTN0XbW+6Lnk/cff9oBIvLlQsuCEETNWGI1VPxRN+
KgZP7GFnYsmHjSGHKCoyPnRi4/zBmbSiBmzmGmRrWO909jl45w0fKhcvCZoRiAAi
Dqkm5Ido1F0fIpO/l4x/GK//rYc/nmFhR7AkrbKaSCVSK8ZYyDcWPw1P5FD5yzjt
qV/BHA5qmv4AN2t8fLryeiMdMnVF0/hUnr3SCxpILj5R9W1fKe1Honc0HdGv6J/p
x3okJMLa8E5MXnisCniGVJa6UX+2jzV81SpA9MnkIh5E7OyeLQ4uzhFzGeVTd5jc
0XOI3b8mq4F4HX+aPzBgZ0I8avS7yVbRvXngfpjCTJgRWkeWN4wggxOYgxljIiHL
YKSnU+IhRHjT4XQMeiv6rsr4WXZAf+hV+SKDcPY/SugaCDfVikmGV4pYMNO0xDNn
CvYEXP6N2G9nSCxLEJZxnPu2DhojK/hrrMnyNCrtzt0K9MtMrBLlfcucqet6aQ8g
FFspds3BA/l1Ywx31DZ4gToWK5YEXGqwHVlLufGE92LgOgbaSfNfq7N2BxLQdosF
7qPgfWp/6acjWV7VlOOYllOtRcSl5G1BrnB1zV/X8t3uDD6GooLLqGXcUT2ZJdap
52LNE7gSRN9y5/m+5D1GdfRuAyxQMn/eSnkLIZbtrwkvXkyPNLj/Ni8KDZlpDmil
umDHspeknbaqHCCx5U8ZAvxB52TdIEyREaLLOWAnJHiuLBrwoXusqPVZpfOLXrXJ
8h46NDTw2egemQJxw4dC/A==
`protect END_PROTECTED
