`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gJeLmXcpEQX8pBrJr/QyEGNgoMTbDx6nJQRplijxU91Fkemuycgo1OKgzQsEgMLM
xbEY48X/ivvdZZVQweE4E9ORK02HkXy1SI+0Hha1Y9IZsuscrI+F7tcAwrr+br+0
vghjXWlnsiJoh0OU36q/lGiBsUUetIEm4Xb0gJtBkXtwozNyjVKwJc7ThK0D2VpF
yjaRJJQHQR7OZP+t62C7ItyAtVxZJX2Z1Adw+RHBz8PRhAj1kqR0i7T+7knwjecH
FFrbUBh3ap/YIjTpdm9NV9Oh6DfN9WGqJLNk8Z+2zb++SLv0yuT5uG9sAsjUUc8d
JbLZVhD+haQQJ+TbmlAu8MNuUc7VEZsi8riXroSEbvp9OcKCWjW0Lja1xpP+uSgP
sviV7ZHGrLYBxXjoYV4CLIGyN3GHww51CwBy2SV1Y4PexOZrcJgfzKde6frZWkrK
aXLBhd/t9iq9vGDCyxxEYEC8EGMhgH10SkgvIytEDrX0JMDunLjw2qYYXQ1ZreEn
JBIQeUjEw45ffuQZrrPBNPCZwvQYO7ZtiV6Kqf7FIpK/LxzxQT+FDoR8vClyVHbQ
+bbpZX4UsZX05Hct33SM11b17MVOZUNxzU03WsSH5cncyF5bHphS5u0I3wdpk3pv
VhfrMVb3DG0VokSl87/6AEJYlNPbV0WF8MVjjQ/wyjKKbwvjDr2HocuQwkbLtGQc
xtu1M7P6tDkVnACXholXeJxQDW8ctJGSFbozQzsJEi1RNsk3B2QJZfYosRid1z8V
+FoUiQ+ngR6+OAcaoKnqbuW6xjWLETk3fG6TqYteEBG5RmMSitEq7Mfs3UWD8Kgh
g37qyd1XmUmz0pxnH3uONKt4xvG2ZRdBjOR1XG966n55I9Y5hPMj6Jj8Q8qNV033
+lo0jqMwmkkOXR7pBfH2vnbSyS/oqkXoP7dXcwrnrVu44CAv51nw2K/ZXqtKGHVp
zlHvdYWt5JU7dCPRQfCZzTd57GUV+90pAqBmOzhQ5TSqiBeNmFoIi2ohD/GxIF1U
C05QXmf+000Se/NuCZ4AVOvkqFwEkQcwcwy/e1p7hp0FHUpZ+UV3k4Yfz95gXo7m
ZIDLglKM0/lVpdyl5lmGTpG4qET8nRrBJsShao8YokJDLaA97525zUnjaBNjczDD
XCDyE2gIoumC0HYgw8RzCtz34KULui4A4AkK6pf9gEjc7WjLMejp7Bkdj6NH3hvG
736xlO2zHZWbGj/lS7oieRoTCHnFp7E9rN45cnrqAl/hc+PRRlmcqSOVCE8ioMIg
wyOI02HSBf4kWbyfp2d92RI4mg4GrxuvcUixHXCO75vRU9+TdmOXdMRodjhFMBsS
kwwQvaiHnyNuyFk3da9S8LGDig98pnQU3Rcvgn0sOMiVrISoLO8c1Z9jyeVIFECj
EPTlvZsn/P6MCuo7f0OnhYGAiBZu3m7sZb82UNBFLIp6sP4TmlC+Y1+OWKk7dVv0
prHj+hL8xDWYTXmtaH0TfnwXLLQxHT8a2kNAS8xXb4Ue5Tz3gXgsD3/rRPqvv0gq
Y6EoB1yARs350LQSyr5BXZ4QHEpxpvta2K7wtbRvP0KRtXzTenVFoSqg/c/EC5dn
emfyhW8NXichLmJg/nbqmCRlyhrLbsVpbWLJ9ROYtfebCq7hpiiMQk7/oi5oYz3f
Da70GcwNZfkuuEJc70uP2mM+ajqATm2IWra0+iN7Fk5AthRf3bYOOkizflTSQ7SS
L9CDxCtfzs26aDAEH4/EDphuPJaGQBMuIeRCA0dTwghz+D2ymXPp4rzxFtDt4F+6
tzKnmEmMLhYBQfoM9QpZS2xGUTunArggEJtEMWDSGYZ2YAMZSAYMpdClZWtsiMBd
oUXjXeGnm2tTYBFmrB98NWHkrZspkUsEQnd0sYak/v8guVGRxra5DK0CmbAWdcrl
tO8gLNvSvCv9MfKYT3Hzag==
`protect END_PROTECTED
