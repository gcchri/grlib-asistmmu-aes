`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PNXpY5J4su2pVCX7dLKay7s94L2e9I8xTm1x4cEqjf6M4Le3SSezv7V2j3knCFeY
U7AGa/I0ztIan7Y+rHMoq+MxkjXI4AFecr1DToouCjLnh86kyy4UH3di2F2aJJ2B
6xbsNiqTNjElrGjjr7biQXcUOcA68ZaWe0EQG4TzqNU6ILCxxZydi7WGW9VGKN8R
fvR0tspKyBk5LWEox2T/ABws79KElEHvknBvIMenJeVaGL3hZExhqClZG6ihPiU0
`protect END_PROTECTED
