`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TLI2YZJxyW/25dfe9Qb3LySFmEmfawTkia+v6rVBxzzHzrXazR7n1Dww/N+v9VK+
LUIrnFomsdI/Y35NXSz2VvUEt7BELNsBUXWLKNbtxkXtRMxi1pSofcI2GmIU+Syw
EHSbNLsuM4jil61N1lmid8jkvrk+BgrluwATjPumeoS/UcxPdazJAbxDmdctzZ1e
0T5xHjtPY/TG3MUgYPuf/gVsRDUareRZsge8336G9rmA6/Ie8zEeYjlSd23vER5v
dVomFhYpTjGc/e84/+O+wihTAXdw7sn+47tJWsjshfpaZrIL77YYj3SZMgVQVMa7
CQyeq5wpzB+xhbP0w1xYK3CHGgn1NAD3hGkYxI6SAt8/SNfaqMTz9vVGIG7LNFeI
+r+qrzZeIg9q8yGNEYNrR51yQu5kOYNpocuneUiKxzlt9dkVgvpmackmW4EGINxL
XZxrySixlpdonRw9J4UaHRy5TYIsjO2tLcG8EGwrGT3NF2UgGoRqpqfU8tVuCyiU
fyzwN3pSdwG9e/kZukGAos8p2BC7Qc4b8KK8OSxZhR/q1HlmfKi0mw9baWEGTGR9
AAYI0wWySD3v/yd/QpIMlBPdrr+TO2hU8iib/WPXFYBisy3TcKPoom1Hc185eE/h
jTOE16uYy9oWerVAhtOE6wG68tLzBY5shrvk5bliO8MOa6dSgrxrCMjP7TW9m7As
d3Zzjw5wW1//iAYkTSkoAynfEYmx2WtsETw++q8a/pOwWIW8U9cLO9gj5xy5oXI5
DJtQh7YnPqFe3iTu+3HaxLU16IxT4wWLxV7KmC8gKVTuiBkPqP1+m6ROlodQMX2o
Rb3BU/9rbg+x2/WFSXMeRaTfUFXhsgjDkinOytH6nuTntSQsHp32oLZK7hMDK0yy
MJ3Viv/l36pXxa11NoDE3VHwVaM1f3g7Wozt50VlsWJANEG/fWhXAidzXoV4eDos
2qaFqpdjH5Y5Ab4Uz05aPOcVVNJOWuFcRpQd/8AT5STt1Y+1O+3nVBLMahv4sUKU
Xo68j9V4/FDPjAw5Bbwnr1gssEeolkOiLlYSm4Pd7FnI9t6iTO0IcGos2z2oCfqt
xMUP6RtXuEa3//pmGa662WF033RNTQ2dzUENlcrYiBmyTD8eGxYT4yJCx2oeFNJT
hzcegQoF5GcVnFG2uB/jIwXrKJ0pWL+kub1C+fr038yQVD4RWpCBxrQln3cdzoQQ
bwZLW7QqQMybvm4n6jA45RdulYX1Se7FrHVFWjZCRUpEgxVIU+/TPMsTcCRWhSNA
SZswC2jKtAlQWkkDviE2jTThK4OuuYVvW689NgpG/h7udwz6h56gaeHPBDIKz7Aq
z6n7wuzwi7g2je1TKG2XbdJIMGhs3xiE6qZxhTtuSfIyFDM8QbEaKBVfDS0aTfHC
S4RNnSzjumd/GzeierGQp+NsUW+uNl9MEpgLr0vQFqZYTHKjXMW9NndRtqyjDdWq
XhhPTFvG+Hd82IWpPMgO0g6MJQHC3zIEVL89hShtMRFYgyGQTWSYYwT2tyIMu4Qe
wi+QWca9O1t2wkxwEEmKXOgZimxYRtpQKUFjNWXD8rngP0Ap3KotFbyld8L0TcKg
TI/52z8+tKZZFfNDxmx5JYMVXXzLtQlBdmTFXWkeVKWs65BKdbSsSg5p3isO+xAT
4RUqzVkqsS3bqaCT7OBc3lXK5z+yZgMU+0z2ULIdNNLFUCMcixV7XJLe+FAkg9Hz
Sbq9LRMOvc5gVjg+AB6TJZAAjg9lj+bsdVfxmUHXO1Cz1EbTV4P2wpsLz1Fvbr23
keDe+uhpHjx3ZqlVj7IQrYHgVeiUBNp/Vv0hfJ+sNl+78ODc2mkchfI0Gcg3iNA+
GFSSnMl7WNS12tFFjFNo8o8xfRFUNbz4oH8E5ezP7eUD7vd3tFn2hb0mVVaCac2a
MyzCkIccTZsgpJ+A5LTeYFm0TOj3Zdii3jvqzghg3hHFfNXFtpjE/WHxy3ZShCec
wIqmhjd9+uHdpAJTe7Z5blj6wtQUKVMXK+siL6xx5NBTidoSt+9TW1m5/Exaq7ce
xL8PQka/TK73HqJgkNFsq78po2lz3/z2Xn50UKhxIBjZIfDb/Pj2xNZn8ugvTrcj
BiCbNmGw72nIOt6Rhk/IF55tpi0zsgPqJjL9Ow8ugDVS/BMoHLTGOer7ahxjGVpr
mbYVrr7qGJLQxfw/OavkmLbSClb7A7RIiqp4biUb7Ag5eNbORiBNkLkHknoHFSPS
s0DxYWKjIriBG96Kaox4LNsqwR7Pb5eTGs1Gz6vVfoVe8UocgP98145kFcYgld8k
So0yBA+fCbX9K1ycCLftxZF66nFPm0vvBh8PyWbcwpHEfn+bTYf8MqbHWXEbZ7He
gEPTrrRvU6uLPAaOQ1r/WpmZYLMYCd6/CeadjXyFTJ3POx1oUjZuRn9BjTUYoiuu
h45ZShf11ZPycdXk7sMJ9AhfnAHpApcUEIgmoifR2gAC1/tEBSw/ojHxrbfMDAfl
dvxN8jJyM8db8qq2rE5Oq1PZ9OQmu2tJzPkvL+AtoLJg67XzWE6aZ45xaEOt5A4V
uWJ9peS903FRDd6hC7XGM3Ah1MNsMaUxSwSz2tzpIxBXf4tyxntMgDhTEYlEPxjI
bjyds6kE3eef3OpOHZ4k/ABhsurZ9iOWhAfsBQvMRsylSfI7rTVmo3z0MD2NM40p
BF2knrZslTgGv2Z71/6XA2gVF3tsFOpZsYkV/qMKGmuJr/EgooU8arqZY+9swWe+
4L2H2fXShx7Y8E3m9l/1NE0o/ZHLEOv9LAht2Iv0ztXEMYBlG178ZZNQhA6GREsw
sr21z7fXm2mIRVhqVIouWHr7artxuxYZt1YwS5nFkxV4JyIJFk+CG+MjXbqkkvBa
BBJTlVh5VIXV00RxJ0o4MNaV4WIxgB4hO7FtjauhnE7eNXnVAXnYxuAwxhHSNLcF
B0ZCpQ24+r5QCnp9J7BFYjGay/TEkTucKQUn2mTTePpI++58zdtdbKh6XhNsAKXW
BxDzFZA2L0e4ct9GRefl4QNhLXnuZAbIjBsH589O3dhxXTL+JcSIwS4SLw9lJwqd
mQPeIqIKmGC+x8YVUed0PrD+cNHLf/HvUrw8DrtgdQYIM03+4tzDsEyreS2Szf10
PQyWQ863eoXojSHCDT8aYS8SNv1mV+kQl9SmOk3/KHEu7jUkilHq1V3lbJbL9VR3
1pRawo0YyAdvSPIZs/40cxv9M28cB65GloYRpI6VsMSt+xyx1UnNDZzEqWu462Yp
A3Py3dYgYkokm5ntrsTI31/mcfAEKAZ0xEyynyTLDyrZw10lb1weJyQA/Tf4tNBF
o6KUD9z+d/Cb9hccmt3U7Xur61hN4lc2GETiNCiQoMOjjnbqzEOml0n4bFy6sXX1
f55LvXaR1Rp3EFAkJiLmGld/DN+/Gf9lZEPvU5Jbq5ww1SjIYuqw6y9ShsmdahD7
cPTUeMfeJ3oAy2spo8kKWd/DW/F8ElqlVIDm9JlItARr3JKkv8HlTK/nufyjxwOk
pFAZ/ECuzMrH2hdSZieR+n0WW6T7LmiaH5dHcWW397vYNhhS1Q/DOXn+BBGiIjQt
ReGlNIgOaIsTIQoczHHcdr/VFvzIM/okSXbrz0Q3knEbZGB0Nm3m8/UEDetwK2Ww
Nrrc1WVv8B/j3wMAKwoc8SG4hnZ9WFWcGV+3bvZ8AF2JNsr/63nkOd+qoHIQcqKp
aSuc86VG+DxwWtAgdNGpuMESOrW4TzQmXjUjvoqZtGiH215xham9CibzRfeqwJrV
veeDs19BEThCmnGwOtxR35DqAxi/KwyRruRhbQDav0JXhyzjkQinqgPRVjQyWvgo
+3aWqySxAkuu2Z7jPtIpBLE0FYCNZwq3YCIM5rlen+kM8VkTpT/jGtEqlA63I5RO
PcBA1wRcnULQ4PKo5lJZoMKD5IWic73xDxN66kEHyos3tMskL5lRKbnz0HEYB5Ez
sxG+5e4kbmy6kFQPuMmfeV/we74VgEkSzDpy+qJIDGTmzPEEU7V6DQDKjELRuUqp
T41e1wWCys5FUTfTCC7WaNoECU+LbzC611bUrY2Ia3L+HeWPa3yUzQAAkzPb5+pw
xEZeFnJdWPzD0OsoGIVeHWScv4+sPwmzbWMPgaVzarddQcMuNTS+V15hwJBx9hzp
z3hVK3IxrSpCbXOuUAiO4gLmxt0hw3OHFOWtMJ56ZFVG1Tnt+qcrIJNxAudj1DRk
/ZD36NlYTzpfC6I59KS7Q4hhvVnFSGbXou6H25RNJ7KRwteWZLBpX2dba5Yq2ts3
F2onPW4Lh77tirqQd1nMbnwyup2hkvLQkNysJB188j5BMqkdtluBx/brSq6kGEkB
tK/t3uUSMDiqbIklkqmCueYgevV+NwSCijzDjSC+yp96gcTU75qhTcD9dEI+lmy4
u7DEiz34+Ihzd2MlrJ/y0FHDuXOLOvC/WvEioYMfRQJASApvURqJrHal/ntH+zF1
CAITKTtBYvGlI+zHCl1xs9RM3zv784PfyBAxh4lqPrmxEeY9FSeHjbrSITQbNm65
4nrH8YbXnkp8ZCJ7mhWedu0eGZmmB2CiBf9W1Q0qSrA6oap1vlkRdUBfRVHBcyTI
xuO9yUbYTia8wSemhYf3cDwLkZQdVum7sBP30NI1Gfjev1Bg/gTtug8idKX8pfKm
8Pcn1UmkcxI0/l1g6Qn4lR1xKaqjm9754zd/dY5LSpfJ+1yZmSjbwAXSnYcYWL1Q
0/iR83oHflVIur+jsSw+EXoLD0u9MRqliCp7lsNNf2ZvkIifKo4wKkcDw3OpP6on
AsJSIvUaOC2U+E967aA7fyuCGFrx9yk2X2Ib/0Eh+2terl9oynXlQWmGTyAvr6vZ
tud8vzNwqtNHRPrmfGI4A35RVW8qyUjXCcqfHuyLaLAI94HgqUqrtyLqlEBU3PTd
I5U2/D1JGZ4kMPlHoLZYHivn+DDUikpljdZtV4zbTOpokr3NLE8P/0FA2VkkeY4A
IidD+VPXIIfCsjTTxmJiwctb8/MA8kNh7faCeffQffd/cefpdEtUsy2AHi6HeEbI
s0K9woD2LBiGFU1AehhBDJ+mFW28HS3CHGveTwtXcQFdf7Z3HYydkZm7XnVOIcxM
jV5yQbQPObwRiOYTbelqzAYiCRU8ITkQrCXw6EzCN24oAH1WjNTmo3ANdmf0/mn6
lwazHJBmr4yFhCavgCsgSSqy1O6iVSDowUv8vcqoizLbCwbG3Bsy2sgnX62byOxT
iovNd/twcWb4+AzcUvZezHIbKB77ducJy13NTfItKETp/JgdCB39eyx/YWaAwW5x
NrL/iQg7j3xwa7vT/sGk7iBKfArXy/BxR+BGLmJNpRgvaXxcacncJK20cIOAVi0n
`protect END_PROTECTED
