`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3BjxQky2Ej3PL80YYzNAcCyV70S2mPU/JAz5XpstFqS9Swir+zcSpFD2CmY5mp6D
tmvuhG8vgmHUR8xnMIpmOuUG4CiVaX6ZyFSfYrDBLnkz8uXcRyF//1N2G0p5+sPo
ixWl0F3yylInq4PxqyW9ZM+TMlTp8O5llsW6HYUb5sNIcvwS870g1BRY+4UhqB5o
Oe5ATtN2i2bRufx3XGDAwjNeBPQR2MvivIposMn1qklYFhUpNomt/7sgkBcVJO3V
KWptRd8ichQ+XP5qeOR4WwXCY5kx7hE3nvbqdXENaoVyXP+At6L+BJKOUMWJL3xv
QO9V595Co2XiJyt+d8+P+1Ia4rzfoNz4WspA3vbea6GM8N3oIrQeQmlqrVmzHbeW
raxZ04pzgAJZQET9YJNYlixz+tRf1AL3e95hV2pWYP1nh0niqr2z4TVZSRj/jvWB
bFpKYjmSkLD0d5eMPD/qSSuE0E9X07lmnSbLFZnavQbkDyxPHztHWctFpVUzve/S
z/9PLdbBPy3IzcIa0GHyq2L6ucEjFZEQ87aIKep//MeZ12+/n1+V0sELdsanzX+z
`protect END_PROTECTED
