`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aov7EWjT0k9GnpEpnYIGOS9Xa+OylyyzgTEdpxmUQd+a8Uj7e3PaXhP12SGF/tev
a4g+G1LRAyrrxoPJGJmBd8EiBUQUYdotPDfE5LC8N8ezPvMUMPUBilmYddjzdkr9
qeZPhQPMmEhjHEOtlTRNU/+Mt4iM1F9AST1opSyPf8RSqGbEB14dR4d17UoungjT
reCQhtpqOW5wmPYTahHIBI99mC3M4bzUM+aeGERrrAtvRLCqE/5U5cUe3BKptUPz
3vbdnD/ZUlgfG3oAm0+YxRxgmJMoUF4nQOFwsAN0cNUI5UF3MuI6Zv0QwBIB616M
kiCjsAXHlQ6/CvjTQ/yahKD8dvnQF9cuQRH3iXvTk4CYdnNgyre5d2qMk0F2Kxcx
fHXHMvC1SbPeZv9/JMA/pmSvVkbXDTxEukJtMP5DjBpvAQRc8uzKGYYh+35fSb8E
F4MHLlUVLrPuPJmwpk33PyuETiN4uzFQoJiTcv2FsYIGk5AH5HlNZq0fm+pveQin
2trmvcN1Bdq/Z0XV78up41G5g4nSJ+m9h/sP7ABMpHcuFCSp4JFpRWt+HeUhMNnP
zAz9zqCZy0/+kZ4GRF7hg/VXD+sDpE2gxfl/SNGJgu2RkPeLXHOq0GmVqFG7p6s1
zai9gEtbT4fyHPEdqOy+dgBnvqxKgkqYIfuX3Evk4vBX9UTF9tNPPl37B/NGJcQR
D5IrqaXdu2qj5p7nyMuf2bkog4uIbVA7i7uwpegA4XF/4i+Hnq0dOH//MGRO5o1r
GlRKVLX50aG/Bzeq3dBAJw/ifd8d041yTN2BzExuZSzILyNtCvptaT6+Kpa/OyNa
pq1SXA0lN77j06ou3QG+lEg9wXifLHPLUkk4EXPMX4NfCUsUjOvTxb/aaNapKHlA
1t8ZWhOPj/xnNWdwJPVvyA==
`protect END_PROTECTED
