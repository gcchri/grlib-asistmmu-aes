`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qBUHb5cPffiwUEwzJiRiiktlyloo9u+xfGBJneEAwXPJk3q7xqzEgtmX9ClNQ/+1
10MqKLgrbXPtqfz8heiSA3q3nU2fLuVoGPACXaum92GN2EAAZoP+DxCu7Xqwq2h5
4nKcx95jTzXw47sQXvs2SzJRujyaeE1YT/8ewizAa/h3fw4LDh7W11zaGq6o4efG
trU9L6sk5fDs9ZT9f1tV1pxQiEYLEB8vtTMo1xoJEEdrapOEFjqNRgyTy9SwnZrf
8hINNsuxL+Dm10nsbNXEYVhXX+0MTtJGPTS4ySs+opIp2kNOPMgoYMI1V3FPFNhp
e0UXzYibvloXKLp6AC9avqWRBJ64u3HVWmiR7Vz/vLfaJGJmjBrir/3pPfE9O9Zd
mx9m2B8HpVx+FwOBNplHGfghYh0xqDXoFq+HNsfUvPqx2UU9ZIeVB+dhFWvLPpei
8+wUMbaZIJR7iyAlLDtHjerF9WBKAKYY8ZT0JyLPwCLVA0vwkfSDPQVzmAaiwS+V
NGicQ+irNM1BCIklX6SajhW4J0myo//rt8V0hlQGcxFR6oGww3rb5w9jg4aYqZbZ
`protect END_PROTECTED
