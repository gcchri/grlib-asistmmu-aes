`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9R35BjO11CvnfGFg/ixla2V8fGBfEjD/xJgDwUCoR4JuFYlM8yLrNRO6tinP5xv7
M2oljq2LiQ0wne/E44lA1OJopUB0z1PGVhD+rJWrbVRJj8F+Xp/f77/hcU8/l6SK
H+TE4HVY9N8pULrc0Moy56MZK03vpunexTEGA0bZhUrN8gTVqbJepxCadPfpeKhn
v3Rc8XLyQQpPMuag54/Syq3HhOfupqF1SWbBdFe3lR+3JHodAJfg65RQzAqGzawv
Du0UdAqkmfo0i08jPHb2gAk144OCbU6oVapGjaLU+TGnnDPstWFK7XET1MT1cTXu
T5g69iswvJ/FHtfNE1kxQCpLbUHKVf4zfvk9zx0TE/HB/qnmX5vs0T6UyD4vo1RI
DeDQtU00YLGXVqHLZkMyXBCVJ4l6YjVUs7QFQHRfp5f+Xs28bN+KhB4/jL5OhQqj
s0YhryeFj5/IBMtkJR/Z9xbXuNaoNstD/QJyEm94i9+U1Z85zwKDyVmfGuIQF4dl
QGz8ZVORIa3ecZncXRlBpj9Ey02YXvVXcptNCxBtvJx1WepicZwe1VM/ORX8gPa0
aPJ9kgsE/4EaaV/mEtT3Jqpr9wZbe9avXNWqGtKIbw7qiUf9CIOwdlQiha/tWUK7
bY+n8bSvEKRkzEIYbaLLx6nc5YZFpA96FIahnlW2+HDiWTjokGSSy1b/OT8fYXV2
qDVhga9ae1GRLwECPI+zAFE1HxVeUJsSLpalu1qNzKXJdRPHfLvoS5guYyO/Hs6S
UwJYXtifb/nMbK87N7l8j5bd6CgjxG8J5cfNagwb7y1TO4cvJrJVpvVHC/0mTzBF
dHalhiWaWO9yz9Ydmh8lmvq3ce0v6Wilb6SnqHurhB/GmouEU1E9ktFjN0y6z7+H
e+qdRKR9qh7FLrUcDlznJThfl77F4GN8Gu3xnmP9448HpYelQwPOBbG7nt7/lDZf
2p1Aav42//bPRKstie/3DWXFpeMZ+MKufqAPIXfG0tTbVW8mxbAxBVvCAAhqkioT
tizuzuTmHRZlsWQt/zMZkNRco1Szt7lEenmMBREGRvBpj7fDO+NQWF4o1fi8a3PF
4DUJiYxDKU0+JHesVRMrbWWXpy2ckbsk7RIfDFqG6xQaBTWt3q+7WtBf+ZgtlnY1
vYfSi9KEoDyETHUQCruAQ1dsA8tX2vsM/FU76HsKmO1azTWXDHxTkfKcHaZV/dE0
NkHevnU7Ll2hegoQbhT1Qp0CSVT5L0MOeRBqqbMJk96QctsX3nydr+W8BJo41bDy
W5NXYKCCup9sp/pIwNbdCMPOISr3JmYUJI+c4v0wbTVuFZ0ytpeWcXoOpB3PMwWe
qtaCkSiNYx/K8+x+0Y1t2dXI8qduTHtGUUZKc6Oy9DVoI27l0mJpJ77cH/lhRMBZ
O0VZ1joorFgxESnRkIP7J8F2VOisDzkSAszDg99loq8ERPWdmbL2bsxwpOXwNsZV
d5RSxLF5OVF4uRMs6jB0qa9HfS+XOJ5EPqUAQ/zsV5NpMmhv5WIagcgC47IJj67s
`protect END_PROTECTED
