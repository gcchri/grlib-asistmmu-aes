`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pYrV6ayNAiRNai9+WDS1woDIBa3qx4ZQ0jBKgxzr4tV3+IcPEanTWlqc8dX7aERa
RvkdLBw6oomlFRgtDdvXnoqVBXVV+fx0neWf29x75uavzdv1mdakGif/yC/UR52B
MC7UVkKMUY87ZxuBXdFPM1UXX17LS7x7NLbTE+q/YNRNk2KJeUNSB1H6O5P/c9Bw
Cp5NSl7lNvojFbubLrdva+q3eYN+svTVm31FmJGVVek1eDYi47UWYTj573Im/Ifg
KfOUUdLm2PNHg9ySQPNnb4hrSMfe8uyyQZoL7bG8OWFpPP1QoLyFa7a0iPAY2gFy
UO+KCqNpbNcpdY0yk3D2b0od+KlIy5ghQHobBOLmmuBe+8DGNMSFlOzc4IWu4sgZ
G7lLm6hnqHNQBAEdilXfO1rsXNVwaRbTMkXNkx3ewYGn6eUqWih4DtidzjfCUPpi
rqNmP/KKQnE9X6d54jmk3VaHEt5Ue6hoL8a8GxRG2ktz5pATEIsb8Fnkn1BHLigd
iEh7Coooo4/Ijf+cS3hstymPhUkxOdjZ9qKzIYm+yH/kBBG/kiT5f3rMCJoSRLWN
wwgKnNX9udtqMNhtY1Jvlb6JrX2/FU4FCiOSqEa94x0rZ3oLgV13G4df8HI7og00
TRDFXmqT6zbFGnZQRwatOyFIM3RpjqPzxzScn20MaVVM5/hOcJTMKmMGC51WA2+5
1/qv2E78g6C0HReeSNJY1CRVmJ2mpoLuD2Kx+fwAlJtBGnTI0hUaNvAttrp2AbUJ
Bz9+w7ksuKWf0n9WOGVAZA3aTNBZGOqL0puEqeflIOgb+51/16FZuy5xLiXRaNqR
yF36K/JPFKijlo89fAbVb8awn+skCb74gVH6vE11IHNsS0zLTBF/lim/cyqfNl7E
ENAU9qBrCrssws0IE3bFnDoiwUzQYsX6oGnR5n2SYGpUrx40HVvn11NUrQe7R5zp
`protect END_PROTECTED
