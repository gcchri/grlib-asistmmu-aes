`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OnwM4/7wD0g5o73pyVTJNexuqWTlcjo2mQ32abMUzLJwrkKk5TqSFkMOfJ90/fRv
6CKwZlKpwHCytYQvbBzCkyq+0j18ja8Be1htJb+d1yDos7WBt5eJzM/HxpL3PDWp
PSTmUFlXo6wBoSNFz6905xOOKY2iKTKS0TyxecJYIHZf0a5/xvdNSQGlTXQoQQTB
II2q11kO6yUbbxBdwAMpZWWpl0RiXr9ExwOkra8f8qC392lXf0fF5/xDYzM/3e+t
PM2hg7NWBow2yP8iopTHpF/kITNbvEPydbSdiS6MZRg=
`protect END_PROTECTED
