`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
esgbznv4rH8QtWYcLaxxk9RoUyvbMhLdRXwe/fuYZe/FtK1bB9R4qQpPnZwbaOpb
Fuou+MimM/zZVHqicL+S1jgeidpU4FDZ2fsHN3z/u/K5vC6RiRuxxVDaLukSzILn
7UG5uQYhhv4fA/rH4ZXvQkvboDLtgzcXQGBsQBHk72gNwllBViomcUbOa+hTW/WZ
S9tTdbuaEGQIesizPgseGifdX7PKb1w2DNLEZ9fN5MaShf+Vbu30DrzMQVNm6Sqe
1Nzku4yIqAMhRusISe6Yxa21CzPFpZTR70yoXF9yITZy8G/4v/QMawLUia+DgHCe
nQw4l0h7ZOtyA8Fi4+b6putnSgIeZAH66moW2f0AAEAJTKuzXBn4LQOVkQWZoh6J
Bi+Pkkl4b+MELuQr+RI8a0Uk52cjGnEFTLQNkwel3zo7+tHiHF6VGSBrktabmzHN
RDgwJPgsyqqYHCn5Om7uG5dNqRcxz34Ep4skm0PfgZSRMlWLrwSqr6mgz6Azp1Rq
zAGpJb0OxBxZNOr97k18WspgtdSzMy/wjdcTW4wL4zZ4NIk2lIGV2oe/jA1svoRJ
9QCxOYC7SdlZHoQ5oWcUTB5F60WUIk3IKUttOm/2sKk848FgHYWugDJMA1LR663f
WZplClBlfNrNHTTiqVFsKDu6RakSHVdJuH0zAXC+iY+bgt2dQuzeH0gtF+DunS/T
`protect END_PROTECTED
