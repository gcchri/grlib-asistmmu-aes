`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sZCWZUvmPrHJ9zcCrjpc/n1WBApUL+eFbRCN1rptLFXu9SCokDcbmNqjJxvWQtSG
JS336YsEClJz5UV74RLIaRqqonXqzeBP4J3jJpD7V951XLvBfuRxB5VvPZxTIVvX
V2x7ffStjQi1t9DrBZCRbWRwZHgYhIF7ljzZSnrIQf6BSJnGb8iKBI7vumOytnQL
3JSvmzx2Nc1Zivu8Tk9Ija5bnarjW8a21DS5hHVq47B6TuKRCWDujQ+xZH4WLVYu
PXWaNch7niKGB0rwESpWERFAy7K0a4PD06+4YmormFLGbFFZJGIHsJNTC0wbdCn9
l5+uSkMVzKriNhI8SpNRvPQp3tUH/FXOs1wjJPWLArM=
`protect END_PROTECTED
