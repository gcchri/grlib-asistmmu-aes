`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jo+JZNcegc69cFa637KxlE0qNnKOB/m83iaTkescibKRSsAgdEaYZutQ8fUrHhvQ
USZp5b5k3W3Qxb5LOwWJWIbJzKui3U/s9/xnphf5zPKvTvDjwLb3ADxAB5W3ojEk
8CLxIQWWMhj+bjsb8PZyRZ0cz1t+QG1zWeI/p+kdxYRRam4JtF64Ml1wSRaDYZ6S
iqZ+U29V8QTelKH19y3NWDB4OOVsw3wILRfnwOas52Ds+WlNNLpCEjSHl6S+58W0
b62uUY7jNA72e12kKTigtP8KkWi4APt424NxPoqxXY7Tdpn3JmxkhLWTiyy/SwzW
YF5avbWW1DdJdVfbPBwswXngfjm5iwr6536cJGXbRgTk4JTcKNBUzMv0PXp4sB8+
GiY0CQNNn4A0CB6lRKLvuK6/THHtrK9OH+tkxXbFuctgDNaeMK+8sH5ghsCuizXX
HiLl4PRhcuCbK77mi+4tgG47XtsWCNuof3YkzQfYXnle7dlF5yKRVATe0wDQ4Pqc
/6cApZZ/9tV0JUeKhHhCjMNtIGboNwIIqIZo2Uzhs57l8X/VQGHQu6zIV6Wg+AH/
tWy5Xm00glzSe1VNUZoT098D/ge7D+OIVyk5zKx15Vm6fGG0kO7vqteSPuwXfPPy
HFc2QovKlIz+FKmveGF1YYxg8ui7kJrDZXuV05X4pqXhXmBTksb1SbrB76yzlpox
flj7VUxgdLXXxO4X851mORwFqLHWXlZTyF/XsuyxlhRYqmevV78VdYCrSyKF3Hz2
0LYsDRyh/Ffv9WhSNE8RyiRE5plQ9s23LncEHa2g4rvqe+X77tRl4HT75ey1uTSb
uD7WJMR5LwPC2imzRAMiD7Yz1kH/bGuMxzpW8ZBeYmaRpk16BgGTM16Y1q+xAbYo
bl5MIfVgKH1z+V5MJwmLDqdG5LfQ7arp6+fmKbtQlLbeZI6UQrn2d5R94eqdRvgZ
PcSi9qTTBybTXvpymRWBIrsdXkinfV/dYj+bAnUpylW9nE2BbR8Nt/h15fFn7IKR
xz8Vs/aAsT6/ZLB2eo/wYfqvbVLr/ZPsY79MnkXIPnv7BnZ80Kl5hC6zAMb/NyYC
vLNBYYx5KH0LNxbOS9zthcjplWCENw262DhOjSAhsghnT7W96+I9KGmnHwkqyJTZ
/cshEAM1+zzYEjjIIm7iiQ82TZchcC82mcM5OiuYU2NMdG+9ZKbyiIzqWMOlvXug
UTZslUm48Cb7rX2Umtjn/egMYdPrefWOoIf5t/xtuC2e2Im+94W3SUR3CGOziE9P
MRORwHuvk7yvFCp5Cdf3n4CfaVaS8agWIkDs4r4jFN+hVTtC6QJD3FPkjR23QEKX
FLGD3eYUPv63JuzSgHW4fDd33Q8Pbr6P64GSVwd26JjhIRQew9dQmfJ6Q0+O4i44
zlbDZVzCDfuVdCvIVDo6V/n/AA05WcIqhw+IE8V61FLHQ/PNtMkIBvmAps6MfIXH
6frkiRO3J2I1HJxhQ55skPUvKz3a4bvC2XYVmSWsM3qkKTmJNCVPZf4edXjAIngt
1B7Tx6tlpz/6H/sCfXS20zae2V86MqPV6iwEDxkj2WAR6FxBqEcnamRr2pL39Rgn
4+0KCZzyt8Phzz4GCGwDYtOJb2/NG2Tsit9fauWAYywrygU5uo8e55NWJCFf207G
kj80GW83dKnJULLOv1ERFjEdfb2tnMkwu67ovid0GXHtWpMGlA54HmhcN9Y0G4UD
AIsXMrWqYdn2AN5bfEr+JyyFM5V8dHMgJHz91n9uXqs7px3SZpQP3oAgZ70YcrqL
eD9y8Zp5gwncnA3+2O6D0R1452QowEub/SYp33bfEAbeZbxdZ+jbaSokEHKZAN8s
QeTOE8CTUih1Bxw/t3VDjIxdHG1iFBr5q8cV3g0jXrNoV8YG3bi4Z2LVyjgSdgMc
r59SgAh0mcoV+UiueIM4wW05eDE+qN18r9hT2I9cMxkv5jr4ayFO4XyoDAOK5rXP
rwpxsH73OFpPftsHkTYWsVA/SMQQuamep999vYRY2nDdorXwQ4N8Zm28GIdT7wj8
GYjzJOdpcN7VRvBxu0UvZI2d8kEy9JQb/yeXXq389h9+/44mqemh4oOnxhL6Ylbu
gIWyFwQ7AAilfj4NvGIjIsQSJLd6/hTGB+dcL2d2aojYlDtpYJvlx2Zfr6vDQtIL
DhM72py5Dc4txYhiEjc3hMCQP/o9gYuvj5F5ZHYWuXiCFYCKuTOcnQob1r2q80O/
pvUOPNza6qYT3efmh8tMfPRUrHQ7Bthns36TvLyoXPKqAU2vnvbecliPLuFN5SOD
xhkIKCgkX5MDJr+bF2ow/4pnUM58ceK3Y6PgJf+/ZIZXxmjlEyFN2oEmn6cs+NWK
1QTof7oQRFfxcspihRE+bWYt8mkW4bDBNcbC+b4Pxj4haoN5IJRb7UlbYnqA1au8
/Gue81O9nvmNWIF3bMH/p1uRGCUxVAG1J/cbaNfgdfGq+SN4uxFukjo/BepIGDA7
JO7uhZb3vRN3pznHWQKURZ/0B4OdpLlE+XVhtnQxitPXlXxtaeoq8+hadv/4ziET
dm2iCLOxv9xVT0WdGWarKCspKe7f9ftDh1GqxGesk1jr9SvCpFSfX1qvXIpIWSOJ
siVZhW0myk2tIQzW59oi/Tb27+4Wv3xxIfg75YNgAgmUkkz1UcehXlhA5Nj+Bc73
K55qDnsaHNSUiCyrB3xUUjNuOjmicH9tWBBp9I4Nbj3nQBPQ7r0gJ5YjgYfve5my
kwjkC4UyGbXNsbZ0hpOpmA7wutW2drmXNHiYzZCZyhqfmfDgxvrUF+tcCqJw+0Tl
lvcRnPdxc0V6zL4kDHDa0BdjSNboojBqyg3rZA0vIi6hK+VVodSJAE25VsaFXS7V
kxJp2SRAVMOHxCHiS4xXQXHGrpGxemqMSMEhny3ho2gEXiSARp6HmExUTymoH4j3
EMl2s0+FGWJowyJ5qsM1gH3MI5i7qi2o05sOgxn747u6z/aj8bS85SjLnHJpntgL
xGKVaSSPoSYMyS6Hk8j2q+3moDn9dnz661adwVOiIq67cB4N/DeHz9gIFW/deyg/
s62yFTdF49mxUH8CRTL8hGBxssj07YdfpfNaaWzy+gIB0m2PLxkLoyRMhl/mkaXq
ne0xcrFvazKdp30RGoxVdXV8IjTZ7upJhalmC/9FOdypz3n68ivJcFtj++M/R+5x
cZCkyV8M4S4lsNS7LUnf6SlxdcUHYvtDkYTaoSV38keKMUDYnuttl6VJUshMzKsE
IujhhOcImxnG2vjx28UJyU1WMw2yK6W9luPUs8O/eSzuFbxUyBh15vxVw9T23bgI
BQxITNLiyR/ywjXUjsiX0YUKGmKgj6rZ6SPMNuWdoSpoXTfvA/5CGubs+72rRd9q
vLQnl0ntRwW0NJJ121sp0DX9k5177QmkGZVSniGNubdHoE0gmw4zLglE6JPjqr72
yhOoZo3eebbtHoiDshiNDOZ9llLRxKkwI+NrK6Una0BUYmjWyptElhfdvxeaJl78
Q0VJHANULTzGrf8V11jhLN6rKazg8WHNvVhdkYMi7oFUFJphdv9NY92E3ddADbXz
q2B0BPCCuG7GCVFBc+G8P0t1DbUQsyVYPSukwXT26EELyp9LUM5J/K10WdXaRLp+
m6nPrdG3RNtys3gPFmF9Kk7WhmBxskYqhR249AY71Pd+QwdBe3fLBRUAp6FaRUa/
buGooq1rBMB2iVKzEJ4F/2BIdYaNVsQEJ5gnVJus6aLuiMsaabCuU8C8e+zecjuA
QYTHiTLtdBqa6FdC5Z8TbZnSvaSmPTi7jItDqc+Sbt0DjFBVReHe/xL0CUDs3Ykn
NMlrLgmNYVfvRn1OwK7SYIAFqyc46LXk9CaPN7Hu+Qp07XAlm9oy3vICRaspdDFt
HlNZshaMn6f3EMDna8yyl29LcjNktAxSG+oNNsRK8DxnKSjuChOg8jHCtkXsDMt8
MUyR9TlAHjwK8+eAZ/eDpowkTuE6E7A+fsmqhttgB9qbkMr3jEeDDyk0MylagOzs
jdGK7XqZkEIxRuXnW/Swwbo8eg3ZRUHA6El+lbcGtrMEs8QElm7T4z9DjOXPzA7P
M6VgWqwO11WS5181+lB05nWy2EyuyE0dYR7zH2GntTIizITx5RdVVTb5uYLz78ED
2630sBTFJ7yTLpFhBtj7hNC2ILjMz3NHhlg9ZJV8SSk9IZDC5z1hRsSfzxTgXYMg
siCYmtkLJK2BwHenW99rY+22hRkGB+0UswAA66+t93ZU8+vADivUQto0PeX5g6xD
NINzV+U+tSLjjhe1r3mhMJj3Qy+C1T9S3on9Guk1d44431cV5ooP13lEL8D23QCn
rb9UgHFDS1+NzS8kbnRkoWwm/MWA7AGad7xIJ4AfhYHijc0xVhcZW0LK7xV2M2JJ
SQN49k5WhRnPoule3fXYVp8QMKdYpUODVgxy93MpaRf8Dp9TIisYr8q07mu7ibtk
HycbPuabVZq8Lvk+8llba8ESTJC2nq5RjtEECznYhg7RduwX7bTd6jFD7v09KkhZ
SoJfk3wBIco5GDM/0D9WtI0jzT1XzdUd1aMiisnv3TWahYwF18m3Ak1J06EI9OMd
rr3aZGta5lNyySPCttdsRCYmpayGLuuAqUC6K90CXc7h1RVsO5Mtn+k+ueeANc5Z
08lzQqjJBlO3mUM9VqWMnFTHpe+RkJBQ5yY8qU7dg/Np8a0ssY9A/YNRB+gxuD7C
gD9rop3JrXJ3pAdwMXaW378adGp/0PoAQ0u9HrTEAHvLa/JPd86Xh/coOi5mHIUJ
3U/d7LhhV4CJCzwODGtoLz5sexz/FKnfgRplcj0ECnJIEVkeKf/o0WpVKFCHlM3A
RyrTXgQJ9xxu3rlYwM4Qo95+hBEmvtDZV0upe9h+aygey5bGRW4SKOz8PtjYw3oD
q1fRzBHmtqwI2RWbLsHmSj5H7+l6np5biFPGE6BhpTDn8K5pMvaB/4133jd1c9q9
eTIttCGQhtVtUyr6ajySNheLojL9DbV2neWYQCLeTRkY09/G9M/VvY7Mmc2p643F
D3GHjXjC9d2myBp32KB+oren7YzIa3Mjg0Y6bHX/q66httaMpEsnDE6ElM7mH/1w
BPLng3kYkE7suE2ZCFY1Bx3YtLan9doUELmzBIpwZchj6pjqgXmGGNn8KK5zD3Mr
mXFiM163gz0SjDt4wQfPRd9OP2ztFdloShlDSGPC/a8xsponE1Ud4M286Hn0b5QU
fMR/RJItpdcVVj7BRyHPqzIKRyBcyYdChnwWQ+drpC8lp0A4mlQWzZC+ZpfqKl1i
553ljsf0uAVuVvXedqMflDNSGd4d4TeOpTzvX7SBNhuLHkBGVbd8ZSyD+u9lK5vY
Y0n7bGPMvhyZHaFyi2MAqoGl2CMiWBy6nww07P0XVh/U3RjOnQerKJI7bgIlQBiZ
nD9F3WeUZup7NcekYOi5yo+HAxuQ+RFJQz2Rhjc10AUjYW6vAaKwD67J3NF91gpq
qd65ejYdx1ywfL/VXbMkT+IPk5POyB2TxxHCYSNGd3polHziAqfWt8+jhX7zR3lj
xfnFn/jkxkZSHxu/2xpaJUHwrWCqk0ilM/SNWEaBBj7liffZwViJB1KoTK8r1RQU
afY1OhUNujHEXbKjojD51UhGybu8D2ITlb1EpLU+14OpOBijHlCFz0A4Uik5XV3l
8N66+x6CCOsxcC0JBuKwJD7YK7TG5yphFzjokRQVKUP6xzRLh6/f1odp+5yAxO3O
gMombj1TiIKK95zzgIQgaUWju0E7lBtAUcAug34OhrhVNekwUH6hL/9ltFrxULxm
L9FQpzeUxtXnH1fKNXtMyddTssdajVkuMp4zE5VEcMke5mOvjbLmcsjaL/jcz2Hc
ctMLx6AzOgPi8l8sW0p5APn266iaf57ete+FrjPeBBAZp+LiHShBRvuzAtjDORBg
DNXhqtHdbDXtugZCibkuHvlwKx1hPvI14qanWk4xRo8wYP4fVjpGlBYEbt/jZ4Nz
UfCtj4dHHV8h4Qd4q1C1mtUO0rqtMtgVZMqZWiKW30sGwLumBaFVzf10G6tsKmOL
t19gJERL/u/lk/comfMlyfMkKyQWm64yxceVbI47kQFhbfgRqLa+p+hQG/u0/GqM
k6G/IWI4XbQggCGlrcOOkwNkdRqJk9SFezvCS5HogOXQGxNuDoSJa+5xbQ72XTpc
N3l+VeWsM/vIra0Dj4u34AqXU+w0ztu61Cj5SAv11VOWEF5+TweNF86luRQbsD/O
5tAgPt9FDScNMOvBR4Ssj07ga41GM/Urjz2w0/hA4i/GjVWGpLv5js07gIChdm4p
PWZ+jRe35NkKn/X83C67ImtZRnr8GA/uPMgypTQSz2bn7hO9bmx+UyyYhBRAxSEr
0TA0NWNgt+wxjEVxWPd2oJOCAp8LjyVfKSh6h0zkjie2nqNxMz9r3A4n9DCgIY8Z
UlS8Oy7bfdoJqlYZpDtwBVK3XLaIWxbPI+ghj73W3Hv7Vp/NKKblHav5PZOfekRh
Gxpst+VJe/JgSjsKQ50sVaohhobE55qRFCnBMSA03ZhxwddE782ar7O90qBusp4a
rRYOFKeZmLPReKIZxPxvc6nNPG0C7l9XlNhBLV+pIFhrDlrd7/G3adi3d05+IrJ6
T+sCRHJ1n4RQoVdmJigSwicDmDfmicIR3aHeRwN9CAF8nqv4R229Pw1fKUwEeVQ3
E7W/CVwFhUtpe/Pn3e5um8MqapXdXmpJhhXOkxBItVs/fH8oOsqn2/4axTY01als
qWsSOmApWYE6sLC4HmwQP/jR4vxJFJhnTdHmhl7bapXKfqKyHIXiAJDJLzATfibe
XvSQDTlh5zipZdNGwnf5VRibUiYdhGxETdAgBwQgv9ZaWk0oFU9b+MDy7Isk/+aH
6sXoU6+sfWIEbPOZ9PqT32cw1927sTI7O2g9dRq4h4xiu74+UkWLZp28J7Jmda06
LSqqvoHqIWtAKd/UFm9iywCjuyZSw0UmrPAoC400MLU66yWvZfA2b83QDXM+iq2i
V8M7q3bIuwiwF7bLhiZfRLbQ7xceabo6YO5SD57NGSvfV+++UxEa9+D3QTLVFQsi
LLuh0WFEEdaXkP8Tgs8vZi9yDCAq0ke/MHKoYvzxI7t5PXmGEfGm2U4oAIxJOwV9
+/Z12GJEKUWNDbeAdV+laooYfEBTDqyTmYNvnmQxLxXwB+E7Wj9eEFOvRfZMPCQA
7VGp6qsrydogGSvXYI3/9CsoTFJ+qzKzLi01chjRKqXzRZEmtLqLZkGf8Xmh+7iV
C+UsWWY5NwBc3FUhAroUVtfCJvExcTAy0Hby6kmNJmNIaxE0xUcS5Ra2qRL5z5Qp
TGEvFvlD7ogIM/2dOGJwrQ7C49CT9KBx3MBfJpXdq8S9MAg259rI1Jl7bA7NYMpf
iozKaRBFkgQqaXpdaOiyrqmZYwNcD5QBj4kzIJDRr8xxDMXlSghA1k4M9BMFpOsv
PefWXrNxXvMiW+lvliJ1a1aqyxZckWQMenSdcA8eBZncmqtkifZ5vhubPaX+EFgB
NljBeruAPoZ8YPBnCOuTeb1so61mExj+E7GLIKPypVvSnMyCS3nWXSSTjRbUTttp
5WAnTUS9qyq0qZsCnaPxzlnZB3p3yR8WRr305fyPshzdKypbyX0VspIVhCqKQZgH
N8ABqt4SymENVmYrmgTz2Oh/20Vln3LI9OAQ5DwrCs16QVk8zJJp3McTTuEkag+f
aAjBR5X1goDWOCe11Bs+i+rJsuCX2pCQ7dHPPgnixQkx4HhmWHpvYYlYs9a46OW+
TfsTS+TsLI2Z1g8pANXMqHcyzzbbn3J9be8aE9OHipSAUgFn0vyvIzGHSuyiiLyx
2FpPsYCVszA5E6kc71cWx7jn4oIelDaW/LRQJT4w5lR4pxo9EOrvUIsN4IkgOgGS
in7r4A1iXtypveT/4jewu1+AFK3RrL21ya/4PmjxviFEYyxNcaUxMt0eGeOECTy8
JtBEydjd4YUXVbKoIZzUbOXhGKbvYrax3KtEAHXdJjAFln+u89bbYghLU7Frp1tI
ErF8rlumfQAR6KiKKC7Nx/8UBHXU9IZM87plfrzrZRr57aEq/tX0QlLTvD95Ca33
ucH8zATqpmwyRmagSDXUQ306sOJCxhD6pppLFdfJhDLSZ7ZpxBVzDotxWRUIpJCS
hzYkh708cYR9AIV7A7HLz0yOCy54OzV8cWLusWCUO2yBcP67f4xU1Hm1rmVpAjlI
2rJxK9QSNQE/0uluHteOz7qBXINlDZH2dglpYIolVSPMNUq+TL2yAZl+9DWdDpms
wKxmXw68JvONT4afsCXZl35BnWbRnlBUVFtelT1TFo1jWBBa+eiLrM5u2mIq6yGT
2yUXyTyx10kY33Eay+GobMW89VlDtwz191jkfvoxC+z1zRSWYN2KSQ/88dOIbf1O
oPBtahdPdwHPY9V+Octa4qD+KGzUKLiAS8zUQMIzQomiLoeQuyf0KSLfOMSZCH9w
SfZUlA6mRzeNBFMjfHXtV5B4lKmWcTMHUm+MxPbjrFYKf3tSPXoWc3R7LtDkTx2Y
Sp7TJwIW4WipcwxdQN5kcwvDQiIOygFjJn2JdamZlXhdR78e91js6lKOlVHU395z
fKmDPvfJMNDZ+si6RZPTTExSub4oihKkbcmpCgG8jXifSgOhQYDY7akMrbCtDrrm
hBWseaLLa+hu61aoB7rR/QEBsr90hESgeUfx/67xniSJdD3N0YxxCDEyf+z+GenO
scPqYGWuB16PpdJeReHyi860NhrFwrS06Ze9Uiy2tldC3jjZxuLAv10AmEzypz3N
AAH40mTIm2hRuLjfmQFmhq9MCdiYmJQeRfJcsB6AuD+Aq0CvAr/LEMT/5lYUo+cl
gvXoviTZ+l92OJtgMIXgEZLV+8VfsYJyBg2499nglRv9CLmzkt6I7mvHX/jVZbcP
S2OKXPQF0YsnPlVFoFaSukylfGf0Kf306lRZeFIlEUaiSGN7VW4sOUOJxMPjbxHs
jI8NLc2ONl2V0f9vHJXtqays5PafXTQJPAXWY7EszQ6kBdHCAeBJJyHZAuAUjTy2
p0cXGRBzMeAm8tmLlLevfYfeB/vjHULQ5G/OZ038+Qx60twReoqppRaxvi57glMj
Jm/r68VHsT0khYLB1TJaNXiM6fafAXLnKNsG/EV3hNO1dVLRiLkF6rRQf8Em6J1i
ISKvs40+xakQsCWZqBmMjU2zKgTamRW5mB0bgspIuiK2Jd5mfsGppjd2+VZLpfjJ
9XnN929H4tqTynjz7Jp6gzn4EOg18csFaT0cPXmNOf1K9Y1jEqKRaKJlBGqaF/LX
FHR6K55lO+xQPfcqsWHHRzEa4RLfvjmxsLyA5vDcUG/qswCL0HmCowtf0ElyB5HL
qEscL6+G8obr7RJ9ErifYbRd/YA9T4Cew0s4KRY2tvRxFAC9cA11DG+knRRWCMOR
b73zbH6HDEKbRXOBvLl1a6IkZzVQgcoHhTMoyk/qZy+J7hg/ykYt1+o/AG2xlTty
ws1pNeIno1M96WlzAZ9dyiFTptuedbJGKQSYiTJmb7aGDK0j7s7kYGMaoWqChYfw
Bay6ADpTKckAShwGT2wMPZQ1I/juq5QcU0D7A4DJzh+/co7EZNvViCtj9GpoyTep
S4j2DakqYAY/HPwC7fKsinstISoe/puTbCpjQ2Er601HTEjahOLYEHh0zwAEL5z9
pZwf62JUYub+WVynDxt3rp9L1F1TGdF6tHsiy+B+ckGUnVpnZ16x2ePmaWJVwQBB
1XA7jm71vm6Nol/Kq3c1rgzUUf+eI/7C1wIxeE0gon0xCx/vjCnCdzyKV6kWfCPv
csz2VK/H0XJyXPirbLHRb50RwNGF/7DauS8FJ3F+sSPH6oXD2CZlzWFlq24pu5Re
/9a67KLjtag2TWfurwuiYwRLxR3goDvuTI36pReE5bcE0WwIEJXlOK/3s7FY9WXG
UvKK4KrsJvZBteY3gzP5A6DUL8xLbadI//RHK9PHZviLVt28WNAKbEKb90LZTm1d
B/CzJ8FXU4iC0wPoYuIj9Zau6XuJ2HZTrCjfKh+y/6eVPPLrIf/Ss/qRlRVuYs79
prWe8ZT0VnE0sFdEPPBjG5+q/WqG5KRb0Fx1T9S7RkO27kH0b7wdn8ppt7foeR6e
p9YHJROPW42aY0wUeiYeMd67JRNsCl+hYVWrY900TqOVKk7Db11V7tS3XH9XBKzH
nSOBKGjJW9zCBOVH+qcC4GguciRaNo3LRoYyxUd8YeaaDn0YeN01b+unWYxBScPT
do+oUpTKMcD8k5X6x058txqD2c9Kcd07X+SWXC5h/fCDsg23FolPxF85+0F+zwZ4
mTq0SmFRUYQduK98H4vz4J1O+GLduyMTCICTsEpf64QFDslRjABR8VSnqMwDKj1T
va0wXs9A97heent2FQ489udW7JTFuMviLdW2Tfl5WyKaMMgUlFH24+pBvQf2o15S
s6qfiL5MkbmYtlqPrWGTsK5Js1/B/J1ogdSPLzx8Vy61e34l1wjw518+fja6qgPz
tXI/oGeR6d/vvvaZKBXxsJgtSn8OG+qFUgvs0SwzU7wOSBtKgW74FwPVyLx+XpwG
2lNjEAZr697hVRRJZy9IT3eNGfmfCbMEUG9AFsAPAwl15Cy0o8mFd6aNk60r8Zvm
Veak6W1zOxBcEJlFiMv6ivZfHQu1yoc9rJI/G56LkNue/qsiG5yHBG0znar+kwG8
06DUcY1uPJmN5Y55/S6ssxfPt6YbWQ3HKCz8ln98Jo1/lyu/NQUebsj2Dbjhwzaw
YV23nNpMpie8VcHXV/6vP8/891FLOIkKAv2HMfVwXvwim3cPk9hQEAUEe9BE1XTF
Xk9NO3vSj5x9oXCMG4y+stENmhB52yd7/sHREPhTKk63fGhn3HX6uNJaBiW6q1Ew
XWN+NH2m9b2M5Vg5mgC1cKQ4dVFZewrIFLjdL4zsrUPfd4U6xAnv6hpF0RcIppur
9d2gpNf0qXVoEhiEcEMhkHgYWaMX3Zy6y++fWES0K0wXyRX2nCLRUelgkH6ik3XQ
TX34DIEluEubkybm9I+WHHlBwtrdiZfmadZiRNP3hJRon/UG2L7SuiEqA4DoR5Sz
aco5331/ZgTj0LksY3f5Kl1D5jjCwFZObKWG5M0B+yBhMbAeUISruFB7CJ3AuhZF
pSyBPHOFiU2ME0VG40Ozoj43cKj/VrAPCsXD5IqRjPOivFE9tbnRCYCDnoP2yD7+
YK0nmzoyPEJuLh0p1iDRXe2i8gtN7gp+iUaq9hmyfGA817+V6YqW2OrqnpZhy/vW
J0mpOHonVcGgEG0J6c/SDM0ZBS2rvxZk+7KNAokgOBTZUR8PxzbMgYzQ/S2prThG
tCrFzimhmswCMvpn7boH9e+u1P2pEyFh8B6XWjeit2WCd3yvXuZePZA6d9BhDECQ
kIBZVbF79Ir5f9W/aftm/aH2C3sOK0Z5eR4s3G0cUkCygEuyCch2SHz/ybBM9zVT
kQ9A37cDaoMoGrZUr+8QAEnaE4LQliNTPnc6W7v07ouNCUu23xcQoc5j6VRHVHAl
CKGnbf+yRIC4GLrkZWqjsyOZ5R4f8ygq+TUcx84Oe2gE9PdBh5sYgkN8CXNxr2a0
3pm9m6Ypj0cPwgBB3xPr9p8NVh9flpIEpfNBO2kUuiwLAiFWjBFaTdeakKJu5dh2
22FTRcTiO5CADF0/DfeYDg5CT/Aq6PkBeYlgMglF1Rup98vOMnSRcdB/FhrsV1yv
r63Wrnu1RLqnZA7/jEeOIMh3RF8B74G8QyHoVdIapga4dDndEfomHnPWpbeJsk0c
eo83GKCpjSTRuYGtE6aNU0wmj3KoqbJsN7oMVKoPCEj53ezpb3dPwWT/hugqBZBV
ByFfVA+Bsx5YOQbRHo1in3tH80mWAk+h2iiKUun9ysLmWJdeE+VPlaZ7jOnGBAJ0
1bO3TCE4haKPHZSox8YtazlQPnLpKbwa9JBxDEDnDjlyzivmuu6Gw1lHsQrrk2Uq
ynbLmb8UZGXUZYlB8w/z5lNgvqW8T28zIK4LphaYpQxoxX6T0fUmDF9bOVCxDHI/
c87mBuHf2WE4OGvelUdya6muRWaCBQDV1NMAywk8RFpQ8VwKXZLGc4ffh78a3OBI
uSqhg+NMg6ShLUyoeiXmqaKtNTFTlSPhVxs68iopGcYIfGT2ZCBfhtI03Gv0tJxy
u04KKzdkPHq2Gm3zzw5jSjk25NNDnFhnELs3imZCUCAFKJt8CHaVTPO/6tg/NBON
MeZmvguNd71sK9YObI7d1SamJvfv3haESFKb1e0aysbsq0aomYBbNrn7BwytWwJm
pW5zrBOVwY+cLpUcfJpK7dpgB7Y2qB7GJ1LeS8kOEM6e5WCDIs0RlpaKLZmRJAh6
dicmuyioORGxgm8W+vVzZx7VKiycdOexAevXx8aupp4Khny4GhCxi3H+XI6pNPNG
kyoQAGUgp4OVuIFg5iBlBgjwTP97mZ6vN4iU7EvGmLuiDAo7hER0o7TGAi1ykfiR
fSalE2CIsDFNNQzla2cUt5mtAjRMtycVx5DfeMCYsjoxmdcjCrBJpRXUrE6MqXxl
pI6YSledV5XqXgVbkcXdd7Lmua7UsmdjGk7hyRl3VDSmtFDmEd7dEFnhP1+zBy3f
BFOPgskiMTmfL+FmxsgX4uhr8jkLSosxfEeRehgqV1d+FruF3hG1zE+VRvWwjr3r
qeb+yt75UHKtpwI+PqzK/uBriKiqtvbeu3sKzrQy2k15yHmixpu0CfrcQB41s6c0
vnUAxgoXvR4iKUCUcp38zixk2Uud2xJFdgPKf0VNM42RK2Dr3cb2hA1Zb2BptaQI
QNCaKH2q8M8x/y/YGWzXEXfqFg8N9Uy8mUXHETB7KXmVK/seCJ1eJ7Mv32IV3MZO
8faYE+xRngCy159X4IrJffSVWtJr8FwpuNi96Z1v9/zilfW8vHKLwcO4JYMTdOpw
68Wd4/stEOp4dRRIO4ekWL5NncayJba7LDimX3Zk23bf0HDcXHtFDF638ywxU8Ba
My3drKcg7Hr8SMa7MRB1ac1BBRRSgnzaS4SbST7AnIGCrpQZmot3tW8w3ae0+XlH
qfww/4qKQ3ROUagZAiHDCabA7Efm0+kgejQzJdA/fvkcft+2/bd5x637zNr4D8Zm
R7EDymd6CD/VGjGcfe1EVObbyiLKA0U0kz5tzwMV+h6g21m0N3seBSnLWxxH72sW
E+MYVahcuww712HV7rWm4izDiL0U8P2DQ9McNwFNni9r5fB2DCUPbPxLLllyLK4R
luxiGWGlo2g8Ggw96XWWbvamV0JL7NDLrCxPvVC112a1uSZpczqxIRhXSDnlz+KI
xkGZwUK7iIGZpno8VqYv1cs/GNZbn3JsYWr2ON6iAgbvxvit1WzqJbTegUkJIDI4
bGeIdGlG2+CBGe7aJmTY+DdcMLzy0Ps4zUAPNjQ335Ue6texaCjW0bTyklLjhaW0
tvVxa5a/AkaSe6+6LoxOJOx27oN0CmqAdSireomW0yHF6kWTxsLsH1Y4P0Acej3y
2mhzq/GP326AcCRJGxNiMDt6t4b80Ns2l0sikvQzeGcuB0te7YssNYu2pjUaUhVe
EvBB6R481PZWM6gauYB00bZOdXFolo0TJyLKqrqarUuUYerC0KVR5P3qvYbv9wLD
GKfI6GSgMehUYnAnY5wj1t1giAP4POMgNJrOm903CaKdiwsU7X4G3JXfASVbGo66
iIuJAadYP8cvSmd82hmwlb+2hhHdS3F2v6jTjVc9+ssOKa4GGREl9f9D0wTooj6a
G+tkWI8OUphxfomw9gsx7nitwoyMuueOfHBHtYXlF0e9DJzih92oWi1N4k1h17oy
xpHaiZHVjlUAEADrNfirzBActY/jO+T0HCjmMeod1fkZuBCdKYgRnk/Pip+Phgu6
OIat4hJmvpuLx3mcwi7I0qzG4bq5Kt5aT6YLhW8bgX27JuunfJjsPDChduVJk21f
8a81IFW4RfxSVV3y4t+sWsK+whGGT6GsY8rFTIEV9ZxF5Kd9XK8nMP6hfvO5Es4m
UlsSiFivPM9YerQfH1sCMgyHEqHWYnmC0/BxmBiyVTd2JGT02e8t53hApcOrQMIq
ML4T6It72R37PzeUx9L+WaJYKdmZMJf1W5RPhx/0hF2KYIsrP6dHsW0VzpBFCXTv
bMQvyX9LjHKbfYI+6P2+47wg7aqYasI5NaoMw5xgJXM3iDRibtECxlA9toO7TLCb
M8CqRkEFSBWf8HPpb0DAP37eAkEOZLtuUwDeHOhe3cx5uwtqL9mKm8+5vgg3hCMi
ounSO5nweaB/vFHnGdDkQ1M/QdHkTe9MzJnnvqhek2Qy9qQVNuqwc1XQ8D6feq4V
I5pczHqKWpy0baSNa6ToBjG9N/10exswkik9RnTzQEkea7uGQ4gDCcQ4lEqBwKaK
DIuTWGjq4VVfGHHDC47gqmhy6dmeDsy9w/A20E6ud1lhi0y+wZIG7CDvGwMZcWiA
hVTHewGw3PpFX3nKJe8QiD0luWG8U54FWo5VtG97+ltJUzp1DJ9wBcAa+jhbnGE5
iphVkuBs5oYaX6UUMztxp7BUyasbvvMfJArgqzedLGWwcdNE5QLhfiyFfaqjnBwW
gOzMBH2/hbw7D93+GmIeMNZ2wqk1awkN+oRnGHOnRQHBemIwKoxuJnPuAdf6qKh+
nMA43PyIf4WmA0ZSS4UO61/gWQWQZ0CiSIAlpSzXsq/dcpU1xS/8ODxqj6xBTp8R
6LFaqK1zkxcUKjOukJxGJQQbI/MCLeTsU2p5RUrjfgdbOOTl8ZwdpImV6wTNV0Qk
HJ1sDwOnI+Lb2xrpfHjGkRGL7987gu+JmvdeofRlPG1uUUEvBYgYeKUV5PmU+WDb
zFre00/jkeTVg9/dF4aN6Zhnny10FsZYX86WElsNVBA7U2bn+1jLj/sr2f6FmI6z
n0+cuJf5SxqGCfTfqRqN3YE/aW2+gA7Rep8szzSs01hUktVeh0PO/KxxgB1nKE5g
Jv82VdEUBOri8Bx17k6vv6QPuq66yG3GvdTGhQ+Cv8Td0mv7m+xwrMDa4ciC7Hv4
S4MkE0ENcsmWJnN/Cm/AVH0Co0L22r6RhPfkvChFTEMUogbiJfU9yY8tOi/2dBHl
ukAtwPP+09rpeIhb2yyqDTs/ycEVP9rIsEli2DzU0qk1X8V2NzZKGvhnN28yB8ls
8rRmIABCt2gUkl4nwkSRLkAGntzGgzKKsZshfEK2QJNKj+AuUbA6XKOmzkvVHZfb
sg3xM8Azqdg1doi99E4x1vk6lgsB3b+FW1FfKIGD+h9A6iKaw3G9J5ZOCvIbH/6J
PT6z78Cg+tSFvJEetXjTQ2/gxN6OcvbsmGHnQQiCPxgTrSxla0h9GQ5KS5lAr4fj
4FVuGiGf9L3myp6XMImF9cqIOtetJoG0O+MEAQcvQ44tbFnjravMNPi24kr7THSF
hMQwCXeCt1qDIIzfFv68QC5FLsam0P4Z9zUJuQZaCAFx0nS/c/7ndH7dYstCSYqv
/V4Wx913IDPeMYVXit9EP4dw25KeGp9NWlVkIQWlFg5x69T9CFRqWyaJZHJSS0L5
hOUCb/veWjOV2wS2ckkgdw7Z4ENiP2tcxiSah6YiAq6qJAcXlV0vkoGc0GtgtGfA
BvIJ+f5GCzyap8+ymegHRdC+IPOaNa3fBdq8UqQuB8k9eS43GknjsFO3j24DY/M2
gGupA3fkBMTTvsqRp+sckEEu/TBT4n4EXAo7+rcN+7FoVqcWv6yUP1gQlM8jYGbZ
NjQRSH2a84LfMJOFKFa7vf1aaR81VQSpmqiKnTjl2DkLpnwl/B7RaC6Fh1zkwbdA
FqcrznH9jNnH0L8++9X46ZkJ4UaTd71qhprnWlRYCBcBIgw5a8zan/zj5vcsQIEs
xmFnhhI8gOKwqURUYT8Zpj3WJAXO0+OJ22Ix3aH2Seu5/p/Dlfy1bG9LTRDYu7sX
XEPBdf7dcWOp9m+RZmF32b22iwB0ajYHtplNDzKBYCTG5xUEQam/3vE1HrbbX34X
fy/RvxbnIgDqSTF7zqvPnkz2uflDT9Xxs245gnsomz0gXPu5f3UNd7sXbOEITBzK
KuJ00+aZpizWnR7gkz9tgcKVyFOIOjMoGkRQuCFiWjC0Rf1+US1qR5ICiO11D5fz
EwKWTjcGVzVtE+CODfQ2l18WmUv3IdzqFWPga+Jzky4FgO1J89cZ/QDVIYYg4qRU
ikZR9NOpLVPLo2RsGTR9tVVsed9/87YQbLEyYDZ/+D2ZWqkmWjUYpeXTdkar42bw
LOw/nqK4m2942AD4g7QFaEsh6rxt/Lp5Y/0m+3Y1uQsMO9iIRxP1lQudpLluiH0I
sCWTyexB2lo1JnVr1wrSNTl6uk/W/HeD8f1EvsKk9mlFgxofR3Ip3bS3KMhY2LEF
M8srN/DxKywCs3ooLotn094Yh4HxMIc/2vHQsL0CIEwqI9W9/XdqjB/3xjfIrmYp
9tCtvdyRj022JQGSFOLWd+9b8l5+qZumZCc+b6ZOV+xI52GrYqPlME+d3iv498nP
8D0eMIlNQ5haynWigpEybi03hBjDYO8Z980BgwrUpJUX5EWBhJVSnDd9QlclkM8F
uhJZzPHRwleBS/HMbJcv/4XkjuVUcloji+PGf8zWGa2sOCBcSpMJrswA3+FNO2Gh
ylDxA8oUB6bCSfuV68EzHvXu2+T5VT/46w6sQ+goqasMa9W4ezDIo9sv6+zGPab0
D1/yrlJQIyLOyS752ClF9ZKBX26z4gIcS0dAqhHzvJv4kfwi8jf+Wsrd630HfeXx
T+cCjXHNSGpXH3/+U5NXw/S7pIAzGgc8N7AAZ4lB7nBXvPdXmvAkr7fdWiezVTId
N8r6XqRhGL0Sv/iA402+Zy429NvgG6W9uRhdNsEJsjSQPECGR/EP0MP1UKWGYgPI
99seTSI5+eTJwR/UxCvwqIpUQaQdkeL41j+r6IqsngR1+QvimYTBnailim9JGFVf
cS78td1SMKH2GAvl22fOydxCArrv/i8wEMMSTXK1sqaZlZ3/BfVxIdZ3qCEpTUUW
OEGpz488shYIEtxwIgRUsZCNUlokkUzaFyfQRDVHK9Xew0a8UzdiEw8W36WHN9Rw
N456v1UjxeLkdHzgvWmJH5N/+JYeuVAX4HRviHVLcRkNhppaVvqzzWDGpscC9l59
D6o+Mt62nlNQSB6FU/p95XEE14jSP1anubOFhFkUHIZ+pn8NYvMH4hToii+Fl/5S
bx8CYPQNXkuTBky4tivFHtcCXxTrzR2zR8tKe9fjgK9Dp+mtm595at0YjmxOqIxZ
13bFMYMC5598xCE2gHQDDBYwqhdSVE+EcAPkItSpv0bKM+EwIl8nocdztv35sPgw
GlcMvrL2EV6ubpv9BQXqs/x2DoM5qemLoRXb2U9WJzzJNUSHhztgjYMJlvP9iORW
dB9lP4r7AftLBUyQhUfH7pTpp2T8cvo/miOr6hO2JqhZLrpqiEHajYIdqVoyW/Ao
Tr97EdWo2RfMTv3zw+g9H6vhj2yErPgaa8G84ARnH/EgK5bXmqS5Y3nWzn5yOXyX
Fce6pqKtMmFeYcs/XMb78DpvxgHZJ4xSuQO2gWu+kf0bsA2uTrXD3LrshGBlRLVe
D3Xct2huLZK85linoa+uNyD7YIysV7y1DBnL7CLmM64h31BH98Jj5+poxxntBRIO
W7jEd2YOqDigdY8rG/nclOLTJthU3rto2VlG/ROLixe4uU5rf/WDrGYgawTdaKzg
Jku6tmqiHecoFMM26YN1V/r6G/04uCcigj3cXXYECW9bm56p7ahohjNNYP3hT2oH
L/LowZ7Uqvz8Hsx7cFQDl3khntPVMxhYCOl4FTcaGcnh0ONRgZtwXvhMSjddigC5
WcY7CWApETJxTBstvZsEvKyLXqy8dOFulhj1peETlN2zoNreaZKpxBvTUDB+UJNN
or4lNHySlQAY9OiwNMqhsDfmpkofXcf2y44U0EBsa25TXGnDeA3F3GFQVMaOSjBd
lgmIsuL0k2HjZyKkiWSdGegxbzz9QvnSkYBvC9gKalEk2YOfRzbFSNX2wLajfbGI
tebnKi0kdNtzBm7iNjjW3pidBv+at84Wk+FJ/n2oR4hnUNfhXqvGFkImwpo23FdJ
7oIaUdhanjdQHuEwl9xcQRiiC1mvfIt5PRTCq772rqubGLGbPdAvUZEfDRckTo9D
6STMjcst/FQF/qz+Jmn9Bt1tlTmEURSDYFSoEl4ZKN7fiQ71TPzJQcNGX3ON+J1m
nO4NoFkv18zBo2qXMdT/6eKsk4+CvirC93r2nrzOqTP7pMPPYi4zfVqXw4LF6c4o
tnibEwqirv826LitMM6Kcgj6zlWMV4nLZclZaQxCAeGXmyC+VZ16TLgB4iklBqfS
mG0gNRmQuDa13CNavOBZnvIWAv5+BznxM1PLZcYEfbyIeLjZKid78LXuYMaldGgm
3edhMgFHNtzjGGn+IxmUTpTo2cariNPKYUrfl33LaGCAMeYlfjnk6+bMsYvCd4Jr
XPhL7K45Bf5sUoGczH9UEubsgl3EfPj+wLk6H1cdMH0Ug+tl4I5Z4EzDACLN2uYq
MSdm6eoyp5ws6Yu+wRHrQZWghYsMmXTrH8loGOAc2U/thBwL+TNp8cCCY3/50yAE
N8kBvjsoXR35SgCLXtf7lc+fitP/DY4g3T4YH8QWwfwZ4EreDYi4pMefop4hOeQc
wkj7h5upFCVD5qtkXfEp8chy1RhzibYvbTl3ZDVK2ZLLX+IW+uurBg1jlfrXx9H7
+mPEbFvCa6KXWppIm9vEIhVpfBoAVLqjNHIvOy0NnCup/m8O0zHO2KExKM9YbPZG
9sIauk6sE49FeRTXn3KPzKFNTqNzmGpGgGoKGXCF94Qlz/j4xw7I06jYYLMckFHX
Vyf7qVuFxgyL8Vv+cnQOoVhLs3zLBNqMAAen0ZINxV+TOGV27nU+rDChrRTZnlAF
ogMJn933SVFeqw1uW0kzlW3w6k2hIEMVi/O6INuHYJCigEbu3IHWAmsBzUNT1I2Z
siIQeaJyCYkIKTGvOyew3ysBSe/hz+Wkw4AEfZRvQWlWfe4LuCc0WtWfhtzoe9Kb
64Hq37xpap09pPB/w78BWqFmScPvA4l/H8cLMfHE5Ek+ijvqENQmiOljXV7cT8Ew
ilT6xV6Bz3cdEKSRhJbFq6GSITpsQeJvK8ySRJeGSJyr0BpOqZXnMdBsXPs5Vm4k
kyvG0pVz1Y88Wih5Qzd3I4y9Q4+uihteoQr/KOoqHb/MeeN6OisleNuXMlKJF4Jn
1T33g60wwXcJiPBqSze6opeZpqmk/GsABI10VUC0qgYQjkM/zzYpHXx39FtPd8ga
nKKKVfPtfUtIJJyaZTyvMZirQvma26dnxsIn5ap6UkLY1oHrtEVfTDiZ1uZKIsLB
w0Tohz3gD0Zhbj0soKv64vP+/j/Orc2DGkhN+XpDYadIdJ9kBPVbG1D2QCls1G/K
DDbvusKK4qxCVZsaIFUDHdVBFrA+gsIzKBru0Kwp2Z1D5pnQxddCvsrhJlRhjTEo
ufyIIDElwJBpV2Ij6/q8RnGfLRX9qBA4QsYGNiu/2FLNRlruJRkMDLxQ6P3CMymS
Kn3lxXGM0BP5Ua/OsWG1ZT0vqZ4nzU/F1BhB9r1HZKjuZ8AhqKp60Q9+J0jChWJj
WM4Ew51eUK1aZGEinmycyd0Qg39BkEp0ol5gLbzNvK3icmLpaLNEnd7B/JNpdjgb
YokPiGhNWKjOkv8Xht1TgTXBsy++rYG3T/V7F1uWFG7v4rneeeNDVB+0/ryhpJev
wlpYm8Dk715/yFoP0FTkiDaSa6WxJbkf6RwEDVYOfGKcqI9CfcKxyNB0pOZR0kr5
6mVc+OjgOqyw7oHvLSNVOEf8PGVmfUUa2OT7vqNSt0DCkM4LdoEW2yy8HAMtFQHb
kai/yhmIyFGJBgmedu7H4c6Y1JraeMF5YbUR+ShDe0Jy8I0SHnTcCZCvJHeVT4TC
AqBQJoOWcCXwCGlbI4ew4B6AsfvAiZS3tEagT9XW+64V5jGu8uAiqwKLBQ9lhWUB
WE7q1xj3iN8F7sofuY8BssNzImZIUBL636TQ4oFxRRH0idzyKs+/khEPothYDO4e
b/QV6dubMDTkYOELd2wHSpOZNTjCa6yTMFGEJKI4O1dWe9TjkD/uCf4zjRIsDx+O
eXxC9XjgApQNpzz9+JC5oQVYDhZo2dxm/287Ro0HjmbHNIlb0hF7R2/8x0HQwo4W
/w1MfYWzBzlcCGIx07fIB2lucGZDHHIrTCdjLUzcVhOkmPckKmDt8YJGoVLt+Y5e
rlnCJkQin5oKVarj6EdlYoeWEY2vyuEYMMP5YY3KQhxxPr0i46ecqp2UORIMdRqX
GVcr0KIDXgT0hMP2da+DXQLmx8ZPE7K/gtt5aYxCcZpY8nOo9Nch3aXnsKRIoQsT
NKGg7W1Wh99PX8e+SHLY5/O9FybDAzWWNu/g4/LXYDVWMHT8ouODUy+LsvHldJCs
iI/PTtEmaqagLy0D3BpBF2EVvU/0cr01mqp68gFPhBXUtiqQG/ZCXv2RKwc0gIu1
udlGInUZ2QTLeWLlORI1xcagcahUd8tB4TodgWtkq0a/Xuyy+upWXTo8xzvwbqhZ
V4dpzlZMvmTxAhsnh4xN+uLzmqm0LbCmhUd+x1iYRXXKxuj3WGViAUa3KSZ9tDEE
CyCK1hEcnorj3WrzbCJr3Mct/ReZvF2tAk6kzXzFMt4asj/FOkxTg/a1cOoCDPxi
HPz3LOcwFFrzIaCnwbzoVBNQwoPEab8ObVa09BQAk4xaw9NJPuTUiFEnLK/7jrAT
aDk7uXsPThpPmJtNrxqZRywfyJAx0vEg46RcAaIVBuXG94V7TltDfY5/d9xWMUjB
g3mqs+Shx/hVbH3x7FIQ/T5n7B11hZP71iw2tgallNX6DkIluvtlgIx6AFJ9uJOq
kAizEBAzB0vbIpqJlUmHlAEE1lMfUW0na7b/fOOCLEYWXQZH7CktyPT7qqSpbtCx
xdCqA5ISfOiY+3iIOsznBelVFbBU2PsZDc1pXrdpWiTcLci071H2d1esV0n5sebL
9SjOzFcvWWfaDYM8BTYoWoFXu54jHhIbZSt9oRcunjxksztpCA735RhAecMQBeL4
L2yX5d7kaa0hUu1X/5go5/t/yncdZPLKtWitCKHp1Sw4KldVffqI4l3MlEbcZq/b
nHnxBAAsFZXl25LkbYF5xgG+ZqKHdKU61AuTYKBYOaEjdbKeXZv5NOsMsatB0qFh
4SITlrHP5SkHJkpQ8UdKJah+Q1b7pLVWDlPme7VRj22TLxy1zL0/MJtrTThbF1ka
XkDe6rcJNnMvdinMSLoXJp/WgE/dNvbdKWrT9N1/pGPtaowRwQSibDh1pS3q071n
9Q9P8r/kTDOshE97oXyJUqRdxWHHRhQtLNm0LftfFMgdR233OH7wXiJzDeGf5utb
n9nB1vZT0bGpCs9/7drsSzk+KODWiEd98W1ril42PxMOTGCl7iiY1fW/IPzty0j1
Ok9+MdrNx49mIAeV26Tun1TqG4Fif3v8B7ibztfwyGWCdi3FLBMHkp6vVGPHDXRm
fk01BsJ9mWmCnAUAmnh4VcknLymX2woNZvNqy6qHCVsYJkG3fJO3oGO265EbdL4C
F721IW4biIxdesVpUptNMpMHpv3NvJdYBnuNyny3DM+pdp4scyLl7idFIeHWqEgc
pxUZ+nlBeKlfPtwgOq0duWLMKXZG8s8hRPzExdCQlMkwIAKgQIImNpEIVh9OHgX/
2rRfEnU+ojJMLoV5niFTz5WGmUpWFEyVNhPdbAPOgyTcs7aqL1N0PhqFHX9JfpZO
hxFqd6rz2uf4NG4gs82o8iAWPSoYmMcYBLnmuFGIo/TScZ2p75aY/BiKfGcXlkyW
4WqROulQtB/n7GK2x0eekSDMu2FResjgZNiQlUDrDWrVZXx7mY40lnd6uBZ+K3iw
44zrKKzdqOHlKZHdRoIacylMNZjcUPMMG7smU8CpLUn/E4mF5wIDR4XYWOmC6I5J
qhIo5ddJ/lnIR3681q+g28/+VWf/mkyk5yBRMScWttwypujMMXYyWWoSBrIsGT2X
zCqbAfAJRpHOtmaEu7P113n//QFwOXaya0h7dhEXnf2gGutUjjIkB374NSbcEg0f
lA8W78W39NJO15bChm8mCu2ahVoaBMS8tJjcT5clEUu9XMKP+4brkGHDH9ip79HG
qbVTNIL7QoPSdplHkXbmmZtpq3bgWXZhkx9p1JeLC/g+rdC2eHDrClq8U7eu3VdZ
65RulIOcIND0MPkoJDVPcRylnHa3/xAWY5A6Zcfn8lm5uPFTOrFyrCUpz7yUR8MT
41RW2JwCVpnTHZ8c6KHlGySeo7PcsK5NU3A6SV9IrJkhxna+BHyQyvDnFl5GiHAR
+TgY6SuUoAXh+J1gEwITUJcyCwwxVF0gQudjudrfgy2uoVo6Pc1/F+c7VOawpXBS
3Me4F0c5Ki2iruEkbk4GIa3Vu8LtYzrtBVcGvJ56iiev174mwQENIhqD+5Xeoz/L
bobqhj/v+eER0e3q1B4BPuphtif2yrRe5o2tL1LzAsoLctylDvqm3xr1oTrXk4W0
X5Ssp8eEuQVBOyxr7nKmVlDyHx5UUE2HoDgPj8hcIi2FsFHCCQcMQ3QwXFJREXh3
olykTrh24OIz39Omk51G/eTyfCJUudot4GSiakdfVGkWD/BHfyUwPOpurEpiwsN5
vqmSGSLVJ/OZS0C9xueEId7lim6xqBcygZLgolQOgDu4LEKxQEKnEJCcnC6OoeDe
va/DzI1dSYVMwkTcETrerI+ZvEp9+xUC8j+U0Dyu6qoP74jdgMcnRXm3ri3tKkrd
01G6A60ur9ovPRhw93uxo7PF2VJU9sS2ASKMn3I58xrHMaTXGZ/xIVh3fEgAPLEF
VLM+UtYwQ9MvWQVLDCvxCuHsRsCq2RtjSwwLgvd1HPAIFL/bVUGZO/AdJL2yOs4Z
Hx2YaUHJhtfg9PJVDWc1wJQXEtJPn7XTX+t7/GZS1o/xGf6Ff6UfeplXbOMzzE60
e+LkNqGMnhP65fjUtrkndEOCz/2FJSbGNVovBDF+XJSD4zc4Gaf9JD7db3+MNVu9
NGtoIVJJNs2K4zeYrdejIUxPC0ZPs9aVD6o0qNU4tsKWMaK1ZfVfalecAiAB6ROq
yvMt4lPQ66sDKIIII1QDlAf9C4QeTCAZnqjlEa6KKxxUBzNLajZqXEmzELBjr7YU
MXtfCTTiUHhTLt49aPHQ+O2YnoRdUiFCNpG2RlUSGjiYqlRTZIleT4MfNKEJjOMn
sut4twkGpST8AwK3d0VpmLKNgWGu5ag9sMECamK5KugN5yIeuPMiC5ym0kgvY04K
yJwaXsA0T7NMfc1vjg91WwAvEud59u3rZ1g1oJJDSOGTuZWaOzowopBNvA1+28LB
9ZLqMnPiHHZrhkq04hIqyG9bFDodpoKla7OkJRCI32UDEAYM1kb06v5RZUc3pMmz
twdoxCMa10wAohCbf//c3OKHuMNTDqhZ2RhjkayEOnhIU7smOE+PtbQACaTOvDkO
FN23X+lGKGJU/5BKE6HUxKF6JpIdDco8j9aDdgDvo7poUf31r6Y09lQitlEVAvL+
ZXSXvmx7usNnTWkwV9AAc5qX76HR3qHR4fwdqfng5mOIWynHiRZcbDl3bJKVpSpM
VdNUhD7OcygPv4rpDuqfOAN+P/sK5hOHmOBlAZiyfpQSM0CwVRq42ct8wkmSL/Zy
22pFhUwo0Lr35eNyXxwgpaUf6MwL7vzwbdaTlAJqTIihAaoaka6Mk4xXm9fFoYVF
HbBUX7P4If8A/qEmYmHxUNKjn2OPqUhNYTvZWGB+yVKdez2Kq3B/2E3qyIJBy2au
G5kO9HGDtLAAsjZ/2smGTX3zdXsfE7G/5h/U4NyK/0y9+6WrDtPzmtaNM0Yg+3VX
kETJz78GWot80m5BgPi8fLpX1vbRaY5Q74pR9ln7i3z3APw8palEaNAhaMAX3H3k
JA/BU2SFrJXmIkSzomDgdbXYrqSVxTv15s8R902ycyK6OYmtgi9VUvL77dm0WlEu
BTxJfxIXlf20An9EZ0VBjv7vAd/6M/4Sq4doE+qF0SLU5ct6h1mbb/IaPdSbbtG1
7tWif4v3MBTeBlPXp7tDfNwymWhnap0bORM/cmtqQeSnvOqx94g18kgRlmEUU6s1
T9/aXe6LMROZuMNMRUd7h12nyA/EfI1VurguNxuAFzaVMU1tP6Eakh65i9mtgM1T
Sx4pPN3L7mjVbUcaz5NHJCQC8Y0jd+Op25cntE/ZE7bZQe/o0w+r+2KbVOxZ64Mx
dHYe+2JEsNgjqYPXlYGITy9k2AOK0qNdnxm+RryEFFsJbzOikb1nznBu96yoUo9d
U3WhDYDlLTC7EixtBU8EKN1xsq6X/d6gGBZvqq/0JzWbVNTavlycOWWRPFr4xc9J
WBAUug/ZmcKEQzvpuPyyJGc2CUKT62mMFtUGLpuw4/arFvdUvtYcw9Jlwb7ChQBl
HvDo+sfIhyH8ge8sNgBwlR563fmX8SSK7+pLYt8eB1bzVIe6w1IGAZzswoAxYDI5
syS1Z1aNGYXQ/WMFWlnnMErYnVwhKVVOjEFm2V1c1JLFhnWhGZRH2XgaxYw744AF
U5+ZslqIyhqGbJ2FQGHwwHlbR8WDzTvaCaAk/Iw5nMRmrzL93fLSNfGdUoy5VosZ
idWrmxWlGoRxJyaXEe4jord68VK7MUWiqzkFqUbWOlxCPFc7utND+C1Ydf8bIBdJ
AO89lX01ziJ157lgbzoLQRDTflFxfg6ZAUA8SOvxEJZXRvkgtwO7fGqPtOe76Vo2
VwB2mQNAQQSxF8kmUnLBXlUYJF43fgNUQnQsjY7yd+7lCzkqs23TR3GWMplLWJmX
xbaFUhXs4YbW9xRi0t0HZ0wkAiXBl3dQtdfs6yYpT4yaxNX5wk0p9Yr60YZ8dG3w
qNB2Kbm0SP2tnDHupgestErR11/fMkLZh/DwZyEAFXOZftj6cFUClF9go2lSNlzt
B4dg1L0lq9+itj2jzADFfk9QK2k/AWhItdi280obNEl7A8LbIYxi7oH7oBQ+DvQv
H24tAANDgsXoqiDLZXR7IKo5SRvFJ7o7wcEzs8nLOtOF7Y7O9KsIdaqhXlhQY9qs
6E+TIBdLfFOzhBcXk4Us7jtg0HumL1MkGQfzUg0/nrc6zekn+08vwcCMLq7/Ei5Y
Iy4De4qqXnQiketG7NLc5S1zeDtghwCNJsD6mzvCvA0PllB00Xxdq6nGnWHerhvy
W9lZWn3J90lQVgw6U/Z0PfxjEVJ/3MRP19Vce32dzaWqxTA8qSKgsGd4j5+BMnbg
aoQHL2oa48n57/iMDQftMvMEHmpkbp4kGSDeipVbdtU0XLQwO+J4zrVXrhOnJA8H
ddiFzd7T3I7ATEYVBpWowG3KhxfqKDPPBACth5Dh4+yBfHh9yM87NFar+ojs28vI
/onRVxrMnKofsD4Z/JB3L33RiDSm8UfAcKale0pEFH2UlgVtpbrL/WP/K5bxlcuV
a/oLTooVYtxd7o0dtFAbG95Y83Pgbvj5YLJv4k6lnQ3DM2fcyHXKWc6RQQ4LZx52
aqTvSP3rDAdK3TqJzh+dDhNOjHbhoS0kuuM2XZSoszuH9/XLa2lsxBz/g2+04h6N
w8cUplTp2jRkA/kOvAdh4wIeC2S0WLqNhA8BoznH3QEuKtu+HQqoIUsCwi1lwkjc
fbu0zswuG/iOwb7SvGZU3cmpY3rNtDZb8c0ilOE4PnlYvvoVvQEF80WoE/W0y45e
BhIeoaQl7MFTUC8tkbzkfAphXsEOrzG18u4bGJ3zv6alqWopSF1i39fzEF58aOF5
rbCwmntzjwYodmokU20Y8IEVTvueOqXUfcTf8yB0Zet2bkJcUTPTj0lBDF2AHOnd
tsNIIvka9djDvtQlZcPoJNK8+BcDQF1NSGjoGGqd/l0CPqt6J41SsnV73wkuBteE
1Z8F39R7f7u3esCM1PWLCsvy0vo4JrYE2e1Ph3XiLW7+qGwUeM6Q4HdcsBy0KER8
lUZ+j8VCLMVaf7hcxN6o5LPUnVhZuykGzoB8QSWrayoHAlGXA3IYOYdEKJgIsgTh
l9Ewe6oGgwO8W4lSjAiI9DcATPFsjdNrt2dhaCOagqrzZy4+YuBIv68bl4dtHeZh
eGLImF8jMmqZ5voyFid6+d3Y9DMT9rpKD+g8kW4mhuTcQPuOSnKo7eSrbixgs1MQ
W/Q6fTGJxVF/T+sWSkOpxq1F20kcgTiFkyob8oj7UNUXFeFMirqqHt4Fuh6EeU2b
69w8b5VgU+5n9xh/FMX+/outJ5j91lOdx1WOtX8FxjQ3gyIJoBwLw03fVP8lyZ+N
ul6XHm+WVClOdXGh6+1EwvGClVCBem4nof2jWmd9zMU8KHSZ3CAZnX9eOAXhkMaX
Zs/HldnUWZ32vYHO4Eu06EclIoYa7G3Pj73HwNx+ob6Bapb1Cra9vAUmVPrcqKXq
9B26Il491G5U+ETBvl8RDCbekkRN+hBJkLpQF0+Ve7qXHY5XnXYP8c3P52dDRb3C
QRWOhh2hZTsrJywixW08JSYLTmlTKi/GDBYvjZXpPjqk3AwNZfn4/MueFz2wpghs
Mxbwk4YPzhFpnPNRhsMAAzeH9uIVrGdmpCvIBq/SByE7Msm1GJ44DaP/399DoN9e
C50UXC8KYFf9Xn8OilSZqZYmkCAB1RBFIz1ijyxK5c8SrmHqi4ndTPPK+s6d15TO
oaZmxFJV6IcjzFUCE4RkBDb2ClUWynDoEsOEun3G18clkydDNJSKKrSYbceNXEN9
3krsYsIysgQrr94qjJdtwY+ofwyxCOBmSfCKN8xrtPU2WSzG9hcMwGRerD+7WCxO
0FkRgDmmhmShJPuCo7HHAhjXMVwHKhwsInrtNNGhdoDS90SthPUm7hlZjjkE1Bp2
5VIjykwoRDk42bX/OvWqf4jDseFrvI8w2ch3k9zEPWiHjq56wCZfQ5wSCIzA2dCH
16nL1LU5U2XZ1rkSe+HdOKdKdrd9gIDLvBhRWtFCpKpnseFG8I9FCX1og9FNpM8J
Qydax6c13NFj18jBeFaIuUYvmQay0jzmSyRBfH0RSS8X3tXlczAirNeoOH98oL3A
J3cBPqnz9jgRoH2oYrAHD8Orr6L5RYRHK1V4OrgUrs/HPzMYBqd/+9u9eazs5Oe+
VHuqGUOk19KRTqgCqZpMX9o5X7BNZsUt+Yce/q41dxaclxpCHWkx4rsZT0FBXN/k
IbinPwGKLtMGMsXSm9omDbwPssnOYg34lxTDW4/distsP/vkb2vzZQqFRe2UTRez
NSW+XT9yb6f+QILOnjJP3l2+W8Zu0ShnacN6lqUF4yhvEsjdeKfMupxKm//R2n/G
DP12yT9l7Yis/rqVQ3DoZnWNB8+ziXHfbMEL3d3+BRDUNVWKfvbZGDpjl1V40Vxw
f+U80vj6dX7U9Vb1qVIk/3dpalTaYb6/sWVXDKB+2XIHiNDqgyx9DverMCO/9UrN
5Y2PPlY7s2048kx7Kh37LoaRKP/HHMhU/gD74584GpeEnST3gNIx7kn0U2cuo4qf
hoQpGiaQzY/9dwE/Ik6CPhO1QYkg9ff6Uiln4CpxJHwRYK6krObiLYJslXtJu9/p
9X8jsyAoNMZTPeNgLcS6RKuHSQzuyM2Sp6wkmWpDGmq3lKrW2JIE6FxygUwCL29N
1QiulatCdvfQMizNK5m0jOnL7a3nqtgNsujDSU9oMCeAMMMKhDaIra1u2moVC8DX
et4wp4u39MRc96sd6VkP53YUAhALZOmYzpyPTF46oMQwlxd3e6cFo4zsryF8YLqh
Q/2zoeqRbnV59+uitq0UNqXGsq6X2aHx6XSWOkxeOOnkcplTZXj7aY6Q8v2BIySX
3Wnme/4xwuxY4b6aftW6/17dFk78+yEY7pNzZ3HzcU60yYWNx4JGRh0LQQ3vkQa+
EsG9dlDWAKxxpAm+j7anpGsb4Zef+HrE1Zean6no4ibwnaQMaCeMIYpZYa48bVLY
W5Jzn3eFKtg+S7xVFOLoeP/KFgN4bBaMgQGCgMFcShcOUWCx+P72lWAmaQEiBD50
6mQ5EXuv8kh8/WpHWsZ2s5ceD947Zg+e2MzLY33/ddhOqbxxJncnYkLE+bW2UABV
gKTYIWbD83vH3ZvbNX1YIpYV03x02UeKmn5KdAuQkR6SjlfbpPPlo3Wc+Tlysxr7
SNrl0JNThwpEOMtCq9Eu8npwggPXo1+Fayk+GQqEvBNA1OwcodhBT1NTpwQRzMbv
94YaFT83LjGNM1dCV+Jdjtbc3ZhPQi5swLJlbSqbJCXpzAQzr6UhWcdAQ/Ck5WyZ
v8FKeXFiIoZJq1hqvil99MCnfDBIKeRNblV+ZbvO5mtO4nec7cLREqKhg3CGvE8i
3uZtcz+4zUWrWNCJh337nPeyWJpHrNHrlu/XrfCuIk0BVkinyOfxuRSZUpzZpaaI
lUy4R8Y/Riifr+vKzSabKucI2a7LrvjMQLhOTrvgkjlHgyu8UkZrD39u/rrs7kq4
YmjPYK2f6mbZ6QwzrTbP7aucw9GXutCn+XYpZ7Cj55WsQeZ+XPQhoSDdyUZUbRNz
lXiAJ/Umd8Bv40Y8qAKnucBViPPyokmiGW3akGXcF3QX4Sk5DSMjXAmLPL+RLp+h
g+y+kYCaDWwXYqlhoj6z6eAhhk91H29J0Xxl1eEDvhbiR6oZyvSXr3v8/QQoZ/8p
qJWup4FOHxcgMl4HVqzMCLFjPeLfo0L0t38FPtAjHdxSlIYF8cq7Yi56kj+cagRj
ggdYiFVCgwXISE/RjjhG5Vawk8vTBulKA2N20RONviJQpqTZ9aaYI5IdEptN6snA
Y4UjxaU+YmgQLaslSs6HaIWE6nXjMQAqwMzL3zI70+RybNQiVuAkc2CRqQDg+ihU
TBDjUmx65v5eWA3kgTa3VZP8g6VQ7Db3v+C414klbxyMsaCjmNSD4fsrL07HUzkV
znjVbWf2ipgFbHiOncREhfU81Cb6l869RU7HHdJBIpdpW9yuqxoEH4sd8Y0DGTaq
oeibp2pLN6/130Wsml4pqw8B0jpRTacNrTPl9jtA98gbCTALxIKOLpwnWI9KyX7w
2zaGGR41lDKtlVhap4Wfi6OmDcUMFmb5fZ9siLUtez0uIwZW7ouk84VXvVFnhNYu
7dkyp7x5eopO7exfHUfBxm9TyQo3DAdBn0EKYIeqNuJQIurU86KHK0s4PsAe0Scu
Hub7RaDtLCsCYBt16ZeVf/RFF15XpxmgusDqq1Efa8upty1fe9NXqwzkUeU77LBb
1dKXW2tdopOvlaPhSU4DYd+/cCsmuzeM1bIZpdjQ1VdNLnxvf+NCuQ2JKXMGMtiR
uPMjWch46hsVo5FbpnDWp7RVQRVnaaMTAyHu9d2ZIM4RW5vcv6Q82lVVpZusXUAi
1ORuS5mPGnGDn1Ozp4+JmucCRFPGjdl654qC9QUemEU326kb3QOxBOaWFUaJ706z
ttDbLxOsYeabem7jWcmgA/YBDSbVt5mZi/PsQV6ccvYWZXUlEgUuHvPSnf9NhRvX
WIdh+JSjRwjfLf8IK2yWt6lvSiAXi0uh3ZjqsxzhFevIK2g+dqJQyRlCnLrwlCQx
VVzWWfCF4ZCpFaW0SlLN0b2KRLaBY+duff8+HvyhVQdm+X4jPMxzXZL2EZOJc/re
h3q1WMsYoXwC2nSS7zNxJ7kKOIBMQi6eGDC7AkjUCE2sQvhqyOAoTHkV51d2hTWh
mmri6dXAC2xnAbxUETEim8k4pEijY71PUupg05uRwKJWmYhw3pB2HrDM74bEJIGh
cNX5uOzt15yfNct0YRyS2U34qFnz5k0ryHSDRiPwKjYhuFKkhHzDs2+YJnLeGh4M
qb1xSK2nobUkOJ9gH/pBlkoMQqx0Ruky1pPaRkFT5bHsZmJVdxaCENbxhD3+PQzF
h/lWVb3bLq82dy5TdVxqhxIADSJRT5FGKdHqivzRY4UQp4O6szb3FQjTNv3l4G8P
bw0tkQRi2sAUMtFVnvYtPhx8n7vMwQfDAgU31/xmiktVG9N3ifFiRYkYfNPCpQKO
0q306Wue8k8YsYhJYIEDpwztHS9VtPRAOZ39ovKy6HO/vMR3/ZSBZXG9ojPL5kzB
JdTaZ509gqcyWXmuQ0jxvt0FKWFf2epNA6aB/rmy8i/6FSlFmNCwY9bXkHvFXy1e
jq9QYYDEJiso/I92WPDhksgQ+SEkPLXUHcstET02FL0JvcumlXSuqboCyTVhNARf
n1/4v3Jo2gdedM2h+IYvNBT6qqrUpFV0B2PLWnA3fxvI9Nr5gJ9sfNtfLDOYmV9m
PRY8YtRhZCN4M53yfkR45BPMx4hLzgBCkc/4YGt/sLs9UU+d9yX0AtAqc7/VzYWK
EgwMMUvGLAbVLyy4GbCFX+8AL9/dtVdolEO5iIA7NgQvIBntU59YJKverixloZoX
okdAfp5W/7VPff6McD1n5b+kZWw1VW1Yr2p0HOsNKCrK6X75OJPvAtu6AQRzQFfH
Ge6FTLCH1szc4ZbUa2zIH/p8OY2g9YNB25P1OwlpENXDhPHuWO9HvJtsPqmm+B1c
O04tB4yRPB09k+Qh5NWsroxZbK5Qq1RzsNXniAi1X4zMRnk3iin5eBeWmlD7vXQJ
gZtvwXJdAc4428PQ7jsdYAxFmePzz12coWsH52+Q5ynNMWVQSXvVfogqagCzZRlx
4jYZH2ReblmbHFVHNHmU49u75zptxX/TYCizCaYN9XKDGKLWWixSl5XgzFQzpth0
dwFwVi2nyUB4ddJGyQFWzr2XQ4oYCJ4P09Bphp1YBS7l41ujVRuY09N6AzyVLey0
dtH2VbJ5YoMRfZ+r8MvTs98YFQG69BA4CGWUAX1nc+tqfyEmqcT2euxr0k683FIm
eOAGjZMLgz03TjqC/dvr9P+C8nwrNyCmQqcKSy4vj96C79x+ZQ+eUzJwd+I8Mt3o
zF0nTKs/25+UIseNvFkS1WovkYA+lrwAnfg/N4QGHU/4W6Bjr1eBpt6Mc5Tg84r5
WwzYNCznIdAPAkdk8rM6EmYcgXS6Z1Mo0JNYeMUHYutP77bZdv8ooj/QwJkS6KYO
jpDo/LOaX3dN5tiCnwmbRPnVOKMn3W4JBDGgie8JhX+kMQH8CjQr0iPvVUDGI6AE
wJ6EqZmG0saiwjgbCE38DFPL+JUjN4TeFGvTxirPkvMAsnO0Tl676768h2pVNH7E
U5XsKeg3kpzX3nWmYBXef6eAfF+swwSvXoc9cJd+KFC/TdMkhE7xaC80HLO2nl2c
S1O9urBVCoMURwrVE86h0c0aTUjKFsEsJzEyhRmzIydzts8HE05Id1SprdCKwsR8
KL4RBdgGVuS3zJHG8ypO5WRtJnyZOuE5HeJVHNX/r03iwjGlOxLjmXTonWl1P3j2
nbba/ODr9wEPoqth1jM/pxiNmt3QXoqg9VcubPJ3g1Lq3q5lFeHitwvLPBx7Q1EH
2ouQqmqxDb6fp/l4USwAvJGnOrC86q8WU5Yp58zzT3auWnEjcBdIbfNxmv1G2KzN
3nQ1tpYeOgEjp7ROF3OsecuglPZ3rG/3S72Gks5rGanWGq38ZZTriWpZFdk8+e0d
c/bQ34Taf0cCdxDZGGYkAayGpivCcX2TQirezM2Ccr+hb+eJFaBVjE9jlegyVYqD
Pj5hrIDtIhQrTsUK28+eGMY7tVOx5rNQd4CZjZKr2zmmUgYWMi9fL8bFl4r0WArA
fEECKzRkf5oUOqM58NiUbu+WX8yENS39AkYtERc/s/uEOZt5aeGURefPuk/ASeR3
1pK06a/+pmflX75uS66RpOBh1z4DDl8T55c2dv+da4diR/Ay6zsoyriIZoq1m1ng
WrK9exayNIQWER3siqldZ+TnhFnjuOzbzPrKNXMMgLSzHkKiYLrAfl5kXKc1djwf
HrqMbJG1Ur4AvQjL5XcMbNRpxplUul9upAa0HA2RAIqOTwsofCOhEMKSFDy32NFj
TF2Ot6O4D0Te9+O1GWtAOqbjW0IYE+ohgnIgxjBJYHIqVHVVnNBSMGl9qxx8zUnw
3JMfcJS9Ed8KdX7T4ztfuUL8WvEc2qI9EAI6ioQeKcNobOLVg77SOBluJv3nia8Y
158o1CiK72xieJKl5fU30FPraDZVXROhC+v30qQSQVhg3EgLoQVNcIbn2bgJ69dl
CfHtN+bVtOeLis5XSGtSGOg+Se58/J/lLlsrwG28qaJT1SZC/PUHc4LB4xdh2Qyk
QatJwS7oFKubnbIzEu5qcFgGn9l8saZWeiyHR1VLkZu6iQkGKRVMAq6UbbgbMaYs
y8AWEN3fbvKpYZXF3bQcHFD3nVrKhcCROeITTppBFF2VhtZajnxOoHKml/ui3uY+
VQnNpyQe2LQ070LVvUvHh0KNGfyPXBI+3nIgs1ZKGlYATrfIA1GsAibd3bwc/JSp
2rvQAi+rtKxU7cFE8yLHUl4luCy+wjiyUQk3E4MZnUYLcJHEkL5xGiZNBaHiHFxE
ccJqJC4tQwEYhgDtkP30URIGOzZ/EEb17zftjc+VGi354bRhqJZQYWkgEwF5JmF0
1IEHRXnGHp232pPpI0U7rjQ52tLG9/i6oUlQNLIxr2VNbA0fiGi/D7qixUI/n267
PNnFm9ZCwfmFim2MH6Z99zQMmHyKmpr+LYWr0T2EQrZYKIyFlx6w2QSoBFJ27yS5
Kw00kmHWoLVMfUZwP01u8FL8pKFxkuyh4VAwxtL2rXe80W89KvNDm4u+dTiu4dEY
BOTtVe4nB9XW1JxEkcYoNMW2T9cXOVN3kiASSLxuvPaVZ6HCmXvmzbms9+FjXRdQ
rgJ88nb790X3ivkmmg0aryS5Tz9pxF15g+4X6YyIri1f/iGgpXHaZoKAOIsd039t
GqH3IsPS9XXZZ4XdnPPdBo5IcOSRMZrh2dUtkRcKFYFZc5SYofGJDzDnWlBEqUbY
LIpe1c7FKMnm49zS/DxkYgVrPHs35i+c9x/IrfIxdMeZQ91s00i/1Y8gZYiMXHdT
SZb+F6k5RF6W3SNOAns1tl1dt/HwwK8zbYMBjrkQ0KWXS6iqztnITy6J/j76Yx3R
G+4AnOObrqIMfEOvRe8dXlto2ccsaSPM7vJcIkpmViiN3O3fw9kBnUvbkKhuZ74O
daw9xfKkJCcH9S70/S+EOvXzOV8IQmgim8VE0NrsHHLlof56J5PYbU7pksk6fw3e
9Z5hU955F9u7+qEarcjSWywnekuBNxMvxknrPhhCurHFfg+97fZM4ghNUZZfWzdZ
H6cpbn+4rb0Xi7GXaaGsPlYiO1ovZBfdSLlz/OS2bnQk70YjeHH1zrKeB8AObSTw
DJaQulBxPOG6N8fHQbbtthc+axx9QTbhb5wajdTMqTQmV97WfNy94fCYjm0hXvfG
Zjx/6S58eZW3znKvG33kJWd3VjSmoOFfxH8qobhLTc42FwQv2K4RfJQCxnFwK7HE
AZc0VCIckHOvmVkIGRUf+qdE7koDL4HKXP+ty7jjrVDmSzIgyiQUZDn8Dw0Cg5Fq
WqVkNzs18RSjvXaXpnmKG3+42PgW4XnIcmRXxUSRlRHz4xpovWtMX1MkFyuM8e6c
ACJoVNFTBLhnXNDoms6/+ABg9xVlTpSXSupeVj2U0Nx7PVh8RUMV/Ua3GrLVvFgK
HTEI8fBNb7PXIAveGBnaRhqoSI87lFZtmFqgNvt+YN4357z2mXU68tv/bEocfa9h
JUQRyfI/N0wbuRsDxhTJgks/t9nWbXjKE0lxyUjB3hvVzET2LjXC41wJ9YP6G8qs
tPN85TpENNzPoFx5482KkHpZJfvnn4+JDoXspGGqDKWMANrCxrxByNwsOx/s6qr5
TbQFQynZW7JV/Zp5IC0Vj2isXCrjuhvqtWLQLnk7Cy6BJcwkUbHVjRkccp/5fHUk
drWoSjlEiWbhCx1fa5aBYtyuM630QYzlDVSNG5qvf6vVfs8K5PGJIr+yWb673PP6
xNi3RENW/hVyEWXBre1wK6M3HLZWW86FVutzdURHI8yUs1EQ2Yv0ODh1t5i16JMs
ysN7BvgWyIZMBen0h/91rJJK7k7kGJgrHWJwwDCQHjTLM+GALWvfvv/lWRN7GzQi
/iq0ZyPRHQ9aFey1IRWbb4HgFR1rWfCNvrAtiNO+WwmTI6XTZf0NvJCYc6htACmj
0NNu3KsQspntaxP57SOb9sC+ZKGAnbq776VtG5+2NGZv5jSExSaZLDEdVswBjN7+
2AVGjPS7giTnf4Gb0KuAaMFMLVXD74wXEWC7ilHhOIytoBKmIbzvOd409V6uIPNs
Hpf3HOak5pXPdr0nV0XkgI7l9ykxxykx/Gs7aIlnNpUS/XJ4rvYmhxWmstwdJqmw
bkUppSoj6ud/rQBdcw0EcH6OOFycx6Ow5jWTv2J6A2Nk/aVRyW9qWTv8QMPMBALk
Ebmt1H5YCPMbGW9whuN9fOTW4mrA0Tjb282VOifZPCX6ZoUphKd9idUGONr1EAdW
TUdYVV9iDDpc5eBnJPzXt+CtLd5H1yRKzaYgrva8krfbRQvvMS3EjXLxUYs2SOLe
zNz98j9ELEkSgqNJkkCdMq3NAhZy+8V6F1DKHvFOVLZIbY5oeXnp+LpFMMzi/V3V
0MYenndeJ7KxEN6Chc25gL9bexEngnNgx4GXX9o69Xw+ZVfLk0pRZwl3Dk73AxEI
fpvbarJh/c67qZpqMHSXpzoOr874n8CIxez48HB/rB3JMKD4XAGRSOS7AzahZeyi
9da8UKRoW1q5//69/x4tJUf7+t9xFBxpjFLqLgYpv4A76DJsFUsvqDl6CmcxY04k
z7F+15fLrD2mRpjNdNhngf6xbVCnDTMW4f/lrUsVRoy8u8aCSRg95jTStUMTKjwb
/d3Mo/Za50PiuE6Q+2sUs9BH963gbw2i35AaKWsIm1VQ40FyduZEykclUEheoVlW
uM7mVFL3LrXBaSpy5losVc69bweTOKGZuQ7c0yfVU8lE215f8XyETonbEkUyOjxg
ScLRFQkYTaN0MUKlSTyh3wjFJWfg3B2A8XfAFBYQjbw/317qyENHEeYKzpSjg2S6
1PmaDyNXr2wQwSPnxZO7GwwGHfMvGKJGNQ4VFqSHPWn78Z/t0Rg8NXdVg9+qWn9N
gVTPyLdaxDRE3/3o7XEmcFWQiEtNtYMkGPizHPfIxBsohoa33uNJeYyVcIuebffL
gMchtrqb1x5G48B24JLIPPoajsK5wOaunHaqNaFYDKlF8pnUiRbC7X3lFrYTjVQN
/IrXd2AdqoyWTLbNNJJj68+q+SzJQu7nZ8Dmk9wFT1qX0PIeavKEb19ZmvRi6q+P
Ar6mx33H55WOVGd2EM0nvF8lvHFVOqZeyy5Cy0SxPTtICFOdi5EgKNdVZDhaYtVN
n/F5lEjFl3KW6D3V9mqA1VM410FoLHhKJAj39a9Z/y24Ms/5WONIdhm4pLqYc3B/
2Qq2eN/5Ut0IeSi3gy++xVzQ81KObJM/YXBIUX2LbSWnIEtielNkQSjL/EvNVaT6
nbCnX5kCJj3lIs5v+YcWL2D0EmKGCsmG+5DEXieE+pMa1H83wN+WzRF4mPVqb7Bd
Zp7XNgD5WQacd9Xf+hZBCgHr8Wca6o2GlC7jdKndA4nDe/xu1VQ4/syc3G/sO5ZU
jf08goY3rjLFpOIKSCtqpAGDa1hidjGKC/oCS9GPS3P6sYhlOCt4Es60ouroLOFV
YGpsTiFo/aBJyF7Vybp4XgWp6widiiIwYIw/JSMzna3QmfkhT7tt4pxu2HdCiZyr
F58VZ9JtQkRZEkmDgCe1QU2P98gNVJTQ/KSR8u8YSWHkOf3bBj1GjLFRb/3fPW8h
if97oQjVkKI4lEpgD51SXfEluznYBM9Y6c77XqcwGD3rhzGep29K52bzubHdfuYp
BDQx8vqOECqoMP1/BXxI3RXhbZsxnScEMH+OcPJ4GmD+rNEoTtyZP+r4H2dBFwM5
50nERSNTiFdGKgdpjNiu3wn6bziauN+dsWrK8KUOa+znmW8XDOkZ8PQFRhmlKoNf
IeBOehGWQqa2+QDugUsNV7SF/qZAkkfmCOklXXmm3ToY7NuMtGfID0KlDlBrKTXO
94Z5F7hq9keFDHrqb/dFPjWB7EApmjXLSN/vcIj/nmps1WzXH/uXKuC6uDXn8Goj
z1SlskU8AvQ0bolfvN6sGPrcqpbfpjEU3/HATYWCpiATLQ5VAkQACdDrd73xZYoa
UmB2NY1iA/kOKjM6pM/lwTMKpi8v3TTGQV2881aeNhyRp50YSQM0y9F0bPguD7Gp
L0ZCNf1EH7pYwjkqDRVjUIRoc9d8s9ZESSvzKeZwPF4Dg11a5sgOjCHxgedeWLzr
hpuIscncSUn/rb7bIiXC0y/PZgwBpbg17GJm2v1MXyQWzHPrRsJT68j+0omvg+uC
0uEJ0GBTsWjdXr6HXyeRs8sjsVWiR2bpcSzBpShCQKG9/J/W5ZOZqoMWdDlBbWVY
GyWfy2owWu/7NvZJJuM4rhpHpmXiZqEbWM5giJdkfAuc3OID4VRoW+zNFgpMPxiZ
QSJCA3iRH/SWkwtRO20cLUGMeFIgk0n7Hi+lFJfZ2rR7856oV3w9VRJ8jkwBwmfM
GbBAJsFhc3Gk3Rxfwp+/Kee43u13xRg9XaPP9rvC2KahY/rswD84ApOg738iG4Nk
H+R/bet5OEW8Pm7Y7v/hAoslHiV7C094vRVZvm8HCEgWO6p7UTRAJl9cJCnuOCWF
Tn3Q5RbZ5Opjc8OzKqLtt90x7FwsGdPaTIU+XQJINkUnf05io6X5dzptO1ZtnOV3
bMstj+feu5XsAKC/Ta8y8xH9CXMlux+H5RyMcakAzF9fHcgL+iZVG2PcxYWkILy7
jpn68rU720xIUcn14BK4z2qoR9y1XKfbekahk2myPfsaj8z35dHkNF69TzUzHMg3
uT4QqnOO7muMhtVGJWv7VkE6vLbmfefkhC1nl5PQBZ2mTQMrlhmt8ywf7uMq1Csb
aU3Wh3mAJL13at8sGQ3l9kimRreGcs1YFivC0BISDxwG2/0tGop2VrUcN6MSUspr
VUVEyiR9iNo8hOHXb5j/9wraG/7S1h9sy2YqLMu16AbWMgmAzpYgPKX5ErvM9hxr
GXHyOIkFclX+VlIeWYzD/qzg8LSvTWUUunwkOlTpxaPb7wgBFfUf1N6GcW8xP+qL
+Cx5nvRpm0SFDBEtx/PP8ATh8vOBAcVirlweDdlBgVmKJOAWwwNWgu4WWos+e1dN
h+KhxgOg+d3gs20JW+Txa5SeMo35TbHvNJUxjQf9C0d1DNnr1drpPJEhTpwj+xNk
BIdLPvGdrlnLq5XyMiC/9WcmDoewBF5uYHHwFtidu+REjLXfK6XiMZfC5+LrA+nH
OZXu6RcMiEmdUPwWLt5YEffbpst1mrXfUM8fmL/r/hwJoEkWkdcQto0PJQr3Dr/N
fhG/i+vz4bwK/iSnEEoBpKYr2NLoLV8WMd5eFVrFJUYYifcxwWEQlNIa0K11stST
nyaC/Zs/kaAM0Mtj29C3uZ/+aEjJ4ThqKzUuFP4zSLfOIabrs5Ew7X9kPT6RXVqU
M51DLfg+yoGhn8thg3mjEzMmtOD/lvg7TDN8+ygNeqSmEafiWo+XmwxmbhERUy79
ySjlPVfoY0mgBIOfbbO5aDJ5a6KCguvrO1Eoh99WnhMUp5a11fbfxmmEm6C9rM/K
ajYrxf95Pdnxu6+oqtI2xzuO1eEhiw/RbrV5HGZx8fOvQ1KC/WMLCvmKn6BU7DpS
Vhc1uj9ZDMAY+yXSL38AYrtx7o2gsz3v+pMEhyeoplXII7Y8rb5m2c6oAnG5pHxX
leTkW8iRyOqiNJfDECyXhZWCWmzrYVuBlRJwULf+0AQzUgqPC6AQKgPdH1EX4pJI
J+cSszWfBZQ4CCaGNobhjIJEOQihYK14iY73G8ye7egtkV1F0FUUEvI1SWKjl54L
aYJkV/X5U8MPegixiN7pevlPe4J1QGAOQZrKQxldutSCcENHLox2Cm5kBMiIvqXv
ug9weIG6llDJGc6Bg9vmx8jq5Ga4zrEtpCY6rgMzomoo+DOfHZaiVKx2oHf9tr4n
pX90KTikooR1uoduq3QGjVabRgc7XbUc5jQbeY+mzA8r7sIkSCP+iM94DTaN3czK
pJ2/dsJitPp4NBHYJgn1SWNWn1RBQgwjwyCFLtg7w622sNRSgpgGE59jmYBItQ11
2zHMGTyrHeLnD/tuFxZi+7N1h8A2oaBBKjD6M/WLG4f6hkAueOOZHRBjgsgse7rV
Tj6hz0Ic7rGwt8HUyYnK5iXU0ORuK+TzP5HnPnVHt44UB3GvULx+JJoolKAZ1suh
BYFacjXHyVkaVQksKGCiwI2euWSqvMT3cxOGpTk73JUMswFNIYtqut6nJdraxOqu
0D55tNZPsT5VSUl9P13Rd0sXi2h7edxso6NSRJpiC68qETghDN6HQq+P/U5fu8qs
kzr4sry81LpE7j83ZrSJhmAWUhYA35FBxkUEmd7KC4LsOHhfo0L9VBgbGDTUCb6k
MpAUj+KaCOpVWv4Qx4CBniHlK3DDEWuQw1+C2P9hoiLjh6o/o/RiYGys/1Xn8Vn+
RvxysUm03VFI23t/l/Bg0+/wSukdnLzm8wdu8ut/RTRVJYTf2pW5zs5+YX+q67RH
+3E0CcaPz1IeDn+BltXOuINI7hj9dwEFmiKZmZcOrCz2JM1Gr4wtgaGpUyVnROGr
75v9o+mupRZ4zlglmhoRpEuzXWWFyg44HyixJrTDxaXXQNirJIuEn+SGKCmDiHCj
tPLscSpYIH3KhEBfw5gAaBI8FDW77m3FpqOdMVLliZbhJOa2xIQfTxXl6IU83bOv
xPVhhnOquTZ3Ml/Kj7LO7w1BMLWwQr7tJPbs3QGFCD6WH4bVHzlymiBuXtaU8gVy
+iY3GPLaNVVfIkB/VxwW1Y5RYPAs8mDS+mzTaVDlDNrrugYydjQs+LAGzCpWyejk
8Qh5phzUI64A8cPuCkpZXtyiS+bwm1wVH7kSxVfb/vqkb9u3t389uqiQiMwPpMKx
z+GmtJ9TworaXJKuLVNNaQOsi6ycHgRkGLbvWWj3zqc+5yjF6GnD+L1vPa7dTrFg
k6OVVmFy+G2TQuN2t3HWn04oPrN1H4cayi5QcT7Yp2hszr+Xg0VSFXj2h1tDZnKX
uY8GIPrPWARUIy8pApx0wZ3oAom2fY3RIG3hr+UI6xxxgzMpB5F7dI0wHiFuHCRh
RRvbntUXU9JXpLH/rctMskKFFkdx6nBiZhgJS7JgFmph7RngPUGupLzNOmQV8CHp
4On+8F3LfPJJlRHqaocijXNQFEqNRTuF4p2atvY+X80PGKvymXHjidtk2onQo7rU
fGB/RV6rgN0pHbvyTEHyrBE8yMskoc9wvLVufQiNuCtt6zuXNTRUOz0UWzw7bAuB
rdHLSoemFqQ3L7jGGuLCAW4ZatugFSx9qUO5ud3YkrgG/OxNY9ZoXSAPAySRPtzV
v5gaGCYd6exma7dMRsz1P7Ao7LaoXx64o4FYw89XHxJr2ELfCeVDAEkclIoTsH3r
j9byyOWwtA10yw1p2dJ198UfVSb0ZDHiPJNZn7udAKR4DAxpZnH9AszkeXzt01QL
bs/JaR74EA2P/rlZwGOat/ALdiWdfBouOxA0Yc2nEJHw9qP6NYaQdDbYVYAlZ2Qx
TxamBn4h0//mGX/2C47st03m8hIkLmCarXRK3IK1F3bPwkEFSahIUHA5j5wvAEVR
QIlOyDnN5Iz3Kui/TkndIcrI1eg4fUDkhbA2hUhcUJvi+WPuPFiXRStYfTduv4Un
yYpLhLkg2/sfGLuGJjXYqLdWpD/O9rsw8muaiLxo5WooFTm68EEF4dDhcbDF27z6
ky7vZcW9b9K8sWzo+oexK43tT4neDICuClM4CiZts/dm8oVpsYJn/9krjCuvg8R0
W71RCJCPLgtRgeGurOhD12pAkM/zfoJhsbhRFlka7rXeS+sB4eb/6dfpv62H4YqL
MO7XdLPZCrdM1ZfGrxOibCM6iYpPTnRfKBh4GXmXtlEZ0WHMod5Z4FQRne/PZ9tA
g8MPpqBdRNLMJj6Y5V5KVc31EPiFoYTcp+Ke65SmRBIMQX9XyRAFWmiAzPW+eJg3
pevYt7mR0TCeRYk9IxqMDI/oIs6ZcN9vae3eZlJh/ISOZHk90q+CneiMwsvlMbUo
EU5RhOJfnNmIgkC4UCtEgMgdj74ZItu2gBYioCdeY2DUHDe3yaMPH6PoKrJ+3NwT
xZkfEoSwo6izZDZp8ogDnlwALli/qSh49ewWobCI0c8RvAox9Wwos3c5sHXP7Sa2
9wL5786MLuBqPMod2YbP3JCT/iXltnYGSaU0jNogydUzol9yuj9u8flX1xYcXsXf
rdylHhgQKY9rkOgriDqxIQEKpzbDjmk2i1naRJAswBhpqUDY9Vvq/yNhsXA3Fzx1
f7lEZSjJ284W0inWuZHFTn00H/Fxykfuekrw2nJK3vhISwzGebwrXCWQ7Azz/YtK
Nc5Sd6NwcMx5gdR9eH3KrWZ0RfmfftzhyONlaI0Z4FmvjOUUp876KSfQ3PkvKj6T
Tl2gYqi8+3QUpr+IG9jQhoqRh25oy7utM8TKuQmKR834YLD08j51V0i6MMR0pIwK
qDev7O2uk5xwJh8/RXEf7GNKa8CmZUHkslWlx+UfdeVp4Mmlz/x5QcR7UUPX25w2
8XcmQKLLwS/q5wBusehPSx0p8ItFi8izcHD4GLwiTV12ZnckRxBFmYhDhIN4pztG
HpjR7HIAKPjhXb6u6PaaDyroVo2EyvqIv/DvcMT7gGRXYrOuIbgT75SSSKkb3+8U
7JKm+EFhI2swwE1DJDUUPId0lRUncYxugv2TprSB2cPdIyCbIXnNj1123wvFrWv1
KxmpyrjAR7UN5Srts584zNUtWnCA170u5q0qkJBOe7pIz2g7Zmdg8GNXlPdmuk9N
d/MBiVqJ5jcY6VGLxIl0NF5O90mmYqzqGPnvyyz8tAtpgYYFGM9XZoihl+rfyu+h
itdMuam8UjkZzRnEUZ/x0QDUTtvdf7sDw2F/yKiinQ4c3Qw7FK1YJ9V+EjB9RZ6+
86qouPXIOci5h6yZ0tYqLAKV92+ypFaWurpTlTUzcsttbxZvsIgYqRLRhd9pwVzY
3kcjBJeBlp/H1iW13Ey/Zex4B8joyrmxTZqt3tklU6Bjq6mO1g3lr8z6kyOpp/9C
gGHcVypaRh5Zq5VIxRg8/av2uhqPRwk4rHIwgvk4vajSjUTh3iXwRTsI0liPF2fE
RVMJ2+rVsdCMgn14AN3Hw4Z65LHVzYKpSKw/g2Wp2+rO6vvp28jfZmlI3VB1N1Sq
2CzR6tpfwBPW/RCXmTLPqPHhuPLZv3zlamZzpc93FziFPvlyg/h5XrTuzAw67sO9
7LoUAv/feAHsADmue7vdJFle/TP7odB0cPRxuYtnC1vZL6i8iEq1noWpZ1aMfypV
FlTEMSWyBj89xriQdTGrrQzArkwmC0k2o2XlX5EPqkMgqFUyVSf5HrHb7AipjAUq
pKbAou+1ycGawJ9j1vmJqkiewQTatJM/FGe/jqIcjGhyYr+zq7F9R6yi8e/BJ5p3
ca06qR7FCE69eFi9M4GZE5rVQKEHVpG9NY4xrIFcDQDX+zFW8QMTWZx0s23H2ILn
b7o2Ec30TlhgGm5ylLMcwWrECoW6WSTwOkis5WLS77ggLAn9cOome67sK7Kt/hcP
zy7hr2Nw9UZWpMWlg0xXvB/YsPRa18bschwdvb+pU+iGJTsZnNNVYniZa+4clpqg
6y2JhXOVjWUNHJJ/HL9k2tMmxvztdS8+eEiT+2fk2qiP72JQQgLaltBRInn3HaKI
IZKbT8ka36xCTDaIlajQkA79i+CaToIM9Kp9w5WgIqeI14lYuUzQXCTbT8m/XDoZ
AudmzCtzLatwNftLI6NxvWlifGSuLbbby3xnVaEETuxzWmqr1kRxdud2LCbL/QHT
ZU7w0frKTaDIRUUwa5U30Qf5bZKxJMY4gLLJR6Wuh9lA3aWFoCD5dsk3g2hR/HqL
5+vavjDpcbze2AUVfRSKKLo4GrDAar30rwO9iUvt+iCcWb8NULscZKjlJwkoK9VE
i/PfMTS3BlKIe/02nFLD+QXWyTBgFU/NZfJ0nK7hpElWSv+QRfLrm6hhZZjZ52OZ
t3HWnaQXLcQTDKL0jyO4msbg4GqPZG617wYM0aiXUk1bOxUK7Q0eeMBRJlMHwCR9
rxsLJ1339m9DRyg1d3UoDrxgge6j0+IlYxs5u0J9OwS57NW/foonYSxdf+7sDNH/
r53P2gKGCRjA7XSTezHYigKctQINqet7+ee3aFCCdPHDDavK/mDYuS/0dw8ZIhmd
RH6mpOoCeL633KN7+jLhHyFt933Ip6R6AjEmiODyfMjxb3ZB4ynZWOw/6FK73HjT
GJapy5NhIzTgl+0CEi8GFrnG2OfOUNr1dZsB5qxL2p9PkLhEFGvcms8fFE7NiZeK
wFS5vbRIp+N7zihBaRjtNRh8EPxCO3AwGFHg7tDYsVVkiZt6BPRdp9xrLvhHehPl
ihXZIRsUobS2tY4c6CY7S/f13kAtJMWw/eB3BBRwMU/iGexU56zT/u5xmuGSiirt
dIhtLfHcKg7uedidw3GRz08d2syC6O9lbjq21BLwdE/5nmpje543Zt2pylSkn0od
CCLswLJCEmT2pds5kWHAXj963P+hEun+5A8xeelWA8n5N5Yh+dC26tHKXlKaRwhn
ZB7itbk5y/pKAwJ19HLHD1Tl2EZbtvh5U8zhlw3M9cb9EzOdFWSMGoh58Mv8mRNz
6VzoM96ElotuXTLBvxuADwQZalos6OLqn09bLE1LSpUyeh9FHpaelvuWhK4uzgjn
+xmRdazD88IE6hwBQUkcygwYcivCCn5dzOff+9x0+n8LZR3vGKUiHKOFFN0gLzyq
3YffPMzk94nVb5cCxKFKtUUiKFKSMm7eKd6PDLntAv74pSCAlcpHV2SpKhyLGf43
diibY3cBau4z15qRB0tKXq7SxZ+FynG0oc3W1o8o8h8JfaN0yX5i65uTWPjsVdE5
grrBshhZoaGwOnc4n+tU7tWk+xjTe4tKtAI6JGKUPS52zDCB86Sjn4Yjf21QP6nQ
RfuJ65jurHRRANaeyJ+H+0CC3G4unLX7KhZp04byXVahbk7Wbqe0jjTBUZiPrIM+
vlCTu2+YZozB011ycfq9oNnIiU8yaMyfZ8UG5bKbTDgSYqJZqvPTgFR72WINoxte
PL52xeSCuYyO+5mWLzhSYfwMmR3jT5iUJU8GJAv6tBLAbhq6yDoggS0H6RDAwPE8
H40hgxbA9ZICJX7fefJoNhXvmNArrEdQSTseY2iOuEz7nqE9wA9NyvZMKhTDbYdr
1yXmAliB2eXKU+F8uXNneiEzpxia5G3yObiCO10+ci90aU8R+oMrdWvcSfnO558l
Jzs9LkSdqRjwRwBgaR2FyCl6FvzRC4q6u5NIQ1ac0812OOr8nT31onRqSN+mxYT/
+x4/s77kwV8lCG/ESahWUDe6bdffhjpB1bkLtSgDwV0CHPrKepD0u/lJbAmg4eyW
Vg+oEZWPeQErAJ7dsaStPIKr+Gv8Ti8RCGBH8HHwgkH2thtfXNx0/Velqem9YdTM
JY8LYQQsfAl1MUlGKkOUlNAiL8mCtz4rp7SdK/ubLXA/KBszmTlWbLqhpg7lYvxr
/TeHCJxD2woONi4Z+SopKHxd8yPicukS6hI0c8dO8pnoWp99be8CX7rdiLgj9t7C
Xy+immZEwlb6C0ih0Rw7I8UaOmTaFrucjDAZ6HwjgpVlaVCzxjHD4yaxzFBCoCgy
1M6DeVCLINlJo41IGKnyi8WcuWSLtJeldN4PRecx20sG/bwrpZHP4bj5msLSC5Sl
EWb379fLYVdEDUtyKf5edGu4KeutMwNVXKC5Iz9KxHjKsE8BtI2WENmVKNlZAUkS
vyzq9WHKYZ9DJ2Dh75QHl2vLkLBfsKMEv0wcQ+GzgKAtuC6QETyTaoTEy/fIqOuE
xZZPazdIfVrDG1scKO7L0r0AqisnkSc/88m9hp2Rj8JMj1qBlneqS3zxWivp4ciZ
yytjOlwM7KgEH85zZqLcDGvlx6c0739VZnDrNGIE+oFwDPHRf0KX87Vtd/3B4EUa
YurYG8DlOhzkpzhVZiO226VKFnrL0KTXAi1jcqOpNXEiYJArCAmhNKtPx06QTkMN
IVTFPC6KN4SPV+Ez7jFB7fK0W8bFQOsUxgggTh3KDP7zfOlT2/4GwilMdzDBZT8f
3sWDfdflyzmGmbnaYXKfElQxDmM94ATkZmvSxj3wva5SOWKPsS9iupZrxRJwhndD
NosQyPNEVPjmTzpnQlRTxj+adQxrsnFyYgF3BDvwnGvnMZUsBssUOFErp2qKX71R
G1n7yD8DGHeg86Ph6UwREQQR86AeaLCCHMyw3TGHHjBBxDfzjhLuJMHwB/TdHM5r
CEvO3q1rmX6P8VjeF89JoOtcpBbSkNND+WXlF26xDQ4N9e41PJpFLh2UcRmxaPj6
n5SwJ5P3EG946zQuOVqVAE3blIAX5/fvbKUMF/c5yrBnAEnCr3o1ZqwKwN3DBVgz
7SnLrnfgoZqp2b+DU96fHdKC2Ogh1wIiRWUobY1TSvbzWgN8As5o9wfjMV7w38Fe
yd3J+inz52L0jcbvtwxEmfsLP85PBix9rUL4n5F/J4vq800ZU/+HfdIgFFKCTZ9j
HyjjdNIGaOd45YtPqaLjSxuRe1rsgH2BxL0Z6p666BfEvH2zDXrFvW1dRSiPfTz+
2LmtBMzh0PV4RFb31m8ahe5d8MTyd2khSVUYzZLHS1+JlmXkXoOEEWesk2TLo8HM
fiVeZzo7G7o6I+9Z5NGTrnhH4tIn0QvYSBQyRoQW3aBGdDFou7j1D3d8a8YnoKvN
a2HrCvh/rpmWgHUdDTSl4zFwVJuQh7ZdHVkpK4RaHr7x03/w4ZCTb5zETBnPISIf
iK0LrUoeebNKMLWVE/Gt7kMEtmzAP7JozuWKMNgeWtCg9GD/y+ocGOaWX8GLTXIb
vGBljzIU6zCGhRqHb/GlqgFAjgtCsFG1j12jUxVFsUhOmPOlwroqB1NWwpXjG4Gt
22SXjbBcoY9gjLU0rorTTi10/c0106X33XukLK4n8VoYcsmzQ2RT1+HBV+fL4WPT
40AThd9gWDP30we/Jtl/a6rc31Mf09GP5WW1Kk3beDJvznV70eD0dyn8Q+ptLri7
MvVNAr3URvyKqdv9XrdpCx1OJYmlyzKNg5lzmxAWxkin9aQxzThXyrVdNUeBpeny
Nz2eZiyf1V5GaeIM7PHPTfVr21wqWw+2ZKR6o5esJj5ppWXdnBTssEfaZojB4cWN
bGORYDMbbFeCoz3MqVwNkTfXRZOn5IMxUvNxOySIuzIxQNnto1OrWelJsE+aD2cR
haHfnFM5m3tfO2xVoSSCblsRFwZil2rt2C836dg+frSe3MvaSbPArnuLiwAZ1QrQ
5xEZXMywdeOgODSvUacZUnfXCTWUOLuXTQLsXkATtTD3W+z7zqNekrEO9a6w+OGd
6UXD41mSPnQOP6vBOb8QyYT6vLd8abOK7mmsEMlxwV0ptfnuC6tNW2IdTGVgYbV8
15lhN81ToYSgigIjCSoUOln1LS+Sk5GrIffi+Xtqk1uRVawKYWlgCNVeK8ikiXWc
WMaHFK0j3jeJBn52/2eqZsHR4PrgZKR8ur1narYJW8ixCl5IzgUT7CJoZhcWa3wb
c38VMOJXwXvq0t1VwmrEn5Dp4I1jyP1jjDE+ELN7Tt0xekUSn8JiuAtHlUWkK1HV
yx0d6ZWi5pUARw3GCIkQCFf8jLejDgPLyVxQH11ODV5b1lfuzLAkMUC2SzWYOe6N
hU08ihqOaqWyMRNs9rm7rjYBWfSzWGbggHgjija6BTk8XjlazNzntg6JXS3S/RvZ
FxIdqzWOirUb7QQwqYha1hiZueiZGwxLOT0aJ9U8HzO/gDEbCxOaU6n8gzSTTagi
ESaVttIjLCKwNDBXHoEtKnVyeD8aLd+dnyFc2YvjIN/9nEsUvgmDb7pDHCA4yS2i
6HR28pEwjva2fuWcp5INIzuLRueo5EUHCJMp7/kykJuiDL4xyDVHDMbcnmXFb5ad
KXJN/zz6o/mJt88aXFOLte6YqDbjT+xyornHCGOmFVfeP339ZY42kb48KIUhwUIW
ONq6AiHT032C4F9Vfurpi6OUDyG3RGUuSTN5qmFMc0WAuM6nIYsG4ixRXd0mhuUz
Bkp1DLCrYfWUTWwNiS/rxndB3YDkOYC6mvd4/GX/PA1d5tM809xcZRO4N+C7qTDF
uToYF2g98knGF92gewi12aAiW/H8OGWwQiDsyrx3KZTbGN3b3wYkbo67saRT5q1T
z2Z1ty3tSa3eCFvOtnwODtF8vHKAzA04DNRgT88+h5+yCEIHSD7nbOYNWwq1O+OY
h1Hn0GcCLxt9dPL8XUfe2v5fMHq2BTbtQTWYQm2qnkOHkwTGi1+2SpiucaZbkWMT
hukk0AwzuYKB3t2yK5YO9cuAn/kA+KQTUxaB0GPpKVUDTmMiKTrMbB++UoreeqrY
rX3XL/IfitBVSPhEGxe0LsdHZ15xNbB7B9/miF5s6RBEEblbAu/BPP2OCk3NdhL2
g9mw/GUPMzvW7HdmWYW/fvY/+e1nkmuC2CEfL7lNOi6tXslPbsvPt5iyiQZFiPji
Y50NsEr915/FfVYW0X6CcljT51ybKyXnKGO799Mp2xIsNPJfWTI3qPE9lngAVgF7
ySUg0T9ZSnjITHvuZux7wsQRcSIaf9aupjr+gz8y5A9XsX/XDJ5CuV9w5/yuSliT
CeOIAhRYslFuoC/mQYgla+IA7aMSfnpAXVNiE+lO7+Nt1xwHDBftXnCvVSsBPxlw
PpWUu83TyJxD4L80vywmpeD9+QK1FOK+cD3doYXViV7MHZCn+PafkgPAE9ZY/b4Z
2qnwIhwXZJMTpfm8xPiVt/PyBrgnQ+P9Xb2mw6wD7PDJcJPS8TDD+qyvQc4NQRbb
CQ3nBJdAimdwM+BB9c9XtjpRDVauDGrW0RrasKU4fERfnh2cKGadtsnaeopu0Nhj
NU9KWILP8cLtpN1E2Ep4zJ2eGcaG8oZAUIeQI6NVviTmxImtTL7RARpKoCI5wvlE
ll+RokKKSXhTxADNLk80ZJqUxw4oo93+1C7g2MNFZNylKuY4DN75VviiQFYBHB8y
NcojdnuawwkCfr0eTbYCdHF5clwZqGbr3QyST5U93yTVnvmT6idm7wIUeGDEHTBt
WJRZQg+1QEEem/K8nEnhua0rX4slXLX+OkfkRgEwQ6K/zhralk5iJqHHv0fk2Aq/
HjaA+ZPXMZr7bNJpTaigVoy6MeWDV3ckve+oXQYWC4A5DLIPFGlz4WyTu+65Qbo2
iTqGA1XdXEu247Y+MiI2Xfye75CoCHX09JsUrtOzd3JGRfaLpzB/X1RcxfKKnOq7
nBaHZwtbQ74p4UkZZ+5OTOBFRG1vnHv4Bm33NkSdTY7XH/rJWVdy0SPJcUZ2bk6v
aO4NuQ4EGI+SMaRYZKWB8NQ9RaQZFtfT4NxCsnuZj7WqSN0egOX2YZvI+Mx+/3+x
pWQXbPF2Io/KtRFEQnmxWjX6lm+lozlEtMy4CVLfSim4b3yHpYO/FdKk91R8q3zL
od9dOdy2KPIeTokQwXpDmMrIJuSCD8VlLOiLwUyUNFCOAwLgI5aRA68QrUgjpyB4
8pi/GIFa6R9UutXkUNt+Ow7Bxo9OmcgEJ2lqZoWJRSOXnhiwp1+3kyCrqs5FrokE
SbLsNfdNe4dB47k3vqRA9MYabulejIQhTDAi5pAGPBymzAGHB8Ffd+J+AUk0xYYb
IjW3fJ1vgTOs5jNeKr2DiT2FYCdQoV471JtmLVLLRNmJUuGNNPGAf35JkBLFOnWR
DVzfv3JripoJvwb7wTlODH6yJnMPXwcQ7BGnodyHnDxmXWpYXRVErxzZDWfgIOtA
fKl1LUCb3WZ4lG0O3oCA097oJpJOmNVQPKhGBCIX/zGtCi9HoAAxf1kSS4vqr6ot
tmrj+/7Q6K2HZlB+0IJ97MsSNJBo1gd9nOYnvR8JU6gMaINVN2r/g1TiYl7HQASN
4+N8VuVE+RRSTpAO2Adxs8sbzvAvtWka3seinwzBLeqpeyPxFJZAUay8AtlHZkdY
gPYmYGTk8bmFRtTJ36wcle0T3AjfTgp2NnmgfZKlpb/9p9p+3EJpFXlAKVqkixWj
BIiKpHakIvc6qg8Hdmfzilixre6AAfWpvScTx2WpciK/17KQb4pjo4V7P9HHKd+p
BEFaf2GsFXI9IjghGea4s8xisE+6ZhT86JMuWXVmUpsygjI5884pXkRU8gtweSUb
n9EKTAVgVWoi5dSyq0Va/QqHgUbaqt+5UXakkmhqthlhix7DZ8PZyjTqFnXRjGYL
ID4njNQeXr0MP4EgvdoJZKOudOMMZczr2EVCcN1HAI4xrvCViJUvxirvifKqWZtb
f2XR0V567GKuefsvrUmJ+Vb1HnlZf8FjWsadbIjVPwUusglg1PxFYKM3feZLduYh
IcD+wbq8Kc215ezqmwzxvFCnTUk2gMlMRbkdNaAnRp2rMEvafeUmNIxz3yVNNmo+
4NlBdM0/vj/IuniZUp4Tafz7uXDkkmOoX7lrmnePeLkPfWmJG7gnBWG8s7+Lce8j
FtDmvV2kNo4yYBcDORUuTPRRIC9x6DFSxGtdkUOfQzes+6DO3SH8sJkHVEy1mG7H
DFztMDijGdyXOdpG1TAaJatvB3TsaXzjIdlL2YnP1aY0j9CqX2D1t/DRoD6rrxYl
RvWp75cK3Xfat6QW7yWy2hOV10DmhDbHds/PFOZuF3jhJdrgfDCek+kz+BTCrIFM
DVPVxZ4nPe0+XhjbRKq2r0leO/BtnK8eW7TTos5NjzYdqXM2Tv754WjdnooEbnUr
K+tAeZIU682GZecvKZYyA9HgjtOpRYY2gKg+Zu/8VoGRzZkKB8cKz8uo2oWuEvVg
2udhV9GIejG51UdfPJozzJl6vA4crlY6+CECAfhZ3YILDr2aHretp5KAl0zh6wIc
/ET0CYkHEgeV3n4lQkLLvTS6i/6lbB8GuOOQtzhSqoxSxjR4osCj/hcsCQFTZbXc
yD5Tjg1zVl3CLj8ZOgJ0QXljLeH5Nv2lB19W9sNT7FYAf3fw6MUzct/NKeEQGw7T
dAEPoIo53b7RPWrsebL7V7n37cTU7QeH54m9gU0+P5y8Sfrro8MqVHh4G1lP6knS
s+r4vBorB9RpMeNaUj6SW89wllaa22kytSkNK6t4TaEVBoUOfd+qIVbWLEH42fyC
QtxvHHOySVNp1/wY5S8dqTjQbx3yh60PqTAa6V+S6jbop+xuxjtXxO638VPP2g+E
YPZM+BKM/1nWiwvCZwZUiRbRk4TWW9vN9zv0GkeycI8+He9Ho0u++boZ6y7waOm+
SaZ2qvtfz9iHj//2JFKLPC8QKFsDDYbxKjBGESPQF505nI2bo46MhHzIdc5kjPDe
d+DuNp9rxiqmCcGYT8x1xKZBa3lQqQPhXzBaEOerAF5CknwmC5JfN1Yh7sAdSxDJ
SLROeI8EPHSkc/bFCbWX2LhVp/UuQxey93lx7b9f8c+beRTrOTc/xhzlDBcelQoe
E9gFB2yH1dy9EVhQmbKKeFW2ajf7INDUbLghjMQP1tmeulSCYd1Lmlum+R+3B+l2
yBEyqrvsdmGzdsQ1ZIKncUArhmkhe8q3RYjN5QU9JKZupp2ZJ2y59Ah3DbZm860V
v+h2JuXLqRJpFZSfHx2lWfgBGOemoCHqFZw0tuSZjtHnoqLH3GwdAoZKPPhSLvFN
b9DFZaMFBe/EUl+ZxJ89k5BlPihT/u4eHWhM8jntLuWuhL+Wb8L5khoTIiK2DEqn
f0t5m7yQmHai/g3I4n7ZWI6ki7vZsbZqabh8qtNuAjK4+Ya0H8rLzxEtf3Rr7zg6
v+Yf9mYFV1igjgvyL7s417BcOx9Lf5eYPvtla3Sgtx8COQ0Q0pAXDu6JHcsDsLWz
+5BJGw7tmtWPaVK3JVXYJL1dhYLYp/LuvltYhDdY3bAfM7294vKrFuf2D9jDn59I
4SqHkFKqg8XGSu2rEX3F3WyouBly4IrJUAvyejEsD2otb0O7Ic1IWVJYR3W9KY7N
cGVLYpDcKhgjauP9SdACP7dyEzJZ0lKPo48doas9tokfmfU9aSTAvkpwar08hR77
ab1vJCnzhWOgZJAEakC2v8JRCy590c/1oUbretfJDG13jEa+0gBPTd8LUC2U8q/V
tFFLcU/V+mrVfg2i/HKtzvrdGC+c9TpLQ0CxmxkaEufW4Yv8Hjz1d2MRA5YlO85C
Ok/s68MY1vFVq8NHFBrZg5QAdxIcke2BPpTBa3cHEgfyCY5deb91S7Mgiruu8ON6
Bsy0/6Bm8Ie7f/3kIKe/49UBxG2XPaK8SrBEuAL6pCJNbw3+7yGhYPZz4tZqp9bl
J/EJjiiEYd7po3BG8U5E2ynX4cueKjq3wag8Uq50UqouBOJJXV5CTIqkRJM7In4V
hlmJQlrBTnhatt3UIoo132JsXr+bHVaLZxyKAkjBjEeH6/O2IP07GgtyMpMthwBH
/WCeDd/bA0rarGKhgA0i8F+MUwWSW6ZMzcDosc6EnXiRmmaEMW5uH+Db3zVfu0uH
6lWFCGRI/y4YCQWCmJqccQksCk//ozY8uuYwFBN/pMYQJ/lC/AnYI4/llbCos9th
OyOx+7HhChyZETsQTq7l8IS+u7bK9fMFHaYbuuG3OP8C/B0HSWcf/xZRvpgz2x+E
Hf6Apihju3AF5ZT5Q1Q7EWdpIgiOaLRScHDKinmn8xI4J94FhDfToo+DwdlKI41h
GFNBzMyP4WuLV8ol3/Iq0WtCMxMS7zgxEOOQuf+cdK/t/gvgrm/fNSZuwx+HB9qW
mwzjvQS9gUS/Eu+9bmv/79+A0yPkJVXAavjRFKfj+2oJkTg/ReQYYTdJukv77uKW
tl0NtgU5as3hnhQcN6KkrbVq6Ovl4XY+TsnYqsyoI5JKgjT1cl2DX2ayNiPxSvUx
hMH1S2APfquL5nsQGRoFyahuTtEQKuvIAcK1iHK8TtlZRwui3g2gVc+fZ7IEp8Hy
YUNXY5ZnO3v5qNfp0/q4nFzIBswV9qHnP1CZDAFG7MQ+i6hwswwgMimbCFDMVjvo
xVW9NX6La3wc7uaApCqAS6qjzrvD/Sv3A2TGyJAw5MUOG1mtFnRq2laoxZD2Iv0p
m0hMjrgPgOS+gzv9wITTEXHAN+27c8hYH6J4HIJA5eVYdSlyISTY8RiJT4Cq5MiC
Er7BIW/kovxwM4WK+9OY2KtMwj7D3oGIs75K4idFi6Sw6MCdnJ6CQxSHj67XhhXx
Xki6mbcX72aqpU6o2VXP83jhj4lXWzuQFVspZzTf6ZW3mf87UgogtWxTtR1tgdeM
xapU3XqYG2WmC/D6okc2P9q59UgUUki8SOujkz13Ydi6oXLwYfu9lDOjAa5qxFMq
roVlwIRSzQWOHWwBAvwj1X9WatAPw/MKQwqqe+R3oAMSHdB9jrMELc9IJMnb3zU1
RSOoSuCIbvjcK8XPs4WKy3FU23Ceet9Rq2CDeRIXikhf/icRD+FpOdwS4DxsQSit
09ob4O6uSVZEcPNJUKyWRSi/hsyKaKsDk5onUvWXjJ6SqxRKCTx5ukGhVlsQafbV
M4b8azo1oI8O+jOsYI6GNQS5JJR+VajE7aWVgVzoNwRp5fRhHnxhcpo17v4TbgT6
BbyOlTXTKPKs0ZGpQVHQvEkCPBk+MXvkS2oa/Q/yCtBaGNoJf/G0JeBNUDk32BQ2
k6kUrgY3j2edRO6u0ABk/qvy9kQzYpisXRNo3wApNvXhtSWpfwUqQIqRuZzfpneg
m655N4m64zKV1bwa/yP6WJ2ELYBCuIbwYXL94rotmbO2b61amoH/JJR7sAjxMtXd
jOKG0gnAYypw7xwCDw22gfVAotS0svMkp+uNJVqkVxRS+sqazD9oT2XWQuEQ9aP3
NsKXTy25/b8pYijfcNnKbTKvMeSsxMIt9hnE8+OSMNRESJcWMJONVY0wYuEabKgp
rp3ZSjtnwg2I3mRB3lY/bmjSYXN1XdZMQApKcLzo7PWfkF/kKkjOg/9D0QsbDwqR
gz3hEMYJZY7SIcW30T1cBlbkY9uzhG91ePgNsC7aiBlW6QzngG6XZ3pnTSZ+wb+D
VuDOuBQEZEUEg55muxPGVKoebWhyXRfoqJc9mOWjalqOUprL1js5vLvEmqVUTlcT
n/r1gSnagAFClnlzZdU/MCnu5lBx1e0CLAT7f/PV/f7YOV2FMVPDv3sJWbtJ3ohF
8cp9wx/n7YeOJnuYTz94SoZtBgUdPTMumx6rkP0SpkcfzzxFOQuXpIklFq0rq8y1
RPo9I9Slzr0JSt4N3HShEn2WMdZGdYbXRVAxYGG9+M1lVyyqqImwiBUd/v0Y6Bys
xqLZmqMxcwZsOtyOkR3j7oCB9FvMKO9u2/6PvRabAAhaNJDvFxWpZyFY3O1VLqkZ
E+Jg4j0f1BwcfgVnudPR9VSRzRSbGx1EPOJ+jBVOAPnHoqr6gFE0enHYE+AAWaQo
gVXc6DHYtQwD7kWeDeq7jSV32x9TCvOhzonTUgRNlXRQFIGluEetM9+Fw2VG23vV
NZIpae0RrcftPSiMUvxuVmkttsN1L8FylTCxXwhZgUJJfF4e/cO0kUNaR8mIQHZQ
m8rczRakEYa4HWYl6Hitd0lHdV2Iozye9SL/1P2CWQx3Tbn/tx02yDEIHumllPIE
rjBW4k6Sd+cH+iP+5bstsP5xaqFUhEzjSiT5k8Q+LM7CVW3/EC0vkAJDtuHRMiDS
lbAoKo11h8nB549uK/L/+3mocVcaBxO/lt4QSFKC2i7c3pi9B748y42OUrX7LIbB
N03hbzAcKq4Zb13eHJBtpzdH8gI0TycPoy+x9HJDGX5V0PK6K/t/HOeFM7xFdKSz
iwHyZs4Mhu6JPB2wUvITsFRNQyS2Ij3GknyEE+HDKv08piuRr90ObV1fPGE036Qu
1IkoxK6VX8deOnRuZL65DNX6UC+8oxKNgAerABkPHqZoFmVhfoMCqiqijQXmsZCl
3rPw15O1FHurJWUfGciV4SUuyD8mJJrxgGb74wO+IgLWI7UUR9CeH2beiCAeG2PJ
X1VuGFrOwhVSt1/6Kq1/qKJSSiGzDIaefu6u2BxE0SavXuR1pbAHqaGFwgggXH1m
8DFSwmxtqUQyLd6h7lSdw5kczEL9mLYjTQoNgHOKIcHRtPkADzJqRJcFoEz6k2WC
aKPm0FxNl2XeTFiQHSSr9arbVXe/rk42nzn2+hBFQikrScWv0pz0eKl+3JbPwgZZ
/RphvNh426/WyvRV2upXoRhj7062YXZGwhhMwHZP6+aaE03DBhECfjYfChWQNjG7
axfDzefjwDmMtSaXerQkSHVe5L4SU+3uO9OiiBGLVJGp6rRfdrZALv9y3Ssq+4k7
ewar5tbrmBcQn0evmaEejK2Fyo0xcTaNag297GumkkXIFmQDBdUV0LaIi4Cy2tXQ
fFpS+Ve5faL3OXHBQZVH5jNMP4OEx1mwbJhQMah/e5bwsy6lSQQ8G8rvdcPLF5ay
08rsPD0CVXUwCtcFekltvYRcJB6ytL6kc7GzM7wZAWtCHNOZ9XYsPBBQ/dPWLPR3
Te1WrA7s5zUX6q9/I92VFHzJLwqmamuF3WIUqoOHoXagu53i4Lc7j2j7z/nzmmET
XYLLURRG2ZBJzRp6Hp2mnojDa0A4t1EMgzDKwMgu1Y3uEZBAewZQw/W7IdjvH9om
XCac4zvkL8ksiqZh9gcz6gg1slnYai4/TY4PvRKGrAEHjtoOf5EOK1V1RaNMrXfm
Li8iZkTAsMBCzAEh0d5JdyK9Bg1nAcpOn3zWokm+wxjxV+Hci3/FhTJR6eLciDcj
l24oL2Oy52Fz5hc7LJX/58wGr7OVJWQFykjI9VSffvuf4kycQi+KPKfTRqrVIt7V
3dXMe32SP7XiFzgWE4rXQmrd1Zbf9VCYb5yRqrsYrRPZkmXadKSVpEpkv5kG5b/z
jMazOwY6MP/tl+zJaEflt3GP3IjnJrAGHZdj7XmbCXoQ74aWw3uFI6bgww1O72vs
ZacbM92dqGy9gRtRx9d/avOfI+lwFejzBfOhT7b0Wxf03B+sJLKUjjtBT0IFYRoj
TiMMDSv8YHHeZ0Kr0Ushld5T4lkGB9FH6wsVhP+W4P36TFjkAkVb2aKMI4aNxG9x
5rxtsE7pwu5GQfO9APBZ3Oy1mqxy9wYKP2MwkXy1fSyJyuAuiSKaCnNbfDJgdaz1
0rReE+nMBxlpCFOHajOeFuafY+QydvN0ytmrddaavr6HuJ7vLgmboJw+dlsQSnpZ
3q0PVZ4pIPD/INCNGbABzyEpscgCr9q98/RBrGqdEtCEa/3llpknd8qaVJJp1vMF
IzFH9kFjMm0/ZhtpzhR7W85UlkOnUZxR0aPvqWqIoRlf7FLC2Vm0KupiEYzUfr+F
kzTBFYMbU5zdQv2d9jIOSTgR+DlQS0+wwTG+qbp2EtWGT0UN6slJKQvILpGYsULL
fI1miWvt0qNqV6RzH5o433WCATcSafkcDOggWohLOOCfXVdbyYzAIy7Gd+ZvdewY
kIgZ+aa6ie/3NNnrI6oIfDcO6Uiizc3YOObTRucbolQFdMZ7XqanEPNx982fnHZq
XiKP5YDj08RFHDKE9DYO4my9xXpq+qtY1cpcWmStUpoa7RXhPxZZrespxJmue3aK
87fexfjXIv+rWXrjZElpXdzJehSWwegqMSEOjHc1j5sNWdqyrMd34hAeBUozXLyQ
X6OlwmNuNNW1SU9nd5h8WrqQUL2e0aRT2vHxUBo+o4MhVSnnFkWB5tkwAzLlDZUp
H7f1d9NjrfaTq26kb+AyZoTljfbmBtF7QXHR8ikLyNIVS4Kdpit49JIkc45X6VGc
0sWzvOJ7GixjdicpG6gisQqp43HdY41Fubn7FVc/ge68r4l9FEnYkOg1U9sMsMht
xB0rizO2IQmCUNbdSBxqfFlpTBFUBz3dZEcncd+xbFb+C+nOlGKuimTHV86I06OZ
GFlNBdrTp+a6YQDDwIvBpUv6oY9TRTCPMg02LIdvihtv7hj2KZAh2+mYW8UusFSN
QKw4lP2LYUj6yJQC2fT8KPyDMkwdszBi27kEJIyoPOJArsy4RPBpwqMTwQPXzOIY
sdIIjLBOr4bSq82JZNtECBrKwT/iZnsTZjaYKuEHPBJsAa228+26CTsYy7JW/LaO
NXXQZzF+/soTb/TWv0rCJXoo6wBUJyCdkDCkqnWfVOqIPajyCN6i8tNa6TRxWSht
piXIte9X8nvtsiS2KL1EN0K75vQoveWgXiqRiv8inp7MV6ECcjvS7PzGUGSEHa1f
sY+7FUpM5dSEloUYRrvnZmz0plF0EiFlxtdoA9sVjaJAJicvsa40ixmPKbR3CkaG
IV/yoDMyzITXrR6Au6tCmEq9aE9ins+4A6YVc3m5nAw/rFHDCnYWcSRHxvqguvRb
BQ5z8R4b/t+WENNZddKk6Y7BKG9oeCthqVA5RrQ5vxYU8ylGobyMyi0DdDb9NCCs
Mz0zxsd7T5G2wyttfOfLkdb5DxUYFr84XHisQ9VgjYdCBS7Se1h0b4GAV5vn6xOh
aYDaAJdNkskeVVc20TvTcDu7cGg9mz7eijOzeGJ7gyOxn3HekBTsqPYni3QyAU3j
YNGPeWuOWVoVotgCZciygGknrtUOkzxFVYszDJ05wd62KtiylECr/JcuqQh2q89t
Xf444WZA4GFKABWPWFXnpwjKTvOSyCdqaJSwk24alR2ecBAVfLWxQTVE/5DYTMC3
Cg903RIf+kjq+yQyfSgEpQhW9BEPxqLFyPDh9ZdAPSqabmE07KuKZJEEv90MmtOc
+oKeD+vd/KDjze0CnSSnuMxGCVqOIFEm5pcOjWUaLwOcLsdJ9Fz2c4FCnKxMw66S
rQjxCc9Uox4ihv3mNRh7UmLQL7Z7f8LtoU22RanyTUULCeQAqW+pPpoPnwtDUvy/
2OS9ni41m3TLieIB4XI6g5kmBfiZFu8LB0MTDKG+MEJaBOLbSA5ZXkIX8wVCSs2f
dFAOqBgOgcZ8OvLG9rjC284UbYGxn0NEAPoaAgs+DrdPQE4pXrhRYYwhoHOAxyw2
8GeqTgCucNwZqZBpPZaijzm86BVesgjI09/gdNviubT8GUrhKoLSPT9gVitzjGbX
ATLoQ97+9ekMB2Cr3+lcECgXarXO74OBaLNVdR3CUvjRXAcVycXXObno1awDnroQ
j8gISJUwI2zsha/ZyswWfkRmOXRHeaxzUFhLaLuzY5A/t4XTcMcudvjOXmD0CCW1
qQDiGFfoVrZiZanr3nx2NuMsDNMiDIi3bylx5uyiDFNgrPD3QuGF1afuuY9KP3nN
ls+0Q83FyIPtg3kLHJxoERdAr8lXEBcV8aY1y8Ne9yQ9XDyYTwBcXZ0Q6DEpk3xV
qUL6qRzeK4ACFHdNVxx+NvI/KTC4k9D6WHStlnoa0unuSSDqO9m1zkwKqi8fr34l
Zr2iIFnSXNaNy2g/I306gjVg4aBE4gcp1IBDkYJqaIls9EDTCc10lVdL3wUoYnjQ
VB1hIGd0JHSjGEC/H5cNflcc8UC5jdojIhtq32AqW54ZRzwhFpPNGzqabYY0KIv/
APFwA62gX8ChcR3O0wtLZS3udgyScPBs/hHKRfVQmfdtG1sphxwoTHLuVmzaokYR
jaK1at5L9b7tjIfjXDm009Cu22kACda+miy3HJOApCGoCTA9ZnUj5kHnkDR+8vHJ
QHIWpUTEHTqc+0zjl3h1RG4cd6wITy39eJwG9cSafIt0uDwtCyE4l0XToTrOI2Gc
JT9lxTAfbulslD7ku9oEQkXvseGqc+eeztpwXZnmLJRMJzv+1F4mYs7hXqZiBQxY
1HdxLrTC8DgvAJq08cpn4xVU8dJ6km+UpKcjOA+zUfRO6hbZWkE6qoNA3ggDymlZ
Y+L8rgczLqlxbJwbglvszzgnRGnsfB2br7gmTS7o7fMicBLKqWG1GhUALQ4hbXuo
iI35xIHMQFYNjPdBo6cMtvLPYVvr3L8Uy1uqlPOJrnFxC112VW5GlURQrxemsKZz
kX7Lu1hcVfAB86llx389VC8TvoO74vxMOPv9sLTFomdcBiimwFrit8v3RbQrfgH0
M8cWqem5duBrFTzvod60C5JoMh1RIPfLraf1be9iHd9Iq8wlUvtK1XWx192ZQ5Jj
JLmn+6zno8r/ySpVrcfYeplrJQ0Ky43+JKCgiXP315F5xDqzmjvGY/AyuAGQMK/P
Y5tfIvxmQ9dZ9n4U2e/Av86TgFdiUnhUfCHH+a0URgACzSbSmPX/OMh4fJSttFL6
/tklpTZpeWZf7pumV4cRRVSHwPRmQBG2w+l9Qt5lmrQkvwkXNoexZsaUQYrrpV9Q
RrY90DL6TFsnjfTmaZGEo2km2ul9+GMCWLkML6PIfrS6RSyeRGuNrohwqLZ9rbOz
Kb3EsBcQ3tjyCHPwveSkY+X19mk8GnthODcbwVUlOcwhNoyI7RWmojqcFy7RzN2F
KxofJg3E+IGkGTR3Rjjl5qfinA/LrFjVZR0DQo+LiVxPcCzgWrAEufya5m8GCfU5
YPZYfITUYSOv1/6Zy6hOp9Uarix1U37WhSePofGY+cWQsitnEDQJIPJ0YgqYKo/P
Rr1SI7iLOcXKpjwpWmgAG0UgOQ7ZOqZaNWaW3s6Xmt7d3G52uUwNJ9GMnD+ZYdDO
UQdB0UbK5YYrfCpB9YaFrvPZoh2ehRapyCJ7PMT1UgGA3qYDbj1x8N/JkzR/DCG+
l1eTXwEjgA9FWHr5sTyaVi7K4J2CJIEXnBjw8jVjEx0ycylHG00N6pAmVU41Hbes
OBdcKpZ3D9WfbB+T2mNZMTNk6m8nKrFlps4PEbsIu76G55vIv+L/7elfFOuftA62
AQw8bu1x6Zf5S+rg8CjCqVJyKCkNlDDkHxUUhmj2l2JTCNHL281n1e9/H7lIKQay
Om2l6BKOHb90AuHu+XJz4TIaWV6Ag4hym8AiQVFcpzNiAhJjrSwqP9frnWUTidPU
IS+g/zdZh/D5z960YrpNL4Lm21+r0A0K4x1dX36qOSbjjQY+gjb6JhMCfobFRcSA
IMDTtSGjyXBiB62PZk8Iu6ymJ8XXI+yjM1z9zw01EY2RiqDhJpxIQWWozZxgsfMR
Z+0ti+ndVfz7xJVNDYPymFhEnWoHX9WixPWdMVXkTwrcu4nuWHVv6dfj57ojob3v
jWJnGInFtJDPCaHdD5p6fikftaW96y4iKMibzi6NJzPnqwi5Lb5dZLZSz/7BClR7
xxyyhgzRnTdn2bJHft56LzO+u+7RvRZclDeSAScV8Q+w3jCKrr/lwet4nAogM/ZX
BDUlXgYCf51TfOJ1M2rpU3m/ppBSXFgL7Yzpb+l4SQH8rMALAqGQnPQ+d8QQehaT
oWwKYPnTmhEmwUjNpsWXMGq40E1eprPRdTAKoENG/u61msvqkq6X7aSEIaMSf3Bs
b2trpDHT3XfIXtElA7DYaR4VSJdM/WF0ykGBlhZRmIWZo02tjHQPncdE6rcBhJWs
y793mZqoDlIwYoD1tyTaS73lNzNBq/UFqAzT/I+BHEwS2NEAaeqkl7oJB03H4R2w
1eb5neBpg+xg7AR7RrG+9zB5zs/Gp3AsEyM0AqKyzktEGJDgV9inQ9IvQlc/wWYu
LXr+rdUmqEubwKDSVArWqnSXhK2NP9H4bHcfvFlVrhb99kQQN9x8OzIAuZKyG43c
5gS+4rSCmDBgRPeZqq6uNzh2ZAXrd8EA55Rx5tsw6rUb4gwGGjTr6TQThHPgt5Dm
/yNVAGcVuBgS4hIUv0l0lGLpU97dwNVJiEqudEQnlQwuk56n39nnrTX2lGazB1WI
oZkRETPY9R1Fa1XZsuvS5SE373tWz0iRrnFw4v4vxcP75lkP5fzA78FB8rcuaVN6
WF3QM1iNv5H83KTPZ37YF7m07kxLRJKn4w2w9ADuAFNWIaBRvIvuJVmG0WqjDri6
R/wd7qhLYWU7KHYv3oaud355om2YXiJxtwG7URt3zFOLYT+zCZO/bals1YocW6bw
DCyqX2gfOTVQtfs1Ana7n6UJFnWu8w+3wKWD3zqN8Uqru+fR9peXi11uP+jU1Kim
Uw1YYEsR+foBnRjMrF9+fjsrWJHYC2NpAU/E8iyb2EniMDrZ3JB4NP15DCluelb8
J5nEfrHcdg0JAuoj/adOmwflQvH6Z/pHXYjnFPmDYFmaCHDAYWppmpYtELVMdeyv
Epg3icuupgHbNsrpuCTuV2Ur+/jL+A58+MxPw4TGVKJGjBPzMAsQQ/Ce/L69iM65
5o32xY3axwkhp2UCi6vCoTQCNwEMCjwPnCxa3NLze945JHeNqHMxZNxvsz/cdrNW
feA9ZWgPh1d+CHwWdt6v8kX2Fh3hM7mwHSzYjTflteQcu2HZNWUH3iR7g9M5MWh6
V6Oiv+SMlsXiM6OOlMoMmX5NiHnlMv6VGq/WncAchXALIGZbOsoLecogSlcgLH6N
nJM+zXVgPtG9j/30ampT2AvA1qocL+1cX4+Wl9MAzueclONdIxlWGDOUdHg4lTLj
hcjwgHjGJTTF/XrImeG4pP2pYbgmj8FUTitexWH0y7vNhc7OdEV1jNlSHMppjzb6
PUyz12PY8Q46lf3LAevxXCafejXR5+efsYVykxhRyDIOD0vnEZwdLLq4GxtYFGxX
0GqK0iHH7VBcy/JvuxEjYu0AA1Pg/2OGTnSXhylHRQD/CnSGZVRp4wkwdej3a3Cm
T5PcdULUu2Cu/ZKiRLBOCaDaUYiCzKk0PYb3OFLt8XiFJ/cXyH/gwpbtaUaHfKBt
aU3UijTdPV2TMHSRW5nIcD9APA6tF33/nPC/an4Q+QD44bJ+qiCQBhuYJGUiDjB5
uaJa7LyQgmiCP5cHMO6kHe5/TdoZE6YaXa5eiXE2IPH/vXyVDWZ3CWklgFkAfSuD
HClIZ3xcq5ecI4qg0sVnpZAmhUTMuAi0CxqfFXHUilXNEWngKgJiQ+PBM9ls4F3n
WcubzR+3CdBPYmUHjGmrRetnAhQwUP8VqUibq5qFHYeR/sDv7O8MTYKgbHiJYkET
uyslis7MHdpGdd3yLA+kc8gO1FnbXQ6R/1tlOUu0PJ3DNjZrG2YRKAj1GY8Se8tP
OOrRTBZhpYFhnMG2gvh1AUN/sR4sH/v6p7Th7AM1saGK6ECvzA3QdLV4edtVKo32
o9yZ0DEq6PrKRz24wegrug1Nd0DSUaFLxNW2smQO6zPJZAe5V4zOvPvcMjdfaZpP
58A1OaMDFTpWO2mJ0Vhce7hP3p4szY8fsSLZTm19DFQDNWgkL7R1j3b2gp+OMzJ1
3x8xp+7t+q4hQ90OG6+b4OXh2IqJzyGNPWgrj5qFVQpc8EpywjQG190wds7SHB30
VAkKbWGXa/oTtelLyoa4M+mK+pfOZAbh1g6DddnPYSTp898ztTppv0MxKULxEi6f
qYpiiaTw0jA1nNywhek8VsmtdwqpvSBc2Tr4gEv5IuJ9rknUF4QU2G+OVzzYUOqZ
0d5KghgT/keAy7vCFP727kIkVpOOdBhummMtjB1XeMnAm3MyMByliMWhAfYFNHhg
Y7DeeeWC77Ev76Cq4fhYh8nQLI0c9Rh7uaRbKY4TxLDRCB5qG8E3ZvH2AU8r3Pl+
pwkGek/1bz2jYpGOs0Enoer0ZFaLaFA0mRb3MP1QIj0eDYKcOpTKdtQdDD6Qcp7q
R6b2TZWSKUPHjc/K5OfiTonbGR5ZFLPGWSOBQ/E0ZKtXShIi+ztaVSAsYhUAiXZX
HCsep534HB+LI7qO8+h/81Xc/ak7Rt7XhLAyvyK6huVH2RIz8DKO3Ek4opNEO/S2
+djdIER6DepSzhpXBgQwbQm6AEy5i2RyKkmfuKGNVg/QHTpYi80KNAo2zGx7dj/z
DplxK0dr1w2unB0otPqpkyMwFSb/z6xPLFL49RWJ8rld6dG6lZxnaNbWVlUyjgeX
PGDZkr6rY6n+UoUWejpEIvIidOu4yw5LyybcgqsSg88TEvXQsRyi0N37XuFsMU8r
5rokBFINbePwKGpg1HqDwnZLsOQem3qW8ZsxQnN9X53qkK9OKepw4gQlbnIMHLxp
otcNWvVQTpqkRvMprUgoQI5e6qxDXsNKoQFfiK1PGTHsYocMYgLYysHbHMzJOmvJ
oFh9NP3ur4iX75sAQs6UWg+5VRb6WtDQ3K/YQns5P1Bqg78X7560qDZyQ1bCDRk3
fBOzC4CtMj9q/gv9qsUdX568kD31t1NpbTxGBFDc3v7+q8kpJmCLIZSfXk6eH4sL
vvfE73vPyqEVA/k6gZ8ujnnBuCCWZpTFeNJwAoOWfalc/wU/GiKvlLajTEKzk8yS
DnKhsNNbmZiJnYcZCtCzdgtil1xeaAxltqA71i+xi7aHZfBCeXoBFD4OpobwMrQg
Td3BxtCVE+t1vqbEgsi8WXSj7OYQCL93KJbxpkL4js2Ak2Bez55Fxltbe+spEsmD
eq8xjp01F+Q9OfMiNn6dWhY8UpEejEmvhscSm3NeK4paVRBhWJ0uli7OLA+EtREL
47zU143sD61mI8eOBzarGNZz4XnMz+Oy3ksbhOKEJBup200P80wOg1Q5GPOKooDY
AIWECFBVs1NVEPCwqG/OoGlVeuyB3woiTp+MhzLtHc23NNxzpTjxzMwba8ogchj4
lU+uLAoQj9V+rAnxyr4Xm/BTaPEu2tihfnlUGpRq4pRjJUdzHH4wvgVqxC/FjKGj
ZkUlGscZbVGPOAXKkXcs/Yqd4eeNLVjF7z77gnX1S0G3RX+W1X9W/Ryz/H5fXqHj
AsnNo6sYO6+Vp2q7KbS4NHiuc1neW5EzfsMhaaGsdydonDqU5Pcyz4c7s017SBwZ
ajB0jT0voa8UvDHB979CuyuDq70AG9Q54qEenzaNFzocR7knlJ7DOA1Cq4ea4Blc
lqWd8+Urkc54f7msVH5VJR9YknxJtucqCVDoafZjek+TTYvzkhptHDp6K52TIS1x
h/kznwesWsMo9ymz9s0oxoKzM9Xj1IjoQj5HPygt57KB4dwCzAXkHZY2o+Kp6Rez
302CNdy7+3PgIDVpN5t2veQdlp6weTxXbw0V3zFS89YQtB/kB3cKd1MuNqtlUm8n
Wzz2S/nT4PMgrIIOHjfbuNZe7aJBcxNZ2RTD2/NSUfPTe8RrBaU475EJpWU7kZvl
mhQae5dJaUpT9uVbC/jEdbD8AYaW/694wmOu/K1paXNdDfNj5UxP20V5W56usKB3
d2PZ7DWXvi4KZ8ca4H3DXZ1PBoOLpy6Dz4cqCU6WT32dd6lww+XRb3nFvKBNQcHe
jmeWdKoXwX9sRlxFPNkoyDC3iBbjLQW163j6KWGMPQnd8bjqd8b7UJ66s461nD0g
Dco0D/T8Uy69hDfQ/bQESdKG0TpgX0TdYCZjsDSIQBb4GIc46OOMxvkAfrcdgqXN
1v7BrabLYb8REYI2jxzShdF164/DbJHrBDpVo0BJaEKnNYiMMEc28mzGrtcJOVgw
sy+odmZPpQTcZCoMWxmhSx3DwfpM8G93nO+iw6MXJqvYRycvkHny6/uXZdCmGQ0b
yP9s3el6M3LfhvxwVQMgwi990yp83E3Ga+AkLLSCnFxaj9mZphz0ahSElPQDlUqL
UAWCu7SPouFvG+Ng8J3lHbQoW3csQvgwSjODew5uRC52+EFYpyxZB0OYW/8Yipyu
VF43IKFEhElkoBjxc9s/ubhmVDI9XqEle6q44G2F6f/kDmI8WmX0AIwWJ6IImulp
xmG0yTw1cj5S2yJUbwikvEL12oEMRqaXSAJZrmQXA6SWA7ywc7IFPqQ37zZsvtGP
UOfg2vLfmCAUIvQ0331yTho0ZeZIj50eAlGO058FwnLaE/Q/tjJct2KGUv/mP5jA
bhZdwD7/qgObEUGfjbJ50iU/FQLbTTKD5W6W7WjaDZKKL41sSisKMgKXRzqPbog8
eO0pet1o+P4Q7uGjc3yvctEQLf5hXqmyAaixAq8cx8BJARRFFLoe0C55FCOfoXMl
KgO/5aGWKJKdAiU/k5recL4Xcrm/oVdRZ1RQlnZACeS2KIDRchMjczYK5k0lgJul
4uab/wXRh9jOHQD3jIfQ8Izv7XQZQ93YuWzSeG86cxh/Nn6UADDc7j2lqHMX2ZSO
bYbhG6NnIZq06mozZ9FUZDOnowPgwOOaxt8as/6WKROAgqp2HorpW1gbPAXhbMLL
EPmHopm/sDKI6VBv5WRiPHlthbv1+6X2gld5fjiq+5YImyxMC692YhrMRAJ6U2C9
snrfwyM6IROwOvAPiStXWic2hlEJslen8ea8F4cGCe+ARxgrfUdIDNFHbpWyeeLn
05pcu7zpqJtVR8gtk+pVRb8FLhE9bd7PHvnKzj1b5h0RrKXRLdeVeu5e9dw3lS7T
fN+UY9amNDGFLNPrVDwSJjkCY++q5IFSRISOvqmXzJ2yiA5rJaTHD9/uCa5YrUXi
8BhAru0SbXDNYNKebXyTw5SRb5L5mckFRWWYs0eXc6AbL97SyQWV+Gfyzx5Pmd3K
VnLDcqmneJOgXAytSMPHXblKggHqBP+hvtfpZ0FteK8/2dGm2erema3xDs8xXw2N
/Jl7WYOMvjXFjoxh3AdUluSJcx31TlD57ACu13DDjXc0n4ABwmk6gyZBp3fRpnM5
9YPM+K2UQzN00XLkvlAgQBCCOBjpiyZdJ6oQGUciihwmLZGZNebV4/muRWdU31wn
AZKzi95oZeuDLROTe/9Q+DgJN2DTPMWxjUs7+bZ45EnvyNhVYf+S1LK2UAk/GpmU
6O5009o1hNE2nAX21yf4xSG4EvgdKt4u2taijm+PN37Xtt637s1p8LylJc7AY5gw
TgGyhVO5RCBbfMJ51A9VqwTawjV09tvubedA05LQEQCyErZpEzNaHjVPJvrqznJP
bKQCNVrceux2nzdf4ZOMMjMhkrBFfzataOwBPcM7KI02PDKR57suzz6ZOCED0bcP
/xBrkkc4ykVnk81uh2CfBj3mLbTELteu9G4T9ro3TexHPT/aAVJR2P/wr/NDfgPd
rx00xMZ/m1E7N1aG6r9S1SbDVI6wJBdw51mYYmLSke8LTwTo0l9A78uEXg/axseN
9/nycq71UEV6TeAXS5lOAOnE4UodMG7yk6a6hQcWfuibWT8pDRheXWNIGA9F2oK1
Eu7qndju4u/h9QfFYd33P9hDuJ/xw7YuEpvHw1Naiq9PCRtHwo7UpQU8QLX6ewv6
jXjoL+ivGtWFfIfAGQp4PZEsZolhYXkjwEX7khqWxlzfXbzc3tbzssBNyNuntKpo
H93F59otELegpkA9ue8S1WIE5s1JgS4WrDFBbQ86YVbA3DykRFjT5OAfCnjRScSv
HZWLGHvfXDzy7dpHQtkQFIP1Wn5gFwbTlJB2rN6fig6LMJ6Npkuf3d4nSEqkAAfw
3p2PANBZBs4tuLWaeuy2Ia+UE+7O/yPtXXeNdFvcLdeg6RvdldEr+FoMdjQL5Ocd
uZshA9ttEv66lHgNA20+Bts7skwLM1VL0rBnTQEK3UxlRdrdJUWfVCWMRhNNyr8Y
bP3T/PQuHdtAM7VhBX2URoomL8XLtBR3Z0v73xaHKEUy3qAvD/pVkpn6YDZPXs6L
X9/U5rW9WMPXsgf8+FdrjDlzQSj6qBUv8/OET1nZT9Yxl7hXu42zOApKUln5oHJb
0KOs8VqOs6NzSNYtgAXX0i0aap8ds59KCCZRMymA9819SmIyywQoMmDk44aVdobP
gK47FRB1JGDaMMy/LqArbAWUNXN4/THjftNcqOl+zF3ZjIbL61qgVQScUqO5gxka
NRFnV+3l9lXMDA+nDuzp5PCR8pBY93rox5iSA5Qgm0SbqIyYzMTEfgjQ8xa2ct31
FKZaRJf5mgbQG/viWrkOga8jPVV0nAbhlIS1QSy471AZw5MBJeUAHlkMkiCGoZ71
dMUC5cMaOMham4Z6I347oK4pPfim2cT+IhpPaXe0jenjwFrUBlQBdfgpS5ymNEuC
/5Ia3VQvVVI6cldue9DnjUiE+acKiDTncUSE278Uzmoe1BgM1leP2rrK+OWerpAF
u9TLutBIHpNzu7gUS+Cla5Z8XIqHlXH5UjNRKCd22lmuCUZ/xXDPOGlSW/UJOf8g
WP10S9sTu3aKlyvVozVsZ4HmQasSqhIaMbivCxdk//VJiyKd2kYUl2NLRe443qQd
k8QTiGFk37I7jCrQpvq23/i67IBF3+UXhZwhzz0jckhlt3ZNrRkGzZnonJxlERpM
51cVgQrx+9NJuWRW+XpwiOmWwSNR7EpoKOV2dF1yx9CHlbmBk1Db52Tv1rLiNjRn
jGpVXihyqpl9/hsKzP9Tkl1OUkseGQUpeGtz4e4MPq9T6pKCsQPHgePLfGR5uWsL
zRoqpohzIIdgI8mdyc6jji00VKBQRRqhsCYGmVKNQQ3CY5liXbEkJzuIvFI8pa6F
s+XGtsJFl6TQAkYjCDiwGbgVUHbzhfP6y1vBv9jFbrIvrMZvjAhgfq3w7yq4OWXf
5r25PkHCs2pLyS9ugWQnEQStP3HKpdSvKmUmHeGY9cEvzY1GQXKaBy6mS8lpZrZU
A2FJj7itarjK6haDSNRTSyPzz+8lAPBUPy7//9J6ukLdE2lqKrZYBeulzJjFMF8d
3uC5hXa4UluIkwmwBdO3ayhMjmreW7Kaw00k/Rp0J+PVSXT1xm7tMYa9FDfQygZZ
4XxxeR7VeYVV3VimBvOwof1AdYnLH9iKoyzj7HOJoR4Y5JMwGFYv3sscr+oRIuwP
G+c4XJrfOifySyIS7WPyN2vQ9RzMGjbNJ+g6Do20Mz7C8VnjDIaTXw/6MgqtuYrb
ogUPmdGI80no3zpacfeSnpy9ywMFkw40BjG37SM49e2A3MrlXN/wyx/vlWMAiEkg
Hzc1lmRslpoiVuwIob1iweFj8Af/HlisZSZQPY3ONhbgmUi3wTvfqkRsJYYb9w/4
StdSP3VSiN8ccjrmWxUNEyRrLHGkGAW48dYeseQe7mYanBqpptWhjl4jLv+/dUiY
0ciSXh5GyI0zMx4Ean5g2NWMHMV3Mt3ftOHtdYQOWVCNbEjh706HnsElCuNOuGYL
uszfK4vWkYmeWLkvIJk9Q/2OOQ4Zo+26CCR1yjvv//s1UAaYqHmKqkd/MsJjwjFl
tJFSb2Fo9Y0/W5Ke8QO41dfHjDWwFXwbdaPd6lDnHg4IlLStfZwKPteQ1bcd7aaf
qcu4ycATlNwSb3yYmxaoKz9CguDCFDcG4UGHP/JrTQulUJd1GQLfJGvGeK6Hfcpb
SHxT9AAa0XMI77yHfrUDcIfouyDrdN5BNs2HbqSHA7NEa/V208R6TqdmMIRxlQBx
VEkFGrAfmSjfx/vZGzowdTbqKKlS2/pQa0Xr/3dmMDezPToR1P934rt4tzATFP5D
cjaVxTUilyd9Bs2swcwk/gVvtuSmAKUDE1oweL7qK2IKMZBeATwWadtSpVxEWysd
sBRFU2XelQkGyh332cs4CE1FYrt19dQGs7cqwDFTovm+Wp7JmjZq4gRzMqol9jVt
wX7a4YNJn2wGyGysPwcwUxfodHixFbntqy4jLOZJzoDajMt6JgMJnf3eeooRriQp
L4zrfUk0ciP82BAdc3epjWc/InkqIz5chAPlO6B1Z+wlTo04sMW5BkG+ag2kNxrz
kpb4LzFMzlC+ARZ3LBBo+4qHX0YyZfvRpfppSyfY8yayxHCPuPiLKD9DB7wtoLh3
WxCm6eeR5rEFssgCXcJuwGlP8bpXggnySz97in+a8+GhLrnJq7uQ+fy6nHQrCaIx
QgNTvXIGlT8ZMpBBjrOMJ77uQXQCrafLxDcYfyINHDDsbPzeQ7xMrgzmheSEm+w8
eZ+2CJPjS/S7Itpw/diSiQAQQX+vFSbr/2qmo4K4sFvBHt7dangpgUQI1uLR2v8Z
AvytIiiY8qsD0iXGxXIIFrfniN8aaxmYzvioJ5gZlTeRtaRzJcrOrHDsMHovD9Qb
4XsMB5W/BP63zcO1TsuPiRkwZlx/zyFhi9zeYWq38yT08aS0cZ8+skoPJ2lA1Zeh
WEEiwhwV2MIUUeS1t2nYVBbmV0/WTF+7DT4Gf55qpT68r6eqN/n6trCvPiceyrIx
fcYDVOhFjFcenNucAOZyk/zNm1epmcYu7MlOwz46hPb+njx6/EpBxGNlYoxV1yK8
qkAUUeKgcMtLIFOLI464UxtTern9znggYBc6snQ2mpvHifDPcyxI88nO9ADKGXJE
DluFLbe6kmgAv2+9Z+jYq0jd5q41LOjt76QLtMAyNHZithzkMBDsl3Q24UYX7OfX
T61yq58Ec7azmTZRVD7xPrzE7/S66IkED8MHLGoqyoGPfNICCK9p+6YtcUGOcynZ
Il4ORSQKuh5vQhZFXLr3lKGJGVm56yNPRUnQUoSV7phOs9/lxnWl77ZHzuswOKfC
JkO5GyEA9meJJCbm6kMPJEuaS5WoA4pTS0iexrejf6c1FCXWxUEh0Oj5CDUZ5sMJ
CDbb0k2PlJ47310NJB9+Bus1t7a9NS0bUxUgx7DW4sRpEJrHO9slGbwgHMvW4OY4
KyTMTCNGyd9+FUr8L8ly3LmbgmdeNmJgImrR8g559WYhJlOX5uV90aZwivThG/oc
lshmYRG8wpvcFEr7HZL8k21MPF4kHAgWK+leVSF7+aoKsWIvz0phBKWs5xUiWfkv
ZHFd8Uz665ef5+rWG8N9jO8BcpXtE59Y06uoY0QufcxPNFCq64Dg9DRjUY+4ejhO
K7kmY4hJTzBi8IgVb1t14xmpnru9jMRlsNT8Ejrz32jwfucfxaXUvG5nTNwtDy3y
O0m1YeabdZBn/oxkXbmla/e+0W5y0CiP1pX4ejUQs04c//bRFcFwIP+tXvABuAmN
IScvxHQ0BhUNjNHV3zjQ/P/Qq53c5auKCP4uhRkjjGCctoLVc+feBw639Z+fx8oV
1x+BOHLzByFZ7HEavOKeRidkxJgCMsyCUXG3kGpgYRdF8ZkBUALecQP518INwzNq
oZF6pT1irC8TIm8rj8EAxfzVPSHp3wqAhaoaezjFCdOtWP6X5314zWj2ijqi1kM0
b/qQwElaISp97zRUI+4XiwSly/Ipbfb5hhGLxX5+B2svr7Hb+z8D2Y5gS3i1Qh67
mFCIf0RINy/QfLo4hFaFO1yL5Oxuu+KesIU0rUCFggvKrxcTqmlKJiR1O8VxgqXM
iJAKcleqJ+6EUjHKzSIFFUpOUeAYgv/SFg8Y676RSaYCumo/bGR8a/Mg5HFLd+GN
xyEGhZgTX9ilZ4Gzg02CnPZ6Kn1NyyHincZxa3z/DmCTV5RehJwwscIoaLNAuzyU
u5CGaOFEmvooVSxm/45Ka4bv8axmNu2P+tEA/GhqDCI0MLfxjfKaQnhZp5YcZZlI
ibt2tpE40Onpn31cHCBJirtDm8CfZJunD0n7Ld/NPnOLAPVBrf1qcewuazQz/9PL
P/TPiY0hWUnFlLahE8eY/dHeyEA6vhTTSNPjIvzuMFUMlGI8Cch3n4C+a8iHkHTx
s4U+quD+qZinENQD7wiyFJTmgM1memO/pQp9EToszjallxAjbbsq/BNeDWDeh9w4
bHWgjjSQ4wHzVTx/XKrIrXAA4gNe8UVDB0zv0b8E5ic5JVQPjccxQFbFCuAunSeF
cLLW/zW8jg+oqilroIRTS9gIluOL2YudYtpOu0xMXNpgFWSqsB2d4KNWn2WiPExI
VmpSlVnmYvwjn7pZQ1CTbgdtkv3WyPicRkFzLVXApqX3iiQGm6aDitzN7cNKJiMk
XwpHgKN5vf9WmK+1wwoTm9ZKdndfqzy7cNWTJUH1sQK66FVMZcPakQd2mWofKpnB
cBmizK78tDfAVewfagkQsWGnYV3vRPgkiWPUWJxkpSxbFqKu8bYtxGBGAcBKJqmh
6qhDJoLV+N/mmfdZNVhhU2eBygB5Afe/sUmvDCgJofXpZQjbl463EksjjDVHip8A
N2YsgQ3MDKBCTva7WsAG5CWAm9eIiW5DjnGA3Jnp55lqYx1wp7QOoervhBsNrJVK
qAOa8DFgwfSWuE0XBQg/u1PB3ObaW8tLv2Owtfmf+GAyu9UsvDIF14YKwWhr1xyL
XWLYQGeh2KufeXV0Y0J3HVDULqqOfjruMkYv2w0bUdhCqHQo5Ox4/4DyvWibbuPU
ssegzV7rP8SgNltLCYUoSSq7Pf/CPiUu7cGwXESZyfue45aZ6+XoLM94qm9IA/kf
11GQ+fRMwDYUWHB6s/Q4AtnF2v/+HtoBgqnQgPQOANdAcVDriLavwU2e3bbFXtY0
YeFQsoGPIUnI/e2TWzGOkbwyC+P7q4aPevbfayjGoYkjS19K2oBJjW1uO3sr6zd5
37opEqoYyrPLbPdMJjF7ChHc9GUrQY748ZVtG+y3ycVaDBvs38K7twcC+M743LGe
2OA0qxFtZNM4OaLwOzzJymB2OYkTiY/r8fAWeAff5BCthd1nr2jVLWxqKW/ua/qJ
ms0NvzLxGfPHJeO3ENLmT9giaW6IrBwiXnCQnG4O6S3H3Yug4FV8rDR7EoK4eOmV
DIqb5mPrkjDiKMTQ29LYmDgD09yJsNnbudlIRKVwX5vIMj6/Ez8nPyWk1yRcdYLA
IZI1w+6U9kHC2ld+UR2adElUUbToaFAmm5s894J0/Rh1WWALDH2Vdgp7wDxPDTKp
6jUcyHq1Cg65UabTtQpC34bUhbVjPxL1c37swJQSjiZkGJMU9ivWrqNNxPX9l0YO
dnF8L3EHpG1gpgnNVVpw0TmW7I+b4mm3G+DsxGRg5EKAmpL64wGXCeSWebph+na/
wyhI4E7j744tk1BFLyUS8xIhCQhMhy3drca6i/swLQdALiqfLyEaeLpSiYSR/TF4
sQbfGPgslbSUb16pVfceZM0RF6BjUMVMHK0ZOqmZavF7naLRWrS0kLoXF+0oF1mU
gMetAlS/eLtyTHvPWWhaX7Di6nySKrZx2yT0vFnQDc/RixgSLMivrBvpRGX3Il06
cbHscA9vGcu3yBCyNCJ29lmsbTxswnWtqVLeiT/xV21mS0FuRsy/z+R0fuTqzglV
ZzlB2zrKXbq96GFMcy7b0/IkZmlu2YAQAJ/pWOdqOW0W4hyP7bEg4hF0n9FvInyD
7zo+2vwQ+y4pXvXCOEtgV2a/NBUH+3+qTV/5SBks6/79KsUcxZy6Ghv/XUwoyRuG
MMZspRZkEr8d0jkwupsBqsRD4IeICWDHaAgmTnHi5pT5hNvP4wLZ51nf79OYzfib
GwiZ/2mdzyQgJ+mewzHtUcatQuvj885NXlMubalH8H+GbImem9+S+xPnLEVvUfYV
Tbeuz2xZwb8kU0y1T/KeosIOHQyntsLJE3gGPmhbG5b3uP8LuUnvb2AXS4gb1MHm
pbtDconDwTfSx33KZJPb6p3AgzQRps+54cycCcZzBEzRoThSFL8SHeQdkeGa52mc
2p9dm0uWGyvMRhrYHAloS1LvIem0U0tlTjRt7Y/NfY8ZhWURmfffhdoIP+Fgiah+
4OWxRRaVIvO1T1bbC/v4YLuArwGj92Y7RZtLDGyVyHDy10E+3UjrxdEaP0YKldtQ
28Prqa0a5T/hCoCKoyRlMp2omhetUMW1SFG7q+ESvuu8BgKN4YCN7favASgRU5Ko
3MlURIaps4t3OlbGTesLZn/VlltvdUBrurqcODMuyHy5WlX4Os5FQgIf7pWTTCgi
2NinuR58kFsYkcYTBjqZhgXvj61grh5sPQWyQjca4bxx+8eJb/ofyRJlWtlMAUfe
63C1XludTmfWw6SA4GmFqvZZnyqH5U3+pKctRRysSAWrxTiEi3UYU9vlFotMAVOa
rXWtiKCEigbaMnrsG0yXAMfrQGEcapMN12wGqMulRysR9B82t/mCgojGwq54grAP
qgwbSoOZ+EDRQnOAoTGQCyxUD0w4bu06n70mhmi69dB58OEnGi/DXVFDvKuCYjhb
EGFsZQnJVlDx3F4Ad4TYaT9jZPGCn7i5O4muGVqITvuUo1/4Q7pqrJVdu20YYKus
+9TNvbgOsRKREpYMikMn55L9R0BxRCA3RLQO8hAMqPpmS5JttjqBxlj6l9WJ+hb6
QGiKbsakh9GelGhQi4mxhFttGtr1TADZIrrUMph856Efj72Jp3f21GPaY3YBWj4P
FPeZ2td6MgBY7OnuQqvjCL1RCwCU0kAX2wIa6iQqPMQk4YMT9iw02BT3+3D2dkxL
8oor2Y2/QjusWt4n0StKqgmwFR5HqFDVALlQrWglIL2PadEEtOvMXPH8AwlXeNZg
N96JUNbXU4LU3erPuC0Yv6krtTEPiHaZo+AwmiPJ2mJbDaVFvV088Xt9e5odBCJV
lkwtqGGCOCHul9YCg3mwQ2aVkeC33BnrNlEiA/ZI0HjgZBMcN9PcFeUk3wOb1FWu
JMEH90Vsvm2cCuTmtySQAsk5HrmfkYQBNSBLuetxpz9bJWFXXGiSFlSePwwDjJlA
t1CrLRzBmERvgFG2rbW+XznfPcWpf9GBX1numqdhzflXYkvKYd2Bgx/IIKyEQXAc
wdtiz7TNGOyMSbtCNz6JbndHrLF6dSUnqe/n1PlwmY/sdAbbTK93gdf5g139opKk
W+l+qi8eQoEh7GqMUQZTn7QiywnnfVNROYtAulhXKZ48SGPKjxFLGNeAPPrX0kiY
20sOjD8Rib77oy4nfUvchCwLBFke6x6uthDXdRNdpFiom9Nen5Btj0X+l3d0R80V
FyA85zOl+/W5Shkj7nWmqvOEOe/Wam+AZZY2OcxiMN4b4XBlSlOK7h6HW8YP2nSA
v68dV6ZfnA1ljovi+uOuzB8CRFIwgd9XdTUYAhlJWS40xgzyeq4Hns1uYdsfRSfs
jbnl93ny5YnUN32wGQTKUnNnupu0xHsNApcw2v4kcsp49iYSXfrWgaRTcm6msoAH
pRhP6wpfufqEWbzWFOGCm55JNs4/sAzDmTZN9vkg3uesa92HrNQPQzJhJNI+l0Jb
yB5W38TkqJ0h1JpCzsxmXmXkYlusKrEUhq3n9W+6YMM4vcUUBDugVE7wO27+ieUD
CWVK8vkV+jjse8+uMJtCDS9U98CQzP326pkwZ2b1gM8xvgmbxkUGw22rkVDoPTyR
VqeMnUr5FMOsiWN4A86gUVgfX9RxfmVZB0BFMuNqtCe5LIN7h7V+kdLTTyl8ba5M
SokQJpMuuczCPTBKi9T6jSLXob9+nKOfaG2o8iCHbmyzQTR6ilrAOwPRwUU19b1P
G0b3sh2c5tC3jeMyM6W0uaiQzrRQtu/ouxvtCX+Sh7aQygSOlGKCEhg5DQqhr34r
TtLTmB3PWF/9PVELymgPslR/57PCCejDucTwbFVcWX4tuIEMNdV503Q+kHzCGMhl
rjizTtlMe17068tQzkWAS6FsIm0FVbTZCFt/Min8IxWQULn8GUssaMpnQu54BQSq
UiTWl+gQuWRDDcrYuAZ/ZS3FQ1yzZ6+F0o6Ae3Tjg8liuVAeI5PPuCoZbmuubSda
XlbCnDh5BJH9pD9w/eAaegdkSRHsVwhqq6k6MSbbjrCbHxtkndUPHLqS5tfqJNHa
XqujTcPRpi15HPpZZYQZolyYY11LQMtvXecRHSIHKsNF9URXOFw/AqzIpo6h2p2j
O+8GViNDDwom+3EgMHdvO44fqHWD0ZQcxTvQz8W6LrFfvRxU1dpM2U6xM6PNvUBz
+mjQhELQyaT/ABAmGwYPiKbZslnSBDqzOOlaHyeDsxRmblqYxQ3YCPbdWAH4Jc+9
MVO9sBwSsRvr1T7kCQIHASgzJwKNG2ioalLkZNHIqizvhJA3YF7L2/J06JeyfNfY
U74znXBW3cu9P0S6AN6m4vq93RdCOauXvng6Vi5C7tEsdJnMRtXUrEzFvXN3ZgjN
vi640LI22RxCbXcko810i9qhjICRwjGLxcWYfC8YHQKXB7XTvhvdSNtdKAaYyTDr
5YCBfSbm+7mP5vEQrp+Bg/5gIwj2zAUn4hPZyWb/K0O9tOhWk23mNIHQfZmErhOH
IeU4uFIFdwSq1amzLQI18b2J9J+OQwZpH4C819FlwZzFWFm9RlxqFtvZUs5I+wK7
+56yMsRY1LeaOdfDee08s0qUmZgnIu9+H2DHCfxwA8gNX8VtKEgfNXozdeg/QCDV
FxCF5Lob3CEIZwIz+fW/QYji3RWtk83MyUWrnKHJ64VimjUYzFZrbWPF5SwLP0oY
w7WYNQCalkXrkLJqR8zxSCoDOeOqY4p3w8aPzHbGQZljmFD4+Pf5Pj0gpgk/zx8a
hEpUq8jCk7FcAMRmQDAqESY+s8Zu9wO72AlovP+1ax78ICy/AMJ/igW3+0Vnb6BZ
wGqA8dfveKClD6SwgWlRkG1BhPth6xpn3I+/KQ4+VgnlNYlnNCVfvHfjvJSj6dJ1
O4x5udNlORe8NbnuS47qlepFG62KWFvZKUBnHsu5cv50Cbn1lfywWly7kvxMvTiW
3q4DkJz1oJSaciuXLhamJwKQOfL1YebWr9tvipAumF3lSpGDChdJXEmER5+7NVTa
3Okaq5BB1LIsrTg6XDAUg2L36AzVw8YhZpgcUzJUJGPD4o4Q4qvFjb5hP+I0sJrs
5nGAjWDbIoGPnfLN0f77iyTntXYcz98YaOn413tPKyuUVwZJjDhxRH7Sd8Sz9C+7
Dv1ClxIQMR+fO3TVlgtsSUb2JuN+PO5Y2S3L9ZbGL/Zz+BMmtrieCkgIWzqCSFx1
jMRdL/2k8nyBYUxxO11GSYJpBDLVTMN7nL1MOcrRqFOnlRm+Y8DTZwdUqvPwYl5b
/BkngkPXxStba5OnsftkP8vJ0DCRC3LQFj6McanmGRbk/bPnnnsjS1gf2jPU/Itf
0tsA7kNVuiSsBVnXh38kkqwtItBAB0kUOL38Y/k76LK143CeCcx05hepNBWIWGKu
4EZJs+uQ8LlFwxMFcYJ93/b5lDV1h3d4elrBqmHEczd4Eh9mXnfelIKx+3bYAucP
FaCHD8k3CbJAwWOXJfo8e2ClNkyMtlFprV05zjodxUnj4x9mSqc/ojxSKLKQUE/a
cYQPte620/iSROdwmJg3gM/Qc6+QcjKwdtIP4nAmsIbSwX2FwC4Q3vsnOraa3c/Y
XRdKoCES6l8IriAPVRjQB5v93yT62mMslQM2C5d7NGaFnvCQDEtAJb4NyVn4zpl3
IScrwq9I3Af5AHkZrXDOlpvE1FeWchSP79LQTFdMK+ZQfYeV66uNehCE1kETUWM0
b5DX+0+7kwduqpze0lqJBRY48vctxTsdU2W8LMzifGkQG2JWMgLh4qKFUzH14boI
jZ39PIKbpIHc7xywEgZEcOGZB8PerLaIstsUc5RXncIdyW8Rc8Mq5lxJyRnXuS9N
KapE9CnAB8eSrkMjjayURnZQeZw4rSVQh4m638OrCPmKDMwVkYUxGmm+1+kFO32E
C3Ph7Utmtd3Sy/fnVmxwKOEw9KzA3xYjElOxzpG++WTSvxh75KeQuB5s8LtVsn5j
cCUGhqy8ANL2FWHMcwQ4BPLkGJmYGh0y1ew0OgWZPtTy3w2mMqS9xyzXqeIeng+f
qqwSoUTjCbvvWtcl/MYe4j+JuX35G/JLo2HkDhgX1IKmsYglOtruU4TlkOP8ALvz
APRZlUbKQ3OxDBKMTL7Z4sU7jfgJPoldp4RvXJ3OaKRK1aMlTbUY1LLOMnw4ytcM
3xsoNOFOyOkuO3zgu7qQ7ox/qBs/55V/W0iWzq8c74hm5jDPoJM0bJXm9HxsI7J1
uQRQQNxxtw7i5Zao8jIu8pgmZsLUDjPbfxlcrNFhGtb59LD77kLq/093R7hqccOV
/FzCix+vmn//i7sXK7M5+PBMoY/8v9AXea2fRF/x1ccA/qKh69hyJnb+FHfd+n1o
zNW8PTIU6wzb2QvvF2JckI+cByttcmSwuLEez01IxwFZshO0RrWq2bYxDIzNo1Mw
jEO1ip8RvUaDkmbaoXUbWfv3Cu55j1OXd6Il4pZVQHv/wok049dNI8B8OzsEt7K/
LyGiKb7btErmyE261GGA+0T6AzC+QMIhjZFKAOPvHR6sm5ZX/kkZvdlq3nvH9xpL
NZz4PazP9zlGs+XM9ly2AFo0H9MZBvkfoVchYjZdyoYt0yCytUzhUbqhzmUMJsWt
VPgZfwzRGp3rUHes9pmX2YLVJvMpkC/zrx+ztZb5ngqn3K7pvDkUcQZCBfYY1DMO
554sk9PX5pXI5+Rjr8dl/9aUOi6so+XCnInEP4wb8i2wo4xQ5Ehtnkm8juafV/GQ
lu5+ahLyc+SPpNZTs+Aps+ObLlFqOzVM7L2EWGMqOL0fNOXPDM1lqM8IkXTPDz8c
0X45q7NGIBqVUPIxVv2fA57bLewW1rT9W5fAhDC7DSekAJlnE2HGw9zlLkXhoYVB
nrNbOctYzZOv7DcAxfo0p9QyPAeg6qSYfbINJtepDVivzzR517qSpUK/66abVMMo
iSq/bWAq9UL7TjQQmk6K3+Ws8ShiXaf6hBb1h72DbgLNi22ME6Qm/EVSGu05WDs+
SFwg1SQ1QoPpiDMusb9UI9z80+d3uloB1xWeDoi3Q5xkqSMUdeULOM+cmiH5bD9d
SfWeNY5vUzLhwA15LSD7gYgkyg6zPUtyVl1fMYkL5G/abk4bpZFmwpR3whlaXlrd
Y3asOjX1wyVUgD9YbWrb3Mw9kDdKW+u0Sivf/QlcoBlTkYh6sp0lItpKTHhbGvHp
g/4GCAEh3nh4rhVLZrfpJs046VrdGG8jMyGfAMkP5xV/cMHK7McZ+EShT31Wavhl
B6SfmMxjmWq5BLWl3vow913Ijq28G8n3cjDHz1avl0mGYujpYi8gevKefFNBE2lh
icq6yOXPHbXo6teanNwKFHyXlnTjH7TEEpGRp+KDd+bEDTB8vXJfuiF11uCpgZmh
uLLMFSoIEMA2GDt1Ueh5rxduHkoRzTTjLuVUfefUTSLkuF51j6FUw1iuouMK4an0
nVaNqCw6B6ZCaUq3254rGZ6WoI4KpIyuwqVVpLictUMmBMZ3Snx2WJVXisKE4mb6
+WLhcHv4i+mFLxLuWBS9dziMGl3p6Vb9y0MO9WebtrLWjUrT/oAMhuV1JDSiu/Iy
7MbofnlmZGA3hD5ftPI6Ba9MljWB6sRjtjyNRBO6upNmNYUmupVvKHPeb4/1iSJG
Uay0IaJhgVMM1hEQhnbUTnEmKeprem53hiSpydGJWRFktLOJj1o32fI89mfcNN2V
9bwcbXVZdps5FwjlLnZCxHcSZjQL1y7PHqtdLPNfJqf50h6oXibw7UVpC1lVmA4x
nPIgsmdRQeKu+ARg4VyEc1zV1/rZ+5OudVV6MtHPbK3ZqRQC0mu6+Z7BdmM3nfit
acYcg3590C3WaNZ17jQ49w3EEKZqT2xq8aWimUlRFppUoSt+tJ3gPZdRPa/x3VdY
jgCtptIbTeK43ovzdQv2/k7FD7qPzgyCBaQJ5bv6AMjaKpirpfgHQTGOUHBmo1F6
yTmQI2LA+3MVUnBzhsA/GgzuMeUT8UCxGusWEICdTbOeQRuGxMT2VB09AxEnR/5D
FIjgf4Fp2nh1i3kLKKuFHZoxFjuFgQKjYk2ZhZ6MwqLDoHGq3rGfBPJYTipS+FEv
4N5CuHKKNXtzU9M2pj7ggcXTzba1JKve1Ws8VHL612v6tf5O5QPkYIIMSKLtFggt
oZPZD9RtAfssM9sbc/9VnEsgKFFD6rln9cqg1ZHPPqzrC8zQvwHenBT8jJBz3WlC
gDeHTkBSs8gCqFRy2CwEsc2AOFkquKQN03iAGODRjG67rhMw4IfKTPFG4o1FZBjP
GNryvmTz3Ue2HRyZc+IOeac2CYPQ2PNL+RlOuQ2f+9XuVxzg9HdMWD5/UCh4BNlQ
E/whPNy3VXo5zn+1DphmUATxEEA0MxDuDSFbwPRk5+jACUUjhm24vYROPh1bAtov
+k2CAoHlZ5U95dAxQVgLKEVVLFXwBxvJN1XqsCc6WVZXjBInaEg2+1+QE/P7onKX
PPsnITiVg1K5vVpESPaIsnibdJbbO53eKinYObIcOor/a0fTgAqbXXT/nGhyXQnr
gv3U7ldg3oIxWJTr9Kzh8DZMwp+hpa85D5AnjY1jDkm30/8tnOh1JXsGQrGNmJjO
rzfCz55vrm7eu3kIuf/dKiyiuduFSlVfgUleeiQDAcC9AsLX+PUGdRCImL1LHPUn
I4CGnHHwVprw2HfiuNdVoZ0nn2R/u9zQQUT4fc4Rk/6imzy2hIFs2IduBX10wqNH
bjUGX1rQup/nmzZ4v0yzSkW67/Cbb3xPq+kiz94ZWQJiXSGvZRXfc2K0LbETtyzc
X7tRkyXhZ3PDAEkClR9VPnAOydhXazl+dSHm3dSizj0iTCMfzMKKfncHWUKDK2Zj
vuNZX1AtJPdSH5hR0r8ILPiPv6CBu8CsW9qzVa30IqgngoN767anfvsbsB+asYBY
p7l4Ycujiu1l9Uc6zQnpyW5FmvKNax2cbuOLUCe0ZRBw+rSBd1DIOm8hCQEjwq+C
nLAeUGmnBlDyR4ITZhdrwHxBc1pNTNQ98vMRjJcpEHVfymGBvTiq0CJb7pRzeRBc
y26bv50z0Sg8AnSsN/WNe6SnXHvJe5BbEZk097KunksbmL5APo1OsGuvRFcoGIkD
D7gSyE7TUY4ChSra+McBiZYBJoH9IXUmdip7ArszjpIPazsGrPXiSOMwU/xyChf/
0PX8kd9DwKE0eV/iNHzZN56NHfD0xclGu04VOvu8Ci7h59TM2H10BNR26682EYrm
7aBP9Tyu49Ah0JE1XCTSeCWQlwlG40+plMbYP0TCMz7MFl+ANV2kGehrlEy54yv2
gDQOkwKGr+anmnwQDrSmNClaChyquYFp0X1+XMgBOhQQBrTcSLN8o5moH5fsiw1u
85BjX/tuedlafmhutHBMZwnkuojvMFfuET2BVpXzaPHttxFdXNhBVswxeL+WMkDG
FvTQFG5WOHIyITT5lUXFjVgpkjzCySWB7AnY/j9xbRgJFU9lgnvzutWv94bjJS7R
+/PUP7lIuUpkuKCSvNQuvdeS7MjpVoDax9hsbNWsddYqQTUJRgJoIxXsWEFqyKUJ
Pc9pisHEoPXqSIVGjt/qM7znGa2fRQJz2R/iBZgTWkIsSuedukS1GxyM69Z6YYVZ
HMBstyCWK/uCZZAqGQNd1SJ7Vf5UHqputLW96rD8F4LjeC2gYHuERiJl5fm8dw4w
rxYHuUYeluC9AWfXyjb8h1eLbE8TWx+2DKxWeKZs1qTN5jpsUmY5L/PR3aRSzDOk
USO0ROFxZL+VfUas5Sii0yUJ3BtKlkxsDn0YcTVG8S2x7QQNDUb186+yokP94s5M
TpGlmAyGtAfKevu1aB3X21Yv2/DNYKYlzNl/Mib5mAC4iqCY3tF1U11UUHTAeYhd
uAR3f5aPuJFLzfNvD+xWcaSaKGzTFv9XhvSmpqWGAgpiioRcqsk8C8IJaMLXyu0+
TAPd+yvhZY3zvza1e7wVVYavBzw6vsEbbO0Bi5cGE9XKn+GZcxQX7kcaI27bxIsM
2XJt5CjkjRpByzcle2uTzKA4so88gjHQ3Q2ycyAjmGsPEPKCH61HHdamRDE+zoK4
i5b21N+AIhrBEzHpg3otGhbMJE0xHlwt0n2XY/6fqu7U7twgxlIRSAltUSjwjENl
buVg4lsLuumpFWQFj15XOt4M3WG7vJwxr8Ap54PZ13n5TQmpdcX+VljV2pEmrrXN
/FWLz/TB2cd3nCLF0tdvV0anAfaRGYHIdTqsTau9HoaV0URuYM0Bzf672A0Jk3ld
QBqdD1IXkpcS8QKD4ZrmihSNdQGYX5+fCeoRzrvF+WxRCE0rxdzTsPYMh8iYEPXp
pLFEpQ3MEXQXSgthMDBewYmCJ7ox+/QcfidgbB4uRZd9PFxhNYabLPfDw0MdEeHI
GTZOKnQPODsr6ML3m9YSykUb9bQhsWCPDbyNIJfiF8xlBlA4TupGs4pCCDBf3fVd
3if2MaqiD7hRIt70gMstUtS5ZRh2Zrw57Bef8Pp9b6PBqnFN5ZVjujIb2VMTfabz
jxFb0OPKtx0cdEgB+h6yLIiddALpZFnti9XwrxcgsRUC6XiwwWeO/cLClggxsFeo
oUFauPmOFDjJAlGAArUlMZjsJtfoV1mOCqwdt0ewi/jYIiA6OzBdSM/V5ayRqQJn
9dqDzo6G7EXKGpT0z6WOa09obDl9HqMMR7zvwVn9XhPVnZ4P4Bw1oMZX2g0hEvwv
EP4WX9s7y9jNGSbWEmfhLa7NmUILSZ8/oCRCcxqNxBh3Juci7bjR3Y4bv555lg8M
ZNpheUwtUFd1AIS5qy7N9+2RytPjREwokHk0V2vrzxkHPNTc7oXZ7G6Zd0dnxFKI
RwDHTJb60wnbAvUOHR5Q9K0DqVAYZKIPZUi5SkBexZtDCcf3Ae4uu6dv4EqHFUEv
kyPJziMeqVlz540CLuv5Ptv7voNtoUhSpn1TZPLuhgd9GFLOm9OzUJlaqtD1pDIn
OCO9tWtHaKeHCZB5PccnXGkv/Rs3kK7d1ZATZCJ6zlseh6fiRDWEo2ktoqYpA2yV
oU7rOuClQy4c4lhW4nssJuaABCupNB3y4VzOeWyPuKyD+TqTKfUyc1whiOcIZyS+
144eipUcitqHG0RDaVyK0vVbFEFpes57F0mLajhaVZhR+bpEM9G8wHPBMQDY1Bp4
QpqIsyfeDDkNwRIYjUiAq80R0LaGeclxOlwGzAF0iZTYDgWiPpIW8BaKjo90lSzh
EkW7j+2dlHd/d0bbuFJ+6fO8RW27DXUJNagqzgNXkf8RyAT8N+fmV+mm/3TbngPX
c5euhuKxpwc8QjNe4WpCMETdePs80jvrCc3ccs0RNu6h/2c3DUrOTMNulpOgK4xf
/aMtn045RfCBW5UGKGTwy0nlvEtSx1OyKywwHgo0xHeix6VZUT9QXsvkpv3h5LmX
JMExRqygTZzbqZwZNzqt2wv2nqecAvRtJNmbspYS0yK0zZfHWCy1UadsRHi7ea9+
z5zrfySLaq3XpXWE3nNEPZ1uegI2Vi6URUneElOX2IqkdrjsFiITOflKyFbgdbGV
lGTzenkfhhZzNxuydUS5qUNgnploQZlz2PaRZQiDQdFLxp1fT3jNKp6sbrfp3cC+
CwUgRxGPW/lqJ8zUej/mdgp3qd4QFLYCtCNSojYvj/9PybVd5uM9RiyRj2MK/kwO
qzDB5p8uoKWaNPM/EGiAl7bIG2zdfY+eHNgAfX1x71YvLUaovPMcepY8rVHQ82Oi
GGkdDJbPZ7yrmN8KKyYrifa2FJjxwyTpEF2aab2on//fZge1C7bFgJh/QJ8DyMmL
pfJglA52J8JLFPDNYN9sT/8xr0S5Lt5yYfgRLz8PVUIhtlzH1CAVtVQvtY5jiG5M
4QBYbm3XEL5phxkgGqXSsy8JqPXvvC+11Lohn1MqxDQBOZRW6erKUWz30Ca9zHZn
+2YJxRGgBsivGxtyyQRp8Ba5++DcBiHqnT1HQsfbzZk4M7d7CDzRUt/chEEIi1cv
xXfllQKinDUbA2fhSam74bxS2Tegp10AeagacXD7RwcoJkiAjbj+e0W3H+zKfI3Z
W6NPiw1MkKxMd3ur7wrcEI3VoLokXA7D5oce3455CL+afxtVFXDBBueXYw7xURgO
r8iEXCsncPoI/S/SfAbQ3K+Yo0baYjdmkztQO8LxdPW2UuMDmDxRvz2zSrIG9zi3
+Vix7xpiXMOMKpTsh1v3zQ8tlrdgLJphS/SlvgHwe/0VRQTUmmXspGopzk29mUhT
uKEiF6tCvdxSEd4YTQn7L2GFZtBmTZeEjeXpu2+LXFBVKo4+8WKSHhaycyPigT2C
1hu65LdtA4zNT2cqMcQYkPo1dO3z6oOILPzzT3Hq+JMWCHxkA0ils4itE1TVHgKZ
lhTCsljS4JOMDr7Iqn2s6nd3rINIn8+0pJb6ChkddPo2uPrvn1ljADXsTHOgl1a0
KkRML5/+ffhxeeLN7sXN0Mw/YXJuc6eukhl7YvMBMK8UO6zQZ1BdZItQDKehgWXG
lyHh053ZleIdrAsU5oDaXqEx+jjgPSDQM4FqPLmmF3npvjMfysEdtDrssvhjXL3s
1A6TrKZ/LnW3dVKGfkz/3dvkjGHk+9stty9xqZY05/ucbYN8/s+CB3Eq2PSkrbQl
aqZ8GrzpN/5U0NT18H22rGvZjc6g9ysSJmASWcmYZBGCCyvN+H1ChbtxSdKpjO3g
E6HavOXpl3dq3APmKbwUsob8EuqLOcVBnp7iEu/L42we6Uemgn2mnYjirPAFxdY4
4UuIKA0LMNY+A5smnuiHn9/58TmqNnIdQ1taJvjYYpvBiAqiG9ju14oPySbcLgiD
CY6mO6UF8olN2OhfVS789fXul/iQ9Q60tYJtQNxsGLqJ7EJ47gpYvxi6PGtv04tH
MIQgRCj5Bl7rss+GAPVb0dshsMAd9LPLyVqBJoJzAt/kBy74OE8yqCcNypC3xyfs
OC9Tc5SJlh7h+LaJNhrZS2+gW3/B0g9M0vMm6L0LOcVMKxvYd7ir3F5s1RCt0u7U
l0fZEyqfQjMeSyVUCh1ejqLE+taq9BW8DoGaEuno7EkjWJumOhysn1jCoXBnz6YC
Og/q79BtZ/K7wKm0Mh2c94IIltGf+VELrhdejEvesZ9eONcZ5UwGIeN0QDvr8taY
k7qCvivEiZwerUtu4TFyKGX6kyv8PLMGd7Xb4ItHZ1AYU392JgbDfeyOE6HoPLZy
e6AyuO1uADdoBuRR9/E+yc4apd2oyw8snxudro+XQyISpIgwImiMXhJzbHARmkxg
ZnqiGIjpRb8T4m5c/iptbpz7blccHN6u0klA8p0QnroQO2SxqBAXrdyPmKWlebKU
HIXzHPM5z/GnVUuYy0W+JG30sihEj1dlLh+WkGRIkBUPB69UBtpeBmjQ10u0/PEN
7MoFkHdV61/OVxuvdIjA4vX2DEVkGPVwFnfCR+bm3wMhuH2rqjYZtSYrwpx8O0QL
ua8wqGr7k90tqfCwsYiHPA==
`protect END_PROTECTED
