`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VOStwdKG+7vNTZkJ0MjMZbCXJ/21k9w9R3aN8YAyiEXr3+j0vqwZrfp9nWbfQWOX
lpG+mMhxtNhjShGEHdtDJagKALr5dVgGyJczXyrn/EGTM+QOMvADzN+hfXkTCsTC
FgZfc57TJ3OZmyCcJa3sINq9v8y+xQe/L6DARBXXXJtvWulbRtJVdq3/QdFdKlLo
5BJrlf6FYmeZl/VsDzk0/Al5GVQOPCyPhx7Avv3YGRsNDYhwfHEs1PoxcecvV2pb
gqekN4uWPWNTsL41MXfW6vWAN7n/75YlMtfFzlbXZkBzVlg2nPvNk0QKBr0cXzWI
hmmZUOvMnItbHujl9vJY+Uy0EKRzvrQjrZA10E1rpSCopek3HYEYUT78pbvVnwR9
6XrmHNWWAy99E7nH21W2ZlHbSIdyDvhUVgfqg0na69VoKy1NJlvsMSDM8JF3rh79
2pJQQjspIFQEVudASI+zR0LWAxCVPkzcz4C0x+NEPLo=
`protect END_PROTECTED
