`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QjcFXmFEk5TOak+7AHesOURSg0EoaxwLK7ixut7vz7Ktx6eicviKWLlU1bkyUtrh
PF75rt4OrN2JNyD7oCWAdbsCLGh+KI9zb4ve08UgUjfKfW9ir/MWr0/+0AVAYdhm
qC3q9+JDbS82pEsx2yZ66hbxMt1a6boT89om9/SSK+fN3CXlRbG8vY4uraCClYDX
5ynXEk62r0XeZTRcv7OzHc+F8wo/yBFSl2KMKENxj8E0m7o+Lqe2TSOslnEArDys
Pht6o+07G1YPsEExNK5XaJ7oaIjUmLXQ2CtckNNqkC4RtWzaESuX8cFBDliFRqLe
CUGUiHOT2qXcTImOjWSb/dMFmgSkrqsPWjkfCzslhnqEszXfbOxm+h1KF5Wv62Aj
e6rPh5Xm2GKdrEMvFPNpRtRP7QVQuf8G7viFiuKJT4kfZkFbZMP1ZXoHqOdHX6eZ
8f1g/uYEBG10lEXyt9ZTCHiEKyckgisf1hQdDkiiwCKoo6CUL15CGNAkl8p/Sz0Q
3Y7WQIEcissdgng/5nDQaQ+zB3+J46BnLwl78wOY/2yweqaFDPwc61YnOWr6gPe4
rNORf90pTS6Ym3Hc7CgvNOfg4j2YBr1WC0zmnjnG5kOBcCRVbp89dyoY/Vey4LTC
r4++AqOpxoh+/Qs+46+oaAUFoMBobzBwwZS4tTpb2PS6XODlpJSyKBDFtpLiTduU
pmjzSFfHXDmMiC4f6gsB/WcZ23p1Dvk7wyXlYWP9Efu/9DU6WsT+HO3RDo7L/psd
YBPEDk8OcsPZ6In3PmYEiA/OwajZvNySMez4Kt0MqNgfpBvVafkybJ01YBDO3Ipz
leSgZDYK1PS06HOmJyyd/gkW2S5/dUPTttUNwbVyTtf+sqINfhFXJbHg/W3jF1ER
x3NI6SqMfpoV75Jyh7yTIX3TCNFuej/dXMqrG7/VECsFn+/NdtUhLEzWEwS9Cshk
TPYSiq6jQxu53QERenKi/ULzU+Vd2PRE4osobbvMxYmM18SdG8ZknTF58EXz5H43
/dT5cE832/csUnsE/mEkBUZI/Qujo1APuPOE5tdTwVAJK8yqawUW/BKZSfLWaDfe
XTsXPtivs9U3ua0PH1fXMA==
`protect END_PROTECTED
