`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SR4zRSk4zFIJdun8BDWNxdbnN9iPoWGp3r10JHIXbwjVvnh3nscg2yehqSdKXthc
LKHgTno9nyvZ/uU/dTLH4pK/TW/KMbRcU5Ap68ydEOV+0tCSHrjweoIENCyORqOU
i4TTpZ14ztSqTKGAkZQLj8TTaR7pnH/A7ifv2ZscjYoTEvXdyzxgnWTRjJ1SOUKI
HnWn9gJAdaoZ4tP12kNmTAxNqN/7gr82lnzPFtEFJt6BK4iprwMyLPbwekJ1lxHs
YQKhlEHKcbC4n1gGJ/HUsgHXQB2cJJ50IksQtMJx6h6GFcsiKv7OlwUavPG8dz0i
+tlcb+2XPbB+BPvWEUwaQyS4Oy58eBmuoOVy1f5uOPv2XNC63ydh6po+b3i+Zdjp
`protect END_PROTECTED
