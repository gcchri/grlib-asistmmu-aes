`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VbvYIJvufv4EZomhZw+niNShvrqy9iPGkS8mwPmfXMpCX6g/ApuPeOSFc38NfBAO
Z0MJ47pXTpfUgniSicJvrf0CgRL3XJw94HbNGdKw3p4JgjoyZlgcn3Mbwby9mKFD
Ubw1KzKY4hHKywGyz/lFlIVViiokxF3bEFX6Z2eHXgXh9OifMHZz0Dc8t5SThqBG
uQznUMgZ1tnp8vPJHnbMKqpskufU1gb1IdJHIsc7EJKWNyeocthsUHb1K4dtQJ+O
jNdnVyGeZb5WltF4pgeH73iqkT8AUKjaX3CyEYUZIAjMxRYPq3lGxdL/rvX03d7n
fwp5ukVLK3wkQ4/inYNB18V55UWN55tz0HiP1eKXubEeBiSFOVsT8hBiQ7AZitVV
Xt05m54xtqNvV5nfuNjbFhp3s7IIy7uh2sO5VsBPsm2AjCYf39KRU8DeaoiDQ0Y4
7WKGtAaGRxkcPlFBnRChNbMVC1vb7/uc1/dwHskIZ5oza9ltp1pVOVnY+3bHfhxm
2g3rDiyzj+AZWLNXwuGOt6Ao4KPs2gTSsiHb/I+2lqk9jpDhtJ/y59nkfBCS99Em
okCldGMKkrMtnANJsdd+c4oVGAVJmSyV0NrB/qh2HdGmGzAUIArl63RPYi148fqC
FHCSYwszSb5y3gyvNCH98WCggkU+e+S6q38R2sZ/7inCghU/oA+1jKvqcEYfuM1o
FDpLFflX+4kgM8tjU3UAWHUTzvFOmjahqgtTQGab6IynhsMGBCarkQe8fX0HbpLD
tUh68jmz3Sm8XUO+avRgFY7jYiR6cKRAGD6PJuOGclz2Gxcdtl9Y6EhNdwd+iHFK
1IHdnvH1AEJd5W5CwyvqUZ39RBHnmgMk3R7FBEB934KELwYxeRrGWQu1M0o6VctJ
MmTJcr4uEGjs5LfBPTeSZqF+R0FWP7BTecSW7hvo/fN25Cp8gOBmSHmOMLpzsLA/
pK2KxOStg1p5nAjd+2RlX0AAIl2NsAeNtGusFERuPIQu8vVhR3OALoKFoxtfaEFG
2J6JOEp95Whq0RF+DV/GFdGdXrc8Pir5QL2pAxypNNCOoPLBWYkBzb13nujhKZw0
ShaS/0crWh5Z2ML//2ZPerSgFSo5fnw04Gq+oFqIHfYeCzXVeyP7Qlmyxl9alKxD
kJhHUkMwhPGw5ha0pKhyK4Zu2Fw1uXDqZAhc7adu4oiQKzS4/Awm+YwnmCVguNK1
VwuSJUj7c5Dafl2cYAH0gVKxVfcfTjdEKJt3W2zNYUdYYoNwCRbP4AT0RMDHlOuF
e0zhmeCsafRcRH+kF5UZM7V6580lrqamMlLmPHP/2BFGZJabRoOV1gH0KHLe9py2
+CUwRdHVJSU2RGhXhtA+DWU5m1xkH6XTH3dw5kipVzaDeP+Lm4Z+8lcFlVtqp5e3
ybiogpCwz37jDN9MY8PeNzSN3Mjf9p2O6WKiduaCOAxx2+MoEDmNLVYtrSOGeWMr
Md3KkS2gGq3QrTXOYzGLnkT6/UNM/mm2i6F2wguCMZifVcVLyIK0GKcOPd9fhPS1
bt0+l2fuKDo1OwkVyq/czyz8ipYdWUdlWtVKZJKuw93/80+4EKz91vfR+8SPCCZ9
mauJA3+I8xHCyqXPhXD2+fGPfTdPc84h+HQUJ9bc90UoNvHLNbB0XXWkQezMeuDv
8USnB+/0M+OgO5xH5WiDIfnGUgKoWoCJDcATD7khtzlSstcIdacQ13g0478XgNPb
V77DRQOVcsA64qpVwuImPF6ooovLUg63Z7/pSLKFUAeFguWsqtPcHLGvn0F8TXsW
291Q0WTILe+MStB4LNDZGXeKSruqg4JqHVv4Hb/0KopDAnqqYStb0yjP99CKwiTr
k/vDVsaGg/bcy5EF7S2CX3h6gXoGyMejKd+nE4bqCR3MTeI9ZklGl+pBpY4bRP1T
vfuDcMbRfkHWRfEgVw3c3eo8vTCSDcXrh5sBELCfpcdlAY3gdZWJnRZwCFaXUOC+
E5Tob/C6MOfL8C2JnpNitePPzG5JLjQt9W7569EpTFcBzY1k15f8yZKXSJVRQhng
KrNYyfPBGTkmxhVDpknHclHHJcCXZDi98hwOyXTWQj9d4lyqGgB6SvJYbx3F5gEB
/GMWrChxqxy2uomWMtUQrVFhqkLH6sze1JYV28htoOy43UWCg2+i2Xm2Qh4X66UA
waM1H8i8QLldKE11a9KjjFht1pB5o18XxBDlM44pd9IrNNxNrtmCCYgCc2cZQAVS
5Ie6LznFeldgDyz52glLylP0/IRyDXpxvoZCoeHfAJIQt1HFBogeOxJbFxwA3Jx6
Hh1LVffK1rD4vyZaWQaJOwOvWQG+Qk+o6KSRZmNI4A4SRiHOUnNK87ElyyimiopB
dPU+Tu+cv5xKENwSjJJfxnq547C9Zs7xb6+ow52YsIv4v2dsSWvU6o8e5QjVMB6o
LOLlo/y9Hl4bceQMntg6SdE9UozqcsgE21abhmabsE0l1oTXQeH7cPOE6lfM8i54
zfbzApbhdlrWJqHXyICcbVk7QI2UgaR/GvhgjBSN8zPq7wNNwLGclggrbrpV4x2y
iL3SLIPVmPGdTPRWauQ2oGuHSv7+iJ4sRr4xFhucD8uPr4DWsN6qAUzuQmY2pQc4
VcFUXl+Ovz18JYBy7IsmCE+B9gbjnu4B6apl4+0i/1uzCqpqyIupCNl5HDZ2+P1f
tFpE26TPBGbLm486Tk2F8odMNKcLxn2cm9YHODHnaSOJXM2/nYzUPYJD2O2B02rQ
CuHAHvhWomGPGWl/hz1E1OZT6bjFio0fEjt0t85F89/hLFFhx5Ov8zJZVOt4VKWk
nYcOzGTsspFDuUf9jchqcKiOGU/7P42Af2/0Bt+5/z8tRINLci3xSPBH97AXA7Vr
EIKd2P9kbcIDBl1LHKSG+/91JkyF+hOoNzpWweKR/H/7WfKICz6q0aYWuYF/vYWc
eKikfp86CwXcy/xgo4RFNtU41mC6vY8O+y7aXUs9uT3tXUCqCVcu0PdDlVMac93A
IWX7wDY0s7L05erXqYBf6byDjadNWN6zc2Z6IcozzuevdVd6V0irhspzraVMv4qn
PVwut6Ffqz707AN5LtmEM3k/eRUJCLsNt/zFrdIsxKxvdU+sJQJtiXCenpWGSFFZ
BwzR+dVDmPBmbNn+7knWO5B3BgskrnhI0V2sB7JV36AdN9tXGYxKcDNKLHDEjFxh
YDofI+pB9ENOEF0Y0sy1qbzJZ89K+x5G/3q+jflcV5w0GQQ4cE+5qsdKrXfS/yTH
evkJAM2XhWZCatemjCpi1m+o2bcztRPnyXeXNcbSjjYPhDKOVl0f1xG1W0A3Qof6
VaUDLX9V7HydLda3mE5xTbbLOj5TiNqH/0CRF/ilD5TJUL4in3/vUfkbQNWIOesS
nMqnVF1I2v0Gq8lEi98Hl8mXG2WitUo/Vi/Zm3ehzye2QSpljkiQEkgSqvyeVXou
RnKZiK3oL6gkoFDL1SJrmIaFD0MmpSzcGpMPztWO7yeM5piWI92BjmKan2tZqpGM
VraH5OqpWG/73iSKobo8+dwiX9h9oA+g13D3gGtrsvdVuGmmHHA6wvNXR7IgXEMC
fCjv0qDzuAfdB9J49Ek8Px7m7Wv6zPyB1XSMcZneAvZ4b77SUpDat55DCZsBsvVQ
lzED+WaXiHPyV9UA7T/pwSfYiO3iui1Wmk9M98mZIn4gEd1sQFu7D3xAt+RV+sPb
5+Ghrjl2GP3tf0M+LfbHLDhSFsgeYi9WnPLVpcygLjXjDZiTxdL/aJo17ZyGss9i
rUwSne5WYhWjf8JWUYJM9112Kdag+q/bLKKnP1tROOR5OAScN5HnMkdunmITxvRw
jGewaHZ1/cQ9Tlw2aXTAy+A0Ie/bjeLSm6dlo2qCFBpPGDBlZbZGPw4uKEA4A50C
Qf27faqimnsWYxbpdRrWrlAiDWw4DpgXGh+T5fftRfvegbK5hZn5LZToXP2TQKOb
TMVTCSPBlsmc8mAioZs2Rh3EOSDsZiqyQ44yoOJVBYkQ2ZNN2QBkpTX6AkQRix0t
Z9GAkD8D8ghVRFK42vidufVI05GPXgV/EYQWksLCgOfqjBywVbS+8n3b82Fzo0nc
oBgNtcPcf8vCIOPXyAFaDQ==
`protect END_PROTECTED
