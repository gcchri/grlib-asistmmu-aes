`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v+w79UXUX4hwlPiXuzqYk3OP0AI1EI8SCA8I1Xe8cuW77JyrLl9xrHFrOmZLCfuC
QdplFd2Y79Fy9MSUbtpv6Lj1PFTwQyIVb0TeYmB0xqJ+KbQyfgzNzlkuQhfgUQD3
zYxWqsyYcgZkQzBMWZNeD+fopdgdnS767AHG87in/3fx9Xs/Bc6O/g6iQ/Wclw5E
DRoFhKqLNju0mFHFc+89DbEm03Z9P1NaabjXNRHlb5bnCsPTbElFpsn7pEBtnQJj
oZONxdOJDvUkke/l8V6IYfMa+lim6vbVyeRcEGJRL9+/yi8nMoZPnG0bNYO22J6g
BY9J1I2HBU0KRv1WaLeU1Yw8Nj73Q2a8bgtzF7qnqUValpJPVV7gijC13E6zxXhm
u5/35+Hw4BsZYbC4pRJMKjobN8vJcClSAdl/a2R22goY7OdCEWyzeyhnv0qvTpSv
3gucJNrne+huk2K58ldWuzDWy6pTHxsJEPlfQJ/FZJd/l0kP/RpJZsOARFNvTA75
Y5+dwzZuxCmnkzgJ73DDcx2Uh21TvbfrOZ2YT+dRFHMiDwl0+ut6BcJ2O6ETjTRA
4mWQb5Cpi68gDfWlahasEGz7RJrAavdwDybUB82MZQEh7i12lK6RpS8QBX1BBwzY
sBMzsS+9hQUh8U7/wQTnd7p5Ygne8zNU3110W0k6JY5mdC2LJWZpDTlVVbC9O3b2
D5Q0F/SNNr/YyDnKA6G33eHvye3uVC3lSW95kEM84qq3XAYyIZOegMmwYecsL0Vc
0kjgwZtalj0aXJLbYAm4CAbQhghF6mM9aMtLbMRFBXuadXpzemdXNAYawV1i19Xk
yFedJyBVybtI6oS8HrmEs+sGA9OSvo0erHX/vogSTRWgWRe3ZQKYhYZY8ROV/M6X
5TpQ/cj2vE3/Cq2q461ZkVLiD//8whx5FNP3cIMGeaNanr5L9ZaxPGIDKBCIGHq8
dU7eUke53YoD209Ri7qm3WwNUbnEupQG7CltrOvvdDgSprv86ZnUXP6/5eLLhVwI
vz16r240GtoLqlKMLIvia8yuHn5qO/8scgq400kxDb9Eu55Tv8cGp/d/jg+DmRkX
huABg08bRXRtObiUY4yFIoNGxw35Zl4xXv7Sa0/v8MgZ1JEd36Gr/kXrUG3LrP3Y
SGRDQqxGHUw+YX66GgmHi2FC723sjk7yBn6IYX7JwVxoSV1pzrYJmhKo2vv/vTR9
2CbKamr2VdQCyQsepKFsZZCVIrld4V340He3AIEK4Mx3/NN3NqUX+2tpxJA3rnAm
`protect END_PROTECTED
