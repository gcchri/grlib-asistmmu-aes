`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QGKO7o+sEkeYXJevAPYWZ3ELkbWrdAz6yALOTaZ5PIF2ykrlqI+EXkhbdEMI2rPX
We6aAHHQHnKccEqPR9sbdcyTkHZL8LZ4BnIMGEJfwW8uGbm3KTLaWZto88mGFgMg
I7kSVGJd5dctTLhx4js81Tp4K62CBPNz6cMMsMtiNojZXCdld2b91IBuXtSODXzq
1e5skyN5Mvft9fBQfjju8hznUJOw6rrBC4mHII2kGQTixGZnC2EkF4sBZQNVBp1v
zlvru+ZUgvT8qRjR+Z3PPg==
`protect END_PROTECTED
