`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s0Y8sUoUrnOB8jk3QfXf0f+sgoBzd33XQWlLC3AIq0f3OJB9pydCqFwOV1f+vOnO
Dpj2g9xhpkoW/14pYm9Tixf3Wt0Wo6f3gVHzApvNzVjl9X+FUvvOTqZ/mMPjUjWj
3sdMyUb3cLHQ2QCIJI0K/mFPu4BIv+lf+EBE2KYXqu73HI0444iComPyWvQWgJM1
XpMU+3zlWhuQpln2SSSaINohTPNankVzVpYxTDgwAvsznfmU2Fh+ivXGZbao/PIG
jwieeOOBx3DxOhPCD/1C/aKwJdNZ9v5G43wwnnT+QbmWWg40IeAU4ptH8czupnvu
QrEMfvrbirhsx0ndFzVKudM09MM1yRdXvB66L30C/5k7xa5eFpd0A2AtiFEdV/YA
Hvs4AvJl1YqW2kevnX5JKvFaYCQwEg2eQZvfIVxTEvj4EX858kGpaVKhkecv+1YN
TuE+Ui3KtrJIl/JF0zg7X5wXfMfMoZ35M50Ia3HnYUwBvGzjND3RySdNS/jPIZdN
63zQXTqDITXNZhkaX4pur81etANEGYW5Y+2lSMhIMigiMqGdc4+RE5sdsBaofqsX
0fEN/c1bE8C/M8gGSxCPwM3+vgmneHmgY1/bDCx8vRTgLI/My0IyJ8ak6pFlkBdn
XvhAyDZNovHvUkFr9JVCEHEpwXUT5oKAP7Dqjmw6ZzzUYYUPN7K/1IQIAsu4jKsT
vMvn/crPs09A6KN0WqhQcHhgm6XF2DXNKsqNfkRjv0kT+l85lZDCuJVYzBFyYLji
FmEQ7v/fvQAV1H9aYByLD+5COh8MII/GuUD8xWnLNIxE7QS6TaeF9Aa/BaM4U5iR
YTD8KSbJHSo7LSK0VCPKlIapReCyuJMTS5FESz8ct0su4aG3Pp+/REkIvUqY9aV1
Mc6Tw5zooaEgBNBuytvkkzi7OOjn0Q+wO2PAQdpJdg7fYWs7CNUSaOs2CnukO1sy
Mg6Bx/o+432C+q05qDvKPT55J8Vvu11yjTOEbFRQ7iS89ThZI1Mpd9YnkQTzE2Km
/8sXHM6jqWJ72sFFs1bXig+41af7UnHCU88iC103h6SDx6qHdd1dW9rwKBUXoB8T
AwXE4UdBe5/gHNuXZX8G8fDA0jRqCcCeZdY/LMfjsxDctMc0olWfwpwxPZWwXTNR
xVrEPdUZI3OmHVqUjDjPRRgekq858EgIrvtOmjeRRYwwk4okKW+yUD5c7BAr23x7
RTZRdhPtrV5+zt9rTLcdTcmlgdUGA4DlsF1SnHRm22lrDk6EPqmS8JIpK+NQ3Dfu
FR++P8xR1+gm23hFJ4J30zqRudU+HlDANa9TF19EkyH3mJRKujYjyJ/+9VoNJQfI
xCtD3wTqiGEWLO38t7l9Spk434LwvodKmRbqiwZ/eDwziFSguXgsNXepEu3rxqSu
3S3wyWbVBoCmF9lu3ioi/uDqWyvefhsroCC+X6eyYIQRoMoX6Z50IFBF1WNDLfFS
zXgiZq2L9HL2OmZFiDNCgfUSglInRwSUZOwwSX6aMzLvz4v2DJ3HBcSPxurxaMGG
9h21hlR9+PNIQHVWr83eKfeiH077oQery6feZrq4i+//EEdVgfVUJb0G/RW8JIFT
vBZFRV3jLq2+Q6QxW/46/EWHtuk626Ubwke0O/5vYxWybpQsVT8b+bCE9grRKxsp
4j3+0jKX7wr21BujPVgzSfRDG9DBIdstDzrl+Zxn2GFlTFVM9Rv4NiXcdE1NMOwb
HmcBuTNR9NMDxEqu4yAlvVQrgAcTtu6TUdH7C05gAfeAbPAnq99UqNfATH0qNLTr
Ly2wnja1xvuk+/4Zof55pu48R2I25rMZdVIZmS+xZyAmXcQ2yfGPfkViZs+xhYNk
kEvSiygocDe0FeQui6AIMwqa+67agxZPNegTrl4ViDP5nalc65X8/JDg+LdkrKdh
z5X2wjkfUhfk8iV/USF0EAL2SqRpaW6wBgC0T8m7kj5kg7gE01xM7Nn+DxgiL3u3
BkIYo64fEsoB4cPZSHbfLfcvuVloAaF8nKWbPbm7Qv5nfZzQbvbn8OCgOrQ6HVR+
gQtELXTLtvotGyWktyXr6NZgicaJ3uKL24Bpl/CocEC1mAFEwACpLPSRd0CtnZ6m
hQXqfCwA1SMJONrQjKCyL3WCTDVoU0lwdIbmtJko5YQ99p31cx9wPlkjdJcljOFc
ro46wkmSxHF4+O7o5jMUj6e6QwjHyPx+4Z3mkrkE7DcpgCGQocvmtwxy1DGXuTxN
1axgQ3OXDQ6dyg3jzvQ9pZILBPX6OUfrdnxhKZUySyrsrlvooJ/XeAnxL4kHYE5E
UJlwfEOdqG9KR+DWilXZx0b4McxXxkDdwyAX8Vt8X44CVC0qG136dtqCg2Tps4u+
KFpAfhNx9OIZl1dHgs+F4EU5XNNkP2uCLKT/E52Gycpk912C94MuExAPn0O2PofE
RyKIbjNZ6vUNflj+zVwGRZYmwF8iQhtAtKujyscdTwneM4nQDq8AuXEMSnEj5tRq
C6FAIBJU9tqFcTh7eUpyHSYze/tZmKSd914gMmP18evi28bmj3c2RNTF+VxuBA7A
CJAtvUD9YGupzQwIpWnZgSzzyp8+Q3p740+aaBF8o4lwLSCFwD5X1xVepOTv9AwY
uX2/oh+1pijiHdAPYyNxsu5aUvSkRPJgbgt2hoIFydzdOkCHz8W2YBIMwRvOl2KS
b4WPQyqxChnjCPtULi0omnvyJxORAkDmboKjFtsH8j3Rr4jou1efIcxfMD8B7wn6
YnqpjAbIxNyJYqp49Xvg7DGvdSapJM04ofHTf2+/YpHEQaJGx8IJFUNqxMNJt37I
4AqNKeSL8Uu+I10AQ41CIZSeZlWCP087x2CfzEs/gZCtxAFntAKX5oXgIpRdonm8
KOUrLpP/vuahzTheEZO62/et9JNL4Ueqll+oyKMFSx3dsGHWcT0baXEAERnad/fT
9Z6q+6DvwW2hMlNWNnwCpHQ+IF+2MWYIQ0Okqjn2n9vNsoC7V0QY0T9GREtP5vig
qPdPliROGJSyP0rHHHaIQzXZc+Qwi9sBtbegrbW3AWms4kv7hzr//lL6IqlHB1fu
nKKmoUDXgBEqV7laOYiS4ekkDohtmwf9b3wBIBodJKbu1TtZbyY5e2L6fWXEiJfL
xrYGoQkVAXrZL6q3Y9rt8MhHtU5WS3UPZZOL/FVceBzgT1g4q0dXcIWfsrAibGIh
Zz38JOYIZpDpA1cxC9z93wDA+drOrbe8475OT9xMr5RWx+vs1zemktpmOWg4rDda
4bZPTaaTDd5+wOV/IWG1FlFjZ6V2d9tIq8l/XVRUpLBO3+KBTNGMNnpjk2/3Aqto
EjC6mLSsYEE/f3XSCmlEtI6av6syZijxcvn7KosIxWI1MLk7lvBwFMbCk/gb+04u
B30IdxnJZAm9EzaaUXMpDfg2VrbuaDDBimsxWItoZEjxRWedFA9HAb4KnUXVXQ/M
W8lu4IEg4G3EjwY/njk8sQ==
`protect END_PROTECTED
