`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BebU3r7oX1U4CobTKqKragMqvVv67KBXDlPq2isBM7dxkJvOeYs0OPhaNFZx5+p5
XE4Wx9Twr/3kGCM7NDMX+zPSDhtMC9S0SGxhathS58CIMly9QdbGxTLRg5/DiXSs
pY+tQaXZ4EGfVBfu2/hQUGV2EvUqZlM4wJCXdovnBEzApsxHPQXSR9SyTcANM1i5
KXQ870yhTB7CsWgCnbRdi4uB4sQRfZvGWyltkGfH5M7cdTnBdeYsacFo59ec+zgC
chWL1YZF/mjEv25h5hVr4I8iVrch9huXh3OtqJsYkY3n1buKv/YX691iz9Y9bhbB
MoeNXRkjMnbUTAgxrClIyZsiIA3zSD6cWgoiRbD9ON2RQdNfT1+zgFHVaUziGOkZ
rdLLYGJpqU5TXVropzXMlbOD1ZikWNPdlnP/9vip90bW0IhHlMY3HZpo3MJ/P3Wq
K9Ep6mL6T/cRnwuRrajbwghTwKWVazSdQ+dmudmYJRkR9lnVSpewi3V5CzLVVXjg
M6DTvj90zmXYNTx22L+Yfo/jUM2fIDqzpBQEDCsuRfTIp1gpD4ASSrurBoq1fChq
RXejsaITlYtfVi0v+xa9tbrahCSv9JPSA3NwMjPreL00QAn1ZDJxckixlTqI6eeW
Qfn9dlMXm3gbTaSIMuZnfAJj35nz/NX5YF+D3tF1lnXBk7xege50voVNEXybZz/j
s1n0gChT04NPGecXqwCzmqa6GH1/ScPm8INQtLn10wvK6yZAEMD1UK3P4cJV2jdZ
EDcd1HnU60S6HiTAj08mzRNWDUx80Saa1qv01n9Uv+opv+AM3BvgNV/aKgRAyFBT
eHgsmRzR/sjGpUoHdA5PhEPA9WjQ9HtTcA5IQcu/51fUOdpwCOghNgpFWlG5rJnW
OiIg2zLXsYYPm1lOlYJvlSxblUof8pHTc5ZLs04FbRqYweklWsO1zlGC0eov5UsK
/t8tZH7KtW9m4Gq9zWfiQg==
`protect END_PROTECTED
