`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k7AdRA936S3ZxpZeEHFukSCVA9//C/rngEZyCoS4CExPmJrT1yll3xlE2AKdSWC4
DoixRq3O4waqbe77UShH04CbaD0sJ4854mYoUF4sJMm9XlL6lItpgNVJs0vQT0Mv
DsFqvkOPPKg4d05szUqbFgqDzpNm9brI+5wq0uKoPl6MRxywaY5F4ka3zM1SMJrb
ZmnsovvUGf+l6x+CwrjDzskXvaSqqivZRUvCpXaFOVfoBPIsYzsfLXKKe98HEkxI
qJWNfO+54cu5LZRukwTZx5iF+wu/f6uaJTcmQW0y5+ejAGwTNbmwDTEJaziIQryK
SptJ/hM8GaF0to1GbOw5CHixuRR7GL+Hvw+Z091yREozA1sS8s8rDOigrFPq6EP1
opoq7mUdmz/N0lzxK7YHfdljE/kQacmT/TgdjrfWoso=
`protect END_PROTECTED
