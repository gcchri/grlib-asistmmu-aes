`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C/9Ck88ihS3O5tzbJQ/ccE1NwGTTd5pyyV6IOkfim8n87oQ84eV0P2Tgm/aiRVo7
pFnFVDt3BIhqK17QVqhHJ4MgQKzc6OUwbZBfGwGs4k8mkDn/DS3qrmy5L6PX6bMf
bQQmtsepCibSayQmEYmy3XXK2O7OOmkAvsLHNAf+RG00FwHEVB31I87qOFmxjPsU
Y7FDHqA5Eynphnn+SP4YJUeTK469dSBFdRKemrmUzMnTkkuQXyiO8lpIoL6aC3mL
zdsdVffWgwXhzKOgpC3wLg+8DcvciXLPRmZNXbqpY+4H4aX7NqD+PAK6YUIVw0KM
pUx5X4T92bRzNG71b2GbRxQ+qdtx6Ob9RTQfLZ/BnxiZO/bAzIByZcfa25i6U8Sk
Xbj/oZ6fHAKyjMvJcAoKkiY7/CGr+3+5QdCFH8XzV0lW64O7RgY35+YB5Qio1Xas
zskI/ar1o5t4G8uEASGQAyqVdgVsLelEwKTSdumlA8g8DRTmNOFcaOIarzI7obYa
FlGHangn2RcftCSepN3Y1gG1g19IFslJSpLl1tK8UwQoyjaW2QvMs9GkNdGR2VE9
euxb++Lk1W5j6mfPzhKiWkRo6NRQEV9Iwp02DmxQvVbtdU9MJ2tynnqCsbOeBjIU
g64dTKdlm24tKCYZmRJM4cXG1R0DxPrqPJPO7fD+QwyKZvruEhldhYFRkQZrwmPd
WDAZheaJBTW00ynv1+3oiygY+XVwZwptf5HbMBduRJHw955Xh5RCosaKM0zkFPHA
71D4UkHvWYm45c+s7Sz5nQ==
`protect END_PROTECTED
