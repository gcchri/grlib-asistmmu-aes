`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bzkjXNRZMeEyXrVJ0Al+MRXpFb1Y65yjnxe4EU/mCmqqOK5uxJ2mVDWT1LiK+9x/
V2EQMvUlTmklKWHzrdGTkjydVWUEj795voI8WBCQ/CtVgDs/ohj4yiV77qtGBUYR
eIcPdCeAfpQAbTPJ0PT5dQ0apqfZ3jbeNLogQg6YXPoUbzsOLw4jTIn4QYhnPszF
qrvZ5syAQeDLTYU4tvvha9OrdOh5JuMUBaVG89X7xOzMxkbLNCx4KSEIZ+qc9cWW
H9dRex6N8EE+1Th/mX3eVR84VPSt4aWXSiHt563MgCisDSyAi8cE67hbEslGGc4m
sorDjb4iv8ZPx27kKqMeFpGvxe7zt2kYjP6TCl2H29KJTtNrpLo6jD+3+eVKWzMh
CwhcGHXu6XnAC5vfqA3EVDVqpirP/EP9Xd3DF3rvMEmw+PXhvSzSztvMSnAJ7MjT
OpqoL9rnNreI5qiGCrdT7GFTKvzIZK1Yr+ln9f2dbxkNsNTrD4IDwD0gAbTMH6AJ
Iv16RwEYEY6Or16eSnuasQ==
`protect END_PROTECTED
