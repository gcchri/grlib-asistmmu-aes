`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SChzU9d+8P3B8EwD3i2gohz0SH+eWWPHkbR9mVJi4yJYJjbcgZULECUdHODjXNn7
wBnm+rh8X1SC/EE1cI5dF6DBWaJkE2ShlIXHIoN0g3fqko3i9hBgO9drKPK/Z6zR
tvgYqRs55cPkz63mzN9/imv9C1YKpE72+s6RBfJFGvUK2SP874TWgVUXDV1yoPx9
/SsIYkWlN4oIP6fjF+VRLcwJxcj7Rihsysce6iW3yAjC68rDsYVlDGOdhArY6vXE
lIssXsI217gDhOKrqqYMIQ==
`protect END_PROTECTED
