`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ucs5u2upCC1vcj/ARBVCtTFQITIT8lE7Ejrv/msd4jDMssdTVthmIRFEDDVUorF2
pg2AbZ7mkOg15s1U5Nl9DOu7ycj+IFJBa59pZiwCKljTI/XvEaM5eadbeIvvC4m8
8sQNqz9AEd1MJU2mZVljKJxQfZEG52ZFbZh+yBkQhRbsQVfmnjAsFYC7KlvxKxlH
NIQ8Qdj0OHNoLHXoLE7Y2jQ3E6KfGQgGGGaH8z6t12XMOllnA+XEIX5RXPQL3/5A
zvS3sP9VLRorRlL6722quKZs3Wfu75acvDtfc9Mzyvjnnn+Xvi+YnaJkoBp8j+rr
dLoL8ALIruHtLafXSVFPMR8juxS5Lfh/BQDj6JLsioor5/xVl3Ny7TFNwb2W6Pwu
IgWw502WL/bmWDMsFp9TnEAVaBwXy1IK+tpioVMLp4lgm2idJdrPmyJmgn/SuZOh
9Kj+C2TfJyqeXkJ6BPgJ8ERGPczBuW9nzyPdO2f9Hy0=
`protect END_PROTECTED
