`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qQemFwU6MobqwWV7hLJ9stPPSA72pqS+tedmyECmXzeJ/oPS6MQiN+/rubcAX1R+
cKbSQ9bGSyTzUT/prWwqnf3YdFYUKl2Mn2ema/se2W4h+Hnac+KlgHk+jpcwe/zx
dZzgifjK7TNrjb8apKPlgquW1MKWqJuv7Qy42USEMHtd5yohUASxBreTor1eBNxV
PtRr74vvhA1Mu8TvveTav1zvli2vq6SaAyAQJmyGOrlBvHYtbCb9iIEcuwNAMNos
gg2Do13+GfmgYocSTdrVUl9vdKmsyIW9Unns/CuUhtqos6EP/pjsiBzEJgwoGoHM
GWospne8Qgih5OgbuCzqXkol4wcO9jHhjXlzzWmakBs0VEq0DPKRStDOJwcDuuH9
lin8lB8W5k5VEhPc9/ykcc+D6VAFljYhs1WAupqPgJI8oAL0VNVX4vn69jI7MQ0W
JR6gTT77nemSBfzBxykF1dzkt0RcGWG2l1LXcftK/Y85KIt3aOaU4Vrdr/N2Bdu0
2zZVhQaldhQyxsv1zGcKOsLGD6F4r1s8Eum+flJPTBl+bV+ru+yR8BAOVryuabDd
G+Q5RVQHzKB1OPkYyabG74QgPk9I4EB6zPBDXLYSqJekmQin39VO0GLjPBNK85sm
hpGFdbD9NKwJ8StGLZZIkwxpW0R7oYuuAZK+v76r29DNsB+aPVUHY1jBCWeQMf1h
mKnIvddIQK7fN5Bu2Z7ypuCLxcLbvVUT08mCROpiysWJWLlS5FUVl8HAa+f1pzgR
cRbSW3hmAnNPRbCTNbbbI4+PlcsT+musBs1eLfYkWPJnWR3jhVwddFhuIiHkYITU
NiWx1mzGsRzFxpDd0Jwyen0BHHc8wT23PfRqqROvMkB5RVxFaWAdp3z+jLQ4GdsB
1dgXvIQiedGAp0yLQeDlrPgxG0xE+8S7RkQAdCHUb+8ZxOkYkCkGagpddZDRikme
`protect END_PROTECTED
