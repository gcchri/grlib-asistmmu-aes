`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ROJjjHemG7TQV0WYYIICPQxFxf7MKfPeZI5L4WEAX9TKHqGSGvFqlkfTNeUMLcuG
NnX0V/Vug00X6I+/eSVGLahdUVwt5kHF5bQ1b1g4T7+o62ihZAmGpAUE5Ud+58aG
Vyg4CUyeVbEHrLMTjqTzVHtyJwlb8hDXiW3fY+Q4Di0cxP7C9dELRoprWzzWSN+a
Tx7OmO0YSbeflR5XD4MW3Hz8Ymx6hrJYEALItI8VSVPS+zQpnLAunm2jOvS4LVYP
j1CXwBUvlP1qidk7aNWfmjLTDtIj4pCJHKbt+B4XsruCmk5nnY7on1fBip0jPt/Z
5z8yD+t0cgbrKnIIcz9K+WXzIlFIC91jPqlQkjz0Vtt1AE7DD9x+Cr0T7vOZmSN4
`protect END_PROTECTED
