`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n7cwKQRcXirkr4D2JyCkILWeGXMWfYsjdgdlScOaKeN/b1q3u5kDDYVO7yrEXbQX
1DtYvOf/oYr62qxcuWMnUT1lnIn2GSUmU03JUgPwrk4vOFGnERJPdy9s9GMzazD2
Es6ZZ7VzB7rbHNhOZXJcltBtC0tPOqq1Jxyb+xMTSHO4XCVTneXXsxuJ4er9MyfO
PG0jmNA8lmSrDKQTsvJvyEtYm7o7yaqUkiboGXhSKun0XqS71WrS/BHQ3v5o1U9U
rglTMVuhRGjl4q/t5akfPaLotR46eq8LoiF7g6HuFDmdQERtNLQd0th9oqz7ay9g
Hy2M/yrbOnyywiLxd/3Msy848W+kQmzB8cdyCeS4EemoYlJGIc4TNS2rLKPYvNiY
6JVlgoiJxnmNRH1nW3k7JF+VGHS5SCxt886r0xdX6mGQGFL+lNVOGoUQJRhmxQiy
gl6bOqIGS0CrTTrpIVD6P7GzaxUDtdqLDu18d1/tDRsbQkzpfGyouPR08svUvgYt
ABWkru0F5NtVGtCl5crU+NN+MDs8b6ukktnmpGJf8FDRJup1QFKxcyJfXbm5sXnx
qhNHfLYi0zlqWLwtcJtCSxt05oC1QyZzwT5Osz2402HxeYPTligqPWXkkJ+z1y9w
/Q8UODhupeGc5OKxEDAfagps7S3qgDhhfq0rMMn9xcnEtVn6gdrXFTfff9psRnMg
jkDFDUIz+DWw7Ha7nRpvzd5KASnDiUq51cQtthWVYgqEA81f/p6vwr6sQyZzX5R8
uRnYiibvo0UFTIwABhQPOJoYSGchfGtial89yA2K3H4GxrLzzu370Bio49cXY/rV
/1+48UOZzSSJy9+MDlAlBrGTrGXwtpZyH9iSm7fm/glSYchA89AbZM5hxDyzG05F
NoBbYbu9H1b2jFwGQWqxiY3BmpU/PnfXzg0n1DqoR8x9uDUpKnTWsqBgz5OqE7bP
0owZd0S2D0vyv9GwZIbUHugP5AvuiH0K8r3d/kAcsZgx01RJz8DR7/kca6pTZ1Vd
gCHaAzkp/Z3LYXRKVNisv4Qgwcmf+UC+4SHL2RKU+tzc7mICKAdaa0tuzeHdeRfz
9FQfk9e90mQzvFhgF94zN9RnkRoPm8+e9IpQmclGrjqCuEDviY5syT/I1h3KhxPJ
/iFFYX5NrUU2fN6kJ1FKVpWly6iZu8QNeaJKhB7q8faudYTTfjUdnIzuRD+hBBRz
07yiSTgAWZUbFgBQXEZbx6oDT/Tj17TAOrxEMQdoYuDPoir2jPPNcthrSBpCs/CA
e7aHiVXHoiMgk1Gt62Mw4wKCvs5CMDMsBRU1NuId/olKcUu9P2cZS5ZKw7B49GFQ
idY9hWD4HXT4IVFlCge30KWbAZRPxOgxhw2eIkirAMqKFpUqP3RBtOTTnC+PA/Of
f11NF7FX0EZKOQQDiSsCq0/vIIAdJlAJ3isaRy03crROz3cfyA3T3UaDBIqR7SQ7
FCA1Lp8pyb3ZZgLJJiZIWVsa/BzOrGPN/YMQsZW7nVgbzjfoprop9PZdR9UICFAh
9KPLEwUBN3NaKBQHmesmU5XLy+/q71e7+Yf44p8GCh+MJ7EtFZwW0fsQvA1YQPVF
4btik8/9v7aSHc3P8HEuuH3GxitVhxhMscV/4dtZesDCf5P7FdA3SjktAH7rBeRe
MsCjmde44AMSf3sOAS/aNWbwHCTgHq45u5OTLKEW6eaLXiM8neDdFqLHyiesaXon
5mQH+06NX7aferUGOmyZzstcgyctmlJrbaZptKAw2itsQvmZzOVU56T0vZ39BpjV
gWMOeVXsBBpiRb0NDR9P0EqRnM/fZO5fcLjHOxsRu5vSz5liJjppEofmEPNjk62r
jOjjUuJaqi53On3wYnfFPbvYfxA6rhWTRF4cQ/tsQx/DlVPKjr/PDIiHq7WVy5pS
oNQ6JFleh52pISYu9M4wRrm3XF851HMMW2YhjB4oDktnohYPo1jN8Di0aibRaGEQ
afn+f07vgsDaQdNdw0Bw+o9yfbLzbyUWaTdY+C6c7sXcfb9+8KuuEjZEWybH7YB3
pT6Tkdp1lCqdG+rYMh+7R9AAnMkV2ifL201nFg9JP97RWhuDo36L6Sym+nbKqqq2
FYFX+SiMguXEhV9g2JODLom2kVyYzv04lafjja7q8Lq2ro17/hwXM7Q7cHl8cozR
CAN6z755DyEJaF4F8mcR0wNcOct1wvqH/OoUfNVZ6OlXUb4Yatj+/ULpCyMCj8iO
ZnErPSOlgDaSUhNpEMUZqB2oXfdgSVGppadujFSKnb6Enbou4wXoli2glvyp9AGw
KyU7hc3X/DXw5SalVH11K8Pb7FCYXnQqSXjV9KLOUvbAzFdkQIX7sgkoytMC4qNd
uwDNsAQDaD3+nhx7PP7zssm6bwIiZ4Bp4mp7mHZYthHclWfQJkC9eby9PaFCI+7L
kTPAOYCa6RyS0/93sYSGFDyGanGYjK3EC9MnFMz0VEBHeQxArTxFinu0q39WvnW9
znFaebMnAnA7JRh34qMNabsWnhSbrb/wKf1RGRi8GZPH8YtMWr8jHP2l1o1a+goK
3pKb60aZB43rIhWl6o9QNPrUxRgvAJK8dI3Jb6eBxDjTcD1qL0bBXos56cbJPnU7
4KxDbfha0RQPqMi/ntpxah9dsc4Tm7rEquCRgw4j4UP7333h7IByqoF9KavtWlc2
dFItCOkQfZkjZ+Z7TerGdeez+1IRPfXv7u+Fw24CTN+9KLWl1rXZK4YTXh/rOIVm
fnAc9SqU/3iIengpxUwell3VvN/GDGQoXir2JA4+p/LWRZVGOPdJkuLXoLEKUKDQ
0+QNezcozUziL+mQc8vP5YZArvdI/Fffk0MkBYMGJA3l7K0ldJtZY0xC0zTQTxlm
gY9YY8OKdpTKIDL3ym+gYcm0sjfSlnUNzZUypEl/kfd62W+I5bPdYpiYrpm0wLKK
xoRvWdLb47RdkYgu5MF9SqwDOFlZYL2oKeOafp0XAqdTasoVieA2ERBMKJbCu8Fw
WnvA7XKJpz827znXKXR+LQVP3SY3ofO+30BJUwCxfQu2dt9jZxLPugO0UWqSJaJF
LO0oNdcU7a650ircalmqxzw8OAt0+SlLBwD6E+DOc15lfAYekDYT2c5ZnsPffRiZ
4p8ZCVkt9v1nQ63DbuCs2BwGw0xetaupk+nTczzVMKS1CglflpGmFc90vQog6qyR
UEtnvTCu13QEDJ3BP3n+2GFqdWqlJR4TdwbzbJl5rMjA3r0bFjr9XInzRCd/+HrA
FQ5J1U1NwbgIv4+tEB8LAijUx84CJQUBMySLg8C+3tOM0+Y2ltWJ0xCJI8BS6ybj
r8Pfo0RLu1A6EGQHqWWJVADHhs210v5EluxigxnOkawnOKQPq9tsa/FZwsYCZv5E
xSiWGLbKvnXlpb2p5ZRXskuzDUJOQ0MQpCW3NNep2JrV/u3a87eaAv1eKfQ29T5C
3JWIHrxzP7IOgYv/jZFu/7FGgqiIkXTijjVqGUygAJpbfEPcUpyVZeSHxJP+u2GN
E8V6uBrJ994zqRhZnZO7UXECV2t7RjAQjmD5hOpwsfZhinIw0pwVYVr7WBxlprF+
gC/oPMlKWkmknK4Qdq9TPLeCegEXsygySFhZUwK6mMr7PYf/f5pzG+Q9ecRDSPyB
zhbAQRS90ADsXCZXxjoDz78SHy4VN8hqnzdbe5zRbWmEFLyVGVIlHE0imvl6EgVP
eW60lzGbRYa6avWpw3kk4twZ+p6qKi3xe/ETUTf21z1QH2Eb9hTuQUScfMceVoRI
EyFbNX9Z3jCG+oqhNduDFH1ibT4qQshyY2kCu3UuwDy3YaH0R7RQ3K9T3fE7312U
Jz4cnOdvUi5xgSpjH5p+QTqR3f9U73eetWKaBAr1U1tkUNsG973RKht5zlsO325s
VgHSVUz6E45/AN8dHn1xdzoRr/ZDYksuWQ3G+MJlzSM8pTn4AYqM4Yanhyv4zOme
Oh3bCI1JVx5T84XExiCzyuatE3Y0J290FxO5ksDgE7cFpmJdUzWSIF6OjHjQiGQN
2L7sjNz+G886JTIKAzwn3GOD73IlmquzdpsRHZQhQto8Mf7DzkkGvfVX+uFVwZIH
qI+1EgCOUlkwPJ/xlnxiIVnhQVli9R05LRE/Dei3HogvYRhyQ1LuhDbswkssKSnY
JLOzvzsL4bWyx3JbhEAfVvDGlXOTZ08kfm9bfa9JTzQl34Dmq02mE5C6qhyCwaHj
2/0FSkkbtPlkkG2tibnMv0hDDZHjpd+kGlA7G3c0LMGbscRLp7UJJMMaGyXNBdbv
h7AyiI1DP9fN+oVUNps3jRFXvM7DSVXLq/b97htf7YiXsjowWLzy0nsY6afySPZ1
YQCEY2ADoCAXOhuqnu43L3vv0Ye4NXvhWXQl6xJjCasVlOx5CFHg3Wih1krIlK8f
DmEKkSPAc4bdUSR/eUmH730vamY9dItmIWG7JlZ33MMi85bo8Bg7tdHqGar2/D6Q
mAFVRA9eUX876O8vlUxVdxH2WoJs63kM1uoh32lHA862zmoXXUWm1ugu0zib7tPI
QBQKjr+CLxf8pUylXJ7CKWSfx+0yyzUwDqKbLDi+JTMO0lw1tTt3kYPXQ8LmhnLV
cI19V6XVWWZ84xXd2/8MHgBx/PR9sR0woobcLRNgDEAXURTzpzdOGLZp0kMGTCPk
SMuYMRm4CU6dizQkPrtAUt1FXWQlj+J3CKiqaq+8+Kgiyt0wEJjEFIhiaBylzqZ2
hByCmXkjT/7vVXslZRk0yo/1Q3bfXLcfoF2j6mUkl7vcsRTRskaWdy/r5ha+MzvP
+cJ1Q7+Nv4x4/Lp7DbIqVY15vepOYWTJCyA7xW/kcoq0fEEnGAmJzDTaGvz1xTkL
9GYqXq4C05vJm0ayTxd95Qg+MFHtmcaAkzKcekSafwAgpcTbv8fLwcbFj1zUoKLt
qX4+RFhJoM/c5FW2FBHZvyDK4q5MHSoASUe3Sp7cTNHsatgcSGQ8RNKeV8gNLy8x
WuMgWj5D0+Z3F5O5uXA3cdR+Tq5qZQjyD/DzTP+7KQEeberYlTvDZyWfDqLvgIZh
AxPP/V4Nji4fZ8dEJOWdCKoi+Ncu4eNEA88G0Xo517KO/HmOGkq/RqEsB69TPNK8
iRsRjIytTHEza16iR22P/EKw+0zYNv+7LWUa0YFQxllKNy9sgaoMNjUOIMkqe+5a
t8SIBnuihBya3ABILojvy8VQsX0kW7Ktv8EIM/NeEvFAgdoOQ506PJU8gooiEs2c
tNL69tkbyloycSr9zpsxkS5O0vhpBpcjmhZ+bI2caCiq3G/mLrUp7IYlioLd3JMA
yBNDX9FKvTzvxHEaP7Q1Q/hDLFQppZaek/hhQWxyanUXkwgAtp30DDN+R9RE3GyQ
ubyJo8gZ2I9tp+/Jsjv/GAUV2OGfdVRJnFWdSNfSZGhcggu4XVIaPHdG14h4dz1d
3HQtt0C6ZiTE7OrJvMBK0ZFX8ATiNgk76KaE81FW4fZQMV/fejzaSbhAsi6LPo6F
mu6/EGb6FcCIQGE3dnm8+i8NDMppt8mvwW9R4NPyeXfbguoVKrCTmG/Co8NBNTlw
OcRiyXQCtX87SpD4HNwOLw6qoHwRKZX9rA5n7p6r0pU8X5I/xegLrH9ihXUaaeJ3
5B6CfbIPEVKvC21gVB932zAhaL2vE36CzEod2r/THozv5tVE4yHqVgWah4ceX8g+
cz2yyn+o4yS+B2U2s1hpzdgprRN2e7Vshte3siQK40/gckqr6vx740k5bIJzhIbl
R6N/eJXUOZYc6uDbwuC3km4DpttYTM9W9t9IBAeC1h7zlI8ET2FYbL/Dfo8yA7tR
0jVBMbaz+yEmSQSDO3NkqV/SFfz/6QSTe7eeYjCO6v46Oh4Z6niAAXK880WqXW4W
cTRYBu0uIqaAwS7kNDrsv1Lh3b9zOgPzxOG9RkoBnKn5BaFhexoihZzeNSR3XnJD
yu6XKxJEXjGU84e/QU4INMzOgd1pYxJtJ5aVBZ71qO8V8jABoMlqgwrqfv/OAyn3
gW3O9CfpO9pTBZk9Nwy0QyZQ5GJcV68PkrbTWvhbF5SKoWBocPo5GLUsF9m1J3ks
nQAv2anvrcbxJtnqyfPWhuzbd7tnfZMJhkmOgEkhxRw6tlWzfxhZ9wHjyfHjjS1d
q10tZcuLAillTZWSZEff3OO2GDiL2IILBRmjlzOGdaz7YKLDsOiz1L42DN/8ufdx
hVXsi0mcdGLg6ll8alnCyoz0CaAZLBjXu8JS0ogxs35t+efEZkdPuYYBPi6lqdWl
BSLYzdI9nPpH0Jo92rljPQ==
`protect END_PROTECTED
