`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3eSOlYB1fa3xylz9KjNIAgxhYm8R6WZqg1lx58fM7A2VPGVKedl/hiBHBMJa86z2
lO0dMIgUIY84dBEUJFRVxtpOMLPzIQ9hBGwgEjGUJgN0oYMSKMIvsQoKyTx8XlEB
i0RWAbdyUysBZmpF5UleyA8ryr9zRqbPGuzuqeN5m+hARqegaYKDwjJsgQ+gjaRj
utWFyNsUXksnrNahlnvK5BF3g6CXhINgaSeGSMtbHoQrqfP0H9/Gk9ibA6sT1hXU
dW2kmoAeoIqDQm0x0s+lizUCp/J+XWzhIlYuSYII9EoDXkmy4a7exiiP3sfwQZMy
wW3sIfBefBN31fR3ClegIFj44URnmVkISKsbNZbfGRrxhgP6g6KbldNJUEggfVRi
eRswQr8DLXWN7ItqqJkgoBRIJTgi1SbiGjFwXGbt9CD07nq64Dg6voZj+RW6p2Hj
+TpERjnuxPGrdC8e8YdKcuMHtWLhSoxpddrgMiPHvKeXqt+T4L35BPjlsqJErmWy
4wDUGlmN/cwNi9ENMf1WYk7i/YLeK+QiakrpbB59tu399To8wDvFkWKzgY2eJJa7
ESC4uJvRTGebSLsAYlAxWjz2SNl4eL7vc/8bhvBV2yGEAy9/VeqKx/HxkUZe9cn9
Q9QwBlLYY29goUPmdMYldA==
`protect END_PROTECTED
