`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Pyn7O+8l7Olqa9jWM3DlFMAy87nJb3hWKCcx1H5imyPqV6p0ozjLNFhcxOiNOHy
alsn9ERB3dyL3jYtgh6yu1yibUj07i+BFv5FUR106GyoNkyJfP+jC2vFdJB9exfB
A6unCSZ2oLbWtCxUB9CAf73ax9TYyYW2BRntoCgWGZwddYAArVqc0kiWTW/XWaGZ
nR5EVgLWtNSBveDgaJ4hhrMB5bUBOpxwmr38H0F2RXc2LQ1oSM1qjQyBM/1Umanw
XEQ3rNaQAQMMToyfTSEfp5phCXnDh/d1apoU5BRiciJwC5v83HqGWlcrfeVVGSYc
2tVfJ8xNmvg9bmVVF6Syt2Knn0QmXaXbWJZDNIn+CIN2zxxoSSYnTri+joRmK8R5
VOo5zCOLNIK3X7Iz4HLh9Dgy7NupUQhVuwNckzIB8ozRjsKRQ92h6GnhdQ+JQlJF
`protect END_PROTECTED
