`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sc0vHDU1RXrxqyvVxWhj0QOD9GRW61rQc8n6MvROkDr5PuiifQm1//yhLaRsAxVu
9DmCJgQAIhGjSFfLy0qjJXo8oAmXfB0WAq6aoZC1U9bXE5B5QDs8LGGcunrThIXt
E+/3c9VJ6B+rG5wmREucDAdOCXAtweZ8aanhxTZT3/kcad/kFpPBM5yVe1IYhnuJ
r6a1zTaarwcAyY9UugNLVU3P0UIgrg2uzh5zys0gbYUQDY1fh2VvZueKF9oV0EZg
x6aZTu021TfuJtgRGHK7MfvVTDRkZyS3JRROhv/9IrC1hMMoYXLkcjy8WYgtctTc
0NpeXR6UtF0f3JrChFxnxU67Ao+lZ3pK4TvtE5cF6FvL7KAgBxmmeh4RQ0B5dQFV
RRWvGgdFmrgzvvpcd06OlTFyTXL5VhURj8gyjJz/bAlS8wlBd0XaDcglk5QS9yoK
oRklYLPWf7VML4QWCbhbYpzMC/KXRofBtYTFFbiuBf0PAZ5EXv50B7J/DJOz/H+I
YnM+AgQxFc2G4XMZhoM2bUcYkn317M9U+Zf5VeTQvZWwSeMcIJRoNEhBJinL4DfR
nibnqH2q5wP6qxx5EzxW9OKimNQfOi03h64Y4W8ddLzPUydkFe1ab94wrLnhFqiV
PKydkF5n/SsE7srzHLBmnstu3QUOABBby+aZqNUxCbJFahhUrUECeuPteRs7Z448
OgJOfAfDti/gNaaGn6If05yCoSfX03atU4bsQvXtElZYnmZlu4IqfRmb06+OBUcN
oyfoM/rbvt0Fu7FPw7joE8f0O1qeX8Qk2wvQgIAAmpnzeakZWYHmjPvhCPGyQh5N
RvcsB4lBNEQjxz5GQopzkK9hmJLU6h69o9YpIJ7yyWOH9W7AqhcURI2umY/q3bVm
`protect END_PROTECTED
