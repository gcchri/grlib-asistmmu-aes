`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g6p3ZsUK9tPtvoWMzAyWnLgEPhD3iQqoPHr9vpz7qJlm6T3yP+RgwMuTob6LNWy7
P97r5+hUKsDVltN7OGN5ea+WsPO05OgvC/Cn/ma3Jtynni/CEUJ7YjcNBmil6CuA
IMmlecTsmcUGWPc9I1UvZNTvXLRmJJ6vTOR211vDCkhLA9wUT2MQRBBscyMmiZt/
XWXH+wLJYkO0zxmbioeK2OZF0pFN2SqS8RavGl5rxBBJhuheRokLEhBye4WfnS5o
d5W72Dfru630AA2MG7Srq39fvcWjp8fVj4v3E6GhExEITbRxHTlSOVWC3ivRii/G
RXGdqrszBa1mDx/Ha7EDTA2wQtFZTBZg6wGZbz4UkqZ80ooYGCaHyV4wGx1RUFgh
BNIHiwprQLipneldfXzpr+cCrJUjypxcZLGdFXBmtEM4o7ZJNDOKXNpsKE5BqObC
`protect END_PROTECTED
