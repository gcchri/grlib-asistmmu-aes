`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bb3jS1PzvBBu/+9A/auYmDS25M09pQBCSuq/Wx2mQYALlutroGgbin0d7rWzyhE4
TFWPjR588SwrbhFpm3athlIOZl1219xyn+z2KVHz19/r7DU+KdVenW+67ii/9ZOS
HYrzBN/U/1uFpJ8eXEVUaAxtqw6J8vxYjGjuNW162ZQ/FjFNQPPVfX0yWx9s4UQh
bWNrxsEKWpgc3w1kbm58eMja3f5p1KbaBkzZPHT/ksiduyDq4IjQ19R+zWCbXE5P
Vs052LoVRIc87RXa9ffifmlmIiNjd1Prom2+ooOhq0jdFGDFxVU2KJVVXMbnj6W+
9vW8UP23AoLHDZw2XB2ykDjfziqo3SPglqVKJ5YePmmkklrsXkBG3/pjY90j1+H2
whu5L0OXoswFhy4lk2y7b2FWTyAf1pLiPoUNlZnI4FVlqGh4D5I6yeXko2MvKUBW
Pvd/FLp3aKa7axpgdjqgsAXSd120WsbaOZLwMEygf0HscqGBs7rcNJ8YqL9j4VdF
5OrbKdPrl6QjVJmuQCCVOFSoULBbLXhzdyjJfktYuyIwpAjbj24Y0Tba+7RJ04fd
I0ejjQ4ayS5YZCTeMKv33zS0lIeGkGFfQ7lRPR6lcgk=
`protect END_PROTECTED
