`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iusk0LUC/shhpn5sPFgdyVaQepXtXFTmXzMaiuf70fxAH/ligCysvfsSWL0eZosl
mmhaLxUBclnaJWPOChyqp4nIBFLjSCdLAovL47rzWO0rVKVMg6cldvsMRIy4XGBq
DvX/1ii4DXcVhKdW+8H2XdwuErrLrHSUpPBP8qSuuW+cg9gcjkcSbazUqkL6AW0k
S1s1j0dq4xparTNvPaYtOPzb5k+/YtPYFDuuU5q+0+ojYeV8C6eD8O/2HRIgp0E5
aYtyy1eD79l8g4l4ggZ94ayxBNB+urVeW4HuJJG8MtQ9o4ZmM7hQl3CNYemRi93/
aedqCi1bIaB7nlhRVoObMv24D52HdXK9EHWpGJCa7hU=
`protect END_PROTECTED
