`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G2Fi59/kQIE9mB8kgy8nZiq2J/SNdVeQ25Y6191IPyuIzqm6wVhD2Yam0WdF0xbV
/JptzP2pdrwFdh4zCWANM9Y0eX3jxGzKWjVjQaGLylp4HL7WB4KP28qaR3ssi+g7
378rnkjq2AcqyDee09v6yfNAS5xrzMRez5xvFX1rh4ik04iSCUHeQ0b6+eEjnMzK
WTOi64VmF2ruuwpg3yO7VjnzOPUePxoA4AHzyNg6qIN6+HeplydxWhzkjNklCkV5
7o+Qy9Evk+3XCv0MlK1fbCFooRlgRLzYTt1ABqTwmdCKO/zUyMMqoeUcz0SA2HTx
jkNjFseS2UGaBiXWqe29IdTg2dgrEWYNAXVHrgD6acA3scGZkc9kYqau+RSwbukC
G3aSnledrx2hXA4jYQa6xByQwrf1Bx1mnacW95f/yty0+094RZ4pN6ASPqO034Xv
FAeZG52F6wAbAj06ZYQ5oVD9ODYzXMWy+Xc4efn9zczCmFkykz62x9/qDto3c3l4
dNWH4A2qdVg1QtYzS8Un7jwkuelTkYj4SSBDdnk8Sh1DjtRJwyKeAnL68quOXymu
EShIpl0pIv8g71sFiC+kiOdTtenu05/x3vJCLSgXOpWegE0gCrdcM5OGbUm90S5C
BIQRXPOWEUTE0oYBrb+5Qn7Xst+vdKupj5LKfSMuQt0r7PAqx5ERiLpNNaIV4ZOV
QmgmPvizp8qDsAtE6LUV4oP9Mp+Kf/5nbJN18HPuoS8xmKKykzX8lEqnE1Ekla5+
pB/jtjaVbQ0N0cjkbLUFVA==
`protect END_PROTECTED
