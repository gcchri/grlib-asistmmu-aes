`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8OhbjD2bBRweKTUPEA5g+fpTTAlFqHo3NNVFMJqSmJ9Tl/BbBxRRXR3JIqm/1j0q
G7SqHVo0RBDPnDqX8+BlcDnX5oCLwaZ23Ww/wZOJsklv1gImAXfqnq3lZ+1JrvbZ
qyYJ2w6jJRnIpO+puT5xHVnjgtt6pm0hDMuWJ5iCkRJ7QBtgbSScYbUxgJ7HW9Ds
SomGK4M89RXHUs2VBEed7iCwPlWj52Zwe+iK3086NSNyoAOrrNGtuYHC+YfHVqSj
jV3dNhMpQz8BJcGO2kUsNH4vA/1woEZRIPz0VIVXA/y/E52BnLqhr9djCti6NaWH
7FTRGCZjp9SxwIRRIs8bKu/4UdXOIpEMTDxRsSnOePvfDznNq84pHAANIy7dwjgU
WmlDLKn5L9H/LErumOnXSkeMdpj2D1WZFWw6BGoCu4Yg/wzWrdxTGKluTEEwmAnJ
vZmzV14sXiCB+MRyFop6oizn/PkqTXKt1IuRbo42u6OyO5TZdKP8DYcRdt4XzuTq
7dGZ2ZL+JoPJ2jNSlZqX/etX7cS3lEuzHpKpghuOKImehd3eAu1YtnDhF13aJCh8
EZV37uJu5tnOWPe7FYhrZkRAtImaLmbI/v0Fh9lV4UqtbOqhbFtaWn8KJhs7VCLk
zzbivHsBZClJtXaq+LoACLPA4nMVz5iww8bpFC9qjMqy3+Wofxe+MDMn7sehO4PQ
ecJc6my2Jge393bkwk+90JZ0Gt58meP1EHrz8gCa0pc8PHCtv5oOrSPAnxKLDtxa
xKRfykYZ9fQAQffcyw9Qg4D2KNDGNF/tG5OD/5LUb7VsQEob/LYS09WLxU+NYYKj
wqirrMDjSjpKHcYnsmSQdhdD+irkBcXLR8VM7jfd+oKfoZCZdbJ9p/oDK0Tk2uGk
3gtA46T3t3i/dU7S0MJcJaUzKQb1iN3IP8QIzFs9w8gtjfj4fN4yGj5zHsjgGb8Z
JkloxtE5Y73qez1h0hMXUxsIxiQpyqnzyrWxntl1om8guRumf1XP49xe/zcOxzEp
UI2YZPaFaMFZ2W8v/tE7iLS+be33maA/UPf+GRVVkVMKuHRdDnTgdq1EEu5gLLCQ
vFJLrPJ1kiYz1yuity9+8vbwaQRB7ABchwInGCMTpLAco7ZDL+xUyKEO+ACcFk0z
1EyoIaQxxJfBgTYnOK0jgvkOhTJkdT0IczXS42YM85EHZGPfmbEhitAWvhu/zFFU
/BJDSxIMJhtwnivGC0t4T8jzx7bt/yQ0ay9ZJY2yQGA0oMZrbegbyZV+4rAZBLMo
DSJg5OotLQZSP1YoBfEknqV3UclycW5cRjyPAJ5IFUL22XY48s67aY1D5AfKSPUF
s4GgMwqWbSx2LxvvB+1Wr3SskmCJDtODaEUwZbpI/YeuVrcTEk8m4VOBdQGJE6rd
wGidyOUaWiP160+Bm26nVfPmqKy1IU9d9BXjPM4b1gXEJ3lG4+7G+e+Rt7+Qbqh1
9bw7Xs2AsW7bib4Ffc6HvjixC9V2EKBD7JzUYd+V9iTL76Pssh0XqQfDbAy7444r
+FuLJVfLDIoFGixOvhT5BibbxTKz7IkPXLC7+ArYXpc5YFWl0x2qMWi4iKn9GKjf
WyiAfwMdpgKBIRnELc6VuKGulfNXh2frhAtIVLCOOPQ8pO3svLegHBvzAZaV4eS6
qmLVBkfcXkZ1Bwb9nQwEmsTJ2zVklznFpwTYDbKS9u1sLL+EubSxK4R71dQWaZoT
UlGTlfm9urNj/LxTwwwSEzOJ75hY3iNq4HLq2dcya7K6sMADNVxKuixj9mRKHS8E
XR0Z0Pt9kd6PnrbF8i0aaY5GSQA6ksFyLWUVEY491tZYNGpVeEeJ2HCglOU434bA
KJfl3zVl/+ivCYu/pGiihFkUjrVunaOTs5ntZkffLQsDNLzSgBE91nPoMyEnTGi/
ORbv06e+69dIbSCw1eEA0Q==
`protect END_PROTECTED
