`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
51ViGGUkWM9ityChpAE2LkPXfO3wnqXz+3kuJxQfDCyj04NN2nFiZPLRuGVyQqj1
FT2hzezNoRgdxTMoekWAtTqNJY84vujoOvk9hNTKlAdYcx/AXIORnBVRPaM7xDol
2Q2vXbziWdfeaPhZFStbDlsZ3ltiDBEeZaBdEKXQl6utGiXSSfsTrnAD9cNa8J6P
+9A6cInwhTbQEld9Jfvt1GuySkLm591rPdaLeFulwHTnPuwkEWbS92K5ruY6JDJ0
v6tP46yL3rTydQg15LY8t1dsI9asdoV81YlCLdphlR/DpvsGjDBzRiu/Fgduxndd
y4ENQ3B2Dpg+MSn8Kw6ZVaWrKyUoHwfPDTh5H5zWVk9giFeF4xUmHz5vVI5rH/7D
P7Tq+DkYGIfH/TSJ8qXvZscfMJ8Rrpp6Xl9A1F3tO+i2eHQ6mW6xCUBEXX/FiDHh
iM44rW78y9uByuqk0xwIbZTIgCkvwmEEqyEV0Z8aIK82Y3PPUE0YU4rwoQ0AqxGm
`protect END_PROTECTED
