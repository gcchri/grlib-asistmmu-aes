`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0rFkU62yFCDP72BJMgldwISW+GbMYtnayqDOQ1B6lFQVLlyR7cO0xRaTKj/iYC3m
eFZjtPgLRasGBoG1RCMQvCUzoIOmqoeXc5Y70f8sFndcfuvZnepHsdVSAAc9y8rk
v/lm5mJvrIVDhij4gAMStZqgfRLO2z8QnLKDHvzUPSaRVD7z5aAoJVwEBfXAo3I9
f+dIBBF0dmSLCKVLFyw86JnxfJFnhFIjJLBnzVoyPY0emRPv0wt97iAKjHr+yRfe
sjmFgXOCKOk7VxWLBSYmZcPkyxII+WRYDbj/7+WGROY2+8v2T56ScyZpxL5/4WLP
bzxFum4Z9Jz95TxIAfuHZAF/4ehN6VzMbEkEy5QQFEGzBi7OX0yQ19Wf9r6AGDHV
jck3hEcP7cieKuz4yj7c4Hz7u7QH1/j2QPI4jg1bFm9tJVaNn27IFa5x508ZrjKU
py0MiuBZMM05XdLtbHjknwt/fDfUYkrYeWbbHjpecvQS2RiENNJwl2e1IFdwqO+R
9qo/6+NZSptNkkrltqqjPfVA6S7CE1u8f1qvjD5l2h7dOkLLl5WEO0qI+XCQy0d1
Zd8jQfZKO5gHGci2rDvw7S2VispfLDGLquDvakZ8a52OoqjOWCnV9uxJ1+xGVIuK
mrWBj0zTUVoMHJZrs3Kme6mtpCNH7FBevB3SQlSui4NFKD9G0EH+ebJvDn5V0o+B
Tn3BaXZMEhv+awPtJGqDgkc5Sm6t8yOH9Rcs9HFYCBbSwpvodR2Zf9OCrRkqT+mR
Psgs6lcbaeG0NfiKMTa1XtiKB8sgF+zFKnKRgTX/Q334Lc20sobdufq6+ntSsTSm
/AWFBwZXWPePWps9AhUXwWbtUvodYH6flYwOzj501nE0vie+1lwRGudlEd/Iirbw
ovU/nCv8ERGVAdBKl1vFdkMg/2RadMzGAWE0quVsgLqHQXzD9QSFINAV6WZffOKR
U0Dc5dbNnJCt0EcnusM6cojBZ3Uu+VJ9asOCkTeerJ8KsZMeYOQNTRmKYuDLh7E0
t2qf+8dvg4vWbnRqIL5f5UbGh98Pm1Fis7aKIw83DF06hwsSOzGYdb//5RUSECIm
ghiIqZ/Du47q3qS2SbdDPImb5rCSw4ztpz86bUMzARuUkUNCYf7qATOXzqoG0sEg
0V5MbL4AYYcSsjW/ggSLLO1ORbV83KO6bx9DtWGmJuLQccEd5DZq7wF1+tdip3sl
l7DK8ApQCVVRYKLH9iN+Q8a2IeIBnBagS6fplpc9kIOgw8kDWMK17XfPTNF2MVVO
8x/Vy6AHLnp/hSXRcCZTyfRbhlKdgTXYi6dEqxBGBX4hVcQr1g7giHZL0Iic/NMD
ZQ3Xm9EMjwNGOr0cUZ1d2ohv94QmB/FnjYZceiYMsgxT7VoyBTZvckkuiZQwl/fa
k/LFwn4raPLa0j9fPw8F75WkQ2n73CWJvTwb+X2sFzi3Lww/VGEH1AEek69zQQp6
vv6J/aTrTtQQm6YRJkZqRhd4ZtBo+lFEl5Tc0WX43gJQMfDMPI5Q3wK1dq3pc5Ef
MrzSYkkCrv7XGhGeOURnLj4s5PvOFD4b3kMr6nHDe11y/Fv0qGLaTykGoegdS083
cTLOUvAzjkY8c/9JSfAhTH1XzmB6a5Gs5UKFfOAwhmj4Ejd/euAZF05LNuxo2/xH
veTd7PrBAcVco1X98ti1jIxtfTTJ0MWZqgs8C7KDyfZpHSBAMjLEL1BreldK+z5Z
MkaPUKwrfO7m2cj7gNvya1V3IQzH39FwpVvChYlBNxyZiEoNS2xoVQrOdousVZge
Sc6jd76KvITB3ORNF2Kn/qFTwJ1F9KesSRCrM2Uxv9MjK6coZdoPIOB7k1AsZV+A
c7uTN+qpTJuAQvoQ46VVkOeWksLNcKN7jnQlgP7OJrjAl644FKkhm+74//PUtQkJ
b13IOL27N52EPnFHW75ixs7mHoGS3soK65SCMakvwVzPWjVu0gugN6GFNzV7R+J0
rY6fDWdjIW8DOz0J+RyALVjGG+u4jdkuzlyfvv9d+v5nVH5vh/ft9ZzeqEm1q5fD
JP+D+V0zFcvXCdxODeW5vcdaWOpxdgsllHiBvt7SjdOPuDTOI3DOPHvKMPmNqnAq
0tipeuBxvb1TTqlwfruRzbuCEsOdTMtvVgDdb2fWjavNVVb1ya2AXRU/tJCkNeYn
z6yGg0oY5ap1UrahsimxMUZsRocRzmx/7dWVOMBR0Vx7zYcSFD5w4yuubihvhdBz
jL3cQ/8mZlePouFK1uEIBjFzgKo7sli7cBScKZDEjvAH24AENV5bW9hZyLwJBzOy
46ONBWeKPobVGxNtYZm5paLENVpybKAFXn7mn3J66VV6hK6ve8KofwlRTMvbuXg2
pQCaC1jpHlB3hNoiTils71JKSDg0wWMZvHk+SKWGu6ImixohZcMFJ5x9dMOgcHMo
7u5GdZridSozdpFVxMkaY5ZjyEVec9T4vA0Kxss+1IL0tD5hqgbqCyx2xxsxXBiS
RrFKfpOl42svurc/j61+hug4kNRTnX7weQA+HDmDm0UuMeGFoYqvUurB7WM7dbCG
GLzciSg/zYJX4lRPRgr0TNHO4u/aaEh58LyKQ6B5Jp0Hk98nK2G6FjDg+ahRKRSH
LEogeVOex8Nprjl0JPWKVNAcg+XvMnmfyyBnrTSDFAfJZX/fRxxi4ZlW8f29MZfg
Stb0XokkdrN4HfKH0qS1syyu0BPua5YiZzMW0vKPZCQ6wjfhhTqUvneJ3xwvSV+T
/vWMlpME6pYNt6iSp/t8OawIgOpK8fLeogOHSLK5605c2MYHfnMopjTEizOpdBCb
IOaxoKBVlYqQW7WigTloUD5FgYSdJiwBY59R5X/Rj67NxUEBNl4h85Yiu+15bKj6
vqzCdOvN4tzDaxoBsc/9oid7RoT3U+wjzBQs6MioCrvFB/vg9/8K5fyA8rDxu/5/
QnznnnK9nns9GcxC614xX+870UM715wiPBqu0c7dr2bprZX5nRMMc8wfia6vvu75
Y3TJXx++EKKrwVEKEFavJfepRaJ10IChUUfmbyZtN/sfo3o5q8Y63Dpt5PKcNMfW
lxOYeVEM+Ft0oB9ApjlEpy388rp7SOz8n7yK4qCqHCiaqmQ+fTYq4fHuL9xisNXW
/Z4DJ+1gIVhUvRHbdN+RGk4L09IP+J/+Lje7BpLPbSQVN79xf+JbTbWsfOleSVcJ
T4gDqN2HNOEwl9dmAcUYdhK4DfS1eJwcGv4hKtFfUqRD+CWJ2jm/WOZgljWllMah
9Z7UsRoySDB82l/2zGW+e+jUDp1k1mOs7LGPIwuEXWEy/w8T946XWeSHl7XWXQla
lMTEle1zE22JydKmlAWQvI3FwBXzV4AMZT4XgrxYIPd0nR5/SE/RLzV2ZoNbjyV6
gXttBTyJYwGlyenaluB8gJ6vLfrx8uL3c6EZ7/wkfUOGbqR9dNEqFqLQG6EKaAMJ
y2Dsysp3nL6NbMyxZNWPqnScvcuD6yK9xyPw+uvsYkrLgqOh8L7EPRmC1rui5EqM
bAFmPg+Z6i/FvXlcy30cwhE2+zp6R5MtqA4AACHQ9qrp5C4iLFANzYSjYeRx4Cy6
wEEhxxy4winqWLWZhKyalWTnnNVFBs5lREeSKo3xesVDlwUfNSgd3KTyG3asyLua
zn8o8VJYuMQm8ynto5AkvSFtn4Csa9NiB9EnDo/JanpgH+85CPccs97geRhDD14G
sAxuQGkz/QMGDaDIeVLlgcZGLWk30HEWq+vDK9hPQD/PuwHobFlmR+Tsdr24iUAo
5KLD3mqAsoxfXa45zU0EY6qEEj9U+LCeDhpB7Yb4SFXt0MR4gHqaoKsgI8n90wif
YsPPKutIl79dr6Y3Hxz3/23di/TKeQeAnFfeQ694AqNThF91aKmqbTmdtPL9klvn
C/i4J/9GsjyV5MTfcx5YY2+Olz98AjbFVCOJgu0WXrM=
`protect END_PROTECTED
