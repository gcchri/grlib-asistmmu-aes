`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MnIJDPs65L+adMyEsuY2+fe7CnIMO3/+mmwwrebkE3zdJIsFyNoONI247T9zyGvr
m2jLfywrEK2F8+b3A8kgYg5lUm/n6NbDPz9Qc4lxTLDmVWSDfH+/MlIZwyoZJwTj
sdtntGXKoSu6/mA33xGW11XXTz952LlagjrHjIEe/d6FrN4aUUxfUhhSUZQQ1dZu
KuYBBNFn1NYxCfJQW2GUiraZiOZnS+AltM/y9JvJs5XKGkCU42sTtB5EpaVBLi7a
x0HTA/1WPdSzwtgIIykYBTSusskafN43TJDZKoWQibprcxtJ2YLAfMb7QFmsPaIK
5Pa8eGlWYL8bzAP144FloQ==
`protect END_PROTECTED
