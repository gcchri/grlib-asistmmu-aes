`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3NQ1UeH16Z/Q2EgStJpXr4DhkV9GJXF0pNVPPwGGUXuLRDMcnxbKR4267Qq4mKZX
wpPVWQFXV+CMBfGe8SOckvwt24LZWpG1eHcfy2r8jkFCKk3Lsze0TGFjqCj2qklX
hbSb8tA0SEYak2CEOUJjOs1lA0GKgKa7o0jahsAxs2KviZoOaLR1bMsOh8FzTSWi
8CxaoWtBb50nzVA806A/SxMtm3yfH3fjBY/+XC14NrRaftsoGjM1UUmCY7WjohYy
ugrZg2aIN390a7sFYsz3Gfyv1WDS8OcRcaENdYWi+FqT4Bn/y3cyTophZwglZxkn
FLEb2V0hsoduLHTn0mHqisCuYO4fPV7xf1hVd8he41lRELOMeiflhGD29vhgY2RP
doy/3/ymbLJwDy576BzhI8gjZa9XxTXoyiyDeN2uFsc/pWudt1vJ3v/Gzg9/7CT2
`protect END_PROTECTED
