`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
34NlapcP4qJAc6gyUeYTamjM/F9Lnmd0akrk3mgx6t8EzU3Tmryb2dVDe8UXBa2m
UXESSvGTDL0+g9lyAWtogcvQydst4Vl47lNDHhhTk4rEx9CFM4/jF4BBSjyo1GLl
wVQlohrAi308AkKrAyY0dyfNLc/cCGvcQXHagAMxUj74oIhYqyaRNRwxqH9V1e6e
rlw0OVhFTuI1EJoM0ZI+33qgKyOG42gcfmNF6j6otlgHE/Ehxnf0MzHNv7CnK7bW
sZXtRzbL4UqiGrdAJGky18BYoRqdwOiQjyb58JvMUAUOwoQc4xgQr9I08AXVMstf
cshWHZqyHwMGhXk9347WEipWo0SWTwuvZdhJMN3S97qZ5jgEHZDBzv4PRU0iaZ8g
`protect END_PROTECTED
