`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ht0JNkIsmtZoVJ7I43jcKXPVq1az8iqxQLXiauie/Oo48wLzwBWMEBwWPCT7STjH
vumwMeNZ4Ex/3zUyrDeOqyJMkk4iBYysDinbYHoZ3TTiqf3p4sguXdhbTbZSm46g
Cwy82Hb7881EKykiStjBI/CwkOPuxg8L5QGrZ8tjBEqSdSSNUa2AE0iRBGGucAvt
Prw4JWYEw731Hvx39Z16eedZNFBBroeqTc6oLwK0C2CClzSGB+lc8P1JtAbEshDI
WQNn1fVT44ZkacjFEY/4OBnfbk65Z7B3LF60k+a9MqIo4/7sdwEfNvs8D7LyQNmy
oFB3QjJmxUBoeqCJMR693YqqJb9ZkbKCXXOL1wbi9rqrNGpGD2k808diV07OEvYH
Cr7TuSn79fGgwk8BBWVe1HK0en/smBlvuxSCkVseonv9z9JCUnICISz9Z/KUOD3v
HadNeXIjg+lLu1OCd8ltnY+pEPGbHOENf4dEFKjR3GS1wHN219noT/YFS1s4Smls
/CKM3rlnXjtkRAwG3CW5Umjw89VtS4Du8fmkOuSIYYCmEj6uNEYJ5jPNcyQaBVT3
D16jYdwwfA1xW9+k2sQ7XO1NBfDNi2/q911bhKLmgH+8MAXf4UXj/TIck2o6ZYHg
mSduEWVsicqkqVOXEPUnW6xEzNBHjkamRHS06uwbn9N+U27RmIYonaADQKg4F0Lh
7+yTPDxrR6RyRT9kTYI9yDFr++RmNJVfS+N+WdquF90gQxRay8euWU0QrU5JXfsm
t4hOm31Wxf/s1JnUDkrEDTW0rYv6ofONs2vhIO6I4J1mwO8cQMacV0hE+KGZ3/Zr
2ttcBMSyuZ5ErS9laK1aY+5cykMkw06kt6gbNBjlkDf/CpFjgJMXNT0EDxdUqWUx
fz9snPcHTODJWX6+Hgt/Ox3zIJY42/MfIySPDOlNOI2t6E0QzMbFgXy9gHNaQoDn
juaorvFDncwKkv4FYlXTVtkTMYh6Q2y3nIBqhz988ay+r9YKNvLNqxWDPiUEhncR
hfqfcJcwyFUhfcnjBDJVYALnZ6lMEg7wH2r4NzMf1yKKAi9wYZSJNyJdfLiWAiyN
YG1J0pSZWqLQsnjw+58FVoKcS4XvvnyldQJSiXn8uPqAVUNQBYnyZG3+ZPd5NMJN
e5LVY3Cq9grtyMw+WaY280ug/fKa6hTfc4PBw7MfIdEmdYFmu7Bjh49ureLcnR8I
OQF1YM5VUvjkcGOHXvfTWA4E6eJcP5LIFwfxQmsmpOjt6cN7AlXf5bMFtXfpAnPb
JETyQJfvLpCU2Jf81TsBobtPfwbjHaZXOecDcElcI5NHvS3E4E3I1ag8Rf3Dp0yJ
pSTb4Eyff48e66P+2bUNOoj8PiG5GkttVvrDCqqafZ1fo5ZOzyfKqUJBaH3xXw+V
5J7oNl0hRCcHPnLrvTRp9B59O4m96j2GAnxsYd1XRpVduxq7guiVeRkxIf8gwYNk
ysmaUFxH0RgajKCiW+yM+aNv9bO4/RTcPE6xHDBZILk=
`protect END_PROTECTED
