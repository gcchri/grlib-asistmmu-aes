`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IuhLFEkKamhjHivtjKhJGNVAuYOmWK/poJN4KlZQHqqvQpuSimD+gojCq6nK6o7g
aK4org9VrSIPqUNAkCXwgMKDaKhE4JC/7YcRdBfY/qjAeas7/LylcvzV169oN9jS
p8NZ2xS0OcbG7m4lHR9JYsrFmiaVS6Sxz2HB6x9vvMOUpoTnR0FQ1YP7sNWJQ+FO
xETNeVGeRYEMNy7LgNg/RhTg+UPE/Yo5nnb1reL5bfeoXArC/Tcev4/2DLJPwybs
uPHIAXqSnSdErb3NPLkGwmX4RHu36BpYafZYfLaQVlNtNbWFlRxcqyDxY3I4z20o
7qSFGEo73NkpVmht3r9ADBVZ8rloPabXdaE7f7HHqQuiGqD2Z6CRSeGdPK76IC7V
wOQ0YjFVqvhsTpS651sRz0p6O/DyWm8EzBOlFPxckadg5jZ3OdbKUTl4FBeroCmU
MpQlnySA3rjRPMf+XSqS0WCsulfZ1jNtpqkqCG8Lgtroe3/gBgiCyDGT32hXxZSB
wWbmgg6tuXhHqlnRvIhDHKOXk9AWZ+FHu/4+g4cyKLoUrW2xg44oJRiLe/Ov6IiN
4lSwpf1QA/dcKIv/jpYp1dbOdDkb+r+6bxTcF52BJsrrGe8Tl65XAOPiEgoQp62P
5u5YORrIgtsRiMRZXKbvCA==
`protect END_PROTECTED
