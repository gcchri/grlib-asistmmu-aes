`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
whWxT9Lj6Gbutms2jzvi42HyuBJwnQ/DoAG5xHNl2XbjNs7IpnHBr0rb6Jz+wOlC
+Se5geiRyYfft8OFVlX8wguj5aWOtF6TlgFFJez+OXtFgXm/TGK7yekjJhUqpcx2
nDHsBLH49gTeyrlr9S2m9ZqWmmsPXaMKkAXrXWon5EIUh/0yreWtDKmbqKNyZH/8
7rhuSVNJNwnYz/9w7r8vuuenVaoxMYnMQN3ETRDIJdOlMpt+QXTh9DdMAmgMjlDh
AF3fPUosq3VIstiHYLypLudOqL1Y/Ek6JVrgAcFLqUNByLBU6Ns0WIZ6Y5qAc5L4
tJRnL09R/c6QIXOak/Tp6mnrNuew7aGFfz+DZ93ZBZ5BP4WnJ2K/panPOV0VOg+B
YMQjcrHtw3MS1O4oNh2Z3qlEuQAkvwfvYrWfH0txaQMD8UMvnsIW3JomeT1Vk1tM
5xzSrrsQK2GbdA1fOrRBQ5j/ycVoA7v6FjKU5RsHsLhlf3YDIL6AYWL9kKWK/b/Z
eUhS2q0kOQFbVKqysouOThLkdtOiq7jEk2+jE9hHo/VFJYZ/e27VNSaBa8fQntq+
sjCXlbnVBV3Ow37b+4mEDbNVG4NBb+xkKYObWqen4oyraZP2WkJKHSWH2x+Yf5d9
bIvVjNEdfehGw26J/jFSzu0PwpvE/KCwdY3QJUPVdFQ8wrbmWBTussAKP97rRgbp
JmRmjExlpENaHvzkXZECDAOqWho2mlr7d8b7bh27t16djLWw5IMDpsULM3lMeuuZ
c3DmLOa7KB4H6LYxKcQ4YNbdtjtmtj0A3lS7W5Hv0xcxk0v2a5WRfeA+oflKqXbP
tRqLZLYhmQEfAuUEG2jkd8JDVW/gq5HqlucSI7IuRfsIQs0MY+EP9Tbs8jSedsAx
wtOiBYa6PpS9oqyKza8cJEAVIFbhNAKdsTT+PH9l7DV1viLjOvWo9hy4P2/eds41
9RIFZWexPYeeeB3zARUjXkg0PFJ5ZAJ0gRp0RBNY9pJ6/af1oqXHit7LfJSo4DuY
44uVM7P0ynjmn4LGW90GBlxMO/U84hkKaSP4mc1ou0UVgyotCU3C5+r2fuk6UxUI
NJnH0NeYE5QgV83gCmNgn6slarYqVDEARZoG71rAHbLy6gZlhxlYAjWZbls0Ingp
4/bW80FOVor2QiiAk56nsTGvGuoXHHF4CpWFK6qOvigTqTUITITSyObVEiOcNReh
04pkfYOeIZDUcjKfHjWauo7cvRQesO95Ey7WlU73Q1Lm3doM2N/p0cur9GGCId2t
Ihr6HpSyeGFb9Uv4dLf9vtV+09PzdZDZaRFj3JTXnC54/Xwpc6VVghTWoOILg+VR
uBukn2cH+3hAppjtNnkAX0778End2SExl3Vg2YNMZSab0lZwxNOSHYNbbdO8WRZ/
oOh0W3N5k2FcVwhKTN7dUbkVBCTJ6rRhJwwWrWCbs/NdjeY3HY1KOi6e/Jv+hqnC
Xe47kxIJIDoJd6Au9/Qb3npXHaFPelxUGEm9nkr6lmgnaIIpYahuJiire+91DjJm
FmH24sSDkbediCMRqQ8Mypcpbwx3TktgHrsznp1X8vyyCHai0bfiCvfFyxmnfrf/
SSfec6Ahd0WusvRxJfsV7uHDw2X7o/oI06jc+t+tDLYmd/K8OsU1xpq40P1BGvoX
k42aHPYXK4d/Cxi7EnCYCnmSTctXaNS1WAlpYHZN5RO/YZZiQCtKQhN35oMwDtxX
yJsCOHLvjhJntA4kc9GS3WcYJuDEc2mHQmra5PDkIoB6M3hUCJ1ekc4bfPUkDW6S
g1LPHn74e8IktcRLMW8QOnOynHKZzPF2FrpUbxSeI1/MLD9/GiRJdvm35TZJX5Kb
s6pMtovXGi/La3NxE6pg1Sl3jaKPn62+ZBagGqfoceU3/a5+3/RjA7OruLl07VYF
We2qWXAshWRLZ7X8o/PJP4hi1RSEBhDteQ/pQvMOhr2kEyOuQFTsBigKEIZeqC86
4AIl94j1lFPvIM6cnzYOuXdIJw67e/spcOvNNPkxvbfsHcAah6YmksPen0DRMkyK
Y7ksyhF6fIv7Gf8Ruhbl7MdLMfYho3iCw7qpUOmahwMTMOHaDmqawf8ODt8SdzTE
deYvlPdy3Ixwv8sOlp6A64xRqHPu1+lb8B5N8PfO4oV7XZqduw7O1JEA2fWvCQMA
3VvuFloE/FRE/KfDWsUcIWBSSABZ0p2hbrlYGoevZshhnF03ZybJUZJCV6lhxfVQ
IeLiAZCCCw2Zw0dhreWqu7a7mfu85oT0oC+qLRXC3XXYyQGvrbsdCFYX9NZCHUKf
ykIFCoTyl8EJievBWKyHmKdh89SOzgQgp79iKGiXiplVOXz0zDECndg9rDYJAVDO
WnvUbAJ+wqLb53Px6Hq+8s+4wkOaXroobQaWB3xPMa1c3z6mebpoMnaxTfjSbIch
coKeGm0Ub5366IJ2xB673JPBxN67SOjUygW47Y/A1ziLdTC3xo02NQKL6KRrWX9n
VBicVZbOaWsDIlVIoPOcKuQgohE9Ch0qLQlWnm+WHglc8Oteqi+UfpGqb3emC80Z
S3wHzWR9EPWzR9TlFx/18izCXmr1swTUzFAmO8zXhdT0+YemGpd0JlrgwBBo/ciH
tJoYbEAYdKYoTO6Kvq+Xtmk9kLSurvSoDeBH9eoznBUoidREhVSjqcWgkoJpTe2Q
geb19erJRFVCK39zz9ECt4BrEZSI22QUhnGPJYbLFNSdLwW71H+zsmf9DDVsRZ9a
7/IpmGWfSqkPqYM9mnZsLanaOrTgaU0/AodYOLFpN0D9VvaI7PXN78D4vGgRWP+9
9Ix5MKSQ3BZgqdF+a27idqb9ZdS9lFfvPjMVHCPzi11eSBIwkSFcLi+srw7auazJ
drFYDEPxWZy2SULBr8FHpKshBUAyRym7flHiMF/LWmB0z8ClBlh+tOksMGigu2r+
yIqqFGn5H8NAYjEONwDmjWg71Pm/h5cd0TD8xf8+tJBk6oCSH6eqE21Nd2TpSGjs
vO3AfMtP9VUhakwbK4RvwvLKYaUxxpPSnjjpm7EiGc9VcY9YK/UCKbKhOvV6zbDn
UfIhLlTS4LSrXpgEgvMalRUY8aeKMe3NDAP8/J1g50p7b9LSBRcOokNGVxLj17bn
bhp6ndMOk/7v76cZGsvueckBg0CymxlgSGTTDoW6+b058HVw3/JJBMYcF/y4cDgJ
Rr4snDCvAhV00L18osvS8Jr+5zUHIrshPGtnLOZrj+wgD73F6e1OeTLsoidKzhGQ
0dT3dwEVgXL/kNgzMdnRjx8D9fMUKB3XZIFYB0dLvRAJZRszSAzopX9/VcW397+m
yXvt0qyqJ9gpanWNHSS9UF397paM+rT6Pfq6PeqzYKBrqJJVk4qQkOJ25eUHVCFd
iii1g6OuGf6eYJBgqHRL5RVclinfuV0QS3b3STziyhp0ATiQq+wDZqm2DvXnS8qh
4oGTJ0h+p/x/clPyLFgH0BCpcMf7uLyNth1bJob5G+KSJaCftbPq5shMG7UoTYYH
ZyOfEmJ9E4TAPtKahdZa1kSlrkeeEkmwZaKL02an+hkh9pQSpH2HbLLRpvZu7xXn
pcvNwZS2kvPCwSyz9RTJDBYSRnEIDru7fYbfuzO5WikAv3/lMoH6qvwNGNJpNpvC
YFZ+hMs9z09kqTkpJu4PdQpeGCePcTq8RVPPVigYpg509i6DML8uVyWXB1LCqGIs
RNz7bJe5m/9EW51Ua3RY4RzESPBtykGlhAsDf5fiicXmtAUNe/6z9+Vam+yty8KW
9g2KKh6kqyMw3JXV77U7AD8m9EefKQhipUIu/CRuf57N7WPGOb5c9alxmHc6/chq
rPjA+14RZGHlNjetQljM0iT4QuUdHIOKBZkeoiNiDxR0u71dgFNezQAtSwyUSIM3
mRPoS9F7ye8Ab6NigftUXUOHZfBod2VYsI5bv7tCQm9orDu5Ij47gaZhAy5gV9UT
mtOrEOR63EyF4+N5PKvxeA==
`protect END_PROTECTED
