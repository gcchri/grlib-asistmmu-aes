`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/PKL+nsiAACZXWqUBiYsz0gYNB7k/52aEp8+qDTvVhXXy59p/wy00gNxuEosIEvO
NLGzHp/TqM7eCZbYJyrw430BoscdZzgyvSshdEx1uxl1p7MdCsGDf8hrTsHGmBAh
bC/oUwuLtDyiQ3R6PseCkZDjrBp1dEjZNJTupG8FXszruwgzT5NeXOO+sasFy7km
ljs6CvAX+rNzsn3vttPpiLooI6DrAH47E/oCMLhAaPuH0gVf8S32kh2Q3qdJwazr
aJqc4pjb8HKsYO71EBkahGJF1IVep328Y3QitU6ncQk/0w/lqFswghQIFLY7UkO/
nEma83bwlH4glxTBmZtiS6e3lRz7moVt78o2yKNzMRmiq7RRc0MzeOjyf2jVQ2L9
jPktcQ6QyNYI0muc2CUDp9F0HqU9RkAOR91zjsXpfl779IrqIi1C5utAoFF+9ry/
BoShHDx4xsHCMh5+GiDwbDwFj6bm+5i/1xkXo+0Nn+L40unm5M/sslOvgNq4raaq
0o+pJGXG3N2sLX7uOTHU8E5/A0B+m34ico+dc4tqyeY8Y6nh8Z7FXk5C8cxzOo60
XBfx/pt/SkSNSrUWr1xJUu9wvZhsQ1LwTWtDzs4GK2phjpnp0AUvMs2QGgzSp0M9
TPD6oQX0Gz37NzKXTOOGEAa4ZLcfzVRvQ1YxPJ8ToeN4ErmZB684HSwTsYpwphDg
d8/zVvn/5pS7RyJoE2OyXF0hAo4zhRIahjDMOXaOPlQV+oZtyuRWKOnqcwRbBbl6
Hwr6mDjtVjTR6bn2yJ3G+w==
`protect END_PROTECTED
