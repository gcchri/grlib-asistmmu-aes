`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oJFlgbg7XEk9W6MQPLZ7b3TJ71z2hYuqJoqnvaMTWwFNhJtLOwmnj2Dpp7VflN1D
QdDo9qZtyT9Ia3OZq2m750cG45RfWFvP6C9jVWEi1/4cV1K6Dom1L1VitR2K6qDm
kOXlVVXnGwUtYXB8pJFtG/17nTHuf8S2laGhfPFAh8P/c4yhhup9HRHJ2uowIVh0
L+377695IehzCIOEL/fLnLyXlZyA3GXle3wANH6QluQfWz8XCjOS0e1er2b7vg8h
cR1eivFK2FkZti3VdHO5NXMcyP0vPhqvl4sjDH3ThW/0b2hMPruPDSrQDsnK4c5V
TAjK1zb4jZUtsoSBdSrhkoNn9tlu5g3CajFTjtTnGQ4GHlBfeubolQ1O78Zdwltg
WGNF6Ib6gV9g2+QqF6b0AJtVYy8Vi5353mv9qIAJ8AfQHWd+qKJdC4rxA6wOoyut
c5NCsJaciqyaVldcvI2Fgw==
`protect END_PROTECTED
