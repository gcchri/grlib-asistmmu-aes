`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V9zfTTlOVzLj4ht1qw0U23Mybip09TJUMd0/nouDiRPiNY5n4lyqowawTcdv2HDI
u4Dx6j3MFObyCBi70J+uBiNFzQIw3BPbJggvheSSeWPXxCub2aKOpAoRkc7eCCYG
b3WwoKQKGbpxoOjFlXXPqkMlLtuOmpoExaXrV2p+Ghf9l7VLsXmjMpFirr9tVAc2
kPkhw7vwZLapeS3mNDIC5LnachKdaor5Sv0esclLxXWe4JES++AKulHoBs4sXBPY
5+ZwGYOcKlrwAQ/+3FS7IvKPWxRhCyb6hH7KVkvMbMF9NnHSqbbSC70NgpyqMb1o
usD+6Pp4KKmjjzfA3/pqL/TLHPGgaZagaq3Jfq/Xq4QDwMIfInZA/edtlcAImOGz
r1thYbRCrbogWHxSLyZBKeqxCedDuy5slslj/WTfnMRYRET/ht3Q9Pg3gCf1ddRs
9cHtNUxIgw43rpVPtm8UCC08OMXChdliA/1jzoMMaoPXSPfJneZmImY7BWhLK+Gv
`protect END_PROTECTED
