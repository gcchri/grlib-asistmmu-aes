`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tr6gvEwfbBc1VmgX199JQ2dj4gEkoI/X4q/WNmlogSi2xfI4/hfRJT74w3KGboli
YeYohP7Nq3u8EvgnViletQqUQxLum5mxxG9felbB4JWO5+TiLzRvDCJnC+exYZF5
JXcfJmQrYPXfrTKPGQk2qfjDnke4lXQvetZSnV1S0Uso9R3Iz7CtODZ1tMGRT68K
0IuvXZYZvNlZxEdRlJ3toeJv6E+jR16auUQxyBk+cmTy3eo4/esd+9icnixTlb1L
GJTFpX5y/c6mpdnrZxXnCE1InZvRhl6bJZpVONSN7vRCv0ka9Nj/mOWUpHii17Pp
Um30X3imdlHsX0vnSvwqjw==
`protect END_PROTECTED
