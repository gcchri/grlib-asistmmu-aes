`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z9j8jRyrcHpX1kxd4Zeg/9xjl5ZlYpNnWo+37t+5MNylS1/iw/50v7tW98tt+8PE
UIFexA8KgS1WAPnAGFVKuZrS0+llrPoTsC2lTdxsfrdqM8fhGnlj77QjN3hjCrFC
ZpDfkYpHUP0tp9dOoa8zBaIatZ2YxMczKYFjcBTM+jlwuQeqggzxlLm7Wll0bNkt
yaPGQfYagEeML2EEoTsj4g+s8RPDPA3y7UfsjgeXwInl7X1NHgzgnKH7hWb8MnOa
B66ReMuquq6fAh7x7gw/DvN3Ry2ZV//aK62wT3r/Sa2eijAj6dLL4xM3Jksp3RDa
aVnilOAD+mrSdIsUcO9KAeEhhBwIvGNcpFU+/zDHecktTILT3BCzcsdOPiO4wLTl
vHJ0CS/Pd5IOmnGhw7awog==
`protect END_PROTECTED
