`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4VEcZAwaC5TDV5mmJXhqwL1pyMKUirFt2l2Vz1DNKEAjwEW9wY1XX+aC6bcL/aub
qgciCWnUiU+MNJ+Il29v/jyG7NP+psGjpeX2E9pJF7pKGfGmU0TWcxgTvY8JNET6
zllH5gFygvGka9eVKqZDc3I0S6r2ZvQaGCeFYMBpEGY3JS3Bm54kSUCG+Yje8P/K
xxv1RPkMUbwL01/StYml8ft9WI7d/xOHtT4leggjwrmbWSK44qFIiXSqyQM9cvc5
JnxzYwHVIUNAOgIQTfNOru062VNRohzEFQhAuc813x6u6XMVXEny6FwERhrkXBAF
24ZMSPdY1xP3xukWeCiJ6jTXMpBbY1HFtG40j5VSYQz8GdEUq7O/77GuRvbUI66Z
`protect END_PROTECTED
