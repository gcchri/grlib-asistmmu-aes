`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jZVw9k86oYQhCKHj0ZKLO0y0IV8iCEN+c+5nRkkMPAIM478haBY2/2S674SjLRxk
JyAXSBsJbXeFO1UgwSFFTohwXqh3R8S+sgEz3HWHwOE6Z/WEuuJYbXlIdmPt4j8w
xoQTDNAMGNm1LjcyyfifKa1IRj+H87r3UxkTsF2gYnGLh63enwImlWvWZp/lT27d
ehUbCVzlWximBnuAbmc4tHr2myN682OR5KmHfdR1wjtyI2z3hBpx6xkBa6Awj6kJ
xxOiv8Zt9+oqLEHeCH2wm9Yvq3CuecrPKkurX3cao/fSap+V99tZsGzAWtQWBHTd
qRCkZAmA+aw9kxGkap81vYaZmoC43VLoM4CFrH7e+9ZsVm6ZrBE5jYxomeeZdr4z
FjKDULk5bO68cKdVfkteBHwwTPHYWhqvBMvxcd4Ju8jq8qrJdUbuAFC6r/5b7XiY
TVRh9qMOUy1AZWKU5NcmpO4I4wxWGuDLXX+mBg4Hk1P/iC3qkVKDBT6p5OoIXckR
cwYEEbVP9l9qa1KZffBz986glKFGKJCjPrPBkSYCVIpOYtL5v8B8mJA2W44H236v
xFtFyUWr17ya2qGXTkDVfmbwMjei+EO0qQ+53+Rso2RFMIzsiI+zPshwppNt2wKB
3PGalh6MxYrgt9T5PA59hGO7a3LNKzFFtwOXQm785mtkAILC5iLEKK0pZ03Ka4lc
qCD0J0WVd7HkSifIGSjZ7g==
`protect END_PROTECTED
