`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aVeqzg6f9gNEHvDF88WUsPOkvXumOM3XbGQ0WPl6ZX+thxuJ29/Q4gI9ggKKXIJR
sCpNIkXYHkoTK3Mko+YKLbitfcguT0gALjrvtqIZx1euWFgXDCROkYmmWlU56b57
Prhs4acxaE1hpbSZSxu+eENUi3+aCavVj3Pbx9BJDai8gBxWFcfiq7cIiyfzUzFd
BBB45pR9wKJQI3h+E4/EukhDhQ75Nqt25qdLfKlX+sUUoZtPC2j9r8N028oNtHP3
D3YMhbdA1j6XNiRKMmVJoRX69szqrAbLaJZlDFI20Eu8/QkYAW5Iw/1x8Ck9Wu6L
WZkpgRJf1nareSHuwxWTkP4Zw9/s1lwnvbk5QTaFpo71zB5fY/PAttqvnmwHAvPk
ghjaGvoeOPVLQJlAbFr2W1t6NeQ16GMpP2rSvhEQuA88PP/pQVUr3PAiepUHPsJW
PNmaTT0wWl1mJiYXN07dbdI/OPvKcyd2a14LOcUScyl6yg5Sjvni2LTlWU7+zR8q
f7C6vpa1z+lqlPTpUY5+AXN8O4ae4aJVqEBmZ4alntO1QYlaEjsqSk1r1WURYAMr
`protect END_PROTECTED
