`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uH1nVSamJWfTGC/AX3FOyDXwyRkNjkF38YzE2E4Nl08Uz56fnUbjAgc3UKzTQ+7z
3vSuK0QggomBTelwftGsJlaMI8bn6sWCYX7z9EGz+0+EBFTu4y+/XUkjxxCLnFOD
Rejcjx3Vxw+liIEIktBCdWff4x6jaBlVmnIRMis2tv3xOb9WjJKAHoDVcUDZTwR6
FUM/+WO7Y+bddiFa9zXquFyDCpnFxZcGgS6JTEUx0eUJkxIBwUXQ/o6ELPBt+eGx
Dn4VHK33lAuaJupF75PayRT2SczaGnihbYT1O9CanCglj4f3VwGJzMhpN1C0IynE
tkGUPCMHMzKi4k2iQVWIJA==
`protect END_PROTECTED
