`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kxH74n7niXenBSedbOEV1zGQSWOqUQM2wYk0sVN4vBUma3V7DPBYjuhFGhUEgUE0
8JzXyfZB/WV3q2BWxlfVEg74K2GlmFzSfMQzdnK7VJpeHr0B8PtjtBbebjXYuCQi
0hrg0FlVWZic9poPLADYwpNDrrh4z0mgHDAkSe6crwy7Qw+RWF2ho1d/fx9SKEHp
IIVrJTe0alLk4ECAsOCPU0/6M341MuzghHB58+fFxCuINgQ9TZuuuuw6fpkAOhkl
rKc6959OjdyjlIGEFeHBnZdoZkG6Uo6nwJ87hVW5qTYvyWCLGwD31v9CCgD4dYf/
55F5jDGhayFgYN7wFkDcTUUUPeZvdYXP5JXZA2ld1A9pECZloPodMBJeW23D1RQg
PD0VaP+AeWGYmfHYBwuWAXEAOeGhBEjZfULNRO5JuLNxooQ4ODS+ePmQ+1v/kU/2
4leFKy5zl0P4bMyWKh3N8ye2Iyzu2gt/P3m+Fbew6UHSXfprlExK8GkE2VQLh0FT
EVhjXSHfmqkHwR/rfz2IrhNjc525XOtzJCTwv9bmyfdrhHovr3M7XppoygxhTgBA
+D8X+Lkd5j2s/0LAdj4Hhqx9RoWzMZquG30CfxjI7wsfY6lBcwYTzMOjxurMTAoW
RaP97wJzTZWhWWGZWJL1a6SSg6OTGQwxMze6q0oDd8fUdFL/YWyTj4CH/KqTATvn
2v31h2gL2d52qaCxlqjpBOlHPnWVGP13Qkhg2xJKMZu6eGDNg47BFVG416JlbBFC
iWXga3phnQ/L3953i9cmkBVYbClrM6PGbEGYpeA3S/PWAWgGCw+EHouBiZnYfVqK
y2AtY4rmYJ9c5EkLhR7HmbAKTufDA95lhsFlHvral6IaF4DDWy9hqW2O0K/UxOsP
ukzoqD69LCQKMu/8ZGbpGOa4wMwDgJSXoTgK++1VadI=
`protect END_PROTECTED
