`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cWvORfdIZ2xo6OkKeAZ8Jl1ftq+7eikf6ZPYC/B2+oGPrjCw0YYkBpiYnZhNbM2g
PDQXFgGQYiynfvz1sOIFlda8fcdTbaiNyo138dBWAKWnyRIDxOPNIijAeYBmc0IM
/1bKBquoy+aWp+yMP6SlrSuNGEeOs4Xf8Ld+/Zrzz3o2BcTj8w32ulsyHymYz4Cy
N9Z2iJStTPQaw5BOiGcxMb/M96ltMYEPUII5L9Qog0i+fY7ypJS0JM07/f/ZePQp
1oyLpyjcxHzAZev1hEwrN+rvgOP2YJyq7aGfDdM3InnQjdyknzak1VN4H8NGPqOX
asM5zwsq4VJEOkZUoOWjuhkHbgR1g7W8m52SgeC8sYmEvrwqS4wQQYUjMNiM7s9L
Sk9Es1luHhbAS9aGKh3h9d6exN1wj6/IELJdkobTysg5qqh+CEr3+MtH/5H5m/xA
43hmppEKv6froogSrujTdnqfUdishR6R/ERPR4gT3UCOg3tAZPe0bt0mPjpt9N2G
`protect END_PROTECTED
