`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pYVa3G9D1OdaQqjTD+YyELQHdDsRvPmovPaeWvnU0jRsQOKsfMH6YbwpqjA0ouhR
bWad/5llkiWNtzMsrhX9QdHmiI1J4GlYs93FDT4VzeEkWMQqLGOq73Ig0jprBSyD
N5xLktuVuLN8d1wMeeCDWGaId4815JeHxACbPd6y/unZvpv62b5T0OQ4GvS2qnc0
5F45YfpxgU2YWX/yxla/mDS5aSomUN6bYrFLBb85yrp+5kl1HQyvzRFSseiZKiZN
s9MpL1kix+vYmKp35cK8Kmv1RfaLpw0KqFhOsl5TEe2LmI/LCmFmI59CMl6fkn0X
oZp3+C/Pdufgtwf5PtGDe7/P86/dwk8g13Ec4et3fERErouQThQ1zgU8UUQtVp1v
`protect END_PROTECTED
