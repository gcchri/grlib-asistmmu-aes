`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kj4F75dHZzQyjjuIWrDe/8HVa6mx18s0xTF1eCs+v41hS8K7otRNJYYYylw4nT1v
5SJEVMIMCI1cc3omUiz0CZU0UQ4RKWO2+1lUBvUZXW7nkp5Pa+ITI2u1YnJ8bhKM
/bHfEJpIgKrnI8dLbYQU4KmZ8IX2f+cvHDRC6d+4i9e3l48G5VT7hTlwSZ8jK+rD
akuczMX39gT6MD4bbnk/sv0ZIrJMZ1aNPJrgIG2DRoTqW2Arn4bYOclprRbCykIC
Mg0jEtsR4vy6ZYLTVC/SMDAuhrj6q/KOD+Jf5ZeA17hTBR0tsNMlLXxgGZyBdz5q
eH7JIrKUJSWd9mUoDggOxP9h/q4gdqdB2FdqcvOW7fv+1D1TBpeE/GRdNu8SLSM9
ElBi7IOhCbj3CYCXM2xhjYwnAaAzc2Ld1m8VFupN47r7oM967nu3CYj28OAX8/oA
CYdzxqc6I/FPRei3F9ydIj9ryFZVUSbK9L3zzzW5RReM0hxINlRerX0u2Nc9UCwl
I/CQMncM41HVX7DzsAAiD6TEVp8OZMOXpCi2HmhN7GrJgSbB/azwKgo7309OXYRA
/aUvXgik1L8v3JfWP4kFto0dsdSG1bv92FtaLl8wJ/PciiavVWadkD7uQODEAJUn
+INFTg9UsvVaffLxhz+62fdoV2OQAZ8DW/zQTmDcLuSd8VuDfg32/d33bK+/cqGU
rac6+z1bt2xa8VPO9KYE8dcNX3MoZmBEImbtOl8uIrguUDxvjKJxBjJa3Y/gFhaL
aRaYhKc1Cn9uQGOEpP6qxUqL48vlCm0HxiLdacbheNh6iuITI7WVfz99B/p+QZpg
JEY+bjriDf+jIoFr3BDm2308fHffpRLEc/P3Q4qIMD938noP2iUD8ryIawcVF7D3
w1Gtpmu7/WLDSvip1mVA3L4A1Qf/uwhFeycmQASyf0iH1Oo+APPHrpj7ZrT/VW74
TSFMKIlv7+s3Gdvi9ClQDMYl0PBJHP1tIYMyuhi/POLt24jRiHAkiUMmGtgD5HZF
OcWJ7SDDogCLDcSSBYRVtV0Ha7h3AvH5W+dlRM3mJrvi2hWwQkEdF79h1Sgm1Vdo
caYWwHhhMiL79+fAGHqjVedrukrHdQXBx4kwEz2tJbN5fSPq1FHmnODhVRXZwBXs
8m773QzRhJfM12Oe3rxaiTcQJZ+UPpAynzLxlBllilC1HA2xb9ge9z+mOuQkptz9
cXrjYUSY9CGsraMpsax1MlpDFLWujHCxsYbHJ9tZqUDjXo69CCmbFBgK2ITrMETy
f+RJdlwov5PZPyJd6RNAU7dsDj1RLV20FIln0MwkBMK9cNtug+uDuhZGxX0elsdj
+e85MnyLfzXMFfyTVyn/EhZDccEpNcU4TNYmHztxClCX6TCY8H8agpo8p7eEAeug
ENJl1TOjCre/VzGri+L5DcGeZc5gVwTBh9Q6wT5/0fKcqSKkWevCd9Puf9FzML+E
vgSXOTj4E5dW+55O/xXQYVHZbi2zk6UP6kRKuptfZ3svLTJKtbTYpAe0F4vtWKDq
pno5Xm0ZccCBIJkRWzTyTyNHZWwlGDIhDf9B7laKikA0WqZJ+Erlft0k/hvYC97t
8Sxcn1Bxf8akv5amViPlID70QI0SxulH1wKr7qNyTt3kLFBtAcSBxPbNt0uQtdq5
3NhD9dgrjdBPh/o3YnAupCsTKk8yCYvWtfJM9yZ6mRflBPjp3sCeydDsh5Ux7Hez
`protect END_PROTECTED
