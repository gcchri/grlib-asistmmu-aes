`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
61+DLQVf1ylNFZmhULpji8qgYo+PT17DM+62m3U+pI+IT02ttjHHNHdiiJuqCajY
i9BXtUOGsCjlTchg82L+ndsyAN5LglsCC4yta5XgAICLCZy3c+eQG66jqB35+uoJ
5wt8QTpntBxlqmGfwZkZK+VW2qKDkOirjazaDqG2pfaOH7ua191Z3ei+anQ2X6dd
atbEyMqqtutQisOn/UcAD7olqDxfOjRUVaotY7JtFJN0oIf2CMpL8rGHLjIDhGWS
fhNy58v3kJkwMLl/leJHVeoKFJKU2MmflKBTui/U+zOxWBY2W3VHFz10k8BDGPnA
h+gIoV22S7F0fwUdRviOV7bOoOEQpWZazo4cKknOqz9HthSUfFbppbf5x79tWTqD
uYyrWGRYCPPyjTb6RSDtVJqn3CdPQXS3eFWHxavS4fsChSizKoHRGX70lKU5X19c
m/y7ndQKCS26JWKo6DiTXJPl5nYnFSrDk/4ySsr1m287sB8UUe2fjnlxoa0SNlEs
Rs8xqERAZ1JOkNbfQuU0pqYxlbTcjf0+zZfGoK8EcGUrEPQWSErhvK4I8b1evRlJ
`protect END_PROTECTED
