`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NDEefzs2DNzlqAcoTiz3SJsdy+2ASr+joj7kR4m5Eve2/Ud4ZRLGAgAWF1l3W/Xp
MEc1dFAL2QupcR3+eyk/NW4EQwrXLMpB/qeKAhTVSxp2JTzh/qwzY/ZcDCtwrCK3
uA93BKTu7uh7Joi48BIPufEntjqaQh7Y/RwEQKknqaHvM7GKOIOBH8yizPhzFtnQ
9YRaxP2DtccfLFlZOZde0N1JLdgMzhMWa0Bt2uGvH/4TE9CQlQavDTqPq1nX8LZo
4D49UtQ5DA/LxKoeTOaNP6ESqUMhpiWv4qy2/7iusPiflmigkUd6HM4f1QCI6/er
7x94yn42IRCdyxpyf8XZFolO2n7nUpQE6MY0rZ8bSP6YDbmu7GRjrslpcH9ejh2p
Kp2HYax5I+uKXYlbxjZe+FsRGUVONklFYB9dMp8bQ9H7ZWuj3coE11lWzZPShJCq
mHaFEcM0t7NJ3bDOaXZC+ybNSuxhHuD4fJd4T1xL6M3c9jyerkc39Gl+0A3P5DcK
cX2SzRIUJNnmuxAZnzHg9jQYpSxz9nPlSGMsAgDjPCfLyaKRdEkqMkpUEPc40UHu
tcc35UYDLiP2zgQjkxxmL/RFK/S684ItPlVaUFLj+8N+TdA2Wu5D86qJZpi3FRwS
Lgy+/oJeBdqtD2mzSjk6MMVXLUf1m0sFI8BMXuqPrxzuKMl7zlHjQkjsZy0OVXQk
FKwWX0miiLjbcwk+FbCLroTJOco5xFr77JE1jPSY/mmsdZ7pQoyiMQhLH0rAvbWI
`protect END_PROTECTED
