`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jENN4RIZZFz0raNfL9UgKE6MHVIAh5kPXxB6PM+v6N6P/jXHRFUw+FrOZGaYN6Uc
TJwINcHcUaLhl9B1u/o9TNTEq8lfneHk4oj07CKzmJW0L2jMaPjzykZTzVxEaeNu
Dd397C+08l2xeAxS1PJxIN7T5sUzBkERcMSPg9qlIz4nhbJmgL1lNJK5fwQxU+VT
wWffhpoBMgGkkynguhFLFXdXgfTYNzBIea0uwFhEHjWGpEY5GNGVNYFBkL2iWTX5
EhEeSByCi1dazNnCo1gXiw==
`protect END_PROTECTED
