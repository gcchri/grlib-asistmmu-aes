`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4tz6+ZuUBmeFS43Oi9qGMGLnmmepShC3+02bOIXV6YvU1UgcL7VNnxJXnpNQK8xC
mzIAddTAhSxNdlr9iHarrge4dZ0FTjXhAfLupZ3pTekRVB+lpBUzYrkD2gNc+zf/
RHMaQqO6Y5RFdfz6WbsRr8DE0fS9R9m6lyYOYBmGuaJh+65/pN6IZFOeCu37eGXC
u621wRDJvXTugNEeCq5PQdNxKOA0f/1l+Ka3b2jqCHyjm+alNk1jb3K6vKVTLJf+
J3QQ1s99pgFXxEAzWCVRUjRGJ+Xf//4+Ob8PBvA5PAlJl3V/Ua/HDhsxw24+TN5M
+C0eME5t/AhuKNuhsJyDnHTsvFSW5jUcBLJ6WZOfxy/XPjnedpnH1oFX3OL7Gp+i
ZoGaWU/tjbdSc7CD6k5utCg/mU66AaUQm1mzX4nLZNATxBEON/OKwugsZG9wD99c
m8AAgvA9P8NtZkFU0KnxZBjQj1oo7xqRIbl1t8GTNd6Gf3ZrSPSP2+tB13PvLi+T
ARsdgESsbGqDPXCp2wgtzc47KnOT37ww/uyPBmnpve08brPBAdW5l85FMNONq8sU
DuQFZMbf5LkzQ7BJzJE8JZJbg23W2iPMLUeySPFNfQw27hz4g/6cbmLNz+tAyQr6
zchREpmShZX2bWrISv0ecqRnul0y3JXFnu+O/2natd7uocVTRLH11Hc4r1D5aSQm
q55BIGRtE6daMDU7QF40cM21lCiGuykV3d4Gigo1K7AWcsd0U9W2K0Te4XCkVtp3
YRXj653ScttTOu7bo64N8Qs76SlMpED1hu6iy6vAUy8pBlMwJeEYcRJ068a86wWL
h+y2ZNwAeZnvpZWEsS1h73pSzS+QrOk5powFI46hCPnz2ehFxhL/FIZmZ76Q7vOP
feRzWmkr+hwsq4BWuSg5ThakQRpmxsaR3Ov2RZZZzSl5xlnkPJSqmfAdp1HFCg+V
SsyVRxOlcvpY87PlcbXrAbH/XsRYkOZCQlUw4AoQi2I2fBkOaGQ4bhgQdRPzVXSz
BMW9b8hRuOIeA3SFMjff/coQEBtRETsOKT2Cot9ynApGd1dU3bWSBuq+97pz0Gio
KVKpGsESFsPP89VqTmB/ts0d6WIgDXV+yUNPJJg7DkcIDl2VLJXHNXsCm5W880PA
AUxGKDQpmuvDlGySge+F/vPQaazvCyicnKUifPJ/RbGyPp7+3WEs/d/np71xe8Ws
2w3Hrws2eZnSzjpLTR8Wf8d5qmuRNl64tSul9izdp91J0Lf5DN5qdLDKPRz2hMPg
kR8jnQfBCnXdWZwMe1aHCPGALGwm60z3CpOHVdZmX60OGyeLc7X8XHO+hxkypeIz
QaV50zA80RYhQP4o1bWF+/Q6K0MM/4vXIZlCm6Y+LNZ15o2jxkfQOOCIdryXzjyq
UBcOFUdBx59DSVy0L3h7Vga3h2WRv6G8Wn6L7LHDyiE8pgQLsrTIvpmG7DJU8Ggm
hMdAXOwKkuqo52xB4IOYnk/i6uDPTuJx9cG9GxUSgn/upl2bgSwh/+PVyGzDiXVG
u6CpNif9wwnkbq5Yyj6a3LxKpKNAWzuNH3MJznHn7MNDFADm7RuhQVjShSdHH26+
/k3hjgBQdv+HO9d2Eg11RcxifxS//GrXiuotjYbym8bqGYxj+OFj4Sk+mu00Rk7C
j34BgAPNBfk51/lTpGTBu9nzVaVGWcsXLX3X2Imj7ovdQWRenigv8kIg4dbE6nQC
fHS6KSENPr9MnNqx3pnjcn6PLnjmf13CaJ43UnEZrU85TaS4OJdKE5AkTt0jS3y3
h5GKKzc+6VTcGJhGRM0rvXSvqnsztKinr2jj22Cqlj3jhh5f9p7I/QFBVhj4l6Ci
`protect END_PROTECTED
