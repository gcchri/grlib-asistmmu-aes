`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ymROQPjEJmmD52Rqo5qiewcegJ1M4qAyRfuq5N5ZmXJGMzn/TwRKwz+QrRn8wH5z
6uMc7lok+KSkU1ZJlXU+pfVAVLXvVNoFExAue0uA7/FdvoxP4HMxtfwrr2dV39j4
2N4kaZc729WJYdZ3ENzqYlWn++NPrLD9tBgGATEmY4uCNv+z1nfxnz8CZzGayxM8
dp46kDLhyHpm1CZLNGoSx0HP5CFUpFIpww+GM2fytLJ8u2Y9KgDCosDw3MPNQpJV
hJtNYrRsU1BTgt1L98obv2oHj6aECKWw3NR+qxoq9yY=
`protect END_PROTECTED
