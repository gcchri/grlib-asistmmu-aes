`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rRv+oxKsox6OdfZnBRlUBPleIDXa7HlchYtXo+ULSntD1jVjs7qEK84JD8sqSXkr
7Tw//4QRkTnDikpRGClcOIGkvc7KmO0hHR6UsjqUhSpzH1u8IVSD3a0+DwHrMKJk
/hEugYmmash0xE6rd3uZjiI4F7/Y52Sp+HKWgcVEsyobH4kELMpivYnNVD4qWLK1
3sokWKbjqrgmOJuDkUQ+TiPYgG7HN80eSexqj7QQ842w4UNYtxKlRL3TyfINZRpY
fM2e9PdBOAkNeRRbuWnlaSfNdPTKU/cLuHnvfQrP+akDgYDQ9NCslhV0OHUzjL2Z
kuo1QAu+B11/8AVc6jA5XZbDhqUxymurX9UT4NoMMIaAvMAbvU99aBS3aPtl6yAh
llWHsDLagTMkTdihzcMHa4L+ReusxpZ40Wzes2hrcJvJ1q3IPZh7X9mC9rsS6f0e
WF5pOSYYMVn60usEK/hJInfwGykInEWHhvxr3e7lavfR77RnIQHAivnJavOr7nN6
tCnrERF9cnezCeLaXUMrafm/mJR6csz+fkOoCkaECnw6upjZjYYFru+0bQIH3Vqj
B5DH+X3Nf8yvVyvdvr3UPyPHNdZcjHR3osX9lT2jcJQSWGrU6OEH6oUtFgCpVu0r
x5AcMzjgNE7soRi+oUBYTuZjDx44AvNYRC5OXbbIGbotOeK/prqDHC+BDT3cN81F
ShuQ6O89GbzJo/kFgzcUY6cuR46RDC9RqYCZ4lhITHY=
`protect END_PROTECTED
