`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bnfw+a8yYapJiO0KuFET5ZU4bwhhqrz2EbMOkzyNIJXWabDhT8UkZ+NgeXdF5B+8
vz5xpb1YPeKTO7K8D97Joxc1d0mo/ToH1l2SthMD9pDE3yqZIJp6eulf1LWczl5n
zGIQ1nCG9HL4UajQXCkqz+zidY5R3AWA6Zc48YiLP9k4bwXLE1Kaxkf8JtXXs9oU
WMoy4duUmszA6W5prwMAZcwIfKsGckxlx4ozfWUUBzUBcFcEc9bBwtkPiQ+T/HgX
iEi2FMZ9EmHG2xQ429cwcvTX6C0p8vICIMW+2e/UBcdbgYleyFqxm3A0tkTjSteq
`protect END_PROTECTED
