`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
urnzVUE8Sqy5ubGTWW9lGtqzEDjFDAo+31wmf+N/EevErvsKqpfPBrKT31XO+JG7
4jOOlaiXSySSpi7vz67KjvPgm5XMKQ3HJSCUmuO0ayh8Y5unGL6xUSa092D09hUa
0ojgjfhX9OcM7H9GScNbR+LtBBs1MO8qZZoKwxe/bP18/DuUowP8vwTEZQrfZC6H
i768q47FMyz/a0HP1myjpiDFiFc501RMpqnguwpv4vFUD/Q3K4BbwDNwihJE5elJ
EqkcNn4RdeZAfSyIP0vuG+MzHEyEBQoXlH3XbJs+botmZ5GLDq9jSJZ9st3QCK3K
Z4kHLe2vQK9g/R/rBQOFPn5smVsprkrS0eK9Ay7OFv+d2aEK3D7iEC1h65qfZWQ2
vjuVuSoavHKDgYn8y1ku4R1oi60jVA0uz+6lnP2n3VY7pvth+UgODK/trWYjx0vO
i828CCGwRuCxGxpD31b40DJAXbPFPOK8Pw3MlUsdHJjVtemnRHMRi3rrER6x2rNm
Rxa5YP+HAtu3jbma4yvH5Wt8yf6a6nz6rI63FspVkf3QNqaaZXU3TYGNFmrqXzBW
tC2YC6j3efYNME8tYzadqGW+Y6VKh8VJk2Zxj63IAa8=
`protect END_PROTECTED
