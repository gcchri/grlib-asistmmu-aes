`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tbLGEFZUMQTUE30sVTFzVTmshBxrFfdllJgqLqJTiwvkXP9/MrCDjZA8eLwJ/vCB
+MwRNMW65EHA4sgqq2TyUNAkGQvgT8QN934LOuLZqmZhIU+qz1nkW6yxRVwWg+pM
JQ5Rz+O8Dq05nTDRTww3C8Ww+SMFrehKKBlGUjnIWsuSdgDcTk8flyo6cQ1deMOF
0QD/4DV/oMEFHvGnto87GFtmE2KmZneIKlEvKCqEclZV9SJtf96P+9m0kvN+IGzC
WWGIjHWKvWTYhDElEWZqKes7ZZiVmSuwzOVUn76mSs3v72r9/0xWRKT7CwFEIvMz
mENIbftXbqfA0dovAHBSIwUjLFTtJT7QuQFlGrtIF3RR49cNSVWv6+NTnTiluy9y
/55shWTFdPC+sDfz/DKdirfNyBGNLHuyl/a2y730bpFYu3RkTBqsOLp/4Rik0Ulq
LhOOI/uCG+w/IUwSvfxH4g==
`protect END_PROTECTED
