`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i1iKz+PU7FgCdh3CL6RVYbsS7aDzl8vutHURabYleTOWRZRvqvkAOVVWgxIeXbZm
oYnz5/bqEftP3STeGlhWoErVfOr93CvItsjHxwwiVFJdBFL6ecvSI+lUNqaOMRuq
cQv7h3IMSGOBk/KBq3sCIjDrhkRuG9H23+kPXO+DmoQDHRMQtkQJJR8bG70Xm2bV
y2oqNGPzltX06yyT563lN1SBsqIiytw/lHgVe9ikfzLklKDkOZEzqK87cw2dfL/m
f0OtqPNmjyDsDAgI3tjxrSUBepzYK4h16ONRFdPS0AdaaRVhLckAro3UIEL+6Efm
3OmKue/F0JPftrmARC3+2Sr3NgidpRJnlykQ0MwTZz9svV0upj1ZmoXtMHcuv/4V
nyBcAShf/ItHb+KFuvQkDPcso6V5fQSVWs6Jl+igmvAYG/ZAwEL8DZu/qqNRHLH+
KNJemIL7cGcpAiPvi5rMfrn7zArwjuUOzzcgZ6MtK6Jfp5yUfPVtS+bdFYGY1snv
rq485rI0UXr3YdWbzinOY/mvtEI3iQ6dGFLEKRqBkbA1Zp7E42cg0fmkvqbU4J95
KVoPEL4lRWFpQmJEnyzoczYI4SzmVtCy8uBaQLhLF89wUyEUGy76ofEhHW2fep3L
79ESEtiRSEmOAYHwbwzgRebZBCosT7AE6wjUS2P2OQgo3lm5zSuDSgmJ9N0ckO5A
/8YZIkWGq6t2L9qcz4/9/w==
`protect END_PROTECTED
