`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wmvjpHN7YxNmWPbsWkx0rJtNpzQLXBnNMeOh/57i2E0WYy5hNc9wPdhX55ZUxcxn
WSUHyz0KkslOyr1+Ih5kKmtS66aBM5ya6dtNm0aHh6TQoegayHFzDWgMQTxX7YKR
+kmhAErPrZ7GmMgf9BrGQLlv85I0nk7wxXQA8gRhfPYtXD4fmd+fkyw1avxVzSkB
AJFaPAJgJePz62KjARwAP//LUjPH25QFCB2WSWkA1F2mTjHt8VarMbx/tiJ9d/jY
fz1w/8w9tAF/UzVauRd9nUaXXHXp0G1vYa7uQyDfWPN1M7ZMj790byuBtFT3jzZJ
BqltcDQ5nlzekWVovOZqgRtMYThJWm9bBpnJRTfkM2lvuXdehEettkwC1GSZAMAi
PN42cWG4K1lchIWH/8mZJWVwS6nf4HM3Gwh9xBTJu2XV4zFrxeM8f+LtGfh1n+sY
I1riQrMTcvoqSEcsFf8mdfK4Ckl2zVYRGIrFGDE5sqKVx+43AAlaKRN+ew7DweHv
ulP//iOqr+Awpr8SV8tZq339FujoVwSdyJu/D+cKUdkaGVlb6GyxpZULgPTwMsC4
iUEzgxFjuFc6pFUGEJc803czYFoaDpiVdfL2Zo51gWrroI7sfPh9MI3klM5ce539
adJlTZqyBltvyQgCh1x4B4xYOkzbn4YFmA5kanQ5R7ks5e+sBvn4ePgBW/7+gP9l
0fEtyU5kQgnf8sBzLXfJlB32KIvEHHmP55zJzHubpVsZMxI5hcvdnkILgcrfGFWV
EDMNyXvl/neqaOR1ky4OlfHYJ+GfXrGIwJT7O4POk/+3AUlK1UOVWrq2iv0ttsEr
ntM6XWflPppQMWkvJkuXWKSa0w3umYwqCsKCuIzw07CMqAlMff/vBlL5eXzO0IDk
ZuWHEzSuhuqebZsxbcUOEhhFO9cqTBk7ClaYkrv9O/uUkiPhRjxdx1gNL6WDW4Pc
3Dlxjeo8QNCaLvVH/cpsgQhM7o+ttQgn6mR9HA7a7+Bv5tWJL7tYvBOjw06LaMk4
8ExIOFV6bWz+WHUQZ+tH/bV9jfPmjBZmyzCk98hu4RoZ9twjAGwQDn3EojBmxFWs
Tf/WSN5m/tArlsJ45Er5Ebwc+6bWYg+wRZP4792chREP2k74avQMGzJeAWJDCqW8
LzMrZvaOmKdQj49XDDTBe13UEPBNXkjQXBJ+RIht1E9pgPL12SgD+CfbaXI87NaS
f1ot2DEZugeEP9pGGv0cCTCRdPPm1qJRItzkBtGGa+Q9NdxWUL5DRtLIcDSHdsTd
auShtHZQ2SbiHBwzxePUXNb+ymXMv5500M5mIAuKHiBd433iZtfrRYHopMpgkWbO
7fCApJGaDKoKWGpTMum+kDxY+mnrOEeJlpvON0gYtg2LoADFRVgwZN9RteX7HKCr
ESv5iLT7osT35Zp9bqEax/J4Ijdj4PwwmwmTbVO60ouvYgQYzm66v7LhtxHTxxAg
cLKvHN17afuUboZ5TZFvb3ZDhkIrfI9p6TQd6Whglgl4Et7GKKyls1mAZ+fFjYsx
s6EZATK263gOKQf4QXQQoYqsojmOR3htOUigG+89cP31SR/+BuI/QtmTK18TRNdq
oKOoZx9SwtICGn6RSNzcR7aDy1y3n2jdB5lU6fOStTV9a0cx9npjE+eFLwtuSObj
iWLw9GPNwj0qwNEc+MtUEU6meUHhAHriuleLYzFtYrzc+qx3G9CBtabwRSxdu3TU
R4yZUJMf8tEXL470HXR3DC0AOWZW/UVzE5ddnrG7xPSdepvejQkFy16DVPLuwWoB
Pz6Q0bdjAk2NFiGxvm1UDc9HfMrfCRT+5jWPe5stMfeje3t5THWg8neKh+OMzE5T
x4O8TFck7WEqzWclvy18dUrvwBPIC3RYvVxFUckd+CowU1wLmz/PyqpogcAD7xS1
j8cJGqTFXhU1O22wEugm09WbaMO9MOry7o4AS1e4VXQYa+8tO5NDoeu9W/Aets+m
Gn9l8RFHKGHRVxrA+bDaJo5QRNqqiGD0yaO/+rFgU6KMjGEIHZqyMi2ngvrt52vU
YG3UVh8indh8N0nxnBub2YlLAmsUEhV3C5yDcZpwsRr9Jix9I5TfZ91PHR2KUspO
O0vEyJUTSPaYv9PcsqcZFoXLZsfBhXg/Ql1/7h/q9rHLxWWzkvqzdyI3wLw/BlEF
d6/oM/COv+BULSLXt1NfREaTfmUogWBucXGRJgA1A351zA8JJqNX7hFdV2sFkEcn
++tMq7kEIXtJRuFjDASByWwLx0y9uEBceUvH9DD35U6xgCnsTp9RpLMFDviyL6B/
Ytlp/jFpLk1xAqhMjqXAZ9XV0ORayN+3r2L+SMkgZXMsWG6A5MAxm+vxSF3guKee
q+3dSVqcaQ0sBN9S71CBGQPgJA9ub7/xnNL3pwR1xnl3pJoDiLstv3vDpNzIUEWm
QEaJ1dvsgOZ/DSG9y6rmNv/rRxs74csC1xbNwh92LC4ema8fVyYjYVzhj5tou3RS
uB0aGD5Y6U0DBknj+wvUCykwUAWAGVnM0FbqS4KkDJ3HboOy7882QH6enJ6d0D35
rUYmABhLzXkjFFTNccE1QNpGO08QmSiBcrDB8dlpgXcWCPVAFKhJAXvx1kNjG5rN
d0YenETuo3DE4RvwxyD2PgeFkDRpkzq3jswbKXruN1GgkB3v/k7QXkzt6zSvBkRl
Xj4AQ93xAWdglIOD3G3acO5HvAg4UXMPOCkrvAsRnBpJhG6jnUjM5oFVFARkp4MR
/U1eGWiq2uIpZ1yPAbkmXsOF+GDoAggatzXktM/wiNeeJlNrw8Q5OVdLxFyQtyUg
68DtIn+woT/BC1r0PynxJMinQpGv3XR/8X3pFhKz1kOaNtc01nnidW43RLpy8PmA
clXxDBSWWCSjJNXj/UXHdACshXwZdaZGNNj4kfsU81lH+u2WMbg4+hwG24nhGzDj
apObfOcPQ2SKSzB8IJA6rvB5Pe7GDDGVb9SBdz68xFnTkP+ylpAJX48RYIH60daV
4nDO3cnQdY3cZysUNA6bny4qjppCBqVTeBmexmFHocoqLonP7IpQDVJ7/tJ/YDBP
80Hj25KlnpnwXMCMYDMYB7oxTUmBh3T0g7APvj4S6EDrqrLkfeJ5ivDNg8LBk4Is
HyNYODe2KVrJK+sEVccl/q9VHWiCNf6c/FPzOF8dReTSFgINMhHA+DiZf6Hqwo67
4P60EE3PWjN7Tga1a7XjKKOodSd9x9RUCqujFfVnCtZsPo4nmFLxenIs7PEJ7vL5
9IJ/Ck3AvKOGsoKlxtiPZxvUmeCY3QF0EbGqf/lrad9pVAdCEqwC2Nd2+7CBarw3
5T5qP9iq2qb3hzjFHoW44vAaLOf3+L8w0ZhCUz1YHaXEevQEN4/ji0YBpxCs4zyD
UsxIwsaXkEi9OG+FQ9UPYaoJu4W7lVBKe6RWe+g8TGZPyY6NoUUHNlb2b7bgSwNI
x3l+NFsxFGUSeRf+hiupeTlW46BMqnZg7oP/61uN82jLAmVKCSpvki4sI/CnBacj
FaMXw9ekxbEjJ8KVN2ZTPZATH3656E1pVJT51NBT3daAOUlYbgg1DWNPqDkwNWV4
FyBjWtoNCWZyIitFFcEz8SDA6R+Oqo4diFWsjkqaQsX0BQ/t+TyKEwcA+zgavmdJ
HYdsACEZNDS2D+b3TYRvXn3VwHpFKgmpYZyKAI9qjEZ/0XcurFVt8S9L/i/9nUNc
beeyybBXD96vywR9Gsk1y6z3mkciPGS1XYDSepNsVjz0zMK8srsgSWzEwtzjc4ic
uD62hZuGYDaLD+cCa5Lbos9QItTsCG/RXruXGB28VO8I+A9QNo1SASryUButhtyw
CJN6obY6z1VFpmbcKpSiNfU/XI5/GajH81DoEQsp4VWmfjUamvNXqU4YbbrlUtIS
yPKnxSDB21ZGlo21BeVV8c3ixfCQG5HAP19HrN4u6EGtxSortAjisYecsPsFo2m9
ZNZ5ah589a/4Z9H2Tnd37TtksQ8Ml3tKQ9lQOpv+/QVLg2G9BejO0Ir/ih3CkBum
0ZorGMkY55RuFfmumpy7UD/wKKwGPrr3TUo/5q05R/Xm8YJEu0NEybW4jNdlAVvg
3tELI34tdiB51d7a+EI3HA9q7uhkyj16uPTcb+eOUs2udyv2Sgpl9GPNujlCH73P
qwONArib636zlQeCImNAXTXFzF5AY3tz/ocgCelFjXvO4rhF5hfPFEABvwSjfsRW
hFaxvA5r2ZpaM4RVyf2BecQo4NLbyFoCjEmu2LHs0RB/3He6FPwGcClt/Gk/giHO
afxB8wMKX1IGLIcD2qpcjQHQ2Fl/wQnA9IqJTPcZrx1CMCFIbPL5s4s43k7BCyXT
MsdLgwiZEI8gH+4LZHUUZJTx+FwgcrttaFQZYKhC3VUDw9eMYeAAJhb44TELFLvu
GvdNMkGkcnVALiFmmbomLHzRehdFeDkpjD2m2aVakZzHemg6AYl7QZmDddDTPlak
hxSwGh/4u2fnKGzonN0q4Bb7Nm6QMsEZJIHZK5xPTtzgPnN1zkJT1OJg7g6qv3jf
pudDIiAqzwDoSzXFiK0dyMuVX0QeerFoMnXhopMuE7o=
`protect END_PROTECTED
