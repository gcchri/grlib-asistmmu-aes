`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kqgNoa58KEJGRqsofNktiNq74E+Wjgcr78IuouB3+mVJoXGM8rHqOSPQCQFBx+09
FsoQDwsQpAU6Q28wxPzKSxq5YO2W+oPKKtLFPocOD2AwSwUyY3wZwAI/iAYoyh45
p2NaQG9hd5BnBwhU2SjtP9Eomr70oVR9JB0z6A35+yfSxrgJEetvyOwd8/cAo6US
cL2aA3b/8pfe45KZC/GRFXXdVOUL7J9EnYuF2bZcsOkMmGmVp3lzp3IuVuqeQ+PN
sd9DQv9DisKkaTLGDacTCPfon6sC0R6505Rr7oL+aMUSqsJp+hlov8kIVnXgFYcW
MH9rHoiNCFkn3mi5K8jPdmNek8utr/dUeWY2TpD+Ci6JwQ9yotw0KHecimVdrIiE
aSbxac7ZNtSTIiglsrbGkzJVDBxoaTpnXx5mYK5w9seyjRTQ3Uej6LrQYb0k589T
MFzgvK3tsPARj0PR4tYQM47Y0nDr8Njg2bOJEoZdd3MLPz8s6LDoTeJbiTqWObm3
5Kc+VbbOUMDQGim6HmafpbxRVX6jSbA8/SkK2SgbMExczwWYJZYZVXUgrjFkI2OQ
i/VEVMmv6HvPXiMhrDijdUEjyFKNMM2PXUM4NzHpYb+jSsnIugQT58LEDEUZBz/2
F2fzXUvyYny4ZGuDnjJPhdtgYEDHvhVmWn94lSYn7lOKfsGPo3kZohGzxF6V2Qxu
HbzIwPjxaSPTR4uJ2WCDzFOH4xOOXMFq8MA2Wgdx4CNeFyVkaUkWYmvk2poW4mrm
PdCDuAN/ViQNv63K6L/udguVZlFPM8jNORZu+HRuBKd8CXkOv1RfJkt2KzgPBoMt
706JVdr9MTl5ElLME9f1b+QeYYIwVo2QDBvnZ+tIn6FTb1sWQHS80IalVyQhh8u7
gjNQALwO1u8YpIlm3alZwCgy1ZvLY69BS3AHYKYKKdZHAnxYumgphfxr5KJDeh4J
PoYUFEntCT7cl8o7XRlVH75qA6PrsF4mkUC+CkgqFWO2a66rz1LSrEnMnCkRV4SW
vKE+agqMbf5HF9kB7lGQWtvzFdfI4vp9+eLJIAstzfVQvskTrRFy1AHD4ocTfMv3
TN0+qZSoxLfiaokgrwodgSl0MPIjvScyXRkyFOdxauADedcUNz2KaBv5DLPkXV5D
tVI3R+Gt9TKXpctEmYQUzSpJjgLOxKFCemvAP8d1IRXccRXlReqYrBgh+5OmxnKg
ONI1KUqVC71d8IcxwKS71maNuPIgKPx0Vrar8y2Yl405luR/d2FOV5T/wYfabRQt
lDVxtu2IDzA+HilvAflfHMj/yLn0zJCT1daUcExfV1bhQE5hK3MBmsap9ap9F7WY
wWuuuDbOF1UlGo1f2Kd36LaJQ7BofOQ/5RLv7zS0rBt/0Qtbuvi7aRVmnMDrydHT
+/cSbGVHMopCuFpU0jAuouThX2iyatL69Mg8bVOEu3yorNa5UqWUkWzmtYD+hW3/
EZdVV+qgWsmiRR8IxEkaNwYRKyRyy203ldg29fhDIl3btvfAiQJej3Gpj3GUiX/Y
kCpwu/27/tjMdHY3f/Shg9ccIw90cDkbyVpazmFqav7x379Br3ATePN4fT/mxELG
2JS0uwTUZ3rT20kwYSfiUC/8J7FZa7Ma/4rvwVuOQ7ESXkXJf8we2e1vL0zN5dlJ
rQeaIt+C+5CFG9tdWpvUEyX0U0R/AYckJRfm5GMvazdbbh1W9x5hz4IWyKaAwOnZ
yp/kY2rAWrFWClmj5W1f99j9Hgu3S6xWJhlu2GXMpw5axz5rZGL3B+o9ARm+UVoi
dBZMxUcMfa8jb4DEZsyjGgXhun3x0z/LpNKi9S7P5NAGYXHFTV+zObXwrF1wUdsa
Xxmq2SYSZ/1ImavcTWXM5ICBNF9x40uimQdtMrn8CxjY6VRC095zPVioRO8ImUdF
50e8hvBht3O9Dnxsys86KtQpmGoOOJTeAinkU7Q8ksZHMvADBNYpkinwGqU34o5p
JJMQsnRDvHYROIVRUr48k7g52O6aSFp49l9fTk4wgwGLXW0M6hRcvotr4AWYzBuf
ROnbY1+U/JaOrxDVLqeF8E5STmBUxx6GRUpV+ynWaYZUMfnGHW1gelBnU/gsg8m9
k/9rp1ANcNxyC2ob4EboXzueMkC5SKjHTf/MEpPd3nsWMgDxpJggTm/EvcsPzn/Q
tLFyRulcQOd3pxv5JArnVvSWa30nQueKZSdQPd3ViUtLVY0g9X7re2gWZlGT7fcI
Q7eTOLPdsWuOSSkO0rpfx122aiduUptB7ScmKyBTLTVtp7Rf+H7tG8zDPWICfFhK
Oz3g54ytv35wzUwF1H4g3vlrKuBgL+rSDEN3JuuuQYjIx1O0lltY5A3tLf418FAD
oyoUnt0uQMc4jRorW+iON54wQ97/Pc56DA0nn1C3i+7G59ZgTweCuROYaW/5o5wq
A9gDcxucfuvsVl5/Fz+eupdox43YT5Ncayd+IJvf/GzE5J6bU4ybqPtg0JDK8B/Q
UCeh6F3sc6vt0LLHVCpH2gI9uzP7JvoUos5q5haR6B3fBIoyS2fx9nk5m6lYzA2w
VzuFI4f9DZxKfTWQc6BObEwGvSrd/8Mm+SOBjgh8PnHtxzb0Sm2x0HKrKOmt33ej
oXkm8hunu+2vkzY8Bw68rDJbRNHOcGvj2XSHu65ACwvUa7lOXBoGWNDBy9n0pkwE
DjjJ9dapDZPlGhkgKCTjg/TwUkxxEnFHOVbCtZLskjxpqKartJckl18Wqqzlt5eK
nW0mXO2s9Jezg3Uu0fHeZI6yYeaeRpTf73f6WtFXGo058Wj+r0+5n7vN2fkeOiXr
G+vKV3ukwXn6FzY5fczKY3apRGNZ7ywDmsC93h2XwGOKyE/oB3JAQr07UZYEwsKN
Z4+LW9PaxQTPXqDxW4erNrQaVe6QTHq7w785wBz7imAn2ziDTQyWVVCHaOCBu8Dy
Wf0Z5J/53r7Nh0hGWADO3Xgzl9/jgj4CjiGGOfRaJ5ursot0ggNHi8i9erZwDsL8
AwJzMTY05KAfUyp9L2rqKNhOXYlJbcsWsXrSf0DlPX3wI3SLuXD+/e7RyhMkwuWJ
KrWyzZRhLf1Vg1CrTBwmB8muwtCSpg/+i7n/FyxkJP4AR86ismjLRqGBO/xvQ7kh
31qPZhDsJCYULREyJg95+2DsvPg4pshYIFWsHEHfoCCy1Bu5c7b57eq/QOL51Xwn
7ecCMJryRosovv3EsTSDqjV171aZ2tJwRBX06eGxaksK8WUBxWU08joG4AKg79y1
+81SPmBR+5koNyxELpb6zLi95ROV1SIizOgj4JQvRmZ+Wa8ulOH6cVrTFYUjvI6T
HGY0h04q2k64dc5+/OQZ1pXu04Zfm07s9XUqeIxKs0PXy/2h+C+3RaBmQa3Yf3iX
sp+C1mR8/ZFJeCenBY6GwAaQcWojWDquCKDD73QtpECuNhTAGsXrL6XT0rICGwW1
CCX/DN53ZuW2xp0gB1sHgJQ7Y0s51Tek8+PRep+X0HBmvCxpOTtO9r5hJmrgTPBm
JIYRC4mAbVYCZNwX78wpTKtgXRsq3jqkfJ9e+e0GRdXq/Pdsrai2hocdYzn/laDv
0JL5ePy3VGRuk4Cqcq/NBLtZ3TmDUQaGd0YtBkqFJaO4B1DZyAGPTL8IdT+Bc8HX
dnLuY5N2ArKYRJ2vWmzTUAqnztn/51LeQx2EBzXYo91GHUeuh6FHYNgVjDDv6qUl
33sE4gVlXem24u4DgKV3pE8KDEkIpqo+P60Q88Zxq3AUZjDXjvx6MytdeM05CYN6
o2AxFmkrOp2+SUFvdeAYMo0uu5x0WMo5qK4IdwnOiRhQwr5z/Gl/qa9EwSbjfFa/
bvd4NpBqc49QapP7Vb4qZB0XgIWsTjZ4Hf/Z1e81wKGkcnmGDmRTF/hIHCplC72l
9ouorLpp3HUU7Hi3ahj0Vr8Ux/uJcXsyjEKW0z2njdvTwtBGxcixX7Lijk0zR4R5
oDI8iZIU9yTQglNpamz0cOxzYShmyrRZz83nCXtrH9jduMeFCdn0+NwPT+FsZPi9
/+n+IjPsYW0z7GPcXc0OfMmLjMesQb8FVNEj2IY/CqOTcgmwM5B8jxdGS8Fl3xIW
Yzhj8aGh6aSWi9tWVnzC4oWP9V5tQM8bbJLfl4f4j79dAysaU49h9jX1EsKz0zan
aQAvcoh7dzB31C4FstDUXYTeNEharKrXUwZmCE6RW9RcRucmhfvU6A4pL+5oTC9p
1gzEpWp3Gx09rv3WL61w0iB0L9KEZKYWtF0tjxlam8BZKbNhbBYZf04cKr2jaisI
Izhcw14LFcpiJ0SZtq0tP4fslb3TAGKxB9We30iE0SKXZOf/CDf3SxssggWsIXbd
5HSWsUvBg2FzDIIgrGDL1ZYvqA160zdxKL9ZTeJQ8OxJjWlFaHm3Far7ZAAFsQxV
yGytyJHlsMcSCI1z4GF1fXjvOVoseGZRYqPENCAebCeWIPOC1+PGFAIZAlOnmcOj
T3Yk43o0r5Bd9jOp2FhqnavCr4nOjeA4R8jYZW9achIqCFSar3rkbnzIOCi33p8D
nTexOBsbnAmIzZce9aNP7xXdw4c+XddL9PgWg1yC+WeuM4X7ratF6VNkWwVBtb6g
7GJgOd/ouLWJ0YSMbaxB2ZLkFSce8P3vVB8BzEwg+LL9rU23XvzgGWbTZvCmgNaZ
EVdkTwHwW/N3qMKzN1VTd7IHcK5z5qirL0KYzp8ph+MjgUTrlZKx9beymoRrifd/
qnLXDkUvVY4RimtziPGPP5a+9WlaCgi9FjnKN+FWNkAi720W25aN0rJQJuKAGtZA
fbL7bySQJ4QpwmiE5UMttICjE7uYZW/7zgOlmR29Y5Z/N2e500RNdcmHiU0VUpV6
XiMhmQxLcSZoguEk47TXSRfLQn9mR85wu/9UfKwueSQcoqmoobUpKlx6nkHOyn6i
9ZWgoNK+leI6krNUPuii65nSJLshtkupelMizA+/XZ2821jD+W2fFdRt0S9BTNOj
02Vevxnn5Zi6NBbBdWeJlsuNCxnYdux4lhQ2/3LEfTpxoklrGJauL7jdIt48OQ/D
zDwMas4OEq+QnUe1LESrB9s+6JxHP5uJu2vEDGgR6H2mCWQQ9saZtMUlNfrwbsrO
j5EeFJfaiqMletzdyHAEVTuUQG2YMI6IMj4wfe4040r4+3cplAsexwTynh3XZQa0
NcQfHi+rykmnUET+rx1lWpTb5RKWl3u2jg/FDGnJIdpn+3emsAfKU5bc5rcz9vAH
3mtQl/BcdLGTjQXKcFBAq31M2Ah4tIjPTXRLCRTlCPy8R76o2KiGG8BAJ8Cdb5qy
MKaYeSSt2Gbcg9bCJLdzAutb+OF7P/prSHL6yv9mynp7iMOeNEeSCWb5ejRjlw9B
6izMM0c5ilRcD0AYwGWhn0RICfmdGW/rXDN6JWrQfTi5IJdXDwuGJe1B33W6Dxr3
2OEfjS0AOPFMzGlIdsls+beTEATy0BRO3UxfyckmhMuvNRyNxXk0FA/hUxN7KbMG
PGcDNn2VJa+JESRBP/JP8w2XLTKy1vhQPJAlwPp9s+xgV3sNqZbL/3E+byNX71R9
NCcEihA3R/NsoIvByS7QvlCZNLr7X4sYHKeipmcqTct29mHVX0esFuyathicpoou
syQKdDpMpnqWg0B9K/45+F4u1yswCfBdi6BsdwTavASk8SlrV4uPdlwsOUyZldHW
6pP0d+ps87FFj3MwEvJCe5vFcB2x3yDO+Y6kCCBh73uld3N5Xs9mEM2YyyIUKWeN
d+JVfU06DphR15n51dxEo3HwqoNSx0gD9l7w1ESyrmhXjff/b/2J9Q89Mr032g9h
Qjxwt5VCEQjUHwmjdBjUPtc0aFDgUx+JbPoCK+UqikysgmAD9t2C70+65qdQc1Ze
10fG7bzWLp0+wvTKOGEajIm9VidajukNsM8OSYnZ6PuKFBcWvKUZvusFgykHugeT
pD17/8QbXaD8yxiI0wdQz6KTDHjc3VGlm8QkWbi3P5meEyGWSNIisj1dMTj6W8dI
aGV6yPumKkMdnr3xXJrXV3n2dleI+oa57Ejz+0tsEiXMFJ7JyVLTvQu/SP6vKHln
Yk9fNbP+IeUyUDD//1CALHwCIJG6tZtiM5SJPp8nA/kNtrIAdztFOWP+yEMEUZnJ
+wq4ZQ2SXsaJpjqNvk+nQz+O5UmjCyfYehGXQAmTiJYJvcURnnHZ1gAWGx8O3pHq
04/ZUlT/62XamHWqozXe41AHb0Fy51P7W/xxQMiSQ9AmzslHkrLLErFblic5UAuc
yPwCAqx5E9eqQ6XyQtVZPF/kKeig/ARj9VXUAAyd22BJq0ITMWRs6ER5COAbAasL
rp8+m119nR55v8Egaq5u6hDLS7DC+WaRjBuF/PlzHpdS6g0FB4RRQAH9xJ5LhTBq
FOXH2U6YBSlZtU6E+qcTOodnvHeaRAFcy0LC0lmsGFKGgMK392fcHDhKUuUMCMoD
w4HPpRm8E9CTLsYvIwK3zsRbSjRniWcWnmdNJUH6K5yxnuG9sBKDMH11w+AXaNcX
Vsb3mGuIKWyZrNJByOBlGxB2JYwK84Hllbh+VfSsO79NbZtKmdKc7v4KvY87Zatf
U5QvsW5RdZnfIdv6oowJLtLZKFDvIKEal8YxgEabCzgJKyapf9JQsDrEFR3Ejemn
2qRwdT/AXIIIsvmtbIYMa8BvdPAbVmvn7bEr3ynuEnOqEh20NngiEgpVmuIqpJlD
x6Pox97c8cID7AjQgYyE8ltcNeJVUnTW4v6RLBaRuiuzTXDMQepQzwNfWxXDkrvg
Mrr1e+FtXMqQ/W++7js39mL4bc6prMdNDBS5r/LLQcKsCR/nFa6PQfCgSEm5DvLp
y9gBm+YGUEgtgbxlPSxSGT46pMz/rC88i3XSvtdgjcUnxcaHz9IR637IQzGdEQhp
22mgwaj2fxhwEaMqukuq7KBhsnCPCnOF8lzd/DdUUpoPiVjvYI8rZGiCUkqksFDs
t2YG4jeeIJKElRE9yInes/GJMsTTo7tLuglyS0Tly01HCc/0vX61TCaiS2KFj4ob
u2styfRjDp/5l8UMim6WAP5cobL01kVb7PuN40WMns67n/vOeyyjW4q2jP8eymBT
au+lGrtjIhrBFxgujCOhkh0f2HNP7yZiq5IPGzWUpEymeELVg5ZzJTZ9kH5J2Dyk
eRK6Cnf4i9Lu1tWpl0dGHlUiNian3yNiz2ngWzl0XY4bmoH3Vk+2yTmXBIgWBeqt
YcLQVWG+UIp/odcc8APY5GUwa3TTZ20SevEAX4EsMG/ey3DzpMgeBhfyhync6Wos
rTeE3/N7ATTCTl8t0JHAObKFzVdh1J7peJeLRBFJsofQsmdgieGBQQt6Xwsf14Fy
coK+OZEt2ViCkk8puPhi59JUDe5VkQ+Oabt11VMpNWSnqgvn0wrB/XS7Hq2F6Mrf
L+MS5xk1gRzgtyPDc5h1MmdaOBUooufZ3YjJrvijKsCT9MKv8wAIcrVig7TU1hA+
RvSqZ8PoWlCekevovIpXOycUUtVNf72q606tGDyDm9Ejnj61PKltcMJGYgYHgHPB
UhK/bWFH6zm70HJ1osANzsOiIZKCxkwnRKv1guf+0qYJrld4R7zKGLsznrxAtXLa
GxdIdmU1kvAPDqqlYrMT2OZoZaBa20Pzy1WodpnFHex9p1Q3Xmcyaz8gocUHjR+c
6mXaLB5Yf1uhe/DoykhtyB3xAlnY8Tst8VHj9birVbdYiJN5SAT07ahYrbQXqb+T
LQQVlcRHCrKMFzoaFeqzCAmdg2JM7abBdA4SlYx/4sXqEBp/iha9jkUJEnq73Ask
XzUSZN5p3MozjlUuXN1WcjUmaIS6AATagSU6O3BqwK9iM8Y8WZW4li4vMTm9p7j1
h15vdFEPU4Xh6vsdEyIIBLovyPZknUVahGGEkfu5TsY73hlsChwGlmbaydTon2+S
GmeY9eFCOS7bWxzXcSKBnDEqCP/vuVDcMbOTfo+uyFYzEMuTfnhsI+HOAzBkpmKP
gCs1O+zYrGHzz8S7Q3adSeeZIFCJd10IJhhRi2/dgXcGzPjnu3V6Lawpt57i6M/X
cXv9vcF92ZiOjiYyPXYxXZ0DcKhEfAn4cFAvfkTp9TwJ5cY0qJn46aWPOvcQn5L7
klRWCKPPnng0wPupKcqo++a6MstnZcenFAynm/h2HlgkmEdFYISSrMqnQ+vIO9S8
Aqvwl+SviXO7vk+4Gn+NEty78V00+J9dL4fvYroq9YEh86rH/U15mGhXw+FgJTM5
3XCHJKgRUGWH0v1kK3rm0GGTFm6uPImndyYpCtw1sJTSTDAksXcvPl816JSQBzgh
PkFItkogTwK4b3at+zezdRE/PfXg7A4dEaQRsMZa7j8=
`protect END_PROTECTED
