`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SsTZFLqmiugXm0rU5ea5Fcs8NQNMeOUh0z9MTdZBvnRJT5hYcXbGmx5eK9Np/EI9
sc1DPdn94nGhRWGqibqZo+ffKYtNJS86yycIgNpm5OuFl5YsRKT3rDoyJDLaqEgj
Gl1K5mM6xS0Dy5YriJvW7YEvztgNMflQE4bweahwawM74ws8inxklQUowebSu+Z7
x+P6xM1sg7SEu3Oe/W5Gp/V8Ccvtbu3mVbJ598a9bSUoVNyXtmCRqd+ZV9cde4da
fDIxaQb3cPcmJC5lS0DqIq9XzTFKhUui1BzvhWORRdyH6brgqwGASUuV3UsMLBfV
lOY/ncNu8lXrV6hXTopwu2xiJ6+EJFX4LRblOLmfV+IovRt1cNp5DZpli/+FUj4j
9/1CnaXcHaOZ5q6ij/BuuAmIzNDC0ts0GHKQJKWcDcY=
`protect END_PROTECTED
