`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qOMDZ0mdrgktwZjmoLommPUtsDjDGDxC1noCWOJLnhr+QZ3hhr9X8L8G1HBiqhYI
RURjqln38++F6aV07udh8pl9I9k4SJE/IJE+qc80knVkvPn1QyLYJUwmhA/nQfj9
MFwao0txtaSnYrwNGnMMzZJxigGiX7vu+4+bH57jA/6LhMQytzYtFLUBf8QFRxQu
sIONcuBJeT2zxhlsob545PKJ8JG58k3li9IDN7Jk7ZM255nSGGZrVRjXZBTlvuqt
Sg7tufLteWlZDpGcurKcEB2UnIQM+1k1SKD3YotFO+V0kov3anGBf5KdnMCv+hl4
fcct0SIj3JYfh4TbVQMPyQRKwhKptgmAvirvQVI5CqscRQPxU3R4zNdlHLufVcK8
FaSuhF5jjMNH7QcSYSyIRc8Fy/qm3W89QmYZgVo/h1EMdSM+W+/zl+Kxez0kaPF6
0dfm4Mwol7Xj1lkmsompm25mld4AQygAmkpu/10/azSh+9tL9i0pTqwlRiP0JPsv
sdz7mM0Kqfu64InecbU/wxbEjIQ8ANghnx6Y85p14Olpbi9V4dj9qAPUWiV1Xhht
AlC/GUPR/ukm6aHV6D1/xxpabi9T/u1ovoziTNMdVTaCs8jQY1pIOrTdB1/qjHuC
FaWYat5+rAqBhpOpHiGM90SymzIXC8mMCmobyUeOc1oLY5viOfaXfznhA9OYDNId
7unbCEKbCWduor7kYNL5mq5fSzxqRME5scYIYT2KoV9ht4iIXoAcvI1c70eRcp19
8Sg6IEWJHUPJKq/E5xOOQA==
`protect END_PROTECTED
