`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4hI8NgxycUh4DnciEzSr6pVQUeJWKw1OD4OygkiB4o5EDkjIQs4gexIJSmqkjMxo
OdCnp/6h3O356/mKXsVhLpWXLwaEiQmsU8cp/d8RHqoDkOl1ltFyRjk0d1HtLh9O
77vbHizOB0kLcHkN0/RBcldeqPcUIH6BGERaxWcq+XxI3RSHi3pmmr0GVoDhyuct
WSGnBh0RCuvTDLk2/zHnn3lUiSncHbPRP0DDnMLVzkFKmL9oTt+8GWAzpHzLZNpL
fb1nnl8pS/00ggSJEptLMGa3qW7oK13iT6Yd/bNErMRHYYh1SfyhYDLtExMqtnxG
Xt2tnmtVLWiiLE3JJp1AdZvpYYmAumdxipxGwJHpnbdUCJiQsvCNjYvGRbKTdaFM
yKB4h6VCY7wCKve67iShH5LVNz6HkiHQHmmqCxXjho4F7A6OvEDPUH7COtrgtg7R
RTrBRZ6HKkkD/z272BPrdkhFa1s2EDVbLmuOddPLDX8wehIo4HBgx6d46DssMZmc
LGj69fO9z8nAZL1eoAytHyIc9W063IngxoeOIdur1MLz26xE/lyHgVPSpxvVOf2+
o5HL1Tukn1gdoAvSMKaL/oJ2uuizA87UK7hF0Ga5VTtKfnLwKG6qDUZJBakH9Yed
aKqSls9f0/TZPL15q/98o+M/I0XF9CEGLiBx+fEgb6k+2ic0rrtckDzOfpztO9PA
q9e5h7eI/Fqz9b3X+QPW6ADrmyq8FEtligBowN28kn+JXn69OS/T3xn9XoyEtyIm
CM5D4Lt76rYLbw4sjd+Py7fwr20/mxB80/usJXK4r5PwBWvzbFTfX8I3Q2JU+jfx
Yg8vHV6TiyqvbtLhKV1TK52J8nSHKR4AoVKs3bNL8JDPNPbbr/ESde6JprmDa/4N
GwLHc0AtpsozxjBKj6hK4S8o5s6K/zBLQumhVKXIkJwD97nkQveRoQby4Gikkj2v
6D425M6de8qg1P1IpW2o3Mv2YZoq4BhtmYxnWNyQL49fweZtN35w91EfxuZXIjaj
wYroUm1fv3Rz+qQmz21bTvmYZERM2JhxOQ2R3WY4wQdBLLnnTMwFOk4qvQbtRUCJ
/VyLXnljByN+Qdr0t4WCZc8iM847Yce4ujry0GVLRnBav2Jz1kgsd3X73b2R2eNW
YV3/cqcIg9iiDeYOLSYngY2VhuDYGIfKFFTGLWzmpVWPFy+pbmvDlUz7CwXx3AnQ
WdMYdY+aQVofUX98Bpgv9tYtpv0VptJ4j0enkT96jM7X9ul8TFWtwUTFad6AqoaE
xVd8CRZRk6lalKa5pxQpKS2lz1xyE9EjM8cdZKkOz4n/2xglg61uoMrnK75/OMC1
Yc7HMyaLYoYTxln4gXaYfpHfngpXVyA0ln8rxjkeP8Hr1rv2IZbGe+KPZcljKc5T
nTUEqb3QwOJvnFeIjx6Oa/vE/Vjd4W2Zn8sqNewpaQK4j+BYB+kRYAFRc1JrgrI+
rtg1N0kFpPeuQPJvVwApgdVviKIOsNwXQv8tz5WjwDRCJsGlNlPkwMCbCGyiBOwJ
Sa7Rn3gncIvQDLK6TjcM83irfmbOMO9XQm9CrYx9+94QseS2dXnxrMLGF21STglK
u/aan8gJ5i9hlwT2bW2D5Z6idSyohbgsbIPSIii+/+QGoDXjsHUQekEbH7ardMbh
wu6mQDvHWn3FC5rEav/kNynEJL8W3tAMrKcs3woZpcsn0FZeEjgU/R9ZOszNAkW1
hDWpAHDYe4CctAB0tlO+/s3Y/Tbb6DI235k7z7J1acWTp30W+IaQsxEwdHc9uh1b
0QQ9jBZWuuiYqjGZpXexQIu4mZsltUVtNjsNil+DykBb96Plph01XvxoXqL49fWO
KRtkWsUNBmCXPQfNvQhbG0kpHG4BaoxqoKhoEx4DjBCa9zqesUIGPX5+K0pwUWrw
8UuuYf0xIZdtVqovzkPOU2lFrZJG9tVGyL17ESk2mcc/9WhA4Lpuvr+NQhXAreWN
/HZnx2OLjnhzjCm17t0jolrwc3Bfw39kwgdEf7Gd2ZLNU4Ii2qQUtO7cFJ8nM7G9
vGkFcdltAlGQOK3F0igO+TrL1+j8HvGS8aci9a05UwxyG2QVDuI2o0JK5osdH4go
HS2oz+LWQgJ7iwWwI5r5rKHzhmrZGxKVbryGXZ7qYcTwjEvgY/YH8rj87QVJFW9V
hKl/w96j+7UY5jXb4+e5ytK1uksrBzB3+k8sbIgEvvFZ03V0cWSdUTIr0XEWH56q
l/Z12Or+jj9fo7N/ThIBA1Qs6CMjxYmH1JRGT4y1mkdIY+kO7/BJZmxu6+irOSe1
ziw1qyhIYVwvkGgT9dC2ZkbGaqMwJXHaSDaz7HdngPkzPz/MkD1m6SEueelTjOnB
wl+waEYEW8NyS6/UXkB8CM+11f6D28SEoqvxk83lXYjEj2dNt/1WyLAGEz1lOFQd
cf8LErIdTwaKKeE0FEHimFXmQ4BuzmNvYPq+fYui0Dnq5pe/dFatessZlqaTIOyA
QRNwld+7csKJp4Xwt8valf5nN/+V91ZN/tIbjyG2mKon1P3PlCAr1VrjMjx57X5S
eYzzAqeJxKMILKROcbB2fynmNR/26U3fJE2tMcEeLMHzNHKLfybO7/MudNvuqjEw
D8gDy1R8mIhqCEHT9ZAhJ1cPVt8RHmkfZUwsQBMW3tvQPOMJUOlLkjETZIAHRqIg
8TK7W/hU+hctMVi0zttKkFJgBJx257B9OTowyRcEXa997iAM80QRdndKBWeBb6nD
jUy6xfta9ch8gMekTLPFIxCPlqjNcokYeoB1/ZLTsrqOV/u/wLQCEkSfoWnpJJGD
99E+l1hU7WHrX70DqiH8eWYElbcU/FUl8BmphpKGrWC57vYQnMfTY7H5Npg3C+8m
9odxR/QSpS2ldSkrQnV1VWBfG/++OTRYdfvk6kTgLn62eDToX3W6+bghUfovcdbf
L3QNRWr0RR4Mumfrom8DQBOFKpJ3dlENQF4udJ1NVHEKPABM3hPzvnAf9/87Zd+m
o7hfkzkSTUAp1kTtrOjWoKkoB4FBKnNDOcA7R65W3CA9QG9g48VXpaAvMJ5oVnRx
EESN5umk8/oi8FUvGcOuRTJTSummE3cO6PsSFCx4vGmRU4fVs29l4AT7lX4/ww9d
Md9aSJ5h53lgIJ/e2wtIXlmJRgEf0Q0pE6xtFcZufWSgIaRQgtnNCePjRifZoAHO
f4IxB/15T0Z0li8NjxbuQpE6YUm6Mq4cc0E31oaU/mfF6oDMDyO5LzZJ+STotfgJ
vvmZmTtf6n/LsLkLW3ssWXUKyIk1aIW3o+nbZPEprUTe5szLVROLSnbe0OOCH/w4
ribHXwlSgqDxJaFaQbA07rDRzkBiaABPU+o1B1nTBjMSGmEWHRnsI6FJXzYWoRUW
eI0q7YKBSs7vwsgKlKis1p6/QRMu2FBCbyBXCOtpIGKZMnXk9wTsTp21Li4CEBr1
jcZpUZxeT9cdOIkFJgZyuxHitBXV9gfMv6bMwI0J30np4Aru8ifgOqp7Q4EznEEK
1gIRm8s2st0t9mwqETVWuCpV8VtcjjvUM0geWkU0Yhf7T2jU0Md2YMqzZgwOXrp4
nrMGHNmzenj2Cf6OWbkvChIIczz+Mne6iP85JLcOkSVqmYzjd2W3koBQpkIhfDjo
barbxZYXy6QXuIR5P05wj+CxlJuqo4fGWC6gJ8WW1KrGZ5rKjxiHf/5lgl5XeBd5
aB2w/vJaLjnHk/814iWz0FSDRJBVC+5gh0/oBpZ6jpiTs7AiJJoblydL4fIIcQix
MHU6lpewvt9mcY3m4gDjyLayXxMNYxaNAeUv1/Fu8LMfW6b4kRnPwTU2M2plY4/3
mFxWyvyvv2kx9lXODo02TQN+PnCbXisVU/Pah3Rmednrz2NY3ARKDXk1IK5flb5V
zmWoWLCgq/WKsz2Yw0StVlTMISukLmE8u7uG+8VB2E/ISy5nOyxoohfa7LWKAmfT
2zX5HlRjMTkNczPohn8ZM3i2ziFnFQtTHznKylnW8xsaTkMuve/6gGpPN5sogBh9
4KYOBkY9aYDJb0cEjvgHvlGB6SVwkN8wgvMnBb97B5Uxy+r7ro4YdSQ2r2YDw/32
iqJ4B8XSSTE7giqVu2yv7Tam5DWYoHk8zbiu/bAqS+sU64K9qUFWvp+QRo+Auk4q
TLToZ0RWBRVLDc0iXTe/MHngOuF8turt04YGmI9AlLlmHQZsU8traYKJfbV5pCCE
9OXjPcn5TjsLi0MbBpOe313l3rOgSEUzOC1TFdCMv3M6RbnPEdNh6rd866EMm0cc
7ZJpDaCpjp2pqjBpaeccgnrmdHRDlu0Sh4jT1hbX/UEkwsgMaBoWX1fCRes/Mlq3
cb2JqomPetGPQlG6Rg4lpJpIG876XR11ZydxK9bgquGVWOiROxDHx4AjaHcXVCVB
sncifbHIbu0gXR8tQUabsqQU0qukzwp43gUjisxUenC85Zt5ZV6DhvtRasmWbU90
/VQsruJH8bEon7fPGZvDmoJHnsm456zxFKzoiuVm98kWn8q2algYX6RUIvkcz5jp
c+tZesixjNJkGPmI9f1lgPd5edVU2gG993vRdjBykHQ1aOlyGj2PoiY3LOj5mm2P
EcoKWKOU3ykQhyEmM/qg2xzSvqIXnMs1EOYs56moVYOhDGdWhrybLoRGrdLB9msu
gN8CqI4snz4dNN7LXIh3YscYDSKFXPX4nH3WmajF6MCLpYz+6/WgXQEVclJpEDfR
0mSHGKfpzI3jIomqPh7GvWH9dPJA9S1SHtLEO2tDKTw0l3ic5oJ0VVoeWP1e4rHP
c4bYvVsS49hnw0iMidZOTJcwoV02YsyHKO4Xx4IbnMrLLkkMr0aMXyquGxzXHvTJ
LOWNAeZ9jCejweLF11+PSwxM3s3jJ3SnjlnFJTyvco/tkIUpefByP3e2IW6odLH3
7FmLx4n0/etK+wWAawFwQTL591kMml4e4RyTxQdROxbi0aV8uc2WxLVxexDgUNwA
a+x9BV2Bu4x47T2t9cGI9fTLq9Hrc7iAzzOZRKSdrXz5DkHR/dgjf4dppbvCW7BQ
iIkAg8bOAs5jMw9+pCg2Rgt/2vU0t+mkdCuxA6l8aWCR0W67BhqBLJ/b+k5mCmmA
xE3cihEMb+BySTGiCe9j2eMe28UVINBK+3U1LveGKE7Zeb03HjN4S6z7eEx4WW1/
FCYvRAtU5S7AzsoFlBkbUIgsEUJXN0PboXVrbXWo7TdWdHrcJosSDcDqUa4UNMMU
w7wsIeOaS1++U/z7BZaOfc82Li9hOmuoKAflQJHViFsjiFA42y2+O95TaI7YYGzX
NPjPX+GsnFcXWpxlBvs3ujAsYs+f7vJvLhY1RKW7bct+GZt0hhNmGgm4s5wmY/JL
PjFRvZUpI6r+M1zFC0Gk3mm9P1zuCpzORPO1kEdtJ7QxjRR1kUtFyiWengCGZdMa
5isHetJ1Q4hrQpdDDQv5OIjftg+KYuBn03j5QxgATzxviObCWvfOTO6JoC+vNp6F
QabCrQyF/B4meCr1NbJSy0hqdE/jdCb7D/7tmVk/8ds47TtqmluGH9xoAoLg24NJ
wODD8RuLOoPp4EQBFlCf7aa/aA44ERrlNvRwKklGLWNFcyz5VQfSTEoACYgJVJIh
+bJ02i/fbblPfw0ATKaKiulNMsRePSM9F94y+5Q/PcdgrlLb7OF7Ugm6U6LxgzRI
xa3W1E9aL+7Q5Ubh/wGx24VNOeIpsA+gM/rV2m9049ZnEgzUbmKF4QP+GYQMDoIn
yvQuVhgclKUHuSgoPY8/GTc1XMhpbG3q/ffDxZBfGg9WyZgceCDZyj6BoiYg6jV3
KBP6tA9RAiIRposud8/+ohZ4qUWvCmrLCFibQGRnY58xbWMTBa4NWPT30diKWc+g
KzH//vZTQVFDla4d4IiiHitJvX5h+GDJvOgtV4mXIbt1rKdXsJlaGvkE+Mmcp26Q
VAo+sowacfxTZwGe0sX4wgDuLM9rWxL2ZIAEWufmJYB7zBrADzF2Jz9tRMZLiu8H
JuBvrWlO0XqXRKra3syyAiDOdUuXDZT34VpFH8p5eLy9Hps+rhb1OSJAe3GIIw/r
RbWTePMxDi16sGttaiNamugedhpE6JK95Xjlj61Nd58AhyZFqgMKERhiFjTFBXyL
OZIB0VDigb8WszCsMIyPJV0xKVy7Jn7qoACbGMnY/n1480It8XYf+bozTTa/mIGy
7QYhX+gE+b1bsHsAlWG+Qxn23XaIrlfJCAdmOvjOsUXsUdZ1eV1/l8+cxtFZ5V1a
aPhs9XBZx2YcwnUY57pVsbFrIbQZ60Kpmj74q40n7vxYEWmj5E5YpIYbZ6W3OtTl
wMmvtTcXRyLsjuR/cZzSSZryAh6t5u3VtojljHW1Ad1MDEFREf98niusKjYLLC4E
+itx1eT3LMjfqgN3RIbnCgJrKDLbdBHbnhJZ5LQ8MN/GgwitosNB4x0eWi7J0byr
LgSjORLoVecxyqKn9ZMZyVYSoFIUgRW1QkomvRWjdyZZv7Ay7BI33tyqbcivWzP6
hbnVc0RYr3n8yv48ZlRnHKGbZZMmkR6SvEBW2extr3F7hZz8D6iqsTEWnk9MUl9V
2g+jhT0smtOgn9m8O4qZzXwrRnbhMOE4jmAMonC5ulSyKXtRPIbwpw0PScI/q8x7
C7DwP2qMnP1QyK1b2v0iN/wQj0/isNCHE6cYBRm0WZC3CJ/PFakPxKXJgSkh9Hrv
aSSwsSE9s7Dw857JPySu0Sn74Intki4Bq+KIfILp4ovLHL9CJRfgKvy/KM1d/lXt
ja+eMNzbrbcH9odDjqmZFpUNyBLEKh7M5uFDmCrA3NO++nNSDD1pIEjIMazuDsGH
4Lw9N9EfwJw1y9W4jle3tHdTUfH0qNg7Ta98UK1qQVZcVDVAo9Tz8HNiezUwNbye
UCxJYZrPVhGBqfo5j9bgzkkKzJ+ObBzs3LjhUwKbCEIuiWD4FoctOTh4OPx3J8AU
7v8d0ERrEqfQzKu+KouKSTQxXJEyRm+rlSqyyV71U2ATWiP+5ryPaTXvYg6r41IZ
WWnudt1IIbNXh8vGrBoOEYiQn+Uepu9nY0mxNArFd80Satw9HqQal34Dj/Rx7nQN
fGCLs3/XZtSYZYMFm8ZV+kSjUwjH7C22kVnODC/P8Qc23IKPreMQgeh9Hs+dSFuj
lqAJy9VlKiLGMxLA/Y2WMS86OR+zHdS2xyBc8HTLNTtM34mtHodrYIwRquZqdQ+k
UC4DTLAagbBFGY7r37XXI/idc6FOHxe37M5E4GcfgpngFp8vW/2TJ1uBpoc1ZKkE
PWIkkJrlnXnJL4Sqn/aIGzvk/FWYhjWbcq7k97zbBujj3S+v7bNllWXPpA2n7pbu
547/2kzq4IxiXM7nL4u2e27UyaJzMv2xnX+v1UEoRDQM6EAXx1dVP3XtuD/6ESj8
g15nnYXgkE1XUIUaYxyAe+To2DaWbJmj/aCzYqHm09GN5rZQD/VaMs/loXy76Mrt
utJ8hXTp6198WLvf5arf+fQSdc+l4UHvikK5t5ARrFjQcMVB2jBM89CwVgL7WqNd
Phg/rhp6i+i92Yq9FqPNJzdkCOZCqXe+U0oTF94y5kLC1wTd9ed9YOAnxi7Tp+s1
83OjmFYA3LWo8TNaIay+R/GkQ4PgfMy6CY3tshPP9IOuL6eB5vo3cHOqZIOqzJEH
F3urvbpq9wxWBU4iHKiFokKBNOf0yAMLTtkuhtPzLe1eUaB5xKbOwjUe6WW4Jx53
Gj4osyQiy1CsRcNF/UX0Ynia8+31qGrJK1Cjq3zTHKDaVPlO1Lpq71m2IqREEmri
bITP0doX0L+HEMotbmEIXBkSW3AGlB5kYZJyCsbmUOVTxfKu9xIXQqQRzOB+CQcV
UkjvzB2PZBiXAm7T6c5m8gqMfvv6ENxJKQIstcg8w/2Ta/8tDh7Q+yBQ8iC4rAU8
vTW4PNN6VBN7l2l8gaLwxXIPQXG24AlpupcpNcOD8l4xpO0f/C//1GUmxL4TjsnI
Il1510YqXC+gJ2ZZzvrNwXH4J2+/WKaQuW4NkS6pW8C0mb1Taf0sT7xD8fFK+NBY
HXvmLkA6Iv5VMUWdJuQfQB1nCrfk5LqU1CT6phgmzRbSE+h5F7I28oY7YjtPAr5f
ceoLvEOx9tvaskCKcbeswzmjqsZw7LiKzMz5T3H41cUnYPAvUO9RjPfpo1teavQQ
yZ1q7OHWgr1NIMqna9A5PsSopdFOhwMXOWuD+lVOA/GROjJG+36s2ILPZlpt80Ws
iCfL5p75sTgPOy7QRcAm+V7vDmSKH1zjgQU51b6L2+5R38vpdYcIwGY1i/0DgwgT
wSKyIv2YJpLr9NItf6Kp5+t0I+38iqjhzDgMmNXIm0KSUYgnMGZgZTj3MOqlrMZh
MBSOc1D25JnUZwxobwdWZxfkcedrqwEsdOamPM7CkfRDlCIszJHkh/DWfiGwvsIx
tAu63Ii+9XmX6QoMirakio0HroVZAEdubLZQZR2W64GmwKAq8gkDZzlQhnUkPBHY
LXrAJ2Q+j4yf0Qui+EXqp0Bqvd6QoFsxZqvCJABURdsmn0BfKW8ybDG8RvcNGaFr
bcwHxMk8ivULQbizO9+Kq/TMbtO0K0j8Qu4uZYdFTRS9UAvaUlc/BEPxK+cxhIug
XVBOuAsXTqFLPcDdZDj2QguckybTpumAwmPBCaixB46HcWkZ74Lbo9iIw5D0ox6Z
Cm5mevEaAmkdSVPkFrO/qFXXKSmkhnmdhNQgDMHqPwygIQ7wT+rbzY2Dy5imx5Hy
iwL8CM6AjWvKM5TQzJbQEeg6N5z9huHWStzkvWSoysF4QBQKEhLjp/DQaMKyyzOd
krfIw1njGrxV62ziLy4IbeJnJnrHJcw+Ttkvqw1pd9kvT8CJNzVXMtS1nFiJv8Yi
RkpEJ2NiES1ZnH5oFK/v+9NG2y/MPaH4sbSyiG3vktK0g65hRYb0orzN9SAEN96U
DZOx7Y1TF1wlqKQgDXHlI3ZBkSrMRfaw0ZnkprUTMY8l4ZBgQ2pgwz1xm0GoQs3p
SKTu/ue040lAxdHkdv2Qn1UlsUR2X/jQrr6JK6HCYYM2mUFdSMNs/ljEKByvby9o
qBphpPY6fs3UTk1FSvVomYy3FZFHfNBbIoCQJVvQXsWf3n+xxCS1STb+QiLBjEKZ
WULK3OktTS6Snncx1fBtWTbzwXwnIVwOYQmEIVJpezsVfjisGFy81KKBDCERgDZB
Kokc+zph1TBzgmK8VT8YKW/05475AWZlsqFHtFWmM+rJaNabJC4+93ODIc2uwrW3
MwC8Y1j3rt2v0HDQj1I+WxcsfQf7DhE1vUkxJLcPMs2dMIvr2N/wTTOGNXejFv/7
SWWg408as5CYsE7NIdBvit0yqrJFiJ+oPGa9ml/PjDtJ4xonegC1lawgtTdRh+yO
2LJMMJwC3EG2jc3oI27a279JrUBgqrPiDi1KCxVPOm8bFZ0aczhAd8YMANbEf+4N
4akgYgol4NmKfzbwWI9OwBQsenRLI4Uze6s0wP97gclm9so+3/R2+xbbmWPInfQX
0tTrre74GcoAx1+WvkLaSc7lIJToQYtU+EQbb5CgJ3xUzNkNUOUAfMbvAkKeIQsD
xv9kS0/wH59tVkk+24Fw0A2HPYEjkVDr0aI+bANrJ7SDUyJmC3RydUWPhh7fsmge
ZAL5IDAUpUoeUznyCcr3FYv24wL19S+4EhM8vOvgPVL8Z53ZQlcFmZZcq6iWKp2t
0fx+zUbM0XbrQ8vQLQ0sJrntagUL9kNl+HTJ64H35HedvY55OzXCRFzabN7j6+/c
8EE8Y27tQJxzKzyok1q+6lou1nS5wkpgBxfE3ti1Y6fEflsQUkfAlG0+4p4AbYK2
dNf9oED1KFLGKImThcoD3XyAfzA9B7G29a2R4ikDO0sZG/+/q783VKcH3Wjee9fS
stNTVSJ8MjjMInwHg357EA47t21F4RGCF+7dWlKtpuzp9nh8xJmEOg0YR+DcSGZj
sARH0/rpvH+8IqbgyX3yUUKkESOM0tIjdZsMFT8QzxuHQHaR1butv2dDYlG8UPSK
xklLoAp+Uk+rB3I0vEelX+NG5gxmwiIhJh/FsLyEUNs2PSD6Dkt7DvjovoFnI3FA
QkaKgUcFH3rbZboH++A2BKYx5nXNEsILOCGL14kAlZwJxhbJ70hpWksNCWgIDhGW
qu6N7056FZED4gPF21yCOti0/iWnoCsWhGmpsMoIgC0Ohy7OipVDG9ZOqgc7MSgK
t2j3cfpwIfBobWaq/c30QwZnCVVNSBkb7Z5ylgs6yunwt+kkWOiQ3uSaDeXU4d3X
D2Ri3iYGfXpLAB5NXjCgff8spXNMm5VcHiXrNpiPvhOQBlc6zs0yqOhMjxGIUe7/
AOkzKntBkoDYpvhhLmLeVakbZRMPsSiLcgklboWhMPhBQDqYjr3p/UgE5sVNPRv9
WcYOu20jl92XKlYxvKkwikIDOwyiQf8igETL9QYj8p5KmVT0ITnk4FDb2WAHqke9
lUImVsLacRdT3cEpwwMFjW4rUqIh00hyXNTtUQl8bHEe88EXqcZWqYMUwJWteKeC
xLLfKC86mFf+3c07z2SE5+ODFyXi/IjWESPUW50tgNwpUIujgVCe7rPzgtRpsh8o
lHbhOWpNIKxhxB4OExO4dMfor5jVTLuemli64Wh2A08Vj4dLgbpTY1MhR7Rwrkxo
00OhEQpcr2VE6lbVObj0ElNwsni7vrewiypUDBHOT/SGkfun4BVGQ4VFtFKPli6S
jLi5lGT6PkzUKp+/3k8/YNETQgCpaLxJRUm4pKiiXlekAt+UKGbw6f9yt0xW3s8C
6dsFJbMmzGZSNAYzw3P3O/MJgD9qJKqW74BtSncmLOAL6CwMn689TNgGrSc6MxWM
dXIvPznit6ffNZhRbKsBnGt6eMm8GVgqNsJdr9aBajDZyBzJCTaTJeVXvVeYmBSu
/hITHWg+aA6Rwi9z+cDEHWUS8FN9VVHzYxIG+pAK4PDdefo+bQTZ68zX5NsMYk8w
Sp9+i1yetbWjRMgWhkbeN6psWPsTfSLRUFowhaBBQowahUG6N6AE5ERBNz/qoJJJ
s/dsjFs42rnz7Nu17/ujabYhl219e+T4yv6itQuDbLLscagn1nyWNSJU+ChZr598
lBxmokyBivswP2wpFF6aa+FQDQ6C5ybOQfP5ZGqq6wQJuZM3gAEVUw90Bs9kOrYO
i1+vsk2HcNF2yTRL3g7QumRipHKKSRYKLnep55zqbutv8mbV4VuAS7J623MoXz6a
eoJqHs2XXMdfZZAXoQsbmbvlpYfnQLoI3LxhHLp5EpG4akdvircsy3TIGRTADbx1
TNQa7wpTtwoTAuCANE/8blkAf9TAF7GI5Sjymxvdztq9ClH/iusGShjXtc+jAsFC
w+g8Q4RR4tEw+9jK/17JITv2bvKtDixEHbNCJgD/mVFUUUDAeN7YdCjX8au3cGw6
UMs1xV7sBnSsQK0HUABdk+K4kKQb23wcg3XkXpybHNYMCJ7HUJhoCgVHzdUPF53D
QJl/D8cO96vi1heLh3jgXbBBidb7lyiRdZYsYb/sv7BFBvbKvHql99zEVRJRJDQy
VQ7uVaUCHaAQJ19ONwrWyVV2tZLm0Xd8zx78HInyhL7/zLyfVXnm5NjxVp7dIflD
3rBmqVWejmAFpGRiyDyS4LVOA1aeOb0Xm76/r87Z7YmD4UVh06aSHHJTrC10z26w
VV3zgLp2rWdNneWbmDuFAm1CZ+nXSc9B7NrumTDdXgHu6wV9Ug8jRdqvvcgPqaXF
lAEona9JGMVVu7v0euxg1lMKWYxew9r1YYkrSfX/bAuxSPpC74/rc8HNFS3s6IDb
6F60r82UPiowXDc4Qk3TYyfi5ryYRh1s4nVtw7YlZ+2TgxThrY0tKTk9MNGbx/KO
SXQPGNrmig56cfwBGaR2d6Ka87T67dQMgqT6+83llEzsQcDB6meNC5OH8AOBBd15
MqtN1kyAX2INkvZihNJc+wGWY3cXbDqQH8hovEo5VAZVvfn65amXZqTQw1kf3qWS
dgvaSrumfyVIRJD7gK6RVHNTtUs1JFD32Mkau5lwsePhxm3IN4f87QO4PRV5iOxc
RZpGpWi0WygCltsquyN6XmguCg2pvMIMLwbCl+vKM0ReuEdhalc2TC38qYs1e69b
Fml2wis2Rye+2omlM027N/vG5DWiyfKH2cfYMAMReVApU/P1PmrcZGczQhH+sPld
5JBqkAi5MvP5uAaoNYmJkkmPPwWlBU7pjHcmUqtNYyRdE3MCvW3BwDk+OGhBe6Hv
yoOZTBoljtpSO7Pq1fortI4vBG2byCoQavitBZSOFRJRszXBmhs1sivZAf4Kuu+Y
ncz6UJwk2acw7aSMzxvYqhpen5UoNK8e7u3KUaXYZlbZ/4vlbEyYKB4njJptsHsp
CfozSLlqMlmWljiU6Qha8rSMPTolD2M2H3pERF1/oqo4DiKS2CziL715C9fESIVC
RUnnyP+YLiEnVWNAJ+XOwfWPZ9wP5YTP8QZtUS/Z/AviPHTQoZldEE+Brq41Iz6y
VNsNcDCZ2Tp48RG3MZ/Kv9PcEOE5JsS1ai0Y5FjyfVsVIYyOOj1DLYat6nStxsmR
CKEZYhDEvlTeD8Es4cpTSSfmo5yZKAwCB5qtxxAokcq+QCpnteib5O650IK6u1zX
ruz4t+JI8UqBypeAEsY6vITjUECM2oFArL3hTmsm/Q2XyPXnnr5FYQID4zIcapW6
Mfas7Wol6R1li1TgthNFsbglmItTqkNF2+WvJ2refPpOu8CoEkVuwQQT88yNMxyC
Ey0Qip1wP6uNor8ywkb793kaTJFuWmtMbayfxkaXfCmTX5BGwDKMMzBMdTXRbseK
xLM6mQLnG2N77nzkYVf8XQfnPTnPXV9ktMRDNN4NNNxNqVekDnIIRWSemf7bNI29
K4KAJxMNhyiyumzwhq2eDtHobT63rNt81RhJg4SrmY/xAIOEW/u8LBBxxNcirT/T
PX25ZOjoO7g/RXqb5sG1Os/+kRhVujx7ueqnUgtMvnVvNfk6A9Z52XwtP3BOsMHe
Wm6hAKbdawp0uUCilVEROR21X79s1kclRsF669CyuOwizCNJ+tAokCKhmAyimcjY
8LQTAVRqhUAGwMQ+47zDt38wXGQw6YW9mrfxRbDFPdIkrBVEFQoRQbVdpM127o7M
4zQr8sIoANxbOozwsoZ1ROW0oPbF+SsLnlELwgISEEkaDApQmVGPajkpbJV/yCi6
PXdeGIKURYQJ5iD8qHoPIkhVvGvEmDcnO4Ch+VnXWEx09/65x2ZDJk9Z1oCS7dDy
SBh6EE41dqTCj3+C9b/biBVk6bJr4UzSLX0UftXtAVs=
`protect END_PROTECTED
