`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qMLiepgzaYTTDA5sO9lYL+78LHeNaBVg1LKq6qfwb6Mw4lkBrlgA//2O8rNb5bGr
P0VgFIsjOchtQ28Og6qyrJ4CzttLWNwnuoVk5TXl1RH9piv9eQ7ZTFoUIDj8qWCd
qDQn7SgFBl5jjvaotQFtfD6dx0G25miiST/IXjtiTIZPOindFt0TN5NS0FN+1W70
DBLwhpPua6l82cKwxEAtFPpqU3hpt3vri/wFmS6HVO/CTqKFoXHiQZ24eJgeORLp
o0PpkGWiguoW126W+MykXZPplqmIPJyUBvpTD96kmNf/KuUTYb1mYgz5+rBbu+M4
7Q0+g0YG5wCpvErMKsH71r2fTc6/IO1EvXfB8EzEjmAxTKW9sI1JHQTU+K0XXQG3
esqfQWXYOcI/aV2i2Dq75fLLwJBEu7mXfiSrSn4sajEb4umgxXqRJyIQ98LoKp4Z
vH3HZuCqaKrhgqwROsuPstc8pvQbFFgmAWwMYJhkDJuyTS3cpN+XC8WGBwn2rcPc
Rgt9B4vf/rzk1C7QyBrTwGxnTjujQrGN1ue+IH2thII0vCuYn2CkyTdsqnEzISzY
tlt5oXu4Ru2+KbHr01B7SeY4V/GWNicMnUwBnvTnsWHS2sS10PsQ2QBMrQJc8V05
lBi07K0NL2SI+XYDSqbJngyOx63MNrxI9wNM/0+7A+i24+n2VI5+m/XjVyeriHh3
Y29xcLi1mg6gFSW25NPlcKIptHwL3AHR48lKU3sck4sRUbU/J6qD3Q0rlyP/gcHr
AY9c3xzwTClmURkEunjWPlyJssLlYTYl+zRcepfqU5uaI53+Bkr/DU5wciu1I2hS
tUFZK2wab7UIfn7H+0GIBz7fyATtc6b+QM4MbEJ8V5dCVT5Kehl+Thhpz+BtE9vk
3o7fonbnR24sc6gpQIINVKgkrgLfC9DEnn5voZyTAkGTJqiwTl/gI5GZS72eC05h
bBLSm8T3eINmCce4RI9lmhHhp4HklQH2E+FHS9KusQt9rbQdvnONZRfHNEu2fLiY
eP97dTLTJMT7bOY+UIbTCTR9dWGY7Grv6bLQuwMygkYM4X8yIm41Pvr6BTKu675B
qDHJDNP9zlh0O8jOyhA0qqGzfQrEwDnb8yvEEcCjbGLzgr9leyOPt4NdMcRSa8Lr
NvYhCUJ8T0EAX3rMON73P3CEdEp6OHp4JK3mIXa0nK8d6bsbmeb8XVpzxQ2nfB/6
t22JeNAOQxKtkvtz14Hk61x00cUEG5R6uEvb9PfXO3NPTsHaKvA052PBj/c0VpoL
uNxh61G5LAAqsiZ4bsh5cFeEYs1c9/iLD+oL4KWBzefGW4TpaCz9PqLha7x/fVv+
PBLu4qjbSMxdTbiXNst2tekZWpQu8+zWijXO23/6CVFFoOcw/ni7CFtwtlUCCJk+
upVfQ3HqIDUlFH9fIMZhNAuZ788YQBdjtj8GbcfcaJg5cz3IZgrmH60i0ts/E1Rf
HwugOamNJrNrlut8Z2oEtZJO90xSiSMxKkvEnOXwmOZLAKsj6tcXKGFv7cU6uRoF
FPvVeCqB79Vv9dnIFkZbxeSPkBb8KAGsBwUzftDHrWxbyl9OqCjHQYeolmC7+jmw
tfP6BzqHHITwn0WBceJtOCV645c+kN3HBEzicniM+GKvGhCXiar4khJo6pwhohmz
QRbOVg7UuFWlnXPSz6LgzgeatIkg91CR4IeDHLB3AJtLrGaDB8CpFzPrWa1oG4NQ
iQll2zS2VNusvpKG68bhXCGPZeGejg3qeJCAHYxRVf4y0xPjeCmce8zehfNHN9RV
w70Yn8Sn3PYQnAQR9wZj0a5+VgOWGe5QxYxjfq7KwAGVc3nvYp6obizxMXniSElA
6AmiPzRqtkZygrx19nrCiztXwqe5jv8mB4bZBdXd08ljR20aA3HKtz7/n5aep6G4
JKUNhzw3Mlkg8ZiEoT1eJSezVi7bDuzy6pde5p5biwnp6e5P6m5O9qa8z2+oe1F5
Rjul5QUSWfhTr474xDXpsTrmgKW+J5yW0WlcsBSX6xFiC6/zkIir9mbFwto04WCn
p9vB7vRMJAQcgLxL4DPBkyALZNaLUBFRGtxQ9POEuwGCz3uNLP5BFkSoWfDmiUn5
Qf0KnnuO2C1pJTrFPJ03SCVU3uFmgqYrS1g6Qs3e34By/pikdkIWaLO06nh+llig
Y5DdFBhClWwwRO1Dr5PnGge5lpABZM2oN/WvOnAKn96X9HYtxAnOiGLdx+30ippw
xvLaIIUzGfjCVXz9l1z8p61wpxa70sejrZySbMm+gVFFskJbhVjLuqDogjSsbGvx
c5p/wWWb2kuA6okBWVS0HUQZKuKeiIdE+8Lq6oapibXbbff2aNGf/fWtJrsAZpqW
kv8qPIolzTBRyd1JmR1+4lc/Mx952apJy3uN1WzmsoIDcb9i/8D1dQiBsotnC2z5
Ngie5swf6I5Ihh7zVZByoSDhxYDek7XTe9Sz6mmBCpT5mLqZMzHllwnHjOD2xxTh
PNe8oWN75j48VMXxSh5saq4bm6+nNhpZXH78QUFjhQIvYmBm5yUhlneEtGHIy6T0
hJXBG1fskObxFCvIlFSVRpk3FdsHAywtwLsUjGP4hW9ppAgV192bmagZuuaPEisr
/7vCL1i44pXxNKtnVrFJjm2rc3EDIdpdqexRo9AVPv2Vldz4wlNARJUYKAk87yW1
wqOMAbL3kdmtPexYRVBSdJuxrg9npH4zQp2K/lqkhlrp4/Qm0eeSBttpjI7t9ZBZ
BfQDL1G10oGCsibswpMLEALZC+GsD7bI5rLXpj38XUyvVRMKzYCpPkddVULeit6b
HgbMkgXEdXfmAIu4No4OYV7g2hbnuxc9DhcB+WobqBUS8t9+fiGKOvL4ln/32nGU
czw9iRnEWN3bWUB00e7naA7ej62dOLyxyLHuc3AbEJJ05h4u+gRQWe6EwlkJ7C1R
0KLPodDI6r6xoRkKE2WYY/ENURPGluSuDBboPdKxmLYzbmUUv1fE1WFw/hjXCOXZ
KJozbnuT1Od1DFE2LVNJVXR1TT5FD2lFqBDMDXsI0kXeWcIuNDVz4SUUccNyjTxF
kuPuJTdelVBRko+IYOlVhFdmeN+W9Sr3w/oyRm2Bu8VSGKml4JQhyBJpKRzbRMw6
5Jge0l4rHtfsfX+jpo/oYkG72sFBLYTEI2ccLXaiEeyp75Yk4z6GspJUR5vp2TYh
TJtFNJXUbPXzs5EiMqreJYTkkGv461Ou5DEhLpb+SDbvcLUQHblC6Dm2vDBhPLLw
eUNKxwB4ESUqMy6XwAFDAAnn/5QmjEdXqovQbUGM+T6XGSTso+JzC5Nl5ywcECNr
frM4sdy0k/G8ddikqetXq9vnxzFIcpLxJAaL6jHK5/98hE3aov7f/nGv/oELim3s
FunSDeBEMxWaVe18xjjipIlKnuT7KEA5TTsVLjDIqf3eowtjLWvCXiF50oqhXZLc
sJ0M7EfL0Vc58QtNQ9qzAVmxPr462wGollK6Lr9vz72D9Gw9QIRZhPTwDBQW73Zo
S9CXG8pxonfRZmjc1gMWtCaSHvXDyU2nqRirdo7FWXrQcYoKG/jW7MC9JORT/oYC
/sWkpvQGMSwZnN6gBaXxt0gYKIdpuCyKSnFrfhFwzruCew8eXFyReKhAQKP/FtgB
fQXT1iE+RS9IBzH1j7ffG/dT1crzIZt4goPnCINBgY0DmyaG/TrWyNP7ZScHuinb
8M/dTA9yG+u5/PGwYd/UXVS9cPlDYItQXSAluMtPj3TJTSqANj6QgXnXyl8T7cC/
j2qTbxtb4zetLN6dWZyErj6xJpvJY3umtTPp2tXHlr+2yMyQeTx/SKLUBP8WJdRK
S2lTj/pCAGReBxA97KfZZce5p9in/QxDiAgl96CMND5vTQX/OagAb0K361o6GXj/
SgkIey1nmYxK2ZcEBEjvz+yPlvqghT68GOCUtj1GunB6A4YEPEBbraNpaXofjnD6
c/gnrd5iwlF3kG6YcfixfgM0x2PxQ5SziQ2tJDOaRxLV0VhZ6DSgyUEtLy5RYBFJ
6ci0ILMilOBoj4D6SLxm58+8xV8aIGABvjUqXl/dNV1oCEiN7Iph9wpcTln9jXKr
0Y3USfPe4OphxElYZORUoMJKXV+w/PbVJmS9sRWQoy83MvZntzPcNpLQ9qCL2A/p
OyJ5czmPYNfjJr35ntS6Xw02NrycqYSYqorFeGqForaskTSZX+CQX+M4H+GmKd2m
NUMgJgSwJdDGX1LKGFa2sW+1Ztev+IDROQl55G6NDGsWClwsLfr1vPTipvQdT3tX
tMe3ArEaWdVDApvpY96138GetyINk59h9N3SevDlrFzS1LeepFbMoY0WtauHpnKF
BHrTyreIaTs+BQr2trDPpDEFPX1WLkcAiZtvAZacdj2edUV0mLlsVvWwI29CCKQw
3XlOiNuIYjYYYKJjqJurxkx6SY2rTAAHlUp0Ooxb4+ziNK4W+gXmOxbCebz5XGG7
AAHT1nwqzSk+uU7boeTSKDOw0NJwqamiWCeqbRMJ+VUtGrqjDxaqW4F+6wqzz93D
/2DApxSdbB1aDso8tJInHEEaArrvcJHAJQ6hAelghn8wSvde7jmhCluYHgPQixAK
0OoQ5WsHUcD5VwB2C1mZaRawid7Gd2pL4ymFaOF46KMRGL2/eqjB5Lhwb1nroxU7
NnD1QMt/V18OYRqHP6/usOZNv+kiuROGax/e1bAZw1kvrgVGEX26TQr6UmeCMlp4
804Hg+xwugz6KWV9vXkwVFy2/rOCsstyApNe+VCekhbuZmcCscdo3pROa0jreM+l
xqkr0soX5yYxttkqVC3kap3ocQBmnyCCsfvrCbgOb0BgO5lN6jvDifKJc6kxoS04
QGmXVrMOG7OG07ngkxHs0XgCanUPR907i2hZvWm4EAMnoORWTLtj+SwtyXoGoYC0
W8UDxg0IdBPmdalfdb0fB5kSpVxRlXjYOWHM+AEBb8WfFuFbKAhVBZyHex9KzS/F
omy4Go6aU+COuPS3r2uAWSy3jGKYut7rvvEDtXMyvw/usQWn3qXprMdMvnKcwpTK
aHx9uoIfkMAkEx2Vt/JacweLtEaPQbBkS3WxH4oqip4YGZ9oTinbo+sR18VdW03Z
tj7r8JxocqsRV9dLltjXzqNXDYbW4stHcvHG0VxVGAq2Rye9GX9N0MrL6ZxCM6/8
VGtgmhfqPBzRwodtBPhhwkJ2sCztREtfmGeFf3XzieG7hv0UkPF/CYaO1u46wiUq
BVAgVJ2vkghnCnqylVhGN27DMnRTVYHqiR48EsnHEeaiqIjEd4aQOE9M34UuZvyr
o5Jgm5fnTWwYLMFvt33VmmnYHSW7MY+pXcBrS60qkI2p3jSjFTuhjBbe4hPyvUA4
IetonuVYXXXPFVWJdC8iz6GrEuzEK0k04A794bwXVh83D3b5DT77U+6EySSO4o/H
bNUIxSsVB0mw8BCMCQbs5SpgOyJdfYjdosD3Ps5fnJrjQkQSo2yJSwpsKWYYU91H
5+m5GBFriUU+QKE1hYBNX1kSTZ7o1mE+m8AVstIqESXt087dql6wde2rgqXpaNJ9
JECHL9W8Op8uw62zW0O80GRCTn4qCGTFsXsCqE08LNu7V+4MpRziMwF7mASTVrJg
Ge9waxZY38QfQgROMgEaBxcIh2MlXKpvYrZswltzFTp79YEl++RcCOTSmI+rqQ1d
UF/9gywLTbxWgWKZOGoATx3SKbi0WfE+q1e4ZLNEiZENIPDx1Pqutp4NWmqU/Bo4
PXymV/QCYohQGk2gYj6Cg1mjf1R5THDLv+dWrdKplBbmHVyCSgK2DIpwvU3QuyCg
AlTCl8y2fooRj6lP6suxxuRSrMLiUxBb1WsJdEQlTZ5VzTTr5/25FtIueBSryg1q
qHb/kz/y5vUj0RsAzNEib+IAuQucKPUNSHljZYgCzFHU2W3Xy4d7POs0bCmNg75R
lwTwVbCCPGMm1Qz3Uk4kJtcjR+ESlAWiWMUvX4QNLVFlfNUXeYL1e4UuJJdAdsJG
0EZreIf5cGEKdYYxn3bb3CxATCJeBK3pDw5TLgNPrjDgaNePqwTE5drn+QTs66ib
P8H2sbOEcxqJcVNK0eSCVsF02TufngyinQiNOJvDnG5WhGD2+nXnPLudr2nj/cIt
mOiL58tdeVwVz3Vcf62uyKjPvkGB/CMAf5hGSDgei1piBPmgan53prnvpXcdQZnd
NOB9LvcZHw578MOVc8Wtsg8PC+A3UyLk7/SzIca2ixrr1/upiHuDiMUZ/aFSdxNJ
JvsAphANBEYRKtVYiTdhIG4e2MK3bFwLnlXcgjmOyPsGNlVutk+/J4tqbvkrPWmX
GrWnalyAEY0xiLeFZOb8u94ip3hNSi9h2dcbuG+b50UURG1r55LXAeGNXWiJzI0v
Na+TSig0jApuy9dqXMkjpRP1LMvuu1OTfEESjmTQHfX5e5+1xjxfVIl9P/FV+DtD
7ipZaHFv0qw0QcykhfV9+eWd20lEgcWOKwamxxoS7M3XoRftDgAw9m3/8zLkAJmv
nWLOxsPYbF8agXK2UnAVSre0DEpQtPRgY63KYmMhliiJ3LignRjzA3agekCJ0Fp8
4rdfYWqP81wXUcQcyluaZn2pVtcczDvT8NykwegO3v1E5BfAbwQnW3KcQBvihrOK
di8/aui+TRo+Fmb/qguAORhZJUQQOhFVuGDCNc5EksdHynos+jYeXXpcTjYrFhpi
1N7dsJVy9IdQY3uKt4Y8p7Wfh2FeROI4M700vBAH0SrPewxFliuMcWZ38wHLYFZE
/F770yKTnhOlEb04t+J/ymzE5C/LgR390STlr401UHO4kmQt3ZQHQzuwRbN4q30D
FLvOhVdDNoNzbgr2eeBOO5E/ZDMP/412z/lMZU0/dsi9jWNTsWhao3lUSp3UPDNs
gMcP38JdjR9FZ0auKKaYzjnN4CunWrG1XsvinqDDfqFgpy720aWUMLxvoEhTLi37
gXRmUzKfXjbCWMAqWbqcFvNa6ee/uRICZbQQzUPvYBJaYMC2dU1OHlsV5BqmZm5F
SI9DJ22Sj6rmmJNkjdXmGB+Ke4VTeB00YMYkFUT0TQD6/9albUkv6XtedDGNUTp/
lCFeU31J+FEa8hyOh6gvn26MOZI41ZrJCu7O8lMk53dndQ+RMamKSmUzrYPEp67R
ZlfO8ekRkosTQGFuBXrIVFxiU+5Zort/4Nip3//86CNUkV1fFwFJ/Yhok4C0/Zf5
RGYBpmuNoUhW36HmDyfzi9VUSSZ2kEeVM6rfJu4RrzjIKiaC/wf/QDOchOAdYUJJ
LVxX37ZsAolCTd/l5kJNAGYeKcYG3GdoHZjH3jQ6/6boCnqkAFOdBB+9zetxtCSK
9updqDPip9TfA2esZG0BBjdxvee7cdLPWrBLxFKXeDgxkkGm6uBLzlwKxZelyC+l
yIDMAwWTXftlKUQAE9zyBd2fqUqSgGSjikGisJB3xQfmJ9Ufm48+v9cOgPBGZ4CI
DRf+7rAD4A7BMyhKQbjviQbK//hfTarhym+a4kXw7mmm/rPPBgtu6AM/glQmeOWx
5JyqzQk/8aVYxefGuosSVdqb92bPKUSO6Tr2NFJIil83EqPQaKKOYC1O5b+P82G2
OlNtR4/zIkn/uCs5arG8HE/P4apywUE4Z6aQGaea5MKUhEYjK0zRWhCxHMluVyev
xwwRxJD9fnrMYcA0pfqfBj5QCJdtLC6A20sxEqKUv2cK4zdgSn97k1kteC4yO5u5
1r0mzKlOhLxR+KFihzzDVoLIG5XRi8zflQ6vxvYxPhYWqcMZdOsBWljyk6+kt0Li
YECS/7OtOr/RMGeJGf5Yf8GZhoXYI6PRpUxB0y+7lMTEc3OYDcnyfnhTnlbhBi3J
vbaypJztjkIyxELppEq6XGD9tHo89QWa0b8aRKcFFln2j4Gom0oner4hK8rSMrOr
kV/g1q8wREdQ0sv3iEe6ezuvSzoS4puraBgje7BEGuESGH6q3AJNVzNvdMmD58VB
IZmoQh+ueLjBTz2t0olC1/6k5qM8qXH2h18U/YeX6D3WqUki/4ZHCuyf6GOQOBBM
zyfWJyYdAtzt0huNgyEpuSlTeTyQGPpwXdelCJrdboo7uwgmRWBfSFBlMUdqhJKf
jQQiqqa0Ij5VwcbSyorgKNhPxbKlfUORGidLV3m0y321Lad/U1gzXpbuMNDYYy+x
XN5jZWtaECfZ/7j6Jl/WX3S5r3GmvDjcIJSu20KhAL0gfrblb8nBz1y/CgI5n7I/
mNDbSyZ9uqnP9HYNMcHd8qyme6jd2qliyCcMUQw8H70MEOSIB17c31/gzPo4eRsM
q6Q23FfzYjXG5BODIzXnKDYuVZMxAfG8d3NGziRoK4aaW8mCHXW8oszhr6gOOXw+
eW9xwY99oKVf5alGnPvejFc1JlWylbL9DmHTzjnxjlIyMelEbsUr3GuX0kjwgIFU
IfU0+NE0PJrdJ6wNAG80XMg4qwJQfbw6OSqWzjBVYjfg8ApSLSDmMzN4KXvzXVh7
LfdcKIaCQBtrzK13zw9bQOWMLjhNxroqN5yfzS15bOcm9yPFn6wMOD+qRTqKYn/+
9PduKPjms8wQbFLbC8Pg927cKoKt/bZc6cDBAcVUWDNFlBCARVZQBRjuwByaegc8
KrRoI5ODd60qATt1VuwkT3fOa/EojEm11jpJ0fymDmqQHPOKjjmYmBw2E/FxVdgr
a8HSSC7GvVr/QXttOQcbpNwueQ4JWzxoDw/2ps8WfXNPanEdxc2/rwaBWFUwCXCA
f10CNdfRibz+u02LryCPxYPjzfBw0UoF1QJzDBiNJvbSTPD4E6pCocunY4tz5+3l
/gY+k0FKub7AfLEOAVQvY2vAjp/rt2cAnvmmeNXMsn94jWNrARsdqrKqBhkWcJcE
UD3mclzOaN1pYnTrRpeSV2WksugGQzUEGbc5fHcORJgZ5sWe64NLYl+GxPXHU6wC
l/JbrpkeX1hXhWbR4dmBw2Uc+2G2/vAN2GWcy+5w4mrTLtdh6gG36eSmyHicTbIm
YROdpYFRv+R7DDPAwZuk4JS0iBK6Vo/A8ROeGyS8jLqCTD6mAk6hpWlu7FrmPwmS
YZnJc8JZnNXBViThdz8oahfgFJcDvdI5tkJV3UHNvzjL04huqJZvRhUzUihewgTh
7DT+ragsZg4/92MTWf+7BGKk1cC45H6+NtX+9IjbQLEItIqrW4c6Ty26cBZocHKU
2EfB0YxGlK6xCa4jKzlRM7RuWZ0mz1MlYe3yV2Er1VnZ+XCEiKcZWqmJcEH7rCAQ
ahfuvRtI4513LvtfXUKhuKSSjiIpjXP8cgU84B4Z1quKl0bPo+hZN2BKpaJQPgMb
vln+zHoPZYHQ0OQYBQtbnkZNREkPAbcfdlsZyVMug4l4Mf+SHS6bd7kiCxs11+P5
r8kiUX7gd/T8M/EuzW0mnwb7vAI1PcFVSs4Bg+K66sTZyGs6gzGwLYfMrXjOrWtq
FKzPn3/nG8pRs0prPzMyy88cZwsrgeveShAtYieXiJnZvnCljmBGCJF8YIXFqKkU
fAYZhI6Ys8wXfqhD4rTh0fKONdHdrcdDV372gjOF/NNEWOCGkoFXlkD8bnGOgJUL
gJg9IFnkFj9VHk9nNqxIBSkTFKurV+71c9ucYlQm/WTwNP0nX//JsNa4pBLeSEnt
XSty12UMWbwjkmJzAeHYgkoTlY0L/ReAIMfGpVwF8kzqcbKS18KzGeGYOsxkAEKu
+HR4mjg7uc58uH3Va3nU3FHvWQG+cmZIWqczJOK8AM44p01xjih4ijaIH4YpyBQ4
t/CfHk3+oF6Jv72sWlcYpAV8/UxTaGjzfEK0u2OvFgABOGDrpE0EyuzBRYhuksMR
nJt5M5CFQ1huYgZJjmuRXEKXZ6y8RbsHbSwy/Lqpo9DQWMGX2rJDRuQr8sBDNQba
2zKdftk9vi6TtyyZ6WsDHXB+TkZGkipAd9vchAzS6TobSYR8kuq6L7muNEqNOPiB
n4niTU9vU92Y7cuuAfvUOHDurbR6Ox1J+kTho930hjGMYs1mgA2AR/of8dzbAdAh
jBlixXBVls70domGEP5kZJ7oslV5xbSEAKSx70vk62CODAm/tnnY0Eb4fDruHcgz
sp3exdjG7/wf8bxNAp2mJmDsEvIZZJX7drXDIWCwYPgU0GxWj0+yjN2L97uPBBWW
IcyqCpGvcLla95lqm8s2bZvxb7Mlm6TAe57diGDKd82kwmWiT9lSk3PrNlCvEehm
ufFZ9sxE8qvjPKs/rwbAJ1GzHzt51q1IuxUy/+xDRP3CU6H+zaUc6PF4h6P4kp1H
ZBmO/KNasPKkmVEt01aZ0tTojXNFozFXBwG6cIuXR7ODd4guchpRIlW3dnrW5QC1
O/Fb9stdxK47IFjCFhRmyO22vXwcXaN2VTKpb2uQswT/8zIwX6tMIXTjQKLSF910
LCyBN+EAWRD3hi+vucA3xXeYy51iriZ32jfROckTgUhTGNL++xxnryjAIyNw4lI/
ny965oANLZ8XOKEo9YgcWSfag2rBFnE321F/ksMAVy4B6eJOIz0UUdU7SgYJqoRr
H7l+bCVu5MiOr2DiSq/RzPryz8wZdrdE7PNq7A0G1Po68MWb+dT5EcJWLP2/IVbe
MFDLzN9IKuYA8iPXhiR47XS0Lat00Gfb1W0w4FTmboCR+MUNsbLz96YgHRibwngg
QbHpR8dBre6vYM3L8LuwxfYQk7UFeENM9DmKncrERE98MgRCJt565o792UQMHKKI
Um3/O17wIiD4jxMqsDGQsnHymN8TRai5DUQhESmXd5SZAmZ/iGLZpRXZza8D2rrg
UoyU7/rmY1z/Je9SrQOo8NR9sKPSGdtNHnZrbCmhkxpUg8RN4jgCYYkaTkr83+o8
37Ww8swvXw80DDh0s3yfcy7scG7PoVzaXj9JVK2zE5ACFPMRmX0ncp56QewHgMY6
V7uEZmr84t6wtrd7eETCdX08Qk3KtNohzj73JAAky/1ppejhGuFG5et+ps3R4haG
hBU2dvmYzSnxCoVlIQ2ak2yYoqOntHLaXfYuUFUKhekxL8rUDAabrkjuXpujktfQ
GLu54+Q8wyttn3IP+gUQVpYaVM7hnE+DZvTVFxl1R5bh2Jt+1jSrGE9FHruesmiF
gn1avzh3Gv6oND3ODJCxFWeg+0mfmQJ4ZlJ7oY/lYZK3U9yitca4fWutnzuJv7BY
6RasTqKk9yZjoWfbBGcFnAR4cSqOb7zYl9QFwWtQE5AfV07OH76xblOGHWSfI4rw
2kX5BVK41FNxx2YNQQqy825H22H7bdbJMWXOXNAlONgAToWenjjtfARqdxNem5HR
II21GVunSY8Jfr2KPND1y8MMl8UT0C3wJIZrPu/dOQ6T9nLCA4gMoR3C7tE63vOQ
CEnu4wzQ9wUfUzz1/KrFTngPer6cEFlLtAvPi404hyl7CZ7EzRHXb2w1UevMkKk3
l5R2HSq8yLcU+G6Kx+RllcRIfbC8GyoQOmZvZeRh7lfLlOHEtz8w/34i0zFdm9nu
87+qSqXTNQU01amTNdfdmDWV+5uh4yte8NPajxsDQ6ZHFsNvogsZw2FS39zCZ1a5
Oy6Jmjj8P3rdvgQz7d1+suz5dyAqCDcucfL3Z9pZWdlMVwTdkciqs3kA4BMDVUNP
BKnU72XVvYjTu1mQ8k5nRU8Di7+haZpIyIZaMCiz+Vx0TrpOpYaQUr150jWwLTg3
54NVmdwQ8NHvxEzCzBPO8lI/A/7oDnF9viszyi+Aq5X2OLd1Kd8c6q+4vnCSVmq9
wlpMBeHYIfQTZgMgWffsBHtWnC5i8nOEpxyzcRx4SrWsfJ7GHK4lkWYivaooJ3ts
AeuKm4SVRCDxnbeoQ5KAV0COLiRtHkAHf9ID1neaSzms/1KoC3tMT1BTS67npe1X
qWppRIQoDTpD/+6UC8gyTUKFCV5DmuOnHrV9AC01f7BZpbsS4Uxfr8ugey+x03k5
vAGHf7BIg3BE+HexsIhdisoD1iYPVjVxwH8D/JXDJFIsdYvGel6h8vR/E5a8mtxi
JskqP5meuuAc10F5ARyDN4b282N87WmoORCWPDygOXLntiaTuYgWkCRUb00/HSyF
85cCtbkF6KpKZFJ4y7G1y+8popRlOAWXXkfrE5D1+UuTrd2K+MnaNcvD1SZmi9JD
SQeeocfL9ly4tc0RTALaRAqkZLoqbQEihxj1bBkku8XIdrUsDR11C5XLmwKW4ULs
99oG13usQeCSY3MPS6GJ8IvxZNlF3Lcd6SBA6GwMaFs/MbQvMXq1UYJACcfcSgbb
3Mp+e0clEGw/o6e0Dh4Yv6Ih25k2D2i3cd/D3IjbwALcDEuiifOARKYjOlF7dJyO
6d2Q5KjeutmWoSKbmRu+OgWCkMSXf1mVlig6htkI6IKbW51eHxVevikJVFMidu6+
6XR1x/RFT5HOGl0NKOy91WVVtBNGo/xbfTq1/onhsWfIN9UDzwFC+4I4r5SFgNsi
sGwlxkIT7L6xA4z6TQD9i6MSJn38m0yqn+PxW9hmSklqXLSniKlgxQ+jrcy+kSKC
/OiMPP69vEHMbBPtTSixzpLjAKM44BmRd0ISKpTt6thPPMADUCvUHOrPGeUpDQ3W
FPEl4KCbuDsPAqtuOWON6bQGjRnJYjbqqckJ3FBe2hskUh0cFRnRBHAcB6R3G7ei
d2vwq0DXabYbYUXSTDFJl4catic1KhnTtQwyWwbVpIELcMsKxCkVEJk/U+jzVWGH
CmALX+k8ZJerz6qefYkS7oOXpWd6v35W1sH60QhBlIfDz1hfPAj1V6HadFmbw+Bf
R5c9fxbd8pxu9oZBbzMk90H+nlsb6FYJ/K0I18xgZICVi8OF3zawPLwxEF4QY3JF
tZhIuKnnnC8elqFw7ubroBgBUV2dSEcqdtrtUDWWOHJ4of4Gk6Dke/ZIdDYsPT6V
tKfl6Vjj47cO/Vhl5UugVg25H36Wr7zrf8b9OP/qpFruAUkMFNcAZu4i+PephCdg
p+R9luOlMGpkcSpoUbmMT5D9LJmdBilBF3Hb2LH2kOXYyXCfdEphzo/o4VZhtdx6
J8ij+ArlARY+d2DI6NaKRKsuxmjZQQv5bgcg72eRB1xvIeT92yW3ihJmU8QOQMI7
knG/9zsiTpFgMP42phS9yw+TavTaRdaX7v6wF8Sz+YOv9QLYFCkwnolTWdGkIEJt
Vacf/Iv/8ntCyQQlO9auiN6Mwyadzr+nt67PwJkFwGoKGTpgnrq+1SueVwrw9kHq
SWEWpAXGKlhhswwmmce9LNVLV4V5342Am1X3SVnoHmrPesTAaczLfmhO5I6bSPtE
XdGfkr4/TSNmqZ9qr17sLRTZmFm6IubelwTBdFJ3N33/Tm1VJFDYtmB3PlIt44s7
c9zaYWNSs5bhuyFu+tnt8qipiXDEIBK/yPzzU0JC9CYVzL5lGMSbf8wZr8IifNTc
mKQuV3AX843a8+eMlug3jAw5otxoEmKjyGKmv34Wn83WMGmsepbe2+zVOAGTw06s
qdDNlJ68cZIdiLiN58DUvkYSFPCOLfsesHDOGpO+YCJ1Q54c+mcCLJhKEj+5w+7j
qNQx3FcbBe8pKBn3U0XMVDfI+2hfu3LEQ2DioMXO3I1ktzusvrMTNfSeK4YDkCrP
Cy4e8+zyIQu4w1VeTwvdWXXpZnN4an/fAunJUjKnUhxuUWIisaMrsQwjf7BxY9NE
edtz+WrNIFbGCtshM0jfBc6sglzYsQNWBPkTRromRlPFcFVIFgDUJBvwCQb06B09
brldXAfu2Z1OFMPC9jfQeGPCZWMOsBnYPiwvjD9Hy1z4nUJUNq02s+4YjAhPT5nE
+twIHUq62BYH40wYAPy0w8fLUCSRiJ+DhpADrd1xG7CZXAAuIjwlthzVCTOIxeh3
PqhY0bQJD0u21PnqwB62W+2LWHINWNMhB1Ii5XcecMYE85Al6fpLxRREpoLnza5Q
wtqsFgKF+YABJAlU5bG01X92ILyTBPFblBXEsnJlW0sGDEkSvcLeEdleFMB/TmsT
9SQlIdQyKAPNM6tbtyGuN6bl2b6Ps5D5gppSqdR0dzE=
`protect END_PROTECTED
