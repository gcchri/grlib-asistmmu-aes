`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dhBpS362ZKko4+2zSWbdZ6imG3BBj2fYjCrs3vA4TGGjyyKudP5UdtqMmp19KfSi
H7u4PZUBEDwGWAqQ9ZMekVLOGSxzIWF5UMQmjtEudCnKAeU/ff8faCqH3osviz9G
RycHiHmCvZsTXfxcHuClJi8udiPAaBsUUlrmaL0Qm84YnVpp9msnnVT1UMOVRDIC
GREzNyjR2E90nLWUD/FpXQz9Z5Bg56Dyvqk6G4DJyKEpto6NgbCUKQJWZU9Paq7w
j3wVXF0FkpWWDoU/S4txLdvPJ+FdNbrUtVouOqND+3uR2NQx9UlLmR5WiFJ2spBr
MYhGu/PKiM7AdHdHdSAC8j323/3O9asjcpaAOlWq3l21ToNwZ+ck//VuGLlHP5Ys
dvNvEY3EmI1tGiFm2FzS971CIAAYV5uIjE8zA3q0VOzL37A8LUcxxkcrgb7PTg9i
MLcEdh7t1Y4liqx+ZyPzhqVVwK4wFgm0b7FGt06oK8P88+huDruk4gHHYn2hUYkr
+KEkzEqv1XVNyQItZn8Y25xamISEPUaFKijHxtGy6lEajyehAfRzkvb7F9VzQ1Qp
TFqHc9ejk2u3CPM84UHxeA==
`protect END_PROTECTED
