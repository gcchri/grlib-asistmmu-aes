`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9All9hRowY4TRHdALzsoXk63jJrEWDJMzQ4BzHsRmTeG4JkQbuAmHvdcWGf1kjYN
Pk9Vfm3L6M15wLn/h22g/Gs5qk6gS3GJp/drNEgD4o5xLa39iRlDEO2BS2lt844G
fCZF5EwUQmBDWUuTLYz0OXSDehCrpA3sJQgaVfob68Z/YpJ+w4FmErREON5OEax7
9H753/UD0zurbDeEriAGSob9ltz+5Ixn+taqXkU0if2xrZWwD6Ny3A/527Knqu7g
A3s3bmV74GHZYecxBB2oOgBxAOXXG9KvuVXPPx9qO/LQ2z7BqSpYsRvRKSTD+vt3
SI99PzKOW2GspDuEDEcn/NFlHiF2dMKEUvZEHYWcUxTsnaxvz8w4ERM38lpczNYu
3CFIlaukrId8Iypi272celHTVHuScjHGV6HsASeqCndtMHhUZUJbVRWTb0bGxvDF
vGbOFIH7PUUk2zke7L6IV+1YENE7o2PaUaU+3KTZPyM6B/4mY4Rhn5AJnuZjYbyi
YJ8sVQ6q2khuqqE5kxr1xnwqMGX0Er2SN/IceK2WwUnqbxWYekNlnc6WK6Kkw7Tf
sZFyZAXp8WSE/M1KKFFOrNHr3yZKj77uaYp12Iv61RPQvwrJnNUBAoGYk/I8wkx5
zT+uEKa4p7F3preNUKzRQjSIa5Q+DlJ2HYCDx13dvXTAXKBVNU2LlX2EJ+xBM1bV
ipyJ9U8SPXKEs0+/4dlB9sS1YfULjmJyuj+L2w7mPM0N4GGWZ4f0yINcPH3zFNOC
lup9snKGtBENQzweGUhyiQ==
`protect END_PROTECTED
