`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tOmKuWWRMb2BTiMIvLmc/nPULJNCrj1kfRAGyBwTeI7v1zFLcEZgq3xtdjdUQIup
Z1CzyKf3cC+nhYKU7IKSnP//3ex1oMoamcxh47/oaaISRO1M3uQ3FCq8KUEhcTV7
vvKTnCyI6YV+nO+4yTqAIwq9Kd4LWmmkEi+8Khl9VjHEbkuBZC+wHaHPaGXPZRUx
yRnYO1cD2fw6PUcYRjZRvKdNDg1Y7DNC0Q3dAExuIKNDAch6i6SalfmLtKxILFkA
/yo3Ru9ylKVYsJR+pWHv/dBFTDOfaltfpa6gD0JCUWwZCb/gx9CxOAVn9khXGeLv
UcMTvimQnViiUho5Qv5dSfKRdNdndfYRUPZxTB/VXqQf0QbJrObzYc/adzF6qIUk
bV5b0B1bGYl7XOgy0DXt1DLCD/eUp6kdYb0mrpNSBS1rI6b0LgDdQP7bxYnHopN1
xqyNOz7X1cHsK2zmbquZI5g7krDN+WDGpWMU04AMeUcpufcBzY95ROgmy9J28q1N
9/WXlA1QT0AnExRfE/Dc7uYk0qMtFQey6dAMvvSpd4fF7qnQ76llzg3fuvKw7Nyr
gHVYpXANNZ73Cj2dpzyQ9sUWAH4jWq0or4TUsbfyU9m0q5YXeEpIXiaF/P/mjF/p
EPnyHTbRVP1tYXCZrn5OmD7Clb6WJlsDsxyChx6WY7v4B27drbChK3NapHTWZONc
5MjD5fpqiDVz2gPae5EMWNiFD4ESIa9R01iLj8r8usqA3gJzubCGfPkhTVG6hLcT
kbIlRMoVUj+9YnEv+/0U/L1+f4NTS4JGbQ4olVtnaQ/KrKDnIiGEy/0aPU/JkTNr
lZN7/dbTM7RqFV4Q/J3oJ876DvSFxwumINNO+GiYruVkyd0kn1klgAkjY6zOJuEv
/wEo0ElLfuFBEjKogE7q5QATCg6PhUyI41UgI44dbVRSrzPt9KTMpsHlO+CAph3K
5vTUIkq/QLYLpppxU+YtZie8turs+ucdmscUPSHuAr1JiuBQJcWIQ5vKqHm+JHQD
/03U120xgvm3R0DYIi/AQ6c4u08Xln4EcknHHx4L+06qxLlSNJopo0Xg3q5mC1fJ
AXL7xZnoCfxpVHp6++N1mz0kUP8cNIQz7PZyILedapQuYDmhaYVVoL8yneaYBV0p
etzTfgaCrD7az1TVh/lud9e6ZM1wRr0xo9zrWDlWE1fDDxJYiidXX42DvNBGK72b
fZJiM9Xu3wna9EKuYPXgqlsdWuHZGhrbwEqlyFthrt54fsP4Mkf/zLfGg1Gqhsc9
Jt4Ck6u7Z+/7XZL0+coYfrP6gyzJK92ZuRb/6ZWE952Ub2Dpz2Zx8IgssT50VG2D
MQgQkHnbXkaVfb6A3Jm0ynMzJk0OzMSjT2DN5bpVB4Lbj6sn97NY2Zq6FBImsRHi
QkMLEsjfPCgwaunsi7E+OACfl7DjFh5N6mOsMvamEIO5RWfhpkMTUl6t+f7qq5vt
egom/zfk3jtdTkOMRwlDweN2MHUvf3dgJrRlrqeU8WSVYgMP/4fBApnbjfzwBhsl
WZg4LXmOph+0Y6xXiP3KudznDmZVbKCQ932srHyaOTTZSqmpV7ZKdbB+92A7bu2Z
diknaZuXvKYSX/vq9qWr+T7+Pl2i6hGsKLcrBJ57d6kpUtXVoiJnWq6t7h9E01hX
DaR6gIQl4+GfHzg75Fx2EIVgD+B3WSRuyBHhSoLzPWH4BtTdwuSP5SsBY3i+R8Dy
7uauoHNhfdxW0GYpz0hyg00IqojD+XBacxRHyK/EPMjTUmrw1ZZ8/y+wVI14Fa0V
JRtasbnIF0OJLF6WzJafAHhoyBoM++g1jrmSk+kU1D79aE/+QFzSzfLQJNOzjs7m
PiXtowRylQr+V4rDgU2rXJ7d72UDjjXpge8YqqIwdtg59Zw6IGel0uoiOfgMgu/y
IfE8LkefRlKpRb/3JC++qVa6Dbl3td4+LXYmspaHAqdV+tTBcand3FjKhrJMcGo+
+aPWxksybl6npGhoEoW/TlpUlDMX4KzG7wjOq7IAW690SowCwJ6b2DWK+98ecMkl
meJ3qYWmi2CFXsVPrATwrFLUkPxm/0tqVpiJYe0nl5vfStGdJMYVJSd2pH4q6bCf
k24dWn5MiQHSOrffhcdnZ/kZbrzHJnXbhtrra00AmVAwCXgWIjYQzWhnOIgcRaF0
1guZhlONjneWmh8M8PsxzW4MG4V4ZplafQ8PIDPe+0eOf8UgXF/C6lI033Jb3n17
kHADSJCfXdptENv5JKgeAbK6PvaBaiQ5rLvEnC5O9I5U2nLf7V5Yna7P4ubuEH2Q
y2qjQ4lKnbV3F/1QnYCOlOXn1o6vH2FG+KzGO1ms+hQ92H4uQRDfrcHrT+zR4x94
p49pB7BZf7rw2oIkVN9jqCN6zK4t0sSSqvGimK/g2lc0wsbxhlem1XCdsIoNibBD
HtAxynRHb35tSFLne1ZtMnQANvJc9OY6iXLUiDLFOy09N37uC5iIadrPcAVJ5FYq
mnVoSmwGt2vyF1f9KSGOp22u2jvgvp3tbQPAWJyYUR7tdIQsh/N4sTV+Zir1fjQG
FgeWeESiGGxEPdN3LkBzTiLJEyC1Nk8uxGV6xxvsQ74fgn1zfDJTB4KfR2R6bz6w
9mizkKlC6a495FgI9614XFZhppuW9trbYpxw145Xzjymi8hcYn16qtryCqfgfZ4b
anFIrB9lipzpo0EopQFHPwlp/jW/l0DWziqC07QK8lZpfAKrBNM5biE6jywZY/K3
oK7dQNCdVeDWexUbFGLZPoKUih33jf+hiwd2I5j+5X7bWQnTcJl0aELd0Tq0cTXG
yj56v/Ahjdbt+2XFioJ2dkhDpwzOYMhXfV34OaXLveeXoThFABxeQOzwThmvptON
57g0nuN80PnZRwame5tvufWUvWaO3RG4twM6NCLCQ9zXVNEAIt2owNbadd89UXU1
x/vReLF4Tr7JWgEbP3VabJ+1Dry4+dt6dJ5+rbHwsrl+b/hdG3y+5CSs3xTRtUTk
Z43jfUA9hmxkk2Hku/Dg4e4vtsBVgBdlapX7UIJ8lBKeg3YFP8peSgO4yCb3aw/l
sIq/PA9Skj5epza4QBlPTlyOHt9gTri4pGriITOymykOkF0fUK7qXFINUoDU8Z9N
w6oduRZzkfJxOfJxNGQm6rf86OPT0F5Fv9mG6ey6peH3lOL2jxTTN1kfE0nSs5fh
FK1MMkkuZh9izCldwsXsjmsYbCRsv5JRieXpT5YyNgs8NVmSCMjIMsLmNCcLiZUH
JC1u5Bw9x2z6Mrji1A/Nl3bC7mVDW5CcZAHM1z1xxhFmmOPhM5AY2FJToSBwBdbK
Z7erRXHRALwy9+rvJLfY8oE6XEe6l7SNNmP1gjq2CmVRPgGQ1L7kCsl4fT9JfbAR
z9lPXQsCvJs3Fx4PI61EeVeaQ24xI0ZnzpjJg4NlbN6MzoTx8S2z5BHje9AeOjTI
CARw/Oxb3PdJNnG2AIlNN0n/pgvtTrhJJKQhSWTDf48K7eEuUk/FVmKJ+KzjK0R3
YPE/ZakQrCQ0fsdpIdKF4L0vklRlWxW/z6xiL0Kv1z9Z7DUNJVxL+2mrGawJEa3u
Eq31y243Jtk4D5NGwzKTS97QCuLJe2vi17ifs2ZdrCj+6a4hWDEVQN/MJoSv/9W8
9oJP35FF7BbTh7HEQegqGk6uSU3qEsfAYTL5z5pe9opJUCF84pTZV+LKjWw3oM36
VDJyd+ryNt2wol2tBjO1NTTS5rvpaZmD/bG/vz2A8xblQSlRQkqpTZ1zv3IueCBc
KEdbBLVQsngtVwYDicMvtLvwtqgw9kBfX+e/e1a1KawjYZN/JV8hhZ3gODozA8j9
hmofbWwS3Grs/I5j+IU4VdvdqCU2cOSqsm82pInkLQoq21dPZTLAJ/+YiFSOztND
Tw6ABrwg1SCZyQD1zMqKfFIVqp4kEAjQZwoGhk2fLJ8ZN65ykWruB9M98faLpY00
VRmX71QtAzDEH9+O5sO8nEZo0B4BJTVMUEfJHZZXGiOamBeSgRkZ3okbgdtb3SiG
i4TnX+moICPCcrOjueMcDsM/NR3segxHbLMIbGT8CgNvORBkS5b1UoZx66qlnZr2
x9vHM7KSG3wg+E0HP6p04atqB5h+rfNdrwGXYEsD+glT06lvmCKNqN/Iy8F4pJmV
rtkCXv0SrO2CRbC/TtkVkzAEUar60eEjaJz4sugnYpMW3fn5GU7PDF+Kqxj/+OQN
4kfKHEkBxfYMBRSWbFoB2Z0Lop6l61Z3atc5jjhzjX5Q7GolzoOxEDYXGTR0op+5
P6z6hUgduDihUOQnqjh0E3fBPbt6qfepPNt9Ghi3IJab/xH3Jc8Uy7UTKihmPo13
2D0HCmscdv6zj3oweUIGzRKvL3JR4nR3fds+m/askIzSEkGVVKqsKmdoy4BYCUFf
KJREVwRllCVcthWARNxrRRI4jz68znKM4auv+RXTXoEiYJ2XIcycEyQNBOJmf4+M
L+LWkAs73flmREtYlGPxRQqNFKIdPj+x/gHWOWNbyvELwZhoBN/in2BomuPr/1/a
vR8P4rD4MjgYzsqFMTs+SBFOQ8iKUN5vhUYasUrY2T2sDEUnHOEsmR9NQW1uJgQx
H1RT5nU1Cjl03f5APWt5zhBkYuN2LetHZTX5N1ypCEgdz/jEg4dW+jsMo7rW3HPb
kjdZtnNHyY/yS3o+l/OuoyNkBYecPtVqSMkyZw/YpO68nf+T1Ji1r1RtA71RwAN9
RVFInzUu8sCI6CB8OPdMf83qVcy9Jmqgi7iMcF2TDMpN1IkIL6/Umgj+hZ8fM6qj
Mjb0liFnXGVFWL1HX3pE3Vb92l8pESfDRSfbfmki60tHRPveEN3WKQy0lLSqzi9F
A2vo0hDWJ4SJ8ZOJT58bzCureqP6pSymdVLElrys2DtQmarnTO9C4Vuo9x2LGCMF
TQfm/IzVWKkdPpoPE+IFmeJTxm3z0Aid77Dyv25oLuDsVUk7cyz+Bym1qlu/Q4Sq
D1SuZRcgctB9t5SGnVo/aETnbvOJ1SKufBdsiQNp6NFG7aulmo3SGcsgHz5wSoDy
DieQllqfHEOoJOHZIEn5PZfS7tL7IaYxbjg7B0r1dyUrm6vwH/GxqYVyGdbJufQh
jHrL55aN1e9u0FsIcA3A1GlL1pptqtoKtYWnuqmpTRs50eJkbT9strQ+XYMGbV1D
76WVfWKS423Hz9Yich4+KmMA2XwuSvrWmUIN0WySoArULKLje8J3v0RDmxek5Lry
Co1ETL7iNIsEeLXMs5cngYninJxTQBT8oU1XJkY8ZQ+q3cevsOm8BgILsWC+cLhj
EKs4w1VmfGijAkKZxa7tALYpZx9Z5SE9YCjMbmjYiGQW3DLCwuoKnGjiJq6aXuzG
d/hAIOIwoX+DpmQl4qdGI2MXJKf6fkKQW2EK9VW9LEW4aFNatDj8ervF1RnHBl2M
P6bf0TA5Kov/0J0xzZhco9aD/QJaHesl3XMGQhNK+bRDk/eo+fG8KM3fTGkmuvcb
hQ2uYBYst+cxG2fH9YDbo4pi7qC7Nb18VehQRPB5+7rLjCJVep1ZhKbqvbLAsfQW
RqLbeGEyKaMwiv8zmkdkkI6nvnwmfMe1qb06o6DM01PohIr9Xta3gJ7u2HQV2lOK
1soklM+NYwD4TMujnm/aO80eKszItCZOhy9blQn/NM7scuGmSvoDCasbuB9Zkxn5
+vWIq3/7x6q5bdxPSZaJcOIBXXGnvatxuIi376cQkKDYksNCV9Y7a3lIBAWW7Ew/
13LtyiU2ewcWNHDk2ODAGyvJ2FDTclRvt34xdtQEiae3Hb4aiQRde72cp2kcegQy
OK+TKQznXJ/POqV6Bt9PIXWXIQvngjrArzgYSGf+ICdm1NAXo04pXJcK8xBCUEpH
p2xxS6cDaFDzBw6g5DBRoRoIURPlAJQ1rZ/aLlM7tqb7MTAgkEQGEPfBIBitN4kA
zk2sRQnOrL6oNLq8RX0iWQML+CjtrbT+WOYhJwg8ENXIPudJN9Zf2l1yzXvl7YiP
dRoHpJCygh/x01KXII4Ox91D6tIlNu9In2dpIuqc+WTTLRIpR1VOlcRxYX2GyikG
NztcjQuFnzo92RN7UGxrd7LQqYIfi7FoFcjIayIe7mcobVopRLvyGEUq6Gd4caTd
D4b+z4foVpnkAycUd/PMYDp86yYwnsilbsYnJ+bSbQ9GnUdYl0aC9YSh61z1esm1
iXg6rXUmtBOdJu6Ol5c4SxnjIkU4RTIKl2KhWFe3+r7Vib1KXCTNwSJg9F/Gz6/o
5E1ToyiV3UfP1hlZHyg98BaIdh+nSoRalKzCrVpGWXHGNTx6wjah6O9FYguzuIdy
r74KVnn0AMCLGFg4b9b9Tyz7ODC39GymcnB/chGysPHQm5ZDSatzgYEDgSD22GZT
mabW9pgPF5yCGZKp8rTSZ6anMwhuAnYediogI1Ga03mJmM74fEtYaY5v4HrZHUVx
cdhYV9wzwLxDfv5GkIM9FO6+OXrUVdM3JShPbPxK8T3dtsffeSDJqaJU/106hZji
yU6xbdLYtyj5Q9E9LpAj14bEP3j+mX8w1+v4io72gQAdybLng/zt8pwmDjwtXrlU
fJtTT1muC651jMChMW8yI/F0i+TW61V/wUgk71zB6wb65usAPwlPqbmUufyq0fUr
kI/lsSawj1JACUixkMMhr4VayGJEbSwRUXI/OmXcte2oWlHpBQjm5RCZ21UfpsG+
ywYXrnimv2sy5Qy6dLQD3oPFwpoXiLoUQWVj5UHEQAj+cVx7blEZNUw2JBKQQR14
2BxBdINM6ADwH/HfxgsDHimWvXrtbuetJzw0tlhAZzFziepdKrPyxykFFymEd8ps
uc9/ZMNgOub6MDQbTpkfbRtadp4VYKFHvq7zWfpuMy5bUIPivYrocUb/ELguxv+c
WPKORfQx6RXdsu5T8HYIkVngl+TlSB4pMECnTtl0/f7phqCRocOdMLESRS0dEyBo
OwcNUOc4brV80YAnuX5FDCZD7c065gk+6Ww+oIciN38E4N8WLk/tirKqNr8dKgzF
If28p+dC/jsz0/p7lq57tf597oLmMtTBnl4fhPOLQFV+2Pp9d4RWE2hFcyql5Fga
MBtpBfj3PmUP/n6hLddva25FXH8DtXKRvGgORRETo5AzZpRDAb3rnDNOUbaYogup
b1pGfPtU1WpTg34vzza3+tok0irM7MiYkYJ5URzhPYmJc2JjvmRm29vWLBzIryV2
X8B4lETmrP6DIMJM5KV0bUdI8Sk2hOBaaMzAoCgnx8coKbEX2YhOFbhDeiMNPRmh
iy2xEGoUWPs/IfC2cJ7bM5VFYV2dlKh6RH84gxsVKrkVc3Z80O2E9pqbwhF2oOlE
Nmi5NcHSpFoI+XPXLtjOrDH7l31tVS0zpKorQt8+UJlcWf6sZ8EV+WLh+58JS6/V
8ghsM1AOOmtt4F6K2p/1bLr3Nq5m4o7w8BiwWtRc9UQPxAvNH61q8AC30W5w7QHK
No9QuxwWKm/kiYoiAM3QK0q3Q5UpgzA2jSMRFkP2fJvd2npPe7HHkNdiyCRYka8l
mscUfcMMsHxrCV8KO6crTJHwy4DMvWk1xI37SyrZMlo=
`protect END_PROTECTED
