`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zINXx783x7RLGvFV92NuPsfqIWOfdspk5vN2Sf45xqEJJUwA7A0YOH2JqJInhdfE
uIkSaHlukco/dKDrCNyknAGWjRsWPGsZBAcyi3uP1bvDE5Fss0VbY+S8jxjosZXP
gya7O19/4U+N3pp6DnUcxozYfDC+zyJDhIJBAvZyE3bz6yk/m5ob/Rw+qXatIkTI
yLwgwjVo3K7Pjl4RMOteBsjVh17CTf/cQo4vK59eDYtM5Ofi3E5zij3dHWer6zpC
C68ApMQ6McEEiMb8RZ1/qWs6Tiv4G8U1nG0IRSHgXa6JsWAkimrufgnD26/eUJD0
vgkHTqzz41wsM+1UVKf5VA==
`protect END_PROTECTED
