`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uNTedt7eJpYAEXNA/ZtJIStlcdhoXAI1w62frSpm21FA6EUNvsopBbhc7yy6bTaM
+Et+sj5VhEhhz9eoeqFewFFZoXHgh2Y/VmkKR/2wP/jz1ybIXyk90WAyFI/OXtGL
6020Fb9uSuVzr9rh1xvsBeF9YGM928dp+pIROXOUc9JgUGB1ZkMzww9Qxm69cHZc
ypZjRDyqnJn9FhkV5whZsqnDem79bxNstDfDYPvWVleKCi/X3cOj/URSwLrJT8is
3DmRKj8I2/dazWNq2wfaIDbABVGHY1GJ78FjuyUGurqWdALAphbthTV+FflwHV+G
SbMx2h3CKUcFHBI/bOvSi8wLo9HfVHl5J74k3CMnWToRjvDMcejpi5Lc1Hpv6xFx
ZKit8jOK9Bv7sbLh0UNSCCRRmlSRD3T5nOvsI4HXnbhtCt02nDELQgJDSov4y1q2
LP7JYRtdoDPwytYE8uV3hQ==
`protect END_PROTECTED
