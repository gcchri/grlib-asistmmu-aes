`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uMed5rKB6oZ0g44BjzfMkw/kyNWE7yBI5mvJITfGvrCYyxQwSLxT/cfgkqCYzXij
WH2asmK9Jnt+kD8THBOrEF9c8b0D+p9aFUg2pNzHWrb7WusXHE35sC4BRLSUjhdA
FpYU2aw+MHnqqJrthnm+LmnG9nN7IMPzI2VGG70j2ACQRCFPTT7eExTH6BxwRjCB
w/OEWZaAg2Elivjyq+qyQ+BdKNzeXHjfq0xaxyb/0j3su3LbksGprTY0LoO40SIn
9+64hfhoTygtzr9m51ONCsp3oiUvuPGLHxUDG8d6INXjJs8VwZqw6yzmmLHUaq27
dE/TIY5aqKhhKU32YopJ8zN1SnQ6ItctkdrJDfMnX4bp5Mk5MLwevK2UXIWkZEna
Ei60hcrTz2X6nUExyfrVhBEl2RQReYbW2XW4ZDt33X4gx1cOpV3myH0wKn/AdWha
DtmMOJ5wuuWJA9dfRRqb6wYSBRQD5bNR4cKiz9gcxKnYupvdYuGT1v8XUCZKwcWD
49scXnS0+hHYyeFIDBwDHeWzdUVZK1KG0BORJoe0wfkHFmrW3sSg8bGWZsmdFmTQ
bYv2N3CoBI5b+qhG0gIfm+q6cb8+ih+YP65AFft9nLB//Ach3XnPGpq2DarMRaiD
bFks5xLt2ZktA0f58G0vTR3KF5x+cHXUEgY8QMpH9mD16IIuE8Y5MUhprR9zmMHu
+5te61ZVho2zrOlPI89HBtBiUFY7smlvk7wsUHQgXy4eY57vQ0YptcqE/6jWxxHR
5w9ZslDsLs86xHi5LF8iY0ThyoBkPyl/nm/3y73sBDNtdeAqQwnLJ80W2PtzOqVM
CHa/2bX110nzLkpXk7m24b3v1QnRTJ5oZRniQKViymZP/TeSZYF2buVG2XuC9zS8
9ZEOdW8ZIztu8Jouz2PJNh2psJHC16tbJKnCJshvrZ7hlz9suHIMkfWYY2owNw6u
7R3doM9qEAkW8K10VjGYmiyxX+mti1GpsJn4BlSCMeaPIAwe6E2n9+Yz7vu9qwKu
dSD1FbQXmoI0ymPBIlwPJDZN22cJI9elCmNwm6cFbPY2/9+QAxu8sp/g4H+E9Qcd
yioz5KV/cB4WcPNi5mccWexCOOy5PA9GRg4lyiyhPaat61kNutN8rfR/wjuZyVrt
1T05o41c2j7BGIvJvZ6HaPmWNk7BddP1Df6C+w6AFkqR+vui0pImYLE5CRqJ9/yi
ETICX5sLL8nWUOhz4HDhpWhZbm7lzF6OcTaUUn4lLM2cD87KYR1ORDK8pBM3BHHT
zDpqUFXtuUDCBKCS9w/djdc6/7tYYtOC/LzsfPGl4PGQgpZCKVRmrOtLo1VDO7So
PDwZLHD5SbsorTG89LL0GjbcofKCW8ueJ1G/+BkuPLupw1BKty/jMpYveCQryvXM
y/OA6eE9wY8RQXPdg0Xa8Rsb14f8381Fj2SY7LfwdUGLay6meTJeCGC5kj7ArhBm
dhtGSVtTj++a4DTOmbPoTlHTbXsbGUha3h9/D8qeE5r2p4P9hs56vmpC6VAfHaRl
Wt6KzEuEFq7rJ3UbDQan6y40ka/buQ08sbAgfHHU4ptw+naUB4V0c7famXRM+I7B
DQY2ICz4JDrq9QgOzgjtuFuAezCIDyKRV84v2wqv8Q1BpBmZyYIUC6SqgVjAu4Ma
`protect END_PROTECTED
