`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uBil2zqhSDk+rdnRFc9VVSf8wyV+2PtUwN1c5TPoiIrRzQzTHMuycXhr9MeeCfT7
ziT6R6Ywo/XXITVCm2gscnjiiRznLKTn12Mg/kS48P+CnPivMZrGcFtTESgrxvcp
kYBGedQbUs3a3NGIS2HSgiuhSFcciERAiTsL/9B1/fb0bLnmHC4h+NFJ9e5NOAe7
4jR/DSD/UM79IA+VzGDqkz8fNy/mA3gmzoGYk1LuekrIGaig5i85/KTPnSWFVgSg
Ldqc98nF7NIM/THJHNm76jGQUzb53WZT9SHQ007U+8pmwj1IiEOp9c5KPb+6ttmo
xo5LD5zcIU5jx/TKW/aGnTlkTV6RXfrpiKZtDNjwrJJIGed7YkMLvmnBY8NtgiDQ
srzvM29+Slak/nEEySfRHufE7q1w+V+VMvODwVfGBkg=
`protect END_PROTECTED
