`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cCTMDABXbRFtwaE/nbjg+PqzOyHcqsa5gzfghn78fS+w8lScyuaJzdk5cnKTsNFT
iOlyXGhzUHNzi0hfWoa1gEdGZyMW0ZpV738gNezQIjhlk8msAzcWkWOhzOQNZWid
f3WEyaRnOJVKGV9AV+jpJvQOjsJTZ9swWWs28ht+tNjHp4S0nIfehwluUr0e7nJU
RbunohPFr+OsalAjXt2U1gPZX/D2Jj9nvyn1bcLRILyErDaQHBTeYJ9rClrzLVhz
Dhvq7v3LwSLpogBYuU8c3h3HhfWKg26oeT/EZpcuwlNDpInKuqzKc3qL+PO7gify
Z553NuZmU1fMeJzaSOxQXrFb2eRPi3NqPOERuSpFc7msLO08fe42/Uq9IuJcJNxz
k52KQ+Gd0+EJN/UX2dGLOhD7ycHSR7ilEDGX6iANYx9hs9bKs5VyA1SB4RFnFMIf
aLT1ln8A2ow0uZM2m9FUZ5sXGdhrzgtlcOK3Qwyqz8bvJE+ZuqA71GdLLu/Y+Wcl
qWJzdfUCQikjzWvQFUla3m8hpIdjyOHWwuFo6ONzd3X2ahuK1bILjhR47EWP443F
D/yN+hnAu4y5KuraxpjfK0P084zpqMe8drf9QYpX2bgnrQrjHq67SXwbSc5R6zEb
y9rHuIx6+2OJpMoiDpcpsFF9Ndzb4M/XUtEwhQh9ad+M0wtSoxtP5KtIo1jL2daD
f601vO9jTCJRlmxdffs3iceBMsfIpY7tXB0e/x6x506+IQ/0UQbKVPFkTqiYB5Nu
WyRtBGru2oCrMT+5pFPccXpPdC59QGLS1bAQWblHe7Izsl6wfp7sjb/XCfyGNyON
POC7QULcqP1ARju1es02fWCnk9tzeNYZuTUX30TdN3pz9t85tTrhY2v/Gdxf5/pv
KMNXRBUMZKVp9+rYeIl+1OXf/Th2CdYo3AjbE9Bef8Bfr5GNhY4f7+TdmKVi+bYK
jaQkGJoz8ZrgDPQryvLt4rqBpctStm0wBu7B9B+uwEIoSj70RMwg2FKlPoCanyFS
BF0lenJygfexRLRWJvYc1Qs07THiFpjIM3axzZtgutG2mjk7mHwFxsVxfQCMfj0z
spI2gkjOWEmwrL+KHMQwtX/eGDMrpuykUUZooPw0bTSgtFq69gZ1yMKu3qMW92BX
8QnYOl/tZxtclDxdkcDyziCkcNAsaf4EBmsaRox3Tsa60v6uL62PsQRHdzXVl6rL
Er+3JxBHBindhwz6Gd8ST5pp0rasWayk3XQxHWIBb0e423Z49g4Zic+RjiwJFb4Q
DngX8ivJ8BaItc8CJYNh/xkI7PGc7pTdOd0SG8PKNM0ASzlAlAoTCFzgxWTZjb4q
jPjaYxZrqynYe4GVp7yqQlcIUlHQqWxpns+mGPBF8uqmzq5Fa9c7dOU4jqm7oKds
0iy/nQwj/ely/HiAca1o/eXWL6L2PedR4bOB0xIkGeYinLde5tu8S9RhrINpanlz
tGBq+TzX1T/eQPIbEyBrlcnXlNydS2WBs8fQ5w3UjcETzPhF5fTwnLjSZWngUwIj
tDBHMUbyqODhgmMDELJgN7acgLhXoajMusadx0nDBaOZ7jWprCP80ryoTEE/8svZ
4lLOka4bBA8vz4am/7Uds2uqMajUaXJBmHGV5H42okYyMZ/kVyeY3hTqlcXDq5E+
B7278oGps/O5RD6UAZHNW0XhmaHdadL4HJmxAemOR3jxZXOHRmbYzVoBScmMa89t
iZRjD2pxBI6K4d66GXVDKZxRxxa2UUFHuDZzQYDXg6GUrJAbbsmHaRhz7vq7N32+
MdediAfw2VK8TzWsUoBB19lfrR6siXEq68rP3gU8II9fr7PeOC3mgJoeqK921mPT
9w6Y39Xs7iTyxvLTNZaT4HvS9N96Tl7FNVT0peh86fNtI8waz7ghShT3witcm7R4
uBBwYYQnuuqVfk+RtmJomnlOFYTmL4fWv9BGcPsRFD6+XEamyK2UdOi8vGqCrx+a
XmYIMj49QDK9lUk532MFFVGSay/sooASdvUd2Y+Mrsz0XpPKcqrVY2s9lHpj5Ist
5peGt07aCLuLAX0Lcvb4I6qYOgu/1/788404vosWXrISYbzuqGJTWJ6YUq71pDI6
nLYmzLMJNdsrQWrDOU9eVv2oWsMrBqKbgjMozuqNndLavowsNs4AoV435f+bHdzH
VRxEOFmLaKWn9Po8SCa0ky0H1X4/J+aRBw+q9EaPp3yX9EEs5umvlr2/Vc035NBE
U3sQ0HMMTudPUe5EQkN9+Zuxa+RrMce8wq7dis1NLQa2rOzm9NaqT1G4x5vX7Vue
hlF2YtQhvXMTiAuFZVg0l1d2+vte/53Q9HfedZAA42ujbviUsbo6TAfoOljqYIgq
yMVXKfTKcHpGzAFjay6jbNjTtre6VGa0/HRzTPwrwFAXtWQDV67f1P6n/NEwuroU
/qJl6RzDVf2D/C8cvl7zEtwm3xFhPobFyH8zt5F3+lncOFg3hqpMVJpfMRExCvSI
ONUKVpk58/amgqMarmrRGOjPl3q6tH8JLsPmr8yMvVXHZ5EthdBAxVPE8j9y5xhK
k/v6wZkQBYNNNcDr5MeE0hG1kTNnCLgyRCfeckO3JuoakeHH5000iWSb5kk2vA2R
XywEQjz78RCGhrT1DiZyvNg1yRqQddPH3Qzb978kSG/fKsFy5qRFQlMH4BxUYslY
ApjG6No9T4sPL8EGBdUPRg==
`protect END_PROTECTED
