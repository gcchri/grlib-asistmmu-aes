`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nydy0v7MxR6HQt9czwEOLoyRbmvFWabI9QWM3p/l2M3mSJKVlU/DoQttCuu/eqE6
88vn3wFbR8OpGk0d1hdQtBcLlbc6HmT9ghYDd0bLbebpJ5YgnnyvCsTJwI6DNWJJ
/eTQIbuGR/8A+AlfNejWrYxTwTE+5R1iw2eDJzcr5U5PXmlfWpxFbKFerTGHRJ5a
cUIV8Ltdsy4RxrrwLjhCmTU4iSKzrou8tYr7A5vfK44zIGp4rvZHPfj4lWH2tnrI
Z6vnnEykchgD9LRpf0J0ZaNanLcJi2WUHhSPanVQrgyTKLQzheNpAaSyHtlpo1/m
kYNs2Laww/4Y2Or4Zhkkag==
`protect END_PROTECTED
