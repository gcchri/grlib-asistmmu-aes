`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HsbIvNGyAE1YcGVdWZsDcD8uIZF5RCrWAkLyrP/C6qTAXunfpkQ0OfuzbuTtqJI8
cNEqNhPWMRQn7VhoGNXzimIQYC+sHLsrIfc4g/DRyoWg72H7AV+WhmvP9imQwGt6
Sz/pJvmaXIs3LR1wD/ldQ8OKhIlf4kCnQzZi5GeHJp/tfqhLdF7mEhHO3h7EiWA8
RMEHvxsyjh8VRcjk254sBmm+0ck7+SzjuimoXG9L2Wbp+zIFielhsF8kNKkYcg9k
jDAdvANa8R0fYAEXIQFYNLCXbt39WNzKI/OpiWI2gKHZFH1uS6R8hAkhVGI4U2er
VZtSKzTixL+ghmzmEiZcscJkMvYDATkkKxVqD/Ki22k48BZR2RJqexAD72z/or2n
nIqwY7slc5v1iu3oVOJ4Tw==
`protect END_PROTECTED
