`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HxV7AOK091xwp9xmlMS5gGy4wgvVzJMSeRVjN+e4rz48d+jb9IOjziUqebTNFoWS
8JF95RBrdJxgYGrlvEBz9sE3kYbcHRI452U8IMPJs1XSNBqvWkvVQytOtTqkFc76
l5CHWe9VNM3wBDi4hW43UydI3/GWXXhDsmXMQ0EvRE9jXhHAETKYd88D8gLthXHg
gm9r7Ug2S6P+qaaJcX4/clCIrfFrjGKLBLlH2c98usrFVMDcVT1lvWk5jBkUWR8K
XGl5RNtDp1Booz3iMP9t/HstZ+9+8Oi10t61NPfI4LXGoWNYcePXT0Ds0HYPqmnh
4GCGQ1vJPwNE+T8U+tNuoA==
`protect END_PROTECTED
