`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VzJEOL/+iO3YnpCjiR8fx27M40eUcO5447lwGonlWIWzPOOp01xVar2vmIsmuY1O
NyT5T2J/SCz3kdGCseXYiE6X5wd6yWpcofppxgF1LiXC2t8u4bB1x5CERH3VJQl5
9OrXWvrkCTLXVyP5BnyDrDPsdH6E3U4io1wke9G5NbSRGgpXdM3/eZ8Xiese4vGP
RkEwel68WPts4r14c7jtghBC8/qR0wl8k3AJN6aSZSzItsCmJLOH0DuAqaWm0o3l
Robm/Ul7dEz6h7vVO2hRXAAwX2xrAkxve9QXjz3hyyZh4cu5J9c6LP0yoMkMYItY
pEtO5fipICK0IxfEikSsAbZwUMpV91my4UKea6w1UpFWsVgHtqKv94/EER4OaGAY
U7T4rtDJ7ku7dyaACiHWlA==
`protect END_PROTECTED
