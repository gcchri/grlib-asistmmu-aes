`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xJvDVc8qULbY25A5yf0iVaf8O10dy5zNyt19PLH6qJN5hruUMzEWQjUx/JVE5lkC
TASkwoWJIC1RXWH0tuJQ10mPnsAuDPtQJ864YVwX/RQClcQ/m4GOTaRcG0fpBs4U
W7rltOA3ZeqOnCY4ZsAOnvy9jHo6N0xKHZLuRc0W56m9mDvXQzrNaGzxFfzH7yup
XiWWe2R8ORDd3nRY7U6pkqYMxUTFrFKVryeQxIrnzewwDXtbE+N99j9I2izDze8b
GUgMONivL5tmHHle7hp0Ua2gUPyj5wURqd8uw+QU/WkPlE7KM32b9YtaTiIbCNR9
f56ZGJoHytMWAh6XoyN8LDhh6iw+YsCdoqbbhRi9aM+/TsTBI5Nf+8Lxi8fi8lmD
FtVsxAegKqh45DsWyaG7FQ==
`protect END_PROTECTED
