`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9fakkoJqqu6QsufkLOB+T9eQxvtKn7AlTfYl2l43ILtWQrIbCJFA0i9yZwa/EB3+
/MvogGpBZv6ZD3AxmZL0+S03HyllF74GufXMx2nms7JfkhXwl18sWXKgkwHk5w8j
p4XHHgaAG0PrRwPjnhiWrzNCgOEp4e0pKsWkBa8rP9GeWQEYu16msaP/KIBbmVAn
pX1heR3ed6IH30wXyFuQz2fgJIcs6L/9SDR/DuH3+an606HfjUOL031+Q8UveVoC
X9ZySUdNnJHQOITxDCxF3Vw9iwPEbi1Ia43xoSdeXMv6xU588JjaL3JYL5IRYBzD
BD2FekGEwifXLG1Hbeea8AfWd4JlQPe4mPS8E4yfcUo0kfEcZUlWT1hsBATNdHC8
IysR9KbBi+lYcck69qcw5LTEMMPZDVWx7Fw791YWDwX90Tz8AFpAoT5YmMWYmHlE
98ONVED4nD4ZG8UVJvabshsG/259BYbWbMNUDDbBBKAs1bCSBNWEYxEtfGIZjngG
8nxVCUshIp15YAq0neHWciQb+GHK1h7sh6lVa7QfMqOHHVoUOgUot6bZuSlHh5P5
GfoWn6FFLUUY31Coltgsol3GNKAulBzr6UKq+B1+zhqErgPb08rDKAH8a+KWAoCl
GDXJCOmafnwskuRsOcryKw==
`protect END_PROTECTED
