`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oIWAphQkSR60eSI+xcRZ3ce1j0E7hOglRoN0SszNic8RCRJ2qcNI4vSfWNyUwf9F
DmBwmSRXMcdfJive9/SP40rdahB9FgXK/j1DOubyeG+oQOuzTrI73WmQB4F7Pwwq
BV5hZ7SnKY8wYrlaDGKmuxS1k/oS8l9glQHXFhx6G2yRv0yJ1eY2DxLGprszBwKI
jDZcKZlTl0gwOUCJfmluk9z/cdtD5Uxh8rdYBRlaSsByzyqXS8kV4ePIKP4OMdjr
IYaFrxN5mZefN5qlBKGdnvYNxdubRVS+p9c02EMuptrtWkAiDmDe4Zku8jdB2hfv
B/pbFdLUaaRC1dcy2+X5CoyoQc6xbrr30CxSAaiHt1uh7NY15w2b4f4dPckcj9kc
CLY48+kH7ZX0zMMQi/bwmMQwPojGtxCRpo7DGsVXdxhUGchb9KdkHoPFiioN5XST
E5+qFGdRoB4NHy+iAsWVt7zqQ8BAKCZN26o51oHBEdqjcO8u+lBTv5GNkbwYnYUf
BsgppacyAMfi8+7zbbpAGm/w5IPR+iU7f56QeHOmKHiC4cNjfyAFQount/bVx2nM
BzS1EewVy6QYjtWCjJ1Z9Pq7CcVfpympzDgn0T7fmipx6sebfLxgS3k6GS5y74wd
beIc/+dlzxV5y/BXKi6K9ytsYNXSrbnJId1q4oZSCmnBV/p4GDVyZQ7AkFXbCeXz
yYGg6nifNI9SdXk3UL5WnDaU5mV92sraOQsEMapeTo6nCDkaNIOo0KObZI/4bc91
/dlBxqrfgLS+uz9dym4V0osL2Ou/ATrol9yDAr2yP3BybY+ZKwi9bw2WcJ/1k2ew
yjBmpi2QHkjrcQdkCTUiJPLTnYJc8gEaBa0itiOZfBsNqRwIe6LQSiy5HQocIXE4
Wpdm06h/RDX1DSFQyfNdSmOE28uMw5S8dWMhqcwmm56QV4IUeiEKS5rRa44T9b3Y
L3+XpDGROFHXkl/x2pT/EJF3zLioV+kaFnNSzFd1qfMhP6ostw27lb9K709rUbTO
xWI6FSKGSy8EOFb8qyaTM3t2X22/jqSa9Kw30N9BDKLf9DUtstwQmNQ9/hXUzFGF
HwIiQf26EOV/uMqvNCialMWhicVlb0ovlCRtdQRVRtmDzUS8dnvF02sRsuavai6Z
xfpUGvyb5XYH+oNeOWIGcSJ9cPh+7ocz+iOTTGqBf1QiSeBJ47PRr3SduqsUcXIa
IhYLwPARJYl4E6/4K17m4UAilQJWgLPOWu2Kee+m68imyKQtYJAMw8dm3+SWQR/R
QHz912usFgTpT5K/aINjEmx1VHyiXYpq2gYIn/A/5xlpWkOufN1flIo3fy3PZlmG
lJgQDTLxejjHpirgbcgEJkM5avF+WVbU4YLqIkxbMpzMIrkpVup4haR4AwVGHPA6
0Z1O+uVyD8TkTLfm9Qjg6lDhb2Zgrk9YJ67aOE0BSpt1fTIB5iz08AU9FmAu1mw/
WZO2oQlIIYHbhqGKujnJbyuHu0cNfF9H4/IjoGla416DgQgRFQajR4SY20YN/QOq
Ev3nSNVCsctLNqBMwzwVfmVqalwsx1cEAxo/UC1mUmSgK9VN2NuI0LonHDuTNPl4
VCKPH2P0s2qJcMoMGfByNu3SSVldwBhnCLW9RAKHjt7Pvr9iWRecdI/lruQNSFVj
+HeX0hiF6IE5iPM5UMGqzQmjYERUgpZb3YzKNsUtjNPxeL2I03JKl31nJVZxT9zt
WYIp0eYZGQMp2w+nha5ppguS7AI53+P6efQrVnoMMhRhJq+DqehiNNlY7MsEqcl6
GWwXnOZKjfmmUABK8eZm5VNWVzZCGYvDxECvMqvm+Kuln1GntcyNoUGzyaa+OTiX
WOC8dE7CGP33RMjvgFGTHluIUT9Xk3LI5CBsI/BpU0PikOj0QNRz7wRs45Lri25/
SEgNpe7sxv1YIqpq8zvWnwGOdrRSNz6DXqGkFOaCWYJNtx05JAW4Y9ge/JXfIqj6
ynvMnj1elAJ6aLVmM9UNT7Zm8065Zv131ud9q1wBdwxc44tgPNgewqKuCS1ctwjL
fk+xbIraB3QWAMCEeh8XeKBtaEJvFAw5DAZbWJ71ZLUf2gF/WEW+MYzr2Wm+tEia
Fj/Pn5UvYjwF6CNUmdPZABE/C9XIsHgral/sj7Or3dDt5Jor7uQNWVTDig4MgOGS
FCxKivy/X/6I2Dq/cXV8Cg==
`protect END_PROTECTED
