`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QTUITtjHw99uyeBENBEoZAEXzzm+Mb+nhEM0NbYJgNPIxIt9CDcMQcG47//lyu8t
LFRNZ990dLaTi7fX6xRkMy4/buI3FsQ7UrcOlh6CP9cisvQTRfNxBiRY49BFGIUJ
YAlW7yXOsRSRKRedwesvkN0na129iFOjSEKiYjPClHIuwCiKUADSWI+004o6keS7
/Posn7BHsQ3sXpd+bFXYctjhGeCYfhEXlo0zX76r7LWe12ZS5TbCrquUf0y6nCoP
kj8CI0QOsdRfdwoiJIXqu7Xhm1/iZxkHuhHPOR3qTlw3gXnry6niSwwDEewl8QIf
AuJtvJ0gvOuqQLawHt7MLRL+WooMexILYNdJ7e29ZEzOzJ2FGsB9DgqpHxObAH7+
8aZA5Ak+tJk0FzE/g4U210cJRL4Tpsp1teePLZD8er+5yoV+9fUZQfngVG6z0OSO
8d/uxUWAJ8UJ8CyGKCO8g4ppVuzhvq+Nv5AkuxrWRLkbEfPPPrhZ6nM7gxaEjkID
pd0Dguij3B7Vz0W2O6wNSzu8QRSGVJX9TQOXowv6nOS6e7b7LOSzSysBL6zTjGQG
uFOmbM9UumDYVi4RYirf13gXXk/0H1xxbF8Jq8GYFB1W+DeyHzsklDZYs2C+dwQB
6DA9Y2dGtCPYULJXfe14gvaq+RE5cFfXviImddfFKPKqtIjf9ggTD4gGA+Snl0cE
tcZWWYzjm8KLIKjXRgSaNVWROMif76FwLLFIpRIF+F1hP/ae5yu8L5g+5YjSfJti
0/k3nBqSpNvRpRGbvbl/dwmRgbGyXT/vrb/XDPWplyyRYOjZgUonChXfQhjnU3Hx
w+TOmf0CyYcMYYsmLgfFFnaZuZzr7v0lMtQMq1yrAGeY4m59m4Cjo2EZwOCxEtLN
jCyLmVi74Nu9jL2RCOYV518M2zVV9SfJHAx8rh55PzoVVNhSbao25qydLMI5gxzb
pol4kcjkIEuF6F26IsakasvKm0fcO4YDJETSosAvdl62uDoumUKrm849rUqE6oCb
vK8LZazS0DgKJkhiZEopTwIKr4PCPcFwwMXS/H14lW786K+PaLZfBIrq9eWGNB6l
lZpzBPIitrVRGaaHJNi9Bz53mPBVzPo299M8WVU9TcFZSiuekqZ6BABj16xEBAP9
fu5woy+u3NbEOc3E3SF3y/BkyIfTxtXbJyDTrofM+CjXrPEukJPFBVbHQzBV7rfy
s8M8B70v67zj6cAvL0AC0WViD0hOllJrBEuqVVOgM1b2lkULiDjSxSbmDntU7vdc
0KP6c4JaUI+ADUEBhntkjxYA38uz89SpT0KuZKDgpzud6yioDEquXhdUnZZpBjbn
Ktlokxp7R8GrE9Se99S0dXbHt3IX9EtH2j3xF/1nMzuZNRwZaJDIX7QENPTJVPTP
5tKrxxkZFz7F55l6IuZkhgUkYlmvKftopU4YR/Bscsw3wGR3WutukkkV2YXE4qju
DN0vG2TrvQI+vQW8H1sjQcB0l5lc/uLVlwWfgsDdTw73qltNOlk6WWMoIfX0N7eA
71DwZfu6TL401SPeCKZECNwpzQ/tXiBk4jayX73lwxP3+ZjiO0nUjQ3WS4kWcNjZ
E1RP4htUdwnfRTnppIEOuNa29hPVqXoLeN6x3AnJCfDd2CR6pzmwBClWUxYuPyUI
2x4UjJJq4KchGzlp0HdRoIhMCspdIjago1pZDePrc4J6edcDF3IDMvJ/7vTSbpB2
QB5cn6M2sedEVEYeYpKClXF6M2oCoVzIyduYVGmZrfZFz2V/76HbB0bp9qFpB1hS
fmGBOKKs7LPe+GEeN0AMaHmGqmHt1yoTzey4BHPNKNwpHSm7oVYmDxQsp4iwcM/t
+QcfiZ8JGhObruRwNktyukTgPHo/LPTPqCzKGLgNi2Z8AjTAhlZIdfWjSyjc/X8D
3gaaYG3F5ZYoPMT0fdVdn/AyYEfhvzZ8T6QTmcG5UmcGCpiVQnOEGqqR5eH7MIIY
Y0+o8JNyCVhzs12vJOoluA0Wo2c6r2vqucqNVKYN9F3lX+IHWj3HJGs7ahQtPUJ5
9BlG5u49Qxu1im1ckNdwVBl0lKjdaPZEItIizPc25qvVtBC+JdI/vk6c+G2Pd+U7
92OI2W4Q4x1irutlCyURh+G37W9hNhOHIRTf1QKL2QtcBe7dWzRVxxiLm5/RCsTk
E/LZOWu7o0/5hvhmILpox2rDDO9o4zTd56vQGflvDpl1p0J5Ph6EKxIHWq3dFM5C
zx4wYmo/sNQISfnfy4T707VkrreKrPm62zuptyIFQH72t78kFbld644Fdrt4hZaB
3O+1vNAGtuODCpXVJ8mF5klBcT9BHVHFPIxX0E134QM/YbY3rJU7p+UqQk8ZMI6U
AHK0TjRf3vp/jeGuk7iO9Er3py6XE8yZzMtvb2Ja5OAo9JQ/en9+D0FLIBHF+mZP
xeOrsYH1iCc7GVBo6QatfHLQyvfwRxhExq7VbIzP7FTM8LgAfL/Gac76J1RMX5gA
m/mRvYZweymzQLFv+Gbu2GS1Zzz8LegtTzXf/vu9z1bM32J5WOogPkUuWbkVJcfv
EB/CPITlvUId+lRwyYSvNb6JrvnDmMU2Cxd7RfRfDMOjIwlSTLUoEib3RRSVnd2a
whmtVnPPIsakBknpoUujQt56W29yr2KJt1u2WK8GspdGsquq7zgiu1vlk+qZGzLq
5+PvPqbQpBkZSBFcdF9qrFQnS9P8OQDMSxzx2mfMyXh8N20YuLpnvr6gSOf1xHlY
cT9/PbnQKKJPYXxoFP37AiuRJBih3sRHBmLuqNOW6lztXswsLXVVDordMVMP7wZD
C5VUHvgFO4M+FlIQAIKFm5+iRnzmltAeyzbeS2tFM9vqgO+IxAGt1uHDNIU0sHMT
hafhIG+jC6sZ1t7bvHSv2XqONxT1TZPk0n+w+CCwdbzqVOGvpSo4anIUHMpON78r
uK0iNTAoZUpzCAnwbryeK4h7GHjrRraiaD4vRPPFB6V88waf00R8xzVLtK5Z9lCx
SWx13Y4qVK4SD5o/3lVhAH3R83vT1DJ2qvnJoCwitloeM5iRhcfp9jAMRKfCHIpc
`protect END_PROTECTED
