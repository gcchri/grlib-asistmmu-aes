`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oBoX84D78f2maUnNIGyvT4To0guI8acHwt7IrOr9T5M3rTUtwyGKiLWmGvLBU0Ge
JxyrbPC2yRoa96LJXMEkiv7ouYlx7IOjpe/FkrmZ6JcBKYuI20+rvafm87a7H4Ma
qW1VSM92XSEBCpgFzkoUnT4ytEQeSKyBPN/gtjJAc3aEXcAHZIK6JzGhjiOv3pFI
xukzXVdqqtbH8xD5odDZO6TTP8IPoaCrYwOdpxG0J4Ml5pMzwByfvtVG2C53T3a6
w4cAsWmLRjExkopx2TXUUt4yx4h/hc5BQLwRyxLf9tuxDR1ARJxgZsYItH0XICn1
WlijtL8oPo20cgIf/zeKYEabHM62EvG3jh3IwPCJmmkwaXZZx5wmrvSylqNmngYQ
uPBqmluj7v9xGp2H9O1sKRq1DRIN3x/KRoSXFvphLQsQANQ9gcE9D8b6l3ZIaY2t
`protect END_PROTECTED
