`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ce+IS2PJDpWGDiihXzKnWwZzV+qh5YpD6N2D6pXF/VBYqKKJ7Y6YK/QuYn9tuZwf
zALUatiKuD4rT8DTVJECcO7DsdjRylJLGH6a8FAAv6lBLDYNUvYkjAzGnzKbH9wq
p1+RMw7+coz3vGdnb6mcd6nI/B4WQHGOkQfnhqWPVsKIw6G7l3lQtJIdPwyQKHvO
+rHEX8Aj9Ems1aDajtg9s10yyNp0wocZbB6O8mHP0WxlT6A8xmyup9bgt3la5hNy
bHcUwb3aTyvd7wiu5nojOddp2dD4OvuiD6u2HjRaLa0+6z0N7aFL0+KW9eilnO5w
S2yP/n8KVJyjSHKDH3+TZxdNRBtJ0uR+IkGfM4Wz3g9LxftDg92drfxO+R0Ny04V
7S/Kr2D2jBmG5LiffgZUx3j9JIVmRvxdcJt9kBTxuUYrbhvvGAzK26OtSN/LoKo5
fejChmkKFRRH1dRlC0hYkFKU8do0G8tdVG9kvAyxO3f7H/rZoRHMl2SJuBr1VTzs
zDsAXUHLOwsl5rDWPb2B2kcbGrIO2u8UL0IHmQ4Zq3wkj3wL0lZLML/+/SLQuMr2
XJ/0i6A5YHg3z2oc1ujPLnXwlhYPWNtwOR1vHyVef2M=
`protect END_PROTECTED
