`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T8fnONJ1abZkceGPeK23HmHU6uKcNdfUpjTzmerbfIYCHk/lXbH4S2SCZllfrYhd
vZHwJzN2ubRVF1LrvLZQaIdOEvAC1voMAID1bcnbHb1GINWjQPc8bf3SW+wHBO5M
D03u0AF32AKPVMrwOPQ5zvlUf5wcrbTZb+KlZX+2twXbo2OacvZ+AlH7YxibBn/8
LAwWpbxFR41YzDeB7y3JsnKR1uFxJA9u7AJVwYyAbTVfaOKb/JI1EEPdzKrTbfmL
olmMrgizU0WJwTyrtVwO0A==
`protect END_PROTECTED
