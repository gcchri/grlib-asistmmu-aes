`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
juPOur8LLIrWV2VAV69dKXFA7G9BLcqZHkYh7VSaaYwnFN/JD8/LTFWE2XX567EZ
UIOxqLagjGPA8il3F/B99C1E/ZEDDF2b/NwusFuF9QflW4xZSZlM8yulp+E9GL4T
5Mk0oqU7ndWErdrO+IqZk1MY1/0u1gvkanG5e21i7SLVPuqNV6k8I4taZqzpyZe0
5+JAv1obPATu7JYJb5p+Z3hIkD3uOz0tH7S+8T/lYX1NtfuWYRu+lk2L/4zcWXQs
PNUqwqf8enHEYT5IJiVTW106XdL1iMRkXfVXF/BKoYsDCyF+GGQCZkafeUGzgVPm
MXBcEJ+iJeV9ixLfSNmBTvp7KN5kTBLPdjvvzWCF84oz1nFcQh57lSMjFruFmRBK
sQQAmGK4iwo0ke2q/6HUVMu3925HX4EC72ap4LyOuNdkt06wQ4z9an+ENYMxZ0T9
`protect END_PROTECTED
