`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zj8dKPX7L3oxf8hlniOud3Qct4zpkLy6XVbrlR8rKO6urNCVERnBtsIDBJf/yYM0
6NFfEGbGQPMvcAmWt4dE3g2+7mioiHpTIjvuRu4+4hoyOtbLBkvFPfLOK3Gm7+ul
qn99VWEcrw3ISa/fjMVePVm1iAiY4Mk4anXBlfUpI2+zj2uP4IE2UR6mxcu0VXi6
XXiVioMBmvIKHCWQCzzIpZfNuzBQzg3n1tTMe4uzG/oc4Y8k9TQ7qbs1nBKryo2a
RApen0s6ud2DNcark/MGCRPAvSHzaB6vJQMWXFdVyH44nOwIaOF0uKxeOn2lK2HF
aS4SjNhevk9z1yPqdp03ZxBF4RdDljayWk1yoQglx/XgQSJoT52PiBy9i76S5NS8
29VSflTR6fyoBl6oftI0ZgmSKTkk1uknUTKLH8t/fIegWN5tvpMUr60dkL7GLGl4
xmyrj1prmsdteA05W5F85jtpjHfYaN9EGLp4gXiILTljSFk0mmggBb3SsPNfyc4H
OP9db/BENeavcAFBdHuVpsDgrPFnW4hvAUay/tgdSXTIBpZIC0GMjY0m0vwVPswW
qzrNNN6ytEOFkAue4C7SxmGfQdDRmk/eEDMQAliIY8L9gtktNrZ/PgVc3YuqmxBE
MNgiuaSyawTYD/uji9/PpgNm+1g9tRE8S5aea/ZIeXCjGOupfIu8sr8Qh18HDq5y
hLNgcofQQbATwa5f3Ye8vsZRjQ3D+KFok2F1lEMzLk6ccS+TcNqJofxgt3x2lIt4
gTCFY8pxm6Rp5HRtc9czF5oD8lNcGybT/wyweOBeNl6dhC9Pd0KjhD45ZEB1BV/z
JGGBduIQ2ZWe33rLyotGuUifSlkzJlo6xU+qVQF6QyFXBTKKPwR2klKAvWyW/f76
kA6tCOKyf+L3GlPPpBDjE8wkttGW9g+NQDyfkk6CJO0lMh2KXX0tEqpUursz00LG
zjeOZ7IhDjrz+HOUskwyYQM2mgaQLEc5SdrREBgTg3RsbngTSrfm7zEV2DNmhe6E
M+cAMlbeVYBpWkM3mRBHy1COyrmG3AyP4Iw29/1CCqwvwdV10zgncIK9XSsm+Fow
CqZW6x8YdkmMGyUNL43+Lz1szFRfu7nDb9z3z6TPC1/EzRyquAIVt0TLs+DzYy9T
VROB/MRsinJTkW+O9+SykRZK9XvkZIvBgFUwDLjn1N89e7BNahTeq8bIUS++PBBR
`protect END_PROTECTED
