`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZBGj+U8yKgeHUNe8YMfrf4K1En4QtDA06RXq2WOHZ7bQIrxJK0Tka9huyFwSm0Jo
6/mg4YfTTtpD50w91n0UFCT+B1ydCV8WNmn1Hx7f02vuiBiX9IQmReReGRj6ZJRv
Q0vd0lN+dB3CX8Wb+hP5S8MHwiQN4Op6WMYq2S0/U9ECWqZj7IxVE972TZbImLM7
S5HxJK4oJaxFLVm0kIBE6qBMvYPXLqp/NvYvjaGDBXJ5Z5Uo6z6i2DC6OUbk1oBe
Z5kbdj+k7w9Eh00Vec+R/OkASGu3RJXQt8JztF5fMs/GU7drrYGbucRNjXNkKb6g
SOMpXKrC51v5sqg3EPMo4linvUFkAtzg/aHipQ41hnwi851Exqtwba5we8YaD0c2
7/k2Lq11ipU5oVZ/p4fxyjOiEn5vOaHhS0TjtGamx3e3/7gXw6I3t7PQMFNMIU93
IBypZtTIDgd4XcdtkmTNRg==
`protect END_PROTECTED
