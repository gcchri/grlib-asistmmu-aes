`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h7QU25u2iqD2LWtMoqaR/aEC/gijIlVzgUuDX2po1OH8k6XMAHeMTyxS4C3495+b
6ac4AqsZ3PxJcjuwZXGbWAOYZ4RNskiPlniufTv78gAQ8ebG0DVNgsSebi9II5ra
KLe1jRLedgv65VCS3TH1ynEwO1j5Sz2fE3zVbdMkJV9psBRUrSUVgCeB9RpLVQ+5
lSugTGKSlKpaBpy3o5YlxKd+MsUYQWJbuaaNBpo/e9Be7cfCv5ZpFUiCpKDIv9SR
gi/nDxtheX90gdD9XsxMEv7o2Zppw8SbWICzyWSWhoqWXQIhch/D0wILkerjMCaD
5GheRX0glKT238rX7Vh6I2EaNZQonADUVQ+xWPZ9BQsZEcD+EAQ7A70CjWG6OGJe
znRFGEOpbVCFMDVd9T9Q6JOYfxLN0LjeL6uURJ4IIUgYkKHjel5BoiGRqZPCAC8B
MfaJ+75boOkVyXUXZ3BJsYXt2nCGfAbz+6zxpj7MMfT1zbF1PsmMV8qGEi0UPsHE
WSEYPxl23Q+9Vw2c5EX7KvwWYbU7GdjOOAo46MJFKyqbTLMCJxzrHoL3EKcP8kKf
hRBdYI4qdjL9coGZT3pJIuk878LZWgQBGpZV8s8qQEg=
`protect END_PROTECTED
