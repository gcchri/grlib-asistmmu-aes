`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/+b5+QVRYHRIeZ/BRjgEU4NOTYtBtnP2bXzRSh0VH+Uau0PhjvbHAu8hTZCgaBiK
kU+CCz/xtJjtRDyXAgJRSzKWTir71lKMwS0MPk4XnqUIvG2qIod9c4K3UTrg6QLN
2Xd6VgITi4f2BhBEz+l0+Lpl4AllAOo/Q3zYiLHeeV0/8RmpJhby8v/0NTW3FE4q
2i2zVZPI9UX3B/JdMKB2JtdPeJyxk1uc4D2SJogS2qWJ7ag+SW1drksS8YxTvCmJ
/tT1YOdV7NlMHaLtRmzqrvW+KOC2uq2btKiTuoHsoYrtHLFqvLOmPo3UMFHLlmIb
`protect END_PROTECTED
