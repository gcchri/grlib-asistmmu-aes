`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4H/VcGIOqG8VjzxlSaILTGn/UfFN08C2L1eGvjmwe4GGSPa5AY5836OoGe2gOrnC
YtbUttWS5lvDzrKFxaQQTx15uDDdVuU2LiIG05bpO7TWsW7w1QXifkFazB2OpHdx
zi7VZ2yPmDxUOEVGI5G899maOdKecpTTU2PzrqZBsJbRBKc14gDrcftdDQZXnIyp
BQflO+ZvULew7tUhNLmyJoHHsEJ2vaE4By3fKjCayPDck1Dpp+GPPzCr3KMyCt30
cR7egmUJoIraJPQXiz3h4vJKpovin/fB8y7SgFu4Yvu6eOyBK0OyqHp+e8bq4wf2
FNiSZBvAKBuDKD7NIxh2kjgR91/47018oXVJSBJiYDSC3vxAoTjvaUaW+jAOw90i
wuJYdQnl+Dj6vyIuyF/jHw==
`protect END_PROTECTED
