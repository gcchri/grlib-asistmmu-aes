`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vjwiDi0s4H40e1zDA45/STXeuYFYmVjQOJX9vVcOJ5kQt8uub13cLeaXY662mDnH
Plmz+qthnDwGgdTINpoUeiFqsRRAc2nvz7aYIRBspSegLv56tplavfWW4//vz+Ex
e9pG7uw/KJxB9fvkdA4M0XeaYXbslbbnjJLq7AOL0QrgMyoAWzpMFm9IVpnDrIrM
Z8kF+eHzIHpRXMTws1F8j5oaAhXQaurqED4TLaMRjOofiC+5EnMVH3y2rcegWN6U
BSfFbr4RsV8k5HqY5z5nbg==
`protect END_PROTECTED
