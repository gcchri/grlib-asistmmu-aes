`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XlJDelDYY0+bn4uZnVlXtm3ayVcS96IFm7KoR5aRIo9HwroZZ8ZUiCtCLeKtzlSV
C9qUuAfTk5I4h2KgYNY6xA1RNJw2GTQtQgZmD3VdgCoxuVNQ/fPRL8wgjNfRcs7f
nzuJSKdZgjvO7bDCGlbW2PqfonGMbD16L8ly99quWroWzZaEWSTXaptUY9FOFIXp
RR1XjzlfZLMgsD6NQPzfVSWCpu8iEcsF9g9bMYK9XbBx2lCbIhb/nRsb0fCI1Bs/
STagSTKKrDuuKNLiVzaKO+b8llLX2ukTh3kbk7VxEptd3lfI12WQ0BOOJJWHeoEZ
ieBJYI2MY8D8dLey2eOol3OWzWX2+nhwoMes9RT+GwyEI4722sxZS8X7nvETL+ZF
lSmKO7aQrXnOq/TfdbzuF8PZsNB3TcdTkiLdu3aUqvCzHl1lrUE3/5HjfLGzF5q2
UIGzaGeNIgppbILX7fciGctWrTc9il7kOUH7esQWU38NtOU8V/nsZylaxVxMT0WH
BZQt/YIHN3UJz7sl7QEBFUqnCaWkj8snfQh9NakaQuJmjGgfPg3VZFi+ituNvfqx
`protect END_PROTECTED
