`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tKxZ+J/98kh4S2tNL7XHOKTaLbcifT/BySjWS6JIP0cUm51Dxxouvf5hRk90D8uZ
jZ3zj0AvVym8OnBxn43GkJPCwR1Cmv2XoxLPw2Cyned0C2ADwWj+TS9IylCW6UsT
7ecm1wVQH+TBGiaV5LoybMEXt4WcJmIx0q3eTdo3k2BOCxiDLg9WVzd++mchtWrz
DNFi/nJMg4HCMF6h6U79HbMFaHKkfEOdYg9Y3SOyMDGNVYsCG7hv4I9ZcxLBh9OP
bXRLQOx52zQmiiv8mPHdBvsH0PlRbYACq/+luo67Iot7dKR59E2bpRNC2NqeO1Rj
Vx1UreDTcRcQzQk2QtuMCtn12sHc77PaiT12zFUb2IiPx+eZrnQh1UWR+fkPSoYe
ckUrprGdJxC3E0AO95MEtwYZwFvaiEAaZLrvVArodIRFOG+nb1oC5yFh1L3Gpz5V
gcQ7St5fKL68ie9a7zZHIv1jcH+4Xd4OKEneBHkdyXOW3er1pp+X5D1S8wwlxHNF
E2xj11INjvrOAOF/ckp81WgLvQojZLZ/SO6G4VYStAYmhUER+6lhwL2PKyLoYwZW
Yp/4Ppz30OBC2UelbWGxUnbx+BrfEOEsxcoVbBFRvcZ5GuIHLRNDbWqz9kSCbssw
6gXxUNcX7XJE0eD4KSjPmCOhy41odminAgUNPRcK8V/HZoiH0+n3AXT9PgYhXTY1
CNTQtmQ3OIVfNOFbwKxZ/V+FKEgiIx/maFrEOkCQqtttNP6akHTQNIUliVjX2g7I
r9irsLmSQ5021OytFoxOSl8BAYLM5FDoLstAWXEEPIA=
`protect END_PROTECTED
