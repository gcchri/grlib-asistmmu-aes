`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5jemzqzmZ/cIMLU0CJsbYj0XT0XcZBkmiRnCZob6yqjqSlFNj2RD1XMTxvndhgnp
dudMAcJtCtsJ1MXIX4qBbGQKN8t5m2Jv1w1cmLJTJ8weV6uTJuD+Mp0IrYbLiY/6
p+I3dB/lvzDHr2PQXmOAKw5ukEo0WFDiZNDA2rHcFGp7JmxbMFjToxlhhjXqFjhQ
1hcQCinzmM6tKefRzlIwjVq6o8e5bTgaudKcdAESsrwxOFcZebry1M2tul6Z4e+X
txbt8JmhsDLfeKbDaekFA7qh53kNFPfGZlkV9hunjDTvJZ/wmldxqTARFZ+4Et45
NxLsZjLCbaM83RWGXrDZt2pBLTs9u04K5s9id3I60AP1Zz1ec7IKyanDA0fLL7tb
qN7QfB7J+RaCW/7ZX5Nj7gdMx2ogw62AdEtQuh1DZa9tKytQBLIe9Js58SWDs4KK
m012g+IDUulitnIF4JooSsR74uMExsHRjM8ArLoqEdMbnVv+H7wu1F8l6DM5okCV
q3+7Gd29+nB/0X8lTtr8RVGt6AsnaAFwbHP7d1MP0fdHCn680KecwgVc27XEUYhd
PkOB2UOVtQFttFu4Ljm5COnEiC1jQC1cXHKJc03KzIz6VTYeHtjrZj7zFeK5D51V
G0OdzLkrKM8uANx2qW3sk6QPd6iJHK6oQOv0C0wNLiWMdK3ALCo8+aR4iZs/rfhl
Jbgd1ninR1aj5aTggRzriVcgCtFiQSji+7ClXpZ4lq0b2riXc8ynBfLOZ5xRFmMc
hC39Eg8tC+F2DffYD8RFIu/3ElvZ0ZAF3YaWp6rWWUJhdrIufUcYiVQMgrxOCOHr
Xztft4v/P4D+PD+8ki0SFec3Yh71nasWzAsVWGOklpIrwjkkCO1Cuo//V8fxmFif
bG0UiBvb/gooHAF0hjPujtBY55v1PYkO10aoIEiH+nwSshNqmsovNJxwmonmL8Ni
82CTikCjmWf9N2ltEJyPOIyn7Yq+LXE71808CChlstMhMGgXvr7k8EEnqtA8iMDU
+otuy4w/UsLergqQkWgRIFhozeOTp0Nmf+hEhlJNko/aAITWq4s8kqcQMNCu8NpH
0PsUVgdB21eznkqJEpC/vKFXk48R+hzsH01D4DQ8+nLg/FyURzvwDHtGbXLGYf8P
9o0htUt9kizSmRpwJlVFN37/B5e6g1xHAJ6fVHvOGngPZh2203Pck1psdD26eLHC
VqPozU/4jHPTbPvtA7/QqBkfNzjIIyZ4ADpnFVXhRJeBXAF9BzB8tvyhlClBYyHa
vIeS249T47GRRbG+4wVzFo7768FT+dvkYQMDAHViMqG95TedOhCR2qtfSDZqHAi4
Ft/W58uuZO0KHtRxZ6wQ25H2BG93AqZwneejcUB4wfBjo6a4DhA+plDeWKb6OCSj
zftmhhsRjz4uiyBGZEaeQ4WNhAw6cfkyPV01OdZG/yIxoGs5+dVaBeL2ETNXKiZz
3mvVMA/dHy9QC1i1aN8X0KOFkvvJxs9g/xbC5HTDQSbj6SaKZfQ+FVZplWj+jsff
k6UU9r4q+ykw0zqlEEn7J/zjS/YhwkBGokUmXTdSs1ySZIvcDP916wg9DG6t5Ro4
G28aRB/GOTGKOFuH9ULCYXpgy/ark68m2KRwLXebx5c3wPGsZWcA1bNfjxg6+hPd
U3YBQzWVSRzK3jvIIjNPgM6IEp3vO24uTR2BBTBRRBxQaIaiPCsUuLJAcwzTkEmw
gmnS+Z+WvvWiPm2T8yEoImTS5TTXi37wpzUSctoRQZilxKsODLOsW/BWhgKhmif2
fqWftVRpyLcQSsLUyJyi39pngK9/xPsZVzyJrQmQO2Kgo232RAZyn07YqPHKk2pE
bgLNGmuij28EPKUFoTS2cZVvD6qlOQj7tcswQ/7NOdf+4w/tTCx8iRm7nItvu0HB
0fD/CrS49sSseWWfWJuf8ttONwov9lrz8UVjN7HeCBxFhyUJEVTNZKH6pmRDQb3K
UczntJOcvTN+qrT5eRy/XvX5wmDOHnQiiksSHgNYupNIoAA/LAg1UzeWAS0yHOaE
YggCb023OF0MX0Mw8GSLhy+352qn/2Kw4sY48VepXtzYZwYO0eQ1WxFMdzBM8pQx
tcUy8yBUj2ZRSVKFy/ISXwbQUT+G0sy+Hxf5bERUrJL3gjHQfijmCuhmAMF8vOc3
hKWlP+C+ABaC09IozyjeSz2Jf/oe+wd0Rr3aU3ju9dNpmVn7aHcU/mXWZfbSVT4s
/jMTiIB5KdWVCeDwthV5BCSus6P7APoaI9Smg6HHmEEalTk+4Pk/0mrLTZZt3RCt
`protect END_PROTECTED
