`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g0XmU+N+iPCkaHVhlbk4XKi5Mp8pwQaUYgk/zJKRfN5zpTporr+mkLUSAOLQuXiZ
60KPOVzwaTbe5KKUwKr1psqK6siKx1du1nfrW4exd0mqFnqv15bASQbF+on2tkuR
paW2jYnevSsz/9hLgha73I+9yh7bIPGUE6wkN4hbac2TxMsaM63rDSIua9SPKUiN
Ji6IHN8wnlOFWVnjf7oxUqRQLYT0iLYUWRMOLFg+urMo7YavQm9cOanXM/8yM0Ps
gzmOvysQ4+VlOEwA+H93XcQUMvTLKICWOAXgSCTKRvcRnVJwg+syS10fCU9Njl30
8NiISvJ/YjUiYBQM/MOREUHzpnBcdFqa9LlMwyctfPdleAv8ZIS7wzPQ4q1FDXen
9kNI5lTcFLdPp7MxIvxO5g==
`protect END_PROTECTED
