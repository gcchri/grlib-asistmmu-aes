`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ibegTU0HmxPheV/h7Jp7Nz4t8pVNZGl8nzCdinTSgiTVUePOiCdzhuX5C+TnLwD7
DQadrnidcWu95lGQAZg8Qgy4jjWJ0qKuTd46NNin0XIYV4aunoiUwOIzXQOiBVxI
Z4JoigsYzlZ4L5GDuFVZf53HKVn0nYj+7vpmHlXcWph5Lluevc4tFB6V+k4dvx4B
rSnC2azvTDys1Ac3++hN+bT8uAeZCtcumjJfdfc0KiW4ZaSDhrbsoIzN7Hy63WV0
+Y+6uKoW5i7uqGh//dhhHkrycTNq9YsjW28XAdmrgTi4Ux8+Kh8fnm0TbRLXHW3H
F1ulsgxJgwcMnpHwD7XBgw==
`protect END_PROTECTED
