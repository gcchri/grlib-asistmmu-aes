`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aunT5kEnozQxCRpkPITHugVcy4FnC5BxSonawTg8l92/YZrvRCNO1Lj9j+GScOsc
VjgHuX4MWVqq8us9Qju4pWDbOhPYEWTWbYw4n4hcwBCZ7Lh6TwAe7I8FaHEvA852
6BFC3bjHcGnslNow53/9EOCnNPlIKpF8txrn5VD6y+rxue9EnwCu358Rf4VbzC01
Kk5AquNLt8FTnGxpDm1bynpC42v2uGLXXyd8uULzPNhybwoutki6ZwXex/XoBwL5
FXuPwTIv9aRHXSE1ar3Lx9Ew7tZeaPnOSbQJx5wEqyPaVluZLOImYul1zk5I0xMd
FKBUCxQ48xOTvwSor4o5BM4PHiHyhBkKhUT0mx5dKoNUENfLBD/1YcReH9p/tBR0
70t4ITOPHB4CTcnAF6Y2BGucnxA2dgx0ffR8coNFKBdSlyXVANbyKOPcIYdLPrAw
Af7RFopRUkcshe931HGDFykCQIp8gC8S7hkU2RDPxtJYfe4Ag+12OaptMMfGBQSw
Nj+5mwcxm9HPDvh6AXxPh87WfmdMA9JTDz2k7VPCUA0kNGTNe0bYu2LjclbMfR47
7hjzGFJgbRRPCd5MtFri5+qtYxiAB2EviSiwkN3PPGzmJLKvItc+nWjBvSb4tGdh
6HJWPlVUdH4DuC4Cpj9l3zK++UuMU+41EZd9e3KyrD/bgks1GRCnuIxJ7gn8GrNc
G+QkGPd+uICK16vxbJAqYVu23GzGTx+NW3cIeYkVn8sZwkLg6UcHGMx8N0l52zRQ
kPL6zVVJF0QwyfRxTTW+XjLJUh1rDEmxR3DuzrHRUhtbd8WNyvuBFB3PYSkwr+x6
hsk1P/AZ8L8T3ElQz95f2F0xpS4z0lCgdFxHzB2r7gi82C8S2ItNB9NsaCqHF7JK
WQLVm6IgrlkoJ/ru5j69qg==
`protect END_PROTECTED
