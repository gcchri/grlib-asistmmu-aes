`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ARq7WyyqSs+gvFwTwOPKVoHFmMFABpbwfE0iwARrnMLKk0E4x/YACMuiWpr8Shht
K40I2aIo9SlnNLCVGLK1clq7uq2BLeLvASpxRVV0tfz4c0Bq2XpyTzLU0C1WLbs9
UHJdU6udorH1h/0ZvJnQY2Bg+Gr+Ol/OxpNTnRosCJp5uMTzYJ1jKIsIdKnoz5hP
s+nFadZ7sq+rvC4111oLWledNQegCIoYKdopwlixvCCPQZC+kub7JyQlwpN7j/V2
wmYr52DR/lGH1URHMnIFfAuvTHXKJGhMFkK2d1Z/kgha9BlTjNJHI2j1rNR5DpdA
ztud1M7O32vza/qI9FE601S66J4cETJ4u2uyutbztW9r9Mde6a8jlKug6j/8QNwJ
xxir/FNbxu4A908rQVfuPhTib94VvepmYxgJs/hyUZu0CQ/jXXljaKBR6eUbb3DE
S/u6dedRwlRXW24e+RY0xWhqN1cmDSmbaejZ8IZvvVHRkt/2kdzn6aoSnWNljLtx
2isdG1UMk0m7ZV75AFS/Bwx1E7OGeBMl0rauZ+enI1iFPytwykBG72874d3E9TV2
f3cOtME73LTrW6fcWJet25xhAvqDSjbxUJ9Tav+ft0xiMSlL5O7bB0ZHTlH/Q8o5
0/elmwSRz4YKFCOjFs4T/KIiDft+ejjsRt+lc9wAqGdM0bbSCAdrjo9ueqNoi+Nk
lqa1t75O5nrT4jTQRVbAfw==
`protect END_PROTECTED
