`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
waz0rXsRz5iUo1lCReXXm0YYO3iSHxGzia87LLPDf+j2P4Z7nv8BE1RHIcgSFbk/
4ETNCqp4wJwlzf8vg5xAStIw4M59McIIY+E27q6l4QDYLPmIjGmXyzx8p8xbo3qk
eOpZFeWv7oFFo8N5hAdxMGUWOFGKhN0n5iv1RHVXp39ICANac766zfnB/G2zVObc
rLXudT/xlPVBhCbuY7wYiOk9pLBq1wAjxerqdiw+BbcX4YHPasArYxefHG24P2VA
BJCaFJDhA6nHxx04SXtth2XWDCzHPm60WqL5PWlg6Wxhkn0Lk9Mc6zShB+Ipa1r6
9A1cxN/hWyr26lF7DO50ZdHL0lffSiTyKNbF2volqva61mH610Fmv29YQ7SOAjMf
4Ico0NGCrm+AfgLnBs/FQcq+0EHu5dHSU5GK7KSe1GkB8n0qx6v3qa7N+rdblmuL
`protect END_PROTECTED
