`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jNqz5fPSD11wG2Z2O08Q+TQTDdbyIswONG6z7armO72Uj3jhszt7dCvME8ND6NjW
A8sM6dXNHxn+/3D7DQsZvEmnw/XKt/cnufceXQ2R9rNoCWdbaDE9EHh/OHU8PAdD
lLkhkVJLvGMM0qBQR5VFQf+8YzFNnAjCSj6je4DB64R/XvDXCqe46i2DLJG0V7AB
IQ0H0vRGUwLGmD1q1j/XVYxyDONkhYI4Ouy7bdkPdgQtKYmnhRece/PgxJ0vYFXU
wZ4sxG5MQiwYHzkLjsF9Lh1ZFRTtu1iRp6Hgxi3P/+xoJxMLXQpMFYOn56hFD7ig
1MNHfQWlaJVM8e48Ift6XbWPLmYMAw+pFeq9mmoFJs4jsrwKYJ8HBfugJmbvAmuy
Tx0bEpInPmB+bd1rilmOOW+wkkNrY7AfJLmT5rqm3ZlS1gMn2WakwQTQwFZ7T3em
wSK/PdwrfLsCLoViNbQqjFOJGaMwzg4OP8+b3Wmu6aPoyfkC54kBfeEqnuOz13Yl
`protect END_PROTECTED
