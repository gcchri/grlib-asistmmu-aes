`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t9+VXwNVqDhRsS0NsXt1RSt9IjUbQbtgiae17bf3T8ypsq3M0YYwv8260Oesb9kQ
VVEu7W+9AgVmbaoM+fSiihLAZTjO0zZocnHYh0p9NJ0lHvL1pOIV/ikrPtDY2NFY
M0XELHpkjfNaI2RPG7rt6JAtB9QJ8cwipbnusfCFrRXETd1U9qYDdvpEr6R3eS32
Y26h701G3BncVPVObGlDiQfB07H5aCPwRGf7DFqThaKKig67lKcbUbTTaDB90tmF
0QQ0kKxxyp5aUtJWu5OUrw==
`protect END_PROTECTED
