`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c7SLs6n63fas4Bcng3T/kp85ED8c+7HHI84BRFurrxA6JNu+d3DW1nljfaytp1du
ZIUySGfTzeRzc42RpsjVosKHwatGxM21mPBoU6znjqPIGi8ZbqJRTnXQSJp2FEsI
Cahe81y6rxA7fmig0QXe1GDCvcH5uCsfWuGQrsudb42+iA4CLTmVMsBYUvyLmEK1
svfsOFaY+gnxXolwc9oyN8exh8XgC2wAao7LfoTz8VYTMhTKvN1mjKJLmjw7a+JD
LyxMJtZm9yWAaZFrUTzQWtkju9KpZWy5vgh+xifvVNAK0IRGtgbxrTPPfCPR22zB
ty1E5nFq/chIdW3vXvXzOjwokdUWA5YdWbNhdcnuTEc+06+/aoYsPRt3OGC1aOE0
74jxbSoo/+NgfQ4hgX/g7w==
`protect END_PROTECTED
