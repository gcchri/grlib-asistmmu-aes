`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fZaJvske0dw1P4XQ9nsGSK78uUQ8g/3AmAI6mBap5to73XQly+GX5kg22c+bGtHD
ZKYr2+QDHwIuxfVc6yF+6s9nICcmbBB/E2aQN5or1BDpR0uix36UV4ByKudC0lMi
GI1kJ7raGPV/1H884UsNFaSn2agn0JQ8XkvutQ2jO7kkLayaIuXNxWhyaItM5vlF
ps+iduUl/pPObCboa+LFiyU2OQuBezzq9oodZytBGQ2+ez8jk8+Mrp5aMs5E0EGz
wLrtelqnOsgcaXZhsptaRdXrAN8SnSaUcV9FUZBaOhCks9eVjma0jKR7HlsgcyXB
n77Z/eIAWSRZkE/qqVhLMD3Wt76+xzyQOHYRrFrj7uRimfm9PtNYhkScKqrdiISV
1shqvGbUpyEiHO3hwWYisEYgSuwbxGnExMRGX3eX4rE=
`protect END_PROTECTED
