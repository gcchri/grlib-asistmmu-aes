`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+CGGHrOebBn8FdLRX9o9RdbP1duqfkH6o4bzoSDbziEXjW/4jiLoMsuVm8LihHRQ
MpWzhLg0Cxp3EgcXuHgTUHbCqb6gFIlOm8xc7c1pV2HcQLD7j73TL3XFinJCtoj1
AJabJU4YJPuETZceysriaEkLxW3JxoJlwof9mtMWyYqO9g5J0X+2Ta+n0xgFd5M2
MGpGnD/1vjNRFxF8pAmFSbpzM3wmg/hwTAGBjfPhN4sJrvbDuT6IG8/yGX4bwXj/
i7Q9rdbC7XQrEswRmf5waQ2dxNOCMmDlSOk8IE4Qx2VYfr+wT3fVVBtK0BZKQcfU
a5UVNIfQKCTbSnj7+70Y/3Sqvb55s9vnB3tDk+kNCpOXmsr3pZSUtYC++UJ0/km0
BqSmoLbJ98Nt1PztTbWkAdj2ZWD+bmx/p7Bm+K873DaaNXHq3NWALEYQi3K+dr7d
0wJwXyLxHGbQz74I4Y9mgs0cAhumnzHwzxQanvyajZP4IkYJZBRKHCuksaCOtjKh
+C15fV4LpP3rjSWvf9CvmI4x7rvvVCoeQJoGTj2bdjSGJn+D2ctbbusawnotlwXj
lENfhq/qDf4npE8XicwbXGfDWILo8laar+yIYjxtOT2Q5ecxxagkuyekFSGlUrF8
593SNUBC0rIr/Y7Q33X2OO3nANGaQVBrokj2RAe5Lgmjp85ytN+hSbuc5ZOLJwB2
ucneNSgJV017XNbW/vb69ylX2l5g1M5Jc5Rx/Ufm5YZjLfc1HtG+2Kim36OVeMzL
fwiaZlgPzIrqIDox5kJ/0FxD/YcCVGuu/7szn1gl4ooSHHboP4v9Mpe0rp06U5Db
JP2oFQTt2REpvT4ms1EH0N3vyx715G/jlrZJg8myn6PBHRcd5ICO6lqZqhzjtYEg
MhLK7hqgelUowA5DpbKwNq9iA6RL4vXYt9YiQHs3iT80qKp4zgkYEG9AbRatgqZ6
aqx81HRlbU6pj1j5Is0RoFZl/RRStv7kVwqVYjMnKvLb1w8qb16vruZpDLYXLEKP
mnJT8+VWo6z7vqvuE0OZQq1fsIX7VSx9gundyt9zOwme9FnNaOSfbPqpSCwdLhcI
y591EPaKqntrLORf0SVkeGQjpwldUZebfi/U1+3dun7m1SZCe79FDyrj8ztVq5IB
Cz9Kj+YmOnMU04xhLc6aTHC/RKJi3UXE/BLcQxMPC6VmmXoiXLRoJszIA8ESDYQ5
`protect END_PROTECTED
