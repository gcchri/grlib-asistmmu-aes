`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FJajMGFCnRFsanJ50pjTzjLDZFE9VZeMrh0zmb+ojL0ZHCSV3t6b4yIICRXKl5br
jHr9d4Q8QE6S+UUEkviGOW630Mn0Bz1ZMZjxwcTZs/7M7GxSUy9xpdApjbkukL94
vcWPcfIwM69cAG7j+oOfOxR8jaE2cyhlItAtKEE8QlyevDrdexAvW1BT4l3GVYfa
HwSGINygFVWilgtRQdX4O2PTntb29Gfxl9xPG1FxQcaO4Bq70AAWOqvsytHIfgqE
kEzk0EvpkJyOyD8PZrc5RnrwXUlnJeoqtYPUC3okDPme5wuvg392xSOHy/ElsqPo
0TpeD9n4slZyOC82FVdkAoSHvIPjoozC/cpyj7Oc38yDU2mmJDxyMuRt40qwUSF6
`protect END_PROTECTED
