`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kdc33RlLXLmUC6NGYpf0o2tFHto0en1IXJZIaddbP9n23be0xbiaemIifS3i9ZW2
yh5Q4JinUzlTuypFlgK81DB4Qs1q+Y5buIve6QGnSQFpHKYdXONiNwnXzcG5GEtH
tvJ71zgnUP+n89Fb4YQR0j6URlF8aYsG4EuN4+zEOoV6uuWKUqdxvloQHYvKTPo4
31S+oJErW1LFp88i2z8Y5rc+77Y4u2X2norBgteD5b2rXLoqx8czGzzQJUHilJ9z
OI2oQKTiDTIstt43hgLqnRxLQfNo6Wc7fSyYGFQdqGAMPj9zcAaqjp+3VFCrrGIC
rJRyXh89dLOB5piF8QkDV/kgWwRPodr7ZehBM7/d3IZ8Ep/xjAsjrRplSmw9pGLE
wPpNp8fjhSDlRyCI+RLqoT/mW+1TAgx3tLBE8uJT1Vw9bRImCYcuV8VkJgjEsTfw
8M6d+63x1mHI2qI/w2b93Q==
`protect END_PROTECTED
