`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nxVqq/U+RtrKneVegd5M16ABOW2bfhUu+Al54h5uyL6sBNQfM/xqOjy1k7VJtz4Z
zdWQcXLSDlxI2GdLIP1q69DIm/uA9UrhSgAbGbVndcLfz+TecFblddC77SurfCbe
c271OIiq6V4S4JJsCndpkDFKt6QmETwtP8HGMrJ1Qp6JMxHGsALs7W88agxnTVzs
2ZLa8Wcs3KuMEC3rZB1SHibmdHXNzhsDUk9wYszFgBjZTiCV5sXe5inTfQawlm6W
42qwwkLG6y0nvEn4JFpWPnaR9HlpfQniVVFUfEFHZDMn3/teMBBEXRoaP25MlJfH
s4MedH8FHaysaV8+Q1nL61chigSiWuhNhzg1JVL52TOaW0aQ3C/zf0G4WnqfTI/t
XYnzKwt/aSHGzLXYPLfT5HK2IeNzwn2q2eMijdGzlRsFxDesr52QlfvAVumHHYyt
`protect END_PROTECTED
