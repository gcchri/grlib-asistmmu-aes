`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Skld/07917z2H/pwDjZfcgdwJiMqyYtpzeAGuOuTVIX8m9HiM70kW0+evSTY77kI
nRZ9iCjS9iR/SOvdViz6kgKC/bdEU1csMB1d0di7DdC3fRKwQTqUviEP562lMkGi
FOxxAP9b3UizRNU82kK8LlkOU1XmzMvbcAXlBw/iqYJyTJX4uPnpNhzRjra1DioG
NDnjpxBLbMfOSMoy5adrIBptFikWlQVf7L6cm9JkDJb5OLPwN7IxeKpiG5LCJ+2H
X/FGpVbye1Wxkh9PpwzkxOo3AQJT0XEms3Se+q5K4PL1QdcWnqJVyV0BI5Ckwl6A
ReVFeTLBjfj0mNcx4jmvW5TQLGiZ92vN9dy1D9Z/mIWZt+4zrs81k+Sa0M4/YkYD
B+yrUwN0TPax0sA7tMas6lwoeqE4uAjDsSAT9b5BV6ZUmwp3e79gkh+TUwmWBwaq
nSCUQfsI4jsFvzQMEWw/oMnO5PXTvxVsjPv+jJNjXDCRagzQLRMEmYaZgoO5pJS5
sB3M7kbJ8PahbZbT0mLU9vWYcJmsZj6kz+S/83ReeemJ8/WINZ6jGuWYeRDbjtU+
EAJIeT7vJOR1+bGFcbOl2K180ubWvU80ZiYFNUR9viE3Eo1BsgvoAjtJi+EBSRFB
15lPQZMUNxvaDXMXTrNuJ41MKZPKucu7dYksuDsPkHe2PvBgLcANn47AjF8Z3f9q
imhio2oCJFlpvi8aLM8hrEzmfXb13s6WEwG47CNpcaW7rPe1zX3JuodifRWNd6pE
BmzMsOYF8NF5K5fhYJUz/sfYDWk8etTkFvct+cXyiUwNoGMhdG6czH1Xq5aMncrT
9ZdWYDVRzPc4vkS7MtWJqEAMO4kTI+9vmx1xOdzriq0Brkvl9KlLQoz9S2jwXl9y
KrNBAaUX6Kf0bm99eyluaK+iD9yi0POuvGyBvRC7n06dORhYEcjwqVBnmOkCdCWw
tMx8mDE7GrZuCkEz8dbmKMPdjCI00h4ohYwyaJKciXFkTIjvv6EhxWIRYRSe9due
6TsUtMjYhTHs0/zayo1vpcXwOrszQgQ2xMkqzSfnyuGBjf7gGaP1wCEzhns89cF2
aIADiBYbzzS8IP6tJggIKLfNfNZqI/ZFsBTpNKJ42BIJkPVtWxFVZ23Zx1GnvPLH
BShNN1zb5fMUF4AOMmhyaCdb51k8LQJxDdIny4KkNt9xmFkrTjh40scGbQRx/WkX
rIWNUWmYEYUapTXODdaMsePPw5fjP8We4x+5zg4H3F9clVPFmM59k/uHaH7giqQd
lvx5LLXk4EpMYpgtBpOjgMc8szOtnIMsXRTr2xQcMAWPqv/qyENOzv9X2IKw4Lzf
HT1eMM3MJJcKdlIKhi6rqXdrbsrw5VtJ7e01RCS5zqaO2uYK/lEVGXSPmC7jqZvf
Bgz81ju07oIFya8xj3A8zA==
`protect END_PROTECTED
