`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8MoAyduVV7YFEs6c9f16Ecd4rAkt9k22g5BjyIAlRdU4nudDqpJIp3eS6j9UrjPo
NnL6fObM9otH/OZP4giyR8kNoa9I92yTDS34qA5UbrHKJEybJamvxFPFXPyWKB/M
KU8K+/tvHWM9rAuYUhvlwQ54s4w6Cs6/cnXsQNWrlrT8j6MsiXIMFEMuFqndK6yo
GPqfara5UBZaT7eK+wZqfTrNGzj121wwMwgb13N3nWtXVAilnFlglONeOESfSz8x
VMSUhRBpRxy2KWzgF++xlY0rZCL1y3meWXJiowdwHWrlWeamVOkJgEZKAU07BkH9
kFT7SzYgo6b/VSXnvX/BO0YULPa+6Q7IqkXLyedZPVbaFzPssc5AZnV0YslCMz91
dmCkWBAS6wkt1w1+PUj4SGJQ7ugW6JwVkVHBB3ZAecd09lKn6vw4OEWuqLB3J5wR
9m4tgjK+eRAhZn1WISoohiyX81YoOvHCmyAwR8y8wR1EBDy2oSS4NlxtxZN1EmwV
F0Z8QqAGA76JHh7fDrKbtetcveE7nD4QXna3UX9WmIRvSdZ38gYlcmw+mB88DLMq
gr5m6DmW9h+lLjXOiWQeo+9EYJbiZwJFrYJ77TJKgXBJrkoO7rajq5RyETtv2x2n
hUr2h0XQNprB60jLgcVCa/v1C96jB8k7wMvqeAMGFq09g98fFZzNLBlT+Nq0KLXo
tQxyVpqmkhia8IcI4/7FahPmu4H0cw7bUT4nOME0f96wSQQuM84Ju+f0llkZI9wR
vM+PE14bL7xT/8Vi/8ynpsx56g6YiB677tdVFIZTmcGcLG2trwHxAeDi+mT26qDc
DTciRT+dDhr5wmJDfK14O3hicyve4J6tpGgNkd1kVz7RLDNkuhTyOYHd/yjQC2o0
h3KPGNHqI9p4N9njJRyLorE7ehCDOFjuV+4GfzePAts/BJ5zJzUG4n25eUP/W6Z9
6BfPBi47m4mtMRQP9P889U+dZJbYRGnmsYdy66gEryCNlLfPsk5yR3xI74UQ5NBp
qAajjwd4dsV/lNq5S0AsPQHbqflaCHKEP0hGkXs2hCiryTCXFJvsQaRs0vY6pdvo
v0yNUWCtmJkHX0laoJel2dyk/CQyGXRCTO8XqaE1viz2GLgBEpD/n2au45DwpjUZ
09VO57vvbNIotnYcC2t0ST50OHeko+01VxzyO720C+42O7wJt9UsxfPrKVPVW1Ns
hfLve2EriDYb7Ro63ttZxf8GlDOFcEFYKTMii6XCm0kMffgpZUjs1ZbDvvxaCqGH
FLL1oKamSftlPNfWddUsKAo5eAzQ8t8pk8Ik7ZIXnM/ZcsRIGq+YV8DKRhv9cWPf
Z0gCPazbiY3cqPorlsgmfXwIqi62xbNV3GtM0SUZuFk92bpXDDFxNlJ7MFAs3V5q
NYLnDPzd0fvRNbS2BI0+R+G4RSo+r3OhUdnuoI+ndo5NXBCVgkleYP3tbmnah3Ux
KB6XiCZ4DyxGApPx+o9d2/AGcXAb7R0fYiTOpO9f06Y4ed36bF/5LRBTrWxyW71o
H6bu9C3HCF2dhGYtkpAJ/mVnvn6kTwkH6HXYwKca5R5qUvetyuHiShjoEoVnQDFy
lXvIQShcBDC83o0req5CZaxtGhrk4dtVUCTVdpoJXvNK59zY68l/qCQ1nK2rRSpl
PFpsLzuv6iXLmOcyk4rtP7OsmvuYVkqgJEx7PlMA4PiOQ3rlOE43QHPJzQ+ba3jP
D2xc+1ADfP7YW6ltz2qX404jFDC2eiXinnO2yekIzvD7QDI2LpQ/UVtEt4MylnpN
XQnipdPk0P3thFXImQLTgAlY8RUPFVpNZk7piqmODtxGHNe6FTky4/TEb5/yG69K
5U1fUTuO1kw+L4i0az/DI/VIWcqKsuvoKOtZSsxnXEw9vR9TgUs6ORuvCM1WY3MW
8Ncf0KLeNPaJNFDTlJY9uGWlq5ysI/yKyjWZvVDaH2Xqry/JTAvNO+LBUVrZ0HDg
znFfBg3FPDzqAat9i6LY2NFcJkPayHH1VofGI5chB4r6br1RR8LUaIdiFEkLdQx4
fgnFiQs0Xh/mUqmPjtxjxjtWDpIRtYXr3JTI9uxlvGoW2pZlkok5begA2hdvsqHN
rb+lDtszTaW93GGTfiQBmi4k3+HHZ7IsBzBCxmSA6F5sz6RelERQopo3PoAFIqom
3O81d7GomBzG6UwVpZVbfwBy/1/3amd0d6t3KoyTBqh/CX7Q+WZfM71mZ1fI5Uc/
cOaVV7Ba6fMosP4di8axFa7br71Q2fSzKfCniX3nWpPSVwu0HxbcWedrnDAN84FG
bcPlt8JmA9tXTQ1T/bSPvt9FVaTCbbLmHqs/+We3L2JOSjUgeXNaTd7tmrrrW8p8
1Q0jHSxfjNxookXCwZEoOmv2b5IF0OYmwSyFefVGIFTxJxZbmFzaQmgjZCddNcSF
0JGy/qlLJ3N1on12fhHpXeJ5X9D4uqoPVZXrGBVbn2tm29bruiTHBMcxXJ3UuIV2
PyTdMC/hxt/ML8awCv3ZFV5ifd0rrSM6LnqnhFa2Ooxji9s1eXQDd8to5wmQRD/E
2J+Xr25uxcB0RtOTkvCaqwwn6B9YgboKrP+uNkhf5Etxjnacs+A+W0ms3vWNarXH
fij2evZQ7b2Cj0Goh6qRlNy8SBDRvDj2a0xVtwYXRsEgo9V0Levhe/6phjEp4W+Z
r2DAGnCPhu6fLXxkhuMEvaPq0IGw4/ekM7Ht6jdZVxHpgOegYxnJCwzkVBoyIJ2V
/L/DBr8fw4qd517uQsGu/e9aUzzR7Ej/aYFfLJ3khDptOph35xCY5f+eR2jMCLky
Nz8L6szjYTSrDBU6hiTk/s6GuAu+SkJrIbA//MLC3cviB22GcEEYGY9NvtmPiclZ
cMlPG7s08L+pL97gUuZjfRV9DOfU+X2qcUpm6u8DW166rwTTvoj1wTdFuuvx0g9w
Z4iFZaCvAWFt5GhfgesMfQovKC11rEuejCwb4CUHjAb27mfcGtTRthaI5aui8kzu
6QE+UBKDhBQZtDNRxNJha1DG7QIORXamOv0+2mk6dA0e+zyf8shglVqNBbsdPew8
hA7AybMTvUyEBFSZajkYCh2Emzl3WASoj12ZKVKEWU57ycNWtKVVqQ/PjBA2z1xb
NS47EY1OOTPi2XWjZfyWTP/IqshB5Ol9m0FxBcEYyy5eakGGnVLnJ578Gyblv5ey
eBlLOg0USQQRR1Q+oae5r0FQSpBFcc+V/DQ92E7wPNPMwNjMK7vqUD4eXCAS3GLn
g+vYkFS0P+IV03ZI8/f/Nb7NY//51DPvOA8dR5kUex45m0x67RpcqHN0vp9uLwWX
zPJERdQWOriCBgrYLViE2KYbMC4EIfbamwLtJv5o7cQoDlwnpa8JaeJIj86tzTay
didzj5P0L5gxIxb95wEVtnl2mVbhFtyEOmr8ucbbQXrZICDmpATN+RDrhvPLIe9L
5oUU6RhZhCqJEQ6lgefA6bLpOwRWjC1Xf84VOUHLif3BsLx8/HD/05z6RgrGMrIV
jlE3L8SgtFwKWaDxwjvoFTCbPWqMzB4tk5oyfGW+us4FElWsLIGVKpxHNrfos28+
jRN4wCVXtk6yodNqF6tX5434wOPYsxs3DZkjRu2D/Z1thwMQ8uo20Pwa1CvaqUkT
wGBZAy7wP3hUh339/b+b3ZTAe4knSzgVtp8pECNTrfLKPpZb0+gb5FqlMBi8sU/H
/DqYGflO4Gw/3gBCzEqVTPmyb0Q1HoaWzKW0KSf3DKdrXQY5d+eTLWok/tkDrNFZ
E3zWuWt+xMWtpF6D7bc9XiB4oT2xYUtCIjdp6G2e/PhztzxltC1U/nVj8EThytdb
S/VWACV/7PtVE1445dQcOezcGBF+20omhv7wXdue+aHtBCushzLOfHDtL9EDHteg
yE8DDSfgHGdmHbOezfSopqDMmGtrOIVP3+HMRa/IBWJ1jmYdPBUZNerm+BbO68H1
xCQOKozQUjj5I4D0dTWlrlXfJMO7u0KOXUsttkHmhqd6UMRwXMLk2/qujZbY3En/
GzgQW4I8suTA7hXiv6icqkzTz4GrPxOaSNw0YiA4HgGRCaFSZ7ygL7emSYvbKN+P
OEw1vUDxQSm4sDGpVSG9K7vKWIa+CIpuGx2O4FiwRysUCIUfo/GKMNdUJ6GRfxsv
0eOSMQIF6Jz2MlzmsDlOd05NcEOv0ZJZ1FKDVA908tU3fON5tcAuTYYWpvjeRj6t
qwBJ248hPqLhJPcwp7YWWrt2TNQMtcahUMLU9sMnhifQ8bUJxm3IjLWer6Je7+D/
2gcYMH2Z8eoQMB//zaaQvkD5SpPLwwnOqBrluiW5k4+M1rAR4BCMA2ZT0Fk2sPYd
Bof7XaJEWDubfWteB0XlC0qblIAEywczyveHlw3HyGnjciDyVwPHPdYyh6/2qkYR
1h9PzwyFzcpqAOEwauHS5Jekcp2sxYjxWSa/JQAh2UoqIMb0MvwvAw9Ws3m9uQ2Z
bgctFbMcuffaxqMhHx5CPXKi894k0fVOUP2ns6fhMO/twhmTH1Xkjv3n5TfyuEAW
VYwReuJpMKyxeVuoVnMR0Y9gttyR9+WOcMyeTMhFMsLcRiHo4smfuDhEClhI+1Jj
abs3szA93eqJnXw+NfuYqsBMlYv50GO19ynUJ15d4pTId7pw8a4KBRDv/go3YgHP
fcuA7e1zMV4BAb1voJIJfV5if3O2ieqyJD/S4GowtFZhaFLRbnrvzU+zutCooyDw
/e3MFVR4af8Z3VmVIfofWPnI9PPovtb7uhciX6/5GiYPc8N6QTx4c9NurXz1tDP7
+Bw3mKXS+3pctIL0m8W4wIA+Mp76DJ+a84cH/LkJkDQ2J5oJhBvphK/sFMV/2zQe
FbyA8ZIHBKdAgpixp2M9H6snHrsPGcUbvSSNCxBj6NCrN3wVQRex7zTsTEjoJrGo
+SkrhbLgPOHZ3PuxzEFayoGZCsoPvLBaebfAzREK/hbCia7zWCzHVvg8k7brFQnz
9/XWZJ5+rj32hq/uhdOLjdPLbKxqjJTW3tQ4jHkTWj/7oULDFmgPuFJiL1PIIGJm
D3yraisPJlzd3olBdRGoR8WLJiVewO5DmPatGoUT2WAJiwCwl8BssXu1k3hf+w6h
nU6dXJPohvsg2GL+jglPpWsqXooegagbzuKSkdC8Z0KCuTZyqwG/NWl6+nYNNFvv
Skki9RUWs/KKM49M+70QH1QxOLjTom5e3llly+VXNilL9datmddN8UPD7VXUK0p6
wWHjcmkqkCl/DJCR1NjVREAshrXwMZZxv/VORJtZy943iO2BpDyfHgViY9FITEMk
K0O1qc2K2tPbPaYbtaDpCcuCUpnhIBjbR1bsvmWszpcHBhsGDqTM/G4A9eAil5iw
J+T5Nq2yJBDNl3+ZcFgJfYndy0XSfs5WR8+8+F1Qb/I=
`protect END_PROTECTED
