`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CjwI66JW22ZSQhGA2hape+/nHyuRMObydZ3XO47FRYObt6UMooNQrsIt7WlTM9yx
sCGrHmKg8WVze38KDGJJD/NOypP+ktj4g/tNEOF33B+abXaLl5SwPdCPk975/ASE
cDCN13yjC66eDi93SxTBFipj29lqhBKnqfI67aXcBIl3hTvLPMUg7a0gR+T0GtUV
caVVeQJC1iPyZtjhl5ryf8DbCzuVj88yynytGAEa1rPnoo13/wNZ6qWkZ03YKVHO
G7aRfYrNzaGJmHDabAqsxo3kZsN5L2238duoXd0TjJs+x+FC8SIlqZFYNDphHypq
f9XeKOoY4glDSjJqoJvSXw==
`protect END_PROTECTED
