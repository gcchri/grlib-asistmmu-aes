`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XSMtJhpnxpj5bPh51IJLf/cKgP2+ktN7tqzmNLCTa+YqWKJJ9jqxkw04zB0XCV/l
/Z3frvqcPfI3crMypDDDrSKRn16ahEEYE2nL/igdDyekC+urcoEwO0aoyuJT8Pjk
+8XqvlFMylVB7vT6mxGaU9N3XoN0ClmBfDtB1JeHlp2CWlbooy71hLV6eex9qIfl
V7yqaFJ8yz5r2d3udCdeyPXcB732U7yhQ/txfEYzbnzq0ce98kfH8CawA98xjpc7
T8JeMRZbBBUd7876CyuBnVUSBoq2KZAbYIFT2VTTpII=
`protect END_PROTECTED
