`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kQlzcKCljIiWUYXVRK/eq3RKL2oadYLjd4pIS1DCBP0lMXDCImqN4SuR/nm2/F3I
fiUuIth/VRAwgw8QxdlOzDouFVD0Bu20RGIKadz4DI+/dghq4njGsc23JxUEDVOI
82fErTin5ZFqEVsyTfpUPCTLevvQvwlgjKCIiYQnW91DCzEOaAudT7qMxF0OwAIi
GxT384Ax5aPoAc/MgcX0s/I3tno0yshK3AmCBv1lmLtcbhXNmZIOYyV21wcp/myk
FgksktR8+SJtrEx2Xn5yoC1PfUDOdXppx25ZvbbHx23cwZYB3nvZ0qhg0KCIVDHA
qbThzrkBUE5t1kY0+KNYKVuhTS2ZTekphxFe94f/9XscUvTTv9gGeyAyoOOgbJlf
tneCx+/NnyaUJdhwzDArEonJLnlJa+QUQlv8rG3I32St4SzwII4olHSpovOdbAqd
HAo+rCEmiJpE48ROCvO+/Ovyt/ghH544eWOqJN51r7XJ608Q3ZRSh7PkQ/60J7Mh
VDcaoSfzFLiTxg1eiZ2f/doyTLKher78DZ95ARtZ/wLG+V6dmrzmHgHetlgcf37j
GPNfORb+m4e3B2t4+kXZ9QxoLFugJcAewzfk0+33DFrnyBjPHnnEbBvqbGLot6PJ
j+6+by3D07oFCCzbhJyjqzAA75y3PLntdriBCy7sXeadpXTZ/FGzuPVKz5scAIXo
9ywqwnYbaQdonwQQKNTZuA==
`protect END_PROTECTED
