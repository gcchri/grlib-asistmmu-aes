`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NLLmLWA4fJO0gdZOssnvlzQK2uHRWjrRTQ8pfV2Pd8SKT3XdZSbO2w+WOU2+2Glj
I08m9RJlyTSp2XzVtM0QZceBJHGiZ/dGkOJ9XdCRF/sV4VL2opf2miKKmGjXpVh4
SMLjAjonG9+i6kkRxlSNeDz71TQc+145kkz+yTzNpXMZcVYVe7di2k5EjCzjI9QO
dvzHDvj8FJmV4jSMlePA6pQF7NCp0ccE///D6Kormg/xl0steW2fcg2oA7vxtc21
lE+/h/2ywZD0SFR0Td0IC+rflNBdwd+y0TpfDI8BYXNEv6A6/1/YgNRUnWXHUShW
Y0CZyGuBPfLy8EWL61MeAgx/M2BVO2bdUzB7E+Yr42WcLMbjuofarrsio4lGvXa4
YMab3iCc0Voqom2unMyly+NJ06mPkp9WDoapjEDQJwNKmM+Ha/PjugseFJt3st1T
eWEug0idgCuUSS3x7ZOa2WTkkLq9TNJXu2SBl6OS3vEuGI+G/0ZHiRChg/ck+5MJ
i/d8CzIX1p5eIZmXhJlE0O3lSTv3IfWzSAN81bkayZSUlRblj3Kh3PmikHNPcxcy
mBdE+zRi2UjSAE/3Hf8HbVt7ByFP6/6ZmNYuu/lhlqHVyj5dwN+2aAB5yBRshCoO
Qx6NpaDO61ZNu9HLmQWqlWB2JaMGhun96UCFu5Afcgzy8pQxA49Jqm+GYKDlpTZ/
jV1oY1dnNOuxh/88iPo1zIDh0j/KHyhMjJGX46eUFzFaaBmYsR5AEWmnYnCY3nyg
trq625Z4CnkVr9QfdVtyXBHI8Tuy/647dsBJ01BfbE7hMK0ySo6Zv4mbDL77y5E3
KitbBRkvvpmJeFYvxxJr6L7j6+uQyMzob+gpqWyL8PQJzdOwIcqGQDo6ZHExq02F
I5+SfT7nNHAzGmlOx4E07pq4+IyJ9J+yACfgdSqgPJbC3tohJH8SX+r8fpkq2yU+
uzzBPospJj6x1/hsaCr2QSyfz0M3/y9EHuuaiwkDHRQfutgEhUdDpsLQlJjwRvX+
pVQrZ7Brz4BkRjThHAw1JIxBuCWlTVD/3RTwwXvM+qxha11m15x2LT+zeJEKTHwh
uHMZpYviPF9+EkDQH4fgo6uRCNj2MoNrWP9my6cOlc/PPJG7aH4hH33k6Sg3s19e
MI8aLu4X3LZZWFi3ToMolfd+6JbwuGoTGiVTVKwBi4t+/kacXzd2yw0nV7c+pc9z
+4WFHuD2+rxDPN87HPqty6jnrCmyLuIMXDHKI0gw9+OnioDXb+vkjwkPwP7ShrHG
6J8oVQZsrYLakBwse18wQfW+wqGwWWQjRD2M4oXpuV5KK+sYha97AXUNwqzsfIkS
C+epXAbtadq9TiqbtvrO0xBG99IXUMxO4NFmJ8qDGekz/NUFBo87CqY8N6DXuM2o
YFzP/LdT23WIM2+tQFbqCb0eAMAmERq5ZzsLvDUWBwAS8TW545SBOCJsSy5565dO
Ouxr3dCQJ7y//Z7GjTotPE2IY0FcxMIhM0nr2H0R+XWXuqQyXnjAMQcguh6ql+cP
46XYRp/M+2UJ4WDdm8hWXktxq8u4dqCnYi3lYvu/yw44JgAWAMSdzhmW3uaKpPbC
md5YotHEgUqLZmQNA4TpX+2/UvkQo1q/S94dyK6K+OcIeVz1h3lLYjaREU7Pz9UT
GevBEfdgW8TPJxi/D/BZElrpHeBsImjI1R9Mg+VLbtqK2rBp5jF8I4l+UO5vdC2L
u5hS5udk20Ro1d4zwYKO4lWb/Bt2P9Z7do1wwbE8TOQT4I8kMhgQS9PDKfGRzNM3
hXiRO4CD/NNNI/uERaDYwOT3iaJiReFTlhkKLpsMJwix0CR8roSM3/pj0/a9uks6
yJpPRw3CsP9i0gYXjB9gjR7zrHIuTM4jQEtn50KOOLibytYmHVJ28EUEumCipRSv
gW528SXbw5u+jKeNN80QYTDTefxjkqc7weJ/ek/xoqqFiFFP77ZB46zvJwI19CPF
y5okPmLiLQ9SoosiQJajHdPMqEwKUEvcKXwxWhfeJ4HPhFOzgJ0pZZFh/qRMfwT3
Es374aZ0CTKirDjpx6SaC6L5BKXq185Pm05lyis/6QNhX1uA9ZDyJv0PHjwDEDhe
ydUGYpfjLiSRkeT3lSyIqe71/mawDUPGhKUG4gYljLnZu2mYlpd5ZLzfKyhl+uJV
q3Tn/5XhQkTHs0achCVDa9ETunRKTla54IO+jOQBnstKmIdZFt8edJqqGBEUBAPD
aS+vBhNe8qfe0Y0HGz6ItUwOP4MjihZEyaTItfJBIki+yPG60fFUupJFVsKffVo2
9JrCxVFVDN8otk02x4ZK/JTpDPx6lo+84rgQOheNfSSDWaj2KpzKK2GkWqUVng4Y
BRUy6YWqOEk552Q6anHZea7tOn00rezmqD1mMbWpAwcEiVDJpzZhjhT2xvI7SA32
ZlCHcPux/WXVI1D5LJ4m9/t+bMVL1um2Qvq3ASqaDQ2Z3SIs3U7FP0G/D/bL/qMj
HkdUZ7C/ViS2H5pzh2XmQi/8KGNpcy1M6FqwXexV8wAWjfXjhscyWZafe+H+v4ji
BOFO1ClKu/JEKB0AyZPj5pd5iVu6xTo0EF3OD62OCgKo4/lutOgGcLj0e4GXQyqg
G8+kR3GBYDZTC2/aK/CH+t2+wR6biy0KGjBHc5WnRll/M3pI+7enW04L//lDw1JZ
/p62DuAI8oW89SDFSj4wDdhT74hqbclAWavD1pgqottRN66gj7KJtWqX491ujpAx
tiU1FFrsml71IgFIhs8VaejHPEzBsc06qVpC5E41yVOV5ZmcNOva2b8PpWJuLVSi
p7aBpgO25Lb74t6IBhoiI95xqfADanXxiZ82p5XUpFGhEBVELP8mLsdoVpLHvVXj
GO7uAUM9h4h1DN7Z7Ht6cXfd2c2Uayg9La/sFlB8XN192dJ4yrtwQMxf37RAYc8U
XM37xzZygh2gLyfUzALbOU4Jq9Y0dm65n4oJU6ljgg3TU060Q/8bXYkNWPP2oWLu
NtC87brj5ZzrPdLS9hzsqPlEwGXhklF8bthdEorncHlYAbUwmKx3jdeEaFPS+H72
lSy0zExswx3xV9UA9xwI1VZpuOQrPzpsQGVUMi8Dpyln+aKOY0uDkQKIrBnTMzRl
JX5PLmFVEGJlARug9cH43fIpUyHgUghF2dW1IwqRsQudXa8+MOOJUxlYSvLge/q8
cXofo6Dr5C363ljclRn+i5adIKTelTdpMHnQ9tJbCwnxhjYa+ul3znBA7rrxMweN
ivYubjEp6IF/b4gXZSNgyfERjxV3mnOmWix3yj+Wp0S8UMvdjxLbUnehkeIE5+dc
CJ7Hf5OGFEMk1R/lERInAojff8HUamwevYYn5maQL4exki8Mm05YAg5uESpHEqUe
SJnAoFHzmMkxGMaC++KDFW9KQvAPC8XTojE4Vcx4XdsnuJHOJ558M2fxH0BjWdQq
F/Y5p69hRUUYdygDDpRZRY7KvExMCD2JprGB2Wl7fds4+ZWRrSzfuiQ9o2uodyVl
NGkxQR+q9yq41VrCTZ4mTitIQbqb84MBMIoD10cwkjM=
`protect END_PROTECTED
