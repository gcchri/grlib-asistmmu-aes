`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
12Tkc+eLAgX6AdFZfSzsapiiFZMYzht7eze1Kr9r8ZSQE6osEHjzpGclON0/08j1
yrVisNBl1udnOH2GytE31kfHTDDrJfOzHEgWIqAJDjz/cyRDn2Ks9eWKkXzAw5Pg
tgLcQHXGYbulrtLRpUQ1U1vuNOKqPPTkSdY9v6h5LOLz0toVhIjOyflo1vgLbWDt
kPXK9n+ETKtm0UlIJFApvkvXfxuNX/RdE5IJa72AdYX6MCd2B+fKekYBt2NzX9e2
oyqeX95CChuyU1J3yH4w4JVaXbaNQkJIqpkDpNd8xjxk6UhF7nT7FlpkjoGn4WKq
aIsYQ4Gx+K+8/yp67uxzPg==
`protect END_PROTECTED
