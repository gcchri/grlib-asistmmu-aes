`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BAoCXZMN9+/RnZ4t3G194kn1c/jBuKj+dpPnJvOXG5VHdBvtKx/ZuGOCy6Q54n6K
M8QdYiP6WogT67fx2OduwRcjcPZgnhYHC4RJmcjih6cri7TRot/XoQSkWejYatdf
iDUFr0ovoCgBtjyO8aDKvYUatprH/3rP1BXfGRpovAHq05qV4qb0etiEM7ddvD6v
k6WJ5Azttt9yle6y047ZuSOR1cX+/P+f7RBEhKFgtjL9TVhD59QL4R1yKDBc8Eqf
vPU7DZdrGbecLolwSc+3pzJQUzf5Yu76j04S46718cYXCdFozI941+xnyvvfWNhI
vU3ZKo72Y9fgNV2m3I0FYd1SvjYfymOw+QRhShdKZfbGgmO1BAi/MqJo0juX1ieY
6eZi15G9kmN9iv/sdEsa1+CjYvXYX3RmBVRjZ0DgoRa5JbG5mT09qIdhxdoEH+2j
IlSrm12NKFEiuoDpt1qSjOkoG+Sv4wv/5EHtr6DbsSG/RDAv5Rn97jsWxlJpGhqC
VdiCm8xpTgvymxzpKQRWQdB3jlhVO/LRgJLeSqL2/wXqnWcwWJc2QmV2cwvjjpxR
sCXuYOC+UxgmFACl1hSAE4lE/+j382LGx9hWZvcs7qB4S8xw+5WFuox2J5BtBdwt
y7s9osPNfafTbLxQySXqZAp++QaUq/e+8I8VsbNbSv4Hi2JDlybTbZ60uPSa4TJP
czFrMmXffhotovMByk6RkjEp7WTi7oh58ooGatZgcjNchjB6ChFWQLPvW2ZU8368
D/tSljNrBgN9TIWdb9mhfxJFthIq2/BihrV5qC+eqF32Y88TBl3kao984c1m7xmh
91sFbb7zt+lwQNvsWEUxhZCXOvxzezymoD4QbJBNldTlgkNrUWwXIhFi/FykVjNe
nOjkY5FSD5Qk+rs8YJHtMxz3uowqhC2m4/vDXuTbBUMmw9tKKYACFbYLwdqr5+YP
gSeN1fRTcfjH0D2NfgjascOQhRkxLQIWynNB+3F6AYokTiY1FN69AAR+LeCa71nZ
L1L3SdwyzvprAivyHFAXYBdyggQxCEXq51DEjz+WvggXBlsQBFiwTgUfNGXdn6Mx
rGhGeoBs5Foqm0nUNSVNUW5IBOEUZzyPcxoEDZbKbsmrRYEM/0lGy6NgkF9eTc0K
nKFv+LkYJ5mxDtk5FrDYC0qVukfhUZVPxKhIIIx72bR0m6FsL11/q8yJA8rydzzZ
DyAqhFMeBAKBEZ8Q8sWXrXzLXykyC18Z0O7IKqiZXf/MzKosb9e+BZdeZb/3sqZo
quvBjRC+jPXwDqx3z+Ucn4bF61I9QBec8typ/C9zzBu8XGbUxjr6VY7lKv+z6uuU
jeXzF9x/hpkvL2lBLz25EpaE4i3iZW2W6v8hc4IS3JhSWMTvjFWyYnnz74+KqMOI
AnaboIul8/frGojMK0jsfVAANmJ4DUpM76aIKz+OstR2tx8rXzt1vXE/GWDsBlRm
dOkET3hRC38Vx81Z0Z3nFFPl3dGw05RsDbxbyjxQMQMOunIr74RE7OZUeqjqOLLn
lR2UR2sy0h09lUVyq7410XByQKFtaQEfAHQDjg6I8LFtkBHBVz1YkNUzkNGIOFcP
i/8XA48VRkJERVeAJFOp/MxRwYBTlegQZycANFfnEHg06RDzU2Fz9ykPmM4n2AYQ
wWNja680h3FTKHIhetaf/0ZsgSxj8YNxDBxngbV18VLORcQY0Aa0E20n1dMQJ+uE
XQfm+tRD345GMtUKkNINDkqJRq1gZ73IrclzQgOZyc60d9B7ng86L8+2WfbiThSc
bpIvrQadcqw+hPVb2gf8ovUFgYiDOsM4gITISsa9L9ERg+CS2gDgLt8mmGr9mgFm
wAHZK7Wvl/7NwZmYyNP+FPFkeY+XTyjaAA/HfISCU3Ha2nTrLNvvOpLvGBVMi01V
t3iRRconPad8YT1lQQKIkdPiwWp5vRYwnNnuoA1vBd/02qJ8K+wx49LozasqPEsV
PDPVRvgmMzQ0BcorERRBuw0OsSTaMODqzN7mmTJyvk6XAIwP5ukmGsNZq/47jMw/
WD+U95ellEtyALPIjY6qZi/Yjd5C8Q6t4LQRVPBxKq970iBLpR0Dr1oHEGe9I80P
I3fPa2MUzoh7Nzhw3xJB6SlQAWW5S5zRZ/gk27s8xdUQrpBjIDuipV7jO/xFPN15
7gXWMzEmK865dTt8C9nGGCZwY+M37tAm1dXLELznsho+1cYH7nbBOz0ChFli1K/9
ld1dIYBvlAW3SO2kQwX8zo/8AWTKPckXx72dOWgIAIqP/Jjrs5x29ayfNo0CRffy
ygrm4ZlhLYfZiz6U7d9nYuXO2qIXLq7EGsL4eMdYUR+1oQwJlVao9Fv/WGsrx64B
B+uL/H9Xj4oi4FmUoJX42AfQeBixPqQmh11SlNJGZp/qgrP4rrN0o58I8y/8I/Iw
oKsJ4j4ZqRTGBapWE1OlkOYcab1nl+JV7BvHI0Wbkk+j2c6IVt4sPZ/BpLYc/7ct
ekI+luN4MI/Egh2uu/Tr10pJ5VihLIsIgNsn/0vZZ9oJW2yhFbdTY8ej4KKB6eI3
JYudr5Wb8n2H8fGZDOfrXF3EES6yTZ22xPl9jsVOT8uU6tQBHNHcpNEwfRDMvj94
ESmyG7Q1oB9jK9tHCvedQIAURKiTxxdEnCbbzg+D6LY8twReszVo/8l6JRSmAJQe
2S07XuxVbiMHJ25krEyVJ79p/4z6vZWgWL92jLS4eAP1DBa9hUP1cNNyZPnG22LO
2xbjgMM1c37E8zp7bdt8Bm8R23QQeI/1AkJb3ogss/wR6UeByjwMo6IiN4RXeS/T
KphPZzOVUjkXlkBMdCJ4p9yjuKvGnGx63x3GfcilDkKkbvtznZeyNSjD8br1Aws/
IbybBnRV5lr4VMOGhiWZB3FvIhqkNn700hA7Kwzowlmd9eHLoo2qPiGBjRVNoXWy
C/C/b1hFyyxFBmRWQS4CDs/6hOpKBN8IHm8ZG0c/5+QOMBqSeiGS4FLdjzHvKsHO
sfaoH1Y0UsLZitNXInp2ambMu4E0X4HvOBQyqYSSh3TxAJyVjx9NkRJJZ0Egkk3q
IuqYNPjgvik3CJcRNNIde6DiivS0tCNEtn3PwnJrRt5bL4yk0x52Q4pcWg229xQ1
DFbZklyuxEJDImLAoyWUh2ATkEonI5SZNyEHswxwqwwCxtqnqU5tn8v1glnAhfIK
Yiij1u25sJd180mNDINEJqBGFq3p3v/4IWfzAdX+apkk05sdsGgmtqJnLlgM3slY
nXeyZV9zD/uN6CdgjaVJvQnzFKq4BsKfGCaLzHlwjh5b/G/ByYEO/IPvOOxEIG3s
9v+c5GDuzVEnebat9vot4ZV6kQS9G1gauUepLhrgmi26zQvmhUeinm079WL/j4rw
IncZczLxFgDuAikUKgFMHAEt/0F6WaCRfcu1U3n1GmYqHC8E7St4P1fJMVgu4vm5
8+ioHfMd0yxsPQ8lMdVfJCzKdYBEvcmwif2VFTv3f1WJaOhEOR0BulbZ8NgorQE6
u+LoFMTosWJEpKNcwKPuT5BNQULtlpZdqBbv6LCoQW3c2GTdDOk23GFi4P0K+R7P
MwbJIoLJeRybOpWB8fDUEsVEcqB6se+dm820zVYGwBk=
`protect END_PROTECTED
