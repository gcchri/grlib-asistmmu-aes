`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uSeZoZXWAUDhjRkRs0vrWCR8PPVgX+Z1Ixn1Dpfmi3UwJKpg+uRZJ4TbwWUilcrO
cOLXFCuMJU5hV9SROhBBWtCiFz7pxJypso8RZcZu1bRsXmFD4QC1lKGh1Ierf3r0
w/PxRXcrxz3+o1Kla7S/pjG35lh0CAZ4iX+BZ2x7HAXCceWrX5/bTUpp0m3PmUZM
8zM6iq95epn7j5Lgl2eCsEIYYbRN0f759IJX24FuklQciVjpnK/Pu8o+uQX+Lg+5
Jl4yMEDB2fIOR3gG4L89hsu3+QPFP4QH6bcRIdMy/T6jfNcM+2mLh002qJN6+x86
`protect END_PROTECTED
