`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vHM48+Cvi1Fr/3/UnHCbq87hqPjrrj0aUtcsXGgrquo4DIIN/WRtkGAq2zQ3b7e2
VoqmX2RSy8yNBwFMgtNXAdFR8fffxdkWvd9rIjxUjH6acjdfj01WtCsZzwBO/W02
E6acF+3ErhO2A5eThTwbdXU2GcFTNt3xOnAkj/zD97I622zuoXrzbGuLD9QoYKuZ
D+lKeJJwVZH5s5frwcJQ2gzGDluXQukpQNMBsGGtPXJtl7jwXHIlBSv5N3pwDBaS
0xvdvhPS03yi/g8YK1p1JTvAvmNA6q/8CnztDmr0zxxMookZZ8ARboVdYIXN/1GB
r/IgdLNYbtFREFHDo8rWeu883g1E/Xf4Wo8LtV0eH6AIVt2jZal6Ac/pHaC5FcUb
qSLGvNvSkfm/ygsRlXbB6tRdmo2S/zENhDB4wVdLbg3MMcV3HytyskVQEu082WF1
Lumv6j4x2NM6MkL7y2yVd4ubCP1ivoiVI68UJcvVKmWAA+zuHiBs1cEhJEhq86uR
BFrGz8gSxuQZuhn7MDZdqQ==
`protect END_PROTECTED
