`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6tTveXlmImj5CwARAEnFuTCjzQXMdEpUY6c6j8bRLkvC7fnzSkQzjtMnUvf5qtkX
DVeU/2Sro4VeOaC+wD7GtCAxu4QylW5q6BGidbDDLMtGRvIAK4mt3gwB7qBYDvOo
T2lFmo4xfubl0LBwfXd71jM2y8G5VdP4slFYHqgog/waJEsL6mj1sfWeomXkfaJc
fV4zB8bDLWYTQ436wEk9GRUg0K08h1yu2ttgRBACtcRZc2eSQI0qEa0lMe2KtVYQ
Dpx4VnZg2IdQJ4BqUgL/bryUvuWSc5qwo4i74rzSlk+Q/5qOAGChOa3610BFPK1x
ip4IHZ5Yd6+kx1gfuTl7c0MvEIAMuzR+F2GOIRmxaEw8KkBaw3XCtyzK+fjyS54j
VAlQHVPCayOAfm++wrDuNFbQxZwRXLZpqxD47upQSkIRGckgeXhuwEPwXVwl/7Dw
Tj+fy4KTgYdjr91bBw8cIjIXfIuzhK6KE6SjvdtroqqBaCtwobV/X6HFvfGAphwt
uimoGVXoh+CTFg/N8OhjyamagsZOdM/Y1T3YfiqS7zuzq2NwZVDWN0IpBKpKieIC
Cvo3Gy8wqSKxBiV45FAQzZkISrtc11rrA1rl5zAb36jFvFjTSmyfJkBHt75SI1h0
PWjedzIZZfZ08xKPmbge71aAZYcZPQHDorLIUgbthNetLG88CcOuqJzcax6e6RD1
sQimeRWjKRmr8I5X93mwoAa5NZ3P5fLsaGjfaEGX7Y8aPAjtZ0YktoV0dwUxWU7F
KziO+pvMefEP8jaksXMp64fokY0xcD+7B3S6V5Fyb56v0SgJqRt3KDvuT8VDG13F
De+VO60dDr9Lvc+8YIJpOuxEAyUDL2zz5YN25PtGkJI3CCZnfOnlvFDe8R52D5D+
NLcnqvnN+R5zTWHKFXRhFRYcArOmJzvey1RXEPVInuvcRTxHqKQzu4G3eBNanfvQ
HNHrYGEFvdn/3WHWFFgvRCdtwH9M9Ha69RGjufhUidhfQ5nP/6G3OAMdnT1s4g1C
1EmXe0bR02oFbyRS+QAGuDgH5F5F7nu2VBce+Qcv++38olY9Khd/c8hujaifWTrP
l6KE4VW5H10D2PueBg3xQZgP8DOzt184wYY0pGwD6OrD3HCuy5qVEfrmArsUyPVB
3Q4dnUeSRr+K7YjMcornAmkF5wqaD95hfcisUHQVxvDMPTq+LyjwMrTGkbZYd54L
gvVN6pxluhOhHZlEkbYuhMZarduNcG7TwoG9oZDFrj9vI0Cu2liivh61vZ4H7d0L
oRqowd2R9W8RdJXoZgpZpU+GYynOmCF7ToIZUnMW1WjGLQy3akP6Otp2CXlnwtjr
KVkKFWaNPeUhFyzBK0RRULM2pw8Q9vQIu8hm0ojS+IER18+zhkVoAk/YKEb1rzVf
yexzOx63NOXmw0Hu0Y/H4bq0DkPkSlKhPdtEXB5dkhHRxGRPi2yPF+ncaK/tZjjU
TcupDj/IPPUs+p/kJBui0wJyo33fFqIQYO/9y7JDnIzvYT3dOqi5UU1kigQQY5wL
iHdc2b0oxJxmkQPiLNQ+ngtmU3rQK4rAq99a5gAzs9STm0WhaI1QBV5ixY9Hoe2F
0BMuITTezFpGunIrt64jRTtMsqqJo3Xdi2NINkjuZaerWzThFOd0ru22Xa63MZUo
tor66r0HIZzT9xbVgjUHY6fOnOmbH+jYp7q56vZzJko8fz1pBYER9AP1i25pZPUu
Fo+R9XxEcVyGfY/TBopdv7ApS2urYMwYdQEccuF+h19zivBZRUkohju2Zf7/7eqN
687DxjNM54fUewk9OLIFo5XzexCAI3XzMmzxuGXDaMDedzuOURAwbRg3VPK0Aaw7
1PL7vanIn4acEcu8kHHl1a7JeMsS2CKfzPo5fnuhEbQ7YVZbqKcwi1U3ZL8lSe1Q
he1o8NPoOIbHsfgNO/evOJ77IbC9dJZT3HTY4zUWRwwL38QLjqItO4YH11O/X5g4
2A7ARaX3ulW6zThjuLFzcpmqP4VuzlTu1DVfxURxlQGCR82hsNdlQ5LfJcTJ+eon
QNrdiatVJy3ex9o2xx7YDr9n2wZcnXlkLmx6Z1hnJ35osEUbVS+876EOffs94ti4
EgxW01bm9H/E5RrckCvZALsYzr+zTUoixwWFqUCmZAoKZGWCfOKSiUwrRyoUBMSl
3mS1S5BuYqG09bRXiC2lLGU7IwudlH0c+G0DdcjyWTFbkXsDOaBuhiYWrw1SbnyP
mJzAfzQ4xCjMr1gs6jrMwyiv6fv85xHCnNenfHbE2z3kcDakge6Ap8IZ5IJig9kO
mEYUAZmHhVE1x24uXa8xWeee13WuRMy/ibaHWeU5dsAY4gTUfRkZ5watiwkG5XjY
lShGqYor3UAmL68MD8hxpqqyYcuxCKi5Gah/kjgH+GrD+fVLPzOJjbhXrFQTTzIE
JotTnuymy7MNDGA5WtdjCMTNxd9pVwmK+/ThMHGy7fXVKcwexeqdYbgEmCLKOy9p
bnR/eRB94qCI6ZdmJihaWjdwSXlqjkAkwjXLCpz3MjUExusWpOgR32fDylhqWueX
/hxcHFRULltZQ12FFaKu4XbMAPe4ZV2+NCdKL6mUQ/PijigPw8xFFuS0TQM1zo9d
LDMJrOvSIFZtkxVojQ63pYrcX64qJtIBRxyJZ1ORGpNZttG9h/QLCV7EzxXwo6J2
ruNMVNuqHmg/bjNlhRQqcgdE0BCV12Sb+wXTcIxAe9Sg7eRqa+RQhUMNonbccgK+
UJArvgytecQnp7jVUxH+hpKKDt60qBWg5UG+Sl4AarcXG/kVKfoU/cVTafWrrGNR
9GPJU5WG5Wm4zWqxn/Ow8w7qs7QfBpN18ZZLUQEWixn5oyadbuz8AgJddshLG9R0
Vrv3IQ7MmS6O3ybQY9zK+RJUhIU6npJnqUBo7oXM52xkrPVXvTJyeQ+bQ/Rf1LNW
yILAP+f6fq0ekOy4Z5HQZz1Ul7vny1Ax1MOngsWN341lGZyzxfBJXk8hjRTQ8E14
B0P9oyKPOO1WTgE1v1JQ0m3XgeA5XqqUqufLmFo9tkh2t64zdIUWWFiR9N7Oa+kk
pEzuWGZRI26KehlsmL9BTMSRg++PnlCW4c407yvs7TWM02QxJdFhZTxJIIM9GCI7
JfTZg+TBwfD2kogT+v4TfRTZBFHifySVWx14c11hpye5ciXd1kNE6rAEeSvI0P41
BCLgZegNO0q2XHoMVBtkKG+QBEgcrmJilBmh56XBRE/R4XRkZj7LmwLu3GD4oMuD
umQfpW9KqvEqUJwdjOMHY6xyCBzSlnZ/bViIh8qAaxn1Bp7jm/rk1wHoeUcEEhwN
Jv8QlOqMhvw+0D629P2NSndABQm4527YBYK/Jus3T1Kzo84pc/g1pcEXcZZwE+AU
u/sH1eHN+Lbvve3lo+2QSDUI7HGyniD+UrmDND6NufQ7G0LxUPNR49Vx7ULBhhvn
N282NeccMnpSGa0FmA9t1xk+xm8tQBRYOexwObNKqEYmaGplZG/h7x/OhYnYaV+K
JIkTacBZVnSRsX/W/l04H6V4F3w4GwhQRh9VQC8lyQsiJqdV69VKq/mT9y5c1IPN
OTpq0BTrEeimeIfEdPDDarMuhxdXWiwxLSChsGjZ4fdq5Y8fBDs0gw6EM+5R7LaQ
pJLh2lOeR84OCzSnV03ISxBNZkwh2BoXeIsRJG5NMKO5hZlbvtjmnMNLHRqlc1el
5EjWTTlw6Bsd025nst3gyT5E9ZiwcH4j8faaUjCwW45F3xRwpoXt7VNz0cdBQtre
pTSoE98xxzjGrYTSBrX2zz3Z+N3RQBHkNyMNwyxgT+QKZ9MohbT32dVKZw1M14g8
n4K7ZfEJXt/elfmWX9pssuB7Ct7isZ5NcqjNgztLvP4s+MjoqWKkZrhWYBuLy9+c
VbRrNkfYIfY/IzDrXphh2Q82LrekKzv32gTIEaC6+7bhrk0I2C7XkCYbMwusc+0v
3/WuaCMQ2dhrITf3sOOgGT+h3nRSCKko9urwtClrZ4ZbYAzum+1guq5vdRev0MxI
NaWaVz89ZWhNQoKmEB4X8+92LOhC3/j19D6Q91HjmgQNaqyJbhX2PQovOhjozvM5
Swcnu7BDjoXAYrznpiII+QwtMpcOsJ/sb2tNjRZ7H/Skgtxv34XaA7eDK14yziik
yjqXEj1VI244jHwwhI4REqk0OU/J0V8fFb6qOFAWFQXS5Adr0TYBwaEEV7JE7xpt
qDTh7Y8wOIuqaTCISXQmgBEA8eAZQkCfRdtn3Mqz/KI2mq5BhOB6Hsbk60tBWNgW
CM32PsORrmWnKA+dlRokWya1EwBlITlthDSDVBOzcX4/GON9gd9t/g0bHZJu0ILM
aejG8Tpve/dXSJgJrRrBmBLo66/xf2M2Or3t4JGslvMkKx/h00hrLOsGy16pv14Y
tRSepyhIzCGgnH2Wj0zGo0ipPlcUEWSVSLPnVqNsz69cZlF3pHsyuVqrZ6a8rtst
JPAwetR+LbhMyFNrDE/Od5E6FTQ4rjGZE3Tt5t9OuHO2ccVYc3dAF2jMULzDlT2H
wWyZrQlMudzBr6/sFQpcerN+WYi+MFaagTwc28xTdAiN7ccetFE6Xe3B5Lopp+8D
hT+XgcNKPTRRsGCIP5vK+siW05lATC9TDGYYPsSmkzRPiOVDrhl9xlZF7i0FD15z
sONm5yqcqmzHpRqexGnRHky0lTjOoWbUB+FqESCeIAGyqW7E+1IQ5vMfl4yjyin5
tszka6NDO1BgZjNhPSRE1m/qkflMzYDqkAPSSSFN+xfoz5On45G1lSN/swvU/xHB
KF69wTAxc4oA/0DxkWmHF1BSDoRcirRBf2JCa94uD1zzi5sevcWvufyp1xgGmvLE
g+NQDI4CqbZH6TPm2am+VHqlUerNUsJUMypPlnI5ky1nflUicm+OTeVMfDURSArD
I/oq2UOON16h+DnMPNAOL3jrZzFh8Mith6GWmbkpslFt0B5R4Fds1pqOTYAzGPi5
pqgBIhrI6RjXSxn05x3aeqz5IYhI0f93ptD9xRz237+M/n6f6wjiYXombpWJxHao
IYUpX2o6hCuLylME9/AAStIlmz/LVnFXBvjWH1Kc3xinghrrQnjmkeXCb+eb1+p1
xcfJxZRf8L2U7oitUubKGz+XtcHMgR3hlPjJ33MwJ1UO6nT2AbSzLHZJ2J0ym16I
fKgxeSX9VFYFvDRMa6+AHkmifE/KUiy9EZEedX6nlWJkmyIjQ0KCfgQwhbdY38n5
aP7cug+H2e/ZhnYA4v8w8SITkT58bFgT/tcZkqkHdQYjvZPQuYH7O4lEJymUt3Qv
gT79aZ21eqCIsq738ViJ1im931R2hVqdBbcuYvolGNlQhnNdl2z5tNQQssEr7/f8
64a+DRkJzj7zLPIC+aykQj5de+LFkxnRkNB05rsZ1CGrz2EYEs9IsEMC0D9xoJIq
CtvSb1oqKgKEOPUT4bgIYZhj1cvM+aSTJJ7ZqJQXCU7YsnQITXyjBH2bOydlZ5Cc
rjZiAYLdIuVCKdwaonnVAS5Puc7iMwC+EZy7eBg6OVo=
`protect END_PROTECTED
