`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aHQv7zqLlPzP/XVysEiHqYtWs6yk/VJ16i5OvSw3ka20JX0k2Nix76tj7OvvYSCh
IcGqSZnxrwya0vyMM4bhc5Sh1SWGInA8nWZ+jPV369RXb0tkiA/v99z6suC8MOWF
hDe8stceNvujUABYfegGn/RsJRlsdn4jsM3RpVMhtIaxAGbJD9J8QNqjMO45F74D
mgn2DkiDZLCreZ6OMwX4pszyEvVUVqeHAKPhaBZfd0XsAVPfSHTr5AKJO7U7/ySd
BnSraPPT332XEPaObA1db+5Qr8NG8UWqS78nTW1ZQL3t80nqwxV4LrF2I9dXvspw
pXbCmZBSf8nCq1LWfqvML0gKyIByGVlI0PWR5hz+hDwQec5/dwsE534dv5bLmdGq
7569Ff+TDrYBh2CTHzDBnsqgnk+x1uGNAOT//3DNoQN0wPylmkWprJPlMffM7wfk
bWjHLvW9MxK7ptd+eDK03muMMZ4RTbfwdJd7/ahwGPzUGldeznZYYA1AaG/s7yzh
ep5Y+/nmYCChZDCJRaJNC7s5ojpvAqhYoroz8BGiK2eXl03rBSjEufAXmWq8JarM
+DZpmKdKMuWPnUGc+3kxrqc5KYv1f/v3BhAXLV3YnbgwLTsdgNO0TuABDGwQN8t0
45YiHbQT0NJamaekusQGHVHjNg03cCI6INBrvRGLIB+RuMSJYy3c4B5LPtRtJ+yN
qGbihSZgQCwWGa8lpO0hRt7B2z/yC5eeRRENbdA3tSCV0+VmbWD1uVmFw1UKS6UV
NK2Tn5kgiNs8IBqIeoxGVStR6SpCVYllCe0yhoT/p76o+XhORUttwHwSuA5VUgfX
uEjysNffOSvaT5920Zji/3LZ8Kq8j7AyNDalpdIc1TdwuMD5DFLpS/fEDi3bhTpb
KSd8wowvnY23V1obHtTeVmYAdH6+ATjLinyWMFLxwrEyNSHmBWQH4o2dlv9eUr4K
BYBfSjaxVJHNm6hgJlPKVrmzQgqp6MYZeNSy4B+b9SFYFZjAvY7buT9zEaBiG+Vv
3jYP6JwK9nT7bCdipJwcvGloEtO7xeqBEgBTu9IkzT890ElZTUTERPgPUP2LA0O0
rDpHjG+ufVEwATyu6QeKdg==
`protect END_PROTECTED
