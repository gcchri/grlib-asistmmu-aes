`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NqxaNSWmLs+s324ve8wMI22r/rwFgDl+v5hqj4stSRFpeoU0USNolp/dYEpkJn+W
rsiABo8vrul0PSDlwgtxy5xduGxZG62QvEKOaNtusykBoSKVevaY8YvcjX9zRH1F
y6BBcaGGgCiVW4wHPxmVvhZ4pLyclnXT9uQzJiVGjSTMMdeJETkJaQZHo+qfVNQu
P6y8OFVQmOyNpEuHqTc2VgxIZCbHCKEc5vPCK9D/Vqbh+haxzMbNQd6EvoB6WbAa
MB9CWxqkMdhnm/uPoqL7ltlnZ1n68yhGfyWcENMvq1A+hvYGoFr+u6/fiyWFpYHA
`protect END_PROTECTED
