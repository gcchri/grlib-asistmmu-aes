`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OyF+cj0MNiVra+X2ADvrwaf7mM81FKxD0xsI+i0o4QSKVp8B4uE1rUBgVX2NqWel
086LD/3Lh4ytX6hnEem8W161iDupcrkjY5zsZf9eJNrauCwpj3iyoF4jnN9TlUGe
ffIRx67LSPvYaP1gaI0gTP5SiYAVBj8YstWNw7aidObtmtRjJ/ZhC5aqdLCnbLIT
ksp6BSlwBwoB5yarBmw9l6w+E8BKZSgfGdmifBXg0Yo+LuK+jg0kB5oFCtWWebtc
DTurVoxAUF5BexOLFspVdEsx4GTSVJ8d3cWY/LPr6P77/SxXoj6Xls6Zc0DTXu68
BkG2j8mFUiR7FVjiekSQZCJNjYsSncNEreOQVoAwGHOtTjXkbX3gImGny6E42ffY
OAAO22LviiwunAPLIOwQ5oyuDBGcidihxCk3WXzsvTg=
`protect END_PROTECTED
