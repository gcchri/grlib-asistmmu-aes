`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3SeCMqVSpR4dYdZBBiDlxVhTQPPQvvfoy066G1+a12hjvJXJupWgyq6UqMimEuRm
YgGPIynhCFkDIH5nf0LUpjNW3jzGOQG/RkFX269SgqTXcVTO8gLkBu8Zpo5CeTBL
zEYXnTYME7so+F6CuWqn/27GPyd88RkZ3uT9YNlM9fr7GmkhqBSW5c35xX9WQnxq
ZyWPfJkr3IIN3KBqtynI0zWMbFCF3mb3U5YAZ9Xvq9sUV4thNS1ERsjWq+btCqkU
JD6V4ITLAPnaFzpH8/M1oiuPStcT7x62U5KNeAyGsquSnf/yYYkbGLOd5YCYT0uf
QmuHOXULGZrzK2y5RKhIHWtHzcb1fCKurr28iWDNuWgc5UpHLkFcu49dn6AgfeQ8
uhF6etTQtJDuQ/HRYOVgkEknPkL+UegJEK5QPnOb1UM/puwrdkFwFQNxiIfQJczv
CxbT9ik8G4DDNk4FHMYd2eVXdekEW6ImbGfHXh6tkN7nOWVMZrtxnx4h2eYmdG16
/a94sbpN9Ye+UVYV6gVtAvnNFwnQJpEPL0M1wu/isEJvAIMMBMMmly1vR5cf7cuT
2SMYHX9inG+UUrPMcQweGonpYEGyk2WW34FWd26dV2ydV5HuMnWzjVdAgThaF80M
nxrg0Hgv5lH0d1KUqRSYluLS6q19S1/zwXPWcckuZtkphormELb9kCPsoNu17HF0
xMlXfqkqEvOBJ7plWmAFIQFzxgUAcRHTBQ/RqT2KzquoM94Pff7O+itmiC4w9xXs
X9UErZnSCD1qgS57tBwzTIu4tnOKJCDVrMQaLFrxK1w6urSYqRX7ilvqIOX54uUo
WmbrBlw53Hzmznwu09DUl3RnxFsLxEbs+yfXvqO97bG/GdDn1ayYFw+tyP+vMG+s
f0gt35c+oeldzgB23/LqNjZAeH0SH9Uyn28nbAar3DXEuaL2GG+9tazKRfQ9d1VH
w/6qS3gvabgIhz8bhehMeXSUaFsUeWwGgqFU+nW3uV+6ikkLVjngw6CNXh6LIyAR
hwpAGbPRWo5rjSwZ94phU9JRarYYBwbEmJAJILMnKyfyVKwDSRkPpD8f2Nrx1Q7E
7ExZIJhYzEoM97rhNc0tH7Dtg/6yXysdR8RUD3qkNmbpAPEM4Cz+JNXcWrllfYrM
apM9WyGPGg+f2hvVstWFKitsU5CNZ08ur3guNNHmxzlI4VdLMM2TLs2rwjGfdiu4
W2v+kct9k42wSaFfn2Sw6hTZnR1PNEeMl6PXJbhwlOo361IyqwZ9mjfzod9Zz3cK
aphwYTh07eoMdx1AfZqCFJ6ehDQ4659QUN1S8aMbH0t//6cIQtdj7Mds2RTJjob4
9dcjCdJtJ5dWrOR1dOX4P+5kVPxB+HAZH1oKJyqmqzhS5A5uCLdSuQm0Q9UD6etX
lnQVY6mjP0X2Ulypyn0OUjfg2nnoR5RDLPFA0/pcc7l7deU878F52wVLkvrLnOr6
DDNEs9sesmHRwvyodTnsA4KfbqGdgglBNTD61aUkBTW/FULoissAtk35dqFMkHn+
6aVjhtag4NQjrAFMQYiwHzOEqhrja4VXDRW0Mb6oB5uKIf8mwWBE0H6tJOYriMBQ
0iAU9U8pNUzpzVoS0obt3lHK2D8VhNp76vf5knn8lVDRAwJufx9uGN3XKAy7up4/
3bIYFI+2H8wlJkD7aTn/PkgV9kesw7GonaZaQXHVpEiD/vp0gcXeO7d3m+P4J05K
H/cy8lJvW7EHDxtGU9a0/rz8c4xNyotxv0fk7spHUcoKopoiOGofGxRwokbWh4nT
7aIECaoJQg6O7j7kcSMHXUgl/36xylzE+/YgSZYHdSbftWEjPY1Sx8GI4hptmQEA
1NiZjAZIuFJ6OPmGdk7z4wIcOViglQzGoOhp/+9CG32yxgP8QmgEOIkJmtNv3kVw
gVCiNzOGXPLNGVhw45dbq1oWRxkxI9ygNvVdZ5BfXhPi/8t5red7aSqn6L975Y76
bccx0GiNYHreckssBqzXREUD4mxvXWrqT+Dr6401qi2gU3hWQGYytU4rScH+MpXU
j5k8xuTWdkhoH91zsQneKz4ov6/Lsy9WZsvvV97pt6VWDkUWunLbN1ljxZOdmcXg
GibKYIWghbo3CIly5v00ifq4sXXxeZjbezkkqrzzcuBPWG/9ZOi36HTFIAxYW5q3
HW2aQkAKBH5JeNJYGzCs2ArOaD4+4SAisluJXCzHLBPaexwDZTqhPsq1F20YQ7gd
b+TPd+Po16HyI+2UHhNYVkx85ZxRyT9l4a4l6yZce4Vt27PhI4RcTdwiGtFfUZ6J
dK6lQjpzYgsZqjmb4SAtyJnqskmB0eF8npLuvQA7FYwp4HT7gAdPVRqJrK7M5hq+
31Ie5YPPAEUSXZAKEOeWWEouU8aZrLzVFM5MCiou+7X3OnmDeola95b3QEMMrw0q
uoncwkLKHJplRbZtXmuA7h3narjT1Ff26fU0OLrHjL0MPpJ8deQPZir5pABbPMe7
HMVKVK6O+E10VVv3RdsJ7qNoyL1Z4LBqY3Vh+W10j0S/Au2ju9JGO9biCwRprzOY
i9fGfWhIa2BFpIDGpQ6ARMy+ZEdKtHTYyHwpUS6uE6F6VNPhK7N3ZvUBifBUhGqa
fJvwERZRkUrDrVtK09SpZHJ30Ck7RxgF3RO8IT+2R9Y9FtyoOWwy91UQK7ZRZPO3
Q9tV7sCMJ4asdYk9skQQ33kF44eibSSG+TT1Ss7f12asQXLiuZ7U4FS6NDZ4mpeu
Ek68TaODVPonexwi91aUAlWqLgPJrriq1Y+uP221rGfYTk/pSXIjAiAiL/VabXmB
+2GT0z3PCcPyZlzCBpnVhkK5N8srXUsPRYLc38il/FfmzERpDgowTrcPV2sBPYX9
SRNkOqmpduAGEbWnDQe3MEEFMhviexIOcIyqNs7gNa5VKSZYa79NRPKoWAm13ka2
fVB2LMHgelGxFFxIpo9diLlNaPzJ/1xtSqJU1luH7Mw5EfwDdsnRRB1Eg9gMJEcn
PUe/iJFgImdN+OHZPwuoHOhNjNOE4bjhcf8YzxnvNi30nXY06YaNL0BlQwLHRYk/
qj8WSt1ezaX82nc1fPW7V4+EzxczQEqCSlf/1BrY5tOAW2+Qc2JkjAmor6w16cWq
w/LGOQjYhIKs/1l2nDHMbDzaboLLPK+VS1hHjY7/60mlt/JHENHt+vpMiUG4VYoQ
48nKBrNM2e6PTZckMH1fxOQW3i1gkOly/Ii21I0K6byD/qcdNOLDY3Cqeyx8+c6O
9gRLVIj1B0FUxwmrevrbDU85aNZnp5B7tfaDCxDNQ2FKZgl09NgG35ghI24o6FpP
BUmi1IVBdpSTecvXUIhkSjhkUR1xPhgK8/YqrObIlsGXhSt+sUW+nT9RpPj5FTZP
lP3tMFOXraX5aEdd6IZqkGZYSQklyQi8aZuJRsfhr5di6YhscHFXVv2he2IXVCAp
BbNS4+aJjEGh0LGb1/VQ3ejCbjoXg6CNeCRW4kqmGo81U2N5D9Wg29pSQS5+eq7O
FshwT5iBT0aDUeK2ObT5ztF05FWL7+zlt8FH3xz2zIZiKhbxxnE8eTXEnlTiTwdL
m2bfYIoOU17HNhPpp1xiNBsFFO00ep2rkes8igFHxF/SvpHD12vsMrL8Lp24Fh7T
DvZ0U1rlrW2fa0r0BvYZCvTgcPSdIAgZ5uBnoPDFiZ7xeq1fZNcxmxACavnTtwwB
9nqjWvMR0rEL5QOqBLwzpanKbuHmoXTyGsGgaMESiYWBU70RqCzD+Wgf1CIL9NgF
bg8GsMKe6TGNwvtjjp8GFV3wz1xSEfuYHCde3euGWP8WUCdDLLk+ugB89V25ucY2
MnwCcCyf/F1Nm1O0/Hr9WIlSJOFh3MbPCARSTkoHDGKyQ0WpXIwey72cl5IfWE08
6HspJCvUOUv7IC3dBJuCSKzcB4856W0zayeWtkpZK785cZmEECqAEeMCmcyXn+HK
Q63+PkrEpaAcWn+0uJ6gQZ1FztYN6BGwcy054+hypuw+2MW9zkzihpYN+0z9kggS
CmnBMXO5kZ5JGrJpTS/O3ErQdH7pqjp0Qn1Uj+WiPWSblJoDZY/QR/Xe9JYnDy04
OArsXB/MKH6mVDtLv30xKSawUeimefBjxPZhNucHADSVa7ROop7Bs0HjZZB51jip
/RYeHHNrmG5ZjAbJa5axoFP3QxCD8o8XZ3mAbpMYMOFdRbWhKZgWNmA9GQ4dnRk1
rgSVlo/r25HBWw5D8n/yNq3sKp+cJwJzvHZTz30rfsaBFDwFpbTyN2Hh1qmOqoaH
qyAyjRQhY3cMf0Fu9fzpSUZwVw+BOmjCVlvR9uxGKDPB9L2Wwvf1pSOyE/HsaL/P
sAPuxQv2ewREhifIIHFJEcrUPmhJN43ejPgfcHrwFhGrnqbvlwnqKpL4B4J2d4It
1Mb3hbtia8mV/n9S85WNRQ/1lgMKyCufz5/mP1OoI9GCC+XjcHjH5YUm0It4IPex
hSrJp07Hu737IJvfdWMfN6pr/siX7G0vtUhEwbSjbfzx7Bn+itwVWZnPcQ/B/1IU
PoMmjzZWEnXsECc2dgWZV8TjvqYGpyIbwWEN7c7UyjQGgh3QCEomLMFU/qP5gimo
v041v/Jv8vZe4treS6ZKIBhPa+nBkQcxblVbwMoHeSn6OpgXS7gfuOCgDHAlKwF0
AxhWpyZlwHnT6SbKf+H5hfWYC7fI1f5gSvxOD8WNg0Cz6j/9fgwPmDsFRlBFajon
TSCMFebvhBD2k8YV+EaGpjvguYadOd3l0JdVp1v+2Ew5ITZxz3+vh50ZcyQWnplB
rOylMYWBJifogna8chZ5xF/xkjAhQHYaNOKqsz3CbDxyKOCPLHLIMAJOxlhyxQVo
eR1l689EeDENJSThPIOcQEGBI11/xYZXtoC+MRs05RTVIVPEQWROtOtNgT4RFujR
etDu5vo+xymfHxVGfZ4g89zb6m53QLjOjGFSJX4NuPDjCVm8o33/IhS4+YQC3pBp
t6mFahEjWkGiZBlcW0mvXHiIt7guWf7jL1JPkF+3xYf9AUFa7OaAoq/9e8yNv9Sw
VzzntaZZeaN9CELhkzUdtdzvHxJn0+MQC1AJ9LJs30QD6jao1j/5TWeKQPT5b3QM
U08i7yKwb1aaTqnAjLIrQyb9waLsXLqgMIvOGJf6h/V7MWqDg+Q/BkmI50trHANr
UvM+flhCl4kKskq1CLiTxyFe6xJQxGoNmvFB/naNlB7ydCwfSp0ARNcHRg7VD9OK
iJGHqfGUIWX38kyAAenPJ7nVt0VN1CfGcQ7r5pSdGNN+SW9sjoACFqiAjGdDPqMF
Ed4Wm4toJZvme1X1JLU8q6gS09SGAxwth2aVnC/trW0PDGFcvxshbZbGIS6nwomn
9AjhLgNpm/sZzL9dX509+BolBUJRhme1xhFHtP8+uxiD4NYcoTNXy82Txr41JXEo
oowfpB4V8dGLs3wkdcQqu8hsWRqri2VDoEutWYxVoNF2tAVs1tEqmJXIJZZTWhqJ
zj30yQvZNk2MIIAiABaj0wCvgw1UC5TQfzV9dU2o6otKDCJYrx/XnOMPMZInaUal
sET7A99Ze6aISK4Fg/9LJ3gw1W0GldZjtO6A3lvkngYT0def4nAI7WUtcisgCLET
7uo0gC0FhaTDUKQ7hq1Yfer6YOi3VPrQiI6B2O9he64O0PDpi++wTenXg5RugyJq
JAlVr7iWBYPsU9XPr8H784UI6xN1drS7ykt0XZWv0UeRg2lDRTlHpRBZq6tmGS5m
lAU60+xGjJ8Y/M/GmozEwrhfIkMpvNa8VIFb8Ccc4eoe08APKTPgMj2iD2RZtm+j
nsaaDQS8irtqNKA5xJmklg3f9eLFmibS3mXYXCA0SM21xu/DecXrHOYte6VHKjWI
WeGav/HjbO79n2RC31b68HbCiGH7/RsJXfxzB3eE3BWPH4U2RxfHOuHu9Ig/eeEc
UJABi82+GfYrKZ1HAoQ1CLUDB4iEOU18CMdLFxtkAjrFySHl8RiWjpnWNLk5QxIm
5aQ8AsS1H5hMBY169ctQXQi56dwqKjZKMH3iIBPDZyAV8if6rH0x0fV5xpFpcjhN
dLTOZusSaxC36+qgYkjIsoYghO8WsKF3GQZ1N46OmxTCpeniBQz/si75mn/PdFsI
ilIGF3ntcoZnjSqGvQHMZE8MCXYr/S9A5czPt4fsKRnKsDxtf+QIRSNu9IKeALb+
SWlH2i0ZOZ+ndHM2nNhWpMdO1NG9BNqnfNjfJPFJ8jKLii1Vku7iYMLReUewg1wW
cyABiExXiMaSq2J4wqfZCU7KkcXt6kEOJtQqEASAGQ17pUwiHwQFgPbo9ve5u4Ld
c3wH9aI1J6k2stcFiGqYLx7V3GTVZh4sy3cc+N9mKEp5e657cmD2iTQcUOfCFhh0
yYH4e3z6GAYwn0p7EcfY8ztU+Wr6M2desit63rAxftr9VV5KN4dPST6y9ubtBf2f
3FDpNEejJ9QmBojXUitRjC6QpAmlhJoD6bfbvHn2/ui1CYzKTAujCdRePowvBRP1
xKtGf8u/Q2LOjH8rb2nTMpviftmD2BI64cQr5wzQUxWPnQXkBwJXXM2Mu8en61VH
Caw1h6U4Ix+M/DBtPAniwbQtUEq7gBKx6sti3xFRTHAnIci1dvlGNJ8n00uj7v8H
9ntI42YpAkQNAZmk6akUvdzRJwLvbS0ZqQT8lXEVA6pjCNRR+Ftkle23YnJMw4KC
TbsszsT7+gz4ruahitO8c2uynPkehAjABary2880tJc0Sxk3xjLGIhHuVHrkF5nH
QBl2lHCKI4glPC2K2xTVomr2DnJ8OKxVyQKBTtwhxqnn8eO4wcdyl/ETPzSYlFU0
bAk6hadw5kj2qKNfPEjGcNMSBJQa8303vRFs+PWvk8sGW5RMvKTKBpEG/rIbWxgJ
hfvMUfE6B7PkcU6iPJnVGWm2koAB1Y0ptntIaL82TnPKA12Q9sdvbwz1clNmYUga
E75cA+uCPLNKkz1LAaEQuC6g7mC9cRdxJK2T03WyGLNMfErb0yLj1o0Pa+RqjYkD
/9br+jXTn9vq/j8Q8t/Jjzz72ee6VG9sP/WqjyIPWlnIamdcd1VqdEBe5rtr6S0F
noCyAhtO+PPHuC7AZRYJpCqaboSTjURQsUsAhTIkujXxi4zuo15PFiHkYENudlOn
uIkNuFfDQ3P1NnsnDCH+rBPU4QYhWk8kK0uWTfQ4COxP5p/cSS/2K/nyk04ltuNz
l4cgQcu9j2XsLTPeDI5XprzIIEknlKTVM5nboE7kgq2C5HaFWNaZrvsW4N8UwVmd
wQqt9iRir9MVlY7fyTf+vSEGcQQ3wDo0WA9YMPN7CR43YYYLQ6ZGcCUIHX0ihsq8
zYZbaYswcxjCr2jB4fOJXt/qJo0KbWAaHOcROk0xpQKNo0xk1LhHV7mIXuW63xny
CISGkZIhSCoFQvfsbM+8SopTf8byu7XiFEsnuk2Nek6GJaWNIdNF2cdWBUk4ranP
V/mPP9TUWBW6BunbwGRLgPTW6Bs4aezjZ+FNing8p9l7AAErR5r2oFc2pM/tftl/
9lMHtvgTSyrtx+YAtVHxWgGv3Z0zITCZ1g5EOG+RD6GrMCqvkFQhdTwdBw1vRR/R
tWZg75DGPTtQpmxi0hRkIWuK4G9hzNUD3B+8+PVH1wHi0isaFVom9XrCwbIfS5US
i++0uGWpl28yqR0M5mwEE0/LZcDch1NKvFGTSIRS0tukcq1+BQS8nIPikOO2wQ8E
Kpokejl6l50Dm5yXA166pR3PFsoXrakta0d91vHl8KRUC9xJt+pz/BsGJI0lIT5m
dBgDnqOQI+PtDxyswGBfJQnBpvoL1s2xY0S11D/xdMK8VZ8LpU8fwmV6SntErlIn
4A7GksWGtlJy3VYeuMdkgNAC1bLxb3dFVPdZnyawHHLI3rIVJlkq2ODIRCggoIPQ
n5iT+d7qAErlxqOF1i+7FJSi2u8cb2jmDt5D616pkTkD2Akyi5cWezXPJQIatrsl
Lqj9/Ngou2+/WXqnbY4SX8iRj+ckqzJstEBeHI32KV3z5MqWv80ZV6VhF8xNmzAW
XC8E2p6xTOuROIN7Q2kqQ5RlnW/QSINUCCe2PtT60yFtdCmYSJBbf+R4/M0oDlER
c2zdhkvkq/y49vYXmnIn62GnX/I+lGAkMu220P2V2XPhBGgxY9OlMeDYi+qTvZlh
dSIeKYe7dhvNY8VVh02cFUJ8IkM3KOiR86O2NDz0MxVTJ6PRAz6rcyzoeBQPrOj4
V5e26/Cpi0gX2YbdgDlO5bPjReoN70xaPO9W2RPF9cnUNUYprigbXDne2XV51gWG
jprQG9WnpwIvIM0w8faiiQ7S0yuZka0tB8aLqGS0InoHgGYmLLuJqoH8L9uXNPN9
JCJ5qKXXlZuBEUq/Cs0ZcZYPweGJXYcHMCE0On5gbcOP0tm9ZSkylRbbJ4vZlY3i
FMwMLMkz7wFfGcQIhrs5JU0T7sHnT63PiB8yXFOo4nKWaJUxLAVdpF2Tv9beR6pA
wEF9HN89v4gzXVVjas5t/wWPYpzmgnhAVOUPRJ2pE1RVAGvkZirij4kOJ8FFrZsL
4lZoogwGL5+mkvuznNuqG4rVzvgRlWpst6u/fzcEYEWgLWwuloKtIrOJHliLyBly
1NUAd6ytsUaRJSO6J0AKMMcA8jfkNHffjdWj9X/NS2kz7wbgW31f6nQ2fgNnQOg9
bi7CcQ47SynWF6Fzf8QNnp+4USUYjy+EVFgQIFMdHakR9rItRkvtAYxQEymAMBaa
1jqWNe2UOZhFSqvlSfY/o1BWtjWVF5MPJbcSz5DuaaCYc2BTVIsKsIY7uB/DJhHZ
zSmGiFhmMrsax8tZiDccDNuadiEi+h/DWemHl2fhWFGJeI+tVYcbpeiu0pWDE+nO
OuDfp3dJCFylFihIZLtfxs+MZ5eExX6ja5lOIgs0IK8VVG0XmfpOIqrwiaJzcscw
93oz7WL2l0ysXFAapjHDmthLU7oJqyJatNj42iF8EM9ntu2najCWuF7P2ejeGArf
9fWn1317C1N2nSK+/qBgb+wrHNrfeNC5DLkPB/oPc7nd0fHhxXlxTZBIEAgEv49/
B/LjNkP8M9l8lSmqGvPa6GcgNlxJyVCGAnqW0jFxULfNfTJBFuhvgJn5k3KM53oh
lUhWUgNDf6QLa4CMg69jBtg8PK0e7C2MBW5e9rE0R5ke8GQ/SnsKXSXhOINI7BXY
la+bU7jZ9VFtvM/IvjN74hhyiJEfQNpxisxsOA31Cd6ri4pYiFx9t4SHAcgDklfh
PoTUpV94E1d+YWeF9o+9agSUqV0+vJyk3/L4kty97KHAE3nxgRE67Gf6JltmUhTp
CtY1Hb9blOVXP5oboN1RlzQDYVQ3L9PelC+9oxvxj+jXwbLylQtlZldtIhityfZn
CDoPfp3btTu/JAZ5utpkCkjgFZF7HkXwk9H+7TiCDHou+CY84umj9Xf2+rd/e4Hn
f/5hNHU0z0Tnsn9iOdgvqM4x90ib1LlWgURdNzo7bleErYpg9DVqCz9i71qTFSNH
3VjbswCGuLNeTnKi5Q+UuT4xph7f6ATUboSgiXtkK6k0h7B2NF5sWI5P59DhBa7V
AevcYwwdx1/YP+j9xb5BgTuw1gs/ijPZvvr5OVmJPtXFCGnAUriSGiE1n2wvHfoX
tpaoBYBOHHUe6LbsuM+ajyE7Gh3iKrKIo9ONcbSZnZ4AXKdjRHbYhxv9tdwmA7iG
N5c696UNgoUzdgZeQ+GrVEmXCiOvPrwTCMSRYyxYp4sBblLDoP7idtIlJlaNyvd2
P84pkRtL+u0M51TQmMl/AEG5BNkQvrR69hCMvDPgLtMAOk6eILGms9U/cANID7gx
wYmzkEPRC5xi1RJmjfGvpgdjEOpGamTxVrgBTnLMssKe1tvX8sH9wudoowY0Cs6v
tn+YWxACGWWHhTOlE4fxFEbqB6oDbNI4G8fhHObtgxOk9PfCemku0N20LPEgH2wY
RMRquY5xA+KXZJgwWK6kTU6MVO58/H1r7JbVHzMgAjDq2/YQlAL3oqk9m7fi+yXZ
bIGzwU+4eQWp+UMjNM9hXm6BOBYH1jRLUCGbiQvhRnA7Hi5WT5Vc6oUtXhjr6Rvm
nyVIRiPEKofeAAiS1bSUqBBswep8A9sl+XeKph/OFuakYEDzNHeg8TDuwMNdSho9
2M9ilpoukhMa4c4h3IpDN4ZeG4EQfCO9NoMcrxayLtngajMGMKn7ImY50MZTe2LM
sKBA/vNuMoNkV/uZa8bk1LLythlOOp8mwgyw7cR0tkuOElwX59Hq2gSIYmTQsazp
Xp0NKs/PsySwB5bjbbPCtGz6sYJI+01qZDWSqQQGUKfL06C5aoC176of5cCoUMFO
d9fXHYqK7ckHfog5OVXJARAoVx5sH/5psWoAiPLCOHsx4jOlyOlJYnQ0tUXAyDYf
NmRCvL/dQ42s4dAuVVzl0ahhsI61pS5tDa3D+6EH9iFGjZZqzht2YSyjQj2O67Ac
80aQ/Nb7dVDi081Qwi/wTFkn8r+VBgXnrdfSEg6ziIhU8RbOtwHsZb4b461fX+1+
0/tdwKzkQ0J+ErL2wENoGU2kptrU7eXm385ingeFkBk5JsS2DuBe8nbZdbrevmHx
RC4h2dvdi4sEZn8+OwzVNMoNR+Hj8bdWiYLX7QC0uZEb2v1UGwQTryFJPC4Jtn/k
1aKUm92Cx3fl/uVy2tZY/EopnGo2NZp0A/oz7E2ALKMSahSRMOMRgrRtzqSqkGBr
VsnbYGayrFA2fGl6qH/iaHKA4LxiDDNp6oFrq3szIzE=
`protect END_PROTECTED
