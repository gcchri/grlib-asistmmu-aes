`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mvqeDqt046F/Pd3Txb4H10f0503Kr4lv9hOrZzbutPquw39ytAVAeg1g23BqIjAA
8dwmEfaPi54JVTgLwi3G/LPtv1AK4N8p8S0iM1h2IAfbmBleYl8oTvnDxSS6ogEP
qP3BXviz0fbx6CJyi/hA4TyrIxlr/sqw6V288PDWMcruLz8XTKfyKsHkxadQr3C4
w5g/HhwE1eDSI9CDqSDp2NMknl9yG9nLf+uCRy8/PcpmHDBeroTwt16KB03/fAnI
AHrewJ2FzqTcnfqOiO502sZY39QqIskqwd1xF8ju0jUrqQ7niVNjQxW778Q8D/Yh
4Dw/UR8pLFRWxm02lG2Ui32L7UkVx7Kgpj2Sc6aQ+cvtMdybKqGTjv66ufs+WwPB
7IikUmlbSWl03UJZyhzqS188cJpNqOYorhfK82GYkeehJW66PnpvJVdOU3X7XRGI
i/E2mOwlu5rJmae97RtKTYMsAPz+jkFhZwPlbq8z254BpqD40TAAfwqDVJff8Ad9
e5JffkT0octM0Sxc8PnzWrutxUhVG5sMPYc1p3wMsvowUNWe9Eo2s4p22rDtvjQM
gzY80VQf2grZrs8dAQfqUWIIL2j0YW62+NoNV1CXbL8=
`protect END_PROTECTED
