`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gXH+us6Nv/KTEJQ+j8Qqq5o8Ysj8gOCgC2Velk/mGr/HjnCzGA6HFg9wMmU/rL18
urNd3pBpTFaik7NFQyhZ3VT0QGObE2dP/xQlZqgTZLoe4w/AZEYG6C//3m3rjUpG
02PT3GBqFCMNogp/aCBJQDRFuJOjDN5i7ao5PCuv2Tv27ka4rM+sZmTA3cy+OpjV
IV86rJIeZqFLc6mxuDxJw+ukzMYABOInO8mt4RHV014NWAwONKXdWkVoqCFSXsSP
EanJTsLG0zFSoAam9yliHXU/hKaChiP/5zo0fatbPhNPpg98/x6I3+XS5tNWEFeo
IMHux9saugmDNDmwzgjr1i2dnz9wvxafW25y6wLR5EUE9x4RbHTrgw5UifSsilH7
0gzZc/E/3R9yHC++vXP9HAw+EfswiQze/z7CMKrrAYMyxDRkMl2VZEAGf/gv1Kck
`protect END_PROTECTED
