`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
txrNSl3Ywq+YmWUl/UDn0E7akjn3UsM1B49otKR9sTQgT0FVvN/DpRG5sQFqFaK7
HJ6jz7zJ3InSdrSWC87+XdJBU5npF5OMKWugsmwUB7DjR0VZOpOcTdhE2GWZ3H04
/zCCETJU9lbOtYlv+aQ7xW/u336vpwtlonUBxqGe3WDZyeNvTr8PTNXsQ70bkgYu
FdDzd8RUzw/GvlV4R4y9eAnOp7sptxU1Z3JsPLZ/r1hhcokXAAsbOweisN+jFoMu
PS6+kWsQNl3jQC7JnHw8sVe4Qk51JaYNMi4ILHhxEDwudeq3IckCNY1YA+n7ysGd
EAASfx5qtRVBGXtlhb7QA0R/aDTqLf1Er3LRT/6zzsvdPGEoSjHd/8ohHgzlYY+N
yQdTQ9vqemxFtwHOr3ffThqOx3iCAPLXzYup7qAeSUhssJCZ8tD/KSmS7GDaV/qy
UcLVglNdOTh3yNI5cORSZ+bDOvJJr3HPsXST9+bRn+kZ9r+szrVMmoOxeGZuapb9
NiPIT5/GbBGB68A2Xqv8IZd7/+RVkbF+kHJWrQjWogP7elXK2OoWbdKCoVdEuz/0
95iMqV63u6PJob11qS5IhTubZAv+21aN6cJPlAF93Q2STXInMbIzIGlQccAqW2uS
ItBE1zdHCHcZM6Ap9fxYmWS4sHz58otfBOAHTrM669qUio4+1rSmIJS4WstIG8yG
k1yCxmHKRFwr0SjzrCjOk/PgN3ttYw5MDudBZtm5++I1+jONXjaQVnHkst8Qikc6
T2UFGraaeYdw6s6jWdAVJ2zQoJFyVjZAhOj1D/86Zp60vZz86PxT3UUxPQSBGTou
oxS/yNzPLcAO/31OtjZSdoTT0VVkd0I/QiqvqDcgIDekL/34hAfAvIBXDgW9WCvK
JUrRT2Z93XZ3u6jUTpzAOtF6JVDU+K6YC02JVmDiPnrHd5LExR9zMOQppykNC9nG
CDGvKs0uphfAjOWJ0dNQ4w==
`protect END_PROTECTED
