`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0FlpBa4CeccEpWPmtjni9JsG7r2/olLQVUWDZ7DvTFXEpXoLVB8Ei5OW99zcZ12y
pPbFpR0LiOH4tBSsR7jYFelMomk7VhzQz5o1vWPjw5Z7KYvlEwohydwHvILvIYCZ
tlI0+mBplJ9Z8OBab/hndrZkXsTxAO1zs8U9sOi7V3sHabZrfY3j3k6VX6t438Ty
L3XloBxfeORNe/evNM0LnzVi40Dh/NpRqkgtaMe3ZceQoyUB/PI5BAGNwY8lPbAL
gtQIkvtN79fle5B6WEoX5TA9yZHIc85tX9oz/d5ICFhrsK7/XqkY+2Vd8WQJwCKu
IrnfYH25/elFg6QSmP2e8u+0HfjCCztp+SKgNB0jItIIomUB3lO9rsYfdz2xjDO2
cdYFA2wvSSkD+L+qggU1UktDu8lzSAqhgo9Lx49dRTU=
`protect END_PROTECTED
