`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XO7a7m8spYOP1ByZeOHfWKcjGFeUIpPnQs6tAWSzVXzdTQdeOErgfN3GBjiFlSfk
y8yEpBZQSosX+XE/RrgRiNn9T85KY9wQefP1GkUnu6DMRYMwTSGtL+YQiAdnyn/2
7+muuHxye8YzwfQ0s5xLKzRHYp2QXh9msOKIf3+eeuQQkMUtl+E4GjX7mQESvrxM
U2NE9wOaZzgZVmZZ6ULdQzMgNSZislRL33bR7qoN90xWFYgCOtrnY5qTSbc3BbwL
Fa1tYCfjbxEwx4JUyQU1wnIINcoSewuZutUDgprRCUW7FghSdDn3hIy1Y4/3ccDN
K5II2sTsEajVGzO7otZONT48ffxlHmysu3xckxBdbXEm/skyHBNWumCzAkgc0pFM
3MdKV4oR3VS9zgY5aCegY+0ZfcU4mDhSWOuPcgXUuJLZX6fd+3VOF2qazIwtQmaH
5BaR2BuWWnx46I165akRSeIl03MHsGsVS++DDbM/yUtYp4EA9bLih46Ye/e5g+Kv
qhWfvbe50Ha0Tix80uAmVu1J79ZCuXOuv4giZJSAFaOS4sFrlbEBLlc7brJEDRNL
`protect END_PROTECTED
