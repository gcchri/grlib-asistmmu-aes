`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mpG9YTmijkZuHQVQ4vjqkYevUPn3LmA1JoVhHXM0UkHSnIaTkNtekv/vtgw5NHxN
UV3GqztING9y3qQJAfBz1+Cll7PxC12rp5YJsTzQ2arqFR/Vn+bu2hptcZ50y8L8
KlnJCJpOt8dGjrFUi++6IWiOKImdjx7xy6NFlvqhBrT1ECsqUJizuKrqLSSoL99J
zgQh65dlfKIvUi++otVA4BX+4G13XkqYXQ0VW0z7ZWXmRMK26P9AlSk+0eGevI+l
ljq9MnFRXZo2QsBsHIuIduhz1X3G8N7Ay288Wb4jKLQ3Okpl7ZQOEZlDj8gbZdZ9
ZPS5XNezFDufzmrJc+p1mqO8JktmX+QijKFQVRhjQS6S495kQbwQ+8YZW7RJULqq
bHMC0vTwtbWx3akxcih7fTGrEKGG6Ehfr9WcZkY8Oeghj3EDthQ1NXKfHD5tPiKa
HsVptbQLTdZwQL2EALwM90TkksoAart3RsrFFCTzjCEMaDvCX7WxwK0uigmGlyMs
VKAGaSCUy1ESODr1sNOLpXhk52u7X4FCl5ScRfnygQI0p3avBBPCNAqSOtPbkYDm
P59EB5vZPmAxHHkken+tZav/mhQW3jYshEA7bX4KM68IL9L30OQpn5UtYmyQQgO5
fnxfwHJARkTN7EtuxCtJVJMwqClaWxG4S9KYzmdai9JlE2hriPstWhsnb2wQ/p3z
iZS5ncmaQIHwXahgQyLN7LC8OYfDZo63sFPBSjPnUavl4q/AAWYlz/e43HckN1pR
NPReTddI14ndiscpTzoD0YRYPNbBsWG/KVAhBWuX1RhTqeG7CpfYjmdvAA56q1p+
MIoa1OAmY5xiEDvTUmrRkGrPieYfvG+iHgJsFyon1QNtO4ha66h0F3ehhZmtOq9g
PaVws8lGpdgti7uKjmi9BbSMUQ5DLavTgndG4u6bXNHDTYubu4rTbxtBIScVTXXc
2jtcJfMfdFsNhJqw7mvrISCxkNNJa8UDr1tcXT3J0WQqtJ5F7E6aeEsrFJuEutER
KJX/gJxHMRwAS7/X7zomWa/sLbIfjlWHbybY70pnxTVzNQCgF1OYIOrq59fgNP91
d2QsoQDXJpGcj4TVveHlekQSDwxapRP7F12mxMGkz2eriqyYysQsQedGE+KZ5TIa
lJUDc4ujf1G3wdOEriVtJlOtkLGphJ17lcW01Prz8U422rBCnn4eCB0JnSAjzcRx
MOkZ+WoBrOXi4jnG6fwXUKq5XPbtd+QNPApMWoSPFQxVpuOO2ObXoERbCIO9o8F4
wWOWlb3FgsUYwAgNZWVZHWusIYqrI6YxqQekuOP4msBQKhr2uVQMzvG40h9L13J0
Z6RWnat+evPQq5PyrNYyNkdTIGm6RtvwqJaerDtecaJA62IJn60Z4GPcDX7VOJ/T
h6FG7HKT/THnykDBExuHu0Ipktjxcj4HcBjuWKTQnUqottXwnbSD8qIVb4j/dWkO
MBHUrZOGKb9K0LSy1wzE6jU5uEMEUcHA82fEjmxW6NxlMh+ysnKsAOJjgRJB8PJW
Y5LOndabnavVsdknI/eJ/026Jufb0j872iJ1CEF8hWBjAGCgT6BVCOCOoi/OhFZ5
+2KV5lV49ncne1tdKFNX6vVvCAZ53kVb60l+uSl529rhefWPeDFjcZDLV2DYp57n
z13e7AjnzIQ6GTLAi7xuWW9s5R8xTM4zehsAwJy8YSyxKNTUYTpKoGJxJUDUrkbU
1hwAqqxYf4uLjBJUnV/Vv7OLtGVHgbQVC3aNaKmW+eA9y43Pkm0XD6cqEuld/G9I
1d1auNwpqXxWc6JMiP2BndMGmTWKG6bO1ctWKVN2SteCqwyPMM8cl1ZHqFto9pXq
AXCismZuL7Bdrbfeotwm8dzmJbpf71/A65y6YZ2oA71i7ExCwi2NO3QWfd4f8Iwh
KTAAg6YhWx+6Vu0yDKBifIemzsHMRZpQ+pTDyOOTdRGXKnVPdgYyXwzZaltB+CXO
90GDGOO5dx77zLdPSwZND+MMX3fKK5+MRBmPIjg2aNa49mdlxRoGrzzsASdg+kjw
gQQ9Htr8kUGUhcawdiqvtKnLLJPZl2GEOL9cNw2FWNhEgu9djYqXaQAmZ2UUFxpI
9N8aISCDaqJslspTXdA7epvayqgwQc/lQe6Kq1gizrHi0hp7G8jJSTrgeIyFDQ59
ytkYBXaHypomgFP1aVezoUl88sN7IXKCRwU4Ds1Fyc+PlJDcsc4zpvkSYgkLBFw5
/Si2zNC3a+Nps1LZYIbcbfMQ3qwTSTK5WmV23agm9mfmdDH3Fj7QFf3VdeWIKoaH
vWiT3EgI+QC2BMyW6D3ItYX9onnLFUE2nt5MORkK9cm9bg86jdcVNEJdTvAais7g
omUnhcgOyh0a0bfkGmb9r1Par0WCMZAfTiePiKfY8MFMwY/iPLd3Ez8r7TFvekJd
uHBPlRFBhYpL1OzV6012xh9LOyvFYg9QCs16fIOIztoV5SVptC+RJpaVNbzGfJ6s
eJD8FIbH7KyybtmYRfH9Jzt1SRwI+yUc1JX2O99uzsYEAK/2uL5wEuza2XUssxA9
v0wPqFRnuAp+w4XCV3XqlWpDFLEFp3qY47BvLvnzIvaWHo7XQ6g7aaoJB3a99aZF
r06Uj81lWws4OU52tYkpurkxAzpqEef26X8+NJj8I7x6hF/s4lmyLZLzNSTuhlkJ
7URzLLqYT4mVpd0STSiVrC0qFvEZpKNnAh0HCnWgBCz9Y7BIoQGTtpqv5rXJE2//
6UZio/istOKgrB+bQZyD+5FF2AtOVklU9w959+SZmiiy4lBfyIyzBsmreMnx0FaD
/j5wBMBtG52yQ+pZZ/IDvHZ2zDmzGbwFmx0yu9rl9GQl7r5D8r/P9G0rh14kFzGt
h8XYRpvkcji3nFPwpvpQugA1MH+VP7QIFsviBgG9zK8z5hasSi4dsQp5emZXc9pA
VVJ5OQ6it4NNpeSLKu1foc+n9GOHOJ8MltnClsgLXeuVqxUkNjOIFsZtFsqJw2mk
e3iiZAeNQaHLkPmaNVlP4PmF13jGuDCqKrRllcDkB17k8jdnAm8Ia+rRPvdIYu95
9GyPBZx42+f7DuyHJjSG6z0Ua1P2Q0quZ1YitXM9QR/BoYjyoN+wOFCiL3ghcKMa
QTYK/3w9MGIkP4Si3Z+kwEjOptM9+EftctDoWluJOv2L5pPKiGA3f0DrAozJ927W
O5aBo8OVpg7opaSZTrLy9HERO7ybY8gXs57c7xLjufffKVHyzCBQxwbBcDchWQph
KAvH8DRAlG8X/Wf8p1vaYnRWjdhroXL0EGCc8f5kDYVGwLXfuQ0xdq9rJhkbvpZl
yGmiu1G4FgcQ+XVXgvezq8mymgGVfZCBv95QdPIi0LyIGyW5yobX+sGAWYQBSwuy
Ze5nKqGWj+aa/DNluPzJ+fD/qphKYRl0diLDplc2VlFiSqK+c4LZllzv2AcsiE2e
b4GFsx2j3SA98hiOrzlmp0oMSKBw1/iyMsjiPGtv+q/79f/8+wwyzaGDg5yHOL0w
NiXVdHMzC0/EwtXx618nLGkMygf/hSeGKXbRGdksQIpeHYO6vPXsnIO1gePQ4kEk
Ge5sC3a9Vu3eCJUi25BTEiy8nyb6x2LuSEwn9UEAJL2GbgsRvIVpJ3MKSZs6dx3P
mKRMxB/gpX9UVcI4pihCHtCCmY5Mx18eUsudozi0sJzRv24PUyA/hEfRcuAvIRdo
glbCQz23Z9+eTfYGszlKuZNnREEZtCXk/7Z1dc5Sc8Lb68hkwu8RZhFJyEN0dlem
2Q4QBR+Zz5wLa6w7ChYsyd2hrWGaYAqSQi9ou7yV8EAHMr2R0ltp3ZZL5EYtgVRp
K9NHsg6gm7D569zuM3SBY8uD93zNTLyAbi0OE0EimlXq65j0fAY++IRdzoNh1TV1
Moh9QgnDOoU7uSqROLshV+PfpPJe5f7iuFWFyRBWAJBb5jovXTt7n6OqaeLrtl+0
yco4CofCtNEMcKe3z0dtcBzw7+Y2q9ZyyiKW2GP47WQd2NCcaX2BvbWcOQslNUCF
/huhbQ2jxI1kBB0RVvzMvHOSf35OQdvKUco9tBU+WsEbpNHt7AMzTwgnNkTdDdnz
iWCu3tAdWHaas5aGJy9T2kqvqsi6/9WOgJEaqdQyT2wrrit/+jOSCAQtFeUjKhjn
SpUbNhK7xt4PKN52p1nY66gRUThnTgEYlUC/doXlbJ/vOt08I+2AQlwb0zMYQm3L
oHc4vrWqd/LLS6jlLj5W4Y+37OWiZLRMVdBEgWl+L33i3qfLwPtlWfwfyjIVMzhP
EC+f4LfNHJBNzfHd03ycNP1HBDbBewHeta9ZiS/gMmhkr8MHKV0FocZbRrGurVMD
DWURiwJsAwmcB6Deewpe6UrtnjfEkCYuZGluz8oMhVdCCFaB2NbFGmdQSJk0YqQG
o23fBOgAJisZm3hE7ODM/dwhspdAPpv388EvYi4xotC0LTo1EkPRME2H9O/UUMlZ
lVtYtNvDKyGdMeFUifW5jl0+uSi2JQYA55JV8TVK26cauMy2mmyJcWqR9lx/jeCk
EGm+U9waTKWaUUKdLGQf+fzHGOSSPUBY80sJJK0705EiHWEWVrAUw+Nk0LfZjzT9
Gvt00jMXmq/bR/PKRAiJgkLIZ3qpdK6CfL+hqVgpxWp/wJV1/1mMe4zkMeH1qz+U
gJg4A89SGJYa6NthjVuUNsnbsOIfh09qwI7/g7rD0b5o6zpTLttHwZmfT4N07DTO
RfM7CkBwEJrqQ0fmGo9r1ocp9ijUevcm2N5+H2TwD7tw73LESyPJ6Ne7l2h36cIz
KqT1ob+bp5Y3sZKostEm6JczFW9f+g6STqLE2qDMpkuR09vmZ6eUKtnF5ZpaLULj
WeG+XX6PYgJNzQWR2cS8zCoBzt75INsIOH9CJ9Z+jmhDO0EUffESXJqYW0KJ/5Zy
rusDJAnyhQBv5D5ez7wm4Kuf8JOPmtAa5GpFIBSSfOJ7vNgopz5XxwRRJ8DBTOa6
jpt4knBzHblHYDoeA7CfNU3g+p09p5ajaqhqZfO0JDl7mku62e3Wpzbr95af9wwj
WTKWBPuCcbAiuqHxULi0Gbukiv0XxD6wBpMtOUTaqlnk8KLPK3172uClVOxKn+RB
rv/zTqHzTem5r4a0En2PSTOgmvOVuhxOIfHP2oI6Hf1VIG7Zmg3t7fchqGewoghe
oEJyj4pBeWxydr6iAFTtRO5xMSZcicw9h+X3r1qEOKQJ0QyezGQ0MICBtdA7dCUo
iFEhQ7h65nrQy2CtOUm+hKvauYUsEfl/Nr/B+VvnT+WGXFPCxvZh8njlrowpuG8V
yFNo3yJBrfnrzlFFjXMWMdY3zZY+e8YV0hZnSPDQI1hFXQuu3iJK1YK2jP6wfzj6
dUv0Odl2akqce7kNGOwWBsq+QVeKCzUDw9ddhmkV9GKXf4uxs0LmtAiuvU3h2gyt
GCopVQHoXeql77Xm+0l68BAc7YL3C4sCrumwoviQegQzAI/J/jhZFCbnH7EOBPkj
lJ8VbI1IXkf2L7xangEuM2XYzhDksqiYwn7FF2GddNQZh7jECZc0GraM2+4/nCNA
LckHgn/lbHwBpzr+/3yYkrTp8P/Iv5WJyqBTHbyPuIJAx0oOZsXA2Z3EZxDiCLis
O9nZH73gMvBXPs0qV57aUTD6kRemW0VhLbqP7NqdkD83LNd4VY3x8Yckq1MGBwQz
x4CL3Qj0khj8upIeIVb4pLTiEBnsK9ih7qz+V71cu9Jw+6jt9Q4KwCxmxFU1NnrC
4PZwu3W+Q1myjKiCGnK/YrZcNvOv8kPqOPu3qSqGBs04d6Wvr+jtJAINL2u8rkw2
E/gL/o14q4ckoJErv5GhmRfgfOB10PVBxtlQEMb/TCTVU93eDsGbu0NFiEXuLsaP
h4f3m1AIC5nAUf8rF16MT7VEbXmUyqi9K0KR2NLLEf5n6B1KdTFn/JexP7S0ZY53
2Bpp5SjrYTvUNlT1SuACZAsvilni7tIYsX+Z8gDLD1Buz5+gMZg1Qbr5BG2/RD9Z
VmLTVrW6AyejSO0Mt9Bm4+YJQuBC37uvlWX5JURBp8REsub9/EOoZkrGqlyzWl7r
P7zaf/msDSXv30G7z6ruwAnvsGgbbu0XjCqMdaEXX+68HHj1WRck5Vzh819/Ds8n
wqABHZcdih7+orA4Z/YwhDEHqXbAlImYvOUgnxKH88zIPv6vX2Txvj0sKwPyhEHn
WqWfD74yyY3z/jM2GQ6ZU5YHA8PhouTupnFx0udBFIJ+wIck2nKnUaf05SwfModG
J5V2B/J++gKu0qsPLhqiiwn/OW9hoCm9lu+N0rCNUrHezYXsVCn1qmfoxAFV/qzJ
jvgYqdOIvImuKWJilF71ZW/LFE+ScTnL5Ww0Temc3oacuDiR+LBxCDtuAnQ4unRC
jMFvTfmyTOoJhkiCwxhJ3/aSOQopgq3wKQLmlGfa+KAjlzKdTEEwheZBzPZchUhE
D8cCPZnkOyUE8HqiEVp3QLGb43AoTYn0ZLi6h1bPhdY3XijTL4FzfL4YnTKUkxpP
tdgoZaomyQ+70UqnPq7TnusYan7Qum2mg6/MvtbBKX+6PZw5IlXEVrbi/P5XvP58
b8KMVp/bZjpwMkDhLgvOh1PA9YwzSyDpSTmty15kJ1MqHsOq2S25SHXaRld9h402
9y/P5LUf8/jDmIvtISEqrRL6vu/D/GFsiw1aKnyteCmsbggD7i33n4+hUVB7fdL9
3eScp+eZx0rJX1sq6/L4uhNYFPIMasbg+ozsb3Cn00AGkysVlNCEKjorpc4kK2pn
j2TfNgktNZzVc816rhvQwA98aISbozSdu59aH8iezHJRyVvjGgkoa3HxycWNTFiW
cxgjbO32HG9ROKGkxAzc6odWwGwndZKLvNV61t1hDC0F7FSN/WMe0wfRETEaAY6h
PPnpV+txMHDbvEigOPwSAm064EOswcTr3eFp5HXfcHJlD4plZMr7ONYoIIfcmHMO
N9ZAt4YsjG5FyfCrxO7X9VACXuzJbR64qjgBzHHRS8iaZ/50sWL6sKt8maKjxbcR
0U1bsZnOdKM6JcTUCF0ZXnQ5pSAJ/cPEKFwQI/HXilkjoaDALLMgP46h14kJ722o
kCgSXtBbQAssqOVbocQWsh/bKIlDfg0M+yPqhBxGt44X0QxIpH1Z+ZtAbQqdHgo2
IGyNnjdNdrl9wad7ZhSihuodBl3f2jiWz+O3c+pQboRwVf75ZD5toQrJ108ltJu7
8O2E11kbxeHVN4bXVHw1Wske1PAs/RQuDSCZ0xXQ7IngwjDDIas5wXDASNJxB0NC
bvQ9gu/Lhw7jMhh0Vx2qFltS5N5uB0yH5mf3Hz6GVc7nzvwr1Dqomp9Df7L0QxnO
OQHSJs6Vht7zqHYvGiZAWu7OfOl77VblmRLI9fuqwIMg+J+Pk3YzTBvIpR7awRMK
90HIwKL6ZtpV5N7gVqvw4NEU/Sx8ZOzGm5dqoMX5+ZzwABcxABLliBECm18VbErB
2lJNAhEGpEydhMHkt5goTYNyahgOMKI6hINSG0TvkTmwY9HSL3B9lzn8YhRp55Dk
AGcGW6PYeWts1ZTLNbXBk+lPbIBS8JsBlectqEzVv7c7L80EvApTG3KZQkIJIu7P
8s6R77rwnjjifrN03XXrqNNKakzf+oe3KuARNguMt9M1H3frKLoh8Ewnu+2/M18D
1ia4s16RixPmdy/VRPm2pfarjpXQPPlTQULOgg7gO4WBRFKJnU4/jeiVvlg9wxZL
5uWfANhAvmZgfCrbKfvBLxdMrCohiS+gjN20tvRwwaWfkHVhdfN2KqMQgm8YWabJ
pcgojB2+g2R1u0Z0A3hg/yd4lFLR1H15bVRM85qi7RmMm6QxYU4OZy+77S7QGU3Y
8wgYs86bIxE2leU+Go/z9NTLLawKbWUI6RI+kGibZoFS1PNKB3AEXTIPkH7sJitz
0y+SyTs87PYlToKrPGhaBK6oJqFSkvdkpZH4jKYZuOQ+GJznOK5Vx65DoTs+lYze
30fOviXjsYyHBlyjsf+0lClUQ5Xl8gn++pO7KW+83Bg3e8zMBAvRo1BQfVwxKGM8
abhyvagN920kwvJXaNhU+orV9cFXxmr4h9ipahPHQrAg3NIyiCI7NvYxROe3/ItL
0+WTPXVQXA6s97LrTSGsvJS7lj9f2TBLUBO8OxRiREXjrg8oXcY/XD5Q6owILrDu
OMF43A5PLq4szCx0F+Q9vWBoD6/Zmg9bAX3n2dmQsZT0RPaek+gC3VwcGm693+td
KHh+kdq5jweWXlyER4iYrvdzKAQmUW3RBhcUM0AvZhjjsJi7nbN9Pi6hvrMlekbd
IFxyFNY3w6xAh25K8QOdRjA3wpnpDX2ivKMG623JPEgRYXc1of21RyaY/Oi56Mla
3rebjNEVV4EJ2R21GWDhvoejnv69IRiRQI1jj81cIhtlj+/p4GH3LjEYV7OKcUoJ
nG7rpz+s1Px8bGYF+RHCajJ0A5LbXT2T6Af3xe0WbiFEhWNVbFuuySpphRyiFzav
/SoNMqAJl9uMpkP0TvjY5E8nKTvIfTGNPVyQm5asMJxxIzOsVi59mFchPKNrhePw
+rs4Nta1EzEYJjzyegyHacjJVsbBqfVXNMihyJhPYPuBDkM+Xtr8rKqbPcpZlBaP
8PXXdqOsNv9KLiU7C8A9ZRUGoUMEJbslUQDj2HPDupnedO+c0973vYZREvAg+Cyh
sZ/4geefM8r8erfTD9YfvJCln04rBxS8BHKzF6yBB4psu+jJUaWThixny3UndMTe
mGPuiOYLYU8uHLCkQ5PJr70W/BAFoaxh49d2viijsfrWHKxzIRbMpwsO4jZ2cYia
sT99wQzVEFmbL9mOtzO040kpRKzKQIbXfCv8r3fhS2WBNpd0xIx1leJThSelf/6V
S/y+cYV6yrRCzRGTwmTfOLJrUsO+GyeB49wMr12zVWTS4U2M1OjagYZH8tMTBXJ3
7cDs/rThQ8JYQTqEneQ2YBJjI6zZzyxVDOFfyX7HJoXf3tym4syvZMEMAjXjrHEz
iTZXQbcPgJU4HzhP0WUponfzgW2LDH1TNzI3H9rItJr0XAwFl/NTyPb5i8PVKTJP
BZD962d2/knkjKm54BMHxn1ZrdrlTw35La8BsxZ0MW0XdbZAz5wv3C7N8ZgtcBwd
06L5fB5r8epH58Ig52g/UKV9d10sCNzQTR5pW17/5AGS2/pcOJur8sLRMZFpF7Ax
nQ2nmSFRjouN5+XT0PDpPLyoRpm3Mr8T44Kl3Csk+lz5TGhiFv1cwh/5n8yrGGA3
eP2TR0IvcB49LuIsohoG6sAH7LVxmm9GBkyBQqQntOhbdXxeWn6tt9hSsDggTlZl
CIWlA1uKIzFUdFXBj7eIj4KBA4MsTST9yxI/oqXcphB1bN15wlbGtkv9M8QxafvB
hCVGLWDO1bTc9SQj0pjsqiyPZrKNNojA6Ytkm0CYjM27X5mfdGdW//KI0tALuUVF
mQSBh1OJyGKf7yrcf8ysKebK/SSBjaR2BIqqizfMx7UvQwivGoXwVeNwQvVn6QmZ
OEj2tUbypnmgZTK5nMiftF+V0tdIH1E/kzu5EXSlyqG2y/enNTvRLs/Tc+oWYTY8
lA1cqanF/enhCqQck4jXQcrTWwaFetIsg6b61octRcfqeYF3ibwpC7ArcnoN/897
q+X8/g9ou0CWzDep09geNwRSZbDY94PiIoKiDf/9FSeEqbvJKxAYzter+24yc+7a
AfVNEZnhQMxoi1FsG/PWmFZwJnviAyRrCWvRFJhxiOqI8UyRLrrXUpICP5yNAhAc
kpiItGMB+ka21dA+fLF/ggtUbb73NcPYOWs+VnOF4uygkAa5EtXLjVYWOZ7Yh9Ou
WsfqialTHoTHw++pNny5ikGfkGCnHpi24Qs/72wSYPaqUYymgh+Z8eUnbgdLLCRg
UV/9rsvtKUW9fpcJKaEKfKWwojfVyIOor4FuHAQhywoY/MYx/ANN/LKBqSbihJqg
JHFSzGkrALbeE0GiIeX7upAq5ih/LPoU59Js273WdGY5QRilMpDcnQxVGJ+5hg+2
OeA7tdHWxPUQEwIqCdeZXZJetJcSjmIpMC0gSvukkPayyZHliMRnfJgZRDr9dR1p
yZbEJdOCHCst1lPeYFmin5M6YIMa73i0tF/JjH3sC/eYV6C0DPjT0MkINUC0vp/R
62bz6/WaJiZJg3Sp8bNcCca24czKom8mKJUhxM/gh6ABPy+sGTSnuok7YEpw8shI
tlxmYnyZLg9XTmwCi5Q7wG/LbpTS2PdD1qZATDkUG+Me4tOs+I8LaIpOUhNAtaoY
T2MLb1wrS7Fms4QXQ8b5O0iJIlhb9fTLHdxSbXenir65iYSImS+4TK9CUKN/NE+3
GU/VaxqCY1R7R5fzWicDq/+ouDtKDQ6Sa/MxsqBxrydkduo0Esj4e1DFZccIG8qj
yPKkgyGO7zcJJWFPnLXq48jsikmfBiRLGPX+E5UB0/qAyoeGnfNY3NBOAxGDYlx5
XXJ5WCJyLaMbGsglFBQ26YWE6/RH8Tiu88ECXSykbUgFk/0+2gG9LVGe4oKRX8x+
fVb3201CpzvREpjAbq80Mluso6RJG9Yu99Qt5lWa44YKbbzDybYQ0ALkERcBdKnz
rImC/k5oZ5OFX7fTx2mBluPnOryFTYs3Nu3zhW36tlMZmcTHxn77mwJyS8ugiXyz
nsJRFuUmDnxNUDs5DA2FD2HS7ioP7bL1qgbMZVwu4l5UmWMTku6hnEsByu94IJDw
bDMgiXx4//gilYgumL+U3Y4xRvmRNhYjrsWUjC4GHuQHwuJuW4hABCMp7+2vNS5x
ReOa8ocXFX7DnGvCHC5zquZm+BtAk+rcUTLrtcY7y99LvF5q1u/VbNdWcsIekrzc
mN/mSu3IWSPZI8OtVJV/1M5LIyP/AjYjNEswiRRdw4afr/Rg5vYCQPVE5ZCBJcvA
Ld0RFCIOoa7Ps0LezP6xCf1ZcG3ylr14wleTotreysF+iwfHSAELc6JD04usufq8
KlYaH5tx1zW4MTrvkqfUY+b+LOsCXo4YD/Yt/miQtdeYdoADgzHlB9kFjWGFsW40
JB6B3vehE4WMMjbUWvi3O8IXAoZ1EeizvQcwdplCdDx8TJzBQOu4V/EYrPkuMVsX
cBh4mJy5zQK1eMdbh0uQFae/lqBiFpphU+3NqkEeE+sdjh4j5IJ1cjM01qXgNfBe
YQ6XicjnkXRM73vBkW/5OucwbK1VJEGvKNAnwFiLM0I10aqX+B8lo5eN1Ib6wFIh
wJnpKjreb3uRtAIR0emgEQcbF52v1Gi+nkHEuWgcbovI/F3WfOym+eT08hc3U159
5OZZRfKoc99wuKMRry1ChdqrSQs61cRhKliGtqJDZ3s5PD5SFkMByjSNzviJuJRY
GWCMei4iYgG5iPQljSFfKVMuBVRuDimK90AvaXOxcUMVa/fbj68cIJCQiOdw5xWK
B7mUdx5J6xXyoOYjTqa64hBBhtRRayqRvYXzkSr5UtedwyMvb58hrEVqR+NTehvT
tWlnsQhc/F7woHgchmPrF0JgGWNm0zPa31+/34AXeROjIdTEDWAJd1BSY9cJNwN0
LufAspeqrtpPTzBOKNZ5VlOoJNWK0DCEtjV3ZNyMqmzBwK24vPTu1/1dM0hccMAW
ZWbCH9DlaLPsA/7AfF+poXN/YJ/jtws3cv2UShoYe5RRzj/I6wVM+rnD9ex4Ucso
t5AIJ/rqr9FRlMEzE6Tyc4eZXOUQaopLZgBW89K/Ul41en3iUI/pZqU3kcIty2Tc
XOnn8nsmrVIzI76NJ5PfpG6eDPz+1Oj0/qltbsjfGxWqeQaQUD1Lihglyw9/xGjy
wxF4LeLJE78PRCX8EQl84E81sZi2p4xBc7iM1npjRaxUgQjWx7BECH3baQd/V5DD
0TXNMJWE2jprbF7rb8QTiJJIigeKF+Dw+0X0P2FTv5bSfFb7Lc+jmRHawtTRwrxn
6yDJe+Bh8NIf6FID+FSv75RdJLAklRCNXIzCD+74/LbbFEKpoNT/P1wOE0abUNyT
o/Y6nhNkwHkTYw3IIKnvIZhZRTQJ8kLj07s1LzZpcKmwiO1xb/9UuxGegYDnBfJh
pVWS3c6LnsIQA7MnSAyDis0WzgnjCjWsU1VEk5Su1lExSfTpb7bdk+hfKpLikk2w
Z/iK8Ht+aXTrU5iKYgB4TPpaSOjoy+292U/H3enHQHG1IZ8w1aPJ9I1zBT4PHX/Q
pfxEOs7oaC83BluodFYIQMKoXdso6cx+CgWodl9UVWkRKBTmZy8KsMYMDWUV9JRJ
iA8WEgpM3zUYLWSyI2jeQOsMsQ5elHm31iykDTrtJYuIl3E/j4dBuWBYW5f3wYwC
cRY+UI7iKm2l1gmgglGDSr7BpSoqa4n9e6QQp6jMreBJDdI+oRkjSAatnzW/Pju4
9cHoYy9ua/nf2AxFTool2m/vDQz6dO17bUgo9ngbpLxr2AbIIgxLBX/9zY72MBCA
M9So2CEFHoEnnr7igSMzKbg1PKUPxzJU1BSuzXLri4OEH4BI39yXYaMQTEuVWaXo
Uk03XMzf8wbo0QqLpZwKtpVX7Dk3Nqw4v6R2gZVg/wMUaOWQTIoIgIjEU/YIBbks
2qtKLQqeNJE0mg8MnI/RJgWSqt00MNrhOkBMM9+u3Iwy7loiXgqX2whRw3IAdPZV
ueWUBJaLNJTSUnV1VcRDssv+1Z5jcG7wNx4qGTrgHn3kTvOrMcfALpfQ5bgXcwaD
kBvw3HvX+ECGFlivXdEftJWd3+ukeE+4H6UdDCC7ayOQvPt7/pHLoKerDQAXmkOS
hFh58a2F9S9plfjYmY+CoNc9mf89JEWorYL2jiOtDfS6wlMv1BMZJ8udYqGU9zhn
6JrefEiXvmF8EsolOS9GswxRybEK2rdfWfaQKzq9CyqBXh43283lEUuI4gjWfx8Z
vof/MVLznBhLmTpt+2yiUR2TEyy3cWQ5ne7T5BfwmWmz6d4lvRFtUJJI1QR89Ftj
8WM11vp8lefyjc3x6UeLL25HlEl5rTYnO09TlKlVD4KHLtoW9NB/5yb0mBBQjIba
5dm1YJnXrGdVB9DMs5wMZAaHOHGjMeUyPA2Ihdk3xcQq+2ILny3jNqt0Vx8fi0Fs
zdITnYL5BETe1fdbP8TwHn6yD0KOBTmumbrDa7ydFIDWXGRT/4ZUqLkszEBIDpVW
2vIeHHmlu5qmsLuQlNADBfTj6nT12+HFc+JprwoAg5Lg1nu2RKUxpEiH8lt5ez/p
6fUQMJk38cKskStcNPaOBSVBP6qTKkXjHcLrSjWnNnk5Rfr1H1Lf+sr5igzBiOpB
UBvmnN0NeCRcpwCbX4/QwzigariISQh9TZW0fJ4aB+Ch1idOFU33dVeTObIpPLcj
xzPqnT+N9PYoKouJCNBQ1PIXhPn8rHexVW101Hg+W2XuUYfe0XBeMEbxFqn+DXjg
oSOZDak/w+UVhv6N1w8h7urAyDUbSm1+EHUGh+c3BQ9nbprxB+xtMCgUreFupXqH
YHK6jMaUQNM56xRklAZYjiGLwncfec3fazujueo/XX7ff34TlIfNTg3vBGKGFQTL
aIBfZ0uwIPoYYMIcxTBRraJ5dDcYQwdtkkRjoJKTSu3k3i+eDsUDBOqC4VC/cSRp
CjNggasMR/ZThd8z2JP0Xsfu0Fnt8+LqURshQKt/5g5veJBsk6dhSCvfTSiOgCLy
QWMcSW6jPwod0OYQlzXs9BB7lIg1OasLYurCzDyUnW4ueKIX710q4qnOm+MafMdt
KVAVVfWMQfM9pf8xll+Tqypcsbid+/Fkz33CJcAtqItkYmhgP9+SYiXeeN+9BYk+
9/P8rDIDYThFFZz2e03CQH3P0QP71lWJ/WHNYwfRYsuI3GJ68xc8MDfTvGGr0j3D
TBMuFnXLH6SrwwMdRLt5TJ2OmT+Qe6CpbqT/u7CeHi3wev/uNYiJJVXaZAnGru5i
vCCAdXitptUlkyZgxgfxGb/rUXARg7jC6CFZ54wMnLnu/gTb62kM8ACMIE9dpm4g
leFH2O0Dur+rGh2u4nvjDAzSzb1MiofeTlHF4qc0f+M3GArlkyiqbLeJ8Dvnu/f7
Y4kEWnnbuDbJYCkhkrlLCucm5XMuVSvZdAA6j9qDt1TvjoByOy2Ra6PpTs3+1Dah
UEN6lXVavyweMbuxT1b2CCR19pyyEO++7K+4jGgkjchFgGL/BAGhAVKfWOKFLMB6
V4aGLVeUxkmn1IY1qkngvTMcw/X9niTZdKqlWnHdiXEDaBVUcAr//PAf8xK0IYE2
OoiCvSp3WqsKcADwnrlupEjOj70hvmnVaiNl05RrOFIhLdaRfSVb+0klSjiCaEg2
FDrnACwAVSQW+28a5yhk/1un5cIDivEb40G7DeY7hI46JJNZKTvx5ODWqAhh+Vo4
FA2xfk701lxXkwe0UMZ6bu4LGRFcq4H++VZRqRI8ptSuacP/iyBz6k+RXQFBXpGU
FXqfjkSpYXH45QYtUufeQHyp+j2PK+X+1+Y44OYsEl0h+DoGzGbP1NsNbQqPrb+4
FDRJiqKWvenjJJNTsPbtFGPCwA0PSPjKbVOH54nsp4gh0F7ec7EkqCahF7Lc3WSg
cgzsQedVvhNeoywuKY+L2wDHM3sdtfnpugB9bs5PXEsivjCz+KNQZdI2wsnJPjgE
a1AXyd4uvl9hs2Je+rCtM62i2cGCIidGAsBPgdPlGURC0oR3UVYkd15p5CwGVmZ2
OzBe8BXKNGueAiB9evRgN1OIJcCiClco/a0LO/jeT1UMfJDfLLYJR0m/7W7k3o8o
poiLwRhntrbye8QBacYRwEtgJE55h43ANqLyzWQyqLaCebpndaMZYHA5ViDmIuaX
ahoSiNg44G0A6FPkqKkLkh0Yfa1LYIGsRQWlgPZSiMW2Oos2e+7P244JhkTjrPr8
En3avwiMNNdd+vIHb2FoFgKKHCs5v6cnMRgqVYhFFBG7g5FrfYntLAbaUT1xwpNn
d0B4/eg3B+SOpGKI7/q0IKPphEgaVV6E9/+8O+sm9X79dmDsc7B0B0nCgJQ774er
LqrhTU4dV1+bnCOQFk9zZNHhYFALnk42jQQkztx0SxGjy21yOBnkpzAqYHP1f5vM
4PppUfDLEb7Zg8COmEXjvw/g8EYtZAqM0fR4JIXtBcroVE9ilnPr0dzEOh9BtKy8
n5xUfzAG4AG89GVk9mA1PB3lRrE5HiCy5xelw6i9hs5ADPMCZ/Xti1txDMrmH08P
6mYYKcfXcsJHmp59m3AIH4FaFcXCchL64azJEMR2pDLL5p8vJ4pDYDWGCZQOHe4x
oMVruQl6FsTSL6CcJ52yXbeM7wGuEYbinzMeSsQM5UamoiE/0Bkmv2IVXxNRKgRj
QbZVib6buwoReOAp47Ic1XMcx+mibp1eaz9Asp5OJM1oobHpT84tt1NETsFqR0PD
3DlyEMkxcb6Ab31Kgl84CFtBC1BYv1HLvbRf48CjD8fmJ93CFFcxB4OgS0inRMSh
ZX2nboLRsJOc/jb2uGWiqpA5FUh7JCEwMnvsUST15a7hIqfQeWzyYnfmra8PGJeR
tJMB+z265bohEVnL45tb9newWkvOtfKcBMtSYKZUK8eKhczTjQ32a585hjCWoeYK
tl59WztG4vp/IYtfc2eVPN8minTWhwYvyxVDb91GV3zu8rxQ/m3svzJk9LweQg+Y
3kOn5UprFiMxDNnL28LNbOWzt+xTfLvynNKc5cK+or6dZmjAnw/MXZ1AUqs7VMTm
g/umbgAf9BarXYt9vHd58+h5wsllvEQkBlRv7VPkUQrZ/o25WbEozDIwhSMkZSow
WxPXoQ4u7pfPkDwm+e2I1MECTlW0slCXiQY3lo0x8G6UJ5SZc2x2xdmo94P97Eye
CJa8cX+2NQ1O9QZTkEi3mXk0W5dabtZel4NBssCFgsb0cg950WooXHaT2REy5Cod
K7TBrLkHT/qyNKEy4AWv5NKifYe2S56jp54ZcxvIVf3t5V1O/GYIaOMBzACAViKs
3Wss7v3//wNta7AfcKHVeUoWFwjgOKG0rZ653UZy6aONGb1hVKW/AUGCy1UZvOzB
9BAeLhE+250HWfpohzwe36cTIUMxLM5b9woExImPa+IH3bW+AW5XINGXuiSEyb4L
sR7URXBJgDugvzmi+6mdkU2kBejmJDcUpekgdcuxaVhCfu6Kqgh350Yo6e3TRxOd
kA4zpYQMIByv+QEgZFhXCBJqV6z1rYPqNgkUW/mGYKAHSsKPIXhA0YhnRzlEB/6k
bVVzgRtOGkgHi6wsVdjxdwHH8U7G+sZ3XmojtUK2E0ZpCeGIzwZetkPpXLxSFSpF
9JyDJFBHyevGYHGqiSjeSWfnQj5yNRk2XpJ2940cOlvbSfjN3jlgNtDJ8s11nKcf
C5Iq6cc0Z5VLeM4xDu72ofS7nJMsfK50cd6fa3WvVq44VSwfDprg03iuGVk22HJ9
0dSQZ4vGZ7XhcEkVMvnZNtcDAaxMzJZbvP+v2IzXhSUmFpqwwsDRsL3aY0Ti9a6L
IQE8EZ+LwXHgtSWsYgimwZFzVVJ1498vai7SWROoxoY7tkFxnzz0WBJD3m40pZ+X
gFINGcgnfj0OSdn4HqrRA6Rod2DSOaYHlagz7gLnwSSgWwMFHCHXZFU9XAt2gOSj
hcBmoi/nkdZ4hbPD0n+AcOuHEmds4r8CwIA01pzXK8RirSeb2puVzhAAeUeN140H
0rH8EugqaWa+JLuqGHsf/DkWILYz32nDNT48feV306r0v4IWDEviXCb6YDGzOnhY
FI9WZIEaE9hSgITFFajUBD1t2UA66gTLfZvlkYPYDkeAMplz2mKIfw/awIL2bxMx
o1Gu/yGdYzSAX1jAGKVeEXcsZ+5xnQOmxJNtXVaD2b080LO2JO9ki1qjFYOx+5Pq
QOqKyqWBXZjeZ6F90Re8tnLNnLbNi6JpR2Hnya0dhiRGAPUty6FqpMHZkB1Eoew9
lgvpNsAhqs+4Yg8dDSQYlNlMo9BgGxS/y5xowjA/1niN7KBIW6EdjbDoInd4Hgmm
uUHwRD9annv3APKiqz9YCHiHkHjOQe5cH1fGOZDvyYlws2gn3NsgD9Yojr/utRJJ
LbXPyB4KijF47j0sXauEctuapdwFjozIWGCQdWaceUKmDokwuJTJfKQS4+Sj9e9+
g36YJ91IiAyGZVBLondLa09+7ultNLxGn0+UbEcGbH0b1R88l9I4/WII3cQZXRRk
5CcgUnwTch5xGmB03/bM2LxksvS4wfK+nzgMr1KYi5KNI4TUT11Wi8v/0lbxc83i
iwvg/TGbebeh4lBzAv/P4xxEwaFQOVUbrRWZWrp2LbDL0TN8Ci6NLFrx6rQ9dMrK
kMREuPCHgY102FjSo5OklE5U/y70eqwNRnMTyvT/9vudKx/XK0s7rt5cneHPVsaZ
id682jng8VXdYLEKB5vZtS+TGQmfvyEp4y1m64bpDLb7YpCWNxVcjAoynQCdeRv5
x9wSQufOajpD3L/sZjmj2jnhnn9eBwm6MAPWEQp6Ivh6QwuPAWu76H27bmqTE1Cx
4ehLididrsKMQaIZC27JOiBzOTjVzt1uk2XGDfNKcIk8MJnqFsJOzx9O98fwUnbb
vazwxQcCMCiza+FnVxsy7QP9l1xmwbhks4mh+uYEh5JHO8iQ+OrvHlHPD9ZarELR
T1SDF5iRMrwTypIOL09qSQGyAP6vwoXTXGFDZof7HBU8e+jdp7axcNT83RnS/ZSP
YkQnZK48fy2vLJPNYQmGUvQIJ/p5n1966304Br3jfH1/+E5oZ0q1TG94IRHIJ4/4
IgM3oiqrOH0gRdJC42ab4+ds6fftKwy8HMGkar6lbfHL+1HBe0YmoSDQLKorjOBw
/6EUjeu3j6vldiT4tF5ilDydKctkC9hiPBgOLg//uEnbzNI7WfYnBOtJWSQnprn2
Wdka8TiRqJrDUXuittCI1xxpVJoruqKQU1xd0zy6wHyWKyl5OdBbexvnK5e5vGaF
qxcf6hD/eRUoWe+I4RaU3B4P9Hm3Bgz9vBzsk868BW8PaQhDvsO6VT3iOO/1TodD
AihtrpbcmtusiHKrJR41JMnnnwudJki+oCVsNLu+2dhhTy1bmIGhhMQZVEV9NOQe
8ZdlHC+2/FzQQCEmwkKgZWEm9TkGwmNlCl/agDep9xqJCPEMsySmTrT75l6GQ6CD
KoKAypSe4bzyRp5M3MXmt7jet/Htv253kBS7PazUMIgDmwQ5eAzc8la2+k6VctMp
sBN2xDmKJDGdM02AvMHWYXEghrmUkqLbSgproA5vBjG6ZwndlSZTQd2QQl5rE3Ef
SqHNW8DiQ9LL/+zaQkoYmzCiHiCVYjJoUEeG64XgOnsaRUxNB/8nXUHrmUi3zLAw
WpudUo5SzCfRczNGchb3LPY1cGlCXpTPGIjDMIdZPChv1dR0BqChAy9mNMirZjRd
55rbRNf3z4BDSQbR0KhCjJO+ymdyfs/ryVqO4j1Qv0vUTmQCH9JjeS6eIY+VywyY
pQSSfjfPVOzHkHZvzr5Hyb7B/W7XhF3CwTR5eoWoB+/5nUJk3L94AstXFJKw6xOz
dyY1x3Fqu02PiXvk0vDd5pJVSZwYHNAvdlJf1PiZtuwJxpvd44WHBp2uei3I+wA3
ZO6j3k7+QMSpScmSVHV8Px7qFsby7V7O0zNnEz1NWsXoqBc8bWCzvm66y81mduI1
Qy6mfYindPfNQnYuk8KfpsV5MeLgE32QwJ5EpQsPUzvtSlKPGUhuyX3H2KwuVOcH
z+OEJkj54cEJog9RE8ph3cwRC3kv8GfGjQedgdh9X9nDqOK4KXVMGaBKG73LD1+U
YjYj0iH0y6E2TEp5B//kGeTgRepZNLZscQjhUbLWcN64knCIryjvh/oJnojL6udD
94KqecYJL2usPQjP8Za99MvlGsBHdyIzSAViCJuTOzqkgoJZ1Fg4NtdCiH/bG1Ct
VO1E4eqWq3hfFD38M27m7PFa1Bta4Xx6Uxfy5nvYMu+azsqlJkWkyC41VVhgdgKW
1lWYaUrs30/+gGQgUo1tEGewQUai2qxtcVouDTUjJ43pC8U7HK1Ddl8jTL9QKXVo
C9GTnQB1FO8G7ahjltCSnw3uDPGlaFFNoKcnx9FXUmuEONr3gC5+WNAoNIawsrcO
VH3zH1ubSHZfti+hYRH0/6uUJM61GMV6ToiBI0Q9xy/Ms/ZYrdW2dXST862Z3bk+
QfmAayPaO7xJYgLpyRv2veGMK9ILi5wMa7tlvNd82BeXV/gs4xM+47hU8rRymsYw
Dr9wVEYJze6+lt150oF9YIZURR8MJa+M8L/toGaJfETXE6vCDKs+ehuLiy1AQ4zE
E/xVRFlc5//f9KgR8ptuXVUQwDxoycNjpfJlD/YyKMGvluTe7QAOlMudQxre2V7z
/x1K+3ZUxAFikqFUR8DZ19gtSDZ1Jc3hHX/S9aRMySV7xvz1t50J5XJxwxdO3JNB
v+URNth368eFi8Qayl3nnsf0IdsGDU38ef7GYYUumm5/hAoLgt/fmN9mcAQBn8as
jvHntTvCITm3mq9kC6F6KGkSNSPH/dCAcCqdWpcdZ1MFkFz5oc7zaBDwq2StbzcL
SsADpvnxGrZj83ypsmqi/Dxga6PohefWVOw8k8kjVMGvmOfb2gcAZuPs5LQ1FTD6
6wvd2nL3y26QG5fOGvVd3M6IZQ+nQdySqO8vRL4dDCr3VAjHqxRyg5Wmt9cH0S3p
yqsnzqUXZZ7bPEc5DrjeJikRHLQLKuQ/4cyH0yg525U1QtpilMRgZcgtzMK3ZZrY
IEuZsUWDgCGJeteU2mXXeSB5a+lFVuB1v1JT3yLaC7D1gIaSUuw6AvrLjMISn6+2
RR2ShgqrwY24New/C53vVcKd4DL9K9L/PrnbnT0bS8YA+KOwWn4cirhfblCgK/BH
rIbShLdUwEA3aVg18VFYtdL7SN1i5+VtnTH9HyZTC1HrWFAu1GgRKSYmQVpdoZu3
J1lbTfXN6z3TOwLBqiJf6ru4SgKqiKFyedDDaeVajJ3Frr8XF1/g6FVsLQKFfOoh
YMQekYin2X6cndwTLZtHFYD0gOELJPSX3kBzKMivZU4QrvTEzZ5ZXnznjPs45hPU
se/junaw4EThrXk9TeYr7b91rS5ndnJrb4K6d2l5lAIjzcyJTgZ9JKwHdXNH/Fqa
d/f+jte5Ohf2ve0ABQKhNxM/BQSUyUfYAoqBEGrzIkgzfaDJbTiHacieDQ9/bJvA
dzrFPYIwC8U91udESX9K9Hg+ScPMX62eNIOXRXGRkBK4CXQzggDJSmwM3WFXa05A
cfkP/z8NVrkHDib+btDwa45o4xM94J321GQlLRaMeUEwA0KChlqU2L+fwefwSsLl
BV6MkwpRTg4lTy0vrniB0nTbOHUgmt1g23r9tq7GrlCitfeX8sqU8nNLL0PpqwpZ
qAqRLy9q9g0M2Zvz4gCNIAXyVaECH5oB6oQH/Ts5rFw4Z7rxM3m4mxqqlWif/PS5
JZfoK/kop1yU8w6kfVlf08iuwklAl09+SyH8cG4s6pYnPfxBYMq1PIA1BaJtUFtU
bQ0C6XQQpkvhOEunhG7y0SCiWcpW1ZJ6dWNE1snh8/wB3MthFYd6V9zs3g9ZR0NT
0AR6jCI3JbodX1EWNkrmxnt7GHxVCjuzpcjHiozv7jbDscf+4aCdCkZRWW8CQJ9w
/OiiIs6FfVfIp9KVFT7YLCyoRk1itUwlMzLYJOQmr4JJl5NeWfZqXdBESwTWHe7L
BGKfpGr/l5cGak3krQL1RNN7GY1noP8ucGEGQ/SFWrUO2z1kpWDNzG64zzIC62gU
az5EU0hAXog1Bkcp16h2cgqpodHphp+dcHWd5JbNf1FTh187+LVDHn9xwsMO9JtD
j56rPHfNa+PMZTDcgXP4i7NLyJxrlNTJ6fnug5RB3TfsnvW4EUUATesTcgA/muSC
xC9XY0qb8bqkDRN0cBe4IJuF25AWYSxR1qN6ebkHwQ0MVXyWPZ4kPSrNIuBQgE1r
E795rOQEGD7lXpggrzIrb+boKytHXnA/2yyCns+owDhpGmmtCsh+VSLtlXIlh66R
2mWgr/dqbzqTcM3Vlpd88fx712QoADaeI//xVjq0ObJAGhUFkrUNfnejMl4QxlGJ
N5tYQuMj2a41Yik66G7en9Yag2B4Wd78GZtBS/KwEq2YDSrCjn1jdpgSaxXM3bww
+z9MqDm6a+Y4I1pE1+/oR0ECc2Eoqbb/eX82/SgnGXJ4sn5m4Pza84MCJ9bMrbqv
ZfhW+4IJga3NdYjpERo5C30QlbVRoCOQ26n644dY8Co18nzO9MqRxBBS5Brs713s
+CyUlsZ3C5gRjaByX1skk6ClPo5GMBgUGmQIGf4vSGn8qfwCTNV17j1objwz7SNT
a+vm54zwGW1c9Tu1ThSw/bmO/A24wvHtOhlY8sM7e1ihHIzdyhT4d335k9OixLB0
toKRpc0oqkDCFum0nE2FRnf0EhIRjfLQvQisyZxIRyo/ylUMxZD3MSzm3O8I/aqZ
VJfQtrjCh3FDQOkO3erur79N9FmTDzCOtOcM0ksLjiM4mawnhWzNs0upcxaPZvsv
mB2zhKEvryNup1zxGMaNa+YFyXtWsbhf994MKZpmDWxd70fSBTYk6UrxlSzXTkfC
jg0iApKX/jTOPBqgK8Iqa3uc0VeoGsfOsFHX0kkHFZYn3deUE10voogT85WYtUz/
XRA+hnmkLzPxigsYOYgHRUFAcqdyd8gZDSQ1Vmtoe5XF0rQhYUQSxcqs5Dy7otgx
R094+1pMK4osuNtHZEHY+B5SPcJPJkREeDrqcXt5sadEtbcwjRFkaFw6b8G+Xv3c
0QrNwv6BwVM3kIhAZTIymcQiUeBqOCm6O/JVpqN7asQTCzit1nJSKeQrhm/1Snds
Zc6P1Gi49/ddkL0uWJe0gHFhV6dMJSGOB5FtaJpcr//bQNpnacwk/9amLmhehMcO
zfd3ODVd4LoXmEcHqmuq38DrrNmgKEYiKRxO6EShSudCiyAU/gW/wR7FU787vvjE
L1I2eRr9YaKoW+4Z08OrPe/+JAbhrU6VlDKztMVMRw5etAvarRW4EUH2puGKx5iY
D2PHX6WQX22INr6bqKOhBRksScDtCXIfdyqFna2Uwv5Ex0ohV514C/+r/J0w9rsw
tW800x6+LkkbbizykfSTBwge1PM7hQ3nxvermBGQ39/CULfqvr4aQpTTjmFkLi48
lCQTfrVSeLKEVdj7YEavparKq+eI8+aXqxPGbc9aZSbKb2EEhL3UcUSFscKlxcVH
xtEbQXge0eANnwA/NZbZxQ7S8ualdIY2rGLgjtq7bn3OybzjMPm1vcqv/qUqRDKE
hxXWzIHCXgdff5Ywf4tDLxoeRZ++UhWx5+ugSuvFN3zgSYB2uMiZYPA+TToN/2rv
FjO7z5rNyV5CN2HzS7oCJHahgeOcC/nhHkaH8FEjQ+kLyzflS9nNjU8HWpe9H34+
S4ZgcLbRTPgwmrz0pe+GhDaWAQWYEQonOyAE8OE2Adw4mPaRRjesd/yu0mor9U8O
qnKFQOrdWvFK32hHtGJZKg3rZVDrVCwOOsxF6jFzm5oJLwNzUwccUGk4eVgA0+Ps
N4mqwquPzTHcv/m+GNGHbnBFmnFIkZeBycO3/fuM+mQxxqU/N4xG89Rh8h6hbJnR
qDcZm2y9H3DD9086IxYG69NAFIpLzlzrwHZfnorXQpgRiIZBnTLkfZU1AH3fRBxl
vjoHdG7ON8kQDbvSkMEWYz8yEbO3GRYIiVwZwppPd7zWWjoOoNwsKmQGX1+2WMCV
dVQT2cnHKUXnKOYR5IderAwoS3PVO6cqeWpZUcdC1GKFhV7ZlmaqsT0q2XPAWh0c
v87j0g9H/u0madC1Y4JOizx87bnLj0t/D5ppsKnB+QVtHE8nQ/pVUfjkUOb7qWAn
CqsjR6GJsjPFKO/Auc8Nbp0RF2fdvCPi8s17gmiBz3xEcttdcVGmvAT29Yii93SM
nSx39FfabYBsIIbrzt+NEKKYSLKDHhk4RkgEgSeTcwVjly+tjcpFFGHPlACgjpAk
d2zqAMmQZX9DJRNUvIlpXujiy65PWkobCS3h3VMkyenXfVPhda4Gp3zMhcWiiMa8
1ihYhxletUq5Keq8c3ko1mq6gIcgknl7Md0n8Dql2yE13DvdrM8ie+xYjnVAbxk4
V1TljYfikQRKWcWEwMhIgs7mGP8DKnBh9jfHDZifz60PE1ITjvq5uMTMuvRJZ6Zb
RGCGsoz6Pd/5GAGlmtunkfnxMFGaLs/3cT/fTRJ57J2BodQTwBCz6IuxmdcWWwV1
YC0rRB9SacHJX7dhQAWr8ayRUtSzKdFon2evcPCWuWjC65Sop4ffY7NqkARHkyow
St0oq3MgEeagEfNOjp/8mYeG0U6MbAlhMRkXIgBAM5VSouNZitxybyNW1t/a1FNR
C+CItg5PFlQ09TkadNLah3VuqlXtokomI3iKfADj0XimypyciqFkjcgKoTU8ehqP
zbc55UD5cw5GPO7NgmKgKP06wSnjnBRryqgZkbmxPAXaXGRZduUzbvm2O7uDOn3d
2d6kHiTJ66v3y+t3u2AKcS4aXFGMZkC7wcPFMWfyeC2bLGTp3fBw4QNaj5hN+nrb
t9NSZZGeZvCvIes01gwmgoY39NcW53oYKz5owifCBGutrmMDxy4ueaZTggk70K89
UUGmU+YSglPHF/IiN1q0ogoCPAd1dz9qnGOCulqhRaT8Si6DNPSiuNYHZBuKiRnP
lmhBRIW/HhzaGtcZWLgrR07JokCwfLszDrN1V2htHyStitdq6gLo1mNU481ey+F/
Eh7NBX0Ky68mUWq0G4cNZNe9Q4fpbBtCj61sG80413aAI2h39g/f+l1hFAsc7vS1
C4KwzXgjKlBwRHNnDzJtVYx9UYttw8Ze+5bKOyfusJ23ZN+yMrBebVtjJ6yXox9U
LFJR+l0Fqp2MeOZa0hV2SBX07pYhFJ85HMfSjNThTo4laSjJp4DIszoGWpAqkwaV
50OeoAmTSdH8Ppe6XUZ+KpvIpW98tcglqNO6TnBq8vos76+Uu4M/AffWfZxNpPV8
pQcAzpHt16YQsE7pQtLxMOCxQwQdurdWtGZGvw3G1c1zd/yfEyvHnsB5xXCtWkcy
PeImqKLAY1e+EvTuxJ0rQPKl5xL/GBaK/q52wKX6ZPfyorwLKDvtPU2kD3vLX4TL
qMEu3CvQuMUPtLG1iIqRPLxcvOL5ba9bR3ghS1ZL6jrCgBhJgq6nNOqeVajdl1m8
P6lLNMFyZVGY1rc77SWItpaP1iJHpRzgnKox8kGsnqJm77LKYQta28m2LEoj7X8f
rrslC8ttJnOtH/pVqMx2X5HuPCqVZj3hREJwoHK0jx3RSo5vqJ/2pUYTds2bU2Ka
IFdG3yQRajBeySq9k+kC76td2QuhBgbY52IQYzedhG9ZOluStHQ6MEmOeWh2cSp3
3KShDsH7UCO5w8493lSeWPqsjH18Z4raCZGCvEKO+NhBkKPrpiqbBggQRw25MmBk
JM0JgtBEtEFoLClWIz2/CyYJUSsLbeV+OUYSbKX/pr7KslPCfS81GF5JEJfRsch6
r1N2iPECFO8Gas0YEf2tlAsyebfry02ImLlmkPoBGgfatVwrT+YvUoczjBaTGRxI
1MxCa7PpBb+FI3Y9PC4tXyrg3w2Ye9RQNjQNbvoYQrW81a/DGXKkSuOIU8ZTkaZf
HvY3CMjdq4Mr2/56mKB6RBJUTFSt2yPxmsriBhS+5BzRT7P7i2aRAjrFDY0zBZ9M
0+AsIxBy6WfjEEdD4SdlJ6s018iFVdpq7TPWxw7sOUR3uOSyqada9/y9nC1xpKlE
/fyKikPzS/va68vgUFnqyqXVb/JvU6ey84LoAWeGZYyOsnB7Rmc9nJYOUpxdcxRV
+5Jn7niaP4bx3MP4ghj7VUIIMRFe+mUKRkOhExv8ykC1GYWDxUfz2tM5P6AgkBvc
cUE0QODkX9qfZ2EqD3jHeQMJs/0IbrMRwmDUUtmeDD1rW1SPK1eMrHJttjbDGSx/
qosh+O56GMaimHbn/jp2Dw/Tc1mde9RkfWdNFPN9xSc/zC7vc5H0v1LHEPoYXQWJ
QdgKQdz4P8ANWnhEarEgvb/u1ynrTAFtLqdapHV2r8rC/+SRlc/gTfX24teO+VXD
ZZ9aK9knsjuJ13+G5z13bxDKpCZ+LnCdLF6VSxrHsHUbk6+7opFDZhkrQubWnM8R
2fj5qu/dIqcxIemgEp+iDLUTWgK3+H0YNLO26QjJphtzBQb1tlEzAOvCYck2WX3A
AWyPvbdZy4jcVmAPTtbv1IaVH7wCrns/4IK9npPEDf6rV5LqMBN2Iv+iOa3ZOvMw
zwjLlhT67IuM+qdjyD6w0nHjG6D4P6hrAc8ZQVEdstvvoh4KWoFl7ZnxoHsfHPw+
IW2FQr7WhWXf55x5G4gVsbs9ft59rBwBcPNcXTQczixt8UttxpLUk/olaRTK7zXi
+pCO8Gla1ovnvmicB2C1fyNFSSNUIYoEwx0TlIuZV2grhFp7XmsT24GE0LCr2mA+
FZ6I0Sb92E7FbMHq1zZnKYV3U5teGj/SQ6z16DLUen+i3eQf1sCHoOMMzqWr+Ylo
aLvpXQ/rtDSfAdLQdKbjpaeHj5kAfu0jQ8x0lvAiO9l+HBmDETzamem1XdhgpzLf
lJgf2YB5KWKO7Q5LpgDek4gAd8x+gUtt8jA+QGcTKInyfPlpftjjzkhqlgVapsYw
4e4nmGzsWAD8TR+JkAyP2xuEPZbex4uKf9MxjJa01jgoQAxgEyWZOmhvpn/uBg+Y
0/l80dar31d30KgtJ1bmwSUyynZzS6vefI3feON1CBTguF6CQRqB2xXn3D/reB+J
puJQkzfSGC7FWEXJkESKt4euDZvSfajHXGqC9s3bEWubUcJfKf5+HcO5/Ka4coCd
eMA66+MwTsr7A97pjYyjencCQqs4bE2nYH3zjXLln1wiWNzyK+8l1UzJF9mdexTc
hgC+yHSwtlOxItYYFtMkfBhc2J3jPYg3gOCC0+OdEKXfvPvojNJ1eGX/SHmN0eNE
0WZ+IqYssiHzltMt+6f/WyXFSqKM3wmut6Rs7GFGr/u4gYpnKt3xvt07xDCYg7Ec
F4tjWdIBv1AF7d3nJoYA/Ee9WQue66wDk+DM9evxYm+5t3QGNI+ButJfgh1IoUYF
TKai/z81+o8u7Q40vlAJ7Go9hm0tM/mhMaIOPKwN1ROVZF0tmZf8ZRP2UW8jpbtx
rNCKkYBjBtfOW8kqVV0GYBdovuhG6gVW3UlnnXAbVrFbqS2bEuS+9b8zX58JTee9
ZDP/9E0RloD08CDybGMdgNZIDSaZIuAzRRpeXc6SyISjYOmkUalNPm1LeueO/afW
3S5CxvshS2tGHFB5W0lAFXmmL5acCvO8sa2iHDfELAnvd0OjSecNWPzyMbT9iC6I
UM+bpSp00aBnOiBh9kEZP7KGyRSMttQWu0SaDFhJzovJK/LTGomXfliJz17rNjA3
VtGl8dq76L/FvIgaf3piEGMm+Ju2g4rUYMAQV0N7loVejq1w4i5rOy3pu/liDqEm
xB83ABq69/FQdP+G8ocIhZwKt2enpigI4CalKJ6hP5KE1u+vqDw94p/BLOZiZpnG
PMJHg1/2nQ55DkE5k1ck+vixx2CLy6Kss93a0hh3l9n96eVkKDtH9Uf7NZEVuPu3
0IxY6IqwSxSO1ho4DagCzYK/oemDoILi6a9j2Zn8IHVP1rn2unS5DhqUBm3P51CD
0k70F+rAtkqPrk4vB3WCRjB6INjZ8DTGXKnS7weQ8tLxS93z0k1xtIsOAnuE1bXT
QwTZnxYosIsGaFmJ3HSW3XQJAWzAegdJzVFEk1i0xWScEnT21Dk5E4687ltwrPy6
xHQN1RvX7cpjjtAkTBWXD1ivIBNIw16On1l4ed+E8TAWYQdRg/evrp2mZk1QrYFG
mJKxLf+nH5xzaiap3swo9PsOn7skUJip0nO6ozyTl12Cx6ARN8xGSxUnsQVNzAB1
Jb/Ygjg3bVnF+onAYtTKVBtO4NeLLuFw1UsZB+DP/S5VO+ZQGW9himMGKRIF/wij
N8ouranOClcSP6ll8DJBvgeN08VURBvqxvhUsaOoJ5CsTvU0PDxYFu6lffRDLLsN
cj2aNHFA6Xir/1PZ91F96U5HWpE8iSdkEpg06sZmLhPrzhEPP81p8372z37tpVRI
FCR6r1NF7wFE3WEeRbsvsHEH3Ddx1rnpJ9CqDycUEqk9xw/vZydui15k0j++KCnH
renVjTcI1nbtYVul/LxTnraOqaPNQS6GZROPlhBTBnipIzMGoIGKlqfzZADhrdck
hez1cjQa1O8rwu/AKgSTTGriznTGsouSOCcsHNqMSR6aJ5q+ggC3VExzRhcjW5kW
BkVAMmnXMzEk6mNcEC2pOozmsZueIlWipgEZb3o+lNk5HAW7uybIVP6r7T64FV9u
hs05P7G8Cv4rKo4s4nyanFgmg/8ByRuEqAFiiEBiCioWY9lW1gF28oNecuck7RqZ
bNF4ei4dkrX86YcKjduGIFMt1lRCA1maII/N4bcg/aDnp3CNcnDaV+PknveAPHHL
iUu8sJPQostD6RTSQFrdZNL2s+EwdP7bDZn3G2rrx+m+QkUofOf59LU0zN6KG2Ra
UgV1zA756ZPwxCUBtIPIqJZvwJ5iIJk8hTbBm5taMHijpzNqYB8tcVUz4OJ7ot3i
1S534n4LZp0RTiQexlOTW3DAV0lQosY8MZPgTIgftV6YO6GstgXBfS/wFPX5/Vt4
tHHUK0eiKy4Ssx9yRuD7rEi4PIz3WVA9dVwd+rECv7hAdthvCltNxNXVPjdXag1H
H0cKQFnFAi1CY8atWvAuqMsibTVB9bQxZVZ1T/JZsgimjr+aTO9HA4b+62EKnFgc
1FuCN1VEDkB4XO4y+W0C6TJgM+PepW5M60LazJ8/exV0DaTh1gjM13pLWuUrLmLw
6PEccc61apbYVbCqfaLOQNyRDVyKHiZSnjtwVXAh50MpE1AAlfx9po2pKfkyFDgX
hFZ9X07hD4mPZL64bBRjyPGzLh01KN4X5BdGvDRmDO0fIaJVT3JntWwOo37AuHvZ
xGubHSyrz/1+tkMhzAGbic4I7nJxbsviUhiQ6+EoLNLVG7ldslzoHps9tauHhqc/
iMVOw0cXgKP98Ytm/xi7T3+uWTQM28TyobFtBKkce3d2Ng1sentpnSMPy/qU+0IB
HQY7Gud3mOlnS4rqmpJJbcsKicxIbx20FjLDUjQfG+8p/MnH0Lfr4JIAUVqQ3fry
5561J3dDMN8GHc06FHAHJgPrq1qREnbGwCkmcIzfZHgcfrpMMO8MmPHCFmmmV+Uy
sjTBqd1cxHcvpnBiJePsnpyZw65nQF7T4kJzayLWhNdUQJRPn+Fl/4sQRoPctN3+
MTHtU2+1fzbgwa62L41PXf0wehi6n3E5/gW7DhHoiH/DNPdvDZ4PAm3ugppun2B4
PlFAbosdAddMEiFTNFvdJ/WefrwPk0btK/Pp61aTKEIzGwuCjkc3YiEyvbIUcNpe
BWTFAu2halIUOt2FIg0A/73APCGhvMCIHZEDRbK+r5dMeMXpqDibhzIblHczMdKY
stw9wSx/jXGM1M67L73mn9U2QClCf7yVB7mcjgpuyPexwBnKdmGVYCjhWx0e+S1t
r0GMUq2n/GxuPWGbxz7w1vEC1UHDe6DyMY/VMNVDWU9fBzVjvbOL1zcCl54dcBZu
upPdRnHAH4sCLmxNXqJWBBMpQPXamTTT7okzUQENsOGj48IK3xKx5Gs6DlIsSZuI
RMYvzGjtPAKGVd4jtNE3/KbV9kmVWlhD56wjYQz4N1M7z9RBT9XVxgiSHiVkqR/C
w9whhFQnHDi30M6ybopGx9lqD+aSPtYHbWX8+yeqEt8rMexsdHxv1eOjR/4yI7vY
53mRgQDOIlKLNeOfCN6ja03+K063rNrlh2sm0p+dTb0VrG2wdJIkpBNObez7xvtk
pYhYZNnYlQMe8Lr5uwgd+tGz95I01szvBkLySm8FxDtwc64QbLF0PcWEnua6Ir7V
5bUt0zgrFzCNlrETEUCWzzxGge/ansDUAe4SMNZApvyiQ1zTPu+Yuo4K6H0cFF1i
P2x3+J6T9E/UIqBwluoM93EQup8AwkLNPWPdzkNNxbFA+PbtgZjxnCRNi/LzWwPe
K0NouaW28BadL4g8vbjCNj9xh5aHPaEU7VtH5Nq9XdVHIxitTKj7C4ILv0d4I+i4
88IWYw06O9PKaVwW7N2ccxoJkNZQz0WHp6ZjYuoDAzZ+JDKxXaUqvXpWKmS1Qvne
hPq011MY5MqovLfxGfI1oXjz4g/Y8//hKbVofFTygu8q2nfY/adM6XPLBHD5MlYJ
6/IiPzWY1ktLUMPDX9aYgMrRTPGoKuTfuzCZUw72OTa9ypj0tru/+l8UHxWAQiHl
U/Re4xhv1VwxpAqHNHTWtoWs4p0PdMpaGsvFTLCgH8s/yVDagKFthivB1YxcOJz1
hQXr5bqqNCqO8iVlxr/AO2lZqWpitaQRpYmdQRhta5kb25CSUFV2aggP+srd4G6n
y6UnvIY+734FAT7UGRyPFlCWEQmHIuB5QKUsIrUAmQiiVB7SAf1mlKeBrLyheNW5
0ifSYKpEY2F+SQuC/E/AoNti+MoFQwBW+yYMkFlmeoN61eqccDHvhyBA1pgoaxg0
ZgDC6OpZ4VHSXXgQD4abtW7aEmNCcKFlhZRn0JUv3j90pUB/tRC4RLncyiFMaafr
GGpJQ8L0f/VD0VCriQpwLLmuSm43Wxcov2Y38jbGAmc4r5nvzP2h0HuJYtdFzSeC
wWy34vtZWgPaXJjf5I3AP6jDqEXzJHy/XUplWBmcZVQN+iY128sT/5/C/vs1h+S7
1DGed4SiQXgGbLa5u42xRiQG6WbFWnGQrA+ocNdkoonIj0PHk00N3dF6iirE0WE5
n/no57eBkDLYixbxBgn29KmQ5aLUy7FwtGd4jV8sIEMdK6REK/AQ1stv62gMgDe8
Z7UnNdf+wiNcatNMznQ8uB1ZwWyO9Wi3NqqXC7UflA4ws0EYSWnHBe74Y1ByVzbE
wH+mVBM5/cLOiMGmqYf4sQguhWsmIW9VnxsrHOtWuPLczumneyu9S4pXPWD+0SzZ
Se6UnwxlZFdZ16EzehcjIppi9iea+v6hX6uG6sIQSDU7LwC7VcTqAa7My7JnS3uA
vAhfosi2nB+5uh7RQTSJTh9sAm/8BLcTNparDfix9SeD6HPgZbSo4lFJv1RlBq7M
Idp7szfwSRqldm4cYq5NXxtPamdRpfqKreCeDE5M8Uz9tVzOuh8pQpurAX7FmSfG
ib1ffCm5dW6l/p+LBnzKSRFTUAKOW7KsDVRUc/+JWHAtdckoxrpBq/lkAOuibg9A
T6I5MRxZ1i017mLqV1mJZuCDRNlF++ALmQiH8TsICqujZhNcWkEDIhxtuq6kPiXV
pDEKhWOcRPShQLdcrkxFs+AFwGvofkVDGNFyZjVyxunaNLzGrDtKTkc3BfkS6Z+N
YC985cPQntusfitIKP0JXmMBwI62F8ghpW9SJR8ODZwKDIy1yQcTdo3C7XF0LyKj
wbWpgy1+aixiNhU6qwJg23sBvJUxbz7h5RYWpdqIEqMUKWGxOSBPNife6eeVTVBf
PR41lIe/NSusPoH8nUsdKxUOFWVFSXzKmjet1dIS3xX1F40FTi5tpie9+Pd471jy
a0HNs0UmBpukpNlIgTR2Yhn/MRADx3uMcy4jtfhsrgamPoSvW7AQOH4ROjitjCNw
aAB89vF32UA037k236kc11aH15f682UjgrxGst6EiYL1XSeClMAalv0HVyyWtkz+
4apHfoLVzKC9VpuP3vyS+L9NB8pnbKHA7kISrEFBt3rFrPEDe4ZSxn6qReFg0sZf
Q2NUKRqE5VCkTKvGcm2XkYR9FhHLFx6aXkhGIduByZoSFRoJvVsh4WiJb+Ivnf3y
F8ae/u8qYIOa2rCfF+9kOc26GtnU12mQATuJ7HQL8LMJK6h93wieXDMQ4iiy7CR4
51kDntnqruYZe2wMOlwEAcVOtPEZ+JabqPvJcLmVectR7w8IvZnp83WTsmxe3qMI
fPfu+N5K/lrE/bkuvngxjBZjqBOx2jQMIN5Iw9ALTpQnzfhn69fwX6udjgk8FWAb
IqewJ6g4/DZ332UmRXNU05640kEEdKS79ccheUfpOhQWix/yt2FQgIiJVwKRyXKA
1tGFbHwu4+r3KnijJcTYeQABKjKrnFkAN6RpX9AWDi47Bf+0sk/ug0TZu2Rd9Qtc
xa8lNUu7WDQpdkKnwmIG8klhQbQbK/GpyYpUSpiWYO3dzfP8GKVhokD7DRSx6+4x
u1HJF5DbtS0BbGC2QJyvBNieM/Qswi/WIVwCQmPFgQDNQRVCcKPIdm/wJ+c3qQwf
YI1Ag07AY8hvPAZFX8w46dLlUEvHq0HGlCnexLDBgtnIy48YE8Ja6H6sc8HtdTN0
ZD5X4YkLompETeIrnwjOEbUNHgSbNAy0EghdPWS0Xq4Cge0HpMda0KGKz8e1W4UL
utMi38vWF9DjMPAS+BdS1w0gXUFqH/MAcYasOl3wTsmjZUidpqRuglk/gb4e4tMr
w6OFczrRK+5icw7afTNfXq7JoE0saYf3L7JSb8uxHSkT32fHjiD4LG/Fi4L9Fpnh
4MNePWhmhiuvvBKRog3JBTFCHajLAHHSfGfmsFt86/L4FouYVwJp2bdH2pfeKbFi
R4/f/ofZ8HRqTPF1fgplAZj5jIYmTbMgxHZL/8jfXKW0AAgVf9MQivYgjVvwtdrW
bb62JhlOCE4eKA8WXwbzx0IOP8Y7QJQZF4OAcA7Kapz9ba6Ods+Iw4Hl3B4C3Rf5
GlBrXeoeGo78PvRXT9gpQ96vM/ClGQBQn1BuVfWugU1Ws/8RB03SA2i3j6mS6HiZ
tyQ965zfB/dO/Ij4WukI7n5wyL6ass9BxgoaJ9q/i7E5OMX3cqWqgyqIbA7H8xGt
87YLgNpK65cpCBW8/bMG4bC7AbdQxi+Hz0Zev37X/684dWX6G/zsjF6F08kcSZSa
8E+qB6SUvPz9Fsyc6BaY0KICOIkjEelHJ9OEICRnmeURnIF0Q9WCtU61FEKlU7+k
uI+J4CIN0WJg6Wb5q44JHNxvsn3vf6JwFQDzobNxgh9bQChUc538mGOLQf+uVbjt
6GJl1kyhZYfXweKvjo4EmBfWDeabgO8ZJxoWe4DeZqt+uzuk2MCARkaXNJmc3x1x
4rbKscwyaKB4Ho5v6AYLC9TNPWxcFF+T5+piz7u4ktrjh2dbZ6b9JWi/T2kSglJj
3WE9db97QqkKgBT29ZOmlO67mOG22eqxiYfrXi5CcWmoamCIW6IZzY6ByCh6PnwH
Aht5Vm5KBOMP7WKJr5LmFlP1kIOi2zSE/uMvcOW32FOy00z0zqAqtAYRHJJzsJrU
jEwipKoQkXF/kXJT7HIY9JmRv7iBM31N6ECSRUyvh2fTfcL6jdKERuqknxeFBURG
D4Syk+xrg4Z2Ym18AuyIWiIJ7mgQvFtWNKwvM79wk9V5b5sP/PwlV9wwuzwofSBl
set2WwTyz3YK/TuHpJN4V2YF2Dlby7kNPP7k7/y3voJDlbRaUSxZt2cGp8wqO0p5
1igIO8a/FIFjqFXaqE2gjPjHXYFMB11g0tHb1MTOrrMeyp1JTtZlRRTjQ1maWJoe
7+s7+t0vJVkK/5p0Nud13URielm42iR0JqefjaeziJxWQCuWLauquqSYXEOVo08c
LF6NOpomm9lnjaYWl+H7/tJYfX+lMGg6sSsOuY/9hM5jXg15f3FauRl3BHASYvG7
9qDMQir4aXBRU9h1kLdv24iIPGOsjWVo6/AopJrafpZx3qYAULLMW4XdM8UriOH+
ju4k/XTCROGk7uO93tJsNSuCY+CroxM5NoM83k90C+URos+OxQnCw0ZNLluXOKtk
gy1UnFenCs7uh1naV4Hy7HRKxX99kv7djPwBP/lPy+5GekFa1UMdEMsrJd4z3B/Y
tucFdGf33cK/kl6YCGpjoNXJcyV2MmIFju5AeeNhhPmNTGIpauJuFMTtwWlmCn3p
1+GFGTi+v8Fqp4bQSUd1nqeREG43SYCskn6aNkU63jdqKUJgVqnhooWztQKnPbUT
7qyYHN0OALsOLBP1sB8IFbOfiCPMarXKHYY2ci2oXT+IXRMVN5vp0Ly3l/SWlJ0n
vpSFyHpAgQ5l/agmClD9SSyFZp6sE3dj4Qr6lhW9WekPj2susK1tKSxopUXWB85q
ss7v0L72HyaBcz3dfxxKRJ0dYCepwHKlLhpgKO2IdbOpr2JewlcaLdIRFbYyOEtm
dBgrWQ8EjNRpU14HSwL6CXUacUrpZirJtsccJrvmQ04LjExW4gxSyrZbAeIX6GAI
QkpkhvK9g2VG3JXljX58Wxpyyu1MLL7PuDfA/EFkU67P+0umOlXgZ5dpXgBcv3NR
0N7TlD4gMRfc6xrdb6Xfl3qLQro28pJsDdOyoWo5EF7csL28O19tlJDmLvwh72AG
IVN0sqEz1OccuEnmQJL5KM+OCAAuj70hCakdD/kV8bsGrp7KBh5NioBhfe4Cvwrm
Isq8t6nDDwMk800JThKLUrlT3kDBTWecFs1NtMQ/GlkZxLhCzL/eWV+94LcU2w1t
`protect END_PROTECTED
