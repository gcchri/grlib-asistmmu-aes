`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UASO96mH+hwRnonthgWg46U1sfihs2T9uG2LtRyI0VN/lRKk8MlPByL8uvHrLY35
MZRqnNL0o/dURAHt/WJouY9t7vTB4DL/DLHWeow5m74LS3Ozt8HxpFLFtXz+xKHx
fyDoB2wIpdfw5MWcrGL1ADF6zhDPJcW+InmuWSh12nHCM0B3MULDK/AklnY7rBY6
DWcw1pFR93+NEWNpqoV0uuzgXuvouuU+vcx0xOxMh9i1X3+UTRGaLafWDXPmuBwH
7Ag0+4yn+s/AqYNYEo1NE0Xi9F4449du5EP8ZSW1wwtbaq0D7NSMuFYcLF2MGdOE
zyk1Vh9QPaSkzveKifwl2fPRIwaxvQhCTA3vFqIgRnE=
`protect END_PROTECTED
