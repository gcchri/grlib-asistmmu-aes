`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KvWYMR5LRctJoBgMGYDm6laE55DhK0HoudAPdyTLRvfz44ZX29stHzj2NIYP5qcy
2X6BuR7HsuQ8IsYF0MS4n9htS9+0xNVpQ3to9KXV5GUOBAI+G0fl4vQWDCZHDPQv
b6HhCalbMyeDnPOVqbWKmUYtxwt2ATexk0vmBv8U11kpREigJPcp5h9sIDvwz5I2
MaA3bBimumogbD3RzSz27Oby9IhAJGSMkZ66xqOX8ycF+B1C+CINdzu+C5/CiZLc
GGqdGkDVONr5sL9fkcjs6Q==
`protect END_PROTECTED
