`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VrQwIk0UZG2NWG2SBbmwMihFihQTzy0tMj9oQx6IqfD+rxYPvcwh0txOhMqAY4yk
i1GesS4wGif0KTeZfXCT4n7oJ2PkdaGntQl0O+lVpEwP3Yv+f/215zEAuees1GuQ
qemAqwUtOhWQGTIJ3mmVCKKG+nvnUBP1mqM1wlRl87tguSnIcm5GF/tlSgUiGHb9
b1QTAujIgfy7lmZNDScGuIiN27y4BYxmBLKS3z97KmdHEGk2ydojh6GFWl+03G+L
JWyogAMrealTnw+/WNLibKj3CQzsO1dF2UFUHRB8On5PMkDl6wDPx+QAnkfuGzVn
LTbVhAtgMaON2tMFJCbomvaGeSzk5UazSr54Y9WEMpNkKwo+pru156it92ZDbTrs
Dhm45yqT3bchpXJRQaSMOM9S7E+winTQb/0ncuImI59JN+qemTiwe6X7xnQLjtBh
CicTrnVCx7BfCtmBC9ELk1S4HUu/Nmt7vOGK6iZ4e9XhRalYhMkGSc/UJaHOmt4h
fnzJ57VsI+YF7zkpAa8FoeWFDMemb4XrJm+bCZrfIM67FJeCY3IcSUfR4E3APx8/
9R7Pa0VkOTEupWTgwYMA+cZwqsIcrYB5N2blJAJ8waFOZ8X7uVg1tIi1i17awwgJ
S+kP/zDeuxcr2uvDkpy3bqixDQlUEvcnjXBqyKIFWtKJJSZI7Jwp5zXf4g1ATQ2c
1qWQ5ZIoPogOVwjWJqR5Wmc/NKvQICVKZsHB8WoqF0Q=
`protect END_PROTECTED
