`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OYW8a2+/NXi/nC+F2UkiRwQ3tM1JgLoQob7dcyvtM+6wmGwQsWNC9CAiqMYVVGgZ
AhBizLGUiuiEEcomaGODs5bs0N7sXD9dq7lGz3u35HrkWB95qguLicGz61dmOyz+
r6QkQy2gE3aJYQSeI9EjtaibYJHKJYmLwrsbGYQlIEAgCb3z0JBmG+wVDfgoMwK8
LP4EmTvnewsLIfIEM/JsHnM5CXRaAztljIh9D0tDoLVEnMu3brxQOApYEN203a09
Nidz6k2t7mdb2SsC5VnvcpiLqxNgrWR4lYjbOCj5V8+TrtQUq2THTvu4u4Tq8Kco
`protect END_PROTECTED
