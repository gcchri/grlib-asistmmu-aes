`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yi/LHgrYvN1kWTY5OZrIOjcQTc/PZHxrHAtwbY9f+C5h/Au1/ybAqV2aTugOfWI+
qgRZPgBQWOB1/IjufT+foN44+7Nc73enF7gRW3zeIb0Mil/RLUn0AAJ/9mq5RQCy
dqgLhHkaUAfaPkPRPo7+6wQJCdYJRp/o2DBiQCJqRR3zgY4I2Gd6lxC3bOfyOFxE
ER7l/4C7M12WSLjDzTioKWmuvFPzKK4q9kEKtyvwJA+GdguYjnowexCmDMZ9cAV+
sFKLWpdzlEF0e41IHtICzB/XwiG7EgNfOvmdPu/vEFEZYYmzbnZPSzy2O4hiJ8Bh
nCzJV9HF5P0q3pvYddVkye9b/T0m1sWRVbUm8Thpu9LUwXPqrNG6m6BRPlU8/A6I
Gv2WarqN2tpZPjOnpUWeCd8DoX1XtNkfrwoaAW+OGxuDDwHbK+zSp4dmJCz16YJZ
pB1hxO9Ac1f6TdC/TZrLk/ZXtoAlSDy/STn8gI34xKt5bmSvUaRfNqOcxGCLku4E
LwSkQ39F7a2wPItA6q4Vsaf71/Uyc//B0OMtASWZQcfqXYO/7uR5+snWGs14pe1C
6JsCY4SOV5ROEbxfRgsoJY3ZCUmoWZmsj8Zkh58lsmdD/piqgDZtn1F/FJXQc42v
yFiNCYentXJogm17WAoVif0RomnNY0mj7dzc3bPMME8=
`protect END_PROTECTED
