`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9PPJpeFVSXuIhbCfFn9EgK4T78ErHg2oB+dyIjiJrzMAMZQvtMeYIQcVBHPRpM+9
uIXlONhFD6DnNFe6qVTxylPzSmFFEO/a9/AQYHIt6C/mXFK3diwMJy7WzeBfDQNR
i1ybZhIwHgAv+18RBy2Fw5ShlAYSZ7/xkZgWoNNQQKKIkAPgEhKDPCXz20C1dGbd
HFt0pj/xy8Yiuc7GcBdVXgvn5VMOaxkcknSlhDE8b47ajS19QSmr7Mmarw/g8/NM
KeerEkksyGuxrg3IlV3EdwVEohof2hNzqSr8nkUBIb0TKDx/r2kH7+bP2y3sZLV3
mbPXj6zMLglpdPBfYho8+0NR+KADkkX4krS++uI7oojWP7zwLgUu8mpVLX3L20B8
oINJ5hoxd8zhSfoHFzTTClUn0Xw1uNaMT2cYI99etmcRA4TJvkxvTYlEpiGI1eUj
LlpAO3p+30N00OLpLCjv9YoSRImdVEv9RVSFxUm25JoeoWY92FTujS7KYhWqclnP
g88KutKSam7fXAw/EcNRc1b2pxU+dk0lrBq1kRyF2v24DenpOiq3NIJqAojZMQdK
lsbUBgkcH4dr9izgLLS4z7VT4yOigTWbIuXn2V/qEL8KRuoDTH5EEOKm07Ei1C+B
RfKJ7Toyd1Mp9JC2Dz6DA+X6Y89VNjzWDzfsoz6wmtXrjCpmkdc5/Vzzj84AN8fJ
dpMvQGUcelzM7EbptQeJz27EiKkkJPxdrl2wJYFotyehQ1Hf62MCVeU02RsdZN82
84aTLXwp8+PXwEbxvcTmM/owXRW8qVX1B66QgbM1oSIoUY6ujPGY89gHspdMnt/B
skqAUOzf9unyYeSsrXg7LzjJwMyNGlbmFg8k7P6dk8GqDJC8h6dnOXiN1eTzXcfn
NYZNvore9Bkr9gCl17mV1TRGFFtcj7vbbdQ3BmjAJz8D0zSd+Zo/ItO/+eRIFSdq
0avOATezSaWiS82dKxNAsdPpb9+uG2z/vYFacMvZbKHUTGEm8sp1ipWtG/Q3oOoY
wDy4X1p4Gg+Gwf5PQW+eVrJL/lUG4yuQsxwRwAxmPg6nSNUpfK31WbEu/IEirxOT
lcBd8Bbm64Rila9iKWyTAZdjQIRY5kDbOZ5874ZSg9lWa7qvqEBWLIeHa8w6zU2G
88D2XANJuIrH6k0apAAxQ2WvDmvpqJom+ntpXuTowyaw/7Qph2gow2v3VT97HZ2N
bn+cDeZY8pJCvNE4VLkvVzgs7cfm6dhapHqN0j5IMfUwK13tfJ5Q7wFMdk/l9Xw4
JdWAg5RdxCnRT3KLrx4Ayay+7Wqn4odaINipY7UshghXEuOQyq2Rl+GMgKuKZONe
oXPvNCCrM1Ojtz54sARPQQLG6WVRjt8HCDaJHP+VppWmO/cpTLEudoACjcMhzJO2
Ze3zf5w4Bs0C8cneFqcSm0V2hCxMhQbsMxaALfBOppJFGrWnDKzlSk0jjAGLSm32
L55PXqHemDLRNHA5NP9pPtHcSWRTVgirJ/uaM1RTPNsAKf0IRwp0VktPmTmBGzG7
gDAY/Z3O+7+CaRH6XGRG/o3ql6rqJ8P9iuHy+x7s437AQLkNCDlndXzEzbyl00bf
zgaWhN+X0mKcooDCfgid9//kPuYBIGwkzSUQOGJtbzX9Sr1gm8uEP0/QmDtmTu/9
DV9ZoLbp+tMdAhbkcdIZY6HlVb5EdlLuxB9j5T1ac0TV69YoLAU8SE928tekDhGf
xGkt059hmQ648r0yB72S+/Px5az6/lCQGFg7RA9IHhtn2aI8IgihL2pyJFTqmiuE
O0WH/T83rlr7zZXKzzTuneMDwARGEk5+ekifsqmXvlI9vqYoZbB+PgI3hlLYqRcU
ChfGs+cWvxTnzBvkJA4gBlW8dAZRaHEmAzH686RbC9mTORlM33mKnWQ6IArf2A/7
ffdUPFzlhlpyG9VeOyp8pMtfH6h2KYrQAxfAIHgwykFUh8c6pFSHdIlOGq2rDHjf
letoFsV4kDlY+qdX8jbeO8Eg2wz3aDlIszDsTQc61B503M65qs3kqeCsjC4TOg2A
kKg6Q/EHAAhFITi6o6bcs7cWV2rQG5mEz+Ru6KVuDyiVZyTVs4TsWvyEkLpoQnMu
XdJ6ontuMIRAo/zEMPlPUty3MkZ3ghe7A7kftAYCVHKWqgO0uSrbjPQPGZkfGDtg
5zJX6wz/cF51LRZA0hYnESuRWslVVO56AW2xS7ysIdMHA1CS9uXTa0S+YBabcZWq
p1O/gK5Nhjn3jSr59j66PWYuV34zrYQjDguYqW26RdM7HaWYnDazXSaqFwwaTkEH
/iepfkt6OXZnQNqShPZy9ED4iGOiADqm9j6GtKwRPm3XDIi4bb7yIIJVpmbnQZQe
MK8x73WjQAZrhl1kvBDHRtqrA519lfVoaYLPLYkjc9fnPohUrp841G3tvUhCjrqg
PD1qG2nlen3Nn5rXY6i39PjGAB7AI2/2ctZ1uwUWJz49bAntSgMNLXmw8Z9HVgNX
/FDrtuDiXk//JeZCmIiWv4FLhMZivhISJLMKxp6QhjRrZlzPUZLR1wJzclPSBRwp
464CspBuTi6YBEkhKwywT5eDskNWHKLP0CQWw29rFFv37l3R+DZrZzIgi55iKKJy
HwRBcPvWt1YkdUDuk7pHbKA6Hh0r/4KeaNBd1oANCq2T7dskhZHgq3ndnCPfXqui
C6/EvBE7xB+fp3k/c9ZL4D22+84ZFtRpZpe2T1guV5TsIX1SBGK/aK4JkJ8rH3Fm
4csK0twSS16ScOYgoHvwH3bUmdOkeLuSW2/OIITkz7xm2DTkx9viQQQgeGDM9G7K
duFbbgoxBZNFLu/I5yA0QBOO7kkZH2+NpaywZpsZH03wWLltyghW2sw/rgEvDCko
ZxGJd5RtWeiFJKmh6ItnTP1fCmvo1ceLi3vzqcVkWTDpMHbtJlidYbRc9lYmtyoz
nSLNFHUPwLPu9YQnkAzgz6p8w/iyw891LFQzYXmlgT3ymWU0B+enCl4eXn+vWJg+
YH7izu+aEeSwk1Z9KCT1YtuNPlX9CaO8GLneTlN51K5bBh7pVlbxG7aXjVh2TOwB
j2X9TJ0x6nfP1TWOTE2dHQ==
`protect END_PROTECTED
