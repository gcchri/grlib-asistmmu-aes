`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
chcVk0uES8jUTJE3pokYRyHsdMyy3Dy8wr2/URtTc0Tc3HQoM2vsvvvE15Bp+ntQ
JgEmvyOW3g/adce+jbCGj3vJN6iUtPU6HtOFSoc/BS0gD7+nAQn5zINaUuXZzKN3
tSgOymnQgox/sBQU81zVRp9YlPz//THTbQcC5MVqtD7bcR9G5Qy4o796b7qDc0uS
QSHMXPXyUVxKQeO5GIIjXHZncsDPfS3PtQd/0i5WUQXdQb9OW4/hHD6dDn6EaAXg
98BS1pQpsRslSZ0qUntoEx/tunkgRQ1kxBO29z3iRkewRaGTSSc4v8BrYpw71fsJ
CbJKwcfxWXIK7aZHPZ9XxYN6CKMlG442W367jDoPa7tzyTOgYNM+VvO7uMvC3mcC
TwdQvmMAzq4iYttIqN2zMnWXhHd1d7usx0RaOVxUuHhQj+h1+FvQMmsT6a9h1kMt
BAy+dIUKSKguFQF/TzkLwX42TnklWlt1OtMsQ4FHY/9ykFi8aed2+HXuyNzkRW2n
kK/siCYyMOh3mUFdxbb9caFW4PZymYeHuI6S2kybQFGSIQN7gFGB9uwYxJhiVbDC
03RqgCCP9UQH5akYn1s8YgecsUi4/+0Hv/ueQmZg8uiq0mtZCeomFZkTpddnEQE3
olyAm+ACjkfkc4VTGMFeP0oeWKaxfso6HF2fHVLHIFeUsr3y3Z50obf7LgMgD7dL
OIjHc/9khNLhRK7a1MhPlJZCon4Kodz1UE5XrslF45ANffsRqGmwU3rlL1cechOR
mo6zrLyd55P3jPuZOIyRxoppMd9Xn/89RpUL7p6Z/9rX7icgVWDiDkevsP9KZBQF
Mzb5oD27PL3POfsbG69fQc3hHwb1Wl5FNAZe/7eQhjKSavB45BTk/6o75XZ4CI2S
kGNgEVBWmNBGqfZCLqz0bp7PZznYP/VFCb5fU+w+5KiLXBxCLyJJx91COM0xEroE
4LFKKztcVJY0pm44y1iETHIpyYnQGDGy4BkCBHByTVO2Mk6/arnZd1aRtp7FWUN7
rCJJrEUipy6KV+Ma/1Hmg0MVvxQmiOFv//j61gYCiShtn7KP1wSbIegxgW2B7NS7
/cXtmgiedYk05VkR20LYkd91dQ2QBtYrZUKwsVKbZZpK2XRs1n2OpD2xoe7wW/Ps
f2MI3r/7myG9zrgIsJ7Ms+qt4EcNV3vpMA9y2Zt4QZSi7WZJXGGgCuGgbkYy70ss
dc3L+3+CLp/I2HB7On88gmA6PSqz/t1jwDp8xClv/+wdug7q2EklABWbps+O2V9s
BGM+8yZziKwwsgbRRuFqZq8RvR8K/clVZHcqrR3kYx8im8opopjx69f57BjYoFd9
zOYV7iRKF0i0rTyabQsxj9WefGiSoRY4EEH+6V1DvCl01uLZ8MDxXUk3Mp/dUucb
wN7dxSBh52B/Y1AXT8qigQZ230KxpJfJ6uNVaTDR0ffjSJtR6JIxbFFTAQ3un827
co6o4MB+4ivO/CUEM95ilkMDqPlZjPQKedW+YnWAaNd98oWLYT6V+9W3MrQO5/hM
`protect END_PROTECTED
