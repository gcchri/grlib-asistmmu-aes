`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q1SLjGB7OInZqTiGkNMkMXCfn6lYYvUTFzntlHJWUwmBdnH7SONX4v0Atb4oaAPb
IUkq0j/c1+3+3yCXc2oZzCr7IMRiYEBKV1ut0wr31izo9Tkyf+64o2156cnJ0IBA
zGHB2w/L0xfnouDEEi6fm5spKk0niveRMaWD9FPDUnPng8+ASn7/mnmhI1nUMsnd
dMLM0RnwDGIaIPgX/S59HlIJu6PhRKOq4lGLCpAGsWxtu/QlI++TcMdOpaMOPgo3
Pnor0Uw0VABw8X1da3Pi/nemL8iVrxi2SEZxRVJ+qSSnL/BGrmWb0lQby1xM2OuS
1qhDuP7FMiD3dx6Rs0uIvLAq5SEbj3jj+c/YUr63ndFmqrD/6u/cLmxDK2/1Zsnv
H9kfFikyZ9y8/Y6ZqjzflmdBcuaiXU0tEav1XJ0I4NymmRdzy0ZRK5gfy6TW891b
Vh6rcNJQxXOfvKZ8z8zFSC0vRmErr9BJYpr1GD3CYXZp6FnUcURRoixsiIRzqXL7
bmgUy61Wx2M3n3cJVzNtlDVpTf9mNxCIZjOvRuX4SvLwECrF4JQDJPLxxp1Cyiyo
+1aWZvCBj79QtyXwbKmhSikSZ6RE31JSqUjAR/dztxd6uLcoNG5FgWVPCulWVLPG
tr2dsVAeIKD0+/YYSuDIBMnVmv/sL1QxRIbMrM9wKKp98gdimjT/SYaCww73BwGh
ycTJWgPu5lhpcBZ0RX4tp+MjXSLwHPY6d6FqGvW/XwV9lYoZIBulbPpzVt6ZdwN1
Izsu+cfCQbpcAvpqVaYt2PJo2wAo9c0+0lS+rG0tYldnQZkZ7K+6c2KEzl/AZveI
IEsdwPqa2ykFGshi8SH4omHAMHZhIVt0JvKfVlvQyeh3D1Z1Di/A2DiOyZyPc/2X
wA3w35lAMMNwhTln27TKk2l8gvIzJixmQO/NVUE4AdvEJwT9smVagIzjvUf8nTHR
XJRn6ewO1yejXZ/mcbONR/y8lXFdlcqLu3HjBL3KBlQ8E9Y5wo/4/dIzDzWQMdgA
8EFsNmYdMNi16+5xaLnukHBKjwh4I3FvXRpBOiDGkB1j7dB1w5agVH2YIioVz/PT
KFV14WzMb5djO8J2S5wJ1o0Kyxljk1goJdTNq36xJdvJccaVPcHh0X9e69exF8TG
Sdr1QCuS8eXTBxN84chu5AqZt5951HxG64DyqlqeCcRnN70a1JilGJhdbHltNkoa
W5yzyc6XdtVevqXyjuwkzSXrjAYPCNyn8ro3R2ZWc05O/bEGGOvVx4818M9dPkNO
QNksTQnzXA83LNqVxrsVFLNP1Pn0dvEeCQfoyb9I697AgFpsWyp3TyOz+jIi6Rpd
5QBqUuLeeNKxohHII3p8I+zezf0Bxdpq5i2s2T7mQWoE8ic5UiSjzyJMUk7ek0Vr
oosImyXo/+zdFeKG6mnEaKBV9M7aQTrN5dpOXYfr16lKXyuXuSRMGLvkLTrIlGZ0
`protect END_PROTECTED
