`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wQMShXGjZJqZGmPzeKCe7q5ZJIAXaDOA8wPiHa0PHCU2wf0ubEp8lPQqjP9qCtAM
DefwcDCxBy+Vzsv+3ikFJGC43jPMYN03/6hcX8NgWnWbmKrj+tL2KMY7bY6svmYL
XGBt0pM8VlXJy2LB9OCCSMQ483eAK4EGTfQBOsjBF1y52irVuvS4dUjEA72m8JSO
qfJYw9NKwy4EWZ7booc6KwR+3vh3G9BIl8OjSvO3E90CgHETI08zRZNuuCFgQl7t
gaZC+5eemd1ykZE8ismzj+L52aD2QrTTYE6gX5j6cLg=
`protect END_PROTECTED
