`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cDyaeE1hwY27pGg0hunlUuMWHLI9Hq8yTdUWLahbtw0OyBIRGDQz0WGgkVmgJbpW
F0TRKqDF2aqPsxIuoAwdaQl99rJuTLVVlaKkYDE30NraydkospYtoDKYeRnnLxmE
ZHoZGmpB8XEFAxvZefA46V0ZHVqhbTmMkFIatc90kZcvGSXWfkjPFFfNgRRkvajn
FKV9wZZDwQiGDb6GmEO6S/2d/sHhSuwhNlDYX9REBlejSUEdJwoRPg3LK77dyDD2
Q0SxSij5QhfXCgcYYES1YSfLcknoxa+ylGJjP0yF1MbaNm4j6ae/Y3ddibO2XRl6
2tua8v382g50ejppZ0vByeWJJzuh1HwdzAPK9CkLYq8jDCm7cKR2teOm2lMawH1A
CKfQATVDCUK1zVDAJYzndcUNYGqa2nvbP1BQJ1eCs7ojP8jfOu8ALbr6P8uuzYM/
yHkAPR/T1yIg5wRIzsgpgnjEXNoU8UdFzFvFmtIf0mQwQn49BVLPQGyFe9NtJmAg
`protect END_PROTECTED
