`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0weL7Xxy4gXa1AF/nAgJ8MjKs21t61yF/LojCb9AgmRHpDjipxLhO4G+kPKQ6bF4
QQaN0Hz7Sl9P4s2/DfVLgJZAmb208ZpOHqIg68Akv8AU6QYCcUj6wqP7VuNKbgVj
1wyJSsKGqn0rFALbWzn3rOpLAXToVsFblFtdtg44zCs6BsjCPHuTwmYIVZWVcS6A
74mV1sH0ldc1Zy+/JroJhpgFPzNoLgyr5VXsQy4hERJBXyMUmFlpV/vE/GysteKQ
0qNd+VsUPxhBbakfeS49ZSt8qRr0EILXLn7kiDNcGminqf7XHoh/56c7tpndzFu8
wgsFDcOfW+4z9Jkztk99dgU3SLeAgb3y+1fu8XE+EsIb+NCYwoku2QV13bRZ7+Kp
ubchleEyWhdYHfhRsZiqN7K14zsZeTVuat0DCrNkHGs=
`protect END_PROTECTED
