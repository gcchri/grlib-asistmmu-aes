`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UlUg5eGz9/tYd0mIFl6BwsiJ9tm2T/ZCNye5bNF1gX5Q2x9Iw9bG2MpRN2DNByLk
1OMaps3kdnIpHtyTwYI6ohsmylC663j69G6XNSd8HgRoZTuE9ys0mI3zzOA6BaWh
/j+leXkJWATf3svniqEMbjqH8CrCaa0bwJspHMnudRs7xAxLxy1M+a5CJqb5Bnrl
GQpnoEiqXxFHtzd0tnepluYBcsejEpeLx79mFA6+E+1pQAKesvSO2F7x+JQPelMh
XrD+ObIJUctBbSgqlQD0hnJ3YXy7OUUlyZSbPncTcEWd+lWKJFVtClNDh59Jf+w7
BDP/iznzCKW3wtkW/x0WiButMrieUBayg+t4R0HqXOEDxihI5pPetrbOaPt6ndHC
dneeMFq4fcA/96ZgLI83nRZzHRFIZP3vzEGrLcy81YE6xJqmmEaKx+bVbn2fhkqP
vIKqDYZpnrMSySiKshIB+/vABDKg9ZOP8oYEd4i3qPgyP07KMSJ/F3t46INU0jlW
1v04VJxYM80H6eR/m4yaWA==
`protect END_PROTECTED
