`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ef213IFUydCgCAy3UxrafWbLEZHqOT4sm3haHEerqaaEB3aGPtYkY93KaQU6BRuL
LtD6zqj2nYNk/+Yku9Br/Eaz+UoHZoDy9bazaAB94TLqaXvKktuRCj9QnrFo1nBi
qIF8mebMccI5WYg75jKraNtvOtQXGRNyeS4+pWlyXzsvHr0MXNHYahqLlxyWgwyB
7S98Y4Tfaql7obVwV3a0/Uq2O80sUwkuM6jd38UAhBUkDvlISsp6glzqGK01j6Uv
0pw786OBkqvSLzHdKFHfk0GfP0c3vsGN66P5XtkD/xCrwoYoxA04XzKWZ/ckE6pO
ZpSAAnxd8xU9lo92Tfiv8w==
`protect END_PROTECTED
