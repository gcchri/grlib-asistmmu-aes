`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3zX5/zrv7HWPD913IMoB6PnBXywHKgBAj9XcRmsEHQkpgKhSZck/tWtEj94foc/E
GfN1s/c2FRtLiME65ke+v/MtIxp58Y2ezDx6rbLp1roQM56IpLu0NZagMYvgEPbx
7HcHvrQQt8XAwLuLt+KOXLKyZRzTn3HSxZy2+7R9WR+woCP26OB+UV0HpXs0UYKu
l0XHgTRY8uc47yt1D1yCaGirN45pKGx+e+QFLzfDQde+Xo/Pq5i79u0LDC2qFfzr
nPFQulmFpNis100MfrYxlpE8JvGquQ73eyVdNaIxoSucGidJbLsU/BPuduCrMAQo
r7eh/VGPVKk1tF88YDqd8mHUN3aKB+pZFhJZ6X9q6hYQ9wZBKJ0EqZ9QeNiGXndn
LCJzv3FfVX6mU/z6Zy+NN9V2SnivaxmlkG0ex3gAj7fjwAZuAIRlAxBXxed0IA2I
f7ga6JRb5w5Cr7Nt9c6u1Ulps6uXbS8md7bLd+qT2iSGzjeYbF42z5XlRc77IBrq
91R6KgTS8rTy+TkzZdPv94CFOYfMPl7qnvuzfwwb40zUyM20LW7pFkQ3IEJPTGbi
7/ri30cOaxXlNWUETVraZ/DN65RQ3ReKhGgzUjk6m/mzTiQwYmiojfX4CLk3gQxS
dUnUDvt2AqgrClovN9wEuNZPwq3zjLUMpjS0gvKuGnbTLwFOLARrxncZ5/nmMcwT
bTxXZXyjdbI0Q8TDJY00KqdIw7rlYb+s4XXWs/efF2yHExc93mrfNdX3VAxZEaTi
P/KaHNBwz944+buWGr811tT3Oda/YoXhOYW8Q5Ixu1RhnTdQSMZGOsvtDFLeZkk+
JnPJHVJxeanYZQSyW3KCWb3nMlI9Li1Cxw5cuTQHN0brLCUpI82c7BTuv3hXSG4Y
9N/d9KGEMmn3qZFEDHCoL08Bk3fAiciuPDOeV/8TaHo=
`protect END_PROTECTED
