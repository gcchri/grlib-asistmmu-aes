`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X7U97pXJdglJZPHAfB+By6on3zZ4GY7tO3mmkIo0aC2tqG9cpReTJGhs1ZQMBnl3
92Qf2TCLF27RKtSZOpYFygZORIsfVHUOdxvMTvu7wg7UKcPg2x0k9AJuLpba/KE9
kcdiTJAakaUj52ZrxLlOYjt5TMa52Q5jKHx2l+/5I1/4qNEZCyFKLV3TG7N6RNHI
orxlYde8hk/K9wSLLDGUIl/3p+wmE9oOiinP4/NUrzZlmpwEgd2vmPuFOvkBNAzM
+F4ovc1diahejb3BRGtU8mJHsRQKOR8AfK14xLBOawwwpsGrtSIeAASDuVGrGkpp
oyM0gsJ2T2rpp+pwhlN4R2kyHTCpbAp9c70c9sk+WgWGQEnU2jyPI1sqQo7ZAt7A
HyghkymXZq9L2OGHpNZA4F0GFkOzlw+hM6KTRlWgCtpguy1/tCqr0jKJIdJYZRDx
3Egip0rsVxiPhMu+9To/LdMbheC7NEYjRj1vNc9mtErxnGVr8lC2BQgu+UGllPzM
btXByqMADxjE2FOwfkSxq1BcxE30scYShNUYUtizaoUqWe9RMsmAbnSs6MkhBSPW
KHym2OnsqFJCWqZcq+21PQ==
`protect END_PROTECTED
