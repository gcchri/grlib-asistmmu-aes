`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j35bpLADtB3nJOpE9UYXdm/sBZysYDB4UhEeD7AW0sJap0Gj0k1WkrsqYhoUS9we
GcSZQxGiag1j8Zn2hp09D7zzjRVomKxY24QJdxHU8RIUr9wxx2izSYOZZmUZDl2m
i1FpNzdi1nIunv2/mQxie/ZkRkbF9u765zMvvr0oNgV/yeHiraUuclSimjc/n2he
6ScE7C0Ey1yxvGQw/NJWglPvPJ8+I2f+gpqnSvZLnevrBK5oJCDwpZ+GrzyrsSF7
8nERdQoyj+cOW3LUUW6Tec3jHc1rMhbzfJmv3TqEQFsmOvomgvOoZTwljQM3yN93
aX6xIgIdPx7EYJ8lMVcDNw==
`protect END_PROTECTED
