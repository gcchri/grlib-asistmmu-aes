`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dMo27CYrhKq4O1ubNznPvPdQ5YbBZruF9QHkXJYhyxn6U5VQf3ZJg/qZCA4VhuLn
AVMKKFVqRVE8nIJ0LspSB9JJMTz8/RGGs8ZZa8ne1L0wHOGaODiFOomv6IOV+dxb
WNTE+CvqYkm7LGWHBYSrPPwMVr5JY4e76C94mx61DWXFJYsZE0ROnm6yW/aWxLfm
o27CTOOVRMXNQTjUnoIM2SpfiKJKq0ETdPNSpF1S4ddZkZjCFOo6QjxeiuvK/JHZ
6p227F0uCZiIdUaH6tpWhJUYm1omNgYGUXCJq7qaUq5NKvOZfUVp09syCDs3JD5X
yujFq/gO28YZC3B26VXOiIMUlLg43Vs+gzx68BpjQP2cBlCf1wvn/AdxUQlEWpG9
ugDr1k3c/Pa8nOtZ56DQZU6r47i2ltOVwGhd1UK3vsQE2nK35AbeU4B8TUTagRR5
kYtDq8bO12J4g0bbALLie/ennyv9eHksKVii5jBpyAfo6awgU7O5ZekFwaFw2RaW
Qk4HooskueMkQWfzsX9caKJ9y86FNMobGieka7GflB0tNc7EOk1lh+lMGrT12UUr
vuHh3NclVO4fmI5Vw0B8CXwGaCgZeZ3rhKKbpnuoX4czMUWsrYb5eA71EdqFlSC9
WZJU55EjnoFhFYD69Nz+J3xTAfx/aPa5nJioTW6PNvzQSXRXIvfsnfJww6C7OHtP
kaDeh8gkslJpFc/hMmTqnL8jZpsckiqzzQv0WEDdmz8GyF0yVg2oNZX9evddwfRb
JJbaH7CXRwPWNsfHX7ZMM+p/gSYEn1RS4dOzpzq3Z8yi2NM9v7n1XXh7uMfpAz6f
lV5uqyAP8SP3z2tI/Y0UoPTo3llxeB4099Lc9ZpldKvn0x/rEWK1QgPLo5fhqdub
AY5wJsuVAcwdKHNCPeeL37GYB6UzZBhCA517gv94YR7usgiiHPGHawdP2YgyCzSf
9fzB9ZVJfMM9NyRZpGCDe9tg7zlblRyHV7ugzW92RDqRQ0J4Uegi0uQQ/Zku8tDq
7jQDMWQ+M6cNNfX43ZBTG16ShT2m+gr8IX0oNIo3QGRM+TCFqPkQw4lBLBcZfVpC
sws/SKi7O+sXJtmRNqid/pEci7iejxXK+FQYzzZnbUZLWcjyUefe5zOkiYl3fVQE
yHCDgMMarxKNjapDEApWu56cgmbJUKpne9XHdgDJtGr+S790qm9q41HlwHlmW0xd
WYSMl3JGfbITdWW8+cv3gtA1V5PMlwFoUAlP1fJwGOaAJ94I/Ev+2JQLt/wTxNXu
QwVLzqtNeCTG7jjHUI0/zh+aOcJ+vNMRfzLICLNLoG5cFXs1RyOtfJ5idwknaBfV
TZut7GxNXVvvSnypCbnOnB23yJTeWm/vm81/R6VIXvPp0Jxjo1iy2S1cTaYQPnx0
ahLhKu66etw696hvIFztWeuOen4Ze7tm4QYNF+bXUEJOElqHC8jiGzdEyFwx93ZM
Avy1tDGSsFNfDGYX/dqMbYgRT3r9Ty0N16l0SPodv+3ObtmSUqhWDdLsDiiD2CP6
ggxc8apb2LH0Lr/Ozdn9ksTpfWVLowT5DaQBeJPVi42iBEL95+pL3EVwCJut91VS
81mJWoqnsWP1G84mzCLD8FwofHXhXQj54taI51VEN7qb/ALxM3Tau/HQ4lOfDajl
pNdMCMqdXIcBAlvDHaAW6bZvvq+w+Tf/rt+kOMq7TceIWTq2+VDcxXpnFmxQDiNj
mUgCAM3zHyLSGaZ0X/Sqz5pkGwH7rzblPu1h3Rv30E+oR41CVKnJPSpMg0N8uuzO
4dx/jrhQgxpY7Sc2qNotcuMdiE1LYGND+C5qdMt8u6HRKQ0dyRDcPScm7SOvf0cb
A/giuglGcqt7AbL7WNyMLqoSUMr5+Qcz1nmki35TC/ZOA9hJg5HJXfnctnHX4+jB
YtYWeVTMITVP6tDlapKqeKGPsgnGINhZTX5HF9YsxmofH/tmug8JHddLj25AoC6n
h6I1hH6JSxHO1F7k7SJcwNzGYYQXKd5gwUOjGay0eQrZTMZfVsUGRlhfC7TT4rT2
iikhTcj9y7mDVYGGHYpVmoOqSg21YKqvUYYaz9Kbw2aKKopfeup+/Pjfwi11GzBJ
p7DJmPGvUBwLHKPFSpgqPtl+gmO7tip8l74XXZXfHw9FIzVibVOCN2yAt4dezw1f
wFHrIiIwZwH2IHbL8qrm3jfQBsBuEfghXfpxdo88xeRLX/1Ivpam8Ri98fDTmK5O
DAYfe+c13rYIDGEZAlE63LM75T03+LEBuiIoT2lu1ItADTmaHoH2v79Y1mjTPT98
Mdyvz543DcxqbADjceRkiuwv6dJa3DVoEL1is7Js0nagGF8y3w1ibMwLL1ggYbuv
BenZC9P6LHOrQnc2TKoBfi8kbM8RLx2Q4B0eMSnG2aK3sTojxFOZFdbL0h2j5vrY
ynJg7eheWO+OiCWZ5LvF1vrOalVZmO+DBss8JN43CSAuPLncnu5KqP1U0ykQeWiC
+RM5uKdaIHFL7daiksS+tzlg1WCmTiP92wJG4qRVch+/T7jV4JKTSef/PFRxyFtF
hIuOm0YnAQE3YmAb2pHicQCd180uVBIPyG8UAMq/xcy1Tk78ulFhE1xEqhtahz9g
blGIJQwMM472cGlaM0gQEexGeLD7q3xm7miB7tYI49Ewh86Bw4PXwoFnv769RwYA
a8hxsXd/lGT5X+gyO5SCZ+Vg/dXGBmS5k19kVWWzkgdyq5Ne5kwCUPH47qSxGJDK
wNL3Eys1bA2gtFi7GHl1W+VoEWS9+ZtbcaLinpfGuj2pvIUxJGNrS6LmrKQeQelS
CIPi/v4EB1wMZ4W+3v2aS1l/HgweCF8kHc+hfhNSwH/xvT7Mas13xhnHmS8lNkQI
uca89H+ia/3Iie/0pvd5/i9rpe414WNizQu4F2JAxCsC9+tVWFsPVEkSqKXZPMzo
AOu+kTOkFDvOs5pEvfzKF8aBSg2ui8yJvtED0wIhSOvJUAHqt9WupOCkpyiaPE/J
OTg67rrKcfOj7TwSU1hNn4ey5mFFjpNlSZid65fdFqnIXOHeHppKmPlC48E4Rmge
+XJx1DEUyFyZ6MRiXmKltOdrdx4EO90FB407ph1XjxPiyeIRjHQPXunykstqLH0S
vCOJe24PsB5tYp2jA762pMC8Tf4BkL7tKGoGruVEnngVlcze9cMTya2FJiTYu8Cz
18LZ16JGyUEmgvRZjrg/OOEGd8CwU1aNMDIGfsWLDxDe0Y2MAQ1KZvGzUN0Z46bD
lKgzfkqlh35mZLf+C+NwfHXcEX3SajeOzt6h29JkQE/D6JVydbs6YObKklXGSV8g
VkmuRiJG/tDu62RR/okmp50v66TB75oUzlb/Z9CATuJ0Zen8WOcBg5jeLyn2h3pL
SK1WzoZUgh/co6BFMwWeSQgd0igMz2dqOW00T9omdhMGRg5zgZoezF46tQpWQIiL
hvK37BkTbl1F9FSZh+Bo4drX5/aovmmXNEUWh5z0p55Xcan5ZERthfaj3rdOccYK
ljfs7+QhJIfN/Q9lNnu+VDwij/jYYYGSvXDAKPVm4XhBfryBC8Wgvj1dk1fsPuvM
EoS1noGfEvrbgEF583ERYg==
`protect END_PROTECTED
