`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HjCeQwmHyxwmp0ypZvPRnLNZO806Qg+RqPWWYtnYjG/2KNbiHCcsQB6Qt7tmvawT
TkVntk7Mz0cfCtLmDntUXIvvX6xIgVf0k9Xl7Dz9ajt/axJLzcHcJTqok9zEF3q8
JiyPAqxMjL92SNIUzkdqSLqXOvp3x8jEbBD+eN/EPsZRn5VicS5ICXFa3yL9tles
wHT+/4qa8wqkk2KSkHAE0aU1rHlsdz91VQG3Quclwj7IqqflchfgWPy+AfTpLRet
5E0o8LNRrRC+Wiukebr7r2G+x8/fTn3ojfp05Y8/aIpwVGU8xQxRnmSoI9XzUasI
dXiAOH0SFayHhxLbYjE+QDgAJeAZne7ftq62Se1kQuhJSTcAVC5ZwD7V5RK0bAYN
uStTu+y7kzCSWB/7UkkKOhZVtTG5LZW/B5bH8L1tx3iMqsCTbeg88Xss3JWdoMPC
56vClN31w5h/CidaFfXjwhBtuelt4atXTd5wV34LvU2c77tI7CH6pQEb4cCuogEO
n1YKocZLhhqfJgAgdlQ2Z+5YW1BUrqyBdP2xBfpXFE6zHkJrDwNIUKB7eR/mDv6D
W+rU71FKGdvQTnUboeQX6cg5krhrnD+Fupt/2mHLgoIaCyxha+vTP4DfPiQEi4h4
mCAqXo9kFjXbYIFS+SKkgaX9TKPbe5h4MYn6OITozUPhJx1FtEJi73F+kOR4WHdz
505BcDnubuPDsGcKDGNvT2dlW/uLv4tVKUWNbPmKRimWjVlNUAF8rHYzGewBMUwf
7ggYh1o4VcZZgKuq6IHbUQobaEWSIpmuFYOcpq0eg1aNOebtsy+sFu+hOduhpEkC
jtCpTeVks+Y2Rrh1sUVYCWBUComzcnR2sLYMFdYzaNh+MtfgwrgDuWBaUf8zY7Z3
p+xx7YVFl/KNYhMx9074F/f1rlSy/wxn9m9faBiV6DoU3ae8AQM3EBSg/1ZqBZ6H
Su+1sRU8P8hyB+sw6BpXXEjDf5vvgYBIZQ6VUo6eONScNbhSqAMP+Gsc9ZCbml1h
U99uYjsT2NOrLBGXx6LiBqxsoGAnuFZwNg7i7HMrFBakmkesZM2vkK8fdgtVyK7E
Xks/maXYJrQ82RJysTYtSc5F+ZWy0oDJ2Dl+1zvLgRh3ioKrybSuf1jk0dwsxFTE
kzXmr1AbYiBCuX6o5DRjZXDF+4bo1matwR435fQNqMrnM8kaBOsJkk9yrqjR1Xi6
8RFMdvUWasbVXaRyorxHDMEoTvPJTKaZCYUm/wK60WanzXz06eJo908fRnpVyhRS
xgAbYID3JuI1qOw+RtxKDQ6rB+CiqEe89h/nEJHRW7ATzGD69TC3IMCmlUW1U7YM
vPHPrRlgRcMXMeI9Y/ELPqZ36jn16yBfAwu2GmOHyQ/TN+y/yOQgFw5/rev9hwhv
JjqMkkpoed63mSrhA+dcaw==
`protect END_PROTECTED
