`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aq1yl5dol/NEfh63hc18DOpaGCgaxlm+zXqCHt+QKKE6XEDpq538zH5D12jE53+s
C0pNFT2iE2WcPifgC9eDEjltMBeDvTMueI+30QZsMOSP1GFdjta3aI+7Wu+45GIC
a5R/v27CCr6k9qleErqWnweAw1IxbbgG5cACLklUQEr+ywZPZoi16km6r3e3mW6r
73blsC1GvQjeOFd0Of74XM2v/IVuLd9b5orEZMdmYJn423351vkfl4oW9c2zDNh/
Jl8fDdTNUGy6WKGL8fBjF3wlsOrFF+h/B0YrEIpUjtduUObN6hzLq0qoi23NHZuI
bgLqFnJDnXcRtAoavehCQT5NFPThV1jKnHadpM0Zq+la1yqxjkLVCK08uw6yLiFP
WexS+5RZYEvku+tdlY7rQdzRJlVx/a2bqV//JpqCcFhGnO5qb7JfTKK78QYtenc0
s28thL1PW8UFCbw8ioKT16hv0Ix1NCcChI1oyXGcLImdn2hPHg0q5LbZlRGpA1w/
nkMOuDuYWQqE+n26zvTOI8haAL23tl8FoEcs9uMOqWLvEcoY/CsC5FTkxKkiUYE+
Tq1nWJ0RlDBt0hOFQE32ITXA28++JPQt/n+H8ivu09zDr8shzfZ0lcIAOt5RNSfI
7NbnIpndouZ2MGxhh10cLfVmIlBYIXwXqsS78PPgwC/goYS6l5twMsVm44FkbOYE
gCjKVCDMT15tsb2OirIz3FiUj2b+S5+Y7Qv74GzWcWgcF7xBxUh5sPP6Mx05VAxc
LGi96SvyQus0+1Ov/KiikTjVvjvxs/8qhZZ9q9aJazEx4pHx9Vok3SLSXwqY0gb8
zUIHYI/Qe30+hxkT/Z/W3VoTL0IWkjqtRxjVmueIQJNzF7dk17cdDV45o4so69mr
q9oTcSPxR0Pk/EIltTadDUpzrmAKSMQnqonDFFC3NIwgbNeJytkWV/s7fApEXZ19
gtITpdYv98+KxbRuW6npXPb6UN+TYTX6HEuz4+WNaHyOVPdPlbDKHuGhcYiEmg7l
rYXAnBO2yQov5VjLLPw3U9vgaih33wO/BQ1k1qNaD3/BEG5Y/C8eOh6jdhJb7piI
9lMH0NGWz4ePuPgCuyX5lw==
`protect END_PROTECTED
