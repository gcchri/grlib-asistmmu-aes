`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5EOp6EGmTP2u3Pb3kDCfjbxWKigxgQ7GqJWnp4vUqId1CM6q9IOg61pHTlLuVBA7
cHt8AS4BWu0YR8WbGBeZ/zs481aI6jeMlYkIKwzzEFAb6qrzwAmrBb1bbC0S1+MC
QS0sfUzEP4tqw9+dkXZ+ZP6YM6gECTJenvRSuiU9WQ0AyQdWadS2bfo0ybbLCYcr
S/gmfGzL5r7ppBW9T7Agf/CUY53RUqsUrDvDOYmVPkr9GXC+AQT7OZcksMmRUwcA
FAUXj80A8HJMnzMIRZ6RPIrXxHoURHp293p7JrviZ2s=
`protect END_PROTECTED
