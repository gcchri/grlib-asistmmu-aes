`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LSgNRFPkszOJHx0L7uC7vPXxoH+PCma4G3JH2/FQvk1vGeqmqiOTE1eB7UetallH
VejxNEXioLHt/ExpBh0CQHKuwURNenNmOmgwuocWBBq57eZqEhRTy4yen2INnSvp
6FTeM5RzSdVOgg6GRKBWfkY5K2vOVTW9BY9yiIf22eydgtJ3mfH5FgNb7wmSiuiS
kYxR0PNGbAT+mb62+VgHfxf0dTu27k6h1yPspQOJuKVJ/6H3oMR/aOVUdUyA+GBa
wTO+KiGw6YUnhBQP8wB6ol5YPIvtrF1KUxkQIEd6Dkpq3QUOHU1se5GZr7JsZ6yG
`protect END_PROTECTED
