`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yTCYgl2BozIHyVLdWmVhv1Adt2e/BcbXLpxAbYH4eFEMa84yduRQCqT68S80fLkr
D/10FDZXcM1KOcMY+ADJIrp0RN/SqG6HnWrGzZ8F++Oh7AX/xVkTl1nBV93o7Znm
FP2t7uUFSlGchclxIJzOuKkNaynEGfY3oUbTGZi68b2LVpC+/y7v9nWbvHCW1Ts5
G59Sc4dESwmZIYhoGzH6RADi/EGYmecPncw1Ev2BoFCkpf5JReIPCGBUSzxYylvO
eM7YHlaH2jTMB9lbcdwj/CfLhGyy+TmSKyPYH7S5XJmSTfuD4btjvYWRCnwTZfnb
mdKEmfqYikNUrkTFnHbsBC2mM2dHuPW6+prEBxfs7zKs/adPlMNqei3lU9jMlNy/
VzwArauJ5pkulUn9quYomWbxjXZO9WU+QlO4fAD8qGKqd9z4AOonKQ2UCnTI2jCg
hJeUdW7jH1HrbXRRnMtVbgo/d5C4GbTLrSIv5JQ5sZpzDj3adhGoyi/VSjT4P08S
FbvVgy1Vbb0jSd6bdJ/SY4es8uVC/5w8aFZac0BcbkQGPv1Kb84hEZQtSPtcJV6y
`protect END_PROTECTED
