`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A/OBVMP3gKLI5RwhwXz+0BlMkbmIDTMkDNgBMnlz7KjUxh6DHKlqZueURyDUJjvL
Er56iuewb8k64vke77I8AUuB1pk0SWpEDwOftgPoihp8YSV/nm1ewKF/ZJL5tsS0
UKlUQsUJ0PAzk78iU6aTNHajlRmOmdH+m1GpGwK99nX3yh4oEq0ZQ0DB2OLOoXca
UxefbQyU2HjEnteZJoNCGeMNapgQaGur9AYVG8nP63/O6rkaeYpltWqxOAwcGLk5
+i8qupieKagoQdQ4Q8obvpMUlGTnDR3m69/t3JoBia8lXqtjSuq3wMqKjLB6qcul
6Ye9ggb8M67uAYEaSWCKJA==
`protect END_PROTECTED
