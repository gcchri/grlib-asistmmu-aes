`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WYxJQydX+rYelRdyVxQmfWE4G64o59yw022wf2Ih9fQYCFvKpAnAF1K7CaIeDizy
nDDHfVHw9+D83bfWodOmMlmJzP/ZE+0xT5LAGr+8fHDGdsj4c+ayZidsMBT+Ox7b
vY3KX5BZ3kspk/0ZFkeRJDpIBnchNZCZRUn0lip5B6/4/HO+mGBJqXpb1SZsOKaV
Fbu/hPc/N6irsen6Y1EUi6vJIe3gFRuHKSn6bPuR5fL1BTJHmLekwOMOXvePO0zO
a+JYgleioKcr8ydKahYgW+JZdKo5a2wf0kU3p3OnLwP90bl9pMfkL+rd0oyS8qr0
cMHE1Yj4IAGWVyDqJ9ez/EfJz3qc1BCooGnaSjDC9iU5kTPEd++BDTVWLyh6a2v4
rTQF7Anp18hk9yq09JC5iqtwTycD1uYwSJWEfOlu9o5Gs0CKR5s1JPJVFJE+J+rz
ycSzIhY0el9EftHUHXxV6d4MnWII/iTRcQNmEdu1QzulobXUgBO7IkCydr9dQ2kr
o/crTZo68gRdJ5QZGa6lIOpOSHTniSpUvKmbPniPD5x8uQoEdL1TL7ZwTczfZkng
uhjVnn0JeP3OestzQOV/RVztNko4H4xSdqCI+hZes1xzshEcYJ8CkjvzdBs41n24
jLq6y2TwPqzSH0MGTecdxDV3VvUjdVlvfztGH8qtKdTH0VUQCJMyInz/iBHgzOZ0
qnDjqfojqKqXH1CcpP2TaIrX2zyt7fdOsjVQkbzh9AgRoL/VTfu9GJCugcBcCrvg
MgtE3wRcHvhLL+BfLNE1ekF2j6MNFqkycXSfsXPOlD8Yfeo55SGV25vXCb/qzS6x
/vz58N4fi8EqseWWhEjBVG0nMt73LnGo+FJlFfYprwljS59lZr2BlvaPwnqVJzK6
gcGqr6TiuHq0RrRhnxElXj+2qAFc+ICz/ErlFW+Ryv/WOp0IWLtTxzSSoZj2pbSU
u7/yVV6EzkuHHldvWuNqn5D0RfS7KoIcU9kwyfZbFxhuXXAKETpIyGdspCeBgV+d
ArpaGiS1g+947Z3TvWQ5PA==
`protect END_PROTECTED
