`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KojobsqAB41A5Yo/hL3nImPygQfKSrZe35pOk/2Uyv4eKMgl/7jrzZ3rJ308h8XO
vubaEBMb99wBZAiMQRio/F64iOcvOaw6NWtN6vUHFC58DmA/MhvE+5rzjMfLN4EA
MH1nY3JOlzBFpt6tamYriLD9RZ9TAAo82nujkmLWyKir3I7FyDNXcpdl4liK3Jxu
MnX5jCaaTST8GCGgm1LbTkk5sgliSQCUM/8yXrfVZGBATbE2ohbi2mCLuDMDqlWD
D/JEAP/DyyRd3jXhUBmB2l99OWFqpRmfQ/p+JVJoaIzxspNMen3niJgUeCdBGxma
EXYi/GhxQBs6CuD6eFpc0MDXIXW+GlaphiqbfjYej3DvamgHPV/Da/nNmNadyybw
isTxa80srmFxgte4xye6yWCqIHUzeINH3AMxODiMJDGFec79ORXxZ5BUKBneM1Nr
yO0vZRHKOIuDZ7IilrWCmvZNdm6W/SP6+mbjFU9QiMZIkZfWE7aiocR8+h8bCWpF
YxYPWqEFBmW+yhNRJIpqR7tyF0CpsuQDD6u4rJkDRQD1OyeISwD/SleCKYz9+ke6
fyrlg6QEuBtNPGw2XG5S2X9Zj6Mcsn3z0x19+D4jdDdCGRqo6HdKBZuBNZSAhfXQ
iZhkFuKYa9WJmE2sV8rmJbyuG0y7G167jVCixELKDJP9cubvkH+bgRUFosS31rmo
KAP4rpmEJr7boNicosOOYmorLAVE2iTGUBEu7WhZ2wHowq4LFWJJlrOT0JJFi1dM
CtkqeGfkVzaWGyFcF9MOtg==
`protect END_PROTECTED
