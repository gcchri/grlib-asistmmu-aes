`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oAyWhFsEfTwVje7IZv1e3/Z65TWVnqnSeWv2+qpevSe7uus8no03u7Nk3v8gkvix
ZNc98vyGvw9Hr3i9Hs78I7s5Jfn1Y+6PPZnGXr0xKREWjMjmPk3Yl4VKszT/gtDX
qqu/cjqISC/y+trSbhaTN3OYshRlbglYiKcoVNmJ9fudIDVswittUJj6kLJaDbuM
Pj8QArf8UZCA43/PicZj78D9CUVuMUjSZjTE3tp0AgwbYvgtue9tKinHZO1SPjy/
mMqhYeDW76sDrktw7xnLls7kQUESWWdf2JESMOMVAaGrVlEJ8CEMHbFf+RmOM60g
QR6hX9xH48Id1VlKxGpwQQ/NKz3Tpfrpf+fhqgPAhCvm+7DFYn8zAd7il7FbPQeK
pBEzA8YbYv3Lo+GpvEAgTPb4u8qwyb3mk6pmKqOa/9PbufaCeiH166sEc4O+Hd+2
`protect END_PROTECTED
