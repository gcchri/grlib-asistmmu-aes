`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+1xoJxmBt48E97K4jYbNB3yMooacSBSllUv2n8wIrM79XlifTLL2wgFSGfMGxXYp
Ugnd1jDXACvGh7gMTlBidBqNhhSfpsiXMQ1HWYp/p1oJA9LBQZf9FpOs/SIL0R4m
v5b8OoJrqkZPso2JEdmJ8i9aEr+PJ8bEorlbHxdMubU5eml25UdqOmiE5dGIod1S
S3bKa5AIFB0OOh4OGrbeC+fKsX9uxws9DWfSjemmKVkbw1SH1eZB5YHsNIu+tk4m
npdT2LTTa9I4JKKe4lyYyO6deXUbZzh/aP6G0X/rpiYWtMe40NAi8EPjc8miYCni
t4ieVkQebILeHcaXIdcHmNrRMz+WKuj1fJndrO+bq1gDXngo/g/1P2cxFrANfAhh
wYtVf3MxbScYn/mlSlBExWXCDW+3AevXMhrXpSYDtfjYJyyVwJSOCK9H9cYXUxud
2UJopJK8LpNYJasOIcGhwju35/6wr0fp7P0pZJl1cdlU7S4Naro8nf1RhUwBie9v
8orgjoLiQQ7tR+zm5RGxXvw1T7vLF/DuK7bFH5f0Jt9X+bbTEKxMx6t6myGJ1Pb8
iMDO58A9ThKZxj/7YwfSgVTTBMUDHmtRsMk4cg8C4IfLSYJLrSV9ZDwmD1SQPA+l
sdbLt05aJSlwNMsWmYC7AnWnR1T5rQsRMUUSjzZlifafMIJtPPaNjombIShzqgIU
Jo+VA5PWBqKD9Ai/y1FKNEu9DS4BhKomfWHlC/nK4GE5Ddo8XaW0FjM7LUjJVuwY
eKt0JURmSgPAvBZGEbBzag==
`protect END_PROTECTED
