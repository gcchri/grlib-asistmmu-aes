`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BtrX2Ns/DdBw8PUIAW7m+VuVrHRxnlnsq3Zgf2O0alUwMWoFbjKnjoXadNDRNCw9
r8sqIBZ5YCwVk+grTW9Ay4G6qbQs4Mj67mlyuuKAqGuzHINXMXMY8jcg/FZvfWpa
mrwMcUInGwzYYS1P5q0KFgnvA9M/pTMs13HJonc8D102484lm3uA3MNdZ3qwDYHa
6XEUyu882z5EhSaNoAVdmZcckGxSE4AW+OD0HdjTMgJHDaS2Y537tBZWTjcAapYQ
j10ficrIt7CpBCl1HmTHqg==
`protect END_PROTECTED
