`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nILLIZAvKQDRXVZK3EC3e6L59pdt9b9XzqZPQUEwzwG+5n9x2MMLKN1gWapXPaK4
aT1shb1mQBanG9W5djdUwov+KKZT4Ae8DV4dMQa6DR8c7wEQSCppyxmBmiFWo7Zb
ThAlC0X17ihIwySdAqLWi2ZaU/8fzy+ZrmA+H3nPhcCaBRFwLXJXl2c3MQRYnjON
kmpZS96BLOgCMAMEwJz4ZyuzloegF0PAvCK6kcgby5bolqBWwvpfwsRs/X2sXcUI
SaRCUf0kU5S2aHmJOXKdfmTuV2l2s4NH5xiPtvISgqjOUjzHevEC5UoNr8LRXdGN
P6OjMJBZckXxIvHgwdvGrOQ8VwC1zdGztu0ebDqQzctPVHIW/pEsTeLOzJ8C+XbU
OBnfIp1S9eftTsingx7btux5U/vNpadEJL1xn71iaSAI4k4IMrfE3FLzgcwMG8ro
DwQ+Zc2XFAFFrm6jsoYVAwOW+SEXy3tgOONythIzwwtY3uqGiBB3zsaDb6yMYv8z
EaHEPfmRIHcAyObED/r+2lAN9S7MFNA5EPQu78OhAQJidMvupaF7bUo2twxFcqSl
eW6rMXutcajUl6rW1baHulAMCoUeC/x0Q1f+c+kdpipccR7O6+6Fr26RO1F2cbFP
yK42YxwRK+HfnksXCaK4IY5mXWtbWypDhmhzmAz9JgMLv0iu8U1gYSLmbEPOb+KV
nM/F1DCaxtGLivUZumrEsMYMVzla380AVJu8U+7heK59P3dJw5daYi2HHlTV+wPu
`protect END_PROTECTED
