`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vHmGuYE0a2VPIULoTO1Tn439imxgmEMCViZ1u00uvJktLk4mTN0qXY6/Yj/jy09Z
49VmljfP4gOC7IZANoNi9fvh1sbpJMVltY0GO+lwtZTWQF0zto6+XNIgUOGQWo28
bGSxM2s0imeDb0J/gn4IAVXa4xem8L1Gfzgg4jrPoYQlTguRA6OSc1Xl/5R1P+yo
6QNnPccVHBF4VKU16b2QKgiqfDoT/uxIEnh0QC6XowhPPhNW8uMDSFY+DPxrimcg
8sbUh8YK5+lAAz0reM2pwkvxIzPCLpB50aMHg7mT92c/Nxh0ZNRe0OEDuPHXhYMF
G0P8/ICHquv9MwhNYrmAkXOBLbOJXNQraBnarOVpharBXsZEnW0VcK1xjUaMQRVd
0W5x53XPIxhdWWPVebBEUfR5yKHfDGPniaDQwWhWf3RtzISBAVSb/mg0HZfZzZNJ
wI4lpjhGASI+gwG5QoQPiXjT/SkobCQB4yrtxHYiqDH3tB0mTjdem+zYo3FLQmZJ
As1t4/0N4VIO5AHw8Pv+HmyDZFYjFFDAswRerQsL5HCwK2Rwp1no810dGG7oH0GW
Dfq38pDcnDrHroaR2nvwGPQu7Hg3MureWzu79kUXVlFiP1JtuvNifblo4Z9rxrDw
NKRTSTEVdoJJ3fp6nX3O31mABNwOVrfzeZIifv8D3doisJQ2rYPtJyIX9kWXqhaT
RVILFLFweNwt6HSIP9Q6gM46pdad2aSJuEnT+JjkRvHrxloq1AAdMbsixBRv/ieF
eNLdDKPE5DHGPTzYEO/ZGloyAtJntBcOP14LjjOnHJXLItZwvz4dItYsfh4DLWfY
0UmEwnsAj9kiBsP3tMCwyExbHBQBsYZlkU4ZKVbfNsAYSAfUHOAkkjo6mHRbzs5b
dC6T/tQgq/Ss3yjydE02qOK4y/XYGHDknQBjqcxqbpX/uKbHhyO+SU+/p42hwrun
`protect END_PROTECTED
