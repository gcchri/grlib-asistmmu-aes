`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pB7ppXNBDDg3yw7awCcbQMXZnOVNgw0NjBwWfba9j+wci65HAXPA8RxK8jhHwjE6
iRnhaUFrTo/4MBJscZzsevj8SpkbgNXfu2GnhybBt8jkFaA1wstN24bc41UAL1gi
vd+H5llqofWhuxSqAEf8kU5E/6RCg3IyfqXnQCAGxD6hORr1oKvt+XGWV5r/N+Cm
yPmYQVmrxvMg5683aumcf9y4bemJO2UW39YhOwwo9ptXjlKRQOgma6H1hN8EqrR/
SoEpvj3xZziMWmdylfisDXpIpmjwdWIv2u7pfvNn9/jPryjOzy9s3bTjSUUfb3uW
WIATWLTIDEp6Lx02LRqQhd4naGSYBbYwINWCk/Z2PUTZf/QrkOipicvhcRIDAvwW
d40GBjAl1f+LXuHofykWeAB1Vps7C2h48DbJKSyW2YVgClnHLsX0iG/d0ElYD1ff
cHvGqWznVAURnfER9Sf7RLBewQaPPc5cKCLTwmmS9fUMWFgszYXS85SxWPGhi2oF
AC97xZzObipdf0XscikbGmQD4NIFP3/H7ba1C6MBrHEFnJUNmWrO1D2FAmPuny/u
OOIzTxrZJN75sKkhxD9vZD5/XqBhUhL9tfuq63ZIISsFQxQd04tRYVszPl6GA0bu
cMYykj60JwKrAgjEH9KZAg==
`protect END_PROTECTED
