`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QRQSsz1hbisIk5/A8OcI8fj0QCa+nohjdyX+TRnaW4D/ENrms3h2h5oPUBK4RuZ0
qjTO5+ycmTHR+j+AOgm8jMk1xLAU4pr0dYPuJnzTM3zRZ1gzPejIGiE5jrApa9iC
SA1WAAemYmQbPyN6e/d75sLVkU0EgIG8W4hCJ9YZDnfyTD/adRDVbvWRvXvNre5I
uTTv/cDgeKX59+PcAttBEw5VW8XNqE6Q03TgSvX6Q7yFFtEGM2a7xO00AdWZ5Pd9
hssWxKf9XQ1fIeD0jd1KDfKvJwRdmkxlE1vlJQ8haEsYNDbEbQPTRBbqETyzh1vi
Ksb1r7bO9amUt4NKY/txgwA9YkNY/slQLzS9iaznuP01467LLEcpDvi3FhohanZN
4Z1wlYL+QBUkZd+VNRYp5Rq8NUd3wAAKnQ8LRkcvr7U1Tr19t8OHhmtWCVQqO4Rw
dHZrHnpKWhLc7tKqIoSxX2BuiKKPAQyz4rWCBgkqLdt3ZgmGEYq8jaJbTnSRtEag
GGtTRGIOben9cTPOsb9lEhWwBwAUWmG4B2L00T1IBiQ2yZ2TqZLi+QUylTmosKLQ
AVCqCaQkZLvQotB0J6QStv0AuUl2hRhD3ihAGOApwhVIk7aQ98/CxwyXFmKsYVFx
0k4vGt0143jEaFiS3fZb3M4nqCUsoNLjhdcD3mbSbAE3a/bkEUq4TjMhYvA89Wen
Jlo4KDFCaX5kdAYQFSG3sTghexpvYg3gnUxqa3pskapbrw/x27XkEtliXsfBMV36
W57JYO7WzRv4BpmrQAwunzVHT5wkDvKsY0WRQdNiuzN1dh1pyQC1dvtQqWSxESQ5
Vi69m9T9A8pBXun8LgNKUM7LUCb3vI1uA6rzOFNya6ONOYu+1jHcy8fQuY5RE5oD
EClAoycHM9xsrVGnqxSI69GX9tvQo7tcv9CnIhpRA//Of/HbLa9eayB9a8g5zhZc
HmqDAIY5zRa2/5fWjmt7yqjtSqbBZWX6C3v0pgNcjtvhehGATv4b/n6Mx9d423+Z
Y5hh/FnC+IGQKvX6c0WS88zxitrtYnRjo/zyD/+xANjatgBhr5JOgPALxyZHXLIJ
eIuliOIIA5RvWnxQ589Ci3wIOCg+yFbeszBiLNHrB+A+39iKkAfzPIzWED7Yc6Up
fZniDY6IhlsrafBgkf4uRfQdODBM8FNAOkS89BfrLATrZOv4jOZz5K2PnhBN7WDT
YNsnr37FCvlUH+CbQLTrJ5xmsht8rT8cwXVUO02QmI1OVHqRbZtcwZw3+XWiI4YM
97jKn1+Fx05tv1Ngu687BGtFUdkGUcr/O0TkS2HNSh1y5TXbZKKxfBKx0vawlqGC
0qeLrNFr9P2PWUr/jQhCLC5OXX4nM01qUTgFGn/VEXZm1DvDFeMhbZ74DwCvMTLW
lESUn1AxhdOat3ozNy2xWoiA1QBES6o6RRgvtQZBMptgBoAYgMk+Iy5ZZEump6hc
rbCbTeN8TEHws9U9Jz9SIQtF4V9NA6FMlIJbVXByIs1BGLG1MmjlXQVfu/NBZwfs
K4V+AJpg3MSb8kK/Wk7x53OK7Cda1xzy1NvAkq3WpxHpvm+knm3IkLKdOnrCAllu
01ZZx+lEIRQg+Ily37FKVaareo5Ytl/Jr7r4R8PiSOzN2sOtCb/NW0oopZ5z4Shy
1WkgdMtYqelhpCEc2vLQ/A==
`protect END_PROTECTED
