`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JV0U2ttZVfe5KAJNFwPP1FBeWPdzdFjr3jEAqDUt1SKu7u8x7RXkpoaf+AMcawEu
E2Tq9c/0dU0VFt1t0lasOl4hk5EVf3WZE3z8YHJErNJ0fzqVsrv43N0qdtKhcVxL
fMPdtzu9EtWRpyuXCqYLknt34Ckts73ib1kVEmt57TecCna2tJ5q6Gvkf+nwy03M
Zb7B8225AfOWsUHTC42EVh+hPGYBBLOETgVKLZw+0wGXVp6s+eHg0a+odRD/gjTj
RfqHp+iAZtVjXXGEazKGkjFlTRwISMjzKI+Fj+o3HTd3gtCMxsfwn9SpUnPmKSC1
bnxggeyFHa3cKFtnE3x+9VCDzup0lOv+CeSdTwExlOyfXrwPajvQkbtFpyofn12E
aNV/srRNISLQyvaTQNcxEO8NIa5W5563rKp3y7d4A9U=
`protect END_PROTECTED
