`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rxhSnbh0q3jyk37BsQ+MUN2CJXoOD1fgYUXEEFve7U4jKjqsTF01SFZJS974v32u
Bp/PNE87Q8Lz3oyC4mkSHaTSR1vDbZJdNxpwlwhqxaW6JmGYRc929kuY7Gw374zA
0t0QpBy2BlLtZ6NO28oiTsx6ejAPVKF/TSb8stjYJAZQFNnoXT69oJxVKE7aBiy+
GXAsCvkI8gPpfto7Gbk5wAB1VZ02Tsy21GMz369+pXla1HiH0tIXeeLLDVAxHtzZ
xwhuosX8Jtp1D932ugHN/N5E4iXTK6MF/4QqAPZYKceWqrmVijDW4+j0LYon6ctY
`protect END_PROTECTED
