`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qHWe9w185fzHr3U/L3Lp+1RSJBcezGE2IKnlmeC4pevylDAl1N9zh21+D3jmiXnH
lv48fzAGX7hPGzv2baqhS+kzE08dq1UpjbuNJamvD0g/T6RLABH1NsnLTOP+SZWO
sLRNMLDo9kpHTyp67/hVzquzpVnRO/BVgOCyQQiBAX+ZyC6o7QezGBK+wR0p1J+9
o3rwaX/93kvnnpqJVxhf2DPb8df6Bb1HSwE/K2s6L4w+kw5Gk91lobprB+5z9u8C
90sZhNpTj0UhPBfEb7kZYi73TLbWqTNUmG4J1J99JPp2psIsBZtVYxB4szZRT9IB
k3HpuQ+L0qUa3ug9K6ejYvvpX9qKSBKyl13m+IZ2ADp8/8yr0YeySwfOU2d+cLYN
1JmplzUOwSKhQhG99ppmyILgK4Y4BzKTAEMxCpnvGvgOSsDxBk89SnXQAa0tBpSL
sWzbUZXbqXkh9FhPzioycXy01BDrSbvT5zDzWq0vUE2d7Wb87Uki8eSjTkqYARqw
E7Z0Bz5nO1P9rqwmBkAnh3EfShXWIZMZX79Ga8gWgukp4pOKGjNJ+zbIAMXiNFK2
cCRIpf5QLMCUmRIE8yhSLp7698rG8rWjxQy+Be4HBALC2c7oE2TLCooUbgXQVZ2q
yD+7R6Q8zPhX17yNQfvcc5nh7I3oe290y3fF+VhjciQIGmJpyGBSD7O1TERW3JeQ
iwSw639mY6rdURfQfvNiue2xT6bom4t6dqghNPVjVmW9HBYPk4eCv71DEe7Mj++u
tutMO4nsoTqjeGF+I65xY+vD8rctCIFTlaaSZbjTC61CiM2kgfU3CDynyH+4g+iy
poyKw6bFDo6ExyBPdMJwB1EbICEntF3Eamjft+GJ1/eLkGgE/Tj9ZJRaS+K430b4
IGj4a1GOjWBlYSrf757XakQgQdi7xFs2JAdc1lf7nEdjK0FVFJ4g2pHNosnM7B0N
ElOPdyNmCnO2K8D6LvjdrP1c+A7kI978edlEAfk88PLzSGUtQAlKpAzPIHcjqYFx
iU8mvw4gUcUaS+aXX18qkd7p7MdLRFGXmf9G/WRyYlSvXXuIAj4Qq+2c2UWMuMFl
3ORodiZkjbmqN0CKcGCWHhfLbzmFsfx/oskeynXy72xkQ/B66tXKM4Eon3MjF+/F
ZBZedbQf1ObJ5z6OT3ynS7XgjupkiPQEWgCjZ8kUVKg8LGx7Td7UnVIwtgNRPG/R
rwm64DL1FA5PTYFoMlTD2wWt9ut3V0qxmnPWUgv7NDL0f70nQFdSxtfBWb+JxM3J
dda1/UJaXf3gclSEgjBF9LEagUqudJH1NzD8Uq0nDv/hnEuM1I1B9x0XkyCOO5di
Gq/YXrb+ysxyMeIYg385AbGJ0agIDMVizgszwhnUh1FB4XPtZN5LQw2+0OXndcva
kUKbnkcox3JG1uOc4eliQCUCmQpHDMHOFKylF+/Ec4N0BAgGsiTjE2tC7YDPBl9y
+b/Nc+RCo7Mhb8GtSEWaUyquUPBDKxNc2byOKTfbFpHAkkuJ4Xf7hjDqx7xyM4zu
S90+K8zClE3TMHfSrB4EpeCNVkjlI19mgkyNIveoB0tEduaMGiT8y5XtnsDvfqHg
`protect END_PROTECTED
