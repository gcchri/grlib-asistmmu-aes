`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c+nMBPwr4Wf4SW6zqJsCsbyD7SST8vlVA15haT9v9s1c7y/8Ad1gEbT5YG2cT6SM
YFBE5Pzx5uGwGsq/EzoK++MsZhyK/0znctUQoeDDR3k2yCkruoackC1gS5cJhB78
wx9+gb42hx8i5BWFSMvV2a9z4cY10EDS9COcBfeDzBz/oSnpaGeTA8fSDwQIU4lz
Xqed3TaSbGfWcuw2J1/PY3HIaSpYOONJVkV/0ci/VCPDfev2PARI/g7ALhRjED7g
zBMSU2kEvGI/WO5LcS8u57sI/zeCBEPjXp5IsrJ/AwXWMrYDx128uxCyXeo0KdwY
CYal/Opdhvkvsikp35HvouHHGRMXvdmPcoocZg3Di3F4IGGp+nv5z7BVtIAsSV49
JV4jILDjXgQ3PjO0dfbLeYhyHoOlrgwHU76UoSEW/Z/GT9zIHzd2BQCzNOIFMTHM
HJGDd9pr1jmAkEvi+x+2KStchAzPOB3o2BKFLpnT7u3YCSpoAzU4HZHm6mNd/60j
Gd5xI2Ezo2tTSrDfZHhOLN4qPYZJOw+kv0czI5KKHyHhMYQoy0s/EHI/B8CCDGtz
Ddfsi+U37grAd7+EkxKPUTF1rMSO53gpOH8r0rtUkBzK9XOQdEh0borB79h3MVlj
Av55RL3BBTXaX2HJvLUSjMWCAIEJzxhT3nFPEO7lF6anKN2O1ULZQLwCTNoSB/sF
5LnQ5aT7OKxEbTPa+gZVHp8FSBlb7RVGZBd8NYhXvtMn9y6kj5eZw6PWRwV5HxJ3
+u1tfG8GGAG7XZjZD8e/Oz1eLw6IsDbFatuHMC3sMuQqlIbvYSIYfgzgDXZiO1os
obb7n8zUCfgu+gKaCgMkMvOkaIa9nHKF0+YDne1u6JS00qX/WpGmPPm2wLWUhlL4
fjf5hyv/LDgS9XZoYjLLtfj7nyVSuQcjqZGQeGRzYP1dpQ9El7QqGjASSr37JF1u
K3OF3I3loZB+cP1+rAJnuqowZIXN1v9T/hvzbaw2YSc517c9MIQJZMD9VRRWzrzE
AqSnVGgr2i0su4Us7FJhPOiXcPtlKfUN2qDPyBYzl1EJSAKQOskARnFyTSN0FAQ5
k3J41gEhOGp6Fnw1qPcI3Sbyn7EXhVXIrwh2/PtbhJaQELnN+wQ9eih9xV+HY7VR
Rk46szpkpy9m3PnwXJut7hfsSX6NJEJwjhopjBh+T6FDWMrKgbZMk5dLS+0ov0L8
ttKaghOVir57+qV9x5NTr+FOEPEGe7kgsAUztK48az3+N6rQHvEbFvtYg0DaVoHM
WJyGRZ8p0XOwxK8riAuKNpSylbphRg34cOfYlo6nBRkWKL4rbv62Bc6Go9p+2kHZ
QdOWVQC8cdkaVCWasRKs+jicCWAB8ht/+3ewE/VoUUBH+fJ+Sxm5kuYP2YF+U1d6
iMA+6ZI0ZywbOJH7/uxpDoklM+sori7Xcw45Yuu8oerK6y5fz5oZOBZINgOF2dY4
uBUE0YJgGV63+66b+o9olMf6+rhUlSZ+q3ZQ4/GtGjZzv5vg0IXZS+zdapQ65u7i
ZfSe4jd3a+rOleWxI0ZzNrMMXsH80Alguwb3XcFYoil92Pc4BFbBdN7K151bVAXS
nPi8yu0B3RaRR6uHUBuMSb2dSw8/gpVePHGzQxk4bVzTvJOknqsbPTqjedtLML8s
zU+LYLuMDLYABlTF4rVLsBaRDfgJL5ho+TM2BGRahZ4tTJDRBaehrQRbrPut7d2R
pgTWGYwKrEzu4bhAAdef7kBywFHrsSqAdrGuftxglwlWiFfvRy3fdQzO0R6X+Rtc
Zm6XCOPp0I1raE0WItrqOpCV3FTeuSpi4+u2AG5k584k7SE0wL36P945/oyFHVMo
xglXjbI/cpCOXaaml0rlSDaP/tGuoqlj04ZPxW67BPaJyfKXzYU/SAPnMBH28yP/
cSlBb1NISqVCdYrIaGXkYrRGKx9qAI0ta/YOT/wPMrE3BG6Kgq4k+wtc9+261glF
TgEyjYQ1aEU+uVKS/hmpuwMCfaeLVfZ8bAUyMvX7vxPNDyXY3dJ+KmfejCvo7WcK
rV3808RQiR2wtdDJort+iecniw+vVQD9QNsm5svJUiJWJocuXzHilsm3cAOwl+3p
bXVn4wA1fwyaLlXwJvAh8VjNO928y7mdNUF+NMx0wBln4xtERVFPaC6DbxDNrCqv
ovJQi12/RoJqPILNkv/mD+ddZtgLZJvU3pAYNKWeALuXjZjq2pEU2sX5cxJBfOv8
HijOqbAo3faGfEPUTh9meJN8Y3qtYVy82HUFFf2T9gv5QMyE+5GDrfZF/e0Lvbi/
aJmsJNrtoWBs88rErNWYR19P6mLMrNfj7pYL/inUfRM/mJBPnflIqmSN6kz04p6w
Z556J5vIwZlEpvKP2GVB78cU7qnTgUiY4XX0ucBmCzN8kreStRHNP5o9EuyUneqJ
vu/FLTaOQtIi9Y9Q9c/glKS+B1t35Cok1azLHgSY0SSQIpFYs2A652ci0+LCpli+
QKEeUSWdJIrxu+h9M4XrZnOhoUYqAbpsbf1s4nogPhSTJKmCqWFmDuyH22LzCLOu
wWTW952d7Vbq4qlT0RLOBPUySof+2BxVmRQ0Q25jOpGO9yibjuFbbzQ5KB1KKEoa
pE814CdAs8AWsMdLpq2mETYzmz/Ui+WgmZiG5QWRR6iWtxPGuWBnfp6p58hrCmsU
5ia93wkwNOsR2lBOz28v0gbEAgAQ0sFCV0KB38wp/YZujyVrYIQjiVUx+jKs9ojk
BCWE1TO32iAxwZHIP2qJhTDvhnow+1quZZhvQKW3G4UjNtTFdXWKS85rqzoLo27i
93/Xr6SgjKkvE0nkiI9xrS7e7Bp9ic+Zm/IR5jM1OlpP68b7RRA5PtEQDGJnwDpp
Im0ht/Rmeh6voNiypREvxA==
`protect END_PROTECTED
