`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C3rN6iX/nBkHufkzP0amShrCcUZOuQ1dLMiGRMpN5MFRBfdQ7j3Ffs1l0R7v0goL
RweB+SGQ1Utj8fGjtmVK5C3Uj3niiNZsK2FTlj51Dd1wSq8xBeitH92jLY9MtHGu
gRTFuLFQOfqDO4hVUl0Al81Duw1NB68Z3yjSxOu0shVGl3SIMa7BspZW0EpVYHuM
hFUSxuh7hGnoWSIpOViQrSuCd4u6meALNjpWvN2rCnw1f7zLt9o/0qhICszSGhka
UtcY5qk6BR7k2NWhGUQfeg==
`protect END_PROTECTED
