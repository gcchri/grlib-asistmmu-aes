`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VpL40IuoojusUgv2wzmL9GcnjVdaaYb2eZbqi9jzBHRX+PmzItdN7p6mvS8Qg6fF
9oaMSpl03JerKNGLuGMmgGNI1cgWBRyYrwLvQgpavS7QtjhTsOM6GVxqnzq9sWez
9WTYde9I7YSOYY/Ozuzumk1GgF0J3NijX35vudRst3X0opYr2D2ZQGzO6g0h3Rs0
6MoK2As5dY9iD4owyQVR8xJf+D1wArmWDgrHBnPOC3IBMWefeQPKhW3ArZ+nSBN9
kxKNdH+5d61QxGFxbfsuo7Nr595U8/JHG5hzWmbrCQw7p8/1goV1d4twzMon2v4n
8KzLkANVtYfzjEFNqckCgByhBQWIVMaGD0aitqkLF8meAt2klxHcTtRPspkrNwty
4vBEyu98gq8yd1wc60LVXfUbk0a94YAeA38hSueZDmopZNtnkcMSi5HJngyzi9uN
uvgU20v/zyaoTjfNiivSPosgzePTcJtArZuWgQH/X2aI6fvgjxZ2bzq7aLD1iFs+
QbzHdWQXIvQc+rqKtR8VV4cgpAGGdPRb+XCll9cA8F5zf7jwPc5jVU/H54LJmb8v
AKfnTE1WJU5vtUq7D6kVbbb/bBQu0avHHtaBhjIaGBMPIKguxRz9Baaqf1GJiB1j
tlZ6rnjoNX9KaEV+CF3BotI8yHIi5JFTyz32zWNeJG4BE26anpXMFwP3YKJ+YZsm
SwE0I1FomhV1dqzjHyk5Uco5DF3IlYBIFCKwIE0hUjE0pK2oCpZbMdlTxkBrN8Te
l2VRGP/xqOfZZu6g29E7NhnZNYaFNSlLk3bpTAKYoaJnjZYi6KY1szl+jSQg6eki
`protect END_PROTECTED
