`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EYgpWBaJbf/F0tlZfd4nPSLjxOltiYREdUW8VuGYBemf8jKIboJNB7nG4OsVkPLO
B+4S6N7ao3BbZ7hRBwOYhjNFUQzTjQ8O8NlH1fK+/Q0PsDQbBNqaEspIU89CUy0q
XxoJeOH+/Ro3FofDaGfZm4QSU6943n6hJad1fVL+hNxGz43Ig/0C81UMJMJiGHM3
Qm0VexpxUD2nKf7JKopDY2LOb7dcaKZQjYix5hgrw7iN5FGfY7o4cQ1qz/QzVgb9
kS55UJa9Ir/bfKzSyriR7TMTkP9LjvC9okfY8Gm8DR9w8TcM3b93osbvVH1Aqw8z
4hUCHORTCeXWE4aEdwwjPcZLJiYh96BYJtQPAwk65ieB/GiaDSgG5aQNfQVHp6fZ
eY+nhM5gR1RaHRp6RnctqLIr7JUByP319icqmZF6f/5az/nMHk4MgfkFV9s+oRtW
NdFXk3tYQWN74FirqcVO895FB1RdliQk2NFdawfqcowyIJchTYTb1QO/D044O8Mi
B5myHKx7eVpgYpzlYZhYbwZL1QYIR04i8o45E1auSXklnMuFR9GTN/BgOXz3fPAK
`protect END_PROTECTED
