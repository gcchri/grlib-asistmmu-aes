`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MTge19Dn2G/h7CZCmtq7eQ0uJePIGQGbP8rHmUvLubfc1bZqLvya0vRn2QT3WjdJ
hVvPwF45SSiTYeVLH7XpI77fc8RNgYtzkUlHz42hLfO3ytwRNZGyI4gz62qMSOme
RYuzzngkCRUawgfxF6/Te+cZEYoXTpjF+h1TYjPflsz+5bCngVqk3CXRzZ4Vc0Bd
cLTLt7KbJQXhVluaRzkrtoVmoKWDyCwsP2l9MW26Vga8zJ1DOUZvtbAu5Y4qKZng
o7jo1IEddgoLz+vS+xKkCZ9xn2aFRzdrATYKiP5Aw5A=
`protect END_PROTECTED
