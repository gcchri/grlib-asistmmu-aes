`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LyPpbQDNLVl9NgEzhpAqCmZT2wquybl35ZXnW6uBdjSRzqVWzz4IvVYgQRvS5KQ1
y3/A/TYTjiUrZCZbTeO9VKT2kOM6+08+3/2DKpwJEtIFYwseMFPyIZB6G29ki+Z9
OtPNtJHeGxNTgda6n5vdh1m9vDVG2+hjA5wkNkyz0671AyMAmOdnfmIVeXCuy4hl
32jH4ohIKwBju6tEjiHz9mwHUH5mZBq2ztL73nKipxpdCB+uJ1WgACeU1ANh5TEF
HIBVzvvm0Jug/GoVJ0o1vn9vlWVWOOu/QcyL9iYCLyDgGnxP8ba+JtYLULkImiSD
2t9899QRDeiL6vL8F51WqsYTDZ5Mwh19OeD8xgJ2bLEE4TDHAS2vhh1/tOKzFRnd
8CaANUkHFT85J7bcyrDP7Bt6J4Xen+2r4PI41gApV6JKLiOsXwctJaaGb9STyq2f
Q41nwCGjtHqT/9mrf3Y4+5ANAflVWi5wV/nRmCfitUDIzRojJ8RlH3ILPn610+w0
5nlRNmrzJk6LKEqhHjRT5GOuRSKmhjpRLJA5Nyz7pSl1D86Vap9Z80YSBoQY0ZlW
OusQsrQO1h2DyIjmnhTxBCQnAp49sw9RSNFauDygzctzS0iB179vREnloWm0m2k+
`protect END_PROTECTED
