`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+4+17sE5AeVJjoPRtyoFpK1ynlwWaf7MgAsuSz8cBguxyDY9Ombhq4ewn3obcXeN
8jzU2zB7P/OjoHVYwoxg3d/1VXWph9OVKKUKdEvehzRGiuvsW5DgNqJVbLjwhs7V
gfbYkDLQBodmABy+nprOI/qTBI5iTFmIxSg5sO5tlWphb2ldJkb4pGfyn6eZln89
6/uhOM+66SrSsqbaQFSSNXO60kLTaUzGyiNyFvWpTxb0+AlDcSDslFFBtnNArPfu
UpLaLPhAA664FdfKX7WFkEXEPDSgKtRAkbjwGC76v+cW6EWFHyvmN5lbox0+lhFE
gBicn37S0xSwms0wPBMFIQ==
`protect END_PROTECTED
