`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LSzIXX0nmcGepA0/WJNMHMOuswjMP/EGu+cIbsZmYJ1Y1/Ld2Cqga/k9NCw+bt8V
Qlp83EWzUiwJzI6O9h9GhC/dnJCt218+iMopMNyJjBvZIFLaXpwnQNcSTJnsEUPP
ddw/crstZnCgZhq4u8XiFDPrVu/5grkM2xF5akHQzXTxm1FPzx/w73ZKikWx4+qu
8p6U+31f00VjMDPZ2bqTCHX70s00dBUwL6kl+puHkbFIEY3w+DrIOgUabU19Yybc
5eSS+qd+idiaFcN3YBSBBeVIj7hY2OvufgnXAb9HrZYG1ae077tgJ1F7Cvby5Owk
CsjJiEwD1jHlBk13B1Lc/JHbcVKsqbVRotFn19J1jkgryVKxTrPsu0komzj+p+yD
gX3wcHOEQf58fFNbNi6Vlm+6gsYmz39S8hoLy33HzZOPcZeP0LuragxoTqJcP8u8
epGl+xkifBc4ou5uSfhVxBlsWvGeIMaVueHHeTljOR2Du8SQavJgdxpNhYAEBuRU
52OUVx6QBYhhSeNf4xQa8utvRV+1M8I/3SMBTiST81lCTlMkaxQRb5lOu1OCdP13
wMkMiVEJ9sEU1Sa8iQt4Tn/qExQbauVksMBpSS8pAjkYAe90QIN1t9UwleDgc8Qd
J/XthgfYZpx8D1piW/GIPJInf2UNfHTO6FostnU7aion9BUiAR4ZUHo2mPMqchpX
NACuF1mnY44hUrO02r0YVDqhXNI0mmITKpCQTl3LkkWLTuwKSQqtLu8GnoAO+mMU
z/IqAOdzmgKTNorLmw8foQ2biJF1L9Uv1up1X+iDnzYE3vGN4n8O/8ANfcOcXOX0
u2wqwXm1nbA7FHEWys3QRDYIh1nS+1qfqIkwDPkP5murX3lklkyHG88cQ08Rxj2R
oxi8XMOt9/4CqVlHljw8Po/GIV6Xg46lvZWmgeW8kd1Qp2LAxFyOYAGZygJsnvqt
0NiKAE6C1RtxtOG+gTEnVc0mfnhY+iWakR9QfQ+1BeFhb9pj1LQWFlKMrWh+vwFo
z2m/li/Np4cWmRRZK3nSf7GCHz+shCxSRpy3mArswmYANSktVVRM8KV3+0Pui1VR
SgjBPgmiYdzAN8/PuZ7YRoUbZY3pBUhASkYyozskd6uEdth7J85wWgNuz0X1BuxC
4KeaxH6dxdhMUlmyWyHG8xjCf89BtelqgzcfgqtZ5r66px+H5ZqOJ8ahz++ZQqlP
50c2FWHoJBhWwpVeCF4qOex5UtYBZX7D3OpDaczG7web0x+TYdXTzHlQFZCEjqy9
2qSYb7PgPwQPT3JdBW6zzGrtfCbdcltfv8GblP973yDlbhecWT91pC8AXAWrFrsW
hg7UVUs+cn11d+9anoN4Is9g5mEtG2q0RaQQdTweJkXIGVRU8/Y6vsJ0/ba1Z6C1
8OfM/Ud4g/JnDluFDmmOrurz7gHNeG7iUhBsTLKzp4x43gMgo4ApM641Seldu8BF
dyAUDK0W9E8Jw96XhJ4pd3nO7kjphbwZjGIGvemp5Ecz9Mcbi6Kv/FQc1Taetsoc
/D4sogVnfSAwMeOdSimQbB9IL03Z7rDD7Qk796Tks8pnQfVp7RKr59NX0kpTRiHR
EgP4jBayUl5utXXAOcFEaRihudiByLbSZQppnKCNmoc7CMHV6MWwbr0zaDaXxJKT
rKAv8Rkb+sYEPX1MAO/4u6jbdwR+VpMAI4uuA0OOrKhEFqfIRxnbTkFOjIDYhxpy
/5M53xMJvugO5SpXWYGtVE7n18Pe3j7ZrJRNX0D/y+nWn0M3sS28sm06BhwYCC7o
pAjmJzog7Zvil1wFmtszlTeSkLhjgNBiTCZMrEBrQa2jHdhAU6SpFYm0MMZJzM5A
sjS2INO640u3zJFkzCel5vXDW+wFV9rkR7jRe7kiqXz7fTgbl1SpO9GQvterpAuZ
vey2GRt1xHvWgxCJA+SpFGTpEkD8FAXUW1HvhJO51EeHl1Ty5qW/NSTeQV0fNp6S
JmXfzjga5iA5RuBZn7XIOPaQw6O6k5l/hDTE6WhRw3PoolQSRDo/11IrpbTCfB/g
0O6h93AKw/dR92VxjdxgBbIm7uuWKg1F47qQJgFzyDc7J/jioONL9I9oyRpZBtIi
5kS1lwsF+01QFd+2eGiHzvBWYO+Kz1z5VFXu2YVpuuVAG4BCGJtMuNGBxySuuH2Y
WknpMzr1P9gf7of+4+FxKzvQ83dFU31uHWtWLCho+AQm+8DrLAjCVhXTbe5wK0ZV
kHmwlL0U2YVClwGZPlS46IG6ShcmkZoGvJnH78jg11Tnp5sjuPYdAKwpTlErCCAf
LjcP2CilsbIHjR6dTIug/UUaLQ0osD4a+F5Mt870MSO8L1i3SHAVUnB5A5g1CuRT
/kOqB+v4/TncNChoIk+XZg5DhfL71dlwtmFnvpXf+6xGPcrzqmko7zcXl2fPmaM9
dOdKJM4Fs2YLRybOjuB4TEvF6S5R+0oIAxbxMXO2a/x1n8rLp5VtBSa2FB9irX9h
Kd8h7HHx+4mCa9dVFRvdGBhMqhHgCHOth4TfUq3PFY/S35PGUbNuoxTgiG6APtph
xJwQiUtTOb9duZjcTpTmuiP1HXGn2bPDT3AshTLfCRAlceynDPlr932bj8x14YWN
LTJlCd1yTkKKk3Itw03ydvfpFLzLwy+UBcJkR9LO2YaofstPB0CdBHhYknHj8acW
9cEVuVH/nG69j0sP9fGqNQQfxBS0AbS3OZsR2mfHWos9bkgoHeKA4GcgPM2QfqYx
DeFuO6CjimIQbTx4nensbusH4lQ2nMxJbt41c9Qpp2YNEY7CnC+VzzsZPpyhux71
TIGCySxFSZco84DDFxELwCuQ3mDSRdeyI68lE/eYFn2Q6WBOuJ+ticnAmCdQibHI
QdwzXbC+QbqgAE6VTJK4ylI5lC9FTcV6KSGftTCfQ32Tfw7Mayx2ecaFFYRQY1aH
B9GN6gt82ETC0Sy2RKubeU7j1CEQJe2RKbPmo1nfwzKPtCbfZlo+j6AxS5cnZSh4
7zoL82l60elO5P23nF2LcSYuL8dG8RTPV3CgBoOvOaIO8jzpTT1kw8oTB6jvTFw+
cYhIiarfH3teHLbk/ckAaTO1IOIvHil8dsnzBXUbx/M0uKAxq8rWNwTiGdDbBbk4
tBZjxZj8t5KW6qy2EY0nDEhRUuVUbGRqhHEp+mc7AYTTaZkwy4d5/fvPmnzIPI9R
`protect END_PROTECTED
