`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M7rfCHK4rvhPUlxM1kEnoo0fvwrz0TIFTAMXCb4tSFS+ZLL6J35x8Hcu2Cb21ote
WhoFdKIpRT0BaZEU42IeIGYuACX6O6qm1I0yv56s5YLt8Nz9XJpph5yLcop9hDcG
VzVrLzYkrDSD8jnF8AQaRC0CXhTl3/XdgyD/IF0woBWCzIdDFRrDAF/Ks1oc23aW
CRQWagSM+muU7r/Ib6JxKNM4Jfeq65w0tePPTSF3rfhoKc3FL7M1P2rr48wXBNGD
YHA6/0utrgUaNSiqp+t3aJGCeKJj3PmgqgSaYmd00jC746/QNjO6xKw/YXwilayY
ayNtMNjX3EQUvQ6EkCN7+m3kWzp7TQh0TA1MvbcQW8bcRa949UtkJWFyVTHhORto
Q8zAMV5XP50hR6H47aHZgkPOp7iWhoFJp98KUy0EZOkzky39h64mpZ4SsLYn2qQN
9K65ADLEDmNoGGQigYQXd1AB4Ff97+Fi8SAafOsXY9J1H+qa0y+MssdnC2aHsMVB
yX0uV2PzRg/+9nDNDi0qUltvpszZBow5b8rD602RaR9EXRTEWBR+TSbf/kPaiKRt
9xL9YrFnHjjX6sVb4LrvIzD51ZjUHtwap4C1Q92ZluMrLkqeCBqOYcG0NC5ppBER
w6LT91Yh+39ZPrHF2X9bMaXDbMW/9dSeHuniUshEa0g=
`protect END_PROTECTED
