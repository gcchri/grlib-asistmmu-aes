`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
puNs75ovb0+AWwKjRq2mdCaYn90lY2eK8lD3tteakqCTY+dMfBvfZRQnSmgBDQ00
6EClPiSpF8RJqL9AMX0C0qoUbzl6sos9pM/XmKQR39nouffq9xTRzO+t+7DNoPC/
3MBuW0AAbGTTVysixbLiUqXm4jHAgcDnOOm+ibcOU4RV2mSOZHDYxirhq9RWoobB
pZiN6K1Ifnnx1TnrpmFwYJYaQ4KeK39ec2GTjQR6pwMzo43dJTrhnBb+VVlGZSMl
gckQCWV43OU+8SVEHRwNnv8LWJmG0QcwNGTc9OhOs0kbRF2S1SqLMtxRfkGKnh5X
Oq+nvNPKF5DEmBfjwV3UeqWeeUdNrtTWG34Ep8PYMQIXCRlDX2IML5OOU85Idv55
Umy+MuZWqBucZ3yEWyqEUECVc0dg08P7kGGNfqrIGoxSkLGdT0oS0QNJS55Kpl7j
RVyoTvqw0W7laWCbecf1RbH5QG3Lt38sRklUgtgy1NBSnAtXwwdFP0M4rmWnyoMJ
EkqtiUIdbo07guUKgOkPtCJPgZGu8hfXbhUz/BrPRkjAI5P2nB64eHkow8sQy8Vs
e9azYGJ6digUPK0pbjo12ugPDqtAO4xW2DEJMU/sE3zne9a7115+AbLivmLaR0T1
pTw5ulVhsIFtPurrRO1N1tRcWS+57Jj+Xa/tu/Bl97I4E042AtEQABHSWsigEa71
d7d8DRfUL1Us3AXtLy1XcrKrReY5vjeH0U6wEoDSkRLlK8Wo5tAnY4HvUVDj4dL4
28n7q8OKdd76MthjD2SnfGMqpJ3rFQYcjIzlplW4Ooodzz0JO969KmxLX5SkpfWW
TvQMdmY67ffT8Szwj7hlqQu+beC5JPja3++nGvUG4U1PSn79Pem2m6DpElVjG2r2
f5LXex3IukE2lHhLp+ZW7YQwLgbd92wWnexaHSSYMgBm49O7ucClk63xKiUheaiN
ht327kYT7KWmeMkWF05GTFHw0SPT2U/EYj8ygqA9rFzpq+OjxMBUxfJZAYxDjYFQ
5QQgf08Ge1n8zlhguwE00Q1MuCeCAI6j4GxT5+FwItQ4xcY0SoQKkc012YIgVI+l
M15uPrrmh5ytf1ABV8xP8eRFXg/VhqiddxGtSRpUlIwgZzVwzPssyVIsDMGCicNE
UlDDZhZ6Fa5Wfk16MdCFlvKO/uKX/F8vuxCxMq3uwD8xx+XF812G9wvKwdmbJHWM
X/uFxSixlkrLUMvJgsUMpz1Iml8tfnwSgOoWgkFcogy1qou27ZZ5tkhm/4oV4weB
igPSmkD4spoduwXL9LgmTE0FKuLkuuQibPeN9U+30zWY4GYHI2/78OUHkx6EEvdq
F0lWLvmxgxUqwGIbykUkDHuOqZ/3BEXp8UJDv+xASgNVHNdluIrj2pLSmnD9PmOd
CllcP01vhb8dTs4w5GpE+AwUH8nKRHAEMMgHeJgdkEGAIjZ/hsiMh7iV8EHa+fUp
HgY40r/SVSlquF7cCpOOOpcQzOrdHJx5fiv59ocgaYRAKczYLBUCSnBIkCjiEyc+
`protect END_PROTECTED
