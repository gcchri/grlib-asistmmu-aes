`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gmel6k51Y2z2yqovjxD0GCZkrNmOUzo/YxHyBUnJRAvA+VLXM/1NYLX8P/LLeTmR
dSeNfvPstF9Yr15kcvvQSiURm4MC+NOF9paqSWoWHHELqoKG+wooT3fbTEqoq8k9
HVi6wvZPWgWv+8+fimyymPUFNUWaQPv8F1dlV2v6xGiCbpCysoFcHIicFcsrovdh
4r2aOgQu1BBtpMwqNkVvTm0g5UBI2d27ssF8cNq5ROgjNygtP3cATJNnuOj5rhY3
ZjX6UF9tYpyjXILDgCRMZJPBzp2BOQMV/19VZT841dvcYhu/DpAVxkD7CYsT9+gg
jyuDvLxZ81jP/Ei4yYR10R49cGH0xZGpg1b28SbyjoFXPh2SOwPsns0RTAcJ4aCY
owbmwgdW7DNtteqjEbOgeLbxltvDjsW7OD6o3V6lT8ZDvnjyavghyvl7yHneMz4T
`protect END_PROTECTED
