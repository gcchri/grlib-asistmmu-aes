`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gvJldwUshe8Bilwcdqk7flqWQ7oaddAKStieA3OQHiiTmLcIFgCwhK22jO1HOo4Z
C8ALnVnPETlA3ALO22oMmpjiF0RjHVnbi6PUdK2564NYNsF//iFOvESuVt6XhP/q
pfCrsaDiJbaIX8nTw/LHl3QE01B0j7/KfNtq+nMHupjulNgPLAdEkOKLIXcCpKGD
1RBCceEO30/VI1ehpFgYUKO5k2NElhqX55oZVU+5B91UHBYcoZDZMMkoNs9f0Ije
Bkxwoca3BN/JGYGTV3mVYNbrNX6Yn1JCCxZj8RsiEGyljhI/B1Idzxu2CgZCddZy
fQdVb1FTF+77x+r5u3cktu565SfJbiyBvYXXhbFs0TTDZ/WWwn439nMjXKBRp5FC
pEe5wkRowKx1NyrlcJsgtA==
`protect END_PROTECTED
