`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FuVVdah6piq8Q1/5hj/4gju3rZBbIyA4K9sdtk/003/QGhl8LgdhJvH9/8p9/nMj
xeG4p32rIeC8xyA6PGaFDOu18pAfMFV3WOxirpemInFzsArqb7zC6y9SRtZaXowV
WTWidRGIWiBfm24WVptn9k1bM17YMWRCie4KblFMG0VTjMnJVEVcbHpq0rJB9cgE
NYfn6eOE+LIQW9UWO2NK5NlPSoLXS+JOkkOjdQooax61iQnlcg0ReBF9u9JYx2eT
guNRmP18gAnQmdLZpIJvw3RqozXmyU49TCBMhRBDkTUKhbcwAITWBuN2c9AFZYBl
PkzlzFtCZPtv5kQQ22kyuO7wz6QUzOF8nk9KEdzHIWYTt87BxunUL5kkDi+kr5WU
2+pHbs+6B6eKXtrH4qOogCrlDWVhpEvRlrnNOnCK+4f1jlVuYE/sZbzfyXDKVrUW
KySDxMqNAxmYBO0bog61954ZwjYpGJgW2kCodAXkreiJUyTlgP7d0C+QTtCha5QW
`protect END_PROTECTED
