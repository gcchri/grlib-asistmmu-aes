`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m/wmgrU+Jhsiw7zDUPqItBPndwGG47vmlQ6PEK+xUUhdSairi60Xe6taSK3ea4jY
kyEQeaeZJ7ubd4/zw3CWrepGAKFclLIwlpnV9H9wk2xtgyJDtc0xeFpaxmlpDNsW
XkJxiC2xIy/wmzemNh1rAQ5cvwAi5TgoAPL3QPzrXmoIrx+4hsfIRUVXZwt+mTQt
O5bwRLjSxAuLfpCjt4XXlS2nkB1L6fWu0WfnRKXc8KyWSDA0QSfwuXerCAS11wLZ
jYLMsxh0VPDAOb1s/pGc6V/etz67gBsSbcXFiibrg/Acfp0/VCL7itN1kQuHyIVU
HxzbwTecdYOvToupWWS8orEV86IObexHBd/+prkJ1x8xbxBXjbUG/j8qErHLXPE5
bJoBJiWGUYI03Y00HpYNTVb94gxxzyp8phPj8SiFzAwnAyRabaX3gO96V6s2D5DP
xoPRBn3edF/ucSzRVtDQjDF2fV+MvqJZR7r6HEXe18iqGtwZsUF0I4aVm46lHBTO
Fk6+wQeG8Qh8V9lhYbco9HFpw/AxO0gSEU5WVE6W0gCfdTCj93sVAHAfVNyl52Ul
BWD6eoeZP5z/rta1zf1PJkqvTAiz49MhpW0KogAchV1/9vUxqJhSg791drJfCIKH
K6OobOHh8qLzo6nqTbFE4ly6b89AS+uQ54mdp+f72VI8UjZ8K7yQwg5MDgogngb7
xwWKcGaXY+PPChOPiGaH6qEnNT4+FGgYAtuEEK714NucixTKf+cL23raQYtTXOn/
nAYJZx/HVgBv43wJJKj95HCr4A4ENeOortexD3atcHQagTNqg25cy9JkcsLo8TgH
qnHBEvLzev2QkkkOwgNV1G+vJ5V47R/KgO0mvbX52wRdlhjdJ+pxfk3t88Dx3MBN
5rGd6VESpG6zchZjaLQ69nFMqosvZ0HoQkbxlWlLs4eQlVXxfdBc4pGzweb969v/
Ju5LFqfQHZ9WV1oytVHyssZBDn1brbP1rAttt6iqO/pdWGm4Fg4xcwdNFR1zwV77
D9LvmT4L0S53ohrh4Q/2s1mWvKCyssZOZKDmBN2PZ5OJppB/hboFAKEE6CDH7803
8gOZlAlrsuiWimWEy5XmDZVDp5jCg0zkuXbTkliOJhwzrl7/Hv0PwtwYwu0drfDA
m0PevYd9wMqzzHM4XXRdVYi9ooRiQXcykBNLyFmzZWSAD9TjRSjk5gBIz7q8/CPF
m4IzoRoWhk+pR1mEzQqjPcfMoOXnZh5R68SgyK7tmr6owCYaoqJk1ufp60+JTIfo
+VL3dyG4ikkFcftHGlG3qGR2It+oB92eKYlJxD6GhfnpQAJIPuOWnfiP3mGTAQCH
WaBk/nk5n7A9fTRshCq8RxoCW9S6AZZyj5su8+IUjcILOoaE07unXZqdvZbR5MUi
9BuG8J3LICxLDXslj1dAAwwghabuZ78vfvmVY14o+OMmlEET8XBqh8JwWb+lof5j
JvIUsk3KRTntWytXjVna5lxQuJMfFv41r812bMYU+J5gjJUDwysQaJV+SIL/sdMk
prAzKcjSRuxczrU16pTYJEXJxDYlGY98PWQGiJB5l0AfwvNbopWTQsQsp1f9HVOt
BiGfjDxgp3oVHqCPUgJakMjjSB7hb9XPEd/mLSLh9cReB8BpqCzZ3QYiD9Jsc3XK
gW9/TznFgr3uLhsuh2QRO+gviG5VD4rrYqvmyxcsYKmCtqToQvltKYZaiF5v4iL9
m5uot6+2rs/rk2gZ4boS18hkY/yAqOR0i3tX08exLesalVW2iFjWeiZDa8ng+pE+
YBHuD+4DCv0V7SD+uARgZzzP2q/9LjmIcYMMPj9rnvExDYZ7tQDA2FQzeugcm0+A
1IywwWcGRb78mFQWYGRXwA0gRf+QDuAnA7DwtQNrB4BC9uG9yrsudpTyGKlc1fba
wC9QhzVqFNz7k1nLBMYvVaszXko8t49AL8dLq09/RjsWzSLGnrp0YUqi7pZ7trmA
XRsSMpdqwukdYoGm3iVPERZ04E2Xpsj2JXSZy7cCnOo2pf5DzhF4AkYelp/UccSW
0jfUFCLIYHuyuTXn/atNP79XkAwM3a6+cq2K57H2sP7RndgN7IgBmRC/0WweA/s7
mumbP0W0DJlLLoYde6dVtUR+t79pFb9u3ULdyghWw44cL8k81oRkP1CSaBBDH5pO
`protect END_PROTECTED
