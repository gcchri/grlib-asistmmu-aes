`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EBrcoV8iRtSXLzGrNbTX7yzOSFLGVREf7T5hfk4UYMkpBE+PbRfslFuypWVnRHsI
kJ8Yq6tF0VOw5BFm9qhzbhh+jRVqV2Ia9tI9zf2QluMP8h6IHWPbmlmh7WuV/WMi
LnutKovh8HYm1CsiUFniDHVuIsS8qFa2lfroOmfOCWPlOsKG9fpCkO0rGFqi7JAs
I/jo6RMnVh/JI9RKP/YohLCUVeNjnTr2d1phtSj6Prh2X9oikXrXU67OtusLnOl/
wO9OI5oijW8MukFwbZugrxqANnWJjJu59YW4vmc47q3UC6hPN849mtdu/F1yJ1U+
gmU3BCcYKhMbjH0vmkxsXQeB+PJio1uVGOqgCJc2pFYkVsmHtA2llA+nnZiy0HyI
VkRqcAIEii3WCeT65TUJSg==
`protect END_PROTECTED
