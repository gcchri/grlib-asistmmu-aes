`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GzgdEAUa8AyKqWE3wU7UlWN6kixLJIBM3uWuYCmio55+we1R/CcCTVBY7UZwh54I
IemANYlGSD+a8YsNGjiF3Gn8Hjjv1zwQJM9HxnoFJ7+8O2I7AtASIlq9ubIQ9bxQ
Pi1ye7+xftbVDk5AhxfrlUuLtiQExjOecvpEq5/aqpKuPe1pZPrphr2Ap9Ymqzuh
w2bCalIZqElf5DWu6hvZtw5n6LbGm8jU2kXGFIK+2haEArcksTNKVSgb8dSEYxty
bvRNgaVHYS819Y9XCnBNIfUxkDX/1xwd+YxCYWZq9FVu/PyAQ26AV2GfYAz5k3Wg
SoAvFEGC10Nq82ppMZzsVgDpO0JJNlFxeVroJJluvDl8ykt9J/5HLxOOt2ZpetUs
PgxP0a163/Fos5KiQPKnNg==
`protect END_PROTECTED
