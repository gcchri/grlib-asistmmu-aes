`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QyZCcgfbw3SxffrLzv7tl+zerAc90xEiZqL2LjXVzfRzd3U9sZAzKhIRTZ+l4BZT
yUqmqtPjAiIKx7q2frJoqaqSj1uqSG4U6NxpwuLqgO/nI/toPsruJcgF9mgDSnL2
i3Gih99pzywi2ZMbXTJU1tKL5AslZObZMIOUMJs1wtrN7S6DkH68pCWZDTIXXmKP
Y+f3XCN21E+KuUL7dauEm1c+9D5asD7Fh7NKoTUA+kZ118FoaBcNIPE4beL1fEmz
gEzjs6Bd6AovVcPqFP4dew==
`protect END_PROTECTED
