`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a2SXaQK4vVEob7aNyNQwHfrCUQwOJ+ESJLknm1QqmcFatDgiZtDpakZdmJTAJeAk
PT8jMtvq2L4wq7qWCcaDKFC9zM/aTn/Lev/74HKoGvapCOIPEaH5vIrHC5xerxy7
m0XPsyxYWJpcb3sfXVdkaO0fncjP1VzRTY9qepCQZgaudcW+MlBtiuXfMMivh7/h
PX2TBbDk/pcQh48837BUqJNlqz6BVBLIZMmHGhxQr707rzc/u+9aN+LQgiQSykPr
VQlPt+tTZW+tQNj57Ar3AhxgxTSSNeOSb7UsE9mMo9Y2CG1ZgGpaLQ5GOF/s2ZAS
9heu/0HsW2QOZwxGxRJrPKaRM5k2DJnLlPUqPKm3l9u++0Hs6jyzkjl6XxnaGXwT
ZjUbgRSPzCkG2p9TDMpUr3RvLFeUtGLK9TL9eJ8syEKuiDawyrjHS9+6RqmmHjSv
nHrNa+GV4OA5CHy743ssW7tPuFI7ff5w/LexoGPmkLmitJIT6GaczyhJdTe5WrfR
ifEcLIh7oBB2RHE7aW5QgnWHxxxVQtwQuxKskZ+UxjzOA3FC1W03eLoJz9Sv2wCz
9saJCPcfBu/7cag+dltKJ/YbD+kihPqX+HewpBMpR9023NkeWZH7pZCPFMXYimkk
j1FuJWe69iWC01LMMp/qJbNucXTARFPheWHmyIf29f8/zjL79fGqd2iICZUJl3p1
xoRDwnW0zvaRslxdOd47Y1AWkhUxXXlGvzYaUi3QTnlCuodrLo+XzHz/+HjfogqQ
yyfA6V78wtkT6aHbMi1WUGNr5FFa1ffWWfgt2EH6NQxOmkvjlkC4UlZ+xX0I+fu4
voHA9b8VzEHFNTTM3cXJnO5b4vh4X7cLHg4Vio/4sMr/fApNdVEUujBXaDZw0l6q
yvZafvQdu4Iw+idASzCeZ0WNK0xY8sENBqTrmrgZg9EcDsbn3V/1E3LE2fLq+7Bf
QyEL9/rLg4B9UTVzYqjrehn5eh4P1cqQI5K7k6IDTw1jo5w0TgYhfhjJPNQJMd3a
Sr09rPFj/PTn4wurNvajM04o64vM/b/a3ejdj28OmJIf4cHhXTjO2X4XBekjLYAR
H9S6wVulClDtjuzJmHedFU+enWhZefnIaSr8/ulkdLnJWzfUh1fUyvQqjsgpmS83
Ua3/v9h6bM9EEcHNMCHTGuy+riwyyiSQ3CVj+1zVqic9nMI7plknDJBwXl7Yhb5q
sJRAbqJHAUtQ0/n/qnk+LQqK4tXqpOFEgxGdka3tXNY=
`protect END_PROTECTED
