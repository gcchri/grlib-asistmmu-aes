`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oqPcBG6HIL/CAHWgZ1UTQjQLUP6DGc4A5AL6mw80RF2vfiU2vWUvVPqZwtpqk4Wv
KyPJ+fjaoWL9vV+IwaRRvNCvFpfcQEvepbW6tV29ga2D7MJOYmz5pqQywL+GPmBm
fhFra59AtKev9EZuUTu2YWTDBHSlIAzarESUmljqizXFFYMlOV13ROP4TGwQhna5
1SgEb8acszBkHGkNWqB0yMLqXxq+vllbK3rEceNsdyhL3v/eaQ76Fs+6uwpBFgwU
UklDLQch0ws1EzV4ze7StKBO4NwyZpx6EfeS9xGaSpUW0gjbWzvtK8UYbQgh3Sg8
+KHQsktB9lZg1qEbAa2xKMWgzBAMmhlWejO1j6+8x3kDI4KY2xe+0303NruFLmI6
tXrEIo6nQ9goMvrwey6OlraaAjQIn0xhUnt0qlfvJNHwVJz1E2bdpDZSKNHT7rYd
MKy+dtrLYK71h7zpPuC5yDQZbuYTV1WJPcD9sa7/G99Ljjb4utmYV9L8A/ghHQ84
`protect END_PROTECTED
