`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lSavKM2J4aPHUv5KvTJ6gfQeeFsdtNprQQmOee0sb76yTy2dRtZTtFuljy6v7lDK
eNtURyKREavldfeTIVscPAmDbSqaBCxwkdu8NZV/LYrWaHpwiraasq/r/onft4kB
emiX3FUDbDJO11tXmSwIj52rL/ZNNvplTl5SgACg42GTCqOA9DIKZjohj29QjT7I
anCcMYyassh5+3Ccwo75LMYgxRO95QhUpOAmenfGwmpN3g1iOXwaTw7mEvNe9wof
mg5OD7rSV/BWnkxhgzC47DzT72E8mt98BVvtwgqIns4t8dWe7EQH+wsCoeHNI4IU
DafMlpswApIi0e0ttijKqCs1Vvik2vRQbJCacACt8DbIZDVbB1Xzm3Vr6qwPNxsC
`protect END_PROTECTED
