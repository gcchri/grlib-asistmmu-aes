`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iFQOZIsAOqLsoJtuDee5WMdjr82CsSGsdmClMQR+0lWcsZtstnvDwObIH86v5yCI
PqwSa4UzjLyMtDd1zwKiYSRUj5t0Mq37McTPtWPUtTURNBBIAdy9jkvy++CSn9nS
rYoTjvdnuG9ryF9gHCTnlg7dQvMBJ8+aLgjgFkEUcxGqNxbXhfg9h6Div/JUQnpj
Veoae8yLKHfi1vriby2QkSN5RPehGVZku2LnuBS9V0cUSCjk/ehPAe0RQcjRwC0u
h62hQiuBydXkObg30AJI/QTwlkC0FBFjMVOKXrAphrkRxq0zkFylGLwHkdbXLArl
1qrkvwGVfzdsJ0EZLu/efZPEH6KvjMPUNmgXAPOtbVsnuFrJkQwH0p+fWKfgzsn3
xyMgxzeUxsGS0iAMkHRiRhRKLONDUXzBi/fWKeJd2gV28tMoLzc+rT/u1DIae3Wq
i9+5fzhgAzp0C4KnWflTzOcixrte83pbbNXLCF+DFycLc6tnlpkXUWVlY2dg+WBX
X540rZCOghoAzkv2CGvC27HuMj+a8RnQytexWjicdE+rLFAAETKzRHp/MEq7GfKb
usdat/xGg8yT/JowZyyvHig8mdhAN10FS/HaNaKck5/a9IpJ/5KusUhJHFtvA/jp
yKKb2lUx/8s7tKdJq8oozYx5uhsnAR5KeQqCDRHsMU1LM/gVeI/fzgbAsVy5Fm9r
`protect END_PROTECTED
