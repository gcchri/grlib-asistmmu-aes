`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nptF6Carf8HwegMfTf3sh0c/CDm9LtnzfJHVF7OgRfWxtGLyXL61fmGJmfMm5dB7
ACSJoZ/Q1WO5oz2F6dL6SNLgbkBFv4OMTdML9WQDtvLmQJNuoRhf4LuRk2NKc5XA
U1SsAAR3UkPO+ddsESPjCZpy34kvrMwqwpQ6PJe4h7t+5XwL63HpgfIDK/lmBHhs
0mteIszticJJoDCHqpAsYYhKpMZgxZATq/jLZmzWofqpChche3i331Rhk3546KA2
oa9N9MvGpC+VDlkdEg0gOV3w7ER0Uq8zjva+I9se2kopLk5iZAs1lv/R9+2wJZch
+bk1IBcG5vrM/8GDyzT8x2D61USply95b6zdVCOkFwpgurEr0/kJ3/+ywH2l2UYa
GOaCbc4Qe7pSEqVZPNCRbbNaxqxyiWnI0Yxblqhx/8tWWa5UcvB+ajWpepyH24eo
BHgJ8LWNJFrP/Mxqmxx7YKFYdKMoUvNbXx7/7mUHy2pLBaE2J7MRqWZS4BmeGUJX
27nJAd055fUPt248yYwt0WSf/VhooZ06cXV7kpSAnyG7iuejihERhmAjwdcR0Oq/
x+34GcE7Czop4sbTngAgmzNhGiRYoZg+bDibgI2kZZ4aUx0ovlgMw+oFQWUkul9n
ilMIphzFpWwOF+ySwtyPTEsmF25jco9DfFWu8dwk9HTCrnXB9F2B2vu1EP6swwLU
VE08Y39Qu44gt159y8sEWF0AvC6TOtbUVqpS2AvanaGxcEztldwNbGRJcXpbX5/h
GrMjKNWd+/DNzx3wg2WxS6/i8eNY2X9BjXwrYjj0Xb9gMXvuQWxFXG26nnqdIdUU
Ap6+l1S+cpRGV+AeF9djeEiLhslpvLO7wUUOvN5ovUw+EBv3ajNY8HZtvgpHfG7z
ZSr4Yzp89ufHjsvDuCZ1U7tOhu7YBD4I+jfu7tFV5x66WFKOCmzERvgnKim7S1Uc
DEqaBNlJtGzBQpdcI0Kgq5UrGoeXQHQGiskt+LFJF53vVCLaZbFLAtevHwYrgcNM
BO4hpMoYmgG8/oZ+Tnaq5NIe2o+sGdfRCjyD6FSc39F4OCH58+YWyM1n78m2a4vk
ncu786ZQVIHfyONhswvwlxTgbp79x+Z/b0kad/JYGu/xpFGkwyPVBfj/Y3+k8U0f
2syyGzkEpe2rD6rdzARflGhhpnPJmopYTHxU6+Xi+Tf4HLGt5W+aF1NT4Zu+1YAz
kchjHZNkuokOIlW0/0zZZN6wMEUPwcCdApKab0HK1YFpYNnZMQ1M6WBLtMV3imgf
7HWI0SFGdYEQYPov2WAjeu5hH4ygXd3H4Lc6/pYp6skmEBg0YpnIh+a/kO1jPtvZ
YNifbEe2BppH2L4rqCRDW8qDYWCQJaIsbDSsjZS8uz7coaXm+1oEaf1zM0JEBKfX
hd1xHFIbAl3bS3lhqhqXTyyMvjd1UhJRlU+2ANpMIezyk53wcIP8kH9jLwHdop2x
3Z849DeXgA9SxstK2NhtZw5kqD+liawMLMAqEDCLD9eJ+oYYc9szxuNwq8GjJVX2
p2ZzGG2AUUSselp9jEVxzh4G7bgNE5LJk580U8fpHohpSgCbBwE//eJ3Cq7oZVpD
TTO9j2eYmvQ9PzD2LzEHNFAN2+2CYZBjuWlPgJvuGbOQhRoGMUZDfo8djzRSaL5o
IzVRX3oHKp9TqqpCk4uivbgWrL+Cyo9ksTwXxvjCQTBbvnDVzwkENOMX1upXJuRC
Dfoa401FVNPCfqs0V5GNGKY1WuyAqXKaZlDv6NwPm1fUo3RRY4q6qmu3aVbuSuK4
Oje7fNqGZh1+t/pzdO4RcONslvFefxjJxtbWbX+CE8ADC9I3jqYzWNLx8Kjfz66z
rZok8rFvEcZgTUtonk0jcjerKFuM7iGRfHYp96p4KmfEKtBHw3ZwMKU8ydjYvDce
zAzVyrbqYKZOZ6m4fR15y1QLzZCXgORG5wHjO89yYizkwgvW5tdb2ib1NCyGmkQ7
OS+GsxGk+gEsL16bSVlGCY2F4dlFHePkAsEhUt7wNMOJu7hP6nl8LNKTSEUkiDON
lIxkc29NB9uFNN8z8BPwG98udaejPyyms7ln3mv0ifGpcZy+YAMaV6Gs1S5h+JJC
UiyLEUWBF6zjLQl3+kU0RqkF6iIehUPMvWeC6Ab20D/+Bh1Qx0HvuGqeXGKnwj4r
qjokrr++BjwhZ1MHX+PjojW88InwlQV/+O7HQsuUXXYgSc5WbQWCyzhyHveiRz2I
xt5eAVCDoj/DuBs5YJu7UG+nCf9q077HvLyp/AyI7A9zoRhewibtL/XCtNm+cmxv
QeqkN8aENzFeHOQ+SyuXKS7FF63d7let8+w0pzWr4ezYngP3dx3cZnBjLN/Po5OQ
LvqO/sOXecAI4Y9/CqRk0WyJbon5mbSMSd5DBQ+mTtSZb3TO8YcBTjZhrNc9gDDW
JgSZcSKYyA9TU757GVV9p/3+2DdfPVmNCzUVbXkbzWttSiJmLg/srNRNCx9s0/oh
5pLJaeAr3m4VAuvmgG77VC+nYiANKUStItWukb1GqBO0KA8GYOJ+HQictyhAVmf5
DsGuKkVX4kY57pOqgYEN2SV6vleW9Og0xj23/wnDUlM0Sn+ZZI49+90adEN7k4Oj
eR6vFxxgB3VBpv2WUn9CoHI1p4qTTycV/MAuUQSb30soLwkxLpiujvoL3b5DbsOt
evSDLOVxK7B+7RDmsyE3o/gL8KGTQx1cfgbYbMNIteY5hYWY4wr/8sBnJwhGgYGP
aJ9Q/Ewohf52f4TDZiwUUGk0ORXD5hXp+p1qjBJua/97xu9VEvnyTMLN++fBnOoQ
He7fc+TLPvcAlqx67wPCawfhnszrBGaphKkMTGJSnlyzfpVbkwT/G/1C4u85cpdR
XfZCGm9ptZXBd3Hq/bnNuONXbqH0k31hXqCCF0g0Eh2KjHrW2yeuKyVfV6VakKtL
z9f9lo6ejC5bXmg9UKUA0rG+CwVU9/FkN4BVw+khc4x3wl+PDVF6IH63HMo5DD91
+PC7HlL24GvGlptQQy6BHIQg+gNuR6F4DJ7CY1gOvgeCViR/WSAsxd3TITp/Sryj
yzPLYjPpTm5LipbUDQn2g8iw57tGT/blj3MT4Mev8tf3fYniP7bX3Tnp1VLHHwsy
vE0hE9Wbl05JT6aSJR06SUWlh+L1Y2SVg0j8nEpUE0Idu83dtFFtWQPP9fncfl7n
y3bExapspA3do6/dmwUjlBUFQqmaozqF9LP8fOhTXUFdKtfCJZZ6b3+JdhuYswcD
tgk+AAs1UbtKVmaxmR1uvcaRoeM4IATz9Be+IvA1Xi4vnFYCx+o5lQbBIeC2igwh
KJ5meYpQ2lpYe/yTAUxdDgW303O1nMrHwWEB9toMi6hEtDz+l76M9qOojUqKeXe1
grAccsHgE0LOs8NCRgzjqxCHF2iTd4YC1ciW8Yn/JqRfPiylInHu5yiPNMjgboDs
pDNhkISxweKrFoJGSVHFyO1n/ThBuPckwjfm/0sF6yRiZ2ROyrOQV2HUNo6skiog
+341b8tR0cs6v37a/0nzZ5yiaeKt/BGaDp+ZHAteROl4YdyurzOyoIVgRBncz/+U
QDj6Tfvn0+yeZ4SMmttzqtey57YKHgiGMwqX4lMWiEkKYuDL2IqdX6LSO1M7gsxy
wiu2+tR/139WSSAF3VQJwiGt69JqYDJgTu0IupIq8jVxa3pftc69KXmIv48v6pLu
nxUuNS/wTfmcjfBYh3GhcFDCKjNQdtBeTPoUEtP7Wafr50qKlst5vOj+XC38nhJE
ob3Vr0KSacl8801fibX2Ltb218xGpHv76UFua1QcaRR9RgR+efBKNx5xdzD1Dejs
RoTQm6kFyFKfLwxyC9zy73MFJv6eHsGUe1K6LVzEPjA++cNaNYaISiIQLQLWP6va
AwkjN9w2nS4IRwjGIo8zsXIomZneAKHYQDYkW5+2xfs2uL+EiJ7L2Y+5o7DIjUJR
G3PrMaPlbx1QNyY0VWqnWPTsjt9kRptfW720a+q3PzxU5Q+kFJYVFil6vAuLIVDX
wLm1j8TEzGP/fODEZkCdBWa8KRSxYaFDQEj4PoCC8cEjg8jFuOpEwURKrH9gHWnE
cmGxjs0iT/vk1qH7yYLoCVi8WvavAEL/MkOcOQvM9FSm5avd40yuFP/0KwX4FWMy
uYbtufErTDdcai4gtQtXCh5u8w2GRiXtwBu2cldUXRCgjp5ZkayX0m8vhRaBiZOf
aasvytVifogIltEjqVH2TkIaasgpfPNqok4rQmSnVIaDnNoXXe4w45JwkBXWoLPe
6n2YNuM8UQfIkTGvuBsG18jjwvY+8nuyNbe31O9gRToNigU1d7HceTBUYffJFNUq
1vbQHu6Vc2IE1R7M1MpknERkHkKJrMn/8WsQQqc21QAi5nSWs+Sz1PIJLmTvSBiu
pIChpSSe6lC1hmn7U36SFybpkf5kuMaxJ29AycyvnvXTGedX6eXeNnlBDT5HJU4S
waOnmQKKoCle/LRyr1RMDJCfiYn6xwkrPuLDSeDnkkIyS261LrAV68uRGEEIITjh
39NDj1f0F7Y0r3dafyJBPRXSVIUhA2tD/IMKVC/0fskUiN5OWhJXmaXiXbDcIN7n
3YQuHPiv9u2DWCafo67T3jtcbejKlAuGiwc6mS0nzcCOIEffKckuBs0yr4CN6Mt4
NPeOSGsSbKPPfBrStwH9ISTH6MNrRL1j24hYT4u0fZJuoDTE5mAMmEd86ogHKw1n
pRnLaycWi7ClERtAHuPn7f0lgHSccUHaHZrCpR9KLd+WAZlj5U+whwNxvLoiL2JL
DDHPSxDcAAnu7QyfJQyvL+CMbFJ6or92ps8kGGVgADZrxf7ghPLcfZNaR7M8AbHQ
UdGgHtJKzfc7fWDJc5OsCtle++LvRZ0uw/xwOGAoly0QPQhlbpRUUe9qH8GVxo6R
jk67T/HNLC4js54OekUNKleWZV/ywS3RmPFJA10k+GWruPxMbQuSsPag0K9s3DSD
oODkTsHJHeYPr9xEuMu0k7RQt2FQWdqO10cDL0dzEGFi7CkrEjZfn+BzJBdN7HNM
gW8cp1Xe60lGmEGTbTOLm6GfzhLoVLHcBVomQuKPbLphM4PA3GO4GXIK+HowYzu/
mvZjbIuwGYYJ674doavtVj3FdwQI0FsFUq+qGboEIzrKcPVKHdjsXTE83TsHMnZR
BSGm18+PfNKio9s3ZFlKRZbF13Qv0EwAW6yks/Nf+jHsa2amEqTdBSxjwNECQShd
knxUaYMfYeQMVMx5exqexy8e5FqIVLhPTYIAvAhZ1PAjoNHuzgpwCY6Uc7jTl3J5
MpXTXH8UpLixHVymaSnlOz+JkiMVR/tIksNaai6i77MEv4iw2DUMMaT9tRTdXDpl
TE/7UxbW+OZmP8XcDUXDPSLWUZK64BXoE81ypM1Xm/J8aF9p/Do7EetzWLo5Jcah
eouQd68RHHbtTixZZP6bSXwlzI2BoGchfbYZsRy1se+mYXVhB1lrBitroAmWBLDf
OmjofcJYWmuVlJYmrRQoseudkmd/zTmJcUVvgCDCMQbFZ1POGBzShh5SyVvrvyKh
3kCYX9VAiTssbwSXKJ4seoddftdBPpYovCOb9WtfrCA1+wMKeZvEucH7ajNaRnPb
OEXvwIyz61w2zOxWbnnK4/lbI0/wUFZINvOWmfwUryHENYbYN8lIVhuwyKzbAuF0
fhoBOuKn3RTHNonrRrXxf2xZvTkLfJB8MdHo4wgvP5VWAgo7XlF8sb3KJ0Sh7Gjp
kUQ5BN44k8t3M+7KocFKxYy3UlmWCtBagWbfvxFPctACiFFkxVrRNwYg1KRped/v
JuG++nMVSpY2buH3SKdVbTCRiSJ2rNWdUUF/BCUGQOQ5COADZE+kjz2LHkTYwFkg
0iDLVM4B8r27lm8ELEMwFyPugt+9c76A4BVA61YkzmOBur/e05AdyZVfoQ2mzUjQ
fskrdG07UkA6VS7LK8wzzoV9iPWJFWkwOfEYLF5Sp1BIS/sotvEjAOT1DzRtqU2Q
oIRLkEKXRXWOwU6TwBofZ+YYM3fRiOgQapl9xmPO1gsTSph5SVXavlOvFRFd97XK
KCYcZiYLqMiNdMhY9pborM6qEirN3dewg4RXUOZebKB3fN6WqxPnNIwjnf5oSGsh
gRmRbZFiBD16IZLCZU7kYg/CFjoVQFiqtkrodl4emUfM3GiidUteb4CIwzShZe2f
J7VuucnuuqtOt2AKB8H8ZIruBBJNTtNAaoahnOfXnXNYcZkGAqkiqrMYLPpKBpyr
aqzxCzXott226QRlcpeI8xqz2kTNWls5V3TEHjkf5EVm/LDX86QKLE+XugGOjD3q
G0y9B5LOes5p6VzcB9Fev/mt1nrbMZCEjERfJbuzGUrDUkhdlTqX0I8GjgQRA0a3
aqhMp5yB5Cfr7B5wkElZyfK58Cn+WvTl5oblETYLKf6JIqY0ENPNlvwxadWvqU4/
1mFlhvU1wYJe6NT4szW5+QHJ+1xlvwggH2Ns37dwqvhEkT9Q0V3z6rJs9bIQvs8l
tqD84SvNCREULH27GjGFa+lJ8jGc5/wFM9jj6+fr9bj+skdIlDeo9R0/6CxRENUB
SXWF/3kIZyk4TKG+5hqWXwb7LOR7i14us9znY9LkXgr72G/XZWloe3IvVb7qekNk
9A5usTeHk8T+wp/gLp99MvqUp8iPUhlynkQNu2vIarOmFe+1C0U7hqeIQowFI7ZG
BodSnRGedyTxTYJgjZfE1o1uh1kgtIyBtheeqNoxVja+vUfyoZTGg0ls3BoqCylf
JSCoT5f85KUmR2C8jk701Nu7Jmbu669N3aPsF+7Yo3VHiKNBUFPpl2sN0R3vXd+g
oSTUGOlXQhKxqtspJWCDgJfTpzbB5kgQ2/Tgi0NcyN9m83kFVdG98LUPlE232yWz
o53Cd4P9kGmqjbyvCF8ZxO2o7mXQhyEhxcNMm4mrz5eKFp6G4EtYtHSr3lKH0lAt
5t4/bw4PN5+Y6ZlLw+l4PgVyGj0KGT1qoxEbLxS+mxKncqeRmlVGHc5YrS3GMpLF
DVzD/0xoSWQ3wNseFPdRlHS48a1ejYxNKDFl3y3Eq/M8ZnMlBB6g9OYzn4Vvxbin
h/ePU70gbY+xdBndKEo1g+0JQdQoP9iKZo1cMW7rTMrwO/yFBgXkPTzYNRq6y2mZ
AKtrZZJRP9aLkPCgC+2ii180lXxqm6CME7WOsSoGKWari7Yki6U1huntmKMItJOB
/bKMnveMMV5Au583j3PQ5NHY0lk9brpV7sqGDizkX+1If++q8wYz2j/LI187GIfu
F3eIlAorklNXAeP48lSE31LYiVvb/vgqPcmSYCVYUh03OmANon5708Fd/cKQoXZ0
wM3MuIJdDJ2/VkXGaPTB7iYCht0FJA9gu7pshfS8MWuL4Fb9zGKIYgkwgQjmMDhI
+wNFT9n61/7GiX++C0pdQhCQUu0hzSF3tMEId6Ynm/hzfJpt4VGl1hqsjSvb/K9L
IhJPqTAhgHQfyzOAu84q9bm1qNj8TypDaCH4gjscOaP4VTOb3UJWJkKf41bJE1nP
4DifTNntbovXVg6As7lpW14MhTjljfO83bIXVkcqZcus8rmSn6/sdzOdu9gEkVFx
/SIc2CdDR9lD7+YW74NWysEkIAQBP/HsXPVwRXOlCLfNUpHVYaZNR1Yb1YINj9qw
oxq2cZ+iMggnZSR23Aaef4S14bR0rjr9u6ZYoMcsC5yaCo1/UeuQxH6CPuNMPpdF
7SXVoLdBUPaoq5QmuQt/lhZv+pCmxej2Oym8T823xXY7o+ElYP4FNEuwF/JQJbLs
lg5NQh24sMxipNRBKL9+VlNZmnJZaOT/0oyqZazE5kTeSVIrLt/PiRltbKtf3//u
9ZtzAzoJRXOUwUPH4HX4kEvwqvA8KeK9bJc6HULdny8jPEkdGYfezrr0sGJBmkzO
5UCo8PtRkSJTjntK63l/05wVyGJZNCBqVk8Xzxzr+MfmrfeAeHQB5EMEBLBlrGPU
AQpugQO6TvN/r6yyvjD0EL6Ghu4ZjaTs/o+E4GYds6c+NyNp5Wn0o+9Yz2yT6iw/
UAFif/avINWBMJo+oyde2kZaStjWyDcbM4mdIxV/Jdvvtxer4K8wUhAuAZLiJNMG
0TccAC3geFZIFJs3fvFXaYG/oNWWF7JltoVERdAK0m97b4prlwjV/OEneZQ+Njbf
S9TtmxN6nqLuZpnNkFv5YA4Xqhs2yr3lE8no1hO8Rp7bCQW0S+UXyHeOBiDh1wMz
DjqiP6skDIAu0ei8Iw+IGt3SLxXJ8z405ZIv9u4jmOHnwIvMTOWyd6sKL1rh48Gi
tqr/Ufmz5w/X1SDJBxLZu8xs5dDOQWuetLiCLApO6c84SdMgy9ovISBYgylXchwo
5Ya+j41bw9MizhKIYZsOYjQwbglaeI5pr2IEu6eIVkKN40Q1cBPDuklK8/jTvGcf
Wtr5sz1j/nlAHtG27gFmIwRcKFIgPtrhlVLsl1aTMEYYupJorCKApey7Y94VU/Yk
mfjS2zTiCQOyl7ANyshW0vm9QKufIfd0n82V6J1Ti7Odwf4IEBtltn+lBeChXpqR
rDLiocMbC0w+SsT32n4Q3iXUw57y2TwbM/A4p7kx8u6qy8ktoYrL5nRakYSZu3CF
k5pKnVVUFlqQCZYhATyXKNPs0rI+CLGLPdqUqDbyTuqUFKLCOtABZ75v8lglYA7l
J502kRdX6TQ7PloIw/vN9n+gVlNOLHiCMelbB4qpNlJIXhUD5rY6T8z9i0j7I0u5
KtzpPBD30Jep5f19Gjot129Zy5QiwPmaaufUuHok25M8UerbJ6q/A7jLaGwX4Ut4
sO2L+LbA4zxEDidAZDU7ETanNqyCk+T0g0J1xfEEjyxSy8e66dO/5R7QfQv5xxxI
nN4UkPKOf9kMw0lfQ4SYk8Q/IZSgA+qcSQJvJ/qXlv1ZH813lzhYhE/Qtrz2Gpca
Yy57QANgBWXPi+MGoVYy/NFItSrlACEixsaJysO0nAdKxWSdo0eobgTXDWPa5J3M
uuUwWM0B3zuBZh53izCGpA==
`protect END_PROTECTED
