`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+VhKk/ZWtaObm8M8WJSSptTcpTlj/3YTbSsEzczQxfC7CYIqIIHEfyu8zsemjq9E
6Slxfo86j8y6DjMT/vYMYV4lYnz5bky9qZv5xn9gwwyFweifXkd19RXBvnpPjvB5
gH51Z+Se2cYmOVYvroFvbzdGps96oDZ1FZFt1Id0C4wX4nqXlS89ONRe73Rps5Ow
ayBSr33AFiJXIlqIDjG/brezoLjw7Tx3kFdREM34sRsh7ltEgxL/Lb2HwZwL7Cb4
RDCoKYdJwFz5cLXUsgWzLjIamkPGpkGdKnS1sNenmEXnoIavML50x/kPO9/Pcsnk
eSHG90mrEr6Jq9fkQ23OonX5JkzZXojTB1cJUW6Wej+7InG9HEVuhLPFGG9Cx1FD
888mA/z1mGiOnlK5cxvGesuesM+lQ/GeRGL9OASWlUPmPM8UY2s59r0lzmlwqHoj
H0df8u3yAA3gA4KsQNwlWwLwR8nhmvN9JsFms/eU0ppjvPDP41JYXMUm6Ncez+YJ
`protect END_PROTECTED
