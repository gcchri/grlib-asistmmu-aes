`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PcctdmtsEEpiIzoQvLV2Nea1VAZOG/aCcSZLUCMqL7KhbJVrVezSyY7s2mnQW6Oi
a7PmUNxhtXncaxyLtMFbZhH7cXiNn+8wLG55I7sVrYSPiP+kdCDHsYIGI0pkJoCH
zdJPTpFJtm9YtBEe/vQlG9DHCQSbAqCJZpO3pGGMI9zi8F01jov9Q5QUnxlDtYWm
PPp99uTqCOVsSP5++iNKYpwzczuyVDKNqsSzqchgXMx6xdyoUNGJtW4MsRe/q1gD
PPl8fEwcBlEF4hRVHwU+ATFso42YVB9jzzrOM6kphFI=
`protect END_PROTECTED
