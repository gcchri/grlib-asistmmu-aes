`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zKhYRA+0yTYGChOEwG7M0jmdGZ/ESq6d8wFvPj99DTTw6eo5OXb0zBOIuUzeNGiS
DX3gm3ORTjlYlJ5plNnnlMt6Ga4M128g+cIGtB829210oO6nCU1OOMjtz4PFjcEJ
T0oXsckI2Pezrw9S/M0JeCB2iaQ4UzzvsuW4PxjYbRG/ywfpm5/u9w4L74gVK1D0
9qGSpiL1FRcR1pH89h4leETj2uTcDFaSwS9193VNfjy79Iqd5MxLdKMdSOhzSo/3
EI55utN+y7NEQvG4cekFaG2zi3ztr/etGTFz1+FYkdz21s+Cuf4rXqftSubULNLN
CHCE7dtQSKyy49idCgmECQfp7Kob267rp+RXldJT8Slaca4t8TZ0HTzte8C1hVzS
DRkbLrW+qDGZxMjS+HjltYYsv/VyPqInnE8mtXjgTnL9BtyTplpYRcKxBQhIuF2k
Ky0eH67zPnXmDvGk1c+Tl+qvoWqM2ENzJ7GWXfOui7Cx5Q8mNWEos54JmvhKoqu0
R3o44OniW0ZdU/+fWaS5TUsYK8Moag7oRqfHMk10k0hSQZDXRxz+urR2cuCriP9O
1uubsQOMhUhiTIywayV5xfAV/NgCMKOS8lidRG0d7NLzav4RbO2HzESFC+xPb/Bw
bVAxoXLn8WPx43gN1a8iwI6rhE1jUX3aF7xu0kx2+dLYfEttGiQGdgFC1Kkusfhs
bk2Nt15ACFtiPRmlWSdAfaz4t888ynSDN7vnh7zt6j7bm26SSj9jhYXMIq/y6Kj0
ugd/wzcYH7YcOjqVI1O6Jw==
`protect END_PROTECTED
