`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9JXXMqwC6m/zQ8CSt9AnIZBqDidcARYFYtR1MerhMyh0qLqk+KR5B0ojQPYkp86q
KMP1QyO4Ch6M456cJHTyqwgLTeawXyP4MEGd8k6oUtsrkOqtapDnLi5dxxqQ602e
grq8R6WlMnHdZDRDKrCMjPfPAgjsepQh+jxzN9lP3HQbtUUZleQxTTxOhC3UzuGe
/cO6qIQimGG4HnvhvyI9XojUtgKRptwvEmd58sgtF9jlHw10ryCk9DN5sBGv0ouo
lZOFPzVqXC58WjYTWZ/4S6ly8uMZBFFYH5jYTUVFr5jOmE9rsvfCSP3Zh/yH0MBG
vG8K9fgMh/a5FGQohhchniDpfmu7+EAl2r/33qmwKNMRkUUkRNQ6zzKx0DPT4+6A
0BSQyNXt07sbZRWWS6BdbA==
`protect END_PROTECTED
