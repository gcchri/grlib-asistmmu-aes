`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qb/IksfnzhuR2OIFVYBRk0RQGcqiu7nPUY4HS6KUCV6J4D+eowCW1CktiyWexhIF
h+ZbkBuqhTb9ZGHfPUwGFGJmg4C97nNpVO24m68WcU8HJO/iMKY9rghdFGcU1stC
TiPT0WERNUkkWkt6U2feVyFhUqIMaV8qU9L1eP5ls/XHGWmdIs7K1qmZNaN3g8BR
LKJBcqcT3TwH3QYAe1gwCJniW8ql242OVRF2j6tT2L9mblVMXmC7GoRjl5/WQ4E/
6hL1cIBKU4saop2AtbUChA4eVMRD5S3Q9FtAp3Sk+072p1yCiaCQ0xixdy7688nv
y8JfJWT44CqbGOzmaC6Pk1ob+ykpiS/BFnd9Nnaw6fl6gFl/25hdgIU9dX8x2Q36
dAwXI+4JISEICHUnvFBdip5xnRZZR1X/m2fd8I6nyJP8vmhsmZa2psREKP3eT+V3
taKrkrwXlX2Ti4N5pPGstRljUEu4l3qHd344AuIgkdH7uuMWLDYkDYq0/HfAImYh
KjzHs1uz65Fj2n+nN8ECATNimhofMIoTV0In/+YD7EFomhVipfIqw1aiE454CN6w
iIqs1fQbW9ZJWMCWvk/D62mfuN8ICkSEkD+aYjHELUugSo1x9hFvg4JFFKIkJQLj
n1gXhGp9z/wrdlJrX/LT/YXkr5JyKkDf3FliEBe63psl5onbZFCagAp3TUlmXWMo
lmyjdawIwZVyqyx+4mg2pzQu1gjL7OzElWQVSTSwBuzNffEA3W/RjSlEzva0A2dz
5FT4LM2cbt8TYMK+x99xMcZ5ZQWiNu+6RxjPmc9QxusmeoK7vq0885L2Zuwb8GYB
sJ5P+LjWAv5pvKy3qC1PCvlt7lL8Qb1SSCy02s1h2p9nocYcoi3AAYbshlUYr7HG
HG0P+OcsyumtBlpjdEgXpgWTL9r0MYDH+yUEl9fozQ1sq1hT38EmTYapXMljZuy6
am956K4YgpxUIgRXu/StwzWbMn4I0jilL/IpCeqbmJ7Al3FKi+WOBLyUvfMj7ntZ
LAmku3UaI13jqSL4xs2VoLR/juK1s4/KlReAevwJniKE3gYK7F6Kwx7hACgDlxCa
EhLweVKS7ldOSPLmi9UOyt15sWzihqPv4pE5Y0l0ZXuUnjp/vuPbJVkOEihNX4ui
X8vBT2u1MuyZvsKrTSE/PzoR7Ye0Hv5HTJ6GQ56RSehOADM8xsatIWs6VzDZqqw0
qieZwhN2Nxk0yCCExy7QoIJESQFQ/8jMqHRRd5CrW/vYiLoxpPvLx/O6fOvXCu1p
x/4HA3QsKNbvqfIx59xl7w==
`protect END_PROTECTED
