`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gmOVqjBapFQEu2921kN/ORXHGm1wF1/g76e0Gc1TkzBJxrKHBd5WMAfCzb05pVlZ
BST896Wys138fCmdJto5idPdo8zfagYJkk88kbRTwjtaXO++gLWc7VtAZUIcRqA+
4VTIK2nmQpHougpl60ogrb+U6KtVnbHQGh3KbQL/4KkMgs1UUzWqDoFY3AU/BS6E
en8wqASgKnTJns6ugfeSfXkZc3VY3GJGAorfK2GcPqRVgLINTLZnbxjtnfJs7Vvl
bjiS+vM7zmkvxNhgg7pUjqPZMghkDILUEv3Si9nB6Ep/7gYLBB7cF6mZUiQXqi4N
zKQuq8WKTeIDBZKdSxWnAx16F1VHx2Gkm8wnhi4FWRexZvtg6XgDBl4s/slvsr0T
3aFSPGqJE+nKxoJIJ9Q2oEHWQUUgpZf3JBrqS9rQpAmHXZz0gvWtF4JA4gqVrx32
C/8CSiMKBDwA27l/rPPM6Lnkl/xdOdHeUJnk6zS/QSCwcXkNpqNIgNmkBN6skdrX
9WlSt7sS0u4m2oMbwAmHJ3Oop3i1WH40G/zGvy8GF1dqqjqPuLB4MgkaMpzBSom6
0URtLB6tBTX6brHWv5S3pqukNTRf+asKuouwDv+MwuKapSdyiI9MUUgyIbf9lEG0
6GqWMynKjrMkGmQkltO734ab9SIF04XyXy1csuGVOllMt/wnMIdi5qZ+JBY2OUnn
DVsGzMH3SPAjTPEvzbD6H+AkUteZbVT7BdvLlgMyxCl+qPJiFAm7jezVTvEhdade
+AepEHqVVhFwmPCHJ4EPyB4mNFuiqmKXvoh7KoPAOFHJCc7L/Zuls9yJQhi4io5x
dhE7I6wsbGJj2SL2B6GyFE+aM2JiU/+wEJyQ58REmQ3FLVQJ4x31zMd9v+bKjhxh
qqiLgNad+KhmGCzFxjuOiUf9lhj9nlSSconV48T7+9bkssJYtQO1ff8v6RGozqzO
kwj/rZ/HjKXdNBKJ1YD2rMEZ9xyFB5rpIDQ1rQ7jgcGCLept15TtsjttEMgc+GBb
iup8rUD90tDh8OHMAYc3Cga55zb2alD1apdv1NVXL+mPWy7N9GyGXCikwy9Busxo
m+DJmsmL2IVs3SObU0Ih62468Tt2/qrk4wm7wGmYZlJRmQnrI5pQZsWwqD+OhvO+
+hoQr3DSAsbk0Me03osuZ0v7YN0JF3RyU1CBsCDik8nZABRODw348NeHD/9IHHF5
ET047tk4P89J6w8IrS3WHa4qEH6L82Ng2FW3GUeGKl5PvBhN6suFRGyc2lN7MYti
Yc/WcGxufoZs7MuFD5Cl2ON/UAIvkUDi4+pFYFn0I3sJqX0/LWjy1byoWLMjb784
hz/d5d3xnpYAJFyBia9apIXUKMhxjI348dPaecTNpfh6gqGNss3BEPCaF7H8dIqd
SOtBoyFe0YI1KOiw6E0ROBU8oocE0GrQYUoiPqz2O7l/R6JbDXaWCzjvM2fL6HVx
wAo9nJhLrF33g41yRbw8g8k7TOvdkGnzec2gzdItg4R/4pGctnOsYZvGlKKocP+2
X66z15R4IfptI90B5/RfYFh2wVw56avnX2VFBsCNDGHwaR2P6B3xEshtDduRjLoO
sQC5DFYaT224IOaZ/W9eswmmLU8EFuorzu8qRozugpMcwvi+51YtVT8BCBkz7YSl
p+ozSeIHDjW+P4SPpkl1YPy2VRCQYvOEpJEt81pigUoJa8yJEZ+LuEdK26n0WhcG
v0Y5ccaASY5vly/WMfYPVEF+EbpRDZI60lV2/DpRZPf6tdQkkSkiFa5z1VKn0hov
X+OfDcA10nGxwHD9bwT8gABa+8NlOxas7J6N0hoMrTkdjjGUt6JjY0Kl6SmmFqBj
t1M970BZl1ETEFA0CcQG+R59os2EXD7KakXE9XaKV0EDQZqLeAoLPlb7EooWjKcF
GDXwYW4Lwbuu0G5H4mpHk5AbMH4uiKhlXi8jG7phncUSAz7UUd7lECH2nAYXDCnc
IkZB8uvJfRErghY+XbAAh+wXcuv7ckzmGaLepsS5RnQbfNB39mJhGjjp7JDON2km
CQHsM0iRyE2Rc9j4YzBKD40363LaWXISWTNHnFeUs5k+PEmtMeq0ylf+Es4ZphKJ
5AlfCrl2CoRjHBlfzZteEgrojIM6MAG74rbiE2X9Lc+HNYs5HSL9IARLQtVj+gck
k8WIHFeTXL4A/5mvlRFy9FXhfZckBi6WL5G8eknWqhJqhS7zl9LB1QirB17G4wIG
JsCCajcYBqSaLqoQ9TF9/PdOrjnfifzJxCR/77Xy04h4dr7FVPvsDkzl54qakV1Y
EWViDW46Fezv1EhAFPmwMBRSsXacwUh9fNelz0FRAIkOUBZDvvuKhUTDt9UQ5GIM
Nftx9pJl1Q5wlKfYM39qcdtuPb/Vj4yXuavkXm9cmWQrsqBBnIEljiXw9SSkJ4Y/
owZSBVDtY1q0n8J+OO4yeaWm8JnxdiZFYznaf8vR0y1OWBuyvYkMSyNAGal/F8M3
GPHrqefGzDKdmYacgVvlgcOymII91BVyuAFRUS/jh47oKNsGbjrpHYwdkChxMKaY
qsj+W/BIqzYniRIzEH2GP6UEs2zv6Vv5Qex1Omk/u98BzC3+DCRlFzwVqOwXZ78g
w0o0eNkJVUYRYK95/t1Ku5psxNEDkbdHtDRc6vDIXzdUyuhVgI2ThdI6XhgnUZYm
GWXKJ+0SlsBRwARoHmWbeAU1LAJ8i/7/TRYwqaxwN9IBiuWHPqtaEGQ2KNBMeMbZ
98aS8d8AMdfcTgREBOJhDsJv8TJ7zPHV1Vl83sFTbbm4cNRFQrgy7ZmoQjKJUKQx
QPL01t6HDw3we77jac1hIs/JCxJRZhDnl2ab4kPsuusY5EKsAAIe9tHeU/lI+Ih4
95pwsbnp+Jy63P0mbpDb1ssmM0sQW2Uj9JMZUj3CsfqXYYllgW9JQKnWILRybQsP
pnWi/gjkMYgfN6eVFpjEpJs+kRIE1ehHugNQhjnPcBwom7QzNtVcA96dALkXL8ug
0rIFy/XwD+aiyFZ5PFf4Lw8AhLI82IG55uCZMWOLM177PzliEFRHIO/5zfHRvDGC
aF03ARqMvCxHM5KyRf/1s8CZbWSXNufKxEwLmtEdpwyx12oFci2tiFVRWlB58p9/
f6axpi+vtKTkMrrsFU6ocqaWogfFNxAjIfUq9fLNGDp7dO/A6nMPurV9Zizhqt1a
nJE36qfDVi5zUiPUdsKEPi6TfwBtUQIcp3W0I/Sk9213xT94eBgfGTUokIG5BezS
B1D1UCVGuaBEr5T9yglz+t4ntqb3s5fpZNcacxPV7AyQ2C0dTQ/sN2NNqBQans6F
aYPSgZwI37I+hHKP5IxvLjrTFnOZ6L9Ee+/gSPSzkWJiclLpkKal/A4qrILJZy1n
AXQoCyDADusnI8ba9zwIJfY9l7KgBeP8I9LPfWLVUq6sQTZ5yrE4b0EXU3W8gOLQ
C0CWyB6FfLxuMbMZkyPSJiRWE0ny5vwcmLk+Kkd8VORPfEuYYkOyI+0eEa6AGSaL
0ePvwhzSsBydBVXHpConpSFilD47962IRr0e39v+BNA4hETuukEtYQwffdqlXoQB
qQ5s1uIA8unCdsm+ceiOPz+EbvDw3bqfqEbOFe+DcwNVAkF6uYtopSE8dPnrpJFD
LV/PeIX3x6DnXPtnOaVs6eYG8BEvA7qLOm4e98lstxbAEl/6OfBoA5n6MfNzp5bB
T6A6V9w5tyk1M8NNUK1ziJP82CT9+nIhlLV9d/ygG9ZItxfD6gV66GY/V4FxT3Fl
RPOZ4toSS/I3i0z2jaPX8H252y9DCvHfMOD4v6TjN9FigpXJEQWtQJ2dkFZPMidM
PZlSGxfxjlgcBOqMoNV8d7JWH9wvwglkyddpZD11rixp+8LQg1/PtmewqgHZvlKR
5JehS0oZL1hnlOKCWZMzYszoeolqirANJ2A60gufC4S6nxEH/VfsAR5vx+tST4wD
GE/I5ygh71E3RtMsRihzCLGBnNEHBUaPZQsEl0YTChprRhZtlBAffAp0JHyDIE8T
iPOR+CovECXngIrcsua7rU93AlGspfnxL+eEayWifLYvgCtSgdz1HMnhPcKQPa41
SFVmIIdub32TWCzur1FCYjnsjrpD2CBQg17kDdi5/97jdADNSXoMJYKw6c+qr/24
oVk3vYqb9gIaArRw1FzspgrHtB5XkLgLu/UJKTa9bBouksHb35vzkk5Sezu4DgDo
5aPvFOd0nLGhCGEfncaFSSetYn1q+L2Hg2rEr3ZTGCkqC/njL2+mJv9j30bE9lUp
BMDLtVHhW1ljgTgsc4kHuaVrXbiDbvDz3vqKV8Efix0gURwTOkpGbNkg+NaOWh/H
HDEPGXqFrlfcBdG0P0XtD6gUtHQw+IMKRcG80CuhdnqNIb9sn30xMHk70aCQlsb4
n/rz56x5xWdQssdv0AHBuw==
`protect END_PROTECTED
