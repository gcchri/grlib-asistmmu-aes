`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g3pjO1jaEbAnj8DjRP7fVRkgK5Kri2XKdPEmcUhnHX+FdlW8hFv4T97VtwMZyzYP
ehByFdNGigkeLcJZ0T+aJWFF0vhUlmQaiLf0WK4rSyg1FzDs8uIyoA6GLYnbmUK/
kH6eJAKlvZNBMJFSokyVS1dOM8IuSlXx259HHLNvfCTBX/Y7/9Gdr5nYUAnSID8Y
cgALT4sztLI38z5FGQ1LsPn588zn1OXQkMb6kOx3M8XKI1A32lUDiWNVpI7Oleck
Pdkf/Bxk8pIDyRqF6eHpzg==
`protect END_PROTECTED
