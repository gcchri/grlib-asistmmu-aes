`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PHEIuW3bj4ml167cbqrbN06iRpozrauIOg/Le6KVLLeHRIcErZCEBuQlGA9dBXXd
HnTnGE0pfzgz8rD6AbaHtbQMhXiXMgzXApqafOef9Gl0ILzS9ta7D24gHJMdx/xo
x9SeESsSkvexzf/HnB9U9lut4fx/pSWvF0Khshun9bIwZoZtLq54QL9dI3Euv4sp
eCqR1jGcfTaeJoN0AxDiIQ45NyPU6z33yYV1eCgjA2tWbbf3mOwszOlA1iFs7utH
u1h72FhbVOyccytVuIqKAdUv7BZAXsHd8SbazB0CI7YtJ5pu1r64qWTsAKApdsKe
Ppf1/7vqxiJ2fZOtOG9CcF0VtK2oRdwAJumAMWMyMWo9jmFfgJ5RyquuovzwRT/i
iyVItDJ88U7CsjKeDNzuU5dF9WmlJd8RdW7uwwhKak+8B3ShQV811anSYWqvzoXW
9kHlliTPCDHTejGxHG/Kx6jfOnxy+t00JERE38DIia4ABs/5SIoKNpLGbxOK3KXx
0VIpzn8Au3lWkTFvEm6pDm9OE/LBjGk0NukN+/N08QJY36N0tI5VJreLSGnNkAX4
79RGRKJAipSN/vc3Js84kfaUFm8k5j+tHicwmHaypPH9PvplWgIx0zOG+Nmst+7p
99EbJqAgJngWaYX4NPc4xVZ1TPWhPzwjivYnQdy4avEFsK3hbAMUdyjkmLZvsGVS
`protect END_PROTECTED
