`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JYqgd7RhG2WLN+uVviSDnnqr536gUtctWp2Qd9aQhOROH0SU8Qe2nLTZM+/JbO6z
ZebmFsCIIETs18jNoZbBtkrB1Qka6IP0k8YJcb38Or3xKpZq5igHm+XAgqci8nTe
HIzi0w7bbjbSH61YvxNGqxwq6/HkHVVg3gV46jgucN+Uitp40GNoflongWWFKCL8
NVsSBWD1O0y60qJLQyHQ2FpQtiDNzFL6XJO85U/O0IulQp7L8IYR+ie1lEvCmh6D
aXfd6DC3FbJEgYQ6Wd9dhOp6a/Hweqaa7erK3k0JcC4bwtJL+BzD0BE3oXGApIPi
NTJlnbygr+Smlp3JhrSHEuhWLTb8xbbrakK3IzRqc3wFkP/Bcl8ECMDERLdLHqCA
DWQMrlnsQQkiQoF9X++J6DEJvpghLDyoAvXOe+pwRDt5kzkmIxdSFBJ2n6HNSTkH
/zeR5lSu76OwMU0wPlLx9BsOxj/fHgXWbK0SOdd9MuWJNOSxweaqmQty6btW1l5Q
g9zAZklFM/dPU3NO+eJNqw==
`protect END_PROTECTED
