`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9yYwe72zj9JvKerCLLsAK1owkper5Kk+/JZrGvNxtUlByi/8qCteFDJ7Qm3IZbQP
QaOa4Cz8ON5DitA8Dpj75AgXhTnryqu4vQPpHjhKovZKt2dt3R/JUufs4La3h/xp
SjAU2AOnyPi3hdmQBOcWPpRs/ZgHXKX/FWb0G8zutO4kXntcC/iTthXWR65s4nVg
nDqAWJOjWd57wZ+EcZw3h/V/nZB3ZZj3IPvPh7e6TvWysEQpobPlIcBc00LXEEps
EfJpEnY095jzwmncmE3vZzBz1pcT9Ecg/2FJx5KR0RHqxmEIK+BtLYbby/yT4xZH
fQGeMtb34tqv6TI/+FDA7WBfNi75OVgEKFSwEPjOIcsSCdc4fpuEmLmCwli9lkvJ
qJmkaImlJ4QABRpLTX8FTCgLy5lESyZo2tPuZ9hoyZk=
`protect END_PROTECTED
