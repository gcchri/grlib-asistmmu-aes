`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P2PpH4iuutWnM74peCpuGryg+8pJz7FUsfY+S+379NjOoVw4vI8r3nBO+uazfmbO
6YFE85Rs2/CM7s9u6B/17tthyhwJIZrI0zRJxG2yMswVadOXzKb7+YbZ9ahJcywT
4NSf8jwyPxU/iOeiTRgLOlLt/YysOXK4LnUeyV0xDika12Pkgso5WjjlK3u+PFQt
NgmA16mD8ah1wqpGKL1O+pVn4PoXP3qqgWhpAFZO6NI9W5SxvW7rh+68lpPYGqSo
VJlkL3B7zlrxj3W1xW+N+1f9ZmBM8+LFmBnckuyfcMNIO7Pw2K+f46n5jsC0RCPP
I9KL+OKrrKI33utsDlX5E+kvqcfkyP7gWVQa+HU8flr4SX/pUY4s6B/QXCGDBQu8
tRa4iTn3vMKttM84rvPYRU3lW34/TvY6mq3jm8EV1wXHS1fpz+LWtVRRtn0fQwSN
yOWGAQcv/qycz8VrqFRx7EKg3GzCAxMFgfaQ2ZvdAeR0ePVQ81hbvDYU5OhBGjhk
sxKGUbh2d7M2fb7+/5hKwsu6tOAvRhh4C2xZ4z1t9kkWN+3G2kBq7UKoKUEPMP3p
kaqZ7bTy2eLtKxT5OzGCBYHo3ul3gsnX1hru/TjgvWdfGWOO7uhef/Nfa0jWkK3w
MK4LgjqAuppnSJzRY6jCCVf59FdacqMVZHPjMs4UK50uSeZe1uQlwF6cjgYGVQaE
H09BTnlF3+mL3PYgfJL3kX3pDXqdC7OZ3iAFmP3y/tO3ASUNvfiyomJSWpG+Zfaz
eL+dZ7wehDTlCHuPgKnxuU2kgk3POriu/G1G02mpHzppEeiN0SBQoWNBhtckHzBY
V3iy4WNpJS1z8ff/LZMdIusBWy68XfCblITkAeOJFjR8NPeQqnBOVhS2Vky1cuTc
+ReE5zRtcJjrmhvcVMz6+g==
`protect END_PROTECTED
