`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aG41OOqMQseA8759en3p0dWMMtaRGD2JT2utmWuPTyo6cczC+pICfjYuR5b37JOT
itoZU/L+LJzSYKJfatnW9tkQpCojvDUk2nyp/slUw1KFsntsUcVCQLRAMSgN8fFk
2ZAgfv8+UOPGtj8RA6HUC6imGcomNilQ232LmpltUw69BFUy6rrSJ/mkBYlj2xQV
t8vaq5CVkzMTwdSuifR+4H85GAhBgijltn6UXgCzwWVSmLnsCDiF7lzDW2UauIaU
TqrSbk4uyqhvXFxy8czEDb0OzG2qw4y1kDJDyn0YKBcIA1hcifZzx+7mb8+iT/Hz
SXT9S+ASOyd+YLGRxJxh3a39LCKFfnzd9txv7+8XLy5Ni/NYRkSGU+s5ej3C0YuP
LR2EfaAASE+8wbNh56W33NHf0WNCy+ISnbZ7THD3+Ls=
`protect END_PROTECTED
