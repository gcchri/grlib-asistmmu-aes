`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lIxtuC1rBmJ6wv0ZYtflCmxArv5dBlvjmZeFrb4xBZ42BVMcDKdht7rsH+O5DRN9
4UeBsMtFhbOvCeoySAVRkWaeSTFlv8FvG2Vlq48sMgUriwXCZbK9eEUEW0AHxwhT
oZRE8RK/zefAvfDxKS9mpUiPGczKLogi80l0cTgj4oqtQu7+xP0XOj6GfBNM43xt
cHxNXW8vVcPnVJX0JElc2TJ35L+pK70gS+qRLl1+7rh8rXKS1nAfSBXRZi5xyRfY
yB4famTpcjz+/97Y7SIEqtMrScbp8o8ggAZxzhNxldnI6HP1+SjWM0YEGGrYHWBc
GihhBvjKyyPQnn9MoY9YDA==
`protect END_PROTECTED
