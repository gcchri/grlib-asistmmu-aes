`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YGwwBFWL2K2hoWAn03U5b//lFg8pfBMA8bZh/sfQqENadNchcpz2hAhyak/bbh85
kpVKpzStk7yRQDaZRXtdEPZ3MDU0ut0zZcHvx+zPaXkxj59YQzUq8nH3KU1UdG2O
5KgKiB8tZ9lhdPyG1aAv5U99zDxcbAvgY95M5dJUDbZlC7//U2PwXC8Gwi+Ny1uw
ra5jfYNpiDT22hqcTGzy+Vcda0d19SB0dp5ymntGHEapFUMIBWqe4OOjuPqOol5x
hjr+AJRvz2c19442U/Oo8Vt1U0ROy+uvhkCxKiZOhEvLsxzpJdCHRhO+ld+GQwzh
jEovm98f+gDrrhe0GX48qipMbBFW00pOJJU0IOkLTwmhziwxG8Ryw28LB3mbVA0W
`protect END_PROTECTED
