`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FmYeETc76PnvxGbW8Dve9XGoO7tC9cvUe2qr9VOp+qbMsDH78DB4XEvHwpw51az/
i9VJWFkW3l8pHC6ORy0eyXNYw4j+yWl6VDxYacnrwuyO2aKs1BhpaBsepcqV4I0v
OkS8yN27MtJhCjsgx4NOI3EOL52/rYoltv1qMU0suEJucy9dDWYue7Dkfxuv4sLR
LATF5GlIOI7H9Lqjy5g1N74rO54euU19iiTvy+5pNz3grfHxKb3+wNeD6YJrBY6P
lY8NK+pL7e0VmnMD920yzYdFNbqMSLlx0YMtRkrFRVQDZ2pFIowGlA8IOsvKeARy
MHb66ZUBlCiooeSP4g3qOivyC6thEFkSsTFgRH88n8VkBikJRN6ghkY+lHG1TqwE
z7tKfULcL/wmB0Xp1+6B7G/JxeI3Ilx4u0zbS1onxsCH6A6H6wRAsnV5TNx/aYfb
Kw9jUArpyBtmlEjF5xZe2NVhJjisE/rvA5tekJoLH/AQ/F/m+ZA2pfz8tM/yiPBL
06cEYL+tB0MZmGLKS9oxmKGD9DTE2n50Iqza/j5DETg=
`protect END_PROTECTED
