`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fjdy9lDv14iHppGHHY+a2DNgDUOIjShvLgA238gk/UTaXXyNI9bigCsD1RY6lMSk
lIPDkVKjXU4C/Y7f16iHBRwo2OMvutqT6nMy3lmUyvbN5F5XCIw7rdlERDw0uKQV
hwqhj996zsJln1GYEMkqvW/ZJa929O0UiSvfXEurwI8lHY6WRphZZM/nTnITcuNa
0OXgbu6NSpGQoH/UQGVsindc0+1eA6mN3PKsdFQLYOya2fgWtsf5btrQFAZX/1Pk
wmIe6VsmQQXofTXMd3HZM+41hQ7P6T+E+kiTtg0FH1WlZ5/D8wjiT/o9zR0zQJUY
VBKC4DvGZQjfCMPsrZARFBG3ftv/rOrdll/3DDOhHszXEbXzN0/nJNN2T4GV/rNH
`protect END_PROTECTED
