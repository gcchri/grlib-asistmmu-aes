`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w3umWPQrBoFJ8KtcO/gVvEfp2gWFNGMJAIieKMQeVEbFAmGE10tckqPsEYqlxLqy
Ehefjur5R75Jv6UveKQs0yJWitCyuMl/LIpEuZblGF5OEZdjTvm+No+Zcj+HIARH
skXA9FTJAlWqzuw3wPr7cu0yn/UdTXRGeuZPhCQL2r1qT+aZELhVZchLHIhIfytH
N743S3CEXL0gVODzBitvqp9U1IU2nhp7j0HNhSBi660/+rwgM0mERzBw65apwL8j
jJHUAn1gDNSSJ1DW65dRCTbXRCg0XtY55+8hx5zWkEsvwiCOWqqj8ixg9M4T00A8
hl2ALy+KugIIo2i9q8YXl95uEYhOPdnBiwmXpJszzwR/IMyygTsmxWATFYrxE136
YOE0iWbZI/FoOcxojcdWuIQnRpOKSV+GRb+Kgg4Ahs4=
`protect END_PROTECTED
