`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m+dojiuCCfM6TofxZHF9wamGYQDO9qyWSuvlKdOIYAUbHxASTQvGWDIYyfbjfUnX
lEXrzAqQIrcxXILwPfsiPWHx2Zl38bRbMLC6D3y+kyw71SwbbMYH8b6AuaA3dJ/q
BbOG6WnqCRIOhisAu4zvyOjghGe0J/BDCXRF55BOaw3gEvzQN//oJm44FPPQrpPE
k6s7DGUnJfjEarHProJmvei3Xc4p2zbNRH0T20+b3d9cuAhLzTSb1bC6hOSjGhVW
/fMriZaOhi12Ic6uR+Y1eS2WAIRgVpxT9qgkbxPNQBSzeSJrk3Yv8NfnCKiEd3qR
`protect END_PROTECTED
