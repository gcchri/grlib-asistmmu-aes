`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R1EjfKj05WFZutVmsaat2s5rPAA5O0sincUSqeW99eOUBsqTq/Uz4rItps4Am0ZM
zaXZHgsDQBQxpWILEoaxTTjKYhPaGt8z3FCsoKsizuQh3gCxGCUcHaChW4aDC3ld
G9TR/U6P4Ws2LZ5xudZGpGMzO09CUzIeDqlnA+5dFKVfTm4lVfRY/GiLmJ11/Z+B
VUGKU4CS2Tn6YMgM0aG1iow/ZtvaUOLjhsV4gPsxXz9UnYqZmYg6FNxtfU3i2Ckq
hZ1fqRU9Ih5Fff460QrYP55qis7SlDCXt/xkWRv1rugzFf1sLow+EtZ+r8Y3bu5Y
KTDtzqRyBjjq7H2S71ZRIBeyovgOCYaC60pKNj4s+f3EkbWmNx0ljV37vDeZhUhN
W407goFwu2HGPVD0fehHcAbxbXTmtSYftkJBjd7Bvt8mxos5z95sDEnbGq92lI+B
6uJWry+V2ptFgAFkkDgh/ULSc7TLrRQCF9Dy4rorWtL5IxrbWWoNhSiffGyFYqll
pSTVGb61eNJgGTokdY841lxJS4tcOiOmxThnOmTlUxFfVVrXI8oj9u/yrXJ2s1PV
ZRiu/GnWPPXG6muPaGozUNht9kuldpzMQ2L1E4BPeXSgJvPySx6/5lJjoi0tvDyr
cawn+n2CF/3/fCdKnzSusJkh/Jpitl1ZvgIWRUP5POoUgr36qg9o93zmo1ZmndVR
iT5Ab7y66vVpHFB185SqoIXNGa+PtgsPgCUnzuKCaHUy2D24s/7QBUovql7joo32
SX34jEd13gcxrW5aJaLRUWhghPjLzVW4KPdCULEso43qwqcE/y2uFl7AC14RuvzF
VemHfQ34BLS655TnBW+c38r18als1xA6huXt+o4hIal7qOMyktx56g0limT1ibkQ
oY9blcGJ8AJH8dEZoyLaMEFXiGlApUKLoWJF2nBqnoAYKrLwv+Bd1IyRHv524JRX
tEnlr+ZI2juwDhPIrEowK7vcIJo7iZXAE2KuXU9ofqXSDThwXBBRB+tZzprd9mT4
lPUz25dAhE30iArrnr5HgQqOGuhTM9f5lflp3zmb8GQfF39N9NqH/++zG8CPRW5b
rIqo6WYMW/PpmVB9SE7fu1FDXmQqdKMc3YjCLeUSWCabaNhdk53I7hYm7IMl3p6J
Ar+gUiu62/TBEzdAjgg3Kbiloi3/fN0KlMD13LgtRwvYMv1YIAM7+388IuuF8B08
8TthmJ1zxPiFTzYjhWtxnAkZeyiEFG7CASNchr2LckGclj26sEm2Ie4Qkz7zr2I7
CDJQI+zObR9lEpJ6grjTugPlGgzdM9DXu/UUgvf4WY3/EiTi7fK3hN95KYyyduoN
XcwzZPxAinLv7WUb7Xm0Wyj4JRLoOAM0kPYv4LSiZJtVYcXZf3FQzahkzzD/F8O8
vz0eK6zckviQpURuL9tGkU3ABY96LI8OwcYoxQbelfDxO1PQttU/quSv2bYhZulc
KsbGuprbM8gX1mid1T+alkId345ONwsKxKMiR5N5hc2S2C+PmsEEvMIhraqy8pJZ
9vWYhwfaYuVrE3bAKMV69i56R/cIVGVnjaywJpNJ5ZYaY99DgpnF9lL7Hzh6Exos
3p2w5B0cpDcQ0cHLWqBA0uUkuXqdjr2d9CYI82op2SSOBs/upVVH3Is4VKqhDHLi
5CX4JLMlk1sUMK/Rjbz3lMYrOz9Z2JJIL3d0LOQtnmdDyE9ScUA7u03mq0IbSLRL
qSVXuZZnadYfk1mJiNDKSe1Ra1or35HUz8jMg3CDS49olkePbeeJV6RmkbuItD8R
MQEdatrwFzkfp1D5NceDj+324OVLn8kFEbS+bHJZwNW1ntin+nz3zMTGNmhuwy51
mLFZrDUG5lHdPv4VEYyq1jsuZPZLnH6eP3ChybeLH/g800duYQy5Hx7DsZB6lFCM
uFv9AArfqnmOTcxKje/K26KsQDrSxPUO0kApFJkQ2PTvLXysi4yGhquhFs7Dylkj
iwu/b8E5y19T6luKefGJvXY5DTMbiwZt0nrVQ8tx8Q9f3Zt3ZwMnIeCp/aIGiLh8
sII/vu2fCHrNm12m0rNv8NzN0RkgqjHMbBd+KyUySPeGQ13afrPgXSSqOVnRQUEe
2reiq3kpTLaGWR9JEz2OmOnJUm4uY2mrIbFBKdjDKpz6Iv2UgqnZ/pSbq7Itb0KY
cBSZ8xYSJ4As7iDr7kRN2BiZwKbUnvATaU3QMILQ2BXNWYFSe6is3zgMreVbqS8+
rT9eyOuLe0B5LkT7cP7At0okpG90+JJyp/mh0YLSR+w=
`protect END_PROTECTED
