`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LBN/aX5omcAlx/ZjdSuyMy2kmoLQh3NLYUsyREuErezM1ZeWZs8myhUkCkUFx7Js
+CE/dRXjVbVNf3YQsNzxRPCTuHBkcYveu66ZIFxmTkbb70fBAYhYYSzCuRDslJdn
cWWpNDGc/v1FT3io1fFdLHFHLeh0ZL82v3iqAhURqZJlhXTDVjbGn078b6knTf5+
uy/aLJiOA2W0OgR4CQQfN0AnfeqZxsQHmm44bNchxAU+TGe6dKL8aP6yCWFbJcTs
HHZAWHaGzhR3YeYO9qtByPiKpZm5gur2zOJ0i+gbST6XeOmZL0y8JnNfvVHUu1Ny
DLdY/cN0FazM18DuR0NPKw==
`protect END_PROTECTED
