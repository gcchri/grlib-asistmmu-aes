`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oAoqIFUg8v2e5Oc75nwQYKrpRYXEsKEOTqgM+HUO8JbkDERxvoVbzRqbK9mEe+Db
4RGdPNqM6n5XfpEZT2uUJPjEhdGRU+RgsQDkJ3nhWE3ZXuvz3A6K1wSI3G3N4Or0
B9sn2RiCPTDhTQAo7WUFj+QYHZOBvnWC5NbrW1oLwbwCqT2CKUWRAgZ24NkQtU2C
LV+C6xG/VGlCwkW+KjnXJ7ZjATOfXTqqWm/f8azmA8/+4J1OKEscjxsenjv/pglO
a2Izk0XWMQA2WmDfd5vac78WGO6hsUO4XG08P+ax1xgOK+46ZcNImrA5R26iW5xu
CqVuVHmKFtxaSoFA/eeAY+nzj8OOk0MOCm8U+FhQ1lNHUe9cI/38SC2FuykHWLvx
gMy97u8lhnybkY5VaC5qy0yqXeJDKLICCbnt8hSWOBUA5e7us8B5MYg2vmj9x+RV
uw5vw43WtciXbv4zSXYf1FkOIUmdAa8KGDZkITVdvfwto1Th0jwHgzj3+jEmEcnD
jin1nkUTcA2spDZ+zPSf2c5+mETYvo/rf3j3E8Y3XPrr2FXjNsjzcK4lFKeMjo8H
0L/sOD0KAW1HBkA0jSPMYuk2W8CtTgRt/Gp/N2/TqAU470Kk8AD3ga324pYbWqLB
El+It1j2l+PMnyLR2MISSde/0Okwrlr08OgUEquRhNGwQ+v3FCYBYOPPPdf+1qXM
0Seycg58GXTT08nbl37Ea8XDSlFR3CjjcMGPRKUOSRIgeqigcTbF9JEUMwn58ViS
tAmX/pUZg+h6CQkmIlRE+l43l4XuiEYCh/ZA0B3QCslogw5znU6lp1Dr18D5aj1Y
WhD5bA6/PEKRC93I/JB2vO899/Lzx+cKRDEiABZtsvRu+9svi/cElkaa0VpLnMT7
SoyTDNOKAxqdgkFbefQLxNnSgHbFC5btsPh6Y1YzzQBZV1seKpcY1LR4r/br18BO
mt7DobHBnlXPqtmLWIc9XAmkMZzwXmNEce/jzy64aazRJMxEMqkUmYbW29bJW/gx
2hrMEEXtZndMl65eNea7PUsjFUURLNibGH2cToH3UjtduEZDXiy57G0Kn2lJikNe
khIV2BHfaHKIMwh/LWAwJhqnKntyBIfz0fME9Gt7VGeAcgEY7xX05SCxtHlPgVqZ
fZ0vfXhhHE+AlTsMhP/9EqLBw3VBZWNF6TZRnzfqYBs3GBL2aItKbSox3Lr1ws6M
O0TnqvV8PqQKlSu+/5Ooo+Sam9k1fLqhNGvV6Ud7Qu5u2GTB1KHKcR9MVYHgqvjg
d0rC+9fHAjn5/WYB96QvzA37j3JfAUkmz2RJx3gvVQXvYoOXROK9NoDdmZ5SZShe
KVPQLVeb4Xk7EBBWiMtpUQA8dArA9/6ylKwoHzjwH9P5RjgMd58sA5kwvlySWp4U
dOg9tUg3tR/gQkjaLgg9keO8xBqM6IbH/oHWLQ+UIeZGsyrclPvFhuiWn3IYP1bH
MT4ZG+t3NS/HaUra2Ox7cWZbcTEMSFmOHvQXs3LE3TOCOuLOsdVeVzSObb9vmhzs
7WKTYnw1VNW1wZONw43ukWXX/QS9ga3/2LS8hg/AOtjeF49T93Mv8VEDwh/gUjHf
sxvOf/ZdUmFNa7/ArFssuV6okMAaFzIv+4+f5B19Hn+Zl93+t2/m1x4E6/mK9AN+
7RmAVvWf6/fnEiE5NDBhsVij/2e+aUjb3qosgbE6LQeTtLa/I2W0KsmqVdrDWMi/
mzCEim7lYsgAi+UPsD9XwQUpTOKEkHLhfBKVM08Ct1QbnJ9MzjYhQwuxiQ6DCGOq
tqygISB+PmxbIcqhLX/Fv3w/fHzvl6LJtroAfB6bUMQ7c5Plf2TRJA6OG4PNd28D
X1YuPJmjwf+WhpfyhpqM+Hk1TOCYOFQTeUzXabSBPO7YD9aHIj5Njp4K6BrV4omQ
lAwAD4mDqsYyLheNS7TG9srSxC30koNIWa8hC0iDNFilOJvdqyQa4cB9jmUfm+Ng
msyZyeC2/IYkqcNaUMwNdAdcAOeCiSYVKC96+AN6L2YIUaMCeQRyyUbKXtYvqpbV
VoChPg0QCMMZtbRfviwHdoNCvEzfTnTGeEvJ3Ozq4UKxgHWmtrz9ukA+NkxKBKKJ
5MlQviQGsq6ApuYec3JKOiBMSUPOHMtn+Aju+gCMiXe6ERuVH8Ns9LZzj+qF3SOp
lQjJxn5voS/EeZPe2x5ZeyDe0lfYpKlIbRY4lxsj23/NECoKhmBNoL0bln6uWI3c
LFS+6yW9dnFAn1Hd2zsANDvVnNC3TVePFaa+QydMZNekpoZIqYchk7hUPhfJcL1e
zWuMxFm4lqGJjkRtbY3JWPT6FYOm1JBjcAXMh0AuViNTAu199bRn9RhZyXpaf3gU
eTVKabXRCMa6RmRWfnbgaaSctRQwfcHcJzg5X34b2UfqcbLRLTtZbJ5X9lU7bIYB
AoeA3Rz1Snn8LihPs1UhohStQDha/sOsVhRI/ck67kTb4Wg3feF8PL2IzFIlRCer
77CvAL8gCwlRiE8Kk8svIbM7F32BX7FThyR1Smf++hL7WrFsWr9oauFqR60aATsT
RFsPdfDl8hx9xyBjBY4XHwnPV8OEUnBESc0rMBa11qgdSmKYFS98/F4HmdFC2n0i
CZfAMe+3RDm+9fUtICeJvxNtVSTyEWLkxZk/4aC0FSn9v0fuym+Jury05SeDDasG
+zf1m6aoiZbeVjCGyS7rNCNaGbx2BOX/JV2EGxESnBtUdGT5bKjrO37aAORH9WQt
/eTIQK2IRKDtd45LcwimfmULNqn/SxaD2pc5Of2qMb2yUIyk8ny46RdStULZOSsM
GOw+osty7OpTRqeRu3qEKYjYoxYiVtTZRNg8lQgM1E/clEjD8LQPmIjP1MaZwPYL
wyC6UG2E2wzzDoGuiTFFzyYklipmvkSlYuWlQmKXrK0Pw3XLLyDzgotJm1SE2Dyj
nVhVCz4avzGL/Y+WEk7xbOQDIMK3cERxcQvS/WN8Scqd0IYNYFjAg9CjFMDYgVSM
LzOCXm4BfjRJTpy7dLM1KR1QtpxVSyg+YJgZlY6+quqDHhoHHoUJxAXANYVwLnUG
2qghqxr+GgV0mXhhs6QB6Y5ZGKk/U74c1TLQowf/wgTD/CDf6ZNlESPSCeBj/Fmq
0m0bGnMgx26QCjL3Zzchig+V0rFe+V8O/aEsLLQFUP4HfGX6uY0UadFdxPvEFYZM
dAdJuzZUssjmFsgQS2h8IdFtqrU5q+EAJy/r7KI08GZPqa3yj/pfZSYqDaVH/1RP
weDvMuyR15ZlnoZjTDzZ3rC11WNfWbBzHRjVyq2SQqxDd8TKS0gSk8eUM5ZGSmcy
LFm/VsJ+jDU2eiUPcx0wgVUPTEvWs9te2DjNT/9EfJ5Ziry2JavFZdI1OYY0Y/sD
5ODtIbsfEa69Bg3goZSesIJCJIg8dU0rCYOQU2i6+RW2Zp8sKRc2O45JNdK1sqqV
HCYjQZEcaUhZvwqo4ghOF1KNFBe/dq5RoOWcZZZAXJfRGQZapO9RCJs/pWgDRyL6
ePtwaggK+CUA833gfKkbqVA99jo0GZRageqgfwO+vkt6ILq465f+p0hwDVZ+BQlV
IvLeQVghOtXahPiepRaw+hbWSVafqNMhgwV6U+pxLlu9grERtYKB6bvRbk4vHBHV
O/Y6FmWYaSSf+iKK1mT2aQk6u5grHnnJSl5iHvfrUgTtpUSSVk6NaviwqscCa8BB
sC/z29liE+6LBxQYjpquvasd/Ce7sukHCJWd5kFgkiDxNZDmr18K7oQYuKFM+43M
bNsWt3VMdDUOH5+qWZAJowhpuWIMJKO4cUz7kTzLrs0/lBIiiy26QtTxZTFjvs6L
kjBDMNpPiHOmyGXKHL5H8yB0/izBJMwui/t5zUCUS7V34QCKhOTwBlRKKcPFNv3/
JZQmzYXR4bddcJieaIBQr55O+u4TJH0DbIBhNsSXFGy6dlRpBhNifAcZHwzg3uFl
a93G4MNo5neQSlzeVCZenh1VhT3UBokRrldDJKtJfN5YVXkmKTaiPyORvv3nofdv
IaaSzXGqdz/txXNhJirA776wz/jbvrfHjFx2kFxxZoRFCaGkpa5tx2hQMP+rWB9U
ONJdfhsw96LdoMUfB8Bbi2JbLmDmstVFMMxs06C6wIlccoYMBS7K55/sN4i6X5VM
D0dzNdTnIcG3OhVpEFG5MV5eNiv9M6qr4K8c2j2MMS9U2AwbosLagW3p/u9pO9/k
nNry2PcqOHkJPKhDPRydBsnGbjYe6B3SgYZUr2b8fTE/Bc7q9FNCREHfXoq6PfvR
/FnwBbS9PajxL2KAyHZgAOIBGE+3C6yPS6Y1GCrH7Und5LHR6flm3OJi8/QZhUBt
3j8v3T0YdhEJL8Klmw81/tiiSQ0tgiVKY+p3m1CKlfn1teygSD/hBuzctW0w2mce
m9mKIeN+LTpGwY8LBRST+wDith6Ar2/k0WVv5by4Wiri7Ru8h8lBG84t+IqTJ7o2
+MVyJzaEsXfaJpX/v5JRS56uCZ5mImt1/BKb2nqFgcTCxb+Fd/urAt5r7zBLgc47
00hLo4UWlrRm/yJMEw6qTL8Hx3pXVJkXkmF2HP26uzN4n6ZGVnr3BMlOyoizDuuS
IP2wwz1P7Enoes9tZbktI3JoVDF4zfrjRmJdhzC1RM8LBFcgHhESkDNm2aOWTTzV
sXen3A9OxtRpZHPff11PDKmFpVjfUG1rR10dnr5C7PPVtmsDpvmCvZf9uBV367LQ
yUyFHPUzsqRoEdxOOAZJeQ/2WVG8a4E0XnfUwNlGz1KPw2Sz2m6Bb2tKrsh36frB
wCPgW5fXQvgw5vHfrbyCNASw/c493/AKf0EuYu5YRA6cmTbIi5slaOyEBvQ8ECLX
/Olde66rWm5wJr72ZGQfKsjL84eXV5wmDUVNnES7uUNbRr1ufzmo2/jaf/UDi4qI
Ltq+aLj7HeDOqUnbGj6UX6ZatMbZ6ZcW/yBJK9T84U60rStRnprEcnPYnfdc47lk
YrUm5mV/WIqUGEhpp/EMVbmSWpzoQbzQLR7C6npRtos4j+6Jnc0AHC2dSFFiOa7n
oSUUl2/X0h5HMYA/f4s4HTsS1uE4zP3baim66kxkj3YWrmbQ8K0ChOiUBk7ghqiW
fiuoO+ltSa822J2DeVj7L/y9VeuCfPAQje+1yp/4+FmfYLAbqupoWCG7Y7hJL6MK
LyZmW2iSSe5XrKatPYoEzphgTPLTCywAf6GFLvfVxrgqcBHtHl1ztTEU0rmJzj0B
vwedPkDWWg6Aayl92frO3lcRJTolVRQvT28gre4+4jHctxmLA3fYfYc728kL/aPQ
jxHv5v5OCxkfR51DyucGNTOt0rrns0vSr4QbnXHKeLuedyRbEp7j+6yru8/zDjMa
wtQB76JzX7hzTQ4UnEosdHzFBGq8SHjCwqJFcRbRwnZU0fF7tN/gjV1aJlcraqIX
3xtH/8TAi0Pofoy6lPLQSeLxl0Qh3YIXv0f9F/K6IqSRCG6sEK9F/tvSGiBcB5wN
gsh+WUa8XZxVanP94pT1hjEqu3ahjyih8SsmBNv7OpljXQR147YQKpIujEwn28x5
LN/PN3WLv10GTAzZ/kzsuAQw2LYoZYbgZmVNKnlSWdRBcEHa7yNnT7yMdqUmhmyM
K7DedZW3dZS2Y2WMR954VK3BM6XPgF1pEgTJ8dhrN0BZSID6YIlhXTVt30m2ZCMV
EJDl117/dcqiyLXjH9K5JJg5QfwB2iAM2oZMCNQRbp7TvRZ1rKGZelhzff0QhBzO
kOg4kOEnkwYO3cdMYonpQoIN6YudbM6gVUgkmNXZHRXT28KKyfSmYqFRvZaxFQsb
GZuHowkvavuDQ2Z5oY/dwPprhhR/8QVBnQDdPzIIXAJtlKYklpNED3e01tzAV9S/
qyAWZ6mXOq/qSSjsqUG4XXOCCAZP5TjosVCMe6nmCTBfZEFt7C0vi7kMH0479lae
02QkS3p7MiQZ0/U8jgdjPlG/nkg5TKprdm3Kh+mUJXyCZcPc6Z7ar5ROXYsEBdEH
vvtT1UA0M2l6Kr9kzxgc9IM9TLtZaqoqbjT3t4P+j7rZNjaaNLxZRwucgl9+Enfd
Q1dj8kpapEoBI9pfCVgfP2zHm4k9msI6m5aDpbuBgMCE8Gm9Fom8kk5RkOKBZthb
ucJ5z7JtU7GkThM0qXsN8dMJMrWvQN+w8a1gXA5tNTBWn6BUY7WLiZ1YflVXGb8X
CLwQXGjmRiGuKsODph4XfnenwDhPqN8ZYbWSgcbJlOxYSVmDtX8jHl3HuSpyHXF+
0ZtzLzNe9axvv+WOf+c6oTrbn6W/PoZxAOm8nbUW3+e/DEnIjdykghG+A/GOjNiq
FD8pKo1/sxuQm8YgTwXBPq2yFbwjbLYToYFpmahHxM4eY9zQBCozbgZxE1UGwaHl
Ugn3xc9CvRmys2hlBP4+VuAWSNicx5L05IKJj2Dy2TDdTX/83UURZtBCrw/pkYh8
5jTrSUFwJFCcO0Excx3lJOqywk3aa+vff0YlBNNSeisYAQ7qgm7VA2SoFw1h/gL5
HVtR2Hh3k1G/CJc8NzTsmPtFJ/RkJWPNchsGJq8GCPWv8T14K1Cgo7+tAXQ/i5zR
jNzYNLQ7ZulDzwXYeNTS8MTiPctWZsRI2J/QOF28grmBH+G8F2xYZdnvPk5zBZPV
TwpQhvSanvVLxDKGYITKzm4tD8A0fkBPTsDiBvML67GAudFfUDnwL0oOH9VLxzWY
SaFHjiN+iEr6gHgPlnvbVmioEQAndn9TOrSvXhObZZzlEd9D7NWxKCxbgLT+jyPM
4nWMxmYkgMw4LQqTZTKhOrHMf5ZUnDDioXZ/+JL5UX1EDz4dlmDUp4tPSwvHZMTG
wfibvOHbu+JIXdOAUaLds18vT6kBhJRx7+WzvC3n0aak+dOe6X17Zmxx1Dz9hz6d
W0NqsTsWjEALkZgWVF0674XktMGLHk1i1m3yTOVmICxkWu5dD+/ld7GR0IZj0QDc
ww29EaPBafpyQ0gk/7u8upJOmj27FuyRK8Xn+XUbmujQHiv32jr/D3qKIEjc+cvh
M1SLmdE7kJcfb3Gsk66L7NXFL7hKABAbjYDBqp3JQcsmv6clyVdrcc35gHATI2BW
abzxCkLCqQvyT2WXI5jDn07xl8EEkK51Huv0DaoTSfwZplOCAz4CzWVxNC++C6S8
jXTgPJ8pzUSMbVTUlSPV8RXXuKnvVs0q81gTpTKv7xsjgCTmNh06bYVb2WYXiJk/
8l2zIASdeUPkx5Vm9Wjg3jtyxTlbOylLA5KbiJnzm1mnX7w5Jz/BgRP/cDm5YrYZ
e6BXJFNMWjLaT6UBpFLn0/jgpoZsrcyQ1h3FtwF5snWgRM1xNyJkvcyhFCRqCQyx
aD4fAh8l3lRvSxic1D5dKRA34T5gl8B2Hq2whpJ2Z7KE/rxeB+EMBMsEz3+uwzg1
Esg0/X6Eb7uQPPvBDAbAUBMO/B2HNvU5vRdogeDNJx1EUYgtYKEhiFE3vRUjhLZ5
au6LNC0Uj4KYx22uakbI8WZf3vsO3XPQWVR2ZSEAj/+svsbdCrKXNzqDfRFgAGXw
iWjyxkLxZBtFuFgXYekUhBnwpzk6D7+378sUhBoDbD80j9orH62IYnzrLEdH1/SH
Q88GlCQl4clW/V6EGNkAaJ1r4lnbKUbhgVZJd+npugxpJthcv7WXocJ7ym3CKz9I
P4IMnSnb7iAYyO4fWmYkX3sljV0Mk4J+7Re03qrSDn/wNj9xpA483dO1+6OtEvXJ
0jKYHSntM6xIxdHBJ0XKREGobDIyXx3UWjlC/K3N/fgXPgcBFUUEVF6ZExm3fAsE
PVib+pf2yHTQsB636RFx0cRHRAU2P8VTxu+VAJ/KLjEbMAgVGEb/CH7kXGiTQDnJ
nzM+nvD6rnf3E1hcvnaXcW4Gfoi1Jo9oX8ri+vZ7BAFK3yi+sMZpNe9Bq19sjpWp
tshUo9RlW5sfl7jqLgo6HlQH7lj2zmQVkza+/N7obqX0tyVM7zFXYJwCKPIWmRvk
HO9t5Pd72Pdbjj/ZDY5HvApNmo0cmN8HmR+MgUvC2tLsgfyIhSOuhSxEtv7VQDmP
shYDXbaFHqNHLRnL/gTbOkeuwloq+U0b+ybSiUSQqsG8QbBFTlLRDlA3YPCdzSPf
4WC1ppRtllsrbVxrBQ9sA48Ur47gj017mO0FirgBASb2w+N0X/SGOcw1rbnK7f+C
VPG53wXM3ZXIF15NH//qe5ZOVF0/fhvtlmlzoKO05thhVHn9O9jJc1a4iUvCEUO5
nuPLwPEUHtCnM+kK5ZQ15dBt3Y55YzK9qssSIWOqcjfsTtyyf9MltpAJYyTc2cq8
Z/V8M4GTjTHjiJZFd63BAu00LEPjM3CPjaY3fgQwHKrKuppud5ZrVN3VWSjIvVUU
PdG5uEAD23kQ0Q9ge2Fh4SvfLfqQlq2f5n0dgiw3ngpyi3mqLiKanzMInSoT+DHe
vjk9YlFvd8gN4EZ1VLx+mdgQMHFSClesYs0kth/qwSAzTkPm1fHW6Ep5vPy7SHoW
AakgLgaBF6FzZ414EnC0Net/yjRkfavemSLamZ2XZ6uKuV2UtxbYaIxIzstjRMgA
s6k/0WUWKsmURUhzzvQCJl1s/TmgtIdzbQvOU8UPLJywZ01B4+OH/5DrkSiLZN5T
LZHwYqg0sEFDiNAyjXnOfhRHckMr3K32Leued4Ev5YE3cYkVP9aPrueLMFjdG6D0
KEvV0Gzt/CFCqE2FCUvxsxqXCDGHhLasxIHjB/auZywJ/WwtBmSsPTthbXGsPji3
5TYFeWiHgeWssxnMLFgxZ/Bwz3EZQFHysfn4hoNv3fnGIt6iPl2tgAV7IzYL6Tix
HhMn85YKoIQHizp5l37/3SfWsfmu5H0yAo8QyyfUHqt/AtYWbDl50NS/G3rH9xjB
IUgJcHGki7WCdp1vdz2Qy4Dieq9ig5w/kCdANnHC9i7ncbnN9HAXFeXd9ZlDWpli
5Z8v3RtW5DfnG/2Ol3Xz0AQobtZFpHVAAgDyAmWaijAAAooy3D4DqoNaEuqIG6N6
p0BJ+IKCx6Kjgsf/EJuxZHkQSymSlePDQPdbxZtM40d9vhkHLFqzJGv1GPA65ALc
r+IwWixqKXACsh0mkOZgFdZObG+2sNTydCwCcW0TgRoTvAOm248Y/SOzv2dl6gWm
WRo72XLkjptWGQyP/NYFx2qag+g2akc44IEDsdEfcgB3vbcixhIWsoPyt6b9v1U4
FeYCrqwg7/R5Atcrn1X8s/AVpqMojbnSA9h2ZXc5gtJ1z9+UVy8hUoMdjRpx9Rda
05DmxxmkrgHxVcOoFZJbh5S9xLOLwGeAkPLKu4R8iZmjsHQiOw+Lns8OgIXDS+R7
uCdt6riTma6pb7qRJ2xWHzhh/FsCH4NYIqMdMWUQcuivtYmdsw2eQ3PXFQVbGVAn
0wGsGcek79AaW0gA7pA+kPKWYuHLzXg9MS/U+nYcOS1xRDfhAUpybhdqRee2C1X7
uyKWi2HeW1pMrV5eCpGy6absHuzkh1VXtguiVyCIJO02Tl0gwXFGymqsj667HXJM
aFVA8Xdy2bTwZWjH99IC6yCf5R6P128slWCqiNFeOZgWah7yAXVuptcMjx3WVGGu
3JfTZN1V81/HtqUgvPaFvEb605l0/ptnxo5ADKGsCMAxQ3qQfMInJEAWwgDRDOvR
8sQMaZGlUaA3/u2AnIU3EItPAaKBH5ioDhL8mNX/PZkeJkLJCCkV8WZfuw1CDMgr
Kswjnom9PAvz48uxnZjGl3T8AV1v1lJ1xK5IUbkhaiFmqw7LDlpo8JFPknew06XX
U8P8+gqHN/R9cO90MHYnP2Ix9sQkYh5QJqz2wl7JJMidQA9zYIFEcKs1nMZGlFx1
U4NvtLkgRy2C9ob4LJML8cXkrVaf9dNmPOtksOzbBZyHtcO7AuT1gm/die3Ryj/x
7Xak2soafJKzg28PrNw/N1wTDoeK9sGAsnZHklwAdbxC+AE2qRJPX+7LSaPW6ReL
YJCWDfmMiDtW6OE6pZPdsy0XkGEBZd4ZMWyEQiUmFKIESO2pFIrIA1o3SmTTUjJk
1VI4oIIcR/M9YXwWNWPYohCrKBEJkXyX+DzDsOnFbxzZe87E/XxPby7xbD/Btmsc
TFGIeiMSJgLgi6nNPDF5gcMvp6HZauG4lkSihhFNE3+Vgfw1ofilQCjp4cRimEwO
Vi4EXdeoxPFFo1mQFVRJm84hp+E6djO5RBbk2bzpX0x3KW4aghyRmytnFaxqJtfc
VXfzg7EXZeS7EgQolKlLgu6rZOlbb3iEkbow8IqZKfTQPWi8iMRpsqkfs+UeW2ri
9R4qU/2XaK7gUvATVOGSuNf0BhIWddAcT9YuhFokP2OlU6kVQE0O9ziWhBNxjy+k
OL8Z6F4fXgCNDKeiczWpOEdd1g0GRMqQMeqUgYrs6xzJx4vXAz3N3P0j+adxGz0R
IZRsixt6Hj5FGqjl9NohbVquPkTsFXzmXTyjoSgU2sZbFg3ld4paa0gZ8ZPDLWQf
rbfcIa2jdVrD5fMOc/1O20RWQHwpJtoC0gugtATQKjcUJIhAVPGctktUE0CPMKjg
hIVpH2590Kt+MKbYpjoYa+i1tV9XHa5PHbpTebUVypq8N8Qt/GVKEBeuBW7K/LJd
ofo1ixnqzVRr9dpRA7FUk/3QnIlG1ZBm/0FQ2ub/sfLYltWW74Lw/FCx1oYwyv3N
Ej9zk5dc8hiAq7MJs6J6eo7sISuSY5644vinxI+AHI8pwBfVREZPGr8+0Ue8Tfz/
jKzHCcJHw11Dyg/db2CtjSCGN/aKLNSSMfoQDRREadSlxm3DywY9moq6/8WF+mBM
aF2u5v2b3aXkBeEKQcEaAkRDZRcMCyRU4+ZtABCj6FtlrdTvpasjcC8SV2jumYu2
PNOIdzqLlaO+ofx8eqzgLYBX4wItpBO784VEgHmHnkXSnkCx3B8DIWwOJtuw5j7J
Z+zseTt8PWTxImND/5tLJDFbvlw0KfrMmtHSuitmJdcPJ47EMF1Ip7PEtEgC5JAt
S1hLPfT5oO+gMieGF13A0AjIKg8rpybEEn5Zg2hZYYWpf9BsPzyOusC39yPM0xnZ
FFFddEO9HiVjmt1w645tn7p3ETxop35AMB7jlbhIuOx9fsfFic40ZxI8HYSM3FXO
4hZ8JsxSQJDSUGz8Ing/Cx5T5M4/9JEHMsCREZTw1W5PSr+HAksRLzhbZT290vWS
ybVqp97vN8XuNffq0HgWOg==
`protect END_PROTECTED
