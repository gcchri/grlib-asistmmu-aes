`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WGsuD4luV0nm6CEWQOH6hsRpfjVjwCgdmeibhjJyXFN2W53NgQQRGcw529CWA4JW
bEBqBpdnkkH1jhLgbsF8fh45Ux5jje6Hsf9vjbDMQpVekl3FnlAG+CIdtL6+oSgZ
c64Xf13lrzw8frmH2PLwY+SZdDPfSoSYiYMcDLbcjCS95EPHGrTxvx4B+Jy7AGS6
co1flfU0k0tYP0iO+v+ELIw4EvLq3jwquJB0Yw4PmlPzsZy8o4Qwxn5InGjmvr52
htyirfqqrd93i1Hh73HkeMBpgN8lyhWlISkSLnIevpQNhkbnITHJ9SljkWd3Idhj
HU2wjDTq1uBCnE7ka2TzKs+xd0RU+B/pKoEQfuywQ6JdHAykbfh/2vJDXrzaGYM5
6jygV4XLPcriqq9UtV/MklNHavtB8i5jknZV2P90j7BeKwoCM78qDGYWwrWRTHCE
`protect END_PROTECTED
