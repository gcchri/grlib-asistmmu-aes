`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UQYQZS9H7ZieRV+4yjwEMHuKwptD82QwWyPYVylWTdeeLCkQXiWs8RYsvEa6BFEY
K0A9jlyNeG9Y2a1X10DAKT0hdmMIvR/dEGI3sQVdhwY5CWHJlPhq93KxjiGRv/e3
nvXf2NlWzQQZDmcOINcrViASHG54MmBKzN+KvodXgp4cGcQ0Ysq5OsEZrRAoSdH/
GIA6Qx99Rft+kuVdeRgDXi+6YhFaF4dB2NzM7IOuc0F+8V+1LXl8+x3BDIchdolo
J8a78VpPrgQhn7H+MxcB9Q==
`protect END_PROTECTED
