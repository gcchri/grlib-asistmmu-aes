`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rPDsvUWksWNtSyXfl/3EJDVDHOVQVAhoV9cAcHEfscbRC5NYNPUgDh4OHMowdCzU
h5Pw5cYODq53VK5MNFG0zUltnQ0gJV6LQN4UfIQhTMXHBbep/yBL5l8qx7BMJpsb
VoW5ZFjQvjfEdCaHXjnHgU2y71LOeQg3EleQXoinXPfzdcnAKe+01JnSuObV8Eln
3sAfExHOfPWLtOoaxBzt27z5XexyT5aPWT1qfwBErmhxGPIx0CQvox767vzJp1sS
XsuCisfZ+j/NKVtwApAqbK2iIWCAIDxFt23wHMhEmReS3jYdz096yLBteDGx63F0
`protect END_PROTECTED
