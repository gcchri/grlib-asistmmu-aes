`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KsiemHBeBOrpi/sUXglfRWMz0SrbqYlQsPVNF195L8LJvb5AHdZN6GKS6XUZYoPM
0OQzMNVmL88KeEi6A1b8A7frGv1I/gW43P0cc6g06cLyQHuYL8OVcHNiL/DCo/Lf
eqBlrbYVbui62kY9Ixe+ZZtp6SL7EOWS4x2l2W6L+dYTju4Vz887QmGuyvGCtstj
t6fAW3hPoG9faQOSDkTRVfu1oLVjK8c3n85wkM9VisFsLAuOCvyrbJZqE1S3I0Ed
mTFgUzViX0P9N3Sea8FeXw==
`protect END_PROTECTED
