`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rYYpWqQDGzbsgnFho+tYpPLMtQq/IWhJsEaBRTCrikc0WuiHUMLxxHPLg/DTem3G
0Wrv0D4s5VoCUFZYiVn3mvObo9cz/YGuGOEwao+u/s1Bemm3edbaJq85eTRqkBs5
5m/Wgq1iqxAaxr+4W5l68PLpFHoy7a8LRxwW2S0aaE4hycO/jf1x4/arxc5K39w2
Dk2/wQr8doF0jwQXC0rtggNXx4P6olmUbY43FaPiZprd52QyWzNlsDm1N7bU1rw2
gNpTiyAe+WjjPe2aTRNS6JFcC+zTqk982/ILmGw5NpQMpK81DF9PZoIKrWrXl045
9gpOHYia8Bo4AdL8lRLGvhK0LhmwTfeXrkYlA9gY+4JrsT7qkM/3u8O3kf1Y9swS
1Dp4e50/yVNBXSGaRj7foJpzMkhvHD7tf5q+lgWgDZE/d2S09Mh6BUzxuC1JA14u
KmIFcL5O3kHVZsgCbNvTvwa1ffHonQOPuy0iPxD/s9Q=
`protect END_PROTECTED
