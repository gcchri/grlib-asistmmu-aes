`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tdLA+rNa7bafBQJqTnaMyH8FMv5MLqAtKg1Z+BpmtuBvXVbQjXpsQPhio/3AQXi+
wcML0AsiC7Ps5yIwQftktkXJbCoCR083csgelrxf4yVSVhotzqf3jTup228CfPfj
vpUNIgQVAguoo4pFLOFFwSxD886k/8XhWzKEBAREpuFI6kUi7YoHuvpR6p5mcIoR
4hmHJ0cRcIxtAXnT3VALWq4CVXDOM0VfH/RdK86hzOI/mtizsq8LUOj3Q8UxCewz
VyRYqqnI24C4GoG6nxQAHg==
`protect END_PROTECTED
