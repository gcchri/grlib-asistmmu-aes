`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u+7ExHRT4dR0TANf3JZryIp5mEUgiMKxiQ9GpDPi5KVO8zwRNXKgbZCmmdeIDTdR
mT3O2H0M+NwafW7NkHlKHqT6BMbv/u3L6dIOa1TEsT7stic9JJxXDvpIytBXW6+1
zYG7xuVXqTg3c8/ayn6K6bUpPmpMxUnxkfi0ptdXppxEquBVgc72mDgSuKw+4x2J
hTKq8Gg9O2lnwy0b+LefvnqfXYaaPq1+WVPALZHQWOfC2/Tc8CJBpqR42TqmKMF+
yOCeFMgbHGOzXlcwKE6iIyKqJ1FypJ5zWFkpPYgH8IT61+Xm/Qy3oHnJJ6DhtWXl
0Lwv+hZKuolngKkCMGKS0kZcjj34Kt2q5aCJ+Ie/1MgBwCqMv7hJEHB6N4U94uBY
8yGG25uag8zRVhl2OQwIUyrcYdjTrvT0PKS/Jlb/+ZlDI5+RMd4zihrhZ6QNTd0b
`protect END_PROTECTED
