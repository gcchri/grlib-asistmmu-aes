`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7+uAUVCUoviCuKYAZjpglsA8E7ih3Wi5oxGTVyu5YZD9qFBAPxhOKz8Eka6LGVm8
9hU9Nixi9Yzymz/Paxaa7bLDri4Z8ZdDHkcbfRzt/6gLJZ21YhWAhmDwbpk8Svc1
avMrp/FukMNrQEZJZ4hXRKTWDD6lOY80jSLpvFRArM5ToscFIRDJGQGJaTV35DuV
hB4p1GpbaPpW41Xn22Y8Q5EQGVURU763ScV7HqFyAF3GbMjiEZpBbxWGWZ8cEmn+
SA4KQpRr3J6WgDrMPR/Xh3y+4psl6zbgJqubqslmY1M=
`protect END_PROTECTED
