`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ves7ErgPEn2XZ3zKgUcZB4oP8Ly7a6+NG8nkfvPzscd5J0kgDbrZjfTzbLZH65IP
rXt+/I5caPiOMlpgGTPy4SRLdZHuGAVeN6eD2/hxlRY9ujs539jCwMc0wTyablhV
FCxfpr6ezHKgO5yNeACs2j9HjDdYnSNE5LfJi4IAfd6F8cXKYr5+S+qXOo8/9p7o
DCXcxyXjITHGFzhmm6ezxWD6aNib1AQNesrfPk3wPFW65ogsiEzdQ1kECb6vnQBX
3/YdN4wv79JWd6CXijfYl50hWilZZyviaduSX+QMErVTOGACK0+pHd+Ea8AFgkJR
e6YebOCSoPZHBR3fkEiZgEpwAVXuX1EvoMqs2XrqJ/HmYOtneqCadCsLSlJVYSiC
GHlVkAu5xAnyJG606jL8THsgEayDXaRoyEfpjNfg3MjXFezCAgu3i+ZAWWVzsiDd
`protect END_PROTECTED
