`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2C/2wa3A43WzCcCG96f/V2fqppY/GBiPqHeoTvzTsBrh2ofx9jeK3yw+ShAIljQ3
F0IZ/vZBzmr6mFpARc/KpCr79u02K2l+gFWJhO8Xlpyczgmr1mZ2+AQYb+pDlqoy
589Hw5K9EgxxA4QomAvDohEai97iEh0sf3/WZ9kXtGJBjUpxfAczOtK61sMB8ZeO
765TFZOAMP+3eAw2w0/DVki+9fGj6yFifdacQ6Nic2jBlL9TT7zCWFpJ+Y4NQ+ep
UgDJt2sajQkWUk5loWhZmKet2Hg0w11vvexoaReumyuC6ipcMAU45qXpvlvomlZg
4stfegmUUkxHALhNjYsvjFHmL8xaY3Wfx5gClLF+QAVqM2lgLKtDGnXrrPdAt/i4
ToT0bZzfDM0uZF8KLOC+1CMrezVd09YO64XqXQOHVXK653y5M7wWXEllqN13ELSz
YJI2l1uOBFdoGgGJ19MC8ra9N5S5i8pKFqeKW4kVGZk=
`protect END_PROTECTED
