`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DP2/Hh9CeLq+NP/O//cF08Mtg+EyI4YFlQtjHUSnPErW39i4ff+jP/aRMiclpSw3
uQjjr2xVvkvuo7PaBEsszFvU3nQu030L0c27NMqdIwkuBe6IAjr/dJkcc2Kk4t4K
sSCmv1GtZgBoSv88Gp1sP53Gw99e/vt4CyMWLcPJcUM4ZEJtvAqo+xIFTXicyf2e
uSpMT6Ev2yajvDDYGLxgFAXdV0rvrf2ja8WnvQvU1lM9/IA4lojPYHDKG/hblfDK
gheDGAW4duLFYGrwLC5TWLu1155q3Afr/kTZFD/khxy94jRrgZp0lkzFboewGN+7
`protect END_PROTECTED
