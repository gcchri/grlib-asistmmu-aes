`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/7m0niaF3jXjvc+E+kdpwkk2IEM2VD0rOfh/TNIuqwiTGb+vNZRWpg417YMwlLJE
g6XkKuP9VygzrGjNnXyDhm154Mf3Dmk1K74NlUSdv5UAhQjALE0F3ZmYS1Kl+DPl
dzCXxmhAZ/eAWFW/9zIr64hwKiMPuYOi9BfSHWZqDH1LCHKvR3ktACSfairMg4KD
AfM9DA1uCFHllTQRjKVmbj7mBZGlkbRUiFL0mugcspu5LouQ3G1qYlzt/VJSDr9U
a4XIP8rqRYw4jTBZTzXS76EtXchE6iryuAEy7woOh1ffNPw+oBuDdhmNVD0BGNGn
8xkHHq2GB1ufkEdCQ1e4MvH90RfPTME3flGg6k9O74RCtSrv5bT5T8+MqIWULDCv
`protect END_PROTECTED
