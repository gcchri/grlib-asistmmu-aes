`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ceYPLByDD/Y6fcfl3cOQPCsBqeoHJpxInUGhKJco6/DM+tbeYC2hFSCVjScwYS6d
dlgpSsmQdLHghfflWrdMYehcdeF8IDNb5htjd2hUJnoJ3r4D4cIiODS5gXgNonK+
X9BFnlIrwrmBwg3nrLlpE5Yzv2ptP+CEkwm9SUZrzsu1zbd2eEhLboAcplXhgplX
L2Mpu2GV1fwqFtyrP6zfbgQk4h1cXi6oup9YvHi9SWx4HVNmk2cO8rBR9J+W9R1Z
J9XoZwV4QNEIcvA+6SZNubMzD12Sdt3ccgWSivREYaSK6YtL7kHcMRWzT5TxhGH+
qnCgZMFeQoq6+drbcSDJ+y6xnAagBDhQvRXAlZZiXWD65QYuIYx1t1trx+tzw0yp
GmtErOfulOd+BFsUzXsPTzAuFv065untvX9xvprtqFWXoIg7RVWND6UqO10+dK8n
3+AloukQHtuNSNx9WP/6kreC0n+cv1PFAs5J5QYkBao5nD+KFEy3CQ21RIfSHpJS
JpbwOhP7HPWvFaXr5GmLwIlmwZNYB0KhDFBdj01yoCAqWIOOnXWrpgB7Tv75lniX
r9ZoQc90VWIh2R9obkuWKHc4tg9ZeGCkUnH3CWNWzuL8YZZ8g955JllwwWvUdVog
I3bMmQ6l+NKTyOq+Z3sTiuZt9w0sVpS4g0w6c4bR9AL9QYd/lrW3B9a3jFewRqjV
zxpWAtrsx/2O90d6GUD5FFXtFhEzAxg+eIhJZ9J6rjuThvqRG2XOWX4w7vu/RDK/
DmgXuGPMYjfZJChzXczgWKOSel3MO/6qrVbMkpKvD0+pe2Roa7HXTuBMOWIrqr1j
UeO3+3eT9+FxNe91exu0c1CHe6B/smO9jJVh3dtCu6E4D9bCLf3ISmrymbD2Fu2L
3XfzSVYZcQaWrHboiD7MiZnwkk/5bOYab71YY2rgb9Z2jBSKUU5jH++q0gTQeBBp
Y7LqJLxKHYWenXsMsTlpHJhxNG6Sgrg3DQt5FW7rmtTqrTbArzXK3d7WTLkCBXqd
ed/RwALptghmapnAqP5YUql0Eck3HVFhFnkz5gXFNVKhpcJnvpOHRjSD/AxlvvXN
jajUzFS1aOrEpb7uRowMh50SiGl1LDGDD8SOuAfyUxcl+LfMs0Cn8PQP2F1nWQVh
42EBlyPFyEZfrnuE1545NZ9M+vaquk9VQ5k8MGRXz5dm1fdOc8gszY2rUIGrYFQ/
VW8+qWjixr0B33DtdtrGGtltaOETBn5Rl9QchDx0RXeJPpLEr9ZqdKs/bqLdZUgY
qtJcJL1suR5HRDPDRrfVAN3vQTIuxFBV0e+uS0GW3MaWO2sjFrTfYVd4hm/nZS50
KsnJ7Ycj5mWVt3XKC1+HyL5AHts6zG4s4rUhI3pjH3bFuwKozb2vR6T0HWxXmadJ
Y4PoRTdaN7+0t2dcR4RyUtM2Kc7AUQeo5GrtzswI7WjgDtbE/qoRQH14T2GRv9mv
UDl5xnf9cIfsOCgYybbNyB9I8OAgdi08jLhjJ6Y5w8cu2drX9xQT4NKRWmMJBqbn
r1XznHkvuSo5m+zeP0g0PmyRrab1ZdqpvF9vbPP9LL4J7ztnrUC0LDT1VdCgvBsZ
fuJ+cRsezqwcgEK7/gjf99kRF9WciOIxIzdu4dS4kTK9RfUYeUPNUY9ELfVsustS
96Wa8t2D8Ix574YKRjdVjBdfy+1OOzu94teNvhLsmJtoHTob7o4cEXwKA8O0CCEu
5MfAQT5/t3Y59jKgF9TorZHE8rE9E171horKF5KWDM/1uMGbMt85EJl2XO0zZ1xg
3OGiMt+BmR+tRnonY/4kUb2GEgY/5EIio0rLlVp3UcY7XAIHaoKwbdyvXRnQ7qoc
ZkZCgz2orTKp6fFk5ZnfeahEJ7yIYxKpFlhl0PeptxyKoPg5i6JWU954hlC+Jf92
Jf64pBrnWhAHyTX04+oDP/oqvSJ82CaXsQ4+SrLa+zWwGPQfSnNA6cljGSBfHjEC
hIgVw00uNEaIv1BZg0tlIg==
`protect END_PROTECTED
