`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6n97XIWV/eNCYB/vIoelIrXhN6Kn0QiIpXZVht44fDayM/ImzTp4A8+UdwIVv+Db
JKTzGViY2+Xmyc+rbDKGNCEyONXv7cP70GS/gviRDDeg1Zy61sZqZL/iT1c9AX67
ajkZbhlrGuQYfCYeVsCk9g/ivGbs0O6IlVtkMJNchj4Tulq5vM7c7oH5++k6bvG8
VjQOnvLIDUFyX3VDlXeBO1zTS0EircPMchedc6N0uVfJ8wz3K3anexjq5VpjDpnw
nwIQT946mrf8yJs7nLcxHsfmq5eBKTwWF6jqiXKGqbdC0oQi52XGha6oEcAdXK4u
hzwE0gTLsggDoUEtGSA+U8eFRrKrLn5g1W+WgE/JumDoZPgJoi8O5eu1mIFiKIqF
WdrXFqwVbF6G3Sw3iFfhQL9E0bRw9M3tohJVYl06WYEeeN3Wkj24Ry03908DYO5n
`protect END_PROTECTED
