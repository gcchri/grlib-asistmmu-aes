`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k72jZQGSzXbmTM0MgB+8EqAjlwuZASiqnZyiQDKsCoCGXlZZWd/xgIjhvdjkCjPc
aaI9k/dYMlUWclfVud+Mz/K34S0mxHqGpECrRBGeHgIRBS72WSRjHTDvrLAob+lr
iEcsfzGXplJL7Br0NJ8pCd82qoqB3/gm4I5SAiwmWpKLLnM4EiG5cjmEYWekP9Ia
gr1u2NK6FpS2DzruytgyLFIR5pnXhrfKdXIKxSFix9QT9/yAU1mDOcjLmStllLDD
w657sO7wrd50BnnrJ5UEu3kOi6Uxa5+uyEqQ+fp87LqVyAYQVqQZxW/76Dc+l7CT
pWi6m+HYaxp5Kr3ytlvs0lvZ7xmOX33qzeALJVVDKmxoLdnpt1KN/qRi0RRKUs66
u9DqRzvA96ZAlXP9bwvGdO1YWP+eqhHz7SlY0efdEVhEa2KGPBi/BmauWMn1Ed3z
bDIXrRtXX2CeDYuTZmECnLSgUN6vKNdmProeHL/fD+T4H0rFcCNL5mpZ+zOsbPTu
7GrfH79naR0WuSxiZjw0fjIJOwdK5u086FSiza307mHW1gZ0WtKWomvLgdmLo4/V
aFvSigxSwdBTyqRXxG7QUNvJrJ2lEDlnHNriEdBRkwK84XCvfYWMK+s90IQrCJuY
Y7h6e/hPecBwB3wjLXCO6UGLWP+seHeYBngZujgtvnSXbzcK7afgjZLx7RL7RhK5
mKOM3vr1gwf9RrVTkBOa94pwhj5POPbPTZi9LzO3sLikEjPoqZCvMaKC0lG3DTcv
5NTrLnbSSPIbR2rar8OAXahoytfSQcQKSZ8EyVn+A34MQKZ8Xo2adtlY+/aEmt90
DptqWNw/vni+ohmvYt84PKl6CfP97RsMGxlZ4lG+HUCL4lcHCviRsBs+adVR61Oz
mbbK1gMKdX0eEjh8hkCnbZuaN0nbd4NtVlHpSvkpQZZw9ZQ0RJ/9+0hn030J2BzB
PFTUS3cg+GkArRfDyhONcZnFmVw6kocL4i4K+NehRwLNmZl04ivQZtCzQHcKz0Vz
Htf85+hvK+RvESXCROGWbyWl4hgX0bcIt0GV3xnXAC7RHpVU+cF9E+Bhai9VNwXE
zEb4pf2uIgA8iMaiuAb+/V39h4AE6AyL/pCSQu7ExJcvzugf53OmWwb1ChJiVx43
oP65NbbJNX2bVx1iDC0PEkx3C1jxxUAB9GdA48WRPkMX7PudYiI1LYDoIRuhCS5l
3hTQkN0jn2CfxMF9LB0OcSi8t34+CMF4VNWa9AxAo4+N8fZJ6wiYhJEm9SQqwX3n
CqTmom6Z6tw9D08vVMFrsLcGzkJxkpwOdGpMs5mhoMsa0/RiRE7o3u+Oo2F7U/et
`protect END_PROTECTED
