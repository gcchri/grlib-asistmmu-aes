`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pjDwHwRZWqfkb309ol7nl/ArLm37/t/v9J98/frRdsxAoM08aJ+OFIe7s6VGLTW5
TOWIIFn3FsCIb0IeGTuzIpfLK7ZxgpExikHDzq3/yiEDs2taESAdfy+GKgJsQaY/
Yg8z1OzUoTaHLubuLAIPgrfFmRPpElVF9NvC6EOZXDddSbIVX749OgxQsMWbdQaX
ZOW7wLD7AYjdAd4NeMqXnWuo/f3aypd7+13F7HewQ6Lurn5DzMp4VhxUD7NqSmoR
8tXJtiWqx9BeCitTtf39X4UtPiJFi6KTFbUn6Ixo0vGDFqCeIRvmwaqNm9S2ZvHL
ojECxHaoXG99jcJYI+Zutg==
`protect END_PROTECTED
