`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cc1n+Jo45q6gp9ErRbav+jXayblBL2xo2y0n7SE9+4SQ+8DZm0a/2ISaoweEchBe
rmfNqtVbGBXqbzFbad25tgkBRm2KRavwW4ZKrGwViKW2Wl2szlMJx3gYuQZMp+3B
sqIBkGq53dW1DKgknGixnpQe20weblENKyxi1ZeAB7pRS2lRjVgnsKvgEW4ZnIIg
35LKgcJvAYLiJUL2dubByiQ9PHx13P9BgxuX6TOZpflVwRWZvVzUpVb1HOsgR8PC
d3CWp+7oPzBvXdzIm/oMcZgPTdY+cr9Z3ho0tFkaTGd9K24uKifZZCd3XwwyoJkZ
0W1Bwc6AjHavLskjQ9Xif1SK0prHhq9fioTp/i4GzpZypzYwR6nFsfsXVtU95PVv
0cwYCETrKc/OU0Rgo0Sx+hkJDnB70QPQtcUrXcMhdvJWTLb/Yo5HLcy0l7BElNhz
M4pSTyLWbe4PFyJfIL1I5R7+jHoNp7whZuG3GoFSbyEDWLe+b1JcfLHfsdtrk7b6
ea6g+ew27nuqNbFHhg+yaQ==
`protect END_PROTECTED
