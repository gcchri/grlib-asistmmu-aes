`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f/UZ5hh8pMREStFQJCjN4YHIqhnIi2VV9FeztTXokSplEVXVYIvwhBqFo0nLF/4M
1pRMR5rtNVz7olGINaVGLs3IWk3RsYjFAN1mAh0Qyc42T2bsZ59me/0dbbFVUO60
DXwiiuX337JRMvWSrIQXP4Fv6+4nCW9LBEOTECP1oWBkDwbyztZfN4GvzTkGy5h1
7m3064WIFR7s+lk+CCkNKoO8rSCzxx00VJZ69ZhqFXfTyyEKaJ0glaCnJph2UI47
1mu+DlhVj4X1DzMKDr64+1Hv0ZLD7dZgyhcOmqOoxyEoJ3DKQv20Ve98365dKcKa
GQZvh19b4jjCM5d1hdpvqTai3cMlCsGOdjyMrKYfRXKIjOaUvOVvluHOHU75RytI
AHx0rpCotBdDma+oppOChNZgYQ0KUMrxswrvtnDQhEFlgJ7xEW5eNkdPC5gaTxVT
wED7NLRlu8vPOCTtSDeijCz8a498C7ObEgqc172V0J1Owz1/lyH8hP7nz7hj2iJR
4e3He24bQxXQgxrJrFju/VZYAt2XS3QI9bidwzi0nW8FmVeprafzLWzWU4oa0jl1
nlZJj549zm8qor/WIqR2WIxAEPeqD5Oue+Ws6Nfd5SEjqeKMW5PuimbvC02N4WES
KIbdK1u17sgS6R4Xu4LXvzGUli3J5aFK6igA72HiWyNpOpDaTp7/FzqV9tMzn908
GkB04YTdkEDhEfyv5p14Lvrwh2vpFGr3kphsbN88dW5iCyqxvqbNQXNh2JgGF7qO
Cpo3xPOkEWF20aj9IA8oVs+pgWfcqmc+bU3VcRB2l0be+AfVI/Kk+Eb7QP+QL+Ki
8FZq3w7VTzW9W8gCyxHAGQ84NbhDZ7fw5Gkqctnn1F18ynlywGVgYlyVdpBpdw8E
cEDopwooQ5WFyfoliyI2fKlGZFRXJJgbXidZODZGeG9YzKqAtN/TzB8TgW9oIs4x
XwMvDDP/Zx6t//PZsVSD+XcDgBbysxF41YBlc8pw0eMvVJ5evOYW/8sfEcugAsuz
qKl7bofKUSI5vo4Aj/QkhGfzm8zBeaNxUTRLmehG5HoOw18pqPZNYEFt/IWKY5+f
O8zHyYfSfZSmZj94/BW8ApDiHbtrmyXapNDSFYig1ILPNTJywFYjwjmMbu+LFKkx
R+Tntyi36kaUtPNg+QCrx8i9oXLszrdScLC0RfUBhLIvZ4mjP4oCbnEYRf1WA6Gg
Q5Wpm4ME1TQI005+q6+o1adO1ERLoZXSPJqk9lWuGgwk4mqhRQDALCQKx7lzpk0F
JZV6ob8Jd+7U4jwJ2nyTxKuvfEXaLslLE5ifzBGmheQOnDEebd80m2+bykCiX0BO
DrggDjgE67SI47n6nV9djfTaQMjmrjejIphB3HxDCRl2roExEwhglPvHuoOLpd3f
kQXrtBFdhfmnUY/dlhzFxtLqGogjgRYAPjO+gOGHmYT57lSNBC5nE6cwIBDwgImH
4fgsviukLvGrA93GAfskcBf56BYv29sC8zFNl2GYisNFtb9Z1UllKXVE+pJDXtP3
JPec1lhAu8kY+2WDh8yybvR2bXmxOyqCunaA6igQnMZBtZglTD9kkccIWzOq40Eh
jg9hiz1irNo4FagmH5n+b8RV583BHircXvWztzbN927ixVQdd3sqm7S3ZSsBhKZU
CuX9x1McnQPxLujdiGqCIXq5IqJvfho7+dYIq/vsh3VBoPsRRbdFOgnzhAYks1OP
XNp4PTJ/BOpdk73ua7IQhySeN9NLIzr+05IfdE3GukDxj0OY1psIY2cwyyuArmdC
iXQxTRVw5wdpHc9hxp4cLOjbVGa0NJMN9zLJc/VGBnzJN31aXTAVRkh1hipgWZI1
ts2J1q3d2CNBXSFRq+WRySlP5whzzyfVJi6pT3K3wRD/v1ZAoSm/lAmM67/RL1dr
Z/Kn/ZS2y7myj7gQTWxcZTVX0YZl5zT8Lv8NPMQLReY7WDQ3Kdilqh8lODHqK+2i
pQEx6Q0pmtbuIDXwjJslSQ7pB37fmljBiKbjXUsdvxagV7cxm61+MHY4MWy91zfC
T36aQpT0WEvHeIT7CHlLZBuc4AOdmQcfH7KPfwDoQkV97VyZpetsLdTdK6th47KK
Krh3y5veIxqF/fy4n+ZgXlS2YBmUMXuBz9S33zMQtbLllLomb7REzg6KVM2OFmbb
13OFOt3jtGyeZDK0k6OdBuwEtP6X+Fx5x3fK32zCPExpZ91das+rQAF5jZJKlOhk
AeXgKOqtqLkhQK+7W2R2/tJunaz2L9dFjggmtTfKoVq9yoXpsDhnhPTLb/NEnLAi
e9ATL/IVv/+aY3ZXYf6s//AHt/dGstgd2K9MVGGh2LBW4hgMp4N6iPHxW68bFow7
dt6aaoLruZr6VDwrMhTPA9oNHbJtSBk6ytMVxrPIW3+gkutx+74koUAC4l+Ftyq6
XOWpKfUqPU7MA9mQw7juEgmGF4CzfGNPzKkolD/nBSAHr4hqiyznIcE/DiVRiYUV
InRv66RSeNdhhTY4P/qu9M6PiOgEoF89o2Awon02PL8KCn4fvb7SQE+nKLOcY7bU
QYd9eK5IBSroAeZ6BC2pDB2MIB1Ci+Y+8Vb+57n09/g/JnHs+U4TmQb3zChGpaW7
8/BSPNYbAhb2+M4vHlIoaHcBME/7XJd0l6da5LvCl+FQv1X5BnvnnVJXjitE4d4N
4Fn9FNBj6KinONWs5swLOsnl5i3fu7TgbIt7Sgvh6e3KjjOlEOQfNivHpvE7wYoL
18bNT4sLPBqpJXM7l/V/hSp6Dkxa/ENIdopY6CSLG+DlGVubX3K3uMhvbvxOo0h+
kw8geJ973uaY0bzblCrYl0LHOffAjfijCSpWoL+L2Dp4OMQKBMj7FqRSfLRdett8
FSi3e8ulP968VC+E/nYM5PkMKHN/NwdXFyqv39NZER0woOf25ukj0UqYAv4DbWj5
ThW8RBfB+tJ79TUsfNScZB1/kiWyL/BSwQnfHNhCart27N7s4uB7NJSH5fw399+F
J4uzmCyoPf58g5BvE8y9P/8flla0RWoS004MGYllcRkrIP/oY9iJ3tMLdm6CAKdQ
DxWLJ3B904CQKY6DsvKHi+FbCZDgUgPcMH3pcDT2ScE24qEgSUYP3pAxmRfXfrtt
DQPg0WutrGwVqrC/BGYJg9RcSP+t7JmY4Tmoq2PUsAJFjdJMFmv/f1sFzkGnBz7N
qtbUG4a25GjTrLhatz2dqIKyd37B4aw91AAttbfeIQVaK86b++eSGdGlUWmnp76x
XjpYyPcBRNsrQXFSgfui9A==
`protect END_PROTECTED
