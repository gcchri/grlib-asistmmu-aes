`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xNIUGFJeuMuDHKv/W684BD6YHH/MqDpRi0Gs/RdE1pknohD43hGr+0XPLHeg3GAG
iHGSkFC2qVwuk10UtOuRG2I1H2p3sdUbM8zafEwquHo3wKmHJLhzQjYg0ltH1saO
y/YlWSPWXfvzrddL25CKSMFxU2/EjqzcAEFXNo033nV24IrcD08QpA9e0+k50DwE
lXaKOwMlRRLmKuZSSHfFq2/A/JohlWvysqXLpzJ0+bDSkUvcbyPj+ojvQIbzfAbv
yx36QRv6u2r3QYzoP0QAUiLRQvZM4hOTvByp6BvWLTl1+IBqcidn+diq6una9gHr
dkT67Cma5nkr2K0bGN7RfCGIo7XVuPul6C8N5LLUYMsn77Ak2LcD38QUJwpCBKAT
lpFa+P04rT/xwfKMnyy7s9k6qlBJiIoEu37qTPEM0+CUQ+fhQsJ1PXYMrrDvsiD6
tKqiOoBvd7A6lRjeCUHoJS3FQJVb6N4oVKDFg1zdyBweBrokQXTl0DcUM2IGG/OH
Ei2fR69lefLvO13DBhaqI8caQ8vv09nzaKMYCp/KLoKZexHubb27IYECx0z878Df
4hm+mnev4JhNEV6f3nfTmH7NIRed1X6iBYpeI7aMQnXeRq623PoE+mEL+0/I6DA0
tyooKE4A9qW28i0B1kpoBcleeyicC8D19UebmBYrGq2lwt4u29Zg1+kEkDvxCoC2
97EyzXlMqntefhD4JQKjB+ZIOQT1uE10hL87mwwqRIifvWmr4KLcpRuOK5Co/km0
dJVttDowhtvGYORO8PLO2+EEtb47HuklNOpcyD54i0OFN2wZV3IS3alcZXrc4hon
XdhCXI1S8ojjVLHF9TmTlivKiZnks61P0GKwLs3bJ82VtfasGNvzbQXQdlGdVFs5
+F4iWqoko87bszDkeN/DMBYk9X3R6BHa5e4WP+TYoEjaHsKu8FIqY8A7FozsyTCr
LQJqzVtiMMzTbkw4JKD30wgEMltvmAhF285IIJXAPbnFpd9Rg0LXS7ah/BlEn4Sq
Ij3kUDCLlizfTy93/II/jCulDjOQIEgwczoanqWIEcNn9gW3fRhp/g0gQRD0xhaa
E/6XUOaAHlIKz9dISyEPYhTMFo283SkoEWCuxiZ3w03ejgP2Y/nBpF/61bpg//5U
wWfA67cwFBg29Og+cVhq50i/JZbD6pq99S2UBzlkzmsY2SXi6GzFM78Ac23357qh
hyeH5jcJxpKLLvvMf0DoQLLuOAhp81W/SwmKHR3DJKKp1atxop98VA42RNirshIG
uVkReD4YL4O5rQVTB8bF0irzkJ2nkuz66SXuMkFNmp5/azBc5Ze4SiaXqL5KeBYV
9aD5du4RgpQ2Tp+B9w+E4zk3qV6nS5StZPhWCvl/QYlVv9o/3zYZw1H/LIa3eoHv
ZMEncOzp2B+i1kGEN1IZ3lmGTuQpekGYF1syxbtTrTGL++QkTg12nPSnSLDbTin8
/Njju7HUiGJJcIBnTMvHy6rPRrZrHN6z0H9jpZX0B2yDXPuK3syId8qG9jPmdKa5
pc+xpuYHSSc2f75kY1Vm3DlPc1y/zF5bku0MWZvJXHHWJZiuMeHIoi1ntvvT/kW4
SXtqIJ2Pn5J8henHXWqQ0KSC2lutRqJ1wR67NP8S1OQJVWJduTmmFSpZZIvI9C1F
YlcxqXcC/mi+sGirvZcdkX3HmouRxLkWCeuKjXBDt+2pqoducEpsGgAUE85x9j46
gRZmOaYT5LIG/F1MMCgU3bvfR3sOxWXDBVaRnP/vo+Wgpe9KrQMruMmAOkV5AWHC
s9RUx+vxC8UpAATtbQXVPHKzulQLQBelvpX+m56dvjJGguWkZa+yJjs+pMeSCNkb
6PfaXfA5N3eK5MdxIWknXkSg1JpFOUNPQSyZhnfxlnO0NTbj59/Ol/xtepUTj2W6
eyEbwXj7XLj5phenRpd+XbZugTCKG/jeoOlOeek1PwsmxmXinABWZJmBH2OXD3gV
BbBPuRoHoH/pXgy/fsZDxAxrH6MvLKCN8ENXncbkExSftYZCj7OqHVWqixqaXq7x
LcHdknxPZu4NCwYROU1TAXByKL/1HfWoVXFVEdh0bEKcDtP/OYoJhWXVnP/Jsp57
qOlVZZAsNVKIT9cQDn9A69NVMRJNijot23CPVgyzV3nCheGzFFacs3X/c/+xYkVe
obAMPdB00OWxYjxrs1rnOZ4mTsB9/Om5EsY7OTIbP9ShmgjKcRaycgYC1pRFT7Zs
K2p8JB0I9ui9jraMqvECU+wiDDClXxYXggPneZaA7t2z4fUXcRlCNu/1PMN5V23s
cC5uVZeBl0rcKTAfPpmG4O84hAMuoeXxGuq7PKEcxAFReIKaW3fmjFURJxla4yMV
QCKQUBV/iINfQuNVxdoEjJMq/MhfOZ7iRm1KWSmdF/BwM3YMgpb7DOhOgf/JWqkx
UvZ+MfuF47jenXkk3tSKvde9ywwkGGGvcRLoMC8H3nQy9FbpVRDdd7yOA0S9ItV1
o2IqnLYmu7IKWyBOi7CAC12wQKRoyJ5iIjv+9VYP9r1wsXN7UxCMfYrTQFJF5iVA
n4jMw0RpnoOmH+w3Eig+Vl07RAZVH8mnSAwPBSn9tDR+aa+lpYn5UVvpbJ0BjlFi
4ih9NfG2SxBC0pyKyYysdtBqzaZG+HGYyO0fBX3SZUzAO90PuarfYV7N6RoKnc0q
iJo3fWBWcrFuqWT10Rf2pf4TI881Xc8/ZK4h3cttld7zf3/DmmyX3m2T2/ghurs3
OwezBo/D/EdMsdTBAaVFPHJMxzkZG6Ei+BviIK6wp62Xs/VvpOybPmojeQ6+WMbU
YuY3X4m3HeFsCISSMyyvYEkmFLj3wmu5JWs+5+SIB5hz3kNukoyJQ8v0Nb1uows3
jrCHYDy/YnTFXRcJsSmdCEgHDd36Hp7htK1zjQtddgszdGKNzPHJLZXxfc9hrTjb
Kfp1bFpLy9FLC2tlxUPQU1rd1Rxe7BB9XOG5YnZBb7MfIjqxIVcWmZM9r4aRrQrW
C0zclStZe9R1B7lHfAM+3sMqwW0RDs/yDeEZ0Z5PwgKKpMcRwte5QbSYryODG0t7
`protect END_PROTECTED
