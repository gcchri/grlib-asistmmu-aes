`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JbtXfbjypU4T/bd1HJk9y+dYENK9PwrbKdCZQ/4Bm+0Igl4Jl/UtLY4uejnB3iDz
p3WTTSEh+Oir5QfhPx+6egPt66Ky/B7R9QK0cKy1eAYg7iNMFkzAj640Ulu1tKLe
Gx0rAro4P4WLwQTryjGmtsXlMDMuVRjh35ckEv8h5GMxZOXTpGwveY1He2vQKs9i
U/VtiUnFHD+sdxar4y1Z903OeHu5WHj4L//Wk3r7MAhihmuLBS8cD6YCxO2qeJj5
lLdoHTJYwq7YLpf8AX6JejxjkvGUnczieUcFtKuQlrQJC4lrqoClwXhw8yHMNRnb
WYmFH0XUO7nP4Gj9FMALvmXzUhKXbP13UVl8b1KtyeYM++mReMHYKIU+ZYdqwKOR
VNKhXNj7AMVhH3JBMO+aumnDA5VtcycdyhuGSgpeWIG3MvNklfT1inZ/BxQBM+Tb
62evythPPzPgs3yy9ET1sUboqbYzdOQHuHB1tiOZ5bqDa67kJBEErGPn0zROTozY
zdJJG69fUzFW9YfRFTDO4RJ1ek3GENZiVHWkaygA8fmST5HiXj9FmALUaTKagtYW
J2U6YpzZ2o3Wt25pXZGYnVMVvexpEAtEYgOtprcEGbtmaPfCnZEHRsgFWt3eLEDD
kfwqf+uhnZvkaJZWx2gVgg==
`protect END_PROTECTED
