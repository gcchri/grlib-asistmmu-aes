`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eX/BXQ5HCPY0Rsf3u831JZXg4UyckfEXoIi7MpEYWjtvRP4Q0UEKRlss9BbAAVat
5SR9uVZmUPv316DKl5W9+iusASx0PBjnae0G4cWGSdF8sIf94+iHm4/7pr4S3ydT
YlsKgi9s792o7Ptcfb+3IJg87lO1hFV02EgJf8BL8n+L+GNXGX4cl/6tkvcUweCo
DKSrAKpJzbGr2VpuHeo3uu5qhGm8sSvywGJzm8DKVSkexbzrPKS5bzc7MNvHL4ED
z4DoMhiOfG5wK67x5cI2ATk2cbP9W7P9vUoqoOzz6Dve1KN/rLQxZudDLNROz8WK
ISGmvEAQ7KsMVCc10FS4E+1HRVI30GpWzC63IC4zEpA8tpkfVweOc0dSYBsZX5iv
pgdQrY8h7sDnZAQZdW99U96lRotfekJDI5YHbwyVYSuIvlfikDbCkWWMtTreADKX
mJCHflS71FYaxGy+iGRpoV0/GPR3rQ/LFKDKC6iManxFcW+TQoWieez8YCwt6oUP
Cd+6xLbJXiRbrUSLrXaxHCMqtbFmBqkZv8IT8OTup9pt3/ndk+iz+MT/UPphZ+VC
Pum9obCzw7RKHtfyZnf3fhlgaUjWzY/FyG9hoT+r+ho=
`protect END_PROTECTED
