`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qtVXkSQeZPPysoJtUtVPZxhGcMD5idfzhpfH0CK0LJlMXyWDk5iaYRj2zWBAsq4F
XAyHNr33Pk0AGkRctePzm0NQkqSoJvyoaMM4X1LsyCkd9yTyHA3aGEGZr4CCm12w
G4yb5a111k2O8XnLtEU0V43GtcKi1td/RkTNbG4O0zdC8O7cBUpGZYt4GzOmK1+3
yPI9h5Q+OZBr/DxgJdh91t/UULuwM+BPuOC7bi30MMh52xI1j8y7/8aQojwd65ut
BqDpBRVsrXhQqkv3vUy8lnWLQSlm7qP7VEVyqH5TrC3rfsQpSkiZvF4qORPmEZ+W
gZQKDRgGJqMW767zkZpYHXxNtPJ03xYtMJyPR0fQxFKYhth+aRtUw4iYJ1gOrSif
9kTva2B2oxRaz8oqjWs5O/7+Cplsciw3JA9sEGvqhGQ64dsT8WI2slxYBz4BPg4a
doNAL5GKaiTTEENx9SY8BQtJPN8PiPkG6JaYxOdZzkA=
`protect END_PROTECTED
