`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bp3h/vmH2o8LL5BUeMqJH5ltNuyK4vd+ToG3MAggOL2+onr0o5Ezic6C+tiL1k2D
fz3NiG6u+g7ERyTrO56qLXHVo2hY6tLHSwCp4cIg9wsTK11a5YT8nIVWHQdnGvBM
YTyjCbB/fgFZQP4H7iXz1uDceNyAAb+64I+oybnN5xy5D+eH0JSGfRxCRFibfrXV
AH1LbCnvi8yJWGztZmFOB0MIN105qhZPHcow0Ve3m+0pszq6oDG/gKctvAUi6HVE
uOHmstwl7U8jYFzpg14D3Tqqf4xUX/SQvSrw++ySybahbvioEOdm3g7pAKvEO6JC
bc3bhpwn17hwOXvY3oaHaoJVP2TuXaQAUuwdHgR/7Adtnsp/Hc8uWoz1s7vMKC2y
D21j/MQoxiOsbd3aLWN0wQtJHbyuhW2PuJpVAlI7PGtQ5/g7Z56S+ORdc8hISC2S
WS75h5WsVkqLiBng7ug3rFaDT4tSAzynkmKLgObH9MsZQcfa8xhSHXJTqDcIQ+W2
P0jBFeiQQ0cBCmRTk8aNo655XsNdVkJ0CUE0m5srnfzO80yekMYq+PSGndnl4Lbq
a0Yho5qhHDh1hWo+6hedWuwQsGemBU4LWvgxCXgCis0JkDsQdwZLFRllmW+e0Pv1
2C+aDLHCSi8Bio38LLOCNEREJ+gFZKuv41odwsZAJRZV/6I315mPppMqaC9m2pqI
7pbiv9/MVdwMyeZEPiPiF9ctfSzo0HNx5Sw1fqv2tuxCRNCwqIFsxskksUquRgSn
Ct+b77ejYxIrp+0cg15kTwGQ/N0/ob6Ww7/B22qpvHaY/uN8vVf/Fn343Sm+i1wS
jToBnQQOfq70gw8TFUW+MCrinuoqZ4V4jVJkpkdXKOXgTFdynzsqXaUU53g4Cmcz
Prg9Cz2wTLhukYXv6dXXXwGdgX+miw4TKiUl1i8mTJw0jJHqWSSQ8zqvfJXxhOM0
LF4cU2ijm3e66OqVPiSB6w==
`protect END_PROTECTED
