`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TGAcLhdyPn1RbbcFQP9p/AxfRULYa1fwLbMdhlM7AWe7UMcnUwAVtL2tfXCrgEHi
iRcWpIvY0W+Fx07JCcmNLTvPcQpT5hjCnjTd95y9WrGWuNXr6eB2o4E2fUffMz5p
UZ4JMAb73DUuRfm5CLOj/Nrin7HyGK3FU8YLOoQlrc8AsSEFt0OTvntUbna2LYiw
5yUg2xfEPpToEwNqpSTAHuVR43xU/mGsJvGnFlkTORIalHTkX5HfdYHzlFImjC4W
a9266noYuRGaRnoJbEXspJAVq9Xq1qywRriT+blqZrO2uBOnbUvLQ89dt1SPC6Vq
McAKL7jWAPx4GHytam1Gx4zWI4VwIJwjC/bKCd4jfWeQDltcWYwInXPCtQ5q7N5s
UXTPpsCxvOi5sc91DIIQCKnmeftUKFmBiL7oZ2zRMxX2Tm4FvPGEx+cLNnLpYgWX
X3xJI/S6PSj2sQyDttyuS+V0pgRAX28owYYxArhN5Imrl9KDaKaS4PgvN2zSa4Bh
u3C4HkFy+nf/PCeFFK+xAMRrPakonqKlmJp3GvJL0ahYxXGyx2nUNxCwVffHXn2w
FQmf09nyuhQ1KAXcZPOAM4M8m0Y1nmfuJVRty6zvhSqFMTPkA9yCXGN0MADDa65/
JDFwTjlMidjvNoHMWkbB9Uydz3wuSCvfYd6YFIC8aRwJiEQjcgeXn4ai3D9P/CPA
p84C5AIBHFSa0qNAVOijwbSfywergiF/pkXnQNSV9nZC93yUQ9pkezD3eDYvVlVM
0Tc2dIpUftBJ3JpoLYI8+vnW3qbNxwcB7a4adg9hCmru6syrMZWAxhhL/80Z1y4R
awj2VM+AlGIH65fz+yvYYus7NVnUk4pmGXowe3JCVTdAMJtIlIvN89WZTdxb3Gw3
6E1ALcqAyuJn4dKkDQiEWhnz26bOUq4ESsIlximLvaHzL8MMBJh5bSpgPgwBcOnG
O57BwqPbyvg9Pi1p+qKSs+jN1+vKTt914hzBa3VL5bkMIWlkXarM6Gr2y0WUkHyE
QnBfK+uS8P0HzH2hqO+VxYj3D3toQ+kLoop5uSgTXfp4A4AdcLi3Wnu/VhlNNNYT
lkwWTxLWK9W5M/kNVlnhNjEELrk9PTHwnvEhTvgyBfuBzbP+9Qd+QWI/M02zStFM
RcqCNaff3g2++jdoNT8z52vdF7TzZGjMGCi7nGqq+FBJr4YrUrLvwVJlaogu9min
k/Ap0aHH60wTV0JwUJkH5Qt+OuMMCeHvMaoAC+t6dE2LtPYB2j9P2DQ3Lx2klwr4
SjEWWub0zGHqN4vXMljtAMDW/3m6BY/LQDOmrNwuqWOQgJm4/5B+pvPvh3Y/dR2B
OKzOAcgiZWgQpHfLL9rWT2sZVgY4oeFaLh+L9l+k5Oa1ZYekTfN5vPbo8yudnMpl
GqyAQat4bH/LhPmY7J1t25/+RzzFmtYivCIk4IqA0BJL7wtyciDFkpfw1LkeVizw
yYoore/1YcSUa8N3cyzBGSMCRg/AyzmFI6giR/Psc8gJwSRdXL5CzcAFfEIK4sfx
21Zz2nxAEoIOQBwR6poCY2lGksq88eve5G3wZLjAe2LW3qOYbJvzA3jpzmgff18c
Z0Bp5//2e7hdvDoBclPQTz4L2NAFQJAqvETFLG6mLPeuEfqCaKNDBSwUwh+Uw0/M
biDTHeG6/DmN8jguPyAblkJVfNe/qrIZaum0UcsXIBiZsWqzXHTyv55JFpuGFQid
gw7CL4oe9vX2Prv/vuC7wBheeONloafdQnqcR47+Hmh/cYrLveNXC9+13VQ4CzXO
h/NrGKEATvhbwxSEgsYkygWgFfdkqz332yE5ofZoPHHhTWGULbXLIoyDz0GvJDOY
jjwjkI+Uc0wFeqRt7Vi591ZhSljCn8nfCNAe/dIIGi25+Rt5e+B0x/ufktAejF54
H5UCd9u0PgSn5V2tLhP7YEU87RF2nN+L8tFlmLJpngWBLFa2M9FiJ0Fd5Z4bHtt+
rjFPT3EX5VpKM9vdwffCtZJVZHVSqNLF4o6tpCRHjXQMilhFh2n9YDYOTB4NRhCb
pVrHqgahxoyuJwrMFU63JXoFQXhtBA7Wwb/dfSsS07qspTeuCZd04dSXSoVlLdFv
nqIeDk41HjB9fbVBLTK/acOWhE5gxSeQ/Fikoc4i/WphDzocrJgt6oOHgJRPj5dq
pvrU/Wl69095KWuA6JRYkH3w0KG5aXR6Dn1Pq12n9HIt4UK4MuuQF3EdzqS+nbOz
6kRFvgNOwV4errKfO8s4XZrurQ+2ZtIipBDO4IG1/OZJaTiATk0mg1iUhZAMyHJw
NbPVyt49UBNpGQeVbmNba/bAUOjVhtf0x+lS8dcfbLUK416YgXv/GsSWLMOuIhee
/c2T1z85fIaG2DV7FD1lXk8u6FpQL8eMm2dyL23F/R7P6J6NXdYF05cvkMsE0yV3
4y/WFfmHhD42GEOuRril4XdKEOZrRlXLVgkArl1ylqNielTm0/6OtMOSdLxT0BMg
/3KPVbrjJkzNBWC3OXKfKBZj2Q+XL56JCsp6Ri7LruTfPlQGLbV9v+7zHslp1SQO
ehgSmfHUSbrojaHUTIDDei0b2fTKffdBiRaIm2SFk+TFrj+1yTVEUbqHRY9T/uNc
26oMvmVKcLQ+wG+dyqrcmc4Ufuk6k/xoqWyosYcNUYbuvAsqUdeIHBszq4xB80R6
FJCLgmzdqohEg7iUY9anvzOIF5CSQvxzg/uQNr7kWLuDyY+TeuobkPjfJ6IsklmR
9AE76k5n9LavxZ7cohULqHUXBoezyozdgbD1c3qVZoedzfX6qm14hrbxsyeFLS4+
f3NnKcZfGtgsdBfwrfclJvokW5Kq1BGBtlRhx00QC2m8lfOr92ScDW1/BTHurmOj
ZCpUcGGdtwLaQs4w7waenecaDqSnn+LsvA3JjpIQaQKqcJTFVydekpYfjxTaz/0M
ZKrpasYT2ypoB+FzvIXoV273qNMyIf2LCuHe17NNNLGkV7XF5bEmvuQitiXW558z
HAuQ+l2VIANfO3RboiDeTB++qUSzDnGKNHFaQ6bBSFfdQ6I92+eqEbOz6aydb6nf
KCQdmGmseiG7SJk9q4d5u3EJdE5QCAllzFkL3u5FZWYhNI6xg8kcE/kQ5eFf+u5h
5QELhF8ctlZCBO0r7jix8po8IEZfjzuMjP9z7F4viJqi59h3xD8zqvhSIeIF9JAf
4IoOUBKNOUbrtW1wMkkXc58BDyEoa8EVXbM02hcsNaBQ1VlIeveyOLe0B7ZENgty
hbbo4w5KUkFc3t2P8FVG1+FokSxt+lPAZAxBaIlOVs4pEAq/6OdCpZTqrPfV/gWb
fryDt8rbIWF77+FCLoOvrIbpEz0kEAiOKOdNA9LJX8vDtr8mp8bsmJihkOl6Imu1
yMjS7GT7PkYTfr4YnFUR6tKSpYYEXV7GGR2htl9JGzKTjSFM0Oy7qvkV28Wk27rw
IXDL2FTDy5sFBdC2CLXdBw==
`protect END_PROTECTED
