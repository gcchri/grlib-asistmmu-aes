`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ohp6d1ZS4YQJYBru6Mu1e68rEu0OK689r+jGNzgU5zPbUt1Q+vLXsjSjGgfpXERj
nRos7HMwaWLK0wNL+udJVO4j1x3anReQOrjSvYCJSq+Hqbn68OEefwEk9WuV013H
/dOXGDDVglEADEsEZUkJfseoHJogAiRD9H5usg6cbgJb4+AuZZHqIZ60Ulk2KxaX
6kRdUGVKwS0myr0kpj+oLSorJ8cRCLl/oJtXaVXxwKwNRN47qXPYovhbAcf7mhhj
WEHbUjd3zvsLHYSFKa7GrhjsM2VYiSxbYPgY895zfjbslvHSKVZ8wQ0KOgPdeSQx
MnpKUZuWYp0pwgluRbi+c0vcHhHPrDERolH127TZbKP/Iq/O5bjvWZpD8jKDQkhu
/pFH+wkseLmQHp4IqBUQ7mxKKvOuCya1WfckCbul275hUCpac8JRNzSnI/rms75b
QSkY5G3raGSG6aKbX0kxznuXuG7lEPd0/HQ2/I0zhEgc00wH4wJGd9SWp3Sz4C0j
BUaEFCcPWy3n+gjJJoPZ00m14Ba+kswT7QKguFh34VUVgwPAfpvPnEwnrYgBb1cY
RzkzHcR6B8BYRbLnFDgzvoiZyynNjKW7N7+HCg+aEU9XhkQV3p00CwhpLKl9WEmu
0JuxE2V6ZZ9lqTZRjJiTg9mTm8zIHdis2906manz6YpzZXWd5+Ncqe47Srh/VEI3
ON9uQ3GjMpDj/CEoe6GYamIHM9x/FWLUr/fvS+uoUCFN+NL9b7pLH7t3xtRJyaXn
QBm7PYmBG2ggef2/z3Uw7UuZihGq5BdPP9SgmSEhx3Gdy0UZZedGGV3+WrrKhkHc
5JDx7/fIklA8N2dAikfJFN92sPduWwtLX0QLO6i4rRvex54tP/v2HL5Ug7c7EF5p
2mzsC6uD4Ry4BDE8ScjLTcMjXG+S4hx3Apx2Sxv9QJ3JRF/5NZGEYvB5LEvLL9Zs
EXhTiOv8R4e2FmMq3yaXcFIEefFXL96sC+fqH57wNp7o9vJmDdrAT8JEsxz7DYC4
/bHwlFJVMSPvjubBvFKdqISxpM+JzzbO/TqYJwoE/Ytoqh0oMA/OwjGaQnojyIGM
0Ae5mjryYCCYyRXd3sW57p51FbMGyOhxIuEXFvYIFbcLFiXCLnn5IW1RjEwNHB7h
7fGs19SOf8eMcEncHYq5ochHAUvu3NChhX3JE8T8iJn8hKCerIH2rmsIQlRIO9RU
SQ4c8eCFneDNYEf9y/neKwdvP8wrQIeEHr4pvvmFrGgLyMAMvlv9NcebeFWq4ok+
`protect END_PROTECTED
