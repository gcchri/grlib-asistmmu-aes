`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vsc5K5WKQgiZlePQx73PpFhRcJyxXqUchs6UHbjw9Ya27Cq/n55td4jBa32TVIFe
vcFENWo8U1Qxb0ZqSaSmjKZ5BdqfaQm+sD/KRcONHFDrXP325oC59JFTFgn3aaRo
3lGMj+Bn3vLX231dbhpU2jTcwRa6zS5UrzvKcgw+MZAviyzRZGb67IEpFPK3Fxx6
iM9mAEGc+m7ptrPbhoDxPN7ZFVYUoRX+LISbhg+PzjjuLs79ktjIdij8P0bdXOY9
2DWrKi22zLthAPbGd1tw1OYvD9EpO67DrH52JcLvjtH1x391sFwA9SPVsPnrVUsJ
WUIJCcGBZzkfHx4dTuk2lybu4m1jfTGXfIzjqa6jbe/StPV8byuuIhV4cFEfTy5V
fgojPLO82Et7F9YZTP1lalBtG3PZgjWVS7+1DRGT0+uoA5eqEs6vtntOnhuKCFb7
344OF100N6N0bDiaKfIZOYub6th4pyXSJZln+4rbElU=
`protect END_PROTECTED
