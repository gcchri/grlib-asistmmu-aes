`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2VqWcYdIdDNL6ZBN9mqgxmERH6MOqPxanBqpciXm2p+xqeK2FH1R+K3pLaj2mwHb
dshVEbPnSSEw1kT6iXhSpGtayw4f2PHKdy/RmoqQp58uOJ4khHaU0T+Ii/fSOtws
sGz9KD1BKAMKDEaUtNXKzaibeAxMuhfZ2x4nW0OUFGiM/Tqu3CH0OPCZ3hZ1JkOt
TNXxMkXRXsy8YTE8u5gnyYaLYKlpXDpbwn8gUDW/9qVJBmGPOWA5nBcOZ6qE3oHi
9MIy/8eCPsqz+fqLWw36uMJF9nP3SlYN+4GcnSmH67yJk+dFjHG+YXdnfoDl3Oll
taTTvOPy7L1PkZmWcEMWwtbog6+2IUGUWDD5Id1PNb9JNx/GJEDR6dInmZxYOSnc
ww7StpEgQtESvqkwG+9+xyGBVWkOoJewF8lX7Ul4+p+jgBJZj0GRWxzDPQOA37K0
8MJYSS9WjVlz/NwR/MLn4A==
`protect END_PROTECTED
