`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bSTHNIFRZ4YNmf4YfhTfZb+7R3Mc7ECc2LvdUw93mBPZ5o+uIcVaD2N5rjCe2DA7
YjD9fEeHptuwvicfP4KHsPdnDoNO9YEnDq2YCOQNcJgowSgMks+Wjcmmt8XUrOds
YrMLzyEq7LNSMrnZDVLubnCZdzxaYP+ul//YcLeaXMWnvhSYKl1KnNhihmpjsToI
W4VTfb5UvoCkrt2JE5J/6vD34e/yifO6BN2iqhxU8ukHpe8W2FAzgZ66Dokfl7md
LN0YVnuBSXsHiMDQBrnvncqF7CeZvp2AdnTHQ7XUTCYuw+HmSpyvYG1NPdl+xs2s
PRX7TYFLgTEaOllt5/NsmbsFIuH3atVSAqhiPoLrd6D3wx15rFyXDUnKEzmYI1zK
sCGjFpO6FBVdIdLkmDKAABYttTKWtc8hZuOh+d0YUJ4=
`protect END_PROTECTED
