`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JtkwMmUN2OdNR54ijFrZIvPTXpGEmmy84Pamje6RxA0Fyae/6KXeQXj34ETQe+Rl
xwiXMZiZ5s2lamSt4BiYDqmgdSl+1jsze0Mgre2fwkCny8BZvQ/ymnDhaDrC4xio
DkaOc9MYQSFMaxT1GdsDVXA433kiO7XMe2l5tNEoTfVkxZ7tc1dR0VH/4q37E4cC
0wHhRw2H9BLW2jg+1ujUlPdAQjDjPO7+XOdhhGVuBr1PfO/UoQKJbBCOFoxYtxXx
kmWxULRQDOG5A7UdloTdUKcYmRakJCIklYzo501A0DiUTvnnr93/82UZCjShM207
bHua40Us4OvjgxcIV6I5PAKUGGgY9jGGVLFLy6PF0cgJKfOmgPngRHzWvKAeOCa6
`protect END_PROTECTED
