`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
exAjuMKpY/zH0b19M1uWzcO4zOFkhT9pDbeRE9rk8j/Mu+Z6SUWJ0/bpSyKPePu2
O9g9ox85ChpU8LZ93I7hndULodHxNps9jg7j6ZOmYPNRk5PBYij5fnIxRYmrmRsm
0nv/LdTEOGWsfqR9OvZjgwIHggt6rGHQ3Mk6b+wX2VYq04iD8svffrudELCvd+CT
G/DS9yl8ZGKu9UNuflHsVyJGBC2deehkI5VO2es9LAXnR0RxWaTLU/Tj3n2ETJhV
O3MsvTyUSl0IgbYv2xBrG7gRnqt1ITdwDpGALRRFrVd4+K368h80+BRRy2QEVv3G
Fo8VLiN1/+JVbkfJp+YQ3LusXYmLL67ixH92A5Aflof8eGWJIT6V70Hv3twcUcYy
0j4BpKUba/ZLBfieUfbmdxgJB57E4W+1ZsCaqk+SUytAz1pME7h2m45qc9E0e5KB
efnrQaM2PdjRdMYlwv9A1wjGw9XxRyxA2ZSPM9Zf9+cXmNW68MDl0mZrxTFf5y5E
QZhCbCTBvaP2nbxOJLlKjIyFsqHyi8VdR0rNZpOS7/Ln4yHyXFkQRyBXKnMgqa35
lm9rKUHKH5G6xigEf+BeiFS11pv9VrkT3rUqRRgsO+EnV64sm2qD8NiOpGtJyslu
1ryE8d8xntU/OO93/qSzQhD6CmlNSfEHAltdg9cDZaE=
`protect END_PROTECTED
