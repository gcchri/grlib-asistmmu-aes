`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c9h2pbg2AAzV+lBy1XShf1G6M+LsopUAAwkfpeV4V6YFPDFEgb47eE5oGVqjGfW4
7t/PRVuzocjFY9zE2GjBXrLKdiLccGPsQ2PJh//44UiTfbN6DXWkWGjuX0Vjr6Aa
6pZwzJIjOpGI5ykyL+1SNiGsczd/HMDYDgUwzvnVkqn6aMETRPN0842hk0Mol74K
K7sz7xt0pRVT1oqW10b8/O8qSSvmiarEfmrBA+uKjj4hqfIIlOQjajkm36zDIPaR
32LaaS1tjjvDHkEWgoXCt84xiUNgKoCB2mloqOng3yx3w76usJNoTKOyIk/U36FS
Xtqcpnim868UeiDM3wEeQvksS5pEuKAXx/CqSvvFONKnA7hgXyTUo6MJ70EOQQoG
eytu+A1GdJrywck9E16qOogkEpo5bjI6WJAlzsiJ1eGMF0v5+KnRmDM3jqgkACq9
b6h7zpYMCBlBTLBUtWCpSo/or6blY9k2CSLt+teAW+fo8kZJcrcGY77snwo7STm9
z+BVgUo0EXibBPhzH2K43GXYB4wt1lLWWPRx+Zudo+KlBkRgV9jmBJa5YfYBSd4U
oqHi9ScYvLPUbtutOJSyXFkWoZymZjZA1Lq0/qsAnWXvBXfxYQmRXgJQlaXgrIz3
pfpX04/nEUYMwgmh8NeepnkD46RRxn2eDILtx7emL0HzGS8Nq9TiKzFyse+CnkhK
JSbvXpygEPPxEV0JuLk2hHU11UCTgHKRtM1SSgXkUgA82jP9HKFtwRFAeRdumVxH
GwiG2hHeCAdzLUKIOjNIGlZF+z9L6K8AG62FuVKyjRjxWKW6Lqtfj8FU61/FnpaQ
NcdB1G3Ay5tUhM+4CoSdbD8x//ZF9wBX+rTwW2hhinyA5LrmsV0mPmzlD/FeBb93
hEisuGQz2qlprkC0axSTH4I+SXZwR63cqWan9TPHoCKZOEdXcDCgg0dCvyB0fiis
g/ZUfc9R0VRg7vUAwf7L3EivI4kV1OtsQbrN0dFPj8JjThqQuCvnQ3GotTq8b/ot
QxinV29RTJzNUyr4FvTt6Eccrm4HIu00QmafUhuuC1JpWOnKoAP7rUM+BlJijRjQ
TybRPt69NFvQ2vGZRhC3AhS/h1eGSlkU52R8QuloiRbP2D5ZwPConw+6bwveI9bq
5bkXdV41KbBurqFIwUrOXSJcMahj7c7Ef+e4b1t/KXmmakoeIouk8fbWDZ0FL4wI
gqOtFhAIi+8LEf25NJ9XYd5drlEvsHISxn6vPI7wycLD4giDfol+lZ7ia6CpSrF2
Xc7oJE4OiUFPF/eElC9dgM8FcPGYVCOdZ+7hYy+DqY03CRyAXYedxVsOWnvbLwmy
OwEv4jsiGJYIGQVYKovkcYIh/6Ni3vb3hOJj84cZadMd7OfHiVw9n8fEkVfPReRq
g6dueYXfEWZJpPqtbkL1pjE62Sj1K3J0xcDNPfCF7QsFArSbZp+gdkSKj+oxGEz7
+k7PVqpUNinmQSS8Dk2ebm5VojWum2YnvkDKkOo3T1HFVlKtxtViOSPF00e7OiX8
X2qOWBbo4eOk7zI/2fE1XGCTKZounoaWZTbDuPEbASXOddDMAw5IAdyK3NnI2QzT
8gK4ud0rR4qG0x8Ivfm+3fAz3k4AH7XfByiW6cwss/lCE7drcaoK3yn9rcmRceut
tbpXspW+oMpQdAyfcPBsZhdF+B9bIam1W2Woke1hagWRS1djTY9AzTG56IRJbSGE
Cx1z3fsbxl+7nlRUviyV1g5q/ZqLzpxlr+2IzgR8sSwtGrHZi3g91thEw8FgSs+1
r4OiQlZSKiLG4DnB6ijQtAn02kgyzosmGTM+K1/H1WKX2Qub43MpF4n28NbVFwzM
YxQroQpiV2xjg3TSD2JhtWC+vNodHYdV5weOIrhMSDsJfg69rGFjf1k8T/X7cxtn
zkpWegJNOp2asOLyOPzpgaBG6Ew/xem6V8dXqOttdsl68MWVGStiad3f+pFPiOQy
uPWnV1WCWEkw6tnLJo6KFGFmtQ2xyUPLAwP4ZjqVaOqAeHVXWna8i1frpQW+XYUo
ccqP2sZpxokfukLvxSl+pZiYqF0xmqSF17IOZVPK/1nfpSZjnaMRREmRU96gACuZ
V+zWYRKmX0nVesHbnER7lPXKGuGgM5zqbaLIq+H5ahnJscH79kj6PCqUQ81sCTV2
3/PRqZ1t0LyumEJA0ib/EcEMgseaE5cVsY6U+zbPgUqqEYJa0S0OxmHgEhqc4Zco
ygC14uVgyZezojRuVNLchqRhWA1RQaeRSUzgC1BU4uREbqMA4E8Y7PMGFxYd0/07
65xCjO4s6beJ8vwqqWEytQ6UBA5JlJeFJyoPWsJkOLGDjyBhhKV01/vYte3VEIIc
8MrhQvQBNx/eIUCzLTX6eNOiFhZTd8I59+JNGe1JRoOsuwWeG3D3zHHxM4p+tG+j
/wg8RQbNe5svvevCrTcAPoOWNlYa3r6EA+08l7m7iE+UorZzEx6caN82HAbshM11
jNg5Qzg1G0izgSPhivbN054/ALWTp/8Aa1RJLJM3K2r927Z0pgFjjwk/Nn/Gn5+o
KcYF8pYTCwpFbpYytXw0FaxWSnQHqt2hBJmEK30ChVCWuJ9oTHxAYXbfI6ac1eMV
SoekiY1Efp5av9WhLywQzPk4o1sWz8IiPepvEBIG94Qd0SlkIdX50Cd8h7oo22c9
2udGggF85G4vqa2rmeVqKLwLq9wTivBv+ulUQO8iHru9outABFVXBveBVIzdEbUy
Bib5C3qCa1T5uOVN0Qfwhjug0jRQKDSpWngOPz6LNp0f307l/XbPpDX0flf/u2qH
ZHUVQUDDdr8JVET51Am5bw4m6fttenmLU00GT2a2ISLcvE09qzUMbDKpYOhknpsW
Hdyv7g6D8NEKGGV+h+nziOxfFJJ9kx/qHE6klMZIVk9upuH5SfakRb6b/ts54aAz
LkcIql4VHJX1zfQGneqMNofAddqLbTnGpJMnnTx7eK3XbSWFCxR2S2gMZnv9GV7/
Pw3AeOTwkeWfv/MgqxUhT1xcOooV3zz2VH2MhlTHQlS0HTkYQnZbFzlt2n82+rvW
HhYy3MpyuGVsJNsxdKKzpTnzgqGF93xxi23rXQZmHT5OYkKSZzHvDhKfebuYRHxx
/NLw3lJCCHpJ4/G/+lax+NjlWoOgFgsYNBMZVp9zJFdKWPhywrmbWgulLMVqh3aT
eOGTacryNBL1p5SnPHDXk9uaVq4QpHSVtqmBSbeyJbWGISgWhjH5aPSXSXqGgr/K
rBp9TvNYF5JDgJwwci/YM8zdfHuK77wj4EKRRJ3GvIsGcAxjOkEknm1mIlW28MCk
uDJGeb2pBXafoaj34yvCPA70YYbaVsyGM0wkf5S8YehuTdD4eFIFLOTs1CKIms17
KZywj9iSjZDm2V6kcW3An4EBBFsVCt+iZJE1QoVie6bQLfX3DJ8QQdVjSWlqlEJp
S3NPIW51Ob00sUTbxhbW3WCyWuCGVSNB3IcA9tazqDQXr1slsL59jvVfexwsCoCR
/Cey6oClTk23xaSPNIpQIIAkT89rt4kewLt8VeT+QAftXesPUUQitiCySyp8cNaG
dAfQLNqVs3o1uw9Us9n2RX5qBodbZEPW/N2uNXtAqvr1KArQOQPkeBUdJcfcPFSY
0Ju8+IT/XMwfp+1wswDByMWO4hhhEAOdMlD5GsUSLLvW4hP7efYHePsTS6kC10Kp
FrVVurSptnUT6debjWbRXIGWiexCwLmJwJ23oL4nYLlLNu5IF9QC17dKYpSbBbk1
qXnpstACbkE8iTJxho8fY7LRfyFAwgPy+Mejn3pYRmTmNZbMCvKv8/XfjQPLxrQP
yGMV8+Xu8P69TPwRPVTAsUSVFclVlni55jwZUyxlgR+t0AcsJINzwSGqb4LmXwuv
mfvHoFy4CFWikZCFmMx/4ZxHXvq/uO1Fb/8PGfoC2hn04Kk+QWXp3zghVLyvDhrr
R5+suyvBLpkrYUIQKjLpsPwl7R8eekZNfHolUPeAOlFBef6po38UZxj63uiZsAkN
Vj6xD9W+PI44051gEXFaIh2gosOAeIqJiLlabbUtP020dYKY29mo8uu1JgqyE0Ck
6UIIP7Wy8uQq6K0yQ584alEpBy1XzPUYVifDJHQ43TK/+bd5UjeaC8tH9FCqyjHm
gou0YaacpmahsmX182oFPABF92cRviBx7SxilUqDpL+3420l9I15LfKd8Ln6gYR7
xwjzfIFC84CgT/0PlpPsXIHUOCi2Q73VgTBUMnjN3+XXqyVs41V/6uRunAm9pIHG
e0Bp9bIcu2EtP9HaUhF0S6NvI+DXbdmqDPXW6V2EDExY7DS0d+VqDZsHwoCEM9LE
SHSVkb5RXayV7OfEbuf/EuM0bAiYflt1VCpLbMwmYEfaa1zkkyKtYS44vpL1JPxz
ViRdJrXuF1VINyDW1Krhnx72C+gJR6BPXOi+6euxFxtEqDcWZlb+JqARewHz39mH
A+HrDe1Az5gzBeMTBvTKyvSNnva7u6bHJjS30aygUKLoVoNWffUhJu7VJxACwhRt
juSP4zC8GxPcwJ9/It1fZGWbWABFyUEy+ZveTfjZxh6s4SAA2MnZW2tZo4KfhCV4
RupRzLIW9vVvR9a2GumpSQuePf3C1GVHFG6UjetqF0xF9mMxfWK8/d4tG/0WSYJw
pODBq+heiLejiO7gxnCFaPsDt+OE4iYqSJQvuBlF8UM5OT/YtzfrlPizIF2+/mZ7
xWwfZ/gP877XK9n4DzXVjDiJpLdHG1Or4UKUnTUqHNLK6DfeNoy92+ADYC9IjECY
zJqtIPSwAyiXybmUb6oPTJ5nwB8McLbNIeoT5MK1P63Poa8u0MCY/3ZJA5iY8Jd7
rK+unqWVOaFWsb9X7/0vH78kNaBMmwwCrQ2CqYoSPNvugPIxmoIlK+r4I9/yUpT3
0oXdC42ekeIaH3AUp5hfplC9/zkUMVuljwzR84EbSUB/ipRMVSe8KlMzAM2ijtuJ
eofuZKIsRUtl6k3XtXeI0i233kbNpMYvbqwe28xiL156Vc28isy8KpCXpHjFHFUs
WrVmPuYoQMjsXPCwyRgvn/H1QuzHbjoKOZva1E3nkGAQdE6wr0fvJaIir4MqJFlj
6frfWNR0HCsDoiPVSXzA6ls0CtNexcIvCKkJ0KYjnRgzcAWuasSpQYTh1zmz7zmc
KnpSCB22A5k8kpNeyI2e0Wh84QlY88s8CRTNo5MQUkCTA8vgHV8oBNqf8bq8ip5G
UwNYpUXd2uKmAoHK4/kYamTC+vKECNNk0v+V5MOr+E/J7hV9d5i56VJAzW0G4nqf
E43Ro+TyvLpC/O+ec0kPQC+B495pXAc5X0SxFU847UazgzzoPAi9+1LoomjdC30Y
EfdseU3RlsfEFX+VrwCQCg/R6hFCg7qVPJlKUurUxLbErj/NhV0pPAN5N+XgJvFm
dWv/xl3FEcWpOt8vlfxnO1fv6Ydw/FdM7WrgV+q2RgAyFK++te2C3zrM0athuWmU
wpL5ACXGtodzLU05vrPT21Mj6fimM/CH2mYwMx2P62ScwqbuPDLYbywgbcuchQ+r
v7lM7RKy1YltS4tdo6hyy5Ek5kIUdfuWSsdfqqF5iEX1USbrs7/9sR3G0cvbylyr
3aEUNpqJDFFbw4A2VrZbiBAcUsD0LPMmHlsz6fi7Nj8QxYAiGepttURjo4EGnnfo
tjWWQUmqqsW6wyjnww0ZU8KEWpLqghBDyl1t+zrpRsDbGuG0S5WEVzdsfWUozH46
LFZ/VtMsZzwUKS9LD9ndVFHu6IZH5Uh+/GyPpXC2y7F3Md8w7fVOVF+rjREAW0qx
K4ssafIwCAEqRrMvwoajJqX5ZV66JChxetv5xHur+JMg47NkbYv0mNo3fL2iOe6j
04stck9rJmL//mH/3sCWbRwkNhKdc5QfFRlqK0cBcT4cF4BVyB1jXDByuODWB8Zb
gjFNqqBYY9opa6I26o6a1EwddqZ0GunOUoWC0TqWCXgHEitlv1PNUu+C0ASRDSxz
N/7FxesmeWT3WdRSpIo5yTvRFb+CU4XASy+0ejINRmgzHxfHoeF4IQHHYJA1Ml2t
KfH+BVtOUZFe7usSNF3nayX+o4l5qWHiIPDcPO0pi0C8wbryar6X5Qe2hvQC2Qhg
s9TZi9CG0+o1Vc6eTHf/g9WEWDF71M/JKf/F/Vm9cMCP8yiFyXyUnAY859D2BvBZ
nqXmRCjtumiSZQJ29TWRu+l8LqNZCpt4Ifxmsk7dwBfdxbzep0w7s9wEOiNZ3hIn
hJfQmX6XW+eYhFUV3t864fxNNGjIKhdcGg9gen7JX806fVHDPA5cL0k5xMEHYLnY
7JU405fz2NyKiiskSjfJtbNB26i9WYN6pGOVS3EUjpj9OmYibR/2RtkZr+h8kt8f
fJqslk4SohCpoRZKAhEpxTDsPePx4USs60RtCRgKz3W6tyMWI2JIbNN+qogIEDTX
T+UaDZ++8zlBR20SCj3aT4sJSz1MScHjs8+Wvzht4HFV4/hOS2K2SgKRA7qhc2Gg
vewP7+cB4EMFyPrAEIX8hCajefDK+8mmNIYlfR0x1WF3nG5UJx4eUZUyFl+SIrJX
JwkLwsYZhypaPc53PjFRUxwg1DVQca0aNpALFG39Syue3zlPcnMqB8J8KdD4SqFI
4Nn0H+m2zoNKpShzSaEO6wiT/FPaAcwXNzhplhesZiOplMopOIUvGF+Ocp3tOyFw
XgscfdyFS5sMGlkeu0tX6+QA45z9OXsSQdeU25NKdBIR3mF51nut3SjG7xvUU2iL
AJWENJpr2huiE/vM3ai9FFawg4+L8Zo6EPl30/mkvu00mgOlElL5DBpZbC281lYW
1WMtTv1U0OzP7R6kxpIMjeVNPkKOyENahf18NXJUk6rDd6znBTNdQb+JtMFpLAya
NZLa3OB9NtIpM7+/63kYyXelkFWRK/Ot8Ea1v+ZLkubKiUg5A/zVLsbkaFlUv8D3
J8Obkq6J+sRsVQV0l+o8MrURK3QAoo1BxSmESv1G8q/L8gKw0o21NYhGoaHujZgf
65yCPmjI+6VGsoV8nndW4+C0YOA4bVwkDmk9MP7cMrO8EeyFIyrYr5O1ZaFFZYfE
SRxkd9DmUJbo+JeLNZMgdVMDCyPPB0tJflnbW5ILD6+QrWqowK2uViKvngmlhVw9
gbf9Mmx7Xgc8Rg1BkY31HOBLRmmusQ1g4RCBHl6csUdQ4s1n5OpbiJ3WYrfDFdGN
fFNZOyMlZ8TxLHjS5jiJpWT7IzJHSD5b56lRI7e7ldX/5uXaBiUNFXvC9DOkoRXO
314u9LSfKpn3pBpSAgLGfmrPJUnR4F8nCwNPSPnWJdUhkeNtdZ4q8vFIn9ObxyDH
LTjqc41p/1c3MMDJaqk8P763Cw4pQQ06WPA7JkNQH1A/TeF1iOmqgIcZTqaaZGdY
SgPmy5rmx418rXrv7krx8a0srV274lDHHn2YELTh9/ThpiQ94QzdUL/SncGhkoyf
ESd6d/o9msHxMnvyZYz8GF/ZnsGGjazT6wk6icu9B8pwWOEwGdqVlhZi/Hp1RhE+
CrUBDZQaaMmsiCqEwev7xK7uK0ucjRG+3oHzslfJtJGSr18jN9HsgW+KHdmyziUP
e4Em6jxvBd+u64yCdQj+Hh8Lvj4MZoEBpo3zK8PeOLgCqqQZRv7px7L0VZT2YYid
wdfVAAZazOX/xm/BZuWFWerf7A8sGL6UBifiGLj4iSUgxb4dsH0kpzqCcyXZTINJ
TIlcx5M9eixh9FrHvvzCzGaNy1QTCGqwqKaJCtIPCPD1uST/+K2teTi1BhBPchiF
0zUKuqPvEtLY7cpY144BLSfwMU0GhP4ZQhs0PIrwpgdZQAi5T7tU8lHbxejfW5Ec
zZb3/j2wEzaahwtib2aDOzUoMisnaUQD+tvTsFy3PEYlpUzGaoWQC3kACklRffQl
bsL6FDvOmpMmHPoRUcWbUFiJ78NROHEE84ff/YUfgPVqR1T3o49AEZJtbtqsa9ZC
FZjtFYTf6xZKscgIkte/PBm+CQspM8Ve9DdPpgT0J6F6MO+xlwO1QltJdGJDYhV2
Yx0frGZK+HodcaGv/+VqpB9CVumiDbm8ClqXfN26DSNY/pxfHJH98digYPZkymLQ
GzW2ZkSlMRPfnGSAyrGbl3JctgmSHpDOnH0p9kshyv8=
`protect END_PROTECTED
