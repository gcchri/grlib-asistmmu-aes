`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w9r3NBKP+yzNjURWcO4m4Hw8cDuCrCNLifBp8i2OYZIPMkEAVjedHjRFVbrRS9N8
xg1PKYFI/CeEkhXjmpVI9z9TJXaC1sLqfEr+vAsg0x+bUZBLM2m6wTPa4WHoUQJu
fUYnOPJs15S/KZFFSnemoWat+Zbu/aieijiJ8Je0umIE90EJLVHn5csDE9CjuWLa
X/G7Dl7lIzZ6FSIKWxVlRnrS0/SBH3gGiNrqcgzqxhdzY+U+5zPD6WjvfbpN2qX0
2IUrIbf7uc8aZ5qTzrUUAmFpPI5lTInW+Dro4zDvsZFRE6jILsVH6RZJ6aEg8Tao
TI+8wWRUIS1APd3qdstd8Al7JZhOQhpfGRJ3mymVXoF/PXpQKfxQeroNuCceQIKp
37t1n68NlCdqtPbHTFKXkSyTEuWVlMfJ4Pnixwi/mIv15X2/W1ocp+/BpPggzue3
9FFZucV17rziocldVKR4vCQVN5C0OH7sF8ulfBs0itPA0BKFbwilfZEcesn+Zewx
IBrBv9GZ2IreChyM3F6K+rTs7z74oGbcp3dXHs+XW3QgXulYp7PbuHHA7mUx4TQY
jlK+QaXdcAO17+e+V4c5SMG4bCCcOyDLOFkyjYyRqJQrHBZlAZy4vJW4+0+5VTSb
oeKgbKmv8iq1aXFRRdVqDM2rwfh/2AGO46uiKuyzJE68h6qc/MQzKANOb5/yFHzb
52rFi9CZzpD5LXjDsGX9AG++SXuNz3kmcoO7F3w0XVM=
`protect END_PROTECTED
