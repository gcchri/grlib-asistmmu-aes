`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ocY2EsAR21hCAHzSnIvq/XdWE0q8C/LE18eygU0kzG/TfYm9Qd37z0eNiXrVHkY7
fjZJujcRafsKlIhOo2xfQAguW0O3rmwn0ZVIM/YY+bjBRIPAwIfJsmyNyHnOgslp
HRhCRurNptFWVo99ipodYyo62yjXFelk9hUTwGv/sbEWd9NefmvlsdVGhaAG5GAj
BtU+wu06zTS1XjnSdX0wBQFCgJU3ZgZcLKVhrp8pw4jHd9Gm8A6EjL3XMvvAo6Xu
kZr2H/rAxGKC9J+IrdjvZ8sviEVfU3UUInF1GZMhgW7fNPg76CsP3S5YrMJtlDtr
+po0ywVOWG1xBjhmaa5RLlqJpsHzXh/NC5meVBvafdjfuFOmLYp84M1fjkRVV42w
jwnfGvfIKaLpmEHJAhSmA5FQueBCuK/vRnpVqkyyde3nAXTyIvGm6+lZ1blfZ6/M
L4kuVwAOqTHjy1rRsWgBZgf0e3wddYO9ZPwpEyerc9Iyt1LmlCrrqsH/ETYxRyx4
Mv2Y2mwrPH/ViPNNWTtOVf1Q62/Y2y3WDNvuD2yis7G2nUpI9OxOHaeDqLxDgosw
DoHEqZ4wnCoHC2jMv5qz5w2u2SdXtuLzaHVof5NtxhvFaTkiZ29hu/9Lp7AfQV5i
WmSUEOiUooZgJHyl81zzTwC91yaTfhDRLLZKJFgdDX3Wfh4EE9EfMdAytWhpDaHU
NWq7/LiR//dS9LAqbDhpIkBKFHWJmB0E4JhTv4UZzOO3mnszfZRIDOQsMfke9X1p
DeWX/kOrBeM+h5VkcxJzbg==
`protect END_PROTECTED
