`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h4moUNzNxoToqkajgU2hERQ+xzCKw5qsXPXJzoq6YmXbcPt0EwNTxws3O8UsFGTm
tkadMx+ytK4eJ4FDCFSWMsl23YiSgnl2N1SkT8PlOpbRbhhfE5RxEgls3wr4kyyr
lQEdm8LNSwVEo/TbuzDxCHspYUyrGqYllaLZry5zjKjQNriEW9GWFRxuiZf31Yrn
MGb7gOAjJDHDgs6UQz6urq0O66CMFnB86Uodsx4Pfuq6Wph3/6TDr9JYhoVNdM+n
UZbW86XTBoogQx8oQMMErckvPs+8GV2eTmDjHFeXXwCs3FFKU+uhDNWOk+emK7r+
86LrJixIwjBLFT9yf+G1cZ9MNgw5aVJRRQYDhh5UDsODYZETgTjtiQYd7gAAhFc7
Ga00833mrkaUB/zpTa7IFOMC6p5ku/2l8sGB8a2fhinLwMfy6+HBtEXc+Rmtgg8R
rRkTfOGHGlpHugAClYapp6+ZlgIPZI8HD2poGmglgO313zEnHfWP6++7/Bw6uBkI
R7oxtiTIcs9ewx672XWfs5myIvoySk+YhHK5ctptaR6vUYxDFvhVnAzfDI4dgefE
g7gelRwOAvj4ESiEyuW+eQ==
`protect END_PROTECTED
