`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o0yoh799pnOnac2K73ks8BgDJkmGKoptHGIgdp2umUVVVfMvo3D/T1z06UzigsSN
jojXgD1y+NiCeZzhnUvHaydZ9VJqm99EpJg16uYI9luNo7MVRuLw8lxGGOF/UDuU
uArU25yJl+rM46zjakboFewyP28eYgSMNs1pNsyJ0dyAW40aQr1nKgowZVqH1kt8
1mZccPDa9RK5hKu6K2kYHPqtLu/S0a676Ygb7D10KgTP1K5dbGp/T9u2BJy3iIOM
9GJTufkTM5QeZusl36fQkw==
`protect END_PROTECTED
