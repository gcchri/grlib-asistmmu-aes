`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jIXnDetm58+7D26lpNv9NCCaYC0BJ1ASk/kIGm46c0Hqg2e6F+LzU6sbmp7MF+B9
KTSt7Jaf/vc21fn2MOfzF/sDMS9jQMdvjPiUQckrGCYzeaQ4uu4ZYjtIDd1s0hvB
NoIavW5/m1YsLI9CzbfCYKllUUNw9L1/j2PXDkDIoS3qNe3cV953xAVXnEgLBgMT
ZQ5WDTod3hRpNNhYVEHKXb1HZaIqc/nPq7If9tk2URD5I01J+yk/EJR7xB/sEJJY
grv/G18fz8kjkQ3cDrW1rqgAUagJqlzgrOhQAhcoXWrHAgHdyU7W52UEX9DpHs8D
Y9tGf2zK33Pni5+dBKR5uWyV5bs3N92z8h47byWMgZo6igoVQJZtprLk8RsRnLwn
rCKAdB0B0v2yM2iUMRTqb/e+Wt/wxp0SEpJJl5qujikkU+74dTTbD/n3r7SBwv0D
Dv3dXhbuNlnHHZ8I0D7oj/9Pa2viRsiIbGDJlmyv5yvPaX41W5zAulxoovaiYHlP
Z3eEN/pX2iwewuuTryjGbVKXqFOHMHrXr6C5LRtvGpLqkJn/yeD8aj0AJqXCgZx2
S06Ny7k66fTvXoyU4nvy6Q+Y8yiRiu9cgssHjAwLJLDc8iRv1BELbPkmJp/uC77B
ylSBzZfK821cut71cfmng0M16Qn397pN0FF5FC46Kfqaj2/+typ+2XSoJPJbulf4
W0CCSO/+Da1Pr5ff/2wt/ulNBCpNZHaRWAyGqZ/DatZQWac2PX3qRcOlU59OKPUO
OX60UhMLYqR7t/8su0ODBaIrB/H1QT/k8TUZEMgspEJlMRUfTv3w1mZ0rlPDn6+c
cO0c3f2bAzn0zFVg4u5R3pne+5EVQ5Fj3mufqhXFtC0loVeXmU7V06xx7EuCfnav
D47FwBnAMD/t8WQcCzhyoCexPUVHKICwj5R71y8JeEofjwdFPaGT7H3yZyyKQslx
5UOCPA70tXCjjEa6JGy3xw==
`protect END_PROTECTED
