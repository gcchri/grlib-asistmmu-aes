`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UM3wCXIECanjJ8SDWtXKq0t7hXzTycjOX8AEH6IxlWLB2jDD7xfAADp3eD/E4Hvh
+bQzQs+htPCWc7IRyItv/Owx78zWeZJSqVUuNp+vPOQa/hYiddh2a54KiFGAcqoi
W2RP9Zn8EBHDdLzKecvKluuWVy9rAyrFvyjGWVVENJr2hgB1asYVaCEk/RlFDgNg
pBi3dQM+TRpukWb+xLIJbYpbvYa1Emi4oSyXEWl6FPT50C/T9kSF/lEsr/76ZVcc
7JAIEv4+w+CZ+0FVXVDZkeviFZNY/wqXTq7nL/HPUAHobCtEIotKwiO+zQ5Y0sLF
cqPOBi8g7yRzzM8fvTeg/cxjRLMiVz3V/VN/UrNXPktCbbx/gX1acRGga4iI3+2Y
4s5tEdwY+rL/zBsbO1v7nw==
`protect END_PROTECTED
