`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Whjf4nntkIjAXitwLE0N+p6wehDPvC5BGRo/m0h37dFlHXbuxPDrOC11ZszU+8hH
FG5AvhaBGMq+0OMtJBuPUjpRVfEEBNanfjLLcO2OdbYtyzYfV+eiewi5gUL9yzkK
4jbCYFSsKuZhCNvGT8Fp6hb5cAgU0TdkscWSQ8nbR0nwuQqndC56RyNCi1gfbzq7
smUmynFOlIQPRROeoi/VlqcN4ub1ly3ZDH+UPbbbnbgMwdFSaoddnvkugbXTigKU
4UPQm4I3qGlq/Bt+sr8Nh3fkDc3UDoNAlLTxIOo+DZsTFWdgtvByPR3Yyl6SAXwp
p1yGU720nO57oOYDjvYC1vhvO6zwnqrZso8eWPM8ojakNw1N81VITaBKFLEBEWl2
ptwsr3P5Is2YUe+n+K1s9lHyZQVPL+/XhpHf6Q7yDauxjlG9AWkgSgoEB2ZGM+y6
zafthcyQCjWCxWZmuoM3TD4RekHB6W5PetaCnqBa3WtIWVrwYR1jdR/d9ZqDvxNu
TDXG4Z5BfAnqfxV3X/8S2KyK8MrBwCvxanekRhU24yloAnzexI9P808r0tVloLwn
Zysx04wUALSb2vGHJHwygCp/KEJ2j6fIe63+gjpBRh0=
`protect END_PROTECTED
