`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0i0dGODT7Q8CLsdkdgcS2DngtgLpMuD1XZl4G0xkETk6gG0TyUmi+TmX5tuS6L8T
ZzmZloPvT+mJrwBwq4dgzpMOH3YLbfUsLH/+2B2FlVTlb+0rdSsDj+rOFOiso2IL
I5gdkGBRcRH5o/xUtsAR0nS+mxLN3iNr79KPefGLDpe3q2hUz8jaHVAeDyj498q2
dVWXysZrb5kEyaUpTNBKUZDn9XgpBGng1IduJEmz2TBkXMKlKJIknHSMVHSWl12d
iRQ+hi6U2DhNpPThFDVQnZowHAuffNhb0UmHB1ODpxtwtpTISi4kpeENPRaKEcTI
3DWv0lCVzi92qbS8rQ6BUnj6CPOQnbVtqzpQ/MJ2P+T+eZ7FjbePWtmz/9IMOMWI
E+yz0oNWU6nNyPNplp3DUK768CfX8VklOAjuED3wI0M=
`protect END_PROTECTED
