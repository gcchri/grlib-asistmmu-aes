`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7wJxijZLdRoZobbDkSqnclKA36Dk1E6a+DAmj7yiQDARltkksho6dKGgu3981X0N
r0orOoDCRFl6TZEBNltxAi+NSj1lZ/4/oMQHvy7yWXXdvFajNnW+lBlALZDUrZ7B
LNnKXQ2zVy9f9el3XmVZNx2sCvtKvulGSU/JpmrXh1NEDqkoIMnrWs4NjjTAL9Ee
zt6/Cuhp1JCwfK4MxujYZEHQgPmbDYgRK69OozsGcUsaAgvvVxj4/aUzX6bQZO67
DwsaaVNXynrgCC2thZC/k/UGv37MMnX6rQvu3Ji8OqhhOnq0jSFtmj3JByH1VgNr
b69ZQZFboJcwT2FuQIqf+T/8FxlM9AP/w48VABc7tLlMYMpecDwr+8iY1FpsEXLN
5cLLsr3pJRLdhMBFl1QQYMKCGqxVDE9bowY3FmLulpQ=
`protect END_PROTECTED
