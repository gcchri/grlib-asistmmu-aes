`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MpMLJ8/YmxKgCPwAo5+jHzNUmPHJhEJSlZdgSCRrUJ3ehL0N9xqTjmcdD+qUA0vt
LI3LYHkfPEBVN6fFAMmA0Xcat1nIITXtgNtdBFbn5Oo3vImM59RJW9zI8l3y9U5N
DkUewJzfCVwu3MM0J5MSH11yzUrTWvnoQGSKvgTLSpAzsvjFTQuL5SqSjkv2+wth
d2NU3Er17RikKHKBKhgTHqRTTqdYP9Dw38MLbqieTz/HBRYjBEKHNfXI/Q1xVsDh
wUk5wqPQlHA2NoZ/JpmUaW22E3WzFoSpDkb2LOShPOw=
`protect END_PROTECTED
