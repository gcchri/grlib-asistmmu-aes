`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+nJ74YogdzBFBpwSBZP6LnYA10x7s1Mo+mysT+fwUHjx9T8I4o6gFM0ujZtM77tL
52WN4JcTKXI3PeX0OpXCJoWg2qx9huWXKKLVhqidl066h+KPG8dFFVH+jihDRaVm
hPZuzEc8BbplfT5fHwOa1JeDm90y0x5Rip/fYpkEL8zLO0CVYGAoxVOKIxCulKKX
Wvb0+JyIDahT/B1eLzlmaSeqWD+XK5GgdiKlyBxMkFjR6QJHFCuTBMzo6xMB9+rq
T7DmH5xJOxVd8FjvcVI0YnexKvHL1smgJx0sueqFBh94ExDVFkycoyuUzdihDNR8
jU0CyhXkdtc4nnebJr0bKw==
`protect END_PROTECTED
