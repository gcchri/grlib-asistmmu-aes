`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T7SO6hTnMONft1Kx0o6kO4rK0+feANms5LoVZ0raqFDjFEd8hI0DcaGbWqwW+Y+o
0foYDBf+MrtPWVJt3lrnoYDhytyeJH2A99AtHpX6SI22zt4glZ2AvxdRQIiNWgGF
8dTcGHXVQYPmOCnxLbmfdHXR8GithPZopiSuhXo9a8Ktn9X18dzNuHYZdM42jd17
/5O0ukb5OjH1WUgDxt0N6X7bixgQSh34u8wl50vg+IJG8+6JS+Np3ZvtvE5T42FI
VRpT4Mmkt7Fc5syIziEBAOu+ozW4BbLXdiTmneAbjNSU5b7kE2kCbnGrdh5oVysq
OLAQUlgPRFBNxZEiS/z0mlIXN7BauIQASQtmaOXLAQ+9RAcPgHA18g2rlMWix5f9
hKHyqVOEZD77JExuBDFvXOKL6KNwkW7joB83F9yaUksOKePi3JCB0CGcJNqGsT3q
9Cut0eu4VsasT9pjNny3X24PocFxtk0rCemHzXdy8nlLv1x8K3DDI2nNp5Cz8Meu
TotIQcqz228AIb//JwiGM3DFFjLB7ndIjZxwEhWTmRu2s7NsN/ARQrFKXbxjfa6F
japwB+fTijmYasD5GSEQogL2wNm7DAN/Z5DUGg26ThsBd+9rgFI9OG4iuWqpQgTz
BS2rkfbLkoOB/2+CPGWKVBOVipThSRpdS/YRD2Ec+ucCwlPgGEc32n8yocfwLbY8
aSlD4ed4CJPcaV3D8Xb0nNgAWLlaDLYUEopm1W31djAhuctE5Vu01vSJFv4lRa6b
LpKusjlKO0bz/3K7yQ7iuxqBZyQxLbiRX74o3P95b/WU3QxQcQP6OD0PUUnAXHdl
lVn8E7pIQS60fof+tlMk4cc+XfhJU2N7KSguT7zp+iW4602aGs66OPge3QOf5S/0
p8FuBdUvAQtQSiwcbFQ6sSX3iGE/pNcKtpgVO64zEgzQqUqFm+N5q3Oyg2QrAPVH
sNAL78Zo7aU+mX462dp+tGKcJjjoxz9PLYsTt5sHpIskEvfaNHjensX+QEXFiTd0
j+YXo5sn9HxJ8QMp7tSnidzFk/zdWFU0E9JHlRfhimWG5TRs/IVKJYPiJY6A4P0c
T9cyQ7XjfWupbgrlPOAvbl0z6JM5SkctZtRPcx6Q5KHoJn7k7fmnlvEx/reWTEBs
BD6sV/ZzlTQu1r790TVAkCpK29GgD+hRBJsBbHi4Z8tvkC8o801Emc2ofr4TJd0e
uUwDia1VC5NRFOYupZ2p2a9Erh2Zwa3WHUNs5zXzmt7PgmDfBQ/aaGJIKIPz0vQC
eRCXmo8IApA5nqWdkv9ZAryUwlhE3ZX0hrkwkMhtT+S3Yi4cG6hjN4i2KD8AdWnz
bbF0sMYQHZIxH3OB17yZvz+tpbL+C25HnimolWjezS8qKLQ1Jp8iEWcEpZdiLZ/b
vGEHJPo8gZSNGW69x8IHhidCAcrYllnaFmLfVdLWE8Ixa5tQ80wvoac9GlOLalnT
4yp11n1DIwnX4DihdiTBHgBJJs7dwrDAZmkzzeOLXLhn9RDK92bc7tc4j6MM6ULx
IOFzGLhqrPxRt9VaZMxNBA==
`protect END_PROTECTED
