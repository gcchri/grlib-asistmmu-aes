`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wno2mkRjWMbwNf19nnT4bmhg0uVcjnAbhTwycywc7D+RDrkvIpDuXDEGqcLH4tlo
6Fei+OYGg+SVXVyxAl5YGk1TsLf241CC3NlpWrW70/zkUUXYs95aS5Z5af2NsAwI
xkiQQ8b60K7G82DzA2BuaejMXKIfYF5SVu6zPBMzpc3EIzngbApfriVq7mWxk0XI
RL6gYNqD21NKi1yh5Xlrl1cg5s5tGR0JOr2plnscp3OXf94XAej3859qqU80xQqJ
IAwOB6v99BSLGM2YIj+y+JI3lmipxajvcafXFtrymDtTufbdGiT6fvUwu3RNz1Ll
3wm4pxxfOIvFFnLNJ3rdctfX1ZbpTa76YexyOzL7FLg=
`protect END_PROTECTED
