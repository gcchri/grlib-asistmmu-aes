`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dLGW6SM4+mSdcQTg3cfgQe5MBSRCanbTg4M21fwfPqWzu9Ks4DOgyXbpZs3Hsq+9
sFmeIWwLhAShfxz3FzyWYLHdYK07YGe2WePxUzeb3M4YE3h7t0nxaSv+5BsI+xmQ
HnvcxQg8ZemuqzwUBGciHtV6EvxOqhOjiV8kYPBrt0YMVbHKOXUJlStLcbGmM+Dj
53qdjPEoc+4KR6BpJlAqxrqOB0JQfe9ISV7PJSjvIDfpV6DhFjAyDNwh2jwP+YsB
yEQenwI6qBewjQFswK7aDm1Uy9A6f0Cddr9dFRllcWZYYR2VDCzx5Iq4gK2yMk+m
zuSJq4FzJIDa65d6HsUY30B9rhqeHh3QqUGdk1oVbyedF2fF0Oq0Todiwx38AWFa
7yXVJJcNlJziMVv6CkihDDk+KKOgKmuLOa0MyEanvP5fWbDWfECXk5QuyNrgJGla
`protect END_PROTECTED
