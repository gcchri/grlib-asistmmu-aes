`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VJQ3icGKwA2/TcTR1BJ9Uez/gMbh1ZN+6VDGGsNF11/n/e16satVW5H7r/2v+6LZ
hEdvcYlGXX0weOXv4A3JoIgHqaXwXITnej23yzpvqkUhKrUmKsbVqEuGyNCuFJye
NVhHD6V6gXkUePoN9Qw0Qc8d5qax3uUZforVwkIcSV9xO8x9FMjYxPVjpyQmrxPy
jrS8H+INH5j2u6S2S02Y+1xfQvh7xd37sFVXHwwRCa+fItwwRgVVzCV7KZJGQU4K
1NczStFod9bdmGrAIqwCp+TlsvY/SfWNpwQ8VEBKmb7TE6HmexJnPhuZ8SDz3cr2
/bodwc1S9oZgh8J9VWnsxUHsEZclchjRgJchUKm/G06FIvk1kdt9jwKYYHxrdu7n
D7lD1e6XsGI9ZoFX10Dgl37xkH66F+CTdvJ7AGo+h9jq3Ci3MUcTWBa21xY8vNtg
gLSbd1OGCB3wSaK7Paqv7kzayUf5bklnPFcz2l8//UBtAli9CrlIsexxd2zbNNnl
NYS1YA5nQSxLham5tHGTt8VEwWdG++AmfkOgADhMZrZMYLtiJ46btVoa53kBhbQc
g+Zak9dOCfwnO4HjR0yGescD+eXqIDC1nQgJvn3oETKgf+cB3kg9epLAbvxtt+/6
v8VOAGreBGYAMAQiASa3dIIemYN0dnImK86gvJ+1CMb7Eo8gbzQPoG82CcA/C5t/
z/FCNVf0q/8/QUvQFaKg+87HSWVKwLabv+3pZA8wNKd3pC1+FblBIC+ZuIZTjjA6
JH02Nuj81knXYvgiBT0ZkmNR9yFK2SgNhl1Gx98+xfWsCSj9AcbnR4BSoBFfIv23
7dzAstwtTqSDGZgiqfq0Ey3oYvdScT9emmRiG3jOXayJr8+EL0dewypQexxoGbRc
AFzXaWDxzpAayCB9SZwryeEaHwppkq+gXNQJIiyZVE7UqfdoCncFKs9iEh2DQfLj
4cK6PMcGKYIAf6vmy4w5c1tW/Z1U2N8MROi6ueYIIMUKYT0hkeOHy5ZT8lmMS72V
SK3NiSOiVJZrQK70MYswDgxHB/lidZvwmqU6tP3PIGVSkZTAU9ZamALmU/3wXTr5
6L6OrtGspt7ZlrK8W5nRG+oi/s8UToj31iS9onDMKXhQXjysZiSvsl2xL+VvfSvi
uEHyDXdlFQm97ZQgg375XxXuqRuGb26NMJdSA406mTfyTeDhQFIujiCSlzhQuljo
CzVeodBbyGkR8bz9gvZVsy7e75UV/EdgOlAV3/APw6I7GUs0LBCFCYzeKIutx/5E
u9UOj+4J4V8jGZIPtDTJNKNKdfcZoiqXR3D4y2guRX+iofSNLv1QL4hhu/Vfc/B4
eAmyAxNVx41Y1mqxWaZNUXYIZpKHqfbxGABD3aG/MmwXIA8i2kfoYl4mMjz2EAdp
iHIZwPQulc4xeakvvChzqdkTMj6wmJynxRzdWVzVm55IUdxp4X9+W7ZJRZkAF6w2
NRtSnqy8/5/ReCJ6MoacdtkzluBDGsfM9btJ4Ii/zOM7DLA6HyQxzL/mOTH9pzSo
+CX0A2zYAdBmlwZtr5MkEjtiOGCQ1HA1EhpgE347jH9MRKsS0tBQHjqDfTsKD3+z
PdMv8YZ3JXZPnWIYxGW9PhPKFgk6FPTf0Gc4QHhxIK1SqmQ3S4JV31r367xJwACW
Qfc6FEV21pZ/X9RK5LhURXY1hYmd2PpXblbY6XNQ7vRcNX1BkOuOnkPcTpqVtPF/
iy8Pisy6HMwBeFWIayRjaPVvoX9bkI4ewHHGABmmFDgJXLNY9cE1DgPIBPXY1Glc
Vb1mSV4elG/vzD6gTP/9SkBGIIujuSd1AF6aActMEsfIbfMGjpaIGJYAu5Bo7A91
swuOMOYB0d+JITMlJh0mQPU4tLA742xA/TKuuM+EdGPcNFGCF6bEUbS7tsYegH1J
vK0/cOudYHt3+ggEvmk/EWixkA8WYm58Q5FX/CEzbItEnCfAPWhWF+hhAouNj4ai
lZrye4U02LzkTlS9+a2Le42q1VKEF9YmeNMLtsjoy9TxqGrdQvZj9QrcR1cQPec8
6HtUQy9dqy/Kkz9c7avtSLaX1ecmospSGMb+Nhcq6FGIeBTskJiUmWctyWJ11Ogl
j+rvntVcG9rKiDeBbbI+tR4i9CKfUFDtBB+Mq/yy0WDNBrLxbDfCRE61kI0k+eFo
gTBuA6lUWqMkQQZ4x/ogD4FnaADuXYRZ5vBVgvxJoG6LKxvGi8T+dTsCpU69+Sjk
A+7CH2DyvnawYh5xWyH4SkQVxCrW2DTznuf04Nghfp4XwjEL/Cie17Of111DnEFC
+HbApqpQp5vix4qShe1w21tDNzTh1vNEZY7y4SnJsDpRVrJAI5ZwBxBxlC7VWvTm
jMUCan0Hai5zBpe55yhkwioTFlBNP2LLmEWUQ2yuJgAySA6hIawPYxcFtuA+Dr8u
RSJCJ1BEsLc01vOHVnZuvZqAuoA+tExk7Tyk4TrW3UmFmHKPRn3/qil+DnnpKM57
38/InQ8MO8c+2SNTqIMnWKsX859V0pCP0S9Y8SBnjavQeNYDBYBnp/iKdRTw73OB
gCVcKJjUS9J2Rrf5pIxGHa+lkEii0nOy3TM82/DFBMfg0lOzMfTerdpCVRIgWBoO
98TVAmWlBZIqigTihEmfhDAld9DSsguVAPCKkLkdfluudhlZLg7/mFPNlnAPXLUV
0tetKPHb3xIC9/TEg2PdW9BL1OTDAOOfLeYTrzgEvW0k+bOYX9bw7PFcScyE66Wb
+sbANtbFOewxwEskFOqGCOp7BNJ4aPm47KPYRMrRuiplg0l3EgQFbtv2gCQIbrTm
afV8PcdJd+AJUHIhy+srt7ikQC77QmxcFHZUd3ijMi/3149xpaswLLyg956FtFf4
6lJZ6gRC40rCzisSCQAWxWRF/huAmoaDabSPpJVPBruukYW660S7VHD9VnYaLcJr
Kxdxk4OWBgeZkIj16EZJYLHxsBzD+gF3kRQAi2PbKpNCq8BSSxzltjKGRP2LETqf
SLbOznb1RQnDdyyWwjHjSVstQqjr2Yxfu6sWZBKE75H2EjoMtukXUpBwbm1rXsE4
GfuWCRQghb/mDqeEgX6bX9gQIUYlgGcCK1nk+uKnIDG6JaXx4pC5oLJzODXRTsSt
wT5PxNGnY4TjZ+c/PpKXZJZOzbVUrBfM5LKHob8o1SGfN6O94ewQmrFTW3EfW3Hc
yO2zDBg8AE3aYkXK5dOu2N6JVI8hZV5dk5V+wSRI26yuMggTAT1XpEOYbDBESR4m
Cf0ilRYplLVK5H7ezZKEBGDqdbrOEVqDsfFUCU9DYDf5F7mzl8DlbJsQ8UR7bZTu
8sjxgP8wEdjCwSPnbsXYTqVf8GECb1ipIh+ssX1O8HvrWckaFtK4uHb26mLnP042
TUjs6HaUW7nENMJxtKuFPdLJ+ho/TRhuIUeqzsdXomS0Q6NZpx9IwSZbkQbcuqc4
u+9ExxF5gMxLupXD8eRcPWXPYfQpBE6ZJSXGsTRwzbnZa3lDE5QcsFRmX/wQnJDd
6FbJ0y/8DwjGNxM0h4W+PRpdmLz5PDwz9Wklo8Kv1QvXH4jHN7OZnCwQhyeXAGct
G+y2+VUUOZj8rudmBCNrsZtvCR9dKo8hUw7mnGeJq8loCU97rrYQ3rVy/cK1gK7n
5BJ3/f8qTXqEy6Uxj7MyFuhqUTcDusflLHixhSOS1qya7mfXg709e+yJcOk9qPt4
Fhin+zPK1v7MBWSbsJAacWdQfCB3LQFr+1HqY3JR9LZMYwt/+ucuiEwgogshcdqq
j2TCqGUlmVqHPBqBILbOb7MEAy+x//lY6BeWoIslc4JL4SL4D+eUFNTvb2BIv4qK
tZPhdaK76QXvRHgJJhrBwXMCiOS3xIAosQLuugAMhXiXS2gOaRGpQVgtg5s1WROp
g8CyRA6hA9yHYeJBV/Ktkz3fFJtFC/h0NPPFbc0jcStkdqFFKMXuf/iRCSyOlC/O
5IWZcmKvxJ00JbtrNv4lRafrAm0TG55nlYe37QAUSMmRhU2y7gylGaiuBhTpcRJk
bYkcEiHZ8CxMV9sSGAnFOGsuDkEEG7KTvwRtV/9NmjLKZ5L4PBO9FjqUPfkuPSIk
vvTBYXnVn5c7ex1F/18rEauHuBQC5CQtI7WbFs960srnqJSs45eInxKVd1z9rGZW
PDV0Ue+pRbHmNcjnFH+u8Wl6yrtuXC65t6RNEBT/NGFzBQMuW4BfJlr+JpFFsMaX
FCFHNXb+qTB3SbR6Bm5FmA/MQ8T6DjAeKCg1+w40X6ZqKm7HJSml0uEGIq//sezZ
d08l+BX3DLuhm6JV6/B9/BlA0BLXYYhDRK1oGaokSISukYX2AoFWAu56OgQweBF7
4VGYjUdM/atNWBdA6cwlleZgRdxHe3Vw0/D0B34pAQ3yAZCnFw6BUUdRd+QWbHdL
jgAnUdN/dk2Yk7jMkf2s0NqFzUdhBrnzOBsq6eHhLSTBrGaX7E7mCyZg1O4/Seel
+fIvtJ77fd0ur2+FapOwUNVdV51s6i9Dm+cJhS6zDZf+m+7+qTQ3IpOcZt7Bjxfm
mNl0uX9ihmvItFVI5WPVLp2Nw9S4uxf1tK7LMuHVNhAKnz7lIDKNyWVZqf7D47iN
AzrdfhT+gLFL45R1yRUDg/ZuZJV8ZQGFFWYUvOyGe+UVPQ9DZhBVBNiWqIvN9aHs
RWlhHNbGEUgBeS/Z2ok8XyYp4TPKiOVqkWGoepnl3pEuhLm9wgnriuemnxTSMTiM
MVyQCKAydQoCL/gNDaaOLSMcztNxzQ7AagNyfPT6rOqISsPzPHijMgVxVAmMN2Q3
iQzqTjyE1UN41v8zRHgpa122XOUWTHrmXzJaGDHqy8Z14NjFm3kTrZWM2GhL6Fdp
4cZxbFdX8sMwutASfe4WVsa+5YgMbggwJIPl0vsnxBD2k7hpo3LAhW+6/8Ujr6O7
WeDlX2K+oN6PAXOUjnyUzCUwfefUslAeq1wDxqGZuVUpMSXOJ8yVzy5iQNjU5Qd9
9+a2mSXGmOJcmkKYV0CAjbsQ9AiLLq0OL0pbm9k9ZhhJkboD0OrSucKxP5plHha3
L8itWRXxwvm6daBaKi+7z30NDvK7fPGN0v9AuNnAlB3bnMnSq3kFfVxbWd3GXCT5
VweTDA1K4lHqYztRH/UQ+UOXwozjHYnWLqnHBsmmI4WH/JGa7QB+CfmFoLN/aJj2
NnS5sWsVNYTJ4yeMFm7mUdLClHWiGCxiKyvLK+7FkmE6UjpFRoJecZdwILH9H4hk
td0NPYMpvNBgEa9KLT5X3ttObXcIP61s5xnDRWrUfOplvCFDWikYZWpGbCJFqGGx
ZiGkJ3CTVM9ypotyZhow8puJiRuSptkQqNVlyM85BYN7bgh5hCS/JHjK9bRVIp4z
a8w2brOpohjyPcqgVX6Z+gbsmwFTwKRXa3/pFWQ3D5fQKawXlH44wN4wSJpqfQ6/
ktTVqr7eAS9PEFjiV++BT93oHN45k0JaTJm0UAk3vP7r6dTBtjbKhr9q3wIAAA9K
hmm/kFPTp/2hXr87MeJawLIKt2TbRsIW4ERw/ogbbSdXEw5mcF40SCA7oLdv7sdI
XTCKmf2ms9j4tUEl3S9I6k0GAbuV+ie7BYxEcBccVssT3Yr9q/gnZUAg0RHgKYBY
d3x8xQVF40IwzIEvEdHi/8QZwfBZQrr0awL1rQyOVHUxKsWETHneqWNvsSyx++Ie
OQKPKIQjvJ65MuyMGFAe9kgbZHLTYcZ6E2HHZ9wHF3k4LKqkome5KHoxJJ2DWQcw
rT3rv/aSe9BctyXsD0rciyfkwizYCIdIRjUR3G1cX3wkT1j0/4c3Xly0EfbZ/hmG
YiEaF19ywvMzPaY/sbiiCFHs8U7H0A+CF24jt/cGBIp3xF8cTvncu5R2iajvPUkP
/XaJdT7uPF9JHKJrQjOORa3TqsRiMfsrYVg7rutlRcOzpPj9dPJWGbS4yghd5Znu
FayjY2uV3zl7Vy3fAAabmjbVh1E8H2Q6vN+PptbnoXTzTwqMhmw2Lh4li2wlJAY/
BzjG6dme6PKYgj+H3O8iZXxLR6md+sgSEYrea7VKDXok3fWjshN5jTCr6zV0HSQk
X7n+Gf0+E2PMpbjtBGfN/RkcOMGxuwGLpc076Gcj8eA9JEbO3srqJwuQBx9Nnz3/
4Td9IOX+N0TUx5MadhnaIJza3nqsS5ekNHg47DYTTZXLWL15t2xCswCJZGsAppl3
BavzgvxCZE+EeZ1OmTex+JmQH3aHSXSF+tVld42chRePPi5z79pIxThbYMxmWhOK
QlUAmb+PblAIHH4gonHdrIF7ldTSGSgcHU9FemvkY9ch3hGb+rLy8K1KuN/trJ2J
eDRhcQ9ShqNURyZt+v67Rvu57vbWz+aZJRXZ4pE5uZtllx5gH/EFq0+51sPH69jb
wC+i4S+H9EG+BBc3uoD4AeBUID0Xtxc1j1vRVSWi6s0p44x0O/uJIzow62qXYLxl
+nORU/sNhLnfrfyefC4SUXXx4MxVwPC3iqTARWvg9WWJzO1Gvk5GyeB8fNveC70c
6gT1YbmcHnY0npR1LwMS7+L1IIL6h5Pao9Sq7dOUUJTQkt16V8f2UPKbKN3im3sh
GgN0PDnlSgn6Uovrixk+tZdROnfa+dWYh6ZqNdT8AOdLT3nrY2kMQJzzSOcyjSaQ
hQCVgX24yGDK3npQkZS57PSuO2yAzU7uxJT2ssXdf6mENNpDX5MG7D/A9glXPpZk
ZKEwpyHmpnodl5IFG2SEGCPZmVv2U2heoypgbUSaF3uN1Zto55Oh5DlZXJzWa0/G
LuIHqxaooQWlZ3iQgUjDtcKJBupHGL3N7VFLsltcnrsqeP2M99gQz7FtvXF7pAvX
yIU3dX0DBysyeljd4HGTjMaF9GlJ6f6s1xjcDfn1wb4p+I7RalSFobbPZMRTp7X8
sjywQ6O5i9aRmiM/e2eC+NQKHu+EM14Id4e9iOqcgRKPmmBP/4xQyjqyxDv8LMGC
2G09W4qMcYKJs7BbMteLnYQ9dDKB2U+MynyxyncC3BRvVuP9SI+Faen94tsJnUgV
KHk+aauz/aKrdNxKNbqCfTKxcwC6bsujQ1TCweUorUfX8eNASxlhFhyVWdL4am3j
N03+E9Cu17IrmWZVU6hbvfQnYv2eaayqU/s6b7PvbjVNXKe00u/tYyeyE7bWTvIj
gzvnrj/ASLPskJ4bkzOmEX0jU/zm0CM4BAl4ZrqsAC1y+g8aYk28Y9xRDKa4/0kT
ziawz0VDH63ItlqMqsb/Gpx9BwG8Bc7ElThVeukQr8GOnxN79Azs08ZRTnq5ziNV
a8MQDJNkXtg+/MDIexHW2oZvAo6Ja9QTdQPqaQCxFcMwJqMenieDyAgRlve5KBlh
aOIJoFJ785G8Zog9KOl3y6tAyWmP6zlo9Usi/8UVaOqgQvtpdxLVSDuEh3C3bMN+
PH4Ahp/DarfbHicZf980Aer1I4VAm7mv/yJxBPp2XSWd5UiataOWfmDnv2OKL9In
tq1q9+FMgRVD9zMS4s+KB7fb//EHUcz+t/SUeawZ/ZwhLhMlu2m/SxapiW3jcLsm
CRHPg0UClT9rtB6EDANrJCSjp4GEG56JMTklifnlmesrF6LMcCwProcmtgTK4fv8
HnYxz7S+rXt3Hp5dv3wlMnTQ73SYkRrtkxuTkWeLfi8ajwBVGeRcU6VFtqYN0FsS
oCTy8DzOx0OTCdkexEY8VU8DxOdBfM0B1GCe2EMNNilnpVAlXH6WWvrDK8UfLItj
/nQ/6kcC1Wtu1ZcKhsSI+azzPLv3PYSSbAcao7fEGGXhJ5fHjZl/TtNWdj1b46go
RyqxOBdRXNyPU+5R17BTe1ZFgcW/8tLcmYC3W33b6Kbxotg59Iv4VLTFrrIMVnK0
Kc/bj2hr+R6s5voxfhBmUFTPtypmXZalXhQCOfbEDSw2ilCa9I6cCZzfrxdGL83P
PIPjzNHPZWWnqFYTaWAjCS2oFFqHMC3LEK39WunLGwk8OPlB0hZRoFaIbSxumJ2w
6Cyf2yCd+SxMQ5G245AAZ1nLWuf4phqHj1SBPDBzs6gWbrKcTVutBZkpyNYLt5Ed
Jz6Oh263i87QRulgPenOYXGZE01N+svwJN+HAHvMO1aOy7ZEvClOxdYD7OfVuIpH
5OoYfpnOmO1iPUqk6MxQ8zW8jb0CjWw/V0cmxTjfwHC8tSK4b0oVi6R9JP1XZYDk
gL8NbkBIElseLRWUlkpq+vU5nDZRYUn5VNdR1fF+pcobXL+IJzVLIBNpgFm490tt
oGzBTjGWzrcX2tkuzxkN0+A1yfqKiOXMPwUEgVjIJ71XafX+P/Bvdcd/WWvbH3Lu
Ps1uqF8A8D8QnBCV8o7ynGVheSypt1bIXApPqGnnZzGT2ebYjf9+br1DmlMaptU0
6U9FHPEonLofj5EdfcvkOAyxi13WMLle9jTf1cutFooZQlf3z3cWwZqdITofEfqj
uPEjWplcJaEYbrcTZ2jT2E5ciIkk5Ffuet39rdh1YMCozpQmdqKELeNs2s6FLOI6
bvlY8GHXCRNEoNWWObAES0bMWMFcVZN7kiahh9L1uMBlWot+5bD0bVEJSD+vLFoj
7haP3onz7rpbtoFYazMoYzJAvqGazPR2AiZItvjSg4wNTKXsAZe/cSZefzmorJ4P
DnzJPKF/Yp6gho5spqZrN9u12kF7C0JDRrMIR11YzpkbOaI9Ucvt8NiO2tCFCcJV
LCTn359O/bLF37i3Q6EuFNY0/5/+bwa0oZAcrEhs7UDG6XZvNEQVl2UnvOEHiIHS
oAxFdyCNZyIbFdC9X5Ol8+U9PaK+sfcKoQwXwsAHt2ayE1FKDuFAthAeqtHcyrq4
QcV2fQLhhHMGFGad2nx/njycUfD1uXIRsNQ0Ec5VGbIO9tNNRSN5/4Okq1q5IhxF
54NN0OU/2+GFjURxsNmhdPvFMizLxnNxOM05jRTAPG/Sj2T/b1F7voFS8Rqhz5a4
VO7ax472vYJabQkyUhaRgsDBtiyE9ha2WwnmrZpbvNw/WoqX51SF/NsYU5JAn6eK
lUYOFVYnYqwx1lkEEYgPqZDWdJ2iXNE5Qm4tsLByhT0n8H0Z9LVmhkdYi5o9uQTh
UMEWb4RsDkZQKXoOhJVh5zPyEZabcYpamGD8TPo+LHzaAnWyfK3mnERS6vj70sdL
zrgCF7yqfeCQZ+0+3qXCHBYAZ4Ep3n93iPmnKVgeslK0YgkWtD2RCngdpZoE8bL2
ME8QHQAM7H5LGXmL+HB/w1xOyJygqazFu0buJswbAPrKhAAnfUzT48COnGVsbuff
taUSFvrMAjgb7PvK5ksix1oPOOO8j4u4pB5woXd6oRWG+CI45IwK/WPDmRofaaK0
aZNEPSG3v3qYUkm+TEOHvbdPPXgAft/oLGflZPglNNQOoeSNa7W3+81zhaOTFTFb
GvoBtJS79djgV1iI5awlhbmpIe4Q8vPCmaye5/cXfWH7Ha7Pisy/heBFigB2r0va
hjWWXfKMQX0flBQCFFZ0dPhGK2+N3geSR8DrrsdWomOQ8Uto1vUlsZ1ya/yaPQFX
s+4dgetKCGPZ5ExCoXbhaZvL2yCBv/FnjoOw32pMn309bVE92QGoiUl4v7NPF2Vr
wk2GjsBDc/6BAODzcNWA0IfC6B1/p9W0fEBvdyR42OF65MazLQSkWuUHdtnd349/
YEUz2uoeqIx86+SZE4+mWQoDjNpDoVLepMeoqS8GqqIqdKNWOh63QUknXTkvbmf4
OkF8Th6Rd52inWoish9L32smpBh0f3EFj8DY4NcoAaTvg5hZCjqP11xbaTfSrATU
WOdREnJ/4a1Yynqyq9krTMVANqPqCZlxL3a1nJlna2pk3Xf4s3+Z9YL6ldK5G0gB
7v8fs6SsdE58sAJNiJSEAUp4kAqgQDoSVDFd+KI3D755eGH6M8eRh/p/G6yQvPdV
9QPcfPoKD0R1tTuKC/pAUuYy2B9kIUKUqFZcxyuAo2fDrCHqg8f+dpBLZvWFYSso
/WTxaVqGw1qnm3asLdvQxbnogbbQtxgfDVcsdkukI+FNpj/SXv4N5hLGgdw2JSQZ
z6EbQNyAra3xJChN7a5mVNovYXqgSRcvYSZ4gJVYeNhnsFT7hIQTh39S0RAmgfex
b7kTkPneDXOGd87plVf+zqhnc1L/20+deTE5hUjFFlawijC3oTjqE014BWD7QRex
VEplpPtzN9lFJscTzMQRFttyD1AnBlExuCtPrEvhd7pB+bIBxH1/Vh6ZwCOTKde9
tqol8GpEA6BfQagn2tHLOZ8C0/6e4ODlPnSyQyCQLBa54fSkioxT3gZrjZ90Pep1
qKqhIvm4B50anurjLksPt02N6ffnDUbMexcV/cOoZOLazswtGK8KMEMnnxM+hmHm
Pj/9VMN6DUPv4LEj6oClKNXMkWaKoD6l2byk3Uw2M5/GbwTC8r81fd7/CiqYLt60
W2SRMiFDVbdpl8deAukdSqi23JvOvHkH9QG2VupnRoKhclsTkiA2dIwarOp3lK3i
91SOTAZJKkQQ7S+uoZI3RudlBWgRXlx+2874YlF6GZ14hORBPks3/5A3EsTwCFwG
2PL1/KrTO1xhAIAoVKxffB8GQp5BXwrF0wkajV0IJpIlt+JAgMqUblAunv2QRzbs
zzRrss6nYilGiZyBYDQfnrPA8cWr4bXCwJ05qIahEDOxWsG9BqL+p30mxX2LJOKl
dD0uzW2osVDkUc+OJ56K0TGvknHZvi1vUm6XlpZMUs0CyUueLWS5oqtspbcryYyx
5S/+Rxaz06JDqkw/ubJwc2ane3XjaPsbZIZ1HmkCzVG3zlfAxOTo8GVXkH+m78CP
c92p2/4ghPq8RZF50LVhO0+v1EDIy76GhjD+Gwrceap0Nmd7yLqU2zI+ng0iyapV
E2wAPNZwhHC2MdPVyAiOcWXsKQRxwGNk57l3223ouxAaCVUL6ymiB3Hw4S3mbA4O
MideX/1nGL0jRf8g7tPc0P+GMw3WKyciJe8uTu31gLJpJMTqnch0KeegDR/b5IFm
GNeSuJHy/jpNruIwn5alkf+Vu6iXH0Duuf03TvF6Cj/ImZRxPEkErN7Ukm+HGxdB
0GIaWnw5fWuXJlO3dp+7lVqwruk+7dx1DF79xqvE7EZlxHKBxoE5+pqS1BsXYsaI
C1fDWsdJiSECHEiTTwKtiL++NV03n/z24sYwkhg8g71IZVi5f8F1VqP8uou1rXm9
B2qW17yIjq9oX57bkVVyQNKnDN0FYfA1Ju4M3pJ27ryBS5yyWtATMyCv1Y5Ypc5i
NOW3nfRVNrJvjGD4L5GYo2WVtKl+A3T+EuurhjP9dQXhCteTAPReV3iiraXlieoL
8OugLSM+FJHMfH44XSYS4yhYAiwCY+G7yr3DLvWt9lAE81r49RIwuzpZN0CU24Ma
qnN3mAYpPIRtS70b0Ww/3e1vF+sXTZALyBuu5nRu0arS+ZSxoIyGJ8ZCIwnhqLXf
ncgVisAyyJd5AvIsHIAlTthZ+L0kmXn3CvLK9nsmEgiUUDwtyJS80wp3Q7JKwMfQ
315bfLhOUy+s+ajcdCohIdUXV3jtKBxHRbXKiBv6SdLoIidTfV2a++zmaNHh95qP
/DmUZfab8i95XHZNum+XE3jBw4FxoNfG5C3m0S0SPHVULx/YHKqAdjj/x618+QzL
5LlcCBe50/lEmZHngZKBCgo0KvQ2C43IPV1dQMv+7rpke6utMQMx4Aso4qTm/5lH
V937R/7eUTNJDkGCw4N83Kg38UYVta01NRGX15c3LIHD+VpQeLYdDOEuzgyS20NT
whsjRshFDZMjIT9opCKBwLbI+p09mnJksqIbpM1Ell0sJfr9OXCFEH3A1032XjA4
LwO69bv9vZYWJ5TFCFRUh4yC1h0WbTK+QZcAULfM2zNJJW1B9nyCNE8AqegTYrv3
E+6/yAZO6w665zfyS9y+mrKtrtDhvUziaofqwnZofGDVBnYZPzd4n+wx/Tig3x0/
d9Q9dIPqxybp7FvNjhBl97tSVzKdZT4e02VI1QE2GscGAXvUi7qlb6H7WAg5DQIL
ivcNK/36UGYPThpwFhBic41yv1bCzgx+VRwvJm2wE1rWsgvSF6yTpVTz1cdD8M9y
Mq/2N1PpwdF5bV4BFoFq5HzD4F0p5rDNZvtchK6nMWKZcSeKbcfA2IounDuxTWyu
qc0AQ6ZciHdut+o6GUFTfJlaxQdPvbw0wvROAsKVsn//iGl+IKafopWfd4keLoHl
Jt4QoR1+K9y64UVLeDzV1vD35woNd6XdSs7J8FR9FF69Rjz9BcLL0mBvaLBG3vBL
NG3Q7j/6KpeZx3zmODG0IC+/AOhGnx1mXclcVAjOvX3e3NI17+6xODvfPPKDbucr
8MbCFfHkZnG4QLr8ln4HfkUAfL8dT3LwUstpTI7Z6rJW7j15t1HLstbcr8VNZgxB
ZyWlQloqqggxjwEkc5W1+RsGgd5l87i5C99cC0smUEbyGCEkvp0pyYWbOyPLrC9g
73WCkTBgUZtrOksFofoxEj9nAQih4wC7YXELRDrtTUUSN7fNpQpV3BCqs0zizOVz
mfokqmnfpE76CvXyS6aX25ui8T38rEYCLS5FOIVJKjmxHj+FOY5PPt9EcE1nPpjW
wd0cxHhJc7yWWqUWfSu8UC0tB8yRh2YammRVj52ocVIhdXadsGvj6P7fkfAPfua5
SnW04IowlV3TNZa4tqW442oKFD1wmXegkA6KJwrlzvyIkS8wOq/qrk/V41Yswmfm
jjPukYvjEsbzrClwIXV6q4qPkPUY3/GuHf6E0RKh0ZgnK4YzTRbbTOQuryb1gBPu
zgN5DexBhn7Bv5FMm9d5AVcxUAP0nJ9hVOTTuQKeEWi2BZIrSh4/ETjK27/WvwJz
pHqVpaOU0qKIwKkr6qNWwNlMVKZDBVfm3f6m808ssG2G2rsJenYZZQJl5LF1YY3G
38RaWUzCwKPm9ICbITyuvl2s/kqMbTWPfX+U0FBMUqBvXZNdf3wxeoGQmcPCdDSc
8zrMu0Sb3ZqfMoLPQESCquOqcX5WqmSuzv5kqZLEAIqzuXElBJXxGt+VBtaJThkj
U9QdcyrWCIGSjK77nlrlc1sP0TNuoo2k00bd86hOhrxvVrqgm3LOP1ZOfqX15G2K
0Z+rszmtANHz7/M8wMk8cCohJmXG6akA4RFU2NMTYJxMfL2v9aT5QVtKjMBFVkJs
JuX3IGrIn4JJLJ9UxfUCLf075JJM8ECvxb5DQRFzF3CpZXFvWQLPQoG9PIEy3Y6I
gE92L691syLgHhzPyJYVwn3YDOGgCVZ5qDBdHo77QrBHwYeCL/RX9ZO10ZwfUqbD
7d0QGmEhkmAuUqk00yR0fbvKtSQySnV9wSD08Di/icUe4YnsB1s+Szv8Bqurb3WI
wCrJLcXIMy5Qf982/yIU3KlmM56Y/5J8EbZy7H4Ldku2R0I4dWWZG+ItR/pNrTWr
wwtSonCdfcn14KBmc4yTosPl1u8eki9qkA24lhUIBEVjM6cNOV0y30BlyvT+CtYH
egUE/oxDqvieDtb9M7SBpI47UPWruzOsZrBv2KiurcdsWQ+TDBfg3iim8uxg+F7u
dyQpPHKKDcS6zEqTBPeo45IMsEYrR3Obeqwdv40zf3cA/PkXhQ7f7oAbWASkmSoK
+BphwfqD83p8LzNV8HuYTew93xFiW9ZGZeS6ysZsw8vLUqSHKuWelkMMWRRyLAwd
Gsq7gvy8kcB9vGtFrJ99ZCMfHt3kQ08j2VRiILdpVww3LTXWrOPkNAeacBH0U3uj
Bh0v5yjXgoEqfO0lzDb4ruuUh/R/fzjBaLAZi6z1pS+we8OEIyE7F3kP7BNGx+53
mpjJazjm9jmIwgfw3kMtLxX4ONhHF9RSaWtj5keV3FesbllWcWT85c7TdopC63Xm
26z6JYX/tlfQg8DFZyNJbAmb7O2jQoZrRLcyc7aneUMP87do6iLmpu3PvDixEVcN
1G7sx92uV/3N2BypElxYsNN1jXrJVI1Zaak059dpOlnqKnFQZo8X5R6h0HtGMbsn
Jxql23boF6DfQkpy/zeq+0uGD1FUoYY11/Tc3wo3bxRSTO3w4dsbIQq7Oy46jaYS
hOXv/6lwDMqzM4wOUGqVXIU08y0jhR0umNKqVqbrB8Q5q+LNWmYv7xzPmHnmb6ME
FVAfg60+5RW2q74uqizztwjH6wzja8XjNVn+Hnp1dtdhqpUdUwzBb1U1E6D0uJoX
Ynv09/ojvtq0BaFjPXKHU41Dd/K4rLoJTS38s19CppkYazNP+Rrw5qKnjulFVi+m
s5uqXWiGK0zxcsYa5k8vQ8fvDvSt7OElHqPevEVPp9fzn7L3o87qa3XHN1aK9sHQ
c9pEY3YFy7BdsSMINcjUwa5aXCX7szVJPX8eFxYgclRAodgZNMMoVUBBfW2RdLsy
phbWZ0uGThKNjQPLUf5+iGkaE18pwQj0tUHmwdVsa86Fbynp/2Re+Xi/my9rN2uX
3b3q/r4mVmo8a30gA0xtIf5vF0Oi1AxOodXZBQvwegr43n3A1FHHvtFJZbnclcbk
QZ2CxgA6N/OLlnJOpkfoVgRO1nRCZoA/VukaJYprAmb9AZr70LVxbSxwk24aerVX
F7QRYtnBCAdzoj65QP4KbSGfmK4IvU+uH4j7NrMVEopQVaO87OuE3f4DGytrDvpU
59pmCPUXLyE1M2INmPQwg6lzlPAMWLdxAXFYVlnvAMWNk9oKOllvGBhjOgqHP08C
GDz7QEyFzlZkoQtDEXB+6g/ktZpDpBqStpS7AJeWzcPyX81otpoKE29M9UMZ9pQY
iJvy1Xy9mkwbH4JMMyE3g9700eHjipqkYu3Yd4udyjccj0kdCHTe1K3WbSwnYFTU
YSPS01PFvqgFPoheJ+U+zgBc4LMk3ZDGCP+kHS9nKTsjEoXdcUQqgDDM3Zur9/oh
tdBtopzhHPy//rreZcrj/zF7i5vUDaxsUQwRU6qiATAXqEkZXum0RGL9vRmPcz9u
+j0L3LNwlbaoYF8u8gqLj6sf+I4enzbevh0vTQS5JsFcVbh1JUuprmy+JaZMUti6
C2nMVcgMcv18Dyi1Rva8jbap3Y/KS0izg8AfkLpy+rlu13ZB1Iog0il+UMtATd+F
zL3+iPo6UOzNffXvv2A2nu0QJEU37IaRfMr9ylKUJP3iMlE2ckdVCL33Tkrzz6/S
VgqEVXOIwpjo1Oh7ZVP0uYqQmmp2MrxUZoLdNwIKsGdDmv+jSvNA9XBLoArwt5b0
R2ZUO75rlzDXdt3rJM/1W/lNrNaE4CWBkiNqOVNcH7eKgVWxqMmsZH0EXvEX/okc
1cvpsqIxwFgDkYKAGdxcsaW3iolg5ufVCxTluT7+DatXwjQGQORiDasar/k6t3Vz
yiNEOJIDwxudzQyUHwsiu/GSfhPcAn8IkIYNz2on9aIphGhboN9ycsdKxcWXg4y4
J01WnILqCP1vyll9B9mmNShUlAmlI8JP8qE4TpH5PbQdAF/RWqUBXzQa8c2P3ybu
/HNBzlgQNthMQ+gzT5oko1hSRZ2D68b/K5SQHayFkafgmktMKB9VHgJxawX7F7gF
HuXxOBuCNlkENeSGP9w74pw4BdeZQqWwFEdk6WSx9WIgf/0+2s1wnkOdjBQvOrDI
Pe4A67ryvFNL+LLbqt0tK5wb4cTmEaCCwrUQqHjX6ytqem9J4l2eSXIh/Z1Q9byK
u/A8qAd9luUaeTGxl2pZTyDrLyJWJR46/GxkWOmYrI3L0kMYuM6cjKz7vhLa9WeS
fBfcGkH7S8KCVJWNsS7IvPpqv9zOGTqHpDeII5rspxcn50Qu5yoXkjpfF7XSDpnC
ZCt96mPnJybcLPqg6eEdXdGXFVDAkD1eC7zbG8mz4PWFBQeIuKmuCC0TsGzBGjKE
ccM7y2wAnVF/5E/PQB4g9b7SauJ/kuWIC5D1Cr3VORs6UdFjUoW31s7ooAjomCWY
w642uKPAzUFThz5ber+TkS9yIw+ZKgZZ46UEakp7wb22yRXXHyy05dq8Xn2qfmpK
7d1V6MRFdxh4cfxsfRx+5T06IUYzEbD3o1PKOatHJRvBvjEJOYTa+ctCJ/vzlj1+
Y1QL1yCYrHCJ2mEbwQBP0/6yzZXtu3iYDv6S0B+0zazlAmBLKnqMfN5WfwL0iPKe
864oaSc/0uNXvnEocU9Kdjg+nx80Qi03dRbreuq5k2je+MhpzWUoqeuW7r8NKC15
PT7/8Qvt42wTQEFJgEeqSw91KeiFQQXkVttR7KeeAxx58IcezrzlAnDHHa9jEwzO
JZEzDMUYEdF08pbGTTBY2PffXjwoD6m9R3RTX4Cg8On1t6MD+zUaRd07htq7Wnif
QlXzmJ8hPkxK7GGahityP71SbQHbhaUr4BGKoNgDoIOitIfNumTOZovHGpztXcK3
4STAO29Pl+4dWGue/NnaYMXfPvCl9gr0hK151eMVciN34g4XzSU6o3gyPJIjdFGV
arIxg/+CbiOSnEbi1sd1MntPaAW0FLrqeoj7bb8WrYDTGqr+RsAcLbZULN0uI1S4
Gud9Ii+T9+fgMSzODHXqnOur7i7rBoxukJPykkcGdiDZ7QoKrLPl6dsD4qfT2v4W
ndpPMtOE02L1XZXqbtD3hsj3fmzszRZ7mc+bIqrl9tovZQPV95JrULvKW6yy7cvR
VTPup0sNOJwpPY4GKzbQtFcO5qS529xsOlBVy3NR+h6jDlEo3D8nVdE0LcxSGPgH
vwOGsTKE7u5t9vhLECYLBi/4J8zkIHccIiPP//8msoHJi/IcflgfoyYFSoaoFUED
fdQpa8xXgL6wTrnOAyQ14bcfhdUX5xEwmHUun0a+HFdfXrk1R/+kKkPfa2RqQCm8
/yT/Swyzn5J4IK2iEQTNTkSzNS6ZpPPUFaTYg+E7xrvulspYHjRG6TtRQ5Er2vSR
Q29rS/HJHT0JW5cDRn0gTSQrsZDVFJTVX352uSqfuAjcdR5uF74csdX5zAdeaHDS
Tin3P3bCVjY6+jk9KLa/F+ctSa0GQHqjOlaEzkaEGvXCKlzkdeXadBg0IdQA/r7R
s1w00ckeFLeMkX4wKC4KFjLoEASjvKoKN63H7gWJnk1d6RaTP4AjGVdbB8qFNCkj
vqD9Q1V/Lg5gocF/eX8J0bSaSDvX/9DOYj5PNN65ST+RmMQ9HHR3ChSQEI81CSYY
EfzyQ/AZ5WSlWipqqMVX39Y2QkVZCH9cBKK4Ec8geshiT2QawoYGLA7WL+e3Xrcz
OnThlvRPe04yevkHwogfN3qqo++1+By3ZOarCA4SNmNYBSJqLrOOudF1kCL0WAV2
hr7bexbuf8db1LEYetc/mGCyCK64bNEPJzwB7pWR7xTTnSAhP8r1FGLMLcemJCy+
iEzwPRsANcgpsIOmOaAYY3uaqbeywQTGu43Yj3Jd7i75t8pZ8m+xYBptvItVd26A
UOaZ1OeLjNjvZCbFvqnAuPvJyUkKUYiWZ4h4kA/lsT+5tn8c2UGWXFF7DYMTMfza
uZnVwPY8WvpT10e4nwzJZtmob3tFYK4SXZyButcM2WsB5NtZglNSKTybkXjnyguY
ugY1Eojs6+Or4V09tZa4frkp7y+J3Xe0RC8wbGl4kjmujdulG3kLiFHIA/jUG4+S
wnyyhUbRDGM7kGT3Oz8wf5/H6HKvQh5Cnii0UtzAO0W1Xdhv8gD+mou175tk8S98
q0bE6goPhWtVYrSrlVOXHQweiOtPEhWDF7T6cNhBmk/VKxkIr+nPJDA5Emxxby0e
I5IY5plFRsk2Uqcp+xc507FpTBgC8LOyJyjW6PsvhoUoxZLWXFfC1dzOgRLvlx0I
FU6W5Su+csz6DcBj9cO1C3h5+oYD5L2OKxnLj4q4N76p5t3mlhE51R/9EFm41OUX
/dsozEdx6xDuT1sdRny6H5cqyfJfyfByaDBykgLvU95POstWWYB25SEnvMdNaIk4
hWig5SsxZSjTQ+K76otiUF7rhaGR/ASrk7x2aCRE1ylZhtdTC0d6v8E1ohVTXZms
W7JSO48GnTOV68kLlOxUpiHzs12Dfhau6MJNHJxHtlQoBmcPfMcWFh+C5qm3Vxq9
Jmr2Uo80RhIooKRGXkHFVc+zI2VcM46Bek+YAjUSoqbbFPK/6hGIzE3n+mtzewhE
JYkmqwLIQxZV7rUeQfQZbK0Y4BSVbIhhWvYn4yqmiXpnmqvgaT6+AH//4dqQ3sjL
n5iqhbPXDvjMbR/2/9kIUR73LJ+KFjkgccfZlgXc6sSFkaXuRCdzOH2f548qHHNF
B/0HermuaPSiy8zm3N+B6nJc1hAawSwYA6qwL/MxEt+Iif9gb3q5QAdGxyyzakGf
XB7o3lxsglhlfo+7XYrpnNaZwmwMER0pY7UaIz5MJjhMqGylg1uE8OzIfEJHHC5/
jvSZHXR6D1mqpzAFPGoMx72VZhoEZ+JS8qXxbnSl2ItWt1LhJQngsF6he8Sy1TRD
q4dw9qFk1NNTcivyPOv4/WMvjscw6mZkdk+eIW5VgfXZ+yrhZMI2kwImyMjU5TXC
qVhgXM6u8VzWNkP3q/hg88y2wINm5ehU2BW21egXG2nMPNfnDE5/WqHiEM1vvaUI
SEdbSCYG7KSL0D3JxI44WCn8R6J8SSqKJtGmKcY5nhqY80lL7Jlmj+boXyZeQnDH
JK1lmGV2PcNbrVEj1fAwPewEhsaVY1YhZF4hl8JiW/YoLrzFiJZfySNYCx7M2yVL
bGXnfSQQDKB/TKtpJtf/IQmCZBWiBh4i4EElg3RHR5qFO/DwOTRApBICAz2D1OUw
VTSOJQCwpIUdc/2NHjaJDKMqnynOBvw9+u5oj6vn0C2rbc1zar2BiMUHdH9uex5d
8AHw5s5xMRt0ZPGVtQqBo4sQ4HibRREzqL5Ly4pcY95Qwf0dDEA3o/62iT51cVv6
CF+eM4xCxrlqTJ0wOxImsAKucp75BYOfhZxFCMKud2nlp4dAQ2dti46UiZcSg2FY
Pz39VwhqcWQjhKg+djSokNkyJs8xEU1ZBVgZlvpVLNE57CHKQPAFAc/tCRbudBXX
UZ8ngb0Ufkfskyl7Row4Yoi83p0JdNBfPBoxg5TeOblU2fbfnSZ8IDbERHBGpLDV
hpoL7x0fMeiEAEL/boffRioccezfwrBA9WWGFY+aLw8Wzw9gcIduHhVSyxwFp3SU
Qksn58BXhq1lTx/LFJN3bZBeyYcVgiC2G/UuE+dg57F3DoJOGSBeaB9duax2OLdG
+s1njDlMwxfaXbuxFyRhmFteF3pcT5XJf+7kYAK1UwR8Tf9UT5E2i21q5feQttt7
q3oY9ku9BBefYfMY7z+Yo7us5O3gXq7pCd2Xo0IaOgYx9nwr/hOknc3a1nx4QFZX
U2XA+Fmz5xFG7HUPxHI0jZVbvqI6chvhCn8G+MGnvxz088lRa0rDmsj/2U7qoVKf
Ngl6hcQZ2y6bHhDZlOvFQYeq+wIeDjsleL6ZCUdJpSmrQYJoBwBHJT/uvrVz14cW
XXfRzP+YlepQ03CQiG5bi72ZQ9xUHEX1HbUNcGHl4u2aVAkGis8zNr3jOeDCjsyL
oAI/zLpFQvbhcSSQC4KrRT5G2nShNBuX6LVr9DdZYxYrWDTrHw1CeUxHziIyyY1f
bX2TwHgIvUSBd8YaQPU2E1LQZLHMkqVZsX6ufkGEDtYLGJp5i7yGZEjcgsAlgYJ5
UZj0h+JnRxlrWXQCki34Nm4iYgFh7ZAf/LDeJSWtRyOOS1GSElWrdZxHMZw3ArBn
mhnVDBLryke2axtLXcA3gqA7UWleb5KIKcl9Yp+ayrEoandtqCNaU/ScuLZDu6EQ
qJs39OgWZ53SnCA/TJzI+8god01pX/sL/b4rGFrqKKwr4NMDfUj2Z7Q47pE5vlO3
HwFg+n3bQLmZH9hXub4Ar5M4Us/rsnhpNgnAjgJ2WL61mSiWtCaxwaTgx0swIEfg
2v9ag9j95XYN/LN2P5pYlUi0Mdwvyy2ePYYa8dkaiEHTzWtl1SFejXv5PJ/RDSQI
KltX0y17gSiiFmOxtRQM+Gj7sl4uLZ00NCu5q1pMowpTHcOKaaBlJeszUEziG+V9
6Vu6FMmlRg3UFDCO596+O3hNbG0NyAMmKzGsiHCBrXkmYfW8hm5o9BsWbnT0qzEE
fGz7mppTOuzfsPCYvAQSIr/xoSODXkyG8NhF1FMniQFjdnspaUE1Ruv/zwAW56O2
tPqsRaWMQv6a4h/OG8tZPHiUa57FLgyHlZlIFQj2eGsaSwxgDcTXYTZHnOurz5pL
o05R00T3J8u8zaYWzw9daUQ3Cl6pP1fXHqujKdaQTePnx+AWC1mxGuLtTfJv5uJD
jTZud3BJklYIqYZ0Xqn0awvz0WYjC9hE71Z4GySkbk0B0QeTloJG0KfotJ9IwYJH
g37a10IVQO5JSHa3m8fBFb7fW7m8eSJRK1iqHbeut+6ExDxAApgewEihv7ADbLz4
wuepcfQzNkswZRkHwULOTUGqbYn1eR/sRWQgVZQ/HgsPRjJmCnjbfQHioivV9hcB
264cgL7OfulAFDgjOcwyCxk4rSppU+fZYUPtWft+Ea7CwM19/ZUlv4rUvT0/9+m6
TkWIs79aGAoaB54X/Tqu0h/vBP1ok3gX4YuCxrqMlsLB2w3uEbjxilMkilPMvpMc
ZHJD1Z1UuGxy0UrHXEwBrc3p5bJbH5/HO12gPUCWHENdjEYxQA+2T5JWOcnGw+ur
BVVTlL5OO197+QYjmpg/pGJ+by12lVyfq4obdMVrTzust0Vshnv6Bx2eUkoLud94
lHWSg/Y8K+baO7o/bThDN31t672FenZj8KuKiNGhehtjaRGaepWKMXf3VWqupWp3
oTqO2skoKFoKV6Cd3RFSijEfOdrn8jF0Psm7DEdVxiXxsyhdp8NXsD+HpCOAGN9w
0ydNd+ftrnZarTrHWXeEi1kBsvXhYY4zITGN30Hgn7w9ev0NeGI93wgFdR4Gufiv
AIY+QK1XwwtuSCqdeyZB9+YjJiMJpjvrtTs7B2x8RL8NClBYyq6LFVImDX5yeVPw
f460vAoqHiPWO26WbZxhGwV0OtWPr6hrkcNBrN8EC0/nt2o2jSzk1oplPBTl6hAD
/y0waB3OfqZ+j8wFNv+rPkFZZTy+YT4xtdv9Kt7M1B/ePKCP9MGd2rqE9fRPCCD6
DduyjJVYuxSZg5wJxK44V5a6BI1BifTNz4qt68IwuIHiUYzhlnL+YPcQNaz+bA6b
JFkeAtWZB5Hddm7ngJjVeBKgsI07neMMgibQVgTR77bnGJ+gBFA+kBI7yH9vBQM7
VjF4Ir8Np8JamdTYFhTe/4JtZgKf7/kc4IGSyDJnXqqsqH28xA9f5/GUH1163hmn
NGND3mi3Zf/A6h8OlxoxHNsbsfgEgj3uJpfoU/JQVLNSWzRr35PYH0CJt2gjpQBy
LNQKVb6Z6W5EyLyFBJjUeeEgPKwzOWQpgJjkC6UeUQsnMffgEgZZiNyUcHo5CHAl
m5RMTOfE9pmOqdHvM5jxrwovcfDfeqsTaiDebahxNpz4OnsQ9dl8ziFD1u34W1Mb
X5YJYUCju3qpPuJTtRL9+dfeK8jC1XyqpU8ZEzsLlZKsYYCQGWFrRZzBWnAOzNO+
CIF5UVNnPSio30bwBeWMPvhUOLcoyjq3DeqCLX6HAvbTU190+eUHqWjY+TL9lhGe
KplIR2xabPWxjvUGMJh9TdiQQAiQe5s/nMG4/fONBvUYt42GkgbbSleabY7vSJD3
RGOfNim6sbpGhs1eC1TrumsVGbJD72mXW30UjSkYsI5dyKHVWshosLvaYUrCq3Iu
t1ddTvY3p4dT3EcAdx8nT4q6qRiAYmqXi1WvpFLeqxHFR6BX6eaSW2FexNWWgOKA
mWRjm1BLkdS30yIQGkjIAj/ZEe9k/Mc7wcuwwmBjM72VPzC/smaaecTOHa6yhJ5k
fAt7SGz8616ugbNzzsZODSX/5nqaHf0TJ+gO0t9wYt+NswcMoUnxbJ3TY/TXxOI8
oqqhJ+gmL6/aK6MXJlAIh61/Qc1SXPoIIN6EZatyjIOZCIESMxBcB9D50MV27iVU
coZRoZtRnxAAHNIQsbVHYe3jAS+tBPjMURXE7oy5zO3A4fPPOug1TwUohWjEnazP
Ix1TmrHijlaw2AHeF/EoE92oVxrwJtm8APpzQs6JK8TxxGgSFa/ITWPzAuIn2UpD
gjU0bVbjPbPeo0qdp6ZweYp4Xp/jP33+kQWdhNlIE29Il288Ar9JNepM+iA82bMz
wJVmFfX8tnmcyRWyeP2canOtcvLnSHenykoJGqtJau7ifDwNbXawE0tX68VqE97r
dL5k9FDGLbPozLk8A1Bl13HVz7GSGHclvbL5O5b7GhAkFyiB8D5exQwM0z7P36TU
Q4rGOtSbhjsbmKJBoFSydy3Uvvc0sZwsGqL1wWt9vRDcf60/re4gz8js7q96nWOX
W9lGpudNSc7VCJLBDI7IdXQSjjVa4R4zLP1qFXXiyNV+R41hKAnvGq6y/VAGSZ17
pu9EtRHhH5E73/IYqFxLP96vm6LrSxKAqWQZen0tmtGFD07tdxJ3yiaVRLcnzqSx
TORvIkX78wNQgJAGrwU230aF8DCvRspbF5wX6DFr09CodLN/QyZnxljr1nA7YdP5
++L91K5CKKkNEPNS322vXmP8QVKtroS67nPnzg4GJnBK8CbCff8j+tpU3bNROjoY
J5g3Mx1aBv85ojdRNLP9zYaCiatBBwMzeEHqFd+P835uOrwb58cSQKYuaED3ToO7
/J8jiQb40Vl0O34bcUNsyTEaW30MdaOmUnl+X8wZA1GJfkcRkvUGkkevUk8fxgqs
fo46VznRbMAQBla8p73Lo27rIzV4WFkfRiKWFVb84o2BmCKQt/lb6wnbQYLMmcCn
gVHyR7PgC5cvWeuJMr1HxRio7WpHlY40uyP6SS6RrX8CjaNpfOO10OsVYNyyyWZC
I4NNpug8nv0ggenIm6MdRA7rm9l386FFqIzopmBNVXH41F1zHcLMJQP/A2eicli1
Mh0yjUwDO4WMs/bfGSB//3pXEL590/kd/VOhhxRlhqznwu8h9ZYkVlItw77hiKrI
sNhiN2V8YY0zUqLEm7NR98IAsghsZkkbNkvyYBvj4R8dcuMhPzvbeK6i2uO1lfso
LRraONktisNwsjvMgKLe0YP1EZv3p2SwZKD3QsKOYFMrJkwIAuEwfUfmHfLAFkyd
zxfLhYQSluE/y0baVmGWzrbyvAqfhcFcJZRnpo9k5p7bICOUiA+an94YCPGxrrPa
5wkvTqXmPM1RZWqHMnYYNAvq90r0hiv2x/HX3Cjkk5rYelUZqprj8yyCqZRCGUiv
Yp/BGTBkIANEJHUTsXP/egZPhKDLJ9eRLKgeK/AfIfTHMW7Aokupi/9Lb9Fwj5AK
+v8wSp77GrXzzPFgsSCnCnmo1gVf2op1FMl/05bdr9EwcSlebzwb+gnTC4zd4OYz
rkOCfo6tnTyI0GL7x6hAIT3aUe1lcVGbpWaoVnmSQ+sFDGGsJj4BXTWU6gXg5qjp
TgbVKm1jmHQB16NROligl+kwUSztc+STWSTQ33z1agDWeuw8Uta+NqCTS1EnMKf/
5BknRgw409wg0RWqmFcR8CzKiMaYcxfpiZ/BecruOk/fTqz1m2nfkcdAlOt/CBTD
e/Lnh8o+CHVvT5qw4dKXBb8l0ffeyKilg0CYu7r16piHxqSSiOnI33EMdFPHdKQd
HmVNqIZRZl5p1A41Zus6ygRu/+tJ1yaEGrzvsyGykzWgCDZJkxyumSem6eWAH19T
8xnklulDiWTaVr1dwoAy/RrW/LXDBXM2V7SWHHAGfquAl/B2zbt1KIqT/xx63hU0
CZOv9J4F4g/1yKM28r+rBDsnvOYjtY0H2iD7tkRdRAatLN+x9OXOc0z+uBu5zTNc
q1woiC0NfU0cRXmBilTRC4o/mtRZOL4GxBRlrDJGFd/7bqi4UzgWaaUwG1uLcBY2
E4y1Bk9gXsl/RR8p2sW+MrelJakBgTxURsoXuT2WqdYPA5u7RT42zpjtMkI7ndHf
XKygiboTjimwRO6ZDsJJbdIP1RQag/2yLMgSwocBu4/DxrL268HbZBcDvYV6rhuq
WIR6lLqqyBgnlzkUFVWFPoqwaOcGPyhy+y/qW442iAEvUH0JvWxMVWBnfq4MtbGn
XIdBhLC37p/6L3OEdA8Cg1O6BAbZzh8oQ9PVZQ80mtjkCmaGKlM51uI/89ZbxWoV
IP8kMmJmcWPsCxo2sYIgl69AicQPhpuhJnhjyCZoSvwpAqV6p64idtrz1e/9gFii
dEWBtuZi/7cotorS7N+8JEADdOhBigYH1UIzwn48L1X9R73y9O0Qztiw+PbRs8mK
HzrsdzO9IxiRQhGbPrIwGevtW5+mIJjjvP724RWkLWmvBD/Y+4oVUXl1NDQxYjIB
6uggpTAw4Vd2xdm7KnXxTFxzgoR0EOQLFTOabiCWJjSbR/iNDEMqLCdayqxX8Z3e
NHj+ImKiDDay8+2nDlibvkqBs4bmqEOf5BgqyHQkx18GGuD3xY6IyI67J5+z1yqo
1xhX/EQ5RImVZvBNs02j+Af4fMYpUb3g8jA6Roc0JzfsIBzIas9z8Y/cHFg/nXHN
hojlXSdoSpqHG7Ecgs1JxAR5hDhQvfDQDnipuvrU8TdO9QwuUdMdy4wRlQ0kipUJ
u0ZOPJGK+w+05h78m7P10a4rsQ5QQqHizwYLX0bY8RU=
`protect END_PROTECTED
