`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
thhNMPaj6j4sRqoNVrNR2rve7WryAdv0zX23Vn/cxk7wgHfXOpE1SBkxCdaFhu6t
CXMmNRVPV8HthXymuq6Jo4BzbpNPBvXV4pcZ/YyhBFH9JwuVU2ReSgajlWmtafSf
93DRRhfR8aGgI3b6cRLt4Td4Hnf3wJubB0vTsMLW4i8AjiE1S58OL1cPs/LVQpxt
02j6wLMeVCJOaOctVJooESfUIbqqKzjsVTFR1484q0QHGRiJEgVjqaTMcRFJm0QT
2I7h45cB2rEznt6Hvcjum+DVDJmcyq5sHqKsN/LpDXCcudkmKmrm2Gle6ZxbdCjO
q4t/3m8Nrnkwbx0iEE8G1NWxztFoPVlUZ+qEoqn/f/42rEWk9n/W0zcpEoBzxZZ7
2XQIFdx2v9YvwX8Gp8v8arba6wlwJjwgY/aJG19lZareCAzSZ1HRrOgE2lO2jhaG
Zl15YA9IuZVyua7D5tcN3BLsUG0nuSmcxiGmAZL77Hsw3f69xlI+FqkEa2NN2g/Y
1HKMNcemcP/LoaCxIHNonWHQu8Zxuip+cZHXstkka/7lx6xLwiCKSnwSA4KPK5LC
k9y1cQvmBWoAJUTLDyIk3w3twNG6IjdfwUD1tpgCUcL4IP8y3/0+NPh8vDUR7oso
O9lWkWm7Q0Us6yeFHFKrohALbBY/YZTSuEPhAxeW/zI5ClWqBYYUPzDVhCaS6j1k
7a8z1LFH7+3Bgvfl8pVfb4z3T+NJCbPF/l7Z0EPJl8eQ4dYS70F11sP/paeMVPPW
t+oSSYLB2Kbry8dHJpekl/NIvN7Viv4cFUock1046sU5uS7ac/355jmStpt478SR
lyZm1y6hTO2EqYqf7TNMAeMnFZ4gyZSvytqoF886VYXTO10biK30L6codWf0z8LL
co6WP6pszrFHz7ZBNdzQiRpKaGtbVfAKm1qUHZkUpxTbg4EJmRURA5IMnyBBN0ik
HiaOPpKjqOiV0Ydgb+DLompNKrdfRiO4WzqKS9gdgUbemSZudlCRK/pZGUDL8rUj
9jdX0glarG1nhtKXHptgVf3IjcUyj+Invjj7EOKTfmWXAK8+ce7XnjN6dtXJW+Zn
innXGeB1UxdtwivYKfF/1CzBigPzaI3vXs5b6bF9ATRu2W6KiqawbY4kEJkjbiSS
NR0Nk3pLb4ehTeRgMF8pTayjw4JjFRFsFJODXDjNqBpQlMrzdXBUKtt7myhuZzZf
cwJdaRMIuOA/4w+HkydaqkOkGXFZe8aO8i7IDvs8M22d2F88P4FGXuEw7eJgtuZb
f9cyCZc8GDE0y+1JsgpStcZjCc0GLWsvcNVHfONWDys33/DqKKUR3f8AzmMfv7au
i1hwYOwme3hkdST6cnMYvvHGUWtOgSrogVdkJzj0/uEYHzIHJSzXjOwwAW9cnShv
hS9jzLFWzEvFBkzimW9QoqM7WBx7Wxc9tN7AxFSCrQDajVG67Vbul2nRwiHtf/AG
afCjnxb4qk0y4QtTNWsJuQaZRZDPtutrObvdcBeHBeYEgLmyAfDHPXgoAuZjHZMG
IcSX1JTzlhkW2xDYMketUITpbOvq5LftjfOVxfCqwJd3gR7T6zH0c2eUYvn6+sj4
rG95QzfnrL1nRvqNmVYINtnVuLv9WTS1xhBc8jJ6zJAm2V1Q1DqEJIAPELMV6lWS
lv+pNOn44OURfKTKKvn7jo/cUQte2M6Xzd9MApS0Iaka7b3d7CK+OBipY+M2YB7M
h6ajGfVWl9qjqbA9mgMlMJKRRu5iB/BQfBgLIHhT+7waTQZ/+bxtJwkkNaWJHxZt
nPphiFqTDYOBrKhY3/aApJLqLhesu9N1HXSOEbLNvbVYBh/X+QLDKmNst+2lvIQ6
mFZWg3P/QOmgfScU4N0Ux9APIT4IjdXsCVBSzx8V+ZwvGoCH7EPoUmPkj723mSCf
pekJuabOze9w5T60Em7+r1fTe9Lda3BPgedbsUf8yjekWv6DxpM97DdN5oJPCJcL
pw7r5bm4t5k2JD8pPVD2D1tPRc8runbFGCqg3GnwLmTPrudPteJ7RDT4lQdeN8vb
7CVx/WSJ3uAWX2GYIycKt5VxJ9BRkIvk5pR2OxHr6TQBx4hQ4lTTCjlarpoWYSlb
qAYiVXm6L+p+ZfHy5vgzFx0goHAQ9zP1CRDkHinxv9Zdg/VylmNBbLzHgIWwD+l5
owHgU8dzk/UZP06fXXYLo44vahWUodIpcIQVf9UPjsNqsU5Zj54SOwPi5dpkGNNG
5SMw7kbqMENm57dtRp/W2vl5ZC5R08T50Vaa4bycIsZWCCtviyvwIozafkjsL/Xt
EZN0jOtmjjDbQP12pZYUqBAP6vJLQwgmY5pi2ZaWfcc13QUCY9u4od8+27H6ro+S
wk8A5nCDeqpG7GgAe25mmyGOWXu6+vLecVCsF2O9e0yrGvwZdPCYM6IaLeiaTYCd
B4SziICWEWPhkJBU0rPkIKu5Lko98kq/lPanSS6188v7liTOUB9aYWZiGjgTXuGM
KawFOPOsNZuAf74GKpjeY8cIr+Yztk6aRVPWrIKvojYD9LuVaG2yphafsqb1RWoz
VXqLQEmE+bgy4tNHuh53OgMeEtFdR3Orw2VLctMrRZyGYLeVzfhqrmvBAAIPcREV
E+xOWHaTNgeGHT8saqBgi792L+0E/r1yw+SoRCrB1IvXv9lP+ZopLkVv/cr6uBk/
Q6VP2dHan5kflqJ+/ctyaS+o0GcoxXLsMRjWA47GUUbBLsSMXbWh5SiyWUXMn7jX
6s3xLL3LumgJH68r3FUeJmgiKYbJTFueZhz0VboKOPkjgoZg4bLsGzgiF2nRIuQl
uLiSuyNwJrgzg/KxTvpFbE+x/w2yalKtXB0Xc9Ymp0BkzP9pReaR4PXRmlbnq6tT
9MpXLUPorDlregiaRxgReqZFkhVXXUVS98wtE3AMmRvcXkEAsHei3YqZbmXeiYQa
Beh2TyPkh/GzWHEyFihjDpznyW3G6FKRgYkQjA8d2AiFyz1POBbuphkUMyvLSfQN
mnR82OwSUsxao/uK/VlnaR2v1VpKOlJRCIJ5Ewz2TxNajORfXkqeYnRO5GmttAc6
ciFBwKj4qy0lbBNo1es72eQZnQH+t37FF4HL9LBhAQ5nh4dZl1K0JMMmX6cI5406
3+G6lAXUwn4ZX6rT805cfAUoQs3laNbI+fQaisH21sOEGgCzZYQsYVdlbrtGKYA2
bCOhVvab0BGIyvkPX2J6N/+b45ZR6inH9gyHi5658Jj8xEam1u6NVBwNRYL3u6y1
zer1tvOCfTE6qtSghzrr0f4mjfN/IwdgKkOtmnvAwBaqpr98qbsA5gMYDhmQPzex
8hqhTg2lzCLkst6AzD18yejChHIDR7hFq/8TJkJSt4OxXK1nk7xqRgZ1QIVCGcqz
EMCJHfbgufnRBzRUGaAuaLZztBTjHjizy8e7hvMeDkKkjiu+J+geQ4ZV5xkOUUAM
wjEDwVzN3lFk8M5KssemCTA9G+zKFjb8Yu6GHjJxrheoHZOZLp7ZIWy5J/pOfMG/
HXx6f8JCnO4fkBhN82abH+FSmcYRE8nEheznMAv238ERqguChWSuGdplRRZdI0UO
QuXduONqDL913sFnb111mnu3+lv728xTFwT3Ak/5zOcVJT3aVI+7zJD81K+f4RRk
0Zt8vTIf6EbSfQ0xSq4UpNfloO7ljV5g+WzhyDq2W5HUddOu7G8NA0R6vLFfu1eu
l/LnfydlFI+6IjJInxL9bJcH/gSmi1dJVM6Xzhw8y+tpadOSToCCV0rIlL7zfMbp
0Cuzr1LHO3/Zf7XtiIh5iW9zuJCeeu6GQR6LxSSnPKn0902au732d6bkaCd3zsgw
bKtYWv4lkwH3+M0y4yAVZ2FG4wDEbMSz/A8XaYldEykplYwJ9dym94qvMzZmuncD
SEcoDrXSR2ECLyh7oqV1pnBYwyT5Od+gbKpwa7lU3IHqlw14c7wVxwblnqFlBc41
0nIeZ+usSVJ8QmrgbWJ/CuBywvMlI605AyOKWkj56eNOzZ/u9yP4GK8jqi9eDRBm
2AQH1/EP3L2szAXSSj6CFWfaA9FG5fk823tveZ9lGCqdAYVPt2/FL2grx2KYtIOP
S0vnkxccp44oFkcUvNKaa3nhIRils8EM4+8eLSyGGsc/6+CD7hz9zLKqlwrZFat3
Q5/zzJMHrl5AMgVHyqT39MDU8gaL+QLhLkkCKPdGXeJ2cELmpS0r3f8PaL6+YMTq
QiWoDjK83OuEpRU6kEYZEr+vSJtnOBYATfT3nZ/zcjtw11Ytv/p36sVacp1jyc7Y
jkl38W6PnfI3Od0z8TKVYKMwB3+wX6gUK40CCNIpD6wEe+E5F+CZjBFYwuw/zT2S
wIKRw9aC+pBvdN1czmUYePNAHcMaNfOq9e4jVNCc2RQ4Wwdf61FZIDdRHjv4zsjo
wU5Qzy9yVBMxXvaSMv7ji2Le1UB9gukY5jM1ZtgfBxGmZXpSwotWTYVoFriCuGdG
ZAnJp9BTtLi6MCsUySs8b5POG/35viisCHMEeO2SZjgSAGyxIi4DiXUMPMyKJpJ9
zZ06DhNFZ6Ucn+Wh3iO29jNH29zoApZ7EJ1yDCNWoQKSCZyzbz4RX2U1Lb/qZHc5
i+L4xW+FHixyYFHDj6XddffzZdsFkGObuBf8YH7TkhqfQVOk3OemtaVxeYPTRkdB
IGI3YH0cJnQpjBsAAcNcqMrbFchzzzlL1PLifu24+rEueKI+ZBNV5WBr1IOdBcY6
pU9O3eOpqY6DmXRwMh0guh5tSlty4kEm0n3cJXvXfPaQKWafvVKxqdlNGm4wj7KQ
mZ2hBhlpOqJI7D6khdiUylqAZL1qP0Nz05al3J7VPRSD8ZUY2bql17/CLtM3eCrS
XZuEj5Pq6NjrutK+Ra/c8igGCWEfU+eVMqOPE3vhNtttccX7amX8CbUcvDtpB5OO
UbpPABhPxMJzk6xrngJepw0oXcSa5luFg6fjV7Q2j3PiGNJ7/0z0XmvnPQI0YLIW
I2oeWwSeuRoOW8OcM82Y5pUNc6VWbH50UmpRg4gowLt1tb39UUZado3Jy3Rg3eq3
opLgtmcRS1t96FpBy/TRVY5+UBIxEx7Kk+HCD2cgsUSfLlrtiL1LPU3P6r9/h32t
jDK6KB6VngRH2mlZ11uLomWuwesp8j7bB25p2I9qw423+IH6SHu52MFfGekxFbbz
FaG21bhQ2jcxYmGHczs36wXkkv0ABaKNcZSU5pg/MR42BQ/DZXTsdfQTkzHAK8nK
ohFHN79v6dCSGPxJdKA8j1wZlzaLRQga1PNnVSk8jsO+FvJORq0jAmZx4ttXeLP2
L97YkcA99x36pDrgAxWMgabW8z0LZlctLzgdUhpeG8tx30OzY6Hs6Mh/CD9+3l2N
7FMHje/AUqlyj/j6YL+2WfWi7CETWqqQBor8hlAOaykYIBa0ZuFhp6+tJE6BmUJv
W85iIfDYpP/po2+VE3IRyw+YmX8p8lF1x5yRzC3YNDO7tlfdofXVjV6e9258iQQV
GyBxI8YlZ0V77F8k8UOU+Q3Siiv7rjkDuRZ0MGSe3cuprRbzYTYZp2zNc9ZcHcY6
QPBV0lVbwaZVuwCxREHY7jKW+p20aDQFsfxIT8ALhHPsogEQGMeAC1x37jA/7IA3
ZnjBEZIqBiYbtUn29sPbXrVg80QnNFK+rXPtChm/XhUImmEc7xC/KhOqG1NIo/GC
WOXPFUpKuhMRPsD3EQzr1NDXqOMvTJ9bt5uPJUVcIFykBQJZAPeVGqNiadEaf+B/
C69AU3HV31KXSTUjVS7UqbnupvnYazCzK+PJY7Gkk7bnRQxrmlgwq1UtbBu34zH9
VzR+ml/H4S+TpEQVtX6BP4mmFNZPr+lzUTD86/7fHa0ok/6wh3aftBmKbxY1dB0V
VtdMKQA82mpiWGKiKtd15VZ+ig7cZWXnxk8KQLbuhZxE9e78+AqcqZj4QjShvEBS
C+vptrvoR1m4+8VPkN/CrQzElf7aszmqVRSmZo7g+eUNIYVqZ6EU6qUEM0xoSjqA
OqTNhdOgN8xQOkIzlVOL7Fc0clfxCQ8fW0+9cGZeJFkB7SGMnxpjT8j5t4rKdg9z
MekA+NpWoOmlWDH/LPPitjCP3+G0UUYxSdhUFYZzdtgpHuGUx4mazhNQCWX+xVrY
ldlxinI5f6FYApksJwXkJQa2cmwz465KuY/4lZ4mrl8rFTtBElALQvBliilU8UXD
hrCKrWSjzXzPePXoId9bSX6Nsnuf5bEzxc/m/Een6VNONn+TxhoAkaTNTgeNyTP0
O0b8K0Dm1s0Unz/XXNqdqyscIb0KkegQmiR67DgjvG4XpcaPUf7q3dQUoWUR227h
d854n7exyI2go6T28NpV0Mhi64cno7D29rBnFv2FPE+fylcaCsbjj1Yc3MCEWyvZ
QcmK2imJk65sbaMagnGCUwbtAfj8cgI4nFtuevTMaJ4XAa+3S9mQ5ZzKFfLck47z
lCOSMY2ocd5TUPNsR9MpqpQnbUkSy0fV6VkKZ5PMS5vlKrkDGOcA9Ul2iStSFBU0
AzxEHJ7lkNhiyL9+OAjMoRLnMh+1IPMqb1FlPa6tFu/1FX3QSx978RvE5LOi8XlY
HcaaMiWl3RaJQxrjYwAjqvsffVury2hjYqG65lkjTkDST6gJs0mIR/4So6d7R2r+
3aVpDlyoT0SxAspOQUnst39191RKogTE+clkBw+bSJFm5YrZqTxDcnF7MeyDoCaL
afJaouDihhD3QJgkvzR61u+dtrYglikkFBUFi8mujgubJAOEziBrv4oci19UhIm+
lrifBIzXLHHPKeiKOsfiDjj02qlCGKGVUJMfMfQcQfzTWloVX/MlKF6Ug3kaMoOL
QmuDGccWlgZOQu0VtWB/qaaAtQvbUhuzsQqQIbvKKAkdL7sJlC8nZXyuSsZMtSkl
DFPqDkwHElSVasMq4DpZHFlNzoMsd3UNmo0b/KCO4ygmw3TC9aemc6JozLTH/H0u
2WbsqRytZLIeyGpQE3i3fO7MyRZtpkO/INzqLtDKa0AiWFwDK27QT6GPE7ZK7j1p
IaFaxkhtwc+B8lD0u4TD1WJeETQJjug09K3Br7u06xv1B0KxDGnuelgi3JsT8JQY
i2Z4kMgSKMNrns8EEYXqCf59RtK708B606SU5VeNNK2zkkw/nCCm7oE6rasw70Dx
BU6IrdfIm6i4RwxKPnCklNm5YXfdn3/3rBcFY3F8B1jPnmMY1rCOW1466L59v2cG
ohxh3YKwCESKjCkyE1DANriMCmQbDbvMP10ukAAmI/gfnuzFKSh+YvG4QMJbdRDt
irg0HAanRreprBcOadfGcj2jVgnw1RDOPaREvdTayu/tqXM6y+qnS5iRmLy7zoc1
NVvcTCwvsOfnYl1EPWTu5LqfOqyaLBY+IADMqPXJrixZSgS5iF7BnKwUSYDEvN2+
XmJ+pLbyYZ5rmWoLCcw7NncDqGIH4UfmkY9cSe/lTY86gzYBmOmgFw7BwN3BQXos
hd3ds9VA87Z53YMQYwe4rwQMkzTjN3ln7rk4BvECNjtFOVUdSo9xYjJXZSFCKIot
yPDRFcd7V50XbWkefFhaTVuEur/Y3gXYwQXkNUEJ64MawvV6eDRveCvnx5SUvbbf
pPzKkMBfKcUGvrJ1ugs2773WXtvy10oT+INs+CwvmjMA533PDqovd0JEdd7Ahemy
vTYjitpCdgB8waNyz9mmG166uGEEWuO5lRFN9t0ZPhR69rf8wHQyCKMIj9Z3C0Rl
rbAQSVbjzxY2FUkF5zPX+LpVcaCDEo5Ra9J5gBlc8m/epgTmlzGSa1ExfSkaqPTW
t88dwhHZPP8L6Oafy8A8IL67wFgo24WcNRZFrbcr/ZGfkASSnXKR3rQvdNmf7YOm
Ur6NDOfpAJ0LECDK5JjeKGOXpbV7XWU7knpkFp5oY4XVsd6I0mFs8WCelQZmLN+/
zxzj17OWgL/Jhj0E/nPfzzKWYsXGyKUsmQidXHSRWK4i8a7qLFM5kZRrAAer7BtH
W3SsVNK9KQX51kNh+5kpn4hK4M6VPVq1CWn9MbV32iuKiP5vbl+UggcukHN0c3TD
hwvrucbAjv6/OsjsNNPy3zRGahe8C1acgx5wDPc287BaSGo5qyDU927ocQsKVZDu
NovGnnF7tCnh8CdoC8tBFU0UEYFlDw0nfqEZCMcHbEdJGr6qBHF2VWGwyly9+CtI
fLW/RA0oEU8bhdP6OMmXv0mYIy2IRq0a12wr60KQ+OCGhk+9pSO5I0tXDCArjynr
jd4tPinmIbIJ5v/pRqlKRYTvuHzgt/29n6YEYZp6RzD83uzb2l+7bcOMTdkTEiLg
MF1oulKqOxXsrdA7Xc6dZG4ohjBry5qbR1hHctTOthL8bJ1Ui+XZ3ioru//jPLkY
qlUK0JxeXFPuCHR0pRK7HBq58oNFNqrWdceut2l7YgMFAfIqQH7U9ZfibE8V8ooG
T62zyOeTGDWBeY8B68ZxsveentTT+awlCpl3AW4eas78sQx9BpRyprZKuK4dpNzG
odMfSM3RSFFhXWYAJ5OvdivT3qVqBX26N0meEZb9xzs1kVLxeLK0i8RYYl1n+Szx
kRz1vKDqdCAX3GilFCkG9YcgGfGZl+Dc8HEUr354s4S8/dDPxsK3yExXUsKA7ESB
vFtDWvStebus0xvoUmx17BLuJ7e51BmpYV/VeL1tw3OZst3MklBKklU1PEpgG4Bj
+A6EHEMUcPVk/IopgBdfjR/3ZN0qtAIF/LbYUT3bmijzJmbwgCdD/1BiQf4PnvfC
J8z0jbRuwF3yOz/pUxnVaj3sGNVVjw/ewNRLwfixTTyNfMYcHQgReO4cOoAdX1kw
+q6a8p/XrX3lyjDAqOj6bCRxqDHErTMinG+y623Gd7dxWRUNLvEbao3M5/oXTkiK
`protect END_PROTECTED
