`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gPfEvXlUUd9/ZZRqjja59vMhMslQ/WGtEkH1Bscm5HseO+brIYom/P4CNDMxpIX0
owUEJyPGD1RKKQkv4bnXIU8P+IWtQpi8FmwCF2VuOlDTBELiYus4ce0K2Iww79O7
MoXjsUg/+gRn00h8h/jzLbRkcoj/nt3UAAE8Gf1pw6IA8iU+d0o2oKYUlxdekqeg
9fk9gCU1vi9sXYAukoq1EYst2qm6vndR24SLepKOs8Gfq4Yxam4Hf0yMHrvDEWqM
iqdaPGpnqR7b7vevLmDxUOqQk5eUV3J/pAHGXnzSDeBa3TTd5YX1bv1rZE/8Zn2L
MDbL1pXa3qwClG/3x8p5Tql+B64XqBQRsYBHiq3r76JLGgDgX1Hb51nvkxW26KpU
OL+wlh3TJA380tlWOCF3NXidye4SPncfTEL8aG+efkmHmZz/OUao+ekOQH58ZhZA
OXg+oXifPdzYvlA/JYN9a6hYNzt69j+ycaOJbNEyqzYYU128JIiwIGmD1qStRzcj
/lAySVC/rO26hBETNFzEYqX739foSfjY/1Q9XHJ64a+ue1hMs1/6gtsyEOASeP5D
kpmoWwcdAWRnStOrMT4XnA==
`protect END_PROTECTED
