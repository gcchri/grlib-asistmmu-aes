`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vY9WhAUomkVvPr6zFuxtA1nmV5acAzvtn9aOjR0oMPitBFbZwwxBC6de2EbFqDng
OTCMLVD525D4TZHyr+pPkOE4FGUWuLwibw0kkjiBnNZEvXzQ3tIc1Hu3Ngc1gbTp
jp0DSypuysdoFmQNveYjZoL2Sfu5xWYrWoGil+fhJs5U7MS7oPaP5y1lszVtbYsF
J4iOt+aAm5CxXamzMPUcJMX6lcGOkYkNjG/0OH+UMVCNZXIwmPzYIEo3F1L0Mltj
K9Z6ji1Hw0lAv8Ogc9aBcyx5+3QU4SfeX0dlP6fEfhDjM5yXVg7xQUxVsTuK/jT3
T3AUyjOdjFKJrGba5Ar4cQ==
`protect END_PROTECTED
