`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OB2i7WKbXCp1llh6s0jQ49jd8Ks1jvOUfxX65ucpwlNTxsWoSmaPXbZao4h5hLq3
poGsR7X8+YF7++3WEEq1QHXLMox2vJwZJy0S2l/RTIg3Y6EaHUWGnM2RBvi3Cdmf
N3xwkPh6XfqDCHqw0PNMUpMIY/eGIXaUx/l0NqCogAaJvAe1rb5YjmLUJTv779xm
Ym5aehzNo2CCO4ULuLNuVneifb4M8D6j0PyoQEUFs3y/iQZnBrTaD9aeVFRI3KT1
mIqZpoxmlSpvLwumWeHi7x2IVDl9tGuBKC1iw15U4RrL+NSq9+5wXhBavPjiDj+l
WWXYf/bCELEfOPpdOzUF/+/z9HsCdZUhiUaZjmgoeR10jgDUXbQKP/GcdZwKAQTs
+jri4annGjD2hMbbIVKFgdAB3HC8WJ436L63XPT8zsiodz9Rb4+K+LICt4pgerF1
yrMp66MuO/sppT0iDy7yZlY4cNClHnzJbrd63MciIVFt65sSy5oENLnqAFS6BpxQ
vpCqcItVcyDFZ7I69OvRa8qBrHV3xUPlUsWdmGoh/loe8aJ/lnls6Och76hCJyw9
SfgJ/a/DkCHWbNVROPUVfAN3t9SQc+om+3mctoOwWftjw6kwrh1Al4gjzh+dtPOB
2/k+mSNVS8nUG8BA060ngqN+UEusrgFloVEvY7PQAQQCbDSWEfhd1Qisc0LIyP40
0ZGLWAa1frWv4hXUCVIxLBdduT1GUYIcN4UvJjhpkKRClOHbirh1e1wGHBwySdcw
zCDSdHHS80GHued6E0BOCVHmIE/up84U+kwM/b+fnYIc+Opkzvhw/s9Rm8V5eEcK
W71wcb/XCe/QMYjMFOUiNZsUGt7g7dgoWoL1V+Yg/mZ/rnIgP4g65/4riONzOvsv
vR5N+sDvho1+p9IpGYA4TWzIBSy8mYNTJ80NKjWs5QTIbuufjy2rO5wwvizm5t+a
WI6OCteyBbVEPX04buEcIs/0Ac78SGwkAxTeGD5AY8mKuSV+iZu4eS1yQU9y3Gqx
nKq59PGKsnLHvHqzOht03VseI2K5kSMEsRcVGwaTQKml/c/2TPv+UOHov2d0h0ov
QNq6fN5LWVFH8toPSJvYcY7xGnTiXKj0GkfsI9nOv1PZDNH++501gk+BLFFCNu8e
bIRZ5QjkAvJ/cptPu/GBZHh7kfAatQm0gN9cj/20vAM=
`protect END_PROTECTED
