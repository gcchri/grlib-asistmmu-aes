`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wA8VVm5687auhWUJxBgZd2PANMQBMwz7JIbHyGAw72DXkfOs4QK635Ah95RvoOhm
YM0do/Y6KmjFRxkT4tDVEfEmhF2iAbPc2Etzmv7Smk5W28jdgcwCZBoZnuLiDHoG
z2qHoiEUKHZhFgISa6ZCGHbj6GwxnZCCpoDuHcVfLxCk+DOx0H5rV8AkxUvJGY3D
eE37nD8RU50yf78mdNGCwSfXZGrhpk1UymxzyxHXQ9OcnfAhLhtEuiiFjBoamE2z
vNLgoh9zoI2PJstDLmc05LxNnv4/m8MXMRuUvM1VcreOA6a7HX7jhxNqbVxML+Ox
gShzNVoizQV9XLJC3q2rvG8sMCSIvftOWZ5DsE27u3XBci1MQ6I3K8VslFhecF0V
nF4KkogTnSdEgjt+sQ2ScprAXYe7OdHfFKJMxRNwMY3iRPu7/jY0qnjPpoJvqTVq
6M/BqrHaqj5CtHTFl6M2qEliuH3fR1ex1yRJ5vhVvK83aTc3uPxG4B0GvsVhJ6Cr
BDPj+20/jys8KZ5Coi1bHzF5u/ZlNGmgS5D6z6Z5CS4XP1GRD8tM56uP5AVOATyo
eh3/ARcep1yA7dqRjmwUj0yoRHdl3XjOZmYFU+AFYwW/1duOIorqkYMavb0nFwfo
6rnsXhtZusk3a2M6kOYWnWUfZsUiAHEXh0IoD0s4WxxSnCSPh2BnFzsZr35b5NFN
dPf7GxJCvwOxJ8YAJ6h7woUD8Ne+9XrHlr4LitPCCEWL9UESdL8bxROniG1Bt5J6
mAXghApSTjeFMCeOzXrvbE6DudFqR2bGntMZEAkUD6FVqqQxYLtL4d97Ry8EVcVX
V0ucvf8cnJ7FP3ojZHbMXddbm33tiJSu8AwLEMbZyJTfehkyCK3jQwJBATI5Ml9y
YNry0WA7tBt3XadmbVtmCoSwQFHZmEpvCHUqszC0DTrZHx75ycxfoWSIRlpYUePG
d7C7Jc0AP5wRzjqn43l6BBUJ1ac529JbDBuflAXgzldoOttXUBH1ySDhrLTNDQok
WWvqonlaXv64a8Ov/Kg/e9cc6vAWYy00pVTk3/O1fHRQTxX10ZvHjVknSRl+Hrro
njDeR/ocx/RSq5ZpKz2x5UUtbADKBVsxYQDTwEJ4i8lNMcTVcVs54vocJSroQW59
0eSre+pHTptE2LXsbjPOgRGQJXZznnznEaJwNU2TBlhuYlKgAdy7+HcY8Io0d1z6
QCgdmoS8nCrVnROiUMvPguOdvDb9ZyrRw8TK2EXV3Kypvx/OZYhV8mrps1v+zdPw
c/H1YQYr3V25GlWGoZpUy1hUL9NskPGY2YEfy2e49dWAdJ7ymAYXuY3G9SyfAoPI
DbCbRQgoyRHSEjfzGNZMnwi+VrO7vRdcoJU1B4itVBlfg7l9lBtUTtktj5AO+oeO
sQY/9lBUE86A39wSsEmhbew6dGWkZj1fK1xHK7hOTAeTN5G4q9KEQGG4nmgAnHHD
GpmgmViylTdMd2e9g40OMx3X1arYCArwums5DLt35nECboaVaYqRtBhCYVtmVhgu
fEogsTMZR/gFui5KS+WAWCBeJADZ/yd38edyvpDhuVcnRBKP6hvGthlIJJ10jRu4
7HU5Ww2bAAoLzhDKNSGP7e6CRBLRP6RgHcDQ6mdLRA9Qi1dod7/7twaklftaouzk
bVtnqCe2vNkItOhFA5fSLrkrxkxOk4qHofnJYtvwJTRS2fBYGeH4quB3V/Sg/Q/O
QtTIctyLD0IlaslkZHePellskzoTyiHiRFw2oHdkCw/9/Meid++sVIiTOcar/s8Z
6OZvElO7+XDIlG6cEY+yh4neTg1lI8bRY/jM9pEBvPShrxk+Jnc9kchCZ5y7Ugkf
Jwf3Dyjm3b+qGNtLYoMHQ98RUHQB4tjCyBIbVyZ/uTwYJUa4/K4MT+4PeFatEYlJ
vJzzQu8OXeHVoMhy0/I1ipH+bWrVZe0lDA1XG+bTuDOlKKkY7EcSmgjLq5STb3gi
KM7dxUYwUcNkdhmj5WuXAyCZIB95+yZWZDInBW1PsusaznGsP6WF7ZRtoIr69jCr
B/hXI0AFlbcDPVZJPeJtilIjt8nYThmEHFfiLxfafpZ4KawLnZr3E7OyeBv5UYHN
3FIH4RoM1udgPPMuHnmZp3Con1PCjLlRkkLyv+06468BPINBYDBdgHlx8v3IH8ft
kQoNZaHqoAX8hem4tHOSpuI3xJO4Mlj1Uosj9UGsAIkXLv5YvZUIQIcclx+hqDUg
bHHOziWGOaZXSbLc0Imr2O39bDjS44eeI9TQYANb9+TwvWh/fiX7cOp/O8H7ie5j
jGgSokIw3+jnuxO3z9I0ySjb2dJZkAtnAs1SiVgpr6D1fg87W2WfAWx36RzXnY8n
gXEaYv9sNUZFC2BBdzNDve0FcYREDBTqKQ+/FJe9D+WIzMlinhvOMvpe7nrhlNA9
Lkmu6kHW5SR5OQVWDoWlNJuM49hTcpbWX3LFZFAxH0w=
`protect END_PROTECTED
