`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rIQW//aSCfB3somu8yTAP202T0T/DVMV9MrMczgA4j5e+mFGP1dSNCK3Po9WlPxZ
LdqV6lcS+m3GrS0CNC6RlTF6bkGZZeux+BZfSGcz1g9OlHid3AIlRYSf2g9GjHQl
7pYFcUtXQqHxlMmiwJyv6JVbclqXlRyqAn2evN3PH4RSK097mOnvWew3TtDlfOPf
fSzOgqX4Gc9FchxE25QkzaoQoRGUKL0mlRmhjvOelZIKk/gVZW4cRNB1AKwe6g5P
wITqBrgPhWshKmKxM1cA0b50uLj2bT3oTNUf9kQ1wINuCTg7v3xDmwCL2e7oh+0Z
`protect END_PROTECTED
