`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tCe529g6fkC3IEyorJGqI1nN3tennsMzUWybTYaYgexZ588AefCyKZbgSrtvnbci
HJ9dzMVYnD4HTfOivZsMIguSqQg2SVttQbU5HRvi+UYE+pFETev6hcKQdJ44PzQy
sO/UOZciCKs59hwqRLwPwCxLmqd13TUO6rjCvnUSzN41ll4yi+0YBjTL5Matd2mS
ezmjzVUvQ1LnK1Keyk5YPEhnO4I9Z8e3UHcH4qEbUeEr6ILeL0V25HRgxwLOYQY6
jjOi7aI8nEFsdu65P7BqmUdQmhPfDcF1fMO2jadh5YQIJjhS5vUBYZqdiieZRkaL
wrVbK8QYuIUtPmnUJEgyd+1LJzECtr3hc2saVKZhiwH1FJR2ypBKA7HQtKHEhXfe
Nk4QGl4ZaBALVyTzavJWqIUu38mcIeL+jPhaDs4fDyzwzJTgPVocJ6bvM3iUG6kH
7zxcDGjAOPwtlrTFj0Xt8m90QLB2Nl46IcBEV4aK8CV4RrWK1bCKcVgmnrXh1cn1
hQ1qEZX+WzE9fdYHV5Ws7XYNQVCssORkpFP2wscsxfn1/eD4rYtz6W/kqAC1nWiz
dNIauovBNN/yAC4aW3Ir9A==
`protect END_PROTECTED
