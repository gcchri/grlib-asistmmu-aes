`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CvlwIhdrb4iRNIBkAqUt3c6kv04jjFKaQhuqJmHe/jZ4hFw8rcXowlwg/4fdMBE3
+Xp9hRfS1cHcerAjw+cn8OEO9YjjHAqiodela63uY0V13CDd8pei5XroiduwhU7v
OUnMOBsnNzkPKaNvzdYSVQV2I18WoS3Y6jShaIfhrDdeY5d+vDsu03Aj8x03QsrM
YAM0PNTTPgz8+8aL6nVF7TcHwUjjh7YLZDLyFxIlRP6H0ZzCZdfd8kGH5HH4GT74
qltjuV/QO5USh+xxE6UQVBty49QTNWrWQAB/lBNO82VsQGM5X0W1doQDjLTj7ILE
qfxe+gUfFgJzifgJ/g9Nu9yk7Gbk/xIpXbDCrEYuMEu5SjwyUTU0zyhKUnZNIYzA
qbMllSH9XwZHi49gyQG9bidrxmMwL+1qbhRWk3jIle+C6+uIMdExlmnf/KMSyF2z
wvmbSvARV0eJjUZCsmfBqWpgc4pdkHIU61/aQmSLwmHIQPSj6ETj840eUcj0srWP
+cHFiUgBrtggmGfKiaJW9TUruvl9GaUbppRuJrqffYU7AxgNlBYUhbfBJ3EKZYGA
a/jv9KC1/O+he85h5TaI3/BcK88syS7dbKYWEaHut7Wcvs3XtH+GUcM+KLWJWz2j
oZtLLmJOIMv7A9b19mL1x7sJ8noYeZLCgmzbjFxa7xky+LZnXhHVfxadYDIaPiBF
4jbwiJGU0yBDJa2/FEQUEnhSLZFXUvQxGgOSnORuWXYmGcIz8JOa8Reywf+TDJz+
OxetM6wUlBAPBJ63JT7O2qfMJl9N+yI0frwFdHwN3NHJBJqMnL/NcBn62UEQKR3W
SQzcU7as+e614/GWGz0qgyJq/CblRd/mFeEwjUifuGFga1n1SwP3dVAz37OMArGv
TKmpKiFDrQ2qaL66tlluDs9bM2wcaDGKcj2aU0a8Vz7iLS6Li2KCC5A1NxZbQ8X6
oCC8ivgm+AF9j8gnZ4SWPnpxXDtcgS6+qdFotFenInqRhZhg6IS7MakY4uy+6hmO
HSbjCrwfWCNtj9A9Vh3NoVC4hvfTxFRoP+xc+xYq2iok1ah8L/AeuHKpByrGFzRz
y4Ui5Q958ScM5+J1sGaOd1tLkAdUXU0igmbFaBKRG34o/kTqXDideuRssP8u7E9U
1UljTMUFwi1C7agtsEWUwQhfNf4vLCMI7RkJXJGTCc3mEFWW3g8VMzt0u0Qi4BRZ
jMrxkxGCykOCGgBNNT+Djv7jzqsXVxu21J8U5ZtRobrvoIhEVxllWAHVk1RsOGw0
dVJocw1sBNrbzNipqmd+6QsyIT+a5gTiCDQQbyRHc7pyvpFkQfxK4l/C2vFf+NyO
+wPDcjGaTPEBZA6mMzYro5G8u2DeOKsMUwVjVDZMrdJzqGoHH+kE1GtRoRpNttYq
AjF79t5AyazHcu72kXemhcc2SaOAmbWhb18fbnM+a1sRgU8WSexyqK6Dxj0Af5Fu
0/yeGCbXFgWzhoU/xNGcTPvXbFNQdeBEmhdWVXbR+m9NexrIW4Whzr6O3RKILr1l
IxcM1qYMRRzkI7KSILo8a3+bRezUPJkBwD3nuAnw2X1sfg+HKAhF3/UpUnsZBfPC
71Huoq6k+3asn/uDzeKigKh2Dhs/PD7Cj0an1Dncy5j2E3xcMs0vcOOTfNBw4Fnx
PyYtV5RY++kXt7qN1Oyzm/wLlGN7NqmPVVU4nZb6N0cB9g6PZh2fBu30UzTAHRlm
UTx5NIuvNQ/tOWS6fUoaknAfYnpUwhvBUDpO7g9VLq7ZLqEliwfSiEN94YBbq8Qd
iC7XOMRYsH88U0uq36VIiGpWRZuBNjusC7O8WHPQr5R5CnriKLo+YjESirmjM7yB
U25HqplqlaIAy6zT5govJsqUjUxXPNkuPFudhsrXmUeYUOlKWfOiIVDd8wbyoodo
c5sYbd4Sazngs146jRdmru/chLlP6/ZHSV0fBrtn74dJo/fZ65t6PQCj5EuFlA2m
d0dDV2P/qYGj7yM7J0zFp5E0FW0nRNoEtvdKiW6R85kMGBbAeUSkbBI4sX1URL9w
Ltx+cB14TMQBp/9CqOjZRVZqu2/bEIF6gUtLXgNuYLZ9ZASmEBCn0YaUU7NM8q37
AbGIDn2rNJ4XjabU6c6lhwwILBAZuEEqM7VaA1Mj4ycI4zxKWHTIN8eIkMbqfTfB
MdxAKxP1MluEyyEdSi2cx34wuhl2yHopb6WKjkdphj4ZWfdYcEPsTAKQo0hymdTz
WT2qr/8FdhCwGmGplNNOuN1GkQ/1fC767cvGi7tHNgTjl6PS7DbydbnRq/nudWnf
eO3FKdpSYfahQBmS9pyNd559an3cakEpvO41Ew3AWXbwMo1ClUGktA09T0AcQozH
gcbbNYW4Fk4kB/9fYQmaZeMHZNg1CVd3L/hMzqcSx4GRTcfIeh2SWRJtj6EMz5Bm
eYvjF6Bb0v+QHzjNBBRh70QN1mZpodG8D4+LFhfweB5vTJHMdCZXoarDnhrmGSb5
lQMqFE2830w8xzYDzRrhvkpPd50OdrNEnS9cYckjzhkTB4xvzbLM/cjsJMeywgPX
wla6umk+LA6trQqf1U2+K23OHxXOP32Ey/uQ4XsSjzIGxfq6GlrbJbW1N+LfmEO3
09KpCmX2UQHmxFZeIvGLutlSGJxFVpjcQVeqnbEJ3jpnTZZ9QLyOpSMcEwv838El
WVstyumNxw8P07iCS/37LHWCHJ5zfUovNgqS2EU124B+y7TZKESeDOQwoJDh/0Ng
QVEdKuHGPhmB/aXdMj+BsuT0ufvcKhSTRO/AXDtFyGKqYXCHUQwQ4QKEVZaTCOyN
s/ZOrw+zCU4u3GuDbEzrnS+qqTLfKANkNCsBVjm3E7IMXslGugocm8rLar56hB2I
gagJLRByacq5qondtWjE0doIIAe12XvyBOkqzyV5ec/l1fSQJD88xlBRfIUclDo/
/cjB5HYqQgrpdUFKRA/gz/i5JgadCOs1FdOSsRAaVe9VL54xwsqmQWgkL2YYu3l6
2F4DogRxc1P7UZ+HZngEmTSeM6MuohuOvTAqs62OIPBumtqaBrHDTz2UGw5OAm1m
m+nAEgX0Tashv7f/Jxd8uMV6soDZ0TTUwEC+SJvRHbIMY71paFJ72S+wariY9LUQ
WnEv86TUoLvz5aNZOEeCFdt/j/ApA0X+saP6kQHGvl+/k3DVCLUE7JWyK1n8Tg+n
li3dNAsoFn0bnWXiKabL1qaNlvce6xxDolDenmgTBNrT9VmExjxuZmNyc0nTUj82
yQnnIieK8IZOtx9ef2CSqixG886cvD/mGdWL1HzVBzKFZ4vn+92Ybtt4fAItNDxX
gKpCeZab7T9d95vTpjhGNeel+WFzjZkfeqYPXoRLHvXZ+Aq8k3SoPnYuWH8/2gJX
4cn44tm4RO9o8Qz9mAl7f/qgNPRLy2diPRJ6+qdLsMGsUDQqbCdeZkTBT391Ssuy
fTos8V5kI56yQcrIl834P2V1uwfYQ2olzG0FDDHulrKs8g6wf219JO/N9OEWYwcS
axNBPMnHVZazoNw2fOfvXA3F1OEWcLAZ7SJByxy0iDlUYHpyecwjnlj8d9yOwnXg
qmfkPuBgICbLGNS1R0QX+K0Fa/AcV41Y4U/CQfsTWLU329OUdGYfS6BSnOSa6NTp
FZ+oEnIm4F2vQblUGdsn2qW8/cpMhRHsrIDVzXqch/Irl151cprwJgODIrdlDH0A
Okbv3ZD+6g8iyzuHRseW+LeeXC7FdpFMG35t0APtcJy1kgFKtw3nkoojmpZoBlBw
uBSFvMWhy+wmNxMGYNcIRdVnkspTmTUdDBCl1YijnNpmxUKJV0DSxQU+SAz0okjR
iavqx5zrhvPnpTUewBPfG1De2ryd0yjnm/sYMD4ZYi+GEyf8aqbQMYHlpUE18rpE
VeOfX1r2ezjLnoMUcsdntV2KAOUobmECcMJrtDYByGu+g9zZuJ43klhIc31X1o9m
sa4GM5OYMat9My+V8oKTPB/CK21vYI2/uAuYXGtxVwa5c0RKsTBbncgy+V0/1LRV
FF4iOg35K2DxBjFpeQfaYxDX4aGg+5tO3S6i45/6D4ldb6hZYTBqTPrPAeZ1st01
jK0KjJ0pbgwz8d5sQtKP33XZohNQsaeu5M3qYTD2pm4ofhlVb9wBojDcHyU9gbTu
R/AZXTHFYH4dVl7mEsw2OZsdjZsGweXgJQTis4aEpO8L85m4an39bcdZoHyBMZjN
q5WH9RBW5oJxoH+B7Y407w9qIWsoM3IsutVKsYJPcCGxLditVxoScIGZK9LZpfk7
1m5GzLUTbTtl4szGcB6wL3wqpC/13ML0Knn3DSc81SfX3mXPXjEb8rhzu5hgxRTq
t/N40qhVyf+SzcpK57M2prO6Yu+nUw0fxkAz7+j66yVhxSWC5buwz7UK+JWIqFy+
5E0TJ+KlEEJRGHA/jS/HvhgX1Wpm4tuHamOG/922+mY91n0bivA78mk3vudWpVgx
OucHRAzUr0AhliXtz/U0uUTihpglMCZ/eI7PmFRzDPGPatzcUyKHcAmSG5zC0L2e
upo9IK/rsjfJSDaGBfvlbW1l2Z3w4LU1BSswMnmzVT5BVoPDRvvhHms0iI7BRSjs
sUJHcL+6V6e4AR6388h8BB58UIpfraFE6Cz0g3JcNAJVOj0ksyyNfwZHKh43puFm
31Bqf44JH1xXtb1uVY4dL02YMhopnBbDB73uCC1p8CvL77AAtjYYwPLDFoa12BP6
oRtRJbvWL/I5CthsqfsK3t1KnEpE+g/YqLx7NVH5EI2w8M2FOZXnJKTlOfmm3HT8
eSt1wzTGmIQweXYoH9F8NpNt6yW2TFIJAi857TM8XzcUR9INvLIErnaImjFdGY+6
uzSTg77yGlzPTCsbz4y4hg6w3UJdfvqGXF14K+F2Uf25ORvYGjV2XpmBbcff24l0
076GxODjWQQy4RqoFHPwwAPE/YZiFgu4ai9DJqZ0RCOiV7//wZDSfjDidR+GTRzx
ieyiSHbL8EbfT7wjYmQyL/gh00mEseR4M08YJGS7ezgzhTh6eS+EwnBVJXoK6wIc
0aDSW2vXcQCyKi50DfrZRkNi/Zcr2xbZ/tkQCONISVicdRcz9ELpbqAYmPP8zPqB
aVJZlVSjoNCi5ifOhe3o5m8dlxdK81+KxLu483eEc7icID9XWUettCo3yC9B0Bgr
Jeyn/f0kbzFCjyKGzqKekOwJFla50idRS3cVioNLuEqvvZi2vlQF95jIHJJLovqI
tPvs/eL1gVgPYBVKEWLGZ3MoYTEyiVSMMt+1KYetA1FmHn+c9fo9C/JZz8+znX/a
9RYuru8a/qMQpFQ3pbuFPkby6z0s1dg94jmFiXK2AGwIG6RMG6JG8Wzxhv56lp1P
JXVnksFZxZFRiObkRpTAlMIOPo6d538U+XY2mefE5UD+UKO7LWQyl7SUUwJTu/74
AqIw2f+DcHH3S4r7cDLnZvERw4X2w6nGKnK9iwjHXPshFOuoa/FfW6LspZcRs2ID
AS0Li6M2iKOD66Oy+CVlSEgAPBtVfnZvzbGWx3bNCEWoXPigW03zq0lM4PVaZtTY
yQyY3GnxCu6HXLMPjKs846bOMgQzCzYyfbEtgxr4hQ9Ws9Q8+R942TdplrUxtzko
p87Pi11JKqXHRo2dslzWkg7/z+bhIkxcw0x6RFwYAFQ=
`protect END_PROTECTED
