`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q742lqJtMV6YUuFeeZ0LYQqBsOG/JPEi9pwHHn4bxY2cCXtOl09eRCRQCQONu5QA
UmyfzIlWJsUk4M/TI6Szz2mmifmDLQ3l4ntKWeYSiGmecpk0z8zjP78QVBC1KCWN
/4qu6Sv8sJ9f14SdOK0YuYVPce71N6a+ifXLX+lUOvfC8z8kw6EFF0ygzwv1ym/+
MrNkl90zSJB0vQKB7eQv4FXDlhdkRVJOCc0FSPyZRyspzDlMSSUPo6TIBvgycS0b
pwoFQfwRn+bHCLqrhp0n7QpdAFzw1jtiY4x/8IfPSRVXj6XP/hrd4sYI0DqGm1ga
B3pABxu9ngRPXDcGA+5sAGfNx0eHihnHp5CzYmOAGJm5yNcUZ79EfdPyJMQo4o83
KuWbPb4IZidFz188Xy49Og==
`protect END_PROTECTED
