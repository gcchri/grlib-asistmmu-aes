`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KheMPt4KE64wNBSChkRxheMLccM7hxoaXkxRup/8fcHRsaJAALI2rRmqgfqvgMRV
rS81IIBuD96GyTVLcEmBCoESyUXp45hbC/Zah6KzYJIlRxr539PyvjgM2xipbv/k
unPGhk4Aqx3ElKxZxS990T3IvFlYBDO98Wf4uqmSL34QES6rOAE8dIQXxKNb44hr
k5+Uj8hY43IRpbNUbWZj484fi3WGjGIa1zGyG+PlYNZFvWfs8UuKPWds+CQg9upt
llHyW8BxCmdAsU9xkxTB9446K1WjAmnE78+Xis1AXSlBlsY3D029MKT/sskFaWCW
wo3t0PzMclNpyS/rz2hrB9S5SWMNGPX0uBO86+Sx/uxPgRlOwWGQUDlObmXoC0IY
EE3P2PyA0SKML2XuRbbzzw==
`protect END_PROTECTED
