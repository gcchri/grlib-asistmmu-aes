`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BHwfVYxBYNsUttB2UEkhtNqNXDiZzvZX4OaYMtBNPyM7hCJciLaeUiah+1QGuu5t
zsIiDKVG6RoMpNp/qI+6CR/t3/EU/SaDmQplbPzKzHG3gFPmSP4Staxvc/aA2BR9
9PSqsQu6Y8SEM61d0w5BHUvHkgre+MYMiZv3V4hPktNK7ZtEjzg6ACZjL87+o46M
1JMgLAKPj76LbC6DjW2EjhefNp88Y6k7/r2lPyLdBH7M9odA4z6nSEbRaMCReUUP
TbWrcQ1mE6es36A0NJmZSCfPzluq5wWXqm7srSKHcOUb58GI8wzR1rPf+oYyJdgI
XASBy1ntTLqcMXyWts3pNrNYzxntddt4D/0hVwwsaXHqpqdbhi9Aj/sBOHDd6KTI
`protect END_PROTECTED
