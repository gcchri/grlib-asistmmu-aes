`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VeXARlXtRPsPLfdzfE19XgjN6UjKyR3Ks8KXma4aZrpwDOmor49CJ/LAftmByQnV
ErlsIhEGk2zs4aEQq7/E/SUfruVKYOmIEvfa0gIy6qql9FCSeyColp5oMooR69BM
MS13yVBY7nCAZc89WGZYyYVIlxJlF1BkN6rqBzvHp/iY3WwxkQAamniaQH2eWTaL
/8iSy6CsHB5AznXDFGL03XVDgxhScJ4ktaRlWgM708N8psQEV7ovY1JV5IcqngsE
h+Fvbuf+osjgb3wl0/lWyPxIPb3ajKcqrvJafo4L9wKBurw+xzqgEFdoLbW458Bp
WkGbuAUeNrYmPrOJpPvymjzYyv7QNmjInB6oTxrev+jiEiZwUHusb3O7bufcsuQA
Cl14k/kkwmIM0ZUYb8YQxVmXR07eA4lFnfdaemA5tFrAlaKCP8EvvOxnTHssaNlL
WAHD859EJcfc1ewps/I48NwovkJ/oChE7NjXa+s9bPJBowklSJU6F95Z4WXdZgwl
czgbwLabDtJpoTlFVyZ43MxJbH79m4zZJ9rgONFCz1HjKOGm9tYgyFNnKgHiBHz3
gY1a5sA3fGlmlTykkju7Ev8OTR4Q0qEvd0CZxeu0/gyDZRMI+AyuUUfRzapSTiE1
`protect END_PROTECTED
