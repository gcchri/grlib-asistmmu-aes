`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1xp4BqQncgfYRM+fMnnkaEo6iZVXnYYoxItZ2UGLmgTqXI6TLjZNrugMBk7CyStS
MttAEb9JQNpHxcrqJaF4yuxsflwm2jy4pZEYUZ3oOidQ9ZKZNFa+1apU3RWFJG9i
pxU7jkeJoI1jBq4Ffnf/HneFt+vkAo9yaVXWbTZyjG6nXB8WMil3GK6VWT4uLU2E
YRlxtOZQYfH/6BqS6/LVUcDDFDo/ag2pXayR+LRXUH/8ZW3Cgs+daOjou1Z3gCd9
Rzo6QdjyiKbM700Sqgx1jVRLNJelRuqqKsACtaRyfFGvMfj7WIOXrxZhRurBE6es
7gj0bdpL2V1a5CM4FBp8BGt4bJ5EMyN6ASI/CAaLp+7gwXyjifzWyV3jsfJ8c7LD
hFihV94W1DxPDFS43I6tXhe2zrFFpz88MAOGHMSsuQS7iComm6nfPyO3ptdztlpw
7B2mS+Vhz11uU0WaqVkJv2SaxiiVfhPjbO9PKMJeWvK0fg44KDE+MnL0OEInNDWm
ERIAXGDSGE8+wjZAPxRsBkPMblXu7JwEkb5ov10GZRJ5vwodVYEIePQ8iGTzXjHl
XwoxzqInQPt/O9i0CMQgzw==
`protect END_PROTECTED
