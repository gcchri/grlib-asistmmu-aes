`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZPQAULwfF3EnTabySo8i4s2seGjlDKMiGu0ruyj1sfl6YDuBRLQIm2AogwKuOthe
u5d0M8tDYuiL0gWN8ukSxfnDETwop69sn1vcfHJ7O2XuUvVAgSfjDFt9D8Lfi7Nu
crt0sIVHwln6A9RYhJ3ROKQOIWfJ+PUcHyav9HRF81wL6ODGM5rzbw4Q245VqTIH
Z3UcUSYaApmNDxxyZpunW3qDNOqz0wqixrAo4fhH6euGsXnUkdftjMVzt1W5ajZO
/DApFwwxNCypf3uHtWMpEWkS0yEimMKRXNWXnfmJQzJZzyC7y/cfDyL76xrfmuno
+p1T6cfJYdBk+LBRoqTBz3Q55D4E3S9OCZFIMdUU3oxs+HG5ZTlOchmyT7VUv5Tt
zckfai9slIRd9+L3OJ9ksS39lYA7fdmM5qgB8INcxHEPvY6mWvqcrk5Tv+/gYuBU
`protect END_PROTECTED
