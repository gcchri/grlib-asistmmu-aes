`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3R72mfplKoqRqGDBU/SORGD5KYGunUzZOuJ35mcFRqJxGQPL2+re3GL8ir2iFcnw
rBuZT8mu6IztRQd3SrEKoA2QZTsUaJ1vSDGQBNl/GPNShmU361Xk8MTPjVMctAvd
mofWT6OtaN92O4wX7pnk7PkY4qDvncb0lK72M3zImmFcmhk7qVl7YUrB8dCB6Dk3
iZP/LOymsb7wFmcFHb5MJ893i0RgSoSNLomZ/D8SlWkPPz5Fw7Auzell9VQ7z2Iw
0JTwXpDlpJtXxkM7GZrzTUyv4NNqPKDvsQxaA3Xe2Jof0EEyQgi+ty7NGjedBt3n
kHWcQKIZcRrPht+CDkRR+9Ff7NLdQetYWITomHAQMQxeOgkbJm5J73W8GZPOVOWF
9XG389o8qFmm500KPAXqiuF5UDvsiPvPlVp8XP2pkik6RgGUUAN1tFyExgsOK34+
3vNYPuPhNvU43P/ivIT25NhPZPKXWqjAECQCri8p2EnB8wwy07G2QS3VILBoOnHf
i83VOGfcuSJJzH4q97m8Iyaj3Vfm1ZipkHKKKMMRvGnqk+XsH/cNdrjShCSFZsWc
sVHAXuRmiNqAk+VMgaZp7p39xgloZqzRslEV24n/i9tJpXNJxyFJ06sAD5+Bcq3X
0C6BZo3nyXXl+ZxJIIrI7g==
`protect END_PROTECTED
