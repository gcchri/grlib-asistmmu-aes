`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jWDpypaVFgR4sAgFRxDew7FIkFTOfWsvSGoIWypcZ1vmUPVTh9Yolp6dn/Yf+gjH
JFNvt48BcRCxKAj7QntfJKfMQmRVl4Q26wtsYr3G1+DuV72hJeo69TArvpAyBWH+
nIq+49DEPXfRhn3mTdi/9HaAc4vuyMIP2CNSnJxO7zji2BkrbZ5b5ncromP2Vdt6
i6/NwTReZWNtQUUOwuRepRkapaL/DDjdk5ZhrB1QrpMlHzECmseG0Dw2YS4gcAGH
T4xXFwc5fMtU/mq2dkCWcw+sfa0Pjv8KyaOPrcJuEoKv7GKfoyoUjgYMhE13H7PC
AAlxKfc//OIDucrd2Ja9oQQUixW04cUXn8G+DawrKcvOGhcXMBoNmQ0xkWArcdyl
h/Ya4jS1cYB6VhbAcMltSwBU+qjW6szC33R94FM3lQmUo6xmBTXURsxsqUAg6eC6
UOlSy1XeoTKBA+QF62+NTqQEM3tPzMe1noChyG48eUEdQMk+D/eJn1RwVvZFJoyY
ZS0dreerSxwrFtvbyxKCUQNm/DkFoQy1tzd8xf4K2fJ0wigtw0hyNPxDwpUuw/Fm
F6zH8boJEMcgdluXjARus6f/UDc5ljMrKfqbVpT7G/LC67QX0fxNa+JjglW0XWNq
8BZlK8QzUlr/4oAdcJnG/IFXcQ2muMSkxJw8g5LzkZAXxF5cwH3Kfsf3/HscMAYT
LvgOVvSuW1Vn1AqUGuo0WoRqwEFcmZjJSJzunb1jpJWAJ5/XpDeRt2XKbEpSBrDY
rFZUTGirM2QG3JIBOFc0myNPCD/Bc+M9RZ+hSAFvERY=
`protect END_PROTECTED
