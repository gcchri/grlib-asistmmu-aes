`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q0rjhbEODOFIDoWYZLgMXbQ2MmRLNjAgCPpV5FQAUN4nskU6ugMAx8noOJCXLgHA
nIWylT6517PdvsRZwHE/R7BWi4syJc4ucOioD19TJbU2dgle1+jjrB022duSuCCg
GD6m6MP7AWUn9ahz7XAEZBfKmqbaRGoIIrBVYwKER8pN3VInQs8T94s0BDmcLaqT
KflNMzs0j50wtZZSEihDqbLW5I47pTM2Ysts5YDEgwlBOQNsj4f9Jt6vrw0FQA+5
mSHeUlsYBRr+X/6AlAZce2+sDG84YkSTx5Datuadb5a9s72hLT/CdLwMy5YX4JO5
Z4myzdS8b/GeDBO27ZltiTQWybdj5J7FBg8skUHRZe10Srl4EEJH9PidL2OHQvud
AQmrR3zvXDhkw+W8lM5tYelBv/5dpHJSLKCmC/6/Pg0oxiLRbxYWQA7NHXvi/k6N
FvoRfm6JdfvauqQVFnR/qHNOLPfkqzLSDMtghwMj8jYx+6E1RceePPe3L7nOnTX0
Flekw9LTo2jSHtaVIqFaQL5FNijeAxeDypp6KWh5NMC7UBcy9oMEwSvsHmj4tpsx
/+Axas2O7zeXB64VWJdZ/HfwDpxDkqVfHXEK0Kw87Av8LS0rSArgNjZco/VPxKiP
kUfjs5D5zvm+0GYv7dbsaD06NJudNEjcrO/j1kqpuB6CbiO3hFA6FyYNdbY26+as
RZAKIDDcv/dUakHvjVi+Ykv5yYYL5BsC5AvaIXqbSN7Zm6Fe54RfJ754XtJV2yLN
D44HVeLV8D6wqL4S2yh0idsEezqVn0ZmMSuRbSwf/uyCGUzPc+w+wybCtwYtWla8
r/ieIOXHtJi6VthPP1FcE83GZFwIJADKChpW1nCMtJQDKMS5GeqfjJL8hEWpqT3J
LG+XtvaN2NLs2ts5rwUE8BKKWuvWw8by+mV+9bGaiy3JmK0KcTvJLYVjBnNSUuL3
JgFfI6KchJe6n/OitXOA5no7v658knXQtMp8EMX1cmcj4gjJ5kZhushBt7d4CdyN
wRZABltkDSXtCRGYqV5r4Q7zrdu25JZEl9+yCguhmPDFjxE+ClHvLjr+LgJB8NPg
7Tz+is9SNDx+didm4bGSmXd++zLnK5MI5OuaKrw8cQZzhgK5o8r4wFFp30gPOVgc
9hZkP7vtYNdoFAZO0xTRi0gVaYd5O25Zt6M654hPAIlciZE+NVXANsDrbyOXandO
fMR0Rfo5GEDIPvHeh2wXKBaXuzs42KzmhYxMlOVHQGIToJOc0MoT28c3Vwg+/Pgj
OTbRZzxFAwJH/aXDKEJP512V5QY06GDOQgqYqaEm1itP2WoggfFEMbgaGsQxuQC2
/JE2wM+tCjINLEdODUBJDFTk71Jsz/1p7BNebN55UFtqT7/RWw+fIxrBt4e4qgUp
yktC65E0Ux/60RtQmobDKMCcnbSuEzrQQ66hZi+LhddfHRbTmdRn/G//VQtq0SBA
nDGxhM6u4PEOAF0oZrQ9WjbRsfxXIDJg16bcjQvuxY+vwBQgNkOI1v41+T5K9TUi
SAgXCXNjQPDoFCR3zZ1XS/ifVSgEUnQLYudOkE5f8G7mZwPlKVqzgVEeOws8sAU8
NeKR3VCi/hVwFdmdeYeUmGHlkU5rGcZ438DrI9bXSy/RLU0um4zdhybw2GX6nta6
w+8OL63bkEebZ9Z2Kc1s7CFU+6IXNbf6pCBL1USV6f3Nah2aOoYMTPhIphhdCkuN
tOKGuruHgbYp5YndDVgtmXWNmwhpGFHx/gDqu0Woqe1hUeWmWL4EXoYx4NGyBEI5
WEn8xmd7UkUWRKZD3+1iF+A4v+EclfWjkJFpHRVABMvXAaEasC0bXRfPnjDzHfRM
/uOWHaeoEcBmyzjNzx6KvNVnwztNZ20jVLO/vvu7ls0gXnRoPw/avdmzvzFX8GUp
JFuwyrvjSOZkyptyZ2432oYO8tv4bebRK1LsBhgeMG/W60IgXxCAsAD9GPxs6XFL
ZRLA6W0pyVvSV2pmTjWMaVjwHB5YULRUYTzFA6A5joBoEoiMG3KyUe9WbmuFaRqa
niCR1IW77rLZl9FEgg5wQokYWqvXmXZFnrnKUjXiRipY/VbOmyiO8+tjOgomVYNz
FkugitpXFQG0Rb77STsQ+t1bAH5TV8+2zUM/rZHr0vSTUNrXV2icFX0AmFkry9wF
YREVyVIHjRu3kViX9ZPq7iYW3aWYfUKGS7jQJUnNsR0VH165httWEFK43W1/Ned1
h0/LZaIxRZLd4GkC+fpNTI+UtyCBPS2pVt9yk3+wmxWF63087qub1JezKVVCSF27
BOCP3YOCFRpUMF4ERR74AW4N78i55sFRGNy5iiw9/QTqT+NxfcsVfdsswSBwapQK
ea/wctGhn/J1h7Z5sEpHp5fK8QOA1b3aFRJ0TGMeYYYXR1l8K33aGuDSQlHsMsPd
LM1jh/11Bgm2p0pVqFEjm32ULctXkKvayLi2KQTOlkh5refkP6jcah7/KevY7/LS
Ox2n7dIS0ahpr2mnyJfGrF4xzGJRejcCrgVl4t7X31NtYAnTDXd6XPWft2hyJBu5
U/GZKQnxQG7tZMC+WtV3BvO6vSKF9/qDZRzVSmUqZlJuZ476xcnRyLFQhzbHCoUH
VBA3A1dnuOmsJ+IEyO6oDh0pFhYhPoIwA5JGZwrgh9d98J2FzJCdUngnHEwyjhWs
l3qgQEkG7yC2koSham7ek9LtpLi3EC6t44Kdbfr/cji8b9l17AZjGfoupVwkgxvV
1fQKhSPSMqYcqFUl3z59BiKjEWt7HEVTmfkM5Bw0dxOSX8XA8fQHhXf5cgb9Mg8c
sS6faq4G+fnH9HQaE6Pq7m9iOvMlcROauVgPm7sqlmCj4LuflTAnWyTuLysXb9kI
NSTTejI4rU7AEWhFU664pinxtS2NSp4vB2TXH/FRaPxNSJD691tVh4w6bER68yuk
1ALuA/12v2APWsSUnBigkxhseilo4lAjZSJgv47ynTQU+AoJPna81g1B8exgyAak
QkaOVXGyOp/UySyYZkn6gICc2l6EevEsoqgbm1Oy5belUiwYm4DY9Eh8S21qnDI3
rpcmnfUO2M0e9FccWWtkoDruKv2wD4F22n1g1SSD9TKUT0QTNd0LjvCK8WJ+Ofk0
JWgeZJ47unkVSXcIkxCjL8J3SPXveCg4nDQMjvYM+lWNgM2Vbc3vLGsqF2Jz2dpt
ReEuxwKobkB4ozEQhLPqDfd8VsHG8HkLflvmE5TnhAh/3NMVg+KInbUFE1KJUZo0
A5Vip+YUy5aCc8pRH6spnSqxDxKfTE4KC6iXG8qdfiEr6lp/bkZ8rnrIcmKoSDYB
CUWE8DwXWekKdyhFiGrfojM/qLDjZ1rRa8qSnXFbdCSBR6Q0pblB3GavgGTuk/6P
nTxzic6oWgLxujGadIGZ74l/lUSm2bXTVs9odsYaHuZq+2L485+jUWayJGhPRdwL
LYHh83yN63BiKhAD6LbbZZDMDDWFmfPShpANOr2OkQOZ0eAYDjNJYbuJjdSxa4u2
cH3gkhvdIavdgClUjysEaJahID67lB+AQh4h1923Q1l3ze1iTpMgBj5tdhTaP+Dw
ZDBe0ADoOwvzRCmFNgcq/XTmpBnvVKVEzjG/crJfHnbNDYOOXDxAc5yoPJxn/gfo
3sw3FL2KAk+8L4FuVp9C7VoSyIXQbUBuhOi9NPdqv7cjnCYHbrH3mLlaZh4tQK+v
UH7s5QuaS+1yPxE0tKOUoyh6oq/vD3tff6h3ywgPeEGIa6sdkH1rogi4RR+TPwAK
3k+Z+GoP/Giw7zGur4zI9SFG9DBJeOJZ7pprdPI2reQTgklX7YGKEaCvsaV07ezk
zAKe8vCaL4E3dr0UQ72ZJr+r8m5BUdvDOo2JchAU8cdWnebR9YDqKe1YjVoQ0VgM
emT1m+60YMp8RgnaeN4UbiKNOpHLVkqesH4smWoS4CCVtqk8DIRHbBqurmbAxccO
Db3W3P3e1MpcNu+VFJHlt1eeU0nytUF1wadBo7Iov60MlD6fKVMaLot7TJAZQ8D9
LR70u56Z1LT2CikJT9h+u1Hiew6UZYpIMkBrLKeiC8t+q0iOYTznafy3IgZQUK4z
4T7Hc+a9TUVSjszEK+s3PRnsBm2jvk3RpYS2aE/pQ8Vb7/JOSF667woQLX4PXs+b
c+3vdjRRuVe28x7JiT1qAoOM7XytU4ImNModdpZ8ITf41W4eaKyAQ005+A2f2d4y
m6QPbYf04Zcf52lAyYv9QptRMxhsQOBwg2tgVLYzqFk6FlSOoXY0/uKzdNypnl3R
FVbH+znOBC+5A7UW3XrE65PcZCKrmw84N1TmunFAHLoU9g/16kqYh41Uzm2ZKypT
jYrU8rt4zb9vAyvxx87DjvIs6GifuvsZe0MO9ePHiQMwzNG/lBN2e7gPFhi6cR6y
zV58Jkz6gr27CTxWzQpN5UQ22u+8nYR2izlha1Nc26gWlA65DwURQqzfndFcfzZJ
rvxrwGSODfh24phAHQGLwCMe7M9RQ5/topxcTiI2hIgo8libt8D3DHZxmeZGD7lF
Q1PDS0Fb9Px3by9T7IB/YKfY1k010ywQqvWGVi3OzZyzM2WVezHkYLVtiU4bGHjk
2zpz61t/Q197SVUU/WYG6xx7jWaXLSM0X3q0YA05HqS6WV/2yMY8ArL0wa04E+mR
fdPoaI7tTEVQtaai2NKv/7cPoEn/iog4YuMRfkMS7n8FE4ScTXiHWAvJd+vzHLRq
R/k8cEYNlZNMzDFoAf1PNKA/xXzc/gccm/te8fVeFLXYitWeZvUE4AzGiSWEEdTi
KwWLrhf2jDilvFx33kDewfknYv6xmgBKWoow6VrigHw1ZD/1SBf+zWxXZ+x994Gi
CwnhoMtXYna0hRQhCIQ/aGuVnm9qGm2BeNZBX1iaFSQcoiqUNP50O/MTiV5RBbDl
LQFGvmHVWOS3nQ4/fyANnaLel2r/VgpaMZ6Xc10nkFgJX83RV8l8XpyKCJSxL9QC
/HVtZ36tLDy48+fq8fzDD4Lcgzbt3Wd5lcUcPi7c7uFgPSyXPoP1Pll28Rw+EfTo
Xe0UHHqJlq0dSKP3ch+vwiy8AaqvPIeHOttC+P1T/MlZAKI/V/OmtubX2KbX3Gxm
WL0KfbkfYkzjwBGFIObt5/26zDUWKbXGNK6fzXYzxUjgp/9QSfSxU6hNLzu/dSYI
OBGiN0F4GDKVBQf5o6mbyHUhpXTEe7azqexYxGcReBSdbOvXFikLHqXYcuEwj3IS
raT91HQ5OXKxm10d3ZPr4lf/t1n6AmcuXZbI0jvxXeGzWw1pny58gdaJYdd9hSFm
7sP3BBRQmKQVDNI9oLH2UNGgyl3XywBF/LEImYkA6Yv4B4YqJSbBchWrC2vy2ExD
KrHmCLoNT640GRmwL0QIVZYu6xMqQe6KtrE9seytJY2N62/3hARlGxQd7pUyj3Vu
CdIbtA1aSygWaHixEnea53iJVSP1ihQ6F8TeXbnH9Fi/0prz1TAVNG6uCBGOjBpF
9t1oz0nq5W/tdugmuyWxmqvDQkmIQ7Sw9wA+DLtFUNhjN70CMR6X2GEwwVOCYlrS
nkwqah8TmiK+H9Mjb6koe9TL3A8ps6UYldjSoUsQ8pWLWrCdUtKM9mogcl6KOfO1
VaAeriBv3DSbtkZPLAUdLxAbTu2e+uaryE1IkchgrqPbgh0lf31WzDqmTh3HKc7U
uQHJqGPJSxFHjiZiR4QAnQSmvqZxQMPFhEKSAzqKrjycSzebgAcpOI7ASV3xnMB6
hUOBttupCE3w+apBpL11qCqzKhC36HMZ1qHyi043kaB0PFX0VtCqOmppHC8bI8iu
r6v7kNKmp5WZVKBLwEi/eIn7tstezwSD7KYe1Lo9tXmn3kA2wmGjgzXYOHYE2Tn7
wJbpWr+8z24qPVGl0r7ZCMr4U85uN6Oj/SgI/q6pyOv0VkoYH0xI//v8WS+dmDij
eo5aoI9MWVgtggLqSzFDD/VMrlmmvI/4SNr0yeWYw5JH2Acq6JxOTeKNlSYKlSBf
k89PG+Z1st5U393WjBJ6YawVNIFSkw27x3I9pIG+DYcAi/8Bdy2MusI30qBDK47j
sJqhSg4CsaLCApl++f31Og16XtRq3oAHCoCXpcrfefs6WVXkM5c5iWDwxbqp3lyH
HC8ES4jCpJgr+11V4zOvC5tSSCxpiZi2kpDehd+XofAuYk236zVvY8NJjA0xyO9D
ajcCW/ZYAR2kKWupF7YB+2IRPZVeyY+0vaNFmWKQ1dKvlJDtjbIGW0+Uwq+PhN/H
Mr7kIdAl52poE3KzlshXFZGo8UACMEK9LL2/Atf8E6H0BnejCtPzYzwvoiwQKJfg
TByay4GzJWy/NMONI9RVYnTM6s4dBPXqyfvsxXpo3wimu2l4Cj0oTnhTUJM83icf
XaX/OVmofqFoEANb9TzYHF8CYk6/xA68jmOdEU/T3KwgdEaVi6mRk5qePvv8M63z
dONVVVcy6+OtqWdL1p2aKALUUhuBF8iq6hSXlCuS/04QZwweu7j87XakoMENixvX
HkwOgxV+46YW77TN7rcYHTN3CYIwnyh3XuLqFd3EW86u4bp3+khYE8K1BZA4pko2
uJK6rNeAvacn2QsnwDH6ljZXg2tGZluLDp1rGgjKOcjpoge9WAS0SmMhO1B+Th7W
Crx0YOU3nKyOrKbP5UxRFC5yoz/jkwlO0W8UKizSqqisSnYlSiYlmzugTlZvd+ln
NAk/LDcxmqM4jlbGCTMuZOdWaVS+HemvHwXv5S2fKqggjhF4B/MNz33Ib4pPe56w
wUzj5R0L9ITrbkGTG5qMVPrkwcWxJA3JoOL2sRe7EqSm/lcjMlKmR2v+0zcbAk7D
9IXn+MH7VjlvrogEAQX4kJ/LV7Ztejr63NIzSEOiUHD5N/awvYXlv/2rPcEb6r7b
ymGXGh9UioniXKNbhpWHCKMvm+wvBj+2wqNQFnyAq1QTZa+VaT4sZXfCIdh7miLu
OIJHqHDCnit4Ta06xKhToCzG5GoZItCuOki+SGpwb3JqBIHa6HEKtqKqYMAcMK6O
/S5rmDtLw9ZU0W5hV4YwUaSS+SfeyvQr/D3akVdn9XDNsR2uLgCXOzP8tVtAuqgn
cRGhOnAuVFKmacYLqG+qQGrigd59JpbNrgi2i37NNfB1ja7IU+Iq2IIiMsPoh668
ZHaFdpYCUZ0og5orqmmmhzmBQHLlPT9I5BEcF0RTqQZXQK7okn1hlDhdCUuAkjd2
RL6QY27SjWUo+0jJz2cyqF9pjFNTYagpz1ajxa6d7nRN9FaIVcHJuPzOlPZTKEU3
Ki/9lWA8EpY2391PL1vvDZDNl4UqKIAoOMlCHb33/ygeuWk+9xNKU+ehs6n9ciHq
WnPuDMCawtiCtWUzwYRhU6RIw9xL3lgP9blrBOuOvl32RonVwt17UrO0A+plt76y
HYVO5w3XQGqqnBWjh4x1KH0bc+NVMV62gmafATHjoKh+hjdyuuzBME45+l0zTvmj
IfcMar41Lem+5tzufTw48Y54zLi+Ssa9V3vXa+d22hnrPlygaqn+WEeQluwQ0GEd
RZY+ysMMvUBOXmbdVpjxV5wLdJaqbcd+b8AppH+MnytPnEUk8sISh9N/RI6scsig
/vO/WQEyrh0s04YuytDiYsKKNJPVOpVAPJGLPqzh1rPWgEkg+rBPvPHsQ6bbqcr1
zdwM9SUoWakVDFVFO8f2y6ZQnJGSPH2Im08QoTvnRHuJ3H16EyWHCvFdl3Ma5UCy
fP+zgA9xsnVUvTfITfhql7XW9GPYvyktOHBuy/p8xPomKNRs7UO5i0rCTq1mZKHc
UIW0aMZdK1Ml0DOyIKh2sEthPtEBNR49DG5QAt1q1ODBg8KNFO/0RQ568FoZOJbo
3QaUqbS6gFbQzstg0wrFzYPpm4Q8WHEAEMwG/wt87WSvEZjPy6MfyLiX28JlZbVF
fNjssbQXGFSEHZ8MwLXCCyabTwVhW5vLsfMfqvtx2J6/KGpHjFp08OPV7Hn1PiTw
pzY4WSQi4v+Kv6rgkcENkHdkUwcoJxmIVv5ZrdUPeXDlh++lYJ25la1ySORp/6mC
3Y8Q0ptdhdZ5hfYvYAEw89q17ANabqnVFnfzoXoS4RKcgQOI6BCJPtMV833uxvRB
LU1kr8by2PqMCumrKqwV5hkarvpPhr4Bs3Y8WxT6OOXM1Ff+wxRoDhzpgJiq8FdF
ER9pnHNOc8ju8WD3nYTgL5A5ZHoq03Ae2UCWEvSjAQpSz3bxsRAh3gjXfKHdsVoq
Pg7G5QRO6QqDU2nwzIREFBkrThMO4eHr2lOtWK0jSVqRPLHgM+B7lB1nZYCQZdDp
vIETAL1/g7Vtk63OKPtFSTEzCkvUU8IdtDiVqcyhJk8c/0six86fh2mkCiq/Ii0H
88n33QDZS567I0fT+4H1/MUnN1t2NiG5alh2/XhjZdBooH3agi61j5IkXjnSoC+R
uEbljRBFYe1s2K4sXLhrcphI/y6PEv7Ffsw7uyCJABZW3oNfwTYaJw7pCA0Xo2Nv
pJsvJo/0jJEI5qpMda6q/ejAwc+M+wvy8GeXhElBhlORhnOVkxbU1wDHRTNKHLKS
Y85lmZwfjt20f5bIyIIJ1Xo/e3ZauV0BFGf+/VaAUu1acbeh8qDwj1uzJ4C/vfUW
Ur0I9Xd7FnJ3lyzSnNQ16CDGCFDV3x2QLt9hXFoC7up5zY3NSfT2/5j51emIa3Nu
QFGWY2h52C8TXW2mNgnUGOvJKAd1hGbPUIdcjpU9mV4bmEKoKHg6Hf3dvGHNh0CP
Fjgij5jCIcg2+0FjMH/Lzqf2Nd5L8nvDaibQXG6C3ppmDqCSZ26ECJmP7pNFej2t
j1eUBrNBVwQXlZS50R9WOWMaNBqd0xZX1nz+TfozP5KQ7YdDqFVSF8F9zWkKnYOm
Kyn7/eIUX+7NK+/YMw7XNZNyS3JVnARKEQ9Rj+9tvTtEMysuYM0zDo15oQfkCSiE
X1rhC2bbcV0OaoNkTJnDiFJI9vG4OspYSvBAQh5hGWUBhRBFGp6RwTWUvf9G7kJ6
zIKMc4m7M67uwdpmCGJ7Pm9jtQD4u04kppbX6d8Jp4p8SPjPXxfqWYYGsDNaDoU9
/u3XXBFGHqtho6wcwqu5jar7uipEemTSQj1d5KEtBh6gLIxmW6CmVmOApYVKIFFZ
npMgb5ImF8KyhRBrGMrNwL2CAdjLmAjc3CzEkQ2PP8ttCuVkXT+AZIwLGUshw4MP
0frQX+UJ0jKLjoVYlk25/yjDbHQYZJhHhojWaRA09sqrDGbtBZPLH3Xi6uTBpbSD
O+Wpeqob2pc0e7mqE2QBIdeXbrj+Cnr4LG1a4bmNeuYWB075gb6uWgKLFoeVkv4n
Dx4lXYCP5M9XmYtxZpSF/3kNCdwwmTt4fGVr+g1+MobAQtnuuAu4bDhDBp+hQ2ep
aAh/UKNCsI4u2kFrHHzxo/bdyEQj38gxrK+HDhPwTV+V9atiw4nomnI1kXwumFoE
KWj8xKlwb7ywmH3a9p4YpDZXeXdpNa43t8eM3k3QPggKDJnXEQuBsASrlqgFdM28
c2kv04HtBCGfGf9Nh1NkSmfddUUxNeUWh81Ri9gkJRxQoCwgC+NsupW+Jlyr8jqH
N/kRAswaNnvUAj/yDrVdRRHtVPQ1UiNBSF56PXVeiDuqX5Kqx82utSFGG6bYHzJB
TkI6YvjTKuFf5UiozWNFpz1CHB2JCRZCmDZjreb2SgMLEu510RFLC/cxxuuNpC/U
imY+7szVmYrB1GQmxCJ2O0rgIsFEFxRq6ge5LE4HK8aAsU0wiLhijwHnHhzUBScH
8JKxuyNceDYwiQPiTmBCzJZ0m8/61peujmHnEWDT+in/Y/KICSqWQ+Tg4pKe0kzF
97MBtc4NHwn+B/FTcWOZTKxsaB8CMjJZ5n5HxTy/Kg6zQmfnFGhYM5FLi340XBUj
EvoGIisF0EVYnI1ocf8bYP/2+0Yr1oGJxF7XXcGbtiHCCMVjFEur7BAW4VGho68L
fOHi1Dnu2qdqMPXSVq1qQunyJoWT03MgkBYWoUJU59gnJYD2mzE6R2G/yDqbsc/V
6qNfRkbged4rVoUNmoDb72QA/2aABHL7nxK3BJz5SlVc3wlqV179zddxxYnsdmn3
z6uk7qcuSxSbbk6rS+h/FYZSuF7eK6hv8uzXZU01Oj2tBFoqq0YLRG1gENmTUbva
QVJKsjzUN2TAOjiPfh291qZizgvNe92CSBxkcaZBnRJsCTp4UDjlJeq8FmkX9vgv
xkK5w8UkLp7LoRl8Jp8TC37BTdBZABhYz+m+2Byuez3Ev1qzFMW1fJ7dQDewP1+O
yqlnzBOIhovU/BNJSAnzpgWVgcwi1/P0RenFZ6B3K6W5O+/hzfWsC92tghZX5Zua
r1e9yUQYqgiZlovDrHKd8TJKuZv4EIOQDN0S1fLjfEr6SglB8+1Sp571dSyhy8nk
kx9k+k0vC4znNzE9A7rfQpDnxW3Sn47aYmo1fyQ2ffHiTx3NvBDdRnK1qzw5J4b+
nHIxIzfY29Pjg1M38UBaXmsnb6FgUYOmUQDygpmj5M24vvfNLFhWOTcMVMIL16KY
LJLLTXX0KsfFYX/VWdd9f3FajhAgPVbseyTP5CYq+ja8XUxrEu+HDx01berZKuUH
IKmRDOpBbhVcJt3EsmVRLxnXmIehcxs1ukBlOxpdhda3RAr6/BTDRy7wpF77G/Lc
ssWniJwykGzebNMuJjMaVrCQKlgodtfRYM737x5kH1yfllVZKqrIGU31yKkRzLmf
BoyRHA3t+E6tvKZLArVqNYhKXkJUA1EtyGxyKGq9i//82iOBRWb2o9ANIjVuFLo6
kRQf6bO5MEVA8d8LQXmuO0US1j+L6rGhJnojyKblOoHfqgvoaSfeENKL8CYuwXtW
GDCS6AvHLvTcmRm36VK5kaXU4AMLlN8bZPqvmm6pwuLJYDvcmdqzWe9LaWa2amvc
8CHrcW7e8R1lCzGCFm9EkgdAMjAhNiU6lL6fDRPHnlc+wpEwcm1ECdGcLZ/rttsP
DJ9dVkHDVwOOSEOpjWxEUghDh83pd3fDKzy8pSQ1LMAslWT6DSZryEEhRRXCKHxg
u6nAvgoJ8mdLq7RHRqsOJuKx45dYGl6Hgpc6LnF/RuF6QkKgG2+o/1ZOtHdkag6e
Qhqw7lUQqEy4ZXvP2mMV6tcJPcUmqlgxDpAnQwd4jQ4qaLccCutUAa2ndUIApYsf
Vu5xzhAGGJMu49o/wt2orhD/cOlYFpuCCfkoYzKsBUFU29l18i7X4al4nYYTdYrH
2a99Ck84lv+XLAjbYtWKiBhU7zodFEw5zK+JZQKL1l+yvzIHIIom6aJ4w98ab0Jc
A2PQlcFt1A4Q/zce5Dl1TvwA0muz7pwaXUslFtPol7PlmTWyAT/5y/wct3eqsvbo
LddC3aU43/o1yNRzFdEU+oMZrI9Ni0pWT9A6mi4UxORbDcngtKUEpRPOsuM31vwU
pbCazdKyQdUWdYb+VmxJH9xyH7Hm8mrCEbGRATX78tv0trBFtNuTiSUDiHVY7Ogq
RyRu+R/8obpGAmEMwVJ/qvHMxN8AnG0w4nNZdn/6Q+8JBeGUGXrOgACpJV1URjlu
+z634tDs4iyodv/6LzKpLOQFc3U6SH5LD10Z34gxinvZdNJRhe5rZGcfgPLdMCyj
YKH/ZfFZpTcYKR+o/QfciU9WanCzFEWxfEXrXBKPoJQ5wS8rrZIRfXvup7B0NSOa
1PJYnkTEQ2wx/jXWdaq765Zzg9+ytGtvGAdxueq/GpYzIw0wLB9TRyfyYLK5KLD5
YES4iHsbqKsqTom4mPxV5ML8M6ZSgrXzJQXxGxCL8JHa1z3lDvgu5o6bXvGq9Dcl
vVRgT82XeL9A3lnv+WyOI/SalahCvtmqeNXJVtZ5UZBidu21DqNZoIlg5MG12T5X
Rv9QMkgcuTdP9fRNKdkeJsQZq7X+ytyHm+Rksc+6/5igwJ4EEPum/AapFclaTdRl
iG2XTR62mH3Brg8L3b1lxG89HuOfT7TBuWgj5Fqe16QqPN4eMfS92nyd9/UuDV22
cPrexrDNq56Nj4LHbGB4dUZtBH7liX35qXKCEYVlvTRmm1/KMBWLzSyt1cmqSE/Y
g0XhUrBB2tV8S7dZzPbX1/5tjfSKvb/WgNxnh6VVoAg0iH2OmrJ52eLLf+4hO415
GP4dlMSQRoDc6hmnPt6eXFT4161i2ODWrc7LsGH/DOmcOO9pME9gLJ9NXozAtIXq
QTV+czZpQUEaibCCtvVhdEdW4O9f1F1EikrutGPeM64abg3N/qt5LECgTl8hb4ra
75hHzMwMwlK9duTs5q6/aeYe03IkzpC4yIfT2OKnOr8eJCqKqwsTUxZRxsVIK/un
qFng5+9OdahCybuH3Svq/kt3p1LJg9QBVcGqdEh2v6a0uYMRQk+Ia1E3KAZdx2KZ
Q6NPBIuf7X8i7WKUmRdZsSbZUj13WrPuz60drI8gVsjEjJLJCBl/PKr//8Kccog9
MtFwQ0GvJCFnWdz8NWoxfrWpikw8k2Npd9uxz2GS1R4eov6EE18ItKDjQgkltLVC
oic0pNFLrpDcyUEFKIXeS0vup5Fzx1CR5mUlBIiDtEDHb5aMlqblP/i6l7oc0Yp/
iqg2DEiWAbSzvQTjOyuHRpYPlM/6HvCZdymHkIGbVEK8v1kc/LbdbFOn+42+1x4l
JcHeGs4cszYmmKRqxcoO1wESLxbJT3h85roXIoM+FuF+CHn6GyZLYxNk/nAbKTkt
nESuD9yQNn8ApSM5N6HELBfdEH52sjNgCEbpgA0SpNx1GQaeqXVhIaEFoHKkGxKN
VUqXGTMfvi9VY2rB+rtetjf2xVh/zuUro6ZwV0KyojvzL1n12uLuhX7vdcCRtd2T
vdnbeHZqMRxWLP6bWqMjfzX8ORKhsvjfuRVanYj+ifclvoxEenQyHL/5CcTXYYnL
HmFEAt/Y/qXOWkUSiaAihsA/x+Kq34ulStNfXmYzBoTDv0yb2DMmBcuDjPvV/Eml
Scw0LqBb+eROmxDNKjR4FwNbIRtcmrABChLIyAfEt8wzZx4xLqtA0l6R69CimW3v
xAhGTCYHFXa2NqMtQVhywoNXjrJv1MIBwbabsIpevPW8XkISfDGhzVky85q5JaSY
jsLpYdRYgZpy3eCO84CPr0zpmvT2+P/b8zekx+GVEnvV4Qnw0S3ccz8rwKuwUaVk
zj5K4tnSd0eehjDWW5pRtQvC6m8U7RddZhgkDaztWvhehIhfAy4MYO3b3SuBIoQo
9WJPA4YLiHGBZiWXcTejPuLa7nUmYcIyLsCbNp42TyeIQUXDBm0jkFQy3YgEkcGt
1L/sMnNnEDOtJYY8RbxCJbY29Mpoko9ZSLz3zdF6m85KDxNPAzafWpu0s6KkOrfH
9lANcWEDo9fZ46vfL+WrzGkrFg55Kx01bmsOguo8PrxF4u6JKMO8REJxg7y/jzrT
alVLAjwUkb3f+jDwnWT6mBsJJzEYP1Dx155JuiPxWnrGfr51d6qvzQoPYXcZnGET
2BHNGENUea4i1vXmLl3QXjtyUJFXXGny42ACWPJIptl8b51LCtFIa1/N3CQvsGpR
+0++f244SMk7UzEcpzzc8EbptC92phF5KLk3NqofkpnPXgTeIBd2Ux+Yb6yaZAbH
sopyX97q8C9scwXaIslkGIO1VIEk/nHKZzmKKjGP5snJhRICFemrkdiGGDb6Bj4W
Mzm3TwbfggvvIvSel5AZNqbhA6Ik3gmlmd2h1kM/PDt23e/ObMbW0/5RSjhrokU/
/zQn7kBz3nASRev4P5WYRChca2MD3GxU/zcYPA9feTlfWY/Ai4JYEMdB5iwfdwvv
f40Oa5oevixNP+PHJ6/EGiTo30214PKavXlwUTYc54B2COhqcUuquZvgIILxOS6L
1yWCvLnhT364Mym5DbJDZN/hULvGM2SOBFDp3XoCZap1H+yKPxRfZk9bgiOrn3Wf
Jo5V9lFQYuuTmkqSPK0aEG93X9XgGX2tm5b8R3NFj/fDHxpxDelsvDYnFacOKv+L
5OaIxtn1NOy1uHpgjHS6xxzD0QRP5skwl/JRAHIHNEar/l7+EGiL7whSkYmxE/ih
HphrwrZ9ESx6d0Euk+7pSyt5c0NKg46uNWG2HSZLXcfO5dvviSsJWrQZCwX0xJ5o
H/FozOgBFhkdtvXKpZ3rjUiKd948CnklDXaaTZamhZrkthcmI/gltRq90/NJncQE
SZdG0sxY5P7teQMXEZrglOxYzu7eSksFoxnpPlGn+oJp8CtMEU2OA7yFy8PqgkJd
Rujg8Yush/gnApoTrz/YpCC2KVosonPj+j72IjWkCthF5RhjKp2cDXKUde/NvLFl
qO+nJhLiM7kfSFKz+TsZbVK9PiVJcKyPX+1OLu0UN6xocAIEA98zAqUASzFXTtqD
Thf/7NFLY0CuOhhheEG9u0HpEFw3/jioAqw04vAjfmBJ3WLd2OYj6nGVTY8cPriM
QpuL51QXZ0zOsklqilk93xrF5I6pvQuQyRzPqwiM3/7toxoaRbheYtqg4LgiUmj+
U9Arc5h/an+vT0xmfxD3Q55VobGOJCccaopinERtd2MjxlcS2I9pEm6plbJ6MKIL
QAnC0JXo4qPAOzQNsjSZAHNgWkCF2bybfBdHdrUQ6iSWUeNOy8mFgdHOr+VL44Ie
rg/1c45nx+r9p5BvAG5GPwstSRxBKa7PmxG7e7lT0KVASzoxcXbTDbFQWeyWSYbW
+uzx6t1pNLxyqoY2tEyKQmuFmukxDSMwNutleBMWS7P74Ue1OU1STf4U1+aeIhLx
Coue7laPLTHNS89qea1rGgrTpFOPo1OQmKsWxXAMEvg2WCUBrWokMowscf9z7Oan
uVokkob5FG/ZzurjXe0/Isn/c8wtZN5V7sIGat9HFroE2exCptbgksTLkuzueCBv
8PEK/NAIf/ooRwTG5Nwx4MtDPfXsXoRwiONcJC6n+AOyOSX1PsdGgZpUrfcG64WY
gEauEr7JipO3zO8EkntEF7RpMg6nKr0Qzvs1FqhcC0edez4tfVjf5CgXCZ1wmqNO
csYxdzoYTGOet4QnyZ3B6Cuqfza1CdW0HX4mHO2ooSyhtwysDNeC5fQmaqYR/+Y/
GvDp71p6XH+pjOiJIPJX5OzPsTZv7pIy8On6JPFji4UZQU7Jub7Qv+tjZiFxrRz0
oUt1aHRf8Sb85OIXmceKrJa/oEtK0RAEDajex4AQO232hNomyJCFICkM8tR5JGWT
cpOJSpsYWgClx6tcPNpD3zAl+s0rufs5g3I3rbzFVTDcAXnWj9Ikwp1XaMTlQVRu
5rhT2gHezMm1RTGzrtpBEPVG9elI95gVfHAMzDY6Mso4VMMzoxxdLdTgagJX8KQg
zbB+sHt5/MQCYHDBRuib/9T7a5O7Ri9O1TIHqlyQg4gbpXtVTFLy5nYbJqgWId0e
+QVmJ0zfFHprBzZSJyC89Uypy43Gs2Ff0HE/APDyegWBx9Kdp6lX7pK/AspJvBNv
i8K49qdddfaM4dM7JP3R7uZwyTnqSnQ97cn1hPvAsl3k2rUcKfu8gfO+WBkQKkbA
g4xc7QMruQREzcYDoGQACKoim53nfjhcClTwPL53f1xnTMLouCgTJjZ9l9/Tiy7M
eDHzTcI5mKZwAveAA5ogJmdhtQMQLxUjCP6tsFK1C/6YDXcGAf9hXoEgLaXfivlj
8IsdMjYmqG4rsDHAxVNlU2MGV5uJhEFSYsTiTuHBFEO/pmvHNYpOf//0PS3EiQZm
TAQT68mIxVoz4BDVZ8korBCGsiWH0BheNImCnd27Spny7nAKIAur8+r8YvpVHuQY
931Bi92OeScW1qBhTygzsjEYYOm9AOYglN57xWPYBr8hXqDgsU3DUej9YWZ9xjFS
/fduwdYrfOtDbWet8u56CvXT7b/F7jolsV+ScxGDDE83kKZknE0X+m84xWVRTXu1
hEPJRaT/cYgYPBwkv3lhWic8TrY/RnNU/bi4Xkm193+YJV+hnB25IMnDr02vEuwp
qTPB5b/oKrVgDmLK+U2vquccRsgieT5ynE4wfqKkdUl/hQioTDvjrkT+sQOThSJ2
T/BxnkuLsdFS1pQ47bPKiossjZOsZDRGhnaBqRxn0OVtaFo5kRRB/ACRVWu+TVTB
DgfdCVPujsU/FjEzuEyEJfVAHoNjcq/KWFXweCcYarmNO+mRnuzqlCck14TtDA3a
gzvr7IjbiXUU6rsQDaZNhiHWgzlDb8Ll1sK2ApCfzAH19VsITpF8HHSl0be0jkly
aTUwbYM71ALXWz37oKhmBxYx9cWjqDX8P+icXiOWyMAB+DYvWYtOmW4CI1AnZD1L
bwgQWU2rJ0qK2MllgzhyiJLaysHO4qKVprh/tanYC9FtCUsxQlrF7r2+7Evj/8aY
cWHkccn1JdQNRBYV+Wl5iVbANrIxi1dhHa2VLeNnjvXC3jMYpCLC6M8I/9lNXdU3
w9rMeMUz6WnjEGDFB6ffadpqyi/cejPgRKpDOvhO6eEuLOSOKk5w7SCB3olpq1aP
uC75G1gFq/eZzhbJBaib0QOaIsr8xqRoaf/UE83xqyqyDUpx1cNrZD5jjvuFeBSr
3Y5DJ1/ezZkxspqMzsX3rhgTwk8qwAIVMC8zhnn8WmZ/ucgKyw2xkdTEEF6tYxay
7Pdwm8CaBYQkSeVyi91uG2dwWwHhy/1sheAYbCNfUyRjuyuqIzx6ceOwxqQ9osFe
wQMLtRh0FNP/57eci1QwdtSKZS7El4HHbk47eohLIapBziwuLLpPST8Mj94N9dlo
ql7t86lwVg7294cUoDI7KLFiBaVJZL4z7VczZXgIY0iQLMh7rGYVGm+CRo4DP99n
gVoV+yk/Q/msZcMrF+ysOEXyQ8a5w0tzGgw0/nXUXTcVaievzf8tV7fjYKC1bwFA
YFJ0LBqebhwR+fKCL7pEOgwffHyUvA9B48oXbseMQ0KWba7MvJPZgddzPsMaKS01
APjYWzSxvy4MB47FB9zdxPbDUTFDDY+ot3Z06mVqlUvS/PjBmVdxoDv2fMobg3eD
U/fSnbd5eEDE/nCcwO2KVt8TxkK/PpAGxX2fg0Cts1cEmy2SUdDWNiItVyhDt0JK
VmjwbcSXfWw0tdQEP4WwriHoQoZVtiuZecwXwZM9c4hY9zOFkL7xn2IE36Gp3J6L
3uwqErRkwPVWU+4bZvHJdo5sT3IosY6PgXUAgyYCtxGos+5H1OlFYVQVYyCaD82C
kuNtYkv9B9960i0zyO0ydrJVLoZ294/AXoXdNXZhKu33umPD4EzzIiTHwvTp/043
f7rZ6TcrECYA0eOQImR6wsojCnT1Fl/9Vy4mnaO/ufCirEx5fG3B9rI7+/+RyMjr
7fJ/+QKts4lYJTMMms+s8/oNcaTnREKhZ+jDwuoWjytBvVPiKtHn+O2oUg94NvL1
x30MxYlwKcNKdDY6Oo4h57MCxaBR4/PkDG2wDGdN1xM5pauICPOr1FTpcAOJ9kvy
Y4uBG2mRAJjCxXzT5AkwMfF6A3S3LCXfo963LRv06EFbJwTWU9ke1kkLIRO9nQPZ
J1tJcC/0r8rlVPU3tQIkKqVcU0eLFBCwPPS+lVvyzQwFllPW0fnDchLSG0wFCegn
JV+gv6BaLV/oWwNnSDjSNMnR84zj/10gKrdE20T/yFPCEThzXI9LBEgecvuB25Uw
xgRslVy15InhZgiH+m3he3Zon3Hr9eR4funvI/x/6631tjiMWlS1OPeIdAMx0i7O
igz3WPG7GZue0gwzNVk0IG+3LVgnMF3OpxLs2+4RopE55hjjeXiCc9NAdtZUTKpE
9JmibKHBk/8wQ1YsRmdacA016mANDyR5TXqybm8UoU+lCsMWiF5TVchCBqQBCmrQ
R/dUxmFWIzP8Y/2pzMa9GjI7mB8jQjjB3C7ZoT5/t4oK2VyvulS1UgafOMiZ0Rhp
JXMJbmpb2aW5pOUIppvbOzuhL3L/Rq/+TAxI3tLACRBxfwfLc+xA4nqULaAcM3Ma
zi3puZAKKGw7X+VntC/FLRy5+y8SbAOUg5OqXE6Lrh6t/yZOCj7keJK03T4LTO4M
u2cpZcCNeTWOsDl/qaJKJ+uihpUF1GQXJTni3JzHcnB/cb01A0xXP/Q3/yju2e5k
Ri9aFHIbSIj+5kg+VizWlh8SohTNz5xy0OkYmuhcY1Iwu7dwAeGG/ajItBUHF+Bl
2m+N5j3gVz6zsgYqfYNeMK2t7OycbLmiiWL3rJWC7tKdcoBxWjmVxgrZkQo9HpTZ
r0W7l4C7Q89UJyJf2aOsUgPlXViouMquAfP2lsok8XQpS18xVCl+ybVOacJDujTt
Se1BJt5VQ6IaLEB65qkuckF1EPDiZ9q7kJH2MsYvp9aYCh+8aR9PY3ZE/F6aF2b3
NmDJMcPSSIyKXtuzt9FD5RcYYBYejwJIFqmoDUuUin6Ti7tpPaCDsleNTAcABp5F
i4M8X1ercFVsVSnuTVNmKF81cxgXYiYo9lZJ4ejTiFhHzX1zPOjYO4YCOMLHu5iQ
dc11Qmg+fytPYz0Vjs8IqnsvPrtxI5FZXgcK1ziBAQ9BqjdqSfo1TDKL/o/0147q
GbtvR3PL0OEZGkdnGhtl/5DM/+FzhFLqIPIqnkZ7q1i+5LluYfh31LguNYuNQGn2
BmMPQSSv3QTMGC/Q6XrBrd3AZj8WqD+XSuZGQWmj/xEGcPdCsPbfictiZU85F4Nz
5793yaqVqzlP5tDOC9nNUpIB5MtnI0jtT/471lO+HnNSYfiQ9KMKLznZ3dLtligb
aVm6KrmipnvNUmNCZ+Kc8gRRl9sMjZXqMRDiFSsRstSElqUa+tNS5XrIhiBAIHCl
XL4JGbu8pbjhcfLZD+52VPaefLjvPrEnSl453jHuy8Y2gh8p3Dbb9XO37pah5urB
sv1dmBEdUj5xefJjTu0x7/Ey5sR3inXXYg6L0SC01VNIkc5JNCp39bRgkqKIaCYx
4HNeP1yKHBQQuad3DialpCt0opA3D1bzl2teJt7H3l4jKikprn5XUqeVTDepCvsY
YrDqo9JNNlncNtgTY2hh/sBZhSbh08U2Ru63F8+yAq3xVbyiNvrnHCdfH/pnPoNK
HpeG/iBS7ae28EOE0TykfkJS92EGwmKDLQ6yDO0gsVJDplf7lhtdeKbLViT5pNVp
H6m68FRUXC/wKLPi8ygxxfeS7bhfY50GOmpoFiOrxqeWai815StbPLIOxBC6KTji
CNoaFuXKUf6oF4Z3IbQZQX8Wflqywtn9uBlOC1cgyvO2VI7aiTILWklLFfsS44aO
zIvK9XAqh+NzXadAZdjSbSNCihaCGPFocp+IBXK1MlfgbqBADBimPlJU40KG6lEz
ECqQVpO8AUJDoTpNpk29yxhXvWI1gfhrAar8N4vRmibTWTEIe4KukzWWfy8jK4Jd
/WqUFcO22LyOy6Bff70tcwi8PomzgkD0xYtO51d94QyGudvZOfF1y6UmGIs9wSIy
85WTgUl2F0gZPOpfZvxsJV/CeMhCcJxR0E6AaqOTYNnI0QLXrQkvafq0ef5Wfp5R
Z15TjxfsVoASkq/Agw6cj6VQc+X0XGKR7/dADAA0fxjSnq/X3Asg5pGZ4nSROusR
oXysqvd+2I6VxZmkkU9HqXItS7IK7EHwYKqXSZzF9j1KuF9autnM0MAFo+o4vvmM
CW2hxBnqHXymn8x3oWYVPsiN/g5yVS1u+OsIXPA5IC937Gl+UhhTSvMDHxMBX3LI
rfpUlN4uS5+sR5Ac/FM81vrew12C6f37qpnzd37/38vcuwLyo0EtpZgRF0kuhjIK
g2+zxJOH8cr19zGsVwRyyDWFWc+SnE9wOzQyGWacUZadw+7+KDHXvyOeG+6dOBnb
WcgGMnxqjUromb/JxGRRXplfW2kC2dwUW3UQoXg7leHKLdXRwcemqlBnJ0nwNYLO
6znFugg92h949LG4vvx4wD59fAdCbqU98JM0rry5r7d9HMnlJpbRTiSttGi6UgI+
xsIZ+BLMMZ2jMx5tKxWfjob7zmkEooYAIQEWcrvJEjGQTX7Y52hXuVvTLC+7XuoZ
SXAb2UKI04NnAJOGWzUx/7bWP0y/eEAZz0ant9IiPpPhYmXenBSwa+FHr0ltuPI3
bN6WaExtXagy72UAmA23QjTe8S0ddGM8b5XXLWy4+QRfsX6NmMdm2Cp/hwM8ed2J
sPNEMsEpcX3mnaQaYp2l3+LhmPlwFTm67wKTqSkqlzSAd1SrgDEGD9h4hhyA9VOq
3SYhhAgrp0oU9oyzno8sXTbtrZr2Jxs3DHccTynskOyTWdx4LiX3IYPSyy6gOj+n
jbAK2OmaeHRQCiyBTEZi17Ay2Y0MAuEjL2hGfUXmNJ+QYwZFnyBjDyo6Q0JTbSy4
OVYBt/l5yTYwaKv4C6+VSv/dVAZ3scu/4F6bdvX7pJQ1nQiFD1RA3hZxYXRA1me5
e2Euv90upb0i7WtGvgcyo9Bv5Hv0COzsqm7M9SI4mcVhsNYKZG0UcGfZ1dc69Ilp
eneSLABcd5lw+4fQHQInFD05SV2JLtsRs3Ag7441Og43Emy0onohGohVhwV72M46
My7scDgVMeyd/oNDmVb46RxoubMBaJU4qTxPjCsKQ5ZZMva+FRGj6fLk2pQUW4mL
uQ4NAaeL+AnOn/S6MPMM6cZ+bRLaHyC7hTU07JcNHXuCqlFbpVth0vzl/nEjDlNF
V4Kec/pkaeVtDSvP6gVM1SmFPbtNnZ7GfwV7H7DvlazRC8R6nh5kikoeiu5Tzzq9
0ndM54uYImglT+8T+kgKczf8UyDPnCVrPjenX8QJDhfqRe0p2UM4Msf7PhXGFV7F
1wlwy7LLLAlcDq4IzDBMg4uTRVp3b26kAq0TKRHzoC/RqhomWUkPVB8jEQALwo1z
43bCHcCgAfEGoyJDHbIsUBAWtfbBjbnK0zZ9GZlxm3cObzlFyd1Q+LWsy4wm25m2
6sX36uyfSlHNJy1F59jhlGI4AEcHipyKmWBgJoj0Xe8YgbjwgEoqP8UuFja1GrCn
tr/75Onq97iQd1W9U0W0VNHvNHoY6YT3ZkmBTjxOTMHsh/qRcQaSxhIjZZkfZMA7
kre7nirqbi2+2r0xpNzxQ0LWpYeFMXv/3DkWdk7MsthJm9JqHhoygsCfEi8P+c3l
vdFc1s5Bg4h77EkDpkfA93LDlk/VDh69KY+9Mpv3zDxzHVGvkROLbgFAtyvXzUe7
qjKkBT7ZFNBW8JJ8eI8wHSqTHFPhl/tmWATFV0JooWI9nY5tQKBNrXtF+UrOU4Nx
/P3rl4V0rWv/Zp/42NZUGIwmUEgCHv7H/ogndoQmuAlIq5J4LfD+Q2f4Wp1iGnnP
CBcAjZF9NsBGio7ZvHUgslK6MuHveNIR7QM9ew7RDiy0Tkr2TFky9jnTlUqROlrY
QN0ALdnb8xIHi+IBVuBqpjQGC12TPmDLrD8wv554FTGvGRi+GcLddKpVVffLc9in
8Xdi9LvBT+GszJFlwQJzfYZ1thOmUV6eb/d5ptNi/oGOQnDQWPWWPMKhUGeCZkZA
6eB7724RVzTSH1S1ZFo5HyRCHJf7In/fXwPgrK/nvrQw8pAPGv0NTsnMjCfEe3Ge
AgUxJo2OBIlPh9JXTT6cMh0KBGHCcOe3rdang8EliDAndSEORFqvwTkPXeuA4emT
E49Ia5rO7hyBLjFCmxsW5HpF7bZTiiaXJiNuKger6TYARHYbJTOGmJVUVUoZF+4h
CBCKdbct+WuyhWVqbm7pFuXctSQ4gVELkgRp99o0NcLfQICUwiismZv8LL53+pSX
k8YUx/iQhG/6AqM2ICCSkQcRYpeo7FZvvJfFzHGvAQ9J3HqAfthAK3VqDqGn13S4
n/u8wD2Szq349t1VJnu6LPS+6lDS3Aq18AXcB3QZvJmArH1Afwiw5ssHgeR4CF/U
vJthG67I1BWVtN6U4nXg7KE5KrSivyevTr3gJjqm3pogKDiPy+4W0YviCOMy0uIV
2OjwSBOCM36ag2XI8AeFMIAqHn5wLaTjFHP4rySnxNGhsebShmc8vrleiuualcAa
N2TvA8xaNsp69tuGsKjH/0aFcS1usPs4E6u90mHea4uRVdztDUeGwstBC9ZO8Snu
SONLcsuo3hE0vV7t1UtlA6dKDAZzRGAJ/uTzkZkmZb9UWoBtqA2u3UtLYvbrNmvU
Dj/dedTXGtZlxaUxaf//DvT6xwHVMo1kPBD/30N59TgSG6e7voxebqZJr+gN+4cE
7cb20u+pkUIKqHpmD0JVdRd5rpUzmLuHD+ZuB1V9trZnaeeY7Ls+I/tyOROdenJn
YQxvFHnyMrP9NWat5XJ+YnjGRlaE2jLeRk9z9dobiw3B6U2wXFrPBulid1b2DC96
gaFqn2j4CQk7icBdZOGTRQlRBd0og3Hjjdn/vLEb3SyCLCfCHW0LoK72tCZpz2fR
cxjADXEp7K/D0ZV4kwRswZrrUBndXJz2PyxE0zSWxLYNmyPaQ4fq2+yyPeyZPEW2
p0MYaEmNCCSuYM6WbeWXzPa6voNCq5NqB7GDJ2SKIXueCYB1peLqFiegwsXugXjn
z70xY568nF+NTeF5obvmoIOvPYeL1fx64xIGZLIt+/Z6zE86YHrUa0QYFN5B1BMX
P60YNv8HXvadd0C1+d64l9JAWYRLBhhx0hdrFVRqGToLofd1XJVpMqiXlHELGwio
D7lI2XBjdocCSxsAHH6TzwEYlZzAGndvBeMrEIB+TRVor9SkNNQw3ViNLkr7MtJD
1iRbbqyKEm9+OJJpgbmR+vgKtEpHxJDGqlvueWZ37WKYngFgapVlAHFr2XUSY0Bg
xXtkCa1UB2qbLTA9fjvNA/v0Haby1B76Fp8pZJgXuoNwdavlDIQQAx4QZaoFnz1q
9wewwGrkQHB3ajcwxy9geMLmGhM2XAqLgTdtnoJZevw6eoMDJmel3XiPab1d2zxt
KJz0PupBk4PfPa+4XWEWN980Efd8Rbrnsfm4UVW7iyQLAM9RKi6gQ0YzPUPmXJ9d
CSvSmOA/ik2dc3qBUPTwcJ0r2N0Hyt4QvIy0k1GZl9N7yWCDDEe9jZ24uCg6W9Jv
lInmCEW0DeDTcI+fxiwTq6mz56CxsnO0sGFbvjZmnPRF6V5Fz/NctebKkpZLQFzR
s3zFJOmTgDFPCaK7nOqopqoqFSykAq/Klj7xekQEy/MJlTHUVzKLRTYheiC82plR
Gkjvl+MvgL8/2ae3AP/pRMSB06AtzvKGkSVS7zN2t3/jHMYGhXuS58eVFKD/yDOn
rBXamM76ED7hSTKM1gAbNBDCLMCVKAadH6GWrv7OizqDF4bj5aOhiMZwvhz2PBrz
nOqobcUEZnJQFdZwDKKnHbTy0HYfd1/v3PdZf++0r3y1U+bzl3NfpH+XY+1gf1Z7
e41mIHl1LfZj+fv2DmdwmmvHgNFBXwxKkiyaph1tvzC28+iK4rjmwCbNaF+NdJoh
123acpthluvQxIq9kLrvClHy2nyna6zscqK5lh8cs3KNV8zgGbKs/ztU6YIAqrKY
tJ+7FCs7910TNyRrORy9Y1oeJiSHgs64+zBIRNtnVOdeXoC+R/c+Cgcx9MSXFIU4
r2wEz+du68tshnYfiD2wJly9/t3L11dCT/v3ADJCn8mRFIrDRe7SBkX0COAnGhFN
qrTRG8LJGfyQvTwBqMcKca+X6ba6TvDRR4h58c7Y3bd7yrxCbwaAb8tj5Pu/A8Bf
NRYI3TfmesvmUdNBle3xcdPnMtj35t0t0RVBrT3wY6VDajd8DTJipg69d1mv1iig
riUcSirBHyK13Cc+DE0Im8SdVuzT/e25DqTELynOkiNiF3X+DdxBkkP6nkEEy8l2
nsfXkdwhKcumWvRWEtm8GpCp7/NSMiKyDlXyXm0u4//zRCuJl9C6HIYd0Xgv8LiL
5ZTRl5H0XFexw2eDXEUbCkR3okbV7fhiS1d3VdE0SBhDMn8qfbJUxU11hgopPojj
dvTzxNBYoqqPawfUZVDaef6uKqUyQSnD7fpTbiUJJiiWxHxi8LguZzclfPgZyG39
yKlDhfcdUWFqyaMZNkPw0KcXk7npnNSHuMs0jG+fyaHL1mGUzGODknsboWm8SiqW
aZz/z6NK/lDhgFqoUlDqAnzzs0lIZTDhyPA5Dz9JqbfZDpd6BVpkHZ6sJGoJ7A8+
EBHNespAwM/G2iyGOnheHg7ibxZrGKoXN1vLyNBWS+frIZTe+zRdHd1EJIFOQZqY
i4diVgL10Bti2OylB0BNNYrAm2GjzDwQgg/kL/atF4Fni2xtdmh8zpTADMtZRBGJ
BDMLGhWxkmH/GxXvhaJendgcAESqlRZL79VJ2IeoeFgvksp0tA23FtL31C3eeh3L
iibJJc0Wy0At50ZGK9DAjCf9xmzAFLSqKWQoaiu5l/5YaEA8Rp3D8lmWZfPHniv6
UbaBeSceAfHPofUapVbTow35TUNaVEGrrkcRO4widWYMYlqvJNmazH1K5LTFyuPw
TV9ZjBiTo6bx+MEsjzaXvwTu/ktgySELLiMlcxio5nUpFnOYHzjnWm5JlcQfAl3k
2FtCmNHJLm1+XOgr67vv3OlGI1o0whsqmy09F3EKCyFf9n7a0TLfymxU6XFhV0vK
Zm03+32r6EpVXRQderRtxc5zfek86GGzkqrWi88MXOpCryIfw5NI/HIQGnNVN0xu
wboyvPzGGF6HFzKrXRYuLi7a8TdNDsTIPy3+g6wa14m1PHIR3B7+0Y6qjQzyRnQ/
Nzm+ZKq1hOjBBgt+7h/znMd6seyhW/7DIA/J7PrRzZh2kUZgwvfYXG41kaWj0rrN
TOhpxupSn26fpNos+giAJroBb3E/SiEmxiWJlumZGencN416CuVvtRW0LQohIw9g
Q93iyoEwY+R9MdL6mEqJqBS0pKahWX/xmCm5JFruuS9Ih8KG0kD2sSqxNt+2MyE/
tO05IsYCT5sYip1A00ORyRjzS+tFbjA+KqVuTaNa9wcsaCYno2JmvU31MGqh6Mdw
QS/o/QJIkfdCjJEbOD7JzC4UofOJyutw/bBQOtjbo2ySgjdVZ+BlDKeXWIBiw3W4
fjjzSkOf0LK0TixZbMT1BsQHtg8VwpZiwBWMgCBk0NDpVti90JG4dDmQeVywjKEa
fB9OiC59k5SefHMHvsA1icOCJUS/k8eUvA6By9cPs18vNz+WV9UnTSHn9kOr8naZ
h043Jojy6EsWh2mF98UI2oocGZ1FfrVJTmZJZJoHy5aiMQ0rtm6ZjfYocSZ52eEB
K+ME1nFjG2B8W2ilg66pZSgKehRHGPhFyG72q3dU2pwNRLMfozesCy8B1g8Y3ruB
MEWwiBlzAsEWmbzOC+TNCdSwiq926ZNeRDz72PElMhegjAAfo97L3maMOGG2ngWa
g7k/+sjDKua4E+5w8Ntme1gFizqi82qYchyi+CexJR/e+HJS0cZjlbtADplzXevV
l2VAMQ3ni+PWmEM1SJhtuLHQus6lklI+VZ2gPUn75x5XPh5BscT9GOD6tAbfELFq
MLoD7Q5KfxI0qYspBbctkYg3S8EwPHBPSJjr5vTPF54Wj1rL+R+VeHvDdZGFx7m3
+rPzWDpEuFLzN/61Dz9PTxB3BSzwqDsRvLGqdoBPUfPid8T9TEShFGIPR4mO4TDw
EuRT17Zsle1OVFCfvJxElk475qHtbT5eyPd3UNqG++YxA4DNG0HwekMDS7IjWOOq
PK7yfyM1JjVIT01NLI3qnDnGTA/6XoW/yMQrhZPUMWm/pL1JIuuS7hNzjuPPyCU8
83hWt7NumFn2BFmcHFWJEJdTOgKo2QeGQ/zcpnoe6xyHBGdwCnsBlbT32UwEqWIG
Eiw64C0/3QQuuQDKV+avtsEg2RC6KuNdQulMZllloTudxzHywfzaJEPzFWtvXmhQ
GH/6bqH0FQPWk3oRPtUa8vl/LNBIy3IV9JiDkrGh3GFPRx+bJszPpY530wnLoES1
5NqPhsGPFFOF4cC45z3gIs4d2n0sRA0RHDOipDifYx29qQHw7M7iI4TSRJAzd6FN
2GeGZytkHYCl2BvrXQgtmQIofA8+t4wULosWY0XCug/VzPiAADhh8rSHgzepebfE
A3g8uM3KivHkveduaIzPwl1RZrmFcAudtlaucUh3cYYTYipBstkZiAkAXIH/Z2S/
bBB6b4XYf4Opp3HCs6r04dd4OIdEawZ6QM02VKzZFAaGTOyW1iHJA6zf5FByLTcn
KHjxpUrFAhCIyVcyMmx459VGQknj8GibQO/1g/diWukFSAjmDC8C1EgE7+rpxVy6
bYd040hUTcpzRIwml3o/c/ATgN2isIPeLgS7RRqm8uaXjIOrcAwlhTGwRhaISQxN
nUcWhEVMEkWrDiZzjz+0kFs60tbLiJNcelwQcF50tvYsI6AKNwCvWwFR+8U5d6GJ
0Yd4z2eE+jxiCB5VimbYoJzR+6rTJmTFZlfq6ePTdCryMJEprYmdi7aVdTp4vnM2
MUkmjf4Nr3mB3gtIMGyFWdooZ0ZhNnm33c3IDQCJPUI97kH+t7zhcPG+DIoCD3+y
1grh5JutCprcUYrxmPzHt/K44zGoGYASzprY0w3hAqL2ZsVaUD3OE2Qb0Hz+U/+o
vQBSUKfNt6+YG9jVaH/Kj9At6Y3jEscNT1OQC+bzfP01fFoJ/h8SwZgkpig9NhTN
z74rsCO+qApXRr9s+wAqP/AVfC7XOFmMiaIbdr2RwkCP+kmefFIA4Hkd8mNL3XqM
ZxxtE/6MbmTuucCRNZIvoBMLNOrzxHwmufGGzlAf8u7uWksqczvPnURJlMFkiDF0
23lsOzNq7NbFHwen3A+HC3RERkV3nac2Vpbz1bcr58Hca5S4LBiu/UHqrjWXSqAr
I9OZfwb9EZyLz7e4Op7s3aGgpnP8Mfur7IS7QvAn/SmFLVUOpwaK2oNwD74NNAOt
PnL3U0Sfq3IBg78MWBivJrPgJuydsQgtjoiD5OH/S+GeAzTJSK1JSW7gWJbwR74o
5odJ/To0EYMhvjCVz0/KrWHzmgQZF6Q5prNAv71p2xJYvAt4aR6lkJ9+lwby5K10
CCAIOzcJbZ5T7+Lftxl+BLFIFsHNAXp670Wr6L3KjulRCoGkXBn+LjvrOAT87TGs
D/PxHq04PmsJPqYuPwtE3VlHetIea+1qiLRyx2qgbzHxtcUMl8c8wlPH/9aRPvB2
/AshAEE9eK5aUPL+c5SndmpNGU6ezKjpZ1lBohBqlVP28AFWtb1rya9UUdv6gv6k
FycRLHoUFxG8I3M4XviTPyDLkvpcjte33XDOB86nsEaxw3Il+CAUEwaLuIxmHo+m
g1mxOvZ/OyS6o9mka0l/fC+ovLZI7l2MOcCGFHc/Bg8cIuivAun+2BO4WRuo3R4y
eNfCe3Lo8c9bl22n1JEOg0/7j8nPBcv/qILFPsY0bRikHTo1q3hUHzmLu3xjWsUx
IrhJaG8onZ0SAufGkCTdiQmnMB+8FLIFlF5XcR+FRL1yqqzuS9OZB+9RYmbM5pwU
S1Wbu2RUKGMNZSwUdRKqiuxfJl8fD3esMOOX1sOXnkNcqybrKxFzpjwRFXm66LeT
D6B+a/bt/Zn7/+DiqdSadxv9+px8/9Sb1Y8s7Ewx568cut16S2X83LinXBw1gVOT
uszvTyI5sabIxy9yyRRqOwbaEtaAK13PRLCXnuVf/RjHVxnyJXvltODrp9VCTPFA
3dUPxLgX0OkRXw+7TQOOJouTUHlN0hd7oKj+0uDHAlwrC8SwZDGlpPv2uXUWLrYG
8d5fThsUgzO6/ywf/id69+m6hMlrZpMEi+EC63fwCm8k9V5MWDeyNBqjzqAy0VTn
MW2mxZjC9hpAqt05JILtSvPeI7BXUX1kwvXOXEwYFt3RNYY7d8BzSr3ovKCs4Bc6
brDnTT3JrPBbp2UGAgUa+T03UOMdoDN6edElwqwV9/DiTgkqLCvOkfBe/0kmLK7m
JqXZYMSmWrcd7xhYAZtgvMdY/sat0Imka+raDk7XtpaQ2m0pxH85WVxKqcax/dwy
Y4sWVaxERS7vQRTaCgAkX9TzcIQyKl5sumbUHi1fRQoG7rA6vjZST1DsigoCaVT6
OGDh5vA+bL1Pqa6nhbijXxTEmL4JNjUcCNgoMdUCPr43O4Ojambgmjd2h5lkFWPk
VGaMmkZQnwvPLpDzi5ddsj/YQ+cLmJfeVV/2WBbLvflHK1G76g2Srzn5ZBlPvMT2
KKFFhkSb7dKHzcJ+IYdNDBKJ8nj5bUFtcbEja6SpHrvUZkVZHM4vhS2Zf2KqMOuA
ukSidAQlm+oc6YLzjnaFc2nJ/3sye+AuY0NH7PuKVsWxQwVM1Ps/Kj/hrxz39Qqc
NPvG3JqSwVE1ulrvcDMWpK9teSzA8o8RS5BszL9ts81pVLH/D8odAXZT4REsSMr2
JL10pmCvxY/FfZVrtGHNTKW29HSSTMytCcgLq7s33qGdRRdBQsdQu3gE0RB0hW/2
TLH51t4xaNJKB+eDV7Bc/n5oImJJyMUFo5UAa3cB4w7+DpCzZEHq90xMBjRBAgMl
Ul4MNrbv4BtNHlHcw2lJkqgC+hFVIRaDfGhlao112bRxowfJ3f9OTc3El21NjqZr
HBqYTGbMJCm8MAmHoIGuxVfiS6XZfl3ISzwoHt+d3zt7Tw60drN0s6fuFN/hbmju
9xjjp/+iBAnSuzFQSWQOTJvqCb4EgSWaTVZ01EG/7GTs1vMuRXAgzI1ud4BN+7H5
BsnEISHhNrp2ETbLyZmHKVHtt5MWDWgAK4fM5UcyUh7HSynfgfZSpJrneqrNqkUe
qblDM7gJboEz1c5qmKMRcOqwiM6vN0uNDYKZTsdw/5hQtxfvuNh5UQm2wapH8Cas
wBBcyM81k+xOToPbH6362zKI/PAQSgDwBg2cCYp2umUvjR6/NW3GKqQRNO4966pV
7zpOhvRNXeFrGdSDLZedDzCTjagX+z7emIBTQ5edNsmek+zm+IxwQVOsaqBEztmK
AZAeN6YmouGjDNbxtkPfRXpYYBfk7nEQzJsCQGGpARR+TAVU3wb0MSxshdPxqtiz
ZcjyYgymLCYtAFq0q3fqt3bxIctVmZ3V+K0mIsydHi3qR+S/UrXEYABIL4Sf5x0I
rPvBDlmEfNClH+JUjWEt0WRq0Py2cFWf+gUD4IZlpbM34sElfMtvrtJvBDnNObdL
Y85hlMrvdV6DYUa/ZxxF/WEPQLDyeTghea+AFcBfh26QeVynkpv91AAonk0zq3FC
xFu7iwfTJt+rdN4oeYz/Y2KDpAljMXSdibFlVEIDvCP3Vb+uRAKXl0D7cF5SkEW0
GNg4YC9CBLfiWsgNGT4XN9w3zxXuIfCl/nt3oi80Dmz54NT0BXK0R2KTpr6oqRmk
EjgQvy0tl6lu8chB3XfnEBELdp7AP7IWZgNZ1nCEiX6em61mFQ/PbLq1E7wCvAY0
0byj5oruO13jjrXR0FnXY9vyClutCWZ/hlOPuNWHFrYfuCbnrqjxnBJSjRXIK3fr
BDVzVzeEK4cnXZMOIqZEb53Az45JXEPQpNJLZoNAe+Kkma2/wfRUBa2XxlVGgxte
5bNx4zQaLipQyC6CrYVxOdfpQFfU7IZDaQVz8RgnidqQPaM741vxBmzeLWkvxpP4
aRNlPvRDEr6X98K9arkTmFMPxLWPMh/9HZuLAF3OqhsNzoYW8cvO4CXBjvsEMijE
dyQxTvF0qlutox3pIl7s2O9NVLJawjMLEPo6tLAXmIqigvlkyS8HzjF15iBAaeXJ
JLhYKzrZpLYhAMqqFuryXtFrfonhSpZze3Fc6QrbP/9X/X58LEYl66s7d5frO9gp
Pjut9AKTp7n9vh5dg6RFImnzbTDg9WkACil/M6Hm6lIXN04+LyMYh0gMQi4/ZWdu
kYfX1nlBPmwnj0L1uHyFwxgApnXQf6ygvpKcaZngp+DtaLzXORt3tWh55ty19zjv
B5tmkTrl8aZQKZo+wBWkt1cIDpXd+VM80OxUNMXtP6GpScClsCDoH8L6sEmWYVEh
Wx3qiViUoc2/TBdyylgRp9B7WC7SlDgEvXGuvB+BDkxUlq0Ck8Yyptmw/V2Jbut7
4p3HY6wKRGw7itOl4AIEmf7ltaH417QqAEvkIuhGz8O72roRTE6oc1YTT2NX/kYH
2PPPhvvACV5uTiSbVAwA5OWvdk9ooLIcMDB80l6mmyIhLEc7gqX1lzvkRjTL57Jq
+Mts5GP5RQ5VwldQbuhHK7zl7YYLibYhGANRcglsa+XJlh7XK5dx69dW0noXdpKw
KLiVLJGfO7M89hYDke+d2nNJcYDGBHCLPMbAk32piOfPu9j6CCbUkXNUFuRlyZdT
f/hDHYVNHfFKJwBGWOBpBFB/C0wO4ESqgop5ZvihlU2Y67q57dD5rB5Dkz7L5LWg
w6t63XBAEgBi8Y7bBk0rrrOujMh1Vw6CpOUw27eluA4YWwZZnoL/hChJhrPU2cO/
QDlKmQ43fHIhs0ypRJJNrV94fV6b4ZDAOW5I8TkvhVOixeTrYXEmxCqHpiTPSowX
uXVPBSwMRgjzN4y4K/T/ppm8yIlHLKQEIx6XhpKF94D29VRITxUlN9nmoF83Vo9/
AAWavJiBAOtGmq62FE/B37E/r6R7woCeuojB4OBb9q/b0YJkHM7vVenUyvtuVP6P
cadRvSJBzXeaq1foNc/HtEFsHuATxa06DjMVYYaXAVJOgo35XDaLt774gXuyGKnq
dqpLyvAxIGjEHDfE4rBcqCEY1f/K8zQB9XHmCLGtZDSP+V6L4Bb+0C1rJUYo46ZT
CAc2RaROdkcsM+BNDiedR//uKa/TOCQNveE4keBBi8u83fjK5p8PUvYZb6qW8G/u
nYLbEdKYQb/+mYVeA6LLgi3tx3nEeJdO/pyvU+q3/K7gjpWCVPTvbRvx0naD75Zh
P2sZs/HunfxPPRXYpC5f77WZttitmcVJNq/ybk2Xsi7o4ze93zzwGFX0QZXacb8u
DuChgKwmixfhzhpM6BVfbg9E/ZMJtLDpoK0yOQg19XKH6xwd7S7hzqoQu+KaL1/x
A9NZdzsCosxQ1ExfOq6909UTVM/ptUfL2xOZP6mmBZdgP1B/SPG6oGjTJbEYlQPv
QBkkIU0HjLnO/3BxFd4v54E1z69drsdffuiH+4lzv1Gkh1bqrYQb41NAxz/d9sin
WK1zhqwXie0RUvb5syUY5slVkomRhh1NfyRVQvuXb2pHewS6XJidkCpvTERqkMV4
XXaJGt6JbeUEAt1bRn3L2XNEQX5Llku7SuI+ivp5XqriJ3Ko2Ggukvg8VkjampMe
sI7SufdjKIXOVRnFLHxhlop30KFW/DH/Q2LW7zavP597SNP08Koxf1eDEHCoVD/z
xfich9VhrUQBbSgqBO5g1BGSW+gSHuSvY8ce9GMNpdWlxpKwY9wYeOTRW8eXNhNv
nflpq4uxM7V/M1z+61kd7WZ2jOzkhzMwhhoUekxBp1/O8rhRjEpIrHFzaEIXmszd
uk8D4a8qmAsUaIdp8MtjQSj+YznlM9dkZsHI5KL1CscBYqRyJGj5tk+pAH01cA5B
8EwDn8+a1HRnf4iG1lRYb9CbnjLho+GoBkfmFTneSguIKU4awPlUje0T96DQ25na
MLwktlm9SjjYDAMOg0fC7bxcWn8XiXg95RMJvx6opDwSHmrpT49ZG02SCU+6WBas
Gdpev6x0d9P8TRhxNAOjq9zGggfbqoF9LcJVDRp77OuXvC4guhUx4l6sniJ+F++M
6iVAN/BDqtE2Up8JWsXTbEFbYPKLSMj0A3FUzfWaTctZCuUtNUZi+I/OvpU+DCf4
ghdgVfqP1q6ulYWVCQrQzDYk9xKADETO4/IJshJpmWIQI+NSAOXo2RnXaFTmwl67
qXumaOH+j7338yO68a+Til1nYbQRkGDFq0bkqf8UJl7pqmTGt1/5W6NTCs9HljLc
p3/hqQwcACZALp4KeRaunxoCiNzwyV4svOJxiHY5fLVnjMCtqfe0vYf56KRez9cq
qb20NK4VzddByzx6hYgSXo60Oy0ABEAGBhEd+LEOL7VgIlZ5/6uCLN6tueBka+2C
TdNjipt2jnwfhBIoBP8E0G8dzFsSMThAwHH7XmY3UC24Mytu8obwkyFv/7abTChR
W2xWvmrNUHqw5NJBBeVBBrdipGk74WQeR+1BNg9GSsBcJ5/bNkCnuqlxgujudtYz
rCk4yDpKcB1WlsWHmML4/6BYiPaxgxvG9FeVdywkObXzDsEIiTUkqqGy0oxMCrQ4
mBaGys3bTpoAuuwQ2o1rL1cG2mEhHrpLnHYp1khAZTsPiPJ9+tLsp/iD0sjPWg9M
VFDQSvXZtEosENUDQZFfTWjg+8uZFdptuUrc+7Un1jKS7lUt1dgrTQwpn7kh3Akh
wscJTxEKkw0ff0uAtAI4RyWx4DtCsyya/9hIwwlFnwdl1P3x4WEm4BH8NfFglzrj
quQokHo3xPdGN5BCtCwTitLR0G1ivFvA8ZHLZ9z4Ul/hcl3f2E1X15sBVTrCSNrM
ld0RZG0B0Ttxle7x7mb7Dvx0I2tPiuRspHceEAjXB/8lDDeF/KbFpza/NLsocc35
HL3Sfgx3idEPsefxP3mWk5wfwR8cDXNerW8mHAPvT3BB4IGy5zGyeAq2XaYGSTBZ
sBSGfwMcr6aGng3Kcb00SzvWEYOXDvfOQ2WZgZ15vDZWEha7x3qXTMjhOqmYPFNb
wzhPPhtsajde8aYn8TEXjaNnF3XOZ5IVSreEBvQZpbJDzd7ISbo9UhMM3O8uIEnK
aLWYsEMcYDOfpFo5fLmh4+3WIPvtbrnsKvF3fljKg6woB80jLCLfliQk9pKqC00s
aO9AAntcjiDzqDANhw6NNNH+4TRJdLy+vwsJl8gRc990L3Y848ro0TmWYxcs/xPM
VxaymcQEBHQT5f/z2zRNJGCFNZ09GKQVi792/Kaq2+niAG09IG17KZD5Mq5dmGyu
BA0vzjvuHlpJ4sU05kC+qxEeyWQaZcuFQVARu5Cn/UYa8ov9xbcNSrj2OXr4f6xj
3nTd7TpsRb83ySZdL864Nx4592eDgAtqZVFZ4fTUAANzZQ6BYhMcwwOsfby1M4ZX
bbANZFjr7cbXane3NOfA57o/A6k2h1aeKTUTAEkGcy3fbltA4vO3c9vOf/ku4eoe
7jSivvVo9JIe741CYM6jaCWNjRvvoqybY90zTrvFbnwir0DFZdf7z3DbAjpuTk5E
8jqHfn9oD2vqOFBf83dyyBM43cI6P6/RNHSK1Q+NK45JKKiH3tVlMuiS0iEMlgC0
0paWzm5Tyjl2zWSRjHOeIU8JrqVbdcQL0WbfyFjKLY/yFK4BusEIOS32N9tjPqkc
daXiRAM6Hy3Of0LZtyn9Dbp+5PXwUqMXmgnSdz63mvHXGgkq/yr5/ADmxEjALJvo
7SNKax5YxSafsmrulyWR+tJFK0K/oRwQ/bl+RNRRSAy08WkI3dSe4+TvhU20XnPp
WLZrfMVWUuHumuEmXjvJwBYEWhaiPxiuUPUsDqTEXGTv4kBNbfXVKpOst9QKGeMh
UI9T2UlEsAZe8XMoWrpbWUFwPe+UAtZmjhhsHlkLi+/TTRQWMM2ZvODwiszvTQ3k
KWUJzvNbs02UklU7bIaOfJxw+yCcxP4IU3kTDAZ5R92SedyZcMatmgcyArHhwaxN
ipTWL3nuCEyJhgXAJe8yKUGanL5uwDh6VyG6PF/DxUa5ajEzyINIMc/EV0fpMyw+
f5lmNdoJ6UTErnw9KO6lUGYrd6vncD/akfjrOsnnFlqClKRlzcJqOTdAG8x7uDQH
UpqOmTk5xLyWi2a/zSnyCY3FNUsuKO5Ib/a3FwFrWVDeNWu+zTsJO3FQfOmTYnCk
W0bEjQqlomz2TLvnaE4AnSzL5KjstTPg9/dxdGsqn561Aa2Q4/v8oQsD+B1Aix5B
82mpUZoKcAGYEK8ZGwcSA2jMILoNV13ai4HlE2TJYEvqffSk6SBrQ1oduIQyA9gs
4ptxxTykxeITHVe8rN7oEllHNGpuePZlTLdCF98z3vZ8KDp6MEYiaIbAq3voU4Yl
CO2t4TKLCbZIYjmfKcu9ytbGkJ+8v3ZWvRhXZXzKcJXwZvU2C5tJyPQRQQjlfpKQ
+gzJAk4YivhyUWFAxFqgdTR8KWEevNCfzxU/KBxBLt/xMoshoZ+EutLt1u6Tyk0S
K32Ao9J9BNQsQJtRaxXudZrxdA1PMC7OZAdmBWmgYjEzs19DMaNa9F5eokPUdMjp
SytQenoBZgDCYPSpM+a5uWCAXmkNrBKxPmRhPMS8o3y5f0mgaCmcQfv/70eOrBq1
6vsWs9i+HD85EIVomd4Dn8iUUtBZuBLIX4iBWe0bwS2eLX9iI7Ovc5DIh8H2bCtS
kzE94EgYdIeeG5hnVUikXByNdu7QKLgUbUdbeAFbveHinguOqFtFwWdrbg1ZWQKJ
SiPeV86DJaYg4jwX0cqAwWb0mU7EyqRzLBt24npuTG1PBpCNVppRD+8Je28cCjgy
uV/6AB4mjIpI1DTJtYb1NSGqYgmXxoyI5PzaJ83coDid+WKU5Tr588E1L4LAFQuR
Cp2vX5XLrozvReJiQmkCUP0rmo3zXgWBIXoIWB9pQELF3m6YhgxJT+0kRWbTZ8tb
2L0Pl+tIP8sEOlejn3Q64SFp/mpBpiZpjDyY9Ug+fo4HGp48/UUht153HgSOpxGd
9FHohN6edamyf4Fe0Td/1q6nwM5lgzh1mGZGBKJJo+GUh3su2TbcAPnD6gx2VcjS
lf+m4VDIMcZ9iVXMfq70DPAv/EvhH1qd7JQgM8JbaWyfCScngO4vHHHdEOe5eYls
4ySIkOoVqZlgpzYjJlB5vcoUNTYcNzZPe3zsYs1FV/n2mnP9EU3Mxa+vUQokXOXO
kODIWZPY2B34rTBbHV3eCUai7rlZlybo67LnuVBJj/Rv+I1ZCRTlzuBgMvwFQZ0u
X5COEbyp1sYh7uXf9zY863EnJFleFFI4GlGw2q/hpYhf5y5bXQGlxw6X0sn5ONZY
baofGBztOHuWPUT+pAuj7LRtgZ2IiOobJBAmtj1GH5fNr4HB2H4ID/MhK0s8EV3w
RII8X3aGl665YqPUg6kTaRjhItI/rCWzPXW2FvRM9p6UbyblhYZOWIyFjDBfj4V5
bBExiV0c4A8VWWbYquvjbBlb5KzrcLsiCV18RcM8mXoJLKe8DEXMNQ2XySYpldmV
XIm9xPNTvurqf2yr8T3weEw15SUk0v/j9MgnSwJqb6VaKVqtgul7GEfE0ytiiPP9
29IWdVgcQUU4cgSPAJbKqIs2REjWKZsHtXifahzhWaSZWTL/F6UpaYiMcN1dsv/q
cA4o685TeIo1qZjT2TssdmCqtHZB+AsmSON2nkevEOqBUgvLv7tkjVy105/LfX6P
vr8eBv+x36bKQOnGm4dpkEJUtfLRoliclz4SuWtPK+otOXfRDCy43rBpwMMf3WY6
R82GxyqrQ81hJ/GoiOASkNidBCwEaPFb83BPpQ8fnquWr0SnKMOYwbGB+eAAlBlT
RiB5aiV2s1XNqvsnGKmbAlyHB9mziUYc0sDLoC5hHYf/ReUOb5eDIIBBTB0xDv+t
hmkoiSbeZkmnmz5VbNB3B1AFsrIbkdyAoNYrtUFssz0hjG9dMADEnSDbND2uxGGM
goTnuQpZuc6bLUG5MW8GZZFNFDvzYpoI3a5iyLL617ZB9j9UxaGLXrHkPtHDlbw9
m2D+GVxK1GSav073SmGYpPdE1sygH6m7HgpHpS4EpfXn/thiIAO49ywzZI6T5AMs
7FSp0mIIeYj6CBvKrc3iHZZHd4QFkAeqh/9HkCkFtQniWw5SiS4uJlqRsYqT/CK4
GshAveX7NHkzeBlsX/pjtlvwitvVEg2lNhWQFYnp97bUJQ2zXtc4gQxkldLk2WaA
8sY5RvF8YE9cBxM0kIvD65loYEGiNP3wYEuQprkIMTrEjxt63i64WgIcixs16D1x
ku4Rb9v+8Nwi4snnoR7XkNAVsKv8xJL54SOT4d1jDkLoCI2JCM/TeUPbeLAoCd9u
clgSD27VX06hfKUIsr6mVEbUyXenxGnwdrd56umO02M4gMhPLL77OF3XqXy+NeOH
u6fDNiNWEmiVfomk2GTKw27dUcu59mnKZ6DQ8i2t0sgaT6PHcahE1EoAvq4K6tvC
fLaCFj2Bkiz63wRYC0W6E0tLZD7OY1vBbvdA1XpwXBo/hqVwG4gS+ofNFu9eySNV
hTDoPFsG6kR3nPEv1kIcyAeBBp2ST+txwRBlDXNmX/puX//te/VkmI+dkuK7UHCl
8Ozrj0nHg88VlN2pVG382/VjZc60Jg0HXPnO4t7W+Oa4FbjWOk2T0fWRyZl15IOI
wUuMI2JDP2J0RnXsqzqEs4CzxPwI4E4birxoO+DRzaOsALF+f25Z6ximDP8iQiL4
OmE2OmsipPTNQ2IDsrcj0KGJb+1ty+5KHEfNdWC1fembyxPUYkG65DjdTdZcvIJv
v5YQ39dqlsJnnZD8Aw0UYWfApWu4V1uDV2sURfybqRbGeUMm5F6nLNTs24SwimHq
Av4bgI4w0746NJXQ7c2XBIMwnpspJeN2uP5ttCgUp7jNbgtSVvt5iBAfmOKhBFQy
slTP+pMvM01XtLtOQ6Rgu02cWIFMq/eMqBndQbXfSupV6KaHEM316qy4BvLhzgmB
FUurR+gw5JGvQWEeCecDuejnPvSV1By+ClvzlmWA7fQN6VGVoe2eF9vQvkjl4NEE
TiFNJvoL5N6jbkfODoLQWnNlmUlBVVlRLLUbMwe9FQUUaTukNLMePNJzliuniYac
WbuZuyaYWMHzcdFrFPNXVjkI0sugFDYVGIUDT0n6Mk/SJmnJQFoXXYYNrSEh5S3d
XdA3NKpRbGSaSX/FVGMCdFPJuEVUZvVpJ9NeJwcUhkzgx2E++q/si7nHnOrPqRnL
x+t0n+SFNkasV86D1ulX9xGx0kmtHkgPhJvPqI+PeKTv/XT+XXQoigQtxD8Q1wZ9
owGZl59m+BXWiyGhuRzzjh2/MT+56ktAsmVVbqjQ0Lig+gisMVsjMhQ8I0Idwhyj
zNAFfL08YQ6plbyRPzbr8hJ03xllCkYNro/2iEYE822TbxfY2qgaDLLY8kwe2vfM
kadVoEi9o7TZIIdtQGYoazP+2kf5ZGgtxmJnYrp1gU2VlFpSVEh0LeH1VYu1vsbx
q/C0vafxfjWUT2vWw7aoN5nbG7jGZPZ3TiRJuiKDuvtc8WmPpl/CtMBs4BvjSTFE
hkkfTivHY6o6ReaJ7i9/hxqYNxoGp4J/VV7Yod7lisTFEYTixNrhuRoiP/B3Xdbh
fJWN1K362LRn5RzyfdRgCKeFVqH+/c/TzM4MQw41NAl1Q3L5zYK+0tPGdDSHRTOu
E4j4r3Kc8msvky5gRvseIHJDdJlk870rWtHEkw6/Z5NZd5Xcejw12PDL/1bs+wYs
8B5gso4Ci8hWx7xzWkuj2Lh3M717szHHmI3VeLlSWW0wZgdnTPaVPpbJ3KpYY8yF
7FB2RghxdWYHuk4/B2GvBPhytgY/74+0YqhA8IhLYbPEjJGwX1UYMgy8BTanbWjF
8BeUR1h5f/y3gOoMRSBYXoPzvpAyes/EdXjHlnHr3ld1B4AthHEu7gxeNOJLFDdX
iADtZkK7uf1Ik+qRC9K1BW0OxfOXBKpa8AeipXYMEC5kHOwpr/8p1KOoYr+U7qYE
CFUVJVr/WmPRnIPiK+RawgtpV+cO2t6VYKQi/8GeTN8kfkTuR5Zq3KikMTbLdsLA
QkE9OzV/ylwGOUrYeD5lb5zErnSX0jRJu227pJLGp25/Y3WQU7hT2aAIZkcjKWJ2
iSQx46FZpPwvPeh+OH8rMf6i7FkDph1ikaBvbShGroRWv7bOirBQTqIl1eHbNQn2
DydPM9Cq2EIct5vSWipph7DJ+cNXG7ANEUDQiAVDvggcpO1wbGEa0PBntsgnCUS4
Yjn1lzDc3JgkiubowzpZX8/jq2bFuP/0pWfEnC3jVh7rQtPPWSjukAE3+G9lkZU8
Z76K5TC9pddcHoumtAf9CZG8he2gBY+JjvQjUu6f+neIJi4vtfj0oPAhB4AgEELN
h+lFIQ/FfrGMbuOfBBuo0l0UcjRcurvak3rDmcy9pO/MHyz1OdcvGNadCEBVihZT
OfdPiHTyarVni6A2vGUV1kshfxx9uCYns98NcgH620LkBfVQQ9mGMI/IXfF1j5wQ
Jwzou+z8ZU/n1fdh7H2S3+/NeU/8Pcpp+t0Ek4zydPvCR9tqefszP1SsDaD+N7Jq
Zb1U4ttuQJDnJzI0Dc5dwU8iMbNxUewreZ1G/49OqLEbw+SSK1T+BBEF39vlCPYf
ckc7F78UGGqsKfL9IugckDoThW2zkgsNVnpYirZWr50lcxJXt7oxFoC6Os4qxQeh
b+ZpdtZKqyGVkiLDDeMYbmc6N3+VpuI6zisGdsPYM/57ydn+gLvFt7rf3hAEwB2E
oY4ob6i7JIvfXsN9j4AHy9d46vHU2YJhm1GD4BcDZfRIEN7Bm+dBkb+SzTcgUbiw
98hTfZYFG0gkt46QavwGa6LxIu9YY1rH6J4ohZXHghmjplAPRslvR/BDOc2GLKUM
jFpsTtmC6G3jDbKXy64fxrAQR2VrU+tbCGwToEZZtnsQrT2G5Lrzsi7zvZf2+UlI
o/CUBe4NCepMiLnGSrnU5eYKLUOmzaGWSPSpeJ5utMCqFAsDcIVbJC71psQy+8t+
AKV//+0ZrMgFzzT+zdOxaDjxsLqMuAYZy5vwSnfgOZGSotOtbwRMTBYeYd9QK9me
/eKXDpvPkiGw6QvR+JTXkxaBrS2n5/I6ZC9W4lDcoY8GvuKKtYnuQRvbhQBkiDTt
5FTtKZgaHh5DeSt+/4wzyqLyboqrzX2Js5H9ZQ/HrRoSPxtZuL892HBBKf9xbk7N
Vow+WuaItejSzvdN2w3R1OBqEScJSuckZrDU2nzXnfCUjXiHYhCukHcVOKQnDwYM
Y+Qe4DXi6j0qAqEeU95InThZ5Vy5zB6qTFGUq/NJzODOTVd6+Is5p0LowdWJaGRu
RpCE2QVbcDzKzqCWAZdPaFzDc3bfQ/eFGJzWyGXUKpe0+uzr4WvUzYjyKHhhdbDf
+CNizW23RFPeCUo33W9reWndHzHZTt+bio+ubyYdzvVbimX5CTjUXiAegS9oxiGR
M1mnz6k5oe0osmDFXjXYDQyG5pngLOf7F3Wvq2JyTp/QRqxQ9w2jrsolYKu+nZxh
TgxKfIx1hWEQNhM6WVlt7tgm+Y/OaCSv2FuHGJwaO45abM54Wqkm+LzUDFHCoxe5
Wz1+TMhYPOyjveMFNyiLA+sInRTFOAM1rUPU8KTzkxkFQH+cDbhHENVZkN9Zs3NN
I/qfeE028y52lP3C5hcGrw7QGgj6lb6DArlVN/Tzv9JwRamOnOYGWhUXce/QqnDw
nuBMexjMJe+WxMyWeCdDYEwGvw6Vmum4UzOX4yK1vgI9zPb7JkPBG/AFFKjw2WxR
9+ve8JpQ2hRbw4vCYNHYAGXxvFR19IVcN+GI7yGmt88R/YPuEy2q8xltd0QFneIC
OtMxaE5Xb5FV6w44v539tR/L5wpR9iKZcUMQ995RLYbQw4nRNC7kZxJ0Ol/jsM/i
4JVHb0PWtL7s//lRFqfvo50w8BgYMzBcmv1uCeHWwkXmC72Fphf2BpGVBLeV3yxR
JnKviswcBRPX7DN4rlrMr9ALhfPG3B6hqp6fz+ZYkqUwGFdzXtxOhCn271TXQdn9
aAdPBn7wdxlMMQUDdkUdHqb5IK5UXn/cqHZoKahZljLMHXM01yaOPMVziG3hCj0m
83IbHIh3xFQ3hCD/O725FybAJjvc50O/mL+ckzRH/4YsBq68iE1qn/nF1dV+to4G
qRP2GfqiD2zM+CZ+U09kU6TFGN4wVlNe5nEEA+3uao+FgHr/CjzJldZecE1DQpup
CUugJXNvJMDS4+PzT304J1i7e1nww62Sz/aJdQIJK4aNJFnRXM4AukC5vLWtiAfE
c7of131d1StdWRNNhR12vI+tHCcuswW1xuLVzQHXNSXbQ14r+AmBvl/Nm3gyNihs
vVQRg0KrFzGANiwFhVamxPfHa9za+MfApKgbz3Dk73PZbc1u7luj5HWOOuIeGThQ
NKSDoJIFVDlsEsTfjU1UQ5sR4NTXDWbiyDhYD/fCZZo8g8xxFRTr8AAgEhIYg0Z6
s2GPjQOEXMviwYbUQw+1W77IGHd7gQfOt6e9EGAf2u4Gfq/AIrPY8+9iASeThj12
mx6A5qp0jv+n9YJf/6ecPkE/72ujUlEo8GEd6TQWAK2CJFD7bxSmq6lSwZYYZSoQ
CJjblN5FLrOShTL7eHZiY9EhNSk9eQT7bsFblLouMcqJr4nxf0xl3Xv4nWvLewCi
CSLNpm3QHlojKc84DQQXW9EG5e44ReYIilZQqgX/RvwzZbMw1FQrj/H/T+GCIgCX
NeVoBx9rELymevMnioe2Qu4p2VSLVmlrh4HI+L8O5AGA2ibUL62I8X/LVQ5n5uZ0
SkG07VAVT6uiQMZYRBzLKzh5xEbt75DYRrfqjSoAriS48x8braBCNGZnGuB0yvJV
qkg3ZN3esLwr/1t+NoFG9QynO6zSNvVCeFrbTQzNZWCEiaJ2CA3NnJn2SPKfs3vV
K4Y3UEprbyZoN4JpgY/VwMBnlbTmhzPNez7BqgQbR9sPH0kkBrGiQnJRNul8j6fJ
lhIr31QeksDUrtreCBNUlHD2N6cDO/G/4LIGrIiapoxLiH9Rs2c4LMoVMybcPbLu
0VFEU3QDST8Xtu6AOBXyMQuNXx66YC0NIdluBsN9nCCiEsCv8WqCon3YTjY0laoy
kdSahoTVpLwAQt2y/zW+W3hnsWaxkd5V+Jik0SHo5ojh8kO766oCuFhHqc3XZlgG
Jqrbx0ipWlL2I/zSUXh2F7MvofY6A23/qftlaOVZOHSICgDChC5WG2TkfJ0SF687
4jV1EE85emQnTIX7AS3v9NBmEOyJ8Zspiep7NAJLAw3QuVQbSPzT/YaXA73zcSh7
o1G76DD1XbWU9E0Xy2kaOpumIcOxe3515fR8neQCyzBNO+HwrxBbB3aYA6QfTFBu
svx6y8BEfep/mc2uhNakJ0GjpH2riaWVTQwpmzY5xxRkiMYKn633RVP6x4Jl0Qx1
T0eG9boi9nHnIr1jn+sjgOnPgI86hfG4tID5RDKWr1/IZb82afGUMk6mWX4urzVs
ifJk7DZXLOpsT/hQS9NCD0DLOcchfzXZP4G5embXz/CBuAcedKlVkn4xAz1S60El
JHvHPY9nUL9bw2v7LURVILbCFTaOuG+d5jp6Tutd4nzbXLYK5Iu2eE86CZpXkGKf
8AcGUf7rSVp5KtZuKHevjfATzNjupFXflJVJK2VQp3x/lqR4JeawzopOL8dfZfjO
MbU65F8YA5ysUHbvjlAzkN92RQlS8+oqf7TDlsxoGAGjng5N+QKCYbXXJGBIA4Js
bzgkAy/l4erbb2DTNFtdgRpEnqZ4JjKQo8kCMJHSxrtKIgrS9wsO8vsfL8FigKfH
/WqrEMNeIedu+ICOJm8SO9hxXbxSoT+70+PNSTYCa/+Oe/145BHOYbghFJ3e40MU
p3Z1FLE0THOfMez/qKaPa2o09aJ0FZbJXYLTtlpRxqO2zewd8ezsCoJh9FktlTMX
Q1VR+vxAlG4ip4dHiAN4F72LHbByEfe72+bViDcxzKQ=
`protect END_PROTECTED
