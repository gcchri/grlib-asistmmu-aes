`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7FG4R2p98kWYA2av4iXfKbcaVnqBRaz+kqU7idc/gwSSMehKalMIBOI6RQrNi0qt
QUzUccWJjTQgt6tmPQfJENStaFEi4tSuMtZeTvDvgGEqdKBCmObxyoQmQB4TguIb
6oyXnWEJRf0GsFHsr81CV+zBgkirbcd9PrEiPcyHIbvK8fbmrW+YytEtvHPSawEA
Cgr9kDic+5FqtJRDFBy6oPaQvzkZGFIXAHOwT/sGeXp8+Especu+MT0yYKFyEPvg
ylto56COtUCC0++ILlg9MrybEgpvNUrJ1rqNqi5AKQ+lvJYN6TyKQts2KVYSMKgp
cXxf7iRP8oNfY/ujv2q8St3q0PrbKxeufuVxv0ljxQuA9sIqf/F+bESnIcYEwTls
+/qJgztsSNvmxkHsK0gh6g==
`protect END_PROTECTED
