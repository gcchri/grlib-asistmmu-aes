`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bFgtysMT+N4x1IZCzFxMR4wdJSQk2iRl9VRt4YZ1R1SzSXLRMokNFhE/wtcROaZj
s+nuhuwZNveDLsyvbwHNqh0KkLhY5genICLb+Bdpi7O37rCjPCfHz50lz1vKHOhM
vU7vJDXTUM7lomjkYjCgPcHtMQP00xXsZ5tedE6N0DV49YkUFSdW4TH1Bfd1T5D5
dXyXtPjdpeaGQffrBn6t5SQYaC1c/M2exGIFqzMBDtvUK+7kHpddkKIQiiwzH3Rt
PV/dRD+hRmpk5lSeMWAvOjA6AC2ou87xCmngIVzEaUmbbotgtX5QR2GYWc+bbLMG
zvHWhatL06IzvHrtlm3N7Ul/etSLt1cl3n6AOanvwFL40YZyqwpTj14Pwh5SNJtT
rddwz+i09uA8UguFo1Hy6fPDPFjowwjjQI3J8otJssY=
`protect END_PROTECTED
