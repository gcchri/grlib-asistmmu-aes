`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Xw3FMMl+FCecJWyTk+hiwnPcbq1DojKtmX9rWg7jdAIWE54dKR6Dtk7UARwlrOc
ViBl5kYeO6t2Lr5ynq8RSD/QwbX7fpH5NsGVRqCNpwaufLCnpMp5I3MmcmwDgUFY
4aP0LUefA0mAf6UKlmOQC0aIMVIeXmi37DTsyVvlbSdG4jcwNa/9iLesQ6cze0n/
DTJl6VnvsW4e8dGQRke0MY6ojdiw/ZURh1jmtQtSCrKqr7L83dmFbKioYfdgWvQU
PCvHMwQZIVxxR55sHLJ4T0sn40tapFZFIK8yXb/WoEl9rBu081lOh21RoAiI+na2
k39mLG4In7n0TxJdcYkrY+UZr80iuXq1L92d8mfVv2UcGT5C7cJ570IKpNjroCRI
0u0ZiyM28iRAhCulOUkgXw==
`protect END_PROTECTED
