`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5o2P3fT+IW76JyQ6GBFhWS4o3QuyINGi1jzVLFBFUIW+GcOGNCj86AwCsw59hjj0
7VhbdJoM/92PYlyg6CI37eAmeTC27XbZ49mg0LMzyr4gG5IjenuPadx375WELnPy
ruMAPHl4srePxHIKg08UIT3f0N5klZDfNGiX64Q6jEnlh433X+lJzntfDjw+UnTn
nYDo0myHYGYCevUqZmeVFPkrkzVvensOhrNB94AOPezPBt2S55uXKomXbvMoNMVA
G+SGpDHogR0e1nRcBZ9/uJ0iwXVeW7HCVWhnAMVq0qyVAWi00qrC19NR/yvfo7YV
1Kgpin/tZUpBEIXQE0PejNV7oZrxycy5ouyh2Yb1Qtmo6DxAj5yQBiPuMJ/m1EQD
2RKoSjlH2uLwI4Vc9MYS7Zft2+c+9g4XoCwAVMiK9z4tkEYsId7LFJNQ9XKpaOMh
`protect END_PROTECTED
