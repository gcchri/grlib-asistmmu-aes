`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o6XV4HMkAjeDOPr9aBqaV/FeayY+JPQx4VCpJuArvH9uu0l0SaQmHxqELqCtO9vZ
2pFEkUXSOMM8SEPoGi0G+Z/uAYui4KnOgwk5A3EpZSgYmDBrTdCxaCu0Qqwt6nnq
clKagOJbEtz9IQo3/4OJinvWA/svl6dBmNgaDZTcbuXAxoFqW3PM5mlsKjbI4dws
pky+lPBaOu0JkgpNaNZ5ZtdyvT5UcDZqmKRTQxPLD6hBXbucnLgNSHSll1+RXD2D
u+awWWw0UKyqQkf/cZxb3MX7ia/fRLERYXWcmmoo7gfI5MdFkaNFIkwRYtm4cX/Y
/5Qr+ByzfotLwAhN3nrpkuGsL0EtHsn2oL+fK7dJl5bWhiYow5b4V/jY5CpWGkrQ
gNzjIu/uAE4OIlKUuBhncPteQVk0XZa4lyG+Gz3FxnhU5ogIsgNAD/97s4vWr9WI
36JxxfQmV0urXY0twqWwik10euuXBmRZVnS8KXE3ZI7BKjIjYScPYAsAaeXBV6AV
4CsCECvdMP7UaFokgyooO+CZu/oKapOTFsfnnKX9tpNyuEtwcCZgwd9M9yHUAmYV
iPXsEfcQKS0CH60BKrPT8NwVh666XIIsrjh+XdyJqKp5AVHcALyxOfh+5sfc4Pjd
Gkl9317l/WVpx6vMX/WFN6QiS1fxMuT51MbhgtEfAAf4pwlC/O/w1FAfz0ZejGkB
lvyzlNgVnPKtaw78Ak170+F8xFssLo10mHz6LrYy2cHCtEt5hNW6T+bOGdVxkB5B
J60QcLYGSxCZdj1+WG84YV8/1xtCKlw/d3X2Fi+ngrVOocvpzo1nZRUea3WyizJC
mqrc31j8Q53Hvb3vV1yd8/llOFxJADMNLOE+njGMb+UB5XYwn1+AOSZVPPjjLhRW
SFUDJZnUWOduOgQaJcs5CCfRvUFeJTeEFBvv26f0UNiVzHYaGn9cHzhBo48eeigX
eOxaJnUm5o24NJ/hawZG0MX+arVG/K0eJhEDWOyd+tvR+I9ZpO1jrJuZu0ONcuoF
52XkDnOxxWy8fqbc67XgnFn6Qe1yja7Iq3K95eSfA5BOZnbKMf27pc1Pu16Kg6PU
6TePF9PF1TI4O62f0WzA8gf3F27Yl5nSl7GtTvJ4IxsLGkwT/cvFJwE3LM4jXbeu
AYr+zviAozemBYMQbe8TR8Couhk1uMGq5pLiuhUvyv1m42qCCk6iSXAEWb2q82xP
OtNLU+ge0GmLfUw7Vqd8HovMcxQuOKI0j5u3sYFy7FTQwnTVEYht0jucVTVUsSTV
k7ZAJLdCPwxvr0Df7zSxisDHbfFW/BIhrdxWzgzr/aiA3diNsTWnPEsVLDGvNhjQ
5TCTzhn4QIy2C621Y51HC+YkAnR7jz+V11k8WOYj2l/ArdE4lK6ZQMnrAGSlJtLW
aeziboaFzqfd8RwuEfbbVoiXwQbZM8Z06sdwh2fLERcU3rD7iyifEKmMoEToXS9X
yK/rs6HVeNp/mSCgqr0uTWLnx9xqXKlAJuGerw9f6iiML1oPNrisxlcix3wv0InT
Af9DiBdapV8LyuYGayKL/8K4Fh7CGjvwrdVdbcT951KhbpWoxI/6jeZZ2z5tSOtd
LfMnND7zCrq2L6ad77rE/eMpt+azKf4UE6mUmRX2bvlHwf5jradx+NKtrjbPJwRk
aI498//sLshRapbjdne0r4kFajXcq37G3kFKURMlo3CyFKAReARJ0He9vW0zgRBZ
K2AiBX30fskmJj19ZubR0vpU5IWnmY6dHPXunSZSiEC4IQMsIhCcgxH3Mb76q6tm
PPM7Y8gKr5lg7eyVpqitkgeHIV/koCT2qzxcKLbh+3+849NOoiHvT2ri0Z4xkpmj
jQfXvq6jKu2oMaFag19bOcQ3mzxs8LYC/cDIXqKZVH3QsTuzwXyOxunnOJ4z8Xov
nT0smUatBc+PeR5LqYv2rtUPLuAU/LyPL7D371E0SdU1pAlAyfVJRAV+TVufPFtI
r/wmiOl+FN0wfmVU7rvaK+UBYKT/GRe6Ky93zOSJ+B13bDf7ZwExzhjDDdn2XKuk
oJ+3ZkEB/Dr0VhzBayz6DE3jAZRoy6q8X4PondWJxcXMlLC2qAJYGUm68sOBBRoI
/v+fuOfR3cqy9hcne3Wh7egicyTiVfu73UBnDKYxb0/YO/q7V3X97NCZVoC5Awln
AbdPVXiJ/q44GrnpafsGtrxGpyPxHKI0TZfb/f4cypoWwoL5xUEGKojB3FvXDb8K
5GdTXTddDYWhbcb01MSUzkO6g3stEuF3or6I3VA3R2ATVAoC9eIOiRrhTlxTQVoQ
lv9PeCnpTV3Ih4RsprhjLf+eueHv3l0uTFpzJ7HefuO8709kN3BfxEG+5xBNw06X
z1+tZ70ryJhNVF8Y8B4L7cgyyWnKtBNwLgyCuCM5e7Pv3bYqtp09AfcHVv9Rft8C
j22BH3G9YcFbKIHeIu9Yj+D5MC6jvJ9X21yQ60eAs7dzO9ylWsY02L7NKDpEnT9Z
COuAuRQWL2Jn9p7SHnSMDe8XDEJT8BUdFZgKqMK4DSGJtBAx32XC2fc320tPQMPj
rOcYzr9MdaC7w4D0yfeM9Q==
`protect END_PROTECTED
