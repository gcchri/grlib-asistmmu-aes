`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YH1Ntco7BGcjiVGWk10wW4JSg1zVBZosI91WMi7K83lv8dc1lAMY4Oxn5zSqUQT5
gK3BiRPIwebIQ5CS0LmRFxw0dx5yfzFhrH75sAlQOwzfYhW2fnTO5LieHdT5fM6c
uficYKeva9xyE9G9PNLmYhWRO7iXm9qvcG3InbRw3DmT2Ezbs/z9ufM7E4u0JGMn
+PFC7MJM9uSSWw86rERCuFUL9a2d8vmObkWzp89qtqmsGNVaN2xdIsmMCfEh8lsi
X2r47WQIVa7EDVrAVRxejz/v5KpKp7V4R1dwusqB1JLWMoLyQPB/HRJkSt1BGkVO
2UtedjXxGNCX/7jyajsUxFnTvDSfd55VyOkJPV3/Lf5ODsLiF1jyTnngL0oVpVQZ
Z5r5u/SEw8e+A18X10QONSqahRGGTSuyo/2rFg9LOvkiNFqpxVSOeOj39iJ+cooz
Yxlp7m59FINWNQqprhvjfgRFLhFyxVvJPsXnodeJCO09J9C8BIiqbMGy5OxsICms
jS/bMsiigFYaE327sxiqxBuTDt/NX76Kpg8alA3kkzW45Yj4SIsDp00WmEbA9knp
IY9WWUlGMb5D/1VL1+3dPN/EXIDLlz1MrvV2QRFGa9rRFBAhzuuHZmKks08JxR9T
PclKf0DTZoDHaoKAfbvOcQ==
`protect END_PROTECTED
