`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
46uljIWFgMI+ztpIgRHMjlcpYXiiLwXYN7N8lGb96a15PUusxHdqO/n0VdE2c21J
Ytz+kkWGQHwuZ8nZhVTpWducYHQ6R+fhorqWJMWh2jeglhcFo6Y1TvIabbQojF5h
/wf7RYAv2cMGIkk5UwRrW74ME4X9XmYTXnP77Py7YQ41viKO0N0SmfX6DRSg1izy
SZqssQC+XkVSZ3MhU2qiwkfu4Xe0/kYkZc7uRoC2N+Iz/rdK441LP0RXRq9UhEAL
AEYkD2Jm/FKHt+vdeCVqaWXC+L3Dq1XcfSdfAK0AZVLyi4ROM04MKjm4Hys67Bbx
QTTOB4aP4KgZFhnmycEw3lzLsQdGvUQ9Lyo4kJkukxw6D7v8e2vUDo+oeeXZGJA0
lTz6y+7h+TLE5kge+BSHrnb22C/K4KXLlRvXicj/2lV51zSmwcQjI9bwUcD18ESS
vHcOmaQjBRaJp5sNH+ORuygMMLf84qCNIBAGLnsp1Hlq0fmg93T1SxWTC6+UCmPS
JUMPkQpS6BvF4PubSwPnyvHINxDPLIQN31mNkZ4hy8+HplIF7GOCYzkgzWTm9Goc
5MBuh9O1NF15PZx/5hgw7340GQdrqDiWkb1E0RTERpEDnpdxfOWkHXPnucvyFIxT
LHDWfS08smnn4Uu3bCdBB+Zbh865pEAtBbSkpJc5JNRWktOjj86FHpAnERuujdPO
Oiiw5DBZNa7pbQbPOSIn7rgXtfKTLNsqeaTiJ6Hf8b27qeWIkTZBsOKmxxLPxwEY
PJ8yonVqy8PwA4S5LiSGqYkLTxH5go4+VN5/z+y++/HQQGOHhQ9zQY0Y9hA8TTRz
5wZ/B6sOr86J4cxlKdHn1lllDCrK2O0/2lIH4/1F9ACLTeV6P/VYb1ce0LmgMXJL
EXcRtS2L3dh/K8ATEduV1JVwHOinzcyqyIkx7Q3Ggacpnl1tDDgVLpOyKiEIiJ7p
qx1DoymwdvJrksX8Ciy0wRz0Gq9RAnvOfLnwMWivt+PcyZxPKZD+glwnMYjT/7J+
VCVmO+Ul4KlggqmCSP+HqWtxKBW9qx9PpfR/oayLZhbTFwNHDmgZbW7gzXi3eItA
Wq7NLMjelnPGwqXp3XY172hDXwVBSylotyOySpcwLPiTQxUKtc+GzWh/lWY+HslN
oJLlx+KppwZom3cOGMDKfrbNLm1xjkGp+Nbm6spg77SV84ffQPd3vpmjkkO4n517
OT899Odzcs14h71EVwiDIoWrGuyye/la/fsSaQUA8zg8Vl6FS6VWZ1pI5OQ3vGOF
KN3kcz6yxMkJQ/tjOWUOqFAdymmOEZnOmtdt3rOLGIkKfVE43T1vuDSeGYbyLm8J
h8wajYT0B4CTk2lrgpQJLt14+do0IO1tTVxJzH10cNT1gxtzp7yIz0wlXGdUdTmz
73YauiY8Cg9HhwAZBtHWCACA6GbOIT7shwjngpBaM2SDdrYWHVwxttkfwJD8tJ+m
UyH39gGvKXXoAMCgVoQF6Sem/6gIN8EUvHLL8Kd8/SrVeLjZNfS/fmgJqAKxTeE9
OkxHBDxDIswEpggeORnYSSN2MaYQC7reThEdqGyy7yAqRhuXgAZDnqq/xidxMtQ7
JM29eSRJJmU+VlzM6Mk6i7wxo7yVC+QeHhub7vtmlWjCKw6qxPdMjucfwjcHq0LA
pOUAtJvvhpNCxlajrVY0x944jxIG09JDJIKJ5J0t27nIoK+yrEhanzDc2T9zEZ15
uMd0RE1o1IT/gtOtzFS0W1mexwxm7G0+pmFG/YfW38kcDNryMZ1Ehxq1BqHZwSRC
cXwIk9xRsPbT17Q3x2JQaMHiMu2qfRbv8YT/U/uIwHLHXu3rTgKXHM1UEZulQX1g
xGZczHhl+TWobl88zRiSPaCQs65hkWmXjg1yZYQ8a3/Mdk+qvNxRBE6mjzoJd7IF
Jdn4SJk9kpFvo2VF2rAJc3bVQJV2E5xf2tMmdiHJJP7H/UT26lhPo6r556xHEUQo
p7zws16JMdDPN/ESCyjd/9LEI3cwuTACiH5xMzntykUQ/j73FICSBJgdbS3MLinA
QZAa5oTyOh8ZdGJsSPT0PAAHMoATWIGHtE0GUC5uIKk3t/cPNZAlkVsDrt02vYj6
WVbuw1BRm20TVW7ABfIqdzzfUxYwfuKMUt7daQikvdDoSzL2AwWzEgUOVPzFedlE
cLC2uJODjT2W3ZtorHNbvbWmu4F8sUEGg9XOVz1IIgxG7ageODx8AGiI8XRysK4F
LTJblid8tfMWtvSREzjIhtROvNuAThMd2rDtVnL8Olu+xFmSPdi4DHErqQClDSfX
b3KcnFRcQO3kfEUBb8Ldw2tI6hJ0++KT4CEuiDmpBi3Zb8eL3ROY4SxUrPztkIbL
cI7kARgeMvfXi36vxHsx0PEBr1YgeC/sLqD+AzGvtGfTR6qaTXXkQAw4Wva+1LMd
7Si4M/zpeCUOd8IJfswIYoWXMTZMKsEEHiBdnbE3KkDdRr84ynqRy23F8VsyzTNT
8kz847SLiJuE5qTrB0tEqF0DmCz21Ep7oric8ETtd821rilDlerqYDdVpoS5kAmk
wv3/2zgI+w4gCSJwSak9gV0yDpYDcBgDu1QKrJVs24h8gEEDQzl7wT5fWOAMzpSy
EDcv18g0SxAr6S9/jjMtYyFXvmBBDx8Gc+CXPK7fat61FrDGJvpGXnFP3lenX4uk
KHanassjNjAqsKRUMk8cOPnsbpqMs2Uvs9ZAe0gO+M2Daev3Tx0mVupgBrm3O40U
wM7rrDjvewPjZDymw5DV5hiLcC3fheJBsGxntWDrValZoqSPXBfODYXL+T2byKtb
J4ApuUf335XkRx2W++/LRcGsnty3Wo8voddtoe+5R9+BUHl8oIUjDAZ1u500B80N
fy+tdWxEBfpQ3jqD1YnovocHGYxEdjxAy/FjlIdn0iQToKE4E3XbpDVPmTLCkFUQ
bi6v/u1dMeSZq0fakq2n8+ciMloD9u2oUoFbrKIt/ns3edDtsbufucxSPuAgftKA
k/kq1F1tnlBgq7vjknH9J+PJijv+cqe5n/2HpucUj62vb1YuEcwnZ0HCxM4IaM5H
iGupg7Ft0qcBPGEzmeGznkwMICR1B7QCD0LeDNd+p32GZ7AziPjYsXdHcEqhphAP
GIhM3EyjD9Nlk9B8VRzTLy8n57bKDEaBXM8ip03exMnBAZWD/xI6ZfjP37hfuCK+
ee1PCp1v6ePBnVS0k7RYtLUzz5a8rej/Af5xrIZ2egZzAPlnn1+p5xzz4GxaBffr
ljMvPK8MtlDRqCZWjaPXU5oBedD4aH0PKamUMGDOvxmRQPk5umIBsuE+PF4ObA+G
U6ugUcEfXhiOIQs5LVzM6n2rPWVF8sJFz51f5x6fJWCe2qFly4YosfRNMEGj18c4
Eer1r/i58RwwB2dRAxUD+RcuTSm/Y+8xKNzaPBy4s4eJqqMmQLpumnNqnH1ssQaT
tI+z7Y6roXafMHykVYanf7nlOhu1ipZpq2di8Vhr5TS1xBMoPPmxTe11kJaNQQKa
RLeG3Sm4pvhCgfaToOCi/cdJie44xVIxL/jvNXSrx5/pBb+6N48ZPnXDWhqd6JBr
VYjetx8Lx3CWvWZjxzdO6bFd6a/CG7vsRzCmkE6sDcUMHtAuObSEM64jizKKs8Ad
7ZZ0/KpoIp8b3sqSdToT9zJEfyf+Rgw0vbDiLsV8Utn8cfqbSiCF7+RGsJHgmDSh
9uVBexOhuESCWaika5l8354kNqeaVvs8c+N3hkTK8dnGiQ5qXuvisKrO+vtXjXA2
YAWT6a7rsvK26n5YzWMRd2exkl3kZQxgZY7txu9ljNNZcvlgmtHTh3yHnO1DI64e
pK3oOEsEKhJe7fQmq4tjYLju7OODsa9x0/yuBU+KjBvwFyyrIzdCPcMrqdJkfjUl
nvJ5CqzqHmAMHCDZ25O+rTTbj21EkbQ0Bslrf5pZqEP/+mTcXKdjSnBOkuFUU8Ra
RBAHI2bMoENIJSIyzKHKTi+F6Tsc3qyUwV7uELYqDSuRkurMDviFv13fy+6IUpff
HmcMXELJSG/KdcHime2ippNa5CR3wvjsR3ySFbuj61TXYSHd12+eCPsPJedFG/Nq
S20YneSxlYY4qzxyCd1BVSV3a4UJo/i19JxM1l5F6RDk4YWpTXcnoKuOKpT8499y
cugk9AcwBzlyAqdOuJmKrlyiRkGUeTUHJLrwDJmPaXQml558nAPHgEflRMFcPuUn
y75FHf6lQF07HPjXOT7tQEiPKvurGfpI3SwatuBuvv8=
`protect END_PROTECTED
