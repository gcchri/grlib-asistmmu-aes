`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I1FPm7L9vG0keLGvR+BKJZMVfxV0d+QMWAG9vnLihW9arG5HTIBQ8M2Jpxr59+03
DlnAC21QS6UumkBOufoNLpjQaw1aEf9rr+bVDnij3DtRckFbx4jjLyTBKejG/Dro
xX05ntkgm4PJ84tdCjd256fabR5SzK93iTJdjtwIrYuPdQ1/9bhcvSmxSKNOrevx
TwWUIgC/crZgyIKpQaSJn5dAa/41HfQsT2T3bmUHf3PXA9U+LnrH0ktanqMXWZTL
cwQy+0EirIXuDCrvL6iCaQX2nT738AhzEWtL8KgwbSADhSRBPWipmbWQA4ArFxFK
YGwD9UM/4KX3k5d5bGzBwaCvVIThv+ohOJg1FOlnCTekgSoG6TOgq5ARMfZARKk7
nxVoLeNlUM32DlH687TwsNDOICFdbZu+hHhpKHPCpF5pdDxvTsrZ4GPfzB/+mPZ7
ijDYpwnOHbun49g8kQzoSTI4bJbMzMz1y47sQFINyOKB6UdA0FmwHS7p++w0oD5+
cCdSEiwn6gtSB3kBH3E6webh9YORa1MLL9Dc6//4Hgqob/tuIZsbOyh21mQIakPg
fw6sB7gxN7Jg/i7eFOa+fNtdx/d3JEeXWLdEZRB/9kI=
`protect END_PROTECTED
