`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x657D3cbpXyQ4N9mC2tip0jugmfrYZL99zLlaZ4viZydLlBYgcSBGhIMD7ACkX7V
qq9bEKrxh6XN8r3hiImvdpvCXAviDoJU2isibQtdTf8FD9q6fgOF5XE2qs4bjuY1
7neTTaS6VmqWdyVDS95CrMlc30YaqxBXTns0M3u7WKhY1cEBFtxS5SbK51IGNE29
5jqehAyCvspIabk4HikA30RytyB0PEL35BaMdrHW1o7N2f47UzwfS5DK2OioDsQz
lMSEB0Dv1YV4/OKuhZgDs80YUezTPlkOgmlDjoJghQ3eZRje8MS4S2MWOfSpPw9R
+KPa0Ghn/yMjNTcWsOZ5DZfT3PNSqVG+cYZjNKOkfLyHwNT9K3Q0u4n4xOmDhSbl
KHWdibCi5gKLPqIlTYLFXVvmxdE258XvaswbuiXgxn9tsAfWFlu7g2Fd4DeIRNwG
R741DOghE63uRML8D50Ps1MElAbvNCaZFtXbVb2TDJtRr5JgnuCW//94WnNZedHi
`protect END_PROTECTED
