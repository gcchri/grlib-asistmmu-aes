`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
POufKtwhs1dCbkPk6zYEXfgQ2r0ou5nH/nQdH04mb++mWzMONNk03/MppFAwHkTb
9V3p3PCRGA1UEBmVxGBJjGdcfdL9ix9e+0pKh0JJ4RkD0yNXOxvIomaxdxgBsWRM
f9u62RmFvpCJDfnKlul4GyvWWCNL3KdipCkEhZp2AQeYNQilSNNQPT9L+JVQGSLU
VNgR1qJ2TTwORYJkPX20WD685xxUm3h/5gVxyPckamjZwfqVwF95pkGeXKWwvBKx
EJkuounvKTFceqcw11uuJf2CrbJcK6jju8KkBnJcQVTPYP/4xyiPFrmg+p/K1XCm
UZEC1AOdGVe/0/NtCB+t5P7yD37HfR8AGn7ENVjB9xQah+XRaCdJjF8Ja3Ssbrel
KYuaxwDemmFw/2Isz4pQLNApl0a5Tvn/D/k93Q27lgumpQUIZhPiVZLmqUl3z2B5
zWS3PHUeEIrRPcMxV/A7eyvzrLFC1KSl9yFgEw6E7+4ZCqdyEwJ3xJ52Oh/yKV96
C4ZnL5WkudmURlPSBcbw52vftLcd4io1PrpdCRsXXf1+haPnv18fN0nMqFDNrGoo
hdmCTLlhLeXR5IfklfmT9Zek/OaaLjckFJ+z9csituHeDlpEPZCcpCeRLa+T4ODt
OvVK4bwN0saD6kXB3poONvEB26TnIOign35WDDi4qyqOS70gOq+E/8pl3WMkbqI2
+9Qe1gjuGQbV9cBQMaAb/nJAmGybhuaIXsRD3fN5d+lkDcSkxgFg2RiyV0Se+Pip
tB0uU3j72EzAuPjLSzeh29uAIT5rFJjd0HpJzaTd2XOSe9KTEdYb6nEoVdk+bSjD
BK9s3/TVDzuae94aKazW2R1Eo+kTu92tT8nqLjeaT2npRqb39gpjzHk0KBIQ9dhY
Fc44fffH5OED0bTJsV5wNFVH4fx+M1YzE0eOYXKYLh45mMhl5Mmn8lh9NfQaSwku
9Jjc8kUupK9h4B1CAMEecAq5EtBAjzMUmYdkQ3W8XvBd3D1DM4fb5h0vJtOUordw
Samv/28AA7REHV9w4+hmD8KfNNEvbYFt+V3XbXoU/6t66210JX0wGVtZocye5h+k
UOqdgU4r0R8fN1qqabtKryoaGpb8DXh5KjNvcAsNt4JqpDAypmWA0O4h/swCp4S9
t56gdMR0BqIiemGOIR8qBnbIUX1Sx/5S7HYyMwESRMmAnkRsM2IaBQAmL+PGmiJs
aXqoXTpwxjCzcGwmCDy6sDNddmSuV+ZizV74JwfDskac41i0Go9MfEMcJXW1J1uW
QYvtlpzlnVnT86zLbCxL1M2OP8VGm+35Uj6GavKHZ0EuCvG/ombq3vd+DcMVkq8E
Zrgnj5eLqlJWjJnDK2b+uGUrnM8yscaD5Kr3bbj/D2yqQECZGg1IglG3iDSBkeFi
qOna59s1zYMcwcTFaoU9U0uljFVYpjA5NybIkvhi2y6vYW4JcPDKZaajjq1aClLU
2wesBRoZ9LHeyMBdZfx9WRdr57x9dntTOnf0lbVJLn2+bAocTWPfLNxRWmmQ1Ysw
ro7I11G0XHCAuLKaU4zjLC8BemTulyddhC5pH2X+mc/iIUhEZsGMOnjUImbAgbAg
wZSLwHz8yKyTJpxuhR+6WgS96vkW0zZn1f+GxQTJdGpIAUmYhS0mjCTBFM+Z5fKP
CUKNBos4EBmTdIGVrNxs0ipiD8QtybvUiGsRNcHvU2CMU674xSfhr2TiHRAnOj/M
yIl2BNMLKLs8M/o3ikZo1Ukh/YGMYhVFj64zJmXopnq5EH6NFuoLF/wiq3agRDLF
K2VjVnNotx62QBlMCIkBwLvjGweEotfKGiAQElkkjt4qWD1AiI3VRduZIyIdHR6a
iQgp5DBRrOXXPxCrFnOnAZqDrE2E5en7Pba46NjbDDkDajzvcB1wizmhoP99I4jU
QhYuuOOOyLP5tGUfeWVMa2pDGUf6/DPGiOuY8i2kVDinWu1gJBGdlqlIkstsM47X
0BbR7GyWKsbdJV/CDxyBWx6Zps9tmvBX1AddoECvo2VgmFhp/yvOU0PFtl/TRKDD
3205J01cD7B14VXU8Nx2bkkGwcSQ9uOL0lIo1Q7/IEkz+zlxiOUvrzwbhaigckfM
byUECGJKS0r6eY6CAhT/tZaGYE2csh9s1klpHqEuPXpnuzVF/ohCUkXuh0ID7HV0
5noucBcjHL3PpZ7KTunjZIUZcqP/b6pBFXQUPfoN3biDBMGMcuH7IVAfmUfb2Olq
KlZ04rWXIlcSfpKcw8eCsNWaomnZR+fTHcIEqUesMVgJJp7hdlrCld5PNZROPfGz
i4f9ikO8lVd3gQanLlCrWy4LZ7HDWCemPMykqeD+AY00VYXKtmN3pvBnDEJq/an7
ygBq9FU+r/re+W4BA7V2A5BaD26F85bubdx13bKtEf930rH6EbiQ+bf7uD8VbEzH
Heb3x3RYtPGIBUyclUz2ykPRZrsNt0Yl0B24o7em1bmUDosXKF6yd4uOIt65Q3u1
G/yLYF7YCJtUVlUBQyeb2BXQa8qWewWqSrLkglyBnBDYRhwnKaSBKiO9CZtIIbbY
uDysYd+u+Pp3hxk0BTO/iVIEav3R275C+P5k1Mkrpj9VZuTTiNUsM5vSc3xra96t
gALX9n+gCaIzgXvP8BS+bVrjVOM+b91oqp/N3XHPxQFMeSXcFSS7o/HVw61i7BLN
wFNppNV3gFuWFiM4wHGYaaEGHnJ26wRKFZDPvumHyF7xapwUfJggSemdS6ssZ8gb
yI/+3iJhMlE+GoI3S6qaBpDDW0VCbDimKzpTKgtIdU4HHqNopjvNjiJWNeQs5DQr
iZBZ0XxZgWRD+73lPe/yO8TfkdCTvZ4EX31uXBKJC0pcdtCp5vEwecb5xnA72vVE
qeHIGPq4Ux9a6u1rRIsIJMLW5JgKDdN2cmo+GW80KpXBwS5/TTX3R2XkF8y8gund
Uh6OdLVAkhuVLFeof8shhCkR20OdU5betsHlQGFUesQF5vPBSG528G0VZM6w8gG/
marmIF6IUehKuzFZjktLe6u5HTm8U/SQtVMBIWyNXkgYmxw/0UUbIgc/OLUsG3Wn
JlXwzYstr7vfUELBODA236qaHaETRbGyRZrzV9VO42Jjug6vCZRvbEiGCu/hGsGb
trhKiil736eCFuxcPkJWKYIo1pzzwMG4pS6IuAQR/jFbUEGRfgcy0Ov2wAmLkqWZ
Cr97eGCwNIlKi2HWCeSqHLyjNk+eJQV5k72ZEMxMcEm6gqClhqKM3aAaoLbmijfW
s7y4NL6ATkanuxkg2zVZ+05jNO0FjgyAaL2EeZHhKkpEyEWKlkZILoCwci8Jn2PL
V/jfgkkJAIV5fyTclYhIsys32Py616rXWMvd4S1wkyGg/WcehztjYuBP+vVJLGkO
7L3STiBmOLVuChjAhkEf96Nd0UujPcvXtmieeXCBeXekpfrndtquoAnrHm7cckL4
BN1rh0yAiRRKZ4MckMGLromwq55+59+9oiOoVrNbyMDtZN+iAgiS0+3g26KoTckr
bpQnWoawH2b74InWA5yIFJdN3p1GHKQQUSjtdGnmtDQQr64xvYZvseqlMeh39Rq2
/HQrj2viWCJmDO0M4i4hwzP0JYxBYLlE+i6W8ZVGvjlvEn7t8gxgduGz6GyBBglO
Gkz14mBthBjpS/e7gFEcnha4IKQpnAoHOtCGsf9PnbqksPZG/rStDU35Bd3VVxJv
iNEtgIGbL43+pDmqt8YlCqqEzK1Wq9mOL0mpjJ+8G95nV5SchiBr45PV137rfMv0
4g6+pHXc9FdyxNLGFD6qOD/g1wkjQ63t4/e6kIJHtnMayFEt84+dyJjcTR2m/3Ok
tiPBBYRczLOFMLj1LW/1dxYLYSsccTJGXXsUwcXhATeTDH5D1zw9swO1ymiIe/pz
jxAO9m5qimFaPy2y8FX3ajgabrDB71kZPqOLRjWEgJXFgu4sW7EtI1Czl53eYl6Q
DukDmozAVnYmWmPT9zTDFkMKLzsKIFqGe7+4X+k9TtaNAr5MG42xKEr+51clFf3l
FDUAy7pYMyoedjpLU8Lc8pl66S7fyV81iHh2QTnAYGxhfB7Np0W/W6loNVN/f9Q7
4k2JbiC+a5wJy3kj3mvGqM1v4M7dZd2iVHLA7yC06wVJ0tWQp5p4YZzKZYmA7Trr
ZAYZ6zKpBzkrs2Mo5IN8IYMdwVuN+L8tH9hBT5eja06mkaYfx7yqlukuCkydEPyL
l6Cd4KqbboZ5ACCl6mf/HmyOEJe1tW6hPqgAsEsHo/Mht1qJVZQbsfo/No9P4AsO
njuzzLCxJLDEDcpFdcCBzRphY7QRlw90n/fj4nb4k3aY1BkkpyqG08nDZ6BGne8R
LJb5pbt4rY/Be/4J+LmMDFL/beR34KVrX99RxD6ZDm37oeSix4+m28pmHpM0Illa
iNcANxFA9fnxMkUlMh0WYFvh6Ei/lg99qzwIDZVWDScbYfKjbEUol/rv5ImjOZ6k
GPyD7uhE26PbAP7pqhJDn5QkBlO12JdZyMCV27+qIWnvvtsJI80xQmil+js60VX/
w2MxFyK1wEP5Uc0svycMXDwwYdrRChdJeiG2cjIdYS85QSxEGJ7646Lei+E9CBZQ
C6kaxfOtsra3jwG1dqQ00dgxxKxOxoIX85T/mhW6R6PYgvGzKJBOPPoBQ2pEkPeL
O5koWf3dx4a40EtXFzvWaKUDeCFFHWFYGxzYYzyYnDc/QMfY+CI5zTmN/ykW2SN2
jiry4KOJ8xNiKkPL4gQdnRRdf25RXbuXANMuucpQcbF2P2rOvknCSqhlC0N2B6rh
Ax1dt8Q+cE9GI10zGTU+b4y2EyqvzcXwq/wEmj2ExCcAFH+nSuut/Rutpz/zi8X1
VbVwah03hycCb6Hqe8heM/7LGQ6nVxZhT3lfFulylBofHA8Jg259Xx4Knpbff1ua
Jm9Cw/gEuNWLcFMMDlEpF34/uZUR5uZN7q9LgQNiMHfxq5sJMI4fFHIGm7rFJk+f
ZGWKmyYSxaiu6/AOaHXTbwOziiggub2XJ1/hv0O3LcE/UBs9btlwzwTf+v9azk+z
W31umFDof3hIdoccijhxVrILDSKT+72R7HJ/tEKK4ckv+vPRlma3+rqm0x0qfhWF
xEKMZ+RE+MrmLJp+As06EmK+4tWyafXL1kw3ID9+scwSfvlTlrC7XsAoEnjHfUrh
X4lQreOdHPT0ZIx0Pjr8nhluPFwAF4gBeOMzbeu+Kx9TFqJNGuLYUFGelKFkD3yQ
mjRmIFY6cZrmNZF78Ljh4uDlyQNxndxhpJMhbhq+vZjnI/MsGTzwSjAU4j3AyCyH
OVOtQ7E70v9lbTwDrEX8ODmOsyG2kvziKMW44IuiGK553aYlMz5J65lb7H3cE42i
NumH4jqljR9fGKeHdDHp+l+QwwlQOdg5YIKVOayxxW1UdlrIisN1OY+4ZakZoIH+
4aGMB8IaaoJMhD+cD2bu9iPG6qUiBqADYS3t4M6Yd5HBtFhbIPuUbp0ZMApg03/u
6IBhnFfqRNu0IJkrv2DAhujyFMHkeiXCmezyrOYMB9YuFtFQYvoTdgKA0PpYvWez
8LfSNQw9zLEJyKgVDOoX68qwJ8qC2Ap2WZwQJmlBuYDuvAscmQAphX2OjprWoYg4
dKHx7cOFatORe2T5CLTf8kffm+MQWkpvqfKyrh0NxkH1wYmKGuy8JmQIsYCBtEuF
zquW749uueB0q9Yg7A9JPAadZbi8/oq6xA1LzOgkOh/1PXaiBl0UpVRsYT/WXedM
BTW0ivWvVzzOSflzkVXZa/jxRV1hPeW3PIkpxOYS8ivBj2+mqdeMTfKmN76eqGCn
gMkrZI9LBk8FVJ21V3NRevakD7AhvShtjNOqQEiZ+bonsZiIO3lIkZMk+FzjdFCp
KOZ9X/9C6VyiTy93JpZAfkuvhawiKKpbCjULNTuB0vjOibxGZ5Eb12FUo0HLgKdP
f3NKva6foL+nW82GjSVe24SNZoFxhW/mj+x7SfBton7VdfSczNF7NN7bBdfb7knY
QUy1x6FaYgeUek2/eN26CGkNMcYPLeIQ1axdemQbQNKIGKV/p+0x2y5yL7In4ZRs
Je6G3aw02DYQWnXPvoIcFE+Ce/0CrVMQ4sK34k8emm6Sr0FF0DtYMkXkFnLQgr/I
rlQXNIH60+VXoD51lT7QjRCwENiy/WlhYy9raJQ57Bc8kvYpAyIvGrkG1fI6IhiE
8B49Tj5g8sH+kh56OW+bZAkTFFrKzM2xBF1BXitVHYYUjuZYgEExZJo2mu3xuUJZ
YhwZaZKswIgu+UtJfQe3XZwgIwVFXLzhDHyZqD+aSdZnU4ciAZK0NX3gMx3ye2Gn
6HuXGWvow2zLdHQ+fbnWxQH3NTK0BehYumwQn/bkb6XZkOlYapcYSUZuiCzxosec
7fPdfwPgvuzh6AfxOmM79I6wMSYsQdVDDpHhXbpFBfhjQQaYEwBz3P8Zed4Ms2/o
RMfkQIPSWBzDSAPdRlcesetKYtvWLZvh/NcM6iIOAO8Lbts3gZ6SvPATXRBGYjQF
3SFailUBUyMs4LdDRUWBn+y7CWEXvzIfozGEnISPN7A7z3IX0oXwM+jCTcW192sH
yTgw4YN4aBo+S4B303IOHs6ams8QZHjNhiPhiso2EjCDwPx8+0lfc62AKHtbVO/A
tI9Kyu8EwBdKfmPsjtmF0sVMcnrvQKxnn7sT4RoxNFvOjl/ZxbYfTxQLMoZXcvjo
Jg86+r0V9DswZ34XRG7BMpdgdqQ/jVU/k7/3/cpwBBM=
`protect END_PROTECTED
