`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g8NrWw+JlCL9bLRNXASiBWfbI8sg1QS0s5e4wT6ovLmtblDC9+7QroA9ooEpU2/N
IYu7GZ8ToWWbWIojiMSqrDLeQWt21Nknv6GIlr52O1BYKGJb1GPBE5sMeMJy71Lw
LkQflWnrmeNieYr9sFWyTLOuVD+sshaH55+10lMqkE2QIGJI++ijSRB6U0raSL3e
KOxQn6DlnnXJUJRd7sjSqaBQ8wSttLtuZskCwOKmyX+GDl2ueBr81Zb+IXWoXRkF
XVcJEDsO8rb2X72TRbVfrwW4+phdcggeS6NmNo2G7/ByGtC0dJOWIKlwWN3vypFV
a3i/I8phQkG7FWppUTXLXT2c3pqvUdSy7Ud3zXUALhRCl6Wmf2N5keKp2hN5GnEW
gKbakTGKyYKM5KKcj14kQRo/4/RXn4cU1SPuycTJEMbylUwU8U6orNraSQLoSMzi
dFWeAlHHgu1H3OCBWnLab47GOsvpZ/j48fDTJbpu+oFkyjV+iTWNjGY9OngAZHHB
f7j2GlHtpKhbgbocCAi0nd3Fr9QbJqTzDQwSub/1u645qjasiZsmk5SNHe0ZPndK
exHX3j6OI1vIJcm1KYriXDgFep1s99gx81AasOp8og0=
`protect END_PROTECTED
