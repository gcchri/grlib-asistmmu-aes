`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R4BOz7Adc+EYySCwAZRH1O+M4SwtuXONPJjMRb2s4HGRXOhAx6qhQyJ/qRoF2fMQ
JxOvCd99KDhirvBEI2H5y+XnlUMqOIhb9J2hbSfrA0ZOT6HTMfWts4doq+kl2v0O
SNmucAvl4r9dAMisDHEjXP7jXxCHk7tlrsOUM9zMFP8/8CkRsUDAocB8FxN1OfEG
SV6V+iTZQy9x9OFHlk/JSZ//9h5FN95+j+k94N7EOPWhyzWOmMNYusgI3tMkakNn
5+RhMhPNFYbSiRKvIrniHA==
`protect END_PROTECTED
