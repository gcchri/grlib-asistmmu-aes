`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rCFNQFMhw8lirR2R/1OUK84GNbUvfRrjevhH3yDOGdF/k5kNi/wghcvHIqlcvlih
MsudH+OCeuGZGcGHrAHVAHVARtspcmqM40lqlEJ+PSs0KwmK8HBjQB55ED305r7x
eOkbLWmdZ2q/Sq+rF9ac6au2QKRWzTxav9MF6BxpGWzC+6RAE8HDYdVl1/GeBg8D
MW10M4VStKDmfnlf5r3QIa6Y6YbsDdHgTaLFerhXi1Nh93hYxyp77q2UzZbtzf5r
keYnaI2Qq8jyWJzbQVKidceXXmMcUHUL00n+NILNVK5PAkpZemClfQiQGd1YUb95
1AsFb+XqoooEdMymU7V9Drk3CKjThXid+6sZd07+Qi5LhrKKnw3RP+H7vYRagXPO
Jd3nNtC4Wab0KrMe66Dd7Q==
`protect END_PROTECTED
