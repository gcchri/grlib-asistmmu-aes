`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E+ElzD4Iw2f493IyFkTeX7oqEpbKG0kUh6uGRacY6DN6faV3qGZtnOEXzYc5A1Oo
cig8qVReNFTzjha29B5dA/m+X5yy8GcbvbWLmEPJvjW8QwHdTOkhsG6YFBufEwwt
N2C/IyTnX2kOAFJX5heC5DlUumgl956sVQjZz9YVDuKtKDvTFolMBCJ9j43ZQ3sc
++7IdNj8WK9i01z8Dmi0IumTnvCw7kgwpjv17vHcJQVriWmmHWp0UbHg+Wdgx6iE
JpCFLR/BfJuhkvIBfjdkUUGxL4inTPY2eGTDePQn+g4pPMyQdyIfSQmamsKjr791
AVM7Tp38Wmk8v9T9Nivuz/kBKKm5mY8qGAwtjklY/N7ZYkkk5cPk0U2s3DxdeC9t
wXW77EpFk5LnWFDnkq8/uGUm6lodn0yy0SymB8S2jkM9isfkwtg25Le6DWIXJYuL
51IUa7e7BqioPmg1ziZ07I2qHKQJy2d+pFr+I7rmx70=
`protect END_PROTECTED
