`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X2J7M6VtjEuMM8xq4PQdHnPgrLhGPrEPr0L5W4lXHhM8DZZZwzYWnFdlPiuPBhN7
I1EIXoY474DVcVr+0//QjHnU64a3Jb0X6mNDN4UKRen2RnBmddtqqyEs+WxQaPJ7
HlovM4XuLegSv9MZVMXidfRuo3611rXNB58xHsrLmqeiaVfOrDvplKBnLc6CXzKM
FkrvrIkrrmZVVdhbDUbyz2UvabV7S95V7VorTATPBQOfKmO0E/pbUem2MlPuPMt/
MAFmKkcwLPQuf9uod6A4469JBaYFUca0pmVXvrynHtVEsgyt/3IAFDs7tLirDpvd
+MSJK5bgdERlxIdu8GYf2q5nwgDl3JKxJl7+8oLBwMftO5e+iJbwtbyIXnRl3qfl
TSl41GigJcRRAvI79FUWOf0szRfZbhs9VPumTBMwIDjl7LSYHrxf7PUIoDkcbSDU
JniB20mpWlJmeIxi+iUXDioOiiZt2Co2e1ujKHq5wcsAMivMCBMt0+2tQLPPuSP4
fadOJAS7GhLRLrBfpWigojojrhconlr1UDJPC5kUOCuVgID1VYB6mqEarHKC6vP8
GztAQKhro+PwyYpogq7mHcp9Nogm3RV7AMMuferIg4OTjUMgAKBRh8sC7ODKRl9W
QxgiGl56wjINoaIjRBhwwXE7CjTFujUp9ki1zeU3J4M=
`protect END_PROTECTED
