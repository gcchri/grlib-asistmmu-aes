`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s1GkoVXnEs1otjcS4rvYVBcm8DKGwajcVwqWIsP2HXWdX8t+c9kCzDcCXa/6fcNy
wJQpQ1JeY4J8NYCjqxJrd8uX3jAc4m9qZYsX0oIHTCYQs6/2jeVVRAe/Fl51jJV8
hh441oBe1X0/IBJGGfKiYxy9JQCrVCYwAY9I4VdEFKMq0vF08ial4z2/DgoRGLHO
fDJpt1A5lgHzpC9CmbXbJl0g8IYWTkhmVEKItf6rX3hXBnxV1oCGn0RD6k3aWKUf
B1yzjv4LE7akv5I1VyAju5gu5UaEi7PnR2ppOPTlhMJ8nvokpW3AnGJwbd8oJ1aB
2rQarREM/aV1nEeDjoNWUvGswaxXQQnppWmZdYlC1p5DbgdlbA8Dv5aSSjIYmkXD
4HBuh2lGL6fVzlWffH6kNhOtDS5uHOh1QQp3e9fdzTutpvnZig2oMfM1jkfLotlj
7Y1JlO0DgwmQDr9QA9ik/CV3ciNpcF11D7Turb0JfLc=
`protect END_PROTECTED
