`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iyhMKLQSzumEhuey3+/FbQ8LSmHHHFuiR4X4noLt3+ggK5KqZ+OkpuDaIsy8lPBP
MlxhWTpcE5NRwiqfG7SRKIWg2iKetCmnx29+z6VbtQESYnMR6nd1GI7Iu/edkk4i
PWPG1cZLPuNIqCMDkvaQ5G1J8KtZejqOihepzZQF3d0HtH4jsUaNpTkVmrM+P3ye
nJOPvQZ5CuNOR2nbLcrfb2rjEH4+nRRAm9VWXTEMKCukMInan26C3/7NQ/D+RyXU
7JG6m7te23rfZHhaP4VShGAsNCivvx/NnVRU7p5vR1QYYEGUjo2ukTc2v3Xgqo9Y
XV4pdV4L98rCo7YF+1JTQxEi0WjdbBTBcBE7JQ3Sq+G2eGVH9surNks2/aB6fz8+
6B+7DTjJEzEyAmjBSsZkR1B6+rS3y4WQyx2QRxNx0QsGE9gP7biT/OyywwXWoiTp
DwIzeLXyvWFENFvOsViuaRYlG+A1pu2Qk+PG/51fW1I=
`protect END_PROTECTED
