`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5biDjzal6iJ3svh1le1kTxGSVBH5EtEGXGIhLMa8x3zT9dUZQcw4xoYv+hWhtrnt
WqbNdIPGWbwVQ9U7DozFWnwC/vJhIwDlGfQofQYB9FdJ25A9kgFB3iLiSe5FNdB7
RzTLhsq2uEEtKER1kNBRk4Z6BmqWO4S/n1kQ6/QH578BFZjS5xQ+4U3cER825IGO
mFrV3T1RRqRTLmGf+YGd7U7kBxNNx+PKDRaxJ34yLE6oDnyD/F3CpmWm2LoTE7ku
pSyLXIlpJzJX5cOO6Ds/Ee3+S67EA2/AI0KH2/A0mGT/jJsn0++D1Cr3IoqMt7GZ
W9BrWz+h9m4jIEmxpD2n59OZL9kZbQHDwYAvFNYmwtv42xbAPHsWg0jQLuRHtX4I
PU3B723u20SqHHdKrAjLoxqS1vRaIQRV0WOaiYTiKPpcHLPVEa1+q0IKhmwahiDN
HcCZxssEsZ1xSt4muUATP11DdfKaH4ucezMyXJdA8UwEqsUqJ9ieHFjroeLn5M2e
4BfQIRJdzqDD9dIX7VuH3AQOlRULWgiH/jiaH4WbARSXjM8+LIq24rddflpMP0Oj
yEWn8mVq16R4c3AWixqi2+pCWj/XJHBD6g41G4WYe4bNRAEft5k+la+tONtTMtG6
NKqcc5InR5QgV3YgFCT3/tkZtWV8ZWuN+PFbuKTzulvNHm50C8iDs74wQWRcHdiH
wNlCaeCPWtwzfeqa5R1g6s8akngXPKNzqaFUmeHwmRf7dSmlw/BC9EkIAn6nADl/
LfbVSjEsEClsvgwE55toAw+ykQuUuWOcUAZ2k2nVuQMp2vfZCre5PnEPfesS8Qs1
4R/1+VF8q/V3GVAInFOUhIOwAsnbU0PXRTq3UnFaP2DevMDGH4kSqbS1OC3EfICN
ku+X9bxc1tJkpFggflS/cQU6et/dGN/16FOYNh+qwtPLQaqwFGuCXaaVgNJ7Yz5J
DmhiGSl89WSpZIvwKR66+GItzJG/R6EVarppzpnIphNgZeKCDKXwwF5vn1g4Z5vB
qee1KH8WhMoePtV/a8c5M4gd3B6hiWV4lRdoeRar/y+3MZ/cPkjDueO3UCj/j31U
O4vYtPIV+mJP3Rzbv/QzybHgqEM/wmVUHdTuKrUK4cYuJzphVVlh+mQgU9YDkPZa
gaJA5a8q1VBoj1SwybLK+M9jZWMkBWyV5TOIzfZ1OE4L8Dzy8GZXd1igLy5vkdP3
ENWVGBiWaDJ+bkyBZsnS/YbHa1gdZautEHog4wYppzgiy/xK5GD/RsrqWlOULXID
MyRegsPNLsQhU7Jd6PewXUWtw/s7zx7T5RViNzaa2AprbFCbnSBnla81gQCAjvrb
J/zrKhB5VCVujzH9mzWsSaSBWGHtmIhMjtReC2S57LmolvehX6vSroBMIkLrapMb
QCr4CBUB0KonQgmVTtekt5tCKb9zU4SA7P0UexBAWh8O7g3KYu3qgeCHfusOFRfB
qNB4BtiaKc3tflJQwZXkby8lp2z9Lvlw0Q2Lr9PdpspZyZ7KjcpCVQrm4KzQvg1t
IGwm7Q3Neqe4CJV4E9f8tYzI9x2I9nDnnOQmKgpHL5ZZVceYErU7n2GfewZCFzfP
lQBODFuPbdG0H2g7+brncvKbucWttL+rZnFMVIaMHlER+xtU1BoQ/moK2dPtnCZ/
yz1Fj6qS/HbZxjJ0kcZAokmE3wDMcvKNUQcpCAfvEoITQPEBOHCG95mCed23JPLL
YspqH4xCc3G3l+M7pMppuxAkKz6GrNb6AZU54UilR8ynX+ssqxlKqTLWunQaPay3
xqHskh4kYaC7FeNxu4T/TWESijlUOyLAq0u0tH3EE+lcf8tGi4ii8C7VYQGm9FAs
HyY2qiYli6uYg2nZbwLt9UGe6s4xT884xK/gqt2ilqJyIbh2ygVJZR44m2N/+JC3
R+y7NKwKGXnFECe1/HYvpbsgVS1O3esNtVMJLpK7wTpFmfQ4rv9IlPchs2wSz+iF
Xnty7hD4NsVCQARl3sAaQA==
`protect END_PROTECTED
