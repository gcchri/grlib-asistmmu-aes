`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GWqu9oXNG8Sx8SsO4DSSovFYl5buMd4YdzTjsM06u8Y/ExxJ9z2KKHd7NsR2ljwr
SZpNMCeWHobCmIggGXvqD6sRA0Xb4YlMeHpn01W2SJlMgZU/rjQAjE5fNkWFo8rD
tw+/bbTA6+gm9wKccy/8jJ0RAGrjp/3COk4YrQsmJAcc5MHYLMFAm3ae9bLWLHDC
CvqMrxvmQNaCJ9zSOhf6F+3Fa8SAjDxgCVcg0ideStv2PdJWxBydnYXUxgvsp48n
eq7uOQPMvEuJRm4CAL9v/J7FTREjJSnINu+bhgggX3wUiWWqzVAqjESysqaMlMde
6FRBSoWC7XzqWB/80tgoZRV/ucpEz9wEc00NO9/Pbz8hP7g3vovl5TgKG9a1Tplj
l2f7NqoTgvuQwkhgXvs5Tit8h0VFVynUYC0wPRMSGGlUOrDXDGzaQ5sBLDx5UWva
LV/gOqgFY/2ZSl0PlrAZoV+AKX79/Lw8GeGfHcxfInDB/y7FTzqRx5QgM74xrrdg
DEMJlExvIwKNYizhKYA4zqwwRjaVpy26lzJ6y84OqsnOGNFnPGFCM1QBTP3bsu/w
/Stx3V2TFay58PAaRS6aIy+aWPpCBbUZ5UIeci4p97vUZu4fKZ5oEwEW70aR7VU+
r2nekQaxZ1dBazNaRTTme6jzJQCNkwVxfBDSl2yodtmKfGKIcmDF+SimhW9gDEFO
QRndjUAeEjyPEsBQ1fIke1OoxGD4huIIgOlE3PkevK1I1NiHLM5woJsvt5GWSInx
BrZrPW/T7Ry0QYgvgJI5kf3Nvv5ZxlssWuDs0oyUCVSfTvV7nW2+QAeeXi067b3F
i2XXc3vugK6yAVZiHKGSBxEe309B1GkydV8ppZtH24nz/jVzyEj+/A9sN6Uesyyp
JCP2IHWx/JGKYHV17TsuDpn65gTTlH8BOWsjpEujszxhmPGUNM7H8OpSKXKYJlvM
gjDb3SfpONtxyjgyBrgOxpSfioUE9tgLy9ZFxFM8xLX8N1U2yzgsSTJrFimLixnO
QUBlxQ1vLQmLQrsVmzI2niP2FosD96Kl9CMFpGsNkyJhuKnSsatKV0Dhn+4rwuLK
SZHAEzl+EOmXeq/9zgCb81qwGIaUI95J3zEW/peg9QqoBWZAxGG6hQvIrhngbBRT
7wfZqGZk45/G+qQXcvgtqjJZ8oUfDIvFeciYLdS+xHakRobMVJ2twA7Nf3M+IHPf
/nlxXflfJthVGZs+fp27WkQBjh0TT1MekSKsKi3RLs5AfTyt6u1mCM6xqikhFpT4
403QIZqrUyGru5lg2qUBfA3LhylGHGd7Pw/JFvcOn4hmPnmv78/D8GO8jixWBOK2
5U3lSUldfqWzGOeSXKnGi7oztEk1vNHi/ly9lb129LKPf7r3gQUON8Ww4XZyCxWX
cMkAAkkzV1iCR326mJ0aLh2OIJvpGgCv9irkeoY96ZraqEYcaabQwMKMQYRrRov9
JHoyl9G2akF7lOsHbFDZnmUppbzUe8OOqyRphxBscIRLdwYf+YSIp+3cceaBeuQr
mKwfrbAegyTNS6/6lNt9xHJM+qLR88Gx+ic9vfbgXsaEXdbUfqw12yqgT3ls+LJ0
Y6cP0z4YBepsA0U3HeUjuQ+6giXtTHusiPIll/IfNhUF/CUQ+benT7bG47Gbe0X7
SRQDiuOno+zKxFzpRxCS8ZGBPThr1sRc5wx6W/GNGeQtw9iNswPFLGnLW3yMnSTs
BBFo/Nhhj4QUEJ8fGQHL4vBwlfshM59XayIeT6oLykzGlNfCRC6IzDWiVPHfKgFo
DW2R5oD225OA8RerVT8EUIU4BkeAjpMEtt1nYVg97X2j/H/Qc5C6oHjOxHshu5ne
5iLMqmbdd3F7gw1Xq3aROyoJVU2ff0b7bXgyqLO5SvHT0MLvOKaRLwFmlARggw78
inzW7guRfao8z0UxIB1qBegHIAhBt7VOj4P3J/szFWyh4uQxe2y2TcDKRA6u6aNf
ki/nhKaZ+jYot6LPq4K9UO6VYHDWRMGdQ8cNQoRRwqhFAsAjDs3wpdGJIDjy/lX9
4HARIuBttCtoOgqwZcsByq/GPy2gmSwLfxuO75vZ5OkYH95cO8QY9q8gd7FbfhIg
ALIa9TWR9pBwqswkjmbkxr84OcLUElLCiU7Ih/15hoJGTfU4yQ9VgOfRnsv5DybY
8lBS/WtjgwyQ13SE6q083uBYj8iaAtXilUHRSk+PIk7q8w4TZjMzm+5RousQG2NV
XNPq+sZwSFTysZw9xGgjJ3OFse8Z8ZqYa+KCVpDjrJnzdxzYuJcIsm1pZjRYfLd5
KAekvHWc9lu8nlfkAu97G+OCY1fV6KAzijHy1z47E8y2Rx40XHIVWWYBybC2co47
yRCbVaLutwto5iYf1INL5PaPNFmuH9BjKMnv31bQBzjIsRUSs6ihS9r15ojhANX7
3Kd5f906/OVYeshjEOHzvEfVMh/CnzrDDaAESh0xm7EweBWVzMt9IDr7NzcnX15m
LSukHRHfV9E2414tpITL09SA2lbLGZGDCBwgZ1WUoRYvQKLjwS/LITsFKOJPYH+T
fr4MNslptZRnbG22QgTsal7Ihx7Dy+FoWLWKJ92Eo5p1y5Vy5p3ADljqf4phC0s1
Bxh7kCQ9QLUnO7LljXeh3Qm2nD+Y537KElxq7SH70r2J/EoAuRWB4NNbAUP+h738
eb2h4eQcldpC51fYzoa0lxpwE6jHyiN21DqmHO8H/uwx4qeV7cT7VBg16r0F/fSY
`protect END_PROTECTED
