`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QE38eDCfPifSEPsHuUOQs92BxNdfa+KceKAfDpH+yZXnI50HhXs+ug73Is0lhmcC
BktkV+vR01wUJzbS0fYjx9OY6jB+2Qfpzl+Y5sC0diRmRaRuhJBnQa0cW/k+nt3O
Aki25Dns7SfpP80qyl12lqjB5yqWx22SI9M2mm9KvFmlOclUP4rWT/NqLaVoSo2n
rPo+uyFeIwHqwensyAuqiYNrJJrNYKvIRgTVDcdVNq2OEXFxL07u5OgzDqpd+6PY
WQFLB3LUTcfxtZqo58BORQ==
`protect END_PROTECTED
