`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TAoK+bEdejJ6ijfJmZZfjzKtQlGoYg9v7GTQg2kT+lg4tttbV+sGbBw1ZJvjqbEH
bSvSxq1bJ07LDNKkssEhaDDtO1GSBFMnvyLAa95DIzXysOwDZVqoIzLYAykkwwFs
JHZAvhd4YTKxQkTP32EWuIM6ULqRL1yAolcZjxw5FXdwoZwPXmVPKx9oG5PCEohe
Cjhx8iGm55bGzqYmlT9eoTcSe+/kYshg6SLmHlcxjuob/9jy643eDTaV7dz6j9LL
7/Ufz6DM20sNBrbmkFN2m/5dnvvsGskZMlhm0gnFFlmKvc88L706SWUbMjylNhmI
5d/rLuhZG7jXVCv1g5hbiXT15mMzHZ6VjrWjS1odk8wpQPMePq0BRctYJClEHHCV
jjwIJqzLiMSIL7D11hrE6Udx+XgjucbELn+rt8/TM4PRYQdffMnIpuCyVsRdp4Gf
WAtXU9lw6Y6kzD4PaT+G3KyciBTOxKz9aHq1C1N24AOnaYLis6jQRmCXcdtWiRJm
F0Qo1j5dJb745DTYVDgDXl+vq7YS6eo/DaaUqDPxqzzxjPdlMzDmmtXzzE0iOYDE
GiFGpWKWmcKJPNHgE5vlnWF/ksCR0rgBIqC9b9QK8Bnqm5bIIAR+iyiMdkE82bzA
Yhd1XrY6KW7rM490nj0LXA==
`protect END_PROTECTED
