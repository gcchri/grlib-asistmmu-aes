`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HlpRbAfkMCwl3PhH1pioNg4mdUCBiI+6Bu+X+NZixsekZRyBY/xZOgsT7nf94aPp
Y+iYAwoBgUzp/SVI3bIUsxPnCR0mXOIQQshexvTEI0AelkZlTeIJmNI/XofpiFTH
ZCk4g/XuT8Q84WU1gM6xifiRDdtjTuUxwxkG43aY2ldC4c4mpg5fLmzpz0dRcKrq
wBPUytWcYIXntzmwOSj88STxEt1Erl6Dbz59G1gfTHE4Q3DqiGxOuH8voDsYQGEu
j1w7lHBa8HXc8rmZG/OzraEmyNnz/TzkHX3bVXYV7Dj1gbnXrdpG3TD+d1F7743w
43Ezhatvo3pXic8oqbx+PvFeEx/0/MdKoKWs6dA4W0pASM8P7M/9hDUaKZbbPPtK
W9CF1D5tonK8578m1ZhGZrXnMJMssi+re1JEiaIHtp5jKKTtKzCKXXJtItoI6JqQ
7+mHvaU280sbKsm0GbZdvQHv7KojpHLI59bxd4d1NzQWyLuIaYAmKRLJjRurO8oh
Ge8GmUU1i5sFr1TnQeAC5K1PRLpxCyTxpyxThjt/ZRPdeGHmwiXEyLhJdmjXWd5w
lV+24XuduI7tKGygj9OIaKGGjy0k35bjtFo4BWD0UQ3DkjYgWWe3wCVLHRPxuOfd
5pN24NFT+QhXT7xSpHFyw4ee4HakMSxawcW76K31q42h5cSi4l6+aE0NXfgka/gb
hs5c00Z9JOZpSikEQUouk3gXnS67z1V9qgcqQfrnJ0WLowTW0Gn6bGulorAWsgs/
FMqzfNpp/EI3fSCgLseMyo7b41VSYeqjzGXjO8PLEdtxJDSMygkziBMfNiSr6CS7
cB5Xfx7pjzpE/s4R0H29nPiZA+Buin3PY3hdKCDQ229IBlV7pxaxsfJ27cJOcwMD
jbTQf4ZvDo/9mnVA8zDp7RLJm3A46M2SynRt9xkjvAEE0J2wTGr0ndN/Wgf4kd7x
kt2JTtfFNhxAALxO8BnYiA==
`protect END_PROTECTED
