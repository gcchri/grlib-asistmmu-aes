`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XyJPrqScu88ddDgVfIsP1QepE74CuPUIoMriOPt/fhqu0oNQQGQZL4lsmXoEBrWn
/HI9HiNBqWAV7eR1HjbF/J5ugiZx5its+UzTTPmGPEWEBtErx9tzyMWtssxf/RtJ
MFp4vgqf4PWLSGs9QLSJOITeX50tGYyLOaqsi28AJMfqeA91olqSB9GmUXaUs6Ka
uPO/nhAoQRn+rxCfTTDnQymoQXLx8UrI5jWYTM1zDp/Jzf17hCrV7QCJ9SiDo5A6
fzsllWC85arIYuv2Z6XdjfCRj9H97Gpkif3h7miwljPyzkHxaLDex1dNN5FPCwZk
`protect END_PROTECTED
