`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lsr8wfqxc7x4yjSUQ8p8+svGOon7nzSPV+pN10rbKumJyeLwo2+JJ1I4H5jrjRhC
eRaNSMXmMKPhj6a04gVTcFBwd+dFXH+XUnt1JCDlDO6xsVMC654E32mJn+xfgpW2
uktGh/+kAJWkduc9lxh/YBVSyQ58FdtQqFmwiquGeNiFsn1Mo6rwAAKDQINZV+3i
hQBcLwNHBxKizcf6CK1tS6ucvyzkDKrBEo8HJk56s6dM/BmWhGAQrmqhW1damyLP
hi6a6L5JOJKlO95EQPg+H2Pc/1u85KQaLWH9zmkaK1GqGKAzFWC5U6TJVL/fevsW
HpUPgGRIddfed+BAekJI4g==
`protect END_PROTECTED
