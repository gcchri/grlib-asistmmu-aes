`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fcjUULwjzBEuugwqTL5G2kgC336X4Ve3JxrL/YuCP5HZ5WTx5HKKDLWt4ULoXobJ
urpOvz0iFlr3b8WOUc0ukCzad85bHss+UHLypfy+iePvDVkQg7b/ukaxNti8cZAX
s1hTG4Gsek3a6muAoxL5jtFRZ1GthWEoh6osVCaLntxlgy1KxYPIT81gy0TQOptw
BDZNw09irkMTHxNSgWJLaS0F3nEHkoUixJwXvmUKnH+hKrT9fIYKs78/dl1CMhp7
/laA2atNVfxKqNDRhYYNpY8xKA456GymalHT4SQk+c99CQti8WSWotQVhCrOQp/f
TNSHQXryw2zsNZmw/n5ia97HW7VxdwosN8DREoRwa8rBOMsjPKzac64OgDPT3Yc4
w5G9HsiWo6Um2UOWd2x7cT4gGF2Zm7Tju91Dx5ctkxyU0VUAj90UfnKLaCeA8D7t
ANV46FX7BegicsJP/eplWxBs7ZzxAandpuLR5r1PzeZYZ0KlYO7e//b3gg1xs57X
QIzNKGJD1NJ0EdKUKLE1MerAXgIjG0tKcP4STF59pG6GRM6pvlixtAV7Wc69EXX9
mNcZe1yH3p2rD89jfIO80p0F90hnhhP/v9WlYbz/SQZAtD6J/AROA+/ZAjdn4XrB
X0ZpTkDoVJjMqnKH27frd/kLyjvfIVRPFC7+Ow940bIW9AACsoFwXvZ1PNSiGbxS
yzVRF3JdVrDpahWQL2lUhac5Vwj/Nu/MUexOUDAwxYjigIt5iG4QX+VFD/NqWdCb
6JntWXRNjTcXDExDX1kJAGiLNpNfH+GyUdI/iHR9v8WFyS8pdKalgjlPw3yz3D1+
KmiNzO5TJ/L1RZpYCjY7oj+yUi6fyWfkU3e804QpQDFPKLJdAJC1eKFX6vGIsy4K
xfp1CaSvLG+nLaRqOgfDXhWoWUMnjO7xJsApNDqoEckl20XrGH/rMsRii1ay2I9u
Wmzz+61ijH6rKHYIcdIByOPRmrreGNey1w97gVizAqB/I7KAQeC+MKBAVGT77Eu4
By2TCLsTKmEpzfkBAXVYNRLgqSIhjoYVcXNK7Vqh1oS+xCZ0EhGJDlS0fFkClk3j
jF/fwromqVS1h4ttVAe4TRsrsfvKsmiBrpQq3vvlXyUPKOGsz4AXJdjustNolDUS
8aeXKseY63xd6iloZZ0PDug5hHTb1Ie4YQdjs6/wReeOhG0AONvY3KAI0XaUlZgz
usJDzOUlcuE1tP1pFLke01XirAKFyyMbztw3TDHGnkuvUC0UCjOI8mJE5okGdDfY
HgMqgVuO232xrm2b+XC47lTpZlu82Vtp3XknRPP4a6LvSPyCFekBlOjh7OglcGsa
mL0IFemtkTWjL4kyV6UsKp2n5VIDaKaZJRWGWF4wjm049sGXNkZT8WZny0++APzB
qHlYTGWJhz65a216d9Q2TDbPdeEGOLe+MXrCiOlxqCxlewiIZqA/KJWulEZ8IsXg
uY9fNaW0N5you70XGx0w1ieaPHxFbThovJUvdEntyeA3YHiZZufPod0WurvavUiF
Zs6H/bMgc0kt+H0CnkT0FCspOfV/8fw5ZX+K+WYeAUOYSdkx7wTGlBZnNnM5usMb
smYbM/Vut+he/TevhW55gFhaeMQcmTzBNcvvMpFYvFtQY8KdJ/J161UAUhm76YbT
bgWrIuBwIexZEk8qtdbiiBg0B0xknNW/116T9wwGO3NHXEXLZEjQ4wEAIETOcUdq
VcwvAy4st7TxK5y9wpmW51XPIMecS7SyqHjoRaDTAjST89YALEDHG0N8cuqExDUa
Tk848096yHnMZy/0YvCuxhR8cU+iE+z4c83ZuJRKH0XHQCBhtC6oECG5onGDP1NJ
mbs0VYVJ1Db/zO5ft/HL7//ZR8nlpG/mlqU15JTK42r88x74xl3SaTla75pn2UTm
GJIg3UfBUIMFZrC+3HMxBkVKTzy8bV+SAqAMeuaM3Hnd1AClN7tjOZi9joD11L0J
vSm+70lTdWlGgoJpZK5MztBcDuu1NfKHc7Kf9oyoMMUYI+lvJYGePcAMklykuuhN
sYdqdI4sbQcPo/cPH4z4dIlS8cKMNkI1lg4igyOitHOHxJRlx6Lz5POBPgGEyySP
v9C/YlFq1KpKPn2/IXbsoCmT2yLQUacJHbPrRQG7/giTn1opHXlEMMAoOvMx8wio
UqoN9O/I0cJ+7zkUrEBty16FAk9fikpQBPpHDxGY7cvr/nV/yM0nSnukSEfuKdTf
5lG/CNVfxhR0U9To1owbdh50XFoFExpL72WC1QzaKFyY2lW2xMjUCBsvEVS6WSjB
EY8qn5zRTkHWzOw+QL69yih6VguyPg/rQ2hyIVHTz+0PU/1K8X3V0ICrUJbd7WOt
pHyjtSSy/leS1b8VIS+qCDn2akE99zBgcNdv2MtB6GKwvyUpcjdTS9aOS7+r2nta
f0+IFSBzYjs/xENpnxGOWh2uRChoWfpwl0Nx/w//YZOM6VCzjRXg6JIeV2fM7HL3
4jloPHwDbvl2aP6KdfsJsLsHlzNuvxB7zKWhe1G+rugd3fusYHiOGktz4E2b3HgZ
CbJwoSjrnRXMtrVXWeyqKf4nGw6fBsBKdoGapcQE6cRoeXs2wJ10S4QQWiTI0u9J
eEjYtlDe+QzyzJt2NsYE5xQF3dW1/uoemawtDW+OII2bTjlXZjOooG2eTG+HaqQw
tuCUZa0yBh4paiWNkjI6T9kceP+WPRBhUdi0StlrrLpja/10hoxXR8IIckNUEXfk
71E9OgZSYlp0wW6UA26o2SmEVE614CwOdBIE9EMi6EdhttMSda3/NcCju7N2OYne
hkGRJU8eGULI5azIuqeh8iczRwmLRPyksOCBrUUgqlOorzS/Uw5zcH/SU719e8BI
52Xs1rl8LJnSCOOlJzEnfXIvra9mW9oS7iiFMZwH4za0U0H+nhaB1fnXpEztXQH5
ZI/Z1tnw+IvPDhiePvegtEE602P9WbGjDsN+W5GOQL4pO3zgS+cQB9/wsFdJLTRx
azQ2xVeln1/wQyQKEB7ExLW/wPJ5jSum3jJpX438LKu+0gEsOTIQ7Ut4ZLkZ6Db8
adn19b1GRIchST4xxCdcUEHl0fUDJjnYRCMszyxZRkQZOT45YUPQYYnCqk3Dx93a
yFvhoEI1G4P0syLAiGqLGGOmqGq6PZ9oaPP71zK8TX14b5VPiI3DfmFcK05S94Ki
mwznbXDNEHee1+O/1zcl5rS0ev59U6Pv8jSdERJ67R3dy+nJQ8i5CYHqc9kBozB8
TDDcjA/EE0wHEHXOkikoyGeBQjI1QaO2viOG1Ind6FltSTWxa2B4//U5bpTUyj7w
7a/mBD2g0xeDvsHOVwxubixDzU39XnYhgFUxuodLjmERZI5nJ9Hdp3Nr6Sh6XA+m
we+QT5n0IwT/NurGoBbInTaxtDMCqLZCPKi+bd2V7i3FebFxln7oqkGUVugrwwl2
ILE3b967Bno1b+57xAdXQCXB//KXiOdb3cR8PXu/VcBSaVATF0BHS61QBJ5BC+Zp
5EcLB64sqSFSobSAhWJEmaVfZSPNYGPKKoGLckF8ol/UWk001ze1bvQ1qGQYs1Vg
CfHWfB0pCaEPlbRByYIZFflB602uNPkbgfHzM690tvEWAxSlxTLBrvHzgwd9xiP5
j8LGUR/Zic+8ggGhwkwof32TUDU/v5g/ST/Zo9tqhvbJammyUFo+K/eQBYHDEdWK
4r+wxN/ImQ1nymMVCVkfGv+RgadF86HEZyKC2d2oZGdS44h13up9/bc91Dnjd/0x
CGGEuB4AWAR0HoG2fxmclF6nmfxVizhrgya3qjj8iYxhiKRYMYqDeTcUWKnIUvgv
CcRmuxsejB6l+U9aZZPHNN+tzXgINmwWEwIXsmf2d1gcSJkL8GvpYSZsPrb/hIZ1
VcayvT4CKI6bcxln/Lz7YaSmDAwl9nObi0LFUJ4dWIYJ2B8OOCCRZaw/HExYZmCX
DM8NVkG3/rm5VWDnbigmUuNF2njUdJzjVhWDJRwrixZaV/Ty1btIl531t0OCi6y+
D0iYKdkGQEJwxlsx+dXCMQx95M7pN64m3ZBEUrYeZxM84/8xsd3J/n87i/aa8B1m
iyNERMnsmjKKj2tDZ/CW6tV6hNmacGa5D8qQR+MmiMQS20pFtEnd5pYlOUpwRb60
OfXTAV2P9Pgds7fvuv8AvLEDUC2iLlM2Hi5j4Z7ff0kNWzaT5yEK5edfCwXYuKPN
yw+xSzNMWj9LCgsCatJP2B5j0te55S1YApinQ+qQnR9JJBFzjxYuqaU6UZqlPdIB
BuaG2jlqjjW25MO4VsO23ng2d7RpAn3QOhNX8QLNCTEnhe5lzofHWhH2a+V7STy+
i6VpgJKT5ykeSH57TxCDOMQc0u9+sdH6DET/DIkq/gFH0T2u30U1ucpu7mDX/Vdg
ryE48cHlxctdNvmHzRuKFcCpcKR0/Xq8kl54KJeeNE4IRluDbUTZiMpBlJNaM+db
WH6qF3GY14Ne5RbRDeuHF/IFxeziACmwVyWnNLsqbCQ3TzMIxx2ytdAzRYaBD7a9
9+qSw8iIsWwoQ6z4cbREM4WJqs+/xoR990MaiAPMYXNsH995uEeRtbmSJQVTbBfc
nkx8FDI082A6POQjdpSa7CeCqQQWmCdWkMYAOGtIBvEazKawCcP3y2MCyKwZxmN0
F1VacsRpmi/WG7AOeqNHN1d7LfajfbAB9ODaH5ugjKqA1ULDdl5dJSChI5yv1Ss0
KE0AUDMl/wAwCD4dsnw9LqTZtYKy05juO2AFpAxYY9XUO2AvVYHGwHyabbbaV+Bj
gwFwH79VRtEzcYsPgdpZBkpzMiTWl30rbksCBH/TFfDVJQ5APhUq/7zHtZS9tfPW
zqVY6U+LjfTIEZRP9QEkEUDS8OeqAOLvDx8DS9Jfa7/kGEVIqBqb5TmyLCJqa7Op
qVdrsICBz4AxgqV5PP/7jvivBFupEAbwMm70bMnOl3CUWznqTSnzt27G6WVEjsW5
xs/4QLplo5CeSHfQjnZidMBgmPb9eb+7CAw7ESne2Vk5GZ14/mHLzmzjhuPoUjp0
Iv375u8NkysBZh036CwceVW5BopjWGYo1JbYDmP2mTaiFELKvqVP2gQKDCfJvXPQ
gDGowwHMediDNDMjqE3MBxxFfs/t1EAYyTSBZmd+wY4fLmgurM9m7EUUsOZ4E4Ww
euFfyowJH8CxItwtdTsS5dmC/SFd432xeNPaM0SPAXVS2qzLX+Be3PGZM2WSRbFW
QCBvFauRJoSwCk9c48thkF7ap/s2DuKKj9UC5C6K11qMj7fh240sNveCAxrUNfEX
bVB88uOAPbO+QLDH9vwqaSmeqfn8qCDxS7qcZzgiqj5tOe5vpniH9uvW336rC35z
yRDXz2kUddWyxxps917vDg==
`protect END_PROTECTED
