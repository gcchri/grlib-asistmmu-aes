`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gDnmPELJ4KPYIixmFxxkVnVZml3YXzStmIgdPZDzVW/OO6/JsqKUIjf4Fd3TtLIa
YEz95WjzqnzVEkLwMqyoJOifsvety+PjFk0kKaZK7wGP6hngP/UrysrXcUubxg5A
G8kRufPkotmn0H/muWGM/O7RMO3B560QN2rIANnF/JSH35mk2pZm2/WikKYCRz1k
SC6YlyXRB9MGT0NATDDw+O15EKKBuvMiRHHu3RphSvwQLTBx82LX7GTVQKf7FhLL
VJZkeyazDq2RtVx5LWnwlhhGwyHvJsSl1ADJeVEyszZ75PJV4XSsEeT9hHiAJ4BJ
kuZ2qyBVuBAOIqdD4y+sn1IOp6E99VYxTuj0/IpsprE=
`protect END_PROTECTED
