`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
thSp3xapt47vnbVzs7dUMy68IwFKi+XMKm0vzm85fJaVQBzpa8+lUzKBMWKlsaiD
3VSfPmm0JnRtSVMKZQVkFbVJXO93J+3smlFiUV1zD8a+S7dt5Gp2G1B+Z3eOEPbc
rVnHQK2wslFmysXXKtAARCRCsZjL71aMHFR/8d60XQ0VStrxeFIPGjJ1u8SiKND5
OmNck7w6+ZfBOyGKRqYpikYVqQO6mZlubg0kCm1RmVNp3TD9gNFCJaWRzHwJ4oM3
DM6uiaP7bAKLKFa1FcbfJm4bnXiTCgvNsmiWudnFhdg8EG12ROhIpJnLT1jjrxKH
aIaWK0NACTWki7xG1mg5lbA5fZu+WycmD5c+4Ep8vaxM+cHK92dT4kjZGuW+cqMS
`protect END_PROTECTED
