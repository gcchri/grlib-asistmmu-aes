`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qCBLr3rJdm2IYZjdNrkRdWzm/6x5IHWwPeApRdEQfche+OKfAccVYaDHEyRhEmxP
Po3Wrv19XronQHqwnjEna3KwYzuUsSRBAqfnoafeJb+INbsf8fK/NZQS/Mx60Eow
9knPJoxOZmgTL3Ifystnaa+mdcxZO7Wdh0QLAE2qAGm8f0BVwWgJ2q5vAll7t7mg
jCOijW/Wb6krMUWK/vvktn1EwMbQb4VDnnDjy58Ge1fxzW2MactQGT84BlPUOeFb
6+COybTLW3BlUoOsltsawT5Kij29m1v86avSeNNnNSiwHpepfi9ThuYwaUnQ0C/o
UbX3jSZ1JwExfNOWnQ1Paw97NSzu0Qx2yaBPO3u/MUdquypivjrJ7Dgq6xV4hGUB
ubWbkdKOFJZNe7hSjsqkC000KlFuHM4L/Bh4BLRhPKlOWs2iLGdZblu4f1fcLQRG
C2Q/pkL3MGOPk9IAOq2DoaKHkLFzAZ8D6yiwxYVzFv+4Gmx8bBeButAkRlWV88dY
mEQMlxsx2PfzNPINUmmvgLXfOhJLTjcQe0bemGS5iMY=
`protect END_PROTECTED
