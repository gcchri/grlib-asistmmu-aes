`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jSfwCHgFFUCpDtnmQM8bzknib6JY25IW6oeJWmPgBOrd6BmAb54+khITkqBiJBRr
01XriduK6tpO4PoOBNxTNkxSEC4FoFHg6+JXKutiWzqsNmed6u8e23yTpXhF5TY/
84U2MQorAUEOMArnn973pFKhLnFNhHcgkJkBcwfjT9cBM+tOqYeSSddFr8G5bjYs
qui8gkHw5zNt6eIIYvzEMzh2yn5EurJ3ACbDTL9+Sh3NYt1ymH/PLpYomNP7bBXt
eRr1E4vMxV0698wxu9MaUY0HM2KiyZMkeT6fFXem4AwpeWT5+16sO0N4CxHskUyD
LUMY+ktQ6rn6I57UAgE3VUIk4u4mx6J4DrGQRVHHJVBLKBbrBfV9edguyB8SN+vJ
ZjdVv/AmwjahMPANn20YiFJ9JlOVt07P1IAEEOM8Cc7tpCyFF+fPJX5p2rBVY/Qc
qimbdOqpToXkT7Vnt9/YZn5xud3Rq+jZN2nT7p2ntDezEN3c3/NrIQcTlbMcFg9F
6esHhQiKMTCIcsTSWXu+llvMzJp/ivqZtxe4/X5gfATCbPxQnlDTqYDVwhoE+fTO
03Tb6ptdhUtprPfVjhtp0bKo7f+xDpyZfOKUx+181FYaa5YuVJ4Uyq8RASX6Uf5L
5ThGcLWk3OreOrp0/cagCt5GVz5KB9sSMhNHhOagtLE3EmS76sHkFzZOrqtltR9O
l4NAgTFw4fwbhIhn68kmK93w6WHgOt7kHM0/6PjKw3pCTJkPS5HcXp+MrB4t0jsM
sV3uWkKCwsKyADKThvICCfKxHxwIQH9HwGAILzFweZweRdTBlecqANf7QZ9LOHI2
p+3q85Flh82/VyTE+stRj5E62g8i3T2nCf8YWmAeSGreHczXjM7Y1AfcYSVugPhj
S5J/iDaXdkKfDttlR70UCCyPnQYqI4clkL8BhsCrg9rK+EomrnUFDblkUdQGnpZ2
iuNNmPc1Nke6s7R+OPxm0Q==
`protect END_PROTECTED
