`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/FSrc3DUb9t58Aw7Ys3LJ0vk1cZRbfmps6KsroV989ejBcqcS6DS2zlGl4zE6eRe
V1cYYvlYxspR1uypfZVtcRMaigKG07hA612wpBb6dnGupkjFYE7CWq5Nij0ybTU8
L9zFms1f5/QE9ZP1X5jkxTwt3hJR4JOTmKpVwjD1+OopMqSPAnHCY8YMimI3fVII
df889ucxwU2AKROijNFvlA+xN8KeqDWkW2omBze+RsFYk4/PPEi0Boo9roxttKAc
/usfYs1D/bhuJZZ8hwe8AwOJr/D6fSnQKB6pEe4ksTYY38Qv6VSlrMRaPfjQgTqp
s0yqB3VD5vgpQd5B6sqCsXqZ2maDR3cULY/j6VzY2oVmhALupb+ttdBLD4K7srjD
be+/6l7FPIcI2xJdroTu5TVShi1ayMqBwlK/aKjrEC77HOdeFV1Si64J72bmzEKr
9tdvHISfcoNGgN67vmpYvhe/RfFVK99Z6UABPpJuO0w=
`protect END_PROTECTED
