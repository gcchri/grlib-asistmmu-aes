`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sQ9//iWXdANDdhGCH+j/UFFnCSu67kVSCMbCDurAoWmqa4hzLCmQpPHfYXcFWnyM
L39DchI4rDKpXd/FyL/4ykcTvzToFzU+iXUJCAiiWGr7qWaUZIOHjQadFdn7EYnj
Zo+L8Fw9cIcRJwYnm5N5o4EDwwATe9yu5xIudjeoBdbkaCyZ0M4nMwKLnBhzbwvj
DTLYXM9uje/kJBgOpfWtCcVEBKycuDvQ61f+YCESu/wpgJsPjWVE4gZ5uhKK27/k
IA4Nsq3lOcbO0loC0qv0x6YixXuFIl8sqmcJR/iOcb5K28fC/Wc30tAhRXPCyEQD
urMLk0FwJMaQm04KdssGGHkNFkR9GFozgCrpwlQUv4EEt88vjAQj0V8qoLIErw1j
nTOaGHZtn/pKFOYtrsltRFXUSWLoCe3pGFE4jM3T1NY=
`protect END_PROTECTED
