`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K5GhPYtn4YJ09zJ5Sm5/XtOxWfyO6mklmQe8gz7QGqWBeizgG25zMLy/B0mPbVXN
8VrbertyUxWpadRie/g8fFx7sOJm5OjtczKSg//poWFZLjHNtSFOqRAfEKzhl7hf
HgYJrk9uTxd0bi82iXkUvzMCx5zm5/NSmaFYWLAw9IKf2xTByFtNUd2vDPFLlE18
Yb8H6qS19wj5xl5ntxVrl2MBtlabGcoCvozyJtygGzay5kZkzjWMvMJXHe+SH8r8
F2ZzkvwYudkxjCIlXH7OTizPRfOJu0nSnqMu7bA1uMx0OOI5o5hH6Y1Pbxx2jSzZ
cBDguW/tOaa0kEsjuuiF5m5gU9EQZmNEQ8jLaqNmOk3JtnQduVV3gmAmrRHK1yxK
y/QlJe4rAYI+lygx8xit4nN7my03pa4mbhnpdfpdubFiDTzNpkZawarRO5EiLAgm
GnmUtHYmweosjbClQbEKFn/qpfehSSvJ92T4NyQNvszyKMiARLw5iHcKpY2G80/A
8m2XWobXqzuk13Cagwwy8MZvFGktN6iRewGv67OYoX+Xdht7PHBX5xVTRvVJlFSx
iUCYEl0jLOMeYnNJhdZ4G4Tvu0e+qxMabeGjF8Uheng8dTMjTBp5WNmbX8dIXksn
JYfY703Yw0IVLQylJ0ykhaxEfqZNfVO1Tk5tQnFRebpHau8gSrxdUMba/4lw+3lC
U2HOzP+T1e5Q3b0B0MA7Gw706ephBK90Hq6VSe0p5NmebO4lvXaeY61PgLyQtf/Z
a8y+QS32zlmqUqsn9qxBKl+sMNPYpTAv1yresoeM6/0RlWkV4MHqBSxavGlAMbU+
L1/4qPoCZI5xKFB62bx6skGCxtu8GbgrhN9NvMG904K+yVkT3+7t4EYi/8BpYemH
ITgyswbChK/AmcMUYmpHHIh9S+B8zTEqrtf3lncimWvIko2GUvn1OXa+E5Fah29d
`protect END_PROTECTED
