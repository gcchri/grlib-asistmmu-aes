`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e2ZYzc0BjxsmWBbgw+PllLdjTGYy9d/D5Vp5FPM9XSKUZbhgirgXLWQzD1EESjQx
wtBYbRqcuGFTdSEU/0wyAyAY6LQqSI07iRvjTWNfmG07UaqtEsyROEFSYmmlvNbe
Egv4AUeatyedkpHuMQ01cK+c0XCPRfsa0Tp7tow/ijMpxlGbdu8JVfIPLWa2SgXD
NKQZaNeJejiPk3vre6f6G5H17lIkf2KFUNPJqzledVB6AueuGCiZsHBxUsJbt4+D
oHCw30Kg4bmDF9nB3S5KIXAOI4LHrSW2sF/KH/yPTIQ4YWNuSUkLoLfG0rRh72j8
b2+S46yNAiHP1YPfgcp5PBoLVcB1CtrNwxoff10Bt/CL0PY6f6s0l5OmQkr0jM1i
EnE2jpKf30FBVdyB3ic4VdRJnlyBMBQmvf9ATgoko3XLDBuh8HUHhZ0/ruymEQxB
0GVJTh98ETBVqHFZ7O9x3UzvooU+vcvTde5JF6GCOE0=
`protect END_PROTECTED
