`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
quoGGPuUnvr6BDk+y+eJGNGlCgJO4N5zQsfIurThTjP8rQu+3KXqdB3gdiQoJcP6
85jd81T5iIA5Rx/i51qODN/J768FjnYnAmqC0fyQTIKQ/KJnjBpIhHWTbBannDFY
ID5WGgdExBYN6FwJy1z0keJejzirCXEp6DMZfQ7SS4Tfux5sp9lu1ds9YEgHDm6s
hEHODfXSic8/ugnrX+KJJvV8CLjx7wHx9vhyT5TVW7Cs3Hqm2ezfsvkRIAsyR2qd
w7B8xacAAYYTPdxATMurh4dTQDPmVy9hyMnBxhov4fukuo4D3rg3JAOisDje9rnk
OHxOTJsr9EmhoMZoc6oSVg==
`protect END_PROTECTED
