`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
871WuqabS3m/ucQDlXx5pOepgsB/RLk6WDqnku+E7qz4w9ug7fzy57Gp0TPWdQ8A
aslTMuSSmgoLkrq2GPu60VOzWHUVgDCV010e3Ex1Cz1ZviP/bu3G/VrNOfkmqOeC
iSp6mETdMrnkcJE8M9rwCAMVlPlA2G3e/2Hn6yM3kp//9y52OMSHERsLfM7RQzhI
Y3kZep6Fjy3i8j8BbSe9TtAIcb53LjkjvRcpJGr9y45jO6Q8g47btZIlD3obuH09
lxhe7HRF2Zzup0u1NFXlJnnAkb2tapY37sXBVrb5Auwf/pBWREsbaoCJSrSpVWtd
y7hFKFfDD3NRN7FAhqJfo/IhMmknrXKKP9b3Z46QgSpFlPBe3IBYw3Te1XZaGDdQ
h1HD/+acxZqaOquj3WPZm890U2zoACspcrQjx6Y46a2KFtuMYI+r9MVqzYDRz1sz
chzjG98KGEBN2J6nQBW/C8AGJTYMCpqYx2MGlyEljh9bv3XlxUjvasiUm35Q9T1c
neVFxtweaZNJP8jHWWjbZSZf/Ffc7RoKbACgtOh3F4pVMUWESGREaXrywr6oz5Uv
3Is/Gy+nCz5XPhY5cRw4Bw==
`protect END_PROTECTED
