`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7vMzN2yxooiWe4gu8uyB1O3ed2RFdLvy5zmdmXzHMv4qxso3zUXt8CtNLZ+iRdQa
8T010+DR0eb+6jsiobrZKjMBdEELvnIvMTiHKGk9U3tMPeG0sSN2j+VfDujqJDwb
L4+tK0L+/eKuZSt8v9VwIoBbNgCOI7sfH6uvXcp7Kuy2PNVCxgN8pqHMDCpCyVzK
tQgPvBCwKxsSI0+B5y829UmW9Cn9gpAR4O3eEOi/EY6bmpgnIQ2M5St02twTa39G
jaCC142Xtu4pZRbH0X43EvGVeQ2HQ2ikB7KnUFBR5/Z2jH3+fOR/GCmetv1yxnSN
IoYiUcON2fuhdNyWwggFJOQckOvb+PiWXTaHFamCUSOI5IFwhv4XbQKDqk+MkkEV
dXLGqSH8SExaoTcR5bTmhUgInxIj0aFTkq6jnOpnLxD7a8bKR5OSIIFw1Kbr400R
mxN9lq0PQ8PfD1k4QNgQurQJsNRsJ/aag6+jmem2mfYcIGFubKTuhoGrUkeDo7Oa
`protect END_PROTECTED
