`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BjKLHcZXQSm9uZkAtuZt/aoh7ZiDFUHHN5yY8nhkF0sclU9a0GS0ghZG8NdBKwpX
Z5KWzXLOqbxpffTMfKS57aUS6qQ5T6D2s+MRxUK38UW8L1LHOaVrcmT7R9+VFlNw
yYYIbu8zHOYc2O34hnaHBVDTMkrB8jBpVEGY7UEGoTKsvrggW7ERpoSJshOfkun2
8aFW7bxwnNYC/Jhy+oNlEzsQdn85mH6trz/bj+f4tn/ASgaNSe4pHLM9J3lwwMkT
P0vsUP0/WtA4mOxXFVQaF9+0fanAPIZyCO0h7BDd3rZPjXTHcvgKzxUZSq7wXjXJ
6/4aX6l5gPW1+LK6nPTuV93oN0P0sDOBh2FbY9FFEIazj5yYlbQ22hSPk8NzWYsj
tvIYEoPgNMJTszCGWPds6JlU7p8oLtUhNYtl87saavO9vxnYwUU3oXA14rh9qEnH
vgqHK3aG1zHAtBDe9r6YmcGPCAbc5mBvLqPhuQpo7UM4DHA602Ry6mRuUZKlJsiM
wZSIMhLqiNWRs556wvc0pA==
`protect END_PROTECTED
