`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jkGyaDlfxwqhwbDeXLITfYcWp/NIAujCaab8YU/NokQCF/xLpPLxMxm/eSpnuyc2
OK3QUMNahJ927uH2ZUM2X31f+EI2k4i901pqCarp1MUTdFeF+n4qLWbbxGrfKmhE
zj2IbcFy/MzjGKXkRbE2TXVtTI3cmYWqmtuifN62VlxC1TI6PL+MOg1bqRxCR1xC
shN6H0Dex8n4gFiyR5QvDKDc3Dm+37H7lJ67hL/GlbzbKS9PvAJfI6Oh3cIS3eYp
t1Gr8xZMRqygkMn0EkCrpJfBwc1tlfP/fMGlp3NDn84nTJLpuYn45cbqKadT1hsy
Esvgz0twECYjLwa4ybQlfjIGQ0/2cucfEIPxElOhSWtqFuf2rTR5sP8y+D8d1bUb
8mc8+QmefqCsakVAzws0SDT1hicDfd3SLpjQZbpV8og4f2YHTWu2ovuxnYIVYwsG
XvHmMBA6UI99wgf6rmUyE5kZOotXXGpN66QHErMCFkT1fLvw67gZ+57hh0ACupx9
KiBxBXGIG2aakxvz3tUIaggsK3a8uuSs9L8pcSX9qMrPXj8h9l+Z/oxJdg0oz/IY
O8SzO9uepuhpIqEGSbAzcud9KZAkv358gpmDSWZNDlEde3htC2dko5nLo6aPlHQF
QradRgPdg+LK6dKOevQsU7Za/7HGEQxb7JJoA+AjA/JcMwWHSpWEMjLkoZ5BGfo+
BoWywouEmn9MZDZekuEN4Qs3MKU0lyN+mx4cDUUtozoHlODZjTramoaCDjcSKLb/
KvkBAIO9MxXB/JOh89GD0a3H7IJZuzJGokcuVlxur1RloiDK+a+gVJlbJl54oob1
iV+oPzyU6EHlJEWe17qrWgPA4DqjSe2PrLcKKST6sASbpg/4FjsvDhXr41PB09Kk
NmDKOmnEYoF5SX4Vgwdcm7mraC9B7J8MtxiK1cSWFqccrUgzMV0knVDUZn31uOoV
X5J62V8tHKOGzVUXEzI1cWmISBLuZV8qAIXA54w0EVh9VaXAitRYRZZal/ZcF/tG
f+UCzBRLAGozFCMlnLWQvKXGV6BLqY4tRvIElo6ZghP4hGP5+Lt9/c3lcqnuoWam
+87QHzoq1+SOhFDvTW43x3aPurLj+XjWRhr0+xVCA9lguLI0wlpO73Ii1S+OkpWs
xLG4FPw0HshOLMIQ4Ajw7g==
`protect END_PROTECTED
