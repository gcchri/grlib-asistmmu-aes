`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UD+Nluvie16RrdsgW1km/dNbR17hxyYSqq546cPBcyCNtpPUDT4VfVikcvzKNCrj
7kZ4+7cRM49DvVewTHxaOdCbh8GZrZC5PJ8s0gxKxZVQGFdX0TP/fJ6CzuxiapFv
Sib+GlJWbGSg7UU+PsTZuEcTxMkj4Ayy4aWqChPp/5YzryCmzIwIcb2TFVYA6v2R
trcu2AuFFuMT1k0QGYCxmEZew+iYW3vPlMM2UOerzmY33YBzo0Y890tyTOIx12MK
eBQMihVEI64/efOavjUqpMOoapXyHN5/nmMDQuIB10LT+Pndl/rW5xFSStGH5s0e
sRFzdCyFw+fhzB0PX1TeRSou06w0FtsPi2AwkxAvzs2RrEX5zFAu0gnxEUi0WDlD
YmMbC5/0kytzsLXkfFJt9yRYZhH3VhoP/Xa/e16wI3NH3Chx8Gf5yO2jUKRv5Fyv
37FEsb/4cXt4tnTr0NJiQmpTtMkgkOGyabFgcFM9tHyOG1wSZaFCKIwZOtwURbad
DYIuIfC0kP4PkBuEnUP+ysLchtEvM84OP1vsSgYNYoPifyvMeRdC5DPcOexktY44
rIk2mH1VJuI4z33zgBO+TVQg8zec1eWOQGUFhJiY916AP1gDJQ/3/49wRo2dZ/JI
hS/CiecAn5O9SFIJH8W0TQ==
`protect END_PROTECTED
