`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l0Mt77DkVlCPSwxCIgM6p3IkM2H++uXRi7B3FB4VtCa4aoPiIwnu5p5mSxVchpyX
VcKraG8o7L8MwgIAdrrOM7AFKnm+K+vVNUCsB5whweZbpgwizDb+7FnrJJRMWWWt
ysuxHfOQyVs68xWd8qLqRdnEIhqPWJx+YOGyfanqFYU0alNoY4eX9dLOh0veEJ81
zkfkkMPRd+z+wXCwtypHT0L4o/hhzmtz31LMgeYQzgB9FoI1ABZBqjDM/IS/M5kz
p11T/2h6J2OETfnhXXIoPQNB9TQpdtUdECpqv2S3GWImRJTuZ5L57YrhFt+2Isd1
6PfxQcE0L/yn/RnzIj+ys+UMNlsZky0/yNrLH5QyXHJJHghVxpEelYvPTAM6irSG
ayvdgazk4LIqpGXUl3R/xZrHeqqR+wf8PuxJtDW4Dh4st/bmVsUXQDZfwHoMVVj9
IBdHueJr5zLx5t0xDPOVSY+80fJxIXBfJnT4pJkZYFTDI1O4iX++pcKQ8jNc9RUk
F19giqZJZdfqLEXPvU9s1izovrQNvaNZ6tOrZYOsZKPkacTBPFEh4WTq1M1zyf5X
1i1ewpoh/HEm3hXigKT9sm4giIhfAXjUE4Ksq4tYVdG9qorf9L+5lo3njZIbCSCA
FhmKs7pfNJC8qH4xhyJBQw==
`protect END_PROTECTED
