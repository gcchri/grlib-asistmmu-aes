`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2XUnUroREiZbbufzDaNaIE5O//PeHtfVYcC7u4rxrBssWyT+ySGp11e/gLYJYf/f
mXf6Gx5OGyaJuFdtL2zD95Zwt1ASMsgIbgJJ3Nx+w35JNn6Qe/Is4ADbcHVHmYzJ
nju+eQx0mpMUM1kuFK27u6Tk2n2vLFOgBERYG6w/HgexWnegaPVEjYWAsL+P0Sgc
HAbHpkGopw+CIGtFuTnQ/wZqIKzStJrZX5Lz9l5YnBsdRrFoPFr2Uxa+jN9CPyjl
1QXzsHDnTKOcZx0Ow0P3HLbCPupXj4OxgQQwKl9EkPhXIGRtEkT6B9V4edmehIWz
H5PXLmc4bb+hXi+Hivc2HUfFDtUyRYWnZtNOrQzF8sHT1yZ1NHGnJQcgoUh3uZvy
c+gsaA574dJoF4rSAy0NJhUTrl2qMq4tU/wgIjcmu7TZNiQWi6+jBeqdJdPeFUF6
dwt+hIS0HQVD3KcqdKG3I38qMmico6KJ+ZmHRpVu0uBmggNXbFc3VqA/kARrzloJ
U/T/hg32GF2wW8YaXJvIjtgiHXAE6a2/q5G/3yKKATHa//4mfqUWGzyM714zFw7f
UntzefPZAAKODhb7A4bqV42f3ePfgbS0WgQJbwtaQR0/U4jenSK49mlZyzcqHWny
8ooDjpa9QV6y/O0q0MfQLNcRqmEFbdMTaDj/UywrrBkz39Jx3ncAuoDEL4AF2oI2
SrEGX+WjZ1AtrJHsAxF0CIYgg4xaJX476jCsFcmMHBq688UTNwK886Do6HG6bk33
CxPorKlzyLID6jncM9iYTP3w3fOeS2LIsAUPM7NP+aClZYo3I1je1+NvspA7HVeI
Rss8fFPOqRVi6JPhqz9ePwd0LeOjevHi1YdF+UZzSxGPYrwRMvoaAICPBw8Yi5ak
ki08wOK/MvKqNzlAzlos6XsUeuinqR6vIPD54K3qvJydmAtu6sXdndwqxHmVD3Jp
fQKdI3mRsXMO0jpZVYDavmewLPAGC8r9JmmXL7GtnzzKnhiCnsM7xCnT3JUbXIV2
7JczktPCVDWSSUkTb0bRs538UzCYllF9eV6xJYCTvehoOenJcekm1D34qTGwfR67
jCnWpQ3loSG4JjionY7QnDxDKjTPG5NikhDvb/VkNmLUhUEANWxhLbqQaq4ETYll
XQk4Iams9NPgRoHCrw+ZT8pLO8utY1d+ehG2SeGG6f3V5UGYS1Un8ZQmlbJtI9+G
zGADWQMPuYSJp/A02CoyirshPrz7GeCVclplxyZ+D8yVZZYqFqcLRIy5/HIfyjxF
0/EDgv8OFdRJBUCZUUeL/g0aEP9u42BNyJ4Z1/qy826ls0VHTWUiVylaHLNnc109
cBqWmif+Cg83uEecik0Xp2d3wt1MNaXKrHQt2XFTIowd3PPACr62ffQXYIbsCZtM
COU3QMrBYMyVWvO6CjFRDI0zXGzx3JIeiOHF3L/HWgH5ZPIXGB+XmXDxjCPBrOXP
afKiJ9gH0wnMAwdjl6PwPAcJ6MWaK5eMXPOotcXEuFD8XVkd191E/2CRSbX7Bqqa
60/fn2tOL7iMpHVU405NWR6nYFqpO2+URt3PYeQJ+0tCRyDyKC2VWRx4VhPvL36R
uxoYSNTRKNS0G5HLic5/IEHnr6ZQzux8d903A0aoAAS06+ji8iqOloD/RvJYrCPo
PEAg1dBTYnX2uGTlXfYIHRfLeJHSAlFVZi2sFJ/523si96EKoZhFcO9FM2FuX9Xw
8S5gatoUQ6v1pawd7IzYcDneSENwrPqMB//cWISfVCdSz8tn9UZC4YC1LoZPFGRu
3pmjppDkFm5N49LdncJRm+smtOxNt/1hgO8RHcJPo9fFXx0k54iOFNh7EmWJ/tWS
N7ouhXGTiDDBIuFj2bX2P0ICQLfPIN8zS2t70Y2l3L49drvReU8e1zmGUTExMXIB
9iBvHjYdmX90B1FuCyk4mPLF81DBdopcnpZCZd8K+U7HzHo72rBscfsNWLilwBs1
S8sv14UBhSGhjhqjqkQPW0Mt3My4l5BGTLmdF/KMdF0xOPpkyQ745By5nRbkvKYW
Ve6iFyZnrHme2Fmzxu9oO7GpcOO0dilJ29RNLL3tUIPmtsrR/rL6l+srGrFrxzE1
PGyt2dMtHITx9Q0bRNiB4Yf7Ivp1U8WiobKIJGvbaTGWAwcf1KgmJX1f917RQFDQ
tB78idHAsQw5/ckh9ggsR4l0TRaiaXTw9BsugZJJIb84uutKnU4W5CeuCzDZnWzo
+J+tX37pq9nbn16S5d3Jj+SclK8p9x3C3rwMTKdXQosvRjRDdmPQ5liqSpDjzQLK
xmhEiULOpKzr6Ok16R1AKaxUNLgS3IYXpxCUjs2UcYtL9xit1knrEsho7mUjsNyO
eMH9LYeVYXUXHIZ433CQE9hpNDYfgtF7SXap778RNHIYGNxD84yTw+vNCXUMeyIj
NPgEF6JADmA+fb6HfBzTfmOlG2VdN2cCa86c+FwJhWqLZN4F1pCQPVsDvpmWAx0g
HXskcjIGZ1GOE1XdPxMx6KJWZ/hSybrb/scwnX680Mf9TwFB5bBDJrFRpagvJiDb
FWyHlBTkXsHLuynGWdZhMhtmdWPO1sOkyOqXJkeUDD63DZLipJf0qotQhVXxKxcf
ahbIYQQ67dcJAIeQFDXDbObNJmqCBGfpjj+VZS5MRWy78Kk0WoTwgNtXwZIu0TEU
x7cectd0UXm/t+g71A0F4De/yRKd67yy1FXSH/hrk4ncXGO343SSR89PGkFswDcv
Hco46yZ/+wuP4EkdoeLUeSHTe0y8QWJ+xiHxW+6qq5ASIr/HiMh/6x4tNaqzHP5G
Xjme/vITTscV2Kjjn2lgYACIKAIL65SMOQ9wBiTYOrHKdrVvQbC0L3g/sEbvSmik
Iw06PDz0/J5O1SpGoxQdKV6v9OLEzBu1uLnW/hd/4ZPNpn+7AUH0aiPGtKvRUpY0
0Xmn3at2oy51IUCl1tZ1CbnBm4PhwLiUvzb3MF7uExSiryGPcYYCmkzwkWZOI0xd
eEm/Rp5mUyWMZ30Q13XCVR9pFfCCyFY9g965l5GVr+C/Ra+ParAhAeFnsdJnuytr
DiAfe4qCf43BA5BzEjdLkq45Sss1gv7OqGh/rXRSnStVl/gLc+HhYkZLggHo978s
sh1Ij3nXR2S5FtvrRh2xTzu25aUoGdVTCCDFeVumZnLKAmCT/TraQnzVNrU+EOya
7tDHBczO4NXFMl+Ax01qIzrmNOLHiSXgXVef7zCj4Ko2PshP8rPvpn47l1eHN+rZ
2F71WRrHHRBh8GmUhwNO6tOzSwxviHLoOpw+avzIORzECStd5IFiZzIPIHlgyHjl
yLI6Ab8HK28mTd8ZTrbSCq7fNsD+6SORJrACwVNKhI9U3t7uqabScsiUaKHLvlcw
9xsT8x9Qb3C4DnZdrV3tDyJXpLWUq7JdN/zkA0tgfKiw26T/as9ynLmlEwnNtIIe
DKLYurSHKIsP3W7G3A3gIEB5OQI8Jj4Nkeyemgy1DceoVPGBruBxTgImTTTLWrUA
ANv/gYSb6PVk1it48wrs4oL8IzPXZr5ruAv1Zr8D7zfHQJZJcrHRd9xTUXjQ/Bsr
cqpT+wVd3N77sStZlRhOs1EkVlrDt8N7QUsH4Lqz6UOU6saOJSr9kKm6WFLTB8RX
AnkXX3J2jqF5ayYImmup8+yBI/sS7yd69PIVtYSse4W5ndpkcW9ZYT+N6T6HK65x
hSUMg2YjaTb/+S5ld1TPslL4D1XFnXoEKq5EhtbNCpsBpmOBjtpWg5rJ4W4bIT87
ltaq8D4J+zawvm4s4skJqhyWAatCKYiekRFrZbmW1VEHB77CzW7pSqbsyKSvQCCf
lWnJv9Sin50mzLLJs/2Th9R7OlSIrIRC1a9ee9Zm4X1QCoM2dELQAN4GzYwX1E3G
GLzAUEedgmChLLAjnScjTE82ZjdxTJ68PHSUpr2/ytVsK5y2XSI6pCAHovq5852n
cTP9e6b0GhYdLPMDgJ5EkilatoomtsU9mcezwY9qso2ZbokNrsK34ibmvDWDGD0s
ZjeeIIU62KQvZewZvnL4+EiAuhP0JX3lGAqNvdUhuNp3h53i+JUoTvTw70HeAoA4
Syp7vgvUXWcH6A4QIOkKKZZpBmDosHFSflAYuLoYKZn5FtBwUWOYStBL85TNKiwv
G79uUpMB8se3mM8K3IzMB9Psva6JYR1Ibog1+KUrpvRs1r/xkCPeUzi0lt7cQq01
trtERpIlmIVaHny0wq4hj6HdNj04/qAqjgSq4VSYQBdUKrA7tvp2wPPNp6qlfPm1
N5J9liHkVmBj/TI3+5pn7+JVKhdYdVieDew/44aGIVcPK+eIdJ+cVLo9mB1i6/iD
/mFRjBpnhEFYh8cYTQattrktlsHPc6WfwjkIK3KO4o8BrPTA4nwIyhbkRFL1Ay2E
H8OPLgAt2NDQ0U4Yjgc8gTRTVQZXQUjMK+hp1tQLWrEQyWEdpQ/o9Xuz3Cn2CB/A
E9mjcU4SGbTwkZqCbURcWNpv3MA+p67pLwg3ZvGoOUNNnSITUr7wyq82YbuFpjXs
7F0FnQpGbpvOW+YIIQqbKYup0g4OzJMAseSbcJgaPg1wfVuzNXHpzSRKEWhGUfXm
ZrnQ9gS1+/LsA7pxMw/FFn5KLwCZ83SJe3j3fEc+RjiGplL4Z01Ae9NKFJ3NQn7P
/nROsRs+MR1ZGq2Y8CYXSTKGU6QpmnEijzL5PJ8wnR4flzoc/RlXQaP+c8RGHYDg
uT11wo/u8eFW6eLufNEK6ES06HLbnfPfAo+i0wtbQrmKp5aWRECpQaqxOwDQy6Ke
rkgLzSDs0m35eQA0uDt3Tjs6edgTWfx3DI6JyccXgXuOyVsgtkpU4/Q8W3W/KOBc
P9DdJVLLMQT+kmfCxmNXnGUxQOhKl3YJ/Pk1J2gapqKnU9iUyZl5zw0eKu3evcxg
CacllrVV4c5hWZcbx0FS9PtpXXjJpR8k8zT/xSgehpXcxHK97e/zz39fnxIarKOM
6z3nsfAByBZeWQbG2gRQvOIb9KmSm7RKmkfeV7fCRyu5jqi+4ioAySp81w/Ah11U
TU7sG+QXQdPFf0w9w1s/NNjE8skJSt8uhrZ3RyhastTbCUSn1TN2gOXhzf0Rn98M
WXCDNnsTFBjJ7UD+iyNtuGwJWvhVegDv3vRYe/BmbF0FyyAN+HOQJaw7g64F6gXZ
Gdmal50Wpnzoe4HcKqD+8LHHLIT3UUXF6ZXuD/2tUcbtAoT4bhoejSCGcbP5/7Bu
TQWBLsrkXPiqv385mHQH6VgIng443waeem2ZUVv/sX5m742jdJKShx02gaTXlB6G
pMC7GFS3hTM/TFNDTGOqqNGzOOep1ubf6x3pAuGs/34GkH8lMQXGvTKHvRaRpxOu
ZHb9VD3TMh2VUhwVjBRJSMqBKAU0It31UFIJryc5CXpn1FvIpIq0bfpzZZKhE/p0
FLuSU3h2EudBruY1kzYEpfM2cxppRjqPEUfB3zC2woyiFUfbxT/XMet6hAmdJu2S
y0KtUzAmv85kf7bdlwXXRessxMiLHMmEOm79gXaqe46YDCHl4oaWfxcZ1yXxhkg+
LCtqCnh053AVL0skV242lb/9DyP4yQsvSYVOGfhOPQvxjGjrqwZoBGcdcaOypsGb
WAwkFDCY7gzeZU/+/Kj40/LLqjdI+MFhYnaX6nGktVbpvk7ZCMcIDJAnVfBZP7+c
BBDExkt3C3dN+aiOuW5h04I1ypg5CLSucXweRuQwthNRELUr5hnpT0dHuFsDNQGf
1ZQaL4nf701tPhjKFo3NqSMqHmUgDEmbodyCn6OEW2Z/BJQcGL+GaFqf8SAHDIxC
xdu5PpGdTR11ZY5ZhZjOzZDzBbVeIcPHrZX8kczrCHncK0kv2bZ10pUt3nrVINZH
0PTjacHQp8pKi2rANnu4q/iMnkKD5E3QAq8f1FCKoX2SdUNk/3kY6yPJEbSRrBPR
zGuWp0VWeHeDxIRSfwh36mGukOXd6d/5zw93QBE8ZOdpMkDrL7NnR5u07vG8xT/5
G/i9EHrZpSnFAeILFLOQIKrEv5kd4zQZ+Pqttlu7cnS7/H34t6kuwptzKHVhhKNQ
rEiksbn7kfzXuq1M2pmE4Qbi+OXx8X6NYjb0cn/yoCM72JavBb8aHceT3a2Z2tsV
uq86p/B6RMvjDwZny1kasfeqtSIbiXUhfE4xx7G3pyVC++/9bZP2PDlBRK/C41Th
nSn3cABrdKF0bd11/Tqvr1teoVYJ5jcrWWAYQrTzZvcfXxJSPsChCiZXzZwhoHvt
/fTq546uggSKIt3RbwFOyxow18OsyGtvZVQeLKjIBhRi0WUpbqTe16mL9DMK1yEl
sAOXS/Qfx+VPgTWWWm87nyfJ5jXFchOqFWOiT6KFrL/tFSJ01OjIhPC0u9VN4aPC
ALjsbCCbYJiJk7LWmoRsDeE15uDQc3OnDhPj9jjabXJ4DL4VKtwZvCicfEpjRHF3
5WolhV6/yotrgjC8F3r4hUNj35af63oDZ9YQFgkt9BdfIDTNv4dT5zlEOF+SrwGq
M3GUrBXTz2V6gupM/udb3OCrQpVIwLykv4Ec37XzxdaB01XxkhCAtAdcn+nw9aVr
EGU12u1e3QoF9RJjaHb8XHFWtTr90mriyqpw8VXIiKHfB1jpE9kEpmaWoaJ2+K2y
gI/PoI0mEJJVmN8o1S5WiyMRrXk3vjmE9rboAYUz4pPuTmRXF41uaneH8ubd1JF8
r4EQxOE9IU075raAkIP/RR20Sc1ArZgnUnCu5YZZAKkouzhtAybKhKwEnhQThQh4
4zcm3/9vi1CaV2R/QhMvWzVAWHoFfPhZHfPloI9X4fY2VvaMfs3jmqyM9f3X5/N6
JbIFt+bap6IiSMHkVWww8ApdILXuvxn24F6rZq0/lsPmubLM3tztXnN6LWFCbSec
x62UaB8YhHB8douGCFlZeCmYOpS51/ZbWuGSMzIz+LUAdboBj6lShgkNocRh0NQB
CxatZy3oFEvLasEBVL0wBUJ4l2owp9afEYfIbB7f8mRQ2a2jW5vMxlSHldOFsNNs
cGS70vVPo9iTVFV9o2BGi0+QVz4mRp5FePWGAnOGrBUEOHgvV/WJjVyVGA5FjD/V
IZpYcDiqIFf/KQwUhYdJqwsRS8VKFuJ6aKDLtUtds03T7mqjKqQTdjxYXCYUh4k/
TBLk7qUOxj21qvdJuTGqPLDz9m1OHOIx7SRo4DeC5FOAUF10SDzVZBxXTqLW1xGm
j6Nsv/7BYyRBTiEdLJwuoChGbp5LvVeedN70ogm7ocUAl85HKpmbMesYhrkGHndl
fzjOwHs+wo+prvxfkG6sd1FxLScbgrApRtlaG71TLsibBYVwaJGQF+eJibeqe03L
N9iBCi6NiHi+oo1Ef45kWScDBfBPtR4h+aGlAHr11uCpNbVVtE/vluD4t6hxwKqm
CN367c30sKN4DAyoHc+StPoBSwpZ1xVNYUqg0ZEck/FotFJYoq3y7EVw/gl+gYcJ
2sxT1z9rv33dM2y8TR70E+VvzewZoyNixAS9V7GPtcQvlM12Yt73jtIVqCas0Coi
lPpHSp7YHeKEgqXvKNcxpDzLOYjFSx5PWTZ/YwlMHIxSgBq/5nlR/dU5F7f3dKqU
WAVvQOR6o0Gq6+yUvUpth71qVYkta3tDmQjuhDslKqn2VIN/E3oXbYsuQUKTew4L
okRYdCAh1fbCH1j2tkWaK/q4G/B+7Rb7QdezQPuKXkKB44VaUkGe+PgC9TPRviyw
KuIdKavTBz5WUWRa2QO9vV0X/6pysyQSER6ekyS+ilSMj7zSoIeq2M/RwNbIrcoV
SP42UbgmkOQM+dD8ERtGf9FZCHHAhQijdE30MipkLmHY+NLybKhFGmE4Gk1m9ECM
egudUw3pKtvKMeXxujWEfFmoVewXHAllppJdm/D/xAIf9K3I7JeHm/SY8+3JbZNG
o0XLbQLKJREVKepw0PEI6CoVJlk5DLdwiasYLUfrwoPSym+UjoqfhR+R5QzuUH+a
jjOsUiWtYIvmE2HJGhnzjZboWjD1KtMP14wvF9JmpKUlkHxAZcDEgjeZMElmLXI2
lXBNVVhaLZBb8R/z4+lxWtk60m4JzoTxC1KLqq/xha0kQn3NKpm5onQNZSCQc8gI
oIDEOxtWL3uqi0y5qeXX63Q6jm/PLqhqQKJexm2p0ahr9vfSN9mtGPVflynM3ods
exz0kzi7C5n92+hFxuiNxBQcEUCaN3TSiGMtOjI6KqMtYPmLV+l0vui9SmXML8rK
Ic16ADX29IT4cHBAXBTLoIqJsRl0wtHl8iNkIOePBzAt6U0PgSIINVWkkXsLr4Dd
iHelyTy5yQP5ZTB7qDTo1yYzS08AG+Mv4rWQaMWglkSRyzfu5ycIoR/WnF5CZwpm
a9u4BYM6Qlovspz8Vd/IcWPRf4ubRqFdQ4FpKypxP6HTFv/wxMrpN5wsNM5D+4UO
YnJrbXuN43Q1I7EI2mIbP18I2YYqR1PrbJmNO0JCPkKQB2RPXjIiok594ZIA6/LK
s/2zDjzi3XITJ/D1joE8u902LfkoewvaFxuwprZB8rvcvh1j5RbCDwavXK2sqWRI
d/puEtPeGxRurb2a0Q/kLODbkNtIUDBiBO1WTvukL38f366+2IFcetLR2X50FmYt
J06QpvDpYAsA3y2S1vesLHfVirffzKt5sS+3uDsV37uGCx3JlhsfcOhyzAeIMD9q
7Up+9d5A5HA97cX/kBWUqY/E4y6FfLlXc0aTTXSl4UmcrQ/Xqf++GUpej+UfFJ7h
9AZwtOh+ximyAskc19dHARt4l6BVL2nCrM1dEvg3UYVQqeFptU7NSgIgtaJqx1kx
KQym1HBJYpxMPR0hLi+KoS7ffO8PgwztGq51Nyxvir+G/mgITUQgDLNM7sljRFJE
1HHAtWLpNW1HMUIJXjYbAfypj3hfRhmgFBNsj1Z6gPxvjfyWsv0/0wBCxqsals0K
TrI3tb78yK4UeyHQgTGxkPEuos51/NjtBOAzatnIZWMnQMwlxwAUbn/OplYVtBVL
AvNrFogBd0IVwDy3BnJmwxM3Fg4pBVsQPr5EO6Nw2kr5BqPtoN/IZ0PoKBr46A1o
NkKp0BMwb0ctgs9fZTLgtq5CblteCDJx3BoVuyfuNJbyTi2CMtYbMIvUgNJ6OT7a
64n0xgnUCDjgmfqolGNS8gV6ZdYmKY3+2ry2KXuZBUY2kwxeuaNmxBUHYD+r+KyM
idq6rim7nT048/msydmHb9o39SblqyrZVvlOl9YzPOfoTwAaUfydTQt5pnrI3Cq/
KkTnl1+zp2VSalM32KgKlZNYm6q9EusK1B+hegeQzdjOij3Hc1exy3Fjd8AlJYkZ
aNdsNL1lvHHD5AhERJwrjppnoUSEY/7XErEGvMaXSRVA1AnYysjmHaB8tDkD4Zmm
7VtYIDgw6jbhmTv59O4KnaKe2rmENt1bhsFFymvIGSmKAuMlHM4LAbpp2K4GZFps
etoKEj+L9HLjsU0VAP/MjDpIdK8pJ/1Dps1AqTZDKJb3qu037IV3nPXBVES2eE6r
lo0SIavRSIouGMHb1gNzqzmE/YKpCr0CrTQ/CrQTrjaRxh37IFoCTu8n2LaPukaQ
855ElVNdNSK2axswXZ+1bezSJ5nGP/uZ0X4uqXffFQtKyPdKEN6UaI1RsEBxweFE
Zj8NHpzRIH5qk4fZYyd/qTlpI0cyAa5dl07Kl1ZUqSsKLnlNYCyvN3QXhGM4aSfH
ifjMaj6fout9zsLXi2UrqcJ0AxSIzYcuvDW/ZBNubkyczA4RWf7Cb7sRRHGZ4DgA
2raH0/zXESeb/n+fyOzoXwKvREinG3Qj3PlQS5GJNY8IHEJrTsLTpWb0R+b3BAfZ
JIBpuApbaPWTr1p0g9paq9EAHK1hT4R8cYDkmzLm1dOGOWCgWHxKHzFeCs8SwOBg
1GAECA9SoDDKGmyMs65tXeOWgYVbNwL5u38loYQykcDYWFn1oh50aSHAfILFJUIv
VRebStHJ8Ucfax4SZdcqyg3CDS3GUz20FFkwKcEAwhsKydkTsfa3UNzlpPsqrlZu
rfw6VJuUSDNXSVTIzRfW8nWh7VSg1rsFUPWwVNRLF1hXKcOVDWs/E9ypYGCfrAeR
FOsEQDaCEnijH2+3+SiV3nVHg1B/L3bAz9cfe1XjgE+qmFqvotyuT5rOuZZiPmDB
6nLXxjfRH239EyO9Y/NXlg4Cv2d5nEnsmCJMIf4n52+5hMslpLMKISzjJNdPujZ7
IeRv0Wews3U6iyuI7eaePgdp46W9oVNT46HRgiD7WJNj/1WWZdG3qe+55AiV7GdD
iNJJY9ym4KOg8kWN0RTBZjlo30AzEsdHPWbiAJU0qBgbavbWH/jBOPPQNRoWj4Cd
3OO2sKn+Dpp49xK+UN1frF8lYvBnz12BJhQecCmLSV/xJbzEdHcS5BmoKC3VAt57
vOvVlXpztqNEZdN3v453LeWczso/Pjnyw0G3Fq4+MHR2Z9AOV1EOfih00fDkAizd
+NaX/VsVGR1PvnKoVJacr7+2R3DoMr6Zd2BODBfM9sGYH7GZjDlVvv7XXck/cKzF
aUKbsid0tou/9oyyiY4H3nnoy8sZFa7dYg0SoDaTngJ+OlEi+pPG7Db2u6HDGmzc
w1cfOnBT2S2Isj8s9s3CPXkxCEY6EIoFyYwjjNE7PiscIgjhS8tggSx/haGZcQBw
5Bix+6EeQtRc4TB5qdVo/sWIHboadyUrgibdKyIeu+8=
`protect END_PROTECTED
