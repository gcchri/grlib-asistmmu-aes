`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jifo6sg7f2cfdg4u4fXz/YM8aploynvY524VHWcEBGd7BRTHGlv6tCe3o7k4LZ+Y
C9eJG7jQBE1In7ETr0GdYxeV5VVuo1WXIdJhGaOUU3AbRsuF0dUSjPpqXPnniJRg
U9W7ZaZdztJPm8xml+hcvhNB1EH88qQiOt/j+a++NtlQKoDzkEoPFU71vgF0JJ4R
ud3B7zSFe3nKsYR5c/giDcR+dFHwAovz4i/L4xzm9/QeEZOAi79yPv2SdaRYNf+y
0VHhuwdrS35t28dh6J1eRg==
`protect END_PROTECTED
