`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fWo3Dcbsj4q2/p9S6zS7I5ZjkYSM8d53G6UyHFQVtIEKKrJ+K5VADXpFxUt3Cwg3
BsX5KLPCYRa0K2spTsxuiwx2ocrj8+XB+JHfGLRJ+aG7G1FzW/29FFs2fwOS8+ZL
l3AR78sQuySRsDL5hpgrqf9RUcHwMHlWkbmmLE8Kiz+yep2dBrrAhKmEyyCsghA2
t5T+p8KvpVQ12wsQ+d92JVYYL5XbJgpUBx9PIMDYJm7SvV8BbyhavFs4eTeY3nyu
Lka03QgZGkUFzQOf42m/ssyavpYRiCj7ANzJjw7n3rqtHBZFdmfM5a61itg2WDpG
vj6h/N6VzbrRvxMbbPQ42hzCDFz2YPE1CrN5BxZIxoluiid3/oPqwubB2R5NrWvQ
l1SL8ohJqA4A0FIIospvjIDk+giHz8wH1NxNQanmMqJpWyuK0GxncnSmmLOhX3oi
IudYtXTQ3Nd55O1wDC0YbiOmNczCNP/9kWhTk12WLHIG124Orb91O/Hs31Qh375G
xfgifKg6+B7eZ22683HhIvu1ja3yRVb+XPaJFnLta+3d7OjCLkff9HzjeKGeBK5X
8MfMl+SZEJerSmjGfUTI7A==
`protect END_PROTECTED
