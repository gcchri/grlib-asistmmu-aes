`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4nboAOoSGrY4GKiQsu8FP2C8BZbtPGRRksl+ub6EU8ztsgO3tWewSyW/kWrTD8fX
bmNG6nfrrtetk0RFlwNa3wbbwWN7RIJQQ8ozNKXBUKbCoBWy2H70/6CDEo57WqYW
aLlynzruc02DXA/XeNUsau6bVRU/QvB5UmiFqjBebTTcNwtRlEJ/XrvBSdiLiUV9
ypki49WVn4b4JVKC4QgngNEFb1kPVGKfP2xwM6cPyhnE3G+atBCmeaZUtzcsIxvs
8RKl10fR4TXteX7t/FE5WwtRLvAr5sjr266vBiVSAqi3eV6boOt3aVtUPFtqQXyt
ccqoGMm1nOLAkzxEhG9vM49bWD47/gJdxbPU4OEuYmiHMqAP6DPWI0HVTHV7m0RT
e7+VXAyeDMYPIDEXzB32WIUnxrjrqpjCCUd1890u8icr4VHVRx8tqpuMo07jlCBk
JXtqnTZhc/Lwl8YeD/RuWXbvijtBMzXZTAYX+wkPnH4dSFayd/Opyp+LTJDNg3wY
A4EkH8KVC3KhqN3erIKAAAP0YIoSjKpWsE/2fntDg6lXOr3DCzccNi0lF6Fm2c+H
mw/u+4wzqdItGRcbjigZzyvo7/HCV/OgMygUo7PEQbb/riUGYmUjbf+YfDkiFOWb
zUExkgGYSBzRiqQoTQJE/aE6J+TVne8vX2psD89qioZDwP2v/SuUP4FPiOPf4r4n
30tswhbAfOEsZCPAZ6hlhi/UmV0HYx2xOxBj77dtUTGAuOuzOUCLFNguLjBk9+GB
F/SXexHHBgGS9sMCVD0xZBI3TNjoCfoAj6s+eQoxLB4EnOXUKuORHJjaCm6EleJy
HDsqqRyKsnr7NMwoGkL7ApimZSdjtDzVcAHoDwb0jl61C8EDRSc+V1+PzW8hEy0E
/yWpxOUyYeSarkmZ0hvCbb0m5F76VrvxxRh1Et1MqZ336l/9ypkUbjsT/WxCkfVr
lGw/lxeB+6f8G0IJJu7h1EysJqFZm7bgQvfJ4dEMUOJVNZFmNT6hVIiwmUrbaAw7
gwzeavunceYexDNVpSA/Xq0SSDFXQ/sljiqmBmoVf+nfNBQUw1Oyhy3WABrMW1ju
zdXYVzsJCVzRP2eoEe4Z//6/TP5SNqIIMQpjSrrs2GCD8+b+GFafpa4frDtSrqti
aBlQB645Ed0y1zjAKZVtpG9dNrBp6j7bpxFHiwye/Cee3psSVjvT5IZMYjZD8hSf
KIvUR4m4wT57eiOuHNf7WyeLQeEDD4QXTOpWLiWLZd3XasXujt/uI6dbcB6x5uhr
37Xh2dSaVP5Cbgqeu3i8RgilVuaV5I/F8ow/5Q9iC7XmKM4wAvHXhYdjoQLaijO4
XRDTktnd8Wm+EDuWVRFjusYf18DTNR1WULK8fv/N+tQ3WkMvjRlYPhdnmoaBUKtB
pTnXuCqp62wIdU1ngKm82OHqDOSdhJTDrdV2eJy8g38eKtSFdAm9NYmgoE08pjW/
BgD7NQ7XGBtOFcw6BKqpXGjLZGIBubs4NEEuWn2JsrZz4MaC8I8eExQw7JFQ7Pol
iuoQ+MwnnW8xkZ5q8sYOVyH/VYTaJpMUD5DyviK44EZFERa1NRFied9uaV+GZYTC
6uvN7vJIQh7lGtkfMbg9YHeiQb82ugHOAIHiqtP3iQnt6t+115WnCI3Cj0sOlNy6
c+Jew09GMmA6ixMXlBjtbGX792rKPpMlvGI6/qZevp2e35CZymQ5m8GxRHCXS3Zf
Gm8kw2iB7lWaiu4umyPhRXSLcSOVbqXnFknUwMbwKIOjVdikR4Nn7rIffqm7r0j3
b5v59xY5GtKQ/WK9KEUl95F7JYC/t4iveZtz3yCu8TbXgo0KVT760jrPxdL68qw9
4Sx0WNpWtyNPX+9nLJRM0NKErf+o9EyAOFVxqCz4AJtWNSWY7a7g+4MolhzzaTqB
h0nnYG+ziG1pjy48Qw30Mmm+ykwtCsLqfa+De7tJKTJrS6g3dSweD+SO32XeYQWJ
TdPJsTquumQRzx9e+bTRfmc+PKYzm5Va0tmRQ2O9hudjeIZjJuTZrDWXNVZSKIdQ
3OegqK5IjPupXi4OAmjU3pSg2hhpREXl7cMiymth+inf+rzPvxZLUq0Ky8hh0e2n
jh0RtmQzMU4ewYHgjDtbZJFCykTD9aBFx4YzHmdC638AhWXH4budYQEpjS5etBaX
qk8FoNAY/CtEM5odO2qMX5d3Q6a4/YW7qLIeUYpck+qHSOzBenNOy5b0Pd7kAlSK
vJYKlGrbE2H0lTdC1400x42U6xbg4t2B/b0L3aaFByscQcwtPNGEdj8UFpieFPJs
mRK4SJy6Xf8gZfEwNmwydrYCdMUCuHkihZryUz48dTLn14V04vZrju1VWGifw1AK
HzY+21otvPmnNSkalTutD4FReJBZ5YxGf4WX/TV3w9ybV5spYTiBOmpE6TqVZhqj
gFI82tpaRYATkW29JA81ndpiCtpqiDW9Eh1KYu2WW2QLjlaMhl77NOy9AhpXJTG7
QZy8XJZhW0U+ElC/NHBRt+oOmPIzIl76OVfTN7GiVea9sOArOPEkk64eIc1BrUCV
lfWz/ohlBBvbSA7FcRckWUI11jPzlnvCi+oaL/gFS/Y3Auoad00CMp8Bju/7hvMh
rSZQ3uFQfdrhumQgiiNYuZujzwKTQkvgfrbxwLIJsBse/vbOA/94kmWAFCF9+aav
TAXawKkj2oUAd5qfGHaDx/7INvoiBmSEHXm+ItZy3l9jBtJP2h5gvdjCnQ1vSSX5
JINc1x7haJP0o6zPZPqj5tJMPSVjONyDM6bV/Xxi3EWPiUdAKb687ALTydaYYEku
tMLCF+WVwzR7hJgDZEGjH4Da8iwDW3tbucapAXpolfta+B0yFnNBqe6CzqJ+F+L5
guf4QcDlNhQQWU2bIWCaKXxgyxgfiRIbd8OWEi5igBdDJutW+/pU5kubNDA7caxT
96jLhOdlM4wFRErai3mxAaPNUFagbXVPdiqn10taqtBUExLFcg+mFkSZzn7J0eve
VwRaccwyGyL2iPVSeSBoH7wTPzRlJJH/BXD0eAohB7jZ/LwuMYH/EghLHeIahEqd
eOKeLFw17LrFM5yHhyQznA0CHIIHADpjDgViKXFvl0j4UZsSfHzHtuKNHH1dtO3w
CxW9uyqeEpsNqMBdh/aBm/eNQx66MgoiALHo3agkF0+45tSXMKvoeVWiSsER4vnI
WZWm1hoWiszMclwGrwC7Mbglfb5oIaYeZ+gstqywEMafqF607V8hnyqGQil1vQgH
uhCAPzM5MBkIRzyXkuihiONoo/7Vvg7YnTxP028Yc451pHgYKayKi7ULZbT+YN6S
HwMxJXcxv5tHIs52L+rhF1tqI4REPlEXXOkG0huuaaUHGg4VLuJiOj51M1E9pNkb
q15xzDoLRG/DZDQ2oAmDAAtBC+/IFt+UOSBZZKJowIO8WBN33LufiuwHjdFaERvK
qRS75v9RwiAopIdGl5LOa+CtJc6sn38Vg5LElRjV9TstdftiiHMAZQzILSSFvDaa
ofvnKWNyP/GQu8u+69HTo5ZlJg+hab3aBjf6Aj0PEo2hrC4yar7J03HsVZNyub75
Xro1r2z0vAK3tCxrXBkVsDTjRRCb+bxRQF55qujwO0hd8rn5P5Cdv6cVS4vKMQK/
Q+dYjk+zEFMdq6s9sS6G1qEA4cnYxIOlI/axQYaKtqYt2LrG3x1+ZPa+xDNgMvka
nuWIUW2xSv+X8/ZROwhZJthE2gYecGylRIi3/Lp0h/XCI1wOl5nzCFZWTN0gIdTY
XI4qih3BBD3D+Lx6dyJ9rb1H0aWohqOFfz+K4JlWDVYC0juDejtj8kS5AgDQBqep
JjtXNV3obKuErpa4g2j9hfGAF9A33uy74zwJyyJsDSWNXKQZ2XfOLljFZayxAKy9
6EFQv+ZQgFF4uXrRS4rluNRb1BO2hoURj7ERnsxK6CoSri4UtyEZVwtxo7eECLrj
yHPWBKB34oMjEe0qcRLxX3ANELZ6PFxBSRiVa+PhxhdUiJvcaZAKX08c9xKiMz9w
ZWGP9qgMA5PO+1cJAl4rFcBIwfm32sURLRK4ORa34vNJ5ad2SKkPzvhFxi4Cqscg
3xuwVMQ0/zFtyZKjZlAb5XYDlTlMmG4ZYQYULaFnJrqu0qHxfopHJCrZXEHbz0bK
4tKpBEZIzyi4oBdSPjZ+iWhMXOTek6zPJqYZMBtXY79s0tJyVZ1aJkhGsL+rOvSI
JBVvay1k/1oEUiLkwChgQohTbzIv2DD/H/WZFhRK2dJ7ZFO9hp9Fm6XuRut7Q7PD
t1E7hnnwooZFGY/SB0N21lbNU6OqEIMFVne44DJwvWZAq4n0Ogwj6b6JxwZY50D2
sOH5eWyDCZ9fehwTSATFXr+Kfy0l4laEh2HpwK+xq1etroxzvxu8mBC2D2zSXsLZ
TL8DovRqzfDA9EdVgpZyVdJmQDKNhuxAx0peQhMzl6s4yrgwMHDWR0V1HOc1TFUA
ZkSiRH0HOluSVwyNyEYE3tR4fWPG+wEc4T4OkYnJkr8wyX+8ImgkLnBMGvO4fWqK
7pJTlCAc02qLTiTaBc7SnOR9oDmC9YA3wGyPv3OuDIru1/B7QMDVyfTbfFajga14
UihUJwNoijTzE6NwMooLPrlalulN3nTWiKygEr+cvUv/ofF5mqCXrHTUcjhy0fx1
lwqTfKWT1mTnd8Ueggs/o3S/EZ7NPBkUO8lFO+HKVR1/m0u/OSvdxzBg0RC/JDc1
j+Q8lRht/3/Duu7AHCAM5LEQHYYWhgmgL9fAmn1Xv7f7fdI0mJO6w4lyBN00Psgv
2k0gGgtEX6zbd136s/3BkjBpNkGkYpKkFFcK1bKKXzMacgsYbv/0u639nKAGVyIe
9XIKD+tSbN/ej5jTivPMQzoQfSef5moQKN0QxAml65Tslz4oHH6eclNjheV8YKnA
jPE54PyNR+WVUsng4W+lQMLTJteAqgrqcgnXLuzSiJGyqWGRZ/UbMex78hlalfLj
VeWg2WFM08/Y7cWifMRkKv8795TObphkAUlA9TLk9XZsFlLMd8aUldpVokwgOfPv
kBHDwyLNlc14t888N157AIUVa1W35FWgmWTvTlugSsTIkWXguzGdbF5BpivPT5+m
2koE805+Rcvrc1NdB9AjgShd+8jRtrfknOodPuAxiRkg8ttP39z9sF+JU+hsgl2C
k1/FqgPNespLWWRkUgtar7rccNnsF02CER9W//XXBd9Mov2VCRhPqZV9Kr63Thvq
HbTnBuYHuwMumnD65oKQbh/KIy5/1SQweH+r0UwWVbgLH5qOruHxdZEyUJmmtJpi
u81j2OaH44aLu/VOOawneC7IqrNQm/3tCCo0ZL7XFP8an6X07SUoyXABrYVuyV2Q
zGcxnDp7CjFy+b6flJThGwOWyc0Nl9RUgzuxu1Fn9QWK2U8GWck4v5z6+JcgvL5x
0c7ZE1n1gXMYFpLrnFwwbT0F8onJ5owPWH3stKHPk8TwzJ6cTVXexxcJ7huhLNAx
V++ng0EDyO9hLm1wLZTTMG71oqlrr8Z7w74c43cdZOOatWWp3rfQO7mzcJxyIBv/
ITv9pZ8j6jGV3/3qZhqkSElWKMAMvSveln9vtreqafAcqTQW76d6ZlusmUwh5rNv
hTESJfQePOWuf6ufgpdWPPxIE/duhkUCZejcpDnFY2+zsY5lQtz9OZlKbNIEp75I
ab/mElwRUlOTcOoL9sfFtVi9ZGCKzH93kiYq1aPs2lKEWdCSuEA294dFKmjyrELX
GEKDqOtDE9D9f3glCWSzsBg+3ef9rB6dtLDhtgKHACOW1dZkMokgpXM4EHYSJMu6
vVVoqAc3qixUDyf4PyeSCSyYjzgQlbfqRFITHaKjzPo43ECIpxJfXoDm23/CE5ne
UF8HE/vD1kPtjOcBnl1qvh3NRzQVFy6Z2y+gzxuKgiP1fPr+NpDcnV7o5KbA3c/R
tlZ+CpTxwleO5X+ZC6k/EkLR82Q2BAaS9wDbnTfk7ofgIQitoaBEIjl5UqXnDYLz
6d6uWu/rKe4Q0hXh4IPaWQBc6z8Dbu1W0Zd2rY9MDVZD80ctBk1nEDRlj1ozoY6V
abFffWiPhTnDCqHUd3FySEOele7hx/XyMBV5301mL3H1nPOYYbSMcdOBZcTlqb8m
TvretRTbBohB3ETJ4xbfgWuIa20TPr5Z7kZQuyXI7gZ1SN3deAZR2B4V8NTBwi8q
nzaF5UnNsm1FYqP1qxM2c3QeAnFGVAJr7iU1qW7N93GufH2cA3b0pODRDHNa/0Lh
2ZJRiyygzWzZXStZgklimYhBEhnt0uW5LnnuquxRILIDCn9RHNvR0hH1InMDi9IH
rwUUIU/WfZH4aB2U62aHSYXW3A90f8494HV+BGmPIBwpNPAUo1UwJpj6gXSan5fj
Bbj4m+VdnEYi/bhPopQJexGpVRfnjB3thZoR138sfEwpiwnJwZ1ahIjFH3C+wYV8
FKwzzyFp0GFEFK/ILnU50zor0G2bc/AeNfPkZl0gKd1J1T6oxEdmjMEnPuncCZoh
wLWU9AfkenB2J6xeiSZq5ZJ2/mXHcyi+TEs16yedwACPC6yOg6XbIefxJU90i2uJ
psowx+dbcqCGRX+arteJI99vDSFBWxCOF23E2L+QHiC9OkNCSTzX2pBLavv4T5X0
TyuEpUF4NvPwAGTtm9G/UdLC4dC+DAihqtogkg+9jHX22pLDkARIRChCul0NZz7a
ULmQMrjRxM2aLdb4oYOtauE0Q+AOPXyDGJNNgAbPOJHoehISyetK0oHTkWyUv2uq
UaBSz4R+KovXwI06O0rePU8u016+AihSRPsyMSyVfZtibc8mZDUN8ey4LIO3oQ0I
Suox8vFXOHjwifH/FkuZJd8nOOAaR4t9uVHx8qj90KRiRXryYmHDWyOaDLpxm1Eh
FL/9VpiTDJjzucZcWPD+1TzVVBZG8iw3sgv5UtpQVwD4yDQcWADz0egj9asrWFfq
MIc88JuEOnyuda7z8DA4Doh6pLwEIFOQ/PK6PCuRKPSmIdXzyQnrl3TGwRXtQPOo
kDn+9UkQxianwbNhh+FZktYZhu2Dic2EgQiRPF3PUe+rNVRCR6sYf0Q8av03309R
jCj0bzGcS68x2k7lKR/dEwsiJr0AZ2i3mM1CXp/Ou9cHkJcwq0OcU8TVyz6RBG6Z
HOOIJKvEr4g9bCVCHkOAP/ak2XJOJiezhlRu4Gh0ungy1iw6walAaAbR2pNXiaWV
61OdQg0f4SqRM9OZC5CnchrYyPy2j91xb4Idyl9bJJCdBCPjez1h3QtZDgbqkC0S
+wLdsLd5Z6tJpq2LzxMhgeiqTR/gPqRRlhJLfuywgKJ+1Bh81OCAIuiEDZCxpL7a
UVMfpv0Es53wqd9szF/QqjvqysxpMZ8qMdVh63ybcL1944dN7CQCPaAba86OqP9j
kQPczfJSLmuM6uB7+6L/Wk18ksK/TGYFbFQo5T8VkhXGEBGKjL5LRkz9ZUXrea2M
6RmFtiI+YcEquYrdUmrN8hXGdtayPnhEViFcFPeC2MoRig4CBBf4EFSMVuMftuuV
STrMWlbkbgIF+uaECX7zflSq06b0a8/Wcge7YrGDVspx4K2XOCNxLrFXKpgB72QJ
lho2ehMpFjMQScmsAPLqegCyJZdjCNlMHRQzKua/OHmob77zAq7tECWAiSs1jwAv
DkBkLrGGl3yUL02Q6u0Pj+QMMTxAu1rdtRer61jonz7D8uegxZR2Wbwpnp04uz3I
Vms/yY8WojPPeCRzVXhYtckysf5eAyHMLLqyp+wUkp6yp4ETcriitqeTBhS6q92p
6mPpYA/5TIthgfInzdD1TEt5Kb1LdvidePPr6rPzaCcN86TXmZvWYPi68crQzH7a
HPDQTMhPB5kR8im2mSZqXU7NwPkruwiTlpYbcWO2WptM+OoBw/TqKqcZN7Nj2xdj
ZbAFePVpDovjB6F23Le8O7dfF5kuPzwEysIWn1LULsaJeCk4Y+ccMgh8DKV8PifS
Tn7hgYVswvbIeDJSDs2feixctOnHtSRliDnuHuBV2Ghq09ZjOszcIFxiPoIfS2NA
m96wHzqJs4t843VfAQNoykFaHOaMX9itS/vDVZvVmxAFPU/oDiGvfpPPMMaNeiSV
58BCFvSzEDRenfoxZybWkMiMza93oYTtFbCer/z0yWAuTJW64CkfqHQeyJhXmVYL
eoXcSUON8sxpjMTqkrkfazd+ecaAcurNAfdgYJH4kLuiY4U0Iu+ZGn8c4jsKvnyz
YCa7aQEps026iT5Mu7TwMLdcIpD3xUC6AflSsBvobHlfllfwlv8FReK4hLGfixqK
GsUpxymz9ec+WVLlLcptqfyZNRNVP443q23BX+STL0hIVndR5b7QgeextYosqr9y
vPyv5l1+9EmrA1KtfoyCa7bIKYsnn9lU9pDXQwedYkEYEAtrm+8zaZaja7st65FZ
wfK31aH7VE9P5IoSiQkPmQ6tm7cFJ5wO5yI9jwJfOsoaGDTuhsQVs+EmSxDw6P85
Cg1lh4L3tH0Mm42PWRQCGnlKNcviJ14YDbbVGqkKxib9LCvbwHToW96QJ49tZPad
NkDNfbJQxB6erXl5MjpxFtjuj+9Y8wCv8kI2tFyoq1gm2Q20cvWv3tHcIUpKJ5LI
Q6CDalHpq5Ayki4igaQ3f7zV0rThNM6jfD8ujIR2e1Q3O/3o5CNSyEj3r9ht6Pq+
nwrldw9RbLAS/8V2xqKhipeCNNiL4305Qs9HCAGco/0bDpvwBHwfkvbq+W+pT7l/
qyHFLCNGt9Zlmys82RxZ+Td2xysoVWgw1H9s40CcqlrGAr7hUMxEib6yVJ9oPUY6
2+iXNdaWHT3Hew/+zDCUdbouX8b8lrvKvbu/nfWPI/6DtFOrazupppvtm3stczLg
5yMnvpqpQRv6prtxCimS+9zwqMx15iXOffvh+vhrPPseZucI5Q+Rg6fJjLAEyQ2T
69lJxDjImCa78kQcjmWcsjyxn0ugXAdwHZ3XzjG6i+59BM7AkNm/x9dAzS5meW0K
DGJzoCS99FIPKAHclXtJVII9kn4jvjgk2qXfHKmcI7vX7Ro4/ZTY1gKUtcDuiEf6
E5F7F9AlV3mkPUpbwjFX4mk9qdDcOk3lS3mbxz1yzdWij4J+X21M+A557NzrmfD1
40xGT2PFu9kMpfc/5nzvOVq3ztsngE3vdiWPnpZOZKyLkjR8tVRNCC1ME5Bi5deA
ny2549CSSmMz/hFX3zbFXFu1MhXvlLRbx+wNLt9aBKRUgj1wIgMnbMW5UIqQUsci
nANzDS8QO0zW2V/OGFtMvv3tUlf9gjnq4cu2Iqu8+GwDxHhd2LhrSgUGPQcVpYd3
4J+/msk2XQvFSuQsIuk3fn2DoLhZlTqN/T00B5+caNAMM2ZdYNBlaZVeb72gNYBN
gdOrxaojij6iH/klUy4DC95NieKcD5fMVaj/cuJ/KpBuWxnPtG6l5p2LTWOhPlET
KPNFUu7JsR+k/vlAFNSWVQmN/1+JJCHXH5T4kms7nmuE+h2a8s8xdzY0LwjjRCig
joIKoplYV+a67ZE5iRCpDDJ9OpZwKwp557NPnO/tQ1Fj6qaYjKA+B7XfbNUFiYSh
dfqebCFZf5mex2Tx4gzzd8rsBSOoYpfLz1BwcVMT4OyafyuXdvFnLDr3anfCLHr6
MlTrvEVaX4T/YgMNFBpr0IEuq90mKJaV8U+kckC5giah37RQuFuMkjhiiJL3/GMj
pUpjJ6Q807NYi66oQLIPyb7MZUir6NvxRh6YtPn6PUXSUZoWPABKEvyYiPAeioei
WrkwWBhNjA4nVwBRtgZOXqrVqsW3Mznc997y+IgSsSlpzkvTMGmeHAf8xZlNs1P4
XOXZXuRI4Kxaip6AkecH1epco3YF5oC7IMDm4+LuhKUEXaFEmlu0OtNaS3/1L+RA
JPKQGLckmwmxwu6lWUYGMP8eW/bz70gkAJaKrZjLE4lQQar4Gaf0iMvFNvCAQ2Cj
amm3F64++CTSwlCxWlJBfvuMM/VIiBibaarSvFp7HUVRSNdf/0cyOB39iiJJQoCJ
utBX5KgW73RJetFjlVNto0aS7VRUM4lFniOCJILquI4AXoTiRSF9rGgP5zKp18w9
JLihkRhasefNdS1nExpmrj/GqE95zYef95AOvOMXKKJxNGL1HWyYSWYzLM3V8o44
TGKHqFF59AxN8MfODcQgOTQkMKUL0mZ+AXqPLZoMS/94LY7G3Ck1PBB5v94nOYZY
TCIr95lSPgXwVSZkipw+oP6QQbfZyFTBDLGMh++AXeOpnBwqzbMjkSoPheA2h0dW
fOllTwcgs+tf0R1gyTn1VqEvUfPJOSXWyhSvywXo6jwpD1V9U1/laPPe8EF+cfgy
d0R5SnTpyxZWEk8gyFOszu7C1ehDVf9cFTMxu9XkMTrvcGFrrGQgin2YjeLzTjxF
NtoTnNwHYrffIlbCUz+BJ8jRc7PB2qdG7L88Z027HT6hFahE7TAVR4HoKi7tMbZM
C+5mDZ79JikD9Iv09IenWvxywrxzrpomT3Y/2phsVzm8Y9+IFqg4BGS5bZ/Ca2xo
yswhBe4YyBXg5jXwXK579WwI026Qr3G/22FY8PlYPXwesJdMHp4A9W8XCFkZB0Kb
Hl6fMrVvaj54UT7D3YQRAF6/uLBtbJytk3pIgQa1YzOg8TNuZOcBUMWT9eNmxci9
J6QRhjBbI97m0R4DZlfcKk1C4G/OffLYgHNi7Fz+J0mYR+3kzrrUOzm3tYf0i4CK
FJcQZVAIkJtXLUuMgAKU+DruoO9sCO64CwZGt2RxQ4CEQTjnqz3XucPWfjE33uSi
M9Dqbzd5M9nx6WJelNvTw2VfnLHDZsfiPVkEON8U0GgCm6DIKWs0KauZ/QzmdeML
/IBZUe0J7ptHTjud7P/pZM5DFJI0w8my7tcwG/2VwfleXiEwgraWaLGcE6aR+Gk7
w1w5+cbKEFElmMoWw69KmVun7Q88bx1WAjeotHojS1LU+mhxzj2WWXDXpKcS4Z05
B8+MWFEAorVjvz9PZpMWraAExuF9TSeCJuw9F6bb1q0MRVBcdYLoYceMWumOvi2V
vnjJt8ZJW8d4q5OZ77nIRW/hO5g4GGYSf6OaPDB8AsbPbYYWqS2XAoleEA3CynhO
hmpUUGkskbAZvcBaJo0rs8VYNfd7sR6AGTKvZJtfJRoenVuBk3EDITPRhaA1+aMn
3y9ZwMSj61I2wKAPyZUwK0dsT6qzT5SgTDoXbd0tm6nQcpkiNQiYLC6dyZPCzmPH
0no/0D9QXZcNcR53eejGAHrf8gqutH/lndUxiU9Il96AjbABGoPXsk7btGE3j2Gn
zkpTXTdflliUKoswsIK7r6Y2jdYk/BjTLJjqSCZH3m8MrTEu79u2ovnTNf1SCO4B
CjlqW8TYT1WKAGxfsyGwCHQ+ySRAdftgfh/gzVk6yzhzL7elVRwV+vglIowqGL/+
LGKjF+j+BAsBsmXTiQMVbJFI9rNyQzXyVDCzs4mrVTAAMAqQhSTG9/qU+74euePZ
oXKoWOE6GrTteWRT/pTHAxgU0CtUgt7yN1cagQZ4zRAI7sxGO1ePbJBNPkJQfR9I
3Q6mnARMZgenKONIB/RhnjAZN7FJ67CrUSr9k5+qnUdu5nVoShKGUJE6ri3Pzds2
nhT2uZmE1MmNwhkmI4qaOJnSFhAK00DAOAQuYQXtwPnZgrU74UMvHLvGxr6o2baC
3oQcJtmVJoY1evaqkewVe4o2cCiMeqOSbI2JP9nLKkilpOyVjw02hIupE7Vlr5Bi
fV4lJ29cmMMRjuZ333iZTpOUGAcQ7Fa6KkqvmUwYH6EDlesFcB59rzJ1yAVGlwh1
dtRiFh8rl7CyGn0oMJsogtL/KNWviJWcVYIWzAE9xlUR83yl4cjitnaayzDQJFDb
uWO9c+wmmQXen667T7GjXCno07mxMA65B8uTO8SQCUy+5im7TyIvxmUZ+Y05OXI4
mvlDixS9hxPZrGgn9CyNgniVlflIBccp0RhFQw22cm29oLwQHwETsI0gOLezWQVi
uFCPL6095BWLA85DeaNXYED31MfeMBH2aCsjcyZ3TLoBNwPLRBBMLTtAwS+ycBmJ
OvayeatqC5qv5A2BSyJEvcRwTbYB2+AS6bTNZNIOv0vRGdRxdQym4wqfl98s+O19
LughOjOYORjhnG0s9Ai4gwXigU3BPguQS8cC5f5cMMsLWO7yoKJxTtECmBGm2pqW
z6JUBOGpOd7Sgi7KkeB1UDpgUAY9zGcfKQdRbosotE679ZY9iMGRK0sYSsI3zF5k
v44/Vd7ta44z9Rf/3uFRzoAW9+G/n1ATN7oEEh9MZFOV4+AflIwsaVC7rk2KqNlE
BSzDhvuQbLrC9KJYkoCr1sYsHbXoWFpq9MWJP9Cw9kgkngSNzx6cfXYdczElfYTE
/Cj4KYCwcU11y6x/Rww41Fmktgo3oKLJMI5yiX9gXbQbh0B/cEKv9sLUEAsqixBy
Uy31kJo/4WLFEqw+Hplhh0LJXuNVBu06ScezQMhqRMsa/4jnqhOBRraNYEVJtjns
qVxBV0jQ/WLU1OGQQot/ppC15KtQ4ZW0WDenmMr/iiLlIGCKt2Rl7dyhTgxJ7RxJ
ccTzLRYaMUHTi9YdyNq6Mss1rq/KjhFsdjibZAp0IGb4bU67KxK8ABdV5NTfjWn7
9tGEUHp8wFpdUtn3pJAuuqKEGr+dzXtqq0oFQpeldOzUcLEO+ekOqs0fpFTwJo3C
iVOczQPI9ZFl4aQdOAk6xnm5QC8iNIsBf3RaXwIXrHHaXzECtTm4CBgp1fo2IHr4
AzgwPDz7kyXldm+PKaJ/d2bPSsqbVNRV/KReIzOJXF6CSqN0/f5svUsNnVxhvBLz
B6MMtbeDjmvKjvD+T6mCYkggC2NV8vcGU0TJ7P+b5WSsQdXBkxV5ZcGan5bXxyrF
yEvSioGKmp4DUBlx3j1CV17hfKwBuiZdReVP/s/64LuyI2koBOWNZr69nOCLHmg2
qSEIpDHTYwk3j1m6HdNw9U/oqevPlLvZxhlgNf/0cOzTmTxdArZhl0VPxuJoG283
/Q/vcFUxQWUIVQXUe+oHRpYz2vL+gmy6IUSL74lgBWPhsqviv7eTgw44GqtnUBxk
0VSnE0ucK/LMkC6EcDv43Xvgti3EwhR8r8jSpPqJEb3TmHWUKlB+pEFTJ0sAjsGN
nicrJIyAQ5/O4AJ9vgyJcs+vnihMjDQwqv9Zh4PonQTn5Q3HkkGGLyJWGtKj6djy
9BeBuyj62sCOB3jzuR7wyq3dQVRf63TEhOfmiWNkIiL5pVbTjQyXrPyiXLjWoFE0
R30AoPyy0TmL0n8YynQdbGVravv3M1E1ykGAiOhfrhGCERwEkInLHmask+rEUK7+
W9ZHgTGnfjdBbo2AmlDgzhe7DrZT4S3/9wHNYKYCgioX+AESejBoFdCq0C56Jx2G
rkHcbBn9CKdKRPbylKjyMb8r8SqPsPsxjiqRzc7dwTuOk3erYXh1WihV/dLW5Sf0
2NUuuZffOv4qan5juzlaGQRmLzM5aKINkA+K2HJLXzXpqlVg806AGCqrdRGr0Gxj
8hZmx1U/I4TPJnkH00VQZ3nLQhL8q55+Yj23KYTGjexyzojCKefSieoR4+Fcajxy
gGfWQz/mR8E1trpZ03n55JV/tQ1vEzVqAr+J8iPrkRRGt8tiOMWHEbe8cQUrbAqK
2rZCsyv1qsrel/0rICxxDqOFkmAsqPvJkaMEm9EsbQ6JAL4H7ndxJfUQsjPgFlEc
F744mUwLmQ2Sqv3DgriWNtvjyry6iOJRXZY1l//4iFwMecxPGzxQ63O80E9aYn1M
DrZX76pg6cdsPpOqtsutbmEeITkNKLJgNG8Fw5ecCDaL24Pdm5B1jv6HxM7Jfejt
c3Iu3k+YJ+B7KsogvjSsTOLYPe6lWle0dEULPTM1dL7J27fxyoa7a5MKFruNS3FB
8Lm5kE+OW6fVGI+jeboZP8in58LImzZHiftm+tTx9hsXa/iy8PzgwkhAAXWBxwSI
u4Xhmrc6+xgfFXdieF3pzsAMdpEjVtNxW5l/WpqQuekYgocdcMt0fp7Dx5/WUpZS
eYww1JleczLIK4xQev1TLBtAwEvr0yPksR0oEU4HoihjVYfqRebvxJmGJDIkaLq1
yforjW7VrMNp7xep5tev1wEmik246WdCposkZ9Seo12vT/6f9Tb35E6XL4QJs2z6
CFjSNUAynkEYTVD+1b5/KLYiV34BSYQjBjAxKx9Wk1gNRqJA7Jpe3bB46N+Q9ssP
fl1xzrpKjIhPCxnwanf4CgnaXT7ovugAgyHLqu7YF0UnrH/srElTJbER2h+ymDmL
2nliGrBhMcnRoIalYsGX7kKmtby2b1fv4eh5vk4oqkPhZeFp5BTNd4azWUd1UwEy
k/Emgii5xc6DYkXdS4AC/et621KqEaLwLt9x6f/cS+M1Mo4T7S54WFIvll1RO/fE
13r7HWAdgm0pj+aGoB3zWuaLR8vBY6xwT5Q1qvxlLE8+0fs5O1fIq5E9Gp1U3gex
JWMW+I1gYsV4/5jj526g8lPGHlZr9BlLFcxyhmKoyISBffQ+r53Cnt5PQmL4lhyq
LUtRFTQ0DsflAfEedRTR/Bx7E5zlcSDz5bxts31wztJkURzHlV/152afe7z3l0hl
/NnLVsf2NaRi9Nkz0P3bFUEkxTZaYXPtou6hcpm/jtIl1W25D7fLGqg7YaecFyl3
CbB7FoTsKTwzLYbAjLbkoxAFpgPmD2AxCYMkX+mecsim4k2CB87ET1FgWkZ0vGFd
DD9fBMQkyavegApQ6BC32Vp2LDV5SqjMVvvneGSjS5AKkBVP12iJ0I4uB9z/Z3To
peXpeXcXt1Mc8jbxAYCsUfvRW/XqjdXwQmrgvKSxX/bLZ5flwJpZ1BFFSj9c4K66
WNeCKXKTSYBJa1E9a75ftKjI2fqhMMlMwNYeXsBq1Bv4reUapVgVP4vto4TxpsYG
rvQLS8hWBtmzXlTjHp8dARVnC2D12KI/ZFEDxtYBQ4SImntcUHdyR0IIvYNEndZX
aqztaHilPG/RXnoEZrgkcuio/aQ5qgVEQnRP3nL78YpJrGtNnwSykck5uJ/1cxM5
knvFn66e8EhdQ2LoPlHe29jM0nSyhOaHjtnLb4bbv5kXx5elJ8p719F1wUiwbRnu
ZeBLIwgCD+/8405nz7h2UjJWSZjZOLWBzcP5ZFfFZvKgM9N6RY9LelKaBoimy6hR
tgT+fR/JTpKoaMbbM7UgaRXVWJuTKSj2p4oFhWkXbcVYp1IvLal+GIrfhMLX1uCH
Srh0oQ3yyaawPvT5baF1E8ycx9gDPAJHevjdenIw81gybjCFCsqGT4TWSo60ptHQ
+gGVXc8TtYgTvy606J+r/xin/GXqOPIt1Ye4ycq6TII5w2kzEnuuNuHrn8xzUPBV
Tp5m2EXRAY0rL1R/bkR1hMfZk76K4TuDvdJVTD/3s5ynbRKTi2s3W9c9oufpO+pk
Xm70EhMaTMEDgy3Zs9y647+RvZuyIS/WQPHBU++rXMKcT+hAMwDMJ90KX4/vBrk3
YZ03fAM9lUivI6B7bhG73AQr6YTkwN90FoL4POylU7BQKVr6dKjSdo8/jF7iqeN8
j8DQhFLdqhgzJ5BsYeNbHUwWoNpaZlINMEkkNztcXRfLsA7yfATOTppFaMJb9nAT
fvzouQ1YrxV5qc3M487lCH2Vjt4Gy5e4WfRSKwcm+Gh4i61sVaGUk4EuQ8WNfpBA
o7yvWF338VKCYSm4bMMb5cwIKFGkwLOFHVzLWn5MGH7WqBFGGt/uAQu6oEOrO9E7
tgc8kKV/wOd6ZkaiJv7DumIU/nL8ziHnvvxQV8rKErywhITFHNaZTFD+FcRw3RjY
4vSw26xa/H9vDoQTaB3DlOJvcI8Q9fwSjc9B7+XvRTvlzNwxFRQxWi7tVU3qmX8d
Ad4eL5GI+TFtGFoEkY2YSmPB84re8TJiwLxd+YRixKXy1GAVrCF6KeGtZCBJgkDq
5r56ReOUiavSCOGFlx8keRwPg4YjG492Ev4wTpfAkhpxD69JuXLTKjnLNDVGW3Ib
z7z5I8wa5/42wNyHWJ3SHNMnZ5SXEzVgZZkZ/OVPHOeALgU2W6llJhm9VutnPZBA
UzBs97gVicUhGD3hRy321SwGaguu6W1v2TB9sSNMKPX781OJiiuxyY4fQgqC5y6E
7U/y8EQtJWYznemdB1xuh4emjps/5PYs0gppd2WNgb7N2F//MwqL9aToTSDfwX5i
Cch6WWHSPxLnJmEXRbrwOulfEmS6M1b6XDaQRkqEgZ0ch6tlttWUp2+AH3H9daJc
YVxmnLeqI9EXtJbiem0qkgYGxTeqyRpBv94KH62r6A19yNoQt0GujoVvW/4OllH9
FLdTw+B6zSR0eIe0Qm55EUzWky6llp7Bj/1Mzfqwk0lJbL64kOpA40TeErxBIvyn
rzMCP9uv08UFl8GUUYF+bGlNDehP7IrtSBNEzAjnVO1vB5tZUyqOt7pBZnBimD4k
CcVuofgNl1Ah56avn7Gb+stWtghcwC1VaMttWU/15qt1mz4tgCDhAAqeyIMzYSB5
mMHZJFYXCsFm2bCKPo6BnH1zwT8GsLhcdYqDf13i3pLbn/paqAy8Sbut4X+I/gPh
c4lksV5MRFqIFc8xJA0qf292Kr+zqZ0cc8zA7pcJiewLgidyYlC4dOWE1Kj1UQ7f
o9ifjYFQsMMgfO4RqbWv0s+sjtTufVNwpYaPtU7w7cNc1NlX6EhQelkMu9JF2h5P
THeG9b0Z3MXXL6kNj80+vSbtFvHXnLVh7FP44h1b8XDVFEYEHUo6XzeUBLOqA8eV
3dbc31K8/TEm3e7jGodn/ystZsVtv3QZfkeHZVZR9eT5aaZv5WSXsIMIAPyEMYhB
ilnBaIMGlTemWlOUTTmtgS9J2xm5JuprN3Q366KYZtWlDtidYZ9KCwCWAWMErLLK
pZaahqPMUswzUVA0YB2b0H2YoBKe6n8h8Ky+t6FdaE4SnOmqEOY+hbJGWhKo4XyD
c8nDn1jnfzKza+rZUwDqHx6iMmyO0nRErJ8dnroDQeILgafUkKBaqKjC3kipykLK
iJrpDBXJaZ7c6GX9gQ3BfkRUk0YGGe0j8Uv9gltKtOvQW9l250E+ybt+1DyzGhty
W59tvwmfH/sJ5GOw7ZlW9yKa/hhjLMjSrt1SgyASpnJjUEfGC8QsXoSXHNjRSpXR
HgzlH7TxWCYrnpzXLw+0UHoOa+1S1bl8ioOosj7SC7UrqhIEsUNk3i321m2xBu+D
vwGN+GViJiTYS7u+ZCYiUuT7/9z5Zob55O961IN4dTEOBF/7TYu3zDFXWth112NT
lJRN1qiabMhf0iigHtpO7x5XnVbl7cEpVhV59YOGFB1Rm78er02mviVIzVsnadqr
uqgSrWygdvkmnFskFWPGPJ+pvD2TcXWWa+O9zzcsP1GDhaKFutwpCcMIInYo2xE7
m7AbiV3bGKfYgBaBIlNT/wI5ABIlo9R4wxQTMpiBtJjyr7zskr4k+TX2CpLmRsZD
xEpalEXajAjTNQBcAe6NHhK9VzUFlgERHLuwrKeThX6vlyM3JqvLLAhsv2mmproX
Xj2kSRHjkCS8WKBWgC0Uie3YXvRiA8G0yn/iLGLKIAkPwzP3hUZ7IZfPEkXzw40S
bINLv7/TDMp3HkJFdegSL8ENrR9XCXmlGWLN/fgH0l0WF3fMuGv5kYg0bnJMun44
hdwXxhY078Ttkp1MeqE+cd2e20VEbs1wspQSCTAgZmduPjKniKoq1sWLRRg65mX3
Kfi/qw96rG/25JvTdsGTtYMTnFaX6sOD4BilTv6qxbj9tlE/GlOVsnKpj4FAkZBq
akqCI2WZR5HMFqQyni/uZ6gXntGIDnYB6WQQk1JenTQCS14NEzuumfniEJSBx0VD
38IP1ofRKag+aWdNMtwdvq0nRlyudBkjo0NgIDaIRbd0KIqOSkmRdcc6gAV4y4UG
PokA6BkmE8Kx8Cmd6kN2qsxB9QJiVtAuafzf/LK/Q8h/6CERdIV+DHvhTB3mXSnr
EAVMI3B8gA7aorMGwu7sR+QZumtNCO+wPZqMwzDznrk7ABZ12CkpKX3lvHTD5uRs
gUdu0LIgJxvlcRKFXWNBcTfADMKlb4ZAhiGYm80e2toBzxnzG9XHCct4v2napuxm
DqkTAo9uulg2TLq4wwJrKfP2yyW5sajdFSK+dqWQ9xbJXSYz1Qaa1uWwfBvgHi1M
Vc6PG0mJUfC6LHDFBvenfDC6CTlQsbB8kc6GxgPGlwuUXqA0YrgCNMLZEQAoBwzD
mciqmvxRyfvupBBiEXOZGEkpNCQWs5QQqq6TgGHQSdk7gJvlpwRPTkcgpvlmTfJ1
7ve7YxClkvGFCjyLrKqxGs8QNnLsU0YNFDpRRQrFYWl8IyPJY2YQr+OwSFNvTJ9+
jUe/11+t56o35XRjxFHhg+53oxT6aECoOcXfjPwx/uuvyTlbswHFbM8elAJcQzFk
WSWzTmsjoPz/dFU91MhnXXkgGCIZviHm7e0plgWTFMU78k8pE5Mu+31o9mc0X+wQ
MSo67h/L5oTc2X2pPk9kMgYfnih9SP7YVc7Q+Xlw466k9/jb/sPZzCKiqvc7N7TZ
WagbZJpIZBVmLwqNcgUr/4ijLDwKhLIHBdZiwc/v1zicD1cF7dqTf+sTaIzM80KS
bNgMsPNyIHedy0rkPe/YnfgjV5vVlj6WMNEvwer2G72bTbR3LjSG5lqG7waVAUHM
eh/C6pc8qa/qDvnHKdPux/w+SqH35gCI+TipHvxtbC/1X5o5y2eagLZmfbq8c/LV
tnT3nexKdctn65TV9w3i+fMwskjB0IwfBHgFGfa2yqpikPbUWcsvGyL9t6f2Ap1+
2hFyFpMlud0Py9Q0WUQ49uaNdPbW4+RSZmhkrJ5GAeJPhd5ppEk9uLHcNHIvYj1l
jatRgx5BzbPmMcLVZSC0OBBq95wucu5mpgl7nCIVY0H7rKWnkRozW6PTyG3JCodH
p1vaQYNy+B5xRV7Z3bk9C4p+A4O8iY0odXHfkzBFvs11e+1M0fTF00HvRZgcqW8Y
v3cUjzktHOxj3PkZna0MM/RKyFUsKvXowDnx7jal3cKDIrPTuluGieZs7X8NDyqO
7KWowJi9YR7U+MZ5YEhLOV3EraegnmAOILEfE0r/YLMCvqZybTNIzOklqs3BEeoy
MFsBHnxEj3fiC16r9EWm55y1p3h66o0pBQHjIo1RGLDZeYw9GlXRTPhCQyRrFMBU
K4VYHDz3x+nyGDOyB2X9ZKbri3d2e226fVmlCQzEZIb+xUlGMC1Y85R7EPwx5o5U
ZP7hRsF1H8LsZEmTr4UGaprxIgOhKKJxP7X1s7FuB8DME6nwIpKqkK16rj/KlwGd
tH7mqSZOMh5YurDqO0zrieHlViT27DsknH2UZ3WHMYpo2CQMrlxq1Tbk1kHbdQsm
e69JEXf0hJy4RTKHK0eN8OCqEwarH3Mh6kVKXhMomo4FOwX15cr4LW0NOZVG7gwh
noe/xTgc6j/hSh69ivHjayGhlTypD5P1SXp0D6kZOZ1X9DtUdjnviOUAd9wpcD/p
mtmv49P1augalPJ3sI1ReOP6kMpeXVKOyhcBIz2/L4hmg48JLV3yUaAcaYXMjy86
hnJIR1Qvo81YSP6YPBu6T7BZxpFfd0NHwBqQcTigUmljYS+nSY/ENzhyrRlZCstN
mS+rDOIVKNcFCs/a+Q0TJ7lkbID2HX4glOgy/KEtSVB8lOI5m2kHTWRj7Xx5b5BR
jD0ayT49KQn3AqImDBzo8ZJb2m0uqLL577Q+ZQeWfRg36lvAChJUbH0F6XGj/EQI
We94x5WknzPBzASHgu94xHYACEitDhe7O5NqFMKpqLzZInSeFRXFgNq8HhDSoYEF
TbJtxEtzcc6dZu/4K8pGIkvrdkpzMJeGdYmql3R7JH94fACMxDtiT0FGMrNp7jIg
2XXcA83SfwRm1QAZ26ttJtVFTxxrwQbt8HdIHkXVmWs4iOb43OnqRZL2j3XGwgVV
sN8Ia6+XzDGowtIJpdWlqfpktccyC4GkwIeVI68dRUFe8zV/QuEEDmQAH1/giPPC
AsOv6z8rO6J/i1zYaFNeUWZfwgcxqyqS61Za63NkkS2ZwRnpbhcJ2Ddc86+Fq7C6
7lsbqlnwhpU1eB98vNqkErnsb0CTjG6lBL4xVTHRuMhSv6omFOH3GLn5X4m/9IgT
TAtq0ankRQr9TXY3ONps16rWV9+wMXINt90FUqIud1+vUJbJGNuF2eEkYwQpwtu6
camBfa1NogDYabFfvkefEnDGvcEjO0zP28+d4CrGFpGf5sxfn0//64+hI7o8/MBb
tZQEaFkIgQLOvgmCv5pFBsTmb8X+0zG3VT2RCV7Cw7W4qQG3UrTeLAyJUQEtBeR7
8to8w3fV0n1S/yLGdzGmqKSpD6ltzm+eIDhRfJoOLgaMyALzgcgafaNwaDGFAWsB
AyKRiuA1OP5cKJTopFC9Up1OxpMWo6yGP/GTVxBzV1T+jQfF2UYs/vyHO5nIbChY
nJkcsxZkg7j/9rqm6gb+MKCaPflmoSCZz96LNjrfXJWdJZkpsCnpzqrMyxEf6RU5
JKlHJqYm2a/uq73mDlEvcCuhFnRRFpJoyEHbdFKE6bMp+YpV9rrhHcYVvOxONORA
E03T4EnUFu8FwA50TDeBlZE5+/EeEbp6q/2y23TnM+nNVNgziSlMakMRw2zZuNti
RqpsVq6KZQdxXrh8+Xec2t7kmRC8OjiL+TKxLucPy1n6rdnt54GrMr8o01dJSjVW
oTqkThj+x+ucUAQuBERZ2EItZkXm3s5GJMsXwpCiYolWNvCiCg7KOLxDdMa3JyZ3
QC4UL9Hz+z6+SecfSzscVGFvAn98HohHHTn0AVLPkNTvQ1yZMplsm+ZNbWf5yaJ4
HNGnPyJY2IoAEJqieLOMzJG/oqLwlAmMmEyVMXMl9q+joGMe2GxGc80qbh1+OtWw
6FlZOaKIl6TDU/w6G9PoOXxgYkSW+JDd95AWFYi8n/UAuh5F+v73bYTEPBskgs4/
PbNRv3iCPnb0c7gnPZh0XMYTLEdKza5XVeBohkFUsvP9PJZS9ItwM5kQCG0M94Dc
jSzIg7g2PD0UE75wOwxYa1LINtbQ+9Yta9FrV1jEjjQ+nPCfADDnUG+hLgmsMc1p
iq4PHgf1+uHAEtqQxidU2eSAJfo1MaObbzTN7KuOGikpGFekaazOFRN0JlYcZEac
D3dOsO5V1NSdEQsNfJjyhqaXv8kRhwdjCqf0Ka1iClmVo6UNbxKTsEFPLU1/sXR+
OmKBjOgJdl+TnWyhmXhKFpwCCP2h0iMJ1j70NcD9l7mROQ5PaYdC5ptSp3Jpt60H
7/Jv2dRAyLPpLioh1UKOydU3Dh05lN79wpNZI/weRzJGJYjfcytZIBSQdUtHk0X+
puftRX15nHvsA1lRQqfF+NW7oU6eMrj4AiylXg9ndr48VUDjbHhoFD4LfjZFXTjd
NcNQ0aN6FOp0PzIfxUQt/Sw0i61QNn6alDWFXjpo0FvOqMRQjzdymgBgaBUswe5E
FAxmX+gYGtvU3oDKTjlyHcyXvEBGwngEWV67VhmLLwCK2WxvMKJI7xlqxAg0WyU0
r52Ctnd+1frZcEZoT0DsAgYbN5+mcZr/HR/3V08MyWa/F1pfRMdse87SQk+sUKEB
AX0jtXZF5r05Ata/kZTWdJi5yVMseat7FhqYDnefjUM1jOcX6WzMC2RwC2KzwvU2
gcagRjXyRuekt3Li7uTd1x1euEOCzPIQSkIJdMSIKauofT0kHGcWSEA3jw2+gk6t
EfaDU8AU7c5IhGyYrZyrWgofl1JK6LlzY32R8hvkzBTfhZ8S7Bo9ZNKnLmlBHenq
f61s4UNjnPYt88laMMvmVo/LcRHS7o6fxi6RziNT9repxjHxBPCPQ0lpqgAugELK
DwlCVqfAcpOvc+VWpL+AY7Wn47D+O6QyXHHjC2ro5yu22c1Zd3umqT9Uy11MxetX
tgUBRPnO4kSCrrpHqWSnMgJXFoOUBJeA7NzErN9dZ+hnKsYeEeurziMMfOiHwLVD
g9yZ3ia1AgBtOcIvTEpArqbQiTDTS+8ZghxXLooIaSjJBzoY5MoEIZ1J6bfpte6v
8PXhuQZHJTk3QzTrAat1HMcjx8Q5UlzipWF9B9r7aWYGphoScVDmhCi2R6MImbdX
kJRMJNNmhTXQ0UMaNhHuKFuDZ8v9BLZmM8vwzkIqeZoIz1s7YFssGIv9l54c/zif
v53Fgb2I0QKZPF26hyo3ahsyTVBM1Z5hDzjLC80b7p7z61HKZXeHuyHGxPMTL7cC
jbPrqP4OX1eBOkrt6RTHqe/zs/l1ZqKMG89fIO73O11jKWWRfx//0TJMd9fCPdT8
zVh2UJVQGmm3pi0T5wcR0CHlsZGYHaQh5As2K4wuIjQdGl4JppvvE11ZBVpWNZaA
cMtEJXZ2JMFJmb0rDzg2BETVCOkb0z3IScUvfinn6pEiv3o+YHfIc4yKYA39AC4z
PcTUEG9DjW+KdWr4+Umo2EHViO2ReJLnWE+OoVLhe7rqmQycWAGRrt/MBLdd42ga
tki20JUvOBXUXTVVa2bOkK1ijIxPjwdkcvJyoYEBQrGNgoGSFDaoRimnfUOetAHi
nJKgfH1mbpnrzHCo4/q5dsStLB88CnRiGk5RECeQItX2T4ZlIeX0ZDCT03Y8FBvM
QYWQZhl/43bZp94yjGXwsSuZJD/rXXp2/TyqTci+9FqxvRbkbpUuMIAL/BmICb0I
inObXQSTLNt+znvf9u0y2TTSmg6qLRoJWhmNRDwVP1DvXJStjD51ocnea3cn3nIf
cMGz5aF2iWOiHgwfnd9TmvwdqXsJpOmoeRVRNMbZpWa9NiMmR5YUhu1Z0TDR60m+
2ECpmMIaYsOOnH6/4SxPbyA5xcalOuzD/qav1QRcXT+36NqE3pdssk1LOzl4xcm9
EOq//L98Yv2YXZApfOn0BhFm4iC5dsOBk0BlH9Iv8mTalg1ZmEKesbaB5+o1UtLS
2ZcKvez1NEJb1ca/66hpEMWwrQd2pSJlWw2mYljwoBdiY1wyZvkgKc4Nx/3czy4U
20cv+Hg56x3vTjQ0sAD0o3AIqwmdUapXtMbAMQ/rRnbMnY2bzPcZeskUrttAy+4y
kkHphC+h8WBvZz0t7nY+uepFvJjchmDu44u/tdOWcWveE2GJaUYg7HOEklgRKeJw
ceD2W+KUlzvX3DtSoEKnpHGHFLVbmx8EPQ3+IZ7NO6fXP0gHO7NWQcDfla9QobWV
jfGnWwmyJ1xRuT59HZQnkpCNT5dQJj67reJ3jrKGK4VXV4gR3mTJHqFBqa8zEGTS
POGn9OORLFYfGR1Kk2qr4IdztTU/iyZLdSmYvHUDYc/6+ml32sbAsCb4yJ1q9KYm
VGKHu59tg+Vmy5lW3i8htf2F+iiqXII/dFpdRJWjG9YdhyUQ7FIkUNx+UghDqZdz
rlKHdgCL0idQEgWsY63p3eRsPFb9Sq2uDgRzLQ49Tl5l8HvQkUiVz8GjIInRKPAh
2n+a4kYVKETFZoIXgNhildHQdpSzOTD6awok5wH+0x/nx4FqrIZPFTh4jYwYxv6j
q1U3rce5OJtJSWdRNVw/AeJg9Gr8aEjHfAVaswo9bFyfVGr3NXHVhS2Cv1Ua7enB
mYrh5JN7p45Y4V3H1HWOyo5Mb1S7OisYmdgR9BUbWgMIZNKHKWg9wO+4zHdQljeE
qrJsglcLEi+4KMEjT+vMr++tOuDzlhPPcG26/mJhEkRTYjFVMKZx6jIwElH4u9Ec
o+dSF4V0bnuFiEhe1fZgdL29M1zXGpd7jom9JsstskCO+LFRsInhYBLKAhfj7db5
WwND9hK2GXcUO82QXG+OkCHIqBVWSvJAhRFnobVZMvb+lRNF1DmoRkvlUPHFWKQe
3SNRyqX7Fu4GGty4xlFcjdmO9dU0mMbebuWg5BkErtoZ0S2ybV3j5Af2uw4vjGYv
YI2dtAeTgd8KTSpeulKcqFvzr/oI7SZ19DFy/R/71UltdU+WE9JtvrPtmszbPzux
ekZXHXYDmmqQuroG0jaP3U4odPag4xYwKwr0VpFESpZm4X/okpCiw7G07q73Y312
rm+vj87/ahQfskpvuDUhW/tEoKDnahG7YuTEh/3b70yphsLsGNqgPqydnuPQ9gOf
CbJx7ZhE+J81UJ7UrYu6NnyY109n5zm+l51lmTiV83ZAx9u6R2VMbhfv++hcMf12
pAMWDj4VwRv+uQtX6NDTWIKtQqbdzeR/wjzBeWwR6mWDhKhth0R+ry/I2tT67/hN
9yAdniCG+x0u3RfKMvIF+9CxnZlocVEYBeNoJYxQnCOdxi2gsDeGt7bgIs/+Dd+b
AZYfnFXHgk6PVERbF8msg04Qo9ouCwbJwn7RF1jGZEmisTEmIs5/wIQO7C8x6/PG
XFjntjsuGvjwf4XOob4iMOqZYhBSOYQVu9CF/3gMCDV7qnIaVbS+uqb5+Kca2iwQ
Vvn4+BaGXh/fSsQqvuwlGo4xoSi1T0ymLdfz9DfJaAH7yX+vub/q9TSLNwEEExhG
zpnl55p42PKUW6dVQa9YhTGglahL7JZtnbpNBSR7iSVAQJAACJ7e++geI9I5U52E
iL48/KTDeacU/kDcw2vjxLMo3+j+cgWPo3VFqyAh5kgbdk2jfsEaY+EmhoWMN3Zh
29SH+WwOXJUlnvBpNIA4+Y1Oc1saFrn4RHxP6tBGGUajCc0+mgxymvEfa96ZACkQ
b3RRI3fdUvtuSM/LrZORq1Xbs8zVB1AYCft6FLtwcDuEuZM/dSSfMsdOPXCUsrwl
hiQte6Gm56xPc0QX/b0p8VQ9YH0SdU6fTgPLBaXccgqNWjhCarT3E2hpKuX0qqLG
h+BomYZxxRzX/gBpmgWxdt78kFbeRbdmCS7kJd5hPquZso0Er0xpGcIN3iVrhrD6
UiGTnQn/wu+wWH96ZemMP7FqHC+5ytAdBrzr08nNOX+osUkWlVCdF/mja0rE6+R2
wraU5cNvmaQ8M9lFNPrnn2Ins5IR24YZG4lwQaddQCgyU4t+syuEVRnJl4b/fF5L
6JkcvnYcg4A2ZcmZPiEOeFp1DR4NwxzpzXFArgqxxYFtxU6rGB0PPdZ26Wr9Sr3X
Q/hI/IdzZLsM9wl53Akg63xs+6mAPvV3EwdpiKRnBmw00XomJrt+NVWRdomnTu90
ZqQ9bIg2sdEjoe64aGh0lEVbqtrekHJF3bfzxYQR/EEtYnnX5TUhNpRGXEO18mFk
KDuovusKC2BznBLTa4wmFrfdnXkeZWUaXg6PEiMScZSR7G7RGmAy1sFhpP9VoLo4
irjGG2qhEn6XdQL1owI1kkRyRWvHi7naFiSzVYrNjX3E8LkMk6E2GxQZsvy6mrEi
GXit+lgfe4UeG6XD7jczpkzghZo47UcgWFKUVIDaA+ffInm9k9O9cMWXW5K3XfNk
kDfcF3nkxi6XcFOLUhs9YScs+E67Ikfd8NZDUZQfCLYn8f39phPmXPkcbDfxvHm/
oSua7vpW1OUnHsCpJvmGnAOqDcfYQKi7vNonkrcLxxLyI2x3++/yApBveUQFPZFT
XMUMcmobPmWVsNpgBBgV+Fi9Q5dPCHGRpI3jZHuTN8w79X0yiafVgdNofA4p0Bp4
4zWNGKx7fITT/iibZkywQIZp4ZDhOZ0sRyGotPZESQhuM0vqHfufziZrDuY1Xpmq
ghnFSUsvOVRfkp8w+FzwqhH/jUL8Y23vAw7I21dwoCDrFkE/N7dZAqJp/fKcKpzQ
Wh+1oD3KMGmtYqOQ9o5Q99FD9zH4Vq4rrjGKjPspAr5MUPEFAl9LGdqpt6+WmTOw
1UAckWQpq3WjXx6+QEBMfWGYa6W+8RIboFfyHgIBD5XfshFJj7ZlcNG4sWCt/4qq
vNnq6u3OX1vUnYPpmgjjsu/4oFWkLW/muklBK3r15BeQJlNfVG/SAMAFgsPiHp4O
M0oGdx9ajVNvssrFZk0epWGEOnkNqATehH9oWghc8jZ9GM33o3oZ0KvGpMY/s3wK
7UcSjw2l72yRRGH0BjL73bIKsjeDr4v648xx54dq8QIQ1AGjzWZeRQT6IHF6s3Ls
9GPe/QINt2l5udLhBTMTP9m8k9IJsXoTbWDjsfSTtzFYPmwmu/vnoSltXYYpeRMA
AdjZWr91B4ydCWK3f77bYhEA9Vng8c51UkVksvaI4b04iYb4YbdlPZitAcb8Avih
udBg5UTqJQpqwJkn2cbMXvy6BrScoCpP8hzJjr/+HxKN1pkxxZcDL9tSb/zrFGyB
GxMhGmwHjcjK1Dt4bUNscYmR0xeFIEEWtpD6lwHD0sFnjqi2PoEO495hDsRcok/f
4Ya74+96YkSyymA/eEQPIc5yCLuQxlFWxZuoDa/ITENuEAnsJEZSEt3Zl5CHGD/O
VhTlOy4/HwmCIINBoZt5rajY3zonT7fsRWZACNydYuS5AhU6WT5FFMowjUNs6qI8
YgdMe4NfgRMJRVRH3IR3wrZ5fqM4Y/jV+fmfICez4+p+TSFldz3Pfefsyxjk32Yk
XSTzIjD1W7A3FHYmjIcC0bWPHhWyXCpy5UeaWT8hCH7l6cFAfQcgHlEuBCBFSWbT
xT5w/aMP3B2B53rXRkrLW3ZIO25pQxl0qftCZWIavwPTzFTJDYB8PZczlkqDd3rK
ieA9iTS5J6Jk4dSHNJKOi9qeIktYcocN8rH+im2vO/IH7jEzANvjXkoEGRV2ohx7
qObJdh1GO0wK5kFyMtG9qKfRlko56az97OmrH4GO9VkjnFx7vXBtDngSwRwavGr7
RDA2Ip6YKQV5tKieyYjs3WiRJ/WohrTfes2t4de7HRm4/bNvmywwQXUEEs8GiNbb
sJ+EUFdeHfi9OdS2u+llGYGsjoImXPFPSfZEr5mWMmvdhLvJhwkva7jnlYR0UJ/z
Hu17XZyhq3mdg8OAjqINL97BbjLC7UMqUWlNqmNug8OpKqaw0Ahz3ad4wD2bxmJ9
TMdDG4Byd+BbZkJf7S8F5w9ufZdhBHo0WbwjWjqbbu8OBXN2TLHyN+mNQUoF5XHx
HXah/HqbuOvCV+oJ8SYtHViz9wWoOFOtg28n0a1UCOFLi/eJNPy/Sj78NXLWuO2y
48aG5OOYnupeXQGtxG+8W4+ior3sh3twD0Vsk33aU9/VkqwKAQocBhcovrjPtS0Z
pqWs7FDZNaxExxVe5gOyg5h+cwCRozY7Ru5TzAatzm+6phIkJLEuXgAJO5Dr77V/
iBSJwfD7/y8PYskSeNiThhdiYqIc7mbo9exo8E3YxbIpXc34Czg2y2GhF1O1OsQc
tBwIYpvKAJIdZgdUWM2bozDEofWia98XTDsM93T7DElrypH17WIS1v7udcbVjGpN
R5NGJMe9B4SHN+XIjo96FEAVjqxT//fepUxQ+zkyBN6pvsc73bwMKXSZFSKXUqFI
sKnjzMhUClOTg1R319ZV2fvS05zEyaSjDMzHSvR8ZhJOhLqYHCeQJXGl8yEVxqYq
Y8TbJq2tMp6g5YsUIb7Ek27j62+3aGgAIM03H2Dx3N5nE+gLMiCAuTd3W2n7h8zc
IQbg0Wh3LZv/sdsBCKI8p5teRYQkIY/TTn20Aara16zcI0MCZ6t+tC8RkAh9Kcpl
ugV0V7TqgblFmizL7o55TNhyTiPZgVk/dFiJgY18h+XUi9eY6zSOu5bv9Vk6hMKa
CHvmwWkaLK38ECTwjtHGqWkcGsp+8EzaB5LXQ5C0XkpGeW2bcWqZtpFc0RlKsqIz
i40N0yUXAjz+ExzCdPDpjs/21KSysCpIpPQEokQHizFPVmG63s6DpcFAWqR1WR/c
JU35ADqO6PyXBsRFMLyVzL1Gxmv9Gy2K9NaAAIAkIYQmb+cnxOxoqVQZk4JD0ahU
Tni2JX9CZVwNp4tGtEdhujWMP7HjcwxpybtUTVkJj1rEZmDiIKyCo6vcJiD81wBr
avGE1yE32vlYKZLrcpLAEYKMvwX/ExAp3SQGSKXTk9UWlo4VI7i//EN450epPQcl
0zMxMrdsuS7UIut20hOORLAz9+qSxLtiPorUpPZKr5zGoOrNrvMbLANpJVwc8mXr
iCk2JrvfsggaJR9OEz3dx4zMsxGCZDrSlwuOfz8BqKDIdKaxlL8jFrjiZ2CSfjiO
1nAGte7NrUvrLxQrf7N53igcm+pamNcYXsNiz7dSOathB8cJaBmXM4ROxQD0Mwif
mAfAaD/KK3RFYqtMPdlmZUg4KK+R2EtJjVjnAqvjRddc9uVKawTZpdOf7BUHVFsW
V/53KSgB5InxR4ygcUrl56ZKOBO1YN2FRBPwi2ehBMYereDq8tccyLpEIP1lIc0j
wnGK4OQ8kKzOGhaQoGwT+bEI0oeJRW7BIyctxEDj9yUhsiPLHb4eTZp0ty1YyZt2
Z+kkaiTpbeBS826AS0nPVPd8cUpdWyJqA4C+DkD7Pi/LsZvyRddu1d9pdRqK+UH+
BARNSK1gHD8cu8BZoj5Jr2DLqaUEB9C6kaAQNU0/Gls7I5p/CTCjedmvkMNoqcKk
v7bZ1r/pWilJZlre0DT9ZkrkTagq+a4HIMG15wLFz4GM/+qy/6w7YB+RwwdXyROx
99tI10B0TURImzzrw12ZAbbSmS6yXJsEFhApQMr+JQZitd7mcEaeofqYuBI9uNdj
8wD6O3N2fLiRhydsfymyZZOGYD3xQoi+1aCZbf4INitIfB46PxBHoTXmr/XbGJx7
/IYNemtHm/lTJh6+tTFPKeiIWBz/gqyT3mzPaJOH+F8RtrtaMWTA/VznReuHh5d6
PVYKdCR/XPX3zEQLK86ugkyZmeXAtFKK6Ogtk69kleYIIHNGXSE/9J+dXyHnT6PO
wVc0+wvJG0SmObQXXF53qjN6aa9jXq9NQPc2ZRs6IbHt8n6DNqW7s8JkJIwivwUx
2t3GHJj5pj0uop1EKRRA1SbtsCW3b3gKcYaN/udkg2UiYGvonG4CYavHlGtsLLas
AWpEN0iDCwTfYlPkdq34PEOcKnOvz32ISyjB4bnc/bPwLhP3IHmH7p6vQUqLBT+W
WXDju6r8STO7gxk5UqxgyuLfWIHlEoyzAaj9AxUkB8Sekp0m+rUpgrWDnbhFfBoI
ga9QjHiY1B3s87VhGSgdjmghYZrOfK31EwnJWC8ywJFvuy4b+2CHcf/OObqCgyDg
70CnNw50rQlprkR4NL6hK4FzdM6dsKCpsZ/w87gcgUQAy2Qn3hMm/wHS/FMpGBAl
GdxMbooDwlgtJgWGP2XornNgBttKX47SJ07cjuCK71V30tf+4LqN6DsWR09o3J6F
20hdZ+e1AfTdM2nINfwWF7uHWWhkoFrBaTFgPqZTq9yzjVcyyig12ll/5L8lQSLr
KaJoz1rZpby2fcCUzhvMw7WXxaLz9DKXrOaI2xvzrPdNWRsY1Lv8wc8hKEnbYYJC
R7UNTHjicO/S3YQtnbabEux0E/2/UgAf/T9/1dMIHICHoPC04vZHdWxvaqyWBsqK
8MtYnztQxladqtMbqtmz0LWwCrv8pwtxIj3dBjdt/QxDDEG8Ckg8iYPIbCdw2GQy
p/ywaIjxKGhMZalP7I3U28PuiQaASmiGjNDc8MPWYPslIUoK8lOus8gW1LMswWm9
3NFTD7rg0Z/YTUsWzOw8bwnUEvAmxsqAqgcuQtMeQC2NsmHitJZNJAvE5MjxcwFU
vGxSVksh82EByC7Fr/UqZOxUx74913zps7vzwlRHjQHsHcYU8hOYxCeIVuuV0Tm4
yLK5GsGdTPbcCZAd1RXuQVCRDMNcKz8UOKiHEc4t5/TBW2fJqBOfjjXHhle7mhi8
bwvq6O7WECSZaww8qP6OMQFkFDfHQ7BSXoVj0CV7bjNLQg3jB3WrZft93gTZrFUK
KACLEp2OO3RpfgX/azAddgBUw5UeWUNOY3izRysEjiw7bc2+tWadZ2mEg665m4On
idtvYalViZccjsGMEGBdK78rG8Do1ZfPRaBYeuRH6DiWRVeI4mTCFZhD07py6hKo
ndCIN3R0kEFW6icACcJSk4K3ByNUxS6bGLaCLtAUxc7vL/1xi89AXCY9f00hp+9W
gKxmvdzeRvoBQvznWUNiVr03jfaObYx7l0cgPJ7lm8CUzIG9vRRiZspUjPRWOuAx
y+LcLR6d49a4E+iUaBT6Ma4PyrPbjij0nUbZg21iMkRi2k4wCJKSLZifKcLLxDvN
kpeilpoRHxvmF7IMMol/Da6VDtTUl+YYfWWvHpq1DW3VPPiWbYWs5vpyCwsiJs7q
crywcb7j1G/gGx3PVHH5bhA4hetAu3Xu+Uer1S9pktTJOH2PvN3KfI7GLDS/JSc8
3myjNRGpD0j3WafdbFVn5oHxxDbX6+7yHiLheGW/8mXfxKz3re9aZKDX6PC5JfWX
6nZ3X1OxWrqb5TBT8IIgxT9H29xxr3jM2Dl7SaTzwRvqsNqNzmVct+qundsjUZrD
2tpDFDO4SJ7CnmJwtcpmF3YTk+NaQ2ZVWJqzeTCvUM3NQ3zYL3ronjNj0iQMYENp
QSFDkod/zsKlGwIu5gzmoZyblmtMRU5LRL/CPqOpJMfFS6b2IbFd+zD12hUCj5zg
uOz567UWi0EFBT/LiIktZTMl8kR4LhufxgDb91lP33CDtSLnWLboHhns8dTiZE+H
SfhGdGiTZvn6ND2u/aG+keBvlPn26XtQyIsjzzmFo7gkO62lgAi12OhT+ppFlzc3
dOUDzj35UzChaObW2KMq8+d9P1GnfR2Z3yq7AO4oRmh5YQkPcyQTctZ9vJQvfqmO
Hz5hlILRexLk3B6Xay7cPNs+rTQnQiuTNgs5GRsEV3tXvTmtOyL2eLyKc7IJDQqP
BqaT5IPGR5dVg2zE8QWEqC5lSLeo7YKiAWLU03niFyM1ddsOXWsRYskMnbPV8uSx
BEhmuGPXK18pFEJhr+ycsJDKEuAKHFsVeYPtc/c08fp9/WHDlwHl8vJLn0lciSrW
lD31FhghfdBBHm6zuc1WYu40Ol6rm+IQozth6MjrZqey/u2e5LLH3s+F4j9E4Z+y
b/kVqIxJjZVPaiANapQ8BNKrf4aIx8eEH8xuuGouZHMP6xBnnygpk4G9FozifEsD
lKFm6rRiGrxfBDOjhkBzHVHkVIg4dKs1tbf4AK9qy7fEj9/U0TPEL8tGnWfKYOwn
A/yX99aXQ+A/wNfYvLdfkCJKaCcGQCiKQTbUu4HfmPehJqppGkOgUTumTWBRnLnN
3z3OnXWfyroMuf6A6URlgIgHb+34LwoBN/4sGzzlgtZuOnK6x5pPyYsbcITg5qSP
7BgduPq2y3xfHgnWUGhEsUWY+r1fMmAXX4VYhuKUw1F3dsYQXrOkoBDid7R9PT6A
g1Fm37ws1sXvR5kQFrIAmihzdTHOpV3j7+xDDZUIDacT9VVgXN2slmM2tGytyN00
bwBYGgKIfQzBEIEDCRVqKQv7Bhlaw4b5NfwdvsVG7oFdwKrORM4sDDeWF4c4JYEA
5/PTcdt6Fov+eleV0b84ylPQYOPCfozWanLj/KJE5FDPkHzdwc3+ZLivT/NRk3GG
+e6hoet4IGLl6cxjZq1GTige1yKYiz74DD8P2ngdzWvVbFAPReeQ/UFQ75oX3EHR
10r3uN3FsjKK2xmATGe9jdcTmAM7mGwTFvf7xUahnf7rN3wibXCZLNRCEC8XSkJ0
wEBV6TkOb2+q+HWfmp38dmvcrMa7cnnn+uldIGfnA82ZdNE/T87Db/IsGe3iddBf
M16aINf4v6qv0aPgIiNMDUQnqH8NwAdrmIDRm0V92XMR0Xn1XL2SeLUwVzNw9CiO
Y+7VRQqx+IYl2oB3+ONU6eyR2a0FcSTQF3Fq4RLmMozyB/IkwAijmFeNL0Y4dXJq
/5/jCASs5LOaNTYV+E7kunlEoLSLNJZtaohvrX8VsB0RgGQ7lMrrbwR4kQh/ZHD+
FZC/snPSurkexHkSlR3hC7Op3f8C6V/leItWMie0/dAnVBgbcktL0a/pVP2ONpCg
Qt0gUMXibPG+i19MYgqgwV9sJdCl6PMARaAkEtAIAXqq6hAlCADCZNOPshd9eZpk
PsSOUCpgtcpjd9olRXg9loWm6IlwUog8aPGy9MbNsOqPUJczD6vE1UIEll6GKEsJ
GVNADllnex4fPwmbyQH5FZe4tjas4fdcFxmkNJVMTVs1kgRpcYTMbStV/UUx/I74
TAW/t2VUnLdaEpphPzvIAu2QL5vXZ/LM+O2VZf1J4N1j48QOnQqFf5VOT+EWnBjH
DN9ZqFsJG5LfMh1ciXs2KUT6FYlccNrEW4z/RTJgbsRw33tZJfyO6oA9zfemZf0r
uI30R6ywpBfxTYdvHWE49fGwxS/wtpjZjG87ndyQ6pPav86FoKIlcZuL8qaMBuUY
eISZNKWOxMewIGF2FMFbiOmfW9OdrI+z+ahLATv0k6VVvlUcB9uxfEhBlb6Q9dXd
JrXIHNZMCpWT9yBWJl7NuerBUjsuVJ9vVJRn/OUPNoVcZdE5exuf21MV+vDVs1t9
e0muhynaKJxKts9zJNFOs/ohopxFmfNy2cbFdbJOsRvXbomb9u109rv0WYIr1EVK
Ox+1t7pQYFvNGEcPoCIotAjknbr0odfrF7OhfMQTYXXlNDa/3Y8eJeKr0jzP1CP3
lGqCPfXDOQXhhskn3Wfx5MqNlBd3aDze0URafvF2JXiKfVSbVSZGeGRiMp19DVPs
VQJysJ1RZoXvG+651MBX1IKF14tfSw1tik7m/f2nB9+5gUrnOBvh5G58HXe6lsHm
NrN6BkivzAOf+ATTG0qjd1H+CiA8vuJKqeRYqoRJDd4cl49o+Utv5MYdHtBAmDhC
FK04/hAnLVDAa/GgC3rvneiNSs/1d4ZPNmL0AG+oDGH6aeNgzJKi2UWUnGH1sC9e
/ktAABSHzU2BUXK3w+lW6a2RaLYumt4K5UmYng9RMv5U9RghTYfIjTbpQzCUbEmq
B5v4u7IQ53I0Xo7q+OFjj9E3X5QlurXrN4V8zRrXKtrH8azxP9wn76YF1ZAwkSbd
mOpIICy88/fmPGL7hra1UO1dqyUZIcajw/BrwTGZldLfN/NzEPOZNCc/h6bv4Eow
6nCbd6NeCG3DxK0sRD+gOiDLm4XEg4YUDv+P/Fiuc+9HvYbvtmqHikr0lN9L4BPx
wwDhtBClXtkN6eZMeoQYgxQlu/74UkSzgxbfeB/OhssAxlxsRYVgZk4POkW5h6W0
xiezfRUuu9TgEoC9G3M1HqJ3jbMOK1lo0A85tt6Sht5TgOzYjqLw3VX9Z7HKiJsg
gE1fml/JXSQXjUb3v1bDwhqnUaeEENzDSUIht3eJIvB+wOSbn/LXyjEM8VLRu1HN
mjFpJGFnSJWQ3JVFvwbke21TM9/1uzRnxjnB51mwpv5ypEI2y6hKaQYxayVes6i9
1qz5OIQD8wVVXZsUKgHW59KIwkV50VGo+dcHqUm5V5NBfE7t10z9/avhjEiTw9Gq
uPhARdZHclYRM1mS0SBOXbcHrlD/rdNScdGewd7wKPSN3QX8jCf9PoQJ/1mHEvBo
yzbTMHPEeY19VywTgqmoMF5tUPKJAorviMawp0s97mt8qeL2D60ppC/7fTvS8O1C
efqQTt3tQ7wxOsSl7LHO4IIVkHMZQlvJC44klTraDld6JVlcWDmIt2RrOSRIghaO
dOC4G/N9oEQ6lOojR+j3GoGFkMTjYKGIoz+FPWxsTU8flOFR5T4HSvdE3NfiNKW8
ilDNY+R/gSkdYwXOn4nWSyGJlPCZ3ZwQr8VAeE1X/ZNMe6TrjSpxDAzeyaqJJXLf
G50LygdKXwHyADY1oM4Ldaobww1YQnDPBj9re3z8mTQ=
`protect END_PROTECTED
