`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xzwdxRS1XskIi6LnWvVFChrNRtsqfhBgkX7ybISZTCsHSBxaZWuXFiHXClHa0KjW
vGeajHbDJCgTqb7eFN7jfLjOlOcQs5yWxV0fZbxqlyeaUfAvgxzp/kYAdkfHCs8V
0Sp792HY7bg5ifyCjj5hsHtX0cYjreCMqVxTqHk2walBHZpX9gBRmWPkPfD2hCQI
Ml5vH7xR+236E72TbD3SgGaHTviWkfEFdVn7uRRuxHjCQObYN38QnlU0BN2Diu08
5F5xqy1Dgvi4HmcaCRDe5Xc6mIFQzN2MX5+yRoUMO397FRA4W5ts9LHRq1b5nHwf
R5UIS8COQttiorB4OfhWtzauUfb4gFYVGHxWFutQVIFCXw4WwcvlCLR63itIVhv4
j+zbRciYe/9rXKipMWVhk81LUApGyi67dwRvQ95cEPZNQfJg+zuaxASRMUud5VJZ
s7CUMsRMiG1QXA/k8EMUQnQtueLQXru2HIx58ANpd3E=
`protect END_PROTECTED
