`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Djh+mhMalPDnk4kqPalz0n3mGf5TDlIpJFT6BCHGxjGO2gLARjvVsRKYCa3gGFe
f3m7i8MDVrbaiJeL3MHhsjgOU8dNjw3oxI4/XSbGNsJpr9QUBvzzrNI8opvP+gjz
zaLXWvTV/qOyIgfMnL4TFxLIYA/+YjPE+Esn+EJKVKtrb7S77GRmsQwKosW+Fr1X
PM5CRwAwphxflNLcWlV0HMb7Do1ttrxpfFBzq+aAaAY8eOmOWDPY3qpAhvHM3rxb
70QMa56M20pMu2SWaMYLC684EsGeaKxut2Mg9HrGu6grFpjPP2/iKmXc0+2OOv/d
eOb3S8Egjpoy6iWI/xDiL+VhX20UB81KU5ZgJdrBiQwcg8WTi7dBN5loeXcPSM3K
MXpiFPMCqBG9YJAnNbN+zQTd+06VoOFwgiEac7znDoWkwNxEmUbca3jCTHfOUkEK
5baZgAl66zwKdAb1DAzKmeWheC67ADsfJdsHf8WqTDCUk8K5VL+WLnhXFjyNKwwk
HmMXldSW0NlJuwwsnMonjj+WddF0KAT94Xt1GrTM/sILRtP9YxAxNi0mjg8Yg+NI
i5H16sOuo1Si7rGyffwfPsWytKS/+RO/Tn/SiNf7ShObq9F92a/Isz/PYGKEp842
LZvafNamF9yu6ADxunOByCsp74MkkehRidQUWa6oK6E0kkW6LSpxVm8GF6koq5QQ
k1/tOXmiL55J2iBh6I0XYtls9z/W8c4xrIPqfvxVauw=
`protect END_PROTECTED
