`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xixyrz/PhaBq/JVf49EILimHuQk/9uejNnCOdeJuBPOVDSJXfwBH48MA7H4TZpEC
ByqvkuTNTpptDF9k1J6bTrQ3ixj7DrqMEWS04Y/ZkRcesQbYluXwP0x8Y8VIupJ/
6jn8+ZDfIMu0MMEwmDUkq3ubzOzCuYzK/6+a08oMGgNgkNt9DOpEHSa16qB0aCGO
gb/L0BgmUn4ULZhwpIU+sRWsFvqnnDUhIWMlJ5Jzy/he/HtTm6ZO1J+eQRsguLat
JHTYEokVvSVIikCD0WoJsVN+o1NMCbB2IvRkRyQVIQNUA2pVmsk37OXeujsm4oMT
o8rPZttbWW+H37eht8O6NFUOBpRwcduHWggAV7kmRn8F+Mheyssq+NE900Q7N6G9
IK/8mpKR5t0LQoLgfGz5Ag==
`protect END_PROTECTED
