`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tYhExTe8owtmZ3R7v1xERymRf9w6rD7MUXvCmrdG3RP8K+aWnzNjYgzqq1+gp15R
TavnZmkUWGN+2ld7mqvLM6ppgvzSRyQaENs0OBJeHmWOLQJ/kybYjmF875zOihfC
kGWfHkkkq0DSry+jcvP1HAYacjbbUiavMmE78xtmQinchIfZY34cPmeeZ4zQkB/o
5z3zHjgK1lL0FEljDcn0l2ikislx3L7Xw+WLdgsEyev/MHiEFyk/QEeOIX84u8mx
fIqKsAsYBPGU4qoN8EGl5Wca1kXRd3eAyBPksfIO9ZfZ5ShK2AVdix8EOMpnjvG4
QRbPL7BOOXamgBYldekFgnT0eW2GFOBYhG2ejfx1A1Pl3nN56DZC0vlLcNoWM/Bv
`protect END_PROTECTED
