`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g+csgaehj5WysjBIu7FhahAezXrErLFB9xGCLSlHPFWHkeqyYPpvOXy3VpcYj1vk
gUQSb8mhnA0IN7Eav0OBBXGvnIRP4vuZQj93tcpy9JiiNYoDMFBERV7gcPeoHfyL
fA7k+gRTrbfrbmaERqAnHIc1gEZJKdAWhBsChX8SaZWpB4YhmVeRoONafdGG1rgt
oeHoiwEyti9HEfqs5Ztm9XkEnXyFzWKGzqmECXPg0sHTRruP8KRVTKb+yehdosXg
LHqbtcRSI1LczfrV+4N5UrrIjHvX21acJG4SAXAH0jSoxYmqq1eXYMPbAwBqptxU
zO6AgUt9tqKOJGtn2qX8TVlkqZRh5ct9Jp5Dratl3S+suUsC+4kwQXLv3S8lbHnU
kiyEX+VW+VQqwU3SsDrUSQ==
`protect END_PROTECTED
