`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6dCb9/QjgrzoR1HfEV9bTnsjGql/JNZpJh2SdVWmg9mFNYn3vlvVIp0uP1hYh6+A
o2IoMnpPiCsMR4mZCHNfvJzyYjeRB6dtjmW4bhOMkMHw9N9DODnFQO7guvQlvTj6
Gu2Khsligdd/3JoHSGXVmxLVFOO81qZ25T2ghsKYEilT404KIjvA7BDWWYPhl0i8
C1Rn3qOZGipKwg9nChkuXOynRnRYsI6noX9dl1Bz7FChceDjWkhMv+yafVwVSMu8
baYSNzLUV68DjpdlS5ZZ24PpiKSZFxFlJ0klDJhsQ8/eHL80fNMjgLMEB3SAMTeG
NCXCtMBmFK4NtsLgxkAK/w==
`protect END_PROTECTED
