`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T0JwiD4qEVfTETgXgHCa+fh9XRyPRSK/WYKbXB0sVMMkKekFIHG5Nm5nwFCosfXv
9+yqw/d4x5PlqdLy18mxYafyVf0NQDNiyrFdmXoKAI4y0sSaxMMsbg1Zx/E5p64M
oBvdoInxZHKRx34R4saozHczoHDhgcnqzGLhQMCQA2M8S27Bz+yn9VuI10mqRAwf
06GqgP0Bgdx7jh7eqHWnzIu+6b5QKrYO8N+a3DUWvN+uwSIYWO0I2dMFkgpipyho
ILyAfOLiM9UvH5ZaxgKcLSbpgSnDciQhzKV6aWN2ZoY5XcSlDw31oapl7fjrUiDB
hyyc5pngUV3wYdxazFA+rj2EHyoA9yAFnIyvRoPTFKPKve+6unX2JgxiDblgfggr
bz5XBZOvqaxga12FHxK68m0XApA559MXP8qjAS5fIjw=
`protect END_PROTECTED
