`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AkyrIHs0h+6kwDijJl4AFqvguyH/2XAuPDO5k6NTSjMElIKQBLJ44nyez0Iiy2bh
AQmJhLTdshruQ9Upc81QVdoGdDTsxi/awVdw6hzuhczkGKLUrSwdtjbRRP9VtHfa
mFCTUlpmYprk2dBXaOJcXz7X3OFh6GNk0Zy5+7xZYXrqcnExjJ+4zBb4AlZK8F4c
r+kgGbEmfYR+rLStWBKdJ68+IAncHFoONKNycQsh/ryfQnebfQO/ahekxWlKyPxg
spkPQkoBeGd+4yVrpoyEYVsI4pT17YNzeXAcluGADs4CZozMnw1wRypSDS71MQv4
sibcZmoQ9eI2EsKZoX+Q9ESKmglt8ry95w2BLOsbTjIVCO5+9bMCTTg3uqjoxsvS
xqFUaoSOqV/42Ow0llWMJzZ6f3zYLZ+FtG0gWFIypwIUzGDM2QX4islpy8pTTYiF
N+24OeEwqbYGrCIyXKLeGMkW+IfVximXCuVLY48TCfmWWxJIqFy6fnsdSlxL1aCd
TauNDRYTFAqjMKtpwueQqsm01cGKz+huswDe1Y2Oxse4oIiNHjxiZIhstU8S+XYb
Edsw2Z9VlbBLK3oiI/rNMhq0GexSuucFglz5YDendrgMsPJrqY0E8tBD817QMAhE
IVoHCDDRzk8BUM9EcnhgTtSVdLuFc3IH3FSHkZc3sAj/mOajqIhIpacntxPoL6Ru
zazcsv4NKknZl2/LtGRUKRHTIAeOKH9upmsVjeOyE/Q18SgsQ509FR5EfLg5BCcZ
bu5n2fr8rDuhMv3bIH6D7wMQdOzoto7SqcNlOZOB/QG9qeBkJVA8Bjj+n2yTyhZZ
QTfmemA2hnLiWeqyUQvaaWaZA4Q3Zk342ptVkFDwyTw1rtVMuZa71MI9BUM5WgCA
rCi4g2KffpF0R9uAWprddzT9rtuMdEe41S+Ii0CgshsvfvTBK9usme006I8VNe0e
FGp1LOZw8h2RKea+jEgKEbvA6w+JcnTfmuJDiTI2rhJ9Oh8kQfhXiLR20YUFryFj
4zQjlpd1+4RykXmq6/ih35qXsUAkEajgpz7Xz80iT3FUrCVJBYMU4+eiK37YV2YW
4uTU5PMfZVZ9potZtSc61k7gLJ5gTP8YAooUDhUQ07kvQ0FdrrAHOkcQ5F07J5mM
3VIlyW5xnYbiNeJyFCCa5nakTQtTe/7DpxldVdM589kcIehrtLLgRyGTBnxrcC0h
r1ONFzEXSXcj4qnF2aurNjL+CQ5rDMUZ+TnHgQ8zNJcAkSAkLLv7oQ63iS3nBrCe
`protect END_PROTECTED
