`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U/gcvKqSiOPDfA9sbXWg2ryv5A3FF67FDD4IOTYLq0GDx/Pa3C3+jLEb6/5hsnaD
KEgZgZ2dshIY2oUnno3iMMzZeln6pFHUwCyjDHS8jVcL4lpeMtruX7o+Vo7WJiJV
p1q133kTuE1uxvQmaX7ZFSFV01HVsgOhL3/uWWNknmwmWHsCwKOkJPXwX+NuBOGM
/uFANufdLbmXxYb0E6MsVqF1sqFNTfdhrG6iYE34FsoD662R8P2LcPXrQ/ZaAki4
Cf08c3/fPgDdIDEkeYUtf6lYEpIwcRfs/uH8IWujTt1F59Fvcf6L/CvEyTwSXQF5
fMIlVL5E7YcjxGsPCCEUkV8n8j0GWwgiZrcKeI3779AUHqo0/LiFlhIEbYvuVbEu
Qwcod0uaOtfXNGQlSvCURUamx8Y4feSKj1h+9E8iViAgU1I7n5lfZ6dOvuDU+Igy
ac4adGE3JCKIiS+4vYrBDl7IsPoaus9NY1lezetM7vteDazFEOxWJNsTxBa2CLGG
Mpw+hBPBEJ4RYOgLoXCmfcQauGr3ovUiIhFQ92UxpOfCs+xItkfzc1kzb2za35Jj
0pHXiE8luDs9dz9vyVndCcxT3uMcbRpsDtH4FHZRXvRxhfn89HNsSyboyYIDCarc
l2xu/q9vBazv9uj6q6fpb+LRddbEWlJBnWVQlrRScCFkQg5dmV4YAF7uQuoQlVWr
jodirJSPrdyOqkI1VS18Wy+U27dBjgpFooz+PiiHlhlK0iZv/LQ2cJMz4YGcD6nz
5K6Fx/43Ajw2CjUAKUnp5gPDCoA5T431cYWPus3ycbYYRFP81sJim2K4E9+vKs57
SGicDBaNRXf7MaOOKySXjW4xkXdgA2Hxz6SQ+GH8YQhY1dVM1DRdhqUgrCI4fKQD
JpMx87oD+m4N6Xyy9tA335V+GoGJuXb5ekTCK4nMjMCmTl0aR88HkxZDS6s8lg6X
Pmz97ORyd2LVXcC97djsLMrntUfDqTujxJ9GRpypCXYfR4VAS6YFsCTS/IUVGjwi
9YJsnhw/W6P0I1iU6YDG57m5X7bk26lkPxMA8RaeUg6kh3WzONIhgX1jzRPfyoy2
xMAoBAZCTLFUUK1M1H0cC0TwPt31v2diurC9d+tb9cxAhF4q82lRBs6GTY0j1Bs0
GV8cWtUUGroHuKHcouP2Wqtfb9UuuOxtAdq5nQp+dBeq7CXXIQPJM9G8db7p1MFF
T8V4icrWCErqcHa7hNy7DNJ+qsAHq+uRywhe1UKad+7ViSYFvD4zUM6D2iMlkuDZ
bvdXrLH5LD/ZRsYlFYeAdWRDK4/7vYt3rTFbDtyzmetsV6qiZBoeti2YMiMBLDU/
+4++fngJGxKXmdNdtrom44ZEDMZSTFuAeJR2OjwlEUmgwFn0v0kBtNOYsSJvx/qM
IvH9kM8sUoY721YbgjkyzknaKkeuxFEnckIjdssxQopSK9ZYp6uo0yFj27qFTh26
MQMtkhtI2zppMf994O9pGFqcXpp0nAK1pko/jlFVvIIFwcaFcot97wFfABdd8JsF
yj3ashSbz8ZzK7LdLIEGo9nynxD3YiVK/cdujt7fRJ3n79Jm/+28MHw5mKHQMKAw
WvYsWHT+tnltg8x0FcwvnUnJVDMmXcYMJg8PSrv7kLh59HJExTql7TLu1n60l9WJ
klEEXIFPaOqOv+HHSlo4Gn+g2eRZhrCjm/UTDXVuj3E=
`protect END_PROTECTED
