`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7jzwlvoWQtY8UAYXZDWittSSSm8ZWjYz83Yw43JjlXezyZGVFvinutK0BkHTuT06
vKCCHF1XM/JTvXay6i5Uf/NisPrp4FTGFYPVrgBryIY83gbZwXe6CYb3n7xOvH1D
WXc7w8CHYgdmn0xgIGjArTdGsK1MWSNygMwwUwytszDbqss09LlULmfiWcEKtBxi
v8vcDErtwpySA+5k/oEyIaqgSUjaJqHXEyIO7MWab5UodnKQ1CeapFpzwVjM8CYf
SzQoz5MjyIb8uSBpVQpNGNnabSLniFQRhIiAZ3cEWYR3KVckD4UZbdPwVucKlO1j
dGkfusQzc/2PHTdqFILb93gwptZZzv5PsNM343PENyi03IltxmfLo4Fomv37qLNq
OlVXKlu0oxat/a8bsPkoEWFi2t7WzO+RgMFeXWdUiVhs7v5n6A/cgFF2f8CM7j1b
Ce40kBoIyu/neoOlO8YTW67DIy2VpYppH/pmcX8rEZfU2UttS/0YWy0p8rUhaW5g
gdC91/+Q5gGlpLMhX4zqcwil3wTs2cxaLeiwPgKCv3C96MXhSDL7QhYQqCbNWc+p
drgV0IjU0yXJ9VbIeLqOC4BulWoMitWNTTLN84ehnE9WazHwOPKn1Mn5iJ1LeOrp
5CsIX9ZSTC1vTDLnP4EveTj7HcfkbjhKMUHXCdBhIQHucuxqgP2Z+LnA/ufNLXRp
9jV1B6tA7ZU7BKJ+9ZbuxfJa8ne0T66BtlpR8O5jfUDQPsHxxwJR1NynBB6sedIj
bu9kyOm5jisk5H9Dg9nqocfaPePKNyFIoNAWhHAc30WXFZqrK9Ntpy+c0o9gQXY0
CDuyWMWshAIlWF+v4Iz1JyWHMYlqg4XnKfd8fAJU/KLR9LA+EwwDPb/8cg+nTjym
U2fuqlflS5PJZtg7LAQbWMWubXZ2+q/VI5jhi0mO73NwBOcVYfExRsNLCBwGcsbt
KQRbGtpLdAMyEl0jXgly+7EasvZqSlddDGgJq2URcnlySuWbjPu3CxDY/i+EVTM4
Z1lMqaBrAp7IpswxHKEgZo7gMNQ5EP6uvMkJ4Hbcz6zpnyZmdacQ0qOLbZCDYYYv
Vhhwd6ruS52fSRQjEdjUqoScT0mMS94FAhZQ3VOe3jabnVMIdveK89rXYuvXQzYV
/Yqbj50wtHujHI4TeLbi7VaulLxvH/Qo7B7BEsxsnfHGcMS83w0rBYzs/bLgdscS
rcAnzIOmN1KDeVVftEpwREBe0k3YVlBamFb04Q6iW5QQSTfM2heK0ekTOkyPeWny
mY2iEutnOog7vXQJeWK0NfT7ICLJURdLGxdGXsSsrpzU1p1n1cCXCczpib72H9kq
Y8cuw2BZglC08meYdMpukBNKOpIYssRGtGexJDXEwSLA/gS/cDQutm2lcFDACYzS
Fu5DBQy2nCRwFkzmkEy1V0cqwDiHgT3wATAd6cqKW/e9sbRmP5EhN4/esZin5VwC
XnmoBVrPs/TI5pjc/Qkrc1AA8wC5YAZeubB3ECCqq+hM2gZxgRRXs/dtRmXJ5/gH
lXzmbvZVwFQMp83XyNOrsUBzcVONJy4jy84q58RgFZv31wQNa0Cc2JccRUY1RteY
6BXNCfkXJUhT4CozQwF/XIonZXAaRZ6bGRPqZ1Kp4G5OWZJbsBmhSrKfsJZsoiNB
AnosvO7MTdpH/ung5VWMx9gWBLi3nBO+tuGT6yy38t32XbteuOtNq7kVOEkNl6IO
3nW3w6DorVsxarpEcVQ2V1/jXChu5kn/Zx6Swtmxvw/eRxHVBk2QUI6An8+0e5Mv
lmjLRObDacMtDvNxnOuSAJGkTw+Fo+jYQaHkk7ZSIBt0hNEEGkDQQ1eXMITX9zgl
`protect END_PROTECTED
