`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iF3zU2lqTe5ddwlQAgZoAvynWTXy+985uRq4i0mRLOlTJxX9HfnU4X008ETcc3Z/
S9U9CNTnyxavVr4hbAJ6kPgL1Kv0wU0nli3dRfgn8oMEhX1xcnu/ODHUkR9BMHOF
e0Gi1t8Db6fQTWbujDZL6Wt8BbCjmuF1m2tdYztpw+omkqNtnH1ARFn/p7tFRXFu
N3korbjtV6EmNuRRcdYJaUZF8YmaljeLOc4qf3oce3MiG/AIJvfVhFYB1AF8lEAb
lRL2q6iAHtJU+72YYA405BUuqLJK65aeG1CoRHAZFu6O7lChn9gfC44rVJQNxsIt
sYfl5FclTY9xH/n9C54ri6NwRoaH6MUaKQQN/8Lx6yng6yR00eicCDPmzb8nCLNG
tblhh3hmjkqkZJpEE1zihijOVIJGkNU2u8HAdQcp9hM=
`protect END_PROTECTED
