`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PvFS0KaUF9Kmab9bLf2WcauAJgaOD1z+v2IelnRqLIfHj8ruZeuxNdcwUXgxwmkx
nqh/S4O3kuhcLa2mBr2X1CUOWWiyTs5TL92pOc8ZUk7YqQ9GwUNJhetcQKU6YeR1
+VeBZhL8ILmX3Zq1YLFrXE1vx5VjpuArK+vKUuKid1OSJSFtKgM+ycAugvAeD4+S
9MsJil1sJ6J5dLvuf7KM4Qa1/5tMFLLEoN3RcVB+Mx9zcPXybmDThlUs7kIceNFq
lmxRHLk2btQHepnSIZRelNM2GCmUa/n5V62amyNVvXv96Kyye15LEl2j0QbSrexP
wTc+l9BFLpAWgvskLPNT9W0Xg5PdPiUqxFBtQPNB/fdXeRpbTLiPhn27xeei7fDY
qvy3qikUqQ0df4PwDZ8/Tj4KWy3tA4MzetsN+DEfdX5QnyiPPIa4evNEPfMihfob
YlS9+2y8xaIYsjb2FmqBmIDac+TY/wmUAVv99+w9DvzYaLOTeoPoL2riTf4br3X0
/+E2hUOLVMvgW0LUviuC9vibW2eWQqSW2DfNatkM9FgPS5I2WEdc2wfUT/GdBXUo
gbmOqr/hYIoiHzKReD7X+cvi3xoctxR/ccJZvcL0inOSq/GoUCdFFe5KSaOkuq+E
ZhtYZ4OqQS/GhKjtxiWoQ9mwW3PjrYGEMU03LJY7LsYjLa3/aj0D18CN9RpewEcM
9FjuQvDrh/sPb94Ey559xnvPZ64iKtAAs/NtQWLXq9ZtDmRYPZO+uMpDphnI9kXG
pVxQ6FwwD5syDRgzSV70/jTf2Sv65AwWT/Rk39R9KZsbaMNvdzL/74dOynHTR2f4
FYYlCDdmbnpNJpUSIqsCrJzLlv/gn8QNlw6mw8bj2DODljywta7FXbhJqQrAX4eH
V13wCKCdt/dp6fuDzVknynOv70YBgQ7XjXre53bgz9Zk+I5u32mD7Rt2YKzMBOYY
nFy/88dF6XoDvEwNl4YnqxEnddnQ9JprTu94ExD4JtUdwxPc+l67ORl5Q/RjfDBd
eQ/ik5AC+MgHjvRJrB17+dGr2rvXRCCouIo+rLz4OKuG/EFBcxVfDcQVNMDxv5f/
u6DETdDHDrm7S8PAnC7nyE+7eDIdaalk/zEj3DbK0QDrSF4gJL4mJhfTcOIhHFbt
L9V5hOzrDf9J7eNll3xk/svzsiQeDkbMXiPc1Um/uOAnHca+yEZtQREyhOgcnEC1
LdkIkr1uIAi9ECG7OcPmcT+7o7I5VIRGvzBLOlJERrRyoYZnjmngMUSDNrLukcoK
lF+UgxM8zJCFneLzvSO74FfzG/Xr9+ezi2VCjhZ49Yax8/NPRWn36T4DnzsrDcT7
LjfF0ol9kR4z/s0kroT461cOWGn+lNavW5BykLIPxBo1xvEMkd+Bjz4dJos/e4WF
+D4gN5aljjGPJRAwgsOzxzNZ86OEbi5dqajV8xgFcTEYKt/G1bPwC/LHpQorpPx4
o4kW0bt/uc6exI/DaSBBaA==
`protect END_PROTECTED
