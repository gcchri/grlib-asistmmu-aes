`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nBE4bbwN11yde+8dJci3TC5pXED8qsF3PlH6kguUziVKpw3ZEg+AqVe7HGF3eBSb
piA/HH19cYH7Qf+J5xbBFCSJvrYAO0/iZ9VgzokWiZLBGpIB2PWJY3pTB5FiiW9J
IJK36qiDQWVmMrLjVe6ZsVkC9bp7P89RodrCoc/RLhdBPFm+cgOxzuUdU40VnWil
Qk9yCvCPklPinmupwnTX2qaIUpm6xGB/c78W4p7w65JNRDDe/n8f4YDpFqT2MAwy
43dds9a3puhLmIWUd8hOl+qHLdOMBjXl+DOUKdhsrhv6QV5is8f9951OAVC8fA/Q
HSH7jKJ8Uh1SSfBuY+gTmQVENpRm4DQYNqBK86y5w8YbEX4cDHNmBQHGMX3SyIMQ
xUygsAKTECbsyu14Lb9SzcEs2omgvCHxSevLLyfWCn4/ApA1FMOr2gC/CetXIKdv
wC84MGfC22Mm1rDAf3ow2SZ8D58ol2lNcyU+vlZKzH0pA2HUmq2x1fy9pKlv+W9+
`protect END_PROTECTED
