`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uJD1E5rA5KDf53fmiX/E8yEj4M5/u1Aa1vnshEhrsjrjS2NF+sDuuPLIweb3Fe94
4+n40Dd1WHengmESJ+PzuBkEZomnqPIH9zI3GKjWJKWma+c5aJSNGQjdOWJh5ZsQ
/YZCFIMkCS3325n4afl6UteYKMSpjxGXyq8o8BrmfnDRuJWfz6u9dP+BdYHscsUb
RE4RaLrlRqPYpukBtySoAM3fD41z/kKYI2oRV6iaJFsfwC8ytNmXiYkaaqaNPeqz
`protect END_PROTECTED
