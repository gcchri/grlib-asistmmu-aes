`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ouiAsy8H6bSDS85mqWMoqPRiSkIlSwqUPl+pqyp0YWvYhxJOZ0+/9mWtXjrXdKO1
FL0e6KmIC2GiDkK+vued5rQ7K9ZHi0nWUECfp3N+lIOYr+45L8mWU9JkFBvUoR4j
Su8WyqTJG2B80Ov7t3UJsCMf4v1vMJwp/s+MbCnzPgXf1xoP+A8Ye0jdefKIR1T8
3POLPE9y2x/1fWT7M8WGNREgM2XVbVAabMJjTT2iK2eyNjBAvnYONbmQa13LX+7c
dUlnFt3VHV1/gfOorixB7yZt/v2RuqcSgpmit+183ibdb+tKMGT3SgvrQZNwgAEa
BKRcK20Fa01Byr3d9MpWzQO8sFtBrxtg4XQZq42yHbPorjkgE7tUzhNSQGOOfshl
LITy2rDs5FAtFJUKHG1KAAfoyGsQtixeRGIZYowY/aFQaZw09VVRfBB7GnAfQs0k
i5KTmmJNrFdJA93EBQBGEPm84sIdAy+9PjmODEUcf40778r4Mwi5jXmGJcpGMQY0
MH+vitxKixXnwTsZXIU02gwKXQFO+jjvwQLXzqqOQBrfNHNbhRMtxBySXdJDL7lG
XSJlWhoXdDBh0QuKndB5EBMxNoKOWovKV5He+TVfY/yN0GHmmPjlb2k3xk08bneG
j7bGQ44TvM7rH2LOT0KMmnKQl95Kknc7K2N3J8pkFzQa+HueLv2dO4NRQByyhgA0
E5BRDFLm6OaxmR/TyaFadSDmm0hr+yJWYHUZ3sI8FGwow1lItLCKnBosfAddAraZ
QQT/2lp5YTD4pUfrl7Fpyif5vG1gszyOZX/BBnImkOTAnp8exX4gE12N6/TSsjx+
hOELa3cgzD7PEMHbUOsYvunhdHD13jGwwgFR0Q9FTQEaRd/l+OELOanJOfUg5Ifb
+bGheVY9ahYaJrcwcSJMiUBsk6m5BtuY0xriT+H0HqhJZTT3PSnn2WVzJeavXOVa
hoH5RckRVY+wuUw9WoKS5i1g2zRO94IohCAZnlgDAmeszuPtivbToVkQJzOJHqID
I2xgyTPMH/TGnnJ3dt3b3JJwoUiY1WqLl2tg6JO4grOvxdZOVWrfinfoFI3rQSxc
v8qbX/qs3fqXw8HgFugt46guxntMMl750j0NQGbSH40rv2vwRmJ0xxsbaXnKIj7Q
llYu0WC3kI7xJEiCXhTEG08T41OTbB1ObRKoq4bFPED7zIw171ZFd+U4KT0TH5Xu
0aP9GtubZFonf0UMKwrSVLS/boL9KpmScrrsynOTGwtO6sjWiqVse5ebXaaQ0ZIT
2OAHWZZI+gnVGnROtIubNC7pYXagvslLxUUXhhIedNP8Z0Vu/zsOx87Xhu42orVs
1rDL6byvvkZhZ3zjAEXzRlaLqinNp9mZxwrvEJoUTCED7rinSnWFWXgdkw8j1v3Q
dd5MsOCa18+rZtjFBioEpVDUJQ6uzsjwG5bbUa8Ffn2nCXUqYQUnpYBcnPBZOMEc
V3E3LQO7cH9p2k6Ztm16atzoC5S2SWqgYKCZBNl9al67SKLz7FQqMDrFoxXQXAKA
IGehUeqt+FgIgMlsnfp+WCAezwEe01gTYLhvYQvBuK2lcvm7htbHBJiA06ax+2V2
3vcRHh6OkFWPg/D5J5KDv9AW8+d6S4fuQ7jsgFnhIWzu0vlYSw2LU2QbcWyzrLE1
R2UmkF6EFKsSyvGn7lxzjSuHtdGMl8nVt3+IuQsnWuwWSiclI0xGOoiASJJBstQE
MOvMWr8bgVnbkE60psT4pK/x+2JRAq8XwSLrN05+eMAYNsw7peAHAqnGWxpCofcu
6OzByADtTPNsR5NY8KOi8hx2BlmhpP/4r/BrKWiIBaNQge7qHWQM4s4OrqWa6J1z
26Fa7Q3IvJvIqxnDiFFJo9sQ0EcmYaFL6G8lXuzXy4MLpmkM6/ZskUEmFOBhOe5x
Ey3y03czA2b9AsgI7IQn921bRgq+tFfJf1LziLAkBWSowRKumfpis7CrxXOTk4RC
mteetShUz0Sd5qox4yH7TNTl3RNeQSWTJZX3lW8diLlaBK9qG2OCjjfuiqZfNG0P
O8ybfT2ld6sFre6a3VwptWHbkXQerQh7chpDQ209M56nikho6b16Mfz89Zgvgy1k
8iA8HT4KoIY+QTknpVrjR4bcXCqNAAIjvd7v1dJ/tIzI6KYANi+IWdc1VKBTXMkB
NwKlcdq0vP0J03v9/TRcnMJNPWKeU7nIwnB9L1jzYGnQSllfOac4lb5O68LD/V6R
ngeHgRl/U+mwBI+VGIqeqBZ80UDSf3H4KZOGN/Zo8a5Z8bmIFF+gHMCDnYRhftY8
5epzEbzt2eEfoMblRUjCHoF/fEEbxhtIhQo3gpFnxFaNuY38C38rbIjy+aq9LiCA
TMa5vGzaoXXzV+X1PiAiMlyVT98gyxvBd79z91DVDqoeGUdulOiQLSkhtan8DV42
HEH59erKJrHHXAdCC+R3td9Wlneud/8pCNZei2VvCxt3Z0VfZzse1+6eCPHI275B
JWTKRfi2nn9SrL6HCtVNs4kALekK9SEKRfncIL0mL5D/3UqfI32idOJ5RS9DB5TY
S72mo27xUUD7rChc1V/UGOfeP+NJRtqweypWuTDjTF1Oc/dJU89jLxrQc6X9EfnS
CV+b9rT4DUSF6nS3saxb+dhZ4DraRiDJLNdpBNVsOimFMPjiyVMs7cM65erug5Zo
s1kLcuqflL4Y29kXAsU7KsVT+bVHwqrWKTI0v4UWX/Ol2BhjtJ6uVOLcJStf257t
CjJCvy2EvQw0mVq4EIb1B2ZFlzO4eK3lXXwzDJnRqhhwiZQS0RiKoSiz2eyhusHU
50zPnQRvNJEXUNje5RX+uGWOBEf5EAwPnJh+heuArXEf6dSTWLx67Eq1kZwhwBm7
2LEm5iFqb/0q6mW7owy9YYsbf+kUsGBmGTQmx/TuwLz2KVY3UyFGMbsbyQJ6VSoR
YUFPYG4yy2hDPp3ytvUek7FO6+MqlYP7k43CIWaJaexcn2NHtG0P76efuIrR5WjE
O/UHQB92taeTXzaZmx6wlks0FKxD+PXYIRp8/jj8OOguLBfR2yv12wzXr9mBKikD
bRpE0350npjWdgV1loiywGtrzEahXxysM9Kv/ooYsCyLIzpAqQutfvIRLjwUoncd
FQ/8Zeah3FEg9xPpgECjcCY3B51FVrBkQQsU2ofzrxilT4A2sEeC00I9liaY/rgJ
o2gDmkxTO++LzhP0q3pULpPvKxpgW8iQS97JA3zPIkwjT8TmiYsbjWKQURO8xRNZ
thQTcYdp1srGa88+LAEIjDLZRkTe1ojBVpy7rihiQwtkdfUeLooRIjXrv3PJCMPT
WMa4aG83Cz0ToTLKq+mJjylM/BNWqBJ8qq5c3bxZzRgqgZdkCWALD+4JiF2pTfDi
99mCjnEr0agYnxMIYSu0nu8BAsGdQdfZ2Y8kzLrMHa+/Oo8fifKsYtCAeFHUmyav
2770HPVBl8kV3jsaLxmwuNRDrdl3zJz8g7W7QSw9x6pO68xM3NtXibUpkSwmc3f1
ih1tsIs5giZQZD7n/dqlWIJN+gWSpM3cUNCRVNdNRh668YWHJ0YVwB2n8JuHo2ql
bYm4J11gp0WV08Q5aykBuu3M1yYBASUhZSgrMTGDk5UaZMBnR1MK1wUWjSWwWfah
S8O8EM8fQL9ej++57G8L90ag5sBxIc3Gcv2Yyztym9Z1RP1UBxbubwPOOme4V1Zv
0atpw13CSw6z5uIpocgdzF0VL4dKRsUujQtDdTbp4Nnk+IxJSjhDps+v01NXoj1Y
YKgZk/eKjVVDQiH9f2CEk2EmSPkSZX9KavH24I57WEcXKYwmvF3KTfar0warlnKR
4JBFsvaoN1txFeayEzGul03MPqSknDTyepyWuuqwAJUFrzTtQETp9kwRInDufEwh
IKIVkvDoKuoh75KHAEruHMecWUxUEV6VEKvLwKYagMH3IHPKdX1SAjsKcAWYiM4F
1/+cHxCBmxSt0epfdAqD9NaAUvFN/pIHfwvtxFoIm0+WJLctWg3FMc09IfoYXQgy
fHRVp7dFfUTKymX5ZYJWJo0H/4arXSzMAVUdBBSZ+AkTfXVivtLlhOkEQlpqF0jz
C2q/URaTkC3HDCEtTAnLWJqs38fnLB0ktnWj6obp5MG+zb6VlEjpXbKJZtbO6EgW
ge2ShAJc954W8KQZ0Ov8NQNL9Bb0kS42KJCAajDfhJ7GtAAwYUFond+fFAIOb8Yp
eeAKVMZXsCaLUTH4nk+Emggv8mmjST6nmMz8IJYYgsfJuLd9A+DrZmk6ZJzRraGl
xWYsH46DnFrTMzJm83ilD9dypHdwCE9kxbDYXoIg49CZMfy9l/+wk8pJMFjR8AlW
zViTWJYoTkFCi/EexRq3Mc5xDSc4QBdR9or7loQ5WgH4lxyB0TBJc48kAyvKL6ly
UnAkGfOwiPgjsa3mxhPxHBoZlHrVTZhUYn3hVi5P9weSlISnJ2l+2ic0jBEYkg1J
3h/GWVfN9VWizJ9SvvHq0AvryLo6R2GYy5a74OP76xCGU9t6UOpH5hcWdbMLdazG
533vwbTzSa0UAoS58k0l523puMG0NdbqdBetcGIO4sUbT6aMTJEabP4kr8DlfYRN
gGbxVxjOzVQD3f8lSEMzBKSXAi2JUFQRJsw2aiVK0crSrE5qdPyofDQSNi9sstgC
Fi5p67D9KzDekiMF5LEQi52pzJiu6NQf0JTDF9/fJLvZVYjZdLfEPuVSykIPaUSK
hI/PlASc7O2regQM2+/bRsT3RUcOlFz0nMSSS+Tp/QVXQsvGj4MWhof9p8fVEgIt
v4u2z2m6DkPglxijMWIYo+KBim3kB/rbwzVLNLf2w9CyCrDES9DHXXR1WUSsKW4Q
yxf6Me9P7G7BW04qFwA4AlMgqDdiyVkpT+E7wbrt8k9VbCk6768Wl50AAjbIaP00
8AnGEurF7fgB5dUhE3gxhyx3dFTr5lZqwXDlpGRFysRpaGOxsuYqcJB7Vu/KinmL
dNpF9sbqsf1KoicyE3KZy4Ffi/mcIP1lt7Ei6y3Ljn80XZX/3amsYFHhCm+HJDat
eGccQUqgZUBBye1vFFxmy6yGgelQYNHVBxw+rO6kZLwpi2HtCp1zTBg85K8/Qvpl
9GBP6tx55LLrPmCSjkBcjIGNLqdMXLKuwKNSLlNeN3+LFpiWDERAGYmYdSET3ERD
pBiTNyxzB0DQvgaq22B8gcrjvi9QI1GEMSsVey68B64xeJJqUcwWV0GnY5B4dsU5
VLe6bkd6XAg8pGrAKv8WV4uJcYVGPlEPG/nMSapzVj0nFYlYQv2kg9HSP3EnoJ9r
/00ESDGPgTv2Ra/H/3ehqCPTrVSb+u/VVtE1ywe0++/ntPcM6xk04z3l9eO9TQyl
Tzv1cUi/t8bVVjl+/U488OtmL+Wi/gnD4WF56jxHPUWkXmoIimQMhA6iTjK55So6
3d4kwhqB7eBxfC+jrMInAbkeuDs22aYOnOClV9FjRfVStu4UNthCcSHdAd+VjaEm
Fh+8vGExkMeTPIYDjV1dFOwNRsPZur9M7KktwdKlZRz/pacTIPbu+xbysHuO3YcO
8TK3YgKX2SWsbAQvNg438cPvP9hv9mhRv7tk2UH50CXG6tXrt3+Viphr8iQBBxFC
3mRW0gK6X/RMAOrD8FOquJjgGMvWuI3hHmZ9oRA8GGFd4DOlmks+7J+4OYCKyUTJ
xg4qz3vuNzHSONshsikgeqCE7eY11ejEhx+0AudSRaQWCXOdokC8y8+qtjdUqpTE
0uZaO0WLBCFSmY4OIBKN1y3MJkHsypVfwVJW9mvmh5UHInwKwk2EpDMZ6oYechCk
wQwvc0ImEbFb5I+UuhmkIKOfVrxovQIwt7Xdp1KEMAp+N0Y2Q8PFhE0oPqKgX4wr
je5k65codyYQqjq6f9FXJc1PsYwRKMXl8HyHwapupbFT+CU9JYdme3z8Aq0ani6R
gdrTdusVlxeZNYve7hFyIMIKqlNRUS9m3Jd/THhdhjovZxAYdB+Q5wXdw4Rb6WCY
ckIaX1UmZb8VDU32CCL1CSBjZfmMiTz5xHDU4fp3zSyjrwx8pqY0O9usy64Tthot
Pxd3z/7hk0ieVurxlPpDQnBpLrAFjMQjZfXQlKmbCfSPPrIVPcFrMwSZbIfVIkbj
MKhu4e8m8HYoW6Htu83ZNgkdX3szUCRmRFtxTM9PvjLRNqwbZrz748DQ9APgFAmS
+z/jUjOh5k+TuCl0LUmSd+4tBc+n8YPR4i5RWx88NsGHvqD+oKMV79qCTwDLt4yb
d+h2aC3/dLMrjTJBzv0j243CCMgrp8aiK/Il1AR18bA1gt50koHzfFaQ7Y0TYvGX
eo1Ixr6VLbwhmr3alT7fy5GDBHfZdBg4c7ErhrqbImPe/B0ZR01pPVeWUePYq3c3
2q+CEirrlrItMcuHM38HDuNkvWnS/9/qOmkP7ZNvZSTAEvTVQnPfPqKsxr23L6lV
9camEeItmFD7D9X4tXXxJIvC1D5pPq2xva8Z38V83DFeK+uR1ktATtAMBHnGP9NF
UFssZdYszI9j2bKk8F7U3xmOXja/DOTZ8jWlBEFwqmCjCZFyWwiMtwa1eBb8WcRK
V8cVgx6ge+qezj9pj/FVgR5Uewau9DabMaLEqklOR9HdhYGAHXtbaGtfc42rBMF5
FgzmLfxPfyZJa1Ix5H38AP4gdaQOrPS2ySjCMrilJyYp/HskmT3HtFsQVDD9lSCE
5BEr1Uz/HHQRL/gf/uvRHqC/eAe5ee6DTTm0Pi26X88JuyhUAf+HJWRgMUyC/D4C
qEA11hoR3C60k5g0tf56kGNgSa4oGks+YkL4HZQXYLHpVS6pJWQQ3fmnvQtoDCkl
6GiN+cPMyPSqCu2sIBoPYpWlQSRP77vk7yVbkw23SpOTJBHSRgSkNmGxk1uvxvYq
pYQEGm9hxP/cA2XcxrdrQLuyxvN8BpPz66NzrFB6rkbeBL03+EKEcs35Ti3jkXIu
eB6l+zhSs6PSPc7+aPXTtgUe1Wnj1Sz+j9DzeXvs7sDhgOcSHdbcgAkttdauMg/+
HaHv882f6FDYq6+7x912hbayNU+YMMudSXFP/6CKlD8jXmyXFDvXa40bJ5S9+sDL
gMAawJnBr8czT4VhxhT1TNsNHBGiwCugcDl1T+Ih0NRQI2g5DTu1VOMn4rzXpsGZ
Rf7SPclMctmhwdms4qjDVMZlIRbiq3tALLPXCNp8g5sZXoI1hpRNROTnBD+T9V25
7ljp55hTyWCZk7spc4M6XIpRAGI1sJ/X2jLmlzffFVjZsQtqfvkPM2BQN90KhLjp
6STjQYiUYvjYKzWCoybzyWcZ3KH+GG8dRBPlFRiZljbdXP9Ygs02RkZhPQh4LTOe
XuZov5GhBEGjHrDl28QgF6Xk2vk9A+HgrgzqsAh9EgnmnaOmvmFrODcnd56c6yyH
qjGUcsRPqd9X6mkhIS9p6z40OSnvxEdY/0T8JCVHXKxaBE/Oplr17uehCI6g9MFx
Zf/tJ9SxeABJMqqWENtGjZLj1A0DaoKgZEmu5/3Q578sDNk1HEbz9zOBsSyPjZw2
2RSkFS17d//wmrlSOX3S4GLe6QtjaLAA1i3szRjQXI4By12p0EBvgidB42y6zXt9
OoBkCFXEWv9F22J0UFC/fL92cWJwFdSyCUIKbrq3qCMtovwWu99HtwaHjsT8k2cG
d2X2JQZll78svf72tcTa5P+fNrMiEdLQUesPTx8HzYYTnjXMqsOEpANWIv1ITF5I
xluF8jUryw8HqHSrXt2M/qYWAuw4UE/atcnhkcZprYFmQncUJsCxXBwP3fzE3Oj9
OFE+rhSRexVnoRihZFA7tmer3YgmvZ3/CQVWrppgJ/LmcCfRN6P5lv9Z/r2+gm7d
3SA6o9OXlQeb2PSOixzgBdkfmv8SqoZ0wTROWoc7TM9KKkc+NIC2I17xQZL75huU
Cpk3zvR1f+HpKsdBHleYv5GBZuTbzqXQlcb9QmJXRS5mIq/yjF7Yu5Xg2G0c/CGn
HW2OY0vEhy4po0iXpzAUG4fyMCYmKlX7DEly9jn2ZpNm2+V2qM0HsOuNY046tFiX
3kx2VilHB5iKNwGc54OltSnMmmgohHZELuC8qYhFQWga6BDS5Dib+PNe3eqoeCK4
L9mvqx1nWDvAH0ul2RNhyOsdS4HOQOffgx4U3F+E1CPJQ//9GEh0Zqx0IS34XHRe
YtzRpgf6Wy/FPGt7vCxb7kOTifEp3IJR2CVxmGe4zViRqPdmwknCabeJCi05P2GI
RPCEjxddzA1kC69cLDchbZIrxNHdo7p+kcoUgI+hnqEEJXfhlrFWzECoFoOCd+61
wS9V9uCGv7MWvbGyrPIeZpRT0JJbwFH9sHpZCEOj/a6VAHjbTyFs7ZStlWcZPZUr
UPamOQNyxIXC1unXsBCDP0k8joSjj4QoJ3Q/2H0VsD7pGY2xsvCXeaqIy5WNPFmY
sqaIhhwQMDAYPRSmGTEHGck+bi1Izc+032xH2SGthZ/5qbXmAxBoN5cgrzGMO3Hb
fjXdHCJm/JnFnJ0JsHlLEuCxl3TS5A944sUh8b7J7AGh67iLESzXSN/fqeh07a5T
Xcjqk4A7fpbqSGyRWZiM4s3xYYSVR80UPiyGgunUA8fZGEyFj1tW1lv9rcYaOPFf
KAQgDMMQUOhTeA/49Vu8F0nzqEDXaG7p3y8QvUtO8x7gqUI7z49GWyHivATglOmJ
gRG+UNEKq5Gw/h7koWXPPR4Jx62A0IhkQRUesFVxGB1oCcrSuxytXLXA1is/TsHD
gldyhuFsb9yxovijYWessn9mI6Mr+toySy7Gf4vpigdWitEKNyd5f8rw5WWDr/z1
sD1z3a5C6Q6dF+jP6NtXJ2MgQF1aseCHehHr2Yp/W2LJZveLPSd+dHlCENiljql+
iNOVzOThDF9gFefM+8EHxFpDupbhfcbsUk5CicE7vCSRXBoRfwmvUuL1lafRp7bz
SG3Q2wnZgHlDGVpqIgSL/cN36D5NE3doctLXrecaUAo18GM6X9ieSDjJLuTr645q
wQ0uEJKNDn98+V81hPaTPyHt9YbndGX9LNggD67hipTOYsUk/M2ox6H8K8UdkBp+
Wb+9cckUaYLGIWJAaPlgw3AYBK/1ArP0AENH/Itlp0jdahwM38EZiaxAOlYeZYTs
XMAnHO4tdNr0mTERpfEFG3izCbHXsdmuGsocO4Lt4BmgSMJtWZgqW1OBT1aikIRD
ZZzn1BECPL2VHxil7bnt/RRwpfM+DHHZYn7ocOGMPxnhLW34EOxzvK8KekB0pUJW
ONZv5aZV6hlj6QnC9JGfeByjYbmJpvs8KIK3HEbv9UvlYE4g0lTCmHd35yj9USVs
UYLooudcfPTnWOe2aSHf6ZIXfiGu7P9Bc15jmsQdNEhvT9iIuN3s0MqNvhJxWZFX
I3oPmdP7tR6hBYGPZe+ErqIChEhcKX2MzUBxx8pPN8iCeQ+R3VZJmWq5vT6vznbw
q2U2Bwkr3rcbi959D+w2riDeCuUFnjTa6F0JSAUvyvm/015MpkNv5jV9vVQGhirH
Z66atSQ7NRFOqEQ1INyNfsl7rBlybx75aExoDruwcJMGHJVI/sgPCaSMpu/94UDr
hx9jCh8Wqe8K9zZAEmtTmJNmwQqoN8Ni0Ak28xcf7Zd6F+mnaJKgmHS9RqePoNtL
S1/FhRDl6Go9QUo1iHsAuCm+Tyy46Qizz+givYI7ED5tZrOY2K/sEgXqHmPF4BHE
VSlI4VbZ0jOQqEC2S4HmJ9tcDolL6w/vCOFSGZkBI1hOezw4jajCQGSX6QnI0l1a
MvD/R/DclSOoYgQiw9AubD6YyKCprchO0D5MYjYhIkx6BNxlUjQ1Y4HkxM1POx4z
dYXUtbO/fSjcqYhPmZAITnApuX7W90vAPk0Dn2CxprXk86eZoG6GP5dZSJHsJ7VH
iNCcRrtuyjDfw0NIh/NL6k0VaTtV6GCL1ElZgeYXnGdnIj8CHK/WXGQCf7B/LeQQ
DpjpnSDuSfOoSQ79xzSVudioleggzbKkIY4FtoHtJnNL6TnNz25Cf0VQn7jRVbKM
XtDpg6o1PjF1FjjbDJ8JI2Y0vzbxbZ72D5+vXtVqIX0YyDK58TTRrj5lOhJqhONw
Kz+wOOhCfLfht11XYfUvMKtBqaYEmPh/u08ugz4wlY0z0jBX3ki/3tWy10UKLTi/
dJ5FFCuqxAawZY0Y0uZmsOxEsO0Y2qQdrt943mqYktCps9W7THL8cN2ivPCd2CFn
qlo9ii+VUy3UneoJyFwnTiNyPFr7VX8DjRGuW+LJILwfxY2Xz9F7yu2SBEQoZD85
8cjnopXK97OpX+EMf7ArgAO+2UAXdDIDhwfZoX85Md4/fbCLOcVq9TGFgnxmpqgr
nrygmdQuU7mcMPBCIHjmAD8gZWMgr/Bva9giOciMLMxXi/LJIawHy/UBEa54CmHM
XyxgOKr8UdlKIpDkX7SagZBChfQjpKAlJhzHb2u/aXhLV6dx6LTv2ivgR6u/yKeG
G91sfggoWoxL8Ex1zVWvkQ==
`protect END_PROTECTED
