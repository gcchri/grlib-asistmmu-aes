`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EGVvW/x1OtwwOvO53M44q9qErwvIhhR2Fskg2yFKzbkMreBdWnO8wn8n8HwYFzkT
Btrs7u/oBWNTlVWCeXnZfCWNipMn6L1TueV0t9mrndJBa3rxXCXqjzuzwsEyJ1G7
uilpEYIB9S5sEt00Nofl7msM5EhS8Q8JxIefuO15FccOgFe7WPvvJTzBlmGqh2Wr
iGOGuvXWE4MK7wmkP0p+ndsY3jq6OaGygxaK2904GoJb+QmFBPsaw27Bjs1xi2qE
GC07R4Tk+4TPQ5PhF3wgu1vL8OHloXrTIYqG+KS2ha+rBliewJdcDWQK6ylQh/WK
tBeUXZVumGZrSDYcApORGtCdhbSRRvj+/GHU5fD3/wk/ENDzN4Ys4u+QTpaKb2zX
iRDJS7isvJgWgb/d638VuIba9ZgA3g2UvUvL7bAdOoc6FwXGUcaZx63EpMfqWHtj
2e5jBVkvMutArGcFeHabWOV2/dnfryzbHeogEK9cc0kq4FjwMlKb541v+hj3A/cg
Xx9wQdlX4CCqbHIdmYfuWVfOmeFDeLvcVfUT7/53YySy3S2+pClFh51VB5XxGYZv
KbcWYdV1D2YyBoqI5/Z1d8S7ZY2h0zoPvA+afcElfbTxt79EqwzDuki4+1edh48o
+qHBmTZnxWF/ZHWIfRkeawNlhYlRiZL2zMSGC96w8v5KRcA/NgUZVZiUMZBi6ytd
f8GPAcf1guVUCQtijwUPr/LQqg4l8GUtcKRUvJI5GrtosJ0f6TPFqwIW77VHPtiQ
oukch+uGPRc/YgVM8xn5j/PNLKaFitWE0km4Sh2liYBVkiYqJcKOupwuOmaJ0w7u
iULXozTkjHwjIrNBycoTXxrCcjBJ/GVXJmUZhuTTt2qZCsYcS/gdib+05844mFeu
jtIs74G8vsDcPYeC4irINb8MnJYCH3taRJdlbxS1H6b2bKF/t7YSlkWIgCtdPGuP
EVALLbNVi0Bc0cp9B77MxWfxxys8Jyemyh60/idMNcX4Ncax8ljKpN//pWnw8mlo
q0AodIcIQZJMU0tJnBBieYT3sUSPuayAH/cjO1zbUnlNaQjCOWPtt3S/eKeRxE0v
w1Lr4wD6KbwH/d4CIRzacCKsD4DkO58qxlgoM/vi+Gg=
`protect END_PROTECTED
