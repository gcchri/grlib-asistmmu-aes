`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qt0XvQovf+8Cu2Izfb6Pv4jVqPeZmAtojd6mK0Oa29NdY5MsmM5jIvJZTGv17qi9
l1VODkyjAhC+RRv/mX8B7L9vFg9dUY3gx5mXq0wOZRI80iIcL3QOwHYiW4E3z3jA
yBITVHGzVE1cVjGHa9XVKgdDJnkv1LOqo9k0yELdQRLp/RXcONea3LYB+YrpxvRs
F9Cs4BcA081tGGb97wsKjX/oKytxeeVu+fsXrQ6PAY41yGuPKas7VJ4t9Gkixd7G
XTJKjDWZx8T8jTn++Ei0kBZ8tJ5yY6W+38uRd6RgiI92bnr1U5lkqh29TW6k77kw
bkOWrVyM+m4DBQP4uR1VSBIpWSEI0G64EN16Na+wfZ6uKEZ3HY/dajawJH3kLPWt
jECAjtUmGNlOTnGaLOU3JMbNgy+ywYaqI0BKprU0RblPAdNSfcxLE4Yb3/CYqZom
d5cfOcXcgwg9phi1jUnVGHennDAq7qtDrpslZ20817vdsjNAaanQcas24ShLL7sM
tcrI9DIzb1mdg7iwaeYhZNmxYlIJ5MC2ccgOeHkIuZNg44ZPMV9nUhV4+0KyEFU9
Mtp7nsHsj3U56ToUy9gybzKw60JCUPO/oPnzENZ0u7i3IMyApV7Tiwf2bmafVXcr
erQy96BEQi417PnpXvjj1dNOKf2vaKv/IVPejZctOtueS2F9B8Q7SPkwcBZAQz8Q
ug7GegIduL4JBDNTeFgoHiq9+3DOa3yYnrqQPGkDEyjliN38mnLrx/LSUVFO2Kvv
h+qPNq/KrOHxJ2R9ZKyhsJY6JohfhpBQF2H1w9k4cjBtmfIWTrJTngCjc8/VCQX9
wDukzQBkQ+QVQNTR4J1w2AORHaTCMRFnNfeJu46/xM1O7dJePvU7WpYyNVJMMrDq
wX0Xmxh9Y+QjE2Qf6DJxE+OhPGsrjgAzM1OoE6k+BTa2vf33mrmofi63+wjLV53o
R+JhbNrjzplyQedi9WKrzSg2TiX+3428PJZCA63zWJzV/MgvxzfmqrNOtkdnhhf3
f/Z45sVgAjHi/oI3UJobia3cA1NlRmaSWRiWY1Rbp4xM2tLXr29VcGn4PjQlZtQ3
V1CWntzib2NljrZt6qnWI4rqRffEOWPO6swYUUiTnmsxwaGFoGJ2Oe8aJnmK2g0V
hLHgAnvjKMhrgfvT8TmsLdZ6joZhhVsc3IE0GJGyW8cvfZvKFCJniCAsDCVgerxJ
m/Sii89CP3uqZLC021yrMzO1eaEyq5zd9Tu47akxtmiy44vKVuGmjmtRJtyWcli9
IayT7zKQpBU9ibf+nJtiivghaAOLcsyQUPOB6dwaUwtJ/xB0LLdVtvaMwxo2lrWW
Q3PUieUJiOBnAgn+qTEP2p0OtNJpfmfKaD6dHp5ZnsM2Y5w9XUrWZiZDiROA7e8e
xsjcjs1rujbtHKAvCsV/lbfV09ZyBarIuhCMPwMWhC39fvwX8SnPdsR3GmsX6OJI
9RjuWrA/w7ropOa/g0Lxp1Y1DweNG4hehXgVfOjrToPuPLeVQU3w9+g2L20M23AD
BIyFSjm6klmmaUH4weVdwCYwqVaD1g7429rsIRsj0lymR+pDOqLyUK8SKUOKNbrA
30gxOmY2sjZRA2Rcgml9tX5PwuBfFaWxwtWCvLG0Ys/A4ee0R3rhzV09pbDwdSMA
9eVT+gdhdVW5JUKVoiw/kTctxJG/qngy/PFD8m29D3XHRDvdiNV2RFF3LSwquPJE
OX/DE/ZbXGZufF1CytUkXAkQ/+feCiCRAKNayjxYFSP6x9j2Wc7R1+SDQYprekzg
3XTvrhsYDOuxNToG/8YCirMh6iw6H2EeLyKsNWHCBsa99ZPrjw8YWkiPkOemUB0w
`protect END_PROTECTED
