`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UhUVCMvZqUvJKx2vp/uniIa004c+CtS/Wz/zQusKiKhOOYUI3FroE60y4/o334lw
sQ0QCLH94xuai5a69r74IhlZ8So9j5O65TnEJqRK7sbWZsAJ0jWidPq2c4m06L1n
NgD8dg3KAeLaoBzEUMaABamsKj0nqeCewjmyzNYVc4jiyN4rJO5Y0pyEjclj9bR7
inaP16UzV+59YKmzurEwYiChO0rQ2BA4XEh1F4dUXWCxlcN1A0i7luG+6F4jhimj
XCcs/8Sk1ecu5UhP4CziTIhrTAyCUIqAmpkFZx+9uu0u9YFs4FXJoZUaY9Q+I2nN
L218FsmyhRUP8wJm3iXvLBcQsXD7MZ0ZGkGDtfegt61wdrqVRFqQ0Jhz460jn9/M
cy5snX9oEQXOVeAK2Em2TOM60Qtl80bsloA9kpcR7Bn+nu8Bs/Iu1JnD26QC9EBv
BemlI9HtxyeYxFiOpt8ybeLgUr4INkCHpKM1ibHXFrtAhCiCLVmTuRDxDJhyoAk0
Ov97aCyxkLK8iHu/zZGdnhLO5JosYB4YfXNgesT4cebwiN/oEO8ZKkt2Ke51Nj91
AnYYyGElTjCyjU6q58BRm1Qokj7aHiFRXejsSKqRvIyOKtPZyuTGLvJt2056ghKk
d/VOiP2YpRvArQ+UBelwtbWSBf9bBgDPuRYOlIpKCa/oQHE1vNNMh1obz9vKbkQY
GPQyVuZxfk5l8aCju+ura9d8DY3bwqZL9EdRLWr5a6sVNkQ7wJAI1cU0GFyGcmNR
lnliztnWcGiTv/7Iqz2wwJE2dDusO+7L0nTKtD/bBZCrT4UfXjaHWh9RUfaJ5QLD
DU8jVpxvB6yxEXAn8PsjRqnLxE2vKugxoOp4eST6u9wW7iTbVESlVdxNvZPAELRy
2j9l45vOLwd8VtDDRgSzGi8WltT+Xj/6Y1ToOf1u6uZx/1oNkcNizi6KuYtU3YWO
UA76I1UtAflkv+y4e0u5VTtqqsx1Up+tibMcYit5PIlgv21qLaYxeP5sllUcFxFQ
0Md0DVZSiRC+Bw1DM8PlKiJv5FWhZTWUu1MDEeObHpTbwFJmX8eUJjGaOhEzwjT7
RdCzUcDS0GjnuEZpUqqcE5nGL/pNH9To+3ruTFPVJESZoTYVuruEXhqhwJk1KHI1
IItRgF07iAjKIDdb9OAjTScwv4oKyU0/hA2mL8OG9CUpM/iaFIwJ97ZwPA4/hyDN
vkeIywtYJEl7eu3I5Je3sd3rMJ+19r7mhWnb5d/H4l5ANGwUrgfAOEfimv/5UAwa
yll+Da82xlvE29smpY0iMJhUI2vE31//XZB+bIljZvMX3ZPcjLtqEqwsgCxypiPN
Wc4Stk9E192guyIGb91aGXjQY1geOdSYJeSryQvU8LMCUr9uNc07vPKLxQDcR/n+
8Jg6HqY+e6OCdb6MRnd9scX5UA2tPjBob3Q7GM0vUzEhPU/c5JV9emtNrUQtnMQt
AQSkNZBuwgwD884Kv6VYf3kEUOetqrr3gtCErmHMLqJpTJiwmWbjrMn1rM1Skoxk
ljnEYw+rjNz4Qt5VwZdftuvkAJgWrFT+1wkTc9eyucQTvJxELsqGeF4/Lqe/MS0n
v3B2AlE0MGbiz5JhOasoRrBKdC9Gmqe26vxAADiFo7RJqNFo/nhwUrYX6S/D4xNA
kd3DnRdna+SJJ92g67aGi8avFwhDWyArjxjKIjUqWLhCBjp2Twq38si+koBaUaw5
u3irzTLqeHdodh1tV7SWRIVrpTVOk5Uz3cTRNS90MqwHF8PArHhXHxQanor+3s84
PneSHJFLljWwxFUfjpuNm7PRsWfLLmeShv8LhUhATr+y3eqPUG19O3o0i3gvrkXQ
hh9Nrdc81qANvQDO5hOGF5LPDkDKv/Y8VBKgl/rXv1UVEGGUFlxlYAjidDb9JoKM
dGUDRFVU/ikdAaM8603Yd1CE1QLwJzPweu2iseyW+j8maKMWcCF35sUaJkDXRA/O
ktX7IeZ2tNPJ7HGt6+aI3ZPsVgd1GwZZdAeBSMc10IQUM7GbXp+OBCOQhcVKeR6A
ewlUsKt4WgQTBCsj0fHfPZdXtOu4qETsKXi15PSG34XajxvoDKV5EDI0Wse9MKa6
JD8w6L+dflEzlSaGh55y4kbSlZhcDXrLTPdyyk+YGmvOT+syYUdlbd4eFbkQtKyY
pFVdAYJxj+ht63TJvtTHma8o4laS5ElXdp5/CB+ZxAfbegIa0fM9+R8WQUV0SwcN
apYKKXcI0P2tpEqu7e4HQ3JJ4gc6dwgtPqL90my8euwzpG+3AuGHommQe+LkHHpz
iZzy9krwgpI65WI/9G14NdBMI3Q7R03OkhutxmvsTxzbBszu9AqitBz3x1B11Bnf
yXhi5OnjdpXB3DX00DXW+gwupi+Gnasb0xek5zNxnk3qJW6WKVSe8pgLqhoIe4mE
b7JasKWstoQypxPkplp0Wa7dw7HA1oy3Lre1XEJTYC6oUm4cqeTg6eytApRDEGZg
+f2L/rYCG+EGRk2hFvbx6Nx3ii9CxaHIlpB2lcyFR6FPsd17TOW6um0Efr7DzCoy
2akN/yIazMScZZZ71GQ63y7EfVcq6cwrtQiuBK9Y3B/84Yna3DFNzlNj+tw1vA6s
JHKTBnZjiJvfmtFrJbw0nlUSRB2EI+BuRocxhNZOXjxMBlFBrLjhzOiBI0PSkfx7
XG+IX91ubLhI/8+Rc6lTbTL8jq4UjO43NYCfQ2x2bIDCB1WJ1aaX9OkDg/7BsDsK
XNcWeOnDDYVM+zNGWHscFeljJAvPcYgkggFfqjNdb96wKxoG5/GM7GS+garxnBqt
lWu/mFr/qWvCRrEXo9fcb94LWvpan4rJTiOoD0ydQUI8n8xLejYL+3am5vrO9MTB
xPxacko+Uj0bPR2ky+fGLcphvU9SN0YUoyAC/6NI5O8+nl/JeMhUJkfcSMGv+zsK
OZxt4xD3Z9hy3H11E77HuqX0jNrcOXZ9TfxIpQnITUckJxd4bT6d6K9KolErEABQ
ilMPwTGM+mXjWORom1YpDu5YrCGSGiAP2F7OgqDH4AIvo524+aSQPkG3DkppZEzp
1nZsPlNGXkNbt2q+0UrXPypHaGDrNpS9FKdvUwdHtSK6m3Q+dUsz8BPeeFmXKUAP
QGuRO2ddA2b4VBsQ5SuCdi4gKNUzN0TWAk68+7cJTb++SCJ5oRrjRiFiqPeSJB23
BNGvo4BmFtTutdip0G7YSQcZTRl8lSCyFf1OnnYIYGiI8gZB1v13ueucOv+Umj1+
s/VcHSwb1vvrAdNuHHjFd7fR57+CfFwkE2VN1Zsz6OlE5QsNxvX/F7BZKRuI0bGJ
w6uGJIRvkpz+GCesbR9KQO5W4s//vwHjzvjOKpnKqwc7gA26GoXiNbl51XC3HW6j
NgDh3a62+ilPHYr8XEGEE0RMkC3JN6zS7M02iUSlQHr5D3hmnSFs7ukaHBmLnHGj
6amQVIex/pIEsPLmYpqS+goFgWwn9mxDcgoYayVRaLGVf8IUepoJSDx0DTsqMzow
XIOyVenV2A8NjSgLJ+8+/Qb8YaA4YvnRWh7EFpGnWi7kZYTrHodoZalN4g7NmY0W
xioz7oNYeRQ/xwvzIA13ygs2ONuAKowKHIyJ5WKWid9zKw/rurTNnPw+k2eYxRby
i17rDvBACigqx0djTBufNriKYn4Mo7IzTGzMTbeJIwf0IZAclowJiL89ReGVsWAE
/Q82O8ytxCT0gSw8msIPx+Hk3JEC1Dl+H2vCwue5uX5OZSFRwbsUCX7XvL8cMjLx
E3P/VkQMen7fdP/p7b16Uk+HkLLRlTB/s/PekhWR34S6+6Opcjt0sToeWafu2HEH
gwfrZY+0A3vuuRBDY8zc8djk8D08i9l0EiQPCPkiDFiIO1l6dj0TNgj83OS3B7Ay
eNyciDpmy0ZaCxndBT+nvKCgXyZz7yw3pQXBqN6r3MD1yt9Py+HkEmR7cKiBWCWP
PN9YKtrmwMnaa7aT2utEs8cmzPh1sFyVg5oP/oB2I0pYtEiMYLkGjBG5BYI9wCfE
mvqytF/GYEdUNz80A+Zc4CRmq8wahxI4fHjRx7NUUIPWeCV56FQqKgOoXDGdb2uC
S+qiW8q8lwiUclLUOz2NM9OR2GvCGznNo5FqLT+3s9eLjrZmmdXA24hG/JbY/zhn
OwLVqlTST9OQs6BdDxrEFkF8cBjwzAoIKkuhPFi1Nm4F70TIPEnPVHw8Pc/nfWbI
VEEqktwhsetCJoY6eCwQb6FYHvQJYLqdyzcvXX/U0hVvpLyvxeN9Tx3Zlgnj7omA
s7j9oWVcgQpNhJfCaCiNr7iDAVPxRnl+7jAO0RyF+elqNXbm/kV1cHHClets7/XO
LcmQLgLqvAaLvRv8eREBwjwAgO1AjRCaT9Y9w6U7eBYuVEAIKi4FJUJd5hZKfbAP
KfypXgoMMyS35uVCCvXPG4z9Cm51Rw023mBfOTzJIrabfUO6NTz9/OI8lQvheED+
v9jKlKELcF4iu1ZrOLB5rvnOZqRJeEh+ayfP+PYDGMCSBVnt1ZbCZpU+1l0+uMbx
AaRsLdBIhYWm3hlHz4Y9TaY7k9bfNZFFA+LBUeFE6DoCPWFgRXr9COj6GI+hht16
7dC0gbR3ujquqTAfKGTG5ev9nlqc/uPoFsaYS746AVpvnUtGIQHipkTxJ7XBtKKU
hZfF5LeX4IfG0JpWIxFF1RTQG7zGwtA6vRUiZjJgIO2ENOMOqey0NWzeDrI7rs2C
OUMZvneGql08N+HsYvdSSMqBBp8fOcdoub/tnOJZaPRPOGF1vBHu9H5e1djEtWxS
fR0C9g5HFnjPg1dbMrXZsThEWFzMPcMJnXvZaFg8eIgcyhWPEL+kWH5o5/HJFd89
nE7MYWLcXfcT/+DMQiNQ7i3MBsnin2aenOxuC3mtMX9DsPhcBbH6kWXn8wxgYkKu
eQNLa9CZvXlKQHBYzn5bzFKo4nWKDyFVHOzKFH3mRPD5HScBVyPJU8CgKpdjQSQo
y2tWt13oB9RGLS29XYghTVXmqpRTYgPwPwdBp69ezagB9XAct2jFSvgVifMoeLIl
dXWr0u5BAA3d4uH/sDmkofnzMRRtxSJpRYfpR21p3LA1AIbSKxI+TKmDApYEu3uj
6n7YSCoc+OcAs+xD1Uahd60ElP2LDrVEsFTl8Saj764DR0zh+dgzfhUVMRafW1pK
0KrXJiOV+coR2ehSMaJI3GpFdFAvsPBMXmkvmnGW07ov4ccjSiW4ttTMeIhdQRYe
0mmgf3ZtdZ6ZRENLACsmp8sB76ljpjDRYx6vlL9JzR2c8F/xZFOOTRNHZGrZ3TJL
kISkbtWxJq3gD2646Za9n3v1JFS6ly5krZogl/Kbct+nWGIPtVRxR5W/MDCwLnRL
HgHyp1br11O/Fpe7QgswbyCzbjun7Bv274NrNRiT3OgeikQezEeGf+z1ZthwzpsS
+OoqPCrz1nukvRli1nHnkag5zWvliMbkBnmySvMCPPmo9j3ZeBWaQIBejajOFfve
zurMR1dP4ZvPTMzaKjCqUTo3hZ7zKs0vP0FhkSa56+qkOySRvW1t7S2omixuY6gO
Qz5QX+WuffKjIWhllGE4uwFldFgTlDAf1ugEfk5MNLEeCwfGSnpvmcKXL+AZtfaW
Bxfb58Tk2P5CWjlhulGI9/MpdUSRCZPeWjyxNGthfzr+i8mCn82lz/Zj9kQkbSA7
M5P7xtryuzmmzwdUP4axzZckDj/gjmZEQyxAP+nj7A//i5WxezFLce5MrFbnj60F
WkIptHyWvKWf+HzbsciHqds7VTzYnJ0Rt3UKPDNjvGnFUhNhlaqKemsHzba8Hr0m
hWJyY7y+bb6fXc7ODwM2uhw/jpbbg5tuXH+zXEs6T1XI0XBiDmeo1HZUE8Km9fZn
TQLO+8NgirYMPkq8Bo/wPZWvsU6BA0xo4KdvxZPozQXV08JFLZoxREW3VePKdCAp
H/0LvomRUoeQqZHcsvcMSCOLkHDP6RS+kqidUw6M2PFfKWgMWTzfPjnwm2wiulWv
PDzHUTV9gBBYTqVW1M2o49C5htW/2fGCuF4DOcSONaXSHLpkX7K9pEg2YjFitjTk
QhUsroIJIA7UGuniIT83YvslEtQHTJ1WJRFPAtXfWCX+Xuep1Mz77DcZa2OCDEG4
Pf/61BVLdwsnTb1/V/jUlWG1KnKE8BXiMDWuYwruojvhkn2ZHHHViBlHrJouynnN
cNQAEXIJttydnGxs6Jj6bRY2HojR6G5+9weHOC8rOIy/Htyb/RTNJofjRbA3MqgN
y2XhA05io3OJ61nvJQGC5sX7nUIU1d3WCHv4yiu4KRco+XpWvOp5H75fS+Kqbibi
cr4oaXGHrkXmThpzcLIncsQUBYVOvqIjOklWFOufiHntP3UBQ4Upki9W7Pz4GvTy
JN7m34qVeRWE6cfGO81GNEBJlnFZ0m2xj5ROy67j0VxnB5GH+hrzx/vpQ14G4k7N
Jhv6xt1qxgzuwybjmD0nI9ISt1eSNuuczhvtiiRrSdXyW/yu1Fy4D1fAjo+y6oZI
rLVOuq2Wx0nFmTmKNtkoiX8dRvFE7JhkN4d966dYaDOYTYVRIqNpcnxkwF3pdjbt
upIl6xQkmHpX9FfH2n0B96MRYsIF8JbyY4ka4bLoS0ZI8P45syRRJUNXALQT+Z0T
o7T3LLWbKzVtMP/chYcIg4/ve9TwTdkCsChzRSsX/SRzkNufK+oDHejT1t2loyJC
4cRt2+rTcMBp2pCqL3GUJ9glK9ph+kwspNxmV5mHpLopbxHBYpbSovgtNNopx1ds
5OxEqOfsr8DbBVZo3hxQJvxQ/qEufNQvLr7ug40OOpN7++LPhu0J4PGydEiqdPjv
AzST0SBs8Ta3/fiCSFrzyZqf7Ay370HS7cYLAQ1xVlejzPp5uk9Lz7rPBW9B7A3s
EyjRJFJg9Ahehf49EWiLt9epqAGb3lU1obcLuZVRs9IwyVcwJaKvFWwG35FN7bDZ
If1hiRiHaAl4BaBv4v8n4elfbmSmjF1a01zj6qu04X3Rd1d3SAVF0Q6YWH49nSEN
pv4roT7wok33R5X3Ynq1/vlF7MMKYJdpBOaX9DdELk/VbXnpwEIN2qM8DuKDpyVO
XL8GOIZEw+AMpI3jYS/4LWigIwMWpRpcsp629oM6nbT8Z9JX3iU1Y7/8l0D1YNyF
AhEOklRtMRFnjbLDUtG91YwX1WDC6HE4OW+iZLPjLqrnzO1mQHrynNJYmHLGsI4G
tO8IR0Oxna8QQHMWRW93WcJ1gcowpfdGx+ms/MMZNEBdoNdfu5n0ptzMxDFZIpzg
yaUjEE3Kq7zvvZLOxFL9Tjv9yW9qFJYrjfhNsuqyUqv1PW4UE9bPczPXyl//SbFm
7aoZWtgTL9G050vqoLAoNrX9dG5OvRcCDOCYKimWaCmEriKezJyscvpIZvimvRfx
rzvy7XZd/zdNGiddRNorQ+UN+mlOsU6jYglzNBfY8ryO4o7+QE5bXTbbBH3aGY99
ZLQZz1xcA2Pyj7K6EaCcZ2SyKUVNQRQZB78/y3nN/o5EnUcYtnnvNKTHUFkoIcEE
V+OqmKD4/roBOM0u5G+xrj7Wd4xqfKbnedpTGT3t29mTJTgD0vU2amBoWmC2SIuU
z5ZoqBQads/k611KJ7pw42KLvgSyo4IsLm32b4XWVypO/F5rmqPVkK2X2Ac5fSj1
dB8HXHFqkjWJt/qWkx7IenazdZvhxPb3qXsIKk6GNdgw+ieUrY4z3voEoiKmgW8c
KQDeIEDcFp1yzJB4Io4RDn8crt+DDzM508vjOnwbuGrGKC/XBhbcd/TFxKzWy9MB
6wnE6BLJ8Ct1s4iTaab9QqIEkqeaboZ7g8P3Zszjw39+ziQSeOMzqjwA2xw1IR8X
Wr+Se46ajFk/YsTjAKfmx+/+v8ZWmrU60fpDIse7vrrcEsohx8Gv8FjZa5P+hNUS
0wJ05JZo7ZMjOuhFg0zo8caAiOn4oEdNqVHVe6R1C+LInRccUP2mOkp7kibErZjj
0L1YtHzQWl4Ea6pRPszVDK2OYd6SUVnfwzLW8XVXpX04wEvwSEvp0G/JvTrgQS/C
iFrFdRrqx/gN9XcVYykfLXbC3a3E4HaTu7lHeFpbRDnvl5J6qUbsiYk8oBLIho+z
6LIllbK0RJurjqSaxt8C6di1qpzm0Jy3tZHIKmrbuvo4y9Q0KH05ouh/yHT0WiBX
nEx44RWQYeu+xLsPwZBadMeS+zDpSOUZcE0LQGzPL1OR2/mNK9vgaABMNlAi0n9T
wQaFCIq9L8oGDLn/HDirhAMqdR81j7m7F7e1TCe4SylGCtZm1s/wV0QkrjIb95QL
XS1dr2WjBM7ANuQ+QB4Gfiy+24Kdiw/2UQmsLzAPk+3rGS49zXhIEKhsMMNKcI8W
8+a/lWRB5UmdovpWjjxGJVjRdE/qVBwJH8+kRMS4GCQgZF46wEbK/VFAUkq8bY9J
vcRazmafHZ4kCqwr65YDuYkafe1bXMDDanSZT7bqGkIbp4qIAeaILLxjZdoyPW8G
RE+XiWaWz3zw+cYkQeUuuHNPyBjT3sZLMj15oy6jborHF+LYnhcPzml88vADeGRH
23xcf1Vz73p3exmjQ5Yil5Phm8fBRbCVyBCWUGN9s8IotfGQPwAMzgBPENfRC0S9
GzBTjOPXDGuuXnfTXHRVEYimkDzLWtjmTLumMzPIOKKDlW6ezw4TrOc6JoWwslV3
/ddgh1wBzmWKn6zROuZqJRHpgUlco5RZW5eKwmwh/tO2Z7uyu1F+ykmbiZZniSrA
olJwVfo2rA86J+1O2vFKoHt0CVVT5a5SQLukjQriI4jaQBoEg9JMYuODKACVQM3j
yfPHAeVIoJlVtA0V82e8lClOcZ6JD6zgmRdT29OIZEmZCJ1LRlR4fPCMANgKfohv
mF811WxdXQpPgqCE1zOLGm7vMjt1yDYO8jGnhnAysWBO3Fngtkp8E8TZg8gT/ioY
CxezwHcGow31Pj+LS+c3jSlMM4Eyebuzxe5kx4zcuCV15XMEdMOajr9TFQpW/t/t
YUqrb0VNQsP5D3QDfzW8Y3CNRgFU8ay19S2wfuSIT+wBtIoNEuto4RTjU0MN6LoG
vdhTKwaJ6zkfvfdRZQRi7f/xXNuqwQL6C/20wVyCpYJijQw4wcbKsgQfTuxDN8kQ
FuwN81mdg3AGQrFTnrTLmy7IVxWvVaTjnuKwcdpTclZ4jr9G6ORrWinYS/ZjeGHm
DKrIfqK6cDp9w0mTmaFrJ3iTgMrRq1j0OCUJwLC6WOee3ACIDywbh1gWrQlIM371
2+WGwaSI8Fxwpka3i7iIQBA8Z1NpB4bP+q9otew/6aqj2WJ2V/XG/HCygwSdmJBk
0kI5F6qBx2kgwwLxTClgiWFbj9IfWM6avwdSJFSbMgEAktCWXZ+55vWSfKwIdslD
NrjouiAannc/ft5ZLfh2HhukMTvHAx0iwoOnyY/eQapSPSaB3ognjh+Y6pv7TpPh
n2Og2lS8HiQIjrXWqXYDwxLnpv9NlOCP9SCTJGeFbUygFSvAbsSGZor1mhMujxuT
9O10uaI+H4QjfrFEQzDlm1imtaHAfnfrHwpuPeedJMfXrNknswr40x5MffyEtPNF
0xm7lCKX1OyaSLCZZfcHeo//2GYN+Jzu+vqxk4Qfg++zZj0LV9tomqpoTwlyDYIT
AKpDfrxakOHM30I3CNvSMgtjIiRqS408q01u94gBRug8zF+4EXOboLBBt50br5R7
kqGAl7p5Da4nlZzmdmOoF7EWX6xfH4f6bsRxtNNgi173xSVBSSWHatZc0O3lY1ys
8wZgt1L3ybupQ+0c5QNsQ5pzxMY4fhJfT3qUhHdWM2SOeEZLec8ZWmcjrVPR6wwc
dznQVw93lQ52cUAMHxqW0ZRZFn8LeleTsWm9t91GdjJQEAfny5XLzemaYK2U4duz
Q0uEmxkmiePlX8/Px7dDW7z4TCuP3Nnxw0aGQHjysrnl+8RMo6E6EQBJtLuwUc36
xJpmBNKAds5sNofPRuLSJTmA5npWaAb7WLvLjdOQsKOnedNzGIAHhWFlQkhBRAcx
0DYSGIYix61pLevWJ8fRvhEfe02qbGtTZz2ERNk8MPwnxDzCBGGoI5sMAHqmLnrA
yrdI//kkyCIekkK6iVkFocRycbaVqAovz5N1jVeOTSHCFRzS/uQHGEWKD0H7A0o+
VlOD5a84knisfMycXc32dYx8JQ1Bz8Luibtc+1+6y1LlVPXSO9sbTViA9orzXSNq
8WZ3pijxZrjZt2/yxht3b3Ej1h3+WujDXixAGXV+IVT1qS0uYnh2xRYdHuOMxDFg
EqqdHS7+b3TQY03D7J0eTao58TQANCa4NQSDvY6zoiVsrynQMziIi1vJtyE57JuJ
W5rfvs4XzjegOjtH/VMY4377QUoZRGC/QXMk54xMrx5lZA15MZkOqxWdCpxZvw2v
SNpJvfQDk7XtigQtK8Sa755P+FIm35PoBdNRUIr3VOtS/SZcJYWlWoVgF7Vukt6w
cnBenJjRnw1QT4PkqJ6ntG+nBwLfrNPZVs3DkO+I304kYi7SWHsrDYfchISQ42Ib
j3Mnky+y8wwGFYjr1a+v97wE5eGbtYoRH3wL60fuj8LJgqA0Bu3YwOY3n9QY24Jc
771yJBGUhhQymuT8wJX1OB2+y5ZXuwnPj8KzmOggQs/+iH+m+1cF+5r2kdwjZYQ+
Z87qCbNcXFzrDFkl0GX0gkfGxQCLtPlJd3Z2yxZP795qoRl2VXNU03TiB74L8mq0
hyUUc24kR5VclPB9uMhcYQhnA4IxUg9Q2OlG1WGx275RDULKC1kebttmjVdCJNO0
xO1G1SCrmfUE5O5MCAHGgGk7Y3UJEbKBbBrrYqyRks4sN4nPDl/sPm7CGMh1+0ZM
vKMfFEcRs9LyQ3c4UrimX1vqz1pUs779Ve1xSxsW77g0OpuiMOEHPb+ZWVviRGIf
1Ih927lrqq0AgWYJ8H7Qeurh80r6WuCkEf99/StEoH85nzT2aIN3E4sa/kN5FGMi
bB0R4H4V4xrkcV9QQNxdKt8iCCOZJvkuZZPu8Jdy6Mu/JqxEsvK+u8Ac/ZSI2vPl
MsaLs+hfhobyleu4NnD54jp9Y0waK+33CpnL7tCMFutr9AKeSZc/3k/+124Soral
RqkswNekr2DeWb/Bgl8ZO0PYlger9qy5hMYvFYdf0ysLYh+h6APzxGC9K+WFbzon
DXi2bBZgmK+POOtIRs5fpmsoWT6aj3ApoBu4uB8K2o3+GqNwXmWCrb5ObqjVztxJ
4+W5Cu7osoBGd5IvMybhoeNa9BToiklozpivkpTZIR0HwooNlmUgfCe7QGbldVBB
Np7N9mO4RtZK19vsh2CbraADQzh7fZHWgQhZlWMAm+hXCv/D5r6up4VM6Rg8pfx/
na7FPcWnRDkXhfzJNyNakzpGZ6hNnqDdQNPXj3smGArGe5HpBifkb6UvjqR3mH6j
FzKCWyJNtI0zQhAFEZYkQT4HCBZ6zVX8N1irDlpaZWT3AYVAtT1mLQy9cAbQ526w
iujrMaNy3pw+cRwNX3Vw5qNE4Ps7UtDTv16jyPxWC6neQcZfJSnInbxK81HX/a6p
r9NnUvWeyc7mAtqcD6GqyeMhACtrvKcwHKMz9kjDLecj93E1/RyOmElJeWCdbRYI
cwLhlyhGocGNYNO5jn8ZP1tkSz7hRJBzsxxzr011HWeK/qGnoipBkGdFrmgWtA9x
gornTEUl3VPFdtLPRqqNfn5AbbRVeppjLO6/Dpz7C+gy5zZu4p8orJChldO7+Vdp
aN00agqqGS74fYoNRvrua3Tm77vhSps8H5esTCPpFg4wpgZh0x9jMjY83UebuG/+
K/SPRxhiA9Xe71XUsuVldZ+/LetZxKcjnLPz7uXxdyKm2EkcTMLdrJUlttIRtrUn
RA+gidFsk9TepqrDrzNTDrnJKX2NuI5tEiBRP7VR4hxsy8hm1sKsE0Ogm4ChTjGI
ll5eZ5fFwdnCkxBgfJXzgC3tVBIfKUwvI/2WH/m18oiLYecOVe1I290RU965Nk3x
raJ9Qa+zgI3sET1GFNLZUrZ1NXBax6Soe601PgUtwar5XG8pQHs4kjHRVAUDCzGZ
mih2fKFXtsrXFj1Axf4Ypfo+zHfrvBmPxommdOKMJZnxcu6BwtwOpxH28RO50pwT
dpq9QGOu4mY6En23OmAfwdcGQhbbsxVqfY6NxKnFFug0USV7NN9ByieJ8nic2IRL
sUOA2pNw2RmsVFDNdoIM2QQf2FnKmbAVeV7ma1JMwx45sEMGyolSthxt+XzkWSg2
ZcLxAHJn7Z7KnA8xas+SbCSTMYxjLU07YJmUFSI3od3CVt0wsphGfqr7VPMG2LUi
O8JV+n63IAoCxPG+i8S1EqW/nP0k9COirxpfhqmvGVrhxwxnPBkQnzRKzJv8HBCH
eCVRMCO4+b5ESVjiwkscBIHl/IgOv4MdeXiDaL5+Msr+x1ip/U+oKeL5kK3jHTIi
cXAPEGGHem4p1XjjYTG0aZmoEvsOtEkBizT53QOU6ybf39DB+Lg6e6gMnCZ5ts8b
Lr+Vtp1vmHEQi2Etl0C77bx4/6IfycP5jUqblACH+KRC6B1bOUZNz3DB4evYEgjR
/MC6mxqL4jAXNAu3gV/jSB4fFOvFrrHJr4raW0edGGEmLajln1ceB5umzn6ph67T
s/tXUdYg3l6hKGrM9exLRCf4Klr00FtAYqJddXqiED53nmYTRktiivOhLiBlP4bC
qsonYN+kYMUQRX4esQ4M3EqxESUAtyFOhq3ETWgUOSibp4EPNIu5JD4r6m8FAPoS
TIIUlr1pGgpAFm+iCta9F6OK2G5bhubhdRNe2U9+p9pRNQ71WGnus6UocnXnMHj1
5QnqBRqGV3vT7YPuT7TU6tyckid6q2C+zbVA+3eRKsRJIB1fciVgva26zWuHqWpK
BWzPl9yKJImLA9/qjBTMLkOKzInSsNeQmtBryCJrgTr1WODKnvj5+dc5Iuhn0K9o
OgyKJKRgMYLYkXVw92nVpG05gO0jBtfmGWN+iHv3vbchkpE2okokUeNRxm1kFfGL
vYuNjs3dIz6YYbz3FY6KiNoNSOaL+347k9FIzkuVe1Q9yZbjauVLcS0RqoKkw3rL
pOJ1LEywkw5WXQOUVxmbEkWnH4B3EJwnixmnXxjf1WNfmRP6de1gGy+tbJK/H7uS
h79Bkxzpa8pooH8bK4pKFKUXAvZ5fSJal66uwmcfShfG9XH71eg51q/FGaDSJwcK
QEIFgqvk/QgTQJhJk9mRrMOPInSqaktCkoK8ELYZwl50M/xJto0iwznagFL6ybR+
B0XtEuTs/+KCGrg9yXVUjHTimC+ChONaE2n38ePaUqX42inbZGBx3u9Tb9inZ5hi
0x+LPnr1zuqLjhzxhwVcq9aPtjsfxZsslMZkf7TnifKFSXQAc2IsQnebUv3FAlE0
y9UFlraCNwd37ztkb2SpcFbUlKTbX09T7fsqbLR0mZiuH3VOwbeaWkI6sm+kaeTt
DBkP4k3CybVYdRKRhSvE0enm4/XWTeZvn9HBPK1D1Io6ycVhn2koL5413FfS+D4o
8TAWAF6dU4sfPAtNdLdpHL4+LkYluUYK8f1y2D5FmvA3VszDFYzkDsldpnWH5yQs
iUyuA/BxuNN6ZqDih9CGazJVuK+Mo8zxtQFrdRlaPK+iXvyOuh8AkXi+5UXxxBEq
gERZaws5/noEv3rJdxg+xH39RtR9TCwn0+FK62re9UcNlSzqruEB8xAqSfG9TGBZ
gLee4q+JE65fnYgjVKSBV7+lTfEbgjFXFGG9eCfgaHFQoQLOc0ps5ibuLfOCQcGj
psgZ9hwYX55i77eC/677KwUgVgH8qT9Wwr4vP11hQQlLUqMkXeaAnAr8N7rq2A1F
LYiujxjomxJQuVByZZS/1RLXxsI1n0nsWVB5ajKDjaiHwqN4yHEIOATd+C3mh8HL
vL1eM5x7yFxw2mz8PiglDfE+Z+TtMwoWbqrk6007WPFqYT5Z7XnHqsL+k1yvoKo3
vR+gvnCKMqcJeH9n0eGy0p7nga1UMTYPR/1DljrnUDfMfUrI0agzzp5a+TTyd271
WuxhOX0brVFohq5R3iguzz1po0g/BKAC2p9Jtq9G1x8sedCOE3gjptahSH35lz1F
a6zjqvJC48TgKHzUMdpMUVJFDma0OvF3cmfmUH9seGecT+Jb+fXQ5fSTmzk8eixo
6vXNve3IxWU/TjcXvTQTLENuLVKm92at0GnQ6ocQlTmtcRTmxCa58/kj8mf/hpCt
io8tiDUY3wy9InjPs+hlW+m/Yk5MvP312GSPZyQdNMPi3UfTx1ZqjHyDP3JOr91B
PhNzZOQ0g9L9rWk3rIPJOZ6c12+LJvMAa25+LBd2vikuTBnGv4rIe963m9aCB6eV
nHTXR/5kQH1V+ydqcnnYU2Rs0icOIZJSla8F0RjkWbjZ9chJxWO9NANFPH3W6dfH
EiNx78Fe3SyC1Dsv57OOsM9V2P0XKe3Zvjdtm0FmMislq2JX538RqxjUOEs6ff41
O13BRE5oCydtlz0Xp3fpnSbSTtjcDP+Upy3XVj+L//wUz6vZ08+Wr+cY3BWNffc6
yWE2JWMlRb+vR8yZj4Z1RWOSvHQZL0J4iaNQPOISAgum0zteuppX/1qdfyrMJ7/r
6MYMr2EBeH1bOWwzmpJsWRzlucd/lmBojNlqgJY112l6U05om8UOqlmWtqRUy4sr
OICYMs9TAEcSnPKTtEp/BPvNKssQks8tJaKzzFqDS8CsU/BTQGhcfIJO5xoHYzA0
tWf+8nSjC/VvDZOYS68Ggej6S6khPL+sSUYBANgOIBqocPtWdQWPAX/7T7l4Xq63
em2CtvUGQsBkZ7upGBxbnlPsmZ+9KNaNRmhlNj3Gf5GWbND6ZHE7gaosx9Rv1apd
FuLK40oS88XR6iQbbfSBcTXpGNpy/ZUMXsGoEZzFkFsPOrf7KlMqIb+ykHEgZv//
BmCzm0O1RG7yX+/eV1iKmxue6wblSrvqPgnql9UNemdrHs6gj8lKsusOYfq1xMaC
sfA1tzgF4bGCUOgydk/ETchPX3KGaU4BGsKytbTPe6xJLYNy1pCZWbE8mB4pmf//
Qdw4lmoLtczu1aBoBjcWUv2w9ODdVFHRuqGmrBOltNhutsqmdrVs8yOSUsCo4P+M
I6/1XlyjjpypBebWnXF+DV+ehOKmvTe54ReYJlPBapNF+Ago8qxeaJoBvhOE0Url
WGntizeulMd2N0ot4EIgDPlr74TW2uSdKAZMsigfXu+rt9gVicWr7p5ML7JumsE/
nkMaWXMTvZkFrZj8r5oX0jCtaSF4F2dICz+mPUst9hhXViyd4wLWG+oBT+ounBzN
nGnqyNlgWtGn0aIQdvCVMw/G4XTKwpj17QpuZjsG1Rqf/ZGfZNBZfBqPLLKCgJZE
dUUjb2V9os+NwBXU3pILvMo4FvlpqBvNsotDG3qrEAIgFUaMCiuFonOKeQOXGF/D
eXmgsSRP3/6pRkhrvpXKEWTSqQeO/aZ9BBeq9plQx2Krj/Px/iZrGSgib5SAKWv+
v8utm0G91s3U74lBZV4F8XQ9Y8nMi8NuAHj/v+J4prcMYfrqu/PyEAFd5n9VOE6C
uQ99KqfwawcmKUw4UV/nq4q6xYzGMdPdybtj+fReVn19tjEKStLuA7v7hrtQ1zEQ
9EC7UyjmgfDPWvgp/oPMgm1XqwEif6iQP0BvRI2AudX3RlpmfglY3qHE//PTQROI
In+llzVX1zkZZlTAv8FEVr1KwTIJlTl8Wdf0yxvluHbCEv+0cnMm1I7oJqc+p0HN
JICLAh1Gz2hZCIwC3AgGYPEpr/ZxU5s/yKHLlHku9cMZ2/6LnwvCFRappKu8lVJ4
B7okFLQwMf+mNNkAEQfTZ/DOV3UMgKoCwDtrmCj+evXYUCf5H2EI3VgyoMkziizA
QJCn5s9ao5kIxG86DlirmNKuzuWFNcHK8aJTV68PzUbiSE0ujJDNfqpnVKjs+F5J
dg/trfyXreVMyrFY+Zzh7Izg9cE1VBCFysQAAmBfBNEpAfnETud6kLHTKr0ccH5D
y0HGj+meBgaG/0xKaJIKksD14P/KYiaAiET7p2pmuLaoQ3TZCXTfglUkvlXdTMb7
gKM6VeYUNeDlW1L+da3swTyIXqwF4AgZPPyyxab7JcU0vvdDo2C7Wj/Kxqa0Kowx
KXcWorv+3PBdV6sGEboG+SVu98Mg8JJyowyx6YR+PW0dwj7AolVbk7BimM4c4MFk
B+FirdXO/u63amVLU3fEZ5vir7/+cq1/YJS3pC9J9ShKie9Yf3k6Ctelbk1JqTKL
rLS4aoT1TKxjLWGcU1m58geAl0HkPQ/YMerW1Xhy4wcyPq3E2/fHivNMZLkLwVvu
JezAwZrDE+eqPhb3y3veTy8UaWAwKwkO0fOcDPIHxGp9qfTtSQBYuYHXBg+rtkYg
9tBRZvHAwxWjFRCDdzGweJXuxH5+6yqgo9ExEJGZNol0QYizxx2ze/7VLQUZ66UJ
2W+msDd3I+bAYc9mk3VwuUZGwc3S5yQP1jgqGExZczcJgFJnGNRvooSLZb+AlXIJ
1jKryN/hsr9McQu+stEDZfJUGiDJMwtLrIjOwlOnusbAURPHeIAsgNamtparY3By
DJzpVYGwowfp1P6QYrZlKTC1CcUzOO441OKAUIFuMC9jNysghiGakQ14n10zHzPf
BKQtIXPtmwXBnN4g9VUgoeplwDM3eaSqxMkwcqTaqd/WnLN+WXjekDW+sz2EeUSl
BVaiY5wh68cfa4rR26S7Y7ZB73CyRNnq51GydgMUEHHj/+T+DBW3HELh+UD7vp2j
2SX86u+PI6uWudq4ITTBxx6oqvvccPL5ZlnFhUg5E2Ajx9k4/xxhOdTe+TaKwPLW
y0jyTi/dQsWXgpVIfxmzCQ5BuGM+mxeUeyK8hepkf/4gefzo3/lOjfuk4AHYw6Jp
Xm4r7LLznvT2jWbz4gK2xUVPTTc1Q9cFF8DWBq7GN7++ByLmLWzMP9eCFlcNX8SU
TF7NXVUJQRb3Dmdoo1yucOmSBohnPK3rs4KLDZVkI/8J1zYF14cg98hNfklOSpp5
+G6L3SwTRNdCDNylBiiuvVldLgYJHvf+FCWYjgZ13OiEeE5ncs7ceRRQ7Sc65bF1
w0psGCSfyJgqqJ1aoOPO08B0Vv6GRdbZULl665fMJIo1ef/S20tZ74JOxJnfLR/4
NTnKQa4FFUntig90sYUA45DSJm6LtqrEHZfRHzQxyYndtQ3z31Bd23U9Yqgk6aZY
q1Uke5rFI5alkly+0ENjcVM9rqs1QifSvxyNy54gD+Ru86dPO1xur7stZKeY5kb1
gs3rH8mRIufVOHpbZhUZJf73h3qLpkE7L0zLQlZwT6DHlAII1ZUuYScPiwyfB6ur
MO/CmHWwD54EwnYmn1Rh1/2aCfk13Xb4xOu1OfdKH01r3VNdDBX8rUXWlov7Aol1
G8FaUJsQCyqKJNjrhmtjxfB81Ri0qEFe9SicZ8ibAm+mMCVdsgLk+0Wh2hQ0xzvf
WwPMiXHIkJgh3Nb1H+pG4GeNclRdHRw6T5hplLveYRMvqcFu5jgTpf36cmcpLupz
U2MIKH9NZsPQN8MrOqVakpF0F8sr4bhCaHgzvG6phgDzjORbidNxV8Wm9Isl/apd
Dmya6VBD4DrGeYRytrZh+uxrnJ51PmkUf+ZVyYCVlVrSYi+Cr7ruS2+CTlZexGO2
LoO83wf73Fj2p5YJ8oUtzbr0/oTueY+0wKwGLf2UD0E=
`protect END_PROTECTED
