`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tfeio9+6BV4DyJ0fwtt9E8Y2EU2NTK/LKkKYIWSzPCFDaRa5lq/QD7CmZQ3f8XeB
q928/6gIV6GqbmElnMwInXEeJ4KmplFQrd7ZX4d+n6813LM/lV4ZQ+yQbNL+mITn
JaKWQ6Y/nwUWfS5NaRBsQTXqosFKYYZFBwVnpDuyAnVBjEjOnao0kU7y4b6+EP3z
ABKDrwaXkwg0TDRWcQ8BbzTfOQ++jy6Tat+J064Wq8IlyJ/94PDpMep+IwNc9k7g
8hSi9mmrUf8iU/hyvbXoLOzaUSXXVi8o18CCpa9rXAOxLAaIY29LwjMmJqp+kUGw
oJ6QiCOk5rdnMc/D5qhLdM2JKhveGja4T8SZozupHjLnhpl7cxqfOfwDFo5aTdKO
JSEcy4oEoBImkdzagc/cLHd4KMIN1n8ACZJII9f/4awXqLu1bpGw1P82xIPQ1hv2
YRP+r2bZFoMxJZABfhv5skxo1PC3MVLGoHt1YOBrz55KCBcv5kUnQEbMtTTUkZX/
eXnJYzcge7vbzppe5QHftcnJea9Hil8bQUm5KXIbkpqdA0z54JcFXWQinju+GkJW
FByWi3ptkZSi46bPPQCAXT5z4EKau0krhbVQOEUtsmw=
`protect END_PROTECTED
