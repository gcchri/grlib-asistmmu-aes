`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BH3+GA2U/TIdkZ0M/HMeizltfdT30XrjsWGydaVvR9V++qFsCl5SVTh+3mIdiiOq
CJJfWxsKO9/7QGmHSckSZseWVXF03DVBFXqFhSbAaSb5JknD9VQla4nnc3ReZgTy
h2Y/qrOna/2v57zOQsqoAEoHLH2FuWnSC3P16sBikhR46li2+MEbnDKVFTzfVqNu
Mb+gneXZ0WpBlH/bt6DWp0rXf0lJSlc+o8yvdHjSDkuM62ffdiXvtCZXNfFtyFnO
61E4NbVpVHUUgMSJzHsLljv3dY7qKnEZeOF3BfT5+EWXmH+Co5gK6Gxpg3s/sR9w
XxEA7RGi+C/WcBCnDLXGQCPUnhGft3o/y/XGNXMb8w9j3+IQHv37du453g2m5HVl
6Jjoy7oRStHDUyIn1ZN465jcahCYUoQ+mB8/ob6t7TXOkO2CbQVUiif0YYFkw5B0
fzcTX9dcFVEKXXrh3bcMQg/5YGKnA9i0CQixQSEA34w=
`protect END_PROTECTED
