`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nM4JLPY2hJnQABhHxIUVv9zrV3mJCybo8gWyovulygQV5Kaz9G0Ts3MolNoyP6yG
1mewo9vO6updrJ0zVkbr2FDT/iQLQ6e2PSI9z5CU/0l+VKdpOHu/04sQNFTaYlGK
Ex1wG2Qx1+sfPwBQ5v6uCWf+Pl5nzKgVkKBs9Hn6raXeqg8i0kCGcD/laePhgM8h
SFJpyosrLhsCDIwFeg/YPwz2Rc9/szwgqW+xv8gUkP5qi0LbMWUJOigccD1i6Tph
i1VahKudSl28hlpK/P3+5A==
`protect END_PROTECTED
