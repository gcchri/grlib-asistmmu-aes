`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qBrCwvl+pvY/yvQ5NUAY2Q0foIneElT8BMYC2+bdGD6tnvpXhhWZ2hOrSBqUSC3n
bDp36dEyhDKG1ShIQ4kw4eqGVx/NXaLEQYEVlywJgdDVYWsiTdt8lpX1lwhmNvM6
7YXruhtphopQw3rJJOj/uVTSLd6nQiVA/gY/b8p0ZSyITGcoUaNjJNLNGYGQaEFM
/JQnSMSWwaeZF+XG3p4tXLreXOaAWgXl+bhyWiQ113S4VoxsIa/6UXg3/iI9Q8f1
lwLWsR09CTythbpSQ1/AatD6JsniCWzTlKTIcJrGCjUXpSVITcqdHEhRzkZu0X0T
08mxhcxAY3v3fZlJ1Eu4hg==
`protect END_PROTECTED
