`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8JFPioQ5ZE3Lbf1tYOYjTStf/wCAb06tZiVDtgs3zwnHFth8oqPMJTz46FY1SSc+
RHJddNa45Ih7CjEa+h20s8wTtmUX0uPfJbmLFYCw9ECZ/j3AtlSYPgVpj2Q21DTG
LEJt/u7CJjbGAL1YT/D2c5BnwJBCxKBWAQyf2J2sps2vTsDflZyAPT9UBAZN+2Fx
k5q+aEclR70oOJTYsbgn/8gUjqFqM8byBYEPK0oaYknvEKdXaCwN1mcoRvewZ1SV
0y6QfsKMSONMeunLTHZ0pbe0c1h+z5NIK2NffyHC19oA5+AKVN1ND2NrFnvd283M
aw0A8JskKW0hJyVAjQf4dZ3F+d1Jgntq//KfgV8nuFXrbwynIap156Anu0ofM6vk
dx4JpudhHqVs3ca/S1YXLlVHNG+A8q3ELq+JoauYhw5BuNrGI36JE+4YlU7fpgsr
UvaMOTTq3uoiSYobSmW8WHuV8F0DuSBOqIS2M3C97qK1Yn+MytOR5N05x2z7blKz
1bY0MrNeTij+EjniZD6XlGOMiYYJOY6sFCE3zdg4Yes1XTaRuks+CzgIb1WedOTW
+Op8ox4abjosOxNLaewveNvWQ94x0LtcaIPAMBctsXA=
`protect END_PROTECTED
