`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XFfWmDcDyRI+fyhGCdVwTJqdJP3cD2ZexJx/GNlqVmMrGkVPZieunrjoKRsGtl1X
nm9vb6C6adUZKuiEfzfsnr8FDXcCdhyYSPWbWi8Mycl6gvxodQYU4EJzrz2vFBy5
aOQViOGsp2jX7IwgzCb8LSCQNCrTDXDnYLSetkPFAAZ9oYjX4uKj4/0MaAjEa6Y1
FD5BgCXNqtB+XqIwQ6IlrP/i4uAP16O56mSAz0WhCBcrN7GyQIubCD4QH87wSnxv
yTmSb7N++ZqqmxwzRq//9ENpfTqc9P72M8xE1cGB1mBnjpvsS1h1ZWidqjq6JRe7
+j4pvNqbB1vvpVJu8r5YQvDZAiGqbYz0tydJvASyRMVa/FzOtwz5N/nIJ1mPTDWC
ld0qWPyPqcZwNoROTP6Pv2d7OD+/XpvICyfdPHD8hwR0Oqm/0d2JT5WnppPt9gWv
`protect END_PROTECTED
