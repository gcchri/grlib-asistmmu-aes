`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BbNt89etIpkDp+12iwFrkVldScEQQZhXEbWB1Zz2tb8IrY9vS8uFIXyMfqRuosgI
ZQKtCG9kOL47eCbs7gc9n7pEcniB8t8l2UtTRlf2g8LPU4ZFFlO/g27qWIPtY9NM
KLuhYAi4cIhIyymrU664Ur+i7m5rjIfyAhdBb9hIW3X7WjuRS7gJWFY1Qoxg3IJI
w44LVxGMK7WUoNU9BXOfqU0JzFmBTBHkVzDZXWUYQqkmTQLJMhk9duwkvTXYpCsA
GNl/Cb2eWbMS1Y29dCPLTA==
`protect END_PROTECTED
