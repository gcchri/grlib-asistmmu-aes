`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b7LbNnP/j1I5Wbd6rGiDnA9ERlfNWKLgDDNHdwW7QQsb0PPUeVCWXWW7fb5Kzl2w
kdf536OTErHGzwnC1n0k/cdZvgEPxdrVgHxfxJTKijbCJNYyLEz9gJLPuhPomoqs
CCcRF0Ks/ccq053n5aChK3ONQac9Hg3Dg72CEOT8adGbs4Zku3v4TQ410KgO9NSj
XdHcUBBQZ8UUDDVmMm7veDwj8n3JOuiu5XucTgBPfZDf+gWd4cLm3ZFaRxnnRass
GymtXOqZ/9xBMYIT7BMsB/hsS2nWygYyzN0hKRtm4nI8yxCDDidqWVhOIkwzgeVZ
DV2nFQDhTFXYRiImKzMlsmTqInkzYwqRY8OGPiLq+pHzKp6H2ALQjHB8J09QVJiR
pC+EIS+JmBDrroj1HWrMQDei5/aQSYZc14G1/9eNraMwh7XSj0R+VOUXVTnWOXyA
6mpBPkV519xKJixBo85+MPCnqHgNa0mUbgx9sGtZIenbs3NbvFMq2U3KSGy6emgv
xXeueZLmRNbXRi+SsmygKzUsI6W6shKTpoNs4oIcib/hjrujvfF6ttVsuf6fBYEk
gJRj4iRauLw14+11UTaSk64lU28pGxTMp7nHXnsKbzAkw+ypb/RD5a4Bnm3IBIoS
H2w0WeGjD7KyAc6kTksMmk/925EhisW0hkE9+Rsv8qde4RhooARPrArbDHviGsNV
PRWqzI/u960lfNBz8SNCGYugN8FNBChg1IYtCowtlf9gLUzlJRGTTVZsvD66dOC6
i3Wl85rHm7zna6GwHPkeNqKlkXcNDhqyTd5MucgBsL9lT80cWJbxhAfuZvaz95p9
RSTb/6Lonjd7vpB/TVq3z33qsK5K8uzejN7WtCH2cHcJ1OeTE3kvE1Yh54XlroIJ
IqZcxQQnQKBnh9ERd08TekLgocP5EHKf4iQCOqvLWpr3zAOh6Cn1IQj9JN3f5HJj
s9CCm3ruSgQW2aILqxlTV9CqJ/kKZb+u/mqIlIYuRilR014MesEhjbTziDOLjDR3
u8bnwyl/ePvHEcHIjzxZspzXfE3DIwnKw/7iDBMyf/PlTC+8U5U1J4e7itcJpAhy
+c1SoxuQsOP3LBoVwhPgHcWqiIoe9vhIcEgFSEIB1D8U1TuTQKa8+078XrbLxLls
vxK2Q+H5r84mrWomHJaOeJGT4CAyM5dDj3lSsLz7oUXkQjfejaL6Nwc8F+ZMJg4F
6LYQNAHPgEzz4iIeceo95b7ueKEMSj7Awi4ijgvVhlQJXXWhR/tdBAjxGX9RRn2x
yHTwo0Mbss1d5TZS5RdxsvVpUBHcVZ4Ec/JjSPNX7+DVYUyZY7MjhWm3V4XRRgXz
2d9RejiwCwsP3nV1vq7rlKdtB+imEvsxOtns3hi3C/8=
`protect END_PROTECTED
