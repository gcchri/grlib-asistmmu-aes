`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1m9bnyGKdIU8BfIywjeVP1C0tWsxx8vZ21lkPX0zbTVuTHCYjCcE0DhduzOxJaaJ
GZ9ocV4oDBwXaS2WjUPheofBUc5WxnCtXrvpE+L9KL1+S9mRIMwSWbj1oeQFevyS
zMYJuAc1SQNZn2fB9m1etejaYjfO96az2eOGMWRKbm79eDu3Bq8oskQK8kjuhH0q
Fkmz4VgLM59g2JBOxXVQOOyDjnaJ9qOiDMmBCUNN3S5cEAlQ1ER8Z/iCFUtRBpCY
fWjzyNDY/necDTKWYfdxy91GD7Fvg9S2ZCQdaU8H7ukJlfkm8RxVYJxumcBqZSfv
761rTR1p69xwnrw2H+KpmXJqRnbR7Ool/+q7p/GEuINJz8kM54uYv3DDEss6QhwQ
yHgaIO1HBHR8vnVMya+Cz2pvxguDYNBkSJ2L4AZIP9Q=
`protect END_PROTECTED
