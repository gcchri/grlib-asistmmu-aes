`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WLNgCULT3wvkASnKNOQJBUWanAWnPW70Xhz/vfbApNv00Gv+MzbnXd4MR5lYN0zI
jmPb07IkOhv/JToLQx72GYS3eEiAbJVp2flBsRgaBXU6MV+mjRpRKzM77vY7AbjO
PqdOYFeYsNBD3XwOQVPBY3J1I0nKJhf9O4MWHgZDhZavAOMcpbdFYob2U4SOmcmJ
PVEqqU72+o1xcVzmauG1BphV6SZ3IabQL18/wh6Al2KdjXq/o4vlNtkjKJ6mCqTc
Iv4LH14LiOsoVf+WXs4wIrWkYEpsd3gnrphI/AptftUzFugqixgtwslRM52Hm8pS
E4pdYuSBwzz4amPPuZchbQ==
`protect END_PROTECTED
