`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vqENpJg72Zz7QkyMabAHjU9RAcfG/kOx9YnDc8XcnEgDYtrOGPsJUj98WfImn/Ms
rvTkTevckbu0W8toP/IcXr3vcL4+ZoCrHxWgiTGCEfvyjvwHXQAJt2CG4cfiEmu1
gXhM6ihPeXqLrsTUxUw4ZwDTkfFoXBCP0EZERKvQwWNiMcatovNIil54m0BdUqsg
7gyvYyVcFnjUAPrj4PfkLPBo2PLYxHvJcz8z99GGkiZuwGRtk+QKkcqjuqmUrcBw
NC4domXlW/2EZR4N1weqDAHcLyUIc93DuwhxknaOxHvPqXnIBraXI5AHQ9Nleqx9
YRaL++9aWXDy3AKOdXGliTDtHrHdhrWy8c5aIBmxqy6rGAmd2pslSACBd5NI97Sz
b5ReysRyVQAhK/gHILzHyzhiujBLSMkI8TmnZ4W7QWcWssOLaZhZiwkD9TC2ppWP
+aDnRMbC3iYgWugzNp6H7g==
`protect END_PROTECTED
