`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yFVEwJts6flPRnFgwgrTr/hbeaGTSNS+WF5h4i9EwsAT9jUskK5zbFp7ikWY4SOc
fWMWba2s+50JCuRayaYNEIvN72TUKT5SZqniIBlFohJEclZyIgBeUbBuKjOa9oLE
lN7WaelPDSOnRWrUGWl3sPI54XQMqa13gIU4A7P4eHl2haMaq6njJm4GlJPmgssx
vZnSnCyRjEukRK7NOVhg5QTuUj0KCgQ2LPTdzOXXd4uSL39JGKtFI1oq2NDOS6AG
XIm2UmSHJghoNc7svIuRuuH+hiMKb8r40pI/8IN+NZ1a6K2K6xjhNnovafS36HrU
1Vy3RuBvI10EjcRMwbEJjpoah0UyJ/l767IQY1bMnOSufUBTbQcW69uq2EyhYLzP
9j0q1HW7+h3opMCgto45RbUL5wUq620l+84fHB9/RL1+ZGv/8YufPedOE9uegGBN
3Cz7CESw8guVD7eBTjXWaSwnXsy8eor64PrWd/RjtX3hxIKxF5koN429tTiHqvtI
yv6qgQ7lqnrrP37Lqkcc9AevjG+2Hhxz18Q0yDGRcaZ1XD2VWWwsYSS9rvymbs1D
mqiXwYXz9G18MQ6MBZO78mhTbMukBUBTZVsJlzp5DurC+BPcFzCik3UVwAq36kSw
rwHkn6ccNQt6ITj0rd9tZg==
`protect END_PROTECTED
