`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1cxiIIvfD7W++8TiglXD3TvzLJrw/ge/83ZXXVMG8eZ8X9vYN6i0CP+AQN0kDhNi
DYznnZZvy0k2L3AYPpeuDQz2UWFYgC1vIPS0MiLf4yD+v03pogW5ZCgJzZODzdbd
l+lxNsdQcToD8j+mLp+2+5IrT82KyHefutYMbY/u5xj3Nk7ozeu5wq8JuxQlc/iA
a9M+KwADjDDfpT9DaBlNgbEiowGYb6kdSewHzoMMyitsjKKaGEf3cnZIrAhEmUbc
ZnVNfMbJG/c6BfiJ8YqtztOAr77ZnNo8GcDeMCl+HPFOJ1gcSAwLEsJcrKb/z4ws
436GYZwxdYk3ZvIhtFFH/jjoCPnzI/38JRQ8lVpc/pN8OMLYQpUAHBHJp/DIFi4x
xDDTH8G1S6yWKFS2juVDKXxLCAlOgJz84uGNbCjaiZ8bPmbw2S9R/WkY88IMJBXq
ZaYKr3r/GPe9xouFw0UDlfyieTylMSttoSDhQzyAY3Br8E3VCmGGlCnf79rSNygT
laubWolfMISqNxcwwvjw5IjleJIju2ZSdxiFmyTMQ6wx+yPFrQ4xsu6eHw1MyCsR
JJ3KjnUvRWgngexRRGS+Ot3CaxV+/iekTgVYTt5cX5uE2sKWdlGIQRpcYa4SQr+d
9Yig4OBgjnnuUzIDSjIZd2Q9iX0quTIGtvzY3EUzHl3rt9kN+bFgRLaR/iwvGz4L
JtAg2YBmu/ltK/iVM/ClkAmMtEQZ3cmH7Y5a4CyveoAHw5j3KncZOwNxo9lY8UJC
u96hGDKLMQmkfD6IfmHXy67mQUBaaz4vPXk5c3rLUxg=
`protect END_PROTECTED
