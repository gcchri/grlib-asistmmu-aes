`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4F20cHeWfociRFVAovfRZTLStMA+OJhHhmzkDznjARUkxLz1tw+aEvY0rr10OL5i
+kz1AkzASRHEOUnf1rXycsFY0276IVZ+nEQaU2VSlqJnw0LTYg4XJ4ZRKGtHSY5L
3LGo4sZVpUw85n8GVhjdeA6oeJLp6CVtOaFkdPfy1c5dlW5T8dm2xqlxo34SEGDm
fH1q4RH0icbU3us7fU0WR10hA4hrzl4XbByF8287OLNH0kseW5vYAWCP6v2W8I3T
jeJKxmwC/kwz9OGPzzzpIKeacyIfvO1dWudXpO3p9Sv5omDdf2E7q8uEeO98XudT
f6b8EML4wA2ja9aODaPLT5FdN5mgg8j5jnwObwx/AuMPbuVfBUp6aLbZelv6h4NW
MVutAsbrk5scxfrkGY3b1nJjCAntb9f7n1Zt/iID7GwodMYlogIqMYyYzYe3tJ2z
+5kbjzo6T1CXtDyK0RNgjXnKPB8RW5Y/UJUehBpQY8xflW2me+2h8Ekd3IQaECDv
7vg5JpiyxCnKOT6HohgMmZRvP0UHZAOHmIq1EOFLWiMBv7unVvg6AFkvuIHAm7v7
Wr8Yl8HfWHX8/IjtXYSDgbEhT00Tn/x/CktREdPBsRAb3PaXb/rJE27ZZA4L6TKl
zasQHOpuPgDBnMXLUBqtqNFO7u/ByZX+p3MtE2EQmDVrTNl55hWchwewaKNu9TKo
h1YkZvikFaTZ1JOxGpzIduufTgoWgv/xnx3vsI4yWehC5blEYC2xpbPr2axuWgRd
z+lNnp+Qg/dsMkQNG3QzduNogEok9WfDKG/7bFcmfI9iazF3CG0hYpat9gkD8PGj
k/UQ9hA7EnI8D9EhcENlFEeyGHUaaxvZC8CuPRfXSbiQZ79W+nikA7WIJzJoEkDF
Gn6RJa9PwgzdofCymNNrkVDmTP33YLlTgLDTp/fwPqgGIfrrNK8k05+NXlwc1W1r
oCmAIBH67OzRBd2w5P/7imcaEduhzTPc8MTPRM6q1r44Cknzgtre2okQW7znv20P
nDRW9MkulBltE4Ehe46ikNaFMlbkvBDnFcVqZDMvHZ+x7ZRUV58vnPb0K7WGkOa+
/yjBQo+269SLrnUNIRDDnlq8CwymgmIqdDl0VFCkZKuImOyT0+RmoHnTx8xg2gNK
MY+csS2FEAiS0GmoV40PoaRiQk+K91aHFyzyuNxct8r/sRunaUdF411MoEExyRA6
iJ+XIPGaj+5ARa6h1+1LAN9DEC599+snFCMcQBoZhyzOvNQKmD053Jpf2yjPkjSW
5j+ltTuaEPns77GlbWF/V++IuvBMLS2SNwO3PUsX5OWmAHJ5nd6SThMpjOKzO5ro
guX5Bz452PgOHjSbztJ8OLpzX8bnCX59/Wwf3joOUEDkhtoCruR4vCiteqpTAlDu
Iw5u3L8xGsHTXJM9+OOnQU77MlhrDYJ8kSBwpSMReBG4mPTH9ezDTvuGQEhVy6IY
g2fFpZPKP4u1F7Ujs4JEq/w+n8Kl6WnjHvHIbAQO62R23rmbX5gSv1RMHgxjmuPV
BtRtTqcg7riNcjTa9ThCQ447dXq2YgmH9uthVHj37Z1naBLZwN7yZPVvjY+IOhk8
+jnp37LtN4Pt3MjAUvUU7MIyem3IUqFodpCnpdsbf+Sk+w3Yd0RZuNRgOrCQhmoM
K6DpEj1i+6AHiwlOByBUAqNsZtRiloWQmK7N5BFEX7hMuELtq/Hut/Kq9Er1oA/P
R8sea4kf/JtmkXvAQZ0o49GnhzBT/Xw0CHtPfbizmaBwW+fYF2nuh7ytNZ1AGpFJ
AR9K3z1D6jvCa2nPBxMrnpb30rzvn/NhNa22IdIxQRucoljXCI/W5X2TBid2uqUn
GFylIn1Jbu9jqXDY8Uf0fvzwZ51f+RlXIGSxAf+hXsslRKRY5H7fGCGxIITtHA7d
qWkBZ82UZ/Vii4QK8vNr9VBZNLhkPGURIE/trcJxzHIMDqxjdFE8xu8Fm/F6qdFf
nuqfzXQOrbei83cGgL/zC28fx1s/yR5/O6vDjmzBQpLEoDYAz+ghwCNFnFtJmgyp
NFjDO2QjvHaZdchQwVbleA==
`protect END_PROTECTED
