`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yTsqi9S7+yzIlNDXyDdIzRlu4nIW0XiZWbRN1JVFv5B3vTaxdtk2EoNKjxcq/arH
n4pj86kjwuK6g8pdYbORoS+JqwypOZ6YODK+oKqKjKe4H3BJPTu/rYctU9B9XQFv
NBr1Qxh/ny5xwBWrttNm5x/eMHja0Yu3YFGDEahnfkepoN3WTGx68R4f4shqS1xQ
eDTIp8yx3GomPIjnWCw6MZcxYdtm3QnC5JmKSECQ2wHHDokSoMjl3B9AwLHcEB7v
a03yvqtZu6xJW3iF6vK4ddu/XYJBlagdMwoipUaQf0dt54uAHMaOj9D/dRCQQ0Z5
M60K/gh2UqxfLjp1nH1Eildb922dPZNx6xtFbXGH28ru7dtlgQg1oSN1sv6YeiKe
f/OA0eOhVCX69UQzGlJ3IHToyXZ29jFg4J4rlxLzkvi3BXgpjEbvXwaF0yClhLvI
pVPRD4RilmZvmaCWjwnerTjw4K9NJbpmI0mlsMDuDx3i7zINXbuL1FghzQTP9WzZ
s2L458XbX1aKnBTFFCXNoeKr3RSpNmu7309NkPuDdBfVjw1/0gjhkRCPBkypCIxv
KiBMoXhhysTk5M2ZhTnYsa4EavzaD16JDOldw6KRN7kAGn+Wc5pqPEz/tVXBCxL4
3KoXJBZt2fkEVLwYt64mi/G3QigVnyYuICaKf29j42X8lWRyStyut4YgojVw0IfM
j+ZjCynDbTbYVZN1LVLPCNeIGiIMKKN48ASWvMXXDcM=
`protect END_PROTECTED
