`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V+sNPvkxxNG7kbnBFz7/PBzsKk1zRMQujufv2+QL6kVdWiMWD64X0Ii0vytnqreH
Jn6jJGyJmfb5n4FOhiVqmx6NxSU5W+Aa0fzzMBREF3RSo+dBK5eoRUjD6BdrxQvc
B/8pC6hthVLM89OKIYVBH82W4WmzhnViYF9qukYnggayzQDPyzNvEDFEO/ysiKPk
waPG+2R4InaYSulAGASuN/dIrD5PgGiMeS7Ll6Cm0TEN3kS8A/47BcaNvjHvPD16
DaLMVuGtzud5/OH3Al6WQDUkOaSkElNvBEg8ViRWKYT9FuOhcrnk9fFfXGifXTqW
d3cVnjsfWdM/S8aSmc/Upw==
`protect END_PROTECTED
