`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PDYO0nAaUKuBhaOyGW9RjUjR5b1tbhAhAs0cXrVsn6P2acoFwsot7VH69Nxairdr
JMdTe+1k8bvKimDxqdOWa4sSCcKvL+lp/rns1JHOA2nYP2LRhtp9I4FkioQBVEdp
Hd6RejIgkc0m6797KrYv5xngA5vPLt99RPNN2KB8Xb97Ozv1gun9eMNxKMDIVbwj
SAIsLSeTPgMbisU8vakptRAX2VsrnEZ5qqoyOeEUPyYUHBo/oULXHMnvabPzzNv2
ovcf7Ca9mxCP3LqyW7NrLmSrNIec+D/brk8YVrSq3MM=
`protect END_PROTECTED
