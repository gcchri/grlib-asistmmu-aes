`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AcK0jG3MS50wwv4wXRrsaIXohfcddSuvC+6KiwJdY5aN5CW0so2GtWGihovRrybL
K47TjQiGUTY/uCzvxz7BJk2o4tkXNx85rwd/U5YfbRLAiefWYKVKPkWXHC8PqZIX
iSNT/HapMXtcJi68qwDjLIba2M+ALBBoa/gmy+CVeTxgYTI/yy/XyiQPexDxxJjp
5ZH0l+2T+ayzrNzEPpaaNYBGEIq8/jDKW9XWsY4UdjLqxXxxKLelpWzv5h+SCpWR
gakx+ti1kh8xeiNd2VlEQOZRgSM1QJO95gXsg9Ak1ht0/v1Yt1LjltAQ/jYZF2Qa
wyAQXQzxtwK0L41TVxNe6C2u0P+9nR44HzfNLFTi6DTbZwJfcbhfxvUMyY/9UZLY
PfwL5vhS4VkW6UBEVT5YKHj92uNitJ/LoaPIBe2Hgoq0nQFHUQkC08gKwDbJhvUi
TtVCq2NX8+hCzm6+eyF32Sitd9bVbtX/0+uaRWxtU63y/GSkytnxo9lLkEWI+LsR
xoasysKDzxXVUHwvGy3X5OI6tJVs9UyVRMx6XDgKt/0SO/AVAHuz7qaUNE4eRLEs
uqP1dsJsjdZ8TdF4N2cb9HjLnPtr4cUAOVr1K6icmlzJUNn+Xyqlu8+6PLE4KGXy
BH9jauaauUEs1hC3+QinwwLrNrVYR0O3u6lqnR9qxPTFO70NDs+zp9eXzxZVvOg4
t6/NNMWKPKw+azU3iAAcyIJH4irCynkQiwiQeGeS1kIRFEjqYS8uiPmT/xN7CLVM
kj0hW37x0tVBuE6pOeGaV7ohlVBEUm1SHNMoE41VgZUvHhSXI0crqb18tHqJe/AJ
sThTrRhTqLTQ9GE7yUZBs6PLygvO1xK9yM4jLUQLkAtM9BRaq6NQ030ImbZjo/Nb
WorYpSxDaj1XiOrWj1K4LK98hgbkfIW3kmn3cR1vPieefVXmTtWthiEd9EQDxLHX
AeZUAhV92NgrfSbR40Y+gESeFt5j+44YLH9DTTd1LnFiYT/HGfJ8krMFfrGtQqrD
1csNjUg8XX5crSFMCR7m6pPJdFdBC8Q0j0DCCOAwgokiIYUJBNimZQJtePno6/R0
3Jitokx7szMd7Agsh+MlmpeV3oulPhYAc9rGor7R7kEVqpEOCgkRRbRYqBCK0SyN
`protect END_PROTECTED
