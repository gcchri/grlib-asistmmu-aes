`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ctaGX0saSi5cV7028Qmt1aqXqXFdEqMvu0sJ9svOIoMNJsJU19AXQ0nBb2+xqTOB
reWq0jlV6odpzKuTYSSWELvmWX56A8FjP/CRU8cKdEXCRoO5tPx4UFBiGDyl+hIt
w2CJ7YVHuLeTZSKwhbcXSffYwCK7wxOPgZOo8aoetY0u7+cR4nElqhaqnw9ZzsgN
6OlJmbmbKAXG1XrJ7BV2MRzcapsc5nmA83kEb8+sPTapTT6h215adXq7SuLP5h7e
UST71pC2y5Hf8SbxiWTj2bMMNEJNkicv7sTE12JeO5XdptqQjPtRdI8cyyAt2CJb
qcmEaCVK8xBjeWG8M6TfMQSw7eTa9d/ev/uT5rOFVKstxaWoR3uNbnEcytmGWp77
e88ANdlbbGkPeSGdwIkYwPSP044zvj59B+nhfWdqB2O5u76GGv0IiJq1Rptt63oW
NDa6oIfob5ThB0FniypR+G0lqtxM8oNZUzG1mCJedFB5XM7p93UdK2XjF7v84gtC
kFaT25qTkWpGuorks93E4BdGEPoARNs1FkmaPgLHPJ+7B+wzhOuxZzCzjDFLruIW
H7PdNrUpr6+d8IWXWp09qcrXsQmQIBbxaQ1ihN/6o3p/O/t6jyACN+wbBBEsCC1P
eekcwrDAhlrKMX6Xa4KqNpWe39xXjJYJHJbMN1Rnvj2QGDXNqBb4dIkYk+pwxHtp
5lSYkRYxZEahciSnK8O2G9/kOqxpjA6Gtlws24Ye5HWTPt7myoj4JmTnSqyaIJp+
q1p78YT1yNr/aYX4IZzSeg==
`protect END_PROTECTED
