`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m6W+lK7K8XR3TYce7NG/h0+Row/I1gQZFSpdepbs/brqEjbwQWne9gvTplSQWL8A
nLgsj6aFXBn+kFhsm3yY5XHwku07vKG7cRGDpldqgbl8agJbGhd4H9qz6Cm8WSjE
X1zr+7GKOYBCdssSakJbVjvtiuHhWprYT1QBFCPEm8SaXY5IoERhZd+Q74/hU/Y7
r+oj3DShjfwJN2MdOep+rTa9+vzFrHQrSThdyMhTNnXPHc46qGNao7ZL/Jr0S2uf
zWGRm6jpEh0NKTrurZ4MN5qf57XNN9BpSnWFCPYYFHCsO/dc0eLHDQaSEWOplG45
naVdLdgeN7Lwqwww9iCxwce2gvgIPSTvCzjJu2PyRQw=
`protect END_PROTECTED
