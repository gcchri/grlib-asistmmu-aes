`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iW6dkJeb6bheaUeJrfwxcO1oXwpFQnZf6cSHO589B6bSEjLu5vCzU9TlMbT6a/C7
1vT5Mq2vHqpkePkgDrWQmosVvkyT2r1LHQFvWLLITXTSOxHFA+pKCpbrxXm78tDk
qorEVbQVreEw7lbBNYNncy7aU7OVEL4GWqUsC9B8A9pL77mCnyB6H/uCgfYFdIm6
wNZTKja4jEsOxyfk+32yVXbpF6UeldmGB0xN06sEXcUkNL9S5ZrDqTDYSDt8To6G
3EHYBeYAlO+TGIPTjxx2YvN16PLjg4CaxWyaMR53ZPU7oGjERWt6e9LEuw5LXL18
SshFqiFsjd4RLf2G0vtCmVoecig7SPMCSYBSyfsvE/ptk4VI3bIGJxvmYi82W9BP
ASpdOQOYu4H/JvYcfHnaEiKoyHH7BiTqAvf2ByG3rGLAz7Klxa/UEiubxPNK5j6J
kwe7CyEVIk5+4DWdv6npC0Q7my5SOZ+Llbq5vzVVhuwBquIsoQZ5w6Q2mT3kF6jN
TfPyIxdggpWliEiDKnLFQvtoDZVovSHSBRbSZ5QJVrTYVgKPjw70khctYSz2bK80
`protect END_PROTECTED
