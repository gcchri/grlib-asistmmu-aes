`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u/SPWM/qRBFawkNEnNhuG2jmyPhXncmGksI3Q46ghd2ZVSJDZhqryqO5WkUkV3aI
q9D8fCx6XdG1tkYf33AP/KhsOXyGercmynB1ILv57dw8COyhRmiyOwIbNgeeYViv
YBIZ6lZ/UeexcnXCtnVHj1vgT2XVGXAJYcCenCxHWEMtPU3jMDd56PcDZmX308Wc
ACnN06gTuc++/v0Nxdkt2wDb6M5aUvponhPLoU75oEu96JT+pX7QFOK24aMgohbq
nFnn9O0W3MDLuZrm8+dLlptAm9gowXj8ep9QkISWUVAPcNasykmc1Ay499ArsU5P
ge/amtpSxzeLKwaCqwDwYjMz1nwwi2a9YJo4ZsL31M5+zVSkWDdis21nZPaXMpKp
Uit2MfSbxwemHBZi6fwtVczEwyffEa8MQfIUTYKwXsLMLth/4N0Vok2c/quDbIWp
Z8r4KSkSNaV8TwD2+x9hFlL7lh9102CeEeZq96q6trP2sXPc0dB0ay7daPKeCv05
0z4VUq+3F11yXt3Le5M9/BSXVE+nvY1h232CH99OqBsF4//u7xZ6uxrvdAnl9g5I
xFS2ecJV0CIVjL4kgtj1NqyYGvk3cc0XMzGIA5q6iRb/aJbCZl1vpJo+U2vQSoAt
R/Udyhx236X4vrMhaRFAzSFeR4XmV0fR/z6kniE3mkn+WRZOWW2/HutBNDDxSbSH
I8oucaXoYp3HfaTShwkhHKBgYMXAjN6anFQxC9YG6zTFnHDYTJ05wyhxsi3mzjuP
NCj1skvdyKRsTwzyjLvY/FJ7oHldRV/dV/qxaQIcmXo3kmrancrF7vrAXfYAynV3
g2D4dMhmqvJxgBcRrewyneOJkY5YWEhuHvIU8je7ckdxN047j7GwgzrPU9+P/NSX
UhzIEt2tkkcnX+KIDIp6qj+ZoSCaerRviLpsGghQ/8j25VBjEfbyaKhsuZ0KPjIW
h9dvAwLxp7RsFTYm/QE9BDLKXB8p2JNvQ4+F4gAEpKrYSVcEAZO9pLOUobDpJ0s9
uraXLM4mfFJgVyITmGcUleK1i3qFEyg1QmTLu5GDkmMZU68h5COCNsu3e0vFIv5J
o6SvitHdwbZQucUHoA6+pJC3d+/pdcmqen37R41NfAqnb565vttJFZrbRV/zcAZa
/phDbfMSPoI5iqDyVc5NufvL1NGbLcUxltfSDGdkbJQNkB4P10DATsNCIM7xQ34V
MgjaOFSaoMCrjCCn1vYp8qo5/0IuE6VSC0kr16fkF24BlE/KPrNMJ5/TQSDPtlJq
aBXvwTx35/2UcsalMmaq/XgE+oD53QpHsHUrfOPeBFjObB8uwiR5pdSBSGJwYZXb
G8BkBJjhGwps4OjDHujg1CBA/QyH+yHWRhl+YukxHZiRjSwJlYu4dyJ6+qF5Qndb
7a7Ri2RmjZTjhYnPiz2wk+hbQlFG2k92EBxGfYkIi3bqPJEZzy7TEYeHphyt6809
tlH/m23INkVPUGTZ80FqRRsWygfyBmkFIFcj+XfW6uHfDqEDiOFGGKhvSEDesyGS
C414PYyMaVG6hPq1eFM7cBwS16hOsn5lMIQWDsYbHV1CNLS/4O9IuwsqGeeUmpGt
18w4yeIG4fVwFaoZd5o6N24ynwyR+k0spqHc6NQT2rLQm+0er/fwWUenbvLBES2d
4yIxvvz5DizfIFRc5A3mN9liLqEVTR/sJG4DYULtqWv3D6nvxKFCHZlDwlh/0vEL
Z3Z/gmbitCeKKhtVPz/b/VYN5BtCs2doyZKJroFZ9/mkFX74EeVQZX0VUU5xWl+t
025fTP0wnepxKbfcjiUIE4fnu4zNy23kBd1tLg+oV8ESp4k0GtQjrZ2JjeX+UXa8
dWx5++58oyuVOsXj+PvaHhCvB+lfxK/Lgyhj3Jd2bxmFMWOTCjmbZKXGOUbinhaj
QS0yHsQMwTPzOI7ndcclMyKiewsFq2t1pno5EcOiIQQvaZtL5hvESYu4vONTP2nX
Vz16gmUJm3+6K6FOrQuNGQ+86A0jsP8jtm9XAO47MyiX5xGvocwmn/5np4TglRTD
nt7e+Vu+GQfg2xuRyFP2JafJQCrYbqOoTXWUUnhQk31Kf3y2GH9JJYJufTskdWCc
qQl1mAOzu4lwH+815pzwGFPNCwJQcpYFKkxnWWEbSA3Ch0sJRG9S7+XWYA+EgPvk
vHuwgXSAJhS5v6qx59LaOiBpJIffn6E+ZGZ03fqmrnHJxWOpCLHnYTlb0JFa/Zst
CzSGXQc6Cs7JKDGcWKkhoBC6sZy7Bcms3lSEKWzoJgSrmtR59h8OhhCTGvCinWpB
cp1JaDT/9rhoAfWzXEiWpIj5f4WDbRYysOWRiYOiG4ql4dyGmD5oYnMxufO2nnsO
63YOA6LffVtMDl1I9ur8Zwmy0Y9+FSUo5M+s3ySAP375ak1Ic2gpUNuvk08cOhvd
ZQaozMmbFUrVpDdeMwIhUHJ6QKK4uMugxJ2OABul269v06G1Juzi0N4dcST8BqOo
3XzS1Ka6iO1HHbFXeDIppcgvBD1LMMPKRqFBnMvz6AZOC+8o3jw8Pd6w1yqbT18R
M5I9Tl5c2dJbnQTg4ErEvqkLt9g6ndQsCtrdvWtCKMKmFQIOSGmmitUkOZU/3wiZ
JH3tsoOX9kyU0mbUdvI6MmyeX5WbT+PC5FWLL/9ftBWMLaGk1aMMvekAJZ42tz2U
eDygbRHQmn6WS0q4XfVk1GZaIAiOc2s0hpQQPGMwvo1XaTnF0Ua12ZmsGM7Y7yH4
YIkL3tB/J2x1E7trx6UgjX5ol9A8x6lzohJth7RPLpShRoN8HPZXX+xiaxR9jtay
NxufexlYhhzxofDFtfLho/LhTVnwbuSW+3wvjfS56YbBaX2aJuHi9SOp7SRVZcaA
ajSV1bRlyKA86ft7Jv3WR5KTHoh7Z9hYgkWqjZzuHJwnYwnlYJOzXX/lAM/ldT7A
bBozbSbm3EandIY/PltxbotWFatnsvgN/lK/4Y6HgJDF+pT2RzhaJS0SHFGGlKUJ
FsyDBoDI4uTVGjwbltBfiGnJyxzrc8OG6YspqFjqln5AhyW7g21f0yylGCzmCAZX
A+wqKMN+nXqpkCRyTkIqjDDHzR3mEAi/DpjOrZkINL5EWUiUKSFHhejTkBwAeNDH
+/ZxiRGkBliy50mNqKu6hoMmvb1Tt4SEFs9x5bHLrVupjZsXLUcRi0Wo6G0GFUSV
kJmsHdQXqHBUOJZPD3+bzZBRKIw8eH9tAlmZXim8kKoKnKKwhfx7D9Iq4MgohYoc
cgwZYyWWUpL07Yi0H4lvimCExUa0FQuqfo1AoR8MMP1qyliZ3Yw77SADc2zexhUC
zZ15r8e9J5Za2DxWJ4e/mIr/OIxyRsOPi3LRakhC4CzkVE84htvXqVvtBiAI+SzO
HCQw3r1hMrN+B4l3GoKUufBvR2YTCYqm2nDhg4EQUTA1y5bi80/tBBdnwkfx6ypJ
IIC7gtOvBP4zJ5iGPlr9JEfuBjfivmvTEtCp93nz5uMi3C5RvWJDGFoP9Ip4UDta
KiO6xpCnZP1v+hFhxkTCDmvruJ3RDEHPC74erODX7TB5Q1UUSZfj3rnNOWQgv8ZW
LZvYAbzyp9tzAYwrzUgrvBWYU5x7LzC5xxU08wnvHp+m+ftAvZacOsyQfzamccS2
9zNBQKzb2ksvFB/qoFq9fupTJVkr+xgOYpvNpwJbUD9sGfPUCg3lOPZ+BQ89p6P2
uZD0g/EKMR9ccQAxG0BSj4g6Jbe1Aww43Lu8UeC2qEwEzCQam2AbLDApgWM8rl+q
uV6PfBTNVrgo6tfvAjoJhH3yXmciUimvK7JGsaSyllhjyDhXht84VEKmxj/cnRNY
qbdQWVXXPmbFMTb844J7JiNo7zAQ0bsD9t2xK/zLy9GnPaQkRYHJeAUrSqAY+c0m
GWThq1gqpDxBswz7DMoL/fbC/A2xypNAv50+YSnyPG/thdqDjjZs7c0/yX5/Xodr
le7Rcauyq8zxuEOzZplXAqM/T3eMxR25Y07P19KP7tTEomigh1Op7Z6YASHvtHgf
472bGVcmckPQ+ypl+7yp10snENineWIO9kJP00rLm+JGi2u0z83aNuf+rjeJUzAF
p84dEFEyG01ZP5Ma7LjcXim5VsS72NfKahMg5KLFwDshezNx1C4nGhRaH9PTmLOr
JcraM7a0RTQjBamvOSFgoE6xgPhrigv7TYXfIPXdkP7rlDxOiah/8tTaJk6mCAqS
r9aBWB6WKiZlcYcQ02mcxJBUgZPbdNzo7cTeb93Y0WNwfpoefzUOTMZlYeqkygmc
HPOO8Mqt01aDwlt+gxYA+Pcyw2Xd78zJTUheX/j8YyAIlsyG+TiIWGm6gVdxXOZ/
lTIkhELHkN0sy699mlx+XwSbb1Cyd6YBRsvqsetKaBpfZ4w4Nbexv7GXAlP8A/P0
k37pRP6w6oVn5gIkMStfh6BvP2xKFLU+wB1R9i952I4vMlaafmBODkbJc5AHc4CD
f1U7+E4zuIxEsC1SUiW9ZOsuxfgyFk2YcNIR6JtcV4xX0tIrQr4A7y9MnTliyw2U
GSxDZnw2fOyKA253n3b46kvB3aYanydZm3Q1C1cMlULSVqUvwbWpoUJAuFcjQTtE
LyiIQk1JNcA+03FYmN5jfn56G7+ESlJlKI8EuXqXwQgEP3mwMuF7Iq8atZSgHxUd
wpieW2j7D/F4hhkR0gU4yX2X8l0GKNEmSHE5aPkQmbbuTTgrDGGHSUwkIwmec4LX
hDfmR6XkpBUUE/TloXyEIfQTGoEFvAUOhUOIOpcQiGYKLKrcUgyry+JuNoQlgirp
ksjOR3hvWRRrixpXF8EYglXenoXgm5/8Bz10W3tRx5W8p/zMtMVdqA5ZI0meQjBk
3PKVvx79KMiS7oY0N5PWJ8mOpR9Qmr+cHByDgH91QrKu2boSfTH1PdaoHBmVg3Z3
WRNiPmrZKBEvwflfbLndhWrfz2YRCohQzcZCB+magjW55gZ2Z6hpR4eEjYHcLG8n
t7p57Q7vscbu2YE0XlyHAvdftByhW9wpuoyDSy+m4p1zQ4THFkCEbR7clJPGHKoW
gsZQnb5m7C23OdMmAMjEjkN0zG80M88fXn7yWqWpii1tqBni6XkXJ7H5H0JISWZv
B8n49bX0JhHy0dBoBkXZb4ugMAWNx5OU2gSXIGVuP+XcI+57z7sIl5VZ+JJddMNV
btK0HJNVUHTedyaplseBS1zmr8CpDB6Q7m8QFqLX7cdBPnX98v55MVaOWg1IRgTa
xs4Mj4bd0vOp6z/c5b3uzDpF0Twg6NYKIvZ3gd+ficFD60kPIeBos8o4YBd/a+gT
awkrLU2PpriaBTIXzPevZQx4NhUVfXfXOBxgO1j4oMm+tGF/Z+8L+06shT8MN0tx
twBkbmoU4Wbh0qVINrPuDovtO9Sr6gnrh8uPO2wqQXKMSvH1pO1aWojuqyOMy8SK
QQtaIuMoglfZ5WV682ohT/zTiqS4Yg5C6cWKc5Sz964v9MLdB6D8PsY90GQGLLsy
3Ishrh1Bvx307wx0Fo0r87KqoZz2KCs2YVPjjTBGJsSTHnbmGlx3bkaRCvdKtIx3
B6MZcEMJIgiFv5B95DeUDFfIsFAEFTQYKuGDb8JA1wKoKh3jv67WLnnJ2Qm0CsCV
Y2fULJY5m3ZDiE4uFoLBDDAFJxsaIFL+r/ctqycH6QP3suZ5IHSKYueBwC8dH4WX
C1gInmYVim8GBR6tsB2HhStTHzA3+GGOr7bhhVpx9+R97vDH94A7G8rZdOwmiW5R
SXv9jdWsdSlU1GmW6/SPcNxoZQHQToxLU8gYyu7CZo5MH8ZQ2cz9GjCb5WZhlew5
tNC0xmcqC9aPrk2Jha0fP7kqiy953Wcqu9dc+vT7RfWCLqkDCPT2Imm3DcR5Mr5h
0QCGvA2R2bUKjMkeMbI6THz1Kx/3WOe1XLYswaKEQ6Z8SfUnbUJion6zM1B9WrJY
KpIk/GgLo0XS1KzAUKV1NLgiqVdzfcke9EP4GruTiEXa5ueBfQYByYb6gGSkQeHj
H4WSSfiDC2alwLS1o34Xo5vJJQTFrwHhWs199gmDIX93b2a7gJq9WxTl5yWZlLm7
B/PIspJl32x2BaTr4pBR7V4NuxpSIVefBt5W72JEo2CdxTMizgT+2tknGcJ3syua
h4kJMEueuzo76Hgg8QD8nf+tM8hfuuJ7WgAsu8dazfwTcvXu+HNavdEMW07ZPnBh
a2HG8yf1CR3bTgMDZ8Nq/rwPNcjaD0K6ORESVzPeLuDe8MfwThNcf/c0zcKbSTJ9
GXTcqAj255NXlCyI2MmtE0zYyK4mc+tZxb+g+AaqaMHI8i4p5ARgOJ/oMmWtVRLp
6A9ab8d1tZUQLPCD1DUTNU4XTFW6y0PzcJcNBGC47ZkHZWPh6WqxlmqRv5Y1EA+a
huyL/4TV5LSy+ZV/oqeMmpdjiOu2Cxmt46ip63Hgg3bEZSDO9GGXWJrLcyRaxPhw
EaMmAF4cKw+J3rudX4bHJAPebw0BcJf6gngMaAJ7pcPU30/X4KsVCLZ1cb7Zf8QT
UJzaKNtBlLUkq5mhmIuU+PGh8o9GKAmvkPRhc2mvr7vwWYgQpiXlmNg3tEcVn0Ha
xwLEQPzPzf0dcd8RuEndsiS6gObm/rErVuA15L5b+RE8pUJeXKXK7HVNCpX6EtoA
gKBYu6wHyatbKXLVkJVKAWMKATy2usg7ahXnXML9dQOic5JiP/Lsm7xUXc5MFiRw
CnaK9gFUd8v3cEw6B0wvFL5VwuykVfcuYUVTU9vvSizL8WC5Nn7mNJeQnokUl6Qm
MlOnKc2SqpFE7GcpqG073ruMJNh5jSm65qP/MelbUAJbOvc+KrIAXfjTpIZGQyGs
sh8uu3Oi/FHxw8Uj9r3n8gC/cy+S1TIMsIQsDNzKTZy6Qhjm4j+i9n4pdRhkwZQ3
Ve5B6TR6SiWjGd9IM5BuYBRagk88dYgnh5+MRq4AHwcWDOza+Bd+J7UcmdwitUdu
cXnkMy81gE9zRefX03Gd8wZ0H2SFMDXAzozoSRrZG9U4wTXNKfa7rE3XpAWuipjh
NgcsT4XWi3Y5crNCvnkktz+0lXEjDCY2o+eAt/K2sPDcrUlAfV7Eg5Lvk429Az/+
j2jDP/1pASFKWfwrCwYmMT3nIvgPOqnczVuBN914NojnvxMjFugnkf4SqjWD7j5h
Uwx4SdfEY6UJj2FykWQYGjpf4OgNooF3YI4sjj8QSC9YvIksonWKuWIOVRcml/jI
E0opUkH36VKXuJa3bgT4BKKuPP3iF3gCuhs3c7i/jfcgvaAohHKlG1+Hbl2mwNJw
cFjOXSOyrPw4ENzD3esURX7Cq9ZZebZkCmDRacL2DRKfU3IyNHWOOOfbJdR12hXC
uYB4Du4iYofSgV/pjEBHMkJUn4zzN0tcmLcc8rsfWPA3ZNSHVIoVHClNNIPskFJS
So7zkS764cEzLHhxD3DBURuWGpvDnzhv8daUmK0tsLYIC9qSHJiJBhHF0+gmyPzM
ieoI3Risrfnlxu/PAPk56leNbLM178UqHTHSBZ/8WN51k5FNfhhFGrsuxyp3hnEo
g7SF8CkAScXjdgGZQULt2cua22xQDPTrE7cc8D18TvG3tV4Es2mNNo5gxbEs5rmu
DbsStNhdGKjRhgLrDE04XhgbGKKiWb8NhmzkSSklPHuSO3GN16VvLn9TNB9k0i4W
jhZVMngDjZt+bHmocuJ0bygp/1Cm9CKMA0/S07jlnQsHBhC7q9bQURIt7hY5ECUJ
08arw/386Ygkac+6FHplDYQNFmHC5zWpcl3sKN1GxRCcPPMPR39R1m2b9YdFCUno
YESPEcCKH4sknf1lbRUNwLP83aUWtQIHOMHijIuqyfaXbHs4TmAD9InwGwsHyYxi
fSOoObPYqFKPkJ59Zv89QQvijUR6k/0peFW5dXMUUqBX/CWKC2H+7wPxuk5sSdcd
Tf1Jo+Ywg7IlJyzLqjgTkv/tCQLljfx3OjWMWvD46aXwQ0CyHpWvDE9Qo9IPwTzJ
yzACd5x7J3wY880Em+yM7XBq5rhJioOGohjm4tk6CrJRNOnzImBsx+A2B7ObLa9E
TOyd0Dxkf8mO5v883j+6vHYzvYj2g43+U2frcebJePtQ72dBcp4i5LigXDqm1pWL
htTLHi3R8flSiSJYFLiyF6aHtjsXJGggC1mYapEkr8MxnI/Mhdp+jo+F88jGx+nQ
5I4METId7mMZYGCsoJvvdXgYpEPmIZ0n64tNGMsHkH53sQSfgEVnEc0F9rp+X/F+
nfxhK7FdL+dGj2xYU1fzKdhoqem/MSfUunFo9fAJMBybaLtZsm0kshy2aXhUWogJ
qPGkmFe8KaYvgweoc5gCh+uzEWWnf+jRV9bgM8jmxZ+muU+pQ+EMQY7muLflyC/c
idwdjF+P7yZZxtMmwbc4VY6VoEMNM22g2MN2eNZtqzjXyD3gZXh4yXf1r75/8l3V
yayd7T2aUPUMeuBRU/0byVFcblI1D856/lesoDrdYwGKEN5rM2gufiL/8T2GIO/+
HaxYisnxB3uCMvAFrBxw3OL9YmhtDVk4gpEA86fX6i1Bf6HgDw33++4JbCsRuOGp
z2BlNy54t2yDktcjW2kMcUGIoIgqIOye+gasL5GZcYv2f/AwrD6RxvxCO54VLUzP
nTH2wh3NbS62iUbTW/HSG64WMudIMjybApgfKX0fTUib6QqgtQLsIN/Ia4TMfeAZ
zOhHNeSERmb83deERXPEyFhyjgUdszQ0j0lx4i5Z5E0fdxmnxj3HSv3QuYjFiJtO
2kzVmxrYu1ey9UVEkdlPaZ4gKCoOchLn1ZN2amPMu1S0XrD7hqf2d0MiW4q/ykFE
bPsjYgt0Lq9aj0djWr4FZgK5+JJSqlWgbumGOA93OC1z7j5QZFiIpZL60sEG/cDJ
5f7gcyb1nQNXqdN7owxArn3hs19W5x3P3yIRc9FlrJSSQ6/LY4I+Msnvb2H4Pw5A
e9mPy62p3TgtC9gds2XqQN5dAHFHTcoJaoxTQcwnlYW+BMIQ13+SkZOKDromqOBw
4R5wmks5xH/P2PbbasdOem2Ummvmpo7vBp7hEgKFuSkvISn+r0vCUNWrOoIOP8n1
eqiXVo0pLRXizMCqfz9q2vlFriJd/Z7+VWQ+0SR3rCsZrSqcP4mvDYV3YyhmndMq
UrOFgix35B9iVZIsWF8o/nDpchUc8PqsyDcIi+Y6wTK9A/eTRwHIK53g9gGONDA4
22XhfEs3vo88fD5hkl4uNAsT3Gn27KX3yl4xcsmnUDuX4St2WB7j70ZhERzabvGO
egzBFpKfx5Kd1+amLhEGmHNmmLdMq7AEG/PMtXbiaVImyUS0AmJm4nepSRDtuO8P
PoCstoUTRoGH6BHG6D+My1xQGzYfo27gW/ifV+NTi36IYVYMMF3eJvoCP7hcnMdu
5I7p0waLFM31fZXJsl/8l4rfIN09lTYIW9yhzb8/RdHhyRD0DY7pAOMyYHQy8GFy
XUaoXGtpwiglukMf1yEh3NmR5qeW96naLtQqkApT1k77F1b/QRBEIVmXCeG9+Um8
0m6wY48zl+AAGpb+l3YxrcG4oBYk5f3TBPYqbb08CwZtCUoR5+AIEhR88XAAJGQm
MFXIvAwdtDy1daDBj2yxmPGy5IvejSevuSckaGU7S5CEoF1XGkgCtiHvpPFjOFmD
QpkQib4lFLkvccqXuEF7poQQg/8thQGFz0thwsY7f5ucc7JJ4qHBEhfQ9crsVJV1
tDAidQ7OS45CqyJ2c8OCEao6BDH7nl+W8gF/pYitX+X60UuWAwcHOW8iY0hLDwmc
qDG+MO/eyw74sBAMl+lwhCtoca2c/CbcUVIycKDf5h75Udh4PS7sEa9JYDth7Ap5
RxeMvuEo74zgPCSQAfEGs96Ot5kwQpY5uQ0+s4LJwplQ73neay1CkpZPzMJeZz45
KdwUktlzhtrsGy2rFmTA71tGRSin78ByauqAC+3eWv1bF5hya2npE59CNoFs41RG
sOegX3Lah9AjNYMcyTkzaedNOs8W6i0TimBipAcDVHC+mSDTPVRSLQ0zC3xNu+uQ
cUBeCaMx8y0qnZW51umWW6bCLSinG5uQERSnZ7i4xMHvbgCj7hyVzTfhbMj/puLH
ho/EHo5aSeyMRY71+vXBKNHkvewLukYDZ2LkPZSM42WsPMVGqjmaNroGRzuNkpVE
7n02nLLo/meRqY+ZUBQt6DMyDikF63cDckF0bdao70FHNzXCmByVcbbUKB8O/Xy7
I6iqNlkPSlAJgLPhmRxDylECAxsBYIzCVw6BRpAshITEEjYnL0uGwlVQD+VUpL5W
XXqyU4Jnyqw3V+p4dDMPcAVPpM3ZEGjusG8aIMv3hYag9Pbww7Q9ewunu6sD/jqE
3xbOQVucRX/U2o/Ft7WW5CJ1d8tx872OO+Z+3VdY0uxN+2+qaiy7/lrj3YCkg0AJ
Z1/WfDc6NDAStbm2P/0y6jMlngPGRg8GMZxiEgW9E4mjE1IH5plYLjM6QuBIZC2C
Dua4vn7hGvir2xYk1uxA+g76l/l1XzlIbPzGLQxwLaIywky3zS8X8vACwgwIRYya
iDrdtNGyANfu8iZsTgU2JoG3X2XNMj0h+LzC1yc1uwMCVjHUBHzex6dzUQ1v8ulo
SR/F8j6l39Od5vn4k7WELShrODY7JUo1TrVMvvb17hBUdKf9FB9iqxLFsd6aNktb
lUQ0+j89A24iU5XGpoca16ZyP/eC2cxxTNzNkf4GL0pD7YJJZp2CSD+OkzjErhw5
yrpvrI4AhaUmsdJZ3Td/Z6KB/lQc5H/kBfytNda67TWk30Nz1NhiuOgpThfBYeC2
M4k+xG7UY5aTpoFs6WJVbAZNEg1z7XOxvpUfkiZ8vXIKZBsfZDX8ftO8ouHbkGvo
iPDuvG3GIXcsjv86g06pIiiEt+cbLreBn9WZX+c47ecuafdM5NYhlxDbmQvYUNBD
qlgj3Cd6JP78gLgjKBFl6MqbrbkkNruVxgdKMuKSyBnF54QWQo9zViBMW8TCQGnQ
m9uwg4OPCZXCHzADqNZ5pgnE+d1i1kW6gTYdXIYIRPisjnmJfAzn8K8ugPQ3R2NR
035GZQQVwmA2FqyI/Nzo3xywDOjNSxBfx5RWPtucRbK6aSz+suU/ScZYGbes5FHh
fdkHSMxf8cQFZA/vIjwD4QpHBj6K3qtxdunlDYNjF6E+UdhgHFwqQzpsVZOdbg6r
jylPno0q0MtdMO5guLbCLy3Un4j9k1gYcMxfRxIIzPc+3ycdSK6ktDXqkj24863z
AlRbqZPzhVefkuNzfexklv9jBZvHC2X0ahz/k+GKRn0qXqzoLo/mI8qJjCri4ekp
qpD/F0PTP5UIYg4f5771OuVUW0z1Hheh+OJKrLLugR7qk71T+lIfECjuG175tPES
WoS65bdDaawvNNmD6jNThAxw0+M+QF+qwynf9aoO66tLLIGXAsoFnuZ7sNwTkSlq
V0UXX8LjbI61KTC8x5gTS0z6VnSUkfkYZWIjoL9gaVbupYNMBoGe6eEUcTsCAJxa
yT8i6njBxzJmc0xl+KAx7eJLsZZyn8im2EzNAqrbkC6q6HAQq/Jb3FfbfvUiUNxT
abROYEDJBw0mYPIavpYQd9vWIeIGIggmc6BoRhE/hn5svpP0BcEDRd7fr8e/YMkY
PVzWoxVWtAXrQ/jOnUh4o2NiUPiBISg9Ey9FSvfOo3R//kyaSD/komrYZk2nzHuG
brVJkf/e9pATR84MH4zutUXJL40utjUij1tpDesAmtz1k3bvynLj9HkQ/RLBffG9
1gjZtwR5xbcgEBYxKb4Bm5DT2tqilJnJnU0/XNGeB3V9shWnzCbDyf6wa9q0TN1j
o13Nav6wdWa+bjtWncEOcZ0cNd4nkFlbZDXnbBtSKOGc+UoWcOtwcowb9QHd5R9R
kZ76jExapgH0HEv0P1I5zwhzB/ma9h0csjqBBCYcsAU0d0CiMmb4s1raQoLEXNB1
mZ9YjDanJkXroaKrAS5QTuzEti5/MGJe8xC25RwzXQRnJ31ZM/vKNDytUjn9YVVc
mbnoUAW3n/OixfoaJlvgsE0A/vnnS9zJBN83kE1f66C5vO+r0nJbBc9+53R3S58/
wNkUe6PALpcXp0A9Ohc13jz0JlPgyPzHgogU9+ZnWT5RgMTiIDkEb5OrZOadP6DW
mYvdCkzOEABtYFHF+vbqsNw74cbUDrmtxUtaEbOlsgyeqyD4QcAKWnoZv6J6IAXT
5jrqur9FEKBzXH7oG6S4CNGRqp/BDOy2RI31EIp4CymTC1HTCEfmuB6N0GvECX+t
fnjzxHH/6Lt6ZYkOwd4pG3btZRU3aoyVPc6gjQ/r4mLA2YOzdLSDWyCerfbWVq6E
QOT8AKdWjM6mV7SyEj8eRrcUJmIueqxqBEocf2tbxUiytfI9m+bZKo2nzZOFOwvT
HkcX/zCyCfgTZne+vAGKtM1Yp9WYdasLfsKR6/mSr6ztT5O4l5oz10sSRh1ydl9/
OXJf2CGqZ73Fs51a9Mvp7rdlBz7LCuHVwR5qv/nAt8htiBvn8RzoJQHIWFb1MaCM
mMU0iTenP3LcKj1LAarL/8Nox/l5NoKFN7pqu5cyBoL4Ss4Q+LwMYEMsMwa0GXdu
oH/4lL2PFIAd5p9YMi97pUFDNvVGXw6+bgWhKDhjMfNO2kQMW5l2B2On9c1YaPyp
bcUiSqMBDhfYQGDsSYWj2fTJq+30jJ0unb3hb/ueUjPGfXC49u+bDozrKAn7MGvK
y8XO9GB+uvmFcgjt1JZ/dDISBExs4ZRL7xlW5OA8tUcKiesCd3AZMwNYJn/W1M4I
6hL3j9+bQhyMWHPViq30OJjJh3EhsE7ziE8xtkmOIs+M+Sp3VsKMqVnIZyUTwg8q
FaK5nF996GIUwJFvsLBFsY54HKXYI1EamCuhPHmR/waVDUXNJqTbzx0mnD4DyG25
X6hQzwVD2VOWLkQf+24bnqO4ERIm0nPxTaBeZmaF4JU3zV3F6h4v7VAnR4/ji5Ua
q/OuVgVJApVdTqFoKGEaINcb+FVCG156H3HbcaZKTh6OlRtOvqseRDrHvGxP8LQ3
AJi1sAbVu5kz45CJUMnBzrK8eamYfmvanPsWanX8LRjqB7Wk2SM4mHjzF/lSwz81
PdSTtNylhw7V6Qs1V4LeqKDCc1/VnbmjcX0sScy/UQzooTaS/Uj0RCzMRUmoqfyu
TpmOCjLhw7q+g/2PdVJEjcO/B9OZhSJgfo+i/c6UNmSt471yIzEdQOn1xCJ5zKoq
NRsQSR7iK/tcwiFD0mas4iWLMUGIG+h8b25gN9PM3fsHA3byA22/1PjYVoQuY0z1
qWED9kcDcLxpI86qZ4t8bavYkuU3OFnhhYr2D1fVja/KwL0vhDShVF3jPCy4alHy
Yv0hquj9r93rRDa2GUw7a81hnZ9ggICEd4EtFhdzK+SEoN2fmYrITjGgi8g474tH
02iH/5HI12onhTXSDYk+ug7MAzETZp3mMkfR0BnITXS65DpLjYua5nQqKZNylJTA
O2SQju3lSsdRa+4CIG6BRwB0eyaaIdsB4jkva+6mk0G5dZaotT9xZT3iT3sYyU/D
cfi+sF/AS/6gj8iw8rrwlukAWhP6ZF5u5BYrruqGmCi5UA3r4Y4RxdLgYzxmoJGd
RUa9WHlafx30+pAPwJD3jpWH6bNd9BPIhl4hwLuXsCkGTrrINRIFE2/J2Fm3T6Ht
v6u6M6K8pCnawLuRNtnM9J1/2GXeyL89UYM9xLSBwmcvitUx8RKHSzhRzvJ+fr/v
H+3lQm3s+AVbc8cvkqBoF70Oy1/QsLo7ESm4hk5vlbN2PVC6Ge4hzKMH4Ez3Nmq5
Rp4wrUcVewvU0QJIDN31AUmI4SjYaS0oyb8reDrD32RdJpJiN5Z+lcivzu6+0DEA
RhhWEVuaQPyNvY9ljK4W4tzE7eVoL7vkX3Rp7kvneTGKihubyBl8pCQBbf1OvmHe
SgxuROqZfA/YJcl1clLtpZuxB4uvGwihzr4vMljd4NUWiHtnhhGjxONH8BNbxH4V
CEH1oLrieUyzSvE2G2e/Q6bhkyXeDyONNMbnzyIH8TDXAVQi92/yw7uKTyZfM7jO
gdivJUc/Ev9Wr1iSmOH5tpvhMLitEiEV5+vCyiAnOqdnGPZfg2IHcxhvYO+J/jVe
7JZG+RHPmZ9mirkevDvEunpYH+QPeqrPL7E2sEEPT7srC7zMjkUBQlm+M3pUm0+Y
HwatQuPojEzs9AeexB0jDFf8aZpS5FY+tL1cUd3lWg5G345vETDoOfl16FXm5gtB
XndPpZxmNGbjn9sk5uJ8GU/0wVbLamN+1xsPNCM1ShxvS0Dp7QejZQmUdNadd40X
xFc9RfiwbIEEcKxOpHm+qxfOYvFE1JWKadBryrwjYKu41yAUaNLv2DRXg3aQZ6oe
nr1s/UOjsWfTdYMKxfqoyAXTLaCuNAcKybQz1k15q1n8luPRHIdYmZDASymWu6KD
/4Z7jOdOB8J1gdvCSl/Ro/EYNbAR1ig5yimRch0gbpk4zlza/51hqiZHEHrn8x8f
XdsklXX3EjIpA+wtSYWr3fi9WPXv2c+bOxduIBtNo1sS2Gsk3R/S+C/vR0qexh6Q
YjjTAIVWdDtCFa/ZvF3FCjTe4kGeS212Pkvmph2xBHTNhrZRQPjK9jEJQpLqO8II
IiVZtaVXvKX2Br3FgOuKR9FmpcfjDls2pQ57+vpQfGtzQJGT/r8vTnIL/OcjWiF0
q6kob88AYog7TDOsgB20uU0Bv9jmdSIZzJrPUsdUMAU+cuBVJOVfFP/GOgSPM6rU
XoiCpys5rDdG6BRaViMhsAOv2cLylKhyIqIlqvtdPAgw9+2TTorQuVLr5pByw/YS
jHo3PhncUYZFDMGHy9ZBWVGPYo+Mli7fwBoCHI1QMCRbkPZ9OVc4Oyo6elZdI1K/
5VeEfM4vrNowDJ2FrvGdmliiSCtRQ9tpBcxvntLXA9xIZIrMAq6NT/Q28hbjimZ4
Uz2XwiABXwnQXA++CE6QExDP4AlgV2STsp5Wufsb2fVqTP+zM6a/ttzngcMxQdt+
DQyWXJy8WjqMhQLgqQLKGRuXJ+dzN/35uuY77Gph4izPXYaT6WKXUj5gbS1p7TS3
yo3w5a0TqagWjYOIMpELkPy7TxRTDnxH6rFESLmA08SWQs/lyWWQI/rjkeiCpk88
`protect END_PROTECTED
