`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lVXfOszhxWBsHsgkQ48UEMS+9KyFlnx/S/VSLtYSzg1L65cWtfR8KhVYLzy8CTYY
HdZZB3XVPp1T974VuW52IqA2nTgotUUL/nrAsgVVaBv/4fgCarDwdSzITEof0iT/
6n9R6ZivfgnpGHLzGgWXpEZCveIFHuku0j/XE+OoOYHsD/uTuhgrKWXQo8hk+dEs
jAJ9NVxd33v89Iaeu9BIpCA7sXogkrGfiUcmriaSEnDyzl9oMXMT1qF8zFG2QAQE
/tof0u5QPocRzjZoMMyQS0p+jyT2T+dwhXpLybC0t96o8+P1slgJxL8uPj/uq5gp
G9ji4CfRsWNrDVZmJo2ARUYmFPtJumKBFI3xi/96xn3KPKR84TxN7BkzxQjeJfrP
zCDyMc/g5bsG8+qjnFjP9lXltoTMlELcQ0zg9RcFusz/yLJ4ppN+o/NAYSTzdux+
EO8Dg2yfVtevB81ZzrHdRKQwX5h1gnB1OfF6rcHe1XUD+odIjlDuEWYLrpQEv1Qk
+PNnb9WkAh8Jmvtx7kJZt9Z3zwT0hN/kdfa98kdfbtJG227O2qFSLwafZZqCrw0D
36ZP5Kz3zdmHy5l8sJSfr87maRPxxBg1KM14w0IP5APJGoOQ5YS/prDDEJB5gH2v
xPVxqLitCyP1xU8DrKbEPQpDHpxMKKkX9CnWq3xTgENKEhzYlIK/VQwd2Py5ff+j
kMhnHhJbfwPGH4UvPmZmr2F375/Z/sZOsT0eLYsTcpdi/UzVOS6+7QF3Jt7xFEmU
RCobUN1hczDSchAG3wGlUw==
`protect END_PROTECTED
