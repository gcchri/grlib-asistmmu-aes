`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p+LW+8hxJHuGSzFCht1vA0O7kB6unacdkLXI0TJTiif+T03swPChLrFfGDTge8qg
OVjh8r+MumKPpNsq4+qwz612kTISfBN9DjVV8nuRs8hmM7Kt4RlJpn1+R4qbTwP0
ccbbxyjy9qXkC17HlzYScG541dj3Vr8JksoAEEdzx11fN0W2HMfR2JqM2pN7TuCC
1Y/kwWYnvxHtDez/noe+3KZSE+LYXCW8MHyi9jgwC/4gLzuvbRVEAHhZAfkns52Y
H6S5Rul7Z5VRvkc43yjprfpKoJ0OvQFnZ1svLdfuK0zSCCN5dxwYFC7jGA78hcFf
yunkoasw6Rnk8tdd2CS9XvbtiReiZItTZYrQGcHJOLSGhluEbWJuJhOyDNwHTOVM
yYU2SucH+tQQmt9BkSMbAcfFTaBH3q42/B8k2TkogPb4r71KllLHk5nXQ8BVP16I
MDOotV6ctLaCxzmS2wU3cZf600ezcbQHPWYGQFDWgQqx2ZUoBRgpwIKtAvExsHfN
`protect END_PROTECTED
