`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A6XU0qWbruj9rK2Myg9itiUsNqP1TVu+SKqN9u20SuAdopW/MSU/v/0Vm6rSrkGO
2dwaJ1kCwndbMMkMCmvorvUEh4/M0VaQ4Lvtv9vmdosuYel5H77kqcFtjr77Y5Xe
qZh8A9RcZn2xhcd0zNfW8VmoEQeiWD85NMq/6bhhpml0qcnromwyy3jIgYP/dUOR
dYtyQIYY0WoXLoNf+6sexlNGW/LTnN5Y0ccEBCs9FiKKmTmt4aAMajxHrK+gFZx6
D8mP0ZRPwJzR9I+8f40S09hlzkTIT3pCmEV/p030p1ikOYwLaShcgv5XWTSb5oSb
Tjq2aJVZjRC92+jyoTpHqen2zqd1PjqN+6UZ2k2xdEw54Zt4PKnh5f085wex2lso
1Z69UiQANwjsaXKaFM3OjV4KaGtsCokWgd02vam++Qn3bZH7gOAbgwlxL8NWdKzw
ltmBReg8XRh29VI2rQYhcvXru9k8uf8LdXRRmGFvnvTHFiAOGT+a2YgJFX9UJ0Da
BgVff9iHqG7Vb0ndB9sYX7KyizWhcCE/CvRMNFTsmNqtXIUozOGDHHzQQv+WE+xY
4rTMjciCMsNUD+k1OvVaSUoH/elFqIk7C4tFBzlgS3Nbpx4nOwF627+BBm0ndRFp
U9sV9L9nJWHOU/ANlXp7hqHtyBoLEnUkLbEyLTyf7q82ZUM/sF1GTK2V6riZuyI6
/oqDgcHd2xiD/TJ6UmnSjYvbAbeh2qsiFYMrXQmnfaW9AVOzaR+Rt9e+/HVsTBrd
X/b2gJTymJhfmQUxwa5L4bknlS46Kb3JJo0FV+o7GH2A1Qv2t7UcJ4O/3FXRRpbM
YY/CM2LWh1GEShfQ+M0AxNs/1S0Pap6NnGBQQ/0VkH+Va4Ha2cc96gJdUG9BKLnW
Kq51JYhdvRxbIn/pmhkG0Chtro+f3gMzTnmQ+mxWf5yI1911zau2eIA0APRBqfbT
92bPy9yihSdMCuEUhxuhvMLt5zIZSQ/0G7zopc3r2vAygCI5LdfQP84Z6q9bDQ0e
+53M0VjPFTta4tfJ3yHR0x2rYnJkesMBUHMtYuqfWncUpWPwdSW451An4lYO/cVZ
Dv5vWMHU3rzuIIMZ/2b3UOGJ0JmgC3HWCmz1CyD9QNpVcGqCVUSpLTqotvYg8BlC
8P0D8jT6ZnP3RgM+4aTf8dRmJgKiiJLfuVjkhg99abl7XQYarPDZc9ZBjdK2ZNrh
ybT/gznX5phpOo5JxdVPO7PvcTG354aq4DuUsvfpv1C+wbiMjYSpoa6C1eY/tYRy
m9/S5KwMo2phybcK6KgIp6MCWymmoqsa0QHZqeqauiHU1J3vcEIRi5MhlnNGYIS8
uxykWGmmy7QxyAJMkRFKj9UN5qn+fMn46TsUBLhWeLjpePwta139p0IsjeWjcoRf
X7i/aWY7q3D1mPYVjF/I5eCRpZlgskJPcZl6gqrsufYwFDOrIvBE+D6KBPuLXkLJ
0y9mC6Br0usTqU72ubTYlJb0VHMOqblCar5tvmQDqCbMkV5/bWKU2ewPC33FdlFs
ascVI2C0/3hyUbu1YNqpSBf/dRHTX/KR5Hma1vU7s3fbTfmP5kmcTeHkICmtt5IN
vXgqGeFSyLtXdlf0ldlY7u3jgTYZzS/ONrFszju/hkIaGHrrLFdZVU5H6XKjfcj0
tFVAfIxA++utl0To4WlZttvQ8OSMGOBxA2nJRmEGvuyXRqpOzCjetqNehmSe+XCa
oOPsv5o1G4OA13b0OjmcbKb7cI8KVF518tZI6zZiDqrKWZm9SSZDlGOmeQ8CgIqS
qjA7B/kAujbRhwLyd5dfO3HkJWaAbGLvfxhxhw3fzDh2nKSVx5gDZPlELJSYM3oi
RoAcGQ0PJ7ySt1sMWItldzv+MeHZRyTECOQkBe6f3uYSGOfBsrBpeL2xs+8G3mk6
FuvX3j0sQH/CL8b1xPqNfgrIxA9uQGl4y6Fhvmnx67k8aZ4BW1JzuvZa/q3vw8Yj
cn8fw9aiXS6oC8STCK565b86nFw2d3HfiY23Hck4+m2N3Q5XbSeCUenhMiwXI70F
u0AsVoV1mR/qsxs0skbYQJqeHnhk7hMlDGSDzqnRbCVU92GrUmipboo1ALKk0BY1
hwW/hsVavF1KcczTn4hDj4AY1Mt5qrJcGrTt38BG4KjdHpq2DaBLqeJZiCOx7wUD
G+qr5WPyMQ5Z/s1eBflyiywQ2cp9mrA5xM8SmdgwVr25cqHa1mK3bacjPU/2DmGz
NEOLrohYP99/sMVsCLFMXq5x1QBAYBp3w9pg+pYL1FReCB2EHPW8tHUMf/U1PRDQ
f4c0eWMYQHdmdBp7RpsSL6jxYfbv6574HaWsDkhjUF0UxBl5MxKMBaqsO4wndDLU
JCaLexquCya3DL6/jdKFYzmWjnP3D4J7ArLiVUE+2cYnKTbImaPneJ9MnQJpMbkS
wZSzcWOAZ94AlxgoVGllDN+xH1vIZoZAAYPkg7h0JG7luUi6ux+jmcPsh//Re8L2
tNKkegnO5+ai8UgLkI+oLjYoJfz/314QdPivnAsQJx9LXJd3z4RSYRGwTsM4UZpI
+BlbmEDhLLPoeqBcvllahiVKPSh9nUS9nKptcBmIYX0DlNhrPAZgeN7eim+emw7q
aEN9LqexKcpoJl7aXJ4lubf4ks0Nm1bzgTZBeXkEGSoY7F+Fz3u+q0MipyZJ031M
vMlFRnRnD4Q7hKaBRQSPFDUzX8PlYi8vWSU7w5uruzMUSjS2K7igcWUkymnTi+AP
RI1JjSxHmCB4/0TH4Hp2h05BaT3xFIrqeOEG1JU+FAy650HDawuXLF+t6S8aYcP+
KtSLl1+wEC3+AItJiY9Uj3CYhm5z92GMepx3vpfc8oMwHYFbzfgK2ZaRj3TQjXKQ
CbP/y0J8I6HQffCzW+UN9oNOq99KWQTk2etN3dAEK7NyaiWf6Uv2WbmGrPLGg1KH
gO6/itY5qVK6taIXTdk+SJp/G3ijR9iiJMNGjmEUjvZM/tjfXgvQQRIhKdE5FRL3
8V9GioFEQIeZJ7HcS+QG9FE6ffplcJFcrtVypJvWqKgsSgOYNdW+rWA5Z3g4anY1
ERS53LyT3yUjR6LC7F96bdrV5LT6CVkVtQ/9ZdsN+0yUV5tiFIXA2Aeiu6AGnjpw
XGfCEmMY0mXqnxWNM1SYtzADIXKuZw40BhHI8v/bLAxSC8LZcOuX+ekmIAHELb4k
vmamLLWcQQRlfY978Z11oWQjVMsAwhr9LUG9XVGU282RUR54Z64H9OcmV93+Byeu
YP8QS34k4Q6lHwmBoEgTTEjCAMAqVT7MgNWE1op0v5wUrKJ2+EgbhFeaQwN27oec
9tsGoouG94RbTgPAal+ObsxtzKWhHxHKToyrFX+Ci43sC42V4GEPZD2HVddOl7Fs
VtrFnVWCEe3cyH1yxMFB7gxlXNvpJilF/1ulAMbW1bbdoFJybaOsjHALuaDywlu7
CVhcLirk/Vv+y7VWyai1IScVhjJmwJxf7mP9mDB1lfihn7UbgEzhue0cgs64R47I
B3eGj8mMUJckFYX27aqDM87DwwIPVwPPQjyMRX90yZVT+V11c0jzFb5YhFrIIC20
EZMB929I0/KwTcL3keLxomN4cN4RH0odcAjPyBGj6ZD8g4QB36/I7quJh55oXbRN
WF5wXiegE31lssrVwIV+lKm37w332MNC3Ic3G/RYYAtQMjAezwUUXDwtylmno593
8REsL67slcYqQrRIsJHIuF9J7eX5PKoWOQFZOs8r2QcT7woVDtb8wIWKrhEcOrxx
LFlT+Giem/u9GjJTExk5B0853I36f7cJAbSrVTDqsuHiWrNjWm0W8r1bP7A8Zovm
7J31hxmch16DC91uD58elVJDyCVw0Rmba3zvU+TwPLRIdurfHseMZf33RnsdNF4+
PXXBnsqxUCCYJEu1sWDWcwVNUwhppyVmwafYVMgL/xQ5VoVnXVcCJLdboqbnMdA7
LKfUWcGwb3x23MgIVkuJIOmAw4s2nVHIAOaBJQ2UMRCmq2/7UanTof87BbfM5Zeg
sqU/ibwHd13yqsip2MMuiKzVUHkvc6/ufUWN+bpXzb67DKvuvSj1GEKuIZY/X574
eLb4xM+S7euvo0ls8Ajn1soT95aQXfYBUo4c2AJDWeOv/7z3NWF0bPCsRX+FWrBv
+JFd/6zPmauqPQZ1Z3JB/w0SisjQoU7FROEyXrpkNW4MfWZO3UBhFZ0+eNc530Cp
GL411WWRUQUw3C2hU7IkImYOI1B7r2Bm3LivxDenPq9LMie9R87UdNQ0pJd0ciLr
8peU3MW8iCOdm+CuP1KApLU0ePBWHsZSaKp+KrsbIVTrlvqDGTe2WcuhPaYTRRp2
TJwOVAyaUctczlFZrHsqFunNI0hHOap60pil8BIQhrQ/9hgHCTo4xLuLCmf7IiCV
E3Hk573DSzfypxJ80e1Aaalqg+UI5KBQeaztoM5sKMUCqdTQXbG4/IeIpQhlQeMW
E2Rh7/yj2OZN83+UdhipRXqTVMLzW3DLTE6zDDVSgzaL3AQVIzKyQSO8+5+TSmyC
tKZW7qbWR3NbNjulZc7KBwg8GaAS/BnyQgIMktFZ2YU9kIt4IgdnmdZ0QNC0l2xx
UiEeXHG06nb3VVmYLn4F2nk9B7Mp6423ya40k4dMUESI4ZXiDPygDTmbjKcQnMil
AmJqFiCPEXbLHCEBryCWjZo2/1NoxKUrrPbTs+xVNDjbY1bnEKXLhM231APGZBWe
/Ekf7JFeok9enzNg4ghMxEBxgxq2cNz4H6S+1RI16Tpv+2+bpsIfoNu4fPqn3NL2
oOGoqrrsvNsEqz0rIet31JixDaCPAzKf03qED2aODTExw1DQE++9EdfzSyrTnDET
7ztWaeYrv9qZpRAsaoOcnx/riOI5NcSwulzSHmV4aL2K6Xa1jgHFCdeYuwPt751C
quL/mulgtjToUMYvfn7ZzEDb06huoZck+eidLOw1bSKoaXnwVZng88u0pkNJUXqS
kGgWEXXi12xXScIr/IIUg9iy68y1n8r6qdNGwDPLBpMuBNfZUbJo+uS7wYVovArt
YvzAaiyqYAOLBwrMFvnPldQXMB0UB+VRIO9EwSXXV2k/od87zIqBBKO7j0DLo4LV
Lb6KZoaz5/ipH9AX1RQEy1ahPolhjYbCh/syqdDZToCIT64nBD0oaOmzrfq289eg
j/4+Q2javOKoGzas+FLoBiGIZlecPTb0WSZKPn4egbw1Qm52Mng1YishB6OzmK4/
suuFE2WLi+e0tnQZ/ws0DNN14rJEvd54GIPZh9rU1oBEt9zSmzEv79XrJlkjobk4
DoekpT6oCG4LMkvXsUw1i1Sf7MQIP3v5oqcZ2omJQ2Vqpx9xPeKFEnyO7zd8YMM9
h+Z8qlObFdl/F+/vy0D7HFISlcXlhjk/F99lb8nIbb6kCUgvBEoDxq4w0BTo03Xz
ngL9bEGvDEVudc7PfLktDXJv9Rm1h6XPZalLTOW3pfF3vfTnnmBO5ivK3Cp3Rcus
uwVlzRmqDgY6IQXmKTLDV+I8uIs/9hB9vru9xAtUrXz7Uk5g5nR0Q6Tdp9vTd8ox
BjMvrZDeM9JgXYHm5N01vk373OcJAXa6ht8xR/B4hMNGpYZa+pwWUv8yU7u9+8G2
QYYgCaBXV2O9uGU1uMRmdx6HirqJteasiaWlwHo6DWpWQj3HTHcPhm8BHfP6CNtD
p3YvuGx/weVGq0JnRmQm1CIkVUqMwn73qvgnPNPnEvrhfh54ryqGiQTVtA1PkYnC
QZw2FL6+bum/depConhCyf4377Eym8lT0+U7YKQNxO7zBccxWGYwdiulj5O9E7mZ
oXIsC/9PIDqoTOXL7qlK+jVoMQm1KBFM6ApkLlWBSkDwW+nZxIm2lMP4Yaegka11
11YvVq1pu9hhSKLRjsvQdzuAPXTkxgUd39G9rRrUrY9ZqjOLY/6bl5uAbHkSRskc
fmX2JitR6W4IekGAaFrci3aLxtcEE17aHS2aL+RfHB69PfpbXl/v9QYkwgsQsdia
TPMBIxtpMsBm0yDCA0RARvOpakE6uaGZFAJr30S4S2EeFC0Y2af3hGHMfNDY65w5
rHkA0+kTf1o7p6P+ND+xB+hgrmCNXfiqjRcDxZ+109yfgIyPuLRYlftnklk7iYUc
TYAQywBpt6J7r5Jw+9c0PaiG92zfyHfSLmqvcdHjMy+RWmR8jsrmhjs7E0NxEdyf
C12t/W12ZrD4fwe5tYtIm4JXF6UJ0iNdCiY86BBgfTYyi+ES6oDydZRV9Q6lHKfx
NaAQYbeL9eTGflkl7nig6s+Dyc3HLCJSJCPfsuJNu6pQZ1PQVJS/30Yt1CfdZFno
6zsZS2soIFSMSqGzGGmJAHo1sq6v48IvwRjFRWsGQmPU8Phg6ujjMLoUD+Cqwpcz
+xPnDFLG+GgfGRO2WcMigvwkF40LXG4GoeLaGhYxaR5JUBIf3iUuuMfQv/gZKjfC
KJV1gusZswky3MnzG+8q/qEprWDEMK+D1XaBj4n0i9yFL/5koUWkuRHVVAb9BRtZ
F7gFPGZUUdVZEX3KZh/93iknq1lglzHdAxr98k0RBameGPGVGtVV+t3Kauc/1H8M
ZpAwDhM3Hm92JFUHjfrCi6NUMkYd/Gju3UoXWNmPAwBZL4UMCMaYVd6bAfk97GSG
6iVmDxI8vcVEokhUvqbx4JYkAqJFG+xixuPosjVboncBNAFaASE6uVt4LHXTJ7Xy
EHkSBr5KRthjSInYf+1OxA==
`protect END_PROTECTED
