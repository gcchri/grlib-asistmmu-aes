`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7b9LO4D6SnWqP3upuula4UDSJqHi4XIKCTNpiKocvSxRDT76+qaWCs6d2SMlBCJb
P2IoF0iBJKEsjLEvCI96ChGVUe2gLi0hyPw8vSlIKj+AO5NyyV5Em9Mpqsd5Padn
WxFk+KzmPNrHG3W5shDSWRd6LJKv+3fn/13z5ihDjzjnWD3zYBBxY0Tc9T8RBCxc
b5XL5lU+mWcoJc6A4vRCDJ9XRm0CeOiV+AEeGwryK/Kl0nI668e5i10AxX/HR2Sv
4yJQwCgUCfMxT7a+gSZFR21hZLxyySnzyiuT57Wh+JE=
`protect END_PROTECTED
