`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hqJzwQgAqjYBXmZl80KUo4xAy6Z8vzHkkURDxmnzGDGC3J3+08muxLxMnVm0Ng44
EuhtT2FcDnzeAk2/D13LoJPzAdNpqQgbuyluhiSq/hKy4gzaee57PgncBkty1DrD
fHGQ9isPttaRm720Al6W9TvpZ0gS2hyUuYFU6e66XA+NUnO6fkE5l9X7LXZU4QAq
sYfbZKoQmtKmfi/yKeVHvGgCNuv9rbeJnRgZkHI/E8WqWXJlP+iDRAaRfEx9QG2O
Y3wQqXlhhmYzBClROh85ncPyguiCMWG0SGsq9wFpR2ay7KtnDJk0XMHSdjhcyl4A
RTmQDVXOaVL5IrH+vLr6DB6Z0s/Cdh+fq/FovO9sJxAvWcUNXDa6+MJQ9l/7JZ6M
QaJnd/+Qv+rs2YxJ683ojDE1tvHFPkh2g6fBcTYN16p4/bS3eSoPBUVLeQmYXNyi
Z5eMgf1Uw5UlUCIXFUUnl4CGnb7sRg2XgeO66JF+1SDQvJWzbCR9CfhOk4IEPAiy
fRFJm8PrlezCdnMCxrbCFysLTTYYlxDCrYzm+GD04VXC4fv1sH68TxM4XnAVPFqF
uY0b2yGQp3ggy7UjJXtceKUmla3ABa8M9Jq0Sg0ig5B6cjH9JH9/cHInswSh4i5W
UxNamIxANJ/F4B5ReDmXAEEfdEnmiYvr+71fDBqe9DYwARUfiLAhtgrL9QmFpjsX
aGM5tJeX2z3+Kt8Fi5VTR6m7UwmBD9a21qtqvW7Cyl55KFg6Tp0VwS0ws3ja3eUA
fza/hgIl96xEcOfqgpmu8Rbnnfgv8rObBe6nrCwRJF0lLUelcaxc+WBUKtUN+D/l
YVYZdfRXQcrYfS6Rk8Dm/8HIzCWJPG7+qDxXwjECsB4bc+uxZ9hbOW9BWUFmTGwR
78Ipmu0oYQK0sSlMdIcpQCp58q8LWqBxgzxGFcwDqKU8ho5JURhfE3h3l6nZALcj
9SJts0M5+yENnmHBB/RUnAZjKoXOXXRkIMxiigY9gz8wxPuMjiqehuuxqFgA81sW
jZphIZDtOi4uNyYPBrnabVXNcpgt9O2OpSCQAWXDGqGkqaGe1U6lJW53wpMWIFlQ
sQi+CaJDC1rckbJxraocCSM0OA7iZ6S5HyLfcyBFr/sGftFvG8E+enPAsZQ+J4lX
ilYvmTG0C718vHKenlY6xQrFv1PvLsad1e4laXdC4wVGunOIajBKz3I4l9jtu8cO
2/wNfdUXORkZcPWRQIO0uzWu2Ij+RjAcxs76M+ae7svrU0j4lI5pImYlONx7rfOI
YtFVRbpKXISJcEgFRQaM8GjIf55W57kcPzFZ7YK+ZnNEx5gSY+FuDAX1nxJQEL/L
krZl9SP0TOHg3gFuOMrpSzXchH95goEGiBay0RQmTZKxSjcr/sNMA6fkxpmV/Mkm
Lz+MIl4cXAncUMNKLQ+i61DzXgRIN5mPmJNrUrDo8TE4Hg2DyGTBpPGbNGFlIf50
3cF4y+aiZztQ7bWv7nfBx8CHG1GesuLNEwZifgZoa4OprNZPxusnE9wlA3d0xokO
ljQQbhksfY/DBQOSsghiUbkVWD/enrqztHah4B0C8ie9mxJ6bRPajI6aZb/zIdPC
zqDKKXa4OovbnC6loWCewGt94EgPMsXVTPjr68JYkt/Vli6VdpxMUknIt0gOdIkl
K89PMexLtrHZktzRBWXHoV3VFGWQn2pguogWcyraXeclmetnP5/YsvR20HOoyAM8
dLoVKB3geezyAVbDHKnaOikhqLzy2cRhHu6AFcYePUbN7yYe/1gGckiRQDN01j7+
HPszwvpbhLsuenvXOTM+any5WNmdjmn6t0oa7sgjONsoyIhRGl2pW+PeAG5UhJBP
p5IP43+yRBAcc7L+pa35UpI4MpZqjWuU7ePohkS0K+uwjrzETLX8N1/ekAyX2EH+
kIWvXE+vtYYVV6q4QODkkE+OKQc+KAFKRbrAtOhvQm9bdULpl/EccBFUp2gK6uMA
XrNNYAuJBx7AD31A2weUf93nvbtCdTbfuU4w6lBvNP1uVCH8RmD6GzfXEDbijeT8
tdpwFRQcUWJn3nTNNeB5CyAr70db+52yq0PEKW9yg0WNUX8/j4ld1h36rvxRnViw
y5GThVBUlneSnwivgVVMhGLFeHeBSY1zGJayBUiN8rHHzxEPPij4mcvPvuypxKto
beP/3hfRnMwdZORYFm6bYceYJEyigtiehc2ZlLmZMu+6J8eidQeZxqAexRIKWNJ1
jgCzGk+wfgPVd0SS55uthgQI8plKT30YQh6dAlo/HjeRQsKvaobOsqG8ufrLiCPK
bASYPNYocNsyb0tzfmwGysgehdiILWtvBMAHGgEfkbLv3LKIevqsAT9TkYG6Vgis
NWC7hyWKoNJ5LqJSX6u9YeeH/9Q2tcKrmpe2AuUvxoFC8O35BoEL/+hswflIqSf1
Qo+yTfyIBXc3CdD81p1qbZlqbuF1fAcFMSlWlo+JPwsT3plrwqNGrXZ0plIrpe4I
Nz9lwn2AnP5N/q72WPKBYqcOnDibeNmrzQgQHaOc7fctlaLjjfDRQrohqXW5cvaq
gMykq6d0luluLdQAMz/yj8rTlqYRN2orR5jg4RPTI+OwEjVbOCfM/+JacSjp2F4j
MT9RNuWvI6DY5Xm5x7BcUSd6RRQc3B7X8DAzjoeJB70f4MIF7u5cAriD7PgVUcEV
iAjfJxOj4FlB6CbdCzIxfqGNu4ws/NHhDVugypa5p0vjYoqDdXhqpMxgaX6E+gVM
Aq0DfOBvsrK5DPUDF9OXWwt7dwYyQ1TbmxBpYXS4wg0dcLR/498Z64G+hkih2ffs
qqJv/UN7nSA6lmAM09I+Ng5QMsqiXfYlc0C/6nvk2yOFgMruC5T/8M5iSTpiz1Fz
YDNm5R2OZ6LxAQncYUtWazrpClKs9xLKZ03aD1mMzibMRnbPYEnYhlvIVokrITd7
5FBJpYAp3DHrzo7vf7j3gM5TolJfjSunIIdYgBpE745hNwqkj35bjllCwVpWpQQB
8TpJ+1X5HIKf25JgVGK0nQahmpqXodayvKbwIvegftw5Q1l47nJg6wssfm0rbIyH
4jF1yqFLNxhHjW+kqWYKsM1z1d6dvZXweQ9F4rcJ970dEzfJgKtR384tlglfh0X/
vJuP8lkMlGaQBtIDfW/86FlMOWYOVc3agopeg1gntWLks13gCm45WWvIwkuPV5SL
FBRVRAoTcka4aLr0u/3yRXNLIXaxcHEDaaJa/xfmfEYU0/rmuag/bWehYZby6uWa
UK3f8FPOwL6v2LYJW7/3GBBGMJiNh5VGzvb0ATiOL5i2odhOZVKcTCRZjvO75ETp
+yVWprXnrl8IC3G4i+reHxHq7HQCmTQwgpowsJxX7e4NJIpYuTOE8kscVnrQtRKl
ArCuLZHW8ZesI3/u/U+UJ1sEPEVGEExVjDUHoDRpVY5C1GGOGOOR7EssYaiMsgOo
4PC922eWdVyIdYQdk2qzV/72vXRWek52h5hBVU/0dpow9uS9fvVGXygJnbpcXSua
yeCMBZhwuu3t0vN8YJvDstnmaRT+8Zop1B6RnRSt3/+MTYBdroWEh2GdqCwkrB+Y
yy70imlz16soZCle4wQ6fxXiHJLaHU6MZuB47VcRxtG1UFCeHm+a32W7V3LIdmlT
QnsMjw4lQ7XQu677pQR85Pm9FbdRdhoLOgY6U30ApQc/X3ns6uunGBcUoIDruoyF
MO9+27fgCf+r9W92Fc1uriHPZURlf0KN6GEuviUiOxzpvuUYWk9ljgp7inR0qJvW
8pzUaQxvE4au7vAq9dS91q2iUbuniPqbTSTki5pRKUY/IF/u1NFZbbC2XC3IGc5v
JYcU3Eky6EnivZ1w6nxPQjlo/yakqSMKD7wW8LxMYbcgNujJ4cv8QFKxJjT9GbW8
vYoXV/NJcKS/t2jsCCHtqEaGJJcFuuMUL4TdnXkEJRldMv7dW/yVUN8Oj/o2qnZk
Y6SqGVtYx3Bj2FXKKXbBdGRXjA6QY5+/Met1tQOu1eSU0veI6RZQn0ZaT7b6x8Sp
iJAaiJIIlZfQdJE7zCfCLLwfBVKiDpYFcZZ5QORaJKUo3+lOHmsiqu1LFv29z8gD
mthveQCLIVIxj7V8N1c/yEQhWztrAuN7gIXhvc+FFOFCrXPosy1wtbPDKSD502Fu
hXLi0zBNrhKEuS+jFnuSnGnDseQkFjQkkQrxsNBSsM+Ibb4QZkkyrp0S5SN+YqjA
JJi6WFe4mJlDoP4ZM9sTAHcxhVVLxyC7WlfMC/eIqtdWBfIvqgl50wVP3p6GuY3F
Q5AwJbU/G6zRsSmsp7yxd+yj9nte/MxIS0Dfi22wvnENoILjSgSWvz3qZHisgrbD
/eA7VV6frDqxmwXFlak8fE9D+InyrAL8twMM4/gV+rz49ppHLkRB+XXxlpi10xJH
b4E3FmceBkZxNgPi8Pf3ARKLChA76DxR1Vit/GiRYbD8j4tG5BOpv1bxT6uGtQJU
5m2ew/P/w3k0UeqoIcFzSSZz1mMOMdwry+JqwYniMv2sFM9Wo//3HOsVgqQair+n
scN/qm6AapqVNMPSOXoF6gNT2ogGHf5c9V3oN5SKsY10FSaqAXlEB1aLcuznnCz9
zKIYMo7ZT1NbYs2cx8exRBkS6OEpe+0DkERLdm2VjF+oKUwaBPqT80XqtUexcb8H
iRwRVhpNQTiiHpLUUBm5L4MDey++cTy/WCmeBP+0FYFUr/0F2zEca4npzVs68x2d
P6VujXLds+N2q1SwkKIP/4c7dL3NTPu0MFPgwySuZcn2Jd9+tWb0o1cp+SdmUi7w
lrnCKH4H+fDOTQWzwsA9UzmdN03UnM92qoo6aGkHJqmspyvpXuC7MZl82QIBQjU2
0nKRYbmhDFuUi9gvRbJOmxLSnFi98fGQuHRvl5OxngJqwSOKuK+QMS+fkE9jVJ6f
WftwYTUgvm3PaKGgbmltbmyXVNY5kxgfUlKH+WVLSTS/DgLJUNnx4NsMuTMXr4GJ
imYXNPT3stEBryV38kXxf+IeOKjxlTIQIVqw3HhehnWFVRTkeYJw6FbCq5ddMa30
homwjOyLlFb0iPs1B8X7PmuS8JpkZDGs1wVM4iQN6IS08XGalXa1fBJNuuzzcjNN
THehESHlUMvrByL5ZGjk+7eYrua9ndEA0y1KfYIcba7NgUMcOQSHT0h63OUKCwCE
0ztD943tAsCRgDZlIn6O6iOoAGi2YqgoJZNeGA8E+skwmkB4cOTHJyDdQ0DwDxLx
XQEPJvOA9aCcf+Xda+zdutq3eApjz5kQYMDXjQJ8fdiIy0xa2HsyDTKDiRhnkBbf
PObgIvdjqkeXGblOYm0O43AD2hmv3Fr0yxXU45Lp1+Y9J/w6cEdxF3hBQL1VVpJM
dkuqeQT5melwkstNv5uSCXedM8NK2ufFnjA90XiQzDw+ax18006BLPPBdhiM4Uwn
IFhSxjlwwk23jHmC/KH7lIoh0AlLimSCG7p9/6d/HLeRV4I0QPa93kLCnbTqcUzU
vIJc6c69QZOIje/1WjwJ/3OI23HSLqHa1fBnzohoMNtKqYzOBgLZFf6UQX6no33z
fYDVE3dNOWbVh1dgYU4qr7fFM/csxAD1EZJn1OveUmln5+yIIyOwsBA3vzjIxg5j
YPNW9Tv9X6tQDBcTls9PT9Or4BZeQTtT04nJ07P5hPWT7tgLscJ55ePhxzquMPO6
zCUHTU76ZDr3X9VuQ9m17l5W3YVJ3/+ZRVWlK73iDn5pOr2RIvezQK0Ua4HHqeCc
iNXcoZwVfVaO4aXh7UobZNd13zW9UHaVGvZx+WUmbRng2gOjNyaNan4TvFbPvBo7
cF2BxbVTkw983GxOv7QlvWcCBqJ40tCFrUMojpGxjRqAjZL3NMSGiocHja7V/DjI
eLKCD3F74/Hg5qPwKF/qohENCZJpTfUVMk/raHJ3w4Joext9ZZaWcsCqE9sYVTxg
ZORzOZgyArW257bJtrqZdFSi7YpcD0+0gMWzCK38hjPce8cZxdjy3MDsBCqJ2zMk
rIhaj80zCZH40HRqcwMXoGkZP+CGu1jMHaGtGccgrDUqWWqJ0A5uueyDALQ6V3o1
/jXPWaR5fzhtApoWcjxHFLiVrqcj12bK3lQFypzlpF61zBW7f17B9TwUwEv8pTwe
dCtQ2BRELKC1Vo7sUQ6OHIdEyaQVSGRMO7d/1MA4vgWxTFa0n4ZoBdWau96vI1OO
n0Xyab+OzlXKu70WvyXmFgGkvZeFT+ExJM3INBtZlIXq5jWTUjjKqInekORC8fbc
Bkhw1HjggIB8YhPfPZqDyvvcnnQndhgphopFnVU9BIdJkt2qoZUzvz4lGDWihuJl
tIIrf6e23DMXyATI9T6NcVd2qsvFTiFQtW9GMOklEMuWW0Y3D9Bmemdg0AmGz5V9
WS3msPyQxeP18/ZaBQ67kIpihW9WY9go9Yjcdsvc23DdxETbG98se6yp0F2j4+/9
yfF1u13xXFeEeXJ5mFrCn35StmGYChk92yCEGMzgWwgDOZ0IfXN7Ni/i/St9rf01
Pcx+D+kOU6zU5goII4nsMjCvnBBr5zogmZEbY3SPgVx8kMlBtp49EwD53gt6lNX8
c1/UMVEdvYNB0oM1/nm8mhmcmQPhCjl5phoCn0CxK1MhB8fgiHeedz6NOa96Fris
GOYOFwysAz/8UHbHTNSp51CSHl6fmg7IJfYTsAm5lYgI2yD1BVgXyt1YVfre89Wt
MLVIRHaTHhiHNKJCxYQwzqNt7n5m/01TgOhi7diHcZit5USTDc5DfpkHB7Gcg4yr
bcyzJ+/mF8xjgAiuOmf9O1TLyr3+60q3G35k4Ao/gJiuyh3bD2C7JE65fip+Yzzt
FDyPpFFiPx44Iymnn3RdXw0cPmLjpmWongPC1gTGhSDyCGNR0CA6P8LsGjkZmu6+
zL+q4ebUMSfGAR5z9UNPcGJlfynUXKeFH8s/c69SuCkUbJEVEmgTCLzpi7mdG4aY
v3BWSImZ0Xv3nMZdkonGxE6vjRO2w9vt0GzuwlDxTrh4RsC9WiR7MbtDhS1XJQSG
RX1yj9IGNImyttRBHpBBXDoTyvhDIJxKV2xr8cakySB5+S5N0xeG3KY/UYj3jGVU
2zsMr/A9dR+7cesc2mSTbH2v1ViDcZ8s00hDP9vQyPDaLY/80p3FKALe5+lkJXGS
C4bWtL9ykcH19D/X0f1aGXWpVPbhMuV6fGbaU26uLmwX7tmkMJMLoD2Cr0jMyj4t
muLuNKwOnris2q7R2nkUB6eNkCkV6EnZqhW39SUeX+RuZz3eEqrdzBZDX4LdHDCt
c4pYSfhd66WQ2+04TBmHI/ji6gQwa+Uq6ruKyYQ8RdM6QH45ICH5co+1iKDQppLV
tRYPXDoT/5dzvnVUdkiG75uVDQNiyiXu0nb4TSKonJehFsZuorX8IENkv4yKQ3tx
r1HvEy9sl5SW5MhmFlhJt3PZcKLrVxtvkgBx3v1awhp9DXRG9YKnanmSChrjUwXJ
KOuO9kyZS9cJJCXpJjcBNj2VnteBV9nGhXs1ywWtGb5cTC8zaZyNhfIeQEqvOeal
BALpEpPGOYyx++dEidA6Aek5LpYFvq0sauprdHajGXWgU1QOOYs6cqfiutjPDPRG
gcVR0hnOK+NxHbOs0i470JHF6XywQfsnwdUgoIRBfj9WO2OXFhYHM+77yCekRPEQ
3BpKhsACqLkSbR7Zc2Mo3MitnpRNmXPYcYo0U4QGlw5SePueIPwGdnHWvqSxbImO
RzbjfPUQjuWMRhmlG2CK76CfoKod8gqdP+B37Up9QNk23/ad1cmJWE9HX1ABs9gk
52Pey+2pS+Ts7MXpRdScDK0wUsjlWGmnTHp3YYRoaWclHdhpVL/g0UR0BC1jEVsO
VJrjo53bSm1SVZdN/9mrKECEz+fMOKtf4kZP0A2Xs1LEHU8ZFasGyl7lP9dsceos
9ziskSKqmG+CtVnhL2ggpAHvJEhxgsEzAYnOcXATnP4xSTLxoN/PYNt3JLduT1Wf
Fba0VR8018xZs+3aB7QIcswhfesCcQSKA2UIyoe0XKQFj7YlBRab1tD/ggFaSOpy
t8IlCfpjOns7yQGwJyJrgwGDBlk33qfPvBachP947QU2CtCzNmF8BsuUIu5SNqn/
7TIV5DCxUOrLuuPcockUrCTFUXhRNzLr2Xyxwc94R3wtKhfWlultV67cZ1eGBGL/
Zv5xgFDU79LmTpqQ4hF9NQtUhXb5XeFFeQUscGw0VjQks+UNHmLaWlGqufbndmE1
6Ap916kAmfEB9GStUrWBlWTUcAEkiDfayb6yO8hEvh3dISBkqY4tB7lm9tmydU0a
f94b/Bq3PGT6GgRPjrh2gzFbGlKJZqnllRIyG53RJvxHGrXC0w3IWmxaE9cRLxUw
3e0mlZYZkV/N0rlrRs7cd5p8wJR90S7xAWDN1eEl2L/Q5aGWEymr9tTOm+sJ2O6x
qNV6o3JKQnTQ7f0nLZREeskpwCaDTM5zCkzSgtrId9OKziUQT5R1khRbOuS0nj7V
k9NuVV7utbOmPtSoUMTJ/lDRBlWeKCLnU2cdh3ZGsGyt667NvbnaPPUjaen0rjVH
LmNfAmgIzgvcjeuvI++ZceBPm9qFV2/BF8obxlytBYCNgF2sr7cvf7iaBjq0zDEf
sXct23fv3vzh0WR15Mm2tWDX6rSxa3/bCJ5GH19XUerf/WHBmAVgQYpPmfwDlzaR
z2A5azK/X5x6AEUXwgh8j3Nd2XaW3hTRBB86BLTKJY7r6UMT7hiNM8wi4vop25fo
jy6lvIOxfO8+P5v6ZSHPBPbYbBdPgCgB2kRz5FrW7qqkSj/6oQVq5rs/Zws0y6ty
KhKZebumV2ZMoKF/eaqOu83A/Zaj5BATmtYgafiSkWV5pEWRseYJxHYkA80YNj3G
lX6CKQ7nMlE6PEYY0CEDAPmQQyWcfkzPlLBl7Y8eIG9XnX6Sziz5iSg3hEL9JZjJ
VAPe0tuW+2rDBYmjZ9HRAnJLj7cazk7LC5eekJcBGajcYKDaW0Lc41k+0lXwQB55
KVl7E/fN8h88j3rxoVTJv0aflvq8ej1pFmNRp3nwHTHCPQOMGrbN4yoA/CanlxF4
Bmehdwr6ifjHyB8IFOCP8AITbmMp2um3sgiJpo9F6DrAJHRbu3f+qKuLLx4ynuVV
jwubNdBQY7XTFnKk4+k+s+AGt3Sd3ayQw9jpJlHtLVZVmBgKDcU1/qzz8nIjgBVu
2C/1ZJE5Pl65DK7lXJhbjjpEwrRTMgw0VtbtCNa0I+hhDBQGGOtKLvAq1ApeTf8S
KHi4CdfE8MSDjUlCJd64XgRJx42x6W1qm7c7Nfz4/LnwP1/RmWoOyeqtYp0aKVhL
gQXwj/hDBlg/6UU2HTl5+q9iRwfbVjbX2puqN3yD/lhPU5d+WnwQR83gXQmY/I4P
Z3IDWdyLC4ryTgfaIzzX20KsCn84Azxo/qFEjblLRCvESo0NPz/vY8EQhKe+pOlj
vLYNz8g8ZY0go2LGzqk9kGuwAzjDr3gzzZjdYOPoapu2McSuGJAtvVl438WOVGbs
AA103XU4os90e95FGf3tlfMDBN7P23UUGTElYnH0jqzTxF9eWvHKD+Z3EL3MadNv
yBZ76Y2h9D1TTAYJcvWS/xgb+sxm/lWZ+RleeyrIVsUe7x/linWf8tfitDnmgWy2
m/dPXv5P2mn2nrUTT4AzxNAAqHg7bk+Fn+ISs0I8Xu8UkY5M0xdjUAQ2fhNzSrvA
X7VvIQkR9U6I78x2TQeFBnByK9mX/QWNhwLI53CT6KXKPK9GY8CRKvIeaXGnt09v
K6JDvI1mrgCIBXnaO4dH92XwVGTiMelp3F5mgI8WsBsAYqP/7wCe1n9Q8dPjuY5E
354WY0M+n9wXsZaZoDWJjz7F2YEXMA2KTwCDEBfADnoM+49hy+uFLaEQgZJ79nUu
C5yKRfZnid2skf5FhtirbuwCA22pvtunEbp5bs20/MEa0yUMxv5fO7cEYwmV80Hc
l0/pbDRhXOFA2WHi9DTfE/jyJZl1Xd797Xm7QdC8hu7mGtz1cBO7dJLHI/8nIx3F
K/LsM+dVVHwCWMa7QyCUIVVvDber1+nvEuati3Kl9TXinpbX2q1/HK4OFAR1tDHR
+dFdd2x06XE9/PAR6t7ptmZSjpELiAyxyB74xH5VMx/6VL+X48NtWGQqVa64Z+gk
ghaA/pG3aOoO2PnofX5GqP/6/6zZ061rSYIVprGmVSXB+dPDMMYGSB+gjl6KkFKd
mwHrj44U2E0eTWM9SaXgK+UZiLrSlxGDwmoa9mJtmmI0h4n/PW5IFTBdnvUESWSz
BvcNOYL6hEWLiHU9FYb0rS5zH3pzvq1jAiTVv2SEcW9n8T3vmCZXiXidP8e59ACp
JbdL64XyAo839gc+kYPQolIWQnNTGLX/d6DeW06FFh69iI4fZbl0SuMttdSeWTBv
5mkDeLPan2h3sZENW0ibQTWVYY2N0KIfFbN/P/75FeQxlI04S6nT5AZNA4pso9mJ
FpBS+iTu23RjfQDCMFlZUKiRLWN6lnFFy8XbZuEqVrriW+ND9muJGtHRo+hDxJok
TdVov3mwyq1Hv/+M0y+2fQZDZZI/NCLboXMHaoG1OTBtCJRJ24FJXn7brzqSoxsM
Oh583muWNlIlFGzAaSVBnSSDvnKPAAyY6JvjnU6KsPCYpepB5L463o60duRyncs2
5ex9lXIBjYv7a5AoTkigEsO392u/vBQPw6xq34LkYy/oeh+V/4UfKNLG7jz2MscN
78S5CDoaLXrcbbV3mTo/2nVT1nWqe11Hhr7lHeBfVIilK5AtUr6zSDxDkgZCLCMz
D9xLHwsCemzox1CqC9ldGI+LDOzTbtib+YLgdrNjil+PqiybcdsyXWWQc2l5VyFu
GcJl+pZAJOIjCNN5kI38D/TWlchs7L846uB+DIupvkgTeKOorZQKLhTOUuhg1SHI
4iH5KmYHuvQsa4h3ypUBOjhl9izePr8s62zJ8/7f5ywElO8KMbLQ6G9mp5g9uDQc
PywQhCJ5cQDeSm5WLNnfiXqbuk4Cl6g9GV38FcHgtwnDGUWP+cXragHG6npbKB8A
ACaZcdrNTkySpI3qPZZlQw==
`protect END_PROTECTED
