`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mDMam9svpcXwCLR04dh1JSPozG3pI2HOyPVkWVhZ9hIkBjdqkuT1C8ORBa/yWpYR
R6dJwgnxMDphYemIWAKcgS3XRuxoU23iL1/tdeELW9JW/r/UbPZGD7c0DreRkW6t
7+qoVT2NQDzXxRVY9vly31P57J5zXFc/Zblh/QOTwPHJ4Opu4qmYCQqUgwE6vwWe
H9ZeYMUfO87BW+8kDz+1qxF0ziysvou56sIkFo0aZ6OZxDGNZ2pvcjneZxUycpg2
PYAoh+E44YFPAP+9AGjC2/52KF1gZ+UzPP+eZ4ilkSsiqR/USRhaCEKiKmb4TXqU
`protect END_PROTECTED
