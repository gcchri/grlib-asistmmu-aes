`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/M0M/mnrz+lakMNcFhz0UAbtRc/BilEmeBWKxizlxw8P8mIII+H1lRu0pmWM36Um
9NVI7T/sb0cH4W9KXHqLG/OpN3WMBf+UxhPw4l5Heom0R3xsHtQW13qI9SSQbfX7
6BLBagw3Dm/CONCdcoTreZPwpWayz12yQi79Z4Xp1YckAtCvZmiaWXaYgjRPSvis
xoJhw4F04PMSxtoFnKZagSeVDrsaADyAANOASLwqug1mVBlgpnhAOHy4uSM36ab8
C6C4AJJ94O5kN0xFWSqwIm4jNPsWpoNh/X9Fz79sGX1oJVbF56yH4mcvUJuEv5Z2
5Q4qWkNgga9fj/tqGNxayAoQ8kxsUUzmKl8EwYQrIq8QpSZNtaeTuTCupU7CxjIN
2qs4wBjSSnjkaFs43n1+5a8JXh85nxYVzolrRHjKjiEKmEJqVhO5WkQ/ick3wXIw
`protect END_PROTECTED
