`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AjDLd+kUdCiITi1boUer7M2z+cjDCaSH9qjLPGkm+eZJBcqlqjQZ2sg9XJLbIn5Q
9KF9P/uh+qCHmn/IRDyc4afoSHJrKMwWAmxTKxugno2yc3vMdmkGyKeHZqToHrox
4SWE/UMO7xnFqHj0NpsslvqNiQ7DdmG049rifIdsz1z84V9IT/oNuCJVbm5efGu4
rnl0z42L0650G7VnCBoAiCcvlBz7SOkvgsDFNEWAZ9qbCil5hCgg7Q2vXjAEPx8j
9Rpa+e7B/n1P7GCq4h4X9LTTlUYSjjTmeJ7OeF4cDD8UiLylzi+JBzd5jAxjdqrH
EGohRWGw4ezzLwUv5RZ2htLwmOImMLf0rHlA9Fe241bs4UGQq/L9WPqR4rjQrL90
T2XtPfNMTXCA9dDCJJjxMW8ETzIbxjoYuzuCNnubbuF5Y6GAFMLc8PKRE7PLrFib
YnzGa+sufEm8sAHCXl68Hn2NYpvwJY3Bh5iDzIKpta7CSs/mSQCi5SNjsbqzbCa9
p4fm1ZoUj1Cig1VLBCpDXo4/jB28OvhMZZijoWGZ2RTfyQ/rXTrBDF5rs8AVmjGX
`protect END_PROTECTED
