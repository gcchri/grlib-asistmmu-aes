`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vqQlNdD+hjyDBA3KzKuPG9yewUobt88jiokcitOd1a/Hs7bUWhPc/ViyO+V99ZB/
GfH5125glo4DgDh+GzfqQ38V8j4EUwLCW3Tcv3iAN8/NA5vxxL4HOgpJntjJPjEy
B7MnoVJO/0P6RLJx+bqKjXdBoOFZqUrvXZ77FaG2m3/M7g58bBt8XgUanhcO7Q/0
OEi2rr4d/fQyFby2AYKuA44JsXnwNYZdXhOZSA0yWjvz7XbY/7PI0cCBvwBNwLeN
n+iIilSTqyy0Px29XJsXFsJhhM2EAKx5VX3Sr85CUkM=
`protect END_PROTECTED
