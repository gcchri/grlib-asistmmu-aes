`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VK11zDljPfisnGCytNoLQ+8l4QtUP45kNe1mGTpFm7FVjYBPS/ljl0CSzo441vrn
iWts3f+rRXA7idQgJ0lOlgkqZ23MXVgp1TslNN4uU8YCWUCqcpId/BrCwMG2xv8t
NLkY4VTPj0uNVckmTpJ263K0fHeJbVg7YINdqTlj/S2MoQJmV/cil03egP/pJ8he
KHcy/uBdatq3NrORqbyZx4prAP+9SIlp9VPIBW+15iWXzXlj7SQkforG/9EGUU9I
SqSFv0J1rrPZ7EzehZ0COhNs/oxbJiUhN6kPeecw5CPoloIIZfM7NHXIjeUZsg7E
gMh+S3Ypv7KtTI0rhJcdbNFLiY5opbbdEsnpz0YXYKu9IKvUVb1j+9DGKghy9dIx
5H6HtI9hgB/ejkkxitJuu/e8l48rPWHk/EiBn7hYRSiGvY2Wgd83uzrMkwBA6xl3
gFifFlUubWkzzAVsCKiZBXpzUE2/lPfVxj4XFCLfc5ZJAJUlyKS4lg4FCDD+IwEb
QPauCsEqiua+Sd6wkDZe5o/4AslCgCVsPe77aZa0yU7vG/DYrS5dKxkApe1CPmti
7Yb6Cxhh5Xk5PIQ7KZriPTQwutXP4Uvz9uiYdo9DOzfGBXPqEF7D0Cv3miQHVNyQ
pjbC7r4fjrJboR4y9o+ymmhQsydpqN6m949ArdPvPzbQD4IsMhO4LI2s5ir6IDn8
R5hijF35Sedkm43Y2mLV3uD4KMPcUylfxBH4hdYOJyri/KjmQUDhxan4Dec42sTg
4wZfSUhLoRTgApzAAq78fiDDOQCpZWKp4nWVTOqSj/zfX5VTj7GktwrGx1bDyOKB
kJaQrSWBvOrq87r9ToG9NuVtgkiIuyXogqEFIsy19ZAoVv/PX+ZXtBlW5lmpPjW/
SGWdeMMbi2WeyuOBOZ68LOYANEn6f2m+oKOINwoCJR/U23dUwzasHwGhxXFuPRKc
0q7czHMiSaA8I3qdlaU1jqJ6ly+n51bRxO6URCYsHcJPTxgOheY1ZAVVjfmMAJeP
zkJcX1i4aZ/uP7/NeO92VbG2+nyKs6NBwkVd94tGJ8EYMIzBlBhqjxVxRIvGHO78
Yk8IA94uLFFaH7pdSGPR0hq2YgRSo2mb05afUES4Jspx1YgTszGgR662ck1cvY9l
RnvGcgn1Uw3/Y1izkqn4Zx0dc74GFg6guc4g9vZ8IQuxlJ6G1iwiEg6F2H6ahajB
Uf8259UsaCa6poPZWxPHy6/vmGZfZiq1hRSKvOaDzZDFQnUH2Jvhjry2gZxNVIJu
9Xn5PV01XEWbeDvH9VKsOEL+T5psB2b8zY0ZtGgwGgLinGmYqE2QPsdgfupvkLWK
a5GuQy75/JzJ5Xp/p1lEmxGyHH6zX7MQyoVa3wEjRt7Xz6o4bEYzFAPqd7LN6cD5
xFlhs2aScyyUNP6BcODRZgRJgu0E9tlWChsDykuskTsWpLDQgNxsyG7tOC8urfKr
Vv3EPPZSrskVAOf7djHoy/S0qLLyS1kviMGD2E/Ew3kp2Mz7xNVizFMnajKAE8o4
3uz1J9Hq4J2NYH681rEh2AHD4Pf1I4OnoqB1P6i/ayp+5NMLW9DNCfS/z8amnanK
1ajujN6eDOKCtnwUn65xDiJPXPQntZq/KZBH+PJ+QZPjYfhEasFe+ukowZ16yYO2
79glQ4kGyuItubBZoWeXj4lTPiM2GLe+n5LmSav6/PJTBHhX5a1xp7x56SQ7KIB5
Bh6gQwL/9r1x3YT50WgUzoLsaAvn2QfFbZB+2oQwIAOyO7rUTWI/PAddbpA4dyQb
4xHvOQdYWIlC6bhm6DQw81yKGRJ1LIccjqDDTbfZLWuSiEnmF0N1GtB8xC10cPDK
xJLpxkdMYwV52BgvnnCmy8VxTobjhbPIqiVyuuuSf74ARQoRhtsl0/gW1F9Fboqc
J0x/Rvdmn9CYff716NSjaE1CH0JfaKe2dtOQ74+3b30DHHv2gHExD39UulLM0E2p
RW0H3aCIc0AZnFEe5o7dW20dWhu3oV5oZ2PmxYumYpWzS3n902oDXGJ80gRecZ6E
P4yxNEjNXLWCm4ASLtUQ5dhDu8IClEXLq6H2Zo7Jwr5itDqGYIH1CTvDfkncq7Zr
FuleGCIzKy7944sOJPeOnnbh0TCGxCwOjWry/BJjY/Oe5C7jdLpwJe0TLQQ7WSDF
WG9M2G4z0Z3R+JBXFQNm6F50iA141ZZtKHvqckLQLfnWKKAPWa+KiKMe4UT7m0FX
JReK/7NNJ3Y2bZwdVwfubDOzvFHmhF8YUIVF9j71in13d4/la8y9bOr1r9OuD3c8
y8jxZWlVIBCK20OkW1Vr21yI2DpVbpKBhpWBKsIBUn/c7lJL+2a1E/uOm6mAUyxF
2S0uKkfPHzUCTjD+DwplyWhVxE6oVVUU7yF6v1xpxtr47FKzh2Qq6ZLtA2+G9VfJ
s2nuf7bJ0x+291blDTUdZpE/qYhR+mPJ1IipTo9lxb5KWMh1phZNdOxyq+KCVy2V
3oL9s4+mOBNtupo/EyjL1xzm7Bogex/ZPqUxGeUVEXN9u9Wfb0pHJ/xYbncaENm2
UAaLfikgfZdkgDrfEEhcNp4kliiF/DM29kF5me0Nf/kd8VW6gZcWXTDlq3TaJlPY
HILruK6GEjbAQtyy/oiKbRCnZ8acSF8sdwoPMIIetxs8uF3pZnKO1bSJa+djfwoW
cfnx0wmvuuZBsHJo9TiK2aeagjnMQswMjucw/Rtx3XeYwE3AFsF9NEPu3wWuAat9
SQa9jezlyjcKP0eTOcRBFid6l7drYb1DX6uBtk2eVi8c1WqirQ/PVk5OdpztRVia
mp7b1GjuDhSC/bqJajKdqvkkjIJ5G24+67LOKWQYmY9gTUwofSXdqARxW8hnzIbX
zT4DvWf9b3gdWk/VxTQrGkXzXBIyQvex1lsmJPVZb+hwbiQXXkhX1iOZiWNm8Ty4
aVpHyH0bGS3cqFntzeCqT0XJFfcXx09I/XlRvVCG8xwUeJYz9/+XNYg5mfYf26Ey
iDGLn+w9OWNNlxn5/2r9HolleUyKv6973N+KsSvY47Bc9H7wlGDe6WxtTGbyyocH
lzuU6dprXAOBCDu9xyN/O29iLbCXdLbkyvNLGFbUW8uNnXXYfWmrSvqNYmREhKFk
9IeHmmPT5Xz5iKYVosmG9SBMuyjSYzGirq67j0gzbASBQMHKb5FH0ly1AZnBksI+
tIqLGDYxjN3OZfBCF+jifyGBF5ZiGyOdXRoR9v11aCvvKH4Nme3ExOxFLQcwwGUh
sw3RRodpZszs+AXZzV4+6WKtnVSlSpHkJMM9236OIPvcs+jSCUOXA96Ine/lyDR0
L1H+wmRB0kuel/q7PoCeJFruf/kkgb5NNrZgu/CRE4oplA/wIQzkxPqfdsNfvnDf
aiyx4S2Akvs20oO/Qhj8ZxUxcqO1/Qc0LLRPM2RaEdTCm8A60AOdhAhEONoJFaQT
qEgQTBza8q/hOT9U/lnpA59NiX05ThmXwvGFmBkyu0eh3Wl+AAGs50VBqt3bn9EX
T2MUO1cJpSbkvn1HRBLukX8TVVYON4obuI/HLokq2JYs4HAWMtXeo9Zv2JvtDImi
O9MxWXDiFLxiBCDGyTTpzMAINLnQ4mJR/dci7ULX5q0D/qksO4WiDlIAWoNdmY1X
g68+my4BjeCwQwxXZ76m3hjsPCu0U3j/w+IQmiOlRa+pE8MpzYW2LGaU5ocbnWAg
HmSlaJTlFMRHOB+gOqXMCEJAhThtVKaAV0kAbtrgJJsWSOrKVZyFXJ1fAMa7mwrE
bHsJSUG8yPboBtnlrAi1KjxNeHzdcdgSqMyOrOLFOwPVFMlVbZJHWYaYzrgcOcbs
OtjTIXR0ugzEcFzar8I1My5FG73bajzvDuhyuFpPLZiyKz1D1CAdqwzLCplj3iVg
4fn8kTKnbSijddg5QdEoMn98jMcd9B/GXoRXhfaBVeA16hbi7Xpbu4rOs5zDFOuL
VZGnvtItZ7YRgGMLn9Rhk5/KAaKCRcGryVBw6L9I4OgdZb6RPvndDRGdiKXrnm82
k3E8QHWmW4SZUynQvVFDZGUi1GHQN88gO+Cw6MgTxqZz5msIBWA755z5g1cmtrIu
G8sH2lzwBPN8ZSx0Bi5cDUS4I+mGfX307yekA58Oco7IPHzVW2c8Sjifdz3N/bDn
KtcWjFng7Yrs8pmtt87HUB8sK86Ls/xh1dq4SREeHNtBBWqioByBNfc1cW8thAeG
FZ6wi+K6zUrpqUdmRtlk+PB/dZWXhfu1j7YEcjZ2anvY6A5Bb7gFkTla+YA+5SFA
g9wA911x3a/DeW0q5O1Ha23uO+A5FHpdErTqFzVYsiCw3FsdRrE1SEu5RG29AdJw
h6Vosq3e4fTWRcUBvqZ82s0Zk+NfNgf0J8tAzYM/VaFRWFNVIZPB2h3ZeL20nFRN
3l4o2Ecl9uj/XLWQA2zFW+WyBhG/HtLcm259YvlYOekPmYCnL7DMoZLVJEY5UvxQ
altBLuOuYTt9PtUTv5mfXwT3OyUIoZfRIfxEXE+Imt/PnL1JvofIEXsCiDRSEzQG
XfqnPvssrLndbLz4OSfy+pFFB4RdJCs+AZ+o5s60SNKv1E7A5U2PTKilZEDaovaw
DAjB+EdiAeqRRnHfpuypS15Z9jxlD1u0MjF1CgrNwMjUFiTU/SwWV0oSmD0jTM/4
3JyR5Caudn66Fy6ENdAxRyL7ThNPd3Z6SEYIdJGv3LVNYcca1KNzsXPw2mAKpnYX
x7RqgBHcgWjGz60UmkMb6b7ZRuJHfwqr+9C2cwOW3yNgL/M7dsOpGcWnUsFmXah2
xZIOXMmrfT9gL20lP2fjWHrkL3fVXC5vqrI9dDz0/dbcts23kRDfSVe2wGKlKEGX
JYUnl6pjyJc7RDd/3h50R3VgS7gQe9mdMC0FvPDbVNDPdMvxNn766cB6WKkaJr6G
K1xl+QkZFYU4HougaGfCMjTew435pz5ugu76r77EbiKY597ck+F3ctu7AnKiyG1T
pQRJwXxZ39iToUJSqvmfffRN0AofFfwWuxB0XuEHYY40LpHU/1J7w4D9hFt7sQTI
s6JdMWKWTDuAabW2Cu3zt6ecS7N11IbD8ZjL96xtM4M=
`protect END_PROTECTED
