`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JyMerH5DoPxc6/FjpUSmIccx/yOHp5gYmTdFbl2WULMRmIAsRFdRHbNJzaw4WDh8
3/uE8FZwiL5F5YfMDpaIEO9fbPeogEgCKUdZzX/Nh+WWb05uHvBUX+MU/oLYp6Oq
iEkp5FwuGniDorC5eaFPx7hdV0o6KuwCtUcoKW0hV8owTrnU1eXVyRL0cxZqnKwc
a6QziI2q609XPRmO1f/0o4QEAlabDbN75ueBjt57LDuGmdw6tfhxPowGpDvMC/Mg
J3mYSdf/nsJgKjZB/RKMDJHBz9P9EpjBJxdp0ggxRw0YCH7wc1EVYXdy6R0t3b8W
yBpmJ717+VZUXtMBUqCrVoglvz2giHjSEhD0BwnnE8vZP0i90pSs590/V7bh8s+V
48eRedcrDSohh2jcRziV8FuG1nlWw02RCu3UaHxi8v1TnJSBr4Rol/USelTCsXxR
`protect END_PROTECTED
