`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XAIClHF0uLqLZARFPdbXq+/jcYnKWPXZjabQATiPMNNoaaItnEQyJvRtiyu/JnoX
OwoQnmv8vUW+HV+svEKnAmC7rp6sl8UUhrEzDPGx3v6su4JoMHOuzgtK9b17aiXA
3afO6giik7CTxdgg/UFt1sG5XHFSvsqWrNhJojA01/huPVOGUy0GdX4M29q/QC4F
sM2/Bssci0zHLBGNfGt3I+1cHU6ILf5gXywm2VhPTQnHwedZH+59GQxVNgjbfxls
Z/RYyYepa+SvpPRnPpJWPTa4JWq7kMjWZV/cJdTgAPrcjuTU+n4GGP/vo4/PgkwL
2ASK4UuCAbMQzvDycN1Xqh3ADYAR9fWP2p4lyqLK3h79PyWKbm4DWKoX7fQrbTP4
3thhME5fXaa6pug0Rw2QGBKJCo+xzvOPSMEk0YBzDwgMmnyoBuwZjc/szkpVNAwO
8otuG1a/7DxDsqewb6/VujvGO1TJAJ30onjqbck3a24KNRSTHrtbt0Y00Db+lTaj
49pWmIIYythKpyhJrpfEtmSEJyshSxFkoSyWs0etI6BBzz8sHVtOEtuELwTkqMGn
+ZmOE1l+EtrVnNtDvVfcAwLGPHkkFM5PvFJgbTH0Ujs=
`protect END_PROTECTED
