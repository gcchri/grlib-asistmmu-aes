`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
USeP02mFQRVchS5JNG4qEbNlluuH4L5jB4hPZ+wPl2LUUjUhcE6/0db74ZTyy5l/
pqN1rmkzeCU08s6TZUifrqW30Z6Sye3yJuUndCHBMF6LsCFKYjW9dp5cfsvTB48r
mOpfTJKHG+5Q6pRSHvTdUjJww/WKN6AGj1e60VFEVtKiTqM0Uv3RJbRajQbf5SaY
185uIMQ1ZS+EaskbHbQ2NaX62tnj7ueFiAZ8DUi4pcdgWac/Zv+++3JEn6W2sbqS
9N36QEdEmWd2cYVTVip28uQTV+NH2i8ju4Mg0++mlele+tRCj2NDUW4Af70Whuw/
kF7uaF1IXLsN8qmf9n0FSlMZ8EwfgCxCbv9Z7bVkYbDe7Q+Arhez3bp1vFpwna+r
`protect END_PROTECTED
