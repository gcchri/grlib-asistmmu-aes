`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OeoGvQ7Mux+Emtzr90zCMIaQHBbRISBmSqznb7d48kwJjFIcGglTFhwHIWlKZJ0A
HHxcT9BJ4V/QUcLelkC2m840xfTQV6wCtxUggmq/GbEK11iioquMeFhJw8K+lvIB
ke9cYiyhq/b37dhJIGtt/pcurEPcb5lw5+b+6eawmvvqc+8hIOBmKV87mdmIdQow
T5jyq+1Us97kXeoIzY7Nq8eSgKxXnxlC+nr6ctCwb82clWbxuAK+7DDDFZJNEmK8
RTsxZozmNXwW7N/oV/a7zxbE/GalarZEJEFskiVoZEaMF88xu4R5usS9ek5c7OJb
`protect END_PROTECTED
