`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qs2ueMvB0W/y842LJyYi0l/UCqdxOmvUvYEC7Nsthjoq0u+wywqxtwTrXzjhg4IK
iyiKGv9/vgC32XEI/MSRbMsaIVc/p4hAvWAemz1WcsK7blkr1alav3vWZNG4kHqI
VN59a54AH2bUYlq3/orSYhsxXS/oMEea4wAhUDmPa94JmXnZIUgrp/Cqolk7jv4k
Zyb1CqZUbT1Fv2YoovwLStvKXpgIKdqcGFFCRyZwDmXH2n/P7RdQwm2VP4gfHO3i
`protect END_PROTECTED
