`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mwCL8gfx0PTHmGV9dh8y0AVcCebJEaIYIrfDNj48+ZJTsaf7YWmWDUpOxFexwnpU
D9baALbft/WfjZZIaLC5sZe/ughiGVRqRbBUdeyeMtuq+XSEductYwbFY0J3+fdB
97XoTFjCj3ipT36bljLh/iSl0ONE/zhp5gzd3VI0XgMMNvF6N45xVFIV7WytAul9
/F9AMRd+dlfu6+TQ8tG4Uv1lKwBQeBgGQs0XqTu6uA2nv8tezROAWLbMs/GcCt+x
bV0Y6r3XfRy4OHkNAxdXMvIGlJvzQQJp1a+tCdVHioEko+QZwkDwPtixgGyIn32p
jyMVxdozVfMzC+LCBAAQeH67KEh4shuwMwg7XO2FZha8JHihaDCgpVvHphCGEe7W
uI+VqTerGOuGmQXU5yydEbyFdUM5OMcPaQkn42Mi47RRuUucqfOubih/h5uCK+BD
3FAT3qn4QeE5iqexVxoZtcCdVDkwNCOMFKmqB6cix1sXWVl6HLAC4OOxI9tvU4bP
oOp6BiwMNo2XkLnbyVaKEKH/8hccNxr2K0x1fxdTPaeo1Kn0x+dO0AvSLlP1uhQk
9Fp3pmWJBf6491hlatiXDEFS/BBy8GYxCP2e4ToXooduXN63ffYxhfRnuuhd8pkn
44sVykcbOOzZAyvV+D6+Z7usUCxtSvfb8uhhRsEDJQ2XlWv9ufZ52ErmeUJU+wTd
22fEYwYrIMJEoTo+oWHcnB5W8vbgjhrtjvrKOeNPP4RkpvY743CRbkGWI8pwKSgb
RZtEIL7U7lnDKxPtCUfh4P6Z4s9dHVGF8Aavdl1vgIn8vyQBDistibBRl8yflGZY
C14wWNaMeAoddkyoino/V4jkm1bBwxw1S+GNrdqFxoqcUyNffbWPN5KExvETdqkm
/xCwRn9maL+3OECBGG1EyWOyy83M38Ar/bIrRZUxNXOes0rkStTUeA2FX10oIcKz
Vr2LfMxOoFm1mBcoypbzNVvDKTTZta2SvwQ+I5nLayuxKfgadSt+dMbVjevbQaoR
QIxvR9j6vRXBjC8b8bF+OR2nIp2omGmqMbOG4l/6rMExKRDF6GNcv/lFkz3pJLB1
VGiB7yMcMX2Wv91Z9hpll8LFHgoE3Im8B9eqWtvof8LFKM4C5yp2OaMKnjlUuskq
L6rhRjQctZiHixfPMexu8grDSIp4k5ZboDirYMGjTDajVeDzIbE1ODuorFCtRBu7
vPBUnVA3+UHhO4/oCBhcH2i2ElDHUC5DVePuXXuYBkpIe4xbrVfxbxFjm7w0ibcL
VkJqURIbGuyOQ5nv6sGmAc5TXwkBOr603mRfLLELVyOO3bHvFji6jp4e9issYhDg
bgweOIOshLjpU5QpLVxf8u/WW8jvPBdbKO7YsRrAWcZVEAJRogzzJBGqztqzNCBK
I/i3S4DOkD51pR8IVAriXtjWU4dFNHnEXDfJc9Ih8dx6tsl9Mgf2eaynPnIe7S5i
YkVNzN37eb0OspIiUdps5vGXxAQ4iU3S9rHOFVE5ZREIDQYF9baV5EJPb6as0Y4I
BWeEfu2OXgSVDSMb8H1MQbv2q9TKZ6MRz7FpDGGwLeXJ96mBYGe5TYqRWw7OnUOV
JRJc9w2xFDJzrENHmbHegtp5OJa8QsuzVkymXD68Ib+iZTKqkBh7SVAZVfN3FbyJ
JkbnmLKLsu4qtxssQ4hNv4/SOKFAdF5a3eSZFGhnqItn6vYaEKBpU3QNqydBprZg
FUWvBCgcZHwzWPenIWS2LqnNOoqlVC/Otflej2h6RTBLL0KF8XrOd8S/Jq99tQyR
LiEflxSPKRsbJyAM8WX+lEpzae3mCyEycPNQIqBMQphOo+dEvsskto2NtLTsRl87
LCIWNztEyvYPjYPv14cGJdy5k7Z2fobQM2Um0zWhhKABxPmPs1VWVh0OewsWKWAO
AlXp0WhHwV1v34B85P0mhSUNCsGhzaR/K7/c6RAo/Cl8OGHLBoxZ2fQoK3WiUPN2
o+JA151IJwixECmSFsH7xtYVSamsssuQiGESHjfd+JJKPUX5kcaI3co8JkO0gqwy
igc1YsRMrD03wlZGhY4sLUSzs+hexHaAGNPCo72oDmjVrJJ3MtG7mn0C1RNv7jjG
i2PwpUhlPoB8CoCVl5DBb3rxULJS8TBVX1A3AAbiZLPbqjYdlAxmQjxyOHcw8qdJ
OhRxtuFsNpufIGNucoFvjI93CFUlw/vFeSzDdqD/Saj/nxpqGcIC7ly8/65lAkpx
Ukh6CQGvpm5K+lkn6am+m880dT3PRKJn4qopmBUIksPdzZCI2g1t3wum1Hjne/xX
xOOFGUeM9tl/zYj1YE622q3l2QdoFVSm5h3E3ssKYaiJTKXvsySuDNerV0ziwlwy
5IemovoLZFTS5U8q3QscV7GM7Wl+2HsM2i/z0Qbr7WdYaYZtPGyQCdEsRFEEKkm4
vf7WzlyFq7v5hk2hvqv+K72SNXuTTQO1rXwrtBuacM2/az8LNja7vUJ4HwQt3pUO
33KtW1E7L5TBo1BdryxSQNJVjZuqBJIFop/BBrVs0fBpgynrYgOONgnejSZFwXiM
uGPeX765tY/8EdYGt9nBJxCMHUROWZalSmpfNftUn+S70+mUxK9GwDkEmh61j0a9
pNQw8fJf5JHvqvIAjJ3L2g0KH9pvpf22N3bGMmpU5bA=
`protect END_PROTECTED
