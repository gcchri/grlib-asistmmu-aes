`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3LbZlQtAtotQ02UTM05FZEHZ56EkvxInNeJAcEZVoLLBBiElGS3i0nuym0I+L5K1
Rgk30upiTwVgzJExp+TYRKhlsVUoltOU6ZmmCZWULy5qyplDt3l9nFcnBffM8Hmq
nPIDbkZbNpEq6Ff8xkPYXLJ5SRodaPQ2nPKfjzbVDnPBDZVqJr7ZJQwJHR+Y0kym
0+xrHL+y6wJizdr0oltpiGsJfcS1kT2mRkTSzM4lLOIUGTq2RB08fHtdcb2Z4Kns
29JuFpNSBJAn638o5/H/JhCivW6HEur4wGWwYH88AJKcf3owBVoMcwsX8cS4T3RK
yliNB42cS5Iyax3Ghf2pHw==
`protect END_PROTECTED
