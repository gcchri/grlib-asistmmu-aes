`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PQUQfiKlgiP9DA0gRUR4eSXRI0We42FBPN6j5GtqfO9qrjfnWjNSBHxofjSKr8QG
24J/4c3U7Z4CUE4l2h2rueNt4xWfIXn5BWZ/ALFzzSJYA0zNLfEsDl67Bf1ZNiMY
UqHx1XBGlmuXA1p5bhf7rNljMFW2efgwmI5OucYIWg5i5MJQ7vctEzTP6T1jm/A+
TKk/WAlbfWI7m9q07kiv/5NHH3m5LYd0n+vt5vPZ6e6PnJM9R3W1qJJFKGnUr5yV
2OOCkIYmFhEMmsm061XAgFMzGgQoWUUz22+kGyGXJKg6wUfeGMgb+zNQIRB9JWRd
HGafq0Qnlk1wsdbGKQo7RqA7ki+fx7VwvX6we/FtZipkZToFfLAfSb1oMB+Y3yQY
CAsROuasamlmqHE42U/gV0MpSHEJrqgQuDUI6v8JmKQqEYoMm6XtBDaFVx7k4HOw
tV9UGvEM4PWQQXmqESLiwQtrmfaUFnQPxbInlYb78BVzcMwkB3Fs0b7k0aRzvBY8
MDyUhkjgJ8HEYNJOdw9E/ZTGCJqQzrOkr3MzGacBf9Ib/25PxwHamy6zsExyWrXY
3ydnUD2vrLeYU9JHVTx62dRYCfY2Gr9YbE4TEFdMEoQ9Suc4M+EOIufhg9wUcjUw
hQJwkPYRDlP8m9rSZ3O+wdOwrGDftI7bOIkJlr2PVjRcFDGnCSrsBdcsadCDg5nF
HN9jt4Y1ozc4+kO6019QHrGXWaaWAySvuHjRzG5/m1hjkucgMnlen3HW7WUOmy4T
nRDM+sDivb0cYg9kLgWloobn4ul1dlml8TlO75BMNqkvG5M3ZE9hg8UhY5ERaHZv
b8aKHTaeQnoGy8RTo2/MGF0aA/oTzE3nkctpFnBfSqCd5GfNAhGUIM1GihkuMget
ivGa7yus31CV89uriMkw1ml2RnZlhJ1YilVqaISEFIecgdiZUyYR86tzuuJTs6kp
`protect END_PROTECTED
