`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mkXAV9UHptyS9bCHy4Ap4PQVsPwBm/QPaZxG1+jfkwxLdBTvzCokQ889Bg5dl013
JsQhRmcQTzJW6kE5gSNs+TyqG6pWSeGzxNCyaY5J08Y+2sCoFBF4dqnXLwjvscMD
0malEtlgq78iILjyVtZ8bFumZNMaPrei8aWIWCUR9yvwN27K8k/Brx0aqg0YIs6l
P3WzsdOKZDcI9ADS5lFJKAtyCQcCbYK2oZ7ONJ4aOy005TLQZFi1Wn8FiOuYKQ+a
rv8CX7ajD3ZM4M2VrJ8993YCjZoA2ZgyDLCEHkPu7BQmFWbj8x05IPlCVbrXvH+2
1cHohslP60iGIgzGPv7C+mwxfYi45BHHZ5FH55HBfgYnjuWcko8OAee4ArRCqgkA
WoqkaaGF36p7dADSDi6XOIV3LY5Wr99DWrEVRDrG02g3dsJJ7VZG1meVCEqYS1tk
Np5vTW3mjARFMFCHtIBmIxUAP4DFvA/u9gzqlzqRoOENxsufUMxBTqcOgculA4zM
y8VzAXnyQlxnJvW0zOx/WbOWm6BrYP48yMciJDokskFRFIl6Z5LL60g8X3NGdTmQ
d74b56VSwb0aSj6PWxRNzMGtUl8Xv8DnhX9RP2lLH68JQdrtDz8agUhb6cU5HNj7
WAteI5Z1eBTLZrMMLrMJMdBkIBAuPvK2MWhZi9q4g/K0vVNb97GSHsy8+igDY8tv
hjZ2g48SBEy6shs/SoRCNbcQOtj459J/Yss7xax6PytJ+vDXM3ZD10+jHj8uDHyF
8UzyYJ7G5TZKQoUaIjnq77RmJJcDw6UhlZwtJdRrOuNwVv4ZKlmivI6lE1NsKlXf
gUBiMSxFEselvthskFrwCv1DT9FzoEu+6EcUOUoWO8nEVxn7rktk70+gqNi1YLu3
8DvpQSfxXsjdKhZWK7WmKKiJ6TCAu7C7BtbSXVoHRIHLLngwSxUpoZ6GuJMIOC4g
H5VBpZQoMFu5NN4jdMWf07UjLMNwNtMAlp/5J0g7+ODt6scHl6vIkpFEyCx6VmL1
BTrhkv5NPp/M5pmAiglzPc9qxwA+ZdoxyhlL8saL5ikzQ1spPC7sgIKMxUGn87So
6zU8Ck0LB/ADCOQTqetcINAEJvZJ6FuDMXTvDmKezSXrtp2UGwRHn7pGOEMabMBX
N3ImKfyTOAG++eTiAyfqBPHqW+YPr2L6+LLUVQtEltPpFyMj2FPbhyJ3pDw1qp2y
6fLk1ayGDepSME0HdxxKjKkpBkuwgJKr0Lw2pX9ByFv/4S50HWoj6l75WNDAMOtD
sFCridtqd0UcMePxix6pvxuU9t4C03bi+E4HPVU9LPeIT2psn3pkqB+RUJb6D+vJ
`protect END_PROTECTED
