`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ecu1XhUgT7mw+8iarIif474i30ver/X4irj17yXaUahmwQtpH4ximaHx4LEhdyUb
7noBNEXrk1gzEAJ4gRY8GpcTXoH/2yOps7pVAjK6U5JoKShXh0sKsz5iZtyDIdpS
gg3Vj6zLe/Q7UXvKNruRuAvHBSWU4lXMQdvDXKvx7gRK4RUxtYcd5CE4KTT2sZH+
pfqXIG9Xq6Tr8wlwtyM+mXUYhOZffFNL0H5+lFvT8CqSFQUyH7YdrpuIBnn7TK1z
th3ku45BmV89rkvhMrkIJ7gF6J/WHAychSvLvsM0G+vmTl9qG3izY0w9tj+de3Sx
BlhTRzz/+lSCcV+8BesPZz3BFePfY1qqvo+CyS9fUWWkpRh5JZL+H7G8geDHy64N
4yEJUW1vkS+TfWNzcUATc5/JVmX9exWx0e/ArArA0x+4W+zJbsH1FnB1GEWu7Wzk
dPYh7kma8rJ/EF8aiHVeSMyNeHaI9YF6+6bs2yxk2T8IB3pf8ZPRw5OUDA7Mn0VI
1nzuvapQy4Hz1j9Mey1krpUdJ+IhuQ0HFX9S32zAA47q1yFiFxH0nXWIF6tPbPkl
TboHwOFJPk6cLkVgVp+kgeLF7uaDgxeukaZQpQvDA/bEi5x3rbTPgtKHnBMex3yF
xecvtvrY7bDM/DUCNpDdQiEf1yFR/26/pj6l8NpHWaGWmVY/+2oqCuhhHPxkpTfL
QCWhJE6ylIWuPMhQDno6/VMR6/2xEJbuxQBUe9OVB/gvfKvPA9nH+feABEaAF6ip
EKkf6ThSAV40dN2dB9nIcQtOqxM4xblceUg54v2NtrMkjgyaG2WDimJ89uztXa2q
FGps65A15p/uVQWg/3go3DzQTgvzwsWuk/u13ocn+5ZiYfgYfUkFaQK1Xg8zoD33
5tOdHUoxFklENJpdqlZlnkpSSo7/HVzjyDUSnYqsGjAlv41QipRq53yKVPn+cmzz
2RpiZJ1a6FOiOaiZ5we/+DCt7cdKxVJtaiyM33NTZa0aKdNcrKPHb4/dG5FEv4QH
fy3fCqXG11A6Vv7GjlxVBRP+Tz+SzBxUMGUtjLt1aqSBa08QnPBYcAfE+lQ/ta0d
LWO5cgocHCuDiKIBx/pILocHzm+cViDv03Sa+qMwggULwj+E+zE51Xo49Ft+4oy5
L5U67eVFzzuqYJS2Jyw2V3DP36dkMzJfH3phmLIqVVckdj+wIg8MCKhksOL/8t1w
OjFy8EqGOnv96uV467P+gIlOJhzgxMIf3ML0+g/BqHpezNyKvlDBJhsz/Le+rYyd
AXCpAOB9Lg2KpzbHx5dJd8rXnqv+DPa2i/iFs4EaaKtkY79CTkfnSQwd/9R7RepT
+KIBUWioGE3AYJ1DzLOiaLUYdPduLGAJj5ZAYTlQzrL1V0/is5XewCwET8fEjURU
fDRKPyxbTZgdg5SnRROPON3udxCj8++Wmt6nfjauA/uDCgZBhDpMUuiheWPciMGE
5xv+QC2Mw7y668ko4uXE+wGEOrspvASdMppeJzsT+dTraUP7/Of2v0oFiA4a4/ac
O9ZN40jnZxUmxUXu6By9nL4kVvrpnSyVQR8AC6vNma0zym+zpYZvGNcxamU+VVvq
ohds+VqodWFToqfTHvaabuNnPPszgY4prJ/A0LEVc8oGL5zg32wq0iUGrLYIc5eg
zy4hiepslXQ8GDjnHJSz2ZZeRkxRjz6EeIT0m8oUi7+PeG189wRjAPN+q1gPsCga
1j0F+ZM4u4oV6+L92WORVXGAZzwjFntOEc6SGFLoqFUwDDEHSXYQusdyE/dbVIDO
MBgdFqRn4Cv+m1HFBtipr08Mhgm6fVKKSTTOcw6A8+ssGKVUiQDnxqjhs/bYDFiY
SZVQDAQdnwvoirUvSlU3mLezmiSr6WIKJOWqmBfZqyeGYEXc6BOehsqzUxpET7/I
BoE/Wek/OqIPbTro4BPR/Eetqkp1PPyo+Yd5rEBS9VcBt/B79pm34RRzxmwD43vq
gqjZ9vvcOhXJIaH4pwuTBoidqjib24DYNLIRgIu4eTqz4nqzh3I2vTSU3nrN2g59
GQhsiIfL4VHgzJWSNb3r6B+REOwSubQAN86IszRl92baFVgXw/aq2LQyBOJCZT9R
sQgOyKiGNW/48rDCZ3vQkndwpC2h5AOxFiSCTHdNMerPv/r+5vam+Z4znNYoyIPf
Zl6iKdN/xJqNvev2ZPxYAVgI7RxfobrOe+8NLOaSW/pXKsspC14p6TL/UHdQtdmI
T0f25+0Ppxhmv2w3vhkhF5eRTuVysOvnatfeod0A8FN4Q0iZu94t72ozPLpXPXjD
D0hnsKx8mBJr0UiCFsnDclvNwaP9J/mBE1ge1q+fPGp8YDioHd6aqbQjQJSmavmE
5yJLY7bw0pZlBB/gR8ZRgJgMOUkBKo1ye2YZpP7UgG2+UkiM4dhtjMuqJeXkkyUN
vVYiahumE8AUnl4uDOq2Z3wvuRMqkUz0TtWcG22odjOx+EXJIFAM5CFtyN1Vst7u
MnNl9kvGfeUaI9ciQuzqXnrRHztxZZLGGB7YZhNBthKHkgPlS3RuoXu00mKGmuC6
sgK0Oqjl36tWUOf72IZ0fb3z8lr5KuOAhzAS2mAAUBNjt+jp/yzVHXose0FMZCcW
z94wsZwZObCYHTSiX1a7gHN7sw2upwNuM53+oPd4UJgRp5nJdjbK/d1l4dDc/xlH
8GMaJEoFu1FNFzB77l8evdon5V4dlVstRhbqdctuWFhh2CBSIr600QlbIKPS5yBZ
5PNCUU2/KVEbo3lTEK68ViVBGRCcChg3Tiu9GSGKbsP+LiwNAaiL6xkBSr7x87c8
bZCCAyjOfTHCBxWN/9OMMZaGnTM/P9O+rVtxvaTrwfbmWZJw31prGnhJUn8lUCXc
9Q3ZjIrcp0PJM9MKl7k2Nsqn1Qsac5XnhPi0x6rwOqT1fZJvTzly9/V7RssD8DaM
9gv1eSWIWuLVhWxYopudUOtLA0PeSVMQ4gJ6rd9n9suTcpGieY5Xru7hcae5qFhn
FlEvHNOrIwmiiV/q2SMN2zD0lkKYzKP18Xn4eBkTt7BWv1p8aF0fC2zxArlgFNL1
b0JB7OIEGjjByne65n7Z6OkMv0eROC9EP5NZ/Q9kcHiiHR6anI3ExK4pmtT0cbzz
vOBeyZAxHLcrIe7mvLavr/8Y8e4sJpLuvh749V5dFffWFfkWRMLyD5KzQmzl+goJ
uf7/Pxv/3lDFPFeBjUyCRmflTRRWiCvQk3c8+d6tgSQxEwD6kfLmr4J4kCmt01JT
XtY1y38dEkK9RoEUobk/nxg6PXeYI3R99EQVRFiJc11hWYt+zTRfHvsltjXIPTC7
Nkah3/9VdWbxd2QMXWJvi7uJTepIexdNxKcsGkUiqN8HmoH//VIkQoFotItqK9cv
jyOnOTSIWG/R4UchT3xmCLnotnAJmM4+xyiGXbjIby6rT5iHvH/Pc5ybMB8fNKJV
R5CXMSyXDOrZ7PvS7XMSabLRNpo7C9aFzshQX8aEpogKBDXeH08SCpjQJ5vg7FUl
hDnQzApjoG7tITKF+l/n/02g1zM6nA9BZIgQqK8VR6FLzKZ+MYhsSE1KYiPdBrhr
aLX+9C45Hpv3lAukJLYfsYd+83o+YkWtbfedO52XzWc3v+4x56avInksUKHXXpFt
0S+mnJnERyDbKyiqXZ5AyQhUB0r0B3t5q7X0Pjr/thJPKIfu/xk/phKgqzlNsquP
OaHZ2BlIM8nd2xf38/nCuiI5CqiHdMna9dW0rjXnA94lqMvaD9lRRCrRiQdCIo5b
+DGZjfhTTfUULNZCsQtqFxhfwPGTUHrf01cmM7B8Pcqss9C6boFiW+IiXFAA7XfL
kUMydr7bAALTX2/rrXPuuiEncL4YrkJiu1rOrODgHPlJMN0oQv4osLG/3Cd0Spik
L4rO4JnuKprBX/OPqlua4fvAPVfEu60kTwq9FmJflD3VeLLiKhNCXM9yrGnX+UkG
0U4dZ644bLLOtbusf4J6qLW7Vk1W8Mij4YvyXXHJKDadGKjxCcUgCXQQtx0kg716
lGY+CIwFutHLst+YGoJKQZOPATeXvhxlZzPH2hqO0XAq0ximjMHOuvN6EUEbSyVn
SiIrQkaDEX1K8NtbusXMVsBtm46nRhHykJrDqcaG3tC3pCG1zkIXTCiGHoWx0UDN
fAm+WJSYAftfG8zahh9qWxTILOUAD7aPn4g1mjPTEHjJ7lQtZllvaSmUAiLVOXjR
Bq6EC8ucJdaBNgC/EvoDfND8SkehdFsrPJHePh9AaGMjOGpFNlBcDOkhMRaiJ4Nk
jfMaOKYe6gWZXjXWLpHKQTpAycf15AEBSbETiYEaT+9MH5Cc+cKn3V9S851G0rin
GYTznLFl8bBf70OG4xXTNViqc4GsN/U0b7nmq6UeYhs12yzckWsbrt4VxASkyCXD
AcxKrGXn6oW4Xc81NMvJXnE0IY0XeUpfWsw7AG1eOv0thtiwAX7Uk4vVOv2k7BfZ
AKpSLOyN9zrdouQ0a0DAtgQFQGReBAc4TLHQyOKxETxY10OXu1uNWPauLze7QPbl
1TmQIa9q5II2ji3VuhF97XX35vlO0EQPxjmdYEJvQkomoujRcMwZ6QprLbvCgdtP
a7kKGKMSG+AmWVpaZaTd1ill9zuk+jmr6RaaBxNfQts7vn4dtrNLGszq+1hDPyij
mr0vFWAxOfgAeUlY3ITKSRzrAlU/oRnjrNhmvZkglAl2Hwl8dR3kf98CVNP2EHLY
U2yhAQNLy9voMjLhxa+fqVaJbxYfHmMOBzmnFAFUNNepBC8TAWgbjFuBaTbnv/x9
Dgl9jrnaVwbpDOxzw2X/yZh/cvr1A2P5dGRBTpoJAyZfrtQmhBa/OyhIfwIYrIhs
5xct0mHTy0N1zKtVz0yHqka6vKCrGMsJOcH2r9afRLpfkNE63UElPesjbf9l8b9E
Z+8GGMCXZy0ycBRzulr2mSAIWye0iO6fcg7g/yYiMOV9DpCSZUUX02xXZ/BxLZ8X
TLjqvsxNj7ZQRcqNjhKdVoWj/YKWTmMvP9zup+Iw+qZlos/W202YRPLJJxqja1rf
UA2hNIjZl2g28LWeY15ssDukZGe9G29M90PMJe0+jqfnn98yHDS/bShjGcIljJe4
mswd1NgxBE8IpOyex52O4rlRdBWt0r2yYGZ0b4Ie2TpZn7g20u5ZJy/OWG1/xP3E
Rfn4TG2ZsX2c7q33GszE9xZhX8JOurEF2ktHVyELe8tjwS+MyKl2ymx+uxtdFUAh
vtf4HrNZ++Rc2OTVZaSMtr6+EEuz4swS/AxxbaWwvDLvMyWg3Gy1JECD2iCGCfW/
EDgHJisP3sHytrJ9C0Zj43zrjm2wFDEtlIah5Yiiw81nJ4kHSmTY+c+tPbQGF4Tn
luAjYMa21PuaEyRb86gwjDK/0r84pMKN+9qcRRV1zCAdmGzSOcs4ap0l5djxEJCt
IvHaCP/s6k1Dbigy9J/OIzP+PG3j/8gIhRFaG/RJBMnDbUWP7Jj8oqiO20iop9tr
3uj6Ufm6YUs5mXm9k1sRylXTmNr0+G0jo9ju+zunllE+EEVaPfo2gyTBiPsUxq4V
eweHs+fjsimyUms2kReTbPm5z3xu7Et895kwRpc3R5wtdFGl6NvZ0MQhkI0P38c2
B6i5Xlk213axM66gMog3cF/N9nxmJ3YpeEBWSjzJeTs1h/OdIskACanX6TiwYJW9
LTyEqrtf0UgfH9d6gyq/LRe0Bt2A3eHJ8KA4aA4nq6uhaojb0CAG/J9Qma/iX6sO
QuyjfpnqPD4Dj4p5ZHlt1D5nanz0cLPZvs2FuMrqE9O14TIdatPA8kis871ic1aV
GHj5uFpVZWvVPL/dy6e79swXmF9vUcQn6FkVSNGbnI/TYkPfKimc1QnPIN7syt4Z
HuhbDV1XbHLBGX9EIp6OJ3yy0WUPSxAdOBPKLnBMrlmK0ynQS+cz5ji7DsA7BEXV
8S3w9sS75ulibzUDcR4WLorxIbNbJPKiQ4ZqLIMp5edaC20nX3dR8ZgtJatKhZH5
8bTd2YPzSU2ZMA6L8od+oEG503sJipBDJeMC+0kK51PjXj/NhIKy20fiXg2dgfuO
vWokBZ61dPSChxLxSkJixztSY9QdcyhuYFEnBbJyfmAfURZubmCUJrUu0hQj/e4G
7MFdZMLod+dk+XJxFIrZRFtszzQxl1PAFyCm8SzEisE4UG3xDJX3wVp0sBqu3lTj
1bYybi8qw1Agk4gcfg3PHyjBir9vumoccMgOzP7qo9yCnRf4VWsuVCll9iRmWTGT
J/PAtX8IbXUU+/Z4WZEjxk33BT8EXz92G32uJhDukIsKYL6pax69SCgGvBDGLIBB
rSsPMb/68pc3eatPrajF2J0LJRnGCubRz5JjUXPzRw/YB3XYpNmdyoE82jwXYeYQ
R/YZuO+hqopj+zlveRHqY7+gTuq7+4RfsbR9LWjOKjtzZfJ9avOwjsN2As6/OGCR
drJyQEupcfEaY+MqS2Zyh4j2axZZfcarr9jV6OMALndoYnz++UCdwf2vogP+D0Eo
DTRGlZyEdhjB4vYJ/wJM1bjD3WTpuGkotucaNpwihn4ndnhmVehOXs6/zyEIplkM
06LuH+s4Enz6PxB/EfXjaRCXKcBlawHlomjfr3AOUyyz4I8noXY7FrCrGK8gHFEj
R4P0gdArisZ/LxM7aPg8sx2BC8TA6ysgIvsbUTDN+lle2VLFWcGLRkUltLxiBjJs
LLZlVj1fRY5OZlvsDqHFjMZttqJtheStyeVqCZ7N14H+QMccecg7Wo9FtlVeo9VH
B9pA2Encl7Mv7lwZesV7tiNZfByvQp2Uz3TQzF3T8/DTz8qC+zmoD445O/vgdhRJ
2QtOH/GJAvmODpFzuqhYCnO4oZYL8xvw7xb7jPfG376vhMxD9V5FoaqmpYcuo/3Z
cttvv8QVB4LyE4utX1TX0eavtczCePfBwKgfajx6Xbv5QC4oCB/ldZVm19Gdns0s
FMb4JIkhlz5SjMZqik+dOYL2dpMdfPiJIvKrqIBqotz88MbqUNO+3BajxIIz3MJw
wsHeRk1oKiWUcCgmBaaqX0waeW66AHg9LgkeAmNTID1j0UjDWzqrqTbnNEZpX3jz
+9rcQW4pl+s+Gvmn9glat1KKT/BSHhGuby6BFDYHuK4MwQ9wWxsrYprWQ/cgUijc
PLoWwBcr6VdnCn0jSFDxvNqkSz3GfTFVsQwOjHtZ/GCCJ24tM8j2Cc5L3sQyW5CA
I9s/OZ9RdZAcAYoWnsmA9kyZGtZNcgzdO2+Z/uoD0lfoJzipEEgFdJgT72yU3bie
LOXWTZgeKWJqbk3xc1BlWlbV49HW1tQmDeOXB6wD6eIZ3CXF0StPbEzbAmj7eI/c
uDk1Vwdot7Zuy5cB6OYOSy0QVLEW3TVNpCEUtaprf/JxemiGkFas6I1tcPyKj53x
2Kpa7bvufNm6wB7LVHC9Ocvs9+c0Su35SebwUukPoczBrZnwehfb4MZmRAsAlD6+
hdFiNIH0c4Di2M5YKyGCCdxOIJmO1IsYN60O1hRsZbs5SJVOULWfUg+4TusjePY+
TSj095LR+nCVlmrZ/+QSMYJHq+xGkgDMuPShdtRWfWH+8xoLzMszje6/Z99DB1aV
XEzElZ6w4jHOIkQNQZqCuaRCDX2ph7S1rVXihUqhg9TRNYA8rM1gLbl9N2YwI5NY
m6WzTMaysZED/NJWFKM7h8h/YE83ngNBOwWx7RkoqitiRd1gPGM20/TmAZkquqXC
h9IpBcDHM6JQ6l8pVqvDUGp6bG8ioL3iIGWFBF+fpcPXT4AnKWTOumRKw/qFbSfu
4jftTx7bNiLxBDgN8TQ15vfqjgMn820t4eD0TwKbePErHmd499Gu/btTdrAI92fS
XC91wIkrgbzC+0055fzV/ycnEWtY/70gBDrS/17HHvqX+3adQNPWUBLNy8hzodsw
a1zJxd4QFHp0Og8i+rEGGuWpJ7IYx1HiRHoMTLqYh0n1e2vnQSrZcPDQaqYAq/su
KC8M9twpL/HvWxBdQqxyt3pXyJ2IC+HNvqyNneon/tMMCSZlK/7SYIqM1+zT2vbo
HguLRGpefT3j6/41+Lz5s/WJd7x+Xfs20I7NxmLCn5aF262hs7TvRwjMvHO0vEIb
AMzrYa+Mh405mXTeMSEFhO3WoQbZ16TCx3H7MUjqp25FGGqQQit2+lIytwUy2YjR
DHe3V0c38cTqs7r3wxjeelv+n9tT1/FyiREEYTw+8GL7nItd2lG1veqSk7vNiPjg
cgdiZBdSo0IjRA9esWbthNUAMMP1C96SZwdfZnzxDc37BFlULATPXSckrpBnnNKl
rUj0bi9qEDBskWiec27uX5ujqYkL2QGpBEOSv4pv5dkADsprHmh2ALAnZL28o1th
1gguToMJpU/rFQFm0aWXDaoSqGVgCzHBj6J4YlHAANN2mq/BaFqtXGjyTgS0E/gB
Xow5iZaDwUrVOhuF/y5onx6X2wbLKqUL6+6+ySdAG+85te0/vbW1IVv5b6Z6Nm+t
pmKfkFN8vD7Ey4GPsuyrm5YGlMaHXNBIVfTkflOaF8tMaQUTtADQW8BodJpcbMBy
lwYBYOcLetkVHh46EtdcZEEdIuMlEwYZVIUcfy8eGgTOP7iGoYoopd5Ic5wnyuFG
urmkHfE5U2H1YYVd/m8KBYx+++8uyAT5BM1q4WZ/TIycXaqu7BKbTeVPY4712nMW
p8kmz4PG9VtavGjwUEcNjfD8jTq6BkOUloHIsAspc4083hy8Uqcge/JzVo2D7QRj
Gl1jgh6vXp5dLidnpHSEkjFmViMsZ7Sq/cJhDKEhRrlx/cz6MwL6vmC5ShAsV/PD
GrNk4h63FpWPLxQJuWFNdciNDz8YyhfsafXQTNx17IcgSfGIPym8KXnqLqcnoNRQ
wINzDaHEnsBVV14epSWumLX6xEVtv+iK17qUcbBSZ3ZymnUHGNYwrkOauK2Np6QN
GREZW3hq0nM7/SsmjswiKmJV6dTEx3kg0aEC63p4zo0cUWz3hq1WvJiqWcgeBTRU
deHlO3J86GLUMENuyoGRxRc2p+/l/NDZlHbhVpyRb7FKWaFBAe5y7FHiG9nwzdpL
hsl2MAn+R/Kk6NZ8QPHRrkSOg8/tU0ioVJODJAcN5VSQx1MR4h3sLbVshexko2Nw
9bRjvrD/Pv6X56BwKjWefvrTAZRps4YJr5ojzwja2Gcl6dkHB1KH+XdSRYZpf/ir
CL3gXAjVdVgB/3Kbu8Cz3zk7NrAY4xv+keL6CWEhCwSTLD/et38rgPxOo8fuk4Hu
RUL9XsKo0h4TxXMQqgvl5dXa63nxpantmqe4PBkKoLUEA/feAssVotwErLUHrrvB
6u1dkj5FQ2zBKw/u6CJwovr/PdkqusGEVWU24bu3q1OFrwVBZggf9Wx2G2wq5FrD
WahUuLTVR/SlkD+yO+5f3aKYnczIBSWem+0oj+bKZfEJBMcURwEK4COL8OYy7hj4
cfP5uTvMj/J4y5khs8iMiYd162ljW3bJ6rvB6Ph6o4YNSW/Akx7MF+7iWGNm3qLK
AKSBdAEqZbWqwdw9yEr4afxKPd0cRjJfcYjLELPSzjtF3aP4MZJuXymImhfQkBB8
bnq2qmFI/QhUYAJdZUCCvRLSRpHXoxCiCtjeRLga+lMqf7D0d3gBBwF5yeTpRfbE
Yja58ye25T1tEyvDeOeMdIl2kpBM5HbKz0syVOVVO9yxX2gGcjWvpy3V/uRyred9
iyrsvYgMBDC4x+76VJl7YLTM4BpabCz2Y/6qi6WL5wk8pNSEmc7ZqF4kawu7VX4C
hucaXHMkRwVx/8K7SNWD61x3ARaRKYwwNw2LNw9cdrT5uBjJxISQpWGfqd8qqtnC
MLxCi/JUR3zRPYV62W6ZhdlPqVZSnBwGL8f1LgeHkFrlXVZqOBfYV9WvgfnJW+Ku
BVdkfGNF515pxWvmhRhCa7RwP7ySWBo0MLwYXhebIfGfEk2LJsfqpzn0OlEY5OrM
ccPSqj5JNtFsdM6S3sCsob2MySUra7BlndDC9vDDvlV6Yoq3GMlEHIhxgUslEuuA
nF6OwwQEaa9bz4AVac5BvUTcPVNDkRFxYPUtlXs49NMk1O/xC0Dq2eIE7u6YAE8N
gyJSZO1bjamifWq+61gbeNdU8tdAZAfVl67q1BiqRWfUQkypicMuxY7G8l0/BNfR
ugvOTp20R/glTSzKGPgO3MRHIvD82a5MU9i2ItxpC7HIdJpXZQYic2K+l2i5VX3L
vXdaKdzThS31cLKmBW9Rt/yyu8GMK1kaTrzRsCHKZGBsTsHuCHE71FGMpLD5pbGm
N5YrDaekgVn2dCTxCVQhoiXs+VmqQ+r9ttCjDZH0zQ8kbQWRvGjPNtZM8WF3l9V3
NZDXnIpUTm9CiQgnidFrYNMjQGH0Y/VloZCi4GyvIzBuzlWVHr2YzLuMmXRez82A
68B/chUb/BxDnruXKpr8aRwTnyN/5d/J+BXzmM/hojiVpq9ia/6OauQllasviqgq
4ZaEzIJtqhDr/bDpZrbOoiFKZdbNI1vAGtRkO1oDq+r+T/bvKtmNWJ95ZFpfm6Yf
fIQgnmIjgKbrR2thmWKSKbLaguT6iGhsBd7lul9CZOs2fwInkNOiExFiX/3i5NV/
D1vv0rx5QwpNSntt9vvevq5TP+fRbHvXTq1rCv9s1E0yqmaPK7oUlpUd99U/RXne
PXi80xH+u7G0myYs8GUTtNudr577PEot7dCIRnK26qlWTGMCZC6FbF87CZUd3TAW
SeTGQn/NSycCSjDznYR1ubzI/pOl0qzXQVKUo/+lWKfRTLhNJJS9shhQMMNaeETb
QpkwuBrJN5RZLFtTlqDoMKuEiroEpzFKdAise3mPupELmdct/3mYl1Q3B30Zk2ZV
LW8Mm6w1XFERXUKhPa5B7mbT9sSXiDFNOTlR/4uQe60umHgz8hOuyS5weK9vEHbv
utUiTcefIvYe07YycgS01tGTeVCAnzZECkKZFJ2UL2ovgvPb4DaHJ9z4Wl8UZDMH
aK5Uzo+copmhBzqhVHNs1ZFcLu/ZiQH+iHuVvl04tZ5vAAPCFavwLt2aE7XLSAW5
ZsHMI/UskPECwxUnUvBQeDln5vXjt00ZUe/91pEdMvaLzSKZiReD0II3gTiielPg
PbEK/aMbmh2uxjpC5jvwsaJgYr1YQyGu6BI5lxC72lPc/AJ8+WqgQ4my3s/vqjvl
/UVa9zxPmbJ+kRfXDSyP0gpAnYYkk/WHqVm6uUqhgqObeKcERX1qVEMbKBiA8xWP
01OK36LyJLH/sH1QrD+OM2OsPcD9uz1E4WbgTsDjA1u+9vFlS21qJfHDLt4jfKuf
tTxHs5zqnhTQdiGER6pKAe9Ojbl6xtnQOG7GNTVZC8Rz1cgswOpAby7s7gC0bN2E
r9btyF3EDKQHmYspr12EPGieTj8hnNZZP6W0qP33l4wJUzjvpNyhRGnjdKI1cVhS
0WXGJt8hlSjMNVFD4KWrySAEEUp6VvFTPcj9/p4es3HqdG4tNj41c+TMLxTaa9GL
dGyPVE0u7pX65JcQMvIJR1v6ZNMrwEAnOYxM7pEUNZQWlgQ4e6RV0eSjGEp7kyH/
aNVPPcTn1CrQR1/izYy+xZoF0rDw3pNosmC8bjHqivg5hCRY1qC6pqeoRNWhs4sO
Zs8iTL/kTBY4yQMu/Ssvr2sWeVPeABTJv8d6VFN1iV6GsKXWtUbg/pB7qTZJeD6d
IDCjMDYdWemVH7iqCzwgl4VJcfQVp9StHdgSyMDcd877Ef1bhIGvWSjd6jiHFKwH
HG0sVxTaX68knMcdWXvGpNturScF3xwo8rV9fFCN9y0AN9dTOmt/L/hSM2ciOC7K
huPFcenPqZIqMNuoFWkgVWaGnsRh8bvq9ii5y0bTnzNMOUqOL/BOISGAQzIUhth+
dmJ/hjecfNC5lTyyj98ur99pH0ETKcV4vlSAxpEnIn+EW+zpUDTUaI90x2VRDfTT
4Ss13cwml03MkW3nVwIEMrJsKXmUMtOww5zTjm2dlrPjxugNjVO+264hu3Dv3IvW
U4ZPwGy4UhgN7d0ZMsl+Bx4EiQv7N8Iwzf0ePWQ211VKzMoYmdTiPnS+xvLs7qbm
mW7vL6nP5atZkXXQTViA+oZ6KwnYH575VgjmYQwV/RtL7MMx9Mf2jeP2/lOyk1W+
S7MQZY9ZifgJq0k0KvSm7bFiompQlKariZuKU9C00gYeslE/zNV3lNnsqyHfvV1O
XG9Uo/pH1eagOJMSjyuDBfVgsdivwVw5XtwmIJ+HvJAH8TfcpZVY5ceuIS3E0HOP
tHcPAsx2HSi2TcNp8BerERg00yulYBLNfpXNYv2yd7RccW5NeVfk9/KZrt+w35/g
S0qM0Q6Ybksgz+PJarK99xES5ejHzu43ft9uyPLevwFsgvxMlk3gItik+3pB7jBF
0MMvi26+b1VIiyrdjtmwT59ZxkUh0KyB1YSE02Jiqi3uNwxWlQeOoU+L41p7Xo/k
KC0JD0zMMbJ5khd6nvZxQAImXb3x32aNfUow29g1xx1XvfmbHqQkY12D0bU4uhUU
NakZMgin5gLD5EM9uQjBt5g9EkZkKDSjBFluLDHsPYRclnzHyr0KmpxOWAVVvQbK
QWa550WGat/oTwLIMDoOT1vnntVFS/CJCIms8JHWzVKr20DgNN0hJ1OI45TM8oVb
Dq83S+N2x36DyfxBdGd1Bf+LWXp2HkMWfNNSuy1jJKePf1R3tehCZceyjE25g4Nn
RNrTCQXL/CMyRvZJyhN6PnIRxjbcbm413191BE53RgtmQTmrcC7hYN2Fa55S9K+s
itjThmlCedSE+rrYLYraX/AC3Zihf4mvraEgSXqPbARQjr/Bl8jurISEfHTs5wk/
ZI8cvNPL+PTUu4MrPeLNQaYX8a5dY12nEpFA1AwkJAKXn9F+JkQ3ZelAm4bOhePY
CLJJRUpnU3w0X7rLdp77iHW05At0LL328Zv/Uft0LJv8zWQUpBwvdIzHQJjkBEnf
tTGg6XDGhJWl41IBDSHA8zkU+yrFXrUOFN62rJbD+4T9kex2otcTXV7GXJya+Vce
M+r3VLz9EzcX8aLukYKjHFA8XDw2gXQB5B+AIJiaIGhIoTrH/6Vd5Tu1ll0rcsY2
fAWncdC5TdoCOEqhJvnVeiyIF4o6Zibh1cnJ8cLt78XLOJpzWWbrFGO0/duqC+OR
KSLYiMXR/DUe6bf20XjBBGK6ndPXhy3RrFPLxM/zezKcMNEOAn72EsrTNN8wwPvS
TyxMPzK+gST1WGZgPn6qANf+aSpiOUpPIwnI3fo81B+WvRJoUuBFZorpILNbK5at
L5HAb4HTE45+wfP4ClpyNQNzUfrY0/UOrahyE9823QmueNlYZjGFT/7G4IezavSM
ERsqf+hZM1SP6X7OMqdeXtiikO0th26S9aoAIH5azSTf5Hxt0/FAzuq7df0lP1bd
vKJiqDoVAEyD5k0utFwpoaA+RtJ2bnR0V8kqAQ2wPqUy/JRhIcw12RcCbAvWPZfl
jMPdz6dOYXzlt9Emsa2oC40R4KM7n/zuizkwxHuzYNnakqa4V2/MWSp2o89tCY2s
TyHAlvgKto9O9CHM8VDhcT4oiD/JWx37x0CUlDApjsrA4IF9kpw9ALhtekLEXnkJ
nZXBDtKvfurV9nfezMgH4ga0toHPFPyAltSDqRoa/Cj2V0KazkGBBacLiVsw/vvm
aG0gfDf3jIRc3wUmOCH+iqLf7hu6qR0TMpiNldSkEZVuOeWiKAMxeEtEqnGda8xA
4FA76GpCt4gZFZEsBqGIwzfq/6MEViYIqS7fMtRkLJX2VZNNpd8FNZ3iX61jwaFf
vphPqeKcDC4wxr8+ZXJQNUJ4AWzrGfERwuH1szzZ2mn6ttDlpnYJ714RAripqCCn
w/k2ALzAkhmEgW+fbueZErXvN78g9khbVgQmDvGqgSpnOID1tefZ/8ypRKv/M8wd
Z+rjdricv8davxOdwkpS+ns6svPJ5yMAHKK2R4ug906ZA1kg465nuUsybimILpSk
QapkM8ydl/bcJbfi+Su42GlRu9veLcs8uJf0NTJ8baFK4lfAKjJXyCnh6+HXfhDu
xQ5wqQHvnQGwFzhJPDXZC2gldjle/+WwQBtadxNiMJ+5Omr+aWhEFXyzN5lIFE3b
UrHeZ4j+4KaNSOqXS8sfT2qudy1vpwWXKgPA9Rzzenqze9qayCR4ekwCby5UQdku
ABmKGGc54L5HOm6VMjSQk56uGnBpC0iRaIpLevnKfpTEI22qqSEahfUESZjya0FU
NrTlOH8tg3Z44fg215kJBFCBn16SJVS4TBVNkYKN9DSxA1L4IcJhwbY3XfZgoKKy
kWYI0hDYjvSh+xSwUeacwoevMW4jFwoH4+5pZ1d7fZKd8wXK5VwSaKOjqbZAXZPV
zOST7deitf0R6IShrgAnEmqW1V5h6OKcHTG2TU0l5e6X1mdZXKApAvBWzl1X0nPu
EFIVTg0lNhU94IXMuhO0kVvY7u+jMnfSCNq4thUD9nfjLQxLzkG0I2iUPLIsK6Lm
a53WXacoptKcI2ElHZY+ZLixOS1FM+wDLuqdQto8AmZVpVCDFO3y5zj449WRJKfC
j34SgPqDp/DimTD5kBBzLx+KAL0szDFpwIXq+hqmEtrv96XvCF1TclOqJbL20zqE
VbTNZh5Z5RrIs4pj65lBIvjSqWYSr8+o9q/u3SVXmIxRnXWjIsZifXBu0Duj5ygG
aYIPvR+i8NJKvjdDcIzc2oFqMOuAz0AyEY4U8MXzcYwjCoBRjmtsspIcVh52dfOA
+NHxjjtjpvwS8TcATZMJc7ywnhagxPZv7/uFStvK2q6QNABK8b3r7sGePHHp9QC0
xP/0MqiR5v6XYAEVfd6VIdaoD37503Dy/3ZKenO5hb9WUfjSoRH0qkL6ZUK5vhxU
A/BvXYYi4gBLhes7PuS+ghywZkHaT7VALfAac7qAeUtFR2SqjvEqE4VJMHjjqha2
NboyEnqn1JWifa+MzOhCi88Ya8zLFcU/IbDcVSrMHArvkovTeQxJy3wKJPF3AaHd
WdiPb788cu7caYQBDnZVmh0Wrg0kcEfGcORXJX600WNTR9SuGwy/2sFI2UsOc/n+
E6CKeoS6byyWT89QpoDET4D36LIlsQ8ambxm7tLdLoA/RU4iFnRxfur+EKEWaowj
50guCQDiuej7dnXffpS62tXURbmvEI6mklukINdF3+xFsV3G9NW96i68AND9yUij
k7TMmqMASq/qJR73PALoT54uUxDMoVlEZo9cIudYAiOQGA8HryjsSPMfoq3Pmfzk
NR2n/n9j/HtOYwkhFSSdhYdTdoqFloN0wjT+HfYguxDqBi7krYWOnG2XpUuIkQI5
XPMML2oUDmeTh+Lbki95Z3u+0bJuZUxn1yOUUylNQ3L0ZnJHQbCq/DvUm0/M4TcH
4GHMQTJ+pws0xX0nSfZQwB+B1IlfOfSsNapbqWq9+REWSiJ0H6o+vEgmRMTjzKyE
5Gf9lRFs2oLZvMIHZKFG8qODfIp9I4+SLP2/P8VoNw6njR6rqPvxJWseYfns1rVF
qmgCO65G7yyMtNYs9r09saljbybeeHBH3HnZQzkmj+x548p6JSHb84fH2QqGR866
M2x6yS64NpxeoT/hvkCM3k3HT4xXkognuOEEayN6jPBMO9T38T42uUfgWQLlubpP
5Q+ohi9DsSxz5pPgnlZkT19AGczSRLf4D0Utn1FPnGwNq3WbtiXCLvym4TV+5gjA
hAsIK7iJCkrGWDg+OciP9wXLYg4G93jPmJ+mCI+1CW+klj1yTAfTqiXlCS4okf7H
1K4f7d6ZwX4PdC+gYyak5freupLU6IGhfcCmpy/NQFAOyD4BKId43MBjY4/4Q0yF
y6ui191PgODYgpvPIgchiWcLNSuCVGzgcMpIxbgXb1B+1Sy5RZMZPG0Vx0MA7F3k
HlgpTYx9ErSq+wWDctP+hgF5Z+mV5efR/gNOY/OA11IMI8puzEzf8zEkQybvukEx
gLBLuP3FbVhlvRBiP33z4hTFgH+0wDI3BB+H35ksMFu+eue3Qhy0orlXAhKfydLe
zGh++WyiPGTT7LZMMPWPBAvjD8zIDxF5yYQxywq4GwBXeOlFYHdkataGMJ59bsxj
+1Iw5jUK2yzrh0TAQJSg7Sx6w2WB/ToK1+fgk7oec0MRVIkttXQ/TPwm3np9ddqB
dPj7YtrA2ZtdcrMADtT5tZlEGe9s5ZXlsa4xKH3h5uAtQ2zgavPB/JowebqD9HvJ
DDPXJ2pNNQ46s9j25Bq79HbHzdPyopvIFvZouLkQmTIUZ6al1NLLFDI4wE61Kz/j
Ox9GkBkMzv+vUiV38rA00kh0xiyjGzOjat0CjpW06JZKjrk/qbvaXxCmtwSVyuf0
QVYL0thyjJCsj/TfBjhCsVsF01Aq7auTiqazTPmh4dzPMMpW41Dg0fwES/Drc/mg
zkTGn/w9cd/8BGbcXR/yq6gc0JdoQLLe81/fTR42ujiNyA47no8z0Iku5CSeAsHM
mlU9M8owW9Kbc2Rd8KJdccTdw4smgc6cb4wSSfwpUVbSmdlLAP2QuLk1hMwUImng
xvN9GDLLt0IrMRa/ha+3sf1OlJam7TffXKhoskgFWlLntBL+jgi+lg76qwXcqD7J
mWz7NDBN7m5ovV2gpxOh6s9Ht+FF+eo2JywctXhkQAjb3r73X8ITrgjo2YXGYzLp
sS/ZJXy6TCQbqYNzWD6eBfse/Bfx/YhRPYk+95j0QsXmKmi1bV6NjZ5+TfxZd2eC
5oP6mpIZyeJyHHgqISHSYc5FlEkVYexJq4kpir50oOYQ6Pikw2rXPUxGiOYTCH8b
58FmtQrJgJAW4AkIUgrO/AooRgfXDzefl6V3Ym4UU6cfoJaY9R6MSAKatp+YDoMD
pZY/bsyu4Sx/MuUD8eWoy6yObw/fi5ozBHX1qpv7U7L/KRD+ZXi8vFRWCfv3Qwo7
Ww3OCPnDOIzaoZGA5m3TGI1RxPqQwV9e8Z+rRzp3PUGR4c8/WH2KlOLGYt3su8BH
atz3sJnqCqwSGMEjhtzUe/iB+GvOaT15mNl/kgUYgtBfqy0duTnB7P57LVmd3fvG
U5pa5GNBLAi7ZQUsQRET3MAWRo4paI3Z/c/4GzLytg2faBSA1pGBXmQT2GnCD4ul
YxWmbJrBojIAYgGFG8Mc/jwbIePTmt1Jb+cbDDU9OE9u7bcgKSWe5VKtGuoFGx3v
NMgy3oLJlhzee1TvOdLZZfAPwYANn43fw3U7oXbwDP6CQ8kO/+xdbm8tvg1v2cAt
wZ23FmFbpbBQKAurh4B2XjL5VDMDDG7BtA8antskfYSWQd6FiJTP3izq8/zr0lyO
GZmoXxxbHiFjSlUer8HoQHjUGdYK+C2mbI+fH3lx1K4hAwMhI25EZHHqyZUDEPYi
so6jyX46tDm35f+ozgscr1MG3DW7K/MRYbuerV14gMQmWF0+qlZX7T6e4m0Ip2Lt
VrO9D+Pht7BIa2tnRNix0DggoxHTXxGOGEQqbFIkh34kmDDTwcKq4DrKMYubLHf3
9qdEIlrzpO6KMXPpqkpgEKSf39hLBZBZy+Yaka1NAM8LZ6GTHjiSpp79q/OHlnJ9
4Lj5W1zWnYO7M5lCECxo0OlE5WpzOjcCbuNtJFH1mNFi0daq1Cqqx57hIBOxQB3c
6QOTsr2kFC8QUz1B4OUImorpAZHTC67p3a7AJiBkEMWUao21hwugVUu5+eL6/YWC
y5hviNHyISXRdEWt/0rSBlH96a0sJKDaUwkmZ9zsqpR15cOfK7YC2Z47CASgvOrr
/EGKSSsSdHwsvxaOkJVbcQxSMk9+wa6OpCs/7OAp7UBwVQFfwpRgBOwhIIssjAib
zfxqh07NUjm8nuAQ8NCP4IRFOKEUBynUyyM08HxVzAhaZFX1Fms02f44HBGgADvV
NJEEtDLN9wd8NjYmFurffad7ZMcHBFjkD9mNMZ7/vPMxSv4+RTOtFRW8wZojS1sr
z6fmI6zhJF7dirJhKVufwc0uL1N+ZkEQO8M9iuc1ytqX13Kh5LblwTd2QhPjXK7u
sFx+Gp6F61m/xzL/0yNwTaYmoDA/CfsfMBl2b6wKUFKRpGydoedjJNAjLLjv2y8K
48ywuORBY4JhUpq5plrl3BSDuPze5AVfJIzFSk43Ut49+nxz64GPtP4CsBHqdeTb
13TazzZPZKz/FU6hFaTHe5pRmycaFaeYbtfRBX4JPviwsQckRbrn6k0BazCHjCvf
z4JX13TRcvFHausv2dCWlUDj+P2zbus6GWNvMRsm5yi++sZYI6kbasszFyFm65J5
5+v2gDJkXJy65C1N5brLYeIB3UY5ifxNVwF4Vhxo6migVeQxf8StlODYLSp/ZgZo
nETea+C1aHmSIO/MZ5jla0SKXGRpKQiu259Tgb8vSetF67dD3mmSv1Q7Qecvzxc8
Vy4XhViI9hsAJWHh+TPDgMlK1kMwEG3NeDk5L0y+ebXqqmfkSgNvKtktQ2CglQ/X
I7MrcW2rU72oJogUnTcnh+d1iFueKode73n/R9xGx++Xgvtuo7blLq3psEpqfEuR
qbJ6JzquMsZyYNpqcJ/wWUtkIu61MBwSpU9XAyfHwkxgf5kUwSdvfCnUYvGONFcy
tqwI3cVLoqBlMFuofkAjIbRA25tXFmx82pzP2WdsvTn6pNBiKH110OaWqGjwefTz
4a0kBt1IxsDlMArNVyoo5KPjl1HFTC44tF6ECSbrl9qk4+4DQyRaU/k8j06rDffG
a4SXOfJyebUiGiIWm91a7MjzlMvaEAXUqQPlf7FcTyqErR4gUg8vzIpFE/QeUTmg
MErFQN42yFriIHYkeQ3URIELzWfqKqSGYg1RFiWOrOAfaZjXfRkPCwAz8iCH8B/N
utE5VuedjN8kpGU4ISKrdn/9BWR+NRclKFvJZ2cFquB+PO1rGmk7OWjqZloFOZjD
UIQoH82bP9cozPcmD7OAVFqKqgMCegsoL3eDiwYbcNzpA3u0hcvlsS6lTk0U/C9O
E/KctC2ApKsHbJbTLEihcswoXoAS0Z7FLVSBqaQaFKqoGowBdLDGgh3VPQn+OSBk
nYM4TS6kZatY7HX6K9HL0XTOB1SFP/LeLnyeRBnRIGedNSRDtdEFgM7fj6MJlzun
6GEKcqLmJ9VoledyYY8QRdfNHV+5DKE5SOYDGmZDxbRHrqPgQSocV7ZnzkDD887Z
Bzm1C+et7aNUho5nmSKJQg2meHSWNmCJSyT1aPZYB2XN+BY8XPpP9JPB84yYaMAh
8GjcJOyW73kAeZR67qOybxaNBqcyeDBBnqKxPgnX6rjhPlLkPS1X5jAaEaCrt57t
SGqUcBnldGrN4wLi7HPyqJmO8HN8B3J8H6Evpb0bweaRDy1+syaA2uHvStfO62Kn
wCLwr8Gw4dmdSpbmM7kl570wzgfUK1nH4MoIHsI+27Fts2YcDbaNpMz3s/f005Od
Z37bm//Xg+gcBO4yeSD3dHMQg0J/NaadZRpe66ghXhDAqlKlf0A5iXP66xBU5hdu
wya2BDKQ+xg+3+CWAI+jMFiwkw7n7MpIZA/ebJp9jpZenmQlBL1xtyPxsKWAPr6F
7eJvCtltkWwo+oO15ZuATvtKmFBkdhHwS1iPeBEW0jOVCOe/yteH8wFvEPft5ynR
7L3kFpH/F1IkllSiEHe//T8vLMzropwVTAw2wCAa5R3Q9FgmoyZD+JsdYhEJcAU8
oq8sv6nZisoqJIUPTSBRPiWymuOinugsrDFnZqzd66Mr+HI2qYfAIHhZVY9X//3n
sz/tXuNtmaak7a3ZcgLcYAYCqyPOhHfd5+/nCqPUnI1ORzHKEVE3m9GG5auPdrae
xTTAfHJn5aPryNauJT81pnS0XaEzQpTgZlL9/ZQI5VT1Xplr49ObbaP+wBQNL9A8
Tnxst4PCuxsF4WWTbsBccTcusXZOHtTtMgm2QwBqa40Nxi2x/IgmWCAZyyQQhILz
F4ON3fJau0juHWCIuUg0gF9c5OYhqemY9N8E5YKFx1A827GwiApIIrLftx20d0KO
sdVfE2uGKPOJzHqemYsj4sAU8+Si3WEEWPbyD+/ZG5/yC3rHmAwqbv6X6Lt/PbD+
SXk41w9WSS19c6Lap+Us/Sh8HuiJK/oRoYo6IJqmWEMu9vWbfgVtlNPR1iNy9BpB
2crJIXospK3lb2eXYak64/RzLJ89e9GeOVDCv9+eOTVBLVOUvUAL60+NBdtRgwW6
n+oQ2eO571NLWYBB+QliMo/PpmSiiMCs4DRJtH3wBnGZAyTs9p+cH0NyZ1YsMwNY
c2fXLPgM0WNiQOKDNlnneDlc9929P9cNOvdhuyZ29WoQb9HBQ3jd0XQTCSAhuhyC
gC/sSPWtK/jm0sRX0TZh5YauKBeCEzbuxn2oLdVLVh/KucEs7xH8Ft7iCDiFwm+5
L73AVOMv5het1KvKoIaSDZaYT+qdEPfwJvtvuzK+v9ZNo1dlbY2DJgZU7AD/P3bT
8fa4Nd1wlV4pg6ZSVyQyEPhHRzgpHkCrnl9DblkjYHKbjlNJMZBsAfUfZVfi2tjl
ScdnnGVZBCOiXB3bL2P91RLKEiaY0NnY73sDn3c+ad9Y5Bh8Zjdx6CY5sD+KD6mJ
mxKHePaXMr5M0XuB1LZV10mn/9M57/I4UwhsYKCmk/XDppVL1IYbAUeBd32KuMGv
9cMMaZHbwhwKj+R4aAzC7Eb4/9CMjvjdFnyRYmAWp6pRqB1kVyQMFVkywjXwuHiT
cjV5Xb0F929DlO3Um/Jkz+AdkmcvP/ZyDMzJNotTL0HcXU/3BXSufShTBNfjCfha
HtdCsJxnsKdLslJ/Gq22DK6fa8+qXSpnpSwuj+jf8TKTwYM6Q28I8jfLph7Y6+0T
wyqeM3zi/mwbyiUDFcj4OpXtTNuzS9VHzkgvNLvAuNeOI7hEGot70xN9SSLelsA4
++nax8ewdTc1zPvsDYDPEc6RQEqztv3qxSdulBKzEOcc5P6sYHKzvaxlYZSyylXh
l31ka4ZJXIGJ1m294GOixGspbdwVRWv5CAqvxfzzTwi6WVJx4Z1x4u016IPn+xFL
8B9n3qbXVZQ1KeAZRzvhfXNuezDXt+xVA7haJh307x2kVkFR4l+cv3bcIKQTwJ5/
mCKXESaqGi5Pes6s6Hbp9pXhQ5bKWdPQbIfaJaewHD7P2CuVeTK+YyxpkSe7/f4x
NXz+7O1oo3SoIiwjidVJzHzEAPd9FBv29qsCoHCs/JLkoeRdqTx1SUq9QO0xwI43
QuCv3EFyLA7mRDtZ+oHN5NU/UOLeZh6mG8Ep/IIOR0ISIm22gGBXrDwTlL+Da5eG
M1xMu5NdWZFyiBEzYxHpZXmYiVjE6nN1RFg+kdc59a+K5OhtzSs0kVRK3hrfBbv9
Aiy2u8leSzmVHThdSUKu9n5nI1lmM7hOQ0phqLJKDZAYS5jXRQwFbz+bjMKV+JzY
9ywYR16dbtpZkf2n8YTufwE+HvaIDwA5ckh2UIpI8WoTF5NrjZPl/R8CPIvXZ1T1
UT1TDAVqF3TqwnlPXJGmDgicTcN4/dWVpz1/Fu1eEexeCwDnnnv7cWgwoq3g6SYB
RcAB1X1aGjOD1dpvs+djqkGR36LYYq0L/WURO4I+ZeOsdkRjLuPiCVERsCSCu1d1
npkYFelvYGYJq+mPvDtSYhIFJbsB4Fi8iFNn+oegSif0kCqiZWLyXkiP3Tfw1DC6
HtFHG/W7zmnMekGotueCPT92dTk5x4TMJ6uaIsID/fgc4vtfnKzqWQoworbFlcT3
c4mW6KZ7sg9JkybIGMaPt8jszF7Ink9Qtj3HzUftb/NPSnuIT7XJOowu+ebesvmf
rJ7t/vRDpsZcccd0FUHoQa6FVVZQpo4b4tX0a5KpCtTIlAJpRKobUnh+KrPQtfde
oelF2SHveK3Mnk6ZS1EWpB4zkUiyqquVOImysAfDhddHPFqCBAoVKDVqEa40x2sD
bNE4/HUD68TdAcySTo9R1H9Eagw3+Ni4sQP7bWnSZiEosIH4UiUf8AG4EWh/rows
WfvYChV4gbaN67sTXc/rEN70LkUQ2LG4ac7SADIyUY2poL+2tRGp4qKpFNXaBuOl
K3oKvlCdSf+XnvAJ6jqxNqMX8j1ekcg/o49QD//vXTU7Q/uQaeP0f/LmjK6LNc2M
cbgipL+XfG7aQCndBtyA6UcOGwOyNM6ydOM9FoYXvAD63KmTOKd3ibneW3Krc89+
+AfBt4x8rBI34vVZcOsBc2ZJo4PcaSN4/tSzC/OBuBCO2gA+3aoxW/f4OxBFJucl
POi6zqPcPqmygPglR2uyTeQRg3NS+P9Y8BE/nHr+b3UxgSps37+WjFmmaavY5MXg
gPt7pL6i1GaIw81jqI8Nz79AiZNPJ79WkQWFkPjqa1S+WPpaBf3abWG5Rm1/oFu/
Zh9h1teQe4IlZ8x0C6WQS+u1Wy4uK7YSqQh9ENgSkvbr7VPdz2jBZOt5K0P7qSWP
vrE/8cURBqzWRi2QkJluwuQW0v/dmC0TiP/OCcrmXSnUIYO9xlvUXwKgJ2Sdgkaf
WO9HPHEOjSsc5kkWzgVfLLzXpN3/JZFNwHr60GdqxEooUlUyCzmmyr5h+W+Y399p
Ert73CPKh6I5DvDDvUvQMGA80HefondJ7JGmsVcvkGwdqljatoRjwtHYG46pm/e1
HeiUABGX7wILc/s/z1oWS/6OrZOQDyHOuoaTHoDgvkDDMK92nVuOPw8tfBp5MnJ5
T5iSTD+7O7hOWTJA6FZH/Ds8VAFZVD/bbiUtGyF0uc25nV5129KubCfB3SRq6Dab
FVttbTQvaIQUHeMZltvgWTvGIdjMKJZTdo5y1fXrwv4ogc9Grx4TpvHL4c6oLVJ2
xjOEkl/kqRLV+y2sRND/V3PLQchZXVXIJ+i1HNBDSA5o4NvzP97BXxW0TPfQftiR
E1PTbG+2SPSsVPE0bzGy1SXdfA1eDx+VMFdHgV4uH3Y1fodbck95g7je+SFb31FV
1P+ecUAe20NV/PQHi/2UAyvxOy44sD5tDcd4uPh+ZaFlQfF0GWvGkhZ/KU1YTAEp
JCVlvF/+yDHSHvm6PJd+XtDvPqNtU2KT5h8vib+742qSLfY3q9ja92udTomtY7My
xAPk4krorVFBB433gGDLk+uPJgDa2REqFhjWhK92+d5bpOhn6xbWJ88trDQXVFJs
q3vu60UL/pn0DrMeBccLUWHduK1zPTbOAGCX383w0DRmoYiXTIBdH2a96OiyOgo1
4pkbmzZ+kvrfYo3s+QTh44AGSCp3ego7keAEETSFUN8AnO0R4BA11FU3Q2uvhuia
Sl9f7Knp0CVRXzrqXV1DaX5qj0T6le+HiEv+yw01kOgEl26hJhdsroBFHUT4RJ9f
zMFJsJdgDxzYMpnT3D0NnuCUi1F4UsUM8N5IPn//0MvSsSOUrf9I0hjFdidm8smn
J8ZO2IvskXF+wX8jb98ihMT62Enk9kUNgL9H9foFCaJD2yn6Owf0FanCRjtWP4Hr
nLUtShcYK8LB4LG8U1riIftnAlUFweRxZCYLwMzozsEHByl5ffaw6b2R8vXBSj0R
UCUfpwDFeprKnZmiKXgJ5R6jrvvJ9BHyEGz9Ad0zy3htOTMJ4MtPTTGbnjJfCKZa
IilYCWMox7NJIlJ6qzfus4Ce8y6gQnhlYLiMLXdXDdk1p/zzjFH4BkfdN/QN+T85
pyoiGCoijYSHX12RTtFcmQzNNsMIC+S8vBoUY9cw9i+wuvn3hz6f1+Amegqup5GC
E9bJcnN5jUxykOXQsipALcembFQxuDGSA4OaYHapplGC8NjPISWRNIdvsfq6HmiQ
OTRchT1GMeZuRDJnAr4Tvv9RFWDAM+W6h64FCLP1Rc8u3wLZOLcilv9CLULJ0hPg
kPlsV7QnK9odjSOeUHRP3Wz9OJRpes8IW/7dMEAP2qWjQtfWIDlEro1yuGN6eOyC
92F6MobWGHYlgLjLew6BlZv0kNKGXpb2l8zenuQ/imzrV5mV0oA4t6CScpp/FiCQ
D6ypCsIvhgRBLGf922x2bq9VtBjfYs6p9Sf/BYCsWYvTyE9X24+XC8GRjMq57eG1
RvMWUVz/U8z/YE/3yINN/IJTVQmErRvatELUApqJjDked0O11HUZY9Po92N7svFj
JaxXujgsUcwhObq/XDQZuxmY6CjwS5T+NJrn6Sl3MEuh/0F5YiyTqdhGliBcrvmL
Kkg2gCQqZ92z76hWKLuHw4NJj9oZja/bxh/1/Mdf1Ai8kWVb7flITgon76g1FIxc
HslgzA7Dm3/V8Vod++PX1hO/ftfdQUgciUmtcQF+PgY8fsd5FJbVZCFyt+8sJslc
i54PpCq0x5gtZ40wJjL1qXAuaAHDkqmkd8XkYtYhG+tc+HfufsDlBw6DTNyvHbTZ
GG8jzrCoo53WO9QOyv1hLklhOXD4xSk431Hpi4C8FSBYhwyIEfmFUTsu21l/tzgR
in+l+ZwLcmTvZmGat1OJ2JzPKBOX85Z1YG054eGC0QEpwD9kcNYPqNmOBxvYMfko
Mn46GlvH9v1rhy3vFSNp2NNgqVTh7b401H3Rscca01+mDNa57NCucKu/mq5Smoyr
g29vxJ2nGqwp4Ex3DaIEeUS6K0u4CBaM8Cx6LF7GTXzSGGlzz5iX1iWaFygmastG
gtAjJ3irkjdSpTegp6kOPXCSpw93L2MAq6DHdaVU9+X4VF9rVnsYu1+aysacv03E
yw7mRSrqrah0HdI9XR+DksqCpk+4bXCICF6YqTtXtQcxOJlclopwuFZ54ns30c2i
EmHPQkhSQLuvGUPqm4Vo20beB0h+aDqfO1YOcwEy5S5/XIAm4JHU9OM2KcTAgyIO
9PP6g67fgOy2R6xIBr+27lFwrBZUiEYtJe9vwEN/06kZid67k6NMQvEATrbCTjhI
XY0tHzJxyV+YFTeYiLEI/sXJVeueuHuTV4iXpVtjl1wI3cJdXGZhALJIufqATjXa
qVYR8RIJ3yC79q9mwTaYpKZB92AVKItsBo3T88C3k1eBFmgJS9caFAmqlbGDQZPX
J8tlJNqpYpa4pxPnkzq2HTJbqxfGMdkB2lU9INJNvKgzxVqkwBGM/HEHrO33ioke
hezDh+QC1hh0G3xWy2KDuKsAmGCrOulGm/l2sAWIktyozGJwK7UAueJGorvVix5b
SEk6YUnm6Rkfki092Jp54w/EjDS5EgZO0D1LqF+XqpaKlQ6exKfCDF2IC4vEwrzZ
yY7IIjN1vwt+YBa9Sp+sAGQRjZweUw0Y72JViX68HxIyC8oLJpxsDreooo1hzT27
MrV42XHgLxsBpS6NgfXR/kErb0hf/3kn2iDJNrGXTUz6fdOGpZNvxb2WuzijXOg3
veoMTUtacRUv5UDEx3ikfJTjcusm/chkE5hRf2FiMysK2TaI6OSNdrqHDzsQByRu
fLjhczA2XtDeIKaf2QVakzJISOlKX5v5PNPV1sAJbf91D0InM8k6Q1qSkKHLUqL1
z1A9xwxF1XTmRR7UghoooiH/OrafxwZjO4LBiIRZonx/NcdKBuiebw0fJ1UfFOmq
qlkLEhtZroB+Kyx1BrXyiv6IDgam9v5kWbokzruodeli9wX/SXYUBTjRB+R7ScRv
UeFptNM++0TaTiTRTfTIw1AJNt5TWacl1fHnfWI7cX1fSrmZS8c7iC/WhMSbzgtD
YbcJvvhoNIxifcuJeX32rfmxy73actwKpR8EUyv6+0+bhkYjbrbuv4fjPO7f4ZhP
pos+csnF9o5QY4zNe+WmHAzrq1L22hbjEqZPsWG8zogbAiwfiu7bBWu8Ej8JUhyX
xYxnFLjMYrCaESX3MDtwj7hpyjMFdvUtMBDG2ZVwI7dekQ7qpKj1UimYI0C3/BJz
YG7aI9HqxIwQoalKIQcOL0uxTBOy+g6tgKLyDzmunO8BPSI9TVKGVZAwAI1QGRlZ
W+JbbRU7I/VJaiEcPVBAb9eVMrLgwvNgwBY9a4f1zqMlTrMUycLue0RYLu+XmBRq
XV5f8IPNXcwpkWNUuE3BrrMkbU+UJfYadyPNwrP5IrWCqZerN/3+yNTuujGtySd7
gopwqGi9XoopcltPQJQqUPHIPEXgZt6PuE5hQbDxj7l2tAGhU9emE/gKgwl1bnWf
Z5GpTXZ22XupW3ektOa7Ks2aiHvPCvwF62VB4Uegt7xkrmoI1I8GQ+diPfMC3Sk8
jTzcGKfRRR6pyYX4TSbdJMkpfxhOuIO/5t8eqsRk/91+xuarJeUNx2uoTf7UMrd5
9QweK6f1q8IzzdOlwHiwufbIwvc7kF0vs36xLeOmfIWFO+G1STIIYuRIoUlpFzRp
eyKvOIbtTaqeQpBOTTr/e5Zd7DLbdydaes3yqBFBhscQJqsq5mUpQsh2CQdQHxIh
sF817wjKLCeJJa21uTgMg6psImGtUpNcMzY3T12VOspkxA/q6b6KyXSeX0aDkJ/X
X0zPUPP2eN5IPqEoM52dGdlNEhkv+qSqGl65tkBMGk0yXz8xXtK7ZljqiMQNhbI3
0ougs4H2WHgnxpfuGjd+vl4ZPNfbhYOBP5sTa7UisbcqEUw4m3usMMEURQPNR1bb
JfjIglxck/MyS1inyyoVv5RtD6CPK5xK1pJf0lhzAEfZR81Og1hwBpDrjOzwdm2d
PqfCR7ldQYm0TwR+ono1ZTy1QNdqwN68D4K3IfKpFSxdU2NugVLOS9049UL+6rPx
YKUgzxHAn66BqFRsTUetlIoHIoANItDw0hLar3LCyu1fwiNyUxvvqZVD9RfXorAl
8/jwC2KnkZtRO6rM9+t426t8sJSUSIbMpnyApiK7TyyGnsJTqBKULbIqM1Dxe3aG
X8tGi+1LsE3Rf4croU9F1VRLjUD10ncA0SLQM2kIw4sR1zv+e8M4SNeuHROC3hFK
XsPNL2u9U6zDsFLikNrq6hw9BHMF48Gl7LvIY8IundBv0T0E5bpvvpOtB8pg2bZX
828u99ouTdQLwpgTmy3TZfM/zyWPkGf/NCuMb98G66uxrEZ1Cl0TUQCNgltXPGWm
KQAhxdEaVUYKnRQNr3sC6/whz583dBIJylzBJUgNgGf9rLzNGor5AgM4g3swiL6S
xKzSbC0SAi1fBlyE87+8kfOPehWYlYlOS6TUsS44IRfML3ROQTRZAeoYMgPnOFbf
arlli7CMm5AS078AxoZcZJwCoL36JB3lvSOyKEKSkmmKEFcd+EX7uLy/CmnIgfgX
3nvPJNDzUVGKjm9OEYlOrDre7VTbuh7PxMA+TQowZW4PimCvdszKqMA/ITw73OzY
Q14nkJ82WsSbXpY6rYU+rH6nxras6Jr8uA1A4iQmMn/8OWDs0kwdxFW31HzjQBpp
V9EEg0muam3QD9669pJ/hbGF3XF63+g9WbsHsNlTWDbNpqGjFTRNSoIsT8+p9BC7
puR39rlaSE8F9k/wjd3cvN2T3ykLpmGKuc9GfRiMif9wgiDEx8wVT6kE9gBwWjlF
FVre3qL9F2W5n5+w+XdW6VTV5wis5UdjuwqTM26ErKPtMgWZXj/yOqnbGCR+moy7
6pXcS7ZuoVKrf+Dq+Mfpc07wt9jAwGMvKb/Q5DBtQv3pW3RvO2tvcpp93tLg8nvn
OLXNuNGzICj5BIU8oDC64CwV/aIf9IIiO/imRremxpJ8EPU93CnmgWOr8N36uSj+
M7Kj0e2CnedbJ2/jgGMU0uB1NoPuXEm/Tzisdh7L9MsJVBdw4Sxkji9N2IsvDlsk
BRENFygcLBBWF3dLkNRcoI00gNtHsbCSXALtyJrX/al3sAhXiuFStEnUhUA5l7CN
bpGyctpkVgW5becDlOot1SruhCybiYs+ItkN21aVNHyrc1+0y9vjH3smXuHmEfrJ
DPbCI8GM53kT7UOEAcf2RNgdm5Q1FOr6ku8cIgyVIKCrCOf/Vf4OyVQ1OUPlU0qj
TY/35yFldHa40QH0i+iu4h++mTjMcimyFkSHf1AohEwjXtq/yW+ZElkLo+9kPWOk
vOqxPHQg8NPHsvKqbnTBepmabzFwXRnmqvoknK+SNpHqQ3ozVIWPIRskHijO+lVk
gRhnelNh03UujrnANy/ExlIk9dURMW4LDcqvRuNao39HesBDjrOy00v963a2i+QM
9mtH48T3k4u9y6Da14IsdOE9Yh309vf1YjDHFmbpb4XUjRIuMMohVm6upuV+Zp6U
H4GQJvdUjHDgac0L6HOveLuh6NW22C9MPKMEfvpatt1AtHwT8Bq83tQLlUQhde/K
RmQebLbJ+krdT7GvZczxWfEppaGewfuh/Zy6Gk0VnM7RG6R+b4w8m39QehxvEFPW
IeTghspLmQpU0L1aKbV0cs3JE2trtEWIdbJqaw7RKhvOITKTAzEss2FqylWLMPkX
LsVfZo6XtC0GP6lOQxiuQsuxMLEwbyIx/yTdAyJiUt3Qa9n3smCSXc9Uc4U6mQ3v
e7dwc0oKNDH4GD9kBttA62FLaxAiyJ/oxXG8aBf7UOLY+DgpsBFbyvnkdW2ilQru
oNMIjf+JapSq+vmioaViVDucR+jbcLBmdqTiSplhK0FOV1R+n1LgC4jThUOnAnFf
0158hiR6Tdy68RbkuUJVzjlVoImjSL5fGUIQbUnLrnI2qUpbcT1+JKoMFG+zLM+3
P+khnjQV2TsdQkc6GhhQBS5v1DrSNbLxeTDPht8JoMhX8TUMTCrmwJP8jJMosHnx
5KMe2I/6ptBZhVwzp0niViJRaCFwy6oagiH0KPLDwTkRfvnZolfI+LzZ4jKb3egP
XiBpc2yWY94mOKNwqBRmDd+ZU7W+Rcvf1O+lRrZhwggGeRZseH44fr9j3teoDcM+
e2Vufj/LNAt0HlKtPTMxJpvWFVaxtmWcqgOVLeeGWuj43cYs3zbubOcn5MEu8moh
Ar8YTtuR3JFKG2AJ4YSbvK1yOGtL+WAF0h2mdPbBd7behRQiSAgmCWThMmNjBTBZ
Ap8HW/AEcIi9nIipa4Qu/0teijCx0PqsHj/7h76H4boTRDZs53FckZxXmmUEcTix
WePY6wzcbTG/X0fyldkBW2pnXl7IBJ3fruY/HTeku2pnSmChLiohsi28G8Dmb5pN
HqgRMCXhzHsEi+C/XoXg0zUzEGyB4ddnjYWbAyEbe8i9dOdeRB0F9LUMSysfv2fx
UgkphcFJd8xHd6HuCt+89jj1qXc67gucQYR0jYfjSKnMcHkX957GtMbX0i3vhpxD
aT1aOmJl1hZRf+DMPweRA/4gJb/jXqtI2qXE2y8MbFv5fVIUZyPQAUfcjheuQlgo
YDfKk1GeEvGi/YE6iTlmcVhi9Xq1DE9NQYej8MoIemNf/pVsLNrQJUwZAwUVBuaa
vOcJy60Rv2cCLWdouoSeksRsB1dXgefG6ccWD69e2ftYAZxmb673++7un2OsnaYF
3xBiDsW9D3EWoBowYH+LdwxfwxnUhKqUZUHDU9vYmkTnjnnyoh6dlzCucj6T1yQs
xc5Ij1/g2h81f2qIN+6UTfvTmoz023YXA6gsZ1jn50tpRgQiRzFMqFzQJGwIbQpt
GWvsF1I7Pvm1eL7EMchQRd+LS1zbfbiMiVVYfDFCPaoLY9+vHNUfgWYmsAnUApap
kRIf6CTJHLCjqgh5rL/ThbYCzJPRs5W95VUgUXkoKJRwB2EhhtVprZ8ZIh3J+H0A
XNqj1GpMx4RVuMC1QTnO1SHQ3GS/3NWfxhpPGu9C45DB/EAlBBdBoXup0zNx5Buc
ol0YdDX/X12kPGAOBRtyLYVlvwysx2Yuo6deRefPBvSOO/9mnyEFszu63it7ZBoP
ZwC7sUBluej9EBqjoJ+hu1jqrqItgUiLAtZ/opwPWNcrT1gixjvIgm57KQGCZmkE
Ut9BfV6B56WVxBVqFBF9Yjr7jCsLlPzLzx7Vkz6Retrg3S7ZPBOsZvdiYfie8WPK
XBDKLjpW42LLUL5dmi0fNX17NQXGhB+fiOx9OEjNMEVj3xRbk4NcNDluZwIlP2/h
kOqKmgLKSNSF4xZT5WOsozKKaxUGuPG1S6p4UrYKQ6a3b0cmi56rW7JjYvWwQW+F
i0ERcsg+bcMLGUJnzkqM8UGrLuKyqX9Yj9ctLJwGdfJdFWF3yU5u8MM2d45W+l9G
U9CoPLT6cXOOEYtpEmh5yH59ac+e2QOoba6uOBSaJed40Su2YbiN8fKuvygcRlB5
Vkhe9ObLRfX+o4E/2+P3L9Vj5/L4X3M+URIwE7OhFd+MS7TDfP9QNtLuXoekkQJ7
dXmpcJutfXeuuGQeJes8W6yzHaEOD4jM9pJWtgRtkt90dDQfc0SnL1dgY+sxjzyP
J0kIS9saPM70BpuE2E7y4kpCgYOp0OLMI5nd2KLuEhUHOM9+dcceB6g1+fgryyF7
e78IsuSGEsDwqZ6OwuSM62kMRDzhTYS/x1vuy0laIs0e8wdrzZPtuZfKer3kwgu5
OKLIZpyW94faEkj7qcmoplOyIM8aYqB8FsOQc+mYa7KmQEZRtl8LiSfFSPDycNjb
nUDyP2aw2RUzX1+oNGki4fdPyMC4Aem0xJn0tljV7vE4ABphXctepDupIsQvmQMx
SKVFqSzQ7i1+bmjEmpUdjOfl6XSUwcO0BfcxTGhBAoPTvMQxqzak58lQC7OefZ2j
XSGcBXq1+Glq+0p4AEhli+rCRQ81Zf+nj5Eh6d1IDfNNAl/5zziCdIRoK3o4EzQA
jVtd/7Sw0SyMf24e3d1ge2xXS+mALVylU2EMvOgFJNewPL4wr1333gIbpeyNfcrj
oDAraGecXw3fVGAPx1wgAj2CMmoi9NjedpsL8+iBC1bUvXMxCCA8f8RrM/9DL2Ou
OZH3HUVJ6ivS3H+SNA/TMGTe4FBAPPqocdRSi4n87VXHpVbGPPwGAig3StR0IPKu
1lgRi8L6VmCZf+R6V9dB42boNI1w0KWGivEMekJL5WLBLj74bcoQ3dqT3QV/+Xb8
3JcqEJ46a7AZVGqMt8iz3V0pZ7AwuaaaKP0VxLli+qlb1VrPRcikLeIJSA33GfmQ
Aizumgv88R94Q2O43kEvvCRHivYpeKyPpOubIK0f6Vu5IFZqqAqi2dIpX++f1XoT
BoaclYuqULIZXjAGYnBRBCanpN8sI66U/CzhzPcEWDO+Hp77SvUjgaIMaVErfafr
LP6qkEh3UbpLXPpyYRun1QkM6psTf54bsyAjmQD03REZey1tYbhlIaioyDY3gWPb
4MDSSTAHVnkJr1uKpc0unplDWSV6LV2VwfTA4qHfZ6BFAeSfR4YEpFdI3lxGKQxq
sctQYsPH46kWQguX/AuzuLOdJ7dWPkVhrc6xionxEK0iD2GpGomkmR+4Rd1nRyJ9
/hgzSGTGphM5OxvloWtoD9LzimbX3Vc18s4d0V4dTlFpeYg/toeA1/+d/Ot9b9Wm
D6a6Xu2R+t6J/hm+Ua1ggS+Q5uCbFIjzPcoRUIlWKKIBaUkE8HNTgF1wOIbCtoU2
c90EWmVCK/yQpMBTpv3P9Q0mospXAIV6cuxHWYa7nrFZT3VtIiVBRoyu9OgJECdG
plPY6SP9alrV6jcI9pli5QFIbbYuBaptLSi7TDnxURKkNEQQLVrOHyEmRBD0BczF
Tda1Nm1BcYOfqNcHBa7S4Kft/FEugvEIcULmon7anGZAVcOAWR06BGbcDZcpgaGc
CPS8KCqVHNHPweojbVSi45m+K80hLvPYujG/cXjKyonBKtjAhqMUN6B+8I5DQPnb
HHzwkaGIk1tgvV4Br02keKPQIgi4cUEbmRT7vgtwUgVNWyHGM9omicJl4hAKUPX/
VY2SgK6nUAhonO+9h70AFlPOi8a9XzFVLeqoxeZnwfrJQbYsrQn+VAC0petlV73Y
IB2Q8+rSAeDVbC5GaSmAZmlFj1VXrwK+4x9JTokAoW5blKQ3Ruist9YYXdNTZH53
QXtNdeFS8E//bYWLtCp6noF1mPJ0k+ztB4M5iIg0zUyKx8QFm+R0cL9ufYdPgITX
mbA+sgAV/4nLAiJhG10kN8W5g16l0abC93IvVGcV7iFqoX+iuP2PvH9bWCRk0SKu
g2ypy5yEQOK1S6tEFzbvMAu4f2XcdvZmT3pCi61KqCwqLsNq3n7eKtssfHaY3Osj
XNoT3OSDOkZrPGyR0+C3HFttscygpHyHfPDuevE8iDDaE+36gy2Xri/wlu6qIyx0
QsG+rdanFNnPPJxz7ak2WZ/K338bXsQxgatfi0kDKF351Fqc8EY6ETBwD8gKNAn1
pNRRgceblpEN/Beym1TinCStinW2h9O7o8xcAHKzXPgEYbvYJscByvlmpnwZTfY7
+e0QfcSEpozEEZiaGFNM8JyjIjrAzlZWoOBi8fosTOVqTRJJiaGOa/E7unUhyhcD
p9tvB22VWRhf3wFlTu13QyrgL7kqsUOUsi/CnH6ZNNA0CW+UgMGGlQl27y8eaxfn
7e4YaJcIvjxNGuKhVtdf07w66+vdUUmc+Yugs5SweL5m/LAHW7BVoMyBPo1RwhT3
yg+cjdD3S+cAyl2kqrxdQvu0kH+e+BjQSxxQ46BozBEYt2olv88hCWUT1w5HB5Bs
/kWkSDrcCw00H2aUMq3thwSaDTjOjDngOOdr9PhrEIB2xNCZkm9R/oRw5oeDynln
U5vkjwfsUl1tcKRnsqkOTIVo7krw7DIIILoo2GNOmiOKckjJm6PUHhwdVw8QUana
PFKQhXE1iKZwbRv6lFBfMwD09QaMdrmn4IjPSFW0+abB3Mq+pjyw6a77iMt4ngAP
kUUiuhTuADXsUJckSHt+Q3Et4Q66Ebbqifuua1OLixrc9FeNXGtRT7Ukj4FYGpME
b4+ImTHyeWkeTk3x+2CY2GmctIHsrOW670ZWV7Kuws2vOYn4Omn06Ujs8ExEjTa1
h6daJxKU0p/E7PDPaNxa+wlnC8Lc38PT5O/3bjfRO21Kq2Xs7Zm8MPPxhXsf24mg
5NNrVzlLr7isp8a/POmFjUSD6K2inBooazKx6DV7dMz57cchV24G3rzYpcWGX7QK
3bNtv7hQkoaQLCxoeO4alqvNfnnDYuOKWaSOj5faVBnJZkGUwokSjCfMIVyMAM0e
P6H62licKlB/g+f2vQ5ogrnid2gDZhbAI9xNWOeH5fdBrpCKa3Pi7SdC5y9Z8xPT
w5UlUyBGDAahbOwUmom6a1G34gwkfjvKt4Mr3PuwP+jtc6ijd74TmKkB97pCtBHu
Iee5xnorZ4D6uXv2mWStr6uzB9JZm2wI4lKhtqf7j3lcfgXnEFChTDwUY45bMOHp
zHAsJMNYSvwegGov0iBOOLh47+4NJxicYAEsL5CuhPuJwpjMMz8lotSGPUtaXWkH
uxFpzpHzoCeXm/pIdM+q2lGYRMPhc/NELaSB8uz52B7CjuPf416+tfvGZapmAdS+
6mMXGPb8Ea4VaX/1j1YxufvVErVNKlk2hRgY7clMMoeL8V9Sinqiv7m7RlloCTsr
79PcGIfSAmI0Drc0rneSFOz8u7o8sSZBJsaiq3RgJOo2PJjfMXqe3apAcZHdQLK6
OfnsnLAjjVuFAes5BeJ04F2gNHZ9VDCTDRs6LvCK3vs6EZgWS9KjOKv2jqeBw/gi
SvNWadlOnPMcE/pfU8Uvht95HGSU+dvc7OWVNRovIn1ZLn5JtQwGo9p1orGF9wl+
vpTZJJSU/obtxXcrPUomFSTzfNOlhxcBRPBn61J/KFi9yNcSxa1dSk5SslGXH6Lm
jRTINwL1TLD4tt82hEwzqUmtqknDguar91IT8xJ+b41O6cTSk0br8QnkD2yDjQ8B
bmlutSBg7MkPhX1HyUR7vFs8lugFth/xCBPFGWzIUp8S6YLRA1otxclI6GbJqoqf
R6gwGkRBRjHkz757lfrxUNzssZcYplOudFPG5BU1u1jHmSFrEbdHfeGywGIAlZyk
n8G/ABs8xFwOEjnZ1zkqhdOl7NZlsttQAvpNabH74WaJN6YtLLe0Wf8PIHE/yb5I
YT1uateg8f3OaahYm8RKtzi94GAzBo3iXFzYGg/TPJEm6y+UsEdEPuYP3eVMIGIX
gSPeoRtJXhVx/JVk33bCJpeUNNxKoy9P1gywUafrD7rXq2xBAaDUm0YFpZnmqImT
NW/IYtY9I1LHtDzkGistSW4ADsBLkCKL/jbYncoLvwKJ3NJSmUSA8hYqPXf8q3x5
0ILtO18k6duLYu/EwiLa4kbj5JahW9IfD9ARGybSylFNhOK9W1fQDPT6OT+eaAaD
nBHpKW7ErQp+MpwBgXcwnKsarXNgB50Q01JW5lJvfhx0s4DAC6Ubb3R9kpBsEfvH
MO84kmKEAvfMib2s5mJObl2LqxicnnV5icm7Qe4H5l+WRuHpU8DWUWXTyq6TR6z9
z92nktkgM/k4y7fjH8M6ddoTepvK1G3P+8+XSGXyKxAYrHXJ2RUngUJhOAqCagm6
tujWe3wGAJb/vwV0WkGWSuxrtfEYDDQPHbL6Io+8adRv0SIrvly2LGGK3+LYMlWM
GY4lWB7QXGRYhAmiCg5SqcbAA/1Ebo6coV3toaJFWoWi1WmSv8HeSj5ZVEMcU5nQ
oTngFOUGlUrLX+B4oKjdX5ODlaCYDvUjgt35+VnijODsuH8C+S/3z/YH37qgkBt9
oAiPVyRTnZJZDVschesm3XoNVRzReY6w2JKzomcDpJr7HBkLj3dYiI1WuqebOrUm
7WGZzqB0pMEr9BbkZG23KQqXwajRc3ybG9Aw9I77NkExhcg9TX9AX/R40Ujfa1Wh
o5DITiHKnm3aQ+48fvI7TyJhpT+jSlhRC5UhuuH5RV7iX60N8L3EwADoVhOApjFC
VYbafe+k8N1KbMPN26HNnjp036Z9qG2xQltoj2yM0zDQ11RyHDo/FUxaGOd0RfIr
O0P3KYDkkjsvkuJsZH7w7zb1s9bSZfkC+1sDcrMYhKJkHGyyQVxrHTIhpkZzUAlQ
OO3QOs0OXgo6g2z1jwCw0k5s0smKnM9qxZMLkordXXZIYb4JGUxqClIoK+pWMH4k
fa30QfsPMp0gBrsnuLukB7kaoSn6HAF8J7umjufpm4xoq2rnhQP9x/O+SbKBnMTI
bXFK55j03SqF3U74/nLmgw5eMLNVT7dxMHS/u7Y77sxkvaO4wZTSq33xl+QdkjbN
SU2SNwV25XUXqDT00bPI4CZFcwVuCGJZHryO78Aorfs+aG4xPSE37VlJ6cVpkdCE
C3XCCb9wN+bm/shpi5p58j95urynIjjbCcNhTgsiRoMuJEuq942nwrUlVNh9PSKB
zY1ljEMZlL0gz0oB31AEV/8esOoUuCsqFbAe5To3i5zC0awzYi6xT1v96fimdC4z
ghe1EKNtQ0LFCNGUU7n7drZkTbFKfqsUjLw4loxcvRpE9/cOegpxqRkNDnpDJ8tI
DIjxAgMXSDxLhwe0wu3Ez1GfQCE5Dqu5Ylko3q2B/EpJoIi7wXwvNe7oKQXqA3+z
rO8XRisv8RJsPrauOan/v6c9ZoDSbOOXayHQqQhYkR13HDInZnW/d3oefyqg4lZN
u8Z5Hd+TWV/HuHgA1RGJurIEL2mLJIv5FPzh9aCtyT/acsU0YHhvr4VB1JrKQ4Dh
5M68+YWFLRbtH28GQ9Ei2U7U2itRPclDHyfUQqH0eeIaWhenEceFVzRPQAclwAVm
0+XjjXthouskS/7oMMv2u1EGGKSUDJ32QH763rHgZtZhBc6b9opTjqe36+qCP2qo
nz9+DyCZb2p9ESxqoRGiIDmd4l8J1NOnSCIQA7WicttvVHu/3z0GGdqE2AbiWxUG
hj81GtDAovSg6+nRi93fb0McUJb6YkIUlcEWM6US+a2guYq3pdxD/pqlEIKKal4n
9VSbPeQvFtyipfJphx5Skf3a6NYpbgzLJUWHABPx0Jcjefys4+hjY8NwJQH3tzHM
arURFf9klrR1i6jcIG8to4exy5UFbY/EhFg+6j+kQlCdWABJVTCUlrxTfQKMSR9N
ZHK52gA902xR1ZgUZctG+FnLcARmhNgyDFdtoBBoR9LEuQZDyRm2/tou+fhwPHdq
QlmWc9rwaJEIi7Ipy1MaKkeKGxkwHFWFZKYrn/kILF0uRhwfrZIf+qKiITS3/W7b
YNwvguh7Vksi2Uoq+Ej0del9TEElLV1Dv0hF+oXiXkvXOzDdNTcXaUDoybfK5kjh
Dw75aknY923O4mmL1mGWY8QCGtojlAK638HILUiNkUMftZ6NSjyLuhX/QsHV0vWt
Efbl2VTXhg+JJ4DPcZ4S8NjxPeT4Ppa4cM/K7LTWL8RFSRU9bJyem+xrO/WH2Gnw
DJn0gdqyyLd3Ti0/y9S+TarNgy5N6Yl+5GJc2on1aCPWAns/gFniK4CJH86oCohU
R6txkuqdx2tRbd5YDS8FbAImVRc2wvIDM5OubfwMrnHhWNLoRc1bXFbw9iKUuUPd
3smk4EELK10QW88IEC0Mc88xvmWmacpnoReeUTV20rbggdbxhmZOPdBaInubfE1/
pulOblr+2QNzsMTHhkZPkewhzG9SVZxX/3w9rxOHRZfitV3HpD6drewEH8RzEDkX
VNjecQawXG4AJEtbkgrjsRMQCI6v/NFAZK9jI4x3PwZspEtX2XdT53NUyp3FbWk5
a6q0rOKdD6y5pZQWlwFPNAqQ5uUPFQnrkxTJQZgx17n0vfIaIXpF8j5nyn1RHoqb
DZEpZbr6YJG6Uos8+ayddMvBksan46OIDIT72T25F/OMkQuKJohcmsIi+Eh5jUQg
tgH0I+jMHNmfu1ZvOsJj2EtAZ9q+YbyMCvfohB2GgsIWjUGsLPDfbgrBhYaQLPL5
TTT1gyNdoWBPh+hpVhZsEwGH3y2TB0yObiOSr6QespPIVXEV1aaLqzDuFzeLRKE+
qOPHt/5kkNLk760q0q5yMzcHHgd8ZUdcic2f2gbKEWUfqv6cISCZ6/xGUBj3p79T
WMTN64rm/1UyMfapC8P7Efwt20C+nOWb2wGFB56cznbF0AslPrT5kPKDtRwvSOUE
gOMSaZIv52kKfG2kGv3XB2kW3bIyTYp8oCTGXmhV6RWDP69jKTesDKmGutkkExIP
AAEw39YoiClv5QosrTtdR2JtlvVH/cgpMBa1z6S6a6HKVRiDMPEHLFTVsqCpQct9
PioqzF/gNaCxpCnclwYmF1mvHhGc5UNKBEr4EIoPALWXhvE8R1huHwOYzOK5VIpj
OcVaAhpjFDUxQJLqMwOalxO7h+wgQ3K8QKx/Xmn5f4B/poY6qUuO04/2bDf5BNch
bTCPcSbv7ZrD+2wjXx6Uz6YKb7KapKrNaly3QncAFM2/yRDjQ7zXjKHShCh7X7Tr
UUx7rpJgPiMf5hU+LChnTP1liN5yee3EypuPIGcZy/Iq69MHlwNBE9AjBUfuJHKs
dVO/eZ/SloJd7iFDB5Enx9D926VVwq9PeDBEMmNubSSraQI7GV1xA8YiJJ1RztWr
guvK2dfOyIwGFXGaEL8Pw1kjHM0a8saGcrA0jTKJ6vjBwWIlUzG4g0cVjEw0R9jK
Sc+FOy/jzHweunuLCb3P4FeISbzhFOz9oMMmSNesUWIFnFHlxE+RFv4NQSXUaRk7
F9gsL4M/6U2inGor8mlyZ8zSbsKYbwXzHbfZQH5P+q+7lKOv3GOerF59Lcu5w0D8
iir+E2tt/ne6y1duGcdOrZYd0qLobj2a1SXMsoi0Jjm73ctGD4N310LOR+fsX4ia
dGMHwsVO+H+T0zV2Mzv4kGdxKrVyYcR6HzDWJK1ckG/3rWGsgCuWshtNvtgpIhc3
EpCN5nFaSSLEf374kjQeNzqCh1Hx+iquQbdzjUHg7P01A63fvpPPdOzZdFX96hXd
2XFN0HDAj7E0z/YfPpEymc5ln81f9IjNt8KQRQ5kEVhXaLmW3+tMSIpJJDkVkDBt
SWiFp+ZIH0VLlbkg9c6u1aBFg7JMLN8ouFMSGut5/r/UL2twL9z4z4l3cG0a5C/E
x5wU1o3lbsCjDgZVZeGtniQOnjuSBh+vgC8CoFzT2ZM6Qzhsf+Rn79oAMFZ9kPlB
r4uMhIsSya6BSBEUFM0YvNt5o5wwq2HcCc8MTwt6avA5O0zZJ+tltVNd+pywYG+L
FoYGR0L9Q//E+cfk5dFWx8qs+dfqMwIE+ehLzZkUOf2LadPo+txf5rLTfi2MZDdX
dmKvfOMDddw9VKIvPF9KyQrET96rseGr427+00b6ByE9WmrQyzIhKgAfBkH9GaSp
nZzudtFbvVJaSOWN76kP9EpWBJbnOxJ/wCNwgg+DR+LfKQ4EVrRrpQwnDiENCFbT
7Fw4uEPyIEXEy0VVL7eXivXXwoA8FXL/AH8neD2LkUyjROMNwo+I5lnJ1YtsdgA+
lCie2p1fnscCN97CE/jNuks4FoKudGczjD5AyL8BCbpve2pIINVdGRSusXcR37Kk
LghCuS8sGelswwVvdhgT9UdKPioReRmWlNog55OCE1wUkqvVaWtNRCdwrPBmqmF3
Nk1OGoZPBrSt5QsJgytBqjGvFHWH5dQ9iE6RZk4Krxmi08aKK/H+DavasUxHgG/1
guisVRNXBen8X8N+AjmD2LTl6T8ABDRUqvYBPd+3Y73hnt8LcK/j8ekgZegb2ddt
iM8bW0QmrBBiJc1nP2RtaxzAL87I8GzlPHQlLM05NXu4Im6VFNk4Rs8Qt6+aGel7
Qfxf9yDrOcuhvHnslj8IQOfGYD/k9Fe4+W0urfCMzgeislNa5CHx0oDxhZE/S3SX
MreIcio4BJ9nUV5dVmVgk8J4i5RU9q00IRQ6zZbbif85/MNk78FlDH3eVuGRfxte
CsCAVwOX63vAMDfn5A5GrEXLRn9m88aoAd09fE1SCMKkIqmflr7CqKQ3Urm4gtBf
0qDy10Jl2/b4Ooa42lO/G38MAzzY0C0CrCYSBC2O1hXFYo1mOMy9LWGJP6nIvGLg
cJ6cdENS+UfN6kMn0Bit557uTRdiSWZi5q0q3d0RQDmlyDM4GkYxbKdKx6NFCWTq
XMq1OuXuIND5X5HP/Y2gdf2rRuXlQKlFVATFoJ/QaHidRgpt8dWrCWEXwklguZ1c
j0MjlK6T959m2nI+MtfAQkLAdw+TT9psrxnS91FoLTzf7S21oMRR+7esgl/P28tu
M0UcM/yXRNY5OafAQakEd4DnulAP6Ue9y5LCQyzApO6LBWv4XpA2dtE3Hrm/Z+3X
fC1TyZa/OlZ0jpOaEuZR1EpHMUSK1NYXaeiO4+3iZifGISSLRH2LrGJfAnMAzkLG
NCHgbHV0iF7pP1BCdK9+BHW+YXLnL+iToc2Cp2sXKwRx+NZWwRpYPI37a+rNV5Wt
Cbu7OWbqkqzLYn2axO9nXTskJW3hYo/L0cdqar/uCU61tmzPLQHjYBrDcBGflzJE
qR2vt6U4/8RSmPZQuHZB41ruFrTNWLnMm+H8yWxHClpQ3mKv58xorf7PBt9A60BY
5vcje0WCuVlfUlRiKDK47gr7CBMcGjR+7+wKsXThEG/32NQ4dq81I+GGYGVm9PAr
ActfFmEQ1kzzMAQhX27uMtxv4b9bz+g85lFPmMMny2IiMsFcpmrr4DxTLgW0w7NS
twqbNUtQ0oQksthK05Nh2EK5xGzOBuNcySo/6vvzBHsGjZkSUs2xsaLJ5YkI8ugp
ppJNDEoUP4BDy2RjSyEWmE+z4JFDn3kyySKQUrXUOE/G36PlQO9i1uNPV6gswZBV
Gh7GX9Zd8bA23PR+9yxUa3fwPm+qBYwi7sV2cQYEjQMiTP8DtIKTtMRcOmz4sqCO
iGhcDG7oH9nslR5j33WcnauMI2F4YpZTZNL6HfzGTostzkwwPJ3jWLFf9aOS3jUo
EpOoH4gqQYy7F9z/RZd2XGOXmtpyybWMolwwtep4JKYUCTlaC6+WM4cyhOW7ek5r
q0mV7waDuEPjCE2k3q4p0T2i3vh/H4aS384PD/VMtw6+4AMXA/GFeAE5JPxC2+Ot
Hjqy6qvfkfEB5bmGKuK9OOw+5hk2+HYw+9y9yoJuaC1fcl6ZSVRYYOeV0AgyByYV
uyad7wz4jJk/BxAOKCNfHZMCq1va3lK0QRfLlZo2TlDwd/T5NyI8tjL7yQPEO6nr
8eCp1zq28ldOGxfwOtIirSgmTnhRU2ryE14N2mhP8K0GIdJjWqInpe9XhI6VZALy
TlhgM8yfMaQ9CnRE1Ku5BHqNeLmAgwpLPRCxBHv5PKdPf/9pcy6ql3H0MQ7lDtrp
XyFtCETvo8VKYntGNvMxlxDVUDDyKzvsk8IvjSNbQoYk8xZqbSjxuxfZLQExDV6z
OP66G3gXMmlUNYm24BQcT+LuTNleI6kRay8Zt0Trdl8vOaapy//f7zTXJNP8dIUW
KJrqDYyr9dwU/EB8a2oU6hgIq5fHo2igofHEdLrvMo31MLhkaXU2o3Lk8i0K0vB3
9IKTVBFCDO6pPURMEP3RQ7SKibmf0wjZ/dqktfvBGcCfzCLR2petM0tit95CMILw
IR4s9M73Jcpvzgxzy1NGaMQSVlA3g3OJOtNn+wiaS5rw6DDaWtGVfkIABkqxsfq7
MwJfgwighMcFQfs8I2jAUbjB8rYkaFldVj6Lyv5sk2w7/BS+rxCPfyddtwCIaxSG
HZZ8pof6bUkeAZt6rcczuc8cqH/Xm6e6UZRTpDcCE2thyrsXnFf2zxFxGpDqJkzF
PGOp0wf1fhXLVt5bYHloYKpbJfI6GWiO/00NG+weHAmd5KrdWFt0lrKN367/uKBp
OdgX6bFMiAnHsv7Dsri9kILxLIchwc1Yu0HtCbCmKM6mtKwNQRex5pB4cWuVxvYn
QbD8nvjdVaPPP0qEI9GasU5XscjeP36Ufkev8/+NFQc1DvrzKuZsva2sSOTun+qk
jM0Ou87dkfa9AWzmYPeiQD072PWsS1ijEr906x/zyRM/IXJUjKi4DRXc9ff8yuRA
82hYs4hGoHvI1DAaYNt1briMg92eQ7IN2cYiz5yX2Lp2FYHbU4YGrA/VEFq+3vRz
z1OKRaBQ3bQgHOuImdrkSjBJ5dY4WsJg4mFD82cJI453zuN8Wr+fcz31sdE0G1jf
K2+s4zrM5WltLBtAln/dzOqf9vQppJfDmiDk2FBbqhdBpTNHZbkke8bWzawIkiiq
4o1obDqqqgea5ISEghLeao6UxHz0VW17YfRISb4amIv4jjPv3ye15ocQI4BJr/rw
GC73MHtrqm5nOmQhlcYrInK/3TD1FNOexnb9+OTqrXy7jYBvjvRbzWSctrLoOPCK
g6FGl9jqGrwYinLV6bEWWUnGxs8a8Vu0XLZXH+gkXQuonqXQXg2eCLfveM+tboNO
7QGBHKXGHnXXQq8SkqykdM/LPtLnGzvTAbkGE2ApqOWmxVEIn5ukc7PjllTphzHI
JSCpcb9R0m14+QDccj93o0PbEeV6wTfICtlVR1BoTFfO174MoOCSQfVsL0FqYv/k
1eUZRxsCOv3yecc6zfFO9Z0q4/Qa7s4wq1HeSVOTXX00BCw66Do6rU+kLeAB7lVB
ASifWiKS7zYgxKeZ9gk9cJi0Jn1NbcN/qEUjWMtVtXJqGckzNgd1JHwnu+WhzK/C
BO7VjuQ/Royf3EgYa30LZ6HXq8fi4KqsI0ccmJ6rQ2PTiFqludQwVpAKQ+8P5Ure
I6PtiKMZOpvBwZkTXwK8IEEgu1gwPROjT07cOaI51R1D1w0UUhayxK5rcaH76gKc
+HT/5Tbp2iSgTNrQEGIq6jJcTWZCOO187L89lwfg74EOMDdeomV6Vfo6Iu1gbuod
0G5a4aYGYZJBxNvtF+1X1F6HL0lymcx++3cxad04sqPROFHSuiT+OBCqWiUR/umx
yjQPITA4sOC9wfpaTwZyHNhob8lKqaAdX+aF+SDSQinZy0nRlPtmh7uvnXrRJSsI
zFlEQrqs656xe4vWP3sS19ASc8eKYWkCxkEd513HxqkXU90bscqyTyuHrTWD1A3J
XwR1PJw1a5ydKYa8raCu6JrF/iSjEPSBoKQT4K5I+lESS62W7L3RcTdT3QsMb+wj
f+0bMb6sqEodf4G/2IYgTUhi5Ygz80T2irAKKPhBc8wHVLIVTVJLOiH0lQ6+Aqrm
zvugygOUF1ZkfC+Jq4TTRx7e4KlskOlOm4g9UmUyOXv4THtD93BfMcGNpV78eNl4
fP31RSQDHq/7iZ/9SS6qnuKbNclkKX4/wIFfdD6yleZX1Kw60hYmtNkWNyak7vSN
VPYvJY+/eEMGeZppOrl6WFOYm3JMIElQKA/w4yJ8zUPsw0Nm3WRYTI/Ht06uzYe1
AtZ0vtzDp/n32n/bwAHtTKu0BiRgNql1mO3Qo9TYK69HRaALzF0DKtX8ayPl4PZn
OmxuFzuLoC9MlZGJQNrzfVNPn5t6DvDHstAYEtWvUutO2/A8dw88Zb/wWqAiWr21
CMSwFwPXRxTCGcxXq547yjINUQbH8DvGj4vbIYgTk5DvVWBAJ5zAg/dc0Ok/IP6V
4kfg6gZPG9bK4DNZzwSMH5pr4gbguU6aGBX0WzHnEiMwKZROtrZqnYlnunxjdqJp
o909x3sYKXrysJ3oBOyjzxcVdiKpeaMRncBUNcToNwRg0uJGfl8IZ3e5eN/3YPSX
7QaPcBAGp0M/Afi51Y5gaEC7ARo2ZMeUFw5bzxmKC1loZVml4v8pw+PUiN66M9bx
joyj2Xy7rwDzmfnVsX24Kfo6S2VS7MrDtkrXrIyOQMZLM8Vkof5pxI9a4HUvhb5r
/OeZOL6trePR3ZzJcA250PlJL2JAWVg0pDi1G1gE0tcCVpfatUdQwI7fD+Fx7Re1
+HLEtrgcAku23cAbHFAfI2MAHAPghWrD/GJI7J8F4GlJcQqou99zneiPcO/e9c4o
stPJBzzBg1A30HGSAxGpGfgA1FkZk6ffRw8kg1rCgPU12jJgUSymVwpVuCm8VpTF
fSIB/Xm9W3uuacDd9tEYo1q530cOcS6W9oxhv7VniSE8AD0KsiD2FZr4BGnJCGMh
sG2D3q5CZ7/jM/0m5oWZnOkGr8Hdn4IYLS5kpjYOD8Tu6Cvb7O0rxPaSdiss0qcK
+Am0oqHxV/iN213j5OVQIT+sNcvu79DDzoi8lJc8Lmb+Fsf/cNUEMOCwQ6TnvKZK
voljcaFy3pFPaGTMfTNbdEs4uTbkm/AMNhMyZFbLeuRpzsS/XFr0Zt8llOYWVAGQ
wqEyYmbAfZHlgvMR6tXVmukWmpv8lUeZmxzZdNH9jCvIiZ4ULLkMpCCEsIo8DgQB
dg+tgvX/FAVegj+Nozdh7Yc6VlOm9JAR0+Yrz1AJhMkCiKex+PdBlg9F683nw4S+
6CZS6FXytWn/xher+ixsOHMEagGg5aJL1dM4noeAmpFCx5f7gOQfzzTvmdplBuRp
aOzVPD5Wgx8a/JVMUfokJddx4aprkTSxYq8YaVlwiIdpcdlatmhbHcZhsEKI7UQV
DA9GSMrCMCOTvktk4ID1Bxh5cO8SL3+yFwwHuxsCTR9btsfcHi7Zjqiuz6q+THDT
8SbpK718+RYNG8vJLa42/kza7LKCv2GlphM2iryYb378k39++Jhevu1RhRnYKF5r
ceojelisX1hY6+CgX3ZSqNe4tmLWhlzNqukIsb6lr1keqU0Qgeyf9O8qJZPPfNmS
jZ5gEOyRkLnLkPJ3Ju0W6PL0//kdAqUxBxO9AgaAtsHkFtov39zcbKcD5ZdIsH0i
ptA8JMiLU/ZW4+IJc67IcGqa0tkDWjugR2iRSAA4gXDeQ5TIn44CMKpshARgBtvB
iuxqngpcTf5HGUp9RzAGg5OMwB0gIgGI/TZpL3Hc0vcNgnPYhNBxPOOtxlhkWhBl
IYZn/X0wyGQ1gDx/M+T1mLPC+1tIbW6lSyOpxrupdrF/ORMyCG5J76dQJZxrwo6N
/75VJqM/KXHMVNwfj6nkIWSy9gUBZCtBQ19M2aqK2/anx7Ta7Qt8EozJmPVM80SI
1BeLb8HI9iomqZAAUCCf5q43sPhoxkLhbj0fP6lll3pLkxfZ8rzwm6DMa9K/WhXb
UQ5j8dzcewgC9ukMRB316A9ZnQgExUrSFFy/DxEBTROwJ53BkTmiBEYnZUNk2Baj
wwbgRLyPktEIw2I4O2r6VtwYlLyuNoUo9loKPEMROU+IOim6kH03Wbt92ETwnAfo
KcuXYay34lcyCnC+tnnvrS8f41G0iIw9vHFIE/o1WV7126pikfrXgIFcv84vXZQ2
H7RqtopLyy1BpfCd5eoxKiQjBPJ1zEAuZXnDSanQgKIMAFz09V03tQLx6CvBUx/J
rKq15KPJKUGS++gD62tmUQ1eHwJXP/vN2rsNELwFIfRygMAoRvJt3uCq9kyDKQbm
+LsnxdgFAsrUI3AX0+bsOra9rpsCvDp8RNnLyGraq7v4gES6/hHRGNR/U7CKp1a3
ik+ttnuRvs0Zgi7TKoofEIw85HDRHwV7tmV9PwJBe2UW4kKhu4Kveyh9WM+Xg1dg
UUAdL6xb5VxUeZfg31vRlT2BFK1NiW0iHeykaah4eG+vc1d6xEH7QW92IGA6gv+3
PalfRkaxrr0xrJa/k0f6XFovjNWTLWpYlZzyecDiNsqPdnft8e5dEfG1LAqmtJVi
2a3hZvzHXypShM7h8o0pdsd0TJZDbW7ANhoEzba5S3u+X8xT+OAbjWNM46UsXznK
BX6VCDjVD9RY+JLBjYXtqIHV6U9TyhLKWfDw8UNcP9Tt2c1iNov15A5nrV1av2oI
5W8srdaoRe0vNySLw46m207i3FxGyAapXdKwxu0A2+OsSBPjy8+03OlA8MHim6su
XWBgES6eOzQPGrL290nGubNrTgcuNrrZdECmCDkx10HmArihcllomezj6pPQ5C6g
aYvRFJiocUM4nRHoEyT+L3tfigTM37/qRzPe3/n5nDXFjfSX/casb4jqu0DzYpq6
C8ve9R5gL99c07h4N8vGSUw2/IOUsPkWmOTEvf2bhjdoNJF3Ukdhr9eCbre7mAYh
dSl3GsQr+gSn2hMchkzI5Vt3TUQlFY+/D45cwNhxulxZuKeL4IuhrFBgi80uNEa8
m8MMV5BE+/gtPZslT6Xae6dSJmjIBiSicnF4T82Xt+cCJLOSeE+VVrNRkRMK5tRZ
GtdtMC6F845lkGgpl1FBccJGyO+NbIP6pKzIQFv8tGfns3yqRt7OZLiTA9rgHy19
1l8pzN1gN0XZJH6Yo9jw6GDUcWjgTDKoK9ZeoOExV14dNC18HbtAAmCNYMwsrm48
XL1yT6uzpvT+2lTUzbAxGMpwtHF9r8it1bhfjBAwMPAxWCe+w2mG0yqpq+8nGa7a
igOIlIlnqIpHiF38ZozRhAkmWBdV8B9KBqZBdxsu0q+oZ0fALp+RP3zcpQNzFdZi
B+uEN9Rmytf60IkxXayUUEYPX8BcKTHMUZhDX77QxyQ/X6Fx94AIy5rHJeqSTGcr
KZ68cBW1i7d0jvGYBjygKggaz5I41osbkai6HMy5Wr7yK2Xjjc06Bjc4pdRWgUCS
4948zAMMHDPiiSp4/fIN9PSjHqWP1uMbnGublvnmPaBqKo6m6fFxZOtxdTYTCdPj
qer3S54xyQdRzytf3bpKb3ZWDqEEgPnF5pGtR3BXTJRc4A3UW7E4yYcWIqeUNWhv
A41vg1wfRw6ot3ZQ/vqiaSOHv0J6+yUtesrOrCBntbz+KB77/xTQmX/V5uzALv8J
OwKz06YemA4C8NTQkr/tFDUU1kmgDm4SWpvI1pFDlGX6qyLgB60qWqZ6qM1DFuEK
r3xaHGSArT7Np/mOpwo+ZoP8BxN8IA6GRKhoS9IbH2kFZzm2nmCnGYncMD9gRwEM
jpRPxp/eMIZ4k7eYJq1MMQvndY28bHhu6MtBE/nVuVox5ZQgH2H3Grrd0oEG/vHv
BUGIP/DFiVSXU25CeILvtF29L6xOOhTWZwQm0b+iqt1gyprtResJKqKhJazXFci5
ObvlZB3T340+66Gv1QDRVRokafP+IBv+vfFBaWJG9QzByMMpmq0YmtgVLNvTP4ul
J69+X+CF6OohQ7aixbEec0Nwk5AFrdyolI99Po/TNSUcpYZwsHxDNSOndqeorAm+
FaPduAjf4V4Zv+fc4uwNT8QgztDU5FaKR0Qf2uktKbqGxzIVBFSSw3xCloa9Ix2j
rZ+hhzjUyv/TFH0bqvZwp6ejBL9dHb24cBRxdiUqYMPF5lO02V+Am0Bw/v53mcqg
5B+Q6kogAJXAKtWOIu+w1XescC8SouuPIfnQthnNKY4AcURiEgnLSGTU2/4KygZo
hUZtS/0IDfd4WDGyLGnbVVC3oB0u3hKUOUdSohHnZKX4k3KJLSv2/0TWsN/QX+O8
pMosxVRQkRmg7mKiM8P+xYk8gmdMw1Dz47k9cHHlY/EYqz/P2/kbYpwZdhYmvVYR
oXQK8XwgWJR3PBmNS6n7Q765I5/rt3FpR2/L6FK1LACvddpmY/4dbuIKNVRnV4DF
jzpCXFAnEqujCQfv8RFVDztHqfcCunils1KUczSsW6fnxf7Lz+GgMbXnSTHscXxO
p0Nt9jhzHmyr9/NhqiUJLJmRM5eSi6voKu4f8wCEQAsFaqHC4dBnu3CJ3uNJQfa3
uzpX5L5QnYoUcT5LUVXFOotrehGcQ40BUlxxycyisKlJ+fY/0greJ0wjSDJisppy
FZdgJt7p0KPASWeepOd6oUb9UWP9hdglTs1i4Bxu5ydbXP75XQtYjIF4diIJ20rw
p4t3iV+hpkzE5JfoWbx9kV4GyAKUklZhC8TssvJKGJ+0gYKM/EfyzOf9giUwuclV
8HC0HXkwrPYbAutJufzFpaAaqOtL3bP7N1dkKmrPHVAfP+q+4josqjjPMfHJq/12
5z1OEfL9pU7BgbzioTSlx+5O0dtDYA0hzM+i7AHAh5p6InfIA6RoNWAxZe9sO5ir
4DBK3INb7qBbvzdOZrRsVItXOlxfrDinDqTkYiK/oUplDVBsTg1sw1PyPJo2e7d8
yBNXM2j17Nc9Vat5jNHWlBUVUNaDzZVsgIp21UGyTUDSLVJoCAUK93IjuFKGqjFe
qM4xVcpFZqP6FRtbeVW6DFasyK/+yVpJe2dfBHa+GD6G6r5D9UL+UV24vUyx0TuB
9LoDfzNu89XSYo/lFLwmH5hFVLgI2MXrM9bEH3njSfgt1CtLoxrtIb/PYvEwLho8
9Yyk73ctoGurrk95ZzgWYbDCGeAkY2VhLKDD2gZFO8Re7SkmfBouxXuFAJJIRGzq
i6kAlWqJyrtJupcZLa88SAYDSjawnUx5vpZKyH1uWwdxh2avok0ROvxVcHSuEX3J
qRcMp7RVQ+LoQb2etZSJ0QYdAO4cxyHSozhzcxw/xnhYJFDXpD/DRSehzKcl0OYy
fRMDJO0U3xzbTl8yO3iGRG0qf/UwkkdUPohRKOyQuMHy7N0StSAxHZafES3trJYX
vQLjiXpgXQFtefm693rIUlZ/HEtji4evN/xueuM/2M0PoEvJqCfk2j3wuBiYGkKL
yeBLIdS9P0oJ/r1iFjDAF7S2+kkLW5oAThMZ3H+J8Zxp4nnNK1toqdrU68Qd4Su4
UVb+0ANTOBK0nvBL5n+VAOBztTegmvSsAtgAXFyiJ9Rlhndm2NZIodR8a3MKYuJp
W3jJJhlcaa5fcGjalIMilqRB6oms3XkYUSAy76tR/VnI3YIZiTvSmqAa0J1pGZGU
GP5MYdffhlCERyn4yRh6R+WdqxemS6jCStP+47wWIC9j9sGo8/c7nbtFakpkM6mF
lm1/ddGwqJLGg5UDcOyVEMDyEIB6UjDib2nIM+EMCbHXr+oHkUHX5KdWL9mB+lQC
9quD1XG4Skv7lL1krT9CHd+0ne+DxEjlXA2nANaWutca0UYP1vm2Xl22dvMQGpF+
AJwJ7l1V9T995mszGE/qC1AbrB6bLeCm25MGyifDcDyZFLXJeVf20TD0gltalF9Y
4IDTZAEWNav5SVzZpfphfCEwIq1DzpO0k0Rf9OpUIBXkSy9bbEc7LdQYfiEycIfU
M8AJAvYhOyvWHJv2SClOecX5t25SUpWkVHc8bBeQbFP2eM9LDdyV2GbL21CtrdSO
wICZ4vK4lS8L4nACdLPDjKjFL2Ec+quGTBbGLkKyxwZXTaSItbZfGAkfzYD3A50y
ci7kx0Adf7Rg+MIXLxMjF32D69UEbK5t8O71Z3ldS1wYWVC7RDrgy5Lzv0fdQU2t
QKt2KGLq/EzAONbcCSirL61+O7wMyIYPR1UHlBa+QZFxzHaDH1fXE2ZIGssgpT7a
Z0Py8maU8TGVKKO+LDibYqY83gmyHf+7WqPhVcqulg8gvgLUe/rICErKEOZNnLpO
ycw94vQ94jQr9CfKyfyUdVOmouDvkhaCpeo+LALfPIjwf2rtcIlkxEeibKW1pozf
+MT4Yo1SHwymZ7XPEU40WRDKIF7q9P9JZh3YOPxEsa7RhJ69SyxGt/UXSTQSU0Jg
SZ/IUTaQlb6/O+7PXd8aXi2qXSNhPPKbLTRtFj6B27x0pVGEnYW5/tW84fF8CDuE
K/xTorV2sAebPI3PTVS8ubpKPetiVZTs2yoNXge3mJI9eowCfQDgJiaZG6cqXVV6
gtIgpn43hehw4wxlsH3n8+sRI4X7twbMj6mTtz1QoL6r+wbn6K2vj7jtYSmkhgK1
ROPTxcZWTv0NzUMdmr4EQbavweTrnAdTswfle/ITB06DW21U80UmiTXEyZU/oEdf
C7z25KhNXsiA94u8OLlh0YL7MJ6J+erQzjYp8kE0vs8wy7+ky6btd0vzwRpQ+xO2
a9d0b3J5MwN7e/5B21hPlLAEYV+x9te0KN9OPSYb+peYL9xtskA/CJJSbY68Ccam
hVxV3Hdc7cp5H3llp2ez5aGjyvzjgHMRpTdk4sixfLO6XYWS3kFmazYNx1og2wAj
JQMZUUKqTrVZ0/xAL8tCRFrAyUKgltf06ajRW5HuHo/lkNFq5zwxOTzTCqX9hdp+
QQhW5M6EcWHNRKmy7vKiLwpQiUDDBoOTJjp16NheHHboeZ9SQ/vjVgOykynbXYaT
Ja9uWWNk64Z+X8ttL9ujlZ+udZMINblR9vKYW03sfNJZK4lgHVJwGfsn1WgG+qz3
uGTHWccaBFkxAnEyAfP3X6ym5XYMRSEutChjtbipxjhIb9+5crvCJeUCOOJ7z2+v
aBBdrWF7Zn7kvAcourYiZk6NfzW3IB+UYjYicyCoqwijR5b66u17qiSJ1DhKFT8j
t3XCxNaJCUk4vlfizOZjGcIjBSNK1RY77cJvENwyid7TcxMGNULeTBipBjVkGWOh
HXBbbxeVZUSz7SYBocNkdrCD8OUJdKL5+6LgKg933UW2QxjSfXMoR8pCcuKrABi5
CvihUTa9XSHvBPJtqS6mAwL5kulPtYPFfKUwoqbs5aFjBKa99+t+D1/pDsQc71oc
t5EbWQuokFh09KDn0Chkf6xpFVhhcY4lEMwD8Q/k1Ckb8qxDqhdrZd4BH8onjfmf
6lncNVnpwBhq/07f+wauaEIejey5GDq8trIiDQTW47RVFLK6UMdveU0bcaz0S4uC
moi/9dTDz7iA+R+v5TjJ26fGixzHhswH4n+8PCqsvtmJueUceMkzAXKQl6GLSjZo
SSvAk1VND/GhI2D3uNCy1D6H5CLrOvDU3MohKBIdzrp+ZJSp1kzfS2tq7H9I6RB2
mdIEldo1XLE6WDoaYjk0lvCfdc4zr+f8/PZ/LXdSkeOih7xu5TlMa9GCjjFgQuuZ
/p1kTV2+oVMFB99ZPbJ2f5EAN/Y7W1SDynzrPzBVUIQBll34XLJs/oxNqo1JFJlf
IzBQfQFqA+pDCSigbbEKiNwmnARLjn4p1zcIYu2be/fhUwABUiKSI3gANthpm0zh
uFeRG+dX/sem9rTZTNXLjCjCZmaxBi6JTVQFkn7vuBZM60uc7Ps/7ZTR/5gY6Tin
lFUob8FT1tAOFMB1jhLSkoIB/rmXbXc9f09lLq2amkZ9YhnAgPIxzfPaAvk4b1qd
U2HjaHW6D7YwEjbLABLpXKm8fiLaQnarDix1nV6acZ6MHlPQKGtG0qvljnpxRoFr
QgcemkAW7gkdO00QtTXQ+iBYvvJcwOKV2VtMfAWhrAfxq7k8EJfYod1QJyTy0+BH
fNILSbxTRvylvducKeJqAlTsfmAf7vLtN1fH68Aftwa+2ZYtySYM46qTUhJ6iETM
AQDjO3qXD+hC6UCVgBcNCn+vLoNKmeiofccbKc4o0zMMDPXQpxuA8/yfxxqG2iRT
kEgfnmJMp34CsyjpRUgpCCKZXGRwAcLOGHnnNbBj2sPdLZdMqRYhUNuWmY/N3qSv
Hh17X1NRsnTMxUsY6NpzZmxahPWjgZbiReEgfNrspHc9kgIbR9adqostkMJ9YPFh
viYAC3lmvZKyf6Q6AhdDniKCEvzz9FxBdw+gkSSG3oLsIQi36TC8uL5hYwmSFPi2
hZ1ghNg5DiZc1nLtwnuzBmwmITVHQxSE2o/SDZgrM7TrdxhFcozBSM52ls0zhjMW
i93x8YXDpOa4i44hBt8vN2Y47lMaebmZKkDJpscVRNBuw1yZF1nXCOEcSle4rnok
9hbr2vSEWeFZ75ln3PFhq4hvYu6pOSvPQbqj3hf4/A0OdJt+D0qb8K849kGGs2dr
mFDNjJcypxfSK9do5PoHURqrHT8xhv0J+/4z2UjzBTnjqNRMr89rLvxahXoVJiR3
NstV8bAMixFh6iGG2tqgKZFg0UKDuuSVBe0aTqVe+CWgzYwJ04gknaFPn3OE5z0e
6PBq5youJl4hjQM5TpQD+hQCCoNl1IRqCz3I+ZRzxcbAdPdnssmmbJ+N3uYQhD70
nrLuV+wBdaYcaHK5smjjWZv/nGN9V+rznaQiAE5Um5lP9b1t4hOvAmq0EYip/Jv5
HjyGLIqo/QQ7IjuCBpqeENfgHGo3cLLK76ZiW0tWGPK6IxfAtzsPXXZhEyFnz+Nw
e5YuZ81KZrptXyIkd/EdSn7AgXKzBBdbC9pN5vmAMb6b5CvOjhqVfH7C822N3Bjt
GX/SNRH6DBmYIaS4jmVWJjH6geS5BEc3ea8GsVTP7B8ngWJD8w2NMyHuxEgH+lIl
BNkx7VsftOcKGspnxjJkHY+subgdJgKPXoE571zQ2pnIMA7pltdvDbbskAtxchOv
UnZYINC3VzhoaXO3yqXp4A6bTTBj2jP8ADFVXUC5KPqZg6giccVa5X6zXeUgDU0n
hpWNAAu50R7qVIPNhVgTpZZF09YcI9b2DDrFgnffdr6db3NJpkmxhlJltKt2tRL+
Ad95wxy5yLOoQ8+QDaDD8CClGpmil8I8+2Z/pfXyI9p2BsZRs1jF5/GrD4gVYoOX
G+Vw6ptLkLfUISqArxaVwrbJOe+dNQ9YJC+V2LP79om6LjDJuYaMdppz4mLcNqHr
FYVU4lfTSOR7c3K6bgtMw8VhSXnhWAgkrUfBry9mxb0T78o7WLYrKL0wFuH8qWvX
wkvwhv4v1FTXDJ5o9VUN7gjCUafZDPKE5W0+dCI0AGFzmtPXFgQqEH7Ee8cCswjl
wQO/JoRK4Xr0hFmWbpHWllXBO2/ERhdSUK3ndQVIkeaIBuG3MQ6w0XsbBfQ0PfwV
yTGtSppTaHVRr/8R4Rr5/1z/25fC82IcIa/eTlqlypfuOyR1LiKsf7oCtQJBbdrj
6+L6nFNHxULwV7S5qNota3b7bvT1QefFyX9eVpbBC7HjjPO9cXw5yPXNVB88R0hW
OhFLToJXZRzvlqmJm4OQA9Q5UuVglBP0R1YlOZkccX1Qrb9Tyxh0Z5OscG4qye8F
xfTnFjooqpz/l1/k5QZGBTuK/ab5/6cbiUQdgxEIGGBUtpgQRsQp9upiuDrq7XOS
SzbUGz2sMbPg9cVcp95ax/uLEojR1/b8f3QJU7asIqSBpDyJx3zx2XMMu7n7SX3K
0g9Jfv5oX9ufbIn6R6hZryYB1JsO7+lHazw2PQA9fpohWo7UwgjF0rRs54Cic3bh
q1PsyhhkAgQoRiHg+TaBllelx3rK/lh+Dq5UFBNx79jvu5GCAZEXoxIBo3/SVa/7
HS3wNsdStd9Z+QgYNKjggdFaMnsLCSxdHPnAsWw1adqkrMxPoue/tZl6O1dPtFDB
N76iGVoDzwr5uFEp5W/KZgIYkGrbqhbMOrkAZ6vvJeJoyXiDrrFr64m80+/55oaj
fOenTOCaK4wU6U/rWtajP33mx2QWuqx2siCxCYjdvUQIk/XG+q7X6ICBWGjr+4Cq
prk0xRxPHRtAbsCnn8L65tm+454C32goRykc1A4ZBbiFgZXxWdKRr5RTmhhhyjAr
yjNNKeTR3XEWBh1qmzBMJpPwqFYpBjAsnBtCrnYFj3kvmcEryDY1qBWDWgIg7N7k
sfmtkF1h0H/eAJ3BdJ1+pbjatK40suFE3UY4lIRFwszD8GD8pawOCaKtSAA5pQTp
sTuLg/Mk7JxFJuBYIU/PT5O9Mt441EIMG5m/h/cSpOZNTtqtyDQYa3IUXDW1Q4ig
wETwr9an96kGubGu1mz7xW3IW6Wimwg4KzikVh3BpItkyLDloVieXNOeZXMcO9QY
qJOkcAUD+LV7zIQPBQe3Vw18tarDoChhgK2huiY/vT4ul9BWxq1M/KGWnmiUBHj9
oQIlQY9iUfjmlT6mjg50bJZHB2CCzhlstkd8LLC1mKJkMtIOSMGNSfLAax41noVK
0VctmLQ1zH56j0Kc1gitGmzuftHoMpcdgPEBo+jXWWiZmHnsqsSTO3cszwGoPXD0
sQszljcVUDfifgD+2gda3JLe85MR5DyjVsOSuQwUnTCy0khi1McArBz7RlKm2MoG
9Efmh/cSDQ6i39LXg7nzsOL8TnvDpMnY4+JH5tBdA9lCuRAXzDHm7ReMjvqReChP
kvVdJ9o/xA6q70DAuk+MaPdNTcXRGvx9FP7XJf3KNu7nScykQSv1WGwGKAUJDO4c
HuTVHAsS21+b+Tfu0P18/G4fe32uKi3SbZo7G1a+lofn3qkWlEsDGgbXDOnCy/PO
AtD2krvr7MKAbeKWyIM2omh+1FDDtFWHZXun/PZinC0RXCS5Nzz1OAbnkApEw6Ha
0sudIbRapNXuW9fUWWqFoIQUpEm45QzIgvhJkD+Q88G5HZeFiNp71DPGxjPY/R+j
NhWz9T7NiXUobIJ/NbT9ed6CbVlN0aoTviQ7ucCAbaIXTFYTCOLVxAH8ZR+LbqD/
uWult2gb+j6aoH5i50gGNunu5xy4ZRRI57YdahwB1/J23NLmEtfU1hewbKVqugHn
dh2sCFNVetX+5S6IfY0iDgD63iTLVjmi2o+yc+Rpi1s5DAudJIqeomjSf4ePTIMr
g71g3cp/RWDOL0tJm0MV2yIJq+dg8Vli1gkfEQn8AjPpKDZsey1iZJGjI69Bp3ag
r9fcgnBk67b2IPQCPJUs7dGs7lERBHYN6gTDTVQq6yAYf8qlHzxMAYJJ/QaBLvOO
k8dhOuxcdLNFBIKHH29f5gDhXYTV/d7dl7z8tccQToAzJa+YtPgmRpPMuy7qnvIy
ovpqMcm8mQmpmH5aN6mxtDidQ3iLBrToAYoDXmyRqSJX/Vby3RLB7bbJgm2Q1wTh
X3ycVwl+eLEaOar/bhu8N7yWyVLZBy7+FTGywVsbqlHOwYQ5NcZAi89xOfysb1ug
AFiCZ4bpc4svCnw6AZcMoDJQCuNp1NEHlp4Q4qOdI2XufyZTLkt1q6t5VwZo2eVr
a31lILCQtlPDj6GZyWzi7/IAVjpfK8ukxGgg+kBn4NV1uNeHaqWd9o/GBc43hw1l
IsrfJl4R53rurjcCd8y3x3LM+JP2vo9TZoxnru39fYBCWlUTng1NK9NozrN6VD8S
4NRAI05S+PP+GHxOsWDFgverjBadl2o+9h4rllHF2YFCqSQxHeOHSBqlVJuJc/DE
+X9/FVHT6w+iHmNLxpHSXvCRVhKZ3yXJwei8rmJEoxxnI3gwnVzVAPZIgll1tn00
KFggtqGlEs0NKgc2QV9MbYlhBAMntVjJq0F/3/GaGhJYg1aa0VMvXwhu8gfeTAwp
y2ca+Ry2CtxzvxmyC4QnB4T0UxLfjDfzzBtaAY3RQKOtf19KwR2maDQ2PlC6Q4IL
gq4kAJaCiz6E4AonSMVczBhC3XuRw39cVXPvFFBmiUnMcR9tuaPhPHAc2/2EpX3Y
Xo6BPTmx/+drB2dhHVYSKQlCpyw/v/c562P/eWBCF/9qvaFjFXZfJJt+QcVcKAQJ
L5vAjRP5J2B2UOTP/uSc16FPQW4Q44vqRvtdCPdK9S9QX9OdgaWmvoR6iyEmfrJl
7EUmWZLJuZdAZopycU1xL+1VkTv7StZz5WgMXzZpzU7oFsYRgA6GcBazvmLlXSef
y1hxVkw8W2qw3+Oze/RnVVESZNZ4ru3lOcmuv/vABWz1OBapkVBIJ+yxpXfMlkY8
Yz0UatKI8MzVlCE79eL/N5k9PGxEM9qrP5htgdckGGaE/Ba7Q1goP/k7/FPFTCkL
heJMbA1BwUznQUgHp0TATaCUYckTmoCmFOSVJLKS//AE/bjX2/4yO/M7Hofo2AJK
ru82GCrwKk63Uxj3uC+w5PYhkOAwlCAVz8Fg/fgDHow3UTm7pJFIDijzvxarON+M
uM0ueZ/u3ADznxJ4R/pfzHYHHakjh830YDT//IP+vnMVex3ObK9EJ93yfpdMHhuQ
Mkq/3VkfHqPFBklid59P+Cfkn7W45LH0UrML3ooEHPNg5yQCvArlgZZLp+cKR0j9
nVs6+wWdI3pLxFKMBXpmTHkF6CAhIeKZewFOO4MWyc97FcXKkn8rDu2wQSLhxDr0
kjtUeVhllG7sT5qDjd0mcZdKBv8FdfdDf6UIKA7KqkoJYUuDHl144sILUkeMASVP
1P46Ojh6P8LnQ9FePzqcWoZd37QV2Ikius0P9hriwoQdkluI/qDs/7luR+BniHJS
qv2Mju4LvwGdp/NlH6KILu6lFXmf6PkODl8eM12Unvv+4+yU1/itPrBGBRZk6c5V
OKn1EY4/OcoRgkR+8FcNxDK3nrF5yHKBBgC9OXaNqurB+WnD/XwponmHRwRSZ+/C
G1pzbMz49w3/8CXIYHPbIFzoPb4vgwZQH8O3/ojAg7vNO+BOBCLTmco6+0A5DEV0
k7a8AlwWWiAbEFvj+KPZVciuHfUpICtXk5iEnYgzi01EsYQm/aykWO5SV5yTZcG7
AP1FUxvdP0dFiBJ0tMg6Yo/P9jfL3EirXtvLp2fnAPmUBbOxaeebo9GqS1/TvAXe
YArS65FONt9VDaU5zSg5dNtadYwUTJAcR3p6Q84xnFFWmY1Q5ON2eJinhAme7vOc
Ito4Q4qGORWYAGLWY5Unb1PdXxYmS+31fMNhyXXGu1INXnK3GWrf+uKFMD/PhSe5
D0SyI42B7YLQgjl2wHkeHwck0JhP2f1fCCXMQI2ANboYW6aIrvhYAxWw36dinpCB
vo7soOiLUKLRkGsaqV78UFzWnih04LNjbrAZtj28j3C1k7iTvwZRQpQ3o7dtKZ2a
eDhWpNwttXSFS1pEMK6JEStGJi8S6Ccc+G6DgCgP6rW/jk29YS8Sbqir6FixKsBp
kBvhn3HVjIBY6KYWHF6C+t8nNbzxLpeCutRsEGu82KIIByOjtjxTn8xPBnXTLbfV
FYRbgd+mgK+qCLP8eYtCyLJL6DfkN6OLA19a+X77qiitz09XS/bkxjAbGB1VKdgm
X01IhO/6y4pF9glKuVzMeaQ+RgJq8daeMO+42OVi/XWiElxRnHZomG7143xMrpAI
Ro0DN4l8YHnqitS7AD0PU5K3MpOQ3Mee/GnGNAwotu+8dgTQ9TdplsNiai5RVrze
gezyh2Aq6MLhclnVVSNsXkUmvty/cFZOOEyUaAKUvXmt/YMfvmB272AYpImAZRV/
2bFHlq0s9Q1Qn+0XH3lKj3uCWrQ/G/MTFXSF9ylDG03mNMtNw5qk6LBOQP/jk24l
/gIKzUh8nsnFd/CNfwiSmarhVy/TEX7LaBqQakdcMO2MDhSBem34HnbD/42uGpv4
pokxK55fHbh3woVIceh0m1rtFiQh9oMNbmKYYvHi+pj7bIKgMk0+bClVNPB5e2Xq
rSeM6DUA6kT38aExSIbY5aD/KQNHAL/3Xs0pMVAnkTv6EFuB2hnGds3s3jH/vPON
VaHS9H+yyNPlh6Kk2RBNY/l6Zi5XAM05qtbhXT5PAKveXbtPuxiwcDnwz62WzMzD
pZBfjIsPgOrWvzSO9Xa2On5i8L3hp/01g5gqEum2o9Dle2Xuu2Dv2CGbt4eEIiHW
lCH3oavsK6nqwsxiQvfpPNU7gU04Lmylz+EXujH2NWHEKBsnKcqXGRkeO1y2yrIz
t4BfcI67SPmw2HYpMTRXRjJ5jMH0RYUCT47oOEvPUOO5JcuLsYgcyn8+cuc//zcD
ibzQ/L+FjXyxitncebaE6q8mLDZ2bukBvWcK6aqKlB/qB1BNAAj45oG2v3fe8hmR
8yY0vi2OCb4wgsi/2KsUBSHArMKtKumG7Lm2e0AeZ8Pqvnx+7kFb73LKmHUWT5mF
TXGXugnSkZ1SeT1ZOz2lLlihs2CAb9VshwPx2bLZ2J024jvEi4NH7G05npWn5sYv
BA0mM2dg2NuQ2OonkiJIcSdFZR983PBD0aHVQKn1BsbCOvVJpEpndzD+2RDcK8Nk
WKGJYFvihc/E6UbtcKuzfJFgmBOyhmAuC1sikjd7lkzwZvto3QRJ7KWs6g0v2vnJ
94RuGcjnYCy5ZsKDMucY6cUKWMFqQGD32AtGDliZXPHJjrr+tcvpEbglZYLxLFF2
7GVaqIq+pgwlCwwRf/v1xiUostw3KjeAKkCeaefqETQlRrhBSXkEV7KDdurl5TuI
RH916qAONsE6pUJF79gx7k5phe1eKw0sXS1/SnBbjRyjNgkOGXG3YcIwHadI4zot
Z0k3KLxEkuTlkcGwkDDVTCN9RUPQa5mYGCL1wFEgb7J5IuSs7ZMcpWbbjh6eIZi/
1SWBAyjS1jdqM+imRq5zZqeEEGLB5z2vlXSTGEFaTycvm6qL6M0fVD3extB66NVz
bb959z5yly9DYrDmDJ3ml75A2lpYYUD86T1+HG4PbOzZL4zhA1t82ZP4GrMWaayf
RXYHM0JED8wGv8Ud++kkKPVPJD5WyO5dl+3ImZd3pksjmNETfunjTq3G9na4kBh6
2/3M1L6wZt7JPRngWN0eFo8XTSjtVe2vBe55j5ACWMbHgYrzYC4+PvWHUfL99ipY
3ZoowDPGXZbdHYgzQwJlmUWfpukivcWMcMe0/Xf1/gik5imyPNQAiGQdpdOv1/I9
o65+L5HnmrbwfpyD75Du+0+RFbqMEstR6eTefCOvp7CBgoJrVDrXSwJmqLn8wrxa
no1q4oSf4S+lVnIcGNUNPBuS9FGzKYHxoT79+VlN1l9+fQAULILAJtz2fKx2b3Y5
uoRs+cpqK6asjquz4rSijp9ETTH84Y+U376C5pNQ1S1gjtTphzyRTRygzPIbFdMI
pxeWtd2PbPPHp5AL5uNEIK58/5Yco4k/aoW+uGnpXOeUEDtvFHq9J5MZOVdgjzWy
rLgycFBYqd9bjdkxga9UUa+jwTtz5ZPJZmMcXNeqKe0u7CoHU3fbVAa5eoVb+erH
0c5k2hynPUfwpGEPgqc/PBvLAuoQ3k1pMgrzEf2gZciEaHsKWkxoKqevZk4+hjaX
yAxPfYxxUua9EQWMuR1iouxqHbjhNce5IZ6y8lK+TU420ZzU8OJpzHPB48+E1IP6
mjKdB/QtaIOmeqKEG8/23EjNamN+OMElNAPpczIxRtTvQmTE3GR85YTgRVdzyUuc
F0R4mv1CDDUqPLCV1XGlTEKwIIhWHKKfN/YhHZt6+DIliIW5XVqcXSPAg+T5Pimh
GPMytwAqugxmGwqbp19EO2GIR2Zi/NhYE1hS4tpIAclgTCaxrkxaWFjOPv2PJEsn
L8m3lcuC3sczz8KUJxa8/UNjDFRELjmwMa/renvAwc8xCjFV/dC6k4nxGIjGV9P6
+n9XPVZ5o1dOwTBqETFEuhPhDKPvsEAddEypcD7Nf5fpzChuqqgrEGJRr/i5SdA8
6kXPNTr4Fj+oq1TtHELH4r0y6m9ClylVhR8x6By5aIp3qRzSqbSobZ23Fr9zouSo
CfAjX/cNSXiasZxhhEav69Anao7ZB7HEcBIDdCFm8cfq6tcIQQdA+XyGspfM58Nl
w8orNDhNH0B9m7ETEbxcMLytS1aFzkcu64Iue3ourLFOA5QVWnuR8VfTVsLIV7YB
Q7gsvfosGXD3yylBNgkwNaw8D1MY8sCxQsELV9Kd2vwpj3rRmn+h/Qd9pQhsZtjn
DyIW/gjMl8gRzikc7eaj8S/YA1RD9iQxexw5I4wtnWK/tXjbkFn6NcZppsswQ91i
v5soMhOb9hpeyCDUd2mH+kVdbkSFuvRTI6jCrwC+x2ntGl/n7flmXxFXWCNi8+nZ
Orsp9H9XCimt2qvvGAlPtsbJNGPIvpj6Y9dQ4IXFNJbv620WP3cNr/HLqNNF+d0c
UJFwJehG0EfRg5NyVAzKJny5MfCP5O7gtk73I4Esl2NxuVF7aU7/uxQ+EaCUInTG
8b1w5AE++KDuleYwJl4P3aLwgbGvMsvxErIllBeXTL/NC2kCX6k8GWFEDeOLPdiO
9K2dluIuYWqmBARTLaxqcdKdZ1gnbHjJDEXWF0kPUkuX4EhNyEbt6xqmT5nC67Pd
J+IC+PgLEgqMOfZzs0KXTEqGWqlfRdKRjWHXewgwWxidMSO4nfQIfV9FzL8Vk3F9
/GJeiiyDVoT0MfO1RoiUUXYeUJ3HiEKs0MMZPVZuqVr0nMX77xjwl58dSVngG8Aj
zCjmlOn/OX7LWlAd5v4fjgg+hfcsCfLmoNyhOs13/cmt+eDWtumG6oR2CErYpmKF
nNJBR/6MpZAGVr8vwnRD0m3WucDzaum+a9aAs5Q9BUPAxukRr51GAo5iougdjS8M
tmMr6Fi9Z0EV8m3npOpaZQbJbsBelta6kFPQv1g/Z4AXPm0EPO31RkNZaXZ6ttG5
M3ldLtkvJVS3TuTTFMXAtuh4oK9SlTIToJO2aJms2aAQSwpeyAerryCpdMU9T652
bntx092XYIZPb8XNkRzR3cESMXQ8w7nzZnKY8vnRQnYXIQZjOEBKSwNM0Yu55dbo
lkY7qtvRkOQo1E3meICSbv04fNSdp1bDQpV9RFAhtY2pvdL5YBN7P6ppHB8mz10F
E4izBBRD7MPcctdoVjyNfZgKopow5AJ2EfyhKp+SijNDnnwuC+vi5hHC7qMcs0J+
t2rqXnjHvIvA/GAHcEu98fyI/NDkQRv7sQtrwLsE9P4sdqi56iB486KYZyGT2WKa
tGGLBwKUwxp6UuNJwA77aSxkvlyd2Z/JrO6rFPG5NafYO1bC7uIM9BJX2vNpjIej
WXprxTav1abaUaWw5qgBirj9gz/bhcEY5yZ1ZFm0pa55DkhRLvL81DqvXtJYPuHt
xuem91kAROOQFLrMDgVCiNvkk1RIODidaRAlii5KAJWwp6DKeQR5PZTFJmAtkCz6
kUld1xv1MBiTniPlwk8tbjOHx6ZWSDUA+if7vtwbDP/CDZnY3cxzJW71lnTJ9n5i
SwEay9OkFdcqhEFCliV5O/SjyRIMss5mjrAkaz1irlsAD7IUOhKpPxfuEmo99dxo
SF5mhxC5ggR1xG4ajUqEY5cMZkmdwVSIo08CUxpclst5Mqwa2zoXdPa854i8YlVh
lgsSoLdpC8BEHkmDKln/zW2QVXX3f3T8otDNjcipOyZt9+YuZQTRW4M8pFo9lzVT
HjUGQmMWnoaaYoqm3/pjnqeV0HrVqVUTbkP74qQvdrdShbZTKZc+BhH5/wZkKNWu
KlVtbJ1KGxUvjMhMtzhN+PFwd5I+NI/Y3R8YDwQ9uV374Thf7K5KCZtmX6UTa5bS
Pn3RdAZRaQSI/g3tFxeZzWJNkGGeY/9uHj7j5wqukF2VPjbCLuRPHVUs1iXWgASZ
+2fRdHDuM84IKqswIkj3w4BizKBjRqzwfNwsv6BSopJ5fJx9ZvVitk0/eUbRz/Da
nqLuIqhr4CftuNmbcHRilPbeTzSI+PMEKeeJ5GLc0FGgcZDTIGOY9Oyww8YLeypy
VVkmSia048kKvsmKeLSNbKAsk5jtDy4UOV3xVvvA/UJiXOawd223QnvmErueOfWI
GtzPae3/Rngmvd5byVVeooQelgm7+/3Y/pzCcwyDusE4jqT3U+h1gt2i7Odj9Iiy
v3mJQT4y3EZioOmFNygVjhwt76PVabOptFX6P7Ah/vJGQ+dVNUSw+3zz6uYqWDkb
jfpHOOd7cvSR+mwqqvWbNAdewc3Vink/wESrB5hDrpK4dt0fRoiIxb7c8CfoYSus
MtKkuCMc4ViwsF49KsMTAEYgzHmh6KIfPgpKqs1oTb7hrzLUBArm5848NOtzfyE/
f13/soNZscVlJH0ywNMuX4qL73nfylBiPoio1mMEE+S6UtQ0snrTnZRPjbxlVf2F
3YOjmA1DCRdO/V+ny1oE26r6PxEE6DlojieyHsu3IhaVhZIRJAfVnwGkmfkradgn
IaNKTjcYl9cNxc6KeQTntjg5vvQ0El7WwIvLPyVQop3stG8of/8MmQenRnmhChuj
WkdswbWd+Sp0ItI99Pb54TMTxM1qrQRzW5yjZ99HwTgzQozJUBSSbviw06R3E3fE
J+Iu4dsfrMK5WwSV3erwUAYkajl3f1D/o4g7UH5msFoMhtqmqgO4fpEUCMifmnDF
L9OxEJZXpslTYH8DSa8Rv73d50AcnqfkdxH79uqkQBYFLlXrfKAp2crFOmpFNYhS
XtmTHS5xrFKELYhRYHVyUtn2zQuQD/swM4c8aeBdkietLixMJsMFKP46Y0kD1w/R
qsWer0NwPc7tc/ctTUwugroBxCOq69WRzvFhLc9BOjkPCYUpcPe5YD7dUNwQryBB
6p2laj5ql9lQqWY/6E/3zwRR10kssEWWRLeBRb6KFd3ZlR+bAi0ojzL79bK2ROgS
azmg9Hez8i4CzQ/No9HxJCyIzzsk0k0WApoeQaHXLI4SFVV80TFGzy121lTJoNS3
fhtICY/xQwUT29vMP4OaHxc7QD9tDLMfp6sev+3/mh7RxbAig8DvKnrGpNUSV12n
YQL4w5a6HCbbxJhJCurFaxbyGIL6KycQmvedhfL3nZx0t/vtOcxMXzxgM+yuSU+B
1RrhwPOv/0I+SgbPaZkC61kBfv8WQ6MVw821fGY9uny2iD2YhOwcLbee7XpOH7it
Urh1ko+z27n+sXuVUfJRqsuHAy0VhhYRz/6KePxtJyUxONbblCqGUDOcVpVfDiqx
tsku/2PsE4SG2++5aGy0RFNexZWQ4RpdcPaJYcD7Cvi0VPfZ5dK6MTNpil6C+6pP
50P3SV1l+lcW2O53FChjApbtaMZfN1jEgUC7vYaMPIHlRsbz97HlQwiFYc1GDJgZ
yCoANsUtn6wLUdqogMy8d205N/+fbW0k0TYl+t+1GBzmki2fkDHdYD6guT4i0zLA
ENLPlwSMnmYEhrd6fGjjgkRYGaUOnbjUvyqA7FK0Bz6BFaZpg87uPi14+SxcLSAF
e0zRqRkxXJSdMKOVGjd0vUroMu7tPmepq+acz5NvfafBIm+lSvmJJECSy81/ORns
IPdgtVoOcqS/rcQod565AeL6CobhJAVD4Z4F2s5Mv7dkie8R1wl8lY9zKvPQ2nBD
yASdKMHR8M0ycGKd4Fl6zjGMT3aV4+4rh4n0eRHltpAVCHPY8S1XA5W8w6AwqIJk
gaG73PP2HNd3oYS5VxR+F+5qA++7wHss8cevnuMkwkhVJxN971s6q/6tJGuFnw4G
yWurWr4HLQlHq9NrTlEWiQ/AVR8Va4VQjsoPebzobolXBSiDqGuUtR/a1FXBgm+b
O8Yg7z552AJRmXrY3TqQVft9SwHNunRTRncAzWgQADXphV34Ys3CViE6PYbwDKwB
86+0dSQDr1bcdHwvwNfkVpUXxaV4aJsX4Lp/ylNMpE5S4a9bjUAZQHvpt8H7YDnX
zejVzvPCqNKzp1PwuQjH+jFFbVyQCuePwigg4pnv6dG2rgDLw0I02nPYS7RBXt7l
li0Sv8VyEiDLNWPwx9TkXGx/k1BHOnsrN2EnJ8qsyZwPaORKgdjmfB5whNHIDyDj
qAwjQMBISEez16JuTfMDB4/izZ6qaOY99MWKmfz5JmDIkL+mew+8iJgUTkSsalsR
G6G1ZOvrpfzdm9yYAxcKA12l2CcaoaCHKPcqWgC2iIbRl/kPPJgTbff81dUpdd1w
6JKqJKMtRiDLD0+vtN63FuVgcFwgZjKbxFyEW4PSYBihcYO0k+1h/kFYcKP5Mv29
Gdb5WXEbQnqJZ/JvGda6nswateAAgL4FoI+ynfMYe1yX+6zpSzmFPvu4ykUDdLHA
mpzNGcut4L7JcdwIUWO5Jvf827P+F9zdw/LufPd6z2zwJ6/42eYgyvNj4BcAUvrx
LoMmS/017MzeMbHZoRe7vLpQHX2qJIEMOFFZ9FGP+lkBvTZTaNV+ETZYTB5pmBFG
f1GOXIbZ/TRfUMdjn9Dd7jIfNQeDTa28V0oJtrnaCiOQjyhM4R4cqW9dVwYICwyI
Pzh0g7eFY19JJ6IsqH4BM+Jycywy4+CJ5nwFAkzCvPYgbaeBnvyXztwy/0f7uGdh
q/1B2rsuam4CDomgTN5aFqwRtr7eZl0iQqQR7YsmCew52Zn4SDsTQjumbHX07hwF
bsKPUzCQXF2XLIA0ATcbIbU1ILTiHEn0bh1tz3SchCa+9J4NLso5IKqcQb3pO1XS
U4EMZBLrA4jmWnZAVx7rCM0dKXFUbh+5yjZyNS+xWlhyLPOAM7r34onq+579Nodf
uJ0JzvrrMLs6rQ7tdUl19uAtO3st018uUKVi1SSRWca3RA5LlEhyg8lRt4/3l718
pQO13CvMm+ku0ukHD0l03V1TYctuOXwQwI/aV+SCSuBgUoAo9F+Bugn3PlvH209H
QZxreeAtphShx7hRH24nzy8rNJ0THlqrBt3z5HgM8p3TvmQ/Ju3hjyA68niQT9Ht
Msya6Zus1iV5JU2mlxnHBZGFxDSi7gyEybV8iPHF98g9FEy77WDvwUlNP+gb7edQ
5RPS1rkm868Mux8FMJmkYf8pEfgm+nhlgYPbbEU8dT6NFmaNqf0duDxayORA5la+
ngLo2ibagDygTtOA/+/n1BXFzDHxPUDOim5+98LmtMDqPDK/UtQUEGj4aPnks1v0
KDqBKQMsFEBDaOB8US5xhpeapesJmpSIvVPq6zVE+Rc79eAPnoQ+w3oTBh6Z9+sg
iM0WVgDH9AV5svKALPe8D6c0zlfOrkIdAqKjrIcPvmlEwtAOtGojWkHpCsIKRsMS
CnjndTw5NtxsJFAy8wkrGBvtCo4KDGnxZgBS22cmLOt/+doGNESNTUVrncMdSPpr
jNukJ3ewpdBL1j/3JarBxBMMYi0ejDUEm/AazHy9qUThZTbT2FosAz1rKCl1flYJ
/xYGy+5dtDMVfSlY/U56DUkmYU+CuUFGpLvrkB4aCHXnjKKiKTKBz9b+t5CU3h8X
ouFzqeq4ye93iUGDYduEWZsQMAWToIsvrpRnl8rY7/CUqX3Qtp1FTTJXkMEJ/6gR
sRkk/+mogXFRebpZ5O/uUdIx6+CXbseEh7ibvvQizdqdCBQnaN7N071yax0MhFoe
VxF7+9hVslg2QhCq/33qVpZ3W9J26n5VdhgYUfMjJHyjlC5EvCceZPYvWTLAK/+E
rpcjHRqzF1ADGv9xASKhMqQRvKdVZqVQxb+JjeRMk2x7gR6Zs6e09snylZNhfDXb
G8XjkpxQTMAoeEQMIosmsdfAb5jruO+QpA1MiLhk+H9MnzClW+5OTeJRIouWn3DP
9/MRrDPkQvMMJNV/5gAvlRXGJHicBltdFrO21A9QOR9cY5obQoZE2Qmgd/6wZuVA
igYZXelQfJeZ6NwNj7xivVCh48cPUs7+RtGZsMrgXAno7aw9mGXhyqQ+nqvxd0lR
NJTLw4meR8kcKenyxrD6syu4VYAS4R5Se7nULObMZEdiY0ILaS+BstYIvgW3T8Xb
YoZbNM0lbsyvQJij8qWR1GbDRJrzdX1LM6sX7vY9lDkpkEkIoVd5uZIWQOxR+RlV
V6p299YZL4Y4rAFWmyrMJLzPD4W/1RWdr3c/gMvqKFoOZulwYYTB+hBBwMWC5JcK
Ir3LU75towWPG214WGt06wF8xe2KNUBWBev9L5RRwI99VnoVNR249PoeQu/u0g8v
yI0REP+8+t08Vc7gJozNyHk1ck2LvQtr50yMP/vRsFOM7f0G0otLuqhqe5quE9U6
KqbN1kdKMoQNRwC5CKlg/G+71QDUlTT2CI56zvswX5ebKUYFu5RtjwilcpRxD/h7
v9+mgvL67xXWEuM6kS6y85H9DFohpoJUxFtuQazR4CiQ6lm/ysMKUadvJoDRg/jF
d282aasFihl1SxwQANwGlfnH7FuXAQlCfg1Tw0FknSBLC6Agiprar5kySw6wOXTn
fY/7E+26QtHhDV6YL0j/NNbeSstcI6EkdP0vvvOqV5dSs6V9kcrWwrR+E4JTupQh
PFugcc6J4m5ZsyX78/HA2qMH56tiu/UM/9JbxTj5RZnSRUqa3+gAh+xmaCx1utWh
efZkqSCAHjPXsvAENKTWEu35gOHmEg2F6F+BlotAAYe2eW+/MMyGZiQQYJ2SbBSx
04n4JgSN9fG6h/VJDXJMYVuhz39OM0uwVPYyOhvuRbYI+LuxtFViMBASNbGP/qb6
VCY46K6LLZvvZZ2bBtvvhZxapWde74x0CDjh1LCoZ9LwHV6V7zA/NxlZe4u+z5Md
83+aNv9odVZWvi+Yv6c6HTaThbC6bvi9uYBTwP5UFCxxzkkiHG5x+u/AbTFVBNi1
PuVqtSVTAA6o7Ve/Kl/ntwzkDqmpzuODksI2vKmN6lauvGVqM0uIUM1FEkYy5X/v
Z9QtucUr9x7FqKvUDk3wNA4PJCDTa6HXwQee1TTl/swXYzfcFLZqso+qjMiRYTe1
lHMrZbFwS/L0idDLNMIjkrPDHqv8C1bIn/2TngaEos/CNpSKTqwWqz2qEnEXZIGW
T19f7n9Sasd5LIopSzYYyTvBrZTUXqkLpyR/G8bsI2W3GKREAx+7cz+qcAPIMinz
2Bbjp7JIAhz9hGdRXb5+UJDkqL4jfFfEacXlC9ayGCcw3SsdUwCzxUgDqeEbOXyP
x9fhKeyrNTDNT+G1rPgiC2WkTmYKrKqbCwvo5RH/FM7dwcomihFbLgktH1PMs4Ep
JLdbUdoTd5coQNxkthgnS8gys53/qUdmKZ3ZV50KGFYuYIVMZPLEixJJsq+QQrYR
uFSw6K77mF7BPayqSyeD5gu/Zcif9VUgkJ3A+jmD0Wl3rQ+2ayou186JCj4Tx+jf
w70hvIBM3X71HfUxormNqNVgU3Wez1ZmNr7aSeloIrKFlZRFsrjrO5zsxugtx84q
ZHmRjNvIP4i6xhURPUug14mnS74MZlohcglutKewa1jL7+CC9XFod34KOCS6dLlw
xEbyg2ZpGCu2Wj/mZOJTQyTT1WG30tqlxRCCyZiUFt8WxGijpqoD5I32p6paT0Sn
5OuDCWLFRGUk5SiueINO7wcLHylpdZyA6loDyh4558LUQynkDzmwJ/my2NTCrgPo
0KQqp1PfXLneMirnXAkk4F8N1TsNzmhscjz6rk0drjyArq/zoCf3mtMod2A32rSZ
CP1feuccW25YecnfOu/CXh7wSlltXjqtbSG6YhXXYQHTa11fCttTvzsxvEJ1SOPJ
abEGZa/gbG5bUOgRog/0JLaV39rCe9x4eu82Ug24m38xrX8bsvwHwDqvzolrK8e5
L4N3xkCVFJodkIiOsR+d0GViHjNx7SY90AZmmPtehLzxTUJcOj4UtkFd9ACsQxWG
ASLGNQ4CrZ6VorfetfEkHu8alk8g82390sTvIlJfA7PCuv824y8FzDj23tnvKtqx
7qR7p10/OhP15n4fCVQTdoDL3M+azFWSdxGqvL1HNXYVFPH3TIFSn2CbED7HMnWz
0rlMSYBjbk0MyEmUjPwbkIrv8y5fhkXcDrFliyHqkCZ2iWMjpzybV3+C+G8DPNBk
xpk9Kj1EUByagzVM8gVuM+o709nJwillY4eWxgY4wRDSci9gyTm7lIP8e4UDyo/Q
rnw1TdWTCLJoB4V723zP0OQbN+VWeguZ8CzGccULRXmhx8V07BEEmeB6AjqG3fgV
zyHabkFAB0FZHQLoO0cDjUFOZTcB/r+Jqm634y1GkPeIOyOxzWwk0Lvu6Kx4ZyJI
pgxhuq8xGYZXfTczqjwVHoZKeIJFkikzbCDSnckf01BEh5nF2FGCfnsw+xIl56K2
xvhIluY0LOnWARtNW4vXBOof4QemieyrLaJZ7QYuvF0sZEpw+AsAfugaBZGP1nqy
KTqtCeKaRBpCGnU9tANzkE6CAXA+SSe1gtkPkQseVxn7/HOzTQ0+wiV6KuqBwD7N
3a0ap35SBq57d9H5O2q3uJWRHwA/yCW6a4B52V2g4OTB1o61mga971OPIajsbb4u
BYdcYHojasaL2lEWxeHePzwQvZxawwBChG1slK8RTMXcMYdQYiQsvQBTf1Kwqtgk
7ulbZ5+GfbFsGHqwcif9SKGcgHryOoCNuDjZagDpXONYAsINYwgo+FHoaRzgX1Q7
GecIVgD8r+EElKl1+lRmpH6RaFIZb40bAhmh1Kz64uGgXVOLJMC4stcghpy+CD5T
XEK7oRoexiSIVNOWHOK9qM/6+TlD61n48e/HPxb71dezWLzdY2jxxDpwpWNXXAMa
eWcEWSXza2SfEBZxX445MU/VQFyGwPXrAXSirmt6VCdMvnt6S14W+WVUTsLuevKH
JpNtIOTRre8D19+01ZXvWpPAHZ6n8J4XSWiTrSUF3sZK/mv24hbQzG4Y6DYr9RaG
2e1lirf0o5H9yioxLWiwSERG7rfjqvdHVJC/POUYYTDZjIHtDbRE0iyLEae9S1GU
bF5L6acpyZ4POD2f/K93WDjbwMMmtevj2LwXsrvyHGLT/oSuVd9Xt5BZtf8zu8gM
kZUHJrrizVv+vp+pHtgbEGZikTELpHozc0xe5A9/4yXNrbi5rbOgZ4cNdTi7IDsv
s73Hf3uGVHNKtPJXF0DgAeoNhhEbNiq1PGbNivNG0gBxlAIyE4vaMAbO4dS+i+uY
QQNpbjtDePZ3ZEzZlZXhHwlE4cYatQoWj4e1Z9CLN+iAA6hISqiFdLyhNahebkwO
I3zgS3Y3h4QP7UqIfD+xh1dKaSVgDxO2t5iwDSbR38km1vjT1hxk9qj/+Rs1Fwc1
XECc5jJHp9zO24VIg8KblSXciNKKfhDv2HZDqA7Jt5WSiP9XaV4vcLBJgQp698co
/qkFSjTxSgns++RU2tXnWYaFMEnjGZ205L37hMD+BdmGHHeBEovXLkBwPF199uRK
pvsVmUc4wn4F7IgQS/Rm4tjCLgnlWjzr40n/6NxQjvkXdKXvDZldGNuZP+TAk38E
cvx/gJNLm7mZ2PMLtBM4VENWrJaIWmx2BW529bSo0rAEs3CpTqSVp+jCl13BNxSg
p0kO+ug4wiKXf+kDH0xC5N0plV9ubzH7G4M/92ojVErXnahJtG944LALGP06SYeF
/Ear5M7Xg/4s24jHTW8LRi9wKNJjvJqndpn0B1WRAJ42Jf60ufetZE2y4ozYU0c2
NaKfop2IWBmTyQvTBfTgoITT2XmgRzVgGko6/e6qrAHSvpA56Ej4qfw50lx+G0O5
hdVMRkNIBwU3IK/rJ6dRSpJrtnctAH+Tpke0MW7/wqY8kMi6DFBmtSSYKavvEMil
VYgAiZb890t507BhpzSMl3a6ObNM3BxTDrGkgXoMP/unqQvba0X3qNeHWgkfpanc
7Dlu54cwuG3FYEZQtg+dRHUxa3xi6rbtB2q6wzfdRwlj5wbaVjORgBBVitXfMaHj
x86BA79vL8vLuVtpNFdO2KKLIK3XX77ZpK2vRdiAvjnVWGvYPlgKmrVM43rpq3ch
SHIY7uSW7izjAIbh6wUyugYX/suu+laobJD9Jsas/EJgdhZq4xxJYg6UqcplPN91
VtQXeXk7iMqZsLFd7jYQw2qdqI/1b8retBupw1AI3OrguT7XddNWFzVetc22iO4J
Jq3zxGZPpM8cn4M5XzZUTa0ACP0MvB9FNmgS1z/aV02jY9C9KrtrW/eyXNH76kA9
f/LqZFNylQ6E6OLYkjYIuSzNF13/4oCeLwsGVh2ORwh5MWbw3gaqIDxPRmS7IrrT
2KoHFEkWvIiENRoUGhzw9A6T1u7HpxXupiwohwc/MSlvbe4qPH8OMpqcMJ6whhhw
mqGtuRsCtfxAZLvszqhcv2PVWE2P98niqo/cOvhlZQZcPdYD87OS2QqttqsFxxUy
xgfC7k1zjltdYUJQ+73M6O+OK1PaevCAwFjQq8kvyDznWWrSOvZ09RI0BYs1SvYA
XcR2/2H8B1CDItpWbf44Xya47TIitHH5eKAQJ5wyk4taMjNOsPodVoH9rF3pZC4M
p3OMI9u1pCx90CEm4GT6F+OaBwcO7ZdDRg7EvfZhZXWg83NSOM+OI7pWJV9lSzMv
UWnSFnJD0L41iP48CK+zHaOXujLQtRCDdJwWqm0IVuarg1ifb4Ep5wpBHbWQaQAM
Ssdt/gTmkTTLr9+RRUH9RZNP3jtHK1VE2mhEU/s35dyDW7tHqUeC7dnH1wT6IrfC
l+s0sZkzFapdgsvyNll1I0LfrbxK8XHk/aeqNzRljymXkfj7GQXbDCbx0fYOqgzD
jabJe079abThsZwM8jMRKyNeH05nws9Ybk4qA9JZg5hFhD0Zd1Wn7mWjBGmSoLJI
gib/DH8TfPJjeNCIBS62vxBUzkliwk8y4rj5qTSphaFr7ZBQa5ksEMQQH9LPKVWz
Ir5rBLqa/WhYZ/ZtHAQ2/v/3QSC2I/d84A1PD3dxQVl7XNph2Tg0/EvV61qY/1Kr
VHErA0nb6Hz+rr1WkOwYzibnImMTE2KqkpWs8Bsjf1sz+JAfrRfz4Qqtzbqy93wu
hnXqEDQ6U23urg6+FHtwBCWCk8vpmamsVz/b4JYyey6XvlDPvwU2MyDMYMnnVhvN
XDrt+RllXJgnQ+dQo4cgUsbAZ/JkU0QCQidlN5H9U4SLPZ9bTCxf7UJf3R4FZ6qq
Zib+d57iMp4qSUanX6s5cZAxDJIE+xDOYID/mZ4ZrBqabZx7Lz4NLvg/wKKWus7K
tRkxPsnvzFUkobikGlibbfSnylwjbcJpEJ+zF4jf09F0m4WDmsNyybOiOl2CzJLp
7TXnifho9B8lKvxi8VJkvSpwI37LpjiK1TwLPwx2UD1eDuXbkwo0588zNWRI96iO
DMtmtl5pXgmyTe7VU4YHhvWutfKtXm4QC/qg1AAW44ep6GHY4VJEjLqjISPql6wv
eKmADGpr4uwjWkEMjTmUr/+3ipuDn1EWCOih5F4V2ZwSJL5jv9Dt1gXxAAI+Ukx4
qb7ZreVDh1GY5sEsjYHssGwPOblt6r83XwglQmmguAOEENVWybKFxb3GhxihJc29
ArQ+q8LkGxFS8ulZj7pXaIogwbSeKQvRE5x4tbOrK3stfUESRZbbkHIHL8U4raQn
0R2v+wl+L2XfcIgchSFe+4l2cFh7gShkOrE98WBXMHodq3spmuud2XwKZqVr/pBe
FxJst43Hd3eZhHZujjvtfVgJOlDMa8DNP/kKQxiqDbfBaN+yIu8PsPJOiDGeG+nN
bQU114PKJ1AkPFQO3JhePp0R4tUZmrpWwByy70R6KhoTmZA2K0DsIgcrEdGXe9yq
xMaodhP8/zUOA1+qzVF0HAD3wa5NtEZ7atlBJc+mczYPRNUPjuNdTNHqwe12Z8yf
paVirfnyB43E/rLp6ZY2fZbsbL/tOqsXAvJBRQton4ugMVooyNOVfqUlFTaRO7fH
E71v8OMlKSPRmCW9Z5ZZVEjQLQSgHbfBcVv661dPiSKNpvKOQCAKX6efwwMe9lYH
zhX0jLEgC73YaskK1AbV2najIKQ032p+ugduJe5IOZ1MtQDEBpNYL38FJkGnMP6d
q6lTLRyUw06riSVxvRELJYi7vLurwhOEKbn3Vfj0whzP16FI3tEVbLY2vEgmjooP
EdBv8UvrYNTYM3eDtKTK8ohp4xvxg+/AqXVgOhBAuPl5MwDJ7nnv+FDYkwBP0JIw
XfDNqoG1zbeej+uTx20wqYQ9vqlPypauaQZHVm0iBU4NTz4QlRbNSqe2YMi+T30P
/yiVtQXZBVTWEp70pyUqmObgJTEnnJ62j4cC4YKNBlGf5ncEER+1pmVZMAPHl1h1
vQ20zN54gzEV9O/7SDfO3Fy//2XHHqH23kqFvcSMG8uKF8Xz/y37+U7waCWo2Kvw
NhBkjWbZtHTJJuSDBgCQwj6Sh+jSnHbHa0rfMs5VfyDjq0MtA7WRNA7ma9Eqd8ah
TlDgpl7Sgg2i/aVsrc+NQ/wyp3kZ7QBoRgw8t9qbJ3AAHj4Y45bCrDnnxMLkC8NW
zp1PrhQS/y3unhBEATYdvpfg+0cDEq4NrCHnnuatrub4+EgN1lITs8EF3eohtsvP
pMXnY4iQYEqZSWp0O8y7lbLzBUomGTw+DmCqN2Fg81NDKYd98Ii2Vw9I9bzLvOdX
qPkG02165zmCRa/hEEgxsq7ZukFXexWs19TvCDx61scFelaU7VQcFwY3PTula1De
0OHcavdNDj4xghnq3nhhQAHndZOm4EfZlx0lb8OO2NBgqK6LNj3fkFjHrdw4b3g7
FOcaD+pOivyWO7dd8XwlmCWb7ZK1d07BC1bTwlilSSFBhaHuLRLldF026SnMeZ2V
VGUdCUvPYXYhqSkSxu0v1C5pr2JBfbEFf8IqsBMessrCStakPQmYPD56q4r7DeQW
+Hd22EGZejLGUxH+q4yYaWUjhaf5WgnD8O/EwmrQ81AhVtubXmGxsF9E9z8hTYli
SbJy+vUjoRK7+zAQLWJ+9D+0dLgj8B4uURW/QkWhO8gp+D+SeQC3ZzRodJFcvyDB
XkijPsh6YGh0zBpm67jF2K1IgpRgJ+zM43QRyqZMhVFa8dWlyUhCzMyISGIG2A+r
yP6PkLIqCia2WQHoywtqffkvh1z82Inv0Gmr+LxKdcyj21b2paQ9quPr04vHDOis
mlm/64mPQDCLCjaRoZ9p/XDnRM3DWSUhl2G3nWK5d+VjXb4wQgM3PsnUVK3CbWNi
rOSnI45xsghSd6fCmvwJNt2atf0ZVn7DL8WojhUpYmz/gOQscptytmUPE5TGJJWZ
qYQdxpV4YxE9fhKxoH5JwU7DKWyki6komtuahOyHWRpyowMwVm2NiUcw9UaNi5CU
i9AF+TLujviQr3LK2hdPRol/MW0OdwMZMHCG/iprQmN7kGp3+t2Wh4MxbTjaViKG
cpW1fmbWIGikV35Aydt/BUSgUSVh7nUrBNm8CJinZvkvP9wSHjDDVkTscEPzCKyn
AYItQCeydX0xIJrrTyWhQQSRFUZU7qakgdaUEziCjnJfOLHp+KDoCyEQntBjwD9y
2CFPFl/3lngoVnljSU2feYctOMn2KOsHltZOv1W7nP501WU0hi3THJVKMnjMIVbL
81kwoTWd+qNNAX+0cNXePyDc15PCN1fB9sF2oyPR7VKf9mq84JfYKWN0F3PiAyOQ
OOZbd/T7IQmcWH3C9za28ut7aNhGtEbHJONugbKWmqQotcDzk/ScOIP/mzs7cLwv
GN3Z30iioNd1yMO8IozVcuxSW0QfVYFbQE0PyTonQY20sCn/9eSJs5AZpmjgb+Yi
1cRirMFrUPngWDuWmTWZvmbcdLrYYjDRYRYlvD5VUbuVDxoklgGO3PWRDKnYD01W
1aKb0EWwtfyELHxnPDn4J164cMJUc8x0QwPdHO7Zg6XBqe5OWqwSyzzZbYoOtWGp
ZFMhPO1wdvJOuYf8sUCOkk7qB0ejpyIu21z3XVWBYNQEITEKWUCdd3gUBfR8tCaF
5evRsmBgU87bG+bDzFSSdkhzzDr05kBRqscgVU9Whdi5z6vPd5dFeHnnzcxipnbw
yhWf+IBgq3TmhZR6OXoFeZcKJZyIQrwsHkrIJ4XMkBrBfslp6pQh+mVCMEGXQTde
LDpJOfLIcFZH6Rkm7AJBQ5Ny5rqosH6O53VYLhvNitH1XxkN2NF+7iSVnVboFoVZ
CxHKygy0brjjpy9vCcaQaq9aElckuACQCU3hYZsNTcFRL5kckvlKZSFZXESp1Tf2
mM1OQd6TRmIAzm4R6yQBgUYhvCwUoYyICkb0NpyIH2IYd8VGLN6YtOmW0Nug8XA9
K24p16FFC1WbFfTLr2swg5Oj47dyhL2HTd2IzyG8+ecD7yfKVr/vwcTk/EDwEuwL
jnXSkQb1bjUXV3dy6IvwGpMa0jbi8oDQkuj5EbbvP87C+ENMWj3+QdOTxyIMlusM
bVziDAIp4R6eoB0A2OsUF4UOi4ZT4zpqcPf4PRGyleUOYPIsCnyNdsqRfQCIVVMB
0Mm22zvx0X0gcdhPFtUrQexUgNflqAXT9A+hOsujVR9bzSuVdpjVKoueenazC4I/
b+Z3ivoueLu5O5RAnrnvrWKxCDuX4fNLQBltTMCWifMcYRQxyvOThHWQ5n0I/d1p
2W/DbK9C78hEtn/EcRDokqhGeVFVGt25+r+uMWl1IWEhqNr14O34iDDmOZR1xz4x
MlIAjGjHdsPG79PodYX8oXUP3AO0ozttrSCVsL9iSBjainsijSy6SM8J8HJKg+Bn
qhdziNRVZ1vc5IKtki/G0+4kHxheseG65FEatpvQ9dMbViq8AeVGpKVGO1KjvkdR
I8uZsUg8r2phzX6OpzdKxcZW/O5LQS9hF3JSpg8/32bW3DuAFLmpOOCg4W+g6Iw7
ydkJBMwv6HBaaJCDzPPyGHgrEvjtZoW7xlgoOfJn4UFybwUz+1fHpkyBfApQEuxM
66XwK2eusCvN8r9Fhf/rMB3MK2jYKo0Sx4jLkoUmNlqRdarIjSIIyw7Q2mXZXCU1
rX9pcrE10lU37yBiu3MwbpfpzzXhKTfQckZIMy2anQQNX6A3L8wvuAz+vNls0AxH
RDnrX3gl9v3IS5ddmbqihCK4s8DJef2tYACVIPxztBwQ9BWDmzryjxF++YvPX3I4
wzf+ncHi31g44vW825qrWnN7q6Z5R7A/8+sZDls/hflAb7c0pV9JE+sgMDZuRbLe
bucg/89fHnMs+O/HqMO+WmVlcmXqzbQeRnLZeJWb023ettHGJThiBOtv0ODNu0YD
XKp4irz691mO/C0QP6kQz2a5pylMVBVAmV168Lo4uUDD05JymhazhuvuwY519iir
IZlyessWKSqcKy4OTpZb7c8W4MML0wwklPNb5xWXljunqiAOHPVV1DqhRzSLevlJ
HzKG5iFV2oep1LJNOaSbJVgesof+rwVMgeg18AN/ghGrPFCCmQfqvwKUGIq0k41B
axxOHctviPfiHIYbIeDJPQ5Ey2TJLhTNEFrASF1nBZp/eKLAU1GR8vfx2SFFPhxK
EFm+Kww8NdPs4y1GcpjXkr+heqa9YH9YtD7pFyZ9fgQJDlX+iwqi01FLujCSTeDq
aB59a6p18V9mMICImSJwfTH1cICV2OKpCkpUMrhIJOaXiexdh4sXBy1WFzqbW900
u8aFSXaxGHnTJoJTmci0AiG1Z+Oo4nqxE7pHIuGvF+ljOKrky9BXJOCnz1l2In+p
07YgpieFvIZjaB/l7UXpz1akM3FWSOrn0/VmW9uOVVo1Z0TiXpOa9WwEYDogtRT/
8+8HTv6+UIucf56NNmmPXN/II0zUc0DXVVhwOI2YFhfyQicbsxfOwusMdDLSDzmj
VjPzFR9Y6X0k5Olz1wt59IU79bmsRcYtl0d9ec8q8VDaUhNRv77x73+56KlOLOKp
DynJRUPlFfISR7HQeABR8fTDBMopzXecus8JsAg4YIgZnL1RolKzD5vL5IAJk7tD
wwpPU+E9LYS1NXsUSd44zSvs5cojyE7zwJkbdxp9XP4gnWus8o3Q8eKE9uV+PPQ7
uIO/NcNBj0ch63DjyyLu27R/6D0cdMs1Vj/cZI10zOjBQ4KyZWafRkMkcaLkJHIU
YHpsGofgShNJPSP6Uq9yMdZahlTAaZ6IbzcxWLfrM2di+eQMIc4VtAZzbZnuuaMG
xK8yVZnM8UW3PBZ2stOJrQICEQK8NGcHa9jq0Xp1FbkBV/sNkpOXIApYm0pAvVgV
tvdL8tFjvjIalMjcuVL4V0bYtl97+UeWdm38RLKY/IRJRm9/clmiSDwl82VRcQuT
hSq6CdC44NHDFGdO/jMgjCJ0aZeqNquLqI58rgHm5Ca+wB39p9JeoBDjbwR4DZUV
len5WHL14e8ZL86Y1VujNjs3uZQAKeAi/ly7SMxbbioGX9eI2wPLH7kgOsQDqk/o
yiyaofOxD4bMf1qqNLZVki5VDc/16qkpopiGYN+DTjLWuRYDvwWcyZuxSfLmqF5T
gLkIUMo6P3sq4z/oAn3su6PdUA38DPK+okCyO4DFnE306i6xdVu6aBBVshtyKY8Y
nvJyI3OrxeP1Rzghyp8WBumbH6EWmEWMX0j+ydGU51M00KMl2GfAUR62qYlRf9wl
Vc62FHItH8kulnO/prGH866g1d/hem+IBBs13EGeyndPoghrB99mWVlPtRoAouOW
VbBvwrIjeIImR5AOTkgqXAt5u6NJdT57E2g/FmUkQMrpgXTnBwgsVN/cR5N8mlzc
2knckkZ+jj4/qppfW/E+OHt+QYCAhr2BJ983VFkdqsWVCjt2sXpe1svBOrvXQy+x
FgCz0ztYRzPIezFNciIxPAPDP3Zr07WncLR7Yx60ytMUfP/Fkb9zLoFFPLaW1ET9
n1eLrAihRab7up1oJng2LI2dW+RAOAB6iRTps2SW7iEEkZDPlmxYSWgOMH4UXvuJ
Ha0x1EgxhtjPZ+9VgEXyl3FCdYKMl6tw5HpOH3f2hl8VrARJDEgmVVg5umeZyAHz
M3oopWx+gwkdZ5l1kNAnstGSFBjbhJg+aZBKfm+uueUq2L1bX8Z1iYP1DOweat8x
7S96R6NyGg0dWaCqU6zI+GHbDqyJDumIl489i1FgrqcJbxYGlqRJYW3z4lRgbg1k
u9Q2DJh42oORI1jeUtJl86hQytNAyse7jy7xvUbtCHuEEPxzZF3D9qv5eraDw3UA
k+4AH/h6PzKVWfb/VZLBm/6F8oifokcDJeZTkk5BnGej/m3NZlPO790N2ggDgsiN
ziGtHtZ5RguhhNzbI2HPJbq0mhxpL1x690N5UEtRaW1kEauVvTBmbof+1uP+4/e0
i2WHWB+Fhv+mKZaHREz/+cKimSdTaOOJH1McrvKVu8DemxTO6G9ZVrxTouObf7F/
t+DAvQmdbr3FOyjb+COk6MqKXcye5O8tpaYJ5SYJrRxklp7CvAUfB594b1CKFJ6T
HGSZG6EmqnSafH88SrhPEtWND8R/K2deV89IdS4uc03MrgHGAC/He9BVTuleeysa
4LPYZP0+Lb1pLe0Bg42V9x0Kb9a5RNZjZLVNarV9Ua/vRgA0XXU0dcsVASRD2gfR
hkDX/+hoM6TyHbJkjfSxp2uMOCh8Csi8f+hDhscAScS+tgfN5djuyqJCNnte7AFU
LZSoJXnNcT31o2P0vjJaT7BwG/3zd5Zacc2LQuph1yHHcs1wbUH1hXYpWTlWOWvA
8ZvDtp1bRdmgBVEuaA7oeLlN46c/Xm/Ci70UNmEXeHbRQoRT6rXfHdJ/h0SM1jf2
ZT4CFAI0JduayjoofYNNioauxT2MXQ7V2czDOWJ0ZWJdbyJeSCpCViykSw7sAfk9
xhgrreoadXCoV7Fnqm0q0Z05DdWamqTNOEqrE69Xqrtgiv3a+H93R0v4YsiNrhJm
XDYy25taaXYWEsIluM6KLWgnryCUWAqRQOVWcf63hW2aFEMUaTCjQ1QvfthC7pwO
4Q9Ej8FgEASmwvfD6xAlkuwjsSoy/EHUu1i2tJ+RrTsiBMw4Q/R+V4P7myNAkIKQ
ag1bcEerIQM4VIRRYBcVjxhYgsOd+7sI9vu18lb5vLtK37goQTslBtbvu+n+GkKM
jvdIK5uZ/rAF3iI1AFEfV6bfGBreJT6nuSAkS9k5ZhQOqCgF5abYLXBF2noUe+LW
vmiF2uN6JJrTfDBblaD61qfscz6Bz2Da15rCWJir9pbi/hRYWnF+Muzxx8sdoxKx
ZLfe1kmJbGNPbrS6g3CvGM2OhnGakVsxZmv121YdH8BcRUMzT0XHu2dt3oSSXg88
q5RWog65tDyMtx0w5em8g4DHk0//cNibCU5dinefQT0gMx4ytTI013QlBSKME2uv
OzyaZ4X9ZtoUtz1XxcJH1Izkq7LmJGMR5RLH8j+ipGcsam/zKk1zdCsAQsOpR/3D
3yhM8TIR91C6Z9rFgCURNFaeQqqmCi0pPvj3DvjU/o7xUr2IUAyEMcRYs0b22Wwv
qCcYJOC6qLkLDQJpClWoM9ToAf3fEN3Ph5EHRO+/ick4kPvUtZ5yFGuta8HBtk2q
Uzh8bAPy/gN3Vyvs902qceFHofBmXM8bv4nshw/g1mOZdntvS0OkWwze2JCVjFo8
MtnJidHcWD8E0+srkr13Ksvhs3IojUjhv8zAVJeIR2J0Sy0lr3Ea/n7Mb94t2gBe
A+i2OxuMLr6KSLaAoo7K/0+hm2FygtxSS0GmAvychP+Lewl7HnkSFst+qAMMXnBt
M1YRWhz3CPnw22cuKePdsoyTvPWSQ91cuasgtjg77j80WVJwj2t1KLSm5lbgDX54
B0wNVhcz9Bn3HnPiMWzX3Q9h+5jEBE6uNRGcsTZgfdlylu8VdU7g7Day6kJ/7fCr
ekdueFL4EwsRPvPca4tNrDs2bGBDPz21LU39/oktRfEyiKS2YE4my60nSbRrs1Rq
D037fSJS0IPzoUcbJxUp7p/R82ZLgaWVLtUeH6owhRbcxXh4tLoC4KRGVQmhxZeb
JGvaKiteeFRew0aRk8tSLh54uz37GOuxVBzechi6lUJ0cF8nxNNTfFmplSI/c3Vz
8fPGg5FJ1zb1ftXpbEgMtYZVWRUEePt4wQfVIVYBANym+L3uRc66GG66FfHNnR+V
DKdKDnxG3zOSZqYPxtmaFo9cScctn5vVv8YVLW/jMCBjnCqDKK4Gx5N1DfDhu/1l
Cfx5EdjycpTnsxEz7dvmldRaB4vGYugz5rAV+1IfzxKJDYaJK3I6CGQUvjEiP5yj
oQtQIWGxg5E69BZ5BG76wjja5ZBT0nbqqez3Ft5mAJQDpBzU47qy/F8Es+FeGwIM
90M8ZzcMGLXwPqEciJaWT9oZc5xELDIqUa+zEqc+bTeyJOAg7J9SUdRoQI7B/lWO
PfscVHWR967EB/DlmA8YRWSh2fAe8eQ+5hINFJJubt+z5C9nBvthEEoPQVlrQ0CB
5ZjWs8fnCv6+5XRpCK9yKDkJem98SN2KO900EbcpGNbFJkTsteQ3+ggSrdox2cGZ
vj7qQ5mZHomacapPrlSaA+F4VBSA7MKJh8qlsokf6p0jhMI6RpeRvSeAdXxfEShV
HEOydXuwzrgedF+MhTu00vxnn3AsKi/xiISAIOEYrvEusulm9S6qFPr2GscBwI0r
+NruEsx1EARbZdjB62eJ3WwIXOUJnmJ1j2V+zzkalwPkhDLyWXHKPo2+MrORI/OG
GVPveIes/km7qdO4h4ZrXJSXoiwVYkH8+4IG8aXx7LVwcru3Dbw2x3tVx9YNxPc7
L4Kvu310YFZ7tm4ekDnsldF2QFd7YFOr3UVtuXhduxUqZTsOVoEOrq810FFhJYNq
w3JNhWrgj3jDDoRR2WQvhOlhVpUPSN7HhOMCUwu7VylXfs4db3CL0bszVMVAGAfl
/blzqZkge6+GvkXeni2RAAAmA0mN7KObxUCeXk7F2fQAeru2JS0I8Hzg1ExZvO9L
a16NckI/ePkvBAjm6K99rN0IJ04yoyO/iIwaU2x4BddfHlfCONrGGy6nanjeR9st
W755M8S3PRFSexo9hJjG49GtEvGRHEdbOl9061RbIrRJAM7XJIUxHgVVl4Y+HRup
JrzB3H4vroY9ul6LRGeKMm73DOtswsISWFzllUjAKh8A6DG960NX4NdCRd7YeenL
JN9uqDmIQdbXUHHSGXdZ4u0rI8Il2aMatar1GIMNE6eWtmdNmV9qSq5OQLpNi30R
yEnHUfHxaQyg/tWlpCSD7m1zTP/Z3XfZz8HTO2lfg1YHUkv8bE7TsjCxydhDoUdV
HDzZii6YvYRSwbZH64H5ENsipv9ttHjMHDsZiwhy5s3su4V2ymM8rTtJ4DEiBiQx
Dql/+KBbU4O16ZRPgwK3U198s1QRk3OtDUoNGoxJtTqxfSxj1SbgBhCjc5vg7r+V
OMZkCDIUlOe+WsIpTAwHfmaPaQNzAob5kx82AsO4JH5pmjHuT46tGpP3m5M1XhUM
izwl9qdv9avtHWMK//JE4x8EdY6YBuNHZh5A8dN3/sRlOa+LjY67/ifQvnMINC3q
F6lnzLcjwqbyksp+JX/rda0e0thwaGQ9wB6X/S44IZvn0SpmAVYD7pLWyVtLgfto
4GZYHAg7kHDToUY2MDGGATMr1USKFEahBiVPYJB3I/Tlbx2JOzgjUQEhdQsDoXbX
j2QDaNpsP8E3OzBkPa/My0w72PB7aBz2TE+SBlqjBKheJtqT1UmKv5lC6yFp804J
Yb8dB3E6xK/EUqynYljZXWYl8peVn/VJa3w/wzWx3YoklCKaOVB26HV19W5iDkXi
oIAgkLmCrbrl4N/9cUQA4yMiSO35eHn9fscjr2rNfJbXRgcAvSRdtJdTchY8DAmr
OmVlbb89x6C8LkJkp7KLJ3IH5KXVO1B5gvj6goYpAMFJ6SKZsM2tmzzeIEYknNdR
DmETeLEWKeCTO92WUOn5XrJHo7TZ5juav+2AmY89bRowltC77pbmH459GnuQydPw
tjs1XNtsQbbPN0vWrztxk1DnNnFAGEXUWSTTu/ARKl7Mng4Wz5inKCbCzzfsx7WK
Nc7ZMk2/zqeO/XOOYTS9Co65hCmGZSzlvXV68s84xNvv0sD0ifsq5cjGkn8aeUcu
ohySbetDwi7dL7mBS1ttAfhrI/bfUdT1aRyf1rN4E2x19EG5KEU2oj8MEMDvTbZf
rPas6XW2fU2V60MvQb/pFQZnJicn1zCew7/B/ra8AOV1j4KDdcNY+SvoM7uCExJI
HHlh3bOjwJOoOPSv3j/feXsx/s26ihkXWZ5U7kzi3BV8S83FTTdKz1+uX29HDgkD
0JZPLiYVRiuQFilcjXro/fq1WP1o1xQ4f0iKZFafrZUtuLXcw1nDUjzYwmMCKPYq
yvx5XM2mdySkyvHn6yk6qFgMW8TfE31rPHAqNV5nITm3XI1B778BZciFhMLZHREC
SBfDDXD6iqYrqysEEK9qpt1AKwnxmbRTftYWI4JYYIxPek6XjPHhiaNqzo/mOFf2
P1qVyD4/BrE7fne817B15W3z0lV2QR9LUREdGF3r798eA7XmDG8K+uoroAJO5Pua
gVK9tl1wpDes5377JobUjRpXGB3G9rjDHOLs493Pr0ofoBPq/SVLd5sqmyAq3dOb
uJRJdhz+e/DA4D36PPWUK9r203rBZHTq/PlfW7otlGpT2S1/t6A+ETRvltp4aLtB
Jjo9ehZ6W9QbIcyts7G4lFj8qfHoR/fsewlpbXXRBc9sCOgH/sMJCq9RHBrnSga4
7IeIsZRN9B6NMHMz+wz8xut1Fk8+6PUjAy+LMVkUwVvujte2+RUwcTQk3afliFM+
5kvCb7scuS6ISBqc8L5voRsrfGDoCRCaThaO/BJQYHEZ+kPe5oRf0HdSyA93oIWn
0S9YTPGJt7A+zAPwjLwCRTCsMEQMbuCwotQozOvGRMW2yllptS1B5rvV/6TMgLUA
zldnd8qyODX6qwcjImgquymCxIql/LbTyApII0l52VjHem/pUEiTRC6iE0KZP77u
9SrAvs7CJ7pS5Q/ZAUb/f6s7Eg5XIQO2MMSJvQq72rvEOAZMHs8NUMzWMZVLtnBY
F+MiaWbAUz7ZNx4rH0llbR/nCZJCM+Wi84do+oz3QGrWSBNnfKjr41mAezAOMkge
IXDZJkpx8hVLN85Rt/lqYko4XIoyQo9HGINSLuoL3KSztfrw3rwhxG9SbET1at/K
cMAY72uAV9QGXv9IsG9heqa43Fa19gGsFJFgB25lsywAg0sk7A6bNw+dnWioCT3k
YBmJGewQi4cGKEZ2QXu2/m+Qjwh0VAG8zU+oKhBnTMpPfpaKmmF8h609TnoKmElW
pMRR0X34Q66RLGvFPFq8yvAtVrmE/ugKC4aybR/KMsLJXgpmQlm+oJmNNs6GsPaA
aNdJwYCxz9UkxzwY8pH2KvGtmasfd8oBiRflb9aQQQ2VzKJzSy2I2OA/NouWZ8D6
0ECsq6hEksatYrVwCCxrTPSOgdJGfxa8l0Wd1ejRYWEp56udxDt14Lv0eokWtfYo
w9EgGGv3X30Lwil/5ymWKYmBuH4Xj/LG/Jxs58cAUxtnHyXCEsxSGj//swQgQqv7
QgtGkcNyVxO2MibPug3VxnEj7cPFqrCgU+y9MsXM0iKW+JI/M6N7Ah/B1y9orLQw
dc7VCOw2f6+V3Pn7+nlBMT71/6U9h7L5jgMwW0jv97d4HELOl6YYHbz+zA5ttU0X
52NErv+QdjLiAFDPXwU2H9ivHs20fsNF8n0m1pjeOQt8JxbfOV3Fb5W1JuxKk9eF
ew2eCJtofYMT+VRfRPEtAlj7we460C4NmUMNvlzaxmYpYk3QK7x6Dev1ughvV/tL
dZNAjH0GkB7c76H9gfoQ9hOkGnE99lcyXnEISaKHrM8a90wNLydM/lFrSwo39eJo
8pC5Jtatt+XG9jnVcLCsL72Eo+edQ/kfOkBaOm/4wGhBtl4cOHcV/uSaILBEvGH0
0KTlyScurAAraQZCzYL0kHUbFJjoIGtYTkFg3EfVvQWUOkMbD72lxZeIRZA18aOV
L7m/UD3+Zbc/NIFNZkSZUlSiEFZzLWUJBqUK9KSrlFTTTEsqdHo9GMtYqVHC9Dn5
cTzJE+3CVvdkPyDvFElgLg4VF6K6uag623yP74RDKKyr9p/LwW1AWHX8QV6h8Qj5
eYQ9x3nf8+FGOGdjEYKjojX062UhRT+hGpFCBnxtvEZwbtbFPikArZVcZQPMkkQQ
d1AXcAcQXq19pbGq+foKTa6fxOdOf+z58V7yj4PKz4U0tcwETu32OaA6KNU5qft8
aLIBgALikhcJeJ9AFsBar9JH5E56nE/k5bk5FOVknUP2PyvkNOSkXPWtLYst0ORo
s7UUSiOPrT5lZ+0GohnK/f0h1EBla+QczFR8rgCQnWsv4/RvMar/uBkYN7/nhJPj
rDhgP5sWlB6RZ3LvaH408lve2+/htF1OT4FccniVMOTRB3RdkscCCUSXCWdZ3chX
K3/HB20JtYwRMPY70J/ih1XdL+KiVyU8qATAoGlYYsYa1ekBUa3VyV2hi+dIKnY/
Z7yYxr0SHdmo8S904lk6w5Yf7ML5WMAgP6OGc3khpTX6Hj4JDKuvHcJGtsfBUPmv
MefdsJELVhuqURTUkw/3d4TGozkWjxpBpqmXxbjiCniE6SyrZqA+er3bwELSFe9R
IMGqfQaGINujRb+yZHXZ9yXY6QhA6QR88cNQmeyTDMmElUUZf7RWEv0Gielf50yu
I5C7PtFEmb4NwkgtdMcegwQrZdyH2FD3thVIEYepl4cCRGSX5Z1cznUMMd5JFxGs
6RcfosSsEt9KIzYKa4FnFUWXww3BXvl9XQGN3Re/NkG4jUJBEEGmJA5VrZvXC8SR
j4RYHMpANIfFjrW7xQxaPx2HANC+yG8klMScUApYXYvPUzhEzdno+3daLdnMEvJb
c+4qqARRAcM+Pc77mi5G1wmWe7cntJlauC+NbRiisCDlHkBj8mRbC6JjXE1D4aPo
Ra4IroiLCAUTYozsIB6y93g5bw9YSxdg7ZezNBXqnbUjI0yAFXGM6TZUyQUugPsd
zitkZ/BfwUIF/FpW3oK+m5eSEEohIUuCdjNal+kn5usAX1WuplpWoXwLxU92ngUY
YSP3VTEZK7Y7cM7416Umgu/tupcJb4QBfyUtthvEiH658OY7OVnABg07HpY5AGDK
5Chkwe2lLKECZX9FQZ9Qlra+HZjO4jNEfZO9+QrnF2+v9cY72GOEv5b+0Mh3okuu
nc/8ByaWlQiLWDehcXj2EyreECnJhdfGF/Sc5+LPMQjh+fl3n/5q6LDoyx06KBdy
/BXNFfOOLW5ZMQG4UUJVTewYVnsTUSePO3fvws6JiOd1WMOi5+oCaKD39AK8x2JH
jBivQXcGCQK9af9qneDf/cN9Jd7xvMy4oujjgfs2zr1Wvp3glSZyJHohgSEoLscn
EFc4h/1zlZlKSIs1dv4yw+XueYkC1/WUP6+VmnSKUoXTPrP0Up5uTVCjCanL4sDp
qTLOzH6NIAcnnLbj+09ubDS5QV4OgyVjV2wn6dk9yKhwNrh2Z/JXrRWTHNCczhP5
T1kikVO6NDfI/EvsvZOFUPi3EPuOQ/nhgz74lhFm8NgWYaPJu5kqdk07xXjhZ1Ix
X+s2zEfBLmqYGidopH2VQu2UreBhlrPntGdxRthX17rIkRrQ2qyQ9tkzGcXbujy7
AnqrVTke/YOop5pSMvmhmWHy6WLoFuPvFb7YM4qZfB6csaJQXA6zjZ3Sckc2qg3W
wGPFf6aC8sj1+vejvX00drRZIUSpt9dk/d9UFw0UlzAYBo/WVtZG2UR9Rn28Lr5k
mzyLyQ3uE1J8+i9dtHNY3lngPzw2kPVMmCYOFbnj7Cg/KWniCN8VO2ud4bYDC6UG
qMaV3+I4ur6KJrBJmqzeCMF/bevcaet0D4VayCw7yuhwSnSLAju2cu44q6dogAT7
U5DRsr5Gw/S9D/mJ30xwatovY0AGsTlIhSkzu390+aoKTj+pZsB1pRes0OTYf2MM
L9rVozyscvCTj78PBqbEAnmp2geXyeu+xoA8IaKyKVntlI16p8Kb3yzMqEEeYhK3
KrcWN6BY8YnXwIvUgML57UiO86v2H6c6Ywoh2TBhE9bIdv0KnbDH1WiuzsUXi/gY
JPXHdzgJpVgT85tNdzi6r8xrjeI+qhrOYljsNxeeV0dmKV0zJpuDoRYZIqPdhtFk
iV1tRfaiw8l8eZK3RrASaUyn2WApO8/kTxQk32djdO5hTPhUsVvmib4hU/DSLyUh
l9R67OnPo7mPFUScBWgGIBHnEPOR4cjDwsp3fFdP/pAW8LCC10S1GO4vEjgL0nwa
Q29m2+5fAN116AiOVnj1Bdg6Ci5m4vAE9bbu49Q2750tJYQoGbmiDPNSN5ODrLy9
gCZCNSwCij6FdetJ2/7xD8QJxGJNPVWPQzFO2+UFXYOo4xpsiCOkLZ/XVBccr9sb
nL8CiTu5gjdMoqXhzP9n0lCjwrN+sbRnWuqnylKKSRGbUP2xlUAL52F7fSXZuH4N
rtqdLdduauoXEEhKA2ZOwYfcpF/vZ8silrHPR8VALgeBwKQVpsIfiK3OvFmXdBun
fXoSjiY8sZW32N7pHLCu11YLAO9/vaUqdAT6CiQE5RS9QSsJVuZBEcbFFdOleiNN
EnFBNKpkPXfBve5EkqX9Ao9lsHfMHNEEGaTSGQdbQCFbXsXrZ856/nBA0H6dE/X4
OrNkkBskAPsMG9ObcBQNRhXcrooZ2Fr8S32OZOVP5u8R1ehTcVZPgQ6myY9S+iY/
fJhzoCKglaySujIKDaCl5V/JQiff9n6IfniPXXbjtKhx7PnqvG9uQt5oEHdKvoXh
3p0cHOUGGLS7YDGKkAjrumkC4/+x6YveL0hipf3eCZXG+j290SHuXelIQyi3GynZ
MUrlZvJ6inA4h8qiY+2K91si9fvLgG20EcHu1qSF2N/rH4K8dqCvC14FXFjWBvz/
zQfxNJWxh1aP7p07uPLXT7WU1F0ZZfeYyi1656mxIZBUgN6YSTo/KA/f7a/pJtVR
UcTNKvyqHmLKe+r/rbqo5JMi7FX+aEVfQQoBbUCiv9ziTbaxUt38vPCT3u0Q/TG7
XNCnKEAwq5IWe7Xw3L8PKAUuv2mY8EghIy9XeABier67hYk+4WjPLE6RrvnNU5Hb
RsmhtN4AmynXRAAWqVyR0K/7aYzUNG4bm7Eiqha3kQHXlag7dfMVEiDch4+ikqaH
kjO9wypikTQL26dh5woEakepdI39YpKXVN2gkBp9M6xLZtE+bloCXnSvaaj3NijB
0p1DXGatYwqKnJnsm3D0NzOVx01Ki4iJyGRKFqN+OIGYj2zuCG45U+/Re5EpS/37
kB5+cVkN/SNNgJOXbfze4fCyMuyjrfIDG+4J8rUw2uD0k65T65RF9nyL+qy4roPT
up0tvINLVDTMCqdcnmy8W2ckbHUUPwkgFRAT702zt1geMVzqkb4+js9h75wpwqRl
fH8fNB2wlwTU+IFFwoJklBb9hLzCq0bCcoVm75gdaLCIzAYPA+v9yR06bOrptZuS
dooCXa6TvH3tK9BIF/R9qGxZEVvumMwjaCEG5vdCqgKlX84wBrqHgPrW5Ec9Cq6S
Kkj/w26rjx/TUSi3Sv3xciFc1TwMkkj913MfNF/QCQrCFpjD4PwcWq8RXBgwwj2V
5it4gyE2RpE7itKgiuEf4ZyicPqmGgK38M4j009EIVxx0bylT58WdvG434FyWJfE
Nd+UaygCdOjuaKVSF+lZEhPaLQsjA2joU1o6AJeD0q8SkQnRroFC9EINv1Ncw2wa
R4doDcNYBrnfBu33a/sgUnoJQeGD2WLbecAwZ0lFq0aqzWsqom3IDZ8na5obcdhy
S8cgCEf7zRFDR9zy3ofai5E2N9ijXOkKdCMz8q5W8/RKcrNUfQuopeO19e8fEU7s
HS+rtDM1gcn6sVgWXAJpR3siBbq65bTHOucsZeXI+PSXhhfwtcckTQF0hG9qGqxj
3cZaiymZcTLRgfUHOC1wMNmB2K4SAUk+wW/aO7tZnTi7yI2PHnxbpiYLuofPuAIE
c5+dqdYGvpWN+xC8hfV4Cvv9XkPlQwx5KXadY86rlF7UmJxUNVejTTafoxNjUEgl
ezRSI3sGXGX6QwUKlWA/T6OjaDToJ/yNCAS6kZVN0h0HRx+c3t7gVmn8Ub66myHl
fPa9sOr43w1zWv5w0byeCfijNVASWlDaTA0zzMGQ0PXaxhkNk6C+o3tDaQcbcm7Y
Fqn9T0lIlZdW9qTp/Mlf+uv+0iaxXbtLxwXjNLrAK0rPESJY3R0Gg+M/XtmVFSFn
dKXrFymhIZZ0OEUELvdg0iiRt/xnTGn9kfZkQKb/Aqexmg1fGjLrvAUAnBi/2t7U
dgMzttWo833Q+LDfUruTqr94ujfu0X1+2dXzP/jWuM+gyn1O4Br8M4uKf3k6Y7kT
W+y56ptkUaahDyNa42+4qNUBa6zGsdMS1vlG7spRDgAoKog1EuzeCbH0XHH3Tfkq
F2U7Wu4O93S7vsjLo8oeN3Wx/jYwxd+UBCJ25ExpdbClp6zpOikF0VbBW0px7ZzE
F6viJ8nTVSGS+TWuFR5F7c0g36DH/Gf7+Oan2ub1tU+pDNbtgjyjPw8dDAn23g04
E8fPp1BKrgmJL/4aaqaRNgLLGnqEeJwH/rOxKtiZZoG8CB5TBw2MQhfOpVx/5FdN
Iw9KqYEBNijNIagg2mbm2PGrVRSOTEewO58Hhw4jRdYdTNsD5YqyO3zCHtT7SNca
bKUx2x1ByYYNI4TjOCSYEKbXRo4AZ8tXmi3lTpYEU2N4VuQVnzh084GaV3Xfil1l
pudjHm7XI2kSPdDaSXaca9nItq/XqCfWFnDicC0JWbvOi2HvfWwOdUlSpIVmru3S
SKgQNotoEMUuiACgc9hmQyj2CDQDEEO30lEDCYr3QE1K3hkJMAt9sTBe7Rt2kHfS
6uA/FItaOAbBQ0I3qujXzcehq0k1Ac50RFVu4i76CMUXv0rxvaRvoLRgIr36/+BP
vKHIebjrIqrakhdwk7MaqQmN7wFTxRjfwCS4rblhKlTMVYTV0JYOJCIgXlUbvkg5
1vE+dGgOBTVL27GQioRX3YXhJTOtfq79xtPpf1o3q3pErwDZDmQkoslFGy5ZWouf
XC45goK7TGE301Z8Qf4R44ag5YWzbW/ZnAVtjjEQSr7bCrgzG73y/BoOCAL8gPrU
s0fDtXELp0qjpIcXBXKcgSX2J9lpF+hDV1Fws+AOzAIBPApTAxcNYBImxLAYVjdy
6zRqf19KGTa42sg/pstvZrSCStP2n0nwTMqrim077EU+wizj2sM6EgCQdYAeMiEW
UGuUlWC3qZmZRV2J2N/KKCGaeRdJF+4Ept2zx1gDoMxTvaCOTlhha94xHpOt2HoO
uhrQ4TSy5/dkFfOk71SYj8tTTT3cu2Scy8rPoavvab3gRDIuOkmr8SGc1YkVL14o
Q9kBrHPl/zsUFhxLUxcithN0ZQCTj6swDF2zy6WvirovDK12WYlh5yjH7obI+kuP
Bgrw1yWRQDW1FChLyuacBAKn1B8K09UWG3cOugRoTWNvIFDAxvwWBI+jw317SBPh
1pfQOBHiqKj/HQ2ktOvKTuMByOqCViDqktVG5VSxrwmL6bqh2t1NaHdRO8WummqU
qe5P5hm+zcShhp/GdIiPoBKa87t/T+7LfTHOSG+whrfpzBbYFoxLjvCuto8bkfhw
suZIE9HFXmY0S/stu+U8y8ZsIGSenFmqeMKIkKdJ84cIiCtzpPS+DFgtGQQNKCEh
I3jaIsYZ6cZEpxKAqqc//LiPxvGIV8gUX0dqRRA859Ek3Ay8ypTEAb6YuIWRz/yf
UJ407/IyXaIGEZlboZUwSP8nJSgDiEwFMnO7p5rWjl9DcXce4ff8B/fX9X2urUKx
+S1uJaXerDvVBw5rHMLP3FaLfVM2SCCiWf1QBsCNflqgfDs9VJDpvJMDddLppF5Y
7NQSS65mdCwqvzmFjp99c+xjcBiaTQmxFSyu7YL3NiKOx85aTKmZ5CYzKIsoL5Rn
y4T1QyfE0ZYvo7eyK0b138Yhm0lH/byHTfcXBzF8zeMEFsqcTtX6y+aODytOiBkz
Or3mympwaTb4vYm3enkt5NHVpXpq1ZfEyjfCxFvX5wo2E7NFuQojZtEYwxva03qk
ZprcxyFnrvqP7lvURcjhVC8OEmzejQHVzdr4S1YPVy94R5zV2KmRHDF6mr6p5UGx
04W0S5Zk+Yq/RImXsfHnQYUGL0NhMePa9YFbWg+ZIJ8M8kypycKr4numfdUB9ott
a67fopykDd59kEwgd1LTgQgoovRETy2vVdESTCRjDWikAQKAiUxBVfgFJ2QYWMJH
Fl5IUlwJK32LQ4hbr5zW6i009nhJd1NHt9e/sQSCsuTnb2L5xWtMrPNBuPWy6X9q
1tjh6aXlPcU9fqYU2nbgqORTtCO5QvbikJgSxJLiQg0CUD+t+yG6n7O976qXsPum
N01cb1n2ef3DZeqvvptBIuqkReCVOr5sr9s9cAdd5wz8BzowbpfhKt7NBM7aA8J+
F4w1Q3OKt5EcVLfGYKgn6r4JxnV9F00WCci4uUpEuU6RrCsP74qJ75GhSQdcACtc
LMkO5+QYJvROTXaZrD+7H50nscUm6K8kWCe+1bSiRjGgSQA4wYezQB9dOSx+PAyk
99zh5kQdjZePVE7w+aAB8ADqD8eHdwkj1ZVIU/rg+xmbz5EwFSxedxC+wMygNy9X
tFnFeyOfurqBuZbBahEofrjgzs7k4QbcvargxEVSNqJfmO32FrLnQwCq4R2Z3bSM
Uunn42nT6KPWx0bVV7hZ/9KWZ9m6FHYJ+WWtKE46e/5LTM1xpCU3qFiqQ/tpmXME
HtH1Vf3ZX+JRlspyzosCNiDqLGqsADEJ8APtT51nnmzd4vxcRXnC5ZIz0HIC4UEl
rhPzQyeYZHzni3JN70sPsmqCFz5Dnic5PXf+NvTnX2B4o6oJXKpf9w1HOMwhbY60
nHOA5iUZj5BWgtu1yM2soo4sZN7rcZjp5X7OxoLuqO8WUHwwSIpb70FRecgYM9K2
pRkaUujFyB+mWjz3RAqezmA53T1bwts5LfQjq4BStdfijz2BbRnO2tG1qN+lOQBd
RP5PKR9M5AmTVvfjLRqRhMQHYPHxaAznSVvfNnYA8o1a6FGKbhC49I63blNRgpDd
9z/U/DSZlg8d5BCco2Zzl1eLURbI6im282/0jx9YyjVKGvPpvy062stW6Iqr2nYV
4Elu6R9EV+9jdmKenbRRrWud9/VDjGFKjHFmESa1WsGYbU5gOkJUHv3QKTeQj90t
+GoE9Su8vtm+maj2rwgo2mNVzrIabtJ9TVcNJMNXAL82OCHigfEpwtWDQDn1RDQX
kkXHFBV+CB3HilZm5gEZG5fCag8sj2fb1qA8Y0wgirSlEgP3v8vUzhiPvAsK8qbm
8EMTigXREjUxy1xi4MZUzD2YCGms6lX+ayoNwqB0YoLeLTldFkMRCelLMbCvMeOl
Eh6pikif0iacW81FMEpQozHrNDgFaqQQRlFblH5+3lU41ahczIa9OYTgbcMJjbGR
Hj9jDsbF38Veu/iALi0iPhwV69wanjyExw1zJizMDRsq1zM+V278jJ8/5VQ/lkPG
XuX022ZYaP9N+EBo3c2AFYcbdnxgjdKMYv6to/P5FMnxetOH5Df7NQDyYAtI+ids
pmmL+w1YWGiKBnXoYe2wTAbdTYSf8Z1gHZrcCqT/bThXo2CaxP9FeqZWVK7hMv0s
lhFZPqJl2b7XgtDewCamH9w0PVc++OwcpFGFMo9jkiHeDI1+cIPw0PNRJQHDNLjo
fhEMZxmGPZStv/1ZAWBqtLLDG+dfriFwFHZAQ4c1mnzo1Dh+ZQTz/MZHd2Y/s56S
GqQCzoVMzyKRkWh9ckkc9a16ZvDKcGcxpA2j5eW6CMkKun8Np4yKe4OzlX3F3IAX
tKUnY0RdClTfhIZUgX5EQ6hQ1qzAbMWKpi7n6mHOzGnSt0ERyK2k0MFZvjqSjZzQ
inVPEY1a007AogjRRq4NQYXzGXW7rAdvkjTDzguda0V459OipwN2Ep/YJ3CEFniV
7cADq5NJsWsiRyfnNDHTb7QCfcgnpb7Iik9nIMmeE2md1B4EQUqK+hzSXjttjVSM
hW4x5sm35sCXNNSmLh/orCBuVvJ0edX5zvS0dsIOfSsuB8f/68F6waFStYuMuzmV
YN/ftc83Vr8RZB/BqLSk//sZ10XC9RoIo3dQoZowOppgLAzar/kkBD9wPeZ0OefC
jN7ZXFvAfaZhVoF1hTnJcrBbGVy5xIjtKVJZY43RXktGULrz0ynho81WcITFmFAP
r1gJPGgLxVkj1i5AIGoaL5uwEh0iN0pJmdb4Yav/IyhJUAGC6sDMT80s5Cexwu/N
L6HUUNNEkORFtz3XTYjVHjq6dlkdnbKad02keRhPPy7aoVISLSURdSbfLXCfn3aH
KB9hi6jypmhR+n5j4BgTo/NTWUdDVmJ+ztp90U+sgEjc4cPuzzS7ORMHR8V2v0on
6i1cL6ucibGorbRoBsH3J4avd35SsX4RV5WzJkRxQLmacLPVPdsNLejX6Ci2L2k3
Xr3ULLrZoFwTC9zSxpUQ/QraHiS4kOFeSdE8Upx9ySFwF2Lz/8YQS9fafxm+UCNl
FCk6z/G0n0hAldagOj8eibQOadGQSV3R2BleFUo1kCeg0FAu6XFi5VVzKrY/NRzF
fSt8u3rI+AMfEpJSH8vhTHajCA63ChHXxStgDt/BOtvgkmxTTZ8IrAf7xwHHd9WK
zl5+z+VtKsycI0JdXDLl/B8CuN+9FawGpXmAWwJiAyUOyn6zc/1h9g3vXVLPnCpd
KQ7SrvXlcV/KbA3ku7S5/SKo6Nsf5FCtru1pKpSfj7OQ6jIlDcb0KDRigFtv/pYG
KQTCuVjh/SjBvODemIhtkStfBKDJLYjoVmLUqenTZxbYlKATVKlUbfpH+g+US1Fy
5TO0R3xtbzpyQWKQFojkGcpCrIbNmrirtB7rFwCKgbvySuGlzPt7LL3r6n6Tm3gZ
2F75bXTh4o9KhscdRbUilqyF9RdyS0g7gMYV8/UPC1HDfE4aIsKoXdeE4mnI27Qe
986bF0pn2EEJOzguBifEn1qHtMTWn1IhKJJYzdXCHjTpPN1UKzbd8QyKqkNlRxBw
SonkB0oIXsRYl5xInTJfSFiF8Y+izpCZJbF4CNs75l4UX2ojmRGuAVqmh/bmLUoT
DHegz2+gdu0Sk/r1VvQdHPRGi98y1XChn9goTAVqLFZvTwDqEN04ahwa482fapIp
Ot+FtbaSLPgvfebOhBNrKxt0jCQW50blDLbSMtpTQ8brBcDzdyToiRk2n6lYWziL
t8XIoENRnFSj3Ep0KhHTXe0C1/1sfSQrm2QLUcNvq+Wbl8BUxp0C9qBVBH54v6dM
IxFphpDvZuwMWiqhJoBKO+9as6xow81s+wt2ZuQdh6zyQLDdeKCxbOperfeIy2DC
JlVccMQPn5tBi5GocPbJ/1J7lnR3LLcFsLoekTZwa8i3YDNEU8hDOFrItBTWEteQ
7EfslPofuqz8X3E11Yok4Y1aLovL+roktq3noE0QRPRjOcAnv26NxkyMdyEc8Z+H
k2rftvDfRLKo+ag98pdxpW7MWHD20GV1Z0fLmlwAbgwq/W1B68xCpLjcOb+ouvza
CykUBi4qesIMmWxBNb+Ilby3cmRE6Jsj1w5YI2MJps5OYnikAVadVELJrKLm5JxI
Q42aEmLV4w1ilyWhzHgn5iYdQLZgWfiXB+3zu/uGi1oPdwAY7m7HRKxZDeredDsz
hesbngi98f9sfEKN70HiF4RPCDn7DklEsk42kIfqWj/yS52WytBq3YrtRreBWxU3
igFJgi76Auf9F0MEYQO2TKtnZyAiXcPETJq98npFN0z/7oOuBZ/7ElOFlldWSBHY
7tUd6E+JGT76D8SLA4wHKzG8ex5MgHExqNWB42jzGkCQCQp0Us+Law7xOIIE+Tp8
p6HpPi9Zs1xBxWOEPqyb4C7D4Y9CSCFaTPazLp46oyk8J2E7G9bJ6H9sIQK2Yl2J
xJsoyeGm0gGdCV/gJA01C9JYQPyOz62ovFNYmTHt/wh3W90b0JWgZPQc8etwXJd3
Mrz5Vdkx+i3O2rlSz8cXfbA7AUK4QYsiKCSt2tMb8FAhBV1JwyyCjNuttVfp3azb
SIWca52cA5++mgq+SdYHp1+M1MKurRfAWHenwzYgI50Hq1k/eVpOvj8AwGbZhci7
EHOguBSvEG+ACp0XOCXaSwPVv1CQrNWqnCy3iviZ2DIhTjLJr7Zu8SVmb1KtskGI
IvwHw1oxcyjKnOBNxfLLGZ5+zHKbB5p7aO3uHzAKg/sr+Ko/tJfdCZw6a4ygY4tb
fAr9kB4RSLmE/3bN399E6f3pwN75eU6r2qGXFEadZpIFGK3fRv4SFNmNZsm0HRKp
SXv0hDYJkEX9qPDSEIKTZW8ZnT+hjBSyJI24woe2hIfC4o5IId14f99xLm+czBTZ
tTN1hGWHhNTwYufyauGQekeiBsiK4YMWxbQZR10VmwbJuGbYXuUsjMB0QOxkjxMm
/MQI6QxRVdpbkCkiVDOF3Y44RydpgmnruwMP1FTMFFbaw6jNYluQV1xNpf90qyoA
7SQQUa2aRhN3IVqeygJUmeATKOcnHzGzVK3DbHxtSsKnCOwzs0BiqcWEPUOM9XBj
p6BII/5g6i3uGK6pYMGs9A35Y0TFwdFr/g8iaM6tbK6G1905QPKrN0vQ86uLc18f
xJ4QdIkZJ9p254HOrPhHvZJBqKe0LcTeSOUZVEJ+eNxxu4+utmrjazSbMap7lppD
gwkJy0EZU6hF9FpV3fwzYJS4R/E49BXe12cu1XULELB80Xy6i1BnNnO+wRLOcWlA
Q5UFJJS7KhIPAv5yq4abjOPJKQHGXo9uzD4P1HwL9dnLr+/ECHZAd+C87XqSqkuJ
pLTb3OMujPE3wWT4Z/3ttC4ZsbD3ZAvxAM9TSIfVSa5mDBHx9JBGqyB1bzBCPeBo
gTnLAvq/tUbSAhA2jpB+kDAp/fey8/aljLMDgo7kngRNuQhW6eW4TlIuo2IRYLEW
mDhU0zdYORGn8cr/9eBa0rDjreVVyeOcjFViCs1Ruu6eW9LjkEA8CjM7wXRJVRb3
AdF+5PO6/4YlgMOQUccBgBUXyD4vlaRq+ibbubOB/4etlgtWOAcM0/PGCYl9azOI
3VVZ8Sjhu2qSCqpEG98o3WKupIQ0mNjI8hGm/JtudbuX6BSAXjxxJpeRZs/RQpe6
3Tf2Inbu9h0nNb+W/wjm2Ezw0DQ4BAKgmmQA7VYtueKEy0XX+Iz+KSbzB+tqqj7x
2fKtcYmbgsTjwhR+ELi4yFVitTgFD8cSTmcUaI4pTukhgK9iTTJ8QcNrI7ksgcmI
AjXE3rVDaK3BBEJfb0eluMHOGDrmJhVDweIb/01VbKp/YWnRcJdm/qKRNSi8oO2g
dTCJgjqS5gTu/dm0DrJAB9z10VO55hvuMG3mUs2Zbjg716lGcJCrAfSe5w7+PYMm
chF2IlvIkbKqC6DpZEdC62M0IQT3MnS+XDgPwJpogGORl89cDUDj1v/2fA3B3F/d
WEXEgc2szEIV5IdkvIgZLaU7BpkaFv2MiI3W4S3PuqOgvg7rN0S7O7BewA2KEbjw
RTYGuQtn+nKzWfQoGjM7O7s/sVuIhaBh9wQojMEHlPA0ugc+zIQiEm3ZvL31XDqp
MC+w2ri8veCiU1tlmnXBwM8T6b1HPLSoWevuHI+qu/fWlsILWJ08+h+XhHU27xMa
p3p1UtP5yOT/y8tfAKJpK1FoRS8WnEqapAOK3+v29QRD2Orl/IBwRciisjMEDxHt
Q93V7NYhhjfXD2MjVBX5UMEQDvEErOGmMbKc1suhCxUOjEq+PgYSIbfAjgSqMYD8
XAtm7B2eYc4joMTtSUH09y5DTODOdjM8imhTsFow6t9vH0Pmk26iSFx0zyvyaiRd
Dvc3kRnlgvmVo3Ulpad7FfQV7nwcuA+a/opSuzKOHEfhxPomxMsV34y46ZzwfdNd
T+p+TyJ+GGtuvpNWgT47G6rKHGNim9V9UTDUk7OfDoouQUJr30ubK476S/SVKz5L
j5EkIxZdvQiiKwWIvvj2iCnPlRYFaVDQbYdkMWZYn3uPtI4dPqXJhmTImpl6ElG1
WVlk5xmvtL0DM+7sdav4RaUSuLu2JVWjjFaWKNlJZp4BoVrRxLixRFdPslApKDki
my9ULDSupeQ4cm7ezKCJ4oZQqoLTwBUvzFGIRKX0wE9jJkXjYaursBkUoejDrkuZ
fXNmXU0fQGSf1u4O7o9X15CEI6/hp7fngo5dTqDAtUkBAc4QDaVSwIs+cKkyF4jj
PsjenE4wLpQ/krnxeNoxwiv6QbFwP0QPweHhq3DXSP5zO+NuEMJQJsoAQqnmnPiU
LB/IITA4eSlRIISn10/2lExM8HsYuB8xyx2EYwtSwTeOnfkSaIRI8AeOLKsHaBRD
qqpNXy60LKTGYve7qHrUAJWSV1MFP3PyxGIPoxp6oTuZQGs7welu6kiWIMTt6xF1
oCczw2OO8nPFOJ+CTuG6JUpncvgMEsS5vRjK1049baUWc6WcIJwt+ydco9ik+Lgz
w96irOqyT2Ec+4O8Rq4lHQoZG+qRoYuxvyDkyl4vP+wA35y/OL5w1f8DxhLOzz/w
kPtBa+5f45E50M0xtSPtU74tYtEorBAV3sltUaJNmAu95zJODUBl2l2Rp8gkQm1V
+Hwsn/K9tXwpFdk7tCZM09CExbNqArju0KWNHRyrBzTOzBtc6nuXiybP7GZUZ9vL
1YMmevAPBJ/WCtZv+/E4h04xRHx7KQ/mtsNli4eN270m3bFcq1oI5gCoLX7uJuhv
tzZP9G7SchY+4UlxMUCV7RYzrokeu4P/92BrztMe8PRhXoAoJfdwJRWEELFL4fm+
85FIg1aAtFAvtqpi7sBzo0mnl/Gb9ItbvIDSE3Xr8h74h8bdjavCUe41z33Efqfo
+fbvtDK4haDc1ByiJjLJekl2TzJVRQQ/PKIFqO2KUoLUWCNj+Mldl/X3UaC5g0oK
oYh27BVYC8mTZjmWgafsLqFLBoH3KWB2jJNOds16dbd+jPW7ac5qDWD8lIFwEx8W
4GkVknzM26l4YDf5W0D9aFwGlVLf9fMutnNcO4k+cOmR1cFy3hR0fgy65Vb/ueqy
jNXkMbK31oSyTWC5a2RGy0qmeVa3CFX1HucK63VeVFaiSJ8NQ0Zonc2XpXf1Wu3w
4sMZpRsVE/v5Gb3bnRlA9VqOAQu8InuuZh6P61oztw7Sp97VbaKTgbP031K8sXsd
iBEdiN6RLDbR39pz10iI1xiHAUccJP5+ZdrCO5XZutDNfrB/4YYiXyXjndRvv18A
JDuESwhM2dRp3h53WOsDtZYbRK7PDTv/+ftiCPbDVBbbqlTZHCp8HCoPzBTfNlWw
UwrlCsa2OvzhPx7KQgGe9rgvFGQnrVi6Hx3RG57glLcHA7CKZsX7HcMUP2sh3C5N
XwFI+29oFD9nKA/q+4O83HOzzkLUS4MwRuifl5s+4d2zLLmZiJrk5cJq6IIoVS9P
3FGAjmc8Md+oKdQQvrlvEaXeoG7w+xK8KSZZV9HhSoExKYVZIlLAw2rfiYj2HqEH
+NGskXbUTGpOSLz1VOJrxdQX0yizxVLFAUv2m4kH+Ow9y111eYJ+T4h2drfn/wUs
413K8IwN/sTb+EFI+8HHYhltxOwA/hEEKpuMSdBs1oybIVtH3FSvgl57N5FKjXlH
n9GEcyGfb/UieetUj60ZvQYJXXTTwXKtcsw++HGhA8i1/3FEhUnlISNms5/v8UBp
7LKvhzVSQeoliKXHBAirSUbzDfbHAhfuhZYGFL0EFjBvpz68/wlnIvDSnLe0kkuD
3QTZiT5gSEn9HblIqo+P3sZ5DXpZ3pkef7aSi3UdHPCzp+AjWiUNTAHeIIOwyhPD
W2oS9aarDwfIi7wpWk9XLjJ5skH2kbLlN3wwrmfZN0PrX4pNw7equ4BcSKSkLrmk
BADKteaobEXfj0RffdaDWu0DvIHq8NmGgLHsTH7YIxRBjTp6hWXnNEhFl6Ar4day
+wbZZZIyVj7kRSXC8zOpKbi6FrMJKipRie9Z5Am0Z2WBlo9EvK+Olsi/GcGXHnzS
HzPBzHoe5E80jYZg//fgph0IOWXY3BZsQgRfhJDkN6FSSw8ndxrmNXtkbbsiCQS8
Cks4ohoV9aD1gy3j72tChEiT3KXzak4IvbIfvRhlMkmSEG+8IL7YXTyPH19W64xW
rU2OvE2Zqe2Vr4Fvm0WT9hxBQbpL9rdUvzbKmGpZ4RVtC9nklHH91WXt9/Z69d1n
hQx1impIX4PIJEI+O5cDBntUjSplHPW5jvfz/IARC78QSXX4iGjCxnHIM275Lz4k
gZ6Utyu8s0TeTj3gWASp25szn+hBq6vZeRGdvYZkup/VhogrUgYT/kEcL882izOr
OLONB1X1wvps/2UL2Nr0Anbc1GmJqxxi9OXDDW6ZByO5M+e18V/00DfhnY9A2rXV
g+BXC7IykIt2rGBgaiEutvNIDbn7IGjZzGStnjR/VXQmZKgrOLRGb9IdmhC3c8za
malFEBhF7gY0JZiLXCZlhBpMI7cxrPI94Vh01i7zhl7J2elXSyG80fkI8TVHT6Pi
lNVKPD9ESe7nh6SunKBHTPME3eViutJ1jWrPdiVevcDcKmYMwRAJprvAITgI2GMS
7/NtGP0uI/nRjiLBNBvHEeZfktTIx418fE/JZ4G0YLyQCPgESrOZoROqYGU7dM76
Vch4gl3K/PFgu7pabAiREQFFS6ZuZdCjhnUlaL4XnXPTaA73ivpgJTfp4Ucb+Fgz
SaVpciRHIEek6PPgiscT7RgD8RHNvbHAi9GjkAGA7SN8c7uasHLeRaS5ujmX/7xm
/duJ8huWQySg7ywNlbAwCL33HfTLgv2WVCrgQD+svORSR85BqE8cXaHTsOdjrmWo
E6NzdtgGm2T0DzFmYM3Km1XwUzjf0T+GRue5/TAR+BK6OC8qFviOkYl3Xf4+DbQC
J861Urw6zy4jAcXKIjXOuCpUvbOPZ5K0lB/vNPko4J66jC4TyPVF8Fxql08Ojwjp
tcwYlK82m8QEIl/3ZTptD1G0iQpjUkY6QB3obOFiW4QoBNNaRqz4JK+lf4jqODjD
VoMlv4T+Xfmcj3qn51RZ0toctaEdRAVHrVja0HoOlX4XDBFTMuBj8nfulyrMOMOa
6yb9Kbawc3T1CCU5rajL5GAkaQn8UeIeaIvkuZTDrnewq6foWWkablf4u6uV37vy
rExxVz/GxQ1/0VpuVxSLm967kmWyYwnJW9Wlz/8dP77qKAPP+i+GwmCX71TJB0HY
YgtuMfv7APZbrdT/0XLLey/yfUHepUeQOAzl7sjBBNfGuEwX4ANLw0rdnVzjwwf3
LWVY00aqGTkdYQbyZ/a/aoNOJLS/8XqaBvc5zb+OqQB5+NkapeJLCdCtmE+LHukM
f5hbtJC5c8lHlT1sp8yDA4ivPY3zNB1WmEBxOrufdZgqaJ8JcNcd11GWmEFkzY3y
zPV5d6J0i2UPVOeOPko9RC0qglT/wiyBbKMZ6vxNs8iUcYEI8S+Nt7kRhLJSFuK1
NKWAeWcgZpVEs6yX7rBS1c/xSOzbjzAi2z+kKBi1IYXKD1DqO52gsec4puCYCwY1
Ce8V5uecTMOpx+kHC2/HT7xDkayPB1QovwYXIrus7xi5IpSl5wcbNENTydxNgxhm
VrIVr/QUzQVlaAWTY9vZV4mYd697V7XyRLAhGPbnCC4+FEI5nkSC8s8HqvCJEbSS
Ucie03danElaaIIbUcyfIBWp8lW4yvtIXRZcR4kPki41BU+8FT+BZ/U9psi3SwnM
+MIZh9pZ3uYup6cIjGTxhORx3ljWorqUCnVJVxs/6wGHkC5zqE0TUedcFrxAKGdf
/IsqAGaWXOsWDAB3aOOzHMBscQiz6pUZyy5vidN243gDjHIeCS0PQlCEFi61N+Ty
4j1MbLGZ02KFfgBl2eL9BsxiAXosf/liZAufEkoeOj9TquPyB7SagduD/LAhSuFY
csxPK3bALluWxaXVBUjIq/ZFMp08r6cEI0gTcCl9Kz2lzfQIau7cPl+RneRZZaHX
KAlLR2Fe8HbX/4nmB6NMBHLH6zyqng8so/A94fH4/xIdXQVQkTH8BsnyMWw/r+aP
XxuPXhkBDbfkVFPq1e6o4QNGCGEYCPcUPoPbY63o4IroVxxpDZRw9+DwvuVxTHdA
orThFLN2KTPLieCxsyYp29m2iakGMfmToJjnOhvKLX670fgUAWQG+xp6155SMpFf
g1fNjULcampy3GMDhUmvvRICpZwOikOYWgLoWWV2wy0uHJt9qhRNWNjqr76PXasq
XznUHzzLwiggqqv2JDKWD1fyMrGWeNj/A4mQvvExtv1C7Cry3LcldjiYcEJ+2+zH
9fHFo3gpfJMtH0ELA9fQ9gqvZmxNb1LxEVEnUwo0GWbuo1yDeu6bEoQ84CrnLB8x
Cv9tsiM4z8FXdL8gjCWt4mjtFH+pkK7n4Dvn35AstfUoTmwxDG9DYUcC9CSfKSPq
Iz61D2wu8dAN+VvUPqAFlBcAh9NFZ+q5yZv1fyuxDHwwflGWQrYeDKbCRxbYI2eB
DKrXY/aazXgevZyIzp/EkAKwmGSxouCAGTKWLNnfJ82eTN73hRNbgRzU71chZa+z
JZXtWkqAyut3f3tY2HnEC6+M3XhQGUkSgkFA1hL+ao0YgAomTkO0RlW/hLN/bIyb
kug0iQxqiN31H8s7xrc66Drp+lzsWfLwxItemrNki9P58N69K5EEfzmAaFfeMYZj
cdAAw4d+MrXKwhHNq1cup8aRwbLlQBhtP3UODVcxh3QAf59n0teLDKs+bWyj2bWY
sYjwNvtT7VS69tlQaPgGGT02oty2RpiA7bmswfh1B1qC4jVzqKgyV6hwRxS9/uJz
DjuI4ul9122vxmRCeA/b4nvx19PAqE4urPnfCrP8kUJnrTW3xpfWrcPReCmKoOQq
FYtBAHCBDvx0B/aN/gesqzh3BDGDY+fEZ+edS6iDpY6A7VqKfLLh44KxQlzJPYLr
fqGKsWgVahChvfLovSOE9BLXQhJXrdyP43eMILunqmYNrWZK9JCs5gu2lk14JEiR
II1BKYGBGlpgeBEczhyC+Bp10VRo/PTsmnQCym8a6s8yhk5uP2HB222YnH9D4xlS
TX4qjmOkwlB13fD3atxJcMUpvbga5FGLY2lY6fumQQ4b3QNVNcW5YhIf6x8aNVhs
GmiErQRdb+K74QQ+ZUT8xW+b4F+rAWbwIfqodjz+ZNhK7MywoznhV3Jig+cUDRu2
yptmaw5bUKk6T7hI5YcbmMTisXzQ5u8CRHclmsW3nntIFznvOToIagoGvgZcCKY9
TW0Wp9M8YHtqTp+JGfcrWfzOlHJEl1C2NBAwPTBNVX+wQK7rk0Gs8jefa7MlL0FI
674IIDVWtr0NSr4nHAFN8BaCxrwvn4xT0GfrtrCXdKfwNTqAffmKMqvRGAOnIkqB
WJfpgAsmUEN0KZCsQwi5RMRG1CWuDysU/9HbJ00QUu/wnzMGeXiP4+iSRFaF+7p5
YxKxS+hEFVnibgUJ2Br8oMXVLU+aAYJwJJd/hCL+0sS0Tt7CiI6D4LTjIs9PkJve
NdXhh2/S29N2r+vJFaMqMj2ypi5PSqVNlc6EI0t7oMKLPD1XltHrowQG+5GPCUJg
xUXYydkMcDwgqqXvY8HkwyEnuolYrLv/0QgdMSNrjiioLugq5tmXb6dYF50yc+E2
ujhxypsmj/pJMqe28NVA5SnIKNrnEGKnck+nPK+6prg=
`protect END_PROTECTED
