`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3iFSUNFOzrP497qB5eDI+HP6wY5u2e1CZQHJQo3MwU1zWdT+7wpA1BIdodRTKLO9
MhhpY0ydNp1ZjdqLhsiv0rKZsu5ae6YOhk0JxHfUHR6togpBL0Pzcg7uWx+6KGEX
gcaoqwHHLdXOtKkZAp4hzBcpus6UYpsYJFWX9ZIlZ30KkOUA32rTlrW2C8PyMECd
CuwvFEk5oyo+ooulITHvONAr+XMxjp6q2U3Byz67oFLlAosoOZabL6TA9AhEpvXV
1TA31f+aLCN8jEKGFQ+ACgZJ0toO7QU9r27pcZJj5iBR9QjIOMyLLuAWPAMqz9Xy
mQB6fXCBzCN+kaA6PSKU3lcSVeZrKPMIr6301TKlk1nmpjzO+KtM49aihbtEGE0O
YTB7hMY1FNzX2g/S7/fH/H/8JokZ4kSH8hlzXB/cNvhGPrkbE7jcLC1J2Mhh7U+d
8UBUW6voYPeVXYk9m/fTsyAWueSc/F6JvLYm1NxzPzRA2+LZQp0WVxNbNKpUDdce
HaJ7gjn3te0qIkjn9jPOGfiE8+hOfDpvU9VcgIPFsw7GV5V7wOLs4kAv4cyeC3Yu
x82qz9FvfDHp3bkh4nCmsgsgm9Jg/SLmJtv/jYir6Rh/6hiZYjKVLA9o9XIKnGky
QnVr22Nzg4KZAuF8+jF21a+BhqXun+5Z/yDps34C5EWrOzDlYgCWpMorizeM3KOD
Z2WNKUxZ0F5RaQRTlGTQp/FCsPw9rDbWanEb8h30D0DNmXGAnhnqGl623M4VGMYy
Nz20XO2AGIQQ58E/8/9hPfIXQYhGmrmth+Z8X27f2JkJeuy4ifFwDgfkNxtyHJPb
ZXwqdAlh4apXq0jm02u0/i8e9/55utCPPD+PXppm0g7zYUqe2hyJQghZLcU31SRR
HDUJhfG11EmHHrPvdwfaC0khYsL2TEVLk6cJXJIRowKzKf6kF2oN/XGDvAKPYpx7
ulubeWuY0Ue/j/0loWrwL6cOWJ1Z2SAgorZa7ZWSj+b2RfIsEHZbMwflwke3XORW
7MFHS8lK8i9fOG6rDZm+kjyyt1TrGOY8v0WjU1iIvizI3FKeq1qyRXMKJWtd0nzD
rr+/y1Pvc5MbaaEEINxrmtKUk/TgWE1npSbHIsyUEkMlPL0GQieH3VBTaVeBgK/e
wzMUTdaBZqG0X3+DbCy2ntz4Kr2f/wzTmzjjrzZUIDYpMjXuf9G/TZAdaDDfo314
AEwleI03dyQN9BbYNJmp3uu9KAldgZEgNhzlAYb5WYJZ7zyj2nbkkHG5zSJMgaS1
kOJe8QpULZLkgLKip2XYfQ/CAT0f8P7U/3yP+eycKB3ViK/3jZRKQVS/aIodLpXM
yu45chzk2/j+XSrZQdKysKEculJcbW6R4Xh6uik2PPTrg+jakn5Eeu2Um8gafGIu
3fq4WA3eHistXJMyA4y+ZejUDtBdAgQgrdYrRlv2zMCKjKqftHbzEFEO0dUUXMkB
kUHDYwWtoWSTYGYj1B7AMZZvkHfgrFhnPQkdrtby1R9vUR2sQdozyK4OPe0Pcgxo
CwRG4dn7AHSyHb5DQg5RM6+SPIkiCafWlMVPePxxgX8Q9RcR4aSXk3N6gHBZMtXR
wqnil5GK+bNgPkN/yzla1KBn3b3/Yd2eK2rUEIgqK7Hy5YF4MHnCs13EDHrMOdzJ
jihPm5NKATdeJuoC5dVarvDuUYHCoMyu0APE4/q+rLJdF8A+98/icHy136lX86TY
BDz3km+6kSuaOCzKLC4pmrt2x8yJlMaIBkdRiegzAV0HHNotej1JZvTlx516QcEM
AK6Too3QeIj7c5UmEVsIPlnWX+uQWz4hZh9Z7TZNx25Ilgd5TMxqt/5vaKfdQ16H
Cd/boO/ZVWyxcAFv4NgSSAyy5HZsyBfK2vQ/vskDtzWD3YMA9TIvACO8jHQHdXiG
`protect END_PROTECTED
