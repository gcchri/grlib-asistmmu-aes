`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lI8tjlpKg6XlpjTKFZFNUaYrBx215erALy9GPgnmPOGL37Bo/+8S2GzXLk4rjBzt
tHk9ZYGew6BtTYEFpbYyo0AXEjjNuPLoIwoJNRKbSWIjVesiZUWh4aYspokGfctl
CtNDBi5RXfgAo7tBxpMjoues2/FTUEN1au/jdcxzwhrfnajp/6vbsIxRRGWaN1Ik
VKDvuLDP/F2ea53JBtGX3zMZE36QiwWR0UN/FlgSave2e30WMsdF6RaiIWNGJnmd
3C2rW9oKK+NvnO7WEh4brh/qOLQ3cZLOOWevfRqIqEj1F/Q30Rg7fcQAHH9HUjTU
OYY8ZwINyr/e+QviKc2+MFQbyZOfqOSoNFv8vUgM+g8gZWnx6eAIZ44PbbFolrwl
vZMsvU7Fv5UBT9ziALrTITijOb49omWSeZ0oDHl6AzWUcOVRbjcgXdKOhLQHPnaR
PBWn8ZirhQo6zIQLg2a93eC3quo43iWvo76Qa4BFfI5Gh//2ZvN8wTafvCNBDSMe
eQkk2oOHoBL8/RNqS2CJlzAbn0dypZRoGhvAzziuNK5/69KhCs3KG0Gew+4WrLFY
GsLEp4Ma38HxeEw/aLkifghViEgT9vtVrl8BmlKsn8QNMnYPAtxG1HHfgM7zgi/O
PjOpaC4So152A2S4L1Rs2jxqcw3lJc2q199NBZ8yAMjYfXvC9ntque/y2+8DTUG7
uQwX6KkdzUKX1BPp+vjHwRbiB2OsX7FMOPwaljAAv9znDI5ZYfx1X78NfauiCsfK
AnEjmA3I+MejoB7tJpP1XzBzrkfzhHuJZgle8hP/GvqLjUgj8LZbHFTvLMC5A0YT
hwsp3jpI3dQG24l6hSbb8V4oFzS6H1E5D9B+AYofHgmV0tEVb4/+7aCJxu4Opwtl
L+InMoaqm5iW8ZstikyozJpxmQbbF5lPl/YVS1ama/fuewqXGenZ4uAir2RNnHT0
589Le7OFOgFfQs6EzlkbI9ggxmC5DtCQm9yrN+AyPPp58dkJvTovGGjxThPRp2Ih
dKjFes43kRaYFZljt0YxgA==
`protect END_PROTECTED
