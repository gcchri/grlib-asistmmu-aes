`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8o+ouv0IQCNp0ZbHG5RfSgSaM8xrsBzwFf7t86BunEeroF0bmfpmS+76mXoJaa9n
ZQNI4ntylCLM3zEyoMh5V4ii4AL6ot/HFppAKqVQTLcw46kcpUqLjtscyvOgjQKs
3ROk+wQe5hp/iaKILXruXiNNpKABorbEVyD3GYwGpXTbjDFigprbxkAiERjvAU7z
RUkSXBg7ui///tc++MvbJJ+MUqr1AEZFC/ERiQs52uFftTYALpBNw6jxpYz38c4i
UY3aAfGEP0ymadgLVFVf9wNpg1NX6dZVT+mVrJi8npsIodkw1ty/AC6YkzCCHdst
l/ZN9iO27SUYNcVku5Qm6r4AY6unMTVS60GsMpZviH+mvFcTkL1/YdxKkBUv2E3H
h0WWxFxRJPYHJZnBCd1ffLr/xmr4cwqkWrzvKkywvHSYblFZY7H1qIB6AsvId4PY
ShIzUHcq+1177z7U4t2HR7H/wKQCVDloUsBPdn211sXC86cdwhYhHmXU658tjYz3
FScJVEKjftYdI4JImo10FEOQoT21Vydsq+N27tYxJB5s8Fi3O2Q42w4ISsmMxsz2
DpZj09FKIwHmF8Rt7pxnUMjWyKt44EYSH3f80/IU31ALiJA8Uvi4PZnf+mtXB1RK
2JL9v/LNPt8aTb0dOBVOKsUmHiWFLF4agnz/VDb+6C6knm5IAUUvfdx5bw4kgyrb
HNltDzvDAbTStN1DpTK+dA==
`protect END_PROTECTED
