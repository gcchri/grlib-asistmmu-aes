`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NKfDzsVaNCfDnlrcjYyiehpNjiWmT99lgSsfzTx3mGkT8v6oe2yTE//Q8jVUtDf3
PjKpYndOs6QrviYuPa6rZQWXY2BMV20U1XHlRYlUxOFQeW7fPqBGzw4JCmQrP0d2
kvIUNAFlQA5Tpsgywi50sUFwWn2njPmfcUvRP8QZZuXl/BwJ1tiU98FhZO4Ef2Ke
YJHwQZd1R7swpk2T2RCofYMeaS4qS7kjsxLXJmWg2tLX5Feqk+uWhLj4AiYreP18
KPWs5hO8yj7aoejDgDOQK5D3ClB5RuBNAf7eTnqAf/bGFCe1pOqtey/Sdn9+M580
7aGAJoPr5aoJ8dMCpIrghdm9F+wxBV6BbhFkphS45OnEtdLxBY71H3Wqw0Kb8RUa
3N+hD+AIjRfykyU2hgZtRtoHLbW5iYnwcqotFwSw5w0fL4XYz8bMBO6WJ5RZRafX
02bzQhiXXFU2W4tHue9om1utxADpIUDPa8tzOu/ukzY=
`protect END_PROTECTED
