`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KqiWXI5dx0GnzEFNehmxTGLCTB3YLVgatjTFKC7Nl22pVAfvRRAbLNlTw8RYm5A9
wHyJ7mQpZWDutjBJSbRwd2DrgULE1wwdAVsnGroCv9/8dileoIk7tJnJZbmWp4jL
/a7wAVg6zUi5TqsU8Et31RTGBmOdZsluYOnCH7W5fOotjo1Cp283mlchBz5mmyV4
L/v6SPxyGldc+/cx/jrI6h437D4EB9ERaxGdw0DDvKkpafutpBxpWEsvhIDk8cdB
7IIGi945pYf+f/mqj2zp5PMd+yjcZPmlmx7996Ja5fL9A9qOrMUhqNjYNBx7oMwF
dYIg0T9kgAo2R/rSAhXyfPEIWn5Ia+kyVIAzbfJIjvgYZDTi0GX0+peTY16nZKlz
Af2rHA0iXzE4SL37+lgT7hoaeUeMjbL5pFnqMJ5HtahL48IFfTIuvp5y+50akLKh
OmO0pONeaodcN1vQ0LLNrtsNALNNz0YYYskmZG/P+EOLdnKod6kgba3GbepBy1/W
TYIncQmZekTNkXacVqP3Fx/Kpnal5h/qYBSV9+lpd/0TaACmlUpOcBnrBEbz3Wv0
tHIrLXNf907wb/4fEapY0YIbiYwkIUHEF8L7Hy4OYwh1Yj5mBwh9XPCCs/i1z1hG
CUnIfIAZfB4Vg9+5yayYd+H3kQdGxfkdbTGiIECTwTIuAM/2pe58QOPGn+Z9rE7s
k9cmJvVYmF1vcSuKjBMlKL8g3NQKpLQkYDSscsJlslf8CRjXb+C0Ztekrn+qtZ/w
ZOGJkY5A1OIQy7bJM06Cn1mmPcWwmx+/bs/LFFmvoxxuNhnI5YXg5yaP75yp7QNS
J4glcTPd/fBK73QaUSJJyUMZ1R62iAFfMIsPlDdVkIPYTMD27eQw90XMLsuqDB+g
MRwWdJcywfubWMvYCkhk1pCw35MyPdwdj/tCBgFlesNr5qC5qSXkG5LTNGobjCP0
AEklsK9Uk/ifTtRgQwArRqlY3gcd/358DqqEBsz7bKOMjTJ8PnM5wNOpF8m/nF8X
YJ/NbT5RnUkfSoOrDqBbg8jSqhHi+6zP2KWFJbFRxzgb8HHe9Kit5C72De3XO12h
FTB4CZMBtRORxCiMh9358zTqvWFRXeIvmWH0CcK5tWcJjp/yeIEoq6X+URwO/Vvg
JNJZ1wNeoegPcU5HOHnnfWc59NGNyv1cmCX7FCbbgNtYXmYASQp/J++mLEb5aVoN
BXEdCyUODrt1c6Umnp6aZXH3zZjdhzvp/3LMg/1sT0VMh+2qUVZLvI2GTCtOZMZ+
bRpcmf/btaSGoLgxGLrZFgKCBBsvB/ob+j7rh1Pwg9XkHPSRMAWbd3d3Qz5T86cH
zkCg/9y1bpOmd3Pm8czkFlAiy6kfdHftedEyc/npqu6m9ZdF5A5uRoB71kTbSJ8Y
GH2zo13+oX1OkKBXGgUWOIDtCcORI0pJXUOPvhg4imPj5QvmbpUKN96i3tgLPWCk
4flFPL1t+rKuUlr38nCoREd2bNmLOE2zIiKFOncXeB/MZffvbBK/HI/pucFMotnE
yhxPbeeny4Gmudd9AP7CGxYHYPXmj5oXOJUxoQw4UpFA56RxQHuRmtYUVNVz77tU
Fxxsx6aX+6Ub81w1yH97K1kqhtS8nec/XbXXNvqGESsUkHfu0BAk22klUTmv6WhG
7sPuER0pZS+vkvO/i34n21EFrt2KWZTf92ffNSsoFj0SCfJvULxXRCh/ve2mBxZm
sP/smFYdToGNNQEXK0jPm2MvuOOyFEC25/sWjI9boF/x1EDahpt/bzecaswVhreN
bDCYW/cJnWr+ZatYNhBFqrJ2z/DBy1w1PdtwOO6LtrcKrwu0e8fxXgIW+G7bL/Eg
FzdSPfdPSBSwwjF7fezNUU+3O7FvBCtqIcQK4V6K59U=
`protect END_PROTECTED
