`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pLUmztnWIe2mVkOVrOvKO6aJ0K7b2ACGjcHkW2sl8hfv3gDBPVlQzCGAqIVForYh
NIOllBsczci/5coCMJeDb1O110PuI966gG3mWyO/D7HxARMKCuYH2Is7hNCa5dq8
2KH9w6HKU3tEQXX6wIp8gCRyGKGcsQENExe8rD3fzYY0gLYeQrJp3PIocrJrfq5P
OUiKm5SF8AFCfnYVrKm548G7ohAHPRveXTffVapq/SM7+PxSdoCyNTLGspHN57ms
jhZka0fJ1JzsA4ZxPA9PL544BZEchkYAUJkB2u9odkoN2GObKyyaayfDyo19qEVl
eyNuC6e5/kG7XeOcexOmXh5nU3BdDyf1YI5EtcyS/ex9pz7J88Itv5A7xEceXovm
jlUNi/3kH+uCGdU6hy+LRqhy7QpOR9sdLpeDwZPfZa6IEkXoLsI9L/2qqnzwZ6Va
IjNshFn6JFpvz7/iBcakqopvsv+z1LD9xua/2S9AE6B+zWCLl7taheT3r74y4wYS
`protect END_PROTECTED
