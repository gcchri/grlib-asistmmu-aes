`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tidIxmVGV1IbsPtI+wHFG/aMWPG5rg//9Vd4Ku0OrCUYXb7d97K20nupOq8Ev1J4
N27gZY0sBVe32qb11X3zrDzStKhUGCujed8jofMvuXa+BVLASTN9fuMW+Be1QNbX
rXkWmxBOeS1q9ByT9ELDQlVpZOe2zfkCHw3or7c2SJLog6dctlkc81Pza8EhqERW
kz9jqJXFJdFCnXu6zaGxqgh4iQkdQ48H/l3iXik+jgP+KZg6davU1A30rZ8XTGug
UDLP6Y28bJYZrc1FR2eReBSVL7zALTcJefo04OQcrXtrCXwpgdGDc7qUbzzPLs3z
VEtmiE8yVYzIKsYMzpYMQ8rPFyQS0dv5j5fDiCi+sWkPo/v0DJ4LpS5US2xTUSNy
eh74okffcdEjpGmiLiVvTlJWiXSIBRdBnsanpQiZdcSG4yKYSwYS2q6b52jehz5A
l02VwfAt/+ITNerrZA41NA==
`protect END_PROTECTED
