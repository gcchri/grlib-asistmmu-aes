`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JI4yEOE5tLXDStUZOTDzFJWFUbGu63JgbwWfYlMVOtjUIy2tanVfBwGClFR0AaVi
jAq8s6Z0VoncpX6SMt2t33tuuTG02G5pa7kQh31WtoJD5CnLM+e6s4vwYV0N7rlT
C8PodeOHd2TQ2z0tH/g8joL9xVM0CDn2uoj5JWwHqTT6eqSDTNUV/dxmTj1nuT2G
QcOtZP0kc4u9RduyQo3oQ8894eKl2gg4mVTOfIIUT+oQX6qMQXsWJFbFgpMOnED5
w3WvYm5eS13bo/C3XQ3Bvi4Xu1MPYQcKyMjwVuKeD5VkjsyRFWbWxq2EolK7kDpo
SKkKojYd5t3OGTJFU8U8YLEA9m2egFpftRgb1d4U92bDm/Z+Cz0pNqxw0aejzKtv
oHKe+hYYloj6ZUpmHq3O0e4TdDn/C/4qPMxm3v7nCmwyEdmmDRTFbPMmvsoskMDy
ItLzmH7Dfybcsshfo4nDL8jbr5EJo63V4tihGn0Xny/VcYe1vYMPIR8Okxlk/ws2
Avx8EjVAi5bOlxFq4LB+5DhroHQFQzmKU5LdqKc5QUGWXITxtw04Y33HdHqAnvxK
pzMJM5nuooaCiB3Q7ugO8k1poAoelli36mKN5EFSAIKDaiorg+aYuRhX5J3lWdJF
1d3nRHC4fHQu5U0AslYP5orZUkqR1ZBGWDGsc2yR7rJsd9N7IdlM9GjSkrVYWwp0
BL36OaBvqVG4LRdPcPXO0VYXSSQt4FV0vLG8jI15DHSVSuGkDDpDxtvH6OJUfle1
ZSHLNLk6tzSEKtIYjEbyYHl+RpFAafGa/5YYhkqo304B/RlTM/j2hrMNHQwia6aZ
e4UUCWuYKJvGeMTHhZMIuSsAhvLvMBF5zR5KoLSP0s0+hYs5GE5hREyM6+/r/Z3U
CWN2PA4OClIPMX4YaQr89KZE3Pyam5QA7mJ80NxRCCfV+KkJ+RAL9w9m8OW9fOum
wnvDn/XsMVOIovWflVFTYD9sIO4YdNSildIfUetQCXFUL9CsmUxzx/gaa5QRI/Yu
wOMOHC8afXKktOiF1Cv4r8yWh1BxEBycJKyjRfkhoqMPo6yN1ilDUa7SA6SAY/CK
1DwGwmTN20ItBcA5UaOTS4GVBDyFxDIDGGh0y26W+wawfUudeXlZLLSG2Z0tFAKa
VLa3Vflp/FHhN+EN+kjb3jd1ujK7dcnOw9lQS8e+LCAgkK+xOKkiXGzlia0uAgF/
UvGidWsz5B37Gknm/s/xYJxgvZ5HCJsJGIRuErQQR4Txjh0nNPvwhP7jN0UdytN2
+f6PxZd/OI0mrSohxfAElTyLxKx+A++IxZz35ai3pcwltY1vPCEI1bXHtmMe5Ha5
No3YPjhOiWKU3nwVTvQyOo+afLpkxjsrHnns4PknJv+6RR8dUxLaYZgRWOGs6kkS
rDfqzOfAGmUdKXghF/228wriyMCOpZgdoKy8anNbW8LWTKSnbLe9QITTXzhAEO+p
UXvfC235ket4VApTGfU2Gyb7lppRahn03cU3HTXyN6xAGzPvyguOyoJFGKjS7vIu
9W8jGneeeyQwZIun2ocJrDhgEcBluYa4s98pbvkEr7fJH2Meq8gqT39SiL9gHtaW
gQbmVD6V5V4Eb0R0UOilEyhJUaGVUFfPziwlfmuM3b3EV7TREgY6KgrcfVQ7kL3P
OHVf7wJHQ/Rqkp4TVIt4sbb/mFFjd/KUaBFVYZVB/Pnrwx9CigG9rPLl8L2lB46W
t0SrZsfjUqu+HzqSSicjPvSRU7LXcCj/bKf8XcVCGOFr32whjK4lysgy81dLNSzx
4GE/WGsR5YoQEQk+U62NevoEm+rZe+IJJmB1h+FCgWOTdcgIF8EV3NEcyun+5JQ4
IF4xH790fe2aYeu0IHMRnyjgUSoy33OoO3fPnP+CIvCjp1eEBASSq3rmsCLjAw58
qDz3ezgDNshtAk8b8m6AtChOjDPISU2sgha6Ql/4i+V5oDkTgFvIhkoIdvAISdQg
wLtCkU7A2VDof5Lps2BmJcFzRddEIOksKu87iR3hNdr3YN1Fs4v85Lbmcy3PM2Ut
9+DV0sqV/2KGJMZx7xevRw==
`protect END_PROTECTED
