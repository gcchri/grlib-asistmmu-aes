`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1bNnjoPuMTCV6Zn1kDwwXz7oJnAdlyPwSt6w0pBZ7aaeN0xYKdkKcU+PaRNq0epC
D6+OQd6oPAUjg8dee2+JiW9hNrcVfj1m7EyhU/oEXBzrTq6u/kciWuwpvF7Qp0wn
n36qto3In4W/98N51FNBxLpI7Pd7m4JbUZVFh5zDhrCJLtZcjKERNG/kOawkdQwf
5Z6POZ5FvmBMgld1NtiRobNo9HEGMz7jHCyrgFlHmcEdEYtRb2POgqtkLGz48ZGr
HXtCWQlDNAZsaT905YH8qQK4kOryQqYWkntHc0J4Un3BUwRrKnm9qJnwpoXlDogT
t3GTQ2eda5Rm2bZ0EkLQDzE0QevAyrXYzcK1zYxbHQAbsHqveQEplUAQD+URRjgM
`protect END_PROTECTED
