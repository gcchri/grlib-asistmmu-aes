`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q/U4f7W9KoO8SdDeLNojgYWWdYIwEueeN9+l4OlAtHHW7c8O7KqfjfUV1L3yCIta
KVPjc2YAe/Al7t/jfSZWF86R8UKNziXprBlFcWItteyXrhd4zr66H0Q3PqEbMFcP
rdTgM7zEINkbkljgRsYIR/WoS0Bg3GWrXOX7a1fxi0uyUGELrQK/KrNBFBvbLYTN
KA+zzYmxRUeyCkoYJ+rfwIsms1SUwbb/y/+S5eJBWqBqqeXwOwgsy5XJyE/w4PbR
lR7JEFNnHBoXIPha+4FYIQbRzgXnM0bJY152IuIEr13yQmjEje9bufthvsmRaXab
vmq+RRbqAaFrG+6V58jBfCLXuQxJB9YUxxdPsFlijp6GKAfYeKNREhAK+TItXHbb
sz5/+aSuYf7BAWVKdhTJ9P7TUNpeaAvz+2CnPxz3UOE=
`protect END_PROTECTED
