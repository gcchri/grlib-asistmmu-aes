`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4AyPwIMr24kX71nIW/ixiD7BnfFm0Mlr1sDVdKryqoC1+YIkfQ11U7sT24dRehSe
vsai+e+BUpCH1ngFUIatCDoo/IsVGKvhsqbHKjKRfwg95W28c5/FDUQx7xbtkYEq
3xvbAI+aJVBd9bWmoTAOm1vTjrRfN0ruws0ApSg3WuFe3Nz1y7y9ixYUkHw5WTmf
hel41Ik91YCMn1TneJM6dg16uQSn0i497qyMPtziVS7mWWpiLEu1Pp5pFBMZ65DJ
PaTzg+pp1uRofZSl3ABUjjCRQ918DGodkDyCKH+TNllerAQJEwgiAysU4kk3vk9V
zIOUmAYwUa9tOmRm0wGElFdIYTxCHuJkX1WWdqcMeIw/He1WZPitZ83n05gxWdUH
/kWS+bQPhFn6yLioGnGlNP2lMJi0Z5Y6fk9yw2eBD1SlgpdbtCq0hafDNloLCrSf
7SaKLQLj5/Fl5NXWvDWZqA==
`protect END_PROTECTED
