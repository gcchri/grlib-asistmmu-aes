`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9yri4GuMKNrO27Ed72sYWEsGjrb2PFyvotDovjJt20+vapjNPjSHFi296pYyauZk
OYDYWuozFlA5m6tIdyVTFfTTUu+lD5LhsiO9noDG3U/l8hLTHvKoz+qwZjQDPGz1
EFouiJOTn+fRY6zAh3u9lUFFGEFShQjOr+rzK/t2Y0+Gw63s8oe4sGzbo1FSgz7G
KCzEsUFy5hvgGe/cQL7SxvHAPnl4xiYX4Ajb2vNDTjRI55ynRJa8zqXrku9EjfMf
w7x3MgGH21ryP4qxbrEbElQ06lhcZhVjqiQ3ddeUipPq2OWjJpXFt0laBY48Qz1B
AKBdnXgffmnrL8XCA+ODsQEDZBDQZ5W6Xd3Odi+UJ+V0sQIqAsodU4pyB1Th5f1h
kPjJU7dE3Rw3CQWJkc4FxQjpLohLugymaQ8edUcgAlltsL2f/4haEQwDYJz/atRB
yxJj48xIo35G/HWi07eH9l8onCxA+Tn2Qt/n5YDI+Hxa3cVTQ/F1dhjgPqNTnnfw
KroLuJil5dgy5fOB3jFnecIi5KsTk4X9vx0qqGO7FjeJ4TWNA7qcExZkH7mRXDwj
PFSUXjcuYBVndcjc9AZP7YtnmuBYhib4x5WlLtjHtt0=
`protect END_PROTECTED
