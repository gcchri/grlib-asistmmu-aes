`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Xvg9muM8ZlVWUOZHdUY7GtU4ZPzxU7KujGxQjDg2b5XNMCVdsMuumeFeoukzVMr
awrHTzpVLetNdvzVGBLe3sB8ouwspenITkCPJpZt8ou45rfDIc+L9g3EZUIb3/sv
/kcnzCoFts/2k4bkcxkj+lEciz9xSDn+oq+2pRSZuUH6QvUdFQd2zT3TDQGWhhEm
2Lo/xbAvbLJlbjRbjViJmT7UoI9tQFDmkklEAADWTImjboilnJzAKw21JujM0KXy
Ub7+e3XI0pMuw+Sxzi42yXV5TvdLgApKVVwqGT/i1BT6SJggmR+u3GsObJ8DI3So
sr0cXKYARegeB04FOC3Rcg==
`protect END_PROTECTED
