`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AE8Fxol/VjMBNcpxxexFipHOMncvI41EiDFhcW9SDWswVHzZP9x9SDVjBLUvm+fy
8g/20qFbciKYWVh274MgczORBUlZPAJnwoMeTzaxCTnWger9Deh2Rlm6hOfRwu/2
giZVPJIvK0yyfxkGurRqoVHVx4goU2NTvc3rd5kpdsCKJ/QTzINiJpOW53u7paj5
gSwyTEcnU9yqunNxrYDDB7h5k7qoKfbJLdCzqCTGtu6F6t245sshoTQZq3hawqMX
Pw79VPX8kybjLyL4s2Emqv4JMMdV9fTLw7UTOfsZ5Hni8AyxTYJVplIiWGqFWDPq
H3d8o1NefWx0CB3Nqlqw/pptFqMPoL39rIbxmL4NkdIhHzLPy3jB2bTJIPztoGj7
ouVIFT64TNB2XWO7KzcE1CMmS1SzPzQ3MglFcmnb7MC0KWai/m3fAaAhTAfgKlc3
PbziniQKv087WjOBKcE8OE0Z38PEG0LZ8GHfLV2swOQXN2evtCNu+4YKVGF91jKG
XZF/7qy6+yYOPkR/MBho1+OuX5a00WEq4p/Gbo/z4q2BU4csN0fivOn57Wte94OL
Y9OGxQZrfRcHsE4Tg3jmlptDoqVn7FSQPO/m7JacvZvaiCNN6moBTXoersDLzAQ6
Om4NwL+wCFqf1Ouju57f3l32oU+u0AUSXsyowx/6JAPGQIi+RrjtbyUqw7c4YfRr
A6WZeTTihPRFE9ofzq2WhdFCrjrahb+ESU98W+kzgCqDv+gsA+iTWTBXUZSGdbBW
o2EC20PA0725EnXPJkmo2q1BI/loFqBJiyoqQG2e7CrYl87nVLPmBLFC2wqpVWjT
wrrgvr9f6IIOO7GcphgTh3zvJ6GUtYrvNPGOsRAw0JOoFINLgilOFag9IfdmRyui
`protect END_PROTECTED
