`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pXEkTYZ6AbrIvkqGggYplV6iwKS4g69ObgmOa5vQNnJ/DOLFGFkY6ICttAiKE8sf
nZ1ddXL6NHPKDYeMTnZASiU/4yYGMmQHw7SpP7qrp53OwpH0XItUorkRTU4RwfQR
W0TzpA91l/fmfRxomIT+8czS/o87QKbA3hOM7588gSJUOzL3RWbcV592jYV9eZHJ
/PkBmmr3rvEFWCXC4OgqUw+6E7rNc/7CdrnlKSLpBDkO0K2jy3ZtGU2mBoXwT0aT
OPNOYigXVsYM5gUm0lXKd/RLyJd6clJEpYT9UHfeek0=
`protect END_PROTECTED
