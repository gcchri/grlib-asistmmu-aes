`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f1RXg7fnQKgH3Zlb6QQ8p744bSL+7mbUOFPqwY3uwLW7r7INhEv6ajn7LTfBZwHK
A/iZ+hfXtQiiouwW3jUX2KiF1dtvtvfzTM1VuW+Uwy6b0EKEkXL3oEtBbxnmsq7d
q1V7PTlztdAmdNy1KRG3o5Z4uFCK2qJlC0JKbdCCFv9L0YIyo6uvgXnhH/mQBC3M
TllYn0IEj3t1SlLD1/Or/CSW7WDUYzjFSdkb81gSCf0Ml7WFfjIoEeoNi/eAo7fZ
gg6HJuyKV92qOJKEPhqRsIfwfZbFpqJEUjRjBP6pf3UTr1tXQOCtrDb6G1Vmy+V1
27JL+aL9OtPrdKGzlG2ddLqfTlwzuHshGF73B+//p91fs+o0hakGy+2IauJiJYbc
/WwctSqh4JmDk6B/EOo+mPhgrfaLGP5sAM/I3dpXgjKa2fRpIT1CFWc/q5mVA9OD
xQgIOs82odGg0hymdMlOlOvd2lfsbZ68Ri2z9kerOG+HR3gf9s/o73QX1IGyk9Hg
P7o1GlLDtAFHyOvEEWfbM5wv0jJCppCyAxvdAwH3xqsGdvTuMlkLRBuELkRDGZwI
7+D+JGfFSQyRi7NQ3+WXspEhz47sDVIzPgqSfZexHLx5QFkF8SLgltIljSkIHoor
hZFTunwAtymgLRlBTn6+PWX+4RqGKeQOrkKdlMy6j7i982IxX6U/8uvmsgGVFeYn
YAZ0MqubLoKBzx0CldtksPBjvfDwdx3zNXtd3JpZP71ZIBBx70RZibcHIVIKEyX3
t5dy2q0BYjp2DSWcUd2wLf0IctW9ueX+w5rM1182IVYtTK+zfvpZLKDcfB24VRa4
i4uTw0I8DkOZTT4v9JzO6w==
`protect END_PROTECTED
