`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w/f8eIHcTqs5iJdr5NPv+gHwbXA4QIF0zB99GEH46ji1Qob036Ws8PvgziqN39fh
zHQlvmi09j/YPf3FpL0P3M2FnHEbVsSiRHxEEOIsgOrLd3L+T+hdOHhPZswucG+v
pz4eCuTTb92N7u7Xuoje7j0IPi7gBLv5NDx1o5PJtDTNk0S9bTSLC3CjwFbjQJfo
OBJF76pxTEoSO64qgIPFj1vtT2S9qsqwOmrOaP7QRTDckuany4GtN/JnFB+uLzWS
t2fIf+n47m0wWLug2u2cANoHQ2wt347cQankb7xyal5Hg5kW2UdhWCNlBfQSuUCR
ttThfncziqq5QiWxx9Hf8z0UPTryZW097ybX/lPiB2CXWVr0qjqAuzadZ3bsYuXn
JpPNw+uPsLCzS+vkdLsVsAyW+ieeTkh9b6ErHINYyAy4s2Tcf2Zf8JYnaYGJaWuL
`protect END_PROTECTED
