`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vMSFVj4iZe8dFt9VmKzYhsO2iVhzHFpfCBLfxO2ZvqN8nXTLZM47Su1Gw0Ztknyq
cbUi28BAvf1COrsvY6ixJXY2xo+NlhjA8FME1o/2aZLW/35/k1Ffu/AFTMUVi/aU
fuYEo4rFzB789pCWSA/r3gxP28HXwnpIKCSG18Tb5lBTInb0RaP1A88ZQPFw2KwY
e5TYMWHSnKaz8BfoBBBdLU3MwgKHztTzOxdMt+rtEQkTtS6CqKeFszqAM13GdN5l
i2Dm9LYOUb7p/QS/nvUsHDWb1GPyvvuHbiOiXwoiunDwePAGmMmqPSKiaynNwxpZ
gD+B42GAt9rm4lAznXpWQgcoxezCuyTOhZH1vvRDKg95dsU5zDZGh1FwiGvVaQjj
LYuP7zoN7I/LK1zUxUB69v38bHp1ihQu1hb8s3CuV/zYlAcGaL6C+Kaq8a/pmlL2
EHAuUUs8qZaBX/I4o7b+rTkyhhKgNb1bur34aNkkQ9fuaOl9Zi2atHhX9/LPMEDj
`protect END_PROTECTED
