`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T36DYasTvOlsyHeNf3RF363e7sLX7A658gGElQhcxJx04gV8+sphjJxOkSeIl+BS
4Zeu1Na/mMdhxgia1I5lICBjld1XFC7LeTOIL2iTVM0jDWk6E2ooY3L8AQrqLLK8
aIEDme6BComCC2lsx6HoUy7ZPlFv3BcwzegLk4bK7JxHwgBeK2xVmyfNpK4iXpng
+xzTf19J3Q3FHwVr7ainCV3ZTva8vkGDwArzRAR/nZxDPppmHGIGHu1r9+FmPUNi
oNsr4+eYEPsrOjZix3UFqUrsX10BI+wBNuT6UXrzFMoaozffgo6hV7FAlT467pvV
ntzDnIV4esUSZ88moDybOkNs6fNe/aMAs/X04LtFJMwVeJWtkFMZA2qmQBKWz83B
Zu6HuAIY/fT7xc57S1nTifYQeB22nvSEdbDEvDRpw97UiW+ugV40Ll+nksO3BQlm
f0Zgk7tFEnoL5wg+wpLw902xwdrucKEY2vATBwjuCaYiNzwD8aE9OZbNAuwJMah+
i/uXeUvCqcdzTIjeHhKi4iFRiBrA0kZpxptl5LHNHN+glGvd/bW3K4KmSIvhjLOx
XPFKLI2Wr6lgGhtwYmcAhYmJ1xFBssohcw29x6GQnC9+jhX0HZK+JeqeF5/HTGSn
0Jkh+p655vG+qsPoiT3S8IhUv36LcP/R8kMnGQHHW/sC2v92DvbSCzMvMPUEDSKl
9RuHzi3YvlFhlpDNjnMUROd7eFQGAaMXaspv5YBTVNbfNGPSOt86dfKcFc5MVLCh
GqRV6kLPxhr2TKtenRRYABHSdMU/0nsK6dSrC2wxtyLtTVvQLmiSItN7lnY6BsWx
BcdIv9O2FJcKda+pkIlKmNQGnwi7ALDzsDqvw05YhGv2qCZPt3uz5FZFBiqGS44N
Ic5HUWi47D+MVVqLqba7Wf6Jpna0iE7Yp/DUqvwa9lqm+oT2K9bJaL7y66kaeeCG
`protect END_PROTECTED
