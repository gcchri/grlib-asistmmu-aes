`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5M3OYEOwM/KlYluUenOFqZxD0nk7HavhprSsk59aJIEMNd0QbLMwLJo/G7hKdsYQ
MHtNu1dfsOYFN6HE3lr5XFyGa2kWbnrn1fcjYsTYJwmGc+Bdirlq1VcY1BSfrjhN
UO9nS0OPsLeZPvND0b1m5PQ5cjf11eNk/dAsWUBeIrl/vCP70wkXw3BoNB0Grl2m
DMTehDRHPP/bd0op69Y/jw==
`protect END_PROTECTED
