`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oz6zOpffnQOBLgjaxQKdI5qNZgrLJs89uCsopWqb3Ci9J003tpVdeoRx61nYq9tW
YoDbl6wq2rqALvU2wYEWZfan3Pvk5Xz97zRgZmogyWzmvdptqZCOPWkaIrCOIGIZ
O4/r8hyRsy9tne+iLoYmyxIa7DkPYtJ/r5y0CaLUHe7oFT2d8IsTBtSh90xkEYHG
LUCa0ZPAIkNHGflQfUqQqYNMftMlZQDW6jdaDXraVcZkkFiLEfBjtPuuuq8V6mod
Y471HLNlUG6YJj9LnPNQ7B2Cnp8bLxsvq/t/o0V8rQzUnHCYng3OpOgh9FptvZyK
wuwDZ7l7VSmgjkd2WmaaPBFMY184RfePcBn+qnPUf6Mu/3PZiL2/WkDRde1XAdk4
5yKdEb9ejspkL9qTTWcNlRcmgdOTSGjYK6OoyqM7U2KCKwkevqMxs+z07J7MOWJL
wnNx5TqAmeBLvG61PZj0pBAZEH4u+ezKNS+VBVqZNxxWihg3Jr8i/iG0V7BB8/Qp
89p1+s0lLGj9+tQomUW7mg70+2khBAQcdaGpNi05Ox8pylNjmXbIjs3KElGxDgmz
SzVzfCbMO5/X+M8MNWSLC4WU/FuHvdOWsmH279xqR98oE2wm+nGgtWDufpUWmOXe
VLVq3mrc9/VXOASEnm4zlXcOSLUgsP58c+gt/D89y02ji69TcfDi6awqn8ZLaRhB
`protect END_PROTECTED
