`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0kHtimfcpMXWx85fo7qGKxk3LWV9v9hr8pLTP+tzzjBQwrTWJDh5Z4YNY889oKdO
t7+bKSiDZp4sSs+5SgFBvwsl+3DLEYNs0HrlBKYT5XePs9gnUd1kiEWNxxuiSdwM
nHVI5F+GVVjm4g4S9/psiqn731BnO5OaUZcmGFCRfcM4XN31s/WGy6gKXip4MazT
BoPt4kM4ugNX9I8uG/SLseZg9Jwz/XWeoL5VngGe2CKiEa5inOKwRxUQ/J/A6WgK
AmpzCLIyNegSajaYpjuLLg==
`protect END_PROTECTED
