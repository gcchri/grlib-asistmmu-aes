`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z84lRiGqWCkg0X4QS/YIyXlQ7PXha35XbDEtER8bwJK+sfGoqtZvZlkiGIioEb9y
fPzL98B8aBjDnMX2ZbOnkKDigFFFKTStkhCCUGBokSJK56OrF9in79G97yfEUo3f
cUddTGOKls7SHtPG4Y7hSgwZPRRDmv871C9XDJKJ5F/2G3ctiOOXoF4dU6QfGIPd
KjIHHFhIgotxbwQLyb0Cd2rn1qcWIpLEBMm2yrmQu+95/Kz9xITUUor38eLECzE8
N/p9MQAnImTV7hgr9jkQ+NPIdhkA7aSfcw1cXyVA2wb7q5UPdIgDHsp+uq0h6lYy
lfmiEABa4Q6aHB2YCux9cRVM/lXEtakkwqwKBNYz6HvZa1WYd0LOnZLTRc1dBW69
I2qUaJCKDmHp070GSx2BW1oG1ZNME6qYfUA3xWeKccI=
`protect END_PROTECTED
