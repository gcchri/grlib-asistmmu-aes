`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
osMJcDc/qLoxdp/TZ64rK+IR4uIo9PwYdcMh7WYPyYWhXqtVt0VuDfGeYXHvsx1w
eoOnUZJ2v3pvEeqfLVuX90xwEWn1qLeccmsR60D2wr9jPoDV0osClW9qJ4LeHTJH
hY5NB1xAnuFSRArT4zkGwzIy7rY1A5MGDJtSuFtQNRuIGbLoqGIZpKQH/CULKXpS
Q/J50K/a0dnfT85O3VnPcgII3oW5V1UsZyeBFuFCzR7UoPj3ZmfV8aQqbDp+18t1
Q/elD3iXA5rfarFsTP7fKuTVVOBgIC1v9ae0ouzwrIAvr4cvvQJimk+afnL8nYwd
LZCwh9KMfwuuFnzwvhQBO4jRk6MYjz6Xbwk4keX8c0oE3kyVEyCfSOwYZNESocgC
DITdLLL9UbnI8fgE/A/lF/7cketAFeT8fzwytUPiscaeNfs+O2j5YQyz21mgtXTG
bBeJbPeMTfUZFnmBmBfPtz2zTt7+IaA8iL43Vi7ubH8ZT470mSa+sTBykxVirDes
PAi/xCG5kmOqb2O9b1RuCjZ6piJnwT8+iVsK/WTWI0Q2uFWqi3CX69dtXxKRE9BK
HfRVpfmwvtN8a3a6Qr2hdgP6NUiIfQGQNDc5RYUqEKPTsFTCOntqlwikGyKj1DDH
Wcahb9ZCjVyqTVNuSYxH0DpnsiSThxC/T66v/+MteaL2WfonToPE7E4w81Lu2Lzd
rrWH7lmomruEcIWAYKmxfWtzWW8Q5NpOT9JKOp0gvkuEnzrNXO6smlAgpXWF3jHg
dGQOeqAKkxCo1rnG/XJe2ZcPWO77EbUC1zsvFKiSiY7TZAaIEPrcpwgXVM/Bk8Wk
XuB3lYymXNSJVETHpqvLm19Mt4NUg0K7K9fPidC982HRwXJQdDRo9EEc33GPXiCk
vnVaJdw7TUDRD4RCkC/AWr7UBY9IF87Eh2DPjF/RxAQzZknviKdVzWtMphoqTrsv
`protect END_PROTECTED
