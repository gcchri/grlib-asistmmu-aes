`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IJRuDZGVelWzgA//qlPOH/5qW+g0JCpr3P5gWGFuZ4OP86pTauSw/5iEUGHfX68H
J2ATIpy33BGU8AugjDsd0n0mEhlruTdLpiFUsAl3hHtED7nQq27owg1izZ4IVk2L
+0a5Dwd9byxvGGCtfNC2/iZZwxK3trmvQ50CxBZuyStq5hj0sIA4subuuGLHe8uH
p7l/U9Hso7X0/thSWRvhQtPjIfUlPSf0hImtiyawxXklkbTM0U9ufD6hXXUZbpF0
+ZbBeS0bsAI0NvIz+g1Z47IP3NSYzGSCSXWoE7nFMiN+3ul84/yMkqv3NT5UudLf
pTxvYgrNupOOzaS+v26YYIxD6onJabZvbaZ0WliQ/ibKSO2hBMPTWj4Hnc4kx6wY
gCIZUT7qrJM2qkwHgLBIAJEuqP2/LPXqy2+K3zwqzevzttuV5fwbBjK2cYUaLTxs
uzMD7pPOD9FUbuM9rC2onkiaNYsbDF39PUISRixe/poo1rcrDe+H8XxB0VWf+ZzM
E8PpknFJ4v5ZXs6Oweh92w==
`protect END_PROTECTED
