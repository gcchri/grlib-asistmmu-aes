`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aDHG2BNeStGoiYEQCgW8emaTS3JO5oicL0Uq6F9kcpauzk8HOj46WduBtQf2o4Js
mDUYRSZYYvTQKBQWn5g+XGmrubwaVAJ7RMMvCacKyOMDGZdqJT7Lc1BqSuW3MCzT
YiFGxGKHj7R9HbSdV/0U9EPWrWCp982X2fgLij3uQwJn6kHkpvPxnae5LSrZ/f8v
wX3aChHk/wPTkHac4Rd8+/e07/1DR5MO+Vi5WOUk/2nGX2ub0eD288ixrYOh3JCu
kKYFPOMUo3QYtl4FfFUGFyKFYvSYxSbkAha+yP4wGJlNaYPSjMOQxK1u3QMS6GKW
LAGQra4R/TRQx1WM9ZIjRjYU24gWVOFFKdyr4j9YDONCiP/0F0paXvGKSHMKqhsz
Qv+2hNvcWo+G4FXVzyAd0A==
`protect END_PROTECTED
