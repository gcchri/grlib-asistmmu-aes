`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DvTVZST5ZFnk7I/W7cUMdh+H3rSzwDzLPv/E3F/o4+WDSIE6J1mqN1c0+KJqw8LV
9N4wFl1i6x7V9J/cXX3yeVWFr1tALigt8Bl6EfW2gIVqZJTOymWud8T3HEy0xKxO
LCZNfPN8Pr6cea6h+jRWsD+ntLJZJ17p8XqGUMgmny2XmAvSzu3X6zbUpen438++
n2Lqgspy+iW+LyMP79i9HdHR18PnhNC5fd5KaWqthbJKBaPgAnd8cHV467YKCS2Z
5HwiJJEWmwT/5crC/32pCH3AYoxoui7LnzhQ8JZCC3UIAeao7s07xUhHWYtgywYV
p/0hXtS5pi305oXBUEz2YChOzoEa/fOq5gXFzRoLWpKHpC48Vq/slveP099UX6AJ
T3rmA3+T4mw3HcnNADIgKUa92aZVG7V7rJI4+/ijocU43rw+YK5CH3MwiPUH2fJ9
mKXLlCNeKMXXdHC21aHltg1RX9xhR7dqjptUIu5Lq8lThJB4qiJDVCSmGYt1wyca
FbmCVflCnIWRG52zu5BhIOdKiH77LlpyD0BuMedAXuz4zQzTuTzaTlDAmzhgr49y
IVh6HMt5Gpdy4FThltfe6usq+Aynr8Oo12VzrUuvBV/jzJ+mPMIO66qVzIjeihzF
GgPY0ZXIK7d0/D57ntOPwRVNckIHfapy7qddU09Z5e7lV5djhBR76VYN8UAcw1Jq
pQ1Js25ZniYBAeiY8kCN3cMC9WNYcoWujO1FstDrICh4CsCD7AvNKBAN10iITHBh
r+5ZmxuPY8kbMjMyeBXraxpiurmIPasJSjD+pMjZ2WcYTsaDSjfckSLC2B0iL4ZS
HOwoV768ddhVHTKA54rh06flJRl9TLyY5AJZhdS4DE3Xeav0cSdmfTJICv356obH
ymw9uHDGwoQzL378eWKx28M28hNji/7dWXz+m2KRWY/wvULopg79fejQDWCQzfd4
tTODxxn+8WXdAKfdSco1wWtNFk5xTt8ZCp2wYS5gu/iKRNM6q+bkLw5ZmG85Lko+
EjjErdrYzUU9Xu1x50/J48g1w8nuoj2C2cYlpSKbhr3ptVQWQffhERP4xQSr5bvN
88FDy/dKf76F/43jDaE/f4HIrU9Q2pTbP8vK2f8nQEM+Uz0pD+c44gIN0XBU46Tj
QWOEh1GxNf00D6nT4kGis9r0Ce6lDnKVKOGRpdWhm9GSa/fhairm4Wz9UzhMtblx
UPZWbGSWjbEFe6+rw37wIPN6uPD+EfKmVqYOPMmtYRaDdzhaFQlqd0mHfpySSwe3
bV6wdrXWc8Q5hH7M06ZJiGWdQmpvpJISauDKVIDQZitihgCqhlMGQ/mNjzqHbHMw
lPK//bFviVY6pBaNV3HjITZszNSXUrnikjTnDt52GuTNjO3eOlClFm19njm+jIua
0OqqAMrqlpobC2rz7kGTgNvT7ObjMujqZRV/3x1Aa1sKKESU+I1CAGglc1YjWLCQ
YrlGEPHVx/8NGryNxFonQ1hRltrRajsIkVJwcOzCmXEvI/SzfFg6jZOIVrSyMtof
ZRI2TkHgjLMwo9/7Y24m2jhKZvAiTMAzOxN1yL0o8uL2lL9izOINpyPFbSRWCu6Q
MbkPbsNsmJatz3atig0sXLBUB/leJEz+LjmXvCayszJclr/F5ZD8wXc0p7vQOyVE
u5VeeEvIxwJhRAJUZ6M2+APqxsaIrwBb68Eq1o/Osf4SLgjq3g97XQYL4cu87oRX
ZhAszkZMiQw4Dq2ayWlFYkKb8TCQG79mZeieO7KGZ403ObfaYgpEyA6kqqEz98Fu
Ayr/FkaIV3josQxYgPVd4xmzHPE5ptfdYpqJHAPk4unqyw9aFeW0Ef+a2tZL1Zwu
SO2aziEgD626+u66DDKBPjOUxja62/78WCuGdgW5ToDWGjQGZ+WdW42iBU28jmsI
TAWuT/sF7E0KCZJQv+2d7VL+vwwvGkzeNUsSX9WN8fqoZmM1BNUnuxAeo97Z3bzj
FOmUs5F2ubNHmv9djU4doZQ5BmUIx4PD/CQ/iJM1AmpL611r+2mI6zaY5lKEAzpz
UxdsM18+b/nnYZTKvmWzITmGlxumKHrIRcpvO0c9HCaWsurA6lx+7piYVibJRHbg
p7DZq6CuoVIpMWDJQunDldzxOrJNN/ogScRywJUx8jZ2nNgGQ0pePfnmqLgrzuWm
9wAkATepn6S+flYnZbTZQoReyNs8so+Ufus55dLOO4m1GYnbSKk1V4vvsQD09P8E
y11z68+Nlih5GRwoK3wjBJQW5FtWsk9ssRUGxt6CzfKVzc/oIjNZuO+1+3LGx0cD
Zzqd5spAquErU8BwbXxg3oMJLIFUHRe/71syPbMDo4baCQP3GKNX5se4yemWZsgF
aAbrEC1LbRQgGy18vhSq+najtCDeZ35O2eZHuufR0C5gb69r+jpzzTxgKEZ4IBnP
vQzdnFkUoqFcUS8XFz2/syLuWqgAgFBc6I3fHXGgJ1YpIapUoYEkXUPXxb/AgEFV
eqOGUz7WY8gbjXl5eYJXhwH90PiP/u5nFFz2rDrXncTFLQvSDSULjlmj+4hwehap
gSsiqkPMUNFqDexX8Bigi2hxTHRDexdH0/pprbdyYP1V9wAn5KJhgGPdJn2kA25d
mTpryHVVVOOZItOCfRbOvusJeijg42HXtRdBy8NJ/jT6x+1cRelVN1ufrSCGS5/C
CWa8kLBAW4IVdhMxeje5aPKr2NjjasD0ifCcdpoh7rLTD2sxQMnoBYGU7XhHHj6o
twnxNJpfu1X2VPbNOX+8bFXkWUWa2xHJielvkHx7Enm+oKmv0kMsV7FwvN0JN8HC
1By5J2tAa0AvmTVNjRUOqyIWBW685Sy71eHY9ZD75CcdMatyA41O+LAPfDufSONP
Cpoi/0o5swsPZFg3XRZOiApeoOYC1YVIvcxdY3vj4z0Etfh7HvHKwpLdRshloRW8
pTLKoYCUwuoDeoz0HcfWvN3hxdUsIdM9VtJyy97+sZBuIiN/PW6ZiyKZ4kU7mu7J
EdvYI/sogAS7CQ+edC1cOCkXcDC7cPq4ejbpwfZAKmzwZCTUjnDMJ0iljYCRekVx
DMKxTSTZUZutOfHimHresW4EmKgvgxzspfqq504XsY3Z6ZPfTPIgQzINuHdj/rNA
7iMPsEIcN+6PyPjK1JGP4+HSBM3STdAPCOCgMqhH9zR0NMAk1L+TP0PgwIIBrc78
Bvo/Iq90vSouTWBctUo8kH8eLj5wPa2amf7KsNkS8Tz/Ob5xeBLRTzeZamhLS7GQ
aE19uw3tDBN6P1DohPbAGg9f4BzAOE8tp3Fl0PPc3gXes2FH6ythpG6glkEXd9ul
wvHQ/Lx+wQWYOnau0T+zlRZduj6YGxtLJunEt6BwyLw8CnU/thfiq+yfbz0JBNYh
sIUlRQMlJqvZvEaW4hz18iOIzQaulxscmBb8XxXdHSoxuZGOIQLEIqYBPFRVmnzH
mei5o/9kSGihDAo1OFywL7hojekZu1jbjPM3u2/Sf0GdXirb9TuU2txBw4j2DDRQ
cLpMOVUhYfQHBvgZxFwba/v0WB19lTIQzjXGaiMMI42m8Y4e0DZUc7YnVQq7HLG1
HFuseR+BndLBdenodETb2ix65OzheGQr1vGRSHIFUWcVXVIHk/ur4xj8A9sZixCb
1lfXR89236HqnDRA+2jh87WxSyrBc3qdBh9h7GIJRZcQp6o/i/+0IUqvkZrT+uIR
BeLdW+Iy1iWyGlyyNTyoVhRVwLaJN0GP05AsJHbiGiCSfVo+48OVIkh3hrJ5LJif
bI8mNXUQFfjYG+NJNlXi7jtuc1/ZvS8+anO8zuPRtlD3OqSCcoy0IcadonCNMLY5
0YHApvA5gkPN4fMcpDibs7VcXl902jQHEt5yY4Wof+oIl61km2/SoUGsItU4Ym2n
nIa/y7eA58uYZM4/CZvoFaxmicSZo+VqbbP6/+W7if9YKXUmZDJgpFtYqX6O3E2r
J0fnWAN6xY3Ql4pNDymEjZrxXx+d7H2qNqO6AldbEAb+1TY3lrGXYsWRYLxnYo4+
Mpba7PTnU1O555zLq9Cr6h1nrWk8+tBFCKRycoi+5wvbZj3ANxw/yR2eJ9ZIH/BX
4dUgAf+HyOPh1OiJ4CNsmacagv4vpj90qU/v8+Ptk9VX85TWeMGfZquVYjQcfXhO
cYcBVYLtATmT/AgUAPkY6Wm1NVvxbYeT4xs7KY6MjShie8f7EzbVGH+RHzHpMjdB
vg34/oReIWrqf12Xx+8YbvrRA7hC1A6mfjlPM3dxdMUaid+aZ8EyYF/hKmiCy6uf
WpZsx1QEu5+L1h4l8u0xhP0P+1+nu9JjhLzXIJtUuJdIexbfIUFWMSA+C1dfF2QV
St5eDHYpQYxBurEQQ7fwa3PTrKx6KKQQn5LnTrwGrW4ivA3mvDW8oUSOA0K/N7Uo
kM74KOa7amJebfOpPA7CWVMzUY+fHuP1l9jLYBj0u3b8xeDW9lRwbuPrYOu5b7DZ
ohGqrbPraLU4goD1/bdkQQZDqBjscoKQtn2dghKZhmQUMozuUe6iM24FQpAJuHBW
zSALWG7XQG8KJmrBH/rl+1hYfBE1HyCD757fw7TG5o6X/JXkIB0NGOfC/GHTY7eJ
UyF0bIrqS2AVfPXlNOh98+GQfdhtKRBqLvMOAitojRdxdHRzWMXtuc5RNlE7dhXt
giT2mLDVQqr/VcYqoV7qpBTLI3jXK7+cZpL5QfjHTTyKt4TPTCFBaMIwCy+ALrJy
PyFg9d9MIUZpG34tbjTWXkL/Z0DqPEVfVi09Rc9fKq6rIYDF7dDWGXhaPv+pNA4P
U9c7HhkKJw3P+bvvJ9uz65uwIXU3iRWyhww0NhFhRPTgv5CDwUkUez/1AxzzYetl
mQil+gaHzCVa1EAKcBRQ8ODVwwdUv4TshIzG4fmY+HfwkpkUA18S2ecphqsMupUq
5nwIhqyswkcY80mWVn1W77kLinZqMGQpIMgro92S+TeleCJ4hD4JI43oOhkd3KeV
degzrRejvaleOA/u30Ca+YhglmCXR6PQF+uif6pVr2NDGwTc1h0JLQ2kfQzjXI/p
8+J0V4KVeSAb7grcK2h3zHVX8rGauNhwl2LHeJbwoktbzqhWyfiNWAlmmSy9876t
ooTdadehQN9zKZrOo6u/HJgis8hi13VU6WZoLtgYzV+9PZApDGl0etgtgdCFDFaz
zrPF8M3KhxUkVbw/rrC6UuKqqsId91yz+XqYY0ooWoCw3Cp0tST4YyhlcWwBQEKE
i3+bz8Bv0HYyIGI5Bd+mb+P9VCg0DOEYoAYuJgv4jnj88FYaUwxMqxAlizDb8PMy
EYF0tn8Tvz6/S01U2dSu7n5DIBWLAfFSvdBAd9mKxBvByokYR1wMw5H+nNMo6GRF
FbnK9cjy55pQftdZokgwNe/siDFcaGxFiP6/qKElSQJz9XXzYmuJfb3ub1Z5VskD
a6JrbSNGYB++7Xvq1QaHhocQtzGUYWeYnR5xwTZyl9Z6plutYNOKOlH3TuUuL+x+
eCDw6Kcy9OruVhgIP95XCa/neuirkZkxgI6VUsuCwGAVbbQXVopBA6yByfdBfpNI
JwW4V/cz8nSJ6Hsal6tvAz6o2rkX9bYVHzobifopA4+6WVexgW1eUehsj2o3GgiQ
kwNtX2gZqbZ41u55aaBcduuG6wWoNHZpSZwrWwa6hV/BvD91rwCHa+gz9vDaExFw
qwMPdDDfMWi5cg15XyQdpbsUp3Y3VEcczkpB0g8+8RUK5LEVF0zh4geEMQZ9rO7g
mK+07PLvYBfYhzQJGjbKdTvkIwBUX6KkMQTyQTDuEYm0DGbpDWy7Y+73G87hJuyi
mF6wmmNhmCAUpxwNzeYz/iIIK8K0K1D5ExPuUG59pu8LG+H7UtORCy/1VY9QSJ5l
vX3v1S5G5rBfyKWMc0dws7VK7cK57O/Vvxak0k6ae7cUgcKyTqlIQMAf8811dn7a
hFH5NKr+BGr6xVd02V9KVAoLGZZvOcsqcRH+b+zh+tH2E4zSFzg+gPIrkRTzMJX8
ADbnClXcpA6A62mGIycuexMiAo/h10f2fskNSajRwAN9i2hJLeATz0PWAmQtzGEe
ph/GiegLF2cQ4RCbesXRhHQVn5Tqglnwk+FV9LZGG08Pfm1dEJyntRaXwuhBueDQ
OVexU4gT1MxBbZ787TCnpGPdVRF2NnTKB2/cSR2oXeZBUOf7GDtpf/orZl1Kbqka
WpLqZQ0tfzLK0Y2Sq0C/LYaZOqfhQ5T8Mqz8x+7FuCdS4ebkXJ4HQcU2FEOp+l7q
lRIehgLY4K4YI0i7QLc/HNm2V4ISvCi2jbVNu+odsEDwb/zy+eOAKHxX7Ksgm88O
RM5FXAjduQFBDN/Ul2AYJxOgZaqT1Pu6Flndb17QwKqmkqwfitIo6EA/W7noGfFv
OhGbieyeGIVIRytrEvqoFmuLb2L4ssTcvwchfUhTZVdeQpR8H6bg9LK6T2PLn3rC
eqVYlk4OsELHmzluLSmYXvgp+LVTbrWlgMjPZgV45a6fG75CcQ+FIagqOt/qxjkF
bybnf5/vRxaQxuW9WHNJy54Lok0mR75Fh1Llc5qNHgdQaCP52qCXB49a4PUyKd6L
zBY73rEKp+Nfi5Xo73+wDgNip+lEgO7igU2xEaJ05udg4057aTP/2Ye9U1vPGcew
Pq9dH1eqIqBVvB4XhwfTnvmyVD3yQTd+ifUTUvH6I6xVk8fpx3Dr11m7t4gS8wQp
Mu/0KP5F2esg/IvM4SOyomwkTXWIhp9lEVihSVaUyRqNOTbgUrg4Gh2DDzAA7nzZ
G2JJ8zLfCsQvRRzbUQ0Wklzv6peN+VMHR2BnxzyoV6qvzJHTwaY/upjYz3sVEwb7
Nt5MIArz/7jhl6+F74WkVdlJ2JuI/cfg59aQBDsrhrX6PGs7PHVDZUmYRKIOlQTJ
fJGvlUnZMUOAdDSJAdVK/wgLJ4RArY7qw9chuzhfFVVg4eFErIMdUqROrao9LMER
UbR/D51jXUbOKEfSRCrhrMbcr8iuFUL0oBW5WoTRPeJjjwvOOhAAmD7mxqKLkuFq
dL49SFL5erf2+vb4gSpOggap7r6o6GkgHXfDkrOPqgZlsVidxuglKaeJmYs5nPnV
ayOY3bVxUn2Mfh/nl2UFIdQFSWRqLL2Qxv0P06/N5y6D5GW3Vv/Qn8C5GKFMYugC
nOzdUYnUIFr0FeM29754Oq2wzLQ0BXcjYZ82muJZumhwa9w0nRIVMFn9CineElX+
5E/aNJ7w5hImgn/BWL5vkA7XN0ACTYv6ZUf9WoUvdy8K+1ycdIXOHpbZNFMYj4Sp
HaIwLKm7oehPZN68rMPHM7dz6zuXm68VDTQrcEJavE1xQqoehXzHae21m2lTXS4q
yiDucCi7HvgHkTwPNTfIoW4ueWygUfccwV7vqPsi8nahEOo0YTxtGytXPBijurR8
a5WySYAig9NcNLvaJWqTnPpmC/b/axpRWZi9SzswSMWp983e1LMy2LSkNbe6FQ00
laccjH6LmQBEfgKo2FpFYMdSf8thK61Ht4x7vSp4MFbHB83XrMQOypWQtKAqsbQ2
lq3bH4xqmtwDvHgbcDC/AqCuNiAlBUmSVbe49psgRjbTvgc15XJsOaKF4CrWjNUa
c1D5chhkSfMconpwiXeFMivjus5kazb/GqtbI+z7/EE8HFPLsGObwIvGMIH0Ade8
fdghJH/E5xLNN2YwLhSpy3PGcOXZQR9GD5Yf/XbROtinCIRZqd9h8ZoAyaix/f5w
kBagMWAnFeQTgO0VuSjH9v+4ZoH1XoYBPjOcmO+iJ27QOjCEjI395GuWq84LXZo1
Wu8P0drzJQ3y1oTxvr4Ug+P3ZMtBNsfOZqTcWBxp57L4WIjpUtE3219ikqoopD4H
5CmFgBuYLZiGXimQrF/Vzw/GvoRZSbe3zjlYOSiZK3dlUxK+ou+kbQ891BL60m5O
dMP0jkvFRBtCMbgXINLMm0e1iMxthL1sSjClIm/cquZ+c7DTxQZRROrUCh5BQ6wR
vjbPMTaEFWN6ezSBICHEzVbCfnqvhYWGLeYpTo1pLpX5nCWU2ZvvgTHVooFFe+oI
MBPB/qYLpojfi1doMwlXZfpFuzX4OcLIbAwlFpddwA6hRQ0lJ9oZyze3NwL5waIW
EJa9O4cl4pb+dReY6UOSc4245e06GaA3wKiCS1PfJbMAzm0xnk5qxH64aFo/r/mk
isUofeQ92FljWLTW4iATjPm7HTLUAeiTM68gdlSfp6b9CfjSCHkW9JXbyGFq4NWa
naU02mhWUpWifNoc7ch4Y2ejZy++zIdnMiiz/RvP/h7pjC98eclTbf4J5csOxbWx
9xG/aaJgL/NOnWNddqT1Dy4yTnjhP4HBZdW9mITho1QtCWyxMXKLwxC0IQszWBuc
xiRUU7/2pVGRw8X8AmY4naJmB2irpHccg/KmXGxV6DxXSW+gpfpkFQilI3EVeVZM
Xuju08JNLQoxzjeKMq5H2cwhWv6x6V1Q6AIeeG/rCFP+Hchg9fsuydGLfqE3onoq
mff5GVdsRw1duLIrnd64JBB4KRmySJXUhKkWBqzj1d+V8tEVcIb1F51abh2OpkUm
5mDn3ejyPSdAQXva0i0AKWkEC32neyfgv7BmcAJEP6GlWbPIU4aewAhXWIzSu9+U
bwwFPsJVf1goMgdNvlJecWzG80oHgwmiQ3TI/IzhyUyO9fKeR8XjG7RCmefkJhV/
VitPZXuB17TYSWPfmV7UXg1n03B7s/v1V8i7Xf8LqG03CkNPgk+ojx63oX+6kxDR
olyYS021HQtwiCWZ9G8HPX1C7a5lJOLfaqez7DuLTF0zEwNdxM4RnzLmvjft1TaQ
iVi48+Zid0IMMa+T+hd5btPgCUXmnZtHoSWOI1/f7RTqgY8iVLplp3Az0tgWmnjp
SFcmchQ91uFwRWI92oZ3Pbnk57UflQwxbkHiH3afRCMs79jzNnbcQJDc4lTXGkth
WqC63PDqN+GC+c0BL7K9JzZXHwo0d++nHL7NgGI3/NitJ2wnwrfYg8mR/P+O17dp
hsANQnFsPtUdDZ1y/73GubchNhK99+Tu3fPuFCxuHk4ZLibEm+lGBdKRCCWOojPg
G/xC1DdjfooKVDmA21ZAXm04jf8iV04Lzbq6+tDXOM3BlBD4lDi0eWCceDLPu6/m
GcBhRKmawgspCfwUTCoEUIJ9ey4FltcVieS9u3+/Ke7HMajKLQPRTD8m1fLZRc2h
VLtKeoPgMzQR5XzKvPws4IudRfLSEzMH04SaDPfaKvKbKChnQG+5ZJNKuACySH90
CVP61dkjjZ1qC2IQWMXeSRBKTZlCMe7BeIF/dQPKKgedgnRXMWehrZYBbOC1O/mB
JhIsAVw7bPmqIZxR50pLTcB93Asbk7G9a9+EgThn5+IyVMw8Dd0N6SQ645cmwwMV
t/8MB4d1QeJ3a2odQJo7Wk8rF8N6M/Vq7tFcOexP3DKpbErNXF1L1Gk9qaOpGxpd
1zGkIzig3TyobbJ5wX4aGwZOEYg+/g1FLyvkTqs/HYSgRAZ38pHsr5byOQjCI37d
/RHyJRh6Rn1+m38UN4qcXztldw4Z8PJKJz7LopHABYX5yskmBOXlUp9LuYm71w7F
xjFC7IYIHVLdmLdBE9Im0f40d39ZjUJJ7sS1rM9iX+QQWRtLmzdmxIa3uiFgAQyn
+xMtz2HPkWa7ColG6YRUyhOCfl3d9Yi5hJtgvYjNDG0Xvm5poaX1dfEge0j3i/Cf
CDhzzViDUH0B1bb8V6XmpO5iDGu6ONyzCFE2F4VCy79FheTcsBNImHpjHHXB0Dg3
zpTRgtS3jw9z30peizURl2hWFQAYvkFByOZ9EywHrte/jUGOUlSlMzV0Bs2/K7RC
V8dCDuT54f9geYQ4W+C92ANSF+0A6dZ98izBz9Tk9U3pJvd+Qz7yHpM8d2vzOXWa
FU7v3UN8Cvz1omUPkupU2H4jlk/YVf2o9rc/b1uabQg0Fa11CyNDOso8zhzOHpX1
Jv1vIoirhSNgMi4QROhLXlR8I4zzQyMRXuhvf1NiMQqcOkiGLCqq0a8iiAQDqvQa
Gy0NMA8s3WVGLkWTNoCroIUObtmmPAZCRLtE02cecGtIztnCWCzLPSqClG3JyWP0
hUs8jPBgf5vkoZ8eTcQjWoPRHHPziW7fYz9HRy1WJxycKEVJSSq2TmTybCLAxu/Q
UwBYW6J/RBYcChxUBAHCOEuoWAhEdnAv/o7CEa+XvYM097np/eNjC19qPL14D4RJ
WawCfb1ctg5oEEw/Xgp4KTcraAOZQlbxYXqKcAzAYpc1WYlDuWvju+LiFDioYfOU
Q/2AfItsLJMZofArgqU/426HQLkKJubTEV8oWIrPMlFaJmLsW2sP8iBrhwxlxBr6
lB2EyMnZh2NOK/7xyCWnGQAnQL0YZ7mWqahR3pB1oC6jqOEPmzCUZKf7rbLXvkRs
jBDCAjNruBwasmgjABpH18HQcJqtDIKz18fi0/uBcUt08BbYSYEi2UrRw+c5T5Qa
SQhJm0SomOmxLbjSSdGvapoJRXc8BHpJAtfw5gczvx+K/m3zGD5xrt6noLUGckDA
h2RHvV9LQC+cQM8tngKNq15aasVxsD0DKeJeH5GPaYMgqhnazMxklvxscenVpkWw
JTG9qS7ohiMmnFz5G8ABeUI+GqTAgFV+XVtLxTMGzRun3PjW6QUoO8HJQzUr3sCg
uHsg8C54z6uB5QIC6p0HLO5RQZox6vsQpfGYITCiVION0ZDaZdy99lk51RUpbFbe
HhV5wfy8jfCRJW5ElpnQ15pUBNs1/ElWK9YSIcyQsLpfG/VVkB5El6qq/tGIAATA
SmorAPvFjhxxDykqcWMNaEKA6KD7yab9373SrYdKmOQpbT9MBsavVtrZ1+7GqI1l
n0p0jwe7YHAhkPj356eoEC2ORGsE1dmPwoPNHmgrA3Inrgqnxv5WU1+D47t/YpXV
6MipBPfMUu4Nqweokg0uVJev9gRwOqAZY3rYWUmXC0dbZ9Sbp1hyAM5lEOfKXmCO
rcUwaAMpSFgVkSbABMrqmZMyyjlSGbR4pCbMAVIYQN2wK1sTIU1wJULrUYJ0yobT
rlRoZA6m38sMP9Qkt7MCZlvcERCiRLy6NocRcT0QMtBy5W6G8dR6qPNyua7+Dq22
ndFwcDUfm8lI66lr+QCt6LnN6DxDjZBGKAE56fqHUs5HJxYFuvCDWTIcjmNevrCJ
a0jwyrIeFhuBUsaAv1O4ggWSAd+tRsGoaY4cEgl4wCSVvIvOfP0jTSEj6NUdA0yC
hLPEkGb/t/1Do84lKIYAJIV8amcD5Z6HB3B90nD1jLwlEFVvcTPbtFePk4Bo28b4
RXxcgHFeJ6HFeybLj7RYfifwXvVf+sS/OVD6GEyWcrD0iUrrIC6Pz1wJcfr+NoQR
8fa+7zYtbKaL1N4HD3/kO3GtPONvigpDs8URu9KaVmO8BirD1IAWuzgFBL0s9SzS
4foz4hKf4gg2I/6awy46AoCO7iX2II7ZtWDoLPtt9cemtOoUidfLhvZnND9tTSnl
q+sT+TqekDnGFudW6l2/tiXtMIlytbBXqCuIOvOmaur8kw5K1lUHBasn8JbyzyMM
eJv2SlNIh2PbPyuTyv+rG+TjXsMdnybhxe/sRtlgD7pRUR2v3BRSgQMwHlbYyqTu
zHDrCc2N0B4IKoImnHOMon7I8V1xFdsQYwFFNqozIm790fdJeU97xwpfk/T79h24
JBGKqYff1DdAl7ZKfaotlz/8betuNkgtWs/IY0BRwc59dNanAtpZCwYj0xEIeAfw
0Jylm3gXfK13p8SkPlScMVuwYWoj/4XsqtkJz1SP8CvwlqA5swZjLklbAIPOqIZ3
QumI1BWrCFsKoY8W08eoRSaSBxmla6hv7FGQFqpDgAT55tIot2L4f+wS/vgeE5/a
qLkAXQsVmfrbQmMy8XaRmrGCKW8vsHTioGfhMTkeohCBDrmGaalZWF5FS0ZYi4/d
1er7RFMylueSQ2eOHOm7iOMK2zxYylD0wRrwI5MCCEEE0Z7VfDywEbxcYhyCbCZ9
oXkIu1I25aKUfLgM+2UaEdRYCiIRTXtR6HZWdbrM2L0joe+dXgjzmp5t3TonlnmP
bC1v6ZGWH9CS5bQHaih8Ehd3MCXfzhovbUUH+lzTZDiv5LigSdigDLZcdmkqTGbh
3zFv6+pJDDAqvRtJBNjvc2myTJvFa5oRRvVs716i7kGtuRinuKqo1u1UdjYOJAVO
tPxkKzd7spE4Q/1b/Pp67b4OHm7PXwymMA3Dk0daCHsiibAhQk7IDgpxOWfMCjm/
rJolGQ3I7XYVisWcBGGDOlYBUDaHfA2zheMglo9toaFGFbbSPhjgBMgTQIlvQ9uY
R1nbhAWwBFuXx0Rm4hP+0i0adR6E19eOaRB2LbRTipKY4GI6jEAVKWXTDVg5nq9Z
0n3gHSSAKdSjjTdPmvAJwBaLBc5w8nrSAZJP57FbROLZt/vB4406bhR4lP/KWjsS
d54EjxUC5Q9z2p6WSNNoZXdQ1hRugd7AdMrEFV2XwprvV/JoI6AtBDFckEKWEbdh
TM7BUDDzP86emVe5ykJ71qUtUC/6PnrdgEg6fe3TfLVDaT3rcNhM6QKEMtAHNm5P
bEAaUU1SQg9zFanpDNf1uZMrEfsdMenKR1flcWs4q7yNceOsyhWDXHMYo1lafXWQ
glQcRiUIzUKgiOu/nbn+7Oq7Qnec/3MG3MxRc7vyJi9Mv/oWgALsrHODj23u7/v7
hODDRrkWJIRPCsT/hhmzbMCCAZMm7VDQap1Xw/t8TFsBnK1XLIlX40XhBcCW8oxM
DqyIQPgczSWnFxaD2PCVWJsT1vMe2TVeziiPwu15CXPzLP806++vfmGl4ttOPQj/
upaXGML9EHs1Nw9olXhnVpqBcOLvoVDZADO/l/s2OKFVmEi1LiJXf+zHMIDdZ/u7
UpMY67npFqokugfj3fEy9mvooRMI8tb/rbJzqwry4kksJO93bGEt2CozC5M7fwEp
s+Z6+sOPsYLSnYGs2i3aHlaaEuygB8/Nw8A3SsIQKG97HdumsGfWI8j8MjLax6Ir
4ErFo3BoH3n5FARDG0ygGIHPTd7UZiO1GOJmqBSeA/F5ycfs0g+f3p1aU+wPZ7Fp
LooYd/jfzDm8kDFXRdtBqMYEoLhDZmRJsvBc+424Tlf3cBqMR8/T/pLbjoVGcu8Q
har4yfIrh+txZXHl+ja2wOvHfMSeeulhy51i+1K/kQtbcO+78j8KlpdMf2S+RVGr
GF2R7YBdw2LG4x/gsUICHWfwabFPBWroD9FJhN7aKIB/ym5nIqVRYp/IN85ogiRP
hEizUEln5xBGCEvq435uBfPDFLnJqHgw7tWjh7SbwXky5BtqDVtKDqo+Fr57SJMW
oTAQa40pV8Nxdg7QQFc2DZ4np9jzYZypReDth+Op0FEOfdyiGYiBIEbDs1zl/Hk7
O2GgNN+AS3F8pi+ylpQUMC3p8scVsJsDBOLc96LBtLxnPN/ttQtc8Y+0HZRpffUV
8rAgFe+oiwihVUIr3eZSLIRoWAnQkjlH9qyxRVF6KPJeEjTueKAAAi5+Nnwi4/ZI
AHb/NxshD5KAUcA2kzCKJWoaiYGVtaELNx4MBES5ZIGx9a1vkoCX+E/uruiv+R5+
/y4/KCTEEHlEq+A5FQ4WmRXQ5t07Ow39PfbO3vZd5DPDvIq/DExmm3fQo4tx1MST
PKk6qeVfgDvZNTKDO8EDwH2GWtAuBd1PBqbYdzv7KhXWSNKtyCPDaVbEfvgFXp0c
+ZSDuRcBY6P+5fVbNtxGa8yDD1SChALnNwSkJHsCtQp7GsaKQ2fWTcx/r9nBSWiq
6lv0VqegslV+bV9UFw2+VR0ZEefXnNIIHunF6xodNtJkVRNqh2bpE4d9Ryr7tXa/
+U4i3JixFlwIKLAGHycHIrzrMhsDjMW9Kujh4leCrwhrojnyvDtVMDNvFJggLznQ
NvLyBTH8ULR2KNawHGg91Jo9+Q2YqiKadr59tWuvRJCy2uZSEDBP392QdstbGvMp
pGls3M1boaDyLTJtR+uVzuQgvFF0xmC1kIFKe60PXT53namXCuXntx0Ks2dpnhlw
JM7O7TfzS2n3BedXjSGASxByDAbl3nF6RDikDNAX5BpvlrF7tfsGl1CVaoWMupv/
NPYlKiQCDtKWDs6tutO/i6G8gcqcPW94w74GCuyp0c3hcsCAM+cSH3Rcd20ZTApF
oWVqcgw0BNTTKTjk4sSlWvgOQRGJGVLYYkaUpZ3dLzhg1FNaUVFXU9Z2emIG815N
fv3PqjS9rEIk5mLQlcUE8s2L8TnhXOVUIPIcEImIuUYZXaSAN6V0Yoa6hNXhen/m
aNe0ErF3P3AelUm+MQEtUyyfFsgg4Pnxn5A82nT7p8JnVQgKAn6KESJbJ7Xr7ORT
BuMuGAFMQXu5vhly6XLMGkyL9WbMoIxna5YtVDr4SnGp1Rxk7A7EYNTJ/MDn3iY3
hpZlCizCvJY9Kuk7sZEm8hchUj2KJxS/Xbgu1E6GyYPW57KQwZUR3ciY1oioFsnW
YZkinxy8puqxrQ65eH4W85v7D2JN1HO8YjslZvwVIiswD8XX5vv0TO7Z+ag3GXFE
BIaKDjS0PQ4rAoziYsNCttMI0ATrpfEHJGVQ7bmYLAPV5AUTf1aaZj8dH8URac0m
tbUliP4kMsdNGeTt+yjJE/aAcGlnAckgt6w9YGnewrpJBreaSHMQQUwt5719nX7b
L+7QYv9zD6ZWQBGE32x2xAxIHx+M2XUOVi9KS3OpalmN0jdl7gLAXL2qYmeOhFVX
YsMeTEpPBDSyq6hWrxF+GfwGG1Qs3wwKSc7IpVDInQxHJ73K8hks8lI/msRFiYft
fTSdrVOIui/akD/kTCxbrWAIF0wQCIX1zuvX1toWFW7TT13VypZuM0yNVzTprh+3
FyFaho4lVfXUjfs4E1meB67ScBcCK2OpgmNFSPiT+YL0TWxtVo5wB2QL3QbEmKZy
ZDrWSC/9oWcyscgUSmS1F/kS6Vvcr0vYxqrNafYhbcet8n3ncMWexUu7jSmGO1ld
SL7LZNB0NMxgvFqqppLLf5V/0ssEof/oD5x8p9lS/zcMh/5EqDLbhx6Ee6utGfAP
oIGhme0mA2g/JkSfs7vVfT7HNaiZvrhn/vuZuWPKYdAzCtfcfux+iWd+Zb+9Er3D
a9eKccu7JS8+IK8DS6XiabLpUsUWbFey6pMBaHmbp9Z2uOnPidtTPexqQzuWvNsD
BUfK4Hg3iLEA+Fvnzx/vctjMt0slekUgSzYImJ9InudPujW0ijKLE1J+qwyJItZe
vlg/h7XSUXTrWoGLI1wJIT8QKoCdLS9AA6FNNkpoT48cfNL117FK/+USZJen9F1C
Sw9IWqieiDxYCABthAy5OOmyJTqD9wFwHNr2Ok3WmQA43ohkov+p3sISHN8+NJmR
amDrEQ4qJZhsirTc1wKpCC9rB/MTF3lnRkSQh8kgQzLg/WCFsKELO00YjXHTZ1pC
hxKrMx+lpGZtasPcwgF+fs4Q92KSFoDXHDnQFE8LsIbSAY2lUpwYh9q8FWzpphb/
MbgioqYTPmej54zDvg+j+nD0fk1UE3QZix837p8p4LBzq7IzOvNUi+6/s8DgVERr
+AJRXjWKeU4A8fvowsR0dmCu9PwhQBNiiqV4pkD+g7uK74q05d1e8jw9DsbaWkwM
GwEAvDAeurAdVtFNWJ0hmFRTJNOWnozVjzMqzQEh9ZiHp+hWcu+GXs2KGPcTXlFh
fCiPX1/27+2tWX+peLlMUS3HcXs6OayxaNE50V70RIdz7hAJ11MxZiEPR8jkBYeL
oegI+DeNewjMLWj3l3e5BBOTUkUm0xVxyk3jlDf8XUJXGy4hpMnSFX6VnmKviTMr
5XacCLEa1lNIGYXfDdyqgoT0wTDymNKkCF/8ESOUH4QxgqVWU/ACKqWC9MuS3L7p
Q2/PdLT7SjQxSsy/MVyRCX62RFkhFzmtPzktkUVwXTJKwOzrNwmFDGaBEh8rlQVQ
vVq8TEAEimcysImoK/kGm8IGSC4OfC/1XY6djvMk1IuL75YSoP/R8c+KzT/zCAub
TigggANmGzUx03elC2wbLLqIpvKO2s95hSE8eElqRTC1eKBnhb4aaAZ8LPomsyb0
E8ZJMHt0q0cfr/esu+9XgKz6BrsEhBQTSiFmIURhI/HBTcW4drrWl8FQlY57lowl
gx6yfqeJwMj9no68iCb8+96F1UjM9y6iV0B9xIC7P6CyrhqR1PyrjrfYnGZerOw3
bgw1I0KG+sAnSX4dJ31QkK3xjmeMzRKmO2M/MsuiPay1ImYgtc8XDVsu6YTXyq1P
unmj71FhQPK5FftnQOQIj4OMM6tXe/XMkzRqmO7GpFDmiyW9f13Zfeso1kPzGS99
cPJHs27upWik3sDwvkloZbgk80gk4o20litd2Td8LWae6JD8woVl/5wKTh5GvfJV
alU4vQX4WynMNRByG/XF5QM8KIiSl1+8ikdrqMUQlJv1/dWdxjQe+qnGx2FXWFkV
QKx4jBAPn8Dmk5zYZbU7hFjoX6FecEWn7Ao6+I0IgXxbJCdpTsuno5IBmeQmArJI
MmnGzUr2Sw77KTfmb1sZxKanW5FohDS2JnasVuI/tgeLi38jTeOUw2BVz+GvmyYG
nUtrVcFkQnEC0nnzMTIcSEjSiAHbXMWobN7HhRgy9KASlskjgZyf/NU6CSARGdng
JdKuKjVPac+1C/8veXQ/XXQQdeCGL8cZgHRG7KaC9CUFzwXBc1nK6lDMZ2EJ3ALT
Y1cIUU+HX3/gOzAfDgNWicxO4yvtzlC0/ne53PSg/fKxiQdHlZ2ibvrzkJcdNO6G
2WRtxkXZsI5uqKM8VA17b/uKO7BDzDky+zYfrIbgLPw9paBpwzOa3nPR0yu8SK3e
lbVdfKt9PedHeJTclpKjtt/hFWq4KCf+OKSYwqXo6KmkwMLOdrDmCOZA5FeYCaBP
3JXqeDQyDi5ug9MZunM1e/tF4lURbyrIeJevzFXRetQuUs1SFSdM5bM/50R2rXig
uhkaxYw8/fbgQfVziPvCZ+/7LKCtnvN+cxrmlMIn93v006WcMI+p/wI/n67Bzer3
4RvJ0DeTHrDFsRxwHfvN5xOTZ/pXvLkJfIobCc1rc5wF1UY+0a5woPK+uV8Kng8+
sJcP53gUD2dwyyZWghH+P2LDPegezFGG0JgMV/aGvGboEBqYuUZctvqlnaeT2+BR
A93gf+LLdZ+PmyEE7OSF2TCrEVjqV4AWEiPxRKQv80TS6j5lBgUSRVo+Pyg5QZgg
cgTrn/DLeWIizjvnBxK4FQijs9MiFl2ks0yCvNDGQvQywy9+ZfD/MtPWVQnNHdjf
1z6PcDTwZbJG58hn/wxRWFFnes5RoTW1oc5sWRnT09cXTE2oT40xz4EHRgAayABe
odgAve2wk+tAa05ZNIU4PaOQuqQTVEhuLOSbDzUDSQ7jejTZmz+atSZqUNLErCPQ
ev2/U4UVPIvmOGsruCbdkYaX/rxrdvmOQ5YtSRM9weSX/e7ZIjpJHEhKbLmwbWP+
CFHCwfC4AkksIgRyhS+XgQyey9h+EBM9gLgp4H/WSjlSYqiw8MVAE+j0gJnD733j
at90tG3XAEeneAVT1dXjO1ITGm6zxzo0zS3U9MoE/b1Gb232pMQZNDno/cQEJ0/f
s1+WeSetYJA53H+EM3hgdUKVZHvBBdfkx+i+XvMsf4f4Q3+TDvsn6+DnJnrLRidt
sbtWv/RJP2HqQiidVb2KIZmvWUy9FgpzEeTQgX8JpIHyTycIhHUU0OZkCKeK6yeQ
w0HKgvAfSLuEoLSApxYzl+lhpio9GpXlM1ITM8/193bvaIuSrxCMoX9nfLrqdj6b
FC8kyfKts5aluUIRyDdLu83Fb+a4qssh+szbAPi5ChgpK9ZuwVpIdetpI+KeJtQE
mhq035xYtfcR2Nll9nFY15Raz8kQM0BPOB+mpda75EtVX5DS6gswuNl2Pehqk1E9
dV2jQgNXJVnO0z8ZFyZZd5co/1nfcFldFUp0ac8t0MtaC3aN0df+DSqC37z+X/MW
mxTKHVfct+W2qP52wkHcxqVYouVRFe4wHfz+OVKq72zsAjtOG7VpMtg0heC27ZAM
Qvzo1FBse+Qi0rFo/fqdvi+10SmWPVkevvcdf9heELNUJmPagaZKB3TQkzvm1Ic4
sSndqLXggPngIBz9hymSIfDbzh1gvYXvn5ZkVpPLbvQVgKcaoAK7GlCC+P/wspMq
9snH8C9pRCOrZmjXIuDeJeqokgCQ5vWlxQz7GCL2zUaLrGb5xKbjbo88Q7l33jGx
6UMKWIyWsaGRCrC7zImRuOlLBl97ZCXCTiT9xXk66PqwcjcZ/yfoWPNa2bgmkN/U
sONEBXT68EmqP80MvWZalTFj5AotW3VVEXWqnlfpUeuxHJMDwrbSXOkez4Cg6RJd
YqHjB4Gc3k5YfCIL1JUCL0Sa2DT4+OxoHrlH2TVL9RFG32I7BNU8fy0LzbW+6g8O
3jfMNqIDUeV9h3TBM0dobBaXE85F3PZtmgh+cGryJXiBb8BnsnaChX7ZJEIdC96e
EOzbf3xd/2r0kxPsv0NJuA==
`protect END_PROTECTED
