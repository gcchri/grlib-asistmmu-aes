`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CvkY1BiaT2hKlnTyp47TMpYAhSjTiBWz0ZLiWb0KQrS8zV7S4GTRx5r1tT0NyFn0
9nuHcv2P6YZQu6kapHahyo0eU3Sre4B2je/Ro941hj3VytkWgXPZ7P1mMLhBxyac
eZK9TZ9Q6Xtsu9He2rMUByX5wIl23f12rXcjEztzDkBs5M6egyCGf1QQofMC2Pz3
TrXngaiqedZUnoxZnTj82+SNCG8lzhR9z4sCo+PFvQOAe3CkdDOkUgiGtmv6uANv
ecwmIkWAlDLpCiCjZJI25RV94jm7RNJi8U5op2SEPZ1x+PE7CwvvOSlFtq1FCekS
tEOh8eFJPNXgaF5H/ebe4pFD9lxCMFpLho581pwXHrTZoRhAXI2bxFOGRPcisvHS
`protect END_PROTECTED
