`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9i0alnCdi6RORaZbS9XH90593xF2eILdxnF9a8eWGSNcjXV3pnmRXR0xFAxhL1vu
RWY0CH83QB9def/7JhUSxS4FwkwHTP21KScQu7uETARLfLQQOfPJI6n3ErHpwDR9
nNgnes+CRBVdpMRAY2g2XYHHn3M0C207KudFd0fKIImrjdDfUVKt8gWv4Gp1XQGb
+SugcE9MJUTsg/zdoalRMPmc7pIbvueY9IXaOg12ONWaE2Mu/fFcKvynfbLex/nW
Z9t9aF+1f3fZUNHc5dzWJPrbcc/GNt8/8QQ4DtwjCaQC+YSCUGLNJCJGsR8bEh1X
FN2RKVJX+DFzKc80PELXPmJtQDVRTwU8CufP1HHCU+EO2dR3FZP68SF/HFVCZ+06
mbbnJIg4WKmd6ArPE9Dpt6FeVLKX96LYQt0aMAWX4AvMvfbrqwHhMhq3kr4lIS0O
Z0BL8jSPtAwtG3TPx038ODzsno6LuSaRCt4XOX8wL9l54y/efSak901eLR6zKR9V
jreZZsqYA+CVCyaL8fkdlGKR0uOwtM/Un3YSL9YcwBAlv598yfNzMTehL1u/DZh+
nfyWINjQ3LHu0rzgaAEyVkx1o4u2njKmfMKMe0ur9hGTdLfMA6uk77tuGzHSP5db
yMiJ/x2PjXdLjHP3VXTnQ+bnXKDqOq8YFFlIWuDTJ64KdWRQOiqRgwuXb9tu+B9h
+OOxMZLqquhDss8idYztiURUQSu+tfr1KShJgpla9W/8yKU7au7KQBsZCiBB18aS
8xedGYjvLUlPGU4f2N9gmbXPB4q++UiHCG8azOsPH1VkAZaoSjwKVbTX3ubJvKCw
dXjzpXlMuzlQUDwMf2WX+gvbfWnH5fI3iqwWfGUiQMx6zKJlYMv6UAM/8BfqQDYj
1t8MkMF9a/agdWQzKC9IpoPtFblvVJnlbD91AMA1zZczqVosckvvORjG1Za3PmXP
KFCq8yOGawZdxMt7KuTyUH7szJeWzrNjUDCHplttmzqF7sJyPjiHjaMURIEjpTAq
xyMKBKQ2Xz4jZV27nJYpL2WAlfBQPFobMeu5vLF86S4KAqC5lC/3gurLa1CWhHmd
oVSeuSDER+lCwFGHuZMQiOOMIVk5RrfyJ7ArOp2f//TUsnoahNQWYM4970/H79Sn
IPXUsT/JdvHFwbOz4XvR6NEsLnmtUXlgBNMbPEYXhhE/6kPPOmoukJtdoMWDwmOa
QQ96uMxrNDTpF7TH6OolUClCPpizd4ZD8rq0QGLPMf4=
`protect END_PROTECTED
