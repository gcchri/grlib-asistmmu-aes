`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uLT4iGacTsjUlsarsQaeUCOr2zAkOIK4q5Hja6gZgZ9CetE78fXXpoLU9kEkMSxp
OR7xPeNsIA1Vb9qfJnZkfkCls6mm1mN3jii+oxsoh53HO1DZxADJVKn2XLvcObcc
U9pp5WU9VGBulzUyw4ssfVL39TE3NLqYxHsooYac3QOHziWCUudhTpS8Ho0GmaZp
IDoy2ZMZ5cp5iphK0ryC5rrliL+vPVc8bwQxH78nlIbN2XZXtHQNR4h44/qIocPU
aAPGhemfdkA3MXF9L3qm6K2z/C7srTuGbQagJq1lXdWJhfsKy7lZF8fBCTKMgx1a
QoblRZTURwpSnvA+XjZZxbTNZyjOxyjZm0PGqUlVLLyiGbmSWVlhQxzlh53ejwhh
Sl3c8QhnNnYB49jZjArscoyPcAyQLAGNOiz1MoxuZN//YST7u8OwsMQOipvhpWeM
5YgSQXuIM39DS0hPz4eJ7o1UcfVIai/nazx/KaKWQf/3ExYdl0yV2AYhy0dQt1W/
J/hKO/hIVXz2CFJnp/IM0A/zYVC6x5AbuAJJYW7nN0QXqUgO0R6FZ4CC7p+dOEnW
RMBMi3HQrdcRYc1wy83h3ZuJgWGyNRNDChvvLParRbL/3tIFVvIa45QzJvUqN5Dx
tLLvBedGDPvZp5Ldf4riEAURDbOMfvDH5u1+lY9Cr3HJsOJNQqIgMaHJnRvJ3tCu
CejCEcCXRbWtp+N23MkQKtj1lUBjaGjeygLIm653156HZi/taOdVYVq6ZvdkFi0k
zryjJ6FK3pcoFYpzBJ23md1d+XH6Okt3VQsmG84a4eszKN6sGmS2EO8ZnUdXvbXu
2HI3oNJn/+cjB1YQe4cE5lS1kFAR1kyVHkPnOD4ZjKHeHprHR9LtzP7DUpi3qB5s
Hojg2RS4U6nmZX0RyQ+IBlgHcgrz61LncQNeCij+E0x95+qjsb/RQZ2B3fuhqZpQ
`protect END_PROTECTED
