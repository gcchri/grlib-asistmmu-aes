`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y4S0A+N8ATlzSdJhbc3Ehbt72vIDjrnOgPRB/KQ2zCjCzCEtET7f/lXOTmVj2/Lq
UzW5+vVHJrKtjcYenf1L5a4SQV0rI10VMHu8/OjeazeymalhyVRAiQX/c3sZXHMT
PUDiph91n+/Br2PMHff8kp9ERw6i24pbzm9xDcrrnoeG4KofkR+Klth3PnhOeG80
5bVxPg0X0rnhfA5Ljv7zlF+FD1nEPHjR4hG/9B/ynVnYkWp9vv+pkMB4bBzR3TLj
mW4ZBcqFxDhGXukoUexteNleOnHu3s1CAUcV4W3IuDW0J9nfO1cWwGJueOcIME2z
JKDX2Ys0yQ2zYG6bXFFXb0YBBfp2mL2V3J+cscCqa3NJ/lO/lBO7Mp60+TCLqHmn
8v/ISboY3b+le8kfyo7vH63+yPKO3puglGxgdUhcQ5WVAufJPqcOQKXI9z9rrh12
`protect END_PROTECTED
