`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UHrwNg2vvYUEXnQER2RSpVGZhZJZZ1bfnvSDpl5taCMwj1ZWZFb6CoxUG/B1er2Q
PSqMbF1w+58mxZdFmn7eM+EZFfDzjTC/OMBEEIZAena8AfsmHfHlM7zIrAV+0h23
3CdqZayXnKoTs3A6SyN9KSYtfAOErN7J7giCjHJjzCsmbRm5tvnASH2vupGDx+Os
O82TakbC05R3W2RvGePeY+1AquVH8HjBkWqMdKooq5S/3GRzvUjqsTzu8dDteMW6
HRNNU9kLhQthEC4435Eviuuw0v4hvvreUV2/mAYIdDBJa7uWSjboBQXMbNxwPDkE
lEE0cbasWYeXF/1ns8p4r8RgXQhy5Rg8JOdt1JlHdQDZsc1E/WKp5kU6GPT2Balv
hr8Xmi1LanK7zkLF6uyDVDlAgqxtQZkTCNojCcjsn6BryfylHAozAomwjXIuzcGm
agarguDhA3t7hlbqXS44s04yohX2mPRGI91VsLBIHqziNm/4r5gLKlY3/rpIVVIl
TE7Z4CqsPGnOTpA68AnR+NgzmuhHU84A1GT1xOcsZbZeu0wkW9N0oM9W0B/zpx+D
95kNbbL0vp+35shmPWAYyu5D8Vr7t7lcT10xbOow94W/WrjdaSJ256tFyPzijd3N
ldDL8uc7abIuVHODJrixnN5PeKzTUIMosAmu7ujMLrEOQsVWqsyWsRv5qTxMkduh
ScHUoNjcYfR4BR7g4dJrGGD5fIzusN7etWZM05HE+qsr95nQMEtdWzOaAoYDSWvo
xrR7gVknjoFtUDlv5ORbjM9xiPzx3DcmTGGYQ5vkjEY92jEsP/9SxBgVn9Dko7ZX
noOXsXxRAjM4flgKBvGxkVpukn3GWOYidG4movmM+AB+Em7mtyYO/aECRfzgO+TA
IXrt1/70EHTIh8vNW4Tjkw==
`protect END_PROTECTED
