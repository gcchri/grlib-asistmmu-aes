`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xbB9Kz1mdD6tlL6WXrfF1nDZUHvdrm/g/rTisf4PQ5Bi3I0uZ+1Es+wfWjP21F+O
b2m+SKxWBBr1NFlYsTzLWkgjUK5oEO8P7Z59XXMsjygpgzJsfDK5PodzIV1rHb9O
gF+QkltCM6GFNtXxN6+V/bSPnPVGHrZba3wwAMSBSc8PQPkn4tJYv59hLfmp4jnK
JMdRykHwjEgW+eZHo6CB3oJcJbZysYDl/xbUacdqk7kYBA0/qgQim76v5RZ0pAAR
FidxoEvMW8aygmxml/r1OM7BdHesVusPeNrQr/4FHeoQ9oQ04X7Hg7GsqJ8fcecE
5xWOZqR7U9Je0KGCBNPz1yTykGY+JiDZ3mTbiinBRiPkt0orpjLKArJniWbkJtMv
U3fNFsaQ8C4K0pEToXr+0gruGJW0pVXwAG0w7npNmFcGT0EhSJ8t7DQQBC+u00OS
`protect END_PROTECTED
