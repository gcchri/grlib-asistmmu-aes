`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I925nlDNNxi0AmdoAHRQrJj3Bxhz+45ztXJthj5bA8qnD7ATalL18JCeGP8c85SG
LIXs/a5CRNnp9i6yYMwxRslwapJFSOXR+unAeMtiM8Mw/1K/HxGOHuhh5iW23byB
9Yx6B4jMcq4vz1fl8Lceif2WyParqD8R9c2NkhwID3YawRhtmMAwz5jF1sxcfmpr
BADvHVGPuaHplk8wtkj85VVNjXTngnj1u616kZxRspS6b/qh75hFDBJdY4emL92Q
R+s5SIZ2ECgR/tDRYab1k1IFQ1gcKjMjJa37kFW+4OAt94CZ92BN/58P94rBLAIN
XfsbKOWaZ2sNIrIQa/tcI/EDnEUp2ap4jQObI1aSoIxQfGRYgIEoCpLAFsn2qRTM
PXTiDpzzc7FWqC6+KMe5cxaD5Z7DIxq42qg/dTKkGOcV3SuJBqRNpeffKvY1nsJe
`protect END_PROTECTED
