`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GIHPTgpHx14q8VFsT4/EH3iBJOt7F/XXmhwhfEOBw+FNAtJJ0xlTu8aA4EQkR6Ra
+jBmIqb63Hkao9M5AYyZZS1T2tOcICE+8Rl1mS1BWSNToUdzuBxRZ7Fshf7H+XxC
M9qs/lU9vUfayNjBlYTPnhHuKt1GsKstMORzCcJvr/bkr1AL1WFeVZs/8GJ1970N
gtgghVs9t3IUCoRAHMLPEcJqhi8ec7Oq+wfWJAZBzU2V9qoON1ddbEr3cYKkUBy0
LMRrJDxsHlVq0+HOM3+Up3DLAglbviemCIA3TqrtZDXaEBFg8uIxm/ubrhZ72ePG
bF9tvDYFFxkeheFK7suPJrYY9300TvoaDPtrBvEaVlLmPSophtQOXNZ/4UJwnGRb
Ss6QJh6YWrOGHbNBhiIx2SXex8W+PTQQt9w/qDOQ0Dfe0YxyikcO+Yx8pNuVCClV
`protect END_PROTECTED
