`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+1GRZQ93muZn9kMUxIDTGZhNG4WWXLlCrw7J5FaJHnBlaCyY9becwNDzTeDd1BdW
B+FyW+VVFkMgPq28FdfKAK6D1Qx5MWK31ZzCVb1AucPyO55RBgS45K81ozFWjokU
8ZSe+J1KH31i+rRZobPqmmClYP1bQ21ZyLHL0edgYQyjzDcxlMdfPTZdcAZIM05d
fOgSnkgxeQ6KpUCrU6Jw/eadqWctixkFsETPaKtaEpJv3CqCgyvHwy4358w5+zmT
UZwMk5OkrwconoszBTGy37BLFj1J3X2QEJJG2Nifq+Kjvdvr3+zLUnQ2k2OV7a//
yQzlse6n9OqLroF5BHsD5b1o56vjTyeF5MzHFzYTpxCSIqB4DcPFnqJMszUSWSPE
1QVZU7P1QdwDhERGDbAYFRLCoLhI3wr0w/gDskyR6Ufe0cPyNzx6KCqFDahHHt8n
fIAnQdje9D0WaiCVRAyrxex+kSLuLa22rrS8696r6Gf0Z+rxJJt18IAZhrdK1RqO
SrDHL6Rco9L3i3ouvhFEGNOoIh14cGi/mkWJkmh8wj54nSWOkTF4i/A8h1clvlfj
WGki3piZBzeHzRHl559wWs7H3nwm/VTpGsG//Dw7j7FIJKlkyhd2qtWJ5m/Tvyx6
nn/T9841XwffjaLKoQELuvIUvvtjXFvgAefjDGr8FIotoXObtNe7KWAKv8qfYBCg
VMscZexWRtjHc+DS40OSkOvrU/3A6IWGYWiZIXr4GAmHVJhNZ+htDweRd0M2EvN/
Wig+3OEPlnQtGElCfBGk0t60xzuvUUvR/oWo4Y45HlKXInRLnrMWUUZhn7qm8z/v
qX44bDG9pZylAVm3i6XUYp3l37K5Zhj3hwi1dyvjn72bUStzrayoRDvh7gPruRGN
LMEQ5kowtZQAjrqd2c6iSwPk/XbT4YITj42eh9zCDFCQQkSc2Rfdy92Fx2Uo3PHg
`protect END_PROTECTED
