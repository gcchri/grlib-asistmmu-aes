`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AzUooeNCBbDUjaSqesgpS+x4vXLfQssHYgN6s8KJhqaicreyg+EmrmP9+Eu87xbw
W4glO2CGy1fMiGVzWvSbmuqV2PJrdwvIejScBlpMY43MyS0z90oUs5gKSD355fD8
d/qwH1iyX4nYviJpRhOLJy5WfJjadCp2L0YBHW0q/ImRd6kVYLh8mzw6q+joOEX4
Kqioy+iTCJvD+idqDyse/bFXokQqRKeHYy/jLGk7KtYnXa/qLnqUEGA6B+GzlRGD
MGvrBQHPDTEaeBoMje8cJkkwWVL1+/eGsC0pWHWrjL8VIIckzaz9QECJ7FwJK51o
L54eB163WTFAha6FbcJxl6/jKH1Oxv7gYeQLDpjX/UsLBtpVc5CI9WI3lP3hov6K
sn8ivF91479dqF0wBva7UPa71gdY2NjbjQUK/d2EFV9CCeULQ5Lc7i18dHKd/d5/
J0IvWiKkKlAABYBcQIY/y0W6PCQvYpyTiNKD2mOfKEF+boxNl+yCoYL90gQdlMHp
VIdkSqdLfTpNEg9eDKk4tLPtME0D/xhcZLg0Gqtw3+g56mKfNjYUBOwHHLEPCJEu
PCJ/jm9DWBeXKkF6lVb2vnuszu/Hb97fr9UUdgznF93cCLB3TugimbzqUwGeA39E
nCqBY5a0vLGo0sB/60ONHVS/ctMauWSlgLTv3LDBdQeum/S+5cysBNfFLtRTcZvm
GoqeRHyILOemNycH+O6fKox7xrIvQ2DtxSMAyJBcOt8IVOjgENUJ3HGQa8lDA87K
sjCPCwdqgzddHFQJhMOVZlFL9uRyHcDD3mBU8VU5EMuUoTNEdIvrG3Deavi9aPn7
2VuaJcsuyBHi7TfE7oEvjUPFhayw6L5gG2qL2iF0hNw+nOxrlkfrwo7x0EmDgDiO
EsT7lE5YKWiav4fQo+1F+rIjkRzmfGJ0aIKG2t6X8odNPBITidhJ5ysKMeJQDgkE
8EheApY2Cf5+JTrOJua7J0dNaxkXFg2ezgULK4rPDQY=
`protect END_PROTECTED
