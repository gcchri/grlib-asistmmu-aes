`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UovAToeUy54a6IY+gF6mxjbhX8uGKB3FLGMMWOlDxOvhMUbzAHGoeVLX7w0mvfrq
xbkp4mNc/hAUfxTo2Acuui6nVqaMJhb9QEyq0jLVidluBC9KhEU2lX6S0yhXHGWL
JAmGG4baibsVu/fVQjalGyLVO5ela4tQLHICOIY7QEcx3soQHLDgJ0HJMMTsS0QQ
31dWzJjFtvyXW2mw4w+uDawrPM+y7tbHseQypw4rmRgeE4sgAp7fPvxqfarPoiZO
RBbtbPid4uEMxM9dJX09apbSsJvq8+h72DWJMMttC/o5bGM3tFx/4KKEmRs9WRP5
frMnAxHRga78elJyYjWJnb9R2sA7ZtYrf3p6jOPB75x7ji0K57W/jwxYqMTYfNXy
RKrbFF7BsykYN04wNBUAFAmit8zpHbd6yIMoOdFyo4BwU5A4G5gBIyh4prnoA+MU
Two5tGxjkY8hFhpGLI/VHtcYfYG0ULHHrQF+zQ58H9OLlmP/AiDbHwyWdpRrLmfU
hGx14ypyCCY2Pj79faIiOECDcXXhWportntTLHK511XW0PSafQJkFYLMHPXDPtrE
X80yr3L8xt8RnvUI9xdcSyb4l9w0bhkk2kgy5Q3JDdONHh/IO8xZk2QfCh5zYP+6
HqYUEtca32PW928fViIrCkhGlh4vhGd5/cN0OnHJHGjuudeYXTj9DRNYkoauf/9T
Fi6FDXq1HeiPOSf830Rcfm9I1RPhpzf199S6fYlwMk3u05M7Aub6KE/kaWRgcOdG
xRVjJQlcuS2jO6JP1ezziLE1PpdrmODVb2uzIiAbMQcQO3NHGsfRY1VjjXeTq/ht
yGP50QbQ+Fm02FurYP/isWql4PWRjb8Vc/MSASY/wXgxLSxjJtWmb4Hu3jBzUhNV
2jtpyPRwt/yMfhDDXnV8p0CfqpnvlmYqmW547zqV6Dv4yss4D9xTgmVtJi4DZO6R
EfZMwZ/kFjpyLILd3IUOn9L8tYHMWtVKpR2rTCwqOpA=
`protect END_PROTECTED
