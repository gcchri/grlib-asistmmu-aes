`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
epo8H9UuNw4KqEGg18ieFS1zYqgPdpj/jbMeRmePJxOPAZLHuy9bVS0jQDL1edW/
fI26Fpxzet0m8Ljo/2GCt80SA76CpfjJU1tcQ/+Kp0TpnqYPt4QUHFrHGizVktM4
9MzEGKbrUeeKcRAGNK8lSRFpLeRcEnJNXp+2yW3T2JuDT0BoueFFNh7Lm46M2xV3
9qA11lNYXnXmk9agWnuuRbaNXyrM97g6GIohWQg2w9Ux0XjJKavyq1dt8s5AYaib
tFvt6wfv4uUZhijXrVu8tyvADCmcifz6xxsaSfIcohQkokcWxNb1zZojm7B44ZD9
wkn8VH3WqNILJVrr3LY4WX/qZJYAI8L8/f1iHXPIuz8=
`protect END_PROTECTED
