`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RNUDgK7bmXtqDQte5iLmZIJBqvMy/wpKwjPNsmiUlkSgQ/RxL/IWJzQCYUGreEvp
3mtEKg7y5mLcCH/Pc1QfTW4Gna4C+XY9TT9lUTGVeBEaYn8CBcJh+uXFZKbAoYdC
fyFb38hn/CdAt2hccx5uFUrf5cwfbCcuh096gL3Oh4r91FkdQcwJaXCh/j5KhVah
pzYPnhO1StH+12zFjVjsAqirjr5K5QCC2+wnY7hfgh6jS4f9jEk64DoDTzLslL8U
l3yl06oDVtmnUMU2UdNFqPKQzCAxCqT/vVlpjrhP/NMAP5FoZFMK5h2QaXomjqzE
pDPqPFOiyAOXqf8FVaUtyFO0En8GoNDPBTLLQvL597YEfv++iH3ehv7kRGjF9ISP
l9eICD2PeZnJdlSCHKA0/Whc2jCjYPTokoVtB/ENC4UvqCsYN0qSatH1a7/f4+zO
M9cDkd3qygbeLgtYGgYejCjyecdoufz7dZkV9qCxIBFPFQBAv0Etu5+IewIluadQ
`protect END_PROTECTED
