`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2fUKKNjy79TAz5pRO78+Q3Q7BMB8SogSLuhGQBZe3Nkm7N50yh/edpKOta+P83B+
yIKg3cY+TnqH0I2mtnTWRvA0BFtCsA4c3O0qFHhkKNEYsz0Q5ORFyW9PEwXPSzpU
9lBRINDDLqzlNsMf5xLs1ITRnPCvJKBVZNxs+wwRm4EsBd/lA5da43MqfSmpJSn0
EufpzK06ZpgaMDcnWfuQjl+DMtozt31fyFxv6/2MNSyzoQ9lB1vcwpq6/6FN48KS
FFSfZITwGdK/8i9+TNCTlRbY7WtP4pBcqMo3WTrHpfsHNldovpaB3y2PEqcOcM+4
1SlMBEml+hITHcubnmXEMJ9h9MMmMdlvwk+c/sZ5AGNM9ITBFaKV4lv4+aRHijiu
`protect END_PROTECTED
