`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d7RztHP+xfu3DJagIDfVDQYHyTkFCpzqkM/sA04TZSyxkq0qQ/GdpcS19NY41N9E
Z0eZCapW7RQqDtrrwCJJBg8SM6PaJM2VTKhVd4H29zOMuxr3uHnOuR8wU8J12izt
OTA5by/zFW7sDe/P3bKiyuae/BCTgoFjF3qQS8yYIxyMpwRQXCL8EhkxDoLW+Fqn
HJY4vx78WcOAksvHswoWzJ1d0Iupcs44E5QOsHTU6RqIzXRoRfBumm/oEwBzgFyL
oB6uqeW9N32X2mjoayiU70VrIDZ7r1XWuSSN544cbjuks4lphLlkjPKUUGCa95mT
rSicjPPfvGCzSVNNzmHLdzEcwFy5NkPOOfHDaLvUDgwtUFwWKip4Pnbs811bBAlb
MtWic5scDuf7rkkvgCX+4p7KAMtlYa636mG8bhAwMlpZX5Uh2d2oEAMJSFFYujeo
C8YVTuZ1FM+cqzxRTLch+c38J9DMTs8NZ3Jw9zVgNai4RC7JMOwhTfzN4JmmiEN1
z+vzQLC/gW8XF7aJWhBYQGb1TuCZ8EsoNxtYxe5qjhfN0UNzZQEcx3AInAPIk/eU
pntNx6Ixh4MY1ZvA+4X8LpTC2ZK+/5D4ZLRL/LN/9dQ=
`protect END_PROTECTED
