`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V6lxbLHVALg3hPIVY+Lwe73JyN3pUyNS9ZUk0B1We39UyZ0uCcpRgusisEbJsPbl
unamciHzP8eEGatldDabPs/KE81f4/DG3iG75ac48VJkI/k4KhThIBBSAU935aSR
un3GWZLdAd1kdRqhwX/sBh3pXrzLLbI42LRPV/Lwmqb77K6lwm771rQN6DqnaG2b
Rnak/4pW3FqfmR8iaYjn/Nb8NDoRSLTHDQcE0MLCBGIwosrQwciiyBMjpeYWCTfV
Vy7XU4XNP2JB4SmeqoYKTRbOi2BtmngRFtZqdwPfmkusmNnmLvsHfUB4HaHYiZsG
SaCTy/nX/qnh4BGpQ6zPM3YOd3lFVsYcEszinWTLNzOYojja0nsOe+3XUm/WzFac
+58UkddeQzBSl/jsfX+B+ds/u2DYTfd+AzXa0KvDpLNDkvl8KMzk6QjfA4qTYIQc
9DfZg8eYXOYfOEW9U+xN/wQ9OaTSP+cGYsdXeZbJeKU3cwrFc/jYkM3QBdOLkq9Y
ptGCTHSYl904cMvd3yblF3qrgtIRr7k9ETSZu3on4ICsBowXxRUL9Dnd56F+Z/zo
2PyQRdA/nW2NbyidvRw7azeep9+KrFYXC13UFiQs/RSuEayZIpYbIEqbbcV8A8dS
nCY2YVvCjSnKe67l/ke7FyA8EhrCsQze22QKeB3ZWS4=
`protect END_PROTECTED
