`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
axW1eIKCHucuoSDYd0wfHVcBFiKpX96+GFDCUz22s81G996E1wyQA41kD5OGV+LC
1rdPQIeH8QVvhgq6ANvZeUvTs7SU+D1D/6HfI/wXCE2iQnIbxADXh9LAltKbMm66
WDOccbchcZ8Z8a9NtW9tdjZpBbImzgc5/wNKl/MnLW/tDRk1CqvrHpIU4DDm/ZZ+
RLN/u0JY8VwLu8pxFw9CJ+sFeKFeleVy62FzsvW2C7XOCeOe/UjOB3aq5zfsY3av
YCgmS7MhQgs1ZMtX0K0TR6hS973Yu6exjkEukrSnzqxQfVwOQ+mS0VBHOJLw23cu
VhUZZeT2le/Nz5kIVdkZ9WbCbLFld7azPlKQ+IWQaKvMVVr94UsaspBkXiQjLzU8
oqpqqlnbs9qWr2Bf+NxkC9Gh0UJCbfXeMQ51KfBTk/LVJE3qNfptnEl60zwzwW8i
ZK5hpiGCxrD5+58Rs8upBUluMevNJwpAxuEdkVOAmgUAVP0OJs1xF4wrc9dYpmjt
AvXP2oDceTBWbhpMiE4atIehBGajZZkVM33FexAU0w6H6+XtDCLjSErSliiKZBWM
qEcrHLiyEbVpt27YQ4XzSPh9Rs/cEfXKMoxIjLf/gYIHFxxV6gkwu+bXvdHDbLwi
NEJo0itc51YZylvO/9JkjCaRfinOw4B7Yi3sdMVKwARF341P/vMf0CCoctCrYAoe
lcVJIE7ufrhg1yG4hWSWJVjXj8eXIh6nNFNbwAEYJ3rkf3zhCENeg//sw91Zrt7e
ibpaPjz/T9tp029kquN1D+dM0GIdx8ios8lBtsUY8Y1uG1GHYXO9gWVpjLVdX/na
aOO+P9tJdICaeUvXLrEXthYGhD3IupEW3ZWkKO/g/6JYa9RUtO6ELG3ouws899st
t0sbtQ727bphZg87AXBKh2G9rBl9tGQyWREktXARjFlgTq324rhrJTUgxKRe5ax9
/dR+NRwNEhuGZaahmOWm2YrtlvVS6B83/7h9Utsp7ZgShl4Ipgq0XLwAIjM0ONXx
zz4Slv8dC7pNiqCD8Jn6v08ff9YECqHFJOLCoY1yZCsa5qXGnRsY/i/QZnuTTwts
5DEC8sHOCS8uD/XdRepoRhA+9ONgnZiEQkBIE4+JPJIIVv/3QA/ggjTTiRDrbzYI
BbutIVgtMqBxJrDzbpfXcz1mutb/6YiUhLP2PIfiKMEnIABmro9sn0jjDPHq9TK3
eN9DQ9Ep8tI997uOLIiJniCWds+Sxn5GKbT9mCU09bJQVYSG5m2XgAz801d1/dlW
QBxLzs4VCltC9HhI1IQSHjWkrGBw0bFFiGYDIT6NQV9hR0AZnmnDfJ5ME9YFy+Bf
Uhq87inIIXuUZrOjLZLEByOlcOi3JV1x5SsKUFQRHqjmKVFKB+3IVGmIoXSn10w5
WkFZN1TEX9AcTMj4j3duXsPQpwgi+M7YwYrnxwEzzZUh8gfNyX31WyLSkktjobzy
SYWiveijDn/MNPc6Bt8Segg7J5B9ldambQlKlkv8TIGgFW2VAa09TJIEUkv6961g
lQKgqSdkiuvVlPFMQBBUTcuwPEQ/nBsPwwB4/Z3fKq+4kfp1Qe/RaK9HAPh/hbyc
fTrCSzg9MDmKtMs0nS8abRfhexMLtdSY3dVZB5RE8Pm/9V9Dr5CKHHf8xPpCmHpf
WzlJAlVIFvPrZdUDahBZStNpTUgD+UTCFDx/sBW9kmLXqNdigNfD5YjPbW0n7F4W
RqBjVHQ2LXZfK2dSch+rthE02jiDIbWYvahxI30pGOWbecbZl8ItjaHJpGenmjlu
hUFBXCJDMdZ8qAkZJmwn69lYBZXMWr/RrFfXGlK6U2O9CyZUwjosZRaP+TpWsu/6
7uFE+qzC88WZdfKQrPmFRPQxEwvn5PZjz3f4HMbbJgNo66VUT0C6aikzlIhA0pVm
XyXn2R/xoO7QjS7blZJviRkvv+rpm29DKLJlqZw2bILVU2EEraDoRzTIQjNzFyFF
SfjmyKJAII62E7L8Do6O4FPXJBMhLnwupS0yeh2SP3iBFLrZHckFJ2XR5eD9Yhb9
5TlWMEL+VX1CFa32Qf09h/kZLyBYK3sp1HQ/EdM0C1UTJ/0RltzsOYMe70k0/UFA
0gCwOtz2ZuVpG1feaw9wvIqsdWdYX4KKzYbEdVQVL+kTEVXAOU93+9+4KPPycfak
rQXBaw1E/fUBtSqbXlE+pa3Fe4yyVHaWfXZ7jq/ABRM=
`protect END_PROTECTED
