`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lq5PMpWKRPenLMiSqMRIsBfAAVbFeSjRq3WoblEwOKcoz08PGMubFXjpg3FS0ie0
oIHhxpifG5cKJchGbBBECo/GGVA3p1LkiL4W/rSKPFH/ihnAQ81Lqd9ougzilmUs
SPcbkyPujFq9QBTvwbg06CFfiLScdM3EzCB4bc3Tx3yOBE/JclMfOPkvyu7+O0y9
9I/pEBwYT4ZZimW4j/KQF3eh2ZhkRcGQWIRSDQ8wwXUgsJbf87yTblim6cmZtC0F
mkxuTYbl8vXY3PAJgCy3uM6/SwXgwwp0UMzAVARGDdg=
`protect END_PROTECTED
