`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GN54Eag527KzDIl2jprD/W6GxlAv5Tfd+vh+htjEzFLATHr5EyN+BOuSotFDwHLT
vmxaIvl5ljdtsoBZZA6SIJ/1H6cmHz4Y/o4BeetWnExB8hXMNuyCIRZy389ZUpJI
CJYJzpv4mwOTJYjO5DNYA2P998TzyFh/P/3GkeNf26fF73BIvGefKRxLR/HxGyNT
QcH0jMCqJMqeqYjFYClWXtPdzEJEGtYE3pCHpk204sIE013lxxxQG3CCBmBLRv2M
/vCKahMhE9IlMFC3CJDi7cEVJhmhvrIfHJdH7BxorvkMk20C4aZqXQtmuTGxye2w
4Ioe0y55X1dI7UnewVx6gOCcAf1JFuXXt5NjaMlfeBLO7qs5roPWFvcvQgStTTEi
rCoMy627/1P5EcXWQCPI/fqBmriTNfmNy38tEqggl8+j36770nHXdblzUU2TdxCj
3As+MX/tLOrTJ+khoLSvox5JBiZS7f1ESGwkVqKcTTjVZ8CiGSpjGjBl1UebpGlG
k7F6xG+Ng7/nEkWDBn9GkfpXARPgwACgod39W/HcfNlC2yTf9tUnA/l7Kvr3ydlb
spojlEEBC9bgHIC/6A9CLAjrBtmXfZ3fmx/6eMzPqwB69oVbc6hoQ4sziEfJ0MY5
V2L6JDvDaI/CzEoHmCq3jA==
`protect END_PROTECTED
