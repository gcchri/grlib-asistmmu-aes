`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rvg5MijXAUod5mCPB2EIMDocxOQG5OsDnhKnAkLMVe5tJyfaKZLYTK3su0/+P7RF
j5lDMdqAzAauQ2xRdzr2ghaZHXXnh/O9Ak4PLN8GwN+9+g1uAsz/jHUUXrvhFadO
o9ThRdRhQ531SHyTOjZHiz3MVBdKDtS1kVtTvjuOK+u9GXfUr7h16R7ZeI71LTf6
YQ6ULrCfMU2+DIvcx2sbwksa+v5lsnfj+EkiUk12Aj93R93iFp1a9D4E+26j/0fM
0kELZARBsqi1HR6dPYjZhimK7dE0D/6LoZFhkU86nYOc4RJDDC9eXMaKbudEA/BG
09eAgkOfx+PL56nZBW0Y++8ykALd6O43cHSr/AdxUmvm735YCqAJtIfKG+cwPgM0
TAN2ITFsOcxTDKoxOceS+0dmJVUpvzSBTpdvdYHwP3153/QENTXCNJFck6FSbBmt
HRPJzyWwAWuv1bh2jjuB7y9iRHVaZl0NLUf1PMH3+jp/kPW9v22UzsC7kz7hKRqj
`protect END_PROTECTED
