`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l7Y6b2YvxfZnSL3h3Mu8SrIaAMQ9b3oA9vWIc+zYUzWsI0Id14HfsbUB9tuqmYzZ
fLzbyXwc2d3gMjRc/M1LvRrL9d9Ua/bgvYyMsWrDrs3JGAi69KGu7srqY/C3lIdr
XZLoL6R4ULyDaIuAuGUfQfpcslfh06D6RLeTcvmdtiL9ydfpXvOLL5bED8ZlcXdw
YCX/r5iLNvty6J2zdBSCCanzHT9b3/W3DoXy0/k74LlIV1FgfudVaH0gdm/20IRh
wC7RD5Vi58nV5zx6rZUFt3hAKCeOR3C/p28oEZ61GF4azw1AeTmB92r8AYIydz2v
JKgtkZ2Up0bFzGAj/zwUv7+hKHcvNC95fplaj9+ZMhlfvMP5sA58/cF98HFMzmWt
ekT6hPEzpbyEcsHjQ2oX0lsSVbK4uBR78c0vqmnyqXc=
`protect END_PROTECTED
