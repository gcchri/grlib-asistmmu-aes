`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WFaulOGM8vDL1SA0AYlmqVlZl0nkitjNphpYRtxcg5OzTrgsepi4uQ9p/twBFmj3
geGxtalz5nzFwzeLturYQtkCLAHLfimmEpmtpIz9k1N3PEUzhLCa4dRrDI9Ibqq9
FsyY9aR9gWu8ZbLWMD/Y/5+CT4eGE0DSXFILRVQ4s0L7bQrevI48zeMJKzv8tlAM
4sRkfi3fDa3W+Q7Mj0/RgvcKOyPhptTn6W5cZJCvUCVjuvz2xf728tZCsTqBkxE6
SiP/5NehV5V4XM9wdcrzCWs+QuzpuoiCNMs2nKy+CxlHBu9B6ZMjhf1CdRx+zUqW
mHTnBqvlmhjEvqfNJB6VJp+dZb6eH1x2y/vu9ZPbFJapFdOY5ComhRA6JDaGZXKd
bR3RkHVexioUMz4XhthxGD8Ftf4bnC0a2xjSq+F2RvtfRQYZ2mmn1Tpf2pu8RMyM
EFH/S7YrsMf2OjtrAJ4ubh8Td59qPJ/63nLXLi3Q0PjRch2d5C9Lm2eleweLpDJA
nyahQsk+WclRPV792s3tc3+MwH2EtRFccJsopxrljiR0uHj1yTm9mWb5HzPqCJ3q
9zqhGhrzc1ViWZrcOdkXqg==
`protect END_PROTECTED
