`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wi6fyqZGSjrk2cIeo6ofWw/nY66c0CYVHE4kJxPQZX7eC7tqmGUnyQpURVOm7BzL
d7FX//lGFqh6ohGHTnACsaDbep1IMqaDNbU+6AFY/VeaZUIzZDmsEiuG6tdzXY4t
dmA4NRX6iLwq9fVTCvZwL389ZrXfh5pOgNc8zXzThuHebjpkMX61b/hOsvSjFPlm
wYETG2o9b0VMHSHZrZdtiSTk2okbLEFNR0Vjuk6k22OxNOZ9rvXQXqQdeTFjai/y
Qq67G6k5SVJ7LDiBkDAGUDj9hmk1sWBA+NrM0h9V9hYX8BGyVJBpuoor/E1Z/bl3
eSqRRr3S9fceZ6f/atR/rqYYpVc457+Wk7YFrC8e8hhNHhCv091BbrQp1FKgZ+c2
brDxJP7rquFPlNvY6iZlWk43MM8p/0/kNO6i9XXeNredlvujt54fFjN3aayq1z7P
bR2wwdJ+J6sCwD8PcS8jp2wT1HUDaG9nSmMeHlyhMlH09/gLhTf1NsrXy+unzGvz
Vi18td8u7j6N78g6X4znkRPCEy2NbTop3h5k1VogCdLFCh8T6BQ1zGmtZzlEQF9f
33YDO8WmWH8eMCXdpCiuBVhJf35xsodrR57sruQfz26glpXyBf9nImUZo1z201+f
zTw9fwQ6NibGvPNQCfpg2iTN3vsoTJ6s0TBLEbKPmo41WfBLTFM0zjWjoDe0Mljc
6bI+UC3T3tVVq7ieO4eb6G3e441gjGTTfDy+zfCW7tKuJTPtylEh3iidrttFJWh/
V4nZQAobqCFBwMVS0lSAJSxCHjCllp/d3cT5YBL1LexnLhbcpiTBaYAA0llO/Iu3
PH/ivciwSsDgAZpNJYVS22GcIm9X6w4tGUndGqqiHyF6E0e7uSBJKc19wpfJ77KL
Usd/6/250Zm2wj63F2Mtu0r+xOYTA1qFdJvAgrUeLG5NtsCnSPJ4XyZlP59pp9Hu
5uzg7egFkn/mM1BEsrSyu3KqHp80uoRhFwOSplgz5x1iTyq5fICs7FwYqkbwjzCa
icGizJaRb29pJleJGKel/MKXi2zxioHmKTlV6RLh9WTSzordBvvfgYa+2rAVCwYB
pbEACWAUmP1aSWt6CS6D3UQHkcxWSz5p+lO9kmQelWTGcCrR1O9VuItqGPO2LxA4
HuJPh5ki6bmqj7zvQPZVBp7295T33cwheZEfh0Yh9pQHn/vz8WniJEdQPP/FqWVZ
XT5IQ9ggeTTtxnxXeGe0ECxKVoui9wKUURmU013vg4XDUJweJcom/VH0E69Z5ILu
0JSLKZlwktGuj674X3lgkOdx+Tf5As/B2fHq3h92Wz2XjR+EQzfVjUfbI/8ojZZa
ucuZc0HGodTMqPipRR98jzWJhBpNe2YCS+OZJPc73fxSe2dhGI5JaVY5owaCK4VO
aFBh/OAQo9dC71bIK9LMa00h7wD9ET7iGpJNPv/bWV7En6svUL87cpmbqh4NZvqh
eFEvb4Etn4ivJJ7vethVBgqVc+WOOoSZMmgupx4qrhK4jBu1Ki4X6A0kz0LF1lmV
OtqI/DPHJSeQx2yuag/TSyqISwifjG+0m/iAHWHxoazuJH+728d8Tx6f3P98Xlgr
MlrP88KMbdPHt0yW6oLSkmrwwXgO6Y5d/f4Zq4K+qEtwr2khtinGMiihlbIq7+5n
ppkdMNN/rye8aw7eYYDorPoHY4ZanE5GAbjLdv4wegtiDtX991LDYUUlLExz3tT9
GEOLDvgCAsO/WN7puFsWhKXO+c5nE4Xw9GPNENzu4RcxSn5/KUy4Q0YGKpXmCbB7
qIqSjTTIisEDD1X56NXkQq/TuSiqTSQ2gFAXX8mlqEZ7U8TDhta7IDga1FS0bUty
ndiSvKo7Op34fh6uExYyc+gg0woMUEVS9GqnRXr9HFBVC7F6JTRx/+u4LuWhlpul
ZsVJ3f/cgYTGNbSqSFTCv9r7nMbbdUpjrg884sNlezolTcae1FhXb5q8di+EsxMJ
coniNPv9ZQ7WKc/dEBghz2obqcZ13hmv48xFUmP2VshkfCH23TP1LmeY0NJOOP90
nHwolrpokn0dX6J+kxVBj/KaN36f89NN1gNsUOKbjERkJEH+OWzBxQKNAS9eDtre
Na+YTZaLMpXc6NEfb8h44vIxf2qvmmN5FdToxDBSXXpLruubhP1hOzOfDBuoHwVT
u32vA4fmv4NRuemCSzl164bI8LEl8Jkd+4mPw1B06/y6qW/VLQtvFghQBmJXpm60
94zGpwE3AjV0Wz9V2wXRawe5mLB/xpZDnP7/tcWdNDgy1EUf2Qw/tRVocV7RhyGJ
Coc/8JLuFSvvSfYGX/mlGbKT8HYkiHfgL/zE+OnHODETZIlas8+4rq2nOibjeGzL
+as7EB9RamCFzV2HhYDAiscXuq6ic/83e6uUCMUyB1vyYkSaAyr26Dq6VSFbZk8K
ljBdfiX/BpBbJdS4JVQTljeySud2aqSZ/HFC/4Cwklt/NJoN8NfDF2eB7f7YTxBD
eI0Pd/2Jn+fP9/prnTDstzqkQ1wzvqvvmrbujdCldVotRzMTuQd1gDs8tdUsTPi/
tEbnY/DfAXYwKX73g+YXnm7dhgRxPvTc4oVs3iA2sQepSp0GU6fO8EhnIVSRRaPs
EvqNdhgfguOQe5q0D6SMl9ibAS/Cge4quT9Y5cWouWVA0y2Fdrum1iXZRlF9/TNU
H3Ro9iDFXceAfmufUUmYHoRXKmYafq+8Eglcv0UulKQsS6kHzWklwWDmEJAQGm8j
5XrS4zlFdm91lBZ2oeTsuV+gunBWkvoH0FeVUcf8BJutslfMCk5bBkmimox4Knte
XIMS5B4IdDerrFIHHOMddIY/MqFdkmv7Y3ci5iezJyJdn+lk4LSOliDTGU5OeRb4
gdpy02r8aPHHInB6yu89bm8Yundk+D9HzXbVjwrD0r4l00BTYyEh4PCve7Cw391M
bfcu2y2GiNhjaaRHEAuQscy7lzywYRDsuma5xLkdj+fkWYb0pJ6QuvlBOuk7aoK6
J2lf2JSw1r4Gkrz3J8DrT7AYbjXwR4MowBjWqRG+R4rGr9kTV51/r4oGhSW3yrVd
3ttA0i1TlG/GBDKtWYMrNFIdut+Ue1gOnNxgHlVTWyBQOVjFaY/8efUKurvyBTvI
LkNkpEvIdBzUagTBusC+LcK0Dj3UiW6pEd+dszfq9hSEKcgEI2ryIPC9T1cQjjDu
LZDrkAsLd4YqgRw373C4V3jf4+tc4U1/XAUfE6umYTvVbWk6gkTP1v06ZHtYguV0
Z1qiEu2kQnNIb/zp88ESP7vUD0UJRaSwaonjV7kV/XUc9K4Af4Pze1iFg/WWiY0B
kkp3GEdGDAA1yPV48pJr0/gcuxEWNxAtMXy+AppTmm73YfbkbxHqVzOVKYj2Q+IF
xRk6G/HmQd6JLlPHn4xYzJ/DNiHGliL63jGwfSYYZuB9lEpogfwr9hx9uF3drz93
oVdrWQ5ggqz4WBqPe2O1vP+0iP8NnSI8WmB3hDHomPTjb6BckJz2MBTQaIZrZOgY
PWOy/6cCx/j+uO5Q6WN8M3hNdcWDbJtwE92XFbVQai3GdHKRVhBgzbVdDmVV1MRG
sOsX7Eth/pIOGq1E3zEv1LvxRi3mutcUUZ8w8oYlRWYS1NCD+pWYcEtJE3Z/nAAT
9DsWUpG96I+JVZ4J4cozBoC0w8Oq6mmWvfDortcL+frxB4PShsrcq4D4b9TCP/bq
EN9UZWl9qSA6WNJdvChMTfYk54CG4WOcP5W6xoeraNqV1IAkCrWQ6LQS0vUc5oG3
vGzX1iVx9LGQrFXgeAmYBm+LL5XCH2dwK2QZjwsIqIK9WONczvUpMusID0Z3TdYK
m7PdkLUftarq8o6qRQr7FTTHjcf+wBAxN03EXMuRHBSvQCykhfKTXmtwONwAqAHw
0ajN3oziDWf8T0RdOFXwUVjA+QNf45qCwQ/loqdkhWqRvuI8WCVOGlSt6/J53tyB
496pBxljsnSbjJFWjFwoR4QWO+SeUB2yQgr2FlEm3EtUKH6AMq/e3XdbdO0XFOLe
uK9nTng/cwhbKngiPtsRvyKTTiwK8fgAMBXLPdwNwsmGl4y0lMCWFXMFRHiSan7J
4DiXWvCiz12M1GYR0Bk7qNauFaHAkd8mpe/MortVj8gKlMpvIYVN3mlM6ik3O3j/
33OkIAijF9j2sFX6YYFZN7A2HgPMhLaaqzmt/xrLCebKDn1UTxj8kIr8dsfGzc7V
MnwzEq3huKNrBxnMIglzfE+xNFW3jdDqKMoNWAeB7cRQCfx7Flc8ervw+vnou4mp
epu9YsMAkndheaQXYUOID6X/h6sEsbFiYv5+awyveKyKOhneb200WeuxZvF4LEGd
vOqJiEWWcfwYH/2EtGotacZJPofh84vndeR/HY/lQl7aV1a5jAuGg3Ru/EfLNwNq
EGnV2NB8gUb6GXBagAwKz9piEVa+R4aMj+vdbVZR5yhyaN8LTnoBDBY+swhyGkbs
EVzq4pdb+Lx/WnppRmMWmTTR59IU9rnstDdLcvVirEFXakHBTHsoAaej5R+Ve1cN
URgF50x4JtO10iXtlgu5r1OhAFSIK0DTgpnMwF5uGe1EM0Iis3c9AfVIVk51eupn
XWyDdL4IAzcgcpA8I2OjD3owWttlUgbWzAE/eElCgoRknvUgt7MYAv7ywigInNcm
33yh2FDN77Iihk85MOsXFn7DpPgRpvz4IMnQ5nufuPgcaI/anQyyr4sqHdSZoK7c
RVsJkTv5+i+XvOc6WvvcTCz/CQPbRXlc0RpamHXFjNzH0uZPxt+JpuYZTqM+HN+w
s0FA72rY4WGYaPBNxJ+qhWjiszClO+mUKvG5zc0gn1N3w8bcTyEkOJ5zMIeRd6zd
mYaZkRyJw5OGsDRxKfQs0yQEAulUAF6PPGL5n0ln0Nai3IcbjD62zlePCth/pmx3
6xykywaFcOwYboTYGEBqjx0Cpcpd/6nwt4+AQpfl4iOqnPU0p8o3RO/KFjLFanF/
VC7P0UZNL8S50LBsSI3wPGy3u2q7NS3uTfSBKBBitz/bgxd1fY5vqBj2VJMNcuDs
QRi7nAceXSXYRxtv7A8ZCS+jYrBiY8YU15XLh2zMdl3uz+1EkTVV/1AnlS7otc9T
ecxqODFHbzFKR3qEC7Xg6Z0B9jUX8zZj64l6c+3xIdcnCvKXT34q4nDO9QUMcIaH
TG+F1cosPB9I4PyVlTvM1aGZeDDDUGDKzCQmz9t0pN9hR3Kkp5dlA18Om4p046sR
IB7LSe77vbWlNbmU9xeFdrzE1gJiijgdMBFQqwqCoulkjmpeb15iAY2gj41yukk1
NeKbBow8zFhRX/1K45KiwLSK/A3gbfvex/HN2otTOKd4z0EPTLn4TWBe8O5ouM3u
pMCb2cUrhT7J36u3KpO6OTM+pIdDje3LNQs4J6nyjXxFC6LqNzgVdhrLtSLXjMn3
cHfCTITRng5FDUJLpp3ciD2wK9BAH45ATp+izHr5p0jf5zf7wI+obXi83ctCnE9H
2CGIydOSGydOjKqp8GsGGa47bS9xjAhhY97YWR5NAUVoAtlYjb/npqCcGxvFSnUU
YNLh8VTxnCJAI2lBIH01a+j/9KQVnGMe3yfJ2oKb4F4N8HPLrIQZdwB6Nfb2+EQr
n5ZCiAGb55FsAtQOGCmqGSUhpo2wvK+CZUN28YP2kriOl2s0dMxOZl7cNCvYcpli
m4MgHgT9XuTN0evJU+oQPx4BXFRFWm/gk2dsi0iARQEiASjnZrcv1VaQw2Oy3vGg
6BMMDWnUXtKM3ZhvNmwyWYBlM5yPLsAZEspdY0+VGd3UHplocj3U/1uGqv0HO31G
YgmFT2dURi1lMF7qldvBPb41pw0p6gtjMODYikoBOWDs2ix20sjZeC3ynr6PHqsl
w0IqY5SukVXUf8TfTM9S0+4GXcJIxSWz2lLib03Z5350+T9Q5Ibr8ajLxDyEiqw2
`protect END_PROTECTED
