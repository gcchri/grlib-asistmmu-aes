`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l06OoxZTkdyUbDgH0SR4CIt5Nd9UmbhRFJ/7n+H9A+m1iI1+YXpRDdG+oxnX3+i1
XPdurdOCjcwgVAY3Lqo8/89yZW/bJIShIRJbCPsle4XcVQ8QiafTstz9T2yXv7Zn
DqWEdlueCs5EXnByT+M1cbg1lxEUtKj/cadqPJdtCfaGZtNGmy14p/yIb3VCMP96
8pJO8HMdofL3lesVJMmKInWi1mr/HxWoT/vj2u42UgcS0q5HehxrgDZ0+AWgjh0B
Balhm99dvXTaFPlhOLgGQ4OPnyJ1QHMCDKyyMlfnaXw5lFyG5uqAA5HnR0JI7lkb
q+nUdqD11qoevZU54MShzwjBr6MNbY802AzauvR3ypdV9EMuZmN4p5gbp97ZMad4
84Htp8NQ3EndhUCRkT1AgpVLJuxWjF4/xr5GphPvBTw=
`protect END_PROTECTED
