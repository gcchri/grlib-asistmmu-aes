`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ehXNbjPV9k/JVm7D9bb4PQtl2/BkuKd68ddRo26Ir2joUB9V0ukeaedk80Hun2U3
5qduXGk0mwDlOXNF9L+cjTtdY4fQkR9kSbYsZcLv03i1NHk08aBsOH0F3oIO4HCg
5BeuUvcB/+dHEMQVC6qI9t/GdQ1XV6J4P1mHWK+sBqH9ha/DrthgYdE9VML4Zega
H7Tp8dTiobOCG28AWPJxeD5rX6zmf492T/GRvJphnP9MJtpgVc+zZoRqV0B2mCGD
+LQsj4MLmxNZVdwKW94JEsOs53c7rwPf1pyL3GRw9Xb1KyjpxUgOzl/Z/WhVcnS2
gITuY1Azkz3deQXKozVVa+pHK1Z2O32xjbIerXVyz/16mvXQrMiGUvIoGZFnRbJJ
T9Ague5LqaavSEkPJCov/1po3lPBcCYpSXNPbFrgmTw=
`protect END_PROTECTED
