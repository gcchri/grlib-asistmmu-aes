`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w7dzuVffhXu9j/3b74Q+3xperwKR6oEmwV/xLgeygd0tBnBD8W1cTv7qSiKp4rM2
fbl+KBEAhIeWDfZWlvaWce8625GPySSiLd4sviTBCPkWtMteNwOkz5k/eMadJ327
m+7MAGxVGyexiQy3zWAzDo1sWy5DC2+iwdGqAD3xn2+gSaXPAM5B4oj9B9xkP4bM
l4yWCGnidX1a78dzA7+8zuQlNUdBkc/SomLaf2JAxITDVJnL+/OnErggS7nvFawk
eWHlmCWK+xuZmYSDmIg6bQ==
`protect END_PROTECTED
