`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bNIprfozbd5lkzDtHWSYT3lrtU3XUPw5EpkxNU3XehaV5iEJ4pVSIEgbRc5Jaia7
nvEh6HSpvWKYcXODJb1fpgkGQuLKcFMtERlPHRaXyDeh3QRcUeTFwXu4wIRZ2jWB
DgahvOkEmYoQMAD5vnpKlQ0gzcuel1FBK//FZBI+NGm8MY6D8Ol6vIwN+2Exblx0
SjQUYvPlsCmQu3Sx5Z7p73Ta1qvLBJYyn9qRm3hlYgE6SPGMVmc7u9pJW6+dain2
s2W8VfeDRiXrXtg4B+LBow/CwyEBfKovsVMuP+lL2/otySdC8QAn+caAqFnXQseo
lyFJIj23bAsD/GOQ54GdK7PWa+PPwCt2p5wxbaC5B345pYZO7wgsRJOtDo+1Q/U3
JFb2z/SD8YCeuNo0eHINa0xSf4y8aeji9DvTxVLB+fk=
`protect END_PROTECTED
