`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JHd4MsH5NTgCjSTuL9QoXDVwabecCKWMPifD+l/XTjHhW0X/qf1qGhOdOrbgfAx0
559x674xvjLA/o/CZyPKZaHRovizCM2l+aUsnTAQDor8WBJ7zpaSasQ2OS8zT/XD
662BoYrbUmS0pzROA61Z6Y62ipgxqrAHDlIYNW2Mp9ruxkdBzyIkPAgT1qrqwVWC
aVZGrnNoOc53kVibaKD0xnrK9Vqa1YA6Qp91+wC8nk7OhFlAcp46iDa6ttmZwzaH
pJlzjJgygTsBFcWsCJ+YUYpazA0s/JtPuDZyh5eFmcMhxqm/6PnWmhgATdSx3aXl
XTv1Ul4uczBC48GCGxoynDWB1nzrOXZ3m1ln77x04xkyR+6Azo/0eZdpG5yDVlIz
SbRRPrsMeMDPHZC4PJucSNtr7bOHhQ/XGncYPVBbj/LLikHEwa1qryUXASJXaWhP
AcEUjJLP2rSHBfRZYCwi9E95JhpvU7NuHS5BeFqxSX+qEcc5SvGyH8+V+PrW1fuN
`protect END_PROTECTED
