`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yp8AnqjIR7eyHPnEnnTG1wFnVl1RzF9uhKfmymsXSBCKaMvINZeO4zRuEO58SQ4z
9QuyFzhBMAScCkeaK3G72hnWIDUABQERjvaHnWb1gHy+d9AXxmqNlNn4O0+Fs1ri
5XNWMopcpGeci74gWRaBRRoz+G0xcat1dZmIPb3uAm73d3h8Ogk2B7NUPNO8sFnn
HNKp1UybVJTVstrzxax6aqj2qM74uX78E9Y1LU6WbbGNM4vpjvwYoj95dUjTu5gV
2WAYvFoVBFjsjYg/7He3X3A2Fa1OxqgtMfg2IGnSGxSAb+UrR/OQ0Sdm6EeNbCun
BWaxXHT3WlihSvpKtxALj2Ooi9L8CeWsoUWj/0O/rotYq+diQ+eNqZUfgzo1U9MO
F7SLvziq5qk7AXqVrbX9JWyUhPCPPqCSzSUs3hlLVQstazbm5LD2rWQ8Zvcxrlsv
jVlWKCFqd8GyNu04I71wDKz8/bHdWWK5EBArZb/N4v4XrUmqQrjQ5fBuZ5giFu7g
whtlFy02FHeVY/jI7EfBITIGX4hqrn2gGfG0bV45ETxwfrqpHLD5APLPfWtZiem/
lYJI+zC9lJsSKiKnxflyL1acPc4CCvu9M/Enoeqm+knb4nc56g6PdXx/YnWwxl7p
3x9fKB+WIcdem3+/vXhZ5zVDyWgSRyoWB85N+u90cRT2QGKhO7SgwncfUCkKa9H2
xroRRW+LCcl78Qwi8E2omRpgdMiDoBn59iGgIgeY3d0yaOYIVmtp8vCtkPg2M7hr
5Sr5L20gkEGYDY9+JBz5oLb/WduPHvknGNuoGR2QbVR/ulRycWm15XTrKwlrGjC+
uHAx+Z2lur2eYEOQMu1hC6pKr50IWL72hzbslH0BotDkIK7Zc1sGvmXdwlPrBNeI
rF00/pENyMcO9VJwYVwJTE1JvGRIlUkyV6IWWFqbdpuy+azQ5BY1sI3v0PQy2H/6
yZUOfhtK9aJUjjyW8IRPMTy8d1wc22Du//sMObGd/++9Y9USKuqnMQ1/bI7nHbOe
54t9MAncWpv4LC276dFP5SKvaGSG/Vx/XHZN0lE4N7Yr2CmpFP5nKH5jOXJX7gzQ
17YJQdAoSP9KLbSzHRjBP0xMXO9S23wq7y2GLxsuAFGM1KvdDJ4Cdn7qRGS6I4fT
OZp92GkNvsep1ht4ZD1Ka0hwXsXPwMwZu/XDNBQTYU+55C9w+KDRZ9DtmOdp8WxF
cxbJlqrtNJ4YqldphNzPW3oRfsO3BC8HbJEX8N1mYjeGpjZ56IwH7CN3AuFrt7WW
ttBtbqa7eN5RO8RvOLr1UQC2Unlu/7ElQsmQfESGA+Jxu2SAzPSFrjLi93ylTiDb
I1mxEkr5UA7GMD3gObA7sS0TjLPAYKaBRorvTEdRrQH8OWzLrraR/7vwIHU4WRlG
ELogapiJ0/1hyO6WA9xVAqbauRrlzl+66wacw08CN/3YGVeGkpDplejOJL2rLsb8
Ju70JCe+q4siYpr/hG7aV4EvON13J1NmY9hYlDUkLmo+WpBiEhvFoi5GQt6RNcGu
kq2YKHVeRd2wB5Inr2Muf0EE3lzJG7qseTYqOlAq1Q+LbUtadkljQtesDtjBHKMj
NWCS7eVksWhc2mp47EgXMtqnsLJNMsitkcdgdUuUbfPoEc8HaAnWs2uG2gaxYAjv
51ktBTmGqlJ/kFCwlYvouDw48UABRIe1FpCkz2TM1GA8LSTtQobuWqVI4AUnnQ/H
5FpPaxvBZ2nqxAL/aJUaVztPCFFDmFtPZbway7sfFjFPDgi5y90XCIRXfJ0cWrHQ
WOz4AvpkUZZpqapxjd5CPD7CsfBvJwUuwZ251jZhjcwawPbBTMmdYtDTZwlaLnwf
zBvQRj39scGCMF4PyK6SWfzjbjRjt+drvLfxPF1DN1BtkChc0oa4BDCErk4eHqCi
McrTusDDHDZtSC49cMZZneCLvxVKIMUrodYP0PX5H85oUSaVvjhobcvrCc5BU+pD
whLskM4FKt19qmcT3vJQkX2Fc0RbowAzhOFxdTOh8ZlERQKkUucyKB0FP7IuQv7D
a2avx+xeG45YAyAYpaBshRY06rW8253iFnhxd41nyT1LRrbrHI3thPCOkAuEHmfF
zsti4IIEZxPb/ZyqXdY6RUtzex6oLXDtTHxN5xVNde99CKHE5FHQNTAP3OXUV6LE
IwuGdMSk8Uuj6K+TYwU8tmkc8NTS9jvQ02raFCyVY8K/jlH/KI7P1+FCo4LOn9eG
byqDhVf+KwdQbU9603flAyK59II+1OVJAsZeFPNDZHcMl1xyglQQjfmigjlMm5UV
FyWn7bja0glopY3GmwY27Ag7Q54oPcAmwFGctVnwtJfe/dVXJyq8NB2nw0BLkJ6v
hdCxZKwMl1U4BQLYgq/TnMGNKRdWwStYh/p1jnaUwlN/ucZJG4YhweVUpV/vb83O
3LPtvgnrGfSwf+7Q4Rqf61aDO0GKd8H1bRDyLLiZNUPvOmJgyOyjS8nDqRfeusOQ
YLH4ii6XZn9NJGbN74eVAon72N+y5wYCL6xngoZDWGEpZa+OQqVMNpEhujpCsyGs
ac3Y/prgnEF7TzAT57KZBIdpvI1jRul5JkEy4ATD5EozK2OLzSgorx3SuUnKC3Si
RCQi8QEFN9rlR/rU7nCrPQw5wI+ah6MZatyvYBYvD1pMrvGRH3WUcsUUqHgtPi3k
qcapqFJ9U5mQ7BcozRD6PvAO0p3DOzB3SKA7e2bQLoye65w2mskSByxU492URt2H
XRP0y+/j//v6gKhxEetI7pfuG84DeyJK0t2PnucExSdwQ5KE7JR9P1oLYCrdtIRl
QVEErhFriXAbO+TfvmRjH95ybIkvLFT532eehuOPEoilw0pM+KXqY6y29zRSDVC2
cSanb+y1eM4Am1Wvti9ltBfDrcfiXcTaiv+GbAg3+xD6vUGH+4fP7uMZzV2MlHXn
6xgDgIL8t9PJiQet+iqm86JhY83mM8pU5V8dyxVyIyGDnZ7IthrU6uy3egxeybEF
XnkRTiGlKDTYj1nsfZl0oxESBPh1cZFoDBNmPfMz5xauWtlgqsr8ORyVifdIGhi0
scqvxVdMxzSEee3s9ggmixABVTJjCNAMoFkNzsJ3Z8vN1Cu6uH/98AWeEpPRsWiU
3k0Pow9gJ/x8+Qy/mhUa4ae3DNONP+mn+JPuveDnGQ0VftELDxaUjSpHtnEvnVkP
wVgGTdT126kXUZjOGwxrCF9k96r/Y7Jn5lz347OJmbBvBT4MnW+dDheoO+vrc7tt
2mFG9mxyExkfVaBZf7TyINeFcu7vvdDY3PNcYoEZgrcsJEoF0hCYEbUES3zYmZ5G
rB1w4OA/HOlZVMGUhNC4AQAnryq6uZGK4OnPOkmSvHoDYnhNtEYMGKjGEkZD2J6Y
gSVGrEBLvVkQ9qvCMWMzlmjvCeE/neFAijU7NWMm8akTQXzHs/xQytW/GXzKsTfS
HtzDYR23gzcPSescyHhpYlFuAvGy4H4RZlVzQDAWYryNbwLE96GBYCpi6RMpaq3L
21lR7WPdEo6XByiB8YcCiRmsStoRlDHBfwm2L0jQKch0zfsTQpHBb04iQIUFZzSs
0XH7C9FEGHomCEHWM8NvZd9B6m8IjC3QKqFfcLkCDkWSkRJcX4YgBRkXk8sPDy+C
/dvouzXJsYoRFRGg7nS6hE2/q1cMpWfNG8Tzs5ts18Ghv7oAQ62qlN3P+X7zcJap
TaCDxOxhtvHlXcz3K8NWEmBzNNkErFSF9JRIaje/hpoSx5VAzrr4ZV3IW40x+hsd
IN8F9j/UdOMb1aKiq+MldX6DtacoEZBxQH294BA/mBaYiNqg7szvUdWG0+yvKOYs
YRyi76O0pzF1a1K7aLxi4l35yxFmg/Uw95LwwpiPt8I3V0lerqrihkcFEIBS4cbi
OhqAwCj5rxz94ReoQIy6S14HpRXx3HdzoxfTQerB65aH7sunyl92ehK5zQPXeoz+
lUZWgn+V2idS4yz9PJSAKbAbPpSOohI8SRMXHlTaIrtNXv2BayioCkmqV2CmF04Y
gjHcN2T992s5wutrRyJg+zSWGsTpkcHBnITrLbhlibr2Fmsejzg3H+CY3AmbFydn
cl6nse3StwN/65gyGTqFg3lzQr8RcxSN6/l99471THNIATlfQ8WhPZDf6JQdinAI
dAutzmzCcOihSllfQLICD5q7dZLA25TjMO1QTTO22eHnXlIkNw5hZcCQqixyeUod
HEPkMIAEMkvL5ArwVuyx4msZr2N4/ncpuRKGKLFJN2T4wE+Y3wB0KCwt99THu3bA
5H8lCOUePhhtFlB3p5XxYagEY5vJbSBYBxfo8Dbi2kBQ+/pT6QhaLRPMr/wfq663
y1uwC1QwGb1PC7mXXQLKTUpsqngyfhlah21aAuUboIP9aqR6DpC10Qmlh2rmU+cf
FxZoJZPN0r6QKLVliVxT1he/WGrtJ4guvOF4PS1UkWY5ddqxCDVXCd/dOamqq/Sp
UKEJol2luXYHS1zfttpqgYYPfd4UWf2aPgD6RR2lsl3zlbMSifxLMqu2appxgvA9
e/i1XkUobu9dAO3HxPzxsq6YF9SpbYIRYQSe1nS8r+m3SyIpSa4lxStmJSeL2Wht
zaOuUCm27XwLG3zYl4YZVgwkAUHxE7Cfo+BE2uE5RcpBoIXfW1fE9tWNKFqmJGlD
+S8nhUlhhGPDLjFK5Nxvhh4A3K9YXRIanSziKPrx8rwig7DSMpBOqDlSgbXncLip
JbCj5xK1mUA6tazFmiM2hzjxwaXT9qsd4xYdRNPKK0wbdSqhha2AFdoJydvpduo8
GoyRsRTLsCLpCb2RnM6r8RjxbOoyd5hNaCzfzpyCCaGSliKTGGV4SjA7fRgVtu3d
DJgU0pQ3RuCEw1sWvN5gJKq1yJpbVm12UA/Yl/W5YaIeNknweAZSHY1dSwJXgUGk
MTCtAD/WckRDXGf6J8QeIqaq+MCgSEatxN0gem8z2nJfM0Dtr9ChYHNRMzEH1cnm
dWmAooT7OnKp37AZ5H1MHz4YK2Ha9gLmRJW+9L3BE9sNFTYTR/ZbVOiTTznqW2VW
bZXsW1NnyXs/ago3jPKBAPCpnYAgyKtBpxXNei+dz8fzldlv0VDKf9yAdpKfLIJJ
4wmC+FaxhNzk2wHN0PLjxYivtBmuj+/d2uUZS4BiMGnZsEJ5jr8NCpArT//LRaR+
m2YnjN6Uhps3kwbeLJOrAKCwRZIw3K4kf4ZexGsb67GmZ39zvO8PxN2PGJP9OcJO
tFgUFJc9XxbvUTT0yMbcJSkAqaIV1XNRwGyS4P5OhLWPXSe2prbs/4E3pv1SBibi
4gDpxLXIEzU8ZLyikPPVD5adbWrYMWJQD+kBNrLNfxPgzC5sQZ62CQ69JRs+T29J
4sdF70APltLc0TnLWUze7Xc8TSv1zNgzMYthUMWsHdhqCtVr1tagItV23d044Ip0
44oB9fnTjlldgPCO1iCKbWJ7rEgGoo++50qMRwa/W2Q59wphslIxItm8+nLGg5ic
AiDn64T6KP48TFzt9qJuXWky/CbXeitQ3G5TKNUi4QOgJqooU8tGRXX7x5UZx/Ys
EOdQQe1soXWvq8nlJ0WACvLWNKY5BCV40lWK9EDXuipf0ZRs+q/N6qXHdm0ktl1F
NowxC9fzEfuIQ3WTInqtkqMBzu4M8hxWHo/TPWYhZ/+bi7NE4KMD4SYjxCWWIzWP
uW74h4Dw6wtrlYlQwi/hYx08eL5f/dPLfWnBWCl8XrBxRX3KWhjzGYrAZ7aOJbiX
0/HKmP0YLbdOHevQCdQfSjKsmi2ADBH4UO3YZqavczOa1+0HFVU7LEPKKBpPyOi2
1URlBn/3tH4xdw3kb0HATzYxNvYM1d4Ckv+T9ReuY62u79SI3nLt2x63G/ZjnoNl
QsgvYIwDI7Tc7ZLIMAUsrs0Mpi84FtvyjcdkzqC8aKA5O1ogGWEPdYBjYVhlzDI3
jFadnDKiSUGLDPgrFhWK17JTUnzXFvNYaAONY3X/zkbbL8t3GdcuDHIjwUyD95yN
orBqrET+qYHqhgAwpivzPgViLR9S4EIr+xcpuG/sYkipYXMDE/wfO/grL9HPHMHp
WVJ6NkApj2ttnhzzNnwM0FMC69HC08Wzw+oXxYmzJMkxaenfu9v4Cv1Xs0nJBcAl
Dvv8z5c8OvVMTL4ZxIa10MGk2+0Czo1nWC8Vr6uZzD+xk2lCvwabOBmEw21zqKD9
+tGL3EYcOy6E5TKaZlQyJAQZSKk55FOxabmIkrC5lxWrGqGl6w/5rbxilCgxIXKc
KNGWwWo/Xx9xaWWfBu+7QFDGvpTgXQzcMEPvDQVa2LBfSGDGjtygLojZAH6wPsr/
PzsUdq50b4CUNactDGCpJc0WaaylOu7X4oZGNFMJnnTABqMQObycK0BrEdWJNgiB
S2MZfBIDLTJ+hNVTvibudeaXtuoX7ORK7/QAaWFrc9biB0QIGIXDZU3rJdaYT0R+
C2N6NEn1reFKJFDL9p4WHvSoE9oOuITgDfcAlNkxjX+M0e1k+GTAcZ/L4h4W5Qo9
Q0qBP4buFLOC1UxS8L2fUlNHhgRHZRkNO91qSC/SENhmYjn1DiYKLbyzu2CxiOsi
AlSEvoYXA5B9mhBejDOGfReL574LwTWKmY/6HeC/A++3uy4tBX446tSHm4sHeH5a
lKVtAHDFzkRPybZX6mrbZqDLXnYntx8z/zJHp9R0C3CmpKtknoyZwBUyiqWXFa9j
nHXaGz2vWaS+fglXDBS3ehwIEK/S+lxZshdQDYmHWYDMSZCLtgiFQ+T+UEIQTnwU
+uDrQZQ3RKgFftsJbJKT/VGy4zTW+El5oC1b7z6ZXj7kk4XYO/2xMzSGWpkOddVL
oqJYB3n9UFof/AtJ7XK3k21SrGWm4+SgRD3Frg+GIoTTlH5WOAaL7i7grX5c4w7Y
k64dvxYM6/bEH/oX9eW5M6uYx4KVn3gWb7fgiPsAUazsFCbvHTSWKL6bh02mF41v
7i9I2+TigiVdWQ5XKOg8T/5yd6Hj6SI9UAQ7UR70gqI1O3vjeju+BzTpPa97sQmw
hl6Tt7aq4Myz5P5sq0LlzAMLlEWSW1bSygpP8NNnVxd1eZ7bBDd2zY+ypGmk+Nb2
TV6F448ZRycpiRl9SeAi/pCszG1RmORUp1+lJWbmQnQlVuR3Z+1R7XFRrjoU/iQ8
HkVhCV5wCnwz2JMzu69oOnpSs66oL4PuL/4sdpKUo9Lo8NPjNVOkfq011nDg1Gyt
2sYHREjT5JRnYgcUp/UxbN6/5Ms9PtPxrx2BSu6xL11Uca8tZmEFBf/8aLddiRtI
i7dtf2A10Z6rzwMEshiJIvzMEU4XeCz5Fuq9mg6nKDHENsb4fdF5o+wBcBOGsO2H
e/ylXeq8M/DnDnBrJpj7GvV4WIvEOcHmK9pF6wvtaw5lIPj6RXFxCWdVanLAR09H
tYPSqHguYtZq6OAMiwINm+1taTI3GnowqutsVmi7RO0KhaNK1oRRMCp0zViix6gw
0zZ2nTO+Nii25bIJ6cKOS+3kN8k9646QHcoQy9NSO3dA6i8qywxB236e5/7BjOHu
iAs219JB5cscs61I1FWeROqurpwdIvVGelnhqxgQs4nh9I3zkf2opJ0XBMMdeYwL
5hNfkspMsDphC8Yfc/lOpxqr0ahvrlu9x6Rc5Qx0dHCa5UfdoQ9/EyUc8kFTqbyQ
p8QNU3+VHL78x4W6NBKBZ6AZZLq2J8P+R+A9PlJujSyQHRyP9L0ZutAtlFmUcpvt
4vPCJpGR+/SzYjdNvi41b1yNgYd91zxdDOQF+XBBc/VjFZ7OTBQKtocA7zik7CLZ
YK3C8HGsX6/i9Y/ixsHU87AVwCtiS3F8wWsPDCkGBDB/FGfMxE+vAjocwf7oSaC/
XBJTmRaBubIoUFhRau6dsy0xLCL7PmI7dyhvpvXeH/NzOS+liIZE/qx/ISTazDFO
xYC4THq2SGgYwSVcknWLTBd0yUkzYnkiGJVxVyo+H4rBrnZLoiSmnyJBpuKbQuq5
HWgtBx/gmZXTLtKfUXCTMmPVU+B62/9yPQpzgJGF9kOd5tZU82L2Y3jKtVKr3vuc
8B4gEL0wRj20zvFjQUH148PqmdplLL+3U1QjHBt5pGyBHwYxIWmRmso5AquiDRj4
4O70wQJW40LxKmy3wcR+Q7RLUK/EBFmy1OhH/byAolfIgeBXpLorJj1jYGqPZ/4J
TRIYraedaa82oNtSPta5Gkt/ViP4E5do0lQ37udSAM5Np89UzXSLea7U/WA5pgzK
TQ+xLkRSXxhFhmWdWbZscKgFfXj/SMjHK2V70Ln5BONlXLsouAGXPMV/Mwk6M8W9
eHKVorxjchEwGUkLPot4dzl+waI/P3xH9mTlPnYwYoQVlTRiVzXvFnv31CeBOFRt
CunlawAmsA/UmO9uVXA7kAdG3JB4yC50WxN+ovvgfPLdk4+3RRMBtuzzn2ER5Eo4
e2E38/xu/1mhgytSjSPgWxHPvIUV3rSK4bjqr+/ZEwI+sK+NrZ1738KzwJdDNgCM
ZKQOJ0WDVGT9BnDoK0aClcwZgnxoJgrJ75QRhNZ5UWzec7TsL9Y1Xn0u5xmjtmTc
WpSQbLE0NsEpm/VblK9mmQ==
`protect END_PROTECTED
