`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
68p5kLvaqOXPqxqEtlXwZrFgD1sR1z3fNVTARZXRHqL5ueQhb8pZNA1DTkHqbiV7
a6TsW8P4WUv/cB5iOaF593qVEFfkz9OL5WG1IrwRCCwEAgkEwyEd9gyMashr4kXg
GrUHfn+SxcK2kvyQpFUvCkZk+4zYMF9zBBUFHNjPDTQ4xGmjvscnTAUWBaulFVX0
t8Z2PkvxjCOX2q5cg3nXojbEC//LQ6cTzD12Lqmhl/DxYAaxwXQgRN1T3OTogAF3
5ws4bqW7bt1LMIHqg9Q5XFavp00AvMHYMP3DNGDaZhNl/HZhPEg4IE15NMshdIBw
BProTVrCXHvPuxCKG+wM+T/Qt+huw7I3TNCHX2JEPw6zM3w5/BliGz+ULrKq7eKo
oUx9N4twSs2M0zIYIsBYl0dHJehS496ahQ8z+LRPoGcjGjrWurILnvnvX1t3dftE
EHek5yLvnawTGbDVgsuytMxL5b/PvvtGCMawwlsxxk6gW+Rts3h0ew8Ce6z1ARhY
joyCgK1PB4f63YDXbd8HhqVKYv+/tKzNegLAelpDzqytsW41/Ywez2YoQt+Z1NQQ
s+WIqyDRo2k8GKE8EutbVI3ggQp9Ju+8/uMCxarQ51SxmnRe0gMo/rbGa5+9J/44
aSHzuWyhyAwipDzlskFsF8dIht9GrpisU9br2PM1JX5eKaS0dhRi8AlZh+lkiqE2
HkYbZZmbs/vCBXslIc5DaW1tLEQQ8RfE8rYGdSUup7X6AFLmew02Op0GyAQg7YYn
6BTyCjApXtgesdoP4VQgRq08OHzz4rDmHcQBS7d30Ug=
`protect END_PROTECTED
