`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XiAYMvCdyZf7DbzDjIcmlv+TLS9TPO1GzV1Q3IESzEsZs5rGvdTjYh8kWHRLPHNL
pLF2Q7IYNo3no7Kyt3MsJfB0uIqLglLln5F6198t+c1lTV7B0M3Fp5jkX6WesUCa
TpyX0fD8QNoaHyTY+lPW0kGJywLb9rjI9eunD8u9v1W54mMBPBylLGN8DzThYAOZ
wvoCeAUkhXNSvg0ebs6N8GHhrHZKrp0oepOEk0UGFEILNM+4KOMfA0JSghcQhx+K
4AN5JHJZEWLgLmKnWp8SVDlJWYplJH9Kyhmv4yDjmlcSTzDDVh0k3W9rQcbs3UvQ
J4oZr5MnJ63DyjOFDYnAaLRVXz0+eQLfkjyG0UeigcF1jzaWIEOestkKQkSJWaX9
N/161mBaX+AOPKp0ZMKxQ5nGxMxKrMNo0jJC4DHTkrs8GkWtfH1xU9hPgqmYe/5t
1ElfwSIVyRbPTGcHdq+7YdLub7ySxcCnYe6Lf+0l0cbRm8bdac1weOD+LZ2TSPZ9
A5Umq42Vgk7kk6xmJNmSW/XHCiNcP2vU9BOHzHvDKy4YV5EdcTH4mLeRk+f7PU/n
ufXAmMo7Km5U8l1y6BJgkWGeKjfRbxyTSElXLOgLGNuZC1mBGUIlsvmS7t0CeMhE
CC0+TWf//RBs+Yk6I68vphN+LyglIt836pa0qwyAqNRxJAOY/zqbmaqL3YDA75yk
1D6urnW0AToVVx39FNRUwLLxX1FxjOoYcfkCXuEXSMMcuZlK2U3937MvqydNxkIV
V8vIt8cXma8NEllU7SJ0NRV2oe4bfNaca5UpEr+3oXHMoYHTmHGz3rec/b/noQsp
vMcgC8Sww6asZtgwxYg5eY40Z6oQrPS52UMvTKbiWoWsvkNicHLyNIdexqn7CDxF
6bntwHN5Vca02uD+PQUUF3c2XZncgGjQvgEBrHtJO7vTbMlw7dp5b8hztmbuDHvm
DeUkp6lRw0/wB02gPQPaX0JjooBOTO0SPnQ0XNaW0xe2i81CY0Y1MxiS5buu4LV4
n2NmU21gkDaACpQ81Ja+7ygAT7prdPkzBSzdaxfXWSa0cVhy2jRrr3kJNdVtJ4pO
5M/WWrdfrXpbq0b6M82KQqThunOpE7HA82JW6gD5xsOXbgWZyYsznTj//9ZGCDfB
r2YlitOcmjTjHo7E71f+M+T0eMwympz1auS547OEyOfISmIWAGmr3f4iyfSaqiaO
BYJuz2uCUNyxMwWICOvCs9BWTLWObQhpxzWNJd9z3XlonxM7Mm7FrCxvwgOJMFSu
YD5mdaSJaP7vFv+2H72IQ7kLqeZZKUVK50XBliIcMOTWieXOE9+jACCeOqIzKnAQ
QWGidRCI1muvP8EhNeO2kwdyq2gWL910DDcYLOFkUkF8mmrn3RVlhHRHviKoBPdW
ZJVBFf9krlOtdo8S7lBkvlNpkrrNAybGKCHzvv/zxKgNDmkz7HMCmffZh6jiT8Nn
hgqw/qx741y0NSfyBvGjzy+DwwsFS0ucZhqrGzIZkZqJ65eaS4Hm8AF5RNuINDLs
klqpV/FuXCieMJnLGKoAX2r6NQbeKGI8e7G6Suph2pWDH2l7I7pwHB1a4cfoQWlG
gEhK3FJu8ruY+ia+qmL5ovbO9p5HmKyMsXBquQsKBwUXGGiyIyzy2bRG75qWPr6m
5ZR+Yt8HQJU8sBU6YGW/vlAtihuSPC5kj0ElzVFhXiSDzYyh087r3zPqbACy0J69
WhJMIRyXijn09CANeLELusBeRbIBk0knozVW53M4FNNpqvOrTIJK4QosMAN6xIO2
JjLW0z4Z7YZam3PQLZ1T8jabHomBXUjqmOecLw1a6y0AcTKdLOUs68ety2kZ0h2Y
oS4DgB/VZbqrEEJF06o6/zgIL0jAfqthEJUgWeQommBOLJKliEzTMWIT/3FLmmYm
H7CA9Y8iBk5dutdv5KENt6/jh2wHdW5xVhfNmeCMsM0ll82P0W5x/XaFtq4viBKA
e7JlIHKEMBqz/R5KZcDk3PFyh8GGpPaSAq9SRjNXYjk36r7KqKD9z2QxEt4OdMYs
fkxtMlXFnhL85GC2rebMlieKGZfq3gZMCfdeBcydYJ5RqhhjuMQWkqlFeDeeyhK9
FTpfrhfSaw1i0ydM6Ezd31vX3l/pchx/9O3EqFcfMpG2r1cSexWhpeNxmq204jTU
pp4mxXJT2Pcdk35CtGR8LMpGR56VHn223a+cfaH4EzPt5HwQhuItGqKK53bshqTe
qSfDUTLYldPfD8yFVBJEBjtWNiOCNo+rm2jpdWnG50B8a947cNDJQ+Pz0dekz5Af
zG2JmYXXSFn2D8o3zOoV4CsO8G+/uRzVD9ptBbGscBqim8EnvIqWNHN41TrALi8v
j5PnZNqM+hC8lMDMXFvI1ho4hUIupwbzJJrlQ9FmvN+h51PGOqv8PDi0F5M+Gwlj
TrXaokWPdTTMy9UvbNvYYKnE3IOd4lPHUoFtBLC0EdwjHKEMHZuhp1E5Sg+eELRk
eJhAjqwLFtJkrtXZ1RGSDjQT6Lt0599WhQ75vqHnOttSTLvOW7j6cUU2DMI8Xas4
i20DfN7amSlL8sW77auCkTcuB9b1yN/n7wzPtifFD7LVHbGRxGa2B+hz7uyamzOm
vFcP6LvY84UGEShHH1xsihkvGtirVu26zGhP8Z3R+6vkRfwo3NqDK8D1+l9wBsmG
qCDmK2nFlW6MT8nvgVndTDXrZGHalh9hBwSyzNr53iD6Vo4meNGXAwddF4E+BJqk
jfR5wyMRQorIppGcgxd6ztCdgET3vwobYIu5XMsuF+Nh4x5bAsp6OLp9OWVxT5yi
kbTpm0zjv5F7vkpqSYl9m/L0wBDTn7eCpE3suFCGrE9rmlYaY5Crq4fvZgOu5jtB
x9r72o9rqhN9ul/+t5gYuAMRZ0j/P+YvOCzxwFhuorfoYEoM2afYwJIKYX8ssVjF
1Iu/a0+6huqK9Rtln1HCzL01VImB+UXhYKWKbcCX5aVVB7RSiTJralKMR6kXInyL
YvHvPs33iUPVFhdyd3oYyFXHw4hB+fdiMUCenS3y1K5fiOadxbL40oA/1qfTpXqF
PQLpijDYNwXVrnnK/5FSvRN/lNJ0HvEJvFznFMaMvLB64u1JjUldV9gQCufkFS3U
NNApWFjcCrN1dvspsKYGbXRkmFOIAC1SOTDMJP7llH7DhReIS89DP4X4GWBJqZTo
oWbBMDr6XlMoHZL6s9F6mqmntI93GjChBuLXP9lFULB+5EkN1OmLrb/d+WXA+INU
IV00d/iDd8eh9zahFU/ZkdUM+pzIg4EavsRT2Gzqbl7vylX5JmjooHoe41rvcHzv
LV4uC7+epVbbOVQ8Pi/aD8xzfoS10gS8Dk6Jk9NpK7trmT8U79JG4iOdjlGipROi
hqh4aPXrEIrMrAOBSEY/xvhUDdQs4+5Qqy8jptCL1lN4ij5mgWfKU1z2zVufIHLS
mKlqE77kbOldTa4kmcG7kqT06AR1I3D7L46Mrm7rAWhDE5PiiMD90IhjmfttAXzL
feVCc1sStzi2AGxCi09swCNjlXKpjvy/1s7WU5bl1OkeEUoV+f07fStAi3DfGpJC
o4tKmfK1REGvVdfBBIRYH02IT5H+kYqxKnXsreU1+JiQrix0DgUO7qfk8DQlXIo7
8r5tQfgTiK+apLOJ/zwocZfzm5+I2MAXeuBjTYC7bnovvJCzu89XjHE3m/8zGNX3
1244jvz5DE6b5Z6cyRBsMnx95zTBZ2O8oUSo1kmpMQcaBIpENyKj19ujV2CDmb1u
ccFpzgutQjYsR0oE/nonJZYENAasrF2Eh/AgXPG7b6fZUOLi11TOJA0c/OPr8UcZ
7Xhg+HRnoNMfcfsXVXKRvMpBrPv20sbBYI2FM0LBdZp5nm2y8i53VuiqN3C4lY76
z2cH/Z3qQ3fepjHSYMHwhWa6eZydh98NlMUcd3f44LEELN4cbuyy9mbllirQRp0Y
oo/KPCQ5ElshRb7NkLFRpxgsn0+W5wqnTwj7DU9Bc7WUsn7M/9FpIHpO2QrJ3W4U
2rtfjoB2iafVvnvtdOpI2UIObDzA3eGuNI18dv4iNz2HJiZGejU/RDIJpRHDt4MC
A1WJ7urfOU8Omwl5JN0qBcWVG6Ycpsm4+ZyH7E08S7kM4UkkZnPls6hhtzZKUXye
dAvnIBamY2PX6vJSGFZb3B6miTUsx4aoNq/qMfWcZV8k0khxo62ePcEb46qMb+3b
IRFZXeleWEk5GdvI+vJeQtvBrk3veKcri4zM9AcuTgvOBN03dztjhV4TvOte7Otu
cjwwSCP4aice04XX2G1MS2uJobeUKkajuTDGolKyC3pIa3nPXhiVazRXkDVL/Yv3
jADSXQ4omp6g3BFUQxetigUz+JfngH4cS93XXEV2w6f16nnySNll5FzdhSJ13lYr
bqBQjRmrpchVg5zHrECsjpw5b6cWVPFQ/Wec78wiFk7ErbfD/Eg4p5IOy8XXMtv2
5bngzCdYt27CGCR5nulzrAai9lJD3veJLBLLi+mHjy5RmpTR6ZAcTiaNu+aNIUce
1GTZLbhCEUwjFBdBffMK1QNIqJljkG/21bkbvavxywfAuK6GKh2+uW6NFeTP6mN7
GoQLi7nWtXqZMgpIxuFrveXLxPr6CVE0mautA6D4X0m2es/yKN1E6+AGuVgDWFBV
Ko11TiDDtCJCM1qhYpekL6pEM6/ARsQ4Yjq7VNl2etk+DsSeU8zP6FeO0DifqkAl
T2vVrQOllt3A2v/dUQLtHDD6kgK2dVJbu+uif/M/jolp5UkgsVwgIYW0wocgy9Y6
fzV6U2+0K4od/LOLDGhtsdqi35daTwCVg7As2edXgC/XZv4d26LKNS/z7eOHht0l
ogwmU+EBLiDA02Q1JHO2L7c+Y60jTtAx7TEcGe/Cgz1p4zVPTuwFrnVtelBaPD2X
SurO5vQ4jOTkyeKbkAKz8/Z7DhxHV13aJXHisePPyQmnZtz21vwIj9Eo+Pm3kpn8
KzwaG8O7SaLcj1MMPdsj8vlB8jNDb+B1jqkIgXV4w3z8VZWD0mNV88dXm4PsXGaw
OQnKfSZa22EDzb3GTfw63RqrfgxLTZ5i9HNSVHpO44mFaG+uMJicpp3JH++NfDMv
qpv/11xEZzTJp0/yTrDg9Dg+73rtSUzQT4mfII07gI/+DpgmfCbrEckXBwcbGMRN
5J8hZdUuAfOzel+/ytO4zOCg56Z2L0VJhc774ZIBvUWaNLmffN9OinMv4cUoO/dr
cucnsDOpYieuqfvbfiCf3EoTw6TzO6yVUYAq3EGdFcVy6qQ1mL6jUWI/fhiJh1ZY
TdhZJP8b2WfJ1Bwu/IrU5AHX5p/BbWECApyAlM090VICm4zPPHCzuH+qHCtgtjVP
OdxM70XlFSgq6/ZfjTUfVYT3+E7uauZvOxWBbbNgn1rf/dfVQqkPazdzR14dAgC0
w9GgDogAvtMIu6w6sM85vqaf4wHinafzFM3Lcl+wVSdzfzeIMoZ2cywyok6AKkWI
jetHtzziHbkEkLmR2sM06Loqy5o0YrtCghPbOphjXcx9XRNnnDiKteOEZhDvsuzE
gzA4hlaOMd8c69+5tmJ2ZjrH89elBmrCakeyzA0CgozkwAh6iyIqpxVzsEULOPqN
EskeTmy+qFt4PUUQhaOtPi/h8Cd/F/vtmLuKQL5RSYVnVRmxSLkBiappFvMd67wf
1TgozC99ooOrwZ8nv7LWJ+3NUrxcKhUo+Wwbiy71p627+F3pLljDCkLTm1rk2WwB
ynXDn4D/6TsOYYomxt5EGqfs4sqqug/Y/Bsf7Zj3LWx72/qPH7j9dYz1ls3gC+T1
lZ5pKO2fFTP8ixLLsKyeWPtjjOyIraABPaDW5RsKROuNeWXh9vTmi+DFQQ5hHk7y
TnVeW0rXrAHMhH+dN7YCPCH0/bsm1MXr46MqtWtmif4RRa3eFxVRcATTy/WFQW9e
EUS2RyKDLzzuIKSFL0Exa3xtIRjM5ftRYxHYsd4lDF64Glb4SReflUj+pgk0JfFR
ey1hiw8c5/EO1oBWJav1xTNSywSgQ93edgt9+6Hp6CnhW2cmSCfvabcR/cELWiaM
Z+clINRge2wDv+b6IG7ZRs1pEMsJmqhKwu+wOoJZ4SnU0JR5osC0+kP+6puPHLgf
JbSawJiBc13zZhm8ydgJOqz8aohMYvo6/MVOr3zw/6g4SADF/fU5ogdueMvDlxqC
RoK9dELxECUHPx9depkYAYGbVQhnM4oCUheuwWfXYgDkQY/ItmElpC/M0QPqVWPq
Y0khgvlFscKTEiwz667nQF7pZpKCvkLU0Jtt1cteSZ2bjnFevWX9PBP5OeOxTxMk
7SPdQty4+ch509072ztcYns1Gw14TP6Zaq3i3PFd/eMiKudlz+H0YeODic1JRCqT
2aEklb++sbtMrGyKUMq58P6TKXYvUtMFPlm76FMVCBIbWbXeNqQ29ZlNNHOhkXI2
mVJ9ritras9Kc9GQ3P5n9rA19bLRnvRo8WBxt0j1Co6QaxWoiTcbdvQ+JFclO1mc
n8138LwOH75BxD+Tb3WfhNwvjZZ/zfdCP04CkSAbwye3vmy0UVKxKgC92OPA0oC4
e0rHJRHFfmzocWAR1Mmj+6Zstmx+t/NU/UXLzD1qZuF7aEGn4No8ZXFwWRKDGr3T
I8ecNgPCc47DIlgnNr/uCoyq3HshSSKeq/uD4tHo0WD6ZgwZasWe4XxNAMCZOUe3
7buhqbbWR1DdzQHGi6Rqvrj98T3gbrjhiFLwHR6BaAMhEB1Y7yKV4Rdp/7a9bVLd
5KZqzhFxVaCfOMrjfQYsQFQC9KcAX+WlXq8+4WONZpmt2BJMytrg4uIAy87nheQn
a7YAJ95OkaxhDNRgqOp+1fzOI2qQxE55iePRqZ79+sedcwmOHk3Ab+oG3wdKLmpO
+DPrsmLHiPVlkX3ztvnPoQlxVylLvz4TxFFnN6CEM2RY/SBkJJQrlLvNOu18tCYh
F71e21/Ka3qzL03rm2PUkaXm8sFkkFATlIsIonzvH9lygq/3aNt6c0IBYTKC3Nwq
pmoAmAouSLDrVbxvXAOwpimpdicHkIZTt+xwAyrYQAE2nMtWg4E/nJa8MZlpv3up
IyQCbrCNFTS6cF1aA5OpMVpMTxPG221LfTvEWKiALfpbse2RSDMvvODbDcEhS24f
WHCyxwwmPY4KA0EY4svyVjyF9xZtd84nwhQo1L5T90VTk0V9Rs/jvqEdQr+X1lwb
wk+YtbKM6JgRULzxnSAibu9HfYVU1mL4OkCUAlS6+sIt3QCweCZQqI8vPCtqzc43
7w536lhFqtt+RnHKfKO1k7gUH2yAUQ11lyMr+Y1r+X5nVDwUYDewQCfj7LWP2SzD
TvfqoiTtBFDB39MaBhLN5XGf0A5nqhBVux/EYphY28CZjEOyq+LJVxtutURx5IWd
inNk7cGUK7m6SJtk7AWa/8FdRmZdE8DhpCwc6RWlVoyLDhSuFFlW550F9P084q7G
8fe8voraqM6aAKzFVMt4OS40x4sFbyIZSR3omQ62fRim3S4/TQgJk/Ns7bP8uqC2
WM+77HYUECcMTPY2kHNRyt839F5KOuiWLm+KtKyR0uTvkOtsgzlrw5v+J9TsPlte
ROhmGzDjnC18LUrL9GWMI8GRePR7gjtUKUKAnF9TJKDbcJqtC3U19ZsHvka2jKcr
oBaHlDKKeFNt870nebFHBxd4vY5ld1wGRn0pBSB48ruhNIbVccrOcMRwrkDCtp5n
En5pGd+pzpxNRf0JCUoG6a83CHDndau8HWUW++sPh63d+nXVxe0ZGKzM3nNP1ndR
pwTkcAyTUgLB6hyIQHgSuBLZh+Meu8HoqtxxXLndcvkP+ZaKogQsDYY7CaSkDEJh
avR9wjKJZp8MhMvJV1EUw6+TYcYzYi9KC2V7dUmp5dq7khHZG9DJ1GsgaSWibHv2
00842dUDA5oZywJntdpfga/uiwDZCCyvGCaqjJHrPI+Rie7C+M5p70ZVab0jCjmj
0lf4TV9WX/e0e4viXrH4At6eM8y7uoMtx3J2tYWNzDvuFZ2Gty6oMLwxN6NR7JDk
QlbuSyhUOfhOaPqOcAjr6hytTZd1cqE82tBG8fyGDxoRrLBuA+JBhH0ys6ynH0H8
xrKzBRiSXRRzS1KRUWspCo/IXCC0IU+axskpAl92HMQh9za/hvA9qLw/SokpNU+Q
Hjsvz1jIW6TJTlkiGiHgEYFyeMBrN8Amhkf3qkQxI2/mO1ebq7ds54iTdkS6iR23
F2qnmv43FWNtgGzOm35oebSfE60B354xYT4r340u4tfHHxYLAsGiyj9rDuAB57NT
kpIiHrtbACPxR6Y8fAls0UxX92L+5wq34/DTAVpxjDsAE0fX8tbAHmY2rNYSHwRU
u6bFilTejvA6W5J+M1nJIfxOkKlupgLhzk0lJAwMNcvfUbr+pAVBS5jaeorawX58
d602y9ngxR9a/wqL+VbDtShNOQ/Q5cbyM72WxJwwAqKtHeU/nKB9sbe852mk4Xn6
5N5P5capJXQdmu3BWDtIeCH+uIzZg10O94QetOpmf8DZNrdZNY5iPXQvMFx+SkUv
66e/lbqPJAA3hxdwv8yP1r5b/ANqqCgh0bTTjnUK09u5kFoDB5AYdw/RwVkmJTsv
qnQDMJd0KDrT/ZZ/kFGZ2OJtSTsCDxMy5WYIG9nxjnETpvq6b0Q42bs7UTMq6ELx
pJ59kDkhl+z/crwdo5NBA/OV2WARqe16cefVK0NuTnFhTdfnpxMOGSkQEqEhDciG
IU/13PCr4IekICxmHNRTie6k2LGRZrQZYyXu5Xxt0DkC0JFIyry+lQdh76NjGZeT
1e/uZSv8ZbTthRJ6v0h1mspy6Rcke3plECMBVwHd8TYamH7uBKd0zIcI3Wkxn2kK
YRRK+K0wDyRgpv4ukaTOSIi6ysZDE6ZE0y/1y458PGKGqqL1Fd43hhguMeqd9BE9
Il7WZdS+yqIUsIFziTtMcjrg6wemLGtuZZHBXhqvW1K5W0uVQj4MQciIVAEpVJiV
Qh3QYzazB5FIKbU52PosaxrxpxL52mcnX3vWz2ddx9oneXZjxGXcbLre5RO37Xtn
rQWe0nv7RWJwvg2Fb8SQCDMgbhBtU9OrR5HX+GWr8TALcUUHDLxiWLFaQoQF182Q
tZSPCL75q/Ljg/16CtoGtNpgghcnp9Ax2rqhQ7USNXMFZwhipWnEygmISkTnzKiq
05L/xHcqnd/oISxojLb1UJ/auaekppo0xITJPzvsMwsLnkBEo68b4rOqcqq64P+j
RSbi6KSOjthhzOcxm0iKsEQCHI4/DGg+BbS48vddH52PwBpQKTP6GR8bbezuFmJ8
elRL3ZD98UeLAQGdvUsv21xTqLJYNoKboyi29+SCgadtSsk4MJFH9dEquwTCuX+1
RyoOVZOra81/w5alFEfUIZIdIYFXhXEU/25RX/VyAJSfHizVkksAxeoPuNo0TjD1
bGkYNmYbWa1+jZTfswOOMU585GvuIIP6LFvS2YmRWkqgCNO4k7an7CiiSrEn/8Im
2uTAeWSRhZiHbQ3PA4PGu/bwFJVI7o8JYAMQ1j66/w0RkY9PzW8vYHPgYLn1rs1X
+wKQW8lwYhtLq89tgNlmw5kYm3ohMgRjwmSL3do4ptzk6mdbyDbY8TUORfJeCHKk
1Cm11oFiykg5m1AXlZxQA3TiQfBGCdZ5j02RcA71BboNIt8arc32ko3OBYsR3/c9
51xgd2x2AFEp6C7cKvDs093KOEG7+YipT/lEI2h4gn8lOZ4dMs5Ls3esl93YieT3
YZbDyyBJaMlpf2KxtjWlZJAC+MUq1SvaXP709upM1qLJA92EPjPt/quqsvTIj1dk
/53PfkuWHXJ4zbAZF8J87s6UuXDZK8XnSEwa11v/MvLqqz9riIWA4nhFfwoLgZIn
KpfBH+Syf9ZrSKjz0xTKhpZPJxaTHD+q6hOQdBAwycHCWh5Z2yW0hl+UOH/EqDzb
PyEIkfVEvIW2gllvtHXARjdLyZVeRFa6Yic4GmkDHB+8tg27DbKFwSmo1lBcRMd8
azXJLpjAYW4UDRIBf6uo9WEWjzWmuAZBCQOrxtdFef7ubfnA5A37EIME0tqnrFqH
veEbaTV5aCGqpgXTZOsvwPdHiNPBmZS2oV5QoeQYH6VWT3dQ+0hWmyQhQVVmWqAz
6hy2qocJG7pSjQkr7ec3qyJ3TnNUrlnnbNUeLEbLjWZ1sIBzS4qLHHshwY4voQtE
xPRdIkvIV4x+Cn//qS5nS2rKLxW+gFJUCZyJh/gNM1nPUhyHz4H8C/AZmsmTH3Sa
tJ85djOYBeYOF8ryQnKsM7ueR8ofbrZIm+f8IWiRo54fkqHWXnmhswoDlU18XdFs
yI5Njh19BxwSOSEAEuCkntXMrxN1Cb0nK/X8tNRShpHe887+Zz/H9CgKpj/LBwT8
PaAgjgQtV5jgkXKGnmraK41qTk3vmWsfiub2O3fJC8pS5DLxuWeOwku+vS+4o6dE
Y8i9btE5gY8Mek6665j/+dKygrPb7oGGmaUYHbOcqkapBpNCh3Td6/J/Xen84SOV
rNOKG5PQaqu2SsiI16dBAV2xZKZSXXVuzfEwSDB9BBWglM9F4CugaeZGTAwfsh4g
ldHQtueu/Q3JFJ3CjObiLszYfP+tbyH1MwCkoKZyGjJJkZv6lK4veQkpjsVPMwE1
fK7VOrvfgzGrJNfiP68OeNxcsCdsXRyUxTr/snfYPL34p6GUpOsr/gYDv60YjZAm
a11Ip0KJNDKEV+flACOLqNTeJrV1UQKdPtryy8T8q8zoyhORju1vy8Ej28ASYb3i
huoabxKG4/tjMwXld5IWdYHwhl5OcySc6de2sQ0MhaDXOTaxpSyJLFSDgNb3ZLkl
8uIKC1aGOboIqeN5wF1X8VPiPJUd/n7XIWnOjjkWIjvvYLo4DP6imqIupbR8NPdD
KlMl+ew/Gt2TKkNcgTPcd/KJiWXMnm86MnVodOAoD2SHNJifchIa2OcM0BHXDN/w
Ey4h5NaX7sUFGqtIcZXpDdh04LRwkDQYxy2mjEZlnZZPvHHdFp3ws8VXh67UCRU/
87D1Ww24GOXotec/FWT7ZoA1Bh0wVe357N5g9lL7GfojvmiG/MW4xKMbs1bxvSGB
fKdN18q+sYgo73zHUDWHQfhB2GbhRQtso+UHqMYQqY9TweXs/1LQdW1QT8Vp1OZv
JJ3r83fZop1LPlJN0wOvdg/hl6ZA7LbjpjtRWpomcMj8gvftlUTSqRprBsw2Amws
H3YoHCnW84TueMjeY6p+G9/BRozAh2zsckl/VGrrweIQ3cSmPQ5Xab94u2NfGVHi
8nrCQb08oMWkSxcrPIEP6USL6uwTnauuO4K+xQeQvoFqPG58+yy6h+gXDrFxVSHc
JZVEMpSmAQRTQtDwhEINOSug0ru4QGE+G2ULK3VJuix7Io9d3yTmxnBRm2/eFHu3
OlPvL00SBvIJeK1ee0rwCyLG/FauN/G1Gi9jzHWvDgNkL1mchaicjuQqL3uh2vEe
dIDwQdPwL/v/nsYVpE5jgUxZD4zpRISZ2gkHNrU91jrZSzsdWDa2D0jv5tt8Txwg
NPg3/7pkZHthmlXLfq/Jr2lPGxJ8xpyhrxRtvA+tEM3KGiHA07bdfyLEOZ9C0dG2
rrCq9iOUZX3uxG96p7upbaMTx69m8aGF4QzY/LuSOiF0AeJAYkq0HIiFRIbmdoBI
iik4G5oltsueaKVUrxwpzmWDnz4eZJ9D1eI4++lVzA0xTaFicCdFLu7OO2OMtlvl
EoW/iH2bHbm4kV/CxZ4vLB4A4n8btDzofW9PcDh4eUd3jUc+Rwsl+ggl4ZipZhsp
kxfUPjRXBqtX2TCbyZChoiuw8L8IrLFnkfrnTK9fqTpsXmmUhGYrC4U6kdAI/jZC
Rx1N6oFQtpGwimyT+uPKcsAiIThLLQcz8+o6yJukeGt6tc0uaMUkdGCxcEIScjQj
zI/uq86hgyFtY8V/P9NZKtElF+K0cT0jcXP5Pr1Pc7mDckbFRmciXIKXIMZiyryX
gtMES+7aW6bBvmSltLzzUfi86qDIgOAWMo8NUX+vqXqYgZzRghXBS7ZWoHa/Xjtr
wojMJAAbSoH0rkMh/4NkCXcXlbrK/J5w5zEGeskUsGdJeZDz6uBvPum63d1x4Ti3
zha9lmVCwzgP1eabYqGby3NPD8lzZpvD7mBuS+vnu3CvgoFBlHaX+fKmkREd0Mhn
xnpVTmUKrhhoPfEjjRVp+kcUeWLOQg2NQh6ShXLqj5x4jcsfnL67FGy+SKU87t5Z
ckuT+DvcJOEWjekEEW0LNJJjl1ErC3hoX3ihkzC6irnJV/J8gC/hNc8eHrtrn6an
JL2lz0RK4fn4wQuSM3O7MtjUsREysWMXnvGGJ1Tuc7Q3fuq07MUrhkSgyUteA7oo
3jK0RCGHZuxLjKe01BiLxxZtKPRIcxQ9ZkDpCiItuXQSmQwjH0Tqdexo1BmUVOze
VXvzdfeHCFE/FQCQJmvi/Qjimfwd6LGD3DoPSZCmseoVqCowQ/LpRhRl38Oz9ARi
yJUGPzUuX8fMjxSwNItH1ZEqCxBZXMHYMILeA+wySQ15VGpUAbLWbfy/shyP11Xi
QzBU9K5Znjg4KjEXc6FebShOnnc1lCaX/jMjOGxs0r/LqQDeLh3TlWKg/9ZFtn0G
ThG0+TPvCeRIBG1/0HGyUoC/drrmEcG/rDkU69/ySNbenwuK+mqCNgeUZIz1ihK2
LvEPNEjhvhwcTTf1EQdYKk9jjGQ5kY6IzMr8GEYLiozQg2ZO/69jfs2Ub0pQeSX7
E12vybrBrq+Md2jXAwzze/h8gTxEdmzGAmtyUKBgfbBSeagsWPZXI7gn1EKkUYxP
d59jKVf/O47KydgV9FYS4Wbn500ViLyH8dezsq8HaqbxuxBcPPMd9v3Kt75XiK4o
r44GjpJcUzz2Os8MCBvol4ZPShJcYY7XmOZE0uq3gOvPbH8vb8DmCE8bxTnT0U0M
AfT/uAZkfMGNnwijmT3C05x3AliCXiT32jK0H2jNLtn4bzC49e2uC5F1x/Ld8M8y
R1z49g3m0RIxWvFCsSRTVFCQ+YDm07vJQ+mY7/Rb9eUXq98f1zTDPAfyBKuo+FQd
Xbt/ICmT0B8TF2du6PsX3nTh0qPv6UX7GqZqr06cfaISknVZMt3oTu/V+2kDr5zm
MkqN7/epkompTmDw3OHFnPIT4gP7UejCGvwAkx2fkVAcaUqaTGFuU+S3JinLuZtJ
0A750xm2DZ+NlIoomczcQZvjji1Q0xXiXd/sJ5bITMF1FefbZnfikhaHqinXH5AL
x4rxrzfnibCFlrSxTgD7CrWGY+gD8ai7LExngFVoMcigkOxNvIaJGI0dI3xh5xi8
zGT3TpiSJzQptjAjuVJLucxMctXigJ3vHy5i0qH6iC4feS8Ojc2BgOsB4PGkeiqZ
nHeETjnnuWEFqmwVY9YB9O8XwrvpvKq3F2tSXfg4L/yiknsMWLg2KUTsHTTT67xt
fWxrP3sAdhPMqp/HwmDQOEAQ8E+moH//7967WI53bJmCJqG7MgPwJrsm7+QKe/XA
k8dCUFLpn7B8UQHz8KzY+xYxHeSvm1kCf7fPdIwX2BogKvsVf0vgs52lQfG9nA6Y
cH0zqWW2u2ufHlPgwOJtuHG1Zh16doCkkDwPKvSCnD50NMgSOr9/vuSmOr9gvZ/5
xIbZ2OZoh7aA6bbU7DCTY0cgeX3okqEqIhoIJhAxblTIWydeXCCVcD09Wb93b1Ul
0e8MaP9UYPlCT0ZjWnVQLy32PtnIwmVq8FsEME0x6fRyT7rOROwoKYI5wZR7Kj22
1YihniGFx6Iok1ZTpX1k3KSFej5ZYskyIoKdKxbMgR9PyRAL8EPbmbaxf6CBX7MD
4SQlQ8W49XEuExuh+tP/DsgXwZhrkmak+1jr3uXmH6nvUsK488RBoEO/3u1TrbA9
TVuaXk/vNu/pURQ7tXmC7hdArQk6dP+34u1jwCNV2pke+SE2OTRrKF9WNZWRsvjp
xSiGHpFQrK6mm85nfhV2My8QRHiZcl7uF8d8G0dFWT5waWGDr8ZLo9ogSVmLOdzn
9JfszguKCWK4PBh2DHYuwFDc4jtp3od+xjZQ9u7vF2A6iE0CA582y8HR62Crjbhh
V42IYxk3WdzXHp30sIgXuphT+y15VbbUjxBdFzXebjKuprQEOodAYo79kX2eAUEW
EQ8o6KgOYX9LVo6EnyyB4JgEVatl3cYQlCyI2WTXlmMBLTa0CcDuiAKxv5N5DkkF
JLpfCar2ywLLT250kKykmrCN240PmlTV0pIWG8Os+YaJmCaDdLMG+1J+RWkDU/lZ
r4G+TDB8y712DI15zrGSqDI6SFHbKRXHRL271AmiFonZtUDE39exJ1N7vffFg+Tn
9nQa0NYikegLh7klKuGfc1hxAkyjQl/mAD+8c0m9I3y3/OVhDeACNiQggevdWWjQ
rEM21+IWPkfRZ3d6G3Or+fnbUWvQuac5QwDsxcN9ow9j+Bm/Vej0cmiT+SW592LK
Pi1prcAVxtFqSSeBhyC2ucPXih/nLU9zrfxwUUCn/mLH4yOZa4sTcFY+F2h1YCoL
JyVh7krI472F+94Oy4buZoquRuo/s6J6olp0OYpJqD6qpq+uzt5MasBaE0zjK6+N
A7gHKktfmcwxFwVz/0b+DoJ2W8+MZsOFQsAUDFKIFER9Vrzms6tkFnnpJQSgDFrZ
oXaWCKqLfZ16+dTUR4y2/auuHtK36x3EHH5V/Q8d2h0D4H789ec3rtkBdZ5PrVsc
rGTvc1JY3m0AYqSabkIaPnTd3Lpz1RzrpSK0JbLGaUpJh6j4+izZMuKQ411PdRpw
bpezygQuESiDtM90d7TvFcNK1nSzapNW0TJDwoEkAG4M0i5+zU4S85s8BD68TRVi
F0x9nGIdDaOp4TTHeD6s8FIUDMqdJ3WEHiPw6Q+tTkg5WdjNNHUOVzUbWWVdacDy
6Mtqy+eyriRQxD38rc9AQB4JC36GOBU6+yXYoQv7o52yHLwSA9ZaLqb9VWcMyuUm
MQFTGHW2WIordmfvwLwpvLbKt8evl9NiLsS6F7jdlV9LPGFHKKocvYUpOnu6mglu
gueFkNpbzKLInX1rWgcu+dGsPDnrG9AnTtFwJx6DZ+cUdc42ISuZL57WpcDG2cpl
6OvxleRR+VrGAsZMd9smPKAY+I57y13+MzPaWcDf33wifyovMZPKGXIrM3kEueO6
7sNchdl4BrUwDYYaqrP9Qi6+PKrnNq9Glr0kZGkf1VhHd05u6Zjk/fGY4ifxaGpa
rgjjD3iyMi5V/WmjvTtQkNwh89fmFwK4Ci/w1SjwHL1RLLRnaRumwjXFbR5Mju23
MNosKkBmNjIt9OJFA/AsleY3fSqshi2o38Z2Yzy856PqxJnBpykIknxSpvGXKO1n
cqtE736Ljgexp/PEEzaF4ZVzy5QzeuupxofqPsvQK8SVeZA981vioSEnRiouQUGf
pr/JNzqP9JzUvNAfsGw3SEHULWN8jlfFGXesN4RQ0o366NitpfT9lv5IPzyvRidA
g4DmlirAJFdWxrm2Cy0mQ/Ym9j/bYztlQShdKkOV8IXDKhzCrDoLxfFN99X7xeuT
9NTroGIAF/WLkhgW1iUqv2KQdD7Ecbvr1NJv63NuwkW3zJ5eBvNEjaeJxvjDhV2F
XV4h+FmYmoOHW0ZA9Az6hD5DxI+SsWCLgXN6PYCJOevF2IbAnFjoN6xbcxB81ytW
vzL3cMfWAkuwEy4DaAPHjd7NQNo/YfWt0hdtYrZI657/S8G3Yw1RRgezpWOeCPXa
mbdRyJ1q2XOS/BYA+PMMVlBMHeXYijOivYkPEuC+Um3bo9OspjSGyKzJtwZFcy6o
UbknEgwUh2BHciIY+y79khr1es3Qu14ZWCmZILSbzFD/nxZbNUht6zgwgOAPNTbs
kklCMaTkERhkD/vJnZ0EwflXtbA+OOz+yhY3su7w90EhTbRSTSYtCXGUp9NE/81L
EMunEyQ3IQzutXpWBSdjzBfNY4YaOXYdT5PNWYNlA5YKfGsgH7wNvcZOpUkT1rG5
ef5pzVNoiD7QVSVvLDbP+NvRGLdCCSseDoGtxyP+8nAttCZQRpMCpCqObROGQJ2o
+NpR6KUF09stbxjITN3YTk0tWr8JfXWCKg8AkK25ZWCaIzW84w8fFbGcbqYqgyhU
xXrxVnthH/YKg0MpxLl0mWP4041PTXBFe74RjR+uPH7PCKwFJ7uQCnpvQPvlv0T5
c2GVbqBeRiavzA2f5sUHOSc2JtG6mO11D3KPWt/sPKSWcXTGAxPVtPPI7JXXfcC8
GwK+SpfFYUAGtu4cHux7RP7gj6NuH2GThbSpDSU83kzisTi2oyhrJA252BDtWB40
aZE6vjQUaron6eyh8qYAdQKE0goD3nRqQt+jt464AiXaR7qfIc5kwdbbyN3wNTMf
0UdkjVv7fQ3Rrz0kLkkuYKR1L4T0qUtAFqDBhG2ElXhhwGEbZmkjERLBMIVk7QAg
/jQyhyO4ME1RiiBI7BKoj6KTicn+U2HonmgUus3PDE+hLsrxtpBQuvEz0uyN2QC4
LfgVEzMivGyCR8crakldM5wU8SWlYYJIXK9sgFPiXokCINCY6l6R53qCeRdezLtU
YAnzHExg9pQ2HK/XpmA+1ZSHZ2kB2ThF8Nke+9jSKrGlyVFd8LPAkAwqbPE2qHE5
vj3V0rmyCIkGEgKakKYx2lStHBgS0oevHH5Iwuz46bU9tBGeQ+ycIlzDnc7w6Dgv
g8rzCoPG+mWLPkq35mywdOl4lVZrh/o4n3Thox8Q6vReIqX750RKsPFypkMoBd2f
2BQqaJPu4IbnbkSY/K6Ae2LgVtdHpPBgvdc6sraH/RTDCZ3+yt9DVvLSbQG6EuF/
V/3HD30OMkIQ7fasicwYK1TxklYob6LXotTglW3CCF/tBjEgO95tYn3DVwwXTqeD
Nj9qYng92YYL76IVlQHYgSxS4VB7YoQLzKQhaOY8mUaqBlMRxNQh21tc2gdGmeAM
UltVI/cx7bnFCZufQvGdVddHGzwDdpHIGc1N+6APyKOB+sRfqPtR/dMduEtpcDZL
dI3fWE5CVDo+Psq6fWyAaFIYtuVT3Tra06jboLnaZhL5WY+Kz+Q0LWm1kCYQwAXa
sw2trhbssNbmfinlVoJCE3IIkp91R4PyAIAlpLFpj48hD+/DNHrhzkr1YUvm20/t
4NdsPpdA0bJqVVBWt0Mxb5oI/4ZOhDn9YlCDtBV28Au8b3OFDSJDfKcX+9gZRt2E
pzVHW4zG5PthD9aPNqQ82ShqEXcmg1Ppx2R3RpLCYjyp36Dhmn4ELM7BMDKNWRzg
3RMDGXN99U5+UrQnHRU1korEF2blCTp8aa45qK1n13Evlv6ujN5XFB8H6/TyQN2d
kacczg5hz/GZbLaWcJDF1k+UFlhy87uz/CGHjBwugcCWb9MLIFMlALGimhmUxSpM
YyAAyMUTVD06gYTYa0btRYDO16PplsndeB3ZZv3J9JnoKfMMwF/ynxkgAinAozrz
I1LI6PNEegfU7sT0MdpL392ovy2ULtJuWKpMd9/pFaWxfTWxMOmiqnSHOa3/lzmr
0w+4heLwtYM/QEeXKtIYRhOOSrszhuUWLYLbl9kQjPsakzl/GAupEYmr/BXNdPPV
A2z1EFx7BvZVhzkYAtYEGZi5RT6Fbscmf6FMeWBdDyrXNsJdQGrAwAOTpGNh34Yq
1eUlrMT/LuCE2/VcgH+3pvsCNDeBQt4JBVWMdZJF7RFUzPDpaoHcvywu+seC2tAE
0DxujBocx1U5tHBfwK3zgbl39vNxA8cAvj7PnU7j95XhQDhYPT4N2s5u/msE6bLl
gCbWcQGgM+tXbA9bMBBs7PxbwYKyKkQrfcSzkGR0YkCWjG0yMcj9sL0Dtmh1pUZL
k8Cc8Eg0he3+71S6NlAIctlZYlRQmnNKrfupINV2w4VFBfHDkV8fqTsH7ouThO7e
Y4yhJiefCt8itoAPYis3yNbFfnocI8lmI5uP3rkmbFJrmUThyWPLL3jhYIH3epmP
U1o37HSTpG7bRj3yax5tA0IOIVuaSzYbLomcMQPJgaDlcu1BZMVmBbbEp7MC+PO3
SBtOP2TB55bsEdO+UNd/WgWLkdwrwwkK1Nl/kVTqO8+w4Ej10PYoWS3GMtwvp3rB
zVF0S8l+Fo1jCoSgat2PIBPHlA5PjbaYGsxCJKgdj0mKDysDh8wrgYtSyX/ScYTD
p6px0ksnoEaJ9/+h8OHjEboElwEWrgjV+0RqRUCNwJeS5GrGFtxSEk1DmZsZiMJw
bZT3WQo8oGnLtuuQZgLNLd2VSKpC53CNXZtrhxsepq3rJdVxvelweMdiI4LKm1KB
5ytLR3nhG4TLCzmWFw3dAJ1M6g/ehQO/s+DasUQ6NCXwlHk8LtBgCOdwa5ovdZ1n
w+67pMsshyOFQ710Wi+4c9rZKBirHW2xQzWMtlKCQ2B3ZbxKsFiGbGnI82CROt/j
ChXPK8eGwAz4NIiINWMiiwmnlrPdb8MhYACk0tmE8HOs1XAgQH+gCsyQvR65W78P
p6v5URkZVRYI7PLgl25qd5EndKWfKz70iuj2WQ7Jr++O/XkholeU0M/vx8UGO14U
GyBIJiY9m9TGYAPIZXA7Rt/ItoKxX5hKu7JmgBSWPLcfbFjGeUXkPHquzC0dUbGs
D+k8SHlxcmDWDFaEU9sgVXgTPBPzrGpIuIFzJzrkAAjn0CMW2pWLjxiKS2Ok74Wn
fAr62TPWjWhLMwaSj9J8WLyLr1lLWIM++eXCBZiXQpdRIYuqk6Ge1TEzzUilbjqa
pxg16Q3a/kixPGmjWqyxUlgEgR5q2aPnlyEFytv4cH1z6LyJQHUJ5vnCwvFpG/e+
1+ka55H33n+b+N0wpwmARMFnhMd6cTUXn3tcuQ/dwiW7vnjaraCU3WgCctydnJVB
zDt/tid1ukC4fp97FYmS0cBYm9opzjf5b59pM3KuXZOH3UP9NdrIhOVuFmSpNnbb
uh2pabpZub27wLfRcdvr57zLnYSJwmeNbAauv2lgemxHfljcQTQsKHLjlV/aL4E/
x8KmAbo5cq6Ey+zTtKLiyRDpoPQlzDsLcWxAS9X7XdEMyuQW8nia+QhO3sLBoMXv
HJslDGeUGvLRVdtYDfw3vZcxxW7LUjmyCblNEtSioW8Igw4zQCQ621Zg4AUO/U98
ElvqlWXrgtHSJ/DEZBRl/TTkB/v+SSvG+CK899Koug9bRRNPAl/W6HrJv+2gYZbA
mA8PzJC8vKAEiBvZlkktmEIuDGWzt+JIMiWoN/VnWN5hw9HpCh364WxT6BxWPXSY
ttcfsgqAA5GHBHmgskxwh6y4RFMP9x7vG0QsVqIXWJVU45g2QeyM/b8fcgqArlXM
paYGAnpUdt06tG5dD3caSo5JFEQNdNGPW055CI+KuqFAkaBcr03Ig42HVYHeX0uJ
NKCUNzAropnnQ1VW358mE/6OXYMa7YRopYiy2vT6s9lCupl02B3kT9DNaSRWfIC3
P3GEyDJT4/a5hzKDG4TMV3LzOXIImvhD0ZRmm55XrCMzp9/sQEzJhQNGpYape4RJ
v2gHF2D8X8hrk7GiRLNKTdxuAhqKf6IF0KWmzAqO158lGibvk7Z79D94GPJ4xSVx
xH7nR3vHRNhhL28bCTArsWiVkxISkDya3zDftrL6vsLI7D9pQ6/4pjGTYAM0Fv9h
EPSZV3NDSJgrYtj2FL1H8h3t1sDsibHDPsSZw4bqfxjPSCcb82p2IFwxpEquo24J
lq+mi5WYperjnqQ0keXx/sdiNsgriDKAvq0GRKzB83MtaP72tXtXJoMqZUwLhKa6
rLirg4CE49tHaHRzgB8C6+5ZISfShZ+d98EiXC6WTiyrZ3sEiM6e1Xx0+mV1Tx38
he/fvcxtKHS+p/30D4VppAjajkoosVb24kDpiw/hJhR1yrAdPKABGNZLX3/p01Kx
oqF9Kao5hsYaLBXbzqb9OIU6I28a8DoYzgXwKimpAv3VUrbgQG7DvqDaIJq+wjbf
MbE6keeI5tahgptmS5XJmQAlShijrCiUc/BHR5At19Ck+VlGv8yU+LZGwiN+xBQw
TVjDLwChzkcUfTfeQRSwSvYbYX0dbj+LoG//MdfalkCank9Zphw8/simRdMXybIc
vuitojE3QZ/kxgw/LQFrgokzSVA06DyGGHKZccKHqRURt71Ruvwe/3dU5fPPA1zb
LVmT8GOfS0/nT6yC2+d2Qq3eD5IOBB490brmuwwKOC09ffca4zWIhbp/502QLOQr
7g+8cr+yEptaM9Uvfzy8uK4iSSrUGFv7EYs+wzQi/Z6kaNj0Lfl9zsNtVBxIBmSb
sQgrC98XyKzjq7UZKK9gojqqDxkSFnVg0B18smzc4FDxWU3o2qyTwl/0ADwCIPe2
5dIDtQzuPD4ZtPjfHoBg9AnyGVGYL315IHTiHlPU30Oly/JEIQvhmAo/h5BhwkPq
pcBegB+SMoQR0zyi1SPRcOxyDXneGXtn0e62WreVy4Yqvotg9303QB+neKKfR0NC
40jZixLaDlRlcLTu1bEiOFU6A+RbxFZ/iyoxSx+cuZ9ZoLeDe29FNCdESabDxjb2
81DLOkmpjSuWD9AU1LsVfv7JAxNViv0renpU/5boTKnVG6YN/tyV1BFh0f/HggoG
piA9dPuey29XFa3QIyjuyyw3vXvN7/G3to9fh2RzoaKf1KASMOL4IObpz5Zmd+r1
mD1VIM2o9OE3/X4jA9Nrm2jKeRVEKA6GjanEsq4Hzk+NKVcKYnCTLZXACRLaLw7s
GqiVRP6KLvHufvcrbZZ7cO4KMaC8n5vc/GKR2YoLEILLUMyRF9mVm2MqeKYYDvzQ
T6B2mShUoGOPuH+WqXlJk0JS1cCFK8qjM2sFikXRX9HUjYfo9pHMPhRx7ipNaDZQ
eKsHAoMcCg2ciR2IL0J6vXuv/yTdtxbWV79dxXrmwuoGVU48tLJfKNLDTqo6+S2n
0fOfkefiFmjuH9PagnMwHGD4jf6lcsa8uzd2rfqIejYjVLA9pj0QxyPUfcJVyiF9
ddPRxRM5QVQeZzjO40/YdMCMOZRpPMbDTSHCq/S65gXUoTJ6kFKULt9kbHyWtjS7
JAtYw/FP5MzpbW5uMEfUH9ieJRtliq7ESFlIg12yImc6KeNO9GfewfFtgkcPtY0x
4dS+rNEF6CHBnT3vbKg4eZJx4ETpUnhoQ2A1frQUvNuBjnrqTlttzrHNpNyaYYa/
Rx2hewokBwJ87oUexHmA95EKNcFGPdKkR5juN/bzuiVypRHLBpGV2VH8n/xdv+5P
iK0CCkauG+jg4Mj9hKQscEkRX+rydPsyDxikU8xvKUZzH/yZVCGpSbU1G1GOC1NK
eGv8Dk8udtBiiL14Xii25a1WZNl0mmRJAqfABD+YRlAxtFMuRZGTYIYSRIFhyWzp
/64zlpvJzYkkIbOUl+locUrPmfg169EfwbS4A79Qu7JBzAddZ7qY4b078cDbhewl
vVngmO7VWncS9jsyd/+mcA==
`protect END_PROTECTED
