`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qt6j3HLcltSTgOVQOpaFkEUfJccWy9dLHQhlJ/Ztp7KtMS7VfbwqUEsc4onzW4DP
91kdFqe/+Vei6rz05cfwkSZJhj+M5ga01crg9S5vSALe52cHJLbNM+tpQOlGcIdw
U9nmh1VVTvU19zWhIgfRgmhXDC7LbnS6po/50ugIlUT4AQMA6ecuuyUk2nIc8mNb
xg8a/xIG5m+pB2Pjy+LDFK7j5wojEqyelgglsBLBSWZ1+Vj9qTsg4y2NAGroQZ6T
olmDnPl+ophMGnqaM+YScVcuwGUpg5+Tgv7s9X0I7G/MH/VokFcE3y2eJnc0cX28
ZHQGuctrP/lg03JpefIWFMIxciTh/wxO9yDVTw90OU0Rme5q8FifOJW8ncU2bYrQ
QD4bwgVnjdTaQnepXMAnEcmkjURtDW3QQMeNv0qEQP3PNG8Ezo5Wgmrj4gYlc7Dd
SM4YuFY63YJoqQ4iNVpiSjyRaaLNc+tXQ8FzRni9fxYMZpqD+AVVBs5HHIhUMXcq
oN6I/ANcSaB47b6C79JMrLHPUxt7MkrcjZfnzzeLORblvTPE7b587qSUw8RwqRZX
qZ4cwYNGv6dxFDSCtwaQoxgSzQMJ6fBFMRRRKoxdfXv1TipKq0oER2t7eSWoTKZg
e21/b9oeunW07zYHz5/fkvfY/fc8EOCk4Gh192rQgUwW0S1E+tz+MpLgJhMUrWMZ
v7tVXdLPLByuMJUkgWgZDMonNcx+Bn2g2HHvTS9P7zYVwqdeNuIKCh5ow0ojTQ91
bUvJVrIkNebJN5aJ3Z5xI0t25o8cvnDzJAXQ8u9M73NkGkX2RMc5CbsqdME9XfAf
TMV666y8bkOEb/4atqLeR5/7EYDuV/28HQNfaE28BraHK8us4+ARt5Me83B+8W/Y
E+k5a99vrKL1cEN0e8P7wwfNDZdLMscKvcdMQfIf+Pfs71oPXy+AL1XUJXuhrTPO
`protect END_PROTECTED
