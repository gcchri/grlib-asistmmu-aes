`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tkcb7TUa/WDrEHhYVigQCESsaf05n+a/LZAY73XL1HnOOCZPekE7XlITNidKrjhg
d8eKIsGa7M0jeNRM14CtKd2zeXVN0aLBsiL2A2FpcaLy8TrdD5F6KVPhftwCjmiE
rqLiuM0J8dC/5fWZC3XxM9PEDCl1R2YPaPykn3pkAQl6ZNSD0mtcE/qlfy1mpjot
tWNfMWP2ta3uiUAXsdy5HYwgvKggH1DOM37vfNLV1eKgUiTRhpCe1hkfmJSBOOyj
ZCeYAJC3OvZvJ2TxIBB/8AD9kEvhWCXDmTkOfaLkY0iQ3kyWG3PKTsgQILdIb5tA
ZfC5pNT9Dw6Eq4TrOwVj2rZZAf8br0Ht0QlvwY8fV0Vlzd5Fj9Wn2SuWbeWgZzaE
00fv0K5rwwgIWbI2uFYIxw==
`protect END_PROTECTED
