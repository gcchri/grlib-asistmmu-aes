`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RUyAtXPnkSqsJBUe4hp6Go0AWnvb1wJZWgXnN7gDypKkrBMZpA9qStfG9H8Cghvu
Lzu/xufs7BZ5XFMHxsw1Grz02ZELQgr0arb2cT+r+uvsP9IJ9PmmBaXW4lQsyvGb
Ed8JI3SDqvzsLZ/j/7sTV2DST9aLKRsbHUHaHCZ/kB/l7n5gIclrFLVFaFVEqGIB
cCuN89wKb2onsK/vtIQJGOnuM7LoHsExgUuewYPx0uyxN9cBSTzc4GDwWPuPi+uO
XJ8Cr5tjWQuawFxJqisYmfyFkTB/BIitdn1q2XdBExOf+ieN1m3MWdBmBQLM9ifW
axZHZ4iyM+E/Fl/rJbewkBMoGCSYkYO4Q53kGqz+b5YJmfVPJorEO+Jy0h3RWMV0
nYuOoo75/q9YvaGAcKax+nOGZFKBHIUzx1N4ovDTTBe4Rm3g4uQk5HCnsK0cjwd2
sL2oUebK5qRpi9C4jLCU7S24wIx0b3bhVGIdiHSk07U=
`protect END_PROTECTED
