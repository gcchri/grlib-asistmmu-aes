`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9odHNA3PXxi7klHUXeeqEzxC4tHbaq4PEIYu1hlTvkIeT9P35KXMwAWHHyfQc/d+
6drXXnFxNItCiDJgQ2xuOiDPB53cvtOZQJkghNIa//G91M85gdFsUy7C0Ey/7xoe
MAkq1SDrbQEJXcXkPMupaQt5mNvFbHUi9J9RnRuzFW8JqSewdJ01qMMV3jMkbyac
EXdG1ujHTiCIjz1b5lweCW0U9xnR2doBD7rgS3QSqLzlpl7plJ8C4xjMjnT5INSK
5bwJDPxar54CJFqX8SK5Ijo3Ja4MyvM3fU83yO7J9QtqUXyHr882myE6FJxuGZU3
uOVmai5ECLmiYFeqdnlsMvYMskzCh9yjSGvjX/3FzEXQ3aWo4837IReRriv9FFgT
3EF0n0SBagX17RAnGi5Q1LXIQYBULTQzcCvIBp0Kpe4kh3MA2uVPj7ZTiMd2YOYP
8ykFqEdBDnUa/h2F2FXlM5cTVNnPAIHpVt5fUjppBGRiR7qggUqOHMpfKEp/GOYx
WX++UiBoZIqU+chkNuu+7zFZyTVuN/jNQFeIPr07jtT0YODGtC+/BeBEkJssIm2l
bdvfzHXpz+LUIfPW/87Iiw==
`protect END_PROTECTED
