`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8kuN7/LnMhusnj6Ntza9LYPXsogDCHsn9gsJtf2jUfXoF+kbunevk6qDpR+t3GG6
UK8YNeUcwjhLg0/REZH4q/cSE92osDvEIUGNSYkX1eq0n3n7BFQB6x38EtpQGnm0
FZ0ZmtOfOj5esrEQsiMR32zCNA+LQMBizyjoFO9TJJjU7xQwn2bea7dRPA3Voj/Q
fyZ3jSsp1h4BLPaPYBS+b44mFFWVJHE9ao7lchMex6g8r/Cyjzm5Uw9VMNanlOz5
Z8tCFfQ90dpB1/jXQRw6sEI7BVQuDkjNBrpKfv4lqbJUJQT0ckxX3EGUBzVJNqTX
PZ8o+rpbyClDQY/DPztKau8ExjmXNibaHEBsbX7kshvYAE+yrraRNgXp9k7xibTh
aKSTije3n/Vf7bFLkXSeq/AFupuy+a+7DDRpPOANKUo=
`protect END_PROTECTED
