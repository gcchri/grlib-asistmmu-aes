`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eBLHqGgkrXoF2m/h5wvW4wzgJY33dBqYrKrlxwVp/QvtBjQK4IUYgjIo4MGvrOB0
Ob0huynrx7XcU1fiPojy/0sGz3jPUJbq0mOxc+ljFi0U92WmeGf7hySvbsg2BpoE
/tv6tHbsjxDEr1gSQWfu1TERHZ6Akatk79vDcEV3P43swWqDJlNRh76feBdyA1Kq
wa1gR36JLF9K6rvmd2MHHs3618ajSsEFKgo71WRAjczmCHJ/BhkCO/rYFbyvvQhS
WQrZk9ZlEPc+Ov2Td96C+vHUpJ9+E3gSl39w7dL4WGqO4HUzrK3sme6Eb5jZl79C
FpOP9nysGkokWvSHBcrkSwQ4gEaaavIaNd5NwGEsL92vB2Ma0Mgu1T5B/avigwpy
GqIE9gXZ9FMXPKXq8ruUSyRW/6TntTw85geA89Ilv5vO00sWuEXoLZXJAm79+pxv
HHRO71XuPwOjNmGTqHcV5VDYJfkHDkMjpXwB63N0ucm3RYczlIwSvn1qOvWhDwsZ
rlf2bRB0FO5AvlMxbR8xAKgegDn8AY1UpbktGD7yzqCSY2RVzsRPDCZOFVkiazhb
uJpCIyFPzUQI1ueVCnXw/CU7FNu++V5x85sNrTREfUKrkDa9jqfrVU5bQ2azYl+S
FZ6VUj2hc5HKseoNHsKwItOwfrrrUT4PQ35lqb8lfTI=
`protect END_PROTECTED
