`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pYmwIJqXpJSa6xw8Fi6FpVj0GvFxaKDoebOqgHNChBC7tSBwlLoTfe7YIApbOb37
fBLJCGDx/L9VHAqJIzZg5cqbUfBNXPW3tpsF+r7AmOfiOGmvzjv8ZWUxdKn2hJA7
sIb6eqivOcJ4DfTW6mWaFBV2/0R6EUJF3ZUIPAhnTQ8uDxWMl/qQFHNviG/YmUks
8nVsIkb+sgz6ByhPbUs/sqNPfzgV54HssssMoaYNZf1D8CGMzozR50irqZ+sksXo
c+z2vZR+WDJoO95pkKmaXXLIf29WbpD2cpOzHSrn6I8CKB3FwoAgHjl0XykuD4Mk
idJ6VmP7tolYa9e5oZUHOw==
`protect END_PROTECTED
