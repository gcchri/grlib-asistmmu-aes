`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W6B3TdqE6xxP81ErWOoWBlNeG6GvzMx65S1o4LaWbz6HvCA0fE1DvyJ2QGMA8m9s
iLhPQRIMo8eiNq8n4/soxJZpFHuwwx4Di3BA24wloVFLPLAR24mM+VrDJo4pqk+T
z4Xr7BUC7CVg0/aazoKaPEuB8TGAL8WUIOtRpH4WxUUsdHyrYWEs+tzJmuwcpTeg
5LUaBTqRcmGZfKRKgOCFPyMBFMp/bwV81rpqXjNaJ1oGFYDOzf1xh4EMlxxFI7ng
j4mWam+oBXqsgCBOGGtT8r2KHe2y7oBHrpwiGbYNUXeo9IZDAkGQk+fnz9BsRV6u
pqOZ/jTEt2ppRomlFwvlNjS8Db49nW5X8hA4jElqIoUm5ZTJLnTIX4BkpNMUWgd/
E1tfTsIdmrhEZVioiceJqIGATjXpyAgHD21SRqJ3fmccz6yqzNDojFRGsLdBMI2g
LKgc06yK0n2PWjHDP5ItMjYYtnKUfshxdVOs11jUcECwxbAN8pPdaJtYvCefQCZ4
T5wWCrH8HTz/iKHvBmoVi/mpwRWAJrJW2c1xpaTNld1Jvpc9P7oQ8t+5Dbb237Vp
9wPT8yMCh6gIQ/fhDJVCkWMNapkgGKDQfhKAsEWtArzwWbU71ZgsVa3ZTrZZqGZY
5ATOudjgC+FWQiBWSv4WA1A7MTgiDuqVJGV2g+4DdQG48r53yf11yWSiBXKxHAYB
aMJlTcy4NxY643Yc1coe33eoeMjfw57YAHMXYoa3VWJarjiNcdAfDFu+VtrveKx7
aeh/ZkSl/4nNEEGkCFUmS7Slu73l59Z6/t9yDTl/PTyygQqFnFsn7j6Er0c6Rf+S
ZVF6U0ITUKBV05/PVXWFF7WGQzu3xgPYkl80VNpErPcRQE9hmNn/i63Vu1prIR2q
uOeT7opoA60ofWyi2OI9OMK/YYZsXrZZN4HTXgax/vwEKE/qatjHaIx9KZWUYAE7
uNE5f6GMfbo53wDd5yR1dtwjujHRZdZ2Z44GSJJ71eLAr7wGDSollfIc3QHNFdIc
53oulDQMCIbowbkGy+Gva/Rb9Mw7L9yb44ZnQv8WpDIPrXpnx5uOlBDKUHSTgKwu
XrmaKMDWVtVA1oByuMv4clJZsFFUqyK+PvKglglcFapr7lhea6siJ4UkEX3Eh+En
7Xo8gpy0mRL6cD6LCtFCAglcZSDS3QwKcWj8ajQwCwYpwDgviKeTjzI3T+piLylV
ev0fCWO6P+Jzy4BKSq7CdSrIiJ819afQPtqEG43bYRfAOf1VlBXgITWPbqZSSScK
RbTWZnPR/iswOazvEDrR0m+ViaM/yDqU9tWC4QKL8eZVrrhGcxcdma6wRZ8zqkLH
9x+S7hbcClca8KNK0wNfnRtTPstbPVGJDJ5+sa0Gkl+FOS+4tALNpMdwIcSo0mGM
eVyi4ybc3c+utwdlwLF2YMB03YUq0n/qMJlrn+keuReTM5tKIUHT0USde0atJK4a
LQ0bqB06BPdh89ZpF5wi/nsx+A/nLMo4PcMRVoTJy+NoskHsZ361luC1RPMDfUrl
r6VLZxsxwH+lyfv39Qn1SRwV6CC8Fv7aM9wZcIrTtvDkWZecM1iC0IPgb2wK0nVy
Ol2qv2Dy6hBG1AQm/xd+Fv0lzzStJ2AOny5FiV3Agws4c28A2hyR5sAiSVBhDssa
U7AxsoJftDz3s6rVJmTngcmAahrl4JYdTIV08tpu+jAYZs7YnXyvV+u0Ggb/Ndtl
cVK+tOm/w3q+0T3l3YCSAhi7jsLrqLrcGufAPmN+pt54cY9F1LqkDraguB5/R2+L
WksXTjcWfGiahCwlDgLS1DSH1Qjalh3S/xSxVi0OhvF5J44ImCUj/79yeF6dSmNM
uwp4OWNyMLEXe+1GdXdh0w/5HDvNiROE1kSBZQsJdC1d+9bOzNW8unFJ+tE5TDD0
zxG8kxB6cFqxCA0Vnf4Go4iNus+cIPmTY92+14oPYDkywNWB43+1sKHTAS7bBhqX
RVImKjyimI8JkgEtKoygI0Ka+VJIuu4x4x+9e0oJS6/gHQn0unHwyqhEQxbb5jVl
9Gli7w3+wBOlnpnfzy7NxfTOV6MqYkh8brr/Uo2s38LESmXBLwIThoc+rBtDEPBQ
0PUMQX0qG55c6Pug0gJaYyokSrVSOgrIxlCFzS1AsgDdxnqjEm+aOjZWkjNzA9Bz
pWrqxi2rX5UC5JnaUcOxerTRfIfi9TEapTkKqvsTCZtSLtj8ek3W5cFNdjhq/fbb
g0RaJEZLhu+JOt53MaJwLmG6ugD3rXVMlBk/A4IcGhsq8Z+DxVYh26Ena/gTIdeA
wlBQ8/c9S88ju3Go7FHFeh9yx+7XDIx9x/WNTTIE8SIBpjs8+SmCJbM0cieJ2wSC
2K6FzYKbsq83zlqYVT/UDhwyEApEBBW83GepHnXqKzFTCJkcBe5U5rsRK9mt1QRg
0bYyro6toVm3TXaTkdNEChIqkc7GxYsxd39NVA+CBtYuTyFdTVdK5aPAgLvSIdix
Sn1Nxh5xMc64uFOhA5pUElfCBlLwfIi2PV9S4ZPLDAWKjC1UROXmAeEI7H+UL69o
rCTBNRsb2OoY3/C+vh7c44vKBNcYATk4mBUWjydd2vC0lGOM+iBFdi6iR4htRe6l
g+b76hh3/i+QuOUbswEXUyFuHstGTzpYvvssVhPYlPKju2huJKqSGFbLoEO70loy
BwFZ4bvn3D33TFj/P9eTMfxUdpSzYcZeEHDft7Cu+FOB6KBbkZtEpXlI5x1FekEd
hufy6n/mJbO8G20Ab3JvsCvBv5q5I9zbXrPlTUTliWcSwydiY0rbnQKis2dL8ydo
PbepjlnrscbX+SZkLGpFtrZOW+WOZ/xAq+/Js7nTdtSJnkIaE4iRFfzHYUK7/kpx
+LnbO87rqByrbv8cCGP4BAe1hSbzzc0upHh7aN/6Zd9JzH5FZjKj6pPcp1kRQ96I
buCPMIVrNKd7JJTSuTNbNkjhvpFwys9OeAcqOBVWhgM6A13/MvFCUPxXU2LDqa8l
1CUd7kmSvbq0XAglHyhLEHAiBnTiJyS4gUuF5WqcS1mdaVmg/HlZQ3AD8zesbCDM
FrWthxIfv/4KyJg8SNmo9mRaH9+p9mxSMQkDomwubE0wvM35Na5EoHhgrN6aMCGF
0cdmavnA+p0l7Q2eSNj0iXkAFCmchO/ZzQuVp4eV7aY5OZhYvw2Emss16u8nqJBR
JU+sxwkTXjB7IL6zbsl3yR57ZKz7gS1kNeQ0xFl8PpfHdu5XAyNiz4zVqi/YxaUK
zLopohXR+3NleiQCeh/EJVrfQytuAyvmg7h9Bslrnf/pwEF+vKgSHPKzuTjvUvhI
myqeHYPUXAZLsbYyFMJaoBeN7xgDy1kpPXrLH6BI6O4TccWK5fKmQDIfZDxrvHoF
0bAmbWo2yLXed/6n3AyqGBzTKr6PS5dfIVaHfkXs5jvmDn+49OgK/SyextJyAyA/
lqTCrSou8KyfvJzlL9pwZRwq0cksI1OVOhtoyXOJtq85bm2kiQaNUVZLRipbzLRP
j9Egh6uXBWoi+07fmpIgnwJYbiaO7Vuy8bndvMW4Q1S7jBSXKcd0ocBIDLwmIjGh
Sk+W0lC7mJ3qsTvgVLNfb4+2ZCamtNCmLfGxdZuRjEXsI/SKdW9tIFg8EOxO4UXh
hLmOHGCmtYXvfV3NJiDf0Enu9fVSz2uT0f+EXys5lIyy39OBJE7oxRi0TdCOnJu9
nLN+2tT1rUX6CcGU8ma1h/Ptg8zMXC+fkgJn7DvV6/LCrG0aV6XDxliHcaVZw+PM
mxPjZw9vZmeIRQOMKFoIcnWtYdRA9zqfRedLuBb7/p2pNC7BUdSNBB2s35aodOoC
U3gfcZXUOcuJvo4Pqh4cvf6JdR+av+nGmjAhGsSuvWS5NPV0nYocy0zigmFXS6al
uRS20kaTuKMYJvbeiQVnJbXtgdhH4bUAYomSe6NN3o4n8lgT+SqvjlN6V4I3dGAT
Gc+fs3Jmi2eOUAomnC+ftfu0eCEvI1UNd9tR1w7ZFqSvwMT80VjPvGCM4wXB1hA0
HXX+eVBErfRuKbMbMSKx9BGKTBLCB4IfzX2a/UIcqHDRQ7YplU/+EkiwRmwiULy8
QK9I+A/wwI+JBnAT6EGLW/G25XYC40UqtXwhQLXV/UEO5EBi8WS47b9TMf4PBssP
Usft+TmC0QPv9appzG0IhE/ethKqifQRtFe4XMdSDQ42ZUy/1U1mezy0ng+ObOwi
EQjxltf88Zjl0pFQespxFCu3cZ+qkQqCHaDUmJ8nBSzt7gqW+q32EvkDvQT+F68g
yWxKHyzbRRRUJREh1UaOsyvxx54pnSYLXDkN6lIeh96maGbBtQ8b1nLt8HRwI1uR
3FITbw1n3sJxewsByNtWa46gaVnKwcSP1F7C687r8bZb/lGg38EjPN25EqpsUDj5
elQJcPQBjLxYTkHcrzskr/8c/gx2npRCBlixYnw1TAF+mUYDIcDGg+juG6DlbdDp
YIwQQyKuaLtA4JvET9qLyZRnJbzTqD33xYLD+aK6NVM6O+UAWkUTJqsWn2TGY3pR
alpOHaAcucdGMJ8eN4tUgxZxQudnu3bj7ljaTloxwNIHy1+gIpU13ipXfw30ao9k
rhk7TUqHPqGTPloZ7t+XNyhIzT+XucXzzGhgBj7sXvF9ZyMFKLOGaEkDw/gVzIG2
bGxkqQNthBFDklnXgM0eWlQK4tMCT+OEL/Dyo9zsducmDi76gwLgjhlwy94WOkcO
`protect END_PROTECTED
