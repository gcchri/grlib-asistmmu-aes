`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kkVKRaE1ltQ6bbCAQvB9nt3ZSs/AWHtOP85k7THfU4KLy3IeSuZ0LEi0aYqGaY8x
S0vjqaXSuHVSW8Qczm600oltnfz/V0eLcya78q4nW5q25GYHqZXUuFwc+JJyQJtr
yJvoc/5CGldPie4HpmXJLhYpMv5iqswHFGTd4Hdqa1sEbSRixjDvPD003P4lHBmU
3QJiAtVq3GI1ogQTvXD3PBgp6Suh3iRi43ekHpJxkvhbljsfJ5OQ0LovHHljoeEN
Lj+FlCllk03ga5cr5m9QGxGzEwQAkpP/WURhCynVs6fOX8FHQnO4KUoAUebx9WE7
vaDnliod4Sbgem7DRdKoWYf4gFKrd1aKZ9spbV9F8GPmU6tIsH9K/uUTZyfkUiTo
`protect END_PROTECTED
