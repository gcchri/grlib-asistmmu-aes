`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6hVUeaQiE9QIR7Z33tbxLm2AMoFlmH20JFG6UYF8uxTKdm0kgHVe5NYwBNCoF/7t
NzhDWOm2JkIpbHMiOlW8pKYiC/+kRYv3tEHdIlU3vRAkvlhcps8kDDRCRLcyUcvn
bVtxXwAMqQ4HLJNfF6SHl0PC70JpPvrmVYyEiVX/ZkK0QEkE6PswN2Ilc0pfuMN9
krOMuFjoxC1s4KpGyjawKeF96ReacQDD6o0pLvZmBi1vYPg4iYWkorllFia+B9cc
Gz0c0/d/gf4aPqSrNC3Y3hOBqrBUJksc8+Rl8AbfaiPBZHBcZFDNRO6yaC/C0x6S
Hwmwuz+tEjx+gDVPl7C/aYWd6xUWgA1fI4HqKc9bT1zIL6ndz/l9Jea8QogEUHf+
qUWe7c8YuhoG0hQeALUBnw==
`protect END_PROTECTED
