`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nnZrJKZzNTA7uP+BFirQEQ78lrnYfYd1Qo6i+5iK4PunPocKT7K6r7+bzhfEs0xU
p1fTP7NX4WiXd6b5oiw+beOlrzSBezDNZP5/9DQ4C/g1fNpVfGJX0MxboZ7enFeY
hwHINJN83OtUdEsZovcEUhypM3nHxQklF9MjMfMKJdWYV+GU2bJiZRvyvJsFo30u
s7m15HO1rI3KD4ZZmiaRupaCeOz5BHv/47eERnPSEybVGLCkNMAR4zXutnI10FSI
BZVPpRXx1GTxh+n6gEUj65/8l1ufsGuDmmIOPTA8cSZdE21IbprFdSqVzNqK3HhD
Wpv4tmecNEEzb+M3nYakw/1pc+eAerQFQpxVXvqaSOZ50gWpAUyKFEutfCN9Svy4
kkkdF85aEU+flLRDL+Z+4ZqtkDniBpGclDsl/fG7R2RmrF3AqMl+3iWKTUSUDPv6
dTAR4w06dQ55VoQGn8UybVM1LLfocs7YQcEauA82d84fC88VviZnfcrVW1YDx9AC
6cPXXWX31OEKHjr+TyldDrwNLzOjf116HsOQNmMc21X25evQnor1HmFWCFsTwRST
pta850k7Un3HUsYDbWy9efLVOojzpNkUiSZcqftWr63d1rhcPpQmKbsCrMPk5QOd
OBozX6Q1eLIKkDO5gVh3JTPKn27x5m/JJK3g6Wyj5Mzm2dL+hFDCo/jchNiTQ1Lk
4Tvr/QTtgmdmiABAJBSX9j7z52TwZ53QU5319Qk1V0VegdjTKtROzjFISE3mzcD4
yRWARPMbamTTeff7A7IdFM3UN+YaJ+lfL0uuMa8Igc8qSkMdp5y1c5MqhL23RKOT
FqXPP3T/IL0C+JRZmRsXjDT0l3zqSkccod2OoiEFrWPdwB7YS7Wg4yh/hUzLo15L
FdDwKd423hB2H7LqceGrcPIR0QW0afxR64J+5A5sTen6hYMAk/lj965X83Tqh7PE
s15N1vmZ+gQggFJBIFQxKWB/iTFuwea3Uam2xRDQ6sl5PI2CRTtk+mb3hnh7+RAV
bSmJxzlljly9AwEbJ8+ogRKLR+F4bNOCNyVIlyM866a4N34/YlTbEasnlbJeDGL7
bDeCorYI5mXWpHSEYPPOJU/q4eJz9m3lhAHfYKKwB1+Ic9MMZYPLpBoZI7LKNyIG
mWP/D5Mc86pLAJeDIXz23RjQMxgzv8c5ABHed0QzdDEvWmmAzehhL7v3VDA4VfQK
OUUbfVgnatl935aMnOxlSzUd1tKd6Kx8Twjb0FnmLy9wXESHiIfEEouA6wnsiprL
/GFXwbQEca8AARbnjx3uUP4PhhOo6BWw7s2zXn1gFDBTr1VITYpxgh/5SYB23RPW
0S2padcS1BoyeTXbZErkavKrTsRiWMzXaCvlql2JM2MhIlPowwy5CmItYL8TS1H2
rUxKSy73zUIJZTBxvk3n4PIOzxlWgzv5E+x3GrgzwUklpzsiZN10cUgORBqMbb6r
hhye6VJo9G8NUylnOXmD7XQ/Scp9T/hbqatpskVHTwT9YjqWrFVjD9j03xMGDL0O
CrllnGpshW5rqH8bcxJqK9hceFlOHhsBMBKbMMyj9IgSvw1eXakZcXBaOix2WzCs
gTvPg0rkypsLrLGuW8QVX1Lz2WEmNZ+kr0BbB/lBHTMSkbwHq8BeJYaUjRh00c+P
zg3Jk4F0eXCI73HuigJEUb32jRapc7jIkGaGDgIANlLiZBjJvJ8eyTx/Wh+dUFRN
Ij+DWAGwQv3AVW26y8E/Vt1/NjeHU5rrZQyTNvq3NWlnKwc1U72q3vNOAsqSTy8g
i1mg6RLqAvo9z4sBQWu5DAU2vX58DIAL372Jf+fCFwVkvSfGH4iB0I+JqEP9kSFX
4e1i+MNess+btZO4RH6Tj0T3B+Q9fHlSE6py0cir6mxnRZQLgFPrcYqXfz/cn/uv
59mcUqCpsOMDPFvHDwysvZdp4uLc0XU4tYob/ttd1KL36FiuHl+k1Gj2nbW9TTNy
y9b5TnSqbYhayna03yLsM0PgtMVFcjBZaiAIQefcBq05VhxlwbAAh7P9sqjH/COO
fdP8qCHFoDNDbIutK4tfFfvctuToXHIbBx7eI6ukVy8=
`protect END_PROTECTED
