`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0aQjkDOZ78q93jiaeu4jzPxjYAQOoyx5b+Cf+uU8H+XclESa+IICbUbk4clUt8/i
FqS1k2ohdJoSFlUIj2YFcOhgAwdG2ssvDBa2RhSMVnS2nYbpMYzGtVONxG5XXhoz
MyTTUMvo3m/YyXznGBGmY6BlQ9EvP/XWFG8ZLykaeaoMyVxuBniCzEJo0Mq2Zt6w
Beus0bwnLZVK6W664aFI4VKzbg4ZUFcOKn0x22duuMc9llTkvlVKPCQkf0g0h/tT
oOEMv7fr4tGZJpuAfGw1Pg==
`protect END_PROTECTED
