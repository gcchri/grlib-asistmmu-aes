`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h8wHuyoB0KsjNXSw+J4LHb2i6xTeZz2BqIELGiSt1wLBofikKoaMV6XS42c8Ms9c
gaedFsqgIyXrkFst2WEHPZXWrBGhryo4FSrGJoU/HEaRjTy4VI5KnT8t6Hn/6JUa
QDJBmMN1pioZ/PNOy40EpKJohFkGCAtfGTM5CmhXil2rXTD1ooRVNVtGWdjU/QBJ
QKUQzBOxwmxReLdpfBg6t9Drn2NtaGvYHkQ2J7CbU8iY1xhr5WqA73XALTw1rkuU
hYuvJnTFLqa/EzHVHCHVMJmtinAh28Hj6/sXRQsrbsY0ZdPCEzy5kwTA8gDr1MTr
fMrULkvuWEHuyyb818f60xP7K4ywZ0Pi7A+sPYhp+BQpAgXvg4r5aa2T6Dk6c2yP
OhKsWZCiwvKIfO2nSpYKqPOPk68w3+QmN3P4sCh39oBk85u0amXkB2fmWhbqD9tJ
DqMyBS/yLFaZnApLS3+30uzpkSgI8+hECDe3yGxJJVWeiMAyvzDwr2hOJTau01GM
6M15N/ceMmeeJcxdGS37/gL/+c2aiIlU5cHe03CiKDj9ZB+9kT1G6Delv8qztJ1B
biwF8iUdY0hiWynmMJ1UCYXjlirB7bIAmBAi5i7W6gs=
`protect END_PROTECTED
