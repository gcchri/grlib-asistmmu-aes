`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ubttgG+JW3Q7RWutOsfGGAfGF8+OzRmeUiwlymcK/IfBtK9wQaK+PJomtdiWkaKE
eChmvLEE2tzoVGwV+FVlgL/k9sqlxePYGwU4wT6BYP60sf39a/eDJEWM+HGPunJb
UVJVEEzrFGko/IJgL1GMCjJ48j0ZKF+rU6BW6vuCgf6Bng+l/Z0tlvNSiX1qidSc
WSgIW7xIIA1R/uFkolIoS3Z9ZYDthxrxAb1s/4ul5CgaJMwdVrTyuStbEmn7ZPFP
1Tmo3qYGXyGmvJIfG4M4LtIsvSx8DGWHc6PGMMiFGeI8n//9e+DyKucs2ygmKMLF
S9QEKYyv0Z43SXmPSLHBmXX18zS9qINBO7yqCv4bu/P94U38W3VTx5yKZsjXVfrN
lXaRIErk2kltBaMXfrwsZ+RPlqDtPDGeKely0RrtW8t78/0AYyxVb0AQnSgzQAwh
67zrpKVH4N3WBLCx0po2dTXtneXKNqdUJMmmacqwTeZMV9GXMHxJM4rZw7s9FVXn
eJxP5tPxi+DhIL4cF6lcKBaap2oj9QCN+YtZ8eJZBju4+6RICCyvohrucALM9i8f
0pE17nwxmjtoGAYbMHNgL3l7oBMlk/MmLsq0v0WiAUP9psAMgQ8v1ihFuEbq3jUD
uYsLX1nd/jlkcsRD6CErl2qbZAdHy6ErPeHFJHhzlx6D6GsPTylE1ybAThMiaGWS
y5vBwSMFtim6kiTgp1KzxOm6A+5wqGaf43Eioulyt6FGnQ+50iHWchEVk/rXYfa1
dptDLOwaxUy7KQUxlfHlfKnr47N6C/uvJ3bONJtULYnZxH6XZn36J4sbH2yChKv5
aQrxvxIx8N9Cxs2RbbfrM/EwawBmV3CkHOE1zqao2037kOKau3DDpVPlO4JNoecH
44H5V8/n2Q7qujdPFA4oBDr8HpO8JCYlD/qgXFxsPmofztHMwSQDndoQgTsOAicd
YKu+vTYtLDiKCTelHqrr0484YrGKe56hS/BgLTKzubd2xGdoVvh7pbNgeZQwlA/0
yTNQybmcyOtGsFGiMHvzwFy3uPZoe1tKKZGPs94hWsWlFo711clyN1LkaDI2T0NC
eqCgnWV8CgBecnKoYQkq1kG7zTiar8AaFahfYm+dg4TiHR5uraqFUo49B+NHB7o2
7cV3fAXa3s1skQSom3qpB7IBffMS9WbgN8Ba2UEAiRSW06dkyXo9/sPCh3A3hR7i
1GweOdpQ3D0J/DtyBYMIvCioCFp5s0AVsjKPBXr7TwOhAP/WycaOKd6+v7pWY5SK
sswRRaGwNUdBbK6CnZCgRc7SH6pZZykD2RikSLZ1yCkpMZ4WEJkzq9TUgK0eYf1B
14uZKY1eJMKbVUe74UbU+vCeFc0yMWnOXuYtRQXiLleHFqFgYmBCGf6wA69VH2M7
rIl0/UW0VBYaheoRIIRDjLR2GoEAJlajsvRr4O8psjfQm4re0XH45XNUjG3M71j3
PxVX0aTK/Pdv4SAvsQLwIzUFAja/Q2hY7FX6oftnVXJkkPW4nWu/01IKUvjOsy1p
aRZs+LB+LNVUT9Vjazb9n00E1pN6eW+YF9RUjteDw5J+Us4F5m5FzYdFxP0watUs
XlVh6jBgFR/0WVnLx1QnVT5rL7iOcWifWhvdGXdMVUncs6RNHDYZppiZhgWckva3
p3gUA8MZl4kXLiwTLEvCatN9RSRe2hxMLzmQ61eUx9cV1EciCM9+thiONgHMlXMi
XvKN8RPGdz4L7NxYZT6wL/QlC0jv/ZQ0hTGPxm0FVc3/RWySD5Vm8tuu6/FkJTfi
yolyN3qzeDx2RJ2TUCVP2NZ/nnMbJa+vJNjHyEMc3G5ZiZSQibIsXns3Y8y4mEeB
k1nb/2D9VHSzjFObPyvIgGcuixGSbANoyB8E5AlYTq+25jV0RD6+rPqoF00bdouS
WDUnTVimIS6pOi3vzydTdJxcK+w8HbTzrROKQ2LgHgo8mKlvPg0f6KW5SKlrQ1Tk
QRNSaaU8Bzs0sXtfHVznq9p83iiVunj5VbeCk9gQbvvQdzWHmBCQnH9qvNHtliyf
otScctwuu252LRrzXU6URoYjmSbHfzbXgv9OyU2J9iHeHuU4Nn4WoI+VOAmWDmRU
KtZHgT9gPzGI2KyLQHOLUAVauBerfjSw1W7aGOfAvFA1NuduZ5IHD3B8MMa8LxBC
SJYhcpbuEK+cHDVfuaXqWJ7BNY9iVpmhcA4ub+iyEWiWWs9rRihZJ5ylY7N8ilo3
6bE0HxC939dCtP7zseS1h3vXKXjLLwENW+KQSZjC/yTWFDPC7ttc3DGkMMScWNoT
04if4k3FIPGfTwqlqJp8hu73K1xSZy9xC6Pm36UEKxRoFXFwTfjoXf1iYSijD4QN
DFjjbczXxr2DWS7edjDwLpD5vO8P3KMCBAekp7RzlqQ4eXn/xYBJwIcqTFkV9pRO
l00+eqO1z3fOhFLRkqjPtyvgweui+uBde0WQcHjzP5ryJBZn0zcN3/YnHkZMl2HF
2U2RIZrUZ9+Zdkm2UvXgFBozKZAXMil2KWarkU7qj9Ud9bypEtz757kCDRpTtaSW
vR5Sl6SKqLphpq3R/HcnJphqzbJoCunJjCGph8fRHl+RPsAOVEYlXRNUZSq5H+9H
MziyDhZe24o6i0hU2lJGw2Opi3aXFDYWoNllTD+tzQf8NxWKKy9+myd49cLLc64x
TBifdDlZ4qh0Lw6fOkeiqP9wl8TaOi+Z2sCB83HaiL4pnX1eRssxoLxHLzqsPMYI
xXQKvxQL1k9PpHZk7NksDrPwScV1qGG0t7IE1guP0IIJlB3prU1mFCer19APripZ
J9oD2rGUiKzYt7ESYncqLbybauDkuPPjd+cYdA0FELUSQb2FmigIJjtAxfXq9vg2
5xUIojaLVxAbKTeCDjPpSzcZly8/mMpGLttfyRdl/MJc6cT+IChe+RuM5u9Hh59t
vvzuD430tlHbqxVtNdHUYiRBzOfmzD6u7u9U/fDjwIc2gQqu0po15SrBC5I4zE3D
jjoq3oIHNdxcN87hPGY89e46fa7pFqL0sy0cXKvvBuX/R3VPuIz6UwBVycUThQCA
1w01WjZc/cfgbtfWxsYeYElvtbtqUG6sfnMwuwspZWZkgQLB/yew1wi0SFVr40Uh
WS2T+drEiDp1AujbkoyLsD4vseXobkmmh5OT7IdEohM=
`protect END_PROTECTED
