`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z66nuy2GtIeQQeblcjpAJZuFol6JRJO/4CQS/b954XyMUxLTk0UwfVU0+6kSUkyh
NlYlkOtJSlUCT1gwevETgm9AdAGfoxuJIM1SY2kEK9K1tL+YkK/fzMvKwmh5l21w
JdRt1Sh44pGDRmCUJGSEPksqUHH0OAJuYClNbO4nZjT+8GIsN0MDhkE1o+4jbyYX
opSMr0UpDWOdEsN5BUN8GqLvUFAGJsdkU7KO3+WjoU6tmwHr7LDZ1LFGVgudrBQy
rvylkI+Lb/sD4Dj7n3CSqXxKdauhvwOIGItAgfdFi+TyC1ptoa9J03LeJzLVd44N
aQW6jjBQGjznlH5efc5hawPcA/HX6v/re76zV3k5z3OddrkiFzqbaoCl2NnxV1Vh
qJMjWvT8F2kNw2Jjs6dEqvNll7JqwHwXPpRR8823Prw=
`protect END_PROTECTED
