`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MOXqzsZkx64QJs7nM/d9qVaRNWgfFznNXB6Zd3G9Ju3iHu1LHxZc1HcM4/9+ssT4
tQhQRM82zSYLiUH6RUDtSdvmQFoMWUbLNVTLfqToGoAZ6dlMjKazeXTvT15NLJ72
sbnj9b2GmQaztsfYFCG3HMC0zbZVwReLw2qkDUE9ARdyoMnEKodtapr8dx5gN0OK
XIQAZdq+XzaZPlMnD4EXxkDsmsN66cRd37AiyzVCcOk94/decpENvPjjUVmiOhN6
JKD7PsChAsxNE1+Pudf2x5pwmg5vgXD22LhIQINbADs7w/StDEcqZTV3nytEnhuU
BWVu6uz+5OlieKAIY+xEtW0MNwe5PkbdlwFsQNOL8vvZ2maxfh6VwnV6HBthUIEe
hIPoBxHwVXAR9YBzyE3+84sB6/A+vBDbVy6MMIfbUpR2nNQd9s+NEusJ4wWMc7sw
aXCrcQYolRCGRgZPq1E8WbahFdVNQLVYrQclyB+4zZ3jW3eRXwXf7gpJR6ZiVR51
qkF4yPMVyRKQAUBz0u/9oSQMKxNpKuup8D3A1z85fvD4YAp3bZwxHQqiwZGCSIyn
JZVNnoOh5714qN6gw2BMCAsGXzMYQ/96N4jkqpmM8BEQDgS5JHAaLMQukmcnEaIL
xwQU/HOB0DtIBm/sTvGYIMgILCHT92Xb9/2pvb6jHyWbrwCNKAsSUjjKUURL5PRM
qBlJY7Y+9htd8cirkISPkadqjKM2WqJ5MNIpKNNyNl622ZZafORYkbju+kCF6tVZ
vggJLWsOzVbtmXKN0kYtH9zEjkNawG+xhSWu45ga9BcFxaOSWAUqIpS41JrajRTl
wHw4Mq5M1z5M8QKl1EUaCsyS+ezHY7oRN4AtSpldn3k+G4pDg3e6P6n61T027zmV
CGo6U6dUQ6nSIvvT1Qh0ksox/O94DofykZio7OcOKzT8xgV52pDLoKFGpKGzhhSZ
`protect END_PROTECTED
