`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GFImqqhtdqlUt8MRrbg/BTo5KpWpJ0V5X+2QK256vk2AnCOGiUOLRzTObE7dFpJE
/RmytyWGl2f81V0t+4R3lmRAIC235z9JZCi6Da/MWFUIgX8fEPppNSNZmDHT+S3k
SE02uSmbU9AZY3e+muxfDgbMeH0CaKOPel4BxYjr1SjE7hYfjrXjlWJIjkeBgSjF
hXMjS5RdWKXJiCLMgQp/9fmfITtcZOKpkESDAQDewxZYJdIqKwlkyw05bzHXFhM3
i/X+jQxxQZStpWGzg+IKdQVdcuZR8dOJqHAw49tEBTaswGSGqk2jduothmaRb2bH
0mIQl9kRvblSLy7xXvStpDBesYwiaZbc2KonkscU8fVVumOnokQtqj1UuxVhRmLH
A9BNmHG9Ru+q3QHow85iVeuNg/Z2LQIi9NahAVNC+Csm1zoa6zeClSVX3MA1fWYv
Jp1lZ1oSZHYgmNqr9hCH80WjbXoukxgzuccQShtd1PywUiTZ5jzzqbUpbonpByXV
7/psSr2NJENZGJ7EAQEsTfufhHSpfy4xJB3YFRvvXmgfvZP/SvDnxCRT01T1Tqqa
2aNXE0Y99qLs6Y/zyIm29023+XMrP0Ud+rPpO6b6LODbPeWUl09TsEnwiwIz6+VZ
60k8oFsOcC05ebpwJ+VWr4/3TA4Z1XUHT6DbXmhAlL28omJXaJFxSzmF/kDX3bCq
kL4MBuj4dQefxCE6a6WnXkwfqCH5p3Y++aUkWOHUXv5v7eqMWfMKreTTfn4Fg4Zg
yvtycQE0pesgYNndIesJsguxZIUIaVAjrUk7iU2iGDGhuUTa4gFkGaal7DOYgnoC
o/2ZnWYJlgctaAl5Zyx9hUF0vPe9KLkOw2QnoAPDyvgvm6jQPxyhg6B9UuOLCJTU
4P599a9DzWcpdLaRZKbIBp+BUzgdSNOnBV9/jOs7KjiNPorPr6Frnswzzrqc5V5j
QXODWFJXsMxGhX9oHCXzHc8PLV/YwdFBwpkvHAgDkSgax61MTnj0L4ar9q+oDiHs
doDlT7htgT5y6mF44gcJvwj3icFXPuQGbYyccaIqkWlehE9hZUhe5JM+Z9wNu9d3
8MMwHKY2LVoJ2yzTQ4qFaGkgQmXJW0dAs6UZ/R8rDMDGudes68Y0bdmk9ViO3v+Z
DABasnyQahUI61CuYWXCxYlvMg5DrUo36Rz09qyUVGTSohsYXFKSH4hugQoBa8oy
/n7zGkP27yMOMoNyHol9ZcX18eAYFq6F44XJCc8lZwM=
`protect END_PROTECTED
