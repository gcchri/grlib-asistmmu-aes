`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YihHSxdAP4mUaDvAFo9aoPLIyGADZPuHjH5HsH/GGSnhetN18uG1SbPB4pWC41vS
3GQkVJyIVkK//N9Xt58t9IZ8LpKmM2lJt1EPGA5JP13AVG88Ed/yDPwtSXKUQuKo
oc7nhz5WdCovARXNNVD5dtM++kpg+Rwg+Gy/rjSwkEeR1SyAURaPp7ET0EZcZyli
AJPI5l+ry8moBgvEGcuJnWkuCfpWnZrZYgmMcEfZlLvQsluWylJXp8fe48omHlxc
OG0jDzvf9DcKc0ZugTeIyQ==
`protect END_PROTECTED
