`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KX02dbGySSzb0fRAKbdEDuayHLE2rgHdUhFaLJ+16snu1CxUla5abcHRrd4CDjBB
QL85zaN4zMmcSImtVfpc3gPZx7cdHoIWO63gnPJq50yiIKHw00MPZoGFU8Dmi9xu
q6Kx0/33jOv7Ts9n+MIZgRDfoJFJt30JPKJsVEynwomik8JqA0t+4ZpHUxdv21M/
oT9GVJqPb3vteUdOfvvRdJtlfTpgiFKrmYAIiZrqVetub3d9GUBuZqAvIN17DXmj
3bS8BsA2YDM7xM7wUfq4/sJxQDLDLe9ibwAsU+O7TErf+O2CoPy/UC9EJEAyrBTs
4U1mQben14lSPr5/FES2aEHbW/EsBsDdM8BjO5zbNx0TePiBwghggv84lDZcMJuP
sZa4K9Y4fC7z2FcZE06nujJaMY4r5gTGP/OIa6fKS/BjYHXiBXHvWort/XFP0NER
cXUqvx+cdFH6AheA/a6BFV1qbYPFAEenbMWS40+vPuPj7hejy2wORKvgsGISgNwH
/L+HAxlZzsbkQrfggHmvfqW2GhOZMC6sfNI5eNgsPvpKQWkOOU82FqOtWQizFsUq
TbefjmJ1lM/FPd2u+Cv7RnsiSxRpUm+/Lw+bleZToOs=
`protect END_PROTECTED
