`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mYrsxikSfLOMvk+tHzErcUWZtNtCKwX4/x9nKY7Jt92KvUVsHeuUCifbXxL1kF2q
Rxqe8uAAx4fvqI4z03ZcQetWGr24C+K6IBWkKjFzQ3WSwp7vyD4TVa+GEx7KQ3un
dcZPcaDbQEB0qAmX6FayHGuecRW29PR/US2p+zZ23SQWKyGXtTgH0mpJSUi3UZF4
VF7OqMQ+MeqH24oxcWi73leqOB2Pgo5PhCRwHBAQFKZSS57+MkqWo4mBq693aFUD
VG2JlgxISV++45ZCKbTlD9ZFhNZxMd/SE1FOUQfOi1I3giX1Nq0Tn8+9NFFUnbG0
GwupCuoBgrFdUjoKmaFBTD5/mAApl8a74Lzp/tTp13VUgvni3Uehwh4GPGw9g+rH
TLjwuXV+EQypJA75FIMPTIozIixX3p+pRpkDfiblksF6fiJkobBCQdPYeC0DRuRB
QAqoChAlL84yh0KDe69Zh6UMXLtM1ERjMJhBxZ9fQdq6Cuk15cdurXw6uaR8QOzg
vHbe5BdSGfRT8nzriKqIIPintO34bjnqaoUlTsanhhw88vMVN+Vu1ksOKSXX9Bxz
QYgft7CAtvCo/NIhFIlajXhewN+AJaS3JMJoJXjNgZK7j01w/OGuv0KSQoA5Br07
t+FvsZ/B/ND0cie7veLxMkwYggyHCFteFDoTQj50AJDHC8O/sjEKZH0jstCidPJB
CNbeUHNSpiCDRpb46ss8KPbxBflyDsrjLtfPUEn8vjrJwgS0ys/pADsS4+Iykuy7
TXzYmaAAWAaAXUUiKe9qIGlFoVAeU2M4wR0WFIDWNHMWdLkJY2bjzOYzmskOdTcl
l86pE3KcRhO0Mku2rKPem2FwMOI3sBfGnkiHM5WtaWjOh4n2K2UB0fLSVITSscTO
yro3C2h9mqiQTHlodw6+Dsx68y5If+1dh7uIHueQKiNaMSK/vHH8T23DEE207a/e
47bXqSKAeH/5KudfAnTSvY1FZq2ayhJhp7Y30rAuF58gm2KM8uoK4NkbFy7K0RZJ
J7GOT18FS2Qx22u5spTDq9QVGcgT/gOSZA7STqhNpPzHEVzULQuaQ/aDTnHpV5+r
JhAh8up+kQEWLUme135BCKS0JS6LwEDP8BnZ+LmHdr76kxEC0vw4+kMSdC1ld6ZO
x3tXVkJiX50lvIzibMv5g44PLZ7M1AEF98fgLj2SXZsZhcUEw4a+ZmT8dNeRBz1Y
HGSmw/h7XeSbuHfIaJl6R8cersMdjwOELtkae5+8vJTZTAMmMOcM4SZeai504U0k
4TPFmqqUhpK3cqwR6jFJsJpqEm23ZfWBmdt9IJ/IzIcSw2kaUF3I0wndRMjU5u8G
ivEnWdOpyEg6ufAC0y1zNz3+tNWh1PPx9pGFOhEqy+yPaI6Fnc3GyxzJ82WjbLH1
u26kqGqFIPuUEu/FQLFSKUth4EhdHUEWPaH+ym1t2JI4TA5RFps4h4rUlRwLdDxr
HtEKzoP+OU7Dfu81IUnbPZGcCB5vVABi17tFPBlnGJtcZBHhCj6Wc6xWdRlJo18Q
8TAxrkYFkkAez3J3IDN+YwgwQXmoxQbMc8tb75gdYNl2B4ZSy8qvJ4Akn/pc9rhb
tDyVPlbDyEqVKm7ro3Lk+4fkmvUlVGfEyBgYEbtpeSgzw5bIt96eNAV50EQwKnxA
FN8m01e1F2xf5QxOomrxKOWUIyg3UtRZk/0qwyWaXOjPsarNiHHnA4V/nDwofSXO
dwNY0l9pEYehke7mxhmSj0i9EgGy9uTnfXksYKNSIA1Ak8jGIhjl95ElrK7gS7mC
NU+j6z7qpAWUyK7NJQxhRi5zx61kjrPXrst9KxEPetfhMgYfSLvGAQCnyb2h5+/8
Cx9Ec3d+cjfyyKFsvHGg0A4UbTlxK1qbWrTQDoImVkq1Epc5SjLTiuiimi3bYN3C
v+ARqFXAJICoQgpF2AAs1W2Da4yMOELiNI/7g+iNpw5u6V0FKlI/gTQTxrtkDsCB
jClhPUH9iH/I+VGHyKP+2EC+cmBas861XG3hVWrg7jirEBOEK5WA8mqr2FhpvQnK
X1usZW69O6N9B/Xp49UwjbRjqAykVtKvevKZXAfKT2z/ZmOyXzW2GLGQW9jeJ44Y
2egA97/ICs5hAUB6WwIvr7mvJK13cuKEcgdZLCtmIsq7qlP687P7AAagM9J+LbfR
+1C4NjBU/VndpSHsYPWJSaMPVs1XnFP6MRGVxAAjQsDY9tRrEGbZt6SForh+Uwdt
0rpCHHih1HSCrzehn/5W48FTs+jtq+C6WmoW4rfvZuV0JaaEN4GFZlxW1jmC097I
FSErYRPmoceD2LMpXBJoKL1uL9MFoglABiaa83LdUdLmBow3oaemdf7G8J9yjb2A
i/RkogjCdZgEVEPL4pic+ygZzhCtarDSuAw01JZi5qGrO/afEL9Fvoc+X71rhFrt
wVEfxVajVxpPwebCHiVUsWjAbaG3VcgMKFpcO8D8hUJdGNBWE+sXFFbrz+6UE5pM
oo/kkMuiWuq3A0wwLa68uuLvo8PB+0nkgq35cUZejRmC/3xkqQWNsZ1DM3jpAHB+
TZklo3p/I6HjW4dcXp5uo5+xLPrWy72YBXgI3G57suYtalKKXc78M9gv9ch0JSFu
uPyc+d7l/KwJ/ScKUSzdziZ0Ikea82jkERL4DfQQHtegIvjAgw7fvz7onKCqoyP5
RiYYNmX3qAdqs8YsEsR8MmW6o88shQctZe1yJmrgb/f30MC4pL0+JbirO67OOw0B
PZy6cmcJnODMxVFLYAzXnccWPTgM6FfReUMYRzuFAPZw8cN6Z1o3vzyTJID5xSh5
pzhaalN3b5f745Ix9V5kEmJ+jg+ixUFvyfhKHJDKqcbnNjP/WL2hyAcbnsKi0fqH
fPoA7PExYpsLTBvfVxIFs9rUfUPlN0t9DUTlISlncYrE9a7EsYQ0+yBUPmAhyQdx
SnxtE3wazmLqRSS59JNs7G7bju4tXFHJl10wE8lyJ3gUcb1wNNCTsnsxJ3wCsNUp
B418JoNryL8IuQQ0B9KsjOZU0J400PzyT9tHyxvVPd3asn8IqlB2YKBlevgyEzim
itL6ESpKEgknvkpQgg53i7Al+oJtBypCI19+Q5CvCNgIZjEypKH0gaSGRrueUdCc
uzEIOiaHOFA4KE3Z/rRHLBnhmOqwWKUevn9H6o1tPMEZnR3QRNzQ81PBh7LrVWeV
FBod4WSRRjvHRJbYFul/LTZvNAzXAFKKNY+3W5ml/zK6r+eb5uiE2hmIEXS18TnF
mfBxvKKtl6gCKOysrpvTLLGrR5eeN3n7LhsibzJFWUvQOVJySiToY/oFvNjxYuAT
pa26+mqfPiSkh9rsmteYXtwUkrUWnYHv2hyVvCyJO+f1Zf3ebPhPdmQPbfrGAMhx
ATHwg0GUCZaLRTvbyXRHv44Bn5OaXZWCEoV5qMi6puhOKe3fCoB9JIMroeQBdxrw
xlIMacZqljBcdiwvobs7rS8JOE23BXZ3S3Ev7qMyIhAAJgcccB+XzDtz0jv2B0tK
2CyOEVbe3FtwCYDVwKgubbeeghp0twt+t63bpA0pxYGDpoZG4iqJW5DVC7/BK5a9
QbkGIMlwprWY+vXSytFcE2HrdLipAGwMHBCon6ShuZre8HI065G6EjVLGJ2tiGa8
m7Ms9p2nHLx5aljs2ffu6PW/mf7valzM3iZAtxcRm8Q7lXcIqEXTEfxzYdqhYnNA
HgCFNjc8T+PqATBhK9PnyN53t9WTt5tqvK9+t+3qgARCnT8PRrhyvtq7tZ9cT2YP
hEXlMMAPGsBc01qBUHzzYZA2mhqZ6O8I3UleVK8RqlMgwR712Yal5iouFVvOgQeS
lvh+DnrRZodYBx5BfE/linykGLTfC9mnU3gWRH8+iY8hH3SwTxxCKBPYgYyKIqSA
oexwGwvdfNojHZB/jaPxUaYrrDqVb6oagU2GFDTpz8siJozdYdBSg2nJRjhpYHv8
a75gZAx1TCiYbgJxhgyvN3ZW1fucjwiiXvVVI5WeP0RvEKeJdGVWP0hlVQa4FKYi
duQPnBSf9IhYqxSBm7LWpNOru2sMunbzmyubeSztKGY1QR1Kiu/KBZ5E4OmAU9vJ
tTCqAqauhbmrsimdl0lMS/W51q5RzoNKLK200eq0Yh1mWlLjYzTZ/IK8wdr0qTOR
6Fbf8atndhDtr6c4eXTcZS0NxQreQhiKkSkv0fCLFHAkJ+tu13o52gTuBEZDi46z
5fFU/Y1bvXoC9yAhFJFIoJ3UwaU+wWImh7OYqcsXPVCPVLsDybwkEb2HIROP6DvJ
Dh0izJL5ZDp6/gXJfAbjXz1AzJlWurdi7GSsZ2bkJyWwBSpojYImiz/FiAPhb8xU
k1me2Q0GGViOj0WoFQLNMOad4Pd4ZpO/QpompP8XoG1h2USR6e0xVkdcLYhRcLff
6wVMkhiEmDyf6mGXOYNFDrKyJMYbBqguwVm4VYRcrt2SHvMol2aZACkl7ixwwf3B
ZafePx2l47vedSWcC0Z34U6beQ77Tg2a6HgcQ1Y/pbd2uM9EFHmx+BpHghc8zS0+
i3IxuSV3N/0bdzrIdyPWi7sDc4ac/6SEfF+Eid2SAVAOd3e6N0xM+fABPa6SGESH
xl3AvABKsD5p3jHSoAzcA6PmPNxwSJSga8P85dlwCWPAoC1Hxv7mAw5XWUCuagsM
K29cww5b1q9V2Ker6SXopk32bBwAf/fkqq8P+UYuTOUpW4ThQ/WE2V/k1JVRUz//
MdRFwKi5aNk6eKYPY18T0WaEWCa40bAvieuw/jaqa2wkwJDa+O5N90bgXkY8ztlQ
PO8hAarzF9XJgl1f3GGUsr5Ico8Wtdsk/Z6Nge0aC5IPEWLjeq5vwSviJh/VqQ9E
1o3YYeAe+tkXtaCDHKu8V8r8VUXvzTa4K+iZIrdQvifHgQuDp10NCrR7yE2x+VJL
r198kRbi7ajvNA343bdQUwY/xQxVh0TCpSwzbZVt38zBlpD/aO1sBDc5lMHP/w+0
akrQtCobOAndlVUq2DM3O6QkH7NRcbnU1p6TUevh3b1w5f+P5WGYcseJHualRcD1
wb5OP5fhVnejkdxm/L7ztUdnKtxCL4kEJ78awQbL7SS82Z6ZSx1yVhkqUzOOXa31
LeWqo7K0lWboZxAg8CiFhSzG8tBvItgIK4XizRY+MN8ahvQlnTbCu/ItkLgbH6hi
mx6wP6ok53O4qxEfL9aMS99AWGyYX9r5X68wcITk5zLwHlOCFKS+d8rJW9gqg5fo
qvRxQ4+dKCviOvM4BkQFGn+DqgT9k9Dxf8/1kbMapORg0syq4sZisMx28y598wTS
a+OikJaEU90R94q2s52aJiP2BwD2+vCRmm0/0Z7SqzPfFmT2b9x4a4/FQrgbZNno
u/RGNRfxS9ksn75MtyshWvePGIPLZtZXa6t6RZUFph5qpflsLyvKcUm+WfAOWgYB
9Ghk89ROiAPraTJ52QZvC89RA12X2gNAvmMQb/X4sgKxhieoWZiXkm3S2MaWCzw+
hSO545Aiiv4j05sMn0zMcMeYEw0h68o4Ik7xYyLJVrBGZnjuSQM2v+4OG1BSNo4L
H0o4zRZRJ2O5izwOvHoItq8+1kPcdJhcKWXyGCP4EYPsyfe+hXEn9W+zIl2w9lyw
uyrOatgUnIUKBaRyYigejfr9UzJViALS8MzkdLRLftktaVPSCUEj3ml5Ihg5j45Z
0vPkqc5zp9L4AiwoJO1fLzsfRTHIcc53B6Og0wQ4SuFAztrxyU3O0GLnRgHiBnQo
+H9K6vjqzk3ZIsJf7QKi6XOMaGe9Es1Tf/S6A+iQKNpDGdplMmK3U1+4l7yeTlTn
ge++Ku6/tBk6cA9OV2clO+1Y8oPWztNXnTh3saWGl0uH1rhmNZxv70bZ0fuTnvOB
3+Jw2XoQ7/xW+ffTkUTh4rxhzA9Tngsx9YH0iApPXCM6qDGrThU5B52vjXW2EezJ
XtRFfLMWjYasfflvlzRc+fZCKLi8YavKgj2kReoCWEbAkdmQCv+lxRUcbBB1uTyi
u+J94Uy1xToOJ8yOMweuZLR8bKp4B+9ECdz7r2Wcr9i4KAPGoNq8RUBBLpA2Driz
AF940MNOnyyrj2GpzpVsp9T1rP5rpO1jimKQTBv+cpiXZFiDp3YqIkpf/1gkUQw8
sU9pe6Ab6SVG/roxK4OwFD+ANmH2QXRjWOpr4v3zuLrLHPiT5QfeCegCT+V3/GQT
EKWMaH8fcgLBVeGG+9BsBWEGi2yZf+hpo7X2dxp7cqQAbY/2p/n8RWB33eQ7ExbO
Pi4GQoEGAU+SNKEJ+QneX3mvPAPSIL6yGB0s6fXdrGU5+GPpYiUlNgqVa4wCvh8p
Hu9cwkq9Ep2WRu+X9uhHZh/IDdxxVT4Tzwg0jFLU/R6gyW6CiiPmDE4cB6qL2AaW
MXsmkfVXl4XFB36+RY1UZ3b+FBbd8sko3RRkHO8ejTgUuLlFVv0Tq6Me7ckhQtp/
eEQoxFxJN330IHTQcZgF9AH7h9DN0Bi7NNPvXb+Yf13gWgQcdypockHn/8VEHdss
wcrPZ4cE6Gfa25ayy0YBP53bpnGkc3XRJ36wqxzWdDWl+MaF0l94bdfnul0rVeRm
bk+xeC5yC8jjp2X4oyMRaWkMX74JWtG8xEqND5IYN67truSqfDWAPvg1dhsj03ki
Wwoej29Uos8YSeSTGjM7UTVVAQCxPPk31d1un5UKvbminqgnSreJPkapoTwmlbnn
zWB8qsAs2KQIQW/y+G9ZsIGnKJlfZ6HlBRu0W62sVYyx12FLTtk4qrDJeS1GhMaP
9pNd7iYnFNLk0Gio4u7ApHoPjjXk0GJZQV2fpyQyz7xZxtiwDRqHecrmqmOtwtid
Ko4gBayxDuKIFBYnHo4rOHbhfBsrcxhDNNrs8ROClfrewULSWWp2rzgLyDWrNavP
M3uKgOE6XDNPjxF5FkcSQhdleUONrwz4LH982JfzHmmYvBtN4R7sbJb5jWZ1HpAx
ZP+WUX7cVTeZVSkien2cwXN8W/rOSaj/MIkU1Bfbzzgm933JjglJBV8BYG6ZXIse
rhfFrb0nfDh1wW0JggEvH0fGmcISBmwy0nZILadixO27sBXmMphs6CApmBGj59+2
x1iGt+qFUG7l6Zjfv9X3XgMljocOOjj9E9mHFtqY9v3d1zsHLqTlrrvJ5vVLPzvZ
w+e3VGM8/yDHMrfaNL7/hWvCk+B6/vC22UiZVsQ8tIYlKE4qjRWwnfe97gQaFYbm
ljT/FNzjKd7cJUYyWBXve82+vic8aGOng1/jS/qehmmDYZ2HMNsNYt7MTbl6EBXA
GW1f2QGmZyklsjPQ4YAWwlPPe9vWnDMm70qT3L8neJfWPhQuKrULfDQ0snsVqQYW
OrUS2cZvVzeA8ridm/M5u/mP7Y/9UTWZQ8O66SSUa/pAxRMoTZfCHKzU7m+s20Rm
glfPfrpUKfWyMPVCBOHAtCrqHhEYCH5CqRrhsGoPQNuF/HWkwVtvJo5oh3WMfduj
EavzDjx6KSAuB9D46H5lAScrcAiRp0tse5izz0o+YOpe//5USKx8kMLqj/b2Mp9U
dP2q5SPdMxHI+b30zvKeFy6W8urG2y5fZ4rBHpR4PF0Zb8fW39/l89LzQzTpsRxg
ahRzopvz1062zRMve3Yv30lTIgG+mSwOr8Ua+MVIOW0faeyPDxufkSSDNi09JNv8
nqF0JXeUAy4UYaLv15AwEGuqnZck9n/Q+BQyYos3Mmab/82p4XAq52rTImA3n2Py
6BaxVpfZSmZD2iqNjJR/qgT/qZ5Kcmv9sPq/WoX6jaBXKWNGUeevbvSIO5ROrSev
9MDEcDoFzEbSQpSGgANCFTuQMi2sDHkIDmEID8nekgoZO785woz6CS+PlNcpQPzy
xGGBY7/Bic8JSoO+7IoTl+VXsMCE1bbHPrWLrNCp3xLUV89p01IPa3wRyMRKi1wV
F7CbV0dzulVkTxQBdvcWuU7gIa8GxMP5U2eFyLc+0RbruLHFZDrpIjvDymDCQmiK
E4IowpiLXtrUU91Xaxs+eijYABl3Q7QayvO8U8mdn4rWA49WP0rF+SrB6Wk3H/W/
aiPkjFqVeZ/CBJ1o/pSSXyVpYDzgSZsQ7JD4eNxKdYVPAQdkx1x6Bt0WMVBv4DuF
5yisqTPIq1CD1En0WGMJGTT4TrNgMSsFYUxNgUyeJUE2VaRTbPvprT3lsXkGqFdi
7X+6gogwZ2NatFp5yms7pvxesa/HorDIGISAWHptA7S6YcddzslEfNZH/bZnouTO
CaC0i5BBZTOjtiDlO4m4vf1jQzTjZDVwBct2pxSYs7dqLgzvFqmdp9gTAxLBC0QW
z5kA+5gXU/8Dfgh9s5ga+VNkdymjCVHaKFFZqcopG+VYJISMp9EA+3KB4D9avO2Z
jl1BuXuTfOoVwcqOw40ANka/Cuzy/7h4lzRiqcBx+IEdAdXpZqSyQ6wiV6Bs4h4l
HMnrHKg8fj1EFZTrpxOrYKkm32+t21eMGOL5iD+5JOpr+xACSNTSsshayTk6W/vl
bXcaVKI/ll9sUwb9CPLMJdJPaYqvrVomkfgPcHkQ+ybvEz81jSL2lL+W7j7IsYSd
bACEdKY3VdrOl88KF7TsBPgvLkBXy3V5mSM4+H5eEuBkSkeSjgCnkQNyBiSQx97t
zxuMEULpLd0yuGr21Kp2Dl+16VmrxSHOtbVNHOgTUeSzKVncnNbHPR14OM4LRah7
JMtJBa9fQDaxtl/DNdmi2o2yg+BA1q7+Uyz4xPJiCR29Gz65VoFAQwVPU1RVrPt4
t8LX361mlf0+yGBZQ4HBS9GbhORuQUgy/nCq5RsqdscKyGQSHsyyuHAK3ISfJrxb
9W5hgkSunIUtp8+zX6LDkUFAKWKO7Wkrh0Pco4YrAB8RD4SWuwJgUfLpS4Olmi4p
Bu1o9Tx/0JpS8uFaL8pP/CqpG6SYh2tYQIEobxulKF4r+yxuVT4cjuEy/A31PhSU
abexcfAbKQAKAGNBlJl5/YRFEP94UnESS0w37XsNWQHBiWYaLtMRUw1dvreELi5d
wKAj4K4PTiMRLUAm+nhkU3BCWjpRH02j3rSzclEJD+BnKUCNCZj7mUS8H49qFoMi
jPghVED7Sm9nw116NKITpexqPaT/oDcLU2CV0Sh9rfdZIVus94x0RiAmBGP0HT/m
odCun9NjHfMgk11rbSQPYVmcEla+PPRXEjEfkckNCg74zDHerwe51f5+sgZaMkNa
FZcX7U07mkYRY73+GhHQBt8sIVAmA0T5X61oVBqp+OvAaDtEY5FHRhaU5zDfg8Ph
P45p9FGwLfjPgf/CcU94rt//ePgHuO1ldBlcYCeSmm7wg/f+6U1SGZ/u4BsrthSF
FgsgcHoLYqi+4SD5oIKpF+UYPMXb+G49VbrPtGJNBV6tNgiwiRYTrfXXLtMSKNZN
Iu79bi105kNCs+zYNWmUU1o3Dt9jJFB9f8FdYbCOFCLQCqL8zhi+TPkaEUpsXTD7
hB/MoFn454r/rtBUD4+5+txVbGQcFo5OwbllGgzCwvXB9l94uqvqwVz/GzHCWBDN
LiXtNR91sYO3SSUhGGePJRBhE+g89rakTU69KwUNj6ro37JxzXax3ozPxUt6uRz9
NP9+vxEN1kci2Pj9CE/tQvt/k0KI5H1mpnIZOdSUgTN2NHoaITTnDE+d5FkGgzd2
KIQ/mTbSSip1eJciRgKXL3zB1Ch6WK/FwMybsg88u/EHvFX68mR4sjBXHCRiXm6G
KlGqHgaw1Wifiv2CERj2Nmy94cKUptD+cJoSijyvwUbkQOfwYe4lP8AKIhBpsa4L
MkQVRCP8MzT3V3/YKtnDW1rbuCf+Ha4nJb04hrLLvdQGU8LzfSbutYTtzaI2DFrg
02fu/MECkakDTZHlJPMlJ3Apypv4qQCcbns6miS0hI3al8dgEO2I3QRgwqnFYCQU
kkoUM89Y6Mhkl+wGfSb6fBDUm0qS9k5x6lcfGMO0gRm97agyGvOPAa8OgNKL9/aX
agQfS0xAP0BmGvuy3dpEHqxsmGeuWTErss2kO8wluOM63dvHryCI+8IFYl0tGE7z
HshAq5s35GRN0XHV3WQd69Poo7He8klKquPlrb/HL4Zkqml3eskAvrShQvdkBXqx
zeL3f1F1UCqzPB3J8/xmB9Jdxl9KP1fzPoC1s++4hnuBJN/FPTciLTVIvMOwiw5H
QDJHgagDgRWveFo4Qwr2Z6mopgelt4/FTvlQRRGgNzPv8BUYjIxninkeJ7nz/y5H
gZhpy4oBOoGrkOXstFM8ieUvRZ6XxyUzyD7ulKb9I1rWyv3mTNZZLymo2NBbPzyw
SqnEa3mJZl0gCc0T5zsRrTAgZhDn7eheGvLzKk13W29/7OdIP5Oe2J4AwekC1NII
gB+9giXeRAyyrwKFZrNsP0u4r+k4fLY125hObWWdY3RUPd5QsoRWDkDnDW0jR9uJ
h+NkCWScWZAF7j7HYEK18x0R+Lpw7ScFV7GIgY6PljRchDDg3cCxr27MvFsHh4Cj
A30Ics8p0wGjDeWqXbF4hArM5cCW7iijcr2WwezTuMqNY8vzf7HXB86+kzbk7Yc+
wrCqCJC1VirIpjrk78sVVB4OzKoowxTa1e9PDIScWvKBRiDtQuVYJHUpxEwgCBkU
t8HRpVHmuvughYC6nJVxvQmD3BqyUUM5ZJ7y9hTzDD5kESgh2FvNfqcncHDV+3Uv
c+I2PLWV20JiZ6q57RHUqfKaMAizXTH5G2D+/UDh21mUqzkGmhZX8ukS9TJYXB07
f+SroBLpg4NobMh+GNzjCXNaly5+ZH3Ou3nCs/xozI+kldLT5pGAQBxnxWuz0Qj/
+gI/Qx3RfRcETK1nP0FDd/BdrNh9Mb7En3qCnL41VctgF1JqXMT7QZTXMVXHT1Zs
HpxhR/Sv62s/KvcGZHLa7vZAwymxQMNkRCMEIrYHGLg/uZEaXyYC/17IfurfmP44
1u+Ie5/WpdNOMBopJANS1WkuvSnh5iWLv3sxD8ovS5JG2cb+uk5lxCmMwWG/X+vB
/+JZfu5qz4StP3Z/o7D979pbls3VFWyUOY2tGPqYnxQ308ncya/ZMQSTVtkkkeE/
uKjkrIiq67Z2wkgB7fexrhLWYru6hzaMENN7qs/VPjrGquksbkDAUBF/AJFG7NRm
CLpWS1GyedFTRjM3ttYf57r13t3AyRTpkcxVUhp64LzfJUcMxr56IyCrjWPxVyCB
0swZ9gQM/jaHXPSWf5uSoDTKIidsaWOPUFLCg5xISOIVtPZ03Vm1fBaE/fSE/5wa
6lBekcrHehITe+3vtgaBrTn0SKM3v9b6RbO6Lk1DxheoSb77VlaA+0b4hz73V8HN
saqvo1M8GHcZ9alPrOXidvbc3sQkEz8qUqfyzjAGNXdE3LxFF+WPibFiJS5Mlo1x
LaPPYlO2P4iHa97KEdz5jW3NaRC1s3D/a4HVAZaeSAI4kdwuzbDlsw1Auh/GAXij
Nhm73SjJFphmLLVKne3S30bsX2mpEJl/MWoUySeMSaR+V6CCWBjQCHbzgxukq/a+
3/xkq3Rnfd9TYv8RGL9B5cAZ2dAEm4qEksNwzz3l6ApZ77hdr3URI3c1m8AlN6qG
xjEbCKy2N/WJ60hzQC62YOm8jtie2cyZO0mX8TnNe/ZZjdEaoLrHpUC7GJlPmus1
3j/cUWJ6FHwPe98qDyKatgXeYc6fNE9wDCVuHVCDoJEsOtKCqYc7yjULjgdyDZzO
e6COcptfgqr/wtTQiAkrnEl9hHAOHhc/niphw9zQ1g0ziNX91IGzKrdEf5YHlm9t
zLmW7MR98aXPQYdnP1lOnnxq26bwuR1y1xatKWWNN0lAzYT3BOMbnNMYsLjo3LDD
xaiRvRiE6Ol/2JBgXuKe9GNH6j7bTaYuhFn3vQ/ICe8IRjSdLclHm3hrMTqMy6NE
M2QNkyNy5Wi2bOQELwHLiMHOptdtvKHjLMVyPXj95Wo7Qf+FetYCwUcwTD0C4fsh
Y8ksQSKp8yJA9I4nXqPmwCvXgEcD3Qvrqkl5SkLhSHaqyJEDYPKyR2pPTgTLNzs5
fHIylKFn5S2O3sbnwRxSCXFcX+GGy6w8HR6pSmwaWh46Ej/NR/I28N9N34dOXAjs
rti1YUpeGYw+dh9Aa/V0HdOw8rIfy4YYObu84rdezX3kQYN0GEF470SsqLOMQO4s
1kVj1p93DvN6+JKePrP+Fx4boQRhdGC118CYp0IlTPEuiGKztui3h9w37+HYbyca
N3w6CBWI2d4Y3q1rMQHa1sYBybRUVrUJzdIJ5Dhon0ebc9qf4T7gjxzEmV+PDD9u
zI+0zeDvpTyryJM0ESJ3ucu8gFqSXzK4/LggRdfuUk37GZQa188Jwc4luKYDbzdK
i/723jkeAyy/KwEaUK3U1DaQnFPWPFJWG8Fubkhwx/lAN026UVzBy2/1NWi6qGZU
WQOs4B0EsuXlchfkZNWn/46zZZoJn1J8HVq3byyjOVGTx0qZvK4xoVFJHeJMMKyu
GMeba8Dq0otZhIGYktZKFgYwjGwMLkzRdB+x2muz/RcMYAYSJil1t2vb0NeCIQ56
8cmLUOOOQS7ZtRYOuPD/FDQ5q7QstZWmdDTVsxxJbtq4ijUJbAhfY7gw5LINK+QT
3M1CQxcz2po8qppx6nA4oszKpbeUxCcZFYbKiedjJTTAlCxCT5kJgOgAvJxaDABo
PXo2vj1QEC9oTDjFWQXKqk+iLxO/XKsnWOSj6FHiJ/RBwt0Sps8w6hua9KQfF/0C
3297hPC0O9MoIxoy1JwDObOZCS5hjFxcC6o+wSzi3ecYmaAT9G2u6E/M3y5su8Fr
Vzw7r//C/gjw5tQPLTB1NjJR0wOqq3SrbyEwp6uGdacADbXiWa6BWTtMmfLk4sVk
LDS0rn1FR5v9E8cSEwBYNFJM2J1XLnzGVHbAZBYB/4Lwnx6IJ35V12O2+ZHy9j/L
Hattd/bK2JYXYpuX+rCvBsqv+376lrclDV9dhlEZQctij7PNRGpCHKi939OEctbS
VuUUMoRC17NaTNY2i+5KEQV5wHAqdSRgE1m8PxAql1fcKXwe9zilI5KjXl6GtvYr
GxzYJRGBQP4rSP7ybSctVFAhY1swniRO9aOtlczP0KAfp27MAvo/4IP+c+7cGXoy
rLrp0+7uppVmqjz0KIXOW8ryZ+oLokAfVgF0j7KLRuhsblrYXQuAPy2qhcQWTkMk
qCLs3m+PM9lam1+qMQsKcEZB4SI1lZT7oV1wvi3WRjZ8aMqtvqonN6g1Wp3gpkiM
g209CCFCG19EjNIHv9UNwP7/ud10I51rl9xbqZCoMpiw/aOFICB2tD4P/jrZjpjP
SW1OUhJdPjwcvU4/zvKZtJtQoV3LKPnxLUS7fuBFiEHfsDjRTqRlVIR5P2JQxvdY
UEI8CWIDOm8BMRQO7wj4qRsAypxVT1ixoXA+lxrdpankyGP6Q5+uZFNqRRmdPtw2
J+Ykp2jSjlrlaY67uSIJex1qmZl8ZeDoZSdYR53XXfZfLrxIKkZtzh339uaeU9v1
FXxZM/2UwQy1nXNuwyELE0E4X+VFWTAVtoID/AJ8rRUc7bzjSX0Rqsjmk2IzdkeJ
a8OUqn6WnTmB0mKNYsrV0HEywSLQ47mNYUnDG5xtlt1FJquP79V7vbGCz0VN/aUb
drCcWQtBQYGzVlxnmTAk4h21cUEynQr9gF6KokbQsGfmpHux7lLxey2gUb7wJ8k3
VSmoS+5G/XzpXXJ/5k5PIicjVVyWIn3hVh3Iu3VM50ib5NVotX1zj/dJWmRofVGz
I7nCBBStx2fH9lCmxa+xRkSBfrUQg2T6XYKDyVFyIRX6bmdUnzHvFk9VD6pM5Nvw
eWzCkylt/NTguwLy2oPvX4Kd7bKPa1f+pK4yRFYCpINuYr5UUulnyDnyCsV/isF0
No6Hl9yx67EiMG4mvW4dy2f61AVbV71xguhoe5BZ/GCZw161QCw4XrhSQ3dEagN8
WAAKlfHXPTszVVHcPgFFWp+3d4twK1zS1dWjy+kkwJnFDdzUMZ25wpVn+WgDUIaM
4f6se803xAu8OQRyL57Rth7HrVQBtNOI1I15s/LZq0aofjRWM5S/qExKEjzjDFTU
yra3tb3CHECNWKtE+19NGuGPfkQvOrk4MXemb6P4fDuj6p81BjgrHycfxYXUEGOk
T8ndHgH2XZVQgkSbPbUuD2gtZOTwRW/H4IXMK+cmcVV9ZtdJMGGBOs1GRw0q9gVO
iZ5vp6bm/TnBb7MBDi9eY3JBuI9SIiMbAqbf3NGITPBeL4izDzclAdNAkpXBjyE1
WhDNFQpLb2fOMQMzhd94G6vAkODOQavs1d+KLw+bSgspxo4vXtvAwRui0ZaOc2mz
M9A9z5vvce2rx/9/K9wut0jj2UVieg45K9Ia7q+UqCe18SDDQSAhjCxKQL9ekNJ7
xdYq5F4nwSERGjrl4fO1n+wN+AK6cWhn96AS/0DDDCN8Y5RX9Vl7OhZlpuALXumQ
mSVoI9j3AiDuyQVLUhIJcZ5uR1edZwXTxMqh50Qy9llLZzmTOdJVXQWJR1i5Uvgb
MGiaAoroCS9a4aSrbgUrtIXhTbWVjLm9n3g/qC4NRPsTwoqsnpuvkb3tP3Kqu62K
4W/4/7EqbcQFYSFCB5gyPiPy5yHQ8Ser/hIxxcdalnYoHgt3DZBBsJ1daL2z2G0K
8VsEm5C9kp0D45mWA7l0qNAdv5rXJgksIYsVpyARWcooGU5N4VIJEbQwu+XEB0J/
uU9A3sV+oglEI+To9d2DUbHkS2FWiSDjiZRfxgF4w++z9lP3yvuIbxRRAigYUpLW
oa3yzQNP7cLNOmeZIMjV0e5ROimCNj2Yrr/kQB3tHSLZBTV+zlmMB84w28Dvz5tm
/p+s1LdZwqdvvQYYSSxJaKwzeJWvr23H2lS3hETiPM8govWh/C/JA2cb0ONhDgBV
zGCZhjjKnyzirrb7V56e96qdjNNh/rlBjHcRRhuNlaJOHmPyVrxR9qJFiwjQ5e6C
AvLUv40V310SoFDsocLLvJ3MR+WWkaJ5eFUNN6pFdByypF24Zw9vd9ubpMxH23Gy
5092iejpd8oF0ITrtFSs8+InW8+g/8vRfXE7s41dGiVRw/Xz0epjdiBD5VJFU5GU
eEvB8mOwdcMuYzREcTv9GvtP8QVTaFNGjMuoyT7/D30TPzSXrvLDW7yuB0JUsR7n
AXW9iDoVipsoBfpj5UsQ4u1uAlsy9j9izpPJA2wSlYEdQtmT+VOTmnJVAApqY0r0
0CMbndXnai6f/5dZDXZh3LRiKzeiyrDxEPz+qVlYl3amskIbYy61W9kg3BBY26BH
tc5wOpaeIfmYxQiUZFkRB7vn8FgWvocxHdDGg0FL2ia7OiHYbeaurr5qx5lk12NX
rhAYdrtWCVfxruQ+FzQMry0i/M6f87c69q/trkPqKyoUCaFKZJJu/zmcLYqqfhOn
/2TgDFHYnOGOu05D/lIgM8NdAKOXov/6Wv59jGjFC2/iPYTrOyMWxkN7iwQJ7iji
xphKUzuDutKlCyCzRvsnvGoH/0gYb/7Y7NChs4m8Mxio7TKc0fdz4t59iSMImJoN
7KYplqfzMf9D780+7p5B5FraBGdEojhMLbjCOdWQihZ/rChb7VSH9OOJopkgEgra
O6oT2R9vNDBosCkflsPd4dR0CeVLCfW3Rm1vJ8oOeTj9w2ipiZdORmbVSSZfLuSP
GM4zk3HDye+5vGo6sZWTTW+KngSgKBgVI7EH4E7nAQXga8ukUs3JFwlM1j/hvQK6
H0juZGIJCYrm5NR5eRKiWNskOZpTMcF3gkHLebPViG2P2qqOc9ARa6i3cV8KCcX5
BVlNTgQTs1/tSHhmvbXTCU7fnGEC6sJsSmG2hwirxp3wyKRsyEThFpXFUvcNva2y
CPWANl0akUuzXHMkXBN60wDgmiXYTvDac5mOputP5EKJw6jiBfINRMvXJs0j2vGT
jcz80J4TRKijnC0l62YLcUfbDFw1Z/igDWF4E7EIA6QiKLQ9aEBbSzvVg0OpkLNx
KJJfxFkjIt5QLNC9WsDyzM0GySDMxeBlF5qCde1b3x4DMOt1VWGSYLHvcjjVUhVO
6C2+dE91tRtcggAWetouJe6tgk8xQfh1PV4FMbGt28ldYyXNYIJdOyiFX/87gl8x
i0cYpRAY7cutO9Sun+8vJzhMFM2ZQ2i+0AgmnON/Hm7A04z8Voj8Ul+vHbi3CG3f
D2N1jH+sNgRdfww0177ATOSvnbTXWkzuOULfakPxWIj0n+ovXN6ZU2uKEIHr7HOO
p1lqCIL6Cf/tc5D40gT0ohEdnpNzsrQNF//fvbPwfnoKfJcGTqqMirMd1bGS5eEh
gixVNu5x72XULqjZVF2Sfs49ANWJMIx1Z+/bE3XreOjgr1V45O/hwSNfiXTdwcAL
4f7bQduhg5XzT5McgwBCXXh4A9wTxWEPUsblO+3a5FF3kx+3ujkOpOGQ6/8gcej2
Cc208xAlx5CONuoNUFpnZMFcWLovWCm3eekPuC/35E41qeMZ1x+QHwjvQ+dx9SAA
aCClA9EHYIXED9r6k63jropCrbf6xQlBoD9M+uD0syZDj1FNvkG8Pum6O9/9YHH3
/N1griCJAGOKQNe7q720E4ypCoHzBYw2UrBMhqC5H4tnVbcet6DR6qewLj6AKm0R
m54c+1FmK5+o9kaxzo0ets4bWZ9OL/a6Q0iabAKCNpus/i3VTtXjxBN3Zr5+DJMn
OAqhPH2DforYsAQa5LsY2+8lIALx10YnRoEz30SQyXTbvRs1F4LaQxgaow49SvER
S0KYbM1eYbdPtjlngCxRLhaShuFx9fqpS4m0I7uEbWNhHxd3XG7yIo1Zl5Yr4SjJ
ytXbzCeu78ZR1agqKPTGacp8sFHelj70KR+I/oCwEn0WH0iSW862vwWa3JQ2TVjy
kijFct4NhZX6K1BAY3rF6UUArdy6iHquvnD3PaozyuVZ1oOZNpF6WMfvV3YrXggR
qqAv8EnEV1zdBZ+g6utMUIXCmyJVR7VJTcuwX1ehy8xGxXsKBGUsfggxyObrYOKM
osCEA6cPuchU2RugZXNZLA+FMSyff2Grbjs94+/Q9LYIf8lt5lmDzi0bitMjQeGK
++EG3DdUNpxy/CENxAKpaJoo7+RgbUVzPLP3TkpXjw/CJ3sO+91fKePBdrhtY1yZ
aNayv24+Ra9eNGdYnRiXQ8dVjuMD7zMvUgJ17qgyLMm5mGWvBK1yOwbNf/svOe4x
WOQq4lccvhUOxUHOPgPAbCjV+n/WoRLoVrBRtKTidqVc9uYgJxJiTvEMknUHbbns
J/dN7oNdRtw5hFquS4lVIoVsFBsukeKH5LnEPAu+tUFzdGsiZAF2YoG1rrLdDG0J
AT+96XsX1LeW8t440sTOen8h1ZSJcnRrpYYGQMH0DR7Qquwc4Q4RLq/RIUexJRHj
AugyEH2LAnXSYA1d3p3g8dpUqGKPDO2/jt+k3OuDKeoj6gFu5IeLFy9guxzXClyH
dodk2uhdGDtbrUWp6dUrp77APIsMVTyb2kwFjdwvZO3cqpxsd3kwFKf1V92sG/EU
6U/Kx6ElyLBbf+47iiVdIYR2ZYMIRP0RgAoPGyKmmPYf3fPjq7WN0eRoL75GP81r
wRxP1u+6ShdcKNl3AymGyl15Xfvld64Da0tJzXV53IgXG3P9MOCZpfsYfcEqcamX
wxyY7aZJ3gQOLMOCQ1OASdBtwDG3CMCsZhv1D515frOpFSNwQuR5mnACPWZqxudU
m9labK33qRJA/Tx3BfBEfk02wzrnGRoWHkC2+Ij9zO8J7niYMv/NaTQVkCx4y8GF
S1eNaqdAsd0/nIQMv46Zs/pqE+lylzpsLiuXekyxHByyI/LaF0QvRe9dobCJ4W9y
W1l9O4pTZlJBlI1MqrdknWlCX+/PAg5kIZBKTqEYsxCwmRfEDM3B0sKPdqY3WG50
RaZ9HmDk+j+MCtsmdXB4aox8aIyzvmRHLeIVhNOxuV5SydSaLUKE0JttlHbGn9mI
q2SqDCGcIR8GaVvRNZO7KXwHx52M41GRJx3NLn/uzZ66e8pVKu9GYWDgaLdYM0PU
1kzVIahPaygxoob9iRGmgUCuievNrrXWEGGlS/7qyy8CEOL4/Mp1qy3PNyjcCbRF
k0d/umyEC+Sot/WOwEyD81FV96MHbmEyUbhfnhazowhsa/ss3DzrzQo69ljOM6sB
SGZy4RoWAvQ7y/PgCyErsDHQdN7KPTxRWjwA1uAXACqFREv8mqwonjf/S3Nxe4Mc
P1xzz3Ubh3GwZ40x2/nue5paMHV2Ca3wVkn0TK6bAphtuVj80bRRU2gxl9F6Yt59
ocNM7RMC7BY6NzdF+T+dIgXSgAwxfkz0+9ihx60x+uf9GDmTa0Sz76bG4CKzw3mn
6CWVu4oMlH5TOoDd0CR/hoc8ohQBZ1/y0l9daoAlFBuY8sZTKjib2RLYE/8AtiKT
Nche8NVG9oSIlhOH1AoCbERFfwEVTLf9GaulN9OnZHX3im3EiNIdYIQTgm6CAA2h
ZeWfXPdvm0MorTo52yTfsiApxLCx2p+92h7arM6WAV6nRcMMD/Cd3JNeurg690IR
KaOT/tAtyavfaO6a0v2NMvbv8cqL4t0ndhNSuYZYELCqIpLSmOCAYHmrycnOU04Y
K439AfMC6G35JtllLOwoBDV1WziaUQumqeCZ4AZ/HxjulrUBmfJKfCOZGoj6qf4M
j3WE48RdArXpaF6EvGF9BeUzvsUtcDLQoshHeF3rMLi3vxfHfN8qQvC0FoTou+23
skUqOZ6jBoNpIRft/u2JpCIw6RUAUYBBmHTq3u4I0Me3Nccnnae5VR+JPhGe+hWD
ttk/oOa7Gasjd/RMGTVW5+j1E16Ran0Pj6eZ1ZODY0fpB6mhhYEdtD3CkVcGQYoq
B/NKsQFy5+aUaXGlGLIqjtCUDG7Kg175UvR/7CVrQAvZxK6nLjgTIPFohJOEjCTE
XLM9G+0733aiSopKjpXlZOiivE4aeR7+Q+6nJ8TnnpuM+4ajbyulLJjNJwqug/tZ
G7RpMuKj0eWIiYBQgNDsx9iPY5JoAsG4IouvpOD9TreXK7VmbIJZ4Z6kyPm4x8pH
NKUDvQyQ+YZsFMFq3/lOA7J48iRdL7qFGrDxXkQ8w1xzj4x1rJVIZO0pCqlh/RVL
mYPyzlxC98nd/5n84idf42sISrEbiQn4N6e4RS4k11NgPA3Fm3z2yMLmWW6sSqy4
zSBWhBDapXKl7bkh3eWXQbmds7vT5/Ji5Ruy3y8ubk+lXsnSK6v/Vr8WyXND2vdr
bwbYXwl+nAqxaq/0FXHF8x5GoXyUu0b/QHhoUcHXpjtlbOe5q62FOH8TMWe4fJ58
UxopXSYsCRRMxic1mRG3j3/f3jBjLDAOUCQumWn+jbfJjwhxk3c3DRctBNwZWRCh
c1Er4Wt+6lFzcbISapZZW8SVcZLD0JrZQ9viH4HH0iOCuSaRlAycxWpYdAp9Y6Og
PIXsLMYkDyZMUhzMAE/LbCgFAkNNc7L08Is1UUrHgFxLoRaMcurx6P+47XiHMGLg
fzLH7KUZwDMkKIjblNZo2Mbn58flp4J0HvSXU7/B0LiD0F+Jx/9AmbDMlloJ62U/
pUGWv1Pqb9tlB7Vc6O+QdQbkuAX+gAuv42bmKVo7oSd4CThDysAS4kQHnA58taf0
Bq/12md3RnqUPokhM93/cgZQm6EW73i8KdFEm+/DcQOhaA1W0WkVJWUvcnnwNfbk
iWEusDS8yffShZCY4d0guH0igjfdnEbqhlrpMczsGX7xP9RENX+LGx2DaZc2qJhH
zU+xJ1Q6HX+mRo0wTIpUZ4s49iZEo2HqUxOvDoC/b8djhWv3x3PtMYdQJFfFLJU0
nqd/H6PrQ2cFKQGH8F5V8xOMYnXzDw5Ur8TKXrvU7JWi3bLsTFZqj6V/rncuXILb
pW6iocRUUXNOx6tLIvqHkSATx6+fs1Q+sHKxQJm7s0ekVx2ujKhp534rHwqabgGB
9CuetqLzt1s3ubRy3usHDfwm10Yh5lOxTMmJV502tGhWK1eV7Pa802lP3xTthaAS
IZTNykK5oK9t1MNvTNgM88OiiaQseqvZpx75bVT9YtxXKVerX4MevOudb3m2ueCm
h0W4GJLNjoqxeVITG2iiKotHZ5X8W1ZWGPF99Rh/Fr27Rvzk9MKBwo3MheVjWYHh
kDXTP/OgkD+N6Cv18PRJ1wDwSdOz0Do4lkVlYDhZNrcUkPMb7pWs4zXy9NnyC8A/
N9VChDIezVLgvoS9VGNpEx0p7AZsj1G5zookcGv0MEdq5jzfW/6MG2X9UW47C0Nn
NmAcPuNuXmH/JbffDGPwiB2oerDZJ7N66BJKiPp+DheTyNfny8OFRJYu0C2jtlPV
XkpUvjBxqHpWIu8q7AHU3Hdx0hd/fF4CwX932FHXpYyTZANziZcEjoEGuVpOzX+r
yTnctOFrQ0TCzXyee+VlbeU/kMZQUpt6E5Brun0sLOFxeCcahax9+MOiRBrTXHQK
78fXhBX/o5dtIaOvZgsmtNtmWNyhk0T7UJh1i+dQWQcJc13OVa1humupuzH3EUPy
AOLwUZV1TxLlsOX/+EJ5dmwu2X5ZwRZYeUPeHFoELZcHgPRl0MhcepnoHlrm6wMN
7YlY9jn0nOmD5Bhmcopk3KuyhGNpEbOT+yzeq/PbqZ6aUJsqahSUGr3NVUwocruN
eMJwhszfRsEJBLDVUEGNV2gytSLdVZBzcgEZzHGbF2foapsbDlVcKMX7+wpHTZoc
cbHvec8WN0C4etLsFvpKOTl0pBM1dxqkwTk2dCOVNM4HGYgVxb2PHbQAbtT9yj1n
BbwqnDKHFT3O3k5rJekG7l8UUnCC75iDBS2hBIJD05nMm7sFhsnY6lQ/4wQG2FD3
+W6EntYAe61624rmRUeEE3yYYtuWAOBiiD+1iB1jgcdaYU7UGUbCAMm68EEBP+h8
66bW7prPUR1FNSrAlp37Q65TjgkoiwGy3EqSHcV9RAeSMpRzr6lnf7HguLlBLLGE
t7SCc5ynyOj7QYS39mJURL7kGs+VyQkXmV/oB9nKdyBMU88OCt/qShW4M0JM6eeb
kQm5ODw6ZiVo35Z3y/FStlmh7tzTHNdiYUWJYwSDmPHd+j3iA3pPBWVKSxFzhqQ7
opJ3apT4Pv3RFMBRqMedOkxUKSD5IxkPL1D16WFIQs3+w+hvapIqlv0zmGeBistB
OmislnvVSCmKkb2oxRQmWpujCf56eHE3vAUWANzYhu5kjTHGxiTM5k9gRsZke2lw
EPD5m9oKjhbLvwTD8A/WDXSuVL8ZEjliixldV7vO656ZOgJ+hrMTvQFsi1GEdfRC
B5nnmELXm0Rz4YgRGCx9q8/4u9ZYQE9a3GIJ6AIIYdhkF6wIq8ty7YyqLi1a2W5E
//MKjv9+3VjIRzzczmPDfNcI5G4nMitT1OyPrpJfmDiCfWSfXD7hKIAARnDBRTSD
9i4XcMq6ua44Tf+GSb8kBOOG/qbz19DA/N2dks0hz181EHmKXxMtwqIqs8U+OFET
o5DV/9hLZKm5bigF6YL44nwH3rPAnz7MmBUXpJA0nvxvXqEedRDHLsbBnasboc6v
PV/lCjf/JHuDjI1B2tqI9CffebHnUNs97yz/w0R22X0=
`protect END_PROTECTED
