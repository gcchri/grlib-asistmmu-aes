`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0hnJseQ2Mh3cDqb77SHyDnOhHG3k0tMVqznn7sJrq2QV6i9vKT4/wVCRwe0Il0kX
fzpK8W0V4BM9rTqDPWWlGUVCJkpNR3bXYoj1RpZfH4u0ic24dz4YfuT0FZ1Tg9IY
Hs8xIcfEJ5o4Jlmgcrfmk6SDquayuOaoz2Nkv4CQnpyju2eY4hQYwDYc2PAn1f2L
1+mSzwcatfrUdadvMDm7Lk4KqLMgQNscH3IlJXen7dwELCJm4V+XYKjpYXC7p2DI
gfIAkQVQInLeaZXvcvz1E85NbRlH0pr0NGYPc7QrTTScA1qvOkewfAS0gnjjRBsb
`protect END_PROTECTED
