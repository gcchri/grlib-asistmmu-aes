`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kGP6t44XZ67/6i+HW71zS1DLcWhla7PkcJ1oOdKIfVzbRR6XFqgf/2J0bl/UA5r5
S1UDUCWdWDKjUf7UOnOq1YMErCMxU/tctni8fGetQKnhULxD6k+IjjzP9ikzEPOG
KDul3ZKW0v+betVg3+JnfXk83G9Nip1JyyQ7i5mAXWTZTevlzMvNNP+kumeqoNrK
ZP6g6lcMjcqBwCNDbW2bvMphrs6A4U+PiuCI0yj+eG7qW7VXuK9UpehGgep2GSEh
KaER551kKZcXnquMTLdlrzoR0HuO34Nvy/ivLhy2XNlHPLSyqYtQxsvWzb6duAHG
MvTyAn9XYs06MZYeTflCWNHXa+Ak5LUkUsfHVAN5fQ1ZXW/vnCZbXblyuqN7uuJa
YuayecMKag382klKqrIaEbfyyomfVKm7foHPVmQaD9G/Q2kz7KvsxmwhhdDBOVN9
`protect END_PROTECTED
