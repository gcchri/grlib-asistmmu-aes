`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hkcfNNRGxhfcNrZjAMZ/u1auWeCESZiaphZE6/wBODWNGs4/fCgSJt5dGgqEinZj
9suUY8u/EPEbHago/70Ognw8QEpQZXR2phP/1Q/AC+gmJKKH6rOT0VS1C9fFiak0
gIi26bjtSip3DlNktxXNJz/el5LMl0YE+EBP7sdwhWyqZatURjtlC+4n8sxEOMis
46PMF62fRoTyCq65GAJ4UMI3DBE6tVwbmJjJY1Xi4XUPFWGMEVnAxTu6V3EafmhG
/mym7w/lZi2C+ZAxf21mSgO2TqOep6Y2j8DCGk/q84RLVAYsIA0lahbmX5b7HjGX
E6oRVDEiXMrWX8XVfzMHJx/qpzXHyKl2MGPnE1sMsDiGaXCHziO4w2HUx/0v7iSa
V9JQ7uumUmKm1ADTeMqQhBOusL2htPQ7k9ylimpEYoWK+691/4qMikZ4xsnfIpwj
i25f8ItAuCmpWvPdmRnuzzKBXfulcw8uexpizubVWK++jkHE5bCGM1fN1OmPqK91
9zzX2u6+N0fDGNKWkU8rnkbwS4zCfBhKL/WKP2AaR1ATY1pN+6ft3o9aijFD0aZW
VDULU1DC0sdJw31QFohOou2LV1dOMITCimp/kL8dp5BAFCx6KWXJYAei4+Jlevba
EWCRVWBrZPMb0DnQHJRoQVBcFJ0EAO34oLfJ9Ml3qpCbdpYEwT9BJq5xgYmGuV4W
LedB3RFuVgDdGZjsDCQwAUqEUwnQLI7gmAm26CIAGGnc9YlYMuQL0hbfggMBJDmr
ukbu3hXo85rDpqXh5IITALuH3oYXSMT5bW3Jnllpeok=
`protect END_PROTECTED
