`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LBQ6RMlD6/5vEYfP+Zq24scm8z7toLG4HM8ZSazm7OpS9JxhJImmkLLNE2Jmnn8k
fP7fZD9XoFHxUuSmrAPu1Be5olwNVtvmWmK14rpvExI96Qk+hkZUSq/XeWfXHF4d
MX1Ky38IhqlL3rVWx9RIvmfN3BDTVocgRAMPePfC1H74GHGVIryO3oR6tMYTyMUk
4UmD1EYLaOL+lEUSkY/nBraM0ukPQMOhmWUGhUiUxGt2yVBrE9KLKDvzEN14sT3R
vOhnacp62TeKEqEeeZf0/JUFxFw5X7U024DqB9msvFkZwLT+T1MMkrijYdYXgF1p
u4bUcqyBKFUvHmEwj5+yrgt0BpFmNWznToAJ4ypAJvM7wR9igfAu+/9Asqo6oagU
LNSpC4nT7S59POJ11a8dX/nWMgRC5w1iYZLXBVZLq7I=
`protect END_PROTECTED
