`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7FN5xcQhSnLh0Fr24ndI4VhZopJ8Y2unV0tsOY1LPTa6qZDoJm+SB0g/n3bpzr6H
QUbEgaMRVT41VKwVWPCCc9VRzsgdhf4rophiY8BNyzgjS3sLjoJcB5XQ2cRzfAOs
gJ50gODo2T1Shmdw3VXipJGkISH6LNQmYyfXZsHpzppfnT5Syo/L7uAWygO0hc8H
pE48cCEi5I8lWFFJXOCk1VXKVeg6GwZ0m7PhTKycY3fb+nqLYMsDNuaevyRUNWju
+myHWtAiSe5xKBVgEFuJNhWqiQkA1xdyMrhjzbMJsbndsA45n+9cK069bXNIynAL
ZVqDn0Usmm3DPwBiwJzYn+BSS6SHUOhDpSakE9C+6C2H56QOoPByspuruNQ8/CdO
jDLvcgS0y9VIMUwc3bFEWE2QsVn2tgdNx8iEGI0Ml7c=
`protect END_PROTECTED
