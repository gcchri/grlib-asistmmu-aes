`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bXHns/KvbaPbxXGPwnafkqQTdAiVwbIqehvYGCA49UAhF9bRoKjbO27kMHPQbA8C
ZblG5pGOcvSRgRW91BEU8UNtZgrTJQdi8oyGjopBeIftr7ZVKNOhicSoqt4E7wuj
gjTF0gqoMv+imB+KKh+86Hp6PqmRC5b6ubGj30cdV4NMdtA8PoLkKyEqNkbAcOsI
e8G1dQtlG4jenaO4/Z118OSiJH3tJraH8XqIfyVGcqDOi7XfHi59WSr2PXv5PhsC
WV1rYtrz9Di8yoncR9BaRnIuqf97t11hH4DT9yP0WjoBqVGqu8H7UVviMJOdfFaS
hx+fMI4BH2V6iIknY+F9Q7/PcSiffg5WvVuPtmBP/5qAKwXSyrPdlRVA7ncNboz4
md2um1TSNDEKtZB7rtAeLK/rQddmg8qhAjuvezXOA1cVp1goWXwApFnyd2tr/49Q
uvhtKpdQ7X/AGA3YzMUwE/ipBlAu+Xcx5Pyg6dzd34iG/K1qDaOUxjF/I7igHvd7
dEd9CYcKgqqidEfoR5RkqIcvYmuRDWUkqL42DSMwBSxOali938NLAWU+fc3KBVlr
WNGo86c3OBTzzVmbmXxC9+A7vZFsyuDfQY46qVRbFLe/mgdFWC3IZ/SFgmfc2HWM
`protect END_PROTECTED
