`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4r3gtv7pTj79yj12CAXTINkGbojV6Rqe/dml4M2Zop8lQ7Qss00if6GyJLFG5i12
w8O57qCLLX1o7X5hS5KpDX+5vNB6ds6EVBQYOPXeq/mDsCQSMRuroV/pgx7xex2r
/Vl8K9YwbjjdeqxNfzspztJ3sBm2s0LZR/amR3AE6q0RFEek8IRaPkCXtKjAHPc9
rwEpR2mhddEfrIn8Bg35mOWghVuW9UoajpYAjVwIJR//8fR1++imV4JR37FE5wtd
DSVh2z5oZU7uAHb5lgn8H9h4JIDXIiwzYe9+IvHPNvY=
`protect END_PROTECTED
