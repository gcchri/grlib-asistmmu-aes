`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bQl8l0Jf+qc7HuA8qEjR/knTAaEh6+JxtVGghrrMJRweP7lONbMv65p2LLqWgCRJ
bbrzc4cftKraksRLfuwo2eICYQ00fK/uoibXS+w8Y048dwo/4/co7bDTlhu1wa0U
tWSl7T3Ksw5eGuwnxySQaZWkK27m35jyYiCo4i+sOppy+mFYEP0Dm+gqnMrfKb+9
k2nAYY73wlr8JJLEY3Tz8WQD+sDg8nmCEXVa7pUlTg070bZ3ilOvsU4Lps6ulkHz
ZVQhovabnJ91GMkpVm7knR0298XF7TY/oEs7IgGQ7QJrwmIT+bSzzlkrghNHIoVw
ahdu2pdqzzeJWite/iuk5ea3MBdRjrsvqSZNgbx4vgCas4ILnfIQjQ53okedK8B/
GcjmvughVRj+sT/dNQ2htSAEudgeYKLKBkYO7ZhyWWq/GDAcfysWm9dCGS7x0CWm
+/u94ZdPPPcXA78swPGqLBIrLWd/izkwXP94maeWX6E3vQ4czyxZEm97gzusKeUW
8repJ1QLz/HrfSyIdsH4L9TPe1WLVdb4FHoZ9BGJl6iaAh9dKNCFzzLQBNWRg1CS
oLmdx7WVbv/yob88x8F1jC/sS0xKw8HbKDoixSnfzg78d+rdS9wXL30KI4FC5Y+t
q7uDBBjhaidQXPjf1WUZaLAueUjqM0fw3H+D8+Zmx17hFfSETzBa8rrYfFg7UNdO
bvKrd+QtC6ckAXtba6rqEW0h3pKhWdQj51GhzMGSfiLWaTHeJIRoFty4zPBVw1fo
OYiKAsI7kd0W+5dX5TXu4hDt0OcE+wYhOo8L+ibP/OQv/E6HlFDrBb1RtVyuKnrj
ddknRjQowH4PGas5iTEzDx0NFYN/1SY4XfHqT8Ay2BHTbcSxvDvuQsPihDwYnnKo
fxDPdBS31FeS9GzITWfVbcauM6vzjYaHmCXcBoMcYl1WxW/eHBlKiXpq58CzZsfL
XFyFjDez/Jc1DeQGh5p9pSoOieYb0QsaCCbvxFjwmTGgc/B2Q4hMQxk1hpYhn9iC
89Hpjkb/JxaRtfYujfVdK+9w5q2lqHm7yJB9ds2Pga926AM1I76jslyD6HMpJQGG
2hMja0+s0R+FXW1s+V+bQaNyeLVISxaoLZH/LsQLdwvbsZJvKmEC7jRzuRGFF7tt
bytK041vzMjxjpcQxVPFUPUAnbjAoEp8TsVCqSs8An1+ykSxQRaOgX+7T9F3S3yT
tUz7xM1nqG/1DI3PVurdAKEh9hB1UkLd29SQZWdimfvAnX7l4w/9y7vOgvm/ebzv
7dtIpEafuDnaYee6ufl+BI/FhxcaomRPfCwO/sw8Ppww8llzy7rNNOZIpF+IbeFo
TsIY1FXCg8+ieKrUDhJX72y/BO4txLdVjN8toiS18ybDgF7tvv+n4XSD77rTqDtf
UgterAu2Dd7v7/3phJGZWLub0Pu8sG1+h5z/hdYaVWhsl210G7dJS0L2Xv2Wjbqq
bmLDWlXhE3Nds3iFKnDH0AjNjjnpjKe5Zlu8otdEmOf6Fat35ftBBBYptaZ6win+
cY6ys83JGUAiCzGjnxFNQ3HfMd1MKOmtV9re9oOMZo7d5pMKeJDXnth4X06NCtvR
XKm3Bm5Aw4/mIT2NwQyGmysE/ctZlBDQXnsFGGqLCJdLaljgqzUwZkTDYE+atw8B
/ku7KbVKL7sgl5LaOFmU+0ZX5KP3yF+7uO94Y8xGXlBR/w3dFNSdCIX+EAKTD38L
GknqYyl/1aowOzRy+slWcEOElnaGL4GMBtxsb8udmrlVs32U6owdDEBTFJd5xwXb
DZFPcQMOtHPP2iAe17I5u5eDl01qdb1BxdYxGciqVZ4LcXvPkqiBFrnDuQJQVLoE
zqOOOGINQXN1HKJpv4j4UcpbOMRnugDp/dk1I2fn2qKlR/DKNWeCbgUVEwa2ClnZ
jtwMb2jk76jbIDfkVvUt95zfceup9UldTYFvByQsxK4BSFUb6afOYQV1G6Dn4kx6
FedXyK08yq+dd1YLJg2ALyojn12HUtQ6jHXCxHpiq2oR2AoON+umWtjoDCKA3tbj
LERiuk1vM0FHgi4Jzqwc1OHbF+GOctciCgqes90k5XI75NZtV62mmpJ5u4kc5dbH
xo1p0uFeu4vy47TBEuSZpbT2CmTnkm4qUEi+PkeYOFE4uUAHmLg9DPMqWxSYYSmB
VPSwwq/rhnjge5LqUIv9hB0Ie9dfp4c97P5y7Ksg2qY5p36L3jTyCpq60LJlM1lr
AxLAcohoUImXmROoswA683US0dm8NyGo0xIF8UkpvXd9YhtIRMBrwlhR6gqVS82G
4A+pATwBiPNnuMI8RbDH8SiGHw40ENg1YlT1bT+3yZkmTNit416PzNSI0WFqbUr5
oRlUH4OxwdUwu4ZRuUt/+31NQwMDc4ZkqIhuBlFOWeUDZ1eKFlsv6yzrrGNSImqz
3T8Yx8CREySbVh384qFgXcHKunk/8iwbTdSfej8g1XDK673AyD/UcttWEWAuBCM/
7dtRkT3eUxAD0V1kyf0YY2e8k0fLysEmZLW+dpJsW4l330W8TFqUlKeTUVx5NaDB
Hnd0L49sgcfF/VS+/0xdhpyKByFoR7ak/n24urjeCIbU1w1vdWO9Qx3ckFkk53s0
/RbGjJdazuAUs3iNsd/IPsuiyvMHrminiyjRKnrLCjOJpBjAl6K8OptHhCQuBCRR
N2XRVQiUzaJGriHSucujsJu/uAviKmQTiPYdar/ffejJEfb19Ys/TEK21tC8ghQB
t0fVOEg5Pqmf00MwuMYQkAby67/LC5G2h/7Q+Epyls8NK0R1sS7+Wf4unGqUZHg+
+XUNxQ5O3+89SouGEzUxDZfRlyslB3b4A1DXPFjvRfqBWLdosilZ1wFtF843Dyc7
5fsOuN0AVxlhwrqmCQN6Qz1A1lipPAPoZkyM7HksAM+k3vpzoxLNizhu31Gv/FEL
ChhwKqOQI+4JJ0cJYJN9B6fBDYqemULXBUlWe0xbBeZ6vsNiTiKuXi0YsXqrEBEt
U9+mQZB8VxYrQiv3wY3Z4F0WTGAKJgczyBXNf3RIdxcfbQPcr4waLpNYNAZraSD2
+jMq0CvwBxzBbrB3Zw8w3OYi78B6xy4Q9zBpGNczohpdFSA3gYxboEfX+mglXFwj
vzC32AqbKu+JOuV7kAnaltWKxICw/uUHPcnbje2+iDYqLMjkP0wiXpqh1WKTegP0
1VDS5tzm9ycWgRqnoD2P2kjJ7GUCm8pwXkCl6ogNXg0an3nWS3ON0HNK5IzAUBox
10f/OGC6ElTgeubNZRyz1uDrdieloOQNfhYdeyxIk78/mwFxtslhr/zfO4RQdS8/
7w9gpGtYOcIRcPccW/4AiFs7EFdZFef1kvh7n4/Zj3ynq2ZZjf1Q37EgC1sgJSlH
crNNp+x5zcwxBCOBWgWv+sJI0qbnIdfCJJP3NL3+PH5RUNl2W1X0WDVfTkTeuLcX
kLr03ofI0bB4Ta9ujkHpUb+BCbcNjXJGenhwGOEEQpjxluBJaGYFPJdu3qI00e9Y
ZOxkc/kLzhmXUV71FSeXghtG07oI62NQITtEDQbKeWO7yezt4VO5YGyKN/PsJgji
iRkughEOmZt2lCPAhF/Ur5QDFUpYtEZ7LIpHwc4r70+FO385XKmqL7EiNFhn/A5y
/kCt6nBn5S+871cSyKy86HxYMX8nmEl8ZGgO9nlqWB0uKy+rf2C0JB7qLB3Kl7rX
Of5kPFebHYs//3ftpYMDup4F3tSS0fBy5wiMUUuu7JI0PCz63z+chabvwHdryknh
fPemcW9B6cBvZBjodn5idGe4BNwliJ+iCXAQiV99am/q8MaNjxyee2PiPijW2/Wx
EFFxpWucULKVPFOz3gwJOICF4AD6L5DbEbYrkLeDd0orPRKakTFhz4g/Sty/tONL
aKc7lBfcREk/Ei55rLc1FMINgNvaXWdTdFyDzJoWNB32Wc49BZTa7TM2VjtQIf0f
fR6FvnjD2efYf92zf0keByD85p2bd5PALqjpktVcToMaf2z0EozD8p5AA0foptNM
BALv07/ZAHH4pVnMKrkVo9f88cIDxM4fS/0ZBLx2HoLHgtToFOhS8pbNjU+ySjOc
Fxxq2hjWLuai8HhbOSsd58nWMz+IatAibyZXkZWk0B8nArRXRPdOlaKDc9+YGN6d
BowctkaWDMS9A5fLBLE0aRDsQIcRZi2tEwEkA53whFZg4IOhGETJ4FLVxhbYrRj4
8fIzokrJMJNhSU0wTjNqShdzYlGw/M8lTbOnjFFLnW48JSMk6H2BEiObzqm45Mvn
6qt3f1TLVM42O4hUBfU4oR88Yfkq7+Z0R/BngeETNWv62S5sfn3zpi+MDAJt3BNE
ECxTlq8Jzs9117/HSdvp1BvHryIjvmV6iaeUBsYODNHXUME3+g9owJj6KxRDhNbA
znMIW+ESgKLfgBhppaTOUaJOLTqsLmyJ7hJmj+ACuNzxc2jXY7yYqsjf/IfjfKqb
bzFDFUukIcgQB0+ELWeXQStx/c71KxekcFNnSF2vSh0PnGUKizX4qSCxUdHxLoPP
449+lYMBLJAThdj4myIqv99jC2kbh2bm1EIObzbf11cHWMim4rz8WUGCiW8deQlP
rxj3KGtt2ZDCXF0HohnQEHdGLPlZzCSO9VH8LPbAJrbf8ML6U31B92pdsvu1GNC6
Nk432K+F8QZglOhvraTRK5iqht+bt4U5qpzQEGd/C6qgFVQo2CLJqMf1l5Wt5pNi
XZTM5QzK74XMhS4tbubvHoooYIv7gFyMPqaGfQ8SZsrnN4ui91RX97HO1RQnUa8n
nx13VCQYrsU0Sw34RHgO4/Hr5rHjiVVMLuT+Hajon2QlGHrzXrN2bdU3WO56cDE5
O5glsSBZf4RZOJh5i56gur1Ytm/sqHGh98HwCd0VSIMLCTps3/4Asx/bTXY4mXIR
c7ZV9BZcVYpZr29/3sne/j/mw2Os8yHzslScFgL3mxqswXkTB5V1mA2fSaVHTooV
oWGDOecPZOQrcSBIBTiRI1LZHDcJHG6Dj6G3ibgXnBgxZbMuzNBEz+FcF3qYvWSa
EAw6IKbvc6phxHjK2YNjIy9EquJ/WBDtkouw8NC1G4b2SoTq10WaiJCsVLe9WcxF
ihbzJaTsFFDOtbmci2thbWVxeBBIUq2LLqRt+Iquuat89y8mN6GYR6RZFFd8fLSw
YxjI9FLBDjXN/qVd9Myc3on0pVfmJfkhb2zwfQceGg4Pl+0QZqw5Cd8NfYDxWgEW
N4TOH0U4nnXMsndqAp3ZfsHs0ZZ3qNjsHqpxAX4YHlvZfXNhXQLoDsfBsesISrHm
4PGpZ6JKyulBwrf1JH80Xw3rWgtQ9gNnHdY3963gV2AOtau86oILAx8nkmx/ITNA
NXUovb1XA0L+Y0zO6svTRSR3xc4CYLQBOBJ1nUTNrN3IwgHLaayE/8powcR6dvBI
AgEmLYi/LxEBInnBB+CKvOMFsOxhgF5nRHZ845AuSrnNkBKm+961lEDlYKBd/XgO
SUsHWYE7oCZcXR/165qp7Tb5VKr84rzrXLQ6wSHAL6HENAVyh0rJI2CDp1wyZdCH
WBEFSHweK8HlymFjK6FfExmTBVOeLP2DiuzmmdOjWCr/rc2FUeq9Ne44WgA+YscP
V3wtDcXLbNIjFhhulWHZKDycI95C0yS7k+gUyDpHyMq6qpW+DmUvJckfwAGhCf2w
N/m/nbQZQC8fkjruYe7cKWZR/noMYdTXX/O+3di/pABlIzMGOcQsvx86Ny/i6gXk
zMlpKz+cFMNNekHoVhbPtVWNeja48SNqE4UQekrjCqpaQY6YmHAXByvZ+d9yADcY
O3R/zE2McLqh+1PJFUr8oXcubjJFbODwQPItEAmq+uM4oMNOnjVJrP5BEOWmOf9w
Gt3ela1T6ZQ28pvkwhKj37oJBhSAE18OEE2UZEpTQpdfUzPcL7lkDJKH/FwuYJey
7gfWnMX6eWSNdp11PmhQbLWWLXrTI+8WFpxBx4bA41U074x3Lq8eTEFK/Cdx8Ldn
vnRX5hBJsDMzLq9EO/TsDfaEbI1uqvLie8qtCHdB9jGk1rS5/es6YxYNB102hAbC
ghmd7sFJ5L1qiSLG4W2TwenNwZ/r6fdp937bTexbbr4mCHz0YjMn6jeRp6m/YEll
dw3Lmib4xQPj0QRaJ9b6evcqwBYO5Ty3rgzjPzCnpbgU5q2KextRasNId7D6MW+W
HSiqwaOx//SXpybtS1Qjrr+8PE9NERXJiNYke6MuFUMwUjFjkj4LuxE0tBlD/5T0
BO658Od8mNcK+l8D8QNND6kdKf3DXzbJEjXULZuWFWODKpFX0n7JRpKMa0deEP8E
KOVDS5eGtinz1M/Z8Ifu3Kuy7k/wzZBNXRAzVqSCm8SnLMmaITiVFIIH12FHTYmD
TmBIAKU5LPqRbVg0hTf+q3M6yFbyBg8mDv3kRKO8jFS2mPxPWWFWReagmIAwIP3V
WU3Ms3ZSMy2n2FZldgbI5GwDKTkkOydaLC63/75kRY7UNsQtC+cbFlcGULwTU+YH
pxigUHozPVoiG/Znth3/MxI8yepXyrH51sHt+kPoqlkN1Blkdq/JOHwMGadia5mq
rJwwGVbY17SBKt/g0eGfCM26dG+zyQ5soV8Qkea2UMCTtNLFgSETj7/5pUYQFRHn
RL/rfSWFknyWtj3Xr3+uc9S1JH1y5+K+WXldhZtd8dkzcfQyI1Fz06gDknEHInkJ
XACcPoqrfRPZU0xjfnqyBxcVbyV4yADZAysJpzFu+nnfKQvwVnhQuWmm975OsPBc
LGKx9srUX/gMHkeb7mR2k6ruSXGJOaZY6Ajm0VyDVHbAoGo7u7KL6w2zoeVrATj3
2QNJDvq20cpfR2h8atfoLeCqK0yXsJFN4t7AR9AecP2Drx7wxYqI7NdE8leqq71+
CN7SOD09QyZclaYv1ezW/QYOdpC6VYn5Msdco3jWiVslEJTJbuKJEohoUUBeuN0R
ccgE6KRa20ymhhTE8C39PkNifHRN64+zI5k99EOcL+1HrWuIMdyfZr793Qr0lWh+
9kDJqpMx86RoKL3Vw9sS+bhgN1rZdgXtR65WZ4bGAWhW1aWm+hokxW4jT57BRKjE
N4GmO61RwTjPHgbPn49Nj/+d05TwCrYXXbndNuKlLG0bkQDs4ZrDB65Rv1dUrh7T
BBsyhYvBv0UP4Xxpl+IyYCXQwqYdzN1oJSP592IPcgVj9cKml07SnLH9AiRvc7AM
sL1frzIWed43yP71PvCW5PPFRAtgjzehAKQyz4gWXxDMuWI3vbwW3vYp04S3m1Y1
LizNANI67ZMjbJVo5OjbAY0/od2GLYSt4SW/E6NNC3GpmZQ1i4iV8bx+G5ngFl4L
Bb1eb3b2Et0JU2b2KkkI5+DNlOZ9avR7Wi9pZONOc7P8y50CHRvrirH/qy/QtVwl
aYxrBwus/GW2sb8LD7xA7BdSeXUdSYhhFKUbtOxCTcT4F4TYV0wznBhoNw5fP+U6
ie6FTj0up/RAxSErxcDWTUIrInhMtuabaDE3tahOQ4XhnApJxWag+6ZR0ROeweb3
GKYlVzh6pNlc+sj035HdOo1KcJ6TVOKEUl6n1YUNBfD4z0nMCrmq2n4+RIN+pOW2
Jf2BYKdMhJUd7tRfK2JLbA6Cs5LhnMwe53Ad5qc8l6PIf4HW0utnOxXmWcG+dPkn
fhhnURbxpkuMtWf1asFBuDCnUdXty21UPgBs+YtUFiCFvK2iqyUMwSrX+/3fmMsA
FsZ793roNicIEunkfdwd+ITvsjfiIxGaQiAld6OfBAlXPzsVrd5vV8tYK8Lv1jUf
Bi9swpsJNbKCGF1SeLPyW5FA3hIqwVPxzVrGrTzdsMnnZbbLwP/nY0f2VWQUoLpG
4m8fgKKUwXHud2O5WtkdNJNhogw/HMkOiSQ2exIyj8yrJ9D0SBBSQkTjTuHoPqqe
/1sTkzlKzK6ZkYNE2tyZRfaRDYB9wRKxgZ9WbWwjCS5xdBqNCOAhdKXCh/s/qJWg
LSk16KYu2qIpQBs66viJUsdHnp1TYk2FeBuoP1cByK0p+trvZuKD95bh5Vbk2NCM
DUYIUh+4d8wU7xWHA/llgP12qYJGPADWXkFZMAZQGJwb8UWMuTuSQAzSH9ULjv31
2U9Ea4lfDgslhv05BlYldt9SnXNB3PaAX0lXH4LfxjC2orsI0iu5YO77M1UTElII
yTlRmYa1lX1Vy4ENiSxiwprbAoSiQEyD1wue8OZMSQvwkpN27J8WnV3KGoAoMdol
hTKsuak8V0YTpFivOXVOXep0u938Iu/k364LiwRNWGG52vzZc7e9ShNstVNjwce8
vF8wdicA2FfYHYQ548KD1u7pVT4lyo6Z3rgjC3mEi+3flAQZXYolTjzfvYbtM5NF
Tpo+aKtaZmwgXd6HQxCxEgEW3byztL2vq4iYuwhWWRUNSEWQQLLyVa3rQfjZssE1
1Je11+rQLjjkn5jJ00+h/5MItERMVEc8ymf2GKNRBXQ5bvlMvPWksD5oLkGYxm8w
eMu8T9awi3rIpGgi3UhIxiJCLe8OLYeCWVgTJlach9C+VUI/mpDALBp/QbXMIOlg
uRUpZiwe0phYP6chRr2o9ehC6b2cnE3rru3Qb2sIGCFsLTgvchpzyUyjF4v4e15U
dBMWe4bBIjNVvZnbzB7f6icmN63+oGr/iACp03AaUCizHgwu1ogbbEbDC5MPmepd
Z4wOELqiZ6ox1sdRzSGcl/fomNTOMtljI8r0NQhxvucB+x/kFjNnHT+n9u9oIM3P
SKzHB97SXGPuubx8TR4znCuUb3ecjENV5i0iimVUQHoFXuaN+5EVrJfPev9Pc9fV
zMFJnwWldgPVaYl+ZU22Rbs0YK/im8EI2tUEM7sdqg3xkiMzrr/JRvzRdbGDdQ1X
IAQ0KDjHx3jEC2Eu83jIGg9o805H+bFa18eWM38ziwT+5uhDAdvU0x/tavMd4Kgn
bRFnhNqpvprgeQ5x0dJHlahLI9HfeCZ/wJ29kZgPn/qZGi6yT6vUbsgn0vQlRbyW
P1LyXRDc27RY84Yiu7GC9/rQiIeWtWPs/q9G0IN+fZ8mwrvFQ+dctuFe4co8wBn9
P2pVnI0F3HGMUVqVpimh+W8zDD9kgYePLWTyRQqKvh4uaN09jQs51RDM5HxMs1SH
iS9PxSSW71KOtsqpULv5h6VE9fk+UiglnJtnRQAKQ2Tf6ENum9pH2z25G6Xxz/+u
AN3XwfB/pjoHxldGbY2Z5JysXoULWw7noBBE0fvxgYSFFs0OV4CZDaEmKY59flqP
r41fBvxgW3qUdO2s7CxHve7f5nqWw4qktqHVTS2O211X/zBzaQg0vZ/Fhkr6Z6R4
WvTccNRDKo+JFol9vt+pgNqCBFWBBsnNJEn2+0Dps5Fy+bCffu/g5LKhyFvoqzSV
rWoK5U6oDTI0A1K4tr+OPI17s2KLnPm8s47AumyeKX5r2EfRFqjLVqMmqHhUsyig
2tLXL1OZn8jitvwCX1Q72S51XqUnVDBqc0mGHyrdhw5OojzwaCetdFgjgd7YoM+J
uYB7CXeeCbphkcDYp3Rl4+Zamkqj6IR2BGwyfjWD5HjmxhSE13xo8JT7UQ7GKWHC
5/GSDkPk//go0YMiqGaea4Fhi+Er0IP7ISolkvaNZoEhXrWrAweEWGyZkXD+EYdR
9XuBZJp7GIry0E2BaGjFcX571x9w/xhdcvOAG9EOgEXy2SXiISMvPdf7X6FLZ6mZ
mMwd7QhOf+ny/RRoHVcEdg5Xyz3+zWU0XpZR9kFGBpHS9Tv24WkmQGsQWgILTHkH
+1jI8Bst/Wv+ii0wt/bZxS8FyZxDOf1zCAc1v9nKTv4J6bxwJ+jBBruv9/UkjV4a
2CPWH5prSkl2gDT7k0uMDW8RpZGTZD2rBPT2u/UG3Pc4iQ/JeXkYgZZSCtyE0CdT
C/1evo3MLIWGZXYKMdEVMC77UBgHqFLPkxbLXO9suBcXVicNCaNL2LqVXBJat/DX
AKpvpeUdHbdnaObfSSEKVIg6gZP6xGSIcmFDl1wkbSjWWbExiuToqLzEFp8l/zxr
ZNLAa3Fwdk95paIMtb1RYf1FqvnM9I7dzLUTvvE2r0RKvJ+A6Hfc+sX0BXZv+74x
wWbsv08WIZtiEaAdFj9K9QTXfdIfbKQWz4HH53dSGepUT6Bfr792LLrHjAWqdZht
2nbnMQ2zmHNHxeObL3tL/Yxj/81JpmXczL6XU/4G2qzN7uiI05ZRO6c/FyX/w5CC
G4sPjh8lyXdJYEvhJSDCaMGtCLN3Kun/NMYT4dEao8Wd3R11VYhjdVN8DnHZ/oKq
t/rjjeQreLpk4LsiPjUCCJlz5Hf7JJ2esGKAu/Hs1/NYMNc7v2Li8l6oNFt73NMH
4Qak9PB9KZKBzrHJW4lGvOQ+7BmJMJBa9lUf4LvJG3kqfo4qucTTN1fjXZojpQU2
pEDQj3YvN9YmDDmdDLGx62VC6BHTpJVVZCL+uOGm+xjHkuHcmg3CX2A8j+6MFHG2
Oalp+2IlglJbxo92GnHv9cCXAqH4tSaxvYGfrN1v6+5/nPiomt4t/aj8uNrT0i9h
Uw0m/KmALJNlocwGCC4ON2O73fYiqT4e4udzmNnFpE3pS3+vNLxeT5zbMWzYqO6U
bOQZ3tEGtNHoJoGHzCh2EC80rNykou3ABxna2dHQOnjvWEAj97+6dr7af68o/Vuf
7vohyd4PT7XTTUWJsJZKZaxaon/mgjBkbByDzClqTM4fhnOLKeK6+ntbiGyX8QBN
DmBy2Jj3FGITTzRZhfA1PPPX+5/5ShQDiSRZ20kclV2ypZINPXXmWNcJV6z6KZls
y/mejGqDis3D2ju/NPZUf+cX9OSaxV+Y6tbDk6yUBjhSXAtgPzcJ0G7nGiNWSA2f
4QtDIbtd5YUcsi4+jCs5dqboa4yBJODrccxyfugBYLW1eric1yx6M7MQma5L0O9U
g8b+AHH/DJPAKPkaecmIuxbJH9AZJqlYrJiQLcPpIGL3JdIdz1YGMVK9NnkkfGaa
AZYpTaqei1pvJjJ00q9y1aG2Y03ogQtXiog+4yYP4Uc+zbV6+DKqI08utnDu3nzh
1lAPpmSnK1VfqXcEwOA5Xyw4QXDLvStKmp0QOSDH6xTPKYAvRs281HPFxNyUvAKV
Ze0Fxz1yHRs/iB66cKYofFDynmZl/FydQXWq0yhshK9Z/AuPuhU1lJ/Q7z6CiNbP
ctofNZRf4CRo6Xfy40iB0aw/pP/7AirwIV5a3zcC5x9BxTAJ35k3TiAXf+bD16XY
Y8DEMZFUs1BuVUyQqxCXP08VrX84DiAnWR0wrcXSxIbLrSwF/A08gwoAY4KL3u94
ZgJh4tC8caHlcmxwMsU830uyQrdNofFK2hiHOds+ty0kGAvioWfrZQmw/3e6BhK+
kYXLDK6JNcIaLKHtSa/UK+zJcDOQ9EG1QG0X+ytwaeJwELNvuOukNcVEICkV4Oof
iwNp9BGqF9TXzQZBdgg8LKhbrqE6riQGdhPavxW6VyfqkVaWWm8ypnCK+T8aABZy
w5r0mj2tBQp3Yu7iEAVzPVKOIU7iBuMAi4gKjQpDVOHHQgPdNf2w9RrcAvz8Hzm6
4vkuV3yhAcgOQ7loZITAMQG+IRQF8tiA8M4Ak52lqWc=
`protect END_PROTECTED
