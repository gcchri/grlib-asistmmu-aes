`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v0KeGYRtttr5M9hN0jZWCC+si7j+lx9l7IQmH1xf+UWmhqo4dv0sabxaiOowQApF
OnJmAmPbP2DTW/NN833SWGusD2ZVoo3Cxbs8GxkfjgsaN3eS/lW2ZebEA9cbNkcg
SYrsARPUo9+HJ8DpYaeAB/Y8id5Blv5/FVmh64cqS9kDxSnnO22u4zbklZlkod9a
foudFDXrKdMDqXzQ0UY3XUmQzZ/BeqsEQKlStbEYf96fsRZrsD7AxWv4RHyv0hrS
uN68UfHYZdjH0qFZADs57PX9z9lfkxjIp0npyishH/tuVh10IW7eKVl11mlLxTaA
ETX0qLhgjgUoO6QeMtw2sYHfU/lxtKorKJwEcJWLoTec5xQfZqKvVcLSx6PlUwUA
JFIsNs9YjfKfpisW/EfHKsygwGeJvqgmU9wX8Np5lWigbavpvnv5RZ2FurQdDik4
DGerdvGDrlzjl/kf41/1OfKs/2POkdAQ/XGd0yT2/oIwKwbSVTKh9m92jLcaEVtc
deHpQGw0HcgQHNXsvHYfCQJU0KXwjxLZ4b+i15P+zHShiUqG3FwNh5lftAUVom7H
ZaE2ptJIwjWcMTx+DWCheQqq9+1euqfyVbNxX+6CF26brzytvmVF3rMf6CY5qbAM
yxArlfzYywLSZmJ9zA2cGkumAmsDphDmV4pTi5v9LYOqrxzsXBusUafttE+a3UAP
TE3T+1hVVJxUja3hjV4TyQ0W1xnVDLpPCi1Jzk1/aBLI8+4Jmnsch12E73ccYvnK
E0yY59q0F6NHXCFWvSNMERtpHYhvg49w4q+rGr7zSU76+Oj4l6fuQkrbcGzugSif
inCa+15M9Bmxywn5JCq7pTb3ADZ+mx8jky+dXCj+ecCX5JIHo3adKgjQM41p/znv
ZmymbPgW9DgUH77MSSP57YFmx+sv75Wb0+FD66f6IhkDAqM4z2KD/270in7B2F+z
STGRYX976hJMQDOO0yonR3BX89SEdVHEVUandm1IJ7pDJvzn/EDBT7poYsc+gZka
Q9n5kIFvex5JikmTCdjJGgWJM/0CGvcso3YfvbvyufYD5TD4llXHgA5VBnzjbwAk
nq1D9IlxU8oIM06+tJLcNbiVgzxzcAdBE49oSkNz+r+Q/dtS1xI4igOb7q5ouBkp
XDgno0NAwJ2JOvNBN3KTov7FPRX2Tmx5n6Hj08DWWgUUtpCRQMjsthAP0x4xb/Lh
SaopladgqywC99chTjcloFnuLt91WnMg8Vw48NbsGOh87YxvHDQx1DpmDDnWOOsJ
GsMOS6kYPgjhj/wB1emjgwOqPWV+AQpQm1lEivdcNCRwfVqkv+Xrn0f5CRxdmeMS
1cWYtXgm/8oa5vGYHksxpA8Pmphqavjp0jKHb4NDadh2KJNwPQrZe9DuP5wvP0hY
Qr7UxOf6vjdGH3+LHOTLVn4WLnSdUssZ6LhrbWyDlmucKdZZPWrGse3ynddC0kkh
YChyNDcZSE8591r86mltAVdtW3mz4LebjyZtSnVuC2xPsbQB45k4E2MhhCn0Bndq
99h8u9OhRXZvdcjgigh4Q4ITPYT1SjnWLsqJUgcfLbktfsqvCGINfecDC3lVm37+
7ytcbABgY6FyBpgSHIZ3okjmI8sGBACDWl+atyO3ZGXuqiSWKw6+HIq5z5BjxafZ
euqsBp0OnkaMovrDpk9Js2/LbpgwYy+wTcSTdCra3KqdybTq53ZuRLDTKelryP7v
2kuoBTX3hof4T3hxxGDYsEOvJ56nUgq/5RdaTkN7J7v+YHrXLrdGOM8xCiiFIl7j
YD9SgwFsI93frnLYhvY0iR/RueLbY67QaESrHWErKBArVT2mQKJJvtZvKhRtQNxh
DNIgncR5fIMb6Gd9IqKD8U1OxXkv4vnMoRHqjyn6kOWy+85ZAlM4Yb77/69BwSLW
0rHQfDGb1Tu1qirgySOo2u3TpAERZeJtPLp18AWVtXnDywq+Vlfi22STQDEfVeyQ
WjNwDjnKdqitff4THd6xuohwCE5QiqZXxEMNc94iVnhJNhNOiC2HWl0ROUvv4r3O
cmQzlXrTZU7OuLLXaE9yCd7duFsIAFXZvjO1wbQQDCBukPFnK3BYRGUTi0fFTfFN
nIVRk69gol/dXqNsMix9bxKKvdPT6QzF+orH8IPN+RamOE8U35PiBIpP5mc/otVv
M6g4mukWVpdwccStG2tnemdaMcZULxwKXGgcjPqYZl/NXpqchAeX1oiyKFG9+AR3
rA3YWfYD6YpT5lLAjvZlEryLE6/+GrtaJvL4vKomz+ZCH7/y5hxwcaAKEra5VpOU
RpFCgIBfLUsNrOA6wFrB8ZwuXAOih5W+7tuEi3Lo/ai+DvQ9HZYfvckj6Ci1HL+D
oHEGM30y4czsIE7IiMAsmKwT6hspXolDY2TL5kjkSv4EkIvdbzzaZ0Zdk+T9knpm
oTjugJ0dok4SSeSPR469kk4ErpoblcSlrRo9936ImHdlo6sSc2KQk3CzL67VYEfM
tq22uzkIUIqx2PHhO9IA4wE0cIGWWm96e5WaZZsTn6MJSqLNxcJ+6U2vIl/v9IBN
k4aRDJVpNWCjnufXAz3OykKRDcQ/Srx9bbsZ6LixjQnIogCRFPw+WyeziQm5+/DH
J7bre2/+D0GpeMZbGd+MRpndhwbaPRe5ptdAtl8ElJRJBbuks4+7wx1kwywR6aVH
kcmCk4jIzbTu5eqcv5jOBVyBrR588OkQ4XTY3tj4ndjRAvWTLzd449kMmEBheq9T
7pWnPn0mKfOSrV87mil6LZkCe02/axe41TdCFTL7x/vdrTPktPW3NgDNgcOEq+oQ
qxT0ps0me1UQrBX81dYpO7rR1bQ5Mko3CxjXMgrlGIyqq5XKlUCaKQerff9DlX5i
wOBB4IxpOlpBLEdwLz1FYnN4z8ILeCKSIKx+nCy6AadC1ZzaBJ9gtpUgjmlohjx7
MOaSm4wf2myMgkvQbJLZDmUAS+IQ1RlWCTCW5qRrjP3jmcAwv+FlML+aSjch0U4q
Sza9HWcpJo9wUzRbYe72pU4lNYyLR9rsFsqUznPMWm+P2rWOPP2KUpyp9xtNIp6l
oJf5LSW/Utvb23IfKOwVkRrEQNU5e7OCLWpCi3YtYEnhO7Wa9AciiauX+ct/5NbM
J6PG4Y/mstS09R635FCt6C0oKs5QnXpqDtpBFwzYyMmOPar7SP8jcKWfCdyuaGqJ
TFO+blbJAJbo1u5TTeZbvf/4hTtItroubR1Qvca1TPT/jhW9Bz1yxn49jF0P3aqM
gj4rgY+5xJ+gjiFVtuRmMj7BwjI0bfL/KJmxE07nfXBLz2MvDRspEULFqPU10tmM
rtZksDOvXpNixWqCUADorG6EdwBK8S4VWhBANrApYzXjTdDSI8b1DxuE+sPeu6mG
7NKmrzrWR7GKWpkwLEZgTn6q4hwi9XQQXF1YH+7MD41AnKzzDKJh1y53Wd/gV8WC
rs17wXu9f6OWHFTrpHjccaHmTTg5iTsWMHUpBl9dCwD3SY7ikrAxdrFH+LdthP7V
28TnPa04QI27gK5mIQ0adSyRUqL1EfBOzJl+Sy6nqIuE86a6UYjQMNmSqWRqCumh
N4FJU0lqOnq60RHP8CAGaHExKIDYLbZH8a4OgWGhmzCN7I2FL2aJDTlIz8HHA55h
t5QQbgDV+Z/nw5AgMJi0QrWauGYomq6hWfvnCCrK6V9RkX5gWplIJhs2DnupcyVO
XcKCeWyPEgGObRKGciKlk/A/9Q4GnQ0FGHwRPSASPpJpNKHZQm3uznkxS/PGRpma
MXS5jVazRetjQXzcoBGkt2dTNMn5fiZOB86tsH+GE7px4H5thGYzM6YREiSc9nuu
nBSfvkiwoEESX/sIwRq8oRjhHuf7ec/VZ0hdmVXfRVYz+EYVVk20RriWZi67fxrI
pMXEGBVB7qah1R6ebHyGyjrW1o3VE6G0bkQB+xQodTOzkvuvmtP1Jp2HepLEFRMs
kgZnXnSmoGQi2kX7uWNvwy5/I68LK/nYEyGN8ilIh98YEyzrD3UEErEP+vVdK4uN
bWRcoGjRJ6C2M/3p2I9D8ych26jJL+6urdAHpkt06N4REcObFJ5388yaxrDKTQID
vfQytg0lbCfwa7oeJlCIUYf1V754qmznraNm2EoKSZEtgYaAw5zh9dOR+7Qx6XQ9
5BbPO1Ivyt7z5eP1H6tPCBXB8dCdcyyxXucqzZqoN06+HMKSneJnZAhhqS+huMz9
OW9dtNeKU2Qw/VsZNttKKOgiOKKeZmCIUlHLYxZo526Xi6KoHyJtpCfaLVJN3WX3
K287EDAqAoMzJ4VAJFZBtJw3quBFw7JxPgRb1aSle94RnKpzQVjj4TfyJLiCFgh7
UdrQAOUyZmV7/i2n4Z741ihNWY2N1SEg8PXRIeEheZ43lq+35brqzwMZ5Wow1jFg
cKLXpAQdXQ9iUzXZGFkyt72MzxsvL+YZSCA4DFgyz7kakTvg1Hd/B8DqozFfW1tF
clGGeZUL44TysL2V4YNjR6feIj0elrnfvaM+4Xg6pQsOwvk0NhANzEbRtTqXs6Ey
V4XIU69MjHiJrgpt/Mqn3kMdSxvEfeWpM0I5U1A/6S5waymAxKCmNv/DwhCZX8gm
pzCjhPNa0/AklY0wusu7Gt5aF/Lh9pOW7ePj1QRsS1ebX5UgmhIn/3CYJOaYZfXE
7VCaFX4HMV1H4foGFSSyAXf0zl3UugQcTkieZCCjwt64iesgs66rIMrZ3qJTG1yv
xnPmgeitKNHbAWzZBSgmZrwUOCbDupPnTsWHauSEB1ACeUF7HduTKMAqCo43OUZm
qZH6mPURC9DGxTLt3STfzM1XBtNhGFRh5f/FynpmXEcmsx4ljWJ1f+wrENl8r9xY
rNzZNxoYlPtZ+ragLo8b35X/pYm+0OxPY5LCKkIQ1dPiWiTle0e8UZXp5Z5CGb+P
/MGdiPrL48db2eOgZtCkSnbuDUmqSPQ9aztp4U3G1I46M0y7YC+FLhau01BRkaid
FUJNE2xXcgmKaJGKcrNFrJiS/7C5EU7a+/geF+98eXl4Bynm0ae8Qn7d1VoNuBM6
Snzczx1BlnlFCZaADV8WoFNn4vQgqp1FBs+vpmGPfjb9TatEvF4HEDBVxKxviH8l
T4yzIyg3/rfTUwcbjs1FLw4sp5lUP68iX9YQ+AMygawFrotgk8a2pf1bXSR7X6g2
9Ae86/20dOF9jQg5U8/Rligf/Sj6ttpKuyrlRUa3tpxm7sGCz5HxGMop2AF5Q6U6
FCFs6XdMKGMniukd8c0rJ2NwnNR5MqbBRmzLYTeE6ZbFVlWJHm5u/Lzc3MuYvvzC
iZ/AkKnrKOj/YWpEUUDpCcuCYfWi/WyALkTuHFnh4MkbKyGTqRmXa3pFQhXdWmK3
CPVBB5ompRQlM3yRD/bRjPLeF6W6uq/JcYU/SxQp26j+alS8qbjnLb5Sd9FTBcjj
QALztqoWH6A4P9zFuo/hnfISA9PjCdasSE5NAcSNvgrP/uQcAlYH30LX6BTVHnZ+
flsmXrEjL9ajq99LSwUfuFgePtXWcnpLmZdE4NKB7yXosJIVSd+va94wub9tFySO
28ynzZZcoR+H2jJXrfkcse9TWpEtgIT7D+4ZiUqL1o4AJamnxdbKwsKnrlpn/EDJ
nwFrbjsI/gFI2Xtkfxfh+wQjVai8i7YDsJYakXcZWyI8KfruFxZhgClg3Dtcd83o
k/7acriArsbNtxk1XWxdOSQJSl/fD7nwUQvyj3G8eMzZvgOqgnu5J9RelmOHA4P+
bGU2S3hgZjWwzNPfmSn8/yTIQAX0KSstUpx89bV8fSVKeo57mG4LSzyBwiCQIbbD
HgFRTsLo4xWeFBeVAIh/4YjonsHfiQ7Dtrp4i2Gka3RZh28VO5HjCKj8NePIaEOw
57Aqk9E27EWGVw7eJDGv78xfUFamWs0Jc5LCsD7hiO7erhj3IvG9OzgpOPNrTE3F
dYrnI8Zzuf/n9EI2vb4Jiy0enQ6XShxSDMCg75KJOXzQpmwMb/Yb73UUN1T2c2PV
UyC3hWzl0Ekm+3+OqEZpgp+VzEYVajcnV00eayNbvIC6/K4WgQNJiw3Uby+pK38F
8DFH94QQBCSMYbok/WZ2DlnA0RD45dxkdjgZY3OdO0dmlADnNJhL+MpaWQrnQzSR
rBd8TS/QpKiBpqNRsE5L2rXBN6RJduaimcwqDNElo/XsBXaSpBsWDbjD2IWmtpu5
A3MHEJsMAlEFpA3Raaqbf3nGOmSKeNr14taHLmyRt8BlEurHv5i86ahlyYLcrPLU
O8QkSMFmty1y4aeOk4bw+SMx9jg9hM+3TFSsX+5BqQeVRCGj41lolF0mLMwrv/Nv
6vz/2L8Ze3bXYvxpmqDVfIBnSOQ94Dz4c3xI0oZaxTqFYL2qwp1yp+HYgHta2heK
VZm6rjWiFKDD8KrSYO5Nj3FivZvUw/0iDHWLVZtIcc3yxeABRCCDBvb8azxXjITp
DZAx+kiuYOzCKLpAYShmqHQDlNLI0H5xzRNteKgMgSSy2Bvqioz76+KmAQKLmTkq
Mjyr11NY0ZT8ZwBqnRoym28fq7ROn4glUSskuXXfmrPKpTUCzrrqBMQaHWsoXKAw
Wm5ASuKGY79QWJUHzINWN5wSQwLqLYFnfMm14M9cv0eRoHWM7bN/8zD++e+AXfEy
QScW42qjtStjnpawBb4Qit79Bkxxxd8hAIgp/4+v5wdlDk1EUm/rqqmLoj5AvxrA
IhLqSHKvGFKB2pYXA8eYcygrJoeerCAxAnfvFCPL6GPxLhXmggL6f0aNabZtPOFH
nbnRd9AF9G2fnqQu0/hhqMs9KANfM0Uw95P4OZqa1lmliTMH2OKDFBV+o7ZK6rV2
e8F3ZYtr23EpfiH6HlVfmNhwvTdj0fB1UleMVLyIpo4zi2kH0E4OqqUkasN2zFgy
u9346RVAVRGZudBskRn8433V7BUEdvMsFYtY9OyqkskdHVUlxq8Xmk7kdbYVyM15
cTx9T4UaU9Td0EkVE0rLZayD4ibn9lbzGqPvYAHNtK5i9wDKL2vJtEXDFHSyH1CO
m9JLfipztDzdBv0dUBMbrHTOxD6i/QI5KjCaa7sUt5gIrSVoMXBOCxlHwdjIXsdT
d9+K26b870MgPRlkB7jaFSrD3gGEt/qLhUG7q3iLHYXdaNNPJVYdId9An8IK1JNW
eYxelBmJ2Q7h98/xTiM50p9Atve7E8rkYVxt0wv7tO1HCgSfpLnjzK4wop4qUgGD
IADouIeBte9zHZihSjuXmGDYoDFeW/2ybZuBsJlNRU3tiXqEi5SK2cstG+MAzHAd
a/QPOMzhq7urO8Pcyjbq4nlMlqEVEXX+gez4AWv3+pz1woR09hlu/8/QPn7ypSPP
GztTN41PWegZIIqA24Hs+VCpQot9aKdt9bbR7CtvWpIRWUVlX4pIkb1SklEftc6/
g9uPbJVMHbqFV1c94SdANkY1mq1gaEWmu6DcFV/rycG0XTN3MNi9+Snv8id6MJ9x
5+M6UajvhZK/z44SflgPH9O+2qvwlXe5A4y5oROFcxPGAy76hI4b8v/ELVo9YW73
OCH/j6YsrttVP2VSL7T2UzsBVXXpaks3gw+E8qv4qOoMHlOWc+b+5hel91NQuIRi
F6EKwDCl0Iba1kYt4bQ8h6h21xAdT4Z7QuAdbgqgn8g+/MooXqoRa+FBCdrZUF3F
Tv4cVbAp7ATlZ5p4dptkkwYekc5WvQCmM+q29UsWXhoPraSrJebyc5/GgxZjQU/S
xqfVJxYrE0cJD0cIPH5o3f7TEQiX40sSD9m/5SwGYTOpVeEk8nB54Pn6fuR46psC
M8zaihNre/vqsZK759oYNgkApqUkhgs0j2r5r6892pSKoh/Nd5JVS6H7xkez5sey
8FfX/s1FaTzDBFHFVdmvhVMvMX647wK5v5SUDL2hvpSYa/iP8jjRSktLH+1bNvfR
/C3pvBwhrOJkaMKtFoDlxs60bqMZwDlzU26neB12RsId+TZmz6wdzMkUEvmat2td
iyTAud968TP88iotaKQzehSmu67wvzCzqh4sDWT9jK6SIH2jVpOL5Oly6hsI6Ez8
aqyN0NZo2uZdqWaqmbb6QXFr7FCcDXbvJIInQoS2ohZTnAaOzpHnCiQZ4VWy8eAj
mJiDuMMF3UbAd0HsqrbKCb7A3bpErG5s+7wNNJY7/RSrUnoN6QziyKTRGDSQl/Uc
23JG3yXU1wd3CJIbGJKda/QDU7CvQseoF50+hf+YcBqNQaD23wnbSGZ7Okmt32wy
WDZRj035OgJ8S2zsfhRoiOuzsD41DjdyZ/db2aI68b7K4msLmSRCXm0iYmgr4Rgr
jHsLjvOYmC63LcInzuf+mAxoMRbgLumy3twG5oKj9WGXpYL+uxR32jNEByu1HrW0
96aqpkdUzXwnpvbnAYUOUWDF4ExuW3fTmVcoXBbRroxEspJT9s9SNW5+s2FZAAeZ
Q+zbc5SAWSRG7TXOJ4H+htTPAjPVZ/+QX/IoR0zvsFj67xF/IQtVcycNVFEK0kwr
e9gKZvcTjdwQOdGpdWZaVFy4WNkqaSuKQG5eEZODWy2XGaTNDoyiCkzHDDLgvwNw
PwD2nYY+Q/IkfoDqV4nNI6hJx5LdlbAG8Sl+0QHrHJa+Y3OzKVp1XoibzZ7fD7Hy
HoItEJfuwnd+PwmGkFe0LGC2CyN+xBGea33Di39CYlYAMpK/UPXth75buzBVHGgF
n6TBaZqawYOKbsQy8LXMzHbshrBz/YuF9yWoXuG2s9EokmBH/Caged3U1yPhQ4Mx
jsIieRH2dwDmfRiAsj4OXfYYDz2whq58Hx/D6ZcLIJNhkskDZoB8cUJAu45pUyDu
oMIbzndcDUwFCflETHQorf+yqV7jzl5ycslK0NMCDHUSwY+C5XpSJHnEKEwBHJDs
uyzdbPDM9uut2MdUoXi7hRwao2nYRxd9RFRcCEZdscXhZADwHCoAuDPvg9Cq7CL4
o4lUWfDqZ+tlEZgO/hxuB6fFgkmINFl25suzUNV2ObOoTJb9izaBRheSgvpvUJI6
WPlFs5obcOdm7eMUn/QdrFlqKr0InVgw4W0YrUHb5qScG4iMQg6iX19ep0ZjjgZw
ee7sJUSmUj96HVdzq3e5yxZMCMOeYTz5GuO4MM5Z/lZtolJ8Z27yn/HJ19KtHr1m
smiQKbar/k9ep0esE9KXJgCZ2LgWR6O2FOHu3eR2Ee+K/X3LguVoXQ4+KbR/6VKh
FFWUtG5f7bT5NH+3NqTzJ6k1ZHHxsHvD8sod8EqdgRsumzBLUuinrWUI3DX12QcU
PRJlVKSopvPyE379gulJJsiLZdFqlYweC/UV0X04rm2DvjWbTB9iQXmmwpf6yYwd
tUdb1AytAhngswAz2XFXA0XSlqU57GDpbOBLjm1goWwkNEywyVja46yo4I62IOp5
sqao0G62rLWDS2hIUOhhEhWZm8aQH+jLtLcRjtLgneoBM8SNIaxfq+lDg7bwnu9J
6mmtEkczrGeVyzYEW1v4hKF5TPRXvtRoOB7fS5ZFncn2e+baOHND3weDzW5sEjUB
rLWC8hkVdEv5YTCKcAegS+YBDL14UZHuZQVi03rejJyMEqvbwzVedj4QETGuV+9t
dYLKzKdTxkYmUDS14wyID5INXQiRbNrKrj/w4Vfiteg3pPFg+HRHJfT+c5bU9RJR
YXzEVpD5xwJTAKHohtBQdmYJQo9Vtn1xmRt2z6En08lFlQBG5K9AGK25muHK2KY9
dn6Ial6xfOoCJF7NC+65vExakQawyoEMYI8+3vpmqqAfZYYPgOWL3TFDCFmIDu1i
SA9f8cxqdglNp0IHFvb7dYADg5EZBQqvBZaeEUWgbTC3x4NCt+RPltQX0mNrmUZ5
BpC1skXfOs9S3jyOYJl19+kDQjB81wgJfvQHwdZ3ZxrlG7qP2fevG9UbUc5HHbkZ
3l0ODSbIQV7wPohDTXdKpnh39dgYQ1y5kB1PYbHMwVAsD4D/gSlnrE5KhZMSKoxI
7iFh1BJCGOFoJeslRl9cLyR6WaOFqmvnPlwBFQL5pxYRpqMqFiDR6PcHsK07jVul
G0uSqhyf2YgI9JPlPyPy0kbhhfb8vdSdlxJZuoVasBmQP1pOMfETKNxHNP1XvZrE
/DIZzxWRI1f1DtGJ3ZQ49Ofs1Y0p7RirCSlXgmdt4MeQWDapZqB6SJE27MWbg2vv
gyEH6xKb4F8zWaBUiV39WVBSEy/6jQHTCpm7KXrMA/JdtRuhxLuV+bQYB4P//Dta
yyy7JXfElIsEM/F6WI2hYMEhfw7uYKdgtkvrxQztw+dGcofS7uyKA3uTq5KsG+Is
9fQNAyBWDkxZ7wn3b9zgdOXfJG5uvaT7TLyi1+1GuzQ+TFP9wSESnoreNpUmxFD0
hcZG4fPewGY20+AlzJf+MmGxTIZhCTDyP2fBFrGBR5X1lHeEle8+fl/AaDBhNvd1
jgPoE385FrVqfkWEEQnas91EmkC1ey4l2dhBNtT/1je534BSM/H2YYPF7tgfrjn0
UKLYjx/GDk1xnfqrOaQJBJgIG8b8F4uUHRHQOmIrqG+xLVtOvdM2Jx2w63K+XODq
HSaYcUbWTlR6bRrQ3cPLyNOo8aUUrn0iJOrMaFnTLJue2bT+/T2sjveOQ2fjmeB9
LJ5mMI+D5KbKKZ7tw15156Lygy9NcQ9D6uk02VY9Uv3OfiS2Xg1kqnroQ09brLHC
BenhkUZOw3Ni2bBuOZz5/JoZoL+9icOWKMcBt6T/kbr6aI7fMyNqUcZ/Btmz66H/
OTkMeexjXqQSGGin1eGXErhchteepCLSzKOucVXU3R67h/V/qow1+0BGSRzOVuZb
CqVPAWpn/p/KT+dVoGHy3zaaUV+2qFn3igibdCAZMdl/zuan1ZTak/UY7p6DbIZz
At3GcWCvIOR74Kh1zHTsaH0NEGEkfugltIIBiFGHWSJFh27aFpLx0UeBSkO56Vva
J9HW1ly51gf6N2PhnooWOUiB8SpcZ8wDlgww9QJc6ADpKvkCIMkro97KBIX5IbBS
sn0d1z0iOBvfrWoOTHNx01ZOmHfxQH/nn99jG543GiyGtdmysNvQuJwKLfFZGtz+
8qYq3rBESJb+MvDL3WRsszdlv3LBGtCKScuYJPqlBgQMvOj9Guiv1wdkMWdr1afI
2gbkr8qeluOLY95mcMotLUSNBiHCphY4WQOoDbpmYJd+8l00PYGGVieiAirpTzxZ
ZmYTdL21dBCPrroEdg+G0EFDaZeDSjpPVwLxn2f12ZjuTm/t6q7SVGZ2GG/vapBw
8SzptrZqeL/mFxmZQxbPFv6OZgWDwa3Yw9stdw4r+HruOT9FB8ZQrfxKIi7TYQMT
AmNv/H1QBON+7COKQ4G+07vxUl98cwq+L75brirzdW8lw5zXCBUUtaMIGSVdOBLI
LTOyXam86n5YLnm3NYOkZMBifNNIhCQyl2XYVE+A4GTKLTprxh0Ty+LBW7IgrwKA
HbDTXz476Ka79iQnE4fXxcATgW2xPhsGjCtyYREe4brJqRHG8M0QzoXapsvNIt8a
V5d7mBV6bpcIWDr6cEk6CtSpnmuYAK3bneI+3tJ8khGznrs4JNb6rxWHznXSL2Ud
kdv9MqO/bmlLQPzFMRAH92N6FE9FqJQSNYrJLvtPHfsF39X6CFfZEGYyWUr2uuJR
biSqsLlsNZa/LTab56xLcKsU/FxYM28Yg2HGzYqj9m8aiCJISHw8SZLgr2d33/GG
wseyzHQcDXlFDbBaeuIMwMn/0VR5ynSV8DhvWhl2mY79UqpFNCFnjHEqna6Tz482
uhUjvhbn/+mo5Nh5Z4JO3PkvALvZOo9/KFPC+nyxaE04b8RlEUkjowoagowEGgCj
EkdsdHIsL33FaqhM137A3clN+U+JTnqzP8EujqYdJdZzRxHX27uQesurtZl9KMwq
r0P1RBoWeCvo1dnBYb6jr9QZ1A8WaftWs7Z6nzrneWsSNIYD1OUmPVxvFqzOXrrS
pLpbTwu+mkgBsVMp9aJpFu5qUqzvY3pFGq3gXX/AJWAmAZ1FrVkfqJPrxBs40j7p
YpXJ3DuXiOrwpPhOVPxoMWlOfzJ/Z/m7ztFMwYpKK8yvagtzwDvOgFCNejUDtYft
FSxWwLvMdKg1RYAfbG6MJ6YbLzyeNkdPHfMrQKPPKOQu/IppfU4joEgHSX+3Uoda
veCr7HiAwqLwM1gMfxbAb7ha9gzxwfc5zhomtHD2O33D8hembq3YinhJU6I2XU+A
gCGppICt9zErqzm91++rd99zZg2mwJCZQMEC8ctw/3xMfmoGyItudCT6Vu5sWD1l
dcgyrbNLXTX1GN1qLEGSHEQnOSMZZkhd16tI7B/hLw2tpCpS1Zea6QVFJmOy8Q+w
GdfaIUC5Ae/3OjnmFWnN5MMRWCLkkySlAIBFdkoKnerevrw6MwxxZDWH4pfaH+6g
Af8qq4k+NT5jfRbUPpN4xr/0Cuok2rwXqKaL7ELrV3mPGy5FDW8qsadukhQqmfW9
vQGS5Zwqe42vVTT5PTYLb4ZeMS+QKO3C+FDGuKios4GmkEHFYn999k7oIvjPpYOa
UpIxXvyckSby6Z9Z2wuvB0eJGHHnzAy77+OllXsnigyU9Pu3cRzDzLlOrLrjQPG6
x2pRqqwv6KXYpW2IvK4IzrKlgSjmf24hp59RceyvLsFw1bxSxALYmNiTrVFtKawq
fNfPoyP9Jk2IDV+DLJCZwKn57pyu8ms/O8VrMg9lualsleyx/gdCuZIqz8wFvbdQ
mX97EtNWACrYFFbdM4BbTNXV0dPYPrElFfpvWKH39sennagQQwkme0eWGivdoRkz
IMo2C1HZjWQU76xPwu+mvCBrIJ7GPYRRKJ5+3xdrb8zonviMaQy/YNih3GJjNWx7
BSKg47Gv1K4C3wOUS/Ebx3GTeKqt7B0fg2kJKhW7aF6JAj8gKjJ4SSTXJE1UpUuZ
sP0WIEz2xT/yvxrO6xY7IdTOcECzu+oQdXiAStk/L/Zw+5JbzdcA0cZRlUSyl1wX
8wToCc/rCdTMa6niBc1oMbi679acwoN9SWYGTJmSKTGhz0K5saE1Xwn7abrEWUcO
EOnjTUDORmqkZvxIQQcpFGDKinoiJ4NTuIHbozvoJbRhW0YCS8hIGr65XDkkHMxy
HSUWt9uP74XPDhmZ/Gp2qvHqkJHtvf8eFht837nvSyITouP5nAt6nTCs5+K5d+V8
xPkRR5K1jUTse1jgL6YOlfe003hjUBRdGYSopuCjgC8cY8uGkH4mv9Jyf+wcUuav
G0zWw6uJKR5p+1sDAgFD1o1UC0zvfp8GcHMlj9PIl9h8VPdxDYy4I69uheJnGPjR
zocEOBZBJ+mKWBdrxJpy/M5UPWktog+SuiwWdmDZhOCDMWP/DXCLRHM82tTqxlCw
ygju6t7JxnO3mzsejWnyhBZHpUOa81M/jOTZ3JBLMDZxsxCcMDvptm8uy94lnOrY
UxAR6kYrF/f0UKcrWt2ffGVWlHsFTY5WtMO3AI8WYC2OBfFerW3WQNtZ+ly3ANwx
Rk6XJLrsgjrm7MdTC8XNv1WwOxwBjVpMOC7dIL22lvjKMMT2U7TmxktWassiq5AX
F3KcWGvhNLTW2IK+d0PxXrI46DOJn0FrDmNORHL6yXrThdtSReqbDSzCT2LSn4f+
aUTtXCQwEcCwuO7XGCj1kW0JuWPoWG0U40wTCHECVogw5/Ow4pOWKtIiV1Sy+/BG
ZvttMg1Uf5L81BX7hN0NwHfIBbZXsq/uWs/kVcehN6rz9gWKl3M8Wn2Pb/t4MCWZ
WkaKG5JjGHRAIQnbR/ktn5BpUMbP9EQvGB5M2gmT66bAJ17BLLqy45HR+5bSVmHK
EbDFM5AIZJKqcvjLLUG56osKWmKQK2sT8fr3uBUYU/MvVEKm0suMSAR43b1bMSrG
kjk8LoosuRK7VomkIesurMSXZg89T5WcFhK1Kfyx7h3HRfyfoZaV7sUOOCVBE4Cl
Or7Qzyoq4LOxeBB46Ijph/tWYS723VA9uHgCseoJ4NGDIlKwjNvd38UkUY6iVR0u
7HpKe+Jysi3te9r+khH37vesqqUOi7ibeo0+UuhP350FspUIp0ABFranurOU+27G
1GkYVkzW2k6m/UZgZFzG1SrQtvMZrLLLyJr4UW4FJ/xFwqfjj4LXckU0AX7v33iH
RvmkdRzGteM+ri7QwlLiAJsO1hxTgAbe8iDK/qjf/tfWhgOY66pAiDWsKpw5Zy2v
fgf/CJQf9pIEVNTD3gNweiBuBhdXHnxBbBdFD4j47VFa+KsJUgGi6+iZQ4Fd3AA7
zHFcwlOvfogvxGDHKawbfFSOZaXcF5N7dEj1Im+vfa8hlim21Pt6vKbGM0ZY0Q+p
dsaUsgk4XPX91C7iv4RHnLygFXkNgvmsJnNMOmH5f2CxPBUNXTxgEmEHUPEE7Oka
hm9geLYHQzrQqgTBfM9iTQ5uUo4rob10DBe3UI1pD0qZNaf9g1X/UK3XbU4ktFqO
kXmNKmtFbzmh1m9t8xjrx1SOwwFNryNZ9ZN8m/8+zpO3RgiA7CAQvkYqDa8dQqtO
ro8SLfRgyht59z7ODIRp1qDLfXo03BJdoZ/Y7+yvyIsFZVyxUaGFgECDXMVWIYLH
Ik0SWrv6PwraYo10LP9oxcivEvwmRCbYXjqnFEf5CcMpJS3tURR90H2lEJ4AlpC/
6NHldzRZB/U/kucyi+XiOUoJIJ+yUYkrOvtu884XEwmOPGOfUjtzwYDS/2pC82f5
To8yLzgJHJZOnDoi+7XqsGIroxGZ9Obv+516hmv2eckYAsjSJjkqnCtLw3ixJrzD
N5Dqxd5Bn+XdCv78LyxsfIwU+nluxqCtT4CQ5DznfxMXAq2kFped0hzxlRrrtQz7
xS/vXv7erahDjdi9BQqphYmzZntCE39HQK8k8yslCSK3yKmtC3iCDf92cqXIJcQ7
xtsi4uV1rQxfvke7XOdiVyuJlIC8nW/JlVSBjBQ7vtzrHnNw6k7Ii6qqlgxPGoc0
c+hh1A08unFrWctrx0+ylXnjHEcyKnXHgSUOu6Fp0E9gj3AL0Ig/Nm07lEl/UVlX
K3gAqBse4VVEt3hfqN5caiVQMoqVrwpp9Wfi6Doy24w2WOf6g2jTY8id094LOwmC
PyZbFW9S1iE37L11tQ03yfv3AbeldSjECdTGgE4Mnlqo5jwNsLDGyYG0GIVLpXxs
AsTrFnomPvso5q8dcxABrxVElwCg7zz5+lOOacox9kB2+VkUeELY+TF5LLJvyUvA
uEMwkiv82AvxjX4JTM/Ek+K47Qb8ojHho6ASL0KQK3V+4sxG//Jgbj4s75HpAPwd
bkBYWr+JRZEyfHc+XDXz35dkEvuJDtyTqaIv26p5gaUa17lSBZumoQ8sSQRGomNV
ooaNCeJWHDRWO/LFj6+988mif2rm30PhADpz9iqdTZZqX7phxkKcA8wFE8D+Wclp
yRdY5tCK6rZ7kcSlSroyf0PMWYLBykxR164Od5FbCjFmx5rMR8AgeDEylIRuMv9m
dq5W/sj12jOgbkVuilpHz+OZF2gLEwaqw0V3ZOI2h5sDkSEmDExVHSDTDqZWVVTJ
3Sh2oX6w6/TsszOXWgkEWD9yoMiEHpXODO1BrELe9qYPjX4NoRrSXmZVd0ycdXqp
Sq/0ykt+ye4scrEXlMpkBuZTwGjU8B764+x1uc3jUYSVVpg6Ko2tR33P6hRgnXOW
3edXBk1aBioAW5ZDboawi/m98L9v+O9wWV867LFj2d5vTuAI3yu1qWpcQrshH2zJ
kmyCpHiBWQMConsGpW4SvwSlwY4bqnREltkPSOgW1/gvhVjlPaH0OvJz/uPVoxVG
e0KaNe317nJcAUllWoshbB0Evrg9pPRHORoRgr52hvyFqcQPJl3BdDw/7aFCROO9
JCmSLH8LIV5HhM/1p/O5BigeZgoGOoxUGlG9dJLuLCpvSPg3vF1ZSN2kxlQ2/dXY
Nw4lXGsYm1lVtL/OtGttYPaTN+WnrwmQl7OMkB428zT8QUVVkzgjvfgdUg4NrGiN
msLR/jD5/BQnc45Ht7sbj3NB3jvkULfoWqLV6VqIB3Ykp8M28xOali7s9CCu5+IC
QG2po5YvF+abosBUYimUNDVGC8dXeAFSaAY6t3DYmHNHzk/CfrtFq7ku36OnnRoe
v59uhSS5+EdmCcP/1QpUn1/jtwN97XYJz/Nt4/7lIoHWCiPBa4SXy0Il70Ux34J+
CclkR3/I+F0lrUCSc2ANijaZczDLyVeFFcO4dABBSQo3suLeGSsbryiGJhf63yz8
UhmTneeRpzuKbVYYg3m0CcHZ4TzvsFcpeunFtZTuBgrlYR/6dBxLYtCBeYCgN6GF
NZTT4Mm4tDlNKND0uFCMPue6xg8faQODaSAD5KsHntIxZGXKaLXGFXsw+TqO42H0
vtnrzFVnB4WRIidTL8tRqz5icrOTXn3tyUDxu0ICQ+arPVIdArncwVpUJ2aZmMor
KD3cWReISw/RJ3/xifXf97+st9ZCB9MBIRoTmw0BfQOClIRX2X3jNTlyvZR3XXIS
7wlahLfZ7nw3n4Ls6uXNtpkBGIE9XFFITbuCKXOEW59WKjhGTYyY0saeC2OeQkj9
+hEZaYUMlCl5fJ7YwthvwpnkyYXMfXJXzET8YqVvHSHzYNuHFpRouNv6a8n/RK40
SoJV5CLKX4d9TP0PQT6PKPNujTecsHV5XZrJBMwtJ90QXmZheASqdha9GL3KuGQS
HPzgbMtavlofNVXN9YUPpQLPmNg7GSde6R+6A0wwMn/awR+3gPQy0lRob837itWA
tiCFhEnZap1vxkCYrd4f51NXiDHaOmoZomBY3AYDhmUyIMvS0U3Dp9PG+cX3bu1K
GnA3hCSwgrWiWlhD4z0riuGgasrtFGRsQOPJ342KRc72Ktithl9MpP6aBxQuo+/Y
45KqCNCVVSSRNhSwMYaxSqwlx4oNxVQs+e075i3JKj9DgoS3YXJM8cAGqcMGIC8q
Y2ACQYfKE/iRneh4gz2rZU9pFjAgAOC5jg54lUJsZd4pMaLyCTtqLl1QJH6l6QMq
ptukvavLLTvfdBRskt45oHSxVP3/72MatlegAOVQgCb6WQ/zk0dE0kY8ktoTlRoP
DD5s7GCzem/LzvwYA9JVUzEcaHGkaHN3vBV9iXZKQKrPl0OX250eQNfRpsx6k0K2
aiM8hbd+FZMs70BCn59x7hT4A2bzM1W6w/qVaTfFx4/fk0Q49K0XBtE2/3PZRDnr
UIvvuSjd7NfLPnBm4JNaEFH8eAbGGmFtBPbuKNGyJl+pzVqDvoxEKeKVaN91uokg
ty7irtco5c624RUe1IHOLUq0+fOIPAeMrOJ10y/aFQtWIjM35gXOzfvRTRGyYahx
CfGUF7N4jFO4aJAUjovjowI2iq4ajpD150GSxRAqtqLrtwOPtE908YucJ/0Rm5EM
XiKjrVwbBrG44+rT6cbIvCGU7N79XZiOuFT/k48Qaz23C/MEcAYccfYXbMOhrR5p
qz1zE+ZtgmPw0snZOA11dhK2BM6jKAXxhomccUJvTPOn1x71PxO5LXP3hxvemk0m
G6VCrnydNd7GDykZaiO2SGu2xgbHoj0rkARO8vhnvf0CQruI46TgpvNBv5sGZjNu
EfIYPCX73Hrl0kY8xBXmjVb+7poBi44UKRpTD3SjAYLG86B+eN5NLc/w/SEYeNW1
iVsdsoFn/ZuLJFKRQrI+dAfXtguEgQZK24nyDB5wc/FaioE8k+38ZMCJEyNhb5WA
Hlb/gAnxHIgRXE3ejtC9LfKQ8D6XEljheeztPlqfTfyrkQYabZ9UWEECZLPl5SHH
nxt7C9eyvu3H6Ck6jkwMN9LQekGEyd4RVandg0PJV3umIi5TVliKbxoRbB7TOrsC
emTpg0bAzpxUkaj83w3xSQLrZP2FCVHXCbxCjBdIB+55wWCmcGDbODIzf++Zq4w2
RD+cKLpRJbYeZISFLN0DQteEQSKJ3qMYBZy7LYMzW3okQqR9ojxY7+wuW84JxEoU
GKDVDk++22ORgqKbIxRa80aPkd+suTNSQpjLFEgS49IbyaNdvpObzFRAF0ZJ/A9w
ayg9MrZnvGBtWqEj/PlrwrSXNxgd+k9/Q5g2T4KW4nF+nmmvncDjhhliMIYk30sB
XuRINUsOL64eH/XGf8DcEAZZU04HRLNoIv/JDNP5bKWl86dvqi9ZFFnjDMU6ehkS
H7zG/bME5oJsibn6uJsUuf4K4haa6ppsaLbiiRSs/X2Vo2i3maXeQy5paW7Jau7N
PaRmz2vyvsCosy6khd2tW0BngiIanE2qn7l7RsF454xOVn7bZ6lK5sPlCYwrjUhd
oosQcJ3A+CSN7oXjEEDsZ8Gj3leePq0oMD6aZo+pdQ1B4XI7Ieyk0wSOvGTbSWyS
L3e9kleKYmHHKP4VFkg/kTxkYFnmG02v+gWgcxtGAgBhgtSHzQw+/r0p2hnLAHej
9L9Q8RUAlCeD8uCiVXnW54QYPD+iXEOuCBaqXYrrbivlxLeNye6+IVIKltikKrmE
J+jO3XuOtPbQmESmaZx3z6gWleD8l0qhCYYEWBU+PQ6SPBIhSUTCiLu+uKaBPXUL
jON/bfPHH97zK/cXrZm4b+WdE2cRttQLRFQzCgwK26qli33snWB24ACELbTuMrA5
cvu1e3xhf2fbGuVnvp7lmdIIgRXIcnPscqzQJwiNAGO7V/VGt4R0u9VhaT/GeYwa
5KpMxGFKCmo6YdV/AlqFjdl21bkeO/F9bFPg7Za8Vzwg2shIkBvvsbHj2pA/BdfD
gi8kB9/YJ8uIxZu9L7NMsij1GRpG4BcJmo40eOQahTKbjAhy/BYEk5p4zvNjVJvW
ROcLjj+O3lmRpVgeOgxU7dOTQ3eopJj4PfxeRX09ygd7WmD9Z+sUJE7AEcdYP01S
y6/6ocMhS8MDVNulSEmF2C1Or1Peun9JM9Vmg9oEpaPK/5f4byZgosBL/AmVpNxo
Y/Qdt2xTpdf7gHRl6GODkZDHHG8MivkGQmk4+AVqbuaigbYTGWlJkiHZ4p7Uj/yY
UFDIKVLFbCPNtuiopEk+Y+C3iQWE7cmyna36WGVkP+JymMwVAFh39XSXBsFKiYhV
Qpy4Pd6B80YI8TpptyR5GXtftI+BL7DJ516MZDp6nkSXtO2XN9Gkz8W3+4sm1/DX
29TOkbu1Pwtg+oX/n/PFL0cuc0uPQrdjFyjfx0a3S5vTqQqa5CrP9aEH/R/Blox9
+MBNYBKSzH6x9p1seclU/sMf3uMsrLSp2iiAHWtM1nOwDQc8L0Snt+mILqm9GXjt
BiAotcgybHxLWyPJZW1rlfFdt+s7SukERgGBovCkaGVjUSED2cMzMdTdD6aCkVP5
eHQX36VGhXXf8YP6KjbQph7VNJratklIFJz/Zdcq8sPCueUPmUftY8aSno0o7CNR
B/6zdf+RzqLQ+oSHDyKSNXPOcjMRo5/8XF4vNlt+itruyLYUoUDf4SaO7o2VhZiq
a32wWy+NRfpIOdxACXlY8R2qvTfMXyH55vUdseX5c+QhEpF+Bm35uj8qTjrHTDpW
3+hfhgHk4YFeMZTpWTBsfc5k9HP6joG0D9F/dAWYi3cIcsSEdK4eBK7BoM+fZ9uL
FBE0IsQnFWsRouznopwjwnKEc6XNL9I7k8YNT0ijN5+SvSJ1J/Z8zEcckg/zPuKm
3sczAlbcb8dken6QI7VU8yWTEkDko24yiwi7+vIweISqcj+BVZ1Y4fAxPDEwVsnZ
FLHl6mfKB2vWR/ui/qd4aAYPk0srbuhSzjDQ6jq/LvBFWpAvEWBAIASb0/YE3M6h
XaVNghakQzmd+yGpLRk2MrOZq5K0YA3f408HrnFuadIMYa2BT5lVd/jjCMXa6CVU
OgQrYidzdedZqaUWO3Pk6xe1NIRCDjWiJWfrI1mRTqK/zfX3brQSaW6JgMMv8ISa
JVqn5iuAUV1zPqiS7zdBO8P4v2orIVmteQNSGkt7Ooa7LGWyA8yNmvRFbbaCLBQz
sCWEv7s/ikVY7MoI5iddAlVLxUHFnPGitw6OH9ueUCzeKnYbQ5VQ3qFKBSMme/fq
JOM0E3BUFBVgRe0LhGVV77nSmQCQ2kQ95l7lgefbCXHq5FUFEUCO0B9uSTDx0VKh
zfsa5NLOLapjkg2bERjxDBiCUhFNM5/R8Cyn5RG9Zvjety5/T8dD4BL+8PD0VmxJ
ojceFLH9IAeyNEANPNNlLrqisPgYwMJX5ZhDwF3c2+zEVthHHAlaigb11e2WlbXp
pMXVufPHN98+OYga2ltLxr9xOB9E87aTbpLLw//Yf46yCDPPFunY/RwGKBEiXUFB
RB6KBYgEE1ngYOzdy2AEPqRAo8L5MU5yItOwJHwimHzWjcwt61MKXTN02/XL3lk8
RHRj+6hD5y9P9jGQmu70lsF8qlgQRJAyGGfplKXFNRnO7h6wQ3vZ3/s2hMxAHE3r
0kbDWfV+gSeJ5cRq6mlJKvjmLTVXjlloqYqgvA2KadgEDQap4fesQg1fwzS4fVmn
j9UcDqgvRv4Mz3jfWdDfn/eRTU8zMyfhEBYr7OplNRPAGungldU/usPiZLycT/sB
3v/MLV3WxQONhoNcQwTc1D4lC861irYSQIasNY6obZu4bylp2OIB1rpE3i52VyhG
P5NBfI5+4H/pawfoXtY7Yof7uxGgmRrfYoxBSV7aptjn6m+gFbZqQcFk/baLyGOI
bTv1c0WOiKZgfOPQJaDN7ygwURtBnFjfbNTLLKPkcnQ9xVBcClHGbfYgu8wZmmf9
Tf4i+ppjNn4kP3lYZwEYaXx7/N0tFs0nNFvjc1KntCgAUgdOLbmSI3jK8Jld35SU
qQoekj7rNTXbnZMnPBkLQm6TJDl4NQTauU7AbxLHLqwzMza8HJTpmCY4Y8ipbdnb
8GyZ/jYsNoKtQboJUsAwOGqMq+FGh60r6UJQB65Xx6JjJOlkRKEWYjYDrfR+pJ/n
31d4GDWELSSfZdmMFEfKJ/80NI3+9J5/9jN/o2xrjvxr80bnVgIwB0QHQ3Au4M4K
D3whWhtFhiolRSFv/Eluna7Fn00erDlrcrUWn5FkugmdQ2tI7kXXIpA+b4iYTrpi
qozeR3/Jt/tT0/MUT4IpDOYd3xxszYgZg0ZZ/2u/134HSMVkzEvI9P6W2SXRYnQ3
d0nBnOhLr1DUF5GvWQVXvu4vW5b7zkIq0K5MJiVPJ+0DAVHtgLFeCEYJDs0QpAVK
Vbr8DZhVhGv+Hg1xD3kNMZ2rhAtiwMU5K/7fQvRUbQ9JS1nlKhBuwZjQmWTcJqw5
XZqwsVTDfE/tSMcY+7F4NXgra6teCoLjfy6g/MvFj0WpXzHJXYCWTt6cWIh0yT3B
nPwQdzdvPDZD5V0ZFWaqNZdrCDuW2DorEmC/Wwdn+KjUYPd73A7yYM8hv1R1JULb
dIe7LfjeH/yHp78yZPLfI6xn9sgqP6g+Hrly4buIrazYRnTMtLN0HmzsX5X/RDMC
3WkkHNNZUIjslTYjB96LzGxzxS6SnWddu8A+jbDcZkzbuut4wcWc0thW9V8Wemmh
lwoYOAYb0SnZjVMs8SG9GpvZIkweHAglJw5SJNu5tRx/hW/zHxMxIaGhmz73xPfC
6A3DbqIMisq1pz4fg70tOsrcxQC9gy8qAvetgpFHZt9hrOclEN5tJosAYC4qJvyu
RwXMbhBFBUq48OmEuUaTXS2EA8vstIEfd0ZjnJs5gpIDjPGfbSCl7SBy24ig+4uK
+ofcd1YLl/ztlThIMofRPr8pwxinHX/AAF2ftK7+/xJa3N3GHA3KdsCoNmsVVW23
qbhIyQc+/W+O2AhGzpCE0Actm+BxvcWb4wcaSghWSX7OJFQTwOVW1C7Hbv9FbZiU
7DZ0yUah/c3S5lcrw+jee1Njh86vYQXk9xl0i+yuS3jb8ptZ10oAAC7LSIORUVRG
/GFViLcyXDnadngxNMyImvQ30sPeCUpxncKjvdlQgcYCDcgxiF60VUqa+ivceapJ
OJ+23hQI/u+q2hq6PvKF0tOBkFGfRLBo6yCJwi1RwUFYPX/hSCc+piPWNOGsJ+2l
edxhRo8cBjs/qdNqGeZcVNO4HjYtpZJul9JQDrMTx8ap31TYAXidPrcZ9LDHHJOQ
LKcADpoBgMtFmEmw2FYfMl3Dlj5cxKEGfnW1UFu7UtzSjmToQb7hpYEWduX44J41
xVVzKGg6m7kyiyWczNLEtmupTeZfnLs4+RfOhFHarK5rN4OWRKFLwnYmQGOgRUBz
9yBb8wJxBO5hXZGXFkiS5w1lfRZAZLgASRAU3oYwDzYPYLZnvumL9yt4rnqfAkMn
mVkzlpGJMnxTu9cZO05XnAfTbjlMpmRNnRfcW4nuIhiJJutQnUxGB7l9RpmAqlAk
2h0EBpSr3BOnZX59tjG1kUHURZuooXWmqnfE2wGGxhXOYgbNZcEIE8mbNC4PCCv6
yKfnymvPeWeICC0OYjN9T6uzOahzfAPI/etr58uJNCkxXh9rl2nKPXu3pMY4LdHp
eDC/7SMMTYfDWnL73958+tb1ovDf81QgEIXxQhhui/kVlAnGy0J8UQk7cXmiIfK9
7K2t+CnvZdtHkAntDibxlX1sJPL+WIM22yxVnV1lSFGphMpKfU6SiSCt3O7JpDev
+3wcIbpmLIOnsO7yyz/jcMQadXBvP774ZJkx0V6e3YQXAZgRjfbPL4LYfkzBSn7N
p6sunibPSiLG8dG5YOf0i6QpJKgZNwodlrq7FG9hicOL0C/zbXqJ7wnS2A2Y52e+
oN0jtsWaoe9tZAjmEBMzjZ4J4m8AeA9LuofZmBQUCry3L3+iDtk5bvrwOuB2xDWP
I91+iAF8+Jnof+XjizbXfNlimH4MpNP8LGtaREokTPuLbg2nVjYqv6p6fPN7nEWZ
yTDDTJxRJdLQWb5H+ACQdtm+UwdGi95ldwESM1m2Rh9pRdyPsyAfeHFGhxalVMvN
juQZOJWsPbwapA3quP/j/hS0I7YT4ZTVzAns2/BPLdpRaF3Q9lJvBoFqfYbWlqQe
tNO/Pu6wdTgKzqy9O/HvujX13Jc24SQKDxYqLprkAWxbUBQgfBniKsx8bsagfoZv
nNa1SqYwPpyFm3xtxmixtu90v2REM+jRTvi6K9NnCaZ8dIhs5Uno55YUoLs+89XK
T+nMMnzTx6YT4h3vwuA+LDahCRa2U+LWSbgJd3nkbDLtIUUAl/GDkgsP/fL+P8QW
ZgBS5XpKkCUIsHbhwmzpsq+NahR3k+cVVY0+vD0CxiHCsABW5KKzLq92PCO/pn83
+VyxoqWhIUY0EIyE/Xv4KHD0iERNegvt3geO+5ZedF3Rd9ELczbNfSiuq5+iwjqC
T/D5dvWZy2gPbzWb0ybzNUc+82g30uyfL8Rj6r5KXUNZywaNfv2vUQEiuI+2lyTt
dVdfB+DYynuZpD5/0u8VLa+So1nurF52hF8rDliM/POxef3iGvnAAO0mKziAoCBR
bj5IKiq17F7IJ/bbFd5TiKwrI3CHct8F+X3AC4kL8hGomFQCmqAUQx+6XOpTBcAJ
1FZvWhMgzvm8w7/PSEZRApOzejoCX2RmmxTp8KqvJsi93ZVmwma0vb9LogWfUBNZ
PK5eWeECv4ouBOGETMK3mnzeWBTkiXuozXpmpnTyag10mzHPlhO8TTafsP1i9EBk
AsiQDF+09nHOkLW6BtbSthAM2g6EUwhsFrr7IdVmvjeHK4v27CJGxW96egDFn6WX
CzsqkcSkjyCg7PgbTpXxbKPsNg2lOIv3i0bw70lCn/5i3lGhC4UAhj0dAlNWlVoi
K0JtyeMIVGDVtuI34cKWHqp4J8/BmrXijvbORvFI9blOJnV5HUhETfv/3yoxmxIj
yxEusJbgelrLe+wWFPS857sEL+/9JBIFTKgK3ODqEuAyS7lGi85ePveNj2O6zfX2
XqBzl3Gcpcx2BjkU9Eq8IN5JE1oTRs6EfRbsA1u6kzAwKr7BydWPO54Q9EhKv3co
78iBLV/fzKznZizvUVxJpgyqeKnnN4jhCc0XzsPp5ihdzQd7v6PDgwOt+SiC3Mil
IpoQ3iqvmulQJjphcCVg5nVBD6mN317GNGPQDrg/bXcsCWR/MkaetAEEqLZ/r7ik
+x/L3GJ8qbM34QPrAfJyrMGbYD5vZs/wHOi+1XgBjJxZu5CVHNGFsMVjQ9P+UzSV
/vf2gR4HIjPcDLGoXLMpM3lxIq9DFuUcxHZEyclFJwpIlixz97iMVTgelcznU/CL
4/XZq3u7oAri3ncqJVHXvitfJhsfZw2Zz5aH2ib7Uh9aHJs2tB68J/NGb/G+uX+C
GrXg6qEEOdIRejVluZDBTj9O5ZtOYi4T6JRVG1/lsyMWE1h13CZ7f7Hgw+NltM0E
PBNvxNxq7ATX9PImLV8MIFqOq03+AnaJ+wrJ3k65F6nX7AbydzUegvmwsLatJtkd
udLZexB0Up7+q6LNoJMyy9lcC0b0JeqViRft2vybQDqZXdvtdsJjdAIBnEqnmVbg
75vSwyXdyWQTUEQQWtEwR8VZuDxs1Qehhu8nWPZbyrxlWUbEd8Vd3ICmhOQSqeTH
cXixs2IkdmFuQbxQL+mcDSJ1OntdyZ951s/Uhx/Pn27IU9bldMl9PtN4nOH4F5Yq
TepDbvfvhDs9jfDYmgIjoK7peXCbbmCsvIJAp0yKl/1/XbFFrKbwAxsK7RY+C3dJ
EQh4mUDZJT6sAkPzwDp5+3THaGFp0QyAteBbC8Xi0VdsbBfVYp8uoOxJD6NVgQ3V
LiOSDwLdC6h10FRIsRgBid0bs1eD6zWqLLa6pj1xkXE8n93rLFpHSA2gSgGrDqBa
S3kyg9FnlLD2W+8JZ4is2KtNOQRgLD3IOUaqF6lqE0aycMmccNxJBGYLZCnMgEFj
B1kExlum271ejzWhc/d8A9hfByYXry6HcQLi/efsDaugqlIqaFu/akjPPNKE7pMh
9e+7FqXJIl3Yp3D7ozIDPMILA+8oTkOX9w7etFCBWuDa38jBCmoqiV1i7KZuHy3D
gPbPRuIcTVMwg8MNZdROB4wd5z/aiRA2VkMgoj6uuslhMF2uOAvbNzMPPWc7Quox
QmiDnNvZMcDEcsZo5y8M7W3WkH8cBAhUTBxrULSx64eld5lkTvSwlEnqO9krOlGO
BEUoyNhx+cxZkFoH1jcDCwsof7vM3rBfs6mGsGNuIIkwysqTEpno7Fj0zYVS9slP
G173Bkt6q/sLeO5KhmPF+g6ncmGdPfp6vqGvdF1MynqB1QTUrW/MK3pWY9V7yq42
AVt+ejsXHGvJXIt0FFAIud/P4Un+NoCiyL2lDYswJUka/ktKIvuELBj2i7ZEJ5kB
tZYsQN8YRLAbPNfue/ePILByfI5X2owGlyflSMTQORrDixnWklE1JnYe57WzEqcN
wL85otpJvmrY/9NHUqwZ6nhidvbG8m+ZfPAxAk6oyWwntnqv5baxJNAd8MEH85Wh
wC33Pq3ayGmCCLXgtuq/+8kf4PnrDHP8hpu58ZQrIFu0xkbmbfk3/hgZ+EMMy+d0
1hy0rJYbJYwgpjwJplKvs2XUtr8i0PsxYPab1BLoG9HMr9jYw18fRXzB74RwKPMb
UYBQ0s1YI9VKh/+SvEwmt+uLQB47c3KxclMRR2gWpbJMvM0B92zFRj7dN+ruXtf2
/c0o6/KhxV297vTEZwn34hxFYLl5eQj035CMjShtl0Z6DrkOreAGjRlNvHBWHEAB
XKQWZR4+dJOddwOd2mrIM8FwVS3sjXJ8wi+RcS2VKArBF0kG0KiYfbalBcZBspbF
WBz4WXIxqCe3TBdkU7Pl7+Ih/dvlkaLyxIdMWZOTrB1XviIG2T+nta3t10Q5vzLe
9SmUsJMzJ2golBkND2L6QxufwGOEx8K19kbPELb3+L9IVHspvAACRxH5Y8b/vEh4
gM3LlDrVKNddPUOTJ6LNGsKvx0rsiItSEXauQpH3baH8B+uUUIsRDJ2n5rNrZGt2
pgbvbqb03KBJSb16WG2+K3Yd+G1UN3Nj3SVInJP7IooQI9o+Tj6z375+L3aMVosg
NYcwijNT84GhevlQ8Wm9IS0wdm72kqx+FqfEZNK1MM5oBtGte66gMiGHKzMTOTNE
FGUr3lGzgbivGI5EU177tNtiGBPHEjkc5XWEFqpy9eNb6TJ5tIdIk/HPmfyPUTR0
ETfrSgrCftK7kyK5L9qT5M9K7Z0fcRVSPnwdbcFA6ucDRk8m56vKRrlKvEeqrzrh
HCIAxJRJwIpnZrBUPw6c8YuH739weNQ9tko/55U/FHGFOvWW+vU17tknklucHM4o
+wp12b44A9qmSQKbmlGY/lhXAGtJcfdCyMdrNYPo3nld0dAUu6IlZxxP8gIK3PDD
Fs5+CZhO72hO361nnY1QqZSXcYdJBP7mxrFCIg8vl5Q6iWpn7aNl2/Ww4W+kjOfw
aRYZmf9KQpTXblD7p84uGRwUJePuciEeoqcWlINrWFKhgSxUyucP6RkJBboKXSKY
atmUOZqL8AE82EfgksYxJ0vr2KMyFWHwLoUjBnfq6DFJsnF4EI+qo00toY2oP8wC
WAkKexvmvdwNUbz9XjvDNKiHI2QgCukEb63s9CLemNQWrwbTreGUlhE1WlcvH5A/
GuVArgr5d6OwKuqYjhd+sC4NJ7sDNI7BN4OBclK88DGU1XnXh2tQv6hIvfbE2m5+
JoBIiK1pQ1dN6gMq9nRWcE5kC6u1Ei5MHJ4HtC5mwCC4JpNA+uSbqLvK028Pk4oF
VerMcdDyeqkpQ1T9Ctnw7S/4MIsX4Eo089lAvZAOm5Vo5SHr6JFa0I/2GGTztj3G
CIgVYS2n9hq3N33SKqTJ5PKbRdhYPl76WW0OVeRXzCIjGpMCboCTzQLrFI/FXap5
zR8pOzQk2pKLUXyjL8fJv7m+0VxJkQt+5wiGAmbnQQenAG5sNiFR4uW8looxZFpV
FAQlXX3c6qA05OsNjpxcNONPkanUb7NSmaK7To0/ln6DI1w0nXxCJUFzRqTmgnaW
1QA8kSbtqtX0MhQZ6KJ8Scg66Nojz1nkqdKXaGSnYIeJUZc58c6NCgLvfrHy1Q8K
bkVsMknA4xe74zhrVH5hWSlTZJBA6Knp4OpizY+XlTIuGXAXM3eU/K4dMDFf1fBQ
cbSqq/sydIympR6q/6FDUvusUM5ro9/RD817y2+adCRyRKlK4rRkN4q+6w7mgEZD
aWBsuKDmWfB0/vsl3lCZF+24EWX8nEkHmYxJ6qqrrziggREc/RqbpvEZA4d75cR8
u06cCDwT63Rgm+lxlPFhm1lTMt50Vijo81MFW+djQDNJQhH8RjY1AJq+bmHKeaY9
D1U82c0YeYWvhKV1XaCbt3l3xzYsUuo81jXxgNsfgjfmTyH5lhb/HymdA2jijhMW
j5HW8lMJPfOpq/0n5709YmkdhJTWLl/l83Llb23lcIBlr7QUGsEN4ACRGEYLLjTh
HFxj6hUZzHz6q6u3x/53X8XlEmP3DUXs+trsQVsaCOFmRbCfSF9ss8Gz0oEePTqo
qbw+cfx27iXvj/qnHt1Fruy5LwpKe9V1fre35OBgAb/rWdwSYaXCMtDwxSFSaGOY
kUyqGdDgiO7WbLM4wpl+5Vfe+GDCgQ3+/Z4GaaDogffgcLRfHNRBobc6GStgE615
RnyE6XbZx/RzIRC716Dhirw8Eob/hqkkV6sP0hkLSEe35lkdpW8c+Ir6hcMNwdl2
LzJ8NZ2U7M8KhEbML6XQLRnaLUVLzaLmBaLho8zbEUhrZ5EdRpYrn+4to8YHRksn
BiLu2XfDmZNc8LKjSdlYSNs+AqxJtOQNvOtY9iwF0sW3mSf/XFZ7thyiMBLmgvFt
WV0QTt5N6Pf9E7cI5G+lCem88N9ynlJgG/oqYGw8lnxSBHxQ9Swe9G73lwCAAysl
1lfdczziAOanvPD5Da+P4DrVL5rwoQQJMMkwL89lBCiXQyHM7gjYyRm6b3wqCDMj
oLdvDAqNlgNz4v9E3IrPQQbHSqwTFLFwnEmFOw7Y4N+2leZT/FIfJQlkKaZau07+
F5QRzUe2zf+4Bnho2/oIVVwLuy9SnwBDa9Kps0tIO8sVe0VR0sb3choAFPquQzE6
IIxh/he9+OxC6He5LPZTNv6LhEQt+hHTGQ12JXziHKKUsNUPZeMVC/O74MhkKPQ1
uENQqsMPcVxwOnLlcXQ+cS7yVHyLsZYELb1OB+39Z/kN8CcijTutPVjrsDRNM6cz
+TQYe5xjLVHA82V7iGZGX116OwcHDAXrSsxFQqWyl51DOkqb/ZkkPRXDKmd/8/9J
rTCDBZMt7DajJC6BAWErk/LQ2lkt1FMDgyJ7V+gUtmZaJGNSg8u+Oj8wpOreCG2R
xGUzf+MR+5qvV/e0ymDS6wj6AqnaBFMHHBXgys6l3Mh88Bqc75NAIMv4J7igQeNf
TCfdfwxlPDnLIZgOR3Hj3Pi1Y+2Ooaxeeb6Bqw+i6rKW0luVpHimTGjontqqGRx7
e0jQuIeTf/5TG777/N6pHLV3ngyTH8IBmh0n5F+NqYec6MMTEz4QUHP0mXOhfsFZ
mN2kZUebo9O26dFKmTFapjiYtihbbN3mNH7s7u1dtBsVzeWJGwfhv6w+OQMjni4n
6aFZzG0KEJF2+N6sIGPP4y4owmtJsX4s1L5EW22Cyax77wdYqy5xYw5VsSOef95N
JXQCe16RSOlH0WKCXKw/qZ+ctY3DU/dWcUAE1lcODC/PK4o5tTAmLUEIsJBmRVI/
I12D2Kn4dXq8Bsb+vHupe83AtIpN2bAptZasQP6mGyCMZepCsizpTxLROt8pmpGF
P/5qx0BM30W/ex+qRk4Y1pWNoBj4QeZbSPlAOrhAt+/3wakPFE0iHaWHHGgU+lFV
TDWxOL0Mm0A4+eg5fybmCBvp032Vp7RcZBqwTAd3+3iNfmcIx1EVt09Hdu2KyS3C
uUQMUIPtT0RuL4E6gTU8wceJW99wvshEgj0yD7L0sWbMtd9QD/nZWNfSKb+6TBvC
p8FOWZ5GaWqKPr94G8t7MgDZaiaA0BtU4h37LN1pI7TJ2k/GT93ASkm8Cs1+3Kkn
iZ098zytcMzZae1v9q7gJnoDF1XUDR+C7Rz8A0f4jGHisD/ASj3SdAK3i/0wNJZA
5rVstdchS6Jety1whpY2IHU5wK3BwANMhqEf7sShmpV2bY/9UoSN9uDhstFwWbw6
UnO4GWqGgNHp1v+xdN0f63AP+o7BRpxxKNWUGYn36g0KzmStFA1csylh3P4KXvmz
9zE0lAFLTWigdZAAhqwUsTF1fSbm0LkCl/qrGR6QJv8fxTsWqekmdi+y5ZIk/RaK
Nu8oArU+oRCwqMc6OBmZXFSoFxXGx6zvzYMukjrcVSqGVJoBD7nVyJxoIsJeoxUg
RFUi8HiliTJ22/LPis5RLDtubkvNxM2ObbN3TT2l+0VEp/ZNJvtGwKuw/TRdKr2Y
p20qo1+Np7WLTAOiYvcqSmJEn5hMBkdYwZsuzKIRHHpsN+uRTG0NwU1k1p2Cekhr
7CmWFc0+xRUti9ty4Nx00vKTV4KNcajzN/ymVEdHfBcYBTit+lVs1hj/PdtIJI5F
XzmM7Murd1km//AqP1w3ldXW2Te/XVavz+Tfcwxl+NLYdVP81S5diJtWQW/s+LC6
Bj6c7H6mC5GaCJsfXktLumWKfORBqdSVS0zI5zvDEkXW/juZCO/bn5dd6n6SHaDL
PRJw7c2oIxSu9g6hgP4g9xvqa6cBrkW4/L1BBLr00nup3TOwCGrPw192HvIIQRSQ
EUd5MTv49BRIYeB9ct2pTTFlQw8gSx19Mdd8YF5RD8p+WnaFi8lqE9ygJXnPJht4
Kaoc0ne1YT4nYJgG4RwYQRAH5sC+KC6A42GzxYrZmics5I8iZixsdo0IsklNUNyZ
RNsCVMpuLP9xEnnjyUuJ8JDTDsKvJAWWlmRNfttySvgiIt6f2M48qdIMi0BmJo7I
uw85ADgC/H2QhQT/gZ0dE641gxWhkSWM7XQLbwUIFUbe2VX9r3Iw84ogZlNc01b9
iL/3kFvkuhnXVJ/HFu34ShlepuPStHwwUTveNqMVoDhv9I3Hh90mxpPSHvvwkXDs
Mw6UHldGVjeTNhys2OlA6txmcJkYKducCSf5UBVknhJ7M5dpmLeUlYlhSfkenQJt
sZ+U4LDirOIWzRZS0OhWxxZPTbx+mWxK8hYB4D+h49qeW0U+vOlLLvYtgBm+9rSS
iShrkqgB64kO+5LPOwkwwWfTn7/H6v+OXnKRh4p2Lz3uBZcQuNxIMwtf66Y/ZSwV
qVNPRr/npcbrMiPmhtrPESLWohA5kU4XCQiVOIBisfYePz4DNZBCNatwpOm538HT
K0HOanyNIHz3RQD7al/yjSvxk79z9C/aDOhc9dlB1t07kl2802NUZLmAxXM7FaJB
eo/St9+SoKRcsBZvUjeNtXosl5KwrpYiESDH+STE6x2hZiD/OkGOrWOXi1jdTqS6
YQJUMva7ST0gYosbkzhJjTKOtf0znYcyXuGk4xr6AKr+0qK8DuKo5zpPrAejZ/eJ
G0AZabpKAlprBn9h0BKeKnrD6jpuCBWwRhyAR2cI1pOqIYbFQ7WxNIOlgzrayP+0
hFXSz0BWE+2ePE+/o+W2kRtGe+RfwLk8kEZB5gRpS1jAxLKXgf6UED1ajVfiuT10
1q8o9Z14+94god+eeHz11AgFimZXjEVcSubJ/f4+6fakXA2T5mbZNThwVSxS05hx
eGqyLop35L5mhSHM2mWRvPS4MMs/a8JKZzv/J2qH3kiBAfzQ3lLd9xeS5vYv42TP
CBNcY62VkHN0xNj87Pa/cgQz8JS31hoh9e9x2vEcdUowwabSyCORXbniSLuhrAdZ
i2pCmyKNx9/rWAM7tEifl0lSv1WycFpPyE9ml+4m5oluCo0j6iFUBw9rLe+G12Mn
A6VyWIWTO3Dm89+KotKozjyhbkZxPNv8S4yBvy5bp+v+NHQx931jKPP924Mx11Q7
r/W3to660Ueqfhvna/8jDdNkgECiBf9d91sl4mOTQeRrvbqtgw+K9P5GXCCFikjM
coCTflPAfHTq+4HaRjLpgrzf9IhTSe57czr9q45vcZPAV/k7c64XHkDNdwuJFgGO
lsQpmIHHhy7eHtOWhCk+/ObIgHGGSXXyvPihXbosMzVaR+p8p724CkV4iWOewvys
OYtcod3joyEh4n27taphliAE4FnVuRNkqvV8CJOG7hrSgyZgDQU2+ALF+ZPWXJhc
DsVTzCaEVMgTuK23U5+JvUFBXHUuScp1ii3kf+68Gw2l1wQ6VJW5mJahQoMGESJs
DvH8315SewsNpMrvsvxVMTR9PIzkc5JFaVFRkraiJwBwGrDExXpuv8X5oEN9ojHr
c7CJTqOApAOz+4JbIYc1v+LuUPJtvhCFJcNW/jRU0mIW6ZXJRgN5GPnAg8BiWFuI
KCyJOPCGtX+zwIqiCRcNar8StScn9fjjAdJ3C0DAfDSMRHVDV9mL0knQNmE/4ota
wfjlo1Hc0J4lAfMgmnvsEe5VdgjE30z194TxEW4XHB7LlcfT+RhknuE+jFEits83
qPyVrU4v5FtJG7zEYk3kKIji1N30bl8duK1sLve9MkOeIMNWrZTyGeh4Vl7gFdGP
EomOVunqcqmPYufBNWyxG45o7g4tP/t9tQowtaI4YcdblCkRe6pKNkyzOaaQ6RvK
IBWBv1D9u3jZEpWZlPJpTzahFP5mggNxAdtbTQB9MUwc5qNt3D3EqNGhxjCsMV15
dgJuNr6BjKPzXFIT7q0+QbQ0/a3s6nNHLDMTxJNXOIVVHR62LVfesnRVYE7AW8zV
VhiFI06AGz6UTvOlQ+1JnC97CAoBoh52MSvuCm8ZThDQwu/+kmbzlMJqBGb9AYwc
GMblGuVqZTkdsswskywvsN93dHNsIJkj6r3FyaSABF32DOZHVibsQ2jAVlAQiZlw
0Kh72HT9siYIwNAziSlvT93R4r5lDdpO9aSIJ9bxgYnGW7//k2E1opAA20BADvQK
gIoJYqIgtr0f4yA8pGDNWGai4nenIpHHTbFMi5+1zUDNA3oANszQdrkSgIrmzZCd
MDiCPdJvEdkVEpHsr3MT/706XDP/3pRJxmFU2StzAud11TrJRjelMQqqhMWRhK5K
xjH2d7v/jivnG35EQLCNSP7cuF94+YV7faM0jSfQr9PaT0/uawzkiZRws1iEQDEU
1Mw5qCwfiaHTXcYU8bweascMv9hqm9PBJUTABxbAs2koAsEfhkR7SHs0X7Cyifey
dqywhQwUEtUKGn+sTrqYUo5jbbb1GkSgHkqZvWlQL1kTYd+bD/A4Ew05rE5rSTMH
9Ayrq64wuoNTHUfc7Sa7Pr/8shHfieznfabfwYcmn4b7CwcPobpvIbeHm0bspzF1
zjAAQxhDIg7Jmkc7CznpGNDKImIpPJ0ZpZcE3SPEqLq+rRwQARMnJJym4NHK45sK
vxoPtkYYiVk6Gf+lXzFW6sOFc0PIUAUbmuB/c6MccCMEMxhtbqBFkhNOWSr9Bnzy
kByOc/BYBb/e16bB1usI3jj4aPRtNQWPvKFV/ViXpIZBgxUZkUWWfL44ez/TLz5o
lea+hWZspQi90mVbuO2rPnV0VBI5zh/7FBzg3eSA3kgbPNgZUdp1Tu+eAsRrjwLc
J9XwGsZek6EPWiT2hZj043fopBy9nTG3mBprPLqKIwuDBj9CpDmYHgzJ0vWKXouX
GxxfwZQV59fc/mhTMs04b99UmTMJrzhvU/DGpkBGQ9MBEdU2JiQsW6wDGa+XS2n/
jDDo4k87afPIu/FoBLR0XPtThgul8Q9H+O80OEbtT1gGTBmwUotCg7hTd7arIRGK
4BB/UzteBABc1cZ2CtXhTkJ3coLt8BdzMmvgZZTVYobd+Q92PrzoRuScBojsHAhV
2gRfQWCVNFSU16rUikW+dfvYmeA/Dz3rQQZZJea3Wm9bZJvkx533i6vu6dThU67o
w4DOO3kL90fZRGjP8S+WVvahk4eNfYEerO6qcM6QIa5WxbUmsGHc37rj/9n8t04q
yLVSdr/ma21wc7FzNOYyBQoQ7IYbavG48qNanc/aser58h+GBjflErx7MyaMjf26
mqQQqomQRJOKiJJ5OLW+O00qblKz4IiX9hwIHZeL0a9b38GInYXrpZ02SYTRA0IH
yzzEjWNpszxi6ba+HL/mbIpvTrbyeimzxis3WJJkqyrRbNo706ocJsH5CpgMUMoV
SMhCfADPTSMzzSopYpO4b5WoCqps7so1jZoCsQOpfBqSZZml+NQqLVCcZaZOyhoc
RhBkbVwsXkW7UUXr7aqSFFOtEJjS/F5lXvPz3Dqv14+o4k4Aq2DpAaGYggLDJKI7
/WzHAneIL3q62cweXbxdai2GnKiesd+hr+HZDYrvaB0wnHxFmT4iLvAqQJNAstQ2
Ay6v1w5tHrXXo2kTg4T2br6JeeNZnpE/5zG/PUQjtfbWF5mDWp+3F+0pdpQ9W/yB
x6emY/DlCe/s+MGsTss8kUKLxPeDyHxAuhzGEHQWCpk+ZIhN5ykxKTyCLYt+Pjgo
PsWWTjPaVMHip0qBgdAvAMfo46xjtVedbB3xkI36ESG/uQBG9vrc/rVJ7ybIQy3E
rNG7fSIQZW9HCoqdHFxmqnDQmDq4DEqe8bDpate7s34EIZxLQRigmZaxg5Nut9ok
/DVwTbarqraVV0Z7uvVG6PWOnXrMQSAhNL6NfLeVF1SBaGU/tmEmQIrmaBXXOn6B
EexJ1L+5B8PJQHVDPGThTrDGI4Qq5/DeOin4jnLdSlO5HqFCuA4KTZedRCFudPTf
zbcsGKtgO35BX9dJ0bdz8oOiEM1sDjRWMXdPoNPqHRLxCxkjHpHQoQfckiY9zZU/
akUWGhzSj27WszkrAKr9Jg==
`protect END_PROTECTED
