`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NVGetOXaLDSWFOVouEcPCXzxmJxu76s1550WIC8FfXLky8BY1eQu0O6gNHIc0nUX
jjDy/vG2nJLZWcZMH00r8ORzj+d/B9xVCzGJfEg/92dbSw0A2wKF0AAslgEWnJcu
P3OtR2nmoGtsAbXDWV7C0BRIr4wyEMb95Wxe1F+TpKsmiUqp/e7jSVV9vILeMrbF
IacmL4P6abdvwAmD7O5FmzZ4ZYwEwGQY3GAcEfSlsfSQZM5ns7yHObFhe0/ogHVH
485GhoWktiHuKPfoJIzeIR1BjrSthTP2/o+FcY9DK2RAfuiFvLcafURtkPkW5ItN
OfuPTembJHIaQXPOAydBiJoS2lj/sdrTxp7/RE1DUJTdvouBVjaQOeklOmCEsUZQ
rMATMe/Xz7FLUVkwaW6Cft4L6BWQH4A7xDHB0bB4g75pI9UCuTQMbmQvYREMe2rz
286AQMB/p7xdruMvuIpmI+c3pg2zGG43y85alUEjbxlxdY/Po2f2WiDqEBKwY5qA
Ey20Ax4+0/nR8NBsxPnZzD+/h3Nj8sb3Io3o/BifUJ0wqYwAvDyelifQSPl7x18v
1ym/jajulRLJjvmDuqZiZA8yo4RyHpNqRIBbMGGJL75Rm1Q6ob/WS4RnRpI6zdav
4BBmLQXMSgluTQFsqqNDsQ==
`protect END_PROTECTED
