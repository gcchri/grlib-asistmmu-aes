`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7wXb2XJQly9MaTTirAvQ2Wl2imWOrZlUY7j2GY9+jIapavG/ZO9HOG5uBdbJTEfB
yJrTQ6vuiyhXkX/24g6n6SNkXdje5FPZmOTSIHCH3gx6VhFWmxbts+GWNtFITyqN
xURJjzcbF1erzTchYaJhxTIz/+j/hYg3oPyGUxPJejSGF0/kope1P5f1lEBMZtAJ
xTnRyqOeHpauaL6bot8Z9fDA2bDiXaN9xe3EBb2vjzGL6tstlqiQ49xwACPy9d45
u0R1EbkP+Iko4rOimMA6drRxwqkzNg23Vy0DPyMSHZLbWGNN40XhQlaY83C9ICxM
j9GJrocKGwwxYENJtgH+xOXpYmuJcQ8UXk/YohHO5AjZyxHphbHCT6ldS1QdBNtJ
TkUujoRIWP+N1Ko/xR60ldQxe/U4as6CyP+10R+XYUh4hRCGwRR/+xSl95sy4Ftv
/fDRVOAqbitft3+fYw5zuV3/907sKn7AnEb/V2jPRHLNH7mc7UFSGMU23eEb4ndd
zKPAzE2D2FJ7DS83itJYSzOEJiEWlOv4nPMfJVdWPyl6x6chapUVfS3fOoMv1i7l
hYHhYjoFUuV3iTbezJeleQsrcDGen7DRHAu2nwmV4o4Tm3wv1PYZ2l64+k+W0N8B
9BXQAET+AsY+sxvo78VTBnnWR/zQcPHFP/bsAjY3mOI=
`protect END_PROTECTED
