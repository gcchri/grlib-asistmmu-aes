`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wzAxl4MWJX04ny7d+D2XaQIpujX9w91y7Sf7bpXjGKQcyjlNXwnDhY913jDNcBKs
qCDQvyRG2kyz8emRDiP2UZxpUvto8gJlNnk1RT4hlQ+RukqLdJgAGebwldt63MJ4
Z5Jw55ca7HGLFDGAmDsU8X4xTDSx68A5nO1FCo4XS9ok0/9qkXToaBaIEqaysfCo
Ul7f6H2uTP6qGYmiYe025M5x+YqbUkvXtmNgSyb29nPi68tbWIkVDdHhK7oMZPd+
X61wHFMKpSy4MIak32EMBBRas3Sb4fkUJLUkmSog+1yiQ9nNinympIOKUPWr04np
dw22Vd2OwxZ+ykfWRDVtb/ZCOUcSJcXp8d+RdSlw7sEKsRg1dme2Hju04sd8PeAA
fNGUWfUW2PIYTqZgAyTjdFlYdCG8s+wm9Zlyc5CNbXWoE1LG1D56F6QJXGKJDunf
ZqSaqVB8zeW8wQS5/xCTHLQQ0aE3gm2k0Ml+e0vAuYCTyDe1WfTpfhohBgZb+rku
0xiE+BEOQYiiQNnkdJWMLxFlm9y7ZS2NLhybrAsj9Jz7wforELr6e4iIzNB/eER0
O9rbroBqyij9QBlphMnwhLX8H3E4+AZ87yf0MomFBuC0zO5JIm5QWu8YCTr6ZYA6
13LK/9HgYBgsFuOYV2ZtnwlBto2iWeBVrFLaf5vnQIpXu0/5sN5pcP4Q2+M8UYyO
nhbNp2WWUaJF+t8iSIA3EjTMyr/xWcQo9en7aFFXlpZp8iFalqRhtWZp5e963GIl
VxRu9xVZH1qvmhWdpNkgTxepsD82xT6PIYPUCpOKSnFcoRjvcAPce5q15vx50AsH
/YYM5NIL1koDggviQ1c0PRCcgmM+mze8iWj0B111ZqesNMv+xy25/vu7iCRYflPo
5ktT0jATxeg00D5sqCWBBAIuFgXQvK6tU2+h5WWV+gSV34kpsW/O7rRvt9/mu2LA
q3GkHmObUsl2a8WAkG2y4W3G8M/q3yF1qNNwdflSXwiKN9Rt9JQ93R8Goq6HaKjs
Z5oAgteu6WZFVdxesOe7ZsmKEWHcFTSARuwDkDxXu67SNJmbBJOf+s5ODFeCfgkA
ol5d2ZQzm2x4krdcRm7dxtSOb1LXRFA2NadGgDo1ILgBaB6dTNtmoRG4832aRynH
qGq1RppIhshJYz/eIDb8N/42B4vxDVfyRew5zW2ZCYJC+2SWIW7WdZrJPHJNsli3
1mMLpjN01E6pClaHz0PnRkA0HK536MQHu3nwZ815vAmbXpvW4a3nJnD8VXlCYjvn
d2U11pMPKLyZNyEBUvVv1MZWbudCfKquSeahMTRNIyK+lciFouCwDA1tYuArcDNU
UxqasN1Wvepx+0Hk3vs5zLH8JTr8jDXLzsmIbb6vzKZD/gnCR2pFL4taHnTWOlsc
QzAbYQNCrxe6u3sZoJeZMPmfOQsritSjIrvn18UqGgQa/I75aTakC3nJgQZ584uE
H2e4ZmuPxdPLQyPrSToqTqdoHh5zOfxIpfnRRSUlwh56HqMyMPcapBftnagDeGkb
z4kT8EYxi+JHIihxlf+cRhhOC5PkqyST9nGR1GFUUQwd4q8KIIfxdliQzT1CmEEx
c0hI8YO9qMBTmuZPmTGt4h5Cpq8QYwDekJaPNXnrwDcBOaHCDEwecVBJEu1VzHp0
3dfmeChAAcAfk0on8U0+JD+PMcp0zrBW6yXRppxS4qjboilLm8JQhL1Goto4q9ej
3YTRRWbv53ofCz9TUClcAMFisJkZa5avqUMtdpoDs3OVO21JQK1kuXow/2Am8WSt
mPZllCHWoKkB8j9jsKgi9y1z64Ik7qRVQnTh9hQ5jHm42jIR4zcn6pz9gNoqJ6g4
PHoLB+PAW70RfNdFjWtaecwkS2AD2liGhGqJWXabElaoiF7SqCwv+Lla+L97ps0d
8Xl6OcVVC8bsG7B8Yk6U/sxkfd+U0TMlEhP9fFEgKp8i26cSwOInY7Rg1olIVh3Y
ofGaSn7vWMzsQAuCu7EbttqD1FSRaPOBzioSdgnKrygJ89dJTwn95aedkg4otlP4
`protect END_PROTECTED
