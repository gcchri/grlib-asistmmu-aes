`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gcbU+biRsrqtUXFC80ok7X85a6G9tmW6J1/PYjjtWm5wTy1rZ5IwZ+v4COJOXQuf
+R0GJRqB+tW/bj2vnouvFgih8RGSHao3dWeFG4LPjDDx6TZqWvXHPhnJeS6Xk0Rk
6RtmN9+Poc11ngR5CDRhpjSDBh/TLeLdVAbHpHklVq9w6v7eG0sZUHaUXrgHUG8f
wK9STpJ4AHFc5AHUEhY1G0EspK9c8xkWbKnDiMGlAC60Wsm6dykhsrgbau/NAtys
/cbxG7rWC/go46O9YEbihjEdY4CoSuTEso/rg5pxogYl/AaNjYJlj8pMjD5IAFyE
`protect END_PROTECTED
