`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zmpCBM/GXNTfKYuOPIvUscBsKaprCe2rvQD+Wpp4mGtUxFFhj6/T0tIdUmI7LUt1
t2kCMSVfDpQIhtoQ43FicJiTk/Q8OuSzCT7jThB3rnQFOfYj1gzvSsdd6TRQYI+I
G31BMrRaksrnfwhOfThiWfqsuu3cO8edcHcfxkH/i3TV+3dWt62xMLP6oDbqjpbi
O7bIn0h0Lt2dLEe2hi5vaGPVknC+i2eTp0Mo83TAvKbJ5ahpjyppHx+kclKisTrO
p+wLJ+irmB509/e5/mN5enN1hFR/NHVgj/IDcemi9JEhzoMpOkKX2KhtgPdksaq5
/hDhJryTcd4IyCR50BYd+ajGWIN5+GY+C8OsHbzjKyMf6wDD2XaI4+1j5velJXEZ
+7ihBwa5UMRcQJ9ZghXcoLg/b+R8XdFt6geO9DWujruZ5Rph7BZC+FRJzqN6sck1
bV4g1FrLeAPMRbdCJB86uabXiUxTzmjWCt4QN7WLOa3Eiwo0M8qFA+q6K8GRHsKE
LRZX1S1e53/kcdHiHb+Xbl5vPxvnpCEE2bfzleb5HTkqGX4Ab68P65nZTgGaJo26
XeFy+F47GSFo6DcKkduGu3ou32er2drGzJ7wHSjza3mC76yqVV1iL5CLnXmyrkAZ
1l+Q/0EGIHmsqUWh3WuNZk8xNPlIoqZS3WyJtZMNIB6hsf6U4oLDKWcQSrDPI6DV
+NznM9AuyQDSJre0XRI90DhkEL8G0ZE3eMD0lexY6HJ19bpKpysFoAI0ZtF0LUhc
J1QENwDOSir3s2QD5IC1WQ==
`protect END_PROTECTED
