`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DVoxYxoGvU/fqux2AzfcpVnqmgKCE9aC7EJQLltrvvx2CR7FxI4+O1IclN5ZTrlM
QhYWPTTCBrzANzGc1NAfk993m8GW6BobJivo5T2TaaYGJzQVZ1bs71OxWdLu6L26
lUFYIeAkgHKeWvhKbqa2FsTweT6e/4uV3juJMzTejseThcscjPXABLYeXrzPHLMo
X4bvFmDEbhHUSveD2/pFrlh44giKH8LEd8GprVwON8ZG66j0tHdYhYRHfgzoV/VF
ptE8LlScFV/Wfn106//kTxnrSsRnATPdeuCrDcpAJkiWQrEzfRaxf9WU1KUqPTYX
S1osoPSK3sb7JiMniPsxqPtoLRCM5KAtwa2qRax/Uks=
`protect END_PROTECTED
