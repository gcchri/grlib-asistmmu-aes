`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8IBxkv22sp1aiCuzDeepTXCZeBdIVC1UvPpvbEU4Nbhh4PTRT9b3LBSRCUbXkWEp
LSVnOhK4rAl7f94pcbzvyQjmijdTglTnPnLk8rM7dNxcNxICWuMN+6ul5VpThjv4
PNRUuiMvTpgNEUnu02DfQEXyoZ5rXppMVy7xe3/c/oedm5g6YYzBiS99p9Q24Xyf
b/X0QtLYqrbh5Bb1PXM/fvIgujPE1WKtiq/tSWM/ApZyDd0T6Aq5d6khhN+BvPUJ
2IysfhAtwiDCWsk8a+MawppwaTVWwHy9fa4xUPUENtf4zntPGClUDRNgCaVJhJXu
+8xUwnjsX5lPO0oDzdMgNb+Mtzu6sSqdE3ZLL3B8zmMLhrqrmZHMIxBZ3Y3k7GOJ
sBP5GdjhqRAGgXEB+OIzZ99GTzcAMPo0buu+15DgUjI=
`protect END_PROTECTED
