`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q1Ddop3PEJItXXZ3aiwSF09nIZ6cTHHoEDf8QZvFJyM1j1R6bFOafFjHrBwDO/tj
M/uQCEbxBDbVo9npGLuTsqAZbZ/UHvEvJsm2H7JVpXxrm4LPxbJ2mocJI2bejdSW
EvLEOY1jsb72lD5X8qcroVSXofjCyKPzfGhu0jtd7hnO9a739lOwzGh1sJX0MreS
Hj+f7JlJ1worzGY+fcv3Em61Eps83aB1pI6m/tEk2kj65bCnbo8JN3fwJ7L+JwAD
Hqsqhj78YDeN61JvbifaWw==
`protect END_PROTECTED
