`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zfbnj3qa+OjdVroUU14eW2MvvkTt8ztLn82fKqc2Zy8G7Zq8TmUVCALFHDqfdCDJ
EgijkhJOkkj1G+7oXyJm3BzwIMhSBIT/Mc+QcoU7hSOo2Or4J+y63BceA9L0h+jl
6Ii4DbpyGcrrFsC+XZHa5bDz4DApEcGg3rwRcq859dWvQj/B7lGAB5MACNa55ASK
VdvuCtTA/PavCVQQ9FjIjG8MpN5ZQn1s7ZgS50+t6O6GBhNaJiBVPsreTcerfhZF
izZ+2h9oygetYVmWUxBumOwNPQ+wtdIJ1e5+nqqCYjvmrF5ftRvWch+Ex/Ok6Og7
DdyfBo6ybX7AKyXBAOE3A3nYHxbxNpMvF58g01sXaQToI0JDgVfXxbbeeKJktUVw
ZJ9nvv08pV34+m2jdXtRmw==
`protect END_PROTECTED
