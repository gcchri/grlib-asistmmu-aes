`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dPB7ubdxqKsG3ZW4GojDs773mN+e3d+Y55ybB86yf/3MApr9rS8bzPeJ3PD2vIZE
w2GBfkPqi7WMiAj0LK1BHI/ZpjWvd7nfz1+VTA7ScwJ8LF+UidZ/VG8JoKnADitE
xRZbcrt3J0GVxSrU7IYHA1Sipm1Bp/5v2DHdBxkPFOxvcBviOeVb2kVO46sQh/+6
aWg5Zqhk4g0OtgHD6TmTjW/JvCUXD2VpAhlRQ1uOppPOeyxtpJeRjGGZyAGmMKMI
syJRia/Zs7CWfckM3RCmb/1aN6o1u3gKnDjvlhBuO6LlPWLSmDXd1nScvq+qjgA3
RSWLfg4Gz+LbnWynK9sON0rDuK9cHe2gtKR/WJXzkN049Ann5BzH9Rh8W5cBdDbn
M2pr2DGDPxQk/5eK28SWbG+KBtWMTjAhF4eN/LpE22ls6O/+T3XSvZsEwzO2JrSC
v9uCVMD0tRZmFaQeLl1XlPW6EVV7gE34Qj/ykxxfy8p97ujZ59BgH81R4a2mDpk4
NH0T6VeG4RSwXuBEnhxTikqaA60uft6U3Q1/kC8drz8Y4cTtRtRBl559LNCCUoLs
8CJXiwshEubCvNJfXEAFGHfhDFszC9S0jqbuLxZDNzNN4AByy/UUHWXMAD/P2pzC
zErrckZbSTnESNdq56CaFLuqZI5OBjRf/z51sE3Wo78UQhvK0wA1C26hmy2Ll7UT
ApvLQMplyR7qErgb3rDqIa68rubkBJ7YONvNm8YGM+7R1Dy7ZNls01muVrsodtPp
/iSxPtDwHpvZDPxsDg/lBb3mXlyxm8vBZXcPngEPOQMRBU7LewqaRzzKprWu9qM0
e7QZJjS3mmctCNWiewsBOGG2XwqdsfC4H+TxerunogLP1fs7azRJJACkj5jPsB/2
Z/LviZ7bUslllKow1liSqwheqMyVHLm3J5Fpnb6b10nALEr2x3JEZZw+oqe6u80v
CBymfQ4gv3OC/6zyRccM5VhGTs3gMShonCp4Cm6RtnHSaSinYSgFC4Znt/l0jU93
i+KfDgHWYN2sv0KfiQYwRPbMeFr/3wcFE+tLj4M8+VkafSYn+zFh9tJBZ5Q8I9op
cq1ESWW4zNPmbcqBCeWXS/k0UVttiWAVRTrPA0YO44Nqm6oYVx8RlE0/qznKpGlx
9ijy6tXoiQQxx+qZjHwm2HCb1IZJYBqq9Q5zO2dV9MhU0gvgfiE5Zstaime5zdIf
TnVj0r9pWBqHTlpDxPZEHM9syRoU4WxdayLWyYOoUATKNDEUB1rrhgP7u8bo0LyT
`protect END_PROTECTED
