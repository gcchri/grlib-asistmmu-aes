`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NlQyvETVVAS5chvA0DWD0UNzrFkg4w0IyVRl2xTi3IMW4JKShdXfNqYROHh9eaQ1
5srDw/i9tVL6Tl5pCkZ2/GJS1+E9bOTBB6v1qkguUTFDWDJDOx4gQfEk2RJvczDM
62XEtsk3qKMi7XnSOtzemxlLOl3zmxKHt2NC4r9kk0ot9ASYQqFXgAjGPJ35zH2f
o3PBhpAOhjAPDlmlS//RqoEPvDmzalfJahP4NxCHSzq/m43UPvyo+Oz7typUeNwV
NBMzkWFSeOlI3NIltzvN5X4gmtSs880dko2ynIsG0Wmxfz1DaWR8JsdrvR7fS7MU
RwiBKWondGPmta+o8bjGBclDxbfv/RY5R3d/rt4kO4wPIMDdXZRSHS3yjhp9bVJH
qv4WQ3GwqYEti7IRV3RyIqVE2lTtXM6MiiKQNuqt5E/f2JDD8fnqcGaVibBnIgQ+
tQisjP6TAMelg1frll75Yh3gmeSvLKkKAsfWPLcQguy5/ww4j4+6c+Idb8jUVQ4c
DlMCETaboEEUbGuMlVb29vdzMRR+a2SY6aL4CUjJnYPq253ttJRlw1Y4G4kWBfNc
KfGSJ7f5TOscbWzhiO/sospT4YphFvBznZLRSyh1wNNtm+CQWD7moU4b3Y7aY3LW
LaAQhaF+uKWPWxnpnlX77Nlt1mcaXB0xkx7cTxRfpXsqyFhZ8Pu4a/t4pCCDwOA9
8NmIjLmS/sjErXTfJpCoodq4vX6bDUX0jeY8AxbQjjJOJJwls7j3d83fRicf0Rmz
sLaasmFPPeDWtSUKNjHj4QTPV2ZBNiz25mftCByBJFq08zohNJkd9gqYDzQW4wrq
ZQdNhv6LgmYMZpbiKTN73l/qcTD/s981vMWe6lvmJr3oiKLvSY4Hf92xFLH8iTAJ
MFpXGJ5bDz3Y4mWedG4Owd68//NVRAqfm0Awg7xWDbegMLLWjLBp+heqe0U3ZEEZ
yRcHQVzPESUwkodxnM7LjD0Mm8CZJpVcPQ5lo+0Fvp5TGnI0fNTwk3+Ri2hffYLu
dqLYW6K3QAusrAluyB/pu39GqFHNi7FfgzvycJZvOuhaCsVaNRO5XOcc8ZwubVMu
PnMFLoU+PBZNscV4OG0uM82CQEVGLnQVvGtYHB8RXGM6bv+ATEETuP8fHOeoL1F8
qIx8i4HdBy51p57H3AR+HQdGCFP4HdSFEUNqOVtpIDn+qPk1BBhlz0MIOWchzfxd
yXadNOnwkY+qHMV/rNlGXohUH5m5AvSOQ56KvDiiVfbh9k6tcbjMB65aRrqTTqxl
Txmfj/UEPcDnWpgF2m9IKHbuBVoM/WAdHcCWZl0QzCYhTALT78UT3rB22zP8hNkS
3LzuaFSM0t4Z5Zi5UesBczRjFgSJmHiFUnBjQeutHw3I/42rrLZ/ZyTYa7pXAord
vz3pTklN8fFgqOlRXRIZe9//x27lJP7Xcgeq9NYhHOjSzpeXm0Vk2WRmGbZdo//1
d1UMHXZQz+5+YmpBAicl4ZR8zv5iyINhUxucJ9zOvM/KGeyfjV6c0rWpi0cRgdVP
vGdayW8UhTaWqNqasTkJp+Jyv5nRKp6qaEb6cHEp3ZFj8UNgiEL8jBEkc953ODAK
XF/ryhEl0g/KpWVrZTWYdAy+1Ub7B/E5J0gY6iBcEfAzY6EMBVAeeercJPexnReJ
B/QCSX0nxFWlX1l0Cxfk5UTvpnf0TDo1qkysuGmPPrV64MNmq27jpXNQZJl2zRaz
WkjhNI4EEKjAzJEhxY1zv4cS6s9QvSXJYe2O6hnAD2xuFnnVBciY1QVDDpw2AAlZ
50RSe37PXp/u8QHP3jQ4uB3V2oFcxBm+JyJpbvtDyXr1Ku7iHLN/+VHNpqeCU6yg
cinMFnzagbnlyEf/hXxPleajU5hNl9w0te78UqmzV2WGAQM+voUTO8e2ERvmPAdq
FmSRSgM7jUpPTytHvg2EYGoyVGgQcYN/XcrnC7SLYfVt8H3uIZFUFssBn9Eq8pfT
m+f//2rdOQeyhuun7ofzbMV12zfiZmCzs1bDolrBr2GL2jicvrrLvkxBQzZRl3b6
ENyRh+HiN9qAisQHhcB6Y//ninaNgA655UPp2SxtjS2Yi1b0579NrH5QMyUkmnoF
sBUVbFrBwyKzuAFd7Z7pbRsiZ/z0lx1uWbGLcdN7yIvNm+e0s0OD76mEbGomiu24
`protect END_PROTECTED
