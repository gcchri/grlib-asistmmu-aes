`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
igx+1bs4OkNc8Dod7sKIkzzuBoNHHK6Dgw4o8InM2eJwwlMaglMwEM3HcTYopoj1
7Pivw+vbivTDAzbFmQctrHcoDqTnO65xGSPCyfTDTqrTbJs2eY9pGhT7S/ni6rBm
4ieLhlGbtIyZnvcKVKMtS1lLyTgCiFbLIiixsPexFkUYjYkKlRyeGpx+KLd4/1Gu
SNf2ll/rIoUUhLTd2A7wFHKb75FEoNUf/hdqjHuA+4/buhmY92SflM0xWhmfhfGc
4AeaX/OG3ZzxRwuspBSZzA6iwCpDY87L6FrMhGcEBetDXLQkCCHnWxW/iv8oAneu
vyb42x4pp2CE56RD5VHHIC4nxphzEnkjjCIOoLyh5KK+TdWNqJ7YK6woZehvIiyD
y5/WfXb0qcpm0nizIv4gB1r7Jvm0UPKdLQ8XY1yZvFHG/U9L64EQxlqglFh+IvBw
y97gVcCsXeBTJzi5hFYznwEY7pbcU9JDflZqdMGu11LLlWqxp3zHvmBczHuKpOhs
cT4qDVRPlVm4W2/HQEPCMm0LXrWjkoSMZwinktiCGXv7yj7DncyreMT97BKYt0oI
6SBZxmzsS73SDxqKG4xBrYWZ8AR+g5WQkNTKC0ki2S2tDBlPmhnNZnnArKRSWXU7
k/Ry/HzLAGXlbhpbAZxkJw==
`protect END_PROTECTED
