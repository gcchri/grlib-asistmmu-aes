`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2cSVSAGhH/MBXgGMvWCXQvoW9Sw0C6Isu9rtaE3DUOr/YiKntgYpDHieO3vjh2aM
ZLoS5Jqk3ClHHb5+/E0YwLif5kF3VhQCfAOxY2hKGhmOuFmlRCmlw+AD3Ka9PWuv
auwDJH/rbph6diHO+UREcmoNIdLyr+0gFA04Wfs60QMZhE/QXicjE4NpmUGy09Hn
JqeOehheZ8phmH+Z1k/0DcdkRwCPdJQ/yu2mxZKqo+Gl40hMpHczvfdeKj+noje/
J+5+w1+JRE+tBcF1txFI8IYcpILqqcV3n2r5qQQf2+rQwFwMirEvp8d5If2mjAeJ
+s4XCyFnOJdnl5lNoYnkKn8ba4vUzZ/lY8YBoD6NcbWuPCyPFFJE78mjSOlJc/0b
HPB/p37OFOaC6/g4zhk8GG0D3L9UnUDJ0zAqRv69SUg1+AZRaVTKaG2NdOVWZnXm
2sBb4P4MBfsAPWnRrxjm1UUUrR5x6Hy77zmpNVt9w8FxFHHOYFkWuX6lxLitm1H5
/l1W2BLfYjyEM/CuCl14ommFL0iiW7UwJ6kALOuO58WScOIvEtGshWBl693NJ1ea
mhlFQxVuc2lUkaPRH6KHJnNLzAGAIs80M9qzbT/+nWJLda+hhmJYprMzwUeZWG6D
AtG39RXbsSzhWZ3bwoolK5/J8mNTsvFl32mnv+FHgNwO3vmT/WxQtSKfpms5RJ3Y
2NY9E1mYMudMdLPg7dK28Y8ldNDqXsRia8KzlkCF9o1J9UEW9MW6VoiTh+pmRKMg
CYKXty7lB0uyZu+Fk/Tefn3mnYAKgtglNU3Ib+bFCmsB7HWEGr8jamrlUCVtohXw
Yt+VqdNGNOYhN2e80PRtu1xhs/650S8Buncqi5YolBIz7fn7Jky1I4+4qkDhn9ky
0MVeYTpQTQ2ocuOdJ2g7pPE9/bLZaEY3BDleVGpPEsWB8zPG6ua1diZrhUxaFYC6
ct9p31/G5fIfBLY0i1EGhxL8kLvUUUddoH9gwIeaK/gIMEu1iJBQrtU9yO2Lxudn
xETBR/XT+QXgJT/pavYlANSlqTTrjp8r+Rtk6T4sOQdB42Ty50tSGzfdL9nRRDJo
AYzqL3LxpkSPkmATUlK09+thFK0ni32tfk1TqtiCau6swrL0tQ7xdxtcyEgjZtsA
PgL2XwFRFPDPyOMdmTw7hUSGG+oDXRSYU2Hl25hxN/3oI9pohgyEhne7kzGDoWD8
ojIemHPq2JYlFWUNjnq0ZUIkAT9hch2Bk4z/tBGm3/4nuzuZ+enA6rI7hiKW5dhZ
plc1Q7M1yZ0nVB5NvI2DPsIDofZxLj1dawH0xxEe73sZzXkEZ4FWuLtdeP8bLaVG
zH0xCEP8R+dni3N+joNrrkXIoL39zPKQ3Op2I7KH3KdX1QcemI4B6Gs+obR8yrXe
dchXDXvSh0y1+Q3CzTCSUsUfnSXGVggH9l5bdtSPJgW/ZoVSEra2HzEjnLPntqU0
AigUEIP7YzAreJAUkwGQJEmi1OIeGqEVDIc/+e2n8ruqt5kjgkuu6PmxCAAbNY8q
1JUD+aUd1+CJe/ECtZ36dXBWNuSMlBbuU0/TDxEHpnkMpAho9iJUsSUpGPZjHNN8
RHmIPPz8NnPnhgvfFE1ecyDNYz6L82rJxiz7kzcN+V+oXfNe6IHx2d0uAjB/vQyN
689hr/hzUKBvzHta+UYDdL9bkxkvlrtRLK9tVoLo/eyA8ChJd6hp/Xi5YOkvWNSB
qAmCqrahEe7s8dOW8Y4NxaT3NlHvrtlUZAvkhjaKXqIE1qE/cfK6zkTO4mxOWyyk
c8T/auXXdpVNuLlyCjg5jk7MYeLzWDGpo0rN3z1nlHs9ZFUkK4eVmvAf3uGsO5fb
5o2LpGxXyCaxD8dUK13mOzWtD4YqCyIgnB9tBrA6lBhuhC2hQDVibwGeD+ZI9gZR
YRTUqY4TmZ0/zMJeYoxp7+zMt3Da81ZPOPFIdRP9k3Qcc/LIr8Co6Kz+3Si6O61U
KjcvoVgtHjiHVfxy7suQLCspKnWxe9Kt6r4260gHWu7rNWPSMf9kwBFuocOb51Ts
7/IelZcgpmfJ5CNf3b+FgwnhHtEZ8yD1hqQN3Jrb/qPa2ioUP2gEki+gv8SOJPBw
2U/7EXIp9nVQ0eRSzC9ABC4g3lEkXO1oy1Q4mFEosXK4d3fGhUzO0orrk32V0bXL
9BsKV+zfd223kdo39eTK9T6kS1lHBdCokys94CH9y2lWTclVS2WGcSjK6tMcqFFz
rA0plnY4JoMOunPcEsjQhOijylOogH9DNkkbMvzjer+z09p6crQH+4RCjR2kbZIV
T8OFaZdEw/8Ze2w2cC7oa1twOL/n8dR0M7sjpCweikiYqx2GLk/tIslGiUlwLq0s
QbYP1+hywLguFuu805AGZVsDfwsAlVAxBmLXCv9OHoA9Lj0LXTSl9N+RhkZ5JoU3
nVblysIhlvemqm5iG8vrBRkcKkwwYU2DBw2jgHLTlYvMB+HKXTQ0U9z3YMs/TL59
wdKx3n27GuM/I70/P9c4yBS63asuAqyGKss7IHi+LxPGcazzqYP9Uwm49D5Pt0Nc
A15y7nMrGFSBoe1n8CS3biZkHHG75l8eIuw/ZAHsWUuE7a9BMw4UgdEEJ8sSAc1L
ASf12H5CAinUe0xnAgf8rug1PM5dySkKKsmgmNnSoXituBUpqTWiqVK4O8r+2Kvm
vz9bA4Z3PHDouytacvKmXEK6S/++KsLe7F8qUthQsktQFHIrqbQS0w/QzspEFRj8
NRgA1vi4ijwJDqjbvukZFxn0kDexwL6nMBfk6GIuOtEQ18vUf/LSIKfQ4SaY2g3t
+zLR7TUqnKpe78m3K5nuxjkNmKBc6eIa8/2Xdqw3X4XShdiXCNIOEYcvEVGgZtNG
nRpgbkuBvFO3QmnL/xkXYBMU+SnOnlClHcHZBfI+OImCCGWbp3bcHxeXLK+C1v7d
nvfrdQ1jnwz+y1R6Uax07j3efyUX4WWPJU1sf+0FdxNwSasVoxgwarUFZw0mc9Vk
4Df86rwRakoHbuzr/PXMhMJBPOmlC0XC4YPgHogw6IlwtDhrlfTFRgxhVnIkIF03
9Fit0Gq7wsp4BRdQRvN2U/U59ohm1PhtrhJcA7K4oXkT1Wn14bc1UnqkWTzdB4Pg
mEItKQS0v+AwkLsDzPpe2xepjiwJM5r0XkxPGC8bv/MrY6aVnru6stLtaTc0csnJ
ZUdJZDCifG7UAa+Qgf5pCl/RchG67x/OArI28N3uUnxdrYYz8SlE9GwZiedxsFyJ
SUhIeAI4uOY3SsAxIEbOubsOWOd1GarQe3KqStyAQ5H6TGnNqGccuT0J43LJsVSg
7p1rvrs5YYtXXFszkJUtekTV727u9DVwwLIy8DWL/u7/7EOkz6RCBlaymMgO8uBL
my8ayk/QYmmcQ/vZCiETzinGhNt43kGkKY34M3U26a4BpmDY1kAKteEGLcJfkjJ5
h6FIRBM9NcDSr7LdV0KK363/9G+qWtuNXyalbu8jIr7Xx9AWVkT+2BAWYPd9zkvk
bU+TFRlR5WHREd305g9zqEf6MLOVl2dckrQlqfIXn4ck30RXa1L9QcrEQI9n+vY+
jS3qPo4oLvDZQ45MX5vWCd6+PIr7mOiw+BrmCrvS4+ywWcWoreghvETD0PNjFxmH
AQVRBm6NVEkuv/ZN54HiS6G4u5koNR/2ByHGT5Q333LTnQOKpaVZOFJg1o+FP+tg
B0ooQFhEQWpRcAmbuvbNv30aZozqTmYNyqQ/kz9ZkuaE6EkLBKsTpneaPjNu51g9
DAI+B68XyUQS4tOjk40/FRsK7o9usrzHzoCQTyIOk5fcLAJiAKE4TzMYVIbVqV7Y
50aJudjV2+OvNR3KLSByJau2QdrSjgPrKgNFMHaOSKaJ1btiqRDsdUvki/LZyanc
a/bKMGeMbRgj87gILifqN57IBqrqwGCTy0/CTrGD529XyFC8kJrINPi4HDmFYPL1
6Cioyqlp/uqQ9r6CLk+S0ZByu0WBfKaws3LXu5evSHro3LqJ5YlR0hOgWjGSdXI3
12cwdQ+u2hM/YW4FXUiPdVb5kUjJr3yhEskGSuFSUIYx584UahOtJJ5bpxtqUaIX
5yBy0vtvtHvLoqbSBlt3xe0tjV/CHGBeUDwOfmIkCt5GF2iO8M3W8ulBp4tkyk2f
WRRVl1T1WwEEByPduh/LGidnIBwDpMT5yZfKUUa8IrNukkK6+3gf2UtxcP9tQT/3
CwmUjQ5uYV7nbtkRHkolp/5TvRaEmx0jOYLBmP1YunHQA7k2FO2RROWrLGsNbr7Y
wVHxFP90V1CHwGt6DGLdWSG86ES+OvQVcoSEonjEs2ICQP3G5M2PQ/AgzC6Xo5Cp
rTfmA66Juxb1kAE+smHUrE/Njlf1YB7scuHym3Wt941xUXmpgqL8Z+/N+TWup/J+
ZlI8YU+nSZpQpDiuqgxTZitgbrKTT2iN4QSV9aNkp871uaKTGcoH99pRTR6m4N5H
UXAY6o5Nw37c7mxgxrAJIMW4UP+hnB69DE512G8LiiZYOCdGdlZ/nmctkf/N44+H
r+apiRi4MN1QHzHqma1nMZ8flpfK5X1KY8EgStJUPC0s6pc43JB4lNgrKvsVo4CR
zzmQcif7Jzn8tuqBJeUwlfRjt/2pX8D0xCqn7+vL72NglMJ/s8p57qF0hY9VXwvX
x/Iw5YN92H6/IGKTOrSV+05ATg/HmL06NFtpQLF6ukbYdoAHTaBhgLdWaE1bObhT
l0NIsH2CP2l4rvmibl+zUz0UjDbzr9W1JPI4rS6h82WGXPfVDVUP0TF8GfldqRER
+2LuhfOxBUk+gcteN/8EPPz8hwHSNZ+6oQgrCLew842mL15Lb4ZmB3pP/A7bMbV/
G6YsodOC0xEuHx838kbvPRHel7MfYDUVMbwn7lfENiiS3q/DplLG00YUMeECJRJI
tAJK1YY7cL6dcEHXdF6ZbcHyMyBoCQyrejamTUcuy4DMwD5xl3EQhHuzfh/M2SP4
AXKtdwIf1X4M9k5PogEF51RSys3ScmAEdoui9jPLl0lDFlbN2Geox45vh5PG0cXx
J69bYetMHkpyskluL2Rsfw09gYe5UsczZljIOkCIWp8JCm5544j5X630GTcnFBDM
JjNiTzjJXvbwUSoJMYgPhyj23IU4zADweG2zTbPzB10ISNi+6hxtyGr/BXhegvDh
+AHbzfIDA1xRvPlYEK9D2Q==
`protect END_PROTECTED
