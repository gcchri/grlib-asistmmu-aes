`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6nj5kpf5GFu7vr3N7Me5s77jd+BoSSeUbFceXlhVEg1kBt1kCVNWvySL3uxDYiVo
QNtYgvqtrZTBPvgr6EZ1rDVNcW2cOhSw0CaVqOv2tMz5uZDyF//zQ0TuDO0Gv0SD
uav3QwgeDbSmi1lAj9ymPpgQF5YIZM6bOkup6msdIGuDe5sIJTHU51V4Y+dy45Az
wKp0PY2rX0080/f6s3cIod7owB5TxIgjKnALCuHaps2KY2nJL1oW3YE53oCt2S1K
HMtOM/WfQgYuLLb+qyFB97ySMko0Rs8da4bRn4vTqpSwXKwLTuTsmGzqI5B3fZcr
k4xBbj3pV5YlsjGgK17P6tGgVT37yiVD0vAvwH1oyfja/sHc5zmCV/MbLk5ugZ/X
h+ikLVDku35rEMX/pNP79JFqjvWmS+qiZJVqnqg42e19wbqAsNh0FLgFoP/O/sXn
GDLECIqI2QdToSfncPgugACjtdh9vzFyGm+ObrfOkcn8wAURNhG5eD9wwKyP1oWS
YVpZ9G9n1lVzNeR2ujXgQYAAtJRMwao+ntRcN79btLNXocAvfHJY0dZ/wDZ7Asew
qXBQzkmyvxLvxvBCxbGSZQB9I8Un4wZocO/vOjsRtyKi6mfI1qM7U4wXWXDpErx8
eBEt98wDVb2N0TffbFeej6h5MkU6lUellwidIENuxuY01b1Fzhp3Fq7ZH1KJYG3N
RHIn9Nun0ODdoT/AywAhGLm48nmHdz6OrUZGI3TkNacyd27RMtVeUHx+dSavGQFk
`protect END_PROTECTED
