`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ifr8llw3XU3cZr3V+nA+d8bASLnnsL8RPAPt3ob/RQjkApawG82w7QxHJ4gAWpzr
wi4cXTYflR2KhMTxtikpbKcXQalDBEsPE+/0OIGQ+qcGELWVLBqPLyQcqYZ3KVhX
qW8nkg+CTnXEdYVrlkrNlgwwls3oclJVHyi12ZVlDFcx+eHR8ca7uNtmhTgyxvYF
dXdB7My11+B4BHHFsFoLfxCMBLMOX730rvc9R69+4nTLV5h+p6y0GAiyscXmplcb
qOuB1Jd7zVO7UmdzKGOzWw==
`protect END_PROTECTED
