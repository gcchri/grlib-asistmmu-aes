`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v/K7acVh6FOPvy/EhLXp92C7sZDjwHkRvxhuTLXmJlgrfwDYE1fFRCm3VDVvZR/q
pL5HGqltTikHObU1ODlMEyUBqRgJ5qFg4Kyz0V5Y0rf4ibUft7pIhWxQqkitRMlh
NR036d6/pqoP4Ag1UbyZPKsmE9LBe8RKuFbu93uSrwPCFhxFhPre6nJx7EH3Itbr
pVRUPHI/Iyk2OcRtrizRZ4kyez6kIFi09Tk8dH4vb5fD0NwbB2yfW2HVBLSQHk8A
yRmIRs9TWIfb36muXJtwaNEdU/6zBqQMSFrL2Ujg0280em7KIBHid+pZLEfI9STO
isYOKZSTOd/+eWOFveAxuH5fnsPClYVjRm2g6BRWzW6qmVyMDIMSc8DxigORN/Gx
I3vuYKYSYg6hayBrQ3L7DTvk1GgUyh4XbiPXCDCB1quesON2WUptoqPbs1dxui7w
rxy23QXEWUFFSt9d+QQ5hOokZcVE6OatmI0PslCnZrhG5RBdNl+1R3iWe0R7l/un
9x4he5VqwaMKcMGh9kpR/K6qvXWdtVbDAUdAKmxg54uYfd3YVCaVmB4pt1S3zPiK
D3oJY3uV682woyrf1tGJcRQHMb2soMVeOMdf97AFzcEDg2Sr/ehWT/GTwEBEFyPg
vQGQMzd2974PhqjdyjA80SlNxSqW8s3r75a7CqMkiMqZEtoz+OtY5Dkx6eRCMoIL
uKQyp7dWK42l2sA6JKflhyUmzuqu7F0shG2vHZcLLzh4qH3bYuFcK5/R1XPMV7Zv
tZgPdOHYLj5Octi7GncesgL+A95WSp1OCb0hIjDDhgtUWVVKDOgsp/NkxlvqHClu
0a3zTmmbWI8lQeBhS4y/jJADEUbMC/I16SpuXSQf226edYaAwfgt9H3w25pGeeZC
1e55ZfoStXypdjIF6/Ob1+m/S6Hg4EuDCcVn0fukvreCQw+TyLFWTB4+jhg0bp8Q
a4w8GqkrO9DyejguY83ifUJG2xkVPMRUTvIZBNDTXyVeGTDtZC3SSiKzXMSSl56r
9JHJD7HZ6A4XTlDFmsHKP9tK7RG4vEM8Qvb+qcseY7wTbLd4CzPf2/v21cVAVkfU
X+E7aeAqj4ft8O+g2r3FIVus60O8O0cfOCAC1t5uXq6HS6uV5qEMkrAiqmVQaWmR
Hi+5s6gS6+xjsN7yqNLBwf/tmFN3C+70+XDEstVnrKju0VoZ2EJuiixM+fGLhRgn
jB+uSgInGJ9mspRga59eA8qNmaYYibWkpJiLUDOva/QVdkuh+Y/qY+B68Y9ZI2k5
UOLxyMYLO3004utPoYBtA9WubAIFhGl5+XLvSy/D2i/8JqU6sn10Xb+EHQwZak8r
y/Xbuzx0xlr73Vlr6F3JlsrkAaMcu+cHxzQIETzX0ZGc8qtAvqxSLSSQGrx8da0T
7MVi6pvas/WSJ8pfQA1boXKiV4YQQ6oE+YbitUM5KNHEmzNplbKF2Bk+6j2PPNwV
thBow7XE7p5WmJmkTstdFce6stGzT78/NFvhnO9W3FYVXskuUd/9DSi/QM4XTu7s
6CXquzP6C/JvjXR3N/Oko8RiqEAoSGslyfrna8VDXF7nKCh6yeQskTZuv5aB7tNL
0y4KJmni9+zWEHGmbJ+UheOU8cdVET07sJdJNjjMwLgGpd4OAqeN+x6d/SNxaXg4
lRtPGge4JGr7kmycJDa1N9LWYaaJTgaCyqzMfqiR4iC7tBmT+iF1tzyLCR6LNQCB
seddrYbV78OQ4rnSXFftWXpfZF3EAAMuUs6uDt7a/VAtgSXN7kubfAQcRDGqnhp4
EN75qW3gOIfBQUJajaFIJyQxu96UL0Fl1x310VP2/hkK6peCxVkDih8pBLaBjGLF
LkZKHfMEPZcI8l6EZ8iwDmpEL92mVAQKCQoLsBd/5Sgg5ZNh+5CqQM79n/ha9+bB
25fvQomO50VGnbPDz4eoNr1kYKNs0x7+i6YQrA2dm10ztnDtgkSGm0xqNdCHtjIW
vuhu/j+1/ZfE1n3KHSohF/HXWy9vNo4ivWeE8hi38/xnQo4QxS2zsxq0gPVZKxNN
UwgutJx58TNqhnYtjLP+VlXcJcmUrS+ye4XW2wWthrFxYtLPAp6PbQlh98FlcYFv
NO53DZy0FqXRQT1iOo3MUEed9yZ1OA98m33VWPlDiG0VNcHHUKIaz0OQXYSrTXio
UKgRf0KrrJEcL4wnkSXK1m48tk/9qelAmRAJHFrj5MgscLq4y7LUYvIOAryrsZRB
6clBhIJFrX+f9OOHi27y0JoG2EZLuX2g/dQA9KE+t5zY6e6D98LRQvsDTu4wUzNg
ErBR2/4baLgbMpuglAwQcX8BluOqS4vOnRfCtDLinQwWz8I0JCFL29yfIJI7mA5i
BR+tojqGehLgetyC3W5YivWcBlhSGh81mhPleUr9UxMr3LERz/vV1vls83FZz3VQ
xGd2S89gE0ivaUOnHdYZTx5zgzkaWpCCUP1KQT+ZHW/ioNcmSYd1YSuq08iAzqmF
nvaIaw3Kb4SHs1CfkQqJpzZJ+jyChqcz1x1bSmGGp58dsUem/AM1o6haaSS+s5Sl
57q7bKdbkhikch6XV/xl8XPVmGXgmx9hZvIBiCxBdmygvEw7/H4wLD5rgk39Mi1V
+BVBpQ/3cT6TBbXTAGjYKbwCiuIOIHeeof5MbPAq1EKNHs0snh5g6M/7GYTRnX92
nrPjt74ZS7gHiNXXbx4cto4mw8sDau1/P6zsrjbpEygEaqlrTCy7fSKNJ2Xq65bQ
aukObF+LxIrWdCopNXl+awflioeKiARYBYJjfC8hkGgGwQWfMxZPV1W4AQyfZEjn
/r+ONg1NMcBUx/aX/FbxqlUm8Dz4yW+wWRhFeO4bUP8FufA1BIseHKOElSwV8GIO
Y+TYSK6F6cTk1PF4M6UPLHacVC8h+hFjMeBcF3ct2+oA+1jtpqEnhzih82RvFka5
B6X8UhstlsH8ErgB03Fq+Tl9LjQFo8j3VvZ6M2lf2zRmiFWvotbikxhXNXcSRkzE
Wv+9K164LGtu/ZDw1Agf6wx1p5N2S38R1roVJXxhYUkNwRPAlM7cAH8MEfzCdAet
4avPJti9EarHGu0AxBGya3Nd+ywdolRcsu1n+VZGI+sT/CVhj0DACfuvIcow4YQz
yAOEaVeclfCmqbst7dSqTLrRtEoKkQx8wBsbABgZR1rGjNodSCFQtW1D8y+R5Xyg
33jmirYXg05KFH4pPzkkFhWm/5C6SZNbGufmtJNN5/aO5TLUYL/KjMPX+yn/v++I
EnGOGXhYF6TahWJh+LS6av5R71/Qi2JAYun7ZBzwfSxk+CzK4tfKRAf6Rq5mF/5A
Y9Sv0XS/F+mGur0hcgnQWaeDIWfPUaJbmQ3N4phNtpNWqdX2BG09nFmmLL+0CM4A
Ul+9UpscTh4B7+GmdhFAcoFFQgOtb8L/oZ3IL8LW0OGsq83n+YJ1lTIVWW5oB9g6
Q1ZcM+LSss8vnN5FmqSqZVRZahMqeo/jcFpED0SjwAP0BS4fzCUQthk7XAOt+qbI
fc9s02gij60v/zNhvPKIPhrBv5uLgBa45N8jrfX5LgoZduLddvdpE08nPonIyTHA
4FxhQhHrWXJuIilMyEYSfmh0CM3sqBK6rW1hWY300WjJBqUOZxCGd0U9ieCOloOj
LNH6+s4cQaoMsGRNt2eGcF36Z0qbWMUCnfgKm2YmYylriu5M0NgYkw0eXppIWrhA
jhGU3Qgh4KV6geed4U4mhOYXCxqjwbwqh1W9F9gSvHkYJY85SkuYkHM66Yoe9YAx
evFK6V9luecv6K8hsSghPN/CO5OfHeXe3u+BQYtXw7ZH5VNUuVp8JdXYveRZmlNx
KDjdTzx+dcigJLgPIw7m35NCX7hlgkzT4Jt/OOeG9Xx1iBJng5CLFLOBG6fYeJLC
g4S8IBJVEtzwxjBEJ5zKDxJRqKmT9t8NwPxvl/a8KlqyX/3hDce5MpK4HIGFfMm3
OVxQtUqSw1KBXX3C0wZ8KI1/IuHxp4akQWw02iOt/WSWKGVjBANqhE7PNCn15/b9
6jOz6pnT+qM9+2BxVS8ilDRfzpLT9iBGM4XZQ6pqtcz6eUlwNMbemVsTNdixTz9f
wzZMG7u8+qtIRf4jlLaBp826CGUU5cMJRTE7LOJixlTQngBjtRm2Julendps4hn2
Nu8djvqsa7ZULJz6vdEpcQUgUp2p/Z6F8zGZ2tI8cTqzRlZ19/QnTpe/PCyLr2Jy
D0d/oYxwv8jP8w7rxb0Xs8aPF9pCo/PXcHfYqauu52XmCDNc164aWRSgdBcTKRIQ
0dbFzz3CT1zQiU9Ey1rRrxNFetJ4jG+ivaNcYEoaodSRCaivBUocVdGGp+3Sfk2X
sG2trKLBqcF6j6R0tgVhTArmNrMWKP9RTDmX14HKRqDyHsNNeGeFo6kaF2ulkn/a
LIPqMg3bUyv1O9y599kC7Hx+edlyF9XIk6SPeHG7vF+gZKq9d/GDhEkNLkZbjbbn
E5SqpDQtMyDg6tyFEbAQEtONaW+P66JSdX6frVvqC39DfHj7LrTxJJ4zgXtCp7Yj
F+NFvlM5zgLyfOFTMSlOOX/WGAWPcX3xJhi15X+7mebXm+z9CT4y31ggNKIzoB3A
LAPN6RWjsB5xYm1F0savxyaaVQ96SECAqRnqiAIuFqtxAEu2gYmfdNDW2qmzNwSF
5PPun9HvCeqE4aOXr2nJHKEBubk4uGqZ4I0m1RhtSVCe1l5vKplebOqFNnU5ow6n
qz5CMzYlnafWCtRr3/lbQiimcPGm/lyq2QryYz8OUSKKJa7XCvFR5wMv8ne1lpD8
4zX8C2IM8viysKdBs4c1476glHz/y1ehtjYc18rXqiKzdOjWfRUnpENkgQc60XHH
eaMyWfv1MhoT68hQH37fwC7oCaQrbJvhivciM5uGcvTDdp7GRRvDGVmg933X5ND/
LDQrixMMGRStWV5D9ddvXO64odQkfCgpEqL0IUX/WM++b8SWW9RK48zKCaoRM8zu
`protect END_PROTECTED
