`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+fSfhFgZ7FKmartgubTSlVrP+sH5K6wNCMdDgIQAm2Tk8b1kUNNRJsRGsUR3SlMQ
99T0u9tuT2xQbHOJiGGxecbKdt12C+fYuROmHWLC5sRtde2icNwc3HfRDpXTSYNp
CmD3Fgf82grEmDl5PRweLdW9wU4t4BSfS5Df4Im1vhuPu9W4TQhuhrrF9bYbH/gI
HYqJPU7TzSpew/z10VV3mb6ImMPiV3U8ybTwu3gBa1cPTFJTjL8wUv6L6T61+5w9
6ClQDAOML5JiDMZJSScHNIDzvemlayJvmSvRsVwrkmAKVE+A+1L3vYUH+ArxPtJW
hnFc+q9YW8aIQKVzEPM+VEb5F+me1K8UHhGRHWD2mV9Vj/1J7K480nkJ5z2znVTl
JjSQjfrTe2Rp4soSCnjKY3QRcJCGzlvN4GPahOFUc0NPrcVkum1/KCWLksCLMNL6
V+ILJAJt8e+0WrDlVEFKD5mHF8768FOZpokT0pA4k+yQgu9gfdgzMwdx2QPrOI5h
/F/Zgtx3lgIfO5F4Bm+r+qaFLysUPTt3kZt8A2VZuuPa9Icx4D40j90CocWblZD2
nBG4wsuYd1pA9CQXasFnYs0kGn8Lz00vydYEDNYl/51iKiy/0/XB3tdPoygcKf3Y
FhQWWTmF8ub18XvMW+SC/Uw2SW+t0Rdhp7UD2Njg6p1SOnGyDk4qkDvfAQR2j/No
jeUjjed1eaUkE4UnDjsNufzooVdX1W3jNp5YLnsTaMFYvIiQCBKwJj3W/ztqin4a
R2jV5AxhLF9s0oOpl5l+W43zUwBu/0Gc7oeCN/HrA4KFH4700Ah9IFt43l0zcjG5
QaozxHr2aiU2urKYPU4Z+JP/yFh2KoxMmo4tnn5VktyXDPE6USPGQtXVVZUlBnMi
6q0ISF+1Bmas6xTC6yNQ8YqGrvA3RcfmLJPW5kWHdfvS+b8vzdpBYYZFAVVaj+TW
zjYB8vB01P6MdEUwExkpvKMCm+c6IaCuZYdLA64DH5EPVVK0RURNtRd18Uepu1/P
jaLGg6xX4CQePLQZFQBCXKnfpVU+m8RBVwcaXgGNiPY5WC03gaG2ifDDTD5G95yD
UsqTuE3IAD7CcA/pTkip/FE3DWmTwE5/4Bh4zVOgA4DhSFulZYxspCJgocp/uoDP
CdezpwxJDWEsdrWnqksczsPJFjQQk3DUx9cYHjm7xoOUkkAsdy3daB10Vxw8SDao
sydL3+PR7usdh/QFYiXnQg38o8yvrlqt/EqL4i3AhzP5QuWhD1/4zmKMalfAUm5J
p8xIKEgd7zUeW35FliKqcjPHkle5JILW6qUP+fbfHwg5yG6Xr5Wc3DltlTyZ9VZY
9n6doRmodbvOcKeWEpk2VEq8TWRWhzzjR+yLGVah1/keYgLsHoCRjIWSQTjkvdrF
7fy6Oxbd6h4xge9V/FnHdnCbRUXwM8eM76W/SeIEQ+ld/JKM4b1J9pAfLVu4EkpV
tqQy30qGG7rXQPJAIZWWifqy1Y3PJWqccu54avzjzjRsmuPxLcMrLtOXSmk05Up1
s2/k1p27fkSHRsb/kFpSvwx0A9z74W24gHoAOXg3kbpOAPKqUgX2zxCRu03E8JYz
NNyl6qjkSMq7l57bzc4IuNwBP+IcgQHg1dySHNWI20UexbtC+q2nGYPpHIgYzm0C
9DkLGwCxsdNLTHCQqBVvoiM+OtcRUzP+51AuwQhajrqy9aDvk64lAASH12hMdSGP
Ys1XPOOQWPAOIVAAArltoQOvHWbGoTSzw9/m3A9hqICI3oPsvK+4gGPvH28AFJTS
Ikv3Z6zKaUPNHz1gpSfNs1j+QXgtUwjYU4sib97opctC4PMzsJ4gddfuqZ95847/
G62XD4OnFsXUiz5cD1QFyM/82yffr5xOE+RDBm+jaO0KoyECFLYtu3FXUJvkMh+g
XzjLXRKpbSi4VYMF098qWGdZvlzRk962lsz/+iZ/DMDeuK+4ArqFg88GG1SsHZoN
UcrjC5Ss9exktT5dn6IGAWUWLFSSfafK/UVrwi0r45S47UJepy5Y1thjecy35HEd
rsHvAxIRdgZ6rr3YKeYfiVqeEJAuoC0D1DIMz91drog0pgJ+a5OQTeADeuZtX51X
OUr+c7C7Tf+uDSPXVby84KFDq5kUkMisJlKT71z2iH/P4N5zrHaUKdocIwmudSxg
L9+8o7aHDYOKJ/uEgWSE6tZqJiqIVh6+jZS/6MemceaTbeNGdjXkJLx09u+8Qp/T
NeH502OBuekI6vgX3vBfHNC9WXt02ZHNGmVaP6A1DXb0fgeWovomw/JWXw6IGBGG
E9vegV+T0QlavyQFWqjvf6OVZg6O4mv2zqTIa+mhpZNqZJhPC49ulS8/MKXnnqLU
512bDUGaUIeNGSaLIxVYb2Z52cHnohdlEJiWxSMTyzYPwMSAgGumd6UQP6Nrj0Jm
xQy5uyQoTK+RW8D5z2PCb1AcfoRMqozqBM4lJKDyeBvE8n+ka9CJUAjmlK3mDLix
DURa9C6mlUn1xN+qXVsKduhPHYF8W1AmZtovQDMAVskDN/CxiWlK8oHqxy2v2u76
QRKVma6jVMtS1DtDRYGM5RwWEVLzSVEIYh4NnWPaVnRHtSoMOqqF+lOH0GG4LdBF
Vvwd93aD4+BynmaWT/10FDp01WPNImbvs0Jthk46cRBDRaiuyxlAwBy3E2tmZlrA
99FeYsNK352V4Y+bgUNUm96wDFHazaU84yI4ICzfUg0ZAQYEcfjAauYf7490Ox7X
hpwwTNK22upV3ASODf+RKeBl3KIh5nC686/EmyRbk0RkGvhr7R9W7a2Kc9fsxU9u
qWrO8Xi8vkmnicjuPdgakXgPksiJgxGFKSoSLwEnpOitBlrA4BH9qp+cAkMiCiM/
6FE7vDWQL8Q+eOQH8LBMoMhd6+x+MFHPwVUgYgr40P9yneMZHdPfpuglsvYH1qC+
dNnKYcYEqTweGVi44my5ZINfD2B/9Y6xtdhlGC0quUU5wfgPONxekqnWDk+NRS/l
xS3IPC86QzLDlorTbmUmF4z6svOv90EDWwHgUMMNozaLg1xK9wzjg2YPvDayOhxT
XTJ08yPapr5i4If4YZrVlRDaD8n8+TRHKJUoteUni7f2BYtDq9b28606RuyP69tx
m2v28V6RbGlT2foAhPER+Pzor2IHUtrIvHfB14lEq6Wf0Gn5BaHm5B1fhS9NTYlr
JNdmZXFesJZJJC0+OI2jCJAMbLkmqMmDso9FbxLJKnx1Lq7x6IwsRCJrg2nVAMfT
RSK6YJDcVukrdomk6l0tGLnhKDCnvi10RcDat1HaDdfXj0WL/4lPAX6fLXduyGHV
k2hA5R7mCbIM+f9wm4KGbJ0gRWi+zFPFqnzmd0b04ejOSjhyK49zWvb9UU7slH+R
VzHWfmZ2Jwe9b43XMKyig/wVCqsC/igIbnN586HF0v+5rN5qgb0YAcQ2k9zqHDh6
R8CDyT2bukDb4eTp56EEGS5r+CaRbYu40BCuCHMH0+adRCNKH/2tmI38s1I6g5vq
xjtnlH8trocaSscfTiSm5nGIuMP56bFzGJnQpjM7jHZBSDUJqkt6DQfJbVOSEhDS
MgJO/+gVkXzNHwTy39EW1Q==
`protect END_PROTECTED
