`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ta8MVtuPeNG1Ur3KleKMY8I+N0S0z8wsMMknk8la1GODXZw93hZ6Y2eua+tKmhAD
SrsxIP4zphbW668DnHZe104JZj0rdsUJ8m3szDvkiDR+HUNy0tZBzFd4NlLqnOJN
R20vvGSZL6PmFyUpLQvOQgvKAyIGqwa3nDzbCh0wPERXv+K45vgvMMxSZrCf4qni
aktMZm5sbPFPWPZ/q0m/ZmdqS93por7HKuMQDeM1qLlHZJ3xxkHpB9YVbODKLokK
ibvpI2f0aWdQOQJRY7cGoTEHqioc1ZJtrPJSosByCNRFQW0P8pqFNvAA6KQCE5eq
fWp91w5/I6icHvbo+pGSDOm9OlVCXN8JlYaGmzIE+urgDkPBvam0wpRAUcr/V3kd
atYfOcE2LpcZ5Xk37E8o2sVDYNkXKbxM8zMwI80x96asAjGpfgYTUo4S9VP2vq/j
KcPo/sYlTPQpRG3nxW2v5MUv03zyLLctQuWEonQ7vlwWde3j37l875ZytuVMNdGv
2BLEXjleOymrVwRFfdFAG0epgcO3SV2qfLz4h+kCetoxQoUwFrzVBQE9nJlxos6T
jORF3lkOx6uUFM08XVIeAmebq4Rt3Vl2kDlSnFVeL6dIiukRykzpoXHYff5Rq6FE
4CwIEPFpgQtY/v4P26d15nt5GK1RsXVKlHzEudSiMA/kq9XGHoYJDlV75/MzJ9KP
ZbLIoCRvWGnkpLYm9VTX0tdvAe4vyrw3IJ5E9k6J0khA4mxaRC41taVGpoZN4KZ3
+RGRC93AjwmpULcuqgByqbSeBcF0GoB7mnQTMnppnJf2c/no8X1Vu/2cU38uJVVz
dobHHkTCXX8gYNEuBxJUTDZdM/eRduXPtRU2GwWDQdNMqqaHsi22PUp7jPaJupFu
73JaqGYWNxW0326eFn8RtZLx5S04C5CLDYsurVMCBM61i9jez0EtjmsXlQ2r7z51
7K6gcqrFeZGZqbqRB/sOfhACmgVfvZoyPbVESL7emQ2yYIXQGnY/vn8BecrjvhvU
dADGiHM3JwtEVpG+STvRCGgIH5yoiQWpmbGNF9FwHXx5mtC/F0Fm2+Wj+afaAipP
OyApY0rhj8BuyOV65hUpGGSzXAkzWIp2NdigNp2Pl+y1Rz3o1VTSDfypBTqVqFoj
jsq5qN8pd/b9lZ9/BJH+VAAX9tTvOlM2yrQw6nHT4RU0BTHO4uGTjJTZwSsqGamG
uKpqrVIWhzEBTJAgjnWI9SirYT8mkW1ijzMPHY+ZZDUXm7l97jvbnjlGbcTIvws9
p9J86zAJ1m3EAzADZ8PJFU60wXoi4DNP926JAut9IB3bVPVaAMaF5Jyd8sZBweAy
99xMth8KsH4GNWhso2k77rm0Az5mmqM1fT5roC09y6IPlV9TsfZTwdSQA5KPHHL+
maecT0VrStubwaBpYtOCoRb9K/7esrI+w7GAP3n40IVxUOjx2aToJrtW3W3eWb5R
XXE7KIBIfslRneXqd/79KEtlLlHjpZg7pSDOwSPDdj7+csvKNy/e1+mCCdTgIWru
IW5Dt6c2quKM7g7Rc1wKUadxZS0y0nJw/Rcjr30HkeduedSzJ55mJSxbnzvKIWgr
6q+QtHn9TagLoJu0O0UMj+Z+6olQWMKykjDcqGRnlKXVSzN5Lo2onrZZ+eHBu+K9
cz6lBepDwxJDMBFv5srs1mY+jeWmuAlUjMqLCGepCGcf3cLH0x/O8qDAQfw4G3uV
FRrrvHLWDisuoJqJuc7BnWS5kTWQmyScOnfCEzbddCOmGzAe3ku8WMPvYNiQH/UX
kYZoG2lv3NVIQj8lKXGmWDZ5DRYgu09C1mML/0a4OE569Df7h7TyhUlUe5dUziMG
OfL+yFxzcSnFxjA0qmCu4TP+ilAGjQGNYTSCDBD6Res3jUlUSqlLapmAu462843l
SJGRFBPldHGTU5snKCO20/ygTSM98YoXzkYvrR/7z+Reh7lC1lMXcU1c2jFWjBJb
QwO38FuB1t7DI4h3CT44YPl/69TqbuNe8bAXwovDATgul/cy0VSs7K59z5I0Cqre
A+yCKc5+R7MHFOfKxAU7Tp1JgvJBx8VWT4mlonvGjAwdynDro1adnp+wSR/Eu79K
zNsxtA5Ijx/531whzN1fF5wRxf6mW1jkpIEEqBN3gZgFyqpKdbj6duWB6Pk29wff
`protect END_PROTECTED
