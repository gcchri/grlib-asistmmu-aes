`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SjzBllySZlHYBPQu8NkNf9MiSPOnPfycSyGSp630kkeKmTNaGxCZhM/nuQrQ2An/
hz7timo73+NW1L8XUmvTv0CRUuvSKNPtzaE4OacbJnBIZ2SMihmicpqy7EHL9ZD9
akg7dIZNg6csNkkPneLRLOWORjphtvz8Z4UE1ecr+G4NFLkg1mm/cz/jElw7xosl
aYNGL7CQdri2NXYdi2jehDghhjh8J2fZ7LOAeqd7eGpJeCv8Ar+fjK/K0/jG+JE7
NiC51x5SWrfkFYAMisn6/jBXj+KVkpeHPOXcLlF3x1dbvEn49+eOdB+uloVlrG39
9oXVgcoeuosaLG3Y4KkNjW5ncpki2/nM9gy4kbn0FUUu61Q6DDy7ldntwpznl7fJ
Ui6xr6nenLujNHyag/zMR5SYBuUQ7BMSUjIfOcURIIRuOzAJb6Jux9mDxElLkJD8
KPMaHt0ICzEs73TLtQLOy9l6+OIo4Jeb48K4NIp9PSOcLX6uSMcHHc9hxn+tEes7
CiUeAUbkvjPMiN7mC718CohYQrSHO2TFYRAR/DZ8PssEt8D1At0mq4Q/ffwLLGUf
6yqde/Yg4NFgKVljPc4/+B9FcpCAnvlj6ifUKkvfaPomD6hwptMZdU9ENEANlZcc
hmXgx4wC81SLTOQPt5rKP96ZMdjnSmDWnDeK8LZZS46/u0q47Qzt0L9/sbQohkHD
1B/FjUX/TjhG5QhNFkg9xnczkwp7BP/BzWsZIc/1wgvuvw1Yq7ZxLXE6idM4OfAC
MyvTaM14XFrbSrQxhS/Nd55OMRShexa4oIz2qglpg07lXgTc68/dbPkPUykK++f3
EtRNOzKxZfNZfqv6xUYm7lxkCORtQWy6Xmc0TvUpzrVkrvPkpkbEZE2m8UhOLyj4
lB31al0HAK0pAx0vHecT1ugqZ5fi/KVc76rZ5bCoEXMotdf18Nuh5HvT2hkWDZgf
7jB9bAI7be3+fmOhnLhrJonzlx0VUG6qJnSFipVFqhniLTyRx0ftyKn+Q4sPBTbf
1AUVY0lY0C4b/VkY6D1CDCxo+5+P1PwC4BYuisCJ4VjL8JUWcZg/bwOJYr4OFU8U
TAQUsSjxXJJ8G7GGqYAfPX15MmxM3LKNmg8onryaBeCwzd4LV18CAacX3WyP3gPx
gjm2gLLqLleIoBBkPReY0z91G6SBChwVB/jMmB82JuJe9JxTZNfx8U0e1B7BSnW3
cyxYgWBPH1Qr6eTm8ht6gHdpVNz52gPW5EaXZx380f+2Y2jXCklNy3NEiqm/B47E
KR2tW7es9WbvxBTRPXrToU0Iiu8PbK2RNvJGawHUj2lzD9o6c8iwfBY4EeiN2bCi
Yuc78+UQ4LEMoPOy1QJUU7sXnne9Qpg5sysglZUR8oHwmWwrhpbaTrsn/hpoiQ76
tt2xn2tvEW/jwGgKa5Z4SHEG0poJ0RkWBXWthZs3QiWBhgb6P03l5ob6R0VN1ORy
NdC6VjjM5t7HNYSnJHxWsT+YSMNeDd+NURLZNWmFDQQpzSpp1jTn7ZN31cm+e6Rs
evIRW8ktNwJOHnXHVZAzCTIQdfrhcmSNyGgmiU0/Eqnma63HA8Otk1WRKryarrOX
JYrM0L58G5FJ8i9twbobEXl68jlWH627N295HvYIrqWR8rgTNlbQ9OWdzgOMlLos
Bp/j4/wbDxY1JDpAUANi5oaZSKyXCzGGVUl7XliERRyJ8xFZZ9njwpn3WH0AIEGv
OfCMGRxQP+2hlVuvOK09/PZ14LlV5Hb9q9iYXzPTWkyeU+rW0573018U4Xk+Vam1
d3OEuhLn560AlVYWCISCaYLaB9f8jgDER9WWey/hlJ7lkJywuYexO/Ed7VIpgXy5
FPrwdJnfceOcA83M837W0OhMY66DpPBFH/v3sgCMiaZc2eyFgkzWCv3C1VIzKxcs
zEk9gq7Hkc9SzsV/fwfQ98kOw3NaNR2AOjDVI924HIqZ+jtded7bSs/kaV9dA8w4
HaZG2aV96YDMfe0JL3lYsQHqtu/4YyN1Pxxk2ECMNEseVOJvHz8tKCweJdJjCyFi
3p1LTUPJ7PWUvWSuimw3/tSUiwMlFJfO2QwEURbR635JRwtGAY1I6MGrrlm68kld
2j24ZYN/6xzv4hyFwUCri8BPw3uRvcF5LM2OLsSXr8kiyGsCVDnmkzNCT3IOcl4M
kpdCWOHed3ZfC+FvT+zWAdQlqCOCXXC/IJbehsPdS4RII1+shyilExtuKh2bLWAs
TO17TkioSFGpcxbi/SqBiOVgwS38IBbVoeACY49QuxOwhYDXJ0eIzUHaQgzBOk3R
y5lm1qApgklwLDBOBL4FXlCFzjxRSZeDkTHnksCRJe4xHdD2AGHVXkyguUtrMeIV
lUU/1iK4c9wwzoR9dY+lCiI3rPKaxpokEmYRa/Tu8+Va7lWswXbnN6g0FTj9AYlN
DkGuUISekddn1u9gR1XUaS58puAx1kFMfxQc4lDXAxNxc+2l68Cp/MTKgPkXWiFI
5yVrJ9QbELwg5S+c3dHJFJaIXUZYgQY4XtUSE1S51vq5BiD9mEWMYwK9wiYk3YqA
EkoqIDI0rjXeeth7agSjZmRwb1xUKoIfN9qROsLy4DOYvZKxoLkI2XgIS/Iz4vqt
X3dwQoyIJ67Hl0R94U+eje56JWEo9GdjSO0v+ieaE7a2WTRKSKClSZLy2zD0g/ep
XAm+Y6vOFg8Hir8ECG1oovP7BLxOM8Yta/6H1CNOnmmj7re6JDuXL56Dn7eJNEKu
rJ0gjW8xCg/XUjapV6JYUiD+R+s0ZUPcez5XXzYjj+7Xqm+9SPdB9eRfus0Eo8Jx
I5MGWL2cew2QmjE+xYUC/VoEx/R/NDR20DrNl9AD2ziwjVWRgHfowKYsIFVX/Lf4
GHqef27sCqJEFR3i+OOkdgkOY2Z+DfkNddBtG4j2i69fSc3RSFJyXGKY6OvHofN9
6L5FOy8AM8ZPU3KXv3l6iDBztYxX4aQtLyZBCQfR7bcKs5NSSM25wVOFV9XKjWuD
k/y5cFEGGf6Y+iWpWeL/LEKFjLjM+uwOxQXWAs7kOHBBoVVQmRV2uVzoH6gQ5wc0
+n0ciNDn4/aveujEO7XmnWz1sONIvJ4zk9IK0JQNp+By6IwitrqfwclMe0LyeVGX
JReenPhAcUEdkyq6SGCGJv1IIRiX+C5oAnLIbyXS1X0tPu/4tn35ggZxtn/PAhHe
S5WsUNyapfGgxWZwczTa9KXmq6JcDuxGrQ/kFpjXIPVpCneuO5M8RG3Ftzh0elCC
eVpS/MNW1qZx5VZsL2YTWzRLX9g74x4AuYbVDJk3UzsHoaESAYnl9DW0s2Z6dK+l
J869Y/wZId4CkPlfll4cpSmV0Pv/m5lNV9etmVFB7puO2LgBX5oYKXHDvZRM5fed
tprpYLN21R/vnnVs178R/cQYCNLIjq04eqMDznOcvr0z94EiVV40hdV2MupfhtFP
+dIqO/XNHNM9rEgjWic/Z2fz7fNmpCq/h3kIF9RW03VWpwL/sB3HmntemOGyy+P4
T5RqFhjKQXx9tVQFTOTyW/ZrhMUX86byKHZ7B/ogpHQPpSipdSbIbnP/gkrC3J2X
3vi9slgOjEoKRz9xKUvLj7w66WV3rdZNU908d9t2wudlj/CF1Ui6CVCvIMSEf3Xc
zItUFM5CtyCBi1FIL+Xh62LbVFVusTk04B7W4xiockEmUEcTYXZ7xcMs7QM2iQOk
rYoUwKuhUvvakFDSKdL08YlvN0X7VSvRaraig2NeGfeYc525M0epe4u7ckB0BCLF
IHz5zzrECYmnWRDSTWGPPOw3eqhpRcDVGsAR9uPO/hTn3zJyRIKTwyRcbtETjqiw
wTIRcxZ4czSqPJztURjZeQwYHKC86rLAAVDyQQaNW71AK+1PPfehQMo2r3Cr3fCd
L9vHsrfqcRkIKzxqmv/fm0W2+hu1Af9MLjVoTIu/sTmTkeBCWB7X8Ne9oajtj0rk
kqZLZ97fVDafXtSfXT7t/J8GGOwFVdns6Y7s85nfVX5HymSP7b8EJv8bTsdUg/YW
Z0rxOvQUE83ClwRaZAFH3RlMb1eHp5kkBz+dIuUJlVNz9aNdm3ooh2UjVoaU/UBe
WxeadDaP4aUeeVoXjFps5pUXm/1YUudOYtWZfl2PxSH2TB38pkysKVbrXHhULmnv
Pa6IE4RthlNwNjCT4ahsLQP0tvCSnGYECtGapCyM1s2E6hon4NkcnPH0M0SMVINY
zi74P9xDtAlXKQz3GV/cSMkT+3cca7H3JNUP2mR/HafRFn8gbXccAbGQpEIQaXuU
Jjkt7smfKevtJT0aMuR33xuFDbnoozUjwUnuaBgKbBqqha73XDzwLeNyA4775TpF
FHBiTVMLQwq0teTyr+ysRXfjDflkcUpCMN1ZDdLpTrlC+fAMy96g76Y1Uvzk/EYS
707EURkOdE2K7vjVeG5qWHhCntZlI79fGqNWTDw3d4fGVvqes9gH32F6h+pldZ6l
LmUJkRnZRsHIanXZZtcKVJXMWvDDOIGYho/lv/78/tSRDrDsLMvg/RPQBG+ACU7K
7sOI1cJlgKc8gRO9U9DfdREzdjxdIxSf0vK1E83TFBchgzh0Si+IG8XftFX0QkDm
zSRNX6dkQgMqVo0lSHzDP8X475LvKNkCWrkBzECPjHqMT5Bx/KqHa+na4noy4P3l
i34V58p93SEZQo5UY7P4qrLfoYxgZOUlqr2tDiKAR11KMQ5gKLY0riCA7aXWeq3+
ivYRH3kbWHKR3LoL3Xkcz3C1fKVJlgQH4WA2vNY3dbgm4KyyYS3evwwoNA8CYoQR
FCTDXw/FCCYEzzFVqNbQNoLAUMRHFxlgT/iL6FQRxKBICwZW9HtbPZ7zqUwl3zUX
1Km/eJmNjQNrY/y+5dRiqEbHcwrcFoUHtqOurpZEwDa4ayMmRecAj8yx+vTpaC+c
1+CNiSpyeSoFcBAbAePsbjYYJ/H5hxLW01osx/j/LTuEIM0QtjztYZFVqOh4GKzf
wIPKGtcYtYFsCtD6+1h9rWlZCzub+maqLvwkzzG7+AkyR/3XTehuxs2j8Hnld7wo
sPytF2Ouy2cD8hb3zCpORu2RjdD3ytVPA8RTRduboU5dKI5tSn2o7EpLMTArWHJD
61gwM29JC64Q/daRnKoURZjG6axU4QGp6INzMWXZ3G4lllVXgHF0T+nELk52TMm9
zhd+P3ypgTLkpmjjoTZtetc1MTsE/BJQrrBx9NoTWJv2D09rTfYybXDM/YIHfmQs
y30DIoLu2gIWx8UmjWawcnZm/9oaO/UlQ6PYiQwUc1gds3XqDROjZ0eeG4LV7y44
wclEuOEwPbqpgI4zLCj7/ePClAkcLBpPABuazKbVregKXQgmb0lpoZv+VYO1fjDQ
7b/uYaTMSqkcL/jmd16RmHEa8wwcUo0XzN/Ac68G4j/r2CXNtWfs8vW5Bq/sY/m8
mO2mTQ8TJK/lGb20DjAIK/zDsUIbM4m3IC9xmer6xNuD8osQGG9HXrAXeP79idQT
QjwGTR/955/2riz5ieT/350UKmibNsCN7yVnerTn4d2t3/dgmP0NsediLkO6gB0c
03PRlL7jSPm6dg1AiYCFCoj1ufqOso5TRtnJdoYbAyAbfscFMQ6PyeX94zQdDII7
Wm/cqZHxsOBITo6OVNNdFyWYzuUEHnLj2q/a4n/fZQVrZ/ke4DSHrav2CgI00IRi
ZiaCvSiz9gZXy2VrPQsf2KV/Rr2Dzl2RTuLTPXXupnkl/jTuDQ8oAoAjZhWrREGc
EZ9cjuo1qWIVPrMQcFHTp1xPD/NlLc+lc7Ew8PcMjl1/6dp8V+CoqpiF0wYWUNSB
0O39t2Xhf18aJyPz1YWLU9qs0SqhEM1bwDeZ4pWDq5kuIcTlEpyBxNf+DBZvOB9i
czHdT3rgqtju1d9MKvfS0BT6C9qVfkg4D5LfSUrdITwcVZc16dHZn+WUeCMdNg6d
O4EdEaDAzhgPa7BgRQ69qp4vqIrxlKe2Hd7AMa5smVF2OYZ2+UcUdjtsMKBhnJbc
0qyEwx+934MUs7fEyfVNZwu++wnQDH6tPq3ks16zPvrzU7oB+5GCmWSjgTzTEoum
fNSNWJ0+7jXanAtfOnuorG9/rTHklVUDzRkEepcYA5vmtMuSuiEPfKfZFppP9WVC
Vi8ObZWF6tC92SKzywYrI5b3hZFS7ZvYn9ipKA/O+/l+1XF6qwE547zOwAekp2pP
lRw/3tYYZInMIXnACYRbcppoSS8J6SZt71EP9VcfDei0ibZvRHNKCGroEeoJR0I8
Pd3QwjrsDvWp+tLx1IlF8lC2lUdNb6m7JbrQu5zeGkTe3N22eF029DZoryiGSnqJ
6yMrIfQ33n1h8IVyE8adf5BoDOnm1awDO2SNEMfcxgEHu6FeMZnFU9DXbWH+ADlx
yMFLC5FM3o62xXapgZJt8RIqSiDTWvuXJyYVjJNQ47N81ngRL37aqULTOquDQ7Co
QkV2qL4hLSdZ4jyCZOEdIJLA0gBezNTKPchJGufsISb4P/sBgk5teasKU4MeDMaZ
X8tgjmVJTVz23u1Ex2gDVfypgSBx3gAL6ruF6i9nmE/NTPNOTPFe/vfain8WXiEw
7md1QtqPPdFujlnAII8sc29hNqUrcBDEGpI7ScsgTmYljEqvJyWVAwEw+nb0BYiP
MqygNleE6Jv9tNKmmx2iKhcOelLCnZWhzBtWoCRHFZ6OxaUhIhlLAGQUgNxrjzqU
TUvGkVqdLpocvSmV1OudlC+IxpwtQZhsTQj6LKTEC4FQ/7yU7kKNiwV/pkG52h9w
vwzBsnp19HRymztupphG+6VGp2t5LTNznPrXwx90G20wWPNlQT0Bh9zHJDHBU/ha
mNRs2XFZtqXyigbEz6ry8lhFzsxcek8paOb7WyyFCOFORKJUEx7ZbwM/YBqPCaId
C6+lu0KBZV7bq2yjMradtlf6chl/iZp9F+sjrh7CmyRoKO6KVYY542Sy+qi6ns5D
lgtoFcfAJAYWVwilHSru8K5Jcv5iyTMIDe9uHLpagxxpZfWIW/og51eeAfkqkHoc
LVJJCbTXE+mCZG+CZlnMf18u5ilv0ZpQj0RjmLX0jHJDU8pd9gMN7JXqUwWJ1tvT
ahjswagHyLDHSDAO33fxpItOkP8G5/F1Jjuwny7NXM17NNR4TVzDtyezhLeeVQNh
VAOk8EwhgWpYuiKeaO1/uh5lh3Oun8XsFg38BlhOFBtDq1JohHGrWon6+dhSOAc/
mxje9UcoVmBjWdMTViMma2UDZ1lc35Pkmx2tRS6NCuY9s94XpIwg96BYACbF+d+L
+guJ+peB/eyE37cO0rdPpzWcDu1MACsrKk/AAvtvovBLuGaZqHaAdDoZ1TaMQXi1
dMKgt2GT9ELVz66CA4NPha9QO9+SXQ17akelFb4zvV4IWi43G4y0FVR7v+GmrgqJ
1TonzAtMOlnGBBWMuE1UEPzAHoHrAIxI5Vdr53LV4V2wA5HhtuOd0YAHhWJ70baq
YLPr2qHMM/9dgDwTeL0JZX5aHAZzDdznEkRTVmWuA1j+MIGklpvJ6RV3Ae2utp3i
3JsNKeoAss8qB8grNAD4gI9pysGN1pDizE2FntIjn0evo/ushKegVdQJT/Rmbtxl
m4/R1M8E26c0siwWdg8UJMn+HPO3uXCJHdfWXNmO3lRX9PtywL9YKUiM4e94T9aH
UMSXJebwC44tU23HzPnxXauA32sot3CPWasWKz4N3VG6SQwUym56nt80sicgk96d
KajAI8PbkAC9izYVEBoU7DvU4bVhRwjP2jgQd2Jgmc3WpqZwKVMi06+TYBHkNqaJ
vgWe1fmBIB5rLR2/++qFnzGZuStaE//Rf+iYZnagX2SADyfV7Qt0YCo81hpm9w7L
25yoG4WZsy0M4WiZXyJKbHMhrbbMvKAMoXe5s6trBL8CCqI7g3aHdjJU3H1o2ulN
sQXl9dvZhoky9D3iYYngQkW+m/39uBIG+658BFPN4nsLzliReM/38AUVIZr1Jft7
z/Hdpb80JV2GQxJJfix7nVHs8Pi7GDBPji6+1XCVmK4CnfKJ03qalsu2aSBZKObm
LxZSOXD6yR6vyqlO5gqOdQMSlMkiVmDIbAwHeYgVBcqCICPPbsFKYPFKCBKMgEZ0
M4AYrA2jJVuMH3bovGDX3LBJqzMG7AgTAXA9Xwf8+oireFWQe91vcuz782KZEwzl
EygA+dX+kaRll/1eF8l5QPkxQ6oG3KnCfIwmV8niln9HUDhAOeHRe8BUP7d1nQmH
5PX12Lw0JlROnJvM7wGB9CJe1g2wSvvRch5DBHBPyYy/n17KyGcsNE1QBby6Q3rU
qipGYlQgMgVCh0GeoQE7GDhIwNT+VbXx7XTMZ2gZ+sXC8KD1crn45hL/nEHbE/9O
LIvWuxlzTpoPwfR2O1Rj3Q783liILwfSlHXk9x63/zVBkSu1umYaMU++IqFvvqBq
hQ2/h3kdNN8TtMibOXugrGc97cClxbhKBU2GHRU8P1pNQfLL3cXe1qs+pne114DS
ObEolzZlLTC+O8M46TD0+nAed8e4SN5Shpge2aEtVvHmYMoAzGcDesqA4S7NIDy0
BZoe+tni1MIoscY84aKX53a0kR1q4hHmhNaJSf3f/IDcVLDsfCu/ACweOFdvFoL5
XR8yZpJdjzSYzSzxcvOmW8Z+pMZj6lXzSQswwmvwwipJZRpN3Zl9hYTP61A2X6Kr
YNGh8/clkW0M6obavFvC5qzoZwugq/4sHvmnOLXvyJUZnh8bKlVq7DC+admCzVIt
Vkrelk2A5hB+pDNQ5qI6jDi8QzWoN629xF9YsQ1RG2zMUEwjMDpyLBj6Sr29D/Hm
W5iUaxYyROX5Y2dgCS2FbvvhWfxgGStLRxbg25i0eF016thw1UGFtY/40nl8oIGd
gd7658DSwHRT4WxgQ+kvK2oBPJW571DyTL0p3jZE04o3j+T7yTDlISjCrYH/zEhO
qa6WEiNAukN4gmo4wGfbaXDG0ZDuBkTY3jL0EfB0QdFsdcFMrdnlDSRDzsBeLJKE
gInM+pmIlVxebtW39BLmAlTuSU4+/QJzpksYYRkBRNUvOVgeBTQlkLL/2LFUiYSK
H9QrhgAH6aEdd67AeKwEfUjfSJFT+aMb+imyR/EsCliikltRUjOXDwHCbwzJ5a7b
xShwkERHrn0/TwFNHlbHFdo0X9KA8Sp02K+WHavb3bD+zX6Or/Syr1ADs222yOHA
T2iWaH+4zyByRpUjFN67dQ8XHzYCKO/pdammOQ8AElPzOZ5KA6Yl85h5IE//tnSG
AQIKMCRIMAXSD//DMSlqxA72F7FHBz9VMt4kdDitQBYZplUIVkFAlr45kN4gExRL
5+5BdgXYl0nJy+ByofL9zmyPkC3aa8E1dRFy9cLuIP6PrW6J5vPIPAio8kD8VyI/
L0Ve7HTJGak+usJv1D27KM2h9klfxSOJynVArYzM5rsTZ3ZSt/9L8DkSBO5ji9Hv
LGsy5JBUG6FB48d2siOKJQkwREbJ4oyEtF8CCxUSzoIjX5Sp1WrmWxmJtfOpVl18
Ni0BqnRVALVIA56fXQzFpCp/+vwVmXaFykqMbU/amQcknOzLOhN9R37xUzQl0DT4
PZOaradwV4awZc/hZ4lWzYiw4Poh6UFwipzoEm6eeoxGJCEQJNiPHzPzx9alq9/P
J4k8PZsfNpjGm3Yd6xq0cdX12KkNLONyMWi3Yg/Hi2HgTyK7+Zx7idOucr2Lq/vq
c+XTZR56AQlJNmIT/PHghEIMr1GdOhUsoVClCNohPsQsRuOJWok7eBUIFXTGlhcr
l0O7EwRzOfh133G9yavCFktWGCw1MutloZUzuKtqIZN3kvLk6R9rnm5eq8Zv1kwE
qKVZSLzP+QgjW113JbHOl7B696GgQXHRCCFXs31hPiVH99HxxbWY6J+fJOrR4DdU
isR6jLkm86ftyGkTwK3TuIa8I/SX+irsUydSZWdY+ouhV2IgCardi0Jp+1i1v1Kv
TMWDlPDChsb7BqxIoj6snt1TCMeRmPwVe/17L2H3eAu2EsXLpjLgQs2zYRnQYu2V
WePK3rHywxWnRgb+qgER2sGg8IsSjT7t7fNrw6AM83Xji5MXwdRC0LvgaTwV5Tv7
mex1cg0KSxP+170TxSWUni8dL/hiKZ5xdijBZVQpBS4/NtNzmHRLXENsocpls2iT
kR1zaBT1y2V0FQxiau2SEEmJp+D0RB+AUFlMZQc05ntiXtqBv3roGpYEIxT0piOv
C/fB96zB7ykoVoQ//yHftJ/5rEaF9OfwYpU6F5zN3HvCPL2qv5MDQaNHjVnlCCmB
3q0ubTE+7pW+zyiJhKFqeRJdHj5iZTJnWW3u77fTNV4MQIW2WbCsHY6B0Ah8bOEj
hgmSiAVWMoGoMM7wSufaQb8mjTPfPYLW34//a9Mx3a8datorpRRf+LpR2KhxzrWd
6VqvuhJLjjC/7sK0ccVjYxXqj6c8bkTLJW8bLXnAV0RB7NV5QuHwEDODoIU99Rti
kjwsdVZ5h8b1AKNOQGxvQPKaqDNMCK7jQk1XD+Lzx0nyowsXWCqke2NdrdYcAH6e
Y19d8wt/JeVoHA7r6+aphBXp9pvd8b3Gv6jj4TU7amyoSDB3J8hnvLO28X0h3/F6
X7OZinbvj6EMe8/11UY+4QFrUwBQH6LxQ4fYbxB10dGTqI9ZdQnKJ76BpwCua9Eb
eyYrHTWotAUxKakmCm/UihbYzn3pHCmVzK1VjNmW+rQHlnIuZrKV35WNPv3TjKlG
jhx661udFHYc7cWzwci3PLjfagojTXQhLPBTWZdZwzAuRlVzVuNO9w0RIz3cxhgX
wrAFi+kAFif8ENl2cHWjzYBuQBCcjXzrTPDrLJYUB6vMqSQQpnVuVQG//GPrsx7I
gaGX7AY5zZFL0L6BRbyjJ5+SEsMu9B1IOm84MctAWbKf0MzNafVuJ5InXX1HGfPs
/WCenMunwHaovH6J4wKcnHZGw0olvSeU7+qUD7R9A3d3BSyHLbQc1NK0imNiNQ5g
6srOEWwEraU3whlStigBW1dUQJwNXlQrKDgJKliYvaeVvKxVzmUdHzXDyhKtHmwJ
ZAlvLZLGs6W493uieA94nh6uKg4Q1uCLHfVeVTGK3+G1hYbY0gIJ5DpWG8iyfj7H
qn8xpkOIJERNagfm13B5d1F/1bWqgZcnCtGeEASpbjj80Ibn3mtKxjHycZMZj9kq
bw82CoDUQWFIW5OwIiXTkSARPigClRvxUAKTy33YIftrBR+1+IbklRhaUn5gb/z9
Vg7zTb2Z8xMnqRYRlWOKn9BBT1dD+VEhDh1DnFYQVfKgfT2DVUPOccyKVY0kq5GI
y4/R98B01VCOIL5lJlVnE8Yrp4M26m2wWPBw3vlXJBufcGxEF1+elS7Ypwy6PAaK
ok7xxL6PsdHHUC25XHTgBOQKn4/0EaimuXVu3X+jYDQODUBZWzDs6gh5vOmj2kpC
FQVCPZ1lTiz7jRxVmE5cb7Se8RbP2U2fgcqszEruIulyNkk5HkCQnDO6jm7vl2YC
OtESzyS7lgS1Z5ytLTcOu9mbHxwls5pB/un+QzQK0/sVeOIbQd/W6dMwWgjpfaay
W4MERP5Rc7lws0EsKv1hPFQsJArXtY87UtIjfl/7iR5bLZBaFEY4SRcmKJS7gLsG
ohMXv6z78TNlb/7zayaLu3ZNTQYt+Fx2GXv4TZAezTm2ShC5v+gkwfgb28lMVUXC
pOoS0rYIh84VSxT9f50T6etPrA/nqfdRCyn9XBpwEcUzc/epwrMoYMekiCT9sNcL
JsxQOJBDTLqjfL5D6p/tnWnMEWM99csvzJDwZMghNreK/1czqYkSlRqKDS+ADofs
CMuzNOP0pSc3L1IzqMCRzYKJrPyC1LDoHgLhDIdoRX0jkpezzIxLHYhQG57WC009
ek+cV7COkptOBycx1EcCvdEjrBXrN2jI1PMMpm+r4Lu7T0OgrSIrHhzbtOy0YpmX
lFlo0JThAkiJX5sfMST/WW7Sj75tActFO2CA9VjI/kwCjx29LTlhE1QzuHFlsH1c
4pQXekvjDmdcqk6dWRFMJM5xl0nNm/uN45TmYxwK4ioo34xfjGANuty+2AXNvaH3
NCK0wH6wb7OUVvzH12eyu/yzJP/9FOG1Z01m8nZEZuhzUsOjSfIowZEgq1RClLK4
60CzNNLqDWAd0j2obz/abI3nQ3rzJmD6wXVyAAIaIOmPsjt8xyciPFoqJKWtOTSv
f0AYQ59cCJV+Kh/mlKl0biKHLK9L9EYf8fG4NkmKLu2kHGr17eZNQxni9EJnmu3C
sRH2G/37gVHdN6+JyHAUwkhYzD9r2uwKEJ5S95AflJ+dUJZ25pcWb2IdXZlNAkBu
EBmmK8Pl0YVQcU5VwU+MbD7MJRV5vTxLPpRaQNILFtH2nAZypjuC5InBB1oBUxHY
5XgSrk/JqJV5FIgwGdKFBrySYr+vYWUrQ4weLfGPp04ChZIQOBcWkGu4zogCm+OT
MpXONBPVuro07BP9J87Ksa2UN7bJZDpR4ld2HNazddNIMfCB72Fqtrd5mZ74s8Ge
um/AE0bJHfIytzhKKClWhcdcJ0KIj5N/d0QiuClx761TtYFCLK1znQxG2znBCUbk
NvAqns+/rN4E+PGtiodaaWpkUss5T7tYmgffW5lXXG6fJUHoR8hpdJtxnDJa8+vx
nhUP5D9SAtYCc6Crj2+1p7S2TkU6gpDQoAELW7sUlBOnGmpVKZF/HiRVEQ37bk82
ZxvE2lz4WhXFIdzgNHMlWlUMxJhbSsQXCkRLetI/ePNMmf/gPxNhDyM2u4TfexRK
vjViCh+o5/QAHXNaNyGQmppLNPTfrXujKC37ood9xTyIwVoNMKTUhEtQApHub6db
2/4K7+DF/OKCLN+sZKiYLikpfULT4TZvVb1oO61IjJw61Z4xIZhJ61k7kDcKraaq
T28itRZUQJKaUHZt6uX2U+d0AxNA5tcw3yMNTQMjOeFf+e4ZHjXHrYOcEBxgDXoM
FpITnnGpcbpn71NNaTaP1CpOYQWheQg/nDf5kQjWNWzyWcXFMBlbxedISNx9VzDs
S7oX+ztnp0eA6c+Dhpl/q88p7VBqWcK/6OWgUmqPEQbaVnTS0vyRlkeVqLGXK9Ef
7VjHF5ReIJbGkdIW7oCFKYfbGlXIiWRxolOk6TbgJqzsiZC/Z0Z35OtKPHL2BYVj
8SBz2MUfPxzEuutJnLUuMvWT3KLBBe3tgSapEJkCHh7ZNywshrqh6Fgq3xBHbCZv
tMnxqUhxWWjIIdX3BCa7pj7swuDk76CjnQRONGF/ljwvkSnyxf15DoINgFPVRiEH
y1uzi/3a9PyiOsrpztEN0Wmu8RYHpEIkZsjg+6Z0AStnCrJHI3wTH/5lnCuC3bHh
4k6oiAUqE2FxdjnSRjFFoPAi1DZS0wbbRASCuWwAdz6eQtHMG7TtVSs7LjhkbZwN
bM+LfOM+nMsj1RddLFBL210oLAsmnNctE3XBRdp7OVpgTFCIAuM+g5hkn5C2KF4P
WfsZrOmqsQvlHFvSzTg3rbjZSf6hTC7pTPAuKLmyhpyLzAsDxoh5FjcD2FlHCtW7
8+VZz4uCmMRECsMWVte+L/4vh6/IzXkptZu4yLltHm3tQPDRIcycGoSBppIzXW7g
XQzO8xnUPbqTh/tTuHUKaDcUumjz9OgO825s37V09xyAjxIWhb4QviJvWP8Mb67R
kBF2M5VESp+GLsYkoJqwhlski2DBbVf7tGhprTYWmIRHfHkyjUFJyMguelFi4ZMx
vHkSOu2eCOgEiU+prhlzaoQRCpZLxOJ2E/H69i9uSiwUTJG6sjaN5qvL+CoV8sz2
5FqSoh4I70Iy2FZioTfwFMV2Wz4e0Lv5AkKj9K88Q3AbuVaeHaK4Cxk4YCzMECHy
Vs7syWxX2zr1ob8j5TDX7eNgPYxbScJ3Q4UShIjG1QsHR2498bDTuUgDXIGUM+w7
hE8cqIPjf4tWm/DD2thMHpKVAj2n1wfwUI49F3uPJsm65BuEICuoy721VLIHFKpT
WBAiLhewu3lX8zZEOABwM9WQZUJijwI/onqG3tY7uqcJS0u0JrePDnDYELvJ0230
vajs8R15OX9y0Fjlaeaaac1TFUb+CCA+0CnVio0bcAQYbZWgRnzXnniW6p1LANAR
CwCtC1woZ+Zh3aiq1FhBGll+CCH0eyy5YxOEGzk13bAlKHP4ygOXhHTJ36xop0Qd
g/QdPWKoN1LACvGr+RhdXVbxiITGCxgGHfBDGuNQ1kAV0Gr6rq3fhclosElZLSFT
7YmT3FTdsyW2teW8yEOAzs7a/3ZjYo0RCMKSC6s5GUfm5nj/LtNNiPwcKVTGbBbV
4QPJgBbdleprFCMH6Y6xMu+FKiCRyeAU5bjyheoNCpbGKpVA0w9oZCqXBJ1LncMg
FfCIW2eGWQkqsSDiGlXHq+TTraCYFC6mKsOR7MorfZKamFx2/A8GJ2oFcs5Pp8Sf
huCsb64OrT1x5pyjbbNWIN3PoyZcixjW9QX1jShZJyAPa00jcFGUSPWh3OXKn14A
aEMPEY+4IRynvVl4OEuUkyqOEvBpBW7r5HAdb/CUDqQlZ0qBXUGM+i3QJCZ4tjsv
KNOYByNEe4be3FtHaZCGk334L/oTsmujkQ5r+FtsJzk3pKTRC7Gg9NA/8E4/rIdW
wd/DmZ/b+eEH4SMNxQG4zXk42DeGNzFSCSRbAO1aX5Gy6eBeVgKAiqz86Ic4yu1a
Q6YkH+nBIJgz5zWC8+sibX42bpPn2l6osTKjwYdLTo2kuLjN6G/bA6JoTUDdSxMK
pHl6cGEaHSKaH1Aimn5zvH6WxHCvx3jJITO67ajIEgsNQFFYRXeYJgEzJwFGrYBI
T1mGbwLkEAoRtbmZisbkZ8S/VYWu77WMgIr2D/5uSKZJxP3n86KNyV2e5EGqTr0z
9VNOmKDLc51snk/o6djni4KelKgh9LlGWhjIV6oJjQJh9uL3EAqXi0sff17yVf75
xGgwOi2omRMvrCrBFf9pBZJudsE2zvGvWmy3+Bratg4cAyZCSQK/L9QLP//cjaVu
ubI2mG/l0U/0NE8KJMNLlNgl9fJZVgeVUopIHCz/CCuULUVXPeFcZb10uW+3UIDd
a8k0l7lw2w/V463GrucyUCi51hK0hYaZxH1zZylMx72zKma8jDNqFbtDlQsIGABm
xyJXLFhX/6e1sJ7vx+l6wc7WCvwwaD22ifPSNNAEL5Gp6QFfytdWo9JaTzfK3EUX
i8b5KFGhLUfde/7Yy5WckjPZx5rFLPg8XxkmsbaPZZ+la/VSKU0pNaxDGeuD3Whs
4hx5SCmcRi38W81kncjjyIj11RXafLwOxu2vU53yjOrxdygApegL1eqD6XiydqwW
nrxszbj/2BpYjlf4B/5qNqL/trcC4KLgmveCsrueeEnsiWsayiuA4ugQG8VVR1AZ
qlgNuzwGMG6PNuHQPHYIvJM6YPPqHQfifHyw+l4NNpn11UrhD+b56lXsWCqzcjmE
ZEe5jelOmiB1fGwt0AvpNnbtOK9O30i4/CWd02xbtCXJz5lGtUmIHLZgbwlcvdP0
3KpeIkqJa8Je34ps39SzpxLXvnSXvfQynBs0aO8AapNF244w6OBF/YT6pXcBhDQh
+iw9mzJGZ7K16VjqZoP3cYvhrLi6diJXGL4t8VQJZnOxVwac0R6G5E8F9K8Sc+PO
4bMvu2T3tQWZDiMTP0FdxxYr5W1xFvy8ON+EiNUz/byAgVtsCP2hEKXy57GQVil0
1Mz0YnuNu9W3OkAeTlOYSotkQ7mtx0jMPlumuqIE9CYLwQTnNqmjmT4v7K9PiC2x
E7z0ohFpJl6C/1Cy+X8Hy+EjOwzNDgBuWHH1XVrBl+Lcg+NdMAQIelm9JOE9URSC
TjIjEC8MsVZwFEiTPl3FQb5rrDSHuPsqmCyeBl/2VVxfdBdhi823GrRkrjQ4QD+u
j5oxaOXA6eohy13gDlHZWueRo4mWQ6wBOxDVMWqQV51EBkK5m6961rAIQWDeoX/2
8WFqx920bC2z4aX6fxF1fXuTqYv37PoWIyTBVeToESRmIJY7ENmOVZ/VAjZH8HyY
TA5j0d5Gqf00YVtJwJNI6rzV5qPhuosjS8tyQRhN1/VT2/FROUtgvtsQLz8MAUW2
kg2HS6rh7mqXb6Smrha7+7/tFGuOiNymwkEb+OGOpF1zxkG551zveTi835g6m0Kg
FoHRTmLBZe4QYBt3DXT2PujaE3rQMtxvDWhkrEjEMC9itGCG9GA4t2xADiBNdEUZ
MZiP2iFkTUWMw2o8e1nh8yWcA1NcoEgnBiNaoZ1QCFXanfn+M1pdvfoSUtCVZnfn
1mRTAobNzTR9HvW+RqjOgeRYGop86FtbcqYmp5zrgJGeYBu8yONE4T66mMeiAq6y
b3fLDcgh5TBqyijDfECruVK2N8BhtsdHIR16KOICOdwq2MkR7UBf2/wPCv3FiXFB
S7zS8d2gWtsDYc3R/cfiCGZ/L/pJnAvF2uoDiUMrZ4BZg1l7fUlrlf7ICskw396z
ghB8i45u31cQJUzj7p7Gu1j3EYDLn8lgyO08V7Gq9YwbucBQYGCGhrkOm/2MBmkH
nv42bbyyPk1Gd7JyWO3tj8sJuoPbKqvz2epeDzpde5pQ/9LaBTGCgWkcST05tF9t
FlgfF6nl+ud/woj4vcbg/dKYB9MaYH9OUfkaDl66DZpMX25otSGzs/+NXgpwfGu+
qKrV6JtzC83sVol0+jR26Ap3p0DEUW2sUhXD62ShAUDdHn4FzIVb5PyFHyNyxlB1
dSGxFRTqh3CFetddl34YEyTGuo7C/ApowQeXw/NA6bgX/4OCOWvSXVHiYtuU929A
RZ2Rq1iugzPCxWHCCgq0SXdewGjehzr0zKefxnabcQJtm5pFF5ttwHc5iu/aQ8em
QCQfhQQBR468U+RJJyow+n1pRwVKyWr5Oi8Ozk1s19VTK3MmQBA7txAsHDpNgbNz
PiPYGHH++Kubkn+2iluVy3r0zkfXPvss7390oi3OyFbO/RbfbEj/ubWA+Q+Y0qmc
2SheodYCz7xEgkcRqLImwPl57X3+XYF9mMznmd3Du87Ny2jnHISchnTLB8FD3IAm
lYcagIzBHD/lKrBiVh5HXiVde9Em//d56Hm7Fd0Bb+2FaD0tHGSOXj6d0cNl72PQ
46FLcqgd5WMreHePXdKHa9Shqtd0iqUJ/iOHCqrma+Lbp1NdGpvrvSL3YHGKaOlq
ibUfDcnd0U3AR5tEKvqgzHdu2BUIi6KVhN/VI0BQnoFesHZHIHYLvv2bnpsDZXmk
OUw9mvgotafKK8Mc3Gn6HtvawZbGuy8sDcYn5V5DC8Rk6k17JVmNlJdqACc29oqe
ZKH3i1UiS2/E+1RAOjKg9+CXJV7sHR54r4OTMszDgfpcLuq+BdT1nfXil68cjYQ/
FwE7OUMFfUdSW+jXAgi8Np9iAxdQtcJ8JqeFP2Q3/PXnLC6lx8u0iQ0fDP27h/am
9NtXy2IdOuzqCjphA380vhYzQx0hQ0XH0nsJk7qFLrt8bcR6rOIumQ048wTXcPAx
l8Blbfk29KYG3OYl8zzvTmX7xfpo4giBcQZrZtROO0Ot6xQNwVWE8C98xhSOq4XA
gxGGvsrbd/a51As1qUEuuUAlmpUXyLDCzDOaA6FD0e/hCg8pW5Lym1h7gXFPIiAk
qDwdqky0tGKeMJKGFyPhf0DOGeproH4eOib46BmJZspcnP8p0maj8UDnPHjhJ+t/
4CL1yzUOKJZQWsFGSIReqo3z6RnXqIdPGXGBmPOT0xSAW9BgShkkgEWAMuiJdWdW
tVqxFeHkr0Kvev0rL6uYu8IhsQ4oyfgdXAhu5dWCCBgO+kDX/pkswhmWNb/5vSh2
HgdFxo26Jri9AZi/0EANPm/pnGKbshJzQjDzUrp77/A2TN6UNPnSS5/BrKE/7D6r
HdF7tARDlqI6BPCosg1F0XG4uqjduY011IHMwJXJ8Jj5lvvHdGB2Qp6O2Ydashef
HosHO5pzc11QIJfzZ6+bzLUf3t/MJaDMIz2jjdJQRisG62y/7C2E3cFQOMjKk+tR
gEXATJmgqdzGuE8AFiNZIQ==
`protect END_PROTECTED
