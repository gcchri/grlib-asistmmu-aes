`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vznxmDcrhU29pOWaHbmsx8slgJCwgNtTIdKigdOcIvGoVAyqgzHeVHkITSw1rGUV
pdS2lt/qnY0dUNf0JfHhTPIlu1VOefSkQkx4gj1Z61jNF8lUor/yg4Nqefj+96IW
Zn6t0SrFakHtQyzy3Am3qyeW3ZKhOXtWUPYutIfW+35AyT9eOl511RV5a4ejr7YZ
VYq/c5BVUMsvpDnCIgdiwNse7splOHQyKcq/WELRJoFRMRGTa++t6BOTd1lHZE1R
Kxs2+1JBv8JOWtLaPtBL/Qmxet3o1MMzmwnPDIaXrjkWQJqIUnHfIRdyeyqoTZ8d
GwbEsVmQXyOXwQLkdgeCvxEGfcQzsGLIxcaIzXoJVjQZemF7O6MXP72oDUJDZIqL
tPW6OOLqLttnxsKXgDAbHk5PmXLq4nGrWXbL7lZ9y5g3aakXiC2Z3sI6CMvtrxb4
DxJEuP3pfOV1fgmfMt/wPb0HpT+ljpWemck39iXPTl9f6vBFxVyAa5upZcexAYpG
h0cwvyc7wA1HtGuSgeMoYMG0tyj/7FV9QwUGbu9p32B53I2cSL3acjjZxozkLUhM
R2yi2wRiHU7MSBKPRA6aLdJ6MeC0U4dR1Hbs1u3vgfJbAu4v36vL0COT58qjJDW0
gL164P3REstKdKMS7o9+fXO/EwXA5ECZkznjMDdnEQEZNAwhp7ok/3sVrBg7K+zb
Fk0PCd2EPVcMcxPTMXhTl1D/I79tBuyDoAHX7ikZwjLAgtdYiyYQjYoXsRkQtE2I
b7Wt+dn8bqQFGFUS5plYUDcWpe+Q2urjDIxKWqYtGqQnjaIXuKOxRe4T1QTQ6LOK
uWxKi5eyDirpGd/jSsTYqP8mTs2yuZfQx2MvZWxO6UIBxed3PoMbW6tZtUbMmlA9
SOj3TVqUnWWhZg0+wwHQKGZ7dhTU1wIHD3xuhMi5f6EoUGa/A29bsu9Qr20z1tCH
OHZsAlqYKUGW7WheGFMrOS1E7MqxKUF0d2ZwBoxOklYDf2oJs3xQijQ9wPbUdot7
NMnFiwpz4LtbIKOOKHQlf+4LJ7bPKV6SscNGFYG7FwLoezCsTdGGAiMtXaCeCHtN
PtPWGcO5RiUtho/slkS+i3tXiVmWYVQtoLo798DFdX+TBf73vNgpYt9FTkgReq1N
b3az/zpH2A0xUXVHktg7Iv42CgRWTlGhKujfFOqDHmbaXVpIVaIt+8yGIy/8AeQY
ZtbmpEBI4PgRAoTV/LYiX2jqlRerP7plDdGN1xeoAqi9o5N4MrSCdMf/L6aFkS/v
tRisoTYk19PioczsnEaaDX8UIRGfHpjMM6Gn43fAOQmGaXs/NHx3rsNWUDFhQzCd
AESiPa1J2SOindzx7i5ac34nNWjI8+L5XpP/rFvgRE4/41ImN3mf2tQ/gMt0w7BL
9RLUxzzPDC8DZdeVmhxHNPLFGxSSjxsCQC5agzv0end8r170Ljpjah+e3vl9H3Qn
sfa7x1Z7MIJRrbjUh5hub3HlVtk4SzN5drtz6MDE9In9wBJD9J5tyCZ+rs2YE94P
1pFIVOsQmpHHmz+/vz/1vSbxyEYzBLDA1aFT4m0F3igilt5QAVh6HbKh/YscktuU
zpazpz/Xi7gQCET4Qai/4SKgccBWZW8HktfVEEPMUqrOHByqkhnz9Wf/WjE1xK+7
78OgglOQsvuW2aViZGb11YeuPJigm4EdnLudKy8qYEd+3cmWx63R2pCQfHVusvtZ
yZcu/yaDKFEI3G7ckMbhppFeB8/8J5wyhh+E9oslfumL+elqCoJsWL72Kd8H8pG9
Wybl7NhlPeMWLKrPZ8VF4u+LM0ozujy75myHBxKCX+yLp8FOF2Gtq58UpIzWSsZG
/aDHweKCKSPbxbEqU6j8jbB/vydZ8Z0j2QvDZiX2HZTJLeR/h3cPzjachdZWiv8j
778kGu4MofECTlSxfDy2Xj2iVdCZEiKymQ/uD1cBqBv7pLaUnNLNHKcON8ca2PCB
2DMm4JCFQLW10NX3V3kN/VRIWFh4iBtT2UhRNd6huTUvHtHYGs4thtyBEuwZYWTi
Gg5hFZaCt7NBHqt0wC8ZFbrnfuVHE6SzO3KKuHUq7WyCqDal90qJbDkQZPoKNXK+
2I2ABEWhlp5AX4OBYtvUVTSqFrZkgOPzp/eZ+b4HFYI7+cQ5KGfIoDPA457ujN7t
dU8BUQov0vmdnCR/XLChb1k99s+1AqIjX17g0sIKom8=
`protect END_PROTECTED
