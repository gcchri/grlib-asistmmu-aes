`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+i2LQLiT+XO1WuXygy57/+9ShsAYNWY0LZ71UiNy6DpTSczt7cnyMaE3okblrkJG
7ubATU6nibMOQ47KetFd36Wuvste1POH2a038h/ihIsrmZcIMeNq/TQ3Qvr6trUi
0KzYTV/jHk/VzFXO2kKc2VV9rQ0fR0cfReGB2F2b58xLnAGfwmUOpElMzqDQs8vm
NGo5YarU4+HplxvYEY3FNUVCQTfyjofM+IL+LIEHwOnhOeU2Xff+cPDwjenSYSso
HRpIxuFFIlTI2J5lPcEYGJ8ut6vHRh7snhn0tCSofZXZW3Xalvqmu/WGzAYKxUY+
LdwnaFvYTUCY1OMgeiGEOqxU5i7+XIITTalk3S+gKSbFZAiMHDk7omXlTZIibmgj
xRdNwX+HcYpgnQ6myk4MBPHJ68WRDaowpCY4qpvcP9eSEDZxzzRvW7CGSddZbV0Q
qSnKndnoXrHysbaduy5uD3CKYY5kKB+f7aKgChrb7MqEarZ8sZybQOfweD1zXVwJ
IXur+0TgO1rQ85JNe5fecrd1HDiQhGQGepje3X/oMYxmlHrUrTquYDDu6JitBKkz
qDfsGr36m4pyda87ZExnaIQ/XeWERUo24AjYsyP064YFQHf3rZDKyC0zF4F125ht
`protect END_PROTECTED
