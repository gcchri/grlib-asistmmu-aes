`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
28PE3T8C9935U8hgtoB2PpJWNDlNGciCURif6Lbz6hc09HQUYa0J47MEn4wA3X98
8VZnWsNhcJdyJoiyHJSXREfdapX/R1NGFnU12qDLOHsIag30sq5jyBHIxPKXL9ez
hzMbb8RdHiUwkpljBaZaV7mLLlg2cOAe10vsnHJ+ZMCjWLQMqI37BN5bMGJf7iZa
rQ/Ed+3uYARfdoeJUxnbUiIr78pekSQwUrR7aG/E6Oyzq80BTh/TvC74djHVYQ2n
azGFQuhT+VhZkI9O8zyx753IuTFQXubjD2Q5sARjybuvbDTSz3s+EzNIMdZxYeJP
meMJOKZyDv3xPyj61QpVMp6qPx3PTWS0vbinYgE2NuZN4A0eOtVWwkdl2BTvjbIF
q2A07xzNleS6K2QnjEwLz9PG72o1L1XSUkPFKiC4rMI=
`protect END_PROTECTED
