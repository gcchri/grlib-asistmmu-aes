`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
euqs2CUyeSVqB1IN40tiyT4BXQzgJKieEasVVHfMV4EjfMwtGumyoG8/+KPKVkPr
e2v0sdylXKMvvFVfc42FIPA6m8bVD0C77wNjk7MqP0SmgtX8+oXNS0vLgES8D2na
Ijo9O+vM/HYzPhqYnNM/ubIC98uZYSVIv5bkzkLlOU0Qj0KQxUkB9odVnTGhTs6Q
NjEgaXMSQ/xgUXZcsKFqqDRVSgBb01CR1c1pPnERyhzuZLIFyb8Z03UE8jlNWo+y
CBA2MBrR+6SyuTrM0o9nlg==
`protect END_PROTECTED
