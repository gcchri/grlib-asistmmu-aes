`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7dWs+m1tUaOGTmwVMgA/64Oh2NAE8gHU1zoUW3OHSanT4PfJvfus1GdK4feqdWJd
MQcMMiANfavcZs1TcLsOJKS+wU09q7wkRYkieU6WM1MuoxWEpyeQ+7URDMDx0+nb
f3yIjMch/LN/eR2SsrcDIq0k7uAld/lXIpu2r3akbm39CZndOsUGbLGZjVFyOWbn
lwCRy23CKlmjom+Jg3T1+mQhWkH/nJn3rnWdQHReWj/d+LIOLdefe38DmiMGTBkF
B9uVqeQt/GKyi8xOaYfYKeyX/fFj9rZfM2sMVTnygRpyZM6BTDRwl0WerjsiIQXf
kmAO2jEvwD2+Qt9RJyv3PYnJS2QoJDQckkUwTYC8MoiOjCxW6g0WCrZKgXjXJ/p9
yuAIeOiWA6aUKT994zkYeWZmVfcDNQwBtQD0MuNCc+8OIMG++OadD8blEDd0STd9
3ECXDao+5ec8EuDSjkgLR5oTiRieYz8NEF4Mb/X2Pwk=
`protect END_PROTECTED
