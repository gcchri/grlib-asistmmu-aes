`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TudVk+8pC7IDbVkNobrgkmqxjUFXbK8VwMRR2dqS0mU8xxX+7Qs3gwRyOagH0vTf
y5Hxv48AGg8u5wHR3fZg1CDdSVhF4YrHKcO5rNIA4BW1hivsfSrQYhKJWpPhDTgL
d0neUm9Q0NH3BAqxpLROd20DNoALuI74xvggcBtORiKrv79r+XI3cJoAWgY7r6bO
a9oNYVxghgbbpr8aWkJCHYSAei05Oqna8zFZvdo5CHdDzdeibZB1Phswhz5Sm7Y1
Wug48aNCYCaXhoAfDJSs9Viq+tpSOxqDhwxK04hhZ50Op1TuGQb1/DLvfOpc+5Iu
yPifAowZZUeMG+AJsnWMSPEDVUS7ieckdc19XMjpqJbpqQ1xg15RbgGjhXd6l3mt
tkB4gp3Ltuu1808SN9SjIQ==
`protect END_PROTECTED
