`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OEMCPW6cG/lHF72jk5zYuSYQCjmFR/R0TQKvH0GqoG2C/k+69MEm3HiBWfyZDAge
Mjwo95cRTsj1g3gcunmsEuDvgjbk3dfWA+KkNyX1lQBpvDP+yqn4vKQo033vZVIA
oRsI6xhS5CfKFhNl3rtl/Q9pq+ugUcp7Dte1xsfSzWC1v68GUDc7oBe23k+yBjlc
QAhP5sgHprPKUuHhSMs3me0FIlh7/vI9bCGHycv6TTXDjmWd/HX7yBXlrh/rBgeb
ycgnAj1p2cCY0LSyV7XG7z0kHvh7FdZXMhA2iNaKC0ncxjkzdE2Ypfm8VtOQ39LY
o5kMNT2yWcur20tCrk/azm6XOdD1qn1yP+NYq+pHJk1g0PFkqBMpRs/9zzSIs9Sz
B4pbYUzQ3vK5xBn5wJPxuWaog43ADRLNHsgpzMqRQznya4AspRNghlCwDlxAtqp2
3sNRHc0ufIKVe6eE2GVIOR8vxFXdKHCJ2+zFExa7sdbQU8XFKp+Fb/k64jhGiM3f
`protect END_PROTECTED
