`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cru6b5nvRtz/FzpBu9sGb9IPLyewj/JG08hFhG4YYSu1IKchHeFAlBKjbxqsXFo8
RAWt2pGtcC/9XyIkKDJg+gJkRE4UbyLh7xqIIsx8S0XA7WI9FxsTkSI5yT1M/Lqu
ndqV4JXTa0jl7S/hBqJAM3+1CYn+8gAwHWAuq5/gpgVt2dfcCT42FH/6y3zQFnm0
0jv+kxCfQh5rOyRITMHsAFVz9VWIPpE1xNR6mTSyhxTcBOEwJu3M4LZaEuqCIPmx
0iU4XCvN9jbNSYmT6yl+0tGgCLvWCgR3kWNk4cCbNrefjOGDYxw2W4mt58LtD9AA
YPuY1ACEL7otRIAUb2LeBO27kJTkz/EtcatGO705zocGDHfMBuyR4s/GbCHMbkfa
8pZmCmzInywKB80NyZV/D5yDQkvGa9mE9/0RbPcT/bD5Yc0zsB6w5uyxi06hkuHW
IJS1kDFLrf66nS/oCqsOm8CGGDgRxzj09Say//o+UR9GhFU1lrFhfZhe/peVS3wX
fo8o9pddV8yA9x7zbQ6b34vU7Ml6Yl6ArxlAla/1q8HWcHKKvIl4dU+X+ADZZwcB
a++4ejO3/pL1tk0sP3UeEXVMOsGHRxiYSVZYXiOYFnHpMW4E+ibXsX8rpQTf/8Tx
wIBRheYUgP8GL7uhBuyY/oJNP0NBPkoFvd+ZFS3+8NiL+2iJ1oZQcWxLPwdOs2gl
yV0wk6y8fC3jb9j49/L8EeJI7BLaUWj7tUA7BOVJsJIzrIW0DTcOMWAsHR4ecqo1
eXuvZQ65W5TiLeJhwyzxMsaFoYiCFKkJ5FqqvEYuhgMatYEw7phui5UbcL56739P
WFdkQVcNfTGQgwM9YDrvPlO9kJ4brk2/OagWFD6NLffTimW1GzWYsvp2grAdzHV7
QQTlSfogZlh/KePqN2/gbPaZEf+lZQ67WMWHQz8E7J5GDjpTUcHCWmId+gZWj9rq
3s5UaQMO9ein1sF4WO04mA==
`protect END_PROTECTED
