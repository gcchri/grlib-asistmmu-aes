`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qWm+d493nx+PDtLvjkz3jJwASt0VXpcM9lRSDTQ5SRItzXE4EosvF8RtQbr8cSPT
0zKwxfaopQ+6s0ovcoVXyAgMlLhBfkOTSf45ksbp5BXPNNU1MHCjBnjFRloItBJy
Et5wp0Y1lCNIKxjVpXN/FxS+ChwxZsjDGh7LS7U02SSZHEytRZMDq5RlUHwthHMI
okMP13s6OCuQ3xLcCHLG/RHp9ywzK2VRhCZZqJG1ipbalfeeTQHZWrNdsxfAl9T/
7YGK5AzI+PT+8dE+iBJpkh8BziVIAkhulzFj4ws6lpsGXk1r62Wh9xNJ6p4d82qj
db+6RIQVFiympBdXFko/scELFcoCg+J2ed8Zk0KuNIwjxImNE5tyFLWQ5IZoRUIh
4HJD23Bq5orlzpczBaNif3hoPY+Jx5qYlcy5zLUSNCwDIW4eeJmQ7tz9uVqOjtER
2hjY6Vi5n1oiiy1II/PQurjkheL0uPTSOhISxI/Dioo=
`protect END_PROTECTED
