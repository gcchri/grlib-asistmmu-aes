`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BMmcn6Eere3QZp6NGitmaDWm6Sf3zlCpXrAknZqCMC6tFqZVL7kslva7XrwEArK9
uLjVqHSPs0GvWx1cZKPL72jzHFtbTwEQzyJsMmJ7F6jr2XdOoGtlO4tV7LWV/k1H
qL/1/x1AwjoSqXQZ73p+GrC2rXJiCNnxBOiRsoYyNmq1knntMWFkRJtAPrQnTuMU
TDrioPTm+mQrFnCYM2sVLaK87Mc1qxDTZPmhobzBLuks6hHLjuB0BopknnS8vo0Y
Wk2U2d2e60z7MChnUGdVHkVZSlimCuQRquRwHGdOrbyr6ah4A3ycfR11GYES3giu
VeQvhofyEFOgODT3Q8Zfw3m/7jXpz3sct4rDzC4fThUvtDckm4uGN0QfcyDPQFCn
g3NXU/fG9riWYI38xlQ+D+ivokAc/AbVWjvNDiBW26xAixRbXzOW5ueqWrt2Vzvr
iNXK1/OnO1SNK4jwKmLMpcctZT2ky0k9WlZT3GA5/9ciAYowr4BSDz+8pcnkgYZ/
i2OAZlvEH1G0V9KtzYCUcUlqKC+9qHbXGzmnGhfB1LDlGCV5yKJjFuTF7sRhy9GP
6+j8onK7pUH15NcE4lkAAxPTL0ttQs6fiu24t1MvBaZqOXJg7OiaMmdgkKgJ9NmI
5kW6HMLMMtH1g1kbKO8Nw0m6Ab0ZAPHmfrMjFMEaRoPQnXG9JqWJsD/0L4gYsuTl
jgdP2cIwtIWajTkid303kMRz3WwDOfV3UDth8Ywh733oUK8g85cjV4OXOYV2bPn/
ec0Y7irqMjRBPULcoic7Ey6m5JFMHgCtiwv5ke1SlAZqngR4iGle3JD2f3vtxxph
0LSGEIdNJ6FstTWNKBzx6U/HucGjhFA9xjfNk84uPnIFL/s5A7MiR3GbccVJOg+i
46HZ/jvQ2po6tIiNoK+exl1uCRLUN0CflKvANM+5CPhZZ4pohfFBooNt6yB4GGSb
ZYVwV6XZapjx6dwFh+hmi/t3YpelB2ap7UiH4z+pf4LQcVf2STmP7Rm39xpEyubT
vJ/9hAr7986MC+fuMbAmXbpbdT2exJYcMbmOmI2ecgtHlCdbvoA6g9rwVURLLLlX
iUdBwlCi6fFIMEaShq/Gjy3ISi7eBWtaMnZjHqFt0I8T2OvmG3HIlyxFIdbFDez1
YoXD7i1c6SuCf4ka1JRk5DDjYBUIhyZ/EEygFUVyviGMByjTgJv3c2Wt7/ctr82W
igAJz6M1RB/NWZxXjRDWSg==
`protect END_PROTECTED
