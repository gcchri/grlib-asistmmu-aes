`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qlXaM4WNe0PSaz0S1RboXh7WGT97BFWpl1TE/RQlP7Sgq3+uLAPfBhnPdO9PVP2F
KhObBMpHH/VEQWYk5WQWSw56eD93ieIqMP8ToGGQ70ewM8wh5IifRZcn4XKOFAAu
9MEnE6mTYPmhprYjIGpdP+pKTCHJPWp9S/LRwckIvKcHZJQiMg7Lq0qA1/W7Dp2X
AcdnL8cHIuJg9tONSi85XEgD0o3ArmdH0RiHalKSqrlBccLH81EOsCLpjqcC7SD6
IhCpV6Os3IhyjcLurBNj8PnIlU2a9F0VMDxIGh0efJ1GolTnzccK04I6WQVKB72E
OsWaQG3uERl1GHdDVEOWNbU/cicq17Bq14TNLVxrAZFBq2Ddr7pXUydH0AnrhuHu
MftuUiQ2lXJF8aL4OlDb1WK5hKe988OIvN8SLr2v/GXhVH9krwFiCuNTM9VM7/mI
fst20Sou9fi0hlRj7W9+RX/xmE+iScdQO/u4GilPtYIVyJapkZTnG+tu42YSs4ci
pylXWLcUnFGeGrZFkcpnD+7UZHYoTnDUqE2z3mrwjAU=
`protect END_PROTECTED
