`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z1LToLyO85MUIUGM1J+alduWcT0fJFfFTw/xPuTyDEXn40wyGZeCxuAfUCxKd/5N
62BNlv1kGmT4jDoCkkbePfJat2j+qmjzuw3hVl/0rsm044YQt+tXZMxdpONJtnGG
FtT+WCuRoglqkc3EgzZA+h9THOVUL0RC+NlQ0Gv3r3HpD6j23WrcMSwxk4ELm8dM
Y4dZlagkfXDEwDhPKHb83Degf6i/4Q6TDumE7xp9/AGwonOyRL/LbrvYreAqBiFT
Z4e3D2KS/BAT9Pz6Zybh5P5RVt578fRj2YjFuXfFzglcnDImBCbcbcuqsv1qa7GK
8+BiRRfz7EUgYcqoEukObLWpTNpAhX+afRprF5075nWTdnXvX83ABkQcMC64qmG0
9qv8aGtrhM9Vp8gouaaVBRrqMyRJQmec3fZXcll5DPfVnqxq5W8Stm6Q5eVUQgAc
cKJwkBcwhWmim5ZjYMd5bk81EsCkg0tAgKLsMZMp5q1/dBg+h+F0txjoVxJUvBPW
wdZDggscjta3U57y8ydzta0Xo7OgFH+o/D9FTjd9ahc=
`protect END_PROTECTED
