`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dr8QcBfWRM5AJbTVplhwSgKJj7EAYBLLaprcq7BgDDai8tmCpvzpYPCmLiDGklkI
JQr6Gb31kBK5w0luG1koMR/jbjLIsEb+8oFngFM7MPYlJHls34+TW1ObaDCZGH+q
q10eyg64TP/airu/pU22JueYE52qdKlz1e/KVESGJHfB8QTbItbdoJZs84EUKN2F
ItXN9gQVyURv7md0BN18yZrTWRuaYJuGyrXBpkWppT+mNCQ3mxmDMGys9gpSoI94
cfOTdr2hEsGGlFC2pLY8oSsOWtuBoF0JWVJMKdNsDP4=
`protect END_PROTECTED
