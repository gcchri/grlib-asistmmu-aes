`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CaVhbUNCPg3ZorS/5g+SQWjHR6QLrsxmZRu5nUSYQdBYVV3qGO1SfSNkM/mtT61f
qgUWnMKyMadoAN09zfwA/lEqIGOMrGbkZndL80JQWHdgVLHsC4uhMPQZZPa5XVhr
wLuj0C+26zsThn7iRGjwic7XrGi/dlSAacvRyoZBP7H35pHXUzS5rVS7nvyunv0/
FOhjQ9iksCRHhVJlZpp0jQ2nViEVl7cryyCkSZ7eCE1K/+7XdaSv/cU6sL8ur3rX
tlXkuv0/vvP2BZ2Uj9OIFYy6RDmOHYymZTWQ18oiWgcj0ZfNjPZKvK1wHoCjH/ff
jESroNQaH3+TFI6671bMJA==
`protect END_PROTECTED
