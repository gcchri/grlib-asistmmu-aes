`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yf4KB2+KqwlTTkrMj19WSG6qeYJMDEaGHsm03rvvb9W5IOxwG0vy+pX1BYzNvNEo
rVCorHMNzTkn8HSPqC8UB7Ws2OzqoSKDH9ifzgBMx/F1vAtSTCbP1NpXgkzA2/wT
OE4roLBEgUAu/YumJ3C6iseFtFds8ha9iJm19DL5Dk7J3YIojgvwWFgCVTk1fDEK
tMLzDhDjHZlOtEjaaRPNQw/rCDNOqEwHEkuh5xhxhT+H15teZsvBBF0eeRRGYezT
8so47gop6JYNJGL/wBH3JG2ZgOhqQ1D0OV7QJtT/D9kup9P/+sHbd1O/hTD0rpTT
nrxpoUHoCtm1Szieqj2RigFvBgd0ShUz0keAfVUMB/1ZXDBlZ/K8Nf6k56xrga3W
4NSq2mF78y4ofwcz1JEo+sUoO/QHKGkXANdY0sO532I=
`protect END_PROTECTED
