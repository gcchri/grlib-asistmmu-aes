`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NfPW9tx7penP0Xkpuuql8/xli6EcG/1hgeart4xBZLMxK/fYRG2zlhqp3iW79G9O
eDQ9OK+pqJyFAza1YQ+JMO3lgbS0hhRDQF4361WGHla3EG/fN+wzvkWBgNoi3MDx
T+bWAfIspiPfnQECJc9x5THAM/1tnBufgTcBYDqwOor9yzPpqHSuU9eLbRJRFzsZ
yT1QDCcq19NrH1EXBBbud8JQ4NrctZD3XtgmpwK5VWlcHvd0ge+CwLuBYbBJxwrD
7vqOWAZyHGg/faxqtuZav0xjH+Bp//wpDF3dM2sl2DfQZDwCDOvZZ+ku60OMif1Y
va9hKVc5OFyy3XfLlAsURcR0xo3akEU0jckEfftNdrpi1uCm/TY2iERjs80WK5rd
3NEMBJFlhwx71Hd0wKGE4g==
`protect END_PROTECTED
