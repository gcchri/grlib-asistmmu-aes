`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RZt7nO5lL8yc/Ctf4HAlIB811jXGHC9nxDdhZOmFfoI2sHcLiDbVTOAnMiPLpebR
//80XtGC8Sd2eTBYHxK/R7zRLCZuyDNs0AoYFfGofxqkrOwgjB+VxaV1a8cutdpI
21UALbK1c/w9UYedsNbeyVPXidZSMxCF3cX12QJUuQVflZBCsroof59/gu2oficP
c20J2UpVWR4KcYyV9xxHUmsl8VnwXD3F8Pd6kRVSmUhN0ZgwtNlOZZ7QP7ttp7vw
y0s93iF2RdTKpS4zDpmSprPmY7IMqj4J/ey8Wx4f6GxVz75SUZHHHMhqggrMPbbT
RGsWAws3YCUejk2JQb+WGVGcoNQuFLMF8oikmT7bvUibtRhNYAu/NNI70nK4AGOl
FZk9mtfRnTrlK5tcTCLuPZODznzprZuWMozwrhH1vr6I0x7Np1PrA2uo8rMvMsE2
6/e8yHUKtAeJHcerZohsGc9zQKH1s1zExpFRbJFy3vOa+cFIZ3RUsg+ivc2Xsyzc
bMI2iVbcIoeL2b3S5ry9SM3gsD26gCY7EP/65cApZlOTic6VXSS81QNxyEidInui
ol88NjgkOT3Cx39aO9bVfwLesj/ap6djh4z93qfvWarU1CABomr0X4++beZdjrjN
EW3An5AXloKdf4CQmn6B5HOMd5OryJzIu/MJbZjPsyfE3M+FI06Eo9VHCDQSrVI0
pR+ROvy3AKc5QgmpWq7Bwwm7o3HNWE+7vR9QPuc0A5Af634VyBDnI+GSpyCGVets
PTJAQq50LU0qdZ6CLMvevGF/28ljMJr7rKcpUVtZUxkNDoT0Nt0XPIz0H2qTBJOs
Hbz17F8BJebjOg/TgB0Azv4t9zAZX433sEHu7YXZQYPjAfTAo++sxFmGZYShZ3bT
+srLLxW/9t5UiUGqtORol5nuOBbs3avfabatwRYH/eqzekys0LXZ8H4Gfh1ShWap
SxMvjX4idefnUnQev3/P0TG11NJksAF1NKKsbq+rQ1Ch3noWZItfMIX46nZ3s5S3
jpsaA80EHLrLpwl2ygzDD2QLIgPWzUsQNjojy1rS2ddqb7RNBhgmdJ5Cfz+wv7qP
CZqL0kLZJYWR3VKQqaipjb5OkfTB3MiBV3f+A8LXXwxFXSB6pOAAfWAk7TpvNI9V
kiW58hXfkdToxw0swyWJXmb4+L0aQY9AWljxT+QeDP4zG3GKSQFLG3Q1hPDUA9SF
0p9eQtyJZrzpmyjtgvYzGhxSFRdrcvPlw60EcX3/FTEamstvPcdCJRTh5ECeNsLP
AfuReyl+xp1uWSabd2bOGuhiz3P3yHSxwpKPQmnfUQWQ1CiLoLHrGkPCxvQ/UD68
RJOaOBR++VHfPFjptZCq3aQg4NcOh3N/g1AaOel3NJsdkKoSZ4yyU9bU/dpXE4f2
4bsYjE8pes/4UgNUTs8sSKqdTeDQ38fgCFhJJRLGnkYcpla/y9sXFYaiCjixgiKn
WcrJGyXOh4+VzpBsXMIUJ1VkTtMqLmc7Z2gPuXGAZIzd/U3hlXzsZfwotQY0Dw5E
YmIEVLOUbPU+dMwdJUI5HUJVOK7l1JoP2HaZ/Am0xJis2nAQBgPkjw8eybPzQYGX
g4SYj3D5X99edsIOCB184aQm2uZqJnRvKCXlpIxml8owzj/Sm1sajTKlB1Ob7NGs
zpNaRuUCOxUIKG+7FueyiuttipHLsDr168MW2PB8DDSlo5TIJ7+qHiavqhJG6rCF
9YtCFJ7n6iNOvpv60V8nb9DWr5RuKlSVR/5Nkfea5aXrmYfpM1+h80+hdwJJ1vMD
hbLUI8pyiXr8dOS+5pVMD771ANAij2M7aCwkUA6BDRZrsLHt2HrUx7szY4YCfRop
LosMmLvyNMdkkgnoUBUKPACHIBCdlhaKTBmFWdu9fYACurTiF6aAVxioYXuxXQMA
urRnZsMaSWNSHBc/P6utHv3d2+CRE8c/Xx3Dnbi6babZBzBXyBKqgltrG3RPbeTs
KZqi9kN0tuuhclXAz7GbGygpMOvDaVUhosFcIdbw5G+h23Tudd2a/+iT6QsG86C7
XZiX5vQt+I/yEHORptRJYW6Nn6N2GIAekri53tiT7AuZ8yTKtXCefVxUTVL2DC/z
dcXvW0pmXyrh/XUqPL0TjUvwqJtqflpoO+5KGN9B7RWLCkvcDNsffhCVN8vV4adk
wxqij/MHTRfPeEjJPZLAVE8WCzJp4QteRHDKKrhHMyYRmQw2e9r1ng/gFlQI6NyM
WbTBrlrUjsK5loi1UhzzB1lnxiqcVZhdSzy4APBgpnqyqAAJ1i4RsshvXi6iTP2T
+l0JzJpSyNdZuYdVOmKeBfcZ1Qoa987zj580jnoz6FytPJAq0k/nYF0DSQARLlPk
c5q94ORAMvrlGFgjRVny5LTKEHk2JJmZpDL0+pXJVcUuDNUVG6rj/nWsNeccxM/q
3WtlTm43CojG5Wsl1OjDsoVPa56iKQLxS6pEJ2+RKfXVOziRQiFLYrYL4kViug+P
vEyE03QgepyCbJgUUYA9R9xfSTQmthcZSH/r5X8sV/OMF9kuB0M6IkraYfqAxbZl
ZnNxWUAw41hMZZ5NlSZ7VQ1z2ySGMBJJhMAD0veNK9VL7EPZuSn0ZqHPBheUKcot
ewRR+Ca+YZt6SNvZJ1sMcrT6CkKb1NiSH4UqsQU0CEXVPKs7/DZuyvUcdr0ElmY8
Pu9smZ+v9h706oH5dff4RxvNtcKCA5WUwyDqCwomCr+JiOBn3s6Tt0v0wPJ70HzV
OeCXFBZKyPD2lpdOs/mREOB9hyKByoytMsHr5ss+134zWk853fqlCu0CuNs1i2eo
gV2hT9x9Fb9u68D0M9XuLW6nTHG0MeLRmPQfpZY4+6OScihJjy5oyGBLdR5HFU8P
Ci4rLoa86IWIs8MulCH4Z7OQYWobHoWFsq8ITWjjm2jm4SAsk3AcSwPXcCKx39MD
dJ1IhpTkPKztPJsFxG/vLa1cQ1X4u/oOv8UUubh3d9Up1JnvMC/DNmSKCCrJyl4g
aDMCpDZhwb8UGI1BVC0JvhCfRVHZo678ah9FDPDi3H5mEOchQ+O7Q/AkEF/ISrhP
aHk/8xjmUxyp330u4QqrQdQesye/dlp5E+ac1zrETDtD/YUWEgcq1S8W92+LmxOC
59xkKQBFfk6E5+FMIfmCrwhxn0a7jYnjBDdq6nWvDRZmgZIYMu4Gyet42wc+KarA
I7hwlCkS7o1tCDhnepf2VeynmoQ/Nq386lFsXZdPpP+p7qKn5IBQnN22jsge11eZ
/l9t+mghZ89KOPzokzAvpYx4Rf7RupgRUP2MctxxTDWxhTKMM1G5pmwlHaXgR63V
dJnlveeZizpxIxgJyUda7PC5sbv7eH5LqZZYw+5M5j2hEAgAmeDymI/ha6OmPdem
D+lwBDIkZJNEtI5X2peNFfCNud1OPMy/96ONhwecxLTd7yUfCsTe0Z5tr5+3sbLV
70EPQlPoDvtKfhh4Lau8/dgx0qmjQ9ouoA2Ij1KeC/kgk/KmvPP6ekI+LQGOBeWf
e2TsfhvwhN0YcYe+iI7laoeyHpwjY0qdbagpqo7NaIPixpbo4MJXd9nTqTVbCe1S
XpfsIxUwDQeUqawpzHYqsR/Q5BS4jta7g1SZmEeZKArpGQgyw3kV6b86BBpGSMfE
n8/soGIE2eQym8qrhnx9ylqoEkOZUoomh0WeETINrmKW5tTAdTDAKQ0dqswBrTW1
k16tuC5ERnBke2mULbv/El0y7GoYdjA7Jvoy6da9NcHCBCm/KI2Id+4EzlUfSXLr
Q5Id9RiQouevdyD+NHYen4yKt90O37hQ4vm1xfzo+/YEh8yhi0HXm6zUHgMtnGJc
ekRgKuMI+kRz5QDxRMZ4whxwowz4oNq+Gf7LOVG5inlGPyvukgvCvlEMh3MPUiv4
gsUPBwEHhAgakEUbrW41sPg0LJ72UW26jSoV6omIqHMvbuNWVxUDsTLHoKjNMYmR
X53o4FZr8FgjYsDk6O2ejU4KdfgN4mYqttxQjx8scW+DsaAKIX8x9sXMuBuujEkb
T1jfKcA5WroCea/kCF/tJTjKg9IMDeq0S2WimonY9IOs8aVVppYkKjqpHhD0yLio
DjzEagDtCLeZL1RSfgkOj35gb7BqQWN/Gl7ahj8Lz2rsRlvRovGVYhkBPDyErWUD
zUxovAX/+/JJYFsAk070a6Ht8Jk5EoDwnKaUbtXHoXR4mbdSMBgiA1xe2VAqNCOf
8gwlxFjz+to2tApkr/rpkGkUpGGjXulqAgamDmyq2Jxa/YnTYljSLM39u3efbxxo
d6xPFfqBiP/cP9SFXHPOZeoObnhNSLFf4qEtspvwQwQiCPyIEhgZsm3fihd7bkB6
fH2t3Jq48Q1bvbtnft+WrPd0EorXVtxKDRRUsjYZNtW92Gz2ShRet+g+GjX/auHu
u5ebNDe95oVSwatXQ5JMv+gnZdYShrYpUjCNjVNWr+0TvoDdR+Yb07hDGxRXAy2/
Ig7VEqxlZN/X465sHJyZ71wUnkIt1Vj4w+xz2Iv9ATh3KMbMSCcTa3ejmyAdfiRl
y2TagSN9LqqXsIl+5KE5M5QL9K02Uq+OQb7xsXShrIic3p0m3/goX+3fi++DvWFf
Yq/MdddtCXSSiQ+EySXdkIXuEj+bTsnPIQqG0z+ajQMbK13q0gk1p7JN6S+Wkk6k
K2aaY4MI55igbivMyDUtg5u9/IrbUNCbPoOeoSXXx/d3SzXIlyTst1ECd6pHSqt9
G/NF3RUGg9KR/6uHqVBH8ASkXS1shAoMAlJXaV3QCGyDSNnR53m0Ba8aHeI+ZtlI
e4faPil/Q76ZvxMQb4aF9ar6+JUoUaDSbRn+XOVy6H5xvbOrBz+Knq3LO07up6KZ
ucTQw1PcwAQrdBnuAXH4kPK/DN60hujJYOp1ho0VC7VX5ECd5QhA+AFWG40Fr7RV
aWCB90EgwlYaLGuK5pvuZUBtrCeTld156gVE+shL2mctms57G1iyZqREHDHs9ujf
6cz6il+vzpkcahN1YRa5zItxuCHhDaGMTfBEMuwtolSYr/1+k4R7VqWDsywCZIQI
Ty1xVvaTnKhoXASHgz8NQoeiDUOna9WtB8C6HRNthqmvKHK9CARmxdoyRIpWFVzB
rBDt89fWSPnC6qJSPxjwtesuJ3K//qxUyTgF4oPGP6Luu2nJw36Y2tLngmbGrs3l
e+FDKPJKY9K21YT7nicV7IhhqeN3owwI9atxgWI504FQY5mNabdtSNDZUK4AE2XW
u2TG+AsMJLS6eS5P+egCMsRomwUItg8iPkDu53PE8X+XrMj0ozSilzw2uhRzVGiB
cJrIcUL+Yp6tw2tJQGHz4zLuGAwJD/sgcdZGYUVntKYYUa0OSmJKxfbRsX1cPXPq
kSk2QeTgQseSAJVPU5GqTbIHP1DQaaMcF7QK16U/ebxvSFaSAkaM0SRAG9k1Dw2b
BW2Pd93BQHQNpf8T/LuP/j/1bTkto0fXy7F6+qQwU61gAOr53CAJ9O/RX8f0SFg+
OtsCGPAKL9RewolEIUeF1N5r4Vj8VSEqQSFCazuCZP/Y7UVp9ZIir1N5JfcnLHpp
dCVILVD4ddwzJ6SN7kF0aWa+bKtqPQdc/MjDYWKV+4e9jTqakVWbBuugTxN3wSnE
iDUVlaMDMIi1mt0m7pt8PIekEKkVZm+V3cPIn3K90Ift299bKypGwMC911p3BKtB
FS7qbeq+8qNuLb0DiozJVK5hAW7KLe725suilIiQCT4OUTy74oNZVTcvdMcH2BOb
QJGEjp+W5u3KQCPDSFeEMELgsStODpXcWCecVDDrKjllyNVxQMKU0o7pAOOJT7Sg
Yx4FjDRVLGX0VVNBG3AwnvWHz1jkXRKlHwIIWyaj8IO3yn4wZgE05//KZ4LbgVti
YIZbPiqlBuDnKM4tSlAKdEQzj9vgdIFUa4M3NuM5adC2GVu2ayVSkm20SiuN0Daw
PoK4wRbslmaflt6Hx6QNVGDMNW11VWyjjoxDgGBIY+Oka0HOGBdD+X9MEgyNJmmk
T9hPGneHkkIebOvZ5tE5jQIYz2gk9KmfoKo5uNOSCywfIuxITvfHqpiTAo77N8kQ
cmkDWzfrBpWObCY7PShaWKnES4T9/eEbHMi5CGFV3XAh+IeyLVMbhm+f22oimIuv
Bs5uaDwfZR4DNwBo2N/MM5NlkhiR97x4zjounQXczNwy5M5VaLLXjwg/5M1xmFvP
35OWWBJPNRKZ7HtMDGX+VkbzZ9TUqqW1PlmR7Foycs0dp19qC32/QHpqyh9xGJML
CQ11fk3jvenbpLNtMSSWrAjTVRa189CyOQvCCttlwqzw07k0aa7Ul2bWf0BV6som
D3LHB6xJlg+BFTbyogzqGGyLjet1x+iDU3xyNKd18MXQS5nuXLzPClhPQclYMQqv
2vsVThRTTxz8DpalmFm8UVAlORkaC3hfmyPSLLW9Zum8pOjodRFinTZesk1b9VfD
riDYpClc2k/Y18wIDxUCUKqrFplNzpUpTkzbCyZp7A6vjrjEHPpkaj8P8IZG07jQ
/QblFxRfhnuNdwnYCJ7o5/7nCPkgXNb/THjIr8NoRG85YbvtT3RGlC4eZNAHIEcv
jp8PX+UyXhzpp4KnLgmtc7kjI+u/nWrmKWWQAnVKQE+5npEwXpSPUd1F5/LPn7ch
gLGEyQKQQE61iqGRtZ2TBaN4CrvmiZMTA7hJ5JH2EBRCAkND7wviIcr6/Elj29iz
CHY3Eh5alLmcMS6UFCOLvX0bs9thKpg5INx9tInay99htLAyYiCySvR6S/FMRMqM
mzVTLOEEvZ8Pas74qI8oRsvoipngZB/6k3flWOylRF5uHAbW9IiB4K5rJQzFjpfW
7BRVvVFeL8DaECSvjW5mhJEAfPD/vl+FyWeMWkk0BmiV7Z6HdgDtjlYJ3nPjC28b
ZjxTHUWimtE8vETZw7ZHLNG8o1mxZpFV8gqRuW3yDBkM8vTbvh4PKQJ5SvX3EYTi
o4HQgOEq0vPnTusMtFq3C4lUMHUV94MArgJe1ZjKqhXNgarx5xWR90qdQY3JjEcZ
Nr1A2eZJRRi8URt5VQiZo6s81eEerf5VYt7JXvhrFKRWOokXmfe0v7tIpgUGG7PP
fG+eDLySPER+XWcTX7cobmdie5MR4NYGQfonueG9VvPaR+sjvXNdKoylOBChIUky
Xt8JL/SO+cpYaRorHUBIN5SC1CHxTXOp0cN+pTAjgaNYETKeknfTPIC671W74lLK
9w3/Fd8Oldqpf4JyB548/kwrH3V/4AdyUYxbvOJV1C92nFnZ9mPnVZ86rx8dkNP4
KK3NC0ycga/QvDP3Cz8a0wLslvs0TmXRUK9ll2QRgEtKNoJakkUnvMrgWmY2b5V+
PCep6ENWZVUV6ZoijMA1gvytnwQn6nEKSrtP6GvNvhgRQ+z9J4ORZG7zV3uszTsk
PS5Nmo2x4hqDVheHx2GluXKRImNt5si+dZ9W6YHQWvF+uveA20xoRNf5/4Igw61U
N8Xz5vjnI5+yLhiVeRATbxAJ/V55Uwu9TJ4gpknbWNH22S74Q8bkvSLFQk0FWZIA
UB8PXR2VV+OQZ5nCN/HBXL8W3YMIuLnFetOftX6obR2IbTEsCCnJIsLSSB4JGFyE
zYzlDQThHqyhyMrsxdHl8AazTjpI4Z5Dcm0YVpkjla0chYmly4CvUc3ifQZoU8ci
39YQK33Tcf8MEqGki7bBDiOLJr4pLTmVrHKWjraGSLnHva0Vs6ON1PgfP3Xa+YCF
oWlKWLuwsoe3ezHseiMkZKfJnKc8ztxcIKAhtwF8RidU0IvpotNcKc9DPj/cLZK8
CllCilxE+2dJB72YNQ5pXIN1tJvxjMN/Iglo6/fsFboo4TIP8nxQUD/xzaJFn+Th
l5FwFploDvHPV3aqQeROy6Arhuv3QDQfM4XYeyW0XtaOGfcFnanHJ95D8ikv8Hhs
xOhxqcxyKTEaifp9r9PgX+OLhKPXyjOfNzggm8M0/jQHZnqZTJvbfaLUUuvJVV0N
IugeBWLo1VoXPEoo8vi3KhJRZ+Gwpi9p7xM0PC/SEZnZL7yNrXklKpJy5Ivli5Xh
3T1/DlbYEfODGStih9oKm/H8VCAiWD1R0Os7VuF+A3ByBNt1c5TVYDCJgBnXTlpa
hGKBBJb9RKwDw/NU/8aaX7cxPazRFRDCWYNx0WyF0ABbtmp9Pxk9P0RUG1qSUg2W
lSdyt/aqLOKe+rYXm1XxOuJW68cTCGZEFu/97f30NQpPFl/H5SDR2kvamdpoNMTt
fv9f6cqoHbWWnxSWRzvKb7Dz0HWEOUz4wy2rk16/KhDVi63L15exocTRo3Ctx/CG
7OaN7Ek2SyiFL73eOnwS1jDjTzkUwtCGuaGnTmzt4LMQbq88fx6Pp2CSGhJrius8
E8IqrCbjHlpyJ5nGjysQ0waoSZ8l1vMtPTAdwYdDbALw9OrCWGGHpY74j2q/itjE
QiCSuLJqAFbQYe/V+lt1YLJAI8B2z0XtNtrBh2lgQ4Vf/XcEjNamOzoKpKPnQPhx
ApVeX9Fl7G/BEXOZIf3BNq+BjIIBrMhgeKif9JvXt3I7grSnK9moWOW8DH0S3qhF
RIYGBI514nUp+wiVRGqc3K5aE9sjNCRuu4YrxsLBrSuno2X+9zVufSvfRtHFWOZL
rFLtwlRX1VvPLnSEaEx04ae7WohyHGCbQTX/TcC36+kseIEXdM3UY/x4uiSmTX+l
XPVFz1Mw9uEMiCr9lOCu9dge/aqfmQeU7i3u21lyaUcOyRzx+op/Ea/BeSEluA4r
HhDlOf/+D4LKtA9t2CYOOSloWt7eFMB9RR9DajrKCO1pX0bSvbXTYpYDGL+hILpI
jCkQN8ktdJWMs0MDUWt6gY2elOZl3jhF6ucVkTIKsQh3oLl0zyss5h7lFK80T8gG
gGvP8puXYbId7u6pbAkvwoETtY4uV6qbmh0Ag7dehNTuLBkBDg6gR9BqPx0sYmkW
46N0OB6FqizpmhbnH22b+yovqnWHrN7bKIXr9Xx+Piyj9lOpS1L3poDgWcn70E3I
cs9LXuwGURkmNaSevB/ELDHINTCJjZrDqLaxFb0oDxdR8cGIawRlfmtsWI5QAXs0
Er7n06zsVFz5dXB5ltzvzBjIA+S3u15SYMx3D1KfnNBi2+/o0novxmbCBxLuAFj8
9rfLI6M5d/1412wCTRQW/hq1aI5g8S3zlzhICxJ5kiZlBChaZwltf0F+WMS+0Oj1
p6Y+f3TxlkQGPhifWiR5ys5QCCE17m0WgVTXdumVGmV8HiabjYjm7+T3x6/Cbja/
VpELIpEDCU+ujgeMZ1GPetQg8P992oofIRfKWfZKPtIl5DyFkMaK0uOKFvMz1mju
eewVteEXgq/kYBpSTzVwN5Gs97wTbzaHPbhy/0EmPfUqRtDqYL7vYJ2GcmYAgnqY
5B7CCC96sYgUbR0ZAd/SqHxfyOYFP2sQEupp1SInuVAVaB11n5fVscw5RuEkWKc+
BFVh3A9XmYQFuJddfARxqettUep5gsP+HlE0u1r2UqmbOC+mzrBWd4I+RXXNFB4e
eF+uqtRoXhY3qS5VtU9Qdxj0HaLq6x+EBPZggVi0WWYx3uCPT9KWlZpIAVa/tFNT
eG6iHGd7KiFwImM+Te0D0C3e6EkZjQ/NHVxNrBAJvyj8Tp+MD43eRDK7BenKLgd4
1QclHC/rWdUFdv8loty9ZlL6+KfYiq3Yu6+Mnb6VU0B8iKJXcCum5cahyfGXjMFS
prXzTfBAvhYQRBwfnNYgl3niFXAX3KKiD8PZkwgujqC3BwNjaeHCP+ziSC96xz/8
wGnj+3zkbpo4G/koOd7rkh9DP47o5S1qZ+pgCfXzQE1EmdEThe3+RLpb4EYbY9h3
drSYq450k725rcSzTiji1VvSnnFKHO2ZAZ7UnR3AcJxsp4eJXHKcBldMi/oDfMq4
Tffl4TWIMybXI+CekqlLHLdxlLgx8hZbGjB2ZMNVEBViRhXnVn/25Aa5e9Fs3WCO
1cKrXPNsow6IEVatZLWcLIoosmuxk9TMblhuo0CXVp/wxX31/Hkv6VLvTkxFv3Js
CAn/CLf+bc0QAFusF7NyXlN+vevv7zb86Rw3qeBAMqO81dm2r91IMG+GvF+d/Ous
54rqhQLfEuMIDgIwEcYxDd8OfRZvoZdajvy/F0lxs2XZN/zJ46edaOo/1mcBAMNO
V3uQPU6K2xOwkddYA+wssG4AHFmZg061X7spSf3aAPM2CXhzvgEaBUmusOVqzvow
qagt+K65x6j/K2NwCKSfw3vZ6v2h6NLkKaT0HSsovQGG1y5cAHIgOG7RXqOTPUGy
fDfDHVtkqzhCG68+T9NOT5rcwUmy0TMz3q3FXR4p3kWJquPZodwchLQGFGe8Tuq6
XSW3QNk6So71M/4fAEJx0ZvhOHT7auJR2buOqZBCT0Nq6Koz1eMWqrC6yNSsSlf5
PKTTpT1Ul6YRSmALp4WLLIK5ArlTeJMGd6DASld4rYpzysT1oPlUuljYiQf/nSye
XVItd169cZQdnj2XyvWzvAd8KZIE5jNd/lfjxESLv31Gr5mWs0aHy268pe5DBXng
pdGRksCIe9HYbrCUpewfeZgLaSrhPqd/7XZHTtkodJeo9Tzrc9WbcWeHnWVxTit7
WQbAYavOB7e3DlASMLbB+ZS9EJhuDbMB49H45kn4nwnpORG0unNyFoFTcKOLrfXJ
5Of/OMdBVHx0q50N59X1fyjjbQGnaJ0/3yHC83yjuWJoQbM5lrYVfP5M/yC+s81R
zwIdQHgAuOzM72GxCB4V8fXr0WR7BYZzZ4psZeOpM3SgY7dSBGKxm6VJFlSq4ltn
XXgwV2qrwdEFlE3LL3Lz+dG4cW3estDC04BL7YZ1YVzARvbQu/8HL8hn9aq8D5UG
WmnwO0Y8z43YuIvtedBxWtAGqWS4Ot2amNdFn9HZqNqpOSWQkODDgINf8rdPYUkp
AROLdK1WJS+xBKhA4lHQ0/xOKVJ5NKetfLFKX/YZ8bt1GHAQgEPtkE6UU/5vblbq
q8BXLZQ6QQ/rOwNzlxC1F0bs40Dp6CjSK50SJfdQS5c0PzGChGO0LlloiNc98RZS
r8847qaJif4Hgs8C9FFGBCoTiQW1j32TsGvZbZKmEm3GyrMydG3oIln2HuQumj0q
X+mqLVFOXTtA6Oq9+WmuP+p5XVnm4bf/v13QEHqhfimjy/fJ8s/eUUqlavDPuKIT
`protect END_PROTECTED
