`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6mQ2syPKNkd/MdaMktB/Qw97ML8uH8xoDnuSmtE+Imna2Me6O50M21wMvNlyCNd6
IbduqadbEQBklyDfdBG/m3nBxKqvg5GAM4DzclXA9oqCMunAciUI453tcIS7NOxf
CdVHl+w4E/+DjTX9AvIktOmGyBh7AEpU9cVhEr6sg+aDo4C86m/LrkAj0G016lvb
s10MCYtLdHZddKNPGQdmix9k9CNsB5YtJ4xx2Z8q0CS2BJL0vism7nmsAgeQAD7r
llmq1bMIK3DXsmkajNtkXQWXhFF1KMeSneRziE6vxt46SwTe/DBVq7lXY/qAJl6r
nRMhAlZuvnj6LzRUqw6PHshsBDykCkhlyCT0yxJEDKB7qtY2lJx+6rkobCaLnUJf
KieVJpcbrPOwWLBioccRamgTxAygd8v5/ZV7nPVuRu/OILOES5BpTPJa5ozhr01b
xUVV+Q9TwfQuy/RJjKK5pniue9MKWhebivCfHRfxLKNliVa4cQkoy6g/udOmv7vP
E6pdJP4KJ+b+W39Gr2HPJvYKMgqucQ2+F+392KwQs3SyI1Yz0Q1Z51LHcgGyomDk
rsT+ArJAbshbRvWvovDgsJ02gXPfIYoROQNDleYG2tVJyiHB8TDGq6pF13YUVHCL
YIa+8FjAnymhqtnUMNoLmKntwNqj+p+C0H9PqQW33Q+FBJRS0Vu9M40akFu/kS4L
1Eb18YXCn4Gz1qSu/mdMw53bX+UavOmEENKXXBg3ZUIj7HHQ91gGAq/JDL6E53wa
emDm46dwpW/4mD4AGuZAOfobK5Q9++0BSTIsfnQlMZv1Um/XkozQe0vLP501ccIw
LIg3egejrwY8ibE4tsAjqeWmj274iZ+329Fbn/TvoTXIaqfIpl9ztEYDagzPcmLJ
`protect END_PROTECTED
