`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4ZTOxzLRfbR7JzUqZN7rNmQUTxWagfQLYYSznHCMePUru0XHjmsv1B0x4vSv8N85
yr8alD4P/6AaYreYbuC11Ghe67E3toybOGKqIaBY/WJK2tsMff9VFCNJ2nt6OW5S
UawbQr2eD0iQnMm7ZNL/i9kcdELDyoKBF7QXtrmLwNdUDHMaGTMfkoE6/7ok1d7Q
6wo/rLv9AIdABsLTiKXHDH08j9jIoJQn+qPUf5Zab7h0J/qrAC9FJ8FAilTLTFgz
SNX037UNRDFAtL+uVe0vKF+nfYz3yHbNNlpa7lSC1QDre02+yxIuXaa1WKJM0rIv
Ws01f1R0LOaV0ogy1pPGg7R3Nf67F264W8pJVv8LQienCSq1BCcSK0wBw5JXWSCv
Sxdu2CI5KTjqFXzZw36IF3Lw5uSpb5w0EWyadCMwW9RrVOwsWI3vRkNFfQkongSZ
xmzadBdvA4L36nmbJ1yikQMFsILkvZXTN54M959C1G3MtBa7BZcjD60fGJMg6ga6
7iSOTbsx8A5t2GUoJCIYr//zvqG6HbtodOSaeH9sq3sD2qCBZKLQTGMP0HcLqAGt
22q8H9YIWwC4oZVZqueHoyKxymc74iGzltlXWXreZQM1SUPOb8dVtqaHFPgwRcNb
RTR1/yRrnTstOmrW5ar3JQDKjGMN3xtJ6KisJTyiM6KcmVSrvC5dKL/nbAuUGmaV
EBqMX1kE+VeFgWqnjw9TSyzvJSCULzrhjO1pSDZaP3A3KF0Bj+51Ogf+2ii1dAih
ese4wTIGa+/zhRzuoFaWzNjJZHimP4Ki4bJreE2tph6/0AGIclO05WzJL/z5KK71
+waHRklyLcRiqckEu4YrHxKBZ8lJxHwaIi5qRktc3ps1daY8yGVDNmEk1nSP12iQ
f22K88RMzzaDlhkcx6fVGFaV/WfR5uHpncH6QVP3kZJmAMHRi0kpnNDOImCqs/ew
C+XILunwNiBNtuWCDFxLPPs2T3o2pxSSSNsKa+UO2oT2NqNMvHRw+FdDPd7TldGd
pAv9vjhR1aZfgH7zKuL9EocGhV9lr3jRXF5OLZGhO7p1vGS5DnkRAc4Df/mlON9T
9MXkq9NJtajZGfCYZZkxEXogqU9vKS/KLc5ZVrZSB8nd78risuIh+4tbTH4Y/K3t
sRd80SeWZPFHWoHj8musJSP2UhaqIzSkRLq2q0Ef2yLmL70xxITjfnGYnD+CraO/
BdVIPw9WhZizeMHcUC0pGaEcmcKPUmoHkWrxL70M/cU347DxnHo4sPhxSjjxs3j3
hk2D+pKtTeTe8OBV01WlsquRgAj5wi7A8gu2IDZs4xiJhNsrGHnmu6zaubewCdGj
Sta3WFejQua9dCiOF8ei8CaUl4LsGUm0disg+S+ab9UiDaWx9afEIHJ4cWrTSXv0
0RUC+ubsLfyyfIoRc+kfokIavqf5TiA3mGVulF0lZ5mS+hee4w+w4vkiknITGP7J
1F7Butg4WkEpWAyBDx+uAhC8FoqMVgbOs2d63TAygE/Ek7nOJccl+Er5/GdvHMdE
OhWR1kf2UocfGPKrB3AQU2tWqkr62XZP0JCXsj9sO96s12pyeHQfF+A2PNOU36e6
R3rkwNPpsTFeDw6otunYedQB3XU/7mNP0bg4AQJX90I1uHTua27XUvpId3SlUTV9
HzlOyBQiG+lajLIHWLh9yKuUaeVZg7YuyHCuv4H5KbpUqyTffrLu5TZFBosUEQJl
YE4zKNUj9Q9ovTpulSRLFw9z48HyrQdYNP+OttD/3TJxmEe26xGWOVrNcvv9iDCZ
oj1cXJzEoySGY/iybiGBrD5rFyia8oNR6+KMM0DMWneGCS0fxaThibZKuE+Pw6fH
IyNWyNUX9iXLgWtDBH6z94wV5pDKDjkYLQpLD17XgMKfK6+p/VwQ/UdZJXXdii2Y
ol3TkU4B58Q6jHHrwKt+HSaY6XHM3imkrGtXzDlMmNefIhU7uQC4SJgfarU8/l56
9mnir3JXzUaWS4xYHYiQamGpq4lAnITNiV4b5OKZJmUnQtw/vJcuWeb7BqJsCXCl
4XDxjEyJmqaPl5Zwej/wuojz1WDU42w6p9xWAjsd8eUJdyrkEEnX398JUBTay1Op
G7MmA8pr3cpwxcMqko3dnYDxLV185Rivhw5HOar5eFQE2T+urBxWGm4mE0OZTdsg
h3s9QT4Rnks5M6csI1Fv4Kd9tzGQLl8qp9u0q2XwsCOZ4OF/w2cBFJ+EfX01lHzm
zADGo2dwEtufHSYh3PjHp8huos0kQ5spwSQIjAbaNUkPXrVy3yamw/a94mGe3FO1
n7W17+X++FhQJm5Fp6IeCfhifFQhLQyXXtmifLYf3oNWEv9ilr1mAFH1c7hI2sgY
LskXW8d9rxKYDNLofV5aLwjZZaTyjb0t52pNLXPASpVqr8fECg5ZOZheSdtJQ80Y
OB7zwBS++ODr0H2UEpI00Sp7ges1jz5C/SpFfW9bYecvS7iKPMj5WaQvv34ckH9/
l3PRlzciD2SQ+AFE3jEtKiFXtQ4jawcGDCd5SXGspXI0McxJAitwOlvg5XVHO03Z
ycR3yIeCOuJArquhwAzjx/t3+SZEzlworPrHrMLUUpvFDG8N4JjNjtX6UX/KCCTT
q35GrJNAtUtWyRIJ4FGvTud90fHNQnuyGjj3VSUUZlOHivhfwnVJx/533E0wjE8V
kR6Vv3vVEfqxK//tgYBgX5w30RYRV5w3fF1SxG2378n+zEPqWGoNYY7Mh3qjpB11
u1usN0MeQ1r/BqqL9ecouZAq8tuIfP4PmWzo8yg9j6FALdcKTrH3uUM5UzV96aJ0
hxZkuUSlIL4G3IzwGBRavRGlMBQ+vCIWBPbqxfbxk9hNJRS1mI2wdAxaMAtSq9Tg
PSFfRcP6E9E69THycVKkxe7MynvW61p0Jwdtm145hIFwY1Ioa5w3X3udhWZ0rBBq
WdGxJhiK/DhpRnksIXQdm08euBukWrT0Nz1XcpBRv3P9e+sdEJrh2ibP/OPZ5ar9
Wk7uVywH25fRmijL1Tmc6wuajrV/kpR/biUtT/2daIGraAWUVuAS92NwKCSaH2qr
CMdzq0m7zSVfRM4RNCVqxGALXUZLWscBS62aPt/xOhVezVTq+EUQUnkFcbWXR1G7
QA+Zv2Fwd2hG/XDY/9uBUGOqZ0rnbw+kUbRnhoNkshLL7HwouXqUecpCmgPokpU2
HGV9kA/CajPvFDK2g909Lc/QlhQubGlJZQMPn7hCnmMDY5hKkKLzPZWbzxcIayxe
YYIp+QMEV1ZO+DBmzERACnQcpSOEOAOwmQEbhhQ8dMMd2EGejKRIndgvfQnSJ9b3
vgqwX0M6LIzHgr4Ik5XxuNt6bxx5UK4kpRFHdsRkBhEY/r2Umy8iCnWl+ErfR5xp
s7SqIYjChpseO9hl8zQvPcacjFky3iCbPA80PwyqkSOR3Gj55sPqLU0sihaB9QjE
fWj4KZGTjJ0K4WdlxRvkhHMVO/E56E8bvOc9PMt8QZs/5vx0dh3D7u2IOa/q5kj3
D9Oi3PM/wLG3X5qC5DiH5xgj1dieehu5+WgoERZPqbDBfxgAS5C/K+TsF6m+ttfa
fjNFnq8QBKiDTB3vuzR6xwPPEOFxYIl3CjMOAf/j5mbuMQn88k6BZTZ08u+tLclB
2uMDJOHE0j+VDD4ors3ULICpxHEbqJ4EO/Hs2zVIiGL3xEKlPID6OdO6h+jleyOl
ID5jqNMQ7Aobr/ViPxjTw4IvHR3dekV6y5G0uUjiPzmUzNBqIjfs0T7QEZPPUG7d
2N4vMNZjK1dcu3HZq8JKoMuSzGqJTqB2pCJzaW/vz50ShlcPH03p7DNUxIOG2Cc2
DUylra14+Y9sc6APs+CRELxt9kSzbqzfVTqwN943lcLvKQJ1rjQtI7ObXRTB7W59
ljU18SbGVXEwvYISJ6Dlh4JgTO9C+cpFBH9BwIpPzQ/eVIL+e7OvLyTYqsuVOccB
jNfFLlcBKtksDgAxWhOZeeoq8zP7P32bRW/vwpI0YfwEk1PkSlBNAvaMh1rfkomt
RK+s2Vn1D9OsOGqREr/PiPagK/oZCq6uBQnIfIb+4zJxV9tebn8DiYUuClB6vs/S
zuqR7tKhc1isZXcPZkH2l6GhOjMF+c9wrEF9eoCSAB+ivtBKCchawhGeFJXzHwWE
qAnVvYUGEBakuN6s9Ry9Mt5GIUm3oOMICBrhEGMZxsEbTgnrepp+YK8NEvBw7eIu
bsnjWI6BRsi1FWnczcTn1iKFj2nwnQnlkz6QVVUGciTsqWoxwq2dSExX3a5tjpq9
e887xzW8XcovuKbhYErx/26AVbo2Ti7I/n5EF4Z3za1sUm8aCLs3z6yVUXnD40B6
3HXst6Sx0b8tLkIKLvmmOPq98b0POU48HSt4Zc5juynWUNMJo7eeggBL68hdPvcV
wt6Bc3M2wQtYcEMx1bVkkT4dcpQopJZlOHXY41z9L7vTMvjWqE+NWtMb/0xtETzY
P4XE/JJx6WRbXJIFIcAacJWTwbXDWutUz89HAHQmGHTjBwIwkRqTmihk8yur0PY/
vj87cxdRQKKekF0fjLpdsKXB8XiqiaiRdG0e3c8TOqqrDpSDRaTrYHlEhUXdjS5e
IDMp6Sewf6LtNpAQzSCCPnw+TYkf/k3imrZtTbu2uN9yySVTnSBqMWsnOtZ7IHw2
q8X8/Q0nfFcYkXuKUSS8oC9WHvey2gafJKdFfAur+x9WNTHDSq/CEdDGHFL8NXyd
KSSTXmBs886j0WUzQessEzgiZ02fJWTMuVyVN5bD34e+pXqILsUKQRk4dA3jES8A
y/r7e9+JjFzb+Qb6+cgMCECJ8TyYuBohwUpe/77Yyiy7iQfxjdKifC+wbVQ20ElR
wA7KseL66EMXXDidlcKH2o8Qe9d478LboJvQNbWctEt3L3FA1F5oqN80q4T9bpzM
yZLoHc9L/Qtz9ksWhkIUM6EVLXTJJdmaKKyDi4sV8egQensVs9om7Klm/yM+ZIr4
3PWh+zoxZt0YbhHdtP6d5wBsl/WTBY/pPZFYg5IgJQOVxoIlSfGDnRTezUEh9QmZ
fWfvit0bNQfJ8M0ZoPPkzF3XJL5MmPsoJQpDIOsLoF8b7RoXUrA0hEVXQ6NFFep7
Kjz9ISyZzxrg2BK+7Gx+L6HTSy8A4hGaK1AmFzjW3sm622LRm0vVC/P6SKMQRd80
53s58fEqFaGyFGoADBvKAZ8npBxsHLe2W9c/xb8au1wWTGnyk9l/qzlubZ+zYh5E
j4r+MPZ01tn9wF84JbddAPHpF33axoisK77W+PmZO3O9RgPKMytJ8RmAZ+Auv8w5
kGkxhxHalHQOuXRRH8aR1j9lQwS6dzsvAI6BnI6UaJWpp5Ri8n41sGGtOhEH1doF
equWgh6Ie3+ZgyJpMTqAvy0W4kcTT3sXI06mS6YyyVhh5C5prx0B9AUwSKrSyuFg
TGY6s0tfJ5OjcboqaNaMU1obsYIg52Zb/Ee9E/8M0s5rDzl4UWuQV0grbUow0pOh
mvGinTpkSe/9Hr2wrGVPeATOA80rwA+Etc3e9boM2j7xMPXTsQp2WNNGsVEAe8Hj
oNEvMixIEJlSrLDPnzzDi9FlA7vNkimIT2h3xaxBdtIZEJa5SVqADWqTmGAohscE
PhZ8yzPELhWSjGZkVrFj53MNSuPG4s5FV89Iz0Iv1iVwRDGmGfOb4Pl8aUU6nuka
+lcH6eubTemsn1La9I1PlJZIdBNj3if2DguQiDaIn5b8deLiXN/b4TbKKCbGwpRH
nx1IGMN1KCiKixxSEm2a5VZhPvmedVXasvsmZgYmKluBhOK74mpv+jqVJU6D/bdj
w5B3Ir9P5cY59Gz7Z1p4pyimTo5Ytanm/uIJyh9TQxCJlj2eVj7eP7yao8b559qh
D7F+VV7zDiHXFe+b4cIrwxTtxm6/wLitMT2MzXDtBxaWV8JnlmTaq7OihV87QRWE
iWaOUrKBel3IUaRajNfzJNT20Wdk68cBq7VPnDMsYUWMsQT4Low9pbHLVM73AS2D
wYtAFJHAAsE+cjaDWqdBvrtUd4IUoRkb0H6TTJ9IGW312WkKSShxIWgaAC00Y2/H
lKOTmEuNLV+uRNRSI6m95JLEqSuIYjV6Pub86Kpza4084P75bfRiHkpJeidjnIIJ
shA/V5RyOlDtr8nZMqKc+xg4QhjbNaPHxIBAz/ESzaOcvtJIOGiEI/q/U/j4BT91
/FBXRt5mug4XnSXWStHjARPdu8C5eUMo/hrLpjqVfdXwdSdaRrkYKKPKtwhu8pUr
pDZLkeLC82z5tTuQhQp6hofn3DypsLbCo8mA5J+VTc/CiCDI3O0KVyHVL3Fk+DhJ
3yhCQtnCzz85sNNRIXKEPnOeGsaoUBSjcYj69GPN5OnsPltor+OWW8VGJ2Jwi2eY
UrC4WImLMZH4aZzm9VNhP+tOCMGiipVlH9onzIG/0ComxU7PUDExR8+fHq+qne/1
kuIforRuQnZ19Z45HCGn4j8P6oq0O9nDdFDXBmPKLd/dnxOpb5fvDHP8e8ee860i
1RRofmlFeAfABPN1KL3D56BY7uAoUtKpP9G9O2vqKkmPQ2pbAMn7dHN3BFDS48YC
FDHGOcbcnGezqZuHp+PkHfBiSTGROmSouO2t+ieI9or4+SFkY/griL+zejKAb6Nm
lrd1o7OOltg2vq3HOQVGo32yzy+NA52YDJgIM6hebg38JsOdNj/p9ruztuySedQA
e+n0StWUmgwu0JumxmFT9mqulVgfn6SBlzaoPWEuRM5Hrc6yKdmXRZnjlv7HKAa/
muuVglDyLBjKoT54hZSKNMOfE6ut0vTwrUB6DKb/8FU6tkFVQj4lxIwmjEoLrE7+
gtlDiTJLUDapR58s5fbLQe7r6TKepI7g1obGvr3zGTEDvfHttr1//Jg4pz8UGDwY
hk0U0U4syjV/EpU1/6z3G6ynOhA2w3mNEq8VNzWM6IPuqkxZBMQ5sVpYDEXZn9eV
Xxigq9sqO5Izg8PMBbWF4CRTlaeUij5Doay7n3zLwS/07HGFzhW1PymgJQ92wdeI
ZbJbkefG/+7f19iv5PYrtIJQs1ScmSzqp2M3v9fSV1IdZ+BKNJvXYegTDIXwayQl
agfuwgHzKScF4TwjpxYlqx2RpNST82kJK4fYBpGFDR/RwJr6v2TqNUNgqX152xF5
TvHEAqSYYGuSWwndmOAosZ6oA0ivUzisrbUZ3+HeXFFvowYQ7YqGU4/4wxx8p5qC
II2YNGoxvxBegb26wafBOYiijyXJr5p0vgVeumq1SCWs4WlekBS2/NpT5+sqBi+L
xuDpeFfyVxiGduYWKbnzyBN+1jw+2BTkqwZ+EUjVAwdDQy1JT9W75UbVhp3Mh2RW
adOdmvv1Y4XFi5Kb1tTQrpr9kXNz8rvMG+72DcFOCfO5kJ3GC+C17K1QgUr/npSk
tHC1INEqxeyrkPW34UPlzgVQ73L1hAZzxobn6KWnJqNqoPgcjsUdDmUB6RfGsbtz
kYhF07VvWj4peCKGeaoMwpd8ZNE/iRteDwAs3zH9jqcuYNZ20vNwQ4ofwij5Z/DJ
tZ210KcCyxa4FUnl1KDjbA8IaDyhB1Q/TqBhRHt/OdFyyNvZo59vbtfC8QNHco1h
tJTTn+7whOiHwKk+bpqdp+DU7wa+mcAJdXS76NtpYUmG00dQRFoG+jkpvsc5eFrr
cQtnEdWTQgORCaPXOHaQ/3u8u6PD9g/tm8DORAMzP2OsJVOJlZwVTDK6OmrKvwvg
Mly27dh0VPvHY8dpl/jyTnuL6FqCfWQOGhGNCyVnp7h8V2ZpE+7oGdWIW/ekuKTa
chwlrsYPu2Nx5sjE05PtDowHQrWNTpYkT8JQXxXI9eDUQiHOFY/M1EjpEXFY8C8u
Wxl/8Pl3ZC/joS2n12DYGMOI+gzJ2Fu4axmyhS7CSdQEoDoj856b+fpz6e7id2jz
HtzVh8vellVx8k8H3MjfvNYS1JL9r5W8ibbi42ZezOyoHWBkcne4HJc8jG3ueOES
SDbwEIdUEvO/GdnyV0eM0EFHdK08fKbCt3IocIAJ4zQxPd7UxHA+dlOoBwPOaBKi
XQbykg3pUoI6WiZwXBEEk1njbZE//t2Nq/p/NSz1FfajiY0jepkp/3au0ojWegNi
qtfHfswk6ix5VCVjf3C9WRrBd86S/ahstRfYB0pNQHco8aKqgTc2yhEEXm+mSr6W
AqZT0cdzAp3qKW5AX7mw8s1YytriDAnp6NO8dsxKvJFVgmiJ0FRUvMhiHIn6BDX3
nHnRcbCr0YFLCgUFXaSlMaDs/F8hqlpf4DqeNndGLs/l2xJd73LotNy0Hgbq7wh4
781RSWbM75QwePN9QgQ/fNg725AXIWVG3P26Sqku5bUT+aDE9gOCRZpxdYHORRNu
R9tkEjWXv9wnkNUBV0yfLnMmc6hzplM0CQdydypsgMmvmf+KomNkrOlwZ03ECe3H
9Gi0c1vMvZLvEZWRKpP9VRPr3IavAqJ3t2nYDyQGXquN4++LVB0U+f5T8BTZf9lg
`protect END_PROTECTED
