`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nJ9Onm/nUt87nIV2P/WVm8A1m00y2mAB3iTnkMSGdq8RgxpLA7mIEvbFM6dhRXlo
0MUhfi4paZf/mu3wLJpNk0s/RAx6u+ZmU3EH11oCktwi5mFgkYrGNJgeqN6IFdCZ
q6V5VK5flp7J3bVa47zXsb+bPY+Met1+WOqWX4/wJW+/np0n9eC4MM5P7EnTo5vF
2EOY49UKo/Pj6P1rWE04++HWyYz/SP2eZ9mFLqkVJWm7/WHe/xunzHIcYOWt3ZYl
/tyu4c1sulHs3iPyOneq/vPeyT0fb9geD9bCEWxqRWxA1/WoKmDDQEels9JzKBCB
44sC1XmlfzElBVJBgoJ8C+2hLmnE/Ho0/hKIJ040GmsXg2sXBeoYEMkHHoE6Wc1M
vAZKhQ7NSzN/USptBcio+EURBIXfUKtteN0k0ZdSRE5laM9I5Km2uLAYyjHAdZU8
w+GAART/Kq582iyZ2i9v1EdAAWa3TGqRKLeiLgCy7QIMWmFGMOWJpJIsSBep8EvU
RoXWoC4y6bcRuNWGvqurO4B/Gu/yt0vTH0InItocQCi/in3Ythxx77VQGu+zTNSx
OWuVTHtbmlUHCQjNCudKPVQOk8QMiRzNiU/jGBfhgC87Ms56HcYGWS7l9u1RnCQt
t2y7LH0bORZ4qQDMq/K0bzMYi1Q9FDd6q0pC7VbQkGSdQhNRKXDnGeu2Ibj2Fm07
85rrpdy9HW435xUm+jycSDNurc68lhRYjHlPLH4qbv6ZischoWCqdD5MLI4zAoji
sBF56uz1IWX7AtyeLZMY3LxMYmxRHpZg02whCBgPYoEbxVN/8YUAsOYg2wR6P0rz
xc7rHRHmAbcAEu7t51asHXOWne+/ZEBjCxD1kr++KwinqbExxuQ4OsXZvQkjIMqt
eyTRBU/idtOJnOElihdYzKSh9GOQY/djv+EUN4UXcFyHrbEnMLwkp8xOr3xM3iZD
puVW3Ssp0CXIq0C8cEEWnOxlQoPuh6AqbSdm958DTG55aiqaZ85xqgDqoko/JwhD
oKA3h1fdbvQH42JVf6FzUppBNMwbQ99gG5EKtfk2a30zBC+VJL5bWnbx6/d1XdAn
MCP7pxYB45sWDkpGt3B/xQKKjCl0RsYgEroZtQzUrMpnr5u3GfxtvplxhcYZE+ZD
O3+azMxCjDY/O/acb+VD48j2guArR9hi+avYB3h2OuBU0pPzcmwxDcI9729SWCin
Atz7A+LFVgiFd6h5dMLURSsc44YrKrjlc+lvXgo2YwpBa5pKnFhlyFxkPdRJhIRS
o/ykX/x/NT3+/H+G2VaVUPxIXftspiLFYgxp+QRTl8JVKhIlXy0D9sqADu7t4IBa
PpUlF4JqrGWMQrFtbOJSwhjPhrf4RK/4HQmYCjxU8Wr5Q2e3JS2ZaQYx1GRJ6lnI
C+4sidzO2MaTjC90vDVuvnec/GGd+BHM/B86ImExn9KfZbeoIktxLbKmRAtE9040
sFbfygmvJ6HrCWlQ0HvTyemzS09By9GsQcbDCXJ6n7ntaaTILAkgqEXkeRhIh5Tb
Uh/yJ5l06dRUQZmRsn4A/txMZ5sNVcA+CrJAj0W5lAVQDPZBIaIQjCujipRZXLJ+
pk/1SHbg1PH3SY6gRDIJGFmf5/ZX7OvyPuarTT8Ex5eLqtxITwi4aV7cjLUiZrxK
jUog2Rqfbwx7dfPwBPJUxcpgfIZJpUZNFEc0rWyIurHjmdzxb8y/lVc5y8qTPiKo
NQBD2cjxKX2BgIO3dotyokEuDPNo6jA9guHr/25l1YiOrIIm2dC0FdBKWZ9OD0oP
uLF4SNAz0XTeIaJnP+PhJqApAyomZ0CMXJ1Ra4TH872kVwtShFAlYnwOYtzVWG45
yaoVHuJ8jS/e3bFE2K6G8rXKvGgQuGJElgCgVglfzV3Bsf3q8y8JMk5JIgEWvUF6
Hkb1NxW60kT3G8b4Uh4Cx32HJYBC0DABLFlqcuUZ6+ZHf1oVWt9sORam8ddZtN+N
9bfQ31rM0CZdFIUWoewxG3Wr48zI28tSClljhFEzSwZ1GIPFxfacqPQgORnuI3Rz
l6zIG68TSssbfbZxwGSmRh11daOqudGF+7n6RV7MNLtQMw70lBKiplVraPxVWwOp
da2vPg/CYy/eW2Ig9OFHEj6Zfl0z4IZBuw7gPMfBml5u6T6m5XIDHp2iA6Qbzg2T
dRy2jm4uylhuJepFa/AqFgabZaSDfw0x5q1Q9CULTL069k+FaAGdqpx2bBNV5JGk
sEL2RCecn/XqOwXv8Jc10mXcajAl5ADTZNJpBpytwM7AafUBb8lAo4KSulLZ4rjV
6pYTnf8n8yQBarktQda9LbN83lgh9DKDlZlpBG1CJzk20k6MW88FDEBLlQMoB073
VJJCmRcngHQlW5+Tcs+ToJJQ0co8kmoaZ5DzsibUj10WC4ArLEq6M3pnIx8pl6nx
Kv0fp9XXuNQiaC3bNY+Q4bWxcTK570i2ZrwOQKqXKqyUDa1q0Lv4eYFOX78JSQ4a
6+JzYBJlu3qsXuIR9gZOWoknnYroFUYknWwbA+PM7QLiz/dOjYr0039T87PPc+nx
9SgHAovjlzV75R004wUsFThW5UJYpu9kSPtTzsMZH8p9ZKPOLBsE/yeCplUjInmJ
ToyiKKgBlYwGAwvJ71XRJvUdlsVY3SpzHKaNKu9LJW9nfEA+jNiQ4SWdINsN4lr/
OkkRmNJD278p13J5NyfK9/FaYqY7ms9MI5S36ngsfo9PAk48tGip9KpuVapwpX7y
8cPSkbzUgucP2C1reavbA+Sqe1WiLYcuobtFZfeceADwk5zdCyIg+XpXPGjV9uET
0cI8QDuula4kbz6fZEmtsnqsYsjR12/jl1iYe482/ZsBeVSJTmei9tej83hEl/ad
PnbiYMQTnuAKpFN6vpZw/DMJ15HKehbMu5AQskVtNmh3wb6BC+0kkSxGms1wZh2b
vnLPz6j6jn2tzvjDC9Bdo9q06a+zNNt4vL0typRWuhFx6ViS3csxsQUTSQgTT7ZY
XNaiDdPz5cEtnx5rFiHzTOid0Quf8LyrG5d+ncfcHnkNVPRbspWy3kC77o7Goa0y
YfYKkqEqF5/nrfsT+rf17M/L+uLcKqDA4cE3791Vjedn38nHfTLRq/xo4Hp4LFrl
Cyipoe7PHgvc55IjFF9rfgX15efOjN+TQa/eedB+D+FGc1BunBltqWwPvL6N9wLX
65EHjhQBu6Yozv4M5EGtQbXSGb696FXIPnLCZA9nJmt/+DF7RZlfUd+YmO2RzzTN
tiOVsGLJWT8Tqn9cIJcA3hmP0w6eCSkIS7rkC7wOxjJChF6zkZ3Xptop7bk2BKDz
rjO78mcyWt0X2qq14B+cUEUanqQVsdinrgVj6W6H97QKCCWOumEauAZEridEOoUM
jywsHXlzY/heMhcPMo4gBg8earTL+Df3ameweW+/QLDq4XDb9SViDBe1aREt5PU3
X5agSeEmF06hJOM+VcurBgwY5eu0hj8IA0BnyNfFlWpzZpPKEY4XwftJJ6LYBF+C
+unKRtoPG9N6ABp0QtltM1+aoXlKL9obR/lYAbTKrUn+f1m+pZTy+tocuaLME9qb
w2k2dlwEfd8Uxd7nE1urZT+h/3kgR02suw6cvbPS227nAD2lJtEEgzNYgymQRByq
tFBpNZwCygePXb4mHy3lngYeiWAotrd+6OJuiy6cvu2vH9WvAJaXcEAlxnPW3vOO
DXYjSWkZZ/SBpCLjQ6FV+x5C1a9t3Y4PZkPQraWcddSkimxWhDuHpfSdFyEh1mZ8
41lrznkVNvHF4c+vOC4kbUf4gmW7fvHMTs0/f9wQDgDCgIFFgMTndnW8OGYQlfzg
YbTYzLkKMhNU2vGkQ+IDKRBZD85oNYH08nEc9P7Nknhbz9mC4Yw26l2NGMru01Dz
Vks7WQRfx/u98K3wO2DIOPha+Mhmcsh5l92fpeGwP/P/odMHyfxlIAVe3yl5oxi0
De40rwoVw3COvFyqw59+Imwpy5OWWkScdrtkT2aponGwW4vHEM2aUWAiL/xEWbGy
fR04q5JqnluwV1vsjaw6aBTonfHhR2NKnof1S8Ij0coY0wDLsE7Nodmc7MVkXHuq
7Vau89Bq8rY4C0hNZZzAtV0RzOpt+cC/6m4XrYpp3I5vjUfuIFfZBZj2TIB4IVrH
rxYb2/KbSS5jYFNe8O9+q+gcM3hfmSexiNEMRrqjBB4+2Mf+8cD5ZA4AuQZtWVOP
EiHG/ycAA5+SxqrNJNoWSMGzwpWAQj6R269VGeMaLl7OwVaTN8qYwwjtgG7Ad7GY
p038sfOqY07OY2ztFNPeNpUWfhKTKEW0HYxNSwy20O+QlU/ub5CPtxTVn6O2zIlc
1cfNzxR7DrscMLaf/qmKOwILpXCBi6kHungINkG9PAAAVy4SwJvWN8w4xhFxkgTS
VmoTAeZcjo+6BtlElEzhtQMjwS9O190SLJYLKTL9chIJkPvOREsm9WrhgOEIVYYP
W1J8va70yVbvaYDicQem/J8oj/ZqAqWrr/M3BSckA1V7+e+o7WSwF23em41P96SJ
7u7+quDIVLwPESgbqON3S9/GWVp3iblv9cgkRQ8GB7v8eezxfL3dSEaE42ew1k7k
E+NxaPjtDeaawgJMCqkbv0BpliTfXuCxABfLC/feR9e62FHZ3yA3Vo19EwEOzz+y
7/dJmD0rMxRT5b6vebF22Ez25v4/T2mLmfrDhMmS8hhMcOCuQQAcHft+a7oGkcS2
c8Eo3UikLPyFMLqnqcG1f4WRj6I8XNUWrcbHOwYTR3kPe9xPsxsLRzyatI7hbAOc
Wtg+MeiCeUJ7zydlX9PTVc2OD7UqnP09a4qCEObgnZhRA4KucaHSjPuefgulJyas
hr2nPqczTnCtywfFNYgj+ES7o3TKgZGHIuVD+BjjLWIBAt3BvEglzeysl4X8NsP4
kwZyt8Pah2vsGNEFJgVz3oof3GRr09qLMS7ezU3xGYzte6Izqd1WjqiUL7MnpLfw
co6a2e/2ZkcO6PASxwVIGWPQ5VnIt/KXD4erYVPlOpiadWVR0t+oqEEosxrlAgGL
heg9yEK1j/wMVdwn0hsx0EPogZD8tF3PMkIlNcwEJjLm2v0XQUCyZhXnmQTk2kxa
x4pWx64XHRkhi/z/WuucbjHLaMLqO/ZvQx3bQux/Z369D4ADr0eQ8eyjxUN54jOk
lewE6YN+CB5liVmZ4VjmTQAMy5vaAjghyiydveHjnMSrKK6i3nUKnGSyn9D4Bmxe
CvBzc2t4T3t22NEVRbJIYvFo9hy4kvxaFbf7FmdXVNjuUjIrCT+1kfENNh5Vdp4M
0Gquk/IHDN/WFH/tDirXX+2P7t4hKMXD6774IFBdoV9cLyYfbM4OUh50msDKV86n
lLOqPBP7ozUxrU+e77pGYQA3xMdzgGTIhnkJ+CbDutvR/FZnkJYhq5EYZi9lACGn
7OpMoZ44vA0BaCF/jsyq+f+fubvWKU0fr6YJkwsBsVbpxNjdhPvqV0W0KnWw6O8q
0Xd0RkCDmM+V49KpaIwf9A388bn6T66JTtcNeIATwH6KFVyWt9lo9He/EwPqTwV8
otm0FI/eu5mjNs9wBNdJwQ/ZdezJ0v5CDA8nQupbYsB4MlLgrUeMUir/w9VMGIqu
WnhL6jwLDP6Udhlarl+XeYybNXCM4p8y4ZSxV8TbcuM7inIR5B7TtVSh1Z6v2lhh
CVzZe44LEXCeoTfk8oimbsFIMiWX0PAbH6aUcBXFMvTgVtQudZbQK+VtAK2kCP8G
Bg7YXPB8cA2dEBV1It3VW2pDv3fvnm53iu/HmziNCZ3Wux8kk6cnzwXEMpk4u+eY
ywSZQSzKAu6SeCBDjmVPo4nEDGCFSFfU6TOUA0qSSeTFlMoysyJZhA3FC059eJgL
IGCuWSlM9ee7H6mp+54wQSNmMVfMEgJtbvPxP1w4e/z/ouZdNPBp1DZbXXiyz4o3
Fu6kmZYWpIqolsdgrfh+RwdtqLPf3Hm/q/e/6dV+bW5omcCaGhZnoyZSxaTai4B0
Nqzh3Uuxts0wGbPb4bJuIkTKpk1qkFwWCDC0nJnoOoUL5lmzGgMVN2u77YR/n90C
YpcGepCJ+53r+AA4yqnkKMLkCKrwD5Roi9F58nAzIDd+4deb/6kH/N0kdEeg5C4v
xHC5Z2V8A8NS33y6CZtXzBea1s4BZLsWbNR5p9YQhd97Fg8COUcvJyMtrIvNW1PT
MyqMy7KQKxZlpYswi8/KYRB8yGKU1mMQdo08ZrEzoeoazVAg/oPdV8BE7XSN3NEL
8s7/hCHYNf/APB8RYJ1AykU5ora8Z/V8mtFDNZWuvIHquVXSuTpbjjwvTgu/Vn1v
MygXTxC/V8+ldcduvP7Lxy4zU6ZSCTszVPBn6AyvJXZTTyc/FjmU1UJob/tGPx1F
2IMPXjPl3JHKJsT3Xok1XTPUNcrEI+0ZapZ//WRcLq5eEYFrSS8ZBfcLFpJkVm94
xKAmZgUwKEIZl/zfNt4e9ZCjj1p4uEhZGl0+zIUpVZZyfeKFSG69FSgftAwMI5lc
9ahPurXFlPFPlF/U8p40fPhuY4vAnlxEBQktxdJAty9XvQCgYN8Zo7vPTQmJSFJN
gCgn9Fz3ilJLIFWFadAHhY4iVrvrLrVmfLkzg/YISS2EAE9btnrdlyi8HKaZqwwD
7WIa7LdrA5CEYJxq4D2WaIIBU1w+UCkPW9/+KUJ+pLr1oGBMd8XSj4y8F27Ov5IE
kkUfj405LMo8p71he+V7clYJjVL5SY/zu7hBScTMrkvAXiA08ctdKYQ8ki0MRIK1
hdQWa1ry2HRbtjGL2dEQoSpi5OoQScrVF/WMHd8nMfe/Lt9vCcBkCy2tHAi84pbC
unURFT+aZTJUyFmKvdWcUPVFMQxerONrgUKpQdI9Zi02c/LxYBex3UKSvjgVow1K
sF9d4NA6+K07IxWPfNnXQlYjIpf784k/7u7pt4X0+636YXyWgkzqrlKRA6uy+U6Z
+NzkufUEiX2yTAXeKihknHjIfzEvgCAmmn5vaLhy01/3HBBs8jK7Qm6sYKqkSTF5
XJFZN3stxp/rtYyIj5ZzbQUGvr+cJWDv87Wgr/adaA7GwH+juimZlQ6kpXxFtpFr
nAI6vw/MhvDvev5kHlVxTwaxIATGMHhJjv0BJZK5fvkhDWqTkmQWXRyNWqRh/eO+
H+CBl9HJu4elTCnbePYa3W7bLU8szz/B6UNWhYevgD5sQ3zLf6AvIm9R9ijJETXZ
gtH0RLSWcXvh8w/P/oix/SB+jTdGugN3RCB7WHFYx0virdJZIAuxbUZken74XKdX
P+s/me7usoa4T600SJIY/imF7zuvDc2YpN/7t5YsEOeX30F9M2H56F7HtGLSeTE3
nAH0NWBfkBryvcw2A5EMJxyO+RbaRDFHgKTXHmgEQKhrxL8bi+Ko/hfNWHV5fdSk
fofO2v2Z0ON3yrIRBCJzUZCeQBNBcdQ8ByzJtm3gb/HBmRCbQYL6PBB2Z12P6L79
/JqUxgZd9Y6VgWoGxmznFm8okopzO065w9BgFMgGFi6/td4dVDK86eQ9IsBbyJ58
SQ1dU3d1Q3UWQpv9keLIqFN2q/jScA/CQ5wdU3CBTcy/FE4I0S7Pr/DnQHFa5pr7
YJT7I2f3KDga3Ds3NHFggVwetGSBYb/VIGTLnC5rrzVhpzLYerjMSV5bfNsh4lFX
yDV5qS4liE6j+Mj7sAS/Qd65zMnEY1QmpkegkcS8Y4qyBr71+vQRckELTv6Tfypg
vE2PaY8o6KmRLKtxO+Zk9z2rCTEPLXGzHtlJ02Q2M5x6ySmXF1eMr8wC2DBNJzOl
kGdDE1szpYrJ9AnKKU0GQfyy2BintOwN01UwdcvhTRAOO2dTaUgHWnDBzeYEfi4/
awZWXhs1AAgWfLIwGC6AzbFDK6wwOlTE97hMc6UjK2MAbik9YPaGy/wuM3267IZW
1lpbtUBK0yAPLhdm4l1EdRxLu0jj7w1PP1pQcaxF5Cpwveyc+v3SEPpU5Sx3Xlo1
3tVMxdIHbTPidMZIvBA2+teA2Wsbnj/3KGHLBxQeb0rkO/4uG+gywFBFaX+Wm9ap
VlW96gcRwAnT7CX8Q1h+Bho2cPr2cpkQA3e5BxIt+dqJSrVZmN7j6kMYSTeFzj/k
RH/p7l6jvCR2351b7FsCzrPZ7EVOPiQnbhHZl0JamT2V/tttJ+rogR+HbcPLsH4H
xxnOU/YTV3fHH0xFcmtr4oaP7jlxb6yorY2l5pa2G8VeYo6w50/gam2TH5Kcijhv
wmlbIVn12889yoPB9CusCRypURjP8vbz1SajZEapfuTj9z1fXSkFnH9CsYhbbHgb
PtgnzHmQZjT8eHk5Jhf3I8uNWVykPSKpsgrVMWNH5KeXEZmEwej2+NfgRDatdcC2
GAxZb2iAirUrVX5u3OpuxIeQ/QN8295zUhsf6dyjP8rK9ZIyj72LWBbkAMWsjT6X
I7pCxb4IbSykBayoz6iGna3wfJASU0xxkp+zuoy07kkuV5O2n8C00o9bY8wlX7JY
a/hOFbdhJTt9edSmsGYP5+QvHX2gqHQV1jE/0YM622q6QAkRxd5aLsNaV5+qZudy
dBiWsj40yOLDN0PiAvbYfIDs37yq6o6el8T9qgVV2Ia/Rhusn4tkgtREcxUK49xL
mK5kUP80TiqDeMDdcSZXr73wtXdYVBHSkuGLpwYo7CI9pYUpbWKYkgdcakH6C25X
LozaizdINRbKJLs+ZlvVK+lOD0VMxROUThelNk0ekYKYD9sffnE/pY+XW1B7oahV
VGtSKRh77cjV1d+tpOjaUd4f+ppFRcfGAcJd7bKwaCxK7JTVwe2bOg6oFaz4Ca5u
7jPEfElVySbe3kHSLj49bhiQm0Cbs6osP0pNA8atTnbT58xkJrieAj5ukMVzTvMD
d0m+BzchTj7vpGZz+y+jgcynwePpMmU4nI85rshKcegTfFKAq8sAKQWBcyxrbid/
9rrYuXxaVHe4ElWuNG90sqBlztGLkxGokXpEKoZ1qzKeRnmSsmrClf4yptV44yVH
IwFumIzgOE7VkQ9Fcs5oN6tfwNuvTYljNfZyGycRxsqA2g9iZU+hCRf9FIuM4rKY
f7PDxPJY3PF2/9QYPN4XqjLaeKjudCBZaOagviFuQfIjBR+dG0pYJVcRIeZqkCZc
OAM5wQB8DIyyfFYVuJtJ3mbNqMvnR+fCKn62P17oaTNsfLV3zNPIwXtN0dEDcXfx
0Ll+q1g/lQZIDwdIgdoGiBcF97+U5G1ylj+dcHUXci45XglKTqRlDGvCjN+K+eGk
50Bws/hkPnmd6Ausunlz/wMB/5lI9s56fvfmDqziMS1X90LDBspRfKelFxe7t+Dp
V7T5WeMt1eui7QjWwxjjlb//ubvl7ATKimU4RVHkR47G9FWbyMdlzWIgOT+jcRNU
A/uIMf9Hibh007Ei+3hQW4Ws4tjjl3BLLSkS6fYLht7dkFgShtfkJ9sheorB0fMC
n4fK94nBzpnFEhwA1u4f/vMnMxli/esAYKppf156mKnsnmeIygLN4G7jahJNwG67
9byYJYWr0Je7EP/A5f/n2jX88jiCSULCjyyCqEtQHRcDQn/n0qmnJGbZIhBfTR2I
GHPuxCVxXE44GQwufyKmcUg/SRcgPyFYAciLrP79Sl2d6ozqIvWQeRutWTk5i5BL
9OBLbMWJZM4m+StdKDMHZJkbSXcWlgw8DxDyJDioCRBzRBfVPHoHj3pAIJntUbtb
NdMdeY1bkq2EnXiEh3lyKI+h+Ec/3KeOTTM9Ft/d0iXmF0b22cjoLrVricvDnR5Z
o4YSHQsdMCkzeGQ1v0mm9IT7Cr9iWPJkjqasS5AfPfD6APvlRFKLquy/NuDRH12Z
g3n/8gTnWS8I5DVd6YEO2iOUg5BjT0/lwgB6VQcUnO9RphKvTumlEeDKqHJ9XO8f
VXp2Vz8/b4v3GKH6NaaJ1yJ5UwPrXjEFs3G6cgbdKFJ3u9oSGRWgc6H+H5t/FZmi
1vcDtrethpyzuGSAEbYDxAr/xPIxJxLZ/QBIvR41f5pe7I6a2+uqm90pirdodEw1
QmhXNINU0TXuW3JoyrJJ//sM5La2qRrkHCxYNabbBhFhYlNg8PHpdT34m54uE56L
PLnmRb0HFRWCI23XRBd+9zJ5OAL+V8SnuGAnsASkqiOUH5jZWTmH+MK/xqsCD8yG
CXY9XGBEkZmCBxp5cWFrW8288G6nvBrmLuJvJEq+S5KIi2IuPJ+cJ8GnEsmTnvMl
3OSjibcJ8pzQf8tvAa792UqoY/+MhQfo7GN7ryYSXPy6Vm0d/Uhymg3cT9YdoGDI
+pvQ7e6QIy64w6AnvSQW6IkQ+rLA8OrhZNFlhX+FziGCrqgElV6QZ6SRj3PT05z7
5KfIWvMvOm1KbYUDNH8QyuuNEGKnb4W7RNaTkzOeM3m7X0F+CzPEowUEuwiZNz+C
YKLGsScvixcxt0NEQF195P7jwLxAZcW/vXphUDPCXTtnbOWMAzzMWrb8d19R8TwQ
XjhZ6QRm4HGvd7qKlUTGFPcH2j0J3UWddm3SsleZVIDzNJCig1wQLeYlSabqI8bA
NOrVnnVUYvAPYPdshN4Ba2jN/HmQiZXNihprfhtXpFFu4go9qGwF34oHhzWhf6ja
Vn+OcQJ8WpgG5zvu75dze1gJ1XeDKJ8VebrEj6gUmOhpzux1p0SwPjonO9ZvQjCl
BCdSTforO4x3D0yrAIf4d7p4NUSmIgrPX2j3NJk9YuRdSPV0PfFoPiJvk9mJ8/xv
CYryYEzHkRnAQCWiU11Os9pJNFZu3M0FYvKsyV8kWMCy9DJywrI5bbNXUU0d+wJT
yYNOX9dnPizXrkgdzuDSyELr7JG7yfLyn2GDTofZ2t/glTobMvx4eVBW9RHmPeRp
uOSxqWY31U+4ZyjDdvv8P1NjFTkdhMP0iOaT08jophjONVPS57i2zr5HyFYqMZft
HTjrD7rzni7qmx7Xn7eFoayI2ApMR2DoiQX6xSPkOxVhB0/3C7S21o/BaENh5q8O
n8hlSib+zyKXXhvNYnQcWBSk5DcRzZx/e20Iy4vZbt9itOobnuGeO8qFjKBqtNr5
16J93tFSvuq2n2MrMdXRxT4dNWFS1R672N2Ha4rkYszDeSG31gItKAWywqEFaHfK
fsp6yp5rpSs51aOo7nHD5WpbxE1cxmRt4tA9idw8K9KStw06IWKunfbM+A0xtCdC
1jU/QL1xi3YlZ9qMF1dImN7yQJNGtUqKOB1Tateyd6ZJ49dQfYHpxVHz4tIzVF8k
pGF13cmIhozw0mzRpsvROnCdEAq9lD3viWOfPYj6ZXGQ7H8bdXVNf2VjA2oj2BaD
s97z1RGVzu8uvnLnUyBRJ/Yv7cjTCs1LkU7jYuYrLBhSTjJOPqKbuxXMXoZqsLgU
W5MwwDNq/B8iqwgOL0tJyy8De3QpVQ5xbYzCniqi4LClCLZ0qwKhQ+xVi1HMYvlg
RcvvmjFvi3EFR7uS9kVQKwFtH14/Kls5R2ZnRhbUZu/pzih9EN1okpZnHM+KWqQT
sEr3W08i+Wx4DTqfTIOFI8D+hP7KM0LrIBAG3pl+/FNjkcZ2J1fcunmbYGMN2O/k
hUSReNXosp+tL8XMhi76jc5sqbz3xv0zuDU/edWhwI5K7iuc1ijlyEAgN5mU2DBJ
J8zwZxQmLOThod2tgtdkBd+/vCuXDd2pQKQ+AQcZgb0F3y1Zd3ojDFHeeL1n4sEC
fTekB/HG/giItieE+czOPOWwzyR7dZOWYZ2PWaaXoE1H+u1mSlyLt5HfgPqx27nb
bJK2Dwepsjyf7XMi0vA7OlPQJ8zFsFyN8BW88w6fX2askl6Ug6TuyOM4l04GCrBt
p4cRdYUa03uajTYjAR8U0dJzbKK/7lFfJe9nrbfdmIT4dJYodjpRW+AokinP+ofC
iyRsGOT7wQ9DncjHvKAgy7XZ3xJKQybpSYMWJCnUVLscrOZuCHSgHKGBLmqS+C3Y
h/Bk5jqCUp+VymBKgNA2vJWGJklUptj7k8BIUEdnDttmUpD6UYOjnzKvrdRDvZ5R
dTTFh9VonADKlJ71KJqBcqgEZmA3cV91tn7lUd4xBN0/CooJXInP8YSEFe8/nPGm
dktyc1uzfiK55GcjnAv5hg81fHsjMEYrRcVQqX8X/zhE8z8RD2zXoSA8gBhYnuC6
blXRpNbOmAV7TU6L3aqfg5BylLkgKUJr/hKnJdEkD5svVh0S2dfn7irlc6hqm8Vj
dzSxZ0zdTu3fSvo+s7oc/7Rctg/Msl09y81aOsbedWb0UKnx3rPqhFhDywneK3Tv
cSeilBSSsCELAv5sBqTo917O67NRP2amk9RgfGHFq0jI0dgJYZ/mWPqZe+Kz9Gtj
B70QWYl/wzP6FY+12f2I61jwxA2aIjdMWc668SDROb24EHoOwvDSmWB7PO4j4pdt
++IOJWwDEG3W0sH2vaDP/8ExMLXcmkV8fO2ChpA6nWj9vQV/s1JMrxzuR0eaKj2m
bqd70usBEcn6P/Ks8M5NQ1Yvey6f88D95QVizlTz+tt85PQMgndKeT8RwjOS+7RF
0wz6eafSSy2ozfcRMROr/VMlxqqC5cZsFJEOCcvJPCmKAL5SKRE954hFJ6OBiJdo
yjWAcEzERAd28vsYFIvTA/wqYGmV+yboEuPhky1ZMwrvKWw+AAdgMqa77PNzMc/3
f59As/QoU/sBcONyPg//GjJaEfqtrRWOZGG2D6mNEg5Dh0QAmC3aFxDLu1N2pC30
3rqbLS9XpXhGGMySAAAeWnQTispGue9SEV6tD52j/pGSnB+6naaa6xUjI65Isb3h
IXGHlP6L6IX0+TE01auxIGMOlalgTjclIFCtHjrHpBBgOTfHpPhfyXiEAButB/qS
+ZgWAqqeNGSyCEkF9yHfKyndJ1H/tXKw4i/Py+VyjfjYqbqfUQ18e2PvI/LFnPE7
V86ZwMj6pQa2zMk9kMcNX0I8IrSa4kmCN/eVoh2g07DHFQa7f8dG2bJo8SeQH4fB
BFK9ylw37vRwGeGjDfde9lHykByMC2qofH9H+zz1pr1nIMzcop5suXOkNouLkkvg
FVkqbMipPt4GRCQ1xwRSTS3f37OCWiGaqHrIiBPy574NWJfESiCyQor2B+DovOpI
B+MoD9WHJ9It+a7VJxew+iixKWWTzBA7oHdAyI66rZCIQERDckzWlnTSXNFVmpMu
v+kZiSUctU15o8DTfCJqi1FBMEu9MYONOrHLOpA14qacBZ9+pW/bYLj5W+D5jo0W
1M7FQa8BF8da5ET5Qy9I3RsLOR39HufV7cxpmsiE+gVl2LSwe8tUNFm+IItBF+qm
0cZ4O6CBfPNeFdeuBMZg5DTgdCwEWTjgUSslna8G1LMEuKlzfuQdmuBqBj2l68Kx
xLtCizFtKBcaq0xx4dHWoNB+zrsGug9LNYzZa9JilciQtQA2u7VsJSgo6EF0mACA
1Yt8MLYqal1e+As+toTnL47QoU4NBbaz0lFhleBkz3u140f+bti5S1GD0doa+y/w
6tlN9Os1wsC2EEFGgw+iHrONd3ZFM55KXJAhfarnrkOSbGBWuoBnSBG1UG7Uyv66
IPSwHw5+Cbu7xeLCYAQI/aGvY6dUQWcUzKJio1GKKf/ZV3IpFgtvVsAFf+VNo5NN
erBDyydbl2YFSHRlkrAa2dOn7emDyLMlWl7y92tERF6VpaZwObQizeoO3PqtciWF
dyLvIU/nMIEucWVIYrVKe5DS2sFzZvaJrnnasCeniztAT0cnSVbM4f7KVeJw/rS3
xr3vxWqGSdS8hqSoYsTMdf0ztdZMWZAV9LCkJ4fAzxUsWgcJqAWgFBbc4Zq0ARfB
c6wm22ot4gYNw5YzrtUaS+APX6ZQ0h0tjpDYeHMN4FAQxAqmbrN9CzAYVhuCxR2N
2OWSuAiYH/lP7HSqpPhpH390zoO5NuX40pWAIM43U1we25jqKaBgNcSibEPemKiQ
KVDloIxsHyQXS4YIzESZMLXq+k61T8kK+VtNO0hSFrVTVXbuv7fMRoeoAfxDpcer
3gZftn9oY4yVpxJhdk4IXyq2iVGsxSDyR2sGxS6TdTW5EyAN67ax6/sSkGdTpvIR
Suq0VwLcz0FUUsE9GEKV/3M+wrlNzkP1ipHgjnrvnBvNbx/ueiA3KYuCCoEgiOVi
dD5lCSIfLQxZJUyLcM/MRbqIcU3xaCoRImIVqw9jEj9FsKKXFzA8JjP/5SL5Maru
cuM/5m7EBzAfDKLpO6JXPQ==
`protect END_PROTECTED
