`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sQmaxCvldSKHa6hxz/1jw7nK6BfTfCZ+JG7C03YvIRidyPsLrHa6KedM7NdP/L+b
sBdoHmhVg4vU2u6X/Hf32RGmSOFHTeofEW7JTZEfBCdBhA97FieFfyXb+NCcGdpH
jDrzG0JjF/GfSZKcBnqnrBZQbcKqxt2/WnYHcZVXhbW+KLOEt6lkpgq1FFtadT4k
SX0KgXTPnL5aCy2p0eiNX6WQPQxjlRHbD3V1QAb26HntSesqacqTe/mtcYbtBdxU
IG8bR9jB2U4gMjQgApjXY9nbYaZS8I5W94dLtXitYhuIft66JoLLdxuk5AhCaET7
/w6zLzfcHVKzgA/Kj+FdZGgiWCSUBkS2BmN0BiaWFyMQVAnDnXjFbSDKocVKzvCs
RLpxU9HODAFfFdxYiiDZYg8YpsaQVcITRnI+EA4djSYziPu1o1//QPp9VVtYWpA4
V/kognr4ZdBCDm3aJ31S9BbGxDh7JvUlpY6LeSfwWaqDDS0wXinuYTq8YUiJrzbj
+NdfZhvreF7zd1vIkG+rRibBl1I7hH3VXeuFi/yY8l8Xu2MQNSP4DaDcHFy3OBCR
pACCkvAjXKXrpi8YsaWx+Sc3flSjgCSNlJoX3f3H9ibe1G+qr+Hr7PVM+DgMttoJ
YfIT38Qd+6zo0XP9/Nc7yT47WZl0lwqFzwZrASllS2+TOozAPrserHg9ELHc1+z5
a32MG8uMO6utpS+DSvYkkyetFLne9LVLZSX/EWwms48/VbbNuEtFfTZZ7tXL67Pk
NM0kSson0OBGI6MqdD8MUtbzov2PEMysSZJjDFF66ItrW9aTU7GIDnFFJpXacSrE
54fGj6AkbGVkCAAmkVOsXBgBP2kDWUmeTHFjYwQUL3oEPavzWAvQaWBvmFiRW6kO
Lu6u4oLELJH6l1iK82fqX3KH1TNMJNgeZSNebuotYo9K6CyPVwDpwLMnNhhaXMuQ
5pUuFF0VHVoiwTk/ZfOJYAeIk9vwJ0eHNGtlZ7H73PheGDnCX79pOzRUhUiakJNx
KmfflRpRhyybnPscAtMCHkA8qkg1X+2Z15P92nYdbuXX4ZepA/gMbfgEqrf/Ppuc
OD0o7y8JmEsP+AoF0bCRMqucA0g7p/MMDm7Oo1RALyv37k9cxmQpKZRMFrSuMgNj
5oeOlrBHoBoR7DILJpQ1bAa2xWH/ik4rJFb5+/uzSr5Bz9TkEK0IEsSRGCuejeu0
lFYurlpMURhY/dHe/A4QEsjCKUXHvB/nxPa30i+uQBHqGY+vno2oi/XR2ZW0f4S3
gzt4NA5elY1ESl0LCW3VFNtnEwMc1OSm6izAtc3u9URnzUfQwQvtAI1iWs4HMDGx
/6yb3OInIsUTK73cyE7ZI9rTY4mqJMH4S+V6lBkNNuJOg6O2IExC8sc1PIjKR182
/4dFmQPND44xksnsXnreNwdYX9mirg5ywmUqsXN8kKEnD91Ay4uU4RcWiXrA/My2
hkegCGGlTK+9XFik3cIwfjmyyxe02XInVh901pYf3uLeZJiRD7QXpa7QyfbF6iGb
4+14A6MV7OdTEoiTcvi0S4htfeY8eytg01sKgMvJJAUcAicVpea6T0WH0qcXRUwL
wpRunwXIRiZpsN/Ar3/FRumyZ7lHkEUZV0CdwOlzfD3D4NAsjd+GQFPSm3ILCgSP
/JIuoDimX8+T4O5d2eSpR9Jl/XHvg674nOHxZx0VNf5ENpDHvcQoAUfskE66TEa+
gBcskagXO368a4g+hLm+RsYLe9FocPFQpXAijKZTA4zOfsx0e3xT4Y/zrhiY+jdK
8hfUDbFAhLc41qOuEcY2tAk4E3npjeVVFUY2bOa3qndiK6N+jnFJspKXbu1ia/NQ
`protect END_PROTECTED
