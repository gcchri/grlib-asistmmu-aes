`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cF4StYXP+iAHl5i4s2j8YwjtVbOOVNFRWkhmyEEZQj4Om8Q4ZlSv8zanGV/Qjgpr
F5T9oT4ST1FN01c2eyDhDtjgXzoSw6kA0pOvNbCaWQ13+ko5PCYYkNXIgvkS/Fht
O3FvBrePjlz448E25bUPR1De+6Ly1Pen8R44WPk0CiSeAEhk79LHhBR+CefnE3Jk
pk4C9fvMB2kXphrxZkq/4h/wUpZ56cerAIhHotKEu/uv0WyAHbAPAkTR5ZaGvQ87
OsXWMVPI2dIPr7J14DY6XkBhcUDM/riLZwGUIP6rrjzmtgHGdxlbNAoE1azzVdSe
OHovn85BlVQn0RcU2NSgGiteG6QwRCRNkSZUnuKhgUMXygrSRV/mOEWllJqYnWjj
93rZSxmqjvCS/jtC5jO8QydPJtUoPhfai97CVvU+E5xTTdG9Z5NP9ZEtLahZ7sU0
cg5amiBBxBbMtZV0IS+loI8ZlHztWcwuYH97aO5H0HBhrTS/DCHjEext3JBB9I1Y
zfnowOi4rLLoUa18OT4ySg==
`protect END_PROTECTED
