`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iDCCsnoV5LCzBestMdyG6iA9xuP3F/7j+qMQV2NNmNqyGQWYbebJs6Tjo8W6Ek88
3Tpj/3+l7M9OrGI4c8vxd2BcAcE03RgeWtxtyqUYrE3fahMlkoxG/BCKpKYSOAX3
0X8GiRN94jew+kP+WryLAsjmgDv036pK9KdfVaJHoN1dixyb+6csgvap6Do4ghBw
3mXl7+QxOOPQHQBxsiy4w0kPdCgAlUjf/1F22Jpt7N+Y9fBNvhuaLG1fIobxrIAj
9+HTywUfgEBj76gVqB0vkg==
`protect END_PROTECTED
