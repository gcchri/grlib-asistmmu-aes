`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W+uVnr4/p3sWHYpFMSjYkSUk+9IKTXCjRhPzCTmq9DhVxh0T9wqnMpHwtz5fn4Mr
26qm6RlXMOp8PP7oXT9hEAVWKHxpyvlS1hrb8RomUQZ600+LUmQKkeWNkNiFOf2T
WDrK/gSxOO0MRG6HJHb4rcPZ+h8lcWf1XV2aIawubAXYqgJyNAXxkItinGkCF+d4
+YfwYsZsVECIKJ0NJjZ9XLubIJ8S9qGhF1UV6fbQsoChNCTjoMntCnd541hA7wTN
sNcG2Bl6VisTXgvW/LRcUG4D7qomp2AxXMv46O1OwY8kPkHNETGQzf4vHR0mp6Mi
/EKepT38fu/Ir2iF8difAKOkSuu0YLgnfTljUEiyIzRMW13LMZ/j/0LHeDwwMtTK
ySl1hmo4qsrubIhXdF4WiOL7+QBU30wGE56O/y2dNNbOeBreDWDzzhImdl0q5ebO
fyWisqRjyR2TYOrIB87LiaX2vfTvp/sF2usmF67AyHJrdkJgAxQ76oKztZ2fV0gi
2G56hCKSBzjgvO0YF5HlZan6yu4fLOZsn1en/p+PUVu6Cs50tw2rhV2p9/qkTx/k
HgMgFq+1jP2gVF7b8itD+0Engiv4ohsJgWQfhXTSoVvMcuCWrTsA9bwTYhgycGPU
EntZHVEdqOL6lWnZ7qCByiti/ffUtEtNVM3xHkM3LFlLNx/WPJeBBTe13uCMVqbC
A+CnUxgFJsqFBjqr20FRl2PPYalcii9X3nmEYFqPRDg8wLoZ7HG+r1y7xWKg/gXW
im9kAVwHyoWkGT53fzV8wzB1WXJGXKOzZ+GGTrCuIoorpRdZXj9u9O7FoFCKYp+3
Nrie28wNQn2cp/ooL+P51otuSBg2Cd8/6eVDeLQokuKiXw87TItvAUs8Z9iO6iOV
34YL7fzAy4/Ed5WGrPzHpUYYUAF9N0TXI5cb3W5QNG7GKr3/I4uVfuGOgwkMAqHB
GDuqXTO49f6eg/ulP+ROfcgnKDU3MRdO0OEBXpZgkzioNDIkcIRO9fkrtLRkuIS/
WMWVyyK3JUe1xvKuLUc8ayu9xfOAhAGCEdshDkWf9Z3wu+O7BcpMqj/JWRFFHjVo
CxM5+OMfuFEiGQcE8+KEF2m+peuUvOo/oQP+AjOlUNldFKMKbVc7aecnnwSUJjHW
uPh5JdThsowlBVYoktYedFktb/6vAIazFnjU6Ui25qeW/VQ1WUzQUwSR5I8F4hM6
In2EyY0FjkiB/etFwl0AM7vovMg92kUfDIZnWT6vgWT76UFKvFIpFclQfhUSk1Q8
wtJmLmNLOwJmtnQ+pUewbZh/uLVMFaafJVsts/EoQpFzUYJMhRA+x5uzb6yBMkwW
S6zNUR1K5PunmvWRoobZ1VVIonJKYaxIH0rtIwK/xdc5M4wVbRJSRXoKHSUrLM5G
N0HBDfIGnQTVQLIoMOzYUALD7g24Fawk7Mnqd2PxxyhkuQt5QwIPab9tMi6fGHZS
BCK60ZCFLLZw6F5+UuOwTM38qGTwFyI+SISnBEVVcMTtPdW3yok9Lw1aZnf/dClB
x173fFa4gFgoxFj0YjEK5F1XdJFSEXFkjDOqOJJOnqWFMcgNx06ICIfuAj5C28oF
EJR+fqi8b/eX9zxQESUCUEDdyV/62JUF5ULAVVU6UAHL93cop/kUnH0WsgoO9LLd
KBfN+J9vvnrAWfYQk6Nn8MMkMo5OnAG1kpc8ivPWQTrp1R4aCBvH/Vf2rVb1wDWw
f7Y/pa6wTsvjyJOLxmNvNU4C9mvn784WcNF5nlMflHmmD2ntiotCiVLmgGjVLkVJ
WJXIc/QSrhlUUqpptNyVrnomyzV7mtuaYHc3qt0hC51CEAZx2so/s2iUd444860A
ITl6mMsK8zf3lFp3Mfwe6UlH2cnbgz3GFGQ8lr0b+/ZHWvmqcgCWhWnX6GkehoJS
4qECMWWuTemPM2zAZII6yYHG/PUoBx7jwuAke0R2H82ovzSTxGIAjUncsuHC7qiN
EtqyAS99ns6RUbgL6GRS700lFM93hiepPr7J0aVQwIOG3l8gONoImnqlftmEuHZ+
CeEp5w/G8e5hySZkGHF8w2sO9mfnfwGGSzLE26FQ7AOFVFgz5TBjLDCw4pL7Xpaw
I1TtydmveCUx30F85qA6kirg3nabruiTNVL1WGVSudTiR9hxc4WCC3Ye7RFj4aq0
E0jR0JrHbCjlqVCFLSUacbjNDCSIEhVHDhO2kLtbROFLiP74GzkFkMxioRoDnZDk
5OElziAQhQtAdsk0C1K6pxrl3khXO1uAYzrxRaROS0HU7J4oKmM0L97fiyRiyifK
oyCaW5Bb2jovyfkYnT0++BzMPF+aS7TtcwOfewjqgT8=
`protect END_PROTECTED
