`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ST24FvBjS5Xy37UhA96J5FBNxB9M6ruQ0dBk14Wri3YDhd2BOvyO9SySSkjjCbEi
2T//a8D0ffbqhwYRJcGuFMYFYMrYGqgUuju1QgLV/mpT6REQqQhCiDpyFqlr21Xr
rnVecMMiCa5NRx6khHUrMV1ym47555lX8QhrRQAJnGZZKmCXs4b1aYMwbCVfdTn0
1K4Z+ZXx3MHuOdObUOLTVUa0vvOKC1NJhmVMDkNIsnA9VL5xco/Kb3aFW+Z5rgHC
isWAFeqXJHn+2VrxQJk4W0Fgtg00Qjh6+60pOSjZrIe4V5c6DQKlqJRL9jqL1qGT
5odY1iAEkbVsLtqjioPu2pro4p1FtQrbYnJFesybeqvWgqpjlgpPCujswVUl12BY
jJ4veqbGsZkEy9IKUS6IClus4ae7SdB8XhpWYAXwroG0sYnWrETtVnyQdnZJS1bV
etPEDGQ9zZrZqKV0dWmIcALeZkIu0yunUevoH84XEGak/6wsJatdW4jXICPoppFM
QUlaG6/49wCzhon3e+3xwpCqv3Bz/1jN+yaoQ6CIbRby0mfZ7Kgjr/s7em5EFCbe
zCFFpx6TddXRplfkcCxV6UXMXOZEcyUKxwOxzeUA1tk8TCt/5/iGn91+DeYD2/+u
tv9TchdrPhdVcduO5wJUyg==
`protect END_PROTECTED
