`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hgSFUGjATWiOtIxBD4HxGURbcsTr3pVbvvQzyv+5jul6ma54/gker53AdOuB/DkN
bazwneHr78kD3U7PHY9fDrnELvk6TYL1gUKtQIyhJZgWqGl+375M2aob8/aGDYv3
t+QnkmjM4rJZE7YVFENKzwUPJErM5G6v1aArA5J/p+IRLUV7waOZdcr9R8HcA8GM
K6NZvUJjeca92pdlk/a+JkHrdOpd7Hj+eHR/wbK3NBJnxsKVkxJ5x+dJFX8ums48
ScIWorlgQeiGAx2FRUqXImKsL5GYRMpTGSoh2NoclDptoznvQN1nusTIfkkcjBi0
mS8RuQ/DPXCezk+MPjJKd7rkr6g1ucoQimFmOVKwFe1yGgI/bqlquEHQ/VbLP7bV
V6TdI2M8kSDCem9YHqZ6Gv6cFPbgsU6VUxKHHS/jaRyTEKGaS9EdE4WpeHqN1mXl
FxuAXd4A5MlZzUyvf3nxqoEKdbcnp5gqM1mDGxq4Z7s=
`protect END_PROTECTED
