`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1kzqMfObYdSewWqMQAx+cShkzUzeVSo4fuJOULqi5Ix11ugqtXFdY4KiLFfpAGHr
W1RdW5JbFDBC+kgVA7D6LE8Vc4osiMsvpRkrbozkZIrFGZcMwczMlqz8xXA7VUDx
ksSofXTv/ygEoaPNR7ObfQWant263Yk2W6bWOJywJzN1YyctlLbhKj56o1IkiL+j
ckD4PWxA0jEV60tuWaOttjxMJWBIiwj5En/wm+nWed86quVKBbahcBjcyTidNQzj
ZqPoLhJ9N1nI8zYe4fyXh5EuOW1w1HBB9Dj0gzSpJmPvM+DWsNxR+rmBvZTsOFEI
aaRiQRI8xMjYwX9dUFVv2o84AkNuVieo+GJ72KSiOxziy0iK/OshFvUEdDb2o3yk
+9HE8voCtgoL+UwfMS3xhyUGcB693WnoUVxvpb4Aye1Sk3Fg8ls+220o9dX9ah9e
BXv37EL/+wesCRznaUbOv/VfjMdlobMvuNilBz+XuuIJVmM9OsX6d+vKvtYx2EV1
jRXAUqvcKNlzETocmycunc/TvtQwHPNkUG3EwwvB/gkIQG86DwzDQ2+yecKT9ATH
slKsFxdKsFR3NRIGSM5Utd0TINLvwnsHYSQXgGdHl/OuV2E6eu2sB4CH37mmoZT5
GQsibWaZRUbRsFlK2M4gzPkCWxux4N/YivFv23hWnLNbAigyUMDYF5AtpUhyQElD
tU7po4GtS5FpPsPblPvVzJxNmYYZ/kS5Mo6qRihyVY8ABykRzWBPLei7F9AA+EJH
n0i7v5o4p1RIjv2qLVDfziELbDJUcK3fH2L4c1+pTE3UfuGp0Q3Ev72HegYQnHj8
`protect END_PROTECTED
