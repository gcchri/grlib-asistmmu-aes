`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nm5BRbw4srVmLE3EOLCdH05aqipRazrU5GV9fxsX1RgTtTlsezdLhVSfJKZ7B1iC
OZEKmBXMZc/jttfOrJC4TuUaMueSc1xQ6oapADpk7gzd49yEQre8UbDRL5lwDfBw
KlPH9IcHrVTQKII7f2kYIXBhxLNPSVaOkwtDBm3PuDPHHL6fAAFawH5oqkM0DZFy
1/wBiDQctfR2gWzQVSJqCFwsxvld5+vyaAn67n0PZbgExadfTJDYpVMe6p77HPWm
+eynQzFJbmR+UsaaPBJLfqoLGsN6K0QpJFCKWKbEGda2+DiiSV46iWrPu7uU0re/
gzbHphtiXkUOZwHJQX/ZN5ueCdmEYsiLcHt6YOTHZzdYbdZAIkg8W6VnE75KkEoc
891k4rAaNrBF0Op5NhzgSyQ2qapdw63d46vAiFOst6kadUNlJs17YxsXrrlcZ29j
SKOjalcOwR7nL0FnoxLD+HvjyNyF0xkZuCETWqJntBhvp6GQGchwLzOWeHASRQPp
/DaF3kfyuPYtPJOknYmFLJrcopyFCt1n/yluFKmTQV/oiSjJkK9a+frPoCRW8gCG
LEzIibPTJLIanjyPVwVqcBs9z8JnObnq4TWdLwS91Kg/smY05oLXVPfV+ojsTxIa
pU3ydhRwkruIcuIAPRdJNN732ayy5PB2K0wsMBHaqiMU5cM+c55RK9A5uQbizdI/
TZ1bKmYWgJoZV3zYBCTu30en/vdCiTMED9H+oCrNpqWOjvIvml/g9pvRQbMXBdlC
8izKXxwRREtbMEbKN48Bytr2K9ltrFKdPSUL32smh/NsJ65bmoJGX9pJgiCq6yVy
WG2gbakNp0TXVd7CDhlfnWqpiwJ8M1q5qcKWlS9v0/gddzU8F7Yn54gthPj7j4NC
PfmWRupy21p9VUWup8kYBH+IemUT+Qm+YJyTNh1bR5byvViVc3ZyW0w3DLJjr6+g
kmwJWmAOQQz9geabp/LNQN0OgvG8nRaQR01SQvtFbGW3C6RLwRZ03/rZbu+Nbhtl
GvUDFurdoun9YFGmXBDrphfrNIMtTkxy1vV2nuMQ8YMYN94lY2iVdOSk7Dy73RIy
BW098rZYILOFu8aW0V1M/mjHJeuLZCnaFwIcakEz6wd7sImOC1nLbULtWe6HVK+t
JAmtPQ0x7R5Npz8Y+ffbtjqVyqnfQfjvPtMQfoq0JuDHM0McBuK2NezQuP/ux/AG
68Kwug8He3rEjEN+3n4wtIOR9YLQEYvFApxA9z54agbIJoG/lRDF7m3Dxugx6Ltc
mxDVwGyJCuH+adzsdpk67pzAuI1NiAfpJnzSanojqCZhhNBbEMwJeMTgkC7xwJPQ
xRqYTonuCxdOqTrMPNHAfo+kYae+YRZYoxFFS8mwidmg5qSY7Z9AScb0Bmz/wvJr
dfGXS7QN0yBgXR+wzjoE2sPfYx1W7qA5U6i4LQ5n18i7/Tnx/LAuRky+K7Q3FY3d
jbdSnW+tCL3EX8ngIxryJ0wjTHPfFdv3YXTko7EKOUQBbjUNmvYeHVsMDCOTWHeK
cRT5RYxm7L+XH56GHMCzz4TI+thyLNA6dwZ6KP0/TWZDSrM2PLRT8ZY0supmxh/P
kb9QsPw66fNG+qiehy0mwfX3PvsXE8/t250BWu1yadY3Rn/0yekdc/BIdb2bWiON
V5wi7QLSaqdGNJMm/mUN32LstgMkDgt0dBJ8gIUWGAGnqdHGjzACfPh1dCB8c02x
E9yL5OYR5k02R1UQI/T/WDHoEuOgCHlnCg3KvFBeGcW5FqZiPc7hrUehZxDbUO+Q
GWAsU0cE1Ws78fFBGzTfL2inRnoXBHzq9S8JJj8jLDhVjfn604e+OQlQsvtE6APk
d5h6pLYBAM2386Af1JziIhNjRq9zAMv3fKjRoUMXh+b2A0uoKuwntq5fHsUB0IhM
xtgcpAt76IDmMycZPG8p+TCGT2uX2ICbGW3sWZVJgUj0vZ1fVx8SOwlHk+qHf4sN
JQ2JaANAcSDpi8GNsX9732R/RXrrGfeiOu03+sKM674ra4u4n5k1lslLc4iff2Ca
U61J3HjKPCL+Dy8luLonaQ==
`protect END_PROTECTED
