`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c1e5o2hRPOkpOM0KO8t9kDcwkEVBH14Rwt5E3tauBQphWoIOvTjyOjJA5TgPZ0I7
W5YZW0E2DmMjfzBU6EzRad6eK/bcL4nczpV+AXnrZ9PoNUNI7Heu2GrRjqvnL2ND
mxPCpwx9itffDOP30AXGsaLP6Zk1m231OLE74iUaaKk+tBQfyMyrMa0QrnuqfIg9
n4wJwXNrr+SaF5XVsdbw77pvKHZ9bhS9NKHT4a2FIpPpS0dL34v3iLnQV8FV5CPP
/aImZPJEtFRpvy+GvER6qWYu2RfaJYS8kva7aCa+b8eVSZIDMHya/URg9+D4LUCK
HKcDZx83INLyIDmZ2e4IFC93Er7z+5NqLvt6MIadEhwU/xNWr+Lz1J6JB7rgFau4
L2SA4PyAXjPLzj19NRTp7KG4DVGc/i76uO94cZdC7Q9/ZYuHM/RRB/yJ4rT4b4En
o0uExe0lf7v3NfI/GahjuC82JuFkZcCQV8uD85MKMj0Rz39XbevA5eteMUVt+Hp4
1/XSrdAjiXCnKLKVVI7SsA==
`protect END_PROTECTED
