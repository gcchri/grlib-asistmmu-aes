`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OlkAZ35Jx9h2kQNEfNA88HT0VgplZ9fHq6ZfGy16X3sArASt4ob5T2zReyERBXuj
2n7+ELoW8PnenN4D0Sz4QUUebEpbeCVyCaAZ3Fp/j6a9XwN2iYpjoSnyRuDAfgJc
tTjn9aIkEBKPrb3og1Z5W5oRbJe7XOmFmGUzf+e+9oasAFeHy3R4vxJOYbDdVopE
+PeBUipD8djtSHqV6Yvrt2X9F3Q+FKjSeqPqInlijWXMa3Iu90J2ziGg7SU+NEiH
HJgF1ZwWb7U+kPWkkhjeA0nb+/XsdmyBiZkXctlq/sg802hn53ajhh74o12JAk+N
SYfNFaJipTD9Pziqjb1EMg==
`protect END_PROTECTED
