`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iPLnjHUSPGS0O039x6jIWTCGOQ1yiJuxADIy1heWXRUdnr+/waw994VqWf1YcR9w
+hD/ys47cnwHc1RgVs7ELY63P3o9RzoSrHi7ryJLPyaDcKpBvcsyMQeccKrC/GCF
vhmw6V2RBMFr+js4WJlIsRXnOqh7zAkYPJ/xnGqCsg0aAKsfK8GnDWWgHBVEOVO/
Iuz4mIj4kWAJeZ4lzZPVS95W9U8/YXtCf9+BsIMx6nSiIJCNE4Tr9P4boeYp/zwC
ixLL3XxWIguoF67cLOAk4LNW8usfpswBaOKqCds8tXl3r1Z5i3f39p/qd5f3rjkg
ysE/PcMX5esAVx41DqcBdlkn9vJZsyocS09ZHwuAPrMXhLKbSFMetcUtz8Q9lvTL
ikTocbBCw6t0zdByfA6naZPlz4Rj46lpWBfIZR69eSGbTWTRUmzuk1zSUM7FucO4
QTFwGV8oZtZZQclYBZvcY9XzDrnSYWN+8ExZDBccNCkDHHp+Kamn0xGB2cjI67Fw
gKy8DiJ+LyZkhBuZLd1X1nTRKnMZGxsVq2C5roUpi1mnxr1TdOlVp5/aziSMI2P1
zxILzdwmRJvQaawPEnrRKRxG3jzloMbhft8f6/Ld7a4=
`protect END_PROTECTED
