`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9EI4fritvMv9dNj9rUoGoxrs+Db6oJpiWg6hIrQcj7bf5bWPeuqfL7hxu5+vSnWE
GDfaJajFBzJKP21jRbCu1V16GCwomDzSqXY9UkGnqQI9RQQr36p5+Uks7hlxzQhW
KrJc4s0WEf277XGR/iriCtoSNMrooNGvVRVtJscr7X+LvVB4dswJ8JPC51VV8oC1
Agw+UOKS+6q4RCmBkRpDe8pqCeIggGIC1WMyy4ZtnfIr6EFDwupItminsi7VX1k0
7rfXs8dnEPNzI3Yj1NjyLCYJSR6TG1Z9oy9r5UaD8z6yj+5tDCPeze70OJ4qgKwg
TwJRemsoAHTbMkjPHHYvNzlYaQteTDv6lbHM/YDtG+KwtdtWOjxoFVF6b3+sIALF
gpEVI5vimrZOU64gLbljP/i7ctBhYWXJ9694gxJoO8X9nMLXc1zb2lzicefpZgM0
v8WDMMO7nshsyKNxs1vf53VXYewnyY5wTL4lEOMPI2DhXbGNyNWnfkCPqk4ufnvD
addW7w7JLTlnkpuMo2gVcl3kRvZeB6SLOuJ2Nkp77gzbWxsV74xC/sytWKeGxJcp
IOKKgwC59Cl3FTp/FRhp5Fmp5zqwDoRl1G+/Wq7tH7VkmXJ5n+I9O88c1dT8jV64
kS3qsND4am8ConZQk+MaZuy7HpCYsg71F0idPtSguxYW7rWcppmeg9LV0JAkhB+7
Jc9HyJm/14QAbfT0jRfaY1sdvOiRNMim7AsTP5XxOIS1enF0LUZNzGGb16/+kyGN
Z/nlA7MtnHTVV6GlJxATEKh6Occ/D3icmjTdKQedq+cNKOTWYLnJXjo/nDbNm/ff
5013FiZ320WR0B6bPXu3f/96ZFjx+fR9vVaYwEx6m1WOOjVOXRbarmM/LQFaB4bI
blj5L1/0Vyml5FM7FhrArHzaBJj+uTJvZXEYKbvFD6To+Wugrv62mBDK0w71wspl
30f5owzUnGD1KLewH/JbfNim3m6yFlzpB2IcLpEa1nTJirK6t+VEFc6k6WCLfCDY
h0qwLAICSGmgfODhf39RUKhrBtUau3VxmXG6UuGvAjR5PiSAjKRDFlIWFzCt4Mar
nW1ZRA6GVx1G2ma7CrIbvdOONlNTmK8wJg4WAODQ8N1+L6/5o5q24X+1qBlUk/jf
MyzTmyKTCHmx8esnOGOuGJZVfJbaFAfhkQnVAOzYo4+NdbBBzKxVY8GnRFRWwIbX
Y3t6F9R06XfGkC3SqjGPqTd016q1q+E5Sal7w72UUenAQfwUx9EmVFIqQnT2JfBb
qdHvQ1IOTnxOfXUgKZUn1YwnymGJ7WT0LuKM/D5nrClJiGl2E82faTlmmWKBYloe
XC9M6ZFbwpbXt3J/t+LvLMaDq+0Hp4m05ov8Sgr+YJH0a5hO0mGGwYkfHPqjikRG
bUdsF96juHvtAcmwluSnGbFXQtzR92gsaRzWAmcsgHdol8TeWh5kpkcCz17aPHBz
oQLVFdVqOzgg/uJJs0GwQa7VK5PXNyzyLdHVIgJxmb25/ZDsAxLAZ+hFQlRM6j3w
pmeseftZofUakhF+wdGyMTxtLJpHBhe7bGeqq+rsEQKnd9JjbkZoX2AF3giC5lL6
5gozpK0zMYq8ipUWsNGYZ4M+PTplfEtdVlOuUHJCW3EI3sFBzEd37RKfqnS1HvRT
VWbyo8knQ6Fy8ptMZ7q1JpRM/ShYgGqlMEE0Se8aJEOkemsqxUHc5og30cQQ3EOP
YiiAS5TkVKz1PvWjOlnnjOmzGj8DNvrGU4YInx5V8Ash9MGhtaHDM2W0T7gMsVjB
Zw8BuKlbf/V+J9+tzMKb0LOrN3rKizMirz+j1lSq+dZ5i+h6iwsPvv9SN6AMxUZw
nTkZ8DDGjiJfAWowiELJOOqVxgFUPVRH/B/8OZPrjf9iugZsqP8hhKNo348PM08w
Lr1Vi8rvG2rlLvyIwhabig==
`protect END_PROTECTED
