`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xi6YhD7HKK8EUAOfM9E2lFjL/PZTvuKzLspTkl7odyYc0kLcRkqYQQ6zD0186fr7
8ewE+UJGogUx+OpudVMEWGcilEUTc1r12hQ6C8OMrK1Xb3sm04tvzyVRvUhQIaeS
WIGXikhDT9TAqar5DDZHsvN6lRhoNJbIs9ILTdYI0GqMpAmlFNlj/imCvyz1ZYr5
vQNIABEc2dj0vIe0WRHplp/FaGdlDpXOtT8GmxT7zaYhibOWFn8vQ0c0eFdvRQ35
LWmDumpOBEIHLAJdItOFx4ZDrFrnnXZXfXnx04xuw8wujPQxcKbdkhdY0twgPKq5
CunBBgXKQVFQ8LezeOBhuAVLOuf+VK41JNNeEWb+oHPR7cxz4E6pc19MJgDzMu19
KCs02CYDCwvM7HvOBF89TgdoYRhsAZW4NfQX8+PGDQ4bqFG6f/ZaLqXyZJ1E73WE
xXW2ODCkjRwEyEW1Ha3ckJknT3v8wNZ6IyVL0QOq/yzHi0hftIwJRWhXYbKYoEMe
VqzNsMB4FAUTlkXUETEgnP8QX+23LZ/CNtBxGseHTrynoPqdeMHeb0nQEk27ptC0
`protect END_PROTECTED
