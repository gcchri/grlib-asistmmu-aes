`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PYz9PdIZJwjB3dw2Alz+RkJ1LUJe7HtGaIVTBdju2mJk8a2YsGPoUdudWoJJGOyx
v9Ctgj4WRllpAqfll3v76ZeGPq0HraQSp/2HuFxjl3dOqdsCDHup1GT2LTGcxmb+
NU0bIEN7VLNgWTJIhAH/Q0ovomWirTkyZx1d2bnwvbqEMTfAvVOKfEuJScwqlmb7
629j0mDKKpXDz7VFcVOXEviEvGmoVulvldOE7i3R9eQY/bornpUN9CnpMHIBfiZI
OGJM7ReEV1QOKmwNQfHLJ7fcRD6EVcDn9/ssqHX/9YHla4bXYcEwDAGyblQZXo6r
S90oSdgFiYnuUNybyJXQWuMN9JJUKPPbD4YrVfsY/YK81g4S4vsOpL/8CtTsmTXq
un6Vp6VO9pBks5ZR2rbTy8ayNdHM8WuLLYjhvMsSwEzrBgu1Z/NBDs3omKEfi60W
MFhsQ5Qxr9DE/S2x7QaRHdY4t4j43b6qM/t8f/AoGuRQTQe24d4Ff/X3RscZmpyP
WSF3V3iadr8rVN084+DeG+VGs9GAYPx5tHFvex2dIQV2Axb2d8IkofO1N4q63yMV
G3tNL6wsZ9Bn5/Kvq96ySxCE5Fe1B6taZLbinrKEOo9yewdXuIeGMvnL07A2G3O1
O9h1hMNoOY5WoWkU2ggOuD5LkI84jsm5Uwsfe7UeSAxTwy3q/tEY+PC0Zp41CXec
xr6HGmG1vZ9E9600bjSkoB2+QmddIbZPQ+IAJv/DDfPYA71pYDg8dc3SkDLL+tBw
kUqjFWqy1/WVrWg9FYCGnVr/Z6BscRNencMP/4cbBoP9VhPakREIRPVmcx7cCeqr
1kI3GWx9vtJiplS1ZspSCGZl9/7XKS4kU5AJSYV0uKJ2q5VuRiZiKcaOC+M1TDVp
bfT4PrVSHrvDFLRV0ljOMpbPmo0MVGopOurwsl1PREfe5kCbQnU0lsC0muj7f7xf
GdMCJj4HKf/XoXCCjX6SxwOJihaIp+t9FiseW4r/RgE=
`protect END_PROTECTED
