`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3J4aoU7hrOh2Nhi/+05cssl+eVSehOo4AjzwNGAS6htoUKBWeZPYh4PltV4ZCHiz
jHaXb3zAblxd7TGjHOnxbbeJJhVbkSQCuBSGbQi9GM14fnBBjdFnNyOTfKaoqEcJ
JWT0l3UUz7EfSyWTeJvNE6OYkJ6LP1HfqrP/J1ZqYp/tNZcM4KGPnS2/Nq3TUCtr
JtgdMM4UbEUK23zDXtnJ+x2Ds2KZVlW62gh1zMzqNRT6TkUuWYb1UIPES6Zur26g
R15UfUZpxQIU8jn+ziWQDiDE+sp+2goYin9aV1Pbd3OXv7aV7TeXkDZf5hlCkU7j
ni6V6JsEWGOQV2eTStgKrdBhHsEOuS7aPDoY2ElS6jGQFqcqw3Rh7TlvKZkLGXyV
U7+IhCzXEyk8Pf52x4ipDVA01uYBuzsz3x5f8YIXUiBAqg4evw6u1wrtK1xmD+Wa
rjQoIQ+ZeEGcjbtcrlCdoEuwlY7LCANY+Y0bT7E3KQzj5pp7V6HaecxjBmIia5Zx
jNhFosN8hqFOVBBa9XXkhs67ArAKlbfMIwtAiETCz1i5vkUCNldUKyis147ddlIR
Zg7VU7+iVGkzewU4hV9V3ug6nd5NZsoxTy619DtYaqFR+rc2mwtGrH9E7DtRH8Vc
mZ5BC6BXh8W/139yOb3ItS6w6zU0FW+ibb1rxz70n/fb0V9/im1hLoobeUgbVkte
7CizcjoaTfVaKhb2QuMf5CfyjlfRnqYnJFF02liOuRUsIQ35mdFQ3N2Qlk1ZCdIi
3Y1H1gNARY160VoAdse9NJQxgfUeNw3OtjD3kl+p8TXiulQtsJYbIF47fnMlp7NT
56DIwSaaselgvweJ6CS+2hd/h3YNHnRxSSYvOdSNbnnnbiw/xihYGCEhf7xxM96q
JynHTC/Gz5sFSmr21pWl6NL/LA5ApqwJOcCBZW/MXXHU9UQ70igJ2fFG8EgtHCQH
IBeyDG2enOk9CgNlE86Bh3f6eY2U3zBn/S54/I/NKvoSHhpFYEwWoroqEO7duuzX
bZsLhrdhl715cFlERtdol0PRnh0HS+pM1jmC9og1gc3tby0Y/bQv54uAEasBLuO8
w44hUmqqXH9va8lcW4lDedy7fAbmBjWa1jK+XVZUDcupB+LHDS/DlxU3QWU8Db36
QTsrksZlXWuAFPCvX7Xu/Bs+yuB3leEjbJVhpaUo8geXobLSeDigcPPLjbYyaE4O
LOAyjdhQqTaMST2uBwwr2oBK6TZIuvB1mxNxS6WOrDZ+3U+NXhWYvGYdB7mPXAKz
IkOvUqGEXO+dOcW1r8E1aLZvMpXBae6JaUJd7I4oEps/fjDlAC6JtNUsFGEaxT7d
awevBpyEpluwIvPq4JguNE2KKcRwtMViZtAHeZGXd2dpq4cQPm6DflS/irSx7njx
Q70RvKAwiqdJ1fH4IAE69hd8a9KIYbqOX1JueEeXfHLEcCFUJnNvnA75UIpYE6SS
sf6VAwXWJKt0+RNHXfnRuDSbBY/BTgESX6rQL7eWUg+yuhUdHlBSHrd+pPg89M+k
3kFZhe3kpRVlG1+DSNtpgJ3kUxXRs2LfYiQuVu4o4R2BhO422V4ueymAyJgU60Ae
ZZ08a85JlCZB/XLXI1tNqDm7piYim+JFyTpt/JTXwlArIPDxhTBDTp6KxFS9bSmk
+rLT0sX4lJ0JcDgpoPNX9XoBVCasoAGZdC/U1E8uFyknDOBVhlA5vGNpcs886fhL
9FIrctqdcuM15Fv/nasjQbOK0fuefjgOATAUbGhxqSYYZgDd9D58OWFyQxihWDet
BFOC6M9ml6r4Zvo2EMvx5EIpkZOuwwqU/M318BiMk+5EBkG9Xdm2Sm2Je3xOz7ga
4mJb7lNEBoVkGd7KAQUA9gAhd56NwqPiSavdNor/R8pRGqy+ZJ/MjNK44hf9uug5
EB8/HW3xqmTebcdobXwh1nobAPZ9Xl1wZwutLkRwcnbTnkwbMOJ7Vi8mIOdRIuQK
JWszl5GLMKXSk3tMqLJV1Vm/pUFMKQUBR7LYFIZlnSs=
`protect END_PROTECTED
