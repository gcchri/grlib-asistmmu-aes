`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TNS/D2vrvHOgNp4qiyaErKaxoFJFMiznSR00l/8IaCp6XKJ4x5qHueTEDLG4z6P3
mTn5p5mrZ/igUYt/PCmND6UXcp6Td3UYkktaqDbKahvwQyGpTK92FELaaQDYLnd9
j1hlspjIqXEccmIHGT4agYr3X5opJk8GpnRNMfIEvM2CfYvRiG3mEDDjoiJw4RnT
ZOE6DEt+wS9DwJQeqv22OkgOAI63Ew989fGKp0TQWOMTrHoskoX3CgzbIWDuPmsM
Pb5T+65Sv1PKgOExl8DYrqwoTuxTne3zaLKlr8fkmGIxcorxgVkuDkVbzhdhbTl4
qRT+kxl/geUTLsx8DP1Gxy7gFjx64fz/2hrHAgfK5FI=
`protect END_PROTECTED
