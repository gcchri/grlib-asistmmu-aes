`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pHYeX3CN+3BpTkCCPESYIW3ZMwXUm6Z+3CYb5/oMaNa/PoR9tmuvXF7sBDWr+9bK
B2sVSWURgkyyko+P6dU+G0dlCbd7oNAW4pzQBSo6IDGEPSwn3M7P8dIwce39vK89
kvyJS0BQMUKqVwoJmcwJE1sXLHVUvDhSO8Ctm5mr6Px1v3RbWfQ14knsIS87v/yG
AaJtYyupvC3KhfC7Jrhc2iIlLf3e1m6jp/qd4bOcnyALpWRAS3jJk2L749r3szus
rSYI+NpPuWJB0TEBGObbP5iA56Gj01uL4wRXLGBkVd9xi1enLxEuUIK0AWrEgszH
l41jBvg+iP6punHvX6rP3d2z1NrsBvjSnq3OfJk7Dz5MC/7aYQ2H+ZhFup3m4eDo
vSlS6HnTKT8Q5n+upp3wzWlbMOmeVVgz4oWCtJTbBiLdhLGc56Z/yL8aemlgHp4O
lEhr1a+AhLg4tgQkc6dEGactvVkbvc3yYevFsUEo+CRhIPG9CYPRYJ9Uxawr+8ow
SF3Xw9TuFTpqeUImTwhRK9WrKOVDcIsJyKuMViheCEkiyDoqZdVLUh4TvqmpeEN1
`protect END_PROTECTED
