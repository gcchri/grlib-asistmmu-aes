`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9DF0MHm0DD8Ty4ZlxpqhE8fzt0zWWQ+IaOoN0vjbxW214NUqQa6kx+1mPCKNQmRv
aUj3QoVYCX3YGUcmsotdTc9h3Az+9IoPVLN27Yx9oNuiMqhGgAhCeycTxVujG+iu
ntyYM8IZ7Lxm2ewmArmeVinZj8ucIhSmMwhCiOktLCV5kApoMSBGo5tJQnTWt8Xg
gCYSVd0ujsfr88lKObcbB5/nD2LbU5BcjLn/q4Rh/d/sgbIy6OYX7gE9rAVGQK8W
Ju0t/0r1f5fPYm3yp0y6FYzGGwCCZsPAOO4BXhGOoQ8YE0/zqAU7FLspjBvYdEAQ
Y6EWLwq/K82MbN0Oqpe10JjnD268wmrBlBnXZgWZ8F5dBd96HWXTkTqbJ/Srha3h
IbA6wnooVxiKxn8ep4erOoTFgCSQNJqiyjtltuPY2BGqYE6DeAZeBUUIvz9X27DF
`protect END_PROTECTED
