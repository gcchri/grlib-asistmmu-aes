`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dGM4ZAvjBFA9DvyJCeVaCTS77QzEIbSmkqWVBR3Va5P9f+E3FJuoHsu/lycBampB
r0glYTFW/o6k/x5QNI5/ju5gRQ9KbGZE52GASULIoXedr8w9FyGsKY0VZMG5NviK
5erdZ3wOi1f7TZIxxJgTuD8+pW+ZXMRrkJS2PYpY2WIewH6ahOOX6t69d3JkNF17
eR+v7K1efzo0SWnFv+qUEq/wBcnhV/yEtzNaeSVLqUk9nrpI5wlNZmUq34eYCDx4
XcvNORGZQ9OgqUmlb7/G2g==
`protect END_PROTECTED
