`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JCaqfFY5te62uTjBvaI4+6vYhYt9YHEbkzh8zB5OgpMdxqXHDdPKZKid4gB1Ccuk
xosNm2sQbVEx8vYZK0qUnLM9A0S/9ParJuXIJdXOtZOAlH8EfCkHvDRDnEKqIp9O
lPN1EANzAU+BwuZaLndcbSnR5DS2KdouWX4d+A3DsUxaahFoJ8GIGBtxr+qJ4tKf
eWjSa2dCLnQS3h2wOj6OEDOJkQd4hyjpot3lYJJGhq0qPHFztA+Lw0e8/wx24ovk
iaHBopfsZ6WGfT3m6dZ1yhIokb2O6Ap5nTH9Ziu5Wm6wtkClBfCy5FwqkHUwgmSy
jBbyIszuMdPaqkNFF0nNvYm2rYoLhllmD12AHevcZ85gegKmvWTSK6vH/2bq5NOw
kAYWrG2iPK4AeLk8iIzHBhdc6IrQOtQcyL3v+ckJACpLlHi7Sin8FjoYixzuLHQN
oKDOA8+luDacONd26AqRDcA5lVLkU7D+wmzi7guGB6+LDNKXk5qKklRDzCki2/Xb
`protect END_PROTECTED
