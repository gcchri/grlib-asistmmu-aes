`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h0wnx0KZnG7HB4uLap12Xa1EqAwdCtYfJRXxTJ5JV5v0AEsk+HZO/qPSHXOiioOB
zSZgNUSJpWVAhUCegRlCixqNXqCFLazxRSiITzohugnUNBXaXZx6XcojzgMVf+Yd
QpVn6fTX3LLS7hG3GKqDLS7lACAEMGb5NoYyL6I0jV1JhcSkHE3JdThgvbD70j9s
GomnltMaXWXDnJt1kIVjLei8+dWSuzYHWYh13OkpdpW5rfd+TueBYhgUFPfKm1LZ
yq9RgE8V2Llkxr/pKH8pTwPjqjuZsU6r5G1zQD++HsrfIrkuJXmSunofLtiJottd
7YSl5a18lxLyKodNAIMVgddYXIucHICbXFR+ygie0sYy6rB+O1beXTKxvF39Jglm
ueO1qyVuz53++VOTVxsdKW+7sA+IoXO68LVUUqot3KF37MWwQkB70eKciu0wxNAN
fA8mnPpzV1PWE/LreLL6x5PB1sTxrJuHeRWEPrJa98NXmufvNjeXmPJG65W9lMFt
DrL8Uws3HlyW6zDovOsJ0UiZGOvnoW/U72KbB/m2LWhohme2GCk2BaEOlQ55IMdY
wNhAU2f5nD4KS/klNdAYlaJI6Wkv5U79/xbrfzMW6c6PuTQAFmmlmwk0+b2xrvQz
zBkRP2d5jiJA8g7Ge6MB4ODirIJ8K5ZVHxqakg6J5H8iy/5xRhKKU6ID02vOrqLx
1bjjCTseZxBvZfKkhkAn+0jTw71Nb/SRl95T1PGaGXWpzNnbdHNP/8d3wWHny7LZ
RKyuR0w1/fMkUj5f8MLE2LnC9k6YC/J2gA2oE/vwG476sg9JNZX/YaDv+2w8gLr6
UgT+vHPADZStKm9VTgNuek6HgM/yBAYge0QwXAJOrwQDgUf1SFUxv3q2GWUCo49n
2nj3/8NrrbOlaTJiYcsEyzvwjv2jDCLsJMSqDsUYGZ4q2nC37r6BCCueEUlsRnW8
MRqFt0Bx1Dmghn7YEM0+NVymL70PHQO3AF6XoyHq4P1sx6JahDV+16RVMms1G92P
F5VC6CjG3lxoUbMzRP05iKA6cFZ2bl7mcDk/Oh/ClAvhGrdBsH/Tv0E5Hx7wVXV1
vQrys3C4l13KzoH/KU0hyw==
`protect END_PROTECTED
