`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uMsRsbp6LxiSMfzL2X1jKnhWC9FlxhnOZXyXGOlGoXNpVIWqx9gJoHQrxZvtwHBK
sp/p7TVdgMk8HZHpo8lLrBPyLKli/+eWEKTEnklxEhbB5jxAvTMhois9VtjPMc0I
5gq7RPF+NOBf4bl8nHGwth9nLxxnTl1FxD/d9gqMe8c7jud82T9G4JV84vGi9/JY
sp0p77ieilI5YbYAW/fRF4foyMocOnv8fZdTp5Y67uzVpFLlClk0bDub11d3FONq
+GLSw8XRq0TkOn/99zWK67I2tcaCLg4AHWtVQVVej6jJm1STMnGQNDVjdFQxRwS4
UUwNarkxZG7Ey92ZUQjxHU0PIkbArMJTGDNME1KgzLSo8Ony+NTUEiU4rC8XirnY
SQbtNhVxcIAGFTvVZpsmMA6Hm1SsxlF/pkMmTEeRpp7nObwV7Ny3pwg1n+SpDnQK
LN0780SYOiglOhUrRHEN/ISPs8IjjYFlcZH2dWiItJUfiK0SA+xD99KlIrGOIKiA
aPgRf5b5gwAMB4EEwtcoxlJ7HIWCEESDwCQfbuuVKVM=
`protect END_PROTECTED
