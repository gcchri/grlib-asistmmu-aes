`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ClDaCmVrhqla4/tain3QSwOri9RhLrALUS+tmD8lK8jGvxpEHmxRdSt34HBqsX6
Ls/i2Bn0ctrCbLWhfqghV3pvDeMVvvX403peNyYnTf5ZFFzy3gsoh7yo1vgHVQ+i
fUVI7atAGP0FwiWHfQcjCzRve1caEOqszlg0xiTtnmT8AFUhx6wbhDDUdkcTfwBQ
5dBc66BGstc/sCAlnY1mKOcXuxU7a2jMl6Xuuo9CLe/N+lduiOVsfBVvrwCoEBJZ
axk8AkZuCnIGnCgwPnsBV+ObXj6Bzup1Uot34LAuszLr553ZlH/xYzCxTmPzGt9c
tDOJ1d7/x2aHbPZ32KUR+1rJ8l7B2WRpCd3Qz0uGR8/4XNd8P3XBOgvEm3i3RpFQ
h6/6QjkS72qbWTOg3XuNQneP5lXIdL+qaR7gmggi2A+tT6oyS+E+i19KiBZMj1bX
agH2IWQqmZHiRzPleLN28BKBXQn1URfksSEcwzONLcXTf4FmKOeNrtdPUDcUUglL
EZgu6Dx81SO++7MHVMt8wJnPipFbFIXcg3uJeMxJKI/l4D3TK/eNu7rsuHr4xK9U
xcqIcdjunnyvaqNxWNpdxvcE4uBDgsLShBz/0zutF/ar+pFhYw6K9DUn2ZJW1upB
GNSWz9hiwkWgLSVhPzOq2VB5PRRdSTCAKjAih3iQF69qognlhnH2H7+Q+axZd+p7
zidh+VVoppr2+JkdccwK5R1lxpkkSlGCxxCfs4xz1X/8CDLiEvlZM/vepYVisAlw
jjwnoQu18RwmXV5q8DSUEKFMu6GAKqsOFyzBhxviUNClNb0DLXPrbo5ChsdzSXT4
V2vhBkSvG7qW9x3QgrzXgYd0PAKK0LaJJBzUhIw1nkJaNhGHRWUSVzWzuFEzfnli
`protect END_PROTECTED
