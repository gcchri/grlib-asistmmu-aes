`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+QTPAAcjuL61x8NfCF/ywx4Cd7CYn36gp6BcfbyjGfH6Z6ZNPXMNT+2g5537zT2V
ZjEdOl+Ivb3lrlE/EI7oWyUq5Pg6KHKf+LPF5fCa9vjkjy9fVaQsKPEIh9h5ed3i
cpNsV4QfvC18ayaRcKuEVz/XeYz0HSMjrH+Jre6+iYrdiyRrurS3UWsntUnuiY2m
sJj+3k10FdMlM/62PxxDY8yhVkWb46uYEc3HCaxO8Aur6/MAk5xSx2nIK2jhgQIG
zwdI0H3HeMo3nFIBD8UdhnN5bdiz6bcTiL7qiAs3IoLJIvr+GhfxCM07mz8OfoPf
UqYDIIhJHjvhjO6/5HUH59TR0TsW7w4XHYJjvdgwTZ+y6yehTJ78kJo7tVVz84Mw
jwp6X3eFi0Ma7lgrIkIaxzZkNIbHw9XAr8Lq903NO319nmiNJbQvvWtQ0AdWrghO
vkZIaPLpHYIks3Mlm6iVpI3evQZXqI3TvIzCFjj9TyparumvZAl3yAZ2U8XWa+Ai
s3Gp4svVHqXHFbBe7PcDcC7Pnz+f+GE2hPXaHjhdjdCwdWlQjkKOcAHvljdESQ4B
6V76Fjzp2GFOCrWFNsyCOf69uEj0mJgsLFX5uA3azJpij5F870GqbPfjp9kkemY/
4sxAMaIYkG7+oKYpu1EMEjm27YDS3HQPqLjldH2gVFTpV+a0kxZ71Wg9BY5/YWhL
wzgDKhlPHAY/7p7ku40hjlVQRmaZeBZcuFHlKy3Xml9bpfF0b1paOb5zgKfxoSEN
enR5i1+1r0kRmzvUVMB+0tV1pQEOerxkD+b/8E8JJkmtSOJVKcWwFxhAz8Z8EQSS
7jHE2q6DseumLnyGNKoBTw==
`protect END_PROTECTED
