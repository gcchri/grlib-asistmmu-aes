`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rRnuxVGBjjaIeRVu3GdwU6wFLpcairLWNslivnK3iR6uusSxt7Dq5hrV0l8HwjQa
Rf6B8oTpMHIsNgPrLC5hXWKrBdJhXl9tXFZSEtmBRhSNYGHHMI89lsH+hcFizDOc
9l+w30QA2v5YCQT+OeNvt8WmEB0/8digdGM9VqbVLCOSQ+fS2XvYWU6VRmYAe0wt
v1bMAN9eeIVDqwnVVKO7SLdV47LNIP6WebUbEX7kD+sZMFIgk/z9LVpf6XbvSrES
hkwU+bguy7UoI/kRx1Im9uk+IMcqVoTsOpwbAlY6LaG23cEQLxxp3nuC77WQlQwD
zW3qR1yEMd2CeqPEaUZtLrpmY2s9Ox/cqyrrDD7zb47s36UXwGmSiKdwlEQJelmv
BNgfNjevZQFpn8JaobQk515n/6V+res2SFBa+LPZTdyswrfG3pCVvXJj6gg27fkz
JLme/cjOGUUJ0D1x6baAdmWUCDprlP+E9C1F3jqEWF/LPm5zS4iKKS5dR/zjXs8X
M6zEt/XFMqfYIXNp6qNXnkGwc3AAKr3g3s272HlQpVzCpuG/rBmYV9bjrS9/lgxx
x3YQqaCDxKsa9P3Q5OK+zleHPkJ+EY6oauTygW8WBbqnCst9l51jQfkyaLZbiCbG
K+GdGRqlNLJLrolvN4TAXFLhd8hsXopDkWRA0N9SfiajF1ClBaMyJ7IScFQoMsXE
JjPqUXvLQyGTYT3zLZePGXHJpA5rypO4gSdasR6rvuUT4ffLxN/UeLQvPqtd8Xsr
u/E9/zvs9DVFNwm5h9Pznv3mZ7LRVCChGQYb7kE2KwFHptGnX4EsFajL76WuvxAx
TZ2TzGm07hfU7jOrt5o62ahLNNuMhuiWQjrsYl8mIKF3LD16gU9Ak67HxzqGWv0y
/qxZ6HlZycS/1cHBxEbVPFpqXtZsJZy3pr7O3szlGAbvYjeTunnokDRYPR5HcgE3
ob45hWLTUGBob34HwUquJevpJLry+AfLLnLrguLBAifEshTYQ63i3JDNbhM9TtX8
JuPcfcdN7zPppLUGxwi5GtZ4p9KNC/oYUayBmgelmE5Diuuy24UjZkh+WTyJxITj
89h/olMIj++OE4JLeoxHFmGddXwpOLCvH6Cc9458Yupp54BtIK395G03g2kI669f
ag7OXb8Aw7RAiI6THmOnVpwnnoWMFKuFFpNQegpIbk0qZRSEWetQtXnF2NY60vui
6rOn/iLqFtqOYmqpUok/Hmk+yoGsOOfN5EA2Gxbl7CXiyzcx3s8AEeAn/+tNH798
pZvgJOAFf8vpUqxM7ez+mgUuBOFy4C62y2V7Ot3vjSZplo7ufbS+Rmb1HI4bjQGf
nc9VtEKQmkvSfbLtrCuUrslBozrhVnSTyuzFPoZebYHZHoN+8Q1Ky/xU4krlvASy
j0kSF5NPqr17M7DP83JiVtkVf517kPFQKNEC3kNQRaX8+xeUi+szA2lg98urqFB8
J73VGZ2xsHpf54DvZxxtSVfJkfQJl91/qJvsgPZTSIn3GEnLsYQ+bWoWzAX0eZDg
bGiFXA3jO+97oWII9Mn182g6EDydy5McfqtOKKm/8ymVLr9OJM0VaR96P1qHOIbh
LQU1abTblHpc4D0GGn3Nduu6uVnHzRzJecCi2QFhrhBnTjJLWChCjqzXoBKRMyTb
MslpkiSg3Uwk8Jxhst1FmIE+GWHhI28eGtAAjruhplDYokcemE2neJRP9VutcEwW
of8Ya3rGvBJ4ZznJzCNrf24/0jHcj6Ex1zn0ga90KQy6ECBVuakWWexb4hGNr3qu
KWL66KfcfdUXbw7pY4dlbiXBI4Z3MhUgILTmIZDqP4yKjXv2E1r9ADLtSBmtYy36
08ghvStCO2DQ2QZ5dIIeKbbeupb9GqBKhyMDI498PGQ2BPpTEquEYT6aZVre+qYm
nY6sSS6HkJFZxtZfiPx2HNtxOg4+tn5Hh1bhrTCpFMsO3RAmeOS0GI6w6H9u5Wgd
4wRFrUQDknqIh0/JJGVj3L9Nb+ZHFGEJmPLDh7LIa1c6TdnmUtrOHu+Vbp3V6z0h
AueCCwPjLI95qhNDcF5/YKgDhv1stsDp50hpQ9LMF/MJU6irSAWefJAZ+0fK/SDD
qfeGFHFRaJizqWwrzgiOBRdiF5IMzlnOD7t3XbMVh5ITKWeZ5z6XKKKi1WKGKiMv
HlYz3SrdHVamnOeBgReqRyb5w6XPYqHJzhFbkzpHT5M0xV4tJQZjnbeKc/ZT4ko7
Sn4krGRWeqntkMpzwBbCxbnBbE6eZ0COM2dxm5MMKG6+VOANlNz1pbHddqM4F/iZ
GZyvnWBukTKvVGjYgvGWlgDlRI/12PHuIINEoe08pfDvW/Id3xNf5ek6BPZ4BO3H
Mnp72gEF8Ub2ZQjQFwX4YdJ2N2BLxlRCIW3LoC/5NrUgpouoe+DNwzUuLNdS4Ioa
iabnzdW4vA0v6pUvkTBNlB5YFrGJf2PeBNXq3eOyNp7plv8hu/Zs90QUKhiPHV15
PNf6HHG6YncxQmOygmpNfcCmha89WDu79v3x/0qewRvQhUkzl3ne5hSvKMCTVn1+
PUKLS8ALH2q+Tyz/MdzKMFvY+Z3EsV7YPjoLYh/jmvskRH1cyB77R0yp31m3vJ6+
d90E7v8M8klmEodvTln+k+fj84R9rB+5qKjcNU97H3dEuomKqBiW55UVJUf43k5b
FZkEVdgZwsHMJmaVQV5767McF7TCccdyP9t/wMcQ4Zs=
`protect END_PROTECTED
