`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oa4niCs3XLs5W6GEbz9kcFurWgA3DF3sDgCMRbzThzgk8ZUbOAFrjsHJJwjKnwgz
kPjVtqhoRLnyvH574FBLuCq7w/xouXNtV2Nv1Ave5iGodTxVYWDF9calxJpbLliD
yZEOwlrFqSTskwNl5oW4iQ1arNSunDue6t8S3fUnwSCAA83YD8n0/OmtG65qJ6KE
nc8ervUe/MTxX7+t3jKJySXao9pVFhAo0JmbpJjNYABW6XkmWdBfuV6w2n0WH1t5
2BBwJ+ybF3nHLALjqKZdTRFBQBo+vFwfYVvCQtKsvmJdUfES8o0EFN/PCv1hlO4N
zRQTDs69gDf4aBBUYJXedcpKD0OwOezz04PPxI9WQbvHZANi2x1s58cir+7oe5ly
V97Dsgn1Y+v+C0QYOJWIXQ==
`protect END_PROTECTED
