`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UWR+WJgykKjYDYEJcbc4tmLAG4K+2ZIkDmgaarfmHn8+3+6zW3RurDzdQ7A6UsgF
8lTkOSYWLxY3nA3MITcqEWhi2D8bgDbVIPKqtlNiSMJEdXTewg3XbpnssHHneJCn
5xyj+5jtMf+JJtrbdu/djFshPURjVALZGKng5GewacWypP497Gmh067bcjbM8qT1
vFoKUOg7YKqmSSQSVouxSsZjNLYQcHBZ1rOrDTzESgvu/brxNT2PpeiomCKyXNG4
m6d3AQgSgegAyWGtsULuKnGGc0jFXKMVfO3HabWZoDSVJnUGII3ePT6iD9onp8xX
kwjJ/mrljYiDzQAKQR6otQ==
`protect END_PROTECTED
