`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
foPh50tQM6JFIYK7ZJAh5HFW1Z3gyw6ssIMU0i85twQ+rSoFde3E4czVqEfhuHnh
WEIwXGOpskL1W+sOIbQ+N+vdCVtsA4e8VoiNmrpTKEfwEneYH/EUaSySxM3F3hHX
e9dg2po495FBFE/1zqzTLNDNvJn5L+OHL6ts041mti558lpZccMlFm4AsOc8OmXM
tf17/d0Jep8zLyRBpzPLCr9majd2Fgt55+3MoKdRmv2A3Bk8RYo1mfSX0GZ/O/FO
cbJWt36NRoSBx0AboN31pNqaGBZzEXwWLbVP5gI4C79m1oVEssYSR1jtEe3bmWzK
zC91u/dAAb8feK6qs52ky+yL732fderpuUbydu3AFbYddp0z7hLrD8n+XMxGNpL0
edptdvnPA616vUJWGETxf4d6/eIR/F+B0BzCst347O7hX5YerAaLqOl5u4zXi7Ws
DN58gNH86cpFNiwj200ITw==
`protect END_PROTECTED
