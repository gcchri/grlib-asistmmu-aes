`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BySKsRtvvCE1wkBtX5uCVNmp2YYY0Ioi9PYR3c0TBZVg7s6FyttQos78EqaAlVmk
UoL5Rw/0MoVqmLAEo+B3wG++fo8GOO580CLdV+Y/w7px/tZLT7kRJZhDptkTogl5
n3sItfNuXXAfKIxvwREtLt87w8TgLBTXv2jbjy4WPclWGbDA2c43kQs3Sbu7uMFl
mLGwYe4pXkAN/8sMi4eJAIkzZP2dhkNWbV3Cn3vtTvYDHlSzlXH+i2xgv8vlfWCg
o1Q+svCzhstbYunZMAluDHw1MLyxOzx/kwCQ2QjeFoP0GDlFe2JuJbBYFqmCg7Y8
THeRb9UzBh6kYn3mCHY75CaFmMpAc1mfPGBlCSksbPZ0F7ldrmJNn6uVVxW7ToTt
B/zO1P6bOnPuPDg8wnAhsQ==
`protect END_PROTECTED
