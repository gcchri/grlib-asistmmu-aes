`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
se9iyj+MvvdBowpLexrqAbaAj+ZM15vaOzZWrnvmZ+wCdqeGwtXIPmhH7ozI4QCM
YaymRZ73ZfJC5gQuGRZEl6raAV137EkkrrkXrD72kP1AJOGTeCRGqzpvrbfn0yX9
LJWrvUqt3QG/7EiBskSDTfagfV1EldRJK8QYWEoJjc6mdAtegjzpzu3y+s2RgeSA
wekqJwfrN+85efYoCD0jNNBfAdAk0Ia7I9LrMzOkNWsXKrXTCEZoJHC12lszjlpW
FltZJwLVFw1zPKIvagUYsSJCJa0Oy6heyYCwvWxQt9Giplzm1DFSCZm9aaVNhXR7
xlnHcxqeC9TEyXU+8gXL1oswvziklQdif2vYJWrYkjJVgOmClMonSuxIU/J+VcJE
TIRu5xf8wT3zHBG1Qm9J9XgH2NHxDlEYP/NBVLhnDz5y0bV7ZC6VgiufeuiSg3vv
`protect END_PROTECTED
