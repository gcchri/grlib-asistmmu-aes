`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4FEmfsOQ2FjXsFHTxUfuq+CL2/sh0MD4EmElaZyJxjxa/hDn19OYKxdQHl26e3JB
nWmr92slO86OymNDvZ8i6VQdG5aQML/iE2aqsh92Ed8zWrGqI6blHXMxV/poQAKa
h9aRhwcyMY8LH9+lLkAIsU1+GLKPSxT0ZfNmuPqpxobdJNOsr9ssuwDRMvXO3DDE
mNfZJmxHyWVB/4Wiy/+wncrC8bIjMe3ALDkgfcxWlXRe+lceE9sphBNQ8aCvAzQ6
4qcQE+U2C8ZDwLbz+Or/SIh5FlhxKBat0aBLo04EAZS4l9Kp3eQHPiMvsz9sYpYb
Iq8gUUasiC5dhXuyZF4MJfeRP7gqy5qIm3TjM1Mgphgrjggd2V7eCbbIzJJuP6cf
A2Uc8ylBRU8d70A0jzQILzy4JCJSOBZ1fQBrH29Hb+0cKDWRgdH5ZJpidn8BAZei
xI7aDPceTc1pK+xaPcRmXDhynm7RQ2d9FDHns8Nq25FMmSWvnVa+LXdAuozlDszy
tfHGRdpZlt72X7whXEZR8VDQAHwitUDogP7tLElejycl40yIy0R0R6eIuaO9SDsE
vSjx+9W6BabWSE3vyKnrtqUX/PeYRh8g9Aukku9RA6Dfqm5sIq5xy8ruH9XR3s12
Jw5N83r5c97q54k4nPqBf5sf7J6NA+dSQx52PcpbyuouzJEIqv4sp53AAvhPFWi1
AJ25xAvJXBtuLSEyupKYBx6uVtpvwdseitz8qWKnaKRfeQPwO4rKvdDNXGvYVvlo
S0ptTTcOEoNIfW9fwcCvgVbwNmT077CmMyL0DobKoIV4x0Jb7Pfg2ioD1C78BZzw
Qlu5CBotevtVYxNfA3EHP9b2r0qD2hovATLVllQVg7a1rkmWUjDCxZkddA95do8H
8OqYr/fMRAHFJ27wgCOzaT6CUibFyBzBeMPMgxKdum/LH3BQa5GMZKDagwC8/sXH
FS4DE8HdBYCAqFy0MGDKGU30+MKfM5S0e+lpkdDFCQOGOZqYdLM5BkiB17uv5DCl
U6CgljbVHLpPfDpbasIVvPY8i/lyTmat7jJWxOiUESnjgz90xIwVkofNVVlTerq8
S/qOnQ2D9VVSM4bMe+AxyBvm4p2UNvsv2AxazeCBVAPNyjONEHtMN4/iCAOvyn7X
07vFhTK7fC6SmncaU2dzDks2vn3CGeBbsF4wfV72P56+HXaPT6uC8YlFzuI4OMFK
6+MzeJlVy/DmtmBLOOWlmP6Gzy/9iuQxmYGY/19i4X9EDlglyAXKhrym4YM6+ro6
xm08ix+nptkFnOZsrwQvMkAwr3Dnv6CcZ9QL+jXRNXAaBUhnfgY01/aZ6lGzw0q1
aZumxSBy+eNkaA0dpbovZJuP62FP/R8Rot2AlnXTjN5jUiuBMIef9s2E2oi6WDiJ
Frt984ox0D7BAO9LKI5PDzdEf1ZxEjz3bJVfqyGsvgoTcS+jdpoDFragOoYUTcsY
5IgOiKXo28bNNz5cLmFHhdwy1XaY578W0s3336fxKsNQarRbo4D6BYzOQJ5Z3cqI
GlXZ4B2NMXo7ELIJYRrvSUSWhua75KNsnZj36FxBUHmDAnX00Lk3033u8f8mRMCU
YLdTtU3GMQj1Bfwoe2tPZa6F5iTxn6VEqFOoB9oQgSxq6H6YBrB4UgK1eHQ6XXH7
q/RI0Yftx8XO1LLe6zLalCnpl+ubD9BfwQexHaB9qI7GHm0ovi2gQ/HptRyn3vZI
JO8zgtSENafaYf9kYNOO8rfPFy441nRXGwqmHuICqs6fc5TWufBfoBXISqelb7TV
ntvWQzlIYXKlF+rZ/lGqTXDr574KThPL/olhyJ47UXht7GaB5JrGFOtUv7WSJsN5
ttJpiNSmsc+KQVLVbORSjmI3wuRXu8f3BwaytpN/Vz3ilxdJdXCzKnEu5ZtLq1u8
jFmXNuSw3vkqshOWqDhZbihohqs0P3jdtj/HmUY6mav8Nyuu2eDuffUvxVNX9Mmh
6D9keB/ky20tkE39a+8Ma6gk0JL0UvdP9fgBOLrNw+d4Osz/3tHViPq3s2gsvcTA
PC0eSYWB1Zc2stOb907W+fXosnhzoiuogcXYJbkIn27VlOlj+5VhGsUSvZj5tmKQ
vjLmcn/BYp5MkRp0ggnkBXRJXd03UX+Pq6jYjY5/U92yA9D0gtCIkBfl2LbR+n5H
bqY2GGgKIyURom3ymhZx+2pfwzMxRhGLFeJ0ztHhkDgGM4QCMok6v9JemYIGBlhQ
RLpIyaMunQ0C2nApjUsZ9aCdh2txeFQTL1ym+3/lLlWzwz8AP2jd/uCKyHgopAdz
GJmTf/Vp33H0q/YUcIhz0J0AF7zoNq8F0od1V3Y5yhKp9h84MX8IJlovQe/u/P0i
BYhJkseildrFlv7rQ9i92yc9VrXEUGlnSEtJ0JxIQ/TyjK3b74eHH3BrJPBTidgo
2RboA1QI34HFqhwKMX0Fo7uTfJJO/oVSkjDVi4Z+Me5eHcHX3Iq9nS/1I6et2j/w
jlJs+QSDZuc6uoh3GpwOKeN7OZZc/11WooHzeQA94wGDbEZpP5cIDsp750XH66Ht
ZenrNqa3qsMOoaN49w5W+gTjHluQo7w+thYhI//HIZdU68i/q49jmb6IGNivnNse
onkqbMT8BFJwivdv73kVVe5V9aVCOJRukl8L3kEg4OSUWKS/GXdAF8mn83493uR/
UKqCu5BS5iTVvfpE3cxfjT0YKPVA9I9WgCbuF1Lq6XdPQc7zG3Z/b7uI4daqYXhw
Sa5808jcoqSTFLKqZVdUueVX2HRtMHkVGl/w7Xy3y6MHH/YdC5jE0yZN1VjBhan4
sju6TlBgDGhvvQWT4C3gfHzwZWOJb6PJlaOykpYMzduESmmD85bFhqRd0rT3ssFt
jVQGbuaitkmXExwR7HV4YOXKGzl3VxzWABqrAS2VvIXUi/qOmkLV3QnvwVbs0Agf
/v58ylhDojLD1olX40JHpTP12T+7diBHdDQcZ5Y/CPRsKm5Wsls+rKt0l6ISkXxu
iTqd+PDY8oLGmGw2BN5Tcx3YCL2PkX9IQ+xHmdgU3dtMAZaAIhz7vg02s/ZAuqAm
y2jGQu9Gr00PGqFljJB75ACpofyeteYKLH9gVQvAMImc5b9O3YG80nPZflFPVKkj
M3pgakb3KYM1uP7oAsgRIQyQGko9CJDex24TNZ1Wwp0qJ0/2Oo+lSigTGl/RVMNM
sJudTU7AhnfpFQoVWoZMOQq3RnjyyQDPQzn4CrsGnC7cqMZx/BfzN/jVRym3RltW
uQQaHp90K0UngDkhckJsNYmiI2q14BNC003/6/VTe0gyphSuafXeD+jtqiVZ+WcS
BcfXSI8D2/pUZdvYw6PUgopMp4XlHUMwQsGXnYLCqFmaVZeaW48zdQNcivv1q+29
biNTVUhZadk2LwkY3It7DshECrheMhWMzSu+LciCgifMmdq+aFQ5SND9lrp0ck8q
YH5YM4btxpHeRiJJ6e60PLBq3zsNCE9HRnoGEBq1mTYZ68QcscRY5mbbsT7qgYVb
qA0GfOakb/CHnZdj/4pK/tRpay1indhtZPZYN71xtFjlLZLGVTmtcVTsWHYnACHC
1WDQBUIVDq/5lL9aOapdl3iQzxUqQeDQIkYhOBr5dCF3aEb3fPfG637wayAK5OM+
H8i9JCvP9FKn+G+sYaApCyHNzcovZh5uIW8yYmQ16KLTKJUAWWQ8lZPx6qmyMUao
C/GyR0BC56PR5UdRLQxfRcQDWhXe5+ZEhRsWrWrbu6ALG0qCF1ZVzUOb35eeJ3KG
jeXaMpBlvc8pr7EKmbltUdPYwgQIes2SoAkQvQPBkhPvRR3Jm2FpilDCa48MXOuJ
55a53hwsdLJGoVykhNtYWg3V+DOM5t3Off8rLJNmAls7sRPcyrfNCuvAvfvhxlh0
y1392ciScdyH25souFoJDFKOv92syE0ZtBKJ7eC3KHXtUn/Wk2tJIuPelT7z48Ay
danMB+Ba3ObS8MCSFVCAp77O3UO5YIDBVJ7ZjuaAz6qA/IUNElMPBlsr6HJqsfwZ
ialU6kkNKkO+j+XBV5MNfkxFdeXuixNtbW3bN4umsNpD5FZWk5KPyWYZUFTn38uP
IbB+LP125bXd/6X7KrlHWYcqHPlLXa8Z/TeRozDMw1M+odvf1TXHte75fHKZ3/QR
7OGglKmT2u4NjFP9tYGzjLyUy8NvwpGnATINrkbd5u4mfMaGWlutLloAe+TVzcvB
UxmDwajNn2p09mYPIx7nlDKxIZaeNk3lA5GxvsPoSO8WsYghTMJeiH2YGMXzf/T8
U/CTibBL5rOdQgTOz9UWQwh/z+S5Pzp+wIE/5+odvzAB/1jgHeJKLow4NXAGH4in
avL9n0KsE8OIjJ9umtLVJlLl202mFNAIU8qeVO/V5bBQpTMmB+mRe/akB0Kgmp9l
QA1XK+2xymcUc608Lhpa5Key5i5e3oOntHe6Txn8Y8O7cZKYvGTTwUk8jz88edPS
T6APCPBm7XEwoOEJYQfw4koUl1EeQ4BOC2dGhf9LaCZ+otjxy1YgA+ppR8ClZ9Al
QhmYKkXV7Fc2gAJHqBZUCAzBTyLGEyG3Cihfq6xeXr8OExW7ZgdjsBGR/Mb2tjVh
a6hYa6rjOHtzlStbtgOdyknDb3tx/yluoxhpcR9vet5YRp+/hC6+0ueJxzVmJAn+
73HG3tVNpuamgIVnu7JGHHQ84CydAZFETH+SW4+CxjlkOc+2E9LbjyP1KBTQSUuE
FT0i1FK7G0sOr/ksg/b/+AdYKnFoNXxMvKD5VfDROkt0sHeAkdFmzsEGXXlCt8TP
sUXBeuN9DummFUnXTdNDosE6tv95ZiWceaMs3x5uybbpreVwLwySn6QEtqE3K5mv
5IouWrb2fSid31nUe80BxnWB3wmUCf8b2pQNcYBF5Lp4X70cq7ZeAC91Z+ffxetH
RuBpPAREDPJ2sJP90Xi3eTcsv41+WbUBlITtMp2/seX9ch3lagX0kd7ZLATmItX9
CwELgfvxR5XKgKMcNv8m1s8dkmI+FA4XgybHGkOkd2bUiDuKSXXpiVcDu8F1l/pD
4bK6dRhENz0s8dygDrvCXaW+ymuYGIa6Vku17lAcD2Qb7xUImJMzyJ0LpZng3awk
nbn+22DMIQ+gc6P6SxbFUA==
`protect END_PROTECTED
