`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wN5fhKE/K403981JBkgMDDjdV0exmEuENgW2W29WcbuDPZP7LPLyU3X19z+Ftula
eojINKi/sWjjF0orwemY7iDsViUa7GuHj8mDU6oZr1LaCF77CRyJhrGEUVh0wkG/
BdGL8OhYWe4nk1Lnxsq92FPQURri/WYHkA3HiqIyF/AvLt8FJ3B8llQqd66PbADa
wkvEcKZQxX6BeJanvzZ+cU2K+C/5IETI6CFeRO4tDoyKFMLzRfMjUCn0EukRwdZp
YVdcGfXSTgbdmntsa3B1I+FK/OQgPp6hHSEDDkCjoWXGX4THJdYoDyLlPAMxlBAJ
PDCuGidYfhngqXmhaUqVycWjzwMRy8PFVuXalgyduI0pFvlxrJM8cLrO07PZzidM
6n+PC544AhK5aFZVTw6fwBdw0wdryA+5aIkKpXrZAjU+sNtf0NGrdFH0p/y111/H
YhM8IXYvT9G/iNCJ/bycVAC9vShSuGHH2u7ZYaoxPBLL0Wa2VHkvOa6GvdFw4n2S
1FWz/e4NL+LPmm+A8F6PzadPjGYi10RnkaLXt5K77oU1ARSygC5jLzbUYAHCSn1E
WfH8YAtBuyYmLwfK7S9QxagY2QxBj8gYgiPH73QN9G27r9HuvzwViTU2yOoZTy28
`protect END_PROTECTED
