`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xrsclbJKr7UtmCb+6PFyXfIaDOWXvsZTDjNXOg4EPb1o7XVf+x/8P7XzA3KIGedE
fZlvn6DglQD8g8zosbCdPnozKDYcRlke1gq0NE0nsi2idCGE/gHm8yOrz9KmSYYB
xpt4/Ryubdp3waiohz9BspYWB4X8CuG0LTfpBidFdgH8hcgEQDJm7rtOeZocBq+2
b4E2OkKXxWUv9cZuQNeGUcFEDEL+3WDTGEFAUG6+KNJK1LMCU4o8Ua+nzHerP0Rs
403ExtbdDGWylh/OGVuEIh36WJZRJgoTvEZXxcFM0dE7sO/NO5WFKyuB0KcQftUR
ZFX1D1Y7w5/X2/OAe2A0jl5pupSylqFojkTX7GRXVKY8mwVEXJ0nkQltXpqoSJfb
HuJuhY59dSR52Owj5FIyP9IOumSyOJ4jW3I1M4ngQrknq2MxISjAoLEgyar/yy0U
v3NGQNXZRWXL1licYScqMv1404NE10twil7MiW3zuv//9xGcKVV/bPGlEIo4A+I+
pKTQlA1NKPWULKY8ybZIa3C+KA/JkBLu2mkoyXyk1oJr5gu2dBRvlppYQjIq3tfi
`protect END_PROTECTED
