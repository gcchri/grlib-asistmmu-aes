`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3mh1kEqs3C+dQAPKzEEazLZXl5R0yEJRbBKXPvQ+2gDnz2lqUku+5F9n1sUKuYuq
RGQGcqW8QKwd0aNSyfouK9ygtee3pQBDp243bY5Ki/e9IQDw1+rVwsewvO190vpD
m+4waucqvr/LRczJARx6kN4vkS8L62LCg9NxKYs49ArTrsZNR4ojER7yTd4UvDZL
UnV02/aebgmr4+1W16b6H1/jkSxt+P42O5GvfFA4YTPG9RuomPldfXlXtV+Y0N8O
qM8IcC92JwfUOZGx53HUYf+YcnM9CnltgfUeEi9G8w03wGN8flwPFtv72nMPhYpj
aTJpangE80nCXD7+hDnusCPRl62dXxpFhOBzCPvR6wxVYi7WtfE6b7o3AN2xH+HP
eI0OfosH/n98Jg1oYGglGg==
`protect END_PROTECTED
