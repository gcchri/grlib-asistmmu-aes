`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LB64rL64Tc9k2rGSEyipCN7/POe1p1lUo0EiRMOCsz8LBbpHoddvSWvKtuXjEsnw
Rhm1fcsuyJE4ddKHyZ0B0YTtTwQvW19yjliRRkCaWD1qIc+WIsDoQwRoMbvhogZw
KyKWfd7LpXJ8WhHK/IOUkDxPB3y+l1G4jwU4n0ciDo3PAvMj5ul/WOSF5H04K6GM
vfdTHLj8ES9VpNzAD9/zPsfI6v/57G/PxxTssVWMfGt+0RisXUPuQbLrwR1WzpPo
3hc2h76ci77dua6QuWpPbac+8WvnFX152nyBiCZCSeiqOySday2nvc/JZ3E3jiU7
JMSEynKZ1x10KZiYNxAE3XPNUSDsJ6qK9vCM1KI/MfFcewe3CRM3lLBqejiVSwRg
kZRqYwZcGikfjtAYbSWvFVFSSPfmQ4UEl0a+wG2UpSVl0/gTDcJOxg0kI/83bqAF
BrHvyVA0VAHyK+lVkwPcVchLVVL8ZuzZHJghd9YeqZV/MhURi3JZx29tqOmK0m0o
TSu89FF93m6yfSn9WfgufIq29teQsDQ8mmE8uc/5pliwKhOKqiz9SBOtcrjeS97O
kvoxvJtnf7BAr79LU0f2mKbnYAPhyM8B71vPe89Rv21iTHslAwg2m9PYSZdbQ2TL
cFahRbvwPEVvjorCTP5e9UPpQ67LHZtuWUlJi4OfjfeIkwYPssq0mN70nbfT/t7f
2ariI85CbjPLqnHf8PJN4xnlUNpXgxoR1FpKSIZKRzt29+R0yb9HGfwt0u7z6QxQ
gjpNYHirxav3mtmqz2+ze13YwM3POp3TNVMxu02yagd5zp4c/2hCfLBrbgO0u5X2
TXuUfvQjyWwGYqcNu8mfPDIy56pzUkp/UTuANKWiKeU6qB8Sc52Yf3YU9eXnUkfc
OuwiUmzxxGuI81dDNr29dDWW9993a6MMoA323UG6Zx2G+BWAA41bGu2a8MuMKQ66
ieqly6fVcA3WAV/vrxbnE0UBDtkSNWyLGtR67LC+Ie9c4Yp5skNt4vtbBrkL76dD
`protect END_PROTECTED
