`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mUN0UDeNX9MbbV8sX9AxvVjH+yOWnEwN8++Q999nqcwiAB4Rp/E+jTgO8QuOPMfu
/4QxA0hkge3lNJbGE6Q8b2ElyjAvSoUKdE8f7HXq01uJHF+dmNEqkN8sC8X/sG2+
GYtQ+ArnlxDGIwt4VFf0eTbrSFUxKEHgQuNm7ubM81mYJ1Ze74n5G/qMG8YFo9Ex
VQ3cuBvwqR0fQ5SnTuTJCTZOLEua1NmLvbqwdnXmYLC9HZNTGwyh1ZzNfAVDE9wx
Dad7s8opswfwGKquVff6nAqMZL0tiLA+Re2yT617KShEqSKRBwtEwkcsk4Q8g4Kz
Z4aGVfhXuhuziOVaFpLnyBoA0mPnwxFxKmFttTd3aBUNayzuSZ1gT+XQvvvo7WtF
NHD1XEh8uXP5crMiwSWVeNk9FlIsRfgCEOSpVldibWM=
`protect END_PROTECTED
