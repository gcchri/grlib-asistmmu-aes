`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9f7vxPp9Uq74EHYo3V0LyF0J513HEZ0BQ2ShztSLsBmt3O9knAWPldtKA7WB0kgZ
HA14ejeADnabD6DgaINdHpLms63y9RZQLgEFsOaYxE0jsFhlMgOXxdKAVQu4TpV4
Ue8oV+OLGILs659fnStFzAV2202427nVL570cvKswjqxbotY2OrMrav3pBh3mjfN
nM2mpXRrOGFP1yC2d40VUGvJ3+6M+hoVxFAXkOiIHG231ytT0IgKx6mWZqjBsEAc
W17fWGDOAHQxHxezEY0sOvqcQ6EFyLP8FiesKbA6rUgRckWKvKjpFfAyyb0Sne9e
DLsb6yPi1ERZvSc+RH8P5GOyfmv3sXGHk75GclMNbh1eP04HjFBBWglrs3+6Gei9
nUW0NMk7wXe9/B1kiE3Lf7W8AQGujpuVqs/nilDl83dEVhbJVrk8p+49S4Hju0fa
`protect END_PROTECTED
