`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C/1bMqH/ba/wM4zdQ4kIU9HrTnVsgccM9PPCL4SAOaLDe0JlIcXvTdHo+zDDz7FN
0s+uqmRkhqkXygkG04uXSuyOEwMA1vCEEbFqPFod/RL6Kq763TXvF9OCxJnM/Fhd
vBiU0PnRZzamZReCVmsCeAlOUXQs2ArRujHTKG0QSB2u6sSj6GlmlEcwdgqu471f
h/Lr5SWYOgeJkNJtWDNJpHxLOPPrxAXelIkQ7gLysI2z5kq218c5ddozOvAVkabp
IPb9rQNywqREylFfmP1T72FPTly2zGEcEvLqMRIeMweFRCCO0TU00MNudS8AvXGR
srz0Yt+U9neXkWpFMcVtlRl7UtQFsoRLbmMbAC5or97hwBsiJX+mpCU2cd9fDxXG
nnq6tzIOS2nWJxE+xJNPErhFblZ6/slPiIj1XyTsN9asQ7sfSWoMLVsHgpf7ZlD+
9eKdRBtOQ90MCZ4jo1plJic+YgoDALLbkOsppU4Qg98=
`protect END_PROTECTED
