`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pgLUtFhWL4nlrOX6aarLVF/zJDN92H0Snb9FAhJ4GigOny94U28kRV5H0G74C1Rg
ct0ZUqIvXe0mc1wMozanwLIpa12jhSuSJ/R7mdJo+R0s1B72dxgkO6VbCsIrkQV6
VopgYfPmHlaXQqi32ZJySOzvrbD5BuSgn53AV919/XGxlphFPV/DtDhriR4se5qM
Tp1Q5J06VXT8ulT+Yb5+/boD54jnQV4JzIndij9Vn1LuEtfe1fX1oCxdxB6/1gSW
IrCFLui51gHuzA6jTpLONHsx9PEOqyHNhARfaG+JnNpyv3No9ZTfPeG9SAvbq4JS
dKd7OL6mWFvHVMOUKxdT30EIqrNKSd/XURF+fd+w86xC5Ru5OjDwlzW0UYzp7X1m
OTjiDf/5K791qIA4uVtsEdKE5XX+W/bv0FgEPXC7YsWMHZnyXk0FNWJg/P6ZJAdP
EmTCogUJz+bvd7PbHBE4dU2w9fkPvk9ZKk4jfH+2nJ2sYq/7+mCd6r3DVbWi+8pu
Dia9CJNOw2RNLf6w/ZGVIu8L3qMTuFBWa/Wnmj5tUvsOr+/A77Jx8pmxqdA9qiLg
8zrtTfR3tN2TTUTS/MccfxqkBmBuFEbpF6KQjURv9owsPGCCDn4d7E3rTbF9/z4Y
rzjlp2G+HjaLFBUfBXCe4qmIhuppoCtPWwS99XFmxkKoCRaLXX2XMMrWvplqIU/E
zyT1XVh7tBLSlD+oAGzOa7QKJ+JgReaFvQ9ilh7uUbhRzX3X5pT+9JvLI43RxyF4
FEpiJP4BYoFtBy7s7IFYYxP1Zqm/8ty/J9fR0oiCZerrX9LpfsmC+sNRxf5tQvMS
fTlzvzUcAD4vXo3YekmK3+W811wAFMIqVJTaA9mocjdatoYdz/+7pnvtkRFiEu5b
a9VHKjyGGi6LIYN7Uslt+5oFc0osLZaYdUJgSgr+ct/ydhrRd34K1q9uW1i+BTlc
1QzXe+maY84uGV//ZG6fLn52lym4Oevfv3PUWFF/l6xMmL3LsvV7RMn2TXsru/h+
GZrSbiQgcyd/W/pIOTUnR/wnXn+r/AlEV2tpW+kpHht7b2gsSd7AqFL5gMujpT3T
J2kabDQYXVykrSb/RHsrzcweKABIyayYHC5XAxoXY/TkqbOWN+xcLaR4eed2tiU6
2MpSEvW0RcUlZSDSkU3HoKNDLw02faKk0/KtRP/Lpb0rrh05ey1x7S+lqFYv9UOW
TN5DeWmUX1egzuxDHkyJAmXRP4EHytaDD1Q3kmcbfAW7JOs+0LXNuRWl+MS0DgMT
CH83RFYsrGNo56Od5Cu4tDFCxKYAQbxqB1rzaDOlb0S1gFTT459YFU0MIEwjsXfV
1EoiVbr4M4IuUNhtu3fL1RIiWecJmyVD9gFLAv3zI5T3T5yH48R0oiR689c0MO2M
pkEO4i+ioaZ7d6ZY8mXyatjaDFV/a+RQ/A/mLqvzUEMaCBgLvbUnPDXuF7XCuoDh
xuNd1hoJBZWu6BAZxU3I31IlU86SK71cIeTwJ0VQ3Xgnif442L3qB/3yLNEBNfCf
rlBCj0340qhGQsfe7iasTEFmez/VJlBq4LQUjJkMe0UuiISXbkSMlp6A7EAEaOzy
YwQJz5d22yK39pHMaJFHEf97pueiI39dTYQ27PhWGISjtmLJXg9WCW5v/e0haPXL
aBx+lJzEZpFSgkOA2Sj7AYKmtDmQ4pAzw7qq6rT6HSJ2KMnX+gttCNlU+En/kFgR
bJssulpRtLLdhN3SCq9FZiq+vLmXoIoJ9YOeasP1iowGpQ3OXgPbsBbi0qXOJx/d
0frQxlgYJkJesgWywKTsLBd0ef8lnfCUhsu2OeWQ3jYUofAZxOUYJtg7JjKsfJkS
9GSQT7PtewETB4TFPsdb0VUQkWSct7YHlqLn7xZvfyOVdZRe+4Ara2AU9DB40hnG
/IDIkysza495GASUUXClDvl61V//eIc2AmhU5xP5f49hN6LZC/lq/kH/GzOHYJQM
Zxz5/ZPrsIMdx4hNgjl42O919NJA+l6RJhb9xDbP+P8DtfFHEmrPn8lUy4jmrv/V
dpUpFtv0Ie0zx0TC8sz3n5mDYWO9wfpZ0DS+tncglflcGWUzOEvqsghuhfdT5JJn
1/TSeBAfVpGHc3sE5FfuSxIpnARLOlNCj3SNxO7H9Ty56xq2n/6ZNAb3fFzM2UY5
/0BZU6Jq4Y92AdUjCNOtISOqKNa+nm2korP8GRT5wXbLwbtGSklbGGoCWHqmsx6e
i6GZgU/tK5qHiUj4RtCztpStc+kfNjuRhEVoS834r1X1ZAEwRbxxhjXjv+CRfqon
4wfnJksuwIb9LpsGz9L8ORtjAO4Pl4vkoHoFmMluJsKmkY+q/NkNGWVG79pZ3akX
ACO4xfqfH9pzf6Eiv7Cd4VHnPmzXlTLqgXv7RsMeNREbsgQCM3xQIjmN6NAFVauH
VhCpRirp1c1SZjEga723VxK9Jr8dRlgTYPsxw4ZKhZuDZhQ3b/VzjojgnSjy5VZe
pcE9e1V5DYp4SYYRpuSzfZ/qADzjLnZ9D/HJ6z3ogIIA3BXFXC4OxTYER1XV8RaB
J6kfC8Y3MshwwGGyBb1wsj/8Vq7RyVZO/KHsDsuap4wi7piznV4DRgXuyL+WbLOL
c2Y6fHIvUF2ufhNF3j8WVNky0maQR0D80Vsk2HHA4FBDvb3dflbuo5SChS09C0BR
F5S97wC+wLv05i3ahvDQKSd7qZzfW1jmBnWObzoXqSGQu6pI04isJX6BtmRheHeB
jK4O/OYjqQK0q9paph4yQpmGPIP0BP5oz6LeqNV/x+AC2yNi7e8+s8YtmqTDGAWy
ly1HlT1flIum2R56NcaJyDfldlVIIYv2LLUCJV4IjS9eLnauDz65lDCIdClxXVRe
wwTL7VG5QGKTMnJAY9dOEtqUouN8MnrfsQwqnF+OEG9I4nZxpmgRRGBI0486KEW7
Jw279z0MyVIX/a5DdRGMzzjT8oX6kVoOMKoC2mcTO7cQ9sP+DtdDjFATcH1098bi
uCKQk8nK9xmXe2UC32sPIjxSyIZF31udQGvXr77CIurcm7iIM4iaRbCYiTNtMWTh
cHbKR8AS2yCcbeeUQdIbS4d+zgbGDo7mdWSvrXzM+VEO6ji7pBj4nyX74riJIhxG
CQmCUb+ZXEruZ+a02P5oSuvg3TkuRzn4bL8FgcMb8OJLX00/LK9Y348CSiR2YyhO
UQH1pB/uk28Gf69zerXVsg==
`protect END_PROTECTED
