`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k+0Fe30dHnYIaoDqbaJIiegdvb3z9EpnpUrnPI7rB+HKPsbFv6ZX/Q0dlX4KxsHK
7Zo9DvdCQTpyIQPvDpNdat9V+0g2Lga+gRcOvJRQh8lrTt5mqCuvrm8rGm0k25rS
Hv0j8xDxiZnjcWzhHEq/Ba8GROScE24dM1utaiDm2ZQOMAfAqNFXYLky7bsgNuT5
CRQCimGveWtyQmzXcWAklbR/vp5BsKTFaCN9IGu+VCmssQaivaYXQ3WIBL8hWovx
aE7qFmRq58GhvY9+X2hZioCxbYN435EGllB9vfgiidADaZ+613aQrtJQGPBzGHX1
0ntM/fMThCjghezUQUGwZB9ZEoSvIqoY2Ft7g8tCR1+onJwSZIzE+Lg0m0a7cDmj
AwNg4S3icCbKrWY7FvZTR9/havo8/kWg/DGiqm5i7cy4dlnTxHJvx55NB1iPl6Th
`protect END_PROTECTED
