`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HupCJsO5Z0e2u6MYH6LlesGHNdBBekBlFqhoMK3BLNnMY7iiIalo8tp/RfmIp7rn
aaVYt6Vh1dnfKlkbl2SZoyxpOvg6Hwji5vlk6GtwEfVWukmTB88FJjKPhf1hQP3B
++7EaCCQNcHqmY7VvubagvAbQpoCBH/dRgtcLavSwrv7wK9V41Gi5XrFoZr4NRsa
sNTrFn5LA38VF/pgLP4yibvjfmGz4kCJm+FNEzOyc7SBKmLWEuQVB+CfDPPGelei
HMd2B//GdMJaXAtu7oKHWL3ZddvLixMvNMqwnOm4NzCFP1BMiPV7NCqW042qvG9Y
WTSiNGrPGBqzNTxQEuPCONnNnMyVqoEdwECG5FjM0+vaC6J298RrD73j1OdjjqPM
Ie8u2WfXYf8gIs85TzXuhym08K9OST5153+eq2rf4KFruDeNaKpmq4MakbAxDJg6
0BkncPZTX7h7Vdev7JAxnFogSnKVQe/wHUv1Kxgl/qJD9rRsunShbVhn6PeeGrn/
ji/osUpNNSdOKEXnLAIos2jsTSXRh+v7aYPpIZUfA/oLY1vHaohctkBXWyAe8/Vb
zZj5HsVjn4eapiKuJNMsACaEPMU6smeVRRXa4qwZfaP8mvkgFuHGknk4M0BzWxZU
rvtPnGjJfxuGl+fA1WvIv2tJNz6TXPQ35zDzUKM2p24yus+sQ6UUr4ro6tDkWN8L
DgLkDp/0Klxfc+6n/lFvbNmQndUk+cSmVhQJc71EdyfU539sK877t7xbo/zxdlF1
BbatCu5DOpI5TlVOWMdnXSyEdoZBgySe8JoZLL/bJPwher2pVxKeCEzKx0C2CeHz
mXqpnTECeuDWEZNWAGb9U0bFwWeFaMjOjDPtebhC8usL3SyzloqXpMfM+7rVfRc4
Cq8CNLNvoMCtcAKqaJvd7fqErWtZvJQ1NZC2vwiv8Kf/icLuPhjN5pSolwLD5YAJ
aijPHsGhYtSbmtZ7YEp5lGZKjlIBZh9yR3xbjGguklHatk8fIR7MTcLV5Ejx2DgE
3AkWaZJ9nWufSqZSxjrbPwzOI7TETDkaDgvgfNWBCzXSlwEUiGddWXF4hqoGSySV
ciUxN5xq/C8MpIsNeppyHxcCfBg2IFrAt+VeuGWRg4rfqbXcIea+8Gpg3fa+y2th
+I1GlufB7Z/pvK964hBPx+xUHDBaE0bLmL8BTwgNI9kCcgi7H1i2L1PEitwn10ET
pe/AoRhmTlmu6IFOo1wkeQruYqQzDNiHl8Tur1hVGOIBmUtckJRxsKlLaey2s4np
V1bL87DlA0bwizJaGkahJAwFJwo15PZcEmo2HKNT7hIBdEK8rAPGeVS1Q7pftJBS
fjvwfxtNlb/vIy8QCpfe+ikl4njIz2X5YcEvUxSJHTjfjfKQQbQbpJKcd41Cri2s
814YUj0vwWOjXj2PDmgIFAsQWT4xZfUshOXsauluNR4A9hUKdkcH7QI0FJ3sGKKg
D76sM5TB6lOYb0taY6Pk6txn97NlwRYTu+5w8oTR36JiTY9Q4dYUdFumMn4sH+8s
D2/54G0YABzpOmBJ19afo16FLH8lUPu2vYm3dffr2tOevxEn6mjR++Q+xMaebN9C
x+LUpW/Wk/HAF4gOwjuF0oGYVZOm/RG4sStHm2MwdVNn1ZQMIOzRt4Os4udDGj2t
aYncypdFWWPVFmkBnZ2ZTF+04paiqzXKs7sycILIr4L3lO2/eZCQAd9oFkZ1WSFY
WajPvs0QibC+qUonjOat15Sc7tBM4eVCsyInU+h6/HkPdH2pcXwe3fNFlBuVmdZb
WYm1eGA5iDK10wvXe0W5SVNmCnafIWEzitrGI6B95N9DnUcN4E1vezUGFefyOjBb
2uATOQlF8ztiZRnWwUf60gK+slBHLcA8rtb7wj6uUYHwxUcSLLRWngCxK/qfwRbu
iZ2BNSXRyb0qxD5Mf/37keQiEDT1kva6nNFGrXgdPKJZeCHZSwc8RXOzrmA+pxZ8
hxXWr9J+Z3nh7zmYcho/T2Kuwx+c+yYF5c2lUMJPkBvQe/Tuknr3qHgfNbxGyC5E
pdYN0TmVxvkRLT1TybVNtG0qUk1gSDdIgmTMlgZxum+X4dKwitMSn1RcGGjSwsRX
bCF5BVuw/wm74hYg+iOEoHg4j791Fqu8le9Tz9R5CbMRCIgnYUeFmYMenQqPvXvL
Rjp30X605tNn5r13cxn1eFp6aGa0FmaMt9EB1Lko28KVXXlsiVRdH/Z9VHS3cn7g
vbIGk203Y4EA5yOMsNrFlq5tVUuTa1ILmYmhlvvaN3SGv2CIK9LUL+o/0Ba4pYx+
5DbPpx9IP6bH/ViJs3Lidyh0n91SwoZ6xFLtdt56jiVT8fA+Rr13/NxMeLU3CkqP
sBqNSkVQ0NR9rOytOXpzQBxH0O3l3QP853LgyhzySzF48bbirOjY30ue+k00lSFM
zXx2IdNCTG73I+R+bcTbCL7qPq2+z8hbK82s3R5ozrLojDNXg9GyQtQb6afFbKh6
6E3l9/icz0WNcq37dJjcO1h6ZqPAm3S4NzTStSueh/AzyMgY3nqGZbvUcthAvmj6
+nojD6xbsy4tNlhusmLtvdRU0G1ihBrd8UjWwCfCyMV1Z2TcQ0Aj4q78gZEN+Xn4
WhE1Pjt2q9AHP0KxeP1esqXQliAXDdnXCN6G4cZDJrL+b2S59vC91WYlC8ve6VO9
NSr2NHvKiN6EvzIPxzZCsNSorYjKdusCirhNAF1ZDGPLvgQsOcczEAbNdEqxVVGV
0X8BzRH4S8o+1/b8iLj7FPlk8F8CZbbjBneM1vN1pN06yS72YnSpcXffZ4qjaMUn
ZC7ZKbaSgolyE8LnXi1CuM8sKvB77t3D29jEvkk77PVLLtEZxbsr3ClpB0MqtWPE
79QwvVvPmNAFZDd3G1q11Eyl6aYWfcdeQLHcA18/WJCROH4cQ0Lc3A/27wIBF0Oo
kIceY+gudDjjtF3C62ClIYJHrm/FtemyXZN8ciHdE6dbDCK9ZgEfcFZcpkjRv/zJ
WGHiBnhU9e+Jn3R0t1zL65cRBAAckDazB7OIYwPENih6sItK1WyBvqVaQNEECLq4
Ww8k8O2cYAT30lONcBJf+OL6d7x9up+pgkVOSK28i6t+4kr9JkPZpP6kBPXW6kQN
Zp3yn+cj4zBq8Xh3dKn3Jgz5vVFzqzcSov6pYjIhNVNqZtGI/Llkn3FjE3Xvyn2c
faYHuUiQV+G5+hfc3cTLMEhU/22tcW8azG/v7/J/a2DaEOOW/RCwVnLEjIbcRoNQ
FSNK4yZQZdg5e63KeRs4fh2NvMMLI12KBQ42X9Kkq8o3d7M0EtTKUbFqORlyHdse
QZsmQDVtiNM7nako/TN246RAJZlZwcLwPCw+ss1obwbJxiArQ9mxzbRxpBETq82m
gKjonNiLZhiFnssBeXK5XkelmZGqeDKv7oyJ9ICfjpbbV/rQIk8lY5IjBnnKpYhw
nK5Vt/CsBwCVtr0WvjaHgzkUMmhNXL+C1/9FrWRlzXcVC9y64r+oZbXaSCsZEZ7W
erCifVcl2IWSKwp0Hky0qa6OREYOnmoSfW9IM5sGl8deHbuBjGF+etNbpZRLKr2T
dT6BuuKkyyu3t1Pfo9ZYetBBI7po9rpc+cZx7YXiO1x9/3gmAjgaZiClgrgQqzZa
jShYql1MpxUa7HUadGoXmesCrZiHW9abXRlndeLLvbHqxpAiqoVTPJjnCnxmtNlC
wgcTCOWflE49X9rd96OlHFgV5NuUHMzLXaig2MotjApqi3H8ZQ+vGfk/TrRQZ5FP
GATcmoOB9+BxyUUhZ/lJLduPWwyIFcp84GTycHsHvhnM589E+eZlIPRm083r/FvG
/9URWsdLD93Ip51jexnBlyS8oxsTH+cwRk4X53bS5Z4efPVfoaLFmhX4VoePsIOP
ALgLRIREvE8S2vVkFax3GLz/acihFSHH0izihLbqSUPYZyK2cl1zLjj5A+pTPwOZ
6YSSthgVgUpgNZDr0nCmC/upVqiyVwwzJTx831TxnmM1Z1fz1hPdV33Ea3dpQctU
lhKaC/b2ca2zcxSzncm24TjXHkkWMbvmW94FLKa4D7+Huylhq/+mEx0na4n8AJZ4
k0Ds3nQ8t2DIQeiNzd6NCXVPS5tlXpzoV7KKKWChWcxNonDEqWtXqk88+DjJYCPD
plj4A/WMCMKauJoKEUznNEzJx2o7iUTyQNn9+Uct/xmS0tam/G7j0UkfOW6IIuVY
H5ExDcLB4coSVqIk7q3vsYXEaxdKFqVU85qnVHoPdh71Nqt2izuuKu6/Cze9C4l+
qZIBoYIih51JK8jib+T1yGTZ4dDpNnJ6mlZA72hwSHRfghwEjR45yybZpcw3nYZr
ghaV30S/ySCFi3hBXd6luJiOdK5dfsI1sZcWvqlS2LmY0sRkqxl1digtILzSsCGT
RSOatNW56IvZxG7BHRN45IxESm0Zj+GpkiztiMacwZgyz8ppxVnnMtTOXtxIrvDj
KjLwtlwEE0fWKH+OLwNqEU65xJ1RONZRLKpO86aBF/YsS5Lff2DtedTi5pBGNE8f
3nYCa62pz7JZ8CpD1BF4RsriXQ5U9yO6c1IAlEwYUc6tzjuHMpT584cQJxcn3Rvm
6gbfge9hbiP0hgn2yBONaO9MGd/x4y1fqGXd7VUwA9usJm9NaHQriKWgpBJaQHOv
Ct8GxhoiPmend880mFWmMCy3Tf4svCGhhjvUUhSITdqW8SyrWb3fMTyRRVVb6LTk
VYzyWVe7mixJUlvX3WSjvoigBHR0FHcr4SIqq8fvdUaaFRShy6B5ViBuqik1XQ4e
TPSJJ5dgm3JbdBr4iGnQjeQrZv/JqgYGiqxI6uE6vXwY7v6C/P0Ec2mlv8aKozna
WsCRfnIdocSlHIGO8zRQrbslLam1MozIZunM3Kdi0xxWTkxOBfGseUdbiWHJER4k
N7cPjDRfyWCJTAdD5JPiUCY24qDGrFCOahZ9OJL0u9qj+GtdrjZ605UCiD/doIJc
bBDlp7TKtm8SI6iESNOGM1KXP0u4dAxcRJa3EyegoU+f5mrmYN4vEK50ojViqN9b
p189fR8e2ICwjJ5gjQ4jTXLKBRINLIEkmwkXU7x7yZ+iaz/bdAbBTvolYeyndoV8
ON3R3TDU3SVh6eG2Y2yNyNrFz6sjgwNrBB8x32fLVmme3JucoU/+b9bYBC5enGiX
RacoH6loGeOcd54KzqraongjZqYx+soaxfx9SHMEPI/4cbuABHAyxkmP64xkPLke
xI3lLL1Cht1vNSv3wF+V7b3gqT541eS+24NkVGF018Wxpwx14REBKy6j8unV/xbp
z9Ycnkrc+amWXB/S0Y8to4RhS15BBdpj/vZzBQIEoz3t6E+RbNwJUfTCsrB5KnWM
sMF88xmpWyCXCZmVQ1o8ku3N4RapSJo9Up4CkLYaFeSp9m1GoF8uwrvSaBkuW36p
R5v/NTBkBG5wHqfcEQ800B5uFYbi7xYqw31lJoDd1/+uaDSAPKFxlCzh5H8ondkK
9m4vc+HfXvWuL5PntMsi4OlrqlZ/ZOlqGWx04ypMgZgDqe3eArhpaNTkFoxb+30u
v+FBPO3iNs9q1RUyvbzI+jPHNFXC/9BEalvqAjYSt2p+t40mXOy+NH9YudFVG9J5
Pzlm32O81/2p5pCvql3n91G9+wK6orRplXQihagM0XPpmZf1OSLiGGFsmHygQhXv
AzWIjhfbCAjMvSBYYK3eF+inwDbAzLfJa3c1MSmC8IbnBXcSqOo/pGK3xh2SHB6/
HZ/TTg3EJY2NOH97d3wZU3zhFBhZkPj7J4KaMp7FwOOFTeqrcITOniiiBjKoMhsb
tCXRSUFs+FyZmwCZGVViZE3zqvrUlaWWKSqT//cNeIjRPBUIBMnzxSfrHo2EDq7b
4oHBjCwblOX60Fy+TNp/BnsobCEL39/sg9tLPWF9Y483Oi15E/JQI1rddl2tcxDC
ASB5VEjg1OIkFIaRa80lw8vgRYmecTxU86wl0RiT4GuGph/9NDd9HsV/aVxaSOG8
ywi4s3UBTfybBDA/RJcmObvjam90DUPdZ7avE4jzVcClEdBjFsXWPYBSf3aQgbw7
jEcxiwXy6rEKV7DogGKrdwIMBTh2PvHfcTPAousj/MUY2YYf+0w7UJ9h5COcWLLK
jycRV/wMz2rfx8YK+IO96Qf0Dee2jImgoAfU08tj418SgFlH92doxCgEjvFAMbCq
gpI1zfo9ar20OILRT9iJk08NNqp+E4F324EkrojHg8Q1K9udlu0aMnZeS642bwv3
hO0ITpzfZN5lb9ohCV9QFQIFOlhvBw88bd+PoxkqOsr5K6Sj0+JcNxe5XnfPf2bs
4qes6JoQITlKbkFgQkuINilZcf4PHZqDYygNVCNbB/skUQumdjueFoaX6hRQrOM7
cImcM65UAaXaKvWsDvPz+Zfc8IbaTWRvophzHruvzGg51cx6m3Pg2WCY0+mVjy1V
DTgbmVdCMawulEE2wstxRDlIb/sNpgCd3e7Xs7dKsCs5+8CGPQeIX6NmJIN8pRFI
k9wOSmB4u84aglBrMVeVqMfc5fXso4Jm0jkr7hgD2EaTCNdFubLqnA+YMdk1VErb
+rPqI5W6QDLcpVsPgey3XVZRheL6wD5v3xysIz97E79R1Py4PYNpvgQDUqTQuSpx
8GAXRyDFqHYWUnZ3Bc9RM1AOu6Q3HkdJWAwzm1Pd7r2WRzgFtTqBC8IWbtDtYxI/
pLzzvyUmDgRYxZG4CY6gojMXQQD4Ibvf7mwzhLFt/iJ4m25auzyAmcM5OhXUmYSM
SsiKD73hD2eLNiexckYCv+MU19wTDzl0nhxJT5Z9y9jb5ef2W8Mc1YSXchbHd1jT
tRSwMGJwZWEXER1eeLrQCEtHwOtNSP4A55g2AxAZoENFH2yvcM1ZOzvHt8way9Ga
Pcvsba0kTrgLXkGJpPWEjVATe+b3+8hDJx/hyjMymEHFPf6Fyzx4EqMWgifH3JMT
quLWnlHxwL9tREH8x8akoM6+B4woymosNhYEMPysSJufZL88Rrd/cryh/1mCPgH0
T4yUXZNgVgB68/lZ4yQIr3lDeDI7MaOxJpesbm0HedAmhl2wJyc08dcsBAG10Lh1
cysrfVsR47Ok9oe/j3Ji7y21+/uOgKmZU+6kNVH+utWpGAculiUQZf9/JB88Cu0v
aa2JIHB1t3XpaqY00IQSnTVXEAtC78HRlR4dm/LNEyQ8Cf025ixTNfVMCJz64Kbj
33j+Yh6cZ8eXl2dJYcqqPWEP7sfhxQuJlJLWazoxpHdMrP0mtpBcFdF8sqqcNKR9
zaSeR2zHzC+13DTnUuFZx6QTw0DrJ2aQjv1BRIfTXhUN4WQe08m8jvKUPr0NNZlM
MproVsNtmSEEkj8ckjPy3XYQzctsQloNUQRCJ5GmVakrGVviPBm6j4idkAq6ik3G
vLckmea2XqPnUXJQ/AdpDYUtf5kfA8JOSkxgrpPxh0A3Pspb4PDLBXKWJqoavRvp
Ow/H1eJHw//ggq9SloM0QO/hA/1C8H0nvHrZiFoUAfrV2+gzOKiQz0nhUbPVceMr
jCBxdhWr44vdTcFmo9PXjVDK6+E0hZ/IHZvPdqn+4tkFfDSyFcyBHNquZg+dip8i
Lj1gcjGjPxmqQn61GOfoLT0T6+TtVLlIbR61q64ECwIWfxhBG3fOY9Ce2gfBqKt0
8YVkiRhwdxZra7g3UhbhkvkGA+vSfIDIg/Bt2mr99gEVvEsAeUWuyu73qqXzyYAA
2CEMyvYBORCjkGdDb/VBIaKVe4TdAFcIzHrVXINOMr3Bjqr7t4CQB/JdatRrPMNz
nBv7tRdtZNmtSDGnZNKugxgNak/jZ81xhuEC5cXh/hlvPczI02kJCsGzGMGs8oIS
i+7VkOb8RkyJtpU49mtkwfLO7W00oSJeN6+oYuO97gAXU+3rI/irDeRxQSofRokc
CTvb0hfuccXyDuuywxxtg3itKi/NjJkC6v20QMPfgW/P4T3GrqTUPWlDIckm9/J+
UAQIXohNVNmYCI6UV6Q02HEmvoO5h+75BRoU67weKxCP/FbiMIcuLglJVltCYHci
EBmEqLYBZKyDpYiGZuiJVRQc8hN2LUJn9CxMJ6uwoIv1hUlZdEj3hMnEHzNc7mYe
tK/az1sA7JosG/ii24fW2OD3/3JJyfAuaWO2bKBdYoDPs8jzCopoAzneo3uQqqv8
OblIDh0pHIkFfEZvfbU9ulA/SHH925AqvNiR8MkQo8tzl1d/qebfEA6su3cYul2q
CvU7ZI8jfBVQpyeumxVnwNdYW7bUNW3cKKi7FA8gsWETghlod24kY53NyDlb18O0
vKa1KIsiNy4qEQRD7z5vUgHMDqP1recrcXaqWeX3rhuVrnOxQ/pFZvQD4JX7pSP3
iqzHknHleewbtPF075fkQIvWxOZ08RKbivvUzkQPdQBxco87rFUlSnM+/mLMVUJj
YWsyBwSnbA05XXzAhwWt/8N2nOsjoyL592VBBck05fk5klrl3VnNf59nxWdWwrn5
vCW+BhFm0Z4jpNPSdVstIInP4FiD259EQLUhJfIBuCh7hO1WqaUUtx9n7ieLelHs
bZ8T6kHbBmKJWfNAFHDCf9rhN6y5Ri5J+LrC7sx5LkcHYtjpObmovjC1iaXUKBu0
xP3vySD2eZHQ5PBmS2rUr5C7qp6iursvfK2BgLwSVgbfVVB8yBYHBykdaNYU6nyW
EiyqfttZevu9PI4VieACYBst7Qj23PP/aV5VZycaw/CdxESBVOs1A+TC+DDOyMzW
yeh0l9oXcX+MNmwUkazASCcJTtYLidXjiUmYEVBhkJ9tA9P63eNR1A/zKxJBCmQI
u5HSWHyb2bRT6lT1r1QOOqnPwpIzMaG1N6QKnTCF/UiqM5FfENq9ulZ9iaLO8JMA
A2+O5FoNmP21jC5yWAu4DV/2oDSjoiB7U+DXy5NAgqr61EHnaZhCGyjv/XEZwF3h
CyXttxkIuqgGH7p2v+UwFgCga9fBsrGT9QDqVGhXt94eVjBqnnj30NprN3sUA4Hl
op5ekWcsarrsSdvvwHmULvfmaSt/qOuoiRBMRAIKqQLLXIyK3kx7wJzC5PN/cmwM
UjVFcAqfnXRpuT9tZC/PAmNkrIM2bYV+mkpSMmTyhLB4M+ni5DIl7vYEpalofhxj
gs52BJKCUgn4ge1UBm1dx9xOnn3p9ktNGOvRUNiaNKOP5QazUku6TwX0jFJ4TZcc
4S8JgYv7qvtiOp9kaLdvtAjNFi8gfWfT+a+eae8Qiw/3rXlc69HmRFJrzNuXA8pw
5P9MO5TT/PbS2eDefByv1LoO+ZjXPfA0ydnFkSdu9cxN5CDhNCJgPIttgZs3J+lw
z1P4s2eWi605nZy5QpJmOvGN8mdtigElSLu9L/u4Jg9wgRV6kK/eKyo7s+t7S1u0
jX5SA9peEGvc72PbkNx36ufcsVq5sgYxKjD3Vv77W/vL+e1pw0DlmWuJoCYm3g76
BsAXBGtCH2E10elQmtgJW0YeErj0tqjKAQMRuFEdab5KxleZJ8bBuHcrmgoWefek
Wr1QMfjLW7q4Qjq0DR9iqDxN9KAC84GHnSVlti5PTrjoag8HoUS+G+ITzeGv22Ik
YN3dRN9WofgUnKdTbSqCn9331halfQKWphstBM95oyjeU+uNidvLnPhxjJtij9aB
TmCB4fCC9iDV3oxFTclF3Ry6bdU6l/OuKtf12TYBe7SWt3lRzcnd6lIZcGuErB33
HBmPE5QfAHfyVFrzoqMmrnAvwGn1fmkzP6vGgxg4HS6lXIdn++Hb46i0h/8+XL12
K2qz+oRl9uvK9wTfOU5ldXT/m1+/pFaDdl+2lLBLa1O2bGGaUkOGCS3evUNGhCNd
jExa5EO3yHWoavNGtBdXrTo1O9ch4kQzWgg222f5FNpCPSX5MAOnS1UwoLt0BL01
xKRlyZxHqAY0vDt2sCmdFAFAB7OEvSJjv6zJZIY/C01fINenphq6SvgOtO9sTlO5
sEWUr82Zc0uh7hGed2HR8Igfgo5gw0wXYLPnuv/iDP82/cYVs8MPCMz6VPx7gr6/
Ytmugc+YVPJqfzIezjwY8aQplEsv2BUZSoUFuJ7uuLEmKyln7PKJPGncacII73Wv
1WB5mjoRCeF/x0q/AOU5KnVExziEef5oyHHyQeXZ/4+FklpHGEqreTCyRo2Niodh
UVAwzDCFecdZftiKEvxLOtzw8S5RO4F7xevy7Jvnu9wlr9I46qWshVF0SrFVwExe
fZaM5MmkDrAT0Ex7S6iZ+QsLYyhkiAPHL39VjrrqiytWJhWmrrsb/25ewnzKVNv4
ausKnH4MdYDGgunvrRzIyDhhan9c8le20TWRqojxmsI/NAhFgqrWzPJQe9H2tWyx
7IfLxZDyL7HbHr2wTLhIR6d8CwM+utsO11Cnf2kGB4zBFipnB68VHAJ0/zAPVNip
paBttiKeokDIi/R5ttfvEScPvQSKTXUZPxkG/mYcLUM6En5IgINuC1l0mwlBiETZ
B2HD1Hsy1rPfDAZmVNUOFjtH44tAMOR66q+Kq0DBft1Hfz16aocHYmZMS8NwcdvM
Vg10wYhF4grmd4mKxWKyeryUU+eishSX1xvi91KuYVLSdUYeNNs9rMEQtp0vtsVU
fr+Biiw4Eb0234wlxXtnP3pEAJprwi1v9Vk82zyV/NkgkSuJo3f6QcmjOk5gR9CF
pUXecyBX82qaN4iYkSqP7JlDdsZTy2h7EDa/ZSqOWkl032VUp1cKLWZVRG/cQoQx
w99eLyqh1px9GusoMynD2EAZHj1kOKGgDHiS39F6O2CBeM/mnDmR2ypudCa1raRc
L9s2pUy7at2dEaJYwnQZWcvvy7nqr/zVKZ1BczMa8u/mp27aM5egRNjDrZmZgIvY
bCnonmCL6owJQ7WNh7i83lvxwV2NEo87OkIVqKGmFkHLLlU/4qiYhUuOOslxjvLl
OrIP2GDFLege9RZiqr4KSztqso6IYXGVMy37Yr4qTQK7CTKAuYxAjfFaVJVdud0Y
qH3qWzeHCxS5S+yxymXvzsx/REETiezsCc5URYV4yT1odjge679/MUrQmW+px6NX
uK+hyUPw7m7cDmu8dQUELtvAzqqhmadYPmnzz+7KoZyduYEYCnkfHZU++5APjUsA
ajuqCCimNkr0cwFZX1ohLkO/SV97K/cDDjn/jmY3yYR9TxtyeAJsnZdX0ZTjWGHS
7g98FR2nnVL3VYSWmsz9zOXs0J316FXMuzStFqYq+a2Sl2xm6avxEyiQrjZR0nhO
1lJYebOToKRdyRt2KQZui26HkQGg9JlBAZ9bdl/+YcBZ5e1ftwlEM3EUUaindTvv
jsGFr1+8oMS/Nf8pvFUedAEc54BtofQdLKcZVio7xzJBMIm+AwOZMdRX+3d7dRjr
p8qZRfH2dIb7yFTeL8buftLTUDvraSY70iF7A+uPm7JByH9FaXAyP+YOcLfLickf
JFC8CEh1Ru+QcKgQuEMpyVVeHUKtiO6yNCvPQKUwWlGcr6NT607Fjh0B+0myTJhc
QI/LCK0a1Ry57zlMNDaM9R3VTQYMdA58YDbprUTPsduNmQKP24kyoFmbrNA4b3ZW
d++p5K1DOW7PnFy4GaLdQWhHsfOO3rKI0+A9QQ1rAYZ5XDt5lyHxiBncF4fp2m3C
bdzKR7SfQ+i/5VS1vZ2PQEN75C3evK9na2jqqwA4nTY5hkrDLQ9BS51oaaG59dZf
ADFqa+HXEmAlLP1CvHziHOUxTk2BvKgSrRcAWEPvD05CB7VRolP6HXCn3VnAb7lP
feAkZxTzMUK+jLtQKinQlAQQWV5GgU0upiEKHgiANlv/ealUuf2WkJr9F1p5pcRa
oCcHuoz+9G8eMh6hg1dvUGzu30tXmu2GpG9JyEeZd1m2NJxMCuyvaJT5CORMrVZQ
6k2pZGOy6iI4iroSYOa//D14yU/SKrtusyyjczH1DmpR1jifupqBQ8JEnd2p+jdb
zRnK03t1/IomYrW5zdXZGP/hSaVr/km2IcTS4+DzAMTTCYJChB1FroI0kNmWk6dG
gAK/4DRm72jfGrYS+cppAqix4NtKsxq70D1xgKOqissmdMc78fULaO2nfppLb5vT
lYKxRz4lk91MRtoX2m7biowc17Ar/rUmhVA0uq5ZP9kwy/2CZQ3tezf/7d9VLCrU
ezoEjfzv0tuvgdBUDY04THexihcbRESEfgmioeybOaelrgKdKa5SpXr9trDf4lul
9Pmttmb3hEYC0v1AGzxfMWf9/CzmTa1D+P9RKARivq7fKiQzT41IsZRHHmdY2RXh
bChYyWRr5TAy2iwj6HorlEwXnanvey2JEh1MjxORm5oXMp9r1oGWqr5Cq2unX/yA
bktHAIJv8Lcc448IFXuSruGn0+MvlI2hfsLAdsj67Z0LfMd6ZKe0Ck7c0ud5Y/4T
LXTjJ2oRSUwHie1YJif2Ma725s6Z4Ec8SjRD6hatzMTJRQsdnVt1OLaJTVGNMB8n
zKlyYQK0Gfjy6GUSHhpXYaBNRDSk6hzSXNQfhRoyv7p/qawB0K5qadSk7dMh3kq1
/uHxjMEaxuPohdcAIVCabbFqgNim+bTZxnjS9Tr2hJe7kX4A1cJmuBFVZau8UzVH
ffICdROOv6USC+vd0AMfzm7axZyj51Pt38MhAZ/2W155CB1t75ZejphNTav16pe5
RrKe7+lCMaPRDraIlcne9NGo2VZQkqm3kN1KzvN0VTyIwePEy5HC4qkLxvy06aQ/
8Gc8jFVqjKSDtFbRM29mzHfp0yg4pNlXzVqXFY9WTuYbwRlHSimUdHrit0cg8f4P
Mrvnl/QciFUXDg1Ara4NxugEJNtsJJq7OEopLeLjrrQXCyEnIemoImF96ZoMbK4U
82eQSsgOK1uJOGD6X1D2MUnmvCs7qrKrCewdKsIoeU+/utaUUy85s5u4N8umfFPC
sM++IlCCqvafz8cwKruQLmJ4jBbcGY1zAAvCyaKfsBMc9IvAq8a4Tc5Vh8C1jmal
cbzEW5JGA07rmWA1Z4MS1JQIxy/HS/XrzfTukX1uQx8X+wFLQjMxp6AnA8djmXV2
U4crocXyOXtEev2vdzMn/kgdk1lGWshb5OcyEY0p5tv7UTDOIgIKJd6+C+AaZvvw
Mrz98mYnPqPhKjCYis9QA86iU2GT3pVcXV1Sw1/g+MtDzDDuqKFtbKS5iQSdG6km
70WTDD4NqV7ZHekRvInphdW7IiTSL5YOGNq7ofuKTpsmrXqS3ZIF3FlKxQhnjQGO
s/aecN88EYGVulR1eLVa15p3ee61ua4KuLTLDKsQUhTjouGsuso9oBeEh8Bqu4BJ
2kHpEp4kX9aBdFCk41BYaUICIys/nb/5M4W8w6rOwWRi03HzDMhsqsCUJCt7L7lr
YCZupkkCHVaKXJLODiVzuWo5fY/4FFinJk28KRDV7zw5hoTb0jIp4B0j6ciQ+42x
E5nVlAcDiRo9y7LURQyquSsgK7af77ld9+7qOV7zd3/RYomAiICF05Glt2gTxm1P
2tuw/KEsCGaY5MLdOp3wjTbcvQee5J406ysGPCaST+C1T5fCPzftCyXHObk27w/b
9XwK5/DUIezYFjZcV+Y7FATxiEbQ0ZbnweZeh5MIERVyHJ5FNwrf+nT4F4+GsDVY
FKdfDUF5ytAwp1NG0WAf5admKovby0694/IcTwd6al9c2vWxBMS8FFDsj8pUCMmB
ulDUaX+3bSRWQ3P6rngaPxC6VSwSuT0O+W/8RgieaWcGANWteDfXf8lXt0MG9rSC
gLkLZzm1UuH83VuNzGwGU772fS8D86AUbT9eLtuTMAr1gRNAow45DszNdHCiADQ1
WDEkV44zSA25B1Dem2eBfHVOKH4ORKCwFbopdwOlQef/gRx0YiPBpa0dhEJIg757
CoaDIKVYvi9GBxkRlTmU9ho4o+Dx1LKF1pzPfkRvxg1iWt0rz5JJb4vH3t2iXn5F
TrItX3CGjYo5YTzfTR+2g9hDX9ES2zHn1aD8iInIc9KndAFk5oAi2bxsG5uEOhHz
9Yh2hcvjQrWS9ysOWuUeytBuaQUnUzsS+smvXHTi7wFJhPurT28CRU7HoudHB9os
+WhMXSYJK6gwcX24jxUIoZkUGAXxz1eJcCmF8DHP/i3jXotAxlUdAgqzJvmdjjpB
mpnO9qFTbRIx7IHWWjskq3vmtO0Y8uSMa2usuYHpoYh583TiBWTx2MovQaipGJIr
VA3OgFBkWZjE0btgvTItvo9ep5OL9Min1k/R/3V+bCk3LM9zo3J4xv3elD4Cy8cm
kp+ptJCcwIrqaMzSwz4kn7lAiefkz+zvI1PsySB+bWxoOggkjncpdMqeYJc9/3VV
aDnxGc+Wlie9hF/GXKNXtBprvQBdlmZmn1mIsuwJ53at63IAeus3s9FWXPZ0Yl6C
MEldPPmblkOruEevN39qV9uQhKcnA1J36jsPNofOPPd1plauaO1j8ya64pV6EBOw
9LCIvXgmu3O51OQ7ho0gtIZHRJW51jAL0lljpMpMNRVEep8BddikcB29gKNFeHYu
Qf1ptuzO1IUG3tMkp7MoElMs6PXCe6Rr6ICfZrnIfnbDOrGrZHLZkSVZRlGnGaRV
fQwq8jvyWn1kU0b4wgxs8dMlpWll8Oxc7zdI+1LdNb9GOd1Kg5s2LU8NsceW92S1
zfVNrY/v8hlnMXEf97afdTnhky+2qaFwdfQaf8zE6/obBGquO6n33DuFk+fbOx8K
5g63KhJ6ETAYdlzaqBBxQYEOfK2Ex4bx9DevlTUvGhTOXc8evpmuNFnIHt2kP++g
5u9zmHKPcGOUgQEe5NHFR24Cu8cFyVDgSslTtlHBvN6dbMxJqrR4IzIs2D7GrSSw
cxNkJuUqOlwGwtiA7Pz+AGjCv1gcpkcE9GIkPdH8SZoEwehbEoRJSdd68IPIup5B
7H7iBih5sbweiDFsbclbyYVKCCGe672cwuvcGgvAc8H8+5d/PR0jKWUDPRO0ZeB7
p0c95VwdN6G4eD3TREY2yXKoDredCVTlWvxQkqkqT8khxSIwOH1zZK5FfEjLvs71
xFV6cZGOrq8jxB2mzEZJLomIJFqLrJEA31mSB0rq+QUi25efbZdMkBb0B3ACNLJ1
yIdyQ37qGA/req9fjNoJthRoZ6WAHlpWWEA6ZPfVsTbiG3YXXhHMTSVZE3DTZSMG
/Kgl9QkH6fI7Zll1NbaSbtJuQjUfJU6wyCHKpQTkg346iQKHNCMroqEa5CFaYz8/
heSlcgtkFrmrQTjZlzWeuQzuRl7E83z8J78HPaV05gerWFgjCu3DsyOrdKxsn1Ej
YIfr9VH0d9hmQZfdjF1Of34odlAOfXAaX7va4kGNrMWrH0w3knHRr/x9yJ0UHwEU
nFc64YF3Y0PwupGWhaFVgLIxBws8IuAtJLQ+FcehLDIAXBIWX3ve+ykGJeICFXuc
dIlhNKoD+ddeZmVCIbaHyYEFZkGyRLkElrgW7hK1MSi+44IuwCiHQN7y+No9shvl
/GhjLKZYbxva4phSIzZidlMtmZiOwwUZR8oahG9sFvoMrv1HQznv00oSehsDoROg
Q2Jx4INmDdbD5GocPw735q4SbbjIsc/QRtG2umz4fltRX39Vrbg5XPry72Q/lSWI
6riueK60+m5BCnPJL8XaxGsbKhyk3+/gYfT4p8acMdRi2zzwtRaIniA6kXaNMWd1
py8ZXmtDaDUVyLwda1GbnYra80NOir2dZqxpW7/qyzpPX1Ns3aevF0bSq8gxJ/Yx
LbMYMfdl3pES8G8K0cVD+eCBze5cNcFalj413scRuae9RHl2fEUULleikW8YDBgu
psvY62mWh6x7RPHgM+iJbMPESGGpZxb+VOON7zncjMvLxX9KGa9Hcqcz1+IEwRBD
QaOf0OcdbPipAk/UjTZlBTy8v8HmX6g3CCgdmBOKeXMxbzHGydhhUkQwKty/bcYK
gti/ikIExLeuxxtls3v5FQkoDCnQjbo+Sw910ijuWr5pPatPlUP8rmRVVLcH8sva
6PStHr3mAjUHCCkii+kA7/LZXi4annxpju33ZcBdSt4ZaGpcEj4F8ztY+G2iWzie
aALsHH2c6PFavC4r4n7VULTlDaxTRxWEx7gYf3t+ihZ88dq0z5wS9jEOo/RGym0j
XbIuGlyci7I99g7gtsIlt/pYvYZYe0s15r/OWXWUA7+Dt+Udh/lnY2AuqjzmQWZb
33VJwQ/Utz+IAkvxMDWbNmQQ7HZq/aJmSzKbxeGD2OmsaIkaNmUSGMu4ud+v2EOR
UQod0IEI7bl5nvoUw8xo4Gl0s3j8smFPDjfdPVAB6gI0HzUXshKg1YOXgNZXyAeV
0IUlxSxsHqJE2YyBwvGBPCHe7qVOtHaQmbbvYO37TY9w16FXnYSCvLwSELpLxpgE
uQ2nzXQfADoFx+tbMPLGawy9z02BoTLG9ICfPvfnrOV8tB4bI5/gRDnPUwGfBmNf
EernEIcGjwJsy64sM8mR3fhQ8oO6GIu40A+1j+7WCYVa2JthcIPiT49rQb5jVmmc
xGPfDv9szGZw76agcyWHfdB4MTBRA6yGlHjSKgARFbR8WKbsTdvQBhStjfIo6iGd
nrzLN8aC0hMGSwzwhD6USuJayHEFjoJnu0zWS+OnVDwk/m3dGnXC2L4CyfBXNvgO
gnEBNhQxP+AGCt6CVckGIRdhQt9LYsEQ0ZdZAXstRTBN89Af4T/wY5ZR5/jo0zbF
V4FMw3Z7CH9BCCq5613UpJP9V5XZzKMjjgmFUoKKx4Mos6QF2OJ/6uC6wX0TIBLm
ciiUvU+zFsFsklijHnfaj8Mgr8zOEMp33yPJs9xMn86G8xb2If/O2ESl08aHt1MV
tTIMLOWEHxjsfECL7HEgNOsMXHSyU016kdIJMqym/em+M8fly0uALbRA3iCTc3Ez
0Y2x65QWflk/r8TBufd4OZmVPV2E4VGLWhRIhsUAEpAvIXMuntxfKNwYAiBQQcen
vr9IUwp3Vx/t/koTd2tkqN8/4c0Xonak9+jk5nY7pFSJ3A01JdxtrAWCj9GtxX4Q
gBmyPdvfbRqYEVayBk1hBKo2+H6Ij5PffwSnEustX5M3TS0kNpDgeK1lKLwz2UpW
yNK5DfmojRydPWwIvKjL3B4PsKJVRXAo3n3AQs+dbuQ5KH7ng8sEITURLwUQFDgJ
vkEr7fzsVT4G6lvXRdCgrMFpBp9Pa6ypOec1By0XE+ncxdLi+gOH6irGgUZrQ2A4
2p6m997TCIuTlHjdWdzQ/783P6vKIoA4q1SfUhSDNFVBqlYSj8qJ/jIiX1nP2YtL
PXxX32ci6lrOCRC/pMNoP4u4WiU3u2B9xL+AOCEG16IoQPh5b+NUbYx8qgeWcMB0
EcX56NC4XQToHiqxttU232d7h5517Y6oiWsxXK55W23zKbtRbYo6bAH8cL1SNXt+
woAhNKJy/+mjwY314I/tTt7KATvzos6PURsCbXNL+SMGX94Xy3uSlwh8nWEgkaQf
x6Wx1TxX37AsLvftE4k6aMUDgiyoqZNbViF7AjYfrRmggDh8vVKM8aU1bQtdzdvU
fFNf/up+ybF8eGePlBGwtMZX3iKHq/mop5tLAXq1SJRHpfaE9bdpclvp3kPVbec5
air8HkY2sl8ztnPIBhgdH6i9u6P7zNwwNogFIs/V5CPo5qblgz4mbSjZMfydC1oY
Y8cCOS28lcMKdC021QShv/mgmponV3RRw8gtogQbpmGnTBzZV+FL/EsKzWPFdJmi
Ody5O8US0ojO2Jl2cyI5HvaGjlrjuL6cN1izlrWwn/URgyKZmc9zBM8PnqzsClQc
M6otZwvTlIOqAXRqstSpXfKpmGGUXBXO2vkiEmZ0rKI/HxbreHbEHqRE/UmHQe4v
8XprHjoA9Vbjuo1e8yM03mAmfJBflRCniUKOHaxJaXxJWr+izlaWCy9w4I4RVyCx
Syi3+Elu9uJYZMb6DBhG/5LEUWgAuD2clIDKS5sKj82+M6ioW4gER7qaonprls0y
tH7rqb1CbaZ4UJp9UcbowxScb+HK030H/SCkz7+OQn4Z4DvSD/2JewK/ROSd9PYm
sNXWALpr8MH70dO03X/eLYjRbenoXxuBwYc04j599jpMINfnipHxgI18JQnykp9/
SmfWSXRWL1U5DNY5VphvSnVGOAy84ID6D5tXg1mAUPT4tfa+vuoXQdvmL8DBQ3wY
1G4Q0rfzYbwixZEcUnG15J6oxj3UwUdkYWJyOpqbDU1v051qxGurweVzC7sfMERh
+8JHI+A+k4lQKQLm+qjcZymv1gUL6bBChNM9cyk3FF/NhA4gUu/skC7H7oIobIrj
f2HUNEq6Snyy5NHmb6zvg0tFnAXLVJZ9YcjtPvyljI7TibbmYSMjdfawXTqQI9uM
Iwr+q/mrEzG1pCGZOUiXm7sEP197XLM/LgkSbV2KPR9cfVcIK8Na7HCiUPgAk1FN
8J6ZhH+YvA/kGj/jCocNNpCqKQUeidLkji/DY5VCukq66GUmHZzzccZunW9kMOH7
N1vuJk3IyT6ZPqK0/lcojJ2JCXFJ4dW2S4lj1azxm2Dqhiw1Ryh7sQHdqNdiV5+F
aJpulueIpQvFnpkvcxRDUMO8Ooj2Z/B23w0DvccmSO3pTcJ4uRfRI5S2wyD/YV5E
ShNpZsTK3LgdZdbT52bAFNOOOQULXHdtTV+b5KuBq5xSGL9dGSQetATSl27R05tX
Kztb2Zk6zE+T6p+FuKRW/mBTBUZDOHonDEWTKAmYVwRNcy4z5+jMgwDAYTcAvBX+
hwXWd3fDuG8lfLDChTyqjtrTlg1QA6nuJSjBOPASB+lcUIGMYEX7qJrv8/6kkCd0
FgVWLPrVnAdyOhowHM/0ueX5dDNkRXHI545eY5A67o4T70IqfWuauu9Ljk8YnQUs
GLPD4PzYvn03KK+K2wDqmeGdRmg9hcUmkfUCb2zNFiXUdG1/qfOr/S4CaBV7F0qj
KsmVkueAuBplmeP3sxm7h7NMd9yiHL0Rv/kJM2aYn0aBvNoyN53xPlVfX992DnwS
sBjSA/jzTM1nuc+RTFUtSFm1XrNjNl+30cCkiZ6CmwEFMNfxcCo3nFEHiFOhyM7K
Uv/5sFoIrbmZeWmx0HPBzRVHQaZcx4N6qBDl+VHQ5bF280fhenBrqi/TtuUQ5rZr
LKDE0ZHnOKNmxatTTJy/D2dcosCjMO0vX6pTdSO4hJmmH9fAiIky5HFIkIyhtptN
RjicMI2JfruWOuiLQ1GoxmXVL50gK/9FLhWvReeKIf7WOM0MHTT8L2+6cE44Px0R
y2SVSnqt0DDdMlSi1r1sK0Il38ZyMiGodthqVi8bMh58P0t3zWJswfIdy57wn/fE
xZAU8mVWlykVCO8t/b0YrT2NnAnHjROxsx08lj0BaicCKIJrtEOIbi+1iYS3cBdL
yC+4CYQRhIMICCWp9RoENaaVzyvKGlVdr3EMn/XOcpvxiwybwId+VxNAfaZ7DyJy
YOPX+9Zio3EAqEen/+TiIzR1v17ovzZ07Hxx1tYwHE3DOh7gaCy4jMwuFBulWEag
lQHUMZbkm0fZ28XNam+6wRjinAk7+EPC675fLqVb1MBTh96QFKmjY9j7LOzXYlZC
srG9zfOo/nhik63vfJNY3ni0HQqdpFgryXzjK3gtMIA2rfcjIM75kZACZyHZOttu
9knydNHNnNv0iXeheD93xdoUIrAiMtYZ2D7AWC4dg3vhqCgKIHO7I+qViDpOLs1B
ZUDZKk5oA2ZEaFX3pZSuD7rqjU27VmVahdfbTzk9Wo4z2e1Wl8CSyXEWE3TxFXZj
51wiswGUcEQLxK/4NGGaRgP6/c32LmytfMED/N+hKUHFIANIn7DzCMHQOworkJOd
6bKqYiPpSDcZV1N+mlse8LS4nynCWSFe4IqcFDNhScD4zjQ5aBm1Xu/YIyDfx8Ht
0MaTJnZdTLnJewX7ONYU2Em94NNhSu3Rw72W6qg/YlSQbZO3owCLoeW+zbzm9RXz
IOkR7+Q+Wq2nqIzcsRFDOHU3NkTzSCa3ddUgJeKTO+g5YZJbQx4BTHvqP8EuVIUb
phPqyZEn/vSeesqrcabcHz7x93Gl+ApkkdxCfwrQbVHV4GRS2nyJaZp2PnwszHC5
2SEgP8sUieM4dCbR+b6zjma0ItpyvB5ASnrx9fxKnQaOErtLNgknpSDCN2b0oBo2
360kBR+tmb2SPkH0XQydowvz2mk8KX9hvAnAPz7PPtkyD+OkO87hPTsfEt4/n2Rk
vqDqjFP6menWJRYN9KT7H1zMsyUa0eRO2iUj76n4aomyBvAYekIG0hJIOnhdWEW6
t7PSjFH3QB/5/5Q0RFWzX9V+I3AnIlcI0Ob114PdElzNTgerjrLZ8S8GYpqfwnNp
NR0+TJYxUYwVVxhVRGjMnbY1vuwydDzWX68pzeB5+lwz7q6QiKOf2cRYP25uW6Ps
FToaigYawwPXLmlKlZc9gj9J5lD0ufc/aNNL/+ZzbHJkXAS1+hPkA2RDUjxbfq0Q
4sPGya0aDiq/E88PrRr6j8+NO5irCcAunKIEbF5sKYTxxxvatbN3G4bHZLJlnWKg
Kv49oZIPv1AQa1sZmiKIOrDKPrWNf6dYAio9B1+l803jSDzDpVWZQrBbc++q3VWC
Ko/WqbGtvCtkHPnU0MomYmVpqYlezcx73g1Qsp1XRS74jJio7MAGDR97ODFdUILA
tyYu3y7eA2VLf5C4A6XKRZzgQPGbdnguiJ9ACTgRcv3SDRkZ8hnffI/mOFTUtZ2+
xyrBCdQPSb0QbWF/eKpombK6gV/3cREwkOFi9d4ofA9nyShLmRPTPWPYUaN2KTYw
7dMIJG/BE7r9qLvRUQdEheLKYtxK/mTf3jL3R3R8Tuy9S2cog1lfugn5yfNpGfd4
Awo1QreKneQEgsRMuTI99S08Kc2iy0rZTqGnhOKyhdtqd35xOrDPOsWAOcwQ76XN
y9WeQZJsdtyUzoK3rBIN2fBtZNnY+6oDWLysTPLYTTJMqE26391j4dlBhR2v0OPx
um5/QxcUHRlPUo9KBl6NR0jBqruahIKMBtGWvEvtJ99kZYSd+0VaD4ILb6dakBHW
Jim2ROUYaLJJCR8jUARtRQ9JTDjF6xtQIOhmP8+GElm9L2DzGWiLNBxCchxMFV1s
VQYlh6fa1kry6n4gwFXbWnUo71dUt2s1eFpbkKKSzGbupAJ6B0sHSCm7Xd/dEK1z
JRwJahoe1zSwRtEigrNgXI81Ru6N6UTzAl5NxgwCbEjVyLWQ2xMuxdMOJFLCjVMC
BkzUhQOsDbVcIuqstrt0vcvX9aHduztbZ3GB5ixPLmocojuerjFMkYHmqUXIO2VP
EQORkg2wPz5PrdbEGNS3U1ZSF99Xbk3UybZbuXW+oLd/3QqVVHK/aAJcgQSYJ8XC
fmy6mW7RJW4kREqacYiv0lE7QhAzi/IOQRBlAvrAfZ/qsC45TX+4IeW0l89EESVg
v45kiyW8zcnnX2qTUmBLeLrCwIEmx+04Fdh+Oht7+f9UA29iqO7BxTslb+jZbJs0
2rco+pEJ1Pb2sBZtoZrG5u82V3weCFE2uFNn+10YKfkaMk6u5P6JGqRqCnUlDYlf
9ufZLs4/XM4DnWuumm+Oxv314p7aDK2X2tWtPuCBTZ/O+VyDvxkI6+zLZxFsuqbA
nTQH65HoxGfEC8SlR6l9G57sU/qZyTD6Wpu1OZG5u1D5lKr/f7Qny/x4DBgaT2YR
OgmK4d+5IVu1S9CUYr8MwvU4VUsp+0O5RhVl2I6WRtgrglWIighNNmQsuN9id8a4
cjpSV4OdgDix+gyQrHRdHbBhaG4xOww9FZ7hWfMhUHaggDMtfyVmQ3K4zxzRZWM+
8lUFt2kr7oH9D0GbfFlDLLW7HGN3s4i4aenD+bn4JYWKYRUi7E4WB2oLzMGS2Gyv
V2xQQBghx1Lk4rXz5VxfVy//rsj46yhTx++A5/dDX1aAd2JidAli6z7hxp5IdiuW
pfR0OoLdG5Mn99iLcGOxmSYyBBFGpM1lOIUIAC1C+P0PT2gThtnayELPm6bvDOO3
oABwxqU+AiSTq4V09oXQm4Wn4FSF6Pzlz26TVhyG5higibKo8J9FeClLM5JxFbjc
4g5uzSr+VdVkUnx59ApbKYPjCXNWivvv4N8v7+7NeZvtfN6eUvZ9C46I6XbImDzt
V/M09d2NX7ZfyL1eApWC8VQcAloEGs8TQRrzbofO1SA65xr1hT4loX2BIueHGiKS
u2Y5+GHN6oMO4DzGFf1WEDf0kYgAfX/SLy+tGdHupb85/PBINxoCDXT5WL4AqxdW
WC8HTJlPDQ5Ll0oBJAiKTETefOUbsao3Kd4o5DawHwsgug/N8RKSCOh3Fy8ejDkT
4br3FNRMU5nQ2EHfGFovT0SKE760dFNO3NbeDeKT5lumcy816rJhDxHZV9UYvSS1
yanEbr/U7IIRzSpsvgYNh2Tz1GZvhFQjSKM4aX8oIWFRtdTuUuY4rWEJRnAq+mQF
plBbINohgoGfTBoNHAyqSziE5HcgzHoABjXi3QsUbt13a6BAA0FUCR78+XN8scI8
ilGk3xblZDYz4jpQssMitnVaykfWwsSzMao+FA/c6u3+LqTN7wXrwugN3w5pP+Wq
VRHOE7bgKjAIBDI+AJ6MQvYs0vVvo46Uz9/AxYHujBo9LUEzfA8KmNz/ywkMrEPA
/V5U0qC8tmwNFOqf1D4CUovdqAblh0mM2fYGydxp4ywVcrwENoF9EOne19gZVVgS
PZjOOxLeJwdRxYW8/LLK4VmA+VRDyJ5YU/hvGnvb+BXyyvrMZSF5bDVHTRfWPtfb
SKq2r5Q7egc87D+o36QUZ0llmGcPQnA6CbkSA/640X7nweJpkgS2pxraPlYBZDIK
6Sb9rgdfjhTfYctN/rRUnd13XGv690Y/3THRtwA9rTU07DGKADj7Uak5XgTypUmX
Hzwv3bedq8da4ZIb9Z0wT1qkLBMiCD+AF0MSw42vogTeRdN0Av+5b8sQAlU0lVwP
pk2+yU9k7kjrTWCr+L+gm7rhevpZCSktHqQw9C/UWex2+8JYUqIBlW8PE+5MnZBM
7yQNTTNTCl0vFIPnPd4RdPe3yDM20m40OhyHugJY2JCVg4r1OhAvJl6BS7oY9Q65
/qvgKRWo5T9bGQ9U+59dAd7JjC+ASXv75SUonEz6logYWRPcMblYhcyzu71lIP9R
X1NMFeYQctJjYU+EUilrPnuardrr2JtnVDG4nuuYdtxqio51xNLZ7dLnRK+eSW6a
FKZqvzJGRS2FK/5SgC3PSGiHWQEkROT0iqueK7vJTNhGt3sGqapVFsEamTSaQfIt
aC1a9Ch3U9UpEhq4y99zBtxP0C8vMD5fo5vIVjni9FBBcodgbMw5enss6DP9sHka
3chqStQ63/hPcZdHtH7ZU0lgSGTvxlvyTXRDwcdTtf4zjHeNtf45bGck1/mNRPmd
MTbp3h2BBbxcDJmmXAUTqI/oxYx6bgurHxF/nK4mwvIHADNSPdlyuUPdfdTg7PPy
PnMZRSQp9usVcGLWZyrJl8tFK0o8UD45v7JI/NhjHCY7khMu5/Co3JrEmHJGXCQ2
4OciS41N2HgzqwQYbAIp9gj9zWQQCoxLKqs2BRevnPDBg26OxWe2Ii+/yYI48N2n
iYHJbpzgisDYlx3z9q5Sxq2X6Sp8fr3UpRknd/DyIGOBvUmnzIWqq11kqlLVdWLj
bYJiMOAHk6wGSZee6B8V6KlSX4r3Ogt8ngzwqDOOZ9vnhd4O4QOTTO2LjpWO6i3p
mFxZ9+N8mmY2AYbpaFHaP8RpohhhKT5n+OFol7mrOjtbvICMyzFhEHvgfbj5SYWZ
PJv6Hn8HxI4viXzoZBpFfxX6Oqj/sX3zKVAUfSBy6ZsFwN4Y5SG3dNWavHsqpM0V
hzROt09Ju47PGzbeC3uvWtF6Ef8P7P30Og5LZU7ura1nzcM9zTjjRLYRvGrU7aOH
KY8REZ+PqS2XMT1+T2gYvE0t7RbLfwC789S0ob7J1FEVI4wOvWxvRBS306IE5z7F
FohwoLo9QNjP9FEr6I8wAI9G/x/Q5Z+R4qB9IoSzUFkbj0pCDVe0u+qhU4/63aM2
znS6yv9XBqZHRv/wkrMXmAbQBX7AXHwdRJYFnEBYzaL3jUt9UlPZqk0QLOeCtB30
Iv27wgzL4Vn4WmmI8yFtMQ8nr1mxjoRG6JcIrpZPMH9g+tkNBxl4y0j0ottnC9ld
8A7y5fpuRtgeC8hOfXBkaHT2fNND5p/+ewJ1U1vII5UbhkhA2XyXOsOs9JNP/0Kn
8Qwtkekl2hBSSc02XJgk7CWpVlsAKqgFNcqJKv5LWSPlBvRNmZ6nePxFlynpLXrO
+HCl2htYv7cJLhHxoUewmQ7Uyy/pjiWZOLq5u1EkOkxR4VPnIWJqyYyu+rNh6Zte
B+NLa1apF/p6J7x13CRWNd+kzNw+nOOa5hqwO9oNMJpFWztEqF1bykrKaCAityv7
pKn7m7i/V9dspchCPa6AqefN00t/ktn6sqfolYQSQgvH75bD2m/DwA4r/ZvDB7P5
9ahMUw5uncGktG5UzAx3DNG+Ie5jQvvRU6jVQIxZM2R1xyoq+jTCuFjw/PRi5mB+
C8urhdW5c+wtGRU56UAzduh5FmY8MUxqWYkk+ScQFZs/ytp+JjnQNsAeV6JMlvYX
vqX1ONOxm/x/VJlDoex2yvtQW67P7otF9HsHA+JDwIrfEi1CRin1rZ0gGynN0THf
xhbIx09BvrKhbhEAZERqENQ7FkBaozWKNDV7+lgqSMuPE+MvFzLuUt66k9YzX2qs
p9Jfpvuv5Gwd/yI0qON60tM48QctJ8ROiQ9HIgd28wf1K5HaMZy0/2Pt96k+1dee
mcFqPhDMzLu3Jt2jHWDyNgV83Zac0DyNotNvfj3sFfTR69scjWF3lXai3WAT07Vd
Ola8r18hxL0mn3VSWIU83+eVicqkVlJAJ0ZoOuDsoK3AKABh0AxGjv5eJCpS+Hdz
BSu19CqcX6DLz6vpHTTgGWyfcm6AsURPl4hcwa3Zvy2RB8I5/U8ibPXkhLWfrNlD
3HPgeqJviNLNExJPrUXKi9FGBVMDLSBPuA0GDR8MbB6Rr3k+eJkWrGkrDctxSlZd
U2FHpLk8gtImPZw/vQ6/qN6p1gwVBTNbXK7A8iWpK14KFnX1qN+1odBgyekhPntl
8FAw1Ly1IWkkkXu9gpXQlJAO+J4H8eU6+xknW6K06PTVM96CLHxbIobohsORExqQ
ESOHNqlgZsUows6/3wX8bZL2vEnkP2n3XU8vpBMI28BTBSKHmR9gqiRVbi1CNuxK
CpNqixyEG96g2mH0z2NPu56+tIno/zY9AxhJv0FygBm6sS8Hqfhjq2UEXozVntMz
CtgyIK88xToKyEdiuKmhbpBtVGC6pv/bgLt5kYKlwTrwusFEX2x1yVMls2gKjes2
7IWqTdhe89UFNbclwQdKpmaatnJ/+JcnbhGQzdDjNAIL6swzJHcvbipIZrVqcISV
8KdNKlKbggN9GdBmTMfXgNVb08XuCFvWBJpbNHoGqwjpryl0x5nfOEkqSwXTlJiB
k+b+2gF9RbgxYQV9I7KYYstDdcBPbDduMLi3Ea/OyiP7JlTG/6hmguP9CvCtv2zH
/7SHvNgDHFEhHNzGFuZ8GtM2p5BRBi5wG2A2qGdX7CsmCcAcyb1nH3Fe3Nps+1TH
2H5AajVdiyN8qviL+dxscc4jCgPW2rSZOCtZFd3DQCX6lvJSxbLANohqHE7uNgdu
dKhAWWw/pCtUrQ3UoNm85qlCdhiRKqsz6biWNaUwqAINIDMj38XiU52WjM32i5Qj
iJcQt7tYxgHdG18w6yWhRS63jGk/LTjA7+e/fwVOwbaBW1+PXKxcWWEbEP9pS5h/
5m+WaC5yRzYGoLMmE5qCN+qGZBovx0ug3j+tiprDQxuGedBDGbc62j07pRmIta4Y
UL3s8XpqU50zMK84E+ZB21U2RON5gHwDGenOaomfXvvFUZ61SElwT9DpGAg14gpw
VgTmI+MYoPij54+eb0FyvkkvfmUqRbzCSDvkPDquP43uiCV4CqYNs/afEXcWPnmx
0cGyy8VtjtBB7YXoE9cbvFvgO4RjPy+M0EEV/W6Y452nartkTzI5zfX3Vxu1+h3o
8s1xa1yBcICD0l2yVksmo7tqta+HaAJz8BGov1KmYJJ1Ftb+8N4MUFdGX/rgLLk5
9LDwKeBZPKVEHVC44yUVxTRYN6ahHV6HLaCdYrRQp6Kwm2VsQqJMHGHNq1zNMTMZ
eg52Ci7ktyFYlXPdDk7hhCZlMGPwtovcYNcbgY0XEEKxpviUrLFrcZbtqqYwDgwI
HqUI20BbsFu10LtxqH9982zxyDTwBEdOMwZnhdxLHlXqhOL73tcXpa7qk23Al7Q4
sLyGt0szRv9qPLUI/cSzt8bXrWuQC4fF9UVUD76n3RSL4XCUJyO8JfUvcIz2KClh
nzSleUiLQd3lQxK1gY2i+SKstfkDU3vhcezxSwhGJUmhNlSFbFkuJ45eTyQB7xNS
XkYDlvbFVKGUuyjDRLiPKN+DNIelw8rzEB5xcxc5s5C/3j1cstI2uF6/3zqaookY
QgZl+w06AD50KfgfjOy5DvLlSAuUYXBFUHYiuTbv7KG3x1yxIz2H57S8G/usCJ68
UNAxQ/bhWQMOCoau5PIa59Ux1E/l22FbMjLxpjpgmOuMxBSx0dVip/zqfL+qFBBM
zUKvu9aoLofHO1RkPld4+VwUR9ertSpMSN1cW+cAEoaqK8fXNA0PIZeZ+Uq0YTEo
Lls/nQdbCFoTUCN9kJy6oodoy2bMIeZpbWr3CV1QPkSkr4tUhd5gYyhADbjKuMPZ
+pxtyrDgJlOU4rtO5X3mZeLTMu4nwF1rKybgZiDSfMSEMnzMWQ3gY6HP0/oTDYOe
0MvCoOQTBBNIoAmA9EWbwkfGxAtrAlWleqxdSZXgPSqJ56N78RuahQG70qFODmoT
E7SxMz2CFG4owy8xwRPKLKdSTmnq3B6js/XhwLLU/uNKG9Jcpbd2MWDBofeWMkfV
BxLgmKhyujoA6X8O6mqP3zp6gnRYKN9Sh5/sL4MxIBYAUxKuI4Z4zOu5G0gFTG+Y
N69IZTO//ldak4hMUpeV4FMRmBkHK6LF+OuCa4IlxDSqjb3jsXFS4IeiYr+te6KH
QLhy4ym1Xcu9TZK0r5SZR4HiKNF+tEIv8QYyAXs0/nreB799X1wgh4PFGuZ4UPrp
P34rtOBe06o3vxMrOkn9RmRvpP9nrGJvK5I8a4guWuzj8uHsWIUCphHgynnzJQP/
6Gf6Ti+IePBfX2O87AtF0jOkhC12kI9D/UfehiESmE+c4HOkvHQCI7RvO0zMFrVN
5ue923m0T//r0VxuRpPKPZElwx59F2kvJGZ+LWaFysyUoiYc4cH30f/uEg8eVge/
pq+GHwlDUbX5PVq2g2iWp4QPZteJOfO1QNJaz7lDM6CTG1c/RFTqArBgrJNcRnu6
IEnX+lEvew0kwar+kM6Aeu5NzWMqn+zu3imlTQYdaS5+GOuMG9bRPR4fbRtcZE+q
owBRGfQ9/HhaCporTVwfnD4xK4VcQ0cyWJ0rytBRps6yDzIXrCxMU2AP83uhuToY
j7xbTv3bvO+RaCLYwaBhUJCoAgPs14P/uo1WvNR9vrfo1cHVNGJhXTdmKJYyepPm
d9opq5zzWtHs1snGPCp4SgzMGrSBCvOvJWwrEs7Z/DxwSLiF4fq7G8Nofe9F+64C
Ze9G1akXs3y5ughGPpESfjwHSdEJtUsnrfWn1y8WoLOoTyE0sNg168cxKD4xsySx
fo8WszR4Hmnt5Bsw5QDl+kxvrgfvnmbWAU1Ab+nZt2I9uqVOgFE5TX8xXITreeB9
MTotuyHqypmgHt3aSvnWI2Iuad9fcG5gtp+cCqmNBEMP1h/FKdCkkziVXkH/uQ0l
aKq0BhmMU1s+xXQzpvTNYqk2x2mvCoMxF3BxE8USuV9a15AGOsowkc4rfWN69Zwc
iOQHPSuIVS2MrSWlHFJMeowjqQZBtTwgXiEAn8oJ4D1cNQYnXZ2K0CA9KpArbP6z
+aKIIulZ1a2X6ABkIWSv7/8LJ2QVPgVNu+HlY5asv6GYJoN/KQ6RTUH4oXs+0RhM
pfMltwEkSX+onEBwEAEAuEuAUAuhruNy1A0hT+fzt2TARxorC1QjGIC02+6+Dcfr
4FJgoBZlXB4NcrbdxM/8esZCWAW7EakscTCd+ewbWYHVLoGZi//XBVkR51PTSymk
6HyonNZKGCTr55iZrAb//jXihcLrUfstXIcQxuYOXQ0jJ4N3adeM9QM5HKriix4v
mev8ql8eo0Ed15+dGWvnJpvJ9a+TO6eofKstW6GBt22TLKLXMOksPbg9ZPuWRc4a
TqFKg4JFR3Q2Zs0cBP2PDZPGMgpNzKHLmN/1/GqAPE6MeLIXuF7eVSV1O49fkWSg
89IZI6kEN//po6eKxjPOL8JFBs2HvAKyjxEMQM2yQ0sjskgr6YmdLU9GbnAePBb6
XWdQcwCyDhohLUvtCTLrIdYJr09Bp1VYlf1lRMqCLqXJPcM5VFLu5JQKjsAYMDh0
KONLTMiEtQ3HSY0D4Py2BHcQFX05QcLl3yzmKk4jpWNjzerFCC/9nTwmL6xUIahW
m7lH6rYU16HvOhJI4pcjXy38MnIpRaWGPVDmismVvTHD35v6Nm0krESba2YwdYEo
JcCfLEPAl57ZFN0ngpnh4xuO1kgX9htWxSczAkqchhF1tibyMw8kFgoS7lz5EUZg
m3orKTyMVpj9blqMx2bQBI67EBF6THD7m2uR5ZTMr2aG1/o0cG7FpjGEjc/lMe23
IXEF8pLOJYvISLq0DL2Qc7sJ4cm6nRioAaxjaVUtpiJZjHC9aX2KdSYF19xnLpdw
Ppv0d+ij2dl8QLKkz9nk+93mFY0Lu39p970+t0HA7LUkfOZIYyMPnnRBavzUw1CK
rjqLJrjsQiF9izemkMRK8inmKx/nOlGHebTTlmbn6FKOa0bBkP4IteKEP/38Yd+4
LxoKvBHwUtue+5NpzKo7N7z1FtS7aiESM2dxiqykimqlczXzXEx/QAAZ7zQ5MJO2
ix9Ur+Q5HHGjG8sLXgMAB9RhqF6UU2sMxLnLH6IqB1xnca6+l5U97O60JIzjtCk6
LFQIomv/m0rYcBy5zEUf3j12ZsBZ+MX99WZl1+dPm5sUDT6Sr1luu42tDsmwOHly
r36AQ2WkpeQOumAbN4hmZxc1hPmUrYP2sHtWI9Hpaayx4+ZtNCi8fTBLyQbFNkTb
4nWoFt5JCo0hfaCw73VUrdnpHOntIQ/PUpIR1Xg4PsySv5K4jc/fnZymlMrzQOEb
4ZZkdb/SmBSevC+flupuugCoy+OOhebHXFrX0K8EiiG6uwgkf3l7vpJ4eoM3MJzn
ubZoeBjUwoMehhpdIanivNH71yC9pwcxuBnhiYyUlznAnMCUKQ8BMgweZDs3tVox
DUpgLFc6+rCwomUbIqzm5U1vP3QzijUrSYBFRymip/FfZzb6s8ntSCxvozj8xa+x
7bGzHKwn/JpCHsRblVtKwBh+FSeE9Tu78oBzt8+BcffDCciMTqi9W/fRxa29/Py2
GRCTcVtYD4VzDwDy31vKytirwRg+geBFcP6bfj4KHwxMBaN0lNOY0ubNbbUDvo6+
ffBeXNAgPmR2BGF8VnAnnltT4PBeYcv5Xhe8Q/kRT1Ws0WqBIawIBKPPQFVytc0c
lG+UkdupQnCE0Ib90GtW5Rz/YKkRJ7lG3REZVKSePG3IOF55Apfd/i7VudadBl3U
MDbBme/vVmaPmbPhDEMQq9sjV5yWx8Qb2C56bU9+TOSmhqSBE126qN6w3y3D5S/G
AsYLYyyvzEMap90SuCJMIwY1R3g/FgRBytaIaWSTIQebWRDBIVflgjzrlx6V/1Lb
EkHY22m0CZA52bOVjbvh7PHCB/eOSqou5xRttsaGee/Kp/qs/qYBN8+OsVk7fHVf
6LNLovqBCRf0TR4/lp0BBQPtp8/Fod1Qpc1aunkQ50oTJH+aEPgYtb5zuenLAoEu
KCh6i4QBIDVvsk8Lislazg66wsiecQ2ICvnBolunjr5SCa1GyBwfw05kr+Art4bQ
2ePZ5As7w6xKN7tv7R8zslEnT/IpbFVKgizNd8AI5BvL+9x2tdH4TXKXyRgX533u
NC299dYHblI/8bFsArzTcSIFn7HFMZ1dt73sdiDZ71gEALyLypodsMmHre1fIyPu
WI10j53fPpezBDUGaGW4JUYkctooO5Oz8RtSAak5zyKh7G6BB4pt9Z2sJwzJxO7Q
E92VJ45ME9R1TC6Bg2fApgw2zWPrA1C44A3peU2En4TLGbvYzy5lwICgKpE2yxl9
Hw58F41+okn4aRQ+gqsIClxN+QEWbVDWNB3fUhTBYMnPlJAjuaxBYTT9f8PnccXn
E2uaoOCVw3doRUwQcqVK4pmlc3DVigYp6AfTxoQiGtXvNqDv+Id2NPuXGa7IvD7E
mSDScG44bL3e8xa7bmeU2m6OwoW1WyKT7y7pYIJggneY0L0jp3Jy1e8hO4U4mXKx
bAZFRX795PepvEM8jJgeluqrqlyL4JJijOJPqnN06DG4mxshmoaDTwMirFDJzaVG
RXr3fVmGSK6gG5WhuftPoYtsKhCcmPpESz7D9+gJ3cDKRtwmHiv4LrvbxMBKsG79
REBzxs4locLbihuhH/+Yqh85gOnxp6f9nH7dTY6Vj3IleL+wi2MF0ld5+4lnIrOY
Tfitedf8t5v4HGVQ8T8c3bvfWPTGhJnTkGlJMCCrlK+kgz5W4ehIwpdKUZ7vCPxy
JBFzDkb+d0wdAxg8yM6+JjvROjTt7X1I1+vl2bsRBkvmfRgQRVbD/2c+RwKkloOD
2mcoRuRSNn7lnDChnYINns7PoOR6em7sKp4uJHcbMS7N4Tg5nNOLSKD4LUHQ+1As
cUG4FD0kLGEqRZF8PK7ReL8WjVSr+s7BSpJaHcfPwfYItZBbDhIQkZFrJRx+RUVV
cqo0ceFAnAtVpc9N11NbiKEyVWx8uR1a46P95+4F/72zJTmJyG5qABy54YMD8NKH
6zrWDbk5QU13unPrwdbUonJGFaKi/u/N1rgcjS7mtGzJ1XrxR1UvxWj+l/LVvQwl
to6pPh42ZIWwsZdh7V409YLdA93h94exknTIrm2safWQ/guFTmoXx4BM4ikc7EWA
Hd7sANNByPJoZtvDokaTfySJSWVajnZTWsR8tDFIORju5gv5do0NG6Q/lzqVvK5Q
VsXqtND4jZDpe6J1q99y6vzV34TYeHWCjFQYNcz4M9/VDSO9LZYE9E5mEm0B/lhh
HL1QOYWgsAhKpDGYoMV6aGPhrmBV54F91VptdqWzntpv1MrYIj2WPz+H9sYzNZD7
yodLZAjh0CFUU5lIUqlFMY/igIR+goqYrPU04LA835E25Jp2VgatKnAH93zHbSVP
qr4uosy2ed9TJwG17uBuNK4IQ7cVcEKDd9zsg96thiET4NVymsKEakBq9+Q1TRYO
HitRcEikWyP2VYpaDYIQAgfK2zr+G9wZBwSV0/xXhzZEC+AF5QsL7qXd/H0dMxp7
sPFrrEP3QrFScdZlnWHkMdBTAdDWOdDm2oIWDFueva5QtMt0kfPZA7lcSqsHck2f
7+nXy08vdmTZuNWwlJXXQ7+Lvp8RqWw/UQq1H2TlmAmMrcJkJDoLXYkIOb/IQ/Sd
Rk0VC9TUy8PebKXzbrPWsj08taVSiwmGFqEf1JkI9z9W0ljeoAEVepwXLTSM09Ef
fh1QLO0TBsgAc+79YXYL8aSkMstILY61v5xXd+MpRXKVabtj/23usXWBGKFpDoM1
PKodprDAxz4rvgDrjzzfGHei90it+Sc1LtRbzKk5rGbJ5ner7ixPstgrLm1uDiyx
CEUkIBzo8EPL9DNzCgSlVPI0qpovNOCnTSIEETqMdz2+nlgqxupZ4JDeITuMnVmD
ybLwdtb6ZGBXNPZtRv0aIVOoO8zq/HoM+5XELJPNlyeJq55yBU6Qit660INqclWv
iLJQXguZ/xj4qti+QSosA6CHG92HFxpw6ikj5bUdQybuzGSvx1x44/YbD+yvezn7
e+yEyx0+WNn39qWAU/tdruGcKIfwIXbOpt56x85OSmKUqWKY8tNRD1sO5n77/ynE
VwfbexhGkjGR2XDqEd7BTvmBhcjURJdPqO3OqHdypPkVeNMPoCnGLlGZz+P2rqmH
ieFlThyRFvQSASW6f/d9QgV1tRphBLQId6kp/AfeV/4ziejeaA9dLXaxt2m+NzjR
yk2tR0mO6Dq/1oWAEDlua/N6Hjk/Ch6rKodwcbXeAdniAYeUCn8YNY0FSbB0Wrdo
GMxogCRAPwuoUOwLZdTo3QfKVXpdnizv8Eu2G/Z1uebPYJCSand+aKDT7EpzkRfD
0wHeNmllkKhOYtWBzc3DDOPydmZGcpsJdS6vfgbha5ppr0R+5sMtnBs66MTm+ZIw
XgwuHmgQSwfvd6R15VJ5JyNpyBrsMSnWx77No7121dZXopPRwg3X+RzgQbcKyqms
LJ6XJjxpqBSr0zuUi5U1In19AfORUlV3hbr1L/KHtx47EVKuwt9er3/ktBgK2MhP
49YkPwFFmnFuvw9YXMuzwkpoTAw5fF5+kvegr8b5mC1HaJm5BslA4B6w7z3U0O8c
z+O1CXRbuv5fIybLbhE4oK4TOj83x0b7YJwC4vd89g/AvpqG6Ke+sXtqGsSb7Ac1
+YJlkor6kNLAAs8oLawmtklmhuVEl63rB95mj7iMr4M9d0NFEN/1Aj0iiAK3xfUc
BgyCXRY2g4RghVH/sWSEgFKHquv52rWrmsWY1NeUjLKkp9EMJAAJV24pLAoHPey9
pHWJBXSKYr1+mTLWvaxmhHtzLbGKQ1aKK2sm9qGHRQ7Lxh4KFVXcA7V8bcxtaFnt
GdSIUT09u7bquS6yUG3aISvq9Ul+3bL0lfc9N0+VaC2Cp5b/NILlY4DzoLh5coKF
uEPeuV+WMG8tpXgGaeNUesekYBun3jt9Mq+2n2Wqca2ABKUb6H/40cPjrVVJMZrM
mpuYBXzOAsX6TXzTIeUmmCMGjtjIUyJm5h+KhrmOskwPDOrDvWEB0eJ8SO11gaKx
4JXIQh17kH91IcG6bkVHNpISgQcM80wflXMLIt9fif17IgqOOGkQ0F7k5cAZJKLD
KSP78q7bT6tEt9tdd0z1AjUYddzohdij2NExdC15NgSpXIzJIJxsZHLLK7cHqrIB
4bCmy2BfHtKV1SLllWfsR3hNigY3s3Ph2+XpjJKhp3oKBilNFfxmm2MTGo08GwA1
BPKhxrXynWAzq0nayNFSTIgkhcYiOz3FaS6GvllfFdxeAykOdn6hUUkU6Am/e+q3
FMjORE2pM67UX83H1Mvgt6D9LxCi5EtZH0J3Z7xOU3EUfgrVq8nbTINF3J6tVY9s
l/aWBxrnzUS9+WSOjIpmfIIRWiDLSaMcgMB2gxsXuHAjK17M1MNY9egOZKgnxOgI
q7es3lo21ByDr/fscAmQuLPOvxYjLbQS9H/Jk0yRo80SEyOF8t2V8AnfpH1SPE1L
Dc0f+lXcni6Ttn7MRXyjQMUXDFBFQjbjrX3ibfA1R9w64ifHwcY2u8qbC7CKlGiF
k4EJd/d/S3U+6bHFUolPlMsJz0WWqNEd/uSCQIEqElQaD7YqpElqNEthCmY5skVr
xBPZUGhiz/WhGQPFqjgMtKkTvA6TqKvBx0GjqZdebOXsR0IupXgh3JimOtVotIUJ
Dpp03WSCDUjP5EDJ0VCFcZHRn4Fs8UWdCyvgX7iCTq2O90Kc2GAw/hcg+JNpXjMG
tUggk9XmAhBIv0juw1OBwt/pdYg8Ug/c/g38t4H2RQexPuFdx18ZxLnukAQHKEXa
zTkFqIYsyaDs5Mp92NghJVcUNZHNxV6/ntHwNLQajbEGWcl2v5X7qieSIpAekqks
bWqmmu08d/DknFTWKrSpyHRoJXpJIL8FaDvM6JBZJqioq1zaiaYBEBUpNpRkgURM
dge6ZkAOLGM/7TIKdZ1fyB6xxBv8KnCjFolSZOysc46o9Dni+gsGYWCk1cceA8xP
TaLrhjV1GQyuXoTIf22X97xPQ/bQ7uJrGMB2rMbzMyl0TnBHaYPNH95Y5XxgTsFe
pYy4YG9SqGjLzD9HFJXeJ0gASW9Fwg/vcCK2yOnEScRIAPEPyT2PXxmvkGLXOBvX
/9na2YQ3/Xmz7dhMLESOFWmz3SC1HCjmmDyfoYmiGvJoqvrGqNEZ7XDE/Ips8AdA
/2EsIQDTZffTHm1oKQIx837I9Kzydrj1O3F+6w8zHwoWvPcCGcfiWLyKRlzGItGT
nLm67gdFDvdSHV+krOh/l/DUPzrhJFHaeWC+PjBMXLkS3Y81CdjCWshLR+7h6/d5
K5UNpZrAOyv3bH1Wc8dJKwY19n3UFJQ3NFxGnyH4E2prM4ICUiCfUfOeEgWEoUzt
Z5pav28msMT6OUItTHR7RGRnvC03PNalnV4biqIfujvGmnJ27XJP6yotXFHASgI5
dpNA4cfrjSeCeyPMgV0O/3ZJwcPGZIc/q5EV1fPWD4tpxHmhR93avm4SSBvlX5zf
GqMnFshfgmdkYNdmkgrjfP7gJrmTHhCQnuybMhSzAx1ZBwxMm6IHPTKNLKzeIvY2
/qnL3dIRmNufpqX7//efP0P4S8QT3rFtYn7EAX1jmzZCkzuxwIfNZ64rWMU/EQLj
+kbrilzaBn9ynVK/O2emnY0Va3X9c10WyEtopYvrieM5B7g97H1zLrbzlw6fb8dD
LUOqBjbmhm3Rel6m+PVYLSvSMr/fEXmV7VjJ4Zc+cP/r0cMb6vSiiSynNdtVE9NT
KrFlxnyThz7d0VARTj5B2YEcNAQGNywga0L5WoiD/zdJ7I2xIOUwQM1MUYTWqvmq
mgHlx4t7o5mO+dOZaBF+huDvqdbe2PhfNm2fvGbKCtc8sazYNbgu0b0np++eUL6r
C3x572PjQ0KT8gfx6BVb7XKtDUBDGpvABcmP78otNfhpnqSsKwf5dMwmdVxQvBhm
7wYpaQ8d1D7TH3ZKgGRckrQhvlDnyTPEXuUtplcsuwioOpgzFVthVbqhRnzm5aZY
IInEhetpnVlAt3G6i4fzjQbX0HwCBB8EF6fO9S1fb2/zeAPeNO0eifjOz9wo/mdK
jHXdw0z2XRXqmIeztKwr1OirNnrFz8x6ACvRdpThOD13rZE7yovW4wJ7p5fMZ+m7
Pan0PkgF792ZtulCalyH0vgZylfx6khpCapi7Git1a8zaIrmlhUHdtNhZY0oQJR+
AaV1Qk5MXacF2V6Bhs6U9p9hIHVKpBE7slcb99+dmxXVsuU0lthdRBtY1PDMiQMD
HNvLgc2EAuawdgoyrgDkpj9g5LQ2pQytYIBuvsiEmzWCy2XNF4nmfO+EV1SDfWn1
1eNWJ7F1x0d9DkQCYgqWemW7ZyF86uqVnfEGtVeFrCLoH0cefIno1bq8CGjeWorG
SjXxuz6+NvpQXTrdowZHyvaNY6ei7/7jeV5ueZ8PZfWjZcEWvkEOTBTUvQGr2H1Y
b6hj10BwGSC2Nzl81aEcFPk/ybuSKs8A19o5xWTXbFClVBCc5dyWPoGyNQOk708A
66qPqvnwzGI4/Lednu7jfS/+I/fGVDmlLDHnEbG2ZRLs+ea8TnFc75pP7v+bb/ka
BxbdvNUZoh2Lywcrwosyt/xE1rN2uXqk8w7S/aN4iOq9xGJrOIhZpvAQ6pEL3cYx
LAko5OPJ+o3Yl9zv1KoxW0toZVjSakLTFgTMpJ1qfEkRjwRLb/4pju5TyUwYcySQ
jElTZXjeuBai++6mEe14kH+pXMxiyw29hJzzzG2GoBB3TE+O/Kgv89/CdntVApAg
u+4HZEs9lSvEyZ3t5modY0g56qXKM0bjBqrk7GspPtxaTQG+wqjZAxHdhjop/Hkh
1cCcu5d74JJcI8ClGuxzCqPVeMtuhVohvNpnX0iGYtDqIxW8CGecf+KVzlOeBCd8
uVMJ4JJrr83IvLKHUf+QnYhJWfmlRtLr1zdr89FMD8NcDsBKen8QO0ffm/qpA0TA
wY+zt4p2D/ZO+YRaPLPG8m931JWPRcxWCtMmZxytz9UY+vRK9oyWej/btCnUaqV9
Xr5JooTb2JfI0spl8z5hKPip8YE51nSOD3Zy+wFUiqpBx1mcNb2zEwoJcbIhqTMO
aF4SXETaLCrNQkUIIwqfIU5zFJNaU20xqfWq/7yieh7PNhL2yfflMZD2IGgtvMu9
xpuFBbXC6XKce3gTjV2dM94kXSZr/FsIeHnx5VREl6ZAMSRjwLwjZ9HMbIa4eaAr
kHD3jThYE/62+o4IGfxGdnSPvx8q9UkNsEMR3OBSB11KIQRSG4MBFhfCOkW1aisc
DvDBKQjgo1dK+jF3Ot1iqFBHDeDUsHefENRYAPSjyMm11H99sSKXkplpMIW2W/pb
kr9v6fx6J2yg1xCt7W9hc9hYN/NPtsKm0/d2Ai3+Fhp5ECUBYgnPtRibpuR4PoUk
hqnrJKK8GXb6SwT7MHSdhT6P3PKIejU0pdPBnEzcMEQq3DufMuy+YxoFHjWNbjr8
0AdL7RY3pqQBYjnqhstSt2tAvC6f+Pz+MDon2SLcBfnj+f0xXOmJv0Xl3U7NmJAc
J9sSejhVoS5pv7lt+2FSsJsEzYjthCpUNqAoPUZ7oGC23B+VbAAGnlPdJYsaVzOQ
4J3tsxsVpQurASZEJsJwp8qPl1YmT2UICvZIccPWnDH57cdqruOERlogGu9dYQ84
nohCCJQwh4Ygj1IlLKwW6kciOftMo6c7ZNtzaW1csQP7qnI0cXhIwZYtzSS2EV1z
Cdsf7EuZ71ZMfWDPu4q+yo/CA2r1w1xKnt1etxwmUX/Vm99/vMrRjpaYNnG41c9E
yq2cXTjCvzrO/ZCvfEatBeVFYPYjnvHmwsKLcaxOigv03T+PMuO57mhqgHEcB/li
jR99evVjPesMs8f+DIK5gYaHoEszkvWXYkjvLRfdKDdbJ5JhpAp7zA3LPWypBlk9
HzpNrbvNFOdg0kavCzP5YFJVjuhIixW4JVJDmBPG1YV/K8yIM3GJk/2de6YNYBpu
X0SrQ1vNk0sAGxBY953UheW88ljvyTtC43fHrZuyaBML3mkyY7Riv/xLJCE/aijR
b5rE38WPCBJaGzShWi69jobZB1g+wujzABmHJZNuoqOHh4QEjjPoPRNoHSQAQ7md
uqONIK4GC3CpIwivNB+Tg4D9RGg50/AiYI+KasZwHMuX5Qz+MzbS+XBxbf4thMUr
Q6c+xsHR9AQiZLAbAogH+Y6Bx9hleK843psv590pLuorLi35nlddpR2KiPlBCl9q
7yU9xVnAkggxuD1CNS/R0K59M+lAdr1TR5k9oC62odDKHVTvLU+0v9m+86672Y3i
41xdD9r7dCi6PexpAPci6+E+/rjBYqbCBWQVMMOdfJ/DeeytMWeMvEuxEDvch1rc
23cWd3H6uz+Mxn4ftHBIpJrAloF510hCvDO8XliJKqBAfQW9ObPMBgvlvUonZ0Jj
2BYEYkasfkRvkrSimtHp0Mod2WEihzRS4O3QHkvkYBGFGjp7PogVEP81GPF7XJdj
MzeLqnM1dqrTMLNnw+nMS2GXgiy6MpkoaO17+ERPhqMyrUwROmwD7ITTbdG7VIog
Cfc1I48FrSrljXk54dNCliXfE4t1v090a7628kxqnff8Cjmp3J1fQQfTzLF6Vw5l
/78a2wQkhZz1PZ6QYSU9+d37ryZ9B0n/J8WhhM96Jo3T3sdUa8To6kefw+s+5m8k
CW9EuvUzkXG3PM1loPLUTYADamZJoA6PACCt8eSa0sPUT3pB9lUPxJ5Dlywh1gDw
9TsxdfEK/sCxjOgg3j7R+g+PKLTE5sBJOKxEkfX0WsddJafpysG1a8tXz0CDUvRx
pG0Ejn2NsvUUtX8LhLqCTArAvlSU/tJpep17JDzoH9bVJ3ROU3++EwKEuY4Gr5hO
2kZ883UMJU4Lw2XkylYMKjLVyjvNeOvjMFMC23/FFUsWm/Y9AXMOnskDfL51O16R
XYjBIANBkxaZXC1siWIEPXaIERBjDszXiWVM1jJTyXjkYiIy1Lqkui41lP7Mhuq9
ilGPVnEFTTBPAFSWFoFe1cA+LZFRvouq1e7PaJNrNq612+LK8Zy/c6NAoV0kD566
0lqELVFFUWDY0aoO0zMkQY1jNqOAT0cfbRwnf1Q1MX9Fwben3QGrcKSGByLAEcod
MRjRojJ+zMjAwVGOhE4exyYxOru2gMa0+AQyrnIQvM8OppXg1O8BKOlRNPE5GHrb
SXI7uZ7spFgk0sdDOZ+gJ87S+XIzEg/S9UOUS4Ivbs9ranCa1yBFY2Mlw6+QFT4F
RinDPKUUrfRvKz+ONrgbDhO1Yaopl9WUQI7WW/fd9ncb+HgRY6b+xtDBwEb4RKiU
ntzWxSY396D6sPvnTL4n8c5JDeugBkcPnwZLTEk19uz77sTHL1HRfY78x8E4L9uf
O22ls1MJVTNJVsNSqAXO8TWEnZK8PLnCONV6OXvjMrbh69WqherqudbhoDCkK1e9
jyp0gGEsuWsk0u74hNZaEpakJTaZbWHqLS6KgB6NxvSjiK479tnDOGvqWQgFrgLz
XGQSBlDguYKuUjyMF62dYSnbB7Dj6iuUwMQKqWSzwC/B10mP+xZ86Ydy8ysjbHAA
0EPdwNdRF3EhPU1mOSmQ06gsD9iMqfXhLyLhHRbdEFXe3fxgxFz57KxAiiC3Nyh3
9ZAfMBWhtKHx8HI10+BCXUu6Q4AabtEuH4r2rAAm/5Wr6ytQUuEpeaQ18CnyJTou
UennJkRazwAHjbuJBKm4ha0hT2DD9tiQ2BYaNQ5B9wEVyC1NdqXqezYtS0u925zN
BYtIrdap/BjdIlCdSQ0ckYXyChXfBOFsKf9mxN8H1vpVJqnavxTCFI+kG6UDK1/F
5G2y5e9h+Z/qkr2Fg0ktzQbVHs3a/y2cIyoLJuC+7B8N5jREQ7XpMFdQXUn7Gqod
HY8WvrmfVLzgNrfHC71gni6NjQ9XJLbO+IpVojG0GOUZeWfyk5rOnj9GVZ42qnqx
23J/HqQ2JG30itfBNAG9MD55o8i421cAX/c6FhYDZrQ3VTRU6K7V7O6niKBp2IFF
nPM1bxsyAZm6mcUzP3aCmmGcvEfuYBBGx9T0oXW3DSDf6YeBSGydAVNn4sZQadaN
HAlLifk2RWcT7I/+bZfWhuYlU37rgxw0LcwDwHoxN6sPOr8d5JTmAm5e5YOIH3bj
JnhgVE8lNyXz1LQlnK5lh3Lby/SFIbhnjZb/lXwiZs2OQX7vQ5HzYzKZhizMn65L
5zT33TjKOG1eSiOmkhmw5nbwxjWHGOlKhDiX4Tzooo5qijtEOA7+y4k0O58g1FH1
8dhp+I0Pxtye1+8WqxnX5A9ejJ1uomAURQ+SqFKH3l3x9LNyGcyN2goeIfNNcj5i
/0Wd4KJarfVTaBOC6wKrCSz0PM8vm7Z7KXq1cm47nH6IELc2bhDLkWNvLNuODzV5
hdUiCvtYFnxWFJZI7YG1AQ0gul4W4njYSZ7PXCHRnxk1BlodCFKyglhXGUlTqFDa
x6AxEv6YzuB5dVOb5Xom45ERLE3BPx2XK6t16GfiCzouNPEMiYJs69TUU+J0+UWO
h0TxglV95DXWL0F48cuneaiOwsr+kMfZCBd/eGc7NIBp7/PVYILnEaNJBGv9MVeS
A6p+ug1kQdrwdYY0ZfPGpTZKmOAaoDsQfWQUnS9TM+58s3gv+hVhYcwOT8MzIfyS
EIG1ygc5QuL1LL5kGCs1va57zcpZdTAjMm6Jeo0et7wgseL1bm8Wik/oK2gk7sPL
A4dec3rR5gtFjlk7JYCisS26qj5XsULP4LBmBrdyVth2dm7tc+cWUln91yh+XLjm
v1Gb6JE91rDr6pbPgGTKRM9+fpXkw8jsJIf7Cqm77kiR7CZHnDgXF8ehaRi/vFiB
3jIRyhiQrR0ILD0F0wQsnb12FWNAYHnicnubLDio0ni5cHLKNbgL2Ni9zGNJPrz9
PUBrwTwg41Cy61WSL3Sotu9KxJCTfZO0K1TIFLY6CGtSNkMDJMY/94+9AmeXHbjq
UoucaNav6WF63q00kYFX9zl7WgCzk+YxxLqm6/sFrpp76hssTZqo51N9d9kxDAfG
8YDwFNk6pSVwlLhLwpqA7SSz8fEyw9Ef87uwWOWiRZG37EuuWPI0GyBjGp40OjUQ
EPYCMB76dErRHr0ryVs2gm8rXujA3L+HxRUKtKUFZFuqluaGryLKKnykvzMPhtUA
rgR+TOxSy0V9TG+FPvrnEaydIqlMrEA9w4fNl1pxIpzgLhsXkngCNkgMxui2nL5u
yb5QqmUhv13CmbP85M7N5jwjCX8KIPPuE26oAm+eiqZPdR+58LxtyYQwhCUYnQeN
w0zl4yAiT9aPGoWLnT+yQnr8cjx3IVEq2OPYB/mkDt37qV3noK8onSzlfjeEYYuT
RLhvcMME5vJrgFygw1GWVCOl2HIz0nd3OAgKqDs//O47K5RGFg73HIqSJn8MF1jc
kolkqiXe1MzRsRO3gfAMqwqSErvXTDnEA+XwsWLms96VQmfWMCbS4a16E6UzDA8I
toyKIWo8ph1iZ4XqRtEGm0D3sBwftRM2NHvYHX+v8bV5A7t6SgJ1Ri3byZSYQL2X
GE6cqiPaySeawxjk/Z7AYrjjBrY5xIexA145TBIB2SNamYy8+BRkicbctqiB6fmt
FLmeboMqtkltQ+0mkmmuEWHKsPP4vUhY9KHWA1f6feTrMOaNYA6boHs8qcD9lmuz
c3PyjkIL7ZweZIVY8zAk83e/7wxTE0z+5OQBlPyJ/UlTqjKb1J91zsw+F168GKqB
t6h7tR83fe+iPNjlA6axDdEYPpJmkbDF1OWBkd03JmHIRwBapt1BFSirPMctJFIN
KuSOVtTEsckI0LrM26/k+se4MWzSbbIN2d16YdpUY+z+qllw+0q78uiWoBEaFAp1
vVqBT3qPkgnykmxUZazzIfxl6SEGLLg8UjgZGQSInR19OTqkV2NcU8VW+KcqM8jc
C5pasmZhsgJd/MJ0Tq29SwoCBk59s4Im+DCYzwVekSvWgQU/I2c+jCbdR8ZsRmNj
SMfG+v6YUQoT2hHbYbSTTDPtePZKouZKj7+Up3ES7KTt3zA73A2y0W9JNQe1zp/T
hjtVXgtmJf16Ry2FH6ybIEnfU9hFElsedJ1bTJSwhzSVo4AZ+9FoHv75+tUh2KjG
4/1Tq6dUq2WOnCPhSXDmBkEpZ2pEXX7MphPAhQqrrrgogVJUfvJ3XKfg3ph59q28
3VJ0G4klmufiaA34Tt8eJXkGHEcQegRzXqT4LbiUBTRE9Ck5L1XX2y2iZpre4wCV
DkWWpuXzD67ghkWC6mgmkB8nwgLoUIEB65tldb4KjPaPajTmJoU3pvYsMiodr9D5
SrE9zi3mTqK47C3nhYCYQGvLlp+v65bP6wxqtggPKf6yPsTo+T532zch14SXXVAV
TzicKA5dSqYyVHlRVwwk8DfCwxMyTTlLSCIFS+kMgqWwlAxMOJKOVwes1KTO4S5T
uCZpVwKMHSNl+848Ij1vmJJqgjiL06ncezUEDvy3beusnE+s1ZM+NL7fVnEkzlio
850eyhvBY7YGY9KqIh2ilEZViKm6wm8O2rEy/J5cXMOXK76xCTChFlOlaRdwzyek
IeJ5S5g/0wjObV/pF6P0OhxIKxTeof4+7Q4dRD+hNV8bTPMz6rC7VP9PdfxSn1aR
lwNySL7JfoqE4s7PiboXPaZmR0USVikA/8WMSYkd78n/yWKy3IvV+LLA67Z2ts+n
1RrBmKwVTVlpttiHf/Pi3c/2pVH6kfTkBQdbF/HNP5I6XIubbWTBbZ0nBEuL+BiY
EvJLXU1sJqd/YEA4e367YbHbjoeDN2lz1AgS3iUKC/EsaDbctxYB2O4mECbNSC9g
dCxzOcoMw5ObbWv9Q7euQAFCtYnNosxUQIk36GKjZ36BIxoyA0L0vsGdypjQ+KTd
hDDhNMXwQvtq1LicjThAPyq57k8g/BhIiXtHgSAm9xN1L9qagSyIxL9pgsMmbOl9
Nbi0Tml6pNePD6XP+FBCpak6Q3ZayAj35TJC793N+6pUvkpNP9m0mjwPnD6kaO/z
Q7f1WBqbOyX65cIANW/KTCdk7uSYoM6TyLyLGfhjsOWMPY8sHNjnTz9knhhmUrCY
/+1kIVvcimT97+fr6xhxNrLn095SJvZ1q00rMChm96QsJpLeJh21hMcv4cjO5WQO
2SR8oFc7Kgt4KlV00BDd1mvaEs6UzrmEl+RkHaPDeEreMIfgD7Wc6CDz01Kv5xE2
1VEi4Bmx/ErS3IwCcBYSEPu4elGpOEaQ1+BCNdUa/DFfMVdGTwAVpMyoTc7C7bhy
NbVhvl0AQJTuyjVzmXXa9o2Cy9vTQjTvWnhZ8bFr0xKaYCx7RsYU2o7u+N1cM7H6
nncM4ijJyDuqvgi86oMcjI4YxB7GvQqnE75kMaP7vWr/FhRUzLW9asXX766nz1KD
IfeQeAiO4jJ2geFHtE7U3J7HLbHbk4C+JjSR3/m6hnoZW4qsAMQ97rw7h7EVsbrx
y0fZkN30c2nzfwDz0134SAhZ+Wg8YoVD88fs41PAeRUbCJDx6e0T/ODQYxe3Yrh0
mhb/vj4DjkAOTL2Qncr84TGxow3FrzvLuKb5+vUTJ86dB3nO2QJYufG5bUGn9jpV
GDCCxtdlmGCjxntYwJsc0ZjOp0Lz0FHZmadxgaLtF50j+6TkSM0PIQeC+s88kEyJ
gXQoyNpEqIRoYAcOARwAth9QP3VxbV9NEfn08B9eOyF25NTdoguzidvoxZ47Zsdf
mUmVUGNcGiyPrM6A6dxfPhEHmw29fS/xzmPfkkRAp+dIVBW/UhiOZx0qgodoEDdj
AD4ONRXifAs2qKi6NAjbtBsBQYf0eAlI2J+pfTGG8qR7sneQF04NUy90uJCMRjDt
8+ZslvtOghbe4WIsr9yleJEVPIMUs3PaWHmB2ml0XmQ7dP3UDjkqxf/MqBlDQKEI
2VL0VzYBNKduHSkItw2H/ib7DSPjxni/k4G4QiUGSi1HokWuKkQgiVZZIu3Be0Jc
cgJ8NVr2LyWLLuZvr4uU3CWzlHjprgztSTcWFaVuYVJAhsgghtTYAbvVpd4kyTMj
JnHsBp/+3aG9NJGYPl3toyulchUSP+Vw76n26Fkp/7Pj/ZAwTgdMmNmBxXe9uKuB
cNV8P4v8uhCkggPlHmk+7IuhJ8Gz6IGsiuIbVBZ6utIAHrwijtqgWRkWgQMn/0MK
16drggtpJYNol2/Kt/aNiR82uIneTkPlt9rwkZ0Yus7qtCe7SAWTtyLmLy2u0Nkv
1wBncrhkcg8mwN418qmqPG4cj0dfrMMeLwkb/Wm1kTIHt+YYOCYLUkCe4f1IT9zO
aEuqckebtzQcZiP/zsfg7VqqmTC9dBM29VCgrFTEBFX1W4ak3zoFMT/kjl+l4esN
dvVGhUCaTgbqa6swmOQdhp4qd8xkmXE+qsM9qsXf1Gfrll2T0Y3NxNaSYKLB9nup
6NKG75gdbIgzeqJKdgoSAX9McyoIPNha6Kc1Q94Wtw4HLXgUqlwuRYqj++LhRt6Q
5tJoEUxbtwPmspJPtS5jRB1/uRVA911SYlooxtqNBFBctEtQ69JLY1jOb8MRu37Y
TAq4hnJyW7ekbAKADawZWsIzfqJ7T9uNmSPKw+ZrNz7bGck0Z4RIiSUEoiVW3wY7
+5OMx+EnPCr6c5bMZtjZvKJtwavLhuFUGDlPBMy+JgZJ95b8o/H2s+RNkZMUzNoD
G7/1oYU3SoGmloXaXxaknE6K3v7xN09+3m9sGONsH4udlU80Wn+Bmjhr9u2O7zB9
u1wnwlJOc514aJpkdXQIn+vHtqTJUWPlsBweGNLAQWIqMHStpoFt8xTpeZZp8iMR
YqOcwY8ZZvQD7oShbaiqQmrbKMk/sfOt8k9QDIfDir5pYEefk6UFPDha1aNAs427
HNp5yIjX1+WaN5vX4/prRQZRkj9rj7Uf0DwJyq+1MfWdWcKDJsUeygWtaldkUR5A
1HiMZOwNPtTzzvFvWRcjXti49cwHqj7jAwvbbu+7qm0yEiabps5aumiXc8020CCt
NIvjcXArc5NhdOvHaA4kiNg1QGU0IHTL13k4hEh+4K8vilE+n+QbAZvasPWEaUDN
OnHKuqqeTiyYFIwZHILhZckjgpoxH265vXu9EQ3CJ18m63AFS9IJvwFQjFGu00TF
aa+xGjGFSxoIkkcc1WDqbDU4xY36erLdccUxzo7OXwx8sGWTcLOVGGhpYts12c6d
uKv/f+3LH21mDzpfnWSGQ0VkLJBZaA+jnQLDSH56fcPoY7VWhAoY9hgr5H3z6Tyl
1AY/PJeiMB42qo4FLePDQJzvgdMDWDsB9UlwQr6ycPnhNDmKB151kLwdViBcbIUr
7auYyIbvWGbx3TTQ9GzIfaKRbNEaST+1g3LLeOjuCnb+Aavil+j8j8MYe27mHw33
rs4+FTc1dGX5iU4k9pxS1IkBOCwSQ1QLiepBsiD9dZE4rT6XZW707P7YS4zFYiXk
7UtRopxDQW+adCUiPWFA7QHBJi6DEPqNoQEN0Ap5QHO6GKl64mUshC4nqFWci0ZW
h+0EQI4CIrGQ2bv+LXm6fJzASeNkMCPAkUnV6wfAhPjz1YpO2o7MLlBe67pvxCN9
0G78/FUzryz4TLfH21ARSWEklLa3MHBM5SYdEe+eaA+gYIBmfW1fkBw1vPqqJmcv
0/BcB97vlw+L9eSZhNXVyzZ4pyXQzbAE1iqHTOEdVFpfwndcbTfJv+arQJcl11va
bAHCvjAehLhzViGPsrE1ETBqkK8BKyrnkQrOBhRXodNDM/hnThA+bZfIzsEK6irs
E3kH5ub0IVuW446Lrbu1awbQiEXySFk/lMP7kX2K0l8cLIN3+wtMJpeuXw44dDoQ
Vh0m9yLdfNB+B8dG13xfJ+aE+QxBnUFVyZR+y64wXYUMA265yMMDGlNlOsgkM2cu
9wXFYYwtiQtaPqNMd1zpuVgNSfV3v4FO49MxToMxCZ8cf1yDJLtwCQKfGPlWmIVI
swiOVFMIX/zGWj8/1+cJDALO0l+hLb6D8dGOaNAwI/exPLCbrklOvQGiNlGtqW8F
Mbzm/bOIH+9Gdfj1NWBuZFecV4w3yUtChY/Ewe6kEsSPlx6b/4zkK0pV52TZjNSy
8HIb0xCdhuMIu4lJ000Fa8ZEV/2KJcDHdh7/TDItLAv0RJE1ewft0zPtLJBp9aL0
Q0A4xDHA30HqLn/ch1kcW2aQjpw3oKP1o/BP+tKcbndMfkrVgVQfMWwB11a4JuUl
M2dUtS2g//Nn4KEz47eklOdoN4fSxhjEGmeZwNyKeqz09ZK+ugjgJ82bfXfN5fq9
Ldo6x4CheA9jRzcgFUXzSV3jm1oalahAID8/RZMfFbfePBsF1YgSUwnXvYXxE/Ql
FGMiiU/Dem+hJ3kQfRWlQs8UWB0+Fh5JDUW2kD7N91H3Lkqc6kUEouxl0NlkqqtL
RN1ym7nBzXz//Nsk+EjtAqCtt4NRAdooz+XVU6Wh2fysAWcEhvWrMzRhIPK+lV+j
wzMGqiPtdCiXXIYFOt4EOEmOG5DsrXPiIMoI/53GedodzKf0t24JyDu3ju93IeNj
Fa7qA9/upiV3k1gskFwAAJCuB8r8QzD+4kj1cX38a93xRY80Qv+lUOIb9rL4IDEE
nCR7k4G1XDytKpVn7n91KUFETNHH9NRE16udZqzG5HAswIpKV6kNd537J24xdLB1
ylEJ3YCuVbdnL0qqcd9IoTCW5LgUJPXUd0SRnnidh2UWYWoI95O9HlPfDEkBrnjC
H/w0VpLIJoQEhUG2FwWTkq8c5JldUSi3EGRT4wq/fzjkMNk4av6sDw90I6iUX8Fp
nPAI52z03xBaSecyO54VAhlwlr4Wcm9FAApKiumc6JkbZioIAjIU1bErOPLYCCkb
vYfdC4ulZQicyYCe9/7dlV0Uoo+EhE5GhFmopIxdaCxsqp9XQlzxE/lnXqBen56F
+21QHQz+s8FLWBI5qr07zAR503lKPnhrFigwxZAc/PTQK8sW5J1bkmFlPcssZRAZ
07wp8ZJeWtsfstmP9uxacncWvRORvRGdk7dwmpWDhAlT0fUxHURgcvJIWKpbrVZz
gmpWHRUiknUZh2VAUTcRYNQFHg9y5H7VOhdGrQRCtFt9uTfi+WsmP1wDU2Mzbo+9
CKWbieqsLIpDBqESnjNGiWkHQn6V+tAZ15f5M9/fgZl6BZx1yQtZxDcOUOjNRtCB
UpACJ/v2XgyLJvQc3RHIKZqAjhzCWqSgKWfMPNOp2WNfVXMXu6tWRwYBZBRP5qCy
jEKZO2JmTjgZpK/2Sc+7x+V98gvF6p4up14Q6FJ4/fUwCuUmlZdeQqekrqpmzIwS
nHthEMd1KL8qDfsMnkMA3lkF6/OnWdZKTD8DRYo77uVZXHmVtQ7EDstWlM1WCaiU
VI8h1Lp5GP89Dh4SkCpwi6RIAVGbjvDT1zYMCJ2P1BucU+IWWCArdPmm8HfLA1U2
L2ZgXbDsWzj80T3vw/0ktTU+5NZPdDNirqZAA4yH1P9jzVdmgNWnvvjTF2tb+a5T
gy7Ms89CSDA7mCO+Jbd7i64R0Rp9cNOg0UnvTAm4DJkA4NW/Tsq3FBvwAj7zbu7G
mgwOJkZoazedpMikcT9Zt4uIoHfHD2zSxKTVqH98U+f8u0k3y8nhi0sJmCxy4pu4
BX+cfkaVFJC380l4pS9tt0klIKpBENBO0J91tz+JsJbGEbUsqeFoPkchsyO/lwuP
SO0bKswSsICPeAotfsHp7l4BW3BvSeIPGTloZ4YoZ9FQhFMskAUHYGialUUxTi48
HOm6wFkyrnbEQgd1aCCggjMchhB2YZL6uLwRIbNW/AoDREn78Ynf+sOieFx+VdRP
wU9MH819IwpZT71KrcpgcFcQimMBkxZ6L9bwpeUlKLymvBsRoStXQ7swK3CH02V0
kyteOSQKNeIJCk5LN4MNpOTOm4H+MTKWrJO7r1shl5wEW6i7pz+ifGlFg28e+d0Q
Q+RYDkGYDET9P8uJHMkKi1WFCznlhv7EINckP4VMO7FER79X6N4YToEZG/AbM8oe
SsYixoYZSc3HeMUN8Jt6HA8kECkJEpg8fTY+ssgYyBLZK8Ac1HVXY+CTTMARGhZu
DDJHeNcXoWtRI1dvmO6cbX6uPpRJ2C0UTkFygpGIW0U+voK3r/12iREjsnEmuUQt
kUboYeBJthx4tuFFPrzfsA+BR+2bCPJrorGM6OQXv42glNlqIiAUZyZLQpVCN1L4
g5WPEURgVQZNTSAz3x9RtfmP0au2sky0hqLBgvfuooDdvvAXi+3t262CrOBkcK9T
L8jP/Vqw+4cd4WwiBnnrqSyOwQy2lIbHjiPF8pIgeYRkn6nwbKxnZht2ZeJWESQT
eU11Lh421e+9sbvyFbyGEeQx2AbOttTH86/ow8GujcdlVSUP4nOv6cSco5vWVdKH
s0Rrublmd6FGML+LBWXHkfrZ99bJTJeg/VgEHmDhxV3Td4W5lOzGcHDLrJjcxjzd
Esxjq6A8iAKBKRlnPfFUF+b7AJSEWx07qYiWgzyFrgvbWVdFaX+1TkDEUY/vxYdt
f1VjaKWr0RhTRUCQR3Gx/9bRmRZ0HSaD4oM7Skm3BKC7oym4wmjX3N3IwyxU0GoH
9+BgORh1+DNN3eJfP9ELf4iuqisaYudtrvBA1SZ4Oik4RQ/Hb+XD20dXrnDJdJ3g
eBb4LczE4swSIiL5hKNoaKt2w4i13uPEWiBpoB7W+sv2Ty5Vm7a7diS8expJoSpx
5RgBfgiWEkbqqfWyA/PjHnNAHCIfqNy9lj1Pwpnak8UGfSPmhvyXkHKDS1tij0Ht
Jyy+XNVUfH/hIn9bK8uQWTxPrKaw6CdXZZJ63GsX0Dq2izrFsLU3B0HaQ7bRYlKq
vZovCOjKednnqkHMGcmA7n1xd6Fla6wRLUV35u0UymOqdLR4/hvTJDLZ8VtADIWj
gMu5HrAA52s46blDoB8yVszQKdRYFsLE0y9uRTf2rH2n9hd27G6MiOjvG2jv/hyU
hFoWdkyklnFV6YLnA+WbYD1gXxG6J+jmGQz8GmaqhYeZxbqkoxrUmk1G7aTOVeMU
g/G0nGtl7t7Muc754NF5hJteszTQSzn7c6wsFjd6yfqRAiGHhyukWUhQb9j6xDpE
YcIFcaINq6bjR5eXyRdndy25kBU3O6TbZLRpAjuRSxGDcHcoOklGCMB5EAjsRi71
jrk2Lcaq/8pLFskAQWGkAhad7XAZITbnujDPB4sBtLMj4A5fHjqle625h1GKCfvk
Mh2s58dG65gfmUyCMy0fBze/Ptp9kI3NGofZXNHNGaIbU7Wfwww33l0tSbz0PqQ4
jiF736tOBGClBhVvHIl73O6LkVPiA879O0Jt3gHX+66KB3RkOYr4GDIWjEQGNQod
bj4k65c9Y2pwRthPnUqi6XJxET68i5V/KkWNmDkG0lUAB1+wQZpo3RQTPXZrp+dm
PiP0CcGLmtpa3q28denccLazWKMyRBRwuniq2kW2AiiCATSESOdWGfGLGrbCsetn
0IhaJ0jAG8YJXyBs6HLFj7qNU0watLqgp7W78TYDrqruSsRJx/s8tBGIZJNnI4fG
hHhd9vT6NMisv217ZFJY88fDJVKSW7TfZZyznGLEmT2L24gbnW4i2P9GveKc+mrB
TJcbEGR+yOcA9LJGYtFjksVDFssboijScMwXMiVSxQg8yQhW5XWNWGVUiuLFdfid
c5spNbrVni7Xg/DUkLYV6eIvhqrIvya2fEeMnEodH8OWMJ9827emTK7rb3WYKHF5
QVsj/eEJP8wzo+qiVLj9TNssfIvQQlPv98PLofKRlvDwtVf5t05r8ZDjvAVClThn
WKN2c9nD4XM5HHxx6StF0L9xl8MZrx61EGINcSAVA0r6RioK6xC35luJVNEHSud3
ZBkoMm/4EP5d2tFx2Y2VjUhKOL94wznVkro+U4MxCHqwNOCSY0ZzvAJ6FhkYHr/E
/YO+fwX333q2kIqQmPVw8eeK4UnYtf9eeNsHHYPBvMlRyTFUjIv8BwCwtCqjksT6
r3lnsPaXY7LnPmKU3rHNjRnvkd1S6Qiuiv4bUwICapI70rgYCL3uXwPbtj/YwP/d
ntqlLw1EO55P2icvYxo7GvynZEXFal3QPLTtTjr6ajgMI+5KH3bfUL11eVjCo19s
4MBmrEzfC4DnTSkI1Ep/MKuTgl1Kn8DnB1a9KdI1kBRSU2zAIMrK9uc5MYHc0ROy
KizpgmTNGXSDPtRthGjxvdFeWlURjsF/lApf5+GN1n2zRd7x7dJJMqmXNV2cX48Z
3fbH4FXnoYTvDc98rkDofQZaVtI7Gr0o/OgVY0r9wHFxsTfGOmJMSnpylwqWSCy6
vITUo0VP7R61BLiIeyyHAG4aD205KVORzreCNXQz3feBPebDBH3ELd4zvIsynvRo
rPpO5QeEoUl2DHA/VdP6lRjQkuoaC9vKY0shyGOqo4Qm+Ld3MoERFPY74ZOrazPS
Ht7LgUeG/hDAL1FZVgP8tfHTIJ4SnohoPBrSaMwk+TnoqzvMB478UYkfjthHYCJ6
n4zWRgvNkNWX44T7gyAm+Jf2fEwSKkDwQVO+k9rkOXCcPKWyj7O6/fw02WjasMPL
N3ZbSVn6sSPkrTZq+/qf6tdlm13DZCuF1HbpSrYrfoX4tq3OAJcB4inRKd2C2cRO
hhs90m6jtyW69VqczDT4oxVwQGaqox+dZBK0dqcPZiFsOiYQNJoRceB2sXZ9IOYc
nfmlQTbLB0nSmm0zaYZjTC6rS3v9nQkDQ1OteF1aJbg2x+RhqY6xlDCuvH7xHaJo
eprZeOxpnBx2BKVptGf/tuzDyBE4Xzp8NmN5Y/eUwUgbiextjfrJ2EhvImV0M+3x
vJa8h1bGmbiCyrbcIjc4GCiFYQoyQb5Gk6003K5Snq7VlpeTk+1qKOmOutjzc9Ol
owMVLaE+0FkIfcSjM7fIUZrBsVADD16+PR8RfazCuJNNXf9b9TORS0zk6hxyrA+t
VGYPv0KV3FOkp12i4AWPzW4Z3wxorlEOg8qutixqjSmmnqC5ZQ47ISb0o+sbjKMv
QHcFhfAJlDbHxS803Ey1DunOmnk9p6WY0nmq/M/Kdv5WzHXq1vMIQ5Y3uBr9g/FU
2Vfc5NBkDhQi4NXDehD1ajV9H1KGGG1mokGmZ3k/8+q/C60pKSK66mzZQm5n5+D4
wHvCrUWucXW0ObOJ0pRPlWjch0nIXK98TXyxra+DXM5Ri0TLP9DWioW643WicOYE
B0gidcWrDdZRN/7FzOaUIVTmzQRCPdSPURidfIVJzXt8WevNl2tZCkxn+lzy3tsW
woezoS7IYejcVdUvQsNuxon8GCda857Tm7f+lVmRJA7auj6V1iitgTmIkEkT5Hb/
hb7n9oA2nAkq6PWpiKoN7nW8ONjD19KYX3Woc+ekyJcHdo8CRvuYmw6lhw7NJ6kc
e9gVZJyTHQ4aO5RjbdD+PqGeH2pH079LFfU+6h8d9h6LhqyQf8gt1x/rziF8ekKd
whorCRjJqxqPkAAqMUDtz3uRm4FYWxQWKVzLOLpwcU1sVqBqT5MsWgmAxRWUzfzv
18R6taid0viWGWgp7xB5O/j5WzXsncngCYkFqwc3lJMcuAeUFCxEzCGl9n6f8Qbl
WmC1Q7RsCIDntlki0V1/VAeKzrnT9IGpLOhYn3STFuMAmulBClYU4ZF57uvUnK5n
Aw4e3DyIcO3JUkhDpX/+ZmU+bywxojKfkPdiHMIpVyj2dMkKDqQZeJ/AKumylyq8
KKJmqNU7uQ78ezkBIhpbp62gMqiAD+nEushM1l4QuZS2OFfliOlGqj9aU/+znuUw
miADhS1BYpQ0NFblPRuKQd5WQOo0xJDI2H2KpLES0uM/9tLU6uHv1jzA3EI2i538
iRq2AR3x89KiXzTgrdBc4atqInvlJMtzvOkR4GhbyqqOqdl3ulw5wG0EIf2JF3Gc
wwij03fmJXg3TUzm/jiiIQLUimC1+xTRoidDGqOfXSzmzfqZwSc0L5kpwNEb9BL7
8qI5Q6pp3LAOeOU/88Z5G+0jzyeqDVZgKcqEZaiPIRIsLiyKx9a+jU1pJ5zpYJ8O
meYw48JsJEE4mn4trHUrjoKlEeoiia0vLvunu3qQX+AAmdt/OWd3OnSnyY/Tljs7
hnVwDY7aI+c8cvyEGYjdbTXA9YJvp7xDmdBAxaNgV+kcpZATlXcofISrne3nyMOm
TBk3EPuiyffvLfJyvZL/A6owml9W+vKvRe1neSHcbUb1qkLtvfSeqgo469XUvXow
EOS3fw7/QRBQbErqbnlBBUEp59gR9BJV5Jdra7h23aShJyH+TyNilpQtvDeJ0L4K
ZFO0ygSKdry94JGtB1I4yR6ZFCwff3W3m9V8gjoxgK9TdNj28OkQIp7v7vt0nyZx
8yhral6k83Q87eBAFL1KKv+q9ratPQKehzUOZAbIvzzqPN8sYlzvqr9qGane2AoG
H9nryMHG35Qc31ytofkaKPqNLU9xiVXxMAFeJ0bVkpl9PcqsLfNCPGmEzKIpyja4
bDj6n012BuDZydlJMoW9z+IYNlRdk5qCHRzQs4bIdaY6T6jQqmfuxcrGULUiYhMZ
IvtRPzwS+UW9bplAH/4wYS9pOG/tpYN5yTqoEicwHjDa2K+Km5EDYTy0pzDhvPR2
EU0j0or5uE0iBFHoyhGK/2sGpKrR6cMeP2uMuUouDIBt5fuzNrERE5NWSVXpPUaJ
2gD911DtMDxGkglfLm0N4QYk18JEj8SByTRy/yMhyZL6X9WNVVZ1kUMb1PR0sMyf
bOGP6Lt/gCcT+GI0/0WpPxm2ft6ctyX1l6gjhNxpr38AKr+DkVRKjI5guqR9naXg
qprz5zltdoDmLc4SsuQxAdbSsvW8v/21KYmF8Bh1heGlcn36Q8+y2pQx1Z70bcxr
NntqMl0eRphWJ9jMnFf+/fjFP0zlWW7iVN0N9aUhEeq2zxa6OPSbhHSLQpm9gmAO
jI626T97EediJVpMR2FWj2qC8fJn8QQYgnuKWTo0GDMkMVyB3+F0436Vs+gQMn/W
baN6n/cGXtd0JJyx+4pgeFxK7Ify9xNbnxgP4OCIgGy/faRqiT/FjDCJcNzhDSJD
ua0xEBvb+xAdBFTtRtjib3Ayv5vAMpBSAn2mpiecoM0ozymS8C7Fk3IE80p1CJh7
XJjwi4AqKsVdz8zsnBGoP6rZE7XVNhmNtivYgQCggquFDDd+ZuL9lCoXabYgAkcp
eN7glM2m9rZzXTAf5V2NM43qFZwqLB0iCg0VTdmmf3/3y/BgG+CLyHQq8mZZ8ut3
2w2wgM43q08KpbPjMLefs+Amnbxntur3/p8aIzKt2pHIY0xB3xQZtwX00u3dauti
LqM1XvcqI4D1NLnShxK+qRTgAYKWe1SxMyl45tmNLWptWOz5kwZl6kVToZzu86W0
cqNLhFLbGqVnNvU0WCgvVe5BjX0TZLBzBCHQpsE4jNK2LUz7TRow/Qeu1GNUzr+l
VBRYpuyQ4h50ZqrJzE6/zfPD1k+I4zHWChbI2DIxe3QF+SU0VtuTrVi1DP2IMbij
YhFb9kwZPUNGErw9hYxtDfWOJEvVUe6mmb09U1St6j0SCEhqCE4PL8czhLsIC+8E
fsFPy9Zkgfq0s0DIUW90P8iF8HoIT6h8jJFS8PhAEtjVfYFDN7lQauhA2kVqswjf
0JwmCPY5S9IKkAh1qq6aQrmecwelIdvWlp3GUPbdkMjI1tyfMwvRbSRxcgaJWngf
vGx2F7HybY9n2ZywhilctjMA+lSYe0EpfPeZQzQNOs5VbyHHE7VSgBWnuzlor0ws
Kkc1fYxZGGml4KIiepqUll5svKMNaDqIdckW+8k0KQ3htlDNUX5vp3GbAikjWJdY
lmErJVdtqWx7ZL4QAUkPpt/zE3uyMp0LjtSRBJ804Ct0vuSW+jmpHWUyI7oRhQx7
zqPddX/SE+zFPsUY6T2bISF4XXwxAbN66UmQbeSIX5j55+trFWC5iIwW6Y4eL+hV
k6fCpn2KrulHj4cB7khaS9fB7Xh9LgSBlhrIUfFV6hMtRibbeFQbv8jsnNKFsU4d
uEMq1PRL7l4p2pcH8a2iw1QsIc0nzNwWxLj5o/oYgBhDZWPuWH+nys6i4WRFhI+P
cwif5lSUgAFN1XcWH0wDP4Kf3gNZfR6wT241D9CsDCgAYnBgSyyTDgqCVCbo6oXK
TMuwWBZFtfrciC5u7EjhAPknG9sxnttBjG2x4MwM9s1puWSgZxBrUC00goIenPmL
msZCemlZIXwSgM4SEDuPGLA8zfEc6u6yK16nd2WmMbjnpma8CcXKF1J6fCcbE5+Q
RpmlNSGNZN7jfGl8Dtbei2VfMeUE6yftIjnOtHivyWGwnRF38BJAU7yKfi1+WoDr
usOaeyxORqoDSfyO1624DQ9pB4imSnR9B0ZTqT+I62Kb4NbbotnSNmOdKHQYvgtO
+phBkgE8S3+YV39CDtF1kMuQxDfT1Yx8l0dGHE3rxchoUmBLNwL484ggF2Ig9WE7
8soCeXwo13uyPQj6hJeJpR+3zV6h3dwPSi5/pzeqckbV+s5B3cSKpamjj0nmghAT
5HTMPY48viBTGhu6ueMJyM03J2ox7HHPi23ruhx/5p6nEJWfdtJlvgZVYVUwwAY2
5aC5bSYLMBgwJJBIM84MuTz+7koYNfmNFuaZJglDerOLDQU8RQnIK8EpEtNKfgM5
bBUjPTkvXT93hDyGncxBpum75lDD/r1N9KHSBIYd+RCcZl007JGmyuZHipLqz7Y7
Bs1AqRjrjo8zWwDpjcQiAJW/6LqENOKMdOJSUs5WZvpQcBalkhD2iiYwhJTgFb1u
elUDqpmKTYB3p+vfnFc3BgZih63mrT+rj1/55JMmifxRGCAljAHhovZtpwHwRcmC
LkLbWyfuTTUw/8ppCAm5yNdwRhMqJKXHoGCOcDfH/2xueqFjz7j5vR6h3NwVlIpT
+n5+fBa1QxgTdCbtKjwk81Jvnxr7TaQpbXVBLg9HVKhD/0uPmtqigcDxMpdFY5GG
U9hdGMsjM/zUNHfDxSvbQXy7VaieaB0Bl/Y9n95WQ0jmGScOC/Vj3HOMb5lfRCon
WgyCMkk+qaNsOKP6OCPhdvpqSbO2I6LQWEPqCDwk2Mj66bvKpyokd8TK+42T4SdD
lTtwwrkI6HQTkg5I8S60T7d1cgGE80qI+XKztmPbkK8OMFIq9LFSDu9/gtA6Arw/
KOXNL3Nz0PcmAXWwIoSeGUTjo6W6TdUPBCuQYoELLasJMYuLQyVNLdCbpUlFY+9s
y26rcEjee2yVqS9EH5GFePUf9Ti1JMuOZon9IqoqWmmmq1q9P2aCcRthdLYxMXQY
Z4f4v5EYMGMjzt83ZzwldpKzCHiqxW0siV5erzBOAjlBP1SKI44n1N9mH7qW6lKB
oxnTPYas4UUZ9a9K6biQiqvEmipba3wKf/JD8c2RrUISHTHemI29UMFIS56whgCL
EzYozxXGgZ6Hu8naMWu/wVuRZ/FZBlNhbH+Pg3sObYFj/iTD5SNp585J1bdQ2Ugs
YHH+2ixaA1IGXaRHMRpbPNAFKmHgsxOlhJ5xEGNLiCbrBL0Jj2VmaXZjKanlUlCo
dp4a15iK5NuxCBqV+1wRi6si5L7gYOBpzs+vVYrPFFj4+3ZVDyQPhgu96feqY7uq
0wdaqymKi+yxTp1tSyuLDmodWUaMpU2jhdKiZILhGiR3G9yoW/gDBAhvTVwPfcAY
oOeR+5DwLUKd0NNeRlyHEgtzba9agFKEynYTwrVcWbC139uZ0mYjyNlN8MVc2I/U
SamJhTiUeyW/wofbXsjbcj3X7UL6qz3P1aXqyB5ZslrRwK97VxCwbQQjHYvV6+xF
Sm8ZE6QNY1usQoqy1ptu9MogHCHvPxgjV0SfOulIXQ47rJSiV791yQDRfjq3kBOW
BaovxvadhkbMQSi52n20Dw==
`protect END_PROTECTED
