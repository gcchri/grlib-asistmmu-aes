`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/uDLoxvsRBpNh2B49KpebN2F3aD6V72AJWqutmdLI1adL7n+W1LCbbgE6eGXr9t8
NSYU/EoeMFtSH4AVK1OLMchI9oAdP9Ng7R5CV220gaEMdf1f1hzHU/jeO73b5Gha
gZMQwNVQMAfK24br2y6SsqTp7mpFGU/5kj/3jO1JQA/CUy+4epIYYYP+6eEslHXO
RhXjaECRQtMANxdfhHC92afCQi/+Y1EPa0qagRYqcVatYRkCOAZXi9d/fSRCYNel
Zy6Zw8xmOcY2bY8HMEfq46DQwEF672UPgek3e/EUOYVeC9VAIDdauoRPQqtI52yG
KhYx8LUrIPefAgjRobm+6opdgB5riNmhRFNgICW7jOhw1zVsofDR2KNG4r1H2hCi
AzcNEGDTKx7sbPEeDDfdnc0eF/yCrN+NQMSsHGPm4cJM20Qt6PQhJVfHbSbUqHXf
`protect END_PROTECTED
