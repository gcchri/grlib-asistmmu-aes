`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5/WE0lBKkFcfNcsxkUhPGRpnDIMEY3pZerv9V89CEQMis4qjfcz2h5SX2HZ+wKG0
ZynPwgfm2wzyXqZoV/6WrUR1S4usmsNDuHj4bmPnea7GMvw4tFRArPZBnMOu+rAu
HVQBQAqn3jk6eW5oedeaJV1fM7lK91/BZjLGLealXKrQ1rnqTSKwpYgG3PTT8Cfs
ypjTifXF88zexVv/wO0HbapZBL4s22afaWPtj7QzceQMR7SDou5wSYD1QVYTWqZC
KtMshSWlcCrboOMN6XF3U0s3O/h7h5R6tUCjYQF+FL26cqwqj9vkOVpyOS5UvjRy
RL3VvY9UOWmr4Ai8MdODfA==
`protect END_PROTECTED
