`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d8Pl0wicsmDEamZLwASo2BojtICpcajf01EObcrXT9uWA/lKOSWWH12CuB86uN1S
cYqq8ZH0DADfV3PTr3KYXger7Cp70KqWhPj6Wzg16NF2Ut5V6MURDIQ9oiGKnhwa
tNs2kT7leit2wwEXYJw7LkbSGtJ8b4qKQzZ+c94xRGAS4YiHk5m473Nf+egoGBY5
euEevbLX8v5ep0Avqyxp5iZu1bfwAvQhs0AxQF0oOcdN8S+YfKsIUP7JDj48IYJp
z9v1FkB94HLiY5BNiyiPqh4VZU4VIYxkKR9fhKymnfBpvKv2/+CulHPMmI1OWvjL
pTo7DhzGwGeiZ282KxR3JVWPvAR62FwGy8KtOJzVz7wOlWVFF0d7mXqgnraAx7VV
+myWK0PYYaazlXsTxR5cHOlyvmQE26Co/pvIC+X6PMtkOprHn7XEhUds3et3kGC6
KaxYHKeyomSEfjWIIHaUxbgPy/xX1S+upjFlBv+NUdJjfTvqtKZhF2l+H1WPk8aS
5t4lbkGMBTY+r+RPsFVSd3MmILZ+dm8Aj1pNxNIHEoi4GkoCyQkkin2bRiW4L9K6
JZYBt7/K7v+4Hhhkq2lxT6/sVouwL8VFNuXNBU9KNp+n436HmPSyaZ2cx+cw5mZ0
RNeOKDx66sd/uLRByQAh7ibEjOaOAmV+COCw8dkDwHHNoVzhTndddvDXiLdBfH9L
sdJ1n/R5wKM56fsoL2xoifJijmvEE+YfA/lichaLEWTRuOw6V0FTRFp8HUuVkmsG
ec3RhdqHJvqGDKBs0Y8S10T/2ZRH22vdLgfSOkolGwJLuXyCPdSxG7x9B2xJ+jeo
1SwjNX1mHaWEdGSYKOu5VDu9g07leq1fREWvLdwVM99dF5Mw3srewVPuZniCp962
OzjFBLLrkTZp4pqei6OLuKOrv4vwoVZeFBSSUe0Dea4ozi2/jfC683mgh+DsyxU1
kOGSEULW4eMz5hj2+C1mJeNaORvrPJaWoU3L2OKdvVBAtosGK6OoDSQuDwhN1BRd
`protect END_PROTECTED
