`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qWQLbjpldbDSNK/E2uoVITPgOGTH4HBPSgMgyyOWqATWY/xACU7wVyGuvdWeDFYx
ISxmvyTNocE80j8ZeZbArwuRZ174zci2+hI0NlrrLOBo/0t9P/XRBBpCZFE2CA/f
8/R0jn63jyGmxeZKGwwVny8xVMG3pTpl11PyEldBttLH53zACF1IKTI7fTWSbAPW
5sWkJ7LfFI22DylwRDbagcQ7fmF+Kkz258sGaipBVZLgdOIfQ+hYridm680XehJv
wptPiyR+dUaVH6h/5rwxUmItRQCy6PAQRytXlptPFks1LO6Q1NbecToyATvanV1m
KKRYXURTQd0MkYFySSJpA/2amba+0rEOLty8qeUcaQykor00gRdv68z896Q8TIVS
Gf6pQuWipx5QPlA0Mk/eJwaDBRMk2py42lqbDieojebTKC/cfTQHBlymYFnF+rOe
ubfpkIkijqm2SkgJtxd3/IVV7yhYqmd5/OYp7udEHSI=
`protect END_PROTECTED
