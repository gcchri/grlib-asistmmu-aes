`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aD7L0IpMCK6d/a07mwrQxGOvBLQy+pQNtLCW5Z+8p9GhE+fUWNkL4l8QbCs36nnH
J+EV2OIeMBu/xmBrzCLlDtcTPP8tu7M+AoCh9EZf4/WaA2UziQ2LDMPE3stNMAOj
LQPzx1a0MbupQw38hruRrkxLSndGIWukdoZOXk+BjR4JfZIg7gtQSeS/f9vZTyMa
f2AyxF6qNOe7I3n+CJPH9t6b+oVz8uPJ6iVrzq2+m9GjO0IzVogdM87kUbGTlJaD
Su6M4MCUWghR+tmr/HxiyA==
`protect END_PROTECTED
