`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YGdNym+BRUZGbqVv0/OtlQjhPcq25D8F344yv0vAvU6qqceS4voybWHuVZ3PeViY
BoWJY2YZi+GJFQmCn1PAbWJRQqvfdsFFb8TflfnnRP6qArWVbEI52f6TuThQY2Ty
+ro6DBDp7fui1IZATNh1S3TVx7fCMb0SqquTWpyGM+j1i0rqvh8ad+qvde1o3xHU
noh89jcjZv8tqNVZ38zUu80g3e+R6Y31QZ7HREnpoKVUkm1nB+O5xKKWNVvZ/bG8
6jTiGIaVHx9426bMt1mnvQxtmhvWTnqf8kr/ZEOdkviVSmlZFkyoX+aLmAQ6jj6d
jU9z8ohZLE6CCGuV37vx0/hWsKbTb1tjRPv3cDqgoNj+kPAwv2PK70kNoXCUgLag
Axwa3Q8EXtRNG50Q85D8Amq2Dxd5DTRWxOEI0ZE0+OVlCP83QpIMYF1+2Wa6DqaH
fDrkY2Xr9c9xdQ0AwOFR6xCkALTCxTjR6aUfn8R6FlYJu2s+q+3PB3h2+78btbuV
42WmdAepGvbWUcLHXB7EHUMMfMy2twdVqhcmvmDvHvo=
`protect END_PROTECTED
