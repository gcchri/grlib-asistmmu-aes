`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6vA/a/LV1XV8sTAt8VO42zCjyYP/r4PeV37E4EdICWWyv5ZW0Slyp7aLR6CXENLE
xrr9QvVhDKVN6q9fs+0LlJfmA5Q5daSY5KW4vez7Gn3jRZRZILaOAjkYjBA0ko1R
1vllOESIkWsPhoTKtAMuASzwPK+AtVlqrYvLsLEkfqt06EjC9nuJIhNdbCUKrvFo
XDkjsbWQ1iJyNPWgHbAnIRNLoirlxUgGdUK3WZMQXFHGUCUGDvTvTBEDhsFIwNsI
CbO6dHwLSuLZQn2VySHDHR7PP7vwA0D/prsDxVdqmjgNcis9jqvqod7Gwrr03Xph
SZ4Ie/qW38sWo8oNVLAi8g==
`protect END_PROTECTED
