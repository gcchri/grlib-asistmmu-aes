`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A69vDLyTbIaHBoVUqTn8nKLjNtIwZEYbPZ6GkQZfANVQbnBx0w8Avq1VVNpfnJuw
ZgnC2p/YiV0QJwWI8C+168ue4HOaHL3nwm0rNUvSa5utlOZahNjCzLlpS3q94XRW
zTfZcowUaPjmyGCdYCganeO6/SyZCAP3vbb/PkS+au6cj2Cm76s+ZiO1TUmq3Pd/
IO51YCpy40kl0XyLkmRcemCuJ8FzmgLCabXVVru/Ni1vcMU+/q/AEEZfTExc3DUq
u+ODCJa7p/TtVvKi9jVQvcXS0/qStQNjRpkLbBiTbsOTpoQ1KwX8MFOVjptl24uE
Tr/XJv92N65oxAnYTEJ+ag==
`protect END_PROTECTED
