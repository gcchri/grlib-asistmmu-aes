`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VdCGlAY3mc4M8sbGDHNsTEeAzJQxL765ra5CDfzeNIv1OSwXdX89OzK/E0Mcn3NS
w9LFucMj1eu8+IU0IYKoK9OZsbbFzaongAuzoLqJXpLJlWeX9pfaBYI08cqpcqpg
JJ7ixSVXLpx5ZHXwm6pktrj5C5jH3oQ7RyLobe/8tsFNV6i8Op74nZLqKdyaYfK3
aZDBalgah8TcOz8VeAXN46OfNrxy7y4DJBl/fJvsISoG2aq2lLWe96xx5Gyx/gq5
EzIYrlmNA8j9TS2g4kpGJjW2zEWq9U2x4XOSKEgWr3zy5yoet922rw8diMJb8anl
MXctjqr2Qz9hO1MijFTw3IPgQPKSJqrlZku/R/MPnieSoOaoNVl90SN38+NZQ5V8
jAEWWfBKJJBKO5s3sT3VOGVsPrhewHb8q1YpikRu+aSRXPyENH5fn1U1V5i7PxmF
ixi0reR98GzvuKJbHZQMyRjEYzghj6m7Afogcd1aaiKChOUVUQzdYs70tQWzvNxb
rEOd2S3SBpGT8VOgWf1A+8HTqiWzszLR1wHJV4kNa95pLrjczlygYyuSmwB7i7KT
tjfEAtynFofyNcKIRUQKqofTALpmGJmQET6Z6bQmuCxCQDpNbI/+3JEeX06uIrZm
JlSGte5iXHCvp3wTpxaapQ==
`protect END_PROTECTED
