`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7eTxpAs+FQvxGJfXd68sdVHoahLmBKN92NugKJ1rIVP5xkVOZZd3UQ4VErc1VDeC
1Eig8x2Y5K960QuX+dUxfcT/E+E2sD5BgPFB0BhuvyUOy2GsUtR6fANxLWhtJRad
e6KbzOHl2Pdym/ZIF6cqx9k4GvlQDY9S6xUZK/+XapBNJA4p7vHhMX7xSHKZE8zJ
tWIRxKj/h3C+Pzaz1C+i6z5J4kVyGXba0d3C+k2CvofGA4EDDQAxGF2jfIDmyK7v
VoVjoShJOmRR4zCvoYFW62tLSoskzWmNeql+yOHUf9U=
`protect END_PROTECTED
