`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
73t41mHrw8yKjR+Rqz9v7jCSkrraVvl516szaSBeRSX4Cymq1spbjxn/I6gMP7jF
QJuSOV3Mz5AEuv4ofFIDOG7Ln3CjPxNXctavyTb+JX3FeoH87yhj+ItgwwOz66Mc
RxJWlpyZI1N8sPnBRMV0pCZuoKxe32O37lrlpzEG2Qlcm3UMHScazadFq5gUuqUz
6ls1sdAuPFsiLFYCtWx8Luf8HUWo5PWTn/bNAvH6wpQ2yVZ5IYwxbhn40be4PJe1
vKVckh5HF8XJxGpdfhAhJm3IwwhcAUtUDphIpdsTUtsjKYI3k/7tOnIySCEiCWoJ
p7ttLtQsO6W4jv7HXqY2/i5RZiD3UGqsa2j/TLcE95PjuhA/Ixbbaghd9Xhd3vZQ
Z40gOztaybTmAtdyOemddaBpIePAPqdLbfvriClxuFhhxazyMgwoa+jC/qODtscP
+V0m+PY8g9zhLBqS6GzFebxEXxSwd9yaacCsls4zBNE0va/ZY12ID099b6L3zr05
F4j/zi/9bpNwJGzg8HYNwtrx8ajJJE0eNvBnGBLqEakaEn9+iG2mknfSzvmaO1xB
9jQpv/utR7W1ZSmq3bHleFvi6YB9NK03PJAlEnV+Lj0=
`protect END_PROTECTED
