`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IkQnJB5yGdpKvMA/cPbBCMXxmjUgUpqmA6hXyqdkqDIZUhEy5bA2dycSCzm5nVr/
5Hb6+wy+h2uryyTS+1Z/l1J3CdZ91YwyYCdxdBNYGQC0+d3heGTsSZm8cSjHO04o
G2RTcmlipMxy8mtIwm2qBbikojw/OsKJx+BQx5OXPLR36loz7j7b+/Z0ZPsjyj+O
hdnrhr4jlzD2jPpPEY19eb9XupM/GpI+ka0RS1HzGaThoSKWlXPjULArN51zpnPV
OTy+JEEaT2XS6WvPco0lp+CI490Zuc877YxH1C4njC2TFqq7pTcVVOvIfZJbR+m5
7COMBcczC+bsmMRKCEI7tuNrBmAz0NTE1jzL6Nf+NO0=
`protect END_PROTECTED
