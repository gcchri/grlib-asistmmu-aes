`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CksCAipIUKkb4Pw9i58VI+vTU2m9d72myyO64NUD5yp1OQFgull3JU4RyX0IpMI+
YT2pj8vxi331jsV6n76PygYFzN/850pq0QXcPjrutS3ACWFPYjtrAf/bgoHbVO1i
TBKuM3h3LA1RT4CCjwYAmqcKz/x2QApT60dmc7P/rtR/doSQ5B5EMYHl4owEra0S
/0PJoTFeau42Hi33apWvPkv6qQferOVeLiTj42Dk7tAGJ92qhOxG7LPdJw6ua6u9
xRBgjeMD7Zd+XIJ+EQkDlEDOjhz7O2YBxE5b68t/jXTw0A7NLPwYFI6pg8MbjeKS
2fXpTW34fD1cR9rhSgS0DGnWpqRG6BULfVhGo74glOfwK5ksZEfwEsDAs5uXX1NG
cxUdYqbkh4CzxLLHHIgM9ZjXxr0UngNYxm7F5Xsvw9HPoRF+URuucU/USiEUy6uV
s3ZF8K566AUDbKg4xV3ZWgnZ1qonlh9mPdleBEWXlsM=
`protect END_PROTECTED
