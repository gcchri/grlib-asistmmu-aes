`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jCEqv1J8CpTXafyNFnAEgByciGbea8+Gy0KI7URM0FntqT7hZmXywl7GCY21jiNM
fzy4Is5XWq6ehbfRPFnKkUZgwpWPP94DC78cAeYgYACzz3De5BWEYePH6Ja97z3E
4H01qSui7Yx7j7uWMbYVTUhtl355stQaf1LD3m00a1aV0E5i6pvAJ0A5UtG8jHwM
SN1GqZpSTZQJkHh8wLLIFTm31Uf0jVL4LClnb2fyChBWFFpyfkm4wvKARRP8KiOq
cxWTpBPnvymKMaUpfglkUipVAwvA1qWOojerFsWe7pUwmndRQRBQJnDNsqEO1lf9
7WKowYVB28sxCvhBj9/KFZvFuNMKssKy718KP2VTTTFOF1k/5ihTMLZCS5bg/yAk
4J85kpEDtXpZFkv9zaHF3ICYDRPBN7Z+PxiCWaCPSnPS7dQjg+P4I4tq+PGCNuZn
XKTdQX9CTxut662u4UY/k6vkTZDyXlHykJuQneU9GsLrdl+1qmcgFM/1nlVbB0UZ
E5qCyGjXhfgys0akdUPovu8auSmevN34t1bstZTFJJI2CWm6KKdArSXzXXGp4/XF
fDtRrQ1TxqG0pyevUPIEIr/OnAIuSchVLqu42ad/GaCeiKjdGznY2xlVyBoonZkj
6i4VzratUE2qRfkLnRG2Uve7lgt5QOi1AE9ou9TQequ67rdkj+52Og35r3H8bDxy
u/2h7QZVY0Xm+xUpLludrzX15bOzJLq5aNoFXvMUlflzVkiDZRZZPWSeIFUHB6wW
APQmbdxghfFzzL5HJ7dyxgIARruqrIFo2heimMPBLUZixOdhDGlfL6ybdL+vo9y3
WDv+3FxrG+0DPeMk1JsxKYzR9FMWRdOe5rsFwW8oErnRYW3umTZTavw+f09JT8lM
XmX2GHjcli/y05AQpX5zAcn9enuJxnLKMl/mcLJ/OT8WMcQjebWd4QfE7OWxTstv
QL1ZAssjZ2hZINYGVJomogS7lx4IAHkyo4gpiJugHkuYyMB28N5ns2AA/Fwje7Bt
zdu7eadoZkthlvYOTJ5N4IQJFIYQPmtlSvksV4Jpiu2SyRjEv1lK8WNZO7iMeJNX
KucDKoVULAaZyqPF1o4rr9IX+Sh+5Vy13Gm6Jdn0/1gMdiOFTNg3VA2OMqSPGfSI
mgRrc8JsYlngB2b7n05yxFmKJAhmnC2SOnw/esGBj9YzKHys2yqtqR11bu38I1W6
X//s3l1+ZkWcfrQcouaBversxiNdQyl2vgM9MLCeK7YQ2y9Ya93oWPdLmYFvuFIY
qD0BdCOize878BFDQ91PnMg08KrGzQfPo6L37O9Od9QPldekJvD0oNAME1rb4ZBo
uNkGicISnPz3y2yEkETL953jrhoRtkjJqRva1nnQgYG9o/JgY0EvFDuD86SAEZO4
GfDRf79pVjAI9aTpScEGmR9RmowEdbQSQh9OdKS0IiARLpv9Bx8iThoGXwS5pPTw
RibV03kGk70kRVsJzk31xLare0WgJ1dLb1PknENUTyd1yhd39Rf9YO7TGaJLNFGY
xOPJzR3CNe+26P3l/evCtfZCXXXDOFOFYwf2ARpPlsm0jskDJPAy0kbqLpDcdTrG
VFA/w+C51rw8mniSIEEScUvruapzDtZKV/F5UAWt50T96IGjQmXLRB5BbgnGc5qq
e53jFETuIrqbxQcRVCJBFfOiFTW8v4DJ8RDfVAgV52C/3ctgf3xXTYpup4ckP52v
cMKyUwgMMwJ91Vg3BufCERcatEpGa0m9G1ywhWiiidVNQ+bTELiixlcolMBQlqjm
KU5MUWQX3L6V8gtNeUPTkP8z2MPUuAcKCjM1yk5TqbgniSVDo9v/uuLNSGPg2OQi
woyvFRiadyaMvW+Cy2y6RA2DMUbuXWjIMJjzZzEP/o0+eIVRwKsrDsjvqRB3N5AY
+v5OX+dUoh2sixUDl1Sbdg417ATSdQZbgwHBu2xyaKvVc+9K+jPkgLd4py38DU/S
rVRU4G6GkOF6bweXDR8UPKYuqX0tv4PbD6S9qMW/f0Rn5Qxsmdk0u+N40S79aAA7
uoQNL0hl3nUVc6EMdKJSFLSFFqKUwZ2dezsEf98xQnHXN1w5MguwwUDzyTiSK4o8
Oa4lewJpN3mI3YXLY1mwxr+KpFXjjVAfICD9hF3j1qepU9OfwUMXW5GZ2CfjmEEI
gyrgNxC32L6inIroIxmjX0/iVY47lGORutxdQatYLuQL832qJcqvLOVJTsHWq6dl
igXiqkhC7Xa507Hk+z07pCcY5uIJN08LhBrBXeYB+STtTHcSJFUgjlfB9D8L2gXG
etdgxHVTJDiWriCU7wKv6h8tbJoeKNN+Amjswa4YjyYYvQOJtXgs0MTFi8QlGviR
cdl5+eVxtsB9T7uWEqUMhVZy1GkIEgnaspxjWZaAGKmTyh6AzT4GOX0s3+18+RTY
Dz/e3xPCOSqFPORKDBAVpOYITu0NZ0ChaXX9R3j58BjAGKVqgJEWF9AaLcC3KOH4
H6mP5vRcCnVwI0zcUWQcb9GKpwKluxCcepP8ODGRTd6z+DH4ag7ArykT4fpR/JEn
grhI84eGGOsH17RQbT9RHuwCII+HHhC5juARSqy8Y9oVnPD/AXMs413JC1pEIBLY
JhEEVWx+8xz6Ig647VMXkqxFulGjzGjk301ZFpauFPel2tue/mW9i3o8DOxIo1v8
Xgim94YqcoZkCV5TyxcLjXViS3ImrJpJqyNInudU5aotldwY44gvxuNbbnXGpwxC
`protect END_PROTECTED
