`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
knPFo8lAIDVelOIMRB6ah5frOc0Rz015y3TURkf6Q0pO0acNUSSi2qY44fhre4Ek
1FA3HVt9TpZACsf4j2wqFfQjt1sA8rm61QSNuAaeI55w875QaS0KveE9itUJOLs4
F4ASyDzVTS7wKwphsrZxWPt8GTbxvReMgG/SLrOXNuMZ1qvNUOPRh3dDewxtlSc+
1eoxor9ZxWgkRzF7CgsrV8qwjdEiiVAm01RCCkoPcR6Ps+qFGFSevuyV+hWM0toN
P7IkfKAJfC9GG91fgB92meQnbpudiSaMbr5ErRNQQmcUhuzWFYLK/cU9QjU5pXQe
oRWw5h9W0r2JrMvm4M7FQEQCj9XnptvNlHmKOQwqukRlZZJsqC66SocdeJr/N0k7
vD3jgEZNoQ8aQSY9y0C/FeUF9NXTxsWc/wkrAbV5IRGBI5WqC5zbxc6GPLpg2Y7W
jVfe5psRZXfzAqTkqJ97ig0FZiuyW9OOCruUmxnp/On8rYUv9+cvkuSHajuwsG4O
UmDSdmv2u9wT78Bl3Hdfg6q6kSLXjB23XE0uJh/vizpvtXqtzpabNIEQIY46W7EZ
9OQyH2VT78KdB6QtguOYlZrlEz1sVBt/LRweouyIuTHlxGQ30Fne2ZtExQiGpArQ
X395g28Sa/JkXhsDOS/EW9eBHdX4lSnnf1Gc14NvPFbb9NzXWQ7Jj3rVavqIgxCc
CkeJz0eAXI1u5zU6p9Ky5oxWKwTVJpYbLn2SJBhShRdtjqp2PlPdd9gAhp1lD29B
ibAX7a44SXCgBkIzWwyV8kMxx9F+7eWw4heRgfotBHyNlWV2nIeb7YQGojH/TmKt
nZUEVJqL77T6r1CkP4lcKW40+E/N16PetgL8u3PWAWrppQ6/UZoLRpjxfDe2Sfmo
snEkYblynES5tJ+PrhVtht4w181Mw15q+xbpss/7MhRCpJkPcE4SniY3s39zWuSz
Mw8jc2oe4kjZ9LMpMpialo9WreVmJjODPWLKBASsiOra/vGdXQP3/pwrn3VE9Eao
FF99f8tGelnaphyZsyx3WwAyUU6lhBnLkaVOZZKIvCsw3FWnO5M019v4hoqR00J1
DFHNUlPu0jRNUf99n5IWzA==
`protect END_PROTECTED
