`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d55dTQyEK8FJgNBM5EseJ/Jr+1YGxNTmJ2aoULwMWhSwJr1yMICBsUlzbEThkr+I
Xrg/DUsaGnObFw4PKz1pjRWDhS3GddqNxQioiXLxmJUQFJIkcYJg9Nq0U4Vb4vCf
xHsNrFQ2NWOO7NzHKETvEXWAkRVOgSemcHWbNMtxpyGs9f6ObatF02yOqist3Ue6
BFNA+JRyfXOonCfeKjOSpmL8TViyMlCOS2aBJz5CDf8h9DVsACSEgS6508vYFME9
tvKn2aI+u1liY4fCdXLtlZoOMZxWko5TcoEdMv+e8AbRMR0I0AwmXRYa6Fub0+O7
/zJ2oeOW8bueUNDDyDR3lYjdySDDCtiGcBDAIONuArRl7mTxx5WjErf4OrRVjWV3
ekOhzkwmmybqheNIvbKLECe6xWt6xeFOVVeo2kcdCFxs2Cyg6YYnPLG2jca7D1dy
QKpAZprtm71xBGF8WNZP/9hsTQzNG3tWhocvnU5iRFP9wu3YMCTWDuPsQU4rdAOX
aH9OSrPEqh8wjAKNqT3eO5wXIhT6GeP7+xSw2jXnW5ROM5qMpGgf5hbifALfbP5d
GIfK8s7M8RxLL6Q+9hr/6+9OChXyZF5iJSQod2vXWCLQZ5l7FBnTp72K8roTCQ/n
RC5uD2bZtwwmJ1/VJg7vzKWQ6dhN7qzsxMmik0hxVNkEYE01ydsiNFwwJMkQe/77
6pMM+LEpesZ4y+VPeHh1Gl6RYpAFYsz+ALYOG95rX1EDK6+3A6IxvCBBKzJAtMCL
fE2jEBYey8E1LOCZcDWoBbAQWsy6ol7jnv1+NFKHyckJNOX3DYnf+Hd+dZonl2yo
FoEtL6JoZMrIVezVA6t8mxVmfjSeNrEUkbzDWiucUcR4EanCxiDCA3UIyMYYOX2c
t+EvxgnNuYtLzLo0o88rGw2/PJxSdF7Mx//OAfa+iq3WeEc+OgnmdeBHd+qImDzm
znZIDipNalI7RshDQSIKL529TJaV+qQza5ga4UbRCH1kD5JpYgAn49nJtefyulLy
T30GFKgxM6eF9RRhvzD0BB3RKmfEWVBN7RmNSDvOnYWC9QJrt5jAf3M6XxY6SnNp
VCNFJBWCOebNsm7WcWE+XEMSnsUn6p5/9N1PQaQ0GQM=
`protect END_PROTECTED
