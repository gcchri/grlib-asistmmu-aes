`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZFLqyfb+jbFbXmrX9Gcr2rG5AsMHMuEe14n+Y+EemG2IfGBKgmL3Jx9o+FoOgFnM
ktKbgkzh/DlwwZnP+dSLFEborcue5hFzXnH9Ngwyt0SbuaMrBrSHB59SrClzSXjX
OF6PZ91T2HcjDR7Bvgwj95jNzH1QBNK96jcu7LUP406HEiLuwlpp7CgYiOL0/H5/
vy7nF+Fn5KHeaNrjCCX812HyjtqYMn3Q8gsG6iMq+brYGul/y0DFJRdh/B3/geJf
Yg7FK/6uj/2dsUwdrWAe/S2UgQz5RjfFffhWt80jG/XgC9b7A73t4obNweyAFzmu
WG3E1QEVCSKvd/yJrV09GM8q05pRaxhzhYQ0VykACIxeLfuXROSxN4blz5jcM/x2
P2D0A/tgR/9ahjC4okGpkPeaK08mIcHIDW+WlytxO7ZvTBrb07IHTkWsRy65PewE
STts7kNYkJCxxVZmGn3tDSHWDplnFP8mzYNGpvOMimYyQeu7xS3FiaCabRgFaiYF
2SSqUnI7P21MnWHxG7D9PLP3ka7NCH7qujDg2kf1hxEZuOMEF9Kb2aztq7CEp9M5
soqTklCrKl4iXnn+PFcn8A==
`protect END_PROTECTED
