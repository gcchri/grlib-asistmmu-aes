`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6X4GJYIl6UWSSc8jfSwxX7Kfox2om4RBkcitCHjbFFgNjUtmAuG5Lw5B17XizZyX
RiYgFvvS51sUcfJuJRhQer7S5eYPks49T6QNN5W5yNKiwKH2gSWaZLhsNabvMMuI
vNQIs90Ec8YTkSoAJbEOPAmQ67UQxz42v5QJaudPJ0y8sdy2zAE6Izeb2Ycl751i
CKHMoV4ynyxVqLsSDjUXy3XkfgqKqbnuA837/9RvZzkBWYPx+mZRGDSuGvhBszhX
yr0Kc88aAQnLxqg3huxj/pQKMqWBzkmn/9jG95RD3++tcIab5Z3MF3HCN+B2ZSx9
sQ6yWBSdrr3MFERzunTGGhrhk2ZFCGKVd0FiqSw0+NNT9qYbH4DvMG71zafYzXrI
Ti8kHql0Yv6rN8c+wvB3nvzWVBMSPL8peA7bfPlnlR2V5unZkcDlIUe+70tDs2RO
NsXVH4oLE70R19pXytjEVYYlvhpe53xDMEEZk6QKo0S14BD3uz7rN2k+uqAF/KvZ
eBWzc4lArBJ+jEb+U8J0rfjp8dUcIKSSfOrJ1dllLQFShAQ+8QeJd+APMy7MHGMm
GMp/jkOzkkqCbOXMJbQeuLNfes5HBqJlS5H8ZcKnTJxaLcVRDA3raANyqHlIhXIE
KIosHiMEMnKsbSeBH96uOgoamOITWk6zG6hpD5deZbhc6LjDgmwOryQ7gSwHKCPw
Tnt9OacHlWAjjEz3CSoE8ZjH6zXGDy1lZ7008DsP6ZfXTgk8JMrvShPkj8r9qbGG
GBammdOXMrd9q7knz+SfuwUSq6aGO3FtfAJIwl3eLGOCtyg+SW+i3J4q6u88V3kU
PPPt/QzF/iVuszR+wY5zamW3LpOhqagwgmt2XFcEmiptbjFTG7sDhYWc9pjvO6Jj
7wectUl1vMt9G8XaiKVtHh09DfEt3WyBpWh6gxGfLnEbEGXAN+reJuN4rRaXVEWq
`protect END_PROTECTED
