`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HEHDehxy559jUkuJs2Qv15IUXFx1/lzbObeSwrbMLvZCke51/ryrgWztfjRRSOIn
AC8tdGWwNaF3tOXQGv5Fljh7tdTXNVLIiXwcLoZcyyFUvJfddEunDm0K1i/F4eha
E62uLWj0lbptMDyWqoHapFgCbMWB8n1IPKtO1yYwqVKFJufiElPwZl8Qlq4KyaYF
51Dh6oveml+PTVqLRJwdMYMOJMJt4Gsl53cqrS4zqKHnc9BeyzH+uozV5yIn80ga
8/35iH3c7lXCilFI51IpaZDOcXCb8/f6WmM7/Jegjpkcm5fMpSJ9AP96yj9TTdNe
40JqYaOsvMG0JPZcwtMt5T1W1pVDeW/j9bfDW3hqaPLjCW6V4g86JG+Qr3C5W7i2
p3vRHdaFGd8me1j2+weOI2U9bv6FD8NZZ5mJi5Guyh+U0xNVNu+bhoO4TrIKE1SV
f4wSKbu51r9DgQHkYLksCvXxAbP8Xowqpv6ztF4kp3NZRHSNn65F696BOqIrmXux
K+8/MsOyYuTPrQgqw1owHezMSh/ILN0AqrEd2ibKEuCriFKgSslBv97Vt6P1Wxz1
jcyHkli8Fo1fSnxGewz/UYYJYtObCUwZEgB+Ov36sI2ifERLvYWh9Q4ivuYwKt+4
NAUGbNxCw0d7iToPTN0+vn/h9d6ZzAChHwr7vn4ibRH0i+xUFVeiN9taJG8vjq4/
dGMa7ChwRaLH096MJUYNhi6vHeO/Uy37VMTPWLrBoSr4WVutgnsmG3U1iz51ETBH
UFkdBDQrOSSgnemc0kg/MqeEJZULwX795QdtPFhrc4Vn6vd9xSSknZiez5iFnVWX
soyE1E5bBj28bjLSsQoIEll8KKzqG4hJ13u6mSBJu0C7rezm5VPFabiVmvqUanwF
rtETfjK/5ICXAYPAFH1YM1ZMK+NreL5FEJAGARxkpARlEf0/xD0Gt9WNmHKLNO+Z
LZHSWDQW5X2VonDr/KwDjAltJ9DPFovaO61SNT2tZCT+1E21yDzjIEBWmqFrurd8
JLLLkVotiLVzQzE9yDSDoJglY3te5zXFbVliO/1AGaOxeNQwi/XQd6MmzYs0ORZ+
XL1kiR/UsAMfoNYgAkw+TRHCV7UirBij7P413g4lcKDIsVefhMHc22NiP69gzNrM
r5gwcNHq0D+ZRu8dUTHuKhoeyxLT+jBQYmYxVUrlhUdq8ZCHOXQwd3GyT2KlzGXy
irdAKE5qxfQ4OkVY81AHdkXe8gzkyqYXUWoqLCGhweFHMk3SPBz7W3ybfedAcxU0
olGi2Oh0KxTAnfOK7gxmZkXFn8ehsWJMld8w2S5hG7SonfUVJ0TVPPnuGz6FlhlL
uDMJnH5QTTrwrG9Pnb9cN1953U/suwhkn+8oGMl8SrvaDNslt5jxgd/mOxlVWOwm
PmJ3hnziupF28fOb9zVISh6N/pRYqvv2twb+z4vhIaZEqawTCUCiLQbN8m8yfUpi
OFlLUsAt1kSkoS4qU0YN2Tb+H7GaF0BDSse13/yclg+7wTAl3MOkE0oHsGfseP2n
q+zpZ49ounVjsQvBYNdUAjg0YTWtOG6Tz+kn2xj6vgIHEFv08M6YMB09U4gmpkm6
OLJIGAzq0ytpj7WQ+MkmWZvHPVUBmWMl85xdDxAE3YtSb6PJp+Ml4ZTQr13tqfwr
8QSfoXTtAtR+PkDNmOTUnvdOPuRSDMEK2mAAcG+iO7KdWjhbjX6njNmKqo6Tjlk7
yGrnHRBe71EsGGsBBb93AcJTHCsAOrjbvsSCld8fqtK0vrl5a0rtx3cbB1cZTECf
whg2seyph6Nm+tOM8K2ghmbosHPnRSSffuX2bwFnj5iDAa8UsyCAQu+C6K7HwULf
ebS5VhBQ5rfrowjWo8z0viNopNcSvRoXpHz/ijhrVegYUNev3Aw2BLRUAeziasqz
gbG7Sit+GPTK/bd/9tN9X1wcwti+YmZYx6LZZXJIW5iuLnjZKHgkENQIN5lzRd0m
2+OEIGRApWrPDKFdKSRU1AkFsB4v7X38aP6pBrIMTvkzPZz8tJWpplc37guoxh1z
ENAHmfpseS5RGI1GSrw+isYXTAnCyTLAt7r+97iCnf2Er4Cczwvyxg/kcjAIdwC/
LIVH035IXr2F/oGWftCV/wAqW6ZCdsTXS/AtFjCByxI7gHsKtZ6kqgx2t0tVzkVP
uZwVl9h5WorHxpdoK+akGwGanUC0vqOHV1zNLa7rpoQUzv+DNbPM+QUHppjEkrRw
9kPxquqnmWdboiZc0lUot7QaIS+EkSMMRExntbSl6k6Jeapb+ble2IeUsDUJEpk8
didE2pO7WkGXTxD2REDYTG+QFCtETev5ZIDdd2LAkZTh9LAeHRRDYmxG9azq/3lh
18B5Mo4767ACub+2ZUSSLkFXMDRIoV0YEgH6zP1DPyrHQSGq3UODpIuMfrF9AjaB
6GD6MYCYShI40HJYLgb4SUITQbiG8skM/MrqNfe8QA40xUU2pXGo+npnNgo9rY8Q
5b9ogTECMvYR0N333fQZ5+7cu8YdFws8p8Q3BHAQzb/hp2vTWp5syc/iP7p7hma5
dx0VLSFEN79bQlq4IBRZlXTAFp7f3NlG8CLGoiJCmpYrqzzh1jnLysTonS/ti22c
l2G0Fv7tGABDuFlx3Yrx2m+J9hsUDOUMfcKYBDtAw95XFE3fYfejMxGHETaSQRk6
OOQmg+ACXb6wSedfcJDkWOkAKm4mS9/LxpiJEVeDLSdwYvK0CqxuE0wWJLW3/gkv
Hdb/cZIYOsjTk7dXu7I1n27wPuMpv2CPA3dWiUvww9H2l0YcEX9cquM1Io6ajGLP
LIZkhEgvKyJFYmDtZ5USigC40UJ8D2wMoG3Ekc6PRkwsmmTk4xBj0yQB6yN8Tv4r
DfIg/96FjKKS2i8ig20IEVcFVct/SoCtHH6hSlnWuZrsKzCxcLy69i236oSo98zQ
jTWfvc3wYoDncRflRTB3dCKwTCUFDW4sORhSDaekewRRtx/QxO/9jXoUjuT7RyOb
7eGgvmxz4SvBwbx9kiMtEXZs7lVSH5vrGQqik67+7Q3DVaS7K4RAeSXzau1XwVaC
C0LTpzK4R+TBDkaEsvvDTcPF9sxT0jUmiwu8obZAEeG8174alrWDafk/i8fjQbLA
VDs9YiH5LBLA0oscpziLOw/4y8V+183RfKuX+tcJTKGwL20fRsmSpwELyEQmbbeW
EYJKnkwaMdYEUJsGZ/KQUoup/QfreluKb+qT6b2YIw4Uk5kipfEy7R656b6lkzGa
DYxsjKHEUF42zVWgK7RhQKj2BvAZAm3XOHNtLpIV8o00BO3VW8/JJPqS71+GiFJV
JR+TQ2U58anVheCwzBDOn+/OIOimaOODTR4P09vsRIVlvZS/Fgb6NgZ3aJJFPCz/
JiiWEHIyQR154w336+ZQWngspgGCbo3/xztfSSV9YA1pU5aLM7+R7OeVR9QzCmSf
U51cvZCe090hx4qWL03gdzCsOyezmEswTA6UnoBJDPAzbGIe/Sv8SfvcVR+iPc6Y
/37UReFiupCc+5ZCW3t7zNMGxcibJhz7b/QUOmtJOBXkL/FPJLu+0zOxJVYS1SJg
HTFjkJmR9Snmc6Yno0D9wmPCHqPack1ktbFxJJU7v0GLrdpI7vjzo6Vty8vNNWga
YxWKnbq84MbyTpyLrrScZH6/QXUn/1L0bmbI8RIo0qcXde1sFiBs2//4Jo9pOup9
j/ncKWTgnooBARliIUxsoe0N/ZEprk5LDhzudHzhcUDg2DHh4Pno3lY86R1nBYAK
P5X6PO0EUiwvVz/rl/PVPz5MmgWqt5MzcDdEqnqASLza3ahuwmbTI+FG/zS4OcvP
H/8ybhSA0+8bAhT8yqAmu1YU6m/Qd8AeQw3skVO+az4QE8buTGe2U5LtIouZAtkP
2ALjBedyq9ZdqTN5qQRFY0eUBlRW56RLNm8uZdNhX6GbcHdWwDVZacmQdunLrkdf
83wwb9dFhyKE4K1kqY3rVXTRdCoGCg+/lG4DhLUG7wGjBQfe4Yq+/KazBmNAIsAA
TU21nbzsUWta1itZz3di4TLN2+OKPIkFTrrzbG79XTnzWqeyNH9op37/XUtWZ/qT
9WqB9zMQIrMQJ8VpZZV+h1HR1xDLlXX94D5rrDGdXJZRj3u7fLI2PKs0PAhJaW7T
i9ItP+OzHLPrTlytmA3WR9V/dGPElgBVlTuel/2AqfyOEx8HiNh0TlasUlHcJqpR
D5fEvYQtng11EM78Ce+HrSpm1jfC5q9hc0qW8sA+SU9sT0iscCQ0B2r9Ei6J6YVh
cAobT6Mo1sajakq+d5u72cp+l3Ew/lO4SP9wLVQa41HN/ZqtBtfTC/L50RF4bCac
E/apCAUpmSJa+0foXnZHYRWCC/WMOCf+ToKGaxQPCFLFQ1bsaHpyq1393X07CBIf
HiKfW0KPTmLA7BK9rn49dRUxslpSOe0wSxIVyZM73qxbE/vkquVNPG0L9d9hTNIA
hQtI7y39gdunIJ8Lw/fH63zSzUzfMyl9bFF48sq2Y4GoBVdjcQkAgJKZ+MWrvNiz
xwbC1/xlBcpGt0uB7vBjAj+xRS9Qzk7qGnHt0o/+su9kHbNwFM4/yMt4Bife9tvT
7I66MFkN8GMmuhviy8kZq/dyOUIfAZt+pga1VjVdPqOS93+/iE7DhfBQM8jcyEwF
j2gLyuW9aBG+h3YBYUCHWXMK9f/NHLMyESJ/H6qxZYpQ232j202ZSenT47yis3I1
uPTb7K+2nXKge2UE5AFoxrcdhi1Zk05zcJO1kqJ/36XJSJz/oL8+xFZkwXW2XoNt
OyIEVU73eRodQ6/4FNkhHRXa9GxeIXwnlrk1w8llgAU=
`protect END_PROTECTED
