`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QHB0ip/XgroGZrjN3TMxncLKhe5cRLn055xbfq7tMyLLuHDT5+ImMMBcUd6izWqb
ZGyIdjIHxwiTT4mtpUh9Pn++pWia9oN0NHfHfdZBWh0Hn1vRogpKlmQyYV47GuFZ
lVSDhavlVCp4RUXfF+090+l4NDsA7c5nCU6iBXYQkFD1NSlT1fwo5w4VDT+6h5Xl
tCWVz8mxqZVwGv5nVpgPwOqYAzKs+G+dDsZc7ob5U+9h5mSQChO5/N94avEnh8NK
caA6oL2RLaqNQq6Ek9y2VpFAx8rt55tHHXQdh7yq98G71MDA56sOHhwig2ZpzovE
S+n3vYiyx5YsCKrnPTIZhBs9EBQ3lC12Nym8MzvJpw098bZakVh36nvrDDgzQN1c
9uWQUXMiE38n2H6cXVJaoNK7GfctBCyb7PcAbtBzO62YXdBMDkeZLY3dauDdYZ4x
TXBLTmUoAkRqm03x4NfjTirUR0YCqmSKrC5c5mrP3QcNw4bIHPuX9gIla91kHz9I
GfhjbMs2+Bk9Lg4nycSkylsHSQFdpbEtxGviVW36whu7CZORYtvC0TwOS49BUnP3
uZLFLabXlfHNlgQaRvpCGQ==
`protect END_PROTECTED
