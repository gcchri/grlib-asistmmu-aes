`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+xfvkyuPGJ0q7Ndnnz6P70E/I0eLxDBVILz0x9I+eLPlw7WhFpOIDQq0HDFNwGd8
NKUKgKiK7DknxL9Ocwz2bsSVJP48m9xJ3vwNS4JnGpfyQLj2Ilw3XU99v+M5ObfE
uf7Du+XitKkDKNCkjYfYpAa47yFd6ItLEbL6dxdkW9GpVhjjjZBsfVWW+Wcx01BK
3xJjQ2Ab1T0K4L8jWRDuFYmYg+QBbAc22uw0zX+WdGI7h7yRPwFOgnUBHt8TAtNC
9DdAspSDmP8mUNl8+XSCVmH9Xx7rVQodhh21VIco4VGRG+tX2vV2RzyJNH2gjdwc
QOYhOnNtiekyjnY3AQgaxTGha/Oqg7tRDWvRMiNgj8UG9nqNih+3h7deWwi0u0+9
MXdiD01Okr4fIq+DXuv/kBSK8as5aWS6dBqk07J4EyGNJrDMpzPJM+SfR0AbCTlN
gHt4oxnSJCPPcVt7c8w51vlN8Btyjilcj3hxDXOnYCA35WVWyIMSiQjAE1uTmntF
sYWQ1nc2bpg+djvYP85k3zs3KHKIOnWuU3Qg/bKrGwo8X7I3huYASK3XWeSHZoE1
WIgKzOEyhcMfxrmWU9MoZ8ky/6VlpGYndyv5xYOQq0qvUIzyJYb1M26nthZSlXC+
aLnohlNy8MtEOwZ0m52QQtpDEb/rUWsXK2tJ+IVdqw1GdlQJ9Nq39m4Ks/5PX/Wb
H4yAsrvWtGRsrivbHi7xD30Hw6DdtAQJhgzUyV6Q5S3Ptc+2NeNuKevU7uTz9W8h
EX6VHBhcDq7QhYZ4ADqzz4eeuWnv8Qvw7uvZq1m9NQ+97LMBghYt8aV0cBLGO40Q
gTgWsJxjTH+1LiAaiAh1JyZKyPTUeaMihKikBdZtoFroYq0NLeRiD7S6tNxza1Lp
1MM0CPse7WeX5wD76/FuNlZhc+hWZECF8tPqz1evSbOJ7N5e5Cv0yGtpqjUUU0pQ
NzMhF6fPeJEjAILWgLd0ZOL8vdyTaC28ueDAj3wK/BkreJ2bqLSH/jUdN4XHI7zc
HxgRLpUpLUadVDCsbOuMNkEzUiSZUWbswLY/fw+iRKFzuE9gfOZD0UVxQZj2hdDw
WoJ9YqByGPcE+QrFCM/eo3yQ7QHj/V0yWU46ni6QGiMApN4PGVdiyaSzgeHL4/57
bzIchQ3JmLeEzTNE1T8Um22GxFtSepBFFQRxaRSkifAIOE7lHhJ6AwOctxpPgLe0
l1DdOaS8ai/AJHUtWo5aSQBzwb8LELjyyaFe5KTEykc=
`protect END_PROTECTED
