`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XD/k/2R58fQ3v1NIZL+Ix1AhXgeIgKWFPFYYV7z1E+YyI+y0vV2xt9MuqOi5qNsr
4DzlXANE6iSt/DiB+UGpdDHYRUL7O5FeLWpiJQGxsgL6mEgszcugtzMbFyzjaS3U
7x0xbX3SEP7zsPTMztjsVqrMy/rwd4tHMtoMnYn5M+jLELL3havgd/8nYDg5Fea2
EcuNDCTCRnoD1VB81zsXlJzDaiDJhLZOJ1NuostlOd92kNZirht7Zj6eI7ZW+k/R
+b1wexHi0+kUeyyCs4GAcIc7Zi4qRU9/b7XaHPNI3ijQErJbH5alne8cXpZsZx1w
UvhqqidOvk6q9T0SZlj6VFNAh0E+0mDU9VwyQ9I1gxuTbRKqEhwvsmrneG/zkyTL
ESrMwdBhXO2NotZHQPW8E7Ejx24H2jhmk5ISqTrnZXvuPmvDsMK6IWVj9ltTq1d0
U2ORNtCG7iRnn0L45bkG5k45DLeUCNay1JiVn2acBjbsGE4bpKtT+4moeVs+SNBn
`protect END_PROTECTED
