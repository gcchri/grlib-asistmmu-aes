`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TSSecx+bVDP59kfowuprRW0oO0O5SurI0b+tnUgWTewfoYShoYPm7KbTmULLZ0Eh
YLDAH3+x/DACdTjgggk/zgOORlRZLd2jzywRAa4P2vk27IXW3D053qgy3vVM6oGz
zNYNHq3ZxY8f617LIcQ2wsuss7cb/Y9Jpol8Yx1gEhu0cdEnqhNtXjLibJvyhs48
iF7hv0uOP8L+EpGIb7hArRXeJPdquaNNhzu72V5mMKQU/zWHCrmIFoIo2+sxY8Ip
nIhJKBRdu2GhTO3BpyWKMAhIGGXqwS38gqDgYqIy1yY=
`protect END_PROTECTED
