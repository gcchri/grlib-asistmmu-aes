`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FN7hLIzUW6cu5Io9T1iHHKOZIrBTkPhd2wMpO2ujuRRjdWA8EqGKCvY2jX7jEFmz
MNmg1GLyl50M34SYRoUe4Q/RLea500ZvBXMUCzEx/0mAQjQdTuC6A9Zy8NloQgbr
qYobzDkMUfTztO+5HrcceOEuxs6AhPHuTjPCDBM6JcuXmbD95yqbJUn4UfXibXFB
lq89j3LhUHUtUufzWozlGTGf2polo5scCIvNnxWd1WPYo+upRxPh9ngoWCc4h8w8
N3MCKhZAySpk6KCG9P6uV2/D2RSek63CQXiPZBxlps3+HD3y3m+NuUubwPmipOSi
rY4/L1xuCf0Tc4RaMsE4Ivv+BiYXJa05oe5WVaC4UW0GiTv3a0AU+3zVjyhFy5Ky
DiDSnPGqTxhoQrLnJci6arYyCwDSkC8bdA1iM15DK43iw1d07LN9Op2erKvZcItT
YV3o3AZdU4D9jncGXI8sC0oYb4gze/ADKujKpJdl1r5VFazn3qWK+9MkOENeI6Gk
PsABBNXMVIADvJb1fEB/pgYD6kZTxfH81xaZptOnsq0JeTFWl1g5y/ed9KxkNf+K
0k2AooV9mRICnVLaEWP5VSADCDoQMJwpxQjVVYSK9NtF56vVqwwuIav3YvhPfdRw
NbVHbpCX9g/6fSk1pJUhAKdl0qDOY1tTW7lJIccs/FFa/GlGw9b4Mkm5QghNt83b
uukZxLy0FKzWvA/JNX9H9MOnAzefkoSliHIWhGEf1bwC/lbIh8H3pPsNqReDv5QC
oyIikHw41hDEgPvHpREpc+R+ah772CyluyqQ2FlOTwiwvA+FLhRQBtWdnTNU0qa4
+6poz0VGXDv38eUbX8tGefKTQw8Ta0r6+FYy9Y8qRRU0ztFUlUsgxW5HF/gvCnXq
B9PSzRXXXm/FKilqtuJ6Md9qRPAd7FQDQlNJzpsaRsZCrBVPQG9VmQwMZhZ4izN7
hE9WGqWt0EcP5Xd6OKYBDn4nC4q5Z7ozBo2oeOLj5otynRlPzeRegxuoJUUBnYZo
1Tn1YF8Ve40VYm0js0Rc4vZuIOLSq2bfO2YSvk24gxKLVycGjnf1+83QGKTRiX50
l0FOTQA8fBVyNm9h+f6OIWqko8D2kkiP8Ew4aqQ81ATdb7Sn2UBeOlRa5jyMG1iZ
mCM5b2mVcXGPzjeCCR63aWbuydx92YOYUirPvhoaYl0YDNuWyoDLqMEWvoaojW/i
qa2HlfLnlcKvl8xss/9MKKAUAecCDiBi4hfASlsiMVu9Gz5q8MhbMdmcS1AC+Q93
AgGvwCgx0hgYNtzHS0z5f19oxeIhPMqVwePTgAIofDIFkSvOl7JdmYfjo9zApJ4C
CKtiWbD1TpW3RmEouoPUrC9F5pZGRSyFvlu1vn1HK8MOa2nnY8JFiC27SOzFs/XK
SoLBKGfBnveOy9qxV4hZrW7hIIfZPcwdHTkR6jJNZAQugZOZH/Wl5u7DB9AnD8aL
JmUoNux6qTakyd03TWLxydDZ3xq4xmtlQhaDrcjVPO5YeOcJDRDTfO+/L3sAiOfl
lAbTGUH4U/IU6WZ2PMV42PLJB2zxGFJUhtd+OS/FSPpDnNyH/GutCVBxxTGOhF6p
OoRu0XhUTd1kMTpR8eFSeOcC+5oFMr2TlADFkPsucyIb22S+ptI06cfd8wUbyZtR
IHgC40SmKQNqMrorozV2LrQCj0JJvpJOA6GTrgikldRlozaWrG3a7xqIEYNhJsVY
PeIz6WAHFyITdrVJ5C+V6eLCMECPLUvaTBeOeZpoxEFPHm5tttyOWxxHeqPerk9T
ywJbBA2Uizc2pnWNCGUAChJnU5Rg+UhY2+/DDgXGzHexbpsqdlQn6vs9UD754atC
xk2+niodPTBAwOTPoA+jlqtZqZMgilv+XndLQR4UPB8Gd3CENR3MCZFsCHLht1LD
p06+7D29v5suoHEDMtw98JarMkruRo5zGIVOtrMfmhzregcFg9l7TGZ68y5SxVex
Uy3F3CQaPFr3kgihZGijQQCGJ76MLZ2WzKGEQNymcUI+ntU/B2Dv0j/zF/2wjQ5A
El8kO1thb/I1Cd3vvr4+0ymkaPXAWebimeBOUb0EYWQ=
`protect END_PROTECTED
