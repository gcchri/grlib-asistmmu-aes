`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ewT0kD9X/7TCkWcnvgRedwbszWI4wlBpp4jGB/qrTbjMp75Gl8+A8FcbGMnfYkkh
lnTgdp5nX34QCpcry5A+qUBXbD5Km/GbIYzj+TLIy5P+DCNHucKxOe8vgZzFAETK
S5eX9CDSEcfhWqNO6LNGCOwxgCnNMrFNj/G/4G/X+tL0nQ+H8JiiELTmg0cPPMc6
Lz3MD0R7PLCLTtvoBhMChMYlmY2i3SglBe4d9TxT/WFxtS9CPKVfv791fAZUG3TH
exogMFgNTFtjrxE0B3tcaS2XMTggl9kUS3ODp8DI1o2TsvqFe2rGYr/sVz5HqpTK
STH1IKd/DVOReUFdpEA5WTcpD61vGA+J2rh89BXA1ed5005qtj+iGocv6o/3D31i
n7ClOHob3ZjjNLqg/5erXiU1LvmOEjoLQbmIRyHeutzU867jyi7kjWkgfLHhn8Mt
L318c8jFKWcJf1TxjgRO2jGFjyNLf4DaCZ6jl67/hri8I7twOWIFm4mFe+P5i+nn
inQ7Khi0Us2mCDLcs7MATH6wZfyf/8akFGgOmpfgKjtPvZlGWO6rKJunFNBQe8L/
1j6pb7EoF2XxHD3wQlq93vrmkpbS071EALtDfhg2lhrAPm1LnaeM6gv30euViBcT
r5v9lt1PzX0P81IiXMoQmBQV1PF5WNTff/410ic+TUpaexNcsANlF1iRKbjnaTYN
/F8vXdNkbyu6bKc23Hh9u8dHnIUsjxrCqhAlFlXAI/NN3va/icYND/2gVUHpdV1/
DMeS9jlaHXwAVzLfmbHwFgPzsCfu4CSdwr3eGyFAi96OXbngbLPa/duEGAtMUJxb
0yo/nY0sDVBzpwk3/drhOjRmCXjDMGmPqWeJYF2I+JWGcoJ9nVcRBNTtBuGzahen
oZxRm4eyPhrhZD5wPp81gSlxPToR7rwaTYMK4c2u9++7DRVyPfUyH/tuHAmcySz+
y2p8V4tCKt5ADLP86Bu8rj5xw1kLsTN/GyO0HJfOrRzFnK8CIDBHM+g5r60rPj4v
M7oxHs5tSYuGIWYAWNAto6NniCfBXJoIG6jQ4TT3cNzyl3dSdu4X1JfOck+l47E1
tJ8prspcsaLuyjbXYn83dn5rEOBzuXuve9Xrr+dtYU6xk3JrSIfiN4eLgOVroPsS
BUhsY5irhNR8rNOUf3fHY0CYrm8kkOTqDlLvlBMFCTHp7lw5RDIc0Ln+oWl+xKDc
7pRj6fQeuPMMCf75o7Tw3ReX/4dqTbkNahYdIzU9LAFDEKVV1ODgpkqos659FX4B
uDc/uYpva7ohu82Pz76K6CNrHyHyIHeGldXabEGN+PyvovY06IiCI5THpPD5dBNS
hbhtscx3df3pdiFaOk1n08AzwMFBq99jDRgJg6z1UEgAxE+xz3WM6gAlVKlvQI74
LRKkRqh/hwaTzHDeE3CXPaDbEh3AopqsliM2VI1N8oDzAQQTBlZP6QLDb5yC3VIB
LFDKHKOUuDdvv1E0696rmRhr2gzogFDlmRfT8AgiZGu3tNP9UX02t/xT97VLKEmw
avJOgRTJU4Zl0wLFE9oh7mnS2rX+dX1hx2H/CuAtUIWF1TOUzLUYpFdRZlM3Kmme
FnBO5t72kLTXq5A3thD18rr/o84casny9PPULjH1jLXNy44mAyg1qVkjKUpAG8sw
9Cokpw9ALn1Q1PXVv4cc2BhqQlXDpcYPyHDSXrMJCH8KUu5d53yJU0yF0B24ECTH
c260SgbvQA54DyMXsCWKyDml5Fh32Kys3e6sCebxB2yN/FPDQ5rEAMQzF0vl1i8p
CYxKTQlW/gs6y6LfDT1JOOUbR3iKsXPSxP6cMM3FompmlhFduyBMuUXey7/KETkn
Np47fi5D63AfGQjW8rWZyzEE4OwF39ovaJbt1cbyHsYmwCg4QAENITZEPoBAqMzN
0h5ZM/PoE2L3E5aSxQTedezX8pzxjsPXY5wvJ5+27M5jymRY5abBZJPcQadjb9Qt
ob/traMZFpn43L6qF7ShNPZucFBwrTlDP/R1b8SQ9sQnKJuvEaOip0b1efmxHVjA
6nfKmN/u6kjkGTMJROvwPYZVTEaT4hjVQB33fxY6FyIytpUthmH1smvzYT6Fn1Hw
Q433ntwUJ6+b1TQkIRjgkXIhVYpLCqx9XBksqlcRzU3bZYfcOgaJYDtbQZoDnCW4
ZawlQnIEuqJBoFQT3Zx/qZAYWI5b4SuiFIJ15MWmdC4ssuM08LgetVOhBBMnrWOD
Eofwk8p7z9jls7LdUhraIdnL+ZL/H2SmuZGz9mP+6tuWttCkCvJRX1vF4/BxgrbV
MZCyfpDA471ejuTVu1Jxf51gUAisJycGf1BCu9ImV1qGiAtLnXm46Y1UQq91kdUy
H8W+FGdn5L3AN/7QfnTPHhioJnXkgsdF3HetmeFo3VQOWhjdWeFm8tLpvUhzKX5K
2JbMMymt6iU1OGP0YigPnv3LHpMsZEpQKd5becPJBFzbAf0p83MFyGR7Fjo4B05u
gbritewVETE4dWSr1buE89nGffh47IPIM50OG235eAda9lbooi/zNNtcFkFTNAii
h1JO1oYXot6zl1TPDEg3HnaVeH14ozRXtbjp/ydoKiDZdP8wVxECkUhv0vDFpFCE
PqP7RIn03IT0Rk+BYT4SXh7uzz28Dic7G9NrsgGrfbs+U0xMK8AJCnel7PW4stCk
VDNEL/pFdp86OyXqY3AX7/IyoliiJbtHBd+5htLiqlVRDtaRRXpRDdhGjuyUdOOu
GERADn7XIUCf8AWebVaw7kELG3LaCLX5uAst5KQYZ1M3IY6C3ONg54AQkggUoI+3
yMBos4gLLqzJx2bh/u98nmTCVLbBGv7PgqczPEIYsjR+AVL9U2gH+0m77Cp7yzC9
ejhUI7cV6kTocqLrHmykZKuWaSEYhXF+AipF82b1oEs9EhcqbQ0Fmgfh7Uoh2eib
Zz3UphzzmogHiET1El+FWrHtI487ASZV6pr2xTutRpcDQ+rQghILSbbxZjiXBsV+
6X0OUo/0TKUmEPXZg1jH8YmymZveZ/Gpv56iZNL7QCdHhCSXYuZ2TxKaZENtn7xJ
1zYrg6FiB1VTzCfCHHIjMroLtup6YAPOBinOXOrp+A0p50czP4W8VvKoAXs+DXgr
7dK9x+fGwCjt4fB0B+yvIAukX2+wDb8xl/UWB9DscyRY7xwdQIKo5QJQp0YXaPyH
4ZdCluaFE9f+pird9ThWsJX63rBMw7/fBXz07+RU2Qv+hhzGr2OmiLuQdz0z8DLX
4dwmph1OqNj4pF5hpJ/0BKJKJjq/aZzC5eWxdK1DdaGl4HkwULYBoXZZRpe+MpTG
c7sOS5Ajm/da9EZC9XYvfPT1cQT3spyDmA+hmpEA5JRs5rkqTkF9QodqQZtF3KCT
fPqFxQDkgJIv9w3WnmJtqRJ7Vthdrt2coX0jIt67JoQEdc/NEenTK4S1elcE95Cq
ojY5+vt1igj/cVFIpccABiz6PadFQ5OG/GzuOUcQHZQVsYMCSWJqhKqCtvPNKgi7
0BYvUTW9gKC4o0CLPwsjsspsDLYYoCuq4B1ZSA5FwMkZ+grKGpDyzhHORlYh5kiX
kF0eiupS5obnVw4PuVIgq3KsE3f2Jf8x+3Cqe9M2sUXH48rR1TglzIv4MNbterE/
fCWhsfFzV5MtEzOGYSGWn1M4+jET6f8PZVgBscWLPSNcnKtrriwiPoGiTIDDjYxZ
Pk62582lBtf2+/sCtOjUFLJi0Joe1qKk+Z1EMnuT+z7hoo0Xccf5D4BuWxO9Y7uY
dRMBxcwNSG7ECFvYJoSusBKPhf+/MvzxHHoKiQOTZDy0E6IXgj7aHycDJSWFn7MV
Dreb6h7IAvw8matB3LV5IHfnzanwJjL/QGStbOaMq0uYvbJHFq+PX8lUo0nIYOil
ZnSEXwYvx02rxUxKa5tiuJ9m7OXDnSdAQu1yFhhLqDxjwJgs12YDA9tJW6r30u1b
pxwYXU38Ii1PWUr25TPHgpuE2rLpL2ffJnAezf86gPCcAQxqqZlXO7zd8uY+HJ9l
Ghte2/HLleaqXGBB4M1VXjT48toS47SeJ8Z6QuX1OG2JxSj1MD64rKSbbFu6qify
g5LnQpDu3Ptzn5P9bZlzL4CIZL+l57GMTRwkrjDvv8YbU6tZp6PAMUTR8UkC9F50
0AmI/bNM4oiLM0LdLOPhlB9uJ+sz4xOVYm71JtkZ2rHgBb5pXLgxq663SBk0bx06
KbWkwHjrhvnw744Q0SYr2Vsq61VDc4pRpdOWIGhHpXUDvi//dtWZLrAqgy4pNYxH
CkqppZDrTx6UKyykDsYUIxPvVqsZqVV3qFQzIKfvdmCErOyTxgnjBtxWbq72X3gf
cFXCJuO2KpccQkSmyc+i04AmW3DRYOVF9VEdhU6s4izTTuVl6uWTtmJIISxGzOFt
ksWwkQ74vrN6hdNQj78SFBPjEbje9FBdtDPP4XAA+96ZtpO4TnlcDpyVoniT9LhW
vIeiO/Tn3GtK8ZhrnCJQ3C9iXdZk7SJls+7vw0jQ210Pk6/IClqsCYhtznbaPCKj
eR3LuHfdQHoBpyTCN/3NJxYkcrJw6x1yO9q/2ggJYsZk5iGbPHx5IRrGNPz9EBLg
QNOR6FOc+sIkW61fWSMpuo935PhVtxeYpmN2QVAMUJQHyDp4wFs9XyJfD7CZCiee
Uyd0CoeDg2miuz5Z4JQWR1RmBIEpCZNSUOx5xtGTrMxKnL2Ljed38DQYOVUWMed0
a2es0VAEKHWU4NsgeYx/tE7wjxsjJ8c9mE9GAyQTt+/0pAM1zWl44mjBax753k8F
kof1MB0brab3jclu4UOusodg8y7cdgaw75t1oKzdZUZfP/P6yY3RPjQ5KHSBGwOx
xg2ou5o5zDRqEjeIwjPUC0SJ+YI+9iQB5v5iNCRJ910X4XPzm82f+9BLbidYr54k
Og+uADsX3GFyPQVEv8Gtm64I9grheHh2hoK38nYFf3Uc4PXWFUcmGSZTEmcYRW64
SCgyiWv2DhmRnNDqvONHMJu22gvEyEIRakrs2nBfuoDMUfFReyrKTNu1bDNnASdm
B5EqYPEYk81m/sjXVb80vcFtZ9/OFj1bqF/EvRzWWCnv0/pb0jwtHFuMSem5HBBw
48CJvU+bw7tmseZjjrxmUViLZxVU7dhOP2qPyTK3OyKAka7w6vzt4wO8c/iqlpGS
BfxFfaS/frTT8DQJeayqejHySt8lYxj/aL6PlFXPDqphDWECiQox2CwDWFpx3vmx
DOTd4+93vQnqWXFx8JNfCBbWTGVBtcZUWqDrKto8UVYUPgd4zCK3BKMHD/mExRTV
GavX5yuDEiRWYWf4IJgO3KBxYpwaTamPU8XToMgQi33Xr97vpJEUClZvPRkbn4VZ
ycc+Un2bEtZOOl9uWo736KNcjCo4lY9dCOooQ7+UT6UUgU4kZU89LBDuxtUx4z4x
rkIWachdb2TH7HAdKfcCp95uZBqH8aSr6qIKOFeOaBMqwVJDQdG63iDiOQoWqAjl
g+/2qF9zD36MScATxoy0SmoARV6Y/hJFTFkn0zt1hXldNZnQv/LjiVPA4emfA9cA
e0HnogkEUVSwnc1FkNro95bR7bUcwzKxhUyu0GivIsuTtg97suOWBnoGO5BODuKa
2HPMuR+UV62YpoDsk/Wx1V0s+oENBJSJjR5hxMN+tS6WgKepHgkmbscjAv0zXt0i
aSJNAAVcR9tdXEFW+oT5RBFo+Kg3Yk/eNY4N3/zi8NvORWf7nu0Ii/T29D2ppWFE
Rg5yDFWL5iez84biZUCqyVox/QVIaO9s4FCZCl0sYqNuBodUkZpnKZFOXFudk8MC
A4YF84esRbLyghTeZgKcZwvyCFHdxMyfCmtm1iedjFxaOa4VXzklFnYFN+R9wSN/
rvYpx0Ju84D8pbMPSNQ6kCeCRA3tU0Efbg8FAKGshr42fJ7+2KxKpfuBSmzTpPGY
frZtrxB+E42tGSXmn9cKVHsxN37AevbslDCjgeYs+X9/vmliMXKfxfEzovIsq4fN
RwD4z0ZUNzvznF68Zp9bunJKHaATF7knBXMj3UPtaWbgcdMCjEoWBvpITKo9M7Bu
kN5rRKyDFPzKsCgvOyZJ6pRJXB0rwSnVsTb2yDfi0ZvGqwefQj3Z2MVZLtPuAQr6
kzhL4rfkLDRp69wLMwH7SdYYyk/mb/kFJA05AO30XPUQcFCvl/MCu8F9ZhPcgGjO
OpI8/UIeDy+dwx25BOd4ZMCJWmRQGdvM1hCIIzAntjg14fCZt8mA6AoclIVsNVKz
JfMOaaSgJUkcU2et3vSqh77yjliuh2MH1UGcq1dtt4i5+forPHGMB68+2S6zjh8K
XImFCgfNFVNpu6wTw31hokHsNYMVEPdB/GF7hI+oPfgaCGS43whfFxvOsFMmQnPa
mJwXxXQfGv1OpS8I4uXq1lNdiGWZYACscGvsnGzFbKdf0Ur7YyIIQfuMvulFaueB
84W1tp7lkFJTY0tbFdLzG16GZEZ+JWYCjM/wzpFDteuFMFuiqPExnLL4337MUDM6
ZbxpAXl4KdwvsH0J/+ZPIY99ZfF+6kZ9eHc3MwCfIKgnNwtgnsOnk12RBLIll877
+GrCKt4YeY26n+DAaLJfnArmACi2TLvohJNs15/mDBn9vID72cdekuJDAdC49G4G
fMqp+FH1/q4rIo7lTwt96I1gT03oB8Xjxb39d3vi94etncF8mnZ8292jr5DFeEJ5
SIsRiy31RGQUKMEwapj2yNhH8RuQB3fteTd72gjzPIJ/2aAIvLupRCZY7NVl6hVH
TPWIxYIdQL1O8Wf7qh2Bpr+/2VUQJa4GEM9Jjd6fyGlL97y6ZbSIDYreehV8Q2PO
m1MYTljjvpewkpFNDt9+eBRwEdHuGDbpuGpsqam+ETKeFJ7ON8qKrc1sbfyERDgq
SrJyQd5krutYQsYb+uwGdT73OxpGptKhj3rYxnB+49l6PAHc9gAQmpFdK1eelKQn
UPyhMUtpMluMq8tBNFhiKGDGLriMDxFuG+WkR8LvxQZe3nYP8PoORTeHh6NSgIDN
3/nO87V2cTX7qETjRhc+F+NSkV78pU08dTVzHaJsK0vu3U+VmnEB56i2Bg9HK/Fo
VzMbnCswtodCr+iY41qYn0YepGGmJS2+LhHn1yurSuvHz2mwVArW4R/zv/NdPf3h
Wjshh1sRGtLBpefG8f7HolD0YShSox7Ef+BvC+rGzXKuQBrWkYwC1lAilJrlSVtR
m9FUid4MnkPJ2mawf/tSWzdB/2nrKzh1cWRpE42GY+X2WGNy2m7ftP70QYUul5/w
chJvwLpWLu8bZFNcw0ACgAr7ZFo4Mhq0wJ5TNxAo3udLUGn3veeO72XJyiWXI/ke
IDGMO4LjMiNGNY5yj6lx9l/tPm9btHvOWq6Xg7/T3dbPFMP4m9bKWR3YxfhnpsLv
1CButfdi0CtG/HnkVAoYY67v8PmZHEhmonWQhFVxKCFHU8UdU/ojJIB2WVJtG79y
CmwQ8OCCzfcG1GIUiPQY4/G1Q06zNoTrcbncK4eltBZ8Md/eCCiwZeSN218xee/H
rOfkhwbGseYB7WYh4ugYkECKD+BibLDcjUaqZEar/cnwQc8ro2Y5pJhpyyOuG2UC
deVIJ37nOO2sQvTnV2Hxb5VrVJKNLtX3+rVR8YElAB133TYZL/eIcaoCdt6nf+6w
eeVcINtFe/1AsUFkaMXIQ4muqMUFYzE+nbBHMx+C9eLDZuETRRziJvDiGw9tOPXB
Ipn6+Ai3Kg1T4cAAZSp7d8qjwoKJR1dI8QcrHsO0KBavnQsOO71uNTsHzJuppo5p
ulwqBKD4EOW8szPC0rC4qOxrUaPF9Tn8aK87Hjs1fRBVkZO4XKjJkPcDj85YoP8T
QqKG/So2bIdE5YU9b7v0BOL0FgUoaP4939XeCw6/WAeFhqB+K3DQaw6A4XKsANSi
sqhmh2u/qZJ6q30Ik9qMrtfAWRmghm0jdBw4A+cUt1AouYmU7sBXmMg0+VSHZ50e
7sWSSrSVdLlad6d59b8nJpSm82dtNz3Wo0dc/l9Qb6WqmkCLmSzm7OQFRL5FBT5Z
9EfR7e7yKGnA7+tfZuOAKH/SYgfZdC5voty/n0F26eo=
`protect END_PROTECTED
