`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E/HiXp9PqkzOwIYPMz5EAz70uSJJwo3uXwESYOZZhW0ZZj84kYbdpHsM+3Rzdsl+
Cj4Ie7NpmYIgvG61bXd/RE6iSHTidB2IaLJk8ScyWWOCC3jtIe1VbEWit4/vjKzE
bp1PE0i3FXBicLZBbOaxtdcbbc85fyIkuE94bxmOVQWT/UmMRDJpa14Kx/AtBwo6
XrMzMfqBFkSZuEUN7yzOsnxktWnJSeQdzp2gKiFTRJh+tTQzms1eNanL1IoTEzVD
dKEOlkWU+WvZG5Zi87DDUdj1aiqbaPoDzWT09U8aB9+10c5cvM9LWuQ91x4TzpnM
/fYhD2PqqWqZFszxuXb+s5id3AKpDaTcsezVg72bjLINnbsxsurbL77D39cdCIyS
+tnZp9EwhhjYmRDejNd+FZtYTOs/KAuZMU6NVFGWD5wegQBBqRo9QFVpT2tc6OO5
FBLCONcZFbxvA64397x6wg==
`protect END_PROTECTED
