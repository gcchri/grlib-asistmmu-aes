`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZnZmp6e3/kJdEKiGxEPM4MwXjF6aBtGkDwSv6aNweI3Qoz5vTiJCgrEJQlsm7I2k
5fyUW2jNisu72CUB1U+QG1iTeffjfVPoKDb91rupRzB8lyScjFbASAxXENGwmC9/
vJRX8h13DmrivHrKXSC+xKmFNrsIMcS20td1s82PCIklhkI27xqGeFUiwOvkL96O
+OKJpKSLx6K2kkwyMSiTQq2HDe+hTeNfkEpenhzzueEWNf9SMht4QfJMg//Fdf5Z
aYhd9sw619K3bpNw92AuCaar9tRjucQ6PLDW66pvyIT/MmAFmrvS6GEV34RIDQRx
PYNfBRch5B8CaEnKeOqsPw==
`protect END_PROTECTED
