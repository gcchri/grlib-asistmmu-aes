`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+hSn/MXctpZPDCxGXXSI0mByxzZfxnnN+GiW/j7Yr28iD8UmpcN/tQDSLsl+QLUX
ibQBK4M8C2DvRVR3LekeeM0tCa0u09eEQiqg4djf8X0slmwNErcFxpw8DFmXOOi6
U9gfLo2xJ9zRrXbWVRdjWeHYW8iaTj9li/hDl6dMtm+eraroXT5GXYjQrXcg4GuE
hPv3qKe/KrkqLFm4+MV92eG1GzBQlJyJ/We/+3rZQ4gASaAw1Ny7wNiDf2EvLp44
e/Lzhg73sALCqbZjWbobegNmgBFwo7bcjd/H6L7e4Lhk7C2rbSMJzVbSNPR4UJaR
GXxAw+uYBeP4N6JPvaGFSg==
`protect END_PROTECTED
