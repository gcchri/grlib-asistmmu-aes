`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+lcFB9qgzOnF6R+82NLq0CmXynLLSi8vAF7FEgQwI7sRWF96Isp8geaYG44gvX+j
Ql+G1pM0dRWN4iPHSwmXmDR20I5QqoCye3/0YrnDIdilACLlpC1OfNoSm03Q/F8G
//oPZMB0x4/vn4lcIn9g32dVqAb3k3yxah+cSPV1M93yyWkg+F/wcNKhzgOIHwsc
43b9+CGp7F/T3IoEAIrAPT9aK/HhP5J98O0M0BtAuQmHmAjN7jLRgtf57lGTrDsh
kyrCQxG4QB/V3XA3Hm0nt0esyAT3IEFIoQR20nbTx8ezO3UBk22HLjsOhXpeYaOm
zPeNnasSQDVDgxzGa4Mh8WeVr7LGNnvIFUqKL8HwwW5bGnos6vtwnIpF9Fe8yRD/
G/oQA+R3TtcWSDXsgryU7/XnT7PNmfGIWCqBV4SARNsiUvXggYdRx3Mh5u+Ic2P+
wVY+6e7RdK3U9yXeH+ZesB1tu2a/S1hjGVJi5MRXdFrP9yJB6yaFe2KGrnXkmN9U
d7pbnI5/e+4GpcZiJBlIZbrDTyCyRdM5DeCTGYoemE2BisiKFtPvgbA2fsIfar5M
NKrcmV9q0lCmnLFeq6avYoSy45/6lx+mYzW2aoRF1AuH7PV8rHSDM4tgz+Mhl5dm
foIFM5j1qX09th1WgVVFnjrewh76g5kJ8UTewX6kdDZzhfaxmsfw56OkdPoC7wFu
mUYfCKeNtqXy5zfrQ2PxSHXwyEWrHUvwllBLkC+s/OWE+odGQkMIEcduMRuRYmZb
L22fGbq1MMOETpm7IJlSWVdRE6XyJmEYmcdGtsfMZk2rbP/gtJV7wIGW87SA7qaW
FQSUEAZmgpmFslPOOe/RqfLJU4a3L5WmoDbQtMDE+6zP6yJY+d0K99PmU00B5UU6
jBpmA/0pjpyYauT2kDrqbEDhdos2MTNjv/S7bD132Ljjv8fnIdATaelDAGiqmtII
eILxnoDm8GihmKuvEKZktQ5unta7bJt3gh4brGEou3CPi9lPg8SNwtlvjzTgv0X5
VrSg8FjEV6LXWgLZP+S57x1HTA5zBc5aWcaq3xd4O78uG8NSY4lXjxRpti8pRSVF
GLwTamx+bQtoTzQoxFlzSIeEJLb2vGDphaNZS9cWLOaKcwh1qF7Av0D5z/nAavUo
uO5zl9N3zOjT3T6bDzsklwxu4zPfdLdF1cumMHzYp2qslZdTlffPYMVnJj65k/Cg
x3isG+DxH4LXm6kxYnbgSe7L9C6DK8lRW3YC6N82rLSoD/0fuH87plUq/0qLDpEF
lt9bjTlFUkZtbr+/wdfhczN1NS59YYkoDBqRGO4xoOmYvMBcCk5fcq70NASq4z4G
yJDprDvFKv5asfTqFyfDMYqZGsD1yjesnAg+w0ZUDngExzY0vljy0j7PKKbk5yZL
HCfRrmcOODhBuaei1tdXwewMD0aEXoKeh5q/8sNo6s7c4DKVtowmP1HG6uFt4mSF
AEAVfIPW7sdR3REPc7mEAwaQi/ohZ1MFyOfdYJ02IM0URLiZKHnaGN3GbGEi+5fU
4XSpcgsadsGQqmuD1N3SyZJDmQe5aSg6cEanl6wkHw0hQHVONhmaNkYx+rr0mVcI
XjEGnRZykGolwvOVvpDY8zZby/XwRkLByXIxRlEgCaY8f8TzNK2zZbeHhsMXFszd
BqzfStkLEoTPYqCxP8X28mEi5LxnsfJgeh0ZVRxyeM1oqprpe43aGxN5AJm+u+QU
wyWCVkiml592sXBmiW7hUOMWzwK96RjPh+kFhatW/Y1zPy6EnexHeqUsgLHiI2PS
dwl8CW2qPL8BrmPOfOm2LYYkZark2k6n62LvGYIv6n7Imm+EljiLUc4B97QOM4mb
T6BR/mVRA4RVQUEFzTVzWpcFsQwEaZkrX9opP+WrMFdr/e/ce6MJ3o56EH2kvO5b
+5LabuXG1nuOhaF05B+hi4liDEqM4UaNrigI5VME7a20TvsoZ9OnYpOr4kTLiqeB
vLX3N45zx9dHof0fOuZMEXB12Tt0iCnbsvzMponiJgf9xyXLSSKWC/+sm7C1Et1e
OIgQsiBm7mGmUClS31TW0rVGoAAbGZ8Qr+rtjJQT1Yffg7JkCjSF83CbbOd0LIv1
IeoqcO/nGhiwGCgEk/hSIdxE+A0tNwk6zpBIQIfPoSa+cTjWZGMoJVGuxPdscnvZ
58BxM9M/3hhVQCnS08PSQvTbYmCviBdeABeou2u7gOBRBgG2h8qYTW653neLQglT
XH9kWnfpvqj/hp7vqUKo83hQX2WpoEWJ/52W7MJn7KzQUHZ6Up71Giq2z9R7M6+L
7UF90DQs7pisD7s2UsWPFiErPD0E2+xUaivEJPgf5ViO26qTVleGZJ3Xthqfeubq
VhNotwcNMc6jiBnkOuhPJz26PqGDqnkRQH3Xd+T7fUzCT2nxPdQqK6AKDS7ElwT9
+86ipDb2xNNagpJwnsrLfSHI/In06LdRmZLFBiznVHVQRMr/6m/APh6ymWJKylEd
1dPBF/5SCU1UKvu9Y48FX/i9PceGq/Za0ETGnO+3b16xbv1393Xn/g0CR26SMwKF
wEMroR93HVZP4w+cevR2WG29yYLxN+ovxeBxDuPwB+QZ3I897cNFUXUvE4PnjOm9
RxBHFMmh2UiNJ661eJpZMj1+veYL6upZ8aabHkc1z1rCdcD2YOIpBeEB7eHfNrIi
EsQGPpgVUvaHscUrSolOipnNvCneGvrJmh14MKWPXeP4mh7biWQ8HLZ4nvxa/0wq
A/4g0NqnBrohHoo7oIaLKgWJboRGP6/szEpvp1H9I8t0w4xQeitg1708CcOh3B81
PlpMko7EgMvop2aNT+CyH8D3vcBt697/F5zHB/H6LXUl2Vcp/R1XDOi7I4mhT4dS
PO8o5MglIMKGCI3Ous1g+/Q0ObVxA6FVkxrgm52eNasnSUWmgWsUd+ePLNJ20xNS
BwMy0eh7itHQdEm3JNO4om3TgWLSHhv5QcJXsLo2HAKIm8ebVN5aS0ae43OyCRhr
a4lIE76satq4BtcY8qO0YgP672zj8ex7nOiVPOxdkvx431p3mUcbiznNtZE69IKx
z4QKYb2MVvYZnn5Payec0HSHMLT5RkQzE5hJd8NytgIN3WeXa8DEusNx/pkEfXCu
dW/1tXaCjiuYo4Ly/+dXP0nb9OWopnEsen0zajMr1geF1cwvjpUsTL54TUTSkf7s
Xk8R39IiPCi3pIdhquua97jQhPHgSplIKZkv1Hm+qZCHF/TADt19ePA0c7eBXACw
YlLtaB6gGJSJQnCsfiXPP/md3aaha8QPwcIgJAmyU175xx8lKcTpFCdazeOznHel
NAsskup7V3SqRLicCs5fYkSQFSWfoG9qfrWhd3UcYYF+c4EAkFEybomiFnmSkOoW
ECCaaJoOX+gND4+z9HFLTIJuDZSuDGiLk0oDzmVbvXLKeSyfBctpCxnKQ8Hmtc+C
l3hspolLNz1lF1meN82giKlS/gjQPWsLGf0qX8B3kdBljBZSEC7vJmDG/d1mrRz6
ecX4mCcWbd+cbiRhR/yK/qorOPkRPxbY/qDg9Od1WhuuUKkw0L8m9LzAWuwNZEq1
FrztBGp9epBeXfCdQJXPRh2lhAVtD7i3BvAOaAQYGMauJXI1QBJVRCRHmfvXYWWR
YU2NsjkVbWOC1MFi48v+0rFVxVUKBs+7egLkRGMsSsILG+NxwyKgx4IECBRbbCpY
8KHnQ3nejCHfRfH3DhnOVH5GP65L+0CdGxT2NDenknuGzpJ4ZawEr0PK15LUSP2O
xN9W6FKlJG6WM+e5kbALNKyWXvJZECDeUx3andpRAfijEqJQOOYt9E1yIHohugnd
k3SuTV7WgmiZPUFt5AwS8ngKAMQU33ZbLrWqUjAHfBqiA7aBmiowo4kxesMXbwR6
0pWBKgYf5PwgnR57km5pjmHvVv98W9o2C0taEjcsA4W2CPjAWGYk9P9UtkuAdU2P
asK272u0uK+/+TImRnv1qPYrcNYO5OiyYENoArUnN4X4dcOicx92jO8kYQPyWA3k
zT55Zr9RsGIhWkYToA2IZmrrhMVLh3L4hz82Rt+Qj4SQ4R02nDC6PgOGCmyTbRgh
EQzQnIek2QPI7HJpp9mT/VrFBHU1Pwrwq2xjB9Lpw4Z3aBke8f49HpfOeMqg8BW3
/h5NVOzmHLmtwXL3Jw77EIo3nH5RWg2Nz09qu5irPV3e2UayAGwGLJlI7sU9HwSw
luUBLejk4hZ4ijhDE7OsKsT/D/iRNv4lrAmvfHcQv2K/4VA2QIaKe47lvVGSLYI9
ddZHqL7nQcsYx29yzoRxbxftCDJ9LWNPn+F81BoUCle+HVRjMnoptz/yc6Iq1d55
MU62MHM3K21XLd55BR7ri6orS+5DmEkeNeHjoAN3HoviI6Vop7oB2EGolR/VyVWG
JjAkXJnYB+ozjYJ99+fqQoYsOys1lcST05UY4/cJzg2cDuugrFchgCMjaP53yPK8
nR/4E3Q/l5PvcLc2ZdZ246x6hXVYHG126nLVcvBhRf09+mo17T2QB2M+N6X0uOFZ
R4C1Oa7ILpkjtZCDFI6hjv3vnJLKmya3Gtv0m5Rfk39jGOehU8R8aqkM4IdTUn9f
E2S3l17vtuQ2WSLmLt5zekII6231F2lcxHPd28tYM4s7G9NMkmSmCPzW/N+ILFNS
6+Nd5tyiG7s0PbmMLWFuBRdxfAVE/ZlqjZjx5yZFKyN8JRJApAYn7RB/7y+GSat0
ruhgVw3oHXcDQds96aye1k/wed86MJ50OQk+c1+E6+swmBgOtpOuOdS3X0qbIfqG
uAx8whVWPo2CW/HTuR3dumtWxXx+MvqotMqPTZreDTExC4W4+hDpTViTFm5p7mbs
UKYrV/f+F0IlBuhuPt+/IaQ28HdBGoxUA7nhqozJlRLAdTO1KhLtoYuyVGKOWOn0
oEzDxd4E1BhyPQh/Hxi4BfMw9CF8U3Qs+NMKt7S4CyXTzAq7CfuHFSZig95p2tFj
670/ALwmdWju7CpSP021yODrthjQzlizhrKr7Ci9yBtDD5FrvDjnzYDSwFi3JCQF
p8Q0WYVbUrsttYBtpXfX9m0USnKhXBUOFAijwFlKSuIJhpeL2Kr9HqoXO6Xd2o9i
s66gzSTEO81TWnvOlFEX2j7QvvpLkdrjsva3UhEpS5SkxAo8w6txcECz2jBjMlhh
s9NtlOwfRNcj7gQHgQXaHtwMCL43j7nVqwyGbLhT31nLQln1+J5l6e372UiVyFzc
2Iensc52ZCrwV0YAr7auNEbcpZbcwq0iRwRDKC4T9jIM9LdfBMDhQAUxcg45XyiD
l2O6PjFf8EzfSSQM9YcVxXvEx9MRA5GsqaV0yCqyGhUSHc2wsOcyenIHiWjV06ZZ
qaNyFvl0ZSzVD5xkBZ70JLD8rx9pF4ariLs+4pVONjj98efx9P+MEmFPls8qWGDW
/veDSUCIE4A0PiG38GaJslanGC/H49ZwJsJFBXX9rsEq6YYj8GdphO6qTxyWEJ+O
cVKD11jQPoNzZuyL/GtyM9ZvxoukY5YEIMh7lP6YlMqxI0OHBkGwvPfjJTz/SGlC
z5mpZMrxEnsqRABU8WotsYWtIpj7539LWtEL04rVMcXXo55p6FUn9gRTEvCrbRtq
9EjO9UrPtI34eEhwVE4nH4DCd7UdGLY7/4/7BNR2fys0CwA7j8HF9TzO1023UKJc
H/+Uh/Tp7FfFu2fJMMTEzKpqEpaqmUx/7HIPivPK2bsW0LTM9HqQo7yjilAP3TNW
AI6o52RsrvcQ/ZQKqvNrBEkVTJSX1RHk2SXa0j/YbfLbNYI6K9av6M0xy3C6eK5/
mS8ZUQ0rZ3iT6YyG/sB0F8l6015srOUmfLPSCXvl3m4nqv1FtbSlvSCHUk9LBR+j
1kFPXzplAKOFlpNEGVGs1MqCLqzpBLHqEkGF1tNc1x9pmAyQL5eUurzO+ZljHTTX
JF8lgXC6j3YPESjvp9fFLEGDiTKEA9LLRXKTaeFzQ5HilradqZFJcJaGBFNNSSur
2vlIKcIkC+y/kNu5akn9f0x8xXDKtGOm01I1BBieOt5hhY3jJdzYdgSLoT83EHwh
kWGVnW6HP/+AW/Hr65JwxJYuMrfOKe/GzS1PXgkZbGPmqUT2VssmtYTxyQ60WEwZ
kD7i2WPVzyknv9I0EMNjzqyazbRSCslGirmkSC6S9tta9LsuPaIsR7ap4kA51d4h
TrDeXDRlNpj2kBMc3ZXobwkUNg7XrnOqTzBE5WmYyoVfErzBT6WQlFonCI/7w9m8
XsrI+B/dHPrZEY3L/Nulsnqaa4UXKi+nzcibQ5yMEdM6+dlg2s7gVMqSbh6BVWcX
Fr6MQoENeZpVhT4XKWKqT8tHA/jFCdZubTyebHljGNI9y/FIKhYb+CUr/DEy374z
22hAq2Jk613xfhg34LFVzDwEeyBVmDJpvfal/qapZ0urTRDJxzD3hSordh9urgIG
HQ8sRBE/YXOsOgyBoFViaMaKPI+LmTKbbiacr+tYVHGz5Kb/G9Ebp4WZ9OlYRsEh
H7e/2GJcqoKoeoJGQirAfX+QU/B2f7cS0Cl/atEhPq4c7Nx5befY88uCfbe6iv0M
vX6oQ9Bgw+jlLxhPFCOgTTvehl5nBxdSlXN7aKSyH9EAWwFnEGnzI4A1Zkg0ctdq
83TlMUrL67IMHL6t77Z5nf7WTd8RU4DnHdBZqruURnoQL7l1ZyNNVJAHgAfmEFLo
SZl1597Ur0Q3zDn8LZrScUtvu5j8LriEu0q1fvplGdcXbkXrgwK81xkOujtYGcpE
ZEIoZ62ZYJEvIEM3EZBd3FapkO4wGn56jnF/4X9C4uvl0ZwgW6OyVVIPRZymx84u
S2IVvPl2Z/7AgWF5m01sgwQMFhzVO1OhlFK1gQzLJinvKs/JkvydOQJ2d0elR/Gk
I3QGW/HKCA9PeHmnlHDimKEb2rykQFXfmOH0SV3f5t3LtWPDp4URAwZUuMwG63pJ
sG/FJCzhfHVqyvd8TVpZi2yEurKhjSx/KqyFHoTqEbukj22j0hsiXSeK8NTtMI+d
8/rIj8Pd2dE0RLtaUOHfXWry9NHp1nERuz85M9OqdnPSRKjDqnc0FTip5tYsYq5/
U4BIwozZzftzavQS3WMpWwiqT4csh+Ox1SEcbEoGPG+PLtNezCJvPyxQxmcJOMhU
plA2Gdk7gECE0J3nITAtzfPk3zJfd+cGXA2mRvJ0Zem2hLk2SK2r3FZqk033OIbi
aXWaodEyyPtcwdzvYFehFNvdQfnBE1B8opP2vDPgiad7dBZEEMZHueqv1Ra4wJl9
7/Qo0jewOCUddUqeF9FLqRcYFSMEkO142UpnAeaSQGuYL1ssI8YM3kyc9op2JdeF
0EjHCAZcKKWRW7/nn9ib2U5tQJG1er33fYjNTWcwEkgkuUfG89G0q/xWNqQZay+O
u2asd9DQ6rqkXzLfXJnIcNWE1MFqipJ8jlHfxjbMPlDJZpPYUQBGA8kM1p1/AWl5
bs8dHBIv388UzwHOvRxaCJDa8e+6cIEtRDy0GW6xQ3KdOTT9QT7XpVjH6SZrE3gp
9qoBuqYoCeg1HI/BM+xAI1WvBoiZ8zxm0AZrV37j0XIyLXJsVcxM4TDT67wSEZdc
njYAGqQ5He9uPCrSEjw6GsPABLxsNMqJaYFv7yrVYb3MDsbUH1vL4m8YaqD3lM3T
NRdksLs8khoEVjzP3rPiaa4tvmrJRvtZsAP+mIIcH9RFnhwZVaMtdk3Mg33EvLa7
fH/TquNalxFW804278M62sCYjnBgdu69x9zINP9kJzSxp4vYhrrvR2+UPwg8hQb3
AU0xWhtDKcfRfq5E5dm53xh9Ym3MY6hTRd2iFhiBaVVplYVGv3uq9EXwziHZKoWQ
cq6t3iWHKdSCPBQ1CVm1AxCHU1Lh0I1BgvELCRDblW9fOu+UD1AkguZe5FAZB5BV
dST/IE/LCWD17xCpLiHaE7noGswRPzf1bng6HPhaEGEs3WwxViNd07wdyfaCK3SD
0KCygWPO/+3XZP3L5ws20rIb7QXeh1SxJlznpC6yPuEfiRzEeHqgwJo3GTSOon8S
VrIGac0DmDy/8j2psv3aqSG1PSATwBwW8CzCyD9OG31FM7JSZDriCjoTcJB32SNX
syGFq381yetU5OAMI+ZZM6Ngh43DQXr7b06veU5KCKfKaXlEWAVd6DwAoL4t73HP
oBCFh2mxhrSmc82/vipxy7zYVNCey2j5ta6llaBcnnp42vHb4EjW9DiUM7FYclv6
KUGw5FiSS6v+eK4glhpO5s1OsOyJpMrdH1YvKiMxF2SvzVIUUeE9StBQLpg/whUJ
okQh/qnw6eDOM7UTVnHj3SOubhRieGTvbc8EBDkXUUJMeTKuEeCfp7BgIui1Xdpw
/B+08xoNs889kIuMwc1DyCNS+ezJJJYdUMTlnRjN4JeDUkpvCx7brTFaDMc6SxZm
v9QnbGNR3ZeILFHZsdjbBS1A+jjBqcmjw9WWJ1tBR/IqU/GA2wEGR3IEVoUCx+JW
IH5E1azPU0hnjG7YsjhDdBr+TWFxIT3drY5DKT/0a8ZQMTvmnuGz+ZGs4RiUieQ/
F1MPzenG0BiH6sSzq+OW6i2m8fO+/OPcWwYiMAKS61Mw3CMSg5rpYlt4RE67ZYDY
RxG4UExr3Ec8p7SSIgyBqwwIUDEAt5V0LA7ssSsu0jy5SU1P75sDaLc+ZNk1T0cB
TEGFjnn/miZ/WELlOsqpg5/IwPoODqjm2jlM3+mGdR6+MOeVcqvsTSOMxcsgpYAW
DP7kpFfJlOJXWlaJEn3rvtDuKwubgeD950qGgs26Tyr9VuqQTSR+0cKy+9/V14XG
amd7Rt4LfS4rDcHqRD8scpy8eBBaQu8nbnyBPtzOMDOerJtZDrBCCH53cm0DbwmB
HI6eVtlqrNBZGbxegmxPE+u303DmhziQyfpjx/f+8VEvDP9+O7aCssDZqFUJTDLU
vegtwTZYo2cbmXKC41+2EH77/KXqADV2IhBCpW48u0DTFts/m0EympG9qxYDWM25
VhrjSSDoaddtzx4bRy93CzEyMWb4dwkd/2DD+FrJgnDTviwXKh9dMz1FFnsBvEEe
S6FNunWAFMaabHo5XuA+EiWvLF9SFiG3elfR3cZFRNl83ABE04X6ovBa3hSXmRCS
ydeH3nLSJicz23Pe3POULIiIJMGkLgQ7ZNwwpJY1miQenFm5LHswqXsrJYgoyJXd
+90oxnGZEgFM9ZV/0kJRK6ju9PHJ86HA2nynUhLeLdsPEG/Ikfz4bi+JMG+dJD9/
Pf9SpDceh2krm4nVPkzgXZyhwpK5+p26jloYyXIad9ii/Du8DeDPYpB5rLpMQpiV
tmWzLkh0I8NsqX5xtVioJwI+LXABXgPPQE6UAH3Gz6HYMTcA3N7Np3apOV+d0sJ9
E+qTzWZv49yTnwPTsLT2glL5puqnwYqqeCGWAtyjCjXYSFeAAw1PVR8tJqenm+DU
NA4wpVAp+X4pkUHhuY+RYzeB2t0hN9k/vEYKfREI2WTZAwayixRpzXGQ8BlKH1xy
EC9EP/2iQZKC8RKhJ7zhln0GNzrtfHKpkE3N0hCi5qH8I1DGOrFGjvp3ZGCY9mFO
bW7hw/MCMLPh0q+zg0ocn9c30VephpZH+PqHAddw6ah7NgCL3iuN5ouzrBmq+7f0
/cgJ0ZZXT19KsEnjNNCcVbOONdyMoqmKXdU56n8cqivlh1NEtbBKnIpN4fZCRqKa
pL/DFNa0yoomUS/T7GzXr5g3cSp8T8Zqt30VW4uque14Uj13tb4zvFPSq93Hn15K
QPjh/3t4i08EeYF4OHPO3Pq5UJ0K2+gJFcIrWHiKIIiIKJZ5gslc4NKHT4707SWl
o0j2Yb/EwmlQZIfKKNdRdlQ/jPPFih9FGJMxTTrFALcDHuu9SyTYQGGIFGJiTlb8
Ei2Z8lt4vfMe6Y7y4ELgnguF0MIpBur002lGhedxWIt6h2s94KfuyhjaqaPKc3kb
g72zs0s7x4Zl+e1Z7TFnpRER4OhApH8BAM2JMbs7CMKg7xQxiwj0Ad0oTaH1j+M/
+kly0FOO9t2L5H5rE924Amk5DIQdIjxCCwoUVQf5LbVwqe5wyDc8YDjqcRKeuiKj
Myj0+o02uHnpzf0I7xpq05mn7Q5d6c9YIctYzR86PljwmJX5najE7UxPQHtSCdit
mssN9qhUDju8ICBqo9OcgdHkAj0fzUwYSrLzW5YTTtUo5xe9mUSRb+pb8b/XZ1PQ
ptLYhyPUIwosrxulb26TC40rAmg/WtvPEgJofOxveJ3DdCPmipnLE+BVSwWKRI4q
qbyxDAUNzxpaX0Y72e5EboQl9kRWYAASA7oNhvcGzMoBZpgusVCoAnNUa2Uvjvt+
Y94o+MU/uS0yYT55twI6j/FFZqDIKX50VjDNUEtQchHckOYuyBcDeD5eC+by5kbO
tx9Km9teLP+HBe1McogiwNWYJ9l+oQSnvLe3xUo1O62FlYKGxKekKV7WzD33+ScG
GcyqS/I02tDK42peJzdV/ly3wxPdDTplt1z+kSpRPTeR39HPXAjWloRYmlik5kE9
ZP39NEHqyIRbIJ7JaG7G+nj/hWY8/S//BmbtK1/C60xdAgcB8jieVaoTPErvyHsr
vQ++NkE8yCpqNzyqU5Y6THg/Pig97k0jJ1i2azv17HFoy2/65GkSChnoGJ59poAM
wqIwNKG/8kl4kaW8HffAY4sNecnBb9BzFzBR6QOmJHGDi+E8Zmkg543z2G5zu7t9
MXe5jtOKZ7simq+bhgeyja00etA1m49s6A9a5wO8mZp//zbqOITIooUzdq4ODxFz
zugIo7iknz9motWznpC3aQ1kdNZC91zmF9Ltvpr2pGw4SoRKD49TrYLJMyvj6ze2
0+r9LS8PYg3nexxlWxf7D8twGTQlbzbkaa9r1tYYnqXYG532M/mi5fu2WaCuXH4k
oZ4+Vlwt43dQynUfLlCTHTIKxQQFSD3lKxwSOGFyr4e9FjKki/Od6MK8YAy+scgK
4Ng5YHayUmTKDoWHnnXIaanHuV7glohjp2pA0kxp6+xTrTtNsNXwyWHbGsrzQKtN
fFkbRwwPX2n14nT4kAi6Ty4qUeDe+e+J2iZ+OqBXmnzoe6ljs6hN3/ueGAmFuFrD
r4PUyQ7U+sQafKcRJ8hBrqhMnKubKJqzPQVpuwxWSaZkXv0z4rycOGXVGhT9w2MJ
7u8RsYCmyNguWoeUQEkxjbz0/bJiXyh9WyX27f1pRLO+JG9LtgGoLiO8VpiY/lwf
2MPGLPO8yO7hbJO6UaDQGFsMdjaYVdt7FD2aJzTR57ajsYUhxQUOtuPksHsJx42a
1ijPYrjKFTftm779ofJtmLuQr2BRhP7ij+GT4glaBlZeHRV3j1neRWIvMjM3JZUY
/yKH9voG29MHcFVktklOEv7fxWXiDl/LYXz5mlUXPpEcqG3MK70VgONSoP5r/WHu
NI3nRe9/0YPX0GRbWt0U6dVRHNdUa9TeH7s107IeImXTZWdPYnYnXRAcSZEvRG7U
Zg1SxuJB2lKKTmF/YDKKLzFvMViGI7/2zHRoRsgpi9tQvA4dMeByW30qhInlQSyT
pw78cxIolSDJYoV/i2PkLQqvnUA0Lk2MmiZAn1/IPumR4jQmZbWQbbl/kbOoXNpd
3YL4YEElKnIMx5HZDSePEMeQW2SEFv6rV60WZW8h0JLI5IWSxUo4EzIDEk8F5CPa
SdVC/WMiabZUomtBC+hUzKTQcfGMvDLi0PJH8SmUTt5TSkrxiCvVhD6/6k4W52XT
W5HAIkpz9au8lNIvRdZ4I/SWX9ln335TCfSjfrT/qBg3Wxh9o5Ba/0Xao2XTH1DZ
7v+VMicUpsF5KTeVLKHfIibwZcXOvWNQKhnY/qXxsOvrdLVg1ZfwC6LGLhHpmE/8
XZy7t5EfJkIOS2GvZ+i+lAmKpg6UhCkY+itjTs/jJrRw1ns5zT9DDXhXu4Rv8pI4
RGlzqEGBOiAfz1BEg4Y17PflNxWAJtWEXgZZwgYWCHqx9YFrInVUCLVOV9BphKQN
4KZuxW3cDU4rmeDe/Fj20S9wwhIHjvSd0Zi/gqYqUJ1c4odjCWwcYRKgJKLCvNlp
deblhxOq5J656jLiuKEKm3KGFwIm3sGnajerRhjA5gDebuJ0OVYvSf6ezO1zIG0K
O3ZizIdpC2XQOozqNfuyeHEGtaWG1tOi71nqKEYs4gewHWXx4Xd9zNS2nzoWqCCK
f+pWUYcqVguiAmSa/us91N0CoTVXjpWcRrcoAfQ797v2Yq+HK6QPL9VUbr5oxJS5
oTVkeNxMeWNvpxzVZoRx6S1flIIazyfZ+orpFmCtAO5pfLH1I+uS2pOjIcE0ndWT
yj7hVsM07MQr1nniamgU5tFh3MHf0BKQ0hYWPcRqoI11ZQKc/UWX3cZZinp/MIcH
3XkPr/xddLE5FVrBL9XMrlFbcdvcz+0HgZvj1rANelzVTb0Rff5o7fbx1s9ngh0m
NjDF3by2dqacgnaaHdnJukQMZaBabawwBLAoOeiBOYuQ7paYN+ZQObVO/0S7RAUU
Gki8e41e0RYD9+UdOH4+VfLqmiwmm3rKISFgogeJbHuVtjJOa1rTsJlU3Qtwpg9U
+04ddcnoK3F01V4yCvJxr/POv7k6v8cMZiLNM4QzMpHvaMNk8xk6FbTk01NlvNaN
pAV/Yp4S3TqILXUVM5oLplGqGuj0riZJSSMYsaw2OEnpXU46VEMDzXRagbQyQu/f
xZA0sk8IMOth9cr7rp96lP+0LHjEmYZfWYCIvbk0MLIcisEH0i6gb/8T1mmS3WDT
5Indn4ECvoAGXQJ5xxC+X6WscxzJAPrRuZmeQpbce0Y+Y5OxrYCRxNyIUpllSd4c
ZbGbqYD+9po3cTsnsACwh8GB78ItAyFBqALB96lCWbRF7xAedHeYZWgkvwvZUxF7
/ZBXKC9QjxcFDNo6AMM28T+ZyA5mLHeaWTZBUDioMnUMpuNy6WszYUbbXQ5Kkc4l
PVhMhMedIPsgal7zgNQJOxLueOUrT8/ySoqh5dae31hhgnko4PyHq5eeIn6pZ323
Kj6gIyv0lsXSgMifmY2o3wc0p1mORL9S6oTrOTV609beU54jepzSC2/g5mcfCAEE
SGNPfhwayOwF2+BMm5FPO24LyrEnJkWgYnM7zVK2oKGg39OBPGA5K059EwLteZ2U
XRdjJHQx/TNsPCZsHtCqMhjAiVihC7qDJMJAE9uq/hWOWZbeLa0wZsuCxNxEEMDl
RW/OKuIvtiEzk6W8vQp7yEJj9KJFMxW4rOcWIzaYUnfeNHU5U3eqJKA0p20uGUsR
7/+ZMsY9kWkAbVN71faWLm9YbfqAeM785rgpf/mOFOoHPvRnQokxWD5fqF2eeeR3
R0RgMeg+pb+QkjMNLd3+9s1ZeJNB5qwqQpZybQEeddGUHST+1mBrTCFD5kjsY5IR
gbxgLPLeyuS/AlEipo4UJIGsjRPkITTKqiCplHwY/A/g3ZWZaZ7cMzcXR3im3bCg
lpynqkhj65DnR5x+OMVYiMEvhpfwrhhz8YW1efVLKyunMF5wmjY5qblUEs/RBXvO
LOH4A6x+5fgMbCU4m0ZpMGQd8HKUdczGJAKqhRDzPd0b+3Lcth7dNUOk0Cjl18MZ
TjLlp7UgeOTO8a1XQKbxtvG2fQZWot0Qv85EnoJztpp2Yxg2UvNE6NI1S15v89+q
SwYQPCFid4Zqfh8aXgbbsUzq4XdhGqPZNXgx4Q4fRgcx7oSkzD8v3q2BWxsjWD6b
E+lsCcQf6RsdCA9BCb8yM8cR5IhP1ucretwvl3hzCVJ4zbUj39tHXBuxS1lajS9u
rygPaqb55+t396+iUASLvlpnDAFU3sYcy1ovKj2jfhXKQuKiWOzwpPsl6YHas5I/
iW6qzBoD47QPeuY5S7xO6S2SGknKrloFiOzAsYJaJe8UlmH3go2sr0FuoYhJLseq
uUS+RqVgWyWKSDUQ8F+Q8lYRNljn1AyjskeEgW63lE5MINTbYpIzq4qjgEWm7ZCf
UxOHudGgzdlvymkU5g8qOkknLmheLf4vPwiE1tptUUojZMI0GUii4cyb/PhzIZ0m
Bt9s0wq2b6RmYQrZz5FYEUBXiKA0X7zmjMltpsXqSm4HamJt44Z5NpBHGbP9zXhX
aCqWHFZFZqUxG6qLpAlVw5cux6kimGoo7CZPlBkb28wxj8+NOeOEdT265h3d+e41
I5/u23079Popv3n0uICCkGX7Eq5NIjHuuacDb9VXnhS74ef1sqAwVPJPGp7jeXZr
rQ05YDS2FvPaUOJjpvHsyj6f2PtFOmfdh0VkjBH5UoXcp5211593jeNNFijbOkPH
g6l5DoKf9Vx0OBrsLZjkgWuKlOIl3txYO+dtyJL3x68KCK0m97MsquhRIF3d8ECW
jrim+9XuHadH/nw34a3D65eqZxLYIz/YEFrhCQ4C3yOZnKiD08kJGPHfK4uMJeRS
oVj7AYbstSYH3EZiTXVeCytBRXHlebzTzr2jXfeLiT1jW1B7Vh5HvGMmLfE86Z4Y
adVEMjbn7eubLMvPcJwvBdEJ3s9WDFslEdsqVb13+OI3Y5QdIlWoOUe+Iqyz9L++
AEY4xCWOxDQHMcvQmC0BQNf3t0Q/3Bi7ci8jszxAE+sfk1YCMjk4VW8wf0dm8qy+
uE4KZDK0g+jzyxADUZSfuEoqPZ9dXK7Z0haL9/1ka624St7dp3DNz7HxqwhilDT6
6RfBE+E3Leus72/UnFbE099+xwIWt90Rzhs2RXjUpgDQD1SNmEUKRvdE4PDgT/fK
UZTuZuKeNX0weYxfhOkSpSN7bVOApr86Adqee8LseNitFiy0I+qvpdPD6Lr+bX/n
MKTCB0OwyEQEuwGU6o16j7+JU52lsS2NYRqgAKDe0+Ep5LrMWKOF3q67zwOuX26q
XR7LMEdny8LskVSutevAgFtv+PC0puxevC/tVtEQ+e8A8GeEXSQojcOmgTqnM0aZ
dpstSmeat+DPN5MsuZ+dxM4tiBPAyNnF5ryx08nHVB3YZUTq3HY8wesPpwkd/QSj
zFuAbPadxKPTVsLQtJV8oWVhYDAlNOmRMEuJmvoeKTCQhR1q58iMx1H+p7JeP3hn
a/HKGvvA7tWnJ2kEeOctJT4vhfA2gnB8SVVHJAqp+pr4aJTpYeCI+/D37quIuBX9
janol7n8boZy1SzoIVfc2kgl7j+AeFIMAZV6PAI7Nm/54u8WSb6XjQbW+Jn3Vbix
kX46mdWAXGCLiIiyFbZp1VlIjcD9sWjiPgYihyCNwQKQpD00nP98EM5KmI5TOYgP
2jox46qoWLaQ1HLUhlqVBRhbE8FIgex19d4pHwJUxQpOwF/5eEb22mDUsOHxUk/L
kZrswjwzAfR9DVrVIjMerHzpBe+JXgekjKCNstzMJ6ZzQZilFmkl5+qHRum8cp3u
jeneihb5Cp59yHB0hYHCHV/m6gQNlc7aZ9kWSad6GG3YrxOSuQOTzLpOH4XI9lMd
P8UsqPHDXL2U26J+BFCP+RqQ8Xb4l5c/NHrd9VOG1V7nRH6KiDEa0SStn9aU0biT
XWUBN3s9vdflbAUWZE3J9Tb5/AJ5kJp42+6U2/DOPmPIHpCHX5D6SSFMoythXcnN
UeIgSulPaAaTWisanxb6SOHCrUfr9Ma3VHOSciQxQsg5dlG7WSX2aFaIlBccjLt4
9I/SWLuf2/H8bL7mAFaCenLCISwb86ht5pC4npVEb+kuyyU25srXVI4NPkJgOxm2
kLaeiKXUbaTLUOUeO/R5rprroZArtwNk8CfpbUSzsEkqWYy+V+1d7klqlc1ZGQPd
0cUPceu7WnbMCMYMQRKVPPgtaLyWLsHDbO0A2adl0bImo9nH5WZxZyOS8MGZiE+C
s+y/eVXCov2Tt7UzUxC2dyj/0usdT0ptbmxmgXnDC9IUL57rGV1DG035aif3k8yZ
50XTQ5BdbWpuhD/27LeG8lwAFsnRu4aFf4+Yu7bo6GL8+n+3GRyXk5oixqIJMh9n
bRHFOtOx4473Gx26uMhgnFwGeO6Rz1aEk75LNhsFAeSWdFJLo39KnYmkJ2QkRbS0
HyRwcsAa+1TI1HfO6oPix/abujPFrukljHHwgMS9912tOaxHaEs4ZA1lVVAOYhHa
aEjx4NKUvNLWlYfv6zrc16AzTyGTWc3txD6RRSlcgbalr8YlgwTCB+okglmhhthW
nHulToKDZH62d1caLJ3SvKOmLlHsU9Lv+yYmCF6nZEmy7kmV/dzpAKLgPt8FfJqT
6CbDzyAz1gpCeCJodBDOqai3802BJII6NmyRswC5ugdp1yfpsKGeB8atBaOQk440
93MbzGpYA9Aom0PuAUThp5z8rkXj/MIf5gPf2ut7AOhCkjoK/JxeXSWO95zsw41w
b1aOhabgfh68PGjMxO0NZSF723RKJVuXsWSHOnJDV/QwKYx5Lyb7pZeGLV60u1jp
MC+mfT1VhLovFZoHMP/LEBna/alw1i+wLQTlwZEQ10JPOlPhAFqkik2CoAz2awOS
9W5GJCsR6eQxLFNRE+PVo7bxjCLZj0vYHgCUDHmNJoSavg2sLC7iaKKYJ9l7M6eJ
EVUpEbPicSJIdWao5g8qwh6eglAgvSXSQpFYQVPKWWd/Zf8/gqNjVtj8qS4sc+Z+
C9KILp2enFdNAzqhG4fdeqyM7FiKWduAgyWTst07o35cs0qUMgfTtdgoUmNSu0C2
vgUq5oQGSbwNwvLuA70UVocbIXps3TwuPbRuAVlkbIZc5rnguit1baunzEsyeb4n
+oVnIirVUoeS3NSCpmn6Z/9CicZ1qU5dvd+2TU4sHYPwvf7TbOM3VOadboArGAxq
FJznnakG2EG2piEzzPv1SbcHdX3E8G/4yjoNDaZwl5ghV6Q/p0P2/ft/oJ35yl2U
VTBf6Ph5QZki/ZMMqOEpFKm3qyrFOJbLPViFd3aAmr41aRzXfRbEl0VCQn+u4DZk
RtBd6PjsiX6hPBwZZOCLkbFPzzqJkK/wspDiTcxqsoBvZveymCwWmDhFcjYoLjp/
LICAT1apCfZsvBxo2hpjCuoAiVyA5v+csyVNX6jIpi1jSaYICqHy8znUj0DqPQIn
VnZZc/p9fyh/R/kUC2/gR17UYPELvIqp3UPOUoZG9WRKn8hAkxy0xGIvljkvnMZ1
eS6+3WhNVxTAVV11rqvBqUD1LyZlvgwmuCLTqBgT6s4A9yCYoZz7vMdmzw6AUiZZ
NkGLJOKAdETCIydqXwt0g0AInKpHoswJu96qL8Clna+kHZOxhBvfLyQY08XGdHPf
xgEznpP44cIHln2a8qHPtaTpuXOga1mtRzpxvkfqPWhuaJCp5mBf5H2l6FhWXlba
Wc9icDoxco869MYPXmNbeWqRff56rVXVdTwFexS97y/Y5is1RSlJw7TNFBdfVRGs
TKx9CPnsiAXLRe2KB7iqxGLD3LXImyzcIQnnJPKEEQ8Kc1y6RlTo5RllbFdR9KEP
pnjHvHBroTPzOg0byfPAcESh45dViWXqJkF9anuNLEl9XAJw5/EbO2JELyFrT0DF
jAjtBwFWlSz8n8R9rvALTQJzjLd62AbmN39XtspKMxUuMaztAUAPL/vDbLXbBXbo
KLo/7h+2cMFjQNP2O7WQvOo/6HQ30x+yZ2O3ocY3lG+yfXFWz9kTfsd6vQtepJ0J
uiHkB7WIi8h2z6gaW+OiO5J2K0qTWjyqhRsvAT5n0ZlAmusbJFFcf26Zez2vOQMk
ebd37BjLRU14DZNuUku9TJGlxQzEIvkad2BvEYOAQaY1wB/xoBqiqZVyB+37tUkY
SRQGus1n9iqTXdksfyA0R9hOPY1xz6mOhxtpa+9UpkM3b8wNo4UZ4IxK+rks6Wli
gtluGEmafZiqNbon2SjL7Qj34pKc0eWTgHYmSMTbmuYwCsjvGCNQR6YHwz43z9BY
fFCbVAxfijqRtz0255jh9LI2ry7VA6bkXRm/P3Htmi0yN5fB+4VlfDBR55ngeCmZ
P3Q8UxDqUN8tqq6p0YR5kumGdzlOntYy4u5uGXa0MpLqdsDwZBBO1gsZAG+zHePM
MiLI0vy54lPPEAb3rwoDNArelqSu4/7q9IQ573Q6LNRNZD6vnKBEDeFG9qGIPoxN
uix1WK4tQF5u002juRGT58cpEap+iotaRQK7x/yOvkoswlvGgjxE9GV/Nkw6jP4D
5PNRHidoDYy2KvzWMCxmRx0K99j1euv38TzzjgcBntTMoDU8zT89p/pkdr+JDaPg
0MBYlMAtdTtmEFiSdoeCd6AN0+LH8PjamNIEnGeCrLLIR+wZdMj0DqwkdTMRRHBH
qIOighaqDf+xrJUGPsy7SQG2XlpOid0vN12eMcCL98cg8TL8G+M2lz2OZjUqqovx
XmbIV4KGxqPCcsYdkWOLAqfCLSpBLdEHoBqMCBh7z80C/YrZDHirYz44GtD8wmgg
M8pYnjGvU8vzZrE+9ZVHChM7sg2LV6ERExGpCQv6wnfckMrSU0MwMS5KVYrxghwm
H5BkAkcfWAaTnYkMSVYQmKqEPhW2rjyGa+EzOLyKBfaPT6AhkDs72NN9G3wXMhWK
yYZ+Fv8ZztpKMhAv/QDpD/VDLOt1hln4hVY+Y75ChCxh2KwLOwi+26SRvd/HL9NM
9mMAWC/31IZSEY3Hzi3TRym9yXYgYUVQW36VGuGGMvLq1meKyOHnnFU2UGenqDE6
TK75YbPy/F/L6ea5JJy8V2Z7PZBR7yrEwugowkyZv+wZnGGyglZWmg5RRHjbcCyE
qiHVqzLYNaJn5ZPiB8c1Kegx9nKnil3wAD7MoKHjxaHc7rC1bk2Z2qRBpsChHha/
O/sai0IrrMvkdG/8fjtBapwPzEtEMutD/JGQKOVozfCHs2Au0TAeFbQdZCBv8a0G
wiW5iphOheFMtIfhPb3o5TNRSgj+zrAIhXe7KBS+m84SRktF+uBgS6aKpfZfOuxW
GXcuNQIiM3RsF2wWnwMJ9humXRxncgAlYXrYxd/EkLaiClkyQVu0I6xxHg8xhBBG
+YRETtxA0GtSYrybwX1csG5s3zMiwOoCP6PWlPnE7CrfWbFLP7B+dos7RWal8PjW
x9K2ATzydKBOiTLXc8YryrEB+c/Hjl4BuLxhHbGCHIhWJ6PJ/wtB041k/She1szg
XY1rGDDwcBuN/GTS85mvWtZ/sdth1sGWTwtYfhjTR6rPiNKoF4xSFUeYv0uyHU0q
0C2HO6jA7l6jjaj16DkDLu+IveMaGMqH08DpbZ3hKlTFIeKdgr6i0iRU0ZBt7la9
BZHUP6Q184j7BY/9AYamRpvQet/AsjhFpDVJPBb3DvEPyiq6WWbg3uJd6CdwgEBF
GKn/HyPq2uce7P30nPV+WwCBkHD+cOyF36HymbnKOm8sUpZomG5W6DqLpCNdzIpj
OH8EIkPn9k4i95B3AYRDtxCms3lsgleKZ1iKuvhW095/oEoZpi8hgwZKL7PLuYLD
w7MYQ/eHmi6yyq9p/oFIdZOZa8+1HNj8wBSwXFyxMxVxzgxHFjnirizCr5CK/4eF
0goNmyyXK/S24c6POEesr2hnGjkj7nw6U8jKk7P5zL/G9DD7TVyaOd/3asBvVsDn
nEpotwXNeEohjx+8yFYxOdNwOG8oUS5zgBGQ03y2Vbp00lGh6GIeaOPEpoHZ3TBw
3PL9uq66N84umYJaAgUdhvaV04znKDKH+nzsNT9eKVAd/9RppOvvG4JVhNNQHxV3
cv3dGp/aS5yr86eD3+jcOJsFaFDeLVSe6SQwnhpppqwiJgtw+g+k3oChFxfcaeKg
8gG/7i1XjELWNhqSV328NIpCiPZeAbq5dmlTzBDDcfBRDeroBDXK7nlrsUQxNrYm
9p06TVbMvEURRbaa3FL+QS8vcvgnFo1ZImzkFJyzygAL4RFdeEzL9yEmDl/TcwhA
aLnrStdLGD9JgzaXACYL+TDJGMkqIj+++4Q2k5DVBm6r92RcUNhtFqwve2AQsz0m
pJIld3EP2OtqtcMO+SFRjPbghEZpbcr2eJJp3IMzV+RfYa0QsAzb8S4+FMinHJPx
7XzhFBGVVc+wntmCNxlojwhBZGh9dSpY/FnPdZKtI3DGQC79jbCcmVF5wofgite8
gTGpc04OOzMf8UbaRksrxgFIw1n+UQ7TH0fIPc4Jk3mqG6+M2RZ0LUClXT7239Jn
cpT0MwxUwcYbKo+cqrUJpGO57knP1yFM8Hsv+uGfAGn3+d+glVhMIk/yMnufe22s
QYMqTA/voiuXR4qifsXbK8P3wSUiOxcYB++aGMo53SoOUSXFg/vws7JbvPWQbui9
AU0ahbnRsulxmdVhzGF895NZZIebqswCont7qlaPTea1BAfP8Or26rvoCTrOrYTF
Yf5aiidwA7BOUtZm4f5LAqtrj6W9bY3jBZeBUGZ5FbitZJBtLLsp7u8y3og373Zb
qFk/an+NQJBVcCcbL3mYv8IxkgN4s0mZ5teJ37EX6yIHR8udiLFqOWOZYpIDf/as
ZvSUgF1ZSGTQNbe66Z6eDeiEHMkdCg89gvnkvMp2t7HUO/5sXRjMp10prcBUFU/J
e+yNYiH+4OpXYP23ejx4TBjFBM1vyvVykDr+CY34ViO94MSB+YAzKdylQLZZmlU4
TWfXzG+tc0nSErts/nlD8FM/10QzwxAx1VOYBXbNWjxt1hPsEfdMYPe2SKQqlJJY
ISt1j3B4ATnVPYi6VFMbx7Cgg/UO0EjU/T87kjqvBDN6PB/gTXiYruYETv+JlROe
e4xbVTCl7IOxhZACNct+gbas0WapUWtCe1w+3MXQt7OQ5GkSZLBkdVQBSLdXEayU
/fGUqai6dmnHEiIVFoqcdsQjpjW4CBprtszcOHA7csow5a32JHxRYCSPUKq7Xfae
HoUbj1kVkCrjTxUT5f//6KZkY5aIYLZRs+G1EyPYRO9JPddGzpeTRhzn24mm9arw
kBQVQlhKBwyUjokWqp6BxLWd8iB0fbe0sQzcpI+r/RAUuZaIdgacdoLEEUYCgWyj
ReuDfeURxJ108KQEW6gF6qPoWrR9XBtvR27c0reuMoAUXR8cmWpsfYSo5QZJEAvi
lwW4BRvQiL0pN5cTtmXxRJL3NJtSIJRFjQfRvujZrMDkBTCao3+C9vjRRmMH04X5
YDXZw8Vzgcx8ZS0AMZaa0NzUVVoh/iQSaUgE8cbn/FwH8uy09y66ImWCBh44IPpX
+XvuvV+erty1HJS2Wvvq2huL/eOZrIIFOEu9k/uXym7bYNdHhcAzblDwij7zImZL
9zKZt7OoTDJTaHTMWvgSeA10UwlZ9Qo/t386pdn8INPEoUJTB0QT53arWj2nI0OF
5jidmPwToiPE1JhzZss+9tLx6f1TssjS5Lekq6++54JyPCIaJtVMpAo5eOoEEUd3
CMQjLMuo758chPxUyIlWTClVbEqySsh9iwrpE/Qj56Jjv9lDI146hh5+j4o2ZZj5
QYAp8ZUYeXXtWgYqRyjl+07FjZtfKG4ofiBl7uuLIJ9SzWXrn0tQPSDcdueW3ZO5
hnuKYJuVuYMJPscRBLbSrCXYP8spESNBrbUv3UP2jnrHvNUCpYF/mDD8zhv4rmc6
PAgm2CJhcppwpjQTgcsaUhx66WR18wRT/nxP4oBUz3i68Od3uuBuGsTjgHMd5E6A
`protect END_PROTECTED
