`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yHQYBkpIGGkPYhaqmMCvhfpFNvRGKcutqinufC0CPj3aqS5jYBEysL2TsM2tDbxW
ArtMOeKNKY8eVENvTahy7fOxGAsrZKWAVAJ4KIKHAfbnuipyXQVhTkjbG21+KZv9
xkOJAH/v6kS6YkApMqYYgVXOCfywbWMG6qg/UT4xgj2kmUF/0NIGod8jbOd9QGp5
AJgdzZc6LmkU+8vPcW2FPxpabPOzql1NCGha8jADtf2uiSnn2v68FUrPAlJFxcV1
xx9nnnAHpDXsRNzNG/3CqapMCAJCWTJ9UYCC5gAzXpblXDI6Bx7HOVtTTgO+AurK
AwdHV1o5poWzpi3CeKzAOrYtoSAql5ZLubxr+qCPJwt07P+YNLm270Z+hwFd8I7d
TbOpNuf4KBenRmW3D4zr8IhWpRs+ggMjp4e+NiGqIFe76OHJ0C0i5rXPNUBhNtA6
W57gx7Zqs8hrKRR0eoV1WHEBzwKzSoi+bOIabF8Y0BqrSJFsqCRvrQ7od60LOzWv
UW66n+wVb1Jgw0JNIDPSpokYVCngSbdcgrEp99lLBLeGAQkk6O+q77qE0EDtzwyD
`protect END_PROTECTED
