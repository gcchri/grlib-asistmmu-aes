`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+32NEOBbHJKbj8PBSWkvFu3w2u7nXQutFcAOO87/u7U2SjZEXARau3Te4sCCLOel
sMqIPLQJwOEl4xbl/o7M7r/CnCOnaQq4Ww6iDjLCYGbt/cWbvQQaXblxvGNZ1RV8
xAkF2XFbM8k5I9fFIGkahHswMbDXiqtgyojWqV1bZMvWs3AhcJ4ap707tYpSmK0g
hTywwpxs8uiP6zqMaFnZJj/1thOV12Q4QEdd44MNStlxxy+SFXbWTzEXXjEDC9Z/
4hUaF9JCLcoQARxKRZ81hkRVHVeK0yRu4EYSQ8gupuJ2d18wAOU4GNUXpNd1oG2d
YMdGYdNCtLrBB23EQlpEgoUVaVSHznomE5rtQIg9Nv58AI8AJVsBih4UwW4tGmGA
zMSQd1YuC+wRj9R8vch37TsLGvK3cQoz8rOQ4uL2pbZoKA2cwmdGPO1SlOT0/hjp
p2C+niNtDP+KMkOfmuGIgu6snvDPrbr07DUHsg2Y1dQ4TZPW3tAy4F2UuxZSaRmc
KCTaczky+I0bC4s+BSpmOKHTU7NNU0AN6pgM/hBwa86hHn/PTzQmxEPBmRpeiSQ3
7UhGpBTICGozq1YI+zDHkqDYdSGtkTH+E55+sV9ydQD7JAxh1hyvZ0KJx7RtptTp
D1iIJ1/D2oVeExPxwcgnc0HvJDrrTvdw/2Ys4RNHoXv2mp500GMDK2LzCHClDW/o
mlZty1nPu4Llpn8yO2YwYcO+CSH99ppg2aV/MsFwEu7dX3cO+VdSTp+jy/gB9MMe
wpARjZIu9PAIPhYGxCVUQ4kTMhsRTIeDXtheyeCrWJMkQXEhVvLWzCQqazF6BI/M
k01vkzaOvLqWR6IP7y9q8xpx65p0Z/C77/dAVQ7dF46gK1cDQWjrOElIYwD3Y++y
PnLXazY/p4/wMiwAgM4/aqB9sqBgWxVfew+zP2efB3MxhFheqIbpAaxzfNRGdzcV
Xnwr/4i1ljgYECHcOV3GWZdjP4NR0+qkpH5XxGu5duX1bOujymmlSQsggAm91D50
iYxzmnpUgndtHCdZ9EVvycQpehA9BW2cs16Zf80b1COnOodwcGggIra65WWsT3cJ
KRjYsoWkabpHD803JJ4LP5wviOnav8nvEqvzMpDMAk6N0esSZYJ1B5WrfS1Xx1Tu
BACNHvSruqmJb5HoRnYI1y+79mvZHK8bznWwYEqtsEarBICSrLaaw/DXUhLewzur
T3VqXs+/ROUPomurb2ShaoFD9tSCQIVJB5ofAYFOh1rmTX51kX1JXNrr/5fhZf8c
eNNXMG33aDI0FV3vWhztTw/KqzJ8V7EuoOLExjj0vClpOcLNhUAG/xa+gP8Ep0wN
x3+euaNWGt3rDLa0khEUry90UrRaFr2LjgCD3LPYo1RPAl7bQktrXI2DzkBx/9PM
GXet0o2wTvhPPEsJjeiRduEdz6dJ+IDIVWktbX4lTk4W/7qjBpDtYNpsBMFcMAZy
DMEnmnM4Cph3LggH5r6avA1yXptQnTn76u9ISAK9orcViX+UbN5tv/K5xMrzL1pt
UTDfyv1AHqGAVURfnQBWHgQ7mJIcGb9ENNGC1JkT9ekyejVDjQC4UygaMY0DyU0j
7jZy//OWQ2QYU3ja7XVxotGWuYJr40JxWs2zqk9Mtyz2wFvgSMpp/Sv2UjBY+BKt
NZmWhkIpvoPXSNhXq2kX4o9jqTVwq3E1C12AJMz4sRmOZm2LWb25+TO4xrO6WQF1
iED3IfAXMOwA91/6V335ljAZZeH9OTzrdsFau1JbCZ1REMl5qkpXGNrFAkHc7hLC
rUIJTKgB3ksVqpZ/aJ8W/jo7O1zIHziDLQGKr+y2CapdwCOfCH9IXeLPm+AWjb8L
racySANfRC11MwfZeOoImlFqT8tgBkkj5cg2hj1x+zGK6s7367sbPTuoULMI0l1f
ef9J9sUTSsGy34ST4Z5Dk2fG72hJmPg9iJWSsgNCzSjqGwwom16pdTx5cP0zDGNo
vmNGiXJRrhtamn5gfA1rUW7dItv8SDY5ZfbiwAKGpoUQdCtLxitbXUTDflc1VDlS
SPnRH4KWvDrBWUacZB2pd2mcnrbgGQUyDSYK7QzimdQc41NHi99SQe9e+eI6d2uS
u8aDyZ8W/gKXjArTj/5lHvluT2L/gbL0cjPbqsh+7gFCVYH/BFlYJs3wwqk0hQvc
GC2jChOHUZUPEeftSN3AqjfokYv82GE+y0sg+a4vb6hsr4CiHR9AKnETDlHiy5c8
5a6O9b1opnlZm2RbtOOGxVo/wY+E20/A9dUk1GB0CGqELTuN6O4y0NPZP7VMFH1N
nIYBx4cvjFY51C4BSIu8Oz0F/Cw+DrSBU10XfDdUg719ZjXXNznTd/OINsOFfadW
u6dzAbpDYmgtW3MJCZ5068jvSiiUQIx8WW0g38K0AraFCqHAoJcVCs/sdft/33MK
hzluvTAPruJB1wZGI/Fa92pfdKwh7+VoHDX1J92F9D6wN8DhB8LSzBMvd6uyJSJw
vpdbVnfd0tNhBiwfq4FxW6ZCp7LbwLJcIMpIG1SREhrZSmNUBTlvMNrCsUvw6Ind
lR9H+akDSI3BikSkWapalhQqZhV1yz5/33wfbIhJ7bVWN7S9q39xMgGs4AgcX8Ie
VFKqkoAZC6iur4ehztziNEuGwrkj6G6WwvyPJPP5POfnEzwPANtRwFCZVyp6+SIS
dSW/CkHtNmX0ND/Y4WyvlSU90zKB7o9eekd3xpJjQbz3HkNFQSn/VskCzXdBYS9x
PrpgN0RO8HsV283E2QqVn8zh8VcrihkiXjEzjARTEtdtfmllCUf3Ua4BVanrsGRQ
ifunrmP/E9OjTQO3ouMyb5qlxZYg4MpOL9kcy/fVra11hanusk06xaonbofTl6A4
YeNFylVhw5Nwxf2l3TaDfKc1MDMZf0BF5qVBIXcNzYBZl2qp3X7Se5GjWigMMIJZ
Qxy6sRwII/baJ8EPRUan3aAEq0g2/tVodnk3rmGv0hFwI563QrMj/ow6sIOkHM9W
O8yhEjllS/3XtqVKT0QJurhqMbJOsO7qff3hEbkWnl4P0Kqh/odV+9ydiFEKdXm5
jcXwBmnXhOVyT0470rJDoqjDgz7ZJAuipbWvG/ep+QyWUBEasTI8P7k4PFstctlW
msxMt10IG8ydyJjXF+COzEimRiHI7hNpou8LtqlDhfHJOB5WrecK/RS/tgCqh688
AZcxgqPp6exRgLf8wD641OQImirtzu6O/F4L/K3ntb3a/fJaea5TSwXZ1GDl2cqA
rErDDBl+D8jxjOz5vd2iVnwdrs2DwURs71J9qnyq8JrCJ3CuKN8TBkSuV+Tqg6xQ
wDmmuBQ4LT/vLBuinXk1etRQYD+tSsGdfmHXDC301GyYH2W+4RBn0+dxbNr1CeLW
A+OY91lCt/n3rVAmNJEXpiorTibPhj9wtj9/dlscYg+NldKfwAXpM6GJnT8DBoOH
1qLor/AjN9Nhsg4H596erYUU7cVnPrsxpiUIbsUvopqhKJhWIpgNMfKLh+GS1ACH
Azi8JDCblpSrBV1oOl1mYlRN/HOvl5+8WWV65oYWSOxdGJvaRhM5sv8W15jZrCkI
YuDQr9aybrAVDI68C0B64Ox1jtqFuSTHDO3FMrnF1kXkbYkteRIComC1Xzn+oTkD
OZJG2RSSObcrA7Z6Yt36izJot3i2wGFzRmYv+gZTyeLmgU2GvGxCpg2fUezIclYg
1PH35muCr9EK06PlX0/r7sy9BFyeX/aBuk2owtwB9N9Kw3zD6Hw74yvPcy3hhFVs
qWeJVPrkTgiM1S+zu3u3veUGGoinlbqn44vFUcBdfYDvVlesIjEgmb2C7fQyhY+W
m9O/eLpBM1Urrwx0lI3pc/P9QFP/ZRLvN5DTdcsawVHMDV1l1sJkObDxhI6TSPz/
6wlTqXIInbmLOuQXAv+FOm/0oCWvqSc/dBFyw6yZ5PJ/VpK1tJI20qrcSUdy2ykB
Erv0uHYoCgLc5BcVmogVBG24FwPMmxWSqNR5+AYHgLRaC9bJTdH/s85EWM/m0VRx
yJJaCc9QMayP+/kPmApFCnxR6aqJk76VHUePPqCS2NFWQLxRx6cM0R+qnqrHYLjV
Fx6FisvWNPrWKtZM6+OhlGT9scTRU3a24cJ2jnjYSRNhjr0/9coRBMHbUQLaMilP
CAEQVuQd7OdY4yY1SEbCvZ+5oOPYkH/PNjqx0beaS0v9CoQ2wrtLgGZ7UvjtkKSQ
+pkEpui08QU28TuC/d07bLDjK3aIS723bG2htBq+x5c9zHp/suFRHHdND8D+p5Ik
0uMjQTcXMsbWU2xmFlGBVKuZg86KlHi/m+JBkkzF242uit+2Q7G/H7kGenKJPzcW
6lsElUGWdSF4yGtGuEjt9m4s/b5BJG0t/g5/llCuLnCTP2KW5FYB9LRDB15C3sAV
HsCqQ38nahNboqTH3ZWya5OvEvZvmQXWzcKtH1772SaepVxwGkUMkZG55BPcDOwZ
ARYXG3hEks5NkdeB3pNO8DRaTqzuxKJ5gBVz5rabK6IKElQdlk7orSz3KFlgkafZ
70Gabj0D6ec1AIJcGmJulsZnRvN/1NiqIxuqyqZEOKteuUrUnmu4ihW0xx3wUvBV
q7czKjVLVd1lwyVovy6Fl3K/DMt+vimhG2HibkNd7HY5R5fYSZv1XVaFD8yUCUsp
NigVOYTheY+7dTC9sL85BlV6keriI9sS0TaaeX6if+UTjOF76s8xwOkV1X2avbiv
yMmdXiqQ4G6IFJJKlV38V4t8SMQqvTIJMELbK9PleA7ZunBFZT+HlWsI2C/yr4wi
0xpraFrRvL7o5P+6lQG5homNPGmYJDOncK/mRUpK0HYeAdSee6rvqBl6cugrJCf6
LzPK00fAfBc0F9RzQtZTqlZ3WqyqfTS0KzZsHk0JB0BoaPsgUck0vWsEaspy0ph7
XTNtPT7AvvuV6h74yS9c+I89xMlHQBk0astYPPqNGRSr8KZ5UMXF1t/X6BAH5cs1
NvXiWDfr2qZVcsPioDELOG7ScwX8WH1zo43o7oL0vFK/YuTrz74ZHjQsyiKJfGAj
M2ojiaVur4u3thtHw5nc19iwhLDnahyoI3uZMb5rRp0O6VGN/+kcSROj3QwH0rGw
6PLyO5BuyqnelzoixHe4YnH6FGbb9Czi1NvWEsjOV9/+dGldcoYaACqDyKjyiyqu
BBXZxdB8I1FLYkBo3amKinuHHPVzUpf26gdU8lI1xcs6c3x3yeE6NYncqB1Hl4yJ
U9BI/zQuxNb4Xee2/T7DcAqQKprq+20RWxJTOMx6EsMjSW09PpKNayMnq8fRNDk7
veNGB2x3skwh8gZUzfvLMNYD2vtX3ccko81EpFvJU1ZVxFL1ytW73U7owlZqTdJd
aUf94LfAgV9MFMeZ1e6to3sPqtwBc+cbjoRB6ZCP2SthCXndMunCqkofSEEYAdww
HV4RcjvacCDzLUtPjqHUNOqEdgmpXXmWs0U2y3fS452OUPdpL9HFoM7BX5AyepiF
xohjeAccnuc0f8OmSTvWOBvCpusKCrimrJbhKcrJXIlJDYD2h8ey25nMdoDvAmyg
zOXcX5Qc/o7wR5NkAcezn34QAF+mdTF8xsQzqG5qkHIOqYSFusCDmQTiY5zgsL3u
bDiNbddShuHXY9IYFUsVtvf1mm1gBRmUze2u895Qk+g+1P3tcJqg5Zd6+5Mz40su
2BOsJb/0C/oqHoby91PrPgFAXeXK+r0cSubrm0+HfomnMA20Lpr24LenUakL/mDs
QwkLwpj6B6RX1qw/BUS/vTaUy8cmBUKShMAozC9XCDrWMF5OM31roxuJTIn9NZd4
I/yTnBo/g08MiPhI5PX0Tp8hl9UeG9HZeUxB4lITFq/wIdjGPqzM1PYL5GHcck94
aJEkm6foB0YOGQXygU5iQ9dTdqY3eEKbCYWWDlcbnkPFbbZZn7DuoMZwwrfcJRCp
GJ4BsMWGYp29/MmKD2L1EJfhPmQp97RwKhAzGqfHWeZcHzaINNgpz/nuAKrxrj2Y
JCFw7q7PI3riQsWV10MVECE6oCbGL2pEprXsh6ObVN0z8t1732N2YSj0MQqhwiNP
kA1Pdzxw6W9E66Ua2kq26uMTNBfDcmuzt6Djs5Hvs5vQnvvWGpAimUCAz0mzpDm0
NDDVoF82r+4OnCIOOeAEPP+tjHyHpX6DT0jmqIpLfhwJ40FiSfK18kQeMkqePjVT
a7YC+/IEZlu70iA5VoAQUGakwWWstna+mHaYb/M4vjKvYV57YCG9nWe3Au5f9yR+
Q3M5Yo2EukulB6EXwZjE5QWKW5Il0MWGB+8/SugmwcYiDfnSUMFXWSEbPB8vaWGF
eQ0skAQWh1ZQHAhuHabY4oxbu00zf0eGtuxy5ct2m+/AikKpADeshT0VrNOWAtje
QZJuhBlruJtrxfaCwan4ss4UAKj7S9aAeZH1D7m9fL2DYP5CY3Aw99upl0REF/0I
uEgC1arQ4vhFtckfQOLpyc90pRap+wTzGFQIkDgg6om6gXbsjPCaU8glEZKKbYOe
0LIPnnJAB5/mte8CRZ6WEzQ57rnzscBKqTFAey3yHbFrsstV4laof13XkWEXk90M
LSLxArLJOaih2KU1ek+jzXPPxskSIocsze3kGcNlj+8QZpmRgVUXKm3VpMjNpRcB
7Ip+2HWHVG3t7RjNjXYSOJOvvD/+p38eAPwG8BpQOnTwLLmpZX4WAuFc3P+okVgM
SFqx4OrYYBRdHq6GaUdkge3YlNo7tdX2h8SDYDytcemIpVHFiNAs1434Wp8jMcQ7
lU6NsqNRxLRP8+FK68TItM/WLjCFXpHDvZ4n/Szf3WDs+gtnZOFuUCejS1YsIN8/
CuW4hyj0RZyviotnmkIi5DccW/Hsugn6otoZIfG4LqQ2ATGbUKjHfeT/djsjSkzo
2HEQZZnkRhmON10Z1a2q7mS+YJvN7emUCYgYOfFSvJ40dYNdkyFJNpm8lU6W8av5
dTmIwYg9uNrjXT/9/5uj9mCltBXhJ4D48DOKYawRW/319AX64b4fYWib93uGU1Qm
W6wwnKKRD8+9oz60eZHoqgjCxQBYS2zzR62tWsfiSvwaYt7s0r+CJ/v+mLmkn8YA
Io8eG6tOVGaxmdWleeUOYNrcY4xZW59WNsANbuwbfB6EWwOQLUVNqH08cqfixlFf
f9/xUdWKRat8UQNBICCiFUnI87SZP14Om6ImMbew6WhX2noa0tEwwR0iso+J1bFd
ZGrkeh++n3d1U+UaZOv5PQSgLOZ9ZB6BS9mh7jmb7yB30NHGyU+ITqnCgIs/5wSN
VU2ZQVacJV88JJhhLa/oqpDLB6Hcm6M2A/8km9kNNi4s5ymKdjtV2qJxQa1OzlWp
h0yUxrsCV8BOGR+8TiHgLIJI+2OUT6BiTUxH1jPOK/0yju1qYk2Fi08nAbJZ3lb7
8MfFKBw8BBZy/LhVGInvf91f44AVgj1l/PeJ1vi3dbkEyqoucgx8vlRgC0wXEBrA
vUA7EwDFOTOcGXvQzyRc5ILeTSFQmqkH/hLWvQn3dCC6J7vZbFqlSTCrq0mn1sg/
G+Us1e5Cx1RENNIbTTd8rV2j9tvPcoahynz7HmZimdCjF3KVOidJOtq5TFAK18F2
94Jp5GFfZuxKKVW6SqoWDFasUq1djrWIdCjiR03h7ZgwIYvvoT8t1WWWNsju7cgt
4TIC5V+YgYbRdVsEdv+vilZsOFF+IXiRpdPhu8jlfp5uI9jW2GnB6XRtRjx+OXPd
0YG8eK1T04tw5t9TWKh4eTvaqmf75A4yp65O3eFeokK4PWvzgtaYDOk5VFo0nZFh
Uf8SoqnqU2NrpCHsASXQLR96z8yBejxI/Gg5E6s6eF2NvKiIGUYmVGXhbwQFPKPQ
vzyaVL+q1YAP3stTbQi2XxLKsB6ADmZeiFfHsXpycOSfntReOpGVqOMBaCpQwawV
WiOvgoNV0/ONhBXlkCd+skTD739+BUuLuII6S31MJAFFgi6IHKZK+DGNhsKfBNIc
rUwoX08WOrt0PSw9SsuJTBF3DrnLmDS+WEK3ex4OHdER/EhJgN+0qFXw22Vrte3p
CS5D5AcHd8e1Sn/fa3Eyew==
`protect END_PROTECTED
