`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LHyQ+K1i2cE1VIPWueCfnnRxRjoNMTILTP1/x9OCQWW/cWkToVcX05CeTxOYNQP6
bHXCamecKOMTFph3wlCbXK4seGIMfDnFDk3DpQCxlpThwAZM1R/XJIDeFNZAJUiI
C3ddsgtacjcVXg9RBtpyatBeZcy9hdZszmF5fR6GS8QFTz19YL4x2Zxwe1V2tJAJ
J2ySGCosighFWQnYCk7ZXtyqwQVGNv1NGdqd0dDMQL/bKXCJV1f+cbpVFz9QZZ77
7nd7+I894XG4koqE9i4I/Q==
`protect END_PROTECTED
