`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HnuMRUscWncjekFojMil4E7fJNk3pg3Hdi5jMOtlNUVT7LxQe8S0MP80QZ8ptyXn
t/0f6LtDDMw/yTtd5y1egMb8/8QnM+Fh1DXuwgil6AyIhWjLDTXZw9gKK1ThiRFn
5bIsFqU5ZtlgXrb/s1ov4f6ucacHRneQZnrbf4dl7xdxys/k9AlaGMbplAQy/kbf
wPrRQ3oXTIi+V37U8M/h2wupZfwvBrDqR+OkZTLhd4f1fSAZOGDw+KnJTW9hfcgF
VmmD1vbmWFnO9LiHJWLcU5FPnLOpPizu/DSv6gYb71utpqip4rGJdEDGEbUJnTV8
FWAZWg6sY/4rwKzJ1osB/GwW4NVaAZyshXRrfpRFeC04An1c+Il49yvRxInGExRG
1mXlvyiku1aYlZiWpUuErOA4T9cSrAClE+Gi/GfI26vAe60sOQc5pmmIs6gcv9mE
`protect END_PROTECTED
