`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZSclvKvosfEFoPki9L4k+BCa85MGCOZGVb1RdzfeeKyAoqIf8S75gQAfRvp20zQA
ALgZo74NCbJFYgxH80uhX8iEBxy+5Qw6oTPJ+HN9g4zDRppFPWDCBQkxKMIXqWOQ
A6YjVm3MZP2NY6dAP91EApOIXQi1ywP63WUJKe85G5NCe7f2AWVGmIy+N792xNuY
12l0qD9Fv94jgaQUwWJzOnLKSsxFT3SBcb7v1jwSDJ9Jz9QZJMjRByjp0u4+2qYv
FpbotczYpYz4A7IL5FHSFtVS1umaO71BKuOm/xLiDk8qYQRW2usHgYRYUW98eLCd
n91jjsGKEqTFHP1VyAUxr/GL3bmMqKx7comPp/D/X4rXJYScp4TiB9T2TAq4FgmX
fF6b0pKNXrwL3q1dQ8guWDSd1xUCvnAqpu1Cf2Rmt3BsQhQMkX4Q/xoeACDEpsig
pjaI22A8+h78Fx1Jc6fggNHP9HdArsbcmrHVKgMpIff5z3sczOSpKIQ7tekHGOVC
wokOehzZTwv4O4JT8+P7Bx/G7flINXGuqHxj3JCGwS+CCVW8YP8LC6PT6lv48lyI
`protect END_PROTECTED
