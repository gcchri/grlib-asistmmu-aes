`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yfcla3C+2zJxoR9gZ2Qfq04fvR9Fi4Z2qLZPsCzZJpC28bjwGF//9u4O8KeI179g
oY8XCZILay+R7vt4OSJOOZ65+GwPaumggTJQyCG3RRqfAz7z19mM16wD+jRMLnJj
nuASIDASqJj2Z8BCLSajNJiJIRm6SOpS/cewRvvdA77WZdcX0WSPQaVtbUndtYhI
UOHu4PjdwwDK3hi9Chw4xOdqMbBJPaHd6Jxi3cuZ7LPa54Q/dn4Hi01UxR4yrQ0R
DK7dngYY4P1uXL5k8m/8DqRZRx21IpgaU3cKLUDX4d6vdH6prNqw8ue0jNcy578f
WQni2kDHjGWgYWbgcXiI3J87PcTXGsjlgZqu0WdexYo=
`protect END_PROTECTED
