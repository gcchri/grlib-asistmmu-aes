`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GGoiXk9WRSj8gEJWRLBZSDs7d1WoYRUFwqYg/Cjk9fvkHgkQJHyjI9gkS+hOoF/R
wboE7xpmPiJlMgyqEgex2OSk3j7zep7we1dkLNHNnASojcBr4BYSLnJiDVT+QDEw
U+KVvTNI2UM3tS27P42RgIdX5jhiRyVCx/zQIjp1UNVZJ+8Zh6pf4p/+o3RHN4Ok
+VQikXN0iB5D8t6fUVk6AU0SDgSqOifsJTuN3lgO09qQpf8PRgy/v5Oxy2L5Yw4N
7R806xZpx0YG1F7nYrq/2Mnaqv4nOkDDGRPk+x7rgh6MEu1pMZL7d7imUnu0OX8E
esI2MR3NNIkZMrweR5WxWmBlabSrHiPaj0YKSoK6hB9h7bJdcUIqmwQCDzM41j0g
hV9funUQxntcS24jcQEyaLZqQXazh8evmxSsrV3n09O4i2mPJo9pzqRYpRsPMVaC
jaWAkyJbryBVboepwwHI26UeR3G+a3YNfxryGZOhEOquFIhDGuhkBw69Fb40pNNv
kpTW2tFILKuBvJNKjZSYFu7tb4yx7D8uat5ohiLFZ5ZuiJHblGJ+ahpLqbZ/bYZn
PFeDbwjuAdiJFIVBA2EMK47qymyUcqI7tSxG4xpWI3k=
`protect END_PROTECTED
