`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kH9nTWYwaIInWjlmKbl/xDX34KFIten1Ca3E3dp1lwsYkqMrm8KvRgY25xZ9KHCL
lNtP1wDfrjVtMTl31C0brHgXO9JgR/aa4hPjz4bNhl/jHUs7Wp01/11VeKQ/vITY
M4Yfry3W/LzyKWHO9Q2QYuikX1wOsfZuZShnsT1wU/HNTuGf26zS3GolEZJdGwIX
r1rYftEbOD4P1awa+MszWpirZiN9BpH1wZeIrWhT5PsbQXRAbG4JUomZFdiB9O50
mymHnEVM9fzTnRKsPgQInxg7nI63XDvbofexS0j9dAqm5y+JPBsFI/Z+C9uEKA+N
D2vOTSio16DJwYVMiRwgufvO+anNpByI5zwPhoBfk1PHpa+JCAU+3GEZQQT2aU+e
xhMB7AnoK+5fnWWQrU+i0iipSP3aye9Eu/Xc8ZjADuDG2ciavXEjfLQYi9VY2VXM
q8nvZWOOiybqdXVA2KrS8H/MXCBLrL+UM9Xbm+TSwrWRmEKtFLPo3VMzypDTJwyu
PLSsoPMJUB42r1IYgL7j1ico1QUqv0J7SPrioSjjkaw=
`protect END_PROTECTED
