`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pG69DscclFUXSNH4SAtYbPlBWzVCjBHxgSCwdRAMN8PVkPzidZgkeOVZkqfA83P2
FXmHhLOB2vC1GU9pIfcs9uZcyQWa6vc2JMNLdpsss+M8jLkdlv8JFTHXbxLdhgJ6
PXHwUrAC3LS2jNj6+gmdKZidPTbwtjccSa9YzYlPsszfUjeO9so62hFW+RA0wJ37
C+7Fa/17FAQbUy88Nu+DzHNBBQCkiMH2pQTzi4VLzksurB8NQp0fn+D4aoGyj6N9
XShbfDp4KGKRl9Sz5P0DjA==
`protect END_PROTECTED
