`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hucTNqzW+sDS+4WCslKOCNo2HDI9HhR1BOZkknUq4SJjhjMjnSM2wkhBOoji6XEv
MoNz+nshI7r+7ZHfZQySSxKWIEdXADoTmmZIqPYwsIhqm1pZcs3MYn+aztt/Z8lZ
Fg9C56359/sJnYi7Ylsm9ANvfDMDtQSwZgBIpZYkqsh5ezeltHzlnYwOxnOxge51
2DkA5epjPOv60L8C3XWi5080HTXrnz0hhlUQrjYeETkYh9JYSwOXUTTs3B3pvnE1
ZvBbzV7FsY62zvZOfF9DULrKN5mf6PNm1FwdaZQ2SjTdF+qCpLvumvruCbDh4xjX
KNunw1pnAvQRnSIxLb4rbgzAx0v/4kVp93Fh3+ouzn4e0MykpSYNbGyQk9boFfkg
YWRy0wkiSRuz9O7ZurBjWhlSNuy5Ajs8GFKk9dXk3vWNSQqZ5Acms9gp32ahhSmw
4YQx2KSnhxjNCcfoLSACA/cIpu3mVoj9q9Rii5eqmFVLf/ivpXHLCZRi1bj+66Kk
K94UVWVkl3eltGHtIGiOhFaKPZPBN1XS56eR24xrYyOUHI5azN1KcBNAZcmy2XvQ
MKf2cGYPpArS3t+/f5xVejjYCCkCpLIArF6nP2pDs8X28ir1pQ2ibbhcxDxCluvv
UtrTFLbcbqrznqPleSB+5C7JYRkMlya3WfREBAgLna34ClWekxPdM7rC/Y+jcd8H
dVBK0vF2KiC4S0M+DVw2rx3CZxLIQB+kzIVifyG2VsjUObrkwonSPnyq80fx6xGz
F6qcxe0YbO+mTxu1tfBI8pPXEd3MHdTj7HPsHYIbDFB2uUQLN3ZsLHVud8sO8kJH
MxZ3mGxKH8gtuFeaHdA+opgBLkyTWEEktk3LFRzzJbXsTlHM4BWHxiNnyu+AO/9u
gPwBNhNBqKGv7VwGUEpaVPGx0EI3L096YIim3V+C9Lw3qtzeWs5vgP9iWihb7nJo
/FB+yge3H9h2yCpEY8kkSP+ygJ87q4wi+BE936VF/X80WpsgIxjHCrbcaE+RyQLG
vnQ5opwtB93H4rJ5wbWXsFBlogt7lo1NCcmgTxAbTL1FWOyLFm6hSOZL94XasTSg
KLt3nS36XeInSdDRfOGkIty+AmL6EOAj4XcRmhF5xAxrFJ7x/70Fm0DW0hdeQwrt
6iiqxX3YJC8a7fHBLATww2XfNUGX+VA5mNOFKDa+kNdBV0YGjRbMiU1T7XDCMmFO
Zr6LYEN05Btn7pgHLFiQ5WvYeNc1W5y7M3VfsSkM2f4h/JkvXF78D8k8aKxR6xoz
M2MKH2+P6n63etpZ4/XecOLwxy2NLQtnPfO32b9T6tbDmnTrc7ZnVqScIa1pTCba
wAaNG+y7jjkivAAx+hoals+uWJ1W3kPN+z2bUi96fxTrnzZ1K5iuc8cj8rAXxnKe
nKBb+/27h8xQlm+7Moq/3J70ZYWNu+plufFYw0DTSfFll5XUhOEdUZGWMQuYCLYr
JPRPHIwa1UZ5ZrwsG9HqymltYVfUV9lnY7f95bcAFN1PidBeNrmRyRTrxCik1YSO
2o2hbc0qdISiJiLM6k+wLn5nqAmmT10eFTRi7UeAFGlURvpEaTCzPM6wparCU4lA
x5zPk+kiqMRMcEHPRXPAxgAfafSMcnNRG8hf9N2MAmXjrCq+7QU8JbEIMAbkcUxz
gNqIlqI0dlQ49eKUs6xOb6dTBl01/fcsuoksJCpwkBaZFv1xVnr0nAyqDvB1cL7Q
`protect END_PROTECTED
