`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gDt/ffPM4qwaKWkdCycYwAcyTVvrfPJ5lQuO/f9sFCif9cfDlh3sbKg1iNy/LokB
IjLxja5lrs3Wqq2/A8Uogo62Ws86FWmLn3z6/7pvAE1iBN5eqBuvz5ceGSGOTMbE
h8JRSVxfKdV7qdDd37aDE9cr5eZaEsCml3SgeeY0lSN9s5vVXvhNEqJt6yRpz+Ec
SvBlIS3UnoHCq3kXc0kE3ts0nAR9y5k1r3wM68aTzft4gFZFCxl1Zm+tk0dYbtLT
4wOR3+SgsOaT/FU8WP7qgolk72PKaaAr+3YbvD7u38bAxeJYEQL7WdC40KnzZgAm
qbOcUi3ZAHIDkbk/FtdorDVAAfDJ1C4rFpXPYWQxk1ei4A0o2soyUkicnExeNlhJ
K6Y3QfYXcpCZQAH3ddNz1DvZb3XEaCd/9X1fk0mLo0ubKe/SewoxNr4nQXxuNxM3
sjPNuCDuiPsMD89voZTdooSwXEIwaI0m6ghfldBMnS7sP36kw7479fhSV2KtGmMz
hwshIo+jvMRirB9pjmPoR/wMrrrrdDRT9DvT7OyAc9ztBrhm7Dj8mMo+jB79vC5o
71v9nMT2zlFikVUGusqSImmHzKIvUbYE1jSov2eS55VAmr7lIrLo6TZugNeNTD/X
qpsmQT8U3qg1YH9na0qln4U746tQ4Q1R+utolFo0ajbt7yHHBkXeQ7DZXfosKueU
YL4TPxo8X+ym08peEPi9Zfe29et5GYqWwSLxIXvDZlHdkgNJgJEyyO35qacxIk45
xI+FNuVztQvM2JRAFot1d8067+jYE02uQWEndYgAr5L7LDGVq6LZf5KoAFK4hpK6
qhwk4CsvfvvwEyafPsmuqE1groHJaOajEoG2JMVlz4hY7zevQjzHZVaSa0E5Pfjr
zF06v3u/FVSoO7MgQyC7KqyKEsLUUl1/2tSJt2m1T3/AptnWba6BT8Zvh7QLk4C2
hD4eW7ympBq+2FE/cxXNyuBxrPI4h1BEDKUGLPGuKAJV63pXeNBpjf09+dPAsaOT
5iY32cZPexst1oADCdgqJikKmCCzBFGbKR4yZY3z/f42F98P7LXYao0bo2nTGECF
cUsV4JCcSwVgLXcAcE1kLrpRm12+Be0LrAG9CcLgonSnEzr5tDzDCFFvgQsETUzG
F6xkbWym4IP7u/LlCRnaZlGIBsCuCWU/O/KGbxk4+ggmcOBPH86bVZlO8oxHsPCW
WuRiAco8pbFnNDGG/56a0Nx5wzlc+0/gRNZnXAR6EUcD81fxpCpL/MO6uvMbsyYq
e5x5i6BV8oNZHPlgS1YCvBho/yBZnSdeJvkXXz05+ImqA9yHE6DHcd1yX6cXULqZ
YapuzmyqQQEfYMn8qtDfYd03E2rO7Mn3pJTE7f4lWgx+5ODi+6qgsp5Tcoq3iOxO
yIeKEi4eismQzydxHUJReUSCg7NnRLMFlHuzmxoI0tsakw/Yc8uhuqCZyXt5f9AL
eSQa8yx15e+lzcr0Gg+zPAzelISzlK2kpuaaV/QcuZ1UiZkHQBWYzktJWUftIi0p
WE2MMU4JuxclAdki/UGbwPvm04QI+qmso9sotjzE6m+QK0l0R0pzQRnDUdMAdsv0
o0dkcvGRg8+HVMv1XhZt+OehCCyCp6+6rRSWDJPS4vYIGwnzXkCH4XYPzCMM9fPY
5mqc1iDdjtW3rtGaTeWDB8hPBkJd2qrlKXb6ZCm2CqzEERcNyv3wKGbpOMf9oBNB
HGAi18t5UQ6Nj7i7DY4Jsvh8b/tYztztnGEUFJi/RKrLWYMgRKbG8XcM9+I2qSvJ
t/F6zwmOJ9dWy4vqIWqq9k7077ioo2C5vkDKhIeNh5qsLFjBTKj81UiGznjBknZP
GrW/lNB+vjfg75YHhd+lrzCQfaE0i0+WsjKrrk2VrNpkfeaHaRXchyiLsWjD7cm9
yPU0KrKlDa1J2GWvhsAa1UtH8BahQYCE+TdGM8nSdAfvY2ZkMS4KjwAOsABIW9cU
aluuFpBj5ytU6WZIH6YNPrn1OId+C/Ly4XzjNq/XHnGb2r29GktwWzCMYqQDDy6z
cCX7b3WU9tA9pJOrjSF2y4yAhWhFfidcS3oeAe5azb7ZZ7yBo7VreNz5MzLtwMJk
HJjr4GfHDD6EvSagBmunxnedy5+SjuL7yj4tNnpgsYtnKVW5UGaOoqSsuC9scZXn
2EX5WB7ljKn4jCaQ2tFgXvrFaXgvmxMyGpAOLVrGT6qXppSjy+0u5Wet+9xklUdL
cqUqGDAV5G3ksv0+yi8/BChBxqPI4s9M80RxBNCSjNJhGX2LdwlYihvauqzbnlk3
rtAKqCGOBNNj/x22UDD4CSHNZqdCKc/5zu54+4vY2yjb4cPKVyUHADbkRCmZlH/2
BXEuMJtj2W0/lMsHHkRIx2/ErrkjnmoHajHlEyRLh6LMFPPAHMpZZGeCmnzp9piN
nwVZmG9jfywhUgqsjTBTYWBDnQXT/beivcSB/NjIH5LcddohhKpE0COwF5eqVebe
h8kIZZUVRBOfquhgea2VFdLX3Nc3aLaC8iDr2O2e4o2Ku07F16n5PXxUS0jmxrEo
xVerce8v8MNpBdybXICUU4jOInyOwoaLRsQB3F8e1TrKdWXfpaE7HaEYzpfzR055
L2LFIzQnpfbCS6k4cDb6eVNPvW0LcY20h/sWGHFTNNOwOWhu6GL5O9fpZnTcRAd5
eqYhGHgPWClm1w95t9UdlrP7GPdeR9mKQqffxzx84/LKhFpEmoRbOV8jLIcH9zws
ddqrWXPJbgmTcwCthj7ULK1PILmcIN80+CNJr6QCwHYKUBhLABziANyBjEMJtvkx
Z5lQ4KZ8UkvbyiS6Rg9mG7sRo0Ydxnlzo10TmeXgnlC3I9MOrn8q7EilIHALDrme
Pj5wiU9WdUgLry4kZInVaF4ZKKBEzS87RegN99SNGGQehDP/jvrPfSTsU2KgKSdW
bcSlC6zFuwtEGKyX1JLL/Mpygg+PTa/S7vu50lzLHqIoM+wy31DV2WiIpaLKdB7r
9AS5eWHlf53xzeeXVJghM+kkeSjNHlgEP5IiTX4ynxj5n/Sc7wXRnjEcZTrsttyy
8JcGJ1n7CHNMGOxQAKhYqjFkariSfKsCFZV4IIeRjhGPQVywW0Xxlg/VzVqRHw+2
gdBoG07E0bBgcdRhy0cV4PJAipDnMonk1i1cz9acVpRDmSKXu7MF1H72ZqJ9cvae
Ot2KTVtZ6T6das1EYd3pxipkuSp0HEJddQzsLf8Fk4X9IcBJms56AlKcNwEyGdXX
iWRvea6x8iMJyl7pgfcXv2WAtO0ke926tE+yedMh0depOdFLlc2PzZP3E8GdPlXo
xN3Cxp1X+kQ/HZnLjqGwAXP9+P0suEtlCLtrGkxr99shVFhkVP6t6LugXi8CP6K1
c1pWIbghwy2omUdfoy8Troa9beBDznZCmhmKfs2zQg8V49x6g3eNySDup/eVsiE7
EgA5lChRd/3vx9EnuvieGbnMmQYuNWblxI7ZhCIvl3VEnmS4bDvPREtEksYplLAz
9tROICMB4cTEYYdjC/KwH6A7oxxeAVgLGZvIwhC2s3E7KP3/UtralUOdPtJrvV4K
M6O0E79FGIKl2d9cYnP9v7omxfkuQYAlXMJGuURr25z48fvlriqmlNNLqF3I3FrS
u+E1M7VPa18SMH/9t9lEXGL2+dVcEpmVF5aEovLymhY4FuDHJUHv5jGReD6Ib/N6
1VRGnFxkN+gLDwUrh/oKrsUuGuSn/Lpb/bqvDEjbSyY1A08Lor41EvVuen98GqGW
egA7+NtL8bkScvNpmzRAeyD6E3ojPr+mvIMlp2reMYA=
`protect END_PROTECTED
