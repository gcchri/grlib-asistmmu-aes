`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l1JH8bQvHMSve3Ngw3/aamPkTkZkT8MEzUGPRRGAgBpsNcV5robICq4F1iDDnVt4
CLZn+CpF1xMquXu9XsF54og6XCPvKJs+KWWJjMJrGGRzwfUb9gi42SAbKVWrW+eS
fn/ztjzyFRW0N9ODWixfW/G3gKMwZNdrZwo5/Eu0AiQKTy3t0Xvk/FvtetJ2X2Wf
rRyWzEPzhqvXGVpk5UFhJy7PT5BAJGyhrmjK4J4poVaSnF9H+iSY8UAX1VgAEx80
YfC1GR7Qyd2nmh6LTuhgOuRUW4vRFlZ/QooI4KM4YhEGWuR8GHdlPw+58I8AiNpu
h9ggKWvu0wTqvolfffumRpRdZLMBjO5r82X3ISqcHhUk8F5w3Z8LWsQ/iAKOM2Ee
5B5hExHd2dYp2m4UO/FOTT0Y70YasCunCQ2lCw2RAygaOUHMk4ykiXnZMba5R1yJ
9RR0l9hDaYB/pfNUigcXWvYp1NVGyPetQLf2OJ6C7I58XcgC6EhpGOsOeKjbl3qx
VqfoxVoXon4YU8MmKRrR+13jEd0FWteg62V9hitekPba1zLh+U5r0GgIvIths723
zAgqADSIDGyuAC+Q3DhvkeQUgqIVXTQ3AHQTRDCrfI1zQrSWRIERGeHm0uxTRrK6
zPT0impkfCXMVIopx3/iCK7yTQ5Mq5P+r3pLEQf/XtQAptXQQ8h9UTKD/XxS4jZz
87zxjf/LCpfmIRmZgk4VhmyjA0o89Gu5HAtoPxsFYgqZdCGRx4cekqEOJarVF9GB
qFSKFP2Uebil/CCr9RvSH0TbWjDfAjiG+wfXqkMMHpTx68wA2OBfGdY4RQcZQEYk
JfsqmPquf7E9gIiGIJbuuLYN3mZfJkNxtRZP1SgIloAIlG1GZNqri4cQpI4heIRh
LWs1JDC/B3J57scQNqomMDdt/fSNI8CNaOIMK6s00BLhptSgV7tN3WUaeXImv1YI
2K9tBZL9n6ngSebZqbQipuPT3y6BOjbohs0R70NnFrPpOy9w5TvSwScZk0gksENR
MPIGQ/RU5duJUuRgDnbfgjFlvwLorr3EMigYd4W2zrNI21LM5Mre0X6vC97ivQfF
dfZnfhaAj7p3NZ3JeEkaOOQV7iKvLaurRwvjH1GFeVHxsFFJDiERbRMiQ2n/+lUq
vob72FKqfbhvJHwT2PnexM8BBPFnYeNj+AkxbTjZDZDSuvZLvPdYLeLx2X1XnYg2
VnktYmq0jDzk9hnQMCDxyzMizvGMnncAGK8heL31fMKIMF/9r8Hu5t2qO2bA9mz5
V9q7tUraz/CsGESI6tyxA4PjVwW2mfgW17Qtlj4gQfxrTJowuZW6y0Ac5CTNxbKm
lvq6s9DkV9WQ3ZPw9jvyISMpcQOwwEUOHKV1X3L0otWB3uuSVRfvsmzlccBMyZBL
OfC6X6A6kNqkcsRw7/nsDvJLx7Sr6lrzgSd1/OarG6abnmZ7rL7uVC3t1E8SGxfk
jhDO+FQrFTTqI9Q8Gq/TVBOnYyoxSmtMCc4QZHH2V1hxn7lvjLbpifxPzL0Hyuxg
+e6oziAQLp270yhnKAjX4LPnJJIeiKuT0MAX1Bt5Fz+6wjwg27sOq7KJc8yf6UoC
g//3+E5H1Jx3c4ZpyJ3EJDQ8fl+dEy2MiRCLX0yL8ivQRA+ru4MXXQKu+IoBEYUP
wcopfY2XNTGQCxOjpSQ/Hwvl69w2K+Kx4ldI96A9/YRGXJ+YIhYER11OMMPt2ju4
kSRlKX47FYxaiF2ckWo8oF+h5dxxgHRt83NQVgs+Sd36A9Lf0d+xZolvTI4d/Bbt
OgkLjJG78zf5f37l35xAv3UbeZ92pkKQ1QBHUii0j2BbvpKEbhZXcWISethSt3kp
y1kJvorstUgkJsvUxnGmt+rkUrDHwMOKbQmcwGY2j1U4fPKKMjVyxdUL3cGt/6dG
t/l2JFCcrn19w0nGmxz3PFCFEUZLlIaZ1wuUHSKW9A9QYRrKY2k83UjwdOmLDC37
Ozl0ONAB53J0zcdmiAJ73ChXbfA/TIkIFqKyQy/Ru6toyN/zP1/hvOgIw2aVPkjI
xSGoP1KhPsYvhqgCcIPMAAUHqKMdluRABRoUp9vaJx76v7rGnew9cGIu/vru66MO
piVBtJNLPNsWJHexgH2R2Ch7D7DFgYriFvPG2GEHj3eDEXSJiUONzF1gvn9z8izm
wT+pwGrKPXjjHlMNVAc8crQEaOWSNv7ICJ4nxJBoZ6WhDTaNxvxAHPo8E/l0PitJ
Bm04NKBGcz1WRBgFhSOLu5rB5uz0XjgQ+ci6otUGWWTKtM36ATG6Ohw/bIA3edju
UHEA8dlExTc8X9dpZ0sTkWkFfIVl1dCJ+AKtPJE6Mdfvm8TOEKGeVwOxGb3VSWyQ
8nuvj0qEJex52fP0VFUThdhzNINaEk/s9CCj0G5uLLrW6VvhO7WdheSYhfkAvbWS
akOWAwkr8XjAk80838R6NNcrYD7cMrqHuxn6SYIniSjXpPQBV6fTHv1U/x1Bq5Al
I3XkPGappOPzh939xOGPFqM1tmNk0fp7eMvXXIlZ3YwklZjdwSZnozp1OnwLcE3r
YpVSB8LjY+frO7YV/AfTQCj5tFZDjRcJaEcpgKFQX5vArlTeoJvsPkvP4cuFmNoT
zfElxW//3aRqWuReV3hqbxrfu+6JFxqBFiwgoq1dBOTGCsFSZDF1PK+U6OPr62KL
URV/9SUfAO13Ur7i7xPU/qFNsvRWfDenRd7YkN9OHQM=
`protect END_PROTECTED
