`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T9oqYbZtfmzlYYl3IOkHK++SebaTbFOZIyXipAFONqlMgKG4fRXs/RNrWsFz68ao
mDxmEh8Aj11Cvj658KlgpGLGD0HkGWQ3h3TIWH6PwVRSe7XZMkHKou8uuHkikVHF
RIIOOjYiN9SWhOeHmMQNT88noRrtDWN+EsvYVi0crbIu12WtpPzO/pMHAUd/PTg1
LBdxVkC88PZ47nxGf8R+r1zEyYJJcyafpIApkRYYKNq6mizqA+oTeIR2Uk+IjXna
74ezSWMzkpgR6wpNTm+N+Nd2Co3yalac7pLFieta41oc6MVL3plOA9jtQpZftEjj
imZ4SYMq1KGk5eVvXdzTZwKzntMz0qNyYEnT2ybN9mRlIbpPcGctcdUXXUcx04E9
RbJU50gYUPkYNv0A1wje7/QiwW9vZB8U/zUWFx/64lapmhjBCxbfA+qDw94WC/4X
z3i3/eav+pzR1thANnd4fDkt07jBzsaqOMURiT3gdZNdXIVIgvF5SRVIv8uGyN5J
Ld0gyenT0fxeALCUgHlJONiqJmXy9nuzk3P6Cfzhc3kPh/oWWzGIg+rdx2lbBtg9
mf4FJCJCL65OH6OFngZb9L6umOes20/7SqJQd+u6Az8uXdTasP8IOnaYIrVoQexL
w6yh19xfTkkqseUWX4YjDQtbg28WeY3QYakq+Uxyb81FkkcCluPiEwGWfU0oB0R4
B7PJHQJIGBTdLzOOHLVoCzH77EW7uyydncP7mGgSl7yF1u/zk75rxOaxkHYoJbY4
9bCdq6ApuL8Wf8qRtrZcU2zsC6z1Or7V3zGNU5q+rrmLSaGAM7sABIjR4E2Y+UoA
ArFWHdNsu6ZEWCvSuu7XmQ==
`protect END_PROTECTED
