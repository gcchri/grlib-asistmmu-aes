`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1U7Pv7TbtLzVlWd+ZofUpWzWP77crYWXMKEO+lZhu6VBa8h9i4pAqPE1tmSwgLyj
cPw0f6RtB0bIr1vLEkMGPZEnzedySpVCYhOi/D/Zolen5U9yrQ3TV2b+XvzEWeJ8
l0iLnHYBk4knSaBl+u0G26Ipmk0GwvRjCCHbPUDYnNsKxIe3nbC3wO3s+ptY5OqU
izgAEEe5we4ggLhlHkU7SveDqlK4R3CqLiWZAUeOLdDwaf7kuBTbOI4jkPZIxRaw
i6sfHSnj+QokKpVrZW3z9+i26MChYWuMQFRIjHU2Tzet1SQFFT7qtq9rdnG4zAyY
xgqvaEZryiojbZ6shL7sPsdY1Co181VRUDa0qj7vl5RShM4bAL+arnaLkVeyALiO
TFjYg1wE/ueJPBBpbcOALBnV1lVofeARKhmLaWBxhqVwa8rNcs0QT3pVu2TgbBkH
tq42of+o9qc+Wnhm15bv/8b1Ns861rTPb+exakfj4ZsyYynGCiD9N8NRtvQgzIsn
JZ8u6sn+A3bcdB1jrDNhtTM51eKny9znVMiePR02IJS8WPueLRPtmKYj+CLs2hyK
Jbe2le1zCwFIH63ors2m2YEewlhmS2x13qAlNZ6SA5DM6Vo4TRQ39mh6+g6rqIrG
LztiXD1FpjatvJcG5uietsZA7aU192xn2JmDLn2GAoFlyaeTPzVN+z6qVC+zhMWE
3UuZFKi2eoBbOdQ6dsaeWFKcfcneY0W0wr7SI0F3yvfIPBY4rzUrwLnGotl6MgOX
06SIoL1VAph9Qjld6juOGvZ5kRfFZfMHyrpmp2hluqs=
`protect END_PROTECTED
