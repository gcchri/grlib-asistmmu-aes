`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
767hBxS21W/VEjYiHcbYNBSvn85gNo3L4TFXZHhpq3XFFRXSLFY0K5I0y8sazcpr
tupMN4X+HFjzDVXOGp/RqWTbPnVfsMMfGqopa9fkeYGOB4LcesNE7eU9empt+re+
ETA+ZJnsgSdussSTLOoknVgRCLY/fo1bpgzZNODZ19sRq9eN151uBIPLncQHO8Cr
dxpMioL8azMU7wMIT38KlA0q71gSJhxoO1ALm0AhBMdo32RoBeOdxQjAwsuYuv+R
d3DuUEoxX9+VFIzjdYEgtIDBJXXSE3L9WlBZQT+bHZ1eVE2HUAfT/SrAmWGULIxF
ZWAQAiiwkgBMezBFVbwvzrcUIt/b5YNhW7KLEdqmC69h8KbzpbnmcKdk99OzHWxe
8FkIcICNyPCL1PKbcc0YGJIhUQ89U9tXWBIHROd3gWTjE33pyCZAHsNphCFW/RCv
peaQbHM3Rago0Cm6o3BuwKX6yAH9L9t7oF0nLvFdYIxA2xQJ4v5K2DYI66ZoU3nr
uSqFiXHoNVhASQVBWWwfBHNxBUxe24KnViMYAWr/0+d0izLw+9nTHUaqSR/856PH
TWrMR83MwubGZWzIraz0dgBSvHBtyADcn1rxcvlBr74JI6iegYmyPEtrYqIzkL3D
tQFDtvj51tsAvBL04UeQ1o87k4X0c0pRlwVValmhalHNd7Ma/E5uqV4tkdDTU4KO
MqKR9fDnpEQ/JsVTX8KxvDhkvTUwGfX9fxN9qlaKfeYlqERo87TRMNs6qp0Nx8Ib
nLZDjGZvTz2orIEC+F8fw0teyYJP4xJKwAUDVspFf72zuYxTr3oQTLK16CQpjbaf
IvxMUTDscRqWPgvVHr2E0quABh7BZzcdihWailNM9fLbUVCgEImRNSm2LTLRUHX6
3WPAYOeJ5L2ZBmhUtgWcGEmemCVPatcGEr79BzJk1uy6SsVJnyhxhOIGpKjIJVos
FMn8Pbby8EaKmJSOeF8f3uifN9putvIdcNCBzpegbmyPwTm/k2OTS8FmmO3i0O8k
niVqp7OaOXuwAPov08D21rvaHIHx5vCUc3vMZ9MQVYc1hCMmSy3PVygJjgwVxdIo
JWO/FaOqN3nRc+HvEucXFHlu8s6x4fidOUb0Q995H4uH7OWc63omS1cFUxYOphcY
BPIm/VlwlqyaJSNq1Bo36g==
`protect END_PROTECTED
