`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kK17gwG1ta4VobuzgSOsKvau+QabpwxVog7pkjhsZU88ECF5B8pHsMetYy2ucQhb
eqNiKIOA2Cam0XZGA5RqQVwGZQsPwYqRHfjuelSGIjuUVMXhuWmyyN/8HhWrD/5S
4knYAjJl/HPEHQ/d34bnkuq5tffhAK0h5GRf/AvJS6tgGPSnQ2vKvu+gV0gs/OOt
hH9Xuze3UOJGN66M48puwOQwVrfWJt/SEkjR3mSlOPJLZRlobSwbhI6mLlA376O+
zEgyc5zHEkbpFKST9yCnjLZDNy83+hYx/46gsdDGHCJcpyY7GrBZt/ird0g3L/y+
qcyf59v77fUGDGtYC3fnvvL59z61Igyz+Ro9zscVeKaIzfWa3nzWHHLl7wQI1Tek
aR+pDWBfVnnsp8I9LROTg0VwmWXaqVIuqurxQkXGISVz170YGI1L+FR6+bN0542M
6u6aoRO3636TT5NWq2yaZSzMJzQoOw8wuy69e321zJP3WXhqeEKhERw4Fg/xMqj/
`protect END_PROTECTED
