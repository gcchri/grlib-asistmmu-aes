`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cMxeATSb9BExPys79BIx3uYy0csCpqiaYHVH/CWlj7XaM63BXmWKfi+iwVEY7PP9
0JbfrAIAAlcGyYxXumyxT2pHtaspzP0wZC1rUHWhjbv738in4dP21+INj37byKt5
IGDeitwNguFWp93QVcaP5sea9cLU+TrJakWTH7UEooKkH3/GopXV6yM7pmPbgMuS
xV/vMd+X79YJBwOZaRXmXk+glVLpLL8qrJL4l21ZDlu5bSHTky+ML+ypW9tJ9H87
/Ojqu0EQ7A2dqXdb+VjAy5LBdWXvdUwfwQmnkERIuhEzOxzMRJBIicyY5eClb334
nODx4ofnfVbKotve0xtpHofFBmxJdoWgRw3CpOvMfvr8cV26lw99u6ApwZuqt+1F
/AJs4BWVJlkpkUgaMM5ROi2Fk8vaeWbB/rwo3ZgOQmabxoovvORmmwbSOh+mXBFt
8NhKerF2hJqfMs2FYGmld5Ydvn2vvNmDizAK9yRPwHvQDpaq+nTyPLZ6IbaXJi7K
rPzfTYUllTS7wK35vMj0dViaW6txBK4zyYMOXvO6tbuSAdp5lmMrXV0krnc5Zdw6
119ag/KAY4iF6MTWPC5FkHOMhIdz0LuWzhSTgT2lq6CoFIcCbdcPR/ea5KAsJabD
p3GrWe18NrdyS4taRoboZO2pYXLKgL2W9V+O6d37/lWKIut2/jNIwVuO0j1SagPy
Hi0pzduqxR++jeQsT7xfaw==
`protect END_PROTECTED
