`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9WfVD2CjbxJjwp1KsHeFJoFYuhiIFzJxP2R+xprrG1GfIbd+fmi8WlDJu/AekRhJ
jsBf0b7UdP3hZ+frSEZgrOYEV4ccmi80zYAXrr0MQukaP2zUlVmxOSIpec2XN5V2
xmiO2NKs9VN0rKPqQQP2P205BhXCh8ejtI4jlhKP8uTLFQwiVh049fNnvHjCWzSt
ZLMMOg1WkpgOyoXLxviRWhbqiWkx+NiHR+2yOnUwoHlvYUYPJVWOpm9ynsYKj5Lr
CRZ4cvKtIwK9GRpiNiQ/4rWu0n4guebYhpfUPYH/ZH9DCrN+aOT+2WmF1FtoJsrI
5IQwH/P9+jiw1/LcJorpBz8HsCbYQ5Gl7NHqNPqyk3sK93afJDGUHR0yjzADtWwS
Q3KWdSNsHfmrWvysHM3kECh0z0z7DY92Pn5cDY7/GwJmUF9qcuUKxgMPlCSEu6Bk
q08MI8iLh4zKb2GyLvW5gAxT2oJDmvFnAYZGL+7UQxLbBw+1nG17kU38UvKicnFq
PfI35LPMuTRgLz3HIvhT356/rnLfwaDlOQA4TuEP2kJQolEPisKvwN+tzz0rqIFl
ebj0SG/QjnvH6H4o7n58FUScc+M1QiK/8c58IqE0lIf5QZ80K/LLm+BRj1/uFhxY
UJCK5x3ZrxW1vqHGAgA39SDBIT03VVMQWkII8EAVZKQ5nw9KVZAd3XPRYNTY3K3m
u5Bqw9xsAv7cV8f/B2HuQk5fBrKw7x1LVeXk5VsLjhSCtoUkUXlqnYdwSdD1SO1R
PbFAZd1+D1toDs0+TZ3N3dXiMvUb7w0TGRBTbHAB1E1GDsmqA8RmaqAquw+mwEej
cIF3v3foWXdmvR4OVNhQYA==
`protect END_PROTECTED
