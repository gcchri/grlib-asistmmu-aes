`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tVt/6ctkWpkdhLwi5sAk42DO38yiSlAlTxtfpA4HXrL1BhGc2u7BbX69huMTSj+N
sCR1gMYrNzJZ1p89WPDV8sFtH0P1m4z7GWB/ut15fA2ceNYoZlR2GyaEiZZDsKNK
No5mZZ/TLUMxFgy0HXrhiDESjAOxn720c6c8YTRVsKBe/Veq815PxamhX52UGLVO
oD/NesXAP8GbT8cXbv1dM56bMtBuq4QgK3h//BrtFLnPYXIQ+L1rYcE+vX5Ifx4Q
gjgy/XGN509jSvvtpeN4x8CS5NNYMt4KMwaK3UbXDDp0B6CsqY1LWEAExWKWjhEs
XqXbI9qKaB4F9RVly8NxLafqSiBc4YZygMBbHvDyBVf+Zz6UrrHqwu59x+NQTHXj
B0BGQSzqo0bQEVLwxnYoEcoBOe1BsqLyCRKzysKCL3dVKtiNeLcrR1EUko+rHG2l
Kxo8VVuXmRTqQY6/Pz1ANnVstuzBEz7B0IFj46ORyqa9G7yFGd1xuqhYtJQ+Y0As
bBz1bvWrtFWV+DGONqH6MGKFNR2m87ad1DmJnT7HJu4/cZKM92jOlEh6Sr0JjFLN
TK15AZ4rq7Vpfg89ClzwhsFg0121hV5jmAZaMbu2/x0Qz3BSYTlmujIlMQdi+4qC
cpT7MYmzQIWnh4CHXi+R6QkSSGHvyThdzwNPZOEtxsZULbRIcueZAw8ZR3aOIMYe
D9APGeKv7SnAYf2aYGsWEycHfKPysCWJ3WGfvgZaYZ3gDZ5/J08Wmh+SBjKTjGMR
Xy+HhWJcieoGgRMj6h834CxLyup3TSXBjOEpSMRepfct/FiSYW/BCAc4r75vzirR
3vgF3Qj7NDpJrbgdNk59hQdmmIw01JsyJZpiIz8piienhlNRVIssPGVoDkVtWrj2
SRdEsrvQcKte+EJf7upBo7FS0jL2BDLO2A7GF9Pmum12tma7TkylPC8zRo4plc0z
KwG0vS4aFtteKArqOgiFSDXQ04Rs1pDW+h43j76ic01ZJmla+dRGU/6Bq9BIrnSg
rv8pGG0pPA13arVBjSuQ1cZVMirNQ7UFJY7RDTJW7djKnlUP8hUPBNwZlRrz8ecQ
Xddyx2rhVMyxdwxP5xrjgc0IrZ/Tls8Ak0h+OFK7XoTBFHlLmJSv4MijPj/fPHev
qKNm0ALbzZkIZ7KooYQznRDm4Ohem3Cipi2MPiyqGiy2voVbiWT9Srkc0BLmdini
nTWNWXE6igs2V0i0buPAprCIGOM1/qkqH0IUZmjWGeo+3CaXJQ7QRxB4JLqae4JS
dsF6/NQowD8s+0r1U/Q/JASJ8KeUm/cguCg7WXNOFvpP2TqegG9oWtHgYeZZgphA
yEeghX2l9fChLjjva/KKsYxyfGiJBHEvCTZKdATMkT6gD9keQ0QiydDdYq2uqYdT
OyPRAcPTyMBrr0526FjEqSLk9af7sd5R7/UmGgl73AOne5nC8qqvNvAOifBLpGbQ
IQhtpbfYkA4GhmysPJfb/YF8+NAX/EVKvtpcflGhFp+NbOxhqA/wv0LXUnY3gE63
47QMtpPESydeg3l0FVuTZIpxB+NQerCt87jY+BbeRHY2kkjpojgKIfQ/f8LUQ9WW
PqdthQS+4wLjNGCO3JuBUvzbyvamXVx0vM1LQd6wpX9r61ELgsS14epcNJW1vDCR
7kI/0JqGCpujQAoE+dpN84vU9Xjn7Nv9cnaFSVub09tjAoMMYAwfMWRjSWDF1Q5t
YNzHUD/BoyTEFJALtu5Sa899rAtYmdPh9zwRuVMIvsjhpGOB8wkIy+/uk1BZdxt4
KQTIPezcRv+on7HAXBOnPAbOvzUZtvYb0tf2oeNXQJ1mMyTfLKw0t6eWyMLBxYK2
XcZUt+/HIVegbj1ToOnjdSQnWwI8YuX1t1LgYuSBvsiKKsCOGoMFqHr/qV8DOdk1
U7gEhoBfNY2fzJfNCFJFD/ma2mJlQf44BcGlaHo4E04lQZmL/4EH6AfU++5V5VYp
2Xks/oCC/ebEYZU/08++KnPLb3brywYT6PYTqJMSIZU0iXG1B2peVXuD4MKivqnu
i04b8hUQP2PXxHiweNfwoVw7BGTH4W7lSdLXw3n6W1gRf6HQb4HwQKdpP6+WBnKR
lQQ/ix+JuEf4lbXiBJ+32F55dcHx65Sx/PX6s0aUWAeyFSbqSDPEMYdzaEF7MEMZ
aPrar9mRjP/JFpW5ZEvw+oMB5XrhYxibDPQyNOzfeIT9TOvVHgyOfKK5VcmQDQ4s
m7yGWc2M8mMfy6RXxLf382yvTEGr9TUAe9rvPxb4iqQMMech8p2bNAG5mwU7nBSO
et9bwoyf8PSBYgrOn7PBGRvr0w6pkPWX6KvfxW+XnbMxqZHJkqUFzrHdA7IjOWey
4t4ZK/kUb8Ni0FwJ906cSPlQ30W98ooVPkm+7/PR5IqgN64KtahTZ1mk4q0xlVXz
mcYGigZDf180hOEOx3mlawhSsnPvQc+fIKsmpmwUEiwvgc9m19VgazxljPMAlxNc
SUmihD2WirY/qCEYLvqojG6mS4Gn8lLh/kisLUQW/baSZXXlZnNCWCvxY21pT7rT
muPP0JzsvSeMqInKBqxUSygzd6mhZPRAkEXNImbjUse0o4ShbDfc3SAmTt/jYXp2
N2vGUoIQ4x7jHBkPELBZtMkX8DrY01ltQXSWt5i+7JrKkkycCVWl84vDb2Er/K0D
XLwXNrjNahP4Lx3bl5G1RTD9PTaqhqD37hggi2pR3HPebRxKQUNr3ebjztHyzG6T
tYyHLR/oVSw9Xb+KVpmaE4f9dk8/suEWJjogNo/DB7hP9OK9PzCXbBE+qTyRZokX
XJAJfYpCTF0i5ymF47Ok/wGklQxdERs6LpUjAtavgkU=
`protect END_PROTECTED
