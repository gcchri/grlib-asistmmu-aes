`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AItc0hkkJJXBEgcYNZPeZ/lMIiNsUMI6xaSMw3PXSQ/viPqnLybTazoedyE4nycF
CYERbVD7637CdNZZiVx8916hV5HHFU6mAWGxxB/QZN/PO35ArAlReF6/F5NVwhKO
4rkX6gjrnxFtCcZ//jWPG0voxnMwzi3zipczU1veuQLhizCsxwrIoYelK0Q1xf6f
0Iae4F+dt0R1nNnXAzeXr4UwdD+Gl7jNFh6gg9sqqmv9JSQUlx5/+btA1bV8D9is
b5RHOEChN4YPRDXrskE/Dou3fdzuxgU7IL0/4LRvSqC88Xnfiv/lgsIX9xCvQZbc
hBunduDIhJ7tT2SLH1+csPogxliBF63XDcCApAIcYlxJcTPH0PWIubRjnJxiTALI
mZW8uwCLWiRFkftVX+ZW8GwZS6r7PjUgx3fUgwtd1W1fyW2W9KJQtftvg+YUNz3b
`protect END_PROTECTED
