`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r6GIQxYgzok+lOUxZuAJYo5xSEqm5poHii/12M0Nz+6KDMVdde4TrqR/743KKuPr
A6q3qnR97+blVr9gUhFC+MZE+Hg2bUlNwj68JYztad67z85bKHfx6uOXxOUuoPJq
+ZGmfbNVHxUzeHjb/vrKELHC6R+UFUaaAmiYj7PrLJIjy4wme9QRID88j8AWxf4T
4lyDe8bxJAdBzJmUrU4EIcPoilcZBBLzDNjBjJnbCVHgtYShIAaW+l8WrG/6VypI
ul45a6l2huilJJe78nLBFMF8QqsBkIgO0Fh0uRa7PQ0GsADpYbTySLkmShatotfJ
iKIX3sAA8AWy6JZFFyqLz20H5VzwumG500/a+/MhI70iQQpc640hbpSF6DXO3tZB
uHESYM3MEnGXdrfF8NYuticBFzFxbf++iG9Z9K1U3hMhVmezHrNq8RCGoLNcZN7W
`protect END_PROTECTED
