`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iMG/kyUysHolrrcp1p+sDjko/5vNt9Tl/+7l+BmWpHDjy7dep9oLJaL3KaUDxsih
PG+TR5I8jhDO3V2J9xuxggSIqWSSJxcTTTEeEx7WF7aUz7zKmKfJ+RiSKDFUTFJj
EnxR5XC2hGpVKBbjcQhZ12fOH1H2MYqKrlVUg3gqpV4PqbliPL/YwwJ0f//go2pA
/h/LPPJn1HnScaHjYHeyD4clAeAWsxSyDFcaoIw9dHOzrI1Gkjp9j8bEs526+n61
nq43orapvPen0LGAkv3codBrmelGOTLpryAizVOpcp3rjzu8Cjtq5DCbU2JmNhKG
SLPKhUKaeM6+Q1ABAkeajzb6r7ap+NVt/kKuSAVITd/9MYYwSmBQBqIA5i0XQddN
6TG23C3oK/ejr74Q1iBugWrSzNR0t+90WyWi6tLEaMizM/8kVk5J9Y3PB35HcMGd
ezw1V9i8l+vniEJWaqERrmc4kTFrhq4pdpgwh9cbuGip3H9mjsGVR+AZuf38k2b4
zOfHQ+ZUWKR1966cO0oFWwMfRxcugsKfGKDmDzxa4Q8d9F7BChYSf0h/ONo+90WK
5cNfQ2tfmba1uBCv9FPwPWsaYYhWJsT6Uo8IbDrRRPbJPg7nAnxpWMnnCvFKZPVh
VAkZMwi2ge3vBUqkCI2W1lJxD6AKJ8bPtXDvFIvCHLnbwhTf82ucbLBLsJrjCLEl
wlWgYQ1QdUnvtGZ4/m1n1w==
`protect END_PROTECTED
