`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bBf5PJLQ1sBaXRcetr7Ex8TxKPa6y3+JhPX6erCz0WhYcua3mLhX8jexULLztBQl
t7QVNO4JGgiT0yaVJCO+qM89/UMoeCGRsQQZi9HOiZ3tjsYcTKFUNfFUrtT0AC04
eq4J38kX5NmBwP0q60Vk8EuYOwoAZubUeYtncdQWfLnHO8PwAsVxi4hHO2gto7t5
4cewjY4asgy67ZmHdW3N8DtZl0RWnZyty7Lq7tWfL4qWVoeCBxWC/wqV7pMOT1Mm
sitUqiGJd8wlvtitOCiZ6zwVIhyKncCRh7JBETtPut9GYrsiX3F2Fy7m3xrCtRku
pkXXnp4UZz2RSGll5KobdnVsj0KAjhvzYfn33YKsUS06xFAjXnFMsX22T2b0yW4a
`protect END_PROTECTED
