`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pXqR3e3r1Wl9/QVIfjEyf8vzbR/S0ISiab01T9b+uNvvYN0wyAo2V8k8zNDnLk9q
0XwG2klXoyvikjwJDV8NBo1SvXwhS7bf3Bph38bQOQXHDT92wWFYrghQ0RC9bBJZ
QDuAvU2ZdNPhpsCon/YHszszuLtHcbDaSJ/qqvIVkfTsya34Raec2S3LNJzU5XaS
CM0hBUBNRljdQKyKuPrS1MnSJJw598upmx88JGKWzHmMGs9AjKuxzdg73pCx8rW9
AWRXx7awsI5N2ELYFh5iuoalKdHIYnDq4DgJTCpfR9+shbSe30XQsbKQr6dXAIo5
YtyYgHMf78H7nGcf4T8/wv8OBH5MJekLGBa6SZRWaaGLHZUGHTVAD8cU/Uk08QL3
UVledjPV2NEVnhQUWf9ghr1ULfycqiARiu77B4LrVXmuQtgND5IyM4FviHfmvFL+
SwTjxEMR8k3bkZ9dZR2E6CKC0hz4riHkp5VksFqSayafrgU78tiBEJc0qFfSHVwn
PbThXyZeycaqP6ZC52KTEoDAm/VZzPcN8wt+U7oFTeyzpvCgHrn7N3hlsSAng7cv
g6ixp6aWv8DOQrqfpeT+oJP2uhs6+bQTzTHmnYor9KX2brnzy2bL0+JNaHfsCy2L
wZk+rd1idbT3KWL7wQ/DtYYfiqjtrVIr/LMj6FJjYC8=
`protect END_PROTECTED
