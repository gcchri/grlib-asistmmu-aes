`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SI15AAuZlLsAorzk/vXj5/rWMWjjOKaRbEuzD55Na8p7EHg8cCKLA+8ixT3QLGfr
mgFqszzqlHEPmYEmwXwS4dYnQApJ0PVZPPo2pcIuYwfqzitlwqzhMfc2XHUzfppA
HEiU3RsBkCrR+Gnv4cVaT08s700qincLLW+aVL0r6eQx5gWKrIeik1zivgqj2AKq
W94JHrcokmQh+0xm7w7neTBXEyh04ama5BChEd3w2AL6D8/lYqTzZC3T7Xg7wPXX
Tht4KtqJEfDlZGR1rqjpfeoU07Y1eGpmBevar+H48EYpIp5umk3eF4VIvpnXro/u
jg0HSv68eaKUCIwb8K4cIX7tz9FkxA70e3NvoRYuwh6eNun1Hm+pcK5A7sqpJWED
lhjd2X4M0gZLFvxGGxOEbPm9HmTv7DUnEU/BmTGLuyhtO8uPve9NnlTKMJXHhZ/J
xr33BxSDOKjm/tM8mJkJYWXGIwDkJk0XT8CnIaO3/t+ELycSH8NBbqzyOSxyKAYZ
`protect END_PROTECTED
