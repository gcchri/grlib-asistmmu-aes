`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b1KGbPBt+KRQDkcunVC/s/D9OZk8ELKiKt6ysBlO/bkN33O02uLapaEMchMPHtl3
C5G0tq+8qtl7N0CyTocbQ3/TQXcWeLxq+ZdseBBn74DdV08WS9UIshb9z01dbcIn
l9Tpvgp0hJf6PB6RJFq+6kUQkyxCq5BmjpyHTrCWb+FPF08iN3IAx0bFueqyensn
C5+wAVpzXRxPxpbgZ5LTBWKvKQRzp0/Omu2WgeriuaKT8bS0QQPooMf9NQbOZlDg
xehLY5ZF9j2+fEfXoPTfTv6BS/+EtbN2bCBxEqGvX8w5bdtA4TpxR4Oq4ZiQ+5tx
2dPXKlIuyBaAaEb5D9n4Qp/6qJYJqp5TxR1OJZkAYf+QqG9pY6jwf/n/63pRRXUI
I9tU14Dk9kAW2JF4Kj1mTKDLXpoX3UDoup9c8qp9c2SQZWrn229NYf3jB+8UlRPp
OGu4IHdxTf98gUe1gGnPgffonnJRveEu2CIKkEdso3s65w2rQF+U1+m+0vKMGNgk
rMvuHu6HK5xYFe3/Py1ASgq5DStCjiLccniWR7wqu0/ViXjwJQd8X6oTyqZdHt43
K7IhKCTgp26hTK47m6I3676k1bM8o1TVobcR7IYfk6p9u3ShS18z49AZo0DaQV0e
7MpHWXLPaQiSCs+scnimWbV7VZxLYL2L81h/qRDAgE0/me0vpN0pe4N5LDmqiOaM
UlcAJ7jDmAFT+Em4/k4DqK6ooMty9zpiPzGaARHgfRC++7tZD2VwrNjQ0ITAQucy
etp4dS4c5pafdljzXVl+LWb9SO1dLiPvhFc5seM7Fk62brAc5s35WaXi4JQB2GlU
oJc6PCrqhNMrRITO9skd+2/ZT9fOybr5f/Z8L737V6oNFaNG5bhqcz0k7EdRpHsB
PetUvxdml4xDdXb16tqEvjNmu11E7y6IGOLPJacP9ZN3Pe/Nhxw7V1wsxcSA/2NG
fEpvgHt2x455+R3tD/E+rjve+bRtLppP6SZzdmZxQ7A=
`protect END_PROTECTED
