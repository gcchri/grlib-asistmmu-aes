`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8r44i8OXo0CKFtnrsVxalIvcqbMJVqe2z5/C1LKqzb/E0LXlRTeHzbCfpEpSXaOK
V0pvDNvIsOqVpyjDSs0SSsto551afba/r1vE7pEtWqy9QMCQ0+5C8PFhUISJC5jp
Oaifzm+5zeZ+6iUO0/H4Cx0IbX67iwvVJKqWM3xBHdIxnZfIQZZAWrp+5uZYEBhn
nsviPIsp7QwhJuziFPccMUqNaZVNHxw0ECcrCyQ3bFundLdcwuJMViCOYmo5SQjz
YbnnIrzhI0dy039dO39Rw6PBLMMBeFAIrHLw5/qeDC3NS1NQPlXfYULobid4DJBz
ZSX0pEzAt7SCQxMU6fotZ6rh2Nkf7j0bP+mg+sRcWqTQPZ8ONLfK87l5PbQwxUjG
brxORnXJB30VlPVs1bjT23W3XU4P3maHbfxlGHjFHKY3SHCo9br2EB+DGVPkS/V8
MX6Vko/9kQQ0JEZR5F8AL8WMH2SbcxR8BSd2UyZR+bLaEHQWhHrVqHUizoOS6g2m
HfZoUKHNCf3LtxHaoPU3C9JoiGe06m/0w7+Y7SGKldqDIdQWDJwNQItLdw0YNcL8
Mck+J5RTfbHNZJr1pRmsxJ17qAezc/yMbn/CLPD+L5e2+XL/jixy1VNQvCsZoGko
1XcoYG1KxUdHSGTG+GO3nyaoWo+STlad1LU5/0f99DrRH/oWYFxcpJp8P3n/ALh2
zw4SShbU9LjgiS6+gWdg6sLOr0ya3R+u4Cu7nlItQATQBXJxwXH5bsFOFaA1W5Kr
HtLzhZwSZFQbKbp25sys/p7HrsR2tML0TrlUi4bY5BLJMxfy+wGgw87oYdm4CLed
G3Pusjup9JP1uMXQVqu1hVMmpvDQec1BMYh+F1Izl/M7wGLgS+sPlQfYWXBz9S3A
hc7McKd72W0Jhgb7kSqFHUAmNicc4HBPdrzixT4H+WXgtpxSwuZWwp9B8nUb8Z98
7tpW7LyJtcYvZeGMfI7o5Jrco7pWP6rV8biwxpciQxWkXvYbk9GjJx5d3GLc0ARq
hVRRbvN26Y1IIUBeFL7lgT+ScHD3xefO4233Xrc3hGkBYc2tx0cl7d6QHgL04KYI
lciXB5FG+4BGpjdiJRCh7Zo9GxnxTjMVwrbpfyDfKOmvJRT5vhNG/lVDSu5ai7ul
0rjpCni2Fe7hZQIB4TvNcEapymxPeJl05sC8puRgsMvVS1YM0TyGBXV6FaSx8lTy
l9UoFnhs8uiLLtoQ5EEGYPOCXSTatjtVwbfhhBJJh+906cW0DifGC+ZpNhHvC0kP
hml3VU57uuhuxXTIpMZevn7LgyPKfQGvRQglYlPWMcx7zu50mxOlk/DI7h2XBlb9
5ZLVvv3/mlvpes7adn1tttnxjv8H7SneabuCyQVWu2bIJHNluG/E/UGnkhavOMTq
DK6JD1z93y5oaUKiMKUv48x0E6cZX5FlUUHoAix+k8zHUYCsq4j7DaqXXSLmkUIn
JWVeIL60TqbY7nomG4URmEM9JrsH9CxqkLVI0ZWWRQiqg+xJ5ZYcmr13h5kBg9fO
sFrnEf/LD5583hvbeElixJW+sUclAFSIa+2eXGp2+tDOO01NAKVcBJfljRSUE2Ws
a/gm2GAphF7alEBX7IzNPj77x+i4t46YsLWPG2vmamMLYSuuZgDC+AHqvFCXs3pR
avxd3UGVov5EGG8ERNyFOXjXm85Vp/D2sF+su+68SRaYWT+J768SbRfxuQ44iIQS
aZQAhXjKJjjNKJmsRtMrJxBr86JZCgf6Q7meAVY7PLJypgrgcpwYGHsnHYmMUI8c
bHPoNzRwBNpKCfr/4jNlqH7BOcy55PbHlap2A4CJsTHqYe3UEpMSoAuMse1LQw6f
N3jac4m2MzAxX9I3je0VH3vBW+ZpI75Gr0ozff4hvAjImqOkTeOzwLJmktCgXT2o
SP0YVXBbIP2GlRZrTiu9ZbcoZHtqREpzPKJ7GKVh9ovDuQwwP5GYtd824Y82KqE5
u4UsNQrFfjltNsSt8TNWr8jyfrYHvGX5GwrF7srJeDPItBhh5/YWHI1piuf9joDK
ve/t1zxBECHbUHZB0mYX7zdJim8atzhdEsG8IJC9gD37tL4AXSbZxwT0uGPUuPfi
F04hNeDNilwR94nRz7h5CLD/Q3iHFDtXrSGGMLUXIrTB/fnMQkh9XP2s2PvQ8qpi
R5LWtbU4A00mQm+Klb/rsinVfQNZIJA9bzbpl6/XZNprkmu3ZEz+P/sy2XdTOvF9
8nSEK4xI/av2cZFDgAAxQQ3uF/vHH4MU7OBKZHjaSwTXGpyY8EnPSBUw7prGF0cw
NHZrwRY+vvt9lBJ7u5ewBFY20qjTfBPvSzR16rzmXi2/H7X/tEkkHMf2WqV5WpBH
oWB4ojfY4W122wrYWEfiy7N6+vsm/g5RI+oPmZmPjiIXhexUmkIMYLUgI0atRDjK
NTX0FgpgkQKmxl+wTKdlOcmkSznXhNP9Ai0E32n1gXJt130+Q3L7HX68zDYtrSzd
Ft0edJb37MwwI4SU9M0vHG5iQFA4rP472NZ/tu+9Tz0OYaStSwn3itNwzkFaccGC
WJeTPfzdcFBvXIOj9jZGu/QjbSfQ4g1Pdtm31X0c9gYtZZfRn0kNIQ3Bwfo7EkxG
fhW35AiOKon2OkM89iI55NbOa90Elsp3IcYF7y/uN1X6zrrmJJusSrsKewBRziac
ktLpjkW4Vnh0zBggp57v2bjEdJE/OzEp+fe9YBSFi3RvBr4Kn+OWvW2u4iPnC4XC
78WsIbb9ZbG0HOCnLnU4v4JuFXAHFXfTeD6REDuFqNKglOV9OlxSLqhDmGBzHpP7
hN/A92tqvjLK0qWxD02PHxAjdumr6KEmMLqx8tMPSN2u5cYKhYL4hQ3pMXRRrleu
IbcUJmendcGWmS7eir4PlyHhy7FcrFzunOfi4gL4EmDYntKLZs2Awv/d/j9x4o+S
ZBxTLkdqp82IxzEaTl2qotNEylppTb2jn0v3q4Cz/b5+ueNwRvPw2WUieOE07XHR
QO0TlQ0AHSIWG62S+c2b4FMQv1VNwlWQkC0kbAPaOovWBC45GpzNNw+dpMLIJ/Nh
jUoa7X4oHmMTd4WX9DrK3+5Tl2B7W2G4AggGsIo76WsF9nEdgIqtGzi1DjMvYUfU
3ZhWd2ANpWyshxZiHKvnPEesrE8EtmxwCoaqbGEKHa+niCCxNnh3O5fJIFcmhzmd
kCn1cu5xjF8K/2RU8NBvh9rhzCeYKovexWfUGVB0DB8xseeVBm//dQJUFLIs8DRo
46Z7QzidP3s5WopjYt4NPTOJuZJuN8Z/JQeACQCEmZXDqu6dzdeMtRmVttLtfvAD
hFvL+0WqU26e7H1ANoEzb/2FpX2SHBPaQ6pBCiJf7bfcERc4LjxoJP2YQAqM9C1j
jK2blIq4dEMmnSnvT7927Amceny4NIsHDAavQCGDVljjWsMF8mCo4TjZ6tAwpSYO
pxslmBnjhbZUuhEcuT3/+bp7Ih0/s9TNqhQwS8m/ks0Mbz+AHGo2ZUEKDJPreWI0
Hi3iy+23U3ZNiQiJCjrNL9EzKpwJxmMKwvgmd6tFX2lp1q/MYjc0z2OsS2yGJfIc
uvkldkDbiXe33E90O5MFpFH5IlS/QWJI8uMQckzphNcjUFDrhri8QBllueUHs9ar
eL/dT19Iysia66uxZVILHzfuBBkfWMzlC6J6YK8rFmadEmY5tKn5MLwCGftUEdIm
fkdPiMDitIgxSu1x1UItzV8+xV993z0zRmqg4fBgKseshZbB3lxpKG/JUyQnm3LP
JUqm6HZtJggb3+OFdqYGbimr3vlwpbiTJZxXzl6jyc8RRnBkmHPEbtsVOKnnCJ85
bw0E2qmBXE+FGj2Km7ufYkssegLRbPLix/dh7M4S/+L/Z2eDIYbNhCM2g/ip2gdC
tmIhzfAwwrdKTkMJuWPt72nZuUdY/aKRLsNYGRZVFNYyoQqdFVd0oRzAxh0oyP7Q
YBOgKml52KB1z4qvTheOiuMIIH9qPkl7crucYXnOPUyWD80zix+9N7d2reU7jAbm
mEmsOLzBX0oDW/i2Gn18hzjvu+e5WhlIs0RnTMfHdnSekeIStGeda0F74iOlt2N9
1wT8J5qMBJ5+x3ap27BSF1fr+vzxmy0BBMy6woLjWoPViwShCF/VorC3pdxeiAsZ
krn4zIlJRC8S4wW+bs+Jqho9OsqUTo/dFCuQ6Ezohtz/MhpCnp4qEQ8S7/l+YQWO
wlHcVHXtKPvcx63SX2jPTk/Fxu6c0+PN/xUeqMlLysMIX2stWpSsXHt6HT/FbTXq
31anSldXCEw6Ab8mMCdUJQUENufu2T2nTRcG0SNDDX5k1vuBd6NEnCQmm546J22l
U54ZH0Qer/gPOKwTgWILbRrz8vqbGY0ZMRIcHdIFzyGmMCQ/VmEzo71jIvHk0iaq
4mJbesB4RqIum+X18EW8bOfSfuMhlkU/k/iH9aPgPYvPbdI+XuP4utwGud/6YgnJ
mtZ3Wq3q2qrtDT5M+xdAflQuTUBahKwnq3nB6r1g3amFrZYjPg2BPKcy5eVnzJj6
5r/EQPNRsidtlVr3wrrkWOIxLsRcKntMWbcOsInVXFx0zHPlsYoKHg9UjWuu7avT
pH99SuchgyDLeE4H7qTlduIJJ3dywmWVlBO9iVKQu54Wm74zX7sXZMpr1qInKJQr
m4koVOWUJz4+43edHWgyJdME/ZZ5sopdtlzGMqAfsqLyNcV0dh22MTS6CBU/39Ju
IFb8hfJKtJBKbDpERmeM/QeXE8nQYFdnBViMsftzsPdkwqxVhCXlNi+Za6gyHSCd
AynAxcB4LsxUFWM+fJ+8SJtHU+K8DkczFuryCpoEyiVJfJQydcqxGAJ1tquzCI/A
Y9PPSXQdE3EJnFwuHBvNen385zXUxsOBRaJ9Y1bWpZp8T87zfjWTsht6o/FLRPpK
Nz5t7GULgYpSQ6TA+1GiwUDEXSZsBG/cRH/EgUn5S8jT4RPg/9faoiNEZlZ6nRkZ
xU+tY5UQkL/Ru2is/4vWtch2xTjM36k9/5yko8+6aL2G8FA20pb87g/jV+CSbEu6
FVa7hppjL9rkHhfu1oond5PnSXty1K6aXvwk+J+1OVoq4tjmaOCA+wIX2uqaEhdQ
l3hoz2kHouYvaSEomHcKNkyaSC6b0ygZLs4+4tACrrAcVUdkS5jvm0PStRcshfdb
N4zWrSKePO3tQ49iSeafg0cVwYpWUmZdzarEeibRvupIJhEg4uFjokdih9xFQfH0
I836bAxjlH6F3734+wRASCJEXhltA2K3h3fodVbCEkbpHuDSeBj/4p3rVFaLc3zI
1x0WCsQyyWrl3Hq/16yRi6KZPzygAnHxHQ0vDLUUjblfK5FFRtEF+6p/La/tw0h0
P8tliFhkAaB6d6Y1LC16RrRl79IfM1mxvGJKPd2P/zl8bX9942dLIew+cxoQixfb
Zr2qFiZdpyW3JuejSrz9riuiLwx228VkskgzOi2FGqCB0UNHU480v1vqrSi/PZUK
5dUw/vaP9AibyR5ZR8bYPj2vgEIhTb+H5a7DMJANmoe8uq76LOlfNkpyTTtGXhbz
vG2V/MhhUxXEJKHqSg619WxTYBXxq2eJc44wdpJ37DPM8bnGFh7PktMLU7+3AvyU
381q6e4o8bREaTWpWmBrcQM3g/QUMclYM5JCWCU2JEJqSs7xGyT5Wj9KUxSzdXpw
iV5btodfcx4rxcxiYaQ99dWuXNiV70XtoN/inKgqlJutGJrd597dyNWLGxmvN4b8
Y6vP/q/NwUsVV+XncG+Lc8dKrSdVsGxdrHboZJ3VZIjU1nSK45q5HuLjeM7D2VOs
/4oZQYz6MEiNLhtr3tCRzTuLqRu+2x22WwT0qZXLndyu+iGGlEPuuSNj5I1gaNUg
FmdLC0RhHWmTkQV8Ty1DPbtmDWcjzekeweKJ+CPYKgax06RpapT1SEAIHFP+VI5O
nFsllD+UoXMpWEY1ReEdWC2SnFswuKjs3jR6DlGfkb6q51RykpInveOoLTnXZNyj
sG55KC1bW0/oqhEWKwKNrlZnv7kZ3aP8MQa3YLfRVxDe+X7CSjdkWR3y1A1ewGXG
O6i0z+xPk7YaiPmsz29bYXuxzwtBip2mHf9vODa0Hr1dF9qTqETb/C5gxY8NxMts
R5MMfjKN8oBtLzIgF4E2NoNTTAAWkgiOpT8HS36WsG1c3wwqJIlmkYBeOvFFt2UA
muCc/BgxvsPjZDhlY7H4///STVkTrjlDjjKlbmyCwcsXiTM4h2apgcan02Hh819q
qJfLh7pRphXY4CrCR1HGKF+y1nkwKRXDenphEFK8k6uyD/xJ+i8OxP2TZ4UaeXbM
Hmdeisvur5xsxwXP14mTIfG9Oaa112dkHQZILZ5vpTYNIXYvNtUEuqruLon9Id2D
NcHbK9eQahG37aDA2WdI7neuAJNtlSW/DkB42U17hP8vaZ1Al7qxM0iMddDeMKxD
eLwnVSYqO6zPOtEoRvj9CLKCyJQk6/BUbYkINEO5eGkDiczVdvhClM80l5O0UUMb
slDRPBE/+JmhR9oi2K0FZQ40W+IqjGvfV+dwj05LJ66hHKjVilpJdz7dNrd36uQn
0LkgDfvAj+9ui0mWEq68/C0rKbHlrQFjE8XpBCxv05WBepD4FokKWAjs+/IXBCVY
6x+IRD83ISVvZxn4sKg14bcVe881PEo2ylHhWU+tLX+rqD128RC07aU4ENjg8rcZ
czjkSpea8g/FRQ+Q3Jsfwtt+iNLZyox/r72wea9d5n4Sa0Zqz1GDz707+Ea8bX2e
L0kCVJohKh1WlsF2EntxtGcxytvEokO9zwtgJ8g0DuU467GzGI7vcupa+VmaYmKu
YDIsUObH/CIuwh10VeO3NwJXcmXud7hcY9PWvaDop8qY6+xq9rwdLb5Sa6Z3Ek9Q
S4BOJiRWr/CTDVgqxkjMsvfbkx6hVrgsxHGbJ9ime/2hJlNzEbslKE4INh690vdx
kgt1lFK5PXrxDG4x/2SQEcUbyizHRRv+/FW5NojEL56hsA1CHPiXayaTE+3wREkk
/33dxcSQL76P1nCHowdT3y7IW6M+qd/WFsYPoSQ7txBa+wWfGOlr/jpe/39NBcPX
30muYEHdT6yCDt/vYqtRLMuApkXyvlZp72oZMdomoDIdUX9FwL/Wts7v6J2GbyvF
NTVU6AEi6D6RE6qzphfCJAhr79XcDSUVza/cmAtbGTVeQv+C+lc0a7WgUC1c/baA
bxl48V4gnP9S4yDx0k5CKLcdXBeZo1AGaG25/riQ1RJ0mm2qSqFTl97CNqEYo4qQ
S7XDZDcb0Aau5sgmJBN36MCtpetPM90FinAyhceLpa54+6j841ZInU72XGzJkTe1
6H9RiJ6QnUZ5dyBIOC7iUAMXBSE4oqkK9VzaJ59Pw6t25ka3cjbGQMb858rO9azd
ZDDQcTw3PCBPeDh51Sij18DxtnVG2sOZxaGkwbn840ShpqHZuaKYlNIh96wMUADd
cPxtyKMh31d6buH54CeMSgcVcIf2cj95AeONhacPkYs9ciXKKiwx+aCGuV4PHyf3
jE6mybrA8gtRA6Mv5NXOPYdI09mmHYlC/IHU87XhrC3vqGnRq3b2QS3ygjAwVAcz
Z+2nZ7ULGBrxqF5XlpmI+nylrUCe0tfTZKmLQfm0urq7LfrVOUWh+KXMQ/XjipVH
5ZXJ5xBm6MGvuJ6NAb+uBc+U9KdHioZ6tY7rXyvZsv14p4kWz1vASRVcicp0Ac6u
qDKCZYjtoqjx6Yr1aRerc8cTfCESgaJZnu5yq8icxc2pbQ7YJers4Zehz3QzyfQD
5xcHIlCGzWox3k7LaZUZWBH6TodPJdNDp9zg64exLx/H4IbwtKbNmdKZZRkTSiBP
M8vg/Bsd0HdXWkLCbGmWiGS0/JRKw+2K6nNhzHSqmNRTHXbJhM1i0TCcCmxzaSNO
z0tWvuLYtP4fS6Icytqq7PCPHguUfsEwl5FcNRXz/48Q79sPzeb9MWe/XQg1u1lV
aDRrVPWv0g/enjv5Squ67DqkThKkyCgTH9q4vD7lHLX03lRmyhowZ80PLmrAS3YO
IeVZfnELXND/fC8S8v9yV0oQ6YXVIyNDtSJzsZ2pLbyoawIpYHLrGW/eFUaM+eOI
VO0QHrPWgLGcX4QoPbdqwIXhEMUwnDZ1nWmTKYUlZlsxCfTcxheyxBeNOmXCkK9J
GgZuS1JIjOsfb6ZsXEOTzgyMMB9dWN7jRHLnfmGkmhbT7deLby/jeaIP2FLChjgr
YRlEOszqiIksJuJ9vzSfJDNrTdxkDNc18/ymE2lXwjJA15YgMbynbrHHUQeuD9To
eGp5FQ2ecti5GEttEmMQBJk/awvPrxoLErUnWlYa7MqpR6BBDDD1px/O93/6IPXn
xgvlSo34Y0tAG6hc6sv6uNDqEM9/WmNKfgJlBpzBbTsY4yb7I/l/hmeKJWX1gpbB
PkX6k9IZVL6eNKdq3Jqn7wLQhmjCc1xfFcXQ50dUksauuPZvs8KYGwSLW23nGWJC
fBfIIWWcRc68DYC8gdY+MrH9+RSXmhqAAzmq5a6tOT3NLvfbCpAE37rDfrIDUSlf
17EZ3NHX6cHA7mrPwMWOwTMa8lzp7aFLv/2CxrThb5FCiN7PasCaMXsgU0qeVUjJ
gpuP6lnbk54u2n4H7tQkGXcsXFM6eryFpaCRb0BjfaXWtqsK2NGlfFQzEc0YGAvt
e+HYaB32tpoeN0RYR4xjqcJLRsDMMq/OHmDlu5xB7S4dPz8KAs2CRvCGnxdzTill
LTBW7kwPZuUpfLx4P43i6LhqtKXLt+ZwJmENv3yP7NXc2Nsl2rP3iiWaoxOpJNRA
uvn6bqSecpiVF8VYw6lz3GQxqcL+Dt26/z+HMfO+VS413YGWHcpw2gMa/D/grRP0
ATRpGk1vmMIWfXZxGmjp1v13Sn4SilYiySvNo69txIQTJL/fgJUiWFgNdag0c4M0
n8GMtVbF44GtT967FLHZ03eOjpfZkEn6p5tUYNBQRWD5xO/KI8/23w/kWBEllSzC
hr1J5NJHddPzjTRApciM12ajoRL9Qv7H35x1JCO8QH1RrdEO4/ioHE0qO8mIe7cx
f6iIY1Z/9SykIP6l7lRFZIelaoGlt/iqaI0rUz9iPuJkgBb5YacX2DC6KMQxPqHQ
t9zNO3zhLLQi9gMlVc0tKFN3X5Iy9lQ89v2YnpEyNHoFApwUUHb3LHNifEinE0W+
apJhs3QXsnHW0egZEvYr8LSgguM0SAYV4EI7ukQRN+02/rph7N8MTGGVk/d6S1xR
/9R70/hcCEQ9Zp1G/LX+uw9MfdEJtStmarAEyGzJVmgkUgbAC2oIkH0rygdsM+0T
CeGLf4HoOA3SmcAJXy56dXDUAKDFCw526BZZkmzgTWySbR9HLbIJPYW8VQXcAIiO
HZZzY3xZYaNSVqo3UH0FNDRnO5kgPikd+BJ9OaVFMkgQFA2V/FmJnkQXJZSTtmig
qFKpu4bUHeG8Vp9gKdnlyUHo4MJ++31/K9DsKjsX7ZLanfdFp02Tj9tiZbKPHCOy
HW2ep4YBDv/RvC4+av6X8/AtN9n6wmEaS3enRHyqHjGk9oEZSb1MKTTOojH1ozjk
DjfZOPmazctm+gUXcLwkh+yWgT1FIsjeJxGMlPJEsBbfmQ/y032WARJA0Ok/sMt7
Y/Zj/K7qDBqNUWo9QIRmfzQeaY4EX3lTjPdjXkdgYVSeisxdRjlfi/7HnjM547hc
4SVq6SK3X95701jV6iVhU4Ifq83t7dfRbC2hZPuo5Sz2RDxGZv7uEW78swQauW+D
Q5+hcu3PP1jxpijgVtk+Ozus1CHJiiLy8d1hgPzmqRlD/DcJD3Uhp8hiSd25jpWy
hPudiS5t5upS1fqIsyt8ozheBIzTfDUJWtfSWO3TNp/070A0kfsqsRmA6TPKgm39
ZRFCJPZEPF/R2RG1tM9q3s82lT2yo3UrbupoK7mV9esdkRLBm0wogQuZKYTAAj8G
QVumyK8Khb3gdjES47USm6LgdQPWOnTbSw+PmQDj0islmDvVNkz4KYODjyK0/YbQ
BDntEd7RFEKlFP2byOm7cGAUt9QuZaNaE2tK9gmrP/U/w3RlRlwgGmMsasl9lcya
UFJX0MSsGuMiZ4BgspRksY6E//Ch6nqiGbyK9VK48mD3pmMZ79f916JoS8K6l9RS
jho3DsPhKT5wiQtijO+8JeRLcF25BlyUW5CNFAVwkm4GC+bFAwGPg7kI5r6K+l84
4fA6QwQl6EHJmk6Gif5dVdZcvzyI+NHC1uzsXmW8bOyaSYR+AX59VEw3rF7uUxVw
W3vrt5drrIUllibJnjEeygGR/F9zL7vJSfi+skel3Gg8yrl07ogBg5fruiP8iqJX
/D0D3EMN9KrcZl443lkgUSb3aBzw4UT/JwsFXPqeGjLVFrH7oTOwNlM8s62gsjSe
AjqDw8R0+Td00Twq9pvMSSQM6RP1zSi3K6OuIy0XhPljlHJGe1GRVGwB6mIE+PZh
/0ErOgLZ5BL+x0J56AsWU711DFwtmPdDPbyMstfpGOJdOczjLwSwXpSCTk7cIIap
dm84+u5TtBGK84qTC/0QJUsug0zdDQMH5GbAkJvf/eoRyun6YLSXq+PlpAm3lz3h
ptaBfxkVhkv/rCbJsGpb85uAJXDJ1IpHD/8BOi06VTLUAtdZ61mk0fVe7iYzEPVA
27dBQTODwsa6KgyTwI3fgGiMFhywR75RjzYqniqw8LZ6WJBuGAIXj+QbKnq56sfH
b7FDb1fSqVpx3bEfJhYFNM5N1ZnCjPxMpvtwVL2oBmMD5ZXBOZs8hXedX1N2z7aI
ab7SvW7wSCrLC2aJ8LlXY9Fw7hwl+LI8Nxs6kKFxx8iSqL4Pf1/xhsUEhhBpBzld
FcAKpT2pz3sYBr6TmZnX3VsYhTgWKYXyxgibqKoVPoEQqFUDvDitM3s4Afcs2+J5
bzbjNKgdnOd+k8zlD4xrk4yG/GVqjGm2MYQJ29i4PAotHgTWojgd3UeSvXU8ausI
PrNISxpPje7kcDgZqL3D1Jv5xZH1qTWaMfy3q5SEpxEupx6hzNf82YzeJbbMVCwR
LfOmh5taEECht0J0fDzZVM6UC1mnY32N0qXKgr4V64+Nv2fryPMexhiaY+8F/KSF
5M8zLmt9dyLmvLNhXc6VrKt3E4+cgaVn4kFz1VqqdRoaRWrnRTH5asqlj2LJiTkG
RQ52oltdggjRpHrQPc4gIQ98T4ameYg42tswEEA9BnLuZ9SEdgq1suUyb68YT7LK
rKo7K1IHfCxJNkB0XzDCaWsaH769dr/I+TcFCZaWeqqHmEDFDkk9HVyWzdMi0BI5
rAXVMFRzpMCUdLe2j3Bgns1hl5JS7XE/cNCMnVHzRjbYs2/EB6sa8RPCge37OpVj
kyMEUZhwo143rEKiZ3cMyYxA1qW5nCqIpn/vSzFSmvBIiq5gcJQoVPmRlDtF/H3Y
SR2EErHf0J14AE/LrODeVAbzxW1mwchcMgPAwBiYW5XXDHCJtzWhwBbdD2VXhcAw
FnbLu3/w9q5r4I1ASMKQnDx7c9uAkwcuy6XT9S1PTyqZFxACtmENaHRjdye2RraC
SyQ/DqsPQ+0gF6OcpJVSJL7EjWjwTiGBTpJRJ/h4RcviZq2FI8b1KsQ0RcQF8y30
MT9F1EkKgxflvuJvzz5T75verp1nob1ScmJKXAdjCzp5lqL83dJSoDHomIsp/7Ji
dNdjOBlv18SD7104ZCuhWDKKaEac5XMmmcPSPAvUG+td8VDRkAmwSY/cdSI7aQxP
B5KEFSu0Rplp6eh4zl2EhAHVeL3KilcwCrioPCYMWsrAyk3kxTG09FwhJfP5lM9u
LAz37OZI3oZx1iP16zLEsKun4LVvN43rBqU/x9yiqIDS3h0ZPKpTnRBtLkE+tfgl
WqTHWZIThYbXu0Zlyj7OKGms2y/c3RDxKtBBgO1KkZUD7xxkvefS+I+/IZPKvcs8
zdgGl1gfUKOEi5un7nG2MijosnjLa4jNHqs3ojyAclaZlVSdnnpJK9y6i9ssHQAG
F6Nxfp3YKNiOz1R7vZii0Roh+t8z1iaUS/+EmmqZ7PmIP5k9GxxyPOAilogXZXtl
Pc1ozM41UwXC1uytBAYq+mzvXZQrQgvMfx9KUxOY4FbvP7oehBjU0u7v6mQB4yyW
XfSRrXwyLpE9Swo/UxvdEQTz9JrenkL7Z3NzDoA5ci/5MT+yjMoosPGFx00oNHRW
EA12Wt5mm+PaWzvqL43V6i20Hzfo4fo0pamn+Us4xU9lfMlePAaf1RIgem5NjbWK
5qiSn1elmkK7p3Ybv8EC4JkpDpX1hCi+N7CwrW3rvevJWb6CXGLeiH79xg97U0yq
6cZwUB745ClxK3h9SPqW5GyUZ6LXvZEZskT+yBiKM2M8cJXiEiEKZiXbPqOLrZEU
DnnBtr+mJ8J5Njipq2aggKeOvhdyHbN1mLM/YADrjUuZvNrvF6+rw3UUS1nvAMQt
e2XVOB2IG6riMmTh0NWRVVaWA66tG07iR1XSApbo/ySGT7T0c/LQLrBkm++z5kcl
GrpCeB8I6MPmUAK1hrXfd6KQEumtK3WhtqCxopc1ylLdfKJ71Ifgp0RBBFKkFFu2
Dtt6OFjC/APsJdAfHI5ll1E7t5tIZiBRcGX9MMzhbguk05I2ftzRFMusz7P4rLhg
vJwwKvtJjTqZzX9CwiZPVnxz+c95Q9OA95S8m6hnofoOSju+d3qTeh4Ff99VEDlz
2oIroTnqKFp66h0R7b5/xB1J5DBVGvVYuyCHxZgvdDVAUdjkKej3VmEHXh+BfyGO
5zkCO6t2h88qmNHv449cK5i5wdjGXlnZlK40Rht66XbNJRwRjUw7dE1dDAsdJnIa
ttZIY3HT6TsQLt3yyIBm9ytJtManklkDkk+JN9f4R5GQB5G54fnxJesvxl2iNRaU
FD4s5LxNqch6YJ98hJYH4ReC8/P+PC6UaYmefyJoBnc9LnSKwdrdHCyAFeeYlq+w
z+ucLYeXDnDUgUW+N7CEb7Qdj0/w7ph24EmTn0AFiTYABUOV6ETGveKYsiHghmi9
URLhI8pD9EeZvlsdUachByqsGmwp03Ycx098zbHb9b8efNtyrDdcXkN3cyHm4j5h
N0d9/Bn0s4xdxE5rP1BW4PWsFrHyx2X/57vokDts6VCG5PH8mA/wpXC90WPdd4Qo
YQbhnVzPiPLo9c/qpprjf+6QubOW2TDj+CoYsXbZoAhQyqTwgyIIxncw/8GLDyft
TP8ZnQGT8yjzP0gtcqvNHJZ/37WbyQJ7E0hUqpu0SY07jeoWEGkH6LHXfV/MPR1M
z2KAa8jX0+unoRa6tCJMkB0+V5CBDudOepvPGzvWFRk=
`protect END_PROTECTED
