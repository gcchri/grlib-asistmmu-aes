`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BEBMcgJg6jn3WbLNLdsZ4pHiBkWM0eL3PWSrwz74Bu+dcS0NJ8aOGFAkdi3z+tKq
QxZ/z2gle6zdyb9EiyoAijQzY0CNi/pdYypT0ccKWbTmpzkLh5PAU8NFS7Vu+0Xr
1BBSkltm+88ORz/ZpDqidoKrVhz4QsFJ89ZBBSJdUnJ28JJxHRsvTCqF9m7upkLR
kQQ6Gj/3+lvd+csgDAdgIdQoXpC3hGfKlyrLBA93CtA70Kejc0J0yjPbRlGNaAJ7
NIXcrFRcTtmm3Q9oCFGR0MpJbdcDmbA/XJW4Q4Qfuq9254sgG1EhwDQRNR4YwBER
3oOAS4QL5Ig8yUfXq3JDbIDFieKe6Irv3uQgL/FK4CyAGgY5aIh7Dk8ccCDS63Ox
9j6oh3wC9v81N79gNeUkp8le3vctE3AuTXfTlSkIeCRdES7ldctrQZdi5s1WE5Nc
kqcNisyx6D5KOnYA4r9bjUzBZz2jH1r1qsbVCd2S8YZzGmFzYAXTGhJFRjygDRf/
S1HrKnwnReGfnTRTIzabDnxtY7Q5u0OOZ/MWjfV7z0KKapJZGIPvSOZsEgSJlzd4
YXe5kYIUL31ZLY2pNoAeMpLeamLVWMu3cc8dyyG6sJ2j+5SlhQOpiQhQbf3y+DN3
sLcaTluxn567LFlpt9jcGBfVrYNn5qFMajLvV2R3vgf5yuuLHbuHXjiGCi8hd7PN
4QA6kAKooxVKZn0xIq0x1ne2XmE11eZothpuwjSmrAYyeSGqY4baiT8CLK1CEliz
HwzpZvW0P8uppIcs+/8sA9FqKwkpQ7bpEOozpT4S2Omvn1WqAlqk+7+vd9lLuTfu
9HSRIN1/HEgSWysly6USLg==
`protect END_PROTECTED
