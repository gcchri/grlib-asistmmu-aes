`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fX1ygo2en5wWvV92oqkje8Nx4tm5kZvBHxHvJiUFVHFjW9rReCWHDbEPefuku6uH
WrQUosYHgNOX70VHrHET2lEP/dtf18UIAHD/OoLvb6L5FO4jYUcc1A+PuuPlXuQI
jkqEEsxCVVGCvdIrO5lh0iQEt9yawnvAezWTYF32Ki+bjPv+w3qfvQhnzDXHRVp4
YE4hwf8oj92NjunZ9KpzO/I5emn1ShUFfhNw7sHsRPvZn5lLJnXYNHgq1rKzid7F
uhF3LILeJVtw8i4m0fD/tf28UlaMgQFv9u9nVzGDwf4DbvbzXXPfblU/W+FZ8gyS
E6gV3a3sARWq97bGrn+FnCvhYU1YPhz88tR8b3DZMOyKS6gphZhJJZRoJcgbyfU6
89ZFcB1HnAkBCpfZxHLElvud562Sz2ltjl25O9MdUiY=
`protect END_PROTECTED
