`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AJlVzPyXKYvxWU9AnkSqanZgYMfZmZC1PG1jmiHGZOgdQd2xjGWT3CiatjJ8l+Zi
6SJjsmUzn7FRbVdH4MFQyilHvikkKDWM/EZ29z3Ummi/QPLPRScQWzn/y2AvaBNm
mUS8mJ3C6x3QuRTDtUi+JDpCAxgzUrpKzn7HMOFl3nrY5bS+1zKanE2FHLIczngQ
/0O0Vkh67ITQLzpPehWhPin56e36KRNqZfVQe6gn9QrSdpC3Z275TJMQMAsj0Y1R
KglBqc7ml83x2PQsy9ff1BfahxBlJwNYJxwAukFZc1364gLT1Mn7Op+sNMMH7IQE
ii/BwktcVfUmDqs9RY1yOWB1eQ02pEkMsHXeYFBM9FMiTgkR7OHPBfwTlqoJYua0
c2bkVvMVga+uqPasIktRNS+/6/+Q1Imzzd3a4WhiNUkf1EdintPwS7PoJmDRIoDu
vq9rCzpemT3yP/y1+xgJSD+Ej+UwrU1PcA5ff3bkKWRaOWk83u6Y5jQxs3OIGwi6
9AE1Vwse8uKd0l22negkSJQt4ZIp6s/MjZrGU5wnuXc2GkEQic5rYeHBgO48mheC
8cXkR2Apizj1W10vAQn4wpLKtkHBkgnEo+HG9/YBnpIKwvKis2QxMCvwKSi07/wl
fYEvjrPW4CNNAuHrvnaQDA==
`protect END_PROTECTED
