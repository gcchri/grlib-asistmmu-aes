`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FAbsge5vfJHrNCrBlWus2WhVaOZga/gU3pD3pyTy0VjLFCw2uZac5WDgp67vB8v2
K8yIvjFTGsXYZot9BkwOAUl3Cg5y0Ox9qrphKY1Zflf/t3pv8wxDo2uMonP+SP8g
a1lVMJoe+W1Fbiu6pREDjxap1/6d2mTtiahlprHssv9dv00T9leYiELWHD4LhAkz
TtEzZdv3JCr5ja12VlO5hHc5FqPSbUgEcC7/JB2+LfjqlA6Q5DM+XN4J9RRIHZcG
V1HJuqmo26bOnKyqVrE56l3NZ41H6iC5xOG8HPUwliipePKBqP4qLIfriPJKhDD2
PJFdWJR9ZqIk0tzQRh1BufuX3bGonAKJosXGdh26OS94guGaDJnvlW3nG5cZEf2n
o3bp4ws/nrpGNw4jDbTHq6yN3vJ/Ymjfk+nlca0nqNeEiPC9eHQwvhC+k944yRMV
ggtGgIQG5q+tLYG8x3yLyfac2qXS4kky9fFUA7QzmZ/o9qVMf82MDV/1qylZXbRF
OOn0XqrV5tc42ylZLuDkK8Zne2ag56jAKWzv41XXiUWSaCNn2/nwTHK7jd5QTWz2
HVGfTYN6v3TAlEdaWmX4etTZRwk/Sb7n0ld5DbDtH0qAh6HP4v7BWN5zmBtdasbw
p14R+FNFlNoXckMf5sYuwbXj7hQZdSQNrqmSzKdD7Nul55GVAFJIHPUmo36WmXIc
PQqKKsRYC3AwthEeHabZhe/WBzF3a3sM1KIphCkQlq2w36sbj9c52rle4jKJMAJb
KfaYrhD+EcV2Djuwuw2IkL2xUhgDh2Fb5lEzrVjqvyzbIncGa7jzbrPGwHlW70bM
krOL1cPo1xY9AMX8sxsj8CDdQvVOKHC+URZtRlJNTwqjIJYy25yshrY9w6pw72/H
V5OhOm+RYcGdD0d1CZnZpmGf4YDiENeowHeG5Mq5/OxTrNgjHt1Y/smf9y/nLhOZ
j+pYAgar38duryHbMLGd9whC7JvjMx3U4vZ29up92zRIjDXXDSRXkmMJQF04u2ke
`protect END_PROTECTED
