`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vvdr5nfTlmVbxAjG9q1/41Y7yWVkZD8VZyieLH58zwNsnRjCSs32Iitp7tyHDOWc
F2sUe8jjdO/cdM7xbCeSchpIHNZSnIcdp7hh5JmyboYJKMk2blMMDP4Jl0oJh4yn
kn32u7tQ8PdkaoLCAyAZf4UG7xUIDUJH9lhVOIHST+ZbglAPZTqz+s7Xbx+yMP25
wGmUi+jVkvaQ9nIsN4Ya5c5VhFC7kkvpukAPJ0VuZrbOlnEQ2gzCIVXWzH8j4mx8
oRqGOji9Gyfn/7i2GXiKG3qHKmRVhKsMqg8RLku6RYcObaIowy5mJ2Bvj/RPaOor
5QpzcD46rRPU0tLVNXfGEDqWs/eMpYNf7VLNxjeEXdG9yBR/xA3d8fyqMUG6JmKM
Lqc133AmOv7auLB2c6peZQ==
`protect END_PROTECTED
