`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vLcgiqJLGQflLFGkFeLV6jHLLrCa7jqo6/FCI9r26IAJ1/rQQVB4ZZrVzGZpGv4V
VlGXmzYCQ2Fbi2bOsnPT8/rG94gxl2smxJk0YCksX/Akg05Ao4wPlRKOKBFytdNA
8m+IZgob0EXibgYQsxG8LL8nHtI1OShRvaXhV9gS4dve1UN4E6OfPY6hWqzm+e90
m3VVdduFK9jbWM4/Bo/Tac2q7jWBG2IM8c/5ciX3Qp4PhBnRXHQC1+SmXjDs9fDu
xXx9WWGQ/W2J9QKNIWTFICvBYC5+6bLum4BNuA4TcfsVmKL2o6U4W2fuGjejOyGm
DiXKiPluFZGMgtTK3HydgzaP42mZFT2zkRsQ0aRwX8fl06ty+DV0UXl/zQ9ARs/E
blxtUi2PvX6LnIBGB1sQv2b/HHu1lEecycmzwxRd8jrMRddKsROcbJJhktyNrogV
OHZl0AsB7RNOlkC9KJb04URlO15WHRHCrkna3ESvJnBJVYHOpm0aeOQyjoQEtfFf
ovC6GkBmDdTY8WAG4lEUvYCuA3YIaXFYYC5xGLFtuZx2IZ5ffdfSH8VE8KW8EDam
eYin2Rvy7WfURoab9OZwKesZwTujuZjpzTxvLhh7he1yg/owgqHC+9ZA0kS8TXzy
fXOlcEdmAtusx8w0Don0FmBz8HknlWopt9bHk3SqxYtgR2+3C+X+tfH1q6ZiHsmu
FbvXlj/D4BHfxJlK7txGGzbc6ytwFMLLyR4xRS1OVvHM/SA0ODjy9VeCv8nRHEkU
iaEH7CypEFV/p9jpSNBQPfLhNtAn67AeliRMknZkGv/1oLpFn9CA+0mGlzJPDjP/
K9kUJFb8eTuMVsjV5J+PC3A/9KFn6wrPGZSppdXNL2tbrfQ3HBzypLcSrnbLw503
0rudY6607y5Dm8vqJv1wgMHyDjxVErCy58B/DP7nhHe1j5XmP1iCJTrVxkXRzc5I
zfbCOKg/PzCV2qa2HluScXtlmol5snlTAKlkJn6YfPNrGYFQ3bQtyA8I6Kqg9MzO
+VUDtu3DKyaBkoFSQY4ogDItIpLpHpMobUb3UJ96A5BYob8IX65s+9/CDs6IYJqs
+Eh3KbaSluOFHXQmpBYPh/5BAfHbltDLlNiXe0hUakCCFTg8gHoWwCDtzv5Ey8vP
`protect END_PROTECTED
