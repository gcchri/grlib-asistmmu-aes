`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cvTuJZOo0eqAtqsrob1wJ8Qj+rOk9tmQ7oUcwEwzhRJ2R86sP7XnoQc1kCf8OLFn
0Wlug9tWe+nOwIEP3EsUkCiRlcz7MZ9uRvC1pai8eca0uUMrncrNmQfu5DRAAyp7
35e84GUbhl+Fymlt2A+CTtBEhrOyg5zxrT3p/Gmf64dRT8OoN5V2erCGN1Q5acIq
XMtfMWsBLADvECRiZfsoHAY7M1cZo0VrUkMIO6lFH/G1z5LoFTIHeU/YNsYjIBps
g6INBjEKnZ6PddAdM08SLwGraeiAfqfqD9td600rqkg7KsjhoXVBIPSFoeOE8uE/
2NHTqzMLlDYVAJVURSEuHI7s1Dx+JLl/6U7U49WSWmQE0FNfpgTkbmJUI4f43cJ1
h1xRl+qEcew8Ewb3WtWanjQ4vIiM0fT2igcE6APmiqNLwVm5CdcYCYGQ8AX579FD
j8EhV4EaeLGuDKL3xTE4mbJiYhKeg51FXP1ptYysX7QsTsi6JGFFBZBY2S6rxFoZ
F81YcUHqZL3upz3cx3pwkummDIwcMlSi/+un0NzmeVj0gPiAgaMCL5j0i0tXTGYO
MZMJALiBxSxljUvsmr8Yq7Re34qLONw4S9AFUpktftMSWdC7ZSpUvxFD5sZMyqNT
bkTXlKKbBe1w5XYVN7+cdee8j4bZELhk8yq+ezinP/lR0bsUQV3ODNfUy+aPGLia
fEHfBFOBv2RWx3ZhERGBs5neuq+wIsLj0kDHP/e+euDAXkk4H01lSFVDd+D86OAA
QD6vLMkV/plHGQaUBtg1D+7r3F6YO1nnqMH0W0fHUfW707MNNDczmCaur4oJYp+R
4xujNdEqAdZmpntsPKl4EHfjRV/Fw0uqgCajkk2mPAg=
`protect END_PROTECTED
