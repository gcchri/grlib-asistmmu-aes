`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PzH8/2HXlgi3C/40+Q4gJHkQL8XCwirO/S0dkRa5TL8a2I+TkLFvx9ckRERIskIb
aTXdeRI9UUOu1aE17U8w6Af4ZZLdkHFblvBlIEw/7Hxg/fsbtQokLNAbr8o52xQb
gl+U2x4yW6GhTy9cisn35SllPPUiy2yTmMLEaeqBMgk2JXvO+MkhCt5FPJVeHy4A
+bPl1nnQXktkBKMQbj61UkSDtXDRPLYncUHyFFYma0agk5E3JbkIdgGcHBxOa3VB
ohHAhmuOGas/DmtePfaA0F4Ieg/wLcgskBFr+lGtMB8qNF/64OQNc4W+YYftwpz2
rat0CfA6p03NEQdJNQ5BIAWqruS9zFe1DsKbHqYKOOVDnhcpxQN4wkSzvW4nfe5a
`protect END_PROTECTED
