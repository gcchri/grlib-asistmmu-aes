`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J8R7PvWkWHyPpR9r12lQtXNZjwfFEMJuKOCeKChxHOBvaIbxFDN229mdZ42BajDd
WsbykcxQ0yS+4S3bWDILJ6tyrA9NclUYop191CXs88ovUeV1I2INeC3HIso4YW7F
M/g2a+7e8UmbmBqOrDKxmT0JbDHzPDw4izS1q+x/0Jrmr2Z28vJDUgxhUOT1Xc1i
oB+Pe+vaBfaC5NhfAMVEgs5b22AjjAr96sMRdKh5z2+MMP1re9ucznwsKOtvSNWm
ltieucDlyqhhX3T8Yk68nex2W7ctvoyX9Q9+lvV7w+c=
`protect END_PROTECTED
