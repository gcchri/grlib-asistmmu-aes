`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e//EZPp5UamMd5Z8RzLBxD4SysESAbilC5/SSxePa2NI2THsbLZ844LQbA3Sxhqf
cRzDDzf+ndb85bLX89o1i6LqV8B8UIvawEYZKKV09ZetkQHkWAtcr9jyk3hSsyq/
Hq4X4Og8cP0fO7Vv3HA2AL+vwVpiCp4tJcBRVIWbiblEmvyKzmFdY9OCVeJbiz2x
H0wM5np//a+Rki8DpsgEkQ5QsVf5vG0bvgEVBYCsRCSRPAeYt+rpH46zXBTkG+No
aVH5NRG47BPiwGee2GEP5HVRuGRBdvEClG8Rq9CMNTV0k/R3W5vBOH9bD7kDQZCU
79wzXXBI7t+0QyQSTR4/jRf4+Lc0yKjnpW7s+JMu1gg998NSZ9/TAyqv0wdgwQJ8
rS77+iccXbmIeVaAC7IiXLmF4znKl/Fs12oVzcAeRJzUoofmOe6aQwTUuBjNvKmZ
fMScuv3OjXX2SNzS4WJDDFvcd9qWZhA4nwJ4HJVr2SxhU4j2PbOZu7JfUM28SqXN
`protect END_PROTECTED
