`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vOFx+MmkUbnp5aA9nJXXTaGQqWj0rgiPImc8eWz6WI6odinkhB2FDPNViiZH1YbY
11DTxlqhpE2QmjeWo//cbWJhY4z6MY+UPDpP5zPQXOq3EMols14aNt3qB2xYiw7o
SemBSLQO+sPlK9E+VsA6KmP5maSNJreAkHrKWCiZGgR6TL8LwsfDMFAHJXrLXiHn
Om/VumKoEKvd4DROQA4Z+Wq2KCcIyxpnyk6K+Zuy7GPAlVKAt72yNEdz/gx1+hbD
vQ0aHuAedahumTLbsay4PTTPysfaIIuPjDbPFSpapFo=
`protect END_PROTECTED
