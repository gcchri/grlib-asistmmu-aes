`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TZpofXY7Tdp9tysogfXJmohp2Yvxe0PLjd2UI4pPZkrL8tpcRbHD/XW8diX++2Tv
OejsNdwtJmfAAEBDF1xuMkV2JXBeb2hY5Jo3jBdz921eKWeNx4ASz+Fprvkeib4L
ROpEJ2uK0NmBNfGJvj1mzSX09Zkm47IRwGOeBNw20Gyc6a7K7KKMd2spcfbmwWtK
fRzhe92vGu3dqr4Zm7FvIMFWnCLEoajKwwchyPoWz/TWCopmdXfkLyEzOYGqrwKX
OBfSQJjdQ/1eWSZoL0lPAiLeso/TdscXOyALEIYRdA2JUxFD0vSBfXwc5nz74WuM
WyC+APYELPvF4oFziskZc6Y6QgZlnI32r4VzxwSNFZ2klYJZz/bKS4IyPvXzUM3+
FaOZuzcQCs4tND8dQEALBRogERTa1wc4C7WvWWq80EbQWG/4y+GZekYMtdw7ftMB
yVxYUtx3lHKQuv7MgCctFMPYDfMsVcolAztJ+Uh3Zix/kk2p/l1K/5qMourYNn1W
B81sqnTr/sWlDbR5cHH2w9Iy3UiB7WLjk0OGVsAb8Xy1+edbJO9B4UeE+3qfigGt
2ligJMNLfbkCqhsFo7HsV1jC/E/2sbayfRjLhKyJBia0tY9tkPboQnkmcVYojdJd
ylOo6VS23wNsdKBtLrJn0Eh/JpdzOcsSEAKo6Qu02pYLoPzVjaPNoxsph6+O/d+7
U2UKMzyDI684e0BY8GGU+rcvexitSv6BIQrXIVvZV5rL0yE/LoINPePcsIMojBDn
hN/V+vJpV0M4id3C7sG8RweDF0FkijZZk7MZGWkNtPnNSBSRUWavM+hn/Bu9SHyP
+smDJ01J/vrVgpFvmKbDO5dqvgXh3Pc/ykAJcZ8ArD2iw+pvL8TR8AT6eGlbUigb
RCARx8HaQ+pysrWD6iUaN6z67RA753/DV9kOqccgc6Lh+xXk0GJkk8K7Sp/huZvT
fJuYWX0ik0L5+0WK/sY+e9F+TCYkZR6yuoJ6FBWq/HIpwxt0qCEMOhz5XpFpsHki
Lj2nFG5Z/r6UVAcQfZTvyQ==
`protect END_PROTECTED
