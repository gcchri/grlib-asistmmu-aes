`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x5XMHzzF3/5NMfletHPHecs8i++F4VGYybx6hOrFLgHPDK1RDtDLsOPCjEWZKu4X
wbMuO8Ie/H+iLE+50fNiESVxN0FveQkHFSxL6J9fQAwuxFZpmGz6pKTt3M7jIzgp
fgG4qWYWEqdV/n1MZbyJPuDpnxz+EXvR+Fn2tiDTyIcROMt7QbS2nBCFky310+v1
NDLvr8IjPaoN2L5goiZ5fZqyq5FQr99Ep/aSiBcA3E1f6El8flNvC6zQ5rycVtjc
xUhIv2vKwNPWiEPZb4wjikzFlpGsRF2RDQBHleGiMW7Z0OjW3OGG209xeJSNHhFn
FpRPYQWYbnxHhTAgUvb+oM+eDNmkFf10zxJBdiFKWV1ULEkwPkYzpW4YJupWFtaL
OlCEDdD5wEYXKvZ33Q51JjaSaP9o0YfyBwxnU6TnOCY=
`protect END_PROTECTED
