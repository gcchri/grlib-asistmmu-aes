`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bdlYKNKbpN5oN9ApEu9hyPjdHX6yiKY8ZQeUBXOqGZ1L2zIjGE25A2oZRSm8aPjH
LHKadh7gimlho8xdsroYeR+bFJxZdocXl4N0nCMIzzXpaPjJxwQD3RxfaH4p9PHx
V1zzGAE8qJIP4y08EDsFnHWiLLI3y/yUduNH4F/taDU2DEkeAUp6gnF2NlzJJetz
gtTCkhjABcaQ5uJll1dIszhVAVNY+EnI9VHSjoIQdA4qW90fohRmvGuDryfP+7xG
sXO0eto10HsTqcnd4vbl3iCTnuxmvlPRUWflVbskDhgOUE8cmqWlpQS99UYusr4W
sRFSZWXgH22O1sQC6ZIPyzy2f/gP9FBKZlG0p9seizxNj68JtFDWZslRdNSuvv7z
aypZ3CpGwf4F7ZsCkssbMsTiOtByia5dOFig3OYOedoPQzBgjIVr7cGsLWMjd514
Ci852QwYVtH4YUK01wl5WviRn6Ra35mlblBO0RxGmJgatvZyO08TSZFO4+GM2Lbb
TiS42WZ/6PycqY32+TiUag==
`protect END_PROTECTED
