`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lL7fPKFPY/apqYKFkWZ6h/rSWz8Hli75AwwQfmnjdjVBqkw6rOnicvH1fcQQCuT/
3Uf8/bEzHiyGSLmHkm3qInx+ve2moMyOCujKAzKDiFlvO0AcQbfaXgSUz2IXLMM9
BFmyjmuK3FSHzOLOFb7PblFa3FjFH4F7UFcCPIy/3B4PLfclVoGYWfAeHzDSfuKZ
TIn6RsVQNf9lxLkkomuM2KFqFHtbUUh7Z3//S6DD3bNdtwfDsQLdMwMUWRMBXOj3
e083hOfgj3WT2g+HKrQ0tnprSz9v3Fppr42+EtxGh/U=
`protect END_PROTECTED
