`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LOhzUWIbR95Md2XvSmRiXwxd+Djch7BCkaOVAk4dgGGmiijdnIRQAHPqmkzJnfT5
NUo3Efyk2nS4vI69RBk3lRndLtcpz6zXaPAHz4srMTUikV3O+hmdGHSYRVVJcTki
/yLdM9lRv1XtxWpEhvI/zQjEcpHAYNVAplBC8NNTE8sgKin78ut5BqQLjEroZ01l
Usc05ufkv49PgfZGMyHDKJDF1fZCJFSiSX3bwcQo4itomOagAxVVjXcYMeqR+uWd
o5yV6PVxaqpVo7HzqjRgVjRg61Xw/pd1kgj3hqI/RDnBy8mzkx1S+qV54ZmMTm6E
RktsdL+WbzIMznkTbWnF/Kdzv1izsxcWj1bWGuwzkhdibQvbft7XVpZdaXax2Cje
auR+PPjfIybI7f9TntIcW+hFe2gbVkF3WD+4GoozcM4ZS+Sve8NccoM1wLRvtUTF
gj01p6QGLrt2OTMhuLDbed7p6T+goOElYtH+ZpCofb0H5kHZMJlK8qBfC2lSfpRX
UHjJ81vO3Z745cn7M3lGcTq+1+YE2RadKgeaJ7xLi3v60K4ZzqoMaUX7PmN8QLkB
V4PV76UHDoHMlqjmNnf/jmoSsJf0OsFH65RyHlLAuqcoQX/w3yI+/wpTb6BUP+a/
3tRiviCGfF+vT3s/KfK2U+9I7oN1WYGTpRv3jzZuauZouGulQQd5xcGgwHTovwNj
WPhP5k5ttVVMriug/0D8n+TLkU5QroqTsriA7oFhvjsUcZGcr5ssGEb7CymuaQ1U
tbncL0PGkF3jjJl9boBCZMzLv1d1iz5ChVEN4yWUq0OhIWOLSZfaw9FjuSXJEDOx
pDBcCV3ypWdBzCBZuUilSNxTjT+zNv3PucSrGH3NFGgTfJKTpvS7sc59zcGsvQKW
vVmiEizho0cbFDBr9WtpofuxH7/cOGR5By9wFYZcEro=
`protect END_PROTECTED
