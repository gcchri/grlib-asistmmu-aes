`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eMWVXaYK3W4bnnD/dJ0Mfherva8/0FYv82hD2CTJsqgyw5unv2UTN+LLS1r3QbRu
INt0BFsfTaeC/ad7TRnU+nwNcO8G8pApZDBTJXjHcmZTQEUCpiXlfqN6fkQ0DVsY
TgkiZ0XClU+lp3gqcMtJohMJ7K7grMANjcYk5Y6hm8dI9/AQM5EcdbnUk1wBEcgf
9+FbfVHKh/URNM1zSQC5ZJe6fMfVYAviHdRowaNwVCjC1atSt22+7VbUUulOth2B
BsnM84hJ3k2rjNHaj1GYmXCb1LbYkXqmph4eXtMnUmuQgLZTQgiXkbQcTArzGtLb
LrGBQLvDdk94FUmMloABMoZRT16ZV8fxhhxCxWcI/Su2hFFkvRhs1UcS13CEDlMo
1lzXq7vdsm6yVYRoyN1AEAzEr7izaUZ36McD+8+Vs79SrqXyAm07FF73HcxAxetF
dS0TmetYs01p7vNzEqkkdVLO9iyZnNkL1m5VRYJnMKrN5Cyxcs+gFdjWStFaHrah
jqTVU09WnFysQ3jncz1u/iHTyBTnHMMZIBjvzO3yABxcaCQCh42WYQil4A8NO7wq
UvLVMqPNGwoEASQN2OK3XGuRtJYTCY0HqZU0brSkFJM=
`protect END_PROTECTED
