`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ms+DZViJ2LOljMVmBsM0CCqZQMOV+Kl0aUwHlTe/8lcKUv+uMTMLh54iML3cL5Rj
QViS4/1JNwHEm0piLKo+Lf+GGJXqKoEHZgbJDpGeOHwJqbFTlpcNJn5EYxgwRDSP
zuHu308fMmFd+i1u9LeeD/HTk1jj1KGZrHY6PUVt8SUi8NvYqY5An2f/+L9eygIV
Qb37n8RBDA4DvBnI5S48ArHHPVzpcXs09dQ+aO31I2pcOxsDU9zFx8XLZ1pYe9ck
AnUav6D90SLSW0aZkkTN8tBXsZSlRXmKd7xNJyFmhjlwbo3xKYd4jhLfzCbyTbO5
c7PwAjipfoSDXJfZ9zB94X+oFoYorlAX6D5xK5GRRRMPBk55LbhjxJHuozabbp9T
DAEMXB5aJ+dwHnDODqizFw==
`protect END_PROTECTED
