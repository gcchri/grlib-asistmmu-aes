`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lDGh2npI2EOL9aXvDcc5I/YIWG9kk4SghGV5bfHHw5kYbfqk6fV1uWaKsi+2i7xV
ETxrL/vpq4aJ1Q7m8ja6YPuit37DXNCujt0EmeWedhRRQlQLCrOPIbuFwF+9AcYW
klX5S58+QNlCpOcx9Aa0sTY+JaGHnWeq7hdRHXht1LptKL+wHA461bnieS7cBB+A
E2nlJ7AwR2gF7/zW0m+tooBd9cI/Rii6pG0L4FI4BzaffnnJEdoxZ+ShATyokRRZ
hbH1f0+1iRMlbC2yh3Ni3Urifc7ekjmKUQhRuP0jyH7yISO2yzb8IQc4VueMS5oI
eKomKOjYFNmH0OLTwz1QBzzMah2sDZrElsy/7B+p2wrJkUzI91/FjxpWcs25x0bq
NVec1RQ9mtfBykjpJpL3vQ+8T8PF+MTYw0MxmM8t/voecLMoPntvytKA3SZB2Pda
0bwEk0wQARmHFOpUcgFPYZX/rbIaszDrXKKeQ9atu7a8aap9f3dzTJDq+pq58yrA
XhjUJuy0qSDUcg6IhHGrIX/xIEypp2APPMJlS6TNnIiHla4T1lzLQWn2lyZMgYRQ
I0Wcy8lyWhfW8JniPvtl7Q==
`protect END_PROTECTED
