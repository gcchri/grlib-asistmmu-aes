`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pmxKoMKHBhqIIaOJW8L+jTLS/UYnpot2T8FHFcwDfAjRqzN7GXWXc7A+I72FYfbq
SD88GV332pI1Zj9F3lksP7jblR2snoszTixEHYOOouLEl5SRjddiNofyDmFEmqQt
GrYX1ryIdOJn2EEOrtGQOeVPW0ssC/OmFS6pUGaKLcC86NyAbucIaejZRA7mA/yk
Lp4WiN0WEA6t+iGGSHnMRxZhGOd1ZTY6odUlIicLw43FIxUq+1Wd3fwN2WruvTu0
AdFGQiEVdCoacAOoy4x+x4hrEc29WIDdVtPvgIm8M32I5+giMBqbCk580I6I0DYI
X/NDVWMOwAN/DUM5PqJzj1ciD39OZ8sVuKUm+j4mOXJtbEg3pIwkYJyH8JQzMdhs
QnV2kdY5l7oSDseczgKVmQ==
`protect END_PROTECTED
