`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hjudH8E3vkpQGwRBFPNBqg8rYH7VCP/E1RyN/4amdzMUB0rrVe0OqKaBnIkkFzpP
Ii8vkRbJ4KF2fqb28q8zzJzL35nTf0a7Fxgn1Q5METZyNGB5xgMc2lWE8Uzg7Dl9
Vw9Vvr+oHpgXe1k2ksb032OtzcCb8ddzbluBG0Kaqka3VsAdS3tgxxK4aCBw+MKX
wB73lxSxHRgkP4xXKpbCuG6sMsGjRll7dmq+FkhRx0GYfIYWhvSVoqGheMtbft8J
84MpR9rAJuEtdjhjHEVaRbbK/CFqEwC0Ays4ttjyp6jNtPW/2weH1a2xEJjaA/i5
zsRLsIYtxwOsBISi1/hR8DJTzj7lbwdSygT7j9OnQuOta68I31M0gv9eAWcAjlNF
KNv02qVp7mzzSLbYr9iqVflyF8B9xEFRp57PtH3DrFgoyR02Htcjt6XyxOwYoNtG
i+boZnf7MntRG59StBM05MFFk/+UKwU+lakVhC0B5QTEja1E6GTl2hNUpTTn2HR0
TLXpPEsGjc42eSShuvzokpVwXQzBw5t3MrGQ6c6/E43noGuvc8l3qR0AALwfjKkv
jBNwaCHEo/Z60CtlMFERx02BkUHn1yaX9uEdwLjNqajbPW3YbhWQ1yqVT2HpBEOE
EGrTBd00fff45CrOYTzRHJD9n5P7pdIrjApsWyvD5kU529f5pM4D0EXWq/zc8Isz
gNlYwGZ35vP0go+A15KrJKH0bCyB5Q2kbfgcyXw5qzWygBUni9AdpDomXpv2b9ZL
AwWPhFkg4S/cDyNdrlqwIojo5YYX3Y/zrvrnzREVDMCsfHiW08t6c3d4gOHGFSzU
KKgtyHxaW9nZk69VrQeH3Gf9MsqyeHQxgXcS1bODCDfoePCD8BXXjBKP7N5HMJXK
pNojJ6vjD9UYcskkHiPqst+mG3Is5zyu0jDh7nyEjvQbfzJXVu2vNl9kKZm1oWSD
4N+8xCQAtZ8sdNE+KbNC5QfZP/cZ1P529Kj3+CeQBxGxWS4hLRtVArN19S5BavS9
GNZ9+vfJ1y6CwL8HuiBbbmjTOLAC+rVuYoMnyVe4gNZBXugoEaRLVutPNoziOOat
x+jpUEmlXXWTvnsuN6vRrkl/XoAqCDkXBohTGIhbf0DGSBtomatDnJAaccQ1gvN6
IITUqbFqgN9cnic/9jfc7xXxukAPB78vDUPfoqhnZVthOmXZfd7/Zkp6W3evsTIx
eqLZC/gGhJJVj0S1rRHA2FDJ8ixoaKpanzpbspt69KilyPTkLgHlIg07lanP/Yb3
fLnRRPRbe29YySi4CqD0jn2o0mXPsFsAtlGU4Za/KBpZ51UpjVBUhxumJnACLxhK
G8RGFfsDHRlQjmjHKRHhNVrO3ye773SMAREZYBD7qUXPoszDbxiPImQRXPryr7lf
+ajfekfr7Za90oQBi9bD3OIT8gTWcAf42spKAbYGhINkOzM9gZM2YPWjTw3Y8Ucs
ZRqpudN04Kp2we4Y4KAqddDTCgUFemirdZuS4VOA5lH3+lM32aCE4eZUMcPjZYNw
O123GagusXqqzIRTHsaNPt9bP75U+ruq+7y6DIeAJbPissPTurE7WWuFp9Qr1qAD
zXYXFLX4C8PABUaSB84jufdFrrOUchAwqtkCLQOxXdf+Hh4Vx4o5N+OlgXGnXQwE
0nL8Iqpsq+b0ySMSwp9Tth8g0dUSQq7X4jVL53/ONizE3XAA5zEgwvEqrzMabJOW
nAeyUgl2OQSHAYQYEw0liXmg0lY1ttLl/sXKjb6/fO5oudWfyv3M2DAz7Nc2GqKD
MzwROfqGCj3Qgerc3hyC17MKj+MLNdG3hLHB4Y2dncDqvWEJ//rn6XM/CM9XXSNx
RqAnc1HgYBzvHhrl/7KNgtLihVuX4b9dDhINohBOuv0t7JltH8V9H0n0Q0WkSuMz
ukmP8MxTYneaq6CtOaykWG/hYKkbWTWF/9am2vK6lUbDSSBqP5wFZZBxGv+V3+dB
mdr3uNLyXGu02IFJcWCgL4Tr8MXc2+cINb5894vVyQW+jQ5Azmcvg1yUhLiYac7y
wZwqhzk4Vr++ccxP03moN1P7rrtmaNaNbUNQj+KaElI=
`protect END_PROTECTED
