`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bpJJIkq0xbCysxJ7s8V/TLV3MKQJOsCnCQWuPRLmmcDkfY9rJMK6W2DsXMybfQuC
Sh121j+0Ruj01nA0d/IXrX2YK6RLePll9pOt6SaXU56nMHr0LSc8RBApzeo6h5rI
dC4v/i4OaLNXLcQSLUgVGYOq314ZL+8FpWXWPIzhUvBQ0SQ0a+H+0mSijF1X96WI
PJTq6snM0T8pVGeF2i/h38TpvLmJVFa5lrgwm9rDk5wE8F4ZCps/aWm3ZoZqU7gq
MWFnrxWgK36XJLMDU6O0++OOz+CGGPLT6EaKZe+FlSEzUpeHnIa3VAcq2NV7+03Y
muWbUNtCRtU0PiP7OqIx48BYVTFItlOE2rqdMs5DAFkmRJDVgUjd6bwNY9vNDgCM
b+jPKR5l3wAG39XnvWabjFJRDliFgKcMR4PkkegBRFDsYfQU4T8DPikrLMCIZu1s
5NHLJIOjfmz7dlqX1C20Wy8pf/Bpkhy0kA5ZCcb7jGCQQJ30yTHii9N3nRJEgECg
QK+pS7meCsenZI5PGlFPwIyfn1OrEtJhNo8E7+D8gvGl+b+vU+qgqzKifaRo/gkk
GAAoZYBNyGikwr493VJ92qrPaZGAt+QVoYbBuYSryYcvs2Aevc1XhsfOyBeyEAb0
10/lxo12pOGjcyts2q0a4SwKCriBnwWHCSNWx81zk9dSQxTgs0GsvVWIfRKySPkR
z14XClnPTmdKJaVr+oHdxZNhP5Tr1vFnKOxTqEoNr95lC/n84FMaLBq3yQe5Id9s
O/CTnO6gJePJCkHl6CcPuAdaBPT1rCRwJSMkeZB8V/idFI7xibjSvYTgtBbtiRem
7OSNNoNsfontQ9h9kzD7hYpGeB1/zkWyNJtWwsFW9vw=
`protect END_PROTECTED
