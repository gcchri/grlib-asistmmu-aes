`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9WvyW3WOOwR360yTVD16vvBQMg8axEzerzzR/IIbnDiZHhor1QvifKiIzzNBhitb
B5hIOsZtsWvLj0geQDvqdlMgwyOGu1gabOLbaMIB8WH43xGoaCUMciyBdP/0tOgV
Zj1iUla9tHmkswaaotzRja/36rwhCkR+iMe+VRQlykot7T5qNaiqpGLiQh/QCobW
q1Bj1h73PLfxp56O+eXYjOfzx2kNvlsncWnk1V9jguIULVgLtRuRxv6VyIhrgd0U
YXqAeZxpxccLr51WePUodg==
`protect END_PROTECTED
