`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P0XFULNeg+9uyYN5xz7Y37wK7rn/lfoU6zSs2C1c9x17LVyXTCNY7xEKBTzBO+/k
n1cwOzmPnd6daI52ivSKnYoKmXHb5DxrRwBADS2oeupOuSwSCVDtMIOy/XlOMQYj
enTzlGfBojMynE4Uh19tdP0+ocHtIVFzBoxNHcCEx7DMGtmBLbDPA0muEVvZPbSJ
ESI2gwHqgrh51iGSv+XWl26XnXdL4W7PE+ZD+OpsjKelw3HHC64T9DSs8efhbEeV
g3w/l+PV6WgTS+0sw0UOY3YVfRbWdZLlZzPZVxzLqD1gY+K1RrKUpZcqGkODusZ1
DB3BMFCkDqsWLshsc/UFWFFvPXCK7XPoNRoLGRUcbQjfKzqupcOB3M5D+aTAJpu6
zuF3JyeuZ+GU68br18a+YdyBzibyGYhw5uIIv8sMBvyvjA7fJruIcltSb93ORTAk
Ealt8OfoCvwVTeUmHehMU0iO86C8PyjLKTXmRBFV7Lo2TZQN9CCF61aKClr09YP/
d3EwbRXBfrR/JibdCxwQ5GRBFU+HA4oUEm/L+d9w0jY3errGVKPBfGUvxET2CKL7
xBJLSIhbzMldiYDD7zQgkZQEgA8adi0BHnj/GoSyRGmLsZUxLvytmMerUXC47nnA
Rhzz5pGJdWWYGy+Ut8TZhmbchxOcWoebWG2AMtGKS7/ZY2kVrD1ASQuGJ0r3S+Cw
Ys6F2IRkO7tpmJ7KJE9H2oC2vj/WDdKbYEdQRFxh/71gXlFgxRHoo/bRKQTzGsYh
iFLCRLO02NTI627Az8PewnVRKMqSUc32fkSEjs0cZ+yFUFuI2k1x1kip9E6lZY4N
TT7q7rveVV/UoLeKuFvISA==
`protect END_PROTECTED
