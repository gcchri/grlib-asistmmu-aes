`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0KUJJrJkeLGtbrux2ns5Kp+375LOVxlcJXJojeJgdTXXRFiIVQhPG8EwDDcRjzM0
eAZd/577JzfNrHTNReUt2K2AcjZJ9erD6hqIum5ULw6JzipKpc1tu1HhAZddVENH
SYk4eAWJjOGuCx3QcI94czkfBLVSi4znYhQbwHCCcrC3pFbYQQuhH5QEAYCqL6wq
tLEXkasNbEHVz4tujzbJ/CoCznjiG2Edaxa72mQKbV3jFdUA3TS3IJsJ19C9V0xd
h2x2EAmGwMtlZPuZNWmwvuKpfr8DKVy15eC7S5wcGLA3RYHY8Upjq2CyUmNNIhz0
o19DPhmqSyAa4n7pPCMok0eNho9/ydMuskdD4KQkF72Z+CyetI/+3ApWINM/Sqge
qxTIZ8opPZvu18Z5B2YGgDJ4NugRnQCbaPnUY6pK/34=
`protect END_PROTECTED
