`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v2MOYihtP1NaT8NMbPMkfeI6LFRVfgy/SGi1wFEpHsKFAQ+ytkUk4tbHvc8wspcR
++z8mFpirVz9uKGCF6XSesaVohvpDAcGeibRKqWZ/LsyI+RKgZoEkA47nJXM8a4E
tMNU0b9MnCYIWeqBGYrQ+ITVnkwgsc+DnTlgRHgvwWveuwkR+idLZFESYPCNxneE
wBjOtvmwfvwlUfwB6TOOyErGyr+GU2df+3PEwbBX8vZe754ADlX7kp0nRTg4hkzW
EzHlxzv3dCyvGOfSMRW2NQ==
`protect END_PROTECTED
