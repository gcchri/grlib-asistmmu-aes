`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9xtMxJdSZwC9Ixj4yGGNfXriiCmEP5IzV2R8/Z2dBrxfdmtdX8zOeTeibLVlnU33
XXdsWbtlsTuNL0T6cB2OwgD8jTdwvqjkrvqp/5QWIQ03hWB3fBgNLgWgkNgv2DHc
qb4hT4bLVUQMKMz/WP756DoqUu8Nlulk+KoJOlwfIPJ+tP1iQDJFD4bUnWq42fNr
DrJX3hSiVWk0+nt9WMgZeKfVUDqhLt6VWj3OB0KUNVOvmGTpnGT//yPPMyh/Xg++
0/thj+c1w1eOMK7pdRJUaFw2qQPwBtAjmyte+QGT7BtIjJMhqtEP5CfaU3A6vSyK
kH8Fp0+f+qS/pGkofXS3czqjLaE7/zCt4PgAwPWHwGbrkjlG7xg1O4IyiBwZyx4m
xym9YZN1Mj1MVuO0drdYOg==
`protect END_PROTECTED
