`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ycypn4ZSsbiBW56k8avBVuo2Zo092Zvvnt06FkI7SuQDGvrCUguuP5/7WFSOO14t
ZnvCBT4Z28gDe9Dd1DIpB8eN8yDjK71AuA3a8HwzkakHvx3bpr9NRh7Q27rtyhDA
L+QMJj24QAT4Ys7T9TDUhT+0Urng7uavXOmgM4ROnEJ9ea6WDg5tNGF4xZMX+wKk
E2u3UhywnzP7Mu5PyZ+JB8GwKXscjX1PAwt4UfTUeWoNdDiXiF9SjFHID/+Se9Ao
UQ4q06PuM58QcmG85aR2c5i1zC/YH5PGdf5c7f7BJAnrmW+RHz+vf5Ob7d7yX+v8
A4lOxe3EgMdv+3jf9Id5pzyIpeFo1RP72fOxoLFCiajfXmQDZ+TZIPjte4BOSFWv
hDbOmJAOShvv18AXEUm2uIRKZa+1vJLoikgDHPjY/jetJQgKvWRG1tr1ZqwR1ZHB
AylqqQJycNeBRI2JBntOrg+YobHlA0yIRAbMM+uk87YIuxa/MdN7GtjbKu81aJNO
pZdQFSU1xKjidxysYqCIP2Oh7Vkx6wb9hqebfvUakjfpxien7MRL3wTpMSJKhKwi
GZPJpqBzHuBzRXkNJt/7mw==
`protect END_PROTECTED
