`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5M91T+wQBgkGHIsApwQdMz6rfKroSxrzNV+mbZuRqRsv+Ilpi86E5/TuwcL5SaZ4
nrbu+407afwzuSchEMmoBrkHS/Gksum/Z/hyTdr2QdQr9J4hf0vabEZzACn7vFvc
N9z/Q6QjrlmEru1x6Bo9p4ON6SAnzyGDIDu5WExyklkKGVJFU5sVrzkS2xhH9dOx
jem7U0/tAj0f4kzyEAqQ+SeWuaDONJqhUXqq7olbKdjaBsbrE9Qhw5293qWLPY6Y
OpCIV8n5tSUNitHrECHAkAkL4RM1/zeBqjq9/7tywWvee4lPc8ZYGw3SwxgFO//d
VYcvMsUxexCfTke+RoeUrJ0fC2goYQK0emHRC2TyAhNLwmI+/TGsIeWKFeSoJChs
aOq1/4mla981RY2sT57sxp6tJ/5qBq3joC0hrYz1DMgrXuHVrJTMCxIhy0vShjEI
k1UmW3+A4ad3r5TWE8A/Q6UOz6i7uUG4TIoMZkn0jWE=
`protect END_PROTECTED
