`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8FrsqQZUkexz2OVCEqNDQ+AMler2o/WKV1GtukRjQe2DfbOUsR/lEwq4mE5LQxZW
xbWKHsqkNQrn9+DuAw6WXWJUdTr6eCPkIj+fQ5K4pnQTMDbYJe4YnVS/VIBGv0r1
c8CgEFsMiKf4n0ulMcpIqhm0m6VJe+DyDFz5h4WBGGqB7E5KICQY23lgrdjra+mM
ghfZtcfgxfdLhFTnYVzxep9Y6vg9oBBGKDaDqeCEioVROQwjfoUFQsPKcaT87YpQ
7cSqnvmaRgNETOmRD7dFBMb75YJ78tvoay79jJnOj42Jj22QGRhyY0B5tWTw0PFn
e9Jn8LE46ozUIzHL4cMeNhuTpBlyXqG3H9K//R3LLVwVtJd+s0tCxv7HJtksPAwE
aek5YN+cMa9UGejdGZdJIw2nbKaJXvD7OjVNzda0OEXS79c6pYTkCNyfyR6/OnlP
m6w6NNnv8piuSYMfoIK9qKORumK1JFXWYsFnw4XxH8ez/yKzNHUAMrtzCk1P27KA
GPMMsUfDDPwg9wvmhY1RXCvYUchY3cvAXhQuuFSjuC969wQhADUPaspydIrmfJcY
Ni8aZP3miHkHDCWGN5XYw/mTF0JKGMLlBDYD4bu/mCU=
`protect END_PROTECTED
