`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nXW1Isd+j31sm9sTGL4YU97ApllDjPtlQtvqfMTgkSJYh4ZjqzqKEBdyREdPLBe0
auqZTmJI/CfRaana7yCpc87jyIHwV1zmfwxUZep/tmsIiFAx+3QW1uNmJxtR5fVO
Q3/QAuBXu1wCS9nUObG+IsF31UQrEVgzY0/RfnZW7Ne4g5UTRTbekfhJK9bseCaW
2S1MzY5oDQE26iudHwzn21T3F9QyrkLKsWr3YhAcnTwgWbomTvAPSwbT66I51Ctd
nWk4AMD7j/oHaNcgwUCOM3TDc8uC1CeUk/r2R5LmQmY8jfRLZ+pmINTx6mPKVVI/
0iXEn8M9qZYkmR9B1GjSyoTLR2bZjLgiMR/LDRygIgUmvAPOX/2jVf68Ju5cBTT4
u2TlOhqIu28B8+uLmem/rxogD4rG8zpLm8nXS7OTndybWR6LVcvoUZUfQ5NdqlnE
5tIjtwMjjiBMk1CSklbKV5YZlb4Asw+GuHYd735i7/A=
`protect END_PROTECTED
