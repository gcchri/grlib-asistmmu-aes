`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h2X9FSY3RtBRJec/5TdWTDRQJbKDaYiRBsYSRhGZuuItDwd6yymBZk5YVo86/75n
1XkgKbRu+G1K/h8RXV3y4IAAL66fA7bjZavIDUkBit9l0rhu4TFwa2lRwushumZa
zl6dpGAjSHhS1KpKF35k09ORBuXOzh/viYxMrKB/mt9GpLCn7+cTc4Eep4AUv0V/
d7HRlc9Jl6yPTN75z1bZOX2jG+56ENCdqOtKP7+MKEkke/sLk9gFrKznqQHlRL3S
cZfh0EKWlovzLJKC4XliDCXlwHoMvfE8wvSK2/GSIES+pY4PgYqyydyJAeC49rTd
WrGw3+hyUuipv2FWQUekNmslbGri8FoJxRvS8EEw8zS2HxMTP1RAQxTq4GthumUk
3UqeS0DCK/f3HMTK5WSjCU4/qBQ/OVyf9dzZaWmG25Ymg9zs0/N/P65x8ZgSJ67S
tHUq+t/Pt0SbXGjvlhltnKEkqSY/EXtiRYUyMG7lKfKOPzfJVuYvx8ocfd0U42vx
61aOa6rDqT5CDjcuZ/zh29eTz8LkW3oKQQZmEmvo0Tc4oTnGr59GEj2kU0mAnZnW
+DJ10TQhHJe7zOEnH+MqaOlQYantcG5ipTsaOA5lZ6GvSPYFB/CS7f2flz13mPG2
/3rmd2INiDzhFN+OvPwCAc9FScVXtHhdPHYUTRQYW2Fvxe3Cg/CwY6UzfycLYD8v
0Q/VxE1Dyh2dq70lg6am2RHTjwsXEH94wuq/VAd+OlXM77NuW8ZiUh/BzNMHzhpP
akQKMni0e6TOptHZ0y96JebrQCGChTa/27CzO4slnAjlZev8KtdFxh0FKsjkifT3
Ckt6rZfj3ohh+jhAY2kyEBe6k7rcldhHUVSljG3qCdDOwgoJjSwpSNRaW81/WrdT
Tn1ZuqJn+l5jf95Es6QgygGj0cHc2qL10xRyuSfckW5SsgXYz+7rfjqd8FVj5k69
I7nSC7mrfwyISp2HqsUmRbJemu92WNJVHERS0G7WqK+WRXlmWfBvHJe4d0yb1jD+
vU57POlPCXAeSXLcPKCwt7jh/8ByMlQMXuU3+PeXFDXBtZ5sjPjxnT5n/W9xjF6m
qMxsan+SZrTJjL5V8GAXFaDdvdxbNmgD5I6zhwQmA0RIhG9iVh9VIpJUvz9SfUh2
F8LLYHOn3WRtkvgck7XG7/oJr+VAs2tmPMrTa2AbsnI+LybBKWQa5AUOyeoswM2w
eEg+Ovdx7JaimBXNIOfjsVkftWGhdZQ7gl7WcUhTIRzhl0vE13Iz9SOwAIYVjVvu
jOYSmsh/5+aB+dKJJ5CUOELC7mud/lMtifI1XM1pamZWr5OjEnCNKNQU9D3akRXJ
pVAiDaOxx4MTVz3fl9hOe29SRE1xtEVa3LhjOLPn3ds3fP9f1AmXfuy4cbyQznGW
zpGZ9zKx2cZB8TnjVpIXvTJzxjzO4sMQJO8AL8WB+3yPjSwXCC7KzKbydm6hwW3v
C6JitE87u+QuBA5DoHXFE/nhRfiDEc40e+2gF/rtYKaDdQXYbZpBmbL4F2gAE1vz
TB1MRjVU5KI60M7kRFBmTD7HljwtYYSsEheQdx6YQeX77/Twd73PJYopc93iIZJu
o+WkOcjrNP1ANYEEcbxRtjGWz889A0GvtTiYnwNsuYtZSihs3tYMJI9ZcA5j3xHl
NpQvYImlzJBF5MICmwTRtBXBcNkDf1aqx/7k3X+dEiq11PMdMWksjAEskBJtrwMj
MT1SFv96SyNJ9es23s8tfiA6NADYUBjbgJQio/7XKa1d5ZUR8SK+2zYKWJ3XJ0IM
088DOacpRUyeCP/zkrLu0BeOw+3Z6fRPIZZV2OueGA/QsyAeQvh5DYkSvHjofu3s
i3ZcTkdtCjaqwST92qWceJp7Yuftcq4Vp5TeFLk4b96r2ihVEZVByPBie1v3eY4K
urrt3q87iwLKvCoroSRyePt8L7X2icSK+ZGwqP4x0Drx/pC7Wr56EK+3PDF48mw2
yqIGqDn175jnWWlyFL2DamIDD/KE8RFCsb4nWS46QIzV/9duqD0NwSUF6a5E8mIw
jIkyGtOSg4GANeEvjB3lt7yGUVsZKDXtyTaDshYlCHkUIR/B7qkFsEoSp/k3PvS0
xkWtXbJwLISgV1p3gl8MVbHHpMmRpqVevN9Icq6Pycte82WM+56IDGJTkQJ938b0
IoEy2Rd/0+Bwn6INXZmIrXWiobc2bj2WAsOy6DznL6PGsyTPu+kKKXE5b8cwJRIU
qJWzIxURxveSW4Nddxszw+JOs+u3rHw93tmSwgkTC5//uNav4oztxZ9pz7L6JVXg
G6yLSq7qjKfSbM9DF05cYpUMe7Nlxpx9rLaec61si+RYeT34ULZHqtENSRO/PK3p
2ctC7IL4w0RC/bfPWHzSxVlUVTCOXA/hJJUNZ10NlNoVaI4JdDfNxun9yNlXzDuP
fk/Eg67GMgG8k9g+kg+BUO4QP/nj+XvimgjWMjXQtETMwNuMu+qQGWfGIw1Jy45q
UFWzcZRXJ0ecgl/0yfLRl1wUmLg0NdZVtwDn77E41rg+eB6HRDENFnC7Biwr3KYA
MpTXu2M9xV1gMRMqrbUJPV+mD3wAwIk7I1NUgRGpMyOXLTK6KLJxUzMaZmsIsTGL
2rhHr14vWF8JCGXH9X5BIY7IsHnBEYhk8GJyV4pjkNS0rzDTHi/qUODH6BQN9nQ6
SiitsXRaM9dhzdYdjwwKIkphDjV8yR7B4VKii8HM8pD8UPGr/0HimJMFnhvxSLZY
ZMBBZKKx8znpMjNCavtlRjYgxofbTYgnOlIA2ln84/7hKWKrMJOrSO6avi4JeTiI
VQBh7hwOuokJs0ef/AlhhbT/Yb97Q19ZJlOJTa+VotfigvQ9e+VtiD7mNmHQ2FBC
3gVywDyYmPx1XaCT5cM74HLTiCdqAg4Ti2ep6go1TmPSv0Q6qxS+ZAqpFFBow7rG
rGHw/kTEreEumI6gpCKvd/cJDj8qBIi9C5H0Srs8vzgoPSuN4GQDwcGieZbe/E/x
177UZI4ARMr9BzjUeYkJgo0/qDwZQPq3WPKg8R6WGRxJ3arjzkzQdMIJyuTshpbF
ygX0e1ZRbtcrb3nP8QS5AWtJxmlHCuukzskXtDNPvz3tlHCAv2ZPjcVsXBf7/EU6
IErIqkG4pHWUC066lxFbJNWExr57nYP4Q2fp4zXfXcsAdnsKjq8RLiqWPJzOu7VX
cjtZPoyckt9CA+Sppz4oGIzpAEjD098aqfP6GVRmPlq3ED3e2PfC8mgq0oJ55FhS
sN0rmFX3gFz1/g19gfW+1/s1/Gpnn358vcjWqvv5appW1kwsEwu93G5WfWQI86Da
MAXmpTjKYxrt4ffBvc4USHgVhs8n1NijfRXKfdNrC7O78Z0uEQVnz2ZdAFFQ5PR9
O+zizMzrqPTuov+4kwgc/Ni250nmWeHd5ngJxnuSPEeoB/vIpkeNcskaXCh8uCQA
sinvqCTHjmBYUrxAT8gAbfM9j+NSVzThA1qCXj0hVaRNaCwjH77AxnM97jHxHPt7
DbG07a1GxR1DV7oIE4K5xw6JR8677vq4kkcYb1WeD6/ecQw26kAWUkTnRXDbrnqx
pom/OXs4IgQY/auqk/h8vtI+zLH5EBRFYrOXvWPRyBgjU4IRSIzcWlDQVfDJkE6W
KQW4NNZ+ZCKdePNY1c6trAwwO6ioPgkAHAJY3jaY9UjWfpq2syaJ0ynP/5Giv48G
Y+JTaJpvC2pm7FZBYPsFuHRIWvQ1ksKafBvau1HxwLBZ2xM7JhxsVshgwLVXX+iz
/n5AegamL8f3781GXiw4QnunN9OOicR8KMB+CS5IIAlGFdwXVYpreiDaLywjbFE8
1HSSUzRp9ZmPTHkI4NrYDSVBeSZoAN2p3Olq4OIrGHPRiFMpcgn0g5f2AlmSPxUT
XmL+r52+8k3wc5GOyADi0Fo9Um5KSgZexhw2aHB7eyGYN5bsnQz1XloAlmu9s6FH
Xwechwf5MJYIn0HW8jyYhwP1KgAvhw3cqxVycFYS8sOzK/u/NcPGjQxF6tzJnjTN
Xi6YMgyG5E+p5ku3qgwNylJfoaz5yWVF2/Jd2aoGOAUiL2ofnzDP63tGkTyEDc0C
gkMAZQP034/UxiwjKZzhTPdNgx7NTt67kIQ+SZCeD6zcyhP+7XoReiT5DYIHl1ZP
xSwczrNUGgm+ZW0hfiZ5pvVgXUpsNwWpi0H8y1oyFekwq7ESST4NI4/2NqUyTuMY
twyhCqnOXz8+rFVQdlQcJx6ywhgLn43q1/0jmEWfkv8AKPWQyp22yqjv5JaU0koQ
BY0q1uR9nswbJCmsaaH7A+dcx+ctfyw2kfif7j9jGwgGNdgRQvLqwc/F4i5660TA
ejgqlXo2Sg7FYysgRLOD+Hc9NRGYeWa3TmY+JmI1t1t3AstVIEbiCTlCETOn98wi
q2sT6Fr0fXQ0rPbps5L7iBdgm/P28hRTPw22TSRIpTLeILmD9Km80nmXJPIBu6Ec
pVOcG0EOgAYxSH+HNbUuUcpnb140GYCAlVlC/5hER9ixMUzNs4lF/iZznbmFQLd2
hoa9X/d3xgpAPZDu0b7VYC4Ib1yXsxF/liamzhwvh1sOHRxUHCJhItCQzbGXZ/Tf
nVfyHp30Oa99VVM1IVCCbVImF4fVXSUQ8fWy/T1gIY1HeiSKwnX92lTGyQJkyWWL
OHAAnjJNpp+7XtWkyPAYINYD6JA0Eu58wWs5bQRMLHuz4l7LDd6ihSZS1BfE9vLe
PFmA6uRAXDP0fkdT1Lr3B/Moz/L0EEqD4joEbAe5DLhwbd0MheHhIobc9dhfyiC/
tG8TCOBLQvHy84UxU2DKxe359N48My+JyiSYwZpmAHZe8i3j5vTAUqWsuYQWsjAm
agTAd+EZUCjQCUoG1bZ1FlX6KRzvi0M/KEJsKik7H+6WXTD1nqE4wbiSpI2RiVtI
/KlhgIBGP0lUFZf4glk/+0ml3YMhXXdnznyH6uKKL0OTPKPWms/4Ay1j48y5WYWC
fpDW+9osJSMnDy8ELSGUe+XmKVQz2wzjRx4ACje5J06vGayWFaYC7n2Tz3u/DxyJ
Af9QcEWtap90v90wPgt6GEoIyVPt0UXaKPT+He3PMKJ2qRGqZL3Rwv8OtEMjYBJt
hrrBHEXyKfkJcHfxgXqGgS6ITo0fdNeuWMgvhKdTtWQavNFuBKf2ljIzQX8BKr4p
IpR7eZtR5k6FBUJ0tAUQyAH/EzEwSy6ircwPYvZNRcdYEVC0Hre9t80n2CZpAK+V
Z0eOibp6koovUPYlxAZ3g2WsixSRvotL4MfPtfYkl97I6eg4LEDrlkgwgfyUijjq
bK4sybB+Li2vXwgc+4E+ZL3ib/3DR4PloCGm+HrC0BNYWTT6YeXsS+JKQ4bI/NqG
IDlSzJlWzoIPOH4bDXPXmxF1C9cPu343UXiHzIu9bePUVufYnmlUzJh1V9+jwfrx
7KUlUVMjSvKCiFPhA1pgTWHuA8HHxyT84iWjyDfk1aJLnvwh+aCYn5rLacksBobK
sGnFLd87qbbY2ZHXJnOp4W3HU+T7EDsTxuQ5sKKjuU/z4C3SVpg5igw9qEulF/JF
mqkAa/qGtSc+/nC+pkIlc+Dy9030mFLPCtuQSldD7eORxXzetWiS6pvpWL7MBTZy
UNGFCfqKW2otHN2fyUylbK8mWAkTKACJB3QpPAC2HIlSlP1JPvWyCsoNEHWSUwpY
rn9oPupPu+hgbGPiz/gsYXGJS2D2FKCkEly+xHfftZzd1XX2Z1g620tC14zHQ6jL
vRpzSR99YWiT5bRDOyZKR8Zu7BLF3rrfr9i2Sh0YYBgWXUSoRNKbLgNu92UD6Sc9
MScN8uAqofYof0dyfLokPxHFtL7Egwg6OfvayP75O4IcdavT52LGlp7xQBAg4EZ3
FJjZRY6MNu2SzC9SC/fYKtaXtumgwNGjL/LoRaIPBF6x4CxvK3R7aR/fBzNszfAF
IzpOvXWjzpjn0J92HeJZe85snqxvJishthRP+0sxyoi/zPHXL4otblqtrqaDmAaZ
W3Bl/G80WaTz6rcikPu118RYzHzEfzYmsy1DngJGC407rf6XQTC28so+4rTqkGBA
J/GTD8XF0rC8FIfU8ZAQdNcW9rgod9sD8PgaMX/sc1g7NRaL1all3EfB4DED+e5v
CT5UBRXPV+lrApiO0lulFY8Tz8z7Dqe3Ll/S+d1mQRjfF/Pkz5dI180b7zav0snk
dopzzfHHy5Gt5SVDBEeAKpNQt+EBry/FQGxyqioyW8i6LKu0tTDWI7H1inrQA5DC
1Jv9AFv/9OAyJtiOTUKFPUJi0ZKiANccYlTBDrCmakKaZHaHlZBGB4yExwF/x5ug
zHDeju/qm042uQxvac5XOOcNbPMTPg+dk3YRN3amkRpMx1AkUPlbRPQ7Hf6GMula
DaRGS9dZJGH0BRkU8l2hjx2h/dbJUohgnL75vH6E4fD7W6dKtsBWmd0Z5ttuuZCM
UYbLtRqcJ+qFFD8LayCEUChpbqm575nXhcXYVD1QG+3CD2GlKRNM9CUox0pnH5sy
qgopzuOQpQJSkuMnBpIP4GfJAVKmB6uDc8ZzYoLG8u2yqDYmAF5qr1Xdpe1fkw1O
w38xAk6hsCnfJjxzlSqF9bm3p84WxWHZBOI5mNPYwpPkIDfcDpd/X7Vw40Y+YQOj
NaHyIVP6PXet9H+sPUqza3ncUQSxZwjZYsZbEE9mMnYx2LoofqEKbdy/3+Ykq8go
RUufcb9y5DJpvZijYDXbtShocpiVXjSKNQ0bapZRmDKIz0NT8DDAoNVvfSFLPKbX
mXf7GNcjhaMmohqU8HyndqEMsVNrDxBeO2vfmKZvkIt0sNl5074gNAb2ztb2OEiz
jxYBKTjNkRVFYqPHRpgAtXPR9RWZNJAj66RQWVPBqnLOKhSWR6RiwDjLViB+mo/d
0eih0aDImwTemTBXC0KJNGvD+QCJRUCbplsk5IjG4CEHg8+BDPjPWavksSxeCGf4
/Ix6XMTeRhSsi7VYmo3liCvZ23OxgGh+RgXOp8kvLfpi79+LYa5h11dRbkIS6nHC
sE8CrGTv3WI+uTcRblLMSJqxjj0hN3ykiSUi9pMZa0j2xMRVPFoLW1FplC3i4nQg
QFgF6izaDg+m/hBQKP448GC5JgJTbhUHQttyoJ2jGmWxjLDTH/Cckf81dQBJt5eh
FogpcfHsyZTHBDTSvTyw4zGMGwKcXAfHQkufF8UIFCS09xICBSr/fVZ4RIq+o7+P
xb7Zb/fvzGo+W/Dh7ew96N/3K+50IC67meN/yAsVyqzjJs0pewa42igyLuIRHfbG
n4cFSiPv/7lFgpbXn/H9aLv7EpjeChFF8fnM1o+ngARAGqbl/NRNGHjq+bVgE2oI
I7Px9sTk/tzGw7VJOLzdLiehCc0But2p2vQ16pxh84BVM0wqG8wImxS+XYWTe0kn
bch/NADV7YLVBZZU9kRetp2rl7QgQbnQGDrXkmj9NG/9qXyaKtZZpi38ieMGDlBA
ekgAS5B3flzlJMLoD0BXSXNUhurVfEMF/jIRKRsQA7bOj5RkYdl6hbKuVNeEoE/6
iR7ZmPprfc1zlMlC1IO4mVRqQkRHy5/ydvfWih2TBxc0qc8M4kuLxkO1660zCBCJ
/BoyCXkdisHibTI2Uejv/XsVtvwWL9CxN9UahOjygEZbOwCJF7x4IMNYJNRrSE8Z
K3LWoWwyLCPeeXffP2zTKw9/oNCk7QcYf2T8sadR20aR1dcXuaoj85hazIxuwUXp
cS8R3ssiZ+4VqmSd8xymer1lknOH4YHaCRC4dN2K26FEP0OXgPPxtXdLvDwywZlv
CLC5TNC7XPeXW2Ek2gxFrsxmDY6YkiAk5vFdewQSTcx5I6Qv8E1hvm8RS7dfLphk
H1+vIQzF2uQjluJFEQMQVGnj2f1h0rdze0P9XuQSyI4U3oy5+GCP9Lz3LPMgYlf3
muFw+c7M1gD65NeO3he+4bpq1g/kXgnHK5kakozzhhPoekIOzQ8UJfWnnxAd9H6s
ND5mWxGQJBtP9SZj9EzFW+Xf0SvNqduEfOEV7WEGFDAAyM8Caaw0PHaxvbPXwIb9
xg6CJ5R5dgkw+3vUZS80Bn8k62ej6ZcuNZsQcY6e8feGqCAbVtenMI3uh3b/XCpl
lqVtoBZWsh5y1shzgqX45mIOC/X9ETjZRWMeskv5BJX2y2OobM3sJgJ+6Ix6xq5X
yfp839b0ZugvsGD4VAvq67uBeVrcsj++YV5FK4tXLprqFjyC6rd/PkKgKNqORPG7
ts2VpcU1OK63Od+H7yeev/ahp1yrTaUZGGlt2B0I2XN4MKMhJwMSWNqxMVxkbe6R
AZdoCmQ8MEXrR1NaZDBbRIvi82A3e4iUSPEhemoBB6a/3EzWoS/ahQSRe1Uo7bb8
tpVO19KbNZdtklwDb4+wDUb1oJMMlabwko2C+YhbAyQTXaBGLcwBQEKAzU5MlAKC
2YzxzURLS2sDg+xlt1zU+aXfg06VRS6UK00w78XVXVjYMTTHnDxYU+9ANbXhjcCv
ubhe+WCMl6sCow2X73WfJcacivOOEdbnMlF+/ZFTMuJcQqm9m+ZDZALpF7tj5fWr
x09lqHXko7etCTCGhOBzcXkzqJ3vbfNXGRL9dirxPbNCra3HZiIKE/eHkSepud81
Ljio3QOggg040mwE5EuUjzbXwLsDLDGJCCEyXzjfLJd87Mv6F1KvQ5cZsAKPRFE2
snx1DhknNYNWIioL5o2F1TPJq+qtybJNd8DDUcJ0qhZo9BYvIJUhAjb+qnoqbkvE
cGJoFPOy2deEClteP5JMemRNCR7icX2PHNqaVA4feUEGytYprAJb87lpsXr2SfNi
PzUzuqdqWztldwwkhvUQUCjpF9ckCw2zqTckhuSAAdQt1WKh+7ljSm5FhZqWVgVB
1jxxvAtCQgKGuP2DXC0Z2To4sZbdmFb+2Hvm8WWqtxFt44qQMymRCBYdWWr5FGnf
NIPuvO8b4KBUxHfnD3YpqAPSuf188x8h/bWozbiVaY4JjmVWVp4rnldpt/Hf3qI/
hI+w3gZDx0BgoT/dY+lb2HnaY6tLOqnwvBTJj/0Txq8Go+gU7I/LZDP2t0Mhedhg
4C021bGkdce8+mzrOW9b28r63DK34dH4+yDlNGBhwBHeF5Tb0rw5PE6oxx1Yi00E
xcP7jAhEcnHsiUUW4AnbUUSh6RSqWyJqiUC8py6EU7PwcmlyKgfVNtOl6E6vw1wf
8QSfrIGe47ytji1+DYJy21OPgpKbagT31vpblIXTGB+Dft8QAWMYLlqj20N30pKM
9huwzJ0YZBnxh+IxuDEa4BcNCO9id8JZDd5fMZZjEPEPenoGUiYWJF6KJCNImvLv
qnu1Y0aMBt640j561k3HvksUxZM8m1WQhdVSCwYAGNH+gn09wRNIp0ZGeBX7miEx
vexyIdJwf0MZrNO8CXdkl6vXwTTYzPmcapRX3dBg2VF1NHy/L1UiTI2Ar+Rx3Pi0
ZS++3+tbZytJyChdbKdwkA5jEzoMVmWFIShCMV2zwd8KG17irCNX7rHpjaH4Xlsj
3tyne0w1EQhdZu4NT0J3SlLqZaZi9BL4c2qvQTTWJ0oXLiCdK9ohvKfrkL1Xb5Uk
QhlC2ALAaCk1e/VqrVZRt6ud/rnuyDKelosIyyETazTZglzNYf+EEi/PGz+EkJNn
8jW5WHI2cf4CrEb7iQQ6MKwrkF9k9g5XuV3l26z8NnPJ2uj7UiV9ykxLk2viMEbo
YutyFdLUDon3HhZgNSqut8m/kgcHgXz8OXYKQQxLlNpym1b9igFcgTrZWqbRaUrB
ToWU+PYtxZT34tJUwYzxkSXNMSUDU4amdYHU0IDaSNzBIlTPiFiQGb4pwZgS+nm7
zlhrekGfnp+tFEfOCeE+nTIrqt243L1X5/J9TNaww4doosQzLXZtJsYM5Ivk6bn8
IZiqP1QxXZ1/GX2sbVGD5qGdxzUH9Z+eHlegWSUZoVUknhc+6TlHQDe4KWTZOM6n
O7vHxnY/360dcIjF92H2s3NGGJ8MLdvN08i5FgvcI+TxZx5elMwVPHvo2ZdkNuu0
CcMD4IJOIA90QGhPNCM1Il66CtgtwPonoRACf0LQB0x7TxQIzjwovR2tQxXlVqJC
X2QSFJ+zwPjlOI1w7hU4v+wyYPteJnE/hQgEcZgwfrzBKOgMLD/n9qUm9xhC1RHV
13ZNHfncYd3pr3/Rwcmm/CjIhN1U01NF3GNjgRTNHviU7JGoH9F7MRFaGXqezn/F
bxT2DXz3qEkEhlyZ/2pU2ueyfJAshNtry7tLprFJT7aF93Oq+IMVLxpXA+fvmJYd
xnet53uX/JmUwRRR5APjxqYC+0TpGGC0ntsdwEiDZp67TPOPAk8YQw5PuUkLm7FX
DtDpV9WsevhULo3j8c353K1jaQYQxP102nev3/ZtGNJ14huGF6mq21VLdmm0BehP
J8LyNi8JcJ0oLNGY7NGZmA5XMnKFD1/buu/AG+/rcHUjpOVd7OqvRqkuJEyJPdo3
v9cRNgLnRRJkCEbYoOlfMw1vUAdpV9wYFA4QBTIw/JRqf8EVit/9wLiWuGqW3+Y1
e8O0V1xyYhOLS0WIsTHhR2FtEgOBTFdEmd271tgrdQHs4YRKiztCePjhODvBq4aq
F3T23MR906gf0y1tes1jKtprxB+a2R4lk2iF+yLnHJEbjvusFKgrX3iQWbWZTflp
AtR4zLuX2e2XQ+neyhAOQMIWekVTBgV9JSahH9X7h39TvzxmWwpVng+XHyS1YFA8
qIk7KOHo/Xax2viy8FbBQ9EMzj+jMdmrRy35T2A+JWCEbiMU+41jkcFMF7UWwQ23
R9OYolNGBiluz2vNvW1Cw8hm/NYkZ6B/Q2Th1+gA12wMJylbHw5mI1w3EiGU0yAd
iUl6MHcUlecNkf2P0lvtQfubHOLxlaYdflYty+uF2vGkSG3da9uz8al2g7lN6YT2
D6XZnLwk0x8u8cJ3iIikFbJi52udyTjqJKpananpKmgobp8TP+PiQmse3N3OSVfQ
xu6PTkcU/wefgqVujIqKkeSH0ixSYsZK5IFI0rXd327tVWo1pqaG41bqGPuMpLQx
1PxL7h12RroCgw3tTcyUlFfkQnJulimG+G6timu9Zir6Gtcazyuqy+lTEepX872A
Cl/wAbxsMhE4KvNS1a9az0LZUY63RAJKWi8/q3pcgrZ2wRDhM32j1zfs5PFW+sEr
B4KWjPZgaeCwGXGHmyKSXBGA991d8OY3Xeaf1MsqSPcMp8VX7T2KU0rp5ezEZKMV
C/PsP8rOIeNJ93U+Ti6jRWoHS6Ks86h0xXO8qEqkOY2MVbb918cw4U+k0WmUbcc8
k3ev9EGIB0LId06tzh6IZmBwWLODLoPeIakO+Gps76GcJ9SDb+REbRNrhiZ+71eh
2nCzImelz+k0DjZjYzBN3HzEXV3joysXXBQ8kuDXPuP3/AZ/nz542Pmy0yXTFBHd
4djJgJ0u1YoGcyT7AWMK+QyHWBABDphs6AUedpmGpR+XkVyLAAExlkkrh39LdU+t
BKx+NMhL2im0mBx/BNxwJThoL8GWX4Yf45sPCCoHZgxMmgS5Zq4l+HQ6t/BRl6Xj
ZMK0PlIrMrhdoBIEByxr1ILSMasRBH++hECyKcdw18w5GVR4mmYcm4mwQCgRVwey
tU1wj844UfW3yiCapQW9q8BMYJ9WZhw2v5A4WyORN9i2kgx2etOrIC1iiR2UuczI
aPX9/galTkzHj6bEzoEozP0O0r+phdVa4gEz5nzWOAwt7VfFh6ks8HGkcWdw/ceb
Is0VsZD4cl4hE0bjcrYJDgIMyJ02rG3toeK+JpgQv7ub283K5y840PUkH4jsSVFX
Kj0TbX+s+V+t9FqNUuJ5AFnTfDnW4qJPeCKrZyx+6fXjCs73j5bys/5/NWnnH4CM
X8pcbLXGzL4KWUxm+uQBjL33Y5dneo0mVdf6u+SkojZ6l09fGSp/8yVIJ5lWPJuX
zU5cGJdRxJh4MGd40p4Iduk13S1uO0B2qFEDM3XirwxFwy4YdBSsd49jMOauVWFW
SGmRYo7q7uJFH1DjiRGzJfdhcsoThvCoKCi26FkEMEX+IcJae0x5pjwwzjUkT3LD
vEeRb2XKw+nRhRv8OrsPXOQFgBtKX6T0YQY0YV8uYVzps3I3HbehqeoBmml957Le
BoSx8bTOYjQKQivoqXw6SFSXx8Jh4wDp2KGlaWMBYy0OUoV2Q2oVfsYsP85P0cKA
7U1ctC8KktlD0NQiDgNFjUe1pk+U9nVIoqBk2E4J52OV9ZxccUUN5p0e+gljN6Gm
RbhBl9ZROVms6d12td6RyDF24oF8IHuZVaR92UiCyyssCL7qeuloQLqRv1et61fO
XYtGWRdsKhPxEJPIA5A70LwrvyUHCv+HqFueOVn7ShIu4wqt4In31+b0cmyB+O8V
8IP7QfQjXbDXNoUJwZSbOh0ixWtBYCKVFFtSabQu06/NpnAApisfrKOQLqCEVnPq
F3RzDJg/729HCXawvjpaGFhRsmvr/1Q/5T8RScJrf9l1PxZiRga72A7YMtpT02Fi
U0vE0zxtHD+5Qv83yST+oue3sSRJgMcNlOlvVZdaKHfSHjdRsIetgzAn0/uD1bJD
y9D7IMZ0kIrr5JGDbaVR7PW8PYejAAuF+5MdJpNiwCvNTtp8WLLu9ZmdXusS2Mdo
WRzMzd/Zoei3L4iear3vbzwFovw5/KcuxRTjeHBpAZErTLxnZTpHzfSDP3Rmk74H
utWumbk3qUW7tNLlpv2mRW7ykpdeirpp7qT3qHUvMS8AabRAAj1c4RT6WCcqArc5
wK39Usa8sBpNQseECFc7YiFOKyJDqoCIs9L3767m4TPNn7pWqJAuon4p6jAUxUlH
gWYtKS34KL/Ei56/HXTxLOW4nzoIVxuDfWDp16MQgzpt261Am2CJuwlhHhetME+t
X7mpVpA7/ojSZiIrw/1+y30niKWx4tqb//9ttF9la/Z1+rey9hAYAs8bjsGP6Elu
Js3DNTZpHqteknr0SEYDuyqXsj5CDXVhmYtiWHoshjZCDUgl47rm72iw3NIvcEY9
H6UxNkLQH4ZGu1Qkd2b4wf84yT64wNZzVjUpz5+0z5MZLz3RwGBZjl4y/2jP7a+i
VOM4VPO27FMS2qc6uPJIt3KQLGCS0+bgiOY3l8kHP7EDFSsu40Ngg8s7IQe3jUHX
JQfKV7idnVUuMBvJaPe0icDUGOSYd0DwDi9QmJeY8oj+P/dq7Wdl8+N2x2yGsI2V
wW6t8gDtGd/ZMQwLM06G85hAtzC+E9uXK0tHk4litD2Iqen3ZI4D6kCZq3IEnl8v
Lj2YzuRiyFBEeekcB/O1AA8Q3urzlL3vkKNL7XH/fO56Q68L8yW8G8tPDJA6CsCR
oa2EzHrsU5EpkmjK/EBQQwzznYw5h1gy4zvCufuIzteA0eVSm8XqKOYlkkyT+OBs
SxU7PFksvTZr+gxw/V6omx0PYY4apLEsDRcBxfFC0nBDXrCp/PJZEFUHDvZLjC3z
D/KZRBQcxnTXm7Gxbp4AYGYkRHri0Fd8CeiTZCPQ0CPaOCZRlarSqScDl5i2m53o
WdEmNxak/KvkBqO98Y3nULvlghT5G2219q32APBqmWk2miY94d6pIuBTP5Ocw80a
kgkOimTssU8wLED8FiFsdttZPg0XXjzQ2j+1XfGs+k3Z+/lMR2aR6o0jIe+kqv2D
kT/3gnaJvKq8wTMn6J3/1/q+uMqHzJ8l9oCKKj9B7h2D4sAHtSuS7Lwv3CUsg2f1
PcZDlM9QiTdg5TKpoGib3ivxn50ixZTAg9dpNVJhggpW+muFsgO9fS+eDnGNjBo7
FDYh+ismbwlgidRN1Rkh9w+2/JpYlGzRUtioG6YGBXpWJsh68MISy/OTPpfdDKCO
245l/MKT+EGz3eXEK6FNm7Gb25agcNVV27QDQTSxoJSl4e0fgjhKmnIZycvAGfph
teLr/eTIYkflGO+EBERHgNushHjR8JhKzD2HyZiYvFAYqrP9U8IR6sa8lBg2nMae
PYoTaOdGq7Ddzq4Pb9maEeaRqC4+A9qPz+NqvJuetMSb+MJ4E1neTghyD+7QbdHZ
F7WLHMlMOeAC7oVnTv4yP2nmO1KBND04317RbBK2M3+sRDXrPMLth4OGVJdDM5PE
CUXrFx42tTv+9wOS8yThJtwYiL8kMfdAOhL7CTAFxf0NS6uZAs+zDlyuyMIynm2k
BlKw2A+Cg1T+c9HiRVogwLsJ6porBWJA2Tp+dX14+E69KkYA4mRFG9Q+StVKD6Sc
IOwik0U5ziO9qPu3b439nvq64uvJDNpGZwuEelYvVLsNx+ud+FBc+9jSeo3exb5I
zb5YdSVrkM/FuWOrf8d7DaLuPK0R2ZoKV3Bh41U4cN6980rW2cBmpHp8BJ5YFXAT
Tbyr8dvZJ1YXjG6aO5/EFnRc3mtl5K9XP6ZUgn0wVIClmUHqJz0rSuZbeTo+qrAz
+e4VDreLHDPeH9ngdxV9CfV6H8sff8iPBbqus5JfZBymcqJ7W4pOmrexhJRVoquH
LcThFTbnl1nLCrHJrFDIGWBzk50K11O5stUEEX2uz9mP3SKoX2qPyHiJuR2zMBeP
sfW8QELWl451YMamJLx8VmLot41ZkFaUKIaClmMdKOQEq16GYV/HpR1v8evuMqN2
zzW8rc751mqUl/PDdtt5YG8oWwjrxQLIr/TB5yuOQkCMZtKXXTtVOdOCcKqF0ziD
Mk094ncB0nF22P91zua6ZrwVoN8r88SOpNMlbCGF7U/MRVO/4CaOJQVzXY3H7+9v
TWmjLOkWVfFH47RXLXjoxATdfusDNQ/UGeqmWEfJdxgUyZmdb4rHzXfhEHqS/mhf
YNmizEy/6x1laMRopMTCzGZ3avfeIDoSKW3niyeFIPYQAz6fdiCl4FqQN292nwPv
3gfGdXovPSvmnnoGsCDkULJkkHoTJxE1HqxnMeYyGnIZQEYTqstzvlIiizegU/JH
kk5LV+2MjCeOLbOECa3M35kgLwW16roipffDADnZ1KqIbNtKvHo3MHoyUm2m7efo
WlnNhQioVBlPxTGUFILEPh5B1umsKv5T3x5ndKx7ImTx2pV90/0PQh3xF1D6LRqm
XSRs4/fyge44Vltm0BCNxcKVjZgVT7J8MvmY1wRzZ8RtyZw2EDrJRMjkveAJAgJu
W+txokzlIszIDg69wWWH3+klrT2n6kUCB53NukLDneJHb5Z8CBfs8nVshhTOj9nH
HIDeUK6HtkkR2UO8/tSn3tknXrk/7aOwnv5fZLkDBUZZHc3lrsYx/awT9OEYXcz/
VMrzXhbbvBVWaa5uqtGkht/PvsdnUTKTRkH/3951K6aKh2HCIa0cjJ4OBR4Ulncb
1x1yqCSbzWlpGKdK0v1N6pIHT8FHsl1AEvTYkJeZ3cXyTvCy79LR8bVEt5gf8062
QAYD363qyUQS7spHidGWIKrysJoXdqjozcZ8gFNJdGFMpc2BooNNcCR+8N4Dp3u6
ZRAT6k2o5G4XgMlErBTeHP5SUgGZJeJvSQ/OpT279bWq/kpQrniVrEfsdlXi626x
p8v6y2+fx3E+YH6dj3URAjlAl5ad8UFyTjP8Sh9WNWflVCTS4CAkhQn6vlOVbb4W
0FUloA/KximGWJVonui/04/kz53nlV93Emvcw1/lseY1x1kD7T8DPUYBnlG/OYxG
IbYYpuQooYSaK/XAkbRrPiflXCoaFH+ub4WHeYN1V3qRZHRtcEznXy2yEgWozltC
3Vw9jzKBDJnlos9ps6RhGYjtJUb9MiS8VdYw6HFjo97Bdi4oTa27iQL3YJGwihe9
ed5BoQG1yTBqvVNzLtcu0h5bMlp58CT6EMjzLk27nEryUMp9P4Lj2QUgRxFFV9Lq
CTxNGKlNnGgcOcWgllYgSckeVpEXvC0L/AhpYxaBfS2HmFJD3TYUhuy/pY+4f7Cj
MQfChGDuz2eecPHWgsnBrWB+RJHXjRy13/LQjE8+oZ5wjEyBuZhhtZQK0taCB+of
NGNmBYcnF+HMJJaSmi5GImc5IOe761E/BQBLgy2SiXYHLpyxrJrFz5muIQkkaqLV
7J85wRRbhCclgQCFCuMGzVzA9uLQZZTIgTGjCWrqidillCeZLsO9Mv6eWa4T5ItS
TWhAJUqHuX1l1a+WOehmxrC5huQxY0RPitId9qInzAu/PKFpfvRRcusW8xVGF57Y
wzk6yHvrJHhrydJras0om8nDS2ZYkOlKRhbT/WSffT5kiPEIT9r7990TfqbV7Msj
+g0peiW4Pga6VhZfUG1ZTnkcZf18TqYeVY+Zm6NPbZ/Ts1SebBLoSsA7y0Xz5VVL
qFjF+CgKR9P0WXRpdwDvTgWmyjVD8OzICu9j33Hcz2hRGY7G3+IwPtuHnd0FPJLJ
L0V0JjH0EJ/YWHrLE9Dz5irAubLMddUS5q8laWAT6+3Rrs69bpOFVtVnQtjFEE0T
OLQVw5wIZta6Y/G7lXLsiRRjWQ3MAUBEXZl+20QqA0KHL+k+Zky2CgNIuZ5wa8iq
hbHal72Rxf3+aO+xHoV3elR9QecQtCL1awVpgcBEp+ieR8CCqQaismczHUHgEm1V
mDcOVZ20tOMO4XAfSHrYdRB2o/G3UC50aTPT0s6hTOE9EMhq0tqB9aec0gk6xumi
gQxh7tE+zxqH8a/r14NxUDTvXeXZQ4MkD/8prZg4wqgbh5VFEQ1CXP5BbLPqdWU+
TzE4puaJsrcwYp8g8uDzUdDncL2mwLCCTQPUo9Dd+cHr6YSHnA3Q+P0QYGmR+hF5
orZRQuWgH6rkHtbPhf0eEbZ02Kg2PJIHbNP1eTrIrye6ZYLrh1E+l/Quxtwt4tDC
rTWM4ih4ULi/Wa9SKyMTJbFq95PwO4KVWu75ixzKjsYKiJua9B3UPJQi+odqYrFt
bZMj1H60FJsRdTAWhm50BNAiVpn/XG1bM574l2f26CDUQ7iJfvWRuDrbS2mrXGJW
8tdc3c+aTs1CorqurzD2O8cdqwaGM3hmifubmZSD9696XrN2JwnVAtBNGsrFJbwy
EwWoitSHMojdvcCP+mm4RDltF7a+crBBrvdInM1BNgfJMfoyAQfn6yppPh18PWBW
fSFdQEPn3FAap/r6BYWuslkhcmAua6Wgj6SllLl1RREHn3gQMO8FwvrDHO2cNsRL
J7tyqqzVCasGMAmTydqDPeXhw1T89H3KfuV8OW9KV7rD4eKUxBlerVTkbF+lVI0W
3LMKvJk6hW+5IQXrBrNXpv0kG1XM1ozlpJe/O5Eq0kxRyxzhAnrTr4J9wNWuYEmM
LT/UPvn+UX5/lhpJuxk1GrUiqzS1pM3O93rZosLhWFWCWaJgzWS4X0/rdNsEPnel
gyN1c3/n+CSYSHV1/UnPNYkCdeczSzcXuZAQK+nz+i0D6PC6BZL2tBuSi1KXWySa
sjsqyEGVBvApvYVlypFe5XgA9QjYG0m4Hf40zdoCoZ6AdXXS8dp6Dp9kabnNHbwQ
8AxNf3LRQo8EtA/xl9I1OCwWHYSu6Jv7PPSIekauMBDwfXIE1zlbxazAwP4XHyB2
1718hnN//IWeFRqGvp9qtxyks9oohWOzHGclQmnJXgGqw8NqEBAJaPypr4XUcckD
5tYv5wnEHiMhq5hiX7IoewI4FDSt3SSs7cncd9p3zVYrQ6KM+um0rLupVprl6Dr7
B9s54b8oCkOivrb/2fv/72PIYrGNJwrY9/OL32sP8I8u5eOUT5Dj12WgpOWRizdO
HnnXDf5KVout3j/Y1mDza1Nq0UuI+XaG01icSOT3xp7lAGPpnTnNfZ375Wq1jSRA
wxvMJr28NPCUtTTAbDviuhqoxAE9YdscHGLaadKWnJg0vdj3lWCyiXyKibi4BLZs
TyqvRAhsRlGavG7TNW3ZM8IELzH97kXAKgzGoF96+MLJyXGUwEVsQZqLQls6qKO+
Qh4ww66Jppgs6MStRXbQPV97mxTfi78ARyZlbvTdRYSRphTfAjsyTU+vts14QAgK
emvmmqvOkBSs8kb6eYsbGgxpFoScFfOf9e79PMUIHPhAPPFTCFcmoIWy+pkV5QnD
PAWwxBsgd9AjHXtZjJ9hG5whh+bSp0rMhXGRckGokpFqR1URAkyhY/cliQFV6U8M
IVlr056WZxvFfW4UaQIaFSMg5yrQsnKrAlIqi36maFt7fgNibjiLsn4FuG6kNC8S
xTlru/Z+Xn44vDsxqN44YNegAyL7vCYwk/wP/fvT6pg4XK7BO2D51TSzXY6WDxCh
fF8TiMDs+jqA1hHmohoWzh9BRhxt4a4zg+rP/6PrFpTzIq0lIK4l2VOg5EdEelbT
DtOS59pWG4WVQGUBS4XkZ4sdTqerLT8LAePH7yY4CptmeWB3ivbUwO2cTsVPvSCt
ySHkDbFOHUyLS7EKK6hPTq6MGlyhculkx3woVw8T+TYqwlkIqWSOywPV26oy7KSk
CgfuOKnAXuPGo4bNbyp6CYzuVb8HNa7CcbulmtGBHsH6kw9pmV1nMeQ5F5f/FwTS
YtwdlYanw6hflnmYmfzPz+bMaOUg2YTKnAtGvDi6K0sz/XavfkHVnacozB3a+JXT
5OWptxh+MyjQZsHGmzwAQX3zSCloGClg32TcnRbUUsRAEQufB6DGv5FQ1R3wYdZZ
LI+eDHq/eGtaDusB/h6NZuG6nElKh/OMA73U9zlsJty+tyZl4lcX3T7CbNYgvMrq
BlfBQzT4SgjcJqkJUARspCZYGkdkWVPnO1Fe8ONjkyuHPtUVQsIw1ED6z1NmH1TN
mjHpbme273w6EIvx/xCviaHTNJTs8pI8/RlXaJY+SA2Mz8ve6J8LXPXlT9pqrURA
wQwIBvvqqX8MVro2FZahDwV/xOzID2noHKB3ZD+RLWLn/QvqMJWaEwirlji25hW8
cZLIcGmafWx31IJnYBISbpcpqRWRXyqHa8RpNOyQ6v65Tr2jIQMlczhHHq3LYfe3
MWt4vsTE4emQQ1/9RsfTfjNfDdXF/uxbXiJBooor1XGgjNJ+/t58tUVjnncchokc
bjjaeR3HuUh29quUUfE0yuVbqN06Bfe5bB4Zd/IhSOfeiBJzN4vvrUwT0eUSrdOX
6D6Z76Lf1IURO8lBxigAJsknJNJB1Yi7faIxQSWOjvlKXhw1t6XDoqHXvhOvwLmV
5kv5ksxgP/DllOTrZa/IKJtWJ8UOSwsjo1b3tuQlG3sMAPa7X84E1MhYLtBL37ei
TQCTVfRe3LNcBj46uEY7Xdow5JE6YCGHAJ3j/kjZiIe9/ASvR0oWTkp743jOdRcH
OFV1rEK4yC3L8WwCiCwnivEPBQx5ihdQbPJiFDa1/u55a9+Xy0f/uuAlE/DO+rqt
5M4jEUyUQARZqSrpU5kpG/q100h/5M51xyxNg4FuT96SulP8zVhwpBl6RDCqXpeN
9+Fu3aUos/8MzdxxhI5FtZ5vvjibmKQ0U8vIk7eLkEEFY0aQlsqRfIX0qJP4CsZp
/vzQY9UxrVW3Tk7rCJfD5iu/KKkaeQnsbrDLLB3MpEGy20Gos1Z6oxHnduopZKWW
E/sUIAZNsABs3pI9M1Pg0aFqdU1ii/B9HaXx69M97vXTeMjeDEHuIwAgqhcgQMD5
ZTwRRhqfTGuTF7jF8GF9GlvGygmp0L+8A2OOqSYd5OKYVEEKzCsQ6FFzxC6EWKVY
ppAihCzqm3+skTKa++UvVB3cvdNH74+LHMymnYIzCU56YOxQ1Cxkc7ePW3/j39AZ
JpROQoN3aEdNz0gPfDefMrWPhmz0/DvxakgtuTnSa26viQdeiLc/axE85SPrTNGy
ntrkgPIRA1fKo0b11aYnfNg8D9vWpqtu1euGezD76RY6vqbciB+S5ZmdOduZWo/2
0aEalvp5omWz9P+mCjh7FKgm7urd8SqVIsiERfXpePYwbObdOHmaSvAz+jfgPgxy
jsoVjs1773V0JkEaU3TAFdrJuNmu4fZpR8jMV9Qh07rOS5Npq72Z5GVFIpdysBcH
C47ImnnluBTtML+CsWfWCAnC341K/X/bznQ1Gj9ZrUYNOXnRe3gAoXL6tsP8xSbP
vJz7+tWcPusdcjJbRd2aICqHHjx/ZONt4XrQ2ECfLAn2Jfjq7BbU96YFebIwZWHW
HXnrQvE1Aoeg8DqEls0Iih4Q+H+LKC4o+x5c5EKb26NnlKGotRprmUrmJfGAln4M
FtJdJ0L8QyZlBZzPbBtf6+KtvSfMPXupqQVbgQWv9k3U+664qvxgZfSku1rEww9G
0Sqi96v5LS43bBqwrMVLbkOfPQ5uJLwoOZLymXS+XcyPcsJG/naoCcmmUcJ+Ukh+
GTb88h5Kb3DK8QCUe4SGB8pKYnPAstKt08M6LEwwivS/q9peWGO1O+b+Ws2Yr7PD
ExX1S0ceQ44jk5UigTrGULGGgN+FVq5QZ3QbyhNZYAzaDQN5EkGFT/Rdz91OcN5X
RKw54merLC024VFUZ3HkctgCSCZk1i3BZCwbGoZYPjY8NgetuDzdt4/sO+PO5zSU
jEjxn6Z3zqIXvQTZUtck0iRXWhGAj45lMEx1c+iuFS2vMF7SYtIFCJ0rPYtCTS6e
WSfETOi4fuQwHdQKR95sW0gMEaXdv+DZnH5/6sR3FXVnJBBb/4H+e9VY0QDVyT66
0v/CzIieMauHB2VgrFsh/qWNAYlBIDywOGmape8yskgs+tsrM38s7cHksyT5xVg3
JgYRCbcwl8d5r/ljHEdNEUMMNA6TE5OX3nKznvRb00y5EGmobk98XWIzVSJHnjQV
T9znSs+reaSfTCk6awv2A88jr2oNAFbzQ+GVa4MXPZxOFDpA1V8GfCzTATFpzfaR
IMVcjoRmGxN3Jjjk1uhr0+PRIzfPCQjOgD/+j2ovC0r4n9ygCVvpgsazWWyuoLgD
ZxXN85+lmAv8aKTgIXQ7ssSqxxuafiwAta2uf7/SwwWZ0rzwZIzUPWteajD3lX6Y
RHHOAi10lBxEXAoLYvV/pbXCxwPwdbnXUSY8Bvtd5nHAZu1JHdZ0b9fAZtZivqnA
B7TaQKfNHvXX34omWPc5GXwnES17efXzGxKuHJJQK7hBtNuINN/kX068pFVY4Rym
UQpLvuO5MfZSmSWMbOc5sMlfqrIKtV3Rp/6FT3HUBsuRIVJc1cPPbB8KgTToeb/M
hWLTkUjSGmaz9hBUF05gCsQng3Vl0G3tlF/lkNPh8W9PeokOYqlOxEyDziHyeZLa
4tXvIGWqQ4ozG2MNSpP/gKszwu7NxaSX33kbIKsJm5S/PlJy9ntirz2XeWHLTJkV
dU2QA8RItWl2u9twskkLYIVPLnGgWk81qN5a6MIKNr8aCpgj2i8lZzdBvQI8XaVK
DyRhxy4bSlghvUByenHtB3pMZvTKoaL9Bory2lAtfjpZWJsu+3zxIxiZjMPNjxeF
3S/+uU54gTXKf73OpY2CP85NBuQkiFJlleReDjxErfWTGEx6gOwW+2W60kYVzc+Y
aYxPSrHQWmn51WyFsx3KCpGAWndxBQ4gEZwPwIc+SlHOxrpI2Ytn4fkuepIIl/gS
lI47daBapYLz++0Fq+QrpCBeH5ubvWxBf6fejionJ8Ul1Fayp3s8sWNWP7jFY1Ss
Zi89dFS0EEFfXZ7mnXxoSangg+xzuE1EWSmjidS1mdPjCWp0uquffec3094wx/DX
IAOxGlGW1VMHC2hKW8dhoLd/G3zkmml/XEH2PVkax2TtHdo6l+8i4+zcc0AtSub4
WBRKlwwQGeyUQKE+9Yl7GsaPlxtNVZ+OAV9eQJJRFfA9mH/5Z37v38g5i8ezwdN/
hdymVYYjP/aEYi47iKXOrjxwa2QLp2DM4lLg9FYY6oVSkdY3+pgT1+yL15cBk306
ErM/LdZo/zSpjAq7iTfgiWRWZJBH+JayrV8du/KVOm2avfazpe3JUpkG7LSK8gXP
JZKbrVjJWcX/btVUAuyvH4xQ+FqL/udNI2W32XpnqgnO+to48K4rMkj3kaAmPMCr
nE9jOBjET/W3HUlqsho8oibrdzJxJU6x0Bp/BOOlmywuMgeIFtlKTNWMsMlYS53Q
//onbZfZdpe5bKL/Jlsx3s/jc9p5PAR7lTrF+SDhHMzZ6gO+1J2WrdczMhTRny46
sj80bjnQ30ZD0T7I+x4uN03GQgPB08BZZLjVwe/Xbg+yjctiiRjBLsMopoRROa4q
oiylL1nl//3iEi7Gkub/fXkNLGWlCFWOeuxSZy8dZZ06cgC9gsOs7HwF7oq+RVom
mi1FP98K8cl41CCrlFhUVtAe2rquomyPscujAeYp24AnIo1ctEdD8W+4hcXIONz3
Zs0PzXyu/D3KZ5JRMGM8xUmL4aE4bUOuT3p4qrAlao8c3RYYiyy5TrFwvAsALLhK
At41KgxZ5HjbiEqNJo4o090/guW5kEtyyNXjsHnn7dSsIBbJ3O1lRkSVFdFdgptp
ZWzVTiC7tWbzcZQ4Fy1GYe5Fog26TZIzLOH1TErrnAus8IUskFDtPR+pI0wGqJA2
FLPr4DoT/GptQcz91YeS3onnngcjAx2lPNpfMmpRgVQSf85fQYGcRXL86FqpMwN2
f7kwLHsbHknrm9FcUtMsRCFRNjzrlXI9Qb8OCt47/LxPbPmWkyNrrAQ3rfblayls
7j7ywYHug29xwcmtbFRsTHc+0GOCvoemMmy228YOjGaEFMCzax3UplyUOluO2I+Q
lv0I4QtcldP2gHMJPAIyXLs+2GSMT/l0cVD0Y1pkhX30wrdPLywgtHe+43Oqa23S
x9OgrFrlZjB7I0mAhotWwvhTChzcXwnMOCsGYeSIjFSX7A6bM4Lp5emxo+6vCzoH
KgmxizK7vcc+fvlV6hrkkh1sHJbQq8kppVVClYnv23Znj3utMqv52QBBuLKS2vAO
CbUHVsNA0cB+aop9yku0l2irt9mNPERiU+ZhJVXOINgJXBaAw7DvrMYOO/t2ZDi2
Z5+Ic5O3AKQPixB0SbXAAjceHTcvamF4zGyrjFtzndwr4eIHB26C2ZS/u9/0KVUE
U1xWJkGd+brcYH+7Zy6qoruiO5G7SYatrMhDN7CSBSSom4+k/fXuLq9y7gVN6vR0
IDZr6d+nPTge28y+HgH3bt3Xb3z2F5qFcSNNy+FMoKfrdOCi+H2nU7NbSvZVLvYK
Bk3PPLMsxjmbLpu2FQOgIGdiN0ykXAYM3QbWv5bDFzrSUvtGEL6gEqJZYn1pbjdu
wTOUeNnPfeAsXW0JqLqUTE+xeSJLJgckm2k0pGqCBH9qc2GLxbJYg4S6qzw1rw62
FfvHloIhGWhmfCYOEZSgewOQ9koIEwGynk4e/wgKJ0/xjPuALmdj3gO+dIjvdvK+
+XJj3FqdmcVoRmCcxc2Oo5r5paJ4bzbFA2oidV5tcJSAYMS7eql2S1gkju1WcBvY
wotcWEy9/F6czscsYvzEvFdj4QRExl1FL/1BiKE6cP5iqaLVumbwBmcbhbEkaHHD
o4Ehg61L0bHuIGSEGnSyI5HA3r4lLjT85TQEDkKIpcujCasB4iE6Lg7LqocQyM6j
WQIPhEiQ0lj2SAkHWpqAuElfnhfCCG7yLQ+z8zFo+uEZ4wHL58LgzjnZuRQ2kSLG
hF6HPjGDlbtkqFWzjLVx7VZ/ZSU3W6DWl4OFG+sdoxtGJdicnD3STdTC6tKQSRDU
VmFfvFWUzdLdjG4ebquBntP4XO2szwJBUS5ilPJC9QbpkK89khvicsu5xiWr6R09
4JfVqV8c9yYx1fyduei7oOgbpQPjMgMb3cjhubh+uBpZWiYZ1jjvkD7C/rD8CmvK
YLWe3But9KNPa5JKJGbeM74ZhlggdMmh1Nm4408SbH6GgT/aDNqSPFQRehA2IRAH
2/xmG1s5H2xGo0lgs/G/HYwZWOZd5GtPhR7n7siSLRBVPSX/I7YG9WIuGNCB+vJ4
WeCKuYMQRYG6Ys6MkNY1nUg3rFaN4ikO3RX91iIhrAEwzmDD+r2OCSwzrHjmhesB
GXE/DnlXS02ZIE96tA7tgHNzHowbM6spVn8UE2Q+jV7SObFXUJ1O+QKfH8oWWV49
YUkYpPP5y0GS3Qp1dQ+EQb80wUczGgH0w3JkwWWk9RCq7xfxJK8z9G+8W9GcxRIl
/kNY0sDN0NuVGnnkScEYRBKFjZQsQDVrtr4xxryjj5yx7YXleqTW1xY5DEWln/Pu
Nfndg1m2XL+IFu6wJZ3tEM0RxbZNbPVSspuvWYKJ3S9IbovEyYz/Hbeq5nK4C1Ml
1c7VTN/DOP1iI2fB9KNTgTYQ0yZaz/S3b8VXHUvzcfuJFz+nkA3PhXq8oYOT07xt
nNd/6XiCPtPzQYbYK5jEJneivWHeDjToXfako0Zlxw44G6omApZ9u6dHKMEk9A2N
wx4G4o34ZMnNrPH4wibIfge8+2yeZ/SBnpjoGkSZBP13WFQaxH8E9kw5GG9se7nw
1Qh8jrQ8H977TrDhnu8RbTyzuTNz5eHgldCw7VdONJZuUg54GOuuTisxiDEIGfWj
PcqAgUwoEB7Ki3yXF/KToYrZhsxlyW1dwLzWTNl2CaM3xhKfRU2AqlX+rQMAQH7G
d2cH4PFW1SrDGbJWYQDMB8gNhjvyPPEo6A6Opt75VQ2qM9jgUfp6vZmRTs1ZLR2/
vQNw1JYRkY5gOU2Uaswkk+gWDf9/zthCNebLhhuXFn9p1w51qgnxjxxV8qfYolhk
5suyyt/69MRU0703T7tdDkglLClwmdG6ueuWLPnHSLpxd+B+1J9lsm0Y/N6kiIPO
RzMVyHJP/wHh1zs633sZhQjXPrGj9mGXDvY0+TBMHGBh6LidWCL3LljHKll3g2OC
i6rygmXdJCY0BcGs0+f0EB1XP3ZCehCXQyb3cTz02tIU9KXwYFmmySfAUOAKVqL6
0aK8zCCno3lP17XC8c/KYJ4jaSu0bstMRGy39CQxmSNEuC8ecJYTIjZtGy8V5x4y
efR6LStT3g0v+chRsY4H6fDyFsfybvixvOPGC3ThipmHrHIPeOrnM3xY8R8/mnxV
nbrJJlv9CWWPnbsJtG10hJ5oVOY7IyqPKKZu4Pi82iu16WV1Xowfwehf4BVl9pqA
5r3QPdGK0shKb45XQWwV8AsDjbRrr2RgKaWOf92cOTe/8Nfa0llCasUPoAYt9IYk
cSgc10tDSnUVAyxtmYPNpDjogjkRYOOC37jfFiPJXuIqvSKt9QoPQ2YxjkU6H+IQ
fTZJ47iqTb4arJEeA6YSKUcpXNihT0vXKZiJ/tE6QL5UzwR+kGhG0x4WEsxmNLsf
1PuNlFGduH+orqTi21ANDkqf4qbp8+9SOHYp1Y0y/55AsNyw+m83oKKHwpWcLRAq
RWrtxY/EfugdEqfwL4+cE0ytTEicXEz75dI126BsNlRdxvohp1Ncup3Iy9nobAfz
SxCD3fnyGwpkhgwhHh2u9neKgJvYHuzBRMEC3HZODznGyvd2OvnMMesFoy8ZSu6H
bZLjkoWYPAQQLYI2togPlDJa90xTFirjXB9p20i+SJ4UXgz/zwoCBdKYCMpx3siA
h85y6TmodO51blMtXvHbEVyxhYznwiVijC6aoF/4ZW7tOF7SxUrHOZ5oaRBLeqy7
SqhIU4vwO3SFHg7eYoxsW2WazxgDXdwW4RRJbJz80JP+PjOuFg2tAmYjwUmBfzDx
6xGeXHOiPc9bp1w9GHjrc3NVT0HHy6UpdCXyE95t2xSOs5yY8ipdJM9tUUxQ0z5U
CV+EOomYYE8cWXJPm5CX3Mo1oqCkSaPMu7r6oegyhXwiK7jNH/lUKNq9rvgzC2lf
oCDYu3ATfnpZX1xgf1Bwc34kJKmfgpsZV9q/8sdTriHjdyPwPb5f/XXxDnw9Ikgs
RLW8OBZSub1I0SpBi7QNLEENEkljrCFURNMzAahleX+JU+OIXh0ecKNHCJBiIMB+
Ni4JFqvXt4zLYO6yPSaEaycAssOh/P6fLShLs7pNeOmoRyDOPoGjS4bIyroXt34k
9LDccmTOirFdNpwIbVM2uRelNM/e8LkWwKdPkSS9UWohn1r2jSGLl0r3AP3e6BNm
+FF4DfAFj/FXfTZROzjD/qkuW/O7b7B/1bsjbhX8hO3M1Q0Q7GJJsSLq5GeEE7H1
eQKNoP9d7WEEGDQhrwo/MDPiS4c/tQ402eyOtQ3BQ+3XZrI+e07Ra9OgzAY/ShUz
NydiV6eD4jatXv6xu9D7hc1ht0iz9djMlBeOGNDNlnZ+aKinMVJXZ70Iyi7I2BWg
+KRyTQoK9uBs4CWVEVPG8L15o42BOvP2e9EgjN/IItOK+iQyxoViwDoULXuqKzmy
1suqboUITFvgGWInkJULd9rtoBEeoHccWAB+Y6WgwfmOdAioAFSjgU8WyOdtWWom
r8VZ0jGa9vKmw9d9DKzLz2CHHsaPTz1iAGR5VSm7tFQapCP/XkzKDkothkECrH0g
XCwywugoCmNIzEwRJKd9GlPSh5NbTVDTl5gByhtfyqe+7ZPDxZmUlXjOroGeSAM6
mnOIPFa7lAJ/aPRjW0SBCTgcPduXbuahIDL4fy4815548nRuoPHJSMvHPcBbD4c1
ttl4+jAPWQ5MZO9VkucXJ1VEw/+JlbUzhls3ELdIRouHKnwXmyToQa6oNv6XJkNQ
CLWnCpikKIS7IsdbN/evYlxbLGsXcuCsDduqR6OYHrbcv7qL3DlFnuBANdIjvr1C
cnY389t9ASB6oIrLEWl5SjvEC2lM2pXlIE62un4qFvMMzQ7XQiHoxX/yxqNA5blQ
/ONj4AJib9KYkzFQr/yJhW0ZBPUt1qQDfaGxtEK36JywUorvuNy0W0DfhGNqYkTN
HBrMsZTwoU1CbrrlIMqPt6D9WBkeQ3RGmGDbQOQ2K7erFea2zmBEKg1mvZPdFsN4
n3tQbFO1I3J9pIEJDJfyTzgcHTRgc4BxDi6tJLi6MUxmL7ipySkDNrGsLyV/oO9g
owQgjvcXqQQ3OjbhWAg4HJt8+0HO5DLTpY7ti9moF96vCMECPDVLlLGO6xht3Z39
7VYh35qAvlcO3mQIWFlNZPHVKkOmUeWQ0jtgBRGuwmYC0vg6kRvI1qfye8fideNp
YIT0VpPq8h0skdsSzxQOxP2ijYVDH1LgQ1+S+gFK73SIMIkT7ARgGLVBJw1Vpk5i
il/c+sF6j3TsQUarRhelUia9wz0vMekUwhV4cO0svuR/ZLAgU8htGEsC7Zcj50E9
u7vN1TRNBODca8ArXUaJd0HQBTtNJYuOkiC0DYbPc428SNIxzS7/RMEMrnDRUbpz
BRAhVlqs6VNJzQK7CM+hgeD98KFDlVzXiI8A6l76X/3or3Ye4vRmubqarhIakbvq
WfHzfQ+ZrFUv4GLKFYwoA87M7QynaXqWIgB6NnGAlaorAP9Loj74niL2vutlfosV
EmhnZ8GuRWAge52BaBuT/FJes8KwOdxNnYvMLXIUfyqqa916faqhCQQ75ov4u7uK
glQ9nd5ska4KUTiheeYHuFAuyXPXxVBflQwSdWQF3tOAHL5WyxIkZtWit76TPQHJ
LqBtA87zt8o86CRbPqmxTdx31o4mVbyWfhj08TNR4iFfCbzdDDlBOUmsIG1rMtwX
+tRieS+aMWvSNQVpc+VeULFA+ip6w21CXwt1v4thI58cCMYUhyFZqGwhqvzPn/Bm
AlEDJGKid/s5Pt0M8nisxEdmoMEasM6bWyaKv8mfmYmWto2ohfIqzF40ef/TiyfX
K1Ucgcb+8+Omf+gsG+GL8I2p7E6/IqdL8h7Djdgr1sn9WM7uQgj/SdZFSLSJEPl4
WeA/p4ocENWkYhdStrVJQhMiRhS+Z6oApTMYFubeuXfkZIa+GCRJvm+aOu+05L0f
8oT3suHdXVYLSjY6fsH7wexs5kuKgae/zB43qN5BsGKDN3sO6CuvsU0Vt7YQO/Mj
n6GApMXZ8XKEdXzHP9serQ7SpeUTRFkDFsWdH+kc/03t9GCJH75KSwSprdjjWvio
xulvXpAdnLRGtVEms2mYiNKkeIgyogg9ABHx0uwo+FP1M6Rblzbe5gVoBF3SkXlX
vJ4DocnmNVuftC/NRiSOoqb/nGaj1RAqPpy7dl8K9UK1hOoBrDyWDGikoPti3wWx
tWTIYViHwKYnHj9wPuLKgR+ZwBTsrdLFCB2JV7RXG8J14K900bVEcH60O8/WUaX9
cr+Th2HthEQj11GD1lCxylmwo9gzobpSw6BNQkSl5ECgUpACzdAuUhvlvK3RA4aK
34kZnxLx++uFH6uaqKsrjXjWvU4JMR2Rv7t0xfs7I8ma9A3NgcanXiDFzDilbNjL
VHTNuj+1QvNifYtBBT+xq8RsDWATbOeHIegY/hXpt1v76uQq90a5EA0epW8LGHZz
PFiB7+aNHz6DaDEYR0jyEvk/MTBlvMnXXA21R/VoqIm1w1850amYhfj+1/YNsYE1
9zAn+x98KRlV8CU1LrJ0nBIIdSRmX/Ku6Lvo1tpd0xcYAFX0OVopLNz4RsMmisjP
GChR7naf5RHBPwh12gDnmVrcasChKUlALOFtQkg0tO4DQamYGCn/rc1J+RGQv9+S
yugrhK87mdozSkS8YD+vrRqNAB8SyeXQzW8L29GSgnDM2ITSM9nf6BgMjdNWCu6p
h8DTTrRVUvPe4HifpPRbt7yfm9CeMRUMpk9c+x0ZWUg4WkTqzHKRwNmS/bEofy0q
nlxuIrGr+55Mrgc6LICKQLr/OsjwBLiwHqojG5PMLvESrM5xBGOyG4o7/c7dyTYW
BiWvOky1+ejixVWW22Fl2vsoxf9gq0uwPOPzGxJ7kvbHhJ4EwV84NbfkVVBSAjnq
4BWpBf7BkSXM8ImBY4ayPX3v00ShKqVPKkssU+oKoCxxXh77NO/LapKmlSA0OTYO
D8uJc3F13fky7oqS26MQ5REAC0lA8c5IeVbe9JDArHc1o2RVeLs4JLThi7/xsZVl
vLY0vv9WZ9D/zQqo8tkIx7vl9tKyR3mAK9P2+ToiVv+6FjEvWe6kZ56gOzX16ABO
FolmkiDtb+2tc2gtDRTfIsJnGz99ixr/4GvKxh1XrYzsVwF5Q7bICAm9VJruyaK5
BMP6gd1WHshwtfuK738A+U53IsO08TylrMdpPQclWTQVbPDv05ujUUqlyrPfcHBa
Xn3apm3NFtIjGV7j34DM7v4NhTxctVG4hXfoCnNdtx6Z0kHJ1gqb9NYZgR6TueK+
OaP1zXg7sYnyF/eJkJ6rzKR7ztVlTiAT9EpqOr6cbjw5S26SobkOfPK3YydJAxrP
Oc8K1vM4VZyVrV4MCP3zJWvGdvKxGQjOjoWr3/eT+o1rDusxJIYd3/j/6BaIVAlI
4+bidAqMC33jVPWv2ZvbHwUMJ7UUJf3uEP9iauYXJnyCA2GCoPfDAqgs1Sm4mr0K
FhRNsBzgVBthXtgmJ3KzA80JWI3b8MfnGmziW6oAZHT+UnPxu2ZGm8wsWzgD8d8l
jquEGDaN+1/GJbt9zW8InS/dD7dIQ/EjUtrQCxJXpXadnwccmYhVSKeKSFmqfOxL
i/TEggkdmnfTLCp28GAY7CAeETYPU2Qz19zLkxaAnQdRud7UhDaNpRBtMS4EsdC+
qfKx8uAwB143GYd4ChocuXUIG6Lf5GdGiJQjcWnIfmjQtCj+5kRp3kBmK25BDv+k
hQ7rsitmJFjgh7S26exmtdAolohW5fQ/AcSgfmbqrE+WlXbnBMENqxQx3wDctGCz
Lj8ehLSFz+SIWfdBueeeqTMMBYSUK0sV2Eylp+Ecc69LZ1RVFhjnhdBPx1B1N/it
APQvw8QejYtOi8ZaIL4MPDgVVHO/LWJCsT4Uko5fSK6yd/4PZattYZlQtCQ4k06C
02/zN6KdJz1pySOF0a68/09F3n3wG5VTaifqi4khVeZYWHy2WM2WMaUyVU3gmOUY
7SKDZ5SC6LzPQConVjfgUdKla+VYcVDxloJE5W+ethwmgkPkIARWmh94y+jYKDq7
r0/Vz6n7AZGlzjMiI9rO3iskRWIKhf4BgKWMO76GjNoCMmqpSHFZ6L9TGlhAKW8F
hg/57ibygr0DPHfjsGuvgnl4nW+GaD0/b1amkO2GcfHGe3HUu0acp78b80xHQved
604TwsNuQxA41OE5oBrj6eY01d2dsii8NVYwJNRz28gRTwa/qzEXIizXL3bSps3R
kYNVfStHLAxIf4xmNWORg2yVZlFtT0yacJraeWz9vjdBRM216u7NobXuRu3jlCmW
sKnKbhv0FTdD7ecvJIziltLMdRrVnIVqAmV7MXC3x+XyhEpFuNj7NRyZnTU38aqW
VVNCa4unSYtQ1XamV7imMpZlQ8rWExfoia/TTUikwIQrWUJhrvCkQfumTwB77yBf
zB7IXbRNiK1MLztjmYJVGKSX2JdxBFmX20Po9wcEECw/MFLr2LYqCwXEH4KcpkwL
ch2bNF7LVVQuyVHJN9G8B5spEHGZKiMpfOxsRJw7JYxrWVFGmMVprJov6DRBB07d
2SKKyLC5M2bjXm0YzCQAVLiXn8cGBsn7ELsctgtBFb8vcYmBj2pmGwBLBJyLsavd
HVYSi7VUqIE1+/mFpZGjGpoKFbQ7ExO0wd6i12iHzDyeUqRTBD7uR+tFjWLC/QOO
87a2N3ymC2spoQZ6Xl7vQaSnJxzHhrGIumu9xPryWYtAI1yIV2JSYg9k0KuKFv5H
VOBA/HmbCCq2wUwm94vzUgU5Qs/6Cf2xlyrT8VgFS4bWvnbyzhZW5x80EcY2eoH4
CG18HasPhBVxItZdhbV6rwcSPTOVlR4OVQKO13RwELASHxsn2Q+0fK2URzMcjM2o
G/3CWI/HlIjDuqw4x9F4Pvt12c55bRV8RoAC8jwNMurnlI0dbWaCMXOu8m8rNLn2
/91FDddZmwRnNac4bFvanCFLFO7k3ES9Zz9ppmlSXbSC4qwT8RXGG/CZychCYBso
uY8dyULgdUPZU8iy0K4AVX9/SRBYWdrDX9Qtr/W3Uvn7FZTJxbJ/uWdpNs+tkYO4
ipX0YuzASIHhjyg2CjhbkldOi/y9S4SzZJZwYPs4IV4n8Kol/XR/HTuwc9dt1xuM
6MDu0mcfiF31oqrHZGu+QfUqeEMsxPbGaxs+1YQ1disPIzwRps+T60e+RqZ8bh5S
VEuTEHEDlU7n4Nyv3n9pn1dgJKuYCrfCSmAuyXbGZS0Te5SyyVvoObYL16fgTfwZ
mzBuW/BezHTZom1Wel1WjuagKEu/tQ+fEvCctCSZzxKB4t3HdSO0QMMLFDxtOc5j
HuXIExveatwQ6Gm9tgQgo2QaukjrStGHrQbpoRVgGtU5qw7PkyMHs4juq4+7in5N
fDSuPDw7KlHpxyAoHI8UoiAYvT/ucaEg0TcNZNKV3wwpeBzbRcZY3A8NLMF+eEhP
C3rtpm+mbAHp/FyVYThDz3wzt1jlUHB+Sm0KpL7o7cyaQXkqD7/VSG21RWo+Hn1z
rMRiuKSMGsLEhXaeh4LeT0NdS7iO80qPg3/na12Y4rUQZeWRpn0APp29m9Rg+DPG
Y4B1mFmwy2vTg9wO5aF3dEju9PtwgoxxqL8+qM+5yffuC203F3/++RlU9wuWqfJs
2hA+B3JtCYcJu20u7Mqg6axpmLlAiJTqZ4O11t3V/jo4gdNzTqZSMNe3aJzFZG1Q
CLj1/M6M7B8sxh3WvG223Wg5/IueDfWEzeiOhDMSh9AvULAfL54gkaGsW2tm7i+S
l0cI2ka+r/UPGCbYYFBR+gnX4rWNzkFCwCPn5gaD/XG+I7u5/vmnBudOBCLZMJpA
X/GwkTdlM+OeVnwF1BnNsBK5xJA5rdK/hWnM4jV25nzspyZz9Nher8IdAVC2SyrT
OZQlyf6whG1/YoaSPeMOwILbzY9f0blM556VSYbIrTcMq2QEALU9pvUJu17KdyAh
ui1Klwsl+LvcnFljo5VkFzYtOdKnvLLrL1fOfY35vnoQjJjN3WQdO1HBWAEXTZ0V
Vy8iNlWJt+qbaTgvC5gxEfHxL3T62EzWAGQZMevOBZ9MSZwUWA+oY+ciNy6/srEd
mMpEZGqDghSU0keQHj2wo0+RLjZWFi9vP4zWUyTsz6sI1psOmCvK4+fTMR0YcsPA
YVQE4PJSvI+fRmu3LaAz1lzrAlRkp1ZyIt8cAcRx2Tv5kAQ08vHS7iO2k9aklevq
3DwW9eRQNOZUZLk9OV7y15Mf6lPEG7zt54bL9yqiGlEFFYoicFyiylWLk/MUDEF2
DswH7RJRhGCkc+NKxOwont8qUwPLnm7ytpz7tImETX8vx4uGI6s6c0b89l5LSrC4
mywzYUiW9mLkqyEqZbBbJjk+Gp880lD7sxCSCtFYG6omI+FP0caBNAv6EvJbsOXQ
wEkGIrLlsFnxDepvGGpnDAEL0reTB0D6WVFJ9955sIpmH4u59BleQzcEPzvmWM0u
7f11PHFTucWO6o8EQHxnNl/UEPS7YAlhg2osmSDoVxA8rVDTCWHwI5vmAlk0Ul7b
tRHvo8HtoY/aEnn558nZVyuGPNip2KiRcdrChGTOPL1UuIVnvyT+tqPUuOSom2Ms
I75ZuLuYxvz5HAhL1BUcIq9WkuPsdKhISvjyXwKVQJX0GJFXH8RSXhVTz/dXIoan
u1RNby6s1wexCDBLiV/JJDQvAeqcWcRNvjK0RiPrpe1LnAMfCMalofCQFmvwFBMJ
dbLxMcDgKx2rT9BnHn+XzeP8i9t0rLkBUTlFa0vdnM2W2DOgbrdNWwTmHV1+xzQm
pthaji2scYSCRRL5mX02/LSM2tDcnS6lLE4LKzWAEs4kxyCYDw2T597ONizoGAy7
FWPVq6Tzw3uNZBHaLfwNPXco3he+bet00U5vsuCOdNR37+AeOosPcmL0LGN+SgXI
lL4+6zbTiFD9iNDUIN3CMEaCNcoOpUWRvOPboPP4y52VLNc7n+IhYxY6VYUDOELV
E5BA2I3nkOeGcQKkDguSykzZjBr0inFLKUVYZSkXg0c2FQsidMaP7WKyTuc69EOw
K821h0WqnQ4maAt0xKzhVmDB/SoYyDvsorHDLByBKscV48+sVklbEbx+PZu6tgsq
6pfisZxLVy0xXt/f8L5O1/471sgsRmHjunw2y7zDR5w0l09Fijm2Eh8mh6BPX/2r
t2hTgsPH14nq/wwsM9Of6vassqj6KXjOnqBO/LDCw6ySyNbPF7J5CbxJRys3rlAv
3Lm/QAj6dY8PuuRn4RzcKp1qm497GTtBMgPQvdOdmOCgDZxrELIXniK2nXB9Yi26
lTZA/5ALrco3WiQl8RAjqAeeRZqPZuzSyuiXr9P4p6GdILZWZ5aSAp4k10MbLHpO
Co4XJhXzALq4FeH0PGnYnPiCcH6NL8vwTvw++ZGYs/ZapeDwfJ9MBdwW/49w+Lcw
Z9rumQSQ7R0syUPNC6JW6ktkYXq49u7S71gv15VjfOdHFSw3CGRKKzq6JrEiZhw8
+hRi1WDvO1UgZ8tp4JN9zkXwmluIKSQAhYFq0dIwe3IXvrXkX5qGQ5dzXt4Xo/b9
9HwwgFRQTaRy4QS6yOMsMCR0lhpSCLodAfSSeI1m1hNFJB8ihwz5gx0g9mvpBKhf
HIVjtC2o8Utg17bcZjVbdB5bq0q5hsJEhoPoYaWEniKQljBHfWWr/yKWAZYHHgct
7mnICSiUcvCQIEk4JrNcynWjnPSs0KbQ4oKHTDs4HC2svDJTfMKbGgT4LCrM9ji0
Jjj5ijNm/toM35AOKMS/i1nn60i+IRp5ZT5KRCxfiy3674kmI97OpJMcrDSStS0/
42WOLd1j7jGtH9K0CPErzGASWw4S+l4zRZsElYGTwLoBD+psURV7qjFfwhETjzB4
OsrmIl/d69+NlWNUy3Y9tjXyuo0h3MiOTcJ/ledsfKs7cBtlYxvo58PP0k6/PAIh
vDMxv+oHfzugmXp5roIsKGUJklDo/3ffDZKUE3z8MeDnPfbZlm/kArVU+7mm+StU
bezDXW3yAslPWLRfNRiMeKboQiWGOEhgkJN/tGvpn+wkjxIizZM/tGHg4umoK7xP
p1Y4DCcd3axLcccDbsqG8qgeXh79wTWqaeq9GubBYIIiicKIryBrvVitExHyxM3V
LdNTZY95/+UrnywmtlyHlYMU2n0XypQZIKW1/eYhyJ49die4+2VR+ZhSCUDnVzfp
MGV/egoiWjHZxML+RHyv/0ocfIxNoYWFRL91bRG8ilVpkxanvPbBAHhQdKZF0EM+
kepPNFbC4VTrbSMYTUdLg5x30PZAhvtxSLoR8IK7qzEwww/mqdnvw/1N07uay4L0
1DCAjUL3p78Qk6/ji1x98pWx57n/EUIBUFWYQ4qG7GXp5SGXuJgadlBug2JUNVz9
bXbzaiK2xz99kT/VcQGyfH49R3y5fT9N3AVUZud8rGvBJqdSpWpV1/rb/VqiW11L
CBFugkAkF/eXOCUihs+3sbwJ/kCsW6r/al8Sv7GEwuQV7PXG9HUcxgadNyAqgur8
1GqNAadEXMptKNnXPNSs4tpAfIePH6+US1/sU4pTj6jcH6+9dCRkY+tsCwFrfVij
7dUg4OrcddrgnuSl7PO/oVpUWg/J3D8jvvAUVO2o0eHdU3J0ldoiVKvZWoiD43oz
sl3dse1I5FlmEIvBtDkQtS9WV4epvnunHp3cyaf93vv3FSZfuZTQ2UXCVDl58lTl
iLtQm778yPlLRAYB+cvh02eDStXg5W722cZRySWuPNE8LoiXGJlaRuHpoIw/kjnM
W+R6fL5xaLzxIwaCGALYaPkqEMnJ5PEQnmolkPD6sYrJva9ULK55uN3j9BB3SMwE
i5iLOfpDWP/nhnzIuh9j+ylIUr3qoz+ufomQO30UAc4EEaU6yy+mPaqJ8RNmzKE5
o1h/Yf31arMFuGunCUmeczoK1FbpFMBkmmToPLvSU8bY+IWQNid/bLa09jlEDboa
UQ79x3/sredO7YO+4m+bnsILjr+F/QQS8AGUtlgY3teBJFDEAAh6FEK7N+ptfx1D
1KSseYq6ctNO965xz7djXJDVaEBRVB60eh3eRADfJYS72psil5El7Nwrai4R4+p3
6A7fD1C8Xvh/LsdxPAmq57TQgPJ3DKJlUcmM4ojwPRKJVigT++ZUYTziLFscGmyn
ildXseGRJiR2V+vwHzjOo15H50ZQ+8ghAHkjafa47fi6fV1id+aYuKh95DyhxCTF
+S7SBM0PQY2qdoG/Lq2yty+Rxm11i2jv0Z1eBW4zwwHiaLMQuN/02+Jp+QUVI4/f
IbjjNlFWQ3mFdjkAOgk8iRq+P9SrdVl4n0Fv3gQKSpiXFKzVWgED+8fF2izXNoC+
XtMKGB6QUgApkXTsum0QopwBQ09aeEryc0G0/f/S7TxWARAqBccVd4LoG49esf5w
2hffN0jiQpVKUUrZLkc2K65jYPJ/PRhlVI2S/B08idPOWmvGT5k04aT7dkC9u08A
iX8Vkruh+TSkrN3Bxt/s5U/qR1Go7uxd4VOLxR0ePIHFNbf7nnl60n1oCcz079NX
r9G0/H6mjQs1aBeGHO+NryErSNWozcUWHvT7rExKHN1tX22k8bPs4x92FDZbVPUm
jN5wNtQJ3qy9z9buTypmk+y625MAbwkR/za6RxItkiKvfYO97v5bgdi8EkDgnfu6
A7t7d6VIk6uWJtNF6JbDZmL/F/WMAKshC9ThdTnkbyn8S4+MQ27A+tvCr0c5Smh4
PaOVBcFbpSNZNN8VygfeUD9rcuIVrkm/xUD4Pi3rIAtCDSnrroZp/9YJXv1ed8VY
Ecntndg8x6NCJLE3GMfWRNLUUMfQ7moAxcccmj5x889HMgPiZkIqRqGkNS9f0gb4
Fo+EtPgOKZXr9XuReX2+sYC3/mNU5TFP6E7Em9goJT09GIgDzSYTK/KszgnnhRtz
aHCI2lXiotPHRcZJvuUQf+BN6PoGLCGXRmPVoQXCZ/3REG4hM2wbydvi2KZ1RctH
xNnjsXps8DfOdbubrUvHQWfNsC8fxQ4Cuf82FctWq8uwyyneEJdgY1sXGUwOJrWh
5qGLyZjFuTqINHZ6ENvt7FKelLKCNBBoZB8yxxoFsROquEsHZeiGuBOYRX1WCHeu
sXvHilFAOq1/ohDH0ja25cTM9r8uWx8SViZkvGE31r2pyRIVgONS902RI66tcdTe
pFItTNaRpdrE1S2jQP/0HDb3nf+4BRtIhHwgh890ZsyN9uKLXUkLNdx40oL4hquO
WyBFyg0CwOv+40ZaR7opFv0anTkRsvyG7m7RO6nVgefOmlsPWPteQBw3+CF8hjbS
cYPyqCIlbrWR6FSVGJX9TJNZt3JM8wKHoSKnYfdKc3wEdrhx7T7xV7oExxvvPi/Z
ZaN380aFA1cw9b066HJaU1r5NyFx+ljuMahSo4jdXMIwa5IpFGUq+UwqNOTftzu/
qMjrT55ewCRMTYdNO5/NKUYLcCy9H9vaVxqN2ApAiSLPWhosOc5BK+VsB7n6m/VF
fX3DzGI+QjWIDIXXV7Yc17+oHc8i3iJDi/LTpNNCn7HqFPzO0xlOSzfme4oPhmgx
RLMJeZd9Abay7aH90u/r3cbEc56aGs+j1oRV8fTr631wy6dQla5QMm3e8tOHfk+3
yve9cQvMYzxageARpb+VELV0hagBUpGy61y+fwcjrBBxyIujhY9KfCzfe4CLE4jb
Zs21kbyz0XlALAQc5TwRSsp22fYK/kDOpeG63jHPOjkN9royahii/kiZGUDaa+g+
UXUmN3gIQcKQFrQqNiZecRR70Pz33qzaS0r6mTvHYHObW/2WzMBaafd+RtmjX3tM
hgkISIjmXX8ejpPtkMkbqAKF7gIaSS+Gq2VxtrO3mBbpVWmRG4CsUjFxlwzVQg76
cKG+venF7UqZdYuOmQbiE4rEhjY/3ARDR0R1bTC1jeaQ4994/nWKJPV8PVm7RUlB
jq6bkxQD7c5CeKqNcQdrbhapG2ZjsO1fwdzkfX3BhS0AleHyoji7m3FE4MTwmTp2
GUH7MfSmfk6g9SwCZrnzT3cNFofHwAWB+SZM95130DSUWzM4EkFcBnqBeU/CWM+J
ISj3PutNWvWHgJ5Kr/Edmb5xLVKc6xWel33yw13+PQylf/4GYJHuTHW1LtMjVMKZ
uP8fKLNe5PK/nBr0hi0vXuHsuluQwBzzWOs8KyOjIkK3X0m9GNfXZGLq1cpOvsgb
NwLk0IZ5xi1rxSik9AZEJNXwuXfjmLyLqOq7Jtkjs62e83vY/EGYi4RZ3eaZqQ4v
RwC1F15k4Q1V4HbiTO8l0MbRn2xKjji41r0rlb8zBz5vtImNR7KYQ7ijlv251YAv
W/GQ+ADkKYtPdbD7oPB0bkVbjbHSpHKGvVipj+mj0CgjW9Pirxlps+9sTs/Eubh1
S9OibArqf/v5JEcEjll5m0qo5W/9Uke2Ix3CzvFQdibWjwNMjc+UscoRbSDzjxPC
u9mFXJhUbtUwgmKPDh07VDqMXNG9bup/Ez4HHSZRz9A1CWZZG0MOElIl3Yi2Nlcx
5YR/KZZRMiZ5JRTwlPBxFtJLPABO1K/OaYHKzDMFBNFnLXoQzsN1Fy5dITtPKXYQ
alaW+acVKgK+bG7Rd1VOi+VabuA3siOchinqq9YpyTjZ99eTT3rhUKdHlBQYMGVq
xNzy0W25suF/ddGlQY+lXjVZr4Wypa//mizrcOwW9+GIUTjSxz3+trx0U2fcyMsk
3OW7uOIGsIZuLILX/PPhbUniqmXHqUJ4Gjy0O6S0GF25HtLJQpDUu2OVJIrxLJS0
G4asq146mjJnq55Eu+Ecm80nRXzyR9SSOpOS7/bpgKq1j3N8QJ6KSLmpB/QSe5c0
5zt9x97CpzrLXm9khvAokdkyore9G3kyOsMnSZb58Fv2giuBBc8BaGnSJHNZNlG2
Pkch6sDQug7ctCyz9wT+ThNegn4+d6Y6TyKhJqqIitzS7r3ItifkbMUaCXSEEfHn
xTzbkY4kGJSiQNm5jtTldK/56/DKpp9tkU5vlp+jZcbCh1rL7oJORt2YyUASli8O
bM26hIdwlHsKtaWMzjTSH/kOCsDD2PmHNSKZCkRjwvrmnXNSzEnai3QShWxd4m/t
PzaBWWQQhbSk5Xinco9aJbocOm/rd1FH+Tuy8RN1yrOwHy0X65Rwxhf+H37kZlBH
xeRu7AAn9ojWu0J5pFI/T7tNGJV/NnjymEmGf6qTFjRxSlejKbm3cIGgiqls5JHT
zGOr/ss2ZRiRV+hD9Vca1eYWPPf4geiurE3K27xT8vpBNWjqWNIP9WoUq/bDekeR
f7QleK4+abW5gfmEeh2031P1mSW4Faf4Kc2W0okDfSNp3621FbqcV1yAKDaOboI4
5EUwD4CIfIydDsTSFAF5hYK1owsjBx44IboPEuhmQmhbVL76Na2+BE9hPHDUlAax
nBKJavyTyns8aFlbXUZ6s03ZfPqTh4BQEp0c1GMtG+qrptE8D3ZkFzUK+bvbNEQ3
aIhUzKbYD1WAjAftJqr/sm4GmNoK9IfVlCIZsvtceuXBm/YkErz05az+gGlpVmdj
gXS0HsmHgem1JIY8R9uynvAb8OU0rrKqCwjGgCK/VZBQgqnPb5sOxsQTV9OU8n0P
H/HZewV89bCKd21zi9TaE5LCya0KKhJaGUzbAEgFYCRX9HiEZ6Id3m438U4v9C+F
wd36yuKPXG00ltPm5jrDeZ1Bazy4FbXCjtDHv3l/PcQUbmX9v7PZ0mzu3sInrWuv
YHM9FjdpG5eoEFGFzc/WuqFcQxtXDZgdqZvDxJzXi6DbYoBGQKKo6TzCVPsQJi6D
8DUwonlJorwACTyJqy15a2FAlWDZ/9EKEoYuUY+9jhoCP0v71QbTyRbXLj5Y+jKV
dsgCWkySSbtUtIMb5hm0shIjqPczpHthhVkkFqhrthEn+jD8rbtMhs1ganSk7UwT
/Y6buim9Uw+IH5wraXqT4it/0NoBTaOkABbhUKy5JvcUH9YFnvwYXjE+Aaj8fA4+
7NpAg2lCPpdVtAjjkCxeyWHtBPE00lJeTpoqt9plYLEuNL32zg0GtnU2UAImJr+t
WLoCbFD6JDEm+zVpT09ehWXAnXbMd7NuISx6Kj26GoSaCTVKr9niH1E4T09NPfNh
Wlq1JfB4oZ0aQ7pQZDlxkNmzlpSMafRZOlhNktMw9ZHPfHmQv1BAS17SLoloGo8t
+ePs7BhTeZesQCK5NhWeG9HbeeBLfSv/l8IwO1ChqS2j9A4spA/+35Bw4rX/Du6g
I3wnbtzdeNK+nQivzmI2NV2HePsSWetdtDJLuVrZug//lkJwx3KacvIs1hVe1ZmI
DcEAY4jgte0FwQYX0q+G2KKyg0QpH357Vo1wswjhJL85c+nWNm9w610PCFeKANOp
AKRA7Djc1RB2idFjn8+HShM/xXqUFN3kq9C5YQle7kja8P632g1YNn3/a2Z8ECwk
Za4oUItsDC8ThQFWJqpR9/7cugkSoNjYFt67TKzgravDRhFZXrL6iYg54xWbi24b
WirlrCdB1aiT4jwowm1ZKXGptNZo2Waj4/bnpliDLaqZWcg1G2M6XKYZb3/Hwboc
/20QCsNpofckchzylI0ImVBvH0oLkQ3+IsppK4VkI5Nsco+Ec9CssU8Qydot7p27
nEU2mjoZVj2oZNrZoE6gjzx9GR38GWXyIMKe40hgVYoEwt8UTtzWY9swVBwN1JCl
XSoOzuCX2ApVb0Nuc6VhHxt3lT5JMQDpgGuo2PcoIWWyzJVxVhy/SgG0jsUy/578
mFVEe+0tfkJENnih6lPFxudaqW+AyZnc6/h9hDwWbDiU+eUHhARuWSL8Zj2RKvMD
+iDK0PpK6w7/q9TbTYQExTNAh0VdsSqRYgNrzqXYED07Otj9wZm3IFu/3gOVf52u
fNrv+tvzdIE9RLOXYvPTeLQ4lylv72eoi67fySNjxzYSrgnjV0g73LAxSWSq135z
4mhDjpXbobIVSrJUCgQA4xHzpbuDFitSwTLAYeHLYlUBfivEfTZ1ag2bb0IqJowr
IPPrbY1VXEJQ/Q3uXh/hjVU01jXj4bTIbLJPrhKXH99tj/18U+zBfj7/wzQ76CHG
rerV+7hQlfnEotTyYbPQqKRHOnL7fG7mbnK10s/IM2zORFfFYIAgTxdseRS7lekN
Rq6Hi4veh4OAR9nGTWjw7Pxa6r8AGvj3jBEtYMWLRnnGLwkcaFx/B7dMaZMdP0VS
xXAJljWyf39Ab6B6muQ7pDFhF9zQpaU9Dq0eAusbNlXgQmDjipTNK+1bE1QVJ0HR
0x9xedaWoPQCOlYIz616SwVc+aST230LESiK50BHhWI/awytJHz/+nNmzhtJBXz9
KrUeVoJOgWVcWhLtUiJHcyiOFk7II8yJjzrx8InV+WajG+4McG3BOpioLgf/3zVl
YItGEIhY/b+6C7azb8oFkK1ImzBcdbWTOeE9MAjtZ0y0UdGqBU1vEkXSuZVnEhI6
2QfZHhpZ/axwKWAPMXtDIfV5JCUva4BRirwIeeiZRaCKXYcww0oU1pWgBnW5jmy9
ZNL550cXLNCRkQLJgKCwALmE2E1h/9AaWh6UoZk5Kxv/4LpiKhopZwvoAf7uQmPK
d+B4sSyQehKm+7k0Hp+Mc/JN/yzVlrIPpsHKP9EjSlKfoFsGzKPU2VOoMJhP9CP+
IL2E8bdaHZyizWtJPYknbhDYH70njf8EE3RLq3ztkC4hdXYu1A8z5YJCcWnsco4x
EyQTVdJOg+Bbx/JnLZZnSA7R0bX11VFXPoGXD5zeKJAALfQDo7QJYU+VYVCr6AbQ
K5HgENizsPFd26+kZCVVIywuo5YZzVSvhZeA9sTLZBcGceLl9/UEBdlEnblkRblk
Kzdhr3H6wXiBPl9Z+kQYb7k0EwZahMTuVg/67SAkGQuqTXzjZUMmYiSHlbswo+EM
Sfhg+0Zi+y/G7Zv834uzucw77HmeUlANhepDsGgruRL5za3DTGRGNyWB+H5xpvUs
pFt/fRSHgbjyRxoX933IrLesy61cMyxuGGb8i/DZe/d1Cga9pOrAKLI0AlpY/HK5
UgV3aTI5pHcOYvuPSlpBYDPnWhA6O5F3PNRCTs8DvDJJFyj6AAPHUjiZ4W+teRoI
Jqf9ZWIGNH7IZhlJqPNecr85lKy44PgeB9vrli3spIl1BiJz2Pz7rlLKwa7pjE0T
ml9EPwbAqaU4ICV3zc13tJ9AwmyL57Nz4SJLJIlvnPWWovTolXqx6IwlVxa6RjFv
/+w6Bj1WYP64D7rqBQ+0831lgmKJakZxUIVab3plPAg5MFyZxEaA2T70ZUAmxKa4
7LlvHSBrP2jzbK3kpRfoaqDmFjqbgTvCtDW7Hpve3T6J8tWjqZqWmdFTqejkgpML
TYW2inD6qFFNU9cR1IUKxqWGcGdrOHhiah0azhRK2CwKzmIO02PFiPV0PtYqC4lI
8kOHlBGyT5s5B0pYOGDT2Faey96Ylk9bS/15xajrC7eEcDRqqgtNdK0G3yGvyq9q
7WwR21hj01aChO05MCPSdsSJ/amOfwlGQ8tjH6stQSGrRPNTReB45xnXPhJCqhI7
XVM4iPnWb2mNH0i9RIDYD1ALceV8lkcsZA+4mXlZa5QexeUqD3f+lkWC9oBlg7t2
TyNEGx6x1cI+4evMQA3GNkE6gx/zv+MUdyR3c1Skwu9+OU0FSKcLOfIBzZR+5tgP
MeM2ioUKkn/Bt7oJ4sLTqCD3sUscbR28GtIRFqDJnohx7ZGAtUgbmCxygCggJBWv
Yq0KNnu9cVjNsiiKwwUHl5DYdvVECDpxjk+0VvNJTYDJlPOhvnXI5xVY1R2fFnaq
wGGlaFmKXM+o22+nNfD0IqpyQn6ytNgrDEa7Jim5H9G+FCJmlJC0eKaqMbSRCZQl
SMwCGCB5B/uWaVj7+yEdk3mvs1fKY8a47hZB/vDhTDFEUb2k3j6uq106K4/PWLZ6
7KCzsBdOiVDxUjwfz21BdiHLgKPN6187Kh7VpCpffseanmjiPNvpBCjeJNkFVbgp
57QOWjSq7hyIYFjBdGRTQL0/xqOGUb4QPa92Mn4GJkwiVu870NLntxnVkxw/8Zc7
QjErdjNl5FEuMrHYV8DyvVvW0irp3kB8Zjfdi/030pIsILNsGPiFGOSUGEU9JJhg
OnK+DXx8abQHOLMpjkZQB6xhQdOCgJVpWTXkyh73ZWRurXP6uKGuXVn73mCVQQfG
MmtLnmHM9gnMu8QvFD1JzzL0NfshL42TV4zGd1HHGPhtFCI4XwMmdx5qMPFBpbvG
UrHmU6+e5j5HZlqIeOU3noyaiJCUvoXZ8ly1hZO4/DuO+EG+YwCUpIzI+oAV+Bea
bccpi/bPPFSIrOA67R8+Ca1hEE+yxvdqPXWfqnMCn/dJZzemeYoisMeDh5tbKXmX
Xt0aHz9d6shVsyYU0prLaHfVCSqF3RMX82IMQHTq6tbl/9WEWZG1MgvRxpkJ0SGn
mv9Z3VVZxX3bgvRL9k+14OvMsOqAgpbm2tLQ9v7AckYI9xQvAplR5SvPJtaERgER
Niqu/V4RmtE6wIOpQM4ZNmAaKSuSv1JBZxOvjZcxv2dE6T3VzDxnmZkRZ81SJKyy
/3velzKjK4OwOpWLC9cB4cZkEz1dWPKvXEyt+Gph/5ACkoQkeD2EJWTHJ56kJq02
m3YaqifJb0mVhcBCmL/N/Px0HTLlw+zsa0oozIt/WZYN1eG6IpgYAMC1CIor6rNT
gQDEt8py6A32LzVWBEYBn508cchuli3sry55lNj26BDDCLR1qHC0GVBVs9540szx
qvuon2iHMqI2Rm4A1rvoi9aTQsEEWttkEDaP0jSPVWnxc0s+Vq/fr7emX0tUEBOb
SufZ7O0VNA4bjNkVJaqsoQP6WLYhGaEwOwApp41eXOJq1Xuvm/bBNG3RLIFyl+iy
IJ7Nl2QOL0IqibqxNROhsheWK86pzTwIPTaCWx7ptFbsPkfmitFUnJmJx7nCiEY0
/fth7bEJ/eT2mZVSYT6qmrp6xU/+PBJLjkexIoEbVmK5rXrQXHQ705b17AeJnJwo
VwGQnccmC+Cly2nC9irq5g==
`protect END_PROTECTED
