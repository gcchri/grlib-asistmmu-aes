`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hyZm4IoGrsS5/op+u85CF6epRHVDKJ4bw/wM5sgTRQsra2aIUMGuq3ArG3N8QtMg
KujYeni4QeoAjDB3x60qyHhlPnGOhoD0H6sSr3+w8gHIVFCYbpwZFzQtC78xt+yz
RzKB/vly4UYYYVIVopPTG9Sv2c60hGQ+DmUmzIy3be/ACav7E+ChMHOXHT2H66ol
0rzP9zPZGqqX2mHjbPOdVdSXDTOm3vzmow54u3KKyPXS7509UgJJURWaVBz7p/Re
nSzP7m9KRDOEM8P6937KmosPd4pRZpSYt2anmEeKppHumNCldv410rHtmGZSGuIG
RDLQEAKl4AYCFFzrLYBRrFklJ55DHOAD/e2rwDZw3eH86UnV/tm9u6mj/yzfwCDH
mDLgW9FakaGw4uZQI8ohRcsRhkLqgzO/FuFuVSxgoFY0a1X0Xn9zcSYaf3tJ917P
UH5Er/S4k36e7+gbQUfNQ+j+KvxWeoAV8+kn4CFpImeZ9mpwb+8E/NSRxOQ9RbAA
lwqq084eoUOmBqg8vhANl1UFac6MeHsNzB6C00MEr7O21Q5PXjWJtUl387EpCfyx
MUvt82pAKiuiM0a5ayuIZO+I6vYocFfkd9KPcKxc5PCJml2TPsY+oYmXb6HzMDue
4qF0okVJyNRwiRcZwb75jVUDVkb4Imm3Vca1Nw70IAin+L6jo34WG7MFUjx7XVAk
bgQPAZibKpnO/2h5FRPw2SNl4w+blOuZF72uWbYGXO0PXHkWhPPrueqt+YxfGrUf
necvkgQHTUjJMQpersWWyJ4B19SqWoQK2d0WY8au6Fkkau93kbtgfmZHEo3uxLDF
P9rvmDjcz0B/N/mrjW1TVNtXLfGk085gv1KclV8YSI5CND+GGsEm7IPKMuASq5/F
A53K6UMOfwGHh5IwOxK6J9U4cpH5gTNjLu8tYw/19kPz2oRVMm6845R94+zwjNRo
n1/BPTJLl+lYqwcavKdDW1xeu/0Qi/Np1s7RridrsyOw5kgDLsNlkR7L8MId6O78
Gn87Os8IRLrVAInN0Sh/LAYGViNmqGL/HNngGUsSjZ1+3ioQX9OXyldNn99/tfoG
3ODfS4It0OVyk3kP9XjqBRZEM+Wklehehkk+FoJ7TzXn8eDcMBL6re97hRCTf4v4
XaoaqRaBot8QKrbqKdF0DtQnBzAGQWj8pmXOLOPvJyO6WUhbV0CpoNC5VAYzxEOE
XRSnwewjRuU0eaEsfpKmZpGkkwaxOFBKMRsOeXpbtc9FBEqy6aDL7M9hGCKWLbBa
4uXSapsxCGPqzO9CSGoE06XOzQTvGMsMDoGBSKpSsCqcnw8WAgT+9iStkY8IJtoz
1QHXhDU5E9MYCO4DjNdglZabA26pTuU1wTx85xH/6CTdcggGR6VjHDqGq4IoySU+
67Ep8VkH9vNbsANNjFwR3NB6ySq4wWbgoO192cI+AHjVE3ErSE5jSVDem88bDBC2
mNz2e2a5NWfP45OEyZ7/g6BHEnu7mqpoZHAWBW84Wluwi7Ie9CgwaoTIGfPNU8m3
Abr9VdZvTeyOe6R9H6AlZgeZ44HVAvjXwXBjTQAcR7kWrt/FzdNU+PITPIfFrLE5
BBUFp0zbnrDi7YOdIH0k0NY2cGgxUGHodT8bsztB8dQjMjypbNhHmIcNgln0cEvP
zTa2rFsXi6aNlQKKvFpa91sCdCHuGON2VDCVD/+r9g1OgWg7A8OZkiJEPg/0pokz
mMV8NqPXPTP/4mKlYdvYP0we5HTQTGas5e3Uh5SySUEwFuE9Ypr5pVDtMcPzB6ti
4ZXrG/AHxAVTDG8yiuRHJJkloOHl9mnMunsbPTmw0LhC8CdRXuet1BvPtK57C9rE
vAmIJ99Z4zkzTDWs/6AgxhqlPFWshoATtKRDuYUc2MUpblEJcmzUq7ZvtRgUlDQC
n5221Bnevg5n1rqW2kXwSBB1RqF3/nKZYDzpDRHtuicLDP/2vHIJXKGNSo+acSBG
V/VOae+6/8/oDqJrBYBJPnMBsgn7EKkV8iD9cUK9U/5Wjf8P+xIeODTR0wU+GsTY
MApy8vvM3HZxSEfUvv4Af5bluoprnPXxUM4OO702Q3ZYQwJEOwsJF3IP9npGJKPE
2cgYpGnESg/3zrAKP1YJBL2G97IyGEi8sQ+X8eLZlDw42XJYwu+ZiN27F9SpPoUn
lk2l1sfQvVwEVcW66ik01vl1Cs9MazSUYsg0zOQ/BPi/ubkhD37up2wnQ8CDXzdx
3BEBzXgaCO34Thi7ZvpPw6mnkjwg6EyVClQN0WKVTzaF58rRSJq0q0BKfauyfPRk
w0L+YpJSQ3SbTKFaLEUQw0DbPdvsq5fGmEza4xR/7GCcNEkHTJS4gtZEN1DUc3Iz
I+nRp656ra0Ls4POHGJNnY7sHc8zUhutNnlJMfoLN61meFsD8F6EwUOx9Jeaut4x
WQtiT7qfY4V0LVgcbMy34Pa2pd7RK0cr3RcrC5mcviVNjcQiMAg3EAwXJckaST9s
Rqb0mh2qiK4RAIywjAMUsSTD4UhqBKhGSA+Tzmh3FXSOs/zH2gS3RCqsT+CgB7Q3
9pN89NepJBM1+CD+x2xK+rKhhB4NlyE2lwTpAWbfkEUBO5W3TYDC0ARO6unxctNq
qhzK9w6cjb3Sh6EuqXSDD01d9P/GSaJYrcV2Gf3/s65NVx86nvA1MbgZUuVtc8KC
0+ewt8kt6TwSE9YgRh5pK7T7IRxLn/ki4DYyQh8HpnN242GRWGrH+41meZSkHtmu
1kdrpgaCOmSHuP3aGSeKKj2rdKf0LH/YXQUAnZolJW8Z0lNQppom5XKkEG+2Gdb3
8uMAJ4qgZasr5a1PvoTGxjFR+ai0lOAbnEmjYHAe0zpa05HAJMtbmKmwtkqYwkxv
AupWsLj6ku6nuQYunRHYDD051TQE+c9+iRa83OsPU8SStuQJz9pnC/t/8lTLoYmt
8T5oBzToaqSY2OqL5RXfK7/JdoNcUj60YlGDsFCFSBfoCgALRwcKEafZQbvfSzLU
OmDjjJCq2eeqB6enKc/v0GbcaTzq1ontyDs3eez9mwXfz1vOwFRyccuZ2EZ0Uvwz
Ej5VeF6iYxLwDqg4uOL3J9XYhd78vyfQVAt5OpHopLQa43mshFcz1bIfXn9OerPg
632B217wsDKQ7V3EWDXQUJExOEcm/5IVPoQYYUzm4zoEIPSZGOKzcHk2DG8Hr2CQ
/wDwRnb3BjEfrzkVxVpzW7qMq8X1gAgfW7oVV0ohOBQhRt+D9KHMz6iRDgBoLIuO
JXnjlQPujiqWKZyUvO8hRTFh741AGV6eBOaVvyb5e8X9fZeAQvo9J63aDclf7DRX
tiGxKscnNyNb9UWXEigBavw+93FVQc1AcTINBxcA1sPciKzoXJzJCzMTGr/6NLLB
iD7/iOgeLqdt49Mc1cZn8AZJFoEbiusi1BKSw2uwPOGLl+l3qkZ2JdIxOFLx2Ckr
kbljKu8F13DvE9crcIcTcyIMVa8YLdd0Cg4aNsLGguwfnhUY0p9okl2WqWjdhDLC
DGukvLBnACv7LdSZAE2+emUNk0UauuU+Q1yXC81OBeVlse29v3iK/iC1swZlxQsY
yKw2rq8d6NLarqWsjEVb+ZjxA9EO+iWV02W8byZjaXkZsZ5AOTNF/Ad+RSeoyW+H
izwS0fJXMJzaMyVCCy7KOzcaOeVG5gAPrKOCnnnsV/Blu5wxXEVsu8F8OZqklu36
1btzhOEBycOXD8QDEIfYZ8OZjOPSIT711W0yhdoI0yZMYttinOYFTTfuWNsjRezr
jsnfiFf/n1z/O5bzPTFu3p96O9UIGdbgurpYPKwgn7DUgfYkZqCVULgBKVQIFNu3
m4MdqaQ9WDLX8vtTLQf21B5JFC8H0EDSr99l7JZlPah/gGkTJQ3BYpVs0Nikj8IN
sL7ycQ+ZhXSJzhxVxBR47g==
`protect END_PROTECTED
