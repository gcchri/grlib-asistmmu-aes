`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sz7+qmJeK5ReN+5zhCRVHPRzPob2InLqv6VUgoQr7IS0Q2ZQ+TaFYNS2ufQC8YKd
htVssVBBJ/GMRM6ytmwjRcqcISgo7Ep39/RGu2iv+sy9MF4JYMntavm8X+U5e43R
IuRLXRdQC+VSmlailyRK25QitHyZV0UARM7RWnIJtmVnqvlZnicRcju04hVN9oXh
ud6uwCqcpnHhdlm3fIhHaOUbswI2CK00OLi5n2Hzm2Sdft+jmkouiq3z6kCi51DO
fe3UJiIMOisZkAg7qszusTVwOWpJpIK3CY/NuZ/Rrck=
`protect END_PROTECTED
