`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pJKIeXqsHe29LPGCR7eo1xhHmYMWIkIHnwHFi8XX4Bn1/t+2M+k6lswBRnkHPzMT
zi+MkPsDaWNGazMuNRa3I7fpZsexHJnqLT97kqfDTqiF/8zTzXW8WOgLrIMjMBtz
fqYrsjYT9Fmq//Xeews6of350HbmujQXkPTIGOdw/o/nFfwKeIJrcUIWrktjJIlv
Uko7022VeaJ61Te5MBNq8MjqdHI0xcZILsZbj8CPljL54AQGJpHBffHeb54HBLxP
yOoPtuYoIeVqYtMt+Xvpv5lLYEkG88YjG+LG2tWnoBpauQx6oBwd7L03J4CO8KKA
7w5VpU88Z1cKmQxjYv6ycQ8iQ28zvy127sK+ykh8RmxvnFuW92PTM+tD+iahCuWW
J5yYZ+fLvLTyYvm9WZ6izp1ItQOJNnF+m7ixHmNgJ+oUrZtqChxxIIAn94K08JBu
xdE7NW4Z0REYLB/2h/CeVJrFCiWD4ZyoFfuL7FM7sk8IYa4WXyYbGKdwHCLk9yQK
`protect END_PROTECTED
