`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mweNH7qX69FzguhWz6bEQLPZIkkTs3fQpPS6XIJ9wwsii9ln3T4RGRweQa9EKEeR
cr+NDrSpXOWj66RKm8n88f1Wip0RpKy6cy8wqXPo4qlf8WyvwrcirT4Mk5zwGtWx
5YIqTmC0nvsF23NSbmDdM0iMWix25oDnLzkbuBZRv5Uyk5RBs8WIKaXIE+X9Qyye
OguMrMrfOSiMukLkRz/K4KXndfzCpq1VGUOwi/U93WELQ1gcDeeumLmzNhnq2b3W
+nNg5GqS5cJklgkgWWLoHvxRQDPlJgfR+2gCCbXNFuJmcCL++XhOnWm2d3+sB8iC
AmNBQC78M9CHsF9UY7aWeeZz1Ykv5oSD3EoUQA1LsoRB8LJXQlFZCAYVbp3THZNo
c58KfB0cmoNQrNJ8FeDtRXBeZnBxn/pswNrSKjhBbtJIIpD+QgX/v5Li45xz+D/F
ZtvFCBhqVuuy0XJg9++3ZgOh159rsAkVRnBqTnYp1uXEEH2kl9+rMwD6t5ImtA+N
WI8UGaXj+Yo2Dy1PCkvXrtpIkMzxBfttDSenb9NBdztQsgSav23+CplMc3wZ7ZIr
Cipq5+k9EC9pqCTdX2Zwv50HZ1jUc+t4TjEJPhL4DHqfffjOJYTbtDwSUZcgyOtg
ccwSqa4CmON59EVMjPiUbCN8qk2VFxZln5+/fj5vHfr+9nmT4e+D2hWTn8BgYrYQ
JrwzE9aceULl8I/BIKV73q1lbbGbBzNU4GMzBoyi8ZY9z6rDS1kVUx1a/hH8gDaO
/ZWvKS8NlugF1lof4eK8HB7m4G7fIm5cFl3h9B97pVwQGh1tzG67reshh+/DMTZS
+229/l5/89Zh8JcTFv+ofQ==
`protect END_PROTECTED
