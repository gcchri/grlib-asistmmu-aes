`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y6DX0nSaHs45fXEPXtkL7tc9F8bQxdeVB+9CMYKkCX4mJ034qPp63jdWaWXiJVip
0P0zivlI2GHUep2iW1YPB1eeOGquSDRLLL3fKUuT6EZTxc+ZEgCViaUzNrKKn45Y
EFWHOp5KK+lclpbOQPmZq4KmrFxneXaDCSTcnsUm3YRbSihupr8N328QleXjfhIe
DPBatxTfHLF7o4vIW11DrjixJKS/pWpusDWVUEUddGjohotgdrakSz7BXabWLJ8w
8Sc5LE/Ax0xv/z08KESZPuN4bBGoTubweaJouXmj0yOURRn5OSEs4ZKNimnZi3nN
nv0nJIOZIo/TeUu5qaP1xRlkZq1MecS4vnA4ESF2smTVH4GJth/eUDGoAD37qvud
0QpU3SVl5icwu2463VErRES3KmXqBMpgTc0Ys1FjlO5XUtG0Jfs55sGMplURc7dW
sqYrCmhWybc0PwOFX2LG1oAz5ffrVHS5W+lJPkR0aOEe2aIIjSKXuVwqNlB1pMj3
e42T8d14JEX8GBJlaDPToxqnF13lPzeUgML78LcTzmTSRTyFJgBdKIO6F5NASzRM
UTk0T027wmdvUmy1Taa3b3YulRVBNXtG+68nVcJ2niBpXCzMzgniL5CX9dhUFoPs
nNLRK9iQf1w//40/oDrdMV4brJzabB07wEEpS3SZPk3OTbwbkF35dgmvw/q1/3u6
aDUEVMfeYosHn0ChAK7mbAQBgu+xVrqkuyVwa7Pu6XQ=
`protect END_PROTECTED
