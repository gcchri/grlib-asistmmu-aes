`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iNxpUlujIYTThOSSX58ojsmdv+/7VyWHPrmgvpCes+l20Uw/ZWnlv9NngsV1Fpep
MYzqSCiRxJsmvq6srnzfw+yMMsxIWXmMTv6Azv+DfwohsOU6HdQwRa7/NkOuICbY
W1HfxtlDua9+4cT8j6VyeBxvlP8DChVn5j1mGqLfpjFOI2yrnM2j0enEUbfrPP/y
KxSmxt0ozkWz0/LFuPOdsFlTgn7wrt8pE4Kni/CrYdhuRtQ1Bl2hd3K1Qy4Q7BSy
0BVaiS9y6PoIIRGP3BYXf8bfOftf8TGwU7mKtpmyQcAo8+Iaw+jcUL8AB9WRnkah
YQ7XGvNOs/Lw1FLVJGXb8aBz7Z4ihRsxTtx+HDplUz55WQGeNui/t286pRNszVuO
t+si21/dzHwjdV7TjegAMxiwHHaS6Lg2pP30k4IZxC7W5JJl14o08fNQRlbk6ju3
PsvpWkWpsZmwFmQX33TynFwh9wf7Xiom7FTSpQlfnl2w5nThDdu6VvtSZ9Cx/uSH
TSDb9kXqcC39pISAkaMj5ttGhPsQWxLCrdM/OVuB2p0WymA0iRsVJLAMVOZQkKWK
YPhILZ+P1V4H4si3oTfR4FJLmeL6S7X4dBxbz4s60K+djrCtB48p6E8oZG5phkvg
mzWFDGmyaDJDkqqfGJREHA6nBJy3Qd/rCUwHIfMutCwXNwBPH780urWJ57G+wJlm
AXE5MNiKlcxFaVrcdK/IzHMZY4tRQXObz6Jnob9X/3OxZjHwuGFlQZo1SAsy50am
0d+9uOEAHzkMHE+b87+oeWo4Eol/dsgfPTMjHimYSvxA3v9jxlmEaO/eZtD7Wyis
IgoFh8W4PwCssWfCA1RBuwqUiXhpgMG03XyC/YOWbw2RB/seHJSJrsFfXUuwJHbb
AkcpcK3GrzLBn7tN/3/uPpUIrU0/54iizFAMrBcara+xlITNiPCaeAVrxXPrR8Ij
GUZPFoYxA5fO7HNQt4Bbggsp5QrjM0ivXd4Kppa0l+HTVDVBEIkOBmMPeQ4DIk0d
cEUQd7qBwxeuK3wQmeHtyc057hlXHw6jqHMnJBLBbZtCi0vhiar7EE0IZFYhHI5w
UAcJkauhLj6JL4okNbeuW5n3D7Ewuuqm4Z/0GwK2vXg=
`protect END_PROTECTED
