`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AFUTdbqSkUaIBY83r/zmwLlEuSvcPtDSpSm4l6QJ5xP84ta5xOxZPzq6JBQTCz2g
AmghVMllNWXFuhoeU2dZ53anf8C90gmIp7/pfOcJV89UZERx+XCedIKJ6jba0Jgq
3xbNxR2e1FVkUmk2GGnnk+SOGv9P8GC3E3034ZvEGnGImr4WDvB7a6ocFsL8IIa2
rG4WrmuDZ/Aqxfn5Mzk0d7hVbbJcTkFDvW+ALYB21cRI4jr9KcGPax2pn1mGyrfc
R7dtoX9rsWRx4CT+IZkRLlMkwOgCPxNmWElzO1u/wFweoF5jiR0pGXVjN5UFSwCc
7janSEyNqH7KRefSbEuNfY9RqvmQ7Yy2gJ9Uf8Pwha6zF4zvvE8d5TUR3ZkiyW4R
Xfp9ChOlnY56hlHgESESnYwpPqEqPsQR1xizPX67/nvajKVP+xZvV0C8ycchOlIr
qrLJ3gQqlFVucVd6dFBeJ72lhtbRvh5TyhyIkudMhvwN4rwzh5S4Q1soDM+yuX1Z
`protect END_PROTECTED
