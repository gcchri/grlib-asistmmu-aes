`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2j9tRgauH0RzWfHZaRzSKjnBCeqtGlctzS9OuNYCbjXa1xS5/YEU8q2Z/9uM3mF7
of4KsE6EkwifQ0A7V8paYxCuWLOUCVzDcNu57C39zy+CvvsmCMvmMYskTEyePJZM
By9GLXL7q+nZq87ly1nTyMMQCCdme2lkissk8MWcNWWjYgub+7RvBwzlvCcg7Fzq
HCxuUxNl4lQyvDZDV47pgTtmSBS1fEOgptUqBm28uOYi+i6pZlbZDVB9Hm2K8Fe8
mH9KgVcPUxhia+w9plrqQ5jde3bNwgHkNs6e7TA0B6r9hGbDY18F0iUCCAHPTCjz
CO7AxEysAhb72NKkIuufrCBRyB9nme1a+RglorjaRxBeTubt4YZfG9rE8xAB2KuB
Oord3w7uhytYSNJAUNeKXJwaCL+8J+k6vQtIOSB63Oum2t3/b3f8FEK0VFWK0NAl
mr061Jd4GXJJbkH10P+hxGvAQ7lN4g0eeMkYz8e3tRSUouqBx0ANJMFOVQ4O+Y4c
t9hIf52WQHgbzUhc+NZF7HPQjgrIe0/CMSQqpeAOwmS7QyO8M4JqcFNS0Pr5gb1s
YYoetlp73Fm16goMbRVCFZGp6FDSYc6YjAWMSC4js4NOyWwIkHpZEp/Rw29uNEAF
PNazsZUCo+3+B9R6jj4c/UYCYCMeOrD/P8RVVaoKlxrvuPLgfFO4BxEs6v5x6nuC
pkysfJ3TWtyuhJJMM1QVYO2S8X0qUWzxNAc9gt5do2lWZvJYbSOZSGjUvcH+c51Q
cGWP/teSi7SO45ycDMedg/Xlz0xbI6JbSXm++KX+d3CHRv2LdnuE3bSLj+qfBmwy
YkFZtfSzD1iIbaxgfX/gXvhrsZoYRRuG3DjL5CNLrSmoNDHqrRLGDpr9ElMMCX6z
s1Rx2d6O6rJ8AjMJMkZkbNKOQIBsenbE8l3QQG7DQw4RUpbsKYjgMURNVdgA3gE7
RTErv4jgDQyQf6nP1a53Et3UnIegDmgZHQuBXv5I3cI9En+798XlXjnKyCa955ns
3kRYYyaH1/z5br2YfzNPK9ORxF3CNcnvFkbzD+6ztAjHqcXS3CSxd2kKsvEni2zb
H9VOLZOrxDwvAxz3x1sT+89KM1hJwrStFLVnglHhaVAloz55wKlvyN5gpcuOXjYB
9P92rEw7wHlyPuX9UDsI7TEYUMnqgCGoKELuRKvsPxAxGgn1B7pimVH4FtCR0ACF
GdnDbxAYHEBpwyzPv/YZtKQb1HsOwP/WkqEmivv5jWSgZSobkhCqTe8uDk5d81OH
3dnVTP1RTlkjKIadBV8oe5i2TIEo5FZS5C+Gk+u3WkCeE7a+2T6EDTajd3X9nPkc
lfwyQMScTv4usotmivrbb5QlppHGtKlBTv+taShOfMhIJV1ErXQQsBBSEu/MEGjM
4A/Hr/wxiGO4yPqVuRAMj9F6k9jl4gbcM+tLl/vwkqOiI2IuFRUSOhfLXZURyvnl
a5RqZcQ7Ld1vLL1LSFS56+AqoGSIs3Ig9tq4vj1EvzJ1vQsGSm/pS6Fdu+xcynpb
YX/m3DOn0PVUre8bYmzjXfhPYrRiuJ14tipL8RfEQ8xral/biQz9T+P8YvbgB886
y/PiLgwfmIYT74q/qFdQ26LjD//JAcRqv6jwdhesSNR96ivmHLAoFMhty4FgYKbx
044VmxTdGT5ZpLdZSiKsix0M/n4X811JmJ63La3WYnwtTej9jEQpCz5gEs9c3L2z
EcITK0Kv630uHCtCs1o/lmOP+GL6Izdf6H/kaiZQtnAlOPMeCuU0iq3niIADaXTT
xM3xYZR8il5+CyKXrosRKV/crBHGQvuPnfvlBKrhIbTg2Csv7zch4Lsp2If0VEb8
6aN9Zgye1L8XQEfG8tSmr/14FW0aBSQeMnaY2eWrCOy9koG1FPVz6/Aro+CuxArO
pBC6f2OhRZib05mdTUc+DAS44XyikqWX3cl7uEQOvWUVOBXI8qPVpjomc1sRLRNY
YrhRUoag+b3kob8SLwDrH9rP0bfZlXymm2TeGfWk/oMrlTwFk4jprGVL1ewKb1KX
fWCBUGpOKdKlKEuLlqpdUEQr+MnEAfxezw5UUm3pNJus0e5ofHOAJd8h8cM4m3vI
drmwl7U5mmYCltk825WiKIuS0M/WLnFcK8XRFUWSB2NCY5krCrnWWHd2xMWK0vST
xOFvlXVzCWIpOGp0hN2B2F9wavNu+j4hvFBFyBywQnwV2UEOkZ3Em1HzIvWMfSbt
DyMxuyebwj/I6RvfbDpPhoCOO5QZJsudt4G3mI+0vC6Fsm0sCJytm7cTPgcO3IR9
sokQBNZ0OBvD8ObozAOq8vVQqzCYh3Zn6p8L11Dtd9Ym57aQcTrKb97dCx1dPmUO
mEx2U1czaUPB2R00oXsgiqmDPKjUhEqx61TKDK7/Om8Hh9PZBDWknNuHaJ+lCbBF
j0W3D8guF6onPz0IOhMhFqnqg5Abou65gLXTkhrfhdBHcfCwMjWauWkE5GsfTQnt
CdWH23szEVAaJdOg39ypEELryAbXS2HfhntVHWtY/cYm579Wbn5WPHGRu0hV4yAi
A2sAHh4ffYyi5f2DVUeKjCgY4h0Palb/BnQZcuK+UNB0sRJJCwj3DoKDBLu2k95+
7Oi7PTVY58DQRvTWp5XK0lix/pgMPCE4szdzWbmPSnphmdIezxyGUddr9eaedZIh
Vj898o75Gxmqes1sR0I87tkTunGtk1AFHRRai5mcj3wAXjItrnAfG8rS7DccSs05
eB9SOndUE26mMqo/vbfNV23YyEzoOsvDWKk22vpzUQ3lqGsZhImbRy+k3HKN295T
ujXHynsrRjyujSO84F6DppOe57Q+koj91zLEFMXh8mL6Wvd6XqTHyjfgyj+NcoNI
gS6p7kpXDAzIOAdH67s5dfzuMQOqkThk8n4u0RZPM6lPwBjtXuhV3WT88z7nsLYv
vXaOUfHjRA8Fkx2zpX1C5clpE2iDio4tLFYRfMI/vm81/BdbMCp93GTpct5kpLpS
Xwag4j1WB93Exqx/G/J8vJECDLZquU9yb5NkY0OtFHa4kEpFfiTjydwoNH+Vf1r0
iJZY+6HrZJQGzA+iWidarqEVd1fuQ9fsR4aIZEvMyvWjjDqVa8uF8Q7vhwDEgXiD
rHeMNRUUWOZ6OqBorfQCtvwAUkX8mXSMMpeUgZwzkOY1R4Ec0jhA23sVmYZ9Nv1s
w5gbMyzfdJRmrDkHMjqhAVKxD6RVTCUzuNMpZR3RJ6I0XObE5P58QEK571lrgP59
6hGMzqBDML0vIXEKbCX+C6u4wD8ghRL6fEDNDKP/RIJfSPZbY59uEdcQhUuqg2Zz
w5P7ZYajYXaNLdjaUW9tLyoPwfOCUXl12O20+VuFMIq9Iqi2jB0VQidL2LNZ9jxM
+lJ9l1gKxf/WikLa6KLoVymmRNgf5j5RcWuM2Vozdgo7bQOatbEpHF0vPZ/O2zs5
+UeEXXFS9lnzOmK/6s1FZTLmEIqEi6jgyAQYGi8IcrndvrmC0FlJKK1kYppEDxYr
FKyjAn8iZMlEz+JvPA7PhbNZbekSzfhbfxB5DMnj0lgoNflpQIrq2PbHL1XyaEJk
Vg7Y+smBAH2EfFDB0wX9YARukpjsq2NpX32WhQGJspQ6IoWfpSrG5BVAVP1q8Q7x
1Q7O3anhshbOzzIP3JQLS1faBJRYQIhPLc38GxwO6t0g3C+2rOWXCXV06ie0Mt5c
0znorq8qFriad9vr9gPcWK5y6Z4qkGn6sxy134zBW9WqY46Myohegt5hYQ3OjMji
`protect END_PROTECTED
