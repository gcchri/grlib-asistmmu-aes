`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YWfOyVQRj7b4nkXf58SvFkwgSOFxNiVul81IuISzDa7dqGaUKzPlX4AyLijR6zST
WkHFnU1vkfR/1usFLPZIsMyPQ2r4R7Sg84eWw4kspE9s/srZX5h1nv3D6x2W1j5w
tbCa8YJmiDL3DeNlVXi+Kv7+HTyapm8Q7FgxNdIfzh3U9w452tLbC3bKYSPjqRPE
It889UEQ23CprR0R7AlJShVLjhYCDbTKHyDZolp/z4F1XbdnHobjKPGNovIX5jKP
D5QBp1Id99K0CtFo8nfHCDTuCX3tDO+wsvyN/nPXqQ2M6BrAgniyx7p8+/F9gHFb
1PNYDjDbmurcGO8Uol1iAP7BlxJSKj37No/QJfqHaD7GV4wmnmA+395bdjMrJjo7
Plk56enYcCASw6Z+DmgRRzbj8Uo4SFzx/bE2D4R4yT+Qnb7letSCBvRkALmnhfjW
8srwn/6Neoc1nwlRzwc4WH8peEGS8T9yMs1b7w0brpUdacOG8Wp5YGox/U5eBrsa
`protect END_PROTECTED
