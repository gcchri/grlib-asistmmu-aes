`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VzcOeKZ9A4cy6Qy2NZtzaz3SL+JPL8sb82G3dyuUZIvXMhWMMBlSM++U4hA/ycUb
Aa0ALtyQBKXnqsREBZYDrwVv4FljJGmrkqFIClgQhVNKj5PI1Hxai85XIbZBHFbT
Y60OBWSbaBuhQbJy+0lA0m79b96bgZYVmImJZVwJYODsTFONwZUi0mVcCW6lSYdR
wYXCJwoZjYHW9rzQbJGe84tSGZdNZ2OnLmI3jhjkofgv0XbdLj3X95nVjEHHV+w9
TnrnawkdBeiFLbf9tolfsvHRMR03HspIVGiuMg02dkRba1ZgGZ2Iac3wZP67ctcY
fSQkAQv39d18ZUh1B2v+exs0GOUGAG3xAFsLJXQE1KD9pT9eflG2HoPucgwTvmLE
OvJ32l2yOS7SjPi0PMYVOE/x7Yp1qiOLa/FG5LX0EANJ1BG/n1gRT1mzERqe/LOm
JTGDG2MSpYWs7CR8SV4jsA==
`protect END_PROTECTED
