`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hjTi8vbnMRC7+tCJKUerf06qJ5pDl5MkX+0o+phf0ofM14K8AwgFv9lXDSdYx4eA
zDcZpk8QkByuoWNurxl6hOEfBiAwC+gP9zpqhO9ueHeuod6hf4wfpVkGzXR990lO
8yfvD4ecr8UTpW2HwK5YXTELKt2Te+6UinTnjRxBcUvVzzHeHDQYXzkCYbEgD2ot
zBTphzUeg9TRcNnFZW3DaicwsBbjAozbH/UZ6801DYGJztWqhAYw2fnQD1vVPVfW
HoGNnfzRCcHIA9TZysCKBUT7aySUr80513bdiU7C2NdPVwcMB34ZZDPk/S04hD0w
8sS+zEbgYE4z749YA/D4e4P1G+nwnb/iPv69c57uZhiq0tqQ6jwLN1ZmfOG/XwMy
mfDERgF85Fi/sQAPtj7e+FfRyYudhCMusatDZpPwdfX7fotFQUpw1ZAs7aBOdR05
hv059YEfNiSkm+TWETgr6XMsrp4U+AebYLDT1wVe5afCZVwxou3ZXiehKN0Jd4L1
hG37I2+XU4u9t6FY1rdW9dOENiZdosX+sEDz74Hp8OGbwTzg7T/B1QcE0Iq5Dtxp
cVL36HxXtxr3uRb9XnvbdjUr3/78xJfQXGe33V/cKeGs9R5jLeA+wpnQ8nJIjDYm
tmyR6BFuB54fp7Nv/B31PRuZ+P06tiF9AYMIjdyYMIxoQSTEvEL0w9WRYvn+V1Pj
0cevwWV4kTPAAEJ2CYPY6jN3riv8v+rmimAupcrZgMLdJDGQOWuK5LQvB3Zgk7ft
WS37Q2/1sV8+EiLK3Td2VsJAdMZOQP+ZPFGJvdk2WKV3I8pLSvvieP7PKDUxg6tV
xAkCVt7ArB0xx+1SbRrqicoZdIdzAx3yUpUfQhbqXSEKuxn+4w2UrKeCRSC/WwmH
69vnGjARn+9pFTDlQ0wo1R61M/uZzm7w8tAGGA01qFS74bgWKTH92qGxUn7y9/nB
8ew0H727Z1HwFXsDBHxZy3nExmHApPOf3sg4Y+UA0f8q12gtXjq/imvzuonmbVKN
V+dUKldtSG3s84riBeMZ2z2cZv/geCJcN3AbmXHJWZb9wD0GOk/VgD9l9in4BKK7
gSvHdaEmZNvhZDUTZFBQiu2UKq7V0kGInR39XyQRdsz++W0K55g2EcazKe4GcJsv
n4nBLEGtPBp52VCuo40dGWaoGxVexezUQkZlxkbiF/3lWrMZMr5y0zde+yy3vsYE
mg29Zl/+xA0/Uzrf3z9VmwZo76g+tx4UaLESw0AsZSb6zEzuSMvHj5DGjkjzCtyM
GLWvfQ3qAiL8ciKb58V64U8aIE3DO9uYWmTFT7Fhroew+8jvZvuMKvpTwxp5/sbd
cR3dWmzJStFzQ9cWO74k+5k89STawzQ/r2hmiG2MGIJrxe+qi5EdyraqEWA+e1cv
Fis9ClGohKCpZdUmBdF3TpDOHf6pTPh9KTd35zmLuT0t/SnMBnJp571+oUzqwlTd
29znaWUvvnX7xTaaUOxHGzukpLYPfUMA6TMxNigPk+uqt9KROrqptQykfjyWQnBJ
K6HmWXWesldkzMz/T7tPYLO75WgnbaAwoOXDog6Zw0zUZPj49fzwa+RtDV0/yXtY
g0uw5IDzpj5JoAEc9DKFkx1b60bpdg80wNeQImECY+WYezKAz6cuLcK3eqeX355f
JH2gL+2v7jN0SdhIiIpK1K6zyQQbeqGupM+OEp/TLe12Sc5zjkOX3DNWFTcbJyJC
oFn7YKxxp68/4aYKwXUiFlni/1V1ZXjzBbpGGU0i2/q9jcxdvbmFrld6dm/QQrd6
2g5Upluf4yrWh9GD7RwZt2wNXoB9PRN3gyOJUaJDo0flUQ02m13BSsVmrHmN1KV3
eoufMmin9rFp+sSUvFox94gywecI5uc/iajiNOMvulqfux9Xl+j/nDRU4CccFkee
ImwvL80/ZpfGMbqjO1NzeTq6Sc4RNM2iyPgFfdglGSu1s1h2FEfG7I/MvbtVyzla
3H9mySDQ8NkqZvQkC+ks6jbh45FKNyswB+usHOSYIMisUknLpHheGthF+zJxPZVK
eSbD3nlHsMGlhwTxP5iBhc2ew4XOhGxE4WcPftD9q5wiSh2Ut9Pbl18+BiMl/SWV
bMTQFFSJ5xJ3a6ci1AJTre5+aD5qLc7q6xwzK8+tHghzXMJrABbZ/9//zjHBLZS/
OkS9lmiEfI1u/LjbKlAHVTxtbPLQwscPJm8h+yRcPPzvEJUglrzLkmGJXNZfTULA
BbTiB61VXKNNHigMGqNfn/n462zQXHSyrH8yjKkuCG5csmhET5mI4+XRsuGE9Zqb
gVV745vNspYPPV6FZWM7QkSqqCrD0KenqUrz0ONkJ4McbucNe9BJbz3tovctsrv6
ja3gIdYLsZxeLp9uT9Y+YqAm9qd1LwFwHr11ZckfYXYFghhmwLGUiRrakCxXVYGK
q0CQp/2Cpel/Zbb/mbRZ4eiIXK9MXG02luEybmR3eH1ZztnLN3WRC5LEXQNGB2ty
CLp5+YlmxRBxnoAa7KEZDQB9f5ctBpXDsaLiDBgstrOrHXppgWXmwzZ/jpb9ZvIr
DHTAo+wpjigNPzOyZ7+PKPlf+C4OFXQTTlvTDF/rb74jhWu3/wKEk98OmHzEaW9e
wwR1UElZAHAi1Rl/e23iAQmxajCS5l93KqZhRfgvo1oJ3RbJyvfQMNbG9gD6j72E
N3PfGiMJCXR8pwIp4gYvw0yVjM8vmGzlme+vFAt4Du/1/D0t40IQyy49noUJXqTV
ILjgkaPZvjajjUoTupYgJ3EJSdvcmbxpHOs2po2dPyu1C5j/ongRF+En4rWjijVL
4BYGQpz7ltl3uaqr7YuuLAkpv4pEm4LQ6h9INBt4gHANUpGJqFtx6SvMIEdmg/a/
InefRDd7ebiCBzPhfa2o3M+oMgQrUYEBLNsgxsEmm5rG+CyTF0cafFn3mi1qTSLx
Ip9EdbnF/K13cq1k2gyisOdXoSfq3CLjz1dmSbLtrANdDHzR/NxOmA9QgYoo+PTG
wNXvG9+6g76mDawYw6cERHVPm+S5oul9wjRxaov/kDIrOMfc/Q9SJtT19WKbk+/8
WaNRrpeDl6IlSmskI/3FPgd986qVH9XTL6J8GMqFblW6r9it+lIzun8yZqPRRNap
J7KhM4f9FJxA1oCev2F3IejykibQFKUxD2msLAlmnQiHUOBJHQSmtpPmpf2mw/+Y
cBKaIoKB2l+YT2CTEziVJOaqWdjWgMnstEaNNx1IwgMfKifaGysVD1cOiwRJ6nia
afXojT3C2ln6JnqQY/28swOXO9+/sPywzrbQ6CPjMLio6WPTybmwJl3UCJRQdWbO
R7dbjTOvokBEkLngSPojKjy8KgJYMN5vlaH3tcdxvJTwrFzjgtPaLfcixsr80u+m
9XlQcPuIDN+LM3gZTIPfB+E8lvcJ+MqX5aq/y5ohwWPvTnz2cKdwvaBx+47B6SM0
wa9bagdU7FXZtlIMh/pG424ed9XmqwlbFILIXaYVUo2v2cyJFzidNamlEdyLUlcv
aTNRks7EL4xrJQ3u2CdBB5RWobq0jN/xuhvLOcPPAuS1/X5qnG5oGu7RBBkemwB+
WoOHls0Xc65jIGj+qbuafhxKfN31B03j+1JWhR1XTLvYKl4ZVKvqcTMk0ZDWDOxE
pOgXZWZusgTIi/8SxjdLpbLx+xb6s2ZoPGiYmDTJ8PySTA248YmKTmiCBBOkOKCg
frr/E+xIQv3XZV9rnZjFWrEP6DUYxqGBcs/C51Vee6UlxocFSfg49ZFXpzHTaikg
FcjBwo7p/nggp0Fh9DJcZjYX1iWh7Je1zcZkFcLsvLSNa01nWBTJ7cm5Rdr8Zy5q
g0nF2A0bUNvhDroccUqiKSnVR6T4xXOl+e4YcQEXbwZXzDCi+U7oHLyiG47PFKWB
8dU7Soy/pydyAcXDScN0el3mMM5w0/dtGpcWFQAkpovgK/qvgzuybkkeEjUq6CvN
Fia+CgganSbwEclBI9E6kaAfAvm309tdWTFTVh7Fs2/qSSpTj9OJx2g8mEWel7DD
7urfx6XnK+oq3RWobcYKnIEiuOw+1wtS02wxf3SduQyNdrwDm//S/TJBdkSrAFYy
q5nU/tWmugP8/5DNerdo7tH5JTwi+k1ZkKxd338IS5x8srEeSTfOn0oVh0jnAkDP
6N0wEu53jlMK1kZd1N2qULBJsbPuvabRQMBSN9McnwK+FKCzakcnUxBT0uCcMmNm
Ub9qJvji8TAmVFJolJCobe8DX6LKJtaWXF+zZAvFmneBO/3Xzm2qsehNarHOADbr
oiktctxyJOm2nXM62fRz7izopq4MujSW1Mh5TlKEvPrnjtNeXoeLofRdkVGwCSd0
7G8FoTrKEwcLA5TZMBPDJwzwsoAv7P69a+MxoWmbTqHtbbrV8hTwjhtiJu51GMD6
F93G+4Yj0Qw707Hd4wSTTI8dQFjYwJFuVFWue9Tlw2oci5dK7jEGRs+Bo9a5Boz4
yfVKAFG6uKJp1jEkMsA/YpuJdqA+DGY1SS1w56+3+48iKQXY89rZK9r2BmncEaNI
WwI62MCUH9CJtKVAVEVdvoXIYminMlK+rb2UR1FRWj/tRXhmDN7WPokutzqmMdyt
tTQS4i5aosFTZv+IEGVybQD0KoKxycQHhQiRuraLkLPY0vCzhlfUFIiMVRH39XGe
4AY/jZEWkdYD8ePVARhZcnkktXMfLHsat9trdj32/Zlz4kOkjMmAoAtqe5f9tOiw
WYY7u996zb0JNIfCeWqwGBS2N4zxBUrTRMIrZHzieD5iRTFF0H8kru6d1qDRTioy
DnBbYCCF/dvhYFUVMs14eQ4wap3H7QWKvmQKcPttgr9EYd+YO/O7z4eq7cl7gMd5
RfF+I6tY/lAeQcLFQBVrvLvxgKxHTbj0jYnBiGoAiPXX6gxwPjlUtnkDr9M5+Awb
`protect END_PROTECTED
