`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cbRMr075hCU34VBz19eLAmpkyvELcOZax1OYkwG7pZqVSH+9OqXyHxhar6wJFlk9
gcqsCu59v5YdM48Hk0Xqwen20E5C2U9RBjv8GbWTlzxGI4KcM2gcP2RshOTF3tLz
0Za8z4gdanr1oYVVByV8flPjNA4I8TUof5cJBCGlH3Ysw/alQGqCFpb81LM3PU/T
BneJvTJT1IbCT/kflA1S2XS7Qwln+ZCOvnvlX1+js2SeW68ZOzKkUp3OIC8CL6ny
fk0+2Wekn3hicph+MjSG0g3zv7pQ341XfDScy6+qszg31bNd6/jhgmOZNMM1ro/Q
kzaz66NiSv09qQh4xq2YwV/uVX7IIA/NUxmjJRMXSZZBnH5eMoXQeUWL4XZWUsw8
NWR2OZFCc/WGUHg7bgo38rWGv92TDsNfLT25/rXuJZylo8C8LH/+KMFCH/y7kI+D
ZSP/vBknZGvA091e73q0oQ==
`protect END_PROTECTED
