`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6UYtR7Md2OGiaa6m9z9Yuz/NBkkatbXy92zuYgz377z8pITYm/2t3lvnEBpBtix+
uRJ58o2ZU/kEx029rHBj/DJU1TtcpT3no85gBr2lCbY0tCpsHtYgj8qslGYSGlo6
tndnQJOycuy7xU9rkMuamutTjSO/gzZT/Xlr3jSa+4V1IlMkHYfXkuM0X/YfAVnU
5ZtkZWCO/EDj/e00E9r6UpeTwqrChLB2BGy+sa2b+cfN9jmmK6fkjfrSfFeBHT0Q
UgsrWINCw5m5HNWbQ2ErFUP7XKo++Ii1EfaZO4r/duD/9aLYXR7ZUbUpQisoxlPV
WbDso5porBuyRky22FvRi+TdmjUHPEOnCbEK5nCc7eDt3SGW0okunDXrqHoi+mqT
8y0D2W7Knq45aO2PiHZvZaJxc8Quchxwy9jPy5BXtmCMmJTy65oTQVdDHlJhaZfu
0amZIQ0MpiweieZlarBxdY2hEfQm4Dc9iFy1/olbYaA=
`protect END_PROTECTED
