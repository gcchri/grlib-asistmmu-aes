`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y6xtfR8MTf2ydUFZrX2lDq2LvSGw9vFDonwCb2htVrkyIDWa6v5MeZpHqME7hzHf
zj8VgShV3sd6W3aL/gV3pljObvlz1CU2rdLMK5Y+lbaf0PSAecEr9OL0mf2biyEy
s1jWFvAJ5QO3doWeiM/M4fTLxR7sHad59e37iNpY8uGfQFIe82dsHaTUrdcMcwbi
HRCDsGcZRaNsCZ6DUbxDe5u7zXAhnnujagAghtJMXoQHXRXSR+9xNqxbVukQsrUJ
tDNI3xzCxr+Pal0+e1ggWEeEqPrG4tRKELrp1mb0LRWYzmHPkluJjbbrfFmPlrN8
z2YsWiRP1GiK7nLN1R+SH6Mi2WMJvnKJnL4NFhOkDMAE4HsEwh2//H471TO+6RwS
EWZ/e1X70gn3EKJDYGZrNg6Qn3rpYvYSlE3O1dx8eHq/ISKB/w8HFWsBH99OVh+F
31Ljq8vs9om8t3Pu+lTLiEoaQuufQ8t7v0N23pc1WPrwiM6y2wSLD9mPwoCbJl7o
lpjEy7JfH7WNDSbrqqiwo9iqbGXCNuQzsHVvJzaU8hlHLplY0PC2A+5DBxx9H9Pt
ujoJw80SkYLcpZOpHBA8BoF+OF0rnj9YN3gP8UY/Ky9yTi/tbBeucsTfI76oGhjS
K+U+PnpagW6gdnwMgf6os/jpQQjAzbgoh+hmhvhi4gASe1QWMH0JmMLvCuDQPt0H
jtSE3gztVNkr1CQ9cw32gXODLtlNm1J0+wJpmmkUwdFuM9Li2uTFvMX7/P3+ILNz
SVd1seoWJdMpCfpfBR+5AYfVLrlbx5bhZVbZtB0IqLdqAIF18X9an13fy82yLy7R
PogSOvI20Kx0pxm5Fq+rsDEbu3qfHey6BVkaWYlJMWJDLYKXa9RIGd7pu7U0lMLi
IoJXGI8zdg11S69lmXx/xTQQSl8uR/hzB3WCO5GyrGh2i5mIrbhFD72zhAJW5H8B
Uiwt2IL8TPhj5y7ncklQdwX2hnXzuiykpKo6sAXRjcsvZToEyIfCLs3ndKd4S0QO
n0DjgvN7w/vs2wmFbLtPZgxmrG1PkHWxJE6sXRyTugVMBX7PUxwK8BvcMjKqv5nM
Ern/qZ6uYK9LU7cmMkIVPJyFJhhdOSH5X4ThiXOZZKofayaiMVw/DWztOHlCTqRn
9Wi4PVuHMSGDSJbrRbgsGb1oqLSKVByZDH2qU/AdxdaTB4j4OVMGgboeTagecxMm
FjYH/5ywkUYOIFsO871d1ue4AVcDLJnfYWQ88noiWBn4+y3bb7S9pgkcFneQmsjw
9HJhyjnWeJB2AJZS9nVDN2Ii0FIUksc4fJ+rZ7VUNtIsOkAnyT6XQmOSlAsC9pIX
bn2zyuJND3u5RDXJGpqzDCzad+y0DFAiFRFlNh9a1Q83kFXnxrm2Skuv4qzpo4gU
g9RAh+49DDrqaW6ytlJjyJcZ+1qSSo+ESkylaSjepDK9YzbXiNzZYQxC83YPrdxT
6L/9SLHnVsxy0Yvf7DLIPiMnipV+KFlN/yLqOe5ibE4nizfU/4MNxbMLCl0m0Ih6
Dp8sudEY0VCA8dj7p966dbZq/1G+etppUC23vVfuMXeKMGjXbxTtQo2ArPvLJh6W
RS71fD5EIeFR4zdFCOwBXPLEiT0ubeEnjS2C1BZR4m6LXg3ZsI/Z3UI7pbGlUISI
t/jD20DIKefWjmw0kU2Bh2yKYadKbiFTgQBqeOozPWChRtBfoUs5LVbhc87GCAYN
XmUmxI4RClmIcKyaHg7vGN9JvgyRL1p9NDh7lqwysv6nSnxgepbYDezY6ap3LA2H
SqxKAStqhwQvImzvOmQvXi1ev+y32wzLdST4AygHABphFFJ282UZy8NyfcVLyMxf
TuHqo7IN3SJ/6hba4mlRnEejgV/+f9zAgC1ATjJg1TDdbpnujYnwunrC/9G6xCQB
1vR4DuR/76FDUmv+pBwIaZNoDbGfo0QzecDxQzs43HI/FLcE0Lg9+01BNz3/lhhx
h9hXUGZvHT1lsWm/lCPLy1hQ9ERQBcz7VVFE+dOoow9gqa7w+D43xqgkF/E3J9hM
zRpteXqBEvw/AzFKAOtRID0zkPTjJh0ufBG2mtj2JnOG5uT72+zPl/nZo3wflgLH
XScR/tqN+M5R0lgbeIrQrzk2d0Er88y9RMhnPARyRKJMPz20gvpfAZNneJ0mtozb
Afb0b8bVix9CnZciQLsA8k4DBoL184Iv7+7m7gkFdt40qAlV9mmJ0QRH6Ulayj4A
lOsbCUyo0uytB7mSBAI3CtuLM2cosxOg9yQCRM9kMiAFfzmxLxwKUDkcFmXOpNMF
yGtOSfCFWlLVfklfdqz+L+Afr48BaHtmWaS9X2t41WTqrfK3w+LHgufiC0ZDMp4R
5xX9uR9jp/cMprA5xvgPE9HpEchiDvskv5d3kDXodZ5/H/h2f5DFd7s7CMaqXyRe
kFD7dAG4OhxIEoenluxUavjwDWH/nab30RsbPtjPXR76EAzhB0B6D5F8RvBAtMUx
T4zMUEOsWW5snBOiBOy4VwinV1i8qeJlF47PriFWSc3Y0baiQ94EwtbdYnzeV+e7
aF31oDaGAFumwZk9MQK0ZdCwwSiZxKdfpstaNtSgp0wYqlE0Vf3Z3AiVXjmxOjVS
55zJU7xSIkCpdzvlTJwiOyFm59aPy/UdlFAgIZQ8e85t+quPmoSL6zfF4WJeNn6g
3VgHqKHdXP5J1c+PvJs6dhrzQsCislPAB3au9esIkQI/yAgdIHhsQCt8i7rI7ciB
2l2lYeXbqKfyUy0RWshIeouYI47e1oUQ5PhXV+q4OHYzA7aiHubjN1OrJ/MuIAxN
X5OTH0YKUTR80z8NL4s55WA6f88Sz1EJ+6kA+qxe27zUtYV3dS9t2KsRxq2lXwEP
cJeZPSyQVvr93nGDjwBkTrkWw2fFiX+uR3iiItHM/v7bstIxe2TZX2mHUXVM+qLE
au5DP4SzVNgW1zoxNaDoC8Pw94+0RujtIAv/UbZiib8y+zdSWIXW4pzd/m/8z7us
UBuzy3znX6rO4Au3tRNM3Lk8f9lprEjqve91x2pzT7PuUAF+TD64n1CgMgHtcjoG
CGmnmuX8khByKmgROh7B5cAH3qDNGtmxvKXJPf55VXEU18Pq46s1h7J/BYSzo4Xt
GJROFYnePP9xkOHKFuMydhfBa9S9IpbxIfcOTMsLWJzcu3b1Ry49Am+8/jXrMOCY
d1WgmUgXaAKndi5mU/ivqp/s7emSYRZshBbtfGC3CH5g/vQHX5XPhmX7PaF3u5i8
2IM4aVdAw7UKGL/rEPlqwiYrHqJlwetaWF2vp5bqlUmxIyR3vUWwutzzLsJXTShy
MTwUFGjomm+wfADbFh/xiK+UMH9SVMRU4ZdmffOo3BUbzJxAcPS5QlUY1mOj4dPV
th5mxTwkO1+OMF8IavBrgbczsv6CkCPjjGKQXoBdRHVELQZNgK1D0YJIrGZGO/O3
elo6IP2rYYJ3MXWr+1EQk9UK2Fg1bg+Sk58kny1hwE4fC6Vf8hmZNuCqw9UBW+jP
WUKOd5beXjTK83GdJNkgprNyOuZS3evgfd5xlmYAAYCIGzJs/ozoHitv3b/yCGIL
YsfjYAIMGvZZCPbB/oDarRUF9rYGo6PFWNeo4LxHie5nJaC3CLxwap+mCQc05SoP
1kw8edP5I40yLUGmWeI0+DrfktXrDKT1EotrYVPpianOFbOR4g9hSnzazGczkrD9
dpv5GKJvW4nBX9MPfWwxjJjQJKLRXt786EkUAO11X9rqNrIGO9sUU73HXxSZYuxL
Cpp7r+7Fy3et6HZvwfXtcjiVeLti5CyfJR1c4lMc8riG7QQAjZ9M1QqAGp7huUtS
m+eGGV5/9dyD5pb2Lu4VtPUBBEmy6e+ji+4rIC0IJc+jnmfSIn+qYDth8U/93mCq
V2pEE2LFgjrs9BpT3elHOCFnPJXtusU3lsi2h4qPx2Y26eYvQXldIioGq91GQWtW
CyRe5NQ4GZ/ivumO5hXzn+jW65eSNQRnUlehs2UppYkY1YRa6zUByhi00VCDX6L3
cSYQA2gGMAA0WghYgNP0dknYki7nlGkbD2n4kQFJXxkRsyz+YTFK0PN1i2jGVa/Z
sUoRvYMbyIn1/2TSMP3C/ppMTOcGQJxRuFl/ji6svoRu3oP0La0SQYTtRmtZ5LtI
yZvhHWn3z7ycJIwHHq1n2Fx2ZUae3hRdVOYhU14OiD+EW3WPmogNrqEqUmthBFQU
F8ZYgEQ80Meh/cd/M4KxoXN9OKX7d8BZ2v1ojr7j//AWuBKNzRmTprXRcDqajsZp
`protect END_PROTECTED
