`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bIwq+Js6QYeJ0cYz4mP6ozMHBnRAhNA2ZqQvBLBrWGEP+sRWmLcjAod0xkVKEFeO
wqC0C9DzVnpkhGtIzWYpUwihNo7gH1gvUOIfOtuWA4T+M7+PlGeoF9OT96a7STjv
uBT7Nc1bXDBcChcWCNc578+KJJuAsdmrJbh9r9pqMgh824rVB0FcgrbVLh6F5o1j
rH8CFj9p5HnmJo0HSnjLcU/h4se6bMlrL5fGd1y15YlVangppD4ymo6Fo1bp+FN3
27ocLnLl8uIfpnKq2GfQ4i9wL2rkHxI+6BtInBlU1084jGU2RWbWF5iKHbiDzIjv
IBZr704nHtxeyelcwYWPeXcrG4tJjsIfp13i/1VZ3yLy4atUh2BOdK+LgfNlVaM7
SsgfluY6jXN0TVeM/FJcTG+ycno1I48JRfrVhlFwDv/Ws1uSMCumhdJupQBDJ6Xo
XGhMiRCAC+94ddyjq5JD1g89VQxklseG9oFEy1SSu7t162pwIk4ByC/Dz8tXzsOF
VMqTdrCPBBHaipVOE6rlYODmtZ+P2ETJBKcTT+E4veyURiXGXW4ItVZZ/9koxAWc
YVXsaGFwGlmg3FPv0EYwpXMGHcFRzuxQSoaQz7ygkhyMGm9G6md+RF5XnQU2yxeY
dUIKZ5edV1keKg8Pu0eKOpwjuOLhVsFX25UEFeao3DA8dlf46BF2ocjdi4P6rR6x
AMdasOqMbzv1S9te1JDUaYWL6tfki0eWSod/gDmT/DVSfsobbAI6Jl1hZHHobmcO
OkWysYNornnEF9MGusu2dPyM6hKVzAbD2WT2/Yk/mIW6t3TvCcZcJ9HxtSE5xMif
5slIzU7mQOvqJioMgKQ9aJ2ozXjRXMZej4tmuc+6CeUqBTjO0Bcme15qDgfFjT81
iDAd9I/JBPThWy/cMqKpag==
`protect END_PROTECTED
