`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
69MyPfUrCPHdK0Tf469C5mstX2GB0sT8AxXOa5TUgZLjfYD7BJXLxAh6yEzwm54l
UThi8txnQJKfJmByFqLKJ7NHWkyFztd4iojMP4DSqEeNW/pcWH63Os1TJF0aTNTp
V5yeraRUBgD15uEqKzzARQC6j5430SixeEVIdzSsvlT32S7Rk4TeBlHYI1y1M1QT
lQLJe30YyY1lWSRTQmYXeSn3pQ6WEXAyvvIL+ZsPZUr8oHbkUQU0RM9XK0iBn6ya
YmNajK6cfrqCsuzdpmWpf3ycUk17iQwcmnQSlwgL1Bs9HAr/keAnUvP45b6UmHe1
1mg/CuaOI8YCibAwH706o8mBkwE0/JjO5wXuWBrYte7qCc2AYx/rG3JNnqbXazNE
Ijr9vDHc7f+aRh+Pr5IShdOSSdjbAyoqPeqZ6oHcUP3UUeVHAvskWkIRte/DCl8e
g6OeyYA63NgCeR1U1XDnn/PDdDjgw6t97fNDDLZWkRTY0vLWEjZL5EvMWVzHOJi4
Z+c6Gk6r0j4F7ilMX5Cycxsfp3qWUQXUAYM0nZfdWZcYY/Hn/4xgheFbkvk63iXZ
WaJOy45RTp6DK0dY6fkgjMvigQganvaCTAxQlkPLC+xzT8kIEl1eagPpJgqrnX+U
gxVeEagpBVjB0l99vHq74/eACPlgQnlCmouqBtknOBR9rC8QaJTg9rP9q9kIwOw1
SkyqJ+VR5Afx3EHEzUNyOiBwKsHwc74tXispmjkf1Mo2h6iECYxm0vFon/lnoLvL
`protect END_PROTECTED
