`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E0JDoNdq6qdIziwCY/MY7xHSgRSnlTHpa9Nn4YCMkvoqWEYSJE/LD12CO8it88FZ
ccSzx7j5LjH7wfmgjPQllnJp8Plydq3d7Fr+IDA5D8zITE1M+ft1LkZ8PNPyeCo9
LZs08DLDH6+Nmkd2NGfnBtppRI6iZrLAgD5hH6hGN1TGchPbQNYy54LGeATSMdzL
kxnYG1GUWnEtdzdj8hDUAyY527miWIjjbjGdq8lVsThDpcgSkzn4T+uu3miAJF41
IJfRSuCq/do4vp6gVSE9LnvXZo4fDzVeV+WHXvrm/Czefkzz7ZpNOEq/Sa/Gpoo/
Xxm1k3Vr+uMtQAwSVAxhdbpNdgzoKqUxij++gx0+ei83ruRvd/YPHvCWR0EgijIh
GqrAenIwiZVoX4ug10XnD8fJf0bLbCyB0/85xOxHzKVd/pmQxU7+gz4/M0QBSQ/p
sHFrN8uzj1Y6lmZ6xWn5bx+ZEXHBltPCjFVYs1ZuXx6P87i0JqhSd1rO2we2kZny
+avyDnfyfoHFCFqaHwIzTRwRoDiQeHeQdjAdJrWF0qM=
`protect END_PROTECTED
