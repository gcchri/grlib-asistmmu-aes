`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jScNsf0yvhjhuPNN8AIgbN9njAKb1WPP6lzKDoN7UVmx9CE1l+8xm4UDd6s5LTA9
lTBPF5edtsJEn9h0e7iis5YypnnCMhZahK+QT5c4XdTu5NJsj/tdc3HZi5UhgmWm
S0BeUcFUGDosUaxb31CR9hoxEh/us/CdoiEMWdhcsOiotqzfxDep6wAyJt5q5exY
3PL9ECfJw+tTm7phvwjgvkrsIo1lAoOcCcg4y5yBUQSj1J+FvY4wdBHeodZyxB8D
Z9SH4jxybTyUIu8NJ5uhYlKamNp3yFfHcuzDgHMkBpghELiPyRE1jeUtTjqYmos1
J2U7jprcgKERd5d/+PN4t0KOOm5i2qO0i/CbvIBNF/2sSVEZ3/rM+2ognC/YMQy8
efIvnHo4ycs7jRj2zwJtSA==
`protect END_PROTECTED
