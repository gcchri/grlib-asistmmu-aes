`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YsibU3znzVHFPEwh1mfgR1dUZixD8YRMfSUEcNOCOCsCYW9tdP1CRnylE2KTEQpO
FWCkb9y21fkeXU5BCmloJZATtxPSu1OsflC1fyRipnONzRIsoVv7DPJt0Vm/MMP8
TDukf833lxEFmASjvihvu/kCU9Ft3H4pf9EZr5hanTfkzlL1ZefdN0qJLru/h5J6
m2/p7r4PgtWeRZpPUyun9wOqx4ypBAvTulT6yCu3HZnCwVcFAW9EOzOB6qRbbM3y
Gcga61hGPOrdnywgss8FtJ0ci4qn5sVX0ZzlfN2fC8Wtuu3+uOo+EeZfxLvrb3d+
OMWxIo/8VCM6JEiONfEJ2g==
`protect END_PROTECTED
