`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fLF60hHraaSFOuoRE0ZlEOPF9RM3Yrmb+PCirI0LtHeTp0v+b5iCuiFFZE6deiPx
Eu7gYZ76KUpNsblN9UGHrzrjNkrnsgHC+96/p/7yAPXf8jZO9A2fd1buV1YdLf/A
CN8tnLRWwxG6dZDi2cx95kpbHtO1ZlVB4R3mEfWBUUcGlHwFciMVYWR4t3JB289W
eQdrVTK/fZ+B+2H6u9BxR9ziaSUKQktoI4jqRzfDHDMbCfFqZPbVfoaHjctyKw7f
dcEB+dj2NcGCUX3WzpB45gOf3s1zVI7zeHi92IR/e1HuzJw5LtljvBGKUrtmwIfp
vzmXlD0OUOZbfIOdqW70thvIOcmjmepFVtWSaqyFsfSP9TxE1p67hVRLO38GwPRH
2bMBYIMMv3IcGSNlrhM3nkENzAXxWZuau2nx6Eus0OiAxanQ5vGgVIOaJAlIzjZ9
nYRpEc3aZoPKhNGrkdJri9nkcf1PUo+F97DjJzlUcwAHUtBhS/7kJ2xkXvOTTYKy
xtvKn1h/VjF8tAVbBzGzXMF6zIkIV1p55MN+hoTPloOc04Rc4S36DlFi0rp3Uqa2
p9hXKueAUpxCg6GCXFtY2Tl19f3fTwFJ3G8vFrgNpV8chvjcv/vOX8Pi66gRMe7a
Kh3j8fD50DZr4SmsOGYl/O0cS4Oqofg0kxhK9UwhcER/Fnjq9Xw8o2CiXP2H8K4K
AG01oULg5CsJfLfj4A5/FVva8aFcKUAhziUNvVAGoGCOQoQ+Utj0T/ezKQnvrQqZ
3Ij7rg/Tt1Xew8mm3u28H/P+9hjd6wsgvUavRduT5CJObGO5gBX50LELMEPJjuN9
/aYL+iOgdosO1jg3TZ0rw8OFcbopUqLoTcWeX/17lhhu0S9O+wPiHrhi9BS+kII5
sqRmEihE3n/GJ+CwJjggDS+pMKyR0wHqxJGo2kbkUjg6TpOsy9NUAAO29Xtm7Gta
LvfcTtNaIu1sY3nWdZwo3w==
`protect END_PROTECTED
