`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hHSTf+MY7VJkKS3ViqiWMBU0x6QjiKZCZW82e3IeBRBhjcKsPCVC62DB/7ul+EEV
NInFe2LYgkWX58lbPVrK2OmOMzsXTrWIYhrokEMIF9Jpuyvb4pLGYL1bQsB5rJrc
MPVaZxi+AFuosVmroRoC0PG5MQ68rXWVbemn4LrB8zv2/MtHSVzyWiv/wdWdM2SC
BCcA7lwvhIvd5szS03PyOqdbLzE3oi8ToxdXIYke/xxEYl2+p5zTtpBqityiWaJl
iZHDKTCPFHQcwk6FOPoPo7+n0BapQTwk119KvMs65iL62rWFLyhl0lUzTowyJfxT
4tA/6lahLn5l79NWU+zEeBxggNQg5tnH2wHFBfAwmcj2aVQYJsnIAz7wzsq2evyO
VFiGQ95fpdqfBmPpJcb1FyxZTV2GSBwO3EqTpM3Y7RlDWV61MaNLsEYfpRxFf9kV
Mq5AzxTMdCwrG44W/SLLzwo0LPfDjQ+4n7t5DRuwPx8J16CKb6OFuh6pgUWuGsoc
QvonWmJ6vs73tZLEBDJyzZD35HeIkHZ8x1BKK8rAZRkO+le9vRylp/yD2+yE5Oba
TFnHfqh/njKX5YlQGcyC2v/DpiZMh+hxgCrNka6ieSdOD1z3FA3qsNnSX3+O4pZ3
ZIG3YDsyWY76vurtDyLTzWBbPTYJvZmMJFJiY9HDZvh1twJ+9aIid6Z0AMTzfBti
2F5NCsMI3zuG2SCZvFupmnWrrac6TbQALwvcMkQARCiMupYESb5hzIq1wtnHvbnZ
fpG4tYYoCedAiHGKYKfAeBGCvOnG+jVm5aHAdSYt/ZhMtGunBwI2btF26tAsP47W
wmYX1WFAhBBTwZkEfXeP2FN2ZLuGYlnRgo6MJ5d3XS/3VI/HkrgxhvN01EEUAdMP
6ZA2V4o/cPhbdw7bXSotEPusaOEdPvVj6IFiiJ4w84oMgCnUVPcoaDE+6YI/6DWd
xtcn/imfa6SBi5Sdfib1U51xABOqi+Kx6hSSQWo2ciO4/PYuIrYS4dr0zxGvqoyP
oKHJ3XNDqocIHvbR9+PHiamjSFaQf527Pcazw4gU1Jgo/LU8S+heAPeM1iPlcXH/
vcyLX98IS9lkfufi+G7OblhsIgAJXmtvaYB7UdoL7vbcAeWxPPFTlt9FudbZ50FJ
53pnVQzko/KH3wh+qF+ZxbSBvikNbhh2pG/TZCcdJOoT0UV8B85y7uWQIW2umTzL
aafa1Z2oirsd0GvYjKx3a4HhWEEaXzLLHGgrg1o2KW3io6fH+JK+xcEDUziPFAk2
IJRUNul6+dd5v9GtUUIvA6fmfjhorckud7uz1yVBNrXh2ZVBwu+IxtME7THi8zse
LWXajT5oSZkQtZfQ67DSklbDkP9bupwg8ceu1bYLG8Ok5yA1e75aeOEKtJPpLidh
AydSVus1DTaZp3TCaDtLa4A3MYM30Lj0AbokRD9cZCTbKTUitbHFJ2qhFNFWYqNx
14Dxy/QWkqzkXDTl1hkuH0mvNA1bw591qK6v9jBHzy0DoWpCQKQm9C3Kjp42xRIB
nHG5bwKUjbfHbfZS6ZUzE/r4BG9VmSxeFF1CuJDV0i/jigTSDJjZ4TckMMEjQJYt
QFa36ZcsqYMVvncqiOGLpBaJHnNotXlwwhbmpJ0scA0BXjzjMzL7vvOpgnw0buc6
uewJFp40Xmkd9/YHIKzLB3FHX0W9V/x7Ul9/H8+ObDh46FSkU/U1JnlD9A7kPQhT
xsD9L4RdjxX8ozV6v4FhBHbGvWEz55UD4ZROvaNw4tVcKJFh4DViLE8wQQIyuoJl
AzfFTlNGdAENhqr7Z/8PFSIGdA4CTRDDf5hnFga/0eP/jcSZWb4Z2/1yJk6N67y2
tnr9iHHaHyNDHpi3gyca5+pRtPsQtzMn1fmKr5kqE9QycF0SPQiJl6FNH/TXMbIz
Cgt3J6z1D9znwFGA+At66w7C5S4ljbn02ndi1iPMcY9aHizhN2x/EItz+AguDEq8
L26GWVGn8T7pplEfDYwUfX2a3mT/MwWpJ4XpGKb4p+XfVFHepFHcE8b7y0H/SHc1
41rCavQ0xujwp3P9wvu4wwca7SHnJjfHZ/Ss23cIpGtH3iTRqj/hzrPrvC+8Vwsb
k5CJP2LeZMZ6fXy8+1ZIN7/954VbkUjZu6RJQRX5pv2CwFGOCGWmS+1Ebqr18mqy
1oYIqsraEt5H9iqIxU77hA7K/Egk8EA66MqHP86T+2IoTJwwfBGl/Ve1O20sE9Ru
c4/WFsztNcEnfafINkG9wqZK0l5zAlcYcrNMQQk3GG+1+E7Ny6IOOwAN6XQZ/kjy
jYwqk/UxH3LXybpOC55loGrwkE9ivPmq7TIT8Hqjj0c=
`protect END_PROTECTED
