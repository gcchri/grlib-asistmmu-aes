`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n49302tebtNEmQYrDbIpRqjAkU+6Cox3EMGGOKR+jTrIJMjufL6VrUTnnZDDAL0o
ckGfAhyS4vvkW+CJNaAAkwt7ywrwCReG5UaWfH5RP0RAgz2Wq2wU3FG3s8HRFwGB
ueJtN/1oNIsydsJxDE356/g7NNH4DA4zWGOg14BQDGN/rWJQxL899O1ZbcqrBOoh
y6PC2IiOFRceUcSqOc81P1B2dafbg5Rn3u6u/8sgCYLY+0/F1unMzPkZOrdqxj5u
eRYpgFnI/D00IYKYdeBTR6iUeBAk4Nd7ysZZMm/+zujmWMEFVQuID6SrQJxmKSm8
LXKzrONYZGTUEj37mevRDKTU+hk+UaYQhTeAEgYaC2fR9DlR/dUgP1Cxj9gZohwU
mEwXNWR6QB/yFdNQDnbXVJPPWitA3VXt8PGWnAuy/c4NtOdXHabGSNB1XZ7bCbP9
PhyjCwTROet++9nFzM2O/CzlZ5uNOxsafv+sfNmB3Mqtylm/avDKuj+hawBubZ62
rOiQ0s053Rd4X5PUw1DG0KyXBk0ucEkt94413wfQPJ9H+svZnIktzpKRVJNVFKgH
9/5NXgSFISfgx8naIKSdrHOrnA35kKAYcFHeYspVYwbRxZZ25/s4jzEzWcI+Gw2R
JQNrcXa/BOwJEap9vc6IPjbNF9iUH4md/Yf0m/9t2AFqNNTr0fXQZMRqhbMTyE5D
i53rBBDZ3d2V5VD47YgKd9ytArRKnIpM+thdC0Q5EESQp+bbb2USfmUjDWOrh2cH
2wn0uX7HZjU2ZaAe+RVCZSb49X/4UXiS6U6dc99jygR34EeEyZ8i6BwyFTifCuU9
LBDDQZ73MTTq4hWHPHETRppCJKfN8VjAxGDknid/niwVuVbCPOxgngunaoiZVdXv
ApKsFKLueWAI3r1bGL0x29+WhNcniuCieSu51pdmb1k0HswMg5q4A5JECui1rhMU
cQgJlQqct4wWywzL8n+nAy6wJyg11w28CmswEnTc5BLCWlSxpoSSm4t+LkT1AhZ3
Wix+WzUJweviwhvC5yCTI1bM5MabKGwi9ww1ihC/fbZAG57Yr5sGLhBSvI/DvnKO
wlV/ewl40ykzuMY6A97+avFzYy5m1qE7T+63JhjrK37CMEIsywI02b0ve3Uy7ZAa
8aU5+1+mVqwXy3e2pd+V908AB+9KGXfHbdyr9cgoZC+b51rrrkrLngNtvFTAkFKY
sD/GntyY0UdZsexu70H8WE0JjVC+YJJRnqVJtEnzrU5yPUFcDB7imxO5zTm5Yqjb
DVBhwKUEIaw0P0tzLuDIUoPk6uQTv1c7C6ykeUTIrP4EHdFcqTGO4Yp4BOdmlMfw
ikvUmj977/aSwzHN97Rav49U2tDMS7t9rFIiK70TiAI0l0a4vdA7ZPcnZxxwOLxZ
7iw6Hj+lQ8goEKtuitGPM0j9mz8jfA1BO4UAg2Rww39qk/Ol4beS6Zgs9R2v+CdY
93e4uT8F55/fx7fsTu984nsqQQDysFt2cDxyTt92woosCot8PGJLqqka0bGaq2PV
8elfvbJDmf7dDXW0fs5Y7kmFW1POwVa9MAQALsLmqtvBV2uj2dAA3qDVVDODKfWP
+9XaziAaLPWOEkIfquOKoWPbBLBcSvh4xr+FHiHoR/mUZ4Dwtu3FwiYrqFW67fmB
brrIRdEf41G61nXqDVw4fTHJYc+aqC0ex7qTbRoRQVp2aq0mlM/ROuSQ6gTZ8I0Y
/8suwY8x8iUMlZmXxHX2BZebboJGBE0OekxrpY0XgT8YYaumr8KM+K5sKim3IoD6
nnEqCRI1t814nRBntdaYbyo2deMCknbDZa5EN+FrVmyAqzmgdNDOMPlnvFw+f5a2
JYyo/nivnOIiKlZmp4tMzA3HFKNHrnB9FwBrGME8uYSxdiFNCvLKtMtJsbAJ8fu5
2EyFcPD28CxBoOci195XryCJ0WFbCDU6XEzv/cnMJyfpyRWW4KG8y03N8Ns7j9ke
PjCHE3/39FNaxE23+y+fsL2OaqDHpR8n//cUIqAe2ZHXdAZBjiG7H55sa6ejiNrU
HYV4tgZbI2BIsvat2U2hXi4wCmCbeXHT4ywPJr0Mda2oh+XCHWzebawbWnCV0QkW
AlJL31XHYrfIbeAKpp12f8Vi1hI2jMKdZyTPi4yflZ7zKlatfE78vRD5bd+39BHJ
/21btKa4PIZ/z/e+moJlW5QiZjVWqVZk6c9A3wyZem3wiPoPsiUIWIorN1decl4J
DYZNhmDC1USEF5vFO/UKeAbOlXLNFtOES+3OXluYTMP5cTiQt2L5yqlEkrJ0P9T2
rdRvsMN0HdCmLF7SWBEKQNCofaI1MuVyY93oCsgWYzY8MKwfjEx9/K3oE0zHmLuk
fHjfCplx4bh2SMtUP4aPJgqDJ1kdzo4xyDU66RdWtX/Fy/PL80CtLTWsMkUnmA4c
1ofk9fbH8DwIl40AQSKQ2X0EwhOxKOiLB71NrSmYWq89nF8L/MLSobRFz8Ruh2JL
aE6nMzFGAbmUTfV68rgMa5QaE0k5rt7w2aDmOJuaaOADRb2dp2e09DsMZc0Ivlvq
4M3aLw3orBilsu7XpVwybVQilcxTMbCauYCPn1Zgn36gcUtsfM7BF2bU3QK5ZYx0
4p8dWOWKlMtOwIorq5gglDtTCejD8LymPbmWEpEQNjcnOxaOd5xhMyJE4pJBmxOe
k0wnptcRcu3Z3DK5iTmrGz+hYYPyGjF32BOmvZzAzb7Zt/AP6HkTG7BQm60dhNHp
OSin7L8gKSILXHophByOE01ASBsGeHlCe4dn9aODqFKHEs9bHzJlj97vK2NoxEoU
zPywHH+AK9yctQMs3oJJEZGWxnf4GldC84D3UwjFcnpf0LpnlFaNlRZ0gZUmVP5x
+a21ooPy49rQLlIKPyQuyRdK4oiPRGhoF1byxGM8aQg/ie37AlkiwNYD8hDzaOkU
yxTp/3XFhUR3A0ZnN4j2t/lr9bN/GlDhgpmMoIe/h7z0ASqE7BA5VEV/WETxD95v
hFbzSxSkBUvd/naRzxgiC1jvbtJVessVSahrNEpDaXWHQru0HAuCPUg6ZweLTZ8c
u5G+sQZxREUOadrEYkSu8k5APma9FGTeYcG50d3QM0z4QLSKo025pHUubTBDtX5l
6mjO7KMljP+mxtAsFsYz3rjcWaSlaai+j2gy1CuOlNxs4QCT9xn0mIKzXZG/zCXe
Q+qfAnq/0bzuM9u7h2Ib+o625VL5IDAvIDvSFzwIvMQBU0RoWyw/5arOCcH9JH6t
EUmSFEvyioXA8+9txKC/fgpPpVUM0YgzxBv8kbQ1fpA7+V1vg3m4lTHbj6O7XA8p
y7EpD6LeK7x8nwp9FY3eKE1+3aOf3XYyn69qNdKt2qLQDSiPp5NfiR7N8/DXgJVK
Po+J+P6A6+94eWTj64gmQqdNYJlzBS9mO4BHmtpLqCXhtmuMmOkUUbOwWh6UicS4
E0jd8mZ+EeJ3lx4B/1HEeQtCbEUPGy6Y6U9Xcl9rK6lof2E8a6QCEDnpsXgTscgj
l1y4+9TADMOlBiLt+0I1j1MOh6UO0p0SRBWnZR5gk10MarXYeGqOBMWvgNQlhGTX
5ZmBRxMVjA42skjyv2riDo4uY4pnvc45wPSGPVaBK1bd8LVdR0iWBEGYMN9cnPiz
aWZRHpbi5BF18HJZQJvjXuR9Y7g5i6D0jtBEiCyFGoTfafWRYsvFHwyPLsjIe2fL
w5+dtholliUVakXYuUBeMcYdETUvxspM0+IxCEfG8CYbeWEzg/4Ns/aizuwgQFHP
3U+a46YgkJd4aphX1qzUorJ1Z86Jiw6T4jMep38burNITkAjJdYle9X1KTjjBSlW
YDeAfXESkH/BqMz7bz7dWkGPmSJtH0v4LqgmvyrsI4DpxeI3eE2qx8yHcu84WzSy
ux1MMb3jZTP6VVqeEx99MJemOUYHa77yt+ajv98MlOy+ne4SA2nfPVLkoj2S7+BY
KlBYlHa0O+URRtEydjyAfMRDhE8U56fFWTs//W88ri9Bt+zeXOuSMAz83bEMuFpW
umkZaYOOn0VsWog8IVnKHQNZ5q/WiaX4LuXtTmZgwEdV0OT3XyQujgw9Rd+uq5Oz
62fOx9OvMsU5L8RaizGkAoKheMJqvlC+7VaEjAEzb1tIQx60q6Udh6JrIrpR7gyX
Bgdg2XJN7720R+0CgeaTxCealxaPhR8EOW58uMXCRtULU1KsvYLZRzOUKGvTVuO+
COmMmLhs3E9NcodQJCC+0rM8up78jt3s8zhN/NcHaV5i/UVbIewPRGjuDLQocO4a
kpqD0rDuCFf0XOoLqzkmJK/Jojvm4KQYpGUfkzvaOembTS/RvAeDOqrGx3F+T3Kx
ITen0H8VRQ660VNc/kOL5cz5iRmVDchyv/JsjuQln6yfqATaIoBQplUyTsbat22e
evsLU80y4ELPwgeLsUB+InVWmz1F4zU1K4C5vYhoUihGLu2J3v62KsWnjpIMduVm
GPzxgKI3NBtLr0gABOUAlUSp0/IEexr8qrzBUsYhGVgDzdCkYfEV8DpOBv2bQw17
7TSpDuRCKMC/TvsHzD7b0YJyzjUXwtoAyFfkDez8sYOIGBR2mCkeES9x0zkRL7UR
wTpXX+tYaMi8HJR1BKBQQfiWK/ScY5gSQ40hBSoxAjkkzrUbWj33AhNSEVyqSSVB
joMSQGQXDZ6ZyvWdXUf+cLN63xwMhD3dhjcSEy9ZJUV6SZvRPs8fugWEm+tCTZbS
JQTyprnPmI8ttnjtPwmnNoeFn4psQFs9IBPkYPWUjjQqphKxkSSIlb4KbSO2ATLA
W8GSJHOJlKKT4cLymKdEFzSGhWNNFsh/zS0tOUokR43/Aa8ooj1AND7k/XnvuuTX
tf23BWlRWV8BFzg57tdI80SI/ppkvf0bJv3hn3IRuzpf10BKRdw0m1n0/0c4lFb0
N9lnF8P17jjxHJ/+Kjqs3jGpaUBnExO/8LsF7Mb3ug0jKcakX9VHKG55cQpBB8jM
344LD2E7h+IfCZr2Tj/i5iimUDW4pjrFR0r8HFpcI4h7jlqasPFncF1vNysTA0mh
Qq9oT3SucixeZopckyp1TT0CDBA/Ia0MpzWKxbyySKdFyIMl9HtkbUxiJcw82N1t
3FkP0tXXP1u4PsI47A7jQ3j4nNtm6XruGJctwKvbz1e0GU72CrHgrN4f+BTEDHba
9yd0qViaWV1UBg125W+I2ZLvSSOqlSOYAfMFEVmF98tN9ySLjDkmToI6nktLrp0H
dPLuYtRT0AekzyeUVuBpcqhA+Ua9VctB1qYxm0luMCIc1ND0DUPgXJONZeZQ402Z
5bbgfDhfTXYxcsNPD8tdKRtGNl45d6PL9ajXhWED0oBbLrTXDNqAZaigTM35sc5U
VxVEvspv/pKSU5v6sv94q882VrIatqomzNmzEE+9goH1F2blvxoVvkXqjJCee2Wz
KEAggjR9ebt/xZWZNRGECygv8cqkLNAAJDCK5MZ8v4IUDqjhPTCzbhsB/qg7ZlGk
WbSAEVsuRrQtOpwuCcjogp6hVm/7BawNXqoGE7KXO8Attqg0KsMVtllvS6c2VjGT
Gze1v4xs6T5RYuNbTqiutVFMHibpwkFiFFBao8Awzy2wJKTi2iZ4TBuRY1ZUfpoS
kY1FS4YvUxnxla/r00pBbZcJQkeL5YKZ5ah0Y+sWT8L0r/JC/0eN1LKmV5uQ3jEx
z/TqMHO+w1KMdUE5LfJBhEIAu2sJK9EcFZh2fzxNx8ImK55WbWBNllHOTlz75CQ1
+s0g58BqHJia6ip25iqUYRzbuOIpkr4ZZ1KdDsdr+WQmvvkRvDbzkFYnZxJOqYrd
uyqOvulLTWC19BCr1QJqJ1cejtmf194Ddgl7YZOSorKd3maYR2/ahrBaxFv4TYpe
JWrHqJT57WdJVJ013aXujIXFAprYaMygrLXf85H/KioNH4au+wl0oZcT7dOsHZkx
EylWNxRPpZuA/0+zxr5azznw1oKWUtjLUOZptQoyCl6m4BaGZOcDkR5l6FuAWcWf
5T2Zisf+x9Zqmgm3V6T5bm5SkYzYelqv2TScJ+urf/QRqTv7u59XjnLVBUxAVYtH
PjgnqzLFOHTAZf9BPrIqljnh6V0K1lz0NOh7dh4D/SnpyY+jty61HFo0bNPH1W9N
dzjoaQoxSwWn2ukg7YtZViqlMD6dokwCkQ4A4i8E0S4YNsu8Iotb/bPPcGA7roEB
0l2u9SJS9UkzvEuB3lx7huXWCzGzsTq0yXfklK89yUBpGjycrYfewAoVBIpoBVO1
a0QLPyP6ayQN0Zj4KvVE4dbu567CtdQHsTgTJ7xyzwlSK2h67mHUxCUWFM+1GDvx
vbdhO7PJ3kgFPDK00T6e07mpDmQl55+BNtbOM5KR5R6FkAAba8WZ19yxBwG1hq3X
ppWnGiwIcgYnSzF7SlfjsV+6Tfes1GGMIm8ss4zB786VW+0RIG817KB/tPZ0ibP7
cdSsAcok2wC67egcLGV1DlQtOLbMmAYNOGmLbSN9Vw+3Y7f9tkK+hJt5OddESRLm
mMG7Y3l4KrHXziF9TcW5AIehVTkv6bpyh/spXui6el3fq9cbDCxWlegPKQ6bmDbM
Or1BjGfsfVfB18WAgUciVNhIKYt3CHesj2ex7fQm2UdLGBGSvCHPZLI0fl94Nci/
XdjC2rdNPOHTb4nMIbuwTrtvCTmAivpdy/f5ugthFH/0LlPSfH6WpKF1+ZPlCD5U
cYwqkghb9YF8DE8idUV4we8ewZOWJ6Jo5YQjh55GoEHYD6WDgDoox9dwp4k2j3CM
XrC3/KjB7EyX3MlMK/Hd69nAu1m0u2K8wA95w7bqAb4RmcrH+8zOMWx65E8s82Eh
6tJyt9/Sydv8Eru5kTsD168K0uaDleDhgvD7CA1/KUEM9nzsKWiJNYIhTyj2AIzd
/S4SR2oDgk1Wf4QyGsGYEV+ytQTEXRQOK7kOFH1ZDCB9eHsIedEYoO6jfieIF2Sn
KuG5A1XKYz2CxYHU+OSDJ/JNYoKQydFq2JpNlK0+gjmoHLcvoiDTAOX1fOxuIcKz
gdGqPPwcBAzXm6OTppnC2uoOjwinYpvFVFgdnlMsARY9L9I03EfK/TCK5zOj7P3V
MStcKwCmDDl+RB6N6ZVZoCPtKKOPx/Ac98GmJsxOZiTEvNJ7OkVw3Z9XxZX6Z+b+
ynVw8SftibPLAEO/lPt9cOy0V+WcwDvYcCbVclG/JFuWv7Jr71t8gXoRRuwouDhk
+zLuThVUmnvw00Pl6bVhMtD6axeYm8OiRYX6m21ESjcmjOj3AxpQH8U4GR5p2zc8
n++BaRof3RT3QpOOYXIt39Q4NFnXSlphC+rxMrbR5ugTG3Cc+w24M3ajE6K3jtGF
9SkwUECyKVgh7GjT2IRPB3YlEi3bmnsNvfqXnMIiIDV6GgpYk8SLV/rTUmeSkEit
8zQD8H9t8OerWwv860jR1zVb/VJuEI87e0X06G45n52aZqKFnZQdnXFFIQNnQOCU
SSyhAsMv2vl17Ov8TyMNZGsT4VaGxD5e3oeVxFf9XN0DAK+/4FcUylXFrMMAKyrl
RcxK84WdxBaLgzAwvFGc2GmSsZTM3qKo0wr2RUIieoaQqt7IjBRbdjL28tpP4Fsa
KP/9GqHCNzwNVBZnecwmgL8fPeCmjupV4+2C3tqOkUra+wOXT6gsHSnVNz7YO4Ya
gsUIJcSx+LoWaBvPfPTJHttLSx7Mk/1W4ZK6roLKkI2YGUYngWHanpEml9xHHnS7
edxM3qgBt9tJXktY5ZWpD7DWmz22EhnBKNYUAIQ+damJvM7UQjXOn65UDL+d8h24
lM/FDk3HcD4WHh0Vljj3hiwG2CXcFCahiAuac/QKRNH98H1iNgKtQ5yiQDVsh7Tm
2Lzn5dMCTcLEW2xI+AJdn6NMfRI1hlYJx8cT4bcSU9f3FoToZem5+0G7nB4F/nkZ
24Au1FiFcP5H+FQm80Kd80BOhprCt2K12ss5LjRzkUhQxlr7i/FSCNxJt/XpYnwU
d7hLtRfsAKREjHRSxjQfLjycHz83PFHNkrgSIgvkvKMOdSldKBXV/0F8s7UppPbn
3C2XDJW2lNUylMgXsaXvpmAt51P6lB/kuuLu8VSgaRO7nDe9zL6tBel/Ah0cG3Se
Ku9gJ1xv84HVyrrtarXfGK701r2B4OasfwT2RowDpdLMAx5NJvLRK528MnmGXefE
E014LaY8hZWK2aC2JYiHEJG9QgCKwB22+Il+K4zj4X6LZKXm9NV/d72u1cDh4qS/
sJeyw/QZ982QfdkE0V4KO4AEkX5c+70a0iqfHrJqWb+JIYRB9gwerCKD27orQ96/
KhraNjlZkrGTfLFJL2PD3IVkC1SJxVasZFV/iTe1Wp2xHgr3P/6c32PZRh21iYHr
0vHTNCaquwkIuHbXBHc+uFrpN+faaNlxVd9v01EC8xs3AZBN1xQ9yB7EqwBOZk3y
vt9FVkHCwvG37tePoBFeBl5FzVKUfcTGerETzRZWYky9nbIFa6j3uyj1CL1RewGS
YThoCc+wf3GKuJblPqBb4xNB4+BUWTlyOujQLEfATs5w6/lg+6OI07VZCS+fwnyG
lccwQXNBJznrf8X2J6pUrNnaaGeyfBPjwNFhs0ldbhRtr96uOKkj5mYZMrbZKgXA
HFZ/OP+n73EUreCoQxkzNftwDUrjyi2HN1KPRN9qA2PsrQYCXw/VXTfcNK6/vZAs
99ZaBAFjuXNUViHqoR+w/odRs5KFYb5rBL0ZWpmInB7n26JzKHEusYWrifkVri8D
BaG7ZoY4oaXaVCLcvN7e63MrRcus6jIbWQg+aYXI0xTsgSddB5Hwcn13o4ABFmpv
diMGElp3L2PlZYdv6YldzCv711zbSAE8NrixHzG/NZ1zgTzlt8aamfb4rRt4vgeM
u5UYegytvTFD9aED64/u2UYHiAifhdE6mb8E3yIkZE6jdr+RmYe9maBC8O80OCZu
xeHxs3YwlxgqDaYz+6S10igK5ZzJkom3t4ZsjngfVASjLR3jYTqx4RueOdKDUC1V
WqKrPFwUcqEjHftXQInZ9c/U6iqW5bEvZSbGvaMx3UbgI8pmLEu7DI4EYMYVklGP
c82p+UZDRXa2GuQXOBqnREjIx83xBuJK1szQAf0zyJEJWT9ryhYfTV1hQUT5gBpZ
7GI0mimBOn+OugBhwuEB8U6LY3eUFOCUXZrEy/aX79bRng+KpgMc5FnHYDlVEmtn
tU3Z0gZNIUdHNrS7c8tn7J2okPh4uN3L3nvQAMLlMyzjXpwQpMv8camzoXLvGnZl
eofz2cXPZM5LeAOntr5ob5Kfx2IjDab7QJbJW8MgPB5a6gwiG7NmyyOntdiplI/z
z096wHLsfzRBXE6x/4Tsn9OQiYbk6pvPw0wc2KrhyaMCt7j+qE8joDp8weiRXD7F
hSiX9hD8bfUoZoRT9V82WEfQ5i+ugL8Fi9o8sb1wNIb/jjaqTpreFWQYqXQUrBCj
m4cp6yiCWULpUDqCbI7YzAJi2sKAUzKRNLutHq2uZ5sH83hja5jd8p5ik1HoteM5
QJqNqgctBo0gfcH1Y4EawujJ7/ZrgRAFjW/pAF7SQ0dedSb09+cEhKwWnW0C0D8i
KN4IbKd60yDMc/C5pLbJ+ukurrvvsZ1Ip9Mr5RYPLWBQp9Neuk3yVOVTvh7tXB2A
SBZ7aNf9zURAl4+KX6l3/a7Q42ro9E0c0JysVD0FctDaGJvjbDmfiy6m9kq9xjGs
Aqt0UyLOwkpKdaePQ+uw/EA0nZtsSbhDFf9W6ursZW6EVLM1Gn2GjUSa9GB2EyyA
R7AzRVFwmUmwbg5f9ZXzlW05ubYdGcCmM3kDFj4abH9dGlzwV9WagG6C7bjyoDNb
eDp+aTE4ZZejVRG8nadeEVPuq3l9N9WL2Cm0SPtCu4ucDz/tM4Zkl/F+mpYOH8P7
nwUF1GpAMZr0/d1nSaq5A5lPL+qmqa2DVzicOCkguBXvjqRK61TIczLB8bc15Yuj
/wKmmfFWkT7sUeiVT4vqPiJC0Ox3Tdn8AY4l9cQ9PHXIyHYmw6I1DMk+Cyyj0zuS
IUNrZPCG90/2JhpLFLS8Vw5yKjfryYcVEXXYkTAeuRGsntqSDm0TAmEfV3TX/qCZ
NM2f8QdBESu7rt+V2xHiSSAvd779Bd+PycwqMW1133vB2p5EIgbw/KdeMnBGeGC1
5z7E7wcQLQkZefrphNlKdDat1KgdNMf6ryfsQtFbkY4DRvEV41t/mRbsAhhOZjaA
WWk5b+/NPZAgv4arFLQ0YqRHKc75JAY4N7C5ckFlofgc7YaoMegg10JOICLFgvWm
HZtJCo91ZPw41D+aruw8COdGFFQBnUOwx7NI6lEyuNa7e9WZ5FSo66dHGZ2jvavo
8pTCzmvQp3UgadmReilIGBz2v+TwRTuC5UwcVSLHvn6f6qWeUQYJaKwt6BgLY+eU
8JATOgaN77CDZiCBM1GUclCRp5QuSHXETUVBwI6gmd+oWmDvjEN7CRlpRT/8lPoy
qor0f4+UykIPcv0hOenXRuPNMUJWVBciMoqllUnjnkQeNU4VCZWS+ZxhlHLynhfh
9CRM0r5owH5asrA+cPq9l6AG7U5xYmTgDR5v2Gb6qbjPiDvTedcT94V4Mrx9Pu7k
zwliQgIXkqGimBcanvoo4sTjG9SEb9eDhYIGj7LDmH0UWsaV1CDJ9nOXnnqCk8jx
GCfKaciAZCBFtM5FjZk5/JDuoWtyLhebrEzrSNpvarCERMfKqdUVyTWPPT0jAeiY
CO7Yjlm9mzKhK1H+dXOVoniAY9/ahSmOeUx8zuuL2H2gFycSn95bs45Eg7iHBSi7
sj/Bx2rgJoxTxsbHIn5louDc4Bc4561QEZSVohfTYBN6fkpztmaQPfrlw70Jvbq/
ajJeL10NfxG1COw+Q5BIktOhbDNhiU89+iACkorbMFtUSsNUfDKzj+GQG0rE9DDA
3Ftto1HOUnMeMfdtfbylqmuM+do23dFCXwTHNJc3QOBtJMPxDl4XNE2aYwn9Lzi/
rCQ5hhKBWCLxyu5yNJEf/odkTYaqIY+iVYuDnyxRip541OASBjVAYQhx0CnwBKOu
Z0Migc0dyJTMsvK20LZ9YaysE1pRTpTMUg+wIlFBEHfCIv6LsXGIh9Aq1PhP0O1T
YxByEqdNJ1ElHkaQKakxSuFMZAH3q916YVsj2L+xT6ZWgun3X90q0vXsxvAHKWz8
mvN+LvPn6D+Pxb2JkcrnVPFipKgwOda60ndMfEOtZf6eMuGTQOQ8DYDnAlxqnq1+
olrcbCRb3XX9lWOmMyIrEQpcslmDcyf8VKtBgrUyFyUg4cV4CB8sxH/x8yXhRnNe
OJeIWTGrdzQL5lvgn1rXlfKb2mW7e44jhTqJL1dumUEawCE8+TuPmqhlwBXc/vcH
WvABu9zaH/29q9PCF/jj1wrmmb+e5yYAuK5vPju9f/cU39A83lX+yjVx5qvi0pSR
pBVzsz/Cn7u0yRWBqTJYGIZWfu8BGXDJ9b3ukgnqdNvzrKPym3YsnHJ/UaYPEyBx
HJg8C3goPndVXxD6HdSSVYz7Ofn0PjDY5++X41L5ueCGKg9S1dXKpOCp5L+8C5IZ
zMVsltyktMX4dOzDtQGgwiHGkdk1v771WBrK8oVj6TRO6APtZcEvl5FLFnbR22eQ
UGTb1kg7j9autM4fPd4pBcUwJF7yw7a+eqqouGtduFOxLpHCCk7eIF4HqlXPbJ3C
qMDBFPlzdaaSfzAVFb3qc/0yi3Ri+rTnIHFgL3A8GBwZDm9tMVQKjCiTDNYvlDhk
MRgHvMj5P7McMLBGlYJSz4P1/0WXYNgkjUtv0fyMXRAN7bCF5pNfbx1PDumogvt3
IjxITg3TRhjuk/gz2Mu/KU+/NRyfmzkgAC46OFPPUsVIWNs5bNJ+nUlkROf2fVT2
GB1mu5YlF+1+h+9wJ103UoeHaKS955NpThhWnUi3g0vzyWXDbteFHZ7Vs2ux5ea3
o0Iz5j9ZNX8OT1HGaPtiPUC5WUMXWNY7d+Q+rqdG0tuGYHAc6QIVVEWFxXv/jQY7
KGdQusTrUYJJIJ0kZ0RvBGqyAm2HWxCWY0k9ZGaJ2Po82wQrmx+6MFagai7gIKhi
RIHB2w4I1D/4eFU75KefKc+1l9F0fRgtn8oVJtGes/5k5QRVBrFDdbjeSAKbclhD
oGGNyah+Kb1rh9btIK+i9FFcKR252A1GbZGIfd7Gdj48YSegZ92d//aZNaHst4qX
777GpDVzg/tisxuu6fas9HlQvG48C2wZdasHQshQm6BlDAt8gecrCPVivmHxd1JN
zpmc9dyKdcTcISk9m7Kw8cEjzQSJKmS4mK1H/ok1+MTR/nt+Zg+hI28ef5Mwc8Cz
bwVZ1wd4T2ODdbB7gjHX0IHgBl0wumIqheqBUru++GImXjOIt7mYMN4MCZbGbSEt
qCBj+BGg8OQWmmPjUJgFOqtzvJBqtYfQx85mHpN6MgnNxpNuoRS2IiqPt7atIRFT
tcfu/8gpmQDeDzgs5lxVfgYuuoDzSfZU/AT191YZ/eAxbC3own08C3L52bJny9qp
K3l/JMCQRyYbUhvqvLF4Xi68tDnQi8TnWJZ2f2Il+5lPydLXi/eua0AxAaOY98qB
Nke41IHq6t18BbRM/ThCLOrPjOgJD2IGsvp7HYvsSvuZhA2DxamJ5Ea2fBDE/XmA
Oq1ess+IBuidV8hwfxaSC7pGmb4OkRi7WTYAhW4rc8+opDDtS7FagjsGG+ihhV56
ukflLBlXb5BP3WO+1Rr4kGW/9mDIl1AarQXtuHKjJHuY29398WQ+RobalRoqkUA1
Te6ogSU0IdwoKlh355+47kjEfany4wWrCb/96SLhRuGgAgIoGR/HnZC1FtaNBGDy
SNaxREioQy9h9LvzwusMvt+yOw6fvO+edIcQkXivJeAkmsRdDfAzeVyRe9hf1kSZ
XkIku40m6KZ1qAyWxFLKDbjzg2OiXyqTnD+PySGkPQAtDPHmhMCGFG6EGT+nQIya
jJgkQtSGjviUFYhPNOSig3E4n/9eHRX/K6b3Te1NUMGYVI4H/BbUD29b/6SCN7C+
lIzqBw/hfz4oulnx1lSgvNoiQpzkUBLooCDxjXdOzOk6o4Yp2MDUsMuBv64wOD50
JIKcWDQ/H3y5o7AFBLZekHslxT16C43/sGEW1Pp5plo58PWc96FzBt6Kwtp6UwBA
Hew5njEOmuZMFcNhosAC8BA6335+HP6lzYIWb/K6Z+PUUrqW4CRZ847Ts3BxePNW
zxWXBZkTsisuYFDu17YWB+CcW+3ehPOAUucxtuOfwcl3l13ixD/NHnhQVk9zjnwS
au7GanQlcc8bi1Pp7M+CVhIWJ2ehAjpmZcjSK5C6mPi68kyDODRrNKjDMdwAB4e6
CIVEQEAneTYsn1E+8njAKinvMhfreOGw+3WartQwhYNLScgMhpcuUoc0j9IjnQo8
qxkQAHmEJvxU2N9qj/p602MrODlLfWghfR19VA+G7NLzVmkd/Y39+72/Pht5sdq/
ZSiBddOF91aT9h2Lym2KoSqOQ0fHsi9GM5TeVjgYbSs0J4ZX3TWPAYOqfk9ed9Hp
eFMMeiu9p2IoIncOe4Tg40JaNamty6kGe4B3U0U3t2XHG5pESky1d9Eo51aisDJC
FXGG+Gf1iLxVmi5BHgVkpopS7c8oGwOCX0P1W5ArEmigAqbWJ7R8EfT0U6jAliaH
lmbv+C60IUuNLRfDEKNx4RRZljQEQc3cX2D0ad3ysYyCHcbGTNrkWIt7jxU3LY8Q
203lgA4PhSWIqV6BTM1IkdLcsc0klT4mxSg0rvhimF4/0V0TdxjYCMgNF/lFPhNk
poS/NZgT6xVdkqqUR3NT7SKNk6gY3jEuMgMTb7BiYw5MVSPlHx+/+DcS8K5y2YHk
ZeSVF0/0vFIlKtvGmMsRRv5okPbDfLsLUMMce5UFhZwnW3+OXdczkXfn4nLikQCx
UEPRTmArWOzNkfdkg71Nx82Oc0cqJh8Uuf+HT1a0BmfZfV/yj/eSDfd0CfGQ35fV
wWTrsIvMDzHwWKdBSQVcZqtW4kFbpwatJgYU7T5uhNQJKnWWKcmwkAGsm40GD4xi
ga+Zx4n+wzViRzj384PzqF0rg0788hR5l4S3403JOh9Vf8R+F2wBxnDvRI7kzDj9
ws/1YAXxuWPYEsEnWUR/ElpN5/s5FXeDaz7c4DVtKkrgWpd4jpwThdasf58fOeDz
uOD+dSPdnf2FV+Q9iJP9VAwrGUnMQBGYtp++KWb0aAEtRW1DtGPLospXBEQlRus/
US3zcSOSz3XekeHAcxkmu4/s2nFLxvX1wDnatGZFeO/aB+ygngffTH5/IDFK6o7z
yHEB7Wa7PMTEHzB+UIHLBYsgpUHRq9udnwUIEub6accW2Fc2PCfT+C0jr7MuhG2i
8eIyAkfGAgt6bVyO/CBJQmrXTtmr3Q9nJAqVKMgvxQXOv4qutLeSEibvn43LEODk
wePVbkRjFMgbL3PyA//kW851iq6bdkCUQRXj3lAg13crGo9KBWhHQMBJhoZv1zPV
kGTMM4OxF9PCEzrv6NyXNagOVokJOSn6B9W4Lt+MmRkdUnI6PPAVPWNDUcUhxCs/
Kpci+lFOhSFnjdefJcdQi0zKHdUzOBlKGxh8N9Yockp1HzQ3J48qIruiQuyo/x7W
whugcIqZJrAf/Z0nW2jz/UVJbjHRe97Oxvk5jigrw6WZNzHTAVox1JcI/I5capY1
px8ACxgOs48O7y6XrJfu0OLdtiyH7+2hBguBCK5rSz+hw7ZYP9xZaXXHGUC+4WM9
N5OiNJA8HezP0lLykInI9lejgNhlIWKGP/78LiXXtSEQbYi34ymrPaiVKIA5J+Ym
ZKKYQ6slYcM6p6r9tr2deWYI+Jfa8yqPDjfqtq9IlJgI1ZLWBgaCrMxQpA+MiUTF
DIkarAUx6U42RbJmLWBvUt/aL2Uf5JnRsErfaxvhVatV0lbvoQeqVg0u8FiMVzhn
610eBR3PkB+0KYgbVp7AnXpi588HBtKu9hn3LS1dWo5cgW843MJLTYiMGzqv7+/B
8HYzRYiHCHCDTH3DB1A8R0i/90zRxl41aQMSHJikgHXSUWP4NlXkvNV9QtZZE5Ch
DRdwBc4yoRAFzaBwasZBK47IV8F/GAl+viBhBMoMdeXisGjUAzmsZgfwkW2iayWb
+/igq/tVxlZUzOuD1HmHWYp4v4tqeCaJSQAlTevnayB8GMLVtJaupbxBnfKnGDHc
W6Z67EY1B7eIW0S3NJIziK22UzHdAZoQ/kUphIkzASeG51vK9eE9CBglQmqy5RY4
Dl4G90MH0fsiERwPWJJH0kKGAKOnydwTygKyulcOOsB+Ydr5Ad5HkuyFGZAl1Ous
UI1PNFeiZxfU6tt66SiUSGKv44o99Lfm/zbWv8aptApf1ASsY6Jzb3tVoXTppC1r
QdsnbfDBkY6Do1WQzgm4crWRfbrxzeAkP2vVHTszXqU5t6T4madfDatpZtd1sugi
aAPcovUz7I3IlIslrYdmGVF9gugqKTuMMeUOxpPXBziLlurDK66rBodtBavCA0tq
ybug/CW86PejPWNXsI2qN6nJA3n/EztQdPiyk1q1BRDIvxjCYpqtcVqJWa2UgMmu
wV9umch4ZyJ1Tj5QCbl96cuSFoXgPAT6KnZCSi/gwC9LXhlXEuyFcqFBc8XRuUDg
Vx5fuA7WEbQbk0oX0lWd2FvvdzxiYl5mVpPTBomAyCnYGQCfhGKxmOjfMgzoyL57
eK+YbIbyUKntLYiSS0Xv6axKyqDM8qZu3RY6kdgCBcRsHn7BhJpfy7C3t6JWrWNy
LFAyXPFWdcWzu29LBYbwlEhudFq6gmoOfkWWevLN3n83P5og+VmPi5t2ZkApDYtn
L7mPdhbquLcQTBVCU99jEj6mgC2vNgS18JOAcMBJcHRIrarVDLOM6J08oOJ3/KHE
09UnXMoWDNsW5pUEac0tALOL7RX+VZPu8fEEKRq7pHbF3+EY9IBWPjE10ALcrXEB
qGsW2c42p1WIQDsR9vqNjYUwyFec44Km6IvKl9W39MXL3a2U+Ww4vQE+yqr+WPsz
OCgWgm3QUHvJ2OfRimHqgwBXAZABa8HKb+QrKLC9+ZBQZFlQ+UYPD0tt14kR1j+6
a9HmVn1Jg83j6hIOOCS9v8tAXAdQtLGgbsJJ9NFZ1RE1V4x1mfV2HM2E21bPguZA
Rpgv2SaZeOHbsKPDlEIasE2QRYcNNc+3fR33hS3VS3GCmI7HOT+vEd6Irj1iUANA
fakfsxu0NUir7RyB5mCiTSz1tRVE1+tIiSkGC9ARJMEYEQXrSNlPBIkrWb/JAR2X
lrzkuyca87hE4cyBr+Ypgc7sB+G72OpbqWk9NtMaVTd/sEiJbTaETHfESkLb3754
eGmUw9zBNUQnBYMHhm0uPBsHr1OsHPcWEvVjrgQYAu99eTgzVgVFGft2E8qfZqKY
1yuXYIlrPVoG+uT02qARfO6HFsHnXvUw2LD/12W1b90E7ucMo/V6B3MIN2asXSac
wbrzOTHVNaPt46W3/hmnkpl5nUpjNNR5GyW9YNg6Kq2mIMYpqQZIRbL035Ju5NuG
JCT2+T0L8BEHjZDevbxWqejVfoR48wMPjG1FR2A+gDk8lv2r4PAdWzJJfHVSCe/P
fdNjWByMWe0C9utQJlbWttpi/9U9elg68Tu3M/4VrQfifXHsHvjIGLAWo666S5WV
cA6hZvNOcx2EfsgbhT7SsrRaSUHkmCN9EXA4RmyECxWyjUUGbxKdB3Er5LvyAIiJ
Z9NwJ5jq/NgKZmoVxaV/jaB/Q4+xBDkjfbp4wd1nY2P2VQfYAntJMkvHn5q/s6rW
1M43MVTb5hShr+s0cjksVUV3VmLEz/EIIlpsB/aytlEX8zfFyLnPubbkKOddb/TG
aHD8+gz/aNVn5Wcnlfsetl7jKjNU8RaKN8peYpI5avXIRnUvO3TpiJvQEZZYQdFu
pZ6ET4vV3A1MmI5FYl1wTaOeJQIKk5LStDEE3FMbICkVCtwxbPpo5C+TW9czlp1/
QMengKdOjWHqxX4q1G7i+bB2fShPnUmArdCHSv2w2/uBXFYT8UfDmdpfE4YDJKv3
tt9KFT/QCgULh1dUg+rKexKZ7U0SkNpCCkU8ZjooTBFjfiwMQbNTljXacVJa5PF3
g2WnROTU/NA7DrzWsWzFXjbw8qRo9NrvtZcGO2tgQyf1yYfjNzPVUTaU4VFK6LMj
FtMytTi84d8ZnmU71Ng9tFTjFcYXVBNYPtwcpYzCOep7WC8w/GNQcn1YIlqtgPjz
JdIEsCpFG9xScnF/8yX4qV9QZjHXfZ7p+mj+/bcdYFoYEWUl87G4qhCspY8mJ2Ln
VfVTcLM6cjERnz/U1Le7JtATjJsoWqIsaFIRBjLc2XVuUB4ho2lWHj8SSrjptqX2
xo4ZBkIldw79TB9pYmst8vsKAAfz+18Ui6u0pcHSf+Y6D6WiQfUYVY9abN6zkFeO
qPfilLdYiVwxiRQzTek4iLmWDmGYtGVozGjbI0JOvwz/c0tiKhZKUSJykUYDrWU9
dUA4e5MpXQzTe039x2zG6vN2aUM5idT3tlsHDz/Le4WHgSmvXpIOAWvs7neqa9dL
lhNpk6D5SZC8xFeUPKRvdPbH/PGiupH2sdhShyT2pfD/ssDQe3EjmOH3EAz12kBw
G4QeaSQZcIScIs380an11SltOcC+rhdx1tAQBBQwn61xHcyrVyeQ397vb93gclRh
wLCi6QH43yIr6s0vtSKVTG5pArZBEDWWTDEBN/kWKNocrRG/R3++FJQkB5z4DH7u
P0Hk0WhuNHcrcpugbs8ZIAfseSdP1qYVja1pN2wC3ztGE1iimVDMCj65aj6uGy3P
YKXXRVxa0ScNsVR5rs4NAIlVJZ35S0RxOU5JZz94cjfn8sP/W78H2aiKYOS2ncQJ
snN/xjFky1UYVU4FFH+hBjj5qEKGFVKqedgNaDJF7tbwOcYOc7gC66niemPzh6Qc
tc/EKyiZqeq6uO2lHwxuvwQub5HxyRD7jbD4Nt0Y+9bO97D8YG8ZDKUy5V49V4c3
AHImiOufsYbi4fTPaloX6vW1M3Sn3oZxiWfq2cE37IfW80aL8W9SjhY5iVRIEWrG
mUTSHnEB17hhT1Q2oci39JLrpFMnQ580pm0SzU4MJUvGGw/7u3PAvm3jYhsh6cs/
OEySsXuN5r1GsdRDI6MX0x/sMadZ6nvxZvGfCY0P9pn0YwSJAzVdcgb88VYCik5n
hbjMejx0ssTDo4B8CjDBQkomwiktEJT+oS/i3rHt1WOzW3ybEU8tZ8IgxoXrS+l8
EdJ8M+ot8g0BeqX6i146KwdIvLDjlRkAj5NtjOkijGg2PPTlyIkuu8mmAtoxhW37
Vgj43Vb3Mq8vgj8S6hphxglay/YD6bJ4oPlT6vXYo7WCdFDOwIMlmmAwBadSsljc
kiDv/QyNSnWrDMGyG8uyMJVytSeSlr5HLhf8yzBqsMTUpIicPslhhsfTkrPKMC3V
YbIFJPfLi/n/rORsbtWnnoPp81hu9I4NsTwZoTLxTvW7HBogDI3dXNGmkM0DwzzS
7oI9D3sCVKATSVdDZKFAonza026KvfpbjfGTepwIY0BxSyXWe2dU3v8G04B8NWnb
fkjjaT+Hp9ogLRUv8Z1doqEUv4OBbgncj2wwIrA9/hJo0MinN1/lMlSoA9J1TCL6
FGHcIbRl6S6snmvOs0jAlTzGwiYKOIcpxTq5qyiS0zQDTU4d9deLabLMmKBs5O2u
XjZNK7amGJ7WKtG0ZiKeeqoE+MOJH+GBovDE7SkKWw03cO18TYKJuwvDSzsPTI2V
TSd+QAY25Ed+JJSo1tsfRsGbdA3u/NIjS4O2iRDG3SFcQ2ohVeqsmgQ3INtNcCa5
/LYqUW644zXmEMGjQl1fErFVZBrSekVUeWInPZrT73leoGihzT9wK3/ctj5HRDVE
GZfYpMQw5++MYRRAoZ2QPY0kYCHHT3gY9RHz/x/1CZGWKwEk+RUTP5xh4VULeO/9
Zgwr6mVUCO5wsx4NuZoLgxU5xTprqoS0BY90VKaTd9b4cV13vKf8AJNsunJCq3de
YeDVRDfJOco+21ewv//TdCb6Ev4b1CtVmc2Huq5bFvVjVELFvo1IYAm9z4Fpmek/
2HjpR+NX8YRFf0bLTvJ4kr78EF6tVK5c9QLCpJf2oQY6ZLutwPP3d3oNl78JAwAD
6r1ahVTtLjqEgQUI+ukyy2oZscGLe4HWEIhZHhqZn5VBze3tyJIXrVm+XU2aLFJq
XeGRX1znIL3N9cmPb2wbe8dxNVvqozvio02apdhwL2Bd8uCYO7HZxREekxTyVKNU
us/bdLqMRJ5jDWkopeUUqV51aCzoKESl5MdawkT6+HP3hT9UmNq0Ze/uXH/06hNf
+vfxdhz8oyg2q8077s55kvZ99GU3xTWo7/GjKy58BkwxyUdX8XX7FCDygNlJOFfR
9M4kP4hrro37wJYLbpm2fQ/4perwroiIsI0lAsaMK6I7FE4r2pfK0kehPgeL6EYL
DEqX/abSnJbODbHOavgScMCPJ6XhBmn4076TIoE76hZ/5b2qRLZglRpSOQXP88aW
EOes0nncSIeLZUqhDXISFyo7iIgNlMHFBE6qL4HVsN78hq4bVCsI3xOYB/nE6sow
ZgIanxCTl0ULmwYILTuUAIFFTbeJsUsmXssrRVkdajwvOQ0+Skr2Njw43R+XgKRi
+ed0x/pLRsRFcSFUHkxf/cry6Wn7UlLuk2fA1JjgwyimNelZ8ZgwCN+lLTZhJvpt
RnFyPD7vL/VXaKocGJMhDXtDBXulWfWbP4pVIgzvqM06psPXP6Gb29qHEt2/duCY
y/orACqwRG+z/JIl79OsfAomIfEacczm6VsuzPOVFalb9Kj5tmCFetz516y4rBwF
vfE4C+uKI6RGtiBaBbfJ8HK+l2We8TrKrE/l77PPLyZQNhmtoSOZYGUtqlERzhDX
uro2yGFhYPfdHAyyTpLNAvIRJFwpwrHffdUEasVVKb438PMyeSOnZW6MwzYUL+lu
igfvuwIuXmSG3oTfQlGQpbOMFuDzIH2YgcZO0Vj+HepI9OxE+siey4a2SqLrZ/4y
H3FdqVx2yOkEoxTMTg3MCBav9dzN/9BvFEdqJluC6PKGxpn//AgIHEW6y77NU2Gy
HEvbzr7C3XsC+bpvOGG2Z7/Yl0RoLb9xWx4+nR16x5hOuQ4SOaPpqf/f22dWv8nY
R090lly4YmYeMd6QcbU0Ey0hByHQzDtYus+mOIHN0pj4q6R4EAwgSQYaupq+HbS7
2Du435j5gKPF2JHQU0qv6DFxZb+guX+b1jWK4OVcJAW522J8lFB4QPtlYwG+Li/D
SiVEMNZga1dwBY5JEXDD7azv7Vzyd3BlMncAj5F8eOFGHkbJrhAzG5O9JTvt2SwU
fAN5TIbmtZ+wr1LJiQ8pU3NSOnb3GoahjfPCs4a2ToWKPC6O7n+dSzZLXBnp7Ufc
x/jXSb6Xm7so5KZ85/TOFTIIUKM+Y+ATiUqK2dro4Pd9/hmiggV7uKLSwGiYCRKT
snIBm5vzWJc70hDR5oyFllRSlZl6SxuUSQuQy0ET3ZtuqORHff7bUwIsNiwCRCsT
m8VmgCJkbc9wPDvWOMr+OIuT26CNL0yOIAxs9AzGGUdA1pIjXvGdl/IAVYqmGXIp
MTpZ3XPiWSC8etV52cBWO1yXTYf+ha0bcntn2UQ1Qm7RYyykhz8KX/C4pPypRelz
j34dSPW5W21vJOAcFCiBUC+mwOb5YgoZO2BA/jAApc3sZ6VDc/KdH79/7ICEpPih
DMpERXHykhZsjS30/MdXae7Bfi711DuCoK0GY1dVRKj6GprK1woojuqJBiGZni+x
bagEWyxHOXFkTuXPZdOiYwRNRwsWj5VJs5o72VLYQAKCeBEPLcShWCSeszm8aHwA
zxLE2Vepr6o2LqHblp31aDDTe1HTlAVmRdnkOjQonjSTRZkscZNuo6hCp7Wsnr/y
7JNpvv/IMuaAuFjYHaGgMr6kAi2azZC62LCR/7MKAiOpJrb1v37Km+RTmFNRItJt
g1YjQvPdsCSufH1e032HEuogSr+uUKr4aK+Oua9ftnfbY9MRDpcdLGst+ZVlhDxQ
18SkFY+9S3S6zAb5xEx/oQ9HB4oQ/rN3/b0ogQqt4I4x5nYsSC8qRtN07hdsMSed
NEtWB6yPzhMozeR5/Ig9XW6tlmAj/mc0KEJMKArkSLE/6MdvSCvTXriNGexbIBB3
lWy6L7bVa6hdmnDv/Hs5MgM9vHHEGb+INiKjB6yUvZ4qX/CnyIaJQ12laaVGtXVf
ez87EOLH4ypDqddk0XsAq6keeyrMRjHlgit8fszVgDljSEfu+2xr2o6YfmE77SbN
kl+9AX6pwVRSVy1mZHo/4oDA85SBkVr84nei+mL4805rPpzS+6XJqQUUcPhaWT+c
00ShBYbQ4cLtfXl0H73XyB9ssKTSw2BAo7O1y7Tm2/O9u/iRInAP2WMY6xhWrpQw
W2CLuEA//AY+PCoLaCP0N5UMxWEEj794m5fClFQ/WaqXyTzXPW+Orlyh8BB+Hpr3
QLnh06wIjfPWECLWUIFjgyzkudtfahwR+Wx16a72NNB/tmai2sqfENYXzRZul6xB
npHkm9cAD1P9S92ifisJ6TfY/vnVGr0BNC1bbFXrFIVSXPUc2dE4le3N9YinTIXe
5suSaK/0hbSOy3TwI+jshRAKM0UaudHXqgiGYpREeCiOOuGaeZZftT+AQiB+GOSA
j9XZZMbcKKRHyU4LwCyYsHdTAdk83R2+v+jn5RH74JXU3h2C5AxN0UnXkkrVnVGU
U9fPh387ABArBQACQElb1c5ID+PemzztBYepzbttYY4NPgBw7iL83drxp62AXIQ/
4itMSbw6taVf8UsHEO3tRDNDEeb1pCsRmrgkGl1d8PPesZXH/mL3rPRJjaOMqs0d
xUexJISa7HtNDpuWBwudqm14UHHgqKMYPyP+LaYAQzw/trf8BKvV2KJwKwe7z/U1
582OhZfTglACtQkpslYaUscwCLZm0MdoVaCtFIe3/YezA2cOb/cGwwEEhEjfxMuc
sfb3S/+mKDBHZ5sAcHSXTEQkhcJlQrZ6mgBnDJrf5KljZfQYk/qtHPD7HLn6G29D
kVnUCj7a/49JL2c5mNIzOHvy4j32tVIizRpdHemxg0YJmkl+ZwqJCJCUC2MYnNy3
2By4aP0RaAjcuffrtSy1h2MAJMs3LgFOO8Wk7U39SDiLfnA/MO7V2c5SJOf8Ztdo
LYEwB8KBdhJZ8owCDeiDc13Ts8+oI/4v4kVPXH+xA+OWqSRAgH1i5824z1X7KmAD
7MONrJA+tcYL7CVGQLL/RwzoHQFIbH2U9pLaLz0uVZ+E1MT4D5tMcsBwy+g28iZw
Jsa816XlB82vHKzAFawFOnwaojQ5VuIv8gy7dNZ7gWleS09Yan9Ea8HMOJeElvIW
VNnMepzjNk8jlJT5LOtd3QiC189ZqPNwMI4I8NuAyDJlvGiSghlhDFnLnBJQLQU+
bc9Qrxzt2a4HmRShSIrUFMsxSM9jbgyRgyd64SJkf6YUT0AEPH85krJzVVGA7Jim
cNi3CDpTF40v4csRlL334FRI7URKW/x7IL4hMhV+40YgLvL9BuRBgDzVZDK6gLNm
6K3bW3Fl8u6wBAuGv6cgh6em4jq4Sd7J8jvksk4APOEbtjLjkGw7Xs0ZCtz2oH0q
BPXpeXaC6/0AFEBIrIPakPsbtjZeg5MTDOZTQFC4Ew7Xbn39rLymza7JpEVJN5fn
5u1sJoDqHBuYjXUbeH2LZ5q7Cys3n1nYokbH3a3oHebftqkx6w1pirw/O87vqtbn
tvp4IoXaFhiZRLFbSIaoWlVHvXNuCdP1xQP6O7JGMSXhoHHXY1Rel3q2FGsgNMAu
nJ1LXR53HkJhy3OgsnAcimFiusIjQDHjT6dryPd6R4hqmhI/rPqKCXt8W0Am8Z54
IAMepn5jB6R+LhOVsjx8pC4jfWHoKdM4A3MXVmBtddyHxxRPe2/zKybHW2bWT//K
v9CCo6leZdZi0V9zEGAiHcN1Lsq4xMHucH6ydTvd65ADK7bAGcv4gUbfRIxryL6X
j98rQlBIZ+eN6duwxHJK2FKjy+cdpPGD+xV9PDyNBYyqOUv0JSTr757q/0XmiteF
rohWT/b8EcL/I2MPJYGkVpDWfeHAqKoT1nS24ysQBiRSOoi2Jqi3zmPqm79CujlG
Y69aO+AmXSzkhi/SqoX4RfGuOk/onaeJeAPW+qZ/ibzhLfe2b2jTRJ/DBUrICy8x
XkmV6Ba5O2r9ptwH/ABmKX9yOCkEUiS/L9yIzH0DpSu4PrvqZhXiPtXTW4I+A4gP
OpUphg67fV5EwhT6bSmXschYcIigMmWW56bPM0q3zn7HJn25ZiwzUilfwe2wwOsR
7/6zZ1S1ZajyR+4I06lVobL6uvNqqY5NFuDrrkacgInA8HEx7+Ke73ApwTU+1bnj
YDmcWE5Mie728YHFDJUrXLIe9wJSvoeDnLEF+pbs28i3d9dkLiD0YAZsAloIQD/A
MRF7LY3Fc3Ur/CYT9gd3v+IYOp1ct4wUqW0rKm4Na55WvjasaTSfuyfwCPeFrAwU
zcx6J6hyS/agZMAr9K2L8cRpmlW0NBFSw7KJLpiv5HarOw+UmatrkWb3fSYD7I5G
O1yvhmeD+GTgdE9KOlJTsqG9Z7Uc51iGVvAQ3gyr9ol275jJ756jXYvZmq8/Ufr/
ZcJw5aKz91F4sYuLN2fjQRHOmbHa/dpdZRngxDxTYXJp/hL7L8rr4ZVRwtndkdVm
2FoVHdOQnnAM4L808GvH9RjoXnmkh+Pf/i6tCqo4ibv4x+vm1ENbo+YdSXO+78hU
Un0U2GuOGolo9hsJDCJn3EVnEZVvPnc6ns40jqGrzU/RotICAiJ7VgnDRl8o3cXB
1QLwReo9iZLNeioO+cmwYYY9O29II07TDxLyEniGRhuTAmK9/KX+Tg7BTlEJfxjf
nYTdPV5BRAuLMtSWQZ9b7fC6LNRdQtQ+jDcy+/liy1LmdsAPFhaNUQO/g6fcKg1C
cKYN9qjRf0fTNvMyr3+3RJPmiXoGyzW8ppE4Q6cOHrHVwe5icRKZN63EP9EJPaJJ
ZkoWdZp4sgnsX1Ejrt/TOEhT5no9ZrdRdWm6dqT+o7pZfPeLx4RUgo6V7OKBw3fb
2/+iDvTkCcm/eD83Nx0KzQLoshYWjM2YWl4M3xexc8RwTCK7IPwszTeDhwE8bC0v
Fiu59787mkN+LX6aR+PM0tMWUQO/65EjHFSWIXiPwsfo7QVO38L18eEQb5olvGZi
tJzK6aui4ITH+lvwuYd8NhDB7681gdfPeSEkGaLDgsoYnw0Tob0eAcvWsWQeb407
2E1zssnCmYNv/czMjJ1ZMGKTZCFniCJ5ldzeXNSHfkaIaauPTlLKsvQCBVrComKq
zCVhP2esi6Ouqw8culRvbe6iW/tnqJNxaN2Psk31tmmbveyHegz2lDpE9xcAw7HB
zlkMmZfV+KiYfJHtmoNvYikQdF3SYrm/rV8EKClHUeKdmA0W9j+ftQX3ClKV50rM
ecXCNAvbRuvXWZufvpjWCP/ML0erSK71i0zISpi6hxLiShMaqJwLJZQR34wKMqEv
Aqvf2dy/XEpFrPd9lCcXoAu0u5Wl0kCFwRpwXHC4yv15t6dvtXu5cVa6qSmyc1ZI
E7bkp2hSsWiRUvHZaYebqnMfUrhii1i1dMZl3wgh5qjZ6YNBKh4QlWE5aCEPVvp+
5LDMbKNmdE2G88vrVAl2uPbZCTjwTcZWHEs5sUmZl8d7kuP1S2aCKw8RsdZpCgIi
5ntIYDgdEFNaYWfqJXZWEfQ5Y8Ir1tPLt1pPReJwU/uxtEnjEYPp9Rm5qZH6T5sK
A0RlzVRQY6Uh3efyXVvLncbui6weTG5bD/4UIxzsg6f1jIIXJTiSNKYcH4EFcucf
yRaPd34mCFQqPYz8dq5ox32Acq6GoJwwTJRYgbSbiEGXO/OHHahpTtAx2SP6sA2N
taumYKwbazeabPOM9xw5qbVnDWKl+EZ3hTuQYiKnsbApzUWmKuULt9uRfSPUUHan
NuUJSym27PzctyJyUGlJtGDQaYmt4ee9FElwgZ97MOYXzhXhTzh8sjl079w7TMrN
hUIK1CmxJaQTEOKkRyOVG0Q2/iu4KSaUgsDmP0Jo4UPffvczhwKlyw9g7ZOZ7UX2
Nf6lJkOQwFy52me9zrfS+iRJgriavQsuOblcWZV7/7/mlp4alQzt9b54/qUGmpg6
7g9IzAV1iOhiiQs4FUyS0IQ920tK67osJjvKAYRiE6RY3BZ/HYj9jCzigxA8kMH8
FlW0531J0FCId4vuOj3ZPWTJdkSOb0sfGbipOoT7I+PPh9hptNifXPMZaCAGcSQ8
QlKYy9/2S2g2kNMTT0duGBKqe6UsQ4POfg075jITzzttPtksSjntfE/jJGaoTP6r
EIS+P5NAd8VdSwX2Ck1o0J33VbVW2CfGGussxU0Y+9Aqi2xOlZrf5jsO/qpifnrT
K1elxS8W5xufwrtPAmj+0S4Xox7yrZlRB5THE6bQY646oa/Ux6vBmMMxmzmKZX1r
xy3ALtQ7tPTrPPYZ8pVQVrhMPKFMPuSfg1lQZXhgLXcpY5vluljeqd4+0crj3Ube
sFcrnoDMSDXVoKo93eJXEZ+GHOtw5LkBHuDT1FKLczHN2P+Q7CBnwLp7yW0lVQHZ
9VebaAxOo7q7q1UASbmqY1+6d/xMyQVT373bugkk1OpZCZX4d1sy4ZBWVI5e57GU
UhssIN7VpclZNspS2R3k3hPFf0+V3p6MQvcBpsDhy5XMBi6aFoeJruVoGoFypEB8
8KrhL3n/Hgxdu9+XPzsPNKMt9b8ftGUtgPx63JTZExDTj4atG+81s9OpN+kaHDRy
CYGYyUHbeJK4L+LW7mbXFeGLFQJbDcW8pzP7K//pVW1eACAdKFqEuWsVlAJeeXKe
BLGwherFKTw+XzPbSjAzW0cuBwrrg3oNTejP2oqnlxzT/D5mnbp/UolR+OTkRWPl
bPpd4mKUxw4Fm5VBHFX6qkYR+CuykN85oE9YGaPHvkgxyONIW8hNCcbKNgc/co1D
8b7DXApp9gNktVJdgUs8MiBLM9h5B7P7b2xjZliWpzITq/HbeYdkeoMopxeyTalg
FiMCLzV+TDpY/KWjOvFpX+XdpG1Re7FFxmVKvwv+Br3hEoaMerybhHLE+pMV+uCi
CwN6jQOEWIIDFyDYBzgrFvu4JT1f0/IlZ0fifbRFuZ/NhMZkpenl3etEFKc0k+aF
1DpIwWHBOBmFD3iBv6Os6baJhOClV9MuA1/KFkOLXBwko5i0lp+e1pGs9u2QqMEZ
NG88tCz1dZo7uMMW3SKTsawb2G4LcyePeDzKtDkis4fxvaahVRoJOsUsUU/5GSnj
fn3NNqZQJXOjeMF/4FRLADUV18B4ccp4Jo6DyPNcE5mET2AxYUMPpvjQTsR1d/6Y
eR+fFXNigp0TUrbNTP5j0IFtZpJoYFux4BWG3ekj94ovwHmI+OJ5uDd/yBHgOvud
x7IpGZbpRYOpZvHezdkYtPIofAxxoYU7Ba1DHQTTuUGiBXb1aaWzUJU3D2FAhM04
twbBbC6EA406gf6vTpymFUEj6+YW0u/7Nt/Yz5O67bI/D+7sk6vOoOBV20xHBM60
Dt2JY4GFZagwsVKB0LwP7v2xNBPOvB1ekdTrRFKJ/c71kiuoTwE7nXcJ8U+ao6wB
MMODS8WQBi1tyKJnkAs5Feg9UJNXsT/FgL/D7C7W0HuoM5ea1zCYFGQ29rNx/9vL
If7QurFSxf3bz08El9rPnJPG8cFs9eEbWEF0FRiIrIcE6yhyzDGxnYg5NXT948wq
FLU9Z6DrJtZEjGEfz6M9kSsBQs3eK4aFiXHc3AyAE4msYnMgPnBmkJQ+TEMPRXUB
XUMn7BkOq067z369K+SfdaCl9SlKbktYpyVh+MzeIFxhng5MXxeJzEWR4ImX8tfs
crsSYjtbLch2A1t3XJgwpvflcdP/KK4P0o6GVI8gWtdxwpboDyRMS5ze89rOb1zS
DM0sUEKmErJO7OqFSDMAXBAhNCZML4YOMQxVkG1ufZi2wZKZVKtJ/1qtJag8/PCz
AjBQXxP5n9Sypme6aN15S8fv832PyYE9vgOV3ZUEmwEqn/NyvRvhhC9k8PoX+TEk
oYv59szPusmckIOn+olEiSaqmfKaztk4iLX6hNvbP9YJrKEyoz7Zq88bs+hdmdP4
HuuJN11/ZLcwqW3LGSNEEhoplZbL2kqcBF3zu4YOWMQafxmd23C/nCVJ4HYxVlJL
r+CDETk3SjdQS3IbsYfmDBU+NPTYohjTEr0hZFSp5Y9sJgfUWWzk1XyjCcxzs9fL
mGmMSntu+0MyRjsQMJus4BVOeYL3tBiarVgcsKTjOC6LO39CreDJ/CVBl3waetvB
66B4vUMyxPTeM4C2HMW2+9pc0SuIt6utWkmSvWCW911VhwXmJ12KCySFMN3P4zyT
zefvDK8rgYU64Lae/O5tscCitczlag4z90F2XIvQL6x09tFDSWklYZzLxvXeZxWa
VX0AkzaXg/Oyp2JdN82cLKfESSW1YmWnDNBoLNmNMDzxEoXe/p2le2w6/C+eMCZV
acj1Eioq2GumhVNZ9KHvCRli1dap96NEmW9uyRbqbPr9RH2xBrWMO3FvJU0DdlLI
c1mXPZ+JR03vvsAjQIXBzcNagiOfs9YVeUPikH6QZKZT+EHlhkToVJLUgB6889Hp
rVLB13nrDXYm8Gegr4A5m68llCC+ITxvcD2kMrR4uDRE3oZ/6SHNjM226medMtm9
GnZNzKRuuzf03r6dVmuPZH70MGPmfRxCB/5gtxIbqId2/Yui4j8A5stsEI1PS41V
XrIK1OKQAZJ+EmhAqxN5PEf7yVpwoPoMxnC+Iul81vztjQ/5wJX3cR94x5cKz2VZ
TcbEYaYhF0Vod0tk0Iw/B+4ANc/tvT99EZu8U9cYfkvyFWGmbl4gt8seqKYjEKrv
sP8Co40cU3Bjv4zlQQz9EHJR0WjpXfTcuLI5h84XUdZbJ2sv1uIT7mwCpJjVxKrw
OGl245WD1POsxrrkG5YRCTPPkLU2GQVFnF34WhkLZNH6KlMt4ui7DqlnLStVd9Ci
+GVys8COO+BsOLDz3/v34SWVYsl/9W4wTWWtotBitA1NlRB5EhPiBBRV5FP7vCde
6xa4G2TujX4wqGYXofOus7xzuwpJzIA/F231c0pwP3woNFz8SRLy+noadWKweSKw
Jc9hgbIiq5zXK4DhTTuENcDN5qoiumXKTIQoBCTjivtyo4GaCsnO2Bj+1s3onWuN
71T/N4nL/JJTCUA2ZAVeeYHP8bvxI3TDmIAwHdZ4t6mFuPNqFmiKefDtmjuJHAuF
aeBPp1IkEJEbKfjjbr9np/uSNOr5GHvAy5Q2mVJH0j5qygEK/DlxrNyP1f7zJpIu
cavJORGjYp1VzoExGF/egpnUbyFINC+yqTKg7Pbt/M08V5nhxsfPekse+lg75rTg
cg8f8k+hwKQUkH8Ie2nldpaQdd+33hmQhH2sZAh7A7hympMdFjx+v/OnfSO245uW
FsJ3WCjKGBOMEuMUmmTQz7DE1vrhRrqVfm50Zk9g+0D3BKT/StAMN317ImMR1tuE
m7DaUGC5qJ4ahHDKAIKpqalImCy53+0Nhrkz8FqpYqAIrQTjBRRWNacIH1e1R64Y
u15O40Kd9iTBSnuzpjtygzscXg13XU+vCrZpgsUDP06hLDoyHHVlnnsjRim5n2IB
078Bz8vzEzvWwgY/ANCm1zCH5IfhlyVcrxXkdtYB3N0QZY9Ycm19/hgzO1BfsUyW
xRxMp7yWSS0AbYkSIsbD11y4ugTIvqjB1rH+4P2RCZguhIalTXX7BQAHF9eij2ZL
3x7hNankuO210xaqvWz1P+DS1AFEVYeI89LZ2wF5Dji1cWIX0Cc4vWZTQd1IbLrH
B0qpl9nZp1hM33zbyAh8Vsgu344H8ht/pfWrpRRluD0pbK240at+LEgHgff8yooE
ua+vg71JwK0lr6sLzLZUrG4OadMedfVY+W8rvaC+LYatNLh152Y8RJjPZ8XF3AqX
S6I3yZcmgEBa6yxFdIxMoSBqVuLoVxT1EOQRVBRuqPluYv0BGHZmFpLd8lKdXpIx
tbyrEQxenyuRPanEJN/dDI7Hmws1/EPCVynO9u9z+d5+bsJI1Ur2k7Nf7Hp2L19I
ImWmEpWhCL/GVOhZXgB9y9JT6FTcHfu0v+jFc4G5DAK+Hb22KdwI693CZX3iaOI9
ENscc8s99XTQYuhyUNiZUpwkJMIUYWqvp9fWMYWB7+QX12AlfS8nyf95DO8DzyNN
LKloRbX5FLV4RHkoo+stsmPSdyvYsmH5IeQSFJ92nX0aFIjABtsKSbvKYg7OJjuw
q3O9LV9gJB293RpZpKy+wEc5G7juktcXtI5k8tjmgLYdq/o6JqzdiK7UwZiD0VHk
Gv8KGAfn7dhvkFL+5ecIpp1KtaXLfAQAj3BfFwWngJUFRY2+aI7IV+UFmyy8+r+4
uoWlz4h42VtgutXjRFyugWwoM/mbM5FVPyyc6DDwIjfnGAk81v7CYqopYbrmXgi9
vYzQLmQ3YuyWyakg67UcX3e9fqYn7iT/KPn6Iz2ujtORFUVzzgR6NzK7Yk/ISUED
TwR+MHkdJIwiUEHsHKH09aFnIS+RkAzqsACYKi5GnRSbqzYbbVOP6u3o49i4QkSA
2Z/hNhdZEL1nOCOpcgU/F6eXsKbSKHCjo2vhjUz3VqpqMrAzrWvYCFZhTLaYqUyF
aFdLmMhglVnHPLLa4hiryRWQ+w1lFdyROt+qJuKdAxRPzMet3PJmQE1jdV4nYTeN
m1HpEJAfClo6AX1doVRu79mWdll8b7BNdTrqn2P9FF8o9VQcmPzw9IuMykhi7gZk
F3G4Eqb6rCcfea41h1zrWQkf8ket7hWn2oOWhtIBbRSFTF+1YSCavcZoHGP7CXuz
zcd7bMy15xdNa6qsyNY3kh3DLTwZ8bC8A97ThsUCUJqU0TZ1Jr1smIr9hguJYDpe
UEOe79qJdj1wOE+GNYbx0U8sPBw1PuXlHY6OjOI0NQUoGf+6RhpVHyqOY2B7KbwT
U0xonpZ3A5tuPWwBPjm+bvpnX7Ql/A248cjTBN8HsDTGev2Mxn38sZTBcIeZeRHs
KMDvTaGvsNKQ0toaMMxoPOBZdD7NM1SnQTbU0p+tgOqPFpRTNFui+f+gjLJOdmBl
1/Lgct0FkfCYXsoYwRb13JS9P+96I7oqEJ8oh30eQOYkLsFYO7Wxjvqv1QR94SNb
BhF4v8WIFGyDSBrfjYNYQ0KzMEF59gKdeK8L+H/d7YxNYKA+0lPdCg+pimrT+3SJ
jbBb6fFhrk1L+f6A3oNpu2439qLyU7nAq8//rFOgEXPlwMQuVs39ctolvCPoyWVh
uknfx3b8TM8fC5mpJmk30+VHUkDbIEy81bFoKkaCIoCieL3W/hLKG1aLwbTXNbB9
f9DQYs/tNTsLS86QidaCdwWwliAfP0b8UdkL6UNSuEjturDxJJqBrQ8HuES8mh+Q
Gi3vmumOYTue5wC5MM3NQjIS9Jun5Wt/IKgw9SM7DO6+yk6KcGA4KwOtTru0jaI2
ssH4M1OmvDWyFQOpkfe9EpWdLo6ikUZU5pK5XRM3G0hxF7WxBqj0OXxl3kKzRsbI
js88Dvzb2QOCXVIdaRuvuXuKJVi5lmwJYiztwKum2hoQTIWoB+8LWuNwRWGUKwub
HVGEklUHytVtG2HALQbXfqBEDmXM7x5CTI0Mm28Ydjc8ASmsuCMP69BP8Ytv/yhV
wdlqPf3e7u2mdAy6oEudSEhNdbZYdkum1aE7xk/7JaBcihSjWiyHCY5uCR6luO8N
cl/Gt11G7wen0U1FwvS/guidLmA24gPe/tgnY3P4XiTsKFF19W7irxBQoQGn+z1v
KowIByjcpMGDWyh+z/9TfXg3elMWwFTJsKJp2RsU/4NjoVlOIxd6A6bGuIkvmL40
HTXgUGtpSOqAxDAIP2cJpmMjtvLiz7KhUSyMZq5tv37fpSnx94Nly8X7qnwSLa51
zByUjl/+d18O4sT17FVt4RPT6Jx4uyNX7BzezRFLtpHhU19AQPEVGOdi7Bx/XrKA
Nt4WO891m8liqLn9lgprPUFf76mgPW8cccgNJ/pqi9reSgCzGOTmTNZYS3I+sx+S
uHm153/SMeTtPrMcVpM6mgDU+z3kwJoWKfogdoURxUaLrbQKGPW6Djn7FJXsDB5e
srsc/w19JreDSsF1DHfKb78ly/Lr+JA99bW8cuZu1y1vnZ6ZgJFCAkimpX1DvBS+
eemd+cmJWOZA5BagqHxiTFch707yvyQTJqCGZ7GACs1jSObcRNeEUP0MZWlx0R9o
mwHATwNqPWiRcHUpG2/YKKrl4v7eL4Zor534H9P6/F/TfwYNLA61SKaPhQmLajQb
6EGiScsW58dVBCnOp7+R7BKQFnKTIpVoaaNV/cVfB8w48Hk393HIoLaAf2rZcvGN
gSFyuIqNQ03PV+jj71E35/Iu3KSK4YoLQLhXptpXArEmJXCOI/P9Jari71FmRmaB
hHLwpuKJfM7ELWcybCteJV92QtN7U3ORXPuNcwYkbHBdyw6x24fPfMrhC8u4WDkO
m99xhvNLM2U2poiuAXB0ldKV2DOLF/bDPsWtVuyObv57O8/1jbMGdR1qNuRZQaB3
M5zkBQzj51g1V+2INmu1ezBdFjwU5NvpoDVTju1trdHRcBPm03cMm6z9efSeyCsG
YblVVFR0xrjWaYr5JU/cGtlxrXQuR1eXafvURTZL1vmTlpVooFJLMIu+movbkJQp
aVcsZps0bQt33aLmI4iUas7bla0thYf/vIqLPnUa9Ze1+qGyZwQ5QZtL5RLPAnZF
xwMssY9JQ0HGzk4ZLvzl2/pWgJrKdJvuyiXHRYoLWNZsxnV6k8jQoK1w44NhgMG7
3V+4z2XeKZ5bOCN2KqsrhhiQ1t0Fnh5x9eTQBj7plutDYLbf5CV1HIAL/o7nhxnw
UlDpOpq4WRIqku8IamiLO1XcCSLF1gQRs6G8B2fYhZf5sBEqWjvYrHATaBHx6l/b
zEcQYIMAlysLm0+6TA6uO+YXIjjdS1oRjUTeJ3ls75Imlm9HsFE01NaFTPNwYV5d
XR9td8o/32/oa5roEFy9e8sruZh/yTVBS4lhu76xhFbr2rZrP4fPKefQ9Y9hQ5ip
wSxQN//ZhedamhmgQ/SdQG0Iik0qByypVpXVFIGM+rJBtBQW5+DnpkttRiPjkg3k
5LufjYMTjSHaZ3BPjEFB08xvnWYR4uqththZ2CGMglYeZQ8vGb+akLgoXsESCCTw
kPQywLFZ8pKUf8EB66NdT1G/St7plTqDc7PnyBbYKDovByuJR+vuv+/fA0r4kF8S
p80qVf6/sRqf3I8MI7FqS/DoU5gL31D7urKeSYOaQFwG3PhNNUhHf4bo2ifDoL/P
Or9fizIiDOojdxLWKs7MnvLmt2zvcbZzWcLdJqzRnV/XcqKwTL6Rc3eu/k9SPBXN
MKpEYcO/ZKnYRNbCLrfv3zzvHw55S2hh83BnojvTOzT8vM2mceeoMW7XzAGLTJ4m
xEbOQrIjQFOfziLg5tJpKImSyniY699N9Zu+JH/L+1D+TG5PF1uZ3FH1E5S1OkV5
R+aIKlbtYPFAaQMq1akShD+xfHZ9+kUx7aTspLYEU4+ZlIl5xhHDq6bPtxYeOjQE
MjJfk9eukSSAvlo3JCSrrtZ1113Ied8jpEh2xgFSfPco9UDGyXgagf/h6fDDZk3g
dIbFWsiyNTQ/ic2Qbuf5gmOs23fluxFQ8WnwnFRf7avg5WDVAPkckUfuoc7nniCz
EUMP7COIXIwlV8B66wdYsvIvFuPHE9UphQoLqxIVOv4pCWBUdC+Gs+d/OfdttyBP
qix+XVpt7n8pQfXjASQtkFui5jeXGQfqRnsdwrVbwYz+KpC/AMbHqiHskA0PDXLp
HugGuCsjn99yI8G8fsKd3kiTob9N0qDezDwPk9JF/gLbiHtKn8/DUMxTIe8UwJkm
Q0H2IM8/+ZrDTwSNKBnFYhzg9ka1sdkMXz9Q5D6mXOpC4WP0Qq3YgMewqyYSmPHU
edTksFUa1C0jeSAOtoMNWaCeC6sJKieNQCP+h0jUggUC8r8Bw19Mb6E4ImVwWvFc
dq/qgI1d4ixGhmQlHi7M3qG/bu+GkanljS7UyOHcC8N9N4ZjmIYEhigHo4B1gWGt
4gMmroBCxQ8liYiByl7breC3aXzLHyn89T+v6zDmclaZEXO7itfVPgjYRujLYX0N
7WTvBexW82oDu7wP+SBRSKPMylOu2XDzwgtis8qIt5WThBAhWC/Ccf1mk97jEz+L
BETEqp/KkOdUBKSOz3xBe+unf6CQRZlk3IwC5/AaOErN2EaIb3fUD+x9BYwh0B9o
fVth6NurQb5/1gAyt5bHtl5uSxDbFGho3hdC910JJiIXsBXeBh9mYMXvSIpa87Fr
Ag25bgAbrLPrNdst2PV4fSNDSI33mUXyQ56vttH1K0FMkvvulNUSL2q5dVWhpwU2
B023R1mdkjneW3/y5/QLhgvK8rMrKn46JTnu3d/V9bKXe1udH+sdDvAYxArU0VhA
mHpp27Xofn0J6rNf+YNQmy0F2YFDU3rGDZ+Cr0NeXWf0ERtQuW/IUJT5GGezqhoG
r+POJ3wdxtykEpFduNGmUcsaad/G82/656lgahEWEoDBVT7GFjcunnF0Orp2wpXH
H4XgufCiqPW/Hnl/0Tf/WfvVlNUAU1+haP1ZBhuQ3rm7ntWjHbLKYogHMWfP+REf
o35ZoRPAq6RtjUqEDErrhktGjPYNYpH3Ew/XgnRSPsZqdmHFoRX4tNpYwdnNvI1v
mDelZRgX6ZJxJrgBR7D1rQN0BObqc+EEYW98FUUfF9RhgT+StRT4cvYWqFFd0dVl
nQGWAO3cYbXd7IX38gK/nLky6rEmsWNU9kCg1Xvllg51ohRNbd0wJ6wB8NQRg53+
baX3J1kkVpLkiL+ewQWJsTQnkCO96qxsx8Co0dsISisu1UTc5lp/bF4BqhShSo2H
1CeypQVqv5sXLiaaw+BpHJ0N/bfTJwndZ6ytt09gradtGjc1GR0B7Pa5dBCFSvOn
Bxei8syUpXmpQP746fr2nDCWEOgLO1/VFhZCFn9H7+nChqMH7OkjitDmprVXnQBP
UH87azcinwDBgF7oIJLGxOsaMwI85ArOp/JWd0Pv0jhQsFrcXlMLByEXzlXaU9mK
KCUJwWHO9RFewS1ZqL4UGP2JTF2ieghmANxpNYiK4P8CYZFLVwA0d69rH6gZ3G6l
8GM/tEV9Vz/V8lDnJx2eeG6CaEPwOtJiR1dfLuRjbrC6HYHSScjqfmIwBJQy5h7+
2ZQoMhcrH64OkHEvnXCtOiVjiOQfSq90zVUy8+oG8e7ILxsmSjxRL6lMp5XkQw7T
6CBTmdAoy/I8NBiJgmozUSvViryINNjBKg+7nBm9dEeFPRhTcsWbtxG5fZFnu207
hgMtUCtUUA9nMgKzMMlaOVK12nQY6R0f5jsd2ZgCJAsFGDG/6XVSldmv29tX58fO
6HfKQOluEVpQar8FuMu60X7QkcP3N64v1fF+HfueYRvHmmJeV4O3MWrgQCqnoVeP
jrrCl+QMa/Lfd7bZ8YBhppfhxWRe5U4rxjdWVQij4SlSmXnwdCYbrAUWs20CGbku
YC5QcW7D5AnDNNQtSuhq2pCWmLXGutrtgGxwQw9maxU0gwkiUua/sjN7GPcRLsXV
7yH1FZ59bOfePqv5eqeuDkOC7tm3HXsM75Ynjj/20XXM1LW9k70EBATOaVlo8D7A
Cloq9UPvl0LUTxaw3guB5QWA41Qnp9Iia7VbGRJuGyomu4OJG0skJE3zzpzxOKW1
AzowJmgOCM5ZM+7EwtaVsctGILl2MvD7v0JI0hVKRjKEkk6dW22BE6B5aFguzKtk
yQhs2/tKIPDq7qqM9xszgU+22FS3NVRMMNqbAwpEHiEu0WlwCk8ZUnWBjxi412d5
Zhng9Ad3lXqrrXA3VmeIvG6o8YkeO2BUgJ4ti7totnKOlAa1lVAHhGMkSkI2Vdue
B5qj/qu/d32pHUegCQ992RiHAhS4pUYlAOWr4JLIs8ymH+ORsgke9skfJj7cihKn
8QKNx29jXvescmUVxa4DLJ6Q3Xu+D6piUAHvLlaUfzjykQ8DKC1TkS84RR1LGdb3
AJvoFkV3k5nqcczATBTR/eeIC9kf5DLeYve2x1fjPZ3l9y0QfMMU9/LWAb239gYD
63jAYxywku51SRgvWexd/q+RKq2BoCnTj15+qIjdarU4wnoXPxYMLlmNrl2S+PFk
sB2GbzS61O9FKxeHdRuMXZBQGh1usbVDca2w21MUppEtiXQK+5iDt+zWV59Mhg/f
fRkOmQFI3I6xpuOdSa2WQ/CSSvuYzKGp/ck3cmgExEko5s5t9DhqR+PaNifFhcyk
AlUeblOzK21wAQw18DF/pPzztfWqzbMjgy3KlnPCfCv5XbuWhANbVpv/j1/PKmYD
IdJTUVe8wuW+fPfKwcYzsoDo36efMfJwOJetj8dSQEFbmVAWUGodth7Krs6v9EcA
if/l3dvybgLkHn1vlFwvJcV6wxYZb2SjUXuATD5bKePSJEzqAWL6ILeZiUnFySWy
umie1C+Xq9ACgUe/ZQzlCZEbxOAFeE73Tc+6oY6Rkm7Mke5Qp025lY3+TToUUgjF
+C7YyMr8og07djGFgZ7Ydvd7D2ppUNpKtgxyFwwO33IEcEfFHFydCNCRtYLGV+G+
DFXXAAGZ3t+h0ReYZ73nSRcwJeaHDKDmruNzwogZKEF/bgxlAnrU92l+uNUzXQuK
QCJuHM1tryBGdE5C0qTA36cdAkbspz+1YLblZrx7LLZKrzmUercOopTSLRLr+h7b
ZjkUAhSllwLLBQcern7q3rQT5BrAtb4Dm14+3IJ+Fd+n55WDttS38VaMSpW33jY4
yc+tiUhCZnOrzuvl8AMT8uilJa08sZVz5NCwnoEmbrVyEBsa4iUzC6FpLaznB3yG
QvY4ZpOuVSRLiLjiWRE7Mbr7TvmwEtRodozuYrDtJNlX+cWBRrEl4AScCgoVTBuO
lisx4bXwGSlTUUpRbwCG5TDD47XzFPSpVYlEK5GfM/aiFrgq36rdmEx9g9RtbNMw
UmFUF9gT/CfHcXw4ATtvzNYm0iBHMX35CwneWr8B+B8C73pZIrR4ZBf26AzKMR3M
GHlFGJihM711Nft6i8SmO3xcpJBQ5Zye6ZmZ5T76q7YIn/LGglmTN4YOMKtsvafN
JRfvYrnouuS740pVclpoM7B4ngf0a1d/Mc98TyGhriw/r4VFZRL1T/U0yXnraJh5
XytzONroUibqB6hytAZk5Vms/IjDIkdikzhXRob7HUU3gIrklotuZhgZD26FxYyN
x/YRLTH5cQfZgNcZdVYN9BeJXIoH+0QuF7TnVx1rcmQ1o1WVwR6yy7VBG0pbklzO
eON0M7cLCvL3ZKzkRi678gf1WVrfZG+HX1yIxjw3qCrRN4SUJ5YykXYum1Ud1PSW
uc+itQlxLuWBfmWZccAnCK4k8Z2nZoLc3+38YrluQKaJzb1hMfYdf9xGhp8JCeec
lD/vJzJXqD8PugGJQG01XNwGHIkNAujIFrpeHntCNtJ4jd5oA4VxRIm04eZQzgnH
W8E68knkpSwjz/DldlnURP0rJZB+2HkeRhnD8WLok0ZiZh7iPqPx3ALOywLEULUl
QuZRtwX9wgVYqmRrCne7GG5DcG7E+PICsx9E3etaDYI66vIzk99dXUWJ1Wjfzgmn
nbSwWjhzEpzZV31Y/ptLdVtA7cSpV6oP4z3+rQPV4Ft9PS35OcN6QAgelpnRCE8a
PDjKCWQBFIa+sjPVE98hgGzWlbcQF0+ft5SKQdQLvQfWKFlH1vr7JamwsfgS68Pb
p975Kmm11RhwCd5dr8AlfSZenGOWwLY3Xk3dcvkUaBcHLZ1Q6l/5nGaj+RQbPvBf
JPUvb+SSCrxzZMtb3W7+qyOMVq64R0zBP1fHoa7gTQarfWE5Jlntn3ZwUJN290Uu
qiNixbCUq/8eyM74lpU/iwlfN68lLkSIszwwNss5aKPjt/OMFxc9XXdS2WK18Qql
+06Dl3ExwjHw/UCMWRi6UDwsgsgJ8+lG7UMPPj92lCqgJTCiYfk6aRV3XBAv5wUz
Ow0FqXeAgviQBn8/+XqJHfEVvOaUTDOcCy4gHugwIEjWP3MUVYHTN9nJkQD12xLr
IFZ0KhIfSXfq1Y8f2RpbnJBckG22rmbWOyRs2JEVu7idpSeTIOhJiZLYy1ZKSU2c
rT1gU+A9B+GAg/TX9K6IGiThHyrO/hcwMsI/wYCrs+tmcKza/BIu3Wq+SM/zDNOv
z+VYpnB70dxvD8zqelKI4bZadPkOfeUeJ82PsOF+KAHe3JUDqftTlmuELyLCOvPF
0UCT1OzF/CQTSYF4GKUAo7SWJrDBs4PqxgKV7Mb8e0tEqMuGMEgRCcUrbzhO+JOo
aQyYzibBqaMrgiuBIVAvoXq1sx4h623YlUwXkiMyTsv8IYA5t/qJXyuB43Q0cZYH
pIxYQa/vGqYQ1CdgNO/RAFaisZ+AX/bBePg9g8kpI6vrJ4t7Puv2piMgASPh1jsq
M7CyMZYN/I5O9AuUR8E3XXFtwtfYq9DgAN3xtk0byey6StFJSmjveQ7Bgu9rsEyE
K6TBg95wvDyUgVyRsSP277cUYBDAWHT6PXnThFbJoLpmESIeIx5ICxIZp6i3sMAD
VbVzoqHXOcSnn2WW94tI1XbNkJFRL85hsxiawyMH92fFIQaEZIoMloBp3NuVon4w
LGz8CmFveAyJnVTV4g/CalZf16pM67DhZHIDAefYZr6kBPGuiUTMG8pJTNR7scod
FPxdzvUOvHghcYjyFQtNdWv1AUKcxMwD1gmY+88ft1Yr5W7gNXDTPwgRaIGUNzzz
QaOArP5n/qLHzbv3Oexp+PJTn5LmwKJ1aSet5oAzDHt4BBa6a14ZtSb4hI094c5l
5za4tjfp5sqfsHHxAtbMjr+7xMRGREchgPxOf3uWF6Rv9EXiMCWnUJIWAoU7RAtV
PWnt/KAiGt2EtlDrXsKjGc/a0b2/7R6KjyIvFr5yA0FXimwzvpkoQufs1G+GqyMY
oOh5IbD/PTwZM4Wf14QR+cfm4pgMA3/U41UeKziVTp5BdgDEYcIJp9sqK4E2WSlT
yb54H91wtOj4QAcmvfcAHkI61lhWi+NWT0NwwJ9HScSw7rsrcMi9aJbiEG7dpHL7
5wJWB66hnqB+naXc5hRuKJaw+3VMRP2yjmC07G4c7T7roG6VRNl3zHCsXW8yV4EM
Bv3bLOf+NOQlNi9QHLDZCAa5R63wOsD0FoHIurOUaohskTkeEsF12Re7It+5R2ma
l1KOGNYT6MX6KHMPzKo7gbwdazuW20d37YE93IHTlXWaXf5pkv0SahgnEVmxapCi
HM0V0niaADyvG7Q9LMYekF5Ell6IW3gaeSOvP1hXpo6w/MjfG9nLSjdTHS2v7fWV
/FPqsarcQgDEOxF71ya/hXXsTXl4DldOe6sLczZ4Nxjm19kl/dir22DIuG76WNPE
aBpkCJjBepoPdrHr0KfCMGlb+7lUXQscHFEUkw/L66HWd6ln8UVO+S8m7A7uBbGL
a0WOnfjJvHP85EbSei0fzXW+p800kSweJN1HKWdTh6JKTIdmwZ5wjLAFcssbOudv
bfKu+kFUGENtAribkLNXDZWXBFg69tXWdfGLWjt6vZV4LjSFLjbp7S21TOecayNQ
3wqfBlx6QqpO9R04Tk/LPXJiDPOcAilfeB8ogllbiFN3IQbgWB/p459JWkgWUhFE
42RBAj4r2L2Edzy5tBzlsU0tNobj/cVGOghnPrpIM7shrtW/bTd2D/klONHhPz7x
atfYjXlQWpgqusqV2/WPnD0E0IrugoPmnmziJlGJd9FsoDHMb0GxlYlJ4l2Aq8jv
ctZYy6kZRRXP0G2pVnAA28hck04M6gWHzPvyclsMlPnYjfkcMLc6t0QUEiVl3zo6
9jQhJfz8fQvXc8/i4Ne/tHKY8sMfNt218YDxn6GNjwpc3XChTiJEND3AvO+o/cts
pU+xpdV432L0c7daZx+xkfCSugYOF/u7C8VCMmpTD1DeBinxVB/d1Azno/2vzyn/
2CdrxDLVZvLc31WxP8yyviJzavjYQ1UTXTdOe4X5XhIWjTr2uE2UZxbP3PBZek8a
2KA4/h5Qe4WkTcg5mid0ro+iIpF6xi3vYj/s38d5GPT7oOyVP5ffUTpCO8xB3hiv
o/BdZY8BcVkiC7x0t1RCu3dK4r7DDC4EP65H8YTpy5kw8p8uOxDbUjBVx81PTIHN
0dmHCHDxZ6pqVw/ZGqP/HU72RVThJEFJfBWEu9mEAH4IOyLJGO8RqfujCHIMa5Rw
j364vj1Gg9ySJmI3Dk326PvQl0rjw2T1q3WdLJUu7oV/FPgEAF80G4b+Id7Y/OzK
ziIQIyWAF1K/aK9l+XAEh46TCcfFi1UzQxB9U1FtwbQbM/7n8nOQlqI2u6jDkZDD
17Z4fRbF6NrbVfvnTt43oo++w8hXVVuRrl9WXpxxhvvc5kInObEUM+I8sZbOYKu2
tEeBwDjd+jStv/7CvuTphaed5lDemZ6IoX7aeZU/6d6Fg5KXTzYve2/Zr0AZwNcb
YSJV91zCwS7oOe83NBJYnM2Ksv+A3it5ye4LdOycNoiKzX4kh0IDAQk327uEpEfU
rZhlAHAygebKcIcxvREZ0Y02zZYBCx81lLy5cimV4364JPaUatFCKF84ex1T+xfp
tVBLBWQMZNOJ8HJjEXqxb8oRbqgK0QXU+JIT6vlHPnhBeMxhSedzreaEdw3AzZM5
iqxwXmtffp7kqYxL5j6qLagb3lWiwc/0rCyL4FwyHe3twSp207Lcs2EyyhNLZbXy
FpgAW0o8KH/OU0VTsyR6y6av/+7mQeKozOgSKD3QzqyhPkdFbHiRcuOPqC+psOYl
h9+z6pDIGRzDeu84M0J+xaJ3NpMpfldJcMjA/71XM+lfLXOVFi8KG2adQoWtFD7P
CnX3Z89WaVV/9AnO+lAqoq+uahutgfat6Iz2p8rITMkOyxHLd+ETJV89kGlwdlPr
7A2p6yD2fQS/ruwBM0QWk196y/tyDfvS0mDBDms5Mg7HwP5zG92VDAa67Cx3QRwC
jVs21XS5irmPO5WMBGE4YmeZE17t/robdpC2UNBGQf/F6Z9Q1go6Xvy/AIhoSci+
1G1QpatjP2iwXcR7EN12n16y06cBinEP9ITn2cHH8lRS/L1ENC+fS5bDi8LuFKQV
EMsGrnaYzg+zkeZJFec2aLXwX7x3lFtMKj1y8V2F5U3JcrglXbue5KMp4PkxRTjA
ZfBI7ICSJG7DjycXL0Wuu3xOd527F5973oNLhLQOIbsL/CuJ34Zp1vPgAdRr0+oF
AdSi13oeV351cReC872Q7KOYR+GvQEUqQ1FFf97doaDxRmy45XqVb8iD0F0y6R4H
DbEe0XN0ZCmxlHZAUcURNPh3vA44+tG2hMR/JExYoggrJs4ZnyruWuX6xGF1IPuq
VHTPW4CLq9fQBv0P634ZrF56VzgoYlU7/x3iTR7L1nc3LIeFYnKzeyyOKSVkzgrA
Mi7L1dqfmRFOEsFO74L0Gq1rI9rwFEv7Ii2WP0PWDkeSRcspE9mbsYN6X954faRb
7ttG77nXMCKuBuf6zlgP9raq8R1kh9JGSBZRK3lahKSLGxlGNoGkK/1OL33MwtGV
dEhMxZt70ghBJd1GsQeoOIHX06uKTcExtLs42zVlHt8HGX0pkM5cX4iO16t29wZc
8tf7w8iW8lynt0JrZrJXSOsLal9cqntQepTeJiVOmdg0lL6/nPZAXg6kxORfiWJZ
OQ8GaCD5wjehX+OSdrvRPCYcsxKNeU+yUbj4pnau3W3sOpsN/6H+Xk8dC+jUEf2K
Fsbd6TEtNgD/zlRYQgKItwDNsVhgCp6IWdi0To+7wDI1ZlcbGjFi/xYtQ0G/0K3m
n5gXDZTIhBqEgZfLaS0ET8oaHqhj042TlbpMI0xcdhwJTMHjseVfmSQN4rR1d51a
xdgryO0ikZsnwxpuOe2U4uB6JpCE3KLcwlxTq+vdCo0GYO5JwGE7o+r6oZZiB7OU
VfaBlf4qUzFmlG6bB+v1JLkzlI5GtiqVUtbg95dTI9DLZoM4wQRYtdrH0EWmztLE
mlMbzA1NkBpF0nt4CBDU/YVtK7CYffZH7Q/oG719RibRap0Bi0PzHebRof0zsLqW
qXx7bex+o1Pxf26erjwxuox2T8wksM6U3zDx9DQTaCK0i2kaTCQBnX7xtXVvy4AV
17AgJllUNjyn6Cz2pRFgKA1RiSESfHVoU3tNTVp88mqVfnkH0IcPGaVGVPxo2x+q
6MSb5YTvkCQx7P1dzNzak9Cd3QZ2wu6ypo0Rq1XV0eV6LxNhUvgMednhD3Swlc/1
xuBef2uUiKLYhpcCqlm/iAmT5amgHBTqA2OMsPhNDx278cq9MffsOvB6Yt/R+4nR
fAbU2rFoZBA/SFjsle8BxOk9h1G83LMSMZabDV9C9Ib9XhOs5Vq6BW4KPnlxa02W
eZkD1cq97jp+rzpr/SF6A+3w6VfZC1bhhlJD3stLzgcSe15ygJnI3mzTTRM4duX4
Ovhhs4YSeBV3fYgXbIiNCSCCYWvKGe23vac5CjMoiEc0Dgj8xKbteeTi7EjLHwyU
JuEMgCXWHpVMOm0GGfJ4/9wf0TBly4B2xcpUDL4wLq2IWUJICR7+6Z4ov1idtPNW
QRP9eyUKdK6Kh/tC8pl8BzUuZBRlCecLhPu2P5NfTo+C632LEP7IeYZnj5MgH84F
piRQyvBo0mneeucJjbzP0Kz9XuKZgi+eIEldw7VOqD0PxwhR57pf2XMPMxZ3vKKx
fLBPet+YOAJ3L8f6wppPemZPKhWsMbly7iIlt3Gg8rcKnrqDHUbvGNgV6iIR8PY+
rKgTdPGPaoLKHwjeNeIeEY/zoLpCsjIJP4EQwvo8Xjq+rYEhkXrKRttOxMFGn9nh
ZHHJVaLinPm9XeZOd/aGl3ve8RbZRVW3Ug3OgAgE5xkLZiVWKbanzWcbiitL9PAX
ewkXncTt53kF59Z2fLKQhDu9JJtQjgrJSohsRraWPx4KXn91C+0fQgbZnXcqS302
Gu3XRJHJwi1lL91Y8lv9xq7CugxMG7KlSvIouhdEd2asiy3j2me5E9Fo06vV7jpk
SV/Q/kOpq381o8DM2xqkI6l9heOqk5IpsiEZ7/+4ZFTdBAQsZ2i8R1VepcLv29KK
sFbmq7wpU3/0Os78I7uVMwIy6e6iSblm1+G0f/cOVV+job0WbtH8oRqd1Rlwfd1b
hGjyQFBqsVrdFB47l9zfJ3ao7pPjiUpI8jd0ZAlALC98woC9Mwn2k3BmfIaNI+zt
xKsdZWRwOFxO205b88e9dq9869WZfjYyP0hQGfK0hppR9hlHl6Hxa94AMS5+LFjU
4OlXXzzz2SpI+nrR1ChfE1f0D/R26EUPYLX1RBfP58KJpmIs/5DmFleXlw8PgpT5
JwAlQYxStOXNUpP6dJqkyMvMIsAhj0IfvUGJDvR07Mlle+2FWaVRg+/saC4P75AQ
wKVDQW/JUkTXiADsDssCsZawdCMkicQR/pPCpyihwwAiagqe81z9I5LpKrTGUl04
kM6FgofueykdviD8iDMLfTgZOjUAfWxgokvMb2RO4/CL1wGeSFCoOw15nrhY4JEY
U+sOgqQSJtq0gAu1jOuPKoPUDA4fXKRXMfs0s3WFaTpBUTG/ZcCo7giOJOnggmzx
UbU923NcQmYO95qNbFhjuc7WJQxnAEGh8cSzaErKB3bh9px4923RT6eCyy2FWsHM
1HXyrph7xc/Wj/jnD+pcW5witlikr4dmH9PCOh1qQnT/x/W1G9UP+EkqM5oX8/CC
8qCaU3BGj7v8alV3I5d94WOmbkA1E5KJYcu9/X4dPxgOF5IjNBYR1676y/DzzGiK
IcoIMUMcqICZh1IjjIGrno+FMTWUFJh+93T9YdITtRsxgxQQ+y2EeVNq8qEhT4V5
2VsnX34n9YRQF2cCny+lxeb1SVjO2R4XuBXHSePeZRyRTx74kezGE6utx53mGJ9k
CzO00zRTLFKLT3GNGPwB/T09SAzgYe63j6ceO5QdFqTX6y/8Y74oMmRh8Oxvgxkf
nMraJ4N35bKtgyoVbJbk/3aQ/M0PZcqWjvBi+ESI/IeoF/SYWfy3dzCRP+e8qUZ+
Ndgq9sxBayjretquqHefnoN2g314gc6BeA+rL+ZKmOqtgf4XUN5OHxSlp6oIhfs0
rZsl8RSn4CL9MmjwInOUw5FYmqYQgQZBr3n6Z/1kf+iJs7hm2hnh/Hmd3a0Wxti8
JH8Q6hGcbiqdsZ3U/Lf0O7oq+sf0/0YR9xDR+TEWLnoTF+CE6AWJXRYeUaxoD360
V0SkjN6Qk15oGPIOX8fKbTqEVtq0ijKrjp6+rDZU3O+AwOW168VuJ3komVo/xFDD
V490w3xRzkCPDzZ3OLcw2p+k+Sq+rZdcm9BmASZfL3YyvkXLsOP9r+cBqeSGay8w
Lk4++kDALO90unI8Ci2yp1kWf3PVYxEXZjGfrQUJmGvlmNVrX9giEh7ImBQYx699
6TZgm+kz8hMIgKZN5k36SBro1dym8VIfaHcdYuIMU2Cxqt95VH/hluyLIEeM91Er
44qFjOHZll5l66k4O8ev80IO9bU1Zq1xVkTfV2Rh1N5aErJJDz8MSaBoGtLImSWD
2j7VgKxk5ykc7NiPkKZm60NPQWkbd7tILo4BBRz1glufseOC50q69boTLMbez58b
2DZopTJFMLqaobIHAfB2SWHvIJXm2tkjDJ5m0v6hLX2iucWcGlhyVM7BCCXgRPvJ
aaE1X1KLXenvw/Ksb+u4AAp8fcX61v3y3DLMMam0EKNV1wXOh6BorZ/t+pfJu7kP
kW/u5SnN+QeVOvBLOBSc9l9c15ZiJJQJjwAH1G/fVoFu9jlxWsw/Zr9xYdYLymFV
KTCB4UkUVi069Q8dokQJZRMMtnVxLCvC6+pvrynKtEwKLMmOvLxnpbd58az9Wwbj
/Gqk5wbyJHpHW06fkXK5v1skVTKcHuEX3NP2B3Vl4/LOJvUHRo2K5TjcCa8CIGei
/u9L5yrZ8sBY74uo3AxMWS56kb2kqlVtnscqiaTdKAvGaaB+zGbPO1NNoSKm1V9T
8Nwunty5jPN8iAN9BXtSqLZG63cVofVx2JfJfQRSeXbR77tcmUd1hLuXNjMDDTJX
nYXanboxPXgjuuwY5DBCTrcm3iLCIiYncPezDSamkA7ZJ4Ncjq60Ugm1PIV3bJnq
ONGcbgtpHeEjp3zDWBVoZ79mUbWYghcsmLuKLThBMqPnH8yR1Va0u/W41aoiCI0G
jlbUFT0Hrbo5pt5uG+cfsdPcE3kaC6t70fQsXFvgNPPARjDHipFKoofz6G9aVzVk
6tbi0YWdCVvwwbelghSsm7JoiHH3HklXwPcNWmj7uW+yWvmv2iVxJcYbWSaghYuS
nVS1LlEr3pp7rkFyzyuObVC16YOFzpl2Fudc4uGbQ4IV8ehGcTfiisDY64s2J6Ik
XQi3tibuJYumR2ssEd4djvc6XeLbZRjW3OQNLwi6OAzf0x5l02EnVflu3Ak6lOKd
unl3GJxQS3YlrKq4ziqEc5zrlrgPMD3v/iaBssoGwc2cq8XmWrBWCLVzotkCJvGM
POkbzFFYQU64jkh2kpNwiwGWCVjPXDYnxpdJOBTsq0WF3YvpZArf7e3TN5DL6CRu
zujjqhhs5fABYIBOqZwhYp7/IBYxhISV8zZIJGp2DCJHvvqIO9hnGcV7VvNv6/dx
mnEhTmGcaBSQ1Ue++ahQYhcgchQKOpqbzLnjD54nIdubz8B1b9477WRK8D4OVDrf
aSOOCOYfLyp80CBX0Xf/XuQgXoEDnRt1zaYRr2ldIGgQvadyLbRUhwtvpfL3OWbR
vqJPTSTJJsGWKAAbl2iLjLG0ZzO3j5aFkiAfSVY7YBw9JRuJtgq6z3cLD2kvlLug
UdXSAKpJVg0LQ98PNz3RtIOCTCrRU0ECwi1c4dYFNrjiCvm6GjVII4N87RyGsPv8
1mo6vhwH0OBVquDJUTzhIwicjrT4mvTNlx4NKQFUCN6d4dCwYFVUSvp0RrtTPPj9
afnPeHDiC8PLJLKUNP1UVRRsQyVZibsqMxIJG477dCfAx4Olh3sfKY6T44euJ5Ty
b3KAfeTVpmZUEM49XemKHEhtcjU4ry/k0Wq6+6jxrLvhFcEjLuSDxH8T3+TkGP1x
s2COTZYH0c74o8yDXNTyODRz1fneblPu9sRcvph8CfSQ/JY+TdKZ8jggpYHDDb1g
+GUJXm/cxGhYq73eHIrRdT8zmj5yj6qIT5ie3XmGspSsf76VTnddHJOd+haTBeOP
KNN5gRXeo8XBEWbMlKvQhROOJ/2FEWc39DjDE3x1hrkud2RgUMH30CHXUbsRERS1
V+7kc1WsmZoEbcn0brdqkFRXrCYyc8v/mGoKlmzvtVcjnAJ3vF7pz2NJqL1+SpXb
/3Jl6lsz3Mn0i8nbmSV9usFrzKvPBVNiBPmXEO+kWpnTu0xetTlF1bntoPSephiR
58qEuWGqOVOm89U/UPDoAzZcFvfEOekgUimRMmjG6Ky5k4mpdYcetvpPUd5sIkEk
vFZL0wu8L9licgwNW2np96zIln17NE7W818ThobYNg6RwNUnqRqaMpCCmXknIQGu
DLOZ5Ob8K8V74BLPbb6QWTrmHeLqKEESWvqMhKYUn+WXYc//rS+VBi/nHLUARyIj
z00GTuH25pkCGRhSaAjHE1YO/29DT3qBuHNborQ7bH+F1/n8tEcv+GyqAyKF3J6f
R0PxrakkE8UwOcIBfXWBq87GN0fuNKfQ7PDbiMqlPWfz2uKda+iGUkkATLrlmTSX
/wclW8WUP3DgtjGXtfYY0nxKa9ixVNnQBgckKknphMrWfB1JJDGs3G5KoTyRk9WG
UPHze1PtpjaktVZ2ytDJ8B/rGiROx9v7X9m3v3FciXs9VT5PR3uRgDpqGmy4mm5S
ihtllsvpPQgBgPHUiN5RF2NL921u38bWdBIdD2f2oYZjeEnYQd/GWv86dVqZanph
1hEafibK1m45ucHH6k8kCpxRvzloeHenrqWqNFj7SDWU+0H5O6AVK9VrT33Hlr10
lKQaIOxeJA+aqN+ZBYz9tZJaHd6zf1AdvYTgpI2SDPuWhyF4FUuse5rVGb61Dhif
9iPfgfImPnscxGw5HfKclO4kzZ23UfMZ2/3Fpz4aHinZ6FtFD43/kmO5f6XHbWSN
Xos6alySj3UADI0zuEsrs95irnmUxYbkBKyOydxmlUVQQFL8XLq8vClf9soqHR5r
LaZ4r7BcnRF+Ozp+yrucR7mzE5su24vUiQuIFPUEifi7YnrZ1W3leWI4xi2CVmb2
enKcgh4sLglrCMmNiXmlEinqXwwl2wEU3tl91vTqQRpM4M48ldwjxTiPQ5r8rAwR
bJzFkHiXUK01oAS9Y94gPm2LwduZnlYfNmnrl27NqQ+NAIC1S6lRUlrAS2eyfF1b
zOD2LbNXZv2jhf787T0234VaFzF7UpHOHa4jiNBQQ57uq7TE+ozeoHSH766zJY4Q
y7TPlzq4tHJ3W1t9byLCPHFNeGz2OUXpDKidAG0RXRmznqKueSbnI5XyzEl769eA
qc4OTkZFnPL67jtafVRd9iF6q45UeghF6rX6zjtGWW7XAogvhdkbL8/Ctu+nR3gH
Ie/00uTs09eY+iuNTmKZg92FDVMfnLSFMwyx4sRV55wOxVMOXorDgJgQfh4uS8Bf
hKjVMKwlBgLO+yB/GxQIqgstCerL8Rk6qBFKSmDhHrxyECa5K4jyqMYpD8A3Tlkq
yr8opUAoBSgTYM41hf2JKaectUPdolKEclOh2rOv9JijWaEfc08/hxpaQRH1p6/r
yN575GubOV+3wkbwDT0fzGnKnr347k+hm145b1U24lfStITfHWAkDkqczYKwd9WO
8VwJdR1Q1fAWLgWs0DDNzTTz9QI67A8HBh+8VtUveNrqDnBnWgr0swL7fIHAP9BR
V1JgH504KsvHwr8HrBRw8UPNBQoRxD7LAIy3K0YD4keBk2CLFpf7RrhlmS8joVdj
bTdGKUBV+LHdzjfMICjtAAKeKsUEYqThQo0Qh2VGylbYmfk736EhZckCIHSFTT1B
1xIOKnCiUyIYyeZQwsD3X1ND6DG/h21Lxj/OlSJBED5ACnAwvKqrYt/Gx6mukePn
h015CSlKi5a1DB6wuGOtURd/4NYy9esI7Ot1+B0V5YRHpXj4w+inkzl+SF7Q+Rfy
8B/5CFM00DiPXbMtWx60/7bcWX4SJjFB3FrvxgN3xrBdjMefPJz8xTOygCeOZsUd
lBP9HQoU+tx4nKehhCyWENOkLKl+J+jxQVm9AuhoLAFnZNyQCkfpxbyuhxSkC+Y/
LUl8mLy2Wl1e/zoQJ6qF70JjIfSFx21jncD9FG1NjafYiBLlwg2TMqWjyw5mWfkj
mwrfSXsaF4bMLyY5UgpSolOTEvmZoHCKbalda2OqUtkO8nH22M+oJJJut6AAA0Et
WD5qre4XdCE7ILptEgVazs6l45kN/QRwJq8vrVOkfXXDWhxf+Dng9jbrAeBlY+1U
LVBEmi7LBTswr3KFtaOeI2cV/Xlrnenr1A6GnFnx7c3PbeEHjpbiIxTtxvcBkeCD
PocsAIdqxig7HfnLjwgDAmJCULf5iewdsDESqs8CQLNnnD9LYuvXanwKfULTWVlj
gWmKET25NUvU7Chzv8FEbCvILrqI/O6uYfSijS39PaUWWs0m0nrR4DHUzl6S4996
aRq3TG4h75PvPMf514WXwlLDjphGQ8+ql1dXRp8+RnAJJA9S2sBCEGIbxpyurPz1
ybEVgPrcvBOzoaQkyprs+Aqrd8TpybPey5kHOuL8N1FqjIfcGuVmDUCUpdHW/P57
q/+HPcaXBGW4Mcyu3IJ/uUKM625yHBna2uyXAmTcp0Dgud3xfLg9sxQ2mo+yt14W
OPY/LU2npeBu4vuqmApGJheyGu0ttApqDACtSTUiSm8K6pFwCEROEMCCUwq9uovF
bVffr6Lr9Jx2sRF4wCAIspfbjcfcrQWPl2tuCoxS2BygZ/nSLk+wJOF16HRD811s
/i0cJsaKP2i+aen/srQHv+8P/3/3qj3XEI2zuGkWbmffuiKNESFtLAsxzcuE5EvT
UjsGbwiF4f7wu4pnGK6wJuMyDhEWhtEBIU8NwleWTaYEmLZg/QugwXF5hSdO7c0e
FbRb1cgCXSRXKJ9WmLvf6kV+qEVolUaOY5vfgjICCF14d8il9zpCwtAZ+W91gusb
i23G/wAN1Od4Vl0Z2l9hdSLgvMv7R6SRC/shiR3H+AM2HbiYjDJ04NDOAD4J7Cs2
RSnjXRDYZPx2/FWjPHN+YaMcHbSH/D2f9ZbKaJCQM3pSDrl36nH9JW/pWj/5j1bM
jonQKzORrvgnKGVS4PbCnf28T3X+p/PqTYV5icCqdZMBwUWR2L+t+8CEWaw+MJ6Z
h5NIProqVVEcYpMZ/bhzWxtpzQRMcTy2JVhOqsAx7F0b3TQjL2fX79BUu6ToRTFe
pGVtZ0I/SaagNRMca7CBJj/qh/L2q4lDIjNuVrmFS4D7i8ZZgUQWSL4sAfbKcTcB
FZwVmx3KOtTOC4lFJ+P0lH6DW36tmMNGdV7NWslxIq6GiO9GA3KbwQG401Oh00fd
GiVv5zIzG6xB2S3bBR5Uz5Tw1cz+jP0e/66SryK4ULojlzKPVDaKTev5My+X0zBY
+lA4o7gKwFu1Sge3I4Dx+KHVLFIX1yLRaPjHxt25T0gB/mOq8lg60W4S4K4Gv1CH
+cDBuXICE4DCCPEQ3SPi6Gto9zbOnKALPH/q+RfC3UpMsVzuy4cwJrlFy5FTVxqv
VnCV6hPb07Jd4aW7484BJ7eE+Hsh4yhV13UlcULYIebxsMrtXwz5OStl5AjVnGg5
/DlFS71E0jFVR9T4ETNO1xFJP6p5hw6JwS269d2Ffsg0/vflhef24gC5YFC+63G0
Cq1dGWidNV7TboLK0/yke8+021+TX1lGox3IYFqBW+rmjcjKcN6wZvB9GSHFQId9
MV1/zqN7YZOamh+ZNHTZ/Hd05RcNZjgr1Nx4dJ/qL8jQPj9uQ7pN1GGdhEhELwzZ
MrsQTiU0XV+PVB7nov6I6ip3meOegTESDxZfQWg4z5DxRewX0sh9WWfbjrnvgY/0
6eu4OzsDbehagU9FSQntsKdYyLibHkFs8qxK5Caj04rNUSywTK5GI0ueL0CYxDva
TbSr1Zaipiekl9Bt6yvnseBC1+i1SdUjVciCxTGVclK2AYvQa2nXFcmbrT077IlJ
c6KcFGS2vfWfpAt2Qs2GrkEIZJUwZZ+kASK5nVGjyvUD6wa/n6glXKgu6CMciL7W
1qOFupk0JhvTPkz7yb/4mqhnPEt1ZneeJ+CBSKT5z9P+JwVn2Za5rA4bIZk2Tp8a
8rtmiDQQ7VfySaEx9UemfREVQD5MbjkM/95Uqs/C7IKlZFWZKsUB+j6FbZ7z0oio
3wRWJ8BhSikJ6Js5dQdQwHGjQaEXvNwNcJToiTJB+vsPi5G1aphXhYb+1VdFX+bM
I6HgHie6Oq6H9m3w/epa7a5Kyd0hwrqJUIa4rs2iEr8332LS1xoMSOXPtXnQo5Ay
KyptVPGSmf0NbQzm7rUeeEtHQ6ClARcrgw9j6JY8+y1w+Q/CrMZRtqhRQZAFuMnR
KPNqx8I1g3E52ODTHURvytTjh9iQKnZCiHF//NQuxv7XhgcnjTOMW2uAny+Q9wO6
gXkrEzThQzntBNLEJUnHaLiFjgFuzHFCBYwqJz9VIKHHHQzfIu4knXO2MO0IkJtf
7N5Zlo8I/fEdFSsDt8cSF1nnk0QGj1WdiSDvPbsr8pS4FuA74rtc8Wx2WGhAinby
0aPmGOe+tbeV7vSYZDDVw5rudWhH4w8NCXZxkJloxy+MqkmVlsqamijy3kQSc8Xa
Y5F9HQrQesX5+TlCbHe1JBQODvjcO9rc/GqMxGtH6wHaCBp8JHmdr2Ag5g/lGeY1
Uwt48saZUjbPJpYUhVQSZ6j1AtWCAApfmVn7PUdFca9gD6D31EBwaZsnqj0AS8HI
BZxqqCOz3Kvi7TvV04jDoAHWgBGf3JMZpZs4YGYN6LydJaO5YkPGd5iCKQ03i7xs
uThDMsmGNR18cxtNpcZ4WqSUSiE5D1hEDjJM01NOx8M7XQgsb8eLkFbbawC4JwWm
h5jTdReqyEJVqOChF4RjfsEfZGdUrKAusD46pAi+f0qF9aE6UFcUmqVnv7fLjm/c
kFEce/xkD7j1UZT6Kv5VzK44nxplHsqc83jrPiPJKUxPI6mUH3xsKdVvIU6Qm6RE
tJ+c02Tv6ZYpgy070yLKGLG4IpQ8YuFV1AF3ioVSbMAwnlHB8t5Oa6RrU2d7/NxW
sfEih6WdwzsUdEcHzRW7ELsG5PDGNRqetM9VktgGoYS4/IL9jbH9uHwACYY7WgSU
j7u8TFSx+aXqXeC4JvzVsPu75mH/jtD/wCjXkFBHuD+d43cFknZ624MFm1Sw7r2N
JTZ4AcTdxWYbjHKz1VBOn99bJ74AgcWLAJkSF/W3k7QLsKuGp6agQ/9a026hLW5z
hiMDJhYCycnluQSyLvKdsk6LpSqApNift7/O8FcMzJFSQOBmrdZ8EMEZ5NHvAvtL
bb75S6GAg6C2ma4yaR+M6UqelYXsSh+z8wcd4XR7VERAsVBr9c9W2uueF1o2DhIn
qCFlNrXHqLeh5wieBLLNFEIHkQzTrcyWcMZJdG5IZeysoy1v9t1sKAjbU0QGUmr/
AkNgqpmV0kgHTRuF+1FPJPNNLZKlkHpFIls6WqKO16kbbZiD8U3IFFFiQ3RsQOqg
1hHER1zOTP15BaSKwzFW+GAe4GnUdyra6RQ/dQfI6dvBeHpoYW17BvC+nqmOiI0J
oB77HQrHAKgwGi+UbYjgGOVWmGOiqjmH/gqJGeMhUrD0oFEXtIQgdUTmzCxEhvrs
9EH2SGBpHG9HfAO5rph/VV8T5l5vHkMAs/3UYx70JYeD3Oa0gdGJ4YKpsKPlIubM
FBk323UQiQSbOU+sqGdNYWxY1edWvooCZQF6S8A64EJcRvU5KGWIZMAtVwFHMKwn
2mtbuSCzeMO1PoF/Q9PhWPHCzfNELB19qpyuBMnHpX3xSDMOMHGIDck5G+uYLrq5
xoOzkfQTUX1pL62KFq34+POq7NwsayIplsYBxSxTwY83O030He8Ie1oqJZtldcA8
T8XwgfI5aUkrOsKOxsJGhQtxr3dFyhTMX1o+yf0cFmlJpe/mTsfpnyEf4qVQGIdA
tAM1ycENY6Qxh9QhLpA4aP/ewAO9j0XRKjqbX+L7IKcqEyKzIHIYLuHPhXzjXyjt
eEHQxcfoO8ZL2iIHkeAflvFyDMq6egAQ4xwhLbNKD4bPeep02srwKvaLGduZbSnd
Dfo0aR+ZSa43Iogv8SV5GV80T24o5Ugetmdd/DuQLw3Y/7izlhcmjVz6QX96ZMz3
dCFJzbcm+EVA9dxChJkPL1ee/tRz2P47jqxh6oQCbg/vY+5bmxM4UkbB5nZvZNXp
Of+vGtTD7PZAEPPAju6J6pbmPlxw88tOv4QdiuEeG2R58/tpEtzCKno1aHbn1Sj2
0npyBbf3WkWPBP54MRqkCX57KSN6msj7Cq28uR+NMQ75/BLbbqdGn0dUNoykfwyt
UbSaz2u2TthLYOTyGPN1vxQpVitohLWQJmjSJ1T3xi/nBI7t5wYtG/pUI2hJpOmb
KPBi7GvjKijE6nPXZk3CMu84yr9SVn5skyRMyXHscN43ITS6zYicCqo/pdETN7G3
GnXQg1sK0YeHvLc4DxE3Cx91irxbhY3lv1o45niTLNX3R2RRQcbR+Cafwdv97AFJ
x3DcVVZ1Re0vaFTPvQB2DrpXmrwSCzsojq7t6aQrAx0gvIaBjF1kO4aS1RjrJDdS
at86dSDBpF1jog7YDTyQcmvDiPjS8KV44GuVGQMQ82gXbmDu8vqeWU7i7FnK0MYP
ttnrJqwEQ4YnNQ2bmgMnI3GltRm3bE7OLhpBQDJe88fDZ+6oGp3QIvJBSYkmKcvX
D6Q/STLZ3ei/gw1tCpS+inxAdXUu3TUqloATRI+QBKWNzO8erjx3p4bcRZxKuzuv
z4WQzFbQowAGu9G3L9ydjpR6MLiqO5fpcIaC+5ftjVmm4xYRicDGJkt3DeQBFhwv
4aKAjVUOJYk2TTSeNiz/LaAlsiwi8Fogo21MMmsmX3F0Iw3hlxg0zrxOXzOg6iHK
S1K07F8iIYfXkR1tpc5E0kMVkCrE/aaDELjm4RacowKnb0Op30je1K8CIXB4FeUs
pYQQSrKuoN5ODjPTXN6Wgs44dx+rM7q0QbymEYXgKiUrZ/9vbH3uuxoqwdgDMA67
7pA5a2a0Za6ftcP5RDHTmhSow3r7cUYRrixpjmqyLugJQhIIc2qaICCe+njdCsiB
hQ+lcJ1mmEpiNEgHq9ODMmWJpHQhdThBOQXLekIwJk9kEzBMBX5GIpGB6OeQFUHc
8VkDBMHefb+jANE98yjj73WbmMdQBRppo5g2wal/mVLF2BelpXWVLNq1g4UWrxC/
nkLX6C23HGaEe41kzV1+qVzu67vjbXTVBrjWBn2AltynsOegdCqbserOqrowc8LH
KVKRmtVFMO+ecLpqUZoHlpqyopgmGjewJNHLE+2ostAVtaLPGcG+x41cwIiiDzQH
AspBSCEi00/QgKncjpgRd1QpbQTC3iUfuSmuUkNJUGcirUBP4eHBdmil/GqYFbH9
CFBzScAKCZsUHx6LM8GEEhCHgH7wT3g6iivodR+35J+FjDBPSsbxY4Z6X11L8Zy3
+FTjtguFy2WibgUz0HbwSdrACFpA4zeetgMW6NQhfXjvj4eb9R5EjsiWjKE38QYz
4wOhXkWuRtuTUTg+oxJqqDiMATVpBgP3PvrgX2cT5HVT0WJjCOwBj8XzaGgg/BAu
nfTuqRE2HQnTTz7hSiGm1P4kuGNdSJLHa5n7afWetRSCmt+9xXvABjh5YJifdTH1
Hj02JUAHEeirAg/uluEvTnD8olUPhL0SshgpxjVUGC2Lkk5octpvlqzN/J7D4Mue
1ZNUUfaoWhjh5vcNO+XDLFhrc9vLyRZrAMim8S7/FjLO9C+eYphtnLbAKmDjlhw6
yNo7L/C7+BC4NpIbTB+4SwYN0u3Y72WfqB9yygCrTMOkIleUP6OCEgWmAC1OMEMK
v2hqG/ANrc8AyDypUaCBxdETvqDrVXwqLn6Wm3OBWSWGlRa4pA6VNhNlglEQBwLj
N4dBfZ56wtVR0aA3p6ns2VeHCyvakvRWk4dh9eS78oeJ/T9+/CdoJqvnop8k6aQV
dqITieIOFnWj+olAISopqn5SObC/y3+s7Tujivosl2KVbpIzA9/qytcCMSWN/LHc
b2yGjovYLplxa81fPh0MRHhURegDJKdXLGpIr9cEEFMsOF5G76iuLb0N6XMiitby
Bhps9AyuB5swpjxzJmWhIOpCSNUpk5AVeLMvCTbnFfieevrkZnn+QFyDoC8rYE1j
QTJxNOX2Hkr0J2/cIamUHJHbGDEWYkaoSR/cgQ/jlYUrzAnrXn649iuapBMxvDDs
MDXxay9bM3QaqfwFapKfy3ZHeYriLst8N3hxxjef7zqoDW0a5QvItaRBdxQLy7fk
1FI4gI+n0/SIa1PToZisjV74F4dsgFB1ojlp7qUdPyKZU+N8Dv73zI9vrS1kkpZz
2xt7P7XKL4eDW/YV/bOmYW8o6bs9b5cYrzHGZ5TCQePwV8yPKh8ceyUosEA4qinZ
pLRDEbYNiecU11gVRNlf40aFNo+v9+98zUmW98WZepivEwuf71dP9TYZej1qESlv
ZzyCoSAR4VonkgSdX6J9HwfSTTXsDYLEhQhBbib7iBqp8t5tXM9f26JA4BcIBi1d
iU4x9+XXLuh99Ihy8AdF/GTwOWqjfWTKkimC9ZqFDj9U98XBgDxUrejs8nUP1oJ3
0KPb3qgNwY1I+q4qdoRKgrzZkAomdJ8VcXH4Tf6zD6l1Y/dVDhPMlNSLSSYf7xBk
9hlFVZw/AuAMUIrInnRXTKGQqmjTnxciUpYYw3sBb51dOzP5V7tarW9vk5qoQMbe
SOQOtVHSJF7PEC95/rnvuAbwszHwYOfXaU+k0TiLRidUNUVRakr+jM1bfF+vQOQm
RRh3CMDxP5EYCWuzvGi8crkFFE9Ag5/H7SkA0xaYXfTOLY2PdAbtYpnSQQ/J+ubq
6LMS6UGemGqL0D7+syJmWM8I9pI/pRlvM9vxbMbBmAqgjDeJPeDay7ZlOrhgc1Rc
b648IX8tr0nc+rLElMxUeTB90DGnUm8xm0wfPqw/yosvdfx2+mZDGduu2dsZHMR8
FBqeep6/feuP/nz8LYke6cewDwHm12wc0pOBmgg0S5UekVfIKN5F3kE7LyigrNWF
Mb+PDRA6R4pnNed6W8/P9tUtevmtuPfX9T2kzVRvJOE+41eEyCtzm4sA7kClDpC3
ZIJkngYExVl+yhj2BVSBTwO6Iu7IODTBzGNcRlI05JxvStCH4/WqrCjJG8Aw+g+L
g7RecCexfF+OC/UWxucM1jDzkw9xqp0DxOgO46vQFHbE8Fa20kiZNRtzRjh3ODSJ
CM0i/44Ls65oFH9wE2lETZ7y06i+1v4OZniA/OU4YC0RwK1KY54L5c0pWyNmZEnv
c8aU67h8FGJKc4ouPQCsMT04LGw3WzaYrE/OgMkeaHapWsJTLGFu1cAphVP8tMjp
OcC23Z8bjztBWYlLMY1e+kxpqzQL3HdkOBOAXLe6BO4pqnyNpLxxsVQJu4L3CwOW
FNr4hfIMu0ezqwgttioPYEbYyum4NzO+u+lRVJNxQCd5XWj29dHAhNdcOV4IHpoF
RuM+2Xcmf0LJZUui5Ugfrik8wymmbVCY9pP92mtaSkBfu/K8TJcnx3jln6ps0PEw
JgWTliJp4p4E4e0CWR9VkyoHTqOvMeYclKQSpQz0N6alMjQeW3f/LDYggAMJD9Pr
Wh8+m2+AUrJOaOxuKfDbG6aP+QPDOAT85LcTbjIDLHZyfqRun61dE/iNCpDMqbCI
8VJa/vHEBVIOWrZOkDIlIKeBrfJ7KTJUNWF74PZovngVVsagDTwncs0mUBfw5M0g
DlxBHOw3JpbPc6vAB8m6urSk96E43oczunGe/osM1ROOXYBIucbGpU5g3pDblOlu
3K/jDfNjmtMMHmGqSa9kzow1eLO6Gt+KKWJkA7NggigrpSpyxjPNZE3ExQY74rmU
xl1NLfhiPzTO81h9/6nbLWW3gYPqEtsd7n3tMdCl8a9/4TyqriaRsSt3FH+e/JBk
bFLS1qcT0I/qifyxPuOpsYhyI0dqCf+xsfxSL6YhTBrbBxpyMVmSVV7s+Zr8SXGW
gng22dHigeAEs/hVlfhXCIIIwQTf1WmHwAEsfyTVxFLPRuSlHtWf5/BL04D8+kU/
MGlSzwWpGD2bVd7/USqAGwgB5IwE5kEf4mQzF1OzyL2Lni3vdw1bjtYiXhHf3y9O
L/Ni1FfXfm9H+sNHVgOrB56i49RReWduH3eS/OBRmasxsrWFyVMAQfwE0v9jKwMH
pPTgsY8kU87LEfhp/kT9FkGXaeOdqeOHc/L0fR/AXwMhHWsEFUFssv3Ezt6Nt2YY
R29GHXjw9/3XM1JGokQfwSRTYXQlrYpJ97uVzoj68usYr8Y7xeE8KMNQxbQUQ00c
srtRR5DISQQ1Evm4YDOwpVGiqfXd2/fdgdePI+kyIFEYf0zU93AfToGs41bb5uIi
iNz2WTJCzYM9xmCv7wNeIAjYx83xnbImRjL+ucRhr1u9earYZNWcREIEW9Coj09h
tdOxjpY6WX7e1RllC/7YY3RW/jktMMdnAyJyE33X4erk3vJB7dWADQesVQKIXBy0
q65tsH4iHTFiSVTDcHaVg83POpjmhLZekDBlJglW7oDReswQlGUXC1iT5f7e+Xud
YNgZD68dLrRnCPyjAybnxe6FweBliBrv7YKmo41aEjVw13+tXOQBsNdauvRu9jK4
HdMFQTQ00MMICUVScgiBUXugDLsF9F2UD9GcYkDhLH/xVmOiTjOpy+eO3Qo4oxhn
RzYavXHIkLZil6DqRVjzxiZhG0vrj41GhXZXJ2iimG438UXLN+axSVV/6/xNP9GN
t9ZSD7i3nGXQ7tbtz6jxIArkH5ili3f1KBQCAadkut+WkwVBFH+SPp0CMrn2BD71
uUsdP3xy9IcN0Fkr8cq54DPMCPWVrumz+KlSaxApA7yGzmZ0IZZoCa4I107iIOAe
5pWjIfLKjNg9OG0IggneVcLiZuKuGW8qRoutJtZeJ4UV5Qdpw7XRlIZ6eBrJseVx
QeblDecLWIc/DhbR9ZuGKOFtwUQpB3nt+w94OQAkKxvC0HuSGYtRdCbAh8nfScya
6/3H6FYf30QT1B5YCoDfV3QxtbGxYVPO6TJ8Sv9mhdgw8N5niJiBjm/RQ8MY1myA
UMx1pSrNWshX1uyN8pOB47DcQj2n1uqzHoXjDYFu8KNgzQrFvMxZ82dv2Kriizzj
0QYRJM2kBV32gL601I2PRDdEFcoiXRALI6UrERjBoNeQSFjP/pt6/OAIKNXjm/Xv
iW9Shtvk0YUcPO0ALauzu1kBBt1jyEYCgerVi2WbgftwPs06LuLOUI257eT7rs7Q
S9PuflIfF6UmNdaXOqoZ8f7pNCtbdwgmsNkbsd0N8oZQTckN16YQmVxQATC2zL6I
gJGaO4x14kufnF8Qd3hefmi+KKsPwPegCub0K2Gt0DIWSpzEmteGofXkyo+MITzv
qBqtp5rSHBEBGInntdagNPAp7i2tckL0dIiZ8gqAdwI3KN0NpFIRixIt0rCKvoVO
Rfl2iqy5OFLMPuhjwUyrLXJin2GdowFC8ByG5axCWPggdsa0yNXqGfmTzzCbkL9g
dFKcgwrpgpUkQLr4/gvYU/ACb07qoAqV0ilDBUE4AEm0aHUbGcbyulDdMWISIUU7
JAl8xRjkeDbmVFmdFCNAM/e/cqcIjEkV5/0UZY6aKbZhnl+HEerKtbEUc0MerThh
jnyVrNwBF1cGmVqjUFQPyrLQc7iEazbFDVOqsFoUWcK1ZxKEUuZrIPLexZ/NR53S
ZOlM52Y6Dkg1JunlaGPBNTL02Mrx3/qewdcDJGOwh7HyX05Ll0/G3MyZAuBrL17I
tmJXu2QSIUgcMOTDO4C64EYzPy6g9SqMT/oO0vh2HqG+ZLLEDJYduQxX2csccdbE
+THQBj6LWHeV+QSwGNIbsdLemZJyumnG7dkWoWVeHeDBOonjaSwtedMzuStqTEy6
aCJVeQWvP243mgjq5DI656q5YR7kWkzeSStMSRwblv+qU6IKVlJ7380e0wG0LlA7
wP3GoFQVWaRLKUqp8/kzoNumJEO3I564gFjfiSNGhLxmce1yTjDxTaQFNPw84Zj1
Z44DqjX0anX+ShjiojVnklASUL+Gyciu7d7BSebekoarV/14CX3Ugh4ne61syCX0
mNrPwYEZdoCEPFz3nnZDYYXG19/RJDRDGcppB7F9ZlW5NXRqt5EZrWATIm97fn2S
r9yoVkzA8x+hp5il1lmJUK4wy0PYpDVnx8UNDf1iyROOJd21bQZM3kXlYN8MVAAg
pAK4gQ5c3db8TDNjsQChxyTG05g7Nsg4UQY5LCfLmX0vXdovckWXdkJOQci1eS62
aWJPAGPpH8AzdevEue2PZmAXAmFuWsbxvS+dpP6zvrKczoLLbMlyuPIb5UA7Yqhl
1KG5ulmpOPVBobsV8gBCesDxMR9bJsRl1uLBIOrGenZGZ7a7RoBsfVMF+cDr1lS1
KUnG3qX28/xhy35Z+7KjSg/BoAise687SPa7XP9Jl4GUWfVcf8VAZWUs4Z8KjQrt
Dbxj1BwCBrzW1cAa5erq6/yJkv5G4n5V2KMxibTTir8bkuhqCl/RLVHbg9ypatLT
i8QQqRfx5zrgRjwOCozInwYONDeOZKuFhZ7Vphq+b46kmEHzTCj/ClOgFPOUNaAQ
IhMpSJR5XKVXWOrVdyGQFyfPfYrHOLj5hQ2/2eAEOqRY33mZlYviU8ZAV3pMS0qG
ycOsCI2ekkHPc+soZuVLed17DGee6aycFDvJyZnGRG/k4bTw6yE/e+N3afe7lpD+
VFKfgZAw02bMXsHwPCpB+c/6EZyA8dEJns+VpOWI5nYU1iVnqou0qwD9YpOPq8ah
nmT/6xYBuSbxN2bJV8MhFwFbET3WeI6u0qSSwq9iQpRY92GY+OXEEzRwd6Bb5IvF
abhJ1uVkK3V/BAMNXtHGa5btpTgLc0KWgvZSkNfYAr5dBEa2yVbKvLdirJBq7cpZ
tkJ5zANTIsjWtwHkZKWoAadIhwcLZ1Vj5xA9v5s2STMISLxl7WAMMQie+wp6ZLia
aY0NKJgbUmLkD4WegAe7Fv7T4ytkdwTtAIMzZ3rEab5yHVZ2CUjR8Y63r7QoYJJc
5hM3SqLv2GqjEIK1nT0OTLBCBbYABCs4+lzO6ehn5q+6RRI7mj4LDHzTHeVnoUWa
DZQN7Fmyh8AFkpRmdoAudik9LGXUcRvnX1MXlUleUm5gpqNMuFFV9CiuACkZ3qBz
Kejn6K/1nPA08PIi/U7xFtd2PuAo3e3tuhol9WUxFEAN4pydFvOPblmser/2KJ1U
ZkZpb3lBta3/pyrXJZeJPIyttnyZ/GB4vaBxaTEXKer1JHLR+ohB3uzX6IhBh7sO
3y+rMKuH+nbTtntCegg0lCEW6jDA3xjHAq1myFwSmj7zJyC1AvHsiHMRGgLn2xfM
jBAmgrnP1f8qm8jrfnzurayxDSh5S4+arSpwl0dolKxpCLi5UdyrvOjj6BcEJ/vG
E4B0So7PkOOziovPO8eMkI9ZioDnbSFI/K65FdVGvJt9FlVkZAuKv6iJfYOiH8ag
DWbAo7OF9YRee32n7XkJDljKHU6Y+X2RyMM9FrSk1TxyxNb/MbXqh7Bci8ObSh9G
ObdMZKHQDMP3GtROgId0ELkdDloItIWko/dnUECa2y48gAWIoZiqVEFegk1huKts
yzYx5XoSZcwoD4BbBev3nK5wz8htsSABVKyNnv5swQTKz+KpdE/4bvAkqKXjLL8J
EgKExnN8lJNGhT9X9DWBqfpZSX3cPRZO9c+I7NAiYBxRZPcTXINX85uct6K8uWZT
onyf1KEIEqtHTBfMKRCTAge1m38EShV60JdVX6rXp4/Ac4HrlATtjkTETweyI/xv
sSVdg4FsY1mrbm716w5KY3uUYhuzJHkYkDuX3XK/PTY3wNoOTmNQ15SAcbTOy1Rb
pxNco3/Npw1FDOjR+5KsVsA6MzfkWkIipzOQqR686PKnzF4i0vCweEAooL0HDlTl
DrBhW/As3JF4OdMTHnE9Zs9afEGacGc2EIq83VX/0g8CU08momeKIKxI5HKT3XSh
CJEUUv0e4WRmWpT1ltmLrxcCms9YKogAzEw6pJprqxZGd4bDB38NHaBPMKodYppR
kboJLB0qXyYqtnjjTKZmPCtJ47GlbrgdfFtz9b2uDgFYSiWCPCAPzCAtPF4JLb8Z
J2icvqXaNZ6Zpz+VxYQFJ87687qCEaySIkv+b7nC23GTS3EKs5GD2ixNkahr/NY5
X52PfwpPPzDTn+X4/ucvVTfjzgU+dTNM+76SyexP4uZBCOMAHFOJ4YNBUj8gUIt4
KbHkREdlLSQdNkhmOtzmOfEwD977oEQ5mux2BPrcbN6eNHzKUQrfGcUIGQrIspZM
GgjzXlWp3PCsuTbN0Q+sc5l5IE0QN6Wz1lFy86uuGLBoPghDwTsKXi2zBzuPLsDb
fGXhv1BnA78+iw+nUpHCTgtJFDWgcZlx2BWwYcNLiyy+dDjcADRDmga/AloPZ1NL
k7+JhLk3ATsY5cv1xHht2TOF8CwOdIt5VaWOkak7RkxVlij8oFnmffAqd0/se/n6
kCZsIG3r3XW2/f2DYMh1hzI8zuArcb+W66Z9nN6zQXpIx23a+WUMsSyA8RDMBzUr
LN9ivvxIWdTn/WO99puFHSEsE1RgnagGdErfE1/AkiDsWzzuOFkirSrkqgbf3eBV
9Ez3YM+eL70ePYzZgimv+OxJ+EssIvxR+GE1RufvTIK/K/9iz4pYbSkUAmaco6Nr
J4TFC353UlKUg3NemxH116OwwenY5XwZU5SusYZkx9KC8jt8GNvxuNeykGAXtYbr
Ogmr6U4k3Higay2I3p8MtLai1D8eG6cNY3ShvJJSZYkdOTqnJsBgTSlGUEVLCBDP
z/mk2LRHQI/QSfZH0yCM3cDak2AJTOo8QTEGhkQ3Bt///wetquWgp9eouS82fwds
/XjZOjoKSddpx1ebVvfmVRCOLJBklq6yiN/p0Vb7jqXUqHr4QC4hnDke5GCscOkf
yDe/48o373x6WmikpXAmypvolHHZp5M7JSPB/ohdU//hs+ZGOwfAlM4AUUSRTCAo
Is6YXsfOemLqowe+3HNiRiLFlK300OziywG6xr3qeo+mo5q+Na5hRNaEwOLTF+LC
O7Z3gAkUKOurclemRp6XG/EikJ4ig8wtOpySiuUS8SvQxDyeHlgUYgrxbIMxPn4l
ipLVZ6YSDbS5GnxHu5kq6WWbF9WPrhFV1yX5zluXaUVZVGTVWlaa1ZxXOC2+K8Cw
UIN2fERDiCXejrmVpd7gpeuFwdL/hJR0YDi9KJ5xJn7VMipiKWRVTbp41Tfzc40l
MXlMjNOERpAHbfzW3mXvLM+1MW1re93vHauokV0UVteJ+d9yEKQb7cuXre0UtsKQ
64VnvaSKK83wwUzISEDlI0R4Ix0iim6P8dGjQH6InztLBhcRynVU8/yqCAil4ZbG
X+JayYaADAv8WzAiOTukVJe3TDUUN1TbgAV4VIV1/f/05rVUMe5ehsS+94l7yQM0
b2KWWQKdnj9PYZ3OIl8eabZRDHUkCm8Y2P1CCspEe0IiX/DbhikvOW+bae47X3/x
i/ljbiJRSanj/UeYWvLWrKj+dd/lFq+BbMrJcaP4Uy0sOKYufKjXzWYBLO8Jq8D/
Eb0Orejn+MSBbVfuYc99ybo33iJveHy/UwXD/eGkHqBox+MDr0SUmz1pSI9hIip7
wO9dJcYjZSvqgfmlxf0L3paLvYB48LvIQWFOiXhncZGNEQ87cyWb37xO80ydZpVK
Mzz3uVKuxICBF4EgFvtE6/fWV/B5ZYWnt6/fFEa2CJepL0b1lIH6m0QkmjVxyHpF
H50Z+veoSFMEIZFPU0ARSdIrRKtUs29AuQPX4Cp1I+I/VxTGwY1KbO+IoF45BD+0
/uteKFjW7pbbmoZp5rELvEA8BrpMBYVUSPTZoetzZoIbgLaQ9ylPesk7IhPc84Ca
vWSlmmo4O+EKyLxpKKO/hUrmy3BTpoVsLdVKjON7JvW20Kc8ZPe1GxqgaNpt/nVn
gxxhrFtxJtiAzLY2V9W9gVvYo8iBrZk5Yc96PWNL8B21IPqVaaTMxbzp9vBKcCSG
WeOk4yv9VRZzxP/eEf4iGvK2jPYq03v6DR221O+FEnYnQNPPune3cvrYY4/mhoHc
rvZh0pjqViK8mviuRUaTBoZWSSZgAZJmlNx6btpY8QSsfiirwlr+YZ+mWhCX9Ez3
VVw4xHH868Guh1Qz/sJmWyVxLaorm+DKypTerZNJWHbLWXF96nJQTmcR9l56QjF5
KOaUfz7O60oLvcS63G+D9TRWVxCoNt6cKVTJMYglk5zt7QMpGUaZcGsa7nHXlOSF
g8GUD7/sPYGlTeAc4Ha04x4511g/0j+gl8whKE+iIjpjuNJeVUsjZFZ3Jo7YwPIC
TmRYJZziFTMnTLjWrAsC3CMZqX4jIKcmF8k4S7VnJ1GHJEfTTK0iZQ4VPC5MXa+z
MGpaM737GgERaLvfPH5aO72hPuwxJJeOvm7ZOFPwinusWBQ1fsNLd8DycWvy+8CP
czlw1o0h/ggNnxXY+sJXYJQViuUFwxmxuaB96lqNcA4rbnYJPXsDM1oGzGXVYOug
cn2G8Uwj+qaWSIegXhQcv7fXKxDUO2+3dWUeSFQvEROXXU3k/TxLPSc8pTS+l52i
9LElOkGqqEgVkU472CEKiqYlVKThmgLah6+UqWx4I/FEp041o4WJ3FLjmEul9hKe
EJHXeeRDJD6QXI+wzt4DRTBdon45IIIM1rbEYtHWg/p0CE4nTZTcqXBj5QeMYrBG
fxmSdTtvjSyP0wcFTkZsLvLDA+uFgatfshgL8t1B5iXf0gsiadIGEk3cy48tWHST
WO/cMo/FBUeSm1k44PpCjxeiQm4UgrPKp5jC/2SAOELNFoYP7IT4f0XaP/GcfeMF
jv4qKnTUXtomjVQJm7qtUXGtz2yxldxSDXoqmfMq9yILACGv84Ikj3CGHiuFlaCz
+OMDvYPzP7NTxKuwhXzDYbt/FUquSU7xXPBn/murXwespKiuWAObK6EHOK/msu09
w319o+ko4QMTvpjCfkERDIB8CbF7QtwDC69Wx3xm3kUgIvY3ySv39XIn3kUyKt5Y
KSZqxHSdUxpbY6EB/Z5BXsDPQGn6SsfnfaP6JISZ5BZWHqH824/5mGMvt1vvKm7t
KpEasLLYXcDPGjrrg+29nV96bado6+86hAJkpcHdRtdFxP4oI8UkUF/wzjqgHIpr
hX1Yi9y6JpxI2ZuiZy/WX/m4yDwBRBgwQEoHU8GNf/y0N2qopaVVSwjvg8pbLfRs
fz0807bFXosm9FfhmVvePBQAWgmLVL8DtG/EiZ3lNYRNsmaJ5f6uu4Pth7QbS0up
KXIE4nO7kHUpUR5txFTCdmtcTZ7ofW/vQmJQ6mU1p04NrL9HSZKXe3im3ddobK2k
yFPym/4RrUOBtzPg7CySmBhPrxMLwfgsnEsMQYveXIUvFUdo4yQAXvcEFhe1a7Iu
I4xvzET0N1QWCtcQxRCoRVsrQZh9VIi6/VCfXwla2tAnsaUWjl8SdGv7HwPk0hGQ
v4LppbqaGKdRp0AAXBn4b3u7E4myUOZMqGfc38hvXpJ4qKXGDB27i7rjlySrvVnm
ouDQbS2a3OFH5eZvYIjexHsRqrbHlaHPwJpHkjMO/T7eKfmsoQ3FWyUu2OCWYYVb
x2fgSDdDda+mQfX5+UI+GG5T8XFpphUJM+VrjIBGlsdVsx6hJFJKwt8ptYdm4e9l
nsHQI5a5E0pC0/huy83CgBMeIN8UDa67pWCC8B6ewtJGa/PopT6oLJM2LHMiOWie
Td4B2PB9DP2DPrsjAI1nQfUpa/1GR1pryjgGDR7cUoyn92bHMXEmMgAtHJDMYQo4
VNSiTiJzNFyJ/NnXMAISJS/WSLnpnTwbeFP779q6l0cRIGD3z2aPMeuMwdaIBTmj
fQdOfRFUqYGDWAOALSBmnaXec615UcursAIknoUZQ/ThM3M4QeGMiw7VWx+FSNHr
CoA19m7eGAPUWBxCFs6gqxnTBrEXruHtmmBcB0mSiVJjQ9da74ZYnXinj4yDBulg
//FNLTBzDNH8nv7ZLNpa8hnorb8GaTcV6rvW6gAn2NcgcaEObOCbY6uCLJNPW3rT
YOlRc/5EL4njxkZ08cJZ78iWWmcUfLc9MOm/zGCJsMsQ/Bb71F31st0pzem2kn77
p+V+VATLMkX7ySDwAi8TdX/h1227LV9/nuUX7TwBgRXZkWerGwu4hNMQC76CUFH9
MO0Zo7Kq042pxWh7GAGAYOeXGhFx6u8LIj0MZfpdFztmiToshq0SA0D8hE2E3ptn
WYFaxUBpQ5l0lupuXnBMuzeZOqVokHGIqNlenMlrxguYNe9pGXEYm2jsIIIcJ1US
FIb/zVbWx44SoW/LsWEqCpwRUTAcXUilXbVGtEvpEo3sdUqSFwTO4snaunUXdxfK
01dJxGrTApj/hwKLP80KjWR9mtLL815NZpujuLTphfYKru+K1XS8LHGcO5BaRdmV
gEKsYgazJqJJQTNviRljpUvheeYv8wiDCfdoQDwBk46Fn4N4CXRkbNGk2tWhH+Z7
3uPQCxTuHKUwTCaZsF9nReI0o7Vca4U44FWjVqiis6eltMUhTOwJzl2MFBHKYU1m
xA356ElV/ADm+Ccc+rTyAQQbrL9x6JS4H+QFjmgHjhS9uJxQKr4rswvegtzN71bn
ICBCTAyb3T1hWNPxKIng0fZayVgnZjC0hDdUwYlHsdXn/joB4/xRbVlPHkJsqeYO
S2DVminNkyrJ4dwgg4jtogp+CHInwAdQTEmpEC+R+Xk09g+wGqIagLNQmJA9KJV6
+D+17yhooDSyPScsHy0LEmEiUuJsPkZDIj1DwWh19a31F8AExMCXAZUwVHYGNUJD
UlJedd+P6uO7lW1CV8x3xAZZCvHlYNl8oB36GhoAcdnrz+Qmqvg2CXtBaTpi+5pA
H8bofJA06obIi8XvMlCCSDrb6okq0Kay9U8KO+dWHPpk88NYTCFTx4nn9uWsK6hA
b87K7gGNicJ9r8ilpgNYGEvlux7YhlIMhhHmVK1W+qf33E/jeVdESx4EWcaIcWe9
FiDyiBrT2jb0118M/hVKqXgcwt5bNkwF9Y52rwA/pGIbpU6gYq1BlSHio7En6XI4
795d9jMSpJHF2C1cx5cBUNBBnbU5S7QQwXnQ7JhNcfoIaCBjJdejT3wgxG8Zgukw
Gb+/Slty1bLHPx0uZ/Hsmm1Pm9oVhjc8mqXvsrJWgYabaFeyAMZvryI2NSwZyv8f
C9q06CmdRB9j/AoeT29wcyZDSl4W6qkeLoZ39Du/XEwQIG2W9u8OxIIvIAveQdQu
GD795uaJX2tRW20Oq1dMcmWODUe6j/OaB039wN0tPi0yll16y0N3VKUGGWfROrEH
aYOUvVUyfiBYwSN9HpTNS++ua3eb8ks5IiqTIOueuWbPwE4tWFemY5CgolXfVpv2
gCy9+9hWaSREqlQ23crILtLQUJi1g0+HtOvYeHlGnMoEzEKBoXMQPTDkhU42lrc0
1bkFq354Esi/iV+mYvevV05J/h2UCAEdCU1tKz5iEqJbhhQu5F8LxhL17HL6Hi/l
Yn0Zv8has7zUQ/P3EdPQELlghcz6hURmbQtG0fiaPW9kV6ULS9BGrZir0Ws6zi46
f8CZEOR5qF9bh+0nGk6VWGHQBIZ2BVYz0g0shW/PlnygwKEC21Git6p068I3q929
vzRbiyKAYEtFlcf6lfaTkhf8VlJpICEmvzhkQY3i3RqJNQ3+LbmruvCiP6l2v36C
g2Ail8QJ5CQKQc5Gzk7wKl33+vNJMWniZFUrcUY1OwZGZ2rJ9csBLMirbvMalX28
ISJ+EM35hZqBC7pRfJITWn5HW0y0WrUsy+3qpwtrljL+Bo5mHPD78p+Gn05xS5T6
u2nRb855uIyheSTjtxJIrc30qUHjxvmJnSRQmMo3E60Ju15CVrmM4eJvoqwwSTKL
bYbJEKsD7NUwiMhdIV4Q0QUFMLajiiUTngDr/HdAWJi2EI09vBDnprx8EVgFMyxu
BWNx8kraJAyI4kO+HRcRwYfSlVmO9USEHZtxF0S1qkNTwOipTRinSJJyRywEDn51
pbizhqyK4RMkSlyAA8Xxk0eZdNYxuYkB33OOIlw1AdfR7TmhLnOvy1Bg4qdJ12qf
Juss6foRHoKMbhZ77zx+WS5S71zUkR9CnIwevEotg3XoHQzC4ZLTaZDu+JMIuH7M
GRjvB4vZVERD3Cv9/NEFwFJZr+44T84PqHYecc1MJMnv4rhte3lLzbQ1SZkTb9k4
ojrVkK0aZ7n7a3JWry7zuLU8d4MHyeUU2mQISl1i9M53FJKs1vqLuhBdZwhDUVd2
FfrB4JoVSx9RfCTPJbX1cMoQNiBMZux5dKyb7QV4TaYNwB8JMAuif1Fpww7EC+ti
SNvkHYFUZeB5SMabvfQdYhTTxWjL0WLGWa01YvjNSYeohCT6Mn1z9WhoFaUTyaFt
ZYvvYk7AxvtiEpL/Ns3nmv7KMkC9YbpGV12/mM7fVP9Vai51oNMtWbkvXNVI3wAn
JxxDp1E0n2nbLwz+/FeRRrzP3+DVPBwG9R+yRR0xnxexdGveHjm74okku3PuDulM
P4cNE1PS+pjkZoA7FYp4TTflKulCVDHLzfmrkQEJLcTCSkvywIRRu0hdERyNqTdl
Y/JiOUw/jce3LiTJ+1cwxaHJb+6megwQ7bq3uGfkWJx9rOXoWF/tOFCkkUiZyuJe
+gSpCvc6mKiPPuPrRYCt5l8ok1PXeJpzZ77Y12iuCDKX1nUbG/6NU4/GCT4JFqeT
HCC3irafsLPXgsd1HZj/5CdHh1zgJoNUIKTT/sVYjxrziRccqh28x5aNIM61OT8v
q6061ncDObBMz73hjLjzYsu9pvhkB53PKPO/VmcNk57qrKHE1TyDZa2QZp7YLYvs
QvRVGLI9l1kkcdz6tzZaUBQzRzgTh/RVHypbbW31ajxTN7XmAOjknNyu7UhFYzbW
Yf+YA6xB5of2DVELazZM756Nf6CfSavvbiKBP9MXRhSF202pSyxXLoGEUbDhHt4A
nejzwLSBwZTvEawYenkGLuPFWzugILsQ/0EQ7y2TE6Y6Ys/wq2XQz6DHZ4NI9AlM
3WLN4MOTCIe+8JBO+yCvZObzhSy0w5Y9xDeUjZJvrzS/HOjwZIpqHptfmNavREKg
hh0qpkD03lk2ReOBXSco03/FbzEBKnlk2KRPbqpdnPyjeUGLenrC0+P9mElvsjOS
mWx5xyvBcdDCTijAN5bzQbMU639MTp4LAheUSRkuiDrMxdqWWqBmYytzrmA73Oac
MRocWOm+zjuwCYlqvnJTj7q9nzR9HtdNDY231US+shlhOHjQB2lPgFPIaDwl3PSR
xugK+yZfraihAacj6lhQaC8zF9kgdme1R4hmpBsQVQ1yT/J0ScOTlH6J7I39+3jg
nrUualDQV9XpoqJWzGFS1I60N1dRQ6BKJauYdgABC0WssvPuIqon2DVSvACmV+W9
2BAJIA3pwNz3GLeB/ttrWWvLm7Jz0wWjfp78KoAPSqhEI0rG8k2o/OmfE+wr9I+E
3dJX/DLgwnyxjBSzSQlD1/oHYyP+Il6TuBJhUnRPmmKOKxFwgT9RZbFbfjDOYo6x
Yq1WKsYm3oeLWZCyFAi0bu8U1YavGlfdgqqf+dcgktDg6aJQGYENMBA3vEumdXS0
qjYOV5g1SuMB53sJQPlBVznsiCatiSKFAtoELF3x/7NpCy2zlUe9S9Fr4CcjrWhc
gPJVTX8BY7tB3WLtcQhNabSzvcUhjKO76YRhjJBeONforJ2pTYDbQ1w8VsT8fjQU
8NPB9fQkXUdHlZMKXQl7OISYA7zVgklWR/aQgWIhAE8FzOxEqS8MoiX8dl+5Y3v0
ZQHn6aU5LY1lbJDAiF5EYG1m1KlZDVERoUzMeIVgTgQ3YF6rj4bXEiv85jTKCmc0
Kbq2gy0YWtAKIiCUiPCpW6rJVKsbNTEapn7URcynMjdp17jRvBeArgy3DqmDXi9M
/wVttkz6KpWQat9l8aNUpWXxtISuoduhensxVUKsJWCVV1W0BadP+MV74TDDEUiM
dyoLPKj4BjwkTQ+MvHx/YxhPYUxYDznjZCFj0dhDLfIC79zk09rt1Oj9+zJ4RV/l
idql2by1q8+UH1x8kj8fWVuOrSzJqcATdzjE9EzmbRiZwv3AmMA/glZlRubZMaU5
gdWDv1AQhbGnyDjYzPiFVMOW4FH8Ph8puMdJaicyoaE+LWVjxkVSf7rLHYrghbRu
GULs5QFrTLo7ljWyJTzGLOCKUg64W+MUhuWFacvTtPk7XxPQOeNEMFLNU1M1NQY8
UMjiUQTlKfp72NJuyyYpOgycauBnJtEiSi9daFEANXj+tx5GAxv2B5dC3PDzffRe
xpoMQZJMr3hQh094a4l+JyGxsubsNtxj0akgWYliYLukHQ8/B+31xNGx+TnVhWd2
7rhHxy5vlwpZ1TT01fx0NhSyDmDH+hu+ynUm6MxJnolNO33z2PTUtVd+gTGhNb0x
HUCEbxyTh8SalfrcslqkdnltRXsE90YNl17aRZqw8RV+J0j+vJ+JtJSOYbFnY3zw
IleHvGXn+UizqV63m+022LPqMzZfjeP8rHMYrcNx8ool7GuhXFQS1UAi5//Ti0Zh
P+y6qc5Vp0cQGnELBFCm+MEKBXhOMsrtOpVDxiFhDJ/SuFDyAa0swoOoaVJfhEYm
vWTwlZ6PXyIO0U4cF/7DJK4JWXeaN+aA7b1/ooGWeXmNWmPgwJNxIy2ITmc1ESuF
5ofVg2dUuBeQFvD2HbrDPeG2n16WKiYm1E3yiew3GL2rf+cI2vF1gQn7kZqD/xUj
E5pM8oFxeIqcdjoQDlGCWSZyNdmT1zcnYCL1KuF9ug+VM1JW59E7aKPnPL/qp1Fv
LQlrjURqnmcouIwXK4UXpvMKvXRf8bey4YNiBZm5o9o5jZThf23d8za7sp6mErjM
8Fzm8EmrOj078Eh5UFm6co+MR55UVhwvYQkFs/9Izd79HJDcrfNcVIrahCtEsElZ
xwugvzoPkOJjDuOPUXCV57O6rlUS8oN6OKPGGy5b4xxGvpco7fLCdWQs1YUYhziF
40eCdgSjaHIeoMPG3EpSu3mSHhJvXtYIHg8clN8KvgW/fjg/PCDvIUl+CD9X9n7+
VzqQ5QSvd6p2vvSc5o3pzsDSsGi3ldVx7bo6zbR6SD7YeJ5uwzoEASb8mJTBrOa0
P68/TpFh/99lE9Sq+QULAURUR1TOqX8DKxTa7nlXGsvHX4Wch8G9h5QrOLb4M1x5
Nz/9thPLfZ/ZfKdK0I7MGykC7erUTfT1RR6/0zRSoQLm3/ZV6P12fD/Wq/CrpG1z
lgfObcQAQxDUhxPvmV+9agWfW1MLmnJD5mYvHHEfoWMQmMAnNplOBhYn31aFyMuw
z7UfEtPTHFFyumGw37PBCOGiVJqrLte+2nMdXeXCbzMXRm4cVxeaf+u55uZo5yEM
nDY5DUryfIX2fOF19BgBQYTsJbzeVGDPPsXwhtS1TQHTIU5YYKW5NOHxArslxEX/
NL2R1+xaOF4FFVmKStDTT1lnia0up48JqZTHV9ALK8dJuPKliyTZebMRrgDlkpOk
yLZW0UKDYmAk1yY2Hiys/WM3HTd/zm6zUpPQZwugIyoV3i6YWc9f7wKi+lQGKu8S
PX6bwErNX238+9vbKfZik+PMr0NgPw98DzSP95VAuDLZ/Z1+J5/NEZlYfmkIyEMa
XAPYSfRbt+THiddGVQGpcmVbg6dxlrLs7V5LWRTPGvabz2cXsAXRibWI12OOttHC
a3pt/6daiN3EsT8sknZCeEvYbKedpE+soJCDPG3A5bTmJPSFGAv8IPljdEiTZ0ar
F5W6s+HqorYfCqmI8FuyIY0zPCbSLVOnI1+wNHwy6VMDp0PjFY9/GSKgIpzlnmyU
/hRqoBctaze/WwuBQFZ44chux7NhPXHz7OlowN1Dd9PE3Ijt8LvSCO4Ld1D5VXot
jqBbBgFeV0Dm0aHl4hbZHaFeswTxw06hnymRlsEFsO+n9eWXz6xGzy86ShKd0gkJ
mh/T7cUdiC3NrTw6xcELvchj78a3oNpNCEJgyr8mvoZe5PzhMGckqbA00692JBDg
v2CFVfsqF1UOdmRCt13CHIQC8hItGrvHNdqJSGYWNDUq3L7P0j2YQisVQODTklKr
w4eCNFVhexsx2Zhp/4Gw20QQKr/Xykf5vl6RTYSCvRnPLHPlaVYgHuGKv8HTEnoy
VQme74oLcZ12uTqiGjbAg1qg9HN8bEfUYdTC/G7+YqJZQwaF/r8OiMhzdHBvYwFq
7bdJBdvBdMukxfGGM3Uc5U1TAlG7A/vCUlf6p1+mjJa8Ah5rPLsjruEVhqRgF74J
ORk9YYU9+f8N1ZMga349/PxvHi7zq2EEY+gCCK2x9DYP9AfLH99pVGtZaDAHsJH3
lKlO8D0yEzyL9W0NC+Qi62le6WYFfaEteRF8hl//1JV6FtKis4VYO6TaiGlMMSSD
RgqOa5BC66tC8ceWUxhHAmusQs2hnJw15lzVK+EE/vIAMfN/idLMZkl85i+5iA6x
2fCYdmTdLWTFRbZkL9h0TdK4nvajqO079DI9RwVI3KAfPHQbzZ/42XjcAs/G5FP3
ZAAy4+wW/YKarhTPdvtZbSgp4fXYFV3sWEWdXTSv+DjPS6WZOudVD9Qd4jALdNsO
9PdDmyuuWQvJNtS9YC4aZSh7iRqG160mE2QzJhgOaAqRuVMShjCnSVRYRFWyYp9t
ZnHb8GjXLo+SoJ6wp66xwVjLAT9adRXOnCfGPPmJfzgMJ5WPB8m+8UHNzOJBZGsd
NsJigDdW2VaA0m4Ecto2a5NgQRouZSJosdxe+UHrdnlBqu4XzB1qKVLoy0X2+RNO
mY8dxUXyf3GCZKnl2pUiybOZshW1ypVGytf7ZffaeEIBiUU6sSpHfj+SKfR2d8Wc
qZ8gT36Of8Mr/sP7igp/y0pa+ZAITbRddLln6OZC3gHSZuDmrX6UbtZ8N6RXFSD3
GcClZmUmh7Lo2B7+S+ZISVAw0EtgMQwHPV6RL+gNtfnvQUSvr3pqRxZ/Rtzr2wQh
sCo5TI8PK3Vgi3cE0OOkLaB7ObN4cAZeMQ6tKBZsiH00ntKRDKuWUx2idVhMojmm
o01vZ5+mfoB2acgu60MmiSRu/YZJo5VVFJGsaPA9+EpupyahozL/qYvHG4wvPACB
mt+3NSwbrjJ+ld1DXkv2yCJJhbTSuGjAOP4Qy2z2azKKA8XYmHbmrWWEBTToKCM+
h/FZh1DdvS2qcwdT56za+k9/UaOvWriNClS00cvsH3gLSu4J/UIR+ETxGW8rAZf6
W/v/MkImmm2szLBhBpOBOobCtfQ1i/DJIjL2tuQRzTnypFI+GMMdq7p7eVvmwjdZ
B28oUlcUcMrSOr0AWOpkd5Vj+FDjnNvpY26ANK6rb/4R+2szUJ7UtXzB2b0TIQhp
uWxgTUMYjeCB7aCuHKt2Lq02giS9cljFk7M1o+uxHJF4OJOl0HtQclHFDCX94I0p
qUbtXWdzAXOFVd2K8aK6bbranDjaYxs9WHYOpASvQqmdPqRP8foZf+v50FZC4fkS
cZ/u98Px0IEwzz6hemOH0m+vGHIxO+N++u/Wh9wtZyOPIUlUPiQjiP5NGHKX9Oec
S/d4V+oMNb40nJa5hKwwlTfVMGg20lqprmSdJxt0hbUZDPEXmgX96OtrpvNSzx/a
cOwpoXSn1NejUcko8Gf/JjPIbQKc8cxvErRPHO6o/veDegLvDuL46iRhg2gIuRyH
3Yjuqx31LBtawDaDisDmDEME3WpSRTCTshKoMaNfneVy0YVJtsHWvVj1Ankn60Pv
eIc+Y0wlxJoOKY0Y/xSvuOL9m55IlaXNSaYkSedVjjxA7VYGhXAv5Afu1b0MXEou
YnKtchipXh5EPCN91P/iPPTnqTn+pHzVmQY9g+Un9LvRwj7LFHbFGCfsaXPUty3I
kDIa8FSS+k2/OrN+WzYlYm8HCJxAJEbkV+1tcN/yRolev0yZTWIIFwGH044alVJl
5Wv7Sz8s9/dVQliwnVIEh+coblnzpDNJuNVRTzF8+E9WJkWqCngDWxdAFuGpVeqc
kwQIhCyYJ87Cqp0Vf1hU3qz+kdS3c3kbo/gHWkfl8/7DReV12V3Oij/OeHjb4Kbs
lvFj40n4PbQLHEGg8hbhFAixSJLQm5bn9JJNR1i5r9UCatSrtBE9o7aCOtbyWt0Z
GPjrYg/Y0tSjUs9wtNirdFVNMAWwDw0CdNimAVWosualcfhIVRAT82OPj4G1fVXb
MadLL8ySqG4AjckuV0Uh0nv/0EXy4rw9ojW827EVo2zk8Cxhxf2NsroL9BeEdVQS
2fgH71pAWqrulx1rJuH0TflcHEOxeQNhd0KBZaiV99CsYHBxDAJTaajGvJpwb8ry
0GgV+j250sUFiRJ4QjuKZnIxOq6Lk1A8JxSjF7FI7nWbTBpHA+IKnSZtES0Eee+k
C+ImlFITa2rnyAqAvZ5s1dGHZ3uwk66a0zmxfD2J1OZQSUHYk1E5yuPqiBPP/eZI
eXpho+vSxmaOFMymIfdDsG+wnLzMFdYz+z0vtZZaycjS+rZId0MgRMBLEiUIu/BH
djUdhPYaSaA/FGwxYrvX31FMkEEQIYTxIHp6OTi4Ogo6knjoSa6s6bq/Hfi0oCi+
vUT2q5CxVtTBgnBRra0nC+b5njQ4ay5xDWMCKsrmAq3ZYaohvH1eURcj0EZs98lw
PDV30USDJZ6YTX93nZfKWN0BTFRQavhWZj853elF71rED9D9gaXJdMZzmxhwp4Ns
VXzLiQP/GX3WRq1an3K7cAwE+uMKayGPcWCHb3EN0ELbWr+r+0MvHjnhyQWB+Vmb
SfI6H4IK+tWU3TQ8IGfMYnqqhWmS4r6tSsYrB+nluXInWaGDw5khqwIVS2flr8EE
DhdQa+IrnykmpMePrdYhK26d4AudCJCnUmmsW0RuAxqFC19zb+ZyyFEMliPGwWB8
01uv+6dTT0SxiUceTneXY4C5QbxTmOMZ5y1GORiDGxPv5geTxM6+ATC1VpFyk2si
dMo21ydW8ksGm/AUjuLeb7dswQFRwF53C8q2ruzugVj9RvtAOMoGBGhT76Q10NtQ
Kw8PlbWMWtj4dJCkkUay+4KwNi488fPT55bdlGU19Yw08LK/fW6HCuPe0cfVuqBU
T/XwW8q/7DdA1RBgnin23mCeGPczfJVn4eh0hduWYVjyeijQhvbvaBLuf4t/1fvA
M0zdfsghAh7ZnsgqfdCV/oOC2XbJSH2uSW3xWrZ7P7ETyNi5szIBrA+Ozu0rlNLW
hWRTp3gAbyjio2zKp0JPxPk1Me+rA/ijqoksdMHZhys478ZjhUNCMvyFn7cXoWUR
n/HgjDwgaTTDtmKy3abXm00SXqoeQmc/nKMdDOGpbkdZ4aucqckuQK3+8bQkh/is
rN0qWf327Hd3oHKiXRrGGqYmqU9LbOg8BjNFAJi88WCBE4wfLtiSMnjuObTNh2s6
PcOxPQcLpdJyEoQvtRSsUzdKca+ZKxeXWzl/FlovLmAKCClW3ZNTtjJwVPwgp/tF
us6PuDp61JPywJH8MfNBZj46bGrLUdIMZDci3hmdzFiq0KrvzktHJtjwWhKDYI5x
BAbe3fq995RNzjANvRM/UBumB2n1rJCHrrLKv+piuUdpLUKdvGuZPK6bFLZroHKK
k6N4Lbmz7dncIFnoCQgn73r+axsG4Qf5/ag6z3GrUDYf4BhvOExwyg6pFs03knB8
hr8dr0xagc8j4rFTqMLTqBPuSqmqU/R7NYEXETdsmDvGNuQaC1wlRIIx3FcM0TrL
k2GnmsP9h807EF9HzKVwmvfN8Hj59DFJFumhoy/F4eVZH6WooQJB9Ws53DhHCZ+w
reAByB2KBy1ZOXQNX3QMnGUJ1lA92V2lFlHoQSVJGDH51RlbQ3/Wgs5ksR2q75nq
brckjwgHVIzq4YcqI+8J0VcnygLvMpebPRWeb9B+ZNPee9GJrqCk7BO4kjyMB9lk
/ybScq+a4QM+60dHRW95J8HdVC+bnYGSF+HZhJkFhPaTm/ksPVo7uOVcoQER1wXj
iMirBpKOoRG2qZAn8bv7Tao5BRIXATwjI/wE9HdCT0MD59zhyowxUs+YwnP5+6rA
qB+hLyPHjEE4zuzqi9g8+KL/jRTA8e2vY4a/XsZCTjLqzYHNzrZ4yrr15r645Th5
fWwk5Vwg8t0zgKsDbsJNO+P78U4pNbSI7wV2B2ZsdDSDJdFQspQNQtws/YcfO5ru
F8jVuxkpB2xp92Dj2dA+zW3/sw5CnvfxyBVYBUka+w3IiZX+eKBCwBglqr3m7gTk
7GuSKypB2v+uCIg9UA4nLd61tDlNGS1k7wyY30XuvorXvKi6nqCohp527ajnWiL8
pyUmzUqBY1W/NmjHMZ9myxDjJZIo+EWUS6VIGxNu22Y5Hy1DXP2cdlgTd5Yv/nb7
PMG1GdR6ThW40pNhCb0zsUoYarRMLhdAHDBerGy8mSPPB/xPgQYZexXVK7RC/G+n
f3jJqxZoMMGUmiYzxcEKszMOoN+WfeEXUjsYw3ha5h5yQgkjbu6FJaE8MRwWkyUR
wveaB7Dm/ankE6JU+2e1fIwqBZKmU5bEhvXUhr4lBaiCKWkPAfS/byD01uGMOc10
AvxrHVffFH8Rsk4aDlueEEdRSPvZ8rQVFHp0c6B5zQlVdytQg3exwEeGQ0+aPoyl
H2PSF87u8sQjWBixURXWm2XYVM2LWrjsrGM0Yq45uoYYgGxYmo8vwjS12bC9D3Kb
r8/Ir562CjYWH7K9Eb5qCxINBhdZIrfKSdhfEWTWUDVwwihxSTWWrhIksRMk2qg5
nexaMshcWWgmsMXUJ4N4d+WgSOjq2qFQlVpIH7jLySs7hUDCGmAoSlyO18ZPSbp7
aBaodJ8rZT2aVa60gtuWdEJmsLgTvbjD6WuwHyXyqlOvsYTrXIMyNypZZ0KhVZ+0
D3O99vGtqDuwl6Sd/AMBXctp6sdeYgPpvJPNbkFLU1dCQ7vLp8It6St+4+KFejPP
e1skm4oXeTrBzReglaAeu84ns8qer6hCGXqkMesTKwmXKi4K+1IwUxxLCOGiiJiD
Sf2m+3eKAJkoCccuXYh/QjwvOKAFVXDnNnnQEGWf01j7RCTqXGjfkWXueNmLprnn
Yh6XJoJtmsC/MqcZ8laTwJlnA2qsn2MWh3BTb2auFHjM9+OdT3REnn4jDkxrnWcY
pMMzdisypqgjXvV34efn1Ec4HqGpJmd8ymnvOlQhVPa4LlrotTX5g100NwzCtHze
lsuClGsCzATfDJGVlRE/gPVhlWWuI6AB68HzCnWs7s3ytQiSPE+WJ6P6SfylevQd
UXhgoACQezI0/QctulC/MuwJDynGWEcbP/oAetkXnhKwr6CE6cU9eWZp2n7ESKAk
9neiMYHhrm1JTiaOH4Wmqf8WiarzGLyceG4X1RMJwx7GHgdoDyYLoguQvgHaeCHO
8Xy3EUnVGfGG+dKlc/5g56bvzYSuYpKh+lzqrfPHJcCbyLVEQOm3PWVaZfZogczT
B4U/ErRsCd7kaqtE6S9w92x/XToEFdrFEBbaNcYXrQvzInTt1CIK/z0R5t22hcqd
sil4qJGcNpnq/tSI86yqOv5uOuHFrHkqTG/JM8sOLicCVML7FsiojzDHJMHHs0W9
kkoqQLJeNVOlMwBj0yzalR/XdnbkN94AvFFFEpgqgMXWvDDSEHNe+CCJXCiWL4R7
jZFq52w3qBxHcxo5yDvRjRrKV3T0xZluvGyGufcDZ3fPtBH9ugRsU6R8PxnRn6Qr
4m6G2ibwAAn4frJhHGQ+3bxT8HYqnW3zSV0vfWe04sFbOpMc4tY35IVLMe7rJkUj
RkNuV7FFQAuxTt/tudVfqiTm+H1QLP5Dx6Qxghl5E0q65dsfu9O7YtvnTixm2Xqr
HsTFEgi4TH8Ts58O+xKlF2b4gjiiSsBeNkvOIYGcsCGy1Bu/FW2DgeJYEojmZdod
DS/YQGTOmu2hu/ex7w63CpE3wnmvTfk6lWvINh1TbsEbQwgZP0k67b6lmhGYplQ4
DLMspBDhyjsn3nkWMHGk9AnH3GtwIKWPstKccNwLH7D/pUOAAFa7qbLW2paVzH8x
zpFEyd7PQtV0YlFjzh4IVkuDAVF8Axx3wyJ+AdZQuaZMVq85SEI5TjF5NMI/RPMB
CS63f+titr5Tn1S3hUGGLU/Q/CBSd6flmo6lmRLD+ETJuY8me2SBUPiM/dpgmoFJ
6we6BwJ2HVwS1GDSnwDGmtI1GTSyXFVEGjJwKHS0zCWQx4yrbGWYxGd97tnlyeZZ
jdITdA43LV7T1FQCMvGBt1ThSewSU5GVKb8hS/cj+mFopoWXBgq8ImRkTIvn1Nfc
iFwOMBhMt5lsnXZOOCwPtZCgC+kbwdvUVrq+FuzBq/HNE/cfXWAf4Tev2rKsdvXA
8m6XsRDqtmnPDWQyKPtDOijQwTliwLmJuTqHnEtTgbcLlBklWHw4X/QSAgxZBrCF
NBxJ1B+npVtSBAjcOPfOLTREL2vdn9u3+/HuXLfFEzi/GkWgDXgnNZvsJcEbSRka
wY0jsO1U7e85KmhXXQFGGCIYREDtUcjA0a6fvl2ta8iVRP3//89BO+jWDtnaRWk7
4jLoej1eLib9sMV7jnvGnNw0k/rAHgSHfwv4EYBw64j0BYUW+1PsNYEUWTQaA1KE
zhIv9isj0cTfNplzFgK37/8bOBWKyzF9uRoSQcPzFjAfxjW/eYASuj37t7nUvNOt
I+8CDdUM4Ph++SRy/cOGkTd4aZ0k7S+Z5qmcFYh/HVlQulJmIskYoFK1wMUUOxVi
/ka1NZ9m/bsXWOeWKdXtHDKt0tvURWYJZfcGZNtaVsmUwgp6OGJfhiTOh5IJvWIc
0UuCJyBb8M+micH8fre6Lla3Vj7IdFIwUgrp9q2jjuIj/KLPvopH36b5SjBQ2JeW
363MHRHNA9xkB/BmQBJFJrNCVupgsEfvMqb/n3v9b66gOcs/90V9PUqYYEFCgf5n
IgrM3jdFu/upPcwAXxsYSzrcurAez3DjM4FyybBNgo0KmzYcjfr1BO9TSJI/W02U
s/pwCD4XAUIrcXcvHPV/K46rsE6+eFALCwyHG8Zoy6/TTz/dlXUvNuRPpOB+GYid
751XYUCzWwIrUut3PmEU+OrlU5XstggYjxZvFLpAnOt08Yul53u2nWXssjarCIzg
/RRu1CPzLOGjzUBy1gC9nBQBBHypw1QTspqcayhlkySbJgOH/md07RQpwAtPnxgk
MFGZxnfnRviaqzoII99kMhaGeTO914Ln4qlfmDIBVqLX1e+rbOR8M4MwAEMlVjKf
4SKtxwWjBZQqpXNuZAa9NCJ9p5F/+i4hU05luceB4EH5l/y9bwcDl5MGfGMPWFKm
U290VFIcWq3eh2fh8Hrdja1kVuB+hXqRpQUCMfnnRDECS/KFQmMyiERobK4ImO0k
mwUTjZJEbaEDO4O2QRfkWOqsG0Axog2hiTPT7l4/F4LyEcg6ww19CIDlAm+Z5/hd
W3grzxKOPT0th9O46D/W14QuosBX+mWNMI0nnD8L98GEQxgPkCAtVcO9o1ZxTMKN
RWz52+CFN0MbPpmjZbK2dHvu7WfKWp2yxG2TZYiUxKIuHiMXNegE3oAxwMu6ySaH
YMipJDF8jFuZaxk4228D+aE04+UvFs7rRmPYmQBGy3yKVSR+on8/PZpBCbvmADRe
iVSbUDok/3dj5pr3S+GP+VSj8BALeM5xPrHVITOXVTto10PtswcGuz0V8CJanRO1
f2LwJit6Idff874OO6nywXjxKLlSsAmBJaVU5jvTvKnO7elPaE4KLHraPDp3dkVx
dp4+iKuTXV9cIV/ubRMeOkh7drUzyvczd5o0syEWajdjH6IIBZ+R9X93SXJgfVbk
2VsmJmifDHpuXXAnzI1BS0zxLQJ9EGBf8c26O1TDt3XonH6UTr5MI0VvESEgGkwq
AG63tn+AJfS0lsq74AgV3F9lmm+PUTAs1efeKvqb/BGLETWO4CMMV38azFViCDfR
7GoPAbKUSzL0lbHU2zigHPNm2Wa6/pF5wO7hYOz1XnxKctOdXQKE1D0rzegcORDS
YVV8vdpHo5iOfKCSNdOiyiPHdBsZjaa9qn7O6U64pPuWfQhKwTGxM2qFkARu7xgQ
zoRdWtE7RRRLBtPI1INnKRK9w7214tO5G4ESlvPbQ4j+vB/9lRjsA/iD2aNssFsx
FTlmcg9uM3KHJkwGvlJlOLnVKTBXCQlX4U0EP31F9W1j8N+5WzzHYmoH6cyOEwpG
PmWZajd2jYNs7+0GPB50iyXB+fNqXMSEeykdD3QN6/sp7fstghKh5WGWv/97ONLG
8D1p41Y4E5QLfWrg6jSYDOSJqNqp2d102XZ3NUgFG8wqlxOaek3AdeZySdCSd2EL
IWMUd3HAYHQfHFLrGSrgn2ibvnCbTdUw5HRspMg+0pM5LBvSGPDjSXYk8/S2dQo/
akRrdva0fe2eHnHDNEf1yD6Q3xP+mHwPpozA9g91+fFyfCvZcqXaszT0Rf9GULah
gNBHFSzlGy9U7f6wf2+6ttuiW8MNq9yfTCM4CZpsklVaqcP0G9ZERNR7NrJCVIvh
j8LHmShEngOBIBJlyTD0LGudXw5VruOquoFey7nzi96sPAIrELQW069HnyLiUgTx
rXVrsxMTcj/egg6X8FSaFKKEsP5CPPTBjyG2OmEdT2M7HW/58gJe8c5ud3GcuJMB
wcPltiVbu+Drj2rRfcSeJgsFq43KV1DXfvkjF8UrH+Aalg8fbFQgSZ06xwIS1psZ
HS9X2Tx+X715nob0uPMxI2bHjbPSk83CjcxHArICsOcOOl6kxrx1vjiio2ewSs7p
BTqSPOIDfTgfqj4ie0JfEH+bf4MmRGEukFzGpcakMPZXaQJsjF3tIS2TzLbNnqcb
/Zjcf7T9ORme5tGGZTDBepwj9HJVT7LtUrddr+oB4wrQG9b1BStLONsVELUfEzdb
MyfVK6qdcSNTbnKnLWmMfOdkftnpGxqVeesyzT5dm/GpFBs1zMZYA3NEudDzzpxh
lOwsQrxMqV7oAddZvPQm2exHJ0YNvZXP8sJ9GsyTyFjSLkBrVUi9Q0mhK+O56HfC
vuA3s65hk1r8ESSXG/tRnX62IoFz/iF6u+R/aUeTB32LINqAMPhFzs223ByukvQ8
qFSeXVzEnovbkXVi7AGm1VKs9IN7P3iLb03oAhj1dfGMDlbgii1BBcTJOU65PyIP
899zz1vTprV0EYIzRy/RL3HHlkNiFEJ2vO9dX8yYB0F0ckLx04kuSeatZUquRzPl
x1NV6HBKV0z4lo3lNoziboyQk2jBsUQ5vL8qqbHgr/WJdH/O3TFbFiaxYfCz1DAM
aS6h+1Jsh4X7/ELngKWEQMrdtydlBGnVUs3zOi+Mz1kNYeQ5dKy4vFQYrNBc1UuW
KZDfSg/yw+IO3o346k4gUxhyp2q2PJlC67m25/1JbKtfBOGPPBPW5Krc39aTACpy
dgfkVjj39hFwzFiHtXRm6atFJwvyFwDMjk5X/0UR2M/kVcmy5A84ID7LGtYIGG7g
v3BU/L91fuXzPnu8Ufu4E/EfSoM04Tg3xRRH7ABk4pL30txMaef93rP6nqzRVfY3
ldO5FJz493hvSOwNZM8lUb3khmvxJBV5RdPQRPWVnKgUqohgpn7Rcv0ok+IsuFaG
Xz3VO8VO/zilw5EV/bIOgl7/D4gaaEQYDecipWqL/3mxy+Gz29sImwfGk1JxoA0/
u4+/sfUEl880LpZZ783NC0c5byISbNBWQnpcov4b1WzNzW5TOkyOZiXtt0rJwf4B
Wv8BsssP3il/c9MpW7cmVntMZuA3XAL8qvR3oTc4WHLwaIG2/rMuiCR0SKuwdtVS
4JAl44BfQz+ACJWoaGbh/vmM6HOTcRlX4LlF9ttqORt1w8b28cZv6AeH7TKBNeJx
YdpRCNBHDxLq2z+c8HU61YL5EJGMOEn9rrJoH/XSxKVhFPnrcHX6Taii8Hb2C57z
WlDDY6RAlgGs9LJL8Jojx4x/uLDOTkmZ1HX9VYZWjNiDM+4dcAO6TCZByaJHqzpY
KocqepQNfnkpR6iE7JGZY3guPRfLT+mNu2PEB+dEAszaYexffUqtCc+/hT09BkI+
j4gvJ/70Gin0oLIcGR04o8s7TPD0rCG4aqRz3dCpcqlwTmWAo7H8bQUYkl65MpIS
Va1yR+RNblrmTtGmBGHReuG4NkHWzzRM9GBBVH4VU9Q6gZYLreDD7gGnTxuGLiD9
lPwN/oWtSAPRcYQl79WQmrLwwMmJPdwynJqmfzPkppvwi7LMzsrJTRG+FTf963Ld
MInqg0LNoP1CQEMOIdukboHy6BjVS4+GTJVNqcWL7EL+KQOfQHgv25nQtqMy5uZG
FAvpxE4tEGmutX5xabVptFKV5tH2SHv8mk8QSMy6SiPuQCq5aqQEUaxycxLT9mUj
USfde16b1MiAQaiwl/lDMsmuxFuTv5fcHS+8W7HbiU5HrHcNbIzbYqAuxtY5nxyV
SUc9zBzXzpUNmyUyT99CBXMe/2nArkmwz5/GdagPb+OZ5ODXm7jFm9s9NtC7iJ1K
SQaphYku4ZAqYTJAXe2g8BBWjNSnA5VUz89gatUeMRResYeKWkgSAz5n6OP5AeQ3
phvFEL9Kcf0IIF809rxcma70bEJZKrlNb8gWV/XnNe11YxivsownMKsc9lNaMcET
1d2AQDDsXYw/7isIPdMnyWDO/faCVEbqJyRlx/Zl0RWpqVIjawxnE/RY111JFgkX
8k6Yff8v4Uxl0Vba9jc7DNYALhEst0L8yvcm2Iut5KKW0fDo+W2ilHRjzzi1Ep+I
EjW6C/HWgBgZeSZKk1AIQ9PIvYS3MpdB511E9Mn67rRyu2s9vvj+3s5LscAJaO6m
pxTeZnkS2SII6AliwOhWSXl0ZUnC+Jz+NXrpLYrHmDQLrUhwifEMTk8W8oSwvuq1
VDQM1B4MFNHy8hUiAK6XVzoBn/PSgiYKkXMym200hwS3lro7w2dOHKDGfry9nOoL
gCa8fadoR6dQTAZQbxFlcW3MlmKhqGPjJ4Y8Ok9y6iO3nZVLcRvXx7UNlCuEY0sV
sNiH1wVb3cgw2d2NyJlH+eZuy4/ccqcNghDQZsr8qO/7FMevpAWSTDX6ZAKOCkXA
v2GrpLIESvBp/EYDqL+w0mx1LYgYbT3LvfXoYyAwxUDS6E8CU9RwkguyPa1p4Ds1
M7eApb3XF3TjzrUrEffSjIFBuVXt6iVWpVK13eboNtLDAuw0gcjz1AHgAnf9m9p9
TraOUdkGMgNSejXBrmrVlshj75HPh42doVdtdLPWArOEvl/eEyOxPnSBol2j2SbN
ivN6FAs3M7XDmMb9ZmD30pUEzJpsUWXXmKhMKJhAe4zmeQjVMFkHwNwc6op5pFTt
6X4MSnR8tOF7OzunKyP/iZlcQDOJjCXc7VzFp7Fs+Z1Cy/RRRMR3OUreFb74L0qm
u6EbnisZSBeze0mzzkaW5NP7Z4ls4XsLw13m26t9XziMvuUPSiCYqBYQ4pKqx1fI
kFchnV75E+8STXbsx++rgXch8oqh9kaA8DZj3Dc/Bu7gcYU0GOaI3jhviSrPVv0i
e5EcoFvPsY+LPCWrqSA3/hk8Ozw3Di0rYcZVtDLJphNsULysSOC2rm0Ty/rbvf0s
pQuRR9fBHJNxAQ34M4IDgsrx1O8UUBIN6wi168/5J5ILwCgz0u3UVq7NKKF8/PMj
pIoI6Bp+G4kt/W8WpimSaxOgs6fSo04KbPefoVIpiQTe8ShjRFxcAKgCTuZVzP4Y
LKOxGm2JoxSNWgafK5b0g6WqnT3eh8SrSpO3kJ9XL6XD3TGNEhOR4w0m4LpyDs0M
fN1hFRPST3WqBjFwXxOflk7hrtH6MwUoqvKxO/7OLhHxzNTvoy+Tt34gWSLHOCq2
FiOLBUnntvj9c1W7Nhz7z0BKSEJGsLnZEa+mKKiGJL+kRovKHTwHe0FQYL1VUNAs
bWxZmej9dOhFrZTVRSRxsKDV4RcimGXBqwkt7cdQHHEMNE2ZZdUDTBL6pwHjwNeP
NGilvHhbj3Da1jqRzPtRCWxrBdP+rGO3KixVXfDzbDQS8Lkkv+Ljiw8kFOWwqSK+
89Z4QSX8JgYTK0QuUf9vr7ytU1nBXkFpjVBroID0fWw61+uNG/+tgnV64ynUnTCE
U/dIB5FHLoDaYOSkhOLJSd84ooJAet+uGOXf2cb7PjYNYR45+woWVjZkHM4Epfg+
tEbDNf6OboS4n6SjSTzutCpHRV8auU2Yf7I5t2RKYDadrGqQD3Td93K6YRwZWYms
/vxZjP0C7raRwzdvT4tFeJj0d/qYSeDjbhyNggUHSFV/QgfzlfsRbddixEjG8qTE
stUNmf7fsFA9/QfwAAdxfXpUMXorYpXTxYrPjR0RP9BW+mWReIuPvCkQ6HbB4UUC
ymsf8ZpV6qrAayH92cCm1NNtIUhBEvpw0+iR/OBMozYpdELpB+jbhiqtnuLRBL+j
+c2g0nVlbTByZM12Ajlf9jN8xoYMdGphGceAhelZ1PkIzdRZdEe94Ehwu/0nCCZ9
mreJXX4N8IcsHcaZS0LFfSG6qXusr4QIoEjz3zHx++6hhQTq6r/hhCqNZayVUSHW
UHit40yL77S+krbDUFXj/5x2UlO+Q5t14PloBebZj4QkQPPRZkKT7x1CsVyVd6xc
0NwqLtXJQK6nTRu+19Zas6g5BT4Qzj5q9gYMBzS9/K2h7ht2RBO3GB3xGmE1hYYP
m9SDpJuLH76V6rrLIj1fAn1KEpt2/RQMJi2xUkCob4klqcxMAUkw0GYBPSvFmjP9
Zqrm0569zCS4TD8ELDnWT13wAOM8q2f7Gbszl4M9dDMP19OzYgcQFJqWJBDshUl0
yLHB4ok4FZzyuBGRC6I+JntFls0Ppw1gQoV5QPMVlBzw3Dy/FyEJsKjUtm25Hmz6
5AFovkbg1w1PbEjCDCMUbkS3FsKquuu//DQgdu3zvmyiEgkkkEJZhM5tjB5OEgxF
CA1BTbyGWK6+w8Vh+k+C3gOui+tLgWGc9MYEMT4KUDUinxZKc0n+TwgfZ6xdUQ9W
Fg8VgTCsp8ozGlPix3FJNzeLRE9UFN8Fu6uzigTHNUaCiLzGA6iVnLtYHSKoQBvA
I0E/867m1BOsos5wqN0BX6ASMieTceYlK2hfefjMAbOY67hPOGD72A/6MtoNCl/D
wEbdS+ba2McQuzDRuY4cFfxbWwo1A0yzawZScF5KQYXSYuFFeLdCmbR++eceO62h
/0q/Prw/u3tRYhcVSk+jzb2QDMb1RyKR5PQ3GcQmq5KcX6aecC7PepMiT9avNRB5
oYu03fDqjgdgtdyGQLxIQovIta9HVGTjlEScc3bsv4Ke4yzWBBS2FFfkWfRSjDPC
NLgsCU6SQPwHz+cHk11cdR6mj6R0mOWCOSERt7TeVdt+oPLx5lELLzHHChe32uhR
h8Bdy53gnSK7wi4EhYgbu49mB8XK+WcW8NHal8lJZq5NsJxF7n46wm0r4bKpoNaH
xX8vN9PyynxOHfUSRe/Rq3W/ik8QdcVCs8MbD1P4nGsEAI+Eh2m1KnFDwHIvgFsD
/ztgwM4XEhSyoZhYP8O6KKKHQwYp4VFVlSFPIqP+yQihvviFO0lzjxF0IUP+6NMz
hGBf+a3D8L4GPxOP1VX7NdKvV9KbnUpyLiA4nJ7qjulUnTPkIgUc+t3GwcB1VHZc
qjEZAVFmxbVRfyr1xnUhHu822avhyfRkGAvY9gidPx2RDoDK+eB/UCwcDtsEw/ru
u8q3LWUrRTb4+4QRSBQRGu07oNmUDoqtC+Xf9l37LQvuyoa41Tcl4rKVL5PHmVtW
mmMrVJlQ0BFF6WkHVCIfMdb5+5S7//UOfOoFVT7HKV1IPb4QZHnLbKBOxBlaq2c2
Ae1gP0FaOG1KFGJDQKJxOhMcXphq6bC93V8BtWFJlOFvhXj7frhb0iKbWtlI2NEl
eaT2nwISxkbSGH5sHgN8KsXk31zpwIeays1LY7oXFOWCyrfw2K1jfpd3zzyw9LIZ
BCjVx4N3fsYhrdOL+VAvjn7/Pe5UhOkkPn/xcNu7vgLs7UpA7lXflwCceywBwuvx
j5o6U8KLCJbMS5aRO6Sgp6A3eqL6GqoGH1GfTVnajTqTFLxGHGehHIxMa1IDcc3d
t6I0fvoCzwvOK1esij4tseHM9zT7gdTUJAHaWnMeTTnt6LFBClTo+jbzhV+I9731
MZTqhYuKE2u2oTEeOXgr1aY09OV02n+OCQ/0iZrq3MWujE7ZDABOFgOQ7unhQGpo
/nawFq/Q3iQWbG17/KN+ZgHeHucb9um6XRbpnijNxJGqWkvz9O1BAEODd2aa9zBX
rtP4QQnaLApwI1DcrOfCnIMO6m4lejRJIy2f2tSU1T8jgjV9eut1F+9UVZJC1NlK
wWFuxPnX8PzWr7eCxJvR/WnUl5tk12uMVglLPtQcFxi8kzaZkrvoCkK9J13N80sZ
f8hAKaFPdUjTRaXyrAP1AD/UWDIQAkHXWZsKtCyu2L+M8smAquotcdNgL+WntH7G
1VDAgJljW+ZuSMMMpRa+M05PADTdWaqLiQUTZdRvaRYnLOeM00aekijywVdGRTET
59Cx1YRaSMgOluufEiwUirvuoCO7Lcmff7VWi5IimQKgpK68x2MZAZNwyeNYtQIN
wmnOp4vR8G2NeJEFw8YZQTTVasBslONkaVpj4PkZ+wQ8tPx4ZmUbvH7htuijT6OL
zuEj4qoVi5UNv5saMOL1ew1TZPd7+3tFxve92i7DhTtFr18ggPe9qdeyooAZa4Wd
7TKvlX4MwM/egYcOT1RjD6wkLDlsVca4SwDhhNib4VrQ8FGJltT4oUkHzRoNwqnH
5taSsjPchFlKoveb4XoNgefwtqlHfcffuJ2mHK/jbh91tFvSVu5pTz3XLuEpYjQ0
X8lPF3d/N9dRxl3pX/laiaGuCkVNduCkSwHACfHN5cknNlq5urc6agEIni3Rmf+K
EfJ6Pc2mIjKplFfhyXMkQJbwi1LDKJ2/40wHgqtp5uy15sbJgxSdJZ+EgfFET8ER
ADIzITgIrjgjqK02hSX7SiceALxNAVzLdgCG5V7rl40vovrfpMI6neUCGKlwIxLT
Wj64rPgZD+Vf3xkT2t5zcgTVUzb/HUe4obvhJnF20rlsKRWfMaV15xBL02cazrYH
ogzfH17QPWYsjgVbEj0QRNGnrg4i39j0xXdfhsb0SGo8x2z+HGTk2BWhTfjVnMCF
SFDgL8ZiqtpkUV2u8uwrk+tYASFxpvf5hCrpTfNJ3ZXTgjaCUftjR1sK0+oXQnT/
bEJTip/JPGVYu6aNnKTmObwY56/8BIpuNWZnVLyV8EGddU+AdK5y+lCfyks0S2D0
V+ZPd5frNJFnfojrUUZb+k8owmbMcF15WMEx5PP0W0M7vUw7GunCGZ/dCaeQjHNc
/Z9kljXSSQpR1SE5uNowzM7cikyMqbbeHHnOwcPKFh643/5n69rVG5QaiSoh/dG3
FgBEYuGp9MKz9IzVvJ2n5SwiITBYBGEK88nBG9AhqIDL9eOqjICzEBNYaDQwZZKg
AZFrrSkErJa8QHETQGXFdvVs0GBD6xaKUFDIoe2ByOh38d3eOYEYCzj1DqNFeoW2
pSvHtL5M7+GhituufNLVpPDjGgYoAj1tcchwMTskWKkiNGRnc78f0qcTN08GXPGN
XPL03NwPYozMAG0StLMMT3RVnfrkdARCkgJ9VwYYlajNCs40hb9opsCu/L08jYDQ
8wt81DYMfBM/fA9NoGp1XscDohWrQ7kjdrtnzlXmiVZATH8AiIx0DuOVLYk4sYru
lr1v7n3RVUSyZIliVlPeIWpM4yo9ATnQPU6Uq5cp6FID10kFoWkolxeaGHTdhoeo
tDqFLDaSsGmBldboxu5bEp7SNrmeKcUY6+r78OBkZ94Wnfy56weGxC+M9QvaE/0a
HDRXOC+Fad8czvLe8kYWoYhnNJUdd9sMAPgsD1/06wNDGtdaOCq1Wfpy34RozfnN
dKHQZMhzVndkF4kXFYMOBlMpI3Z/AKgsiHvihhNU9ho11PUOmTIqfCv9A+oGXCfi
belHD1jv08FnwaAM5lbg6/m7mNMKsVZvv/L+2HsvGaCh6JDR5vcGhR4KU7wsSQNu
Xt8R7Ee7MZTI3HaCg6wmz8xig7bPLqKjV0sQULlpq4R8UTPJ6fX/6+oOxmHRIeL0
XeTonwNtcMBmDIBsLyleO2QZHWc+Zrnl1Ok11HdS3y0qHmeOpOIC/rb22scAMS4h
w/eBKaH1NT5or60iVWwzTByGYU16OInPs9vVVXnb+32xZUQ5WK+BJ7BZ0VKz6V6D
Sw6FecQHACSUTRYQHx3vm6CAQmX4HhqILw3IktbI9PKIK2m1JHVX5cKaoZlCEcaB
`protect END_PROTECTED
