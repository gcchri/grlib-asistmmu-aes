`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7c+vrmDbi7ikAiaY1FPB0KdHKC4LRL32S4lx0ix4wPTu1hIe38AtMX9b1iNHZyMh
FLvxqjnyzFhvZ/becRpD7DDLC4zzkJaQg1MNHY6DvSvLbnbGaQVBaqjjrXIToo91
oIR01LK2/yQRhdEd2E9LamcwlBtjZ3kYkaiRb/WsbipDkoctsqo/s2lnsGD93uNJ
Q+NCloYQPg1m8Rm/hfjE3BMsy/0sX80ys7z6uKQNhLWevQFW4n90wZo0XcoGizJG
W79cpJA11OO20CnK65mI14ueZgEfLZwgTw/XKchPDDh89Fz6v5SRcgH3RsHWxuBL
SlgRv07zl/HZwnHHTeRbqRsDrDUe/q/c7UHMbRthBjM4ZVKTboRnPNdhlhTRM6Xq
g8wSnuHh701P+yckK0pfpp7YnASpLVs6d8R1gMrXMtl7+mGCErxNQXfN+4u2FlDd
tCLVIbHGETGzFhfc9hkWYqYFPTkrONZZhBSvZN9HwJNTenBntJlcWwloM+cKgi7+
v7kqwXZNyYnHFuVJn8OvquwrAkpVzCWxcGphugcCFx1wB1BTJqx4GdfZj0Gy1ZUH
axO1STZqJ2Jt2JudBInpDh27QvpFMtwy6IkIkSuv2dxcgPHvhzXq7QRybovNRLBC
yeIWlRe/r2zndQPUUxdExi1ohzsAWwKqjf26PAKYME3x3sEQORa2Vh2MeUicSAGA
XMjBGxKxWG0nsPgEbED3hBCtBh/1bCTomi2I2+DAG17aFZ780ZM5TQrurJ0BfUZ6
HBQRhInaHneKJTb30od54dV5+p/inGpC0vS3nG4ziJJC7bC+YIcL53vsryNFZ7Iv
c8+2h6603KHNHrH7am7eIUWM2/lOzRxacGclNOToLMaj8cjDnr90FRYO35qve02S
tLZJUBeAbvHLTQa+1jm0hkbS4p9tajVJzfxmplgtf/3hrkqNVc1duvE1FFoMh0f0
KitU8J3cbuRR34aOh0eAF6TRJpHHPFZzvh5r7zFA7STNLe4aqTUoSDSG/4bILFrw
hGUJLT3i/tS9EeBUClMiqYG2tE1wKqkOw1p5I5OQspZK1HcO6WdDDl9DFYjb4btr
eM9QM/+N3H7f4B8ar81KVdfUGufS1R5lJZAEO019WBUPnDDkCw/HzkJAjPX+Zo2h
uN1kJ4bD07pDGHSHaoDi55xD4n7YrS4w3Tr8xE3bVV8g2zWmmGsAlAyEgGmeI07E
MOf/R26+edTBmgllrJPzRpaIWK8AHtOW0FkOnHEIWZfrfyyBxG0qclgrsOnpZnw5
T6Xq797c5NRXxeP+3ZL/Ij1Tfc7rzZJIcK5XZ10F0gQhf51okf3MqE0qDJ9lASv9
amUiLC9ljQuzPSjVh4GyE3/YQk4FMfPzg0X61HSqQ4gcrgX8p0aJNKl/6ti7/pQw
3rXV1G5GfbRA9thZE650fs2WM7l5jl/nQJcda7/uDoy+ylrx9xjqgdWGXPFAt8nH
sfQNxkumZ3A0eWlMhy4q21K0fxgJrET1Uc6a0zPmOEbrNjdIDM8zkdQbtjgjc76F
f7SblQsGkudaHmPqitnoS4I6ptJPL/lma4sO/V5dxH9j3kC8Jwc+ZWX/6TWRKb4I
uYftHpt5JANlcRGJVPSAihwOlb+4px37G5ESexi48SAoyaJ38VGSvXxgpJUO1+3+
Eg25NhPxEUoEaHycjQQB8CNb2Ej6gL5Tj0MKbGMxg8PfR9bKso21yVbMwcow+Gz+
ko5G8yqdXRzml8JsR3bCXQh1n5EwKlcph9cOLdSJcaj+Xfkz1nCoDdvN+8VLBpJJ
p70HbzatQDIqn9ifGl7TDWkCTdA8GA02H5dmmnA263cH9XRtKR1LUVe6/tg1TTXL
SzHCIvLMMMOJ7X0kMDRg7xy2pskiD3LwYGPgzBCaEiiOjqj/d62JagB0jUHcikm8
WPuCPmZbTW+e9YWHFk4tqxSKbsP0ySPzTSwR+h1dTv//U0rtDg/CgQyBM4XiyLzc
8Dmulr2TgtF+xA4iLuYf7zXVkecqUD5C0w+H66DJDiRZ66IHsJBLWMaZiXn2x6W4
rLd9n8Ws/YhTDzP1Oqic3sWxZCqC+JHKntEMmXcz2rU648SAGf7VOtF+3xCuPJ9G
UJJDQeropCl7J+Xs0FIhxzC7Z/KEOqHf1eSejWOSy+QhY+N+DsC1DAsIKciTQs6E
MGxNnj3uQNjV8gktYrMrj7zAoBOpRQDRIuI1Vb28VBG2hmisciHKQN+O25oSBTaA
O65q1rezkOH0psQkfULUfJdlsXlWalOhbAn5pBtq0EVIeqY8k+ZNL9RXXztxiz0s
ENbf7TnxXwYkfIgBGDKQdfA3hJiOP4EBOFJiiBQb7QhZp/m5egOJmtM6MG7uG6j/
VUZCeICsNTpwbVk+ag5Xk+ldnd96lwyWN073UYhE3YWc/gLKTOPQJd/F3XdLQ18x
kQcmWNH9J8Pryt93e7lZnH4TY0rsJvMmggFGoCRoIN/NJFvwR2DCN3+qtV9bujap
4Evow1sp92qi41eiyBtj3hk1Tz53XMbroWrcvRqb4K3YMSwcKiJlbXd8xMYqpcxk
GTQyIIBCQqNKDjELUDBvN6bkW1bRLVckiERzpCoiV5fumpmyO6yDsG9bIFbhArpW
WaXBK9MLytSlKxlgLDN/mGitj+j1+X1CHrUTZVuDTEFTGfYjQL1/8JIwCSdNlbRc
jK+sMoDMs9WNuCCgCyerJqYQ5B0xknFRfEfrsL/LaWV3zNwjbfnwdw9Rf0iS6bxg
9ZHX8iZcugbpnybmezWy75DSD71dPFD99Adphypa0+0E0f8I/q3j8McUWYDofNf7
5ArgYonAkGVrGOo5BsOCFgPoUmYWqFUpz091BIiUvTnR2wOixM0Zwu0fO0QluFK0
kqbxM97JqZHyPg4xXy5mKzmmdmKtbr8dMjTGKu4fWkGhc91xVkBxzCWr6vHcoqag
xuloSxdqkMPoCyM2KLgMuA4rZoHVGVo86sHXgzrlxdQt1axOU2nQR/WbSuNhhQ2f
8ZORsbdaqdD9XvAzX4ZUnscRlnmztZvAxNWUaM3SIeeR0CQeZ0UsZHcIPJX0pr8o
P3rhmZpCiTD2Wt3IHnk+cKI3RMHFr2mcbu0BPzjRo/FOXSTO5w/nL8CqLXZdBXoK
Jx0QWXmMrX7q+AP3mivOprsW+J9lhkuLHDuTqnNkNh/DKnDX69efxAMm+/DRTQeu
avxTlIVjgSDji+/IEqBhmcoX7EyywAD+qzq1Qf0xXeQj/M7uKKw5w99O+/Sm23QE
P//VS2oJFBFUS029pl3LBYAFc6S4lYGs+Yjd18MYftoxPB9/ACl/7hYlqXTQX9H9
82g+wU2NhWJFBNIpbHSG/KDbx5n99OMb5cebwUvR9mvSVJ/EiXpxkgOjzBp+d0/S
pWY+CrQCSwqLjbTyLdpJ8gwfiFaLm0wSQWMKbrFKYz8th6afFE92hQoKjHxRA1wU
ROZy1+aK8RO7OOuholr8R654EZQfAY4da3GpePygHvLmf1MPTXqYNp1m/Qw34nIa
FMKm5sNi6UliLENkUxVQ1UrfEBELYmzfladA6JpfKtJ5/pZ16YWNGsqVlnb6pbjv
wqc8DD5CfLdZGW7Lu6Wbl/JZwv2knH37b/G7/J5D62bjors7TS1tgqss2EaAaquV
nXWcSHfrq51VXx+F9O/XGrDwWeZn96WnbocboZ9fDS6vpzIpNzoF2gR77lZe+ZgG
DchxSHRKQsb5TItRh1lQZoHWtTgHQQjSUC8KmbSLwy4+LoptbXcvIvEo5Xm7Q+lw
jvMsxnJ/lYw8wvFpTbnpCb82K21eOWjYNS6OHWzghvFFNFGZeMBHPKYHUcghU9+e
FHkLvG7JWv2/9Bi0IxdeVRegChvcRsP5wCVCzL7Al+gDxiKF5rKouVkzr1WpDEs/
mX9KfVsNRJgFGbrLkC9A4bqXXqmzwfmm5Odgje2qQywtnphmjqt1mDsvGgf5yMiB
xeRDFZk+A/9g3exXC/CBIthwKDePEBHuOqNC2mIoCjfWock6ORYk9DxZICMNGHl+
RA7q5bR0Xv99PYo545F1NxlH7JJ/FLgV8ruUuBJahR3Y4sFgweLiNG14ng1IQAyp
F2fxCal1rXrXfGNDdLc76OhezrerGb3MVt+1n1iFlZf4CXtoRthYiqlWYSMHvEGw
rOxNb//OEx9u6is8fC8PhGsDlbBh+lZ6mKQ5UJBXiauAC+fw7SCogbeZsK+dq2r+
+Ze9fbA7UD4beov/WB4cLtwQvb9LVNL8WPw0mpBrEUL1MI9Scpb21IONBzxNWL70
FvgE6BbR2IQ3T+nfe0uwB6ZBIaBweHwZJROHTAfwrlhJyuYLikyBQ1JO7TZ7DyNY
2bO1jqtKekn4LicESlNiU3cOI0d0ngHlIG9OP/qR2ZqMHL6AC4NUPlfo6MVuvFlr
BuVOuWMJubd4fdVjh5keeTQQO39/nr1ZlGVhysbfniAm9Z6Tx+8K4SVJmY5QAgmw
W17Q3i2/oUy+WGGR46r/ynSbVnx0FvmRAb5AB7KCtx06plplfgf5Ww9DJyMosm8j
hc0gicyoOE8Ldu1mMbfhjYn2eh1PHQQD4ryu/JnOKoAmTDlXF6XdqXCB+atR889y
4HIVhMfu4H1ufy49ayiPlwNnDICE9GyFP4PtqBZGmXCDgTZzdX2+/WpR9CUJIq9S
TzErJZ97NjAwYoEDo3K5Dpmnme1+lWYL3ejdVjIjvhzkbE/IzQcJdjWOV3blUWbo
527QECWXx4t9MOziOPJ1NErtwm2HCXdsGBcQrFlYOrZJ3sHkcMEaZI6L1F31Nt+/
clhsCzpsGDSSnNxJhxVxmxF3IRCU91ROUcT3nAm8tZiQhf6vqwzLjF1AhCgi7ZMv
6aMU1836sk92nrICARkf8koCeaG5tsNoYhTeMmape+kQ41BGPfGdnpZmXn7yEd/q
1JPpd5f/nEPoWjcQf1blZ43Qila6qM+Ajlk/fWfq9uzgey9h3QjJ7+ysA9Z5RTyh
GAcIssjzPsDCbofbDhDPw9uM+xQfOxEDxJxf+2q5GIkCXSSpgmAeMiJlcxDNLBH3
S8WzfbYtM+cLNzW7sC0qvmm4C2tjOrkeSLazaob4V/C3YWxOUkgO7ClCeLBCKetS
Zfk9AJhjhgaokqju94OedymWsoSq3+uEv49jmkb9TmuxsGOq8/ucq7OWv4hoGerv
LJprkd5HSwQ9m88XDSsA5sAZjzIYDsjKWjOXsw6sg8HrGmVkTqQEd72P7y+dH8uP
rzx5XgkbW4KoawgFNbuHlAysXUxVxh0ow4Mo29+jThmtCcWibF5N+rXib1WLOrNV
u/WChSDrhFO3qIH2Sktr/bdKSaLJqapt0jAQuQjZRdjqjd2/3tkXKeaJYkRQRPSG
S8ocYM6VB7LCY89MgcpiiP9Q0fqk3lSOBo/ILeQ0061JG9Mn8DQL7tUCTgyuiltw
enFhYvCs1O7g2cHKMmMF1R+1zEekvB3x7CVuNVqoJ7AvBItp4j97TZmvSKofpP9O
nz2TAkE50eeNENgLZAR3KkvjzGBt4CowSfddIl5JOficWsdycRuJgYD/N8XNkdEL
IVuxkExmsj+sn/h56feYyh5s3u4+iEd5u3PKbM3zNAZCxoWEZwNFTDHlhA3Qy1L6
rJ6j0gPS8gRNvJXylCwazO04/HfVVdd65F9zE1CmKepi+fmJYeLVBK3E1u0S+Jgc
Ifp6bcg5u3PvbIVfE7AC/raz6/GuRFYRtxZVMNmGIew9m3Q7xn2uIj9L5cpRe1Y1
ais8D6ZKWg9GOftBtdxcA+JvTwtBH7FZdiJetSzK7sGoFWfXjgITcD1xcNafg6Rk
ZOOre4dKSS14mDvD1Mso2VNJAQ0sp26jUPSuHwCngqhnrFBxSvDHJKDVvhbiis+d
0h0DLeyrV8nRAV4xf/b6ow7ghqdq0VB9HIh7OJq2qPd6EaHTmoI3u8Nj/JCAahDj
kJV2SUShx3NJbJnw74wB7jcMpVeUvoo+6ho4Rh450XuZL2QTfNSvcOtfqy2dMGuH
hCExluCQzvWkkLtC09QT2DVjUbTjPQNPXnt3JxfjNiFHa7qZTUnNL0JRv04P/n/3
UN29+kvUYpndg6Vf8mc7sOFfD4FngPXyIrpDafuV3lDPWm2cEdc4EfYkF2wD2YI/
qYsQg3Ag6H3HWietZT5bS9dQI8uDVW22PvXX2opQMpF15VgLAQUGaJBe7ku7ATUW
ahOyxlqc2PUtifSjt7Iagpkk3R9slNC5iJuJVDnCCce2DcI+bjmQtxPEcRAdf587
xkWTt0Jkjqu+Ny7qsceuCCHZgMmgOsRpiaMHP454a8QsbHeWnWggE4oI95Y87M1D
tjpl9ewf9DNJnIj3RehAlnPR9ttIYML63N+R8+HvLmHMo3J5+sKeVhHRVrVsGAW7
dtbuanEtgHXnFfVcBvlfwtrIhRovFtqtzkwNwbnT/4DmA9rG4rgUFeypsUzes/JR
gWJFvc2gwqK8x4IHsiwUbvAAMVpALRSsXDr9EebKxclipnJ68zH00LuFw4iB3lxe
1helNA9gr9mRQDFxuU/ber2+yAO9JTUDBBuF0lAp+zPdnHmRxJrSh9EWiLL10iHZ
g/Qh78wedXT/Js0pBxj/AHmNLQ/yXBFq/b54AxFQRptsWlwcqyusCMxnjxz1nzRo
bq2URGfjpmeuZ3gGNs7aHcaSTsh1lGu8VZ8A1cfTGkaCWoHSjx5T/v5gg3iF9lhl
7cdFFCdpfCMjy/VHidmqBMjkxVowabMLynHx80bIutHfD6VcIHOZPr9Ni/hYcAy6
DHZ4s9IaDSjIRMTfduWJqLzicAOJDeR4RYiY6q9GEyUBd47yGg/cAS22znqUsmbR
Q7ATZZiWP2jF9bH3LCCAZUQ81NjZfjLpj0jaUPm8KBJQF2nwuB/UAPHtR3by7ltP
ircbhTrMoZG/jV+f+loABTaZgoDx6SqfYgAc3c83wVvHo+2N4nB+FBd9IwyCeMG7
VnLBdhTZyHtqFYRyUWWA4ahi2FC/PxR3EHxqceuJdsexTgEMhocQjxGdGXj0eogD
YVhxw7FeEv1zU1CKp0FsLJVAl2CatvndE3sB5vLavB6ZS4Enmulekf8lfIqSNYtx
UOV4QUrWqyAVqkMUHRNEjh9fybLHe4YW0a9ELJ0mQTtBxcFyBMUwq2GzbWPphngU
A+1asxMBXdq2b7lHRnns8vTA3o++NBTUaiWlWHsD4SowsYS8pbzwgzPqFNk42Cfg
K9H+ebCKwy+cAA5lR+Ya83r0QDudyFq665lgfUt7hOES+Nrzv1H4tAcqRGT9ENaf
McBYK4y7VgiLdh2cjMnsYsg+JxJ0VF88gvuqm2cJZy9TkaeXNuVTj8xBfLrcObw3
D2b0QltLXV0n3JHIXyXIY+68v3fQj1//J57p7TtLSJ9bDgoce5/N4CPC+SWMvg07
76/1V3FOgbgEjaYGwFfhaohI4kfC/mhytf8h+Z7whPfljX7kE7NMs0f/B3zX2ccM
RbG/srk7ahsm0R4NazVroe18Kq5e+PvfJxY72bBXB2P8qWvR5dJcIo8AukdcWGIy
DJSeeeRu0T7Ku5KUMbPnZAlDNpoP95CS+7AgPvKVKEMohJtvM79GCCN/HqLX+//O
2NCii9pjOqSBx+shrlBfA1r4i4UqxUV8UROz6vTLum4wmjNEi+Zo7jpJDzXFZhqb
AVasd0Rfug4biNemYBD7B0ONSTW3GMRp9+/zAYzETmzNPByk7rmTxgQIGnvUtMa3
R4zufn4bqTtT9dIVs9jTZ7ssU26VMYHSCGZE6ESN4PVfb4bqSNS5tuPMZqOFtx0R
uBtRYDnaSbGa5ASwLAQWZYSgKTgJwTUv2rdBTe3YiMmOfwzxfwwu313pkPYdMOSi
NABFd0rmKhm1wnjI0U4v7251HraZL3/8VhKWeBDtl51Fb390DGGNxNaMTZRsoxAt
xkmk1CNdw6rRfN6GML2KueJQ+2V8+pSetuhFDmohSFT5Q+UIqTBXh0HBS14Yvn5x
2KndVKHYI64KUZbapAOK3WBya3qJ9WauaCveIIxf8/+PFn2jtT2Pxx1l1dupYYvI
Q3qwm87vDzCqG/x2LgmNjym0lJsS3vhzXX3xJiP+0cgDI5VgWVypE1C5byIFAgh+
/ez6Wg++NE4N+xrq0A9K3M0uFsChTm+z6cnSjb3gZ6eUogkjzB7yqUI25jGvjkBr
BcWhhkCxZlyM2I+3Zy+mSTGqJoU6L108Px/dJBegOReesAYDYQwHbCAjLLG3P0M3
aQq3skDQeXfjgIdjVKhefyjdAutaFkSB4QWqcgZVj0nOespxg2tVMa/+Jym7g7ot
QA7+b7pIQixP/sMf6UsSQIuy3+Gv9kCgXQQiOS9ufU5NNam65I65Fmeonq28KlN2
4yWDDMIL1FESBeUkJRTeWo6JAF5hC7ARyxoequLNmviKkbiPQhhxNF46ZeVr8Xtl
P0KKjH/jbgiMC4YUfTseyCOac0a1gqWDrBoRt0vfsOVxc9uOPUFg1tXjNHhCbCxj
nWNy1RFPrS6fuhBIGcxch5rc90m/r8ANN+8RTdLAQFSYovBkYsT5jwRqyBbSxEW8
J/ZSipteu8gQ7xB+TZIk8XNSXkntTw3bTFoqGYcA1pAa42c/+CC/+AqDjY/6dUfH
uCOWA3cBo4SI67Pn8HZjsvFBsdhZXHDLOrMAhpGIjbUSgc+Oszr86t5KRQjZvRSS
ryWbHfREh+AuHai4UP+/Hvsqm46tMOoBpoLT04OC69bSGp96dEBfkY8E7oppbjEi
t/7MWD5mQutYnVUEMBQLMOCWgyZ3nwHCkp3utWAbtXOUp3Wx5oizGwAU5PSfvZ/e
CrK/iKbS1Y/flFNew8/P7sY4leItypj94FAYBfPsA1jCpqRL6ghgWshtf9HQ75m1
JH/9k+f10i8HT+CFfwJkRwFgGu0PaF/c7y8HT8EuBVBZisOXGvhJyKrdyAeKpwxl
eR1XGtPExInL1Psq83H3T4dc7WGFKiIS/mdPVz8FxCe08bEpYdTl6k0TC+m3z5nZ
iysOcB60eMRAHx/DWH10H57ukb3/nYWWyCAtidmZBzcqDyBU8Fy0TJte6fjZa5lt
zNePr+tddCvXQd99C0VOWSHQHfzfyW+PUH5AGz+X+pRVi4owN88+ceHd/MDzrJOL
VlOuuWD43XmfgMX/NuLNcWabi2o8egQxJ317/nhiPt7EVvjjACiFRcbWlgNnczEn
BUe/KyPO6HkqxZDbv10Bdq5JM1qjNlo2iIZt78qGv8fUh2h2NQUuScnwhx4D4p2O
ohNqoE2OaioaLEfSzALKwv6YaKKdg4kmclvomtXDtSA3urAbtRHjmA5LFMtKE4oY
3HxmP4Crp20AmtbmsmxpYs6M2anWDbnUHKHoWuzAoRNr2JLyoD86liubIzJ7G37X
V/K2uk4FDdPCZcjiLJ2/qJ8g1hrTe+Kbh365MuA8Rc4hlSRMUwgHZ2qku4yLcXD6
xtfVa8ZR5eavB5Pb3jN9vfllmL1eWTZUJiQCAWs9Lm0hgEiu7JYIa7vfKQpfQWnO
Qn8HQ0p51NFk5hnhrsAj+JJG/vtUQyhp/cw9b9Mp2lFrKAt1yJIg3ve0OnHofCta
lDSgYwNiyh1Eo+YczjIPUTp8SrfmD7CIKpKduN9KRrzGa0jasNVYHxxr0uzbPMbW
uWAsi3MGEgSVP0JWVGThCUOIjFFLKSOFJhgXFape81oR6mfCE2u1bbY4whK++04d
j1SZMOyb7HXvfL+jKIc49xC6iMbrWWdDLkaxmHcCftDeY/fxsMR+ftnjywN/70Js
B3noh8KajK7ymvRPd9I17Up8GuDkAqII1PSn5AKjMZO0+8iW/1kQFZxtFZyfn3i2
p0mowX0QWN0FOGdwFLEVRJBTU7JYqAo4EbOmw1QM+q0UUZAWhW+qpX0ThNXOBQmx
RiXIR4RtV+Lx8XU3T0qnK/lq/Z82XiWUS7g9lY0DxOJel0pYmFZUhynZQL2qkQzl
nGh7f5YphftB7H1RYu9Rc+/oOh95toP+XGacKXGUyPsKRlcHxyCBagx92tkfHVtr
wM5dOMPc3Iw+OCispd83T5poL7GOQ6HPk2sZSTxnBjRfueamyuoQ4gIS3nyHBm4E
rsg5+BFVlUYHJT2al4smE7Wu8z+6IXS0VV2zUgz/ArOTCk4HAegGDsiSLuXwSXio
CbxcJmDlbXU9HJEAxcBtbEDio0BWdUY4qpkg84yID44xdDUZJajreekZsmEM55kF
0HO7Hqoi7QV/p2E0ggH500XBPv3MGI2pq9e+mV+m3gLVO9nqZpzj4UZQOWgnUyLC
rgAV3SnVYRaDemZBB4a6ht3iuv7xaN9Yq8/KI+o+8MA7V06s8bsD7yLt7DqfLqm0
N6GgwklrWuJlfhWCOj0v8HBylhp1h4GJgQ5vc1frkW9JvgxcGsDE9XWYyHL2/KMa
vP78ByRVJn6aEiQn+lRYKbRVXVAUuBw0Qg+obaxWo246QiOFv8I1ARLczbf2O891
B+Kkwk4f+KmqwsbHTOR15hhpbZ7YT8/vtJz8HxkRyx5LjjdtZyn4InmVljzlr5Xn
Qq7xJZ1vh67SUzJtEYZWzwHuqs2IAsZwvAZM0G7K+LXteyB47BaC2AikQQlkU2cu
geiosIY2kykkJN3YtWzasWXaoAistcLQUBAlhFrnojXi10pYoGousM6RjnGLhNLP
NhDFE13wlSC+0R3/YzSxtWfbL7IRAteO2YdPrmaevTWGiHdvZBTfXzfyTPmOjxLy
9Fx6xZviIOx5f0kLzu4gdsaKeJfdGmYFgopI1NhhFA1OhgNHnjuSmbd9T+v4rOpP
BPiAJaIL3s5ESmspFUaJhUNu2hutbSQYzB7EfZ2EXPPPaP2dLojEr7/R0kqnQXsJ
B0o8CbUWILX8sAGk21+L2ue5ylpz3WvG4GftdWrWh/Tk9hoD+ifP61RyvHWOZnJa
VTLwVjF2ijC+16qMDb45k+l07+KfHHpMfejiiXCjTTOFiKqwKBXC+xGHhEvHrUDV
mLkc6aLsGeqMhYHcMqBRSqpgW2x+hYjnJZSlaw7yoQQ5TnZJQeQXsixBgyEILCap
mp+G/lEjqii5oTt3SA1cnHgWua/yyiTN/BP1Z4vqgOmbn6xH/c28FqvqhhF80g+2
i2oogLg/NtyDOpM0l8BAOmsUbTZiEpBZuIEuyziNEz78O3vIHRNCF+Yod+H0hfp4
ITEa55li7PZcmUSGRD2lfSQ2/w3dDTFSYkdInW9sT/XeSmnxXYZMtalnNtZDV1O5
oCNE4Iw9qh+r3dNl3jTur0TkgcexYn+FbyFHQdSc/a3DTnOZ0nPp2avmd36kjRVr
WyfNgMS92ivdcwritk98YR0mgp05cUXp2SSJcxaTcUa4YiWaXfyrG23V8G2jUWgz
MhtQbBb5FNwvvWHq1phP5g1H7b97dPizJhko2c7HXYxud4yrSAQLt/UU1//11WOe
1w+YZUC4qG02aE/CDwiEpkGJzvLnR5gu43O2tzOEUfdFUZXfSe/WpGcBtj/F95T3
cnn9HtMc+CheR4ZSAVQFIAs6Dt5vjmYjY8485GpRcrLC0tEo6hFsur2fMBC/gzH3
d40kHs7d29oO2uy6rzR9hCkhgtDORX+kQtjtwliljJ4J5F3sIYjhuMPtJnuq7kgY
7jUHgqkeG0DSJGQVlV+4TNZLMcJ3Thyin9BtvMjhBoBjhq/4iWQ4wo8drTf2fjDR
MC16VPWE2p8OvgTWm+AwV0CNjOoLUphNdFZ034CuI6BzcXv0JH4pVUGjrgPmS+SE
pO/jnw+s2dnzs192z9yatWrXUox4gBd5huZitSnl/ewt55rM6+/Lt2vGSF4O1Qn5
GI85yUDyyBnCU6dtzL3bDX9tKEaedvzDeAMY+t/tPpTrofMw4fF9d+XG7O2NLUcJ
11f6p4siXf9PvsKFA7qQz21wol3SljLkjjwlbm7wA2OFTXjZ+btp0ZNpAXzJFCTN
/SxHeXyN0EwJeJaFB8RYIto84QP2GXW5GinW+vpmIrdIlRSQ5UVUJFjIdznobu7o
u5GoD88r4QyURZFh6DsWWewRkjXs9JZxu8AhDak8LLtBNVtW/5bpK9j8F2/WZYCO
Sin+44LmpO1SjFelS/mRf+gKdHnqsxhzv1muqoTyqxeZkl6gyg14vQox6TaF8v4c
npZE9qoBxrfM0ZRX2JaS3zfkn/s1GZee2vIJ+cTA57fFAx8fOT9OqVj1NH+KCl+h
uvw0VtDwOIc3CUT436jSNTXBx+6zwgyT9S3G79k5WZe4KutE8cJEGU6fyUCScHjL
Ku02pIDP5Wz07NGzVbLFDbujgCbNigrcPjU5bml25/Hdrz3GuGT0WanubiX7L3CL
fnCVqTuGxOsdtoGeVvr3wpBroxC3eJHQpO59LbvfKHadCW9iDiiv7zPgYsRAF0o/
Nh3TL2r/JTg1c9zlCuClPUVBsDUdPZyYxbHW7PdvCvvIz500jRhHRaaWh+16AVDY
ekNASHJOAf9C8SXPJqyCuRmr4Bh5oDsBe1vyZM09OOeAb8g0v3wu6HeBef+/T97M
DFpDVHaI7O2IuwHAI1qP9g/uQ08z8UQrDTGfcO+62s+UzeIMDldcuhD6QCPJq4+K
VV9tttmlwLYbv+sAk5jyKCVDqolJd+FNyCcMQiMfLGQXpIB0W5X2NsQml++CBpPS
hRC+hmzDbJtuFKv+QklKrkQZ3Og7q5ZjIASauumVqjRk2X85LOlGD8HK14csC2bG
UM7+WBGxXVOI8Hc+FOkI44wOTLHB1jin1MpEffzjB1tySDkp5V2zRAcwoK2T1kSa
sXN9dRH74oPLAm0jdwCfol1ztu0t6/bfo46DTJ9sz1J5sTxpy6HB/K7cBFfXfVR0
ofN47TUvHriFQ4wENnkk4ygMbsJMHIdYsFB5f3Bl45h9ofW6rpYtKAMfR37Zw/Qz
Np4t3lhjAsTDdMqxjLCVdJVJJiDICx8Gkt0Adq6wrBB1A4rEpjknnQVPwAQ5PO0Y
iD8vzVnIFdVvNVHmPOnsNq79t7yrCUIU5/JPGLTqlx3X3Gf3I0QMdI7lmJpGifCC
ku/obTFTGTQEKCr8+vHuInK1KqjOKVyF8wZtxv/DPPdgnWbFGQ9FjxEBe/q5NCXZ
QGC/tOuMRrUFZ8Mb/gIw7w70F6ZjcMmTyWu4PU0EukWcuBmPEk7OR18QqMAa//kV
o1VJBDuXxo064rHvG1Kt15XOSVu6KZLdSM6VvvB3upF/vaPAy1UqR/vxeAOM6wj0
MSmww6hJM6pwob1Gmq6ndIa0G6Ewrtc2BIMsxxeyffJvAamRWUpPHeoTTP5kvi7C
tdGEhHuSAuZRJCSU+WdiyjuI3rDgics1mt1Xx73rbF+i2LF5/fnlqMrRZeG8zJN2
lqqzcokEeYEXq1DGPmGliOIVrNyWBQd/eQUltFlXy51/jEdhVqhKQJs2GSO+Opab
gaMmX2GTID2WdaaeKyMsdSBJdUBf10e0C4zxePUdzBRaIlIWx3vo9tM2jiI6ckh+
Kd6Ol3rQK3VXctLp2eA0JJzxAb6fCUasOpPKLhtT8YB37NllGrJCwQ2mv8IxKFeO
vwN5HlqDXGkmgRZaLCg7KJfFEW+PARNHl9wfjzfyH2bVyMzKlvQR3AEGl6Cs4nRC
F58DXcFY8zopDfznYaC6MlqTL5b+YHd5Ktd8RBLOUzDdSUaJbCk7V84XF+jVgJhM
+KERsTZE1WMme5W4ckgsFvmZ7uQq/ZIz1O2QDSzY9WtadLURnrGe0aHTms5PO4/T
fbMkgEDhTubvQxhFAzMloQ2ap5KCYt8Gh147yHfKvvP5E+aMbYiQnnQXobCj1XiJ
6utmwjsAkSdJ0Vika0N7Pj3TdheL3YgupsbSOgJb0lBryw9hesTjoYdur21hv4OT
UGPgzO3tlZsVS+cXa+QWBbctY9cchcKlorAf3TmPDH8X8N93fOf3XO2NdAwnUt6I
14G9VRN9CyzuM3WiMN0buVNu+jKPlbxvf525Puj40mJlHFcAFfxa5jyUtkWtSErH
URTSFD0dIP5EWRp74hVKr4I5bbrzohA1IiqDQBUONLqHcXqixmR6vTqxGHbrdWrX
ZAG5Q9TNmWuKvtL32fL0Y+Q6Dl5hXUNFcIS6AXfh5ACTZ/WJliBHOSCf94C7Wh3Q
PowaAXAboLpS8Dk5vslrqb3/Y4cdmEyR8itN0rZFO/CYqHycgvW4JnUlSqLeLudN
Utr9FxWZDXXFYRHUoT1f3lppw50cpX1/OG48LIfVgnAuaO5zjyv0+17waaNhti9X
8Cie3zuKhfbSVGs/LZKCCjbcJeLoM2J9yUc+2Oe8g3O6sZza1XhDc6ZYSUog+YId
nUNgE08M/1Bwux8kZ2ZIryySwVhchHXgfJEvo66X5YEtPRcGsNfura8E1sjQQwIz
fCalZBibMNCdGrSZxNYE+rFvpPDqkJas2RqJx6XS0HM9q7tpdrQEOyOoFGlCUOvq
ecBQ97NfEarwVlyyCCDmSVv6lXbM4mllZkDYIBxRgDBex3H4TwX7EwEDjwg+7ZyV
USUZJpJzcjA/9+d5AvnWkA53M0kqZHeBcNvwanSvMuaQR8k+YGo/YwQ45Gx4oti9
w+gGh7BoQw/OaiXiPFdMcwBTIVXahgAXYql5xx2inBDkq8V75L+oVmnYv1g/YRVG
o7eQew2ASonF4rGPVK9iyye0cEuxqMGvs22kznYFw3o9/Bt208LiDn2YvdZj5lrs
XPhliTMPDx8CdHShTVcMlIMlG8GDu2FX2db/7loptE6D2lZ5r8WJHvJFG8jbZVia
5z0vMxkJIq3yo5Slka082Osu/rLsmqh/2rsk9FqS3GVKTzv4lygTJWRXKp1goM3l
62Kcj7P85kMFX9iSMiivirv8qr0rC+eO24QuJrvdf5/Sm1byKF79BTpdeKjB2r8Y
TRH+A8lnabrFyV/v6DKtHet6Ctk18zLcq56Vm9vShi4ZPv1GHHJcr8Bart47jLzG
60iXXoFwUY2KemCSFEDJVdizVaK/Xv5RdIGL5D2cDWnvqrr134VQIGz1iyVCdncP
Sd6fTi2zDYm+hWO9FJwsVouA+AA2KYA0uIMHMK0441qWQXLZV25zLDKk2dN0nArv
CilWYfXhkLq15R8qS6CJcb51aEb3D6tHsuJ18GxlkhNwiphYGZqix8ZGIPUxClgZ
tOU/rs/+f6RFkU8T6QzKGe10C5bTdeJV9/0ZSokbc7hrFyJAhCwDRQh+TDwh9n77
+e0854J0q1rit1HawZUOcwac4nJzTkrag7Ku+4q2tAr4z2i14uAeJ23WcCMAjPwd
jECrGVM7MriuKj3As/qhOvQH/FE2OBFth2pJ9tD8Hbqx8d1VOxNJNRQuUdeISB96
rp3GfVmk/QomeIdr/fH+A5wWp2FeZfaJp2qXqio36B9o9EGmaGN2A9DUvs49AjrK
dvTwUNd56aBn36QR4XWOXF4gaBMC/4+71Ute1kAlHlFHJRAq0uwybMzpd9Z8BGOc
lIHwYFY+60uAAe7YSeKQ4p694ktRaOBO1BC/YPYML8SHqyFlc002OJ2/0LWIVTnj
XZxo6y7JOk0UmkAuP8lphza2vmEkG7/rnDInmD/GICaDvHsWHQ9irhH4wpPkKE4P
9WcZz0UaCocZ1KzE+VrVL1cICulXCBQjLZz78vDCYslFIsPr+mOrKjgE18q4yYDO
96THgkKsgMAygTfXpRvzM0fOxcn0MsSI3cDb4SedZiMQEFEHsImFx/SdNEM/162V
2kwMowrK7a2GTnbxih/ayTj6eqgHvwvf0bxL8jxL1OFjz99VEe1AWUH4PLMlXVg7
X5X/dwDC8kGX8cTfEl4oPypZrFeUcqxjymES13Bg5Ia1KyloKWrq3Lkb5lojQYZo
0IBBGVQsBS2XgzYXYYPyxiNkK0mt6531itYtHiTbYK4SDHVBza09JLNPQyhySYJJ
UbYvbcDaXVGr2MwXmO6kjiRM8BwrikPWO2K3nVAXrnK86Z2LyCOTgnZFfSj1Nf31
yG802wXyNwFvKoJPXlIXfRsB1siaYHWWBdIIIiNhbb89EeYADWyDTvz6w+DPo/ow
qaXadobyd+QEuPg3QELLcuu3XOqkAzvwnpbuBAIC4civa8Q0GcMSirhG/59+Ew9J
LkIAEEh3ruzod8VZpWU5y4z3tLDpKH4iWMXAdE5C1FCqTXZsuaN5CNy8KDNkY0GX
EpIDivawk9u2RMrD3Ihpiv7vJAaP5e1akY1Dcw7ixLUZT9B7J3qCE7md7z6Q4Mfu
28NC4J3nQPnEYwoGEkdT5TOGhz0EgawH3t7FXVUpzVtozyTLKQJKnAsZfhRYruz/
u5lZ8tIiJRYIDspdE46uS26ipmPw9DgZ49NZAeUS3NaPK1RnoXSGbm88edzU7pdU
IyGYxSLjtH/eDXrNeD7cRJIFihzrvuWjat6j/EPGwOO8YDhoYiOOF7CH9EJNSaQr
TAbhog7+dNOAxXoY1YM7lJAX+bBoMhUeTrdEOIaWSWkvzwFFobYhLBYwVg4LYh93
KK5zLd8OXLj2zTHz84AB+I5EoqJk2uu2XWAN3kTGlxP431AmRrKJwBMvIy+Sv/T2
C7PYaws3q3slJ9zUxUv3G3tNAZOk7tKPtKY2T/XPdi+I6i5zFJ8pObjHbHkouCjG
OTMPEZa0A4sfPlJ+0HL87NTWoXG236cM2HmKPbHM6BfrS6l69rh4lT1rZq8Xz4M0
MCxMx7vIXmbge/mGSF34KC17s/LWw4ZswQaZWOZHWhWR1d1WGJJcS6OkD79TvL7j
YwGsrxvUOQni7IDsCyKyVerX9Q/RuJf6N10RoUoGmfgNRNOUQDkJ3BF2wlaXFE2q
cpco+u/n+pgjOqws2s8XNN8BLy3Tx06U3uXJxK5wneGPBHnIAeUDlGlP3qXAAOfK
kgNY9pJKbkDIXB4bKYB0QlEHIrKC+6Wwcl6L3VUsH1YjqWgUZr/45OtabzqfPVG0
pIZNllIwKZBE4tm4NJooAXlQOT5f7Y3cc5mfZsPAI/1TBPqduba+YSpGXef64woz
zYEyaDBcnFF81UEZpzXQesgFe1WlNrsSLbqQoPbWo4Erk48FpS8ElPovVWAwze8K
W/MP9i8sGbDPZgnrUGm+0slX0v212FVFXT4N+JGWXroHmaz0aojxTeDFpC/nYodC
Fz+hHu6uoo+/+wzRzUCE+E0Crwz36i6fbZYe5rhY/YP0WUaso1L8G40QAPsphh+H
aIZKO44uDNPsDDIce7u+6ZxF68j3nDrsP/6ZUCWLFICTjvd1/Yzont9aDhQMjV5h
T3tSNfMwK0AlD/yAQKXzaQ4zVFwdd4JWuPRIyWyqh0Pz8Iu4+COB+FDO8LjLrtLf
o7g8+DBSZx2mABB/1Pg/MVT+zWATLXMRF3/QjCCb4n79FZHSYvlVMFisi08dkpjA
6MBOTlJ0GsJqOwFC0I++jnTIKHvuSvb82FOpUtBgTCbqhI5J8+szJPF7y/2LBILk
UHr7lXISXIDycBctX3Wnf43raxUvRAnoEUiMLo46IAvCGvgwFVSy/NhCmyfuvOha
va5/BTlQuS0q95WyVPxM2ytAwj2HrVTn1Yh3t09xQgPZhPDab8W5Ln6x2QZKchm8
cLTTaivMnqdtLyQvDVWqQNnYMKOFL8T2gKyLKAhgYeBVpMI/I8EJfIGZLdQp22mb
R7QHBs48nSjGOXl+JnYpNUZcFlV4Z/6wq5K6ya/YjfNoDMwdoTRtsCBoS9hCqYPt
/0yQuS0x01hmkgtLxOTQFsvSuP/Ai5yStP5p4aDhyzB7dIyJGwQJx+xI94lxLXj2
2zCM1teNldmcDVNcEWy0bIwb89okcb144WaZNdF/3MLeV9B0MhNTJQLCiVtxgf1Z
8xsN2h4Jy2A/nbjlVTtY9D4wNdehZvzJyLzJZNfs7h/JM4rHIK01FG+R2Rx3xXiu
xevDKfIA26LLCkBqFf1tuxmUzLzsLIvFtBtauXSQ1gpf/1RlsPiAVfu8AwVNel3F
SCAOfI4qiITQcIC7afL0r3+13O9zQIBwk4RL2VReLE/RItK+nxbzdmEG9NYJLfIv
hkwXyYo6RkUJz291qQiPIHCLqt02GTL30wgKlwjWxXsQ3fUXNgW3phVa3FZ1eSZL
cxEuDQyCmHDWxFlFPgUV7KXgH6UmO8YKN32ipgxzk99BeahSMOo2sfxvYpVWQnLr
J6fO2GrEs8bjP3bV70VNj4risevJbNQAkqDIf6UqGo9LTd8Hx8knS6DpV+FbtXf5
VrFW3XF6uinT/EyJ6PExI/PmCOB2RQRhQLekjUZJfIcTRD3FQ8k5cN98zgARVHC3
33Mej6KMP9K6/imLLf8Ba0vpIvK4gI7wq8aq2LFxdU6p09zAPNC12W0Q7ASRMGYF
yhWPU2uUOUu3+D2Odsxb1eGALBPOmZoNmSowelps1qtMooSMYWemLzB13+XqGPL7
q+JrH/HhCjhr2C8fJh/CYez4MRVepD+XJlqRpYl9+dq4H5Ze65kK84lTSy/cV34q
3PB0FoqldSBVIzTUZJEMto/DOm5WL5iCH1r1+31p2TUtmR9mEG6uMNW5xRS+i/pv
Mc9xhWaheJro+BzIKaZEjnsEiDtOss+7CrlVPUNDFY6WBXuD2wRKDqvnXAIE+m1R
jlDm2z3YZgBVrPl2F6RkxV7UnBhlkoaScHwndhMIytzrteQ6pw31JXmMLkdoHtW6
shfO7mKD3ci0O64R+aiu9D382ulUv2vJ60m5+A9xC/GSw6qBhFGkqBI1vbH3kOJR
nVI9p8w3NRJ/FQcAmlYeJNGIi+bZ6W9Z8qxoxiJFgJPRLbaq+PQeorU9qkO5ZqgI
GlYI09CbifYP0Fi2vPQy5URTEFy9MuWU7L2qsfC8GjzVrChU6eXdb0K1uknbaX4N
M3TFGascM4AtT+6AMZTB4rvVyeutXlYG5WKlXxTB3eN6RbsYoOStGqcfYyMIwR3E
1mLZcFD3DgTsZyCDB1bYl8OC1ZqXOQ8f/JyaylkdAAXs9i0DPBvhoz0BgnFPTD6q
FzTbMIjkq97I7iwbAJ5Byt3s9oAPTjxR5CNq+JzKZczkUr+WfmN7aXtrYcilVolC
yioYk3bRnM1H96mDpwE7onFMd8NMMXClftKnOdvpmgk8V4Y7Vc1ODk0Y8fTxafKx
8eZF8Z1lwBJ3crVyBFahQSYDEEuhsBVOderh6YseOTJdObVoKbS7MPRRRI22/EW/
TDpZ8M97MIN6BisbtI36Jxznko0n0hzSox6abASyzUTcpV35h/jal0qoZoU8JfkL
O0OREkS1vonA3/ocXkYKWsvn9KJi0dZUEsIeNY9QYZZoDzTVVvOYaebbZD+9WRH6
naJwEM6wAIezdbRzd/T21SKhiXhH66PQeAwLgZEorQjTYuB5feJQmdnuoK/Dz8A4
HH/ZRQPXFcJQdf3a/vyPq9+0pWRMSy4t3ypkfuCs4SsW971BQsY1Zbd0gyAUCran
eXP3d7GH0bRv8wsJ6PYu0hTGH02nximtBHDed9GSggFhYk+vUbYDWQK02cQGFUFG
Fy9hkbdMvGoPRkNGGMrpTg/5NLqIM/6Pweqm5KA6xDej/VulKNEMUgJ/w9+DRkHp
TYE2DkfH5hbhXs+Y9SoBHkrzWtxGL1R6mDi1Wp+aZ1T1tc5oCi3II9+qXOAYIurT
fPLECGcym0Q4ShpiRWU5Dhz9m7o6F/N31JRni4VDlq9U5g93EUwZyww/Y2kqLPXM
WFyeijE6hiylsPZgNy6OjUy64Pu7xpT7orSje5hoEFnftjJQf1xkEyWVzrx34m/F
YpgSuJSNe0RK+vIRYrAVIUfAvsnZx9Jmw6kK6nCLW2aDZqSxJ5y8+eB+AtAQYoX4
wTmtoJHa/byUygSK1HbSSYbra+Wgx95HkjlDOhvLpQHJf/fbEKn1IBtUXj1+vS+s
AcEgu6CaogNJJ4ZS6hQp2VReKWZaZyLDaGNGvzVp0sLLmNwoW+XVjAWtTWIUwSLd
/OuWUmOhYaVtA8x3JbZ1hUFZwjrNgMlKcjtiiMbn7nXD5O5FaATBauJHq16Wgvy/
+8F9Bw7s8vB8JSASesykxFgJAoKLHPmuAB2kshahVe4dUCzWT57oPgEX11K7uDhM
YtdX2uMNOLToP9FnLq1xUwvEGEmcBxff5nvuytr6g/80VgPS7c6NjnFOYFXEKWh0
9jkw0HmCDJg9DRfFLfNZ2pIkt5J9k/+2OTKwet/BMhRrplofOlwZTZpIJpNal0Cd
eZdU8SYmPQRhU7AAbTxlgGb/Oe8HT1w3ev0ji0rU8vwv6GD2E1DHyPhkAvRVY0QU
Vqxy9sRqy0C3UuVAFCf2kQNp1FKg3+kHmSgcU4AOcoLjf9CEmdV1m10rLQ6nbCug
T6bzOXDD+zXAkXIcFNyPxdXI7i0YSFlBS7Bgo2WOir2XPbu00MSozd2J07oNP86F
q54yYCTfNrvoPRF3LEojzrcoUKhP8B86AEWXYBzEvx7AC1/0j+OfTQZlKFYvuOtf
sc5WgOxGo5SeHF7oefCLe6Apk6zdfyX7iv4gY3OX4KBjsVZ1agmX5vkEKJg0dhzt
t+E3kDhyi3JPKUhtPg4omgLO5E7M9CW95jex9y0oVTIHRf+AJn+MBh0ci4gMOGCr
IX8SmsLVQFlgH2Xp0O6Ta1dJSp+xtoTyLSkKksEItOz9yofNabWxG/YTC3fyTuIA
hZQYL1+ijHfuijeRYpiqnq54H24fXtm8wuzf06wDetxQJp1poWwwYLyYkct3N+Zv
E1p0NzvsaJg9T+/sYKRUstFQccHHJM1+zjEeWby9RG3LCEVOyZZ06CBeipYxRm2m
sEej/ywHmEqk11EmuR/4GI18xbQRBMe4QvCiiXfqsxoVj5VX5qiElO3aktmUcxl4
4tH21qsiKHeE2qctwc/Egf+DWzo8yQkEWRZchHGRwdKLdtGL307QczaXCtbzQEPK
1lxAfSOm8NhcrR/oWbknJeu1S1fBX448P+Td11a2of1lYK8CENqCukTopv4NqUw5
XqSLsI0KVCBYeMGvUVXLTsLkNtL105jTC3IjA1CcirsZskS7HDKAFigQEp095Pb5
7knhtG+TRpz83mYtUKppQA3ND9BqWLqt+GM29y+LPFLiUNlZxQ1qCYdJx8LOqK1S
YfYyi+8Burw+6/fOW07ic7qdG5zTHoa+Qc9s5WdFFum+ca+2gJCrrPf7npFZU/c3
oh8Wl7dpnQrDP/k/9Slu8aESIUVRxMAuIDaW9fzpKnGanXSUgatEMES/9J4kgt3v
J2iVqaWwS3/m162UWkth6PaWBA+D9QxRKLHA5vFAO0eM0oPiIGMm8pRyRSbKaaAZ
NuFDk9HjefMnyPVL+YxslXZZG3meFx3UY534Rpc61KKQJPb6lI0VVLSGhr8KfNkg
khamlzFqTFkwvzqPrFWVvv/NRd777rB0Jdug7V+0iVO9PGikU9/+EhuQH5a/Y8sW
d4IAHrkB+GLOsEpM/pFBadeMecSpXTISKipvrcuxrXl1VACxDxz3iVigvtj/kGjg
I2VeymJbAoV8LX2Hi9PpGTueK+2LnwLgva+b5Qg7q3Uk+eKxx2CGEXAZje4YR/sH
0sQ637cnT9XpvD0Fq69qrNxl2O4BHjG+IxxjeKdK0aHkTkcxt+GFvx7k+HB9Hl2K
ESg+YSf1FP9lDpdhWVgZKDTOf2dzxg1TUpyMEDbQolkSVKI5T2xSVt8U5tx2E8pz
PDxvellQxGMzq7bzW4qp+dnE0+F2U9z83mhjtht3bBsJMK8Rf4JOh/ET3h8ioQ63
6vWR8EkDXYQK7ySrLKljGbyfaWfwQ+M674ysTlh24jtBFq5zA21P3S4NTLfPcGwQ
ym8+xuYDeLLku3Zpxp1uAWoOmqK9hDgWEFA/EZi7eD4s0LUxh+DMo5xodUD3Lfk5
4Szzxnv9W7qLxXqHNQe3RPl6qWnl7kr1btZV/C/rBuK1opm31jeUCZjlJLpPnQmn
Oy/8esZq+fiz3TvJ6WOJKIbP68TU7W7UVkR3VK6CW09SSsQ1l/iUc2w60VC+2jvW
e11Klto3OZPBeZrkIDn+2FoJlqugUZ1nSR97+H3T6x0GgqEQZ5cuqsFa+eIn+bjx
ZuSvGs1pNdstSqA7qFQC0ukKfgP1g+atGmDGaNLev/CV6a0zPS5emW5kXSb2c0js
5kALR+SBBFW+aj/Ss7/H4/A4vYdlwz3KlWovTfhr2viM2GovaDoCbrwieBMmTG7N
1eEdpFlhuppP6WpAVQQgjs9OYweNqRbndjd4kot30FD19W0KfTVcjZbA01xWrMn+
eqVO7mNOCJgF1IQ9pi9NPzv5pRTi8nUUAqdQVLnI2vv+9SOm69HG+er6hyqYj6xR
tSDToUJfvfJCUFAb4OcMGRLA68zQk1WYjgHiG19I5EVIgucwI3sJd4EG55PHQT0Q
eowIY+KUy14XKqykvJFSyNj18QDxk/QRluwKILzZNZSXLGMa1MmDhqX0au3hFhzw
uEUL9f2Jin+7M/7U97az4gACJjvntZptCx2efoLvrdPj7uCa9lsMMiwctU9JrHEo
FQWhFz81RuvYcxx0jk0yDwVTTzMAqajPSI98aPKbqLOhgS/tNzs9h9anJWQhU6u1
JgnNnY/q7PqH241dOuc6K2aMIXN5MOieiLoejjEZIAhyXKMC+Nv9ZrPG9RNqNhoH
MK4gl0WHaxpaT9DYgt7RXt36vh75DSFeUZsgdxzaqVyh1t97LDsDgmQgCx+TmHw4
QyzXkwc+52Kwunx/t2UCFYJdELb1p892XoA4VFKG4Byw0xS6bhXjdNHpet8j+wU6
zCasnItpXf4G+D7xe5eT5u+2dNr8vd4aKkzTMjsrviAEoMUE4+SnvCfLZ7oNa3CH
priIWad4cx4KtJR8tzv40mLJfbREDv0ibObDM/cba88Zd8DjqAsDNAZNy6IrNaSA
3YVTil6vo7sDzYacKjupb/aOnvuHxnwtOgTZpORWC1HNjmqMmKv8HlHnuzoj5yL8
olP2TfXL9LX49RyZ9yCvqHNuFEpy+OB1SYR1a+ZZmZwC2hoOffWbs46iCxvDIgfq
MRwogarwdD9KTF+zAG3b1sWbuXa9HYMBUL4GPnxo8R6X3opMYlGAs3OTA6l7GvmY
1tjh/q6b53l8U5URAvPxfwVT8C0bFnyRqKqx6ce80lYTGovvu9k4FS9spgs5O1yE
9usgPUtGidLEAlZo385FOyBi3rxVDpLOBUGLhMMsE3BkgGVofyRkFVnWmym1jTe/
88QbRJJwnVYUBUCOFZJZMnfcYxIiN8PYQecGZS3qBr86HCpSSk9qoVDxU05kuvOe
PwjQPV0no8+9j0+B+bpr0Rc46zJB5lLyAGb6igWRsIgKRI1ndC5wAxeny3wMPm6y
8MUH5pCWrxEiA+4ZZUeIO6rihYNEQZlbyFGrcYZ5AqYizoDt0BeJGQ9+56F+hjY3
mLrD8We0NGrxam81SJRu0Bi5nAigR9HNUtrqu0o/BkPqeUFC6WA6imT+co60cl0o
mI/SGeY4Dedv/vlAPkoiMR6WNkNgKxgSzh2gu02CqCqI/YCWj40edB5E3/r1KqgE
vsnF0125NPhv0D1nQJCAlzeHOOX7LRIRZvDkjOVn7qIxzYREExAH4YF8BmLQnO98
fd4RoS8OGeRFWdizsvOt7/2pnqhj4mLg/y5SJ2KmGt8q+N2u61X1YP5Lx2i73nZh
g0g6nKa0E09SbyHwm9ht8RPwroUMVuA829DrBPn5vLvuDDiHsEHLr06fkQmIpT/X
p3s/Ja4QpBKze9s7kPrRvMx0KtDPtIXD3qXCwNKt4TIkUlfHqKN96SGk1qJkaex0
b//pnampHlaSuI1uTX8Sae3cmko25yuhCTMdpGLvVfmvrpmJM0cHGl1/g7hdlXTx
UPKyCJbC2q8rxoGzf+vvu7+JIeg6rqY7v4GvSYAWETd0cveDNLNdxH6UqUFBCS5v
He79aTm+ivUxokUg9rlNmhPaWCLNz5AQEKhcBNHLZ9voaXbN/PpcLuAZUmefofZj
qe3pbRM33s/xVFOrKHI6I7PcqO6rxUQ5lTH0+NGGsb6Ff2LMh/1imjKobbVSF50k
O9k9wrspxn9XH3K2wJrU0eNH5Ev5I1ZyHefagIBSK4CHR2yb6wkVlJ1lKiamab8z
n2gitc10Xwof17A3sm1owX5DP9kC2/kkS/lZlRWmcAkkX/ElJS7rYsIsGRDgjrz2
ucYcesqEzEfCBbtJwmvTyV+5ps3z5Wm15L6QyeNFJmxUeTC6vRNblRhaa2I8LbdE
ZNy/zFw/SRIO1qlYte9ZyYn/45yE0DmVEvG/eIzGmH467kdxxnwMNU82RUFgigwq
jH+ckhiBRKFghZNFdi1JbPJHa7gSE2yWaNkRhZBWwWgn7fATUHJ5KhHMUx5hrfe1
tgJ69nUTxypGJqIAkBuodg0WyVVUm/av9U3OtuEtbMnUWx2FkXsFetLQm8CnA9Xp
rWWmFwzVWbBw36ZiVL8hFoynGVPeArSnpvfpUdEcDG2f14IclKznzaI6Lx+Phuog
yd+/ivUQXZWf1hX0UCNaMfCcRg6F/T8y6x65fvmDvlhRymA0JUt8AY0TRFuDxJ+D
xSSyfkRCBm0cZ7fLIZKloWccnTos/z9PWNiS2eaQ4ADro/7KLjIinHAvCP5plL0Z
PrriZadaKu0wz7/BfFLg3Fmf1lSkOk/xJdFJhDbCZ+xcwbCJS30BsUTs57MdhiNW
BLu2rY0CJbftbnzGMDRfW3lY+KvWQkg6wRscoGBGolWOVqioaBig8aIRHTMKseyj
mBuSCW8u+wG9QD8az/lrVfEMmYy5e8x2dd27/3JfdICv4K3J/SjUepirMY2yjp0R
zh29t903QPK9afHZc6gcC9FWPsSzp1C1dyPvpTw27oyRu+UPPAMk0yWKCAAZItr8
pz/bkLz5zcSBQXruopLpSWnj9fAn+9yn5W+N4P/ZpA3fU4wpmKgvC/kUOPlcui/o
sM7XEWV1orVUGjykQcYDFV/ykWMfmdX4kgODy3pj7PCG5fH3dhmk+60UkjEDVTcn
ujRKVY8DTGXXC4DDsuzJqmBa8rYQrIYKxPw5q6c50pUBJuN4heNjjfRfZmUEbUMQ
ZGzL2V8gZ80ASxygNJsaqqw133tS8ss+g8NdCbSK19uEtq3+PAngGubBBVjj+YZl
e6a2bosJuyuYaMTgjn+2QnEVqOzlaoIECtC2Wl4sgyY2sfvXzzYpfjqCzPNquHxX
kmAG5/KFg4SRVKdefWi2ELasR9Gbrd6c6h39W50lnf84jJtCE27z6SW8o5h6gRss
clKKPN96mPQJIu/1h0bpeFNy1tdb2uECmZkNfkWYpCqETAWxPw+m6sIAzxhXB/gw
hmOIEVtQnPmz2JiCr4AHgDHXR7ayZMcFU5H1Aiv9YiNhqeObqCpYnHtmSuCTBAaG
tGJKDzfSVV4OQH09tIFtmuoAaXoxOJzQpVpDt/4/nI8/cNgX9Tzs7IKuwRHWjQSp
8jJnnpAGeVzfiPbAVheuq6Z2jgHKVUuPtKR79o/6KzWlcTZOGbda5FFlDxQfLIO8
ithwC8k9ZT6RLngND7T926RTVQq4XDGRxbtUZaQQ0Mwj9QyFqWTj/iIkZ3fPX8tl
lINlLS+9tGQXww1cIJwVn0cM84xuerGg175vZcz3UGuNt6F9Og7GNSwpM6ujdTis
IPtGoDyReW+CLejHUolVggaknPv99jsRXbjYGqRLzbXt2uq5/lqLzDG8M2dVr/iE
CfoBEBQhYzrAW2x0aKB3v0g8r624s8xwgVipCaf3Jeg4ch+7q1zg0g+5LmO2Gfy3
/AnmF/nUGPqK3ZCKJYqpJX1pJDtnAzf53BAxIZFGNSnraS2DoU5/ODd5a+ILtvW3
J7OcEf1aXujc882uQbUgKDo2X/Qzyor5AwJA/iwqaZq2B41pqs4dAWDVon7fnBRs
wi/Q6VtzKXHX5ovRznCr+oscdON4RTvkiROG0Ktfiz/1ViJri8L4OUNnzG7eCMSH
X/zzMm6dAOgwpiDukdK0DCRWfrFpIjKdpytMI/ruZPwMv+uTxv1SVloFoftmBXu/
TJb645IOPhFiQLlE9PPMP1lbMRcosUt8Tl+qtg/ie2vOygg9kaj/gWINGlczon0o
NuGFkh+byH/0j9/bIjDQKzltQrpZWrIoUwj7Btmau2RUKO/RZgETf53R+09YsCwY
Wi6rHt4pz83SFPGbu5oQz/9x0/ni0GhIjRR04N/3xVpahN5Rrzq5v7O+G3Oe3+/m
j3lg2TIVKdgJM6O0xFwUgF0cUhsUT+O0exrM1dWsdaytPh8MgR80Po+ZgMrE2AdQ
cHhUQxHINdx+Qaqg/q/QB+a2xVkDZoOCQm0/hV4ke/OVIrjxB/2fLB1n4g1bSKUf
ky8jiq5H9kWo8CBxHMRdDkU9kbcajH8OH93W5HHWNiMYGCqWo/LAlPgoyNT3yAYr
hHcYJ/vHDgdZJjnzTP+ldXZGGJd3dInc4IPWbwHJ5JF23GaFCDEyO8nLhX4ER39l
RlLtvXQkN9Zv3Iqcx9K5IboOyf7JdjQx6at4lTIvu1G8SmSGRA51z/YBAD3xJAi7
V6Yfnv7Rxa4O4VGfqb+jLQ2WD6NNCWor0Mu5tPEVyqGau1ca8tRCl7mqJ/uMd9yK
BXfDi1fGPbzlNriGWusZmQ6bFe+KtzwNxG47Nf9VcFNiibHq7fYrK45piJqlOGbL
9wDbnBOg7Bi/FQLpLU5AGh1LAFsHyr4+BxzYjnMPHgWb8K/EKQ8gZHv3fuYy+pas
hGfARq6RIx2t49nSBf4ehdvGL8VZwapIhRTA1pGndUTFRorU75hy+Q6yZnKEj2nh
WlNl7VWZyfvxLWtJ44BHPA0EeH4tN+pD/S2KH3Rkh5P688CCgFl1qiRmpHEYjRCt
vxy5VvZmac/XvwZ29wrq/i8uTQxt/CVkF4+bq0aKp2oX8Yf0go5qz3OEhBuw4MNK
P5rTKVq9fblxhbvdQAtLfsiRYzRY0c7ZMpjow/Ph5SPnhIaRx8b6+WlWwXxXzQaw
BDZE493GwfJYxAocs4/k9Z4RTvuca8J9Y5POgJsOJCTZaV/nIJ6KmF+ZAboIbsxC
uJQxd+W5ora/0rFH+0nssmitLQJovTngJHwR59pN/y6oiJYImhzeyui1Ybd9nPeX
i9rF74AlsErz4AuwfY25l9ZR+u9sInukwj65KRlzJfr2fDfZjVX+SsCj78FpkuLk
OlL/qP54QXgpgjSfZU0b3V8OQ4/FPUsigAJq+gecp/LODCulPsIhrNjusryLp6HB
GfXzrPFfvJ8wH2BMyoeBT7nz6aaFNxyULLyUetfADWrf8xbam6Pz4yg/3p2vt+Bb
EYFE2/jHp+QDcTwLi/JlM8WGvTuLW8qE32cehAz/sQ7tmkpTZxmmfAj6iWkL/230
Cne10ntuijsRlyldhwmm2why2nK8aEktOUKLvKorkOlNsCL5anCQkKO8fKxVDsbs
Wj+W/lMfe08ZfY5hU/+Ot12xOOtJpq3wmbGvIvmhbVa+w9J7ofBMok9kw3QAZB9/
l3D2KUtM7Xbpc8rzeFCr+zegou6nR8ljTXbNP67Rd2yombHucIlnPU0cMaTDb8NH
yC/Q6C8txaaLgzSFy+j87Ftlo8FS/HEK1Cof4X+kbkSfvyxQPzezAIvc+1pJlXwi
/gIfoDYPYUHAI7SyCwJC7tjUiyutJ3TGtpg36ECzVBcfdbIllkHuGnQa3+/ynHU5
JcwGgPEKeeZb1rW9ssrun9OnFetAxqVrtzyObIOMHZvovEwKEvQYi3/87fj94sa6
EfEoGBM+XFZNKrrXyNtgS84GFmbS2zRb9SdxWVKE4lcCIJwu5ccTlIlGxvKc7rNP
FQKtkPrBRFwYQsTw7gD6ijuszNgBEXCW3m7Sa9h3sjwHCnfqCVDLnei5W2wtshYt
xHdipGnR8AZRkN9SmkhxKSaTAQictWwkLb7juVwPznBOcgjQlTPFhO4z39lGvZOI
4amTfglhWzM5ZvfwAFOBJicgLyQ/j5RN5ZcKFtxm3fMECIibkCPlF63VC1tnG+00
4MHB4u7N95k80aQl0nPczpDBukf1MX0K+Dh+pWWpaTfKDXYJkLpxQ1T+zr6XpJY5
BGUHO77n9D01nK65j37oE3YR+yQfB/ocCJYypqWryCocTEYoF2BOkFKfkc/2F+5E
SFo44ZHc9iM3oozJ/DaEa7vkxUhMiBnnPFe+MWZt7Ms0wh48K47+qVASzePD/FA/
u8Br6Ag8RUlitW48zjkqZzr2qugqgz61f+csVBs44jU+jtRaa0gmrQiYA5ouvcCV
hPL5GNfFlt3pKWoWDr0L2WYCLV012wMtwT1Eqi3v6pP+O0tUr2OpkCHmlibjXvkG
o/797SR3HpWom9RL74r8e8Ocn30EBJ13aPWsgKF3bZl7RdC83ddZ88kJJrug+KRv
qSNlmj+b1umMRgUF9Y8DXL943xNq8T5580o+2yDmap4NCJsWO5YwS4GziDjNVgXW
YTm2wPGISGbWULH8zJsJZSE4vPcGOQVK3jfndW+s+FzYCrhuS51m+KOVKEo1TIT8
bgzjL8zXjpe4RX5oHDl65yrs3TYFdNKNocG5iqTLNLQfLHxsOtc6duhuxlPIFwux
/ecv90rHpARmOqu+QGdaDIw6dK361hmWTce+AGe+rThsaAI9ZAzsDCIGZRN8o0h/
sCJDI8KCMsEd9O69nlrU0voIY618amXTlXq0ellj2VVFDFhJnz9Mz4LO1AkNINVk
XOAnsKsEm7AW58uYkT+NRwAOL/sPmsou2pw9A9VzfjMUk7NJHli4/brXlCwQVnvK
72OqevGmHXQLJl6SrRC4WnHjwEgwNRnd3pnN0rEEPvfytUpLq+OB9P+KjpvmGBqE
CPvEZZaaqcvv0LK5bJGorirWAylNL4qD09SW6kLJa+DmFALhgW6poSsq3iGrskyV
Vkajb7eHMpE2Brfp3hiCAYL8m3PSlwkfitA9TCWaxCT07fNLU5m0uqcmoJS+cSp+
npSPC+pdQCSFjLJlta31u0vCXpgE/fcjjAZ9INettNk5SLj9bREpyt285sAfWWzi
aeL/SIp/bQMS0FeHbI0ddh1R6p88PCEEYjYE0jkj4a8M9suuJCFy3MXGXP+f0XV2
H1NxUZmHwolUwMFfylVfZrBnnBKMalSNLVBh5bHxUCGzRYGX+IafOFP0Wike7mTC
+EWIT4JNzvWuhosCnMzxBf3czQuw34Nhq+88mgguSBgGeFj9/TtXPEA6sHALdGwH
+X1NB4WHS/S4bYjkXVI60OwlJYYdIO/IBDAtqO95YbJBUQkk9l3fLu46hOMxKYd5
0vpV9xrWtAs3Bl2COHGB1us4zpaOzeAq7UyWU8TmFEW5REi0HdSOZ2Y+0wzUcNNt
g0m5v9/neCoTV+k3v7SGH6uEgHtS+/uIVrcRVFOhvCVA8o7wSudA23s73Hqvj9zh
Un6aDQ261x94U/ul82y+wzBYIhb9TavxpyeAPd1QwOy+89DAJbRUetwULX09IWqU
1YLrGwiVLYXxSBSwPI20ODHet/mGNPvphXSoqEjrmrT/o5uDgoHhvNM9m2wcEgrW
wlrsNtngROkY2RfLANAuJTiZaNdrONDwwWKyGaBKjjseSQMqYacjzhesDTiJFpM6
xpb51LjEjHH1oF8noiRq0n+sPxBoS52L97mIYtTcGD3l2EEAMyYtu23PU+P1Y+Wv
UH+WucflraDPHR2QA/9gP6J5Kf9CMVhdX8npS8hAmLzCfO7LQwacWX1fBdHXb8tW
x1Zx4WG3bI4/m3TrbHXSAYF8FxCQJqTfsy6cIL90h+zy3512iHEMSaX6oSt6pC4I
XqwfdBXeDrEu5dP7At8xwoIHTQANsV8a/F7WiTeFQFzXAdCi913ng758TCqMSanB
vyZmaPZ9F47gIeYHRp66CR3wyVAKzHTdWF5cf9ugJbs7Y87GEf0ar7Wn3Jmt0gtZ
kLJ1Ro/cT1Naf9qiCJ9RCiz6bBkjowo+ed6EnUhJ3iyYFgGXb3AJTFpMJfMD1wev
oo+66jvx+RbEZcAZ58RsiLKUHX4nnKTTL/cLWp584zsdwDHdj+sQeAEm7afb89+z
MAToMMRYtrn/IYdGrE7gfLooRc87L2U9BaDkTb2LBgahqvhZM6+XogwpTEJnj8kb
MfVXccca5om6FW9TsUYqyqMH0YwubQ/p2zsdohaBL2Ec8V1doVMW/1ARQrtjDX6M
BuVQZYxV/eeXFPAgTDQMGd6Mj42LL/GxU2GZz/oTbzSA9BXNmj6ByzwM2WhTplpz
ExiV76BnHC0BeENh0kxUcB3S59poRHEvxvCVsYDvoT1hvCgeRlDSmafcMl0RvPRT
RYCxh2vcSgyGO8hUDI4ulojjkFkeKlKf1e+PeeyIyv8J0T+S0k3HXp/Cs9FxxV2D
CWLBQF4jW+dR7W9DQzpBuY0+SXBlydmXrTF0PVfVpFs0kd9iSK8GrBLTFPjpjJeU
+jbbVokaeY35ZUe1iDIDshtw/FDkuku3kEhmzlqkC7v75q6aZ2zX3Qw+bRzzJTrK
p4dM2WwIjTP0oXFsqc1Nv0WszCfCKoNUHZKExG8f3O9t3Ab6g0F8lvM7Aqq3U2qU
pyqv8NE9wc8cQvlij1W4QLfuaeB0asJbpAzxDzlsc5QXIw1dXeyqERM7p1TILPyu
tWC/gWt0YwrZ+ONaLBRB6DvQME8FYLyccO8bsnT8E+HQou4pBplA1sd32dx7wxu3
tew68xm4Ib2ipRvhz68TXFffui3GpI0DXLcg8KH4zfTRbD0KjBksGrjHgC9+CxEU
qlgyw/+YL2XefujNl4/hC+eE0d+y0ZN+pG0Gd+sdvPxbyJidLg4TwMbzBsLJSzV7
odcuuJs2ShZhWnTaYp8pfUp9xtoo5uFVya+KiwFoehNHndJRRQsySDYuMi2u40Et
Q089umgjayfNK17frF/cQJxmT04d34YVV7MGdnj163p+sc0H7ld6wXAYkTnZ2pVF
ZB5ZsnVYMh7Hy0zBDI8H9RrWInOmMoXu5jp+8nnGYjczA/uy2W5SCMvUCXcj3+HD
Fj+goyMZPzsaEdau82AbjpCUlZ4ABUmSuH+Mcri8GaaZyrg1uJMFjSpRyp44kayD
bDksjobvKDJF8GL/CXApxqeCv53HfwafNsCVK4kzDPaMuG82J5Rm16ILXiFHMYED
Dvgwbf/5WWC+O+cDcQWr57oaXIrsnpUUO6S77I+3DTI0QpxLvsWhrAGPo5Do5Pkg
Vsnrd2nsRABu6y2KuXkPTSuUrZUdHuWMo0XJQmP48u+QwQ7eBKdqJu6DUJ492jYL
VzmOtdAMTqT7x+zA6dvDarUlMm3KyxdCgqie4SjY6YL7ffsJ2WGsMtoCJcQ8RnTU
Bc/ZcGaUronO93FJZ5B4noWtv/fXVuQorKU8VPNPMEHCpcp87O1LW2nXEhKk7zHT
cvMpDBaPsMe9AF3SjRcfAJPiXyt45hxnE2Ye00IyoBX5IFCGzwB3SAR4heZ05Lbu
n9p3ra05wTpusbBiCmX8894/Us9N09WEAcXcx2gYAR5HyxF4t7Vr1dSAiIINsl2l
+mmDD6njP6spM14hSR0Qq6wWqvdLN760SyImERDh/RNmKU8Q+GeHPTxZaM7c1gxg
U8KCyhsGFIApQBw33pRsypnEwOSJHiGwEx5VRMOXe1ziX8gf24B9gxKKR1g+9su2
Ad53eZMaZrtxMvCPHXt9JL8EifPnFwGd2gUk0+r8DaYFPa3RvibgvvzaBenzzqAh
Mk5vAfbkmVR76waVz1TD9ilHnWpZ2mVOgllsmAS54WAfJhXk0kaOtYD0AEJijsYv
sJ3ckPTHTObax3mEUpfwSYfYo/n6WMD1YvSVTsr03ViLgdKDzMQU0//fVeDG2tHj
Yd6UNtJB05ZfjADe52XbXPoUUjj37bjl4kdhIVthz0VcQ5vFoI0PQBSwyPlWskoC
JAbdwRl2KUuD6Yeu+R8m5OGTrnAwLku9Fipa/+9CG00WIsMOFIjo0tWYyPnyMTzV
J5D55lUF8AFcJ0ONFB/AaozP1cv13cX+VcurVKqf+Y653Oxgk+NTIYTwdlUYfUpe
LJNt3xMyOV/g4K/+PgNCFE5OzV0C2MF/7/9f6jy+xhLKWDLibHbZFzOTWA3CISXP
`protect END_PROTECTED
