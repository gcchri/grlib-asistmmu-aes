`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nxaAfV43phFc+EKexd3Ge1Wy1wjnp7rBCfO89A0lmjvQhnqBbGzkhdGUn74Y1wBN
Dwma84AAKzEN9vWyQJS3XxzfPvAroQf/3XiIXfkmBHinVeYmZ5bhoHO7DRi1nvK8
Hh4mZZdDqv033jNGnynn4pGi7UYxd3V165PgnknhFPgTxFuGvUSpv1ZpMxhJjYx2
/E/NrCeRjJ2M8clusrmm2qdSp0gjmuQDB3ka3HSP2R3XcZ2w0ry810aY3oHvQIdV
ACuQopTVJb0n0oDk0r8yvwGkmGkGWsmn5dEVJT8kXLkffTCcAmUe7MD96SqeNmOx
pekMzTrRp7DEeGaEQ36EhuorkNCmDezmszpQv2/FykKzqTxBEmLOnyHjCzvz6W5D
qhsEvHJoxlfpaeeDrXitrqbofz1WlrzYz/AkcpK+C9p8k4jKl4xgFtnEc3+vX9il
psvtZnhXp4v2GOaKDNmYMw==
`protect END_PROTECTED
