`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dA9uhJ3x5SlSRI+y3fUJ5SMEAGHKIB6B82M0KoTjI/agLP2paLMaMMiT/81n6QpV
EEWCXiXlDOdmKlKZChztAnmQdJp+q7VocuILah6R0me4mGedQqVuGrf2UXBwQT5U
mJc2CxTer9oMmYTFnq28iObDvdTL5bla9UvIGpSZ/vDoW9VJBQfTo8LqXsnksxiq
TjzixcgNwYr9j2ru4Fso/f4nlVYrXcO+/jO6pqyVKjmbvrT1ejYZcNz99+q6BCG3
DM/ARmS6cDAmWwdUQt+OCACGmN5ttThldB4MgLNHpSn52/W24p0PGL1PQ4TwPYRt
VV4iRJSq8ue1mRSOe3dpT6zizbzUZrKaGCMvEHdegeQgPY7mgM61CWKFBzBjYiGn
ix7Wtu0EeSn7C1CurykWutYVl18tfLHle+/+xkXg9VolhjXB/Vp4v06swdr+EZmA
GNtmesWZ8LiJgXnXFVVYUEXuuwcG22t429oDcnoiJpW3IErMNMI4k63/yirEtxUt
xQcIkM0pBSkM9CIUhJrTn9zywY2Yilb2dy8wEQSsKsPkp39unEG9AXqfVC29egB2
9V1xCMT5p2eqH/peyCw9hTzCSVDop2O8ZfqA8hJfpwU9R/zEA7ipHv52AKAuVSRN
5hit3q9mZQUjOaQFPhzuVbYGVTq2zW7bprO8F/uGvo9rzUCH1veVmcqhG6vzng0q
VyBTGOVGc2DB/IQYqVVN8fhv9+JSTyGoweDxViBGwdSzwc/PXth0OvNhXsV17JL6
9Do2q7PZcrXntSTLh5NLom0FV9+nJyVaVzwocRIlhJdxSVNBv7k29ASTSRM0VOxF
0BeRc98ngB198hWxOJWbX65ZtIV5GwcQiKmnHDPpGZVbwnT3lnLCnQYQpZqj5D9q
/O431qGqBylXSHdsBmCtKwgHM2Z4EzaI6P5F5Boc0EZRT+u9B5Q614I8b4K4du1z
5mfG1FiQN7FEgYaclkgyGsC9yGi3xSWjye0Dcr6dJ97fQcHC12WI/UcdxJ0Oh+ws
hCAeudL9fvSB7cU/LeweN/IM7VjEBIIn7OccRBHnCoDM0xTANwwD1oIea7JcVSo+
8/UzQYB6AXmrhDrHHFuZk8zHvip8oMBuV1xPzBzDWVk70kohsf34dIRyF3Ik4dii
N5O1K4rP19YW+6WANo/fmU7d44uo9C5Cvzf9B2/n/R3UQotn8qmxzdDTfzN9f+46
uHdNfBhEdYJlqVckOpEw9c4s09AbN8M9UycKakenyQNIvBWgvE3BGYIWT4E3WuL7
vOvjVQ0PYVXJD8yo6EnCplYkSnnzg0HuJo4CzaX1MefqrOeb7zflrgWl89BeK7Fe
0iDWqG/ND41zZBLm2X5dth4Rku0WreSOKLU9fre9oDornhT8LcsQGPvn0ZPhSSXt
e0aFrKdv8rGAFLv+/njJzagnlBkINM5l/jS/3w7swssOhAngaXd3q2EwkgHfmVgN
VRhOsq4bmsZjFReRsnE+PSoWHr5WhOxdgdPoaR6hloxWyFDn4gF+EdW57iGEOn/A
CHNJk6ZuVL/vAIkAtm9jbbaKQqTFTFMILCXlFdAcJ+i2WsBK0k0HOTL/nUXWpcsU
2pH8rm4mI12CGuOqsGzDkgEduY8DhAAjv1Hj2dYpMQE65z8z3R1iPTLiPRhbIbbm
OOyGV/Hy8Dv8tfBW/QrFAb1jwFeLjB1j8aXfQM7Le4HjFEKFm3B2ue9xOFz14x+Q
FmcSAJKz3CoN6LY9vRiMXGP+t/JiQ4qF3UzD2voLAefIU8eVoDwOC9KFKHnUgGab
5otxn2VwkyqGpYZ3wRV8BQI5Lq9a2vQnvyD5UAgDelIGu7fKtgI93fjbZ49hUv6g
Cgx6KL3ifw3ArsNccyCuNgW64n5FHo1lI0nk1wSlxtViQBjIGib9aIIGA7qqSi7T
yfjaQe7wQr+ibvjDxRL8XQWbCg8L3DkPHKvV/ytKIA3KkSg42Qbr4MTKD7hvu6Pb
3qWq/bn8Wj2MykD8UaK9oPhm0efRyRSYPXJYik/ShUMM7lQZCiEKDiCddlGLm+lC
jqH0ZvODzdmnvH1Xunm2gvi2L2Ol+bubXTcymv6H0xfbgcKT2UCJRexu+FYR6BKj
zQIfRBFE9Ig3iotg3gDdji6uzYwgvBGAKpe91fGj06zh/omlE0Wh4ILY85s4GeEJ
22AReZ5CePRY/LJnDK0fMpBUW60HC8Yb3B2Bi6wFFNqGilQVDIZHuKSswdMpzs3d
t/dyameghtOc/MJH6eoyUcsyzFK4DM1pe9rndLfPNriDqYlZVy3QS0ulXwNQqDTG
BwZwbTTWKO5Y98QKsBQmUNUYpTpbtxNmpFMqJmcgY35hNIpyMqwupywYtNvglx06
JK8Qpl82lkC1FZZZgbD9afqSTEFbvpnSyjOMnbd4PaZiVnt3ho5L/5zTbTJQZg/8
4BrF91cqchJwtudxHvZbWpScGgrb19qqqPVjX1txKp4XtJKnD7aF1zLbknu0FHI8
LMIpvj1drsksQ53ncEMoraSO4oDgTgk8uiwGw6RLmJPyENggbiCt+o+OxbuhM5Fi
sstSU+sjSOPXEglzYHaSB+SlZ4/0QYWZ5qfvq8P90YKjubrL7L0GOY86psiN1RVx
HjSlGFBDBOeTeX6HbiHhh3Ulc46/EOEwya9D60ET2LEi8S0Y1IAzO6QFi2OQy/hM
K9i18UmFrtw7YZMGYqfCUuTcpTjmtTeHF6Donp1s0Z5d2zsivs+v6pKTHbEYTw8V
kUA/ubhPVlrpwojVCpvy1e72b05PB2rz6iHifC/Y5cs=
`protect END_PROTECTED
