`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TOG9Zp4YtjtzYO/NCJTcgPt0kNFlLWFTx6C7L2SDG0nJK8t+IbHK5G1l64vJCtlx
geBbyVDd3O8nUXF++swmtUfdhFLQ3w4tUbkG/EL5X8a7BwsB4tUpwFbVsz47zGnI
yDnBFp/CQkY148kAEVAuIGsB6LBWcrrqg3hgO7rudeTcGuFU1fv3tPEM+tbzODYm
uYqmQPE1gp61F5LmD1/zQ4ftr3sCjtUWEmBdP5MQw2mK2UT9Z6/TdHRslqKTLzAb
QOt0t9jeBG1BmcCe8FqXyAYOmXu5R4NTQIePMjm9f3wzI778vBqQGV2575nVdHPD
oag6AyU9HSQ8SO1EWixe4w==
`protect END_PROTECTED
