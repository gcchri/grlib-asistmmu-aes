`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QB5PvNEjINRl+e4AsY0Pd3gDKE1kn4yB3F4Euf8ql/EvcEmRNYtUw1Ed6DfECQwZ
LkA1dnU1WaSwFb48wr1UtExUAA6EmwFuihvEcQ3GhGXuG3Vx9HUkIhJ/a0O1sARv
KImY5+5HvVdCk8bgh0ztvnfTTBlp9+kEYyfbVNlBIXzca4klOZGzPm3ywtSuc+Zv
sugIs05YCooyVhCPIX/2RUU92HNtXnuWMY2izsPUBVl2j9zKVTsPJ9wsmndcpwjI
6Nsz39jQkCYIrvC17Ojux6X4RF3ucydZOizYxqwAqz/owOc4nNWmbNHutxKqWfap
xfWuGFZqb3uqQT93i3hq1fXnATKf2fBh2ujgV+9SyVPT8eMavREEptFHfgQh+JkI
oFncqSfUJMrdHyuwtKSke6mUDEhGk/fXlyxHrN4yzaSmVKROu8kVjLmA0GvXkPsF
3FSpneCjK77BTAJSODc4bngjkutD5Fj2PWuL2oAU1V0=
`protect END_PROTECTED
