`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vnEkipLF/whw57lfScbp3/Rq+sNKWpSBbtcDQ1EV5nPVI8U8jt5enkolpew70v2+
vh0gXw3/hQaU9R52GzXqm4hJ515MmTAu969Wfo26fN5dztc0rBbP8Ov9SrSqWA0a
bJstAWRlZMPJVnCAb39CJCmP4oPRPamy9r4pPcTqYBjOvzgYwuwK4JGQaF+7GrXP
TOLlrZjv3m6MkLcY9uECm06lBj6dS6SjpIz6UrRsdygT/ZSkMHd6h64L/6DwnY0z
/ReKa5BGEASjUXeBffyG9X/PmUPtWWQ5TG6xESzwtMBnklkL9ILRRDFE1HTF6W1l
ES9CnJP6Per019JqGzP0uKRl/SroSKumqzX9YEf1p02it7Sp/iEecOJOGqlh1RRx
BQrU3whQxSDKxxz1ai71FbIbG96s0MLPgVjc3PBwM1nW3+fBgShIeiPyGSelgsht
Hxdu5QZ93Z588ZDCxkeGpls27Uz3VSoLyof0RB/REaWMsWTvhRraGXP5ehgrR2rR
FIfyWTEsyeJH9Qr7VUpquiv19oCF3kIRxFq49cSxSvtDbsepWHOFNWR2Vy6SB1eE
7/njZ0mqTmQIciBtpUEzOxA4WtmVUCickg8VwPOyBBnXTj66cKliwhbB2UwCrsQ2
taV7bGahzcPrtU69ZrE4WWRyYzw+xZPi7J+9/OysEoLUGwXouCVS6JhY5EfnbEyU
SHQhcHSSU4e1cQJA6W7eG03S4xtDY234D2b0Q+kBc3+SahT6AOGoGsK7f7vImtA1
rAjdbxePov/JcY0ChBaPxAL/YPAB4mpGvMzJcLVjHvDpvr+KNd3mup9KRS+kQXiW
zxgRZc7mCm/1rzUcdKkmC049Cpg9BMaPQGFPjLmLrXvgZUbrQVqLEt4InYnBW9U0
MjszVMPAoIjQarNN1m5twH3hhCtIOTkDTL47BdR6koT+Vm1/xlWh/s5YjOEOeHs0
ezzacLz6R9JTTmGra3J5pk31WQRf3h2vrQUM9fm0/zwokcY3wzvpN3dpjcUOSXXM
Uo8Q3Q1o9ESeKbbKXYkYxgZy3Db6Tc30b9nQ6dfAUkKBQH6na2GlC2tUA2i2Ig09
ocrHz7i8GGneCNCUojEB2sTl1mLkcEEtYRn0eCF3ASoJx2JoVYSs2hSQoISMGZWr
nlQYS/waGhIkByTvfhrJR+x9tm8W4NP441ys1LHW3vIb4/kOL5+/q0E3C5InNlN+
7MlkboLZRTGDYWr+DSiUfcEblo1U/eDNXkEIN2VvaFOPAUz6ygORVuuNuwmqEciR
7XXAFgbfjdW0nKMEVQwsNOdhI6yaKxEIdrvCaQLqLxWQKkkyjJZ9GyrBDrFoknGq
oiDNDqkHgz7Q6N62nwWNXD6xVy1lexaFVuCOLDh3NO+aJKdIEgdVCsY1PfwOhriU
kG5KfknjrXvZtB7A+RCnge7jNp6kEEp4VYO1SGLVJ9PZFGM04fIYPiljVKa5R2/L
c9wi1XtLGczy0MVzLGFXAyfxgNvw2WhMYNzM+phqkNeZWjkTm5Rj3Rm04YaExCwB
wJ3QRESSIM38NF+ZcIAMe+LFzTe+B1DoPPLThZlwaWZAihMUZh8f+eIRp7pT6USi
LNe6EhSfAKbYG7t0YMJQ/J2eW0AuzAgTleSLAKlUql55z5vVs866Xf9V48taDuAW
BY+2lhrDy5T9+e4cMmfxAfhtal2AmdH2RM+uAotoEpMQTN4ZX9sfHgFAT/V9T0p7
J6o0pRpBjJXK7EtYZoBGMIPRkcCy9Ivui5P5GziOYsUTic5C7l6urAPZG29N9ovm
LrezmUJ1vuOZZrrSSaQ94SKmTFeBu5HHfsizhdeZpYwt2Ddlsdl3AzeGTbonK20m
xwBL6VEj46LrlUJiZBnWmu25+/8Ehc2sBR9NZwYJILVu2G8My0EC9dJQVCHr6+Zp
35FYWrIQ2JwSjcXtTilzNkTHdCPv+askfZRDEeu+cKCfWuY35A2uCYCyBDQmklS/
k51yzy4nhd0076ESER4XMP+TEEMzGAEK998/I3lT1U+hTFy/2g7qFU5tEwIv9ykk
Q4E83iz7E8q8b9HFY8hgyMrJfuxbs6gUXJ1IYuuhu/Dmxau8cSwU9V/ByHUqaCBg
6GBokivGamA1PuL2k80fIB2Q4YlM06tIXuc4umx52yTCTn2BG3PIh1D3sFa9xZpy
uD1SlQF9Tsyg5QVJRNpLcXVxg0krUtBLLNWqzQpUEl2AdatCcnWnjapfu7xR5T/E
4g6H4EuohMtyPfshQu0LJ3SJvy+1LTwk9D4lvUrYbHXiaFCGTxYfR4gTcn10rA+M
k5lGMhXVg5F+cy+QAXul6fbFZ4K4yWTAEIsr93envF2mbnnGgAP57pe0xBMn5/Pa
WcSz5x9OaDavpRAdYkVqqEoVw9oUiD1ygXBUE18G/h0ZNyN/MpOIe29nxrSPE++U
VuZgrvX/mecirHAfr7fGowCWwvnb/FtAw3t1wslLEb/vA42t6xIfQM7H21OPJZvu
qxS7N6Ttx8zZp2TMIs7xunAWrCfyY8JD13ZniOIF4ztSs9C+uk7LPXNww/26kl09
cPSYMkxu5/5FAFKnJgsJN7S+IZwkvQ/EPmyIHeeMXw3mO8ve2guN2jjaozmPKcm3
ui6yQHfp3ghuJW9cLfyIfVVhIXxq/7a4we3XW3A9kyX5SWjZO78tUG9Rzqn6ifCB
WsBehSChiFgo2wqn4FkJEfEcJ3N7q+fgOiFt9wYfcBYVfPl6QabsBLnxNl44HAsL
ovmDQj6y2S6Ceb5JDuBpUt61F70FnuCw2DqLnRPswN78BwUPuwmlbzlXrtRjT0JN
RR77p5x9RstACbeVFo7FaIU/OdliL1LaPgfnZditK4PFPxkpHWumkqp1Uw9eJ+8X
CEq2ACPz/BY4c3JVayLxTKXGJwXVXpcmh9EcWsSLR5MXTbi4t4ag8k0x6Y9izwh7
/it6YooKhDauiaeRJmNwjUSB8wiI1L17zyqZamgIF0z1InTwiyKB6A4dJWi3EvOa
+yYCVJ4FOsT8wV7tXD0e07OCB8YK5qeY+5fUdW36hw+uO/6faMa3m9emsm3+oXXp
+6AEYChwhbvXwBdvStcXwX0tXEUgZuMb+iv8SAa7tlEsO6krvCXIjSVE7bkSKKZ6
C458QqkLu6PvQH5aCBfrhHYQwGOe3uDdP/zj9aCf+rzlzndW/RFK+G6az8BRF2Em
SppGQhXBS8nDyIF0e9Ne7ztUzZc7nEzy4dC3iK+97fLJkfiC5yXuE5FJUXeEaemz
N3Mqx4DwTNN8HXj0NowiGZh2Rj0VKrq3wIpzt9bHSdMRMMtRK35eqqTaqTHPELfb
YM960N7eEqVbN+GI2RuJJCwhFvlGo/rjkaawi70mA3X+g3hPg9U4PUIQBREbmahh
cjEwOYaWWxh5KFLHawefMiuqPSi/JOPNEZAXpSYzg3Y9pHf0VRegue4wrwZl8XzI
BGvl3u9cazyerRov0ehD1WwGbuPnke8kwJ8yBVK5ihQm7akVuv+COB1DuRTj1ZVv
sPyjmOQI/W4TnxbL6MGc83krkwpUs/LbpDGoxWCEd/eLHRLibUfDrHbWXE3rPK2+
DG3hy6TsdajtoHCzDiAEhRN9RDNsIj9Xcb9fsDYqKeZGDmRFdsAQvnZoi5X90nFl
XCNrmfudSPkaMv3uLXm/xuXMcDL3U6d5Vb39soA1CfyivlKrap2Zv7GDcCtuFQQS
CTq6hmM+nnXvB3BuBToWv6bY5Tb7exhTChOhojxx740JGhOOeOGejUilDIUPRc3A
QmRm2JRjbXH8uvq2YMccPGjdaGvdbJpnfbCfslIzp2PhDXbZCKD6jvCZQsaatt0U
GTH4PuYeHYLa5DD7AEEPQguWvUkeDt/vmDYLl9gIPnxYE7rFDo2CiG7QFp3DiP+4
uk+ScrxLkFCmgPz4sYFyjX/KVPsz15Cqmr8EDr8VWsy2sS5hz3xQec/eEEvRwZIe
g17vfZn4U8g/5qO6s1/usG2beUAkol+KX52ySNeruslXm3DHF/Q7e+nX5q2TLXdh
BEggMW94X8OL3/CSthzwNMFZmNUYB3TAvy+48N8TnjZFHhxd4kZAGe9SxhaUQJ2B
N34tRFXHKggbCFwFpJOMgYRCj9FS1I/PdOB0i1k2sszGEakmwSWjhK8yEKZ2bxur
c0kjh1zbSHGFJ524uxS8E979ZitOiXAo81KAq1Oxs2p3TzbN5ycDNYK0GE6IKz3x
cN8TMPXqh1X9Ase0oeXRblK0maYp0fayG8yBaryL37D1l3Nck2o8Y29tJulDf6wQ
GYsegKJUoWVBP7E7LpKxAmI4O4N8JMEO6CVTyG09EEjm1E7NqeWRnj7po2WWXNua
/T3LbuunceO4OxhBrXTMDwp7ElKlqOeJ8zZ/smGel4wn8nk8N3T4NRRkXM/Sr0aK
YjDGc2sl5RGyxZTgPT+WT0eChYLK3pIqcYr5FZX/IdDEzeMXJUDUs0l+ZTZo1yFo
HMEqnrOYWqr7SPBzD6fZ9GMbHPx5rlU9Jy+0S0u/D1Z4pQiLZDzTJbrNb5Rolcmy
6iwFNfqbhi/U6Zk+5yBl+sKRnlJfBak+RwOlVJE2j4GAkwN+P/8mkr2IznhpZdiq
q49yz7mIc2p9jB1KHWkXSk5C0SXTdhSa9/TPdZgI6mhp9r3GD6CRd8nHQxlG88OJ
hohVyTUjR9XMmoZQOtVvP+/R7ckYg4qMekSUOWTYRLhDX9Gmq6oaF2L/iLkcCVqv
0ArcCr1qZAN0cESNvUPZWWdjJVeSGjDwE8Qsl+ZZ3+MY70vqh6njWwTHNGJrMaAR
ZSSBfOU9RxQ+er42LuNXx6ZjjNFSV9Jy9Ntz710Ak+hGmeYKnE68azCPPST0tKIi
P0BrVtozfYnVrj8z0bD0a1XlydPtUFXMhHIWMEtLmgq+434q11wJ9kEw2AwYzNA+
EgOFxGvj6CFNHYfNjFCvZBJwiDrcLNZ6X0qttqmWRG+TgvTHesuMoxqAYrnygxDY
1n37MpXKU8xOIW0UXJRqK2tR+nir6qbooCOZnDlJnhLbmjcqms6MAPI79NDmqQmS
+z8VsgKXAOCDlPnL2XKxxen2FRl5y0ygCJQ/Jk4Z6O6YzMyfSeabOkXVnJJgN2F3
p3tpSEFMK2BEKAJNnbKPK7GRknufJg6Ee7xoFXC4Iuh2CN53g7NSTus2PC4Ne18u
BtyxAgT09MiyonXRGj0KAPU+J3jq43wnSgBUqcQXc1uWQi2qCM7kx0ZePLppl5xn
+ZzIYyNAapsSBCYNCNsp2kKqGCIuH+qV+hpXUeO2+SvqUx3MwD4KZxhUn225Lk/h
V4ncWWGVr6YFPF44zy2qMbgPBpQ//yEBICxJAQ9gydD6xjCXdR6rYFaBOHI5AoKN
/8FJX7QyQkI/ZBVXq5VqoXkZ2JdUBBGJu7EtBWPwyggyYAY9CpO4ybLxZ6qeGss6
FrTFGglufj/HRH2/rLxShMds9m2897yz2Vs8ia8E/SOWaHEXufJJZRqvujwfVX95
fT9aYYxZyDruqCSJpRVZ17+G9CVDMAgOPdoxjhG003YEpoXKefyYweIbYVNMVn+A
7FQb5vREz/dbRwoHN8cK7gePkzHtGsjDkJ/jgdbIK+ql2TaNG86SJIrUmp3DrJIJ
aVfB/151GKDb+mKSxdfHyf8z02qToMR5Cnsees7IJaWnN8vurTX9TudrcGSik71o
8+rh94yKJwUFl66tFkVHyh0aQgNJN/YVcA1S/mewc84yVuZl5Th1vZk8897lxpvU
d0MweH92wcGUzVGXTcI8Ob00DrvLaMbf8WfQ34njU7ZefKnrcYfMr5djIJMxYWgO
HdUYSXrWu1yLhdHbSIPotkxwHlE+MyE7fnBu9YiBcnFQXH24O6tUq0usxA9Nn+UD
RLAQ9WNSZQkgUpezSKRQkZv22DZaLtDvM7bDWT2zfFxdXD0m4ZlEfYggFEzXS25/
tDmYJp4YX0zH7s/n4OqFiCra7L0iWVeA9qdNBRw4nkoON1dR8oTJwBCl06sOaCi/
Z+7wP/EgYVraKm8dDfvfNy1GKil228ckjLGKf6JhZ1hnViV8M1P5u9hQfSqCG5Oh
/D/v6d4z1ih0JDY9tV1E8SrUaiYvAQcrlwiSqkzpoDfApHllxi524hnlQrPOUiQw
xD0OdFYgaxgQyfY1NUOoXCLfGzvfDxJ++3hKNNNi0gmqpAsgQ+nSgRmu+0+wjnnC
UzRhDLfe+m36dBYo+oQiafZ68Q6VZd2+SeAKENkVXCrEXNBrMmuFcowEX1WJ5YGg
E1rCycaSzfk7tDVcYL5NcwMkL/ULkLnxK+x5P5qwMQPGpDih4xY14hW4IFnPbbYp
y/x5hFu1YKCltyDttnDk/zFASVcBKUj+c+aDLMangx0UBj1g9yaYqEp5kcD5/Q+4
ZhOR+Q/xX2RfmsCAUHrNKQdaFHH4Mdhi4jH36D8oeZUVa4/9Gs3w26Z0DmRTuoOe
4V2xdfJZZe3p4iszq4ExxwjfyilSboA5w5uc3whN3YU8BfKANsGgC0bwLtV6+O0I
MKi8VsGUwjK5XDm4x380X23Ts6OrDWQ5LWTUSKkFrwjdkSDdqoWtmpDiyI1GmayA
ZQR49F3j54xyBWSetSdB+tk5kbDD+WKc/vRSw8zaYsqeTUNWMT9NL4SvzIJmOZ8A
neuw1dOctSXFJ8bXaoxFkconhk9G3wBZZy43ibfxkGypgjRDPHdm9A2gwzlr/AzS
6XRuo1GYb3yr+ifyk2XqewhWu6Sm+5mC/dGgZN/GNip5d9rJkHVTugDYGYnUvogX
cqk2qx0hUDotKgL4r910oNTboMuoy4wqcUeacmdlIeVCHEreSSUYe87vslz6txo4
CYm99A6M+lJlLW8K3tQyP+xWs1w2NBZEalfOAPBxDlRvNwwglgLEr9HJslyt1GQ4
hS9xbuNLeO4ynfMzGvmixUsdX7aCQn5fcYbQRPIYYPaMR/8WqL2oD2aXDKSbWxXa
rCnbcH6suTk7ABje1N8fF9tRY4MPueU67SYWz1pQgEFIqwvmhipKncjUjZcdQsgQ
UWsl7NBZul+OgUMruSBGoDmJsH4qFvEsMo5GZehCzJtPPSshXSbOAnR+ZhPUPQcz
MT3TfGgSC8+q0TPjibtMY6mh1MuK3VJlqEZKF2fq7kAI083V+ij6CGKJto9fT0hc
ja8IkSgI/Tfv6/iHsXYW/0h9rSd3rzNN1ySGeASSPqA=
`protect END_PROTECTED
