`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oGgqEH7bEbuXZVlPUDmMq0XZK37lCoB7Al/cVwTVnoZUcYrQ8B8oRvJRGhEd2y84
iLaSVdHOynhFFYPh2LzEWoRmueopDMboBJJucsYOTWimhNg0tUgeon+WGUjS21kD
O2nRI2qVmx4i4InecLhYMB1OFADusi4KwZfmoyFoj7Hv3P/pWZ+sOLhGXPqVRtpz
zR2K4Cf/yHtboyAZrwDUE3kJzxpfMeLVHni2eLI3MV9G1upwgL2xXVChUZlaN6Zm
V7YPi0IxaOBfIzQ5bxvyfzKhAGOSk2LbpoXQsI6c0Mqi3R3aSUeUu3aiTvgPZ5Ex
YcGTph8CEmgUB9mSnhv6SmyUSzTkMnNABVXvrnkgFVKpJArSg8cAqlOlliZU+NNc
8xtu1yQAz6fxg1IslhoapLqRCYHjCQiJF6texrc/zFfKt7PisNpTDXa6otweL+CQ
vt3cEzoQfkcjJM5ligkhUujCFikUhqDOrsnqsfDQZlYixyaQ6+JeC6q3XDHv5XId
kUhQAeejUyEo4DXBUWGrPXUvujf9KIWa4n2hI1Cxj37PQYud6srO6a3MWOTIRT1Z
dgHHn4jVrlCk6ZeRalSm2snsBzcmbdbLS7L+0DzBaXBGoqVnDgQ6MiuKyS9K4d3f
tas0V5c2y1i3qwLk0ABd3sdRQd/swBqSTMS2VfRwQa5Yxnwu1fcXMNA0pTAb0OaO
CGf6nUOIY/MBpKf8D63rzA==
`protect END_PROTECTED
