`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RCzOUMsL0ybzRh7IBhUJSaTReawWE5TpdlTcZaNy6N47yxoXgaYAE2KViJsxubqX
2if/6kqMCXawMMCboNONMiYU94D12L7ZO0h+IPj3ntQ6GMMNUXaJLnPXclBhQjL8
NrOx0elcxdqsmJYAsfD5A63V9sy8JTj/4bJLXYqJJm8gHZ+C2tNuP8VEtAjqwczK
F4Su+xqdixQuv+BOCqnnY0IgtLyZWY2LzjFBLGCS95RfI/oT5+lCsHRZDbo+Kl9X
6x2kitTIwTO5PURdj0Ho2CTUGjUSE0gYYpd4ETVofx3joAGO/ZhbRVu2Qi6d3win
ZjMzDEyYIcYYtWUcq/ZW4UvZmgDOkRV71jBHa2mWQw/8/GR7WU1qtmyOLiGsw+yr
dfEoUapjdAHTae4Qx76NDVOM9pEGNG6bKNxyfJuuvOdnxLsE7U2CcWYilKvNFA/l
/tlREswPys4D7NkeRdfuBd5FAG9fsS8IVVVE7lU/T+ITHguJSYjsczqA4ufVG2ga
cMnK/d5SS7Ky55QDLG/eRfLiuaDPA2ENlazArtNnZzXOqsxL1rwWhCNqhTScA0ho
NwBXH0Q/Mq1mIRgxY6v8qaCjWALR9A4vu3z8JO8UOViSptOT/MKK6hofWpB7/SmF
7Iv+McMm16i+vo/zqCmsk2o+jvw7bVr5FLQZ9s/XO0rc4Rg7pG0VFW8Ua4T7hLtX
8iuXX85hO6uBhvw62AmzdeZP6iGSZ6rXGbt4hUWOmY5jvK8r4u3nGvo+19W65GYp
`protect END_PROTECTED
