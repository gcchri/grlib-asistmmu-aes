`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pBc77WYDAX6CFo087mqs9k55SVB/mStOrc2fo5xi9sBge+XvYTbtlPeIn3ofyzeV
EW51SoipMcJRHAGw/9yC87wZ37/bINFQsJ1mmPMFg4B3vt1K4zyKULkDwNkSz3MT
q6Q5Kn2ZWwjVcgP5b5hoRinjRmGjUnYQ3Gdlf1PMePmnhLoyUgsIqCTzUnDglWsO
yxKp/BC7eheAQjqnX6PLKCB2eA889X6747mAE0L/iObvsA6J/FYw/2/n0qgtvXoV
JeKDLiJvzfjcu4l6SBkXc5yWpbfTO4XDwtd4CmxZfpMfoFVpbdFzh17aaT6PaM06
mAnxQchkhXcvS7PdySFNF2N2r0W28epRhJhae6oDa6BrgO+Ao5P9rNlMpM2Zit9R
AYypuEBeohhJ0ApqyKgtDrsbumNiiulTPE/HE0xDb4tKM0RvMzrpbrLSZtMm9ZoC
0uZRPCeARxwk6dMbnVDkj+K7F/5gRJc4nMo9Nd2Q13//+NnZCdtlc7u6CQLdOevc
RJiW8pzff9C36ckTuYeXmp+x8m3ivs8wV22+aGxHpPekmlC1M0i6oaNpUAvWJkEz
PZXGE2i3IdpM/9rrLrpj7lZFp4W5DdDYMRPGuTK37myAufkZvN9kdRrZuo2H1pPt
n7p4L0qQx4UOZxRNHoE+F/3hwXTe1yjK8eBq2/2nlfueF/xUhjYXw9kaD8KAXD/F
kNPdQV7YJy02K6GjliV6H8O9swq3ovz4kFGze+lR/N8zpra0ojvNJIU+U7lzf13p
xKf2aVonjNWFFC2kUoUp0wsfwAM+rDrZKg7N3TmB7DQLK/zVvaPqg/gwxbv5Ohlp
uI0ECLldPmqx4NAepopBzkQmDrM9wHWS019dMvkNV7Eq65Y5oZGHx8qzppT7m1ym
D7FEsMDaCqW+M5O/il3id9rJbeG/ypY0rySuENZ8vzs/wOQIR7K7EiPUe/s3VVnR
TKVsVH7aPiL7ARdJLviwPWw2mZrJobUBgJVI4zoyBzD/qNgmFYDCBkx1lHkezNLg
ZUvXc7p/ZXg3mRnyaYpSfpMLcxCDckQvuEhAYGoYc5baByj5VUY0gZlXDageV1wn
mswkiCi7h4k19rFQPJUWv71MDoM3ihek3mjg/H+F82gsrqH1wWErsU1qyyUcDCyV
j24qYQ0TtqXyc5PfzBDcz6HVGo69pPrRMk4E099YhpAlNIbkCtkbIqpPwvqX2aW4
qEhKM595KmRksGEJVQIQmQAN3h7RlLiQuxu8G3p06wJFiMKQ7CCupBaaCndunE82
SinbN7CP28ipwmv47p1G7FjcBNM3LQoWqtzsrGCZKqBXKHPeVkF8M4QiRAQfkqBp
E8uEcU6G+uV9jkdbtfEnMCzEUs7VelKJXeiFSOTo3m5EI1j6gBYVPKoqRF+zaO8A
oWkoAu2IWWgsfGzVFFsuCetp/ZAUiT9hl5svWhQt+aaP2+iiPv58Z1/XXTFbVT8l
MnEFpwSDugjt+ew+dwg7BAKd5jA1yWpOo1eVLvfBN115I5I8xpGirkLDcVIo2vT3
q9/FYvLkiBvviIeVIZtpN6EyXB6WNmUt+PlusXdIvbNMUJWQ55QnTDfRLG2Kpcre
oo/a7LGswt644sj5ZkbKukRW6Wc9QlZGwmmBcppLafgDZ3BaY2uqTFqDoIHqtHsu
CnHVK83qC6PO8F82oK+2UMIR92zTIN+VawCOaaR9DnLA507Cfw5qpeJ9cJ0bS77/
31EAi8bdSnZ7+9LjU25qEjTTI1ajVLBESy9WJjcWBf3Lwq05uCAo+wWi+hjr4TGy
OUgzxATmJvQ0hMWB4qOe5ds1W2QSL4XUtudd/igRSNfUM+Qrp2VFoKhx3eM1HjjF
JBTGbzbMKGoR2WmYw4hxu5orsLgpGp0bRucF3AbbQdYJ7eASHwPK5fptSs7BjW32
B38YgoMwkHiSdsJJjvljidPbwt8M52M7EWcJ6N7HjTwVeHfA1Dpo2tEG30CgXeCM
UIs6dZkVloTDH5LlWeOFdIqqlAB/rsD+imahgKTr1SIq084guXHay8IPTavG/kDy
kxhfJQwt4Il5r0I1SsTdzHYzLlqaU+GB7Let5KstYIx3sus/Qmgz7H6SnklPY9Vx
bE3uLwXnIz92FxcD8VuEVDpOnEHjR7kwrJyNT4w1YARCy3ngfJiD8vAsRhdfGI+3
44tWMQzlTMUXA6/zxP3AUxPL9QB2ECmxSdo8pjBXvfog+DdmoulHQxpDkDuQIdYl
GJgRgMYFKb8y4Ywb0sPnDbCdS4+11O/XEKtKqoOqp3vW44jO54uRiojnd4CcFDk1
NStGknuL7zkKiHpPRVhlkZSAjR6iGmSGE+UNTYW6pntrl/6VeEhtatB5vJZbCLIE
hXsfpQVvKWgsQ9enHXWsPAeSO0fZtp20R6AjBWUc8RcUExIkslv0uYM+jNH3ZWKo
ZyZ+zdHSU6OzJII92rfnnaX1tAFuDcoMLPjkoorcM9Shk+0eKrJyPKD/0phNYhU6
wvzAjw8A+h/d/kNdZKrTVVvDWw6NnqkT9vwnHLlqv3Oh5zC2IDoBYNG2cw052onE
zNrhPhgk5ZfrljCXSqV1DKSpe6F8TtZf3jMJ8cBhlAIALMvrHCrwlUBLkZxkE7+v
8bLSAZQoRl8hJplEzSV5KEl6o5DYb9gYPHuqoHPBTGIBTt9RCE5R4E2c4B1WoaAb
KGm5Jd+4Gv0gFDrcvMkl0EE6Bzq8oYWBr+EE8AkOOIZvKPjBjCcU8ew0OGiEqW9d
ua2Yv9p9f8+R+GUgelyW+kcX9CrU/Y6SdQqis0fyr2SLwhwhsozzV5spI3jL6tVM
+VlhlGSHZxYVIFHdAtDYWbkBnA6AJg1MCM/IlbAqC4uZIlSVFtrQOOLtzoFvpNil
tbLj9xXhsD6ujMV6+Zb3h/NcdDSHsYIG7N2lttUVLkkA5up1/tMIu13HjTD1rsic
TnEB6vcgJXyiI8n13ysRwM8le4EJ37JCFxFPYz3sLdOePGO3yqan+1ayMxXC6kW1
Ka7Yn22YsS55U9J7vfEQnCnaUkvOz02LsJkTa8maCeqNLIF2uXc+Mdo2NcHi5iix
3tG/l04lSwGGaQVSdxdpfgamizpNpgWFhjkxINxq7OmHOaAx9/BMpVLdmpC9AjsL
X7zD+j2CIRoVP2OVBmaYSR+0jll1IfhVW+yIjU+oRZa5nvWikKGhqT96vUU+sQqW
tQRyL4RCw7BBhMCP6zLpndw2zy02yvmsq9CexB0PJCx171brThnsRDSqmO5Mz75o
C+GkCtmO3iC7MMD035kCvSbxvNHbF3uxYh97mdfA7RWIbueLt3r0Fc1lpCWaKTzP
3LNQt1FLDr4zdb854yVBrIZUI4qV8cKJjawEEuLf0ZSjkf6VEdLENy6aTL52D2df
chjGz28tYjvhp6Fj8wulgJiSm1gjKLBotNyhKeWmPNiyrqBQpGbZVTaipnKj9PT4
Kzo9sCEKiEtffaJGvlXZ/bZQ73OhRU1/HM3lmdl9vagyvcYNTlYADg4CYAsdQJOa
kXWzycYiqnLrlfMNdzAUGyQMsZ0f0rp2PO2V0DqYadsTsEKh8oERS5JMoq2mZUYQ
gudCt+BqUkiXHy4rNmmRIUt4kiJNKO0Yg4/yS6bXUlYDhu1TCnPg9Yx6OHi4b8XS
C/PYcFfJHn3gjwzozJm4SP09e0YYLOvKn70eCKLhty1Bf/Fc5sASD5SRhepqMR1G
jjQUj95AkkIdEbCjv6cHDMU0MnyXMKYTPScFLgagew0hLPTESofnxRHKbxrLJmNg
uTt4oJLd7b7WqM21tLQKoh+1jsyMOd7yJNsKauMudk0+EW4vddJ/m3HTaP32TosS
VMBDDKSx7qSPm2LSAIme1p+Xp8A5sk9ZeoJJBQwal5OYsjpCvWa6HVCFsDxm9UJT
wh39yQSOKnbk6859X18O8C+CJCZd0mvoxbCH6GPbJ0EUAm+FMmRI6yCCPlxPbNWJ
Ng4/JN/tJtfixyC9HLbGLkRfXpMS1QijFvW1y6IURNeA+jOtxivD3Awnc/m5J2te
Kv3M5mrukHbtoaXjGt6/vTMfZHSEFz/BwlnYg1Zl3znRDuIQm+Glk0iNm667501/
QnHySBbG0c4hYy+HWZVY7Kb33wc0fx2caR/Lg+nq/zAj5cAXjItO50ydi1UEUEYI
ImgAv8jd9EWfU8fFawyRWeqgEkngHSrBrGoWZ13I5wF86EHmZoyKVvUcLMVgI01G
TRUy8xh05jIgXLGiAP4U8B/5y6pXYc3MbbaNfj5ru34Nrwj1pmJH3kdBKr+rysq/
ylfOdzyb07T9MON89tc+R3uffQwQGRQQWHR1kIOxAOm1wkD6nYvR43NunGbMC+Id
2JWsmsSpAx1Nm1MLrlUqmCyX5IwhdCmnSZE8doVL8NtlGRk2HSqlAzdIj9V8W93q
4uxhEi1NmUjpcXAzX5Y++BGUIrIKzhakTwj6vxzmmO7Q1VFMyEfAjFC61KwIu4vo
nBLV8rtraQeyl6iIfkRX6Y909hVey2vAPZYwZv9wW1z6J+Le5DZlAtwWDzhtGmsR
r2dr3B12UQlNe1PclAAuQxotSkM2uTWiUq09c8W4C2CScZ2dwEXWhIlus5opd73r
2BGbY4cNZyIoZs7KHRtddEcZInCk/LkiWUWYLXn91Y1tce3+Rvg2D5XgDqHcm56P
4R5qETGEkp50qFIeaOSnsTTZO00MN7agO3FZu4AEWLP7B8KLEWQJSUjQtnVGNdAs
b1jkefuZcb43XaYIV32IVH5dqwvgE2xuVRQK9JfuBMayOtMWvs8pGbEYapvMQVBL
HXl2n/a/895tvgCdfxzx1ZsaEYolFEPHzcHZGO8r2xhxDvPDLwMIBW6djPrWXbzB
HSC4U39OH0A+hL9dVdePnIoR354Af2lltx/hGFIOWUzNkus0n7c1oCWLZ+TEGIYo
EN/UD5J1go02cZmWnoyiKA1K0FwYrwvKb+9KN7PlvAGdM43ExI7TZTS9W9ZHbQtF
onGMuI4Z2Z7LgaSPYqjT7jJMn7854oVDoTK8UwzpcpJ81b8gbUo2K90xgxRi4LYm
pvzm6N289HDbUmUs/DmnbY637ZjLbl6MMDhhrQIbuCmBnPSnpBI9GPoTK6Q3tN+O
q/tJVamJi86nczpcx2cTP+OvgBhor/ZiC77IxsYcBOWxh8oL61vX2b001gCAtdbO
PHjH2oKbqsZjEXFdMyRVJ3VGmIORA5LuV16lJrNHnpsSzhqi6nCaO9+hse67df5V
01C5ba4fzPEyOT+/fAZjOfR/sJ8IcgD2ARANy1okdmSsBCMxFrl8B3FMmk0Hdgoe
O7ASNqOoPELkHzIdTdge5Y5blTb2qqhipu6U4aqaT2rzIH8RPYiIZ8Hc10fUssLB
e/l6Xp2s49Ij0pRR9eMLoHl2eLvR6c1ba11cF6OF5c0bl01UlJ9UUhdMlqzUHgC6
KTmgmCvDO/ZDyqGlBrh1BlUBpDhPsVV6t96yW5hOnU1UvNgqCHvtubVax/UFDeLz
qP6A5buGpP8I/Ghd5wF69mdlVTChyxkpW1mr0gPAKSHLwTSz/l2Ez0dPUuhim+me
4CYcjVQa3ssi0WIACVZQSM2M20uCHu+47kvgrmm/nEiYP8g1aYiw2vvNPGsfuuoo
q0LSxRwBg/NGxLaGQDxZCgcZjvTxLR7hNMDmU4BPgIXURLc8KuKnkQOrJhxoERZh
+9yMpVc+heyJgLnfsFlRsPgVqXmpB40EC6aJ2klMXSO4SOlMf4yH7nH4EUXmG5ij
ZY0FPhn2PAaZw6Qj/QFS7rGIqJn4yzwKM163x1wuLmEQuJTzDUO97iididDwgtNL
myRmG3HQwCubnbG6uhBLY0nZ2hOWkLz/4g+9BlEGiqxQ7MnEJl4U//K74UShifDM
NIOM9aTl68ZghjztzqIvTA9GNBUlkImD3sYpifxTmExj86U9SvMEk84J1UnRy0HC
kFrNabsohzpQqgSIQvWS4tiJQBxMwB5aH94omS3vwdu5OUtTEx2izLhGIOUybvgh
adTp5O784+qBdHW+gjSF34UgbLtv9/0bWQnprqSoTSuvOL8/lZLzFIL/spIhEPbs
WaKiP2OgvfwU4T6JOWJJ0PdM1MykxeGhXkcLqNUxGCgYJfLKkAyL2ueq+yJxqKJK
IsMB8rVhItfgfcCN+D/NGA==
`protect END_PROTECTED
