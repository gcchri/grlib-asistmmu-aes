`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c3tn6UAnwu0S8yrh/hutgF20HGjQRKP7thmyoDulBsT7n8+6r8vB5k6BB3aENWcz
xB61MXLztrWXxEicQuMVjsuc0zt+YD9VQwYEAhcxhid1WLLJCyC9y7GNAqPa+Wkl
H4GDtgqsPJK0OO2B2bCE/ZWh4hBNI+xKo6t8O2tAoKMgGPvE33f62dx/XwQy+WgQ
m/KQGeyEFBYw6g4e2TcTJ2Zj8ksGmxIX4MkBb3JuNpMY0+snhl139FwVfU8FYlw6
qg7hE2sXk4dcco0l3lZqyKcEFVCmMG878/A9dRmYXPelEthuYIwJ7vg06AaHCusd
4z67I4E8W9HrdZdCzXfdat91JlSJ45EzrRBR7yNzQ7xFCfYpT2ZYGfory8iy9UKr
nYTn21uVwV4Vj8fQYuzrMS1845FrwtTWC6WSrfWUOWdhwdjyofTUt5XQUhfRCCZF
sHkxW1kj+DDWkvjyTog/TZAEfCcobMCzPS8hoXVQLTDFcU6IRtECPSZ54cFtap4J
S5ZXC+uO/mXOrZbWXEW0bI65R30rsbKI53sp59KEc4kFbg8Kzp1Fbdh7t53GQQir
DXncetCIvf6Y1flDmMxyvCnuxIDShqFZPk9CW1lWzqu3ruKl8OeZw9ii2cRqeFEm
P7T55OwyPi2JgB7h8rAH1eGhbNg1xrOH34wh1kofIHxDNHll8lqsI5sfkSC6fbdq
bHWANICS4loVD8TaKb92K+xb5p4tP8olRwx5i2E2suRQnzECytPuy4B0zWTh1Sq1
CIV/SMp8Q/e026aXxqM4BeNA0DqwQQb9HvoqcNBtxOR706XgH//YnJyxWsJSENqC
rtyTBX7eHRBXCusEkGQ1TDk8z9I4JmNZ2rRpYIx5PNXd1QpHdMyNFHkE0mjUC03T
uX1vIlgibDIOTqu0K4Jr3JqnNoJmO6e2SLGJqLXPMgVXMZvmkmJPaswSg01vVeTW
7Hgr+/R+DhDQr2jlFCb1yudknsX6o3FtlFiesfE8R/G5KNNk8d8tYiwnPSVI8hLO
TNbtzWRdbjZTzHvTBHm7+YiUPCJ7YgBQ0AhEw0W+WDsx4e/Z6zY33WrFGCm0ilr8
ByMtOI8MOyhvU3QzDnZqBA==
`protect END_PROTECTED
