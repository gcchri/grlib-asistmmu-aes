`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uOrp6kes01O6oZ0NaXX2DuMHzV8HFKZQIxK/pIxMgwX5D+nfvKamVBSSRR7YDfVu
OA7QCjv4mlEasgxdcRfLyt2rT/1DXBBkn1ciWxzUnB/DN4p52roEBVlyWvVXqj7M
p+6VuQv3KCu1sdjLl+Su83TzhKxfLFyDs0Q4VVV95rLRxIYnIJup7S3VOtKrmnku
qJ5+quDWVsqNBoYpfRfe9iMfu2w5hEUbeB0/ofhaMqfa9sF/IS8yKztVxeA2scEi
H8dMF02DmwKVfx2EV7PReIQ1Ep7jfN+x3py2MSyCC6hz8VqWje/pbePf8knvdV8M
wFj/io9drjb+oLbknSUOUVAJdpSQe7SCyL2gtTaRif1q7NyXMMPDIWWTmlHaFOlw
l3GK4C50f6WTLB0HAoSuN1UAZQUrmqUC7YF5Xjpwwf/hNPG0qTVUvq9YIt08fiC1
/YyWcCeg5ozgADe5sMaRa0rPk1dnGHQQrqqSWklCqe3hlT1xY/oyB7Ay/kMdYhY3
jOOSLv1AT/fayCqOZk+Q8UBvUs/IilGF968wba7F8rXKaA0b5ZpEnBskUiEhqapz
xiR4+6tyzyRRyxhGNQmvcuBIeKSDfol121CvPplkBCVVxy+F2h7jeLKFN3KBKKUz
ui49IO3Q3nh7nodocZadsGEkCgBGnPREITFyfo5SCla4Zg18KQd/KqIAEMop6m/+
saurxtmqm0+bhq5NNo2w5jhNsxZ6MlS7M7efa9h72yd+3nT4tHUN3Cp9MISR6R+u
hOeEIMJwD4vN49zRZzYepJoJugAInEltY6ez2eYVVJWvhQX76f6RAjnE/3wMPTNq
l+Tu7lY5nuZWG8e4wUg9Ok0RTxsoubG0q8jz7FbgtBYt9kdrNp8GLHdcQ+qWSDvV
JAwFV7q7DsGhA01Y8j6odLeQev/klHwzcUZ9/kWMZaAUzhGgoMavPeTsZRMcwoO6
K1tvP9C5e/5iwCDjPuvTYkEXjKt9fhZD7sNhaE0v3XMZA4/qy7yzLY/Oged7TLHx
Ok5QnDFTfWPFH9W8U1eqtLwXSaqMX3p/rtVqlbU6lKVNrihNdXGH9yaZJ6joeqfY
M1iVzms1NwjLrIeYTNWWfOPBYVtsfenyL2uh4ixyfETcAf/PQpd+Ek8U92mKtphP
1BUyDcz25Cj3HJvaLENITiCPnwhGUyC7kcmGiZu2v3rih/W3DiwZ+ODh/SVOZioH
q8VhzmS9ad1dGtG/Y/xlhWU+HdpTNBzwb0ibyDJKDRVTlP/5q727Y4KAygoCZ9VN
r9BSwksS3iEc4QrLU5LBPCDJSbqMFBah/RKrcifDOjjarFYeLH+7zbRQEZa/BkAe
7DNIvQd4cLN4OQZBjkuLQzN9slgn94g8Ps3Yxm6nLO7iuvcXynBMnGruwmGgE149
a3rIE0zCIcg6gphVFCmy7aX+VoYwvnRfXwznxWsI92oyXNN28tEa1YgSfor9BOmj
CA2vTEzkLtXVTi50BRdajPMy+TZy7PZ6CmMRbHzDQRTnuqsHJ0gIW7LTp0Zk/dJW
ZKXel5TKrSv2xUTHfi8R/VDL5aGVjAm4vaPHG99J6/N7sashL5pzv+KdOzBY9Pp8
avM/9cv7KMfLFtQE+dMCwA8nQ+AzJJd0khBBCTGL0nEb8lIpHuQuyf1X7UAQa5h2
CcIIifB74O6TWmmBuDmG+/wrDltsTfRuFxhVZ2d9UrJH86rQJVkerFnvPZhG6wR3
gZBMyq7fQsG6QTXoCYAtmR0wwWZeW+I83GmdndqR5SSC+Xh743hbhoy3TaBP1wo9
mF988BfCYo9S12iduvS5ho7IIOOb0Nw6IWK8N1FNahiuavJzt907X3O04B2cuooZ
esfyZVozQYSPI3oKc/Yc3oPEL/4pzl4uTOzcLHGlZoAJpUZohuCF8GAApKRnU4GS
oaR1eYHLe37mTB2hw55/qFi1TFWr0WLHE604ItnUsk1YUCzK46rx0MfwodEwdwFP
7/RO6GL8OxoC7itZ/x0inVd+JLTs14qUgoURLA/fK3xnGhQbw73IwPNw3thdaYFo
rs4vyY+522f18Js1EM8kXjlt9Xpgk06hp/H0d+esw0s3rN3VD/oiuraw4kOWOS/d
QsqKYnjDrRjnaM+3hcAqC8ZksOobVZdHUYOARmshOAPLk+edzVby7cYkbCp2GsWs
CykwB7Nuh5JJ8zA1NWkc+LdDHBGcE0KXAKsNII+CtS28pGcNbKc6alJ5Gt9qGkY7
uKwpeuq43FXYQVfgtlBLYi9jn6I0BWppBKHYyBG4IxqM2TF01hs7vdqf7odvVdnK
F94dxalGQcwemrKjEn4WexPFVbD6Opi2IIePXSnjLhszwdb2sgtxZJYW7rgZN6qf
0vBuJbf+gal9W9vCFmbBW0+c0Fg10OnbMJgBcRMhtzPZJQU0UMfUjUaSmTxW8mYy
irxU2BJRMi0nQ4zV7c2U3ibCnfff1FQ04mXFaizqJ39+U7hGaYi8f0V/3t8occz4
ps6LPCGDKzjiVwx09i0M1STzZT6OYB4u1Ae8pRRyTdPoIDcldrP/+sRvqMKFLsw8
V89bO6DjDyfh3u8tWEUtc8koPnH6JYyN2g2mDr1ppkQ7NHRCoMY0G0sp9oR5E3AE
r3vUeIxMX+Ag/vv5TEDeMgYv5CFeEoEmGxpYqtDl7jeHqCN5KUVJSEBvao9jxzto
M3EtJr515oOvK6B2QdYyRaikK9THY/2E3j+8U39EonkhVQU7kR4Ok4hNgwE71wqZ
cLkg4PZG/Hfxt9jl0t10Qog+JYN9/SYdluqi9qbHEr7Gs5KDGKXNmDrfAFq+At5o
dHeXuwq7U6vr/nsktd5rdPuYPW4ST99FsNC6JgJaz9+JjDcNw3RC5TwW3poL4Y//
FAHVXnPk0UnFslPhJpCMSIR66rH8K2q0xvnTADSBZQgmGSSCl49ZdYgJ3CdI06vd
DXeRZqCidca3pgKU26iDMGEbGqqzvqku8U2H8VcIgXGR+VqFarWWwe7606MJ9Txo
eniRd/y0A9gERxBmjtZQQYn3flgh7EkQT3Jm1sElpOX/e2HM+lWX9j/9cGeAEgWp
QvxhPInFFVCnq6a/5ReIcHl55Su9mU3XHYAgao8tVX1PoPCHvmA9iyV3KZ66omD3
t9Rn76efp06TtypDiM5pxSCkpc4wxbFHSZvItQnKQVnsVvzNGnnRWwp0cEX+kfIZ
7qVN9npE3nOm15FglE6X80a7ZWrebrhWC1Rq7U7Q3gIEo3OUk/s388pADkjVJJ1g
S37BSdhmA8Y0VwoX7FRhxEkLJzw6su+dYsnCTq0+7mMq1OafzOA+185lpY9JXXL5
ORuLiCuBeSxuBYpN2udIIFxsEz1d0UYMYLgfjKtzrJZSECI0BN+Q19FJZecRAaRS
DY8Syn62w4UN/5LIklEpYvwk8js8R8QZR764L2bExVpc9f9nJJE1LWmdxR+6yXKE
bMmmBlhCb1DU9FPnc7QJkPGUY5SJR/rRswzuw5iBfPkp4JqkG1K+XhFjgcoCkz1T
pkbVl5ZBHt296aKiR1TFlrG8JLnsoP96paQBfwGB0RfOVF+BpdkMKyVIDw/Tsice
uW9IqciATHyPY0Own22wEFBxzetOZwYsyRkPXZHTK0SZ8WinODqIaChIoWTrAE96
1xWZgyFEkCam2j9sSg97o6gHHlvhD6RRi6W/oB92JmHvPhSvQOMDMPFE1LnkS4gK
4clEkflqUm4lAg9ExwUud09DobTTNbceCK9co/iiQORkMBKxLy4ciBDSc2u//rF3
eHr+6iLy/B3EC+mB25+1iTCpSMpzJIooOCyMHsR+azoGvSlpxqhTQ/twYI3w5eds
XPkKJfwzbzB0Z6iNTtaoDDLTRii4DoqkZLR9w/lqQV3+bm8Ba/VLARn5vJyzlRRQ
IIX3mWUJToD19dgjdJUbaGjbuwUTebDQFBnJfhoFwqyTlVxdQ6S8Lr/gBH9iNd+h
vHnwskp+D6GI9+SswQvQ96a+w305qCTdwhuf7QIADQ+Qvz96/OXxqdTg/3FgqEgh
PoS2ZZFVoyIuV31tUxlWJs2FSm149GniURbqkXDryLiKFMw1Anp7gapYCoru8dMH
7cG3FkXkfMeFgmuL+LLZFyxohNrijfo7aXEGI2Ll+0lUeufIAyRN9cFvvgj7Syru
DXF41li9SvFtQN4Qkb45WejP/7lRpQ3Bf+kHyvl7tuiIBLJdRbvGNQuHEB3NmEhd
gy51iJ8C22qQg90JVYQXGsyXFqS296Y+IIIGVRkbE5p/mRFBVRSKYR58CkKoj81b
bXkKMVrKW6afkLVK7CS/FwxI5+KLAR8swj5hCqOkr3TG66fSfFxwZ6KaSarYp3re
DIcpBFAlnaxhcXx6jCxCuWIOEsxmqiYresUSrP/iTy7of+8FUEeV/xhW+4i5/a3y
EYNCggyUaUpdPfwcQ+W7Q6XP6pZVVVcTFhVnUnXLkZOq4HW1GypM7kxEu1SHtCpC
BQf3LlxQoiSdGC4dfalwHyXlkFQVsH3B2NoceyGInlr16o+MToJF7oBm2aeT0mK9
D62KRLm1uRhAanrOWMrKrmb3kouweowwmqWzz4pYx7qsJtjQkGWeYHW5WjazaRZV
VM7gknL8bGcL1wfQlmz+gC48boNjiugDjz/Q9IyHj36US5c6Ilu3wYDcgl+WU15I
8iDSEcOIG/1KwvqoP+Pr3JwdX5azL1UWPuR3tBJWtLfmOWX6z+ts2RLSRFk0g1Zs
Wwpi1B2ZqiLz4ELMROua7nhMrAa2/CyurkPEqZp5rVXwYdQZe/dU0LGJ2LNbSuDp
CdTJkFYZScV9OvTAGbDRxFz7Pq6YnFp8PICGUY/pc60/Je/oUPSRb2Sk/OIXyzbs
W1S7ImcWdmUMxUTTrhaVmCKlBy+6vUKoZ3/LVOAceFhK/Bj56+Kk2hLWypaaE2sY
3NzJ+iFtf4EOo8Icbs4eiJnh47FIwnZmOmtPabhlXhFVkxTwbPkvz2e018EdLe5a
GDeh+XVdiN277Kp7u3uL/vQZ0Ues0y6Bj1WQtNrVzXQTt9H3MCTT5Ij/CHWmE8ol
8l6BRZqhJ8+lOUWloqAd2DqfnLU4vpAjkHOug175uT3phppBU0bx7h+Bri+DcxQQ
34yaf+vBXtUypM3dsGulxOvjvyXApAwyqPWuRA4CzocC93pfuBmq8pAIl0RzTAB4
oULncmATg8O0s9i5Mp6rwNl2Y9+gnT23VKbrqHgfHhiMtQGJEOLfp9xliCJ2mC29
1y7gTtgoxreTBgK9NqjiUvcJMrUIkj8ieJoaUn695u8eJ1UPcWr+EH5LVjsBDqQW
1VCU+aw/AkKMi1qsxuOVrKHKg/5LbxmszOxSTL5TEasHjTAMIifMt1jCHkBeSohQ
oaotRkeq17pUMdTeIuc9LINwy81iEorZ25kCam35EIEQfAUjLlvSFBjQGzeosCrJ
nKYLXti806cecKX/4VkQMb90AjoNVocblUUdC0Asgyf9ZWwTpitf/uDjLgejEJ/C
6Ep7dKV0RTQXBAHUdJVo78vj/c34J2jdhBFtOhPyZvbBwq8/7pefH2GKTpXtVBDp
odokRrL2Zr+EqHpvnop5ZahFTAl4AaZjro26A9HQYfT5vQAguEc80RUOprHjK3Sy
n+erDiXst9xPolkFlTtffelOElF5Oqck5cdklkQGWBvmAzM0abB+dV6qwigDqiBL
/uefU6AKgGWuH1ocabOSa2+ydnLLKCi33QtQG8YVE5V/uAGN/7TVKn3GsdyZUu6U
rq6H5fFgprX06WpGVaHaqwOFhVczc1WTASabODZzrWQcFmP4dHZZMkKKjlPndvrp
PAUyLPRiwzb6PbUyydeXiBjmzCYRsKRfDrcBXRXnH/CN3xh2DD6aOCB4WNBQR0EF
f1nQuPPXOqnoNZ/VmJd3gMRE/1rOkKHasaD6ydCKalzXXYQbKwf6YE2ARjEDba7I
2bG0bIvX4BSvEGQIBoxh1AkJHPCwOU7Pi+KY3RbfueCPy0CIxqZtE82Jjrxf/8jE
YdIK8lSZXtF0ygpRr4iC7YyCoKtjKH6KhZsnV5eXoBiYWPU+1uTUIiCuVZWXcm8M
ev3DoGWgf6vXSbtNZdaluAD/4qaEKS8exFSwB1vLFfAcoPWRpo8Vak7Z4+atuZW5
ichnLtycM8aFSq6VsG81uXd5EQejhM/F2E9GPESSA1T3E5fR4uV/PdtYBAOqtdrE
Jj5XSJFeyfZJX29+Ftp+7/ixolH0X9sleS1PNk0uzVLUFsXRitf6MVj6iUZL9yYQ
EqQWrKCtWwBBRbIAiSWFfqTqNUZOnGtX7pvHNEkyXohmAX/bKWd1x5XzY2oAmTk0
tOZoZ7dUyT8+5ApqFbe8S13oXls3HeAEaPHeeWb1Bq6FRJZw0mZEpNeOiJmHwMqo
bclw5kHTQbia7mFgjzCn39f/wDwM/+JxwiYhkw9YEaGG6kNYg7CgSF8Os2VgzmvK
k/O/H8qpC2l728lQlZAvfjk8tgNkIHzas+XZFi099GuGId3s65Sc8cjm/JtXeqnb
t6e7dRs7c5VV5LsZ1oVuAVvl/1pBwzypWbo/lejZ3E717KButM+viQVvgVNVR8Q2
DYEGylBYutxh4QbFZupjtABrQERgUWJ7PNhcaxzxSGcTeFe92XKW0MXFGbO2acI2
W7e3UyWMr22TES1y82xzXqvhDC4NJ/TLaXAJEKCdnQautUtJ7mxUkorrHzltcyWo
gS3ao2KxspKsBdspPHAdgI0Je7QUKImsesEk11tqA8/GLUBAGa6y1B+meO6nTMyi
+yDhnhDYchOGanlhCPTgWBSA+cvlCNMRtld0G3VQn7q6ICcE3D4ceRLP8WYsZZI7
k/iixQ+fluqxYNVcbrMfwcT2tl+5N3I/XIKFHUyVZKjRVZN50iQNueFSVrYP5OEL
6nhMu+rwTHLaUTaTEybopZuPbSh2fjZYsq5YCjTuRJgb/YmFtQ+jUT1X+3ZO/v+/
Q/B5PJz/BP+QPp57ZUc4mKwlUIpPCeYWqpIHDDETzoEgwNZigTUdcI35r7hAUf1Z
dA9m56Fgw1907RR7NJnlDsiDThsBrSVxuzbLEx00BvFoD0jJGs4nQFSjPEQJ11sR
HR58kjKRamKEnjf8YTv4i7IeuEB33vBtDhubFThdyCsmEYfTZ/Z5FMgFbZ9h3FZV
dENC+iDVHoLvSYcpv0TS6j4TEfAZE5e0/a73I3oZkaoDYS/BPe+ihAPJvtSlR4yv
BA6Iozc9s+76W2X54noqXIDYzytg05Uegy71gJnG52bsoGnUiSj7+vUsgjI/Ehwc
TemEntZsRlZF4dz12QK/q8FdwvqGA7gWuKxDQE85IY+x63cQOhTKBQSyL9Iu6Q99
Aw59AXVLcC6/AWnhy2xoFbxZ2CwtDrGi0BijrIEw+R2tyAWCD+yXrlJySevJlb9D
XaZ4SDE5F+Ep4HG9cnl6ia2f4lEiaU+pt2LIlXb0V6Af7b2vLEoywhBSUq/6ksAD
saFCaVyhHQ5YVc6yDWxIuSY+UcwJGAIAUJBGpnV1tRI68ieWU1xJ27vvU5C8BfL5
KG4ezuPMu8H6vHqm+fvbTTlEjrui+uyap43hJXbgqKttb5wOzAYmmidQD/JDRXVx
T2+CCogE4FygZHRXOraRuVuP3gdSzZY54oevOo4H3rphfKcOU46cIqmTbP/RIDMg
saTmRvEjiZxVOdaecFGYCMlAcVapiHgFqNGZXFL1nIDTDCeJyR/z4V8TZd+HAZJU
czDLwyDQpyQcXAyP8Q1yGZLVEzwxpT7MzyleWD6m9NuYGOf5zQ8WJWecHJrXJwm/
o3hJO0N7TzxSaAAh0YfNHPm4fL+VB2ES2muOb0cJiks93LrgM/RDhUjH3HTqYJBS
8J6C9eDGGUno190ndhA0XBLqFd3IdPjzW5HIt4dHeZH3gcdyYGzuBo9UMRLmOIeo
bCwUA/SCrQHLck6YVAWgzx5XhDKzg7Y3feBEC+tO2ure7OWhANCBtq9u89qlwfH6
7cpsEPPd7xFVez7lJNa3vF8LAs31Gotuvi8v/azpkDTjIV1XDYVxWsdZ9wrEBHVJ
ROB3jp61Bp+B4aJsuxYBK5m4QQ4xIpQ6YL/su7mMmlAqx22Zg2Dy1yX8GkDUpnTn
2wo4Hb7DowxNToCJznowLgaXQurCH7YxrsvAl0sj+VFeEH+ZFHoNfGTy2TvJkLA6
GvUxJp64JQ7DSCkEFyX2GGkVGvoaKHS/ooPRLUwxncXp9JY+dsy0WPzOqCi1stoA
bNRjq5YoL6u8Sr0DXWe57jBfjMBCBinnA7+QXQD6J8yB7yTbew/GWDwuXr2d/IVN
O/D2Y6gu/K+2RQnVWwJ0uKpvEgcXF6qkSHGmqj0zz1HL/qbf2Zlhd0owTmP1yCno
OMxO+RmsyCQEpoUQpegwrhhejdX5t3uozNwjnvs8qs0N7Fn0glS2ebm+11udHfsf
aagWWN6eSKnLRat86D+DuMaWHERke71q4Ud71IVpkxPGeQ4FGzSbD5kJgg6TRZuZ
9EmPUF0WRYUSQfmNtDXOvvmV/m4EAE81/B+xlBOezRHDptUVzqpie4VQk7BcS4Jm
uOH+8bUBluCPydnTXmaIzG395wVU9zq09zPUu9YhStw/+MKeW0TuP0z3FhI+kDcf
xqzzAHFSwrBffxwS+eNI032mKm8x6oWwypmAuury7QKi5MwH8gJ2k5K8Rw0VcZL7
DtvQAtCGefpUuP91W7xtAn9NK9vWsVi6BoX3qfugoXhNLeE5loTWf//GfoRpZYvP
zTVN8o06J0Bjcrh4KWny3mjgBbox/URe8ZMix2QE6YqpeCFUjrQ+QDbOZnf2TfzM
OVfrWa2tC6oPcpWFEnz9tIAnqYs8BpNZdua7w3XIkR/YWFN3XCguvVSHTevvw6s2
A0JQnH+yAVG4qxXxn3/tIKWO22dCipgNjcdaE578Rrt5iVdZEcbpze5JGHC8dao/
ggTT85PV8HlU15rZIpmaIh4H6UBmGNqnpC17hYW9Ub23rLb5gEyHuFJPk3fSpdOD
/XRg7yhN6jP+kA9AdfHkAckKOIewcYpOAbLoU+7Xv+XmrTXoAHq0omXKBRX7ddik
vn00d+V9xoguvzrzlu6O+lcs7298cQLELHRrBS8miuAPW4C40zX2oZ4VikRKV3KT
eVCbgZXB6cys5e7tJLtzCKFE05wsMbUA96iPP23w4LJcMpBglZvvMuQSSxnqSMjt
qMXDLUfiXCvy9iyyYw4QcJSrSbPN4R44WhWaqdgUIAGVY3ecBmCi0fGCQbk9kVoj
0Q3DUP2o+wCfnbQ+cmLzWs+bM5oCgl/rWSDVz38lSAJNZxqtOOTS5NQuqUMrqkqg
+g7tz33Ix0Ml/t3gQIRwjeY6vwx/YlXwJP7bx0Mv2/Kq2Yy+Z7xf74JvfnbCT0Jf
Td+xGu9qjWs6xH25z7M7NlWDh79/g3jS435saXBucNCS5eoQAia2+g5BvUcpDXpq
nUxo7NzfBxd12Do3YCOpdo61hcgrZWxrWG567BtMrHvCk60+yHNWjbzoeh1LnB7R
sJrWX7KUIOK+tJBCzM8p9H8/h1sMHJFaqur90LZAgk/4UFbOPPidZ/oPzSxs1L02
5+O3P6kQlR2HLQgcyMMn6v+sycOn0xTf0JOz59T2SnsHxZz+eNLHVX4NRkyXOKCi
FZ9EasH/cbFoW3PMUnbwxgzI+XCaTQuk/IS+O166Yi6X/3s6v/IU7erHxuNgR/00
5R4KnbEwS7+rrzT5XDRsLXWy+816g0aF4rVj+ImHefDG6IxFWp0FGT1SeBkSJEWY
EXsY6Kkr7TP+z87Og/+FVzGQow7zSeejmUXA1xK3pbWphWcv+TvqrBL4+hbMMglP
U4ZeVgQwYNrbFrv0EtVUJKCRREJAcDYqovGOd1vN0wADjTqI00YutC8lwnD7eXwd
plj0n1a9uU7siYXvfEYyPL5HaGfVbgX2j8ngKH1/MLXZNY8koZA6hJFM2mCkxILp
UmWMrEce0HHkvzFYQd5RN5U1BIN3qOyfnwaIuLVo3H5T5DtHcHGc9uWGNW3wmecZ
ZMc5vbUU0yQinBD/v+4gCaISU+D4W2dFy7VAu2nFtA6d9V05UNMHV0+VFyo58T7e
fx3k+zRJJuLU846bkDm3QGWfuAyn7rnMV4JrPcGdBWikTnQG+5woLRQA/FA/aKdf
isdGlw/wsUPF8pqrf4+PznRwT4mBtNA+zTI9k/y28CWkXXSXfOoLpKH8dv8ctUGD
7oXYRpPitUJcTNX6k3mnMpR1UJ71/zpKvDGUsEmgLRm62EUEIKXJ6v/6wGGBez/H
Db/LN2Nxe0zm+gH0VqJtSoauGvXJnyag91UvOOYp/YVwVKvWgiw3U4tLyYxxC35o
7radWqomY2wpyvXTIkLfkGsTGvxC/NudAYeeEPdRxkxrIw+niymHs4CBwHFLQ66G
6FFEWm+SIQ7sid+4kOQvpSis/oVdD+qQ0P/PVWAwBCVEfX7LQ1r/NTTRzCdlIkjo
E8EwzUTZ5jDNZmtFmKLHJq0XLVs+gDav49KQCtaZ2B9eXwAnrFOHEzX6ny8t8lqd
IFGPN0hE75GkdVnFBPUptKsVf0PTGFR9z6F7k895RXjkfp0CC9QBO5ar5htdenmT
5L1v0KU7a3j3hjXqftG6VJxfk1jkW5XZ+m4sHFSM8bRIMqlOCwIT91q8Vrv+aWGC
LD/d+nKoFeFpNCga4lGd7t4lEDrEMieXM+cn+9+H3V1qPF1ByRxK82SHVtLyPvRQ
opLkE9LNYpsT3ZaXZuxWf+ZrPu1O5FboKJefUwhmeli1zEHwQOGXwS5LNN7dz1is
szLOMZWGdz5T7z0cuwsjgr6GhSeKy8uSBDkCtUUlZj22YdZek/YFhduE+J/PTaYI
FMtOlZbFj0+DQVYCFGo+QAFsTR/vprUNyRT8bCxuWvtDF5I/UJQVcoXDIgLIyUu/
1FoWmLmcxTYoHn646aVlWnp+ztPIFnxIL3RkHdviVLGEx7iin4tQoi3kn8TuDqEH
lM+eFzydK5Pb9fznKzdtpCrzbaUSYyz+tXC/zinkexOEZ6eIFbCc4wA1DhcpLKhQ
/bF/WajsbqcSZQzlXuq0lDyifQ5q+7zAc94hC2j3B5fQXfZ/gujouS9419c1dOur
XMJQak4O8rUH1DPUCyJlzIrshtzyJrAXR2pf/ndr9K5JHvtWDVCzoMMtuOYJpT1w
tDKvxXTilkY7I1uDSUd9DxcBJekjgNaMCVzHxVNPIZUHCdcVwC5kDu5avgM8PFR3
JghXe+8tiG2WlwaHRG1toxrevuB8swZicKaeLGsKzh1Wi7hUFoZu9LBXaKRRbM1u
wB2LPVahhe/TQmXirjbJ6Yi8lYye/NfXzAJ8U04mVUAtylzsSktUelH73LrYxi1u
02Wfpm7LXxYv6T6q2SDzufSH4/t5fPLmjv1yXJZC8wXGBaGUJz0QEZfj+mqCB3aq
SsEgCZsOAdt67I01wmA8KYD0lzHcdr5hjAP239FNAbBsr+ZYtzdue5S9kOBo7Hcq
sShaMijC6oi4MJBUTp+ZFh25j01i3ilu7ygIvavTYg45NWOPEfaF/t1CRjncP4Im
hfbvmHF0XYGk/KAcxOBN5BOH72x2e1a4BKGa6O+U/tO9g8NDjy23+WfBRQK0MwZr
fR4YsAWUQcyXiwiuGxSr1pfPH/dADkEPUV4z+D8LwAge1aetVEpXUHD8UU8RZn5v
5EKzij9TSUDESrvAZU18IBnKJvs3YzmXuQ5xg6RxpAF2HsUSOtTc9YwxeFqtUFs3
OogGyaeNQYFJR/tsncW8v6zG/8PkvyZz9aNJIjFh8uJcTUPcRQ9KSvO8ti5YlWua
LqFEO/o9UG1b7ViFkWkF13GFPf2UFpfg8LDLk8WQKxqA4TeNfkX67VAXnDcZktBa
LAkoPpV67E1heQTlOxB5K+Qpva6ieHn4kfDTrYXNV/HaEPeR5qzRqwNeMQfQbosa
1KYWvPObhT9MMTJ591QEAf80rlV8RVWn5FUd+72S1i0WbGRxan5fWldh1DXGxXeq
iWX7c+/Hmta/VXyIOIdvWhARI0HMfRWaF9gVZl5eF1QDxceHXLkYpobreEQqMor/
eZQ+MiRB5y4y9XVZWZoLdayArGpCrRvQ6sS8cTvMCm35Zfd9L+yp5M5n8+IKufq7
5t+Tb3VFaVbL+Kie6CgPa6u4gMIx4baAYNP9T2cIOtnS/4K5ASGnctsVJOIrKgs9
4NRKzQpsKjCXpVOdD7bUdEtkOP2p5sJgpFPE5MOb0JOEW/kL+aE62mGKixJ/mgcV
D2nfMEYO5a6abMwhtkYgh/JOBrv+qOf4TYyvxlk6g3dqQZk6lolq5yv+bmMMDSpE
5+tATlms9Ynlh8jIdiQ8qMk4siUeqBA4E/lP3wd0KVonxqaUcwXNMDuT4BzR1Td1
bUzDNwecoTcMO39FQDhjUEQp7a1ekgQeZC62n9TQ0RBQS37BNAFipe8mv3afiQBN
FFWzGVkTCMcF3HRmytUMMjUsWlaK6xdFykibJ7EmfEPVWZ9jaSNo0Oq63PZ9qduB
BY6AvvkpGUXsMUMQ6rWos2ySGdAQHy2wqYlMJrDDr9jRkzETxNRfmXkk4RkR5xis
CDe5LSmCCdNTlMyjpNALVbqO0UAZ4CzHuGXtRYQR5cle0A63T41kYeiWDidqPwZk
DzLjxzkUmZejlwtDLZ15B2lCIct22x/hkoS9NwNnI4Tu70U1wG9hyItYi8jNLrn6
/qWr+hjss2FPCy53S3BocZqQOX9GgKZoUNGw7vhpCC7PUPBWQbszrNsqSAf9JK5i
3iTBjkX1R6FUYcyZsU5YTZam+O4PBBJ4O815LSdPrwPIQ8LWE/KORXgCbyzTngC1
I+slgFDfq2NgJcNjSJpvcyDs1M23F3TPaLXgF+CBEQ+BUKOaENmr0bP8H6Sk2kFW
d2EKUzvkxqRBifsUihOaAl1Htk7Ij3zCyk7aMkUW0kacpeJu6U+wo2hr2+EqJ1vh
D4BeRut/0pRQO+/b0iJ/QmcWi4OPWVCBWjhsaCLeVBtnSAFQhM6VL4eWN6YfU2ef
3oXDG8iF0H/GRGYDLESlxleecho/j0/JBs+AiU3VWYw0jspp9LI6yOO9QOMhQvtW
O8txzQ7ratqShxfN0/iT3+6YALse8JMiEBOpoQ9iC5ttoRdGPq4RS3idP3ZV3wZd
Va3dTDDsickeNdRME/Hbl0eJ7hbVOFfIWSmyZ9ZAOsCawWE9KntmPgNYmHiYbRDn
TZDBQc9IOx3HNHTjBDwHq90WeZe0hZ2Roer0eP/gHx01MnmRKtWPniw37VPQ/qjo
oDEGRwgSkNKBNvhh5qCizH6fJT5Fdsky6hdVR5f7/1mmeii3d0kYz+96SeBocCm6
Lbm6bzDNJO464JDYGyHQDfJEgGeUNmh4YRBZhJsdRbPYXcYXbuUcStJaDPxC4o+v
rgoqFirG2U/vaqhq2VSyqv8Vt+tiErFsyO7GUAm0O4sZAvYm4R/f7RxrJVjTgZJF
YxmRgm3/6llQJywMvo8lgo5+A504LhoPE/vJ3LcSXDKksLhpRP609epyLgIOFqmr
htek6Bez2rhdGCWY6IZjCgbLXmdYjNv6XkcTL6o0jixBOzJrZ8pktSJ/OVdOrN+Z
J56F9788sol1J0SM2pwWvikyHXssXwlC/uwjcitrxEvPcCFn2cB1cy8C3JndBwcj
HUvQTHv8NPrUZJe8yFLhcdaM035NE1OOW0POB0fJm/DpBfQV6xmHOxFtjuboP58D
cZKRnwYRuD5R/5lbZDfE6ENVoCwQBRMi05u2mWJ/5YG08nbMY9zl8ulS/qBinePW
ZSA8nx+hUFbFuKdhvRVQIpjXpZaskNJIWhOweijB2sX5Jvn0QvO6N0mAKtW6wDgn
8GTvuaER80NBtPXZk3FZmgtTdeQjzrCToqIGRo8WUUNyNena0chrCe4My2HLuPI8
zStVElMR+UQ9lXok2Xy+PSoBEXoVvJV9+uZ/+imc12cxs2dZBDhwLzxlOHrJwUqe
KCqKwkvVp8zuZxX6279L8NTxRAnxYpuPmU7pV4eEHf8UVSCrL+kCveq2Z69E8yTj
y2NZxE+atperSbVW1se4IN0uBSoaHRabaO1AdfiWYdNLvdSFEZw+9HQ/292+3s2a
whZqqac/DFlE/GesvHY06D2JwSNG50kP45B1uUvkY/ZcpELZm1O4A2FGkQcfLQJb
i3pxpDN11/MYOkJy1884HaNuneojUKx8te2pwNqJcDYsE+r7/Y8XN42ofSB3TYrp
zhVi1sz6ZhFXsk4EU0zTFZJRU2l1rBlgzqGzyUAgfwQB2kfIXqOYqtgcAfcQij2Z
vU+971S+yf2CsP0exdOzJNzquIftgJjbcw3MYgRNzk6Mh7b1MWhlgePSEx8yFNpv
s/95nGmh8aHEFQekg9tP5xBvuH1SHJVbExk30inZOXmuu3k4molQz/10fD8ddovV
h+PNF24usFEcMU7wQ683DHOxF3lDIS4mopDdmU/eSRwRriTaUsHMziZNYCctYUKi
CH/pdGfHbAo95+cy8L2U5PE7qZzsf5/PRB1ZvI+H1EbhW9PCo40ZSWv4KG/8MWG8
XQcrOa5KUFWfkUAMPLSUAzK9f7YvXG3kG4qoDla8xStojdeXg10yICtpaflZmOqG
wgG2jhNwqIZ/wrKgeTsTkkXxq4KRqLeAdoGviqnRabhsyn09QoMMSGpa0P3P/Yks
7ntU40NcFsk6l7QqyJFkFtY3RI8GLBpFkw/K0KbiUanL6pN1xC3Z4cRMYNPIgG1D
YPgZpbmvpArlUY8vnMNwP+0vwKxSd/cQfo0sldy6DtsPEwWsjcAx71YnOkkZgzH6
OGc1KsIdeVFG1ikqmcjF3Pq0Y9QMuiNc0/bArHhQT5PfPLWWI+B79NGLXPR2OPj1
5JvCL2+9TObLCjUu97OPac6awaHkGutZ8QYj9tDzVvMt8N+8b8Y8h2303a49H2VX
a4y7PYM4dQoOirHhygBl4/OOmOsoM2rzJQhIkyzr52K8WAjtLRY07EMaUtsRQO7F
DY/oLGO5GMWfxHWEtnULVGmPjn9yyGjsfqzDld+EkaCYjRvJzhpHdhrwiKI1Xrnl
YFfR6SawUCpxzdnlCtebY0yINjHmKq7wYrN7AgXUl2+qQgIb7B3dFscjFAESn+ui
9s9A4HncILxpYY0sC8AlBGO8Q8Hf1d9lVOw1jnldAn01ogqQf4hgrG9w0yO8qK++
GaSdqxkuJlpga6zmVPxrvSpxFmBsJ9vjwusXWJ9j6gCR4CHtAETB8g60Qsi9QgwQ
0WeHTU6HBzWrksHyKbzoIepNCgoYcwaMogh7y2snjSv9VUNsBReQsQDy6CsgZgBZ
8eNW/M+k4EohzXAqA+3jQUxl0BZ4pksBdgvOAPYF1I7lCmd4x7fObe7bgZqzqGvP
Mng1PNPcJ3oS5vUCENVrsljHkK6A0OqPH1PFmHwpSEV22ws3z49h4WlRIkOcLY/p
g0LgQmzrgj+AJ08FxoeEq45AUNSRIXrThWj2/UEm7eZxAbwgHA3LWi82L0wMUI4b
yPwzEDnZVHxHfH29qpj4kdoFiM/shBJ63aQDiYnyIxNWkippch3egyu//UjvrVOn
m811zGvo9Me0FmkCfJv7WHG6K+7l8Z7hctEvuLwoB54lQWhQIDFKghmiHPtE4x94
OFmG9xMocqSarSFc6ulgFYGX59maXz8q6iga8Wd5YGbZndsmTB2L2u//pWnVMC3T
Twn3wZXzDCa5efq+9MGxahOm0Zk8SKpAYib+b15sJHqTuRh67Nj9G/K8iIp7ZKab
udwlfIWArW0v5HwMUINlas+OHeGKsGH1JTHmz+stC5zpBnWNLGOflwL7TQF0BVvG
U5GCq17J3oobHcCSqX8ePxa20PWFLWNaSm3XyB8AXiXuz5NYiU21eYKuOxrWshUZ
JX0dp4TF71CDzbUNujtIFKjK7ZewcAhk4LSp1DURRNFsr5K+dG1U+dZgQU7gVFiZ
G5bRp0PcjQa/EP5RyPhUoHD25SaG1nFndHqMUrC48foclE/ZoZKK19b6d4MKz9OW
aOP334zqkWf0Dlh+jGUaneJrprO2Ej4bzx7wpZmG67NPoRhvhZx8Tmy7ZQEuI7oB
Xd8nn+A36z5bgIW1F4r4I+RJ9p43LFtPxaVWkyG2dkTzekkUnBvExzXGgsu2D9Gj
e19TzTj22j/YbDWeKRIjkLz7Ubge5PMNVhioQFoDYhcv96atffKecJ5uD1k++Zb0
/Pe+k29Tri5+EeSaXBH1l1GzJwfAuLHlCxtALxtQJizRE7RY12T5HYyfx1As9C4J
dLgzRG83VmMWfxBi7UxHUzoMqc84zHctNAk+0RWFn9KZvEcYqKygnmU+UPnMy01D
TDkszptSr30gzFvY2awoGARSCzES/NM9JdmHdhmJBmzX2XGWMjUPaYAEVluLKY1b
zN7+MZxaTSVWlaF8iiuauC+DnhTk3ClYOr6vE3E7/f/6vAkLvhzPFUpZIcRSe77Q
jhbZM+PVlgds9qWkC6TRi1o411zps/1pkBN0nkw9v8f5OgFcTincY7Sd+CHm9nF7
4nybeh4I6d1NL9cWp92dx5NRw4h2N5/F1UTybVRsIZmxKci7tiBrwe7TA33KwAQy
wWjPNUz8OqbSJbFWpR6D+hrdawWVO6jI3MaTj3m8pIPxDe+HA4LIgdzKoZD5jpTi
D8VRGhfWDsH4fBue9w8G42aJD08cUKxbJdyPUyN08cd7kR4XUFrPXe6JDFqBnmnk
UlzXCyWC8nqMtjxdTMft62m3hnYmxMHduFZ6l0QTsnjztwp8GxfksQw2bSdgbeam
EoqMHi0ad3vksZmfyZiy5vG6jQp3jMdHjqBRNgXwv6AxENlAPYzuTufQ8lPAD3Dc
VwXQOFQG7IVVPWZ40RaLnjk7ZVnPpzjVzLITQaWxcOPTa3LVXr/Xwv1QwfMsrRK9
1k4hJh3xujvo0uWuAbl9OWtAlqrh18ywJiunB41JWlj+0adxv461OaclVGWS0B2l
uDrAUDJdPIwf7M8k74Ivs9uzBoASDcccFNqFRAhRJWvbqiygd7fR9R+WrzhwUNW3
Q3fCLKDAl05afju8zzQLkCUAqpM1AtUazJgcygQaXCXArM30OTjf2xc16Jnih6+t
3alfPTvmWbGcFCSHH6dpIz/rDcQCtJaNSVlb3P/UAiA9y4/CHR/UATsSJFHerk/W
xm5Aw48L+Jw20TUfmq3ywHPOdznPyg3gT+BeYKGlLN7WJ7Xb1/DbWD2zdXhevKNF
oEzGhu4geJDbM/ws+G8QkBdL7dlwBwkDKPmX+4/Vlb8hkbYhmVtbJnsdJcWS+fUV
rlwQn+sr9WR9w3t0JX5zp1PqpAhOTWaDDZwla7EYAzCZoZ8zIocJ+h7xGyLLG+5R
uJRCIDaWL0zmaOfZ08iDucauqZBeM0O/EVRRVB5ctApMn9TiZJBmSiynobGJ36Oj
BTSVEro9N0gCv3qNb6wsnUqcTnMdk2ocJqHLrEbyOVy76jQkvwQ4nXsoyz5FJoJv
OlM0vqxWMT1lEyyDLkK2iKvT1qadIY5iiMAw1X0dZvOccT+7g9yW5xA7NClTznnO
KNdEaQY5LZo4/8smZa9YXhXnEnf/wHToM+Z7iqRmOOSxfjMsCqHImGqgnIsOHtqA
lV3QlVXpGSJl7wD2Lq0SrpjN95Fe1PNKifUBm6K6G6qhjdjJAcajskMY6hKfuy0a
SZ56nTMYPbzZMOCBTOoE8m0MkokN/wggiKM61urYoDPrtkVmI44d1S2qBdawkula
t4iTtj//s0f9ANeOCTwrf5vaxIe0Kwwzi10sY5BsN5yu53BkpFk0YxhehPwAi4kP
Ilzofuq34b2dyh4n+YpBoJYicbASV15GC3ybdOFgatddZglJZTQlxzjdCK0SIqev
74BsjHv3J2AFBDOZIw5m82eNCgZZCjpGjnP5ylFt4QtRgQNVowreBOA6LWxvqDDY
NgFsaDZ0ZUJ6zMECtJbstxmvjI6LQDGN6xS8CC+bxOl4ra0e4w9qpuEuVFy/FM69
3HEv/BjSq0Ih9LjjfzFG4k4Msi+9FKQOrqQCPndR7KWtJVz0Gt6BtJFQvg3nT18H
86Ksl6ItPhdNtsJoz0ImKeydR9iqu8g2Ncvkk3iV7x3CQ+NSPGckJcYJNJHwLHF3
4NVt7yaCjht3r+/qzw/uhy9gMy+aHVypt74Sw7Syli9eHn+nY57ZPHUzULmQPhS2
YwpnM9CmXYzn3dzzM2Dm/mSA32mde8AXzFf4tABpwilKIB06gVOJ+igNT3QGJehL
Kaog3eLMlmOxpIRUydsld8NwhkzHP8TTqLugzga4cMniTdWbsb25RUT4S7EIaUks
gsGEMCOZ6MfFYCCs0J+D/m29u7/OFfCkeuAvl3Ng+dLoX8hsIseDzCnr+69iUA03
wa0M8+2yJjPXGR0qq/yIqu5sY7jKc8c5K25E7p6j5B6PmjMcU+GIMfpAB1QwWc8P
pNINFqc29iVnIAcku5Fin2MCZGkBCnh3YNwMKadhpW4f8AJh6vV+5iWa13EbPwE8
E2ftMPbZdzOVpam2HcXAIRkWup6tWN9mrKsEABJAdGCy2piJUIEGg2t/1y8+4p7E
J9HlzeHhrXGasjHKyyoMG3+SrLZxBsfMpa6SVB4lF2c0d6XzaFvc8MjRpLxpWtvx
uqbZZfUfwhzS9OhUNZGcX+Vs99viqsLFIqHrIG04Jr09YWHapDC6IBKmPEyMFxpJ
zY8CirfGkoZBWl8WxiLIbEYRuNA4YYkQo0WRdy90+WhvLDF/hXzJj2TUB2p7x1Ay
0etIYPuxxpmyKJpd4XpQwfib1PC7ao0opS/E9IkXmIxuQBeOzrufNdrtBed+RMPl
YslkBN0rhxuJ0Dfe3iVDLVrbir3+uwRditNfQF/Lt7xPh+351UixuVIyWy7gjwtL
r4fAlKXl1yAQA0sAV0sWmy0jxdrrHC8a3//zaAIVXMUJ/rJZh5OxMsbi26bC0+wI
oSEbtKbRPYpUU3L07h0gFCZQkqz6CjsYy8t0tuzI7H8ccaIe5tW9turgymzMPVAM
FV9ahCVVAfkM9LH/UiWQqiSmOiMLx1rA7XMT55+6NTt7VKE30TvSfsgpzkWQa8Jb
E2CMQ+YiP9y7njOOfQEEwuikPvMCnSa68hUBPdvSJzKG15ZYf5Ryvw1ZWEA64gut
Dk/eAmb3hPioGYmft9TROIT8isFd9M0d25lObgFD17nQnZOZSmv2NDnZUaICymBd
s6xSwIZnaDqFEIrWKxwPTvq+jaE5t5Ydf1qBAWd20CJCoXz7cgumFJ6aoPoQNDhX
SnOxi/KSzqANi+u7RCYvmlqnclBOUJ22sz4sRingq8T6e0tVxNT1IspY48FrkK10
f+odSAuRHzDjrCQnaqLE/u5iyXqJTcfiONX0MeZ3qZQFqlnfX2imtPzgn7ixjXgc
Fd9vqfxeSi/S1TTwK+qpYl9AUVJ2MdQo2rYw4sIjtPSx16UAqRvShMcKpEc1VeA/
C2uKB4WceD9ahB87V/Xu2IHqg9ScekmayoTiZz6FZXLhkXbbpXVZsAnosh/Kq+Wm
19pjf6c0O5PL2TtNIPrWdk0/VjYdGhLy9SaXTfF0DyGe6Lx0fx6weOzimnZAsAzn
jNj2/Jrv+uxLtq5JwVKFIrXGgaxzsCA9EnYMobftvjvAo3T2J0wbuFlLq4du6jZm
p0VON6GRr5kxG4rBB8Qeass3BN41gO3wEoaF+Xq/utHFQGe20Y26yILsxEXjdpMe
SZVaQcUyvMHV39GH5zsztABXnLeiEwK4GgK/I/+Z7HQp1sw8FZX5w8Rr9d3Sq95v
Oap019/7ja4jU4zxPeQ5l/vfCBW3MoWzz+BAImZ2UPbGhdTE9bjYBMb7I8HJN36d
LPtriO8eE2yPOIdmhhb3SjbUEvCkqKp9qVeJ17tTvT0Ct+qUf9ECc0t9IwXUoSRH
l9q4LJhdMu5iuAG9bndLXxDY7/cVCFMOa9sn/nuyAbBXNvKFD1IyYY6AAJhum/19
QqfKlrP6lYzhr52cT6zrs9O4w2jfJRp4Gk4R3CUMhy0LaCbOdnGahLXurDjzTffb
gpGtRLl94NPspmXIWZkg9jw1FvGXClYmIRMWQV3yTaoLinSIpXL/c+hxlkgvXJzR
BpyWv9/3BPKlPmyRM6Z+Bi4CMtUUz0fBFykpWT6DnBhSKsaxxr3FK24JaqsccQtJ
mkCXir2H7R8/gshyDd4WHlo+P6U24WQVrnu2clmSUBVSZc017xaG23nN3yuQcJ5X
aZDmMjmpWZSmKmh2Pc/y4s3Yotq9Rq5xT8AKzTAFE6P7xtMrLwewL/kCYRQPZQkz
DcVCyOvXN5LO04CQ4Q+OJEqaL+OGWqJ8hSAmAVb/0yu4wjxRCMwJWwnVQ4vrZHth
7HtfcvHAKHyFRsN9JLN/55h3161GcTYvZCy5x6DvyEJC5OJAbX7ODIl3Q5x+Hiqd
V8UsK3vkeHhyLqePCwo/Ilp6XhscbEEk4ADBa9zH3WP2jnW64SjL79+3bqy66Xql
46XkEyZdhGz2QT/5LuVhekerh+Qz7N1Juyo+FXXxUlsASRZBl9Ootat77vp+GPQo
L6+Oj0l7O5zcuQl5aCaTXZJd3omKOkqlw5iuhyPCwaGcbrNsIsn4Phli+e1owmW8
v7kj4hKirKWQR0PqrVwkom/qVnQ8qTtM/JAeALI3Tsh2ksfrYxBM36X2vyA2D2gO
cK8M4NTp6mMIKh7/Zs98m4IdjbG5gANwTHE9vDAR+2Eg+rXvn3XTOctw5DCiJXok
k1HHFjPjgr6Ahe55IUvXpNMFjefYz5lyBRsEOIzh1BQqzqkd/MHv9awpBeWe2gBi
6AetWvUk/A5Tqz2WQf+pbf6ayk16HcCzxyD0Froobr0WIJWVtNOFFEMmGOEakIgi
vvFt4F5ZVLWMTV8KN7YeGHFw72qusO0nOFe5TcFFnWJAs/Cv8vwlT4l2ELjwXkNf
MYAfRumeKxWIlC29MeGtFMAdrj3QAp9bTywKKxXG3c8B9Y8CJxtTK7NDjGhla4To
otUzR4uB2P03HJ+WUk9Iwd6HuFcKTgyFyarchHx36xeIue6vaU0AQsfoSbxHMWmv
v5YeShETWIfJET2EN1NLgFAz6W8FJnYDuhjzvUSRaMO3PUuPOL8LDb3UNTPqrv2A
mfSqXIyomHAbg/EP4tmVEhSiX11k6c7HGge6+KItfvDN5Yyhzk0WcrdxOWIeX2T7
KPAW2ntA1fzCh3Fk0nfUyALx2/2mpx4n+3TX/w646GLK8EOm+PJFa8QB46dacxB9
5NNc7nl76vQ18dm9iSIVL0nP0rUmWHnP850+gO5WR9qlQ1lNaiW3GEh69FsV51BT
6nXm/lUEaF6UXNSBEzAt4Zi4fr3dpYAYWDij3WOyEmqPyUt7O9Sr5fLTZCZdp235
m+lmG/2GxpdIrKgDg9tELfkY+bUUi7MOhcistusHaBKarlFZbpodTA5QyOjIT/NB
gUfMpBPLpVRI/55ThVrSeMQ+7oApRZMzwv/1bvl0WtFFKcKkW+j0brvyPKk+ZXEx
I3R5gyDrkJ+5A8eDI0q2HMEIRz/MCKjSxpkhom/wmg4RHHeoUdtH6mKe27+2mWAM
A7ixOBPqPCZtdkEtUb36L4vatmvWuiGVGlhjOICBPeECtbFnfhgWuGJu4bthJzAQ
TvhEHEkMy8dnjw5K/ixzt8R5ulBEocvSyTOEuaypXB6lKjo7kO3GmJL01k6Xdlfs
X3TdSjNNiE+vUGLfTVcDqM9VDIZTE5GH3ACP5V4qNbwp6VXlKK2daMt2354+/7I/
qb2hFbPdOwu0zw5F6sigCN8juVEQdgA1E4JXM51j8TimSpz853GX6gxJjK7Gm7SU
9cPmuqOYPM2ftoWjyzmneYqwHakjlZ2pKRCSuVxywmHxyk+gIdcmW1KvkACCkZqU
I/vLRkzrTUpUkMJZqNLTP8ciVOztL1U/QaqR0UcYMfJ1NTAQaDkA3hfIL6WTm8Qz
atGr1WRBWZlX0FMxiDgTYW2x591yz+PRSMCOHaTEc7lAE4QH4dgs5ws1/YyvvjjB
qdkwwjgpT2V6MeWQnPxKNqU28AYtoyINOcJfsPpG/e4mCa1l+sMLJXGYuC2Gx0Tv
xDqeDMaW9q+rlmOQ2hdnS4MeK51+ab8V1QF3+75DYE0HsAHeP2tqNDr9UqOsbRzW
Sl8nDKo2yN9KIbb5fmvvF+NcFoRWeZj7eeiIOigERDe0LGnqyTjQO1KNse4N/7I1
mjRVudNbhY4tSgAgn3ttt6AcliYqR2cGnC7zA3TTvg0PFGJ1A/Toncdxcm+XW1pj
pZYMXed+Tj2nbHjBr+SB7v9QXSJBi0keRYfMXJfbKRXftgOlP2xA9WZHANieGBQe
UhN4rJ9OWyiuXYVu8zNhzIHcgFigGZtV+oat5tdCKDTLIU3Dk2VCPV2e4FevlUl5
4cTSy/aP92EK1HZX+ZBG5YkSQtyvfg8VQqVs0ZWCZP+fMI5BQnBh9ZBAIVq2vm6c
gwX71b+Dj7fncNOqJ/KudJFz4J/ckPlCVjewScRx8+j2Z4YFA7m0KuTgOTWtxmCv
B/Y9DHXJ4nf4Z0uIUyQQVum/6tp+9p8taDfZQLeQ7ehoV9cqWXyVUoghPdjzDJ3l
vrnRqM75glFQus8rss9cvpAfTLyFmnUKkXN+pRdUTmxlLb9fBKSJSDkSwaC0kMDW
THOh4Tg7v90BRs3KEMpZ1/i6vX1cw5UMTI2NGqtVFy3mDONv8lPIzh/wDkknYaje
llCqF3AXuf8RyO1PWUhKBQFGRiU8NA4KXd9tpP1u/+XT0VsgPrtU/aZ6Pjgy8/Cb
GXGS7zPl77NHl+KLFpyWrms38leNdrOLuvrBV7d3KiRpRleYEI7ep44M5kzy4WH3
ycLUwfu1qQHxhlMFT1gheEslU0oKaXMhcsZRHcn1UJh4fPXvkRCwsw6C805tSyBi
yVAyfimXwn2CJPdccFHMYrcte0GaxPd7qEx3pgaaCMZRAx83ttGrVYDvEIXGOQzk
r9edXLO9sxvjU06zl7J2rzSfc6bKtIliQ3Y1DKHZMpvd5Srr5ZHokfGo30OiaaB5
eYvnugro7mOgOiLW3mpfSUdJY/gQ40E1DNGAyfgMIIqvSXWHberif91Pg2jO0FEk
drxmiWyRWGZlxehgpWWLf2s8OXRLly3l+3ZlWFJi9nN3j1WW6eLJhJz/4Vhk99iq
BC0BYfUkuMgN6uakdUDIjws5wMXAN5aXyNzTa77WnteQK0+AiXEcbroKBoJyFC1W
W0+lLxNfJDiIYkTaGr5nc1oaGkvcjD0iAWspNWt4EFY2LgeCpfmoSZaI9zq3uFc0
4ce7Tw6jSp4FOLOFt/lNLXut+ZAQvn5n8mO98rXIOAmg5VPp63eqZ1hVASRqsfnp
EJd1/JXy8LutwBAwnJT3HdZ68QS+XrsF0gJZsVOqKflgI5aYNA4R/UqT+DNi2uOw
49gdUUMh+IXJEXQML3bU2U09jvOZv/h3FAf9QZNw7PTebzHpcXzBFt1ixbsDsPdT
+a8HmYo3yMK3y2ql4TywqvXvHwIiMOS86tKW6FLei9hLmhFJ+b5VtobC8chy0PSL
ZfxSIqb4wK6HC2G1cuSUg06XFD9CknLhIe44Q8+0mI3mv1PuSXhEa946gR0EbUuW
mRHvHLSshojqL0RiT93r82hAVuLvphhWo4GHyKgaV51/RDK6F2xkokVr2cJV2oHv
RwQWKIPZP4puoPefL0fNr2yJVmsJnu1fCvt93hHPukxSljAcqp+9+xSRapifpWTK
gQa2XmVmeLVFG7mRNbHCgg4R6sn6XI7LGT9n+0vsfIhWJum3ss/L8aCgwZ3HGe8x
T2zNnaSg/l/gSTX6xIdVqVZ/pGi0iUrpM1NVHnybkSc6wWdpKucuWut2lIC6YmVh
Xk7IWWn2OJaWDXs/kY20o95C/4xs22X/34tLikqoxRtZO56s1J7imNpMRzRf6NUz
/y52FAgeeIxrtwtLIP/TeN5Xi/D229JSsPBa1abHHCqgvYO4lVkX4URVWnzcJDsk
pHVLhpS8eXRxDIoZtBcrMm+f/xj2CYUhdommrKXYfQUHpoCxxUGh8L9PZAlsMkV/
YtXPmOP6rzWZ0TAv+jrV/OScEG5aEmHgdEvCA+nWIDwgviK6Q/QSdML8U7woDtpy
o9RmlD/7nCw8N6Xf/sl2rMxWO8UepYH9QpL0KT7N9VxP/zckXlIcFIyTtDqOOUNR
9DIOmmLVVPZ+9wPoL1ELR6IpxK75PtkBVwd3jdUJEuxnw2r9PgibjPGhC+YuVeMU
TYGoC+6MmL+ucCjsYtmlimp0zE3Q+hA3fS41LO6yFrzo7rrW5qOHPiyC3uzHS9Lx
HeNwsL3HjuOach5tXv5B1ndsCOM7r0QpcAoeY0KFq/+NVi4X0Vz7LTWM09vvixxI
GbM9uaJ/TEvYeLCNDt64zgp7cDWFj0PhfG52BPHUUOX0NmkRG27Dw5Gn0lv943FQ
vOoxN3PRyBh3XHtWbddxo7ir9B6mgLJZCpAb4BqHwGqLGPcEvdl4fwtvbiJD14sy
aujwVl2KZGzCK2ebnmg/LBb/mjvUmsgyxn7R4ahXtB21M6qGwMC1Ejb+DJ6sZzz5
nPvcCACJkh4smvKihbplApLMe/MPhoWMd8qI5YoswBbZvIRkbYXpEbSKp+YMzdk+
o5ZOOxEqITitca+v7SVHhELOEDQU6BkhVeSgdfKjz6pMUPKMFFxPqwxk2SGb/pw3
GHD/tCb5YKMZfPWTgb/K6yxEM0d/jNTGXVqKXvI4A/1RO5q7F9V8+RlO+FxmJaC8
xMa23Mkpf8eKLk+tna+2ZOYYm2zdJHUOzWwQkZf7YghZe/OWWXiD4xgYls8//Ins
H5B3dLIV/Hr5F6U4k2+LdRM1k6XsIvfXqjzYI2rYMp/5U3t7NYYvrTWa9tzicthS
OBnj+SRkOgRFBpHWTvfY0WvKdfP7Sv4UXnrD3NGyw6kTGNDg7lt/te1pgUlxdAyf
+LfBioXk5IZCGoQ7ItkyG7rhJJaWrs67J7fH37XiqQLq9iz65M+hOA2irpoL8Dql
9/dxs3ETRZu15La5poOnXU/gEToTI1P2mDLXDG46l90G2cr/RQgat5OsM58oz/SO
XJVns0G0bAoNCCnh76spiekpM4C+YKSr/mE9c5C73tkeaYVGqN1Z7XHWGFJ1opsS
bPkxmq5T7hxHyY5CobpRHszl+jbQ5028eG8dYiua8BVEq2SudJWk52q0KUIJReYs
fxRTlsbtKJaGZP0Zz94V02VPTbYcaBdT3sg1h9ygodAV42FM20cXkzs6z1NZmFCq
8Kd4Rsr2tHsP+kCO0+eg/XoeYqvXvsOEJG3zUUt+orD5jzf5jOAf8RoIaM9vy20b
071994jNohoBbILeUahtM/SYeQMxzKCCfzJqrMYV12ATycrueil5A3ahiBirrTvu
SMOvC4GAoC+Wqv3u4DTUzWEb0MO72mnWgqHMWulKjQuZ6ViteX4BEeAfxA8mnDjN
o3DqyQWXPxj+358YJo9b8YFP24OPQnqcXW+cMv/jpwp/mW+tcFyYVW1tGzCjdeJx
T5/RVsuf9GGfG4MW4Bhkc71vMHd41TWEMDLFK8iAjGcU8eOGbZX1Al6buJw4R4ux
sWZL1/7C7SoVbSO4PzErDwNpgSJW2kYJXOGR/EL1tGrK5YFnHXTcwcM0Bmolhvgk
5NUBPTh2cYJ1tDapgvK2AqOxIOhPPb8H/AMqYu5mWeC4k1EcTHrV7/M2YLgcIRC2
qd9h4VsHr60I3MFymkzAYjaYPLuJwtT5DeJbrM4R/6Oan+WeQY1zzaPYJyfzftiq
c4KZ3fx9TlEywYlcolzrUU7A2SjVwr9rAQ1nh04aJYT5ucKfofufjXwsmLIFiVqd
2ToCAb+09ewxq8kGc5B3ly6lsVpH/OPOKqrEc8GdNcwxvkieUowOmmnA9wFZSEip
DhvD8AN2EMJAIP7H4Xb38aWyosioF3LryGeMJL+CawBn/gaW9mxULeZPe6i5RqFG
luNC+InVBgX3B1ql/4tqgj50POK/27WxLngTgInu4BbqJzlTyzXDGKPhnU8PWuV3
K90qCHH7AyuPcktobqHUffsnPslov1N1jSHr2EmfwUwtGJPAqb8cW/YzDbOqApyX
asxnFlO55At41NfHDIE5H9cabSwTNvb8J3k2BSoGvhVGqUKmqpMXnnUUFrK9pP87
HcAXIbW/3HMKHbOHQjE1WevK0O5Xbuv58asheKjOISz0c/bxekvEUJg1M2MHQNT+
URFe/3EIfKQSntdJCm3Csn7ScedXsD7vEy4Jk95yX15QJKZawgs6T7PURg1FeLs4
MNArbkoL38GzMqiP4Reswg0zSC7N5A+TH/x2SeQkU6BKOJZ9u6KV9On2aOrXzTi8
175oJgiLqwcsk3sbmToQ8q3OiVwrizrfRdP3FCyU4O4uWYOzz3sBROTbErgEt+Oe
hQbasq9vzNUu+suY+IpMWJvEa02qxsWaLXyhK6GE10+f8QvBLsneaPEilSS2AdJh
tDHx+ULfVmpLFgQ3kQmVRAPGi8M7lQOUeKtLHGj0OecCe6Waudi4eyuyFkwtMVMU
e8qguKCWNxjHXrxfLkRZa00UAFMIbz+p8gAZtvLE8r/gBrSCB0zDzaBOAemove8U
mzJwZedaMEMUBCgfIkZFOzx6h1b42VTokhgTRerDrN8h8RVRzPAU/jcTQsCFt8Yu
Kg8I5QWVkWQCjVc7qAC5ev6LPj9opfGphqi7B9pDKD0rokjh05mAjzga7BivtLl8
rxCSuJvfWYkRcOH9yTVjtDEdHAxGWa6V42e4JhZu3/3wV9+VjS4Mo4qp3POgg6gO
Ir35ObFsbKyTs+EgMll032Ru5oC+BakKao0Era9oyyaAP474QqUoLZ1UgM5rSVjZ
0Sv4FoLKtqYQ7rMKE+iM8Ky/bum95ft6ev6khWPnkScJIt4nohHczzBlpE2r+dI7
5uJUlOqTO5Lj5Yj1i4I8Lxiy631MiK5bkQz9wHfy/jlyRbWeVLc6i3mNvyFtXdNf
PGNvmF3JcgRASfTwTArBCaQWKeeJuCup8np+vzDjCFNNOQj/XydwbRa55vqAY22D
wb3X13SPQbtkOdYIGDMvKPCGRY439jdh7caWZKu0enaTI8gulccF/C9M/+RLGC8Z
C2zI3xu67hBInkAXKPFMJjggg3m1iZy38RTlyfhvwzb/C5pQxHPoLbGYOV9YAc2B
lcC0ALewrd9ZmG2YR4L1AnmRrifX1FD54RyX5TaLXCdNFjpUsSXw+49YYL4uhA2q
kAatVy3kbi26Q9i76hp9hpBG1KVFv5bqw3hKCbHsMUv+VPn2yhWZpkWo3ZMiwR1t
q/7q5jC8ekohrsixy3i768YeU2O/3vgKsdkqFnImnNkWP5wTmsmieGrxrU138P20
MlaUIpv4/HqUDq5eK5gGr9HsPg8fF3Sdww40cmc7QoyO77U1VSy9lt5vKSqU2s5V
/fikbDEdcgao0DkxD9jsWAEZ2WKp+M4Qt81nKGtmrd+uiFdTwpAN1nlGDzOVaDFN
30nH4/73iqYbcEg67Q7Vd/RB1lmQBoDVn4Uxe4gR4LBfqKIPNryohcsGESQN5a1l
LBHzXf2Ok73Zhcc5OLBpv7klDcp7y5gLlPh1xqeIUw/Tv4WWvnN22Re6VylyZXnA
Pcmo3rwwSNH6wqnuQRNb6wITzJ4HvCgYjGXubiyPicn9KHzC7OSzGgeC7+eze2AE
8JCyEGCaJTX+WWstYFtUH9Myqi0OJP99YwprYJdnbyneV0gtSV/XCCLvou5FwCds
0BKVhNID3GgFk7NBtakESu+dBmD6OcmucxrJL6zDXescOFKvT6B0KLes//MsFJov
pj9n03kD6qGJneeIsHR48vDML21LdiMxMCI01/yiCsUDcQVMJXYa+P9L20QW0UPY
jUUvM+rv94e/EcaAwcJUw7RO49znZu8VNZQVUT5r6FKimjzbSV/1PaPKDSwpb07Z
BHF5tl020NnQrd/+yog0x2VQc4msBsXe5n231lGtcRjNowKmhWrYhAp2ZdPEBJCu
OSgYHnAfFQEgRBDKbE6/uom0IeqMG1rBmcF6szaVcty3GLPWrysW50L0Thb2n07Z
eqRAEvt/X7IxuCLXinjBi8owZk7v1HAhRhSE2PsljhyvnFRq36ej+LyZU3+f/xPS
JtdbMQXZzRD4L6IwxuY3UDmB9w5gdSMrrmBBuCg5PKRDQpUiCZ+nH0C9iZ89pxev
2r4wnoY0obG3vqktiVnhlxiR9Z0WGlyQV3TBePIDGSVz7gudZqHlkK5Z0A4CTF7Q
3JDsRuFrbYYU8JEGyzgH8pz76gTrcpruwiOfpBLJvakKTtm24WxO0pE1PHwRXXvR
l70Mz2IoaulD+LlMhgtVUbfJw/IhPOuOYx2j1GSdv8rt8zkH4dhPFO4ldPd1ph1K
vW0zIj7kHMxWnZCfph+BwA8ucsaQnPE72YKcMZ12MtslOOXYD7BvGKoyAlU8Vll8
1gbv6cD7Bes0XxK/VN3blN1Mr9NcTiGaRMtiaJyNNpXMAv+F02WPrxoY3SVumFGK
RcodsJtPbmfNvA9nVz8VcnDwaWwjRfxzPSUcn7lSZkXhh4usrvJ4Fah5e4h2eAyB
f2KHPWcViYMG0qycoD909W2XCE/7e3+RPU84zT+zocTOmuEkxnFynDTkGxDCZEDU
iKPoYWMbhZuaimeuZy21waKjIOgBrk+CkOjlmFbzs2vRP8VDEnK5Btw74EP01dUg
zT9GpbtsIbov1MpGY3t2RV56rYeNcSFBE3fZi8kBWz1Y09qnOTY021li6jRqIYqG
PJVF3NMmkc1p9yrx/XzaO8YGQiCyki/e51UgJNpHyaL35UEfi7Z6GrjjSakXWhmv
0qA4guCSzbH3IlWnBzFNJQlI0In5XOQeBCK0DDZzZCJxlR+UGnniYsf7lMc3M5w5
6J6RTCp8TXGAZulHQ4Cc3r1s5PWZG0Xb0OHONA4KZvhg1VkMsgpmQhreXY5K47i7
g7OOvYKcvRdaaKh6wJCiikKi5kko8CKM40BJaywPUv/ILdSnbFLbK7lW/gZRAs6V
xJtVL+/R4UaZ+diHm0DaJRsz4szzmaN5/eRp64ckOv9IoKKVPhcJKj5c9/QVs1a3
438yiWrf/ry8vvkCEuT66ekbLbIP9XPO5Bhld+7qYX234ap6ngvhJSz2RrQ78uUB
g1ZzaonKf65Q2p/roCjufwDtn30NeKphJda/o5MoWk5NVSNW3O2qdr80M3utQ261
WWlGhRoYqPxa0gHR5bNLiL1jO1OeS1OvAhdJXI1Uf54NObjsX985ZFN81eoEpnTI
JqC6+/3z5l3lx0sGBkTNBMkb5YEnadX71TsiQzpBasVPL1vMJjyYvKA4lmSpJEC5
uZ7ivY7fdcAhsgYCEwOXTlm5l/XRJRSGEsLIT4l4YSJ+735J4AeJwxatXJPRkEZ/
cf2CvVtfwcGDxqj68pv29euGu0cCfMLl82Rc/Gr5i6HqYBRXgdVRWk5iUB5Clfhy
ga5pEZAXPH+bK7dMxc/p/HgnxCpxTd8SkTdnz6LX3ULXlvebUdQBXjUVUa9DGnFu
EYaLFDpkGBp9GjV8JrYlRbdPAQr71blTfBhABON/ENQEj2qsxA1NCYxmZW6owZM9
+IayL1sf7bK/KlV6swcUOVr/LPy7IRjy0PKqCZ3NP+vzt6/7m8j+LE7iIyrzElSz
obfcYv0QRlEzikNXAVlOPBcVtBARHMlKv9lxhLOUjirI5kCKr/fjnJMHrotws9a0
SZAQQfV0O0gkRx87kezl9IHjmbwqmUvMutJEWpclfAJOMKAYjfmLttLm8zh3DUXG
O6vUpYzwMSZAhVOcDkEjzJ36c8RPUsyEREAcAhGRYFBbtUH9wRNIAvBU3QPGR4sL
NoRzMO/cB2B9KOMEY9H4t4lqtknmfGwdlFjvuP6un4y/JtCJ6rNIBAdISSpCPWPd
xD2cGwMFsK0pFcirUJU7H2s9f1DkUdufr66NbPMpiJcDwqr1Jqz9tckXbIW2+1R9
xcE4cp0oG+mn0rhnotjlb05hCNv9XsZC5JvRyOCMlNzt0dxUgQi4iizGvXustzQ4
nEI3TPsLCXnU6WB9l0F3qtNdLtm/Q1EYeke9ZwX6Db12S9oVbo8fhRmQNOrpWSh7
pNpMnj7b0bSQG4qNM0BE0Y7uo0/B7bysEJBhG7NK0dBwTOa+ed3QlvLd4JLhHoo8
bWAe55o9w3vgSCEaL/ES9PJArTKQn16VchoNiW+7fIJ8+CEK4aEilhMCcA7Vsmmn
FYvBcjKqgkWhncqAHNm5PjTOlag9eUpP40TDkHHVYWbz19bUkmCKYzjuL/3j4Zlg
ktHmWWJbqr+Ypc7c/Y/lGWEQGakFlBC4TiJ/tdZXRx0VqLtiD51GW2+7SVZWH47K
oNY0ebm/9oYQR+Ab2VQDvzLg8VfBGTgUujxfWpcjIsrtqhNyYyxLLjfyca63HFkm
lgRCat2oYc+sSyVKpz2VXtu4T7k+bPhVpgH/F/GWPj8SfTOnsMDLsYZZWpoio1p9
0YQewdRgL6TskZIzXfr0BX5UxAo+LWh+nCbzBCP0qLAp/mSrEZOSNGzvzet9VXMC
3ELZkMaUvfvoy7+1G+LFqIuHm18XjKwXIJUeRF+J3fXzfCaoyZPVA3OEpMWfvFqG
v66HbcYdhAO7p3ovuZy/5iMXjdswX1HaqWthcuE+eoBJKAWPMROarf7E1XwPIR4a
0MWwgYq5pImuF7D5HPYViRotcGsBU+z7pD5oNgb1VmRHcgvWZh4Aw/pU1Uf6kk8z
88vtTMdhQoEtoYc/SxAfcC461H32C6e49lZ7ruEcQHdYEYi4WKVuxnynClolImxv
jDYFTYRLrvL+wyc7gSwZToxRjObXK3EgJXbe0DJqmiqY9icxohGsSkx0xU3Lmxty
CCUGCuWO4cQRuuABLtPCOqQLaHI1VcRo5oePjzbu6q/RFnn45ULov3AXWoR3j5gI
RBhbIwJOPueU3rGBSFUnrQyIq3okq5oZVMy6fVnsboA2iPdCwCyU5wRe55Y6JAXW
17ERTRh5cGV1glyPLZnsjohH/Gp6wxB+NWB6KZRtyBWL0aZPwsSZtc+Bd+zfoaxB
7qwPhg6+fmWzsrd1bEyvjFkwlb3nJVYSNkHftUqB0dfW9ZUkvwlQIF31ulNQFWJX
wyCLeRLxxXW37d5gLuqp6dOS9yhZqqIcHz2nfM1o4qjJkrB59EFR6uhH9sk0AYvq
CSG6f5Xb3LAOeRQlcLh3mYkYm857Rv4ooWgzIrgNWavJQQFhKlihtPqzYAhhvOH7
Wj3muMwDsLswLxqsp8pYndZiEULj8VrEZyTY46GkhF1HvxvqzOmqLxipXt+MN+EY
ADNkVODmiAWbLXTjbuFP8el58NVYR/od2dNl0xcb259S5wOhXKJlO6NBTfKjFK9A
UqQc0/JhF6ZK6ogSjY6URkIoLaXz3+9KiUpYDNxgQ6gClJ7rmcTw5gNAUu2dRZVY
6GPp5ZN4AHsuQxiIbExdl2uJCFYuNi0fNSzK+iVvsh6z4ggihwSRfZ03b94LCqx+
IBXL6SWoRqlnsgQJdyN6sxnS/Epja4V+flkB9wT0aJk+SjrSfw4x3ncSmzYU83G6
5171KXBmO1fBxAOxGYQ7I/ka9HGn1JEBMHM1qBMhv7rdwI5LpHS+E8Mfgs+bmdW5
PEJWT8YNuPlyfkguXubRq75snEAynHNj2TLDMPXB9RI6G7U4qG+VaQHFRah2u3Eg
K+b601fNErIPzLRGwjkc8ZnZW5gq6Y4odjz4q1BadllKCPL5oN2I1+WFHsV5Z/3i
/zsefv//HyVhC2xX2MwiZOrf5uXFnkw1vpfeX0BtD4cSeoEskT33pkaihjIBwbZd
pFu4ZoGymt9BFPa9u0elsCm8N+oAZtFbaQJ6TlXOzBQGd8ql7cH2Hx0Oaq3k1N12
H7kHn6cLkXgx7R7RarznjoqjtiNtwzv8WT7IbKhGiAI1DSX33DOfoaTRTGQeasp4
gi+x27m/nFAl3YmJcY5y3n375LAOnc0Qy7HyLSMFQ/xrzw+8iOdfIQFYrEuQF1cQ
zlSniezieREyeKH+TLrwojVxBWybK9z2rPrIswYqyblbu80PEaGzC6/Jpl0aPa0D
UkjlRk8Q0bdFh5F0RZQ+9DBMsA1GFWx3EEoaxI8vn/8WptcJc0Fc8NWzSWecarPH
29QX6dovO/Gi0j9lynkzTN5BJprRo5ukMMEScHwM5suf8ge9VNTUDPgEgDZoK9Do
Wyg6vqXExHSzSZrtWpWVkJpdgFsBL7DDSlfanK11uAB+gRD1dhuSK7nvCgibzwmg
l2OZXXrN6frmTtrXAwomBQAPX/1E4FCv7QyjvNqZ5+BMc55I4BiJgCSqCiS7BybF
+Tj8BUDi6gSmknB4q4iunHm5Cqssy10k08bsNLp+QIzjb1Qopi060u3lMguoacNu
opVD1+FNGyY6C+EKr+40cHbNcls8QcOzbC2suSrTg30IwgpODl7c+V2J/5hkfCUH
dd5NY0h6jmq/A9RPcWDSecO3xhyYeYYRrDuVnBAK40XUy2VdgUxvSib9lCGa5mtH
IP7txg5AUjSBFkgPzUs71irj/qFJTO2GVyR7ulJKB/cAZd5+b3qjnZa/mg6czHhV
BtKc4MYnD136gyvFXIyPFyiDevBXJzv1rj2l04606zK+8hVc6uE/SewwqPIPanyo
YHaMsLKA+R9J8EcWiJRbByqw+rzoVjApzfLEydqO5MQZSTX6YzTxW0iPgIa4LjZQ
RokrYmZxz9vko7NYBDU7yPef/ag9AY6r1Ca01zA616hgaRMatCDXPLWeBKUEs5f6
dv8mLLuIMbgxEiTKJU0Za+HQtx6zsa72NRBp9hoo2Nbur3oX82PvdbzeqMBSajtx
ojGpi/Lk375oYWlVGUcPTztIj/ut6MV9h6VoBPrubKdLMraqSODdkDDN1fkOOxMH
MuAAXzwzS0/tYbdNGmDEtSJ9En/L9RpnqRAeHbFHcMCVOThjLIYE4kWDdvnkUBkA
uGuseTytRIlWu07wKD1E1D74EgYqFkQOt8dFHkdvcG1H+co8TD+xXiWvg+DeY+F1
lI5Vtn/FUhNtAflImwfFSHCPQ7U6Gpyj0cubgN0EoJZXX86owhPjk9fjgVYR8/wL
XVRlfF4NFeDtWCahWtnyCccR8PFleGglC+yg1Zs6asS9zhnOR3FTDyr5FdzxXJ43
vKKFR8fBa2vC9PgTFnyeOTOyUqzLtcQZwJCcqY+MJffc2G9tp04yXVAcdHBhxCg/
0PJEO8F813r+dVDBp9BAfTUGnUoCBXLrzBWInaMWS7AIWgxI5pZK53E7OdoGqpqT
spK64keMM9HykiQ78V27Hq4BNh4XpYWzaXWPCShEkHgf3JF7CTioxIq+BAufqVlc
0aa74Bj51785HwAun4jrcRoORyb9MPFJR4zA8/6qrJcNNSHszDZmdD2ha+Nc9iIB
vT0y+rr4D1bYKCRcdCl/aLV2mztpVneUSATnlapdT/Aqd2ccsDWu2Fl6t9DaOmlP
Uu0thrKa2CSoFf2on1P9wkIxwM/LpBv1GI0UJTIgjkblPzGa2UFWgVtdsIO9U5B4
Hfutj3ISwdDoGsNY/yxB0rRpHOnT1fDaJ1VniAcxwLoaCPjppFZv28hh0nc6ShSw
KueARR19QLm1facl7QT9FJJPE2CQg5Svm7Sgf+kKk3ApgKgkw/5EmOAvPgsSaLTa
0ykZFe1uxoUo0eQob5lVBPUTXigxRoU7COTnYXsyynRBZMJ7JyXz719GA3xDKJnQ
Hjb6h+K21iKJkM10+7fkqL+cY0cOx2OzbczAFzlEyxnbtJi1tLpQWTV7PZWq6Q1T
r8in30gtYn5+BYIUBGEMcjbVCUVHGYn4mGn2m0YQN+7lsSKvBbHMd9ZS1Pi9PtFG
z184Sbs4QekgEJ7fwzJLkE7HVgGybU8CX1SMurDAfutj3sBxO3y+JS/2fc119Tya
RgpO6jD0M7DtDIbMt7TB+ceH+1UqPM4FfVdfMy3ubBpLrxOo9D4V+XNe8ZT/tu+H
3lC++m7ujJs7WyZRsYNYYIVHZPIlS4cM5XurY4gV20ZU5F4zyJRx/zY0nVrUONyB
YvyD7z/wJvojSpts58xpnT0yL8BkwO709x4DjF2V8yArIofpbfghu/ibC5RnYE4E
KmpLE5Jx9x+vImUiF+vnrknmiIyBN7Vo1E2W2gEJf6ftgA+QEHQfYz23CB34yo91
x/SaNi8AFKgbbpGuU56JnI+gIPBtb2zvY1T1jHY/CaqEgLoplC9eEHwnPgRcLpdP
cjaqnPtbv6J98gHzPCgXPvfSzMUmoGevgl6CC5cciGkcB+zgM6JpfBU468c1rAYP
zkfu6DftQ40ejbXMSch0LoWqIaYxIC+GueH7fgQ72Q8XG2Lp9aVbvCbN6yDWMF42
/+cJiLFXLnkId1Fip8mtvno1SlCLgqxAWpz6kP1eoXD+Mr+D6kLl2WbqY7gRlxtc
vvgwptcqy8N0utJ76Tpc8YorleSyhbwsiVvihupUX+rVyy3oRHe8AXptE4eQOF4V
9DCPiUCh4v6VSdx95t9bNA/rgnmMbYUsUPKZJwZXThGbUgDXMYAGEFq+nbrO7Etg
/sR30Go2buIT/cHpMcaaqUL8pXGQoy0RpPPqb4/06fBZe2LcUnm+79ganeRUohs2
Cfg0xlR/WKp7y0BLSZMsA+/MggODjHMtqgG6X6Uil+iNN5PF44mQVJpUnrK4dwB3
Q4kygWZZ+GejlKcuRtxoIFLjrFYI0iumR1axizRy9G0CxeU2qpU+Bx6UyaMYljRy
ilMSFgJATM8/B3zxP7QqO6bcmcfx/STOsmL9insh3HU/S9fh7cVkfLMQS9fdc7EY
3/SXG7hdiQB2Mgh6/Wtj9HOFBmskIkwHGxJypm+4mQ8jGla7fkjCAIhW93wcFXdS
/LXU3mjgrfcGFVCFQCFwbQxAuU0mMGUYw3lv7boZGVAwoG7r3kgm9R4CB3oj/Fe6
xXXBcMwsUCM91TCT5hspyqWODmyTFHDfhiYwFdPGW9diZbw3ObDni+YByjC0JXxW
2yTqxpAXTB6ev7tP40G8qZapyIQJOFhrJgl2j+HcwapJ+jc12JZYWKJdexcFtX+Y
QB6HMB8UBfci/mzz4wqhYlOisAU+cLC9QmXKuzFZpmsRDXZfxGJVJsYfF5xBp5EA
UvrnFE+slvabz63YDPpqmZOnb1tYPCqU9MeT/mG29pn52ZI5NuhqwGSzXRRsyteB
W4Uul37tTDfqQ6fj75llcSlS04aTRVtGIVC4HSx5PUEPUqV0vFuYvPrKwy2pjmTs
6f4ocpqmmfU2CG/6qf2WXlDIwwICtEwvMKSdNW4IirAk+YVIqYyA0YvLs1g0KKEE
v7c/uAFxSYveERQHxBDS9p4XBxwG+4rUmdlf/dhskO8SS+jHGrsEhb6FEqtpOTzf
HQbrzW6aNLBOmmS++vF7bMIlIQeIL5KdOhqJqUH1PXK7+a22HXlvzM5FAtQau5ec
eWZ4gaU3uF1lJb6C+qpEQhAT5XPhJGOVWT+6It3NU2YjGHd7xQzeb9UCHZTGIByi
BOqJhAl15bZA+4LdoFGIOlTPt2pn0h7etNs8RWi+GPTzikBhPaGhRqeSw4gkAS5v
p23i1jDHwhBZQ2SB4akjiQF3ytg7cM7eKA06qnCbLbVVSs96gL0RKs2jJhph/ycQ
GPESF+ZBDrt0phE8V+DEXdcs/65TCIolz9ACHE1ErK/of3PYiIwZVt2JUUBBwYAf
ZmkErg4nV+p8wBtROhMgruidzhtddn6ZFI8PhmulL2CwhEO1bXZj7pfxa4cxFprJ
EHpxsI8DQw0Bp8CWZmMsKIQ92Yy6t0EB3Dqo13NOZKMSR0raX9zYvL45wMO/clzf
VQW7nsG2vjdd8DeVYRGyKRMH0v5lJx3PHMUurBImoReD+8T0HiN3Pg2gtY0r5KGa
HEL0uTa8HDxWkJSugv8lZTVA/vIUjCLnBt/2k4WrkhDhGeHQGcUGmofjiGzi/83y
iEjlSBRGOpzCUAKLVpWnBc7OEVhCYM5iql7ljSotONXW31hkrNc1STv7gWSd9gHP
aXR2+PNB7VS1FjhuJOYKQvxDYCfgnml7GzI5Uo2txtk8GSWjko9mWrZlQwX00zca
f2H4Ubrg5Qi7CDa4XGKCOIlPI5mZ+nzHDGJ6BIp/bVwvQTMvbCLgz9AEf5D4m5xw
38OICBt9AQu/rGfZPfdipShJcTwem2cQVv4CpHtv0fjO5e8rdyWB5SomgIi0mtI+
uedUXuN9jgkDpTNXrW1SUEO0D4VGLywCPuIOtddJe140za0uzGQp+RtYt0+w/VDS
qq7tWtvcCKGAPWtUM54p6eiUNv16wyuEMfQ1ndfuJVMDdin0mY3j5qivWyytNf/H
FQOhvh2YCDpqg68CZ27dlNyEb/ZNQn5PKu33EgHTejdPFDTMsbIWCxRMcmtwnGep
TIt9kWVaSzco/vG3szh0sjvr7pPfGwGqdOIaSTvkInFeSTwDee/Y6//nKUFSTLYv
QqgEoJqYtHrB8YgELpBGPtjSaHtIqggRJ28ZP6EQ+J7XMpwvY9PgrUW2VnuzfOqT
cgJG7yv1WaU4hijvMyB+T4LBaBHsqRseWEY4G3Br6mRf4+pu9fsZf3ylltTggLuf
nXr/Tncu3hEM0arvdLh+nqDl6c/rMqjG49nUpRFvlqMUYupw9Fjj95N/FcfT9f2+
/V5jj1rcMqT+53LTHQojhkLUg8RKzlVyb76aEkx1O/frQJp7YUbEWEORCBAEJWNE
M29l+ontk/bv6WUWyKSBXwqrYxKK6vETqRwzwNIwNYWFW+IgGrzoWudpiYvoaZrZ
Ma8WEw2hdmAK0G/VYN2VcQf239kWuQFAJonnWgDa0JWnghC2gqrObRw09Qvp4mcX
pJSjKzmEslR7JfyxcYRz1yyC1/UgJWciCiqFGEXghvvU33G2QEVhxmWNStAwpJhT
YZ1fo8nhmsdm0PvZhEmqW/+t8wYofoeGoIQs612RZTu5D5t56el1yET83PypYuZh
vvFuvscWroi4NajIneDDN8890h6ymDgakIyOrlVdxoDq57/GVZjd22Nl8v0LHGfc
TgdpxZtiubvwcg5NlBacpvfKYgdfluXCx+DWkvgqJfufL81cxRc4czwM7ebbr4GP
SMC2LaMriu4taSpmF486bUcUGTu23jAszchZt1M5spwqCH+wJMN1yjsi1vfswupG
KkQQmVUEy2Bwp2UAtZYbwf9RLVZoMrrj+CKaS9SMHOFoLTKJWOKJ19ZVIhtoY9wP
h8upcGyu4NrqlX2iFuNI1rAFZIE8NJeCq5Batdkf3y5wfkXLPYS22+Gd6E5VFDma
dLkU5lFgoTRd+9m/yrcJaPQLAq6zpmvgNegls35qegSWNu36s4b3IP34Nn1rCoNT
ChctS8TFG0vjYMrrmwuHX1GTAmG3djDZ4K1Qol+2LVoqkVDl8ysZTP1UXVk9/qJ9
aUtVQQznH96sJCPYoNKBnACLUEdkAD6ECvmoBDXM3ga9FtPoOjJeV9JjwkhnFwIq
vcQoZsEkOtpecll0eE9yUUslxDEQecIZD9fOMV4Y9jwRPcNgoo5D0a+i9PCEpAwp
opfBALcoUsGVqgBuRcjR5o/2hmowQNjat6aZ7TDWyresFThdnV6W81OAv9aXYfBa
YNkn2FTSXuAiyGvpAESuBsfFK4Vj8l8ThfpjEq7pNBswMWtWqPb5SJI58cAvxQNT
vBKIl0MmL9aDkn6mHrHq7zOlbqrJ68pGVhZne8AIKqzoXl12LreSGL2zuL4zuJw5
d9mZWfJHIp3253Ad23NdAycp9kgvze3swyy3jdHcUIKbJrbIRIcshh5g8S+b8Ge7
T41NoCfZM6CCZkjyobWSIDgNYcJkDXJ8iUHIdI687ykeblvOQjmkwBgnwwlOrYp6
znoB8xzVRsmoElY5iy+SYEV533180n56EtA9MXNZd8d7njuQt6mugMDQgZbXhP2f
olCBpnBb8D3Jn05B6gyvYmM3/AM3/Mc6ad4Z1z6OlgauScIgYzK6/IHuQ1DAiGV8
/dqzm89umOyV6ioE7dPwanSzlf0r8dqsDLzYtQl5i15Ap/hHPHFWNtDIS3fcbdSv
KgBb+giBMCWDNtR6zKcjehzZeAPJYc+aZAACN4RR+WARHKfr1eIAnPuQt8vqfNYV
n9T8pI2mMS86aag0zPE8Lg7Kr/9xLM4T2xzEdXpBRBqN2+DDrNC1rwFD/ZRaU59r
1Lxg8extSR0saSgLoXsKKCGX+srYr12wgvJR+sqfCrJT3TNFVGpuvkKB7pg89UBX
XUAhOClIgyZ/+T45ac8vPi9HcTtNopIuf+7HJc1Ir3Ega+wNXd+prZKLypxFu6OG
Bhighcq2UppGV8V8/wVwgcL2cgAGO7PjqsrZz9FlqC0Swnx2OIbTIg2eujGTRSNP
p4vEptJFJ1Jl3qtB3GoDc4j5YkNx0Wx3G8+MlvdM2iLkH95mwkp30S7S6W/6fEKP
hz+kOeEMP57VtEJsHDWMzgL77PSgpuSTgMG1DkqmXJfTQ7eQJNEw/o8WMU1hK1bu
X26K6eJ76duMl10JEP00zjhISYe2OG+zAtg6AZXm7zWcD2pn7IfFax57JKeW/QEc
WE9SfHJXnfYaiiZC/OWqU92HtJnj6y+1nGscJNybfMw6w+g8oCv85kDDUCpn47Zy
4H3XXkHQmJPO5uIjEJ9u21K85j8Rhy1WMn5USk7aamu19VX5MytBwUxqhZwhn7hM
XWNbMwQ2TXl+7HUdnBavwhxX7zG+GVsKU37LEIO4YCV4iSrazw/RmcBD+rjUPVvQ
AiNxNPglUOR76FHnpiUr4c7XMNQUtashTnK4PhUIUwdD1e4+W/pi1n9Nzkbe7fc1
bf+dWqomW/J1myV2FjNHF4kVN9BSHY8GCZ4mnX2QcR+DeunV0vk1ZJ6O+qi9Qv0a
UTh88jZgYsmpe+VBat6GT4uyWwRt0HEOrQlFynER0AXO3tIMEOXWkYSrBW2sEB3Q
rWEphkCEJX8+7bc1b5XVP696QXROgttLT3p3u2biq19ihkKufWAiMtOH0GxA+ISk
Z2GpiSKkpZA/AC75cjpa3fU3E7Xvkd8ZLWN9mATnG3yKoC9XWTah1BgBvqo25YIB
lwIgocaQ9wZEMevUCySoqEMqQq2ooaveQb7tINOMyXLMVR0xxrGHoOCIQ0m7EKuc
6cl/m3ndyvCDDPIcRb25J/U63WcX0rRBc3cxJu/XfKtjEkBBRG8sezX1lg9aX/k9
XdE/96xAyaIA4WA3RHBzJ8u4NehmTU9kRDkFUjoFersEFYV3pvGV+JE7Ioa4Iu+o
zuf0EkbLo0p5NzRHil+uX+tUayULA7yJ7rZL+o0yctihmTCxbpjIP/zaQjafVk6K
cu6hZGRdJigUtG6zv9UfOD4gIANb22vTVKjjoCNngjw6xG8tYwOEWKN/j6Yvt7TQ
jMTknTTjObct1BCiPXHkoHoixJHKM5tOzESNa9uufTTeIZ90qbGkhWPgIzzq5nrk
yPe+QQCRcngLxQPZPXhuggiBJxkbSYujb6TiIdmYkPrkr9QZ5v5FiEOSKK8B3LQN
Lpj2R3n8/PtWi+CyXI+ok7ySo+75MepbImxszf0JDiY335qLsyPIGj+XPcDRCXCL
bDobZunA0ltd0M05RVA15ElUOxT7KfD0N+s9wgN0zZogSql1tOchtv9lWdDaCnCY
/J0hicIgUyRpfL/uHvVM9BkaVwfgqkb66MS7WBzL5pSoA2grtXrYuPg1frz95xd2
NcrCdCvMMTohjVh4lp+6TNd4HDmmGTuNBxymXQ7hlLPHK57qH7FbKxdyVfhAjeMz
5g4DrhKpFFAo1GIHPWuyXwyaVfANteDCY834NE0Tu/IojztNRc+MXVBirKI/aLu5
Bri9glovn8k1CtImp+TiVQLPgkKVrnAj0WEpl6qZlHTizg/gyp/76l2G5scDgETK
HqrcbvNfgerNBMV69FqIQdC039eibN2W+46jqXy9mHbIS05+HXQWOW7nX5/ZOfpH
1/If/kUF1w3V6EP8A7IyuiIbZDYVk2Ksg6fn0J5kob49BOx1N+IsKpaQhOmDymkV
oLLKD4yd9yxTaONdV8om5Zfuw7C6bCmKZ7e3ZkwflWmnyWlGeHKxdEhlrdW0BPly
COcTA/MbeOaXIjLeHxaxs2kjdAfhP7shwOjgFUnTx+tQY1gqxs84bRIqGZv9QgSt
BBFR/3n3pk6zHchce5nCYk6CGfA9y2vBapWazHE2uTOSMywnksfEMOxVXtXxWYD/
qRX770NLTBhxtmoQifHTwEo5ixTrz8xkh6imzAbeO8KsQRnMtoTxxZxev7e8a57D
hYu92AvFkEqaja/X+0WCRF3uSxTlHG36blmrGDkiLaclj+sRu46aShqG2ZHysYXr
/PFY4iNWdT0OqDEbQN3zZmNsXPwNGkuGLUD4DrIRXFx9pnWOgGdhPefUn8VnJwM1
gtENJr/KbdaLaZ8y6kkTUUc9g3B/YCI1Jys0aAxvg/QK0f0tTYM8tWr4wGNn2wdS
LloPZjjk0kyGiPmgPZYI69l5q582f4v0Gj1ocmXBzW4pRyIMLdmw/OVvjvkQV4kd
NyPXJ09Yz8UxGoy5GtxkaucJpYLwlICGSsHGBFib+lfcq8OGbxuiGxcP8rDMQA6S
7mGaccuRlH0hecuNN++NvNfPuyuR4oBt9KjW22PDYJfAfffX7OoaGETEUMmmTp21
ivmL6DhhFxghQrLTJnMEF2F6hGmkZuzpoX0dgi9sE2LUcvZeLVp566fKN97yH2/4
8FGPoa2MqRncULD/EuT3oyAjHFJePDcMnbjl7kJUK4MgWelXPPbwjNP797iFnkFD
veHYMcyo02OE3iXfyEAqZ82LtHThi4STPTm9C9wiA8ouRIpyyUI2kfipe8YT1Ko5
cdNF0/AnCyukOJw1fQgtRB7i71oZYBQf679YWZn2zmosDufHdSr05fb9KTCNoLwb
0l6D/DNoCwRruSUpNzGhu8uOyzmJCdWdn9tgD3JmkIkKPiIN2wT4VLtCfsuZWu8D
VjXhcXnRMy40cvBqtHrA7CQ6D6cZVu2hPLJWw4+yIsQpp0GCeyvho8xnRDqChpE6
BboFByTG7vD7cTptquEr22WDTgWHyvbg7/WZxQHu2JFmQ1KmOSysEGOO6a6Dw+zX
VIjDkHUJcsfi5Cr1sRXRaMaTlq/7uBjwq0ZnlN2qdhXRxO5bKKeBRYNFg1Gz6vQp
mBtKfN3GHOTKX/R/ReGEOX0rjnYWoqyYqPEXOsQu3Hziptet7v7H3M1YXfQP8YfB
6NuyDNP8eSTiXn+BTTSuD9uUXq1m2d+sMJIkW+SThk3k9G8kbvKw7xdUQp4cy46d
CKKhqZnzKeTCaMK4eHi6yeBJ6/XOdcbj4F6pxotJcgj7yNWIe23zoQJ5jzQxVQL7
afTZBmZfQKHdV+dU3rippbKAUAfvwN5HNtNBRL/MX0xSFIFQCZ5uzDNXWKHmjCR2
ED6q6oV5U6axXkzL8IuxKoilU21xHSyB0/dFkCCjaHvFyVQX/LVFZVL6+ZbRtbhZ
LNS9HcSEIfOTsZcAmOqA/SEburfU09WXZRjzBDeh9JAsQV/nfmG03fSR28aRYYgJ
jJDBJzxBwweig8zxFtJtRRvjKpCs6VFwsVqsRjsQwTMKV11lDzo0UoXmnsAxSiDy
wmOFiDwjhdqbdbqOZf4X68lAYLhGDLtnQqfrBm2jFKZYCb57aOTfeTo78eMuX5De
w6g3gVGaQ8EwuHRMGahhNMrP7zxc7067LWdjBTIGU5OSUFDqcM1xYUi3XHNct/Ym
ggaXfyt08sJIyYaxI+XOvvPQGQRbQhsMzvQKLRF0+d54zqPcK0xDrUreuq+hH92h
bRhTcsnmPktU7vkwcAooeqWWtmy6bVYnDAEo5wG69+4H173a9aOzG8JoyippRByl
HKUyr/iP/gywjQlDHtnn2RbhcPN9hpFwNV0i0l9jVBucCvhg0OHePbxOKZ5rrjuV
4faP4G2q76RPOAGXoLMWYwJ3XxDq0NBEACccR7rsRWH3KY59qs9Wwk1H/mr0HYeD
DfAOWFDEqhVfSO+NRZlLmHquSALS2X5IvGlsFmOP+3S7RSjAPwWQAlTU+oK/hy6f
PgbwHqa1gE/vd2LUHBNsaZfUNB6n///CB2CezpB2XSDGvrDfDvJ9CPbPNJYkmkLb
FV+bHOHVvSE9603ZsUIdD/Mh4c1yOCch2fsION4LJzG2j3ZibM0bJzek3vy1Q/bs
S40tWJwl/GvJcyRi2COMeqH4a3ZdwVEhyloPO1F/zn1iDk2GXIImFTCacwjIcMLH
7MysoMgvOBOVN9jKFt2hmFQ6rn3khNs5Rp2rkKk/yvaKEcALCzAug1xUpR93yZ5R
voosbtkml/CIQAsZT3dOOlJZj7LPzyBw26Bnc6bOR3Gedahdlw/IW2TCA9LMJFIf
XNxAzvD/2Po47XqCc20kbK2931TAitIcuSUMRoyKU9AKrHKYrQhHpql0ARNntzHU
DrB9N/oz//eoWFD1SIuSzDgbPX5ktmvlED6qgSDzkllc8sStfdkKmZIY2ksS4rHV
gnsZAhw4n9PDSvhFjzD9LEFMGgP+o6SQNYMxU4RkprTQYxI0p47GbVZwnjwSt+1Q
mPgegQ/ioftRUsbIV52TYxz6BlDKRDUzLchv4ZaDcFv8q9ZkDjCk8wSVJUOoqXD6
4ltDqOpR2o887I18la5gCxrRgJFBjLJFZ1P6uweao1iS3MjNwRsGwIIiBZgqNsTA
o+4uSzQJ5Q+RfRF8NFlLnAv/8PqdEjtdsJzDCY78vM+XBmqhVkhEdGd0hRPPvG6B
FHuJMhE26vw33j/57BaJxiDacHZeqib92OlcX57TFpaqsTNOHCNao71uDHN8WdkU
ugiayia/VasqlY7EJJSlNpUzFWj7I3qW5D2pEkn8ZMRCHhKx74pFkLNOP93QnKTK
PoxerLlxXbW1tB8ndOaiPnLss0ZMt+JguT8nplW9qmIOvmgfn6tcAzscmcy4aVsV
BUio0FstKWD3P+eoENiQI/YV6IliUeiu9XBK18RrprAnbLeSqeqh0HpCSyb9OVQG
f+iBDQa+4qm2HkgUBAEXpdK62cbIEq9wTSJko2ApcDrPxPcwHuAaATkjA+M3vkfW
D0axwvjI6vW3RqWib7cd/DeI4CTjfFg5CocUIsszeChUatPsQSppzFoSZH74p3/4
4FCbfvJ+i3elqaU67XwgrBSoUoBKlqKeHFfCNJ0S0ni+pJwv6JiLmmuG1PGJrocH
s+9a80InBxMrIkl/nzDGoO8X3EDJ+KjR8cQME5utpHdpY0Iy/f96DtJ1OySkHIzT
2rJbg2vU8vO1UTKIJUK/T9pcFCVLQVDi7kdtn+G1n0N3CH1Lhh/2JI0Rlm131h3V
BOwPG6KngpqTfHXw/nSbkIsJNVsb7iXy08bSHEvY3K/k8Je5K08wv9cZx4Gr7Olw
zwHb8I/EepE6hsbL2JwKQaAonPGRPpNYtqfBlM7ymv78c7mx5aWJzBXj5uEf27SR
eosP1pMzkNM6xQqg8/w3JCjrVFxd+5oH/nyxBDPaF0oZIZ/YarXmB2EI2IRkuyP5
kU7xFiRUJO4rJ3YdNceaKRhuv4j1eze9yETTUsJ49KMVoodJxCIAotygy0gY8b5X
6LNWvfrzfDa93FTQxWIBFXZHsYPDwKpThq9Fap1QTbLkRsgnr5f/GyyA769PDev9
9hAYRvts4LJWh0Olw+b9iLLDDRwJEx+lCAPtKCMYTtIArVSIGe17vagV0UGNhOEz
yKLl3zCSwhRIdWIhYJ0WcRwLtPn4GY49hpwL4xcLdK9xkZZZpL0psspNpkVa6Kjq
cg2d+gqBH4/ngsjrZAvkuJyRkMGP5lEWvKyuwo2MzkzIl7Hs8rb2avIQsNnx7zII
mkTav9mMxnJt269eKuuhkVG55aslMXmyKatOdYZ2nDpshrWxoj7tlTPEI9dgjl1X
Pjjh9Bac3YgT7xgqdKwEVWVShB8xxdHtuQY3ogb/6Fv40+WNxafRydiYVEU+Pmhb
DlYvK+gT1cJQnBcPJjGKFInWvEZ+/jHlnzKPkOMsUawxBBc1cp3frAkH1I2EalNd
4rOYULGGmdFeSzr69ZRrjrpQtgsFJyMYbFWGY05oFHc3i6b0UcYFqhoKqumrzxW6
HlFT5eQlnuj/M06DBIvuQ1ARC19LmMRO+9/lNfXIEHx53It2OcBAl54HbV0LuLY9
szSAGIQJ9FvozLPVngx1VTKCV5PXZQe+1kDpZyaQkwV1hFlmk4nubALmBGHKHUB7
Qx+cUZEVjAtHEbZW++HdkEwZHMPgXk7BgkjqHsT7fOLKxA3ZXpTDByFq7Xh5expD
PdqA2+JuW03pChfMhWptSmJbj+7H77HBify6GJddrWgFuvs4QLxANJluVMV+3zJI
MIoQRiO8tHd3+8GZcEWAZTzyhey/xQ1h2K325yTgAhs4KQfTx1DGOJ5ssMIFvQcW
da8z1k+zdrlUfc2s4ttRV9BhZmXEiGoJJiniVRwB1f2opCNtxmvgQN404hJ44JiD
gZuXWhommqEu9eNoEWPf/B4Y/0eashO5VIisv9g34G6CoCi2TCHl3NmbV+ePZ0z/
`protect END_PROTECTED
