`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CQnWLPAoVCt++Di7bl+2ohSGhhlmf/ZgwPEeDqtj7kXA6nRjBdjLV74ChUBItzzQ
kjAvAUUwa6MggqcygfOOEaEff113sUIQnkfKGVsUeR7v45kq5VW/sAu/pwCf9mSo
Uot74lVTf8PUcU8uxH4AF1wa6XRv1kWBeoDPkaOx3ER005hsxMIVsZ4HMSgGJKPk
S0HiLQxByKMt/GuB+9bjsKH8url9/kkTpiPimShXC0qhxHUK2rS7ZAKOKF0618LP
+2J3tMIO/8CHN2tc84O098aFfpBA1MAjQblTjvAlZESlcC04ygWKKHMGFxde7JTo
+DE0sQPgh9cOyHkUQEbD+SlanyKeQ+SjzjOg35T89RiWQqaGOv4i+dhGyqp/wWIM
EVaakx2qSlpiM9V6SPP+AMQ09wc9UypM92CiwHdrhBSrqbwbmeEn/UwBU9mD9IDd
tJLEYztszclD617PXSSIbZdGxr8vbGR8jM25Yk1+3fg5DvPYSuDS5g6wodwC9sV1
JMB3YlnWOWdPmt3RBqJGcbo5bbbC37VexHFxY5dSJgHlxVYTsQkKdp+Fl0T1jDwU
Vx4CTS3em6+4od/8arUqb3WB3YZzjxjmkAjw7S/8oc9hviQdBX0xl0+/hjaEHUml
ORCmx7yC/oFm7PG3FKSH3ocHKizzmO4LM99KaQZFwMyNEjleAl24K/2uA0oGLXH+
/WadhEBu/cs5kiUNziGCyg==
`protect END_PROTECTED
