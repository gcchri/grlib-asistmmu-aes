`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wk2u+tlJx7172v+dhQE3We+JpD9/RBZ/37ULTDjY+80CH7EAOZq4y9xNSlXhMNRZ
cZM9w1g0wr9wTBJWmMO8bmiVmVfGvLsm2Ise95kaakZ1ZwaRwN7Qwp9NfeMGRS41
FyxrfTZcodk+M8msKXdg/kUoGlzjb9ZTdkJkHXs7yvDQXP4P2CJQGqLEEpS0Gafr
3H2tvpiR8zriZaoeTBnLIDU6WyRRUyQ8sHIOkyVsLNUAsxfBAM8dE8SUWufiqYUm
bzLtTaOdmZahVsALez//Lp7bAV7m8HtazqxpP4u35tIUZHC4QGMsEdyGZFW3WoIl
`protect END_PROTECTED
