`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SXCOG26xzDRgKNOwjE/UNkIhbfUPt9ZFwt9RNPh7IhzLGM54dI1sppSYabjsoeyU
3wJp1l855cPhRZlWnujsWE17U57/ji5j1n7hfP/IPqpOMZzSw7j3R/fO1XlP/PmI
aAQ0ed1pNgEHDLIHyNXTaCNSMFz6BeTCS73arIX7TjQEJrA7zF/kZFRs8q8bHby6
DLo76h5m/vHzl34ZxhE8mSUJtCoK8COTPXMZaIVcM4i52kyXqU1laEF3gbtrQIzh
tZtzHN3HuHQvx64kVt5l5D9ZliQiB12KBxtx8gi8vy6VJZst8zRjcmTRedISlSAo
0wqko44P8yim3ph+6fImM3SYThSAPONQP6Kjcxt1VBNtk8xK7Zz0JyGEXZO4tI9m
rTQYc27ZD9aq37NptUxKbDiXs8uFvF98mq0YC/z2gIHDOg0piaK/9vgnzlYDkimg
b78rgxbfALTJY95DW90VxNdCa+ezZ7Gfw20IceC1byLoQO+IOw70kyuFkMHuQ7el
gNKve6ohEEMTpj6tGY2St4EupnC5YDl0h7znH6eJ8oZBapcXhaCxMo5BzeMu7g8N
P4eOdtYwx7T0ZIhIBkoDZ5cPNUJ0MSHR3iuwLKjbrSFhMvTHCXm8riUnBnzQBhna
SvWAZcm9YgfBpYYMV7dxqjoyKrS6fUqGMcjJk0JQdZcF44LS2nfDH35W5ROrmNMR
ioqso46mvC4NEg4nO+Dkmg==
`protect END_PROTECTED
