`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L3+TV1dihV+PHmjBCFuw+b5Hlmm4rSO9m4ERHTSqrkLQEvR7J4he/aITZW6k/Z6t
po7nVH6FIuAS9c4psNE+j1vP27vyaZxaZIn1El4Duz8FmOmynWsiWyVo4svCx/gC
EPZQJ5x6Kp7w67XMVhXFAsYnakdSL/ZL3KDF+SKAxcf3oFnIYlOoJ2HSkCOmE7gI
gSeHWpzKR9WUe2vmhAE6byGwQs4hXqkfnHmcwmhhGSr0YG1GWiiskSvgF+MjPqoO
g7TnPcjL2KOwAWiqnRhF9GhfptVWgV4zf0VtpXVtBJHBG0/ndZijXxQxlUkyu7AZ
F2rB5vo+T/yxxaCqtsgnWDERTizCsrhz1GRri36CL+lEw6a/DwMUVAph5MFMVUoi
hksGVg36t6/UcYzV96gDqUdvqcC+3ckqUTFvCjU+ESwnWLAUV6dXFrP4n8Aozr/3
Ek8gbIjVxhpTbpiHXW0S0wX+pLknHVC/kd94xA4tX1ykLTb8pPkDueFnJJjNhqJ0
onQeFjQZddXGBMw0B81HQeNqo5CjCnwbvxgWzhWI7onkJcgvil0vKEdZpjMX7YbW
`protect END_PROTECTED
