`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iqbnOUcIdydw+/WJZaFTl1WHBwK99VtSFXNXVD2vvz6cKVnyKaXYPzci0PelkGkc
VdreJUkd8ibnkZGDTwjCHVofD0EEZAXXPe8yjKiTsrO32fr+FmQlVdaVhyhxgieO
xqMUT0fcGQhEMtuZSTy+tmYsJ5Ijr1gVuowodHZZHi+13pRvUoMelmYAgkmdCX9k
ZJog/9oVRgIebm6aMrh69g4xLjIWND7fYQRWoPITP6mwYdUrIzLMnAD/s6P0o048
pLgTRzQ0oatAxxonwV5sTy4EZr+rz3BKwAZ6s9hILLHKLS0cBAqT8crlMGqTFXZ+
mgrr0ulGpm1jU073wpdGJyQZLBKsNVCDKYUcx2AnEQfFGove8DLiS8jhtoGXq0v0
kkBtJspZISZ7iKsXwUC0973BdvWQAzBxozI53pBNvBoZRV+UAzopMkqbAORxxZSQ
VPXlPGFNedq86gfxc3ydhJ2X1Q1PwSoLFHIMQzOWnKeuz6KIYZ3GiaI8WcU7Mamr
tJ6FmVCSMEqNrKhWJcZpyw8ZTAmVhPeZNESd6z9KIlXnK+rFxCZRBzKt8dyEeifV
i8jTuFfFrQudbZB2nxl/wY8tX4O9i8XC8TvBIj6Qn5lxiAYMKA4NkTPH1tDFtWLb
ZfaXN4+GyPyMt4wcYtU7cAvmGW1xS1vFvbPs9eXjz+6oXgIcJY53WNaR0/8ifo7c
yRTcMoXu1WWiBqkX5k+GrsmhfKE3aURhfmv9dkS1uCAVnI8djgSCf29HAmG5K6jb
ixluz1EYKOWN3QWOgaV94P+ZR9Ado+IIbfkKvxhfM7jm11WWFaWOqbMn9G9J5Hwd
126Kdh8tK7AZC+yQMxGcnhPs1vL7JXZJe7XqDL8p3V5Ka8ANtop3qHWhuBr+xK9x
8GafedPaTPORp6Pmx8498viqn2UNAAhBjQA2ziCxZgTwNQU0QYT0LAWQOUuwVBKD
`protect END_PROTECTED
