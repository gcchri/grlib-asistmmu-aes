`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g0AGBTBYnvjrv6Jk4qEq45rkZ69KWtaSsGXa4rK36GMhVB+W0gpNZpuBb5ghv5c0
1Ir2Tib3N7bvY66LIw5ki9V35TNODMF23FN9KhV1A4kGR1hFDOLVTmqnIZA71Q/j
6Hnh/LpNBeDDs2qq/BtxxcTsa5TxmW7aTOaTCkIkOt1HgrVdJhkAjAwLHd8dTPK8
/1XjgyN5379MRx+LVRqsTLFpnO6ba0kDlvqmvAZ/eol9kmfPQWqoihZc4uSBPgaD
BOyeS4/XmZHxeZJ2KhQEHXeuIXs+uAwYSlNYuYz/f6ng2ww11GZMf2hQGLiNPsVW
lz0RP+OXyrAT5Gp5lW+F+S5e9G1M3vp7uSG5GE9nDYsGe2orSDZfFyDZfAGiPWmu
WPVzDcg6H1bEm3LnjJCJOT7+DsR6GaZUwpH7sHKk07o=
`protect END_PROTECTED
