`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dpciUBU4PQDjO6TII3+r3GdSzAlwnUg3s5rhqUVDOToVuYqB7bSZkbgOjpMVlmuK
mt8rWb+YEPutDgWcB4y2lA2N2U3xDHXcLuqql6lcQY7j1DutMRgTdjalhTzwmwfq
u7zcfM5doa1FJ7xOsEa8yMNOHpVZgz8xX6m3zLhIe6hMN+XtbC83GKtxlGW6ajoz
y17vKmrk/F6DY5LnvY1f36g0xAPWJionOW6Mvl5qjTg5dGJ43H2jEme8FDP3zHFD
xQ7o18dBPW2v3oI2M25BlsQ5X3z2p8OVooFznoPrDytKeX2UhdzLC9hk11xIA0ff
K46dNv0InVcyBIW+UsBGaxXoWcxSQx37VtfGmarVIjcqvYzCTWWJ3h8OAbO31mXF
`protect END_PROTECTED
