`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DjSkqA+kh/h+Q0xd7dXqFTACZP+wFc5dyEoYioPdsmz+hO0vqHf7PqjlrAuMJ2Nd
ZY+lLXsX3jtaVjwCnC4aKZnGPGVDzDU4OyUIw/AmCQQISijzMHu386ugLURnCtro
wv2Kzya+pspSBR1llKa1JJMRkerMUrRlmOvzdBtINtyuBdA2mTGlosAN68Ua6TeA
BGNApourykSPkzenT/u8/uvYgw1CDPdzHjWiEDNkTdwMSa1LybVqntvRygwBJOf/
Xm/lkm/CbyyDdc7mX9693IUiudTzgfQzZUTBUCCKSNktB2afVI6s5VCW6OnYhes7
k4CPO8C+tmCuviI6Uw7pAZpOmJjC6krsh0NDVghrficMw6m5/Xp4qG5VL380J3KF
pD1JztXWCMX4qYtCgD4aLNR5X210hHtzy2dG1WYuuQvQW6yzYaIumwZ3ywc6AMXD
Y/4mjsdJYtUi182XVHwaSVgyi/N0Enl56/5E7tZ8YdwXbiw8JL5QfpnwrsyFQt1K
lcqKg329l4TItuF4boAhCfUuRPGmyNw1cdr1GrhTLcfZrlaXFUNMIJH9PaJegwER
cRDwmfTCFNu13YvWgQdsExTkRaUTQo7yuFlhZgLSk8i+yZLWdCev3eALgeJPADTB
IPHjn9PgZc2UY4exqrY3MlAuQXgA6jADszYW8cxoBowsYUdzIgtM2vqpvRASpgV1
3VCfBXSn4ckHz6SOlFuopBGGCV6Ux0p7+MjyjN4jY1HI/SHxcxxi+P4GYoNfjAp6
fA1ATN9CBy6ohWwphQAMszymJic7X0TROnf6Q0ahiw0j4bxOd7+X2uM54yheCpHW
SDGqizt28Zyih23DCsq8E690wc1TsKyx2i/TTcyTlf8f2Uuv/e+7X2Blisk53Xmc
AKfbTMl+Pdy1/bO5Q6q9RABh6kvZolbGHYq82rZxCf521VCyRq81QJxiE8Xzu2Ag
1Vc3qp3SaZRmm9VNHIiWeSojwB0RFPMiO7eGLhuN0D2f17S1nrxxPiDHw3QHI5fd
IRc62NRf2j6asQ9ZM+iL2XnmhoziP+xJhjZcNDlsKltjvgi8Us8LDCd7And0fk0u
g9+c1f/Yu557P6AZ51Vguy/l1oYgi3wCnPZvSujkk/h7DBYc8HRGKXTcoL48/0Tc
9nJ645HntL7t7b7L8cdhkaOt6QIQI9nmVnsE63k9SkEgB5QZcZgl3V1cP0XJr2ui
9yQ82kjJ88Zdn2asz7dbnS5K3xDjMbJxtGi6qr38bZC4vz2LMAb0o3fBILwrTjn1
4MNY0+Don+rbeC1AcorJZ+prZIkKrk5pN5r7smesnEqnfJxnNRQuDuS9bXIXwbQx
qcNIsJfhgFZoLmZQpYUu/rxdIVgGFmFQxiuhnwgO1pyGc7J5xCLId/PRl1DDSulA
5o1A2/7/xsozE0LPxPa21++OVHMb1PSWmnMYnWkb/3IRCYcXbnyx9lHHS50QqeNY
8OXG29F2VRVFn366yGSJ82vjtdaVVEiGE6pSV+XzY6mGzO7Ovoy7Nia1AtaOB5of
+XD6ZS+4DKGAAqH2FlhRrzXaErjMx3bEKjlbjq4RGCv+mVRT54KBk+nfno0I0QOU
kCJvKjDBi7oM+2adZobBB1sHMKeObTGkMU4hCy1tEdZ812gmV0miO5t6Ki+gBW5S
0HCxcvPf/gWGHmhXbhMXMplI5r5jQmDNECr74mRM8WcJem6OgPoObQ71Fji10EAe
QOHXe4e9pwFHYOCwo3qMtGE6Hz2CVPeihDTIw0YxliQfn8Tcy4ANf+LRZMylAnmG
6KWDukfSC6bpgcKL6aUFYf6ixSS9XaimZRcZGWaB2nwbCyj95nWOQ8MKebQqGbLR
83xb07/Gfv5vDQASxR5LCHUSET+aOm8RlaJ1Th6F91Anc1jMdHlfpWk93xxoI71v
NWy2GHgRCvreKUZCHGe4tRfnWq2LVe7gZHVGEiHN1T6LsG3XNgoqJkEg9K0zKE6Q
7Y7WNNw8FW9S8ey32I8OszrQoPab6DpthgJCMrrz3qAL3wSVRS74KtPWz9XwWOJD
eibatmGXWmbBPKic/GGRtAHE02IHZYLGvh7ZvIdxE+a6kWHAKVuBPQxBZmzAs9MS
UQJgIaEpfHs7nFEGlZFjkyrctfcEdJ5ZmHSgDmCfah/5g+sNkKMnk/vCNIHC2Y/5
DuglZrh5WJZG5gbOSc4nQ2hQEIxwULLAjBwNxd+2yvWJpo6A2IzSrKY1izNULENk
81XlyzGpZxj1YGe2eDE6ZNcncVhfyvYtaEVtZjmyiAtjMqxfsGZV+FJR1oM2Wi+E
O6+fZcUwWZpRFGB/3P9QRTfA7YgkJz67ITQoO/MePXegvC2wN6l71nYzdkIAfo3U
MYCkh3nzL1M7xSFH6hizAXipf7M2l7A6BVKXJqOPqsD+m/1i+EOc9vd8nmgdkdFe
jiK2J4McQkJvU3DiIpX/XbaBWWec8uxlAFSMhw4w5PMFKCiT1h+kqe2WEMFO0nos
xwps3wcn4JFqwGgaPcdliHFvrbvYZWCsgXgrZ07PqiDQw2zj0WxdFdr6F7FMMx3I
NnpV7FFczBhHNj9wXA7T8gKxg4x987PBjWDIy65ZNrSpN8lzIShF93slaUaPYnog
6OoRWKHGtTZNR7/aXNobX72OU93PIC2scmJuNoCJU+1YJIMR8oyIa6cEmc3QVau8
eDOnm+NIJi0OTtJ5dXj6m3ZANzZMAZDwYaYmJIcEBrfH4xzzpYGPhtOkf0A3c1Xr
frAFalZeWeZHpGmGj5+hZbCaM++l6DGV8QyFwzFsWg68vMOWbzJrDqpFILn0vggy
rvT4xX5txbdvQltvUNujBpFWg9cHCG5rKcojRlx3OoAwfxmlKG0MSfOZtvON2OoS
PNwrQqaPNBKr9lRp+LNAsamyBr42tfmv8Kl0RQhdgWUNcCYKNgLq2Y9LE6nwVaIY
T4O23Ges8wyMnKL0qN8OFa81HIdMPeUFI8n1FsfiNAVVOcI97HCB8/LGLHWi0CtG
ocqfssS1QxUXGIapw6SrbIMej0YsV4l+gCCEwWmI8FoxUci1O6CWYY90+X27wkl0
qLXq3q3bOPGRa+R0Ou1oQjqjwYVlAdVQpkeDya+/6nO5sj87ASJI5kPxfkzzsdl4
Yp6FBR3xLgoyYH19TsEY/O+OLFbDK8ue25kWemZ+/OKCd/DfFOwXLYOBtB63b8de
ErVSQbziCTSBH0nyRA/OHIdO0zSb4ZCWP3TO6KNkJAbUhURk7JfJbzOm0SKkr3O0
RjqpPK2L6ruaN/ne5jO7bKJAD7J6B+uvkHreI5SztQYkahPMt3AX5kSbEBdM/r6H
6zURq8VgidpCGqqLoRNnxlF9q2/Mi+8uS46J/iyAtV0woBqkQlexFuW/VwkECupA
0ppd5fzWNUHeeoczeFXFTuQG8vQW716sNyt8AED1ORUBajpGwxxsTQnaqAZWQ3Wl
pJzgQ3TPVTKQT4gho86ZrGvk1SKHzanqdFH8hKckzwNMsajkk4ZDAoCH4scJZYDs
r36U7PYIAViM4R/2mhGa6ZiPVjbEmF7cmEUggenoFlZb2a6jGC3A0NSjYnS6aIeN
jopechQ9aq/2QDpdCTRIua/ANuL187rvghf/ZIJGGyNQDEs2LFv8F5BiRHBQoboe
k2IdaxnVDf4jXI8VeUR+GI6RHHpjbyWt9IYspeFJ1350iTSwoaN1+zf22/UdEn8g
cNKrMrMgQtdr5ihT0hctxfPa+5Zk4x6fRe9NIEvZNZV8oDRcS9m09uLsgDINvNsm
iCg2HoHKb51WhakdQRhuH/zAkHuuh2skcbJvj1o6MNDSoCIL+lEmT4bdRQgljd2K
VFsyG5azeq1PadQx/urhNKTu6ZdjvSHXyKvK1u/VBvgSRZdwEhws725fk0+l1qGx
9p3Sm+z5jrRJWcB2Us4mvoO4fkSck2uQ30YTCiQ361tidQlQoMQN7gAcvmhNm/X1
u7E4B8ItKr0dxJyET/muLPqOBi3QssncLtwiMpCgRnz9uscfsF/NfrWNR+4LSi55
Kr5KM84+irXOt4LkUNf58MDqP1GfHmKsQC7AwB/F6HpTTPA07m4uJbWoHRQp3Zrm
ZNfYTSaGpej2wkeD9KoFvJqB3lCoT16qFWMUbjHifPO1oc6OPlU6CAplYETIqNri
DSXhZTmMDKTkce+YBdD6U1qPEl/P3I0OqBx+BPbnq0XKiIliRYcZMUejKR/eh0h1
+9mrBD4dDmfYrYA2rP5jy6gl37/5ZcAjAQKy+ZQOEOvYhldo56acfOcrhPGNSbv8
NvYyAzorMQi8yCC3o62Gpies84Ke+jIl8qAYPJIae5Y2Hjr7I6tGVjGNXsZIldrd
Wu3Ct/5tXAD4DYt9fqZ04tKyrkD++LK+p8EIe0907sVbTmBjhlM08vVkbJ0Nqaep
ukeT8ryQ6v86UrVqEJJ8SFo0LEpFdE+IL5fI6UlFZgvQRb680f/vExOWb6J+SscB
YC/h+9j639h1/3MftSHK7JkMr8IYfikYL75Ky0v63KPy6loWQVbtCvCwYnhRbACK
PomRdyGg7dNDlvRpp9HMiM+HDFqcyKmv1WbOV+qUMOtA+OmeAkAdGLP7DyN5Evwc
PXGISdE36iDGJuUq/3JYJyYguxPIKX/tryNjH7qGNpberLcot4uJLX0vTDUmJfNc
MSssXUn0FhL1OJIRWDa7sA==
`protect END_PROTECTED
