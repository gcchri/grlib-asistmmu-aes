`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uB/M9zlEvU6pNsawnEVJdA0VBY1fZ8RjiuMfIx8PjHGyxMYkuhN0tvXrwIJDEINr
+t/bwAFsv5LEPuHpTDcJVgHuYGZx7mso2hje0oYHK1ktKypWPbyGykE7jObA1VK2
YNqEX7R+ERCp0AHNnwhUihjOtrU9vJ3mh2jr/lY+6NNW9/ion+1+c9PvDALW1iUy
ayBkHtiUz7J7TL9JvyNbE6qIERIdM40UeqdlVY5u1KPSY4/VowZrOOiFvPDsecBh
7Hv6RexbCdCiOrL14Pu/FAD2q5IeeUiu8awhP2MFGTo/A132Vs+KyOSZlcgsKuyj
5T4ePoUh396xquq/oNMC/YAx+yxFwhEqgXMwIZokgallL1Z1HzI7bmU4za8YUCKC
moTo6cvATClRjHLt4bBu1HMx2Z7BD3c11RUhDjzNGa2Eg2JYy9k0WslTDnN5ccm6
ygwJC2YrFOzQ/TFE8J7UoOHulfwlLXlDqbGKfKSMj9ekH5sQduzx2gaT+JVxgx8G
QTRrRZPTPFTpc6geuyufli7AebIL+H/f9ETmrsnCM36wI3PyzqkHxx66u7PXCS9v
yabZiwdGfcyYKAs8YJrhdFT4jblfcCGuEzpPVEA12B4+YaTIDnSVsCIaYND6hhIZ
nFGWak7ZUvpq9B2dm46/QQmko9vNAiKyntnj5Y+qwGKT1LKVYSjxKGPQlbRj9A81
+u4HgSu4lTobRxZXB30WBIrInSUBHdaqUxOvblmnJ0NJ6AvEUwdM9nAaiGtBIeFQ
B8vyhH0DdCbM2ZHzUpsLWMrbdZyCF5EYRmJXO+Cjb+YCfDTwFfC2X6bIjyCbA2jl
xUBijKe0bCn7JjA1/ihNXQDjBlPKslae5LcZ3aaFr6QRWZDB+jMxeQSqPD7MrlgE
QugICi76WVq4cBvhELqNEIRRTJJRrCx/ybepQFV670rDIXYbinN7ZoFZzaLGfb4G
8KmIbbOjPRVdwVIgxMLmnzE57bDm6WCOk1RxxP88Rg78FxXx8FJImkUGhr/pL+6H
I2Ib/x0Tai8a7ifhttIFWjy9+mBW9iq1nSv3vnq1I4HuJqlcveJuDzq8mph5EQ6h
5TGrjGyLP8II/TM/j+IOAdeTLey/GiWrOMPjbYRSzsdIBkYuwmKqfLoR+H3brKY5
hanjr7NPXhsy/RqYVGRNbJ99nwfccAISmp9PxcZfpm6unQ6dDU+iikHXDtD2qMOX
SF99Z6OE1kuqUDjvfpl1MhANon25dl4Bpb4On/pqr0f4nkkcKIJ6iTPMu53mv8S5
BeesRvvZKJUILl9nE3todoATGXDYpbn/s4P6Ml6C552UTKzvmsv1mloyb9wtN5Xt
nn/ksH7PR59EIm/T9Dws/qqp8tZYFNea8WxXg1Jh88OOuu6SPdMkEgOBI1k1WVJa
sq9Uz/WuRa+BrMbGkeQX4D9d+o0paRLtR/4MN8bEFvhOr4g+/UyNWba8yccopZ4j
p3FGEEhrfRwj8Ci5AYHj7CiM1t7utnZakJwO2STPb6SkXcp4MYjEfj5NEgelo6hu
mwZpLU48jI2CyTbJu5EfdFbL5CMPEeTSY3X8LNzmxsKSFTQ8KfCOzeppC1nABJef
yvOVcajLX17lDzwh93vhEhPT9OtLAabemsk58puXg9hdYbPgcqaKVh++VnLMp/Yc
QwB7980AL1EYg3PtzVENVmw8m2sdzf4LPHEaN8mUy0kbt4Wbh4s7CfzzUmvw7u6W
wFwuixSXVyvAPRMtrORcSDb6/U6UNEf/0x0kuMp/pG8DX04qkbi1R6QRNuVXvpMJ
opMyh3r4X03qbadQ2r0oviUiN/Ag9LxtyfHzBy8l+7e5Gha28MUm+GIuBoJsgX9R
3ScnwG0FCuv6WOIlN7Zfy7mW0JupYHToAda9bm2+CBPD8UR8SgRvVGudBskeUO0+
ZT+gd3FrkcDLs+s6HNGCQXAFWW/p9R6WOGSbAvPhZvuwfD4eg/mD99txu6P+J/9p
E7sf/ESeave9PMJnnPGXIQcgY15lmOua7f7GC0rVfnSfU33cT/Meh8rJmUsLWsqd
lLlqVj+kz2A5eZR02dp1Tq7qhP/HzKsX6TUy+PFYgzsZ/L4G7XE9L8ytq0aKuvU+
pIQjAeat6pL7ntnKAbb2TzzMmAJZNCyoDvAarkC1/i3y8pcVSYKe4CDPNlHsFJeK
X6sHq/gDroRu/k2lVcPtS4lsUDTKEtc+VHRywrwjIx8twxyijFpy4QTF1Sa52xLY
ZhSNK6qCTVEGMlLOhM7eJC9SHhwi0FRKA1XOCRQ/FjEDeKSgtPG6MAPM2hCRCVKq
CR6aIsYvpfKXqhzAugu+X/Yhy3ctz721tBJ6p6iymkP5u34abfjARuCxgF2Y1EEP
X0K399uWSoLRlCElcoOvvwd1gdNTq4r4sTpnU5izwiIou53o8jdQ3bQpmthaVgXh
Qd83YD73eGefH/MU1YanKpTeDw1uh0x6ZvCTnt8sn1LKikaL5lr79v4ZVgiw4xZo
ZiqYAO4WJT90k9fC6ISFCKllAb/ySx1gY1ltA1bpJqC7Uz4QBBoh1Yp66DShLK5z
MykyVtle+du+arBNC/cysLSIKtsvOO9oh8SZGgMNlj0+xQENB52uqByFcFT6j003
wcTZhtp3KvC3n112k18rDDlg0RIHZRKFmNm1JEN6JjGuPf5xL7XN282lXN/57LgB
VbqYeLRJ34uM1iiEA5yEuCMJ4IqsadRZp/JlPR2tnG0fUb46STcrz3m0/ODvGoBK
yT+Sr2VFtTsrqL3SGkoS3dfT7paM6zF12r1z6gLAbK+xGIUht7SPnWkk0xzksznz
w2SCApDdjF68LUIPlPi2IsvX7geBYqMsBtNqBlm9cyPYbM7Z4zF1jQ+fKXZFLycC
8fyMf0CrCv1vf4fYjtQBp8hgVqVPJyKQQJzc0a/h1/jfPsvYTJTW2p7fsFkqninV
KPbOIWWRLcSHj5Cb0+h8DggrBbGamQuYY2SYPrvmLprVT7h071kaLZC0ZaPAQS/C
uqePWQ6glgKtYxBlbRJtaGEJOEZ8QyeX6O8qd17+ts2H33vtowu2rNGx8bo3M3jo
jCEhWcFUF4b+xd4eVbCVCBhem5RxrK2qvtCTLK9gG7V0Y4BWlQ0MbYY3yFJnw3yI
vOK3k3mC5IwQCX6wPmkcQNR8dUKRmdjZcaY/W/UEN2j828sIqRK0E0qrhbNH4T6e
b37bTi/kbXthncVUoYDKBF8RzD9Q6cdEw2VM3jOn+vC0BwJrJfWRCmxP8LG+gr6R
AKO0WO5yqp3hAu54nnak7WBHs1e7pNCUlO7YiU5Ke+oFUGemAQuFPqFuwNVS6k+A
1bLr+lHG8fhDaS0f1qunynDbKaXGGAFhuZ4WjMwGz4gQ2+jUCCGSR+SrtNIuZve2
h6xCzZBSKXiSokxYvHbDM4DP0/hItA6590HKOUdIufpa0GUuqKSmb6sn1c71YiF+
fxRrDhJKXOaO6wsz/LJ8BOUUhBLq703Aj0sj+roLdesmNbc8wFkFuZjFn6JD4J3A
7lWPJGmVv7c3TFWMmiJpgA8mXyATjwtHk4G0C8VTywAme5FXuTNFy5bmWSdhgmzS
4wzu1WHMIAKFps8wCVkP3WGgjCV8pdG3VsR2pHAl53rfmEovFHCymGsTsRKg/jqj
k3D137h9wT9vuGPeG2Ib9ju6SYoVPSRdaYUuRR5aSOUx+5Zkc4LL12wMQ+ALY3ag
qZYdxv+iQaTzblNJs8ACIOoJNh6ytd8XXyjwZZOoLd99+2DgqkdAO5NTtAty315P
akFRz+DbTEETBZqKiWLWoe2Cacq7Y73ZKeuFeBmRkUsvlY+l99ogaGCOxVgAT+an
/otOmO18/tMsrSUDzf0QfbqWezv9JCQwmK3586M9xxxe2oF+SBGvXCu5XOqIzlqW
sZUN6JjJoUl5YB0xlfVqupTTzFfBza6gqN5pdH4zQQtKyf1WjOAjOuVs1qBsiaOb
FCRJuX/6zUM1V3KQ9cQUCi3i/XrJ7VQcwdr5XV1BPFg+jDCIYXF7aVL0bMquCN5M
SoRIcgBURJ+2GMjl4m8lLr7Dz+FSJhGKNgtu4Sk9XYP3l6bcyfW8lYbyd14KGT5R
RFOjYl6UkPrAgBYHhlUyXiJ1uyqwWtHfz6Ps0MscG20SSkrP2tvDmbjlfTVE1GiV
yRs4KdbPb29LJQvoirxJZVhQuhfEFP6n3WiViuHYvyuiUAHBXlmStfSHNMSCP/Ph
4cEE0581B+5GykKF0X25cnN0OaO/049DhQWOuiV0mEpzJnVEPdA4QMYMXc4+4MiD
2NS1iuKg1wVVURqtUpoxiYdnQAcCt0pi43a0lG33Iu2KTi49Nxr2CiCKHgl4tL12
wd8WuERvkqpG+28OMxam73bGE9lZxkJLr7yjONW4X8QD8YEw+6sLiBVpkDnI9CMw
Qy2DSfynHQxAnwbHpZhXm6W8vMm1/7NvkTgp2fEZq4a/rSSTEyqr2OrDqGYxfK4G
Hiyws5dohxT9+ld8pG/auG2lzQFRvKiEyr7qTrC+/mbZ4QQX361t++thGovpFS/L
66MZWa+8OLv68UP+XlckJbzZjL3J0ek29ENTJ8hBhROGED5FCGNmAy71Ls1RIFh3
CY3qoKorhtEqbSMl1cdDR7LWgKqzodz0sYWrDqamISwXamS8zpf/GbE4ythoGXS9
SfByW4YpuoddAJOchKVtTsD9GXTUvIc+oHg9Sb4nWF8dGHqSKH13Yuc+bbVqIIGl
r9hBlvUHPa6RhJNoNMj+PSYzDn3NFEvHdc/oFpBqjy52wZgQXhIZJQVeO6PKj6j8
vEPi0d63+vAPeVeSx0TDj8G/9+UY98fOWsXCeAk4HNfkuPojz+hJv7QfupKOBdnk
qOdZtqZ5e/bDjJtCcvGPjO/seMJcCHHcf9M1Y12d7QX8DsxBgcrw9zeZxvN2s9SB
CN2wVdQmvYrTLlo7rPENWd5V9etpd5iqASrMges5MgnIGnslEB0LvepTULN+DPKu
MI+MWTLuGfBFv3jCGTyzFXD1VJwHn0OAoQ82Jtr00nnMVy2V8Zud94nyqUWf08cV
sqdG9NGwYCB3qKBJXYoImhdvz6oTrxRYpwafSdPjh/6nvPnGpC/rWBx+ateGVPVM
iUKJkFVntFMFhqXfUVN9pvVd09r/XmeandCHOBh0iS0MPr6hvgateJabp8zCncve
UlNB1bPIb6nouGO7T3f/32/yPmVsx+XPbfSIu1u15l4vfxHH3KmFYHYGRSPWuUmS
LcpdQKqMnqq1Pas2Oxpj8q37XX4vXF2BNckQQwH65/hDFxxUZy+LyLvdAY7Udg9k
JQr5Q3aDRmKY1+Tskh6pyhGvOFqqSK14al1xHp5tm264LWKSApUfWB33OishkkTv
vv1aqCJWk7mSxDZthlQ5Jdpsb0jxuyW3VZLAb/w4NrHdOuHR6JvQpFPd0oIUCCXd
XK1IBQQLNogaf0GQJ3TqVp0ZR5HFR3nqku2NOBJqoElLxomorWHx33WMng2q3dDg
nAMlxloFMA2NZDJsNq836sJKT00eXqRyqv0acqS2E0k96nQVEBn5VbappbYe8q+k
IiwR/xBXTI0RWkevnEb0mO8aQngjUHuq8ynyO8iG+bry7/nTv7uMJKY19s7Ov9aZ
FftyOD0om81iYXnXDQ5m0NKjCft+gv8MWK6PTDPZhYBY9veLEYpSu7B8MldBShHX
GSp26pZerUwLF08yWuljeYwaf/UrQNaQY9DDm2KynqzmukirRKNPZN53AkcXFZkh
fTbUCmKG0F3U2sZltAsY1i69f9QyMCipA4Dub0NQwVjeXoFhdKKHj2QOHqe78Mbw
V6pFyJNkUI9u1VLBefjJC4squRmt/RueCqLNn8tOVLeLzrRSwqvUNP7Zc9mJ/Mtz
e+o81r4AQ6I+85nbQ0yt2lU84iDga2QEHYISRyi3xPN+0lp055tMrGM4KXHTLGwf
0ioborg3I6EZMFnjS8eSQS64JmeXAYBwCGobLGhyKto4gK+HfDcF8qcSShxwLdka
AlvqnwYElFznKfBCA3VmUmOMLgPvxkFI1kj8ZpziQgoomnktqx5XnR782MQeeHD8
vR5OSwCLHCc4fjChcFNf3riWbeDsmzxNMdIE7Xr+5TH6U+ACIKPL5hxRe+X9nxcA
8ikBiSxyZa/St39xtzsH2OjR0xf9CWXHPy1YtdmSQ8ZcXfNLZ+7doINMu/Gxe61v
nX4t7uiJePuwQSso9Zc4OTJrEbQSzCAwaQ9OGmgnv17l1QAfly6Srn5nj+UzFX9I
W2IvmzvHl79WvDRm84gejBhCrMhsmjjxG4bFNnSPrVQ6pR2VVkT43Rsbf4+kzvI9
HxUJz/Y4M5luzJfHudD31WThwUtbV0lD6UssEAjZg6boIWPQAFiXLhnPmhaeK/u2
WzdI4r2wBzybH2xaLepezVlXAPUaonnyI6A3iFvrOvikfxfP5Ee+TYRJCqkWb2Y6
1TC21UT3Awy5+0Bva3L9HHZYfnnpVFOr3t16q/pfMTCixZnGA3LlXFiZtrd4eig9
hNomTLQHs1xJH+m1pjYc4IvYR4xcvhIF1bUxRk1Kb9JRYSkaB2X1eK8MbddR25Wl
G8j3svd61qOzW1T9VWBtJVL376xl4PqjRO4/673ZlNhzkikionglx1MdslpfvyWZ
Bi6cf3Al4J2rCQXqCjHF39dHK9xKtlM5mRG0C0nUnsnacU/zIHsBy/sARy/tJ3pR
N9esp2lsyVA4+EASp7RVxxbns1SNcqU5cIopv/QrmELWNq703MqE5aOBmR/RsXJx
T6v7GITCm/LmYg7maElOdYVyCE+WqJ8VPvjWOXANR8SYWrMoo2LITc1rvkb5Ou9e
sH8PAdS0AmwpDEO0DycAOT1p9J1U1CUphZHreB9IbY3ImVXuiW31RLZPyPbis59+
la6SwVmV4ZlcpI+90L8Otyfakd7Em7lpPIdU3XmYCQbxUrGnRoOzMS91P+bI0UwF
rnOp6CrOBpPE26y6Y4apAGq71RVrph1hWmVqzBmkSD+vEViFqJq99M5MP+SoUsaM
OrCLK+9zRpqASdrib8HnjIjvMMtdhnhiHKMqR2GnuC3U9GSSRX+dw731Qql02W2c
995cIT77aRreHNPkNL5A0UcwjXe/HLri2I+5+V9GgprWvQMNUCiyaFhhX/b9mMJ8
Ilb/M0Jdp/02w56sz1dyyWq4WB2DpRiZwJhBRdFfSGTbbao0hg4bCbDWS1Ig12i9
btFt8CswbeuAp8+XwatntlCHqRFvFSPqU2E3YqJCoc7SazdG/6zUGP5+A5odYhfv
FHlYT6KH4m3SuDe/GnPKIvZBSehVavOsOox21sMelavhtoIlLwOVsgd8qRt8D0ji
VthZ8T0YHkprGhZflqr9/NRJiUYb3eMYWnFIUJDRQKH9YnBgbixPeDtLg78q7XDU
dAR+/S2bJF0WcXCqwKVCQ4jbDIXj4z4MesaIwWipdlCdnIcTPcghm9NRypV91FvD
dF1uQC/tboi8KZc2gvsilhrDEKHn22bufj8CqLubbcSmIcF3oRIHxD7YpkKhTu21
SwRl7lFBc8mqLwXdHm65aTISkUnmsKMaTrJffKv6AxRefxSGBvigQ768OgrvV+T/
yNxGZo6c8dYDn0k2RhiQ/W+4oAWyMFxdqJOKGdiEuZITj4gSpH4f2RRJi2h8mxpF
5xMVt2uTMkv2OKjDiJQCj+u9jyz/IEt/e3dJSuggwY5GmLyQKviLGYc8ONdDV+gB
RcsfOmD4wf0vc6knqr7Uf00duncf2oHq0U/kfCDAVzW+In+fsrlMs/klIQlSzDKg
m/Qq+DfW6aaDo9VAwwRJ2SOgUvcGtsnB5bABxLApnTaBAa1PRggKsLVXrDeEJ1I3
9RYvRgH6uXaqakRxD0KSyj8jB75G4JL5mMiI7LFh4Ioeuj/WR4cYaHmCr1sR5lWG
fMpancXy+hgD683ygCm7S+2AOtGg7oJu6M9j7qKH98jo6lcCl5pWn61XLcc+ziXj
yeluZza9PPrn1GNPTiTq8kRtmFcGhhOs/QW4vkffB4/Xr7ZMAjPd9oJboUGv+lHF
5sL1maKS30NkgeflkkiqwhXvtnoPVFeVS0vEL76xxTGC5iWN5X6HPk7YF44HYUPo
i0K5qb/uqgkJCO3B9jC5xv2hBhKcPeELgTjPextG2lkfDVKXR3rt3SlZaj+YhuNq
ENLeXBc7U2jMeXXVu4ToQgdbIcTb8XSu5mgbGszxNtW12eqZDdJRDTOy8ffkS9Lu
zIy6C3iIb0IWTmNp+OBSMDsL1kl7ky2OjaURj/bpcn5FtVKPb9xwmcOds9ZprbwP
1XX0RR9m8DVSUNivvaBahn37TX+KiL4+MauN98Pe3raxmRi1rgu0sYIlUI9s2YXe
dLbOIaWbpkUyp3DXTOkVtJBE3yYyOKKY0B35yTjDMpzaXf8AUbrKknVa1OJg/R2x
BTAH/jpeVOS6RXznYVfYNe7S46zR5FIlUA9kweAXBkFvhHHMpSsAJopyvM4iiNqY
GDsVS9F7uwecUvxSFkS34FbHjKG3o9uYqCWJhTkZj5LIVgFFHzaWwDAWICrvVqnd
Ne3p/dUJwNtfdX1mbjdaebD+yP1xb46mSWvqlNXyAHSFuKR57A0tUpTCL7JCa8Zd
HTu5GgKMBRAWZd6LA9iBWswh2LykYNZOtiBFH7GK9Z98SpyCGhXVu8qdKlHQ0C0A
Eooevik3fFDyUzoi4TKdL1r6Az1Wd9oGpNp0QKGvHYa5xSDcbiW73VqukWgaRFtR
wH6zdskU09mCAAsGcStEGKLoGbyZSv8lDtnQO51m/WTt6yRRKi2LsvfN0hbFeCNA
L05+rMavWgjaP4PhsdhrZsAl9LRsTfi83Rzg+vXA8ljC5TdIcf6sU8g7m5d79d8b
VEd8Na0+0tv+prPmSpEAzRklXQYnlpYKScNKzOr+xpbu7Cdz1E0bgD42ya0+cLuO
8Qtw+PHgwUTevOK8T8/0DXHhqJPOJHgHhhLCNJpXulrkQm4InrI+yS/3zme9Wub5
OoASRYZ0ass31KLS4tZp7Ff1Mk28JGgLkZ9eVHE9MTijyRehsGv6IJuQipoR+TXM
u3la5u92oMmcThAEaIRGIvTRyGbpc6JrzEcrk5i7N/GeYgJ9Zc7Be0xRZD83Yk/6
pzUM1/QLIl3lnkrBN5sr7tLvtgMRtjVIcwZvr+EsKXup6R0CrlK03NId63ox95l4
F6K/IiTlDsZS3s+Of8eekswgGEFNf6xQUEmlalPLiDc3vWotArr/VZvHaRXKkarf
6oS3Y5gu4ZLp46IwgjFeiQWrR+pbST7ZxYBTFdFAyXutIfSzfWlJcmhEn2VoSKQK
PEd/TV/e343SiATs+4vHaTrmk102ahaHYzxl9AJdUVROkyQaZjHCCGi5V2zoNZ73
aut1L7yz/4hqKJTrmioFA34GTnvAOXaNwIwN03pfBQIpxeDTtHxQDXBX/X+Q5abK
186Bpjp9Q4PzKM1USht/WYw21v4O55iQ/V/nBaA2+1mq578chY299+NAhC9GOlNi
ZI7lAKBkKcptkDEHj9N60gd00lvaoCBMaThxKEZTf0VbGxThEVzYCUoIvn3M69ap
q1KDB8QBKTP+2EaZMem3eAFPSIgiwWN2dbC3rvvrFzNDUI1UNSvWHxUxBCm4lk0K
gs6z6gLPzpHQeSizKvGo3YKce9W1eLnn5iYh4fI5nFIy2YKuX9p0NhPdNWqOQC9V
okWVOIpY0roXEP2bBJlYJbhhZnbYdQ+uky8xxY4cf6HMzaG0N5ocjBzE78kFKXf2
scJ/cKADxJ6WM0g2RJbTcXYIXnzoSDsUuEkglrqHnu1yrHqcuKjDs+k2O1UMyCtV
u522JXW7ChIu5EjvXWXD7SKErpJVxtfX8m4DOXxpNL33nl0V5ekLH4g/d3g0g3/j
/EHVhYFZ+2il2sFAH6YlHkmxBWt6yaefjUpqPzwFYYaa2KGBIhTGZpQL9kJp4Ea/
ke/t/46JNAhL96yIAXsgufYxXiZenVbmoMs7nBk/uS9R4hBqHFy3I7FwY0PJiDZK
r0Sg9qu3BE7zfcBcdRnFSB0/8ct0UedB3wPDBStajyvDPxp2HmwJKomd0fvaQs3q
dMD7ziOyH31+JhGXG3K2wkCzfb3+5CZFYHX/TnOCZY3C1Sp1hUICbgXdtGVa+m8y
kgH4GS/wY/qj728vEoAnwiSpnpwPqnv0OCS8PF/2uUbUt+QRjgDq3ccfhCUa1+jS
WWqAyxD2dCQFHEL7X0pqlK1/zG+BQ2ywnVtbOBIYb9PCprK+W8dyzEMkrvy/jPQM
rhuB4V5KnkustoTOxae+1Sk6wfPhCxlQWFDfhYnAqcfX0aiH/6tzZRDoNKZyQC/E
/zyZyE+cS/9oQqFFCTbTlB99G1Yd1pO247VGZi6jOiDW1r8pIqbsjTks/hulnwYn
r0EBK3cmagMAo5Ud/MfZuprt/YR1oT2Lq6EEb5a0Avb5juTpXsOZ3jOTjJzh9wmU
e7NvX76IxMuLa1zbaRq1hWt+mVMAI+jIrg0dawtVh+zYMi3CotY5nDKdi8lnt3H+
l4in9vYqG68LDAvCHNZTuF/LjQPkqiHDyhKGKILWfLd7R/vesd5thr+XVI17wIjo
5mCuXZ1u4udDKgOnUkEjW5OENhDNDoWrzn3CxEAIXHzoV8JSxYNo8Fmb2KqmuOtU
AZt/81MS7UcSGKN1JewpCH33lI7XLWE+ZiDms2XCzQKpxX76r6ywGJ2uCxK7I3mj
fwHtr7aPD4axonGYQVTru6dVgZzJNNocT+VLQDVy19ULKjRKuXpkD0Sa3bFzymeS
bfcRQrOh9R88pvSKMNpTYy0O9fplGzm5YdTVKzwxFnERThz46ZnQjkhPB+tup+8a
8RD7YRrEEFW2WuibuI7Rym/f3fh0uRCy+PQKsH4UgWkCLdt7kZZb1rSzcR77p7X6
XnWq16TYyQlcV4wg/1YquBREQhrzTlEGQ9fynhyspIeHG+sH4En2J7MJRuJETPZP
yMvkxndOhYJxl3WwhFyhYyxuFb/Q2D5QlM3TLDTnp0ZdLFAR4PVmzvgA4h2kk5i2
g2fwvu3fYd8iZloAQW7+6J56lRHdeK0cy7gbIRIj9IpKzrWhrztsXjOyRkdjCik7
+9lIrjMlDcJM5M0sZnm00BqEYzflOPTpMqRKcfIn4XIy363v2ZtbqxTXtdery6mM
o6yxAbdxmAzmgu2f5wCb426yqycezk9Hnts+es3N69j88GsRd47BNjY7sQK7sJyf
VI7UnnYiDRx4NKhQfidC7Z0PvJdeiyvSB4t2bcKjWJjFY9wm6ArqcPwZ4MVzfVkg
77XZ+Hv3ilo9Y802YznUd4QDEG4vWJbe8kdFBFodZGfJv0zaOlb0BAdcI/he6V0e
xKOhUMZoaG/nM2WkVpl5/EKkM4j95KS2sAZKt8GE/R5JK3Cb9R1U33y39ILQqYsP
5b9Da8AErXlZezWY1hhVJX4atfSTh76a1hOuNXAUr03Va/jDm/348IUm64aworq3
mWj4hyDGZM2J7qikEk2jSV/5wvSBzku0klSC2KCq4jTa0b4wcy5fnVwrKixZKt15
uES+1LDb5+OY8Dby6IF2nksk2A8U3ps5TdmLFonvAIS56L7JKNKmFHGG/4NVjUXf
rOjWnO5AnCUCjPVUgZWGzH+oAOEA0oWTyUC88ARvt74t+PnnasOWOje1AwStyvr/
AGbPjbbN22jiZymgHGK7PqtWWKmcZmOkZLR9cCpT5rg/MkX/jrCcDmXHcmmOOkVw
ALdB96MTPvIG8AYUqfk44rJoMR8iVHBXDft6K5AmN6ngbrP5L6iQz9R15s9Thqr2
p34Sk0hcC9cUcrXLPm4QHOAkkGphwxwuLHJYx29Jzaq4vaSkM3y58H2HBjeiVuRD
MVoDj7m4t2/MB4asJZJZ2q0W+7BiXydMK1DkCtQ828dO9yQZgEE3Wx93cNx2pp9i
8TOZgePwrhpbwTtYBfF1FGbJBE/znES4MTEHWpbEenHtzQM92PYwOTRG4QfTPThw
Xs8HFNfLQ2FIHDAkGk7wd9NpkzwM5vfDl0ocH3ygOr9axAB3G+J07/fkZ+PEdwmX
E/UaMMbi2qmjH6hNfFSOMWc5ewWgzHs5KaiSgh6usF/ockx16xNZAfhI/o9NouiY
n6QPPhKi3Acdns0bhqCYIRR0djF1rOWaBeZHEAmWV0vSCw14bXfYYAS8q9WpaqGq
XzGgsqPcaVztqtMWVkAxKwy/Y7qvkmmO7toShlZ2mVNazhl/B3LoCTSOLSTmCXqg
d3F9eJSczES+j19NIYC61REvDVfp/4ZHwZJjrjSRdYZwRnJLiZYs6WDsHUQqoGAS
V/nshVvmm5fF4EWah/Luk7KGTzFolFAuKDTty5LQ5ZaA+ICevmxe9nMutlF1oOV3
GObfjG1MFNVF/0SW51dOp+A5mM6HkhCg0DmO4U7fDu/zkOF7tyZLnKf7ArEySm7f
9dT/6I1NwBA19s59TP1JFrr7uGqBRherr0WFtsYUER3f72+nt8pOwv7fcM8878dL
dI8pT+97o3bwzW+aeDEcuWHYZfzvCdEWdPC13WpCO4yLXtAPG2AxgL8R5eW3Xh9z
bqLCMIMgEa0b8SRSkXCXwI/jNmuJpYNSDXY/BgadzB3p+93W85oqgGbMs4+3heCw
FWeaixrYEyr2kYQkxOkRUDoGQUmLjUz18rEFCPvxSvc0+sBdOmaefLGOHxLNvvo6
pLzf6b73Q0U/rGXMxdOt03aWvT+Qmq6KUn2jtdSw59IWakOjCTs8HpqA7UsBQaZR
84+j/uR3LpxwHfkYcPCw4J9lurtNSHG4KLqnkuxOToyCUdnM9a4MxEazxAtcwDfe
JMOxlGzubATtazBI1xvMvrhtvmlJ8eHx9KG8dxCEBnNpzYMBt9++Ov04pgHfTusN
4TpJWY28600ppq6J7qeEJ4i6VbM/aCiLMa3LYXgQWg1dw48M5ToJ+KG7YGkUF3li
egMUufaieyYW/Kjege/Fb0twByIvuhgFkDe8z/akNheOQ2Jqrreor+qY0GmXrpiv
b3yfj82ljVBD4SFDf9VldVrzhtoG+B0c3lhowyzHuamd9PHExI5SQvfOMuABNe8x
+jd9gsHUrH/snBWtXEEVIFxszlqgyMIN5JXg6R4GIIz+EyE8+gRH0idbDQQ2fyR0
Cadg0g+Kx9LlYkUjaPp2Bn0TWOSqfKtY1JKq8DUhoMuCjCCXUFoOfVYJpIAj+gZp
c//Hu+OnKzK86CDAKdxpRrtFrX3Illff80iNttUUUYgQVrVdOvIOoF72B2fn1kNX
cF5yCAirO9oLJ93CQktExPNHu28Rb+5Yg0bsRBLuXgyQU9/cxI+L0U9PDxH6xIwB
5z+f8oX+g+FWIXW7lLWJMdOflCRcf4Ui9gbxsFMSvVjIuoLI9ShMIEeTfP1VfWFp
ZaF+BEX0XewR4kzCrcZxvZogejwb9awFHO2FoYw9XRU6N6FZrI+5FJue/TiRj5+Z
iG0G0CJPp74beGahI4U4gzA4NQgLvr36/EZ4nR0tctCwT3G7zQh1OOb7zsOtUGJW
OqO0zUFItrhCXCO/bwEs0sMR5GSUdqj1iGWkwQpmTEgXo4zgi6ExDCthttnx/FKU
2zPjeW5zyC2RVp4DuyljXow2JeE/6WfAZbbZ85zwZc5SiLo0vOBIH0kHe1GhCpbk
s/j95NZRSj4bnpks15fnr0L9EbvDSGc/26Kxl8bt02qcaTHss2QuQx7e2RoAo86a
9Is/V+BWNseBuxCMIzJx2ilavB5IeCDfJBccyFEedHrPRJ3tPfcWiG+NoGf68ZdK
GDEAZc9ivZeC3K4cQkDV04AteifpMeLVlC9q00OhWA9rHrQS92/aWHrDCKRm0PEe
grQgMPSpsGhdvVG9gw6nmnZuY8Cy8h2/7igKODJL5JhXQAUOzV2307au5nOsu06A
QG1oGkfbnpOctesgXPNxz0z5MSl1FB/06LnKgRuZd3OSk7hbm/gpySFz2CloA8x0
ivGuQvwulhShpnwSzrMzLQiYdLjviBKQbPQ7vo6rthQHjQx9rEAb2Lczrcf0JG1n
X75h2ZmPHEqm5deGuR+2n7i+svS6/8WwOBVH6tKHpBLxfy0hSZu6drRHdicy0U1g
2AjiIUp6GeogpCmYb2CRnUXgbykqnRV1qtENJ0UL/rPkuhvHp085oFGyXLKNHFH8
usxs011cNhOUnZ8LueQ6X7Qs2s+6Jsk99j9e5qIXBH/CC2TRQjhpXE1N9rpljQgQ
s2BJXqBcMfNG8979Sn/H2xM45qyJYnszdGSQbs2GazFD1WdrWSo+rFD8gW5XrBPn
lF+ysovdX5aqmDFjL+TLcBq+o4ayfnOGCRSFPyDQ00q+b1OBH8uGIXaIDlzsfPY9
sVts2E//rIi51LrMNO9slH3Pu+HSEEdLzaA+NPP6Sr+qXjlScz22CRzZz6pslgYl
tB8FWdSLshfjZrFz8T8PhqR+3LzVODOGtXihFpbSa2uxNRY0vs4I7b3txiqk2s50
BI7dzByY1CW0IBv1A192FP5ciSJSp95CGPjwU7sR5iMUlNN1NEqe69FTiZmBUK2V
Jnb+qfjAvYQcce/q0y28UjLbVQNxNhIMSyWU4vgI+XnPaLA5c5RTCogBCjZgxVgB
e9nSOSmtmLGXqVSH3oaMLRyuOYxahlKn+r1Wv7s6rQkIYQE0/8mfkkr7z6A4G3uA
kmhxBGgAI+F4wiwQah9lXjxpcjlWCCkPFlLNfi9yO+gqoQbH0JKj0nQF5MHgDUbi
XpDJMJkZkYbRoXPBRF+yyOYbYurtuKnuhDAmK4Y3rhUCZ+5Mke3eCZ6giiOg3BaN
RTYJFPxrnW3rc5moa6W1mJletfwrXfOO3E7KnhTQKrA68aTei8q3DdMETWdtITVz
UO1GQ+nEo5H7GjTsSlqfi82ptqzZbbOgkNg4Ux23x+mavcdy+ekJHBhHoD0oMKSc
VAKrpZivqFmr2cDvrNsGcK8cRRog6chIHCLNiumXbD62Qi5EntA9nZs+QZzR8ANg
VwKmpW2gka1uIbfKiO0iJiUMOHTClW23T2jmHy8pnbi864Go8l/BLYf8rtgI86Gc
BvlXlqCKmXZvEoIKsmmLKBv1NICgxu/mHB56JMRpUlO96nysoOzS1M1IruwCbqV6
aPGUI3o20F3GvMtFo+QBMcJsS8YS78xnl/kIx1AOl9/i/eX1uCcDnD3Ei4ztYPhm
mFFeZsirbJwbxDr1peFFbsex3V8I7eqy8Vrp82UVt9IJOtIn2iSC4kxHz6J4vukL
UjIEvVPzfypSGVd2kYeTzLFYHO0wp5UvqU9eRQeUCzBGAMWUcWnFAbsKiN8DJqMJ
6ZAO/6sdnr/9NML/bUisaUs5ttAKC3QDYrrzTH2XgvYr5YgPgz1Y57sEelxUMsoV
M3bbj/vgfhwij/WRV3BJzqTgJtHuaEhqtOQUYqClxAKo1FUSu0T1xkVD/VJ29e1X
mejP5m7FsjTjcQ2bo71zS8kgRJKXhX0inzvXVjtC2tWd0umxqVuFGpnco6lkDsUm
mRS1d9N172vmS2Bwdvma3LZWGDCH6n3GObV3+S+sitRIfHNzXQyA0TuXVurtrbRt
spTY8O1W8RDXRs6Ty4SRFsUJLfFxyl2G5BLf6qrAdSTN5jPFFBrUQN8PI8wDsFqt
6JgsOpjeIyEiB53/kT4/bpNVJiel37LNksPaVjsJLnmjd3urujPv73A1EOcv3WVL
41EzlzISWbVRZf6e9GMx+WLgWZMuKhzCxl6rqOfBJNKGg7CrPp9WMpZJrw6ci3oR
ZGSQkvGi29RM8DumQwBKRLb+wi/kgBxp2ywabpG/pNtbnuhBcoV7RSHfwOc/r4NG
Rnfk2SdRRtkYJIy1VNF31n/20+6ySR5qsIDTgzeg8A5wmaOI5FidfjnJKVKVq9A1
7ZzMOvxJXuCxdpY05xk3EUw+8tTXXc8ZKpK9gNZ3Kx/rptHkzkiYvl+KOnsMdvDw
9iANxFYZTMCn+8kzk4Tul2kKYAzj4xjkw/JgeEgel8YEUMmjj4LIYXVKfS+HSCLX
3E0fW7hG4udPl35vnmwz6Z+sx/XG8AKuBne5t0qhL37EdBBgzXMXsTaJWobs1FXb
vkdgRcmnTz4cLTT8rTOgKVzeG+JoXBwZN0J9leDwEWdNU8QdI54OIXFrniGB6yLy
+ZbHQ/UmjSsc8bxkHYomGYHQihAY6gQtlBw2hczjp7tw/8oOrhg4j5IYLgWMNysE
gdgFZ4RF230N92EOwUSRdJvjpPfD2uisujqgnLCWNskCXGiKNxyb25EHKtYkd1lO
HLO3P9ySK1C0fxK+SNPjzHcJi/tu74leq0H++Vc3VJvzY/69evlK2+Wa4J9YNjhV
6zdK6g+29a8wIgExXrU2nA3yiNZY7keCR2nqdtbKNy22nbNHIBPD2/Hyn9HCAh0j
tQenvj6JzF75NYN++ZTq1MNmf7xnMYMZfLSZuE/kK6aJGGw3sj87xZrp1Ir/toci
7N9GKDgHxELTkCDiI7xvx8pKLE2O9h/rWmoXUZHudkJ9IMuvyYzaexnltyVRLCs9
34Q5kLcy1kIc/pZb6gSv7hjDsB9cNwcLqv8feTfASIFB5gbyb8huSDtAMy+lticj
0hP8zSqJSjI2TF/TKKDIMr7OVjRAWLSyWzs43E8n2h9s02J1VuQxFMbMrefs+kRO
rutQvYPmmnM665Lz0hPdr2HvbKnZ34/rj3h6RGIUwe+nUTokl2Ui3fKhzZfpJsN8
8C9maHAvugSpnQvw1Ox97WDidPFmWDFfcLixpZWj6ZRRV6SxFeWBQuPUs/3iO2TN
fh2O3h1zyN048L22OBmFh/IXqJCtd70j5eyyrmn+vBDmniEnCPPgCp+HWo4UhabI
IMT8sCo8+Nz6DmbulaGzQ7cNbbg+9Na4UaGZ4RW130qyWhe5LEhXwTSfHVUAjWmF
8YVInCLeGsKUB8YY4vCDutZwZv6GvQI89welP2+/1TBRtJIlAzHkWyVVQua7bbhs
UxsDI+/LBaAgLb9lRmUXHCnYM6Tgif3JajcazV6FaY8Sfc19toxYIinTrIPPF81A
LO3y0brtgHqkUs7gAM+7xkVixYzek+a4aG6Yu5Yi52g=
`protect END_PROTECTED
