`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i2pwa2azRaHaXTnEjBofXRNPc5e5A7xXXZmZllxoUljyWTkx989WcPi+5UHTWcQD
uQyxOFOqJeBkuHOLoAvubvDVeGmBAtscAnkS0x6ECJ3DHHxhERiE+AEMB1XiREPn
YoAJ8Uydy7P40+XZT03oUoOe36TCLFEijhFXqsZlIY9qWVqOLgI8yJK8pzbqin2e
eoGBnpJwhzkXD9XF3h2IMWayYdiEOyQkY1zPUW2uhpbWVnLEI72P3QkqAoSMvLFh
pwb4nfPMH0BWcQIylzTG5YnaCKmpHikaS+oBeacfFlIgkGHOFK/Upwwq/0XxpUPO
fuc+4PYlajAlnG+2qMDxybIuuewtMX2eW9Zz7oKBP6llmg5IeDyRJcV0Go3VW83e
l+4EsF/MzVwn1DkrVN9FR1Z5QE+nP1Y3220zMdK9oWCFZFvRQPH9WyaebzXGorzP
GUKV38aM+N/Z7F109StGoSDnTcVA4bnaIsHxaUzpujjEveT2Czd3HyR8iwWnQT12
L5QC7A36KryLjPYhNq1gL5ibWXU1MeOyTsIczR11BZT3vRxlWdA1Om1ld845WN/f
Uhs0E3pOxU0gzFdgXHtcx0luVbAkJ7K4mJGgMOh7AfnfeS22XBHeKs9Hg5/KtSnT
U5cWvSO+kuY8x6c4k5bqXAY0YNhSZK+OotTYUQUmQyIo010M02XUtYx5MJj31c/+
6U8O8KZ657jEt1Ij2v7wfhPMmTywBNUz73VhqzZukBtlxZ5JMBwgoMKOHy7ieNd3
d5mYRUfPvyLEAUMnpmG6hOlqgvxtPcbLU3v7SoVwBL9qER1lwMFH/C+0nCSl8JCA
5S6zloTg3m0XFJsOVWm4m2Fq1EZa49mxOJLOcX8CMibsdSuENjdIhzXFBAeYoTlU
or2q1HYXZjgtTviDmWShsXJDsQWuSMleR0WhH0+QAjp+xcQxRPFbduf4QChKxYij
R1rIrv2/d4aHQliLVSzcYYuMoEHW+kovrXV6XJsakz3xxDteEHduuElGKiskld/Z
OMdVUUBHXMBPsgzKpwjn8EjmhETv5ok5xSwW+H5Wc1ZzUjS9OWs8YbMXIfAIGtIg
jALrD47k14vbydA+joWS9LSDo1O0CWQCxCYAIezslymd4jxuNgDCw+Xx0dI4IarF
+jj9ztq1pg60mwtLHovQkcEKb/EBDq+uvpE5IxijvT1eeViboDw/L7PuuTZQkWJ7
pY8VoqMjqHAYJNHG8OsluOJGctbrfTEPmZymjC/rINtiIXGurlnzqoUFxbEHGxsQ
e6MT34xv8EJqnW4xVFB3wI72EArLphzYMAZHQLWRQ8PlNAqo6TnsQmd+p33W94qU
qkQzlDMAUCoIIWr3zPhJwP6Rv/08js9+69ufexbTgJjfBL3u1/vRZWfZbgzmXVsz
EBj1hqUx3Dot0NIljEIzaAuaiOzvto+uKKLDezs0mr5tdcnmDPgL8kROl6PdeA2Q
O79WpMfvHW8RVK8gNDC/PaDGeX4U56aEuk8Y0dO1LU7Fm1zWajY0FwCWFQo62TE9
ph+U8UHJX6XJh6jRoV3JITYoes/U6nR6loSwjFw2e/TaOqFVdVwEbJPETU/EXNbg
AQjSlklb1ezcxnW0YaZaNjUR5JMiUyormVyJW7zckdj74CK+FDQfMNpeuKqKGYTI
mdYk73ENPOsp8/tpG+MWzz48iRVqHQBpDarQmF0t4J3fUUWkhgoe0a5o2ashc218
pUrL7/txEZqF1VPrfE5Ubsw0QW6PGhrpYa5k2We8C83/8NJH60pK3/EnYVZAKFYc
6655f6fAejuyLv5JVFyaYO/Uaa3P6nyyOMeUFZKhWAo1/p6mjUg6BcpJPVxrEnZt
eowSc0FvxAWJEK3yrRiB5dSymUsCX6RLbEVnIgphF7h0ekluzom6PVhBzlNUDcda
5hklI3Hiq8/jjNrHaZlDNYBwh6Gkmb5tYMcEcw67+lCGNpFamIWyfuhctSt9oDYC
UUejwsQJKyNW9PcB+puW0GDgTuwd8aUbC9ZQjRQYPGMkI1BCLHxOy0+kXe27TT78
ler5/uJo3cxkPofLgLmM+c4PYZYCWZPNXeNyuqFWELpeu1brUxWIMR8jl44/x6Jv
TMu8rmH+TxtijUu0DQyYt8i251Q5RyimgFHaT4YOe6fsT6baYVRHLg9hU6zAXakS
IXiQ8C9uDrJrK5oK7XQgy5CE2wDbWI3QiWR3GX2ztRmIPPlnjWUd3BgbJHX/g1qc
9NbF9YExHOkOuDIdexXmbrq8r7D2DCIP0nrwietooQo509rUsnN0FjNpEtd//VWX
HY5KNd57Xmpc5gqQQs+RiePMfDiRqmpMxmKaOmZO6sQNnnyFldqXLh/VkTGhwg1P
pml9leFW+pZBL9uWXB4/IBoTa6sVl+Jdl3rzI3fdOV0Ke4DLVHgO7KrgL1BZzQpO
HXoHZklPwssmwuWfYGlvXZjqqc5BwyQhZ2yp11Ev0jL+/moiIBQabm3Ug12bJu8z
0cXSXP+4pcwenCp37uLBLaUNHb83gT68telXgD5j1pU7eR3eIf2OPyORfRgW3jeo
UPneQKF8+FC0lLzaLUGaGQ2OSuHpdsDpT5PfShFu0xoHKNpNY7N6aQE9GLFbtEFK
N6J/Gh/VD0TZ7+qevUDHV1KCi3/NMwy9nCYWdgCsQ/BqHu8n9ho0mYJ8ChGPTBwm
aEQdrx49bXXgFBhJvPzX7VkjLmzpRC/VulV7W1+DPJsC1+S0x6ftPN9NY288p+ZD
UyQHgTSzzKnnr8mhPDnR4ZubPlkVeY86+RtUpWMsyTZw+ngxZQz7vdRTSlhE+eYv
r9MCJJg3e6O+yUgvpwh9MtRQ0mjTY2LwyCBiMn91VephJlOqDuXtA0+hAT/Qf4ob
biFsQFuDNRK2D8CVuOd3DwlDSw6MwJMRuYhAmS70HopPeYLRIdtQKar87z9umC38
FLHT2MWBg7oo3PC4zx6UVtgqIgkOBARBub9K/qUg/iyt8cISw8bHNsbdoXc2DyPu
i4boUwpnXp9QuYrL/HH2SDpwjk0Y9ce/Ep5WlAhdLrYpwLLzkMvTLPMscNbd2Ilg
5b9By7PMAYmHA4Z9XLNj44jmfVARzBK1ZQO1WRtoF+MDY0oOtAKqS5ggJUhbYVrk
PNhQHkO0NezRjx7DtCaBPsxrF/z7/35QDn0fI/khhw/EeN2uJ///tTqr60ewKbzN
R7nK31dq7IKbWJK+ojJpGeNzzAA3A8GJ2mBiFuuYKHPxKn+bB+isERt0OZoEgS40
7JaDN2vG7HzxZ/w9DHEmJRB0pHGewLtTj4Y4bsMQfgPOQUgiJkcAUrNPFUNXQYdU
CBR3tcMSuvskW6G03IPyVj+zSB++Cw3Y6f+cODYxvZ5KFHZksrXe32VMHZqNFWmb
KhyUHznEamzpt720agglJ97ptUIliMXw7Tp1XzT5ZZ7XhXqiCJs9dDfEkCHwZ/us
fjx9CMvsMya/m+Pwfboy5krEcvgEpwIuzXSWiA3L/kkQmkENdk4JGMqyNwPhAH43
eVZUDuVfsRhWfoDZayNjcod7cTOzLSNRqXC7390juv9spxFGJllve4Pe9DJjtcFZ
YVEUKHK3GFh86G2xkCltc+tOfUR0n0UFU35JkD6e8KvNGqezOH635xKk1i79ABeN
wTXJ9PM5dTkx0eAK4uG7ZQ8nEfPy72eXdWJCjlFdCzd6qoRfkIPwOBlo6HlhJzJy
0+IPRpdPUu6hVOy8D8bZrnFzleOEb9tjfffGZodlajFWgj6WFDbBh96AslAtOODa
81QH2pCj2HW6j/oYTYIKUk0aE1aLvWlxwxVXp0n52QauABwqKpsFQ4Ye3ogoKOu5
ecS2rLIblKJVTEDFUztQrXwjEro2484cDvLSRfYqFmpDMesvO8QSCc/ZSSswqDk8
aCMMSEm6UGQCYeQWNuOKORh/E4mDMd4nvyIhdJ/RJSiRcOM0+SZ8R1qX6e9Q7bs2
uuN1E/j9rOZWmnfd6I1u+XXrBwgxl3DOjqoqSN43eu61Qh7YVvSMtAaNi5PFnRNF
8vtbl5wEH0i69v29+BnFBdm5trjmxQCPodQcf8g1hyKPaMEhbFIJ5jHK16qhj3L9
QaE9kPTFOBW+rEDNm4GJnTx6vD48tuhZGS7eTuK9QbcKPmVu2kINUYLZcEXSVYsx
I+Ock2wtVcjJ/hBxyU/jJs/fF/ehFP6hdglDhyo7rxK8m9h8nSG7UlhCLHS92kXx
yy0QkPReU8K2bvQJhAhfGKW+L+tayTVbTqEK+UZ4R4u8oG3Cn3Zg3n3b8oyorwdr
XQe2zyRRsX9Oy1Oo/hw8wivllFpn2a/SizMiavc6RU87aizCW2h2M5DNUNA3FtKp
7ETNeRr0A/dnJoIKQ89PFmebPc56DGCOT+t/XRkkWZNfL6H2jzBjQz2hQJWnDI96
kJhcxsbC7HIRKMv35396R9eZNmJRJvz6KIPfj0neMR0Bz3ORbkMljWQuKkggtkX5
QE1oOh6vdt1f9te77TPtPqnTRo3w0LVqLOSn/BTuz2SOZ7lwJe46FvW9PaERX9Nf
zNDeJUmazGJIAVaa/IWy0tCKZ3L7B52dNRF4KC2It7AJVOlD5Bf+E3FTzo15CXTz
d8NDiMi4FcIeqrzd2GPwd0e61sfcpv7SnofwgEwz7slCxvjX++APhblJPAPEvjhi
slKCePOG1p6q/1rU7k0vQvAfOOrWXAHD8gd/21f8pGbe85xzALGF4zABFMqGa3mK
LxTmC8dWijXSa+9ur8IvDYdqvNdy4i+tiD/iF9guSaLRtl9HsMOd+S8EkSQ7cTmc
S7MrE0OtU9pPGbMtD3GEWxZOD285RtRIVFDGkw463zzogGp8EUqvII80EaoT1z4N
NLNGC1cnDAhHp7Y04d9bt5+SAbWy3pMkR+7wXuzZnsx8BGJXxsZU0s764QLmrRCW
V75vhQ6RmprnAhWOr6KlZWiBC2a45WmHL/yAOZPdRzjSWyZICUcsCb8K/uPdxMm4
/+CgT9OhMyoL5qeoJp/RxBconh1kU9oRjT99iN48x2tBeEmcDJAiq7R0wTJ27J8T
cDo0Wq0SzTBN/u1Yi2MSd1XkNpP686kU7/ULxZ6loWc3bgVrJCQH4y6mscqWodmQ
ldfVfieBsgkxvIKS/KlnWXUUaw8SjlT8HoURLa17crRpfx1v+0hLTDLR6S8B6QTQ
IZcC4NJ71SF3tH041zHICxsKXeqLEw7DiK8gZ82LjRv85HgBxx0QabQXv0P0tVWF
2xbvvAMY64Wz5WULaoDmkj4H4xaG/Tv1DPyXrOp7G1vlCmj+FWqz8/u1DkgCw8vv
qXqLLudufqigkfYuVYBVdSERDBcgbQ5wF/fPMy2WS2mHAYstdsCz7XEcSDGRB5NH
D2Q63wxweZxEUny9LjqSRYRl1yx1E2I0xd9Ava13fefXqyzOVsSakGwsYou/PFzH
4jmRpeuHKlihqsZu2GyHnw0svjXvPyjlDJX4PIE1WKgPfzN0DMAMPB9WBxm+tjBv
OAKaD2q+SMDDgpS2oUsvpoclE+bJvHUZNu7ORej+poo1hZF3sJfLDyFiQhL37Qp7
CX4yjNfy+BzqgTvI5jLCzX6BfuxxLPWCRIQGBHjW68HdzPiOe+RkUTYQBd+DKXx8
/ZFhabimsRdr2Nh+KXVqguvnng30ZRE3Q9YTSKibbt8emI9NN4VflnKlW9cS4yBT
ngLx8MtYlP5mCyyqoEKfPGfcEuk4MZ//bY12GjDOawO7FHru63DkLL6zU2VGxQtg
Y0gudKQslwD6ZTlKyqpn3U4cjfp+RBykReH+HfzMlBrBQWeals8502EuAOJhKCf+
G872DsFdESsWFSiqEbcMZoyMXTAXhZsImhinSwdOxTpP36CNUCqqQCW/TiZCCVP8
oZDkW2+8cwgoyarmV6GiN1AwKoAoGVRYr99GjYGfpJBbwWRyOVV3CPOiVd0yGnY2
EW+Wa5NVZaX2W1OnK/o2opNPZXH7LleLa2dqN1Ogkmmn1HF4v+shjWe2X5vaK7uB
26i+cPvsRieT4jASGAQwlaGQ+yD2gDB63yZ5ZU4mK+3BQxIEHNGXCUUXuoJu+AuY
GT0eHOrKaQO22V/RfWoJmugZBNmuynhPTk99dlvPXE+YoJDUqa73gTAChdH2Zu03
9AQWCi//hvI7aidF0CAiNO8U2OxUFGq7ndr+FD+3Mcmb6XIPNs7ePqlwmcJEwKAK
JBgF2anHJ4E/gmcvT7Mu9yuou/odujXs5xem3R4SRkt+qdZLjqzLYRZPpQSzMnDf
Cvb6Dn4rx7+wViHBLcaCYE4AxNF/gMKkYF4wd/eCRbqoQFl7uPizn3uE5I5hQUqM
t8gmzgHst36LUuIyHa69UdzpNT2BzpsdGuvoQjjSLoRWPCrAMr+q/I0mOYqyAz59
4y/d5MPbdY3RD1r7IjHwsEvF2xu9zxQCbynyctT3c+nL/OBA4gfbbIqkDWj3OwEr
rtEfX9hWCnixrN3+4tIggwq7qsU7LSXX9hOhWmTXGvgGLf9Pu3o0/a+THkgYpuds
JHnlbCseHvp5HjQNc/xHJ3D+MI54+x2AevnB6tkW7Zk3eIrrkn6tlYSHPlvFnMK5
M2ENdt9rVz+qeCJBkBxfNv7HqIPQZgQMyL1hJD29zXI4+auujcqBF6qo7QdspBaL
nGoSa/iujfntrOC1xBS2FBOkOlc+zUoRGBWY69ujwnzeEhdg+ICoc/rOv7x3wjbD
MDXM2wIi3i9tWfkDER9xgSIF8W2ACV3kgMkom6dqSX3anJXjsEfx5K5IZ6kN/lsY
wu/gL7rc1AEOQSjk1NG/A5Cx90F8q4vdk+/svgPeEgzRuhGtlPKRHZl9I4KGB/Vz
aB+8lNWEkUKu6dudIc6M4rb8IDEfDDNAZ+zIDdfvHnptQFZ4KrSGO2rSwThfbI/m
fW9jHEMBxCgO8H1jHxhCdJWN9g2rA2Y1dR4P2PCuN0/I4FwnjVqZ1jxaQXAdgNjp
H5bFwJxOqKxH9U7H2lMnKPO+Gpk0QEAoVhNsVuNXf/lVvgc3ag5jUMNt5QCKSMJI
GZdrGZspJKz18F5bptiE/Nos7SrTRHz2YRqp7gOg2J15PK2FIizPJIa9U4a3DBNd
J0hTD90mdU5DBlIOvxAonxtwu2Fjk7y/p//WLkQESrSJv0i8oawmzfLx0zTUlHrq
878YtIKOvxok3mGuILnhcg==
`protect END_PROTECTED
