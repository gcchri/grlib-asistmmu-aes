`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V15mfQrIB/Z93ivqWDnvHT46JhgIOh48t8V9HM2yIJVF6EwpEehvr+efw2K80jm4
aolJec0feJ9TIPEq12zWCfw7rq5sF//8CuPi/zUwD2WcU1B8XyZpogG7HDKGdSCC
ImHXgmzv3Tqss+OnjflQdibimYyG6HfMof8sKSchhfug1iPs9KkujimmbBhe+gwQ
gAaftVkxw9xJRSk280uqZaJtNQwgqp3T+Q+ocNtAcokY3QOsVThOQP3Kia2YssJo
xfarIKug5WcC7rmKKVFCFDIR4k8cu5C2jMmcbKWDGAB06oRRUGVKBvhW1b+eJQna
VYeuIh/cKPI9+OFgO6aOHd2FPeUsKVjHnxF8usX7gYIz9uwjCh1GYupRpRUyzOJM
lPJKzPBl5Wu1L2tvXUH+v94ZNYai6hgl9zXxT4oJ6jga7MvZt9tmZwb5Qwo2+W1A
jxCFoKw6QafDmrpuZ2i38fOTFwKTwfpY6JMpE/bQ3TIphAtwpWaq7k82w1lctOCo
FyMiiHxXrAgPjmHztjQn818gXFFn9j6mMngccc6bGZqqe+z2EU/ic7o8dOWAXogI
jLCPvXzhi3AGPoaPnUHfy4o88c5sMIF9iaWCWWlLr9ny2DlurGSXWFGYu0IhUqvB
jz+udj/eC6q3jXluIUb0wkBEUT1nr8fPdhIvsk1R49tMsC3HOSyRH43Ief0oHHzJ
pKfxtZ3dr/VDwxsitUQo23Bv2ZpKQB3ClO2qkjYFLlO0HwpGmzt2YR/kwv4p9oCw
60sS+B8h/yyxg7GtUElZ/+mnIkVOtbUAqittzfJ96//vw1i5cpqL5mVwHYqtRBia
GWsVW6cuf9RKBLZUy8xdmlhtIIMe857RrHYePB0DIbzea8NuSYKr8HNt1UuVD2i9
F8IfyhuMNlcyWWria2aLOw==
`protect END_PROTECTED
