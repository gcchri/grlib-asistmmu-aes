`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pOT2AXE0ArfzNbDgzszficy9xCzVVB+8QB3eyf3aYip9SrgPz/M6Wgagq14alT8q
M57Nf8GATg+OfaogHn/4oGuTRVxTmOHe8mTIGY8VAHxp2+TfDnF4usD4euRMZW4x
02H4QK6hTgc/PLJ1TydBAqBYdbEWDLtagacWEfIH6UFMMOGM69jp9O/zGvUzextZ
Ppatg3eIZ/iPbkNQo6czn/ImKZDvc+KWE0qjVg5QvF1+jo0/bCzrjCfC1dg0yBAJ
N7eQT68PLS0rSNe/prGYbUaI0LbqJ0Mop4fDGLmlNxGs2qonAlUR8om8GtTvXeMQ
2S3O85UoUHlMTESJpUKo/3ndNCHSjO+jBdHMmjJbRZx+q4mTHgrmuaZyK/eMX7tY
QNL0qVxogloeeDn4XMwEpwwaJnpf81nsSL9MFEopxuL+OrBES9oNcQyUogzr//Lv
WjXxOMQF20whI2BdOjK/99P9xKT5NmXNrNhzZEnMTMvogxZ5n+is9Ro2GlpF5RE3
ajO8K6oDGAL4nukbN+CL6GsEL+7hJLW9fV89GciYxt1PDCfOX+J0xSHb6Jmcab8l
VL4u19/isTgtAF8BmBNeH5mTO+7F/OLsYJBSiYEIqyXJIrdkRQqVwGuy/A3rPjPZ
681xgIUQoKkqfgRJ//F7zfTC1d0xOEtBaP7x36tih9LaPFRhxevmg+TpyhNXG2vk
`protect END_PROTECTED
