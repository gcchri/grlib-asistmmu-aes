`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fv2xmPgQxhQyq3nx79B7GxYvGxoMIRcbzsoI9lififiaWYPI/2/aZD6oW6PJcOaU
JNI+6pge39PrEBDMmrRfSVVnnuEOq7t6aLhuj1eee2lKWbxujFuLYRMNNq7be6Eq
FWaioyYXzUh10shM+9YFW3ErSKn4vlhuokG7oUcPOoPEkJ1Yv7fmq58Cpn92HXh8
G258B39dw06kkcnaMjJ5v2ZUXDSE55SMRaw+eNING6fi88jVVXrCOLFf9SV1ZGf3
DNRDiBNGJkTH3dqcQfrkhiuwUQQdV8W7DzVUvQjI2Pmerp+kmYebMlawvWqO9k7x
j6VjBdnnBqoUilC8yeFGKk706RVSDr5bQs7FsJd6PnJj+Lv2vcj53bacqRhoLmXb
yAyykCXdofdHKF0BoZgDF7WqbwGO7DCQvWcPJ5nT+iYNL3DLFto7MtFk0HD/KjhB
dwvq3xk4p2bEYuZ47UjzlBfUKybIcnVxwnKBYF4bwshI1dsLBkd1onoRmDEDaIvo
2Mj8zjfC1iY7lwBH/UIpNB/oPFqy82op/icluDAhtoiUd1DcSB49mLoU2AwNefYb
yCTFMJVBD2pglIslEKPEl2QBkmg/iKJGO+w5pXjsnxEDV7Td+8EL4kRdNF8XHNTL
Q760zAQdpx9w69Gp3i2c/Z15M2rRM0S59EkSDVQxIkeaKZmBljs4btZ/B8excZ3A
Dqw0Qti0UCzOi5ZPW3r8JTxiVmfoeyPCi298R77wIrJeN2I8dgAu+jVGqgGcB3Eo
g+zxgafXabS66Sw9YqFKMrFd/dGMxwcuWLgRNNsEJwoohck11tdA1fyZqo8wau6z
7JTmfZpgB+bSDNdAKbdIydTAVGcfLjrftsUnBCas4uFG9M+X5DPWlh8m7c8Cm2oJ
SjQvSzQhrHq243xv+J5t0Yu1qUT2nbhrG03Ec1vhtR1rygNHGQCv3Hmiucx/8SXH
n1DaZ/6TMC6ETJBJ73ghdFMmbxS6yzVf2iLgwt7ZObqIJdHQg9yh0TSHiNLuhkyF
2pBHKlkgJoc5a1admaTd2DjAabqoaDND2bW6DDwldieIXwG2eGXgrUieewduOHfY
4Vlq6H780HOCc82+qiQU9sZnuAg6o3B2k7eUFA6a1W5JkCGejktt8dU/OSwqSrKA
K3a5aDAlrQEpQc/BtczSIPS47W1N6CjRL3KIvHx/xffW180/Ck/edtNUReCUmiaJ
OnzKVER/IkWxgiN99qdz+quBSOHN+eXKRvSeea6K5JZrUQg1WUc3KxK0ljDHpNK4
JqGXw2HsBKboiNs4Xn7RX7UNeHC4PkfjqdkdtBP+5gPXb59oRA/QFl8AkJXjN0gM
w1Xe9ndS6N5JcqZJG6dxIE4kVkShBlho8WMHELhVII2Tu6JQPOtBKRNTwfdtDx/X
zOjSAdaxspxGM3wEgsL4EUiKtU699Drvl/3JVXbvVyc8nZkPQY6FIR/CGYXfVOmU
3s29Gq0AWWuwxkrgLTT06MvFnVsuFqlGIPgkRhkLtEDDQpiz54ySnoygyRC1iCht
8jVrsjwg+Tex0xKksB3N8Rvpoam9Be0METHCKaQ/7Of9u6719HdcT3+9EJoQmDQH
jJlVMzllEvW6oE2GUkVwl+zHGlUT5xWnMwXrrRZdNUcWlny+h3P71LuvKtiP9OpN
KZTkn48FPtlVTAjaOpm8kJz74ov8u+0QUxOiAskVwdd+lgGblzIESozwXA57rFPz
PTwLi/izLNTuiAz8qee5N7ftxX2prk113VDy9M15FEd7SxHUnQZ27+BzaRvG38bH
Wupc7cDMU8ttD0rAKLh9FvZs1HjG/8NtgOBjBw3RQ4pVmvQ5J0GrgAKmws7xgE6Y
psRVnFZleL/DXaYyfOnZoqiKXKyrzbi5AHUnk9SjTHhL1UXOvAqiyWk8PtUZ6Qwr
A/+NUqif5Z5JW7kqAnJ6TGHrVB85bZBd5phvnU/rqkUlqj3rTb5iiu4Q78vGaJ/d
117MIyn3ak1i0APToDMUMxNbU05JqkQ2lmtmu0To06QeAIVdkkcL+9eJBVueqVX3
6JoE9uPVrJsK8ZJYLTDL0ZLdJraags+9uQVr8vMt+uyXtHJbnj97XoqBF4oILM5w
Tpgn4MsYds9MpMroag3SifaclDDt1+unrhGseldk7fsGTE5tdfuRcSHJ/Dhd30Ve
YuCieE6S/XxOSQgK2TwD1BMcgo/u/YID4R+HUfmNgdHycEkOXNkNgSs68Uk/v0Ja
wojaQ5Ujy0pTm4Wu6RXkEaC3Ge6O1kW1pzeuVpf/HcTCKI1bttyu9wmdHgZOVOZp
M4dC9VFKdk1Wm+sLW4T+T2Gub/ss0XlkbFac8oBV44OalktOV6yYnqW/MqlRl5rt
DPqxYFE2+/2E8h7uAJ1doxLTvytx2HZqUli/Sfal/IV5YLAjXaJ5/YoOFmOk1EES
HcU0UvwVa5AGRaV7vp+poaa9ehoZDsVSzWnPPcgzwhFQ4aqx6GYYBv7oYucHS8+p
8zqhTfcmNlSQZNERXPYsxblutMcdJLX7yZdQx7Y+R9Oz2YtXMGNGWBDVV1Ltgzzt
xEgF63apCx60Kfy/fD5e31rnvsNSFiFwfZAL4nWX90YlmhhEfh2FqDoGNytnIKCo
WwR466IXkP14KSBAbPGMTHHYi7owMpAOqj/5fU9ikILI+5k7dgbE1nEj09SUo2r3
LhnNQKsVqzCpzQktu1qQNfzT7A11VYBmtNvIkI87UX8XGMJyFON+fsu8CoWO0hPU
Cm7TC34ZfdTZhZ9Dk0xRuIvJIcnCI2rtkHwBER7iayciYZqgE8z2NPmIu7DLqQy6
X4kHO/DX5coP24loI2oxcj9mFFBzKD+evyDyDKtICECQcDHgfXFawYFD0EHq4cjv
BgP/UCXiyMysPxxgP++eA5QYmSy4+rsx+7zOuWd063dd6Lvma4WnRxy2SErRtPae
mI9sEHOwUFI1qz7vf3NmY/7HIlcHnahNRUsfJI7y+q5k2rKc3ikTlueM0waq/9DK
X7qfTx6K6ACjDASSjaoGylxCEVXzV3CdEfKUDeoC4aXEz41XrK2rkxFIVbrVzgvP
DhCZHAwODWLJAtzdCQL50pgmfMSKMvRLzV4aN35LNO9QcGEdIByQas8a1WLxE6i5
1ppKGw58HfTTtLBfHX4ICpJrZisOn846hDrGFBmqZbm2BVhCFL/7Hb9arfSZ4YPo
jykMAa9SyHHXC0nKsqD6Ke9qh9CcHyF0ZY4YB8k76AExN3fEsGQ/R9nWLg3XT/iC
Xfu+kmclztkA5xO6u5Nnfhb4+E3rXzfMqRvGTNDnMsWGM5Ap3U/7ezlcQ0syq7zI
R+5hKyB+fJv30GgnpwKzdhLdLW+EBBwAaeNWMQwhWU3gXoTCTClzFFzkZC76Lv0V
8zzbTz0Z5LKWbCPZBxj4oIvmz2VwnNZXYWCQezCrRL8i15b9wYmGkQt9CEbQhyni
h1cOXdZHeLHqD6awUtj92myECN2n7RXyr+iSB6zd/EtE3InjfLMEV9zE0ogAxgaI
09yTHNwhSqpDoqCnLWVPmW42ZPJZgEeldRg/UiKYU3vmFfuWs+Lcbpa3oZq2MC0t
ylGtJK2wYQbQdQgKLXGbJ+yDayamuMktwSZfqbJn5QWvGCDP6ByPl3kKKOzXrL79
IOlLI473YvBFoh6owyfYuD8fpIU4rd4ALr/gPskvSJnDnoDCy4KghAHJRh6viTIe
2R0g3EVqfOMuPWiq2lHfjBw8QCjx27KgyGC96zbRQvk01tFwEIO5j8vlWzx1H/Oz
EmSVDzKfXBobV4u0qrGmP2M3Hdrs2LmMpt0ZMGKa/S8OTqOYMKKjVw9ZJGOexTHf
48M13uUbNE8QROSMRjaEtfXxcib+BwfKyCVP8s44LBI5PLIouPeX9nRlBOKMF+8q
8UegVpJNuFnGpN+7Bu+9Y4NpL/lLO0mAc7TQnoAWoe754dAJB2u94BAbUzOhq0D5
Vd8uxei9zzbj1F+DFU1aXRbYAx3OBdZgeNPBs8R4OtY96uM40Df/GrFNBJ9o8w96
5CwznmvbAQehrCZpUyk1L9kug3koP7mrR89A+MrVKbFBK9zjQr0HuB/tkI5x9iG3
3oN3Pj+Cn9eg+oLJFTePPjOivyV1Q917I9g71MVunBvENgWsMulY8CLoAt2kScpC
WgdY9FP6xm1pGTONc9pnv/wHcmE/HX8EmzQyHYgec7zaXvPX+sJD5FhzEkUreUIg
snFYPW//Ve66G0zQTR35yXYcQirUXF76JF611GprcNcqWJSV2Fh+6ByVBkWiF2ni
FDvWNtqjdDB1LAiFh4Q5SZ9Rv8800WrR0hE7Sabzm+9mogRWy1y3oIUyCScz6kPS
2l5U83HzCR5seBEdjx7wuV52QqZwmmOvbgMi63wfGWvkBRjDMfmBAE6bMaAG3B5c
NGOR4Hsr0jMzPz7xqxojF9bi0Rfgbq0b9642iPiZiuEHixWUGdhw4HKSxdjjsAEh
fqrbhYyFLwJdcVwaCU5J61q1tpXO12TppLRMEA21zthLRUVrd68dyMw8/DRhkfJw
ut0d73BLOTO+3PqWxqAbs7CYHHsZayaQFAjh59HfrK87V8FV5P3cBtO+1KfcPc6O
sMGUwWGpEeU+YJdiZeDeIFzW/swh660jOYWCTALHsvBbPrXLO1BLA0ntb3ENi4Fw
2RyQ+jEKBQg/nmhxK6cdLZ/X8u2KgrtVlY5Vxv1jo89V+OGhKiDMzrnc1ip6oQkV
`protect END_PROTECTED
