`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6v/1LmfD3bIL2PXmPDfY3HvAeXj8dmFw/nBWQzl2DMx5NROVGe7qTEBlFWya4fCN
PIJ9b6SBfjeNu7U7SYPr7n9Hl/tcib7Y6YEquawG9o0VhhsaJVcKB/Lq/Bu8NnG7
03ngW5E0UqFUpjkQoBMuoLsy5xZPYS1bAWuQQ8ZrhSdsVcgDOqmogF18PLoZQZcJ
rYHAVph0x+IFkSCC+gnkL0/x7u4mYudAcWZi8PJXxW6xPhUlrXvfhuImvT/coPzc
o+3u2DdrD5yCEi1x/fsmS4YCwSWj5I33h2GCLpbfxHBRbOpA4z26NVpESRATHbSK
1QD+Cjqpt4cp/560KM91ooZIIYoFetwM39VdsJE5QuLCtyZlfc2VGjHWW1luQwXM
h0Zby946zYH2JRmsZ82H1IUP9YejUIcaI2NEWXEryA89gHe0RtU/hRBGfgIsOi7Y
2D+CrWXMsEBFwKr1GUUJsIFZWOfiUFh7a1lDPpLFnOO8iZfuyEQLl7fO2J9mnISx
/2WI/ikolVpH0IWb4I6Hcby0VuIayGDQ6HNQI0UlS5uhg7zEyTWsvV3f2vkONCw8
Sp8KpxAYWhS1S7pH3DjyzXwIRU2qKmBXc5rCWWItN5PWMd80Kg9TPeAfzNnx/BIJ
m0S6v4jK/uvmYznJt1uJE6x1M8a9UnyT+PBRFYRAx8oI2oFdapy4rMn0qU1bakQl
g2sakTEmNgd6fxKjSFinGL2nD+uAejf9MGY90ME24qsyxwB7doVawW6fGJxB2ZNL
4yMYUVgXyxqkjtzdF4W+jGVr34EO9yxocNaJ5HSDuX8IL+hBs83mqe9S1m6O3KVj
wsr33bm2LQvxXQQUA2YoKJWS4qImmlWu/8B1lTtsocShwSkmwIQ9bM6ECb+sun5t
g2oQ01G6LBoRtX5BXm5k3+V7SoaFDIvFLOHsXz3qn2C4rdDLlsA4G0V5xXTmUXWe
On55kKY7DwAT2O61ih+4RLM5uO5144qOkfjKE/f4bymN6HGd75uRhYMTdX9ct3Bz
ijFIXw95FLxKO9y8ZermfubMtVrfKARQUpc0Os8gh8Dd25QkRnThAxsR2fhZ7YUD
QavQGPW99Iq7cMgL5LqDYKapHkGfApAq+uOkKuYPiv0=
`protect END_PROTECTED
