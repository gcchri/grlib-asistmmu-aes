`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
06aLKtF535TDd8GZ4lBRBFqU59Mc8qZi8oOe/U4UM5gqUIkaURPXbXdf64/qDch+
y2AOzF8Ju5R9EgEa6a8SwYHG4CUyZC1R7MBdUOLRgm2PKelxBJZbOiWl8dT9nVtV
dO6cDNdWvtNdUOPKspOAqUAYO4BcV02p60hcChTv4k3Y+iZ4NakgY+deSGnzl7WY
Qv2fxiSvxRlmtvxYK4W2/lPViIpCA3mOeVoZtZ2EZroJKaXlLRbY3LXoiuIx1rB5
rjT9IRKjBtM0/St4OzfweDJNLQ1HiKrqiS6IZD1h0gsMS44Yoo/E9uO7Tp5Z1/YF
ak6QGAj0dlDlSFmyXDjDueEFZsDTIaXjxBBJ6TcLVyIbHu1uZ0tAgY6Mubufyubb
32Pl95xi9jTDZe1DsPFZjOmCtWYmEetVIINN5gqQvbJl224PtGruSswNxJ7/iDKh
8Q6cZUBwWzYK1IVMrf1Jx0pJhJ4i4q+bgxicUguXiyAklaVxKSWDo6tVCjCchuzK
6jJRl/mv0jHrWyrBAlTMxLH0/ZqSHgQ0aR/wQZvWDez9rYAxYmnmZTb4RT4JBAuR
cGXhB0DL/c6FmsWiLpsJUiho+pxO7x0Wk/NIWvh7jkxskzKFvTNhot03wImkW1Ob
9WSLcRvuu7yvFOOMJwOvMwThWcsOCJa50GY1zkSLDRZA1wg4jKs2yFr8KOjkVcxD
TY+Ot6qUwavbgI2T0zVYnu6OdV0de0aJNMv58HwAxG5ax97Dup3p+LsvmQ16Q4Zr
GGyUhQToTlTz8C4mB/n/ryi7UMKpeODSkkSiX4u9RWwT/Vf8KJXq1LXp7IbEPD21
2zMeaGn1UpJsz1OIkxSWU2Kn4S7cbrTzw8iQVGZMjDJx/xoukWKlG1pwd/zdC6h0
hF8hVeNgIa92C0AyyoP2I4JqBI16odjJnAcYaI+1vrByGqU65l/TPaMWx4nWyo1V
86VdW4xIR+D4LT06Yz3ZninWRxWYKj++UobJTurS0Sf9I/3HgE7e1GSQzfJ6GeBR
euPuuNN9jckdLXCTBkgfviu0VBD6YFSEUviffP8l2/ho6nfuHg5++9nnQ9YS1/m4
UayyvGAO5odMjGpglQ7LfzWxuXL+942vVozihGFxRT501v8CmI91zPGsc4Jw1Baf
0yhViWYDQLFY2vQKvZO5lBuoywsCUhGsar8WS5c2nuR1pGjX1uRe7r0Wida1fhaT
5QoduFb0VoDK88SlSiL2HWo2uvIBYQ6+NGaaaEQ4uUIrW3LRHiL07dyemCaQ4YJI
`protect END_PROTECTED
