`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BhSzE/a6GxHNDUkwTazW+DXqNssVu/qZCY0OjeeRGDCiYeII5IXUxYE/eTr46Kle
em9jbPw+/B2XVSE8Kyk6/FxRGVaJ9s0Nme8L5tyZgdIdWYi/VP9KrfRmCez6US1a
smNSvk3vDdLK8u7WgUqH6b6AKpL0nT9rPzxvGM84f9plV+tmXa1vHyGgHnxxOcc1
5ugu9UacDARKmjDtKZiQSJ4GRIG1URrVATt+DSRYu4euV8/1KJiuelGAjK6ByoMT
izHwFFHFieMN03Dr2EK9T+mHC9XbVQGwLd1OHaPaBnyMaVjvKGobMTRokwprZyVr
vf1iapjlHFWaIpLBYCIbUpAkwiZH7Vr2EtQ+Fy4UrpExXdjJrTjRladzmTl76RqT
AxMI+8AkglEvgd3F7hXdYSmFvB3vETMbwZOSxVjR0SwErvuhCo/NNaAloW8x4ajH
d9OuFStvB3EMUeoRdQ0WiN58r8zeB4YRbwkcWzEm/RiDPHHM7QXES8cYOpgXvCZB
STgORFirg/K0azi7AA60G4PeJFAKk4lESkboWQJaVkYmqtnpeYtxOsQtpsym3XvW
pJFc5CJlHD//kR3A8Gfk2LmnJ/fF1m+Zqp4/C6QzFoY55g8+EMImG5Lb086gKaH2
CXu+R8l9yCn0hTbJAKyV8kvomsWAlSj+fEU7tN6f0SK4tyu2G7QI0r/pH587t9tR
3G2CcRGjM5Lx3jP9B/cX+Q==
`protect END_PROTECTED
