`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I+rWdzkkbs77m7xJt1lawlE9cHBpM7WDEOG7/Np2Sbd9S5OPdkQYIzxO20r/MJFp
WHs3SiAX0l/Fsd3mwTgqppg/5H23Nc3ks5Th7MMApNvm2XwliiiJCVBMPcWMqTo9
/WX2EbsiIwBZttu6i2NEzEM2a3M3d2pPCu/ljCgw1ILfFLtN6bJSqANpgpI29qlt
cqS1+qWLA4PedWqn7qeXy16BGt4iSYc8qSdDATA6e0t9X/CiWnRm8iOAgEn3RrIV
KuKrRjI7si3WbQyY5cSVuxDiFXrfBZvZ4b+qTW3j/pshIvX+qeBWdwaOZnQyu/5L
qofSFbpr24mEFID/XnYbea7rrznFiCx2/Pk2YWB6FGPnRyR65MWgJ2YPw7Zs4o8/
r5He0ywSNWLIdNSp1Iw60BVMwL5d8EumKjB9az+yulEbvrICidaiOYx7S6vjQUGU
Qom285XFVTpegDyd+PvT/nTMa0VZ9mTv4qjPkHw1j/2XFnUdpZwzy+bZlwkyUdeh
LWPwwQz0rivbokWWBY/xCkEZFiQQ+zZVDwWTeZhN/Xg=
`protect END_PROTECTED
