`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n6y/1DR7C9ypMfboG+1/YaRLlHjISX45jN4bRrOjCg6QACZgcMMOrPJWVbDP862W
At9il1Gy/hGvKgAt8OrTZn0o8OuRiUKeIwJMW6kI6lKAswGSNhnsWHvmU3Y32Jt6
d0zdeSoGTb9uxKpWUvS2tulR81UbLqV5v5eipVgIRaWryMxy05MzbokJEKoUe0gu
lzO/2UzpIupvAGJ3zd/YfcchEoMAv3o3itj12dnLLiinzlrY9V1VRyOxpdF/gSl9
LItOGMktfO5Alm8Bj1/ug0hADpjINgMOQPnC+pa0ObygJMdzTca4KIfwDV5RX+V1
CfqWfeINk5NaoX7PAcxvUmuuT0K5SmiA1QoDWYJDwpNgwFLmsml7vS5tA+Ov2B/E
LlFNhsb9T2UbFkrJHD8oL4Wxsw6O9JMuIG8yko3VdMPffpTTYBGE5EkTvLFWbGY0
Yv5blDKOKx2sA6OPzn/PorzviztzrsQtVHMuY1VnM1NxqU8N0UGgjSGv8zCT7qpm
jfnwPhFR6yUNUYW3ZvZF/nGQYYXWeqigx5JRDc6MKTSbK4vW2EUfplDfzfGjSGus
bkzEPA1k8MtoFHzoiofNVdj3pD5m+SM4/GsoQ1o2dL+zHMhu0nupARgCxqcUhcNP
79IyyJFK6kBFUSPLtJSi7FVM+6qFakQ4MMjyhIIZ65K6chUsaBvj9fgGFvBVrFVt
mK1kdBidJRcoXSyLBIMwT78RmbdIHgaHq9n75uI1yKhfITY0HrzdYM1ATHwCN34F
tnwiZDxeXRiHsj3oonvdXr0RAR957bbYETzQbe+Jg8jCF47FvGXdglWyMYk/4xTs
1DWfBzGl09S0NTdvGhww5jFsugnspjeHAj+FW8J4pz5HAq7PEvi7ZWI9ao+ZY2vo
UYj1yi8YE+QU57CJGjLF/uBncgBwO6SAtW+jRnTiuZnSgnzYmva17D2jIMgwD/E/
QmR3jHCThKuI5nV+zZvXdsJYoBg+TOMUgmh6JfwNDwhH9jW3qvjJ9BSZoXDBdx4x
iMl0kYxUiLA0qQzzBO160HHbLqBerFYLv70gXiFx+EaqvNnMe+RiiJu11nUjJOe4
StxfgsVtPaoMMx4Dq1rew08gpyoFczNdwtPjw807OSNlQKTou5ketcEEqGn+vZN6
SzKHxMKGhIm1Psuva++jdalCXwmudPxGG/m2HPpZoRt/vBQCHBacru/X7L/hwSeA
kktAFl6CHVnJYTaT7SxUOAkDSVwliwrr64tXkz8xvMt8vxxXaTH5ouDdwwh9eCK3
iQL9DMlTLOqtrWdH1x2r5EFfls2OoeYQuMAqpLjJltcnwxrDCrjjYzwUaIoAOC66
pJn+uN2NFRasdi+vD9HZ9sAhiaVJdPezK2CUKcGjPI734vM4oIoL3m9QrVsJ7wXX
orue7QDr5u6c6RrfBrCHvsLYyo9FG0Hy3uVB3yKZKmql8IgEuABsYcQk0Qu72YYt
iyN6gIM2q6BL3RCL0s/l+U1FMO6WZV5uono6Q9P4vhnH0b0Tq2AecfTcGlXF2xQR
q3EDUCtI2OAfjDmOsw/eRt+RrsQDs8Stn44PCCe9rILf/1mZkQ9YORag2UoDxKX+
f/g/G7o+PyZWTT+wnIpfSrH49zH5qtysm3TXeEYTnltP2+wRbtrtKnOD+REBsrsw
6pJhg8qSjvI3fxcqeaOB6UErQgqn3Bpvg/CyHaI4H3nPkc5cEC5PmQomLoAGt57J
/0qkAAU8Few7OaBtBLGVfif1e4A1h5emWmd8xI4/SFiFqE+rfQw1pmG1mKvLJUMM
NfYqXdobhkVz9xATSmU2aT4CIZUOyAUe5yiDkVHSUR+w4eyIBdHOfJSB0pd81E7q
pr+1v0gta6EsNaskFdtUxzoIsLEptAv/dLCRoOYNZnspBLm3Rylvtt5mb3Icl9PH
H1Ktn321jJT5kmrT7GCAG2zKNzhMWhZfztwMBBfyVvqR6xOIcZ1qOE4GrH1F3CGS
mNQzY5fFy5t/xq945P6ZI1BV2NKXQcYjZJPZJyuCvoc8ftZKgg+7F4mljk0UVnSB
wID2ztAYrbPPI2X2mfMhvbEmYhQB9tkCIL+neh1WZwmPQioEZgnJYY/KwGF/geTV
vw7QruRNJ5sGI9YiHCl/Ygj02hWLpQAqAWijkHqsxM+JMSFziP7dZkNxqhrgfqrl
cWcN2WtwhVslmd09l59Uh5qbkIuLLGdTteCyPB9Ev/ev1TVKiitf6f8ikproGXCq
ct4Hv+gkkk/6ydHaJ5A/kaMH+l7+H7nPHa/T9mlvtb/fMJ9KxBOTVYMXaCjmzHZK
dwp92Q1yp91drjnrgorS5OArWsPRYqYiFpYQuedBk2rwKNPC72oCqw4v3O0wDIRk
umOMMnHzBTBAenK0KS07ITR5YtzypQ1vgfmi5hu1aIaw/Be3+J6sEBgU4Hpg2wpK
RUH02jLZWU40EUJQGHewQfBnTKYa3WrIhCGKEGiF5VIPjhssv0ch/HqeOCGCKO3G
LnrPwMvkdfVxe9T0R5sdOaVzJj3qAPo8X9ut+lk4HEgkX4VtWpCUpal2dQHn1hkC
bp10NWTyc4kw52I0vNCotZOKhaQ2POr/zkucfBHRreUlLXe6G39C6ROGPpgaPAzP
CPkTxqHGPV2orWX8Zq0hN4AwciIfEE6AiUVYF4wIN2GFtyJT7AoHBU18sc8wIw49
FiPfbLTGLecwasIX9HtFGYAB4s+SlWdejtYDAoIUUie5BiCG9AmK+vkSwnZr7TCc
RVUglKyXyczIyZUZfE2Qk90B4pBy5BMJrMf7yssNwSLXD+cSBg9gju0ROnRsh5kt
9t+q0I4fP1iB+PnQAu+N6E9YD6qA7LwpjJvHXJaihd3utp3+AAJsczmNV4xLdE3I
7MDjPABpXquDTK+QS8FWC2w371za1EUdlcHZJ50tvIzvVEZH21zud4TyjYA2+eSm
JBcXMa6OMF4j6SJ4pxN8QVh4yOYj3H6ztTAcbT/zLCwULWI+OnYU+I0Jn4ICx/PE
SekFPKzerKpFgAfZoVDAfdmCsqqYNcaL29oie8PQgxcS5QFYEwXtJ0dCbO8IstSw
1jLebMUS00jHDN3FSBvfj41mKzEvtJytcLB4pFVuSVk1TEg36RFsE/SvvLLsz6xy
kCT70hrB9er8K+YoZ4EIaBuD1GZ0HmFpVUBDQeQ3A7nrk5xo2RfOx49gNYLVFNk4
i8IF9g51IWuKGEaaY4+63s87ssGZ7n1qMY9gWT4VOJOgC7eEMpEqOWZdSc+GYZai
WKZpRA3pFxkHr94pN6AXtofNucwdI0tuh25dN4pTDVKGm2AJqN/DRmCnwiw5eqKG
6MYxUcFrqRO6ZU78/gmFWKZ6OVqTHE2LMRJcKctEiGPxoKu/k1YNq4JT0HslUcUc
ORwkZQ8AtD+6GSwUynZYuAgjUlNhriMXDqCgCsGMRcU/crf5z2MqyMfMSvyZPQcJ
eCpYzNiQ3wcibq4jubwULlghcACACHIiYFWN6GtnL0uGbv3E7R0AMevD/Cb2k+dd
n65YS6LCiLu5lzwMPdZYcPXil0kUaqOM819ArFl0UkxYs7Fb3JyqQ6y5pZ7falpW
HWGvhxlR/KyHjjjyBXZO+XP5zrzLMUuOUWTT1Mp4mafYp8NpVVxO2RN7X378rrEL
V0rVh+6iZ4mC3pvrTKdqv1r1hRRJSiMvUczWEPdbgUo/4rUExLH+lm6pTtg8gamL
eOus/cWXh6vKA9qex0JPvWDNU+zEcMqXtS9n5llgJpB1qm5EFyFEfpNGfmpVyhja
XFr4IPy2LQiSjiHk2M1Mdnuru0dC4HPN5/FjfR93yCYvrjZOTaLWcvxN5oGIgIM7
lACXmjir2TfuvLKbJG+ZdfDwuBXPxzTukCsGhynhEHBbUOGtwLrG8C3w3PqotKqe
mus8/G5GlN0LMv+fKL4w9HDBLmXR3ye2Nrg1+ATzsFbPDj6iedKQ5VBHCn0+DyYU
HRyKfSxU15zTihB8wfBDHQLp6baRiXaj87TTmCu4spcGmFwcITvvaCwIg+vhl4NC
yAbK6iBuJxXVW6T4egUqIb36rRxxS9H5ZRaHvTeVUr98PfdQteDKlJDTy5h4+XRX
FVIkTln+ILq/dzIuYIjCqcQcVnHnfcJI4eVoHUvwYKLaOuZgZKtgKUzt6WaHgcBa
uLvRWHyXyO8ncaz2c1HLVaS4UYqHPpDYIewPGCZS5Y+PfAa0yVuBqwmTg/BqVADH
hdr488W/rJ+v7zSkf06fnaIaYWCkzVcMIDLeYJUVRpgYLapFzwZrw+GdpfBTbjsR
EoUk66wyppE+0jYCw1fgE0ewaAvDTyybUv+TnXT/36ptPIJL+7i7dHOg6ACuLv0a
xKoCRuLdZh2oYONoOOFMZ6yUiyX7IcDeTdF8MBpUqqzjvg9W47sZMJuVVy+jlJtM
nL26Ji5oYjkb6D1eJmduynq7ryyD/icgoKDvKuXzh+gKkgYCXKK1DdgsVATFQAAI
obKh17XEf9smPhApiQd5UrGAemh5vPhr4pQP5UUNs73pR7B1H25fa3IYc8Pn9LVR
zemLbcLhLvSvfq2C+R54SVS0IQn7V4W+DWBIJnTwGEOid44WMlgC52vLgcCem5R1
9NEn8dye/rLnykfzEzfvh3aGO3hcDUepnXAYAHogVCuQ/30aXRQsycqnFhK9VypH
A4oaML9JWkZ5EGtlHFu061nhHPe7jazplYEHdfOs/ntcq1H3dGZcO2hLHPi/xVUc
Ry+oifrLa0hWWYyHxibBFd4ex2Bwxm3XeeG99eBgh519YT9d2xzqAjqrBPzSSXWH
t7ZuW2kD4hY0QiPf57yoHQnWellhQuAru8pPpHh4AvKn5Znr0GSOxlOouetkHsyA
u6aJWMojhfaxh6l60DUSzGiDENoqOVRqO/QIMXv1WKPoaTsAomQ87A1dWPWhoKXN
UIFG//ZUJzzAUbiA1d+s3ltDu93GP9jxV6DAYdwX4s/NBN/1QGA5JxEedpMquvOt
06ThFG69xSHT2nt/fCLnIVyexn5Y0a9a6B0hp8gg2YXxoV6aoJVfaZJMam0eXZij
sVj2arqaHcyWrdjy0xcxhSiKbN61kxM3AT+nWKvln+lm80I62NnZFebEKKpKAuoE
TpaNIBjaiAKdW7ZfEnp8arGbyRWuBlnxFQX+MdRrcLv4mXzCjrmy00TP6cGwbMfR
5ga8y5YjRx3bOr5/K47DaqWmHfBiSOv/IfnvjoU6MHrFrCSbVYbckacG3l/khc7A
hYlcK9VDp9mlpuuahGsPPX1Q7S9yAsU3njkCmyCDBK/m3Oi+ID2AThFj/d19kcoB
gHJp9BVwrY3nZC/4E/cOFNBAJ2SAaC6DdinV0T4wnfVxIRW5I7fLwmuSbLoB8z1b
WH2BnfDhxobNWMMxxo9a6z4WmU+k79fTYmPi1y4nd1l3Xu0wQrZ1Wz/oklfFIitJ
swH/Wvq4FgRoMcCQXMOS+wfohytamyrHdGI5bQdddN05kR4FyNLGJH/IJwsZzkfj
Tw4iM5UN0T+VNSxyhsV3gGbsREc5mI9gfuEtYCvHnY61kasyAvRT2jMOoMO529vM
TCIRshly3UXqjlcLEZoLvAlD3dVZN9jUdyh7Zq/gqV3cmJBjcNuN00c6cYEDa2/M
PV7yudLtAkHSASQ427hw5shOvs/5sv9DnNwdtaHXzw0nYMoZaoUcnbpU1VQVrNzs
8AAGmOeb24Uspqn+GaFlEytvZ1seSI8VJw5SqMCxT7ogeIbW2wGt5qSSJKuDLO83
l3GO+VNsVbAYpQCR/2Pw7eVWWx85F66TvsAfZvh3p3FWqBNCSUUemEgrHBzwtPG2
uFUVnzGePEP4pYDLtblZOEOxdKGWnB5ElMW2Ety9vxgAaZVizR/nf8WqRb+iRoqP
hLUsULhLiUnewZqj4PKhhCDzEeysoKPOyaw2esf8sRXZT2YqIj99kvdsQEdWDM8S
JuiPt/8nV0ZfKOpNghJdy5MMGQtyCJDdy49Z79c5D52FFI37sHSHFbBAY+ipc5iS
fjGnhoSZsOeieEt5LcjKnsmyb/5sOf/t3zZvFRY4M63kRLUfhBwMkjezg1Iee242
wYxKxG9+L+/wwy5Puxxzm2iMHLy1cFLU4mb5KA2Nm928w3oFZcfDPZr8eCkoJ68D
B2zocXTKnyIST1xdwec2x+2Dn3/7fEA6ijCxciDW8pKVdCv/HhN6hCD6rxkyrgyP
CZAEfi8FpV0MFWQBrV92uPUQj7R4KPZlmSgQ3qijkQDXriAn9vp8Yder9Ku/StvO
3WZY4ZU6r4ujq28gIBIOyckmSarIScVpVbtUDVpTjqF758LkvxQSO5JXaHepM73p
dKlKZcEgKyq6ODmZ7WZ4kBBWPpB05Mi/+WAvSmS1QlxcDArAzeWVE5AVJ9AW83XT
JQp+RObOg4YD398VGwD1S/W1o4fnHMS9YFzNdwnR9W7U3HKQ2ftosarL6jRKZujN
ZsUSnw5lYWrbqhaw3RNo+2M4FR0e/gUYRt8hpaszP5AfPfGk0VPjzC4zxAYEuzcR
bYW3H3+n/x+AT8TQZ/nAR5t9EnVYvv/uKIItpJWDWMYoQXO6BXBDcrLFX5FCu0oa
UVKpwFZGDgYf6lb9YgyeBNpZHoeY9Cp8RZDZh9tTO/Guisz+87Pmsp0QiC7S4plu
nC1EGVD5fO36Cdk9a5cz7x0UT2s0KreH+G0RNrLzCKbCGIlARdqRDirneg/LSazQ
qrDpbcv/43jlRSsPKN9eqSoDSNoDLxP62nOVbymgg9GF3CaRkSW3Gft3DTmzsC9m
EC48kA1vyLaIj4KYWQMbeIvE7r+euIhLtENyJizBt8fa2tCDVyTxN9sKjwGl1N8P
BwalSGDPVqaCFgOlls5Q7+ulnOh/oRdKgunFL5dMqNbDTyq1YOEcbgt4XIaboGtH
oET7qmmJmFLPTtanfbbiZ24EZDBJ2Z7eM1i3tTaOHEMeIxGmUTjn90ZM/cOP3chn
UoyVLfS22rKu+5IgD+wXumPw2Z9p7EmHsdG8B0re5i3RyQvMyvFg4ilUTOR3bVOU
QFmWto9tQhLVW0RxcSW1l+Ne3ldAUklfnXHKC71o+tmB9EVrAftRmNTTX3RescSQ
ZQENDMAqbtBDJ9gRG3ZA8587hBy/WhheVDiJWVUoyH3DvXEv9I73m0tK7ne7Aqdo
fN9fAud+7AHnqZu+Uc1X9Z+b2YJMit76M9YLyFxsCMHppE9ij3FP6QoQ3WGonSBL
20M4KwnvuJ5/SmCeu+KHQXZZLK9INo5TIthD6tBzOBxw64CHb7wKmK3xxchIWUQy
EQyvFAK5hRfNYiciwp8Wn+c86FcSL6h5phkLESEmyIHMYSl9d/PEimzbyr/RCXFd
vWlzY1MMZY7woG9NmhJfJduZskGRMvS0s4sbHOCl16NiqzzJIBkUpWixdDm56snD
FvhqMksXS+aL0b/S8f5jXcIFg2WmnwOnTqmQkqNfdohH6HciKcH4kggBkRouWBpl
i9hTD/Te6X+qX++WvRhRz7M2xT9scX8waqyIPgZ15nHcif6lBA2b4YGXCYHgoE2Q
JpYIXj+CYhX+buIsIyETQeeDlvMDCn0YIUdADC66GbuTylH9n4aOsXvpu1QQc7js
Q1FpF8TmEW74keTdZipmCdIRoSgJIWDQKhbCnv2bZrQnNVhsZF1Aft7Qcpxp0Ugw
wAZF5RAuknZI0y4P/OB7WSIhpMFDoecpuDJ6QEq7ud59n+hSjBmqDQcAZt6ldmfc
G9fOyvYaNNn5qWxo5IfwQ8V03PJAIXs7dnfCtSlAku2hCAHw+BdwoWDntHiEsBxo
x8tiu+0uISRubeF5jI+hHi6rEK6/W6g+w5KU03CsdU7rIlJY3TEoCX9wNn+OtdGo
l72DEy0mpReoCN/e4YxKPAP3QpNm7jTXEBfI0s9KC8bxWVqrSZt5LDP+UAoDiCs4
6BHmw0ivV4AXxwx3E7jLZCE2G21n6NVMTGVEvUlu/4HSU/rQRcWRacsq2hew8SRA
CGiWHraHuQfuw+cmafVa/5WnZE+WBEbeNYLnlykxRmOheiYRQXeVjrFTaB+XRsC/
Kj9bZKiKp6bPZNi2NgIbQMgGER893iulBsUXjhLZgH34rD04VA3UwsQqLXnpAu8q
SldpxJskAfk6gbOn5Z28VrlI/loOskEBMuMPhmRK0O9iJdjdHs+d2YSuyuYtDqHx
HWFYPuXqE+kNq6InJ2ZX2WU8Hb1hI8NGSoPk4lnzO+F3jQ3kglCAk/laAvWVFjLF
qb79oeOyMOI2kwNANw714/ttQZy3MuNq0WFu63R48hk4y41Mx9QTExRhDvI6YUKp
abBQbX+ZUTjoaYcOsRnmehREkNs/rGRlrusb/5A1pa9vCbaJqP3Xs8mAh05mlZEx
4gsPwxk/jyIZXwxLL5oGepVh2Et8wIgkJ5knPwdZwCF9sKycWx+fHL26VVIwPEhW
9ExYWqPs0LbGrkbK12/khH6hcDPpnoTrNyeSN1gD1w7HB6XkNkDv76GczZMxWBxn
Nr+RuoHOOMeZI45RjrsvuJ3Iuh2amEPk+La0sy9DBZTBLEieC45GswVBOU0dGtpX
Tf1cR+ygXhVRKqUF80W29yU1j3HZlrc6Krfaw/0esM8V6ZjQ4KX/Zcgix3cEN7WH
+QMe66x1M7fKmttI/+Ue4MzsN1+onPFESwi0RoOvnEOE05YhftimF2abkppOWQgb
jFfcUJbxBGMjQQOBQbv/vLdtTrrOCGWGcRE/AFHbZ5/73BxtqkhIygkQLMikmQpl
IDrwXfUZ0ESLQJv+yBEh0tDbThCRt/Sqxpq/hHCkb2Heko3/qaENf+VCvvqlvD+Z
AXp32JBfCOJAwiOrU0on819F1zoA6koaniWFVDKvlkNtplAXIfRZdvAW75Ix4pxh
l5FNJaK86VN6Kz39tE9HI1+cuKR0sUWdoKVDNPA8iW0+mPVo8zr8egEYarvvNX0S
r0GeRWB6mrBogdDs76TLvKDYTKmtR8IjUkjjTaPWMKDnAAOCEHTJo/ZgErktlfOB
6E6APEB9U+oO0OydEncwLnraC4VzY1MB+gmLVRpRkWAhhYiuNfpidtuzmPBoRjTd
nnWB6PoW4VCEYZYkvlEJwjiLFaFJ+ELqPZEZqLyPHsmPyNLw7JHgYjgsWt7SZudu
t9hxzQnXGRI2pGNq4YWIurzVXE3p7w0zhyvBF2Kn23qJspjMkag5b7afq8pvnD/G
cJmh4MbVlby6f+NV+xHRcGsHQUjBctUTQo11S5BXgLXMzb7Kmvjuy36cUGP/oRRE
9AnIvRjvlAW+mmzXWma+tN8h0bWLObqh0dmTcCocN3A5soiLPj7E4sOTzWDV7QHa
kdlK0zWBWBOMtxrMmizxZq7PFXKGlulKGlt0M+w3w2Uf55glyYmRWJhUNZ7MuPsi
IsWgV2cXJNWrMPb71OCPabwexG2LDqvoMiAjVSVH8t95oW8uSq/7O0SONG6mFxZ6
NuQxKX/bXloZ445TGsAV8vh42j5fMXbjCW2qP8trzLLMbGarxVbSFH7jx+cTxT+o
I/7Z9Oxp1nbHsX9GOUoifIh/EOFPIddd8gRrS3tEjTjYrGfLnVX9fTaPO4U8082c
dU9hN/yr10mK6wv4DtSWpRzKh4TvvfDEOeOOKO+V/n0ZTfQz9wbSUWw2n4sIRlXD
G0MuiGRW4qjy8mHCFswXYafmZA/hzKzD6JY2JtjQjfK0RQDLFuyTtmKZKgd9N+sr
g6seUUJAv4EFM+ccUmkLVIHP7mPTaNU2hPZfZUa+BO6UNuMZxV0eTBvBRGotELQ5
Url9mjuOf4qI/yLeLGZgE9NVMo/oQGxtRtQEcIT4CcmpUj574GQJrgA0D1XfR81P
aizeJzv8ekqVVelRMY7e0xRRzk1HaY+5PAer2OvofLjqBnaXIquFqNxEBSNk5pkO
XacTJzOaHqPn7yCiE0Ljzo75K8Qoos9Wh6MLurw4Z0SHcRFPm2h85qxoXNPaQWjq
FC1uQvIsS96JcCta9mvqKoTOwg1Jg4bHh6rZsen0PVTR18QPEHDkVrCbb/XUvRdj
f+OhQ++UG3B6cT05jNTsfOR75fEKZ4RRm626xaSI/k+ihWYHD4FpX/evSYmaV3gr
8Cn8OKKfS/lZ7ZUx/2xlnThlMzYyxiikyYMNg8ltgmlUoIloP78P0tf+qc3awaAh
OEzWiWFCYjeNNBCpvkalZmwZKCAJWaNJiPgCJjeHhpdozg3MrvEoReblOn0h7Um5
mGhK2Ozn7ONVcEDBXO+PNUumM9NXkdrr3+oH9uDLxGlstU1lGhNGbc8uBeT+SZN4
sWX5fGv3sMsaWt0t+HCiRve7syBO45/oVPApdfPGZnVCkbgknxSM0pMNUjbxecsa
EJ39f40mDTcvFjAgX5iVEScZINrlMVgEVhr6+x48hn8H90i6jZgYfPBxeo0EYLE2
NCVxwCBtMaTHTNcetOM1kincV8vtMb+U7HILmYeHdxtlOGuGzu7IBdSzmxCJaU8g
nqBwL7ioj7o9QXDXmxGxZDT0vlPBLNJbM/f2AEP6VxD40Gt1qvqbn792W6jgXX8+
DIc7UL+cEAoJqmr5PNanb4U2gSIDCr1sLhig4BvIQsN9AU8/zpwgV1iRYOIiKgG1
OJNMDiQ5OjfetNintBi2HMwm2xN3KMB84teNSGuQGEGsWqWMletTUfYZmCjijBEA
XKixx7EwqShKeeJQvyTQfe6bBMY+eA2yjuH4Q+LyoSZpuhMlIsFbDN3Mv9RYbB3/
fOOgjHTBsqaOAn1ox5Tmd6JEjhdp6uuhJQnjf8jGGEoBCm9BKFittSZ7snMoPGip
eOdEJ28HUmvkgmQkX/4q3b21H/j+DcNiRdBbUpOYhTTSu5PE93Y5GTauDybu2DZk
SxNcCCUPL5dZtJgkDKQTHfUTb6WjLW152Z1w/3MvwZiaGRCD+B7PDqhQuT1KKe2j
HJyLU76udg2aY17J994uem2cv5+ejPbTh5nH2ZaZZQ/hYNtIZGqU1cAEO4mqrfqF
rJUhVSd4i93jNf0ZpBTF+6epwTxhQ/6uJ+2FiHo3EFFEmntqvZFAoiBczKezfUY/
x2QuCe3w+jUzg9LLkY6xpy1eXuH0AOOaJz8pAer28ls7BZyEXLTieXNiy/zsJrjO
yqEAiB5J0EigMfeEZ4AWna1jFVG08F+0GMki2Rcq9k6HM/1WU2Kum472bPO5lTUb
y0KORLSJ2FXJf4UDvUv966VqeKq9n+wVL/uZB63EhfiHjk7hNPSzqsmnlSLWKEyM
Ht0mcT7Gct4/yuNVjQut5YNBwckA/6wJMm04YdLepDOiq7g7/ogy1cXQ2eiMb7bA
S0amktikjOrCb/e6W5sjdpkByuiphCo2GrbMQ72/lm60WlS9TqTNg3iSUaxfqxK+
7Oh3gGAJy5c7Fe2ZckE2rDbsWkc+7Wh2EHVl0G9tIWbtTlEywGv+O2oj93YHrfQ0
H1QYRH85G435gFhgq+/Zsvd22E3j5fKDXdPCO8EtQvspusd+EVVIcmP4OFz2F540
SFoLOLiKhE9hVPul3wfdMLS+diOW+dEbqe6YLVpzvpFxJG/K6PX1aBPRayAuFpH6
CpU/iOH19btKcFMwPFF7aCcrME6+bWQLxR1QOWV+fEomJgSYkJnUVSCYLdf4Zr6j
KMTc3nMh4NH1bjr/BCuwX9SCqpipRFnKvYcRtpBoMkWlQCv1eTbEtEcs92Uwe+EU
98EWu2pnVU11EP9S3Z9jSaihHQAjKok3qWQUIylfF9GvhE8k1cFA2OGD/IlXMz/v
+1ML+5HnS6eEuC3exjbN1FSbeNgzJ+ApMDArhFp94xg0ZToqDEMhB1bC4zf2D6tb
IsLRTNS/5WL8J1/UXxbyIxMOxJZRFemquIiSKzo8jEMJxfyC+ur3ESnP3PIj/sBg
g8oS5Q82e5ybXm7PyjmMg/VoGajdhYl43eF/lSztLarESXQ6M0ueYYUwOxCqVGe/
lBvkB6jzywc+PWuYcC+gNjeY4IOA9XKrzcq9/gOL5gTooBA49YHwuRu/6SwWKz27
e896SNNU3ARuT2iHW3ugZVW/tKDvUuoPXyiGXa5ELtEF8y6cQ58FU/ZJ/44AV2sn
Ziyf3vyuZygPT4l3mm/S68Ujh2BI0uDtywYIseEWBLS8dCln5ByioOlo1HTVIf+e
x2kj1EXex8MixETPDE4sXChkYZD9y9z/S+74G/un/GTrtLqD34EBn4jn9A37xfVb
VhvgLSh7xG/aPBprB8jZnOVuX6qjbPSV1DF3OP2J6d+pYbxlABANxibjzpN+/wj+
87IHDPVmY3V0o7o+qMIdyJL0CdjLgvVjqZOnOYZ+P58tZS7FaW5hzfkUbo7hdHVM
uarG+s/RHG51RpgmVxm5xPPEjnE908Cfas+lsiDUt8k0Luq5KBRdFwsl2AVNTnL5
9K0WfFuw29ADkNJoRBfJ26rtJpL3V7tzOUrOKQn4TGDvOe8B8wLaBKOz+tGoIlU4
fiQVcTTmpHJhH6TpY0K0WQ2feb1aXICLQsiuijfLLrE0AspILTXZKZdTHYi5oYXf
zzbBj52OiwMd5oWcHlTJBn1B/Mz5EAALSpmM+sei1MI98hYFV+fyjzfAzmCfoNIg
yqDftVcb7krWY+r9jou8M5DGL9foR0unNcHR5Fp2JPU=
`protect END_PROTECTED
