`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B32JpP+ih+x26cFmzoMmjQKncRB63ecrljm0YYLpIQdxHuOyshcHYClgPaKvifEj
tw7aBNgeAPdJzOPA6j+6BS8aWVozqzKHwA4KyUXohaxZpb2YwtisNn/xDTEkUoj4
rAf16GfD0OY6zn0jtsQ5GWeVhCmMIWAEZiT3OsZjeyBQQXUBGwG1nFxCogvbHil4
ruoxyn/uahK5qey9IXKYNHfGNe/INHibWmPMUXGGyxnRrdxUcKcC57ZeSAImMYHT
WBygVGAsShBWJdCriAt0W0T+iHeT82a9f4Q7rj3+T1ci6TS7Ujzbi5kFvBg4syGS
lxOWIjR158dhkyoJrR9HEOA9KlsjNj0DIeXbcbYUf4xVqZfVTPYYBAiU+dGXYhDU
nPDz5zo3JpnP9+RfzGOI7g==
`protect END_PROTECTED
