`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5l8Q4LTE6yWsIIsLFr82f6e1g3A+GqDiGVdXXZsDAG2gfwM+S305/clOzL7yFgaq
animgC01lZtvK9DdCx6pNhqzf3h8ILDwXHYKet8/OC6hseohd5uZ/NVQoQYIvx/g
MzSopujatqOOAP4GKgkeJzCMrYTVHCawRS9jxr55oPKdgLAd5eless2c5gLirQUw
maAQ3lfH41zfoM/tNpWib3ybZr63mqwA6fzPpPXT8VYYzezw7vyaBzcivx9trqvf
CilcLfFBpeWNX+BKmReAZTr5QhP+hbuYTM9JwJZyqjLXE3X1VTk7T0kSH3cuul8j
fpIK+Tgvd80Qw6/tMvpEqNCvItELSR6+HczIvdNIz5j/nCNAvlbgh1FWlwaRa+Tz
I7s8q6SfpSUV+y7f0hp6BgEoxfC/LtJa1PtM+Cnm7/6+fmR8W1Q/tm/aVMysBC5S
L5q3/gGXBtFGPiYWNflSe3Lrnp9sZHg702NbuKwt66qPSljMUajyNdnW/B9C26wZ
6ibQHc567oMY8TxWpeNhjRXYPCkWEQidsnIUCpIC4Q8L5Gq2cjVgDc052dcWf2nV
TqCrlt2TWR0N+LaBI/PGSUUmzJh1gIzSUmYQvwqXw0VN1d4RiDD6RAXm90/dumk4
libeZCICUo3ek6Yfk5Z/NvN4ym8+2oHrMNugy3AKzlLAshsvE9r/FA7N8+FNABxO
fSPE5iDPVnuQnA9Hl9VVj/Dl8MmkwBBw9oIfD2CuBh1XzShJbNI5CGTS5jCmSRLX
UwLLfvtPisX82ebU+AqVBPo7OcxKIDaYb6D6gFsibkwF8qJs8fmheWbQ5M6160cp
FHjBQOekr25ZCh6B5mUMn4VoqthFLst368mafpzOb/oAnq5asls1VlYL8eAfqKT4
ncuCAvdFcK1SlheLsfIepQ==
`protect END_PROTECTED
