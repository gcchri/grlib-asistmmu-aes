`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1EnQlh73VXwg5LqiGueHamDwjUvWJlF/dsZjSEraNi5dI51oGsnojxH/nj7TvowN
X6J2oLowVvnkUYEFUqqpZZ8V3orrmREm2lMgxRM049u8cmbbYePRtSQQhcXIRMe+
Um2A6MGwICSjEVOYo5bZS5A/3AR0MZhQaB55K4mLsiclY8NGptPOyM/JQ0TLSYBP
8Be6nr8Zx0pvIe+XmFWWJvteQjNc+4xaSlzINHnVfM8momfUViSM/YBo5XOQcuAU
IUSKuA7gJZ5UYdCvaPRe5xNsDNaBYT/30oYYXA+wz+Kuclc1O5GZI62C8sgXNU+R
haYBFaiU85VShJs0fuguyH0MTUUxBZ9z18IQgt7EMUjCW323DARbHEDVTDgp2zzg
`protect END_PROTECTED
