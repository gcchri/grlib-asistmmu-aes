`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z0I9qm6SwUFyRPswD/JKuXccC/WzwIXLaWY36U/erZIJEssrmptfFAa2sQsq4ran
lQKQU2xVx9/OFtkv+o2QDIYInNrHQCZxQ7znjQCNDgpiavNkAXP/Cf3uAom6fKcC
Qx0nQ1EAthrxfKxzJihfSkCV2udAgU3wOg63cFQ+ggi0WdYkvwnnTPaRX6XQ/GGt
jg6jcfbeu2gh1M3O24MQAzehB/NwNKZtFt45RqtjzEoCKAfGwzVho5eW8cAgjmzx
qxV1FS2LmO/HUT88LNBF+BOr65ob4oy1IUW044Ra0pISrtZZtjKe1wYES0TUkqef
ZO5c+hIKl6MbqvoegTrRe08DqNpQqaDTHVNGy3Z1nCxSfJjAFOxsd1SaVH8hc7Zy
4JA4KaZrgE9xSjyZ8CojmA==
`protect END_PROTECTED
