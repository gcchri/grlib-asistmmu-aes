`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yOKG6m49NTUMOgdCYRiODlGpRPaLOAv4RzVbdyfa3sbBkNkMjkkm5/faU+037XGv
F07z8S2lsXMceyrDpoigaY+6ED6KeCF4QVYlBS07mu/zMzfyWx8JSSG2uGV5N+vl
Ts75+bvaKnjsglHOumjEEZlGlDcVHcu0QWQhcXoRUjwxp9JAsqv8d7WJMYHSPoc1
HODBO/YpFky/T82i1yBaUeeXv938/TM1zc8rbC/F0VTR03wlCOHgPYRwG7N0bsjc
D5HgRcwGwilntKSSIfzqUQ==
`protect END_PROTECTED
