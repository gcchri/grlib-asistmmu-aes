`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kPmQ8xC2drsQL79izys9fQp6ta85C8hQM84XkMZsuewJ5FlSb7PHgbS5/lxY+Uvt
AuQk88r+yWYWsbum77SAyBsxMkzGMLhiqfsY04yozGFNUbapjHy8kLC+B1fbpEfP
cSOviaz0AucSgZ9Fa74tP/4PtSMm5aCat0YNSmF9AGWESqVuoo5vSzeW7pYxqr+6
gfNvL1ptHypYZlm0MVvUJ3YvEUR7hbe2NATTuX7kgDANmFUBvgjmF/swi/VJmwma
k+/xa5rB4jbYWnoB6NZdGNIIF9PMMXhU9cXRl3+iQD1hLPhrG1fpB8PJFc0w0iww
KHd4/Wqv7ZIW9nf2BYGGNA==
`protect END_PROTECTED
