`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UEqEdTcKmiNKWHSLAcYzndbj+83vrZN8Q5Ck3skVgJZLm3/4pPpUZpf6/DQLQ/xx
lGGqknHxKRoIXAyPmgrQFmNwijxWN6OeRKyAFt14SEMjjuWr/ZV4OopoGuuR/M6t
RnTCSwIO4NoJbP1B5hRC3rdEa6W2NFyXEBstqxe4bT9/9gG0tv/pacLTJm9liFht
GeNkvM2vOyp3kRx/GG4SbSMwAOpLfBcD6l/OnLJq/w/4vZApCsjYn2Fsu4zOhU5O
Xh9i25Gmy60HXBSu8nzXpzOzKJkFu1kp11JGLzX0NW4NZwGs1H6Y04Dy+L+d4HzR
cAwrX2K0BdQoPhAiORyMHrVsi7xM7Zia6DOkDDUWV8L0NOqdAHRgXNbgpHW20vVr
aB3Do7PT6rP6PLQQzrUblDSaboGGuWXaqjTf1zJ1ei8d/GeG//CHqFizWbtu8Psk
9rNhtGSY+4UrunewTJZLIBwEojB0FtL9P4yB7QXll1N5uHwocDrPWf6+XFxqpxis
SX6GrJqmIOn4pe4bMkRWR+htfy86AhZVqp3eQuUmYCvV23D1TBYJt0jRsQQHRN3x
dFgUFfwaKLYHpngOQVtneMJPeI+k7HWCuvk67zAEbAxIUfC/8tdA+QEyZJ6gLOBm
p1y697e5uStHIamzJXkxIQ==
`protect END_PROTECTED
