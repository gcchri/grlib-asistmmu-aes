`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LR9Grt7hFlrMHaKts8dWWBg/hQ22QhYB/1Rwojo7hiC8UpRSn5JbKGV5Hal4NT1n
ogcM+sMBsB7Jfg6FQEJFfAnA3FwgMjwcUCnW94qvtg7lUZLsUZ5ov9naWLvHpqFa
mLasE8d8L/SvSm4JCVOXAJmm0hnuo9B3du0NJ5Z8ovU2X0CPiizWrJnnDlhgsEJm
G0tPOU8C26ZxhL7kh/U1HVZniFrknfvExbwV5jyVY8/GDi1u4utzrob12rQxmgjd
t9ItFIY2ECMG2C5ygymM3rihPJKi3hOjEz4tjJGOW8frh+SNEu+gqwWN5knZmj6v
DWLucyqW/0P/M2PvMIPfgvIpKN4O3pcbBOzXtWX3Ib4O/OAdELZfDMs8cnCvDZkZ
kOA2QhWQ4wXt2MKDe5Bq8vnuc5ZrHQh2HbkpFnZ3MuG+HI32+N9sA3cW2xVF+Co5
E/lKmrIf99tTTBEHWYuqF6ItrVWXW9M46mJZfXhkOPouPt6FwRZhY4CBxHPKcgGt
GPhnEDJjoNnVP7Q4CZw9ANvsfPCJMFDpP+2WHfnLiig=
`protect END_PROTECTED
