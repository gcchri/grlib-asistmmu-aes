`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NQopptsqTnaTp9yG6UjcGIKUlrZ4kxJaGeW3XGRk8R90tIvgT/fNyFdK1fDOASMD
kk8LNOFInCENRnV5k8p3nhJbUY1lwNOuqNXApAvdG/XEMDcdx530ySQDwNf4+8zv
2ViGN7W3PV9rNxFBpdU2Q3pSvmgLz9ayIDkisouePnwa2Eeqkttz6QJoppkDxp2h
4G5wVtiPEQaUqpRIJAcBvAXliH/uffYlsiaITFrS3cDDk3VX9PhjC0FqqmDssDcS
goG9QW0Dl7AXgp2Q+Y/AeIci+eMgbJsjbenXf4EYd66o75AwxmeezzyvGdpxiAPW
1xJLRlKn9cZ25IqHrKZYL7QqxjKanSPo0Mz5brUWjUY06c4m394D6kYOsMKNg8PK
KbFSLKjxB0U86rmU5Vq+4bqo+XExhu8/qb6tsUjvtfR0x2F5R3a5eY1S3TMq/HG4
`protect END_PROTECTED
