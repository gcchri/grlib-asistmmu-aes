`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C5F+ePI+q5Euqvh9IEN5uBoNFh3y9bDN0w5CGViEoVa3rZqaiPZri4pKBWByADUK
DvSus131ig1GbgYYkATonYCxU3i3H0sXoRL01iyeyNJTXLBXdbdl5DvR27luGrHg
56RANDGR2p84iYCYstX2SxWxGrtGXq9Y2x0UI7udm/lUUnccE4YFZr6HpCIGHxoB
39UMrgcXFulgKmzLu8zFPMW5UQyDNDFCslIJJRySJrrG8zphKcZe9eqGWo7SOxzt
XX4CpSObc1isi4eygguuNWZakSRjCzgSGuRBtEdtapSD+/M6Kfw0VO3GoHJdzOYq
R/SHFm5a94v0kPgP7K37jHAe0KkJY+2ffRWJ9NNTuU9eOXOoUcSxIgXDtxGG0mNd
Pp0O1oVRrlerpF/7VuhkDvpCuz+c3Ft9kE8AVlg3laDbYSIrg8cCWPTRoPBUAv9T
YxS/E+W4mb6d0aiMBIoZLkK66OGgHuRkHZpzY2bi06nKcox5EJqIEZuwPmJzvVsA
avVQF1JaxB6QIi5fRyD/kGloEhqrahFmT9QlcYHx0B+bPvZKz2KG4sB366pNagQF
B23pk/8zyE7+8jkSVSuOLCzK38lq3e+PrvlbjfPHXKiH0MdT8Bnpt7+M83MNDnrI
6U8wDQLioMrXfCYSk5Yh8m2QbnXPf6n/LEMX7FxzWAaj08gWUReOHhznxviSZdib
h3O31CzAePXTVQuyamVH4/UeaFs85y0Ok/EcFJloVO5Og20rjJym2ZlOR6yTnd7J
`protect END_PROTECTED
