`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LKmvLoJ6qloN029mI0tds60Xon218LD90Q+5Z4ifrnZrQZTdzCaIWG2nyZ35KQsp
50VifoXnROSxYyL4e+IEUIFRZOcs/wUlionhJlJVDqIAR5VVeDrHztBoDHT85pBh
n4HSyTqPs4loGfnM0Tc+FNplCt7Lao+3gqx52wMW6QwGDHrptYCwHHL0DGrO4hUA
X1bbkPEG2NBzQS/sbuz2sNf1Lf1FSiyoHJAE3M97sqPo1PwTeMUwC2WGZAi6vJPi
A9ruyUw8S12evlNEjP4q6ST6JtwU3Tpy+aEwwkJ8tnL+Gaix+K0meC2C2Rjv8YMC
vGldjRftjyfO1OKZPTdAou3cLbh2oGPQNRKaGSglUHl5C1SJed2O5Ab+s5tqYlkN
hsoRhT+fDxLpZxxi3914zineIkU/L0kuJlG7nxjK49pWseSu/UaCZt4InjuM2R2+
`protect END_PROTECTED
