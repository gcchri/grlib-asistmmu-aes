`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FaRRYWuA6TXzO0j9UuPBX3wv+TEIUhkuCPm82Odio+XlrN034sYc/uDasaV97sa1
XuhMaW2UxJyJ+fyhzHfi1Fx5h8yzNAH6sQorW66VhqBFspfH79pPm2y70Wrl6ft+
2aoB9HUcCknoQnn+SLpNJGT24cWB7wf1jpsKjUXzPxnFnxudffYCPwK+5Z/QLu8g
btwPLPE9At1e1Wv4ItxKBj5qk7OAGIvs+ZqbUYOD7DYo7yB6vnV2BN3pnUsgqs9U
ARHvb+0R5eNTurSiy6KazNBcEzofDzJ1uv4N+jO1YUUKhbTA1+rfpCqmVnhC4mhN
IBA+ssbsj3afmdo0fX/CK4vALlylCi3WyTCnBkNI9lk=
`protect END_PROTECTED
