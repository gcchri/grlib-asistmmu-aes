`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fh8hQZuwb/jaWfa2tuNRjgC1JhJZHSAwm0chuTa3IKw0od4Cm9H9Ik6FLHhTfBZp
53dId4Lo/bYzKOsCksFbtlQ0iOwoUTreiqDyF2QMOMRD7KQeQAgtjrTjLzXjlTO6
tctK0nYFjxfL3FkOZ2UJcXsvqp/3RISwZ70vsTZht7hsj/HjoygiXN+0sTNt7Myv
ByhEOXKv4/Jq3ZtqXSxYOGM6Oym7F+1DanzOIqH7Z14ypOxRkobukSZ0qZr+bzXQ
tXdhupri7q78UCZuJqP05OpslFbe3TJymPdDK3zNTgF/3/TUL/WmFBju5NPuV9jU
aSm9oCqKdMhXpxXRS7x62G3i4uaXWl1nauHa1RGSJi8ZA/fKctJ2wEnZRTJNzP70
wFxuI2K3OCkSPpNLTyj4Jw0Ul0HXIJEM55Nh47eByAgYqLjg0DQjYP3+f0pfwk0T
PmOSE1w8fJrQZky6Gnuljb1c3Kh4xRfLlUZJInmLQmTYje1IRymRVC2XakZka+mF
4xl7dq3+5BbuYj4A1/uKBPMzEA47C1j7duDape0+wBz9Mxt5YgYjJHdvWfRcsGHL
P+8pogok794N/nT6JTcpNrxlisIipplSU8LcFaQqyAXnTzeIuXi/5LAqQ9jRPAVT
vJnSlPJx0xCor5bgsjxDVLpVBKb4lA3V61vBwNSTVMKHczqmNzWtfwi5WkmUlDQY
jXuQzozXs9TANJlTYJgukYl2cpJZ+F84fDaQ1VYHu1KFjvJJSbnyBCksNz5OPIit
hTqo3n/RCVQ/IuuPXLqzAm6ZS0b/XZv/BkjTu5yoE4CkF+AAaSGkeo1Nb1knDoKN
r8IvvkrmvA5QUULHdNvlqQ==
`protect END_PROTECTED
