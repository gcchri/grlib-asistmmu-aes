`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FF0Pfo9Wd5h9gtoOl3osT3GYCIfQd+qCkYcbqKI6uTfAuR3RmALHKHamN9UBwSiy
3he3csyYlPcVh8zHjCgxQ36QPSLdFBCNAEUQLwUuH9y3mBzYarm/TQW96yE9X8fy
a+ULHVLatj8ApAhMPoXtgfiH5M5uIJxnx+bJZT+c8hzhekdwr9xqQ1X+Lk56QAFk
psgnzLpldOCnBo8KQD6avbKEHIBlxVgcrUAwpGmZU7jsA4ps8OyiBWH8nh4vcAwM
fr38Pv5meq6WPrWaA7gwNh4OSaToyau3rPPfQPAjP0r0PFWM9ooYPib1u7aooGUf
ASb5luKSfH7xEMCFORhxdQ==
`protect END_PROTECTED
