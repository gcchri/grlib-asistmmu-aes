`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r+XWv/FI1SPgoDQLiqVEw3bOgUsjP1dJ/4rocdnQlH/YBk72D8zZXNV8MTslQF2+
eC0HP5DQAzM5F/LpX1dvNAR+5mYKknQ+dFslB7Hdjo6fC4rhYrbXkw+hdvDZSIzF
XGeWezYpba/t6K0KJmdNESLATVbR562rw2uKGIt4GfEq7QEM0f3QS72Xr1vnv89y
+mFHh9/PAw9CQLYCPQxBFb05WbJ46RBKMB6kOc6Mt6rHBUqLAPuGNBXrFJ+t8x8t
cDatLovM0lyxTejYoADql78sqdSSmOLpOSdnfPh/Hag3YEa33LMc4QePwoXV8ZUo
3FbZVLLKzwG4hEsO6MJzEHK/B0iDxQu4wXGezNDEFK2/2Y/4823oSH1eqn/zoMnJ
7HJBEuTR2FK2J/DxQRe59ZtVbHVsKknEZNOn1UK/TmyLAX2xzr9K6stXQA8Th/Zk
arABpi1oDjYB1XwUCSnREjuwE6DZgSO8IlO8HDkJeZK9QtYpm/zJ1PCWChAgEDp2
b0ruoJJdc8rapznbY0MfZsziQFQ2bU77rERQBcdln25Ves9v2lMc6GusrFLCuUQE
SgwOwG1k9oa0bbo6oHw7uh7C0V3zun/QRt4znuOUvWeCmAH+0WfdWmcRnHYmU7bb
`protect END_PROTECTED
