`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mc1+QRZpgURLfKeEnRbM5L1XxB8bmUnQSRmuAx3h2h4XuXhlE/wZwFR7FcCQAsDg
njSp5fZSPL6o0aQTb54uvGqSg35B+RSmvqWnACaLVabUyhyVY9mewlkglwu81Y+X
K5eBvDdWgnTd9C8qBnKkC1hEB/OA/cjbHzFKZyO/J0c2VIDr+4lfOv1cjw1nwAdu
isosVdciSMeune0x8CPkI738V5N+BV2H9TRdohCxkQhaeDdH+ssKUa667nNBWezf
hyFhP27mc+LunloUUkfbHO+e+7/fy1+K2zB1mwugczBzjgELJ8Ns9tQZiv8yUCEA
YTMCtaKIcOKx79dBR2t8dPVQv/qmCiI/OFfIsjTboLMEd23/WmIws3pUZ0RuGqCf
fppfX4Z7QLKepMEiQwnI7wYs0+O1fxKajcHnXN7tZLc1W81XaQMkH3ZNS3hlaRRN
PEz8toNA+j6FXlB2X6kGk4/VyGE4hi6JQPwK5FeHIll2W+copP0GL/HuKv7u/qUC
MQ9HWmDKfxkt6I8kjNCC1uwtQUWMm/Wd2fSg5MC5W1dlvAE+96isDaCTsaAfPsPe
Kg+ZXdKjGcWdDvCoHw39qOwye/jrzosFXIuKOCiSI7XdPgMSL4LvuUKLa3wVpsJs
bFQxicJ3nni2+6nOlbD0J4qefZ3FNe5hPeSp0DzCD36G2ejOEfyGooD2IGoWmyug
Lw1tkIfFjkR2jFBKTSEQbFVaq6Nx6TA6rj3uoFeDqmdFp78iQvZyCk+cjRTZxCJK
NKB97YgC/MRSl3I3pw//q2tGKzPPI+T9Hk+EgZZoLiWiMbtKolb42sz0i0Eo/8wG
MxfQmu2fagQ/kafiNHDmmBQz5dPgGsL1dqc2woILm2o=
`protect END_PROTECTED
