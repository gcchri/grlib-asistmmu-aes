`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O0f1sPKFCaMsHEFhNAhN/RJt89FiuLVG34oB4Q+xhNBZ0E9mXJ/hNrKc6Rs8kcbb
IaTJ4yyjN41fzXbpdCahvqrj8vjjWJli4mPrSwayrEuna+lCKRkPQObA9aZ3hXrs
ALD8X7WCby/3V5ttfs0EmkCMZ7fp+pEr+1WfG3hinj0osBr3I4RacIR8NSW5WrRm
UshpjS2bPXkjiyJfKKmnaANj8y/GCjeEyT0o0mjC/pvf6g63NwNwb2Ou47h9I8Xg
p7C+8T64dKoTDuvRV659jV9EJl8Yeg8e4jgwJMs+8IMQ4eMje07S3CnTS0ierpbb
aWiJy9+u6PiaxlgVAsD5mPohFY7Paqx3eCSBG+H/LgjjFYJpG1rZi3IAc5A5qj2/
aZZZSSDTyVIHjHkCbjx0cPTbxMNu5+cqcmA8Mj0NSMMY5uQj4nyD2Ixz7NK21GR4
0YbWp9qPQbs8oPqFUUnKwirCBtsTZ5AeoElsQktUHq3abMpwzDeZkGFFBIO1Xw7X
WXprV7vtt30dVgh+bEdUFbGJWd4ePIKRbaKhY77xUO2ty9MPkO9figp78Ms4DTkM
zs2nV2fafKNPzqoKABbGTDTYXDTmTSsGZeX+7h+9LzJ0Ki1Tkpx9zjQQ+1mA0nwQ
YFFqmtTF1oUxMOLAWYQKw/BTogt88chawfabZuO59BNNt//3wfeSvxgx5x1vORp+
c2dsZwzb8LEwg85TPF61kLcETxAn2L9dyi1c/75Z1R/OE2+NyB2B62w1lM5j3+As
W24wCdzwMy9b2Fa8Kz9troFwcVu63K+gKi7xTQ7OKniWt9cfjNjh7RtuSybw5hkW
`protect END_PROTECTED
