`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kwwZq3sYzOa8tFI9F2GaQxMwu8g1X8nR2m8gJ+rTVCVlD7zbqljfDBGxbvl9iwSH
B227scOlE7Pi071V8uOEACeF3kkkCbsdWBbIwDIS0zzPlyDVXuGZWvin/bTRCasv
PtRHBjLg2aqH9B6fSOLC2mG+y33rUzvceaItcy5JQLHoj0qUHvfsguLjapac3z6g
+NIu/qB9m5+oO92EaLUFW0PhqxhYgBoekcAOha2T5/d9FT7aQtXcrpkK9i6BXu6f
ZcYVUlrlZrFR3vq/XBc8HoBiBk874mdbovbsHSnTq+uSIi6JAJeO1nFBSYWGp2wb
kaa8bATOOTN6YKVX/aOH9qHe70V1/O0vgqkhSchlUfy4iTlKRwk5bF8dbNtvX1Uv
RalMyVaCiipD+EPmmwcBVA==
`protect END_PROTECTED
