`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r9iob1ddYT2F0Vi/CCNANf+mJYs0/mqg2/XFbxOf3Bth3h0e7DgbX1FKbkzla+FI
8/HeBywwGvtCrA4GpTUuasVRCKw9KfFXzTT4hfUKvVMZ7FFsnSyLBfPErXETEseV
zAsKn847yms0QDZ5jv5OaNP87ouWP3DCcL+GbrLm6isu5PFpIxqvwuB6dFbzcAz1
Tf2yj/gBTu51nYo06FZQ+QRmmGK524DCt4n8UNav0Yt7yvJOKJb4JYHOjhLTZxAJ
cLGvhKKBeLstOLjOHkZbWGJxpDhKa/iBoMwBFbba82KwBo17i0dIGO960TA1Iw5u
rAXBsX82mqD7H1bqRroQnvVDV43RqRM1jHRVnulMEC71+SD3/ej5zOSiez5qAaPQ
+GkpyDrPLz5taigTeM+qTxzueEBmvZ9OjRWFm2Lv9Lym7VHK+rvWmn20S8MxqIWB
XZJnTBhnpJJmMv0ID84Nq/hG2PrA9x+65sTLnymFyIzEF590QOj9FWslyim+nuF3
Se3udk1XsJRarjmQy+WoroM829RXd9VI0nruqN+OYSXd/nvhvaF6DxbyWlMY2Nwy
sLpxwbjfTIl5tNzmRxdGRCgjg9JJA8/7PbPxQ5/+vPHZ9M3meM1P6jHw7+WA5zUP
5oyaxpRHxLX3IMJPfXwhuotMX4YG7Kd/zarFOHSFxJt6KwOMfuMck4Dy2obp0O41
+UYJrKmqvQN30pmGVQTv6LDu7Gv16Gg7XuL/dfJte+zZ8sVoe2M+HsJf/rSOrx6s
jt+rYP4DD1pxMh16nVgaCaYYI3iLPsHpdg+JQhTZDTS5+HpfaqslsRODaRdgmFXA
1VBIB8f0yeNvTw+I47OABYuzeX77PZvRf0Hg5c1z5/6+tfbKIELF9SUBshuRAyJO
2Fi+lo1vzkvMbrvoIsWhcuWKwnefHhtwkYzQCWLQ/4IMSSGCCS/Z0M65D1KWHg1x
KtNtz0TsGmTYAvO4yEURvkn3NSJYPnSzJTSmeTltRFYCsIFBkojBsuhEUndl66t1
`protect END_PROTECTED
