`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7m1w0j7XxGwcB62obbEgu3sp+WxdKyGl84og0GT9SO+NNWqrBjSCthQ/RMgNNGMd
6A96H9L3CQp1S56jCjTbTulzOvnP5M84oZ6pKYS4vbieZOBYH0EChkV2c86q3fdn
agSPahj2UfJChOJjRo4FNEgV4Q/7HmJOHklZu4YwRGWGaKbbAqw6dTjwd0p3PPyL
WASLBok5jQpgca0JBmg9vl+sol3dUxTWD/M2enhC3xhbUECDbn0/6FJ8ufZcSyM8
9Uu+W73H5alBQq2HRSgbdA==
`protect END_PROTECTED
