`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PiW45wpk2GjdixwmurAufX4YBeXqjcapSUjpdt4+h/gES+ZoM6kxGG0MM402fDI+
biBF4kbu8YPF2ElH8mlm5XKpYjrXZgV2KZsvX/rxgCrBp+Mfb8zez8zkGtT9r+mQ
Z2tDGkfDlM/eC86Xovvvo0mun1M2EZygJXZUIgWPb5mquYVRkP+fe7wyRksyBtO1
rH8wKNd5vTXVAFc9DS9cG9PC1ToOmk08de8im5GRIXnZZBbria7wpihMhy6/dfu/
gLGIT29wn4+4M3lD6En9Kse49S3pD8uJCd8EHWnVC6ts1ARZuv5E8yxbDHSJ7zlj
tXVDJ9xv5W+Awxjqg49pNxU4n+l4mZhwZQZXESqJTLmSe6FdBWt5bnB/MRAEdgio
1KxDWaFbmWM0YRXSMSiemedWKs4PwSJfBQiJ4DW6XdU9QNXO0BBDondIcV6Bpa2R
megm4Yocj28WyTlDFp7sZ6Ky6wMWEo9I3hHVSMJcPrDT4cMf4seQuVtptSoOmh58
+PhtOxqfKpQFP+I7RJgzj25MLku1HhHkBYxfzUuFzOtYJBmo96pSjxkP5NQcQOLq
oUxe3dPQ17GeAJR9oLj39Db0ue/Y2MjutDMzGWgnipB77og1ovFN4mJ8ZDfJZzFS
/Cqdi5uzVdK2a+cICmov36daWH4AD2m9UHMh7LQYnqYh/urC/G+eDZU54Juchb2h
Db+Z5os8QHfwUJE/fcUqEaQ+bPaIAU2036QIVQDk9CFloUqMtpjgcUfcCY2g+tWC
i37InF8ZRxiFCKTA65p03Z6GJMWeHGltQt5b3yhaOh6IgTSn+XusgOQflHJKNcSq
k+w7/1CKdQmh9CFaulsG3mYpAayjOlHJquY9priieVeoZkF4Nzecj3q1b6mqQhCl
84m+YEB7QjBg0LIjTPOnOFne3Y6F6zXFUY36nT1dBGs0qgaG098GrXUcNgiEEzoj
W7jDVyp5laC9SFBC1UskoHiLHUKI0dkIF7W2iFeWcKiOgMTjgLRkOTgl319H5IsN
45VFUEcOnesFU1F+ezuMl9+GGNgvmDsQfrSR7oEIHrJv685seTQgsMVNxCOPcMtG
XinN+0fouxA6odsvev7qGtWznyOv0KRmMslknpIC4zqWg/hGDYTckh16repObq4s
8FEj3do8W1Dws71KXcnWgscZkPo7+oYM3DagH0nGNTih3s8/ofY1IyJJKZPiu6Ch
gBEppGhxrJSpdcuyxlqXK+MEoDBfqRKIz4k0xdF70s1A4eEUwsmRmx73dIpCXEgu
kKIoVSsJMcOiRjdcm/z2+8xXtJZ4CtASMdBei6LGJyRi1DNMIu031Wo5E3ik0VzG
tsvBUdt7vmJ3Q5UZbXKNMUHqxo6fnEo2dEMIWmFfvBY3PUD28lD/DPeWpaF4ZV/w
TSnMamtD/fomyTLe+6E2gIppNSbZkKIFcmJr/f5RILyjznfVn+mW9H0F+haYAedn
e2/c+gF5E9CwHNbN1AHt4DNT8n7yd8/zoFInEayJYqY=
`protect END_PROTECTED
