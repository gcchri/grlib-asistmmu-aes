`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F4deItuyjfHJisAzxthYxbKF3uxs7U+SIlwD50mnIk2TrvyV39hppbEuphjIy73N
Y9WUQTtzrLMrP4DFPoHFlDLXn6zCoFIGMCRqiFEd6IDhGdnBw/il0/OHYPEP448v
P7YGm3DCK7ylyJpe0fyaHHspfoEPK34CtI5DenrTfszrm87tFFHljqFIG6HChttG
XkgYzEuH1P6ytJIlmj/7w84neKdhc8wbSBXrh769AKdj29NqlxQTKoSCKP4MQI+K
cv8AxeatopRtqzYlQXp3oQZplOma9jiL1Wabo65v4v9dk/vpcJt5YfgungxLZ4D2
cwNfHN0cWaT8iE9hVOqLY99G0WkCAas3RjrRJQ7F2KG3M1lFA96Lm47ukMQtVI2m
2ncKQ5c2T2pqJcrsVm/OjX6ayT+4P+kEzpFhwkTReBpR0LvRIOdS0VK9vshsjhBG
5HDJ+Lld/0be35AM6TFj3VNCtEOsmwGh/0knPjuhFYSet9cFjTYY203ZjDJ1ON01
P7LP+AxtW73ptbqxU2OYKCFkdG6hJFlZlWNfic8cRJOJiyY0Nm4/Iw90WdScrIHd
Ta2ObwAocIG7824lpb3vpcsNdiWaXEBTcvabgV7+Bigm6DoS1iNUWdpMMEwFJyFh
GNH8XLkeWc8DS6cxYKg1V8N5EgwoMxrVdfp3Tcl96UFe6bw9XNVsxczN7IE7ZkSg
q7YxyTTT4ri2ZwMg4MQ2hYMVAOIlhj25uQ57kdZCGyCCMydc5VEGooR7euqWRt/c
pKMyzGZd+YowWavrSTFZB071I5tMHHbi/RQC2plOHP8Vat9VQrujI6sgvUaCdxxl
RvGrpfXS+r9WQ0M5KN0S9l6QDQiIseLPQN4twFBfjWqX/PqMkL0pMmBtqA5kVSpp
/711X3EgcZ3cSv9jhiaORIO6iqdYNS2CP+QK655MTNrJv3YmW/OXBxHR8BiezcVh
xM09jsWSf8Aj9unJPoFKkU1JzViJqNzG99Bq7NwkWgieIRcmOJF85cgmh+oDn9FU
B+2rUFqWUD8S+yzCk6pWDGzGkTraisdfoBGH3ksncU+xTgvWXLci1uOyNu/S5Wr3
HLv15S9OAYZRroKBk15TQyWenDqko8dee9aBidg43acOc40o/sX3jatBvf7AT8mn
hV92Q3pheHs9tjCEpewPh8xRO5+vkWgck8MZgDRYh11iMGbcbmtOqHhywsR4ZSpm
2v4j7gPmoSgYrtw2a/iUrNY+9klFyDW0eC9Is2z9KTy4TCNA97ZYjrV1cy6iueQZ
MmzvOS0+VrH1DUgZJNGu/R+2jxtdpX1P4JDivZ1wOx54osbeY96WrMsE10mkc0g7
kXXIw2GRu7vcnfOA2JIqc9BdWkRQJkOIB/+Kx9tPaT5Tm74BwJtvsMRYeIyXZfKv
YowxDDCgv7zLff8bTt7K3WB/XYc27nymOJ4Y8t+Foo8K5tROmZ1cOCgDHuwCP+PH
BffRRw1fUe92gyzF6SIKbQ5fynN0EozbJRNsi2W2EaO/dduoHKp94ZAZ9sMRB1qQ
TL85e20oaBwaPA70AlWH/a4Jd7RPAJO5F7l3jpF0zlG7s0OXKDYu4bi8yOYZjoxE
pr1bUaW3Q6Me16lxWRbWxicgRDCdyzDkfq18NQJPY7qJj1qTw4dvi3DNaZcVOOSv
t/hGyh6Km75PJQ0LSEYBsqU0eutiU8FI6ZhZlGvvQEXwBHBtiel2Hvxw8kmGWcuK
2JSLlUidu5Rs5FNSIulcyTXA+uXRrZF0INJIV7tggeTcDbhyXiYsvddILrTTpYY/
mWRmxgmfUhRppMsV9Pt7QIyat7VU+6+tCCi09sbo+5W/d+zJFuc9ebRfC/6X69l/
alfV584Am33yarlfSk3pyzZZhdy8VAnp6TU04Luszn8k34VR7sGcufOcLoztZupG
+WMOSSm5sGCzWVmGjifm1NTamiwxdkf2U7xA4NII1f26VIVfF58oMl7hGbHmaLTs
bOIGRPkqPrqKnVskFDu4ifPy36PkFNDHWospcQ3NHpW2MWp6iLZ67cfeFgKgl4aQ
ohz8fElwnLca+VHjRsnmQdppbfDQh560VUmyfffgdH5PTGkEeAb4Ber5duzquGaq
u6f5ObrfsAGiU1JZXtUtzBmi9+VtvIg2hAXgmCTHoFyVRkFtPRNL2w8WYy+N8kqr
CPmkCpRRZwkPYLM+z3PL24CEDaFEskTPIKSTNjpLJtUW8X2mHa3GhSBFclGkpHZ3
rP/vvITA4CQJ9oh4PUorFBaYZq1YnF/ueGD8kOzeY8FlMWF1/mfB7Lngw7v8/wy9
TdvtwPeqTL0zLQ73KIq5aRFGVlsfVO43kbR06TYdN6ymRiwgHlm2oGdwn1glvBU4
CT1r4iNclblcpKiREKJYNSiNb3IEGxHvVzXFAcm1lGLW6UvAyaG9KFehQay93oYA
eq2unHcJRRwQCJrbNWkpRdo+x95LKYKV9ql4lQl+tNob2HEwr+KXd6qNW0PV2gu7
o3PqiPVT8YNEk4ksX6LIupri265A+DlAOafjN9H9zQ+eM/MB4411MP9cHfrpVtdq
mCjMXQYXVdQHSpxR0nb49YnwWPnVmEvzHv0RihPFznXtz8bhEA18i8v7KF/lkhPB
ooS1kNZ7QciSfMYcmOgv9GVW96U5Iidllo3avmXm0gZ34HTYTLQ93xUq0OtR90uh
Oad0CbMqC9Ipm+VGA8CZAnfreNGfmvrTouHWqwjonItxt8oSCQScuhAeUyTcG7Ti
kmJcuO77Rs7LTyjom2a5yB1RKx1DGc2SVm8QvElginuuOfL6zWGJ2rsESCFmtPgt
fCpnkp634oym7On4jjAWQz0GovW+R5OsLNSkVTm3vHAWP0trnexvY3QUm39zaIeR
Eveu0UvLho5y0LvK9Ox/OedBikVNUjJMwbmUejTyiGorbR1iifklMjE2huwZ81v2
oCKRBvXNpYZGDV3HrP3CS3LbtYVYi0lb1OhHYJ7IVx2mbjuhxp4/gdTgPOJYaENE
UUUb7d/7XAbWdtOMlUW5c/BXzK61zbYpn/ny7YF8xJoPbGiLZZyBS3w2vKbBFASs
P2p6w8xwHBVQw9MvllyljfBAS+MePwoiZ0Xzn3VgrSEUPyGGACS7RKYAxHWr2DqO
Mp6CTsu0IhaIR7bh/jll79uJ2QnjmUxBJ+L9juoLzbTpIe+dacHolPEucUdm5Phm
8gn5trlvUsJj0d/AYDeQjusjPyqRTis/WmN3HmD0BRGVtTpp1tngXBBNjoS1YEp+
mWc4Ogw5T75FbMxuOjdQ55SGlQoifql7pYDJBUpAV5B/+COCpBqN3NtoKfxM972Y
HAP+ya1Fpq/fSX+2xc7BVGJ5ED7PNQzrm+EGRaA3mSXxJ8p6CAVXCi5icjG99cXm
OoA4hfp/q2gdG63tmpP2e1BjPfL4D12Gr1WryP/2/6+VmjrFMRfrEEk/fYOYSRGW
H9TlUPhe4PVp2zd9gUxq03WILCLQKjv9rYkbamIu93T3FgM1kIihDFQxBHsFZ4D0
StfLxawjvjBgtWlIGPfa6sZiW6pqUaheimYr1LiAkipGiUbX+7v+NFyMlCzxqDnl
4mcfjl/uznr2+oVdF+97iAXTNPcVvqEoI7hGzkNhwvxiBFAJbAYbJLTBsWCVdPV7
W4I2XiQRovBSQX8378P+LdjU+yR9CEZ4Zppw/y0Ry5DbXrAl9c7Q13ZW+n5uPxV6
X4Ii0FQ8EtsbypwW8JmTzCtit1Qjl8YciO8b2KYgw3raya2Up7m/a0TibrJuAwzG
uskeTHR+lfP82aXS5Q2EG1XneUk72Rbb3QIIDhhfEcuhv1ct6pS9Xpi7tISHlNKC
IGFoNKoXLl0LPip/A+tDCzhcObUZ4X4w0VPVoXJRNeomxZiWcOynIXSsK6zIAKst
OqdHxlPHPZEKpFMvDdC+1nMhpPmAHDmHXxiwnr2JBEL7f3M5EKNOBsw1ic5JiFQc
oPVUfYC6X/K9WWXvNAZA+F35AsmQRjK8orZB7awvTg5hgYYp5IhMXbRxNYrxHHgw
pGde2SBcPUR7Xm2kZsmcFDzEcPFq3bq1Smy6lp6fjF7Gl3djT7lBtUbdAq2S9wws
9FlEATXk7UUXwU+u+DWkpdr3pwMN6JzlLPJl0PndB3XtQIM4qH6CmFhKY9zzXRXU
iReXiaKt7kC8X8s5gtedtMMRk7MqwxWmrCoYHWGmeJ6Vik58JntchF4SIuZ+BK5q
uxdmAR7YWoA/E7SRehC7gAjrI9ROMPi+qEUbpvKyziWUS68IHLZHYwwMmE5PGWhJ
hqLPhcMtju/hO/5YD3+RmaERQL7L4xjEy/HgBWqE1o9rKOlJuE0cVXxIujtL/jxL
gdgvWzCUkyrXDap/F9NNoESqsCtD8hMsZJEdTZFZt66xOUy7MCqjgIC8nyQkWlwE
ZKdX1Bq1imbfKmTzRzarXH+ER4uy47qHr1aMtA42AqGg1BkXAtEno3N480xGxSLs
q4Ce/qCokSZ//2dDAANXkP1fzawkJIYhv0wywkOQGK1eD2vHcOMfyVqPkT5Xqg/P
/gUXTRBC+gyl40x4ppAVrXN1spBeQbnNAT9AXdLn2Rg0AsCCaVu9t6wsk7TmKamr
AzDT+eE87I8azulVckieDs9nl/Q4omyJ4SO1TVR4g9zzui3qRCTyRiASbKkOFuq7
Y6WWdvMw5X8VD9OxPBizk+kG6TFh0GZG0a2W5UowfNeAmuJzC8pt3KruJmwatyew
FurbgdphElkOsXS2AfYMWfN/Zyz4EoWh358T2vVZFo035y0z/Rqzqr9779Dvy2o4
USDn7R8LUl+8o0qR5GK002HkS/IW9xB+L05FGw9bcfkNCUrQ2AFWxOHyTyRIa2A6
MyV2wpjM3XEEb0jSht7QN9DmCJjLykQvI3mZ5ELRcs1s/F/uT5K+KAeWNqJazGni
PusuXV+vhayVcovxRcIHOHguhsCLl6sIvz8azIHpZTW2brfhCEe788cKCgbd6gtD
af0FaTFYP3uLFGGLadkmA0f1Adx5Jb8rhwwGD1KTHN0hf1s9xV2sF9/j/Kfsqecc
/v6zXyeASTInl3h43opvI5J3JRYky3w2TFeQfDP/d3s2sRmdt49W2FS2xC9oP619
tpdq+zkdv+XegUHqgOqanXUZEc1ebwO9xzktwsIxhqrar/U8//aT/sc7m3J3TrBa
w/cycROanwJ/+P1Rnj+wUj37r9+u+tCn1cgBy3P35EtTIwzcUFKg7LpJiTQq8Gus
UMX3BVIQgoDeUOBYvqwVKRTjOcX8mEjKwKwWpEDUsAUZx7Buev79Rra/6elIFD5t
yuDaMJR+vAd5YgOP5R8cI4Lz4jqklloK8S70uEDFXi77obg/n2YzBjduSwPodGcL
qMMT9WMufSSj4Ru0XMlnIDSRWU5pQOkY1tMgyYXLcvVy2pF7it0a7q0GUby1mMyD
SgKqkM1vvRLO/kWYin0MouarXs8nHeZ0j9kiSfRzd3PwlpHXic7/ce+Td7m7JXV7
722nWBazf2vskU4AJUXzp1KR5rpLxOojlw/pDy+Ogfk4VVyKZ1HUvlKJdbg0HVj0
S8dbhpNNeji+jVfUDDoiVJ07lZ0rFyg3YTr7PPFRTIJy7Nesc14VGWv5wp+zGCU2
Wq0WgFIE+cyDfgSQnbPCGi81aIZRP010EaSkhGb3BcJG49xGKAUeIhh3iuhEsvA9
02ljoel6jiOqenohPizTcIszNCwOj/1oRdAY6MJ49ibL/qZNc7kiXYsxgyBwfm5s
N89O5CfgkThTY6V3Ap4LxulDaYvjk1YWdIlVQNX4T21/sIZKZzs81udUEx/ezLyG
8bP4gIE4Re9XUHhThBJcNhuWDnNa6jyN63+np0fsbqtFhvCDXasbtWmJgo3cJPe8
u1KDyTn+PT7U2HNfzrVvZ1Z6qBJ4KHtiVG+MRP9OBTz80JmM2QYaKqE2ljMNWdtG
rSB+W0dQ9lVpfRYLxIPuyvVYkFTp0ILYDL2uT8RNvCfefuIy0q09vpK678oL/ouX
63I6BJQbgps9/dnLS6yLZMWf953vAx3uxXUvFu5CXlO5YsVtm0T4ufnx49n9le+m
DAu2BvxN857D2xDIDxSDQXHywAHYcwH8syXmuS9B3Xmu5WU3e28ESTn8LASB4dzA
i9I6sA8fjFbPyJoPtqWOM0LHMuGMHPbD2nvvh/jHEOq1TTjtn+xxUbKqIcZQUrBK
SuS1b3ypAPCYiAjXoHgUgzfncOC43cJ0Kx1dKIzb3TLFiwvy0X59qFMLCjFJQ2q8
bNI6NmQpt2UidFZ/Ti3pN8OlfxQe4ux0em45ub123QCHxK+33WknlHih0yOSGKL7
y8vmx+T8jD+x1mzeemedAeWqurIA5oesYFPFulF5T+rr6z2JMpaJkgUF6WtRoAVv
snJKePEO50g5ma2et2x1Muv9Ikf2765C09ac1jh8ouL8IAyRDoxg+39YgP987sM7
0GxmHtSCYhnYHOCstl3SGLypI/DrAc16t682rtAc2wBFwB1w6fgGBdKlWLDUAsh3
Dvej+FOfR1Fz7BWKq4OZL9oRoYi5E95pDb53PrVVF/B9pwXkXYvbu4Ze+ZZ6A25f
ZPZMyJrjmcB5dQCTESkLWsu3PA0seYJeZ4vnfxxE1jpWoLdtMIxnQBxLGrL2LHHs
6LH39Iupptx96WTXYKuDm70R5+oMk6dDSnW3nh15mbJKZmGOYeGbb60aRnJmjBSa
eAPscyNNLy9dGLeywFzmFHekAqyPkwTkzCoA/Y8em2gft2wu5CYIrTSU5/gCv4F+
EWbKGqwY3Q76WV5PJQhfsbrG8dX4WyoqTlN/7DpJQLnNOQBUj6LKY8SzJ6VuSuh4
bJGsGR8LCSU71eOHpxXRtpsFOWuKsVFI5p02qlvoPch0m20kWTWXYKpEucDNqvXd
X8X5jmm/QKbcc2LVnAz4+z/VuKq/IS+0Dc5ykcUr6ungeqJG1VE276ktNfY41OPr
viIimKJShgzXBFpZqCkBRfsQM8Lywf66RKBnMKZ0jTF9BsqCSTgcX1bTVzadEbcg
D2H1r1kMa4ZD7utty8ur1d6RmDqGGN9LDQHe5PXKAIzA1+mLzsMCr96upN8kkZO1
iyPEQ0iUtDJeKFBSDrL9X7JV/15A33RzWW7XQf4rnU4k4rOSBDE86xXyVH5dHtEa
37b24KAH4YCKvhkrFkWLga7CCoS4ZhyMAJqUGe9QmQc1+v6E3t/l9LbB8HPEvoa+
zK/FIvu71JIH5xlJ8hZr3ZuCh1fgUA0jsW3CJROMgucGazxxZGnfBzggO7IFGp9k
8S1aP9UeHqsE9bnrfi8rYH58U3TpI6roZby8Dld2N9xVsA1o7Yda8E4cigyfmx6X
GD2RXWMfiA9u7/I3D/0Jnnj9jceet6aPcNreERbm6zahwCOOkUkN3WHlE9M/0fHe
sZVBdx0QtIUOq6SHY0nOT1uiOHLfixnD3PMDKkJlBd+a67dySA0buYbGNNjveve1
tgWCzFlAsOosHZQ0FVHVRWOkzZpG8sJN4cAaPxDYkY6ofWOhQ2LuSYgpHwUrBsWQ
rYYge03iwfbyWyl/amdwDaxLq7/rwCzzKSVT3Z0Lm5oEKoJygA/eBxncLdM3WL72
L9hM0oLQ56WduF+f7LVT6DvYpKMD6xVxOOOmFEu0GM+d2pZezPPpHDfqlaTYLpWe
uvzSE05FpjTNmzcR/Hvx8/GhfuoM1Bu/ImGQV+wp20XG7cZpRMKECJRipLbftPrg
sWgpWeCrznKanLFuFMjSNbUeqv68CLcP1SWzLEfvKOZO/9COK2eJxw7VecNdVEI9
D6aLzli0Qc+vTATyDJV6Zym5ZwgR2834VUTDrZrYZkVG3rFgxuxPfvlQuBqVkxc7
NyW16rZ8/nor3xVO+17q2ZHOTQXV99wPrVUphw3PdbPHuREYzzHNIGXlcPGXpDPr
Xaq+tOvkh7ydrZyqQ0l1UA+IvNmiOQO5ZHcs5CZlaD3M5zsmxeSBsMlv7N5eg3EI
u9WHCcafLTG8EohcTfR9r8JahAaCrILprfRaaM2f60WF1W9GmqE65S/sP20RQYWY
FMm8eud6RxurXaI75wnTuG0nNhuVNEdHUYZYWFBvMBff+b5HxcuSP9qNqcmE3YwA
tlyWTBva8Q9GjFUjRNttkvawvXho2/RiHj1rsc6x4xJ49XH29D7807gse1jPxZhQ
i/JBtrJ1SEiGDNWqFI4zcqH9nb4PLp252zUd/jIUR0qrbUTuBDvYVy0z5s7YVzTZ
zLueauOHdCD9aCegvPN9LNO7xn2vsfwzHR6CGEdpF7StjfTt0X2YYTYVbFcCYGVy
AXJ3wkEdvwvQDjXOt+p/wg1cKVwKC8RNkT1d+d1m7CjhrrirzLLKdnWiRYT8PgCE
5MEu/7xMg7DXfQS6O4w9aThRQ+nWp3WFFOpV9VO2b9lZICfCk9WpXM/Q//uv6gx0
oJRrRS+UkYNywZYCY6gfpBYFC9MX8iJw+M22ltKEeMyntCvkjw4WJcaKovMZl6y6
eESJGdTAOYBwzP/SUDKrnKfBJbntTiFn8PMy4Aml7P/AvTDp6rQHkAObhLaA3HGB
VlsCrds1dyt2G4qjl6QLJeUG/sEIFL5++OVJOI6MDeDdNmGM6+riKKp1vWSBWDZa
V+0TDNQnzDUkZoTIgKpFMfXvz0iq4KmNDOqGesmyYvugBZZ8KdSXy6ODPrtlA6zm
u6NO5dbuC2VPpRbnE5kj2s2V+OYQDrM9Ei2stgQBneIukxRkqMZGSkemKs0OgYP7
vLkAmiDZIQ1bz2GzC/zZgbyLkAoaSSQMXaOXlSHNJdZKF6xb3cpx7gsCVB/rAEUr
PokKoEeI92s9bv7rxau6yACxU2KQhTSqGFxPgtnnGLyE3Oc/gyvJ6uWDfwKpFvVO
hYtGlGndqBFgp6p5fXWQiZoysmRdi+50N+iroGUt7Xj8agI8GXGjVlzwRjY03Wdy
idIM+9wQAlijwXEJ2XVQKVNW5OWsvIIh9P9pCec4w/DaT7NWKxhH1xRe6W58N0sX
yBIePrbdB3ctpco9GhAWYSbaCCrr/BcFnKE8yUSkPkx5/AxhYzerxNLdNiUMjofw
zdby1ge1/HvTUzFeFHcAJD2LEv5dbO1zpLSugdp9NORp7mont8AmLyxNwxcX4sHt
hlrcSJV+w0JqEgffnf/2HoU0hAfyfipIpK4FdxbT77QcRm6DbkeR6D3Qge4cJsBQ
MG6sc7VHFlvW6+ycRzld6TQJKHQ3AeQlgrpA/C93QBFTAc/qiPrTO5+8ln2YB7E1
3sLW4oWIIgAUCqt5hXJG78o2/VypKCmRg4dXX/OngdsWPFoSqVntIm3d7Q27ec4X
gS+YGwyMde6P45jYDPhv8EzjngdZfxJ+BNtwrkJ79elvenmwNLXpCqONqI0FLJri
3BR28T9QPWMBJiroT283mozQOfigLfZC3/dLuS0CWMYrJpkD5wxfgw0/6wNBZccg
`protect END_PROTECTED
