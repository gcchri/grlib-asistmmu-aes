`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZrQGVKanqg4EvveuO9UxyYW1R19RGTgdAhws1jtqw2ks1vgdgIAv1y9GL7AGTsus
qlK5+41Zmqyt30uWipJw145Xsf6q048gbJ3oZL+B4ksThN+xyB4MLarAkzCom681
uVXMVMYb4o2ZRmciYJj52Az/FIiAZvMZ7m7LY+ov2n4WmXJZ6rbMnA8A+wMX87ZY
l/wCMhrRUpIUqpc2i4KAMAdT4ror4g9IsoEUdWVc8vTsNaDaLyAEtFfKuXC33O6L
ZpfY+abRmEtcdpyO/JrcZCy0wV51GkZL5J92dXci+SDbh20zo08MFxN/TFuoViZI
r475j3bNzNMWOUGfqGz68qvdF7S0acy8++14QeGgQLEgpkxaiZzUTA98zDWaKwdO
LvD4te2oigbAlrvOTU2vI4BMPwQmeADW7lIN+mXRPgb5kXiRWMzdfwz36gK+Zh1A
wLfc99QfXfEoYICQQqR+oEGCeqemqHcw6BU7L33uIwzsRHW8XGeNstCsEyyhuzSx
`protect END_PROTECTED
