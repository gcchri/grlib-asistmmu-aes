`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UuTB7/m0l5EhBkq7LIeb+QMdCCZF7KYAMEeRmnSantb3/TSakxEa/fhDAC7RNPu2
RVKLTMo4KQknaR12MEQNtkDULK3nqN0oRM+fOlfGch2+qX+WGKj7geEym5iotVcl
2dnnHkKpg3gXZAr+dQQxYtAal9+HeY4SbukLIYJJlXWRayL7FG8xx+BJieCszAub
mUnM/2cNbGopu5wuE99OmZnzuZDDNs2NrS+4Sm4wwTz4WNq5CQXROJkyB5xhHjpT
FDw2b+Yhd1brtYtqJ4ykW4zFPvLwRhu2ZjT2qas2KrvOVqTZHmrT0GQ0gYh/KP2X
MPMGkXeVxwnpJKgYGsmi8kg7LkojcA5Titcmpy7EyLk=
`protect END_PROTECTED
