`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D+QgbJOItOKSejIGfYdEXUeWUNvnjTVKCUZbBoXEwUp3+n21yJsDkFRgF5DTrc3u
HnPr7CQ96q9BBOvpBGc8C7d/3GQ0BG+QvD4IyEfnQ7f7v4h15U98WimmRwhQ0ELE
3jI5UEwfpQ5M76DtGfocDxDwxv4EkjIsOECjmxQsRNOdsDPFVfasyRxBg8C+CTdX
NYDSUe9xigMuftI/M6xyzRuV9fTCtqFVIugnsWynw9iH5EyWyHCpa4nZiK5snVow
u+jMeKPQi5j2ceM/+MDTsVvii5kbH4AUYZJL8dcwk4g/3fDnfgN/ZLDDnuXHF9kX
Be6E4/1ITuFirfSin+dHpVINuaVUzww/p8k/0Tpc8N1QisQGF0kXujNSk/irR7nT
852pl+M7S18bzotye2toIA==
`protect END_PROTECTED
