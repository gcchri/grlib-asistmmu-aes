`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
065Lm0WL5koYsVNjq4zaL0On6qAH8kNmMk7EReUjjAPV7vubvJwAlJzMnBzWUEph
N8L8BmI7Kze3vj8FzLPZQjp2Z0FUhuBgtSWVSihyyxSF2cPfP03Undrxx9dYQ8L0
WH1HjZNTlHlsSlTRem4DELogB1tiDidKnMCTavxpmwo+X+g6q0iVDYxui+Q7/4Oo
L2qTCmzUyA1w1wv6SQcyxfX3orLMntXMzQCUv+mGrhPrCsXXUfN2WgYLTEXyG0m2
PFU8EUbi89B5uTp58Yp+xALWo9XCdotWGUL0ELDCasbbISha8JBDnzVHbN2mo9CC
Vab6M2isPWrZ9FGSkBSWpeXtMp6FQ/ifeTIX03kE8/GJ7btC51G4VnukjGsFRszS
IuEf262fjJTm1LAViwG4pxKwrfYT7EhrJm4kgToxawVew1T8tJ1NIyzt0e3yo6Ly
73B8sf+RzHq9e5U1V55lllawVnYjDwIfK8oAuRhbZKsausNlNUnQDFlcJOZkXwtB
RrPAU4JcYsv/CW92eHpjjEDhknpnXjrfkLMzZIMADnnjuxUTUcNiFWhmKaojT1BQ
/w7WPDX84HF/f3hcQTci8c9nHg+F7Kjnsm18bWu4BTT+aQ4+UCdi/FFSnuq6bnJY
HyJduvHH78SToes2b5nYiq/vOkwI+LHHywvf76dNjMx/g/y0lNb9Ps/4M4D//V3e
z8LdmnXO6vTckhDhQf+0B/v8IYVB+c/iulZVlQJv588JUTO0zoc2pcNRKiVGqyDH
c3OGpU+NCisUk/gpj+hkBEFZC44UO1cxawBdzVogexw=
`protect END_PROTECTED
