`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6lg9nYtzOQYlHMuNaQKAU6tZFKreTx2NGBRSRlRqlpWYOGTOgPc3hHpWoMDKL+/u
yCE+T1lXKizp78u1gBCj3aUywyWItyMJ4qtJNjnQUe5JUCpgDKYUTeLFNl4h/O90
evBABXW9oaNZsD+WrHVgsx4kP6JKhy0xXRw2d29AVrK5u0affhrqGPu0reFQNM85
OpT94W8vKKLDlAiEsIPVf2AoIDjuqBCa7LDB5Y+kwvHtsv+QUK4gSQpvKd3/vHPW
/OkvJnRXVDDJw2V6bML242JfCS+TPmGpBZspjsZABpH0c5GrRALlKQ41+lYnsjS9
aCmpD+34woEf8Cy31nwJASNDDGOrIXRn1iTkYlV0ppLEWPwUyZP1ZNqqq5UVwmdN
6kiFOLk9m/qtX9hi1hEGjg==
`protect END_PROTECTED
