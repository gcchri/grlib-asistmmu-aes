`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+k/TglNSDSEkhI50DOgw538Dl5TaKfnyHWtZf4kvTCEYUPx5u+FdiSSPkYoCvg1N
fQ27M8YMZKe8jXxACRUMHempNctyA4+SHN/NQ/Kxpnsk8aBv0sEWHxP/y0Cf1+W7
xCZB+oZuK28ZFUTZEzXu51ikr49XpDkChs0jCy0Pdr7QMDnp2x7zWHs+t3pLOi2U
hs5DETFq6SUW5wLsF8yVUpbYT/iorlskBNavH40qMuaTbu/RFUxYMLtE6wjVnZpO
Tg5QLJRhgWAaolnDEXY+ZxaP8LfHDmiSM4zudcDfpukBTZyCNe19xEfGKCTRVOB3
utiYz+y7573MKrt0oP810TSF6qMZvTXBWzxW+clU49wCw88ggaJRYg7iQJRfgnN+
`protect END_PROTECTED
