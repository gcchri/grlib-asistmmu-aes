`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/xdq8E5mgt6ZC3m+joCacyajS/hTWNjPGvNw3gq+P1p5moJqOojbd35RRpFsIBGl
JtVO325X8GGud801Q2LeNzCYbQ5LsCw9fAlwq3XXG8YSkCAqMXCh6Sezehys7NfE
QafRncQ0V0KvsG92Tr1/iQU4UKo7vOlL8TzqjTkSRmkekz1dyCFyxaG2tWyprUX/
A2YglUMrevFZssg3FoPuVnzjQkyFdCZk7d80bEoPr1adRDlHJkCepZp3pVQ46mDl
5GJdo29V95loUbbNEHJr+NnuqlRJoAGC/l5+5KHJwXin50MrP1vmSu8FUlBPO1bc
hNmcyH4q6OaStXFru1/GRbb8TfZom2lsYGv1invUlnb145+6BHHZfPD/6IJBsqU+
5EV1RcSjn/lSz9CPmZ+9n3vscXMhdT7+Ph4YzjNG9ToxzkNn0QoaPl66/eK9DiGR
`protect END_PROTECTED
