`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vojuQXRGaSmL2QqiryxiwCwQDxAjOcU7YkTA8EU4NermZnZq66t8Nky5R5BYscIz
5Qdr53udrw9nhJ+3gj+rXnIHhVVJvC13iRl8+mGc3XK2iyUtUnnwKZA8ACQaA/Wh
3ELxKzUhhqnRqx4GHHLedsGXyAKDnH6WSTztZmdsXdzwMgMEOjtzl0jMzfOTfC81
2lKEXLyxZg1GPd7vqawpR00t86ULpuKDNQM5ecDVI2O/eHJvc9vwIHMtV1XPGGez
KNjoeQs/V78wLS3Y3oNtD+EX57tMpQhKi3Pw4vNzm91+dRcGxC9oGj0t2kTDhfM5
Qe+UW411L4v1eOgCqYYfIAGiTDVT28Sq/nzKjYJSAhYR801hpMvKtw8d3n/YX8rf
v/m+s7akRgAj0Gu/DqwP10O3li4wyp9k1ssW5a50iG6sPuF/gJutvGS3pR8mPzbt
/tqPzjtwoJudPQXtdS0W1BDLn/EUcQksWp47M0xUi04o5Rg65iaM0G69jTNfx0VV
3PDUn7wcsYh0TS+ra/iucI298NFLszrGCEURfDicqcyywyQidNE7WPDHU1cLHyEz
Lq2uZSuNTzL7EjUgSAv6808DFgcJ38nwqk1lLoYeYwf35U3OCwIcd8sR2q2kcZ7Y
X0f/UMKsiV3IkR2UEf6k821QaQRbplAC/KQ4tjrOM4zJq78uDA26Tfmu4g+PdGkS
uiwbJldcm4Zu6TKHg0E6ArdKPPFkYL1rBKflMj99Y14QqPB4/UWGJYeKtvBaylZq
zlDmrKKQyqXT7CbriBpKALVvm3cwQALVFMQ8umpibbaAPbwWK2ZgTNRuw02YXOiX
CqZtu2V94KvGrJV9LBh61FRIc3IJY04gIxg2Hrdo2ffUztt1OZz/7EaLpQSpv3eq
aBwLSEf/uLrClX3D6B2f/vN4VmpS/rgKKsKX7OlbIwOUx0ycLCToWwsAfBKXwpV+
Ynsb+DPwx8mB6fp2sPEkDELYBSiZ4IPCCZUmCjRMbnY+JeO7XTAueDny72UlsyKF
`protect END_PROTECTED
