`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qaeFK3YF8TipIWYHCHUxYpFdTwcuepCsZvz/Ft6Ri81T5J3i08+Hr9ezzn/H959f
6EqRh4OkR2bXuPVFQ/wh05w2DSl0kFQ796Zt/4HSzBcs0eXMZK/nv8PWwv06MRZA
03aXe338sA2NPAG/x3I0G2TrAhWDsrb3v92Qb7uqli+u4zHw8NRwKkv2ODaxZysC
PAuC7xJfpCgY8cM8lD97kIHnohlxmssS6f1el67GOsV/5fro29HvglPiWAsC0HcM
MiapHQPUz+/fstGsYtxvT/XkLVfwv2AiimHdmHDqDyQzpnJVqGJmzJUMgxkaPXIO
bl3k2bdYLzEUqBkPKMamzIDzWjrxBXtVaX/gwM/h4h1A4IYNz5MbdXgAbIE1SZ3h
GPBeSxGCza9NuZ/pbipxETORD4zZoCkreCv42pspbjDcvjV9ctCs9iDllIHysqWn
WGw4/RTNJQZDpVLJOXfiim4JHp/N5bvu1AxNUjEDcgfde0o06AFdt+50chV2ueTX
sXsB6kDWhUwa3t2YSiGD8zw+CTkIi8oEqt4wOqXbPOe5zESSoCTu5c1qwfzhfp9C
7tAM5tBD6t4Lygt8bonuF8VL3qo1+cqtjwoqNRKQm0eLUmfXN0bUrswmZRR1dyVz
E0Q5OB5qiQCoufjITqVvGSh4FqIY56NwEIQRaaxQ/+zarGzku0pb/aGCDuLAxUov
tudPUolfKLdC45oek2DHKzzwmxZQu/c7Hb2JKVxofr0L6bxtbaHtj5aSZBcf3DF6
fVzaeg9ED14JDY4KCulFdbrutOz1WsHPHLo0+WLdYrA1SFa+efcMn6D+mvY9ydiS
GEF1fFDH1k82oY8wnEJBeMJ7Ac3ePKKlk5s+4oc7PLyds8mOLGpS1qhGK/hZf5Yw
JGONVP5d5W2EQcx7o2yWYHw4rAJhIfT54iu9AB4o3mJcYoLdzbpMbnjwn3xbKhfv
F2tsX1jpz3lctcc89ghVJ7u0GikBq1mOcCs9CqvFUuCIlZYSdifhr+npv76FsBpU
atoicT6yGqGEN8w49nw16IU8WnuFTXJOp30c1tTmLHwy6Kh5O/1SAcyjmTKHYJ4G
1VHfvbG8RLwJ5C6IHLMgEq5Wp8bR47xc/iS94jZNjhpX9karBXqlyzKt7ABao0C+
`protect END_PROTECTED
