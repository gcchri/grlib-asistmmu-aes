`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IDe3Q9SmCx/MguraoOwbOOdJ6rFWlZ/HS+tgVXCZf3RA1FRvSzM08D6sS++yRRn2
Mx5URKTye5T0UdnW+5DFmwzzhkkyxJFU47+F9OXSHZAkYHeiUK6csDqm+yUDa5Th
eKcK0JDIfaH4SL3KtBhuNa6aw9DyeydGuB2kE0dHlkIIMv9KNF1x3Jurs4hhAivl
2tMsnj1PK6jeOd5Fu57k9SmBBOcvBzlxSso81lGXvhbkHfxr80PEefpXCHpcNBlF
oTeDUf1MAbFhSXUUmk51sJB2fUH+Bxp3y3oBC3i0aJUG5yBCyjBpsb3AvgAhw/mm
ozf+koRjx168IbPHvQ4Ux2XbpS/AZjjACdhPWFBYcgPr9iyrlrDEFEHcofo1i3WO
aQIdBtgpy4diZDm9FsKGygZIO8PBUhUTjFPkc6U31naWUiBSiTnrKOzXKZKPUF2a
Rlz0Ix1z6B3R7OT2Z8hysH7o04bWRyLCFDMNHkshJoQde1lpd35QzBiua6snYdZ3
TL2cFaagblQCUssKhOgieMD98R9aULkO3cDj8QoMOJqT/AM39SmmpG9WEnCn2aw0
+Q/r2cW5q7M/oZPLjkUN+Ht3D64IV9wkqQ9L0EFZ2Py0X+IDxmQJZsbq6u94/d5C
zhNmctSdd9Vga+Pa1pqwuNviOZ9hmYaLhL8iBU+kmYRf1eQPUzKDU+UXOOy7CrSp
lgcJP50VEMxzd4ILsTJa7Vup/MPCKZmN8jt+vdADhm4O61DSGYEgGcCV0XcQV1pT
/GicyLIoQdK5SnjD14gZny/vprN0XxRbP2ZaaHwAfnd7lrHD4GGLmIsG96t/Bn1O
Xhe/ewUGxVnjtIFIvekNL26Ym8H3QlHjO/WnaeZiMZ1Jg4R8G883yIlKayr3Fwf0
KGZbx0SS9ZUZSsYILQ6q3gX0HXu0UKsW3SJndD1kMLsvREAO85KRo05qUC313SfW
zPXxfFtKXv8BW8EiHnghEnrSOsKYVBKVhCPktdaLzGhxe16UM0XLlWfzUkUrObX6
GvuZDDSGm5hVQ4U3drgB4+5jijMJV+nFBME4gV2UKMQ5fu1kb/aZXHLpZ2blzJbs
h0U7Cawcz78P9ejcJM6ODUDCFmEo/a5nPpnFgBgH0A2UUI30+qr2730MHiAhFEIq
8Rc8hDlRf7o1FDUn0Hn9NLMuYWjGVdzQ3EKWFFhcfMBSUAyhRxvcmUO7ZHerQ4gX
Biie1D5830t3E+FVUQC1nYY1FRDNzwSQXHQ1UP1io8JrJbmcVKFAi+FVeVD/31Iu
RrTW5I9W/n4bWGZFRbbM1gRzRKH1X0MsR9uFX43weTXFbAK8ymm0kMM6FjMMY/wG
MBe0707Tn/CipUQmidDQM15JGFsKJUFsD4BPx+AydSWDkCh4g549SWYbvwSdMpFr
lcuTAh/VkBwml93Pm5cdqQjH2u/ftMWEEyfZpOgBcYQdaKqtrnGqRrZdhIFSm6ix
SuPNKyZZ+74f+gDMF3/gT4PeO3i/7r35NcRO9PXBdUHlASAdH1JeGgZcYxLqLFBL
aj8NpCy4wUDW4p3anzfdhS53u9RM8fFJ7m2uX4HpC4fDzCDxHxFo8McxTHmK8xh+
7boLmS3OZ2vE7z5YXN8k/VvNLXbbZPkKCx0rBMbQqmepim/z2iw6qPFRDAkSGt3G
PVhcVI16LgThmc+bbfHIhy675I8cO6IM9zcde3zf48cTVvH2/nfI+FzGtBWrH+xE
qJHjKulOsQSzvBJKn7d71TmNGYThNIOoe5VAokwpqxrIK+sl43a6DwL3Lt+H8ooL
h4Bm82HVbFQpOzqKddyd6xqz86mGYM7Flbesdt7iN4ixBVLo1Nz+khiO/x8/MPRs
ijeGPYnkX3oql/GGIvIaKmGdYOJv9C3V5H39qpMRqt3oloDAmphGvjCtsSshBXIO
L1tD3yD5i70tFV5lpvdlKpWG+mtb8bBxKfL66BWsfEn7nC7AtMdcAUgPDY5xkJV2
goPtPv7wJ7WBPhO4m4039YoPWuOwE1jE0ic6vRX7s6QEjeByGvz4qDUu1TJmlLAW
mNiWY23Uiy2znHiba4n6YpiMH0gPfivNaBrO7kuc0GxoOlA4eaUTd32e3wzZeMga
6fwwCNw6Lg1zRhpStY1XqXO+dkuKQOdnDGedxXJfFdmwDNy1n33/WE59Q7jCnmrW
5USUHJ2JvO4JGbK8zqdDL4FdNBfgQT7P0kKCKFqQSF44xUwaRFgmFclqYw9JW+QD
NFZsHIkub1n/03p68p1J9L2r0PjOMw65S53HWftuQ2hHspt+P4MaR3Hn9CHLHzWt
Mt5qBULdiGoInauJQY2Olqf5ignXgY/riCMYYAC1Cp4rppeMJzoMyVqSNnEwZ0z1
sXRz8TFUxJMzSokRYtAejVRwO5gDHFq3zx0Dn2+q5pX1qkx8jprQRVMFe48e7s3p
U+Gfjs1sUZ/c9zUF6vjwS5ENTGydsjDnLdORKY8sfVP0CSbJ+JbPOAA6xBzo7Es3
4NWlGu4hzhZsuXXaRE023Ls/ARNOAdwSGpqj87oB9JmFLSLEDXvxcmiH3N+LE5JT
wD2jtxnHTu/KFdLtv+5Iq05JZrY7YPBSUA/McwvyOhzz3c5rXm+nqPv0DP+3JMTc
MTzuPiNflvdrJ4PsKZ6MW3MGnp1CFZVI4kYWEB5hIMqA59fiYTrPubs81YQoT7JR
9xt1Zznl7c5VDhEnxj/qij+UyiMVkMkBa4O3sQq6zzAIqrDcbAlOzxZsR4XumyLh
grPe6Zja/AuPGnwtjKfS/cZQCO4SaDCIPqWP07nA0UUchHJojQoRaUCvcaWdTot5
1tTR8UoB353WrIy2VWi8aN7GflQxkRVmxCM/JzgKoMskMEpM4eaWjC+6NFryICMj
tZs+dmotuyQ0KSQcwj8abYsoT0y1x+i26ni50Ixf828=
`protect END_PROTECTED
