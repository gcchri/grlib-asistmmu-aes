`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zi15EW7zJkO9o+cXvDWRTMyY6WvmDteSXuOqa1IyQJAaX2faHfPjExf8tDStHVm9
bQpwU/lv/s3Lqb08BlJmJZJnwynbigURqz2WrzHezNecJtdGVpZCXNaKTPSPErrB
G/T8GdUhYabdj7pNPRWkwswwDUsWmjJE05PLCmhUh6jU0GMM35IZwCvaiL07rOSj
wxr0tLffrIAMLwTkBmLxSsLOLIhruKR3u74MMT+exIJBlgC1USSvwqPmWFCSMpUf
EC6hmUF0/avJRNYHFB8zojv2MG/s66azQ5YU3FEBxhYHW3cc2W88/8XBVceQZZkc
9v80AFN1EArjUJsD6uQofkzVlYpeGDtisjvjGLC8FMcbVdnSjxZhh+GgVOB5LZbc
cebcq7p+JOruLPIfTjr9o9kP7mzgh7MutennXa+W53nKYxPHZ76CTeoxESXpOsMn
MoViwpQC0KXffzPHGIF6jxHQFiB9KxS0ukg1L/H37MwDKw3OtNp4zypQ91uLVzLU
RQI/XGljwDtaiwG/enNOml/8Nqt8qVVwA4EvYfqkBmha0JdAe7OdwyJT7TW3WiCI
zODReCedQ8YMsYebA/u5KN3QV4/o42ctomX93x3df0dN1iCVaQTVV0Ivzqf/SmFn
efctGvVvAn4J3p2a99bwxbbQkteAPCXPnfXlOcVbUMN6AoVGu/feh6SfYMYceSz3
`protect END_PROTECTED
