`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zv+5FMGHpoXTVlaXEKTcNuwnIh2flQDUS6JgSoYJfdYZZXGI6hCoRcYX7GN6FjMb
rGTcdqsNSrtLA3QDe/h/ZJlJ1bPUilnQfoVewX6YfFOCugGyLoJ2buIyU1jN9rGP
uNtUtK8Al7H2CmmHYoRENvWaiWYwgSPh1bBBMgvISW/uqKH4w9oz5J9w7K3R+vj+
lBFDlYA3Eefo/A2750voCs+jhA71kh4JbqICDyuSrwzTNtzjxTeKpFBs3mEA4GSX
DMd2bqJxLmrPwdVsmy1jcXnqSr24em99hwqgYbT0DTrpO1qfe2zeHkpO32k/TzRQ
CrYUp23RLWGVVbe5FNBqDr3OFjp02+iMzvHNrTZdPjg=
`protect END_PROTECTED
