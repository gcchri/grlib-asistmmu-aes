`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3uDEwkSz0iTplln0tT1sHLPsZLYJ/SyfErvE4jvWpNOY2clpBPQ8r4Xif2zcRol0
E8jA+TWaOvueC/R9j/19gX8WkaqmhSubJcRYu15Kg5oARDlO5icyNfR4fp/eMOyf
1w0AUs7uvkt6owvaLyuFveDepxUvhzlZhLMASUuncWGCFTFO/2mwExIB7iYqKldk
WPkC2p9Ef8+Ft+Tzc8d5oCbg9wGP3XIm8Z1u21yhYyYUsUj7SoKH9u++tK+fKYXM
mCARyWLgmM0omcX9lsEykJXHEHsgDuA+5MycjlKE/nYx+xlk9PlTbv64Tr0e9MYk
jvxDWcdPgLl2w6s1IxLzH15lpGxGjP/beLuqlX6dW/BwNysRNogxrkU9V3LqrfCy
B9jt+wqTK+MQ+DoXh8tpzf+OEkV1MESGUdKdjnAqTXwmOAuzfMIO3+y9zGvxOq60
pLS927hBMJMeLcNZXaexGttjZu/LInh3kw9vWYsCvcpjgI+AoN173CKZv/yvPJ0T
MAWCivb4pd+LGM55c1jnuHxiumtODCD+u0fM+Zh0njYMwLDdxo5aM8SUEIpVIz1Z
K9kBSs07w0NGEeBs82KZMWED9P49EVR0y6pnOibv/mvCIYkBh2AJismvhVQ686GJ
Q8vpDP8vMhTLdXUN3pJBrU9vUJfy69tiKKAaKBh0O9jMYLdScv5jU9jlpBYu0eSq
/TqjjOzVq5X3NLU6aEBaWi6HinKlW/46b0b/nbdxtnh1OdimCrPVdWuplUS85aGN
eAJiYiqjJw+pJj0/ISSNI8B/6QiaqTxur+/tNCFUDU5OozdytM2v7SiTgt0QJpl8
fJcIm3Lc+UOB66qAbffRv7vIoxKRQ9T/+4phGW713TSvn66yd8lqixzULa959797
P84jRAmH7Gcw3Xudu8bEXBQE5XsnJV76lQQZBnoTnI90AbMVj003vB9NIFjt6+9I
fu/sMzWbyjbX3pNiuou0MXR2xlpzB1s0/wRXjGmqB3A=
`protect END_PROTECTED
