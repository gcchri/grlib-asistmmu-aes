`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p+WwzjLiBJdxQxOXhcy7vM3wUZH6ewSOnA0+9Kab8r+IUdnFN00hTBSlYHWUqvw2
6GG5hM5yxsMOIlnPPVxlf3We+Uldtklem7NNADFFLBRv7Q8zK4j7DSVVwX5Vlgzg
QjrbRXNBMQKs/P3E/ylVgbHWrh+evXTHXDKYw4fuWNb5Yw0bJXRk2p3OzvRr7CSI
HEgC5ukFuVBspna6rlyr6cTiSaFVEBsG35cJCrD7x49S0wH7AYC5boGX3ilE0Tak
K4ThNWHL7LfT5tv9q8vYTScFzKEzrclUHWVflOTYzvO2G2hunCLM8Ev9vNNO+BIG
BH9NQzQQ7nuMwKFN23YVEJx5rgDRYuqvvH0+A5OvOn8iaRzEm9Dfwv5s4jTNXKM+
cN3/1+zKlhaIZBGSHtBUUqoDYqb9dkOXeAWDzygksPtUgW7QZo7X3meGidtWMDQv
h0DrAV6hpegs8P8HlSs2jO4v/NJu3tpHgEQB69KZTuf51nWcDCENeWbejoEwCSdH
jgIutLcTAwxfe/841/ZyjuYZJhUA7kPRzDWnDbFpOdldvm6yWD/BxzIq7vIiMjXW
tH04igStJUZX09u8nsMhrCdNKarJoJ/NWcbX+5SZyTsM0oOFX4eS+qrajD8KqZyL
R6U4sqIW5RndLE/DGGjLD0q5zLvQPAvKFqYxRaVM9Lhv3OBwurj90CalY5B0SkyG
1WCZEFAEAO8qjReA3ynfA1b9hFaNcUmXV6sFSqE7paUnWcRF+d4zWoqfk+8wP1qN
lOcAOrex271CNTW1wVTRP8zKjeQHUYyzHdwMbeM/VDGSM50tWMY+3MlZ2btq+1xO
8BCB//IIDI16+5jldsjQLHCQ4IbQtngpdt7x5FJPMBHbsGNYfTEKXNl5CNu+B13m
EAUsQkzcFc+SjSn8ip88Sg==
`protect END_PROTECTED
