`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YnCHOXJkEqWdPeSdYS/c2K9oAYZ2gJktmmfTQzyhSjK31dfvVhcrhaOvFedqHzJy
MgqNvpOCf7QCBzulE+sb/PQ9QkHkXwG71mgv87dhw3qY5pg+kulkquvYm7QvEGdI
pl4Nb0+uFVW7cXOViR46TzQ1Z/FZtJv8eopfJCScwUm4CvQrnmvugZBxCuGbHPJB
+fwPiPrcYPPy1tVYgiv/p52508ZwXLq/Q516bZV52tQdqPsxoG64nnVfE9AllsP4
j2UUuiipIaC7lF2fr09nw3obDt9d2A+FjnYNnpOJkP7igckwt1zVF12o5sZkxq3/
nFpkHr400BQq2C4dFncwmTj/1AmvEQjzdwS2eDmBCGJKHdGg1Zbn+gRZ4Gcqg7Fh
duOZgcAm8w+6/1vWfJkG1n6S0erZMrpJTEXSjlRROao7AyREAW5kvdQLtt5Fi2FW
7o1OAP5yiDy970A+i/XwNGPlk5RHHLkbBblZ85tQPUx16ywO/5bJoe11ydJsSBSl
9MKegfOrtkauYB+OhU6flR2PoTZpbgptmYYuG5rj5XIaCq3Qaez9jYH5KOwhgPBt
t6alWCgUuBbJ3Fps5RGEIbVHUm0m6Wty8Iyn+b8XbNI2gf12tBrtpLd5rJF15pfM
RgIzT0jKbUtYpJZKIy5d/8+Wv+uHEFhY7JBU6ZknU1xCH29Tg8M6jGOJtyZVAn/h
TtXro2U4gGNdcnPsQvhlFxtnr4MKHjJTy/h4P2POOb0WYItY+DGhajCNmSbu8Xr+
GznCEZJ5mKXbysilS150xOISe6M5Vvhr+s4SjANj9NXrRyaf9g2SxroSfte/MsOi
xzUVmSwEOljDiL6T0mnkD2puUh5Xp8Hsg2/WParXmVgycsGGjKl8UpTCJTN5Gju7
pfCFa7kH0MZozLi9zxPMKZzBFqr6rxmfYJSEwLxMJoY8ShN5SQEI5m5YZ00etJLJ
z4pNiG/ZDRdY17MGa18Hdyzi73lDlrJzRxx+phtFC5uG5Mjrrz5/i2q5Cy5CxZYC
`protect END_PROTECTED
