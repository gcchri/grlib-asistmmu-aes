`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6UGqTRD4DgJxXicTSS70JfVQwHm3ZhDmK2Wr42vPHGyv93xkMbptWSTLwCn7eVC3
4N9otpQkVK67mL7P73l5ZLVyJh7UKGpSCpOOZLoajDEewT/2Ew9fSarowVCdBF5H
PMJLGcpZIaqvH0asvd/O9bFEwkyMmY4ljl4B+ElAIWNdi+deyVCNb9Cg964PTpFq
hNtrrjWbr1V8XLrL6C9ErJRS9JRJakXwIYBM5yrz8uO56LaP4wq+8v6GO8VfbrYG
mJT5ZcTRIU29KXbpGZSeriKWESzqwZuB202EeIJDhe4NP4kccUzc6fItf9ppLG0u
nNw9rhESQh381vqJABTCS4QE76ZCL5QebVbq8ee18c0UcIS53vf5hxjBMIanDaCF
dw+Vd+uxg6G/ivnffWpojGqzGP3QaH8BkP2fDQQDXK9MwlC6e+RddqlRyLvJGmUe
`protect END_PROTECTED
