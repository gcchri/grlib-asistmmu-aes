`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iWud99jTw6cMF9BsfkwPSa2O9i43SDDJ7X9WpG7uTjT8ZTppQZiEc4ASfNzXcCRG
CUNHTokl3O0W4qZaFZPM8sMIvkwhnnDLugnFZfIA0Dsv1lIvi95OMjOMWItFP10g
NkHbBszimi3UPNMZI0dB7TliOT1o2+nx5fsBHx5wG7oSgX438JzWOmsY7OYTqRY3
MYgpQVIOSLSJkDLZ1vF7Ej0SSfTSgBE/c1FBXR0vG9ILDUyPFS/Az1sewb3YCuAq
23LQ/9NSGCgKmSiVVlYMLaxtwW8vr3h3gbSILEpAtYF3OOWmhr6l2zrnAA/Dy6vV
U3XztTob9g8+kQOsNOVbYAiafUZKGTWULR15LbTdDrs/Nd5cktscMMpYal8Rgvf8
09zhc3Kc741IeAPS7vwvKE1RtYq0dVdSVVazRKbNKQ8jF2gLdn3FBhkjMiY2g8FT
`protect END_PROTECTED
