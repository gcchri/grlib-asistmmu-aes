`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rxa6KDyyoK0RPCdIM6KRNQ6z0lyp7o9WBDFiX11N2k10o64h3LSQcBbWOrhxGAaZ
LB7GkwJWXbvRlH7Fcr/8y4tgkGGoDcwIbEokIuxezi8G8h/ZHF8W3MI3dJ/GEgxO
mkEIJ5tt11k9PGQidrjRjEpC5wHfqiqOwM59BPrLW7AeP3DPkNZC2v/9L85D7yHx
A2hMLyOq1npf7lGR04/tPFECnk7Fo73SfJgX1BlQGQHEAGjjIpGAXrVAYJ73QmCU
R6aiaLN3ZVUcaXi2mYubpnTy0ZCijFJ2SI6OJjQbCrnBaL/BwAJp2SGVCB4/lxSy
aeWdvsL9hDd0zJlXEv6SPfIMEc7qVDhyDt++LIYUKkJySzKNvT89e5KZUexL5vw1
wPlZZK3kuzorjR/IfPGaaWGQpzX+JFCK66MoFadTNMdgn1M2DMejvk9g2HjdPIKr
iGSwPVM+PSQqEpvG9eSrWyNPnS7VSopsDQaDGYhoPq0ughY08XGqg+7gVnLqui2c
PXql5OTVn861Ez/hp5AD4anDuqY65jPMwtYU38bmmyVhxO9ejqnKkxbMBl1QrvVG
EaaGjpJCi3jxgRXiUdGZuqKgphBVICFzFwoN+/i06xLe7aOO3jkLBP/SbHkHEVHE
hsbV6CFfF9vPBCsFOALVPLxDP8jL/mtr3PLoPCmR61QysL5M9f8MbpNopQtzalgQ
wuv/+ruQNzmlPl4XyyT0zLxc+Aur+R98F7N7NuzlOLdDdS0CoK1ZTjM3MfXf48Ye
m2bLZeR1kTqYlB36ukiZR8X2H4jPYUFmRb0UTb+Te0Qpu5PPIH9+xY24Pq8cOQw6
hXtbcNXYdxfU9Ga3YFB+oel/GshzLE3LaP1PCFwlBsJPWxZ86OWA6ngOMwqG8oG5
ToOG16XHQV5d3R0tFw0GDzhIDllxj0DsnpWv/Hj5jWlgzgIZZkT2vbkGZ4W7Lsaz
he4xCaETovfOi7i1KMrU2bbjBYW/q3wtVNKc73JLHg0LCtd2ZeWR/nWevktCY8WM
pAP3UKPtCSLrwpajl16hzOt5J6AIQ+xhc38XoTKPrgSZabzdhPuDPioCUfJtOug4
EPe9ex/GDl9mSPv5dl0AcsTVNWbKE1IR67H3fC14sH+jW6P9tTwuF4AaH/Sc031W
YTgtoORSPcyPvidXgYXYVaH6//6rsxYCTuEazJcegUEuY6NzOCGL4FWrTRnw4TTH
U206AcfvE4w6Sd14u7u3YElxHwVmBOM+Rv1Duu41SxOXus08QaKjLOM/xxXwL6HL
UBKOyaBXL43CNd4Iad9G8FN5QpHvItpxEpPRjuVA5AJXUZr7Xs8OrK9IwLfzCnNn
x86AF2foswghgrXxdzckV1c9sJTuvb7WQYaZU9ugYDU4epVUujgEaGvJDxghPFyZ
CntIe7o4d1vJqFU0i+zv/M6sdjuoMTav6mEKxafapFfLOv6/YLF6FLOQvmAn7OM8
Z9jEPBd4orgqHD8XSFoIr892PO6388vBg1jsZ7NXZkY3EgGo5Ou7Veq0JorNblGm
iStEEcoF3BKPYwUZDn2iYoQ2v4alyKnWct1K18h24avAoUesyJs9b7H0INDzq00f
hdKB7ZbTpOekhQbxUM0NZMKy2BD4oYo7+UIvffEc6qm3fWTmi5kAZjyEC4ubCFvR
XqQ0B/Da9YEmlPSs+jhvr32+s/A+2lBJczfQAMvuprnnSfxBOlFs0U0S0dK5aeMv
IMuNRv+PnPAvADvQkMYhtz78Fn2J+79l5zI00YGyQQVOrMIMYOHvi53K9Hud8/pd
Sq/5CwtDp/4eslyZn0V5QI7YxcWRkJJkwPP/B1ilcOcr/atYvmM9UW6btZi5MIbE
dcE8OuLYNLi+VcENAZUQofBTMmIGHT7qkZOZTOIg4Ad0aTqg2er24jBo9/r9jQAB
/oJgDMF+iKDWlcxViKMyMB19n6/CSREvQOlSlW64zDlRou27qgM17r1e2EyVL53x
orGKJkI703Z9oNL+T3j286SOm7JMIlugE6LdMhsC0g3zfzLikP4LMyAfh31X+tgb
aXRhkiJ+Ro9StXMdfOCUolA3pb5MKKlPss4xOs84fuIjoRG8aCb4bqFYkrh+VxxI
Xl0tgqjli5vtT3fRAoRvju/Qx6meqLElEcwCG63k5pdv5jVo7b8NNezoEuGQkD5m
bOCQm1Rm96xlc5gb6ljKkRXqk4yEehx4MFqglO5Jx3FTvp98afRYYqaLrw/z0L7J
7luedQjFkHMzrBBlUVXycsprVYUs+eP9YtJIq2nYlwHgKPCigJx+y/WWZkC+U8qH
s5KsexpChqLr2wRMmAcJ2g8JnRIDrSV+QdeQyToKS2usd2qhHBMr6KA4l4LoHeAH
YecA+RIgZm+M7qhv5PnJWyeDIh0fK1T1YbjpUUlIBhv/z7hCZ0nbZTXCJmm9ej4y
7jKScZq6u2rXyisap1Ex2y6rRj7p50riPD2latb14zysrRc4wdQPtpHXHTg/Jz4A
loLTVCRpN0KcrcpFkCAlSmAsGzPDpKaGgIciu32sZ5LVHogmUqME3Ou1Bbvmxd1r
ovZpMUuiLjuCQOqQjIYN+dURs0OhOmNC2jeont52qsCdOCAZVz2+5HPN7aYdik1k
gTEpYWCW+DgT+kKKU2ObmxkVhYZ6IbyVP9O8XW8DQXHbB+opsAKx9icxYEdn0Al3
Kr7gBou7xlR2INEV4DzUrbr0NvBoZwMJoO9Z58Ba5smdeIHjDFvmJyv3XG4TnzsI
wX3PhDB7FAZsHBUKv4RL0aihJz1Cos8onWDZFjGjFuS4AZQ5IpIxXra3G0/NyXr8
CgNhUHRB2FjaKybKZjsyM0i737rlz9XOCxr2D7RwgGxFANhav/Kact9ifZGimePY
YFa5sN1zehfD3qMRaVZi2Cca/vz6IeQaBNuDYm+40m+DJpZ3o8qptis9vg/GrmgV
nE9DcqhQMroI6h97b1oaH21X9cPvUy/y3FG0t6/1HN7mHuBIz4mZD2xb3F4jMcoV
+1xsYCCl3Y0FCEJQmGG4MSx7Nc2P5DVEEybdrCfvW+YqFPSvPRQovp4viSWbtE+9
LQyRUyymPoKHEH4Jyw36anYRBePOr7OwU/TDbBitvwsq4zkn/vNvI7ES8pWVtnK/
FUSVXk4RozR7pAYJWnf/KtM1D/ojDehFyVjCyHt8jDqUCEIFlOvBx2Zlepp+Z3nl
yqHYoQlTWzoSS50w4vKVSuN0Lf3pz4QPDhbyryjWSKU=
`protect END_PROTECTED
