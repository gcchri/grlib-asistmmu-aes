`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WrM3HfuK09q8T4U3XqYwvEcjOebmMGHcPbxU0XPtYcTFInafJPjxf42l0etS+63+
5ipnjwoV59SOv3dsvMt1ORmG16v781AX96EPeLfxWfMydjOyPxzBDsPgAa9zKGxT
La8i6tCKwsS6V/jC1c0K7YabHwM4e2Ce9mdvm8p0vhwltNqa336pP3xwsjmvIwRW
sQgdIHy4Xcg3W7UPkXhQg4MAkNdjHMAGoVv1P+99qqVOp2CrNTAKkeLK4p2SS32N
T64a98PsMCZf5uRISeto9MQ0r3jzGk1TDO8tJ9kSxxprs+rTi7WixyCkdlfy7nBh
jtJgtvAWsct838qQ2Uup/bjbgX+n81X7V+ulYtjCet/lXqnYy+efDfEXkxY7PRAh
slOxNJ/A7I4O/le9fdBle5z/UrhVC3JsgtImtnReu/p7s2doFkHxFDfy5Ac0hd6U
zYRN3gk1Q7XenApHPf6nfBIqL6LhV+rLRymZXt27ofA=
`protect END_PROTECTED
