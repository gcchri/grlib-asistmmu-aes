`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xQOtXj+d0JzaynsEPD0bji29PV2rwotlNLelU5DRM3F2O9FVAfwUVcg+80nvcjBb
eNOZTgpeto7o3Paj4JsKjuS6bBFcqF4egcpVw97PwIYdqGTz1X10cWn7iaKSjOnk
b/8l8r32pBNDt3+pEMXdnd2Te+kgGT3nbsPr/PfS3YCe03lUdCJ/Pa7yBD0zRhvm
2bj+GyDtkiti3V3EV1eGTYNdxjGZmbyErRzu/CcqMrdDJSSMXdg+6xHKzPtluPp6
U6H3mk91ca91D/rGh4aZGjR1DWOuw2mhd6fnw8Vix/PIVrL7d1jdgg04vcu1CRAy
ff70DCjZk0ly8z/p9TmakErH7iSGHFhWxCZ9ZQTc/aM4O3fl96Dh/78bFHGAAxwz
mJ4wm7YkbuGd1ZKAr0H3hYXLAWlpI7tYwnXruJ6uOxv0wbzN7PNrGhsz8Dz2t5w/
jr90CYV7Y66g1BfyJgC3+KIGalMbvQvUF9VPRrez3m8jc0WsMHiqAKzNCCWgv/rH
kTB/po4JVCqJoa6ZeYfjIQ==
`protect END_PROTECTED
