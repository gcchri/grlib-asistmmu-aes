`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n5Few4Qd3OMf4fhU9lVDBXs8e31bQXgyBjb92CF9O6Vy9WWWt3RUMUO1JRPlZpmh
dk6Uybo57+//thzPH3je1lVAPwlebqq0IcB/bRLDxqjtbw8gr0jUgNM1XbwFaggE
iSZJYKmTn2J3RBiphNvl/j4fzhSHAkVsZFTS4NeHERHskai9gKpWl6myHC6ZlUxC
FJg2N0W5AihtvkAfEGnozhUDhXidg8HdLj+ElHFsLmwXkvHkbsyvdJqmH380GT+W
Uh0KfoGo2/uTG5cWM44zmQW+aE5ak/Ye/AWBtt6JER/T/1DB6M7kmogi0vFYKhgO
c/mn7/ypfF4DHYQWuzNHMtYA4HtXyvPoFD5eByDHrJcZ/vdgiY1IVYa6eLsmKQEY
3J07tO8ppzTLVqkzqluh7LKqeSm0W8D98o/wLl/BkgR1ZnBL2Aly2F84sG2FDdI5
2lI4TzfBiVeUBjzIjrn+GBX0qBaAQeRObwHUGrP9aKJU7H4RwAVvSwT7GOwjWJ5o
5OTFERkYpvVp6qHJmeferIkwOuI+eD64eMzHQAdVWU32D776Oqkcg9xqYUfU0HSv
3po7GgX1UMJ4aJZGNuq5rxpjy5TD/7PU+wHenqngTUwdpbfmMUN+FmlLAfqS8W+H
SPGpMhui3S5fO+nNZdluP9GmAqf0SvgQW5ZociPIKZJ6Ya7N8MsJokiKMbYX+fsI
b5ACtjRPEa1LXlxpypGLaLz1DuKrAljdT/HE3mpj3leqIrkJ/E39xSgXfVubskOd
/uG+mfmtvhmzgrpw68tPrw0KSGXft2yhG6iYL5k5RWGWpo5r0ELEgv3fX9WQ2Kv7
L4q3h21RTZw+MRK2lHOpo48BAVhzuVZffEu+Iz5WNkAh0vz3aDD9C2rYcg5i7z2w
lmOz9pQNkQl7BotMoj/yIVOYmH2x03Pppo+HWjgJ0M92DzyiGnkwg9JVn/Fss//N
pf+ehK4I3pP6EuP5w8p0nPbJ8ddx4QNw15FxK0J0wrxrDNGYKR5UKXOn7ET8NKdh
fYJVDVJZ4sgBGQuBE6tKodEkWyifM6KXUHxD+c1DwlI=
`protect END_PROTECTED
