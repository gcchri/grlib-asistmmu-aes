`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Pwb+n4gy4kHW5wCe+LevTNjYgA5OI42ZE3EZu572ti43zU1cxZQ8Vx6iKyGEL5d
uhOEuw0B/GkO9z5xjhLrrFkeEM/e6RpDjexOnH2vg/QUZXQrY3edeP7ojLWsTiOY
XFeB9mwGozNIrJXrPjkeOioaTMaNz6TyZrT5PVeBpT5LXohVli/T3lTN6HFYbeRe
JNBekGgv5xo/mDFcyjiREuYWENDfJwwbBfdGYwbBVO+Pv6MjrAVIEwZqxO+/jQhX
K65fVC8TrpTA9EjbtHbVXuCopEZPtiyC8aghYhUgT/pkeRnnkfcRasldwONmsSED
kX0qhnVepiu50DATRFIREwHsZfI4J4aQbCovOsWC6vqKDNRejN6E8zm44/c4E7eh
UDdC3mzlzfqNoSIxWbjHhQ==
`protect END_PROTECTED
