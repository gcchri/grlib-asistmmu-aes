`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9YB3HqJcDajWGwfIjaQCIaEPyZIk97sWob3bTrRWnAjB3APIYK9l+9ibegot2yFO
oy1te1lvh8Y2LSePc41thSJDoLnQK7KYWNkJsU7RrSatOufjFJeiysLu0fYd6/6+
oTvloPw3LqM/xE7ArjtneVvB7UMFBGmvIU/av7fsnkwXo6LJjIpEj9S6gQpSGXkF
gGgrHDjlP3zLZJQALz7CRR6fF6H/rdOwZaMPJ2ZF88x3lZLoj+QfTF8Wo1w10owG
K4nyUHdDN+OykEJOMN1h7wKTlDl8Ql77NemPTAJpEBsQl1FzTIEB2cQJ/0BR610k
OMa/hUyblV4Y6dkvyTiFjr1C9HVKYr0xSmSAveX2fbI5UlHuAxVP7AcygqeYOqlg
pyld6HprHfnzahFFGGm/tAri2HeKwZFLiVH9eci13UGxAg+d/JyKtFUxUs9NzfY/
zo/2PDvsejT0q/zeHuMijv4LwSrKKuWxu0SwxQyUbfBq8MtCqhfc4oWZ7HA21vj2
MVmWyj0ofXiKJkwJpbPQDm0yRfxzfVS44r/39WkTRM4uyOA2GowcIScmOMCABpms
b+m2N/iDjH7/RlmSI4Mqk1Qt6beDI3ujcSdovv1v+HTNZzDkFR4h96RcppWDyD3P
lZ9SnQ5aufzK8lED1mZEoUl8ilg+Fs65euZMHJTtb6aQIuw7SBdCkCg3L4wjkEbo
x0gXy5sWcpYT/BQ6AqXKx7todU4ORbKdXAh/0Y/HBMfQOxQicZmEnFlzbS+gfxjs
+0SjO97FF1z1/JqZzSqB3lWnyRk8ZsHiv5dU7RnapWkrzK10LdVa5qdhRiHh4zhV
hvbl2lIg3lvEhpOnKhqDHNIslea0U7Fa8bMcTMiN01xBSIt85OwkeRcnbgNSZJ95
MMGlE2N7OYahZkAJrtm0WkPlWPzI8n/9wVU3A7nQHB5OmwVC7WF67dbClKDqq2AC
vLVtVsMs0ZJr+fPuccAWX3HtPApZyApd+WbNzOr3nZlAQKpe7Vns4Z8rXeOgQNBS
9cMkFFi5hsKW6ZTDajsdFz9JLN/z6SURl+9zzC641NaVO1KG3g9YGw2HlhcNuIYc
eOgApFGywpHzwJVBG7C8g9e2tUMz8H+lOoZ6QJ78yG4NbP99l+ieaaR9cGbZIbq7
v9Dzub3q1INvwphBBTXI2RzDEv+6pLM0IXBsj9/APTRR7sINlrC7AR5diVsI9U8Q
Po5b6d4AqTqfQ5vyJOctFtPs76oiMvcXVLIA7qLhMzNbIxt3bClUD9xBkv9TWQGM
aa5fPLxqTFyxDE/UfvESBVrwZEMjqdsybRck0PXPYWVIJxoXHr/ihYPXeozw0RGH
8bNP0qbwJ+CbrHv8opR/N1W78nbdX2fWm9YUqvDc2XscAlp/sk9k/USph3tfpBig
HTXuHOzBnaHika8ozsSCZ6fWkdv2rvV5v64VkLyLyEuFHgc8XKamGLXqZqRH4OAQ
Z6RhMSTnFRDjQf2vjp3nf4iig/EPqUQs6oC9ReCWxVmv9I5JNfgqHrSY3ToVYcRr
rrLPNyIHkErpTJjQ5okaZ+bdyUIPFpeQAg+OfIDGGz3YlFna+pSrdQg9HcjYUnXE
8fkBzH1OC6FoBfp/fupYMmJnU9I0dXxkNs4KvoCacmOoSsBbMtEo5RHN+uG1UOzk
x/rCQTq55u84RFBG3xU1DZPLD2GpNaGuCLn+FvlvkaJuaKwZsI3UlF5sBxYweaY0
TGn9i5PAtAvqWeXFsFXhxuNKZ4sygZy8u1KpPI8Y1T+yrDpIgDxHEOQ8uxZ+5mXk
Y3gPNSM/+NC78JZAxvU02LLASEzT7TQWDM2P1EcpfE6Zwkf8DUHVnT6a/j4nLrO0
SS2zWRMd31K1GscDAMFw5T+y8mBSBpm0y/9rYpiPuVuBsd1iToBfEeJgxv7S2x+z
3aKnxVTmhHeT+IihRzLTzM4gfDifQyQshg4g3TPgYDBMzCM/GzBemGO0Ioh1RcY+
a2tOwqbuVrHm5JhH2bpCwPokWSlfPHL45Ekn53IqzXtaeOkC+yAvbAcpBaHjb8kQ
Pe9eWJfqUQezK+PgT91Vvzyb6tAi3pXCXGR1mxu2piYHkKZynfRRk5tUcSHTtXJ8
`protect END_PROTECTED
