`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FSXqlFyaKGOwGf0gOvb6qz2kZGgfd4srHv5Yjk/UcmUjrUEx5yU/ZqPDEQK50jjC
fUzn34NqT3qbAHf20dP3t3azRl0I1PjNbcdbNCKWOUfJ0xrrvR//OZ9Zifo05zX8
k24SE69FYxCYFqIBg0E5kuvzJ2AHM7NgrNS2M3rCWO+mDeIcilep9bgL8f1bb3Mb
i3L/3wvFt7abjjXJLn+Jmc2kI5mmKic69jFTw+uWCa++KLZNgh3vsNqBFqWaFkDx
0RuPK/B6HUkYBMkP6NMULmoRA9coHCda5kHsT/RMWaQmvB6wGrpAVSc7+wWCsRFE
K56olBlJSezw5vZf1YF7dgx4kqYV80NFixFN7rRd2Sv9W0rKXQOj1wPlw0i4Rcfa
gJWr1dhzI+482yhLix50a0id5puTLfEizctfCMa3zgMxjKHXmfgjRrY9hUj5GxEI
n+3zbCoY8raGgYdrH3i9zHccV+4PMYwO+aDyG739VAQ12QFe0K2DEnuuVRxy5BRr
`protect END_PROTECTED
