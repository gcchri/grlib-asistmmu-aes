`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b8AERKyoIaQAb0LkazN/Qh+tiFxU5oAyYE5iEG42TWK8wIeWwX0ck7wsxXF5HXmr
/Jr0E0+R+o1SlKjc7I7OEkb8yL+ocne/D6UvP01Pv0JvunYmCfKKDypvZNwFsjs/
KMGuvlKDz3E1ib8aBtm3YErSE/RVyk1szqSa3L5fnYINyGoB+VmNNFbW7swbuurf
zJU/MWNifTW8qV85WrHOImhLIRczNDDtgfCskIhiTbznelWZhqkKK3iBDojSu19Q
aCl+y/9LdAfL5VJCIysyPzHvsVXN8Sn7vsv8ffTFyyAJLlwTbwpe2wdiZcyErVRm
i52N+rO1r/ifLKv9zY2+/hN7+UG0VfZlVH15tp0zXZ7juv1n1uXtHXsIS94vFnYY
UqIcR49kie9DeGBZ2JFsmi/gvEfc0Q+wfkg3TM6kfiF4dQin6BKZ1NaJh4BDNXGx
uU/B4cVpZk4+1SNkl2Ymq4NHcxF7YoQmOU8CmqEbaS7drIePWfF8jnWnKRzjAVZ9
Afa6/xOLlCP/etMvfCshlSvZgX0PJ2Ul/TVRsNrP6NzpGq5goLTnZiqMaXEnJalR
6yPjfkrLJ4O1D5loY+K97V/zvsttp3A5c2wpj1nWt5KOOxq86T/6Rnb1OSjHxp1Y
V7BbE5Om5GBtbYvjSoxqzrB8u+auWLBOVfEwRnsK2R4rWcv4mpJFLQH9zTILXXp+
MgcOlDJp5nljvhI/nxjYXiQVhDkzeINFG4BXCYYpUV/xqVLFVtimt+iHQac7d/41
zmH1ayXhNoErFBta8loNng==
`protect END_PROTECTED
