`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oMyqZn3+ElZMO5/4rfMeBUd7Es6n0Gj2AYuh567/xYPffEEsuQ8jyImwZa34++HM
FykJAXGKLf8QT8s1BZUHHei/hrd9J6VDBoiQgXJQaOkeml9y+w1naXjPjCKv2DEK
p8umYVflgWErpllTrzmYA6UnstsuQ+fSwf5d2lz7TGrxrzphl1nKgdupMek2PaGM
H8iAPwAKvkob+vx/b/AFy1sy2ZyX3YCK8OjyH3j/4gcOjo466+W+8BTA3pXyNJKC
XBkQuUdIJlWdxHS5Pq9bfFyzn5ow0sZhhq70r7WiHA+DlBrf5hUm2fQMrG1+yucw
Xt54g24cAuf1npF6ZabawuNmfiopEvk6ekem/lF/jXKVL53nLrpWT1+1HCKZwRaI
djqX35uilpawe2QWQttokYwVbHcfDaFisBs/m57LNBnIcehtgLOKpnxV2WuhOJuW
V0q/HG6ApD3f3TObSGEFfCqkQnFva8ejjRm0Ae+tC9SLP/ZfotiNfs3/WwdVyZ+D
7SPZkWscRnjkyMiCN/u1IIo0w4LHyy0NosVAZ5EdaEMn9QHMROKQNjSEWMawRZY2
XhZakIuetAnGSKh6RtriaWPOtxDlL2V+ix8xD2xXKz2ig/mPnPe2ZUOEVfVTJ3r5
tFkuJmd4ZlffwPMwTwZnv6d9fOsCa92+Ts89/h6F4DQlDqGW9oF/rDLgv3Baksk8
r9GsBXXGL25xYKOJa8MNVYPVtjBUokVi2exTH5JNUZbjHj/I/tKnkqM/O0U4SrhY
6upYjqe95Wjim4rHXr1zA8hk4kr0LnuAO4QwaSGmELs2QzhLc+zh5AeYKqV62axE
CZLqSZ/iA+ZviL5MKwQnslJYJ7vsnJEN4lyN5kTUZMcN/1WIg0YzBG9QpZu3Yv0Y
2HBfZDtTCmxt7Xgy3TNzV49i3exxAilrzq2YK7l1VuqgdzxZ5/HTwukrTLZXgmpj
SpcUGflmw2QzzID38iYEoZFFn31RuXRvIWZLMPk9sPwEZOa0d7wRvuKMqZWCxlUx
QSvpism36oeEIMFte5GcmMcTmQFtiy1+76UfoI5XS95T0jF7HEQH1WgBrH68dHUT
Gi5y4XGurMaDUWBgkqwMkcMzMZM7uAgt1n3fHbg74AVgZqkBnZ8jCRDLXYm1Lpzc
MrVwGmPetH8S64Yx+B+dHYQSC3QX+Qc5wA4JZ1NK/tSP4UmB8ESCRLqQU7IVK8RW
yjA06UX1WXv5Bg7gCwoKU7ruULHrjuvgLt5Jnhcp8hDM2OKgO4ILfLamqb3gmrWI
2RFo7eHIo6gOvVrNXPglWy+4OltW3vrWMK4cjHYl3KsDPFsBQRNPxow4W+ZMuB32
DE3cyBK37ysJgFdeBvrUtgUtcn61+kPRLGoSfssFEgalpwkaSKOikiPqpoTvBSDR
q45ghy+Sruw4HFHd6gQgOCba2k1UMOc7m8RsrRh3WcXNJVFoB3BQ7xK1GRWZQZA0
0+Ni5Fo+SZXf3D8n61cJwT38nUtqTYTm5LSBUBkKo7JQgj9zpOJ0Bxu4MtMVgqRt
VYMc0nFVGo4qPJpH3CxukiqSNIYaWj+e3s00LQ+WnF66Rx1anFN42YBE3CcqA1zS
c2Yz2FnBPsj4L/OqfKMoECz3PNWavh+hmhkU/hlcOtxUkGhlCL66M9sd528vegmf
5LHeDYdR9V0csgn27Bef8Izpb+GveuOgcn3cELeFZ1vfI9FKXWajqXwOnMkq5XJX
yr1/4d9eN+eAsic/sO4fho08iQkhJqmVppunZHGfMndyqNChSvQVtFnGV2qRzXDj
3U8KOx/Ox4ZbsVmyYAgZ9/ZxXVUwbU+kMkLSzlp72G2DggpvgeuG25I6sSLdPnYf
J8yRQzs4zwnSUv54S0iQhQ9QHMWqIAeb+MWqf8B1T4f43ClkyAaEYrCKSeVWvzS1
g6XafP5ZyuvcyizIJNtyHhcqiSm6NzMY4PcxS3ixGF0B7Qw1mDu4XalsknVOAyrz
t3E1H35ZwEoGswUk17xEvdCM8JgQMtXUgL4bqXhi75EY3+lml5BBIbKUs6vPRwuh
tCCRXOPQBZJx3sN4ihaMx72ZRMVb1DYM2YdLtCaQ90JrTop+7Tdxq/yjSInjUJMh
96zzhDKnBRfRQyXRAP6+QNuvQ1NChcFgC+L/ktrb96azkeISlGtp5ryvMz7ryyjB
NREXminiMfBtVzoCUK4+4mbGrBudShg+7v0ZF/Xmcl/+YLcwKw/A3fCS+5epEr29
k3GUuQRsTkmDxFFuQmMoFTHNU945hy4a9mk8QSfK07xPgBmIafYIMgqgQJeUODje
49c5aF12di03J+fnNN/20oA+EgQwauUi0IlTvUbwLu4+MsDKKWg6Y1BiymT1YjtI
PRaZRFk2+eijfoP4b3eamVkM+I0SXNDj4pBKto+Yf/sUlzrpbGC7/kiejYz3n4o3
nkOEqr+WHLRydICBuP9bOCsqF8F0ecbk7yYjOdRTzGEbcduMffe27ryKnEFgvUQS
YojklCDrF48M1ZzGa1QVwDVNOrbO63yW0WH/5TE9qo54theoSPK01QVZsebf6z2B
0ZVFt3UrTvhMeLXkbs5MHBRLedGM3cmS/n67tVd72+kWwPIxwiHWltMc5aKc0cjn
bNDXVTX21Wz7UsC7bdY0GlW71OaaOvt/xStP/m2oXtKe3+oHK+D6d62GfWJCXC5w
7fbLFEnR/ksxb9nTnpLBvInU+8VO3Bq40opQ0eY0DkmHsmZ2NLmYW8/eBbPMDBGn
s/gHPxjYNq46GLI/FdkrFd4d883T+CSyz06iCsanG25fUiSjyxVpM/UPxqJIPnp1
GIWuSdPgdQpG1xYgOB8zIi+jIqspI7UJOhIFfghdUZNvRDzi6o8xGDtpY6JdSWIj
Lz3Xezh8E3G13t7aFg+0rEXEY/rz2wFDFCxh2ox4jYqjcAfWDcY63kVv6C0cYXp6
5u6XjjssAyPnLQl93xDph/jhZvHI8JWwVxFnDcWz6LbQGcJ1FA6Q5IluVfb6Mqxm
DWiJh6pGa0eCcMeQWY1OTn3O57CyKN70dkTlIALK0to5zJzPeLdO+EQftbAKzVfQ
RZd/1TZzitsrxoHHGHKZrW8K96mE18eM60+YG1JHR277mag0QeMu5bHAgkGOtOI0
yehjG6Px/72r/biwfqdETJrCAC/UFhK9QPh6yd2D68Ik5XVaUcZ5+kAIsA0SjCu7
Gnn8B6EMcKHc/GiMBicbQiQ7+Ivrhq1xBOLwilIl+Ztmq2IcGCe5XWsL6P6bPzrE
3mDW6aj55EhIt0hDXHM93RNSNpNBOGnLg3XsyrvSrF42MVxG+UAJ5hHATBep4NxR
wz8fqSvGqw/CC1GA7gYoCUwfry7vYgb+3SIO3Pdj2nCUrKjpUibr4aw4C4GY4YcR
ztW2x0l0jWxbX0NCJLu2ZqYfQu6JUCdyE09X/N79kfDjneNXBNz/vCVhJd5wA2nY
zwtfXyslyn2aEMivunsh/iASZERCnb0S9lbjfvRviH/qnKolyrMyWR36IKL99EtC
MNcdTdIiHrIl4RRMlt0ciS9bJst2ng4+woyzk92lvbjnsnXEKvXCZ/GcL5lggrOW
bMkU5Kv4JCW4tWTY1UkTxSSALWHQecr03gEjJBuYqN6dHUIdFJo6mnWbfWn+TSoC
xG+W2S78oALyxW6apXWQ2946Wag8+AjFk7QYHS7yKH6i5NE2f0rHP2PIys7VLb49
LSkAqRjCRWv4ljVgKRoDEfxGFrKLvSltC/7VdXGbdMWpCtNwT+h1pk+1byu7nJOY
V0cW4hSyua+NsCbNI89NPZl7rFIT2J0xn1mj0sUFz0tQJ4JCvxefpWW3z7XV/92q
Nfthd/E2f8DLh9o7GKNPRzwlMSng5HVoQkI2eHIgc/ud8Ghm+PpE0idTtE9ZLbT/
zlZJPA0lRKKNLWrRPpFwTISfRFWSD9EFSoNOTxD0H+LUOzwPFBODbqfuxRCCJXp7
8mCuaD3aDJ4N1xmAMf+1Pje/TQQxll2m4EMLlKMEBFIGvjvYN2x1Fj2E358N/meY
7+nhQfbs6ulXeuy51PdeklVaC2/WY+8w3u70SnVDbe1S1Zm7bqzxxqnG0ezt86u8
ye1/inWAr4EfNJsVWsciOvEEn7+biMUp3OyRMyyuyLTtfBRLfrT5NQrZbA4+euHL
Et4mtkXbTLpg2vf7FdFngjiFSHCXPiLopjGu8sQqMRuNLc580LYGh/iqCYG+diKv
Gc5eexRjHSPripr7BhP46YP879XfZK6KsE45ozUzzE09sosBR09G9Uqufq8PBFNY
641wyQYtalRrtDAY4Mjy+0m2V3y0nlB4rtP/rFKkomvkbAU0jzdqM8McZdSdDJE4
ObCZsSaC+TXNU5CRuXgLAI2IZTFjoVLeRl4Y8J0971lO78K0+LQtSgutYuxyqaZa
2J/EfkZ2pFRascfWbPkWSYgugth8BGCyl7cmra6O/QM+pjp9sQsJWPAd1+bQ2cfH
ykouIcWUTsRKhkFF2O9EC3hjFX+vpIAZJkkwC8ri4becyHlLB+38DBfTgXbDu7jY
hrvZYyt7XD7PyoRXPCr1VrzrcrcysDemZF9GNiOSEvl4O97pwPpqRTljN/39xeEO
0x7hRmt1nidEzACggtxMIHiFjx8agMLAdnESXBtbNqR8vXppi83GOEnGLXpQWs/k
geu/MQg5xyluf7jcfIf4JSbPz9NyHjD/cSTzg1RUHuhyPzU6ZiR5S1swP3sF3zaO
sswFKhV6LS7xMJdgFKuGmmtEUx8GIhELlibhe6XSyqCr25XZDFCGiwWP8Ap5YwL/
DhdblxOCRm7KvPNtcCnuJTr/L9E02U1GSfIG9D6q9fPXOC+ZQrCiKhKjSiwi4on2
SEESZ1UKWfczhHj2WCnXbd7yThcUYAw+Zaq2y+YSLs6vzEeHIgwsQFGVHg3Mi1/N
zX5zzXmB2BORiaQ54xrRPvKOTjTWzqDW9n8v/rPvpmCZ8pvZFuxPq3fUgaI9mMSS
OaqtdMBCY4jfNc+RzQn4t8ezo+nQicnXcK0vatxyPsczPSXyFCSfL6kzyq+AkIl4
moALre34y7TsfUSo3MNOuZz8CniA12Zr53xICqQasgeUawzCtG1EAFJFT3f7U0fa
vYxqM7dkQRMcmE2kXy3al0Gi4d7HFTkSngLhtsmy1EYsKKoMnlraZ7FkHHrI6yGn
x+/qh6FLSx2B6EqpFPOTshLBlzzfGEKoocS8p3YceX9EtCHh/K16d6gJSZUUGcQf
YkiXcCDvaaswGJbaHqZeBhZNzubj31Bn5o69/FlkyV7Np5lKS9FnKZBzkEUxh3FI
JiXMIwkVdFUKQEKpYIYN/aqF+RL/VbHNsR5447PuRutRq4s6JReRzWWS2E83mSg0
roYV3f6Jht/PliaFpKWTU+VLvFqJCvlPJCgcQoOPLg/gcY0aDzRiM0fLeZ9j1K+G
2vRpB5QmFDylhB4zqu/dSmkZy4chIVCRTTAjmM2IJBAu17SF+snqJBLHmKO0qo8Q
C2UEYGOXTqv1rVoR08dyfSMDXuZgP11gIeM9QLguPuK/nsR7CyAglpemYBbHmTw3
m9xsJRJH0Q5oQWXWNvCJfbC9PaW5Ju4e8G3U4pHfcb5QExOb1Dm9D1a4tZbHb0zp
4mwhsTjwVfHXNDyyddldjzhl3SF8Yj7QNQq7iM0gQrLT//Av7KbK6ALA+B2hlcLD
fl60aXqhFy/olcMThZhb1O7+vZ7CuH5hcJy+ZoYMNiWyUZd2ooKl5Of4zUYuz0ZT
qD7532qYbtCHJVc/ecXk5VM9JheoXjR09AcXEqa8dXH2/fJchqokeAnZjufgowa2
sqqW3wOTBIU3c/uWpVm6zuSX29oY+jPcMlFiZEb3PLhgW/Sp0CjKGzjnrGS6jixU
CpiFK9PC4ky6y/PNOTKk0rVYyBu+w43nYcxfGNJjmig5NY9I9P8BQhzthYDox8gp
S4cfRRzIUS+p7UKcLXwwY1J50SpKDdCUPEFYMsBZAllMq1y20qkRdt0FZBs0WL89
/DooPZWWdaw8ZRy0Rp76YTmJIzIMvJobNVpxwfM9Dv88iAdfmljJWQp55dE6iTFW
xto6lD+TFEXXERWmmapsO2Z92VfBRTPXaORFbrPnIQ7Whqlj9ueOLKT8Ze6E2ElK
93JSSOYmH15XK6QVqUQaDI+vHc72awwRmCGpPaghtoGrUOfcoXphSY9dRmN6G7zs
GbGvXNPj5dURHCPKGidD9YOQQq1/vL+1m+9qiKVGSt1FA/FtHRvO/YTXloNTCQzk
YvoMNY/bAUFfm9Byzx8yD/YVtwJgTXFgezzen03DXonZE/ZjM/BxRZt3dDCDOUxj
i7Ehf3MOP+eSmIavtkHKcECR35bYmnzLs/xkqiHSqsGkl/LDUeVz2zufgEjWwsuk
wks7pHn3nhDywY/RVqrpbFdpBvZ8imXV8mHA73NEjlp2rUU8IYG9/6Ktq9sweDm7
FTld7Voyz4KBPRGBZOBIsptuk94yt7BXp5wYBZkwCEUsVA+fAK7CHkXNLp3dJ3S3
vHBNeQsIPN8EsH97r2/0o7Yabu26OsX7Xe+Guw5jTJdNsj0SZ2UMZtz04QpZvjDI
oZOt/bsRhtswbYWeqPWyu6iObdrm1LdGV6iAgy6uzLm/wLrfcTdmH4OzLQKjAfMi
vjSIOfd4Vk6jKXo1hnL1wmZGMz9W+TP5o+JPYZBgH7NIWofAW4h14pgGkbxZN1ok
FPwOh7bYligHQg+Lo1QD/UiKIuGLMrmG0v9sNl7rebxdp1kJc7IKOKA0pslke+Qt
WX+ZIeQIo8k8lN7fq+2JEGJ7AS+BxsFf/nXJ3K/i+VS8KGYLHgkbSQhY5R3u0y+/
RWKNms/VSFQlmrG5nFcFRA0tb7RaCgawnoMKKrtTIF80WJpINQxluJp7RPlwQ746
t8zGAqZXFRluk87Q+en6f3ZX5OTL/YPmRnRJw1wjphyG3Q7soAMAPvvZKAu2JD/A
hKDB1z46CXpA625EEq2YFLDlQnM5H86N+fmRKVdjdrhVH6sa/3HQix0iKqSxpl2a
z16UGoTz+ET+VwAFUaHc+iARlCK1+cLkldXDvb7C+7/AA78EKft0XV0tcC8Wnp3g
iMIsbgXtowuQBjFi72qoCMtTQjXi9Dln18qlL/uU3C3AM4zCoj6FnRRBpsj2n1TV
L+rabz01QinEPCUpEXFvBE9Kqes05XV8fMKJZvaLfRGdfVH2q9GH5nWJvkfgD+/y
uRlS78O3NEUmDRCw7o/HodI3JaIqbqqu/zueG0/EQlnnXmLicVvlkDHcfCH3+SPg
BomiQgTWWQlUuUma12gpt3teAbfdVF8204E3OFQ5fGB1OtK1xRYsS/BwL88sb1xr
zk2jslquVnUh5+eejrai9Up2C6kf6u9vr/D7bvpmNfvnt+3UEUwPHFvCLMHzRWMB
zZT64yLF5u/BQE2ioSJVAmE4Aq0ka58bJdQk0u0anIR27JwnIUXy/bpZvTnVzOn1
JjWhiD4vB0s3A3FERBN9xbNN3d22xKcAbU5kLxwFUpSTxVLsYNKAqpUtm0p3cqdh
av5cbT57mZVgP9X0k5dh7ioWubqZ1NdpnlpvYZ4wVdIiy48Tq6OFiBJMOb8kWJdL
re/y6U1LEQdsY7k7ti2A3tYP+k5rKlDKgkueX3ViUMRwePQmg2WB7XyxL1no1C0j
sIZtWSPWmLsm9n66zcCfG1zw3RmGtn1mhqcyUTjsykUEKTV3AfXcDqISu8ytOqwj
sDgcq9AyncvNJvCZzzRGAZHXEuagNX+ad+E5qRbiEi3SMBAWKH39e1t3IOujrhHK
3EM7oW77qxyEp9R/AK7IIOr1aFUSn09jMOjN/zOPJd6ouK6FccSxXpbi3RxcDKuO
CpEdwW2wQk67nZB1nRrl9XwqQzQ/AZnfKVDtLWqJ96BVldcdYfar2uKgAXAbRTcv
3vXYRlILprvJ+MtR1muPgR+b42osDJYFoetw1TgR+MLe9s0woHkdxtudKpxntD/B
ZNotyfPAKMmKNyUVQ5GV3aiviqyf4xL/HziaKEul51vJY8mysqkTMQtercBIQbI5
kdOCvPox/4r3MNmhG/ReRlh1jvAZ/JJ4O7FjS7ZnK84vG5qHbg9zCNHyb4VArBWO
HFosvRdo3clfxgT5wm2TaTUfNPhmAhvCG2S5DJo5c6tM2BE/DXvqOwZuS4q/jYBj
bhTK5ZkBFllAi1a3rv2Ql6MQYkvRxty2mS2alH91Rvd/S5w02X1OIHrxD+rZL4mK
8fYmE7ALaBPpWYmH20yAc/52AsaIecoXVkpQJSTUOLCAwOuxZQn4XDUtQLtMHxXV
p5X2QsOQrJ//QgoZl+DDTgapIYkzZaNZVCjwDQK8jrFCN9OrlR/i8vOsEasLJI+l
cdyC9TmBB10hrnQD8xV1IIdqQNCx6udaXKz5C+w3v+V/sO8BdG8lzdyqgcoKqq0H
xHXuogARUmdKI8aOx/1omVG04tTedGYDjZ+BdhCIuj2EINB66vZ//9Xj0pkkaXZI
Qis7PLSVxdbMiYLUkS9RUch1s/Lhn5WaG/7k7dEt6fr4u66nNWu7EHJu+D8qWMVL
dFSNmgJTdYz19YC8cSM6ulhEBrV/N6PBrXQkqUsGPEQt9PvFBF5yOlkydfKoDK3C
aGvAGhra+vGTLKAo0VSohctbNoFZP+It9FNeWyTjUL10vvPhpierRBV7J6FUD3xI
bD4Nx1BC7yXdm92J/XH9be9dwwhOR0OvBmGyxr0Y29OWbzIakwvc300Dk+hvW8LM
kDGZ48RVxdhS69yEj0c1BV3knG8LT0RkR0CW4GO6kSyPOfA9eH6NtAGhxLkhr99/
47gZEvFYvHPCxbBejtcvopK5ygwBTH3ejllzQV6OZxcMVta2qz8CD5E9X0U7WhwO
9DPu3N7o69ttQf45x1gNRe6g1+xmrEZRAsCfQIIqVxNBCN9giBCauRxgrgB5UBDB
GabAlvQL5KrtdM6imqpKmo/QHM8wMQ7TpcdqDGhZRyhPdkFXZSMGiOwEZJcM9kUY
oFIyEn/0zmv/ljMMp5P0AMafcX+gX0/meb3ajGY4XCLPSheGxVv35oK7SmLJ+Zwy
LgYRDTLbDt82zrNQA6WUZbtQ9lnAg8n59BujwNDGNgS/KTRmldo13gsQJVdKtiqj
SGx7jD/TlohkaME1VA4LzHgnN29WlREElPPcww2DvA4JuLJP6uOvftXWgYXCjdeS
LzO/aVe+L9omf6c2kaOxgmpt7/9Y47crE5gP3Qe/AZG/4lD7nNjzdcuK2cJfB7t7
TR1bm2+pJl8v/nCRn1YSPEma0+uTtmSROJlKSe1KMkSu1uLcNaAeEXldzEN0XC+0
v37V727aKsq8DksCbH1EggPTgBDfV6KUGvfnHFZl/NRQ/gtfklSKYCZr11pKdgEd
R5STJ9aEREY+tdfjdwM95zo50wMoXNqzHDofq5YXkWkJB2YS6G08hS0xsqNUMrsl
5avVqVSotqtX4/T0+BWBIS3TzSBHmJJbYe0bMPT/i17Wnz5moRa+8eflP4j1g1QH
5+var0+G3vjS6AGGwn27a3O/LkNlt1QMNMw2Bq5EQQx5Ul5Yp9l0mu7xN/4/qzUK
Y+u2YnyGp0kvdMJvDspFlwqKqSBPvV+TDZdRA0qIMVrbs83GsGd39kllJBBMZ5G2
0xKAfpF+OVJ4zHTu5SnWGSHYznW7Cen+vtpjXSqS6Li3LMPvG8DIdLQWGnhr07p3
g5Z5JIajRO4LNgNcdx/l4AhuLez8QjtJ5uhnp6XQc2JMt0tjEG7rPR4r5yTMqo8W
8VfygZy/V5+1lLP8mphg/g==
`protect END_PROTECTED
