`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dyu7ART6Joac/CJ6/39VDq9oRfJPDTMafwx54bUTAhEnXrxBSzX575Hy7AMiy0Aw
qrYWrs9dD07XU3cpzH2OwDagS+YYkod5IsGX98Zvqw8b4L9B628k0kRlLho6nYuI
S3gMjDmqRr95IRcZxdaRiLeZ6VekSbxW/e+kuwb/DzOsyP8t8OXhWp7G65Wfy3Du
KYWv9AwpHEmMfLADTv7tcbVmtwzyUZIb0ul8R3/5XMYOpBIEEnMJCIVGLLr1oGvF
zCYj7CPLbniT0BTlPjNuROUrNO+ertRtCSg0/aV2Xc6Mm6dgNxQEpnjkW7ifM32b
lOnCozJDhkiC4xakMKrxGyB702EOL3roU9QzRpGCn9Z9iCkDs7nreLsiYRPO/Fhl
Cs6udVEUXgotK5lkt4bgFDDvmjuH5JspXVPXZkYtxwcQ/4L6g64IxyLKJIpZHidX
NUuC9hgK1m/MSvsR7AXveXAFeBgR3wziart47aQ2MD9fEMGW0WEHbOPvjiwmTpAr
vNt+AbesI/WyrCodEdFfm00ZeVDvUUMzAaSJfV3SIhVX5H96awIKgL33zK2aImkw
rokr1kQskWAk0mPOMe/LYC82rkfZSGR4aXFZle/2zkZKsPs/xmHCz2lYj0/grwF+
IK4U+TYqPDCizgeE1Qqml73tKvAzf9ZfKlpzZ8eBSswjyu4VUe0dedslE6SPQQS8
DdN/LboCwTsviqLobGyXUDyw3tpTTT4PIKYVA7ZR7HhG02qfvYK8vSpdQxPNDFiy
8ptTaNo58nJfOSmjoqrK1yjm/NtYb/1cjAreSI4MCLdEy+JTk9tWluaqNMqyFc39
4xc+BuNAmzqKrpnk2RPMQGWjn2fcIRlt+aDJx61ama6Ezsk1inevjcWhS9c0dwTR
+LGPK8IYhhWdCgYaZT6AqfWTOW8m2Abz6POk4vCIaRm3L9XoKvYEeCuiJQ2wnqIj
7+3wle8hWLWqfwMvxJTltEzC0HFuo+bN1SJC5oFCFO2YTmy1vLPEo/r9c9lSASMR
F8FYtLeqD7/zItnJkwSbUF1ke7SBQW+5kuadIK4cMZjuqkQBqKMOwCFl0xl7l8pL
WYMPB9chWOOWpJFJk3pBvipcZM//YLk5V+CqqyRQVD8qc5pE5Oo/BOfJHoFreQ21
K4zZGlBpTTDWSLPqlvZsPSpj7x8aneNysphjDl3+PFywCulJJX3jFpQ90BdHLA1w
u1z+UesbSq6kDYoU55ytc+U+jCng0QembTwpK21CCADNTxFCuTFhis0nscmo0kvG
5U10Cyko0PG2bMbbkJF8iUNFWD0XVX1wVm63kpXuqIBXhDyZ2BYU9BKkcIEVxJCt
YkLQv2LD8QtY/zzzrb2enM6zWnoSudO7s5p5tIU1LDhcpUAauuKkyz7JGXFJG3So
I1dglmaVqO7XMQr/9Ozl2VvuCi42aWudkt1ONgHETIUq+vLgjY06S3XoMWRZrV4x
iHoT/AZHMfm1Z+BLbu4vhDGiSByrZNzucNeb5j0e4pJQ22TPj/uzDktPCNCyVB4/
1OeLi+mkwC80kFSjP+pLXzrbKQwz9duiXFcOjQE+0qIDetGIirW+VU4tneA1QngN
5G2DeN9yKJKyJiFsipJ54qkjAq/ee05qRYSH82+G7CByhiNoi6cidh2qLdyyXME5
wADKeQnt03/+zGMIbp9ijfErUxhQ3e0UH/cmpbtMoInSjYwuWrSXiZ3ab2nhAz3v
Lohu1VHhvR+8NyioQIVNKhvCwOUqk6aVK0y9+PoA0x46Q8tlA6ujJbZanigUVixP
lE1P8twRMe54DbPXfrP+DajlyOpYW24TSoCu81Z1F6/ofhetoN817XpvLdiHulTr
OIwJ620+bCcxWAZg4ic+tEQAX5En6Dfy/Y4R1vy9W5BG8Hsxasg0hmi1KN+1WT7C
M790OeVORFURALD4rX6hAj2oe9wuSCaiYQ5CxqJ330pqZSWdG6PJzdbsBX0Z82dK
pUf5yYqI7KJTsllmlfr22AubPv2707sSJSQJftKeI4gr9RJZyGfAO5zCwa03DTw5
llmv5GsMligiQLw891j1rHA0d3emaJp0WCTIWdRwtGQ3AEuxgW+2V884vv+O6YNo
v0qEolldjoRrBiDKf4suQs4SPs7kMsWOefgY3hnSQPifeVga6hxJscQ/Zwx7HQxn
V/ebIEqbjLmnDrSqcc/OcIsKZJeO85icMiBv/jWr9s+h/G1aaUGRh0PVMILhAW+8
5PNxlQqvguFPozqT0p7Ac02uHiAbvlDnkmAsQVN4Jn8ddYKkDSAzfpHVbN+zSZ28
k4dOHOVK16FZzJ6QDHjvzdP1gBU/QkAO5wf2wFtsaRg+I5qzdxxq7H9eBuU7UeNO
0gL7TA4kf8qu+dCxdP77b8J24563y5pwmpSlhCOYkCyvKBx5qOnDLsecK2fiYOjB
n3SLYPE+zFKwI7sETYdgnQoAVwoWck101xfr/tL1vx45g+vud+Js/Ld/o5lObOxE
kbiTkr0Xg0c7IR8XeE5x7m1k6boS6CK2lAHmtvCg2gNwl9IjqeqlY8vkk0/RBrOm
3Awu5CaMcHnyTnI3Myjf58gyi8Q/2N+I7FtO/hg0SKiyiQWiUC27KXItksDqhdBI
//DGs9NQYqZC5APPf8ARqsJkiQXJsSiKKyA1oKY1nrJhbH4jMIWa7P9D1ch5ek01
bvp7P20YDUNxpR4eEgmpQhnRmnPVaWAzZgeg//icKQ+fNZD3SYOob5DgAsmXkbHs
YWCuFn5ccAaGvPRlDy0etfdzOf897IaqdE4vdAy14XStfmfY9YtNfIBylLzzWTHU
RAFbqF9w7Om9iTx39DH1THyWdQx62lInxW/C72PEqmuK4XMbNmw2mCnKg85XlTyZ
ePkVxQdOc8dyNXUiYOKJ//gk8ldN/Qa5F91uSTTWCTmG9ZY44ZFO12D2tOotOCIz
u9ptgCbfAst0KtjVAghFvtyjnaWkYabR6yI5j4niQBKCT57xD1mrXJNs7TzMlN5G
BgFnVlQSApbkFagSYVLPZvJ1zSElPINOuDV/JDmkLBDM1Sop6S/0j9I7xsLa7zIx
EdLbsev3wBKYh1Jlg3385Q==
`protect END_PROTECTED
