`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EKLDn9w3x1RVi7EZptZ9HJo3uD3ZzpPIqPPKE9WGE998/jbonH12ZfmD1gaGrkE1
fGST7sAUi+E9fX3AcnsOmEG2NuLI3t1IyWgQLR8K0rbOYn98NuzZ29Ie1fgiybeW
Lhr46kMCftk5imo+0IIiqp+3kpOSoleVTXjcj2fH+p6VG1o6S18QiUrPfMo1AH/0
d+kg8tDUFHtfWVInL+rtuTYcMAHkd9HEKkea8mIo54vM8ULbXjAqpZ1ZnotRSH9q
fDljokKzaDV/t8vGJsD97/Ji9ggJNWlr7183v4XV5+SocCgtaXCAOWtDqmLEcF3x
G14Ug7mc2YbSql4wU53RdP9Q9R832nikdKHrBiTDBZPBwxK1vJxAEpkTqmEiu1dr
wya6MyfnfVaORbjC1+xgfMSb91ZjQDry7P0J3KHQqiign3gs0qSs7vMPbeEyCjh6
wR1Y6Ct6tO4TKBrPKa+GRR/n/7glHIAocCZP9c0Jb8NiH1f4X3qRa261sHb0rUy9
3ZwXedR4BQa2+sUJ8EDwda7DJl26Krc4lAEiVD6i3GDGZDZgFVaC4muDODBlNuwy
EN2Ou45+711OK3LlDw0/l5Gq9bHBxrk9KagN2nfwPjk=
`protect END_PROTECTED
