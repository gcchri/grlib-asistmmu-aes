`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2aZg/m7fTG4DXcK+4SgYBFAlzYBPZ8cjb8zInmcH3CE1vsRt9MUXrcLL7cNjIqF0
7bY9xIWlI+TWte5K/N8i8ZnbycS2Uu32zTQv0zJMyF3Yq4OdjAXCaEnK5roOGFTu
PZyLl3QlzLnkWMtEHKucRZ97xqt7Hz8kxEXJbHDwIWivQwmOpfQfeCyJ1y5cwy9k
IUxLEF6KYIgDO6hTiFqqu3lVzQNejc72NTJ0WXeJ2hMMN4cKa7izJFu5wPAsPVP5
VrtZyTdHma8q2hkJiXYiwkdVVRM44nU8yj6U+l45KvYDA/+792mDsbyLDu3oQAsZ
dt4QQ4FyxhQRNfhD3Cojr51+H0oCAG6ftBiQRY7b3E66NeX3052lkVxRqJBr4lfm
w6lE+rL/9JnFft2i9fEXtJUyVcOa9WdozitupVmueDSIYCy71xAzQYTPeYox4P0E
4uaLRBjSRVAMqPTZly2qJZOKvpN9ucWYace752hCg2HaaMjYOz71crGhiz3Nk1iU
CN3BdoSdul1XA1ITOpBV8Pwv3wEMK7sHc7jc/jkn5r8WchTPBa0rVJ/PnLlfBjfh
kN8vjIU2ljBrEzhWMewJ46Rm+Gr4bAJNwVG+fRT7QwXyLU4I/vXAZ6vG4uUHe3wO
QueMf+Db/e3deWNyo0GtI9olf90uBKBfk2IA+zg+fYY12mFy8Iz1ZsGTfH0kJ09A
zVlfREkRh9eavMPgjHfE+n3M9Le5KZL2Xq1tOoYqDzfD8Lda88Su36/SuKpbsUGd
F/CJmyu0dN9Xbxjs6nmeCiokVwOfn+sOGOjvvC1i6W6VfZihiyicZZufzG3znUrZ
w0Y8XqQocCK4ohwUdu2JqYROfejBSt/1G5UEiInD6HMDvLNr27ofNH9Kz4HNYs2q
8hGXdvfh8NrB5E3hXG7/WBBZpeLPj2AsbxB9pheVvT7qn3jAZONEAv2SS54FeIkK
RZWctYtp8TygMxBBO+AjP5n7HZfZQ3R1agV0q6tSbLLBjYXw1TqXjryZlLk1L4i4
NwTXee5fGeJqefZRwYrsH/fwYzdi3VEjXqZfCpY08UlVQSHgSdIiWIT3bXZtk+XE
HjFb2jizp2co+qJ+a6XCEXE4CoEfKIL+k4AARW7fM13s7yFoZ2uOVtsk7ttNuYG1
2e0EZDiIZ119QVAr1nHbiypp8ZzjYRMlIf5LYWiO6D7AyBvClI/++eWXdxONU5T+
BCiPzPP8Z6yO5/9qTBC6MNmZKvqR72cSfEtBB05FRdz5mGscwPai8JoAB5N0c0pW
ecjgBvlrY9lbzDSTUAhYpuk3gTEz1xaaAKqde8r8iHKk/ILjr3z+zpj+MgL33tx7
Yi9fG+2PbZQvZ7VjYoOQNS42vZ85iaWLYFJt0eViI76WacqPHI0VhAJwrXKIGyh6
PNJVh8RSi4i+8/FInnr6RLY+yBNWQr01auzCC5GS5vTnoQnoopewBdE8KV2ZHiqq
Plf6tLKh/CPeG4HTtvJ331aX9nun4kf9sbVkdDSCJnNNCdXf3n6qPqGbQWGPHg7v
d682jtyymdgJ25HG6E10cTdcW3Mk3jdLqet5zjgviDGgOPSy3EIbNs/smCmgLrZH
iOwLVkiuZ8ly7sKfK/R0ffCo8DUrqa2GqsELRaRs0CBQd6K0aD5NHD4PYbaeUAYz
4EPeJKdgM9advJQQpaniNp78Fz7QpQ+NUDApYH34XV57cIIr6oXy8RveeGf0G2QO
lf9sziFapDScAuXKA8bCGHI35eZitOgSVtEdlD9dz0+rXDwPR98t7pNpzvYsSmYe
9dDZupdUzo5C4DBZc1QWkNj2q53I8qUl/zWWp/h7f2D6TCf6uH6y7rAuucY/jVwm
a4FymZJvmrVbvVyTYwxFKj9jyPIfYnbyY3fHPOItOsygOubPMM264SvjA9hBP83I
Pp4O/jU3lMfJxrWrmDUePNwK7WcBXstA8uoCbGJhrKT8sh7lHhYP7ZbNSFvevV5C
nY7LlC+jdhKnDevwkggGGDddEjhJIw9ir5Siy9f6QBi2XHh/2APxZvuwSQgQ/qLK
Wqf5KOQxlWCV2BNoDmRE8+E5oT0PuUU/QTwMQOQQ0EwBTBhv5IYa7sduPpqf/1aL
QvTwU4m84Vp+Xpn9VdpaxwBJfiXy0NW7Uyxlb08Hb2RTmspzYB8ma9+biOjsgIru
At7fkYNbsuBGcnqS0jYWadt7sTeLybXOd9DE4VjssMr3+ZMgQZQEIYqw4g3r6WlD
qbQh9nIHX4cgjRYs2O0qEEncI73HhhSGMjR93XxXzFedxkc4qqLHxFgI3yifmYM6
KiqpNN+oBM7w4jhA9ebAg2FVdCQFx+bO+5SzVCaBM/ZaJ9Y42PUySQV/lskT7Rlx
XAH3EFg8W9jUsMbSBChk9qRcwZPEqC23v97cdjJvLQEN4GRZykKa6hKtSoHANF8v
U5X4S/tfjxtp4g+cbYTMVg==
`protect END_PROTECTED
