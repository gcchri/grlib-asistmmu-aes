`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bwr2nHtR+zn4k8BEp/gE69ANUXChFW9lBMNklRPZf3fAqD8IMl6xy6uPZtLZ/+ak
5TYwuwRnhpf3LuiYra4CbHl864IpcHq+brTtVn7eq8NN4tDPkz26DrlBseZB+imY
/Mo2O4uE0t3Rz+QGjXiN5p2NGXWXF0vMY+e02BTnueTyVmag2xFHzsrgRERUh0hE
4pkqoIfqvGcKgCzRTb4/DHHySLr1EiipRlVhpFMUHHC0InJV0jhdgaMmUYIIEKUw
xs8TcfKOOiBzo5UTQJpwEg==
`protect END_PROTECTED
