`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kXXR22v97gg62M7uomfT1w/D+tGK4zArN18dMBV8xkc0jEtrzt0JMgbSrJF8tatl
gJQry5dPTVuHl9Mphk4vvCCWYBYC08wapMmpDwbFVtDt+OQphNpDMzhy7LgkvWMX
5rxOzuJXrUYj0wH7y3u3L/hw5cdKmwvgBgzIzFaRyd2zSdt5c3gL2dhrfJziUQVx
hcj1k/7RDWcp8PvYIatIor4ohvf9Ke9kwZhxt5IGAHoZAgi/gyHNq6nm6VwiAYoz
QAfW9gyZ6fZhAzA3i++PIBWvYPGNTjxvktv4AXeGwulN5niipswNLBfvK6/vD9sW
mUcNXuCcYPVjUVTB2GQhnMRDznqeVZzTiP4XLmQcGw1kMMR4ZF7BKfAboXVRgfYN
o0KJHHB5H2mwa1tNx2PQbveLNdnv3aXfm6/FAMFaZIW6K6H3LHX+BUeCZ3tSf4Wj
5mQx0RmVu7iVHM1v62Uu0iu9TQ8lH0Em8yZnH+Z68m+CgtiX675Y+/ra1ckJgirP
VDc4pD7qKVjtJl1cNG130IxZWepp9Zej0v7HzclleIx5moAvUJzGWqPdtYg+m1Yb
UBF8X7zwbPuArhUAHXHxnQ2Q/7xq9mhLeyG3UnSlS/g35cp4qJVk1t4OvAxllwUE
se1dnKgvbfefNKy8aIICZwSIz6EmB/VjMdASDxCOIDLIrDEeUPBvRwEotLvJZWhN
8U9tSdVTr0PCe5hz0ZBeiPprfU/HeC4SZ+ieuYObXq7lvLLSEhammrpNu/SLBtHk
133qaKJ4KHMwgwxBA6ftxzranUTzWkOozjZx+8WBSd27TwhAeckvaooiQnPc4FPd
bnHxn2oI67jvw2XmjiZe6rWWq7cjUgwzpRvlr0uAPdThyKtnoeWjkD2PQQ4fqPqR
GWBnYmI1f+v7dgb6V/picEm97LTN7IlNoH/Bera6qkdwMN8ShpsZ9rRj1Z0a73dt
4SFCtOyFlFFQ9Zkf3PQdOQNZtGKSu77WN7ya+DQuw22OCgxaXnj48JKAHcy4e745
RlfHra5rcGpa1IhEGsE2K+4MSp4bzOhSm0PDXedagLDAp+dGr/ADHnJCDOW0hz7o
fo9QjXdKEoNxR3ZxbDk8/VH117ylrV96biXJyKXKgSmrK3DM8JtC0D73YbaPTgr3
FmpwGIc2xXRL+mznl8YiugGhgZnad+zvK2OOsuZIUwXHdLz3LI8zrCYxbdHv5vH6
f/XwBKUx68hNvyfseAhWV8pRx2ceWVweyncrZBgcxKR4bPACQkH/0Kz4gQbBDZlE
`protect END_PROTECTED
