`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m7NYRbA0hZFzxFaoLJ+ljSx/t27DwHf1iA5uEXN30aWIoxdZkDC/h68QVYzKOt5u
9bPltIOOx9D0zYwDLx6m9bsMMEaM/nGVPdGc2OzWUm5MZ/4ardrxWBn/X7l/t68b
9XMjRzOXSXGF9QIEZSiDoOf1Ujfh98a7/cQyZd9swLs4FsiHDfNS8/q/7Evjaxj5
JmeI10hkBhxOXiQWZbQPLZvskdpx+7nerzwTmiknQ/S62SaZTjSG+Vll/IaW+VMh
HeRJOJqkfzNDP92KH1gWsHDOBHONS5hMdR5JooJ/pI5jzLkqA8Hx4hEOrx4b/L2P
4iiyb3wmISwbbsAGwH08H2IkajQjcrTfp1pxcglRG31j044Byk2kyFl5wmc3aN9D
oNmFrNlu1QonqF7+oeOnwaQtfqU0PjsEK+StLHUeoXdodm8DoMbVOahgtZdqkREA
qHlRAkUn8qT7GRr2iQIvR1cA5DF87K55kBTt7MD6knNoNX0DyQ25F4skgTpLi6gI
RK7XTZ2Np6JAt7V9w3FiyLU4ZMzdsHpd9X7UFka/uXbvKLjXBKqkRuUVzAy63myC
vHb4Vha3heyEsq/efVwuMi/oGJtIrE+/S/SwtgqfucdrrnRyyWb6zINvkBNuNWyG
GYso5NHIuXG09EWdmKTC1IraP5ECFeAYrVIBFp7EBdfRDrj8n48EJ63zNFBOScbJ
IENQizZ1oOOgwZwWOt3diJnykh3xAZQJ1QxySeuHTOPauHEwkZwTjWuuHe0nB0S4
QF2WNuF5XZWuSYrrFWOrq4ENkNHBO38msio0XoVoj3CAAkTw0bJAU/LtdllOWbmK
EJBTh7WVlcMa33FvvMsTaRSBULORtmV8iqu1LW1GAwTsL+TApOSkOK1ngwDuzzNe
tn3jRiyVpa5/XyDdz+ki4gemCA5bphsjfAosPquYIIdRObVtVu4yvjaFsx+zl5AG
N8EeveVr+ZoFhg8O/AdOwYnaFrfLi5ws0B1TFHfsfaewQ2m+TojFj0dFva/l7Csv
Tc1HB69Xg85QyA+cxzE1IUTzVn2Y4eW0UHjntOB7krbLiAixC/Y8VwCTfRB2LD83
XOH/xe8RLlMhch9yxZ68W49+08AO35W4MBoipJoHbqbHDNTSsNlzVibP5C0ii2sD
62Bcax2cJRYlC1UOe+KEGnCfw2ESW0rpp3f/F0dRByse1oZ+0703ofUoWUG1BfNJ
vaEnZDptjVfT9Axqey/lra4EsXosMSakWUPCiOmmdiPJ4StZn/r19IMOZ81M6pXK
Za5xh8XmEwX+me4y7LlTmxcVDOcp+IFhAJ3tSWtANvmfbTMkUGQIj+2fDdgPTaEm
5cHgA5PoUeTJUqsBeKd2sfHz0gLYY+QYZtCSSQkwyEPS+MHOEOIR/g0WSelqhndy
PT1jMD0lCXXqNsdMA2aQHMWsTm3B/SiVtYKlUvXoNcEDHYDGnfJbzObz8L0cGuRl
gmiBcEa9GWyQ1G7/8lDm2PBRhWdrzChR3uw4n6i/mZvZNCkCvUB1HBHVcagJ89dA
W5/u2y1p6TlVDfK8q983oLc897XEx0U9pP2BsefKEr3npFG+JhRS7HRUX4P+H7Ny
TqnsHbno7NCd7Yubw1FGS/yB2OGmpzXlk3AbZTYTXOd6pTZNyqZgUWAym+3FAEx9
lKKOV/0hofPbwVzdTmclTdqHIcEiBGAlrP4OF99q/pQif68Ujb3RjwVrLcgnSvpj
qen4VmlEyCYZvQDxupZJNuaVMMYHY+2DI4uinIpmlx0W4/jM2tfo4Q00ngHuKKcR
E4uZY8zpQlk01umZTQQs7/rO8YzbZuYrHU8Yxb9T48XnHLdsMzazd+1GcqnxAyOx
57D0aJwwC3WkLmHI+B8lvvliSyXcdGRIdaA17N5dTu/56g8Ex0pa/OePP7qqAv09
PWsuFERFQEHkcbLnaEAxqs4v/aZwTU4J5b48CRw5dXnObPztWS9ggeKlXnacwfVU
8xn9D7liVYwjSA6Sgaf/a/EPc+5JcaB63cF7jU1idOnEKBiVJZcXaSYu4pSme/3F
opWBH4Q1tePXdY5MJPcWok2FAgzd8/ZUfFXSpp/NXJvXBbQ4HPrF/bz6FO8olpbE
Rt30sUIzQ1nh9OB7gjz2yt1GfI5ZWe8+5oE00Xekv8gxChPrM3bNEtNS6qSNBIW+
of0ku2luaObLlrL347bYEAtyoCfAMyeppL8GUPSb2/NOwlJwEqC57EQPm3OtwlRO
KRiabxuHLP1WKFjbOlhmo7LHOn16icI3848YeJFcZG6nodIjMhFGYh1VIBZ8VOAI
++jG9f0BcorygU/6GchUZrhqFDGPZrdlYxH7a+1bLahjfhEzuhKtCUrtrvlEk1B0
ppfsL7Xf8CVIqAvyBpNX40rTCAWKMGa+o+5EuT923B+rukH21XBWgTdRqKohYp3Z
H7ai9wVx3J/j3qSnkEXniOMoAQNY5N4OdW44bOOXo8Xef/RO3cdvzEWb3AfcDpMk
oIv/lx1BOiIuGK5dvH0m/K6DCI1vWuihOtcb0304reEF13fnzxeMYD3vC1gpVLSu
iNB/2g2F1b6H7lU6Ln37m4cptJho9z1ZwBD6Pvo664uoAEzFonZtqleDipb/0EiJ
8bPXHRqI9xsYA4XzNSllo5vCWpXyWbIcuxklt2mUnqc46L9TISbHDN9fWRa2sqmT
Ev/9y6f6LyPD8MUn4QB3awsRHK5h3KbpCtjhDrdIOLFPfTwEBDG7E3DhbuyL8yLk
yb0UU1eZm4lpuG3qsBNRTzg4qJzLx0tdZbjOZc7u5Zcm7r6F5uh1uf5HBxKef6O3
hddnqiwkBBE3H/3af55qe8X3q0NzpvQSl83YCNZAErlKfHmHIOS4ngCj0mKVKNd9
v09hTe9gk6GzfYkiRvvaYc3fVkZkwlgvIjc8OHPQu1dwAw2bq49kY7allFNa6UbT
PP5VHzjEMwqH8k+TRNdKxo6C0bVc0UQ2+3JGNa5IM53agLv7brXKwCk8sZH8/Cq7
40B43NSpSDRFq8zqjyTokKVodkYQIhZ71Leo1GIZO+FioaeGYQBUjS9WWzlM/+Eo
bTAUjsxoTf2zgzOpR+EYXcQJfJO5OuBOGPREX6eb7VrjhgrfF47f9mq94mnI+nTm
x+Qg5+wgEYVhJJGJ8HvBGYU3549FnIBjrUsDTLGQ8XMusMluaw7GNwejgdfC1M8/
8yXXqrG/fh3lx+BZA4lacLe+bINJz2z1dsyfrX+J0CBSINU+51afdkxQZV52xiDf
3eaPZg4Jq/mmDA/JXGs6thq5QVyxGeam8VtFM8oydD0=
`protect END_PROTECTED
