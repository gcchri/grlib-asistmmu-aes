`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kULKtM11pJvjWZj1jDfa0b3gwdcYxsHOW/NSymBNJHfyP9sH9YwXEgHfjcEHwQ4p
yP2EjNPEEE5n0cGQ0NNYMxpkwHtod6vNiDoCOPOb0YvtRraBHNEo9SXCtYcdaO+O
l85DlGi+ZoQmuCWukXp4xUib04UvGjO7wQODmjMvZn30Nb+eQqGCf5KId1U01hSk
EKn4/sclOT+BjeDEqs1D2VNp6PyKdDC4H4oQ6MjGB+TNXt/nfl1oFam8DYMpENaA
Lf+oszkMkvCMff00f8MZYaixhejTqt+1W0O9xsUuQOPh+SbXFp8FpX2p/RYzbU48
aUc8CKfEbft+f5XB3shaiNLaLtCiTXSlXxJxzKN9LNDswvK8g8OlnKIjc4gOu+Ir
4KFrjhIci1+vSWgiZraRPiX7GyB0jg/Dz2lZbaT924iMVV7aZV+oTZPCbP8Io4FP
4SmeLrfVMMhINvxRlc8b/Xbmz3WCzBuWiwxM53dbZ9DOHiguQ6erf2nrqw3/Gtry
306bbvhNorgVZBldCKaAoA==
`protect END_PROTECTED
