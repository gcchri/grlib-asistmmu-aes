`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xVtVOcwQZqxYyS1IosGNpH922UNrpcyr6Ka/600gmyuPgiOEPuMNwUrv5rMqU3xk
+Vpf0AuLE1iSibDLFiWV7xDUEBanRQ3t9qI2q6DAZlQe2FuRBNBWTQoxc9TFCdPd
z7Z25JAPNf2mrSXTdxaNj7TFFxKxMcNEh6XREOb8v5QxFvETcJ5rl8Wz9oRvN1pj
Nt/SK0NgrJ40ihcwgKK3sO4D9M02jFDONSoVbWiWf75Vp5O7UrxyBxIqbmlaTSLL
zysH2nrHxg2+kl9GfGfDaqcSPW7RVAMnbr/SmepAOVuDsNRkxaVGZ3qWMgcPmIA0
oC9jgNrmGo0iu+6Lj87bmmJDEmTAgfw/ysiQP6drSIBg2gf9q+ELF+YROD/q4pLL
oUH2UtHSQVIQ9FcMcaoGBxsqE+817vmG9roI8dETlQCPgbXZl3nfsnmtoyRbOWm9
YumfaBmEY/cuVRij/HzobzHQIT/rP7JaCbbgx2lp7QYaXeKMvxt/h8CUaMHboKFw
+RxGB4jyLsy8wcE+edwvUQ27ErIBUTAVPTb7rXP4GhNL0wl1AlmvRhLcLW+McNAv
hWz8sxorQ04qZPSaBfTKhDbclC1dV37gp9TvD6HN2RtACJ0Bj3rfj7uNFERQ3DJS
RPF/XNKkIwydH+G7ZQ/C9Robgngswwtc6V6OZHzQuRk2PptoEAQn6I1XGPecOXnE
14Ylcm6kQBemypyw0zEclihF8KGU54diI/aHOSrt8n//RAqw4r+4hckBQj9w5LOw
55zieYuEjNv+qmpgrYE+wQyCLLptesmIC4daq/uj2I+4pwgXtm6rh29k+Ehb4Lxg
bL0EwiYnv9vbGk/GjPGRuct1SGWSRSAmgBOPQOXWzbrw00mvJUbViwAmey4zrY34
+mxwzPjP65nalwc9CENS5FZjOGo+TvGEiyMMCHw45FeAQVu+EXyhGGjKUM7/jI64
ckUhBHFK7/ICvWeBo2pH+5dOnLLTM5bIqMyve5azb0hjlVGX4b0gFGMRQklfFpe9
GajNTIu2Ogy+aGF8UtqHGDYAfiR+7+wKDyHJgHc5dNBn6s8FDKodTr0e/qsJwiCn
Iw9kQnUQDopVDDlu+IL9XGe1Isz82m9I8K+afvgeYoG7xqKDPnYV0Qj9yr8rEItR
JkcwJXzEALc26/f7Ep1khPIOHefgcwDh1s90qGUYPgCLiJSnnxr/TvQ7DC2yNn3H
3b3sKNscWmz1XHkSQdlP4IHXj+IMAjydF6jsYWdbYyiLjeA+mEi/RDyc73NyHVty
AqoaNNKofo0mbvmbCwRemfT1R8HEixWyRU6zzy+OI+3H/SERRDTVmm+fI/Whty/V
vJzRnXl3ubUrKmL4z8npeRt6r9nTEHzQoQxIqSmAynpH0yCkEgRDE6VqVmF/gyiY
RF815xDOW6OZKZYDjcdN9rslZ7RCGk1tiTOa/60WvHXpiiLHEDT511ZBhVb9KWef
pUhiGIaj9EnbvnxS3hA9ybY/1uk+hxwTV5e+OsOOCVk6t/I4LqljAvchBVJDeus8
JFpK4I9o00PqNbjvtvnj6k+ae7PMbScQC4K1kMrOx5R3//8KYZOtm0G5qtGCsozy
nvZeIQMQ8pN9rGLZhAzf1kRSMRA0dxTG3it3ruYZcyUhGQT42I1ixRkfVPJslc+Z
y/FS/f+hTKqhbGtGpphI/vsWR2glm403vaWcTezpnrS+YYbu7NZb0aV4qSDqqPzj
DInOkS3AVfJggx88l+m1ErVS4Zm+xc/eD1AHKycm29kD7ullkV1a7gDrFYfhBb5S
Igfjz9mH7rfReUUnbH0QNh7y0FSwqdlWZ+iO3HtDC/ISQVXBk3z2nMOJYN8DUk3T
qckPKPaiMi3NLh44kCUYUF5J5JO4Vjkkfo+parGRaabGhghpBzPexXDXxYoa97tx
gYbbu4KI1UtDmDgyGrmOAUzfNwsCJzsPadLRuqvKR+JtSswx4aqydHWnV5a6RWvq
DsRp5/HSxHT9Q1oAd8gYTAXEMs49TNgVEAVVV1UQo1/6fUg/ZSpvG0N/pyUYFLoE
F5zpKpLCzGqnJPtWw5E/E8PSH5C/rO5ScznI6g6k7Pr9Qu4bKPHV9sVA/7CCL82Y
75dK8aKRMgSHOF3DBmqWADAVNE+6PFu2af/CcjGYJMupK+jWU6VloslKSEUHFLZS
ahZMtd9WJov0q9dhXuqMNexLqy5S0vTM4080kGPAa12+GpX9zeEjof8B4WdCGbyf
Fv14TxEeuyjM58QwcNwMgNAYPVc4GpUMNIetnqFUgh1cLyUKRIX1inIPifD1sgQx
hXuIn2/6QHdpHjdJAtNaOHHjGdDifJI0IV2uPjAB4j70pRAjqkC6LMueDCeKacA5
DmvSNhUI96uDaAQe31AXiivl/zRDR9pWUpEjdrrLs2JUJGJWpEoarkpzypBaif9a
6AB2dq2dOCv+Ks+rrElnSJr8QY9lF/psJeaWQTrzbuuid+UTvpxAd3sLm1wa/fmD
bgZKiygkw/Vu96LmbHJhxcEngbxTxHNQmURmXEwZmiL7CsDdugZqwHlTRlRZWVUW
Og1uXZhbqkkgghbyqHL/fLQi6mm3c6qKbin9OvOTLYyOH6nLpnTzs3QUYsWb1hUI
Yog4upLp3IWDt44eY2Mq7x3IvSzqPTB7artl3FGegE7LxbiLBYiy6WKI30o1h7zH
qx4EPCVwBi3WUJaEjMxODe4l65TwJrnhQTNEdKQVaQgl7wskQ/ZuMz4Lmkba/Li/
6pWPf9iatcyShL5bIvJUcm7uT2ib1BFT/0CsDLlS87Nz3N/97ykYv1EQn/6tnfAk
5CrrMagqxpZ6ZROjI5qeSuF/v1q7fIeHsUyZ2jKUeeD2GqKbGQPMY2TY6Kms7wvo
PBPZfloG/lpEpR7Ww1U5Hi+FSGRpOLN5/7B1veVgT5dZGJV17l9ADvjJzLCqqOEh
ysMBSijFMktgkWdXEKoJcCT9hb48mEzDt1pcqZS2KFMcrlcV+dZ+F+lm7SGhbYxg
qeJWadz/x+mxMOZ6jzgdtV+7Zhdq/d4Rbm3RLyx1uFPsJ9C3FMBLabCirE62yx1t
AoblSFtzT7nDYdwdtzEUqdLBOzjjwO5d3w8e6T8mhhekc1l23uv4u7+ukNhMdT4o
wJ02RAeWfmd+s/G2ELv3cDWut2tcV6edOZ80LUEwzwOU9DA+ZUYe10xpjYnlMfXj
HQ3zvYX6Cbx8Hy7wpMguRzIdWjypBvR46CRBzGXG/zjbGghbdnq/MPacV3MOeW57
b7H/1P8kvYg0VaUTU6ZstX9yXlkpyHQRTMIV46oU6wjZIaFO1hXN0WWAHyTQP8yd
URHH+ozHyolkuMYLOuLsCp8ch3/XWIlKxzlnz6WbtCb7A84o2aoWzCjLPc611/jI
h97kzp8pK/stQZuoFxST8wP3/0uvb1ofWSY3cMZqExbXghuWDjZllTaPm0rCm+Wa
8ceiTCMuqXYjfsRGK1N49kOe8O+Qzao3/ue8nngBV5Gx6+r2BFn5RjZgsJoV6EhB
u6hgTkpOLlZC0td7Q1N0D+iZNEPKOYKrzzQdpHmr8VaMRtO8Mu71kKZcb6sj3txC
HP0wbvbAV1OOF9txbQUi6//S624O4QHjzzp9+6s6To484CsvrzRnRU5nYEKq8SQJ
kiY9rBeW7NmYyjaY6H8bYqAOV/0DuNMJ7WWJq1u/c32If2eMLRMQhPQfwqWyHf0P
16NizwMvmEUkszQBEAKU1sFzHJlpE/mK2trhCIgGvRikytB+GZwdYzcGRTcSgR45
+N3SxeYyeRQ++vNuAyhnKEo0bhHuVntPU590gfsileqBbRy4umKK7I8rQ3VHfRCG
N8xeIzTH+YSliZjJ0VpRp7hhudGiUZXfzuc0HYwN6lXRnXSBaeW6tIgWVWdkPXy5
anoN3RrwWwVJJw5PvLmqlTVqjESw0TxfJ0nWcYITr1YWwztDWRdbF3M3pNM8Z88Y
SmKuG725plpXSXfH8vh9xW799cDbVauAWm5RFwMm854abFcGpZAdZUoUbAY92vdR
I9asZfg/5ox7mAvmR70BMO84CWW48hmP88rXlQSe3CNTvPzYg50KQ1/u3ojruWwm
ovT4Pynm+viceeMLWQYPu2tjC/aRUg4q8fcy/OGcsZJznv8/ZagNZJUOlgi/1xe9
AjPSut322Ue2JKSf/D5gjCjVjxl3Gk85dldw4W3xgLitY50mv53KBo8S+oNje9Z9
32ePG2dlV5PpS48jW44u3rXIHb0YWnvOsxEINfO1RD5NBKg/7528OJACo3PF4Su9
QK+Mn8GuI2fLLHZfHq387HcMehPtRFp8Tjz5w7B0QJpXrYpeLuFxaIZMyXQz5vlx
FO2pc2AxjSoJ2j9HOTHrfiipcxqvGfOUrAHf8DFBayPG5V+pwt1OapqFkHHbbGkM
oGD6xsNMPebrz8fsSe2vqdOrTdoPI7QtOVoYB/xPju3Agz49FVCkJHFPoPJnI/Se
/Wp1VhkrePL1QUJTbqHtNUlFpiZ+OkVWqY3JgiTrDmQKmZ/Gugtc8SuXd8jTYT2X
/JLFFjw4mO8Td7cn+U4gab6nVRBWKyZeHeVF57N4gkMpP4PDjDVw4X+h8SZcKFPk
PVPKCu/oXDCfIbNprQcHSyg8vWjhWUFoblqHfObwY9NSvfZu5fILbGiwTSVkLbr3
GY7rGit231nQtRPBkjDf2IgNZ96syxfZZENPXmmMax6mqQyki2af9/baRoWCOemo
+hC+R5S4ESiPRKBFzyBvKLMHWSwjabihx3aKFjXBR2IH8nhN816ivQQanUxHgZRp
4+KGp/AHOhPlrJHRm2jnVo3Hz77/A1Rfbt5q1QwMvynZwSoLn07h9O9FvQvyhsaM
wdodc9gNXCrtR+o9exgQ+2Qp94g6PGE8UZkGV6lbr0L6aig8p9Mkfs3gwzlAusBu
Ui9eyp/q/iW5xCSRwOKO7jIdpz/WVNXfwykfYwzg3gpEL/lHjavWtkvQnrQRZFJX
l4ihTlS8iwGTfZ2TXeCqGEE1uyvqVicuiyqwTtLmdSnxXB/XiH117kuKmn/sL1C5
3k4fwOlO6ahIc/iH+t7rZaQ4w5osjV3ZmDIfSsZwMqiKm24TguRZJ52RZroISN/b
vheNlfaJ7oFTrBcbHvtse/Wz6xXCI4x+H2AXVd4rmKmHbc2EqlVLPQCce90uE3xZ
t62LWSLPzJ1xmWOniZoKc9/+bXVxfysIHzGaedOUBxDFuFU0nowZL6Qxvkhl9Pfv
vAsrd2iRJCGh16l/6IMPKrO6bq+A2hrOrtuIcozl0N3Bp2vfHfCF+nkVy6TK68TP
vjJWZXV07PRWcRmzlI/2Eu5sXOUMLXuxcWC3XHJi+Iq0L/V+eNOknti3ovjylK9P
UB/dhn1vhHV5W3PtaSmHw2FV674n2ICy7XK23ypmvZcyfIO3HZWPp7dF39bVyEbo
605+bQeB2Q1994TIjESn2EqFYHrI4Kz8/CKCkUGf6AzlwZ8pFGcXvqsOLhCp6OBU
738/vxgemeISq/fWotISnqFMqwRomXsItP7pWf3fbm8txVK5/gf7NWXrH/9trLaY
w9ILl8OfgX8UhVObvLmKBcm/O/o3O5IWDg1alrvITma86YS8lLqa89/7QD1TmmjZ
8BcfW9y6FjXDTmrdUbn+hR3c14I5o60MDTzYxDME3r0lR1pkN662SXAe865h8hA3
IiEtWoKQLpgP60bJ1fcFrTY4NiHh9+3Gk1JJ8k2w52+gIPsJZO7MZ5B12ysjAWRW
KEMfuZnuPdyjKIdBKVpCHY5L8fqSVOuHUeTFwQ0ym4jlE7W2C/h9AUP117rXIVgd
0KiOWiUO3e/3phy1kB061WSSxd3Vc2D4su1R2Fi3Op2b5oCLpz5xKVUHR0Htd85n
QhSxqA4AZ4cxD+8ubui5AlMU9NMzmC98ZhIHHfFp3I6l+qZ7+q5tvoXyfddnWigm
UBwI/LLdT96mu2k3E4Nn78H9cQKrHGK/xM+gH1ON7aC2CPJWHiy0eN6CpYTa2/hI
hia3VeLZLigHlG9AyVx24gO/DsZVeVsAt1Ffk9azC9DvzxA7zwfCqsPbR5sGSeOk
K3/4vLfaEOFqTMtVcvnFRvl1RD7rdSrx2R1tCL1WP3C8FiFhUj0lOpQ+phGGnYRM
Z4HS745WqUp0NJhg6kIA+H6/DKoIMiOWm2HQv1rLFGdozz4rnU4sxtPBmj9DqG6Q
Uoky7Hc4nBNP9zetsyLt6SXppmTuEtsOhqiz9pTEkUSDi1W3csYSkAyZEWPZ49CS
rEl0fGrwQIQxOjE4Lj0cE/rrPAGRrwpBbzX5caYQQzcbz8Vrd0YcPp3R4307AM3D
8Au5gaU8+1fUW3xzHCpwd58+qLRD3pbSdkrRmc8DAJIrp7S35TfutpN00SAwd7qs
rpHwdYqrnIIrKWqM4ZlXETx/Vdy1X8we103t2NY/CWIguGvoMcVf8e1DsXqfNGae
pMyxLzHANwu8hxnKdIvw5Ah2su3EGeNZGbXsuXHinmT6Zk4rNeQuye/gUin8+d/Y
oJVQ8JB9A3o6roqkVQcco5RlxpiEmjJbpR3Kh3dwB4B6R16KqN2xXEtdo1y92yC7
2BqyoLkBGy3cFDK3vA76gsUGopnTfrKRkqZRBTl+2VZc9mEdW8nht2bquslUuvkB
p953wgZYk8V87zrBVLcz5dkW1G86PuJP06Yj8l5aLbSCzIuoqSmYBoKiFMQdD3/e
jrn0MhlEr4ZN/ndrmhtP1KOnCtDJBoDNVeDzz+RDviY57yuleWlb9GqzmIiLZoeG
CmXYTSYypQei9Bb01IGdx3qaOyHLxa0L0waf2Dftw7aP+RxrYTYOBRf+ioEgREI0
XTPTAjwvaoImyiwMQjhT6CLjG8phVpuqdcTRHDSciQBbHQGexm7aMqSHc1TjnGRz
0iUtMbhUYrPIdPK0kExF8KEDvFi6Zf6Ly2MmbALaUgjYWbWy41tpYDhT5c+r5njx
mUAXcgbwIcgL1aWMKZt8cpI+tpaMSkeLIBAIi7LLL8h6Biy8UB2IOJ/Rv3hDHz05
X/gWVTSPWT1l9gZ0EXmxirtX7nq0QzLxejVeYicW+FzZMKFJY6p40vlwznttH/aC
s/jST3GoGNXUrUu7DTVK7YAEuYfEUaFv+0gA2+L2fakTHF9TGonq1PN+qp//+nJ4
X8qvBj3lmGFoGzih2TAWDP1JMq5mz28JeLoM/BmDfIf1fkBxF/WAAqMO4ZFtrXIZ
V6b8A5sIhit0lnM4uxwm0sNCoFs513v5ONnWxsAh/vjB7YUULR9GyzgR0hFjskqJ
1D05FvaoBt9tc/wvoToakoT4QWgt0gczByC19aHfW/xsOVNk++Uls0e12FKgl1fx
5JM+fqeOhfVzrcdGfrkj/p87XlTnJJEetbDSisf6xHxsyGNa5RQc31fPTL0nI9gY
+gIEBB4AMKVgmrIsRD32vTQIjAOiFq4qRBCj2Y3tO5QyNkPQ9pDiUoCVJLSIXuGX
M87ILInFyC0QbH4PO+zwfZkSU/ovhIKk/Fl+kXjyHXNI3QUXEZ0v1KHIB3YepvKP
UijeYUqU1vxfEFkgtFJKLmvkADpYdZfwyVBTRvwi29arMuGbHbrOt+OpLVjwT4l2
4ZMK2xMEkzz7nAKtpLT2u5gHbMHaAVAt6nmVTQDT/E1ckSCfBR+15fEG4rWfltMG
GU2t5SJBew4J+9utSFXLcqooVxwEL6UypA8AOA9jl5cFrBZu+SFC7SMRwbebvk73
5PHInuMam5f2t+FxwC4uAXQVtIDZC2Cw+UstTqR/yBYhu4NH7YTgBlUfMZd6sFJf
wYtlvlUqQAD2Ywp/azDfu6M4FSuUe40nRmE0FJCWvjVscQSHeiKlhwrQDngBqLYY
ExNCRip0msLvtJRYuoAEyPebXs1M1fLNKsKSjhOQySUuZIu92FaLo69uMrm0QbDV
dIYuu5gVv+cgKsxO5mS8sxw5OXuuOfZPYjdWidS2cxoXZzvsueaILHNL+v+8efZR
xhTg0SLrasfqg0ahyODDM6FZdkh9Oc/w+Rjf7GrQp1SQsGFkNLL02GLK/lsKqjqN
FeSCBlzc/+NUzZvAe5dg1KJjKfpSiZqotaXZ72RQmzOXUuqTMhOiJDY8dJyM+9s0
to7mlIaM05ivHWSF6n2M4EDz+tSFuVDd6Ko9Pd64aq/Ve8S4PMJvLr3dtHxKtVxJ
TPyzLubrqgs1WGiy/lN7eVtHeyZKSgxyoXMFsOW/1wsDWeCjvTLKBJQl8GXb8kUi
oohNK/xqoHOBRTLwSRu8rtx3f2rfwsbONuZdS685HqmmvkCTpzUTlgxdjvkxcUYX
vt7fvJlSANLVlXGPGm1mQ9rHEMw3O5vq9rfUULrVs7JiuXt9cVc1uH4/RvhdCcum
LM6jPSCbetb8pXH6w0thWZKoCCaOJB8DxHPvLq5D0dXTSLzfRnabqGCYz+8b+8X1
Mzv8EYYMz7C8qTk3f0VyEs/TkF6eqxRnGSkl5uvi5DaJdMJwXpvdi4oakEz94Ur4
Et+8mTDVYZ/WPG09ASc3c5sisI4RYaQfuPHe+PMJE4ow//5MqHkZwZrWSQD7ZRAZ
z5upAtF5bveQHo0mltjDZKkB0YNW8HeDNeQ+d74cuKdkuTtN++dp0JpI/OyfNd62
mDkpA4HYRS0JE1C6zXkQyzFPb/zXLl1RJz75xeFuxneIIGEnvAkCv8DmpZcDPfE4
t8xA/BsQrHd4oNTi0xfLdFcAPPdXl2WMD9x1Ap6UZOqJ5O//RBeI2+43+yezsNiS
TVxvybcg4c3fpICAELNhmRJE16mWPWOkb8xuKBOVhiwob5VGq84z4b7i767Lj65r
wJaDb3CBrqcM05uzIEDiyQi+6HtUfgX197zx27boVZC6av7zJ5N9sIRp9KW3CKXG
Qju4ehaWrzwPyijqmzlxtP77n1pOKOybNhglmoblHY9COFMb9/3V4CiQIey6G2Bl
dVVlfSUviCDOWC2K/W0xw0Vjnf60f+TUSImqd5tHDHISjKrVFB8XrskmgGJDCZQ0
S7kV78xYKgOLC4CHMcXRRrGq5sYjPmgCjXISU1kkaw3JD+JpFljk+cDqZRiwsefH
WVf1CV7EOuR8Vjoo+3LJ3xir6Vb7esf7mQKKsLU3UvYZsKR7KRqrdkFADnKMsJpp
9ByQjmT1zogcn3p0FoK4ms45Pdsy1IELi/JtJ0hGTN3MvrXjJRQ041urDaMQONQo
XiumYf+TpuFiKG/s/zK1qFEHOB687m0g52eOqZM9C/IiEWswgiQUaxC8tBFt/oOh
fLkAO4JqJVJoaUTRxO+gSlDsLAHOSuy2UxYNyzQRY+d9h4GeV+uArjCNoLAsFfVn
s5rjdnv8wye9qqM0LU7SP6GXpj1vl1Wur848QhQiAmOrXpKQQk6ziIrIno+EET/0
rBn+ncg7OmSEMvK+JvHNlUdFSyVLVOMBB3RrlA1lKdgWfwTp4EJeqj9RVKnAvKZi
glUp+aiYrT/1MW6NzR4w+Kz1UNT+147Di1lIR2/8APWXz5nN/PqRey+0ogsscqk6
gt13NBw3bKODf9MoEh6iBGPK3jKR7SF9K74zBFirKqi0eOjOGUOgwKZ5lHjLf/cb
RjtVMJyg31h6h68WUJF1HAa/vlgS9n9kRE/iiysa7pvKGYFcFZsK05tZ6EV5yeJZ
EX/ekCfFmHeHFMRVeyY5rsSDZipRiSwcRtE4AOpjumD0grCq8sZ7+0r9NaUXW1qS
4EELwdCBK0CTK6zkDIewClyIcQvU8t8ObhJ2hvMj8VgLKB61Rae4/osvKTP/wgQ1
3mVDdUw0ks75ImkEPglPBs9Zikd/R3a1I4WSb5zh2/pPFLkPwBpoRznhDPHAOZeS
HfeOXqWmgAb6iSjj53uNl4cMg7oVpaur/M5pjUmWZaTs3f2XwVrb4u0/+XdvzMR/
frRW5jodtwKr8b2xFhNMLiq59WDVRRy6VlsN5PzK9rs6/aNUk11uledlbb8wodLv
vUEn23Wvvho3uU6YOVIW0q9m46LX0GRKQLFjdLuKfqq2t8jIzj2JrnJ50d8J22JM
NoXBci1KIZaeRu4IKlKNoXGk2vO3YQYydheA/zOXE5ypzje2bMyvZCrjB/R6AIJ7
/O/0B0XNW4uLI1Y5LGSKV6pew7pkY8+ZmSjVlQY2uAKL0jxSu9sOXfmpONaCZ91b
LqAHKC5Q56+Q+Ogz7KNoFobAMItt0DPKH/J6VZi61MmBSw5BVjAqZtcD9wCU2KlK
OuyRB1/5QdeRmrljyEjl7TQYdbzk3mci+WvZjxwyPUf1TEwAryVlkjXpAZylbrMD
L8vwTZW8s5bhyQlpUH06SM9UegeLz6kVIQ8prJaQQpvF55D3Wqgx0+9K5OfFsan7
QGG+aySS+IJ6kpeOF0diHjvNnxobJryvcs1OSXM1R/CWq6DYEuEvSNNwn620VWRO
4N8Hj4uIt+/17agMPDGb049tnMM2iGqnRshFwNXo4w+/4qNallmahD2G/HwCm4Jp
k0wX+Rm5msvQtkgkQ8Se9SrYvaNJJPPIO5/XAlA2Gtp7N+Gce/iC770sxFvRTwuL
BgySs8z0t66mYNz8KwRg4lyYY4faSEOLqyL4mz4uHPt2RkSvKzhv60UEVt6BB/sg
G9iFYHi5TNAVJ7VPDzzMj/py+cUevqLUxudJMgA1k7KeX/eV8wmmiji1KZvnfeST
EsqB0ZEfFK54iz02Qc89LTU2urioMaG6SxbsFB+ELfLhwG5KEhTUYWWtkrftfsSz
j1QRKQsBjzkrRFhPjgWi2g1xs5jiLMJYUqUnUPRi/AC5S39Rc5Gxm2Rr4hX5Rdbt
IosVO3hGhFEtjuOPTbhX0A+04S82ka4sjQ1Z/W7Cj37c3BtxvyX/Aj4XQtI/96O6
hAUsWZ0RxXkQbyPmzKJZWHIwyRSy2/kpYwqjiy2ZwyzqXvbrrUR7YfB3zUkYTuxw
sANRO4JsGCuUv+Np2r3oZ4yPUeagWN8l494Lc4fJGhx2PgJ1DCXfgGvBncfePYum
0S6uuAdWzwVtu/1alaVZiIOy66Qy0SpIleXwANJsi5G0zcpaWahkwF+URDaEYUyu
gQKYa5eeDJsWSf1bsJggTBjRZk/dO2SpnZwg59tkQPFPTEpXHwr5tRpJKaLohBhp
YDqxu8HBFSl3E528hvE4Tc57y5I4yljXBhs2BDnZ74Cqu2zhR/IXQxlWEAfv4acD
gsC3A+IT09Ts7qn/FUGVmD97kb8pnuarhJhJ8lVvHTcgPtqj4bNd5TjMavk3E9TR
1ntx8Im9WiSTqhfGFNWhWnsHlATv9llUmOhGYmXyqVbEIeaZ3tEV9nTRj2zBFV03
g2Pqrene2yAVhBBnZdc44MPauCwmSUbi2dEPd1NvTb3IExGzGWON+U6PhLG0XtR/
lbmtPWFm9Q/PJlA57ky7103haq3VLUMxU91IhKmuZv/zlpzop0DkivZSZbAAYt2r
SYEltsrxaNENZ629ltRLrGY+M8NyE/enIKGuZMb+S2WHZa2as8Fk5ontQexY13f2
IiKfxw1nQGsQ99SXGEUUR0EuLSCjfajEf1UCUKvNNjcsFwzyvQJE19ekjV7UYhvt
cCTdObaoXbjsmTN6QZSd366dBibOLFHiLccgEc16L7MlYimcFlJl+QgNz3s79ypf
cS3r6trXBPMgQtSrDkct4DqLOP+PEoJpTwfnO8V4UkDev9vsUQXPa1+NjKlC5MyM
3Jlyww7qnXpfO489Pkat1aSIIYFVitUYWMImVB8YibQIzJoK7H83cZ1Q075A045M
dvkAL5o5SZ6CXYVmJyWRYXts+3E41bBsxCw43aGXkcIxa7A+jZLErau3PndeTBMf
bQ0dvCSdK350OaArobveT9cx3UyTytNbDsYmcHTePmCj6UEZTXLiR3SysO+arCkF
gyWaaFM5tAv0PgvAr7xCTH+NDWQ+A3sfzNy1QQo7LQpbh5fgNA1MojaZTAXLXY2p
OVkSAYMdZTrIwMLZ3p5hvfMW+CJxYQWUOf/GE9LVUeEZ+F2kR/CrWf+AazDhjNU/
5zL+MABtrj7z/ngownLgjPuFSTnZbQKfxYIiNLR/MWqoViAoKmlMo3HzL5TGdQbH
Do4v93ytsg4OzGCXc6GBvkbWLQvPgFCL1B2qYV82bHwUWRdxUtyYfsRs8ZLja73K
IHCPa7nwU8qhjSAo+TDrA0OKG9NTq9J02znbIrfGYTHk0LeRKylmie7lX4WrRXih
1ii+oOmt4gy98IBRlN0WjQhucsq69cq1XPDRLLE3zo9GzRuS/omIFv8W36lxN/9J
kQA/O7bfFL8DGBaodCGys20A2dnt9SMcrBGb06Xahn3CXOOYNsKFE1EFpUsjSf2W
l6tLJSBx4mf1/bxD6g3B9xB3sqI7UiISX3I8EmSbgIrXXp2SFUcHHw3IBDe0mwPr
GZC2BdYLvs4rD0hJPyuLgh8aEUQihB8G37aFktxW3pLCoR6PI9BnUhAud7u0YCCc
e31CvJcp3V835CWwPx2gyhCjqclt3bfKfbvz/QXzO6w5wqUQGvqlN8HdcBXi26Bl
OGrf2H6E4K/nKEgV7X0VgZK3QcKy6/cBWuM3jK2M5KGelsHjibf4MyqUjRcMYDTP
w1+eJ9tNphK7z/JuVTIrFy08F/kpPYN5UL3h0N/6+RJvLrBoi9zkyU+MwZT/wu9e
Uq9pKh7xXV0x7qabb5utQNOIrdHiZBVP6fwfgsxEwwXhPM3rFydsWtNtiVHzdMJm
/oGXzoqEGrt/a4VFgHJGZNpFxC5Ix/bA+Ba+WlpQ1EYKOS96XNs71IiuvFNMN65p
by+ZrV2YRYpQpExlpTU/xy3eTYbj8+4RiU84K7OEffrrqXdkOEbzWszxvLPLXgyW
LK8spmOfhwJfu6/yQ7lWymNjPxb5o9+kQF411WKDa0VNB6bmiXGpweNoMFv6bYe6
3830juVAMVXVqW3udrqn5m+DfMcvPmPWVfIg9BWCXNXG4UVW+7DTtTEh3uKIaodv
QY7VJPwIZ++A3oZeOpsmboA9mrEw2m2OwzJqz8EZ6O1Ah1RcNG3DOMbmRyZX6P6n
W2iYUf9oPyhqiBfT97ZzL4alHUjt/0QhkwuoSkKwdzRcLvhoa2LYBLuXFcMZiMys
OmdRe1sFl60fAjNGPLVeEPa1Wu20GKKDW5Aqpyy/GSK2UEI3L534GVCMzF8Pgl8n
vSVWVnFOyf+2E2C2XFfcVS50rnsEKJDlHOiwkBsm498XKrp3+B8q6Wxj6zRxmYt9
1WMSBxrvbVQ1ZGxanWrajtcQBhvC/w7A4ogLTUCvbBTDzM+th6o6WrBWtuTLgA8p
zPKK7KFyXOvNCX4XD93+8G8f7UW6unUxoR7fxnJICjK+WlxBwmi0+btZJa9g8MJO
CyFJtj9UZnL6xbTUctX+0bBWII2d/t8VN5GITUEKicUg3WhFRUqzFTa/jAH987ZG
mXtZ3TmUM/hK6rCHLcRNoa6Rt5m78DWZLz1lmtN+4DjpppBeqZNHJb2dHqttpF7F
duS4bVu0NRIV8BZ5+ycPnG7DgIuoBeniWuIKRt/XC8QBVL54zR+QbYh6kZzs05Cq
F7oolrmqehseYJH7N7LiVeJZG7hB4ILYAtiKNZ46jQ7S5+biitSTtlH0Gb+d+G/z
68qqUIAXpVIPCQC3AJT99xQ3M8kUMVu4ip3wNqvBabAQRSOR5twQihc2WZuH//tM
mJJUaXgnsvUT5DUnLXUBDnLzlLTELCP2CVk3Nx4T6i/JT/yM9Roll+qHzy4vPcOz
sEro5oROm7v55zt9KB/cwxzYk49BDiRFY/Z+Vka/MWnOq9ytJy4XsLWjmBsmWMug
2tu7RJw1PjHiDGls8cpuUlbDW0xWs7ncawfaD6DRIyCN4qWoZ6ME/AqB4kabxVRW
be6UTEECdhWAcbnKa6vI7o/WZX6ZriC/DtZODZbaAyVSFAYoVnJw0e/bdEQQIK+0
02YiBr76R+KUCOTpFkxtIysoWrw2ng0XxWHwnKCxtFwW8zSVXPERBfHDeLUfNCh4
1Lfh4med/DeOr8iglNh+5zxSMWMmK3JNQp65IGZXRKiARtDr0NFvSpdcGwzz84NB
c6GAJtDFtZFyCtmgOIkWqykGgWNwxBb2V/eU0ZCG6fstugLIsz/1AmM/mVp63gfQ
8CWL+++przt/+XSrqH7XDIc7o26Cq3ZXRCSlR5TWniBbrJn7LZbNZ1hzAn36vRTz
FgTnfgu9igsABjvwdYzK+qg//SUjVKh6ZqwDajd2ABELOH2Q3f9QSVQJ9se36veP
hSeNim7HC2OVYTUapW2s7LBilK1J1gkcDvDdeKIlQASqTQ1c8MSidvU2joAKzjFl
CUddm6+XD5PNAMKd6vRs3f9w4gEbHYpiKU28Z6+kjvX2FdwynHdzvF8oC/ym3urC
9n2EvNxOSBTk3i1GU8JfMrW9CpfcghWuSeH4WqbUdxTYneIH1+wELn9+4MZoOuXP
5IbqMlFSGSckS1Kk3xOasGiMgUtItPKqVxu9Eil7zBus9svS9NnOtewWGIzb7t7B
IDopjyj+Edt3AxsBGsfuQ5rQcDcULsx7m204CPa8mA7OhU6dmlLovRnoKdawwOKY
JeOVyAJoeCWnV18ohBjB+YYTaVvUoMZfUDBK4sNr9WVNUgPH8zkRHZUHDVW/x1vU
5vdcAC9mu0jJPdXewctWjId52oE1HiZhuBnedzH3wCwoAHnvDgBE+rJOFfWYr/wZ
laqNwKjl3voRRd9oDsJuD4QaaziV6puXEwu6ZfRf3HB59pl2VhVhZ494Enq0sdsV
yyRpJoNQ3pv+x0zkbtcvbsvliUBMpONJ8Llg1qAE56QakyrTwy4SDUfE4HRn3MH3
ldYg9YQMDzoRUt3vnHRdpB4duN4atjGDFWZ0vQWxeQWqEOA3ovzwgVdq34+o+UHq
nsZ7tSnRypVRCBA6M1tEjralNbOT5MmB+u1/1S2fsc7z5NHDwvKK4/aFmMKGlEtz
kdJgCfbl17tDDgb8IU0pqRKkxvWGXazGq8fvIoeYtdahX9K96HgY/cQwIeWl+GCJ
x5UgMav+wTTTJWIZCXy19x5HjybxqkqnWPJU+VDWsOAhza5vxYv2Yi9TDdTdZi0Q
RitQ4/i+Ai/lz0fvZv9fg+YK485ru7INeya9CfVPbw3zqflJcsHvCS7em58FB1De
OGq8r7uSv3MP9K5apRHxcisJx1u7d+1Wob6PPqcV5ctHgA8pn/+7AGDtvkRIV8oK
loqi9MaEz9HnzjAMmOglbX50cgnX2B4Ww71/6sl8IZeiC/iz5scL7Z1DdJDprSZA
OzrXgwD8dLxMqDftaWgnuGwWKZvBibTqGi6XreJkChpZNPqIk7/apnGUYla+3451
O4MdLDcVcDl+pf5NaQ1U4kySsSM+ADjsgd03eXRvgmaVmrCrV50soMEHzBTKE1v2
+eoNB27bsZQnrbTZ0rFwV/o30ndB3dLGbPApZ2hkbF4s96RbqYUBW1ffK+gpw+a/
Y4K46vK71Rx4Y0XQwu62F4xcpqXteAe4QoJRCfJiR4/TLHnONk0CsB+avpZkGelC
yJQaunk2thvywdZrsUXV+VIL+o4mtqh45qloaatmCKJhwDIsLYPtAmXw1VIgkcf+
wIbJDKiCO/dCmxo3j7T4B4grkCvtJRVPy0t9k9jLQ2mx7i2jDeppbHQIW26JGw2D
/QQBk4Pse9e1xlp6Siz2sHP1plUXn7hvk0xqIGDcGYYSlW1HQSxlHtl7xKMTmM//
dFGYVhGzxAfFRXMBwgLgl0IQGszcG0CVWTJSat2jfsPuFja+kYLfETi72a7VmPMZ
DdYJy12XUtLm2/0DqpM9N4djscpOWGrrdoxspAodTWZnqDWN0amGVYKKGxUAQYBU
m5PBSNHK2k5knR34uF4RwbEE5gopIva15A9Z/rvGpX/r2HrWpMMsIsHyBMo1vvsy
5GzJlqT5QwKaweHOpNkdKe2lHcYN3v8/ghxMNEr5sm/CKIHU11JcTC0dtT+onAx4
k+5OjxWbt2Bbbot8k/Wyfgxdv/TgLCrOpA2jj7BA+7Vz6xQdtS5YrUceD180ZvKB
SmJsAiWPxSCbS3tdy2G3LXXcqlb0ILy0Ro7CC3m+2fsVRmh+cregLLNK107PS+kU
eAR3ZW4ZfucH7hUYfYQ+EN7AupOjKRtbRngReac+ldZ/0G1//Pt4R4S+yyTASKuf
nOEpMJmacUN6lg6eRUGl7FY85cdOTk1LZPMT7BFLqYgeh8t41GJXC3kDeXP/HLLQ
vDHqQiraVy0abvo2PuA+DcXdFSKCeThQii3oBV0b6XepJvMsKJkQwEzISJSNATab
L2U1gj6kT7bNIb1vZ/YVso+PChC6RvyLsxXEMWAaZvKxn1TSTHOvmCH7T7NcKApR
rS0pJ+NZBPtq3WwslBsDCJA+FErmnM/jFZgFBmAfjH1yP7s2Eqq+NZTe+odJt60g
M6eYExiAD17j/ADtPY33HvZ1crFCvjZuxm7isWzEBVbsBbbO7DpzIYpVdzmF8Anc
CPYpN3AcgaRKHFmd0V1LDvmbZtNsiLiguwOmS34tVKS1bSiR4KhJWkxrfBFFB7Tu
IAJ7Rzp2YAUHZCw6T3DKDughNfA9Bc+k3j6/wL9Ud390+FuOctOeC3CqxvfOPmpN
7SRIy29mpojTCPXDkyam7I8T9CUfBSLAH7dzMH5OcQUlqeYdBI5qtOCHBjYy/FFC
b2Ut+ZbTdZP02a14FgwsGjovtUsYQfsV34FQA6FqBjobEt1HaP7JfmmOm7Cn1kYg
9DvaOJASm51os5FfcHlNKZ0jStJ3e1gRb+RAupK3rsvUu2J4l3eNDmh7G/15HQkL
Ag5hZPQhxWniGDjznXylUrhxCEfXt0N0uqDdowzj/r+WPVhNJxoVjIqMjXcl9rO/
U6H5JZ7PpYmDPyFMQA2HEADpnZ78Bbtugu8sFojlQl36Tl9J6zyxdeslNTajXeRm
VQEQrzWlR8s7TT6hHgIySV1USJ+Z4i4CKAO3Vi4TXzqQ2V1lwYc4qiHYBLCQVA0C
fCaTMEudXp/EzPvqfp6gE8JXw2rK4xMQrtvebq9JsXwlQGaVWRmwD/Rz8wQuassV
yR1IY5aRoLTG6UmHOXHxYPK0jLeGicb0xyGMYJJ3OTWSwuDQCetLCSCPXLtTtq62
peuKUi0HGf0OyyCZXQnOi6yMs+W9l+Scw9skcs2zee09smjnTheq6ifYo5yZCJVs
MxOlKmzXi+AzMpEwBfKmuqPcfhXs+kq5Qx1cMrXcsU9oaw0jlFCF9sz6jkbjBscs
m+m+wbn4d/Wn+DTOdYxsVIqhDA9dDJKDlY5FwUDs/iAQSm+mxg9cQhKzkix2KCMC
4yTLjjzZ+fSOA8rAJSPNgA8N0Q4orq3k8gVzlfjHIq7jH0TynFHEgLKTdbR8DU/I
qUIZKYbOf+3N6KyZonThaYiq7/r2DjisWTKpg4hZc9BaJSal+I9UOHRXPPcGLXV9
zfKyFOSAnp6XhohvFUENlczZIrgOlJKYIzOGuaNc3Y21GYtRZzHyPTvPVn+bpNlf
ivanlUrALtSm44tFKlSOoWoyrr6PyBwMb3hbDmPrX1JsFk7mp1arOHHeKWMGIWMr
4JniVDi6jaL3xeBRMVUbwu4cVzNDpQvjPymK6vIeiZEuPkBFW4Yc/REgnK8T9maX
KlDSlgd864paaetCXfpkvps0lFcVSDaO9B7YHJlc6N3Fg0lY9bYF6hbJBE40ftCi
/MmogIO776N+Wu7aErt5Eywirmpznvk1oScYqBMALY8kUqrfDYCRPGXaIyCKjB8n
4Y8XMuAv7gqQ4YRN9c9Xr66TWRaZfCyYdCHcRV14AkUHYMDTyiKGqzg18afJ2zl3
qEiuJeonQ6c+LoId+rq9Dn21GXNiyg4SjiWeF7nlsLS7/tvBtrWFu9qhEiKeWf2P
DDX9Fw93VZlYuB9v5tLDXgdmIQBl7sGrYV/X9PntpzXH4PB3C19sxJqMkTm9UTiW
ngBhZ5fATXcENojJa2GVKTPn5nQSgV9A1HbFFrcvLPBi0seORW9b1OLTaGZi/qcy
JSGBqY4FP2JsWtbhDH2x9hmLfdEvsu65XUBg8lez3luxIWqcGqiOAGrf5CSao2j2
PAWLqj7YkjUP7k0owQIVqd0QZL6APpOdtOcRu4gYz0rjp5MH3P6s1B+8A8YSFVbv
XujrpZmRq19cHBQefklcfJXivW/9TWX3BSMESeOS48YyIyvtLVH+IAnovdahHbHG
fRqom9sbJyF2+0lrg+pVVSeVANGAF3CVAPVh5JUlVWGkatwsKZH8WY35ZIxpfwaG
8KzYPeqOz4R/+dpXd1EB+7E450T3/nccaPW864AuMpX8Dv/MGnIO/U+L+g4w2v9o
xjH2OB0pJi+Z8H/xgwB9fZ5uRmaHcx7r4YUWfkNqNVsv02UrIgQjTRuZWtZaai4h
gqD95LMhEpzDOCKwKWJTnArv91vFpBqMwddBe7Ad0iD+yjP5gZtV4ht9z4MrD8qb
RJNbXhbnSUs0VgNt7uNppz/aV4FkLxBxGeELb4WtkUFhoN7Hk/IoF03j2Uv6hudr
ZeLh7k3l4v+77dDTYvnK+s5rQ2A20mwQCq3pqb2RaEnTWYG5TG8XxH1M3YWvECzp
WBDEz8XcQ8jiVMp1UC5i6+MCcPKRY+gE+ATUHypTt/rlJLf2LFoe3+Ob7ye3zCrn
rwu6vit9BNvDLDwJd/G/6Rcxgowe5dLBk+k9OdgKOCx2azVTmbvBunEE/gnmRni4
YGITBBK89YvhpOKaIWRk1l611wUWZzQ7ov5MllXj4jSMxzSgbXhkVuMiAys2Aasd
rkHVA//QlnEBksOg/EF0cyJXbklHFlj2mD00YiHW2fM1AgaOyfiG9xqBHu/qkL+b
YAVXre/qykeOMqUwof7fcQqXwepqrO3XojGqjmeE3dpT74VrhfHy/2bU06Mlv0vS
h8QFoKeivVPZTRM3wqwHmVQ1J2J+gvwOcXN9JFWygYUCfjPFg1eEaW4CR42UCbfx
6JmZGx+7UlRiy38fqHqV5fF7EgWCvmiMxfJUeulKBe4HHwhQwEFNXy/yno9Dydtc
C9dCZmB+g3jklX3Ohz3y3P0hDOnTTG57MxKixnfqOfehZsiJ2rGyanTRa1btzZMZ
AxsocXICFec9tI+1hx3Cet+npqEwyT3eb3WjW1CmoVptEyVTKjEsmHgW1/puvbXO
k/MZAu/ZMSHuh6XQwxJvDBPLLnuTBrXUNr+luc9T0Kn2Ghp2w+2zuAlC3u4CbceI
Nir5zkwt+D05rLCsTKvmjnNjSMDz8tBd0nMqIGVUww/ygeTUp/uJnXy6XP34/xj2
Mtr+NP/vTQCsMy4G5sB78NL2/ZkcDH2sZ5VFo1Cgd2IdyITnFAp3/kyWJxhMqdKY
BnthSVuXSMNzCQ+a0h0yafj1X6QuBGyuA+uFXhI4u0IssVx7oyolSl6dVQXjJNYN
lNuYZoeUoqZOznSDElXmIplGfIkkz+IFgxeUOg9F0dhZWIM4BCxeSs1Sozjpg4QF
Fg52YIlvp8PG+3uUQkomdkcKfOIADzE5q8w7Jg02w5Cab5ctwVe9IRZiEpiJL6m9
qys5FmwBZeK5J6P170200pCmDffb3UlsPnWcxiaNLr8G8023j6q/lxmMawBpK/2M
W35+BZzsJHD5QMV1GwepSt5SF0RjDEl/6EeMOM5y51R2pAL6mtwTe+tl4Tw/7UH2
Fu08nDQ6MlBpQ4uZv0Vq5HLXLE+t7cRCT4mj+GW8EBqpjhCz6LEsJxrC1qv5KxWx
7gtHKc9n2RHRfUB5zs1fj8XWct8Xo3vKrsKX3zP3kxDxcsJPyASvdFRzswUAslEd
CdSJgQVoX+LY++tAaRsQUsjuQQsXsiMREaBj7iigd1PNWrDUmLan5xjoXjmYD9Bv
p7exmXhcjGOATp8Ih5jXnI/bEhSG+BGv0t4yhG/HxiieK2VptGp7hniSqBLRkESq
bYq2+Y2cIRRVdF+nsQcbncdvRcdqO2UoesUOlztfIQXjNvHhGnI6sdE7GBThvMWc
l4Cy+MY8AEh/mLM1YwJDVIysDka3zvZ2+rLx2RztoKQK2ZCYypXdWoPFAGs9UzBG
0bUH+hgKXCzE+mVkdSP1kM9abGq+FO89OCl/WpfNLzXSxSiNztsUsrpjVQ9A3hwH
sX32IDANIvoAqgQ9TTKlfdzQ9ynlx0pFDupob/e++tiAf7R2+r9t0s4ko8M1IdAH
KpMO2bTf65thG29ZsCPKH+OksOBV1917vNyW89tbSpGGNAH2mbjIMwNYDhcRfER8
QxCwQxiG8MoJXNTogoAlpyarrpnHf7DsOgC9LZqvRqYuKiv0Ut24kHYYGkxoTnt9
TKImqNXG+T3YGFq1wfZyz2QgT1ico0xDH21wvVM+wz9KIO0qirbxkS8nnLPb+KUM
yq5d2nT1kUDAR+AyIWhS9IqGoogPlnf4NuQ+5fL8r2x7t6IbwlsQ+Sj9IzuOTaCz
qGTbQxmFqIhIb/0SWG5D056XJDK7XEsGT/z+LoO7pvB6InXmYvEceRKoPj7Ix6HP
`protect END_PROTECTED
