`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DA6K75jHR9z9KhEsOJJfti5EgOjZfV8SX6H5dbqlbRbwGK1gZrpumLlOuM2/FFFa
HOAxrQVq1m42+LR0ljTtQwi3hT0RcSJSYXd904F75PU3XTYGqLclqBB+dRAni7M0
r9ajB/7o4swcyFi3VXaXSqmXyO7i9OfodY9qL3F2WtU0StFEbaNJludAYmglwyCk
1llLxWL5khk9YY3+e+72M+OA5s1ayrqdRLKkCdyUsI1G9NyDddkOEDeXVH9AEwX5
rcG5/O+ZSVEDkXyF4GxLx3wM2aNL8bbAdL4puUjhVWPGxQCRW7RROTwFeosNrcNf
p/xpTENr+xRWDiEvn9sIMZ8l9XhgGp6dvockfZGZ+2QFeYmc1q4BlYDd31q3yZyT
n7f1iQEBLohmfB4NusB4N8uuA31SvJe4hdCbBFBGvHDjXn7y8SYaLEXfj+zmmJpz
0AJfmjNw4/AF+oyLQDAXWDfQwrNAD1/jMiBXV1c2Hk8hviFCyVL/oS+k0pFKH+XW
U01L+5QiKVG61MnPZA/Z3BIjrd4jGD1vsVIo1ry+JC0SbTza93NPBGJc0tMiLF5T
HCTy28E/S2bpm6wGofbyw0EA3kf3Zkcre5FJ9WRvD87O23rWJIkcGv3yEvv85/Qd
ACTXKu/YxTC+TlkHItNjXSXioOgxk811X+hybc4ejNp3IOrQrpNK68fxisZG91jD
zz46ZsLcgmuko5BrkiaPYl8p37t0NEtfp0nPog7tklLwObq0RtFYfS55uJYuUZR5
NB40MGvlKKr/rJzWQvro1dXsqtDNKHE0gPIywkPoDIoUFoHdUb4xavwjjMT/81Fk
VyFCIFIRXZq//REuZVZ9BjxbgmAjC7CAfqPJXblylp2mTIvHKYkuaHh71c3Xfksz
`protect END_PROTECTED
