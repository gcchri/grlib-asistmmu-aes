`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XQ9zJC+ENPJUOKo78Fae/C896ZKZtiFI59Gb527TQMsbhuWZ/xc65e7uG8w/2cPS
90hiryaCbgSgsrgoUzxnOwnzwLzR49OXitKx6hqYPd8UZMPjWoOdv6FRY/14RQ73
oGYV5YMDJ2yz0lZS3rcQNuFX4VyMzudVur2Db8Rn5c0h25CsVpBfVqlfIz7LhwEi
Meu5GV0eS9vDze8yKWFT0wq9nWeJEIdre/qi4GVWROqoT93bGnhg/rzScdeuY1QP
Kp/mz2qb+8NybV6+1uaNH9mLYtsum23um8STvL2lMixIr3nr5zaYBnzu+7b7dkye
jr0vTvVtTugMRlcVWTyLfv2Cx2NFjLRO4y2Voe2IJK9qJWyUmI/Y/swECNHe5nUd
KJg5P+g0JvyQVfnHO5+iG6w/N0bLFVP3tpecsrdgeBk=
`protect END_PROTECTED
