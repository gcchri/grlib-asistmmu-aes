`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pF5CyMdsjo4wX61n7DI3NSwz2MXKInCGMIUON39c0/qTzKLmNdV75+dXkansC+sJ
oN8SdckwA8SmdSyG0oFW1kpShIv3nPbdQEE4RdfJNZdcyRe7hplwuEBkGRJbRl64
7fh0Ev4TSvuKTuAnt6JWz1d8oP0ZgVEZICkipMOsFXDkp6tcT+5LknZ3etJtX2lf
ajR95Knoz3a8Rcp3BvDjPIyWwqSzawgeEZkqxzohBaObzHpBKaG7bbwV+kvxKAOg
AD657lCCERk0zK6vJebXeN7oqxxJ97Zh/H02KuiBk79qMoplAgglQnNTMGbFVdF4
RDShBosnyqtQh6sNHTcnezmS5IZ13ApoDSWkApFwtuLC2cOX8UOFRxwrh9fFDOGZ
jjJvgk/0kgZhnfEElhz6U6d5PVkAw2EfbaIWaSvdS14VpRg/VMYLH0IaLI77ddqy
BVZAZ3uy6OepP+KfWBgtuYx6TzkSXEvkpS87jMPH24Kt9fab7R0KbPlaZCVBAkRg
JfZJzkgMe79QTNZC9FEYrCUhKnzZri7XL4kGYXr40jU2VQebiqp88fpbQcsubEWp
MyKpxYqOdpW75x+fJeZqrIOEpEtdSLlpNGxa7d4MEhJ5ap0/V8amr6zr6RMSUNa+
VkYU0nre3yFsk4K/COdYFxGAwdBieX3auVqqbUu08f+WQ9Zq9dtzdQZRG1QsSJVi
HjlPRl3xo9XZ07rPaTm5JX8c8/3g74ZkUdrgYBVeNYOlygEzm5KgOhBihNtKIcTl
ItLnI8CgRIFs+7c1JcQ85BaSZzIBPJzo4g0n+CTa6wopLW0aVGdtiLNQsRENYggN
EagItPudt8DG88QlpCSEmh4tXDYuy+dXE/3fV4xqPso2BTh2uIZ0SJIvfqWMHGoC
NkuwrXDbJwk9VKu+TRQkHQhn1eQlJ6KckISh9EkwD+Iv+no90uMEmTgSbWdJwEZU
A2UKRFjnjavlXGR3/Q0LdkAMiphPn/gYpMEWgxJcFuXBSJeZRz4ZX8ohXNq1kbMw
ug8sDzYKc32YKiqWiyhm7N0ul3B5ciJUMCwWli/KJYh6cCQeISBWVlUyTT4fq/yk
cCi10YTqYIp+OuyXo/Xdb3lQemt/TxRmFq4erJanXq0x9p9oSGOcGrJWiIwQsT4u
kX6jgxNS2QUuhIXm+m3R3GFDVdTCTsmuaaLwm61BC+X+xpGJvN2bmoFnFO4ou9Re
Mxps0dLPyQZ0YFWpQWXOVcOqIkRZl2bS9Am7h2EPfXVbOSlEFSYLmYhtNVjrxD7H
taqfCKE0Zb1XuqNpmTg7oMRokwGXcwkSkiI2eqju4HL7qTMF25B78hdHmAXA5Msj
Zry0kR0ojGwgkqxeLmykM5VYTF+JfHUkasjC0PntDr95QuShNhEgaynZfVnaoqU3
FePzmGX/BN+3sriBNhvyz2dv9IwSIc1F3WBM8AJDXB+ODtC8JzqbsPG3S2woRR6h
q30BPVrDHc84faYWEeePqnSs1Zm4+w+cHVxJz7rnbgD6z6E8yY0MSEpaMTuRJSDb
cn2z+niZ/GqozgXV5suhVR+qwFM/YzOeOS1Z0/LSKYkTwaWztO2bIS5iE/RgnG0C
9R0Ly5MLxO2IB8//vMlFjCkYg/mKRFFGslwn+/Sx9MLvjR0uWNRl50pqw5V9w9+U
uElPKJsm14PTBdbNvBpbZVtNsmkjye+QWIEfiDVaMYm/XfkdE/rKG/VKbX1NgLHY
Nj49chzVLJjj8hcf9L3Uoj88Dc+L+9e7w/rd8tvTYj5Fxn4LcBPmoF64sLaZmCfW
4EByxUQhcD9hokRip+2WsgOuuy9kQ+wmwz+UT5lxxkUPzGZnGyvLTGsvjD1BHXIH
Cx5tLh/pzn+T51wJAqmRgw==
`protect END_PROTECTED
