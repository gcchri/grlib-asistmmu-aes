`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
obmlQbnRtHDazi82kDbChCDkrltzlOIy5c9B1OmMTZ/wWXhdxkxtLnvBrOj8W20K
qJcebWcV0I3eWwTF5a593DIPZTLHq5PmizRdPvl8ryBsrx0bk/b7RNjV3J+BP2Ch
Gnd5uM16ZiOPwHOrnCKDgIy2dTk1JYB1YYT5q9Pe0k3hO+I0aYa/ZPkguBBn5IwQ
KxisYeNAFAVx8sYll3dgFvFak2BpkUqvrQMJc8vFoiV+UNhqfNfNuOqR3abQeqmS
WygtYWohOY7dSbiXS6KzMtXSPL5rbYCPWMbZDSHDb8p47B9hFufDH/radpGk51ZV
`protect END_PROTECTED
