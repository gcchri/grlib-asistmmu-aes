`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lcVR6eU6w8cOpEY7vJHbEpLzs2cGPDuh5N6rKzbqKHiaH4whdCxMWcy5MGRCXff8
cSsGQEWVr4XdP/FMcDfGDD1LG5Rm9wYnTWUSHibyx2OkNHuaCTj5NnuDTKkp6YFl
EydkB44jKDdAbyFzsWzRrXZXxbfOQ2V31j5rIfsnj351wBXPKDibdF/XSg0uNZUA
cN/DF7OTFBvPcMd99qqH3Y15VCjCn/UNC15o7xTPDDMlryguYZ++92z/TeU/7j4U
j12s2e/MxIKNYMsUVzcP270Yzo7UkDu5LCUs/t4a6Klg2SucOENB104KpyMupQrb
DzVJpws+N2OJxL+G5DklYIQ//+rZ+qs8/q6gv9Y+y393nIMWjcJHuteqiMi0MFod
IaWrP7tIJ7WrJhbqUQcUJtBBO09Majc8cI+BWMtpg3kNGNbmg02RWV35+r8DSMKI
jWuq3Ck6IxsL2IKfKx9o3KCcYNdMJFNFTYb6b5Yasjc=
`protect END_PROTECTED
