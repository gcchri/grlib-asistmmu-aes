`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pwGG9Se12KLgbTy9FQE8XyjHQT/jXbARjYbVQM+BPqUaAO4XNAsVvYiHA5uxWLba
ZXiFHEA3HctJvnxBzKCJurFzOTrpaBqoMeaK9oLgPQ5ggKQYDuuGIyGWmlIJZ8vc
IZaEVhQ6NlBrjVHfgGXTTgWRNt1SHHbLOfYS3i/t4dgrUJ2hinfG4Dr/Hyqtc5l4
ffsBcMmvAeUeGFw+ZiXuBlG2owIFVLt5pirA0s6JdJvOKiUx6z/ANt1VUCP0gXbE
a9ouLksDc9FMEsduZthLj+X7C6EFY4UKxQroYy6DZdIm7ErVp5TFK7K+qjvAiidL
F4yeA3tPM0yWQHtV1PQFtmS0nxu7/kPQNp5VBDx4aZQuZD6Vaq6VVvHU10XBgVCu
AJAgU55bfpa6UHaLbUMt8Zd0AohWV8fU7n+aCnHuViaMRPn/tRxg5RxyeN2Zqugy
4f+UjU6uO28Vf5wuh9o8WW+PxVJUcUVbwTfoaokd6Me+7vijq9vDWrKw0vHtCrQo
z3q0E2qeaCR1bhT77C6MItsOsUq4OmovTSQtUlWuheOab9MsOrRLff8EQaTMEcYb
u6I5Up9vvzly3AcAT2cWXtX1MHKMUkjGvVg8CtsflDEavh9eQ+FOIVOuVBIcaCOj
hEU0D95ycmyqkAolhPt8Zg1O6eUkH1S6hQ8Ml1Ngxeof3y861Jts5jCocTwgm6AA
`protect END_PROTECTED
