`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SSM7ZOPOLuwH00r8PfyAYIsAQQXT8BC/JG2UWSwa8625M755O29Pwb8HWw5oA5zc
5lASL7Zj2Gj7Ds2Wb9OqHQYroKOQRXGTgXpTO/JIyRcVBa1YVVZiAOH58uJyGp4q
bWbtbEJcribchzJR2YxzlLVZnnsfcbXuNPyXHUaHu1lYzwRd6FFHXEdkJTuCgcVu
7k5a28j1VJ1PHcvgC/vk6uwgqSqDxw0FZAZVJmWJzOBL9xteZQEB6MBKCqy+gKxO
fOs/QZdOMWDCzG/juU1yAr0f0UIvTzG1CAwcHMi/BTRp7wbJiJ0hu8bFqJjc4BKs
rSdzaTFbfvbYdjxhhKGvUlNwLwfOMHd61+TFAVR85HAkpaZH4/Jl6hdyyA7usYZv
/MRFKqWrBiNqqqSK8QoSRlMptXf6+LwBWAmqxR2/CRlAU7Oe+XYanP2JKE6qh4mF
`protect END_PROTECTED
