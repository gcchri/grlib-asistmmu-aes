`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+GP/EVXeg2ff8c4GGXIeSCjIFe4DC50pFdcxUgqSH/uG7ni4HJtkZPqjntIgBO4a
+eo1FuUYjQXx+1YH0XoA2UG7axilz90IGkSYN8fcH4FL2gUoY9VMHGL6tKDPJVcr
bVELd7TpZkOdMXxoFyDAWxubYzDVva/NY5gTWUrjCw2GNXNf3l91aW3RYcwexX7L
8GPkK/tOaLGkCHIKoLSdBuj5IDOA9kVJrwib0SnXA9NTvOnJIiZrCPkYfiApD7ZS
ozmG+ONoFp+FA2yyi8/anVAWhcPemZ+q4UfetcVQqIwv3K769FXnyb3tGao92mh/
NM1xOd8AR3Og8jphGgSkRkjbOrD42U5FIjaRXeb5+VPwrSDH85LgPV+mek0bunsY
Xz1/oRz6IzdnbsxFvLx7jeIyPRX3kL6dFWOopeWwpNMkwJWXQcD99HHCI26ySh2h
GlJB6Rfa/kqvJVr9SMZVIwg1sCeiBqkecyq6td9k9QI=
`protect END_PROTECTED
