`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7PG7ao8166iZCd8Hk+mq0GWHbboSuiFk0aVXom/U+4bhMAwkiaOKy/S3J/agU9ip
Lif1Zg4uDHYmYofAp2y9pMeolh4r4RdK4urp0CHKPxTe1nWQ8wKZikqO5gRhR8bt
E3MKMRcTeD6v8Yhjg+5egGg65yg5YIhXWjOIT70kniaZVygWT2TZ9QvGo7Gf/9nu
c8F4tECuRa6J9Lg+80uL9XFoPL8fGC9+PMQPxL0szDVbjoC2rpdW8ZGf0h+jIPei
ODL2xDOuEnx0qYMWS4dL8IPPnIDEQ8+ioPR8u/rHQ0MBzC1Yv9bkofj16lQ03FF+
YRpXShD2JoISaTLDcyrfOMG0UeyCGHamhiu5Odu6DARWkR1/Nkb/De6OFswVwSw1
ERHhWcBsY7i+58zdcOU2OO3KdNEkvq1djofDr3wfQWU=
`protect END_PROTECTED
