`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W6Mzyx3Tiif7be9dvSxe//k7qf9TKKtV+6l6lrOPbewYIE9Wn5LlI06jCu6nE07u
gBbQm1JSO4zvbdSr1WiwUnwFFVklBOcSBURt0tYQ8OK9kjbwPyZmFFt7QTytvAbI
jsd7GmjhQNFbFEWho34u4VAXNrdFZfUDiUQlOJKabD79bVnP0jBeNwFs4mtMg/GV
KMsO+7ZccWIuPqNIJF4Wcebh9TSjLxshY7zxzgkuW/VgfjNkvZyjoJmTLS2zD1QP
wrSy4ChLPNua2VvR9plqqI1VwdTLHqOfm/+VaOdTBdCN9xmpDpths5ct/EbYIKMs
66y/tWJEJpx5UEuaE4TRFMvw2pmX4e//ldeioIk2JmuS0V+WAHD1A8aN1hNxtZ2h
NRcvaSoSFU/6+OEDvH0OGisdtUFfXPvapRZbWqcK0j0J4tamg3Mm2AQYLDf+FTtK
5LZoCiV+r4zADmo8/1l3NXx4PKrf6DD0ANdqXXeWqSPOpSUxMPY2DmLNLSj2cH86
TKMoiXI5/pcnQZ7pTdB2PQG12TK11pGo+gZPsEEkGub9cozZinsJC0PQSzpdl5l2
zYDcRtCim4mRJ3s/FFY8hQ==
`protect END_PROTECTED
