`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
md3LEzSxD5EzmAHWIktYnI+05SIIOMy/jImBJB32iHl37GxfeF6d6ZKX0Z0ozqQh
7lk/xqmhla0AP+P+6HvyAPKXPd9b2gGYuwrYZhbCN/YnNKFm45TrfOmkQCwuT0Su
MyI7chatoQjereqpme7+D3pZYpP2Mh1GFGQSV0CDkxDbzUbn/oHO5WANRDKOaCUP
7aA7FT69mK7D2kZf9D9RDKji8zF7zPmB8jQmyXwmGIBNXNHx8vhkt9m4WbNJgRyX
6hpqLHawzbnykFOH5nIMJ9niJ7NZth54jntrSAvnftJutmkAgu6ntjY0z+3OjWeV
S0X6wJlpVi8Zw7VrKOoWkpuPI6zpKOXVn/YHuTUeQ7x42QeCaOnzZLMYmKDhh7Mr
HGpKFzdTMo0F0wlFS+dre5/v5L/7/KdK0M1oFD6LJYLXs+oHbyrEbY7YyERNA+uT
Qm2WYZz9+HIbz5sOO+/XxCPhxXOqOMJv4S2vv+ic7SuKjMdWm2qfMkVS+5IFwHL+
Ve1tzmqh9URP6eAfqCDr0Ac9R+KQGNTtLb5Xi2hQkWnpBOamWEtBBON6iXY+CZnM
MMt+lux8w1iiro5zVhgCepKRfJjCQN9rXtl1YGX0MkcpUZutESzzE0ed9rR44ZYR
+wq03voGPD7GWxK41Qxf54EWs2Z1dTGssGUOIbd+tao=
`protect END_PROTECTED
