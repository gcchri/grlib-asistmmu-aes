`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t2a+gVTPOmVQ5StONvf8qDVZidBBtNAzEeabk5tf3PEXQg+iyaDJiPxrtDksvCGI
K/63Hodyp09s5k5a5lhOqDmoVbve8mIcToLi15RtJACSRTbt1+8WG96JKoDmHQea
rr6cUeVRYSSYeB9OHyIIWQtotgdyL6/XPf+kfy2AVaQ9FKNfb8hyLrIQgLbNXQnV
fBql6URtR6WmVWHbjikBjXxQPIvHuANGwimWMuprKbMnX+IjayrfSuRD6FX0xd+T
OsAWl1F3uo0mTbQ0Fr/RMpJsF4Fp6BV64SXnwnhjPAhg88N8egO/x4tgvhBEfVwj
Zaq1n8bURoiyqV7D9wF2RMS49B7nTTEW5HbySHDK56KGzX90mcS35Md6eMac3afQ
DcvsRH2+CO4bqa1U1mDUP/CoiWZFZpP3rt9WhP9AbEAK5AqwopmXVr82E4rwUQhj
WWsiYIKjHw7tDdE1qesI2BbVKV72dRqYeqFKEeL+dPbwXAY0/YajsPJ5++if0dWc
KVIUzIvezBTV0zIBhnh3ByQhBizcS/ZPUFvIHCPMtP3sXjak4zNh16jfp4+LwVly
Y1NsGpWAtokJYNrbNohlYdJlsOWX5mlaRbh3syQNIEGgiL5ZRzD+fIwWjTYfjnJr
J/FhhZxh+vlfr0p7itNv9A==
`protect END_PROTECTED
