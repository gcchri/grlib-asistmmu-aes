`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C1jP0hJgBxfxlH7xh6yQvmS2Qj9UYEUZafHGviJpUWkmw4X3sSSCTW14zJL+a+9k
NuhY88P7nWMP84RuzjLX/Vu8RQpwXfXQGyvi9vMie2KFam+HS4ZAhWOxzZb2D/uy
7JIcoNW+K/ibOtWDb3pxpjFn6yLm4TEHKNNZb1vlAu3+tG7ahUpWeREMnSGUFsRo
gh8wn9MV020eNRrEgvtpt6yfanCzXRzBbUE8blZcC8GYE7AIfdR6rbCDkvGYfqmZ
a6BPkYUiH63IfADCtsiRuuiqQ0RVUkqW0FcfzwH6j4k=
`protect END_PROTECTED
