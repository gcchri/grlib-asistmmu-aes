`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wB5CkYkKipQ1Pu2zGKowj00gPgvG0Ezaxx9WHA3DizmW5fxe7hLfxyKxy3UtWYek
o1O+RI82xaHsRex1NcX485zqLo4wQ5Mkk8D5xKRY/X0UlX6MDNB0OHFmpnZWwU+B
6H73bXOEoAJJaRah2J+c8CSSYWucMfjRIBjcB8ByzHnhGeiBULXENTTVRiNpeCSW
cmyEhrucLvXQ4NsoSGvcEVRBfIlBvJm9bNEhUZp00nVTqm1Ck3kaafjcPqYImDAj
C2/t78tJo7MGGliLAWL1JHa7lh8l6z1yrT3aqTbF6wYxfW3dkmAFVq9znb5k4sxH
r27qd9TKyIxgVA1x3Eju1XWjShMxqka6yG4fObnAosYBWg53lNTTrD1D+KtyV/j5
9zcug4Ax/MMctlPSY6r3CsvXHbHsOHer4kdn6i1ZKNZN0NUY/4yhrXBAByoks2NC
3uSIQ4WhYR5eLOUdgPYEVLu2/EBQHBrszG6eXW9nJKUzj/6YFNw86k7OCUg49XVz
8KSKxV7QBmQRyrlmjOBia4Vq7QPBQCaeP4tGrilSwP+OTOEs1nDaqCdAnWBwqjWB
lr4Jx88jSPc93WhdZ2FDRRDEAqk7y8zW42exGKnPTtg=
`protect END_PROTECTED
