`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ftS1Srqbpu9OcDFUOY8YXBYmlf5tTP/WxL65+C191bzUyK2OFQ9LaC+Zf0sdxPKf
bnbyAEiOiT5HTGHmWxGDJC66CC9hXKVj+hC59JEqjBZZslLwFZgmX1a59GeCfYZK
xmbcrwMm6SJ1hzOi6wGP/5veI9VNTUYVGaP4ZKvHKKwWmPjiUYQpAe3R9oydxVYs
SDvJIQMfetzR2djPuW9JDPIwV4stA9J3WDj8+b7caRnEd9TqPWiRThI9cG6XgCPK
N0RxTwWkJLL45uLQDHjJdM/p3nP9g0HG6oS2QtgWoDHOw7/UcGLCeaMlXLy4hEqw
LF0cacp7bmgM7DCFXZDPvGsgFDe3RVJBzi6td1fyMZe0AUaysx8c+ho5vDhDXyvm
6dE76axJpNjdrdaLVxRC9Fr8PEGjyjcr98tCfeTkr0fZS5IrPi0ANcHvJbd/YKRG
PWlQql7PNT2Imqm5xH/C0ShxQYTeFjmw9JZAtqffIv9ifsYhk4Owi3JBs5ROorN5
6xqwUPtvhryRQinjhWQbQvg8SgKB71ZsRDpW5cDBvuk=
`protect END_PROTECTED
