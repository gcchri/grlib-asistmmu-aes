`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oxO03azNC9mDC5TjFvOBSi/X+oxZo09G/JVzYgT2GVOmqfl6QrrSg5jON1HA0zxD
YiK4woKuRWVUYH5SGw3iyXX98r/WroIromFmT3DHQzs0beM/3FINNvXoRy7Z9yOv
V0AL3aBbyW8XvKtL/kRYsztVhdw0hweiu541YCawC1N+pLv6eIqdRhpa/ei3juHU
E6pMRDFCtiioXcPjikcZMPD8RB1EUQDJJDVwP8zIsy4Nmlex+gkt0vBiSaheHZsj
u8CtPLGj/iyP9atUjHR4Sw==
`protect END_PROTECTED
