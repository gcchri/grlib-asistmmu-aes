`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XEC4jxv16kk9QBV7/n9Np1WYftSlOrl8Adg0J+fFI6UqU/Iln18h7zwBWdpnFQ+k
VaqZbA//ehHpmpDTNDnXc6uC3qDk+xDQOm3lO+ee2/N/BsWsQ9aFTHavXOxyCHpS
Wq79JMUwLvH9ajnsE4WJeekJErg7J+y9Yf6MTcQmXBC5aStHq+8EL1DkVHbEvhdP
cDWKhyJwn7gyLVvyGkg1WEb0r0+52xr1FAC3gbz6Y55go61pYdS4A8DYWmcBldtF
ti0fr7hYqBs6PALauZKlSNUvt6vso0aApdYiTheJU3hjPqC2TdhV2n9fVJwfMxZS
gYgJZk8GAVP1QDNS7AdCClbM3bJYC2Ifa7zLew2on3ftob+1J3ybKOzDlAVLg3xE
Thaw9TLu0LmkjMyWMVJuq2yXQ2P7aWkNjQzlV2D/xEDK4VemIRQ3EUJ8y6FORcW0
nNCSag4tDv3u/lkPB/17V4zFphZitroXj358Mz68/zXFD1wJzy5kSYtLLAI7aqv1
/m/B2aYxjxwQAZtY9Xpm0yH4OnNetVsx/irjDpZ600kVZLcRIImd1jF9loMmQgsC
B6V0ZUXwao1UVmOHRnWpF/ZBrQKCkfn8KzwgtTVmWzkQ3KAWOUtwq2dNH+su1Nd9
LxH3l3KHrURuZ1gfu75pgtC31qhqUa0U7gc6OVTwOXSuUM9s2vgJTLgtIMFNBvcx
Ydlmscy7AGJOZz+Un+j2l55YBiR9L9S1NnJqwWkICsUjur6cWmos+jaULfHBb6cU
tY933aX0BBDL8IeCYe1PrkXdKOW1w+8Qj9pRubYS//HuVwseJmmnJ8oQxAJwHuh7
qU/4JBMrgfBgyua4eo9KgaGAERse63IApIiozrx+jF+JbS+Y158zk/jhNkmTsnYp
8vLbOlklPSbvyQTfCUmomCp/FLNDgFhuA1JajPIwVWs9dPi0TGk8amlYDtgSCxCX
oDSfOsN+wRJwluUjzISlBmutwTf5K+QRN381+6yIVWtxcwsSduy71UimeWUprRdJ
78EOJJXSo5P87cVrID05CL+PtaXcIe3hL4zQqKj9OyM03rUhru4uJqdS6Hf0YPbK
zAbVMyhNxbcI0iAEHDF3uhCG5VL9K9yDR1lDjNVIxFCVS1Xtbvl1Zg82+g3J2uiV
V+anAPezFENEJ6FgOIZ9NoMKDWZTqrn0i4Eg3e5PLx+F1NN37VdpwUJkK9oiyF9d
pF8otrXS8UOm7CQwd4Cll6mKhTrozVxZyvJML45jKwK5y517MQHRxEEJ+00Ygag5
rWBRqVhCLTGNIdoL8InyyBrD0SNjO4mijt8muS6Ntf9D2Huh8hdfIG0IZwzoKxzV
eiZQsUypgy/eBVXfjoF6TIHHWVxMEZivsFTpvyjA01FDc14VLup1Nqp2pVoGFU6s
Bq4PKLgcsAE7Au3bsA6qYxhsDT50lSyAYDS5nq8GX4KaJIGmnCDy4ALzSMgHv8f+
MpRVMZ2BoeHgV+eudbtBfcgLgVtBRl1F9MkGR19z/deHwqt9CJ9CqRjGYIfjhuoB
`protect END_PROTECTED
