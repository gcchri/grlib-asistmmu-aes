`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D4hoTXqpTAgLiCzdN18R4LtLGIn4ufpY1u/hH4MMrX9gKk9aYcwabSfnYSaT2zaK
nV+GBVv+l2/yntMX9L+ixhdw7encqJJDmFWlnLUVE0GkNVeL1Ykb+CPX0i38w2Sj
W2OgIzfpxUkoGrCwAxvaudhAoLpI+B4gqglu3IdUccSzZfxMBnhHKa85KH6MxTJX
WY9FeC8eYNIHr8Hs1SsCa4eQ+7drI7XtoHrtkhFoUFbv7A7H4oOsV59TSN/AmOPw
nirrqHet5+qVy+exsoYXNe9P1X8/173oxtB/5NnqrLFFLor+OZeII2KSQJCFLaTv
4pffUlR9IjdathLYSfEbP/ZBCr3tWWNYl1AT3izUjmGfoMP93hipsHyNiZrYMtT9
`protect END_PROTECTED
