`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IUesTlIrIhuys7w02UjQc2mLUN73pUAAWM7Oj021hExG8SjUy1JHdF0A8eD+D9aV
tGWVHsz3GBuLY8mrQ4dHINNdH2y71q9Fminz6JpadPRXl70N/HiGADI4zQN2bkpZ
84O0ypcC1Dy99VAOxIh62nOasKYwFUCsE2iYjtzm+RtSSSd6AUHAvb+59CDzYRx+
QWUJXJpVhoMyLmMgN9xqMDGPl3VfqDR0RMsNwrTIgv0gSWCmvIMXwfVKK5byxmbq
YwcD+EJU4WUfirFpFSRdmp8LeU2p8oNr1OYVLLsVYzKhO2Dpgunw3N9g0NMvSSld
gm3oCc2ft3EozKde1InaVV+1Si/UFDvx04WZckslsejfpLla+QBg9PSCY/yWfAJo
ONkiTxqCNpen8CpPA5mkBK3jlBQJo35+iAyFxdAeUb3dk/Ag2kVxZFsc51VV2/Cm
VQMbu5AKoMp0dNCVDoofxp8JGvCaRHvOmtcLBnMPsdGa3xNAEzmtaa7a7oEJj+Hj
`protect END_PROTECTED
