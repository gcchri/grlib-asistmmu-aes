`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cAvZSluA3n6tceLTebNAOkvi4qHggfIZ1nclvcj+9hrA8vs5IaZjuRpxRi1eesAc
441y9djUoo4gVk76aBytpb2jo738h4JQZhMbSc6eFNGeTPFrnIQzX7hS7BCK2nIo
uzrwIOYAtb7uegRuCr8lwILKrCKIhTxejpgp1PTZXsyiAd4CtTEXz/rF1wFSbBiU
YchzlL5f7qehr1P/amm6g1RY86n9p//qdeoVWTrSPelKStlVpX+w09wUICLsYw3J
ntyhvVYvA+fkWDEa4EL8UOVqEVDqJvUpjuuwGwrs8VcBsq+8i00tgPJpppPbszO3
C4hzFWmz/A9aRgO4vaH39zlLSRYoF9qrG11ftPhwB61YPDxnG0YT5JpaLPVlW4ca
DVoYEV3kkv8YHm+B9cL5a9Xt6HVHt28DhPUxgj2j5UbeL3TTrLBl0upRJqicEffJ
FYC9e6BNWYqzbMpRGy1T99C28pYRpGZgEo57SVvQRdTND868HbyjoxgYbAqB2gOc
/D1h8aavIycoqaGOMeQdFJ2N5MogCPez76He4JljG5h4H/V8HulzdMr0uJMBtEDA
cWCp3jRyVJPRfEUOuWMJKnrik/Bu0ZCG34kCfiqo9KAG2HptJaoGZ1nj0XKFOKAQ
FP31TkPk1T+wmb/CmAh9asLle/8VAJJtKmCrLgzSU2DoqdTOqikhg5gMHTNk9dd8
AvwjiGnucNXB/z4P7iT9I9ZTe/9vKwsj5DlGcGFXwUvYngjIV4EKf8haNq5XVZyy
AmhjcplMf2AkpBm7skyc+veUxn6/zcZ8QrjvXmJDKT8DeWbGZMPc6zQVkqnbAPhH
3/h8Y2eI/38LySSEkHjPCqUZwXhEBZ2GTpRsLF28JcKilhCeD+kGV8uSS5Skqnbb
hg/7eRYUQo8AMKiq8MoIcq0tPavW90uCxawt2qdmcBJbpNJn3plYatvyPBmrCb0t
twmkRai67qCBTg5XRmUbI+dwtBp6FpVgeix17uPohL0PJfQQwxBkVEON3WwL1hiQ
a+pv3j46HUE99zsI4Jck5P+GjXUVqHHu9MgLWRfUhwflA2BnKD3KY9KzV3+pBPVH
nIogvZfMG4NV0YiFhSSJ3dT/UqVp32s5PpabFMgo4IUBbXgw2WIfS/D4zaLMv5Cc
Nb8BXWdFtRWQtgKKAH/Vmlbn9AchxVQ8jkQQaWDrmEXarWFau1vaQxOckULrhZ1t
sZyi+IlbicTTAzWkG482N8A8/4U15ecQUymkM29LzBZD2aeFYk/Lo6jtbmHwphgK
FJ2oTZ9c0xKMXNv8/ldqcnKCiyOCyCp/PbgaTLEOMlPmUptW3V+C2oenQUDhGuTg
UXW434qdrWgW+a9tWQYrud1yZdusJ2sJW/J+7YurKxJHzpYVcuvf41eWuGv9qVfI
f3A8/2HN1PjPGO3Plnc4HBJxZc1kmeTQPFd2YzLigr5UTBJg318bYVOWv+8tUw17
IC0joQYfDSNlgSGOSWy7h6KOl27v8ii8bJEJIPQjiE3lZCenRmmcNxtIilUHZ/mi
SA3ViVoErSetvNjVsvskydUJScSOC7LSaBdw5O6bSJ6iEzK+e6uO/PcH57LQ9EuQ
8japtjHaNEXpkkvSJ+wR3SWQI/iDSKJJorRSDU7Xge8i7RAam2bMN+TJM7ABWda/
XWxGbLV54uCI+BqDFXivDgoXx9KXzVV+Bx0ygPz/de4NTbc6dRN7kEZYMXzszubC
UlVWrPFDoWbF2fwBKRFEq3VmmaWkL/TMUfDWgfF9gX3+uU3oTnzlRpirC1dOk4q6
bSMvgI3E1F8BkEfnbJ8k5qgpbJRH0bkemq4wp4lxSFZmGgQlGVAyqPZvpvJTpEQo
19jgdmhpQ8OsVTZvkr/1I96Lp02sb47pu4e2D2pBppfC8EGPIf7oXGV9Xau7rEDf
3YG1DO4xFgFdHz9DPXjetPe0lMu7WPLo054PTAVO2krtUQ0n3JvrMUuwcRW2Kaym
lcHD4cgvjC2ldRUDh4jjaWoukvzaLpV/VPVUW+vg/dgxK7kOflMwQqdJJPzY87Pm
Nurz1o9g2DIe3Ee8pLfBMgwSEb121cZwiE/q/DOAm/L6ObGrCKZhrhAoKtIJMhre
JU+Cj1G2BCWCUKyEx6HJlsIHhYf71jiw288UlLitW6R3RHpLyzRP5bKoMzoJ6clC
Ml1kQ9jAOUtIdyyBOPi+hcd/a6DhV23hGT8ULBlThzxa0YLLNcaLp+HLPBxPfVjK
9/YBCoJc5pJzz9ed9E+uq8PVONveKiJuMX95yOWk8YfrWoHZ9yaH+4nezQy70hoW
7TaaLY4Sf3s9xZ7HAT3FI4Fq3u3ltsQkugVLlr1iL2G3dmCElRNcJkGjaTBXzRtI
vVTga27+eNv6BfpPDZVftsgoCTgL7TKENmyHXPsMEl1dijkS797qKIrOv7qkQJgo
ConTObcdblbuc3t2jWb0CcYAzOtF5/EPteVLJwB13VwZIXAmGKdbFpuJivliLMll
VsHbQMnEH94V1deb/x+7WXH58D4QV9UCN0EcXNjA3hkAPtJNDftTTsF6vVdDQlgM
SEDfk/2xkFLHZ35ybJkH70gtr62dBjL1fOlJiHIeq4V8kX5K8ANp7Ztm7iXFWMN0
cTMJ/6psjyhfmZdQ/Nre2FfPD1yE+3ldoTNdJ1E1n556h2Kfjoq8tcELYf5WCzv/
HzIMfp2bV0PdA/uIqGgSrTxGdaukNp1sM81ov5KRpu/SsQK0i9G8MsX22jp7tmBx
yv6gVJuzWYc1h8DxabhPlEauNM1TEZvXbtavkeAMl5ASFvCmeL2Q+Hj+xKpZV2Xy
Dg0LkARXi9UTyOIY0K2i2XahK29go6OJWLqWJ0EIk1mFpZ2k/qS/wEh5FLr5zKjk
yko+TcCDgRkXI2GnNK8NYJEk8ENcrHQqbT0PSfaMRG99dNYXvm2hyraiEXP/2Bym
X40DY2G1ZCO7oISaPx1ZF0MhIouxnsPg3hQ5UYlF8jZXiNfq0yJKzH1+0TbAGr9q
ptTyo54srcjcc9la3r9usBuPCKUy/89tByaGMR+S3/Ryb45dPh9B7OPjhpJJFi4y
33QE8XwEPjyYHBgqEEtkF9EaTwwOMXBk/ATcQ1pv7o81vOflISsmkGDSpYfJzMiG
SR5cWOQgavXCQ8a0TtnlR8JPKBaOjlSnonsuw7Och+b4Vqnv5jACSPhZOcU3+BdE
wNokzLJDYgtD5PBtPhTs+JExyBSEcxJLDcbBem1ax3v28ZpXfFCvFiYf33mhmkxA
e+PqrmMAVmhPvFUs+iyd3+V1JxpPjRCoxzApJ1nURAsLxpJOuY1y+BtHjL01NCsW
UcfAqsqXFL3kyhzExTEuQlZE6VPgN1u3oTFKWKrNInh6bdfU7Jj6O9SJrB4h0e5a
pP5AkbLLsXuc7oWASPZArgRjnRJ6ZUZO2TBNzGjkqgkFaVoNee6t0ZK/iBUUIjuc
MuiTFZj6hvoGzr/Kdh2pkQ+1vFv9FnbkQOaTOFmfJ32QMg+XGs4TztYKQwJ5IBzn
AgZXD805BLAm4IJMG+7Ay9+UquoZmpz1m97u1fPaU0Zgx/09FEAstQS8OLPfuydW
yms9b+E3H/K1fBos6e2dhPz8ACsM+bW8Mo1wemVQkMpeF++0FBDjA4G16P/FUEhY
BKsOB3zRjR+oz/vRcVA3cgHiPv0C7tZjLGWBUh+POuo5op21Jzqosxwjk1v8o/t0
ncoeOly3pCba1/gqhOtwmqyR7nD4Fxd0wemn8/SCUbe/q+3pWMui49odLLMNNlmN
1WLJYUaN9JGG3RuAhKTHQv7Cff3NtZztSedbol4Cr0mPdxNNTB37LghzlXJZ92E6
24fmsd31/k7aRF4eJ1sVQaNl5JVxFxquGXBKGmNuRnXPBQEej+vDQ4j0ISCDautx
lBRCVm3obFlhpJvPuXaCoMwSI4UHtcYIVFYACGKHjyOi0F3LVW/OJ9zblAPY0sXm
v9AxfUveulSyx8Xf9Adh/ip8wkNjrRMulYGDj9SnpTyszdpeaSNVKB/1dJBizVet
fsTQeY1BxeN4cTW+Z7HnLiYlCjvicOpuXduHHCywIO2LQKTVjQBw4jxOQkOxRNh+
cU4RnJ5FToL7PhtzX1y2ZBo0OE3QKvBAZFetzhCTeZGPvh2CXxJ/S7JLBLWJVI/r
S4LrLMA5UQBldLAKnzLQElKsOv4CZEZ0g2fcIuWoGCpfh9YAJcoedb842ITLoWhF
7QhBQQ5hlGoyoUg3v77gNxFa6qO+4lgmuPfFDlwnSo0RNAiEHviQDwMzjXfTbim5
wgxSSt17ponEIh9j7b7m5jQDVJ1jRWyOKpQLdbLBGDSKmeeoOut2xhxux6A1C2rk
SLhAvfbHfOsBgusEsWEruh81OSA5uRxDlUJib+amQveJV7rGapcKefxsgrCn3YR7
k3C5ochPrG4UVVq7u+U82Ohebr3lRSJvdh37mJHmq3U5AbzYitK/Ji4k0Qj4lhGI
XutsgRs/j91NFLUjmc35THX73iHYJzOQPoRUSuWxMmiML/6JTG0kD8r8fKO6wuHb
T1AOsRlUlw7ZpnNfs89OIyjGsSMztYZmoI+Y2ylzaQYz35h3r3Z1sZOrbnbbA/Ur
0rBKXZdeMhAHSaSxRg5PtcDtaynuNTL7LQbtw+O89zo9J54HPwJFSj6HXT4+cMsu
nZ5OzPdd4lyx6Msa5M/7H2ZC9430RaX082Vk1igCvWJGQ3JQb6qiRQ80+7KJXoxm
Pf++pYq3V+go8qnQRFeow5cHOt4WsD07CJMwkW8U+f8/Hh/9pvlaYO1ZFw9xqSuu
jig/DuC0PTMAIhyJ4hOpX1Y6VeN3B0viGZtC0zRzeUCS99yhmiCMd0uByWfnqH/Y
iQ0edFZY/wl+vw5SH/KSB3yCpSCGUA6v3WlpmhqTIvbpyZGw6biIFYtn6KdtpWFs
qYt1khfsUN+66UlxOLwskO8GcazLrBYnHgvO7Fu1I1X1uCeExAifERaJELwOdAwk
WMsGSiIiEyZjtHL01S93D6s5k7pNj0weLNFr55D/8JMc1QoW6lv08dLUuGW8uk8+
6F25UzPBGyH8rF1oNpvqguPNeprJBo0JFbpcG4mTvN2x/f6Bpg4P79lK3iDWMe2h
7r/fSsgrOf4K0kbTbf5q8zbHeI/70TSi4fnPHMzKJi+IP6UXBMckoVVtIGLY8K1P
2ml8xufYlJWLhWCaX/RgHNUMWipBHmHk8ryDzpCkbXuZqqucWzoiVvwgzf1a5wN4
5KCG0n79afOMs6f0idda8pNiifO1uAmXkCOYELhtUtsF/d4sacy1EcoRED90KN9L
V/7+jHIf/nAt6bAkr4cQtuIZJFS1nNk0vCD8wV2D2X5IGLOeQWZPb2aM6xgDB/qR
rg09ujdtWxRbU1TsNwmyNG7bWHs6BCy1pXYH0QPH3O7cVncK74FJgAeLw8ArTLRH
ROjL+0w+EbsOWN6bfjcb5ZEHTKARKk1MQzofjEL7DsOuz920eZBsvndJxBICuUDU
azC5HTqc0l6VNSUgMQv1I7OSoTknSNiU/BMVHAtmHlhbqSYUn+9GLCWEaHyICUCC
ZE2SVuUmk9Vo8M0IJsnbYpmAaW3s61sdYrGyPk3vtZcCouRf6S2kPjvQCwpLzjz6
Jj+o7nTHWM9UTAFkvzAyJDj2Usj4ja4cCkkn5N3QQDgYvUZjvwczJnlvbFLqQRkg
4AkfoN3CWhXLVaDWKF5t4GC8r3hmWr6mmXopDhJeLe+CAxMUouCbK6/YId83fTQp
QTFwj6gD4UPNeaf11eaSW8PbInCK47V7FrkPJQBXtKb/YTdbufSX7QgqQvIT7aKq
s4/DF3dTyx0w9hKp2fptMzTrJpwk76kWf01p9ptRMCIm1ihHFD8DTZOQH6KWbTTW
/ouWSPiKXEm31Fz/wlfOKZwIM99K3tqav88/AOysukbQVExoyWm5m3+PjSoKp0YR
s41m0VR59dFpXl6qt5abVI2eo0JDoKumQOXCOyeKHI6ArQ4ovBGNqSeGiH8jx98k
ikoPms/Ri24hDA90i7g9i8cfHgrCO3ybgSPhiN8uJ/PHfL3EF1pR+UsA1Q/dNiyH
GXLX1W8BIhP3tSaJ3gS7au8+jAtiNeFLW0GlrxEpuqAgK3Jp7ThXU2Yiwum02Gy/
3d6vYv6kXL4fMooeg2GodJTCHKDE5smO+L+ckkT47rrpJjnyeXU5/Qv55bJZz6Nx
a6xlu3m9huV63Q4JnlLz1lsAVE00zoZSuKhocD+URgGcM2px2LrljbHXSocamCGV
d6DXk7TZCQePbPOwLdQNUJLynYQdQGkvEn/a0UC4irdsUDXFSldpS8EW1eKmG5N+
lIjE44nF/ARDSu0I6ymoWgk+rWMqlDYzEaTDrMUAnOBd9LSvcyYMqpKC6MiJ8AQq
ocKEohyiEDEHettk0HCeUOyT5tragYmbUdt+s+2+i3ZwOdzVWhjiMmRpF87erltO
6M2Zkpv+HjxowNY4pP5sw648UZ4drh+gJYnIJ9Fl1SSRc4971bYZKK6ewKQ3xfhX
BDhVv9fN0Q2mjAOMbbY/7PEb6Ui06C7vsc4D5KUUSXFgwH3R1BSHdE/rWmEV5Zhh
cCyKXTDb0gNfWsQlzxjGr4DWOGTOeZ0U+wOXKCRY2YvjwkuaesC/eBlmPPqNOqAw
qmN0VhiyF3u6thJgckVY77gzfeWnDr4VVQLiiuO0iVm1zoLaQix/Za21XaXkp5MM
aV6zm/lgiSAfOtoe7i9isyFlHBCGI2L1TuIPnZWjI6QFYR00Sp4QfJiktfgdZfnc
ZWlV54gmm4KpSaj1HuLmVs9437Q2u1Npe+23mNq8Gq4xleLUbcebqP8UEJ6p+ubG
d3cyYhwGQjJAHTtg5/lvGJw1VVex8XO3rZvJh/qnw/z5MHI/WkOor4veBeBlYSlt
qLTwT8Km8GW94JMKyKaQyfsh1gSNhWNFs6xYzSCZ+1LQf1odnBpLeOWm6AFzzWrR
nQ5EzBU0NBXkpqqwiFxU+WeWfSps7xMHsSzPz4vqQi9lnMpF8spPjofglKEkxEJH
CEF5yR/4bkkQhrgZRoVTobm1uXa+IeztdvFnRYRi2dBNY8tor0lrQjUjZW5l3tIl
QxNAuLKa51tfH80QWXzy6zAPw81pNWyd9sSm5tVlgyzEI1FCFgLsJzmzyQMIMQSI
Xl7DiDIrnBGH4O2YzTffH0W7Jp7FOJHEy1LzRIHU2q7EOlBNlI/ZcR/ulglxZ9z+
tDP+cKtyiqiXzgjvvsmPeaWq2HIdVhutmT3WzE9s/tJMIyFwnRTFrMYEQkKq+4Ck
VSmGPll59WeFBerG99KilO5kg8PjsnGNapK/hx0tlwRxYULPc/zjr5e9J0ggQNSP
PX32fuIxZkW7YSVjJWECaKAW6pdQR9LfDAMuvznnZZwp/ZdYSyCjq0snPEIyETqM
Mj/Rsa0eUmCLf7PGmv+qyDzDcnBV54cv66tegDMIDawqqn/A/8aNXUVZnxDxxVUH
5+uCH3nvsdProg24e4WEIETiKMsWfkKZGnk3uQJ1/BvsDqWikfdD3Q66BeCtwLGB
sj9ZWLnxa3Vw0VJbSCts+RptcTv1Fj3+CJGVXlx3K3CtOCY+jQlbFP3GcAm4e/VS
5h5YUG5p22HdH2M2X0ZU3PrHE3srl1sRcO3aYZqm3whgHo988SEaEQohXj29DdI2
aVU11kCw2nk79Pkk5/lrq8GNXk/UTAWLMnHCFIjpjc0Dmgxk+863X6wtwDlgnRFH
9TbhWSvDGTkloiIdXIrlhYZZrMZBbTNfRWAKxBs0baOP2VmF7epWKClJM1dujSlH
MJbzHN1lVmO9tRMErAmN5+adXvXDaZvrF0UxRjBLf534f6JChYupiroPtqjJJerK
GTXUbXo0QKufRgNJZjjYCqsTUBX0vfYdDRuGjsGdpRObCESdvnxmp/TPctASLkPb
48YxYJboCZzDCkeaFvvPDH04qdFbQ/oXW+qxEaSDXV8bjPFvRE6UIVjMtw8elwgi
xnNTSaZp/cHV/roNG7VwF+A00H0SGUY/dHdqoeF+OQ4yjmiFifPeKh7Au4ejt7iS
AXvmrmVMwyNdpnvx833pl8/K1A+SLalxvThGOX5xF/RTPCTqrP/LGswp6NFcKqin
ATSodQx65ommdfnmX3PBSd2W585KbJy1T4AX7B7M5q0wG5V5sTlROEdP3J+IsuuJ
HUI9ueFJH/x3shwTuAk58CTZR88iWe61HqqKSGHH/QMRZGBTdWwjN0UJjt8z+Sns
zzyiHqlvGN3FPmeOHOCacA5VrNSdKnNvGs2uXNgyBJLK8WiUk4iFzkGPXDoFAf0A
c4d5tvVZMYfgcDHiu3xlQcz0K18qVvkUug/aKJDsoH9Q64GDq+v55tnT+4w0JC5h
/uPk2xo5ItwgrMM2JJc8gE6xxMc9ghs5hNxlO0ofkFPzDZKdH9HzxrJPgG7j6BGN
P+fp4rQyTILi1/byo7xlMb7sk97Fa/U5uQSup8g3L1mgK3ia7/9a69uJD1166UXz
JadA3z4Ra4Rba1d/G7127za1k5vL1xT1l5A/6Wv9r9aKgaGPjTvz65TbMb1RFFPe
dRyFPt6mKXKOJLlpDa7t9nOWfMWotRJ35qdDYM6ACItsMt3HaZEzrO1WO8eSnf2t
5V7ifW1BLMTUKVpbY9ZwvL5AekNAmMANfpotBfWXvA/oJsBbBNXwtGeuQNeRfuiW
BuvKdEUgfSR5NwDNwNo/uksLpu4UXI5pOeiroV2R5PI4U8OA9Du3YWXhlTFmsHiG
nQu3lwvK033v6ZvBb7CItjtz6pbA/AMLWddWogvuuG47Fj1kO/vrq84aJLro2GU2
GQ20ljpYySTu4Q1nmdpyS5i8ZfFMEE7toqQb9r0cPF+cMRwjJNjF0bArfglDg02f
P3ObIRxfDhozk4cQ9sfAA1Wk6wbw6Nenbt3IW5JKhWhDoRqjWqNIR2jVGVwKidRz
83t2Yw+/1OJg2Zp8WSuDJD51tAUnQ+vmWO/2lQdu4VyM93bvP0ghmFt47qccVfom
sgTObLud7VCZ1Qq7FFkrWaKFZZRCyRULz1QvGIzgbUz4SUWWO/vHkz9pHWafCMT+
Bo8Rk0mqnQ+Vp9xMC+Lh3VYFEKXAnSgIY0kEkq0x6eJyyHFWlAZuLYRJoVCORf1m
LXzvC7txg+SVGX+YVpnOm4w4eUkaqLmhy9lLR6t8ja/U8Ld+HsF1bMHSaGUMJMyn
debHpCwwm52Gmm+FlnoZ/oh7FuLqlf9+1uqG7fmJwPX3lwjB+PUB53QlkE07URKE
RegZ0FjlTeIYsOy6Jcezwl3VeBTP5K40D08jjd7RpF+QY3uQmfRG80CLH5lIq+tO
QWh+GAoaQ1VFRjw7kzVqkx7PG/1di1IwMVvvm0QWlxaYOvBF3huQIIIDixkr0bm/
5ujxEWkcWonNXf7i6OlMcZGrVBMPPzFLyvMSJCiXtjiDBkiJjd9ifXmlk82/ahFB
p2Nrr3EjzVp3Zj9oFkH2wpJ3BnNwMmgx3aTHxvFZiOrk1PeoZl3YTTfwQIRCbia6
/Ks28buuo/PcB1r5Ci1AOgHXhseWoGRv5Xmt60OxqODq5OmWY5u2DiJNfyLAys1U
wKH3GOhMmVlpr0XwTgyYJ1CIPvtxu85UL2S+R5/YbOVpoWffXbUawJ6D/W0jLxiO
VwMkSvxZj2weXMqtFJimIoYI23StgggEoBkrUs3B7Upjv4NzMPFzEumaYp4gb91l
RyN24Sdm49NEdtfw5LTGWcBUunnTszljZ/9TxhnYrTv4i9fVai8rEGrPTyE+XjeT
eaRVxAOPICIYUw+rsicrQs0JbIM1qp9oT1qB6c0LKk+Wt04axjFpDDdaoan/ReMo
37vcdbfbj1zuDeCbG6+/CvXvk3kvp2HhddxM5akQJsdz/56K3jMfUTHS7iLiQNvQ
s037fJs/nK2JjwnjLQCHMweH1wwwHJJwWA7kuSZfdPNgbBjAgq1RW0DeoGwvpBOk
95q7giM1MIgAjY/qNkxnjZjif4ZsgT27WV0VoRbqFak4CBaGckp7ROhWzj8Z8DhZ
WYbV/9EOabdwmo7XJd2Rj7Tre8UvLQ5RHNAoxwEnwx2CdG+edb1AvSH6Ly/oQisv
rusQ2Zu0HBQ5BDtS/8xCMn4COs5x8QSrCkT/8cFnbcDEHUyH2Nk6zd8xV6jntgI/
ay1/GeMq4rLper1+bhaLwpRppUYN8uV1bIa7C6MECXbw8Aye146Rb+F1wd/DOgDf
QJc8B4Heex5Ov1Z7jX9gvQj39vg+Oopgm2NG5t9Zsa6k9d3jlQ0WmDXuydM/3kSx
NIDULMXrq3bYGKXFTYC06DidRsqNuKDIB8xfkatOHcZdp2Aciskvr3mC59gbPUVb
oSlcpA868JJ5Y/0aV2LICWrCbiSpfCJ6A67hXQuPfXSEj6NklmBi0AYAzSRNwwer
ZkGqf/fyO/ZfK9lTXcodE3oe00ap2zDMvj3+to1M5ILqTTpBS/Ca25w1o5jF3o6K
yLF8mB0tveGULFCvxMvJ2cPod0W+ySacH3CsU3DqsX82f5lxxCdzDanKTie0Q/Cw
hK2uxzpM7FAQJMYDFTlUrH8jWztlUGsNfulqKIccwXeknnLzbGTPCvUw1pzhRsau
jF4gtsaEzaprmaQSqjlZKEr+gslLUe5E2/nvoj8P6cnu+51ZRhMCpmwxllIyowMQ
HhLC5av918ERj6EsdE53Ol4GtMlPsZ8QeownH9JAgJ9dAXvJPQaXyq6HESTyjcJU
dZhvn4GYoj/g/teneVFvSHgTqZ46whIRVvSlt9iX7ofsVadTr65d/unX6Xx04MJF
qvbp8VnSVCjZnLMQKFgdWtpWJ5C/CBNGYTAw5BDBLR9RDf71FFEfYNMY7V/O8Obw
jxgcK0b3D+oPWN+J5OVKr/AlU2pDbsSTthX6HPxZaY/shPZbKdLYrHl1Fx12i2WM
AzyqMZZfQ2SrIX7MqPVM9+35NmUmTwJFWlFiC+lZYTk0kh2WqeG3SFCS36uuJy+H
H6whL41eeb3wvWiPVhSg3/kE2KX2NyBgFvR0IqmvmdWEXVdbbqoBDluI5zt5+5uA
zW3XB5jBz1yaNIyGLnT4COE+uoumUG9bqeR8/rWgl4kbnmKlEtmAbAm+pr+fhguh
bZu9Sl0nkvwm5lqVd99Yup1ot6UHBoLX7bgXsGgmzx4Xd+WxRnwpRebs7ei76kpH
Pd+LKWhbc5h/edRqY2a1gekc4qkJ7DYPlg37uT4ZLKMDCa59sWRddGWGcEX7MBqH
H3MCfofWD6pBnUCADKd8u27cY6l7vAf7KVI0iSZFIUOXBB1opN74+MxgbVAqFp1Z
Yi321jFtiq0/G8xhWbtMBal+bn6sY1+Jqqsd5YVXiPZCE7NNmqoXA5/1cly4ny+u
zvG3aYOFquVJkuteWudESsLRf0PzmycjS7hBNh6V4Zd/UpdPfQM83PU9T6TmuEdU
dLIIsRtM0lW5PHVOuC7Nj6WajfJ/oNCbC4y+CE/cycaKwU0a5XCdvVxSBwI7OhGV
dxWUOjdOoivH74DPeX4fnWZE9/9m3+ojUNzSb6oL0MvEVaz9Tcl8F8MpQaJUHEiv
8urGtJZnqicLkoScSRT4Lw0De7Adni1lM9Wc9rl0iLqMeX8jqd/ZvtlNz4FX1nN3
uC+neAiGncxbt9IcmNjxc0DeggrJv1zmKNnricyIvjXU7BjewWPXJrNny3XXt3rJ
ilvgXja5atfGUq2U+pJpO19zsqTk7pQfBoI+UBhfUm4umecSXq1BEP3Joyw/WzPe
inQzft6cf06ldDlCQ7GwjTqsMiHNV9zWn+sT2koGCSU7TtqLph6BJGr71PGOKGxL
JGkHen7WKaTIedwkZUVUIICrDVzYz0gqBYWFL+NKSJM9Z7v6D9qAQ48u2MR+2wUD
kjya9BhaYMLyxyFkIoEWtADVSJ0Ql/96Wi6WpNM6CM/Civ9dqrEDDqFKDm3T+RCj
cP23cabRBi+rVqNj4BnhCioiImlj1FQzA9F6Ak4+tvM3mlGoRf0YlToyboGLU0a9
MhPAq80JxMG8tUTC0HhQU/bm14fi/RmSpVmABpV3tFgPeg/xTCWYyAhJzktl6eg6
/flOOPS/cJNepSsYGuUe7zFV1MmZh1o7KaRVbAWO17kfnH803fRLyJEoHUKpPvcE
u31+DC27yWKnrcayxUbzOyY2sIGnQOu0mxvF9vDHtCbfHy+VHCKvyep1xcaus4jq
ouKIxePgV5lb76BCTw5oQBq2h9oWPnnUIjkTvm1DNskYwHuY21SSjhW1FNj3kDsg
ofQ/fY/wo4dT2vmY0pWnkXNnxtl0jb0awEigX4eWLp60dTk/Dd1XCXpww81h33wt
DG/ilK6NRTB4scFGTE/0DWJYExSnSRJa02VB55ueGv/z7KvxLItFDeQQCvJUHYZC
So0k/V/Md29bCz3Qx9D+TKhxGv+vfPAcdQEbHYisBQ/BWV05tW0U1EtbQX6Dlr83
946kc8OHXRMZC79fcY2ozRQrjjyTepA/8eRMSb3XhYfDQ8aGz7b8oeFTrmBDZ3JP
PRbH18/yfN3EdoqxGqJGUcR15sPJUHVcZxSW3Emg+BBqjxaUiDwY+sUL474qg1/Z
u1nMZmZlrWIGRcP0/YHNiHRTV8uJ4P/fCNUUFB5bmB/taDGYdVylLVirXpG1Y17Z
IxzSRbYTbBQuHFw0iirZnHJ3LgSdzzf78TmnVPZpOHMgRe4t6F3hrUnFNgUkp7Wp
eCeU1+YiKP5sfWmlUSmUicBLHo05yfjIbvFmfe8RVKOqrdySbOLmfv1nmnf4JPGV
5iwAq6eLP0JjgV+tNi5Cy7UgB1NSEpY7qjsyIJeFhYUT32JHOVzoj4x1/4BKtw2e
Qcx9FSR4DpfohdlQRAQqo0crS57TzMKlSSqeTsEa+zHp0xfbyJ59RL17YzkK7+OT
Q7I8MYOlOeld8G0pZUYzxWqyA07hdPI7wHoYaLlevbrkdqnqIjvjq9GZLW+G1d2J
BkAhPG19Tq6A2VfwHovAzQGxiBcLWm76DXIM/K0jOp0jyEDHtOkBeFbFuIY7LUy2
WXzR0ARDBctRj6che+idVCATo37sEc39DwJ+rhW9x0jpJE/vyJAn8PIE2ocYEfi7
vAFkcOCeT4sxBKDcn4UPmzmO7vYvIJuSB4h2mFpsIQbqTHHPEiq7zu7wZfPuFi2i
jDIewA+fHlYE9SGal61upz11X0BHk+i4lELtnuvm4PI1lHoyYMmqoHjX2+xSLwz2
WT6CfMNX5jScZQUaRz1zoJcRY7/287k5z3zrh69cfbGDYvsAfBseAjHeTrJ6X/b+
DTdTeHTSFq8fG6CMv/JmTTSVLYL5m7sKFBngrMez0+E9lucovjZbU4OjI/xADscr
8igIE9GldG52QZGDg3DgTqWe9ERQsEgZLO8JQfWdlwHujIDf726hATrw2+EBBdb6
7LydeuSCOtxg454bNfxFssoB2182yw8WwbPyUicKOZhZbEaVhP9N7KVftH/FtlOf
6I2HV6yDhDG/mIw9dCJ2tX+ryVOyJ5tJk8I2PtTGlYHotoa8lqaTOJ4tAwtiIIgT
27Fs/nqbcjtqeYlejlTbjYeHozQWw5pvIpkGBGgzPNr4QxP39RjQ0cKHxAG5HlF/
2CjJcCAJrtxCFAQlErsk0JKOPB0u+hmi87x5Hss7BVOhHWJ+Fu61kamFp8sxWoyP
ehbJAxv2G2A2PFrnw48yi40od4AcsZ8CphUiKfKJPnnFuSoDsB0SKF7LaJ8w/uvh
BlYC6672riv31SEohHaA+VDO4n+oEeXNDZewo0ThQUym1t0QH9v2cazTEf63xuIO
UTF9+0H+5aY+D6iUg4ZitGFExZGweNTDH/iEEOH/N8IZ5reL/4ojxAD3B7rHxHCp
9gDSS3uVmclzsz0IIJGCwgTkRBZSkzuolpXODrE/T+zAUifLnX2C+ukpL5Wyrho1
M6AdjtzhGYA//5+OYjEHuxFXEqAEp8+TkD9taNsWGF/YODguJHP0unlhvC1qRpxq
Y87Ku85ICm8QIrBSg+ywtC+mbAUMg4WSayZ/Ni55/vnW2I42Cg2rZ+yyOpfMzp/Y
jk+LKFhIm52aJC1E08rL6ChP52YucSiYJzoFPce1PZgzjFLqwUHJjUB70oPC76by
f8tqO5TfMwz4txbywMgTmPn8KrJB4YT/++S5M4VmMz4UVyXeYNeyJJXN0N0ZIL8b
/I6Bdk5tIa/wSa0HYF2wPevkP01SejxbazkNG/sHV8/XLZZ5QOtHWpmh90TTTDhz
xNzbJvTZQHARpfH/I0AzsBn01P84J+QrLbqwaIwrPhH4Fm/lX89beT1pvXOrRXDt
TD9Gv3dvJ31XWZ8HHfoeRfRnqhSEVnJdYZwUgupBUh2k6sV1ohIz/xRGuQGHbeui
YR08BVPK5bXflHuCLIbL/DOOWxJT5+oP607xDWbBsgMnvnRXEGuKHpK27TdNdJrT
bx9ENi97fZmZYzGJDPcCuXlAeRddu/jJnmK8ZyeZ+Rxl71Un8+my0R0NvBHz4b9X
yNzC2y41DDIFaVElDurEH1D789dofHxG/5PL4wRcsbsJNRI700LoNthx8ZYJ69Bm
FpIt8AkuHraOFrwyxQ5acldp8GWN23MamfyBvLFGo+1ab224aPpmWOWl6Bi+0p/S
1wb95E6eqglM9ARBe0PoFsC6IBImsokd704VNOklYOYgc0kc4X0x5DapeB5qPBDu
WpUYwqUYGS+FPhZxMbrY1QBY6LMDEglBop/YfeZ/CvVdJdtAu3rNyf7A1aDiP3tl
JkHP2AbPRkDO3p8zA/CiqoInThfoZKvAypRIWR1C/bMts9tY7fX1zW8YFhs2iSM/
Y7Bue/F+5AD24DhbJVaNGm3nGK1ogEoUXXDA1cHFfO+jakdBV4k94zsxxyxYpM91
adbsjb4va2FB1Gw5sdirvAcHwNh99XB52HqZEp8x1Ok/VcBR8cHNhrkkPn9/RVoL
nZBqRHkKwCKL8966021toZZmVSDR4cdGpcfGNumlWld1X1l48Vho76qjaAmyAvhT
r72sX+c36gBJMzHAeqWXw0DoyllWhhVMI59n/eGr157A3jz6tKG4inO6z2KLC2fV
xUUGWNIETVVC0SnWQc9h+xMBLToGEgN8PJ4K3IqjdQIyBiXfdJidx/myo9yeczhT
mVyBdWM8PGMKd7EWVY3Cm2DkgtdQIxSVLGOoZlBQD7DQKnm3WumvYmZSuuz6+FsA
ube+RL4a/bxY7vZ6fmLirJaRlEJPA/cPTExav+i8p/HfQFCN4iv3SJtNJLZ5rPiu
vuNhovzcCahh5cEN/JwmTF8gtIA//Ki17XOuf5dBl048K/n72bU+6R+oMHveXadb
MMJPXe89k2cijih+r0DIFmiNrCO6NzhaHms/ktMeF2VpkyruiTZZvyXR11gRKmvT
0g+RBZzl+C9iVvR5K7e8BA1mEVaJzNotyqTjeMuAEIEO1Jy98dO6GQRPACz/RY6T
BQ2BVXFoFMl2AiBx/XWutBYQXqt5pQUpkLjDI8bHUst7jKlaQg/+I+1WcAs5tZul
mp/ziTuBVHSqoENhT4UgaXNhTo46ARnzoD+8Qx8/Al92sQR7VsxXRQVhkWJK+DYl
OOIXGGJxLwFoElpKvifuSzDtzXJbBw+XjKYikmM9qbK/dR7gNVfXWdohy8cP3eON
gUThOkJwEGvgSYHlRq2S6pMMuClfckgOEg9YB8ZscsNUPD3TuDBRZR2hRqm1z1KT
8zWzrwKKJU/Mw9G4g6cKPJVh8jTm5HI9hnOQsp8PTCMXc8bJ1HByoOqcf5RQtaDY
yFK/r/GrHOo8dwKqBWNQ05tZaYe/CpAZM4KeShE4sfa6O/8bf4dr4mpMnc7m1edn
gwbx0tTWMPHMB/KgExLinILHu1P2aUPU3bGLIfnEK1z0ZleTiwJbdiTnw9dVW0oc
nB3tUZOM4HPws7PJYJe6mT5vhb7H/0Whz1bveeJxvjxj8sGZGOXVBwvMy710ta5x
ebd0JD64B5Qa1dfzcb8Mc0mSbkY+FJapadTt8n3bGmvG2cOiGbruGhnuiZkGr3q1
7Hju08IxnGfgCvYYZK+EOKOfHnuuCNMcSRVSbyYIDZAgh0mPhtPOdczXdH77R85T
2LwUDlPjkVx7luX5WYbkq/QG+iylpihUcJajG/GLgIlmzXKz/ntEn/kkdg/jSMD2
BSqKIpQPp/6wRhUcW3A4KFs3IA/hzmcgQ60E1HrxvB5NjQ6F1XesceKD6DuLbOi7
euKxPL1uOPUM8HC/f8v+XRL27tOVpBadZ4uWGFiye1nNPpJvVE22PaiKecv5y8mz
S/3s1FZruJ15lSrJecbPTDo+ZmYewrPiPKhU89u1Bo9w6ttSgKrJ5uFl6+l1Cvxg
CD2W3iVAJD/VyuG4diHQDxNMFrZ14bR88hriWrMDs6JLByM7iiiL1Qi6t6Q457xp
wBVBH02IqnpItp0m/GR32PjM4W7ej1+bLg9y2JyQy1eoYMfR7A8xD+cCq+l83nYd
/dn0cW8b3DLEhKQ+sR6U9kiP4x85FfryGp4+8ScTZhId2OEUE6NKgxe6dcu65NW9
BlerM9JzmOlK0fctbGu38A7ReE1DZjUoqBX6NfNRg7RkiSL8tGhrrs6hLFsdVccx
TJ3bqcll2n9Lm5kwqhvPzwE62bwAKRgEYY38/16/zwaGblriVAT8iVrbNlhZy15x
SlrcLO6VbEpDaPc1FII2mYDGuKOHSUT9zBkZc1TLzNKJ0A1mXgwXhFK4mKJDALRm
0P90CU64zhzIjUPUnkzyam7iuGt+Tx46vy5nKRtFs/ZPpzYqy6M2RN9n+OInAuTp
j0MQ/YReyEifpKJF0s76mUr4ZxIadVE5LDghkW4sxSDRPQN5BRSxsuEFyIpmojcX
pTzxKDK1vP5Vo8m7SZ3dnJpGJOK949lUtXnfb/5JckZOuhJ8RfF6ve1QO2QNAZAx
uBxk4vU2sy+hYb9ubd4wqzNXEWOoP9l0wlwEYoXiFMHWoWmRkWAzjpCK2jj+kBFS
aYNA9C1gjt5TBp02jTvuWXQqTO2fDtDFKkv58O0Kl+qO+ntT0ZVKKHqyt2tTxkZv
n/sXdd2zrdmkXS9fuddxkAQFuMbJip51tO4XWz5mfSyqmtTfPWO27GqfeP13bWOb
B9VEzhPjZsh7ZKSnO7t2lQ9tadN2FPDe6Ccj8fpOaW0oxVOZgeBlHIptwztx7lKh
ZB8Q9SxEeSGkOQ1TyD8wc+B51RvIPUuB/mLZYyu67UY260PwJQjvYmzjPOHj9kyi
sk1J5LI1CDyrEr5JLUQtupcTSxIuKJrd6TTHzWCvojmME1985JKgvbhxoO/q3Kxq
CtmM5NntOFMBjpfHA9/0VtPg1mKNRf3W4148X5KCWI6TDDu60KDr6EvaqRj1Y919
pp7LUeQRsaskP9+I5AZjWukU6prTeq78TlBQUZxeNuR6tmlE5VJS8vVf/8Tg4Vpf
X3zu8/qrSmT14EzfviYSLegfpXqjLc2M0p3iwQb6MSKdUGEuFE4tAYqU+ULdNRzZ
xHGvCYM9v8lm/wIDqcFF32V586kYMKOUdak67T8Q7mfO0OOHkIU2/9uV/dDMt468
moWydzimDm4hkxfZGKGuPtjAN4TKtwh2h4kuPt2kHf2J3ILW9usZlqdW2IXkyBj1
5APkMObRDS/dggQGLFI7nBUjkV1ASSot3DA8FqRkruDIpuJmVgiCFodxbKQvveYW
hQXgrCGr9+XRXd+l+FtLa7v8TS8DqvBJwYZzRO82Y/DHJbgHARaAWCPf4eB5n/gU
WRqZYHFoz81hyr0IHcucxOnaybddDl+F5XzHpSCsEteckxAC9TJoGgVch30/6u0Z
0P2tV8XjpMyLbQUr97iqFX6v5w55sDuBDoyP83ZVx6lFi+AqMBetMoYPtTIe5+jv
/QwvgAvbhVtqKXHA+byGCgO+ZOhX3jZS2dfxz9mYN049Kfz7ol5mQE6UZst6xf89
lXjIQ64taa7Qk/BLC4+JNIQaxTpjeuIRpvW4LO7Dh/TLbdoTnflT22HUdIFc4WlD
FZr1m0/e6h4AgG5BE9oDODRNF4BdimwqYiSsk3F5/uJYiI744HA0JFFLpVwY5dSb
62uiWiKXAEVsNzBNYCvYSSbPHV8rgBCqr/h9qClgmLuIjmO8DZzuNDB6sF1+NXQz
wrGOtRH7oCV3ClaBcip/kxUx0sMbfjnZQbrcCrufL7w1649sTapaiUekKruMYC4/
1BwOPSvJqctmfKVUNXRvKx8EVZJRIAKB8N39jfRAbX0z8bWZOEAxRc26Or8p00cR
cLzQtngpO6atA81uW855aI6hJVPYaMaOgbzxevXaAH5VQKOJyy4M8KyKpSCvuN64
T9Hu7x9KmkiSsKcGprJKIdsM3qo7E7cHw5VmjNvRerBABTSz2GJ/GkIy7wrHSnHb
muGfW3fXsOghs4GVl+6KG6Bc1HwBRs1w7BE4QrjIATg2GevnsRamns5jJ754Z4tm
kOp8H70+Dyfi/ZdyvGvHN+SQBTtJkb1rth17/cMvxj/9Gn64iRAKCht0Aq0pio07
9wBQT5QgqO/ODRaEPJbWC6dnnLGzeyRROl0ugBwV+tMbf4GxLWj4APf0YTo61i9Q
KK6z3acQ2Futw3FgcQdqM7FWochnYWXTcLjb/a1Ir+QBllaGeIXkjBbZ9Q4ECYq0
L7UwwXPKD61qcaNLoIGQzU5RnKRvLcSJ9LqV8o6joeyDTSi4TlRTRzp2FbwmMs8C
0CJyImMwgWLisfji1xIPsbvlsEeUJhLW2YVm7c8R19eHJXS6YwU8/IdoxYq+9eAC
8RwN/zkxm7uzoZm1rBr2yBNSUZP6qh5vmMA2cvYQpk/d5NZ++Y2CiE6oRL7nDiki
D6qjT2qK6nyWVMavi1qL/zIxsAeveSUFWqqgShKtVCX94uGyJ5uRZwl2r/GXKs5k
YqG3X4SRbaLzxAcJcOXnCO5aGodlrs9VfBiKBgHh/oRTNy+k+03YezubanON/ZYj
1OqkjvFUAliGvQyVIe3E1L5xogFRYZlhjOwEY5nFeiV011xG1CqlT4yfwC+Rbr7A
+lxxYtsTIAX6jjbE3Vu9DAa139zRt/zKIe3ilcN9yiXqMKhzqii2pzgmhEUy09AX
DKd0QZp1vuuKswrPRviiVff+Th9HHQzgU7QPozun+B0TUIQDUMK6jXKPr6JhW3je
60QvGIwg1z/Fh0Y+UQE4DHpRWXlXxmXLpo0wRiG8/FsdIfhldPUx1KwDDx3Ra10D
wbgXrtEI4/pl+FKNGW6pMYGO4hiBH8f7DkpeiVoq7psS+VcHrL6aTRE5jgbe17aH
w2Wc5WWvXrZ9GBFbMiQ8suGuSPZCAz6oCoAeWmnZbxsgzVUCi/kJm9ZELiK/A4GM
FhKUVxHG71bDJlyir+dsvk03QtPHhqxbolpVrdOofMw9ZruAdhrfPH15xoVZPkgR
OwjBq8mNeQlic6Y6tvH9Xk5HIsj2N/FvIpHLt+vxKYFB7eyMcIQvj0hza6J4yHol
Y6+hAGxCymWu3Li6s+zpb7sDdBDqqEiwA8UzmD6qWUreyvR0nASVGXk1e1Qn5xgm
lZ1C/+rFRbbCx56aCKCkAi3jQwVvnVpNjHtPR1l41MhHsNa9kTqM+nZD2Q5Lx383
GSzRMY8bX7oj2+F6BP8xon9R9AtfJStnrvsn9Ojkvgmu+Ic3mQF18rJ1C5dSQFhc
m6D4CzhOg8nC7UCWQ9ylVbcDAAPXvciOrk2YOjNoR4MlzxFKVlGC9zVovW7l1O6s
1mAauzu2S32B/8UpAmWrhi2TPmofseLKdqvyo8adzJ5z45d/tVXGsrlZVGbGGMK9
cXqOfxhjyFHd58hmL/9j2yAXSBJ4hkwQ1B6uAIFT0mX+2y9BpBwjo8CrOl8pp+ir
V1BmKQ7x6JJ6SuJf/JxLSGfiDVfkEx4vnnh2iDtQOcaOArsF7Vqoj2r/hUS88lSx
pTrYtXD4ZVFoNkIn5KCY/0mCAvwPJwVORfi7CqcESJEVWpnAzas2ANsgQ0BY25dE
Ncy5ghhKpFWaxPuEwD5x48sbB58ElCoWbQZKVbX08dZOSbsqndRRQvWLn1B483W1
ZOaV3V+Nfb+CPQEZS/vj9zg4hC6VyYDrBjOaoX/1X7nrWBiwLOMzKsUDkwkvkRmw
Qb23jK+Db+N4TN3/PQ9KQLZVjOjuwLhP171piJXynzezSXaXZtJNWhnUvvanNTCM
fvzM5Qv9tQy37Arrz3jhKVHXFNztKlwYJqiN20MIlRQ4h09pys0OcPYuw/kHYSXU
VrfeS8wgbbLQ3c3SPPFL81GAcQ82CbMOgF2GqbBU0qmUHTbY9mx6oHdo/2cZZJUj
iD7r1j0elPQ7wIKQ3CpgnPC8xQGA+tb/YvbzJhQB4ZidbYt9V002lnp9BQ76xtAS
1L39I7w2Gq4sX4rJ3roNdpU0KEqYiSszBlI7HnsF1a64oaFZPjxGSUAWDCcwQkBB
h8Izq8hP9pNt1AXMCyj3Dn2rzt11iJHa29pPIuKJpQ0smKvRZr/yB/s6UA71imgN
HrqC6wjrfQTZkXfvQd+tc1gQNaJz+03MGJT7uH0tgzPmfH8EXlksymi/Q5/nsE9p
daZnGc5c3j2HKHlaXlfk4yNHlJef33EnC3LnnB9Zefjw4u7jwhEZ5ekUZ9upwgmZ
lTEgE2MKMDYOexUXbUenUq8+lvmgInDAfO7U7Voa5dECO1Tyz7CNV26SZW8K3Fp+
wBTDQoeiEEwT5pl2w9kwdkJwxvtdJanlVu/PdfFqlvP2VR9f/CgWYdIAylD9wApk
i15ADqG6B6NnAYhctxMW9WR97ZeVmxjIIHZkjZSuHjvrevGLFNp8ZUKv/vWRnwS7
h3hl2aOQYSrSbCZPWTTA8UFLmylRBe/bw29UFrJDm4luaevgl/Fe7aHGAh4M1SK7
K+aB+LycHpN9pifHrcTY22T4r5lHHToCSvyH9I66EURzRId2uPQBQ8RTAkMeyIZd
5Fa/2Y4ad0E9naP5KcrxkYVUGHhHuwvj5xZb4KIg/kfIepH11Ij93rW6PJC9u0zb
6LCUiQmGgFIyl44fC9T+/AMZ8H+hWj2I67HecMeVv4gIhG+gwnUw4cbSpQ4HTpKR
mh6gO3Vd9xGrVgCF3REyzHlM9OMH5TwNUEQwu0+RVePwhZxaPekAA7HhoA8T9XnM
KViWSODjNHZnQn+CtqjLi/3pCjXpemhV3D/ZqAzLcITAC2EGGDH4IHxX2me/gBFy
ijSIylpPkMKTqURKN1A9VuTgeTaLS4yj5wpSOqxNCaKzUI/6p9t7E5gTNlKkRbw+
uWPHczbmVjEANAHImi894/LClbCDSqstPqzPfyqLGteeSHX4E/OjBWMyBGt7fxOl
2vH9MglHUYcLhFiE8w6bWtozoFIRSh/gbRPQDaqJqKUnG+aGCkR8khcv5qXUIyLP
SC2bf5/LDM07dR7eTt9Di4IzbR8PgXOXknPs+EStV8+qFkSbmqBPqksonG98HOkJ
vJQ4tkfO5LYgnB7mtTqh8vGAo2u5Mw1U0XOc9t4XfXt1OKuOdCRLAplYjPrfeo4s
iimF7/OZluGid2RF9lc2JVhXvBZ/v7jZ/WH2OMZdqcdKZjUSH6G2imX+UI+YYUUo
Rl/wJ0fD3mKLQ1cFKhWme/RVEO4h2BihDHkzza9YPptVHgDAq4ejmA6nidHdrLVj
ZmYExLtWYecHILBFMbl3VoWov4kY0ll64EckPNzisjh63XG/hyz3WUuzbdjpABYH
Y7q43zVTpgPbAldhGE5vKAmxCuq3Ui/0shKAmvsm4C6tZUid70wLBlCN/iMvYrtz
02KP3UlXt5ErbE/jB4wUlDV4R5SOWXfeHkYF73Qp+V37RcJJKVcy9P4njeEmg379
9eWozUcVC3m1zEaQrLVyueZl8K7A7wvtN3vmAHpSimr+q4RGygl6s7dhupQdoxox
jScRZIVM680K0ufGMfHNf0csMz71CJNatDpRA2BAM9iiYptdgRUuYM4jw7UetBID
RfRUOZZlH1eDlrZ6oRUQroNeVwqgH64FnVWtyrVB1bQN/rrWBzBmtLkASH2hy+bv
QkT1cqT9mBb+hKbkiFRb3Kt3at56w8VIiEQfI8FZhmFvNBSN0qTaxHiwr/u3bs4/
gG/oTlWlGoIUInhqWxiAEyuuli5DIBiD2QCBcNuHkFjaVHb0O+88c+T5pO0I+yKQ
RQx8pyJokdX5l64C4CCe82zAWO8r0mvLc2kM9ponqzWNE4klRI9TjZTBPE5uS4br
OFS99F2iTM+Cx4+y4DjTM7TgQ4QKauZFz+ahRVN3KSnTjA+YM1mMRRJa5KDVPJu7
xqByP7BBFa7nCSkwHZFnrNX9prBtefQ+hV/dDGA6KH2a+sArq5HUiKkrKQVlm89z
govz/2k1BLJ00pSJvWpaMQSTWHfHc0NT1Mth7WyNhzK1bdsPBOprivyUJLkqj2v0
dbqEdL1LJoJKerL26Cb/tzfy/TEd6G2CPHKu/9XaWQoihKzqbDszC7/fH3/i/b25
MCkQT1uuIcU1EeG+yx0TdmUVHXuC4KJiF9q46u94oZ9sVg71/X5NWIuViGo1/x33
tNKmqpuZp7ijI+FKQyFwoMdLiK2om8SOY930HPUqEEGVhKetuGyQAA8Y268cWmXR
0k8WDtlqp3EkkZ5wnEIbiGDulP9IZbqOU+YfeKrFuxjCEEKVRTAZRP/MGJKr/COA
vwmvFH9Yx0eZhbrR+Tpji4BmxY+detU301/VQSD1SEELGHoN7zrVKfjuforMnxjY
EGtJAnoDbMn1tRIuUvwPCXFacp8QvjhtobJNMOMV2IzE6aikH3S+4Oo551NCsCpe
t5xVrlirX947j10cbFgGNUf59Yx/2VRcWeDyxZKc4YXIN+k1L/Ut9ju8vfwFwtyq
tmyG/Xrf/yDM2QmxCrFtDvxmz3auAcdtqnuGXrJpdvfY/0aYottVE+YgNCeuiHlu
KZD8gZhAfWdgITp3ED8GeIH4MBrWlD2HzBrU/bxhjhVfeoyx4y9W5tkGsULUlWc/
8TtV7kZNkWhQbY1IMuxOouj0G5z3lgcxxgNcvwZvEeCIPiABCor1j21IN3GyqpwU
JS8a8S4oK5qpcaLjBNGfrv/aYd1ZlXWHkeMWM3nBjzIhmZm5EPiN/yZlK/ztodNn
u0eRLX3Ki1p6QRth10IU4+ywGBZfCwHc8OoRFQvnIdaklnKp82Cwar7lX3iyphiC
dOpCgFTJIOZBHG17Q+dnRJsB00+NxLjhQwcJb35PCYr4K9GIWFDruApD+jk32yU3
RmQjbMqBH9BV/N/bFdiLGGQWBXbVTfCfDFWX9p9DjuBdbZG0ueCCgyjGQf/P4rV8
e3Vd2UzbPPjsyzClJdkZXPWBmrgUyjK/Vv2ZB+KJaA2GAGd/8xriHZKh1kpuc0j7
udxkkRqwBJ2+whsUCN3bQKrE8+4I41yW94bor4l4D2Ccj2EzoIJZm1IyOv76sDiQ
zL7E8NgF1t1MLZAVmEmgbX3QxpTzYeSxosGIoaMtPynVi2mSN35ehpVh80UuJTwF
ifk3q2izXunGNST34nyI4Rse7N2rfCjzTsQn7Fk8Vax95Ur3gV4dYfwRIpoH894n
y+Nr2OXGf3icMeVKpgpZhl+RE2198LFcTE7XCvHQsmR85m9/kJolynEBUzeD6zgF
saU/kMai53l4Hp0L8QR2T/PsUoJSOfq51HgUmOHXso7sFwc22KqfRJ8MSFnAngB1
B/wzUVbxMl8W+H23LcysoKyXNXn47Wy2weMhKSsZc5m72T99NXZQqHRhXH5jj9fh
jhD/NLlBo55M3Bp5/SgpTJ8m1AX7do8NBDdmg6s9ux8RicKFHCqTfW9LYw0Z1UiW
0ytZ8VvBG0cjHVGaxx00wlUGMB3uloiVBdeTcupqe2Y8EbIjnpB17uwLsplkOsj+
YRAZkGbwdnQEyXZ1/LhWUBp6yxNfq4wRzsd4XGV6BZNmbsAas8asWzDl2Npmn94F
BPUI4qnMqMUJ1W/82OQDyiF1qUf0HNxka5aQyHSHr7DDdIskvy/mh6U3CEXHaeQx
RjIk7noHqozH4WQFUJfb8DAYpLK45wUljQqGsrNbwTBhbaFLt+FD+CPEDmSVe/Qk
s3IV5X/fHwg7HJYb8IhynWWx+ekK6hoa8rU6OReSaMQ/6np6sm/1BEBxH6UIDMk5
zBpUS8blKv6bI4P5n67L9YX1o7aleiniq+LS1t9beYcXpFGuczedQZ91hA1QbQm3
xg6APYoM1onD6utb/2uU/nxyZDoMuCg5Lyh7UikY8TNeCE0Vve0h7NhXecRlfMI7
2RX9ok1TnRFehbB8XhZo7ggk+/s8qLzBASBz+0AFm3T2icwiizlI//Nunittx4OU
87pdydjlPAjmgpSTV5Ob5Wo8sZCE2JE2cuP99of7GxYNv0CZfO7kVB45S11UBU2d
RXp9UN38b2qc455xt+zlSx52f5Wj42jXArE0a7S6ccsD4vnkSlsVURQq9IlVPpcq
MzO4lL6WbDCw2M3vFPyrrXVE7fnz/JXa0A/b9lTY9y9Z2pYgBcmDRytkARDQCta8
t5giIztWE8MGE4oX8ICzt88cHVJzxltrBz/B9rvKPMetrlEKc4Bx9MCcObhkbx2b
8Vd36sPhk1o+bFtxV/ZYkwW9CAaQjVG1jOqbEJXHT+0UmZ/SD+SXICGznHlcbRR2
COvtgWJkLA5o/K6ydLvlq+MLmL5cysUiTR6O+YtCxzvH3pGjMTFauSCpmIcZ3cA0
BTN30BHXuR7j7aRBGgmHB7kTff0YqMYKR+UaNT9FXI5Vaeemb0Bdg9oNtNfg9cHT
5DBwVCR1cYUz43nCklLXsK3Rp937jlOhuELCbgz5IBDD4c1l//2yq25/f+aRC/aV
61RkUeKTclJllsdZ4peGbugCGUiFaavNCcCDn7YhVnrRVEtpUcRuDvKUu70Bwa/1
e4QosfmPXikpgW3P6Z49NQNZXYvpvhGv9IPvkCfE9PO1KuwsUCJ+HrKKT7QByjKq
5tULsnFEpM8HqI+f96I2tVWsKqo9SsXyicZ9OhvNlFV51QjQbF8raWgqQ1NlgZ2p
In4P5xs3OQtoDrjmxuDsXqcVdVbgKpByYdTHYYpIy8xMRMlOhTtVUBRvLvYtZZq+
F3u8Zy8vJNU4PwQZXMg2DUzRWFhRNDaMDxqz4u6C3NUC/6wmtRcaYE916JbVSAMp
lWxOGWA8+WDFM4l7B8lIX5d4nAxpBE5dO6U0PpBjdTdzGLBysSoW+KQGIBGXIuZQ
7ml71n/fO+8DSPe9dxLU2o/qRNHuZoiRONQ+70ybTork2MdY9LgJeSYYbMzG0pHY
jYZ4yunaV+r8N9WAlBTSHYry96RAdZxzC3il2v05bVDlHgMNVXazPhSFONxNC1De
TUcVdkcyqjDaC//HWdy9pRXeuj/pTD4By59sie4xuciRuJTrhJnvVeEPE6vLksPE
I+6MwGIUKbT4TtOhIb6mcNcbR3TSuUPAbTNlnFriog1sq5yczyUk450yJyKWjMdE
ZcwMpUUupmMZHk5O+fk1ByQppb5b8PPHfgGXWsg/iX3byG02U7WCBi2NUz1F1E7r
ThCBl5EOa0YRdEIEFWHM8LVKNPLkmYdOt+C1MaCw0jz08BBwXxFOq2XGBjffhV76
kmTrqrLvgB2J3FvlZycW6yhPjHj4W4XEHogVoVoqvjZ7/bHqLofMT48CHcwzF9Sd
M6Dy6XOcGb5CjnyWiP92WbIE6ersd0KCCM3l2UAAquS6qiZETjQWsDRUa0GEs0WB
w8sNhweVxqKN056l0mhfMfP/U7SlQ/xBnwrO11KrbxIq615J2L/pqNRzP1xyfd2d
mwPuWQMXhQ76+pvGmcWAmq5mcDJ5LWLwFvvpykq1nzoCODORpQ/uY89hepHo2UuS
9M/PFBLdrCqlFm1wNRTnanMr1J7cdD512osO7Wk6T1rc7V53zRMtgg5QpQZze5bx
TAb6YZ8r1uXj/d6lFYNVG/auII7j+liHwFvb2gOFQsxPsJ8mMowq/wJuvVp2xgTZ
32rT5Oi+uVa+2rGvqvfHj6C6vTfNuzXKiIfcKgjAUTVi4b/PZWf9igrVBKbBaW23
SMrxTe+v+IjMjJpUKdmsthhzcv7eGHOLgRhwZik/35snw7CB5x09ElWuy0gyutZJ
QeWNnEKheZ8AJl+GOwMxPBaczcUlAFE09NfdRxsRHwEsCeiEyHaRo3uq/jIfk4fo
iNgyAKgtEaIZCogRG8y7Yswve4d8CfzxyaPbsHxNbV+z+6Z7hzaI7BmQI+ImUh9C
nUm/He28h/x69kys2henQ8hUAzq1LDk+ehWc/wyLU4MkOkN6mzleAr9M+YL39rmV
KZJGBB8QCloxd9E3DxaQWpSntFsBz4o41Lenhj7x1dYU9n6kXX0m1QG4RvOHYXCo
+eXDoSl+46J8I43D/m4Mrdse9ScPpL65eIaOgR73a1v7XmGW0WmiMMtfDNpsi0VK
xuOWyMv/7NMYQa9wzSqG2FkN4ncAYydL5JDSm4PK7DBZ08G3yXswpRiMvi32mdJI
u12V8Ehq2eNObFKKcJEYfPmd/Ur8aLao2g+/UZ3pB25oAfTkh17zUxHdTS0uqcnf
LoEQ5ilnBSh3FV97OlfV7P5dYfeW66GUot9AqFNGGONlZI/YvcHy6bmm9FSjwpAj
XdPgj5o3pXQJctEFx0+rLhk68WlXmcaT2dK7GjSALIBaQs4bpK5fmGNwKvAceufB
V0mGNcFnmsYH7IFeMGdWupEFw0mk/mtZWJ1m1CdJGvBpuqYFGK3W1TG+li1OpHax
TE7HcX/xvz/h/tcFdP+OSsXM4o5IW9/P5huQmSaTTYZeFUxIge1orND/ZcteZYyp
MHAHi8ME8sE87iJWO/EN+jiksrFtTqzE4rhkxbhvU23ZAVLZSj5rPY9kLb6SC9ys
anMsyj2RUxM11tWmmEJTXQKAWPAIp0SfWKirVW8nAuaSb+ZIptD7bNSCQQGupDoK
lAzbYaJwF51TrbG76+7eccJyYuerkm4QKXygq2hKBV0NyZUB7ycRA48xeIOeYm/6
RwZdamzL8UrmBqLBtEAJ98SSq26GhUSqcbco2GYGxGyjKw7kNWwxneN9EVHpPTJJ
HVAC2w5GxfCUYqQWoH/djZTknI1pDcutvYHqXiN1vtyt1w/A5XbKI92IuShbXfHW
77FOKSGH640vytnwHW2zc8gqPpmoTLA1Q70l3I5Lwfn6EDSgx5oCkKyl7ELL0DTQ
63Mn4Y5Fzq5CqWHziIqLEJQTWauSBp4aMHxgSsgxnzLwpnLLnMASohQZJ4nbBMHu
RCYkmujRZvE7HjhK+j2A1ggqhxcAWktdQ0qCyFClTqClfyznB/8F5hFhLs9Bk2G0
YlNAuSUJJu/ly4X2tcF8A4T8lZuozOOypnVqtEb5EnKY/fPovrPvCdNafjy+jxpl
JxJok8TGS9devNjNP04OKgrJaXRRHpCMSyd1jxsUfW2pO5AxH3E/acKsnTPcyMKh
8VR4xeQ95Qo7mG7KlvAsFlOwVBMiXI7E+umydR7yYbYhfXyiDuA96oIdSnP65aea
m5GilwXaFOoSjlDNh4Hen/JAYWDMIFtVhHRWuJ2jCMDfFil1VwMQjmEOgfWGTImE
EflHoh4Sn28tFz9XUVxCjczFPlFzKT2A2JfNoasAt1swxP5puZb9LhiJS4dXaM4O
y7m+FZ4hXtZC6QKKQHyKuiTSSIooDJPII0Inw0aheC72olfqY3yz1YzbG5l1f5GT
B3c9CJRCAC5AtSJ70DNmoMAn/wh4LCtef/D4jCmmh5UKWVTsAh8l6BJ+d7oBSJNg
n15T+aV1OCfhm8IBK/crbJao4Io++Thbx4LCOYWxyHHTSrJ+hlWxBU0a7f8rphJc
vG7fvKj4s0wktk11XoKMzNk/T6UCvvy+14qwxKT3FgGlViOqpM+XOVrnC+t8E0ZV
8MqFqCMHFWD4h4evYYxXXRywFCf2SeudRpTKNmm6AX5eJH6Dz+KhehyyriTOypt+
fRmV5cFBVYNAlMJ0NgIzovYbKXROESPLmZgjD7XUOGkmjmnlo7bMF95k/Ze9wppK
VIMRm9r7D2U/4tvkJr/o+VpcEaiBIJqRi6FETsR92tR4A8vX7XFirdGz1N2lv+EI
CVoSb2OBKQXYu9qxLDUuiK1E1b7slBw0AFbcXCAwAHLA+bilvTranf7kDLDUD+AG
KT/kJED6ba6WcLH91FauofE9rQyyMu8qKVxSb3QbPDDVFrVzHQDIUbN2pSSQ9qTy
zSMATdTJtxTbfiPTtZwKTjyqag4GtMh/1XqEWPdpjsBNRnItFDmL8DXU3symqAMD
EFqAMvq3vblGRheeYZ9Tp3IPQI3hUxHJmU4x9c4rk2U8PaAdTzMwzYYMj2CCACjX
0O4paHyKOcCkXZ005cCLHMbGe814nNyLmuSuwADArJQm/EB+hr7a1t2CssAT+Ciw
WFV4uKz7Fcmv2BsTWT0kqekY6RwfusKjk7M+ETJt54x/rHo4oVsJDotRBo+xF4az
di466pl/cvVv0wXKBRn8ELZMw194Qi4Wn96TB8SNRigUuSpA2hSXfj8lV7bsj1VG
CkLd6ES3vySLMiuLlAPVIgpo3qzvRhvajp3C6yhUikRdA9Vv+XdnG/qx/lnvGdQr
DzJJwWGwcJEMZh/ISTa6sSpQlgof8jaOGzxhe8GWqEYV3SDkWTWTglXoXL6XsmZg
wI76KyCQldbvTRU22TcJmZeAoTkSRZ8lDLS8F9NKWqFQx2ySqVQSXipCJLXdhfS8
H74uGiZ0Zb8k2dcOQIaM7+eAE1YTLpQt8yrClaRsRar8Hwl0m3Asq3D8xO3cODhp
D9T8NGVRb0XYI/8FSNOZKQ1epEY+NBaDsSobLOLzWK57Vx4CYlP+ZctmhCol/+ff
7CZ5bthHcVAOjPzns7FUvPAQTTbkPmLTGkPlZRvncE74ZSN6Qw9vAI0RLHEl1UNg
g7lJpik43sYKEVONpZ8qfG7sSFS43nGjM8WjM27gSwDaxXmiEdIGAaxzNk9Yf6Xr
whnIArX8zVnTcK7cwc3BqA2tsMnfacGmVzzYosDYBGM7c8l/A3PrjhicB4jp3EkP
ybkA+YSBQ5+Mq/fPq8fcYWSgjXis4O361D0S0KWsSo/UAyi4oOSuFdoATpmm3NTf
`protect END_PROTECTED
