`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sg56thhjUFiKNswffKOxWeR8ayMR71bcHhnK9vHA+0SAvmZhBcoEXepzz0fac28K
FhA9I5rTrHjcu3BghvBnyackeiioxsPgqZ5iQDteglTesH2+0hJKarwnox3M4m/1
l+MPFzflSCeuBj7Vot0xN3klQFu3622upY/rGRAfUornTCxW2MD2OEDpRq7J3mRm
S036PLcPlLT1NVvg5wumgtA8xfX2Rixt6Z8iEEje7KADo3cuZ7AsM+SoLBlcBSWr
UnxyccSa6YcFpBpyd+eHmwDrDqyx2W9UhhZtzaa6bJnlw60spdKjsdaMVtTFswiF
l7gfSrPfg1qdpq7G3hMiCJ86VnbfyqwECYI5M0uUC5oIrNbL2ni452XABS33J9RH
K0BjJtmth+vRh3mjRmduAWLxJjhRF8rGPuLrxuFHMIkTSO51fJe7UZGH2WgNi0ey
b9zIjGwQXu2fUJyaFsuOAGSE0Okhe654j0ZVcOeRFekPW/wjIYGwmkNOgVw8u9yN
Y9eBsQr/ygwbPtArbctGQK9P73JCj6eFpN0RtdeVRsE/j2Sj59fnbS0i/BVszFzK
5PFhXs12x5OwV1eXrvl7BRctLpBDRWTE1k5JaDgpJcTDEAmM0fyquZhLgm/rT2pk
CzpKmDJRVd2lIZD0xqzWoA==
`protect END_PROTECTED
