`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wPKOZbNiiHcqc07PfKrl46eim0oNygdSKW+VYpajLLnETCg0cpfhtItHOgvyqgQp
EqO73MN/qZ4leFlhbC0WVt1ydghzJ0rXC1qDYpay8Sox3+WyfIU7QALJ+/t0nBwA
6sgXREEj4/OHU3f1DzvGTmEd6Bu17sFFNKxd8sWlqiBd5mKkWa89fDv8tQGiPFXN
ctyJCgOWyf3ATCJq5BTbNrjBRPOq5IGI9lV69sCa1iHSZuo7PNgRgTe+aFZwhs1O
R1kaVqsacdtNe65YeVF8765V17+za8Mm/2MAZdfNZvOYX7XPcB49/VOvA5C/9sqy
KyVgDh28wm/WKJ37depQD46BZfFZds56Z8ldTjlO8l8fVc+xs6proRu/R4Sdfvax
8GyTbbt8bju0Y0J7j3GLRqrGG7RZghw2i1Dxkv5YQQypDEovVlZ4m3RZEZ4JTwEQ
DE+wtRokhd1oECA+GVZn/swfpQZS6KGUPn50VIeL+9rs4nN1gO7vWicgHt+SDf9V
o5q/62MOh6KjExExAp1hUGIKqNiJHfToguec59HMiOAYGt5Fa8+oCEkoMZADwYq4
Bk6MF7i+82HfUXYGl+eV7jtXdpC/0GSQl7N28fMQrtBZ0JPEFctXUjzdCqlydVAE
/W29/ucBJmr9dhyT72oSHj1akWfkBUYWnXDzmKpWMUPYDRHUZitzl5ByviRSjuAj
5/qlw/G3jyvCWCAmBnmssx7U/PmKXhQvBwsR+41by1y97Rl+k8HjQc3hg5IfLUP+
KGq+E8zybjq7kmICd8pcwV0mLTFXf0o0t/bKapho/lr7TM9NclIMwiqTVZc/GumX
bqbXcglrifViRWbZsu9d6WlUY5mWtG3eZzm+0feBQryalVPi35qnHg2Ry++1pa+a
hQW5egLyWsgsKEzS2OU5QhI/AbZ/O3yy1OjhgJQ1JkDW4P/QDmW9hw/RomrBY8qu
Rfj6/UgO6AAx7477MEXZMyt1/JkLDCfzTyXAVOgAV9lCiMn+UNYz00dmXC//8ID4
vqajk4oqvqDrXdPwis6/CVq3QwXj7/KYdpvwrlyLJNOUCoDWLojU8TOL23mGhHsW
ElNbCZTMxSY5mA6nArCdrtOWwESe9HusJRIQZUTXgHpcAO6KN8iibLeVZ2Npkpsh
73tqxwo5sIaDhlSOxO8WvaITGP8T0N0g33AHJcOE3T9/5lr6rh9UsKgtgT1ek1C9
pYwiEP9K7lx3l/oqVjMyBPatZ25FVgK69tZxyw5TpeTLPE6Dw6G/MF/SgPBYwXnl
vJulbqcIlInHXXx72cL//lq+H8fcSygytUkcWR4PPVL58MINce4AuH+okZXxKkwh
dohAyAsbT/dVhEc8sTxxIjPGRetGD+Ss7HXSm/ka/Ae2xwWOGCUnhA2T6brdP4Gt
tPPGwEpUpJpoC83j7bA+vnoiUpNS+v0VKywrR348OTjqtzN8lO0u6ukugPTa5qZn
gVdEZ061kYArPYxmuzt4sy5xDtv2bMfn5JVI1pTPK+XrLTjEszyQI8eDV0tOIlBx
wpGT7iUX2yIxd322gCPGHLcGQUXCkH7kRYRa/OEYSv3a60a8SEBvElkKiE6RScXh
7dA21qLpLzG9zIOSZnIOZ7Gw4cqFaAg2Hje5AO2liP7WjrWUBRDy3wiARYYykaWK
O+XA4vZGLBbC5mFawQhySLYYDE8bVC0R0qwSURxViSNAUA8neb7lpjw6LiOEJlkt
bp9hT9wWUp3Lc8dLYThSKPombuoRmDB/tMZcJgGK814g0JQt94zHGrjYIf6CcU9m
Ii2pm/bfoD8Oe1p0wWWPNaaEjtqJzW0LzCnipZPVINGqgi89VZUE/zl9fyU5FDQw
seX5uKqUXgHpnhd8YUcAKRxoSvPMI+qOB2vS1NJ5WU0mkXAERuI61jnXL9UGoFp9
dik6pVYOdVVF15sp9rZm23Qm6VcmXs59KgOpPSmxeVPKnxKJt5J+O424HxX2ryn+
sDwNiP6AImwtOwRE3mOEsEr2eMy+DdI+tx2gMS/IHbh6Rc7WKs5pq+IeCOiLoyKA
DXvijo0+UTnh2L2jSEuojY2qsMYigmXEMkaxPhIVpqFJ/bXyQ103taQu1AGrVDtq
h8TadGRSwNx2kE/RFspxMSDTRT072x87AQr/sgbOiPF/dDSgas1+a87rSWWx6Bkr
75ByMn2iGox6xQ3Qh5VfxAYcXP3035JqcBeWtUV2YxuLafhQeQ/AxuMdzkzeSTaP
+LVRNDixhHBQLzrd/FlWgkxcuDh3J8nu57JiEk66hoC+Huw7wUSK9OvqQWh8P0cy
idFp8jBxThfcvmUrATZGrFnwFatmP8EUocZpTZilcMxv7ZQsnDRsu69iN0LOc38W
ZUTnnTArA+0bF3PBwS0qpVTQPlEe++FST8Dy46rWEq0RkU/7y+duNylhbhPCpX7b
nYolmpGEH+js+s5HpTpQOVsnsa9pBwq02Xk+V8SaPmJMfHIKBMs3IcQEf87pJ5Gl
BVhFnpP8nQB7Fb5CK5xS4lQIlnoUwc0JxCQw17hZb9owwg/4FFb0w+keP7c24Uu6
CIaRadf50Dz5h8TaHtKdCjt9gB26cHPng3Oa3XvadBLrKjxIFcfT3xyOamUQphVg
Xwa20xL1OHEWTQS3MrTWSFC/i+vGFHZq2hBsFA8hAbC1qAjER+KjrvY4dM1nv7Kn
IaH0IHcrUIdlNbppPdJHHeFJF3RoOifKNVadz3QDrTo4jyw7iYdoiToeFjEfaLlN
JfBmM5Qwx2cAhm/tRJ1JT2e1jUvAlL6S2/+G/V1A4GyLCT24CQCNoHWXo30QLZQ3
6MaYiqwPbAxDJZu3mHakdVVDdiSYnLcCwnpZzCVl8Hw+AwfRCkiR+/bRelDD2AzO
DM3hKAIt1k0ocExDMjmF36uM8iIpeeRSbkP7AUs26KO8s/X8LbqIeg3QXA4Q/YaY
/d0UCdOrab7LcvKy8rHJBR2sdHwfUlVOLZoaLNqywbyed/yg39RkXgcVXETqWC1o
aSXJ0RtP3kczLsJIo3wnC10xsHxeOMDoXvbrfVfOhPalfgeEnUwEbXwn9S5na2As
0n3CqZawYD80V58uz+mwFkXdQQjAQ+ZdtWlRhBiCQqBkd8r6Fl0EjBJLEiHy2uJZ
ErqVI9UPvaX8s1ItMVAus1/pWDQauH3yYapqxklr83cP0QTOE+HsodgpdvvwE1FZ
1XjrA8bDNB3bMNkcBXcaXN/eG+gfNqny49JwCV7VaK/v3GSm9di1UK4oHImnV/FF
sTIssyv6DAvSwXe2jFH/o0NGhtvJDJiUJfI0/US+ZpU2IS0ZsDzGAUmFRKfwKC1T
1hrSqUVwM75IgKdNth1F+xGYCIbWpi/tXTgvQ6QMd+DthEsQi4MhgO10XuxxkqEW
3GCrN9Z1MyfkQpVk8D8McGkZGMMBo+tfwZcnPCKoqSWbxeo28iyawFtdvgnvfQME
Tlcvp/YgC6FXZ+TzMDnPh+qZYxXuzNzejJPIkMEiOmlWHhymvsRw5t77MnvKggiu
vjk3zg1hXRRb60Oci+Z3NIMlhm0m9C+ypYIv6Vr+mIiTyMzbRJnzpCvCEyFXY4qX
nL5KXrI+mDB297u6Ds+imtwJPAyhgJvu0U5/dsdkM18BAFysXUfImW6nMpjmR6yB
TCZvBFhFFjNtrpJ0BC88b0J70A368yZRwA/+yeXbrvq3lH+iOF/l6ZIGfeSiWFR8
YbDg5hQItiu9Fsph1S8BQ33ChOljSz+29GUZzbiqAU+bzs5L0UjgZsZICmnu/oI3
YTmNa0jiEU3o8zX0ukYMBCztuZebLLCvZIc5C+043zcJu6gGUQ5u3bOQODEpAr9y
FJ0CRwEz8xIzUWfBnizCeom4xcFR1trDx/APxvq+O9DUXgq5kd3vxC1gDbefxe2z
9edfvE4kKZFst0uDBila2z0p4MQU5pncRAvz5vOgj3OynjwJP3wKqsBRmGRNH4+j
5Rgg//fyNGx3iMCM9NKmEL1W/UGjybyf4U81BKgsY60nzwTuR++s9/wCHrW2aRz6
uHH26hu2agg5e6ZZLwaAq/yCZauOUNt+DmWyFb6IF0IvPA17BVGCHZ3rGXvfXPoK
edecfF9dGkUDP/YOGUuhANoOXl0Bmn0EJn5VdJiafgCCJJvUtdp3h9+7x8XkclTB
EfrgJAWIP8H4oGqJpLSLgwCE77eLcvVn09SrjNGpztu6MxFyrgK3/AY67DZyjCkk
7t60JSm9ZkPA6XN/6Sny4Oe23Xkt9IVEUB8enKSQQ5HqdlXlMGLDbAbVTK6dT+fS
PXlq1CP7hvoA5o+s+5OfCNWLUNwBtGnxNh9VgzmG/uR21n8n9gZJVxEYRxGDnLpN
hR+NK50TPAVnVujGDqVscYX3KWEeF/wiIS0yQPyATecirXgAsj78/LbY2skW52zO
Ub52qUUel2QEC4b+E++Y4J96T4k/4KIcEOX5GPCJVh5ctunftM8fiqKMaKBHF6aB
+CvSCcI6gsKtwbYxoENt8dMUqSQRuHCxqyU7wxowEzyDRAjZEm9FlC23VzYk487u
LJ+SSVkWkXvMQwH6jaRVC+dJl4H/akP4tklWu2qHOiwEUIvc7zY9Ibe0Kk/UaEx5
Q157lIRWDo56sQJBW7c5cSbdih8bY+abIXikpUy8mJBrCtjtxYDVINHKfrsRCHin
Xj3CFQaXvToYD4Su0M+yaFGYgdCYr4KXRzJU/uIh/MFN90HaU27NdBx5vVMSkVAj
lmx/pt7Rjh1baCwT9SpKU3EPKmPZ3kfNmV7Ht6FCXQA2twfDNtg+Z6MrlpOlCE3D
ZBNdNZwTABZ241N2ZPXbkSk976VWhF140YZIbA5WnfHoCGqf0QQ72PL9iTBdC/Zk
/L5ceb8KzINa+ureh53ytbxjvlek3p0wczVFY/2OTb68ChS4GqGHvTycCB/9+c+b
d6TGB1O/YQYT4LaYJ8Tf/e72xHlVtoViwGAVDpzRp7aUuFgw2O6T0zZYn5vvB15I
9HYz+SUZn6qeCzfQ8iZoV5kC85NraFQjGCDh7+RHTB7ht2ncbhuI/09YREbiDdcK
JFnqZzXo7b7J6hzVjhwj72rdarx69O/HuA80fkEHoYUjj+7Xinf+u4AmucqtodqQ
v8y0XhuZ/codek3gSqfz2M7glZorC+y81IfKF7bal/DNCV8rJPlO99S2RJvpJ+u1
zF+8iGWaN91KxfxRkWElP37nKySqbQigNR6cJb6DeJVbil8O0OwOF02SCMnL2o77
a9jx/3IcZ6hARZUA5/CX3n5dyOmqQRUOIRVBn+JAjEEKeWyYHae0toEq6xzfvXmS
OljwpCGXjGesNVX1DBO1Ij5t1VDdBZwDoS3Wok4hRIwO+p4Jf9+PrHlPu1wjZXO0
7VrAw+ljLd1GIxtTBEJVZglf5TDrk8N5+GMxM2M/9iQvHe6X4T1Qg6E5VHyjhrkO
yG8xUTYNkBoMU08YGU8W/kpi4KJB8jYMB092r+MNFx0wykBNyYfmYKaRN1abDCBW
P5jdGUw94pit3HWQkTr9EAUO3QcAVmQqxtC61PzOTvzx+wA5ZEPOFkJoel/mDVkN
L4ajlRp5iLqz74C8wdM2FBwvbjMJlpIeaOXPMDbnV301pjwgj9vd1BB+gOf2Fmoq
TVevidpBViuVZ481+nvw3eKjyqAKtg2AuNTKdmhE6iaGb3IeKYB8XfGvQPTl+WdZ
Xl2uIHAdW9rqTbSg8UFkE9kPAQPiFDv0mEfu2EgaHOQFb04TvTA5SVZ3dTbd790I
e2GeLvNISr+KwpwgrcGcnBbSxZljPRhoJMiBgz15LYUF50LsVldsNsFxie63ZOuW
7O3lq9WzjYg1IQ7rlgv3Xz4GXIbyogA7tZOd83YtDPoemad3OH2lfkq4ZaE91Aup
Az5TIEmZfLSWP36zW6fRoeverl+1XqTZmhoIeB3EFeGtvioIAAJvOZmM8EViGIBq
jzxLWv8IRSXvJ+3MU0zXAt0kv4v505+e6Sf1ErIpx99QS0HgdBBGy5ZXuw0G1zXl
T16lGdKHWeDU5jk/LnnsmevmgmqP9IW+cR2GuNh70aL3QrHDsCrftX2L/zZq8Vln
UmEMn+gO1aFo5ThKvoE1Zz4F4bKaMWVnRx1ayMIfF8I+bjoLmrFqXY7NiB2X/uY8
cMLhNmCypsuhV5G047fUj+SJF+iU0Wgh/CWD4UDVtMQGTQ/wn8T8UJBpFMrCJxcL
Y9BudA0Lw/pMjGMmV+KvVhY2xOtWgm3JORHqlgkDwsdYRD4CrXEytsj7laXI+BdE
NG9134zW/VruDwOzQHNgX6oF0tslVL9d9LB3lxbOUZe2xXl6noBiLym3+kPSXjgB
m/yJL2/teJQaEng8LqWk1hUKZWVDVl74dMGiK0QbjcmNUJDcWnD1E+HplOfSoX/i
OEIwj2JQ3XHcKjB057kz0TqHHTwL/q0ndd0Ia/3VtzlQ8de3le/okQsPytZmLnT3
g9NaS/TXgh/tqwd8PshnBR0sb06amqbXOenHQpuPHZJDlIEKGL1awNIbNfdeVGKz
t8Mv1fXwvH22CWO0mdUvBR/RU0874jxONLiVKytZ2Dp+5fW0X1Mai8XyF4ENfMUp
2ErCc4/gWMQVlzMkkIvH3YPYt0UiqPcR6OWhmUiuZ0W9GcvaLx9QOfV9c1rNRg4B
t+mjtbMkG5TGDwt91BoRqNZ1kuLwmgkA43eMU3yKY4vOivvi/N51+MZAWtUj+nHx
FlbZ2YE/PYuIP3OtBmnUWt13G1jaX/5f2A9cIHH/uhOcs2wKNLl/LvrnoDSi6VIZ
5eMd/b8oMj5gDoUjCA1EUfV5Xjri4mUYJr77IBEsOB6G38LP69UpHan1CK7EyOGo
SnQm5tGH1VIhtvhBnHR1Gm6aRvG9fZETRZ5s++yR4CV+7VxV20deZ3aZM5Qif8pB
2LJpoRgziWWNlCq42slAenR79Jkjrin4KJIw0p4zWIoKDgjhVhYhRXYosQLaO7/z
NuC6mVvyhijNEhbKTDI4t3v9WjDjD+wOSnIGZwBQmoNimxK8wxyhT9dowPekfI4y
DDXBF2xJmXNJVwWOaUAHl2qZU9bce9FSrdF41ID3GDFSOo6aEG6tLcXpJAfS73X0
R7lXiGo1Ellh5xGlxs+HNLby97+vK32JngkQRPAsPrMh3buznjJQ0/hDgGiiXF/4
MFlkomtVdZCAaM8f3E95I9XDv9H6/MNp8lcbcOvt0OzYNGHXcfYktciz5iBDvORG
7LpxQlv82n8QNvvyiNFHKjsPX2AOBOM26YMDI/4Xx4oh98jvpfSeqkh9lirequQk
yem0nZB53Ghmmsl+1XnS3GphMVAg8NQMxJIeM+MLCQUVvXhi4QJT6WgPLjn4rnHQ
5EOjxVaqpx8yBD+tD5iacaW+c3fS86qBPy4ha2tjrgf8kDr1CRVSY2c/HabgKW/u
ZPIt6FR03KLnJ1hGXsR4DEcnb7ioi0xZzq3P+L3tuFrlVKzZYzyyhap5GQyc3QV3
3U/+McOXzJIM76k8V0AuTKosYE9lyq+A36AKm+mBVclyjGzcNxG8uU2Kg7QdaHWd
1qyBIUj9/N5tYAoXPuw8ma0hfl90CdZkXwkQdFPeBA1JR9uWpHUJwchk0NUtH2W+
C3xB0G+bCp0YqCItU7On+5wXAGp4ikVzCzX6OajWpJvnp1OIyNWWIBQn6ycT6wwL
LxQRPUztdKEmJPvE9gvgS4Iu6T32nfl7LlR8xc6jfp65TcIvd+dk0nUSXh+VEtkW
1kPuGoniLKm6lrepXhZYGKSH80zRK9qok5f7dycWJ4Gu72PpZX/tWYb0Inmg7qGd
UBclPtj75odhfT5sW3RtmAu7aAcDfTLY2eshHdWDkaQIk07ALLQYQELAjquut264
AOsvw4Dfkm0l+Cg+wl7YbjhqojqtHSSis6Lk+UjEzqlO/qRQTJPzj1LeE+o/NzTR
uWLwcvAC8tVtlARUq7x3NbNBA4zRFO8KkcbDPP1F23HxzMgQHB9J79NolwVJecVA
QS6GsC2sxe/E1YjHpK42IDK32q6cgMDuRQDNCh+SxmU5r+ju/ffVz15LxcRGwMxY
qOvGHyAHKZaFA4JNsx1laNLvVHpg8A3FQjxr/1Q9EeR76yjReGSX1hr1B4imz2cU
AZDQ/QF1NZNoB4/jQkS/BVGQ0fwbZOf/IoBel24+8J5CSnIrovH7mBMq2WHAgYoU
AaD5W6fXLsf4j26DbMyxJaVeCMetJ7n9HlQYhAjiPSuVtt+XSsFglnc8RdzilE9x
Ilu1uYXqtdz4s4OUEz9NWl9N8PKMVGDWIVedkBX0IlnbvOA1NRBoY9SbYQ3XPnVB
QMrMYhEHekkSxhlGhVVFgunx6wt27Gj9ctuujPL5ZlA5AvgslNpg2XHiKPjC1ngo
jjZVj+heTht1FZHrNUuIzWsNjgncDJQ01AYhpHgvdQ8+40YfU3ymZMw4m+Yvbr4S
MvRlqAOaVg5xTx0DPpQxlyzwPDxnsgh7OHTMwFxzZvfz4AR5Vvlnrc6oI4QZ1zO6
Nh1REDntHKTn0oh5sFP0Mwr7leVJdOUAhv5ECBOBy2EZurGbi8i/olRawMFJSYSD
9fpqUFohSoVL/7/cOc3ZY5+2YXlgbXwLXbfdrvID4Khbn1oVaj7WeE3OO4RqjO/c
P3O1DlTy4GZ5Lq5DVMlm4YcT3gaulxFl7MftWYBqKC4uKTCyTu0uqfOSixHOd5zE
3QXNUTo5Y1ILGBplO8/59Mtnur1RThjKDZGqRTZDabUcmeuJPKTlv4UJ+fiAUlpg
KvO+Nr6rFz1MJRLdT07JFiIrEjkqxKV7tD8CPwQQQgIQ+VMfbDW5cdvoj+ZWVidK
jj7tgLwRUMEhQ9/J6Zwsh/lhynnNw4H+OoZHLKNgRd08jY1ROOZWB9VHZL7fM6V+
a3qAwhxgiKoQM2S0pPGLoBjU/LlMpHy/vbsx3n4qfussEgJXWqCz8CeI584LoWwk
wB5nFOr++3SGzgmRS6Tjz65XwLWVqquzySACvzhS/AosY480hREV0+NlmUCKWdE4
iIX0Va8/tfIm57kuj3lSCsIWbG3K8ZPJQBb3hf2ptB/jci5bnFS4g2riRxKDfTmP
6QZanWUsT1J2B40kIvbl3iTpjXrdWGeszCY3rYF4FuBCby+5BwIsibvMDH8U3yGd
gQaCeGf95aqXT2oa4Z2F941lh2IO9kwhwvsEMZnBHVoFmHLSs3+mC5siBNLRIGm3
hIuSFbpEHzzTDNDy7ofZFcfCVkzBGDvt9R9O823SnRJlxtYM7XJCWS8X/QEguKo/
Uzaotuxu9Ci2v9RKuLWmbXzAjZCq/fXFj5YVq8ab7XHMjckMvhPK9VnO49saLhvD
aI27/e7OnBkdMS9lZSeDFg//14w1qgtw4RTkO9CX4lGFrIdaBYRtozmPGU5Xx09l
pL1o/lnQh7grPvTG/YUIyeElLKIn+GSvX+Y+ciMJzLa8BstcbeO7ti2iAspyRA4d
YklUzTyeI1tSZ1eEKy4MTRANTmjaFHJCHlDeHTnlau68rFSjry+MevgOlheGN7jA
lyucShSpWWGr+JhKZ7ZQbKl3SeScxdorKp/VFBBf2Z+t5ryw7j9ZIwfAxHfyNEKe
a7rzWfqyIBFKtUjU7n0UJ6VSVE0Y8o2+ZImwPiVo/qIkOGgpDha51yUcLnkBJOZi
p+Ao1+mCx0yWzkukuGdPF0X0GLJPxLovXE7WIlYjzlM+2EciYR+0ZgEygFx4eX3U
tdeQ/EHtL6+Lcq0RMtWu4nfMDbkwMur1jDVLZcl9v9VIk9omg15vrDTG9Xx/Ut6t
+3aaEiwMLMlWeF6PjhWFtRgdnmpB48ciYNlTw+7LZPic0U7OHiDWB4171fohZtWz
9RDb8/eeIbtOa/cOPyS2ASQjqvQArPA0SMLOfPu4ipk5JO1boMuksZMkv7/43LD6
HYXdPzfWdNpQVybc9/2IRHLB9JhC3vp/EYAALP4ls28g5YVAls9aY3dQTXqoLYi2
yPFRon6G9c3HdTMLKMMMfKj6A9oVI8gcm+0ltwuJ4BNKd8NzHH+KoOnbwvpQy4u0
LCB76Ll/KSXcFoaV3dR/G+9XmYHDzd1d37hy/fgrM9jNFJAQ8RzPW0dmetHQdFgx
U+XcAMTv/FDvTlKyDtGOL6RoJ0+GAjMQpe+zbw7dVDze/tf89WXlQbRyF3bfh793
6E5hKj2EEmTdUYqgsB3Pj46oM8cVUymcyqgCC6xH1fYIA+F6NicMpeNvf4008J/+
XiSJR8rXPrD889+rD84WoagVowcag8F1ULabj5xvD47ADVYPJJymb5eftZnJHlY8
zHk7XFbUaiQndIMxWEVcHF3wTA/IiuF4d3A3r4XsPfU4EaBBjKGEwk1m0pJWYSKR
CigAyU5MK2PxBPDk0Pll+VfHuntuSeULq2HJLM/Le265IFPmeyrDwKnmFkhf3EK2
YYaK1qrwFetMP8GKqpFrkdd+zKlKxZbsExWVSq5b+6A3JseX6CQxsWoG8LYxm8Km
+OysamY1SMlGN9VIth1s2EzkbGjQ6zBq3nDSxJ4wlvsJId78b+9OWShkpX5vYPwI
8qZowXj89KsgfNxK/gqFYmv5TAYya4S1/TQ3ozGeqI37kPSNLO/KjGTO6E+ti/5w
TWAl6NtcgnzDuTkRT/1BWs0uh5EoMFcgP4Qd5QCH3U96s5dGG7GF9Y6XdsP7YOtb
MJlV/aZEEtl82v68Fq4SmeGvjBFKOOF3xeaviIQSUA90R3ST2/cKuuyZUoFYLnp7
gsU1YQkcdkHLaj2q/VzsJ7C9G04Ee5ZV562sSmquO3mfujq77YLjI0enwch7l3kI
3+Prj+KUS/9YNIMdZctsRbTkwatVbp2cQZ66BwnpqWNut4zl0zJRZU6KGenIoGDS
xIzKpLQZNS5bYTHPXC4yUMAgbrYtEiGqQATQgvhXsvSmdUOaaxyUeFSILyXIgqJ5
HxSIPBkv9/mZd6iw603GfRkP3JsDfg5p8lRk9V5NSYD4DdJKB791NlrILHUMIQZ3
otXKW4MirhrgbkSjfxWnCG8NUjcbtzNlqlqbf1vmnrXCBFadxcL0Aze2fMG+NUW2
x8pNI7qz8fTvGU20d/gvZQL3eT5LQHcCcSmITP/nK9yMh7xhE1Hol0xLJ2Lg1woS
9snQ5CZNT2dK0VLkiW/Sg8R19ZeQYYyoZg/QjNn8CImWnhkCO4yB1yLnXyf1X2OM
i8azTJ2ykcZANuwzmDdKbl7GNFg3QHp3GLdDmwzKgC1FPSJIN1fqknUdAobisFlh
sxImitPpnEcvVAkaCxvStkzN0Wvr44NbZ3jgvH3beS3f7UcUmi+BaEaatdfIW7nP
NC7ThWMclX6bnQXZ6i33gBaKfdfYceKT1+hUp8uL/qtt9qBSedtPnBf5zNjCPxxT
/lPEFsOu1c94uBxTbiWE56+FJLEHyyB2nnJyPDRBNHds8bwCtJAgTpKawuHnd8jz
MfMS6YKsaRnawTae5dkrRNBjb0Z0uy6CXcV58OA44itdzeYdI47v/L/ujVRkESld
TEvdo1wDjO9DljR0eGVabnZuIdmHEOXm+sosv8HTZ+gDUeCpCwhxyrlJQPFGQGok
sUMw4Szq4AcqkDKc+Bmxw/qHv4EDZgX+UGuOh7NVg7WZ3jebvFiY6boI70RS0Tul
0ogJezPRkSqFhq+TOQ54btyfvqRc4hRWjJ36nRJZW0xrzqXsDoYnaGEA0QdqGucz
e4Ybne8usOqSF6snFcMMWkg1VENp7coP5x3EtafUpVbrpzCmqkVeMkq3EMNnNb09
S9O8nMYaSVUEZVH5AP0U1pzDuAi/5h5CoNTJHT0gc0o/5pRrHDvAJIf+CPmZnWez
fA9a0zoruSKPfpeCYmwrb1/B8LLq41fFKHioT/o6socbmUAK4g4MyR9/eQ+31Jlx
CL6v/kG6BX38K0jo+XiTxWle585zb1ti6SB/qbd6L1+c02hwjO0haEZ0QAfq6NDT
p9kIPtzW7As01ZcND4vM5QOn34sYUUYpqVWpV4rxJinZIv+w99qZk8GlYjkdXnsz
CfAIBz+/NTfo8cecrFzAZ2IM2OaWgpqGBc8gS6TKu41iRhi13VVwmMjFEuvWrjXR
6W6SqghXrAqX6wl/v1g4QyhwYDRULir7l6H06BzYUUenveknHvyH7po3RP7G71p9
PiTXo2Lj33COxLEsAPdQd6P6i/cMrhw3/p/4f/A6rEQ/usvBspcKBKg6mQpYEj4p
66RCbbtW/tSzNFlOwq9FuDdDRAudG+kefP+mm/WNsROBQ7SkrNOCp1iq8z7hb3tH
5/q27M9ToNon+ur0Ti9/R43cupWWHhbGd2B38zS8VvPzcYHxRrKywNvds1HONuHj
D3f/56pNKtTflzMQ1xQ4VTYVpDzcMyPonkQ8/3wt0eDtbthHawhGNaSME+NoSdjp
QJgQgWQ5jkWB6Pzicub9U4ilsnwDWpw00k4mJRkh3h4G/nsiklkzcTOlUjVjlVyH
8YzP6h5ZoYtI1W4cV4dyGdd0+/7Tji3ppk0ehyKUUEVA5/SfFmgTTA5v362tIPef
wM9PWWd0t/YnxxTlQ+VaY+wMKBYH2PdovUMtrnQj2yqpSoqilvcmmEZPJfNBnyO2
s+IZK223Ksm7M/caTP3xhuSmjJXF46m9mWbpxs6712GapqexSjem67UTI8zqn9cw
AhLfKy1MoChJJ1gpkrwGvAIIkj30iaX6iGF2TqVuYTcm/9i9KDuPVKgZelC1cUc1
LxLnDQFYLsYiGpabUmNDtc6CxOBeR/PGRZkPzEXgwxM=
`protect END_PROTECTED
