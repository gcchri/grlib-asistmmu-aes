`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R2XJ4IoW+GZv/5+OcENJY3/ReUOxDun5b2yd+wgDceg+64PGORrDhvwtO6NAHpdI
90V5ixFtRz1vA/lUSvPiwS4+KpsuvGal/WW45gOwJcqb+e4P6joShL+h79wroadL
pw7X7ImAAZT4DPqc2leIC9N29pNM35LZ6FqgVBrHPAMcQJKLSfDSATzd6enStSbb
MRqsCakw3j3HcQ9TNCPWEtONkow1VFETZNu8CcThVxbIrJLSIn6uGnbfG7WHUMN3
vejZ8KN+Kb62P9nDUCw8HQJH1LgIWknX4SoMknUcAduxEAnQ4thA4roWyjUE1HzA
VOCDcC0gwhNr4R/SzJNkCoUZld7OeQANWlR3Kn7eVSCNC6O/7Z+UC71Wml91IekF
fDMbqg/auu6jFvgliGCQOfDTN7x4pDIR4NKqPrit2pwbGqU8Sx3rOYe+dKD999x6
mx8S+njhGWtdSzqxrkFIT+WbczwrLeh0C92MtJBlhbY3m7SR3UNHMLoZbvg8sGpe
pN5Jh+osUuKn2ruA8QZPUdnVZ65sRLWXZpHeYPygEuOOQp6UdIDFuHR/H03aRPI5
MiUwX8ISaRTJ6B4NWrjB2ErOlnerG+c86/LDlqzrgqzTM2k0v3WmX9zx9Gj3gM1Q
u7k05BIT1bGlxcDHLP++G6bil8NAg1kgHFZ5A51Hl9DoA28DFO4gFB/e5B21yIx6
st6oss653bXf0dDlWXoBK6M0CAZ1sC69gm1c8lvyHrjB4yHCDm8mbndLo87MmXhb
0rJy+PSWMjcmJjSuc9CIFiQJyN5bd1rFS8RzukZ6qifIqDL1RYAAkXVpeiuDf5u0
heYsdtsxUjkj02mydzllxIt+b49MKEYJ1iJKOkk18GP3ZpsIpx0iyfHrWFGFpJHo
W+pgKQ/EKkIwry6QXiovTB2yuOJfBS5sxc2jCtj8LHq5Bd3VMKEZ3rQ0Db/ZugK/
RTc/nd4g4Okd1GM9gOzPkfg7rEvt2gxDG9J/Jr3TFmHIWeKdwAtAZW494VSWZRV1
6YA3C2aSnThhA/AN3sTi6lIHyMMjBa3l1a9YRpLNsBwM/2ii0nE6GDaI/ll7Q8gp
egz5BPMSACSfifIJxVuX3NqpRSJqOSH2sLqwHGcHth0gxX15EUB/jRe+nQ4ogDAz
hDe9y5PK9LAdrXbhLVbVI0JT0Nj48CUTSJ5eIWRoEnKFNiSIZtX/tz9Rt1ar1beR
VX+E4vYD5gwNEVIZ6gbSndcU2jZD9nIx3BVdGAN/KU4RzDpQAsr1sbG6SLRjO8f+
GRfsSZ5d4MAMadoj0OyJDZnXiPec9hXcc1GoAAzGOpHFmQq56GUgzcdpqfZw9S2t
U3s0RPlOgVoOAgqbtamtvTZUXwWymRpsG6y7ge2P+N/2rpplSOori3W2K0piBIdh
VqFjScPxfJd6gu7PZyh3DK2EVvBNcIbAA5DLM4jV2MeHJodUW3B/++I+uWQeGzwh
K45pK9WH3ecsTIyRi6nzDjkbVRh0glslboMHcFuP8+3cjW9Ey9rEH0vgNkzPMnKp
x2plHxVTdHIVdRfoEa6AYd94O7+8ja5yI88AmJry6H84+mBFlyo1ai4/RHodinVf
5IdD2gxFOnxBGvm2xYe2voxyBA9SfL8BwvKcJD9SvQ4+vpDFc5KzJ2bCwGMiFyig
l/5OePnfQd7HJokk3Yw/nIoAtmXPJOMc4GQujJmh/6kPQjdHLwf1ArxZn0j0JR1l
HnZqOpG7g2xcoMkL00/ZyD/r4UUzbmCukdcTAd7j1hBcpchfLDN6L1M5+3lrmn5l
sD2Fp4ja/PX5ixfAM2K2KWbZAyK4BvBjmH+OqC2c7cOtUWR2I7kG49cGhDB3jX3L
gqY0pfgXFLvlUicvTxOtBA99aC7JVnhHZQYjB8jES2Kj6dI0jyFzYJvjqvtRzqv5
y+pJmNLVL9FDYtw2AzbEo0pHRzX3VuFDVPXZ5sM9GfujvpAdRMtpIcPvqN8vsbfO
CFPHCcboYJzuBsmLewosStPRDLR6P3KbPOhsEpfeqAxBKZER5aTJhE5rikrWsYfN
LULhhBFKYKJD1Xbifyjutynh70+My2zW4gqZgBwK67B/srONULVMoo8FQFrRJiiD
kLdHgQo+qsLzM9qbOFG6qR3UlVGUPXa5cnEEiRW0dbz6wo1j/75j/Wn6IXDI0QBx
NuMfwvs3rxJmOvdM+DflRsQVYDG44qXYdlgtxZjtKqU05fbKS6mbWp2FQh9uEJ/f
ESyrSqXFB8+BlV9D+2rkSN4creu6Aj1hJJ2pZl2QZTueSmzEeHjbG74HmWuM8M5a
DmsXesKFw49veWfoLqvTrf6lngj8ikRqOaKtFWQU4CyIptItqaGysTAXiInIWi2G
neH3PyB9vJWoucHdCuu/rSbKT9TrkEXw0HqQF2z+vEXElmcjUI0rdHuKUNjvkeUp
cCp2v+aiZkr0CkFeHyesHvvwHjfBPa7R+m6+zVEBSCGooDYX+aChTGiCZLX8clTH
eSg37I+spS/EaPVog7pgZF8M/cNV5945gFs/0ZSry7MXyIA3oUJrzPHmMepwDVx/
f/CgLUVupYEZ/UBm8In5DThsH5KeWNHbC9IxBFW8iCwTgq1nUEkanGDAFFeUQA0C
P7QLbYZSTm948dYYD7gncgXqpob+4YuDzEvr3ub9SCP4rqQ0uQkY3geI9MzuO3Ix
pL/K7cEgpuxYHkGvrO5dy2NLBExGqe7VahgUlfWpimfskljJcjVtfZtihV17HVcG
2XU36CP7LB1xYUAtJoXj/UQzkHCAmGpm+XzEpWdt6tjm/Ctf5+LuA7OV18JO+qmY
lqeDDWxBvxJr4SzVUQ1lp41sHnUrwUSE6O2SBiVtyEO+DN67NkI7Jn3Hl9ZNmrYK
uXaTe/Z9HO1x3vPjmGCpqOF7jUJiEdO/lR3Ex4AhyZoIaMSxGC2LATspD+GCKF37
6aGgczvZ3c3Vb7/rNkGm4AoGCDAHiXYacZdCIOzTBikRuCeZ/T3JQ0urWK6BViFK
+VLG2FEXVzBcJewcJ7Fs7m3J0HkvTUmC7YuMxV85ZvLtyBZVGu5pAg+jhN9f54Xg
lTBzoSHTZiwniIbd6Dh5Ml0b/54psP8kPDOVKpjgqFJ8rN0qV2U1EnhTZX50qU8I
wJh2iVHuIjODYrOK5OiRpThgZruK/V1GsF62dk/WXiDndhzj9ysOsrB8vh5mSyjv
QmZPDUIR4SlqjvgHAaDLDkd0msgXAnzyDJnT+MWQ19oyQ85JOaCS6ZhWPs0pl35o
N+IXDpItoPWv3vTn9pG35eAsD27qDH976eqFDbz3i9XYURbMY2/ENDUQZexbuF/o
hZ8T6tveBw93k2bDCa0szpkoN6tezMM3Wf3LXBZYIP24A7hP7tGZoJ/BX0hS920L
kRiINmHHeykP3QctwAWAwtIfXhfYG5lW//YnBWGqYBg9LR2E/udHV2fkmOcitcHL
bMarWow6uAiU0jfpVQWEIrNSKrTHi6Ar4i40TsCB/I84AxK+0JCr/1QcgMe4M1wz
E7tvFRQeUNOvyempB6aXSUKOcK9J1rvmKCfrurbYeJrio2bVaayhPCZeRCch/3nr
BAT9+ounqBwIrNZ7Q4XpzV159pbGp3ZztiatNtrFMPYi2ob/0B26i6185f2Ajw4x
2PwAZ2xKJS3wGMhbLtXs9Tnn46F4XJl6ez2qz3vZkBYFwwjHwvyGYzwY+WlPDVs5
ywVwvxi6CJ9JmzMB8Po1vDz/x915+t+i9KT35HF85XNGV0Q2IPV8x4ntUgyRgdWh
pGANNZBcGO1+umHGN+htiy/iQyoaBaxc41oaSXjgfnMkZFKCbtkWEBncGaihPGzT
xx5ogavUfXmhGMZlW4ZN4HkAsduZGNBHpA9Dda4tx6pHaYKnb35gWtZho/wcrXeG
lA2hw97oObsAwF8CUFK4v1hc3GbYxhJKd5+49MJHNOG4z1X9erK0SBrR3u4F6LXU
gmJ54d3kuWXRxcscBqG8XpXA9sq7c7r3pJphJuxgRYSiJ4EA4D/Z5Q5xrINAC3TU
vVs7qzkNf6kxfSv3s1E0JVDMVTVzlu5NkTQZiUFwpcufXCtx8ToCtRwUaXwCLVWx
UvMNZrGp6AirdNCLsxA6onN0uyHMPBP1cQbpRah7F7zCD0XiGHnOhHtEn+iV0SLL
lbhemT7X64f9IhWj31vNBuDrfRiVvqHyrlTcycPbqLKWJeVq4yASe23C5UCF0mF1
ftQ+msinHDZc9nS2XXHNm6St580F3S8QZvhi5ENOxvD4UvkfENH875S9+gVXk1dA
ya1Ky4I9Aph+IzTw9hVwsnEM6PKRpfLfA3iPU3wBTOq5L5BvnkgCZ1TBvVvTrXgU
Vam1cWu1BNMtTwuisxfwital0/FsOM6Wz9od8oXkk9cwwUE0dtl5tHX8pbijg7zS
eAFA7cMmXAFSmrtP4qxxAXas/pQ+2cAQKzPlwSlErY7q1xVix0+UyIFrW9qPNVgl
unoQoi4SbjfeT13CmAJYMmo0o2l1N0xOXxV2Qc1+7xQxdxiPKfa9NnY/AaZUNXsT
K1mBzcBkT2Ex6AYrJZFVglyUTO/NBFFtuxrrlNy6lK0tc+RbT02FaNgBieUkNjHM
9ozBKp0dmV20Isf8GXQIX49wIxOeZobFejFQlnkUAMUkHAXAt/XNnZ392Tdv1MtJ
sfs17oQmS1zRna/eKU+e+WnGoyWAjtpMqFYuCfLh7QOI3uysTmKKzeuoCAxuNXod
NIs0eYhjl5Hu5tLBYkaW6qyIKO/h07BIdbzsn/ceRxwbgT8Rttu7FL6dTC+WV09X
yqHifobULRfrk7vtfP0fBtBt4kcZJ3qyjrmX78pXWqE7pNZ2qiRKgmL5cIfAPhUb
uG+9eJ1M1GMsta/h7eqY4yO4WjjbkEF4NU9jXI9CQ1tSuxkLWUWDTrKEPJfBzdzI
4fVj4Lc1Xy09UVdSADhp4X1Wn0ax/eWkoqMCiaknbNBl4UahUHULd0fGG+UEAsWM
QnLZyhBMLquQnpOSF+pEI7SuhFqC9u1P1INkd/nKOy4fmC6Vx1mgZVJ9aRED/yAq
4eWqtlEilbzsg/tU87QHGIXqpzGsywL3lGL1qmDs3vqutCDJGRobhac2WGIHUQXx
KMqvP8qG7UGdgDJOS9AH91KvEDuRNb57Vut1RXt1ppzcJsB/hiakDEGi4NGcLkzN
owWx3Q8C3naZr3n02Enu3ixTb6fu2AZDFNg8LiS0Jc5XidHccLuclmzYA0+n0Cpi
tbEyivkjMMAWjvNFqVXQ8iGZ16MmKwThoAkrkvzcMfaYX9WaJ6Nl8aUrr5joKD+K
6RKDqWWykSL9nnhEsHojb9v2MHpDuq4W8faJAgkfPwi04UVhfBGt3np9RxtFr14j
jcjN/J2hi/nn1k5PM/wpcVc4i6FoAL5/ks4uEcm3RJj1T27HneOlMEoTAeEjNe2a
DCyNvW00WsHUIwtyH1qjQIHpeWkk2qRcqx2tRDC2XqMlbAvGhzrPLPemBPJN/xxF
RO/BDV8xMj4haFxZNXDDqtd42QIdNhJwJJ+XIAOwnpBeWrv2QwbWkx6JuGScG+7d
P070Z8Osmb0UTGm4yDmgXJX+0jk3O9ouSXtRaJpCcOq48ZbI9YoNcoTdx6BZLW1N
CAmnyO/Vd7niM3lbHHRyuVZ1t9YSHDVHw2dU5H+8k+z6EhqON1Ej73Y1XWbXGyyu
SpocTnxpGV0N+wUnU4wxTMaoRD0czqUVyX6GIXNTXdIaMwmBJwYmhTv7VT67uYWD
FAJugplP2MiDMke/pIcGpNCr6L6csgBKqhgjCZKOPahrk/rpNTH76JM4DJP2AbhA
omLJ7TTI0VwvZA6JEOPmmBQBqEjVqwPN8rpgGRl6qE7Eum57VfBfH5UmxE/ANC+c
F5O6jK7t/ehaHLChCE+rqFQ8LIarZ2p2H5CiTGgbk1MHuihhWjZQmoOGLwpoQl3Z
DTMx8ZFCl2R20jYyAQOz94Gdu9/ezVX7hrMRncrAtx1ZfTCmtEVuV73mddi697xw
wqPu3p0IkpbisZMr3w0XbWZMMGvwpVkBp8DfxSf6/keNEAKyjea9gnFvtgBSg60T
Gf8a8QAIWXuzcbEzV9Hwnndbpo1mfoTw37zePmjx7M0WkIBCOKzaNIQxKnGw/Vfq
Tfi0VfUrw/vH4ml/uGvyeYGujv/P5nvq5azisNiCYlxQC4tc6TePUp9xr6F9GI1v
lWF4Ad6Br1mrNx8dV5B/YG8xJ6J7gz6ygCRuS0koGUs4WlKiz85m/PBjwvigSkKV
UZKMrK/x9KjI4Yww0cxIElu2qLP+DwqSd/8Nld54oiRgSCIHl1vCtnYXLM2xBjla
QvKTKuFOciT+nf1GVVzArdXKQwdBxxPW9FshSX0BcRtYRkv+XANBPpgWD4o8ybAe
FvoroHNqLf0O3lnettuhrqFMAssFJnqZqrJK5mAdzCVktmsgwpUBQ/WJ73hLBkX7
RkYfR4JFHz7ESqvnQPrBefKoWNEFYsSpVU1rfGNnFvyuXxpNKkOg09ky7Ex2i/HE
yJWEmqePkicOBHVqW6r//LpB2Fiz4dfi7ZohGrFjjcRWkt+Xr+l3jA2/YU/g8Lva
NdpxIbam5cCcef2V6FJfIq7DOcWQpmAdWng4/mCDTyGaku4hppRDmm+IpyrZ55nJ
urHhKp9Mfo3TQp7d4TnOim3rxehSimGm8FUqgyAcawmd4EyrxNAp2dEpe/v6upQa
rDVFiXszVNVDkoBUnADXGfbicWWiZ5+czuIuMehIgY2wXAfmytPaFzQ+3LDS3Hym
UnClVY4FkposTmjqQkAwm/aOur1aubwzjIVWe/syU+w9P/KPaqzQUHhXiVt5qgKd
TAUQtWfFa1+XR+/gJa2gWFos4BJXrYqGZVZDYbSDY7Ar3JeZj2Z//B0qX7PL/KEA
qdDvsqsMKOhmFeybOR73J+aIaLP9NZuN/mMZTCgkAhFNe3jhNl/m7V2C7a7bMMUi
cLtKoiMDzZLAz+mihg1Ffrly45ftJLg3ijBu1d3ZBwvCVxxKNl4huNweRS83BWPS
dGXqI35vECpPjrVccvlPyMiUho+fBdt8nWEmFzY0TgrvBn+09Xb9wsRharX8mICl
aGStV7MLK109cqNTJ7zMFhlGlc0WLdwX9YhMPe4z2+XCWC6X/zWX0OztfNdltySR
CDeXa/VLU29bkbBnkBuExVu/o2s6d62AkZHDNueGU/tbUbz+eLKbKgtc+EzF4YpY
ZsPUem7KFUxcizyE1xI+GOuTUPr9xNV3XC0IUDXEh1OdSPW7yuy2y9WxIfDlmVl3
kGxB5NyQ/dzjPCYjytyOxgKqi4EwHJcaeu0mKpTu56sB8Sk6Z95cQJAZ8kt4f1VV
x9wupLJHlza0wfP/DtdoaVk/BHSEx4NgvtaXCBq9LOjQnCjztWJwE5vInbLj2mkh
JaQ1YMTPg/b9TDAIdR+fG25umzK61YRj1dO6hGkehM27B7Ck+fLgIpeXPkQBkf99
nGSE1tOkgeJbT9mIJiEtusNfAnsa9YtT/yjm9JnYL9MYNs9CuUk27uJrzkJn6htj
eJQdThOc8RHZchRsVo+XNLQvuDhAEjzJT3B8lhBMHIUukPql3RiiD2m/3yQgM8YY
S/TUJonTfEC7X2dv0/PiTVQe2gddfgG3fy/BHylhaAsxKO9XQGwdcqASaEed2gb0
4aNiOM7BtQnoOBWmRF6DYIN8h7kjWD53ZhVe/6ET0kToCUe8KRfEwg+nghDALqNr
7ZsQy+EdYuicTmiidzDREDyfuihtq2L9jBjRX/k2ts3toz8rfckegJTEU7J9zmVE
FPYT4X4IcxpdAU0DuZ79n5EisWuG9Tvqoedt7GkqOtOfYcOF3s35HibPzy67QTwM
nkuO3V0UYNrVUH/d2u7w7SCxHZRShaPHGEf6pkQazE3WxauJ3yCM9eI/c3iv16Uf
cRQmwfGlS+9tMQLrhUYLVkvoHBTTnpOYYu86djlG1+fe0bKm0nfXhSwuDzI5HXqN
6OV+hSB8yMtw8PeXYPmYzLgeG15bwqGBdVdjt73bYHff27Hh01h2+DLJK3wCrbXw
x3+xo39vG04526tZkBq5ylyvP1EuZ/GnM9FZf3PbvsKJgVqAhrznMfMKTzov6CZc
o+/cDdx4dGkjaC+JFwC8hMnHMK30UDNlQ2HPUitaaIUasKVQwTmZ2urVl3u2nSfy
l5NIGJcQTbHlvPbN22RPwHyZYe9X9Usp0LU20vKtOSS1msO6HBMAdDv+5nMAWBoh
T2+BtpUAAnZ/9PqqYYmg4sEHHbO3L1Sp1HfGgNd/nZ+rs1y7VCVe74+L7iFEqp5s
0MndF9Rf6n/UdYLbs+S0RxlVnpri9SoZoI37/kjuEOo4+wIKFF/EHtjlsdogzPoa
L7FglOcyDdKs8VziuJjMOsUmWNGTr8C2sfHaynjfgOqOhmXwHDZEh4N3axQceLye
IhrnlQyuawU7+aiqfb3ExV9jRxbldqIqE+kYUc2EpehJTLJoJea1FMcznPveDzQS
y4eTB2HXYAumiiihbEjjBf4CbAccH85pMVE787q5zFTxA10j/WOQwDNE5qAlhmTr
l/g+AC1tQsAcUDtlO57SkhBRGlzpOSSlQtsPlnXuEmuhVLHQAb3GKMU4AWzYKuE+
sDwUxB8j0s9JLRPsMhah/olT4X+wh0Knzww1YR19A+uqOi06P3ptmtKQuxYVX3cg
YoG+oSBFq0QX8+6Ypi5sbRBZHUxnhP5BniH1xX8zr7+/ITYkGsuXw57T5P4UI7qx
0hP4mI5Anin3Uyj/4tMW7+5ZMP8tJ45VC0fpop/vuUX8SzZDwLwljhXFysibrnn5
sDQtWQKVqpswd+3K9W8mgsDF0GOjPJgWUfufTKeuj5NJC1L5aDYUhqmWnKTKTKLc
rrRpTpdPDNls7VVlGL3K53r+O5Ggg/ZeLqmYnusUJPHa3xFL6dvi3B59JCVMWBcQ
2f9KivAtu1M7Ak0Nb4yM/dJZPBSFwm6Yk7NT5SBwBJePosqhHymlvPJ4gXSFFmY4
c7TlonCF3pn8NxlR1u4aTiZ4mT2lFPvb2THs0xCUymIYvckN+MLvMiYOW2JeIJqk
MIrnf05PG9crXK5T7HfxWHkB0Si5ztk8g9ipwU6sLCTRHI99KKp/nXUsxulS/sJI
Lma5IX9KihejxMpPIU753Yl6Gy3r/hnCCnTEJpOPZjUxrP02AXKTWPs8SrajeAax
pe137yEXb3IG/PY4SxFwYYiW62Xb6khypFVSremeutRmPWkD4/NF+oOaArqF3SLX
wRQfaHx1syStqZeqnmrR0IYlgip1pnz40ezb01zi5FJrUURtjjLH8mwb0JQBYteQ
AGmH8JdN6WaMmijqIjSyiKI5iR9GneuABJCN5s0cFyVBNXWNAWh5yD30w6XCmX5Z
lIoQ94pMBKQj6pp8ahrQYkuaFePWnRNsoz2kP57b+LU2Ya9VIOopgku/SCEAkxVp
sNf0Ll4Sp+LnsvAEMKaUelEkspW0Yc1ZQqcy/X9yfejJAXEnFUyhX1OcjGfPQLDV
co82uI/pgh/DkRE60QwnlopZ1LL+2pInH2+47xfey/0RYc2G1UqQjhZYExeTo9ok
1Oh6nZuHc28AfEv/Z7oK8ROBeuxKaQex+NbLMgXraFUzUe+6UvSLqoP0eBYsdPZV
AYeX4TRH20bnhbfcW7y+GPS7qzSn5flTO2dlb4lIG89lVBb7SKdOXhWBcvTKcCe9
VGi2ncgPJrLRyJjPXoGqT31BQ8AtOsruTfFLsKAoNmlBtNb12oQTbhN088Cf6pca
jixAZBvYN6CVQMYtir02aouGlYtpFwV3c5rorKVXAbzTG7/fprX7irTohZEJu1sS
ERA0gB0FPHmMtHT86u3k/sunNol7KzbjZRtoAZCly1cIF+FX/qD8rBXbq7yMjCkQ
QHAoNcawQCks5PRjZae1tmqDU9wYsIUpAm2TflbeZ2ESwsReIDcn+ma8L0dxDbyS
4SUNYKu60BQdVyiUrmwo7i8BTGi2z1qRtoCkr0gn9DP2lS3UhQULBFvdNfvUCpsi
673a9jk2z8pt0XDk/iDRFI6Dl8DYnRDw4lSTBHIi71cnFqW2Jm27vaT6NjfcVXjW
GKZnT9v90kc4RW4dnbdWJgjLt4YtKOezTdNByJTnQUuCmxNwI0B8+ogobOt/MOBC
jRQLhkqgg64s0br0LbtfNlpNRDimOLlXzOVp8RUp5k6dCbYCpU3XlIZd8ull0ous
fpHgefM8/WTVIu9IR5uKcOGrXBWT8mfy19ePLg2AxVPqrlrc6pXIyL3BXTnoR2i/
D5syIyD7FfEfbn0L7cxBKZgfrhBEIotZzhOq8ZVG8u/6qPLOMSLMYrixAF5H27YI
NpXRnLHgQ5IKbCnMJpp5DNzHQqszwGkEVCD9IHUtEiYtvXp1nWVkAl2OUDfYHaFa
wU0dTA91qja3bNNbeg6byypZox/vDnTQbsVNuvGfyW07VBiRDJfupic3MjeiJqs4
7VBcqECQECgBxNXvRqI7lv6bRY48PzdpF+77tr09bWS4UMqmI1ItGg22+mlwzTYO
RjHW3zZAB/BL0TblI2Zryk48H+6Bn39rbdH23pTjgvM8xfPvMqPLvi+/Nqy98GGG
blmeHXb5B9ObkghRm+R3o0z3GkNmf4ncal0LVsAjlMB77bxos9v84idHFOdPfQj8
HPRRVSzeGDrhhHIBi9Ao1pdX0NG9bNBzQqyOt+amyXc8Sts29oeYFPJh57Z41L6v
fN+/vriTpj+8b7KJri054kWnbBYOciRn5HVR8sLjfeCQU4wBPXDARAQ1TYjcDd94
jLq/WWZPSRiQppdnl9/Jw3Ft9pCKe7kBvVMl4kPf0o/N7ggaHqbQXOn5CEwYzvyZ
kESCgpnfrzAFGcC4r/K2M1qbdFU30EH5mnCQwmENlTvIX2PrqC6Gxx1kCccQjbEu
mleEFxSB62VqKrTpBW2+fmrTMeI9l9RdosGsBZGXAEWaGizW/w1T60XywZNcEJ1+
7NEBnYghxkKWN26rIWEULhGyebwViCqnZoMhwlnvT5rDEFzu/h57EZHt1RUtfq3z
pEUwG+o0yYbAR9v4u16PNHhJJMAHfj58WIOOPwxBB0t88q4eak+55polppgMXLdi
01iCy5+7fsKnifWUz0xL12a0S7whWaK0qsQq++VF7ye4yewLf3b/S+jMWLzWqROM
iuVIUP1pgr8WdRqxM2jcBY8KZ0kLGpsXpQ0J0RAX/HKR3Wn11llyGTDnO6UcDmL0
YlfMC5ysqaQpL+BML8PK/5PmtQ/GJKutP9jFOlr6hKEJqOuebdk67VVfVuu1BEU/
AlNBq89R4NH0g9/uX2YXe1oTlppLlEsRRQGWNfLy+hxZnIiVBaVOd83Gusdbh22X
4DdS8HiYaBqEOBkybqqzBivItM/4V0ISHytgGiAJNnPTnAsAceqFfre+ue/xrOPV
uJS5/FLvqLbkqPYSb7i1a3GXGYMULr3dMW6u5HFQbqO5/Dipgo8QEQwibC4AXWiQ
SPghxYFhhGi6eI283O2ns3lz3vh6yusnReIjsGr3/+nMNsI9eR/PQn3yVzAxlTgZ
0ug9dken0PrHRSWGBYt+xCazcGK/L6iYJMGbpbmxc3CumgOpe5V3BXjBKBQDhji8
TQQld9/v1hUunEOA7k+kHfXyd1G0bcd1vQ5hHzTVs9d/fvAKk91ovtdDmFjucDoK
1K5rs5zrk32lMEi3FI0y23S+EM+RtatKGWboH6pxhC2m9ZQpqWyy0zztJYLrKdGD
aujTuOnJfDhb0lDpDGuZJPu+uC2+rTHtp4uhBeNvpfOsZHCGZKYEw7Kpjvk05QC5
vUrUaAern0BcXIQWZdD/SLnbE76e/jOt442g03YK2Dl2n9BNRDLQN/Roa/N1hLoL
4rHQe7rCkfdIC3pmeZ7D/35CtAFDWk7E0G7QMsSAO8lwfUymsXlorurYuRrZeh4j
tBU9KG7OW05abPayHD61tsxCqSUK93xnpxLQfhwpsP44S21Ug2nL/931uwDpCfSi
xix6aWiJR6UU5aNNHsa4B7fQG7eaUkSK54kG//hao7C9ikbdEZzQhnSlZQsSeBRr
tHjdej9VVIhYvyHzotXbon0xG1RcBFnTpLrOwIVw6nX2mOLseJD4cgcSJ7TdWJLf
ooFJJSqGGlY0sHbjZg3iRnUBGd+56OX/gob21GAN7PMPRcTqhpMxNU1OM39rgNWw
0vG3/52tFhjY1kQlf6tmvsUrW3/yYQpr2sdAKJmLJ72/j5QkmvNuBdvG5us3pwl4
MFXM6uBfjS++hNVnLz/hWs/VFXk3fXHrUzcoIHPV/WagaRhHqQsT10qv0Tbgmf06
wtw1mJuCRkyXPWt81+fMZw==
`protect END_PROTECTED
