`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W8gUBtQDJmoa68haM7FoQ0jv+ZT7SPhclOSVdvCG17quAcdlMPGHLzUF52pHP4Az
44F1RcRw44bkxq5Dxn+ILDQ8oDeADG9MLGt5UlnsR8QGGxRYjal0eMO8qTqa/0fH
1PMvEjxHuPWkhj7Op8KfbdIZe/a0a1R75t0BFT1whc3wjIc9aA47DA8Gaf2LGTKv
y1i2sVvGnIR/F2b8jW7EYbjcE9jg5JFrhR35wRZetej7ffJB+Gl5RyMGF/Cbve+4
ZpRR3Ds+Pdu+U/762IYo9v6SJzbe3k2VSlCdDAUZVv+FDMuMghLLlZwg5/ScBgdj
bNpml9FJtcFltvLew1Sshp8/15TeZVqDhVQ3pqXZL6I5zXlQYYmJuXQTwNz/oJ2G
J7mjcvm/ogI6J8iTC8tCMFgA85NkjYwVALp/K+iJpniNEhGkdY/F4UJezDs7toY/
54Ky2LJFbp5OELNmnik3JSd5AoKwnZ/NLFGDJVqcgw+cEzA7yXwyDTmSrsqN4lMP
8PiX5bRPdLzXEQcWMpFL70zDwWxFg2O8SOdlsdZxE+QcWgx12sS/H497cncEEHBW
ADfZzVuMJ0i05jmIm/6DlDXJXORP5oKfkRG+Pfu+giWhPPKMJJ5gbQZSRX0oe0r7
0GKLkHLpzUDbAiU3lrpHWy39HlKORMDe3jkNXB5xSFjx/aYbitbUqmRsycpHtL7D
ztdvApiAVC4W1NuEMzAkN+06IbCsEaE2hEg60oNZjAIWY/gcdvML9OQxhradEQIY
Jjek1bH6qfSBpFVGcRs4fAqbQcMcuWfdyC3Aq4v83H8FmfsVN+al39jQXRRamLBl
j0WvnOFNltriwxHWAG8hTFBCtDENTzGvXqQMqqFq002IbXV9tk03pr0pucheS5Tk
tQ0AUXqO6BAN46Giqo3ehIcieWLZhGeYIRE1CvvN+iH4cOkN+ws6yiq7CFgDZFdv
Nw1C7+cUOouLeV3zQ3g7mWbBr6tzW3/ineRUZAbbgsKI+jHrwVT8mgxo4IgIoT3e
s3JRPzJk4TRPoB4DKjjO6LWFBgKMp4Eil5dUJHIuTBnW3PdaL5SyK0/9+8Q81Qit
pLVGZVGuFhAq5TZRaeuilizIuPhV2SZ65ub+gUjqJfcmsfnj0sb1mcbZzRVpRQFa
nBMJ8Z5mNbI41xWXavJ6hWnzGxzhE+J5ei127duSb7rODuxT8yQ9uxUkCdczCuqw
ySNv2Y6JOR8NJNmapNYKkwpi4OoMJMd9+UMNDjGE35H5sTvTMhNZGjSSR/sztvtx
lttuZk72LsQgKHIkA9b9bTR4NFNDZsgEnVrlFerCkqgrlFkQ2RsOGVDuowS8sG8s
tsRH9UL64sLGOOeqpNshvmi+zPCd44E/6dm7izzYb5TBEeZsiIQGhrRmVrBvWuMU
CdZlZpOJeh0u61oCyeaVykZmpsPnql2dUMr9kYS3cGslLWeizXbvoW/Ck1mi836v
5wztZ9AUzbMIpS6inpaRRGvB3qFAVSyW5CTC8t3leZHlx+w8d1FN1mBI4l+gvsJi
uCJzgrhs9RPhFhialATOQg4xTKrkzmm9VHAPYRbI/c+aOYP3TYeyRYOqIhIYySVk
VDcuKASLkqh0QCGIDrLQ78QsncdwZ6wpd5RYrDsOKnVjSdMHyvchPYqcoRpas1rr
nCi8Ru2/38Ct4OXgsDNy4yoW7ZqgPf4JBuJIN0oC6Zs251RqxrKOLBv2l8WcLsoE
Kq7s4cs6fSF3QHwKPkMNWm34aSPYdzlO4+AXFJwkAADFhixhgkSd6GNxgkx0xG91
mA9rBgLzZ51SPK+BBAfweWHdZKgABSRTUDaOGcRbDmcpzrU8+2WNpAf7SHMbUiMM
80vFwJOeOFE5v8xiy2H4lSijd8XU+E39ueYW6T6HpCekx64TavGgwjjlmwc18qLX
s6iGN5ZCGcSSl2hi7twrQqmPUcPgoxYyN4gkuKpxwOUkQnB2UXAm7wmPpBSc562o
J0DHhJ2MyYHg6To1c3z3K6vtujMEYWulkXRSGq++MUgoGuWkI1mZPJe8aZTr3Iiv
FgVk5PHA48Lf3/00JNILOFmb3jx6k+eWzGrOXpgTwHZ/NiiFWJ0ZO0/G5mphhEUn
9J2geQsHE8GA3PxU/6qcCcZwohIkKOr8jvcryygeKNzLVJxRZWDvwooESP8XEO/G
zeKj3HceSMwN0zrq7sD6f8l+8sM/XvZVbau64x3l2JXU32XpcsZmBPed/7Tq2V3Y
uGNiTsEibV1oT4ZZADTcTzrfvlKlKyX1Yq0y7HeFF+bSSCiazrUlNPtp/C47LvSU
b9I6wvtCcHadLTsYEEcLWtou3yEe9lEr59YwzplDVPD8ZBYktVd5+o2yDAuRbQv3
Jb/bWNCty3b6VK5WJoaV8dC80zLFjF4yLD/ENkNPXSkyQIz2dDyQRIdutQa76yXR
+iFdj8Mgai3qZOb3sIA+l4k8IrLzpbRmdKJCvejbkvsdlU1UOzDs34S/bHtL/K9I
iNlXhlF4MSiBUzICPfdXfQYWT6vU+CEriFSimb7hc66J75075jI/T6COJkFNYqwY
HRHJtxUD1UE6UsxFDinl/TTMOJoVV8jqbTtHRhxxG43sF8eFKbUFWxJn9VJ9zd9A
YaHDYEq3B1Od9Cr2XrqPU5npBz92X7+PwY4Hf004iMckDDuV55r89RtROFtJQPmI
XF+njnT2v3rB5j1tTgW+puWmBD2xoQbtlw7UJOEjeCAJ5/WexTuhJwCgdCQ4lkqU
R9o5ZrvfkZ+aYoE/B6wMEacNw6qY2K89A1TeyXSDF/5qy8z9irAKD6ScZvRfzIJ0
dV3HnJYPLYwyDQp0WXyE/nkYE730AhhpUYQS2WoV94Ensp56JHX7YFMzn/L+BGeC
1/TODIgbEM3XCzRzh1gFBg66nGnXoLgZQPa4DAApHR5EDNSg46uH4RlsvtSNObs0
eQZL4XbFE8L8+OVhZ4fYLTZNeLJwKWhKLP8IY9AjEC1Pph8HAL0L3LZZX3ujTkCu
uLq2HijXYd2DwZgxJbCjRTddP27CFzdvSdZgoDILoqGEdNoRm9Oy/wTozObY4X9O
xodi1FnbI4Sm0JpZ015FlvVXU4hjAOhuPH9uqVaHTBhEsIwqL3oJGLeHsZAwR2xt
4KCStn9YqIxQ3/ZFb1h6iZjc1BF/8cUTSmIB0jd4VEEh+O2vUeIdqCc/LrRp4Qkc
GDOu747w2/YHnynubLYo0FuU8aEcOnNVoMUaSOu4brdHn30Ch4CrRXb/2ndX/Hu/
P9MhJLxou3sUs6bN40EGRhH1cCpDX8ULIIGmhCJJZM6vLrejk1i1hgxbdBQBZof4
kXHQ7yU+4voi1Xgr+vBM3Cnz0NvQ5KIe8rlxn38Dfkiflif4tSuYM6amjW+gJS+N
0jpBJNABdXMVJ72iXaVpLxbkRYDlbIBtSB9v6zqqAfhlSLZhkvj03O3zDQeVf+Sy
Q7Q03AD9mhGTgbusQbxi09/kAmue7VRgkPJV9sWEIsY=
`protect END_PROTECTED
