`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3ql4kApdGwpjnikQqtYzcxXFdRrYgH5Bwcl/Dd3cd/o1idjOyoeWAAb92Qnyv4oq
2JlKPQ/hllfeQkpyJvf6pLt/6Zy7GWDcYQDch72jnGn5mypC+ZfT0QinCorap9y8
jtuqXvyOs19tmQoVbLQgpA4+qfNe1M86MNTXSPO6/wUsnsPIx+FFNXZ3OtRVxauv
C7Ax7jWEnUp3FhegmF09K29N0mbcoDHgtVy+QoDoS6IpshVjM9zSqvqrHzGqkzXe
ZGsXVmOemedsz1qj9TzAwoGa0YvLMHj3yT08L7Uqc9Jdbgl4wxxdu+7sr8N7/9p3
u3UnYvIgcAWpUzESudqkhvi17SRqrTO3yhgGJ6CaVtxSSZaVHL7BkbHjaAY4rHvR
XvIO5x1k6thzZIAG1NZWJiI7txCTZz825v/LAYVzXP1IrbJdvepHa0kTvVWBU6oK
VGz2v6AIYqpg7rTbDfvdJklOEQ8qPLE76kTcztGmV74upzTkx+eDR7kz/We6RCzZ
Z6s29WpCdd51sYt6LJGDc9kqcz1nQuLlwvKUzyo9+hUIZGRtoOVjXGGKEHtlDz5j
nVLjzqfxfrqmKlvKPcFOOow2lMlUSrqy0lgtMpSK1Di8eu1Ih5S7lSZI3WRv3D0S
sexzeFasDWCBWae5u+3jNihZugocMsvCVIRYgZlaTZcq3Rwy/Vn6UMthJ8TeHgqE
F7z2nSJWfunJ/UjA+OFWPCLXx4p2th7NIpCfKPQwQ7JR9Gs9hIkyXOor9jUz0ura
aIXCxEQbuUmaZWRIXkJOqAl7S2q6HAcZu97EwK+1Is7lWcgt9w8v9sXQ7NnDWkMt
+n3b3lzP4xSfXEEHpOIIpvoDD2/GerSWz4uuZ+WMgOEU+WM+LpcIxbv8tD0ebrR1
kJSTXWIJmwC9fh/DT/kRrNXxq20CemsjD+WyZOryopp3W0gVvE/ciQrQUt5q9e5O
FYWMBYACpgyZUbiZsJ5FLVOsBrEtDLobB50wpE2A8gzcp7d4xUAQkpSzhy1W3FrA
iLSIuSu4ctX9w+cWHqQesJagKIszn/SzUnwngtqgiT7brpSRgDXZIbnaAQ8k5phV
nClYQ34f6+rgX0qqY/o7ohKpswUaF86VbsMFIFCwxn3OadJr30yAfVboRGS4NGtp
X1WS1UJqAD6ZzRKJRHsWHep/z2HuhIg8n67XCRLmkF62ppBsb3BJNw9SiE7Sa1OQ
UXmupMRfLgcsoVskr7HT3vaxDH+d7yMEnstT+EMZHjqHkApY2SkRUsYFI8eHO1MK
ZqMvjoHAhNYjh8+qe/+XlMXkOu9pSgehaIQh3vQoWCpBstyf89D5wvtqHjsw0KLK
ZCVKxHF2JB1/8awm1HGpx/bvxXFu0s7CWUmE/8UvDdO6RqKF2lH47nCH6i8JRXsW
0URJHQgz8rKgpbG2XjYG1g==
`protect END_PROTECTED
