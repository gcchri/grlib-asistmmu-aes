`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OObjO2plpy3av4GMtMM2DD1w2bkPH2Iaibg8ARBJLncbt69/8Msncqg+k2L3tKSk
kMXZixPsk28fNYj8EP3mDES+eSM/cAgKMJUxih+nHlA+qPLc0DU4jH05NLh9aX+d
zIRcex+754WSuxGFh01rsbRmH4wZUFPLYaw2QB0+gQi816bsXGLZ7jfUnBi5106N
rZcnBjSdonlmegPxYUd1RYxK5tP83hRHwD9Gi2FsEDzIINBWyUiaJ5r/l7DfRnzv
VznV4pFt6SlKhmgHXrzRVlLhELCi96PznQHCfeGFIP2VpCLwcvR4JCcXlnjEBPFa
ttavrQJ1hkmZtU+NH0Gbyr64p9xw0IKT4e2OR7jl8tjNdJpvQ+IVS9abQ8kk+GaC
f//+J7vlr4kKR+WB6eLanB9KUrR6LPQpTvTEm0hBuacQnQTWkzD6yQ45YHzbzOsA
MBbrsVVA1BVGNrj7n54W2aOqgG3dOtHmjtMA+HyXv8kKryAGMysdE5UqFO5tu6d0
tRRFIY0wm1wQS2/iXJ+pFQ==
`protect END_PROTECTED
