`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hximl7Da6qiOj7XXFJ516tpHlNb993PDnQlXlMbrZqN3xA/GVFDuyFhpdw90ljWf
u5tgrd2oDSS7t+eDf6s2GjbNRryBHMiXKR82k/ZMRP0Vm2pGVjEkNm2FmuitHJeH
ZwbzcAb/ev6wFA9QLSx2AsE92DM17BpZsCZGskjNNbGTTzX/ViGuQvji5fuBqAzS
QI6elN+O41YA4Fs84JtSuRXZkg427hbJLY3A/N+N0MRULowzrhq5W9Z18IeZduIq
1YWUuB/SlseEA9dNLf35KCwCLaOrSI+VMKCESMgFQEG66tflodhd3bHkmbpHE8hm
tK0sTCgQC/u8RwSXh70ki8SQGb0uUliWcdCBVSppcVr8uNb+VKNuQTXtAE+Q6ush
SDQ0LLNPC5bHp/ogr1JQfD6x85Wc8Dx8AQAPzche6PkSMTRwIp4j6xms+AWNN4IW
qODVT5XkcHq3iMXGB4uMJtMzFphtmxIybVJMxheia1xXOYzIIg7n7+gd420rs0NI
1e3H44g4Vge0gWYBVh1pNvRa0MEqPnttUoFo0CCvXFrI5ronmR8FQToraDehuCuf
n/FxJTZbP0K3Wkhu413ZwX1s9ZTlhSLlH5RnYysTHlk88ncpJHhDcec0mpCNg75h
VfKaOAP0R+e4amVfTnmBve/mOo6Uo6qL9NfRCGQGQ4lQQYApA8U9kF0Q7HVQ7CCe
lfXtWQsOV2foicC3y7LuikdTiYrOyg53bEmhdHEkMKWmQuwvuTZBiDJzpxGeVLR6
2IRQeOWqEySbdhFeMxaBtN/5Wz51LCaXNk/KRC7rBXTYSnCCCFxTQVmbgSnpKO/C
exQt5aKm+EkSm5CnlKFDyk1eZsaR2Yn0cAddB6NygTF2ZhIsNzvjLunrBfR2nORA
Lo8vxyhG/6wssqCiYgjcTEM+R720JJz8be2+KVjbczc5x03Fm5lBO4jdrcUNY6pL
kvIxTDg/VNIbc+PEXKnrbCi4oO3mic4o8OtxjXobTYwo3oH/6FbCBfAa5z2JCQ65
`protect END_PROTECTED
