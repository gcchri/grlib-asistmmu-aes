`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SdJLheJ+KwudhLIuaZttfGbmuOYa0GF18B5LfPwEhOXnVkw1dL0WRgTYycbjfiTD
0iWyijM4l/XzKS9DihiP0pviZ4OLucnQk1lcsYVmOTOYnv22B91qTdbOzxjs9S+T
tFdqz+lexHfchCIvsx2Sd8LeiqVT2SgFJy4WxK/JGmgWVNt+RaURGzgJk0aXfCMZ
HNeMHjWtq89AQvnr5iNvdNyVz9dCFlT8TFYqhV/ektbZtWSoqUjWKnJnXO6uwKGi
4u58g3a811F95U/BSE3aNhCRi/dtGFowF1Q2ds/Mhfh0zoLWG2iG0yIbHO+CIDNk
6yaxKotO1uytpXLueNH/+zhODjdg9g8EaXKUTu13sh6hqxBcQBWBPmrxwkKQq17j
C9njYeWdXjWQp+ClXeNPI24mIEAyANR8ld/C8PyrWbosez18lhDs2ZQXVZfAA8Z5
PdFyCsdajUrUKkSsQm40XCLPOFeHZugJd/JShXYcR4GcePM7XpHeh/7LaL9wKWBU
wKtveufLjfdcO04fV0WzhPRvOf5RKR1Blj8wQdd3NhMNSWlq0R6fOcrG9QRxWwFX
Dw0VJRAM4kxhAZcAeTTAN3y63v3aasQ3H1H9UxL8TO+8AogsTSN+WzicEPY9z/ql
TqAjGg03PcegasubQWjcwP8vuyagYziMGGUC1EZDpHj17/KsEdQMmIvj1clQTiUf
BO3j5dM1dnIfH9N6K2tZ+Oeh/1U1OxYIIsdzDI3tC+U=
`protect END_PROTECTED
