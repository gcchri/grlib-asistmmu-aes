`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/EKD3T5n4oy5V7YVBZAOcECWlWnOjGzfZi8ev47wRyx4w7Cm9zQC/wBEjUhDSEhj
We/KlSbqMb5yWi14PHX1vwk4lJ740RtvP1Hc7SZMpkEKWG9yOwt4W4dq/Ay1JgqE
9bvdfRc6X5S8FJBm9R+1vH/Qt6BlwsBQ2j5lUTP1HMIoVYsy+xR0G0QlMKUeZnzT
BvBK40aVoAOy7+51fKadkSaUVz/wLXYztYgFWB12JU5SPwCUC0yM0BAGp2ZFpmCv
1bptKO2pWizmgdD4Wn344voFyESzyIGG+BjASAWg9lau5d6RiCJf6PGzLKetDqau
75dtdhTkBN3rPDHmvaPWJgExZB/Kw2joqqjJ1ti9uIT3TOX2cN+79nkPOaPcDqyC
hkldkCrXDw4qGKwBeukMUcdKAQKLIO3KjdN7EQ2gR/m719OeWKqPYJVxaLX8KB6W
no95MtX/U8/DWCiVdkmuaTGKtpQU+zLmPSXKd9L4nDrqUMeIWzJeZlok8hZAOfv8
yg/sPWKPuoTqdjEnSTT1rARumGjTysVLLTQ0asKefeU=
`protect END_PROTECTED
