`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WlW7cHA7pIY/sX0Om0Md4zQ6pwRy3E4JOpRREgY90M25xsn7GlCCfM9ElLFZp5lG
orFEyp9pJ8qFgq5c5ZXMngbIS1zjRxSvG9fPHDuoi4zHMbgDO8r/m8UaF0qfInr+
ETt/7YnPWiAMoRDLGIRgI4rbKz/6WR/tnU9CQ0VA28b4cU6zXZULfu4nANTm+gCE
f4+I+OsSJUjoY0Ad5zaMjIEITOyT9Sy6GbKQEEZ/TmLahokM1OizVAjy4dWKhX1X
SJA9RMUxnYkM/g45NpSsel9K+8clQJZ7KrMzJF9hUbV11P0ynZGhDa6ZpdMth0aV
RYEUDI8OiyZH1DmmflemtpxoS68nwL1WD6u1VYbjXQeCcbS/nnzUziDNB2/H43u5
DuZ1NPgUHnjnDofmDSAQ4IPZBCr2o/9KLzqJgiO1XU6JSnipSDXbKgnCoNEwhp62
`protect END_PROTECTED
