`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jqB5z9ptO1fM0iHBbd3AXHgCLKlxKAX+eqnipsnE+26XdTgUdbsumh0GBtZuOcTd
/69GDj2Bj6Gmwo0YTomFbihP6D+F4LIy0tYalm3Bi7gfvHKx19+lwv/K3Kr/VcB3
k/YkfLfeypnb69dEHUzNY+1VoHBtE84m6DDLs5YzrW4jB5rNE7/VElJBSgNgMYUJ
eS/nU4mZpQzd7PTDMl2/TW+HG+x0ubF7MQYcqqgI9lkOYKUetR9goWP7X5ChhZtp
MLcrMZZvCZakYi5CnB6Jn8TabnQ0IOYpEY2bshFPkFK+6hd2dMqhyGSyJH1lJAjT
HlVnDLC0Rr0lk0yx+tarybMLEZMBfwAXePPDk6+NPnI8A6wBIMSoIGsfnGR1saHv
WKdeNfoYLRODASAjdg2y38jEKjpMI2wjmIfcVX9bVi0HDh7Igbl6xUwfxMJ7ce6W
9WJeilbUNd2rv5e5n36K2dRD7nwuQC3kxfaUAYm7lUZ8JOOwntwPGl0L5QFw+xV5
3ckbUac/iOwU8plX7i5MxrkDM8HmQpKjOa6oyzWvaAnFWqFWrCInoM2Yrzpqf4sg
pb8qUQL9BKRiv/2Isi7tysDhGtmYPgJub0+Dt8AV0t8KWfamz/NUjIzhUpCEY2KC
1WjIhp6whLNpkt9gxuyBzsD5fi8CImrzKRPXpNNT2EICbpiwHBO6vJEQ4FAj+LVP
Dk4SaEIxIgU9AH/KS6yctCpb2PCVCAHJMPnD3tNWrUuoekeRCg6e1pBRoZS6yv9n
a0zIYMcFQDlhakG1AerhfQ==
`protect END_PROTECTED
