`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aIyC/PClgKOS3w4nHWT1k60rdj/FYMfof7NCc49bheFSKXTK4xbjvpseE/kb8J8g
9h9OrwtoHIUzKObfzwMDSeuh6Hou5MxypoQq9oYxVoQqVWpcw6c4I5A2WQyPQO1b
FjNilUlOFxrGCVLYUohrx2Gj/CVtCZa0danJX9+Jgsp0ixE/cfWkpZ2NVpk0vhBu
EnW6csclFvnMX3XhFPGkXM1TOppcr4XP2fpA6/IQMdKRfZhxs/SG8BXs/v8hpL9+
QwRKrB+PFott0UU/tEj3AP3yafi/on3PEAy7lIbiRpekxIQ+5oqSMGrS743Bvc1w
/wfU5dMDgKooeNrhEf9pIkptkky9aT/m8P6jo14h2ja3/lZ5Q7BPu8BIWe9aKQga
hBwwcbspm43e3S0DP6p1wpQq5h/A7DHvD6PAZ50NntgncqvdB6rKMku2lLjF9LNM
yZLl5WFFbmZtossscaPfhbtoFzy+4uzSVy8Q30QWJJihjIcA0GPS3D2E+xh7CUjK
tm9omeincRdJeWt0rs4W044kZwI9QDm/qYQYw/MxSXNGKjuTU0gujLJ05VXNSjHW
a8Ckd5AkT3tXLNuoCaYyG04Q5Up8sLiwlTbPlLpUInX558MS1SF3nvNxM8vLFI+B
K2XrRJdqxatFpBCKvpxuEDtKLAoEmREed+BerEh/jiDqw9Y0jT9tT3mx1OH5rOJm
hSuMlLH4Ui+f7gMiabvLJh0mtP1wmo+vn0dbB53+FYvfmBlSLiMDRLo9WgwWPcfd
SAeE5JKE+gkoBPs2nBBG3cR0xRs0lQEhy8ZbIBZOE3Uvh9XWfd0oYp4DcQtUkjeH
VFT0obqXcERL67EDbYLCrgPkI0JvWzUtVpciLXmI22nQML44HGLqH41zI1mJkqEA
yOYfYJI+Iu3PmETAUKfsunaD9O1m04XJWU21djD3vZKK7FXiFOakVohD0/MLs7Un
lG2ZeMeeBGB7Yxx4rM85yho8wI8BC3qede3CNE6lQaEWGl6RKIHN/1YbJOg8EZsr
hR6KQQng2AJE8JvUrvDr1uzQPK2qlWul/Y6vZWk7S+I=
`protect END_PROTECTED
