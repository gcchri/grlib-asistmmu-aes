`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uui5v9OZiiqhCuhRe4y2anrMMlNfb486MECPv3Z6EsamckpoxeqKD+YW5hI0znco
5MhmZPopBqkiED4BjkrGviIuLGDi0WtOgnFhMi770ZHN2mukAzNID3XvOMdpT4iX
hkupLMjgAN0pbNVpoQMJNLDf5znodXDrnhstz5yOwEvwgqooaaFxHrxMny5NAw4V
bhJsMy8VL6s3DOxnN0RjMa2JuAvlYA9acBFM7EsJK31rpIsnm2kfnL07dGPUvBxh
3KP3QY+hlcPPRvlRAfg5HVd9abMNRbhWuIjAPwzqOM1/fbT/fyvh9yyOqZCrwH5W
54uhe4m41MI19kmFlhlAlZzw4c1dPN1W57xZv/wEF7Fl7TF86JsNGz0JEwu+WAs0
ANRB3ALoF0INlIDVcJl7J5gB6I1tfejIhvmAv9tUj6JHAUxnTgLHKyQzks6lpvHd
8yrXmCP0u2DbI4J38xe1VKkmxXyvKvNOxd8Gk46KxDG+UC6bag0D8SZRIqwHs0f5
`protect END_PROTECTED
