`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Hb1hmUVhIiwPK+Majwc75pttdZ/ddvISoQSW21mv/BskyEQ+05n0nZF4JBRf2kc
5CmF1ItkcgC/fntoDwmGjhYFZSZ0k4+5tzIhEZjWNIwqWYqKLiE2cmraiZRLeLVy
0LnmhF3UaLjDPy7tCrFrA+4Eh8EoJsYmkJ4OCA317TDnR2m0AduZLrVDFFVBmwuc
f2Y/osDZ4wsfymnXklWdubvpAu1ouZP9HCbN7qQS/Edub2sOtCh1LhvcHMBbN5NX
GIH+fFm1KQkKUYqL5tQJniICvF9MBEXMUI6FRwmzysAHimQEBdGdchrkrmMKhvSl
Y2I8xNPVLBlnYwtE3aQ7dfRXXmOWFk6PDNOW9CrSu9ftbmcf1Z7EQmEwaC7Q8RUN
RqtphzG2RTD2nxVsJOHFpWcDnz/zbu8IBuHU9dM9wH4uLI28ud9Uu6qmhbHEs6Qq
IF4HEBQH0YnF6KhVwvy+YaERgHdQQEl+NDujrx3SYby21PLrux4vBwh8Ij9zCo6U
`protect END_PROTECTED
