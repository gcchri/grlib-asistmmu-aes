`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hn/qqOSaPYWNbZnsuZUkcNvgyTGv2Lj3g0fNURWFO+ZdH2BoBQmbDOWKDYM+YSV8
1ZebWzqtKqg1crVn/Ru926qkyB3U0JBLQoEajo3VzbOGLyETb7/AwzERrzqNZhW8
U2txPXa5B3tCUlCNdTQD2f3z4CuFHgrNx57KjCKXYLqG8PPVJJFbo3TMEi1KK73T
+cTvXrJL9ev/+tDjVMtaQBNzRezt2ikq+8XiUugN8eXC063Xffjqows5yLrkgs9g
2QE/024uJxzmF1BqALb15oZC/LLiYGRgeGfNKW1D+as+ACxO8Vp7jD4kGA6JmH/S
XuLCnSfY2TiNTshYMI87yEXZbBcsgwwhGo3Kk11v80+77HgVNLo/O6RVjzIZVTtp
KyVnEZJRSAOwhDeTVuRGPVXIRrl8dBiHC7lzrI0iKETdpzFB4hjKIs9GEGNOItzI
cRMs3n64Gm/imX+jswKcNOa0jWO/+Qn0ZC4MVjYCBS4WVTgp7GUCeZ7S4YvfiV88
dyEFCIdE/QHh4eVxYFElaU5vzGc48bkYFkgzAVPDYtH42AXqTDwx4pyHu8YH1s2H
zWYQmJof0DEX3cPF9JpdBCHPzbnpBrevQhLfcicpL+n5S6KU7eq3eHJ0j9jYt0nG
RZKiQIjyeXSOcppQw35LTA==
`protect END_PROTECTED
