`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DQV6wJ83t3Tl/pv70Mbg8aw4RCzPxl2upUoOFnLCaOxwfeSm7rCF/LaRac031wm4
8jTuumvk8ubAs3jWuvcBmxcIb572tVWqKQGnFw+jI4EuAH76CLWpRf0CSbc8vnrf
3sipb+Mc3aeaDXlpG3OviAmwcwoi2IFE6IpI2FpfWR01i8fsVhpOL97EiAvjxg/g
XuU6mzy5oL8nfMB/gWR5/XYkgvhl3XHA3r2Z/0jxlAUuZlfKgGETpqmHVNpX3bxx
hM4Hn1d4By8uTJLtkR8JZqIWjsrqipVn3PRU79I0CR0tK9s1syHgRqELGEmIXXl8
svT+xV2OtMslFJnAPHziZWCEQJZPZG5+8ZJmo/2byDfBT3/OKs/FTpwuLQ297OTO
Sjf5SexwZHZDHGRO7d4xFg==
`protect END_PROTECTED
