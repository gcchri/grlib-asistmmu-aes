`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wvokggDCuf7p4A9d7+U7s5bZcZqzVQY4S6FPSOGHdJsIancQKCLTFixDzm3N4563
p4DJyrN98p+MVqL8rL5L9revTseHI69qtC5UFSh8EZ6caLj76WlQzujETFCr4SKp
LpI76cDPFG0YZT0BarMTxFN17/S6JY2WeWzeftB/CWvIIsRY6hRji+PLDML0Xlle
8SdtI6UE1H8cx5ed4bPZtJHLeJJaH+3hEwtYwLBiXjvYKEfTNwXdSA1JduTsabwn
eXEaIOufVNkH369tCxXFrs6FnmFEwBAC0r1ehkO25whUUS8hnu6gUqa4pfoHEEVc
Tum5vUON8catB9Sggpy6yQKR83MB5JKgaM4XgsWVpWLzN94lhoOEQEjWA+MzjkSX
fDKj9NjV2cMz6dbNqytaCa1XYgI/RH5LQwnZLDHclD0=
`protect END_PROTECTED
