`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SLjKrr88Gx9LKIZCQMyqpYfcQ2Qs+b7JpU9T4IIptIQhwnZiPtq/LKnAQan/s3Ah
EqWCxiJBYqJOMND44XJmQ1B8gCboQMk4wuc8fIe/3+G3JzgP8zd95R16s5VcQ9+R
LrCSLqun50K6ywVg4qNsJIQKijz0uWD6vldXRII9qWHcTXp54yKjzy282WMwvTof
uvXX3KR3Mh1M0jNOO6eQmfBHZv5INuF1sM6SizuC6xph6+YqMQX1oUf5TyOGL4cM
etGjnmGaM0790I4PEAi60hMs4VUGb/othZ82E6DTH3LdrV9dqIbi1ycT0rDau63G
1EgXDMOMNvIBAQAx4fQR1R38Y0Mb4qArLCkwMlObKjzZQUXkqn4XuMAavz0Y2q6J
TaCeCZCl/ShiDS4gj3s5xgcrLiLzdISaEZj7XYb+qWvg9QVrINgTM0Fxiiagoz6H
zWjqYqTf/XaI87JGwU2ZUkvUMXMzzvvyPqE6XaZVHbjn55c5UcOkv8d04dtOLv73
`protect END_PROTECTED
