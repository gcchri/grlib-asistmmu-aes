`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L3mVhTZTbf//TnuwckxkDgJwomYTCW8k5RHaWzge88haAgP6cQgPfWQAnVs3yh9s
BqQunLNoE/CYcB/Xnc+Nlsyl2lBcFUWkEeKQcbt7JUYuTnXgvEmLWPx0EKwJrag1
3Vn8bL7HbkwQOoVE+mKjyL2uCHv4RrIVVmQ5322TTLstpLnJhHirG5vrDk+samuv
2N0iBkI4ufJ/F+PJIqThIR0Vb5elkUfkK8mwMw+o7AkeUEcg5dr4ZAXZZ0vNF/hf
/xcFMa+npoVARpiwqHKcOJG8C67Z6cEXh1AnHg0ahpAGt0iDYpRZy4AS1wgfSef9
oN8OSS/gjhdhDeW1uFcrHSx55NoaYEjzlPu8SQp5Kwgc+ttLwCPpNrHzhCdL0caS
mRU0cvRKeUEPxr9CWTMVSNsOZMcQwnIIUUobDHaYyCEpk8x4J35fxbnMuKQfc2U6
4IKPJLYKfPF99HdgMtz6R+VyzrukuonH2huniOPouSfeng+2EXR1ltUzbpTcbhB7
D0sueDTvE5QLkfUE9ik+evOROtNxR16sA9ryNgrBb6nFrJuYJlvqnd2Atr8bCcxD
O8ZA/TdeJDBhRm6t8Zkuz30Y0geGtBmfFqDybQNPf3Yau6YYpVb1BDBSjNdcidgw
Trhh2VTTnlVqI6ZD1q/MROBNT8AGp6QiJbvxH1NYqfdAEX5AbhvLni6v7TD5H6PU
n2+H6ERMb8I7XhbBeo0TCd77FDMAKJBwEj7PMNNhyCi9kpNulajAefoIElIIIGyR
xhp9AxDUiLN9Kzk4SlIHcbIql5CjQNnohCjbxH3qfExva2kxrgE9P2FYJC8TgQEs
erB2+zWxIql6D5O4KSfrScew/ta5jaa6LtHbvoFLrYmcukKOFkoLqayJ5wpNLxn9
Tv1Er6qQTtlZ4zU+Zqq4aE5Cm5tCrtbrtga6WoSobrC7wJzDKSCZO90R4OKRctuZ
g+Z95or5DcvSNaJfvfV6mEb8/sz67N75PFiHRQe8YuoujR8XgLAKUNusIsIHirrW
1shwzLjS+zds4pmdIAq32LLoIMm5lxId0YnNS4nS9Pcr5s5TyaeETT1ucLdn96/4
XR0N2eNXcgwBEOCNvyEl+/eqPz2hO2BGoRInQFsuPSZ8lmz+WYTlqznY2BwnkyvL
32GDGMbBiHjCz4Hr9HaYZfI0aTwCZIiQ+Vg0+nsEHCTEI0oPgACfGeq7zDPjItHs
2ZeaRx1ffrjkGkAVWB1HxmlCw8/+KV4WQJHiYw8yM+fi+DJ9XHesqrg+YnHKka6v
Qeyb9VTVwp6lmsMjzbpCHObvF0CkAVK7DKjDubbtPPKdSuye/LEz2r7K36KbX6Cm
ngHtBmPAc1PFTrkXOt6gsACrzzkV2MzxlHJRtAJ3/MKm/B+xRruVfx14SZQMO67Z
cPHlXdJPIYTFzGXPHu6sPPwlM9u1aqWQkm18sjAO6hROWTA1lKK/Eizfn3ahLQUN
+4CQyPzCIkzFRiZZqkkEKn9y4NiOkejTMF22PERHeLjchRa6QrTyMIxsXHrQG1ou
Cu0OhVvnXJ9N8keRiMiC7gmVK6QgnFJtGkypgnoIN/Fc09QMs5ltnqvGFLQhhhLB
LpZq/q7j7RIHHUdI0P11EPEQu2G5J5oJFo9G+LzwxWzWlNOJoZK+HKEcdpgFXcbv
N1FJ8Y1KBBEQme2LuoC8JJ/0QW4rpAn8si0C+ApgzhnJhPcVMhPo92yRUo2R06H6
dSA3H+oz0AhbO8uQUyUzJHViZIdpVoqvnwN2+YYAEjksS9qzEhZBuf2ak0lDcMGj
3W27QTywX7D9ZAobOxrmTG3dCujtulrGj/7Y0YywewRbcgBrwyHXbFdlBDH7yzxL
Fl0A0tk8SG22uTVHyZtP0xq9zHUhZ6NC2u7lZ9r/L8zMsO7/b+UPOZ297YNPiIUo
7TEa1L37x8xBu/QDgFewcorSOBMMXT4i+ta6VT7zdGT4FjkpJK9Mw36Tszm92Cav
6TLp44q4T1DUet6vsfUf/06kD0N6sByHIoCaOkT5NuWMYZ3sp6aaGAUc3xUxd+Yw
GZzwOGAN16qnWecDyJ5nlKVh29DhyQ7ns+sBnRIFQ/9L5/fBXaHgL0zqOnRnjFNJ
VXoXRpKXTFafzD1foGjF6lskSySEgrqZk/OfDaXTDS0JLaCI/Cs3zgDIr78CJWwu
IULiMBL+6qoWoNYgYOOG9ohvH88Z9jlE/ebv3/DvaaBfu4inT06OnX7rWN4K1Wd6
pfE1wVSkGS8Ombyewkc52p//hQNtJyd70WrdBp/YFQ5lnVfbGGUXafOxZ2NxksuY
v7aaz6++FFA+jAvj5PCimrOJTvhdQZOWWIJ8tt5pBi4ozRLLhU9XkG2hYUnI8F8V
Hqo5co41HN/CE/y03VZU+DMAiP28a6RnIMo9d0YOslxej0QqDuJzrqF7ai6m1YxM
c1a9Sz7k2Zc/DmW8t24v61U3rCkVVzw3u0arl2scnTnhYQ3/hKr1L+yFfgsRXKa+
ztvsGj0QOW1LOl1hO+ZNwsOVe1bbs8hNWtRaH4MM7beujz7GOvKiyKXUeDk1BWN3
CbUMmdDFtPtI5D9d5nID1Qbe/V4uWtgQrp3epydY/OShjJDNTcDl9j0Xnvaq26Bs
BeZ1z5oa/oGttrVLtarkxcNpyZZBhgyvSdOe9ctwzSYutbPoa4pAXMfMRFoibXjS
txbZdXDcevKJH1oz2Wi1yhRGLAq5JgTj/sH8A8sRP+8DiqxehaHv9rB2gbhDpVVp
70xM82u4/CrmLeZLpXDMd9V9lFXA1OaSABBy6VFcVV1xBzB7xt12AAiLMzp/LAtm
KbQpGbYJ/J0J9q3T1b9DbeL5enEjsiYDNpjtOqdWQAevuWDIw+nQl3997S/fcvPn
T5eJhqa51yJ1EUOAG2nhP/EKSqnwb9eHnbv7IRCQn07q5Fbt6CMGbLT6qYzSi1lL
`protect END_PROTECTED
