`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V7K6bQ8k8g593/FeKJhsscYBfVsNeYQbxPlqH6C0Wa8BqVr/Oky/DW8x2cfoHfn4
g0kI1+L97DT43NqqURDh1RfND6Y41uZamg9jXndOZTsrYBq6fKuETnchiGEUmLS2
cCLeSzOzvCAcQOwBBvt7oSe8X1QQjLj7RPz+HSVbF+oEa+6NVOY7E6gYHJQ1qSK3
ZknSZoBdO3eb8wyolbB7u0zidCnubTB/sCsFER9WrnnZA11WwaJVM87yNdNiqwlG
6XvzkvijZHB1cVNkVAx/YHgjubz6ceI9XZdZ2SEvYris4Ekx7NCAtXJfAqZjlX8K
nWzAtZdYJ+GzOrQVLeMY3OG5nfAqIEgS4c3HVwODj9I=
`protect END_PROTECTED
