`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HdblRWFeI4W9yAhmM+USDLbxnikD6vdmF+OgEvXRaQFQ9L+A9ygNy+Uv9X8y1pE+
4c1v/hM3ePHXax2trAWJBH4slk/0TOwMcHZa+iXFIUhSMfrvQMKb0ga6EXWSNokJ
uP4NKwDzn7ei4lgu9+a9kNtm+dze7qnHSqdVVLuyuUrgc/dHJV00DjfziIS7/6HT
bX33Ji6EPcI16a3JkAy/RXJfIAyppCfWfGsDfu/EZv6HBawiywhHnBFqHUOEwScy
8ryn4ENyxWxG4UHKNUKNU2UcRBP65HbyVMTZj56HMEaFptm/9lAhXxneA0x9JWFc
MC7XtCc5tkeEZ+JqqQTT1Nw/f3gKGF/n72MpiXGRMC/Nysf7bMWY65yVxKHUkKOU
WRVJhHWSmpRLrs6ce9XQZQO7voPN+qpxu5EZkBAAXdlJXSH1bd5rFfjbpXxcZ1wJ
gebFLdMl22pTnbn4XHckdA==
`protect END_PROTECTED
