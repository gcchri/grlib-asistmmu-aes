`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hJPBsR0D328qvFjhjrgXXnVKBsH/hHqU82MBbFQ7AbR+6I7YROIwrepZjNKOAquC
2rWyhKt4tgrn7bW8APwgmDIdlaw08d6VGLk6FCKdNzK9ZYXd/ZN4oI4LXZLFyOFc
DWO6FQ9UgUkjvtku6sVDIMJ7MloOITntsUPRoT2r93/OHjcgoS9JNk+GewjK8RTK
TPCKU4weMPUv5lh+Ccv0kQfhWoT/KK3FIDbILBOtZfR2EMZMt/2/91k5oD/0k7OX
0R5Cu2EwHRM7tf4X+uMNlG1+9QcbYnWGKYuzEmyEZxiwxxyEXDpNJMm82xNdq3W4
GVmuRdmre5scvoId3MNGRBFYImlm4/tUZLvGN0NsH91vb7RI7bJ2V497lXs/qLKj
WN6DGXBZy+A9bV8MiwWOzVvxrPCA+idPRzUbWtOVhXCp2I4rL5WvcxOXd/muXuAN
`protect END_PROTECTED
