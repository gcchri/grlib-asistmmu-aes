`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hrnXm00WMTJVriHpDjlVeYnoU/crLcWfx1FMS/qKFnVXDR/jACMyroRt+1Ya0Gtg
lNtkYfRxwfcAYooTCoOH3jaRYmi1hoSbR1pdd9oHJqMDp7ChHuvdxzQNbUiMx6Dm
6XyCXKGQaKh75n66jVrV4NPm1RMQmW08t7BD0PhNZb1+j0n2Osh3sGwjtgyjgpiL
zTRt3Uj/vhvn0rr7MoX5u7ok7y6775844QywNQhgmpegZFZnH4gaKvN38B5h6DCr
mYmwAqNF3yJ1423gqawG/56Wb5+cDNmauSrlrwXy+2/vmZLDBlIXqHOLhL7A6dDz
17fuok75SjI3H2cFZ+fiyjiS4W86gsKlpSpXj21Ep1t8Pa+jzGHIfZyMElkSIr+m
5lczFNgsmMlyDtojA19ruMZbgJMBqfdUuSqlRzCXyi/ElScR//m7LhF3kkbkzRLN
HLEH2RSNM4GqlVxQCwWyHZz0e0i79OU8fj7kLYdxB4xjaD+Gp5iPb4hTCxAvoX8k
ZrjCEndQSdn0K+rIuP33rHkHucWhBhMKd+V1yKrfcPwtjpUOYC982yUERgmmjUnL
X4Y6yKdM0EOPTCScBnmlIwwDNhxQ1ebpLph5FsFP4MGV+p6peb21owh0CMpep7eL
YKgeRd+pClYc1dJ4JpKfs3f3T80QKD11y2fgASOjtqrW2sBQ/K++gSjLOB2drsXn
aEYDhzjkVtzUvUS2akKBvgY4x6lR47+l8gCIZr6fkllkhH5VHTmBndSNZ/fz1spt
U+Ycd8FK67AAhbe1++w/NPGWVFXsYrokLUwa00oeIMlOq2sJhAhglFCkJgvodXs1
zGjaD3RhdFPB7RSX3ok95P1AYTpmEHjbOQOzvn9kVJoQmvlLuH3l9Tg7GlxJIvB7
xt6xnwW4UOEAG4lAC82vCddnMko+ZlzTGY9DVs2TPFZWDg72IbCOeVJ2DrBpPYa4
hKxv2d5fi3FBBQ7Hx/wgu70thHgNxRvJR96Yz4Bj2irOX5qQSQIzoNqrF75rHAUO
z7y6Y9q3M1QOJ6fVzyvs/36IysqyxEqfY7gj2QzxnpwVPPzswaKIpRILhqpGSXpM
s+Dkf/vLYIB6YmVimu4EurQ6F2SjRykitkZs0Irr174Xr7dqo3RNA8gLxvao5NSY
RI4z7ct6NpVGC9JSSszzawGqEZwZWev8yDexdgLEhNjmDQvrwLCq6/HVE//fsKhd
7VtRUaSswH9rj/ytEcgHrTvASAw5jePLMcu+O1U4ucuiqUY/4T84lLfcr6E0JuMf
OUg0U5H3SmUpu3FS+2Cr1WTnZ1L8zuVZEzvelOMSI0Sjo7xH1n5ELIsNcZuTdI7Q
4jcZGEw3FsAM17ASM2JcurgVSvT75G9N37xLdIuiEDto0ZLC5F4ZXcQOu75gjltW
8rOF1PN9I3T1UlogzSing2Xi6mtcAEr/+zOZmXCVKeboYIekSy3Gn/kobHvNtlj5
YkN27L9xsbzzvxYt0VnpGWcNadBaCnWhS1dgrDMcQIWFwKLhQB6z6+TDWaITn6e+
qjWZwk2hOT7VQLvHeqHIeGPtO+vFzi0AhGkjDml+oF6tm7q5Q4E+kFqfeIXeY5lQ
89InHe+/mGxw+J3uT0QMoN09j8czrDw7PLtGhOdavyP3Utc7LHtE2cgqbZt4Qqj5
WQLz22JH4vRrumkUfE8qsujVlwjfvQgzXW5ZIO0/WQq2fyoc7iERS6u82Y6iD7Ld
/nGICBWSXh4RITzuIiNmiUhEXrbZUd1DgtaAaoAXo5qaZ2ouI5QqTksrkOMGEorN
/5a5z9WVWy578U9q/mv3ZkoNzJ64CS3oTi6dS5eIg+ewegLv7Sn6iIumDZ6QmntK
PWEPgznOXNpF8FkPBxJzDoNzCU11HhtqN4o8lxrpW47oSL8saSn+HnRWu31VOhAG
lseZwsq8EgGvhVWOI/zW0QJ9WpJal+3NipR9P7nHXrpZ2XuGJF+hpwnTTuIEJF93
oCoJxCDEGqZhBVPUA/S/9MZ+0RsAE73+3C6C6pnEF8o+oTN0gllURFzTMo706jfD
4luP5udAR5htrZH9uNKqgXtwKBLvi8Z/MFQTaxcwpUV3SeFz5jkQtTrmx9mww3Mr
+MAcIUsHsyiiGHEbP50eoOHsJ/VJiSQNnqZ2TF7sLcOGQE2ANY77rRg3782LUnV8
iWWL6eFHF/BWzia9+RIBVRo8UwHzZQa2XAc13qdnRDsT3YuP+TaVKHZLjhyAdQ9i
yAaQEKXq2hSvDfrfZ2pUHhS5SdnxDut43woGGbOoLy1S4y3dGbN0sTfDSTQs1fQK
QgmeKpSLvCwJ6SJleE9Db/Vgvpg0kL6srst0aeyjULbMyooyf+XYURfjdku+f+oY
MgtJDJ1+d0UAAtS+euyWwNeqNMeyU2B52U1u+NUYldvmrLGY8KuGL1HEp3Y2Lo3Z
DxUR7JIFHrsaKK/1s3xSjfCAF4QS5fm8XtOgXSoMjlbRyy5nrUj0vlcrg393TCQi
VrTZok7O5syTvCj2Bj7EyJ1SQf+uSAczuvUjXERB8zdKS5w6OUAumkJKqduRVjOT
JfgcHb4LIToHFBhAcRsvbxWOcPepstB8oADfjWcMfUBuEKAlfrqtC7DaxdFg6cGZ
hvUXPnjsiHmjbZguXAinE1sXeDEsl9PXQwWhUnmbbZ3F6LRtE4GTakvI3c19rQfd
5tFhU+W01JRmOSxeTzLPTP32yk/7CjBUFVlTFTkuAA7ytRLbvbRQqxVQbbB+5Tlb
i3OfLrzMYL7MZOHa458gfnikLKPH5X/SssRdf+KTgzy9cIhjV4oJ9CX/OIckT91t
Z0SswEDdbH14kr5QE/u0mXzTThatC7HgZOdXRDxz36NYARdoSiYxwDpvIvBkitTF
S6r8yi1PMHI+UHmm9VKeyw/V5MD+rgKCl1Ki04G/BtyPvE7DlIoOlV+9TzEc7SAK
ego9ngjTXpLRPTbjMmx7eSDjjD8VHfhmTlHqDx6/2Ub2BAzQLGLmhuFpuBNNcC58
P10gYkrOMwuyKwlLC6ls3pazqtA/EQLQk55zURRN/8lHbI3QhJOAaanSADlK+dd2
vlopODlMf3ZhKRgKlDWN/7EDg0tS32+vuC9JR0yEnGXKzek838h/m8KzUjtwwlfu
nMp26jMFVZlhF9CN0SaZE9DT7+MoGPxjTk8Gy0mje1HnkPomqHLtHIrIEKb1ixOj
B4z1YnfJw7KJPRO7//YSOLVuFu89RmVmV9NBw/MgRWjYYHHbOzggc0FVgpJH5eJe
24CzZXlfbkzWDMSS0vS1QbP9g8neiriz/y1ww7M9/fHjLmwqRj6HCcfXQ3oz6GOA
LaYXOK7V82uT84VVWd0sodRfBAtpb/CO9DDZGU4lSuW5vhcC5TQl+MCQIHOZtsV6
0t2KOoNtY6A+jqTPFf6hC4MlSVxOZ0otoWXSmossXyz4JiwtZKt3Ft4ej+Zm5otf
SKG/yhbaWy1jBDwGnLVQAvGlH/Sl8XaYTioQWqK6tXY8HC8RP8tEa6h7VmbK7fqt
6RCLQ+MlG5rjT/ozdB77FPN71Rm+dswEKzzqVwwMYWkFOp7ThZ+hGhYKiODeNKfb
CyAgpDVgkiqawaiHmnsMPMsFHmJUHOJJjHO5MvcNk0BI94t7BfCAq7/AdLGGasML
67p/zrC2a53mywOJ+VEmQcssUYAyQDJX4sl8bWjaEZNUOoDMnVvagcEnJLhs+ax5
lxKYGoH1O6dwqNCCl1tkzZ+LYCnW17eu59AjH6+HMYF27B/+c3wUKK81otHKiFpj
CekudcbohNIoI66xtpMoj6DQtTJjHc1o99V9sOesNvj3aUk5pDKkqLnHyvpI6T0o
uwW7VeH/sXizl2COc+zEmbXNyrrdnpiSL31+9LKPgqGm2CHxirASFMzYio/ylmLK
dWGT7Bt0+rTU9psixRU/ZLDzryTAarhlNF3FeYsYb8k7DjdPL0nS21Qiq7taNv38
IqDhkpRv/2LMGtKtwHQok/kJY0HzqPA1GHFG3cK1gXuFYFlUDR/9s9l29OjZ17/R
kADx8BjWPvaWRGEq6NEP3BuVftOWjnk87LaIf0+AGqTS1Tr2bC5wO2i9+p7f+Nwq
nARFKC7BixuSWsWtk25DMzlirLQN26rn/plRUugyTDU1TZYPyYKJNeJyd1xEy0kw
/j7/TeDIaQDMOS3xslWbdDF66ysY+06RCt0dXu9pyw4KA6ORc+pWwbzrGIuqAiSi
MEp994G3UYlwAzFyCBoLRpkVoYXLWZNa2/KoU7sNkgFCXsd8Vs8fdZbSq6+kP31s
JYKO3lJiNxDpWLzxnpcGe/c5l3ZIjfxwTl+rcxGceOwDj+iDm9qhRTldCe942GzR
2fuyAh5V8QIGwZ4MRnSR9MpuntvGWjPzlPFs1A9G8IJ2Z/KWhkl+z/3vsKa42jyE
sI5By5v9W645+kQeXKOkOkCyS47m0r1mRHgz6HkpzboU4PeRU4DqiI0CYu+1HaYM
K+zMOuzNvN+2PGYu2tGyHi2VZYOhbRX5hjGlew5W7Ah7Td0mui970oJ3l65Xk/wU
br5MLCn50I48IIEwXdEWCIMPh5iw2KqaOTK8pzPCJnFlxXmmU4c81IDnrnPOSGvr
6bUauGlpqlea04VUuvTO0cSXBPOLgpZbR2ifoSuZPyuOdSI03hvwK4Q0/oEL6P46
7uNbMXeNw44fiCoLegqUuLznxcvwFE5568gBn94eLwStnN4wYNzZY5TYmT/1X0IO
4DF6frdsgRXKXz9fwRKESpXgbL2whcpEOGrIB6Q2iCgl1Uu6cH4/fFcIFs0Z9mz5
olnIEHHEzaEkCj1qWqCxOd5pShPYf4203Rf0hFc6E2oJWHZ4EfyNRvZsC0ul8Jul
pVicJHMyXlDvxMV/+A/EjRYLrS3TUYyRmWsbZOA0lgokpV6oC0CcUJSnoWhOHNiB
fAla0fjMI3WQHwCroYibndZTMukUASpOJBL4NJoIh6a2kcRon9MHvYJ8A17dG8vO
h1AeLzCIzz4LT/dw16W7AFA3WaBIO8aFmiBgWM1pVbYPoVQ9Lw/mIEvN/ay56RkA
0DUPRrSS7OoIHF+iopmOf8fPqNwznIjpEQyZ46gfSj2DDBOSO6fwNR408NWodhRW
KX2DpPKu6Zr02yweaa7EG/oSJQMrH3jk/kGm9VOQFfCJPuVngzFh5OhxI1HLJ9mi
QPQyFAlqzfy1wiWsSe0oXncaQr8M3bSzGFpA4eV4PFPUOSNP2L9yRwRIAED6ak/Y
siKAWmPgh4EiiuAU1q+9w/UYlAFIBT/M2g0Fksq+WDNK0kzNmnc/sKnaRasgBFaJ
5li391H6PtyhfVhZM16dvqIw7zf6S/Qp3Mv6Rq+JIO0=
`protect END_PROTECTED
