`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i13WTOvO5wiXEJrqlUQ2B0hrgEumRoGnm/3F/LbKknzgkzGP27YCKC20MhosEU9K
u/FuiaiTJPp7MKsXYakZe2OZ8sWCi+/iBq7BBnyw82edr8s+Pv6URfAZrBy4hCRc
vvgPqu1rp8XuUR8OK+obWXRjHI+aKL+CFUwDvRRu+tVpF6puPBZfHJb8gXob8f1Q
quwy2ZrOfAsH6/pkoQNh4cyadpkIHyEMFndwZVMjR1cnp9rxdCwcrTh0QSm8+6pB
BcpIx+4h4+ZaX3B5KYNq5HvYdB826g0G8fz8FaIRf+CLsWmKgTdkAsNXkCTO1WY8
Zb17TTzz1crhjr1peqqVMOFyEWhk9zI19nIYtF0F/TbigS9sMh4Hxl2dY8MoJlVu
5S7sW0CJmGf0D8H3Nwdks6zxj75Wu5ir1qfjnd2AmFay0yUd0T0hl1dD1MfQJu6P
wsKI/UErWaXe5sQ7rq5Xe/0KkaefR6UaJKkn52abaGeL1GmHgEN3Pn59TWuwAQZ/
ABDPgmBB4FC+ikHmDRSWuffTppo0wo2HtwrFYk0N7fuB+R/2WHX9//U4aIoEwJOc
+XjO0hwayNHQEvqrFawu15ppQs9AqZePIYq7hqewXdof5G0EPnT3ckuGhsZn3xEz
`protect END_PROTECTED
