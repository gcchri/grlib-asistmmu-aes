`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3lTHqSbjFDHJfZXyh3U02tK0f8lKeqt/PWomhDWbBcy5v4su/ppaCVGv1nd8FRDm
VtiPV0XdYu+gMSC5jLekYwWDzNhKV4tYtW9vH/lATHIhLlVp3FkarDogFzrPRU6s
BBcnz4tEw4uQt4XyWBPSF3+mSESV2Cbd5qdAmduqa8CQRismw3uxs63cgR74z2Lh
PUxRkzF7R0pptlApJ4cAWCg/OQeyxQXiE11axU32h1sCE0XMp8llW9M8Rr201C/g
6wbZSwNy3tmEpdDxVZxJJu4Cz/nTbH77wQvDO7a5bVyWNLoTr6qi4V/J1SQzvJ0y
hRfd6ksuOx9QMEWjbnWyrpnhC3s1QHlf4g5dCQ9jTbA4wpIF+AG+JQnzcmyOHVMu
Mno/BgyzbfUI5v6EfBpQcGzTuWb4txaFgf9ApQwVweHfSPStsl1PPJolIcFb/ezE
S4Zdi+VnaBACwEnpuOsPclrUewGSklDEqFm9STHQR6sPHIJqiFqW9piMVsC/LHzW
`protect END_PROTECTED
