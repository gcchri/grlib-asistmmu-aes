`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aooCs+78VFGCT6xFniH0acpooWL0oadJ7dsCVPPmM/kQrB8Yqz5rUBNqIahOssqm
tSFibeIGliMSoRUYf1dzO00u3zz24FjVU8D0OBH1yy5crq2iWS6dsAOGdKYSD9Xg
RlfsigCvvRs15iXCzRHPmkDvBXzSBrUqK58rdPJ/oi14xcNah1bEy+WtdVALIcd5
qihoB+TG0BdO1aJ0u4SusDzmgMO7HFLIDk7Cafoep2GIMJySgpO+qWMtBnXM0qOS
E6MgmZjdJixIqY2HIV3rcw0vd890QnxjRzrSERs411HOEFqHgZ62B2TPHqBDYk+6
ceGd97JyZysDw8wXRKe1CjE+PZHNSjGZ4leyVWlWPVip7TUZv4ksAMS8ZmN4ZWl8
eH6F7eGoO5jPuePpYzF695VyH3G/xPXfIyueXVug2wBkjlzPzaU+RxnrZpvHCZKj
fAZPHLKQx5HzfKzbjduarPDOIQugbBIZmn/tmAf8XMyrKiJCRObxMR5tUx3gQDhp
+Z3OLcD6s0SwRR2cyGDUo2wiQ5mK3yYPWb5RvrWKyqA=
`protect END_PROTECTED
