`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gpdv8zOrWu7lcqRjliVG6eLi3nvcNCp2dtLu3bjXa/sIwWzewfUHYdvRU5iTxakp
IwKdJ8Kh3fOYriQnWnY/Y6CeLglI8nQIDpS4Kg6ug+Ni6eOH8lWoGMFAgo4PXyk2
Ma0WZsuXLOeyRRenjB1fp65sJYYMPwjQyw0xjMYGUnnwmZsdwvD50vOC+sX19zF0
/vKp9lPfpZG2j7Pd+79zPLl7tm7wv0U/oU/zg/KoKBYbdmhuc8QqUH2yUN8jLWRL
s7ysSk6k8ObQgNSUqzYY/L4UF/e43+di4q/aGSzZWoL09YovVXjIN0fK7n/SyPTF
AJ4b52m2d1Xl/vzNsxkBldc92ffj4ft8esxV5FfAcPgBpQWjDQl8BzkjgJQRGwyc
kfnQIDdhwKrsOL5HUh2QpNwX2wtb93rQAeTr0hv0/ggKviQupwgtz25VILWF58Wt
jYDQ+qeQ9+pMOXhXJ7YdhcgYHN5iqbBPvjH4vZq4vAzl6bMKHCWF+UYIzZ6Q/G0B
cQU7AeBW/fh7steRRL7sFgJwrkJJVAj0GQx2WRhF4p1iaZkVUwfm0a0siIGbNMgU
j/+uLUjqgez3ulX4II/puweZnF6+ThPb/WsmssxGmf3qF5r8pnk+YCZr9KqiT9R4
R6aMj+1/1nLcI+ZGPfeXJ4c2DIUW5MdgaqsR9jP7bI2zIb5Lp7hLvszJ8GlhQX42
uE3RYBBcI1ky4xN+G0FKDASLHzMsGvWyFxuccPRGpbKYaZ1dxpeHLN1nzF1Mq2sQ
qfbV5hhnFjC3UBpJTmw/p/4Q8pTzwVGZ/2Ht1wEBgenm6bnEszoeTT27yd/plpHS
MBbfSptSVrRRqP6So3MqviAx31MS9Tm1cwXmwEdVDUMabxosaYj1l6urPdjsVyNq
rnvO/SGvVlBzLe3MUqrCu1D0KirgdQHGeMunBi9QX1Bv58KQt24MeeE48xZcCWiS
UpJiOcHuk8asRIXFV0BHicUXWPi4GCL4gdCkxxdmgg99+Ls9DWyHtO8cuX4BSjGs
SbJuHOf3rLuDmG+YBL2oV4s35kklqty4PkpOX3aqrw23UCZd3WT8XHprDkYgv50D
RE55lryq2RpsXuMrglAuOxVcDQFyv4CJf7PIdIsNaViwYRozeFbi7i0AAy7dKc4d
ukv7qPWbZwMjkZzA20hTgnK0p1N15Sx+mA6mpHBnMlPErrvrX2Gx/hBlwQpZA8mf
HQrPANwJBZmWqRKlh4fDk9jzm1j+6Dq54gErH0rpmKuRI1CSaJjA10MUYYi7xryk
Wb0PEllSkTZffZxoTa2m6F4A1KYTw50boJlpzen2XCQgYLWjX1+x3QwR2W8CTwI4
SknsiOmwOPYMvcNNP78HVfHhN0Ixb2bCCkxiRXteKlWnSbO7mNIS4x7K3WZXP6Xd
AzkRcVuldFsQScjWiBtdjZlGNoY9k67bBhn3KRxXjVLTSc8SNiHfq4mkk+k2Wl7i
WynR2xYpqjpEE4+97OSJUpB/nnq+F/QwATxO43Oupc50nL6UVip8CxaZxRFm5c8K
P3LWQoS6P9dBwpLxIqvQDAdYj6xSSAXLGAci+Ch0uTYPk5BTiFvcUca2ZlMihNFp
SdrzwYhShMOJJyw8yDKFDOgGECdSKYntpgEKp8GT7TTYnw4erIxzeH8HlgZLJ84v
BIvibGoONsQs1StiBRItupLBmUHcPPwd2BpVaI91AL8F4NvlkYQHAUmp2ZtgAZgQ
2aSyVLJvG4kreYC7hfZnNXlBxAwRjrcP73UBwOiY9RApo9lqcO5qTkayA4vq6KLW
fv+QYOND3zNMxjPhgcwSWtPhZ+HXTem4h4XBmRWQh7rWaXsU/rS+oVmetP3+G88g
V0sdI6RhrZLL7UnG9mnC+vEs3tVplm5m+1agiU4Vf5SR13pTn83KLDNa43G2mdWp
Gj+jyMql4nRxn+VxWx+5dXZJFpi8i5Iol9fLMBI0rpsSV9i/pfx4t56VhJBuqDNO
CShbcs1hiUjLwQaTgPh/I+7JSvw9YHKkhjPwzKK7HHZUYmJpx99Qnfuba3UySIru
w376U3N66ovACBNDKIok5p2XkvijTQ5kSgOEOB8+LhT11XIyVyDiqsTFbmwoi5dD
ex1LW8Brp8pM1SBDIfNmNqbxCD5yM4NRHpYofnc7JYhAxVSx7D1hUpxL4EuwLmFJ
Sg28j9rbPpxws91Vpe3cqdfTmvz2/+BMwsJM06ZlrZYbUfCcXDGiyqa+5pYVM4nb
x/jPf4KgM9bpvNVseZ1SRCG0lp8qdzNydql1Sfl7Dh+kupacmzsGuJWJaKyta5vn
riEVRQ2juT+aRtSMEoYEYcmXsjo4oAGdNEQlvubbl7uqbIIqgbrNF/az1Fwqb91X
f0JGiWAVcKHI/2c1iu++dK+MukogjvhIjnt0wmZbo1Ivf1cEWjOIpkAZtxoukXb5
z1iB0h2FjRcmLkeW5l80ZVZKh29A7jJMtjB7NRtW5SV4blHnRxWLiNOp2ECULSkz
f8mfJ6gDKrLi2E8rTVymvcRpXKcCXfYFEr6TWcXxdnxBKbgNc/SoBuPhGn63Q6ZC
a6Vl4eaG/upnXCKWTZT6clk5kTswzMBWM4ruJjTFpYxUkDHZZVQ0Pf7rsFjLRYZQ
`protect END_PROTECTED
