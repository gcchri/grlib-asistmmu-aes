`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ecjNnahVTftpwXPPw5U75MLQE3mIpn/XhTOtH9glqMmpRWAGqLgPeheFKi0CsvTY
Mk85lFKp/nwle5Ryg1eQfiQe04qsMerkc8y6TKsob8YAAvbl0zZW1st2KdUrNfrF
RnX8xuodUmbWB/1g0e0J6YmpwKEpCUkg5gI0VlugRS0ZkP+10WB3TXkghO41Ivqt
Q3qLBIS5SiNWlrG4nmyGVRYngYBWibxNWTZ8Oso+0BDoHRUTi/cvsFc3l7IrGFto
qSdMo88SKLHM332j9cU7RvmuzpqldYgtI3LA7x87K51x7xyhiJjQtncVKnYO7McM
ZDKr/Gx1YcD+6NHVjgCktc0WUoNksjGwJXBHL7DsBOoSOr9M67E+BBDJW/akLGWB
bke27hFBfxiO8qbNO+hHVkwI3Ml5+wVOVA03WIruNnJRv1SaOZrvExaaArNsex9y
lnoRmjStZ0zZC7pjQ6RptrfRi+SD/QAc43Z/KxiSYBEuWVbISAuuFwAzBpK5XwEL
aMEr/VbWmDgss/8RJrHMwUfTozzkgY0G7y1tjCjbwmQ/TEJ6THa6FLEjTp7AxPre
Hd6ZnQOIuv78mN/YZK9gbJSsrW3XxoNeMeJHiC9yntZ1ip+R15cjtOPnUpbqrcJz
o2uvlGjfedVo7Gc8InsB6SS9YjGHN/VuRnzs9qC9ZUZC/h2xMrwOSoZQqUVGr59u
`protect END_PROTECTED
