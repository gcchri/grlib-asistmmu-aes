`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
839qi73EmqL41QOP0i0EmgMTQzqCy69Es1CaDh49+PcgLQ2KmrJax7acbMH201lz
jS4gbQSnAWU9c/ENWjIyBW9kNbmvzId/jHWVkDzjepmCabpDP/h+vc73Ns6Oh3M4
RO7yam0CR76bIGJgGtMw317gf3kAAAHuGBWugxdk34LDOYdhkNNdlC30eSy5NIxt
8HB1/qrrYU46Fgx/1pa3MVj8pEMDuAYtVQV2OPlYHwQEkbLRTO7zCITKbh2x3KNS
tUy7CxU7ZoSnI9JLnNeBAO5+q8Ssm8BA17/qPndCBwXxFwsqA7zh57XTs/7xy01x
KvjUF2YL2/COmwWsfFyUAk+9s2bA5j5Hw1LpGeNkBHEUZX53n2K7JPKegswr9lKN
W7dBMbBcMEUq7mGifWjN9Xdq0Al6ikhqm7uLadNemacggsDktkx2eMKnACOXlnjN
iYO2KDx8OtaB+H8apO2Pm01Pu/hNJWYfFlQf1yXxOOmm8E4Kv6qRPMVi8OmjjVjg
A3KdKF7tSxyLL0J0iVdW1Q==
`protect END_PROTECTED
