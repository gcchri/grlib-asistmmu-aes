`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
utPuPZaAriJ+CSgMyrLvX3nMoZnvVuOhSTOa1ubpBlmwj6kLTpVeh/l2fsJ8D+bf
up1jQmByLRZHsEIyfTL+SlVez3Znyoa374lftkZee5RTn0QDfU7sPrtu5GiYtK8N
sftjRx6kXprkXtSC6vt/JWTaw5sUI/etCe68KGDsUvMLIFgdjiXkFio1XKX7MXoc
K/xuElTM3D7H8EN1007nHbKP2SCXhwxY4iL8Y0VB57pvqe5k+NyR/b0XeCFkTVcE
4flWl05X086U1KjgYTx6WWMLCD8nTFnu/VxkI7b+ReIaHUhLqNpp4QIA+xq0ER71
TusdTXmsezNh+y8atuICwRjJjQpijSfPto4w1Ddkm2y0HonO+VSznhMtZlOqnFrK
a8lgDOApkTv2WJ/gZa8WWEDl1f2t7lwNQ2tZnELPN5nkBBa6GrgEnLLl7Fg5amHx
gyJE+u9PE/Itfsi2IjumGlVD8MI0v33RFrVFhoFoMJPSrUhDt73beyYrybR6X8qs
bFHZ6V/RPJCz7Aj+uDBo8gIKMHdUt5WECJOIVqEvM1UFcSIfemlljm9k0ea+8VJb
b1LUKrGkgS5Q1KmLw+3ppGfD5PuicuakjEa51UOcKxvrsi96cLNE0SfQtZZ7vonW
eNiTMsPiufCD8l3rrXkMH3ZwgSZDUEStk2cL3YEZxfPEbMKlg4yQyiz59QwUR9LB
4yUlcWl0rzaAGT01WifzzakozkmdZ7sQR0EoLXV5RV4KXvI3wiX+bVGypNfomh0o
kzx3tJQs1OpKjaIsZPkIRk8ZHHD86iq/e3+2qCHbbuhtbCkTLSjI8XaARnMEAwUD
haAN4xAdwDZ2GbQH5EffadeoBVihjcanC1tNtHzpj5+n6++AQ+akwmw/eIRM8SBE
q6fpbJdPRDup+zpAQK2DLjaDVhooKMUmD9BuoV2W9peHwrVGSVI29D0H7lzcYDwf
GEBl/Cfba6bbCsRKRhYQg28t8OCw2IvLulwUJz+oaD8fb0cYIr7GtPzEXrNiM3Nf
+3L7QdNmRxYBQ8Vb5TlVRMXLof/pTYyul2JIOeuw7iGh6lSs2wshNLcPoCMNBwI3
T7MnkY86JUM5a91NXwtyIeQw21Ld/79GjWGw5Dj1NE1rOCg9gSqJqsLo48E7qPgy
7NI0GaeyXF0ZS6Kt9em3tJSd5S/zLPH22wW5fuZbC5vXQUzfdq7IldwBzTZ+dFgb
y1THRgpcjlUtuQTGUxF99kfMg8ADYMTfn/HtTCKUxV9643GlZjPZjN5Mi1UdjT/Y
KO47SC0DWVY3FMGqX4Foj7epXw9lVew5gCUWyQ8zozdYlRlyMV7GydL0ZXKr1usB
VZzm97Lyxrvmd3qdJVA8tLHRLJL8dZ82O4mllxfRe4DKluYGyI7lnsxVM4Yl9Kyu
bR29tsbuLP9TJV64al7rz9Gzu02j5XbDwBWDkb7qPVRekjOxQ4BuBzTr5fG6J0BN
D9iwC/hoHtz4JTZey7VeJs9ey1FJAQpw09TIdiV3zaFBialZU58JPod4AJCLsquw
13/uqiVnzCzt3BChxVC2bAkA0iQjAtdWPJ7o6dme9/cU+Tq1c6Jq7QlyFEIurUdi
dI2oF3IaSD/iOrCeMEK1YvzZF5vBqpy6dgDZinWesCpeYw1ZYKLeEvuGFip9hN/T
Vm6iB/VrMts9K9p7VrGipMFAIgqF0zZCSlkHUS3vRChuBzbqtnO6PylEHMfUDvQ+
us4a6CjtGvzmbz4tyP/x0AmncdJEfmkkLmnDeOdGu62sYPjh3SPh5iINHyb3S+tF
1yHWbafThc3hCDF5q3eFL7paH3LSl55YNoRmnq1JMCdYlFtK9/exRdVwoZz7WLZZ
2UolS57NGrbesCm9IRoUh1PazwIdZY7Gaxkqb3EnHcuL8MQfjmFiIp6yoP5kAcI9
YAB/C15uyf934TZmttK+Q4bRlMuN2CK134mJ/bSvSasooSJr3Q832BPpBhWtKpjR
jmQE4xrscZWYrHJiHnZ8Bj5mWpv0HMz7RpRPr9ol5TNCX8tCBpdG5WRs02T+oYzt
OYPM0RPDO2rzVap1o3Jx1N7Wxg0zg6arnQ7jFmi+cvKlGYPiNxVyYud60tNS0J7/
XvPGpo73FO8Nns9TcRXma3hN/zV7kHq2P/nTs2O0aJVnxVXJ4z97dk7EfDL3WNyP
sD8rxhRflgzvTk1bqw/PNisWMIDpCK8OKu3cB8nnPlF4RRX4TPkRqUzNOLhcqKFg
GHvFzpT+fTtUWxYmnCUkcwP+fEqYSiRq67sKKrhWcbyDE5CgHW8v98sW1UTRC5UR
APCYG08JXdrHbQg3TJV3nzpi/OBdbclHD5mkIekQJnyR1Fg3auM2kWfeeLsaY5Wi
l2g3sKBn0ptSpZ5oRNWwbl5Jyu5uGajTu2+VArojR9JCC8co5C9nkOaML9BSiT7d
fYg+9+zGCbLUuOfTftt4NHjidDN5dJPE1oHo2FJeYODbJ2jcY/P0dV49ST+IyZ4N
dZxPsP4W3OpLpC41aeXxZT4a28DZB8fAaquyVWWlkAK5ocdnh5mLJzVaH6YVWKCA
6w7ry5UX47sfTE9nNCuMTo830vzjsjtxPDPcu3ZdRl30OUj/AKltJCXn7N3RbOXP
kfjQMPmtTXKUEJshdlgzaQLtVIOR/jScqjMBhgXi0AseChUJgSlUfwFDlbbob1dq
wZIAW/OSqruPctcp+/5i9oK2Arkc8CwTflDfK9/DWYuDv9D+gGxx22yj7IUk3aQJ
/0SUQo3IhH8Q/7eWQzi7bsiOQxLcAsfLhTFD9QXq5aOF3HiEgqDBWlVcxT41x7MH
2+lsZfwrodgkc/MZ5p9N6M+hYnPnzebNOTjx+GzcuonGOYLFA2CJaOtFkyxZi7oT
uo0TtHsjB2bUpb+t0qUA312GTZen4aLSMJZ9wuaN5yQLDb+JxSG2iqOj1QYbgJJ9
NGtzghZuZjH1A6i2TwQ6uwrvrQqPJvREG1rSCNUMGK8xJ5yq4iMk4D4AJGePEwdX
bbTmZplCAojYYihAy7sX+GJ+rRlP4dFAfeSOx5sTXpk+jpZOQwu9M6xI6HMTc+cb
FobE/ALzgUyr6V3TLhBo3vwfmRJpRHgbkZjLB2cVIQLYmRZLSa1zxuODnwr886Op
JR8Y46EjPCw8ZgP+vfv+wI6UdHyih9SMTd1masuviMLG93bgtXkmYGHH1sgD+Qci
OUseGdWAzsYqgHeSwUrSXpfYYoIzLtaGoyAgFTMiePoarPhkL4d0y4JFKlYLVsxW
TsDcVFCGd/7UVBidkkCd27YRaKXko/5aoYKse/HyZRWLcbog/GOik5UEM6J3uG5R
OKvKYnGHzbMhZ8trT3Ko4SwPpEhbQuMaPLKiOkrIDZvWKXN2g9L4T/0l7tRCliTr
PevI/6XpB0giRLtFgEMgoxwdRAD0B8QnRblkUyF9ruG1pzzcD+q2PDnWWYD8mlPd
nNZkqjdkMxh4CiJccoUG2HkvXNkt1+65NzgnDhNDwYZE8ZNSjI+XnZ/pKq9l+FUk
24VHuUOMA0MeHNzF2Orq8I+c871Mu0eEE5j+mDK13XBbXKrs5I/IZuGG+6mx4KiH
Xfbg+eyKdb/xfuT0pAGGl11ubSVkWif6/xbOBj4DyA5XRrbAiClOpLfOxCHOMlfX
ITDsnt7RYz/otsegAUcsV18W9HcXYmYEJQYP3v20eAKWgyFhcCCeIlCHaM/LxOSl
fTuPOKumkVGE+eqcvsSQ2vZ/e5XutysVdcE/VpbV1Wsa1W1LV+vj7+rd0EWniqZb
6y4+pAxtXkWbgiSBq4PzOw==
`protect END_PROTECTED
