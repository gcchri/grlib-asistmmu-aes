`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+iAunpLdQwxdkVVM3CXVL6bnUxfDfliRC9g4AETjCEVgG78uOU97N/sesjJNEHUl
9lzuaVOZjF93krqO+iXmYhSxOyfnexTP86xImO6SNTi5wbTFBB+lXNMGCJau6OVR
dzicxon+Rq1yIfpty/THYqJw04xgTZUUURUDIUz/CJEsAnryUNEscKD1CCI+gbYD
7q24Jp5XvtqN7I8odR9XA5TEdf04fZbwDHDL4geALfQhe/a2s5lp02/dYZw1bPok
aueImH62x4V7B80jN9ZbrXdR2CYfzAkzd+EB1B6MABhmaBXBR1646lC819itZegT
N35CxvT5MR/bu6kH23WsLI3pbJoUJq+ipNumG7QDBajqEj4jvbvcKAAGFyZ0FFy6
lqp/+MHiMNCPudV8uWbfypZfRT65zXMWOkshfarPHSswFMFxK9iDf4M0m3XyoWtN
kYTEZKOEHIkOhHZCtiAAJ3LDPP7Q2FdQGa35nL+DZqWaPby7XKbM7JOBI5veZOVP
1c8BACv2xIXf9Cj0iBPTKe85VZUWRexMh5n48DrQdQ0yNKSPsODbyCi2cokgfTyP
u3HSv1YqaLKG4wFRkrGm/MU8UswHbYCg+zfHCHaYl7waTdz0eiZzHTgPe3yzMqWf
ZJc7s2ajSP6+xgdyi3z4P+Sr6IedwY3zZRjfnZ7pTRY9HwmBYXIZWAPhkFOt0N1X
O8AYJzF+oJf+acwxaNH+GZ3oaCre2+jEmsqqPcJyRIF5nczza+OIsk15G49CCbBd
+0BPzAFkihpzbd0dMxxzvKudctAYi8hwokGrjYLtKU/gA4I+VZETxyuCNifjxe5T
hEt0GtXRh4YuCMfrjo6W5PovXcbdrMo9wrDYWCubf6UCcKPqnEM//l4fhqOTIJrz
l2cuZbUe+SDzZl4drkfQELG94k85v7ppRrdpcVjguEMT3TIXo80IgfP4UV2y0I8Z
d1VDuXFIyIjyN4RS0CRrtvUzRy6+eaBAxVQqiTHoKIq2ome+fyDxg8LAm4PuQ1hv
3nPKAOxWzxMsif0Cp56CDifGh8oSuOcLmoQuZufivHx65cvMimRaeaP64iPXaAcT
dyE/naYfxQmWjQ+Qj0hScYoqWfCY2YuEHNXHOKxUHl+y4NJERO32eSx0YzjAXx3F
D4V/vS0cVIarMfnCgCR60lqRxNuxmGAiesWqpYnSz9NpMDx1U77r3isGtIp5AeiY
OojmgLyBZoNvbEXimcGpmTEoje4b7/QtluCGIdY/LCahp1EIpxWuoDMQ7TzXe8fo
RcWHGWx42Vj1G0huEoOGsnzvIkd5H65wAk52COtuBN4PhegRAT1wZWCeKDE+OvM+
WEbYo3rfx22K9Z4DT242niukFXt5EDJ/mD9u1YWzJYEzS2BQGr3ydDvDZrFSBntL
rxyPrheMyWjl4lnIaV52P7aMRrCVOZg33up1Cv5IMtoSFst4fOXlYMfcUrurXSWT
pkSNY6s9wpDiCGB9GXZeRU+uDnVmcmD2DkA//5PEjIZRbklQH89l9KY9Izgl3jJF
SW+7sXv8UUdv/OWGogyniOOg7v67DvCsvCHR7xpYwlHnlI6Qdo0nTQH9fV+OYNip
8c73Iz8voNuhd64rXTndhO/pfe/KhkR41Yho5jGEL+vRcNd5B8Tf6xWOa2uurrWD
BovBTTKreIec1f8uJgzBsDIcYZkkGmcLx368G/rODehRBCmeCcJ/EGA+8B4wm37y
XFx22PC9FofRH1r2XlEx2yifZ6TluV8yANonDNwl1kkC/uTNmJ8OSzLh+BEGgUxm
qV8lvIL8sGCi05EC6wV5XRx3kAZeCitrYvTTxfiMCmgI4cADRENY29Tfmdf9ETVW
PuZHJ+SPiHlNL2BlyMxuXJgtocTccG8dgu+uaol3dg8V5RPIZhdNq4pyTI6w/AgP
qC2hpGmObjyHIz/gjNPW4toEurg2UP4klHfbOjJ/lIVSsR5+Wv1er8bURHydTQxw
ZZYR/CSneI6LHbedf/o06Pk4FJ1Ba59kEzOYXtpiD2CGw/ESpw6uglX+73VLSMbp
gPbebTrKib4/udowBMqaDR32HgYX7RAyxAK2KjHkBZZaaDoRO3DLq4J5AGS02VJh
ghJ59MdtlFqqX/v8vWFzgtb+3Y/ZgrShKnNc/4DGyKeFmB4lHu63YtKIHr7fx4DN
BKRAze52dOxHPjjRcR6EhlSaBNDMyDt8BUuPNOSMYagAX/rQZ8JctixduB2EGq7S
Go67U7GiUcaMtRUh2ZlHyG9mjTLx21ujlMvxU6evwcBeqzw6RaPzOtiqQa0q+/Gy
Za7tTSgU8ugnDMP8p+S8Fl/sodQW3qmgonY6sU8I+hQuMtm+bTo/HxwO1LlK9yYQ
Kfa0a2EbDiiR9yew/DfwXgnuNYw1lJRpdH517UWJSAjAgVDOlYqCKF5xAkmL5XSD
Eau9RxqhpVnh2vFe2oErDUMz4jOOiGNjQBgRy1jpANrItuRAmYY5L/Gq6Bf34S/g
gstgVLqPF19iZbbCUcFMSPT7Z+Hu0xBTlaUDLEll5Z8wJRExfkulFm+PwRvZDBXG
C/zGr0kpxe/n+0XULSICJiudWMejFXwjyeeTjLkRw9S8vmvypijXawTudSIt1Ijo
TqPHjHXpbexu/JxUrq7QaNUCZ5zHgW11TZEUr7Epa++IYulZMxIIMFeakVqLeGAF
zYoqRyjgkIxLYcwDbVZNUUesXS9jBQnL5gKT11hnFufb5JX8v9ex4POgDpYq5MZ5
ItIL2kAqHxSKEuegR//SDROFfoVI4OngW8ldQXF1r8GeTWm91+L96eaaT419QXLH
ed6n+8GVQEuvdmtmm0MNy86tG5zavc3nKSDIfZ3anHSlFYuPXXecI3X/5MF9K88b
HxONV/xHXvbWIFi00XsC3NMgy1bDbsOyGL0gZmQbNZ9dMOJD3xYeOybhNbuv08fK
YWCz1NWBFDFQOa91hpX9IKvodSH/tbKto2YafpTHEsjERafkkICcXnnnDbdPPwnl
ElzXSk/FC43hYmc+C826k+uwjIpaYIQLH5JEJMx6eFOYbu/ezi2jrVNDQ597zHet
pmBfpqI7ZP87nVpwnZwD/xZ+oHlW85j3eTSNrOhv0SW8W8+W+acvFDowFk7gFyMm
wkO9j37KCc2yQVhaq2OX4RjBqJAt7aPGBI43PWVvCRouekXjPgRr8TDUKb8zIYpn
nSEoU4a1k+F8IjKFPWbA0pfrNbq8RIllIeBpniUyxDWd+gxpujsfSifF2X5LGx+p
hEJLKezLT48hMj0dxf8+k703N7RdTpTNncRmeCJYmZ48ZSGRH/l3+6NlsmOXNN83
DeZQVCmGI4pUU32YbOVIYxKEZF149OkDnWBt6AaDJn6J+qfiTcvDgopI8OkBvEOT
7HMhbLAelxthZ+O6YQthMBQ2i8BiZks/7M7tp+TGiQ0wNsfF4qGGtRQ8RG0UXAqN
coDyiV81OvzGXT+xBOnbMLgp214porxCxFEtUJWq5Hu8L/aBdX0gK6pDsAHKdkyh
NIa7XcUZSIY2ahSuhxDmPAZkNznvZFJiiDwkjWW0RjLYXbP/pbOyqlMcLpjPexKa
VSffvGhyZcnx3FNQspuj+/IB6tKWubvyy7ZvrCKEzbIUmOuobgCLeuqTRZxvNren
2A5Jk+QNGNPR75IyhSfHJF0tQB5RaCLMxr74lLSeptFcO+ltdmnOQO3EO8wi8lHc
iJZJc/+t293LfdRNmLbqfJ+Q5Jx3igI9D/ly6KD8TukmzhV+dqzx6ruhrNuxh54B
xXFBNNVccSaEgCZadsZ5psGTa3bxKDBmC/wo4DRxtgAra3Tk/K4EutTac52jP1yR
FT4A0jPnzEkt+OjX7tqxr4fuBvRUqGB+tG/gcySXbydDamhoZvDePGJoZ/po21Eb
Msa+uUofeqjygHHX1m/5dIMQBY0M578DJ+FAOu8NLMPO1ouQTtSPfXbNYrag9yXx
uFA4bPXKrHiafy10Cs4LbnQyycA6TDViV/sJjNDdxTMW3aQdXW/Nvx4FVxycS0FL
/z6fjQJQvTDpuaBWv0D1AbGR4QEkyfcYf28/+fetS5Xu6RkQ7j9UsJ3N86yFvlR0
mdCQBXMhXihHvg9GKMzceDZ9DU9S/nsnpH/Z7WkT/rinVfHrQ3x/axy4NObPNfku
pXJSlzVE3ekHNqj5vfegvvoBR7MPDkusREtW1TwrTxpStGnjpv7ZivblY0qQDJDX
7giV7WkpN5S6lDtBc2SBE2adH+iFiBLrXUdZFMNZDmoY7ECPo54IrMTUW6AMngDl
tD6EvIcSBX36kqVxufId2k5vuJs6YI2tEKn8LYFcBboWOik4YfKE3k9sciSvYxqY
01aQYBrtMG68V46R1MyuVfoX+fwnIe4GIpsR1vUmj/HUH3nyG2miNYppR312WT4n
/XoP+Wl6Cxm0m5sXv7WyhVArhczg60creladmpHjzmQwMx3yjDtDiIBO9nba1MRD
3MJKzaaGy4So0/USJ/xsuOcRVUaEgeab34KT5Tp4SPo95Vy+jpVYfadOHe5g8Ts0
pJJ5JAXV/eBEwvgfhlDS+b+3st5c+wNigs6AO6UXp51G71d5WbDlT8pNSUzRyk44
qmdRKRXTFKuzks1zhHPNPjPh2oBlDehiTxjnxosQ+afNLM97BWKsrRrZIJMlRjW3
QLO/+LyScNA2mJOOqbvISz/fct3V7VDMWfC+tmrSLV1/sqCOU0X/bQV9e3rJko4A
hTEO3zh9HvqbCfZalPITm2boLg16K5Xl4Do4T+MraMbUQdKwgQKnCDGgDzLxigUG
fj2KYws166wGxtR0VDUu35Z1zg3NKRElEAf6Aa9upnfQ3p0KiROasCkqA77e4N0K
jMUiWDUeqNfX0+9ib8dQL5Zx4eSrqsQIecQTopnMX7e3AMw5Z03cEPity8re9Fon
96GMHKZguiPjmyszJ3irrhXdy1pe/Z2rstT7ldeQAMc8TrSkY2q6iZMCIJuOJ6xu
tPJlxNB2CVSsXxQcuu2ECCjvsr6kHchtTrUXwD75fKWbuoeti6Em7kIlAKcF1krj
uzTZng9T9L3RtzcM5/ym8SEWFFEcp2rlweP2H6vrdOMBN8OAEpHYsYms/RgjyUxD
8tvnIuB+fK7TYi8P33IiYFU+0H1F2gDHycgUE5Bh7ceeZGTIv57cUCvzZBQe0hZH
bHo6TldXuBbykTm4lVEcYnSc/VEUCpqhSp8CIKgyf+L2+oU0jRGT5cXbOr2a5iZ5
RUQjiRy9OkefdOHRSi3jXSEDWFV5ArDfieaP60nkAdPqS3tVAUrhXniUWuo8lEl2
eujr0zP37sPgP/bo6DV2CvafuQVCggBJATIxNiGb+Jm9TzNvoqez2P15OZIARnRJ
tdDFuRl+W+1h1V1tmeLVnEBcE6QUo8Zy/3rvXSi046JwBthZ7AXRyuFmc1sIKPHG
5iZ4YP1xZkM4MKaJ2/+Gl3MGQ/JHRWVbSUT5B6p8G5xhsOONJpHOT+lMt0g+7yX2
V1t7qekNVW3HwpU1sC3zwj5DGtxIu9pz2J7LPr824c8+7MkMvxtJy1sk1LsPA8aS
QavNcBY8jEOlrSPYj6A+6HWUj3lTWpxCc/JPRBVbQHMegPKPGaE2jtPl0g/VSrzb
tP/E+njj2ZwqOKCpEzVgtjzNCOpm91qBV4FEZnSzk1kmW7AP0hs+4OViP+XKdFLk
cbMtmHx6FYkclJ2jBscpYM9wh+a0k9epCApkkUFnES/lI0QPk6BjooR1ciVjdxqi
2TVNUI+LO2JEmbCQZlVT1We8w2VuSh80IJHAQQtKhfD0lLfEDPdzlZwsBzQ341uq
4NQs58jjoUIKO7aNQuTTqCduQqG+4vliEA2CTeTViHkhA7iG7TSyxDY8R5LcCREq
/pIZXD3cxyeJBWUzO6Ct4vYxIOvCyKUxie5EYeThIqkEOKM26+njUDkQLlrGlWQ7
2YtcBBcVO1l681SaCSmCEQhtI3q+06VbajrN1BCalvX8VDXLjXikkU0pwfvGYQSV
ElNgU/omTVFBfWi4KDKR3ITXLQjOvp+TSX3LOqHPiPi6UTYYxbj8L8uLl0ghbNVx
O4X2T6ujGWNwli3t3eliva7+ueC7Y4yGP7Xb+MbPPZz66LldTAdHe4jvLZ70Yrqd
NRUmZ3oYV2CwvSCv/4qNGKb88HBWXxn7MaJnWzbqNsx8RdbsCtfYwOhxS39qlb+S
pp+f8HVUuVPxJHKkRK53C6LLbS7RoRvn6Nf7BWWQhQKLX/BUsEXJBr1MbKTXxRwZ
Xd6IUZwsmXourGseEheHm9glCjhX0xYMBfk8y2l0GV/TDKgY+wR202RU2BBpAm7X
7rAZPCsU5jPypz6L90amCc+Yt0q6JN1aGSxFRcm9rvANlZ4sYGgF4lcIzcXQfIC7
tpVK5RDYMqTzcU0E/d3A68CjtiuDsY/MJgm3YVi9KZp98BMZboMs8jEvXaE/a8tQ
GxCnRNST/3u9S/xmsY1VyFF53VPmmWU34UkuE892EKJ9KmOn3uhNL2yVDCBGE1HH
QOpnicroUZDe6vAUrkOIKM2uT0TCGjQK1BMpdijsPDfASobpvJs7FqIqsjmk+DSY
oRiAgHpzsbAiHfpCnV5YFsxrTXX3NF3VU5ngWCxy9cp2IkVwmGW8qjohfsp838PI
yeWS3mEX6cdx5v1h3g+c7fwdUu/DLmPydS96HvJdxLob0Wv6qoe39SL/afVYRNnS
x0THxGFFp7LP0MkyIXagWal+RcLlqqTgAoGn1MnRlTYLkUNBnYT46oXf6kOwHZ+/
u1BZHCucMLQO2PnynmVdfrqnT6eoHcsTKgaOdUW5IlokbsuAlF2oDWJJOfXRSxJd
VYUBHUKV26jVYN0UwfNGWqqwARILJiorUKvI/q8L3qudo3XB4/BWaQYOPgHzajsE
akdrlCNuMq/wlXlZPF/ZA3+xrV9AeaswfJM07n/TSQhdnWbEBpQm1IPHcTVGJopu
0thfTRUhT6IXDZQ4WSHpjexLzxZt7hEFcpHKmY56JktjSHJILVEPQUlO2gUJRmKt
Fi5pBMdWdpXYv4mC1kkOtcbh2CjmXBMpAs1qcag5ISJmz1IBy2pBKk1XUmGw+OXu
HA3DOtZbTv6nzKLMaN01/JuK0j0+p09/CLXTOidpYOTTklbYHIknZJNmzKLDiXr4
SnBr485Xr5SjUkzWkYd9V76Khkg1TxGchaMbV+kMpc7GkoSKaOvg98FqWvS0VG/z
cps2wLv1Ri5fCWSbYRB2njL8e/uVk29xtI2+tSSlxsGgVvVh80eFxnWiQZGHUlh5
84shtnpL0trr9MkRVqKJH1RriW0yeNREvFcJj7xKsdWNwHRlQixH+RbFYJAbfyUg
5RpEGIbS5ujBN9hOLxxSEiWO/7v52VGnGteY30tVdvd0OANJU0S5/U3P1c4jZxHt
BvXzzoCuhnumvveijI77KXJHTsKKuZNlIUyyLkC+ap3dAQYn4/cfdhvLDUi6kS8L
sqGcAsz8YlDNDCUnE4NhPqafvrOABO7ZqNHobXZrKdkStZmEVL5QDyNUP19smtoa
5funCLrby82l7RhPUq18Q3RB7NQ1n4HQIi8yzKIEzbTsSIMJinEpVsYYxW+O4xTJ
7h4OYfDX8ZRuXljU2I2j8tL9Q1N5z10h9wrlbahxHu1WuGD1TIbg/dsKazP8HmxW
BfGUVmCcqHcgVpPb0FdebBhvk65cTX4aSmuW6cEG8HdC94+/y149PjHvbijbGmsL
e6WhYGyf5jI8gESJWEDhylCxUIPDysUuZTPNmGdvVPELEHoEXqTQ1efOpSoqAoxb
Wvrt1PU3YZAmtbqes0DRTytV6roP45YpZplRV0+k1/YPrmQih73IHV+U3J9moqI7
956gXZMHzD5/t87u3NCSU68x/w722K/niwtJZ+qpIUGHsRioVGGuY0WWeo+MhoOU
id9KsBvdCvCuB6RJpzs06J8PrJbYHyZc3tt6JG6T9peOZ1nEhx6TtTNtvqqtszIy
3BlhDEsPgOwwRTb/W+OB250tYym+8vk4LmoKzMcXxaIOtsJQmo9URUva5uNI1X/b
YBQy0DLm0WfNI8MDMOo1gjnQCNRSO+XpM3+fNsJbfSQeaEz/GFUi64GiyFPv8i6m
zg98bbiwmNHN5k+12IRfKT18VlbVrfr5Ms2w5XqxW0P+veDEMcZOdoG4Pu61VmKt
L4m7x64f8x7DOr3PQhGFoMVxqd3crkFFNLYcT8XYL8cA+UxJym4RPe/+qHTRN3uR
Uaqwbj7SqrdEEcOFjGRIuSXGNrtiepekseQLuPaikeorHJtPgZUAxFqOc+dGAwjw
RtMP1toiE9rLIIumWzPryNpT4qW1NnZpQoKn9cPffIz92Q46W4ISJMmyM9lW5ywb
JQGJr5nBkcsYDv4my9X0v2YCJTeyWSUph3GndspeE60SxjOwwM9BlwX+Jk0ubuhK
a+EbKWVCJvPI9fdN3KS96SxLKtl9KJmZXJZ4CD6BEDsQnYk+4WKkM9VLNM+QwPMQ
IG8mmLpjf6v15C9mp8a6HMCjTKXTCOwo9NrH+yR5e70R7QbvvBec8kFQECn1aQ55
ObSGIs10AfXRKn3mnu2JJplfkBnJgnBWYzKeN5oKBx8EhWTzq5XsACtz4UPEAcjl
hnnlHNE/u0RCJUNgXP5lNPm3LVQ7RdtaeXuyBUfCxkGt77267GQ5hfn9oYqHUFpC
LyyRsDx80TXBgM5Jgw1hmWhNA9/mLRiybEb0gnFxNsQUMKmIfjaMFtqq7OFiKEPm
6d2yfPNueCX/KcXb5CPk13mKPS6SHXK1wa0Xst4eludSN6kHrn2WiadRzm7l3tQk
aLum19Xg7FpYDl0e0NKPmq3Bk18oqkEFR0GfFxTXow7ecYQRco3h7zS5RvtIhEfC
lwXvt+0VGu9ZwLfyvnf60CBxDl3PGPRvumH0GK7bQw5AiMpL59V1BxHNOb5mtQpW
A2xgvp841uE/48CsCDZbpdl1mCsAhITa8iiuL9dbK0Ty80Q3IcD/QsDU2VCBbyEv
uTd5YUFjjLkw8Txl6uWVylga0JgP90SIVKDAd43a5e1V3KjrVnDJeAfZcj0Oq/XS
56WocUTHMg9cTP85lGNCyrcMP+ONNI5paZDglK8yIVSmPfzMYKrWwipFd0YOsFxv
Xj9yjI45+dhmQORnEoisSloZdK64cEXZ+xPP2/BTTWgwF117OOJOEQ6VB1nQ3Xz/
H/gAwP1DtJmNQ0KZR1O6Yb/hFAMTuEMOSseKyuaJsdXsobigyCHo/OxM+OhfL0Ch
5vhAI03OXFkTdCu4NSuGq6TMIJeUCxJbJmgDeGZmZ575tOtWcw9/T9MtNRzMymNv
BTrRHc+kIPRXCJDp3HR481EfVZKleD4UIJ+BgUL6Xu2De7WPm2Vd560isfU081dW
h+YzgKAtqAdOklgwNtwWnygksU1ZPlpCCJ7S6pjXoUex5b+5+p8NostMTGmZ3I2a
Re1G6ZcTkCZD+9HMyQG6TMdg539WLDfda33d2o5JDJou45nb3UQq1JsHdJa5a9sQ
E8s064SBr2jNwneUh6DOfsKdGn793qGVroPeXOv9vNyKE6sVwt6p6qo4XxVWCPjv
1TrbjWZkp1Fo55VF12OXpY9kuKggYtUPjx28YY4fX4PJo+T7wExy/Q+gadJ6qtnn
0tDR3+XSEQGDqmhPdnTCFXlChduTxUsuzqHldXh3og7qTqChqVyeA/lZ7uv75OgO
S/DmAnneShOrvx/pvIAmQKbUqsf3N4Pamb3KFOUzoMVePHJ5S/9oL/DVfX7oIxCs
0B4dBtusryIr0fPs3ZFG3vz9NiOQsSOFkT2vssJkhd+cj8+BjDjY9Xy5Vtcc5nnz
GDuw5AVAGZTHILrvi6VtH4fVsKFV4xkekG4nCNVc5XgRNFGpk+IpiNWCWEr9gYlu
68ipd38ZKZTEQzDGS/RjA1tQG727YHCfisIM+zDR5OWf1XeVA8uRg+l5m6dY4Rpa
T1/x3SOE4NTs9Ytlw4Qs6T+9f4FpRlNgVsY09YzYavyBCT5L6KHNbI821pCG10ul
n8zx4tP/OymcU/RNMKAB00MqO5GZdSDsS2ZzVOnH11kWDItEhspBR/iyELDS+ZvZ
qTTG0nn1bJ9ZE5kgkMou8m8/qJEW2oFCPae6fWRcvg4oX94TPk8tX+uqLO1VDX9c
8U/lIQ8r8L5VYZKUf0awfRTEoi6fX76mUX+PPExQLd+/+exF2rHzK5iHynuYBfMV
/0qwIMEnIcV6qB2F5v7pIg76vNAkxkFpA+FNOpl1gsanGS1OLVS7DAY6Zf33pPx3
t883zGLIChp48l9iPmIZOjkhs72WkOJBQWIVURhWOcqUDB5gAZWm0zVBmCp+9Yav
vavpUTDFXWOlV6GRC0J1io7qSXPGkuOPR9fEY02ZAWOun6ugWLEf71JiwJ1RaVRS
gT/3q1rQRr/dERpuf2EzRzTGBOkaGayrLHMscwTjjPl6evX+MqobVKZcUJFFSTM7
9m6ogQil0XIp6/sYbzY3n2qO8Npc6AlEkLDHSIKhDpv/rmkiA9xIo1EJEoWSoj2I
RZ0hHEoyiFvykDjXkg5ljZBrNjMSx+xT1QIMYBmPrHentp4fRjhnFF51fE8/hfUF
3oQwyr5ZYsYiqs+wLrAzxPOSWx4CCoVFdQzxd/L0RKgoVmhjNJ1vEpDSFVx6hp4B
XygO02Z4GwPXXtvqgbJ3Vl4fc0cCyyE2x9uBFhk69t48tw+4+v9clIlCg3NfKlEu
3n6MJ40H9jao6rfTo0E/qqpAeAzVHUzD5VkG6hPo8J4iw0KAdURMgadJ+dxGnjhN
o/ZNwTxL30ssDhUZtq5XHM49uoYulaENz/WnNapWe44hy3RGjsBD3l0RohOSxktw
rmFv01R0rq8kto44aaZQNxUkfq97QIzjLuWEiXgQThLmQepxd794M1iir0Gf24UL
Vu3SkFxk97iMkLntKog/+M6Rf2r/ZAkiGn55hjf8Jr6jpBqZ29dtIohXvYOReu0/
3XSVcqeGXVFIsxF6ZLfUBFF3xOkqI3TLNRyA/Ajd8xA9KzsE4vBtbDyaB7RjEcME
n7SXBFeP4BUCqdGgVKuZiPI2AeK8i6Ye0jvaSdXZETKANIAQ1hWzuf2z0PfPSXZi
A4ik6odfM0IegVYCwJI/ahJYOHsOiTsOuxj0mclr8IEgLrBRYXmWQPWCFTJVAOHj
0nHxajZBE+qaeB7P7SzqwRGzZ+imaPvoTQ3O0cpY+KKYC/aJ4ebTyNKo5bxnQkRJ
kV/vrecP+1YCX4TKXdJXKJ02dIxKW9Pi9Y6ZtDRGyf5ukwndVTzZzCtvOmhYkOwK
7H/CxTukn5gmZMLCWTv4TwszZLDVdg7d+M57BFBcAUJMwvhc4PDePwgq89sCukaq
OHixCF5OaAFo5Z73xhpFoCS3iYaeebuvrdS3wj0rPWHOljofKeIOW54Bgd40xCeN
MS9j8N1wHpnSIniyjjsgSt4PNpQUf2RkF630t3i2VCQdl6Ro06flDtLXjtZzgGpk
a+BivyMkrSN2DBe67MI3aeuOSTLtOCvyfaGxbuRTAF1fxK+0AdhbtgC+EluSjPBf
V/2mTE4X4sG5nOF5NgqF/PhXCOc62FOdGLONSYQakEvO9kmKcBJglwxswNC5Jz8u
WLnAsag7lXy/tU3/qSMrLFcpbo5wu9ZCjhlf845j7fbK95kxXHsTJ0eALxntZz8X
kQ2OaxcYvA1ZAj3mVYAit4RWgFlUFcfEyWATAprY3Fs+UGmTx4QMLgwR/xGmJNIQ
DQ0nzxgo0Q/N8Ystq5zbkkJmqtQNt1i+q6WNGx4AvEUduun8Jx7qtfaW4C7X9U/S
LQIC8Q0SIN3JawuL+afsxdNVyHjyFjpoKvFnuL+dl13BfFjmcyPrKg1iEJohaAjg
YtAmItQQ1o7ctFjvLSEewCLdZSfSRD6LM1bA7hB7Kr4BNG1ns13ibewC5vEgMzwe
uKu9XIe/12ousj0+RYeoxeEeN/UBCBHIqMvCjQ2gxFA6Tvb28hupdnuPmFuq4oS3
n/fyTlgRnt/BkO+TJmaWT3jlCeqUPTVprwzYPYCyZIJWeyPoZoJUjccAB09dwHC8
zAUORDf7ocz2Blezao7PH9AqEqzkK3Zf1OFSGmmyw2oJBO191dMIJJ0RyTlkHBCf
LSfFR/wb2tskZdCX9BsDhx8+UaW4xl+/uWTwdmbuwK3twcvziZsPEyf9pJX7iEmb
MBH383WKqgmPxd3DtZBalsToelQO2//+57kPvdzqNYO1shGK4saEeHzL/yLONfmN
CagOofEv8aQ/TWP3X+U4EzfIAzUykCQFBP04Ir6tIhvr0mODTzQB4fHba6BDM3uI
xlBB9LpCexqstb/Ac+8j1tYnFOYnwK0yaP1vSMi8OWRHX3y98IFgHRPawdid1XoR
0kcv93uiBWtoli1BDOtVQkIdZvjIWRqIbrglbsZlgvGMtR2F3TR1o32c15bVXd7R
dim8LvwoLQrK1zGrLq/72gc3sajH/dJER1ECX/Mp08MeMy5mbrRqouvNDlHI3CeW
0qg/0bz3w5rCUyaBb2BPUTi+KHabOwziEpRw6ww9qqC4Hno3J7bKrfMGtISunfXa
0EoQYdBp4VxCQK+vOnd3joEpybxw/dqqH+wyji+4Q+OK7nREaEESxy1SCbV7ssHo
D2a7duRBOBCRwEODfBbuCfAcfY54s8J3gegGBWn2nYY+NW2dvC+R65l43gX7raZR
S0o4Wf4KA3d+cBZDWHhtDDqkupVcYm7GJrhBZP+MXM6GZeFxjotmKSMsxTpH2LnP
j5Y8APmfexyxHdCxPejcZQlEJmAxCOT1lrxBbu84/VHyqohGC0Td507E5MamhxRc
YtlgVRTGCHsO7DwV5ueYenFGyQe8oQ6L5oofsa2exhydabO1Pa9QzsM0JNrDzr9z
7vWzYdyKbqiYyvr6njChAfQ2liNMl6yBmDYuBYRiL5g+fsetpRJ6O7su3Wt0za3V
s7tlUvY5CBr4Xv4LYfXIrkQub0tV+EI/nXmbWvKeS30twXEY+IwVNYA6D5wSA/Qm
dCPGC4oeDkH2OFTHUQzeyl4prVKAYayJWQIxsM3Q/b0FvXLKsg6h/729eBdR3rAF
qKkELsen6fFRj2m2qj3S9W722NV6uEOEDfvnsXZNJ3XevUZKijzIbWJJW7h0Qi7L
yRyHf6L1+97O1Wv0jqY3iI5KJm57qmjUULdSyGV4tIPj3FQi/datgO3Jx0mbL0he
Zs0i5OSmNzgwCYfBqufsvM5xg5UFNMQPzlk4Nurg8gy0mOpP0laKAIElf8nAXsbd
Ce1BFlU4yIh45929VXCWD4G7BfUElkDWYvFse3qoUbYIAk8GeDPWa9T1TGi7Cqjm
/y7SBeeQyPA72ie5zVs6HYPzXyVzlZlOyxYXcDS83B2baIgdyx0CzfHcKclfq09w
QA15/yAXba1kuYI3fAI34toPsruWIcG+iU4HeUIKHfpzacEjH834LQEBCHEM8xOK
X0GO8P1Ovg3pRoJKvB+9xCH92ol5GhzMWgvHVLiR/eJRtKYrpRZVCqIei0q7DQjB
KcwnvzZFubvEzrJP1I9mXjw/UDTm5WnRcdRTarovdm0iwCly5QtBEz5CDFw8p3AT
2EALq47rBnu1lpWE3+ozZhMKMF0J6v8/aNKLi7Htae5rmrEfC3Q7GIfxmvM/eRHY
xKsYyL7hSZNSL3BmU4k6hfq+LfKKHkup0GE2SD1XOl6qxwJ6MIauxooteuuxYcA1
5LhKul0gHkSXhmpriM/W7uMwK/csfi1MLh12Jslib4JVbofxr6xHbOMunoPKRwJn
/FRB4ElbjwcFLub7B7JXv3ogrJQBcLgMquzXD+8y0BPlSVi2ukjr+X8pPx0uVSJz
8J+11yT2fQkSE2HKolScfsFixLrS5o9HSNK1Y3SNHGmghZuQQq20PC4n2QxUQctO
JC1zlgKCwXLeA5UPRzMr6BzedRe4uLCJ3k23ICTpXYLpAbflMSCez7NzAEvPGblO
bQzwi5AIAC5yU4rM7DQVJeCblYOXtfBQRfgeo+vi0b7xlVw09foJrY3gOAzsBRki
SRPD2XGqzfFNFqLk2yxZ6ZhRe4CZJFBJX+2n7fR/jXqmKa91nKFe4BPBH5GfU59L
Rv9X28H4nYcwsXuVbztrTjOkmQxrFqAxmG3bICuXWPI+qXm59leSSjW0uFuXfBsU
5D3S9U2f0xaLDrvuNCvuGBnZGt1TB/vzSeP+HGxacXGB0jK7vOClE07FUy+q12lP
4+ERMXDXvK2be5dwbAIzaQYKwAHChNOaC3e1bb4C4JPzQxWaER1uMpT3rhBnb/8V
zhz8XLcUlZHVOLYwc4GRzExVov9cJVspdMnLZ00cWxXv64NH5xFiq7GoqCa3A56L
s6e992/DJWTTYLJZyyJF2ZgwqIwD7b4b+Xu4hXQV6FJO5D5nXl1mmRTVBMI+rod+
HuZUZBTxXHN8ePvyeb9tMXRF+rqgHzRSVZUqjVMBrnamgxW/V7OY5iO35xYckUwL
onCV9JIPw1KuOpE03ZK8EHmOMfpSXl2TNIuWDErGPbxzmAdcw/1GkX4/gyGsNRxu
4c1b+BKZt2pa6UVeJH9jGkVHyo8xQ/u/RlZVSEkrHORWElNh8QILw3U+gRthLotf
NrbWeL4G0tn8M/uy0wd9P2N+PxJl5HXq1nCOulaSMSZwISqHT7vVHE3m1gt3d7NC
WwwYUtZtEAPTzvzHAuhJkyChNYv0oNzi6y2pwqF9GRirk+84qjc5skrQwWJ73BWJ
Uty/zzf6n/sxUPzPaqBL6y2zlN7AedhVEaKWpEFloEEJb0UsQ4KtzDMHBG3yyHV3
MBzBArLQDYupsNx45PDN9uc3stRtW69G3661bRc/ecXEFjBGY7lUMl5QsLx3IBqv
iz7/7whjtNEvOYhMC1ct9Sno1+ONz8KVHgSYaT/ejQbKGdNrPRkZxXaRjK6ugVrT
flA+hiGAinVgQvnvml+lhpsH743cTk0AJ73yFSexvCe/3vy3fN1/p5Sw5kPxpwUR
e0l9tYEHcGZgMPlT8UkG9IBWmeBeg+1BWhuSnO4QaipO4z152tN0Ts8p3equBUZG
SLJkpKxOnrxhGmpMvGEmzhSENxIgDxalSX1pXhqHOJaQA/y2nnIhGi1V/UwQU7Jd
lPn41nAAVtRomlCN9jCOs2Uf+P9RUmez1Gh7M3hKnakrqqLYeryYAI9pBlItfFy+
MQNtXPbKHVlQ8Is9YQ4rKsRSlDMB2yZWMeOmM0uxquOPGmY04uOr9QCxSHjFFPaA
j0J3zHroiI5GK8YY3sBCO2ERwlQeWk1NvEEj5YHXVrGJIhoOMpixerUZDQgYagB8
y++QhUIg0p8gYA7Y4ZiMpr24GsZ2RKYYZBNqoCfT7dHFcuGKwjtrrthMmTLJtUpC
LpI/hhmDqZ/JFokr1aBH1MYqPPJnRCubvQVl/MM+pdtEA6Qm1G4qursuHsLjRP5V
dCkxxo5KQB1i0zN79FjN/HkIthQqMTwr8pg1J0soh4rReQz2zoIKwzytLgsB8IUv
KpacWOCI013/8DU+QLuSREe3d94QvFtKF8vCQx0VRKkMU+K/NUtd0MZo0OzRM9Nv
NxhEuhsEYpvvZl58oWeZuPcCPv/TG3/ZEHjB/pGH8NebynTxJqKorsQJiRFahMDo
quml7dh1a1Dp+VhYZh4G6QE6PhCOMfTCtGjQIawHwRyr0YpKlytEd7WbXH58pbOD
Fa6Mq9NeEgTvHfEoRhwxdXL9PhOQ+g7gq72T1LifVy4FsfpB47rNj9aWAzZpuz0a
VJOYL46DPsN/Yrx3N/pODy9WxmsCQK63VVvX49eWTcY0rUiPDqGI/t5AZJ3nRmYk
OsuwUmE4CMgx+li3iHMbWWVEdkXK5J9RfQxixkNYgLZiJ59+XqA97q2Zb230o6Qn
rxGr28ivk3ZAArmBcl/jSN58W3oGkXAHZHJW3zNwv2vPz3c01xC+GhC5E7fGaTzv
kAi2ZXlKZSTmy0y6GKnG/CaqUJK5zcsYp61tD21AebtArv2hdYHDtGspeeC0JriN
JycFhXgLLqH67xCzVAhu6J4vrTUGhC8D49gVLJlMJ16fZexpYTF/C4UcKuaGsBnI
wUHKbCog5dPPZlTeMrrAmFtDUE9g/ZH2AiEb4VQWxzQv/A69bVvHY+uf470lsTrV
FCZ1qBOZ5uX95U1/R7GE1yu3MEQb8dLSGz+l5fgfA1W7eWZYWKohh+F+hygcNCek
eWsN1OYJyyX3OTiXWZYrWDQn0V2kOa6aJhSwlWSETeBPpmfwFgWiRtFJCwAJRFgs
Qozks1fH/XqslpOEe1SMOIDbiFMK8fIfyV3B/wAax0sl8+N7I0VQeo8PxSEVz3pe
Y+fgH076/PDR3W6wzjfYJqPSsL4vTa/rJRBL8JS7/TBq3tn4fWOjA78hGILkY+NA
9OGxENATCi9DNEd0getAE3q18Az/LHP4u2nAFAW/hNE9ihZoqrDCvD3Eus1c5OlH
cqUwXZKqetjSvxyBSsP8Zhna+yTek6CIsvj4KJx/8Ym1yBCV3nr07e2HTNasfBZc
uz77XeweOJeQbItBTcvr1pRWcjpBXQ54DCsGRpV/Wn5CtYETyEuHPQ73Z8F06H0q
LTHrkxDpo6R5+VTRqKYH/FvGZIC/poFaHDvo+hFpEX+tVw2pbEeKrFlMoTjGVqok
fv+UgVtaUENQMp1aXB0wHFs2XTOYXZUVLNaNHwfVQ1m9lqKEpvVLbmVQdhZZQfXu
gWs8DKYI43mXH6lyztgmlGj7H175bmuxGI/LDRQ/X5ZTYxIFum6nua/pCg42FioA
fxV5JRasNCTjB9i9lgL7Dd7J7vRMabpdY2Hx98kOWIOUvdKx7GjpJcz/V7hXD4MJ
pV5XTSnK7xNyO1zHtp3qK+g/4G5n64dVr+TTqwZ+nvtF+7qA0IlpYinOm77o5Uv2
B3TC9CXqErgT0T0g6kIt6k1N951EB1nAwbMxQnPRTYbEojj0924JgF4RQz7xPyXA
jwDOOUam8eGNV7DFL34z8YpH1otDgb48AV5zOjPvpQpH4J0lE7/fuBwBeAfbEx0F
NfWA1SAb41ttpYQ/OQOtU2if6RrzRWVoUj5tsSNhgBmEyDTAqEEqnQ5onjuU6V2C
Xdvt3HXefWmhwvFEdfhe9NPf+e484c6WTdyC+c8UArnNguA+yvpmUAGWEpfaFUnA
XuLlNHTXngqrmyoXFXoLrk2UQaqPJoF7/FdlhAZrbIDnmLDwN9xAvWVfRaT25I9v
l5jstgt262qD++tpTEUunNmKnd/lbjKJu8BcgntRrFoaBi/XMAtheBs1wHUIp46d
Ko3e9VRp4p4MEKDj4fIU6KhwXqwHfz3TLw83DEpxJ/PnXdidd/cZep4G+A/s9aLh
WJTrIpwcrawB0NGfEZjKOa7bmIeN1/9PM4Eh2Ez8LFKRe+6TLe1Qu9im7Rl3pPVD
7QO9uJayjs3ssrrxVGT6qFsWFKSw5F3Nq/s7hz26LD+KVaLjS3btNRzEiUz9ewu3
gIYMnx7fgNiDV/Eb8KnewaabcqgjW7f2sbFz85Ttae/uuo08xkMrMDMKnW9slx01
pzTmPwIXtZMHnnGlwEZ/wJWpAYQl6yY/xYlaei/7tiwhW5IyItycTsTbkAnllHZi
jTBV6QFtj7AcF83LGaftKil7emqCQrbBtdEYMggNMMa0UUdpBqltHlkMJyifvyh/
Hu5S3XBOHVrJmUtGsff4SaTZxkJiXw6oC7xirTqqV2z9UyFupEyw8qGYdL7cPp2E
lZhabzl2swEhaPQL8ad5euzRC+xMD+MV7X/IFuD+AqsgCDt7UmuTllJw7AFFwZY+
/fAkU1MBQKceVxZ/Hh7tjfPAgxd3OPG3efWoVdfQIU6PliL+b5/TliurLF+LSk1R
DhaCP5pwTEzYBDeKBLjHXNyufg+xrrTypZukgTZJd5cBjnqwADO/T0qKsW2gqq0o
AtSI95RjVXeSn7oA8raxjSicsTK5SUGVX1zdXxtylSHf58+nSXt6nRKW4FLUSoJg
xZuBZY7bMXT/SuO3pjmSpjYtObXVplp1YUzLpHqq+IMvZZefP90SZhFxrQqS66aY
6K4zYKC7x48d2P8CxvJSlRzyQt+/B5HrNaAGNFjEZVSQz5S/Oi9is18P3FZsLvlX
qkf+hvMGl6lRgaAwkDm5wPkZ97EuETIbw65rJcPi22RhqW4x2bDTQU+33TsfAGXl
p70TD4MVlmuYuZwNFhBZfqgEO0iZP8Jzi+/y+FhT322Caan+kVPaR7CZ0NUYr0eH
W288cPq1T3ZE7FUQCF1V5hw2mhwp/dAm3yuEXupAKX3qy9RjDtPvGtOknPcGOZRr
k9JTP2LtpinrSgyK2WbvjQtHtSTXIkhhAAMzj1UxfYengr3783Vwq3yWPCb69D6K
zy3GgJAweobTK0lFEBU/UrILsN2oQQO6Gzn1pIKxJoMPrAgZUyfCwWPl7p93VLui
81lEbg5d0JbHyy8XIpXyp0StlL/x7xceHP1NsiTTDIk+FvQCfyQYcM5UsuIZd46q
9CPwMjzlpAohlf936f5DK9NGzIm/ncFeBHup07JHv3u9ERC7NZ7J5RyYwudCj45g
9i/BjcU9uQ5dahHmgf18j1D2R5NjJDCIt5y7B7vPgVn3IvYTyoWkdam/h0hEibSN
B0Njr78hCGT9OrqVWD/4yhCFWhg7jGW0PboEQAExjeOPXDdxXusGmJ8mobgN3z01
bvSPhaZbVwEQHutho1MGnDZ03J8QK1rR4ZT+OewHzOqNagXIZTilIM9ZACbHyoF7
vjCfuFV3cjWPTY94R3Wybj7mTysYLh+odWChxmyLAVZ8Xji34SpA/kOjpc3OodJc
7u7qDLRNkYpB4ufG06HN+E1tr2xs0WNjXb4aw68jgSwewbUN5/Dz+2W6cpI+Yh+C
osu2C9rj3XDDv+wMHK3Hand9GbRr7grtaenqKlfP2LoAnSfo+jh/v1nGmank4sUh
Rqo649AcZIWJiqow1XBkU7VNgfONHJXv1SDP+0fQH0GSv/FVIFqV1TchGXLOnKOx
JCc0ixpl9onIpKOrTDOUaCphu/gJPRq/J6Bj+NJihQqKLPL991aFLOL9bmP5FSMD
/DiwnEpaopjfpqGA9TOZ8U0Tc/R7iAY9uo9qoDUTFRr5nqNmyk1ejj4eJBPybeT2
lqVxDrFlLXbaZ9VEGws8J26XYY7/pDIR/uj2a96+7vvN9npUf9qBHfGeme+z6td8
CQMoS8EdM3+ht/oNbu3G6NW66dFpOKd4NOxM73eGcHxKxytkl+YbYwok1pqLpPyf
fxaf/2cC4YxyGUw3JH8e6vsUJaMx8SYGWVnrrFCtxaDSnXcWoGpoEVSgfkU+xvKb
xAPMRhqg3zo/qS0UAjWHtVYdFa7P3wpnEOqKOKu4/SoNwEkK/wmBVF2rSSB+gUYl
6KgTpKUISdvEgvUeuzYNagwBQQ7cwW3Njbzgw9Urubn4LvPvjfnVRBFsIIrVv8/K
qy3EuyjvOhwQvB3kT/EmeIo14Aqop2NWDG27iBILE57w66O51KPQhLhBuht+NsYC
sUZAfEME8mSApWLfVrI1SnLxARLWoDl0S0r27PF2sFaIfq6mJeR8TKSUgLTOkJib
ljHl7mf4ZuDg7vyd8/0fLZB4VPNELyrUxCoiTqxAvMRviJ7WRaB/kRW2XDyqb9b1
/q0Wu2o+40mUQbh7HMXBEbzzDmhtwP461kx93NWVmP8Pq9F2powiYqmBS5sfBIZO
7ewVcFUUV38zcS3weQqT7PJQ0OpPm5L1av6ncoGELZd8KA0XF6EePTd2ZxdCo5/h
J2jK8QlaCqVnG7OBil6IAp+alLifT2cy/j+xl1z/WnaN6d1c2EQIOjWQ6s2Xh47n
lpBwzzeA/y6WMVaP6O1dXg7K/Kbnf9J5Ic3e04h0i7d6e886XlqQGpXkFblTL+1a
cCGrzPsCkPZN4sv9xTxkH/EvvEXEQS56hhBgu0grEIVaDhGXjZV7++Vgvag72gae
QdybpsPmk1k/29jrdKcDK8uRkII29mqJS+59VjddikN/UPESMdZ6lwNKawQqCTnp
JsrtAtUWQThkOPQNmPGBXBThb7EAxbPJT6O7LdH31R2xgb9/aUdHlns818uk6ZMf
/HIE6eINRhJLKzBfPJUv1RMpwqgBZN6f/miuy6swZLbfoWZyGb0nEGoPcC9VLjf+
C1lB6KuHI//iz2AHLJWU0i+w0I9D1To4GtrHdtLPsnacmfA1Sqi1B8lqr+IioKxq
crsP3TBChYY11ynYBes2UUkTHVtlmoODt0JRJWvnTAx5J/nhd/k5kZhl2hxmz6hL
6G+pDlzMMLw6NybjSd6t1yEl/wYKGSejNHzWDdbHmTq+/oITN0vW7ehE+xpjoc4q
L+8sxZtI3NI/oZk9r/C5LJH9kQATN5vPXR/2E4PZ2B36q5d/e9ArI/XKuiPwr015
yLcwf+uNPiuPKPPXE4eK4E5l47UsNROSXd/nlEPRWjoJbRy9wh3WNF/9XLFE+qFj
ZurVssqNpChPtv06O4A6+rS4KqhgzBpWlXO0wQzNseUBOF8SbAuh7DOEPYuX617k
Cjol2OB5VRQpwK9A7YRDMbDQfYv5BMJNFtIFPfFGGrkC4JKtr2JiY+0//ooeRIlt
v3ceq8PRpDWIe5FZ1FQ46r1CeZ7UQ6MODCx7E+PAKYZuoY9GvWDLFZB++7osyPSl
2y74rAF7DJXQVCfl2lmXrlDD0wlri78knZibYQcb8U0xzohJSUpnPMgIE+JCFhyO
hmkvpmQ24he7+MEg+wm7mu9ZnnaHxJnVMl4LmY1EOyGFgh983I+wEcPNoRarHx99
q4dTZdBqdXsGnh0uxO6zWaRWISUPe/1B+KBnLn2kObNnQFNGcMFZczc2viJyCpUn
dQG8G1KchNlhZ2krqUrCL5zeOuhzwiWQjfsh2kczx9q5satsnmtRiAj6WNKisGCi
TfDkL/R+lcccSERIt5baDae+pP5kj7Zhm0oTg1Z9MG0DcDRQVvGz+ukbY2EfBzSp
nY7NQMZnZ9TnfiZCfoW5Qdqvki8bjdfC918QNncUHUY4T7Uwry9vDT43yQivVbYd
IZYoa2ne/v32T0t7IPn/ehLJBKQ5reabxxDGX9plIPTfyyzy5bkjV9bEPPonmCoq
NM9UqJ3nAFkaBhAJak+2X+cmowA8GHOmicnd4fQBJ63ZdsUunmMJuQFRdscx1kOZ
FlS+ihTR/g+5xKtdQROze2QpStXukWoSZG16WtitLWeM0mZuu++FwZtcQE5NFOjC
4PV2fHSkGjVpwpSRx4vAek+YscoTYrHfiwtTFpPVIPYPFhjdkB7SbOP/6C30h6mP
u5SzHOQNikPO9ZLA/Xoc7OXLM1w/CkfDpzitb0SAjgCwPjMiX4y14dtGLWbHxCpd
huBklfYOLCwBgTBPaX3OdWHoK/1oQWOqK9xr1pxn4TvT4UjGIpMDfsY/g/V0MV5d
+DJFUOPhdSkvYaePOqnW/nPysHBdYTMSCPap99O2cZtiZHYXXq0DlGWGpDIOFRHB
J7iuXb76g4eAmWo/r5WLigrB4i+UA1ihle+8xLpi6UHkBoZ91lVPYz6+mAE6xguy
pS90bYTt2R3w2dekMTcaU9WBZmP5X9xvgJFbap2GgQVANu+XzCOLZafbFS5MdEX3
wWK6Vvm3XRb7PH7AcUwuhSzztFtWlFRr7iJZWpkFrymdYDD+YD7/fgtYlJeMX5U+
m8PlCBMqvbcmvh8NrcX6xAr6Py0eKxSBoFQZFp8O5HR5/4r+cWmEbujIkNsC7/aF
tQ6+wY8E3abbOo3L6jk3Xhvui+4hRt35FKz0/bx3gFUgnjGDAw3t88yWPrIECgCu
sBV9W6kiVUrhIM3v2WYh5Qjpq9vhh2Gr6oz4yO7bVSez03DhEJh0xM/fcwbe3dIp
izMYN7XCry+3sqczAaSS9DyJmf5Ve5QsQr7JZijOjFaKfkeuQMPQISgdp/6rudOI
oEJkh+QmXTXb0dPpjB+2PqCe/++nIfdw9glF06RIXWmxRWYDfIzekOhZsukcw9vt
SoX4pF0QEnFFnEShN49OMaE3C6QBdbHu8Dkc7158BpHZ+zyDMM8HzWfQJqD1Hafc
HJXnqGQ33Dr+9metdH7ez4cFNsULfzTXEdmf2vDw7cIcwq4wMMKY/zfq0nOm1E8p
OhmWtI4JEFwRz861k6O265ju5fAi6OD6PyWRHkYdMDiljKyWe06t5Xbg1Q5qehu9
p0mM+Z+k8NSpbOiI9Sjte6BSxW64QV3I5Cp8GSWOH5z4pcLHEgpTwbk3K55G9Zre
05LTmP8xr6rdk22z4bZhS07J6es5nzDtAvR9kPIWOocJReDu9VjkfRhuz//sHuD9
uqVpDDgnrKdmXyL7rfneXnNE2DXafMnTl6HP8BF2+MngOqD5Om2TdZuW1+rnoJHo
ACaLBtULFi4qZejxsaMh56p6sQS97ntJldIocbYeHsPsL3G44EpL8fGvEM1JBMSk
nYNJiMBK4Wk63vrcS6wchNENohKEDsVeGmebQgsuAK9nZMrH1yTfx1GC1J3e26kW
IbBim8afe2p01zStkNHO7WMFCkddWCJV9vgjR0yY2SPb7HIz/0fgi+6omgBt3HHr
8Vek0Ngdl0Fxx14iX4zDWpLmK15wV1VTKDv4LEDleBrHWGtzLJWwwIEsLzG4wuDj
PqBAIv6OZ06Ta8/98BABy/pmEAzSehIPg2FE0sIeJsTYE37tfxUUZs41nHu/M5GG
nj+uc9Tn3gPKfO6MRDzYI6J5X7M/5jqlKcEwVnzFz/pJyTMbNdSM9kO3vk8WKf91
YNyRVuQDmeZy+n/ndykyUuWrubKZPi09gpWi3VqyHK6sSy6FYRwp7dbKuuIuSK7u
6VB2M05vifCKGONgQ6kOzXrizAdLtpLJXMhNGcqtpdXPM6F7e8ROfJuACDAj/qNE
QvIKspMhDisLQHt2c7mL05yguRv/uC/piKjaR/dwr2nX5X1T1GBuqTQk08wqIdqy
oYpfxZVaVhOoYwvksP+OWOJqa41B7yYAaBr9jw/6Iw9VWThiuVMU7gbzpa4wQgcQ
nG1z4L5NZcK0zysZH2xqb1cCK4E8dkkMGRnv3iIJx3Rtr8e/rEB6QyZrq4XrD0rf
j7CTdCcgJE0TzTR0R6lRbrJLvZIVqnIcSg5McpQD6PSgIEmevzP3qHrmhhhlo2M4
ZIJZDIBDUQtfCkY5VGzDeAcXtGHZ/OGjzeLibljRCyy7tgWv3IHgvV4JETn2OYbJ
JxsbhHJ+RbgXuRG8rlPe1SmysHM7GKhjAleK+NHx8DHakhgDRG/910vm+CzcrJmU
TdKA7o3i62+rVlhx64FOgdY7Wa2yed1otY+bxcThhErRQ8zxtw+8EW9jg92Z5PCY
m+rw+Hkjsk8khE+XZtAGNit3XOcNElG5lnp2b4fBSWK4slPm23z7vc3G9kPIJ9fF
RofPqcNZ6BWNQgSk/MQ3FtUI7zD4xJ/hBhjpJVyW+9djIebGd5pum8sDpeKZBsWe
azOlskE+Yhj9wgw+D8fFrNuIX6vEIgNHR3hNo7chCMGoZZTJ/PpCa91MLPyXKIIg
KCHcNeKsZ10aFtUq3xbufv3Hr6yx2GrJ7KOFdLJA3TFpBrn2cezHmKkpiQPNBAP4
vd8ZkppzrV+udFRO49ngYosaG0aT018aRMsOKX+bDkMggiyDk4eECBOKQ40Cn1OH
lF2yaxxRS7tOs3oFLQ786Y3Ee6T9rE6q7OmqieffQEw44F4MPHnX2/stSP+FYHWT
3OlHBMrqf1I+1cUtcM6UjEf/0w+qnyua3dtpSipScxEvyQVZvNVA5eFbz4dA9vl/
9XchDgQwCd4MFT+swoFfdkg+oBndY+tdrkX7ys7sYbrwtGwPhhMyI1NoMRlsdyFx
rlGUkv2TASDJ/SYacAzRNrY8Xg30d7ry6NarkHmRe6XbWDVqv7Hs/ejU9FXZB4jg
1LYzpMmpprdrd1deeGn5+k1g6cghWdGNXalAubB3ebqlSszH0sphlbrTrpLwZTZo
odi8296N1b8DvUvLHITz2Cp9Qa+krSrShfDUMWdMocwk5tGqTtKz1OaCsevjzAj1
wtd5jjf2XNr1LT7/UONJqJtvh+NoxnP0YDGWYxvabmEEhAyZBLuPX9GAylI8erbI
5ZTgQz2Ji2pGEyFXk1P28/kbJjcZXMJo8y/3aLF8Mq6EgtfEYqB0OvndaRTki1d0
M9TO2iiNrczik2/l7mfUOHw2myf2tKkVzGIi3wQPI9TRPXnqgYqtx6PknKnWJkUf
FR0+pzUFk33o67BJSoZlWb1uXARxQ32s/zIeO2XkA0k+xK5QCATg8scBGG3xtv4J
IOXrFtUQIUtas1q8cLr7csRC+eEQQeJ7gGI2JjBsd89GkMNKb7wtHUOk0exbgXXC
N1bnJ4vXn64p67AhxGaN9plFmZFLfR64U8btfHo2hoz4SnwSYF+is+EeZNOuZyPh
vk0Lpc5MRdGGj5s3qzTq4zZ+oDDVbXkRm6UzF1t0JTIUFGzjkpztuW0G0p+upKk6
v3BPDpvGY9Ut/3LDwOkjL+KDQlgEerYz2d183Lkg8aIQ5MwMUgULs3Wv0bVGP7lh
nFNoLPap78Slnwx7nLtE+lpxr2Jnd6a6nEO/L0o21NuLcfudzal6NbElcu+wjr7Q
VLJxcB0exiIdFP2M/wlHa+Huz3JwG3HmNLeyvSO9RJf3yY8pvtU8VqxLGUydAgLQ
H6zPE/F7kehDfEvJgEc6o7cKQvkBLRTbXpwfXRzqYiM6p5gvkTMaLlULzbOZJtci
NBcTQ0/rHRzVjdyAy79GNFHgpjrkp3oyNLkYkquuuAg6U3BKg5ghZwsCQ7cfYP7q
sJ3hgs+R4MHZjuYDP1Wi8ILeu3D42A2YNN4oPjEvG/AjXct7gSnsY4Ey9i8PX1Fu
TSmcY7wYhVFxpHLT73JP1KoQWsIQqhU2qeEwqRQ7nnxplQh0wOelLHWGJG5tuK19
I636gaiJMm17SqGmx7FJ4mg91ReM8VRUJ2c0p3t6E/rPQl7rhGszY/UyXnjA5D+/
ZcVIHZmyOl6+v+0iF3jivX5nya3mVrJqze3Fx4eAcWscjA5UKAgKK25XnYT57m6j
ih7Ec36h3cHv5WXC/RJhtFGsJ4yvkwcpsYXf7T25u6wgzP2pceqCssavWg77phFh
CD2gYa1efcmmMYu7pidYSllyfOEthL5vmTBeJPcH/CwGoqXEbx0YdX6m1sfOA87r
ys47C6ioYJHTi61Qg8/JSj/8blJvQNSxHfrWQ+HTUaFKXn9MvK9q5hxreaKj7XhN
zYjDAIOt+SDxtbpW7kiMCzYubVgmUuWvQsoOsqFndOLy4aws/wvvI7BUB+VzUc3U
voOfdVDDyQhJBOrnWR77fhAMo2PZlszaPaTV6N+vEApiGn3t99BxFpBGmKFmKs/q
IEqMWdRrheuphfOxDS5aNZE9jV8+9D5hK6x/Y7LXgv5PDJQDpiNW7Y7PPOVLs+/i
fL6QXDPJpPbmgGi/aYSWgczh/T/0NsAYP3CfYnYEu4L9PjjM19JGqvvc52DqwS26
Afjb+CH+f0/K+2NA2cwQF1WsVE44g4WVAhvxRkIff2j1XaIXzD9+LpVqx20TvIcQ
LCmsX+UOCwYXNd48nJGVo8oZojZbW0vrRKRkuYUNLYq2X1jjq2hJX7uYntCKdzUj
v71PhT/Em0Hpuuf2uUZkY9HQ2Dm+BbNJB54c6VhE+cwSoh5bhoozD3wvDoq7Cpwr
T4wrCBf8+QegVQTcVdlSH3pZg3EPBCapnoPrkbJAkbq8/K0TWVI2/awhMayqhdsk
G/Z7S00qGo0DLqPoUBZew86JaEjaSz+X+VJ4vNUT66FK5jt8E/ULaWj9jw0jGLs6
NfZot9P26+VOrVDIdSWd+x+g2s0VBG4And5gXNFgws1eTYL7WfG4odQ/0PRLjpfy
EnCtug7xONnFnx1jgw0vy7eIApGcZCoreNDJCJY5hnBP7yoWiw8sTxhqLxpT6/CK
z2mm9YENNN1b2CKeNdELGgW7ViAj/xy6zdJYZrVCVYMbJG6vDxwqkgA9xGy0lZOT
3rX8TRjYEHC0eR1NYzoVG46Eywxxnt0wyD6A3BeD+Bdtn0yajzybkOuNo6p3NJPU
hu1zwZa3duXg0x+3zezIkRW16UJH5/B8dTE/bgZGOskWgaxJ+sGmHZp3nGY1/6fm
jiDgYCdMhdN6y9wipkHficBY510kF9buF2TBlt+lF/3UXoAKqJMY/Ki+KgpoXEAL
kOheldt8ee6egrUsImwSjmiuRRvx5A0hoaKbX3FibNLD+VjT7KkU+4QTsuH3pDRt
XcK2Ln9jj7nMF7VaGugd9vwyM5Bpnn/iF8tmJ2UihAzFUtcDrCrahNu7Tppl35sb
rquZCtYunsxL/PTaaZMaTaYdKA9hGgOmk12915g4mYE5hDQy5vFnki4qNGDeX7Hn
H+WfYNEhLGE9CWDCfxkhqEREJVteO10xMayRsjhn4D9VZzfRO8KAequpN9pFxRor
YrVn78YtiTtwwt33WoooXR20Su8fBG4CChnmjwkkHR3ougB162QA9G2QahPhFKI8
0JzGLnIIoLiW0QApMX2NlqZ/qfSD32MxY8WmhwRvB8L8VoUba85zoRT/sPIVD5PT
svtrlVTB+Q8qcWXVfpZSJz6eNSE905ONoHnks9RhqlnHSm17yDK4wdkFP++rX1kM
7egBX9JeKAEHy2xSkY+QGhMsZm6+YqRwpu1T28tTv0GFjdqMZTiIzJicVykPVkKY
j2eemGK73685ojR2jCmZ5z37lltcRi76WmUnPBjzLgjNFiebFGv/kE1QDA+39Q1K
+bQQmIO8RvL/f/fTsGl7JOH+Pc9l11mAirqJDl8W1eErLpZEDG6ploxd8srFwKbl
8i1S4aIJRjIteM1nLOOViA+xgLQ95ypdIFIg+AFqCwwVfuoNUW3zN20FQVz5UTVi
KWVjocfnRTSNWIpySUyfndz1QwiwN7fYgrmyUXvQLURjD6S1q8J2Ykwp0C6ystpT
mht/JbVPZS5Me8bUHBsHql5UjdA1KaB41aBXO1ohQB9+YxIRHiiPsAOcYFrL2gHf
bi+Koreg09elXwiwD2TnNRXmziFOn3RFhVbVMG7lx301P9Vea7f1E2BaTa+L5ZU4
8DbDnowlUjAj7j12o2k5j+BBdQQVHNhTs3p8w76CiEK+vZA/uRY1/fWFDrMZ8TpT
P5JJ+vHfZbN4TBXiaRJPRgsT4WbiE8ojApPYX5rt5wp9uIJvXDLUqxVDhZylILv+
+MBkmgCo4/karuoc3Mj47Mvekz9Z1MCefl2hN0lImfeNr2ftAZzdIAYa8hPBVpNc
/ONWJenXgQO/fJugkai9R41e0oDpWeB37RT/eQ4LSrXVAsUSd48nafAWqzAPH9RI
mOhH0WFr2ep9q+Yq6nhR9iB5Lhqi6hYYpPVoESMQFILqwpaYiwt8+cRV9GQ/gBCV
s1u7rxdSyIIoOJ3dLC9d1xefKeQ4fyd4MOEPtFpGPHDozZwYTY7FayuIBXQbh4LW
6QjkcUkfGC9CgiTCvZBz2k/zTL6AeAnFhg4ztTUy/tdKmuwqOekXsYY1DAPGGNtg
jMaRX/IWu21jFGVB1mguT7I99qi1pAp7UEwUouRJbNslR94uh2bS+ax9Z7Zwl0QQ
e2arkyjdkRLq5eVXUZHf6PdiMfzuCaZdzPjpsI/IRW3sTArnIN1BoK0K9ivGvBfx
TxaUUpa7wnL8E7I1o1woF29jGma4BELG7G3GBWCrqIVZdfWgytgzddyS/u6Wl3qo
tHIBpr3Dcmlv6CExXtxolLD5vcINNo2vB3MErPDQqmZgyglr25faxccVa2H7p6vR
kXTGE+DmJhxvzMWG3WhP0/rVjFGmPABK2z1F/DhYcHR1fHyrf3cf3+frbinn+JUI
5lbpMrhxvsFT0hjCNst2SNATdb8iCos+Lbmh94QkTMEDjiyGcUrng2jbMKb6uUps
GpQevNG+Eijqe6PabevyIibCdq6tArwpG/FEQKX2JFJQVC93lSWaCU98Lzl5/jLM
mDzevL54txXBEyY3qPztAdOigPAXVQ+5cft9mpFGVYZ1OeDweuD68iEw3UWYOoNo
pkWOBNFErQu5yn0tDffT1dQrLD13JHlwfkoE+NzKyCNwwGXtbwolUSvxdyEcgMu7
JeO51fO3+oOwDbOQ0oW34cf1bOi9JijPR3gguybYmX/f++3/rtylvPAeMxyjl3G7
MDC5t6VPyGXxiIgt1OwXyxrJuV2TrJZe9TERcw+4U+fdf8OAkAu5GcilBo9RuFdV
duZMmC/NG1onOeeo0AZefFxecKXKGGB2mjjvtR2S9QUcfuwv6/B203vVnaa/wzer
c7RILYT8BVBX28qv0ZM5JDiKdyufyXSJjv/G2fFEEzjljXVDuaH3XM4m05GjPnBE
0YN+OHOK2J/zY6P9wX2N2zmF+agKmRVBFqR08rkprIUN7ZKjXLYjSp2wT8d6hulx
JzMszQRp9TuIJg7BLn73aEmK98GaHiqhRNyRgswI6xOOukASeLr6KA6+g92ihF5Q
YyZRCPZNGYQlnjwoXLyR0p/g0fpzZRwWnTm2Z00cNz7VkfqM+358oogekaF4oZze
eyni5jZtsx7v9c4qBps2VBy877k8h5wZFHFvuCi3y7k3WfUwqYGwSZpmQKH72Ied
1YUUXPCDDV4+tBVn4WEeUB7dtABTwjvnxLzCacgFoFLhlmW9/dpEKX1yDn/HfiQA
spDwqB92pqEOGNvvFCv7GWQxdMgPpcZ/e6EAkTzjEfZMxcgXXFqwaIuOA8BVNTNr
X5UiFjObvkIiApzpyrRNbgnh8fmG427z67SQO1Ul9Y64Lgk19mMi9VSmkTYFXrqT
0NGXBxjUWLwMCjpEKBKKSG1KzR9q7I+YZ4a7g4SAs3lIu/HxZDZD+3eMZKz44oMS
r8/Q5KK59UOeYYwqiJUlpfPKW1Y1e0cTTVWh+s6L6jrHFY/Pxt7UXjOJ93X8GKHm
7tYYnoSofQlC4JvlAX1eGR6USOV7VX6NzPySbD972S/zXPZhwGvS6ki2OD5Ugqle
gweD7N4W6h4ue4L1ucr1dowRvDLC6BQhIr3XdAm4JBSIuvoFtkg6NyEwe6gOf4s0
zMhIQfP9Cqw9mnNm8wdDpN41MBZmCyjLtibN3SoR8ALYOsAVf+1ru8fG0wzN5nUD
cmDDV4FmxCsiCobw48AWsW9BLOiVjWyOdhTeGL6SHsndRWTImtkti4KBpjqNOwyT
Xxc9S+POrg+toMwrlZm3EzlwtsCXUAZ3Y/ALzMzZW+nWCZr3VIu5BaQ6XRnXdaQr
RX2G9XJIWHqfTEslGC7yGyEp/popgOZhHhaliJxIA+KRX04sj7jJSkE4gZQLCl+b
Ol0ukQtcWHv9EY8Cbsc8C/8WlsXJmG3fXcT5m9L8yP+7cyUU14tPwLiBH3jJ5PWo
Qn5rz81Wwy3pQL5tptAKCi/cnjeeiyZltLsmzhX5p9wyif9sqKoT9AFRvLlMvklG
AABuDYbyt7NkkLlfIbDYcKyhH3iwN/YLiWVWbFd9uuHYZXJ0M9lbgBMcZVlWQrvD
JK281mlzaXA2QfYj+DK2lMjks40H9Zv4Tk0yUxHzGqIo19z37t1LPrJB+zR5Nmrp
L6XhoIqOeVyyoErZSqBGF0C45hdGerFHwv4VxfaKRoGEJ+N+4QpveX9ZySe7ccmj
kWHvDijIW1y5RtDHtBGg2WJtAcvutFjsge6Um31r0p4fGcc5sDyPnW4/7QH8JGOD
agwOlYhRxpkWJjVCtPpthVu9NqYWCwUWSRcJ+Qb5Dndmpx54VS9mFklXIoPC2lst
emIM7pD0Q+aRkdNEMVoF5xz85Lva9EuYmiL3DPdpRoX07qXyZPYrikSu8hU9qd+t
6j/GGDLUYRh1cWR+kjJYDOSR9djQEl7WK3PjwQKLsOVBX/hIzd9npUfGFl0+y13o
BGB0MvLEXmnpXRhmdt56IvyJRtbo+1byP3UUteWA1D/jzjyi520z8sBQM7laa9Yc
9grKZyLx770ov4zfNxSI7pzL0IJlQ5ywacwumYd1Y7nKEVXQoR5oMYP+k6GTItbe
IjkfgDTn+XNfAVU/wJiwYx7I/KHeBV7p7hwu6lTREisrFNrS4L9V3u8mTB5fE0EB
n+1YvedYJpkhburTM8FlQA6MrSGmMO3sur+JvufXSUMY6+SsXGAPw6AMnbyWy2FW
EwkuVE0702imayJhqviM4s+ld4iWFhF6T0/3TXadxU3d1d6a8F2/Qs84BDFtE01D
LWrN0+l+cje6ocD4I3bajyseph7EzqRg5VTlR07CV05VpYQL4knUt3D+jRdVk95C
reA8hPDTIi0F9+rZROoI2i9SbaWKRLX3D0k5xoBgvyzF9sDMlxrEKq87d0Tn5BmL
uzPPRdTy5HuAk775aB7DT8EJGxH30AYbo6HOpznghvsuBN4Ra5OtuPfP8VtFIzte
7D+1abDYv/b5wnukmeNsl3+a5hPeXzUw6EaR8/4GmssypnJTjEcotiU8+yj/dyAp
HCqmue5K0mmLctsCZnU8f0CPPAOiu7rYl8ZCHIPwqNR0EOMx8uhJ/yfwQbcrzlTc
vvEn857BxcPNkwe3b0jnRVxQK4zdUfCXIY9S1CU26NbVYeod8NlkrQGCG3ni5gmU
oMabWVAROqZXQSFojagnNTQ0d4jC0vUx3s6LS5EYqPrvx3t6SRIUCCJC8keMbuyP
5M9YuuAMSNHTB4EqQbN/zbhOS09uoO8cc0BIMeZrUX/Q7rvkv6+1Pig2tYhiOOWV
7aPdBOK8aLRK9BFzjOL9MhxpQcxPFreL69vXN2L4GxBcKhSFLAoIOMuob5zig7OU
8QPDCG4kZxcdLEVzF20gbBIG8JwiSGyCK3a/MMot0o/YDRgBg3z08hTO3wMAh3cX
2S2ZYnrfchDcI4RLqWLewrCgTDOg3BwgbA0ZyZJm2QGzysZT3FQ7V3lpyEC8jiKO
Hj3YnbueG3rXH19Rriag8XYGTfT3Q99qeiERMi7uOA7f/hXSak0cpZrgsEZnKNuU
YlL50wqi5IHAqxxkiVLr5QRCGHO6mJLOO0U2Nn+8Kty/C38KiFQ64j9eC3xF36OX
M2fcZdMUs0NhP4M8o/SSTw33xA6/FXnRU7OqWx4Xl1iVRyAd8vFIJ0I6/qgfY9ze
GILnrSfJW4MLd99cPwiLsLvxcDjdwjtvIg8mxj8Fiz3ugVwooMF9i+f256Ct/nqK
kvTuBPPFQpTHawrfkkG6a4ApTzfOxfJ24rpIYEQ/5+9SxKWZM8j8d9fvxbKqZ036
+gpul8cFBLGkGLco0rBrlqONEPfT8XN+TxqVz1jA6h3py5TyC0E1W5L+92xK3UmK
ZwjbO0ZRf6VsZN28ETiZOyqZuE8UJFiAfrDlA3QznjWyVhxqOpNo3JKKjqzeCYA+
Re90effiVogotY8y7i1RtHn+EG4N1f+fjyDP/U51AfUK2AW3MHUtMtslUgzRnlD+
oJFfePpiNmgBko8CBsm2pqlPzxQBe0WoffyCiZF5Gp08puA6HE+VvMx1GVEEhTKr
qqQPTo1EUWmeb/roX8dHMGE9pGT5LHAMaW44sTp4hx7TKHdA2DzOeqWDxODZFRwL
YKZGRlwyRfuS5F6s48VlACrWYfloQLUqRo1cgFxtM4eGCisjphuSELDsKBPrmbUe
Seyk6+Qehhuk+7XxsGqi7dbsXbPO9LmuSzJ0nXXXTsEXbIWNy/kBhrrUSoNqzIMu
9SZcJA4mdEsiiS0eNf7eoKCYfOum1OX2ZIsDnaM4joGcCG3/2d6K6l4yBIwRcsTK
II3sNQanW4HDU53KnnE/GTBPmfTO+Rzjaomw0ZrDz/1ydQFHA1FbEtCVhJ/Icqrv
r1DxqzizR6LJKIQe51Kq/G1pNHbkHimcWuFEAyLcN8RXHdvtdu+ZgD4ii7iBSJfF
oE/lDXWaFa1epcHZiXGY9yZ6Drk+mPypVIgI0AwkULoOzqdX1l6+Fg3f60RpWjG5
jXx/poxxaJeqh/dbaaRfZzDwqPPRINc4rNyXBHFSGP6/62DF1Siy7DdWGui1YmDx
eTd210pQLM12jQxQhvZiZRU3Z1sMCwbOOdAAw28S0xlcv6Zihk+O199knYEKF/Tz
/HsT3s7zN3c3omdW9VBOn9p4oniI5TQD/8Ln0GxlqI6F3hVAmcmuv2TbrBBGPhHI
+EuLKR7bfJccyEKqQOznnN05jbEx3WjwvH9lW8nWcV6dHm3gQGTH8Lp1L5JNbdFO
mvUHiMN0fD/6wgaFKKnTUC21XQfaXphVghDGuvGQyBnm1Xn8E7uLnKa/7v7yZw+l
HKdk4q0OukWvfUL8vkR09HtpNOZBqqYY7JtT3XA2L7wwpxjOGVXl/DGzNHYxfNNy
asmhpQR9RBcC+iiL8plLnAVZwa76jYYRHDxleafcRN6GWqnI5nNivpPXyYmt6BU2
33xM4Sc+dspp3XQ8RqHsJusv3jt1i4CwwAzJDnArjc5e7wj/TwRJ8ZhsYbTB/KaO
OU5aTRDOjacFGUQ11fk/cMHw2VioppcYdfLuLtwopnnol8wZ312j+sGlUccjvzMO
ni9lnAgGh9J8Fti/U87uagYj0bGQF/Xm5omGNA0umfZPZ9jfm5HtozDXXj4CM4Uw
BcyuXltXIC7oqX2gvGrQB3/AhM6G9IYYHojiC+WPS1LBMSLhjuEDBzPX2q4lO7Il
2uU7cJf6DOHkyrHQbpDAu4e2G/+y2fGeG8YkYDGkWJASar3oFsB4bGhbAWCMXikG
WpXFNqR2jm2m1b3Bp8Eiod7cwBkf8Msf6TG/MbM6DzStFLYoBH0US4iUi/Aq5Fcv
QfYqDyIdRWAlHErJ5LCgLI0GMbTwBah4PJ3FTGrZxJ1a1s+X67vOx4J74T5OcAK1
Rg+RoTMdgD5Fx2Djwja/FChaHK87QeY3r4FAotuOeCrTB4hZHDMaOXHqKkeHluQy
Lk4FtuGhLL0tBInvKvL5Q1h4aaGGvl3PfE8VG5NvCSZ0px54Jn83Thcdmu+ltQAx
8sLiIUuLWWHOtDiBXdFitbPpJtXNgorbbpx8S5rAAkHgNeOKQm/5zI38hBOBfYO6
VH9mr7nEmUo+JbVeXnjl0DS+5k4ifqHv9yhbvFfEqgkr/CWErbZAhcqWFSPMZbPw
gA4KgIrERO0nActgrnds8ixuGEr8uoCzH8NtqQP9l7Ex+at1zr3FCaTbW+TlIJ+7
4RCBw5JsmNzJfyshnfcsHobZFy7fSFLMTHKV+Q9gcCzvLO2uiVxNlgS1DsIJJcXi
LIITtmftBWqTREDYrFaWOb7p2qfasORMSwbUOESOweki3NECArRCukDTgjXIfxNv
VqTdNwi5nRoyQTQtSgdMXFseGxby4yY5lKDzZdvbBUhzzGPdQEs+5kFfnszq8nAf
UijUYCD+ETVnKc9+CicHl8fgKPnL2nR02ShTHKWiI2tdBDYX7RWH7Hdu88B01P7Z
ogdvDFNbJNsiV4ZCxVvNVijiDV2uzXfIiGxAZ9cziRuaY0wucSk8va20xaRdSIaN
83NgL70m/MGe0ANx5mWIAh2TIC1F8V1TMJbk0aAlUYl2HFuAzLIV+X3dPFZ54bKs
Zig/+M5zXEp8rTUs4adRxW+1gEepth5ExphvuDgTNYqZgCGnVn2hjE4Px8+JJnVR
LZNQK5pOg1YSQVG4vyGBnzY6DuWcVZyDP5yoStKGAPzl50b/ed02HQ59paUkVyVQ
sUUerHdspP5zrNoAg0Blaa8WbB23AzdhyffdZRSGgfd7p5MJo1Ti6SwSNb1wOVNV
P1ntyTqBUEFqQPgCLbAaqDWd9XgUJzrZjHXX7XDE8dnVkHlEzIV1oDmLBXrVK4Eo
6Cl2QAF/rNu0twzkTJdPfEwkSJ17Zhrn8gJ93NqSFntmlUFLtPR52p2BSQp/dwVj
Tc12mnHSlCZlZhIqNtjHIphHzbqiGRylvVGJWdG/AzzAJBHwo8SPBFucN0SHZnYn
uSwEI3NlA2mLaFxsmqF2PDWkP2KtWDUehcM9R6cMY4Iyk0DICYGUgdX2eP1V+CIf
uPpq4a0/9TvaVA/3njeqpsAyZWiK9Dmj1km5UJh95o1QysSZfEqamXblJj8Hy/iN
lyqOs0PfMOQUF5Ku87ckK7nJqHo1Fw8SdWQ94IMm9Ssz+E2IBB4uuskqFvYE9jmz
AZVWKnee1WU5XalzYwdHbrWqTJuK+3N+/ZkOp++Waywyxyw6DaVVDz2k2VIZeumX
vP8gymwOfaAbCvOnRRa42NmqAejrAxe2D8c+Ovuohafg441LwdC5T4s6PVXuGaiL
ylL6JEMPn5rRxZ8t6xLKwBx7olqam7X+x3lOQrZrB+j+PSDI87rWuN6U9eOf6MQD
soEF4JNdj2XVcmhEsPCDO3s3IIuhSmBCJSpE2v9GhDfivHkx4FGkURfbXwrPDaPf
uucc/Xfkg2Y8rymxxd9+9ZQMS7ZzgTckTweKnTLpZrAIO5JZQy9zyuecOGHhz2Xm
MwtfAJWBJLZGdLHfl2HwRts/t8gyeB4xGlcjuxcdnW/joEfh8sfos7UujlfDVSzh
02IUK5JDn0q55ZE0qGAENooMDk0ux8Qa48RKx2/PLMqXykL9QmkHl/2LVsfKkysG
EynwbBIVLgsC9sN9jb6jQL4SC7BATPUPfCzxPTFpTORedRDxOCE5/h/i7oRtv+3f
ZA6iRllg/ETEyY11HQImmFTIx0YQ9L86B5lQWD/KW596lATlCK4hxXQOvEee0VVn
5qfZYFSRC2/+BxmUUd2LoseaUFYPs0NwLGb/whwUec+tdpDr5dRHOISIRQ8dqFSv
J9Ozjrgx27AsHvy2kTTEoC0wu9aVGxRhpg6NLfKsiJl4+XzpnDkoHrTFhFaV5CSZ
slUlJIAKulaHx9rKaUma5eL+a8HkHT4T6X5MTWKeMbdBb3dh0mpAWuYc0W0Lg3Z/
On2EeiFzPtenDH8kv/uFdQKhrbGpNo/BMHBCDX/PNQGrnvERT4Yd+MoPMonQfkWB
VEZeKYIKAjxJx70fNVvP+77/kz7gjKfvzEw7EbE9oV3JzHBfcUbDEqFkeYlxyyI4
Tq1srN+Eiv7mUlrlNl0FbyiekL3RMM5sDCwxjj/3C3IFVhacrBFb1tP3tFEGvkyO
Xg3cNFkppJxzABXca3x9xHCE2yjP2ITNihQpdqFqtz5+BDKGqJLC6WGxy3obaZUk
o53OkJ/8rM0PzfCwAprGDoowGhVO7tEzeToA+dIT/UgriQAdaEjzxXGmNGCev3Bm
x0G7xDMDDSd43Hl+L0XOpZQnMb2xAEN1Y5zjmSvr1t9gNlMQovVe9l2M+jLRMRZn
E4Aa4wFN5Bm/jz/jSLxqOUJRYX/NNTN3bjWoOlZJlSQdPyJAFmSOH3/DikPnDEDt
DlOwaWeBSae0JQOLTjCNPhZ8DIsc0s11zm//WNJWCS0CCPRwUrRrJ7hLksLJ1Ba8
FPyib9b/PcbOliVbxIDdK1IGk01EY0WQIKEN/h3qLwEyfbfXxNaFdgoDfTgaABPt
VO8znUpCWX7fvLiaHpTiSDavXVeEqoqluZnFoxtPRa4n5DdU+2yDUiuMOjHfgUbt
HDY9/yOy1gv+gDJAnYCLLvuM/IOvfjhda30EYdu4vJoSDCdt7w/iVBGiGOIQGDH5
+/7J3KE8/8x8T5dMr5LtrAticgc20lxIlPPfWMeiQn9/4ldt+D1qHb/cHB53OgRL
6MZd8BbTeAWYKobYicGXCjvPAV5AidVd9FzbtEuG57q/+LoQIDNvsnXwQEL8WgdM
tD71GF4RxmOlfHmpWu/ICWV51MxpET5taZzY3wyeIFCZWEJsjqIKjQZIUiuu4+KM
1B9Dqs7/gZ3Q1ZV5soEPKG86e7S7A+5AYA6z5yeJKKxKwZQ+cS/YQyRXB3/btMYb
Kw08m/M3mj8iy0L2oCa2yMNjd2jlxEPKxattB6+0gLRlsI8gpTknQ07ZXmZbrrz3
Wng+VG/RrHaXlBg1glzs2D4BkYSnTIu5K0+wRZ1LaWUNDxuvXR9s05kPqW5uPudk
mpjxPQcOvgRM1PC3oiIKNIVIh/1Nx2uZVrX+DF+mdn7rfp8jH77Jq3mT2OUKVddF
5+7UG2R9yV5hJPfpXxIGPaCwB7kaCNl9weilE7W8ueASbHPvG4XsNhNk8Q2Q+t5q
n3Rc+cFjhCICmmjmuI7ybfRFKZ/bvDbHt9Mi5W7rXgOK6evq3jkrUmaU+SQLlM+Q
pPwZ7gnp49Be/ksVPgaBWoXbh/ZBSrUQJ6vfFlONPb0Y2VOALdFy0XyMjmZ9M26j
bzraJhkwOYIfyQQZhkBtbPT3rO8Fp6lgLvjUZER8m9sbxJIndqcq3VeTdPDv5tqF
ZKypy9kHd4buI1pCCc9NOA15rG2c46m17a78kLqhpuqzv+Mb1x7ERReljANU3Ns3
yWzsGCduoQugsVPSWWUJ+wogYb/1g/7rxGukRlbmYWUJgaGpPi++I3O7MpQNFAVE
Jp46VNAtUwUH57JkYUtQzUJf3BtbuU1ww9m++qtespJWRR9Vb9zLDBqCMrKX2n0P
tC2hUiHgRKPctKnX8JAzdHRxlu+cCro7xFo4E22CWPh02Vs4JKPgaoyWcNr2WVD7
BNYC6/cwgCgSQECr3LqoBeKVE8Bq2w1fzXGPXyuIPI4mZuwHKqbDVQtmq2KGREMz
1rURDi+xDQAsstYvWeQYADDpXhYMaIR4SzQLoyaOWlPbLnlxpY15eDVCpxoRhTck
XbmXk1ZoRzlNEvJNJtaVObchpqZE115TeSidc+l2DE9siONBp/C0V8Emxo1S8CNT
Xbnm/qZNZWE26js59dBJljxV0O5K46mYdMJOjIfl8//1NmLaZXNWFKRiCfIcaaYy
Iqy7lHiOvrLsWtPEC1X5B4WDjIAfrlv8b+VGogOO1I1Jlr2bV2glicGlgrkGORPv
qbYZBlRLjBx1yAuanSrly/15xQAR32pl+2GB/WJilD+Q2YWayzKMfM3h98E/jApO
MI6LGxgGYiIiEwoJ8K23ZvGjIPR2Njrd86QDny/7nRwRQJAcmVAXmOB4oyjllPLX
UXhHMa7cBPrAkYAeRTnsUIu9up60cyWHOi6MhNPp4/el1gcvWSqbwzdnie+8sNmG
YeZmw7icI6fxMZe64+4oSvQstHWeAaE4PCYl9sBf8+Q6TUcQdOIe0/XZkfA2wGHI
gXynAwvJkyDGnyPB8TXYazjNvFrB5zkO8HL4SQFd+vnRegVZSxj+Uj++q2D7pkvq
7u9RUpe6djO77/+NJPs7sWbnyGs4JMwS2ZroEB/rqAr91mle/cG/X0+qOz6MkLU0
HJD4Y8MctPrsvJw/3or8vLdxnujqfh39y+gf2TRE+bVKbq5adXxOxxZoLpNvp8Gj
XcK3ceHCc9XRGELpPAZGgEMM1t1zTr6eaN3dRWSpBrSuO+zoWhWquzguwTId+GpQ
ABXV7Qqwz0etnRC/yQaTOwfxEAaw1nlGPW2XrEz1sR/wGPq7wW/iXyZZubbIAPu2
G/nMiJbkbZknzjpf8DGoGH2yiuiT4+ScDgW4ht1JNLxk7O7/LnRhWHlxHsESZwGq
DvN60mBCIjEPydP9EsBol+O38y77L5DMxlm1/9XXaX6CQ9+AcahQTzvr/Jep3uiQ
+Ykf3viFIKMFcvJXRkmJohdsRIlHI3vxJIxHwgxDn2XIlzDZcb7mJ8HpaZAaZ9vr
N6IIAqfL8YCUgERgAgZsQ+2Gx4FFCft9eFaUi2o4usGCBoB7M55fGgFl3qN780UT
uBVcCrWJHJIq2LQ+6fsuH25IVamazyRYg1+Fu9Mmdy9SVFLAG1G/bJTCwbksOp8a
SPZGEoxg4+rHzvWMMHc7DXZFtcqJ1G/uGCxGpsSuxq9Ub0lbKw8t8jBYSYOBhrzn
QZlCigtYYH2nTZ0nY5rmqWA8DOlRo/yvl5+DEAt8jZygCaXw5bwIuq9WmrfDZob1
9uoYbvkuLFVkM+wVxu+AEThvtPjA6KbieAOnPK4+ImzGB3JRk0ugPqmBj7zQA8wQ
skctkgcspmbC8foSP264o4238yBJRxW7q6R8omJcd7JzlPuw6GMEliTN9T8b7dmd
/h00DE766SzaNl5OkyELUOgh8PnZma36j8WC+GMNcX51+EENbCa1iBb/m5mOFCkn
gkVD8HIO+qVTJbRJYe1ZP01YBbBmm85zlJv+jV6YGIcdOP/pgvc7F5c1QrmR2EkS
iYYlcMbBouW9xBcfW5CfgJUf/B6tSxZjylJWI33CC8Mc0GReihRAsEOCHpDMET3A
Gmv5IJSd0xN6m/2RpKH5BLKzqNakYDN5zH/uYxGHNqOjZCJYEs0w8YTv1+kASMXn
MT0FqDQH8af8buvAkwyNwgUgUvIu9PIZdNn2VWh1MKVL3RM/aRKj6hwpJx+WTMvF
t00R94QQpKlVaQg/9dhOeNdhJxdtgST9i4gLkIEhwveoYgC64Hb+f8NgXqUOsJJE
LZMtQZInSvRJizx2d5sJPK8N8zojeLN65/fyjea9jMHoTTjnJ7WqcfxkUw39W4SC
jvpF6oN/VrVwy1opG/T7XQ2QXVmgJVg9d2oiGnX69XP38Q1GDp4rnU+ZJgu0/dyR
4ByGUljGEYaMdNSIkrVnMHWUnNtngC2TiQlui5Kc4/Vpp06wpOPFs7y1HNch4uiT
ogiVmN6J/kSYSuev0n2+0c/CZzbnp3gg8TQQDBpzbPrSQhaRh631ZVB60IVuupkp
581RLBagCCO2Xb++SCkSYs1d8c46UEdQSh4SM1b/A3vpZF0gioHc33XJhaqzGyH1
QCNBcJrla3TMAW35ZmIb4nhc8UA9AVcjUPcBpfN63gbZmk+ivRSuYkKAFadB/MPZ
ulEgqSBeTC4eCEBG2ruNG740rpJI1YJbl9R87yTAbQLV2jLueUl1PZEl7yLG8mN+
E3d6mEA4E/qEuMsh7fnTqAnMcs8kkpnSsYwkMWJVz9097b7MwH12nEEbU6qL401y
wihUyjiVqha+I6KKvA/uP6HcMaBFRci+xHxZ9papAgH0skkyS1lZAyHHEvREq5v3
TXEEDgdjfITJ5j2MZxVPU/x7XNYrw1MEx/4lCS7MOA/SnvtZ0inbmjpUaQoO/RwS
hYP/J0UEjvk6h4hal8N3uKeaY28QOIWPp5xvdMDp5nZxlN8FpoRR+KyKnf4kB7Ax
Ucc1Wm/fc+iKQ+07CFJTbxGk+/5WBdFEbDw8p6aTwTOPYOojoLNOsZsM9ijD8UR0
lZpzsfeLlgGW+wKkgPY5kAjMEyehrpdFMr5wCOI4LEFet1NHpaLpx7H9+gVtGlCS
QY40c0YTRM8CFkZp3qsAsosyaWFvOsdkVqC4lccxDz4z/kLGW2Jj9YX7QRQsPNE+
Bc/5GmcZeGFjtbIZQyVWFWxHuy0YJtvgoQsRb7UZXHY8LrZeeOU8sFZCrHvvH9tM
IAlw5O5Jy4OyBFdCJc+x8VjG010wvzOIjBSddJbis63WjVVvduI/sNMzXiBE3bnD
MNvjQo3ETbafw4EJOqQk+wcVeCAOkKoXJK5ht8zX23xn1pj70j9fgToPqPaPwynJ
K9LE/tJWqzT+u3ge5t994EQQlTKedgzmuHVmkdQXiwyufjJCt/SIxWB/Llo8/ETA
EiytfUaQmvvUAoO7YpXyacAMqvj6CVwhl2mM/B9D+5JZ8J6E3hNsdCi04FtdtsX5
rnYgVDAXZTU8fF0GQ17u4zSW/RxWI+eu1GUR6TOZe6dxdWaHBpb6JKsO/Y+mhn2C
sURbh67WI4FvCzY0QGqmFoZwfeGQgLGIYx5wz1npm3VxGNQeCOn8DmGUAbGgOocr
aj5rCeetUQd5iGLY0MTg9SuktNL/quwnOa/fULclwr5B2tcUkeQdjZ30AQTfEcgQ
JowacBsqbjpjaPS8CwUMAk9wKeXraXx45Xo0bPdqRqKKJrpRBVj/gP0LmLJw0/6g
iA8QrPSgEoSaFX63nTDES8i76zBs5qVzuooXSIuE9T9YtB3NbFHdnfnjLJxzTccU
Kh3b+mfu3mEhMjDLol/Z1/SIaI1VvoWDKTU5UnWkB17NmoqcBmf7sbGpUIfg2zEi
hP7yyzLsLxSGxmWJw1zPLLs76yUy31yDelI5AJ8gvOuUXV7jjqVEl+BP3iL24fR7
NLY5mpVFF5mc+kARUk4Nz7oPZjJv+njKZ9QJVMyCT6JrCesX5GDUxTo3fT7gbeX/
2Kyl/CpXdRERUfQopip3UWJ+jk5DdzTAzURIzsnrBl+SCP2af/X3seFkwtTRqMqO
nQWK7WHaZ87EkMVmFi9lSaXwkFUvaYyllEWSGC5BRnjJ7vJgUxwT+wU3lwwetxwv
+9c2M8Zwth2paIVDvl7tXcTsNbC4GcgIMQkKrR9fgFwqTGj+yP/AmS8WghMHzzrv
fjZjoscmtMh9DrZeANkAzOEcfvTDuv7B6OOs9fhPzpG/0kj9zTEiDIoR3+E6Je8V
GLu6uTNgayx5EeAHnFqQ10OfztE0UvO2k3nXxfRBy8C9vVwuJM6GpKkCHl4XX/hR
asqZj7BvbTHS8sDSg/0VzIRQCy5Vwz1RGO+TF4UWwJxJBGDVgXmny8HHqbyEZWay
0GqgvJI2r0pEqh/O1pTF6Wr0+xwddSgw7/EsOQIApK/DIunw7KXWh8sKavO0qCKa
D+iluKvosP07s3gz/gtVp8GVgSwM2xLVeL3XgGQyd4eXLrT5DbV+uIALH+60SwnE
bHueiHageSOCBlkjVUvdf570hjgisV940gdRalY8ODSd3I249PT/HKLMFjqHeyBb
UTv8TJtPZc7JmJa9jBSCvypMPJfjT3fSWI+4EVtWFRq97AuPG0v8FTncScSj2+Qf
5m61cSK4iFqx/fzkmjVX/sQIyy1GO1Ho3N7tBwnDHkd/agOjCb3ua7saF3kLSDb+
4RDSBmLZxgvMBfeyeG4vflQnQyvFzlJyQJ96W64DKnP+YvGkvpV32YOZmbihCWbw
Ez5wiQNBGcFZBW9zQQ++2Nqyt0OddXBJXEfGUdmHSbBL2Pr7Zu0UPKiS21ZIeDHh
Rc49WnUfA23e669DXCCHchOxWzKTFGpD+uboaPU2Q1uzdV6AcC36MZji8+zjx38J
RRQPyMf6JRqc9k/57j4VlLBehdwzB30nQzzqvjzjFVdCD1TqY74jQsGsFD5ELMlC
P7GDVaQoFenqeL748jOj1cPSghktSF9Fu9XzGP0fAp0ofPnUOpZcUW7vigcU7D8u
Pzdl3dNw17RClJUaVKLY9K9JDVgFP63ilH7Z0AWxsdlnoo2TBATyZ86GTI6JH9c5
tjkclpJ5E470Pfd1zz5mLNrkP5nMoPe4GfVjAhJITO5CeP09Ii4wiWO0f1lHUREp
jkpAoF2AZ0l4b+IHChFVxbHJO8cCFVzUWIJLUfLQm9T8Z35CJUr4REJ7oi+9QHxm
hDuIgvDr3bZTPaAvPTmrJO4dLsXWwUqwqVQIVy+SjLlY4vbMCuqkFcq4dpEkSANp
8J15rgG7BXGJOsPbywtxRKy8rNf0Oo4I38epsUDA1NA1gCOnohrbMlG2aCm+YlM7
7MiTviQaujoCxUnZDfanusyCs3H9lkwAeG9eXQdHh2fENvvkm1XuEG7vNuYGdKQ4
UYsBvjpORhqIlvToQYIE4pKpDvqYyzh9w+/KkLFLcpIvGhdFrjbmKwW5eHmrus4b
a3QCFD2Zxrth829M6olY9Mn6Oq05E/qA8eqbwy6DV1rxZPjozUEO4pS0KvU9ZdYG
epdpK/eNIa6Qc4GjX54JcujGs84Xa2PIkZLUuGL6IUOA8Uc6nt83/f0WW7iYsPeW
UcCaNpdz3YnjHuiqzG/3vfSgygt0nEmLNNICKg6X35TIhdGhfhO5+cEQ97WM3/g3
9pxCpcyTBXSdg2eeqky3uIoJwANjT+boRGfCkB8g9wJL4aEegs8WgPMRmFb9yMmy
6pIlnayNxomZC/dAP6cSxdjUQ64nNTpmxCQNEbvJaAGN55RHu0vep+rtMcryj6/8
54quQ5pj8d0FN7Pz9Y3d1ZKrFeNbtSLo9z2h5urLarl2WGyuCyOx1UfDdivxHk3k
lj83GdtEzscyqqNBSk6BDQtEN13axNBTvBYz+xlTasDUFxtLoIw1h/203G4KGeue
WwtogdCidkBqhHD3qpI3WbX9l+p8t5ZDqafqtVDhOzLjlHOvySGA7Jg/JErNUljV
knmQS3HhMkSshi5qU/DUmMLRZOXoSPk7z0z0/cerCi2uy36d4/tcxOgvQyylZi8s
R8fjhki381kBDoY9s91EN//VK2lAu/dcZq9iUP4cr1t6L3e30qXe+X+LX+OXa8En
L4J3F4+N9ftyUNUzJRxCzZ1c/O3wNCGdyNv2HmfJTM3NPovOv5cjJngfylnWnn3t
QLTS5yX4iGrJu/bleI42YbKLYMyuxdQgJDKhGTfUGNImjYB9uL7NzfoVI2ZU4yQs
Ki8GfitNzOCu88Yp4z/nO0uO+7G2t9OkbXez9pG3fru5UaZCb5TdSHHYyiKdA0Ch
fxwfTWH8gkp/IrDADg+ZVv9ZCoSsEbSSVKGTd7VCBjCzAMIFS3/1aFELPsLd/J8B
3jCNiTNqxdoZ5PE6NCSxzQY1aKV8Ss8hvmRdk2F/x9j+Oj5pZImGvutJSkqHn1NG
qZIakf/W1yxUXmP/S0fIrgmorMcFLxISpW94Cp+E6Hzx4mwymUxY8sNpiiuqNmKM
4TisnsDpq8JXzJSZZxm5N60GE3Q66stE6+xIFlyBQh8LrdP1Zh/UWLYknOo4c8ei
DUtqvYsdYWQO0tj2zvV0DlnuBcF39CK9iJjWopwPFcSWj+b/h3rGU99nfGc6E8V7
lCSukA1jlCd4XixgecVeO8ooYrLWSCZTRAWwLkj2QmuiaEFJkZ3zMxnH+1+UjlD9
L3tDA7OGOqqF+FeLhDXetsT9GySVUa0MT8TOlLNYKj+L6zaoFOVlinb4tx4+OAwl
PeBg6JXbwVLjBDNMijeeRuuJmeNmaq/FEQw/EFVriUjlVZoyIYG02qiIniUJ2oQ0
ATCMydKctPl7vCxGKvEolTxEnJxRglRRMWK749339q7SOeD53r6i22AcJjAXPlJO
D4dqvFrTU9P7FOIRjH4FThBzzYCa5x382i3YMtAHXo46Rk0OokeUQoYCqyq+uJcD
+5h48baipK0Wkc2Lx4IY7QonCw6pFyuLx/e/ZcwjrzU9fbzAfB/qu6Pi+PEpqddL
hQ4zoJVGG+oholfbAKItCqoDA6D32bPDs66BqefSlMwEh7QF7HwdpRGCIU2EYTWr
FldO6Mfvvn1EgkYE7pSgjH+E1TT6HpuC3X16E9zEnl/LD2Kzb54dTMzrGq+Ixo+g
YjOpiIeM1gyzUlRaNQSg4KJWOcExxRM/TUQH6WaRTunUZqWe/UATE4BuQZvOuKRI
j79JdDZxxpBywXlb6LQo3q7R9DzbUYJ48uiFx1LtdukA1tvocrcf4dfEbZEF+Nza
AaMpk96HmT2kw/cMWaMAxlWtvRBws5EzNy0BgAAysBbPeuTL9JzQ1rY5UbLoz+Q+
zGBn8LO4AhJ/rFceO472jBavQTsxpoC9C3IXxohZxo9o9paphRNlAkPEn3rr3fTH
pW+bl7A30ZVEXGurTSvqxBrdhy/dxotlBI62n52hdPebB9q0Qb0hQWGWXFqFunYl
ZnfjuL65nGgwsZCTVUo89xcpSlEPqKZdbFa/1pP5CkkXW+az9Zgim+9hgrSKJmXz
4YfWDeV3RDZrlLPkf8C8YBJy1LDQfWT2t9kja4qYVrEMePvKYh1gACGpsQySzmfP
+pWLVOaz3RM2BucsFQB5E6XbCqF325S7hzwFy5AaN2Myc+UbAylJQ1FXrj2GLRei
aSlcFWqIss1eC5N/JGf0ZdC2BYuExUF1oULasew2RGgtD5peP5wJhBBos8m6TKRr
XFOWroNVeh027K9nxVeYQZcVJHpVAv9Gi66v8qrDl1yUqegU0DCsQfNet3rGmKrE
RDfu7kbaXyAH1d1yrx3aWqydDiPwSyqqzHV16Ky4KEKiUxHocUxT/2XtjT/0/56/
zkZDLjFC8garsDKnBcoGc/hNPMpr3P0wWkebOk0YRbtBhsCgzPMJllUw3BJn84aU
0gc5goax/NUnqTGMj+ijFJ07Oa7gMPCTT8pbzwop4zofekGIuwu+W4CeFeteF+YE
GS447UQfE1+4XEaIGhdAbLYp4Csg7E40SLuc9YUGcV22/K0eKr17lugkSr8Tmo9z
pux2xroBVL9lIA5BZWzk7Brg1ZXT84KSsTIOCA9mg5Jf6vzJiZWn4uy/bXife8FY
Q2KJVY9bOUpfaO+HdGKMWUHLDU0sla3Q5wUrSKf1dJ3b4Z1it2Ba/s/1VtgLQIvv
WyC3I+tKNkdizZ512Y1lECHjJ9m2O1Of0Js4u1wDcST7K0jwC3zrizpfx+AbGw8C
zqJZg8qVak/Wm5VlOCGUNlFYuYGWgZUpziy8f60wC0Wsi+KVlqrmQ/ttBPkqnMBr
mfumC+gVcP9cI1StLKdYEvdNg1ZAvYAwGspkbxHoz/B95mnS41KppWNtXNcX/efX
oJG17H9yf5nQBL1BABjTZ6fGBItFkE8ButpTv+ASUgcGmK/FcN3uL+ddStmigPHa
6Z0hCYS13366thskUeiW0v+Fnx3lN9pXkbNrxOpN8RT2juOkU6en0JO1StMbAo/3
1DlREcFHpwFgEgFruK/5ci8S1QRfFN/bUN14Y9yskjMDjcJQ6W4QN3wsr9sWhnhz
3+jMCAhccEM5fTRESfyfrj203IF3gUnrtn/F5CDd9ef360Vw6aa9tE0pYZzCL0Do
CfWUayCAoFG6NiFK6iSU88CmnAs+SJu0UPflCe3DD3syry2NaFsXkiOWhKw4+GEf
irgsXW0Kc5aC3pLVXHnnxZkQzPu43pMJ8OmPnKtRbtudKLVMhysXWD7lNzjPZQMK
c0ToCwf88Gmbmne2n9TR4VcCnZ9mo9OUqgk3qBqgJBIgOVhDYUyaqkGD7En/Tcm9
1dlHxpKFmbsDP8+63y0H0usKGluh0EW8t8sfHBmxsPO/GoJ5Q/zB58rzBOoXiz1A
Jln19MPGpyQ5E6Tya2nt6kZkN1QB5GO+J7SS1XVtkjrngbddp//FEOZbt1J0A/n4
94MxPELvlS+X5ZHxYlthGsP1gCkMpMQl3e1UyI8bTSWgd5icO8KbhovNGEAx1hmh
+xVa9GWMBdcxXUvJMv+3z6b5vgbihu6oVpf3VZstiHu59s8746cewElNRxGPOQ89
BtwvW59GTrQZ8mRrxVabnCygkNzmy80HFGyCMVsX1HYL9435hHS57qwLGdl4+cng
lJ8ZP/FGQm0jkrlgfbM2RXgP1sMsgr0lG+xxNJcmRZusuLA6Pv1CroW+CGVdbxPd
KH0rRBwu07J3gpwNRLe1HZCkCl8S4l0VQb6zWWiBpdM+72/o3jllykuaJF4BQWCt
ps081TFlAww34xrrHB8HAA5OgtwYQl+hYiymrLxPKtABIWApov7Fq1wXBS6lSgHr
LrBhJ2TkJqatY6So8XPIg0FaWbm7Zi/CnK0JVEdqutxGo3fzin63hVS7t9Dfv6Cd
Hc5DtZKX5b6E7o8kMnM4tsN9/fHcRLyUWcTIzDQ4FU3TBfHMTtA8jLVyFIpIVAJz
Bo9mkEWoBkenPwI0hxNiyRI3894E/cLgC2GTwKkGRWwuK+7oQynXGwGtif0s9YRR
M84eCuSV2yQprXXSYxxoPS2RMlbg1v/96RC+oORNsDFlXNRCJqOElI71gn1ipeWL
eV8yaYqWITui1oSM7p4MCNK5txDdaNTBqVyNtETGw6R8g5w43eOSVr9ephlmoTgy
Ar39cCphbd9TZnGEMR+Rj9DWL20p08FEQsuY30u+oKktSfDqqt4pI57kISMy8Xy1
bGwYQFqJx6wkR5A08+z1wbNHFPIVS0XIRgu4y1wqQRDb3cz2K2wCBxzHXO6OyrbT
2KrjyMDNEaMb+rn0HVmC3OUPyyqcer7V/OtDmXWDexsOo2baNr5dlHXOR3qxRZm6
JWZFLKgzHOTdtiuupBJJqo4QNt43028cuX7/hErUiLvfIZqbeqtIe5jFUzNC6jlQ
yKychy8VeReocUZ9THgl4Gf7mzO6o37JP4t/kxeGrv15wb/rkZJZtnIKy+8qZwr3
yYKKgBr2ukMZaIeCgUg+iv8CSKX7y3QetUVxpHiTpI3pwGULE2GyQCda05ZB6l5y
fVo+O8/zdKcIr+K+Ydl7ghbV0z1SQ9Gw7le5DBv7BFbaRRJsf+efcZDfLCUjdIP5
J0bA1Z9wBOweoJna/0g3RFwm2HgPnGONeJX7xdehAmWMav2GG1YTJzy9E6YhXyrC
TOWaoM/NpYL11pnX7dxBPyvIHS6/B/A5Jb5XaTH+FHvHWYA6rorhv33Z6hQa5DOq
CUxpVbpWXYd1hmy5UvTgX+VeKIybdMos8l8fW/J0gQmALjyNPW0bCbUXFQKbUSo2
s9550VpPla3b0d75/Fhyt5JdkfcPfzadcbe30rwdcvDX7+6+QaU8mgk6iehdop/1
u3ifbzQsXo8hOeKHB4ofE4OKoYzTzKiG7NPsaS1OSLwKPMdkWpJpca0V2B+/LJaa
u3JqCGerBI8uim9wxMsQq/Sxo0syzSmewoEaryhSmaFJVfgX0NklbzgJLpS8lc80
/7rYXm0epiUyc6w4Qh6XlGR6/eIABGI13e83ATsmZPyLRP5ZPeYYASU2rbOEkC1t
57lYj1d0d2nG2MUsmatzXMUHmapwxxqIxFw1wf4SNY8IAO4OAUGTtwJOC1mZp4Sm
Dtp0QQLP1JZmuEFqw65gAfnz7zMUzDn3whgK1k8u5fFk5JZa1IfPvCfwHThdgpLz
u6mlD3txOI0gcQ3g1D0WrwuVGV1dr2o+XG5yPHbDEM/XVNGFnrG9/ECltuD+QUW6
zLWIVUPcx6l6kgILNip0mrFTwjzuxa81qtJTh4BlSxmcyzG/oi3gZ0xpF9iovXZb
Epf0Pa4dAMiXfdLU7JMORr5W3yicCPAk6fm+TdU5FQrGIk/r4QdhXS1MxB7DhxBJ
tam0gn19OpxjQh6e59q+BARE55/cHFwfS12tbAmaWd1xUPwbexfdfPvG6xDJDfVP
aGo9DA6M4CIXuBguqDqsu6wAR5atTnfsTsiQWA5njR0wcsxSE5FnQyl28zr0B+vZ
7FJPIcQpHhET9y0zg3tabqQIgSYx1iC8PF1MWQxtyDd2ztC059pl+2mDIUTiLkPE
30GkiY1cFr7BMgf4AkTxMA4gN3cxkpBZiHJEjqHDwRSWfISlOAmQO8tZ1qi3hySy
E9yDvBc4SX9h0/HuSpHG5GEIl99nQ2cuMPhKz0K1w9HO/TKVxyg9XlhG4wknlZYJ
vTi/4LKu/QqJckDK4T0flLnb/LbgKNiKWG/b2Pv5Eh5JIdJgCJja+zY2R0UFVtry
UoT5cvge/4qhxv4mCMCqj+VQBRpEG3h8/jEyw5v6NCf+8iDiuzw2vd6xwhpLp/4r
5VtYFdGd1liT5fsu+npG9XxV/ZAScwG86fFekRpXb7G9X8C7WH5b1PNq5C9Xzyt4
DXYRtvMy7CufdxJxHqQqyM7YLEMVxhG3kvP+Bcet21E4ZlHriifC0A7AG7PZAs09
9TDQH6t3L6d7o0JaFSD3WY+VhyQVB33nfQvJAeZjpgo6CwQQsL3vm9p3yKrej1VI
TlRzJanWhQicxlTxuKTlKsscPY97LZemCorPTWsSMVyZYgaaciHuRRuMfWjuuY+7
UNdbxErpvq4+hCfJLDBwOA3a0SxS8zrlHJbT/1nRfsEA1La9YGU9A4cbpqdcEqiq
XlQ6Ll4byY1r7BJKWD+twGvD3yI1/2mTrCIeysKTvMkHhbW1OXlXp5poko98a8gn
I4BBp592uLH4jTyhIm4v47Wx5OfZOM6HPTVi1RESaZXPLOopMsBkkC1+4qk1E2ij
PxUPUuwZcxec9Vmd90s9uDx9JC5ewPBhQP/s9cmkJl4R8AVH0Q2c6Xo+Ax3tfKal
Lb6ydI+zk9gmh+TjMcSxNgPQ6c7NSTw+01QsIrTIEOCs8xM5bR0N+cVsuCLd5zQ7
Ag8Vv7La2IwWiSmUXCC4RnN7s3t/1NYrodqrDOZuldzLjwIYVntAYfC0qClsIG7H
cDiKd7TeNaFsl7AUx2X7s4vHpExXTLsW8Bsofq9JdcKfYsR01VigDocAbb03KsH8
tkIUk80BTG0UjWAw+WtAS0FJqgSbeC+mUWiDXLcbCXWbXdzA4yPAV6LIVEzi/DgK
HNL1vYWDbL0VWsMH8Q1XbLfYTtF++QUG0QL4WBWpvsIzPbIfuJjAJX21RPk6TCwe
g8tdveC5lI2DizB5OqRiXZ8L/mclOpSQjsgtzAkFgr5msGiu+t/CsLXakwebK7kX
nVSpKiZaTpXciOHIeTdbON1KtawBQgKWldkuDAquJJnYqsB/jPCAZoas0HFi5KAu
DzTOCYgmzqTpZu6ZNSHceyYTKzHhJLkxmoeRAGYr2tx6jaKc1c+LLfgdaFHjvFz1
EJWYI1HKHg/jGSeeaEsYZl2d1KtHiaJnmRsfpFMxkmoSsHwrjQPAAyhwhixy/tgy
yFxCXdV0jRcpNnVeHCLZSckDdSyzgvA4LSeAzcy5PP68HhX8XdBScKipWKbH1jFC
kuFDIOvUhfzFAOW+Bq5dUd886Ll4NZS7ByT6OzP8zRdxMcsge0mWgrEo+IoQQK5j
ANQFY5sDCO2wutCOaMRlIkkkgBWXVz1s3cbNLVz0AT/tIk6fG25NKsDbuI4oyMvU
3dd3DFAxcruKODpJxrq9VfJGucJv8yru6sdiRM/mDl2TQX8nENKGY0H0J4P3hyB+
nSA0ZIA0s0VIBcIttC8sCwDV8mSLRIBNCirSWaZDY9V6DsyKjuiqx5fiahBhVVvh
pk+frEQkWF7HgZ0vNRupf0lKSpiYMmU+ZRDgN1Xl6dt8SnAVf8xprX4AW8VPwPfD
kFTBEnghLXIEE698Ju4+zAzUOLiUoUcsQ+4j4mfDtH6DLQWVZd2HHmJHynrAGpDp
su73Vs9/YY2XTdAoVFh+E3swLmtnU7w4LfIkVxPdY86OlXPWsE8n4vEyPI8/h6CB
VrA6pp+Bdn5J+WP2uf7CjcZAJjosxnJe8jfsBzHVWsNzikofRZb5QcT+LML5vXQ7
WkA1XNuVjNJR6imT+yojrhdIjVqGl5rGLeFK/uBbjorz7la+4VUSam8acv1dul0K
eb6PWatWxKAwB/xJqH08fcrTysYdkpYl+RFn9B7Nf6dnpWsS4LdyVASAeeIFA/t4
0xRIFtq/Kbo8R8cznfsqLizf6KaXTUPvNNISYP+BVvFC5IyeudcVR5nRSlTtYY4u
BRwJQo6KVBFYWJMDDM1XKf7ZbpwjNCazErApAMZepU2agCsk+l+MYIo92afeZPMM
rEdnP4ABaXkziYF15Xd1d2L1ceRKWzAuZzTeO++KmXTvxuwsNYPyiSvKCFSvjBMb
qIudbJ7jRteVIoE+wo4w3x1lWMpiIjzIJAf+SS3ke8JF83/uP+Fj8cgqn3yoFQYa
32T1gsO+79SK++rgu3iR4ODEI70mcmf4j6rVD70Jq0WN90kmYPVB9BaJaTM3/at0
0XSK1qizGJgNNrGKeAbgYI4WVzJvNSPIK3xctbiEhB4b0exCBzvBTpaWcOBrSEL1
FSyCj8U1QZSuX57kKUkL9kmRsAbEgyEifWqp0iroV75gAhatm4BCBV8d2gmIwqHV
aSZUw9bzTFZIhLSUfmGHm0TCk3ogsjFFcG5sfum0+684Mj2st4fYYdCN0zpGXoea
sN81LUE6fMyrhcwoTLyZ0Vv10AU3uPIOCnIl3wmMAz7BhvxJQxNSCjX3OOSsKkkC
jweHl14pyTzOw6tOf3n2ftb+jf8DnTSMH8eM6Px3Q9v7WJ4olf1smMDQv6H5YWKz
gTiwF9tAy/eKMUZhXOtYs5LOnZsHb6keBmwLHQehOR0pFn3pSQLz/R7NKwaNCaoz
VcyR15cXfnFJ3oSg2uxz/FvGrD0Sq1ugL1X2OwdU9uJqc2sPNQrQHMu7nFe36BOQ
zuLHLadIy0RYmDvMuZzCnMUEtdpiWKkIM9PI32rVixFm3IpmhMBWrxdF5cNQamIU
QPUA0p4qphQZc1Cy/hWss7ALsVTxCSfnSBr3kVX549XDc/6tSGPlnL31NcNbOLfe
ciS1i9KdHI+jcmY9A477R9FOR7TP/vngE5h1lJKdCi0vjHarMZEINsI0+L40C04b
HGiu98hE/nKeKNKVbX6XRtWDPQTjC3Zy7iRxVUuMbKq5LPMuw6l9+AKGaunPuAke
RKCPhF/BitauGUaW5HZ5/KPrWBq2hklvC+H6+aUdQOr3IBRKrk7Z/W3U3S9Ba+5r
dOK7d8biXeS78Nat/YfnElH1VMkiiOlDosjG49hFcn2Vgzl60Zsiz0h2CwNxbxlk
+dyNRTXmpnoZTmpa7KyDOs8zSUffbKKe0rJ5DDY76lD2ftWJDfxekqsqAIcbmDcd
5XJ2GNduqKPGbJh2JfIiqUqxEOfCab6EDdEAeSf5yGr77c6Hh9NFwZNImc5T7Ocx
mHyTMCPMUWSzTwlaPuo/CPzgBt+6S8Wi6XoCZwIxl7xpj70U5MC4nb4ALGvktmSz
o5xq7rSSfEfH6QSZ5I2ReSSaYxKUR+joCMEsiKux8cRgtHVE5xrphRYdsmmaksPy
lleT81cwwTua+7wMkimbHihOTBq+/5Df+5kYBmeO+wwneFxP/1CHr9kVEeRspBM+
iMU4baaS4QVgoFKFnQ5azjJ8Z9JlHGeBaCpCz8oC+QdXy1W1tYZkR4qus3QNoyAw
/FZq7K8P3ken0q0G8SXFd4M0a82k6LWHbf67AtDIgGEnRkp9PZ6hExK1/G3H+DcV
xgazC5cqkPJY1uNtA2YwbufrK0wT09TGhFIY65W13ixaPNwz4c6zgohHPMqbFOyx
PWu69GPhpXMS7Xlfi6kHjULe7JuJlj2n7jqaWlmoheFt+xGYZo/YNmc87OZjmx8U
epcVg0lJVxHq5Z4eIsa8dUjKFcCqqAMQYX+kgrVAdvAgksvOtEkLr5jpSNWpgmdE
rhn6tK0QgV0VRN//b6PUCKKKJT5p4MGtMcAphsmwmUeWOK9gKjmBMe6KnRmS9SUs
oVdd7WzaOOaBSDlbnqEDxwlB8Q86LxtIGdtVgrnxUkgwZM6wKBdTqDSoiGH6htmr
IFX0dZTfyIqp/j5/1mE3dyHJDfGsJLjIDiU9RwG/tDgfY/tMGczQEZZEREWHj1Wx
vV8wVa4ESN/suhMieWNkGhQ6jHqS6LrNbEOO0Yyi+bYmGwVk/Ea5p18Om5Q9tXOx
d0+PJOWRGGkDCtZfVbKF4uWtyKL8L9bV2ithgCauZeW3oLQNezWTJrh+LfN+bEhj
szT5agjh58RjDfpOdApL8e7mzp8V4ABu72aBZf4kLlJzCcfOAf6kANwQabEBV9qp
aKqsuI/zYRio3DL1+Vue4ND+E9WtCVOAbw76Z1BlnBmLPTjX88E+yRzF4B2e7NIk
nVZU/8YzIs5UEFmiBVtyju2SyObNDh6L/SSiU7CSUs0kaJURWfhCHh8EkI+UrEXW
CJiUTCE4alAD1b6xUcSPu9+JBjyHLMPO708oqJgo2xEWwqGX6lOVJP60D1HD+MeV
8tEE41k62nfIRoXTMMQd2b1juABD8vJTkqrQP8pfEacXz2dYZ4brFh7KsoUvSQg6
5EqvOAKpV/zj7JxJAeqR0X7fD3nZcBg2HJ841g+DsJY6TTEXBymOoB2dn6h7j4dG
EHeyghtrvdRp9u3s9bqADsk/vt74NvN3DCxMwJsLyo/aT2u+Ri35j6IAcKb33bln
dKMDn+T4rOa9Md+7EH8gQzvEutWwimPZIOxE4hbwflac/FlvZeInsGJynobe4xgm
VXS20mmcjA/2CDkn4Hoz9XyUQi6RcNw9694/7X7KieS/iPAyfci71KGOWUgWb/jN
0hkGNCUE8g1vgrDuBdjdTE5Ld5MZ0q6K2ZCgVz9lT5lR5NV56+fi4hi1WICwncrI
Y8ROxHccHCJnzm4+Xdxbm0uxhzHKznCDbxv433EdIaBRW8P2PPXeCV984JfS+OQR
LTx/yb2AM9rMQlgBdTm8OHCc/1p/bZk6CeHupM9EUPjjzJcQAX1BUtW0UEvTe3GP
vc2UYMftsH4SZju0Y7Ny+A75WWsrvKBCEr8lgIoz/PK7egbDSXutNeJWtS1ckDsP
ZU0+YW8Ou1ou1zu/RKh4EqRBvLey6WJpljQ4nTAAhxGarok70zG3/x2PQ2tsmGXt
ZMtacZMex2sZJUq7tWuEqT9bIY0GiW0/gfBUEP0oA2YZlSXalOQyWYZmrbFnomvp
fQgdKWzcpZE45aM2Q3PuJL3ctVgchCBoNFT4/ymWupMZV2FdjbalfuaZxa9cyeCR
oktZvL5ek8iTS0yGCfj5Qc2NHEAIwyzxPSewI+hVcNWauw494EdjCS4XGdo5tHBv
FDiEGF1USJ7DgLG/SGww7dMJOQJvj/3F+Wsk0+Nd0SOMiz+wKF6ZAiHjpFUizaZO
K8RpWBoBL9d2gFjoI4Xars55e2ndElTBjk5M6efGIsKYsTz6zN3J//JzZPfXbqAR
a36QG7x5wjh/vqs3lgwbKj5WjqHi/0tdGC9rcFNhLK66qGEecQ4qxptFcLZC80bd
0mSrhQOVU4Ktb/CTDvMiSBpAU8e9PJWOeaBQSV0q1tRBn6N/5Qn04Zg6WTHQzlOb
xW8XUflqkDmNOcSlUXYpGgjLov2b7CgJ+zod0QZa7hmB1W8ivpNOhxCYRdNmfzRd
1L/oYUPn+zrxsHv5uYv8RpytN94G77GjVsT6b+pHUGlAi8QwS90faJ5JpfjMeyOL
An0GtOcfg5VLKWhtoXFN7PlB9HCuNsy3Pz79BCMK1iFDT31AgHBha/31O4FvnJ9N
R43jdmrIV3d4g6kOdx7ka0ZlHKSBpszqHH26In7RS839rgbukc177iXmOgCTV1mk
A7iOlrSQsbcM15/7Q3QqgIOg2eAZLCKANYGNKcIdo91n7jaYRyRKn3R3rkIZp83T
Nld1R35nP5q1q6nFHNJPJ02EPAdNY4HNQaKXZanM022QZUhxaNncJ/TCoBz/+yL7
8Y9QS4+VczA6Uv3WYyVt8M3RRXx7PMVAH5aML9Y2HXKTq6N5t1o9Q5DLaH/V3vrb
GBMoilJrGc6GJRsL0PzGiVYAOOcZHGgQHeaXn2o1yDjpB2K2EoCUy1tJlkg9Uf0y
+5R40D1067VytQ8fw5lWLWl9LQhf3VZIp2owWh3VrilQC1Hfs3qCYWEujKJYG7cq
HNiK137odaZGs9WX+D9M/eKeMsPS6uK9LCdBjg4YjUmuQsJLA6bl+NsDNJIGb5bO
0b6s3lAJpw+x9lIiJmbq+teDl2LMzVyTmPoTsjTZSSolHkSmZnRaLRezvl5qlGEu
YS10Z+AnNPKGSAmgvA+oeYRStIfbaJBfWq6sgb3A01cDOMdm8M4ou0gdB9qWGDRt
0c3V0sA9GpaD7SMz/qkwbOXzdx3oppo9KQREUL91dwee0YY4XJiobwZWxaf9DM57
x9Uo/X2hzpn9d1oMdWjG6m7U6dlc/uYYb1SErxAYrkFN5rLUfDoXCUM5CbMiQlQw
dTJEMfG3VtZPjCOT7Y43sJtmkYxO+xAPceNyqFoIXkQOq3OkTYQ8iy8mc9iybp/f
hYxEdwUfDR5tlRIf5oePRmcFZ8EWWVJzcNv81g/6tzKilWj/SluONxVQL7bnBe53
rSbQatFbpo0LRMJu7Qt08fcLB6l2uLhq1KBd5M6SuPaLMVLn4ZM2rj6zKD6yHQdJ
7xM0WG00dlhrVDsBP2kDYjpG+DOM7f9fiVo5XR/kLKSYbvtUTlGwy2ZnvcVucxSG
uV+GIDZPJdZPlXJkObdMqtyWl3voWoYi0KZ0PyaQmf7B+NvRdoG0XaLxWxrl2HhS
+MUmKFVvhRcAl7a458G+Ir4NllWrAEADGq+rwVXxuOUnjvneaO+wxAaH4VxEy81a
laoogH0rQjs4CIiD6k6wpT3XK4wxmJUivpc6Z4rKtVdbhM5r7QuzC3fThZ1eo+Cg
lO6A+Mjnf69Vb5o0K/soPyk/1IuvYAtwYl6VyV9N3/95kLj6fOkkofvjrDgHjsuE
b94WWqa+sIdvdTvecXSoBEd8ak/wc10h/wTfayeYcMSnDqzD9ntt1Vk2+fYxf5EJ
6nZ6USKANy+YqKlV207jkjmNjj+RAvuLcb/kdNhxbpooCubNiIDJoXbAhiQdKBpa
ZHgk1NkxmnaWDMG7ZY0u19oZmIy0tpJqrDPSfjrR1OuLbgtlZ5NCD9A/V07gGYox
wNEz5sTUIuzRbvJLL8sZOyjlQ1jX3KvlHJCkp4nZvh18W8OUy3i/rYhltq3y3sJV
gHNcmcaeD9hsR/636McjYMEkIiF/oyoVs89L2bc0NwCcUxMWf9xEunVleCbWkmX/
07kzYindacRewwTGgJsQe1DHxvrYWIqE46YlM9Ei4az5h7Xur0KPO6Oi1A012dWY
YhVWULnd6WUmwlE+SYD8hVVb3mJ5TUItRTq9u3ztcEBr5yZC6l9juJMk1ddKTlop
mRNvXLcDdomWI6RtfyrYvfeKlLe57y5LEImXD46OzmYXkMFpxtcMLaOIl1gMToDc
lFr9TF6d9CyEFpLcVRDQeENEzglQn9pdhIln2sYU9/gmcFp+J0dHpP7PnEiiEsiz
tc/5NMsq0/aYdCIpsJClaPPvUdM78vNErWvc3GGslIje8xCD0M60QjRplqF9MU7y
dYMy2Ji6pj3RCuuJ4pqLqvfJT1uH8TeFKp3Kkc1a9k3cMh3oTxh8shTWYWM0QB1u
S5ifrqroq74hOqnzlUE3mlpKyLioDDoNFyolSshWazik/dme8t5wz8wKpS70QwJ4
qehCJV4rUsJFC+4G7G+eEAhmUFofapZ/C2q4LhZt22NmvrD8eCoNk3FPXk0izKNm
7YWT+ykGneCoDkuoHGk331Am61dofbLBDUe+ETEZv5yUoK/xFhFzcs4wAiqpLxut
rpOTirptJ2ftw5HjFJA/VxaTI9IyH0bHhBuHYF7CJoZbc2HrvhnnitB9atIlS0W4
MTqBE0kAjYfZGnFW3FXEIC3Uxs51WX6bUMZNJOStWukzv+TrFiH7zo/XBn99b/Cv
S0CsZ3o5lqquU5bGgcQuChdJRzjRjFl0kbazr0gL8j5vHsLxGi7b1Ao+dpDvnDPE
pYTEwNwd+s171YG0JvGUC7fICGARqqi4dGyQiyPH9RE46Y65A6ALRMDFqKWD9h2I
ywUkKRNTelpENhZp1d6OT0W+HG7H4LWaJ+7bqZBmSnWgRiHE8xbvPZ663k8nGIMl
IAEsIA57El87L4rmHyO3NKDynDpkaqfmhqSDrbhDgQoHr0NPTFyy79hshQ1Ln1O7
oHd879RDoPrt2AZTDk7cfdeFkSAaFNwaCCMyrIRsVd6K3Aak20H2iN9iNraHYNpJ
Z2njSgqfP0NLV7z8o7to4ktIDiKgA7cndLTlg5mDEbqIouxF9nVMpnUzhnDzvsaE
chY5sClbyfa1REj1UfxAC6WxJPLZOmGG/5KgyKe7CM0FqLbN5yLmKMmBpXdXZ2Vx
7T/y/KSEyTdfYT5m1W15v7y9iwKyKxd37qhie8Ssprk62e+8oSttiJyfUhaHslug
20t7iTY5WeoImUpKFfXcFJTbhMqULUX671otE5+aueYxYzDLJf326RBn2sH2HkeB
ZfoPot6EISNyc5PT/++nSyriWAqd6Rx8JujmM1iJThGq/lowaq/R8VdCk2pkVbKs
YyQl0QR1vzlQrKgMGT5f1pUF17N+8wNMbIwK4Du9OXhHuI+JCyvkNUfAyUynk5Ft
DvzQBEwPajRlE58Khl0rnUDgx/Yx0TAiFJcunzMks5CckdCAADSfOTYuqYI7LFKm
hADFqwoDhynuXPf7rxxHODhkz3VALdLvBY4DygxHpiztxZsOkudYZhL1OG01aJjv
bxiYqWsjvc0Z5tCq1JFGcIznPwyQu1iZJ+r7eZVNFBQokxoa5q3S2B64DyMXfeyX
wKo6wraT8tikOqOKabtOGtJDsG5L+JlPK94pGhrvEowjSOxPZGAnMFWfOYKj7+uh
UHEvNNz9yPNPKQrpCcn/0xmUUR0S91qvsrWanT6XrcQvjiBl5wRUsYHvk/xJT2xH
3VtgN31NxjFmYXhzK6DXzMmV5mEXBz1gtPiISJ94viV1AVuNVR3qUd8AGGfrxKax
IGDSqGX3VIhKUn8h6kjVOXIGBhwcq65THopMWXPy3fU2muw1rJugE/AL7tz9vJ5G
GQbfirh+0b5fmr0xRkBJmohZeaDvmd5PDObr8g80KxJrRcAvQuFpWc5xpggkowbt
dhMW7mZYbtr0p69ubElbn8ClwD4gkdqLJ/3jzQf/znzxeAn0DjQrW+sIx7BgbOrv
B1dgXaX7m1Cqe23duc+fj62bM/EBukShBPmwhTZ/RsNwRChNffhT4Xn/3H548eWB
QBxcwdGva+yZaeH/FCLp0uqmBFrAyMIuI64JcSgtxzEM5/DTP/NzPZ/F8V/MIxMg
Ly7OxgpZXJmYX16pGa3+/7V9H4w2nDdXRmFJ4a63uz/8DRl3FU2k346KJK+V6lBM
56E0Rh6AGoDOcSz/58pa9gmCu4o62GB8/KI5nxkA7POdqXypBCCTemLIIKBAT5UX
7FkBDAEr3/AN3GS4VcwsP7ZdJvN26Oh+PcVwjXGlqz3TZJyHaOfdtWIaDUBC4pWh
njnTehbdini+s8lojEPVVaDN9yK9vgL9pbBU+LOhJvS7WQul0UxOPFj9UMsZfZjf
7xfmO3Kepvc62mT8nhT0WydmqQQ94rOedA2yL9WN5PzvEGXHSs9b3O8X0mwaRjeL
CbUPbyN3/EQsu30yo4JdIiPSYyMHygeREggH1YOcZNR11p5GpRvYl3oxhmHxTrU0
frUkN/Nz2+Uk+ltEHHkVPYMcmwIMJ5iaa1eNHMe9wk2N4HjH29o2+ntsjTkjGWwt
4d1F7TeQEdWliiTa2D88NqKKrt0xeMLab1XFBsK809d1So4bagBSIVPK8Qr+FnN5
EQXPN0VHzj+gACQ5qg7M4tm6UPOea/Ldtup08s9u7AmwymJfgnXT3vZDlpgfJXiG
/nT1tJEvCM25dou6OyvGdRVoBhjdONY98FLYsoUCqC49cRxCduSbSA72nipT1vQT
lPqtn9TyZyMpvu5MOp075P3sYh0cvjpndkcXhoNAFvw9kFo9Ru/szfDIHDslKGup
fiMfKQkM1u9JD3/6CFm8krje48NXunZaXm8sk6Xt4qmgKkCatHPy9K/5asc126y1
KMRX7Cx/uANb7qv3F1z2RYy5CP8R1l/F/IX9FYVGKN9y/3h5Da/qdvmXiBwYbJ/z
lLkSpiAG6n2s85mfNWqzxfR8/Kh0LLv+BkMOMD7gfez9ZHnlpl9U25NTOFi5cQB/
zxhwcVI2/ZCME2UquRF00H8laIspqIkn6Tp3STVSNr7viNZwRAUwiqMaPoEM7NEi
LLAk1znqLE5kZC67S/UW21DuFcCtQ0QuBjxdeIokE3gAXuXYBZ4H2Q6qjyTCxTSR
MqBK91l5OdYiE18/z1TffQCac8jN9ase+gl2cRV2/BUwr5xv6LABmVS/3G8coPiu
AJCNOY68JE4eEkSDsruv5PDGc3G7uFXTFfvwmK6fjqxtaIaIKLrwpw8889huR8ue
2jwP2WVuy/ByTIGFEBq13ocZvXs25X9SwlDI7+pGjqs4wr5/R2mD9oCSLPeZI89C
nZKej4DjzhsDCS/FTufiMihYX9uUkLrqGqNpI0VrUcTUX3D5xnNMJRIVToT3vdnI
1OGg4VKyVbDsI1wzyIFX6VDp5uPwh/R3pW5kbAVJymH5ncfnxGCFo5AM+BAJd2pj
IgiLFiMcrBUDQYUqmnqqSkGtpynPmC6EAzVA2+DgyjVJtQM4nMZCOqvN+H5VEymp
dqghPuCWmztHfShYe/bbY5B1Fd4L3tgbhsfb7q1Pc586J2dX6abpkz3WLLUTIczt
pf5LbwE2BR1wr+L1CPSgZF6W2zG4XGewQzhxh4RZAIjGFOoEOWrcds2c2OqQQChp
1nWQMJuFRPFRae0xQEV07xPF6BqKLPDMnz1yzUL+12DXo4d3N6sSbZkKJG/YVRt2
2uq+KmWQ1WRz70XHIVpMpWwdMkSC8ppNNViicNF85RrxmzGGnoSN4pGQpZ/T0vZM
AzW98jxWLN3wKXuV/dL/6tBEirJN0tZzY58lImJ269EhfVjyjzLJqVWK86qHffI8
IvzAbNi+6k/WyAVW8QaLPBfLZJa4SoP+zhbtAsFdOb7FIRswtciWS2Idx9PSUWwP
4+O0WNAQNPjl8v25H5z32WNCkLD8gvfTKfF46IE1m8rSR2QWcH9+WCNKtA4fYdxi
RJWJe0HSiGsc+nixLgRmrx1BqhHEIgfn67m+7i3QA4VXCH+h8awOQxi+z5uY80y3
tkbi9CkhjpazF/4Afo5KKdU7B0IMAnhkUK7rtin40yNeYh2BJwSrQOa68Qwc4B72
AcIBveXokCaIk1/69bkhYx3qdqHHsPWE1fXVfcrFluaXSr20nW3ywLM5F+/j0kXk
L5KYS22f0MCfnwBZGdd+CYcwIohFns+l8XLWax+cQER2xOdt8dEEDwTf9nEtLO7k
qYvyo08BZW739M99meoOSfX3apQavG0ApvlbLnZbLlrKFVmLL+Po6lqZTuhKW6om
KLTq57uaga2E8Cq/xanRqBoW9pbFfPwKkk6dDLdOduzy1190TRVtYeiyWTGWRr0U
T6QdGSMrTZB8+mrwQKtvkUhBqjD7oUtfrrZtOtXaIOwoIRjK9Pqo50g0FqOE9QcH
S0YdN6O8BYgktL6hegcIO6Q1L9GHygNGjAyEspkEiOKZrecqZ/COZpa4v7W3hveY
nZ6jYHU+DdEtoTtOb79G9sJDSxagMv7TdctN8EIxc5UwQH9QkfGBKHM6Crci3wRf
QXlDoMqeRWuAY2gSnwQXoTbfkX2w3WBoomCqFEcgyHXQgzr5MGNi7DI5EoNF/iQr
8nIbiD+S7fssYU81ZU+pVVm1+emx+HANhGDSfBsYg5uebCDLf6DSKwsdLXJu7sKi
0Enj8RMBD4VXfQzZ0bj4gwBcfVOe7Xtc1MOVycjni93EJHfwNraTUIzyHK5ON9dr
wPYBU5H8LQz21BTBvFVQGS121bCSkh98TyfEmANV36yervCCAvB1aTgwvwoY6S1f
23wJJDA7H+75sAs7+76NPjzX5Ft+rUMuNvuSD2diceSwT0i65/oA67QuWXWhU8eR
uw6Aqo/C1cwskAOaJGPcfaofhgW5345p6iQCWQryI6y68smi3i977sta8gWSYBKj
Q/m6ig11bi28O2QGEnuEJqwoF0SBiLlN6XIdY79RPB8VYmEZcRXyJrgMAkG5rACY
eKbiFR4Tokj1N93NsmGgc4LZC5eQAxxrMBU7KW4NclZ+WcHab10fznniq/IyLUUx
VwXSwM8MMn6en22uPY2pJLUgpsJeHz2kvmJ4VXIC747wMZrfbgBV5XPX6qjR27o3
WLjQrmc5f2Dv2UVmJcE2pd/llGSBWpRQVVX/VfhSHpEAWAcMKcQEDKY616E/wGxN
Eyu+G5I4GoUS/XiO/oxAN+/K5Nh49jCbQ6MHLeh70u6bQyzOkWODa+HUe7kHQRP1
xOqwubP/7WAgpWcyEG5Mm3f9UWeWeEr8yklynvyP/mjDAwoHgT7a/LuXWLoP2/Jh
zddsAEqnWXWJXG4BFyZmbVKvTedGeTPvyyUEGAXGad6NfqRry7uEOpSi04PYuXdm
uFrVmCFsn51yimt+nXkUTlUupgoZa6CUOobRL2//ll4ZdqqkPTvBaucFuERg9Bv8
c5Zym30dsUzyX9SxjrftwkpKT0+8SvKJxgdmXwRSm3Jc5862+VUAPtT4lHwxwDuN
ihTBvL5iIQFR1J1QEFRbADMVL2ZDrYYJiKC8TPZOx+prOvJlNqGIrNgqXS3XmsYj
W2In0IZaY/EQ0x98mMGfQsu7NzPu/p3Ay7dP2JoWXT3WjZqRu3b7lWykyVk5/Irc
9UqvIZqbIig36IGxSOaqEXuZsNiVDUUbvXXjrDebkofHlQVvIcYlyISOs0M11htd
Gl7doqS/0TkBVNNuggHzXddHBRTeU0ye3urI+3i9o70CvyAwDVDwhEYUQBQrc8yn
I7htDltAk5yt8vvUHlk6Tk9EMLav/9fOS4elLhJg5pC820LM09oSzVI2fNiZiF2N
4D34ehZpobrTQ9+KCjHryE7VSEkjuPQm2pkq69hnr21vrl9J1uPIjWRyb5i1uU4J
c+6KxaJCVetg3fxg+Z1MAnwUeUMG55pGvnM1mUFoXOUYKphylr/o6yRRGI0muJA0
ZjJJB5TyszQ98zFxA3SuRJcPkolgJtIr30DJrFVQS0CBsEcmAzEm38VyOFvjDMVY
pqV+p6VjCUHZzrkY35DLgWhthTz3MueyVSSyjX5eRnzXr3/O7ruM4KZ18fhOlBlG
hjkK9tcVG0YX9S2EEsSUB79bUXpMWCYSDjmltXVvOPyieHt8yqIjrsny0/M0OKxH
MC5nKjZLUDBCieqp2puVLx2WetFHlF6IMSpG7lo5lFZ2a8xTSiKTID0yfQKZNhFO
RDu5TdHERsyz3qHPZ3wMq/rI2HB9mJMa206vc5uHCZBeeIlysGJ3e5qqLOrykA/s
ve38gE3W5poDMlzd5TEXZ+hbc0AZdwKzbTY87TK5ETA+6L8gd5jQqezo5Q2PLqJJ
stZZMJ5I8DVZIFm6i3M9aQaAyN5nLTqV6+S78f5F0WMRSBQn2mZq+ptqqpvS+7sb
TcghZLCb6RUdBMhe+az0dIjnK4qaemnocYG/o8chaXvXmepsddQ1KVQWkzaCyMy+
MaWhnKVkEmIAU92sfz3o2xF9fspqxrnwPUawG2CNH2jruJfZLGv1Fgoq2cSBJVbJ
Df9w44Rv1o7JtJFAQP5TuWZJTpLBk0dVUSWbRXT3Al2DmgSVB5k81xAXFuaulT+5
y3x1xoI8mtaugh6lrZrnHC9iAQOVcxqpWZEsZCvL8jx6rraBybx8JMe+s9YKlfE+
81hNgMTKClUoAzUB8tb1eC/15LMUP/sN0VRK40HPzXa1rwxMbsyScataK/9oTngt
rDdGJnqYB2CSO2GDWDH/gSRDvM/bwOk4Xd2S9kzxxHxzdJU3/6tONB1j9ANsx+Vm
6HrragETtr2IZIokAVvNRR5kniRxEBOm/VbNpdzX5bw8v6frnTJ8Abc5qDkNPQsT
L6n6wcYsvJ5OENiIJ5v0VVlfxZtOwlaaRIoNN2Q2nNIWxyNHlM9KO/modeZeCnVz
owubKhe6q83QAFxErGcWfA==
`protect END_PROTECTED
