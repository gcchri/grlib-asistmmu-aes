`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WmZN5EJu7B4yED/BrWQPv7bK7r7E+8uwJ9A5nTsJEV9vQwoFQgmNcxIzdA/8iWoC
BHurG4G4lt6hDl29cuBajQpMR+XzvNLIE7lu8PfWGsrd/Kx2uB+bFGkTYp5RDuiz
qiqIKCKR76qBTpiXsHuNP9gj9XxNUcANmPeLJnTXhxVzbdYKiMKWRurotGUpEGTI
rtD0WskI51XEtHggKV/0XmrbUfYklhZDXDjtE9Hr9bS7DwbtA74Oj5DG5WD6TYO5
kfVyWXnKfCd88biygNW7R2lWM+A0MZid/loTO61qr9tkdB2BSsI5896TLPMOzCFF
KWE32DFb05MVxbQH/JBtFCA/uSrEyeBpzNrcBphs9Xdx4PdKE5nuSbBagvQID30g
VqNmN84NvxGtuJ8GgMwtpFHjNfnvI8KwCn0706GciZAWzQqwYOy5CaC0f8Axlxwa
9c+AKZYuowGxVXlI1ZKCjXkgWg/9+YbayTOiXf1yS/cLOwWBFw+5VMp2pVyCZ5nc
ZomJOBO41Xi+pGo7g4KaQBzwp363r2daCCsaeWDKG/3Dln0CyCppE8BjmyPGDUJ6
OU5o/bc7zjlc9lywn7D8JOoQzGklwNc+S6zB0D9sVukxQp2V6X2n5xRhDUj29ImD
LN2IhA5pOQkbVQoPPBIkMxxdb36F34LSvWA1GP5PN6W/9AwSdWP8+vey9V7SjKqP
n7Ta+IsEqhXw70I6Oz4uWhTv83vJS1I/cg3V4YsPnL5xsRdDBAHGprqG/AA1IczJ
2cIVXbBjQRJj2POiUiUP894qbLshhIMCGCD0xdiNO4wMeu4jowlz3qSFsMSM+Jw9
yzGzaeJtYeAodXQKk7Uzw7tD/okNtQnmdIvU/vafpr+/3ojSh9f+p0slZAFP+Ey/
fCJU2G2Z78dbHIJ7jQ1fP7CV7scZAumjzaTdv8PGXYdNWmum6a+nsYAlDq3Zt3z1
4iGm8/XlS34C/dugMskoaxtr3cgcjCWcXku6MrF4miPCm0p/wsnEXdxDTXmVk+W/
IU8wd3X0ikszbWgESrKe9PhIX7VTZgqLHo4hBdjloXAnhWxrmktZnrasAAPe/Mn9
FiqLOskgsiK7UPaSag6k/Ma6TIHCXcLp264xzL3+2lad+fvj/IWm3UR3KqeLPT7d
VmqujhR5X6j9d75RfSSCYtnqs6BXni3lq08KZgOreaFJddLcocNBVrI69LZ9fjX9
ACLsWggatNTev+0IBh2Ney0ATri+bQG6+4iS+t5+4zQTVFFLvEw8+xWN8Lf69OwK
/5yjjPeBZDSOcfgeC+a39htNPp1H00c0bLXnOMuZ0++/mifPYAmOXQBxqR4Tmz56
57rie7trw5+/YflPqB8YF0F+3S35/lSX3URIHQlZi2+OUg+m61pbhGtq9EuLF5jL
7krioEMqPlF8rWvjQqrf8MZQImgk0Ke7rqmZCgOUV3MkXOdbvnmUUPQYY0EMYOG0
OGvcp9Ag+hb5P5997b0xmlhdHy5+v5AnAX4/bNUFUDx6634HLYSEnarOLb6a4rdK
geX2eacQVNUkxy5WjfeUkK0isQA3gWsB+vMypNemQkTEDASQddDF1tM6VngGVbKy
KX6Ap2B5oE97lPZViA66adwLMVHEbsZG6VW4XeyJd9AE0MyWr/FmbOHeypkzwYYD
JexNNs++1ucjSNKHUGaO2Ugad41ksvOSIfcISyledR/vH5y787xFhZPxRGr0MIMy
fqgkJaS62qVzt00SYv4ZOUJsS+/bdrBOhMSJmoZqI8CYbh4NcOOzqSJmR42vEbKP
9ovhAgAExXR9U0e0NNfM3EsO5eszYh57sXldoCCf5n0B2t2hTuXXu0zcPw3+YQIP
/D0M8WPWkluy78qRjrLxQCo0EEj4HPvFxAUo/9HSoXRpoIos9pRvpoXgQAFC360K
BB7vP+GgiFqsI5Mu5dI6EVM31W5ZekimcV8j70jcdKMzw767LLqyg38MA6EdX63K
X5j7DEjOHBWmVX6Cbd+0CDOSHR37sMUgTqDpV01lqYcL8SVSyD7hNPGqAB/yaoc7
Wl3WZbmUt5guHAKGKurvyVHAL99Vmu7QQIeVyEUi+x/HYK9BZphGTsJaxJA69eUt
SC2v6z6HbRTya+Le0l3wVTe7/Wx7xlYiz6lYQE8Rvqq5FbAd79gC1yDD0YVoR12j
GTwu0vswO1vo4y8m1ZRw6Xo/RymMPs4qXx8c6uFwkelwxPtolgh46HRswoXk/Fyq
x6gEgdGayw1oTvy6bprHnD95jQ3BV+ocjGw2vG+nSMkv9xWXc7zzSmj23nNZ93tD
qOuAXDsKbOBUayp18RFtchCBEhumb/6Pw3VLD11CvQFtz/HQsHpiVAwvAdGJN+DV
R2Fz10n12l5rjED826RtaKvpZLnKB7WbaFePxTDB8WgSoPq2NXIXu4VNpIxgGRkZ
lJb6n+fJUDfISp7A/vs3xVmbgmb8RiQ/yHygP10E973rVgwbx/bjRClqnkYphJem
XWdBYp2i7VwJaxJouodaC8XdJkiO8vToXfeO3o0DLp0Pfp1Hij9JVG6B8Y6nL11o
Qw/QTGE9x+WW8b+CnKdJcm1mdsafbgxPkTiNUgBgNBNE8VGWUAvXmq9ya14inTUF
7uDoCRmgijeZg6WEE76tUVtn9OOUDie7gM9rqj+jyQL4sTRb2JlhVIDmClfQLHUd
oHJXKM7OOlajM8Xm87CSOC0j4tSeFm9D/zW0ikRou2wl+4Ez6I7Ar4YVETMTQtUj
4Xdc0WUz9zcL5wejhsZOmBghu1i3P2UBuY7itPn7mmKBiKnUTyrTJ3LHQ8uwS442
kDhFwd7BPRApy9IbGFUt+8SgJ8JU6kdDwl8v6uLeuNNnbJTtHJqJjV0vQ8r4QHh7
eGTW+Ogy8h8k990JdgiQ4MyEKp71RdjTgtVYvFKCU0jnHU9nADFrhjV0ycU9xHXx
ZhtgISGfOVaJm46jbPJpFZWy68f2YcxIMCDwAd1GK8JwAjfLiEcqjHnx/mkC9Emp
IO/89+XUVTfB9ZDE0mhwYQX+s8cbSzopsLL/71F3ZnXa3MDbm+r3OGRnUMqZ7rvG
BNTAD67ocDU77+E3w/YfY493r8Vdi9OFCKP8OzBaBQ4g4tBDwT/n3COKBLiMbGvS
KxF6kxdv54Pllc9nFkTsKhEPYxdaK7Xoq6wQdK6f+cLL1jnga5ZnLxhzeagtxDv/
v6FYpaADRl/AWoLaxXtUDFt3R2StlkfR7Qigl//6agyDUoRBSdRjq+rXxDUVbtMa
3THPZnGrTvY5xL9YVIiqFZJ9GCe6ia2l2l0MFHz/T8A7fyOGv/Uf31M7I81UbdPk
1KBZ4v4UyUa56aygdxGjfjHO3+QwLUmAsFP8WCf9LFGL81hBExt6UEAoBH9eedeK
7+2DzE2NXfMum74aRl55+YcHtckNRtGrMWI3fEmYTYqJkIKZP1JvOdlnLsNdMOK7
RSoiK4cI5bAkWBkZoNkZouI26IDxg9zu3gAc03zITBK0/SnYNPoPxYUDgkFoksc+
trvnSCANPQ6JRCr7YFna9gXqUwdv6altsIF12IYIsdUbjaFmRgBG4ZtqouGclPsO
nKTTTjJMHP5236rg9mJBUS81uFQlnF8n/ZRg4SHo/tG15S+fC+nkwG0tM3FX+tfk
itC4mvFFIVul4Cl2QL6nBSo14wTjq8pWBSKozRrMnS7t8O+WmWhop+khRjDhb8T0
gyb7UcbmsiqiBwZtpPaOPhdoQ1E7ImMbaP06ciL0Pscsz5UiSQBDd++NXJYmpqZe
Q7urxhFo4TxrpBzkQPQeG1CZ7lMmhyfkqYvWondvGp/39x++D/EGIJui/X8ryxTq
IOexNLgdMQlR4PwDjlv9fwcxCJfYT8OL/rM1mE+zyDPIZiuEHv02ilkKE47G211K
hOYBUzEQgO7LqrZWZZrHHykkqvssh3Hm+YAYD/Nkj+mdUpqBsz8eOfpXjypgNAni
4TOs+40e+oJsDxwl+bXsaDCxD9iJXPPDuecMaY7DDr2Tkxk1iGeAD5oJyRHwSXXU
mVYQG/5FdT/6RJv4rIIFjdllvxY8wik6xkf3sS2tozyyFFI55M8hG+gAO9F3bog6
LA3vtKJxWX8UoKSnq+EQMZrsc9WhjagdKrBa8H5g3wBkYepH1d3ltQAv0ZfYlp5s
wl07DlWckfRmFf6Ivlm02RPkZAk7BMQOPxS3tq1ICLwjT/QVFHzkXUrh9RWEwJ4F
Xd0LmLikG+f+hxOgNmBPFmXT4EWcpQ+9IdAoo4gspYqWOMFn5G4BV6Ttj82AwtGF
VH0ZlH0mE1hiUOP9Swr/YfaXkysu9gsQL6pw5QR+YYUPFHiEZiOzakYIfytToDzT
qIAE6YKbV4KRYryiK3S1vUxGJ3aomtbqfpo0ze0dGbvFADkpdQbgSVPaMYK5mQSs
uYhto3QhyDfvj/rXz5JmKoJSim6VuK8CXPW1rY+sbumwQ4hVQ0WGila6y7PPBJMO
3Kf03TeN2rVwwf1pqL3CiOZMxSneux7s5TLPFXHWT4UNT+jS68H/0kTzx4tvJMLt
Uts+4mIb3fah8spLUHCwFLVldX5vYve9419UrmveAFcoDREy3lG5JMhdLVrWEbYq
aBLEZ+kgQCOVxumE/5Z1yzurIYO3yeX9pv7sqvjFcvp2ha1MPuK7+7V9ESR7X4hc
IclClkvuSQvCxumMr4dzoLF02gdk928N0Qrdfo5nUjI17FLaHnY6MI6UsCFCHBuO
o+xNtUoCEKMzqICH3JIh/nANN+KZbeDBsAMi+7pJ0R6rZ206S2hNUWRUW+Jtobw3
oRffF/Xl9Zg0aE8W5MiUuZsHy6EfI9mt9QOxWJdGAYfmr657+hy2C3sEc2jNjz3d
CEQQnLunDXbzjBxwNME1leycZBONSdoMlT7eesSvuobQtJxxddZZX4DZcZxoA8/r
9DU3fW9rMUH+QrJcSpd9RMdSigRHqeFuIWuQ5iK4HFqUC4g40Tmzq9OUhp+83Pvj
Tja577MpnIMbupN6Z+M90x7eT/5uFO8CxxAsQQn+iBgF9ydhXzNbngQcrGMMvB+I
SHsGwkMpQRo5hvPVi76bp2YS52Y//6C26NQ9VrOH+CU8PSMjuYL55DDfEt/U69Ss
f1ht+ct9dc5pkPK9aphqLAUfY0iphV5JjSeas5j91qgnbSE3mC/QTZK7A1bKHzbx
1q9cbXdQvuxdHgKRP10NCQFykcMdsXc5BTvY4+95njkbgs5S/HMX28vjzuza7NQm
gkFTuUznWZhU4Z4Pr18+h5xELiHc8+xOJNKBjbT9/ojK5XgrFTHb0R35K1CX0pZX
uVj5RGwfj8V8tp4exCJwDroMeoC3PFTdGDKyaujoYDbHMA+5V5cpJ8jJBfIslaWg
krEb+mm2CHwqGbAFdLy2Z2xDfuMTny6w8Set5VCrI/JgbWqqRmUN0ECy/di2YT9P
bEp+x/cwTLjaUuVVGVNHYMNDTXw0F2zG6jh5X/LoKMFr4qpek8bLWI0xA5zMH9w5
uhZ/ReksrCbLWdwg94TlJwDaQSelQQLxAiZM/bB+BxgnBO3/9qEbwgFhUzg4vy2a
2UUP3/52axiP8GR+JM/v/4SVD3+exEnVf1wNZ/PXtnmYKnQChC10UMI/FFD7cPal
1z8wsahVllVFFk6rWxM//TJdnxIVIu56S2BuWJhxu65oMvYsf4qtleVI0VZmv4OA
bMCvND7wog9kXmSqBWRDocySVq8SPG2FqbLZX6vueohRP1DueuWymE6VK/3Ef8b9
AbM7hlT0rJI0CXlmE/9mTspZJvRGGUafDgBYr+KNoYfQxUKA+u8WgQOBu6rnld0/
Zi5lmswgPVhdxf3PZfztt5Lc32Ka/4ud3ajzyNA9588aq0ir+T+WLHFJLxDPAn1i
mt05JSEL3OUgiXlDBfi7WVDZlBAGaQTqZEAcwrA+N2hH6eJJ6Kw1pug2dIjMJ7EF
phqjBTAl2A1glygYYSzdjZrLYXZNMpJwG1Be6AWT1V5i/v0vucjxycdlHZtUTZM6
CIAc9tZeuRPBrugQVZVygrqw7oYK+r/hc0fS9SWIsqL9BpTQdXLExLNW1YMGvQRZ
NuSaR/AtuoUsKoEliMyHufz859fE3lJSA6ctqrmoKVY+ax2U4OhngMWGyTAb95ff
pMXnTalZJehui7w3uXUjuEeo1rU9SRHmgn8sOfK9+sfoggnQqLhDfMMGcC6r4ngz
eLeDs6V+y6r3olpM3THtznpjrfznbUEy1/eztcAhhw0h20mjG6tZL8XziOIYpFhV
Lb7AquFv0oUxJr16z9fC/LApMuNFa9HU45Ijaompd5S52sgMo2Ilti7FSms3Grzb
sJG8lO7ifEw3CsZCzQzW3URAZjyZtXFBsHGwVC1wiV5+45UDzflc57aM5hpyxz1g
GHt9HYnK6/a/g7qyuyoGHrbn6KQwqr8so/l43+/P05HrvMoDwcaybFi+UxCkZy/G
lc1qjMBmG/M6pehQfkuc/SuQarfHc8i7BAifc8gzbCKIrRbL7aJfWdnSo97AjD9p
JXr7tjf7Iv11At82Qmu/6TlhSnkLyk4Ci4pqm/9wPRXSJgirKtGECNx4zoEgDT1e
lzjTNmdBr7/yrnbBmyiPhrLvu9xY/k2x3qIj2xKMevtiSzAZbsMSslBj4s+pRTSA
xZbb3e3noEcp1sF9TxuGDVz2Hr0Hn+0jU9MveqW81GRIHRQMydgDK54/Q6R8PYGi
a/+astSWOtFB8ncjqJBk0Y1Kf2/xqMF+Cg+tADtRy6b5CHjBSaLIcR7jM/fZSUGO
7WNs3jt3nlsK35vGAaW2KUPSmBxyFKHdQGZWOfQu0HjDrzQFXpf0wSOwmA6mgZx9
MOh00l0zP3DktHuKs1ZrZ5XEqJUMMs37N1kQgi+NKbpHJEm6P8MzmevvlWy9k2o4
dnoeDANdQlwiBdK6Y1r0F5jBolt0MmYDj977glIlRfw2PiL6/QQxHpIQvvMS4z1/
je8iSCdkkWeiRNnAwChviDQc/8HROsTjoTSwhPI2VrRTBUFB58rgjm59vxfD8PP0
CcCBeb+bB2FUqGyArtxZCnpptLSMAR9eofKcuI8RH0tiup6WMjVtAxqGlZWbp7s1
Naxrewhh9uVuPvOALVZQ1UoLKnypjO6m1yFqEsgvqSz4jMZYyLi2F7AsrFhOvbYg
S1S9aDRY67Y1hbBLXcTbqpTmKL9BppzKEvtP5gaI8E9NpcwQ6wbAH+r1mTybrpXl
f6wvqpnHFBNSOu2QXhDe6/7Ts/m35CmcqofBsajAtSgKqDQyA/3L+DRODiafkpkk
dIS3H4waoz7iCSpZjmfeDW2EUO7hOh3cS3/NMwC2OugxptZulFOXTlyrnZ8LGzSj
qQvlUyYfi59I+QfRDTpWZSO3KqvDmyCLYAfz0MNLBH9od04qLJiCNzj0UaeBOmWR
Z8wdOqCCBQ9b8y51M0/EYkTKGDkgtmhFxwpLSkVieL6w0iHSj9QLmVmDfCClfjQr
rcuWlkVf9bs2bv8PI6b/qI4SlKRIBVQczR+TMWeQWXlnrL95knI5qtHsfdQoFZkN
Zly08/K4L6ezcxIb9yZb9ptROlAa0gipJe46g/SgvT5UEWVx0vkrtlrbSSEsVQFP
ZiJAVVi2u7fJe+CqlHyB8jzqehS91hACbujHBiJVxYAbkH4PUh99SmpvVRLY6pHD
48W/qR38D4zy+Ri+6CYF+z8IcFaUNkrRRJQnBeUQZBl+15aVY2FClEYS1Y9JqEyK
TRl99lGuaRMfTQCRXkfKe+FO6Ljq3UqIa1JLubPru+qHsQGHIoOCQLjM1U4ktr5f
lMHVjHc/UkqbYHoiCC5gm93u/rY9WNne2j4sDbp78C26hgPwL90jhS6TAxJiHtaT
tZ/R97LFQwePXcAQv4Iasmf4dNAaIM6LEH0KtisWR4kjh8FunUTFpjkC6fI2+reE
xnehmRtWMdPitu67luA6gFlv1dBnSBLVmPepPCXjH4Bg42EvUNgN2JECz9wNMSXR
oH2GDtgKz9mim7welz+SuF7EVKaElNJDcLHkgRJpyhN2tSlfFtVEltyDXYQ0FxbT
iMvtuLqrOdnJJODWCliLItwlTZb5wOiWOxL7MHuodk46RnAdkxyT8HONuD/KQt+P
wxmU4dV1t1kyKLnrkcjwjsMUL6H2xUC1A4RBqLuO97RJkNWyou5Jh7yArDp2mOdS
sV+MJH3t28ydnvDhMoQ71ai1n+j+d80vZaEZAxwwzsHC4AL/AA8y6wNahwy2M+jD
a3tnhT2toKkrLd0IeSNFQDx5010qkuQNWgswdI8NQRrUpzrAutx3pRE5HNifugpB
1qG+EratdJxoBiF+NXAjl/5ob1NYV9U9NjjV1GX7DSpgCZUBG/asCQyNuMOxrprh
JQYW85m2arKAAVzb366m/Bln1d4M9DcVUEfTbbcKX1YLqOGvngpgGid4kVXpMyug
kGQam6r67ZoA5gHotQgH47IGRMN4T7byjK8WDeEJhyWYkI69ekA1TT0BivsRTSQz
x08sT/bbgWdUG+L2hWCToojwC/1OAAPX8XIpcHY37Z4vC/Qk/vAfPEuVSs+68yhL
/Gm2VL2kn8TZALZRaU6MXqi8OXoZxd/F84sK4Ne7LDYhnKHzs01v0a07wg8sNqiz
w9dbzkzJJLukpey2MC9+MSeLUWOtmiRyhjVNN+diZ3nrRSE9DyUvFOeR7AOL9GNe
BThhPUU/5XAc6tv3sOQI68iyjzOtUYcPV8UUPjQHFL6VAjGpJ8pfbFbazMJGt/9g
8IxJN9esfk52qFW35zZDLl2yykjwxkyD7aCCaqYkVR8XltBy+j3Yjo1TG8nRx4Tt
7N7a8Av2+6ZzeHaQGtXQAm3IPXjQ/2KbX0J3Wn0sxTlHaUNA0UTkSagnjFLyKLZu
e81JIwxKG6aNEVJCN0QTt3Mx6I4tkzCfwLKTdFicxEMjM9+WL93jdGgq5r59WW3Q
FRUGRqR2E7EoojaFu3Nl7XJt8TWX+mY6pqyFhdItDKDJjnxk3Gchfx4cETXAWo9W
PSFUCgqqXMT2js10vTJ9+fXHYYxbKS7fXmtgJqlugp7BhxJz3j7Gay+9LrnNzxUK
pPvstwvQnk5ohcwgI2lh+4H/UX8nhF8NGWHlBgbgexEocNAYdb//3Dkjq8mC0hzi
ae3v4NIQpClO3cJF88ZQIIID8b3SaK2HXEP/RT9CAAEXXwypMw9/cPW+q52GOP68
hcK8dUDgL45Srb3BWQO/adxwxWYI8lDuNd6D0h2ppKLlIKhpXNFPg+vUaG2OWZLT
rQrBx9XG5W2w1GSnFhCZE7zR4MFa0TwYiyqRPRqapCti+B4ysXkuLfMzuh/va57v
VQEopGVht2i0rudPxqVMyc7saDhqUK+tYc8Wt7478wZe68zIReZuUoCoUTItFgg+
3V/rH1SGEupKRwQ6zE7QUyLaOWvz73UA8AVkzTVsH1aI2vhMs5rVUdvWFjsevSIH
9+kkYenf3ybXfbqeWgrKugeilZdL3jZgS3ZtDwjVOAXux8LqeTx7yVds6YBkqm+8
THKrgcuRU9ZJX7TWnPfEaSwc8cPMNmYVRb5kQkmQ3d4fyF0TJM5HICqA7RhyxsUo
QV8QWXwYkSz1AIjzCLh3LX6ody2OC0GFfGu3OQpR5OtXD0aC9K/xBOLrnFd3Ck9z
zALcH12UEbBvuvIANnjTVOBBBrEat4ndrLvaNxBSY0gK196Pojrpn6jIUxo5ABJK
pPdbZyxzrFASCJCaMS8dGYx+TQNTMUdBnVHiFadVkfaUjINK7LjltpK8/yvYV3mO
MNOg2L4eaD7S8shAn0tuxw==
`protect END_PROTECTED
