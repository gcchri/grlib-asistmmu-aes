`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LwZIAeMKue7Qengi/bcZAH2ceSFNwwCS/epSF9o7QndIV1fhiHbba0GN8uoX1nG0
VN9GeDEt3gbkeeFOibEnw+0xIoXQNWkKHM/o3Er44Cm81+GVSYdb4xM5ljAgDZhJ
g0GbGHFcUXns3JaNbTqfwb5wPX0GY7cTR78tOM5Vc5HwDRAR4oloQZYm+mhj9c6G
PKjgwz0OWYLOv2+XgLEd6yFHtcDSSQidtITT3HVzhmHsjaf0hrT2JgJjWi//zBYR
43QA7gndcQMrFd06EGxV80NrJu1jBGn50yaVbfsSHEwfqJrjFKaQi/NkNJDYQo+j
W2htQTkd3tTsgUSReLlNbMjJQptzM3cbRxGW5lJeaAt/aYPrFWwoBSsLd/erh7/7
pnSOH6IaRqZopssNr3J/ttvEWLpGyMOGy+CsQXZcc0Ec5kMJMKi8BLmXhizTvC2H
k93F8dASQ2BtPQY9d+aLhI7QEu46spgT6q19hrF5MOogWc9STCLbTzJsKW52Ecl1
yMkckbnAVHYYpHOUKoAbSyJZ0UfvIXded5fOfeyYL9fKhL2WO3+ZfF92LQOZYLf2
kR1NiaPLBACapmGeWnO3MLpBrOAqsWWYPb8w19GKycV7/FrNLBLIyYiqpJBFWXvF
5/mQL/oshaZnl84+7G6bcX+WCLTg/YYwpaZz4V6Oz/0oMWhHqVaEJoOw6rV4Q4B6
m/ubm/zWz0FUXhjuF2SLUXgNl1yl1xBF8h9vlqe8p8/iCnJfxBVXR2CgrThxO/Sy
nfQZmLbOFGjMH5T+nBif+4bmuUPPf0RTsh1YnuZ68FvOgUCJeaxvpQZTy4mgJ3eq
cXHPrAhR3nvID0dBbyCVmaWr9V4SJ2bYeHzUK1Cun9MDGoPiXMV9tEu7fvy6iM7X
vJOD9i0invnMPWVpT/YCvsu0Q2sbUr7+NEpklUuXkf7udPROSKNEoj8B1Z4vNS72
qJU8z7XTlJPrOlSRE1ZiR5tjkJ2K9t+O+bbNEr5b42T1KcK+u9hYcgD34fVXMRCH
nA7uH6BaIfpvfMnSLgkUB2163Vg1wgHjJw3wA01DaqpGl6orblFt/EHcX5/7ettW
gzsfYHjFRFNbb9raiGJyb8P3UAFUFP5wnMhlC4H5sg3dhL3Ufv9zPQciQXJrWltQ
xaMyPYhkzQqVk4knKUet/HAbPO82/7iRMFSf4quD+CbFL2H0PHHBr1J64/4qV3p4
wq3Z7vxUin3rdYxbTQGlTRpMvlqVBVSTsM5mpSRf5AM=
`protect END_PROTECTED
