`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cbCi2SbhLiksRToz6I1YcXjngxm/Dj7h+dixPLe/atmiGY5GZIWZBKiJ9YhtdNe7
IaycFujRUx8/g1S2Wwk7JUyPKM929oRRJHt1cmWnAV2Jr1Gdk21OhcYl9o6FBPx2
zgWH0n5NSy+WI/QRAWquqtZgbUgHxxSp6Cl7EDTcHF+9qHZkTGUcm/xLSyBprevz
XP5ztQCTqmqib0K3NwdM9FZQ928uV9kg6rNi2mNCtQvP0JXN41gEw2wpaQfOV2/y
uGbmtzPsRN+PZh26u8+KwpHVqmEcEpWjmfuMP0uLiVLZp1oxnlr3k1llU8FLcMmr
Y1LnCF+en0gUs+1UXtUQe09H2TOIGlejuc8J19S57wnha3U0jetJncwJQI3aRPSH
1R3jhsoPerI7K5tXh/6udCwmPHKcMO5NJmh7PdxiCrY=
`protect END_PROTECTED
