`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AGX+3LXltHKKvFwkV7ozqcs8jyGm0qcnlIL0hJ9i9EKFzU6x2lgyqwXhvKHcVsyT
SNMV6zHPHOZ+dra9H+fLifcaitEmFe3cM4psEwhcY1oPs21ttfjMx+SGPzmMbWv/
Wy4MlpD8kFeUt0fZSZXGLqAHYSk2lYOgc7C937iKod+D33i3tFNzQ5bV/wSl6SdW
UjYXbW6eVRzlypooPx/7rVpajoh4DAycEWZopAv588UZ8BNxbmx8qENnAtIHZvbd
jmzFzKKHqmYtbNI8MEHECBH+jkyOvHoW8YN6r4yO7BhRxdXGQo9dc23IoAFFqd8b
yyyQ2In/C8YYMeZXHTYNRiivb+yyIGxEeJLJB9zF8r5B/hwLZdDHGnDw5uLNW6lK
4BAvx5NIDpZ1NIwgDRRaFfMZT8XEhxqdXIA1eAsPJhevgOW+MxBrDPOJnb6veAVq
FgVLfnvcFzKTUXES16UKGCMmt/3kX7YvqqCeSx6y8YN0MbHlLu4Fu6ft3jX6cI2P
cnU/EPXg+uQQQf4yMAOoAX2u3oP9QD5IMiDnOnEEgxZYyfxBqjpN6cFQnMV/8QN+
i3DN3R1vpRV8KQEkd/uM24AgU9l692mnAQFjYBRGQyewwQbNCDO3CYIb4WuxRIHF
9PJwkhiNKA8UWaOEYo4zUd9XIAIRZyUA3+wrXFvmzVkDWibuSp0sxL3dgk/FHebi
raPoiHV0qJgMNZ/BEsic3Rhh112YIgjNu8rmEyHSSNQnzbof2oS8DswzWnqfED5R
LsYb3zcuEGaSuYW0c47ygvHsjYKEtpSTEURuOCQ+mNw8vW4M7Z3a4MZnrI7bDgES
Zp0cexqyIShHsAU3n/kyAb+T5wxAvxiKPqSzzjcPSmHi5MSO/nS4nJlKRnSBxfs5
zEyEw3JvzZ/3h9pjvA7GjMjOL2e6Ui2tZIKvrWl+FU6DeCbVLOO/ABF8i39WpDTq
`protect END_PROTECTED
