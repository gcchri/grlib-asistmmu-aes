`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BKgBR/sTRyOj+VNqYI911VwbUT3gbUJsvzh9//iAbwxzJHB8VRsgtgGzXFKg6xo3
T0HSzs4LiaXiesxUyvDpzKIfu97qu0cTzdTm8a6CpO/el0lhTvdmwE2llTWB4dUP
KOUA9RWa5d3diihfdiO6fL4W+d7e0xiTk/wpZ4TFNzDYa5+Cp/S1XNginwKgqy2l
vxyuQAzRjqGVPIUTUszOzPLXY+mUPm7ZZzcQFNOPpFehXWyXJv8pDAwgdNlRUPZD
rxqIR7T83bzBK/S4l8zkEMQKLHrUUTP/S0pEZCKNfDDmAVyCtmjJwRX5JPh3RMNc
g/N1kY3lWkmte0ikfUQxTnHwd5gFO2uPkve/IeWCgFcKaj6waVvTQvzCKXwXdDfb
jbCEoylwnK6//en7W2Lgs/ogeeZQOIlEumKM9tmDccg=
`protect END_PROTECTED
