`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a7cI/2xfYgAgHiqmXe59p+jubUQbPSQ+laubVS/drliETgJz++v69MkQZHDUO/fp
PWT6f10kpyzT27pFMn4Jrmzji6/CWEp8omXQJxa8UqCUQOMrXb1bWm+2au04rMx7
hNbyJPeWUarM4VaWCkLD/bIS9fI9d5TyZsa4vTgaTWAGhRlIjGDlH5m1qEGrH6An
mCAPBDwh+uN+a8cr7k0Rh8GcQF3STDnohT9jLLraHakLAbQruxNb+42PW9NmO5QY
`protect END_PROTECTED
