`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k32L+fdQHCmUEhQLyI1AkYCvbFiMKvr4qjpPEdAwVi2uuERrw/kwMNu4S/3b7Pe8
6qfRgygB9CIlcSKBXPXi20HMh1mhwdXH7y0s+txYZnt7Rj6Vb/vshg52Qm79gFyg
kCalbyKtwhJApM4EqdPDwpg3xcf4VrdX8hO2JySrnf29dPY2To+COWks6Ysnppf4
hzkYv/PtLiA6OXKxW1z5OvgTxVIHQWDwYnSo0a+AxEx1aIMqk9IWyP+OwedlwfYY
612w0wsuPqufBNlhArvgClkS37fnf+daBBQmY8f4+If1/emOAh59CkwMbgM7uf/W
gCq/XO1b0Ll+2Eun41JJYzKUatxBIIEvdpWEqHRlKevRMUQgmv7HqUSnLn+WLRVX
mNtGB6cv7MBa/7DrK52b+8Q4HVwQ2QwLLQId3mY7CeqRyorkh+urDKey/7wNVVye
Y+PYelqut9z39p6o3UsGIKk47VusImcUpDVRIYwN7IdGETiwWWGiVk6WiaGfnP1Z
q+KTjc9HT1VkNUspA5V30yIV4E+33nK9LKNteuPgHQhs+llCivoTQo0cxkkFY30T
8qMpYOByWp8i7UHMvzLZ5RkmXos6DJZTFBDIiuuU2ivDD+jP/Gwovp0NIcXX0iJk
8hyE+1wwSGJroVNdN/foGv0rCaygYkToIBC5TSl5wk7EKZ6fV7BjlBYy07F4QLsx
pToKvh2AvCP4dY/jqcMjHrpPn8IEbuKBUarICfSo/kTyRqZ2qtwYYcMqFWu7sLrF
tMZf2hBw5GAAz3GanTD4FLND62IBX+PTzwntxiOqJILMlfGPEvRrKeYqKsgfdamR
VF7+f0PotJnwJkzIxcX0LR5Yb2t7g47kmQWoKXeLPxffy71QW3EItD4AZilZdoaq
LbApKlvuJvWBxTxnLZjKuwe9IX3PYHAvshX9IkFfNQslOje9+K+ABaSAFlbRoAZ9
WSq2FnK4lIcKxVCUPwKCziP0B5xfNKbtK/QgxAocM06n4LkWGUARu+9Z66c6OOMz
q3YF1NI2aKKKdWIbxm7D4yUFROyEmpIahMXIbz9r+f97I5f+o/ta7LbrnDYP3Tmc
GtNB82NiuvPvCB+rg3NV9eoq7wi2JWh3z4WTN9WVl6Kuaxdtssv3VeUtoJI56ORS
rG0ceYszfZXge3Vq7PykF8joPSPJDdnuJTUyAI7KX92TCShXDdoU12zsoDE5Woxj
ChvBIdJDzQCwpCL9WFUQ6pjwgA44xI2AsAZXpxP+t/qtNAvR8Q1SGZ7XKfm9YefE
`protect END_PROTECTED
