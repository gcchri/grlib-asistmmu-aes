`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jsRw4TLhIWoZe53h8SaN0CN5f6+CMDC2Gwmj0d+7iiHCKSeEaRVVGkBQl/Sqk5H9
X4SJd21NOG/zHmhHP/SXOVZMs9kvrUkkXqOxBPtTdbsin0V+LGkeHQFxzC5CpUUL
37Ki0iFz2aNFt6ymScrB6c6plvebaJCKfoEc+mgmNSoJGPP+vkkk9PK+0/p7Zefk
fYrJDZMqOOQibQGICiQKsRZU3LqiUahAm4P6+lTX2ZstC7oHeofm7k0KhUqciT4n
YxQgqNo8k6NZrYuAgPy07Rdv22ec6Cn6eyaTdBuP+xF6MIJhAEex26STA2vuu0w6
VN/hJ4YAp9LhnnBub1dTCg0qiSo9V+ISxxeslFyLAwdMzqjvoGXIgAfMMYE8V+cg
Mi6XSMJ0f8orYbE80w8n6dMqpjApN2KNRcll12TYUGurwLZIo8aeXQyRymjyPtxm
2nzfl0bTBzfgmUHJT7O07668WePChnmGH+9pClzTbQg=
`protect END_PROTECTED
