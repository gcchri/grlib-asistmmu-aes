`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZnOM8BJdtSfWtemS6YoisSVnJMx5+gRzfoqHgbQkGTE5PaCqos/jEa4RnGEni9ij
m39kZPJA2Er+agN92Q46Q+JjgUP9Gz8aCrJkQYuYNn9t0Up905jJ68Q0JCR3ZrkG
pwM3fhzSMBlWt54tSKQOQWYaQnHTB8b51uN4DW6kYAPKheKKs/xsmP43S2JrJDAf
TojDP5wg60YBwmDOghaTLd9xUWNcmLf2mQQO7hdY6mpMgA0/yKcqEwNSi7vlvwRU
YP1YAEhTctWyROWNTVp2u8KZqd0QOyj1CjhYlPt5K5VKlMqFarbq3H7Gm9liuUw7
oIOmqrz0Pw0SiAQcjtJZ9oitsb56U3MX1UkY2RZj1nHNgF+f7goZSQZkwriX9PRL
x1lGV2PUTC4Emw6LZJI52k5PGSoHuUyzxH8YhkQnaIiHMc5akZ5sisVoWDirZxYh
wW9buQwILd2d8OmBJhv8RTxZw9MFh12XuMlPS4hdGL00zn7MYRYkPcRr8dQ786QX
eSe+BZnooesdX6IQIiNxoyX1Tq0lFVuk3UkL11lp2KvdCmJouaMTI9PjGs1YHUgB
4aOWcDugwaUfZiyBLmh+gq0XWczov7PI6XiAM8T1JllVm/AOnlqu+FkGEsYzSAiy
0dZJbmL9gBJR4dy5Skv3WKsMMaKlp1oWn9Z1fTi23yAIkKjDccdG8JvVE4APZ+wv
VGGo9FObPpVbhWwezwQYYul1jE17IpdT08g40X+wPszNpj6DwvJ5FO5n6tr0wTY8
hDP8nz4XufjZpIM0qaQCIsFWcqtzR/rYBBuspNNVeS/HzpIgefhxbxOm+EC0iHhn
v5kznjgy/hZ6mAxfD+26QSPPLHsynOR+ZnyDaHiPm6Mb7LmPadOdsr8SOA96RH4O
xuJ9x/nSJxXAIyJlyxnUiQ==
`protect END_PROTECTED
