`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/NkflydEZZkyhaCgYy+zWswE9NFw3dv85hissr+Ymac8whMDF8bko62J/UeDmL8E
Ldq2juSLmHu94yIaxdHIPKCGvgCE2bRnHCJ6JZro4n0MYFlD7Wx42lWw9mlwj9yD
/AXGsety9gAru5ujPulQI9Fv8GILpc5K+EZHPh0Hhk75nhcOP0BBD5MoiGrJRqs9
U8xg9srkNelgPLnis4HqH81I/seSB5rqRolR1XarTYdzCUlqpTCQOsFIDruJufPk
oSjiO7olGdehfY6BYXD1zKoDf0Tk/deVCBk6JlCGMBhpemSuxSUYR0AF+8gn0fSA
bap2paMumYwpKN4TpsK4AH3KwE8cbwnsnIrJBkj3jSZa7Jt8eFAGPhxFmh/Sv0SC
0eRFg6Ml33HZiboCbRwfCg==
`protect END_PROTECTED
