`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kCWdeO6+n12nT0wfRgwoo38DEu1MsebouvKBaeS6G4cyZgR5FQvT15MEw1zSyihZ
onHeNhBmab47OMgJ3K0WImCNrwju0BtA0GngUZVmzehOxbBKlba+KT7hMMUajBEm
gXs5FppS3nDRm31gee+teiankwn6KuYyGi6IuI1QmssJ2+caeDSMkfb6zOsxlg1T
TnYQnWAsGyRQ0OSCURRxzyyL0w6oxHFiXw8C0gIJesx5aQdTbRHBU+DMkNDVJR93
AzvZLSOoBGS/NlAnc1kGrMSEDDY9Lq0uoWeumAkonYAeaOEmfpchq8uqf1ubuCmL
zFGwFcsjv1DNHiTwKKRVWASQTOXHOBMPY8iOaO+T9RqvOQ5qZ2CofIb4OrPkhmJi
UdXBsezeDjHDRb3zJrs+76r+493D7iaWpijNU73QWfwcCaxg/gLXd8p3DHnCgDET
Ej7VdlAeqw96TVVyAyZ3fBe2Mooagf+TqKGjQE3jtJgC2nE6O0RDZotB2hiRJ+1r
L4ltPASVxrn36Rw9pLQKNwLrOb54/iH6j2jcpYxlzDvYC+f61fy2TG8qA0fTo96p
Z21SdzdaXDM8janjbaFQW92KV8iwViIWtmfdqXteaRwyC0dzEKY+gikYwK7wkX+c
`protect END_PROTECTED
