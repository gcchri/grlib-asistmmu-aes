`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bEnKugvjA4Qe4/zLU0cZAHJo+YCRo6UowUkm4aUu2gkoyNIPlbmcJCt+6QZCt1/7
MuyBcRC/GW149dizx8KTunBTvKNXYhge7sRzbw0ysnsqxigSPSWWaXZP6yq4ELhF
0kFeoEI59tM0kE/+dxpoAjtpp+U+5DpXxCspwUakaIVzcPR6WF92tfy7zW0MYuN6
1Cr5MW8ynONXVqiBwTaNGn8O5OX/CM1Y/7yD8uYTSJ9FLvhDtsAnqpfY4SwNECJR
RuqYKNW6whPsAaLU67bZdgwsfE+g05dwwsgZla5rNZK6Sgg+/yzoTte6E8A20u0h
ck58q2gfU8XFedGkWdH3BoagHrM9MQFs9CJjQBXsYohD6Od1u+Mx4EQMrQfI8foD
g8+DzX7Sv70SY3IXdSwvqBJdPThzw6lQKEHwTKMCnERL4Qm9LJwF2Xe+qguwi3lo
ayOvKFbYJxxmzbnkOkIWb2bZZT994vMsoG1qMhbtGlavWc4Bq4eekZbXv8Ssftps
IxIRc5pemJXDDCMeLy+ILnd9FY7daRw4KhDKIgVKEEI8+aOtKQRCCOmH2HjGBl4J
JRU0mx4pP6kboqocKfwOUnG79yDWbTB+yBaUHvrrgkDvgId09FOLkSoy6H7AwvGr
SjNGn2ushKhEUtyrPucdeg==
`protect END_PROTECTED
