`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ybs2rkNiDpnwOGzOwm+/ZeHSPc/YNDWk+1nifFS5Q4yiweqERE2HGj80vb4smgA6
OQtRcUIrFnWyfyIStr/Fp6elJcfYfnFPyj2105IdgCoZf1/0Yafhgkw+sgJFZhRs
TunVt79wZs6uusz4CVVajroRuTflaPCpmKsJRQSsr92Vt41WnXliEl6+W/eQUWd6
O8qLCnb3LAPa/F2V2xcSL3xoZyHHM46opvJNw6L8aTXlEY1ByPuXQoYIPYIAvh1h
DsuFkqRmcPaPqzmg1ZMBLEdcyTpbKjMiRF+LxA2Yp8lBNF+tP9HEyBEo9CuTZuXy
sQfIezI0KVn4HwTPnHXxreqPE/EMXi2hEN1XTx25BP8=
`protect END_PROTECTED
