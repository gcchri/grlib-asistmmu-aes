`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LL4KgsenhFp5PpwuRdK8edMYEbppgA1YFzUTaMiG0zOVUAMlFfiSZkNput5YVJob
hg5bNlELNruOWIAYl4czaaiQ41TeTCATSMGmn9Reu6zObzdCF5EzfEkTgbs+j//z
hxdh+nguFMHanED3i8HWZyB2tZnTu3PJSTDzNyiCum8ECaovWFir3TRb2+0EbA8v
0rsYglFxZulQ7g55C5UV7lRG05lTG42l7YN5q6+PQCXoZM7dHrPtIx06hj5YuCaH
9qGOJRpBjFgzIx3WmSELJ776GwcefXOgHhCFUHQkCFkQ9GUiFhr5xRNQ0KNGKrd/
WZIL4bmrW0aHAFPBA09qQxplHJAUdURVZS/yY7JKN9DEUeDcAUgyd13sj7+MRDPD
hFja9fuhaFc1uMzrISmTHw==
`protect END_PROTECTED
