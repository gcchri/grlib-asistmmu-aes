`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NRcojGtb9XlRVcqLX9Ai3ka9BtwIebmbuuXj/Zpw5fCl+y1Ajw6kN4Z60lDCb0dS
ULg+AlUX/wdryJ8g6JWWog/ZykBp9t8HZ/sbn7ggK1JWMNbIHNdjNolktUfJaAZk
KRMy9u8c+iixq70m5vkOEOHHqUgKdW8vvYYyBy1gbGH8pk18asVg8Xveda3sGxwM
Q1zXN/PdcV5flmj5wG4kbxXPfjR4ROU5Oj1NBJWZdQ/jUjpcxVZzHlzeVakGDahz
JXYKN9p0QLlVKa0o0ievj27lVoU415W00Hmwomz9PHTMsXisQs7yqfvtDlA2sqlr
G8bUV9e0E4U51yiDdW78cm6TRwHppNdaHxcCmfHG1ZYymMd6B6c8y/kn09YTpS5R
TWBdXym+gnwxsVova86gkaUE7rWJMmx3G7mC6nU1MeRBvJtaOQZOtXWT4s5NogyF
bp5OHGZjpx/DMzrhLf9IQhtW8l8D9kDSLI81j8TdG+C4Rdl6DweiLztb/Y4gvB0C
IciA3JAM4odKL3Lam0NIy1Ixi9N/KYmvdP2VnDRsUtsj8V5kTzFMKwqjqLWBRNx9
aWiFeiyNNq5FxzBj2PzJ0HSrCF2S1okd/CRdrndrwC0dDBx4e2MBUSOZ5TOK60q0
B3Sy9voFb0M22ogu48clBBOJ/emyMiRmzwG/nrSDRnvqgqktFthURTxVXQU1Y/VM
NEmqGUUtW2HgOEtvg/RBpIduzeTdtQPQB+zRnewG73yXdUZW5PUCTkzOjrC+Kfa3
`protect END_PROTECTED
