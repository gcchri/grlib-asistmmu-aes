`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xcwi3zdHHTe0KvNf7WaZWrz0ZyZXfuUKO51s0Z4Rqs8VjccLXqQF0evhyN59RW+u
mejM2CJ8zW/DP3iDxXSofZ1qgSdyLmtMHjTn1RxERBDYmerZpTuOxUW7Tr1D6Gy2
CthFptkMvpFrqauLSKa+TMxvGKdyMlp8ehNhonsFXbX2igTTfSD0Z7yUI0Srdbj/
lQkdvNJFqrSA9QrRlckRRbdR9Yq1c8qkQVlSbxhIwnxiAFFtgyHjn5UeEDEUOcSb
poj7b/blDOQCXm/LzmbKubPUEpb5soeVZj0hpL63mKJajaqoOEDKPuzYdAMOhsIb
v7BSOUyocI3a04IUmuDHK0pCHN0kcczzShj6LjHenvigVaYuM/9zuvq82Sc0wh01
PXpxLHUbwBA/rdupDwBhpA0s3hGk+NulgdFhy/H5MWkLiyDleEJIyYU7noH2qaOZ
aI1e4xamjnoXD+fUwpF45Bywf8hPLJ1lUI+jHs7PP2odVUSskcy4RLw0brOpSg7e
fpGtYhCYIH0lwJl6+GJPZBAPxo5rug8OasNVroLV9phxFRgIUjrdm+lNz6Yp/Hw4
vLxLU0MSs4vW79ws5zFEvz0uw2hbSX7G17RVrxPnLQzwJERRMIWZkwDt8GzAVfcb
DxpMM66yov/mOJzQP6P0AcmRYviNKxe6o/5T1vtUsfx/cbmNtyP31XYIchf5G/X7
DOHs4wwX4kGGeBQ6i+pGkZzh7pVdxCo9vbVqYbhHH/IhiW4BkZdLfl4eqT7SEyRP
pMmzUywXpHgCBEdmviNm9PBHhU3XsfEcrEYCv3U10a949iLiUWVKTc4RlO5Pud1E
6Ey61NPgcHozyBTogmzC0wr8GpYu9aewQHqbTe6vpbtaKA0XyPUKX+bifrBuMwKu
zv4r3VVa/AfL6BCgs3ol2ZHIxN5U9AFNgdlC5dhm8HSeQVIqZW1IXCpuEzSFnob0
fLa5ooXEnHgCgFsWA74SNfVCxfwco2AKTtmE0tMKKVVjqKmCEj6lr29PR9uE8h+0
9kR5xXn8DZ1wTcKNjzXg72Vue3aS2ZdqkpuQbMvnwHbQnk6zbfBAxKlN9yi5KckH
Q4S6DSZz+Ua3qaAzCgnKD3WMOr7Ejt/QiUqrDr2sVYXjIJ0lfhuAddRX4Uv0LWtT
EBSc45M+XdrHk+FO1SN6lJ4Gmt88+oVdQyDjvZ3/ANU9x1PFxiedjaNZAGZryQgQ
8/eWhSv2QXKX7cYjYDuam1qGy7gawtlTpzKof5KZpfpAsUobx8YAA4fNDdj20FpH
8Si9tJnQj1ePGczG12sGm+c4orCDo/GWBnMrtJqKy8CDo2vUccoiWR3+lsO6CNhy
`protect END_PROTECTED
