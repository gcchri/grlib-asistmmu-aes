`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8IXVR37QAdFAlGx2dCh5+auJBA6/SqPivuRinLxCgDqmIhnvcmGjMOTz0a/WeVfz
dyG7h7PIujeEgaBgCepiou51+6JenUcYSHVPJYykbPoIE9kc1gejmEjhd4u8WFrR
70VvOIUxZssNYT5s9OJRG3fFI3zXpZSgwj9ighYZp4vc2PXWUfHvrgLVAHAcUbn4
WTuOwUqRWP3fG1i/9xhsG94StdCzBJ9l9EUqQF3zuGboH9xwbkbnT8iYHu/uXESg
/4oBT++QU14G5cNynCRkhtKBXh8f0/aPVtb595DDsuY7yl0ZL51rumi5FmHoNT/2
6/9Uq1yD9339O1+qyWmQfQ==
`protect END_PROTECTED
