`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ySW+k62ufXc5HApj8e0NqdWpM0v0R5QmTngLufohBUSHUjNnajO5aNJg06Xv/hBq
WLeW2SQlV1mF9AAhNVXa81Lqemj9E5a8ys4WCb634cd7HRS4kajpbTcnbvpb+DjW
Rp1uGScAl2/fzxeOWqH21scftw4Udstz5+s05qPaDkzvStUD8LJLvYm5h03wwboa
/2a9JqNPZzAVa2iXa0o6rBCaV9pjfJfqdKnb9USor3Gh9CmPs3NuvmzvRZv4Wj76
7daeuF+pfCYd9cZI6hsCVpHONVXgvTeRUAcyafEfnmaWtz8zZVzeSdErjOmJCPVg
MWJMOlOi6aO0EDOqW7thXFZbz/5bA5vfAoKOt7MvStlQ6qJv8jhPICYi2j5Bz4IZ
9ZfUQeaQpHx7ouHvtCGZasPHR54dFMWHM9Dwce0S8gk+SQ06z5yrIm7phEZucs9v
aDwaKLRZc3UNGHM8JMmqXY3f9aGmGGXMTntwSa0zXztxnLbCIwpb6Cx/mtr8vIRu
Bt1aQ1qFwQNrpssgJwhUOjZ7MOpDFgl1kFkuG5nYhgS1eaxICubG9eAqxP1gW6kc
9yaHnjVHx8s9iBH98Sn35MQ50bWZehyf0/TFZyJxEEBqB9zU8ZTswCLtn58K+uLU
CZTmDpllkCCu77zZRergYV4qj2wfzdhfaThB5sbHK7iz2QWMPG0bgO002SEVu9oW
LhkKYWb+s0NQg8r+NcATa3n6VzOxadlE7AWLBiwMe1+YoYHPsoHIFZuYTtAora0a
ehbw/SAnJnTNKzLdslKUhwm4Y+VLzk5e3XDs8QNfTxeouWkXES3sRDhW5eftbgxr
81eOcEFyHBnNR0cEqrcaGYzeb66+J4IukfSEyveLrctP40gy68bvNrWQwHyz6Wv9
NKAiSqRJJiq6Riiv4edJJe90ZdZ9GEUju3P26BdEv0ddcfDFpJ7rw0IXFyd81xih
Ymk2Nj1WaS83fPjFHQ73Ao5O5XnaiTm/hDAMIwf4E9ZrB/W85nYyEbfK0dOlmyVX
+i5A8EkrCvVeFX1kNFoOhOELpcgH6Lkw1P8oLa9PlJLy17YjqX20uf79XNMWMwJ9
`protect END_PROTECTED
