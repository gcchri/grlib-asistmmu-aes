`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U145VsTMrb7HrwnXKyEDEfU+SfJqI66tEwgWZAGbLrIK188HPAFJPGVsw5UmB9xF
q+33xhKs7Rg5S5gN09SIiy8G6DudgGt1nvkwruQ5nF3zeyOK7pzH8X6krNwEpwPa
kVUH0AUDgLnj+BgypMTfiparJc4QJjgcqx5wbSYvrLPhoiJiARtiIX6F8pLVJfN8
XkUeofxxs2WGTjndNz3Pxb7sU/o/UNYw1DOQQYONFNmDCaw/3u/vqqsuvQxbeMfq
iX7xcqeefs0jTlpRYD+IWRPwy/Py/4V5QcBUMK9kF1qaxN2fnkCfYYQPT/DjfFnC
60Sh6499Nd43lflyykFkv7IC8ik4UF5ftJv/1zEwtBmh2ddH9ZN5uPBvxjWSMDwD
1uzFRJD1HBRKci816VC5LZW+urtC9vPSXFScO7urcblJmM8H+hYZMqv5Qjxv/3wC
VEj4SxQdgtSSzes+VsSJn7I4Je4KZhsffQswwzet3ACH+Lq1uhUcHL7ibnVP/eGk
hFuA2zJfnZmN9ohtjhJkbMq4DmnwcaxcF5IExTZO1xlsSGgbMJh+Jw8CF0Blp3gt
1IDXUxsJdjFCbwCm9vsNffQQ6FBvx97+U/KClnhZYv6eKc5lcaqS5LU6JOMP2Vn7
Su8+HYDKvJn4q42t7ClPp06gSGTxxaNeF9OLj7hfo0J0lIb92KV1gz1XkzFHjxtQ
uToW2Y1zvaItJYSPT2m7BUdgBZ+TeDh/upKR2cRKiOFN9scsC8/+VCBninM/x9bw
6lOrkNA5fwJtn8PUbnvIfzE91HcltJHJFS++w+nuUtp7NixiDYam3U0E2R1mMS54
JEZMZwdMteCW1go1B7JRuA==
`protect END_PROTECTED
