`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KofUcNWfwNhQvavPm68ZVRW2VScSMnmCfRWFFHboZlk8sHaLT+IwRgKnyZkPEUpd
ladLW0ZXE4NspuBND7brU5X/H4+eieoNaknKZoVR/osApQCX3FPeQOSDmUmPDizW
ZawqegzaYx4EN0Fax/emz7bynTbfGizGgRGhMdCkRGudmk2h75AQRXUdqUWojPmK
zIFwui+dp7MUCqQ1OUNkwhI4G9bRRE3hBBnCNbVUHjJgeRB48iAkL1kT3ijTJLx7
SKPO8Bir0CkuJHYB4cuHpebJ9gNUMLJjsh/WIa7mgDJdpEFz9ypbOGGwf1f7J14q
JSOcVVUSN75t8Ga5t4bPvQOy2ZOiOdfpQNoPWTHym6eWNua5jwUzQjgUY2bJTO5P
tqdnfQ55tnQw2p4rMsmTbNZPSBVrwuu7xlYzdS7MEWsDyM/ovWj1BCXagmRhimUh
luRwgXS+L6Z7vwHc2nImRjVQEGO9CIcD6x70rDBpzwkbBRKqR9BT3m5ufncZIn6Q
5A3kiqsjt+EVUMhBVeCW7hhxS4SA6BrwdPCOsUWRKUVAOboFBZs1mKwhlkvJ0yaI
IvJ45AYOpQ7hdU4LI/VvRr344RDetWvpFU8+dvfn2qmTKrMfQMN/957aoUegUnlP
yXMRk8Tsw+JVpnBrE2jrWScB1Wln23ClSLt407lIMuazgXdFakHsiiRJBjRN6S2R
vSwNAmMXl1GVAAENo571e4uym1vFBwCNXa7rYcMrmnH9xioIXyRXaPyJM1ri2Ilu
KkzBoW9w8VQsTwSRO8SIaAmbXJI4RAxlRm6oFQCHhfJVlkL61PVmJcnz1e6DE+Iv
U/CwwghlKijR8GSu1dGbF16WRppDHLTHPCidIkKzuimmVY2Z+MjX/NyHeIp04STK
JgfzPCY0FeXlHDelH4pbCPL3nZxr04Rg8YBGltL5yGxME1muictS5WxrcpqDuiXP
wuKG1/cRdAtJ0a0z41UuAjXX+QE4OnLXB8YNv7iwtM87/JhgrN9/ikJjeoCbPCkU
fgf3js4c+QugnHxnTEQrzOu4fGrHjhbDz/QFua+2O/ftm9DryGioqib7EbeVRMPk
BLhb4Qx5WHM0ruqSlAf2XVg2qJkWIeoX+SOEx4Q5fW4QhjkKdDovPrW8wqZTDhkY
kZDe08REPoEHKOwin8bsOhWNK3nfZl3BHB4NoLjneTGD22PWxzdxxGFplji7VmcK
/WzbyZKnkg8apjft0s3f+qOFJ8IJedn+3DKFU2uv9B+fvpHDHqxdyOm85sy2pIXD
px3ZH4hsow8yBpyJ88r0iI/pFzaHE5NEtqnun6ZJmJwGhtrooPj3QzX16vtvNOqE
oA8VTRVW8S7KNcuUS6BP+BP976+kkyj4K2zgh3jRLSM4zeKCoBGfXIImT+e+whYF
n42wQEDVAsDRmkbToi5FQnP0iNdjs8kQQA5pexWCVe/6SEj9mrfLZBIytzV6slvi
/l2YnQSJOeK6NzXqKZUW83Dpx3NILQBx/dUlF5znWwY4ihajewIVxMcRNBfBqO6c
kpfmc/yptIEOC+RCRpmdmi6lFwi+BKZnuwBNaSLc8F3HBCx2tBA1W+XDFWA8La5o
oIn5bud0yS4TnHgc6PSP3xsJtbQEMiFdrOAsukhFaDmXH5HCyWy7dsM6FVbu+z9Q
0EYZgIJbg4KwxTmoEiqeJFRI3L+/IxBkRkMcQtxxrkuXK1wkhcVud5yXrJt876rN
UeoRGLgs5gcBEdzRVt6JLTBef9dO/YWkjYR6pfJ974rzsSvE5mLtr+JX6ovXwIU6
MARA4lpECpxyo5qqwmmiHJFswIvADkknx5iMzzg4my2xb0FZ96IcKyLzPkbCeA3s
lVqfAuSeZhOq9fOoQktfKkH2VnI4OyR854r9NDWa2+4xXMoXXZl2MedH4sxmsaCE
jamfyxfraXxe7OGw+RYGaxDc2+qK0hwtCbnWr6OsVir6CVT1ZOx26XnUWLkxQR+x
xWYfczFdxgYonamykEMyVPwTEflHMqhdYjRNDirXkieIuXW7NsKVzLGKYZfVIXYs
ZXjp5WN2iAYV9QnYUoizRz2DrVLyhWiVhNZKhT04tJFQTbq641vbBSxzsyyLaOSp
Vxb+dOcd49Un/H80/+9piKavTGM3Jt9uMiSvwbcDrgaYw11isVgvxUvr5ERtv6pd
Wqp86ZejWpqVm4gp9OF6lJlAMfoF95EqrsYhUJrb4S32A76X0Tw86b9wmKh+LtHj
2gd0DGiz3JP/Hcuv0qaT1kN0TDKGTpCDSR6lnNIFC7Ea7yJxOY9pU2QviI6wfAin
CU3f+rhbnxbKMtV+nIq6jTQs6B8PUpJfwbEVBeiaL/DFdfbgHdSykyxzEFq1sjY2
CGFTBDcPyrP859fTmAED8TrhLJVLFVkTW+La2rMIDr9kNpU5rS4Y8saI4pHOub3Z
uWmTw8G/cYI6LFw5NfSDZ6t5BDACbLM1KhzN7ju2nZoCovIsNfTt7Aq8fseXoHQS
kbVLyddVhixz+cT01I/69fs/HCh1dAWF4X8ThVbQ6/nVKkqBhT2hQg5v+J9+NHG5
4QmPf59jaKytmp9A8l954UaOltH28kIAkgIUqgIuzc9WzT1LnH8cvQuJAsnNWJAa
SSGCW53FYdR8JkqW7Uf5ml7HxgfyVGo7KL3y15QkAWthXoYPbuAzzE5s7akUpuW4
MsM1PzDJTttlVgEe4xgtLZeOy8UGvr635nsimUqJ7QwwJtFsc0PrcBDKD5OE7HOA
zJn4DQuQJvCqi+lIM9cadsrYq/X7Rv8rHucNx7u7vL8kvxX7RCA3yZ2VUJr5Z8Ml
1Ys5ZSE8FF5pUpsxPpAYszq9PMEpWC7Qq0Fut5Mguu64B1XLpQpWXaFP+jXBVC1R
K8LkQAwajn+45dSrfN+++08Tii6gZIUeZ1y9MbBYKrdpe0/ggx0GlTu6lUTwvuuq
iiXhsaTsIVoFxPayYhloCppdfnVDS04eNbgG+JTy1Wwbtw84ZPQseP8VvipyRtst
N/Iu4DYwi3fdxzHwNA7BY4S7g9VjN8ZyTHVldYd7OV6a3/vMvNqo3eE7mCBdD/DK
RTCKAz/2jtGLtd+HOCFZPd+baHV8uxpHhctYhyMbihhqz0oo9n1fN2v1SJaapByG
ud+HZaOLrGuJHE63LOgkc9FQD8Sa0yRhLSpN0EWOK/Bc3UAFHVBYlxuSJTfsB0jy
QPBPsQAP4GhsniFYw+19Bk/v30dxfvCuLEeL15KTARFVa/1Jt8aPeDcEdFqijnaI
RxBCv57ldL7inpBipJLqxUkeWmaFNquiTnpFyj+zZLWUKu5GIqGs4Y8uwlXiJl97
f+t07JTHMHS4+P6SUgMGQoyQCjCewDK66w1gJ8ZgEMiFyUSI01P3eGviK7hEv/xQ
dUXAqYPA3znufqeUfgqME2BLzyNeBLQtOPLCL1bYU0+jbsh+9ZeIsKJnmQrPPZZJ
nTaQhAXSfQC6+JmM/xDGzWOOb+LYMAGdmsC5IEpPjCAgdbCyLJ+JhAPH447dheg+
DbsbUdNtaM+FAMKaRe4PYeamoqaaEP/y4C+Ti5/tb5i0iElcH2SwYYS3nd/aa06s
s8H9g4Gx6q2/dOOVbqvmngxgFJ6XnV0+1a+LIscLZjSAZprVu9ulfVZNzLnnFNkX
MMRWJ17ezeES2+H5+4qsubDoIjL+fAv1iO5bi9jPa5cI8nk/iuLx3iOvCFb447ID
92Hx6yY3oxNwfVWhJP7XO7GPzya5h0eK6FZzwGgIheYzsoV+O6M5MKmbIjgTdxT0
Fd72umZsLD0B19YsRlBrGqd5vcWzPsNt6Aa8JjmKdQ4LBO38+ymoT6mVD0wnfgu2
u6mrnI5IC+SF7hyHbiRfrlyIwc0/X5vEhy+s7W1h8tes70yZoEpjappIgGuhDWXX
xVzzGwf/JdlF/CAPrLNssTFp6wEwxwxfd0dh9b5kZotbfRId2WUNomJuO3ji6RTd
cYu+8FqZ/aWBWVv07aHGx10TeGaPSr+bhsX3UIJZNH3PDciB+EM2iSEEOfBzwBY9
YSJBlJaXf7b/AxQzmOT7Fu2nFIOUNG97RLp+Eb7Ag3kj6Ekb1d+VQQcX7/DRQJoF
RDBH69jArZwNAvC8VOB2Vx7dTXIUA6duZPWHu2FviNNueBBhC8uyUsFQ/9XWu3G7
0bxqgbfdu6qXGwzq63ZdX5DZzChdYvmETIjfNHWc3gTmgBRUZP9GCXNH8PHHRVes
hW/+DrLH4hGQHMGvSn6dQsnE5eW1yBhr4LbqQ2ruRNMa1wpaRJUdmGJv/PbvT/UR
xfXKlcEbJz1GNJpoZB5/k0C0CXHzHOHu7uh4AbdZIxd+Y6aJGgAFET2OPy2A5Pw+
B38AXuzUSCakmREYC5IKeVSPhbyVufIHYDEScZZ3eDUqN/Yvo073TJSKYMNwsueE
nQoYUew2bKKkbtVlzL2UkDTpismKM3eqknLk2gSkbync+2UXSt1TorkUkDxbJphT
J90eLu5SBA9RYiheNTLkXGsIL+JNYy5W04EIIRM27wLr3dWKtPt9e1ZMo74a22q2
Q+UsLa669uDT3CKsae7HB9d8f8/dGTVc2phaZX2C7D8LL2ywpB3eoUPV0zthsbpr
qLzzvDEmkZqMhTQWO6uLG7e7q6DdRRKD2zU4ozD45za8c3x4RJaJXInOsV8eLEDi
5p75u5P3aC+T/dJ/zujB6tEn9G2y/zRYhbGPahpgpiTgrkuIROtiK9oEHQL00N22
23vDzosVYoApLtYOhncx5RnGYQuP/zLhMI11xcsyxXV+9WFKI3+ip5oEtqcL86h3
vs+mZs4iit+uT8nYu73BhVOaNa22OQ+s0T1Dx5YDH4x85YNR/fsXYma2gNi+WkwD
1fFP7GZ/dQTEEoNrGz527w==
`protect END_PROTECTED
