`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
61rCwRKGWObcn4TO3v7X/I+jWk/z53cB0TIw46txFdUJDvlydWGEMR2nS79R6Vm5
315NW7wWx8pFUWyS5bMqHI9JJh6nWy64H5d9FNYdwZI9+RDB3LBHIvqnMfxk5VwX
Jiu7VyHwpAa68UZdjJXSRvS07rDkqhM4Qoy1cJC5ilK74rSw/8yCGjnycPVcNToI
Y95Fg/E9U9c1vjHGKe/r9PZ6INax/Ug3+evKL5dctZMLW9IpjKmX/n+dpsOET77U
h5049WEDyGLcVIRbXEyz3yZ0GYcdedogqMKfbKFpJEUMDc5/PeDSJGmWFL4D3f/D
/0zCLDxogCe/AeDaQjU11CLxRU3j4thkYP46MsE6YCv9mJ+F1VMwlAzzwqQf9bea
ayhnJaQRPbQY9Fo6tB/u3/tWBWgSDUyraJ4KwHvXiuz4Job/Dz2uVejqwd5ND0nR
yXUJZhfcysmSkLbCA/bFJcBnYL7lO0Nvp1co0fQ55Ng=
`protect END_PROTECTED
