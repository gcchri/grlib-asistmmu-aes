`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qmTSY4AhqiOVb7wRetw16hw9JPGuzChDEIHXik73SiN3luJMch8liWmHnzdvgjbH
pcoXHGRYTvM2QABsyy+TZ2GscYF1ZilunMOFVdwc6DAz1plM+3HiYRcFf04jr+ch
MIbJ8GEn7ZlNa6v17O8sXfXvUgQZ7gTH37+mEsjP/pCEOylCD1PRAuzNJi5nK2HJ
f6azyMMMe78v99BGU/8+VD518gotbnFzrnFrB484e010LKtmoDqQRQcLLruNSWdg
RqOKczdpIIjnGB2PlSTJinid3DVBqkXgc+xweP3ll+WS2GQUUY6zuxM+lTsgNoNb
jy7Hw1TVxfjMyy0/7WmsZYmckm6qxQdBMBjBmkGLT/zqgrzDg3yETYv0gyHWOp9c
J9N660zsrPjoIgb+bmINiEB2FA6EKFcLwlnNMQmiWIS804lltKcojepQx8qoxWlz
c+5IgWf777HwzAQhdelhmePMSFwMk03Ylkaxd3Kp/onKPZkjlR3RCYY/P1DvTY60
`protect END_PROTECTED
