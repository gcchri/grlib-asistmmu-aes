`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gbXVxoLrqfaLVWWUB9KKzTN/NTcvSIST0tr1fslANs3ci1aGb98fZ98nP8NUTn6R
Y7frryliePKEDhSKAO4jd8/T/Hlgyq+8BUlDzigGt0dlTlIowFOO6we7LJuFmiyo
Q3VyY5oBYiWLZO9GOYa6wvtoJ7KycbsbUTS2/EJNnA1z9W75FgDUC+jKvA9nkMkm
LG3Q7/jR+wTo4xNRaIZ0Q2X93+NijPEfj8u17Oq7rjuBlvz2jX72i7iBU1pT9n8d
7IY3lo2sd+HCw2UTtkMIRtpQN1QZqTDh61Dw9MRUua7paW0fglIlH0FufFZ6buoM
u+mUgHq9LHqMeJvfGzuMn2QgwY07q+gjBfkG0e38S6RLxpGHG2S7HvMkB34J0q9y
`protect END_PROTECTED
