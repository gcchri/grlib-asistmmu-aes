`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1vcPAkaTqNqhK21AqHI5yvWhQkdC5PrPCA4zhFQah5fFN69XwMoiBWqu6HW2GRhn
VQansgI8UMWMzyLlYayk6Sktk48+35zglLXt/UoVl8L9iPax66QNpiuBI1969bgB
PezTMmtIq01gEPrJHkTTtxcNLbL7FoxvlUQ8LyV/XJkiNW9O+hEW0nCzjOz6VQY3
uH76kA4zgAoUVLxUhJSnzLbSxDB0/zS7lHUr8B5guajGyRtQIO26NwVrPvqiR3R6
LC1JNsH8v4ZTxw1lx+GFTBNRWPkw5tlA+BlTjM4kb+l3U7h+dtEyoF/ouxKDIOtI
unuc5AvqScxCytLySMpwxUjwolkCCQzVi3/sl90teqv7pNF2nApkASbEb2ey/9np
awslgcsR8FLy9kkSPgbrwKtb1+tVF43pJUFMT1iH2t+XrQRSNAUl6JIow1F0kX9s
gxoxbi9cvDxnzadFa5Y1sYNL7JuDSE0/2W6pQRTwWiM=
`protect END_PROTECTED
