`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wh2bVRMH9GIO1XVhsmRfkge37IGVN/OJ5XO7muGKDbzsDeuu1vhtofh3wEar/9YR
Ac5TB7voUarkMW8CDCHJboxVYCp7kRl6c3J/W6fjxSDonaGsFb6Jk730LxqE3G1t
xQhB8sb+52mQe6grKOhDrmKeC6Nh6TtP5IAbYOBHFgk1dsBlCUR6+rkyJfY7i5Um
9a6zIHNNiOlDssHv5n0bRM+nNno4Di+HcRnEEAR+1ZYsgJr5v8/fwjTyh2sIL76S
st91BZoW5IpZRZEqLKYmVRDZ1kWcDJEi20gld7bpjnPn201J2pz2sgj6g7FRaeUn
xRP2M2E/KKWqSXdAurn4cfcbvJ1gBddK6G/dOii6ltI=
`protect END_PROTECTED
