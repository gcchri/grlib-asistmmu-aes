`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ToiP5+h+V8NI6ZRnMp+iw1vXAdHr6HPtXV9SDy5sErs0fsizQ+8DiLxrXtG/2vNk
MCvHcPXe6t6CcgLukRci1NIGkz9ChLDTq2BkRi8Sffq7P8RnQlFDI81TcTV5Q7G7
NM4Cue2AGS1PsXX4Ae5DAIgNU/TH5EMUzuK6eCqOgmFBXZdwRJfmtJjQOg2SZI9t
qZel6f09GF8VvyvVdcDgOov4+xAgmju4y/0tKjscynxE2/X+iinTCBW6dWt+4NzY
z2ceg7kZeDHIzf1/iZM1eSPyThen9Q1LQlIYDrqqChe0xqWcmsHp31Hmm+rTkRdA
z6Z1oR9uR5796AGsO+dIdcRser8dHmVEP1WEv/kSsinsXA60ARgM6VUhthLJot2p
VyUzl7YOpwD94aKmFdLLVH2ByrP9R7wXT8f4osqvyu/IX3o7drta2BNJ0xZTkXUO
`protect END_PROTECTED
