`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WHky5nmizNRcEjTw+3eJr4S0iWrTJmZHs8n4U+BirTw6k8OGHfqt6LgTnVC6o12A
+tIbj6jSkH/PUt2iJ8lIN52o+IOGSRXhMcSUorYTBMRWncp6SJhPxThMCwork6GU
xUreQFnAQx41nMFHlHH88M0Zoy8xJau75+K/727YCljev0GS4d3DmErG8/DjuFKQ
k/zVKcIVJxgA36byiVVhJaiC2EgRgCtYtZhWQAfgbyuBB/+lvbzMWkmMdrB7BOks
GVBFigNY+to1vmvz1QcnQ8xisRcLKu+p6AL0ikPEtxRPJzbECCcUnjfZexG6tr7Q
iI3kHX0alHuFSkwjJKvQth+zAaVThpLicVBm2cNGEf3pZEOc/BE5oxzb1LFLi7Cq
aJJgzZupZhmyx46T8SueHLdy51YENq0lr1z5aM6mGrzmW9++M9sDQKJBAGb2SYuo
5OAkV5pQcEMcpuKJEv/CNX4cMWfdcjCC6cOHmDe8WnAUeGiYRLgMrAstIpJOEkwY
lpO6ROYI3qJSrMh3ROtftPYfZHGaDaC6CMkZnnM4/1APXQdABXdM4WCqCV/ETSrJ
`protect END_PROTECTED
