`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X3K/DaGrPAOzsvykAYp2ecXw3ghJ34m2IXSrmHaBH+Y4GmWeIjpHtVYf+jNUq2ut
8eSN7nXA5GB9/MaasXFU946oZmisB7TKMV6GhDObjYdby4J/V6tdOAEWcX5dxXBL
A+9PsOGVQgZR12zAfYWUc5ncyh1CX7SeBolhY4Hz0OgJH77tTWvH0Ekb6WShn4ik
QjT+iSA8YteQEPLMq5FUx/aWQ7QzHHwzeWpLHdfXr/yXLJzlL8E2dH4gicx5f1Ld
2CBXWREPNPS7QpXJ9vjtJex7z6zlOK+xHaXWBFemNouNJxwz+Wx3ebRlOTLEu5VD
hlzVwa8qjIDfIXD1xVZnddbJGF7+6lrCuh9OxKUTeqP2EgJIF0H3t14VfBERbSei
h0LofJgCZiVmhSXFuuYjfhiTryOsIAeS9hdyqIdwuWQ3SELk2+FWkDUnAqAm6UBE
YlZmgvMZ2In6RFKn7OdEHG8koY7fNSXwwrncSCn/7Oz/mZyN4A9GuPbX0AfnEDBh
ZkmYC988bZmOAkDP8lQ4xlPPOL+kW3+mWV6i/zjN7vBz3L0GILg3W5gdNkOpdu7G
2BuOEtpbdXMzj2pSMay0QbChRbSLzlqZqA4NEQnxxm0xRccrgzDWgzt8+OIKfIgQ
w2+aOSYB9eqIHc/PwgnRWJMQ1yImpZP7CYH+FA5Y+qA=
`protect END_PROTECTED
