`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2V5gpACN5x4DUn2SPx379xM4Ua24IicmTnES+GQNmbax8IGvIdu9H/756a2Crb9T
md1S0BgCwtRzb7atc3FI5806NsKHHInfsdOyYuWYeqp5QheaHlnOhqm7cqDWAE68
a3i9zpg3x+DzTMS8aTM99omQp/VRMK0nRiocBXiJVGyNN49Ce9zfMgnTFLK41/0U
8umLHLwIjgIAs6TaeQ0t2cMVRSgTxva+nG3GxBC5GJ8Ap6giW/yrOtAlZ/K6ID8L
FwwoaDfHon7IWmLVmBd1DV7nNSh144XFSJFoZ90wmtRynFJRhKVlaM+Rit6fgjal
Scp9CmJ/orAJKDSEoaD8aPysMGvn5pScaxlgbff7hm03P63X0mDRSzvA2T8ygxko
+fzdgBFS2O+LlpdmKJ6jjJsk0h7dXSUKwS7tMbxQ5SvXup+uNKeKZzgtvu70UZ1B
Lb5puCmlBOHNgvKbg8jhq6rFvdb1pSuoo4rILJT/8RHHFA/LCrnCL85SE0NFKlR3
L2h7xERl4jDjsZYrc+kfgsN1RXhC0ahS29oBNtoqq8RXCr6wnIRl/GQ61seud0xJ
wt5aIY8fs+OJmPH1BsFn1ufh0D9tcfsOFy3OWtsgMxHSKKbQm4FyzTp2zc3UE/6w
sd39P+H/ZiwMFNJO3+zTozkh82p1S0759n+MtY+DRTo=
`protect END_PROTECTED
