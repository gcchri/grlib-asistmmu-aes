`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cSHzV9aN5+YMMEKA1CT7l+qrv6Mgnd/m5JqKx9B54WAaU9byLbelK/kr7AL51o69
hNc4aT8ki+xAu8Pfp6t8i1jLvGTUStBLHxfizPz9W/+B4L7J7KxDkgGh8+cg2fm+
U+olDxFuOk/PZOtxQ9c6YdQniwGbJHwDqKYt5n9AaPe376M87mp/HtqYqZjXgtcz
Q7Smtvop5ijHp0K4B0tsDAYCVu5RH9Ac0wLvhqKz1HM=
`protect END_PROTECTED
