`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JAvlC+EwC8gufjB+ykHx7sDCXt5E0wUGrpwqfqQMTPqC+zmLr2IHii0/MD2EmUwX
IGRT3n4cGWVgCy9BN7wJY6x+uDS06IeUJ8N/uGVQMLpMt9tBnrmJkrXdm/eVMLD4
hBbEM9dh4yWDQuhe0Pu/WptofZr0kCA5v/xXa3f8CGx2u1Iw+uCe7TE/yik7yC8x
KAtCCvdACbe8CnAge7DjXBXtic4E8Fb6eVR1nxltD2IMiO2m/fz7f5Va8xylYVxf
MCwb2jZrIgAmZbexV01/tw1RuYTNYVgufq+xjMQsU3fd9+plzWoRHQ9A9Ns13AQV
`protect END_PROTECTED
