`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z9z9klZsdcM153gKufmI2/1mxXSzz3cUJnYT7Ez0ZlJPSUfL31Xx19QUChhLsVBi
A8tuswsOLmBt7sA44CjTy7phKhocVIt8tSrZyR4IRljXIFqcnGr7PR0vT3aY2g3m
eefNgGKLsVQk21leXpGzmuTrkY6fLZ/Rgvjpiq7lVdTULR8uXfZmLQIdfaSQXYFK
yv5uos3gRdwL2Pf3BJ6VCEBGXg4juNLEijz0YmJduT1sj8tJKvF68lBf+wP1HXOW
Vn8b6xaeWiTgZ41hlNEhIoNU3957VRPU0DlmTWIjl0Hemi3Oix5YesU2sXgHy5t9
5D3WIT/AzmhytcuHQrQMgjMbi6drcbvdqVf2Kdcxt50BD6CdiBFXNjBk8xOM7lOW
4DGovkKvgyxIlt1asHQCU6IxbB0EBRWVXSXHkEyoZfmQ08cSDub1pVA4fqfU8iPy
32Kp4pTQuq46gTy4uiu0UhcwFOVhqaVvvcFq0lrX0msmE8aXEthcQDn+4fDDj8n/
3dbiHoFTeW/9GwuRAAxR/0CkZT9oJ1jJH1y2h+qVOq48r702Ip/6g2KBeqSfpkEF
j8umc10TscryPq+U0gyqkGMf2U04O3SDvN78J3bhM3cnJ03j+Le8rBbSsPCrYIDC
Of9x127iXFivHohPvk+KhBCdnJ5fAzyuokX5E3WpQI5cP8bPfIK9bqT2fCVKvgUz
k4fpgX04xN6lBEb9NR725caU5r8smb13WjZWhBwQWNzTr6WYae85xXNE6g5pTbEd
rD4abL1Z3IWjgu5Iks3pu08klBKP4+Ex8fw2AwVIAaA9kOAeaXZ9BwMVeG6PvRA+
`protect END_PROTECTED
