`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GPq8I85kkdEb7HXbdGo7nPE+2q7rhZL1Pv/c141odtdbmT3id/hjbe7nvvlSJAE0
vDVLL/iAD7bEEnDSWG5AAv9s3cZdO0gJc48X6IhH7W6iMgeDREoaV3aY6yqZ91Eh
ch9afb6bvwoNZ13OI3MU+GKq8zF1eAfB/IYMqUcltxJzXb01y01H8NdGImW8QlgQ
PxSGh0o2eWGsLEKMd5h03cVExGUYfBfThqIpkoZGIFsNtfUiBlvmi7MNo6SLgAPU
fe8Aa59Z16a3rgZJspVJzbRcE82ZO1LpAjdsy0nf5LZ4o9J3fkUSYyHZCrW+qODT
+Jc03rBXMe2c39DvjEYgnaUaxDpsE/XeqKh7NCLEJjJ2ejTGGh5AUppcwFHkJfQE
C0+I8dCYaQSMq95m5IikOm0UijvekHRAkUHzYIw5Y/MoefSm/FOPbEN7NyVSWtin
N3JP1BNXyzTGxoRoCs6Gpjc0yuaBOFK1rUB7V3iZHqPjKbLZDAShVm/aSosdLPpT
cLT8LRvlZWF2HswxwLZ2vrM4F6N8ctL6tyd/LUaVmV1XZ8uyxaVwEXcTZV6l0Ae0
7Ak7MlixFIaw77NEH/sBlSrbuSA5utg2Q+7NDLinc+BUP4Cnx0DiMSjRGXpm9lGI
OshIKLg8j8VcvaMrudnOBP2CQgyWFbk/cJsxvhnvA9zh38n4aM5GgDC1kgJyzBjt
tu2LNBbk5SIb3e5yjupjqSA8OaURmLB/RClekhWqi4GxT4hNWaf1v3Rm+bAbpsqQ
kvXpbMzGl+nYmQFca2oQ00yqZvYLJzYMFW5V5XXCdvvECNPeS1O3LhR7uOFh0ISC
WKeJovLbRi27Abpe7Fnk3FTLPBT/gPKeDx4G9724dHil+npR4wC29prZp4eMj00U
lBriQTY8JIroJX1q2OE2Br0UwKkj6dncWBShi9AWTvAaGSYOT+VGXxWn1hpoiIdC
pRItJ4s6K1oaOcOJqPEe3MwDIBV6S3WPjsSo9QVnVc63yarSNbk1XdcXyOwcf/qG
TKgGpGoGOxsQ2JnGIdHdMRY6vfonrl+vNwpUhKgMn3hOazge03MExhRM5R+bZOcV
ZdlTwyavj6e6b8OiyYuLQuTG1PMBGaXfEl6t4DHisS9g1l8fc5YNXtEmGGLK7NrD
r2W9u7/x4V8zDQOo2K4dQcrOsaAgsuCiHzU6HqGYUcKoTElJ3c65gBgyq8jlwDzj
PT9QXPs6M4opnSWTXhOgTfHzYdrJRyIXPRYGYjsC4U4Tw7Pas3e1mbK00P0dr54s
tL64r/mzW4wCbnbwtvPPbGAEqFqb+OSiqGIwqpwNoU4a++MC0xs42BAucc5CTRod
xDDOuLmc2QIv1L/r2N95DNS+N16HjK4rGyKEgroPbm8Zv8BCqWjCjFi7qA/Z+dLT
ODa0mcWLMiOgPNaG18FQBqKHfbU8iSQ5i+VsrrMKwStzD727+rqSa8pvbha6mHAl
MIKTAxhnkY4KkA2bTA3UG1zvYp9pgHfH6cQMZzuPHdP8WImyr27dseijKNmR74w4
676CQmYPck/fDpaPzTUifOXY72maKLMktZKuz1BfNIhOGEeJQqukFvpXriz3GTf6
ggHGKU8f1O0loVK68fNLbWg9a0zqLzcmWn7Z7dGrAzgy0F/iQt0o6MD2H9hN4rtK
VAoqUpAIDq3OLDCooim8zJVj+ojMhii3A61v/V5wwjNevSW1CaS7SWZ8GJVkJ5dH
A33Pkgd6LFQw0wglj7iDa5MqkB4gTXK3br9Apx8c9KrJ23eBBFq5V2hlgFweeXVu
6g2/iq/eyAz3VlTpKXAJbFqU0hGwMRyC00NJjU8EGEOMcLIc3WeC2C58sBGMenME
HT+qHjXMWjoCKmuTy/GGdFOvm9W2I9zZwafaoHgIBmiYTX/CjaHNuwQ5TpwOatAi
aIonqkyePM5uJvyql9t5YxZ7sig5AYUzm7YlZOAVjj0zKkP3FDJ7dvw3v0v3oJFV
RKbmAnbKE+ZVbfiMKY7rByK0kKaHd2uYg373P0JGZMz/UFGls8wxWV1sjUmsYmjX
qe2M4iWA20BOIfWmpeK9NzOF/kIiIlYFeTDPKBeGIqJTvrKN0OfMPhtkLnmiAaXe
q2OMTkwZdPxRin/rAWtD8w7irLlGvFpP160gAnxy4cEzFQakvRhck13h4E8nHXsd
LafFgQaO/lKy7CpYbGVAjp//OpUn3BSVaSrHhb9KXS36QY6LV66D5AXnHBXf3c0N
00tHsnMNRWeqYufQiXNcZticpMJL1cOxfpB+IO8J6Jx5CaBROks0K008mlXm0NSH
o59vyGZaGj1+b5C+cwv28WHqdufTY+++XLJH4p39No9EvyoOSCadXBGrqBapu3W+
jbpOCDO5sR6553/1TR2nVWZYurrxzHdnt42aWpqAG2R77i8k2Csf9wXVrF0oM00X
ZvxmDSEttDGNf71QJEzKPlR2+w+sVAR80rV7+JRa+NaVGpMGfpomAOniue7HZRy6
C9B/WvHziA068dE+8PdOjey+3oEKmuXMvhkWvUYniRx6pwM14qpIVnO83s8YHmDC
LHgdrPYd0JphyWjyU8XpljqqIBfwcOcdAK1ZJFWaolmFhGMzmeCdiHOg1YhvK00J
di+wFdAD4GqnRO6lEj80E6MaCOkGJWdQUazAOBors6ddxZFs/1pjj720DrbuASTm
w9+Z++HO1aIaRTTFdylpOaWyNRIRIIylXU7iaUbjGbo4FgRP7w5Xe3jPcb5RyyTY
7lmuo5UjHt4ADOX9pAxG6FN2F9m54Kbkf5LxqGOnWqRjize4+79bUkypwDmkBWIb
kp1ZptK3CGukWKpnURGsZDrJXcZWfuYSxOm/6PfrTSPaJQGAQO2xEzwTh4QM1WOe
Cw8QrbGs+ieEiE7qPHO5IeZ8Hwe69omTNJZaSo3jVy6/6c+RIBbT07bg4rrRpY96
im2d5LxmPjX3znuRtnILQhj4JCxfHrxU3CmDq3OSf1nzhDF4eA7GCrNFxH7FuKtK
vNwuamQ3fBdRs846oZltav/5KyqKCkZXj96b7t7khHJ6u68bIRJIl4Jtbijg51jt
i/PP9g2R4TIpE9w/aj7vlnfdZXzrtbvVpAkII4aopzJS0DsbdcM2wroPlieQ9FLX
KMO+blzjn9yZsALE1ya4DQTsCqrCmyHX8mIzvc5Fuyxy+dgO0UBXgMO7lgfH3/PB
8CJQMV/mgYYuq03+ykgw7GAHF5AuQ5cQ4nFSzdIGZNIkXswH58QJyvmIYaxNaGRa
bPvVdocQ7GVKwDGrAJAqESe2p+mvVogLHcqglwn7MkpuUuYicqS+jmIbgr68R9my
n/Squmwnar9eRy8ZdzoHx3+91ewrPu7M8lSnIQ38KzFXUSrRCvmkispuB9QCZ3So
DAF6vbOnOQS4MAlTfuoAwkVJXO/syHNOjn4FOt760ce10MTJ9mk0xgIuRtrl3v/e
fuJoQYsJW+c47f56hlb4V+dExzN6NAk0Lg4eBAjr4uYFm/O+QV55Qu2GuKNCX7pt
hAu+mG/tx04GdLnYeWwnjiduCNJZdFGosIZ89iVB+8d1iMJ6s+WUbQLJ1KcbPmP9
KgIy/LD/a8r3rTdo/CGI9r+f7jySqufK6ysQCt7oxChYx8wKMsm09MC8FvCoxhCc
QseSTmzeP/ICrHwm/TKPLSx7fMqW0wHnGTR+N3691c7B2T34HOHE49YPhJnZTFMw
Rc+SN5NgXpuTS5uLfH07lhxnZZ8wai5JmlT8B1u8IAUETGZfnorzjQqz2dFYX/yq
D/RdEuhbiqPgrDWo0HPp2Nzc8hzXet+nNC83o7dyEI7LeBhBFfKpDESlRdg8DEQc
j3GjtJlwSndNFYsfFEPCmU9zyBWFtb9lHWYvDTIAvmdS8gqDKGiZqJxEvUxZzWQ5
EnBsA9k9ejTmg0W2h1dzXYFxMQTJ2QlsuSKBrl4rj6WhMrWQXylMaI1O1KqasAvR
uEQP6xB4SgDNv3SPo/O15sUc68N47p2OTKrdChACzEDffvo3KqJwQ/XqivXf/Icn
WFGn14jb3xjM54c/fEoqUQo5G6A5F1H7dGqAldZ13s92+Tk32fHqPEW47JK3u61I
WHD+GXDMTihvMd+EjCjDDMiB8ZIFSod+7sJhtX4W+OK1skLVcx6ZlhpOqkTtjxgG
tR3kNOUtSqYSXubJmAft7nexMMm57PpUNgZ1fx7UYjy3AX6y/lfIJuwz+I85r592
2TP+auJ5+0jBJOzExm92QPfMoP9yr9zDtn4KRKamefETDAndeaNua1WTqXe8QE7B
cFB+b0mdgMN3Rv+/QCndrXkti+gVfIpc4vKlaMf8qvkAa9IIhXT1aUpHxpAYq60t
QGjitIH/tND1Eh2SnLKCNmavL+RZztgnjpV8DmaPh3k90suT8aOO6epHcXDrjll/
WpSjk85UU+SHzndTAPgBG0b5/T78/96Uu06B9WJD+MCFISjAg80lEr6qGUmSP0Az
MsJCiPJwIceQ9c5yI5bJEuiMQhIYKHpa2fdcZY4LgMtpzLD7KYkAoyEsupRKUMuW
xOBYa8qr1O4gSvcZPlJJ6WR6fgCVoXbx+VTEh36RcVgW+Yx3B1JOUNiUKJZU5ggo
Lk6ZDww1PSnM4LBGRLwzKwkpzQ5mSC3sgMH/Jnp9vGO3ZjSyy39AEW8NyXpUcKT3
oPWf2fftUgDV6pbfAQDPIzx06k4b4WTufffDYrRstkeXmaBrv1ohc8C/QcOUwrIY
XSa2DFNUhRVTYHFuclcykLA7fwusBDfRNTo0klEoCTxgHB2GBqNAP5nnTVnW743f
j3/9VetZ0BW3njH9NpYgzx/sv4qjDMhGLyn0g7qwBlReBEiXvs4iBj43MzPkD4g6
4XwIH7X5AgVyCTO5lX2U2+5WttAT0/kfp8Z4anBqcUHXxCI0UFGkpjSRIO666PKy
apT5hotP3rf9wZwb5i2Q8o1HvxHQezriq9nj/VQqrlBkglWfb4Twp/cFw5/eU8gb
tAfK85l8i8F+tUu5652+NrfTXGzXzDphFC21sG/DEuldAeaFbhZZRV+kzXPICgOq
X5LSt2QDlwMNifbLLP7PUqp1S1aDPugLF8JeXuSf5i2omqdiSsbcBq0S52N5gMOy
egyb3io1BLV4peHxbXPz3+EzYzrSCb/sngx5fkMX32NYC626t+Gg+QqAZRn+8qI/
n4RgHSOb8EhvwuClHLNyxrKl8u102tVbowsZyEEn2H/KNxeLlM9L/PqiAbvB5Umg
Vc07L1n1ZDspHFjJlP276tCm2aWJ60cCvwTjS3VI4a27GqrqkHAhN5Df+y7uikPk
UITszErsxdoAw9YMX57YRhSx8DE8DuwZTyHvJxpMNvkIdGkPRHc1czfK0BX/7LF7
M2UOYfYYq/Vd+LNvapT55Y3X4XFJircCGwYSZYnmn5nOZJyRZax+GX/JWP6UISkV
1fa3pEFmILNFFiFeyCds8JBOqPX4/IPQZCFSdK/dKlJnOjwKmoo6xOGBH27qJgiH
6pfo97FRji5nJMZq+UXfi/OEt10LmYVZCs1z/vxNQDmZ4LGdv9gPxFAMXH10p/cg
5cdQLxIB1njTLZFkzTOgFaoF3FM9RcUxhJJQRcUysNpcyQ3KGbY5GoX+2Zg0G5MU
w/SGdusA+lkxUpb32UO/QEdj1x2jRMrVJEBx8Jy9ipDeEfC5Z7EysoTG82R6fbBK
1p+pxppqyYyC86fFiL3OXOj1XDgfBpyUghmKUKbBYxUHHGcU2SKe3qAxh4MjLgws
9wiPyFWp75KwPbCcZnnxbOJI5RNbdIqB53AIish79d2tdeaIUIep80+p4y4EZjR1
ckdyZDDk/OoGg5WBrDVA7SANwkDtZ/83hfk/hRZ3pt7flrFVLMcahhYWcqpoaE76
le9NSNHuKKy/GFDTQGXMCb4yRkao2Ch7Y9n7oiHHwgXe9vocqbBT30G8sFoMXYjP
cRXbF5BtPjlET16a8TJVwFNPgOhkPhWZix7ZyoViGBWQLtrX0xeymPvHo2WAtfSh
Zgoi7hw1maxM7t7wZofgSDxmua+ewfmWx/APxbJhGb+bYvuA7DGu4vdpvylRCiQK
3iuiCL4wSDwvJWi97CVCScACnKAFu+e22kNeYKX5kcmNoLOGWyjjv7ErqblejRrC
gNyjeHKmh8Av3EDMhXOHDWV5UPOjOU6g1r05qdFsiXMm1fS5a8ap8JOOYa80PPJd
rzM6j5Z8mY7sk3xZoWB7F2yNDvsMNsplIoM5dGyFvDe4fE0oh4GgotA8q/mzRHsW
4Tej9jvrJEeFktiXo/xyuy4/HR2OGub0evkGa99c2YNgr0mMQSNYdCBVPJs7Pied
97xBWYipySYKbZplbhjjw+Ap/XT2IXKusbEnwMZBIXXc9LSGTLKPmGY0TGoNqlH4
B7PP7aujEGLddOz1eZ0q9VQvHG1n+s1uX3SWR5qdCRA2XAARKPgT2TwbcqKQzYsn
cfDbMipnuJq2EKh0uQ0+6Sce63aogwjWQ/Yr8sHsGCN/RaCmjr4YKhSWbUxE6jRx
q/1aQ2IK6o8Hu3rwTtOiUFhaoINYQyk1L0v7HERQF3FSGdBlqhP/OI/ZYzmhObEP
aRPqPtYdLOwVtB2Wc/HsOPV/mv9ip4OHnhF7+YCcgbU3hR3KpF7LICjxKrbHonJQ
Z2sllPlkRqd8H8SpgN7hcxxe8X0ZFqjCx0LNdilLQLopGRbJIHni6gqP3EldQ5rF
Qh5k63g749mxwQeM+PaDz3fQZfUrIDXjmpP04AY2GyfsQI+SKUlgEhBmvVD6V9y+
OiTNBSA8VlIX1zVCzsekLOZdXXQE+NfPX65ucPwmHDrF2aCzf3XLITTZ+Z1XKU2v
0e3ewG+IBckNLMe300Szj4bvJ0yaPTeNX96K0aJrPBTpUV96DauQ3CLDqdKCTN9F
qVTG7hsaeF8jVsLVF08QPqjsVoyP+BCq6Je8+nStl5o43VHIQ5o1gVEhWL9PY5JB
d5daSq7oRzUSrEkX2Q46R9HMiPIhd/4ipxrUVAOWqfcSNzAM1fD01aY18zRL54UO
RIXugtvdo5HpqtUtwq01QpBGgOUj7St8x5iHjmLt0+X7k8ftZY9FcNZKpY3QQCsz
L2dmjqudIvTNspxM5CCKxxzd5Uw6BT3dtPqgOpXPtLpoz7VO/OAYSlK/+KONHVU0
FZqZKUNkbdGHlNYMtZEoq0yxT85R+TC/ueQyT0Or3NySe5Y+VO9PEcHBv75D00yJ
JNvPDzmY8Xg2Bo9z9DxMks8K6MxJ9eV7x/7pyC5YmbX3/weFh6C5yUxXzbrr3ZB+
K5DsQSpbzt8xGWfHBS2XEuOiWMuxy/AAFm3k4f/9taf8DNYZz12rCFTQGlVrQRYf
9hoBzkbh4dbXPON22OYg4ZXnPtQ4WpMrDEG71BGWSlJ1afgkr7W2OFAnmJN6F2Oc
9nFe6n8cGjr/gQxrk1ZI2R2elTA69jpqehv5j8zREozccJazq30ECAHu25hlMVmA
pVAg2cK15JI9ACXV0bvxwDKTxYbQ7rpUsJGIZhwsZYRCi1UVDTHqJ5ngsYuDnsrV
g1iS4DDrcSX6UnhXAAGLmH76fktasDuJLFSbngP/b7R8N3u09OY7f14B0baa4T4K
tDrFgTd84RpUpDSxhTgbhisVt5+JmhoDlEND9/yk/UAt8G/CeW8wM1M0W82I0AZ3
SbTEdQAOVAkbyS6gUcAhzh7PUKJJC9Xoztj+CvYAKAoEejHQJxvCflmtr4ppD3wP
vIz7JCeM/PQNjG6tffKEXLBgkqtJqQxErGcIdvpfINSoFDAznhaDZvXuHMkmU05L
QAhWk4Wo7ejGIC5n29V1u/0YTgohxjXORa+9rswSSryCibUhsIGG6k2DGun2l3xp
yJBoOwv6c48F4LDPSjIwbgoyxu3cEN9RRQmZ7LvMeDm/2mOyaP0RDgKXxu1/csKf
+D1YrDwEu7lR47YqFI76QD15X4iCu4UgDBYMI2NK1UXiOWr2zzJdqxc/maAgKX1w
DSdF17oC6AG//00OQJ5c6LkzVVCuENJZSbMalIIX3iEWzGtiFsGCeFkjdIvwQEWt
g4vn7XRWnpcl/Hc4+7VuG3AVcDKgPAdSa0MYCEZO228PQovNIHaVpwQT5NEgHJyi
VtDc5aRo3+6pRpn8p6Mhq8OSz73bc6LHsTE//6FpqCxxNNJMYBxcm4Cs21V4YSNr
kNpP9SxYLfZGni0akwZxIAbUE1UQvz1AmHBSW0hA1gS49s6+GnlRftIlsBLwJ0Ff
KkZwtVl7hnTW+irv1ZAYSJ6xS+TY1jl210e7cUV/g1+FZRSveb6SupvrmJN9NIFz
wpEAbhSssQkA9CyTSwGZXxZr8biT9yISQxvxDzGpBn7ULwSimK3cTQLj+fUPn1Ha
jzaeTeSuZoLRb3LZ0PLv721LsYAi6iyYftxFXbExFxoyovJ43Yq2vL0edNWdlk+0
nCcdPL2PHBiBPk555klr4INvxUlZdryFLaQw4iAzLuxmyP5kdmlsKf9fpW89wGqp
`protect END_PROTECTED
