`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Bq88s9HNTt5MB34kY5hXg0f5PZ4iW8q5vYAfSdIeqbJoOve1GElp5q5Gn7LWTsV
SfRwooQsA1rIzCgpZcNoEHy+qhK0hA4xvXNj6wuOL2aVsV7/Pq/bsdDVKjkgHKKZ
CcOSJqbTkEKEMG7zq5gNdKvnyxBvqZC2lnVqMxTC6hYm2o4hAVhpdANsap/fHU3l
b0kp1w5ynqCHZlPshQKdbw13TH8NqfJTAHEYzjBiJM/QysGVvU+D8a2ksTnnLF60
yUp7NOMB0NvvnC/G7iX5VIYrYM0kiPcY/jFkJTH1LIy11GGnI9IH9izk3Rkrvt73
`protect END_PROTECTED
