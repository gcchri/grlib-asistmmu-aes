`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V1RInC20qzqPfkppSLF90NdzkYJPDB79k5IP/ANL8q8PO8Q+7Nj0s5Uy/n/g+pDX
gQ2+HpzE8jnqSlmAjow0tsKOzoMWCzxpQSoQ3g9YzrV+0vjyVNh0566H8J8h0rzy
23Mzm1LYkVPQlZjhE1Ywpym/PY0HEV1SKkorAM0zS9ovIeIV/yVW0pmXY8Kt7TWK
d6Bg0I+guMwtH722HBR3nsfJ52Ih/JKW6x7KfgOqHsh5naCx1RqUPbSbQaC2qmnD
m8Cvzuj0UjFmga1Tq6mj/SpS9c073Q4Knp+bQ69jhLlmfq22ZCHyCMXetEYRBZpo
TtLj7nhF24/KzFiNmu+KZ5wJkqHnWUV0I3XaqX0SIWipPqJvRyxKMpprGWyL2SGR
3OtOXu8Q1xjSu1YfD+FwfBU4IbG7ljAYiynoJzOUp2N7H0YhIBhp4m36+dsbDt24
KoBiDrI22KpUcH0pZjNLk8UhSNyAqcUxealVVaL9eJ8YXMLsXl36LxIk6amSiiLf
QchKB4UTwqSlf2wwaB23KEVlCEGhVq2jBvO3NNuwu6tLKjPGhewYZj942jwh8F37
Z7jZc0+/0Yiw4T4s4PUfPpYDvdo8vBNunerjUnGAEV6Ce3CfxenO5of6xGPwUK9Y
kDMnx2sXTe65yAlebT5jqNlgZP8nVXH6vyk1tJWhzd1twGwgzSYTJ5u/1cSDBm6t
n3bW0m+a7LN5iZw6z7El/GdN1Ho3b8Ju1h5icCryx6dueJMpvnex1TiwWfBlaYH+
18vWsV3uHQty0eKoBjT7MlpK9UzAO84GFud3v6sljDtW4JjnM799PbOg5h5AY+9V
rNvaz4yR3wGcBp7EiwNVA2ErpkQrERurdqE/bxCIZIqTDYFT3BeT/wBY3wEHsYRO
Tjue5obQ9crvE1gyA9PmgZMNEisUJIdg5J3H8MI+tMlK++kMGxsMs0DjGGcw/+VG
XJMwLUSknCtUQWAwoOX2c3VJG5Aa+BRZqu7VBQYGMiPQf9GV1Vu7u86vbQxZL2wU
pXIwsgU4+FBaLKAZJJQiEQaKhK5jVksQIZ6qK72+0/i81rRN9iwteuj7VBWv2Nz6
551pa+WQP1K7YD6/4a61hW3txO5EftsoOlVV7SL903jQVbFvej21vzNUYYmAVbdI
kAA/pNhoEh3qBqVV3Urkhyg7xqFfSup46ZSWroD61VrwwP6KM5Jom6xZke0GZgkl
R67gubGyhwtOQP/Xf64lCmuElc//AZerkpOUXrqtF8xJU20eTWVhZsmo0X/es0gH
jKeIKhkF+fvJlh1qN3REbyjsLuYUgv25SgY4EO3DuaGHULoNPx9Dpa3BNWJVaZaM
8QhDOzpdNwEXncOqEJAkSSO02aZAM3THd3MB87LWoUQHV1AA1KweufJ/dO+hd2k5
alET5Gf/ezGf5YurCsA/NuRLDck5RIwhTXpmmkT77zdxs3uvPXVwNcCdiNw7Dmu/
1RNcoRVtfNE2Oi77z1MWXLu7euK5dNiSSpmDuOCnlx3jtEr5EA9EGFkhsRD0/hZc
FsjTYQ88nLD6zC41WveJ70B/kY7VY8Y+0fhL8jhENtL/ATV7draFzIyDTcHSD33G
yXFjx7YhiqeKnxzsdDDQeKqNu9+HBUXsOSdA2ZOhJTXs0j/7ZJm/DEXZkdWf6wqO
Xa0Q/UpHgXrwnM98WM26GSnZPfSb1ipRCGNIOLEuTM6eWr8owEYMPK2oQU0Vp8qi
5GxWrX67fzpO9+Pbw5yr2Rmyy1UowcZpwDBbqG0C+Bp60fF7pPsnwjC+rYsg52Wn
n7+XCnNM+TROyA7Kqmia9AEirNpTbIPTlx2hML43PU2Xw2GCH7PGK/kFS7RCjx8s
AYdMbM+x7NDjsbietFXP+mgTGnKxVw3DmhuA/UfgQZOkZnBnXiVoDw35hEA0bF24
z0tMXL+b3FVlB4z94b/5r3S8PnMhMfmiqALkSFtXiNGNbr9ihAiC4deV4awYYNth
jibIpdpBsLcyTHlxBcU0EZJ/scqUrnoee748Pjrt2gRFe9Km3auH949eazFWYyfA
WTx3WLtzleYi2fWQX1VeOyhkV/2hpfrRvovLvNRmhtfG9f+TFslaLF6XT2wdbVAq
qtbQpf5HQKJiOMRgVEfAHDLgEz+BW19LR/TH/fK9XNw5NbJX/ytjZI7Rj09Q8QNu
1O2EEaWaINrsUv4VDxwX6T9utxhDUAAM5LxWQBXLYjn/wuxNUoIdHg0TNl80U9GE
eIKuYtnpGqp1D+Fnq7ddPRntk7VAcYcJqJvlzpTkNMIiE2ZGYorldeQrn5NxgOwy
I2DH2X8STITuZTNByhmDa/Qvtb1QTaGG1J93TBCQAik=
`protect END_PROTECTED
