`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZQrDSPUGtp4JorbfxGHxdOcEP1Jdvzha3JvAiMGd+ibWexUU1m3iEBMOuv/nVlGC
q0CsPUzMIGEZ5KypgM5DiMADnhUVKCNU0FLP4MYOg27blGI90r7uxRg2i4VCTegE
sTx3DkKm56FQYu6YYgDNVIRTtMKFPJ31VjzHUyBDgXoz+cyTs5Me0wj6uExQ8iIr
MpkvcQOt3PSoWSsP2LLkThVHFcqrG4lirWkvl6g/ByaQY9xhyYvZJhGT3r2hv2y1
1QYESWx7tO4biVIycDquFyhrDUmwB7YNOR2lTAeAO3oHGRl+SkbBOgh9UnaUKgiv
pIpBkJDx/o7Em2HOUApmEepvtvFij4s+0ybUOMZsrmWvgwyM3jjiRzumO1vP7VQG
VolM4fyyY4tkXyrBZsiY95PyzxB+CNJjxn3u/0AlNIkhKSC3G7+PH/2j8iSkk8Ia
lCcLOQ5B5VkWo5wEQa1nd3zlwn3ZzyhQ/j/XpkHgGfqSjd0zfCGeYrnPoV1NYl3p
LDw82fM7c/t8Ke9kghFajQ63Ga+2f479WaSp8dqYEms2iWy2gSAofbNj4rnqg9Uq
ePxUvPW1yymCdtKLnV6p2wXCEYxemzHhs+97i/nZPYA=
`protect END_PROTECTED
