`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vry0G5V1AzuH5N/uDcRzu7mltJCqIY9VXGklMGvhFnz/l6YMB3ZZnfllU4W+b33L
pV/gF/a42SBBKDw7LYxapUSHMLbPtSA+Q3Fy6BQM68TEraBd2eqrNQ4deTsUWsS0
DtpsDKLA25BHH4+2VBtcKz3HB/quLcaMk+QZlTZYl2SYOuAw3c0uQ7n45JZVC7JW
eQwGFwL5a5jzBngcgGUDku323/tO+5b/QEzth7NPHNlU01he3p3dBkx5JDAxwiQA
EOUQWP/XlbvGybK9LIAm1O0LpcI8folxX36JEHBOhLHmT7nj2AdyB2ayBJ6ouKZC
kBZPhWI2FN+8XyLkzm7JdEGpPqeUvkVdH/FEE9/+XDPrb7fUcUnBpri7r6lTvG7F
gNkyy+z1DF+2p3pI5wMBYHNCI0Bn3oVuAkoNDiJO+tezFjVnc01yzBUCga6AzAct
QdBXmRUcErK09ZpHvKs/TsJL7pA46JAkb9hW2WGucilcp4jvSepxv3ITYKjlsmoi
`protect END_PROTECTED
