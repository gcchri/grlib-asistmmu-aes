`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g+3PYlPOUimUxg+4kLI+LjYsxm3UkoZTBoBlRGT0ZYdccawrmIxl0gAVIPusXHZB
REx+rnkI1a1oVqXqr31Dzf/D5THsGHv7zRDGMWfkBPbsm5PtjlSia9YfNwXs+sDD
Q6U9cvVzEVgR9pfHGBsHRLaEt1vvvVPbcq3xtv2h6INvxiUywULiB9lDyfb2EZSo
sAnfAMNnYbyIB85QClZdkt2LZ6FlZQ9Tmuw+VIHmSszPJX26EGr5LI3r/SNP1V1r
3XznshzSM4BpJw9Hl0SOf1pugGwnolU+jG5cKvLpTVxX0nrs+rw1rFaAeYJKhV+D
zyKXzZvex89HtaLTc4igBWcEYm2YvucSv0HJ02Qucf8TssRvNDrnxuM+314nSKRw
6yoGCgXpCu0XTp1uLbW0m2f4wCRK1QxdJ2L2zKm9gvTOwUh4MbEF9PAMHZS/+Qoc
jwmt6SlQy4zl6qq/2kT5GzJNIpm3CCzZiyNVoyRPsmQ8czsDMIEjU9zg/b3Squmg
DlvMFjheze0A9SN0R5R39NwZB3UHBQwy8LUUevf1Kzqk7CYXXBagaFf+YzKX3AU7
yZ0dz65VOL94lOzcE0ZH+mWtUHMIluJTljLFDRci/x3+L1SFlz91sndEW5A147Po
W7AehB/BnFHhsLYLmY6cSqSxKdcsGPgOn1hZEZxIvGjNIGv2iHNmXALfGgI42p83
Q9G4lppXEePt8sHFLeUmi2/WPHuBqvT6FTPcvROWzgk=
`protect END_PROTECTED
