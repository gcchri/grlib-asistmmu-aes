`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C3y9xPNHCaTPCEa+ZYUd7nM0suIrUg4YqvjLVFXS31n6z6WGFEsU3x6PCa31Y8U8
7usjAvZgwJPKwCTe0hby4TdK6inc2E4zqL/Os8ngdhRMOiO2BDouMYDZ4+ClM8ey
BXy51Qw8tL/txyu6PX2OQoqg0I2+GVWRnHfV8O8AKSXmetHk798rESM5dLQT2cBc
Wre7EmWh/qGB+zxnkL8bxgzwTlQZnUajChTsCZaR2oS9tdMLtEYbQOp+lwmEpmD/
wEsoWdT2d1KWjyVCIX6S6PXw/E+6j/MvB+AvxjKOtjY=
`protect END_PROTECTED
