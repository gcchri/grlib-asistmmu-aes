`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K0cUlFUIxKoAUrdQ7XmLqPSvcKtlJCKW2qXVv+7R76iauUN59qnkY8uQuaVWdd7N
RwgurMlkdUaxl+DYJPFl+SWgaDdph5rs4HtnIA6nxfpslnWvUc8VCewkgNPtkarl
UQWgvmTrlQki9GOcg28r+oYrsCOv6Y5n5Viq+OuOBOsPFxb3omzfpy+RS2lTXjLS
YwgHxzVkPZ5uE9RbHdKWqhdUJQ8bxhU9sHtwNov24N3hZa4qjrDEeHzrvG1nfByg
TGopTSjPvECqDjABJmmByiyIOvWuPZpyZV2aTSPAhC8uhOdcBDL2BzNCmN7oXSZ0
`protect END_PROTECTED
