`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a8Wpg13ng8neMNvvaPyr2k6ieii2MVR1ZCGMM8/8dipMnXXfS+V/XDSlV+UqJZm5
0LWSiMNQWZKHi/uzm3c82kVkC1GTjyJ0aIkmagsZUfuV1gfsRjq78sAtNNctkvCx
vHtGnUCcw+dDzAau0qRvrsZbTCWJJxH0sy1kxJpUFI+HuMKekSMIfjYjxXWAXONi
9Vmfwlqwz/jrzN8aYg4YS7V7ESk+6flI8wtVx6l8LFNhSB37t1CkG0ElpI4kt5hd
2+n7Iy/hnWrcHYkjUhRNYy4ECzGgcXJreTB8pxSBuwX1TQpKuDESeFwXsAuyPYxx
JfFSZVy49b+DS5Yf98PZq1regxqUUS8wwUyzj916W11JOqLcd6nYcr+Z2AaJ0Yf2
HmHLmyL2M0+TDHdHsmNww8Pif1952wfYfn8LicRCqysO+VwvKZHaA+f5leaRxluj
KsD/lx1LJ9U4HAZ/q32E2tjDwHxkvvBrCCl2insIFH9vIs3UdLgabFIjhRE4AJue
3UIY6Se47n8FuSD8ALN38vUNDfXv074CE8APCNTt9E5edFCQvZtSY6R2l6xbsXN5
DHGuprgFjBrHUtCHu+2Hsr0soYZ0FhaT0b+mKhNadsB9Tj+UFbBTqsTG7+l7W9g2
18SAR6yw6ccB2QKFh43DXhPty/TrCKP/2LdWfJ0GPnI=
`protect END_PROTECTED
