`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RI9ka/oZ8pd9PykKAbPE2VZZU4fj9WkVtDpO+qxEaTUGq8jcW8MH1AxuLEsSUDam
mZjNa5G7iNgttB7P9XMSVG39A7SFnr4nyHjnxX/KcIcEOArRY4AtxsXa8tlnw+0S
qWMu65Gpa5lsF1BtHH59VvcGZMyxo1cjpxmojekZB4yG379XaD8WSt18DGOwP8gc
BFuubbUh/4hdk1754pJKXE1BXPyMDz7q6T36ziENXroG28f07GuvBwCcODjjJWuf
i3C1bRHvVWnImM7qg+MHGTXXu4hxa3xMM4ZamToobOmqEUevSa15hpHgjyEXO/Ou
bPaoxSRXcOP5YM2ps3i9jAKoLYT3bIu++VcWqPgRHHf3/Tx7cRPrDaen4SmGN/md
gi67BjEJmJ5+t0RFzAb4idc2KCDsEhMW5tBASyjycIdlrjgiMNGNAQpFfY4OEbH/
FLia84mZZAP0mvENlxUq1tL8Wvzao6VlSvqsTmMuzhJdLtnRyFmTKrT8N8E83r7/
bOhkgTe4vCKMV75KpUpBb8ap7zI+10jtcAqkxPie86NIn3nzOdO//cQE5CgA0ML0
PIiF191cDYQUz3/8LVdmaDXoPdHkxhxbd11X7XQvRokk1aP09zdRnTiP+HtTfETI
GimP93CTo3lDO49SQZmRYtAjDlngwbvSiBKJoXy071wj0Ta3Sz6hN42gngN+4igo
cfeBjo7191ejb6TtTsZriNJgPz7qPJU/j2MvNwi35nGI202yc8E6ky+SbNZLUb4I
R8TPdNKJjfkGDZw/PBWpxy57ht5JsxBnR5Yb4sc+RwLGfAO4Fnj2DwvufizoyAgM
t/qu0tMYIF+nxxpR6zgGMtKfmcGeGHsgTsFoJwmX05NuGTZvQ/cCO4FwBFW1umC9
MWxzezGbLWv38F7zgW8s1YUki6S3Fv+0TfMsXSzeviqiS4506TQkYAkIPG/PoTwD
y7ntAVbkm/OikyR6s2io9svv2Ut2pGPz3ogBfVp5Cb8IrAnwL76EnuGhHbxJhKAr
TcHSVu5qPIlNozQwRm1qyGVHavOkg3Vt/8kf23zh/S9NXiQxxYOoDez2KZQqV7GW
DTMaZleN6GQN/54BaeesWOaXZ8OQFr0PT9Ow3RhDbqHA5g8KJAF4oc+HM9K3JGgo
dFkLjm+m2aptPohXnOEu6krJCcmpUHYhdxfh7tSYuYuP54ZROlBkyGIImn9wJHTv
tvWMv1+/FF9eRxLa9SVdV3TKGh7ivQ+AHe8SUk9aXyEf/UDVXh9EacVznD0Iek7t
cKtUSGZzyNU+kx/7eiF9tZcYXYG31/DPWLJLsm2x3BC1BXUnqM/7Ugtjy+pZGqW1
rRa6mPu/GWnMalTJsfBK3AVc2g99zDkX25CLFON5s5qpT7/8GZ4FLaj7uh3u1LeB
8+wjZCBEDtfO1Bxe4hiArmUVkCQyKWbzxPZgJVb4X6y1UwdTIy3FYImEve1W5Aah
tQbRcr12IaPEp8hMqywEvzMXHpXX9B3XqzuLRISFVmbAsAJSYA8nhyOI4VBIZa09
jUrnaMzZJJqI7xMqVqXUd78Mh08X5t7hX+a4Ik4crNSZfvC40vE/LDT5LaInSTQf
oC+Nt6mPJbu3CqdIcp5GNlvdroRoianLfCGvnkCwhEciIdBNmCgQKPkbFtdYkPj0
2vSr69Yd+eBvjfVWmnlvXPehXTucerFJeX6qbPDZpWhYZeX738Mix0Ox7zfcln9u
LTvOS6zTbuaoR1EgxtMG/cRPom61U+WpvS1t67qpKH1oc+wcmO0MHYF7h/DyjgsA
HtsWfY5SNHagh8/EsKDg7LHCVCqH7I4uuib5krjvQNHbPz32Bb4CAfMaI8BSWogS
A7hE7x6Drly2RHtuYmDkIvl4ifAQLV0lzeDEFHkaOXV459r/5OP3N8iK8ZdOCnUq
4pCh8dMmHmgvF1nJQ0ApzU7NiflJZ3G7wZmNCuaBKU56qhSFfHdpEMoaepCQdosq
S+Z5k3Or8cV07SUUNO2PUHVTHyn/+Ceb7BTrQrHmyuanJuYkSdf5aOryqRsxQMIi
dmcmK1MjOMAnRVJQZyISKw7wEzIOlNgA0YrJvAGinarSTLTLV1XrIcViSayH4YnX
e2CNGf8HoB3xeW2WKt1dTt8fqBAQiTMONI4t+6J7RyW3RUba77PUXWYwa/gELLJR
70wMbYtnz4eOhk5wF9hQNM4YQmsbGitvwf382RI4mNUMM+GFxyfVSAsB1uYGOa7y
vdN9L5ihXV6CMIY+cI9EcGcXhBLkse2TwQgE8kSZEcHUc78Rn9CjOiLwOW6rB8AW
xXl27XMoYIcTGhb4qravWMc51rDDNXKWbhs9mcM97MM3jxr3SHjEA3IQloJkn5Cj
hIxHgM+pPtzWRYsg30qx+Jpx0Xax6EztcBkmw3JRqBQ35jLCbqP7UUIdVUxnpYZQ
DfvJA7q8NR9lju+DEDxa2s9j2cCiwsgveyAI4ZjcfGIVgj32pAaFOStgALjPEdkn
/oltARKpSusinO/BR0tL8n4KIw+netubFCLyDVZXC1WFt8IY4YwfbFMD5rpMvo0X
CsKquDmNKwxSGuy6XPAxJkeRgMnqCYB6yhQMuaTZYHMPjXCu/YvaSty/0Yogl8Hm
19g6210+2OjKeeqNBAyv9KJSQHr4aPGCkzkonEmj13WLy+MOVeat3mWRaJu9KoqZ
`protect END_PROTECTED
