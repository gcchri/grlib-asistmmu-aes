`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L57VMhXiQrT6ZuzpkAx7JqwLUikWZzaTLmE+3II0aWNO4X96TU4q3nYwbqXW+F9w
OVXFvbnLnTIAl6Dg3rJV6SERXhNEaCKBB6OIltnS9B4ZKJ19vHdr5x1ZYJ5dqWNZ
ZbhKHQKVFUwTdeaa2qd73i7isffvtz87krwKCk7TTnQ/WR/zFY1gLvsKQDquftqb
x41qmo8GK/aKZUHF6rBEdzYUAtd1FVRCyWzpkw3iEoNZ/ClcQKeOO+D9UeNRXfNb
T1xK2lg1yhxMNUYoNcQ+pBML+Xwat1IeoWnJzf9uCK9ic74T4wJ4jN46LWLXxi7d
WIkDoWIjJPA1gqv7Tpdm+Enf6viEIjrPz75BMsLhRa6K7ASWEzYf6G+o7AZv3gnx
4rDGiRka3n7CQ65TVophQQ4+TThvFKkdycgBmH6g0asVgJPe2IkpWG74mCvYpDbO
7tOuxjGrzvPW3Cr6qOJXUFRlFq91EiEArjXZ5Kdh8sLj1cJZrUkgqPZAnlibBUoU
`protect END_PROTECTED
