`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0EXauFe7UN8iNzfHmKHM3sssVzCSCksIc4H/FJLCW+J7Bq/K2JDQ3yjPK+7CXVVz
1H3hFDA4x+dxsq4Fm+ZAKguLmw15DROefe/FC2WLfE+779I/uiTZd5MGmAg5CFBu
pvBnhiuypf8oMj7iLJpLWTMsPAf2D8Zyg7mYpI+bb2xuH+qT/NS35+mTNyLhidla
cy6xSMerFbIhcqr+9tTI+W4hlRLT/ljA1vyye+YnhxP3QClQ0jyhu+5IxOnbMIxg
O/3FpV/RM7yIJzXTIdMNxR3zzn6WByP036X9bjrfJ9CBj4zKc92zATJEM+4bhswm
qsgAPqaJlgWMNRmCic3mSCI/dGsTNw/RfQlC4ImadrJ/q95SZ1YeKCE/YCxFc8bV
jEfTVGr8YhkKxIxlXyEQPoVRbfyLeeuSjoQJCGAd9zMZNrEdsGYGMnhBxUD9XFuR
8L1LdcnHXWo0WjKcKpLzat0jJHQCJebsxDPT6+2CTZQnoSECzjCht5JheRIYi3Ix
oqC36hAfK4Mr6b/AaMHZR+UJEnhQ4AF2LiT8Q3kPFzItGMgw1XCbKPcY7AyA/HEK
wQS5d+D6wxpvZgMTIvr1d2iZ+bfxyXggcn3lOaY2p7EF6Pg23P+/VZ/gAer4WzVx
SUe8ZJmL+VeEXOdjs1P541o58xPPgQCTbuZOyy71p0FpGXP4Je0Jyx4Yu4mUCLQj
iI5JetPXIl1eqZCU8E/KQsexpzKwmrRvHlNlVe6zT3Y=
`protect END_PROTECTED
