`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mRr6vyIt99zZhVqq1w3vb9L67i0x61PAGZMKoFo/gB1IlAdiYwVN5TLnO6u+kzfk
WtdR7WzU3/5Eir4q8/mQKx6c+wJNaWJ6dkczZ7udqrQmdtrJm7rkcrpdx+CzKVvq
brpmIs/p6iF1z6Mom0clwvqZSMt1/TMwyMAZVsJxMHhQp24k1XPpa7m+HKSz3LS3
7/PHHWwOybZ5QfReJkz8v4QjaiBJye4qoxwaiKCEzGs9v62hwSyYhBX9kl6yH1YO
PM3dO96ezn+wtdYzeBpUAZ8ghZHBz2y13hkEWfwn+Nk=
`protect END_PROTECTED
