`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6xgP0/pMLbNHb8LDnLmFYqNQ4N9zy804/qmZbUXnSDIN3EAres5oVqEoTd4cymGz
HR9F4mxiVM4HFAPQhB05JzLTEJtEnfPbORhJEDuSVu10bRuilIrqDhjNh+Kv1l8b
gEAG83mIJnxumCkKvX60WWUJ7Uyu0PoPByig88nPPgQoV+w68a3r9oT/3p/tH+iG
GHckISFi9sBXPcAPoiy3D1J7yiObPwMhIARPnnZuOmSQ8VFe1gVs1uv+92dk1DMU
HM84mHyr1ReVzCUzynjlUq7v0Cg+0PTa8lgfjlNwbl804CI/bGAcrXlcIVSk24+y
7UeUB6x7cps1wBXXp5y6qsTGgxuuj6VJxCda1raynrdbmis+WBS+XRCrYaJs1mkB
zjviq8m9EYzHfe66jBVd/Mn9WtDya1WL4RA73dIzvPkbKyVTYvcmUr+z6cgvLHCs
/ybxJ4Fj3FxYNvt5upAquePw3WwerCACSb4oCevJyr1xm+Ljf7p8GdLuK8OzQ8AY
oSxGOXZbXXGvynMsxcm9lxyfdGKRmQZ9T5aEMzifzAV0WBmczD7WHNoufOQpyGo4
hOroN/ig2LI0wGFCyZLCIzQhet94jAv4BNFuiivjxaDYYl0QmWL6tEhbAkZcCMdW
oIKCN0uqtV6+5Lf0XfxvbncMdpqXu5rR4y0KfzimsEstFjFb9Bn8WViaDUYsFgit
aP5ocalnakaJUWCOD6h3Xpxw05jcEo9gmxwjYtYkivjQuCp+CtDThIlLwOGTQDLc
5Xi69YHnJROEnzL6Ataovq8YJdVFX1yoYh3mb8lQNfm8CazddaAfkRcbU3Og+FXT
QBieRBA1C+kAMrUiTF3rmObsuKSrdwviIFEX00BB8nrVciOBbAK3ioU12w/iLxto
Q3Sv+XH1scWG4nwG/faiE+HCXZqPD3l8+hSW0nmN+YqQCZY3IcjZxNATCiB3QqyZ
dHiaRqMabUKpXEpzhV2PAqIt0+3tQwmRkEVPnIheuHcKV8DsZNj3bQRbZ49Zk7i0
Wyg9iVMN10f1WXIEObtYA3g8T3f3cWEXpG5s8TEMRMmhd32Sd79W7pO08N/rgPii
mQA05tgX70b+5EIyIhzl82pMAbLGzLjxQOZkMRq0f3tk//DzYm4d/r9ZqriAOLeX
H9iyXJo6v+qzQDS7oyndmm736TiBrTkfx8PuP8iUNO88YKrxxNI7/zlibw9+JyPw
52Z1R+fzO3nn2LgV90nuVZUicUuINthnzHvFPqVdjvchQRH8TwC31dvJ6/evpJ0i
ZOAs/Eue8AliLwQYu5i2evT6DFwPCSCCxLr2aCyHZ2+Yre6PolcQ+jwMbhGmutVc
UCm/rjaqenC+VIhLfsAC7rQSZiepUeLyFckKIovvBOhCB+XLt6vrOqM7u+LVjOWz
E/pC7aXlkv3QVJ03v0swTIVeFG8GhmJ0hORvssTfCBRUsfNL58gHKDflb2/SibQR
LwChHrK7YKNtVu+LhAedf/Nqa8R2AHhMzPm/2SpkqT+ZaclLRhZiRshwVxPfVQVY
rtJR8MbVIgKJFRVn42hUwX8mPngE+16jwjUBqZswJ3J40k8r3YyZAjkC+lI/veMj
g5hNfXBu9J7M9sHI1DnVHjc0kZrQr9aJIgXx3JK9jpLmKRz68YpJv1LJdcTFr7RW
bWKtiSeUMs2jlKpDxM/nW/NIo0r0Ywzur4Hmqzjj148+8a/q/PY8n82f5zHjjew/
ZniaBKfpc8Zw8puRCZ0GCpMpBkUmTt0ts1LL1BwA8aKFVKwAAqh/pA5PsWt+8HAH
ZBm1kbYoKrQxFJy6eHzTyi5zasOezMND6hexmcQrqmy8vDcf/Suwp/NSNdNPmSE5
AbHHtM477QxyQ6kN8tTaEP0a/WtuTX5XJF5AABta12JxYXmoshuJ0Kn8lhdzQwki
sK0Ac8ej5v2nzZ49h7brR22GA+1nTEYhjS4W1e8BEZsw+YgXKKc5c/LtStluB49g
RENhN1iah0u2AYE4w3fmlP1Z/kMsIfaxb/KIOITO5yQlBoJ6oAIB/wB+ijlQqNK+
YzQp2Tkswokq1bs6+Vxi4gPu3Lr+4Fkq9lbg66lAbIPN4JafgZMXAlauX2wVJ/3U
2H69LK9hb/uWdDzwDkdIUMkGo5AcPYH8xtZ93LkVbzkjrLMgi5plpyFvCyqT5gMM
U5AgP8n6DhaLplVy+r8mrmt9A7uhcwX58yurVrAzQfV9OhehHwypwZp3P48E1yGU
gXLIEPcT9EckgNy+OpbIt1taj7GIglalpMQg9I6bSC7HL60WwxLdO+F6GKZHmuoK
3eoQ4Rk2jGzeYy0IMLWn/eLzNZlQj0H9xd+9ZA0YFM4tLiW7iqzIl3rxHLmYzsn2
3GvVxf3XYVBer+eTFqGoO0+Jk7+Zl1eEMulZ37i+77eA6LI5X6PTWoFkfmmROLGc
uYdICxCGbZICT7MRCYgxQp31aEYmccjgr33/8lPbb5WvNy0fuuDT0A9a15hTFvQx
ppWTjfyTsDTzOYpTCeTYvo+qm4Fq8f6HXMTZIcp3tWjO99bFy3Xjagci/mHm4Ptr
3SKZlyO+Ts6MHKpBFVC/+uXvmrwbm/CE5SRoYu+5Uc6LmncIn+AmV/BpxH4h0zrd
BxHCkmEIhzeMOuMsuiB8z6P2wxIpv0YNe2HCMSRPgTLLocE2FlzwdKbHgMP82bMW
Kfg4csdqYFOw7N2SykxO6dsrgZ/4fVZUmYdQ7UUMNbCXQUeCiWVwgQKrIcMv+98E
6Aw2m+6JNJCx6GGzgn/AxUVpN3ObFr6NVM198L4s/ccb7eAV3HL9uejXhi9ZByB1
te8qKcMhQOJsatAtFCXImwK9ndPoWZzbwENRjdkhAq/WnnEvW0j0BBpapLwgjBt3
TYvSTLfqrAqFiS7HMGzJ7nSMmInSIxlq3cQgIOv4czuJmTAgBuqEF5Ko60mOOZCi
bt/SkY3s4RFhcecbIQgTasIxp8FdM0iFa7v6gd0Yanw2McCjGn/GxcegA1eORUcF
FZt1+oxF6PE4ou9xjZuzrLV35cFKydiNiWTHY6IeO4cxahf1SeMKCIZhTsRSXpd8
dme4mpC99Uj95/x+sHI+4mkoRpxczGoR3bLIqUpy8CDKuI6YG2MvlkPNt7j23m9S
/stpT9Nd7FXr+H+l7WeKQ/7EYl/VTzuc/89py87H8yptDaGKx3cWEd75xzLaENEV
jf98R8cPYLcFlX/a1BLus3ByZBcWvX7a2R61N4NVOTXaqmZ8W88cUbq6M2YZ1YOD
kz0It4SdKFUkRf2U7n4pu5yEmWW2gZXRQdWIPh1fL/I1Bggpq1aNuRgj/izU3HOL
4IJLQbdgRnS48SetNlkx0dFEjc2C6LwS0QvJbRXqUiw6+aPKAlkp2x5wrLGXdVx5
Lhiz+iIBVoCchtQ6a9jM9Vr5GLuv2eM8w5FL0SxAOsaEzKEeJ8skB09T4f0uF5Ek
pZEaMSz45FKEYcXN7NC2ExXn6AINg7riqvhMV3eRNihS/vHxjYy3Prrg5pUHJgjG
oQ/6Ul6bSZ8MG5TNYLtfFJnV/e1FWYNuzJpG8xcnJadSa7sR6Jz7Z3hWUTSA2XXh
4Hue3ZQvKjwlxlk4lnbzJsw+3zaGwel/FqYHSU1m4TdV5c75ZV/rXTETHXVEcH0g
aZ2cOEJ2D4nzLTg6MJoRUnUZp4MumlPwZrglxfMBEj5ExHho4z4XPfoRU6/NKVjB
pdVDcvThMix6LkGRM7EzN/1OdyFI8UlJi+HTerm/RCwx+a5gfjJqrL7usaHPV7Hk
V/E1SXS/uPCH2Bdd3IRv/iGikK4sHaDnTd6JmTS9QKOddkDtwXGF0eNtJMX/KJl3
+mR7hzpoi2hdHWjGO4HG1zZrsWiYgkRsv0App+g7QWY6sMVkR/FORZHl5N6xTwRu
gvQWM04KfB0B8UAnxmtrivo2mtiA8ic6gzQ8RAxCTzGd9JvhfVCD1vmcpAKp428m
4PpYg7ry0hMdI4CXc3+tKmHCySttwkFicKa1thxZ06vILm2k9+jwpMVW+NR4vGoN
aD6pT7LzET8iN9Rbj+IpbzgwU291MVRJw9GeHu0hwCZLxJUjh34uoXfYrl6mMKAM
f1uHs0xCXUCLyHLxQB1U6rk+n71XH/tD/6Vy7qdVGkt/JITJ2PVhtmIctIPyv6Sl
GpPGR77+ctEEcyRnx9XuGnPRg8itxTrW1pzPJG1A9TTuJgGt7zKewZ/PPGVgkXpL
A+Fr81iVwAvIbtVRE+qur5jSnjj9WwMvLlKFIYd1Ew65QYUnTFlWpMPL/tPjYHUD
U61mxV+gQA1MnhjwDWjd0MMzh88d1nRKy9uiD8qVua6eCBr9TECRIOIu0urI1KiT
8c1Qf2jCQQzbO7MU1ian557ZeS9rxFSz3PFdzbodPjS31zPpP5UJZMgWEmv8UaBb
WajyP5GFn1VWTqmlBV8hsrPhLMoisogshYCKp4JYh1nyHQ1cic0sbtycRganoPw0
vHBpAnB5fmGBssKNyPYk16AynDRO/DdbcXKY6dRQaZxpm4SsIGDtASBxog5VA5zu
42dOI0wKNcJPs+alaxNc2gYijskWJR3ZXzFbiE1REzROtU3rRxc4pw5K5Ujr87Wb
jw8EpXxw094b6bbYe6uxx5qCMA37DLPk6vuuwhXMKnEMs7uxdEemW90d/zsUU+b0
OpwKQ7Rc7mrWyp/XXcd3RrqyYCNhwGTM6uXr3JiouOPj+X9YXr+3HjApO3ArSYdK
PaSpiPVmdbMODgrnW4Lx/VJ7uXYiQRmZMy2I6+d7vEM0gp6IF8U6VRjvJk7OmLMx
m+uto2l5+MvjugAirpsnG9p5cB5mVTMspb5vDykHX7tsEVhrlcYVhH3Oj04htjCE
aqCdRYOpdgTWkuPeVhQ51P8NlHRFjuyHH2DUJs4xjTCSG31XV+tfZg7Cx/cOQwfT
IUPSKLV/UztGH61lB1kYmeC6GbD3oA0qXYAGx2K2k1FQ1VoTZbO9XBftZPOacwWS
VG/S568d4bYjWcOnEssYn8mi4MdIig7TZZaQlYZLvW2XmFl6BKEAaSG4UbVt2yzt
pV/Ty4J2lxReJDDJ+Kx7YB4oeNzZZfRYd+xKUKDfpsxqtmwXqbJzVfZp9EXFZ0LP
OjaRe748t9kZ6JoHlzLFluiWJld/VW4Hsnw6C0zwGLrxBZnn0vMOouuamvoK+IJy
SrRLUIJBbXhCK9R8ADJJhjT9gUlIkBtg9qtCUSJFr2pCS2nu6HAuJNpCCYlzlH8f
LG03RBJQaVhFMOw7GqDyJPrBaFWuTpWbB1/g9G21stGE2J7G1q25juGF+56P0Dlh
DvI3svFBXNxK2AKHMkzjXLV/Pz5ZFy96Vih5CqAW5n8WCaHLWwvJQ9JMjEgUxesB
1NZowCRPcnFTHQPT3gAZAvKW8LdzT8rOsq6Ak+N6ofoAGZcanvCZmV8AaAh9nQjN
rwhMhMN6xuCtwMZJMA9yL4NpZKoox5uWZacTFR1Bs/vBN+UNCpXWNL4zAYxTHMFd
iUkPEjhi80fbOLwHcGgnCoxx0zuL/xYQ+EoUEPQc+eLs1Na4yJsXP5LE8VUWfvXM
6G+IiBbLoBgcP6z2yAz0r2aoUty09ZhJHUyMPLueX0GqvqYP3H4yiQI6tqrH0UCc
bI9acbIVj1B7fZORfW/igEe9zkaqB8dfy2R8BcacAv3oJ5Xpndyl2rrQV//g2H/y
JV/mbGdfhG/RZwS6IMQjVUQvxlTNLWLyLh+asueYBNOuxBV0FmBXfd+mrqN/qdcu
LEDUHAGeUji+SfPvqw9NoMZWnfRu+rNjWg9Y2Wvrm2mbosFAvg4t0L4ZxjLfjYd6
QDVq7JmNrGzhJUJRYSkRgsOCJR9H+h0NdEQJ1/e1RlXO53xC19kT8+O9UTTa4sOZ
fEL+wRs4V8beBVp5a6Nip1OAvlIhIwRObFlp0j/Z1WE3zoRW3/b6cpTHtAYAvHgr
GqCZRiiDYWUkRa0Onz0Cb8kdXp0iMg8vFWok+Ejd58Egbv4yrhET2nHWspLPwXUf
24RQbOS2q+fTll4Oxhr1hpc+mJ+eXuIkOeR+Y67sjUgLkiuAusCUspAMmKGNyhUi
4p8o75+X/ohh4ZOEdoeC7xEEjjxXQwQZ7SaY/6PXx9Fl1yeHe+Ts6nJWfcSq0kd0
DT4st5vUX1RCRbNuhSOV+rs5a55iBGA9iQbKO19fAUa6z2w3JmEtGJqKC4oa6Zc+
MFmMdyYC0nerV2cN6AEkoAUvU9Pm26V2wlsu3z7LkwPeIhCs3OGs5T5W85/f4+6N
TSrJQJgKhS+rKjT9U/WrGpMo44VVpmzR9Y2z5c2bBxgAlDzj29KTV6imb+UGTrUu
Vk10haXgwL9+NdAKq3JFfW+N/vw+BAjvDsAXEycFxjDIDvzflLC4VF3QxocYkxHL
lVY/1oH4mGQ5Se87hGq+GAx+f/yZ4KYNLjtPv8qaSklVW+zIknNQ4Q1IDZGwY+P1
Kb0QGCTQVWKyS3d8n+FDpg==
`protect END_PROTECTED
