`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BsroDeyePnZSZFer+/JOrZgXCKLQcBIWyudarolfTEPf0CVHoBfMwuj4l8xIilLW
MyYe0SmB/oLoWG1Ft4CFy0aea91EPBEriRSyXzV2eGM8OhDgT31HwJk9/OgF/IqY
IqnlBqqKTtuKoy8QLyEagOE3ZlpxRh1GErSmFgxWXsewSdAQxTtoaZHe8tZINd97
1AM/UuHVK213a5RA2vIiARpMOLxOFwS7wsMgjXWg7jrNdG1TiTaEVJ/hdwlSE0Ef
0gFB/qiEntUVFauNFFKCmm0ry+/g9e6hLBk9tBh7urk22egXswmgKYuk8H27SdYk
uuJHods4i/Ap0cBgbtdKK4eJ6hfQKVnhSx7FWTINuZVqWv3phdSeFeXsh1o3yvR1
E9Erl7L0FVh5r5lIfBB2YSSM3pZDVh2X5uocOeXUsAKiYOQi/VhbwuZ93FIqj1BD
BmyGZZyjQfQOWfWpGvapEToJWSkuEitOajd3RmixUjVd7QbNMhCNmjxe9siVusAv
OG0EY1fLNmUz9UooZDv37Q4C/ueK57qRiL7unGtALlvG5v2gpP8AJxAWJtd5iFsD
W51ZwsJF7w9tHcafKqOodhTEm8buzSVdFD40jFoafQ0eTCIC7Av92mg14vIfRCVT
7lr3nsC3bF8BL+46F6ICtbY2APMeE3U584T86qqL3lBBeP4lCLlzaKOGFwdUk0SZ
Ghklz8pEY/VyHz3JuOCZisIibONBGKUUKR1goBExnZwBqh52TLar21LNoVFjWnEL
oS+1Tqq+G/gttnua56WansjL4c1fzBND3APBHGHwauUYrJ6yMmOxE0hL3oT4efUw
GH+7L92FdHu9nwPWhimzZvLhnMoFE1VJU+t5T8cRebru+G/uTOfrVGv6upodhvnV
rW+XwkVk7G/32WuLYpADw6SgrlBfCSkgNgoupS3/nWcsGRjF49X1LnsIRhwzeVs+
jIWAJcXd7/lsulyO5HhqMQqXCByvhXIoLLm3z201FCUDTdfNa1JY6RjqrdmIPuF/
Eccl8C9O8/IGgzuGjFyCbqSyBBhQ/XlN5Zpajz6aR3leNWF//fOP7J46fvbzSpoy
JekBDDnU5NDIye02yuatlT5c6CM9RJSub8YjzID9IXnYqfnRXkOQ+Kg02ev0gQX2
lKrz55IhmV0SmbMQ2yhbJtcsRMVEToblIzp4gVvfUtQDwNUSu7gt43KKNgtomR3v
M4VkofXCwv0C6Ec0VODNVYuc+9GqxhNZzS7B+efdSBbsXx+V8gTc+9X2M9Lq75B6
v3xmpXPCYzMHZRjMOHWvUboQzmU+Tf08nuPspacFCcsDV/ptvzcxGCYniUhtjUoz
/D/aG6Po1tTfnQpMaU80OLamXMX/vEHjd2SHl4uIv6NnLqQRQWmZR+3wJNxaH3gw
mxG8YNbBbsbAwFzygSG2AphQbt8XHKWfxw6M1uX8RhbiaebFijqSjd2oh0O4in+l
Ah+Ix3kYl0N4/rGsNY/bm26CrL7eOvNR7FUbqOqNk6sV2tSDKtslwDEcNmLKsCe+
uqXs9Fx7Z92r4IDZHacYrlC+GLL9laVM6I+FgxKojFJkcwDmwJd4Fe3Of2+pr1wT
IPJXFMJcKhvH0wOcbPM20aHXbl+LS1heC5KIBYwUYNkwwms094N3Wm8bTPRiUaDG
z5c7Fl2CIDxOuBRjyX3xXS2iZyganCWI5EAtHEkkyC2moXMu9XliGCgF/+ufniKC
hQZOULdlDn9H0np46bkWWNOBINjmXxu55hWJlTu9TXhLGnnRU4nBFQyJXzDXMXWk
tuAcpYuEUDHGyWSzLQtqRIbTEbBqfNdeNfuq3cgkiTt8zRzbpwaQ127KBEeIOczp
uoXgh+FzP/yNRl8/ZDvuW87llf4L/QYewrIzlvdRd6FB4Bnl/viadI12FSCAGRLk
CxMDxCA9eW1z3+mu2u0dwlg/q3ki0b43IB0AnY0psg4vLfiGrkjiQPgn56fwjIY/
jSV0GFqBv+BPlwBZpG+SUh6NbK76KvttZ9g3SlTWNjwa0QpKpGc1EJpxnAc7eTD6
`protect END_PROTECTED
