`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9RjSO03itKwLvErNoOQEj6r7AoaqiTHmATSkgLUYh8Hk0X2fRwu3uWc8twDVs0Qw
G4WcdS6MSDe8hs+myfJDbj1WoNTFSXqFdpSNNn/H4eUkBaFDJX4YEysGkOvL3ot9
XrRF567JOjUmr8NV77YbgX8q6Wv4dEhING0QJMYKT116nFSdxnSToDzlMVYBLBMj
y6kLC+cg+OM3wLiWzlkktCwAfNwY189Qt//L2Nmb0NHRQ4sAW5Koc6VU8ZqjdCwG
Ys+793eHs4+jDWzvRo01y3z6y9crI9OYJ6JttJ4x6KnF3cr84Dzk60M6ol6oYnkZ
F2TpXjeLxLukWCf3oVaDad3IMqoTcZhh+z4m6BsrNRKHnndpl0x02l9ULTtNuAyS
XgCaZGzXwBdkSFF7Ps5e4mOuKuuecHwLbR1P0DpmBaQjM2rBjNYHi5s1qGpy5uHP
mjNs80KlAJTZ55vA2VltEhYV4b1rpWvU6+8FJdeyJTQhFbSFulHrB9jvy1fTv1bK
3PFb1xkDup4zA1XGNlXlfyqwNPEiTaMsMRn8rKogxVN6+kf8CQvVlfbJPoX9h4Bd
AB4WOYEi72aFymwKYwXtmOYyFlNt64z+8RHtYMWzx/M=
`protect END_PROTECTED
