`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wSwO/8L/bDk0UuyOkW/tXe8bh8fd3XtTtXJ7UVC5G4harIskjEi0UhiVLcA4N7LU
Wdk589db3KkWPKXNT6gjwJmyNFCkCP8Rhe0aGGOR0TUS2kLXK47g6JxjeO8qri0q
fsl0Ir/kSbBuKpvhkwnv+1gSw7htbd8jjH8qENv5RNjDry0Kd8aNWoP4kGlHfwcg
jfA7cK1BwZ2aO5O9NIj0lb1gIM0ijIVmwbquI2nCwkHMSpocQ6xlNqsgFRlnlrF+
hwe7dR14CzDYGwP1pSmudEw4zaEy/35aqnH4TbKXcsQ=
`protect END_PROTECTED
