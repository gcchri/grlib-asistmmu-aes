`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rZoqz+Bpvpc97jTlDOx9AuZMgNaEZBcWXIm7rWL7l/ONZax1Gek7YCX0pSOrKKfC
eWcvqGXVRTgimO64D8Jm/9mrccPwdMGs1DRk9D3bD2ldSUuPRWlgj2h5UUSFQMYD
OeuDmemUSecvrQeMFCnydh7IEkO5kSAUYO15jyPdgGRkoEbCL4E1SYb148pc8dUw
kJy8tpAMddTN25/SZxYWv5FTOumTkyZgyxpoHQlchXIax0t7I2iYUT8Bt/6U6vx8
6jJEd/Fu92Pf2Lf9RXNO3xAcL0vYXnK2wc4m9v5SNHHZ9303oN1Lo1RPIFT5BqoW
yiXyLRTYOZTl69QCgq5mz2tnEdvx3Ro8zszzfxhwiCx6vQdvNWBjFeCMEVIwA6yR
schZmUElmGa0VSK8qUsQ9HfqaCjRx+Nqgdtjf1T3qnU=
`protect END_PROTECTED
