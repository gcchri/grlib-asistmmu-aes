`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NW7USViThrmbl8gp3l0Af+8VUXSRBUb2GtKA9g082prOxLKrMkieGL3ZDWOLQ1U4
FYdGqE03g86qr7tb5beJCtM/2qcjykPLe1U14PkurDWchIaXMzR8LJCFyBA3UvID
zoqkCHkiATxU1R3XNa7UvQ7AeX0VbNiGU1Q8z67pVyeW+iHXfH2IQEIkJal0YgRP
ThdIROlEESo0aFQgSxlwypqAmyp01EdvHNi4Rmjdv2CzMl5EZeTWGW7cN8vDA3n8
iwKnwmC/qy1O7nJ1y/VdMQG++UKs42U635Ac5NHgfQAgZeaIURBW/B/GUEoX2/HY
rA2wteGPl8B2uJOnitGJwTJaLnYJI9cWyA+BMySw9jS1xo6t3i8tztWR7FavIqXz
`protect END_PROTECTED
