`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qt2X6rkdObZCnb/HMydYa/vO62cyY6pdi205b5dBxwWW7o5jy/CiQ7xrAxQXyPOF
4axwnR39FBTscQoGIoPod2tZ9mvtdGLsA/cL0DzXfpHz4Y07VKr3M0P7VlmM9QMm
zh8n90n6AXtDdBJ6vWb8v6GiKINOLnuwCWECyS6mVSTZQdVW4lJjzwmmmd82NDVf
GtI4OOZhq1L1t9P13MChuqeXHW4drkxWF4//v9T+tNe0Fj2UPuc01NbBZMpVVXp6
1HYA5txMScVR7LxuGwwocZuTI6PG79u9pbHOPMSNFyxvlLxk+/MIC1UaT7Z5maEM
LlBBNE8QYeimr1u3/FHy5WD19fugrw02bnef6nwi75dGH98wmBgxA+PfeMnfwFni
`protect END_PROTECTED
