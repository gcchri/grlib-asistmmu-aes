`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3hSt7yvaPHUnHGqZyNliLR5eibhc6X/GRKQdhzHR1b+h1VBMY6C//BWTn6rEUDoZ
bx+Wst9V2XlVQ8xUYyQbyhYG6DJXyUMg1+P8rCvXRigE9Sicz5LZfXxpLac5MGX+
/8Z8k7wJ/23zmyFr9HWmsCNrdBuwBIJ9oV1QY6fLAKlVbVPUpBfG3mrjUruBH501
BkpwYvq84nxkPVIj7GsxjCSdQhdFGeg9vdl56fV/RxhVIWUcsQ+yiFruY+QZfTXK
BInfwW+ZoLVzAGQ+rZERewOWzZMADbDn9sg3X+qLqRisNxfMl0cJsFda4mnO0oaH
+nPLjgmQ/O1EOzucQY9vntPmzyOWU7QoKU7u1LX8mH7FAMr3m//fIAu+Ez2EjBDG
XK+ViofLCsgavVbpRkWxQFrZNlv5p/P74JXZvsFkUI9Zz2lQ5qw9ZsbkSrkLtbbz
xWp66rm91tigW1lcXO83nARlz9SYr1Sg1ymun1US8+U2pqLvm/E/I3gG+Mw0vm4I
FNjS3O4kMdtsMtWIJ12WlIoBies1EF3OfAKAS3xFP8iEHZ72GKd+vs8i/F8DimMW
h26o5YqTOGx9wFypWX6d20ImaNsSWggNnfOd6+lAdZvlZG+dbumd1GEew/Qd/v/p
lhPnikqXxu+6ksvFNnoX/gQcIjALobKGo41XaqRqksih81VJD1dpYzCWNynvqFke
lrYf5zPC1t9biBUzs9dd6tSNs0DG1I4QUxvSl54IjR63PAItKah495Ts/mKMIxCZ
cv61xSFbMJy0zq5B1az0jw==
`protect END_PROTECTED
