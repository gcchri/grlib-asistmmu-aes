`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gY8Lb9OXWJQLsTjGImzF5whvuZOBH7nW+RqVDM2La6fmKrEzXEQfsjtdUHypOjIu
WAMeH7CvfSoUqQgzghz1HW1qPK57IUZg4ZoYcHrBIQ1RQhtOUirXBaYCcxGf6QSR
g6leFTinxa+WrY62lOoQSnG7pAD9Vh7ddS7nHWWYXoqANKMblBxWad7UrF0U7obR
6O9qWOgpbatZ4BJkC9dgIDeVOeUTtN9Ho8/5SFUeF7yml6y9JouWzvM3XjoOhbB7
k+CjavR8pMZIv5jPBrLHlrmtTJEOmkMMb+BwclDhgzQ6L3pwh1qRU1FSTZTIqaRN
Io+QHJYRbr1F3a/ybXCiRoRx3v4XQaW/j1vad3EqELhKaSJWtHO5jGdKa5J83Job
x9IyrFt4TiywhVAipMWbOHySEbpCM1Yf8IuejnsuUFk=
`protect END_PROTECTED
