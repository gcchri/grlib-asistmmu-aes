`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OKij+bi4IOoAYn+n5/UXUYLfDQmuNGFfs533WR9hwHNf417+bxzGVXOgM+OEihE8
F7FfO/utr/f0DfR5DLkO1afTfEjo7cIYeZSCBTaSJJ6FmM9jQen67qqPllOkSnt4
OzQ5NkReYOShrQZ9zXDviqPg8bUkAF8J2gDd8mIxMSaiUXMgrf58pjUc21K2+xfB
V+CeMQusll817EZNKzgDYhkVkNpx4Is/6w0XPg9/TE3EeuyZfkiCoeRBPMSagj5g
vBBr84P2Z3BjyWFmKMsUJpXIomz3MpaZmxLip0SiqM2WtpjDa3MAVwvw5mzPRpFW
TijKDgBlahyl/98xTcGL3ZOVigDco6QI0GTOF6M0F78P+sCK9bi+GyvP6nTrEFP7
4gFWBgizn1xwnwe8feHwszvdqFpYfgDOYVIUva8CPPgscA30gelS0wQuzSP8eMNQ
Qt6+goE2aTNdre5H7Yk8aO6chkVYrqvl+Ly/BNRFcDdBlAHZgFhmu0en+cuArN14
d8eAj+YhUWoKLECPsT61fq9Dy+NDjzroB7Jbv9Egc7ZtOjS9pvLyl1iGgWFCG3IH
imFVI9C/NC6xMs35zxe8IxDIDz65/oD1FWf/GuIUxiVzopNX4FLckPl7s/KJA48k
pL3Kf2vqOy+MeBCntdMMtHMPa0fOTuxOvpcmC3B3Sn3YUi19a0+ef4lBub2wgxbH
9QXUnbCJkaMhaDA/60yxt/2G/zt05FR2t7THtWds99I2jIOg9iAjNh2dsFPzTnql
NUciZgV5V3MtC/q2qUpXEAnkzqxq7wt/l6hWTSG6qsEEGLVmzhOXrDqcD3PPQd35
bQ1i6W3pjaAR2IC2loBsoOqcMWPfgyzuenDON1lvEMNfK6kcdR6P7zk0WrVHaH38
/x7ujD3iv9YXhc25b9EG8YBcDmZ3kOhVYrumfPutFwm7kEM6rY35yeg/qoXAQkfg
h9mrqbZaBgGJ+Hq0IUWDSg1GuKeSdHz/3LmteQ29MaDdHPtJnIZLFdA/Y+kUzrhP
2alzYNTkW+mHPm5F5DwNyIUObXi3thKu9uAMVUQ9DUbvtgvr3yES9Hm64vfMUh/m
iAslrJ1/unYcyt2uodcvyqkdY6hL4RmaRm3yVE5T66EF0ayB3aUeIKwx7Z2PLM0K
RnYQvs8gcwoU4xvcyGjP9n0iV6SBZ1kHs+t7cvYQi2hbjBuyyhNjqL/OeAuefd1t
8Ilrhxwy5vwSiYCxpXJvgRMTLgetZ0+ZTlnqZ96V5j/I+4t9H6h71uwiWMuKbwD8
wAAUyWXEFDXaINeuf2FNMpwDkwLkLOC6G3olJyDGpCbbxjrqtK6oE1g1EtbeZ/+t
Xr+wJJVYu2F6oyrMZ+AegRvcX4bgrkoOjH5ukoSmYqDQp9NNwX0tzXrYgJ5vpWy6
zwGhHOYuKiII0VVJ8S8aSYIPnaBL1vGPXn0P3BHpkRJ+xY7Y0qEK4uFdgIzUJFnt
FEktB9bm0QSEi9g9wfC6b4z8MiTO8PQOm/SEUblgmahmTExCTQOd9CtZdMIPIvv/
WBwb9BaklwCJF2QUsMkJ9vy9cccf8c6H8L366PPz7LjlZw0/Qnf7WvCEjf7XLkqH
xKNyfFgmHykFnCku+8Dnsy7r9z0mPnROBFp/aJGwSVGpTmyC1tvMtBdL9ceikEJj
Lsp0Fa1kRrtIWu7yCKwQv9xpRRNScPprlqfqSfE/ZZTHrkjW1YSCpqWHHVaQ7Qhj
O+EwhifupI5FotxuLUlvJYqqFgbwjqTAp7ESWSQwRSWhDSvb38v/kOVBrNmB4h/6
oLKZSbOPQia/KCu4BL7Zzp4Sr1EYPSv/atdeFXs2SxMRXg5xCst1W8/CvUePcfcI
su8c/I2W/JOHrPgWvKDQgNWU97VJndZLlEW4utzJYPEglyaQb7T73VPMQbGbE5VU
9ZZZlbQyFr05r+wep+hiGeECuLww4t0DZd5AQV10g1+nyPbknyivLNFay9vjXhNV
rmT/eyupYeLz6D/OW4Hd1X4GAVvfo1ASx0H8JCpJwEpZfCJl5HBP1FvWaio+BA0j
FUkkGbij0JIgnwThY9qcC1tDjIAcuHixJLlzgfHmWnyAfDX1V5ozzvMS2QVJQ8N0
KiwjPjIU1Jkga3x6DdX+iQxcu9Ti8+lnmErKwxBUHLcCZH0T3i0nWjqPktZo3JzD
Ybt8+kKjnrmcyhn2JwqOWw2HzOm3lw2A8fxj80mFPfRqbH7Yx5ZfnqK8w0sEdM+q
c91bqn9L3PhtztYbSiq1jMyEtO9gg1cOqBVNh/MeAEbVdLTXvtr4GYCkfqAjH4Ji
/japjSzJ6zJElCUDFecYmOxQruMFCNKm6c+TOqH+gnOpTERl1HIMbw/vdmdsU3Gk
zwZLv5toU9wIUqnPmv4XCM/4BNJd4NpZjNE/2asTSq7t+5oxZQrIQAjyEb7Nnp7j
/YigUCD3P260zTVAmzj5EOslGKobIFF/rq4eZRVZp/M5jOUH4KXTBtew/Wc2urcw
j9nvNALoisJXk/BghzraNURbHBV3x9KwBjokyJZ7glzzK/Ju5qL6tuIM3JF3a+cc
rhS7/Fg213i4ubANdBeCmE68YuYV7jwtLjtrtc7x+hplACQpJkno2y8qUmcT4feE
GaEE3edE2wVDnnEDqeBQfjcWBNPBY7RI+QI3M7B55r9LTMXyyhg6KYFpvtJlzOTe
FJeXQGOKrp4RjX+O8DaOiUhaxKZvd8A5UyK0eUBxr0NVZqTy0t+oMYlC97T7lXGp
oiGwmy6yhbW4SIsoK2DoKQ8rh2ZmQGQtsA1P2lVQsbrkyQ+pssGnDGrZ/o6J/t3j
HQkvkVF1eCG0QG6yzOhzzH3hH2x2d63uPWWdM9OeP+rKCPBfhvcCtvI75v47wR7/
9Li9POfPdMdJdAR6PV2btv4TgdYgaVRQ6q/7O/MB9x+vZ9nXSc3wT1TrTUytaPWr
6VYD9zLVwcqdvsOBPhYq0HbaPAaEzL3fJP/8PS43+3s/4zdGAjUe33PRZ7obSmDd
arrUINQW/zumiyEH82I39+/Q9FK4E3cIdfXjdPe49virnh4upkDAGhbaOPaSkhtz
iQ8ed/6jyAp6C+SKyR4UwMGx5qWs63/hbgRjHXBl0Bs6TATvZh/jiJb7C/NYikhR
aIbuOLEPaPgOYT2HN3nPg5sLPD7xMoJ4sbMMm0yW3cq5JyPQC8UX8bTEPiaqDmdh
V7dGFJoyCJy9lwMYs4TxKLt3OGVA1Akmx5vDma9R1BI+KOREUVUtDaZbVWsVfXLR
r/e80M/KElv2AUNQfE86FmQuNL1iO4IH45yOXZnqAnQ2AEtwwroM9rcHYr3UI1FW
08JPoLfRbAprg0WQdu3TENBwH/iXfUhsBSPcZEh53Fsy8aAOZpfyWfLyONbLBmlJ
YW8eNIsggSOeYCGwZ+uX4Zgo8WZzZpvOe2nfwMYq5Tn9YSQlIgdvAPvJ+YKbepzY
Ge2soCgB+xebaVdfmCsnGfhKsgr//dADaCG2Oe9v4EQA7CXLFCWsfYb7DIi2v7AX
QnvHmgom7B6sbTuDRBXqvHSp/xe53o1ZMa0og3VdQ7PKeh/0YhReNuXyuajz+6DE
1wZSqLMYXjzb4aynmjsJnQ7exH/H6kWjCaQTpj6+gck=
`protect END_PROTECTED
