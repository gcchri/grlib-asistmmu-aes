`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oE5hlU8xkTI6IKH6QYsN7CUA6EviISsIBnDREQ1obhwq65Q7IbHJeuEFrACU7l6z
d1VyhQgI1+gBgMlyHGEWg/iQxG7aCygfGmdtzcOYSxF104k7GE1klgRDTbFxRkBs
1YsK936fFsKJ4/ypj3v1UWUUu+1kHCbV7NFGzseuyuBf/9Dplmunb6jvuohb19iJ
7IXV1ib726Kjpfj/1w41xwF9CikDIlPgrYM6TuQLhdr7D4m7EW9C4NmTqRXXpjk8
EuFk6xqf04yqcJ8XhdSGMd/zcdI/Lzrbza10QuAM2UDZfYV8ZPRyXmUC3WUKN+o3
cMarDYYHHFDhkbinLuxsMA==
`protect END_PROTECTED
