`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qxFvXjpxuHUIfeoXqfudF1z7+hOuA7zXXdTTHUKk2Md802nLUpCaA9hVsH/UMso3
G5Gh1pam8bMw2+rjqBZSE/MPhJBCl4U22PrJW30HrIGqnQjMCuVI61N52jQNAjRH
OfR7p/ije34TNIyx9MnJSpElMQzP3GJtyFqQ/yRfsL2XWNfEDwlPZOoPI4/DkIXQ
frXoYlvRiXxZrGUNJHOAobVM+vRbjqP/NidI1PJn9ECS1dNES95Wk3diZZLNPx+V
z8b38WqumJx9FPGlscxQoId67dN+LajzxulFWcAvofRX+AP16ZbgXj09nIb6aLcv
bnzOWf6bRBDvvDbEnR2WkZJ+eq4qkKRerP+wHh54jQD6vXSic2vt0l6vOiiQo4PS
g7rNtomcPX6BkrhG9t0YrniAh7yiAFgNlD6c6izpNZmHu7t0UBUeCq+w4uQ9lZxW
`protect END_PROTECTED
