`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UKGUSuFRvGo82pBy546xmSWgOKtbXqlA3b1OOy7MVL8m8Bip5/pg7xDxo0t2H1RS
C7pLV7r+dYEiDec3Epd2ZakJCNmBYBN7hCeN8g0qXD74kfZZeB1zPcrLivIbI2D0
0Yt1nNxbD0FmHnnCzToJNwHsdSojDPmYvBnMvJat09PDS2xDTkmgyneLQk1uDuzw
0QnwAhU9Mw3YdvLaQL3ahCm3YWl0gntCtArpfS3mYSl5bwRhvo/57QiY5aBSWx9W
ndIABaXu+u7mETCkJQVGHdPZthCoLNO20AmsmngMcQG5ZxVTJdOt9XQjP1pOvRqB
3iz5lKb16LrNOodiHrw8KRL8HMg0Ko4kmGCNDp0M6u3Df2oHpDtu5B3JwMNQtO1w
xkvY+pDZdC7UDoE4JaF3zQ==
`protect END_PROTECTED
