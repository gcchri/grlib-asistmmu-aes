`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ikVpUlmBADG8tHCLvQqbwLCVVEkuMzDPZhKTvGLAPQIpGKz8P8gVbxjV1/gtVYwm
zAvEgROopLloPuoFO9/9bqTGrnIFHgHD5j48rpNIABTp32iTxRo8low7jqXbnkeM
aAwWy8BCrLBBJ72wDYqhBEUVQSpmPiykvqz8c+3STsHGZX7U9hgKBFwAaagBtPAD
yxpeGgE1JUGxM/wkevOC480IeU0eaOkQLQ+BpeFFtY3NlQKd/dPS+DDFx1yezWYy
kzxP/LvlXcloZsA0ZtkV6rb4P7UXGz/CZFjWuD6q8KPEX0okVxO6OxtuoytMsMTH
r7tdYFahFbHh+3Xq2bJCSA==
`protect END_PROTECTED
