`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/gnRR6PEM4hjWTd/2WjtcqxF9b1Q7z3XSv7BLL/XNwinnHmDKGjMhxaH87dvmD/V
fcy6b/OldD67MebmIL5Ft03C2o6M3nwx4FHfU7gP0J446xodKAQkpyrwLSPrV7dC
ANFQ3xLDJO4GC7Qk7GI9Ij1u07ndkY3hoT4Ff+9860lJbRFL5UnxBEhpcc4eIULU
moGayXKvpvNuw6GY/AW9dyCnmc4A7mzhOM6AmGwYb3tN4/dD4zEvILb99aaOYXz3
2gcmEKzRdVp50k5k+Hs7d68B4XF2DdSdMJl69BBtJfN+lh2GZGNgForXgEMrT8c+
5x/55eEhORSCCU2QKFIP7dltm0DWe3/uAm5zoCfdwpUtZYvtWx6WVryvGsA8gCgm
yIhfb81yeiVYYtS/cdcP3vmxluN8M7i7MRqoaPR4yj4ulMDIyTcKbVDc0vj0aYx6
BWFJ/0m9Jv9oIwUv8bLBTPFON03it7KfXpF/nN3SRYslpCgmnLwtCQW8TWU8tHe1
THujeDrKel4rhBwBiHfEF5GQHe+CfdhSmIf6txn6uo3FOawZkUk5+JUjawmYB4Wo
+7CEDSU6AY+6eupxl0SByAtPwq1XdhJq0gapR4L7ZmOet758f1jNSSNUJ73arGWh
`protect END_PROTECTED
