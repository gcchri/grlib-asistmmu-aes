`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KIPUOKYasN1Sgco7WQBUp68s4FM1BY6S9DoZR1ZaV00DF9t2aiIFUpsLXCEpgrOA
+r+8Ht30s1evd3AGPnFTZpAXX4XY/SgEHwzd03jyGFwYuLupZuXDzAXAWE0NrYsg
tM+7ag0AsD1Z6b23ZmHFR0ruXEdVE6LXJ6rDUbvdnbzWjhmZnNwCY5fLWAZ+reqk
hZdYBurX0A0J5zDjikBlPUi1cIxBZup23MeElpUNYolAfqB2aUHf6uX2ODTRaBxy
gJ9gGCejsITKxil5z+5GpU9IxRfv0MW4eOprtT9i3D/YRA83g6uBYrg9/vRWpqmy
nEBRdUa7mSM8Kzc6jAWdl1VthrTffmQKNhO79YZAg9nW4lH2Ty4Bbrc5UXRkE753
newxbAwYZqAYiURVU28kmMN8jeZgzkqsXSn+CrUa0c1tzICridp/SZvlQGEd3ZdJ
mpZ+h7GWbKsgBS6g2dXCx1+5M/T1tQxafBtuqazthJjfGGXOGO1H86K669SM0lDi
Io71FuLIiXReXzrKhEb2yPIIiYPbH6HP5XZ+KCfBs1uepIeKX/8GxWH4p7/9PhRh
pl0Qia5gqXYW2c6X+Rz1Tuqz4rO8RtCzcE6a+gr8GE5yVpbH2zBkN5ad9liRlPse
e/Uvq4RJLyXe/0zcNYMN6pVawnOoZioB2RVmNmPpRNLS+Tn/mIfQW8iluwpFmIw4
f3S8919qEioivrA/27ACIUp4CPrvpXU+zyiHHlU/AR22zRlEUOrGqRfOU8rNEPuD
CLn2p76QZZOs4B669eRDCtHQEqteTT2RoivDdG5gVnalKncXLwMiasJxAaoBkaiU
5VytKNI+v4MJ2O56BY5Rgv+HpXBHCw+caFUYDsDkim33o/EBoIS4Mna4y8pKlo4u
6JV9yglHc3LZl5dK4lIkbtGq0nwx2KyGJ8c/hlUIhUBfuyoztZwjZ+6atKV+XiIw
qqzLZDdFnowL5GRjW8YGz2GFyyj+bHeIUorWgzNmicp1F+QVtFbZYZh1EjNe1zIH
Rwzgz9JqvEY2mYa3cIFf/Emmu+WlEC+gBMnewD1+gWWlPHgn/k+4WcB3P21dN+OA
C+cnTX3/z4F15mMKhWg9Dp3EXc4z7O46zeIoJoB0tayWeImwvN7PtGxZ3b75Ecc6
oGNt2E31TLE+D4lH5chDpRp4DD9k2xSS5Eo274LIvVbdXHxnB9DNiVqk0+6egcOf
Wni7hiWgvyIQzBeX0XnPu7VIy2Ps375FBinSPccrCX3hhAf7Nox32c6q+5TO8LUI
WbyutleKKeGo3zK+ICw+3Kgp/YIBmuJYddB9+dNDKKst7LjfCXCAhDQwwGjrfZ7x
1LWeggLbRxWpeL62+4M/46mCFkY70eazTqjvapQ+E0F/s9w2YZx3Bo70eucfs/mf
jNPr4YdY/sMZ/0gigyV9rPja4VBym7TY+Z/cLEWvoQUX6pZMEJuQsT4vkOOeu5Br
Q0bw/yxw6Q965+rgEDJLMfZdTKfXFym1dIPf2Wb5PShiw6rbme3x4jZhK7RNa5Gb
`protect END_PROTECTED
