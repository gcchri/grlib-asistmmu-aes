`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yV1ElX2MMYNamoVlw5b9Eq5+ZhHmDbbP6zHU/5RcmNIZZAjai8nnaS2UVaRWUDoI
gSeXSiYEM43EG9mDjKI9arPScQJeskv9M5LsPSI79VfLntPCH2XKiFF2k/slEpaE
PULSxfOIOJIlqTW0Mujb1lbQWRA4xGnu1TUcxQtc3KMlfHwjBC3bCoq535SVo7gZ
xUAvqJQpks9ysYJiofJLEWbTLRKSxLBKkZgUS8BuHFHsc/uX/eAbFv3v6xJDTiJw
Xyu+Y8jhO6atqTaaJkskDhYGfxrVjLjTSDrU0CeRGF6HUKoF2OUkjovkuCUnnsrb
WT43yk4fTCL/fDXUb7KHoWUASdeHnS5wmLtol11uzjNVRXn0SbXmWpDvaY+mWgGh
bIvbuu2iJAhcO4vsVuWQRQra+pnyeryC/gyW6Q0hLm9fxz6MUAbNrmWCtsP39uXC
DVu56QzOkBO/Lv6euDQiNDjGHtjlf8bQVuSrIwtKAoWj2f3AFh20NDa995eyrb4l
Qg9GLY9qPvLgcLpQBcV10iWdB7EtNisUvqh9zRAykp15Jgg+Md84MaNEWgRwoy2i
EXY0CxiUdGTHARODE8wKtHDKMIMl5FHYecHT3SMa4Vs=
`protect END_PROTECTED
