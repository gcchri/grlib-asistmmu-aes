`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oo3lkQeSpmmopxDYixm/rspGpKUIHmQ+g2MerAKQPcasgFjIXxekEdlpouYwiW4C
kNWEmqYX95vAp1YowhOj3S3NEyWp67dLMmm9XN8gzmo6IZWAm81/HTuApCaPgjKG
fo0ldeCbAchOwH6UVqbSX0Of/TCGw+4Mk+Oy2GR8CxTYk5g8+jfmxQB32lJq99rC
k8qY6AlVq0dPxJU1XFHjxFz505OgBEOxcnDbGu/M2bKn5kBHLzHqP7m9qY1cdvnu
o9A0OjzMtHERLoKXS0TteSEoxXuCzDljUOCAoAVL2FS8/S4rPjn34QV4t/E6a4Mg
SRzALqB9BW+BWNtIUdh2mg==
`protect END_PROTECTED
