`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B3f2/Tc54yjax7ruWE7pN5qmae0P3/PLZo9l7ZhO9V8hfEWT/LdZxEMpdFK5Cd+f
Y6r6ObWDWqkpc/T6YP3mfm+Oepgb2OOkhXe6bIe1fBfynQsWrlYF/ZKLytRYXUXl
BxOBNx9alQvfLGla2aFHfymmggJGyIbsYSjjPbU1JyyokfT60KkQTzfvNnDKVh7+
vYNr61dvuu7HN5lDSheCsS5h5aBjozt08FnDIs0yQKO9pQLyQn/gWCCgBAQcddoJ
waFk4HUM3UeIU5lp/ztEgdWFZrNCTtg/ROQkDIEkGejfp426GArrL+DlgAtvNAK5
P7yBtGkDjUM6yUJ7XhUGyC2EYvfc6evOLNvvOrCJAg0hVqVBtMQWlS3om2v50X8D
dQBgiLuGfNKRuA5LJ7+jomSdCNd/KrJ1ZOGHvNot1arEnptX5mEeeXYR/5mTqgqQ
N0Ba98ZzPQYSOtY+ypWnOuylOuSIrS2U/4MXHmk4GzTOyrCxspANydmVmn3wrxlE
+ZVxfdoxaZx7wMH5sLtNQMVgFUjgzyYjKsuV0dZiGsySml6fXm3avhOVGPNTuBUA
uVbCWQWb3GX7TQYjKsOS2eXR5rNV36Vy4AS+G3VkmdMwBM4FauVaj4PEVOadPe2r
AqXWkcRwSnVuAj1bSLJbzqi06grblXBcloNAeQtc+6JMWzCIxwIh8BMeSnFCTXeS
u5aWY+LZSjZxQ/n3yeP6CSyjblXnPn1ncM0ogs5+XSagYeC8DUWCm6o3ywyQSnns
qcUJdI7qbKZHhEICjF1G8MQfDuh/ajrv+flchYBv6XnejPfljN8YWhu+8A7uJ7dd
zuO2JMR24ENQBWd0qKb8lMY+K7UToCk38vHPCWYTb4YBdRXT+NUqYndEdTl2BEw3
U4DTkgz4JCTLYvVjIweqmykD/hi5Cvdh3OGzPwZ+4l3uLE+5Hyk9H6RvuHTZkupW
pxuYR6XhHRKbR6BrDMhd30BnxqhjrBUNbk/IjqP4Xnfr8QqEs9KL5qvfXe4phkdO
FdSPlr+sgNARNbBOh9Env3YnUxXNIAu1a6w1C+pjYEJyCyc+yuxMRyqyme4bIUX9
GJx/KsUx9rvNDU9g3SxGeywzcBEK1bMJqralbD8isBDlHFb8Mv0xZ19LSlFSG/+F
Z+hezYp4nKLMFpTkf6w6s1HocHCX10UGlEo3zCReRLk=
`protect END_PROTECTED
