`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pQo11RrtoZfe0Gm1Td1SreO2Qg9rYepPXgc32JYFdWNKtlFTNkxvx2vm6A3VnbwQ
j7Iv3pSLxkE42fe3/800kILTIX5ASOubJS6wRQX+S4Kthj49ew3euABRELXzHBlQ
Upa0aFTpspRtM/AeBFJ/XoCvRkRfixUnBec/r+h+bVEBJgxIk3IefMgIoZmVleC5
9+tclKlYabgIy60kHKSpa5CQskTBZz1hkz54wP17ulX+U4fiLR8s6br7KYz9/Y5s
1X51xXSpUdlCGpSCkbSfJysReZFUmPqnrXTgDzZ1lIE=
`protect END_PROTECTED
