`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IRkUF6Crf7VIlsL7g1YTYZVlOmR6f9cewNYVe+9ivr6SuKypTNP4gvGY91MXh0em
wYyF5V3RS8BpRvy9Lu3vUrnVsU2tTNlTuLzhjuVxTWXXrnCCQallatz6J8CTkUtt
DUmnAsjq1OHsOEgUQkoFnWmC/EdTyijRItb67+FrO+I+s6UbTg3DCHjy3tk1Qszu
scvNdk0422SrqaSR0Flp+fTj0mf5QcexcSNLDKK/B8Cok0xI3xaqSG8XbQpwcD/U
i4E+7+bt14pFWXSEoKUmnnnaf4zltrS8Z3tUYFkjZjoOfljmzW2oWm5HN3Ys7wp2
J8y6b+g3jy2Ifd6/0ir2ueWj83yHJeDDRio7Jbs5H9asVe9d59DdGd8yU2wvPZBI
`protect END_PROTECTED
