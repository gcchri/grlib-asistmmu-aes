`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tB043A5Gg/zR+eLU3egiwwEHCa6lfIU7TRyyt7lFSJ2h6TAFKiXQUlCDO3hlmQjq
whoh0E2dDyA8rqBH+lkEaUq3FFMJWeJEXuRpD3ynJwIESSShhkJ15e0m8GXfpEVX
JLQF0UUlShZS0NESUeIjy4roKtv+JGLnxWU0F5Pa5weFZBhvhSv1FraIRVPWoKbK
NTc5bTtEXq/cHKZ1LFi+lSz9aCbMcuVm2Otpdlawe3sJElkRus2bEMZ1elLRQ2h5
b6nQTZNj8o0y2eNxYMYih3M6NyDCEZ6GhFXYDqTfGun1YXi++aOmdrrEO9sOLuJX
K/Lud3cgW1ZHmMBep4B71IXfh8P1879l+7UsfURquz7auY6+yW+MbvOmfShewUhG
kHYmssugVNZrIs/f+7r2SsqsFy4mfByDWpSuWshAetq8LxzMXZ+KeovniIvKkOtu
+v10CRxd3kNGR10qG81B3k8BAPv62E5uoLfmD2GGHkN7GhPMzrCSGXWIYnZR+QsN
1ZVUgGGIswGP9t7eO0V0xaIK+6RPu4amgspE3g7AJZfjE9Y2JEV+cqpjb7DwbFXy
4PoIA8nR6lrCUebRjHVumgDW6zbg3s0HBvM4XApw/lvL1tEYoWNF034wmxbdK2JA
FvUFp61Nk1cHw6YkAMUYYO1bHQjO6CxphJE0o7z9Ge7VU+yrBKiCdkfXt291e7mt
OYETWL67PiM/dsjdRmlQYluBZymuL5jTbj2/eko9KfJNTQfdkHllBzmowwg+BzLN
DMayU/BxXjqIrga1HohDCvCaL3EiXFnO1oRn72TZBrDvP4HjyJfTglc8DedqWzZH
0Kk2+vafWYheWj0ZOGV+QNlHuo8U02pNHExy6uD9muMMzfCXlg79Fk85j1rkftom
XItDcfnfrDsuCBFppK7ZQaNCGHxzcQEZAY76+jstqfMc0IZV0pfZgflUEvq5WQZH
y0WC9AohwdzL3J/D5XcUwxDfDphi9x2/kmpAhEKSBoUn5Wju+dh51HjOb24wHtBE
Pw+Q5gLwdVrXfynY520E4/o6DYNrgRkzhi5tSHmBE0+vmhTy541KmsQNbx17EtPb
fy0jiayn4kfJgacPM4FZ40qmNW2rCeQs7Nu3kcLgZZNbWtBu2Hm1tyoQwvel2Gad
9GZFHSjr+OmcaE6mJZHDvcwIGG0VQsNy+cC0h7dovAG6OUa/b9HVum26qALSe1xE
iGz2KUy+HCEWH77ejHuYvcqAx8RUx3uEU9+rV7ydUpef/KYfLCMqW4LdWtDpuuhw
16YKVT8olLPkA24eKcxvay3XSDESv9VYIAMPyDy+73/Ibr+X0mo8urPMYC81w8UX
iNQJESwggAdnFZoZpPuK2wHbODcW65Vl675WGdxk8acvNTiq+hufeTWN7rSyI05z
f9sx8hef8zEttfvVKR+vhNJ37zqUh2ZXWLejqwOioHH7zIIbYz9V9jt3fAznTKFL
j1MDopQb96q5ruYrMYVFPenynxM617zoWCKQz+52T8/a+wqo6aGI932ZzhUpLidU
ay6poqx+qVRJL0AUGJjq2SFsjkc+smm/mPL13lIUaYEtiSnljVP35KhZwxYKqwK+
rBjyA7pfLI9xJTBW7V/Itro8wL3tY0+0eo40JZWzola1e3G/1MQUxwfydkc1Hef1
96SVSU2x4e2isNBYdIvkkS3OAHVsv8YSiDD5pDqWyMJ14cx856dvHglzX2jsPIB3
gnMc0SDbO/zAdNxpRXNoIa2xFMgWZMOqPb2YD3dCqOp2JaQGJnvtV2FBGOsYvkmv
WlZ6IYrzePw9TCKbtbJDyXSGxw4B+LJhJ05JYHgweCTQXfPbMmVhOuy/VxHhjMw1
YcOruQBXy3eWn87nxYSs5uKGuQ/1G9O2u9DYWXL158XqwppKGecVlGJx2rEAjwUz
fNiwxGuytSs/K44O79B0B8HFcAU2aQzwJrkpBPW5bPYiTUcATFm//SQuwZw/fLjt
0XDbrbOdcgACa7X3oG6rMN0x2RIMt2fSJnUIMNySYIQmYDGBhzUw4G02wogs+8JS
lQ2yJWEnUkvfksWHqu9CVCL1RVM5KN7t0KSzz79eFbVFqTzckFlWI8uOC7NREaIT
AsXpwe9eIhbGIgJ3/bZqakpbaXbj4reJXjYpY0frWpkqR38Qc2PXWJ1bnxF353l6
ApbbF0rSEPkUC0Qc2rpNWBD0G/XNUjjWmQ6Ch2YgQAFSgyOgvLpaQ+QlJGxTLlV0
miMWKEGCzulH9Bu2RPXfh89hzPkcCyCLQRHs8iCTBDafSEOGHVcr4yZUwfT4mekp
IBnkspsAB1DHftvO+frAZxUSxltgSB3JCM1Wmi+Y3jvhfeEGckGrkKSrEs/BjHhq
hq5L2naoHK6MnX9bqpp5NR4Q+6+IQXR96BJK8GSFPHbq8KXKgjUWU7Ff1sxw2oRO
lu4p9JX02jWAiF7yqNg1GI0mv3vuM8g0KXu3tmFXwA+5+GZrOZZfvzCwFjm01eWu
ZgTEcf7q4JTZOfApiOtOrp3VaxfzgnqkfOB3up0NL5yGr8nEanqW+QO218FmWS6H
ABvkzv6Dzbic5DC1+iZzFmsEJi46LZUgwn8zqQmGpiNfSKtxfUI2TetTt+fF41ja
qmf8OvInw/m9IP414MHf3+ewRhX/kJV1jbAvF3iCedge7s3gJVK15mXhdeCwpgRn
gRCPcE81B/qlQhQykO4fMGTkB9ymGrkCxIL+MJNYGnNDVzARGA8aMNjMVEMX0req
qUbBKjw91NqW3pE4pzoDBqt3QmzRImY8KhuDLd7aFIpFL+zUzFT0Sf9qVpvpxsdb
xhQ+m0Fnl9NuqAtZLetTVrbaOIdyrLbtcJfA7UKIzvhPiAL0OuUAxaJmDWYTrZlb
fJLgA+kveFWaZZHpqMTg3Ko6JoBDZ6JgLPXTobbWlQKrZXG+qqER9MaHoN99ed3m
ZMp37Z2RXtdPDrZvIxd+oZRpnW3hZTcd9K23wzuZ+tMTasJKsY5eaIhvNhu9kYt1
CBFaJxrE22zh/rzVc7xjYbDb3GEJcZVRBXDnP4wMGusJBJVeq+iVXP/mr/3zrlbZ
3owoS5dsAvhcpmia/zAKsbMfnrMxKYosx5wcVBwsXvT1DBoJtAZuql1H8c5bvaqB
tsEi546eoIWnl/7oaxSAT9fi8jeQfDro3/BpMi1k7w/Gn5c9ZEDTt8LOFaJ2O9lD
K+2R5SQG8wxSYkIKSFznwI7QFSMJZNjSOUr4lr29uN8URTpV+1Sah63rwlnmIJ/N
PfsTDnWWiRpMiyP05aNe5EetNloLou0GPulcfFKa8MdWTusuD4VHx9zO+0R7ZDKP
sDZQ0fKodLjmHIw7CqtldxVzgMLTDNzMk8yJAgAWymE1oQAPEGf4+yp2W3QUypvl
FqImW63Dv1T/D8Jyqt/81FFOi7fRr+HJrfpQCAGvfGDzuHoc/1Snhapeqwm4Ru39
phH376T178qZ6NXRf4aY0I0zMuoS9qVoMWG8mzIp92k3ZM9JA6pgDqhyah4z6eiP
lLuixyOzmtLCE/pJ1Wm52ZdSVe2eRvohroGJL1rPhm2ijMrE/+Fx7SEUzHnew8Ba
hgdfXYr5IyyyROGzCIKXFP5iFY+VNsbdTsl/DOFPFk7uGTow+Nrf7d1XidU3AaGA
eRYTc/Sv2F6p6Hc4d6M7WScOa/VxnDnTA+5Q5HOCjJny9cP3o8cb1vEjuWxOx1PA
ofcP6Cycz5KeTF3Kxi/+9wxfQyPOp+Q+USDK+0XhgBD9QyL50kwd8HnaWUXw8TmN
malVt4v1av54PA1P6T1zpdgqI8FXyJ3q6wgNhD8akob+xFGoFh+JdmzY5uEyxaAY
IcHPc7essnT4S41djG3BD9BSug/0NL/m5yFSHsvsnPBaoC7he1yc81D3Rmjwwa4c
PuSeMeSL7/+AcOHvuChdKA1hrP55WaOmDNMf0dO7sc1jD4vAeKFchV7ExCjfjXE9
5zzVLQyb8PlxRlR/FNEq3XBPc0I9RfBM7tjdoeOqdvO0W4oOrvDyDTcmSVBFycbI
XDJf0eq1qbnC3hpOAyz882FQCdP6IuShFg32HzU+Z3Vl8cB1Wc2AIJUFZkQktrTs
xAXivCjLdOpG9Bd2eZgVs8AK6/ky4qdNT0+1fpE6sNvEMLZcUb4XUo1jqzd3F99q
cFbT+s07+qqXvrdGj6YdqkxeA0WVDZUT7J4J8V3YpBmbeBQx0D7u1sHhbLnjnJ56
eK4sZn+APcoEY6LAkx79K9HtISKAotrKxxRGEDkQ5z1UQStPPI9hD+JBerxuRayx
aYAhUXp52ywruhR1eB/nwjmrSvOvhjEO6w9Ugl2enUxLRXiGWvSEMLpJTpwcGQ31
Ozrw0VyBNNNG/Z6j6peah4y0eICBr2aC3oPingHvqXpNkaVSdjQ4fgLYF7VKd2mY
sT6m+uz1FpJ8rQ0J+AJjFwiRzUmQscDpZF55jKnoOHrguffLNKfdfVKKm+IauEMI
8KSmbBDzuQBaN3yW/9Dkn6MOBaxlKJSg8w0yg4UDbBvh3oeGzU8R6BFngFmz+9M8
V1L1PrVD3cglHxwFxVFOaKxuPOmoe0BH9B0T2PGSJxN0ndPkiKtko5ezkeDFGeG3
nrPDwcXzsFikuxykObZ+eYtbrDrsZWwFfmTA2Fp6ersilhXa9ZGre/fc8dnuDTl9
Bc7DdY0Pl5Ru0VdYdyNfLFXDM5IeGLmE6N+mPhz0bEQ1bvnIMTHHgX4bv/+hLrUC
BmgNNkmsZ4X8T0Ym0pChFWFLnsztAo/OWynUESEsqjHoX/Ccdo9TgvqJKVcdoFth
shc4odOoRq8/1ybp95Lehf4t0JMaJ2G/hbuY7JlkgPTt5Pgb7PlkEXjaMZ0kKps2
ZQDYGRBgyOBLNUNwzOvS/MhPulZIhOBuTOfUtgl2ySZgE6yhn8zRzfst76Vbbt4F
qEGXsR5zScJcBE8MH61L18BDeZmGxI5lpcm2uHJp/mazfE4fxRqwpqeF2qfa7y47
tvNYYBuji56zA3QJWPEPw1baJT+bjiwg8BhlgAA4Svlu6htThvZn8cQqRaWMuIzY
GeR7Vzr/O4NiHdEABHQwbn6RyV1S430tztLAB9HywsIzvxwVaUJ+aWRWBEzXz4O8
DgOBXb3J40udgDjMiGgmymdYIXNelvf1MuCJD3BOXAuoLyFfc5PzSQtx9kn4vs+Y
Pr74AW8DZ13qe0fmltNSO1ImRn8ljWFCx+m8h9vBbsVuZ6DJWoiwZ0UAHwh2dzXB
akn+ZQjmx6iS+ERp59QjpUQKF1zFGyVS3azCjzhkW65w9/fjSbKWImaNk8EAxPr/
mWIj0vbZsymgu/m57a7HTZ84dF4SBMF3pKUfL9r/cNsWZlIqGzNAYqnu17pZsq20
kWdFysBaLREVPRnbZsAHAbjOMDDD/Noc4y5kXuPIg1Sapr1FLjbivVZEJq442Mmv
Ek4Q1N8XeLnXDSSKxKILGAU6XTKFceO+befTRiegEQyf78MhAkixTZ0mX17VDixI
5HVSM2p2zpXbltKacAiGQfobNctZoaiW51N59UuwJWKjeEj4S29snyJ3ZeTS8Yk8
t7RK6bJDQAloRRlL0YMM4pWnTxmzgthWrWQFtO5nqCeMu80QpBHTi5m9NIG33xNb
383kdTpLIEgwKBpeB1WcBNaVUFCYcAammpIYCRx9rDQ7jihFpj++pUrOp3H24m5U
E77fV6mXwo28847f645s79bbg23Ljf05rGXC0iCIhkzCc7TUNMIdJKkiP/+B9C4x
GG6oxsVA4S9e1WmERL8WlD/N4EqWoFIPL17hurRwhKKvdcBxVImZjmR126G/2bDk
4ul82QAOghPMweBGnNvTpC4cwdJDbglch7Kjg05fq50K4Z1PyEsxWTb0VzJVpeNT
JFcDslFwemB26JPWbTrXJmG+iSL8+QatuNfXg8s/FXtUNSPtkU/Jqlx2W77EUIUT
0gkHlYFoYWfveXEbO/OY/2gX+7a+RRgDNLtX3RtbSdo0jwganHx6DHSRT9PMNxhR
hasvG8S2D/qXzY7ohOfVmcv34F42dhgr+4PHObQJb53f0ERgLK54hg64bwihTHpW
WDrZBagYtaccmMextMQ1sE7tTvZqwJcRmDC39MkVFt3J6hxuMPO6+KVDVuyoaqRu
0SF49xXPezJ7dCxEbJacWueXFaAXbyKBmsevlzw/74K3vcKU7fecKlwxdIumYMxv
PL5ULwgFoVIKY6L7+k5IYtH9x/BhxhXZgW+zOFG7ki/d4zW2dIYyuKQSocLO9mVp
6ensSP26ELwOq6rRT/gbmfk2sjbcygXZrMHscD/OXnVXqm/leJ5E6IsHv3uxE/Tn
LC4Ed4js8vRBZ1Yuwax7sxMi3Us8CR3OpCTbRuUvydVrMysrdKMkid6qTPXLfmhB
NpMQWJOXDfvW33pDO4WOw5fJ5rPVAumBg91y+O9SL5PJ6NlTOltR4xbyOw1G+Wvj
I33ZNhlNp2e8MIS1wVW7oJfXYvOWp52kHdIDsrEYQwLd+bi/q+wB67juj1lznyHn
KOF/anfNY3ROqu71A3NB73kwQpruocgXZCEfbQ813J36UTj+K1UCrm+27UtUpSx6
BB5AxknM+av6f/LadWhnN3D0RBd302kNQxfxKNLbueqKoYNHjnWxn3FqawF5dPQ5
CiDfkbv5tAcRp1Q05l8NJWXzRe57eC1vE1fGdn3srSWb2rIBKcSRWNtWt2BfmDfh
EihF+wJRmbSsOffAlw9ushK8zGUlEhlA3cto9xwCzpWFEDivnGtGPWo33MCpd11e
lfsivEPWP+Q3dNtwzl52bedx23p52MznWZgjj7hbfeehv3BPBmJkwxw2A2mfgshY
lcGiNeeaMFLOuvfqKMKqzv5tS4bviJTXQKph1tlddKR+F9UK/ur3bJiyZwYlZmlu
ogMeYvPEs7HokcxvvWixUS2vav/ITspA9kWGYEYhRGseiyS/LkR5ErFcrsTtqiFh
pJFTokeXYJpznO3EZoTZoCZdXl0kFaTFNOroTnwF/hr37bGA3AU5i4PqLYARwcHH
LBfHxqw/rYdQjKA/W9hVc0xFpUOmm5nELi0Gc2W4XiDeq0n+lFsHGFu7taSyA9wQ
yDK3HR+JnSuTLNmJjyaFKc/UCft4VEVG5bQHNIGoVuUFyItSnz8vXeY2W1r2tMl4
bKldSJbCO7uEi+s/6U8/Wtq3cCP2BEW+RmGK/qny7/HozWH1keOWdv5QF1nNNPmP
V0sHJsACvKg9tjAK71rvyuLIYL2Gh5mlGvRkrGKRD4+bgWM7ihx4q3H+MaJuwoIC
qO1dHUnBDLYptlb/7dJ4fbARB5/IZ/9bSYMMOCQ+0DGIaFor8WnvgZCZxBMsSoUL
FSRnSz5OfTX+bKp0//21lnrSBu9BlWoLuqHSn/s3MiPvuZldbsJ1VFjFZM8lNxXN
a6MV/uaeJ7/b/W/xVFWehGo7jB7bK/gzGVBC8xCVcRF6fT0toWOMgyCDls8z7Y9m
1gevEWKAcT/xsN6A+o2yxpeYPmrIFF1oiE7+Voa+9njxYc0X98C4pJ5ZBPqXSCwm
SGuA1n3dUP1JGSa8jQ+1CNyDcNffgc/6ZH9qi6UmCepwD+H9ZtihvUkHnKsP144z
gDcIvrPHIBVbl8A1KfKY6IxQY1P5REv5C52AzbmgJicXh6ke5yTFG76rgY5lrqxR
t/FD1U6BvlxWqUxPHG0FLUpoVAluygMxNPGtLrJBBKqSJHE+22ZAbHyjSjpbGOC7
1hDNzrDj7XVQICnAbI2nE1s2marviVRxrK7kqVx562JgmRaHXdTag9doIrgS8IIL
9chnn15SyOCBP9VGJADB2ye4nzlleotImTcA2J+MOV29XO42oO834+ENbkQx07wj
V3HbOJDQaEc8n0pC/a5XFb8Qq4WTpEXCpSWZ1XYMPX1Pzu7t34aOuT7hxlO4lhM4
xbmw+pTCdnLEQ8Oxp3nFLRVdL1gCMys4hdk4aAiLemS+9x1rF70UZL5Kq9ClIQIr
OD4+jDc4lNe46k2OaJpLothsHmykBCcTewh8X4Dd+dem9GOrq1dKQFf2vogElAyA
Sq3A6rj84iAZY1JQAODLfUFqJwt9bsh5qVelKbUfmq/wWFLP06xC0KP2wnNlY+ws
Vwlq6en5bnisj7X57Qs8dL4wTguBn17Ym34lVw6sZfpPq1lkFqGNdGySXIHeAI6+
/fXqJNZwlSP52XSfcEUYh/qlgxVJERqjMsBYOrTLn2E+D/jactm5B2csALLxwCZM
fqD2NS1Qu9r93fo0jpOt2pKdcKURTVWz5r49NxRNoJ/h+Ktr5xtyVzFRv8YBpxMC
wOwDnIojgHrs2Z/E3LP/gV3FjgyL79SL1Ca7t0Ursp+DJ39emQKSq/VGSA2uUJMu
iArzvOkSE1S59Ynkd2NYcAKe86BdHXqTIsmi806LQ6RO5dLK+Wy33ti4F5JxqsQW
W3r3ZD+ewfM/VN2Qoimty6pSBCeg8jiJ15wckwkrSSXQAyEmdrh6EUtTLY9XEBoS
r1+IU6dv/baBd//6dA/OYic2U2eDqP0sDI6l19UuirU70kgGp7ygMvYcgyBUYEPm
WcRd2dOl8nJwLUJ7/NTO/d9su2TKZgrpS6od+o0FpqXKxWNwBzbUq+YmtHvxk9sA
UXfAdagWxw6Yvqlsmom8EhkC5j9pv0mbG9reef3mKgp+0drA+kq4pjDF4NuQSeUQ
m6LVgTdaT6HWyo7DuTJPv7ZTi+3q9mUjwuQVd/eNktjnC7COFgoWs6/mPhogR95C
HEZJoCzZ9wmu1LLoCPUWoxGPDI6DLclpAxhzHybF9BByyXb3EIv6zULGVrX7lHt6
ysj+sXTA32aL0uvxsMUc9ySPCb+p5E6hgxGstSYHZq07xdA0UsDRyzfePbszDPcb
F0+kUZiEmIa3/2AUJsXnvzsQlqq7yoBEldKbb+WBCKvkVPcz+lk1QHLsIC689Czw
+N3+z6sLphaIuvBs2tJWaJs8l1frQ18LeEMmcMlRfgyTldz0iFtnnLFVobHONZ7Q
lu80MP8z3oVQnUrHHot9kkj5CCmSEMeaGNdO+w5+yNKbX4NDH7AW8bFoPgLQaqvC
DLxv9SG6Wh/keyjsvLrSr+xPuoO+xtRWQJk8E5IZvwxjnhkSRLrijhwB+LCXNQ8u
agPrDX2YO4G9lJVaO+qpAqJI0AC00fOvnEiued8TB2xhDhn7EiWre4/AU6/VgWDK
mph81TcehAA2ln5TQXIH7Uelz76/rf3tL0/ITa8EpDh9WrEuxy27b9j7pO0kuIHN
RyvIqUoZGlZqK19oKu45IPAievSoiUtZ24KjNdEvBL3/DrQEjXpkGsRJUNPEyIYD
5nRpFGponFPgssX1YdPjlRsojryC05kJ/5ABv+2P5PBOanN65DaqI/Ex+RCbBGYL
pyvedXeMTZVjXKVLSXdPZFPlG+e7WIjrLjzbpG3EGT3shF+f9QIPiKXoaOnE0qa2
SdT2RoxIRrtA3Mab6cOfTi0SweCW4gl96g79lf/UOye1S+vrCkYt7pOopVXinf/A
d3Eh/th2U7OhaFrXMjNvWGn6hkFV/sgiCUrZMagrmWbVVCeUfE7iQABal241Vl6s
uKdfjbZjcN79WP3hgSxqwano/wR5OVHaR7n9A0BiTDJ8bdaPDHtiQfMd/aTVYp+1
w+sL4HdDjPj3EwfpAmVIn5RThgwbWQR98nUHKV2YKVOdzreOCGB5KPXQYJANFe7E
oQglpV2MxwtojljVVhyREsGRb/hYv6KDHOf6p8dxwZwgtYc34lKIcO3dpTdR80i1
xQnAqt/Y3F9r1P7ZoeYHqrqWkGfB7NOx7RpUE5lLIqgvuPFPi6U9gCL8xQ3N5nYo
nAeiQ9jP82m+q6CRWE0yn7el2B2KwjcS2izeD18jTiYWOOQv/y17o7mnby2oKmOo
mC0F/QeM/CenZIMYGa7q7KKMb/GjDW4Xn1PACUjRYqPgRuIt25MQjUVCI5KI2RU6
3eraI27BGBKm61bOZtfksVM3p1wHfIU4gC/Nv3b2Z1wgBrPWZvREVc2NYamRNRci
3fWI5sj2tOcFuk6cbifzoHHZ52+YMVzwxtu+Z+wvsx/1CPbw5WbcBlh423yWNaEk
GeQD5et2JuBJmUGn7ZkRzAANx/t+WgVY/sqoNste1dv7j5Za/9acRBl4VOIdNEMY
+7cOfl+pxoh0/iTi2fVCCIGnqB8CJ/Dm8acfsCcJuYCO12nC+EfFHSBDFHRl9pwl
NHd9rjQitRsBFS/ZVliTJSmsH8Uc3Gp6zGtm+PpYYECO2OXJae8tVxLunJrmSDRl
jTN8aw9CC4TYmwQzVhQWWqPX/6G7EuNuQWrAxD0geU4VJhEEFVvNuZ5ciOszSoGg
768hABXtQ5l0aBUjayoNnhy3EIm607tRawxelk66yYPqijYkL0qFDgocKHCZhcwB
7C5r3Wc0UhltlQSAFeEZONThwROwxUgfje7gHBvJX5zxj8zgjn4ueIQpbfVDlIk1
wQBmgYUofvUztya9cj4MxysfIvLHsJPWzmvo2m2qoPZEhM4ME1nMXte+OP+POtxr
bCaVbVw5zsncx7P3v30ZuMuY4pB91zDsmvnoMSlhEXHt3+c1jIbSqm/eC50I2b0M
CAPobTKTdTdX1m+fJKQhwOreXiTBxUweFt4JrFPq+l+arPjtKQAV9f+XK6BwCmHi
2gUgjOv4MfYMLMxoVHFEXCAn7paf/OSYHO8dpsewmeGhTQsTfbvrK2efy/JtIJ08
ccCyy1NwQwmPrExCNnfutHFPrwyHm6xEjvr7FmE10BtMkNz/CScpT9IEPLG+RrtU
Jn8VbERy2H14Utv9nhVmSC53uu/zLO2zad5VjxU+kYYfNP6riJWx/S/ZAllOW8PD
V/KuRcG4ihD06RjtjtTtk35F/0iPo5GMcfKbhuAsdRbn3ndYpgxMgDp+pRjJvPci
0DMdULazY1b7KheCytNdcNqOXfZVpoDLUsU1nr9fgfuaF3IXnnMFLOUBTwMdzHCa
TUiZUIBVbZAIFaUjZaDr/mQRjc1na+8zEMZjiXxiH1zeWINUbsVNBpNmpqhG/+9b
QujwuU6CcLRf2wzxslScQNveDjEYO3FeIhi62BhKWcCRZKID+g1rLlSZEdDnGpot
iHOk8QyE3JBoZkEz099u/PV/k9C63+0kFU222v64BpJj5BRYuYRi1lIZkwSoQaxu
7ix6eh1qFMv5YTl0BM4B4sE9CjLzZ8Ulk92mc0OVe7No5DunFS0qqML5K2fPEMGN
Nr76eCUqv9Bhd031+6mfP50LhiYn2jEJbDr0f69NrMbnUfmr9L1EVs12AlYo1vjT
gWYeiN/M35fRs7Jmsou6BvlDbcPpj3fTZVXyD+ADarlNsX7EZnayzKhTDzmEV+0K
dq3qofKStGMPbg9pRm0jiDx6Nlf353HXplIvN/pxWutks0crcEANS3dxRjZUUwJ+
XvdcK2I7I+givO5Sfbo0NT6W9lWvNzZ0BeKxxcjNUIqrtJnjuHw91zFDXXApLRF+
cuWI4Mp47IklHFgzsaprjqF6yO1LdREYjP9UF7tGPlHRuAc248VcKCpQCyyAgkZ/
vz7iZ9iNxJz5y1sQPUlfS01H0ILlSfm1zg2+tLH8IZoXI6skG2Apz1UuRxJMkrmj
ohhlbvA+hjCyJVxUUQz30uJJUI0232hfJXlGEWa62Hp1SAyxNdB7PlFXMafcO/Tk
5J1IbYeT+lE+F3IURDSnZeJON8VZRPdHoxzUl3AtP4hKWR9IKvc0VeXtwIj6QJLR
cOrCEiV6vmAAw0zedt3wmgIMCPppxfbXBONxNNw+RpjxqTCz3e8a5xRHkYTyWMSw
+iAlyCZ36LP1TMAaCBfjiAnJBxF9f/xcxwS+ldOcIBcARdu/PYReXBcQHAyyzPi7
VCUX8050bTCTUPt2iJMdyuTgewhLkv6Kux71jXK/I+TCzLvI9wI/kXPEQSQV/P8j
nF4E3KESyzvSHFCaxswoPzeYMLiUNT2yUP1Qc/SQeOAGu7x54rk5796Ic4dYu6Rq
/xtLlU81I9IgV52unYz4uurYWH7+E6gxQDbIIe8Yvc+caec2Hk/pN0goW1Sro34y
QxFfGYHDITKnPkSNfLoKrY9Rbja4m+eB/Dp0nPMI7E+3xAg9ayZ8u+gvqQmk/3I4
kMCc+SI2wjbGYjEEvXWwnLN4Qkr70ae+WQbD/1mB9qkOIfIyneHNGUSGeaEl7h9R
GYuErHMlKlbZb1BioGIFva3oLPclGNiq0MRtMVQpvo6cNogkDEzolyrnUQob5MWG
4ZZh5BT9/CDPcqkcvW4wOdaapci1ndxhXeNmIDjQLzVQPFoT5AFeQpmbh9jX873a
ca0k3qLVBik7dGHbk9CTdYSHY6aWVXW7S6HE2p+gMAgxBpju9K5QNxPk/7ET2TSw
8zvdXYjzRO5sQrqw5BeiPryWtUPTpC/mp1Q32VTRT07dknT63RyIbeqqJKIXhDCL
QbjE/tl70VmONTcgtxF/0CjDNfPIa29xmG+9Mqh1sGQ6G/yK6SFdM1IpqRyDIWFd
0yTg9WnxrXItgDtHMVY5PK49p5B9CgvbAwo7C/SpLkAx1HTED2Xi7i61mHSd8lMD
UXdCL2k8OTI9DEP3P3BeTbXgJJcs0nUuSfycu0A+7rzYd19jA0oG6dxNNjEa2Vnr
LVegIoAydCDvCNHNeRUob0rW/1rHvt6qr4dL4MTOXcbn+tMhGpnY84sP+iyRjkud
BbsEB1tAvo+NMcSrLWKthhsBIUJqAHCxswiapqrTL/0ziw4/vO8mvhg25GRxdYY9
x+vgozG7zONs4y0MeJRdE9EgyrnFMxV2Y2Kqc7zRFhGCA4IoMxhX7eAH/cz8pQJy
65Qu5jeKUCdeiB9lZ98E04/CYeJyQwJCffe1wHgJMfBQqoW5K7Ld8viskSK2iNyD
2iGOvTjMl9YMZGtyEBP02xPFbZdoyVJ3XvqbidpXQx4hhQKDbzmxvqnaaREYSmxq
+MLayCKoiWFgSbTRc1uLEVeCgXgcJdnUjbJzePkR4fjWvpDPE8gQ5h8FBj0iTNAP
L/scjQQSmF1co6punfsu5Pjujsen0jngHC85HZaWDJ6IX9fqYa743xgmrEdfY41v
/pIJKK3bo4vnTi0K0jgxHg+8BPOEutsxA198DkzU0/m+wOAVT43QhgWqv6UU/P8L
hOSn4EYnS7HylLE5qzzqgr3lBAgiRs3PP/9n91o7XNFwmL6NOQDDftGoQgX8cPBm
7ZswpcSyR8Ur/uAwKofcbq4S66aFHsAdg02jCLVWg2Hp1QANJUjpMagw1cj1cHJO
Lkbx9BMuIAhUYFgIsixzN6M/D48S67+JqitKSvGWNv6B1Dn3iSDWwohEVGWCyeuq
jhEwxAAQOif+kHwkngvNp1bxrenfisnIhNQ+8W/K+lfDyLhk2jut668b3ENrOYIV
qGlbZNtwlQZdXTx3k/0oKr8WmxHaKbkMp+gPGdUCdXMkoUkwNqG0GGxdSqele6hF
Sif1jDneLuYXajSzHZ7ujNPCT8l2GVVbqEyWC943eoWAtyee5YNx+PpnXQAgCrUz
ym6VK6+54oQGX6ebyRGNoB1nIYc/r1EqadZvb5yigUupz9onUk4X8302DEBDKTcb
k4p7I/Ynw61QSkG9K1YbWe2TMA9yHr20+U1vO713smLxA7xg1J1h+7TGVTTuMqon
V97RrqXTycVJ+lSJFDdOrUnHetdKja7CvtrCOmiqH1DDfHlLdcxDYNIBjL2wqdDd
yiiUqVu1j2xTS0x8rMWyRdeENKOOT35yyg7frXMcCaJKA9PbuIzE1uYHJxFhs2/f
ThNaTZjMRcfu2GhoWhGH8MWaySlMij+eQx46X0muqVuQYDWzFGuaS0O/oXA/JJIp
DUaDWLasYhSdn1v1q+PfF080K4jX6dP6yXgvCBJ97Wy1STwrW/BJ8MwIKB9gxehb
NIWfkuNrh+d/KTOQNllnHx2Qw0JECXIHM9gQj5FMYKhLV6H3C9/3BaQQ0sjFs4FN
R1DF8XZmSdUhfm2Va+C9q5+n48RxFVGuY62uTDl7Z0hjY9Bo/ywTt/VUBqgf2brZ
eVE4es3Z8WHPPspD0lZoO7dPrD3ts0Oh395dnwq4JDBaWh0iu7vlRj75PVoeN+dj
Wvwz4XvqFHJV4JukMm7f/R63dNPNrqmd3I+rqkl+AX7WcLAbgSzIas09o1rdEb/4
ER7VoN1q/qtkeOPZ0kNvPMB+y6fSq8CRT8toFOQDeQ7FgZqcsMaBcgvKNzhGMRiF
xn0WN2qD4lTmoi4HZBvCNgHoapV7XkXTvZ3xuV6thHrv3tNLVQfEqNMjVw8tz4hw
3CcrKHc5XbCWvuIZd5TMZbJoAc4dtVBJJkjU35Ht+mcXiLOMyz+fl5eHK3Q/bHMb
C+Oh3djxCEGuV/IKrqHyzzQDWYdFb0hAab/gdjchW6XjMePhG0r5Sf3G0I5Ijisa
fP+e5plR9nR26csTj3dyF+Oz0dQRFs3gtCXwfPw8Dp5AoYeHj6lGcxWWbzPQZtPV
lM6VjoxosJM10LfwPufk0CvUfxJKPfv/lsaJLyKh+4WYyj16ozMaR17zbtLpynKL
VTEmpB/C8QgHI2LyAuNfqdyd3Nm2U0p4/BHTPKVn4o0eh6yaSjZxWBg6reKi6LjE
+Wg0oydHJHFqtGPX/m8f038Fo7CQxDpq+jwDvU3yHa/XQLneB72SfFlMsUFY/Mfk
VtM579F17Db30zKSANSnn6RdWnme2O5t8vwdRghp8071dhr/bNmwkLIHgkgYazkl
ejqNRrQVEYs/Tj/UqUhpjRvzVAD2lBkUGT0V6zAjk6sC1yqHv5r4vnNuYMU159dI
T6mF2GSvSR+KAeand1uYe3YKME8+ZTiHqwCFiaqJAc3yDqEJ1BmqsjgdUEZMxN54
WMnOr+cvriplJzuJ3gLOYe0mWBN8te4XsPifurQexfjlR9hfJOIjW50PYP3+Tj1r
QeRS1maO3e2jzyBBuuIYfRZrpbpyld+mtJBRMOKlPlsA2PQEs2CyGZ/qOc2qVkhc
Hi/weuO5KEqc+2bgakXCXMXqq1iT5IDkCbHUGvU0LYyQB8od8yAgD1rELesnmHWr
eJTnWCfG2QUzjjz/ruUhIe7jq/yY7tzUsESaEzexVomO7Xb+SldD0h5aO6fR9pJ+
cWXvMqcxQlk76wWHff1L0V20CxbPmrWe7JhBjEBLgIism9JpxR30YonzMO6Y9FZ0
yKfolcQP8HWpCMhTGU1Erbkk2TqmNmUAlvoYvteQZ43N16BXwU8j+ds3Qu0CPEtn
v6Uoj7zOeMIqA7wqIo7+2+5eumM7qyL9Wtg+JR+mlkpS2l4IgHKHFnq6zEvpjVdD
GnXHhogwBNlC4AVdcMwjVZJZkSXNTPteOv1eE1ndMg6vJX8CWdWtzLhpU0hG8hEe
096kwuzS5S7FD+DCVycCeLtsrP6+SCAC0Wnnqde0cFdR1vyqkZciLHtZfqwYfQe0
8hftseSeoqV2LkX554TnRkx770F71O9jAZakO6Qtz46dkL/8sKNYvF9Ueng6pz0P
ZQqralf/mvcwGyXxJlFOW0PpGZuxoIEzyL1p7Pz7eyAfN5Bj0/qMd8qbbZJMp2sr
WExkgeigFAua7hcjUGfojMPsRoy5exwoj9vb8Xqwk16fXlcjVeoiMJ6KQxPuU/6U
0PUvJnw5JdLxZ92Lh/S3eJDglmo5TDKqYh9BNYWbY70vkIPRP2uvgb8dxaIJlxBk
cxaT7iaK+LoT8Coq2mR7qveiE1mfikn8R+zPhaZZCfPl7/UfC67C4v6Ho4T1SkNU
nuqxewi3MN0kN+xJUj8EUGDdlaTxaKAgtY9WUcnWv0j26uLM8d3zakRWuDYO3MPj
sYoSED8EKqtHHmXPgzZEr9i6lS3KrHgsj4QsanuMVnun4hhq2yj1RSvycaFAco+G
qMmQDXrDWL8uK8U4CrHGjC8BrkWJdx0i0jHjThW0JTpzl5yI5XxXJrcLrO6AeEgj
IZVPlhWgKfxLBhCWc2LNVi1XyylZTY9SOTDrtJvnJ+RsJTKOnbogKJTvFRCmiBF0
Lea3w+ghZq+YJ5xH/RQ/QVRRg9/RCYKsXmWBjCaDO6vj2VmXxmAM5S6TfMPTszk0
jNuomP0mF8cAhFfjWUHqIAqwDzpf6o1I2rIB9XCFixdVF0goKjDB45kN/5HUi3DS
JXXjMSd/dPC89E6mCZVqVWoVISJNU875c7VaFw7wQaldFOf1rjMzGGXBv+cvqkLB
asWtbw/5amIb5SBRMilibPSYEdEY5pcy2nDloAcAeC0DxWNTeM2RGkGT8IQHy+K/
WnRmfv2taDeL4CitgDfXs9qiGZJ6Bg2fqMgwenvOj+vEUj8F+FiUMxHJaiAzc4ih
RynZ0dx2pbjll2D78KvyvzBxiLRPgwRzSnbOvU23Bq8ThHAFdKa0TYEMS40nRwid
jk9KmAeTYHHjcc48OKp+IQjMDHYOo0ix4s+YVyVe8vvC/jhy8i0fKTsNEBsMLSEN
umPfZnFrsByPR3WjqSc183LX14MmM2CkPjEGvFkAMyBMijsOL3ElSV9SZtG7VkNK
uho8MovsM1WHdiFrUzLGnrLW9dk4FSiLQ0t2e4bMOVHuVJBIdYJwsz8rvMk9/eiW
j0LjCMCw9wZ19jyowHZ9ZF7ffTVj1Q/A1UUjRa4jLKPfDt8Szu7DUSr3grBAjXMT
lfUZ7bPyNOsyXTqkbp0zFf1N4eqcHcDUreGdXqiyNk4eX7V0PqacNzft1DHTcg5W
awkJS/8uyRLGlh8JT0eP1QXQhOkNO4SdSAa2Qyr1221ECozAqNzTS8rt3IvcHvnv
ZXG4Jir6/qJUgHWFqd7g29bctxlSRIbfbJix3RyoaBZxYHlzYjPi5eriDJAYfVIx
E+TkGR4tS4Uz/OYQwhBvtSjEhikr7cAfU+cjkMlIQVri0y4rH+lakcIykPavtcwi
NtrhHhQGqhtB2DBc8APtWrxjjysL8kT5O4bECMeADFp02TAv24NbocfOB1RZDrTz
i4RhJzvUsgM9k0YvGWYtZj7sR6qOfe1kce479KdT/PBh/xVVCPIu73QVpCoiBRaX
YZJ7EmgQAAYBBHB85Hsy1y6Kv+65faU50D9B6A3vv1Mh9K/0r1AR0btjKAmsnRJh
OLmwD6/g7Wtolnvwc0M9ePrgbgPpxtKyCl/3BzL8ILrOU3aMDpmSSLn7Tu/B7JoP
eoTwJQWcTd4IYwX6DkM1hlsdZUP31PmdQD+Cd5buH4l8JRz3KWqnBc82AU/LQsgl
Hy7dCDAv8ij13ZROPY5QMCQY1BWTSew9XmF0t5+aA3lph3/yB0Cpyz3fl0CobHe/
TJNimKMNc8OIlGHBjgmMBEUHScm4yCjhlOFr8XaNomaBPm8Z29xoaDr+UK6ra3rw
n3xB/6vSEPnFS1J4eJ/GklJlP3dGfarZqvkB5KknNUawRnu8V972qrRk2QthN/Qj
4f2vGfyjJGlHgnAmebEkWFg/JXSl4+1HAe5EZaP8Lp3WDWdOjbr2sXQU3eNFnInZ
IUhOsPun5NpgrePhho6/aFfz1otuGI2BjzuHP2tAB+qcsqxi3Tvy9vZUI/hQuviF
OncYiaVCvHmLv1+MF5WaWHbpQr3bGsdj6gam2Fh21gNZXebFVaAa4fl4qiLvV3ax
x2y7OZq58uO4/hhztUxggaupSOTCh4Z7Dgb+pk7TXtQacYaFadWhb+oqgzlLQqWF
Y+zuXiCxanFywkek57gUiMDo+vVAgc8I75BDFdZiWHIaotO5NxRex05l7sOJxfss
ySlm4jK4dE+kXVcc7s4KTGRcts9Er67dilvarpAzz6pQAnSdYrAnX7uZOwvyVxGT
SHG32hpQFP6qH8C+DxUowG6EGdfI+cYyum+Dj1+SHqFTDKr2dpm/rUUXPLDrDJ4E
kJ9h4n5Zto73k6jnLTlXeoXcYN6TMhbqxR2R4KbCmYe3Es78WmGTiELEbDB377V0
0igteB80pVBj8A+mF+yzM6fYmvElXMp2xGK5BU/5++jf0IQx595+giXp4Ab0YY4r
hgS1sb9wHx52k22BZVbagRyxhO023rdYef8cQSzNOKFdeLLiToGdrWuwqAPGdEDM
Dcq75A8MzGZlMv+4/3aETG7/kRcahhzgNUAire7Ii+A2TaJj2sLXYmtY9RveA5o8
Pw22LUC1k1lSSUjdYp9c9rDvftoXPpUTj/X9vGF2czNkW57/I3IXZdlUhQHWo90+
1BH/2UGzf8YWiqGyJuUZFBcJsJQa1AB+hEJ/7dbGiOqjqHlXQU85B3GOWqtUWdN6
N92MFnqsykI5UKOdpFgqqnrIjtI5bWTW/uAIfwvDv4tYeWpFeLsIo5uSq4pjJfbX
XOJqEAFxyGhJDgWtHeoO7ZSdOF3Hh53b5Ib5ESCrfzzBtAViRCjVvTGsKa5wsqLG
aKXtLyqiR9SHCmiP3ibfOCROJfj7QmXH12NWzrHgG44dLTtUoqX6Ckq1df3GU0Yl
H8D35I1bCiYjhdsexme+ZFd6etzCRhVAT/GRv4s5xkzi49hD5KE7Us6bw4pcpxIB
Q6FsWo/2YoHfSi39CVK1/wvakFL8IU1Ak4zjPzksc9htj6E3LLzvxkgdvOfDnEku
1wAxtXIpPTfVw47tpYT6xzWbZ/3cxc9R07HusEdYq5F+vz6WVgF90EPLlYoPvVJY
ggygkbVGF1s7JwwDOJzqWiGZJT7f8IHt3Q+TU3LouE1gFqv48CV4NE7vE2k6ttpQ
L2GxjrGqdebnVL/xFgK9a+3+cYYFXXcnRWWHDjCK4rEZpsrxI9fpStGZEm6puDTB
yHhhsgAH1r5bUTmg3ZGpiGeOt5kxSUb1FwBl0mjEorxHp9DtO7KrP6aohTsUyxqm
1TIjD8JzVwcGQ33BS/rt74eE1bxkejY6DEMkMoYQbdJuYqfdHxhxQRyID0eYHNTY
aiDKPogiVYSjmDSKn1VSTURQJD7HiAGzwOvdk5NbAUm8KjN2q8J7vr1vL7wMvQLJ
CnTg8yY71xPDlc+Ynxmlet+ZNc3a33UaJvj9NSj9fvqeg3DKU0resoyTEd5r7mVN
BBnIxpyyGg1TsY6oCI8twHsPdlwB4vXM1Ztu+FrWP3T7v3+nDIHPGJKZVQ6tHWSf
Nzug/FPvyh+URHRi2+hrrx92FGk/CVNs8Qnd6ym5EN85CysBXj/eho6dPPUnH6/D
ISQTyxS3f+6HovywiNRYFI2KiMjyBCzkB65Q/orXeTw=
`protect END_PROTECTED
