`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D367ivdBBzIQb5IL06TlvgIzpa8AnF6gyVTAonhf0lBPJs8yuFWDYAgEWhPascgx
GoW5nz6g0W3CM/axZtcF+0ovq66LBO2cAEWwmpwm1YSMZG+PNuWwr4ajlgnpd/B+
2w7ajOenrn2hW+504ZnmJU89WZ9eO+ptjj/ZgEC/qEdEAV2wuy83Z4ZQ6NZecyql
FfF58EptWFnVyjnBl32rAS7iQF/Ri7RnCWPoglo3j5+2tTGuCWZj7wZJuI0r8RjX
dclHUxShwJViiVhHFXQFkjGOEev2EcSMv0uVne84b5/Ek5cupPhymWjfKjgaNoFe
`protect END_PROTECTED
