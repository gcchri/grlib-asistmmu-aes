`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pr8GpHu+VSOG85d3fCCACab3QYRCrUO49RBPwpAoJfItzB+Uk789ZRQd63viPQIA
UXjPL+AnYGgu+0EQVtksc7rhnBVukKGh70ynoceF2FjOlbft2CrwMGjMJzMrf6Y0
ycFBpGX2ja5Xa16JSirNUbsbY5y7MsYM7+DWqZI6j+qo1K8Mx5zvFc9NH8hXnoiM
EFGb03tMgaxiy9O6ye+AUEz43gjLGVI3aD9L9Y+tn7KKy1FTFSdPx7tEoP5pAS2C
XhIWlQRJYlp90Ot8Fujs/XgmBpnD8GhXyeJcR8ULfhxDfQhpLXTQBN7V/Bq7BhjT
R4Qaa4MO8UoTZ/eHaYgLa8xZDBUKvmAMThnlhDCXzBDII3ONYq/E7yYMvGKbHKYF
+n48G2zaCdNEgqk6h45Z/6QaPISdT8M/TlTABgmudr7InbJt/bS8MGgE+oQ6fG6R
qv2f0cB3OSpoYXaABCPxcg==
`protect END_PROTECTED
