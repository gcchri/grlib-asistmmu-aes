`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AlDhpuH1YGLZ3WdwHKzb0+JyhpAy9QAB7SbnRFYpD25RcN1z1F9bJ692RYxA4i6C
Dt5R3CxwYMBY+KxYnoSzlE6CmZIiL5dY/ccKZjug0M6wquCF7EqTxyJ8tu89EvQ5
2LNVZTwVr4WPI6sTgUPFf5e3jUXgr/SaIQ+/UHOUruTGD9/rBHIjzFw3xvgA3aoS
pbNgcTXRTp8IITKU9gyr46jcYgGSaMlQtbsyRLwpXXIYYQkcBTOjBIag/qMmdDUX
dvCSRun3ZJK7ujzihbd+aAjpXTfeLDTC4BbYckcspBwQHCfJflwG+1JzhnJOHM7k
D8mPuxk+6f51ghZ/Gvoz+vy0MfymbiJYq/beLwQ1ImFYy12OVfz42psDEZHA/ppi
n9BywfpUsSiONpdApJWprRG5zOrxqG1KWF5j+VZdW31+wtbBvlvrqybYZGmvd3+Z
a+SaxswLdQGlUEgw/vHyCVcysN1EFMbxMCnQjwVRhJ7s9R7n6piN6XI1miOJoVqs
CBF6y4MVbXbsuAVjuEqUqu5or+z86GFOr09GhDOHiCHq5rfi8ej+uNVBt5ALSpBX
Y0g0/coNDImNkvArqnIjbA4sOSm37A3ebMPIzapjbFmO/i7/V1OaTWov1kh3zNJ1
KnMNPPlTdKuh3ctB/x+4N94LwPkEzLRN54bDt2g3XsrP7Y/GVNh21ZyAABee/9ep
x1v5HwFliJUEEhNS4/11zrGnaOwdypcqrb6KYve3DqY+3fiXiK6IMkiv4s06o9po
GVmQdd8MhpTfgYJdKuemQwXFORKEycok/12lkBuK3XgqiWmOxIDMP/2+OZ4RqtZu
4qk5CR6b5gdnVyY8FshrsWSf5ZfLKEQw+y0QM3UN1PgF1knuHKxuJAgfRjaPWzEC
qldXuJqLT7Yn/9WHEIGYtlM7IONsD0nTO3Fmm9FmFqS3u18iy6oRIxaJi1gjpglK
rVjjhFXefpJSVT0wN6NGVBIPDfJYObIVIpjTODNr735KuV6bIZf4dgHGE3Jimvdh
tfHyopqgP153AhuXEdfK2f9NILJu5aCjnTjLncWKfI/W5T2DFpaIuvvSd0jY9+uK
YL+Tz2JwoagcvVDgHAbXjuxh9/Sy4ZsC0MxnSGX3QMBXCn5d7UppC1llNChE6SDS
qYi7bupQ9i1HZTNewlgTawbK594+PX8KsTQBH49jMrEtbjT40stN/XAcuratvy7t
MoYfvOoSRDYT3sI16qAtTJWIRFLxndCEL1xmodDIdSRSAQx/J5omJtpzP4I2jUAS
ri/NLmNq0/N6da7lMb9bQIl659OUeANvp7wwwtyPyuqu3WQ1wlERsqTfdQeiyHCT
SKEart+ILQWd7v3+ay0kPHiGgJtkmaqtQqzLJxomhJ4XLyH4NmFjPcQFCr/gClpo
Av2K4UkU58NfWg++xfpWMWpnxxcm7UTytcSIP3FRKEkUeSkF6qh/ce4jzFrwKNkB
Tlz/mb+y0QCXiFaEEWNZ/xgpEOdeDM+bzVljPcANYUDbIW4C72GixF7qeEjiONrG
JkcAE/LX13cEpAS4UXTje1Dcox5xJmzNafLvyjJRghPSl9znu7Wm+uZyE9/xJu8+
XrK0qTN6UkFBA0/VkP40faayoeZ7KJUZBP6jiQo02jaXwkRDBWEKarioSJcyu7Qh
AV6NiX0Dhn1P2ENGWNtiUWdT8T5fg8XDUJ75vERlCW/RxSgmuPjEb6H3CtKxJx+6
Q47bcd6bRLWcRNqgQyLdtCkr9zr7i1kA5TxIyuKmd5fORJLzl48NOSjt0UKhhKlq
6nn9Z5XCo43M2xDjmCWV+JZn1IT7NtRZGv9F/0NT0cf3VfSQZAzdgoScS3ik8fEX
`protect END_PROTECTED
