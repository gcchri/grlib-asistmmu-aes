`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uy+HNrCGUX2PLXSnvkv+hPumoAD+v7SUUDCcCd3adeBA9A0syEKvcmzbLQRT/BBf
fzaYaTEaA0Gize9DssVl/cWe65u6es1z7/SCm2EMwB4BG2gDtatgLjG8Chd40DIf
AdPua2HOKc/qYK3Uup+OQaLzM0x0K4a6gxW7ymIIaZEfNAaO7n+WFdbJi3zo7j9X
H9s6iC67MhPznM49QsK3Cumr2hKh6bB1rzpXmE17L7mqXwyetCG0kgtJDY0bpO9D
ffB0VrFgTlW0rZdF1QQM5TNNyPYTlWwJ1bKUPHvXUnjdkOH0zFtSG01mLARKyocC
eYSFYyzYqten1QA28mH6/Ob9ovKQnaEsvzrPJNgZke0IJwPXwm1FEZgM2EJzW2pk
P0zLwsRrdMIgee2wndoH/A==
`protect END_PROTECTED
