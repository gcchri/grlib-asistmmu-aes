`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6WO1/Z+vYwcUrlYqbcgNKog7r8fZstzciJsmlXtQiI9UB/gJ+txRUrhPpRvBRh7k
2Aaqi+4bDL+N8Z3T5K+LrnQIiHbwYLtXoFfRRdeZJnwlvmkpONN+0xRLBM37twKG
skzkUKgJkyukC9Cn6Nnd37AUj29i+c2qzceSrCgxAQSTeVEBlyasa6ToivsxQ8o6
uloQFwrtQbYGu+bdoh+gur74n9ZbS+ytn2G1CeU5ZMAEgJ7+icSXHWcdp7nIX9uv
PfrN6SacKjT/usKo9ntVUo9uNtYXkZlOkNqmwYgdJtI=
`protect END_PROTECTED
