`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r+qYWQ0QZkUMvakohEfO4rxxhm111Dad4O2GLvOt/oX9ikMAEB580YjmvK3iJm0+
udd142BoIUswK4kzq6AMfACG9HXD8R/qmnbXTXLqd7oZD23McE5BXNN2zi8Rk0CF
hChGZy+SGAf1xzVNox54b3LOy8W1ZO9j4pQ2nHvgs0x+GdT9YOlzokZ3L7kuXbGf
A00P5BSMBhrvtB96O1cjAhGpdg3OPzDWm4TsgZLxY2cOTAs+ZXZPipTp1nZRqGr3
BMU0+8BTJOrQTPz1NXLt7I+nA1xO8gravIBAS/sYRP8=
`protect END_PROTECTED
