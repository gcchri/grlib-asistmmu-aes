`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+gPM1cl9zHvlFms/9YjA260v9M5x46p1l/mIht7FdBrH/hGFqGDY1f6/ipaAOz6C
NhkUCUM1pZaf3BzXSK3USS7/Ear/uhNsLwL61CxSCrWw43cQ2RL/VaxXCn4adyZV
Jg01ZgeuQ/9XtpfO8u7CslTO74J4LwacVt3R/EVnwJCtgJpk3ixEw5iLnauN8A3e
7/8T63LPHFw/ok7AaTLsFIbJQsmrQDYxm9XgyVwUpfk8vC+LUCdStPXkL/M3XEpy
QSDYwgb7xXR0NMi3X4bq+i0Cd/cWGl9tUDZ8CUyss0uVgHuGlG6f7GolLfwnTixY
iVVz7QQpqgUWTkc55UPxeLSgkHI1SOVTI2NAqay+eM+Jeyj8klLw8gNMYOpHuVQB
KTLT+5QZcTDrLK8vT+vWlBkVg6EsNJSk2Bo8F0vLXh6nMCerU3JfXWwZ0XZl0nun
8JtQY7elOOkNDJFVzwJBLV+1mXW8qQ1ofTUa8AeGfPmRNcGyBTf+8ADCP2iAFvUt
QFFLCQBstzWqSd1tsMHHlUAOvOCAE45jIAlLDLt3H6bliVBCQOc4c52R1w9j//ZB
o/E6s+Wo+xXt8nvhpeVZc+pAEwkDGfM3j9Qsn1m4/uDIRyIB6MYacXyr1Rf4nb4g
w94VV5WMWZFR0uEpZcr81v+yQtUSeWwaroCJUAp6w4pzxYieFKulcGkSJqpaGHJM
oJqLBDSDZV1F2c7dMKn5hZNhoTtI0vCGM1uVwc+tduFp8mXde6etnqd3tca1a20q
FB8loKpJTNgk/ZOocGOja07JvDhEFIT6V9foSeuqC+knBfYKZoqHzONnR0zNq0ro
th/gK46gkAmC99c3/gAPRI33kDULWe8akYqn+zSc/D7LPYtH4R758A1MmAMDgoYi
Ft7s+WDkmxnEC71Q+Rp0dM5v7TR0c5BnE/GZw6Q6n9iLpfF2ggdKFyoNM2PVqtcE
GCo+Spdf/7wLr2ZW7RbOTVy/gFSE2cC+/aEsAwxvxTI+AQ30PVY+Xh56poAcgwRD
y32IONQcVSfe5vqHBRco79I9kMWf347f9QXWsg+4Bxf7K2/c2lRVXyXNA+6hRzuU
yWfxaOwgBlU6RC67N9BCsKooleaA6q8GTB+yj2DnF9T815e8TBUFT10AdIy2yrp1
NohH7r8vjfcLGFUge6UA1T107oQE3amCVqvllL8CQ4/d9A6enhkWEO0rPZfT3CAO
hEN41pB/xqZiXgFYGQud/2zNX1XMju37AZKLNYLrxXfZotS3bJuboOILHD9TmCCY
Y0X1f2THWFj2mcIifeBgksSl81Ca+/n+X+DgIn5pmWs/kkS7VZGBJbCggxHPWLO+
lYCqwWnaCpB6GNKmDKyvsrqCpnIDv/k+gSh02+LRNiNbbPXzVEz61M69cAIaSDSn
BESII7OX8lWvTsHZuYOJjLtuw7CKPq3/6H1Ps2+woZJV5Bz/qHkXxqKwMDkW7tKD
klZ9IbIDSmX1CWYnuS/hEHJjBkQ70dpOp0tx3DNjORERhrMfuouWlvGYkTX+DIfg
c0TA5HQct/UU7x0pPBj41+FtmjSj89r/vGp/vW8OvGLZdE/DmJo7KZcj2OEU+sZq
LZLli8JGtmAKpLum4eYt7ogsdPlhKs6OJUtV/zVJc9bw0ypLrNbbWOPLMfnEVN/B
ry+hUIUYAliJa5xMrDCGPkfqTp+Bnat0wfWyiK0lY1Q5oWG7CD49s+RVZZQQKtsn
pq6pmyH+wl1/OBpBUBOcrqafwwxQwtB6ezTpun44soAy55MKhAZKLSH+qvZ73R27
lvenPRvKIummcPRHf09zN1u44WkSF8lPaTOBFG440aP1NpIN0ffGOxVS2SKFWQyR
FopCdjfz0SNoMSViag7NfuYhbt8wXGze+sPVMOwCvc11vIVWylXneOPtmuuXx7TC
i1GqdGBKqCvVY+oEbcRzNRNjD8p6kq9dFg4JYjjaJAlbE900LN+vb8zhlgxdmyY2
FRqfFnALHDC0OM+22NZq0vhoJKOcG8FU9DJqzDxeCHNLsypJuFmdZHIGvHaWIhen
qJsFwuur6ijUvaSooxn7ZbZWzXFCMuB7LWXkNnfYsu+uKhFBkuYJxP07NG4jS401
I03dnooFF1/e9li2IXmdPIdamRbr2Hi/ZzlAH/Coo1q1timF761t06L8bdMlopBr
Xa2ahSRHgFKH/59bo06sDeSuSFT3qzq8I6QlT9C73VK8CtpLrM+Ed2wnKn3O1/0s
ct5oizEMKhceZvMmWavguDoavCdhh5jUQ9bYQif7O3WirdSx2Nx7+qJnnH6HZMkB
zFgHh/WEhVGpRqVC8/xNDSE6v/vwK4avQ4yCJieWrU627cDq+UDJM4iz1JHkJ/Ss
Nw0+64nFYhbGfgHvKoPXik98ZskKh2MAJDQXp9lIJVgPebcEKHNdf0znc82tKUlz
AtQ5obgTPLUyqvq1tG2Ukg6NTxfyiLuxyFUC+i+G0f3r/wr3jcKCEa9H4E4SafH4
enQaO9DyAUbnKM/xZ39Ny0MDNMBDwgLZJFwOhsEkzKwGOuLk8n1fHmRWNssCY3i9
jKbjBQmWTPJGv+qcw/UQX7zkNXPoD0G+vamY6aI2HxfCrfR7BbY4krd8MVH1sDba
QrHCruK5amhTgonRTOnhGPsYxoK8xILu054Hb9PisT6IyUirHVMttDEVrOx5in6h
7UbbXwDJeFCkuzdvsJY2VmnoSlLBzOYQl5mMeV/0Q0XFPUYU++lghwzrjEk+sXbG
FDc554jjWpU7PYtQ+YO0vIPPYLpBZRjL8+YG3pVXcnWESUBwdiR7OKcGuM3vmynZ
zke4d+ChFjg9T0Miq2y+PyzN+8OJm2+DQWdm7ABO3nAFKhCZq4qUt3+XFmGEFQ1B
cfU0y7+ZYamVQZWo8mliGDLHxi3qafpDhYdJDRbi+6SMhZKFj01IcWrzNM3+4oMD
+8abLkTj55d/AlYHbTlog9j04AftPOqGNDyv0M280f7ljE08ZoN5w7tC+Yx1S2DM
U8atLWja0/rkRVdX9edoCHMGRuTUQ1u1oz1ri4I5XTcIBtQo5Jdr1lAZEiJUMFMk
8IyhFwYkyDq2+3XLU+IrApLW8rGLzY8pgZjM4fQ7XoBbZy9JKR8i74r3gn4mH7Hh
DOl0bb5a26ehik/sO0XD6ElAOwPJ17c1aQraT0QFXwiSh2rH7+5RKk3WiQxaGKo4
LQr1F0a9uQUtJIsA0m6v2Wao7y1BN9YfqbUZLJoxy2ibMhWPVU0LW7Uz8GSurs1u
RsXh9yfZfuMdUhI9AygnbmzdgjX4Uy0FioWJnKr99hXmnfq8JT/hfYLS3thahuf6
JDNApmtEzin74NE29ZXjj5fga/JTG6GUy8ahWJJsx21SgQmJqTvBERzr3geKqAO4
M9L384M0nMdzxJ/6vRnyZIZNA04rk/NaNhzM5VAa+bGmxM2FgLpy0c8qPaQjIHoS
G+iP3/vdWC/kF/9fuWoOITrND+AjV+e0pVeRlMZsKuXm8hdQhmZppOTP8LBS9lvf
ZtvgRIswMnJETqbPmdOEqGVoJIzgyr7PJG6v+QJLKW1IcuTedOL8i4o/Ak/2xy/g
aAVt6vTRPxLoJb23W/OgFvUBOSs8AuLED1paHUOgduBAHHoFC/QELLdZFRhvFYgF
OubveUjM7VhcxXPPOaR2jQCMrn+qczoBUfk1rFqRmHT3PuYqb+IrPmAdv7MkDVbz
xTgqrHbZQVRxpEZRnTkri8qDYyWg0uPqj7bPmxuHGDQqKQqzHF+5D+hKYoNEbFGu
Tf+66Nct6zPJJbhbrIPPJo0eunJpiV3idL4Ms1x32Fx7eByymG+EV6R4Kra3zu4x
GF1zJMlwn6q7A5z3UD7kC7LH23tfM6tHPKVk5RUCf1CBm4qkKs7IHzxzq1NbZOVX
863fTPGz5DnHhPly3I8nzRWvXR2uG/eWemRi6/viqdssmmQztT3vYD23WSQtdA3m
fEJZbn8ir2AWgtn8WYNU+5IAK7hbIqapFIds85OqgUkJtwLkixbc0ScOxV0mxbaC
1Z6MscdF9JiDKodgUo/ddAI6TORCcFspZ9qrx18bElX6c+YJUCml7oNQ+Oxhza0j
7KClA6qwkDrPX78CZ8z/ihgxmU7Q0EK/Ww/qrbQ3FalI6k0Xe2Dzz95Ha26M2xPm
lRRyImK7OX77rWgI945+tBLvKluHuVwJ5vwc873k1d474z3WrEa1B70sIyrWldTh
JoV8uZgqZuNjI6+IlGEI9fgqKqYl5XJl7fP8PGPgppfCINe6V+ltNj0Mn7Psl458
o6A2zPOo4E7Ei4E5ltPEgAMM/aoax6OFNVejtp/vaArl7r9sjX0ObxECRxxe7PY6
FiXqI0k2k8La1DImN/5svBjWt+hibar9i5djYXgpdiQjLZZ/pbO+VrqLt6Wgg/Bl
U8hm5TpP+qfJnODtqmizJ/267pJMOyi3qkxG0KK7pm5+T7qWpvvVVqujN68myFTo
rGj7RwhIMioNUXx7Rnh/Agt8sXpNkLY5WWCBnITQny/EMgfMod0ihop5+coYypDD
SzkdnFwQKXpeMFCLv8m2yILbM9vXQVMeGnJZo45gBkACo39ztHYX/38ax/j78PXz
XDrGuDCSIOEE4ulUgojPviqADZ2U022eXXrgL2QMuhXvcl24CTMwBt+XihzjKneE
x65AqREh4w+c7E5sAY12+o/o5Mr++Pz0M86rIEr3ToL7wcqg1yX65GD4cCn9JF50
8Ib65a6qQTmlwT5EdJarl6tCIukSMJ/GJ5r/GVsjQguAJpprVUGksJgH4NzyoZEM
lZvwkj898z2gdyfqr2mZ7Vwxplrxu5d1OJb53DG2BEyAnfXBCmOm7jMrP+45+82V
CLXJBjYd8cO1m/Rl/WE4QWAdmCE2XjrMQHBxJg6VXmrmEdgslDb4Yk25w2skGzRv
bTAGERmcZvvYJSOxIkfwLsHTrLUrUBy9rUX3eTCRCX6TPENKhXTXoeCv+qhviPiQ
3FXmd296fEUEaOAOiemIhvxSngI8sjXpIGIP2nCThjv/dyaolaQ0ezqmAw8BHy4n
UvrS3HEkyyg5/FlO/FVgWxCONN/R/t6WtjU3HqWj//PnAOryTyhBXen/ssV3SCdU
U7eybwOcRl/jaYBLvNOGwUBULPEahFQ1UIlOCl507PwinqArdB5TcL9kCPXLyNuj
O2FCDjIM+ZzwbqoXQz/uZaUJcWnU5JcCpv2C2diW1ZRTi2dkpxNMTtLQMlFItR/m
cfMaj4rZHLCNZ6FsMnjbJOvRexKWPJJR0uyqrQHE7vbL1sxiPS97I/yPdT8zPCED
Iy0JuGgTfPG4PhhUyoW+X9NYkoI3akMfpiIFtbIA+DAlFx8VUAxdizjopJq1OmuV
t505CFZOjzEjWb9sexLD1vGkJtUBRQCGURWB3BA+q54kxXs7P+jvHNOpjHFl80vE
m1K+gbY1KSy4kS4+o++qeOqaoHoZDS1zLHMOObHQGPgDJ+qmY4Jye2xb6OGlYV8g
YKCtAJPudFU/e1zmuuhaqpTgK/RXtRqaTOfW1qK8x1itTNqIaa+FRpdDmS5AdfZi
1cG1fQiIND45WP6jRbwMpm2zgKg7sx+YZq8TVKeISVBHN9Z3VqVp2q6Oo/3yGoLw
spRId6JgJFK2Mhnck7G8gIZA8YzMmZxiOP+CWtTOOVeBLnAEqgseB6lQLUJHlF8u
n5rRAbkKnH1VfEWWKuceNyohvnLsaJsOchj6zrlsn5A=
`protect END_PROTECTED
