`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8p7/6VsfM7f7m1oQwdN5aIh1/bac/goIGj7iWpUkl0y6ppSQleONZW1ky3vneV+3
FN/OQbsVzy/wbFm68GCGQj5WLtK6ujq43c/PIrRghS0idBEeNWb+0NXTUyYkuz6t
rsRPWDEAjwEkR92KnkPeTxvqFY0b4YAhjy4Xw7J5DLpJJ4TZNmx9pTrc0Qz9PtTS
8/VgoJ3K9oai/dIS1HsEu65Ji3q8gQ9Q5RvNYH3wb3T2Zu2a/AKMfgZrnoKGxBT6
mfean7GkanC8vNLeF/IaLHp1mowe4/WNfsFf4L/vyPV6603B9H27cERpvY6CKnsv
TH/Pmp+dZ43uF4VIQHVyrcyygm9k+CKvTwAZdldoOr7XkKXAeWf7cOHGbEQ0h+YM
xj1838HlDmbuhq4fC9ujtXi7oAbSkM4NIET55YUlSdzGalF0XHv5DdLKQFu3x0T8
qe10Hywev2tYHJpDIUCJ1bX+k5zfqGNIimvANKZ492uV3vMK/hmsYRJ3Z8xTeqGI
9/Kfkdr2kLx+fF3vlKKq56wuEdQOz4tTESazUyN/xGM+L2Jc+UYuswM5sK2lntwT
2TSdqcrAcbs5Tzfz6VFu70N2u3iGNYpVp6yBjRRHyCMx5LPo3fYow8HFjr3Jmr+Q
gZEgMUdAbjYsnHZC45LH3OG2opCzaGKthOi2nGuHiM0wHqZUBZJLRKXWSYcI013G
t7ISodiSXZdVj00UPIC42Uwsoq5hA9r9gCjKD+EB6U486G18WodS/4HK9/qXEEP8
aXFq5ZJ2x2DFtO45QqXof1BKvT/BTmsEvPUSvk0h1mZIacl6Z1TqLBQ9AAAALq0W
yjCPxF+geelYKcIDHHleZmAh01yH+fACd50IvP6iCBHv9rsUgQjsaIooIWSJqAzn
3mR+ZTb8Wlo0n4h7TwdqcR6um88VYh6u8RJmRZHbyTBwHd/62wF5VheOLa8Xeb47
TvmdL5F7uR//qnJIDvg+VM4U9Ga5lFt26ll4lwFcBfTUjxhwE1De//mqHRP8FDIm
F1g/QICwcqm7pL51ROLywXQKVC2VjfWNJuM15Q39V6vWnnl42TcwgFVRk0dCuFoz
hbFO3BdlynVgSua+T/wbiQqCNKo+g2cSfZJpOpctErIrFFU+CA0ovRB8PLCaNbIc
gzDFRZk/VO7lGG9MYut6I2R03uwHnAvwCX7G1bMULqXTPcXAf03dKzsySMZIPe6l
AWI25gtLX33XXrkrPl1bnSCzAPREAIfAvVB3To0d2slJKaLpPrIPSWDh3b7ZuR2P
zSuyLlRGNVjyvgO4uscWMWbCTONSVQtO9bBQ76rdMCjgLhQRzfHPWtIYQFlWu4M9
n1fRZAMoTQF6rqIXwoKnBKRTZCtLWGVUqAUCDfSsa+rJbbnO5wB/aIv3rSYuvAL9
jcdZq58ojBS7hK6b8/zl/FmSEbZkwVAUP3fV0BwZX2RsUWJKepvVjLQm+i26eymL
8vxgMzuxi6rvV2dHUl1f5JRLHw9uhN2z/hpqWtiLWrBxwWjUR4MMxlml2PP/kvQH
fSPtPwUIkwBjNjmMPiddlm9g/twIw5pU136E1CW4c/dXSUpHijsbky8DbNDWOH5r
thhxmzE4hDdoQDld7J3su35NB7w6Th8U2mtx8OqyjUlbQDdCLbI7aZLVenbg5MSN
u7g4HWkPWEsmby24dxND5/7wcKcD6cBCI11YcNFDxpqOE6wPtVCz5ad1Dc7or3J5
uzgSyetxWt3mpF8gRfbnyccCJVFH4t5KaeuFHxI1fcHG8bCZ2zNxo2RSb93emGMk
BGlTp2fN4yynfGS5/cnAqCHN0bY2EKCAkgZc6QjhLCZWRfvQoTqtVDWQj3xjtweQ
dp1wwEPgksnlPh/DRxUv3FqrmG60v9YAI08n7UUmbIs=
`protect END_PROTECTED
