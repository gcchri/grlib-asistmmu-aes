`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Uwks6SjRXCNsB/nCYyoOehcQDyR9Vdwy1IMLTzj8nj4md5AZdoqZR0fCFUhWpn0
MCMgQUG00no8tVJa6zyro4H/7385dWxRwYGKWh9OOpMJXGpuri4IUB/nW9e4xQRH
4ZOi4SAun0QFinyxuyy3kHElG8KYbjLJILJUb7opUdf5y1RVx0Viwv4ZcQMa4kgs
q5TLlNzXxEYQu2F0gYLwDc465qpS6cLYLSPMWJ5cjkI=
`protect END_PROTECTED
