`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0KQt+5K+eX7xmqVzguu80bH+bs/idjANkwL2V5otwPDTJ45SvN3/G4NfYx1ZDiU/
XPpeA0hj21nH5G1obDnHWkkDJSjm703bD33g6eiQTQMKmVRnaI0n6sDqRS51h1J3
NFQXHgspyzM51sQbZ7caVi37COmfzCe9ICdmMjsabb4Uc5xasrkFy3ZSMU5PwGrb
A/NmQQWxoBzq7tubflYyBjtcQZ78QlWWHD6MdHVtfkKDwEZkoWTcUoSvN0QXrXnb
vSBiV1U5MM77LdQlnAnv20vDH8rtIGaDULwmkmoyvjiNL5W9a5VKlBXRIqtP9nHk
GFnznog3HTKwd19Trk0J3TrXmrXvTkqjUCNHGK+qFEHECCCNBLffPtt4FTIlnyJF
bQpEI29eZ9EAuaJ1JJZSe9CWHERCJKVapvi4BSOl1BgoPKq43nJs09HTl6wbSKUU
BNUCljR/klh8s3teR0LNxJAzbC/PtpJGlRWbuBT3BeHUWhEfpL2eqPMDOsD1AJz8
mbUwO9aKZo1CVsSM4PcXi8QxOxa0YslaWHiEBq8bB4Evs6iYST7n+ZhiTFzCGDLL
PGwrovkHJiVcVlmtYCxNj3UNmO9Uw6t/0SVwL1gs2BrOZWTANlgtGaaWftDSk6OB
jJRxJuMAp1wPGP8Q02uHbumb2O4bNP//B8wMurpuy/89zzsG6MiMayrWdFJcbWvd
c32lPnbsobAUbUzORP2SWa5hBJYJ1HKmOhoKVgIiApXhNkZJZ3SNAr7ZEbHy+qnH
oxIYSdwqLwuNbnqYIODe1/koKBABayCcVQ7kIfBFqofqVaA1kNc9mGNInx+U5UMY
yqzj4mpEhindj8WWJ0kAi4q63jt6BfMy66nL+rjAA8QqZZkqD30f40exxHRb9Tvw
l8bj2e5Eb7slzN7Qo2ZdSdT4nRaVyVEn/OHrUT6rSps6Va1YRrZhdDzifGqwjg4D
FXFfmeSxOUY4ngcajFRqFs2grgxsFECudx5JtKZOwlNMxZHIqQcjzTtQ9xP1aqjK
qVmM/YprKTm7UTqBKrilg/R0qFXHey332Qg8+uS0cSCHZViOKKkhKULPkWGOUj/G
y4JE2W/9AqgTCaDybwJjP0ReQnpLbZ62ZtxGyDnb61n3ZFx9Iwno/scDeABxXdWr
/ZVmWuK/icviMB+09f+kQw43Mxe0NlABhaf50rbG0COjOkK4BkEHSbiTxbOYaL3i
lKSPC3KWHbhNv0PTUHqmFxkJ9ItTeX1B+gjUM/E/QdX1Qy+kEvckTXmiK+iVvu6i
QNgweqs8W/VMkH2srirJedWLFLpaBRLlqwEFgtsj/aZ5DLwwrid8co2PuhrbTAyx
HPcTqBC/k4BcAwtL2PAvH2+Dcd+GiLlCm+ZGjCdnVdC7yu0d3ti1svY5VVASO1wW
pb9cc7YB/NF8cTBRvO0oTos4mDg1EnXmxMYCccX+nBrdGvIXtp3eFFXhZo/lhXzP
N7bFrFFOviQQbwW1yZVFEg+fLUmI35K5eK4U4IHgv2aTS8Ktjxdsm8B6XL7EoW1J
FFAOkb0boDmkSeApr4Dgle1LGopvac48NyA8W/5FVLSHiL5IjNGBGhxGdBB3z8Qv
23c+2XKd4dxeOT8WPMN7p+eM3+wZHGBgVkAITTbDBacWcS+jwiNW1ygyTp6d9TCd
9uMHdGU4Xr8oGELqOhjvrgIOruDg11LQJXgioYROpNdOE7eT0IhVuyZO3xt+eqTA
FmF5GudNOzRelJ80AX8lmF5yO3E8Mowgvy+GsSmfvaGsWzD9mk5AUrtsZqXUgvQX
djAkAurX2lmpNPbrOhaySeiCdXg2MSmyLjHrK+rBgA6QMCvTU0LgIDnIoHVFQoJP
JfenWuTntW7n7XMghc65cMscrh5XMuwCEu4xWOMdmtAY7OLD1Kz7TjNXG8ywlblh
jwtenKsV/DuH8INCPa0TjL4Iie0Jo0XDGvWz5JL9PLnXTibZpCw+SFnYmJSEWsKR
JhQmDO+yeLcEewoPNsOdV79cIcspeEN0Bngw6/M7HRg=
`protect END_PROTECTED
