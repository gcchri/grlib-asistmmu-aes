`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dg0KUopTQeA7xGd7DP93IuZXD8+qNchGpAvjWqMwMCgse5NNf/hDowf1L+dOUKqy
QgKGNuuwGaFsYzX9GMtlfx7qMgcVle7QvL5XU8h24jVgPm+cWIPWWkSu9jdlfVXv
CXsUtAzM3pr+2ASnLs9wV2Wp79FZOSm7AwEgzpDV/XCqyhmi2v9kGWWgvjaR19i2
lOPOATPZQu70yEowrmfNVpE0Aic+FLWhx2XBRWyB0q4moVRRsBqPESV7I/e+TG37
IwXbeUp819GlL44gIuz8XBUZzO3FtXXDCl6k6u1HaVzt9H+fq9eExA2EQEiOGKS2
wGHbazj3EWDLyU6XF4f6kPmaEgLGE2pTetCLBkW4InIB1Y7WOorpa9K9jKFnxXvC
6pz9lWSr+GSKAjZJ1RQPxu7RSOrPtnKfT6LI5QuLrHyNm5Xu36n9IytoR+GuxfTr
`protect END_PROTECTED
