`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zu+R/3QcAEDjan0vSSRu6VuGqdbnOGqcjiwuCYdXc9czegBdJidsRorUDi05eCSU
7EhZYzVvCXHGT4mxpCQfnvuc/EKDcVAGUvr4NOUHOBftEqKLDIjO3L3pn1/r/+AZ
UCPrm1dhu3X1mfKdVg2xEtkbkV8wuzIrQ3tMLQaw2qut5KHRlirqVDcH4d1yh6I/
dRgQibWb0n15melI585omDSADIXdfa1GYe5EgzkoNzQY7nxh0g6ZAD1EwKXodt3o
VidfOGHJHgnH+JW+EFYduYpM+UNWB0vfMU2pDdpmVM5aoWIW7ZKOqjKUDY4rC9sx
RdbvVvalsGpSdLc9L0ys3g==
`protect END_PROTECTED
