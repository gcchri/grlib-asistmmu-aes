`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tYW/bJXMEE2gM22iyhmDhgZ7SkYRYb68p8K+JL/JgQ0KtBGgXiKHKSXP50xJ1y+E
L8cV4D5lYIENAe8cZis4WHHoyjcFK3o8ebN+kZq4AtPPmIDvs0rwO6Xbd9ZPufUn
lxNQwt97PyGaNua2JLmoYhFXp532XqYYZjsPRhYaWVT5FparubqOMva4+UfscUTn
GgqH2VC013qFjrzAHppzKFI6olp0te9o2TgkZfhzlK8ke5b7fFbNpd2MP2RkAS+v
thWfPrEJCfIRpgl+HUKl/wrfOir7h2Nti8W/qPXs+hyGWIBi0W4ts63upDpP7c4z
txLn9PWvBdho4VgwvjfYtWzOga5rzhy6gLxITNV5oadYHEiT8rpRigh+SKRsq+My
g9Mx9k0AAOsebyzsJCx37knI40HcvcTc5YQ6O3kAsAGAUfu7l2Fz6qU/Yc5Ut0D8
n523Mm+5tU7qzk/Rs2Fn461Laq4gaNHUi/845pc6EzZPJ5C/O6X5cbQ7ZUmMiKbl
7mquZL1BjveaLrKdKUTQOdSEHu2oyQ3M13SLdbqqPe3+SF+754lxUznIYBrpxzQC
ZWI3SLyQ53QqS9BQFUXIl/xyDUK36sHsatliLlPpUr0=
`protect END_PROTECTED
