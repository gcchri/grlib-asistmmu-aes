`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OllAGEXwZ+OqRAmhyAj7FPT8kB/p+70nRAO2mr8U3gYv4amPh7xecxs8Hw9mHjym
Fv+Own9zu9d7H701K0dy0vux+hzni1cm3cJJ+wmnipEI4RaNBcLn6mfXzRLASXZs
gWNdIzQFzq0IScS4y+XHnlFUuSj5EkPFA9aLBPJMZCe134uc4If6kAbXSjeWL1lx
RqeksHPA0gw6I3D+eNBkOumgB1QXliZ5tsK6pxrEIKRGp7Fn2r/vruON+AFAQkLs
JjImqEVypnlZ+ceRuTc4x3PBk07jOLHPPaks7pVcQTpQ5Jdyen5vwVMxA3Bk0M/B
ET9uNwRPsW9StR9fBJHf71QiBZPJwFw4tgOEuXw1nClqN95j2k5/nj8xQXXoYBih
5CV1NWDaWjeTXxZZ8XEUEduvjcTDWEdnScOczzZiMDwmCykeqUomI6iyLItxccyK
gi92YZJQiloNaAobwB1g+0o4mBonPqdoZEKkjhcBDsmjip5mkojE2AIP7be8qtm3
fm2+LcXSKkXZd7wQvZ/zU7EmXuccoL2xVKE4rx6tpZSoS8kF399eyhtEMYA/MEzY
TlYoLmyg4xR+KmmU9EDw3vOaLRxNuudXtHBD173gK6MoDU4017uLcXtNmtH0noSJ
opoaEGMFLQYZh2oLQ3gWnqQmedqXCuP1GfofTNrUYNBOdVzogJSopRjzLKejOXRb
wLN4ReZhDgvJ3n8TfdayH7+Im7Df61OcEafgf2EPBxG/uIpimjDIbzUwrAP6McG1
KrqA9U4YrcWRPKAxp6ddTNUwjxg3UCavUQi8awDtBbHOLD29EeDzdXnlQe37M6RU
FvqWosvs3K5UjIveJfkZqI0IgFzPlcwy7rvK0cQV6Yb009SubhGPklNiPWgQWnbZ
`protect END_PROTECTED
