`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IHhHuGLslL6KpwKK056ASGXbILqfSDmy5KLlChSu5sfMIMlZ6P2gCCN7lvxzohof
zUwMlSadQS6pez+sPzyIUiLyGPlMMNRuQrV+MiMdbj59165CZu8RZc6LCK6YVx77
/p7c+zHXPDD+FTxkn8gNE21DIbvQVME2jzhhaRZc+7IWe0ammEwvRxeOLZTLIgpD
MZUyeHhfPtf9lKA45xMtjGRI660ze69Jl6Spjs9Zx/0Zlqzqb0iuclqem7akeCsW
Q5it1jnPb+UXG1kwMHzmNQ==
`protect END_PROTECTED
