`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UVCKX0d35oKBfHzRPafHc5tDDbXj0+hS3gB1mb7G8lSR+/HAiiG4PRHJ5qFpI0wl
Spube6zY9sQy/6iUZtQHLTn1awLKZoFvZt2noBvC95qksxL2Qy5762Z+Jy6rsD9Y
1dB2zcLHS9bem4MyCuPzKMpuxuAx7Es25D2aPEWigviMzpW6P05EThejdGM+tpw3
rErUjHnPiZQZMA77G27zrXzQdN1bFIh/T+HtmOYm1P4mui4UR9NWXZX/wrG2k+DE
gaFzksjT9vQtLEGHJzUfpAqI3M7V06RhTBrUfZ3R1kMZPwTjGhtSNluNU3ATydq2
K0uGk9+tDjh/fbp86kDz928wjWh/2mBoglMVuuhItuZicyEQw0BKUouJziQeCAOQ
pt59FSSRECwrroj6NOz7JpZvfO9Qm9eExMy6rRADoJyy+vIQCoDzkaqWq/G/Otkr
LVl9xdVaDsrOi+Qm8V7BJE1azexUVfpqd02WUhFt3NpPwiFOvzwji6TIesdv2qF9
BXUDIMrTC8t9tFvc/M+gJsdl8WMsMuWzjfuUQxVRURcNnygv+LxdFI2HFV6dpO58
bZNg1pvAG4grhc2Dk3pN3n64zxCjxqed1D5qxmakEFJSV8EBr47VfaiAOaJhsd4h
qDcIkgqGoheyYhrzOzfisbePvpOjrMql63tV58McAYqQ4zuwSHK2l5m30r4rux2/
lxP1Q1nk1/XcLjEn3/ZRK00aZ4fdYQ3TDUH9YWOWihlr38BMUbQuF0M3MHVWayAa
cNGKXy4QI6/slnUoh/Zjna+sRcv6ANMTO7MBtAZoznxwhj/798kEr4qurR6qN6Xt
8sPeTJGHJVx3D62ba5CQFrqUXCvUzEK1hTZjSaErPlLQ672hwxfkzgj5NfGVWqxf
EnHJdHCXPTnGYppBTBeInKsgcexS5axvEdpFAHYd6x9NG8YUbABiSMN8CgS63MoX
VlloDf14teQEQ1bMrzv3sVYmFHjIt6ch91LdaSqylVw4TRsFVNoG2dhubvlhIhY1
FeYN1d/Er1E+zvKzQ5H9iuPtzpQcCEd1U5cM0F5GT3E6qVxPxs/e23laGvRBAGuy
EO/jo99LPo8MXv5azHznlnkJwM5dsrWfSvS++iuKKV8AOEFnaU+jacEpNTfZcsy3
PNmtOPTo6Tcn1cwMi/eiPV7ZvCh+d1f0k7jd7wqZZbT6XswAwj6gARxxIBsTcMFc
im2r/E5/ywAMBCG/iCuSgfl3lzi7vtFQ4sq9g2Y1C+Zr9xPFT778LyOHRx9lDeAy
QFPkxBfMChX3Zhdu2MmSBF+IWwWxkrepFgDHzdV2y1uskUCXaBA3mSyHjnrkWExj
PsKEKcdypILl1ZeZ5+OInH4fTSmpek8SV7zCTzTCbHGORFyUllKcv3hKIvRkXYp2
XzS2GB6Djto7o5cZjIx3A54kQZWLs27dwGAtMChKeev3xE5QjGf3zQtU/+97eAZV
QxEyTHVqrQzem9MWwhG2UwQnNAfmRmK7wNGHt/ryrhl66zDlzeTZ4Q5+I3H0Fifg
19CL4KKvs99OechEsvN8YAXVwS/8YhTXxCcm9W9CU50+L8hZ+14kGXNMSzBL5vmZ
`protect END_PROTECTED
