`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6XV05+9i9MHIZkIJBIztxSe6efqCiz2LJhekKigmNxLpvRuDSSkXFoXgZgtcQdSs
qILgDO/5S9kOVlSajgfgB1Nr8aFSKZhr83KqEJL2j1e0+CYG6aRIzVJ+w8tThefR
xuJ5Q6yUrYq/sKBu54wFfAbAOzVD8zaDweRZzCB/pAtDJgTTl8PNbKLBK+wwnERZ
7FRzbozDAjHBTtHnYrnFUHnKdzx0Pf7DiS5DwK4brM1gfGegZj2XxFgn1NEiQarv
QHd8waPuHlfqq1KXRozdEtsskU53zD6UVE41UsVjnEs=
`protect END_PROTECTED
