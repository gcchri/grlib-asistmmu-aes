`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VkBePcV0fhuTpJOaTarE4fuDmvS+uii3UeDQlJzl2/+RvU8xi13lPY4IimExgYEl
3HKdIqeLpxI11aq7y4JvRu9opGfsqM/YJtOlkn82TUzDdLtRwovvDCjrma7Af25F
c4vkHog7GIBHUWnVQQX88NogO236PDjq4TcuSW8JAcWYlVLNaAtQJy1evlb8SVnw
/bID8/urkm+LT9aUqT8NNxyVnheSFeN4OuRIls24n4O1osXnC4LM+TtQc8qi4c07
BeJf8AfNE1kUjoqSTXuf7oGnW3paYBn8twGWXM7zU/E=
`protect END_PROTECTED
