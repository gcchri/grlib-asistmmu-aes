`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dJXkZTIxhWHxA7DkJNKT7NXIngMo3r1dyRCltvKoEBqtgr1JZn8xzPocgfrW+tqA
EK3F+0XX7P5CU23fm8B83jmpO6z2uv8bXl8I+JsdkgpsP6hqp5E/rsvO4oh6yTAj
Jw6viE1aLQLi11k06HfFt3RIVOTLaNhdg2CH0n/l+ZaT0Von6IQzFZS4R3/DmsM9
uPMs0yC7yEwuK37ta3YoaDIAW/b/jxn6vhtCubbVLLuub9z/rctTUpqN399MOcTR
o6zPo0wjRVfjqL8GnHV62wEQYnMz4HVTFcfWro9XY6uPvmyFu45LqwMhKo/S+U0d
R7PqZJCxRjHpRaxIeS8Jj3t04f+/jNAoAhMVpgaeSJEdNwB6rL3qucEyzIfSn27W
ruF0MLqFAn+8rHfnzsyal6824JWybHb6ixeQUboEpMo=
`protect END_PROTECTED
