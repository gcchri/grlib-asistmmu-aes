`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EX7eVn470ScPBubjhc/EDTG5+cXFRipi89cOsqBE/MVQiQCEq/aUpv+aO1Di0WpY
VwX3qk+WqUkdmjMeJGSmCRTvbsQGwh3SBDY2CHw2Fj8ssf5Q7Qiibu7vPL1edrar
H9xWdw/NrA0Yca8WRGA4RHhmL/djGnq6JMQauduDMeaIbW6GZwLitnqPxcQbf8BH
s2gpWdJwuFc45fjeAzaQ1lGnK/ibfw/J7znBUfYXTpPM9iTSwWb2TCPJlr1TB09i
oaBVsAeahycMUzdkXuH2GDWWJu0SBWhWt0SBrD5Yw/KyfA1lQebMsAJH5UOtGVUI
XLjWvVav0FfrQnG7dI86AZoKp1Grnb9cxQUgRyD6bJbom0qgeE03ZdP0UI7uYVQG
THhnk0SemacEzpQMhJ+P8GwiHhdsY4R2IgkWHH5xrOw=
`protect END_PROTECTED
