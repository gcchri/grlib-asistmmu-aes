`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lgUigBeXvHZd0v+sIm+rZCPUpe1B9gigJdw+jeQA9+gLSJ/LSIo4/QnTMYQCreCV
JKDWf1SmErJ6Y7Hb1dB/3qb4lEIh8RtxoW/m/Ap/NRDWkHciUxEV1+GQ9wSJx6io
M813P5slFHplsp1YVEvXElR2Ws+q2IG9LhdXIbR4nwkedmZEjDFtEQn2jN+xbdad
XLwksgKB2W45V0hHDcFPGwCI1FxsuwDC0RRoup2GmhHxAlP1/O4rYju0a9QKUk8n
11E9Wt+6rP86hi8DmrDUJBbjH62vNq7fyt1crQ34eAKSXRHK7AQ0UDbwq/oER7Ar
rZMrIT7SBW0Z7tZb6gXvcfMp7SkVypoVYnpsmBnCpwvWQRRi/0gGZQ3gUaWBe2iF
6Q0oTO3C9KcvKSaI0CwnzEzit87BKJqDQiML9rJpKCYa6DK9rHORaOoys8o3a6/K
JXRZToSLv7Jbge59GYVxlZFOWgxD6/t5A936OP5mo6GNaoGjChSmtOO6beWHibV5
yXO90aVE5ov1zCXS/PfSZnc9q8JTyM8SR4E2Ugc9/n1vChsmla722LYUWi2jzfZO
K363YD00Xh3csE5/o848IEjhsRnTgVy0ob/0KV/KR14=
`protect END_PROTECTED
