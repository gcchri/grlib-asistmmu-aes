`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cf2NbxsBPrDRqhAc1pQ/7K/wWilICQ6YrNll4zQnBLJqt41CXml06F5rP+LNPEYZ
mDLNkJSrLS+JWGgrcGBKaWvOF9kjCtpB1I2PDJO80VSDSuCsqV0UgynAX4laY+lD
gZJLYAHypqveQ6XqEPAkfLQfC5xw6MpzYZnXyuAF9xiJlwee+dDKH2Ev5OHfYrz5
k5xBn1fMMKUbty61nuJHSTXbKZLTAzEI9oGDaH5duB0iXBNutJM7rerzFEAVPduf
Vn59rfxnPoas+XxgTvUHy3Ci99UkeItA9hIFituTkLWHj0pgjOmuhD210wTIzwOS
b/9nGvG2ESt01KM+85uwTA==
`protect END_PROTECTED
