`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+eWj2rLcdq4HpFo45NgfybavkgcAlrX1qlYEn5/sQ/s08xRMvLgx/dv0c8VfQVxp
q2lQaPVg6iIX3g32a6541chh9AEh7V+CJYRwIZwqMgeJZ95JJfQ6cC/LizhfVdxV
UPJnI7XjRlF5Y/YrQNmCbfrMdFfUquRtCdOTHXAkKKfcSB17KLQTm8Mwon4x7/w3
A9SPEPX+PgJsuwWx/618DH2YEd5838HcxHiDeLN7yqi32bfStzYKSTNdKuR907cG
NNgp++2NOUM9oIP7751jbQMAKzKT6WQOMzmoEHD0SGVay6JgKuiPDQgNkOgf+pvp
JnpZjBJWs5GuKLiJm0AyHXAw6wBW/WgZ859PLgyUJNlv3w6UNdumT5WU042y9zqx
aD9nxt13/LDYTuKHG7kNTZdsAMnwRAVB2Vb4sJwIUpKNWvwdzO6U2B/VZNgd30Yt
5tukUtl71oldPZ5mpcuJ2kguWSwrn5aVaVQPUhLXgjE=
`protect END_PROTECTED
