`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IvURmXO+hTSfR2qFQgofwUnsJoO46Yp0ADSJLiuCWPGA8OdBzw7O7/3EXcVxDTxt
xh67Ig5M9c7xlnqvzgeLFAHHQ1nS5bOHxn9hJHh8PKLYxqp88K9TjSxP0XF+nZqv
/TtfZFrWXpwgoG3SOMHptH5TVsrvyLIhNYl967D04VYki9jrS4KwSyxdUvs3kbWF
oZIYiJ9RjTepAyd1jtT6rKpPAVeVp93aLhuzN1Tk1Iqm4EmUU2UwWiMQM5Srrcbx
RQsn4a+yXd0P3NCTL8cvMAkWYc/nKWlsfVE8o+VTQJEbZqdSvyPbjlJ0ic2j4QVX
5abroNg0mm0FzCzeHDXRxFoC3QFrUq0GiYoOtyCiVWIP7wj/0GkFRPgrL7xLhJ/q
2VbZJaJL5WZcwI0e/wnt7ykJOLxpKoWF8TMZtkUbeMagv0iN/wpfxZnH6LOe5ikN
NIodLHudoMdudUJ3Kk2vZQ==
`protect END_PROTECTED
