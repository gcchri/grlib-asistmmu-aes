`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j3lbaWGrJtsyUMv7id3SfAg2vhtAa4YyycQk5rkAx++eaFXEh+oqJAdN4e3eV87C
rCK41eXP/1QQO3hcAwEYVVVqbWDAJYtV2mqHC80tjfRqb2mmmTq9K/bo7TUzqduz
Sja3/WGA0TxKDt4rTCskaNnPXpvRj+EPQ+QfBSQw3mWkO1SpfJ2Oi/1leMTA0G9l
RgoMo5/+HfW0tcaUaSzGvwkw1anGYGLtEXIPxIGLrDZtb9LRweHODp/rY+9sdcQc
jW+hHgGFDHZYadnNy0hiThUCFRCP665moFLso58AXTtD9WuHQ6W8vtu4zMVocXlI
euFzaHDoydKAuP85wGnZRj6IOb/YvQ3pg+/5OFN5rnhSsmX29gwD4ELZiYb3rPEp
bpxw3aZWcFWId6jd9sge6ARBadsRLTpEF37w+zZqinI=
`protect END_PROTECTED
