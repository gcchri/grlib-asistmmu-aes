`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OIH8C2SIXaduYOSZCOde2G/qeQ1Am6RFTu2fnMKn4UNWdLiNdOqO6YMFuZwQl9xS
Q6zevXjGkTQXnwYA0atNJQLmIGmn0c8J03+SEvWwhTbjX7Bc9DiXxxeQSaNByjgj
tdkeshPKdHS67sZVmrEuWr5Cx33X0htNyicjgCA1Jhrvnr1/j4IqJbfwcHO6SFIW
Pqqj1A9OVX0CljMRFZmNjbtCALNTami+xutuzTulFvNzDfuYewmLJbtBpnGZxBXx
VrPeRG8OUOn/FbzEjyFLccAQ30Sns6uzDu0bAvH5RxcWJZHDuKMd04ZK0YiAYBbG
m0HY95D/UF/I6Um+7gMzudvSGUaO/cU6mfiMNvdGQrtx8DQ5D2sq8DN224Bni9Ub
RHOjwfX36VP2ff/RBDkmyTwT1X9qUmezVXuWonQuVUA5io+1A/GP2L62mx3Emsna
DsgcXEkjStw5Jeh/JcMcqiGAdzlVot4/F8z9o6CN2cV8suUgrtuggrSVSn9STPMA
8tINctgC+8RD8+74tkOykxsR4amzoV5V9l2k0hAIFSKhvKH/CrgDO9DnNrgmKU9U
CyVsI719Uhqi8gGyNV+o11YCQe1FndNWdaalQ+y8NxiHJaluRZJ+4Wqz2D6Le9FP
QG2pC09SbIhClr0jfuuNCA01NAIKeFG8T1Xa3uEOP1cIeP85Pe42Y243maG+taiK
Kb4kL5g84S/hM/kpBM2E2HYt3aAyCSqDeji6UC0l6z5ZRLCzR4bo12U3ihYmiE5X
JnqWC9SkTwQv64Sp9HIIkKcramdh8bliZQ2ERcxPODyHSkIosOfcHEETXJDXSzFS
S/VXRvNY8+YjmAVuTr062iJO/PBlBs01c/A0lOniRg4+VBPfjEYCwHzEM0gvQcdY
3wrcxA5tFPPaFY6ZyEARUYmJAUtO+Rb7nrk7hT6eD9mAcVpfsno5pQj6JJ4o6SKp
+yX9Y5kpgbIT2oQsnt4fvOtlnTcHLdoMIxKgV4ZqtBymtY9+sGj3Mw7PiPNxqw6/
ChEK3XVIIXA5y1UizQY/+mLAWuUkbtLoEGk9A6nq6//PyBV6lRWm8Z+k0wRK7INT
ehvHu31XFRb+cmdu03g1d773XYTXzfQrkT20r04cGOGU7fwoZpu3vSVsif7McUbm
soMrV7nBDNsI9iG+4mCLArIrivFR23B3L3HR0UPrGV3H5wrucuwJYAW09bVKvbqQ
UfjQ5Ps9gwmXGaqETuQ89Z/WEp9UdzQvNXj+/Z1OM/l5voEWjiNqNNwnJPaqf5z/
9qcJFFZpfUacxDc7sgkAbBQMTxDe5zEf0jZFsmrCwHU/9Y+7NTtxgOwYguTovUGI
MylW/V5nSIYnMzG/obgXwYWn/McwF5+SYru+cPjZBTwlUnbgL6OV0b+8LaWyg/UX
q6gABG/G4hYO2XuvLhIeUEkUWAKV11oi5hh5OX3Rr9M5Fj5eeve0v5BzJixkXe8R
lABdWvKR5PiXvyW0M7DIhlchNmaJM6Vaz3TEsral9OZfsMds8iQwaMMq7wCNRsbo
oVnYhVuca7CBZKSRgioo101SZplpiGAdynieSIwyTFWM4jz7DYOL3CUox66DLYAk
ftf9vUklkh1Yz3TfZUR6/eTftACvBHHWutBOwLgQrKXh24ssByeudYhUxDKrwmru
cotzcOD29QEhcvhJKRlnpC+UoPQqtPgyEmjwPnIbcbOflA89hC5aXevVClBDpF+j
1F8Y23VQ4dbvTzTUG3VCOw==
`protect END_PROTECTED
