`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aYaW8q4FR5SFU09hL3fMAq87diBLsppkPJzrek0Nuu9HRMmV3WdWucWVxyXGpBe0
ko4P+x/EC2udUFNAOEDL8z81A1QPA/JJnL0N7gn5rFGslofv7uaYwIZ3D3z+6wVU
66TZzIMxvwpR/qqgoxmDJcfISOJRNzgKTixxCQapUU2lYjSij1q5qB0zjBCEWmNl
Uu84MT6QtKIMhJNOn0A5OX/EvdovJr9s3H0m6QPyQoKPLAjPAm9eXNygRervrvVU
Gb6YcFUnMIu8KsQXXO2KEc359wOQE6Hy/tE8LvIkT/43K/xmFUSHfA57kl+CvNiQ
RxbazlWQV33t7P3hr9SdsI6HyfaCbSZPHHa8AjODZyBNgVu9S3hpx5P/Hv7RZmF8
6RcSFDPFf1z9HmXFcn+fs04GVwLbBjEDveSdIg2gtN2uBMoXC/1i17eVwsxMo8+s
qxWWsd6e+a/E9+o5XO2hYpYxarZ3IibT/uwZvdIpSZ8wCm1vdsQbiNJZHCFp6UfH
dBRspDVrHsrbUc/i+nUNxo6g2GqekIZ5plCj2HMtaO9TArM2ivWaUSZIzeDCCJ5M
jN8Qg5L5oQIeog8tBBw+bF8Mj8g+f/DqefT/I/0YqxU6GMxWjLfniDeSHCDTrPIj
DGnv3DZv1q1vqszLQRESjKPITDtV3n4AP6YyAUDBFs0=
`protect END_PROTECTED
