`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qSdDY4s0Hjo0IzTz8bWM433Vs2Jb57Y/iBLSjFLnRxGB4EYNkTmsF08/jdlIT+ya
BwJgpjCK4m8wAOT0/wmzm8DlAg1BzpzNvHLBeEqmyMlL9gE8HRQHkS+EMnLfR8T5
+HkqV3psQcHaYni4Vcviuy4/QByDvM3H89lc65OG1bjrOqHzjYtfNCyZ5N8ijrpZ
JHUs5+S0oqe33RBHflxVWJ9/TSwSt/4PXVKbVdARsfgRRd+5HNViK2e93SDGVpT1
55SBt21cmOfYT176yltF7fn5PGQAaz3xfsI1jCfSmEUJtRkiHxizu55KyLav96dO
f7FV0frNumwpZK37/oWBJ6lWtUd5TgKtR9+x/421ozI5CT179rB4+osBt4CfQcsj
eoN6RdI/n33WM1iT1VWpMg==
`protect END_PROTECTED
