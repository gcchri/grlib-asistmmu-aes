`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SavqMJdz9sGXMXWEWbbM6HjEI95nRhdHo4KABgXk+tDcLvWZn5zdRW/BYQ9K5RCj
f/CvLz5a9kdnuj+QACuxoi2ymVBCUysUSbQPIVLQrJMdbuLrOYKpLmcZNrmN6X1S
EhHrB36jaIxEq5koxh5gw+CAvGq+RjyPOSu6+3Q5/OkR86szpNwDnRKvQcAQ0qNZ
4Pl9YNT9pF8DgP4YAv//AZKSRIK3FuTA+kYpxHdqk651EPBBKKWCVXEgo3vNeW14
kiGjN8iSHQDcwTnpVpzt0lx1ZQHDcFzPUIwZShlo3cO1Z0WuPfBC3m3nIqCwQ5/q
ubx9GEXy2KDOoHsS8fUMdrD6TD5LK4DfawbL7ueulpZfUmPBjxznj/4J1q0E/xTw
+A6qfpvPvl4IlxYG1L+GHwt7ggfcNIadmLyzdrlbFHoE9WhHNtgwdSZ2l0bN8WdR
Idx0vQ0scjz1PKsu7U75MBff/RdEjk7Pb4LDujedazj1b28kzX163vibf6YDWAXe
HHwmaEzGFwpLAP9iBV1WRtLhiIB/5w7zE5MwwhCPB+q6VTCKcOJhjExdrmvj6QS7
`protect END_PROTECTED
