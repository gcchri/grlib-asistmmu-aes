`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h3Ov4Oafc7pMNrF6MHVaguf3a2YuPC7o9jBONXVVlIPMcP3+rcmeSgIngpCbqK3o
IJJiMezqr5y21H9fwkwK0omZ79ZQCbzER0aA+rtf4PBil4+8sSmtXXo3FopiOELX
03Xf/6OFUCYm1zRZ0c5ZVL4s5UK5AcyE3AwlU0kdNJlQf+vEgzGwivFZg70iaB3b
tzezkqqj+/FwWr6EOl5znw8j+7MNC2GOBqVAiBv2it5jnttKhqfO0HEGglHcBTvQ
VBxCB9+OV8333Nl24hnfkUBtRInodRj3AUJwiaBH3XJzRyt0O4ZRai29nalUhHcv
01HmeLAQjkveCZsMo2is2pTgPNVr9KIlTjq642zQqxIvueKOH3MYEPAfmOUKOEYE
jKbSezGzDTkvd5p6CwBo1w==
`protect END_PROTECTED
