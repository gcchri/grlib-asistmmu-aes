`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Gw4HZNDp262jDvDgn8Yp+6mDVvOMaw3DNYhYeD+7oGEJf1LZS12UP+VAAUwaOJP
o0A29Ivga+681ryRhxd0hgV/7Xbv+tLpzlkdqLOnjVY8zTcb0U6j6f0ofjaTFtYd
z+1aJD2d3M0YNxwBMwOpRz8+EwCp35vDraFx7X6zXC3nCzKURiH/qAizucKAFdyA
zX0hl8OgHjxCcrhMTeIHLDYPUtomBkv5KmHK40hH/GUBpr8RFovqstNtuztLpNEX
UONPmFnvvtcRpmzXwGOx1QnY/66QBm2BzvUsisJrqlYBZOgWTb9kd5rWwIymP2Ax
KA/JUyS+M7HTIOd77C+6B5q4wlGH46/wtDKFhFu0yntIrmi2ZeLQlhwZqETl6AGE
3QeyP53KjODymBER++GdLuWOY17RsyTfLZscUqOXU7rRj/GHtm1ClowKJhd81JEc
8TGx2TItxZ8eQzUKUGBRrMSzdD2oBXmODmyYXZqvWBu8RCtHgWKuFTqsbAUMO6rF
cliWnWIpFTOpgVmbOPHLjxEzDauZ+b87+VAV0EdKMWnZIMGkMz9CARk4ipdw6UGN
`protect END_PROTECTED
