`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dhKJkG/jmMXdILGNVaD/IaM/YiiNs23bjYTjZggDF6aVCaZN4fTMdHNJmvmVvn/A
LYf+c8z4ejsOFvtplPoqVUpykE6hhSVi3H1L3efVavF0SqqMasrJ9DOVIO8F6YG1
5mlWjq79xibzS4I7Ry1CeCHgXFSQK+ClVU2qoePd0RlJWNmcjsgv+mRrnSpuWklr
4nQMwO8J73w8YXxlk/sLT0tfzsAB/Bjamhsv+xOeg8uUVqDf9gLmWQael8Z/0Fhu
UvffjFAqBlPpOoLnReBG64eR014hveVoKvymifBXxj4=
`protect END_PROTECTED
