`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ua59A/1XdEI6tLZOz8z7dw+qvSdYKSHKNa9r9KptTBqS0psPaZ8rp9yQEka4smwL
l8+JwOHVu5ZB9WUDxvAnRCCeQHoi5XJnbjOwG6qYJ1tWWWfOaqWKXxUZzG0V4u8L
xjIP8GxK8NGbiHX6PPlZ00nqVcjqTwEIz+AwkTjppFIQdujBIgeJvoIAXPHwsvwR
vLf45ztUw9wp372B5t+yppL9UQy+9JYsXIZjek4+32t46z+CyUOk2LXQE/L2mdwl
oBlvF6CuAxNNqhawRLntv2tVkMODpFRXUS0dJCP99igqIHkDE4KHDnoLuWlpYA2D
iHOXizeLkMzNXuTuPDQitQ==
`protect END_PROTECTED
