`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oW2DCoE1oXGV0zB23kMikoJy5yfxoegPw1JZIulpo8xTuKSnbQZBrxhWBPOdq5Yl
fCUBLhefZ0eDxCKaGpMu/ri/QfFxMMlc52+drknNyoyEIYWIjkM7TN53puJnfC4y
ML9fUvkgVIAgs+neoqJ8S4cp+szIaQ5z1GHMFwqdrM6DcUQtLmrItMJL6UZMf6G2
sWfyMqIL4KrFttpWB7CIQ+OrfGTl/A4cJzD8Xkiq+rgGGHYeH8OxUwX56eYYgOzv
pMm5sBJyB6/hdM2uIlMZhYENWoT5KSoFoC3fR0MTTxbVQ/O1UFsykbBLSPeamvFd
7Kj7r25QI6dXRK3QkmmqAg==
`protect END_PROTECTED
