`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4/o15r+DCfHPn+Vvpp075Cy7F+z58+QivWrE8YwnF32gmCqDSAvAbVwfY4nrt7FM
HRpayH4761KH3ivL8vqjxD+J0r9eFIknm92Paca4RM5DhDf0ny4SW2Y770ZAWiuk
F4TCgcSYItmBAVxp/6DXytMxymM8gP1MQo5BXXU1BvpDqmzGO02elcMVBsK7gXLY
jqjG7kUOTagT31zQjVaZMG2r9tnzn9h0xnnxQGnMYWnBCf9K1qv7ZoeOlrP/DxXT
Ezt3wVVKHIuvIKbQczbc+sU++81ZcIezNrN1FwUphfn/mksQZLwefzrSzFZaZh4F
89O5EbCRpBaVcxZlKuNPctzEQtE6jgSEF4X0CMLPzY5fPaMlQtFA/4mFK7sxWBJJ
rjNj2f9VGjbpW9SKZIpyOjuJMQcHFI6orawNFY8Q7JTXsr9VW1+NyHkVoCgkYaYU
N5p8MazHzwMO7jkfXdWz+a9XzQ5BmzhsMoWNqo/+0GPK97teR68fvvMJfKJ5TqYx
d5DazkVUDc+HIChoU5LRMB70qB8uD2P4H8oE6sjWljay5OsZWjrSUo2cnMNgpJlP
FC6f0268IULWRMySjRr0x5eJeUzCU8C+07/J4535EcsSpwLJWIJyOYjGnZFQTdMk
7r4IllgyaX3lRstwj7f3u4vImPLPoZpidrkxEIo4Aq4H9qCCswukjgqTeyblT9WF
VGrtp/JJrjX9P4J72Xq6zZosYoCII4UewwI3L8m/We5FpYfZxg/lis4NeuM+RAsD
3x5ZzfWZ1papTTCDhL68Ig7UhZSeIjd8CCp7qU7SZqZkTTlM9KGsAxmmevtmeJH3
TdD1oOtPZBxqMBO9IYPtw7z8IpZ5v+nFy/88gfT4dWPpBc9x//FknyI5A0gNSOZI
CVZ+RaT5nr+qAZ0eEqq4Fwc4F0g6qXB27tWpOo6ip2C+fAk1LyGdjLoTqqDpJaXz
kSotPsLvq009v4xnfuhfMiVVDP9gI2AZawvbDgK8pdtFhf8qpf/Cv4+YgLDnx39D
DaZKI0Ha7mUfcD/3MKcShtnWZfNHchmZchnNFPWq5JWoc6Sg/AcJEi+vwuVgJnLc
PLCYDqPAAXH1u/I0kOgPCm2PF1rvkX0ujWYLOj/MNyH+ieyYuNh3SqZx1erxPymV
DIjHewXw3HDKoWrW5eG66vqzNDlk2AZGd3muAI4sEXGtTVdDQ4Sfka4St/2WGU2T
Dv99jya/M9c2rFg8IS9jhavHZY9G2kbzPqPcetrLnZYgOiAuyjMKSr3oSOYBduxT
jruZoV6k4eBSFcC56JyZGlXgpsiLuKLzVf8Js/03AjIGWOa/MB30hArAOnZw3kHR
XpAl6IiQutGmG+0YeLlhLn4M/LnMELuoZAeZ+X9ZwrflEOgihd6t0WZnU82vfmuB
ARcG8U8xCpQpwQ7gA8pEDRdHhvJU6vvqIyygZdeIxiNp0hxJuCWCHxmbhi6JMLTO
xm/5l22S7yuL/kA6bGenYd6fR7VsECZEYasEzmoZDcIZ7asaw3dsho3rosxIrJwt
uJ2q1tbBkYI7fh3f4reMnzP3dA6O3MnNRV3Kiuy8Z9TmUVv1enx3LFmttg2+8Wdf
ylgcmxubcoglSJr1bVEQ7e8E+FvNkTgFkpoQodMolYGhXHA7cjJQLPcgP8Wg1bCs
/tPMXwGJMZSbLbiIV+cMR+rje43I04QOu54EYbGuqMYpY2KEO16w2dMWua7D+4sD
YF2s+I5OsZTutkf5TcHNfqxlm+ruZGkYbmVWPDu2aVczhE4U5ksalI4QPABUylGG
rnLf6SJHQq50VUIopHBK/PqFQKdqof9yVBNAqZbLf55GdY0a9Qvme+AGMuGiRhSx
2R49qHCo9sMqiEd6Gd2njNxOWE8QFk8+4l2OEZsyOaHq7MYC5X8ZZOBIcuACr27l
fkhXVE41NaI+HB2x7nAqF0qWM2Q+JDXkcP2P5CBBkTL8OQgYVUUqzIDX56dKOqn9
YChUHFrpBdwvijUWfsrAZR/KUq3s1DwqM2yUF5RjZcb+59azZV+IvJnkQU8L1J96
aOFdmxc7gAfaBep6LtypqXY+/rEWc8SNOqsptwvfYVi8haPMRRC7JyJhRuUdAJ2F
ajXGGi9WWVRfFjPzeCXRgYRpefzE1vioRUzcr9woixkvdSQ+csqTwrDzMDBdxDDk
wNf7cBAlMaElZRgRlNa31xSdION9DHX/dzokUVTfZAVl1957cwP3WArlHuStTo+C
IZ9l97nYyMcn7D4EM6jadk0xgK3f+pqEye50NDvhlky1XHpV/l708+4h/NQCRYpg
kvDFFimmUcWeXDUE6c8VpfMvpVVzs59zFFJax45hOWudWpA2DSg19gyxGYapvtdS
VWYLovxMpOakGFthBNiQgVFGZA/WMzXXFBYE2wHln3mPGL3xlqP+Cah/+7CrR+2t
/hnBJG+oOXbsCEV060QkI4SPg6BK7vqqjH6afELitTqWycpd2m/g5kmYzd8IUmBo
p8pl8A+QJx/3p7J2r44r6ETF/r8r5Ik7xvgjRhLIYtS5RneGiDnfAwqoCjo6m5Id
zjD8fhjKRMtAHbu4dwfA0I0f+ml8H0Qic5vLvJQmQ3xH6CtVxDDPgL2950VT/6fD
ZsgbFY9fZS0K9mVmM+jMMdZKOMJvfEscmJxeK45HOunxLNtZVPBGXb3L1TAfShr8
4k62Vl4o8WpEWn7l12dvbQWSl2G+u6jonVgh35stHNnD96xlqSjCZDw5Y7xzwxYS
6uN3cf1JSSxzjE5t16Otr5dYTFvknv8yHs4rF7F5ccDnxVsaBybwPwSwFAU1b7Dw
kt7iznEk1WMvZgRfAbRjrcc8cAKv7P+npS0Z4bDkhjVTG5ljwmT//T2A36gBWr+g
mdg5jLqC4zJE5ygORy7WtA+Liu3Apxn2arqYOCnHTNOpSmCsSeJDZQlcgs6MfrUQ
ibL/1+aAKIHPcmO2qG76Hz37iqoNCSS3i8aVnUY6nFI=
`protect END_PROTECTED
