`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UzIG7udvFrqrj14qQvF+9TX9oxAGQimIktrnQmNCKz5vDtlURRWc6kTTjLMcaKIR
2wFnEVJI5MOIdOcj8qYUQ4tg9ALFtI3znP2RoHanHY8TY1iyBY88wKGlTH6e75lc
01m4zxu3zLijJW0mY9K7arDghZWMFfoOpilLk8K0hLPkgylymijzqaDGQdEkma1c
3fQfXPJpMO8RaRMMWoi9hDMM2ZmMpvaKboxcxWwrz0adpyNfyHvMXyckhooCmc0Y
XffB1IwwS3kKDmp+1c3mRw==
`protect END_PROTECTED
