`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r00ZMW9i3Ub6PHRMvAeYAle85DmKIhePGUp4pTXDtTkc6Oy6nZkO0tMGzPFoxnXM
tiaAJ0CWiIzVbYDXSy3o3RrdVorGKaCupYFM/Y49L8zHWJYU5co0kdFKsiy4Ak0b
65y9HpKWK/tH7NW7+XkjQhIo2rtVo+NFwCed0nJSTtzyODfYvegQZiLEZ63pdjAe
vxYg8HvvGn08qzRUfjVjCcgim4P6hjnsseN1c1DauDyN7tyvfqwCZxO2XWrj+upK
xA5hlyZbFpIQXWUpqWBTToMcM+enBrx6ilqP0FyaKos=
`protect END_PROTECTED
