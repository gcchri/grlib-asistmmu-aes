`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5gBVDfG9PIphUrhB2T4wy7AOLaaZotVzOXBv5LTkdOITX1czME+VG65B+Clb1r7Z
0WCqZx1g6XkztqSw5gDwWck1Sx4BUs5xXh+dXodwEc80i9NsSCF4thTcviXXqU5e
kDgCQWGxhY/M322/AxsXk5vXFKb9cC75Elk6zMNjOErGIrXJC+MEKiLlv4IKLNUB
dXbHHXRnczpKc/d/ePRWRrEEzbjoHlNJ/tOfSRc/ackF6ba9SK3dIbZD5tcHUz7d
CxC/HN0t44EhboFhzcwhgtPCzY9A/OXP0zRVJn0YgwS3AhsERTicYzP1ndKy5o5T
oIdAyi2cM83UbjXlcjX2f0yBjlehKn6XqyUoCBeZto3NHvmCrlQkFS9NU3b+/qOL
1SnFS84S8u69wugTwNUv81u7tHWn/Fsp7ev2MjcEsyiEr8v3Z18oDwUPldYJ0/4m
vkMH7g2bSv3NlUzRJwc2TNw0tcsYZTs1qxAFX7LlDqmacwjwDUxWVsvgS5nWt8Wo
`protect END_PROTECTED
