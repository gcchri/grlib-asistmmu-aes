`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2hl/thbc0Qxo5kQXge96K+Ab2+R2jd7PoFNMbUriUh2hjkkeQSBvCTD6OhgY3BPe
CEkkJ6kJ20fAfBys63rxT5Xgdn0nIsaJr9j+X0yQmIGQDv1cQyOM3u04p12vTOCY
L3bgUbYlEDziWRCyoAtcdFUuWVECysCex5RPANT3TPShhYvRg2TOgX+LRPh3XdZ3
xN0tkiUIRIag4lCP2ufP28vuaDk7f1DANj7Hkzfkwhsl7SD3EUFBnV3B8yb4H7lb
Nvc3y5yChzSGnn9YWQW3tXxQGwIM+KFgVSbdnA7iTXQIaK9G6j4x3UBW6vyiLDBg
gPOi7dZe2KJF2zgxuGAmBGvOeEc0Dl4PL/F9T3kVI7Lxe0Gg0fgLwfhHY8zoYGmN
lRk6EKzBsqNjQl4mtWe0wzZmBDZ0ERFA6179Z7weV9YRKT9gKil3kLzJn9fdQF33
qL6ef6gYUwlwoRfNAD6IF2QvITBWW3nFPs6DrR8eQOyckDv526aX7udQl4UegntK
+04Ama3Rb921e9NL0sH33oX8LeQAUzM1W7pph4G6NzP9bwKSKLgG1iIAWMyPS2Jt
7HvSOk3eydck8rpAjnmRrqnBKZSojMDDaTfVHPIVNbH4jDziZrdczNtVE2VAMcej
sPTcyPjiDUnVqOJP7WBrlgJP4yusxNyQT5chXwuFqIBgSnFrgEK9ftttvZuueQBn
dt+c5wzdtC1d8FEJSQxAE3IAlZksNa7tAwi7ROIbeCp7uX4rUFG84m7yRtahKasf
Mo0/hC8+mfJd3G0z8g/PlUB+uBuRew2/OCbwCgObpullpPkb1OS8DiB5z8H6ESIn
vHdXWq7DGyxgdjp6bkIctQ==
`protect END_PROTECTED
