`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p342CWGeyA0h6IGGI13oLJxBOrRX9cgmIf28P6wI68gFyA/s5SXYU2Q2Xxtgv55g
mmsR95VqfpccCFUmQ9/2eLtH3IkhdmO2MTLSh6pMBBfmJmDS95JXD6bp8dyz2QQH
2j70AdLmBbuK9Awa5DjaXQ9yvodsCH/dJMPoOZ2WxVUMedAUYj6UyYUVOTFvjRYu
GrJUDaWEJxrGxMzirzzdJaLTPlGEXDyHjaLR2XbKTg4nOQsT8kOVHsHcQSIXD8N+
vjFrnC6OOfECryPkkCPz1cxhenZSyHHxtdxYguq5Z0wzZUOn6zpRGhxjEot7jfJg
`protect END_PROTECTED
