`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LaV2BhPmOj4ppXSc+IqboIfKWnP3ML9AoKaWg6iqw+Fvxr/nxdbXHREw41Ex8Jyc
6mdMIXuP5cRnCtKwP4Y0kNqu7POWDBA/GExXzP8JZIKma1FBiAxNtP5E9YuwQoMT
A1F+QqQjtWZrtuWoega1oDjkP2N9WiAh8Ta/1c8iVGHGQXktG7YJmDJa6InYxWDf
KXKdZjSM23+NckJrNzJbWSI2Zl4yLiZ0U2C98Y4lZpwp8JrV7J63t7kjNF+K3zcR
76syoOWSLwutWCMBfVwCXjTc9txiCjKoDyVQcfy7DYPufkhuo+MwdyFZX4r4A00N
se/OfJKZ1z5LRIuvZI3ckIbRISqwwjnoJHwdyJxOmbG4YI/n3x2wD95pDl9pZLh4
eaqBd6e53U8yCA5GpkbcU1I2m0rKMT24nuySqeQDAz0OOta5LLOVuSuCKmq2HVgF
gdT6gz/SrKNlifReccjINm9cHVaysh3jUFlVdYtRWQBSb6Gr3pZ0JM41wnMIfGTO
RlijtSPQg8+iYG+KUOqcD5H86kV9ux2nvAE+fxwaMmqsJBIGnilf2AaQ7uWrW62h
vGXMsZ6n5U1RHfFLrxv2VATvI83f/G7+rANJ/RlUw7B8GW2bif4EbxA5Aw9McpfV
WaOBCBmtKcU7BBMh1O/74gMbQ7iPVJQFFqqXSxEAdscoQd1kKXwku3HDm2dDhyot
Z+f4MSlY6H70BBvTK5zDwVVoLfKuZjS0YJ8QV2uQMMvzvvfSaaC2BkRuWllzWJut
zSNif6QAd3knK7iF9BeFLoX8tb/DsVzrmqEJqUVgXbi5yyHw3dOxcm8Tw01n3Aq+
VRFReY854CKT+0ctbnTl8DqV69bhP0APZPMv2LMkYRV9FYWsfNBMhNensdQ5kw6f
bDUm3bIFTv+2yTv/ICeEkIYqjwFILo44B6rRj9BR1bG6jzrn+OJ7azt3BXPw5NJt
TGwpZBx2dqwrfAqqcUbOZT3tOXrb2mZl+3iwhwxKvTH0eXh1ursu0MjTIYOawQwS
a0jIx6vE81Djz8zggW1CWA==
`protect END_PROTECTED
