`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r2b39xxamys7nL4GlBTI/LaRcCTGoedRdcgsimZXM3LP/obZh+EhzxcPtWcLB7YA
2OxyQsbWcARLZQZGCoIBeCcu4bKa/GTGAbdF3onemP38o1cUKGSHM1mQ6g6hNp1T
4a8IIbFJBXPHVJufJW80gxKEmSokMiZMCUZx6hDwFi/kT/jsWK7TtjGGqqRETyhX
72ldMPgojtieYGAuPN7A5s7PxlewFLcXBEdk2CpWq52Wwqa+tOw1U6cHzKmIEFjj
e3/F8SlqHZcOJvc2mym+VKp/p+2MpgvFKDM/yoOccrkyLYOKI93aQAyo2XLNDise
1kqHN+lmfjxCixeLg7fwBf8+zI/Hg7BIif0kp497jJlYjevTfy4xtR/piojTfNnW
KHYlqLL1gXJSvygIxZCXRczDsj5pdVPb/REWZYbyyn9e+kNQ2x0dcLLaOOXLBXh9
iFg/c6YO1qMaRRRurbwrk0sEye2CiG5atk53XG8wOcJXvS9M84WqIsLMX9gKp6lv
RYtHrhVd8BcRtFpQWyFx3QnyboPdmpt2hv37dEhd1dJkykZ1MfzCM6BYKWfRg2Do
N8crqNmkw/k4K6xnUblhDHUtX2Z0EhENNCkz8vrqUD4aQlA6SSnvXssbiDdG+d18
NB39Awq87yvqcj2F4PmKSvj6tWK9mE+gWGyjWH8f6bddTxiptulXznwiVJ48WnHe
SySaCn1hrSJDYSCzt4fb4QALA09TeheW23vEKaIXOCDvb5S4+xVYerd+ge7Mi1ZJ
1nzJ55jwS7+DM7QNXqu/xEqzZs7J4kKq5nI/PMoe7sIhNX6JIv1DNeXOiVhzmpK9
eVEXQM/JRX6vAPVOh5YeMQc75/DxpndezdR/XpMbOXj7C5s/nVHE6Zl5GogGwIBn
A2SZp+mEl7hFg67fv2H025MCdUhYPbaawjmtPiQlv+LwaOgeOfyDdgsTtyd2Ytn6
32yEemUWsUZrPrJRI9UXqa/aoUq7osCgu38o5oxAQXD/d6XPO8aSF2sui8f3G4Ds
dYyuAoQd+ckPYddTz6UkNCZ7H2ph19+TYPS9VmKNQvk7BnAuIE2f2PXHf3AVN+9a
3LQda7zVQAxT3zD3cyN2Uz91f+1+yj5aij1T1GwnW+g=
`protect END_PROTECTED
