`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
frNHKjUjPw3KKKeokvYsPNcQXQtH1G9Tt02ab9yef3SOH7xCor98dONrPdPmRTfc
6n5ObRNNjFp7NBcNTjaq81XkzsR9KzLZ25dXBhhuzBqUBbFJc8oXcTWRw+Yi6o3M
pJ8+ziwsbWEOXha+/kw9cxRvTFRKiWX9+PEDLZ9WqhAO21a+rGiO0uXxh8RUzlp2
j/PYEPdqoiGqb7UeDfj4CTQdKH6EEowp6ZxF/BAupCayn3VBR1PZsxTIIeu+Fvbj
myEPXO7q5td2aPs2zcT8+WXKe1nqL2TrDw1DuiQO+kLC8aDgy8iNRTStj4IU8ThC
yF8fN47e+mWhJSx31bifVZWklLYfllXow0TMsxHttWJnX1yKI0igq3D1G5VX2Ous
ABJ2Y/p3j5oQ8SIQMyz79vxDwsQbzjs5DevT3jUsrOX0f3613RvU5aHjHcXn7J/X
Ww3dCyIqk7FlekCTVCGzqsju5VOF/KDShkS1ypVsdpUZkeYg+1QY+b0HurJdD0SR
Bqu52ubW3dYZ+Y1tdkxeLJ02l/A52mYHv31c7Oo8YL7vyLUsaMP3azAxj4+YVX9e
2FKIxGCFLxogx80wiuOkv+9z5p35Kkvitf104wrdPi8IHkgEE1bBFOEfUDu288oj
I7MSyAuKeKYYed/dbp9TK3nLbHEzv233PgTI5LlIoHEqFtVvHkGNa9DdVwh96uiU
uRnwzwXG5LZu1Y5WuMsU2xPll0ZpxxU4Q45Fq05L0VZO6cPxS1upjMhLf42vhaVr
XuqcuMW0VXxyB7ahjxc96Gv5QMlNJ1CnGBLumAJ3Inn2iA4i1OUGE1flgCuJ98Dq
HZdyc+ms4GDcTHq5oLHLU29aHB7Q9xal5DyqqwJixYfEt3HqluSbE6SJn9e7Us66
VtYTNKNpPMOvpNmay5TfzWwGyMWfFny0ZjQKXneLy8o2CHRwZMAuD1oswJb6O9e6
hk8CcL14UdJBDKisnlFT3dYiA6eGn/IOP0f6rIhf/G/tkng8K/GV4SZMSFvBvhT/
5GMxsYrazt7QNVoG1wvjNIdCAudsm2SDsrEvtikFq5zbZ9U4/gul6D8snHzqKNg0
xxl0RWslkps1M9r/qySmY9GQI80LM5Ggeyq9dGhdtGyM39Hot+0k9frZQ3Kwsfgt
8Uxo+xaKj4RiKUr3nzzO4JYjXVRFw6rh2LndPm0PtqPxSI56sztSdtU59USu7WQD
8txoFFPzt6w2AG4y4DT5uv2QzGuAfbCFesfq1/lbscnJIxzKKTbd219Bohsvj1+r
uGigRFj1wrSKhvDc/pv5Y+4JGXflCvlX1yURPekXJ40xYKzjV8oDuOLsZ73tDdfD
i3FIfY2uH01m3Bppjga2W04VkfL1O71DfPtIif/qSzEUJywJcTOavzdpdZecrDBC
ARo9oGBRh6PdeWupgpX++DERCThppIF1J9kPOaAW0KzTX/V0lN5n67L8uHbNAL3t
wklyL7ifAwf7lH9vCeR9b0KYjRwpYYiHeiaUgzlV8skXphhSCTwOgbSbVsUNC8A7
GMX+NSeRC0JktmrgUzMdefLsmMsnwIv3/2hPu00kRKoHf5klR3+fA0NJAIL2wrNt
0lV8HWMMVg6W3RRnm3HP9MLIDhNxW5TMj3rHoR2zqvpOukM1Jki1fp1HaMvsh8cU
D7MB2SevWiugQbdjr87CsbDf7XpDxMUxh8TTwfEEVnodmR7xBS6XGer0lBt26GKb
gRqSvltukGcDB0Ax4zoKNRBwFzbSe77bkuyXoTIZqtp8bP1V03QQfxYqXdUiUsrZ
Mt0qoCGNeBS4CN90q9gaSUVxl88UWoaPkka79sxQImmKJSe8vJP2NdokQ6HZRJ4e
yNG3yggq804tQbwes128CbJMLAdWvLH3L1dn21HCRITqtiWkyfqjK0egVhPeVnyT
Zb8HJou0r+dNcd5M8X628ghkJtifFBr1uujD6eLTc1ZUIHYW4+HsHSqAjfyYHjyO
zXCg3/pyIP3wflEp4kOtqwkYEn6cpbBKR5ss5t+93cZkd7Z2XzYkdxKy3HvmXTn0
Th42rC7XetesImGqfOB4DfY5QL3eV/lgSr/dFLU9crZb7GZ4PXd1sBCGUKxnJPnZ
3sVn9nfT4BA3zLEFtVRw1A==
`protect END_PROTECTED
