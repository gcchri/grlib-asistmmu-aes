`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r4a9TLsW8NO6iGE98C2OiaZZjJPx1RfmtIJ5cMMGXsvbs+8qR77t13L1hM3RyVOz
6kn9mxaI5Cg8n7XvtR8VeY7m0/TLtpD2VrwByk+PeMi1On2kxYR5CAuGvJprVyuh
40lecrHUzl7D/v1WXLXAE7kJa1y4DimVniX55rZ57y6XJD7LIBb/HUmeXUy54heF
2h5Ho6RuXqrM3X8PSHfLeWQXjt1NId/XFw2N8iti4PGW1rd5P2Zo9oVOoCujVss1
sBILyxUuVlEcb4Rj4u67pxeyE40s7p0jed0U7agOLrU=
`protect END_PROTECTED
