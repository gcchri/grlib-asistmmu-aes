`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F/JupWEF/l54ag402FrJNx7cDbk5cFWRCDDphkPqzudDfMPe68UI7tlEkOz03Kf5
3LddOSSxN8GJFwWj2PvlLICBaSaaBN/QCKqvMwuxCszkDs+41VT9V8U1SLJQtftk
FIG7tsFOhm3LLbAPWRlhGc98OuvUwjz8YgGBCm9Wicqhnc58UNPoiKZ2OtLAassD
No+4aTJ/5HFYrbL06C11ONn2jbWQJjVbuTlrRTizqUynJX33E/+MBfrcR43vergk
`protect END_PROTECTED
