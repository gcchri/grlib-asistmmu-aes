`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3XnKWcpoGlCIHUXh7BWYrEGKuBSA1HSCZXHL7X0ylmpUo9IAJC9GlnJvI5jFB3c6
zR9Rloi6+s28p2UQCk6V5mLcJ48jV7y+2YK9SGmZMaZ2CJ69W0G4M0PqGqbM7i5v
CKYLfKnzTI3ftFCdzwW2KdqwYxBjVOHLwQqkHdHVi57g/okpiVFksEB8tI7CMiqe
MGHCUOVGbPuZSxAj5lmjVq1auzBd3yaOps+DUp/B3MN0Sm/Jtii1RtesFTN3qOxd
/ahH0x16AJK275dKKxPmNRDsXIGl5ljtWTWR4Aa3pZpRuZOOQ2HVeBXNEKvKLHsv
SYGXVGVBX79fJA6/MY931/jLiQFjptFWfgbYr2Av1nrMlj04ekvteA3KLDDtBPOl
JrUD9E9ZrSJeEd1ORI31u9Q6UYJ/4xIuy8PFA02MhKoZ+7KJ34PFHOhYTJkGtla5
cxn2i1nlQAJsEuoIsa5wCFxQP3T78GzlFk4hg0taEiitXRBVyovY6ix5brs7B3K2
Jj+lT+flpNvAzQdqtUUUyEFkA0ovmKQHuo9UyQUR7KUUJDvxGDEerHE52f9NJ9Hl
Xxd74l336A0eXFgososZfBNfBdOApTVPn8d7cx+xWjlJJnypOpNpcRHZe3DRVv5A
3bfNqiuZSZ6T2bLZWKjB6fOkiJGv3T4Uh4c/iJwWab21/oN2BbJO2zxBIN83hFDW
CX5uFM7yBMcM7KARo+DVgXD9+4yfQz3ej2LvfwE7BQo=
`protect END_PROTECTED
