`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GGc9NsO5njoUdkrJVidmA3345n2h0e0wS5nFJcT6QSrIth/U3vNGlT4w4mfkmPSZ
I/YaGXRMGJIozteBFufKDJM3SnYoUmZScB61f3PoCPlogXl8x+1IqPJ+ZekkJFII
b+/WxEWI38YACsBSAnBCpimzJN1rmWqxVTtd8+FRSZ7ZIxdt1gMJTawWXow1c7q7
LbQOvqd04tc4BmBChND1gcq3F6+WGJMByxdN/fNzL/GOnBMhOcdffjF2xs5AZdGp
DwiyeKMvHlpXbv9Wb1uj4Hw1NmBY6qzmnxXm2SmsIzmaTkfsSl+UaWm7y2Q5fqFi
jJgUjX6Qbf3JA8oRpKG7oGIwHEnrDd8AhsVbKLD6pkyIIE1MM6hcik2PtBRsaGvf
GTIEqlqPjSQF32eZNWYba/BD/FneoUs9NGdhYBkgzQPRNfcsbyNkfOvSZg/DFVAl
/g2ZrXdRREI+9tekcjOtKTGFwQkTPMkDyNTmm+lesQk6bR9SvqzVurwf1B+DITWq
uVQhD6nxu9aeCdxDFbZ3CXZUmfQhlwssfuglD93TmLufp0mM/BUUNV4gq0YE48kh
h4DAZGs6vEv/MS4WBP9xmHQupypsaOEzzcF8/1unWtg=
`protect END_PROTECTED
