`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jnRZRe4rDnVrVoZ5WfK+lX/dvCaNxKF+obxLqH+Fco0P1I7PVpBkAzqC+FoCC8pZ
zmjwJO6qbg9VWUTKZhUOulWEFUeSHmzas/1AD329c7HgsueEj8AxNCCTgM2sAtAo
RPV9fU2MYZj1h7MIek0KgFSMZaVnZ8don4b0tPGKqmUOZMLgnIwLV1NaJPfH+V3d
iVCXRYMJvbM2CQFs40hvbhAmCW4+t1ohbVTgiP3RgEGiV+ybcpSffL8PWzoOSA60
SsZLoqrNTJKY+Vb8uFxwVAXyDsjKlgTeJBCdWXSzn65T0S/HDgAeWxHNGlco1P5J
GXvHBp1EPMRJUrniKFB7a0eoZ31HnIQU+1uHwUIblHdOxbBgGBVRh6HKykOlJV0v
m0Q6TgW+W6GTRfD8jPnK9dst+XFFWqRXkgRZBwml49ERE7F/Zq47VKd7LkX0yKh/
nq/JhdwEmNJcD9DALqII22JiWFbMHHPhmstcxCXZm0jvOcoQW+26wnhPq2sohQ1A
LKmrs/UXGCUji2+2+r4UPgcmx/QRq7XCfLZQ/DdK52cjEe1JY36Yi+pZioeFBMEv
eCopHe8IwkSy+k8npaDMVxBsldaqhbmSZ0kvHvVwhf0sBD0269GQKpTiQZ7B92aC
1bFP66LhOhdrMl/nhTkhj4WAOuAdbHOl7c22q35eYEFr5LqhxQsf1YcjsL1zytoB
eMFwfUiQBhj/06SjyqsIeYO6ZCxvIWDTl+cijGcQATDM+d7aMgOncXfM+utSCwFV
jzVOi3J9/MaxYstFsVjHG/NOI9xZS1L5Unc+FK7vE8W/0goN4VIZzaNTBDBiR3uY
i/tVLw0NdhwR/cd/wHz84jjHuB89qJptjai/Vk7+9rhFMu8Lam+Xq9fT1RJ/ZYrt
e4uIVn/kLTuHIQE+Osywlbjeoe4jImyIXgWmFkk6Qdi5HXcPDG/h5YrD1hT8tC3G
i49XWpVs5/t679gDQznxhYvSZF28lQ6mYFJaj2q904tf+DyNABMGfPXhYSzMPO1A
pDXs9J2n7Lr2NQ/N+jeGvEDiyM8IXDc2dNS1NY2Jj0TciIXES5ljyjSy2TzIKr64
S1leLQRIinhkxTe61bd3Ht1203M92GzKekFkcPSO3IdC8sAUNSyJUJbSGgh6XK11
sYeNGei3ZZ1rbRCd4YcmysMjjbn7SMn86IoqtLjpMYyx49ss6K/57kGf2tvBNXAJ
coPz1T05fyRnSXUi8PXlqua5x0Ga3ORBXNUY/+KK6RN1WNltoIxI/VTuiaA1jv98
y3RCUMmFCYVBAhgUxgW0XmNwmKWz1M+s7rUR0XFXacAiwa9DOvCptL9Aw9ChWwsl
wnRUzupptLUXECfmmwrC+bzoKYFF2IadqV3fezdlCbe53IASPwux0gHHvnUkljhY
ao7vpa05XNcHLWJxRpB2sif4amdN5AHz1dZJgTkX5NGe6KB7CE3JB5dueSzCIP+x
X4Nb94/JC1JRZgRMIk6ebGFKXf8LmN8vcPjk7L3rpFPznTWVosYRSMJ4oiJjCOUV
tTkWxYuhHQEWvZ5qpp4y2HmrOFDSHOw8xch/z5Q2hiQ=
`protect END_PROTECTED
