`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f3fnSlSlJF/+Wq/RufibyAR6llJDBAf4v7hEsAbeaTZHfdo6BhFK71NhAs2YU2u6
6e+tRcHTjPsjAeBi6kcfDkPYJDFUfZLBwrNvBD2NvPdErLzhrK4ogyvO5nSUVYAS
VfHNf2t6N7EV3aZZ0ZDG/VxdJS31sm7Nwu8jPGxgmIjw5vDRjHmKT0XdDKD0awEn
hjXLFnpbg96IE/fPu8hXTa9fq6uWo995jRCIKt6ikf5DmcDKOFkPr5Vj6j2SlKh9
7BapD3NJxhWgsu+6liDfOehd357SCdtHbMdr6DV8yhnvdTS6fmr19dcl2CjdISTF
zBz3/QcLS4cfpxtIArKkCFANmK2IHtpiRQw57IMZnXwJEsxp65/kk2MexCD+bpAA
/2Xrp3Dhh6OxwMIW4HH8MDhnEsJR0yLi1XQLQ8gyX+4=
`protect END_PROTECTED
