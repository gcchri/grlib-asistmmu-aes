`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QZfkN4jabODPKZAerPujfqNQyPvl4TRoXh/7vZOP5Bn6+SmALHlPzbxIAiTVlErg
1AT6Mfjo3+0epcuWlBYKElZRSRKxyrQ53xCYQW83C/bv3s2jkcdgCgn46QD1mdln
l7uS6Zub+mxlmsbh0ZBjBhWdoAJjxy1SshpJxNcCvnu61O0RGPmW8aumgEC4PopM
oxv3tVL2uvaUjDFFp3llKHxP/F1djLFIpe+L7hFqKKANZN+x16zVRZTrEvNfK633
KdnB/C0sF6Gyrns/xfrXoCXimHV/AbnZkY011+l0EN7GTQy8TL8B8t5sapCpbXwp
yD8meW/K9VpII9ybZmScPA==
`protect END_PROTECTED
