`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/6VzKK09b7kSEk4MEDMrsiTOgfB7yL4RqciiMxhN84Zm6hZLb8WcwZkjszSUsett
NqyR0VWmDtiIOG5DG4IhgXYOmUPtuiukqMdRn9uE3MM/w8Yq9Ha8EvSA/cdEFyqx
fBM0zzrVP05xvSRG4x+d6TeiCknO2ijBw4Sysnc5KsXbV2YAI0koZy/HIFX8lg07
+S//Vvf2SwUuODeqHGMrXjrTPK5dPbRDXOgeYgVdoxl0CwVve34HpTARn5cbsDS0
Foli01G0fPL6o3GlEnZMQJ0zQdH5JaBfnzxZ9SISnC2NPBvO0y420GGnr8jYh01N
6XstD7QGy59i9V8114Nkjrph/iVkB5Dbp+cKy7PBZ5I5XaBkPwQ8byFxpVNwM1m5
hiHpXxjbPWM+dfyAHOc347mTtDIFdu7WzQcje+Y9dBiz4sF7OLR5x57PgzJCYSFg
Kt1rM1eq1BF0Gj2Gdmr6Jc1B8ePslqqdcT8Y+RRWZ5FP4I5UJ94aGmT2E7rt+uc0
Q+LEqppp4buwmMMtE95Frqru2OWAaGfy9gwM2JpldpkMh6eiQy/vxt6/74yhNNMN
h6I6TTLphS6Ag9nH3Tck2YtvH5iqu/yP19DZWIbTnuovgmm77RJehLCx1iKbVHYE
bAAdAg9d7FvuWxqfByHUeF4ydOJn0SDmTbeIlgg3Mryli2gr5HwefMPcW2gTKQtc
7tAdNMQcfMofqQmrBbUcUlVAETchU6XHv9A4X8gLK1PWvIv5v9Ic6U4eEv3eS9VW
gD4/EZduOQDu4ruD6ufNpg+qI62XaxkGdBqMJWPRijUJbk9bJxVRHVV3ZTKASJl/
jU288LahFBQeYIvaX4Pn8RSxYczaPStEA6BNa9nyQS1dsCfniZPVRPUkCYSwWdU0
k/pQ8Fz0YBb3AVhqgliq9LMBKNINuZ5DlJBqPb1af14Fbl8V4WbYUbu852gFd69y
qvlXXIhgMoK7OpBKH+FRMUKVdbcZMyufFh84Dblb5X0bRARue1UBoQRw2Nt79vxD
`protect END_PROTECTED
