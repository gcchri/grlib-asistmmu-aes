`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
34UvNiwggna1IVPWgyTgO32UR5i0V7jWHueefq/av/jYrdA9F3sZ7Xr9CdzhZe/l
hD27pDnJF5ljfOkP7w5iewSTrl3acnOWzAcpGW7VazDwml40AbUtwmvumtrKrsXh
WSiLf0wdxM4PJQ8KiKLqJt95PWUXwLpzstgIoPfRR2a3NrXnZ5xrHkzha489yGvU
TK1NW7qfrE++QWmjjVblinymhzLOk2xXE/ykB7viaAKMr5mc00dfygoMhna6n9EK
`protect END_PROTECTED
