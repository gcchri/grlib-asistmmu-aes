`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZLki5Cux/1dkgejOaOkX8rdfAv9w78FY8Jt4H7y+biUycBaGZx0jFu6JCVUeV8/T
s/isS5abiXq+YMgMDAeaQ7ACJmIQrKpduU1EONDofWNPpiH0EG2+lEYEKxY18Y49
93cOnk7aZ8QtlTAk3+B+mJ+KfotCKFPThn83X0SpXx8iRwhtNdvgEOPntekqifTe
cT0fKZD/v+k9c7jn7bT91zvkVBCIDS1jMnOyN05hgJfRFAXup9oC5X1hjp3eLy4v
xbdCQFeuFxlTB+ch18u/0TiLbYS19Uk0tdBhGGYBxOq4yIk1VdjHN8J3JTLiKK2j
`protect END_PROTECTED
