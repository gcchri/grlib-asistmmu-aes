`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DF7mcXyt1Hc1SxqwMWHfu+sD+AX8xRri1xkeUtLXFoP82XZCsKjY2RgljiX5yQGp
PGMr5ZF+7FgOcLhH8SUem5YnXiD0ZyJGSxXlnM85yDSmJbBMoONdgN8VcTnEQn2z
8I06YW6kpd/DEAliLAMEEeV3eBkQe74TC9LbdOjZNyjXUpp+pCU5l2fRU6rW/4s5
I+V/2sLIoXkyBGbfuoo+fI4hISQebzkJOKUhR+3Z1MjSRJ4ABEO4eHH+XKIu+oDm
rJU/A/Udf5X21M1ZYRDKqaYCqi9AcE03FXv7Ly2YPOhREzMqjQtvIDnXSCryAoMd
sf2+VKWBF6aKOZko4MdaEbE2XJ+xHuFOFZ6L8SkK+14FAjo/MZbp/kC74hKsRct5
b3nsP+3VtR2hCLAs06OYWKMX0mKHZAzcShR9a6/uDGRIUsG045ic/MsESSBiDlDs
N+mBmNbIi+koSMEgGIBpclca8qu7+6Ej60ZC1rVuG5ljPmlmQHiDcK3coZ5N2BmT
oOjrQIEAKgDBGSE6Uo/RU8BMdF6IhtmLkeU08opqFJs8kMtObPYD5n1jNhBabf1z
`protect END_PROTECTED
