`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T2r7Cn6U/o13aLSBxiVK2o0Up2cHgKpglBX4XhHm2+OaDPQmweq4bK9yiRUyl+3r
70N/uRHRr9J3eqyMnfjFQRnyCuIuNUCMmOszuBxfBLZ2J63aO55inS23GGrVWOLF
YwCfEsGcuzsxgP4wyh5QbvQ6o/kQ3Nx5u7Nh30dsMk++ePn60IEBi7jrfOHodseH
1K6B/0JrmE6O47idK9LesF1f+231DpGG5deRCMaKn7/sA0gzdVD7dDMNxQxO+RbE
nb1+TiVpt1XYNUyoxYyGC/JiDBfOnlpX9ruR1PZMmez+7/G6Hu/Kz8S9ro2z9FPc
8rs5rnAG+0QFhxi80TY6TQ==
`protect END_PROTECTED
