`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lgrWRXEQPj8AtwMkRAuuid8sz6De5hoK0BurQY1PWKEY0pBfmDUN6WR+lht94PDi
LN2y40R6uXGMQf+AlMQs2vh0damDWyRn7vE2vc5K23WZQ303QJITnVNmnUkujdqO
/TeIyzXrZBwU7hC0Lo/jC7y2RkqfMRI7uXYm/du13ZjBuOGSYvxTmGORNOEhfBBA
NgbJXSqUTG61op9QLeZhf2d7vOut0ulK4uMQoyO0bIovtJsWg0wxpW+/wKpe/hKO
aCd8HOffa5YMVoZudqhA/d0nY/ezWTPLHarPufXreUjUqeYFA+6hWE2MkwkCZGDb
rbPdvar4IYIauZl5a87DFXUz2P583Ykhj68mFpqvWPlpiz+FFcL1Zu1DuqJnjPhx
92NtqmxPhCvtEm/aZJCvlrZMpaXATqXbxbAraBdmVGRnZmYPQa9rSveqxKJ3D+vf
2+1H/5eXNyLuoZ01ToT8VhZY9bp+UPmdysfUOON3CvTkZnhPfRHdlBDkL7dI8Ycu
vpowRBkHDbV018pm2X9rOvi0RUQ3xNMvsgicc/aCaV0YhaLCPV6KnaHAs99WFGIm
qigusEbVBjQLtkaymZ7gd5HIJfY4jEdU9nLiTJA6zcveGj+dacf+4pdkwLyPQme+
bjFmFNlMXo322dY6FObjtRYnJAXxGSlkEY1dV5AFIgMeU96Oj3obCZFBc6joi9BR
3efhVqx4HDc6zlQ9yjJWG+eAzdsWkTnInCk79S3Yyjhq5YjjZjvS0OxiZD309/8L
pCeKNC0D3ZfUSosLowWtfDtARPFDLqNnWzFigwVDTqkAfssIXWb0bI5kWOVzVYVk
1y54+8WrukZvIf6n6/OCoOGyNLDvdFrpZ0/YUjobD0LJr+1IqVzN9PLD7GAgfJ25
iVTgJFs2F2jiXiA8SUroRRNWWvGIqB90M8+fxGviilG65JbuexYJEDEtzK7+zIww
`protect END_PROTECTED
