`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yE+TlUQoWtw7a96mG8PyBQfbm8nA3vn9CrdIbcptPkhYNUDuauCkGjVJCTc1+p8D
Jz6jAJ7i/pGFDWcfY6YKCyKbyAKfajSwnWPz1LwKjqP+AP326Dvd70LP4tvWGrFI
sP4V0fUdZjkCHlDz0nIB1tSLZY5BTG6dXv+B3eDvzW4mzRfek1faixnbvLYp8mq3
pcCOiAtc2gCHC3+FoVSxpYh9GKpKJZ9vUX5tWROeesFFDxgWGkzvl+He1Ex/E/0k
V9NMfnFyPrNbXFuUJoVhkTptY0sQ0h/1gFX21uu8weMn+KFdchPidfwrJfQQcBIN
ylgzUyEVbEhfe+/FpgDATu8Xfu+5UCdh/Dg5CureC9esPRMQusWcYEGek7xkWEPM
OxJejlK1cBmxgwtlWQ0Z8o6ihwZGYHy6BHTAdXabjQ+J59Y/0POr8GtAoLZPD+Jh
hvmOJgX1lH3AWyd6bqFTt2dJeQLdfcIthfptUHpIo3GIZYEqO18CD2/u5Q/Bt4Aj
YMYVCJi0ZAPSyfAquLHL1DsY778YjWFX3LsFnNcp3y9GOj1S2Duhcg3niYCwLQRP
/y4HNQxtI1/5td87t+Kt6FPftFGSQf7Q8dVI1YPTPKm1IxP8SpwFAs5ayr70UrzX
Jkb7zTvwb1xZypDN4vzKyXNga0Nx2yoY5fbcZT+cnUr/4M4OARw6aHBk4RPSiSkt
6qIDTRC4pm7hxN+MzUQtGAnQqKNED9sV4clbA7vqL71zDJ02IKMM3ugrl63taXA7
1Uk3/W/SSesh+yJwx8BhYauv/bdiqzh8/j2Q9AUFu6ebxR4sEP26KL4LyAYjyKbV
PcUo2ZH/PuLrsDECifDBGNhi2SHNHQI2VLqN3JMXJEDiv3veQ4JjwnUStW6qVLl3
sSnjodlLfpEGxlJucM2tybkwzz3Pc8EP3oSUH3PcEhjnAZUDlLzZ31zan5ssT9tl
vmlpXd84dBVCN9l982ObTcXKxyYsGU7RHLCifDQ+XBlZqYYV9AiSjeGd5o3+BJ0B
TgN1DCIiXr8Hqt1ItA+sgzkvTGsyZZQTIJu2Cv1kvE1pVIZzMxROw1+CUqGAFXDK
o/0WWjDEXirrn6IHCz4C/CsAZ0Yb2eyYafwTbxmvpBNW5oSodl9vp1xuUfadzzww
vjJPO4Sv3ItznhhI2N9shkk7Dbb1oOb9LEa4D8inqGE+IjzVvfdzReBgLWDyhoOz
Rbz4Ln6dMIbsT647PxDpEtNRKICA5I9ZHtEgEZqm23BV5XGCAgCscQf5tLqPDeWM
KIW7tNcxdQVODWPwOnmIw7O5jzOSOuZ5hLLAjvDSFHpuFPCwbfWaTJW49mplJ0iC
lfWHJFOCxaVKKky4ltOJw51iFMhqb76gW0X/YQtOpKaN1mMFk1nWtKvYX8sW89kg
qebGAc+zyV4d78JXHSaZ36nLs4H118s4EyFmiOLY5Hae8KyYpK7Nil09CefXJf+6
R3aRndDCgzjXN8GxulgFcf0gjFg3jRDMURzQkj3tDo4L5CYreNUqtri9HvQW08c7
`protect END_PROTECTED
