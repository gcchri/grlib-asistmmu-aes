`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HMjVbEg8RKQRncCy2u5qHF2YqyZSzlxHX3lzzZUsnwgmg3P33vekcX9fiZ9GxxJf
M+v1PhlArqlfrKste1auEMxAAqhay1LDYS7o3tSporja/o6aBKoh5Wppbc4Z26PT
KN+2PvqV/zBBmXuRlvZwj6EUftMUzibbwT8/xQ1pAXKwjM3dIA4/UWUEmhLo4PNj
hp/K5lA3bogOX9XFqmpW4q2rekG5KmV6zx1rzH+pe2Yp2DKCxTSEoA33RHdsVFcG
mBmPAOltMdQRDjaJwGI8YIMdfbZH8unu6Qu0BTPJA/lgmH+qKcnNj2+XsjeSMUE3
4VRlR2vZv5x6f8Ojtlxf+xkiSdmUE3oYxluaEBcNDV5XS9rXytPRIsJZWeqkzHrt
uexvvM0WjN1PNrw4fDJJgOtw8gM7Ap3nQ1OIvVtytlkC77jnGKy4Tu4mCs3cogP6
`protect END_PROTECTED
