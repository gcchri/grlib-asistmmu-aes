`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PqHR72qsFXE5hvpYTevnKtiNF2nSkmyLIwW1ZoYrLPmFq3FHJVmxICz8SjHUf8di
duNydPyLX3bo5eW3WPoaRwi1Jkd4EATgLMngmWcAm0Yufqf2/tsGJg7AE9g893qx
UE3bjut8t4BD2SZG8BG79t5nk4Lx6cDHiO0W/ejE/WbzzojS3/aqSLB0j1zfNpK3
umEJOPsAUb60RYG++mxo2hQtER7qkOtDnCZ9s/cw129o56ewVDvp2oGkQFLWWIUZ
rfThgJVXUrdXq4h2INKk5d8HxSEi9BTJ5/vz5c/rdDKlbq/yfRgSRhMr71PTq08w
J6WSvS9PnD5sXtMXaS+0DMwXl0Mw8etvgDq2CvBpgz5Idi397D7M05gXt8BCO6FI
C9xVJnO/mabuZX0+lg7a8eMfIqlG49jzMfvvrrezx8XSnMsL8LLCtJ2tWu2f2hLF
7+w6nlJgRKitXdA+h8LUzLufl2ioAZvu870+PB66MQi0VdLgRNp2jLwTQpMWMPmn
m9Q3e/txr4tUE2MdhyE6DeOWWWF2djw4JFMcaWb6WxLP+NjWK1P4PCZCxmbnYDuQ
F79LdF6FnmKhYWr3owZUbcjMw6tBGi0m+v7Sc8WsCjCY+cA7StImsb2VJ8262I5W
DDtQT/2qJtmFtD7+x6JKWhPEJse+PFxnlu35kWIaAEFp9TaFNkqMEGKbxHQG0tn/
9Fx5j2ye3dpi6Or7i/MILETzNYoC1X2A0uIXWsIp+5CmZsnuFoX3IwQkTbwnZCfk
TzqsP34EBNFRhu1ZehL/64V8EFs7QEKtTAOHU0rnatgXdcfTeIqgPSALh0zpUju/
Xkcd1+RNySm6xvkEPU6Ls8bGrQS+wUGXkBFCkYIgBK1YTlg16eFBaunihAtKllQ0
7+4IU9JOyc9orXQ3dQnI9N2SURueDz24JsfAXLkRZl2q/kWi3LnIgtQZeLeGVEZ6
Wof7L03EOQvgMmkKqYoHxksf39gUGIHhYjddrBjjqJhSDJaSxvEHxdPskFDTjdjK
au8MhrthJkqWo9pAN0C357i6igaaYmTPGOHNH2Z7QUfRUMKwf0vodB2zdEcEVhgF
DhMHKWnZGkL4Ib2+TaiVeTJi8cySsHd0QuVSUAk8XAu3cOb2LkccN2oKjJpLyREi
9LWuoNGFXj4BIfguFsOuprZdg/kuj//ktwftHK8Z4Afz/QjsX5bc/5bllVZJnmLE
0GtE7OWp2tMKbfJP1V9/jcXlU3y2Jy33y03IcETMMnVIOlnaxzSL/UEyIb6jWZ8g
YzSinKZ+nlxnViQbAiMy/4ZSTpohOfH6yrPePP0cOYX2huD6G4MJ8cheuCOzD0ba
Wt05mYhyC+WFD+yoOIhTvuU1yy6CnpUQHbBUvwNvh1bXnBeDqrYTOmOXb05zi6jb
F8haDw2f9iMdO5p+GnQ6O2tjIKb/Y06Infi6XhjHytJxbszw4G+QhOEnJcUy37Mg
r2qZbomcckGXLcU5rgtWaJFoRC4M1G4m9HMU2SnCDVzfoSqK+drrswfKzZPfXaWm
YL+GiPPqtvuZJubyg7i6lrtC4dgEIS+rn8R1PKF9Ca80DZ9yvWkJlLP7mzus5nYH
n522taRwPdz3lpJCtcCxqpR9vaTwUIJntHObdiQwFIqfNkgnR3c8ZiiuWRhu+6Xo
YOnvhKrXBoFq8vMshRdb1bWRNri6dGM4rUhwFLMREKj26AgGoKmd9mZICwqR0XEx
hZ0tZHN3JqpwX0qvO4RexszYtoYUmscEAOu6lzfiNBTX7kzWLD/VUZ4P2qDUdmnK
gwFDUTn5wAfUqTmtTWd6TXDvexnGKcs1aiH8YEgrTrexsHviToS2WSVfXki8nbuo
femZg9pc5pd4BdkPmgkVxfPZlKMn1AtBCkdxtejtVjRVIY8UEuwSIIszjDiqduaX
ejydbWvkx8VrDoaXhiuJ5/uHZOajOUR5aPRMCaZzkXL6lQ/8ln6JqK8eBiVATLWR
dfe6JV6nzrZJfzC7Z7J33iDAFAhNjgqRuyxi7qmFAha4euusl/zxQUmvoOmB3tVr
FqR+WkwXxyaCySOdb4k2348SCEp/Wwy0uGcHnhZWL0dcdrmkjra1YWiO6RbcA3UI
HSZs3k9d1ytCFStYYpEyX/nB3T69u4KuhQEm10ipe/dhX+gHdQ+IsmEChyANcyvA
XUSbSHlLu6dir9M6Wzlnt3+AHRMmWb0IoR7awtkNabJDyFzC0V06qGDCWcEFAphP
nwfvb+2OSE5J7MkG4uL/jt4J1wCaCHaoOJTMiAEsFHRb1+o96lqhh3mtU9X6dnux
cz05Qb1gfQdX8a1/da+Bd155v8Rzf5/DFBJRWbgBDUZdsplJOGYJMvfmp0+6sp3A
iyAFWitTlmFKkX0w8RnPqUga/w1zFQNGpQ3cIGxCvM910oLEwT1LfPQf7J2I8gmr
kcWhXUM2fbeSOVMHa9IZ0KssNqzWX7SaSaKhsOko5trT1fLKwE1TaWbS1x2RP/CS
zyk6qGkOrQpSZ2bsJ5xVkw==
`protect END_PROTECTED
