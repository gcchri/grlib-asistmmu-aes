`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UtGThJexO04PG3AWbuj+OLpMJDgD8mtmSW9MOL2HI4sThuTkN+r2CNsl3uqZzgB7
4SyPca3gwsODIfPryztiZLIPDDh7SAztcYlQp3Qjuh/ktGAajurckCanPcurGOi0
sT+hJsmDe4yyaa2i1nLM4xvh6v3gyKTksEyNROaf3u+6zcrshOvIE/tYgpxtpBcC
TAk/W7cvX/wkxFhwGO0YbYZXm6PtlIAD+E14n+sgvhzg7WZodTdrgi3Ca45YRGUV
+OuBcJftWH/WiZpLLbgEeIbbn0SND+53GF3ACLU4sBULM24Q5pGG6CVCn9BXcYmD
BHGr6pwAAKt6kRqgYDWx5YU4JbDatVkjmvDtz19LS/VIbuLiHohV5u0IBq/nc99n
ZyqQBXBAHKERb/0JOslHMjvgilsbigf4inMXRB6a/Vne/KUhaGl2/kxeip1uSeRo
DaB0SJV43VYxVj2cb8xDL9U5VeXKTQYD+Asp06hTU6kHoN1v9BpZE1s5aAPwBpOs
UAwYsCdg8De96QXiPBp2Xok8pN2iSIuyQbEHlOGpcS5B7x2x5pbGHJi7HXfUpTCi
uGPuVnoJAbdTvcsw5R/izKGD8WVCEJVLQquIadP40LpKFU7g8iFOuTtau5vO5OdG
eD1qu3VyGj4veoJU3niRpcjMp/5l8gibmkYYTflOAFqyU9LUJ+jFEAMpuJHwMD8l
`protect END_PROTECTED
