`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QrsFz1tOAjPk3qfDYIcZCWwDSgyDB15IHyI0oU8Mbusd9qyvXZrcZUKaKZ8lUkUE
vpAfvaCaggikMb3BJb4SSGQR51WZT8btjiz6/EzNBzRnTbP1p8KNs6F/AoMUxATF
vn6aP94royEqr/SXPSX35oHWVpi/cjDH74WhAJTMzeH+xDOepNqo1wD2oW00rTwY
7O+gcpCNIROnDLPfVKOb9uOg6k9CzhLlw92cnUuaU0djRWfpKQYFDXr6LmnjXPsu
Edqc30VxeQGw1t6ijjGn942HVCEX8IZuIQfNinzsOtGTtIcXtEX1SP3x8V5+btrd
NI41Oi2dGVDG+PDPSq8jggwnV2+2enWIOLJV6739JFRutvcKGSbTiwtOwPnJk4i1
rJVnV0GoqGgqfbvMPn2rZYlcZBGnXAvm93IEXQ2LhtgdWUlsKXjGZBGVy78+CP4K
yctO7WogYOhXdmZdLpikuDcM+mUgg2xy5x0Sj0Kbi8L6RI2xBuxJbDkuPfvZruGE
iNQ1a5q0bzU6homCg3/XiUS0NIPUdXeiMu7D0lRFkIW7U225ErAXaLs4h5viXMPy
5TB4DZI3h/q1fymyD/z7KNofCd0O3NVMjMMVV6XofQqUTCeoYsg+rbZim0lfNLIE
1JmowDDowgk4FC0oJD43bw==
`protect END_PROTECTED
