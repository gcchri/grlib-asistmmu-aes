`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
voKq+HiYp3iVw31QcHYteNYQ5eRNmRst98sPJ0IDZ1XYWfi3p7yEkzmyV5ni8ZnE
fMZRZmXBYr6tTK54pHaCR8dyz8MjzSqofBMa6hTvKFy6H6Ea8sVuc5FmiW3i3cUy
HFaf0L0HBE+gPq2ByiR5f5+tW3BKPgkgs4VSzDsbzFWjHMsaTHryZHW69poOGBQc
cLHNmQysTzd2i+SD78t9pyZn9DChzUcAMPSNSeg8Nmmhv0LAMzwnerKsAYryw0Ij
doYUY3JJXPZwGMSFGr2gz/dhlAnSKjP8mZ2IZlKPRNbEAtHhxX9xUnKEGvHqS3a3
Xa2o+JZCXIG7hm0sMf+79G7LReHHHPGnBDwOUbUM4BhgLGvbu1cfxawXHUdWUor5
I7W8s9TxsEFcs3rgjphTzZEeZT3QY0LJghD8q+ynqL0pjqCIEj3t9K3vhDYTMzmH
pvt/AQnVdcsHxltDZVloNbvKTCReH+Endn2DKsJ6lzIlIvMxe4/pe/ewGiz+it7H
uKMPMsnpH4OFf775LGyNExbXz2BtlOGHUXDxBtVlC3mW3MOx7YJLDILbsL7vdaP9
1ri9/k509QpFXQEAVxp6HmJ/4oZYG0phOoQG6ExIRHJF7pBlMBNxMdx43GSf93oT
2AjOtUSlLkvEdrFTX30CJQ==
`protect END_PROTECTED
