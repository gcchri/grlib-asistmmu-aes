`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/LGr+3N6I7jITJhHYx90Wj3GxxVmz0aNF9ma95FhnnVjbsbpvV6ljk2pV2dgRKJO
6tNgPw3zeDO6fIOBNYVA2q0rACrq/YTcoTlrWtJPdqL3qNLWRIlpv7bDeOcx1+8g
V6jQ0yrF//IJcKASjcliCzya02WW4BvfGgY1x9fuuhHcCYXYQZrgcOFFl92g1Q73
RTG082hj6WV0CEfb90cfS/rpIX8/mGETjVm56q7Ng0XWkeM2xsGdo1wySac8bmmz
BtwxVC9SzdYDXZAtJr4+CiMzYxoOJXHZFWzU7zP1B/yLJ8nGTYniLOLzRTbKZlmO
tZ+heZl+Mjb4D5QH6/AHVi8WzmQUIO8H2Hbn7iIBoAP8N0iVLHsjFIP/6Qd85qm3
l8RHZ9SHuRUKnmDLDKYHemEyXLf7nCfDlZC1JcR0jhMgxa6rsiKjLkQKIu10ejac
lktuLy0E2h4XbXC+HQVmcpUusmU3Q+mnqVVZB52xYa4r1ws5kxUP4rCneTXrIVeE
`protect END_PROTECTED
