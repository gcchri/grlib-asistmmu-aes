`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N3wjkxlC16OdjyayBOgclYozYod9IEJNNPublsgYqKpquV0Mvq8XWba0wehN8SDl
cgWLnfS+teIn/+f47We/s+Dhju8855goY85BT0Zgqj3i2zxfm5zpFZlUftX3YQXQ
6Xyf3VKz7zoZ7VmbOz+RLa41nd7KtK3zcuHzz7lj87s4gMgScrkaA0+h6FsbZvY5
Xrm4u8NqdbllG3pnI4stHeqItZqs/op785qJ7jTnSS1NeaRZsb3K7R5meIYJ1O8h
qXUJhVFkRLroCyhW2QsnwudGCO47iXSwlXHrkGW7WLxzGu6/ilw6ZbSqJ2SvdKkO
EcZOCmpFQAjOt3YpvJKDWFE+2h5c4ccZn/dcZb0oeVhZOm8jRFFWff1hsT0SytBj
hS831XI16rRT56h6i6Fb8Cj/+ek8HItydWAZ1JbPI49vPi5/QpE3DuRy6r0fbEFG
BlOtDQ3jSRdUQgXZ8tufq3EOBqWPwVKkbMON1uRM0Lc=
`protect END_PROTECTED
