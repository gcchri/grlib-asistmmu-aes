`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6/Xqg5UfSHfJyai1pdO1XQgDsKocEFGzX7jdym6nZ7KN+5E/+bR4+QsJDchG/Z91
r1lLAoOCO04BOkY0sb+ubIvyfN2pDn7bIyQpenIj9N+ASS/+KGpfwndK7LuxoCBJ
6r9BRSsPO/kuIvU0bD2VnVZCmGCc2/zfh8vMc1Cf531UtT3OeFAIbSHdo2LS7Gru
OwN8WYGy4TZLhNGQbcSiLsjEJPxJFrqNRSBAqbwd1GAjpjFlC/VNr5CA+o/inF7c
d2mBQp3z+hA7qooiiytTGJLfqjfK/QRKlCcpaUK1ekRGANbTg1OMHO7NguDoMcP6
oJ/WBVd7UGqM9ImwU63Ul7aMjF+MldRaOYcqIb/sCjru8xfu5waA24JQXMfRTnOg
92rjyfwYaBCctz/eKUOSwUXBXXycmOLf5YHPr+lNGvSI/1Q2cadYYhSacQO0Q5bL
Il0XlsCA5B4RK+nVBBIcU93pHCCL6dvFm+DszzLw3DU=
`protect END_PROTECTED
