`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yZnWRybyDLUWlb5/q8idLSf2DJkrGVm5L8y7HludZpz/UlB8aR1XkSVA9fd7iW1k
rC/5JL/XnUpITBejkvfArsQ2kWeV1fRdcO5H4YI+PGWH9c8t+cJfAat9o3Ih04jf
ch8yP69YxQE7Y1hb72DOMeZkz3WsiqTJTg8qZG9zga8595tgUQCWziLOKQvIBq5D
SWrdD65RGmoS63WuvdOua4DgRBY5DZ5fCfWq3+PRekG5fWMuoCkGH7KZUONp10ZO
huw8Em0JxFBmw9k6/MOzOw==
`protect END_PROTECTED
