`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ry8Egdlyxtur92RYSgub0nmVBaa4wb4ltzvS2q6cHyOyNU6X6ZenepBQhgKkQzI/
aFV+c2sUf1LERX5OynWW76ahLQruhPeEpsjjiM81+jJyoR/JK1I6LzVALtmo1Az2
DQERMNsT2xkxSK8AgEBsOnmWpUm/LztTPhgc1/71Ib7y1omhQdDHCzxt+x0gAcdE
YgrmhDJLOk6Y3FX7D6WTQysyaFiiCdcfyIbkAeJ7GwD4YvblyzmwKVOB8JPCuLCl
tgpSLCMiNqd+Yry0O8aZLMo/ObaI1nZ/EFerJVwhBCQDy7+GpkMmNiJwaAJz8l2C
LoNbvX6PCfesEjzbkIJx1syxV5HCTERNZA06UDn7HnLTodScpShUx8mxF7BwNqxw
QMyd8B7WNn0FLmC4i+eFIysKUfL7Gjf2RJlTZEN3zt8VqHnCNSo9aoMvWHriUEoF
dgBrOymqLQbSDMQKdSCKhR9p2p5hWtjlrgyBF/Z/IRdG/eYtRfKDz6TRT9jjosBq
gqdSJsCK0ql9KYNvzWyRpw==
`protect END_PROTECTED
