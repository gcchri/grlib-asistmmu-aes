`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qds5SZ2z5AB5U0moBxQ6r6N62Kvvt/A0O6CpmGjOk6PkUvjwytrOjIUNuWw8Ie3u
qCv7xHfGm1B5iSKpA1diNkgwE5aqNdWhYnP/mILPGISBSX7btTr28jboedRs2PNd
F+wI3BmlSCSm4+o2Vs9sECC/iR+Hx0R/aWlrgEEVrrXSuoX6f4u63AT53EBZZgXp
ZEuhb97KUeZ81oBf5S4i8WRSlSuzm9pc4daOjZwGXjKCy/ribJWhjM6fWbORGZVq
KW4xNduF/rXgjKxcMJyFMQfPNeJuoKbugouxYEvB9g3JcFofk49VHMFyjNWxtyqB
6+Tj3oK07Z1Z0fsSxsFdblehQOOFC7ZSX+da101o9Gw4Zi4YGzII5O1w/qhwGnGz
3id/EmnBRCPzmo+CmN9u5chIFyKYPS8wlu5vgox7a/DMpVnpvWynmtta4i8ASLAr
HVFtOXJ9VBOp9mjg9CKYmMvkwCXyjWEDdfGZdo+uj1dljo9nHAmjGBgLEk/vw04z
PAJs+QOeSSrUytXc8PzkBCbnKxI/1AYcGDuceWFYgO/+lXAvQFHh1S+3hHI2QyBi
W95Mzq8/hWS+9ZcXksKv1ali3OvFu5mblIBFmOVwreOGjSw5l9cne7ENjg00ephf
bPdepvXjxN8gtDXrD74vPaNZVPw4S9q9QZ2xLlS0Ip9PlOTcUu7H6/BPASC9Ejn2
9JQmE/RtJFaYEMiIpz7XWnkHbCQaBkTu3Fke7QdE31wbdP4zLNXTYmCOlxCwHL/8
VfyNYbOobmk5nfjTWbcNav98LdSU0/R1VkdVPOiv/jZbmDD7UHpAHqrvoU4IO06K
rOehXKSP7Yi8PVlZxS5WvbdgVC+3mTXtqPiDDAgi394CECVF45JRaNUjn8sG4Owk
efQg6eiigO3WzvptmcRG5B6KFbf/F1J4U1jxV9o2FhSsGDMzkR/ufZyvhOH/r1ZY
lTol+40J0pYkgXcej+9UV1ku/oAVHt3eELB8W+kFU9x6g+pdtohbHhsTaeTGWQ6c
xQ2EMez99m+WzgrGCDjoNCp7tsxIdyNzyIUXeHllv+KxXuPBENNjqUi+Lewpxxjp
rKoQGUhmTQMukcdtOMmNt4SrYgGI01sE091reCPIpXqqQkzCkBDtvchQVqYfAmsp
IDOSGUftPT80gfh6xax3MG6I/5ujQkRvthUKZW0HjccpcKCo5KWR6fyUjeNGrBMq
AFbnAdYtah1PjSTAW2zvycra4VxZ+ELNQKtmj6er/uPUmHqTZEwAQBiDA4K1+beI
HHn15FXIVeeItw2EN71Y8FGGjJo5HqSf6lkFk7/s085aDzWPsg2IfGn/7Wc6vSVf
sbWjNro2TjtKWJuUolX6m6OIb0qcCq/pfCXl8SXbya3ZvJzmQPlREQn/V9yeTR4Y
2rhKjSM3v76OVmuzHtxj+Ul6ScLRIGad0SMoDjSjMPaQAsIqdnBExM3ip/wfX/Ih
C5gG9M/gGW0xKUj6F/eqIzsFnskWx6OfYwkhN9jR7ZImUMyTed7cYvwWfjKGUWjS
lVSS/gYXKvD+0/h1v5KEunUYNyROHrDTkDA2nz9j9IPj+xBtfYVMimgIEaqClnWF
bJzqjqt8H+ov3ECzRh1PB9UeiwQrPN1POItRXQOp7gqwwq79uub4fuz1lXfk+q7o
y6miei8Vt1Pgft98dpN+YTmlCW9aL4FmEgMosyFrJh1kN0Go1HqFA4P+Lia3alSh
zyxRxP4Brs42JFTudc5UHD2uEIHOZ+yE1h+qyWlDzMFKKiM8Jfo3Atv+0FuKx+/p
zrpq933MYApnTXUTYSCNICepqxpQWH2/byyvjn70OQlJ5QSqM1wjF0eRxqnaQUld
EWufKMa/Lk156ieDsis5iHW9JvBSyyAkGQA6rE8RbBRit+Evxqoy116hNjeHQyR3
olrfJUeuUdJsFRjf/O/fJ/kPoIRup1mzWpNN7BH182+tzOR3nHfqG9IDe1QosWEg
mNbKHO3TaaJdvMUTvRnZn/ajGCGouiFfBeXuNle1FpQiqdeeibQuDqHj09lIG6xA
AoT6UL43DP5LHQfg06swcBdpEZ12q+TKwZqw6YX6LHUzAnOa9xHfoWaESESc/PdL
tRrkIjbWiRs4CUwkB/5AHmWTVtRKpiDK+B1dEYj4hefoUc/sKzCRuocAuHhzGrqS
6ekeOhZw3a2HwZHx4+RjF1saVDlGqMr09LrzYBVUhb7ctwq6vKZQxlYb+Z/DV3y3
aWuY7Bn6CE5A6/3pklZB1MeqDYT/NfJ9w/WrOvdGT63trgD6FHhxUh9F54JRNgXK
zsBq+8s3WOun16zBaOmL9OWEWHzfLm/7xb3XFATDJxmO9+nWCM57SXM2gvbMnSuK
quJb+AyOMDDWTmtzuTKE1O39/aWo10VAesdRnhc8F6eco8hHYTwfX8AkAgD3lqOw
ZdNWCJ+ZkaVjRz++oEYLQRfV4+zJay5Jp/+626iJPof5p9Hfw9KCOYvJsWls/nlB
Qyz/nYRsaoimf5iXFGzk608S275Utl6O4GSGHx+6ovgxTSjuOOosuFRN0/TjPGAL
msXjjS4EzTZ8dPZGPN4KBc/MISPiodEg77p+2EW6gOb8mQPCwcYhb9E4cEwbCVr1
03Rx4nojm1+BTVP1M4Hq5wodptvtEZN/l4rg6BYHslAIXH1Og25xeWOomBQmhEo3
YaBTtu8nFhc7/qB1vA+Q9QNQbD2BtVqQhvlLA+uP8T0b4nIiI5d7Cm8Vfv2+Jaac
cM/9qRSmvkZraA3HrhyVrcXTw25QeOoh6sNjmwvDvtY6pGS274ZARm8SGZC4XL8G
4Ys0mdqxXtnRUNnh13C9SFGrUNw187EkSy7sQXY2iVwUDJRwvjct+Sqjaqe9f/C2
XalWu5O27yGG+rqDKHxn8Ap/0WJzdQWqA/QuGOrALopKeR3RcrDAXo1jPP0+TtO7
4DUmwXTwFjal998kva/+oPTM3sllzFNOjorBlis3s95FEPoUaAUDipNq/4s6mYCn
oeXdg0ohboPIRlG0mwyi2F9bg5yF/uLSUqQ/2zMwSKgyqVHOrbDuBqHV3kFPc4/9
ewLqRXO+67sNZrFKqRihI4kOC5r6T6rw41fy3YtLhN1sfeNdfynulrZn05He644K
Bilc82AfayRo48kZo5JuDNB1c6V6LFV2gFT6KiRFnO1rnc4yGZ4N9Hvp2Vr5dFrH
ulsqg0legKy26OmVe1N8NnK0swl1dDDsrnEaZSXMOYiX3qPJNaAgtXi99pzrVogc
9pAMx6Va2NKEW8ul4pOZ5WWzd1gP4EuLTRlohq+8udXaEf763b0Ju3gewYUZflPD
K/1y89Ar2I/ISmT82xkz93cTn83jIwyx0ORGE6JPW8YvDWklhc+VCetG/GJFYKFc
iZfGP3NFmpUc/JCChbTGi7T80h6mOEulXcpqyNig3NGbU7QfTuyF0AWVIRYO+ma8
igGJEEkOZr/ZUybBkkyjjsmNkgiVoprYGtOmSN3iRw4ydNUEWuZcoSd8mrSfMdQK
shBcOJRPpWnE/Sgs1SNDZG0JOqfn0RQy0kuViHRhucgPFniC85jyeUvmt/qn3D14
AKkQgfDc7Way089Tl8SpCf/46h/plQ3FAv6HeMZt/hx/nZ/DHW8/GD6dG8sjf6Qa
HZw8t7+axksfv1A7wQYZWqPeFPHaO7m++JzqaP0a+M7LFSShgz3GaIOA+fd9AnXo
XM5O1WyPp+4K0oy+JzpQiI7EtjU1ANNBhzEO3oSXG2RAoaWFM7COscHDKYQfJnmM
Lm9sbRM7+wnuwmpEH31Lw+6lodNqqSdRiuGZe+NMAGlepR4nu7Ad4mGzVfEs3ftm
P4N9ZOTEAWbFRZM9XLK8q5guSUG9Fbio7LAwGGuBhkpshJzj6myUeBcHvOgf+6td
ncBk8VOg9eX165l0W3fgtyMiDSZKg4NyluhPY3+5hfOC7tiTjZiEVWOpnLXRSTz8
J4xnFvKJOI76F+jajV2ez7j/7NbipT5V/nWixf8lsbJzvZRfge/Wkp8zHFxFtnZo
dC6GfySoQb1ciEwMNg6uQJnOliewL4KEnvVkheyLCmjuCrcvzdBxys9BSgVrWjbL
4ssB1vHGhXUR8Y3Bwsg31bzpM7wWCiux9hDvx783QMDNq94cVdvzTnwGTYIaEAw9
e/YBloIuGTEkef78OGbO2x0N2x5cKb379Su3iGKLweuJlNhk3QRVxQ1iq7VVIstu
AMe2w5sLMeWZT6uS+68xUXN06HYpHo1ugeMN/2AMigOB+/kri/qA72DobWTmlT0X
sDA80SaqU4XeZAlcH4sHXJkuEmTBcE3y6GNP8KQpmgELZSNtz2OTQJqOW4X3eTjD
2/6L1I/q5V9CYMJbsIyl4/hc9PeIzCMmTnY5e2sk6olBoRvh1+/7iR/tdjnEPwjR
G/v/6Pyobf7WYCw1BmcjrMUrZ1+HTgdZ8ljbkHyl465NfVcxGl2fPpdhelTTqAdg
rwm58/vfnFqjdlYRC6vt7JzeEaSutO0VFH138UingONgnSbdBjq5eMcf9l0soInx
oerCaRrCB4uMBwCu2HI0Bt2lP//T3CXqYM492fj0M1eejKtiyDGZ2pi70eMH9CHI
huX02U7bAH/LqUn7VlxgBsoVJIyJstH5BdAte6/yYpmSZCyOUughq1rK/n2pBpld
02tYArwnjqkk3lXnZEjYYW22s90tb5MqkLGcLjhMPAaUhaz+Sz7tqS1kkNvpnjCu
rPm4Mnk5digvizLhr+qbTQUP8d3kiNESoZ72VJ7TmhvnZAmbkv94XX+QLdbSfu2V
wiIFCO7bixsdNqrc3wj5ho08Xl54aPCcIuBDGTYNKA3DO83Gx8CkuDNd+ZZc7FQS
h7c3vw7AEAv9pJmesHDcTQAmIBjb9pgMve4QnibJYsQ2fK0j8X9LpIBLvTwTQMMx
9M9X3UfgHNQh08GIpmafm4uiVNPBvtSwTBmzOv39OxGRVtD9VcvO9gtCGkwEFkkA
7sE0o2mAB3fB4zj6dMaLPgcw4o0y6kY1aaTuDyFEYWVYETpiuXC37iUMgGLOdA2V
we/zibj94SoX4PhNs9aeFcdgnxp2Z16zuyb2D3cr8tKaVzlHwK/Nzi/jw1WNopWN
m9wPVLJG2oBSi4uza6tZiaVaUxPKUFm9WJw5y0gwOH+K6g5TW3qBxpkjLaDbqk27
+og3h72RVjrlISVmx2XnAwV2PFYTjnVCZIe9L0hsxYC4AxetfpaomRBNTR7L7taM
hKEqBc/imBG74+cpuW430zcA/bDibPDbLldIdhhZhFobwFS+ZFw0eGF53kn0GEex
h3h8s98gXn8duDWGFnsFE5xsOprLDGYgEn+4eZfQ04MXi4r9Ep49+1U6Uq67/idT
sokPGJXZ7rrPevrLE0VCLkd73FVI9Vsiyu6QIJCh0Bhwm/C4R4T6OEWvgKxazqBc
Ki6B8wXKoDpRXd58+dXhfJmzz5RGgtTiJmMu/q7g/r6YnAmMpjxpczmSQHj/m3LF
OKrC6pmYna1BhDSwLot95b8byz9LKuHJ3DJEG6H2RvjxEZ7izIHrPAyS4Uyv5zWK
1VQdfo7FNQa+29MLb2uNLINU9Ys5KJBN7CttSsQ6bSZQyeSGp5/ZeNCKnUBoK0Pb
JYqyPu6tU6jd2szinqVRgOyAEZU1dRV2VX0tszwcCyVh0SF/3KTnxudhdlBjb/mG
qGUiNe2tA4voaUGlGRX3g8MHIhlRET+v5yi1yiq4Js1JWPBaM22J43RqITz9TBjm
j7/C5fkk4fNjm6aXZAsSejRdpk3pQxuGqhLi3cuMIBOWOdKGqOlGsl+gP9FWPo35
vWbn9b7sSNWxNt68NGHBtlKEsvQsxvkjbvOaRaziAqDbXbl9yKicc/H7pqiuw3nq
QKdXoCNvIGdxDSD0AFsdTtDw+qpDCRGvBslIT7ISis2kalD6894lq+hQUEtLMIG8
2utJ0pS+hPKSSV8/A1MPYrOhRlx9GE8nUWnNKL/3VAuwu1LXeVwQBqzh6sA9sOeN
ZT68VexZK07yskrAdsAVReKwWMwUIwrfSbHije/WdGCQHmsXv/KM7fHTzI0CFXPb
tcJ0axAMmFPXjkX8PoTJGsLHu6a8skgtlZT0J9imDFxh+BftgEzI9rblV3sZkQAe
f1OyhE2MClHdiTSDbqA6YNpBF9LmMAEqAm/46Ymq5ymD5GkIOultPeOxKDKw8qXT
i1WJhYM1OPezurZs85RIRktYNi2P8SZDL1tF36jBz9+Xu1KwYPmHJjoxQi8/yHLd
Go/s3KAqIe21PIbkke4bXzqLxEZGidC+Kl05siqUfueageTsDFjXbwEVkykPD1RG
x4bnZmqGFmNV7Q34/RCs5HFME98APmweDxsW+HVWfK95QtqLDFbWr/VGR06/745n
ADT5iBez3xaJs2JzdLNJiYL9PPeRCjeUudHXjP7opH24U97p1fzRjAZA92eUnCij
W3nwD1DAdmEctny/Iyr1eMjomDEtstsuEII7F/DfEobQ0S5qQP6XOd6lYwt36jUv
GG2JR1hKiG1tmkuKIFbk8Oa32KHMDlV7BIwd3sB2HMcehSFooYBT1R/o+MVQ+oRS
Xench/+isqGY64Xa+GwvUZSU715dordK8aPTR+dDSvTH2yeR5H3fbb6ujTZ+nsBC
7s9t5E7hxKtgKvBg4+vNN7Rf9s/dbDCgxMSdBWmDHj9iFm/n6l0ZhCdNh4EjjW1p
iX0xs4e7mnaCCqC7WmGi9zdJBM4wm1DBOhK+AqYgwKhk1fzDkN8nITBO1GlRrwtr
5Xu9d+D5GADn7zKXjlOsrciHs/hgpggReLBDpIPi62vHTeReUNxs7zR4jDKT/Tc2
7dbDFflWBuloGTcN+O+4rsaAU6jJifFpDb9OSoxBlrN6gBFEwjQRi7Cii2Z8y63b
Sq3cPvAOvBjec66zmKCVXhNC/bOBctKMaO9sXWBh7oqkKPPkPioO1+xrj5HmQ1Ur
EHmPEOhKV7HgT254Igw7iMouQ+Y66PhdD9z8kHPzTSmSMhX70ujebjtysq4qNgTO
8Yk4PKlQX5pzD56RgY5vbpfkAqW0Si9XGcETiOHWXbEXzzYluxcx6QFHewRUfsB8
iTBw2GmBa9hfB3n6SpfLVWM4EMstrTCAwy3Sq5gp87i0Hw3knk77arFf7bR0uX5I
MqlKoQ9xjqs7dZ9Mw56dVffbZ5Qp3n34H++YwsIBSRBaKpEUxeyMJNxV3Bv3LPK+
mvX0Nd99utBYTdWl7s/ticdPKKJx9xl4SYjLtNvaJC0K6PXhyjtDW64vi+aF6ALw
aZGalIUpOMI0OaxvypE4AIY1zdUs9NeWnzyi7W3aHgKJvXMr/IgPtvs/L0yVZ9LR
39T5KcggflbasIaWzUfQ4wi/3RJdvW5PUu304wyPWvPsSvMawcBgFDTbdF2UTKQe
S/ieZzGMKM+jhhLTH6mUOZDDErjGQVOYzx9uoAm9uecExuxsjKORmDp4puipENJ2
zzoCa+LcnX7ygyfWSR5aNbrUb/h0oHN6fFidxL50ukiIxL2BVX6Rl5nhtZ85ZnO5
WEABhDy27BH0JIW7T5s5R8m3Dv9TmPLLF38KO+Lmkptzq+qeNYo6HMu5zN+UcHQ+
rm3rkHwdlyWg6i1nQziVdFtljZG5W0dWjpiCfqIGo8PYW1NuvQ0A6gYRNFOI+lq/
6dffr0NxoSK1qhgk1jPvh8kPGd4DQCW4x0zMxzT4Jzd8xb+gU+EtjuBor4qI7p8G
U7+LbBQ4ChAWOaEf2nhQQDNowh0v6J+IAidxbO2Llffm4Elw1rm2sYXfDaRioSYm
yS9owHKBw5Rkh7rfsEPCmNDQXMgiaSPw81TXTJDss/MhdBNTEi7Z2mcguUNVV95O
6jsmVHjQdyl9YLIIfrayazOqF7hFJqvybmqlT9GDLcZMvqygwTzQ7WYFZ4TGmD2X
An8/7hj9hVWUyUwXAIXoAhx49vAs/vf82gQapX3B7mmaytItCaHzKgQM6+hvbiBN
bnxwHhHda8XR1mNg4hlOSteLxG8bHJwLWarhK/wHK/HaZRu56vuBhYk2EX1yuSM1
ByQkX7rM/FBJ9V9EMZ04bKrgGIQdA0D3F+qbhUJ7fbajQWECJ359g8uW9NzJmKkU
K9SFaxmU4cj1SN+lS3IAx3gPybwTMvt/0oRjk4WKkoo=
`protect END_PROTECTED
