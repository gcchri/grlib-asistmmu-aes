`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aC73yosUerVufhVZ8zgkfHs5RVuW7yCSBqrEXMY8o64IrX8xS7ugcQvkgVX/Mkpj
q1BHdojY/hfw+sANTlUKUoS9tjoAjEwYyXIJb8IJ1XNryVOymurXA+4rT1b6T0Oz
S2v//V1DbGB6N8PNty1Z6WGeY/vYbr9MsnRf89HmpQAR2rEAF49/0rmGVCZMMsAD
K/ypMdlSozwQPxuB+aTdeg1qQlWUZ6lZKo4OZ5ZPzN+ugwSKYEVe6IbcowSj7Yrr
ePzDDTnVPS/u5pbhXskNFRjJf7WRdu0gLuNAf/GsGRxM6qdx3Z2QBJOr3Oc7M9Iy
6mKOZCs265IeyNQ7jJW3a4L6tW1SEAVfMWzi/w/+L/k9H/B3y7TvbPggjiTDKOjh
A1/+FkVGVLXRS+ptvUnC5KhsTLUBJBLC4Fl0Xj2AbWWTa6n6/34LuVLhFlig/BFe
ceipqd0ggdoPU79XSdlefMOm7wuJSryqLsH+b9N2oDOQ705LA+YyzIXcxl+t6A+w
K7T86EHSSJFDyhhqe/T5jcnYVYGEsYcR8IN8BPK6xmpNf8kj1MAB+uDSirT3qSB4
`protect END_PROTECTED
