`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NZHooVM71KWNwiRhGcXAxxQQck88IYihD/y3eEVJ/zOx+RSoAq4ZyiHeiIXVg0LR
VTdU7+2q+Wf2OawqN118uBfVE4YLTHBnQ7GrDQm5gTM4HoriPJB5ezBwnHpXBlCT
wJ46N9z8CvK/ySeeKgUWzFbNAxB5j/Tnz58fLB+zwrW80gsD4OPidX1Islxp5urz
h8WIGN13Z9sn9sC09y5FV3HHf4OjYNTIiE8hHqQbxpiyx8D1dObTOU9+EpN3EDD7
BkY3ypRCKFnOkII+WeHbXxQ9W81ASdvsZ0BlRJ58v+GfN2IPOeHSsxkGab8A4+6v
WoTpdqGCGS2kUsRhahOehHCr0Xi50boA6fs90AxJSEFvmYIKFk8RmtUUz8+J92fP
kd0llv0Q00WLk0C5lLhl2qNggxstFcGuYEadRDHaxIy1bZ1/Z0aqy46ZjiaLncKP
xxZmqXyJ0UzL4vA4Qe4mKldmyjgQ7HxuKbLeptv3X30V6BMLNiWvX71fVXsuo6XB
m9rDsYT/Gss5zJ5xwmQO/ul1W0tI300B9cO54ttn0aXVqkjL/IxNO200fjdgcNHr
3uQ3dcslG8K2cldFbX9sEA==
`protect END_PROTECTED
