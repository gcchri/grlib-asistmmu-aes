`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Yy3zYk+esikR4F9dwcwCeqhutvRiaBvbdl2Dl5mO4ziHGcPme78aBpfVxvmdDHY
nC3dOFD0fM5thNvmKnIV9ymlw1NlqvDuIrQgYmdFZ/UXZNh1fAq5UY9ZQgjctLMI
+gxRTfVFGPDhbhMhzCtw7sojNwlBfVJTkjaRMaX0v82pyCdk5Jd+161K1PMmMZHE
rGvAksmGXfV1zRBkAtjhssqLHNuuXuQ2I4JaPhz2n/GWbp5UYVTc1FPEwBfRwq6D
OR2oYqCcEVqeoqvY0S68l8V7gQgJ+gbaH6wPsh6qKvQYx8xuR0+HxoqfPXcUDITP
/ZVCOMcbgzpmESMbyLgoGwyHd4lmh9MWxOP4HeIGzTeJ82Qe3JEStrrfbrbx4EoL
X0X8TbZaxeS6EFUIzCB3M+JjGzh8tT5lvDKUGc4JO8N2UjXRvU6kHLTl8CIgzwvH
HN8D3Vq7loaHIeZh3QU48jrUo0sPYH8aHTjVff7gZKMk6ag0Np/WdGtAxEIO7DCt
1OkWExv8RHUt85MgErLQL5+PhK08zQZA6lAqR7VTIGPZ9pni5ePDm9Dl+OvlKrIr
6srQEAYbuTHEq2pLU3pTnBEylIe7mzfZuwBSeAr9W/giPixQrpm4Y0tV2hCO6jih
EzAeyp5CWIIg8rKsepZUNhMI40ATrNMtt5lbo9mfFVUZeqI7pczJRrN7/COYMBpW
Z4XvySSxwFOFXfNtfCFQB9Lly1jCLvA/V/tz2vcEiIRy8hUSurReb27mMfPfd3V9
uXEr6cpmb+U8lJWX89MUWCfXg1sfALq7+7MdUWZtsXeWuiuVhJzE+US41kB/TTtp
o5/tlUA3j8aLwwc5Ck21u5DU0IyvacUVuxf60d+fpvs=
`protect END_PROTECTED
