`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ap7LAkpjC2Ch5/Xk6jZ9XQ/89leyfsHnUw3Ial/Tn0F6bfCmAdPRAqttPOw19ZGh
xQ8MvQNejdaVQbtmSRJigPpq0xf7rWEcW3vSw2EUQMj8hW2jA8rF+9jglHWlgtUU
k2TplSmdPDENcLKusS61MAIz5q7+6YiV+Qz8LONXDrgFbjMplx6JyxqaMM8Alifu
UDKo7heYA9FjizSFQiaXF9QQXp1pfkVKzi8N0jVq5sWVyGajifN2HaBAVuGxJ9ck
K6ynW90gYK3/oWxOQI++c5v1BKSN61XDIZ6I4oTj7kGUG1qnrHKtpKodxK0nBWxS
M8jPYb5gmWnIxrrRUWbLlj/6pXXmWaMk3I58SnJJZNHKUfje9L+tEAxcLJp8T4Oi
bV5lDVgiuhEPJetRkqQlWU8IeSvBTKZlls/ELUMpKvc=
`protect END_PROTECTED
