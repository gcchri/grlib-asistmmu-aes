`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UlHi02dem0wIcABLM4z3VYAGpRyRrex6jzqiIdr4HRh8tMhi5WrLHyLvscgnrexB
7m5hEbDQcpDzpjf9s7k0eb6m1UExuP9O62+juhA6ECwk6Wi4dgM6GFmuh5cLmpKB
9mxV6dj0K2T0ICF8v/iPLHL4xQf9kolY2Hk7jya+9e21wX9VVbuDcLDJN6t6MNVL
MBPzhdrj1pZZAtN9OhDkin9CpyTZxQ8aDZhMzn1zmfxvQxiYlRdChhxqA7GptJ22
hd+JYRh1Kn1jThSJ8Ae7wmM+cGce0y7tIOXZ+t4TP1amUw3bB+QD1ZJCSRbWY7m3
t26AWiHHoKVTiq6DF6KvAfvcz1C6BTgJzHbu6ugPsXinwzhotjDReSWPWTFFjSTa
iik39izqevcg6gxMTOT0hLlFpE1TCVIhttHTEiaG6EA=
`protect END_PROTECTED
