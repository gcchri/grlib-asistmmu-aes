`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sEcjl7/RmgKxl87KXvlbAWJsiUlvwJZwmS6Fm1aL53UjAOdHAsorM1LKkFA4g1LN
37e4MKe0rdGtIMdtOik1LcZ32sN+D1B5bJ7mH/Z6ZUrCqMA9FTEEXJ9618Tu6QwE
I8lAULecs4J7kVwBHNsmGnzNcpHAsJ6ZaIHh24rugrY6o0HioF19zErsDJGPbhjm
G+XUNyxNCrGv+brz+IHSOrWnrsK8zbUZEN9v/iYs07GC6PkDwrHZN+NB0ldsw5Jj
Bk1WT8ZDMhJIWJxkr/YwYcFHDJWgEocOkRy9G+UMOyZU2nDFEFK5wLWk+EA7zSFu
0Gmkf/2ayTiRAmagj4vA5pAJ2SbO3htftrn+rzwPSBgtDBRWFJG124PGlC0QYX8P
cxXbcjYhMhtc1imrDF6BsJNEZ0XomX10lSHjMO+mibsQCQGGur8tITh8jNNjAHWW
miOI5MZsFY1tpvsfqLtKO6zjRGjHHLgZO9AMZsz/7Hf7pSy7hicNicy4Fc6rGHyt
9NJU9iIJyTQzxj0AXwzh6DxwnBcoM+/ZIVGXZ4ipFvzcqNJFkoxwhXsxiBtzEVMB
LAbwC0m+YhhU0IPCbIRq5yCVEY9gmAM762oe2qyN6kk=
`protect END_PROTECTED
