`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nxOyt6OOq4MKBaVvX30+CPL+ckpz0QHPF52krkmDlpb1DoeplmGdRHYI3eyEs5PL
hyzf929dIUo9GyWdSH3b5V1f949HF0Okrj0IFT7PRY1EIz+dXmPo2k5M59B2jG7z
RDB1cSMLhy9ZWu2V63prnmb1qS/LvXxEtBCSsaKBrciSswIoapLKAYiP0mkJYDGi
M83Q7lDahY1VQ4V+bDwFJDyQCSgSo5Bdb/XK2ROJG+x1Vn8c5gJjXwhkhoqff3z4
IJLxiQp2WF4sQf3MwfvXHFQNZgq+8aCi9/Xa+uS+Klxpd884nuLZzE2TuH844xw5
QNNi3HiJu8bhzgPPshwxhqGjCiJI7q4oQnDpmyK8XR30dPU4MUC7yC2+cGgrdZC0
cuqhT7pL+3u7S6tdq7IseS89AROca10zox8Z8itgyQU=
`protect END_PROTECTED
