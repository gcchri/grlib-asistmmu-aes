`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aopNSdQElXIDgvf0I7HFRszC42e2DMZtWStXDEszU9DQmH7DoOwpdamo3pT4yIhW
TlBL5Zf5K8kRk3CgQzm8DCDFsel3JvW6tr6wjnLVL3IjFcC1yKXZV6PDCj7qFeVJ
6uSYyz65QoWf9DBSmatZOTqdni8pTz1Hz+Dxpk2RBaw+DM5fr6mXavvFTiCrUQyi
W+NuiyuIVYRntaweXdrKVsvwP+BipFiWCDxS5jThNifz5rIzQbWRYObgCkCp0JCy
gJmiNezFg/+jgcmDCivVr8QXibk3IIYiRjYewBgVrzGLN1c4BvuVvYxl93WFTf82
`protect END_PROTECTED
