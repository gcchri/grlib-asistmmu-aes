`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bbIL8VimKBbcp+cYYac9Octz8ZOYaT/6VCu7nZFhHX6N/npvnxoYeHwe1NReSO9I
eoERfkDeovdNAJSmEVu0HI/oksEAXglx2NIMQrVFM+PFKbJGh+5oAITUMHUgmZtr
a44lUhVabNPJcVM4jy7wVGScBpNgVgWQyOcmf2GD7I+PG80ou7IbRz0ZlBEfgsJ8
LaSWLoUn4CgCPDbN8zmi+VDa5sTTAUItmHur+ds+9h6v8kTUa3w0wQFPJwrl5vj/
dGGKiNrnvLL2g/ILyfWAz+q3VjJoQduKKLaQxnK47wJ6ig2PbqvrE8iLn7vSWHsa
Kr/VXT2ylUBYyYylnXQB8mopi4BoFop21G3WRe7zzSYAB+vS1q1VYEDlHXd4ScdS
iQscu/zR9EVxxqra/Voo6z3tcXS0iViOhqzoW8IcyXoI0dBn0tg/Cg/34FSyP1Rp
sUfisAoj7cdvksTClSI4y2DaeTA06Oa+Piq+DTtXn9IQ9clZcHxvXawZ7+4SLW+K
cAcPPl/J61Bmw9tjsDTRxnB3H//7uwh6cAyVIjdeWOQUu5m8lp2/7IDwzfsLJm1g
z4gpN71DNbLJmwuM832UYuiY1g4trGFgQ2/2FR5Mv0IhYMHpX1+MUlsatA0y16bF
lu3DNSRBSgMap/IQk5mYbMLmwI75FwRYmwkhgW7rcNj991gSDeWc1wNjuf2dctQI
tJXAXrv5RyGkQhojj9uw6RK1Knj8AZOAFlm+lYRtZiSfmhtWWtF4tk2vfPMNTgeP
09dxayWpw3QzxXOmNH9faAtXwDp9WjRxhMBODR3BwdzX7bwvNmLufEwnZvLK7Vx0
UDTgbHZMQfteAhBlR98sC75Sdl5QhakgHr/D3RsFvM77z67UTXDytHLkzjhHxtdJ
uR4ctZXoqZ8NabiyFR4SqWiJ8S2GMZSh86k6YpyJWm0UhBdQotZidig91smYFfVO
oalOYTxrAPoerbCuNw7nt4XJHqX+nAASuL1ZvjqqH1ihEMHwJ0bAl02W3grod/ea
1HFGwbugM8jmd6FYBbJhJB4t8FNX4o1xS1GIovuQkEVpvMI/oOWhEwrubLpU/os1
nWessqraRJVGTAc7smfEZUsBhyL0Wu95eG5V5gWY6eHgPDbarPf51T1FGxwamU0K
6+/7gbOUO4ZXwHJRHTntbofTAg1C983kRfKh8zSU05MlV/nx8sxIBr4N2a0pML3f
nlDM9k177N5AdUcfAoCziO7k7Hdbfr/ayNuD2cXsfMt7CRwxCbBJIduxFyQzfWJU
dMDzx39hdPv0175LXlufw1clUG3LCxrq3c3DXkBXkRhBkAb+TwkG5i0tAZ5c3RSO
J+db9arV1yAMsPRqB4bnSvTfPdFiEjVDI5E5MbwvQ9xOUcoX4LK/fMxHgz43W8p8
5tCcE6m7M7G6e37k9v5MfiscrsHgu+NAa0Zi0Ljttxwt6RxtrbTKoeSwdpSM3eo/
IY06ypZVqYvDCMqh2KPoThZSVet7O6MIUJFy4t5d8pU+vhFrAIKvp6bGXN/4nk7l
FrgHBhK1DG3pagDo/Bs5sTbv/FfU8ABHTFVANcptsZCzp/sMb8c21mr+F24WsWmh
8ze4sDuOM13Zi0qufV6TF2vlYfe9l9HZ//NAu9XsaOoN5bVds1XXDt1zCf2kCAu0
FWzsV59ZQCfG2uM0I6LnFvCl0XoEeCQMeIjVYMu40MEMNducFnL/Zy2ARfamk2t8
4H9pI/yU9Qd+7yy1J4z3iZQeUvgL4UY+1QK4sutnaC1oIRVZHihcmCzwWvbrPLu0
HotjJJP4JN6UKwcbyLdfrN1hWlLZQRfGKI8PehmAtExLoHFhmS+HpnuVefHFUZm2
ej4TbNUCN9AUEWAZNFQSfPDlFl5g2Pf59i3IWNvByTd+NKzEW1MoexuFj8mxVjWN
b6TU9PJqXTBRm90CDWbvUxHuW/cL5qhfIJNbMy2c1MCpvhGGzY26FAC5355LX5jH
2O74CZG/YPfKDYkFe757t3kINUM2sc1kmtTAd8ocO/ypuB9rG6pRstMnMaRe1xAu
76H+cx0TovO94Izzvz3t+rST5YnaFKkvjs6Kzgknjts9ZYOAVJcxCglutAF4MPYv
EiL8qqOp9euMoP6W7EJlTA52ipK/Z3g99pGTJZd0Q6p0Z90Nxwh8ODkvBjCoB+E7
0zibqN808GYaNPop987StAqwiDW8dSZ1IJ+jMtF/dnO5gyhBo2wZslX69evtHWPA
MDxTMNPFBKywm4IrdkW64sg/D4+f0NfEAupEGB0LfM010ZjiELDDGmoN1FXEsw6F
Uwyvo8XQ1un734ydGqbWHHTT2xnPY1482TAYiO1Wseco9ohfgEGHHKiSJYi+ZI4b
ivLMR5cnd978l0bw8klBKrqgjHNhQg3shtLkPlQjRN5SG6j2hPBV2j/i4h/QfvHo
GwIZizX0EwSz0X/Qq8SChqNalCp7+SwB0D8e96hzUDFxH7emKKEDcdBkYMtjglV0
f39PSKy2HAksievmXg8yKuy2qymaaGx4nzBtYpK8E1Khsdrpz/7ff3qTMkOQz4IM
b5/Tzs3n5C5ZcNr5wGOHXRB+EjONFWCPDtLDOBWIPBju92gBC6vUNmDybHRhIePa
sorYaWclXcbHoJIo/ib+44BKZ6p84U+w5PMDrQLfnnlqLzvZy+kVocl8SwMju/Hn
lyUyzLoqfQU16GjX41m0wuAcDU4IcXgnJo2jZs6IW4hfHRIwBV7i55KzR70tONeb
h4Om4b4ewwa6YGp/qqMlUf4ZirTSBT3mH3m7QBID84zmJ7iQ6olLZeL7IB5mzb/J
IgJ8axGsNv17I5KWbSnBpj4JlUrix6qwiw1WfUnEd7B3v/v6vh/BBO38iRZ+Y/GB
mbOvrINtyemvgL1iXZjCkzkS9Yuio6xC2rRWcg1U2LPlwN/H2QxMP6vqLVxDqIjS
lPse9yzAMx179AGxD5Jt/cXZZ9w1Jh3wNqcnJq9qLqhwUUGxularDGVDUug2iYAP
f4CSI82u/GwXT0PwehL7M5mYElF9/hpEE5UTPoFqntGxg5RIeh1IEDmFQ9NpRaeW
/gV0HqIefCFK+GEfWpJPjVVnTrR2voCwYbzJzjx2BzINr3veE3pyKRCaOwi5y1AQ
d6htJ7HliS4BdGM1hx5HVJHDFkOmnA4f9mYpFlS1EixA7tLv70aGYm+VThp47axb
VYoh1CKQo/RgbqkG7wqbUItjjvtaIwQwMTM6JouCAh8s0irKRLt5LoSNkewHaEog
FsabawpXYcx4VJtP48+X4Gf957DmNlFcIOhJr09f25PaIer5SjbqU9SdlATOSLUH
5E1qi4gEooDBXK6H7hwkWatITZSjAhg2C4L6XcBEQ1TE9dHra566wBZNVPB51k6R
9cIsNjdwRcVch9C6Md+yCvV+s7stE9DNy/3gFAskG/FpzfdR6opPe+RLtZgP+X8z
JQ/vI0KhL6inAtNnWPpZ31E/lHwr2G3bAL/gv2V1wBM0N6JoFFYAarByL5EqBv/3
ss27XFPxTIBlSetZyNaVlSggjebA/SxCOsmkV5E7w3RMfMBH6FTQ6WUze0TNDAGj
YsvIqJ7Sy9ZM5m9tOR7jqdC9c13YI3OT02u0QIPuBuf6uTD0H07piT7GA7LSMaj3
6xhdT5wytGpOQ0BKYT4opvYR1QtshY0iJewBrqQYflg5y0g7naFsYhxtQqw2wFnh
dQdZuw7h8ZZ4C6HrbksMh7qxJlF7Uu+gRXTQJDswZnqpFukVESLH0CUt60rg4HMm
sfwbtQIDw6JvfJJT4XdHoLmriKO9KOgZ9kDcLoSUWWziBqPm9ndonmSKc+PZ51EJ
qyKw7wIg2aG+eyGZg8RGtXSgt5e7EpmF5eKiM8cPcV3JWQ0ziV0vEHsEOamdcfPS
d7ZwmiSh5S8QjljAIVCMqCWvvC91doEsBskZe8/ihj2j89tjO3aed/as4nrw48Lp
w+lZUDAxKhJeLzMjK7qgaPBQhyOvxXeZHIDpJlnmo/uKf+CTsEBp2llzG9oDnhAT
MVcCmxMBpyJY3gQQNMl+Y+33Q9U8fdkejOfG19O/wBcodOT3lm0zdcxalhVEcDy1
MQ8mljbmzts2dD20THSMs4GB39K6/guAMS34lAWeXsS0JAFWHHLqZI8SVpeUy8AW
/zfPVaCK05OSYao7e65WJSqZDnPze2hOuxG/y4WFBs3azNXXoVlwVzpFQUH6L1S9
k9FkTaN52hPIYnMgau3YZgl4Wj7fkLivIevy2gdqRL2QyESkIGizppljczZoabIC
amBJT90P6Gz5yhEMoI8qut9AesaXxDs9T5AecBtTaQVkzrp5h1ATbUHEXd3Y6iTX
hL2paNZTH4oUCtr6vpw4yD3KDZNHm7ofuubdT3klqhcjylW9/k1zeiGezGC77ugp
NsBSO0MQRYz93X5Nl2t447wBtRm3Bwr65ltLt1iYATjK8wcm7+LExRnbudldyUA3
9WTClbjkb1lKUKUIjfyEmmeyixBpu9qhbDkQei92kKcHDYcnETQUiGaVgYa3Yl5x
TkhsccVlOdKOzaJ5CWwgD4U8bETIgvx2cVd0nypLVyZp3jIR3VfoGuU0P3BMCCGp
EYmb0eNeyfuTh/Iym+isaAmqWoARwGBEaA1t3b7KtpO0peIzSayANGIKRF3BvIZS
SK2JRLqMXDWay1zLhzedjYzfDCCXk8x5VLhJQN2cBQJDGT/dfWG8ZJfie9itaj8T
DAmOnQTdjO3MtleB8/+xPY2BocGbadqEZrZopwiugoY0xxkIhTPyNAeFZgklPoP5
rNQKc6+EH29GjaRZC36tyV1pn5I9Waa+K1n9CSr6060LlW9nh5RaG+k0MjZbRU9V
/vcrPSEXuY4QJUtgcYddYPnrN+C/NnjLoLwxVd6uct971E354xU1dpic1vrJ3UIO
xYDoWA1JEzd627FDQt9b18UBfXbxc09Zo22+GLDvGxrgbjTV4l8I9cxAFLYfv5U/
OWTJYWnzc5sDoXc8Vp/bQnRwNWMD0Gq81BjWVW6EUyKKIAjyJMTOvCr1HFMcpXkJ
6dP0XC8hgIc5iGLK39KtGZHy79W6dXxYEWWqPqPJvA+dlZC9rmp2VlXEna51HLe7
EiDuUvDq1Xc2c3F4tUqE5L2z1HC4DAJT9U0LA2ZtKQWuNn1e4/3+DViHPBCTicSs
vkSiGJ71iN2TPFP8qr8/xNxcV53ftn80Sb6yMwCExWitjIA0LwQH94xOVfd73Eq2
D7xM9hJMpZFcOomMP1nuZBVg9l8L5R+Er8Yj7I4US3qfadhGxHuRZqwZ6oTyk4qa
z6eQnT5PbTECh98mDucGuM9bLn8IuKYixrufIb746H2tbtDiLs+CRZDvuA+CHlx0
ypsr8JHi1jJZUR6OixvSdBgi5xuHrZxeUr44wb5NJnvNyG2aoKMA/UB+Qr2UPqWG
ceNSBKhquKY0Juk+riZEdMGhfz0wDuVcKKQlYJ8NUOL0y6V/naSp6HIqhsg/RiXI
+FiCCISl2D6W2mybMzKLoDF1xVKb1C/f4KkhY0hzLzoaZu5NyPXQPhet0n7UPI4p
L1SiqC/7psSpY35P7vTXwEQ05Le2N5pjdlgxS6/GjpjzKy1s0cHovCNOjqnsKa6f
qgJjvnqVU3NvbWq6K8oGYYrWtUVBRk7I3EvP1xvpj2SBWNBBzrcI+FTqpowsq2KL
HiiHWosIhUrd+TdpMr8UKQmDmPSylDZJfQKN0sXp7of+LwWCIblH0icbVnU4kgn8
tQzMD5o4XpldKHlM59dZqcJ7uI3Cxy4p5vfWZS3rcaxRLhLjOPR9OF2Ck1ojHx3P
BakpDY3oHphBGp+Lz/jf0sO6qPhwk+QVZkSrF10CuFIXXryjUKoAJl9GmYhVU/9Z
AR2OIZrIvnzsVcDXYwsa2ATx3Hd5lEmtgii+HbqFvnKUtlul4miX0+quaKQ6DjeY
OVjxpcsdkzZph6wLNE3d4nDj7BNqzrsEhBN5cVQFaN28lIi28ixVCIdmC4Kynx8E
8f9p8N10+ILvAAWceV/4fxD3+0DQOhnH5Nht0+0uWRX0q00y1j1BPbszqxs2z7UG
gJ98fAFRJooWQQtSn8b2yKGehEjpfQD7dvUVv4T6c23qqB+fkHZPqf3C14YQ6CJy
rcNy59TZHdy1tnZQGvwLKp3BJKJgaD+cSUIefnbnDZYh0BN9EnnLhCpBEyTA6/t5
06+DH4DSTMxSdRZb/2J1mdFAQlpmE82eglfOvCN7JuG+3XZle0PmNPxakEb7RMvy
TLW2UnLxVtyKFeic+9adAjIB3H6bVTXdP+1hGEsPft1prqXm/oE7JRPbPMr4xDkY
IhtM+q9BaZvA3aeo1HQMANMgko3V1OHSWht2ynptnhkQ5Yx7a4KOhOr+/wtfLn0t
T5tBxxKR/CTIAZN/fuW9fz2hKJOjfwl9XgaZNLyfEiip0Y4xfaDLCDFaHcCwvrnN
IdpWCfSx4+5t2AYJZKqhuvHtFCTAWZrkPO+69eGcFNUQEk2A5Jzj6mPBaQ5nZxYs
M6neZ3haglY7r2DKtTYdVyBrgk2a5In1djA6SRK7OsDID2leQxIyeyp6Ehm4BDph
vGDSDvBQHDXhw9ryXbqwM3L8/UqOMpFP9GqZvpn14qL1CSy/ypPgVKzfRg/IRoYq
K0zg+zvxLcaeSozSkUdLNzMwUNeSGJyBz9CxCP75iKYgh4DdRaUgQGWmaqVrUy7I
W2wvZwMsGcWOMF7SVUlfyMSaKwhh8ViohGRmQs0OCz60tS0CPuwAlQW2Enm9Xl/A
fe1h+Htx0u46nJbom+GzwQuF2s8F8zWtt9Dnz0r8UnQQcnB3b1OmDLm2sIpcU13i
SAm3V/ZrTbT7S1SRFhUgtwnUVmvmR/M0t0IJ2O3t9pnT1dWXBD1ym3mpueqlPsTs
vW1ISzUOxuczZYhjgrg9AhSPGks/F5aQmf9JVMalpohVemEwPvEIAiOyb2QyR/kw
HRQcMwn5nHr4z3QtZQF1Thq3Soa4iT4YbNcNGmy6Py2TE6TtentuPVSRXSrmlgNH
I8b5NY6418Tn/IxJ/qzo8+1AD9reVrQmw2HRU483Pn3LoGhUaIQuJl/kqV0Jdvw1
prizwuarF656uDmk9MxMSpQK6jxOhW9LnXKJhk5A/3/wME3b4QYe8XMtMGjzEebJ
itBDMjWQ1gzxHQUOgqRXrWqJ3qdObIL6E/rWtMecY/ijRaEOeqRFN63JHpn7KDa1
5wcDh5f+3T4Pj7B0SKJ4NLSzTrdEtHXp07pmXzqnT7X2zeHxwHyud9z77h4D2m9+
yEVI+3Xxu6aTDVbZ2vovYDxZ1rBf8Tto6tjKkfTRaKE1PhISMsFXb3blEf9qWpyA
jeLfPkyqSRogJhRIOFRkelD/iBSDbdkRop25FqJgc6Lsb3VKyfRCi8c1cLI40ALk
HZWrFoKSYNSzzyn/rd7TO3HMrgg8CIVCDZuKYkFpl7ibvTO9vpzC/t5Tp1/kapuh
crVALFPr4Vow3dr+/yyxP5DvtGXzT1iXTMiXd8BRyZYngUAy4R0YW0BYOVsqahD6
IdcdFbG1zgPMS0Ycl9RT3uUaLEI5aKjG0Bd8rwEDVi4/W1qPdn6WcdiVqW1HF2Q9
M5BV4XAX+/60TmYGhmZkeXLs/rYnpDAhWYatuuiMpOAkGnuX7HFMeZ4HbvQw+3Qb
JUGLWnT+sXl2z4jHiaYQqSJW9YocGabbFUGY+oQIPVBrKVgn/qgQlqs9nhly0Jl8
fEooSqUdHPr/VL3A+TaNCbV6bRSbhrAaMdYuVypX8UtkCQZH7g2yGzW0JaaZcbku
OTqU4RLZ3ibDBP0+igcEn/RTM7NzMWp1qzelksKN9rMEb1SwcSjiEtAZ8Cdkooqa
JRYw3T+eb9KXD66JQyPGPr00joXBDS6oqnF0hNQpvxSwGkpYGn81r1O7wR9BpKqL
w7zFOVKDE3u/O4VLaUM5Qbzwvd54mJGFEpdJrF6tmBG0ZpnfI4mLBuypAWQ4tabS
P1cIk6CGCH1rj3O7GZ/oJPNKCnwjggbR8qB3rVApV/EnCW44Z9c2Av8b6jtFtSUR
DGRim8UFEScaYaQinz+468uDBIu18ZZnBsDxJAaK8imRzuiJfCCn6cURFHXxRvXb
WlWnCtrwVLa6D3wMcdso5PB+z/fHdtRBrCsHGDGh+RDXLtokzQprNTpGfNCnvO/r
KainoXjTuUafaPQc+ijmW+FNH0Q/G24B6fO6+286C2PmlmBwORFYSPbJA5dvV2ua
h0JyTF/KHzeq2AGmI9AmYItT3DyGp/Io9IlSOUVa8eMHrjWIwUFUX4aT0nghh0cw
cVz6Z7l0foMcEU7SZoQndodCy1mUnOaDjpHzjEic5mHSZ0bwUUXyN+52jg0tcfME
rQtxw7mKx2EuIX1fJm0BA27LFM6ESH0qyUttpIRKoN6wieb3FijuDxXRHIRfKJMC
3nTlyylpA9KvjayCzni/oIUmjD5v5br07Co2UgzVojaqw75wsVxDG5R2Z1V41JEm
YmcFpaj25XuMp87m+CklOTiVKNeTK0NHbt7U1YU15+TeBWC3qMhe3+rZ69LVluky
GLO9qJNzXEGKQXpT4T1g1hwEuDag03h9KjOq1kELMaEI6adh71lYdlUQI1ipm7ND
oji+giziNMhqN67eKnAZLst1xPGOWXYkSp4pqYTP9A3ZEKOBBh/roYiIXrcJw4I8
EZI061dYffuHzMnAlMEe/ZnfYq1MlJgXxVpxDH+h7BzjoMRatHV6X7wtYhvS1Hej
U1e7dvXjkTbJ2leZTN11fezzAQKwyGNFmtRooqd+/bYC1uwkS+6NN8lwkgg7GiST
AIclbbn2ZAPlXyj11QvidbOavRPvQpWj60nUZVHAGEIO6iWF0HDwQ4O+mnME61jx
6H1j85Zg40BtNN8t4EvYPVRndhEJtCa7U85C6MQMfAYzEcLUSVMooZj2BbFP3MMp
5rYHa3pMbj8/wZ1qYJbiz+VtICSHucxTH6UbNzB+pcL8oPIZH023w83ahT4ZFNI6
OaMmGN6lkma1DazLe60gyYnn8S4mlJ10ZMujnj0e74lbDEe5PmxjkGSmj4gZ8dA4
cV8mkQtBGo5LP34HkADmj3/LH1hnPcJ7kD+YbRRGWCDFOuNIWjozRt9G8qSCNmu5
uin6LEpAlUtN5IHlsEOVLGNkWJhJAckzq4s/e2vP9R1nnhIxf2t62qoRSMSDTX9I
FexfHZBKcVPff1JT+/YmmCVeWCYOzWxGXkzDJ70sXRpqHArzk/FEqKOIfTMZyiZ3
xpGZQcRPMw2IKTez4nd3ttf6QI0PJTzAHCm+V/Vm6JotU3PyhVHa8ubo6h2KV5pR
ZPLG5Bb52rd1ZTvWHS3jFFgv+1B7i9wJ7AlJy09wvbKJqJHK+xFihwfo/FIxp39R
H2MkOagQH1CYArxOUR+7qbYCCdRfhbeH4WtHZMrdaLW2B+hJCPoqqa60x3RJ33Qo
KdQFLA5aJQPfyiD9a6xVh+hevBiHMKpeXxVbPOToykEpfj/omvj6ZeKhp9ACv35K
0bccbWHVcAfHJZW6sh0kiiXKT3eJtBTrigRqFbzBi8S/IeiuSy+hI8XX7Ns5ZjGB
8Kywiuw+CpWf86vhR8JgIckpDU4pV61/6GkD6DascFJzhoLfUnOHSgk7HKaO8MYa
gh5Pj9NkP2SJVBXWvaq/6ZmNFBIAgdI+E1xTIEMUT/6OiHLuuTOBum7CYg03iH0L
i0yotjRS/Vo3TcZS+nBjpxXZfgYIV0MqsBtXMRB56mgpcFPpT8sICeTbXeN7ekMN
3nHbU4ZFcXk1dhAAInYlsVhMJMuKJUvxDTUCU8zZ7m30LNGgOy0aBi6s7IZNcxKZ
GSwYsIMDMwVPOXICBP0JRSEsR6iW+aP/Wrgn2ffiDNCIEulvaYi1K9GwjWJUS8+X
BkaTuWhw1/FGzHVxJwqOtFTnNt0NLC6axoPF0w3PbBdgP03bUiO+Bz4wW+XDQolY
YkqRLTbVP7NrDcOR7B7r/wql7DeDHll4oLicVNlJwfc5AJVv7Q6IFCX5mIsJF6Lg
W/j35hpffrUJ54r3yYNw/rJUrDqQb99KJbJk/dzXs+FF4oTUUPwTkDvtut0CF/Vw
J45yBIM0QAsftQ2kP9EAZ5mfV0hVvmbj2VVqXrPlkoSVbWNbiwVXLGaDDYvnXP7y
W5fYc5b5REEWFt5YpDG780Aqz/18qcGOq2pLBKEp+rO0PHlb2cI9pPrFvduxilkx
cnzLyxIszbElFlFL/f7WGSWDm2sJQat1zhIka90FPeY/v4cex6ZD56Vy/qD6Hq4P
fRULdi2QBZiazeUB24xPlAeZ+yL4xjRo4BEVc4vkwwZjLvfar/RmIR2HbpF2czew
eOLdegIKvSPQ1qJ1kBjbDtXWdDvg2g9OkXFCyl+ZSExTh9OG/pey4Vl+QQylBnBu
OZ1JurHBHijqSZTFDXAUK+AUW+MGyOzF+2FG8LhUz8cNRd9NWQj2dDfBHLMiA24C
y/PMjDbUrvHHEXlSy4FjgOrH+8IEJUJGWrWh/ifv08QhSI8fvhTqftfAKeMh92EJ
G+mSdR9DKPMnF5wyR10M9gfeA5NtVk8dCYC2VqcR1dkK5FsTrrxuQPnzNumkR9K8
BdoNJOZW4eqCIXwrBeCATDu6JP50k2UFXcnhmXTB80T9pe73KgZnVRp4AFe4xqOk
M2B8hnyXnHNh2i9oL8jAqv6MMqYJGP7GSLrkzuJgn7lIqmQ9s9bP74FJj6CSdyVr
q/sNUE7k1dWrJK5+DQRiNbrq6EQOc/gKiC/r0g0govpJ7VHZkEmmikj2DyOpPBtf
Mvq9ExyhCChoa9OrPD1CWUrygzSANym2+qsCJlW2x9XEVwP79bvuj80v4A3KX/KF
xhB3J5rzEvO4rJqQnNYao1hAbFMjNm4wNBynNhbnA5xIuAvhetIqZA1eP7JFCSAV
K9b9eWBGT+YnBU4nWdxD3bx1fWMxANoJEcp03ycWAf5meK5fXETSvebEas9p9mTf
xu4kmIHHUE2HYdsPJL6kfjP8Z9eC4aVxZUyvXEUvMxIciz8gpALzNf6dg9e7q0bv
39AqwQGhbJAIhJ8Bii/fPWCA/A5H6xWvfbQdU4uVY3/RWYMrbudhZppb0O13ZsuK
EeA40VU0eZZHq1/kUBiEFFWVW0R7/rayemonlMW/9+acJj60WbMGemjK3brwMeP/
f1VUpIkUTM/vqUhd98H7Fv8tbpo0aRrcUUkaKJ0FmRq7gtBgSMXWxANDi+jtRmK6
0iT455QJUEPWB95kkKutww72VNzmpMgyAXH8UWAmsx42YiQDEqk5DkGTG+WMGTTo
l/pwBf6ozEwqGRJboT9KBUKVAVoscVqhrtD9hotfHZL7ca3yCrOyyxQderzxOlOp
wdDhUFjmS7IxAuoRk56QjuaVmFoVldjisU2FAvtNPWDOGudnMFOp6hEj48xoUneU
6sz0NFO1W+OL9uYCNAKwAIdMWmrn8+Xmfp8Qy6b4T1hQqAevdwbETyGpTF+412ZT
Lxt208eReNuW1eV6UT85kc99RoFtvAYXcCIDZ1aNn+VKPZQkX2SOLm1ouqmMET6S
HbKLG6USsy9mR349l+FD1YIAhzLphsfQi7T0I1Ab9GqOLpRdm5WKMv968cVK9ui2
d/V1IwmW7Y9HDGFwJHmIK2Mcz8WX4g6c/pu7BvTP9q0NzWw7BYQt3moilR3i6C+Q
12FGa0MP2moZXJ1RLgfBx0f5Q92PKUh+mcqDBCd04EE98GPm/+G9mw/FEnGw4mIh
RmIb21FmqDCTR9Ke0/oL1HZFqNhmwwg3hKkG8tpllig5IqIg/+D9wb3KI3bFAgOS
Muj1KQVdnrsYJv0BxoXqX9zA66KmX8t+7oKMf8cFoi++kHLRBDtK/eUzlsLJBrwE
k1Q/j/KKRuDcbCKH6UwjBQyF/CRguSVqZ8QlvCAuhE1YFypm+EBvp8FMlCWU+eRi
P3nD08wRkDSj0zALG7SYzZfihXgKjsqxZVYunHkMCCkV9Jl27TdjQ5lGCYMvr/Ym
T1rhRWx80bRU6yA24VNs5zIWrV0YYLbCIQIFXh6eOZSqaAifo7+PFbMxdbwYeDoA
Hefo7rYBjHv/sA1/JBn1r0/uqFWD1vIyf/qDWc0ZEOBHWGbSmt7Yk9ZnxUFwfRfu
DIT8bVdCDeMBpsyHz21Rqoj4Mbh7nlkhOG2W2gtOCq/FNAVljvpxlyIiUNm71y9q
7+MJD8FUV+pd63DerztL3lnyXJrNezaP/gOLRnToC1HPckEn52BSbh/YVd+qxz/c
UBH8T2DgzXv3YDRw0blXppZgKYyvewfneglw44AKi1QMSmeE9K0rQsSCh80dTS1a
OK/X3BZoRkKnIrIqi2QUtJu8T3YBZpk0Dj9RPyUpFv3pZpmTY3CeMDErWvR6Qffr
3wjMEmr53dEiBCc8WCxdnQQVcSVIsOK3sOFFhfqdGilICinobcdkl7DmDQCdXmsY
a0zeNksccOt9ctdrRYEpH3zhkrwAE6aVkWF+RkfxB9Fu9wvEQRF8z5bBJAmLMRKZ
D/H5anuk9L9xF1gTf3YTNeW66UCc0yjuaWmxK4gYRcxiTY7eL2L8URUmoisYTdSc
k0qqDtTEDt2LlPRLFYpn0mxJ7Q1ra58GYoerlf66oS+MAUs0AEqLufFYrEohwOcU
LZgeIV2KR5Sfeus8NIvyd/K5PCLhm8ll64otzr2j84zWOK0kAnBrx72LmBKb192O
L8VtAw5EVOT2PiRD6SjbJtGEIH8X2deLBO6bwmOnuItQmLWRGwdbqXoziOVG3tx4
Bw2vWwbr21X96Mhx4o0xoKMsu68vCOGzE3TqN7c0LOVuaD+XrcWsrScT/lkZwj21
umP3nwJWSmN0KfRejv4JyFnh0vp5IO8JFUFqXrmRGq1QL+K7tQ0iwdrFcbrsHzyW
s5g5fB7qocPpNfBp7NC86DxevjHH4QLHx0e8bXnvshrbB7PgCJ1eqkZqRv4XzCTW
B7ng8Zmn8YHAhTw5kacXEgW3L6CIqOGQ2pPvkuvsIGgSM0YKVrbytWkkAvu5kCV1
khaEdSylp9c3fvqsWj334PSnxT1QGHf26WCkzJU2fvQ19BZ89FT/mliNnZVB10RJ
LT0Q52odM9+imA9837Ez4/NFdMi/J1P2jO7V/mOs5g4+nNKhphVKPmx61Tzqa3GB
nCkif+oOGBcU6tqk1xvkoXcYcB+M6f81D8OfueCNnDunVAGZfVlhfzxP8CmsiKNj
WdwQnMftNh4ZUW+VyQAbYWpvQAV+6hp0vztOiQjPLVtAMnEwiOmJG9EoKYWOKdPZ
TUEmarx6NIlTgd69uAFDAjcG26q7//UvuaiSMepmrHizEyuQnIjq2QtXwvZKNYtm
jAPsZhqRIgR+aiqPuysXaczkVoLRmtp5nTdvL+JqImXM6vY8hhjyrfZoTmtl8T1i
+N1dTA8KcgjHlMdseUvemetOnZzOmlAt0oi4e4ZRJ9JowMWUoBvT1rrUHLbBLc/l
H4Ib6fZgcIc8/4lyhF/7mx5vBDIYganbS+HzNddswRNjoQMH0kTKGzlfWYf65HFc
AS2AWNXfhfCHq1glYkSlqfCRFSrs/aNFrcN+iQ45v3k0pVuhZFr3SUSB8sPVfNIv
aCQ9UWZ77sCb9XA40lupYDrQ32Oe8D4+ARSFz1KPSTIVBlviRtGtiLZxbLoIwtOE
8oQQIJjXadG0uDD2bMeufA3KdljZaIPVpStQH6FvUWgX7fnaE/9+dwPS6U/U0fLM
yHPdgyc2HIyA9VeoUPfSPdfzwdy9twninqhELXewr2tMxbFOuWYwE5Ptc1r/uY35
VNMFtzMxHB4aJsgA7eMo+6LYURL5bOJtvGZ9ZVH1dyQCA6MsOv1uJEmPqwdso5Ew
6X0NDBRf0ZwDk6hpVyTdISaexJOwRsG57Z0et/YmmoIZaqJt7xc88i+OVGqVkTA0
oHT1IP6bcHoNNE3azzWwYRfq5yT/Jaz+earVYFW9k/M6OStUSubhbFMV8gOhoGS/
asJmmZ7jMaemwb1KnJAwW7CfiOHNoYtrhYkEe/IbgSHpQCjbE7FaDZR+ael5Ra4+
AbZfX0hxwb5vSSGLr3Bpxz1ZE37U12wHWUvcZZlPf0SyZcqTfmwoJdsRRFIutW6Q
fB4THoAhuQkqfszQviO8xGIUkp0gP+jmDGVkfTNVmYbh2EELex5rssi6tAs25tqR
+HuDHJfX7BfBmFThouldlgaho2WorZe0vZBBwCIGFrF0mt4SJgT1H+Jbc/H2xKuV
NlyyvX4KcT2W97iHnMLqtKLGr7dR8uStq3ZbvyLn5Y5W2SgWbD5VXPVp5Fc8PucK
02Sw1Pu5aKOHk5KYHvu/dwRmJvALtyCsOEmByre5dYo=
`protect END_PROTECTED
