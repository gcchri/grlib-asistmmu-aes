`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f/6SrwJJ5yyb80BRLQwcF/yUhw+Xm6Qq1KNb06JrYIPRg80f4fNucXNrxHDBX8a1
IIpLLk0e1um0+E5d86WrDxwSAORpwO2Cp54hakfCVPbF7/ICDTgLDoEN8ev7zGTp
/7SrweG454HBI7Kq+9lTXVJ67UggF2wy918/gRD/ES4ifTmq/Hf8q2nwdZqMCv4a
hDvtI+YH8I3gkjRWp4aSgNj/JK8ukF+7OhNHJkq5QlkymtjzujNSxeez48F4HcaQ
R+TBL4cG0Hj2enB1eg2jCWZSJJBEJ3yns0vSNexbxgN+nOK53hcIMpdv6YTKruTE
Yvo0mDxCz/JNAsqeusFAGccuvR+Np3dcJb3/nuzrdPi9UyAgldREOhTTCN6Oao3Y
mtT8ws6sgBd7QBCEhowCW8SziQ+2kXXJxtlA65ORe2KOHqIWj3U4Z/mny5m58GGD
QZb0QBt7EYXORR/DsfgCZGVFM2FTS1AMkfuaf0x6/kNhxT8AEPoSrFqpohgCAbon
t0A+OYkNRg1lt9JMk22GhtUCOH1KiXqr8il3rqNUQBM=
`protect END_PROTECTED
