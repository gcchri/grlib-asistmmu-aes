`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nnC0kHpunQwEQUAPsMPiWrt8AU22fryX4WQh5HuCtQL/7wM5wCADxQ6taq37gEe+
N9rSwwe9ogUeNhoqwvdVXG88iV4EHG2jXeliT3eJRHQ308l2QhHNQl2/j1TcHp1s
oPja9ygG+z6bjhd9Zn8vsLx0IOp2s0kyBkJHOhx4E8F3YEsertDKcgOZujdfTphx
0Q1o1fVE2MiEJbxp/XEqh6Lpwb5q+Bh90EsvmykxxxL8ErY7jltvrdaI78lpwIuZ
UvB72Kb7ZFrC/sc2+MMoGsThpnAmBvmgDcEDG+Tg/HCU9K4GCqRMGLyotX5zjVn8
iUP4ZDVP6r80NVUe4yidb/zhi4FnqGKfoUh8Ie71dlGneoL34FLH/0lvjogPlHWw
tLX2Y9jboinqtVuAQkWaoF82sbNXrc9l80ra7sK11dISuIq0rj9i4QCoONqbCFQz
DrhsP9HqgPW8ekynWIDECYfo5A70c9Svb4mpvperTMe3nBBW1GvCtqh60zlOkfzG
/eIolI7cVTFliShK3vVZpEfaKuKonjX4ZKlUxBxnFT638QDIyKgA3iihCl1unM6u
`protect END_PROTECTED
