`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nLUjFG06ILfQNJFjyKxRNvEpmRhUcnQa91QSdgnQmhcbPFfJHBnh5CZZkOZcgyYg
JorrtmFH4/J33tXlOm4pcCHrisTm5+VbPNvwql0aJtb0I7uwQF6D/ahufPIGgNrl
mD/0A/J28LAErYUxct7w1n8iqF+TIody1Rw3AifGKWqHt9YOya+SpgkryBML4I5D
esZshgxKtZACOu6I6bKlkxePC7kQm2bVmNtxLriNXf6mqT96UTQhbR3MRrn3dQeq
6s95gC2GY3vtYmW39/4fifRmSrL6iITR/9hoSePgk7+zGJj7QuUpwESVR/Q0InSG
6AdVj6iIq7YW8af2zxDMjPWyre9Kmh79uRswCpwLvuFekLMOxaG9qLh4fXslrwm6
uksvsQajWVVzf/a2Jtag4P44ehY5grFBby+0x+KyUNo/JZOHd/D5y0NOVrl+FCWp
0ZLGxIac+MSbXNCmGnPoRe4rdIKzjFSoRbiJJXOa7sknsnNvd5tnkyaa3VUEQQb1
QDZZB7BCApjaHlOOxu7urFSnMXInXhe9Nl9se2S9Luqn1fL6BgKrhhDXytW2b8aL
R8tK2x/ZJv3kg6P83qn4u7Pm5X0eNcJAnlkL52YhQ5vTmH2XCkU7FaK1EEk53IBW
qIyJVyBWZ9ubNI5IrAHHTMCCwP2FTihw8yMG7s43PKBefdomXCEA+Z5v73n/rwO3
WS8iFgBeEWS1b1bHggF29ea5iP1IgOJwuQKYCshiCDeAaWErRMYfyKYaB8n6Rv3N
UyLfBndeRvBy7y9p58drCA==
`protect END_PROTECTED
