`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9PYTOoxQf8TyXufomUT2JzUMZRkWvfKIU6mroL3ktydt/ywzz372n7dGyGRVtOa+
R6OCYR4CD/OzGWQ+CJAdIGcVeptS3ALylSEitvCTsergg17R8wx34Zn86CANlliY
rOv3LGtgcgiUvvIxrhVgWHajRISg11c/dMlF1skhEdAHp0/+VdYDSwcC4GQObZQU
hT+LmBPO7pPHz43jFdHnYDu0jS++wLc6AXNEX2N2uMVT9FRrE3LOrm3p8c3DNSvP
IWizlWm0oNYDX5x2gCxC/Y+bfGX/ABbV4C/2w9YlGA7kRMrPO+HHsky1V1gVY59n
QvawnlvgdByXV8426OGWWY68FT4vWAN6zhL/UYea7YZpKj40KKB8oAWqW9bdmIQW
NkODYMfKSBmJSfQbZr1yCZLvMyLnXepSafF99qDGZst+tEq7O81sfjxwChZD0Bre
O2sHvU3a5WpqdhNSVOgn/DilU2gRmbNbX6VsVVCh+IvECV01MpcRJtYpkee+Klx+
UPoYprhg0ufh2jMyp4oR/iK+nJ+/HX6Si7ZEqHMFijvffmT4AbLMK0iGdRWHSSRW
Pm2CsR8xf4ChrggQiEY2N3vVSSKNuyBM05C00wWw2qB0abrNaHVC4sPlxZ8c0EUN
4vNZinbolBzUDVUIUfSAxDr4dSuE/FeiVEbBfJfKM1Arr/A9BqulCfLAtn0rnhnU
M/FBH2HFyA4Ej62pB6UDFCqGu5WqFZZojBv32dqiACAIcQT4Jx/VbLGklJK4Ofi9
IBXz+MlG7AP+/HoVyqLAN8ZJwyCO/qpqdazZRvtobtVYz7NfTM9miWpURAbQ3X43
8YoVR+oZrEzt/mmr/DwxJe7EiHoQv2SojEKSWdM+GHYGN9DbkBgSdt+U4MqRQonl
qcyZWLttYucGka6Vxx69dii4gMBcs4YFg13b+b5rLOTDba8Nr94jgPwoGxXyD+Ey
zPV9Bp9s91TloSjNiU5ZZ/4vor3g2e80NXqLgm2hvp2V3pKO3/5esq5H+5aXxZtG
WtVh7DRwAane7mIAtvXmt6wl25A4R5mRQRlBSeA3oxswjdYzpz8OJBzvMnDgdM4J
`protect END_PROTECTED
