`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4iKRHVV+zyUgQWTAeHEFRc+KfKxzi1B8rqcf7Y4EIwen7xrtgvByOZSoi9YihsoJ
CdOeKppBDST47Y4w5SdAStddwgIenYxpLeUUf/kPa+uHF+2muidp+90KJqNuj5OF
aqGeM7PaQIQcKtUcSKbrEHz+JnO8O20L9SMfthQ6qCjA+lnjO6rGJpGJB/2Jyqvq
VbaPeXKrlMN3pNYqr9mJKF1/gcoTsxXwJVf+506jsjqqFrobB3xMR23XkZP1p+3a
p4ohQ0DVKZRPJhD866ljxEhR0mRRDVfnnHirAXe2RpYVsL9Gf+5/HSxZwPqWDlKC
ybhKZ+iyRKb6X2ByyHBFdZf7o60frJyA5IwjvEwmi7FGg82SsqpuRYsN4WrvDCpz
d3qRoKM6sswTF3gfS07WFuRKoE5wpUYV3jEsaK3RNNwE14QmCin54ZUvHvdHpWH0
`protect END_PROTECTED
