`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bD+BChb5JLFmqNZQ9OkrLZQuh5+jV8I83zpMnOTGPWRAhA7A6hKaAisnFaIOLXYF
RPcP/Mup25Ou2xsFyuRV9qtt+lvrf2CF7/AuiEtiJzFOHEEEP335KKap8/S1CjNe
EWE/wZV6+s6hwGQTUfR8rxtWLDMWV6VcwJUypi0pQGLFBvEdbv7y/f2emeubFfQo
Ji+W9IEe4Szpbr00mHh94wCTAYzrlt2oH59xbRVQtnmmtLqgDTnLVoa2K5ElZwtr
`protect END_PROTECTED
