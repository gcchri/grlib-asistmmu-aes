`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kf+SKf+2v4m3+6PHvU5cJvLyYaIQGjaERtXgEwly4gWO9r0Rz2mfa7Fw2F4c6FQG
+LC2uveJ2rvAN5TWQSv1S6OiAXEJ9t73A86ngP6pu02xFAYmWtlpJb2N/dyPgVvZ
n0PqWTmt+6XzHFF1N7EmNCzmV4v7urhrAsZIk2cxNJxDWk7Na6jlCB8+F/nntQOK
LE0Knm5vOQpbsqch8MsQaj2NsUyvuADHaM0G8EcASxfReEhIyr+SCc18d6wgNXCx
zsMxLaVCQ/AHHhb8EBEwRnA7zTSZfzLOICPymtnN+K8B0cycZiaGF8SVJgMysvOD
nKLSmLys+X2F6t0LbVvSmvHQg6UMhUV45Rq/ZZ//L4Zv9vsrkiHP5rLVQ4WafF9L
xyXuT83Tyo6WntUxCjbg9Zwu1eGT1ZsFCH3GrKfPN5Cjn5K19lkBhu7OOfEpPdKL
LAySdzggj/4YRJUuMAc235CE/OMvLsLn/rmtr0r0pqA=
`protect END_PROTECTED
