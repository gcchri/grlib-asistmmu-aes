`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MWXnQ3Gio4xrcdfmHdr00SBWSPu5hPS6n8dk+fxFFvC3YjHMRy16kKNssLITPkup
une9wz8HIGo45s/sYPIWokVYpCv3jKzAs5UuLqZOuqZmbB+NrXk1m2+o/Hn8fb7v
u0itMypfCpUejvPBAvVDbVOARoCJ43M4n3DJZkOiUSe1FWMnQMFGch8D2+ijveYd
cgp+vFwoLjizYum2fBGF1bd6563TzzZhVBkwDXJOSP8leSiF1o91YD1Dc9RidECN
iVudX3o9VM2qSGdxKZB6VQ==
`protect END_PROTECTED
