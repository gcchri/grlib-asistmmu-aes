`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vxaOthkzaERcYCK65wIb2FPt+ktc+HDwH5wyNpbh/cl5E/qu4ub62dSh5Oad3ka8
HiOe+k9udqEnBy4i7SX3ZiMFK5uxzjZz7flRJQAcyL/accBem2Afgqy0hkktIbYK
mmfy8A9EFzEtUOpMIhnLSzAFty5tzJgZJu2v3lyc6HIbTtd+G/8dzX2f4ilMxYX1
TDNkFqrQ1656k1WcfuJNWkKaHTkb4Arq/UdIUTjNSEjKGUHlD80zokyo6o8PwDJ+
gQf91V4bDN1DKf123KG/uK4uWeZXdBWuKc98qZzzq0jnQJCmVt83LDl5AZB6xc2a
spLaFYapC6YSd+1UnFBxC9Hccqnh/03uf37B5o/B4LAoi4ZkDMwm7d2dOsOlHjy8
6qkhYUZItIdT9KEDDm8VVlOi6s+v+fUBqSKemT9QbvHjja7/LJIlFcxjk3KOcPAf
L2FD/QAE/mpyp1TC1ZWXf2KAJ0I37p1aCP+8hKUX9R1EhgzFwBGMpp55uXSBie80
OIZpHPgy15Qc+lhWxbheNMhIle7B8zFrLIzfJhxia+csNja1m4bAMtsvP/RG2ph7
WL86XXcLL95jlFFb9tniJL9vpoQtr1MjQnR0++cy8q0JfHNkn/7+bMvoC9eEeTH6
dS47ZxbB6s8RsK1IfQSe289cEed9tRbCLKB5gvDcRZWL+NibFfw5G1SHQ5xKi10S
k1ySBij4ln0paNsq/+kD6gcwvGfpoGL0Komk+IjuUgoWduVcGb3WFLlzUTJmXg58
A58qdd5yUjUGWCZACfblZuNMfvtHU2caqE/l3+e98XduPnwR8VmrR4SPi0wJjE0m
nHZYP+dQotQWEZW62UaRgXEkvREuTl2snlDJCcjRTPPHu0l9yi66Y8rVgD2glez9
XNvzQuvwJuUAn3tUGU9HBXwDFlMOgeuiebqO/VkiIoWj87eSqZTGTKNKurrJnFK8
4e2i4MdCMGQ3S+Rb5aMy1BYz7ol0aNEhsrPmUfTaif1IDvaW/6dO/WeNHxx9fjBV
prBBnP2Q36bsNR8Fv4dGqXuBHSzBKJmtb6mQCl/GM/tQcfdT1UtfntwtlwCoSgL+
lct+oubm3h52DMg6j/tWwndn5rUjuzIMAuK0X52lnrkIaGxnemCKV9AcwMmuk0Yk
uJlW3uWwXC/rfz1HQh30WsaVm4b1o0WIzkr2L3nVJHq/oB6BLP+ilggeisEH58AZ
dW6F02q8RViARVke4FYFSdQbCgqz/agCAQI6v5SwtER8M0VFeLrfay5qmw8B4pUY
GAPrpjP3KsKgV5vYTH+4LOsPvRchG4WhclXk9cBfBoIH3jXKEvB6OSFsaLtDpLiV
IomfwCFZ9TrYSCk2nLvQHQgh7UhmpwC91tK8aFXL2CZQzQhn82MCla2stzrhNMNm
hJTACQuvr2O5k2zoxkBXXqvNiCftxJ13/CfDXMLZ+ssoeWmyLm1dq6K781Rjgb0p
Tlp9jLGoLsO2Y2UN19oLVovr7n2ijHCzTF4I2vTFzeKHmife3m//keOkeFY35TRL
ilH4oYprEO5BXVaLpXGz1DRQINHtcmZ7Oe8rsognx2tpca41IhNR0VEg89BbPc4v
yO9hXFuUXsT5kS7XS3RyXEFk79DM0WuPkFSzYVuGAqLfN2el/rKEL4pRbSnCTYG5
9aUY6RaQbaWADVJmaiNLWAfAALiuF7llWiqHByPrpznFTRThUquDJaw5jHXVTSqa
E5SGjX7KPObVoL6920A2RMt4HOYuO4fYGTSQqOBP3NuiXNzLoufSjrHuvoexK7HE
W/832/jzcq00dnBeD9enT4LQ9qy5/VVXsFX4/LG45GIoddpIAdOmZSj37JrJgiiZ
hqqDQZMfSsl3h2XY/7rPLROX8Ba3SIPyGWQLToZX32V5Qzw+rPx86KH9NFp7cg/u
Ed/VrPpfM2py/48Pz2YPRzwGkEfnpb3kTKYUDVmJDJEViqcWRk1pe9NtrtHgNoX5
5L9aTJuQjvt/UdyDpAJNhlZ/85S5jvWBF9w29uZcJXIwiNu0gkUB8+IiU6sr0kqX
xmfyvS3kZk04q4bYhc/pFG7+7XOSHClilJtw1dby/k0wBF977T5bf8Z+pp2qQiJX
4eNranUmcnm0JYCd7h7MyYRHioXq0YNiJ9XUglkyf/Dhr9x+a/HMdVnV00EjwUI+
4NqkzIpiX+KGfTqGN3Sbe8lWV3Q9eaFXKSnbDM31k5hYqKQLCettgCO6s6hf5YhV
q3ZS1ay79IfcPMns1dft0TrXLgz/EEubOl7Z9RF/0u0m3klblQRsFZQWu4MEenVh
kcwlrqYpI+JYWXGgU4R2ynzLJfgy8Yg7nt/jzOdmFcDiBi2k04fuSYHA2V2ny0ap
/0y4cCsFZrRaMncacBNCNb/VCJF5S6KVaggVirpSsbNiaM0JxdSbMrby7K6+g+k9
MzGWXvpt9X6XSWGq1goov/+GDOD7g40OyI3xiO9W+7vJBG/oDzuzpsl55iEHZ2h9
EqMfrK6/Hkjil5ciB97yEUlT1GhneJ13sbWfXiY2MomDrULKl5DB1pmjRHbtQAUx
9WdQLXeve9AKUYu+ew+WRXzUSXpw/EFX6XVW0qZJfaVg0N7cMs5aPBQfMj1lVE7U
MO0Awh4hE0/5iz1MpG4pkJMHEjPrsIpG7zxvmMWXzjGWYr6ApCsy5+LHhpiZ7P0P
df+RSI09jNxEKD9YrKk+utCXcQuNdwHWxVfS6DPvxDGZjcu7pad3XaCIRXDtD3Ch
0IhbJ04OWD4mklWBLitZQuwa6UHoACsRTGqXYLk/7+OyWPTQO1vKlat4iN/Q7Wr8
j/do1U0STsgEEnzxinay5/gxdieDUljR8RFQ/eiU1ro5lnJGwM1YxNsp3rTns5Xs
KhJtTYyUn+D/mviKQy8cd1CW3y1faBzOyYucblDrz4Je2usxIIJtjuIgrtiyjcDk
+9/c/ga75mj03idWx8ElqorKcK+/Gy4404AJx0M//OkUto5b/nm9d/gNJVRng1Zj
dhm/0SLJSDkr4BQIxR59LwUnq00JLGlI05fCKLgeOWBfcOs+fe5jv1qRrEHmXoGo
1nLGTLW10kYRjGsrbkeS69IsURI++5Z4lA7kjZWydh7J4mmtu6J3ZBTHcktaM6C3
zjQThBSYcm4HTbZo1V6FwAvD4+1BFZlH0cqiSWMILXLnGznaPccddKvFGuCcOjJd
JlOddJAqPKhJhepuMZIx8q+gnNEei2W6Nxyq3wYI8Z8zKLVu5tLV0fP9gmPFfixG
+m+ChOlpqmlD/AB4Vc16IrIegujIZPOfXuMwmsUaas8eI8zd2Z5qYcOBFX2hDnbg
QNDGmhNNn0lKX4AmdbPibFqiJplyM9g//SuWa22WfEvW3Nhs4heNlpf9kXXNOLXl
1kH6Cz/CkpEaEs9Zf4Jqe+Y2ZGMntMLhnurSuf+ONp7gr9ZyleUA71bZ3iZEjr1r
rDt9jfH/YFzfdqsIqLiKffcVju1aU7CLgeVBvyydhp7svOzUpUqLRqnIeKVhxuEW
HGXHhBOeERW2dMuMb3YoDK0LoKUZMKlSbiiTyZ8mPz+Mgr0S+Io07jTkhDLr9ZnC
uXhoMpMEWWhwTIIbbaWlNme+sPifNGfzPX2JbItuCtdepl3LppgnMQcPbOAQhUza
9WyZqVxYxaqc26BOAXyHrHVm+xcQGK+aRyyl8NoKk5KmD5LDiyhvi68BjvUF0SAo
2r64naRtpElOzuQ0BwpJOdtx7IvkoxD/vUFjRRhQ0FzNNnA1otgL0f29e+KenJu2
FNL7X6H7mEQ4C8OmGEy+5l0VXkOmoyUqT5eYi34WDaCECgKnl7sskmwJ3ppvwOwx
l9MVjL2C1kiUXNgucb++MDzALZ+us5KHFh+So9MlazCrk14WJEKEFGgiYUTftfHB
51xskOZWSD1U1AYYYwYoxydLMgquYqOLGOqiJVK3XV803S1mY994I0GwtfTNG4oZ
+xfnXYpimfFF10By0YOjOw2pFDmpVNMGkxf9st62f3tHe2VU2Vw1BavxNR0WYNcR
J8lp6a8JqFbIBp36CHgi686Mc6xO1cmrdwxcLqOTV66iwnKdRBV+fTr+La+fm0V4
1BTL3wZr8R9beDJIs0SsD2ZQ+E4RcEZGktaBYkAoQAO/AJ29bc3qjKXtcP19qjtl
9/bigYR8ym3MFCRVoJC7EpN9jixK+5olP1mna0tNim7NYQuPIEhgi3yHm/DfRX+D
T5SSccKTphgoH11wdhiDjlnJGC0D8Xl3H5lVv7uBsOxVKdhM/8k5PwLVBOfUrkMf
lxYc6BGccMHmvBLBEMyz5nLXejhG7tE6CJdGAp0fzPegApAEwU6mkUoNOmFWcrTe
yRs4O+8nwV+hpvDkiUP8zyKNxA/0YpDUH6KOYron26giE01Z1ilBIIG/vZoTO2dD
edld080oSauPIHWBMK18UotxbPVNweC1I6S7NEUorkwD7jLN6uEIfjAgY+QYdAc9
ROxNOvgra0sWudGKp+B2ueOtJNa2ZlrlFVoopNlS6a9d0rSAK1u3XSRcjrt2bjs5
1QOFT8DD5O7ow9pqOVhP55//oBQOgZqVHIJCBUGhLfY32cNugDx9j4qyzqLNwjjC
+MFIPJEXPvsm/S0lyu8Czciyfrbv7XkbDF1YQtxN7AuTkyULMGeDBdxlKfTD7HLM
634WdPPpWuag/TfN4f1QqCGqm7k8FWj58AAYvWoGsBOVAGwONSba7eUBd223GIzn
ZSs5ux/lbq0pPnoedL0rJpW6d9goCCht+UfjE7KCIgwbjph6v0lIvKQ+oCnJFWR9
0ak0yqSHY1xXrl3c9MJvb9+aL/kjwXIX3ZILqCOyLbBmRQt1BbZWi+ZWrj+ZJFGP
JrUdK5ompTGkEgk+9+je8Y/BrQF3CI8Dj04bV5Cx4iqYKyP0+cs8n90TTQ/yXhqU
kSlKxzvJDN1QyRomRX1xA+WIafsnPM0al045EWNOaRLjpNwG+XA7dyC2ps16ADDj
WzA7+eNmL2AN/E5IRd077MMr1S2PNmSmyErozkzinmhfWDEpqniaVXXrG3b75Xje
6NPA1YKqKyCAqLVAUvnSNqV/NEsQoqoUXiXgRSJayYF2sWtEy7xHh4EUqxMAyA+r
sX68gsIbAVorKGF1a6LeknRrK7wQiLcPhkGbP9UWpsqURY5QgTD3lrrVGWdR46lt
Mtw8n5boBgkP0mM4zLhWxokzRgbWNckJRc7Cgj0lt7VSYWRusq3Dl6mXUmXaWb5j
CV2RqGFl4IeMqHYFz8wsSqNpQ0bClaAf2zfvVfaAPGlDN3dGhAc/J4CxszHGz33p
Ch6mKJlxFaEugrLoyp87VuX27xAZGrQhCDS1WOlYp8JuP+7sOI6ecDTtzdDlfOCR
fEJ3msyTYu/4LR0dyfTe6FPH5Y5AiRx4M5RzZJ77N2c732U3olhd0m+L5G/CYGKw
CArJhxvXsTYA0h2dEkXPaz1KOzbk1kxNBD1Wk3AzVuLhtfl35KSnvn5WeaX5wk80
pYYYut+4Dz9/jtcP40QKD7u4aPIAyyYLcFBBlmgsXwZxRewZZZvRWQLhIkVPZDF+
vN1kkcXO0jBAn7UcKcNoUm88XJ4ehGYkxs7HqJ3EZppC4ojPNl1g734fBHSeyejk
RI5qLpwovN/ntuW4qga/ETzeI4tJ1I2pf8U48AJpmGFIIboRf+bRfIiRUr0d4rQF
lU23ZW8eOhxREoU0Ea7TqHrfxOgrJ6+YxC9UWJEwOLZZ02KNw3BI3lo/GK47UMXO
ZJj0OCb3/MJARW25Wi7SD7CZYlO9C+uELvVRpSJM/1+1NpfX72jAwW9VV/Fq5tSE
qbn+HAu2L/F4FwS+3TadQHUKf+YwXaXBkg8GBuWAoE/flcBL6H3toytHg45+uoSd
wL7pKP0XXbjOFj0fNc8xHS3IznwMV+2tHu6mhKqgwilN2geGnXgq0XcA44Dfc9Dd
3RCh549GTkIcjMoIpi2decaZQJ3ES4XVVYVTSIL0iUSv5iNN0Y7wf0O9HvaRuv57
y91DfWZtITGomzsupjTtJMGcEC4uUp5rWvsjldtxY4hzo88rr4nDRwAJwa5Y6Cz+
YmvhWSr1A/n0kSWfl0VWQy9VuvHKTNZb3JkyufjNxfaEW9b4ios7dOA3/80EehUJ
Vuql6+FEzSvAQrPkCyV5RrVH5HRnEZmv9CPl0hh5hktCPTFREexgeClJf4gKDY0i
cSy5+Onck2GPmOBHUUL8A0VEm0jhu3YajJoM08TA+MCjfVX7u7P6nqodr5KgGbH5
0X0beDOTCqM3wudJS/+nUMokINaOoCaKeDaikJTwmXmQYyl1oMj5pNSKS6i1Dogi
Z7BGafxqK88Ywg0ze+I7R3fXkIbaXzghcei+5ed/ls4kxHrsG3iRbA6dGlZ9ORBo
o16nXHct6ftepDTOr4q0u6oA960hrlhs61ZywoUJVrkiQSGssxhMnzYObmrUDmdI
OnGdMsyLNCAlZw2W/EYGsMklYRO6NqEvSVH8Cu5XPIXiOiwhoD8YlbBna81dqLcR
W2/cPqWqv2E63hY+DcJkKdyb2nPojm4Jxw+AOcczITLsgVyCSunO8HgWdENVbfKJ
tESBLx6A82A6qJalghKHWobUU4k+zjxdrKvm66RUBww=
`protect END_PROTECTED
