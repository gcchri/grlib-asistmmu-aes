`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QEvNWEPfbhEdCWUW9VSraujgwX49greZKzI9bXUdtbNo6t60pyMQ+sKjkVACgo71
i4RngUduaquyUX82N3HR7g1cSglQWIK3aFzkYaK11d8PYVe1FWKwCi+L/jiiA0ow
u3k+0eNMmwOhgroz2tvuUjHyRU2St79zHJuLh/3eQ6dU0ggGHmGmXyEo3KnNuqqC
o/g/JoDjAwGr8+aeuRrQsNALeyZGB51AZhBySxLzL9Is3XraVqC02BDHaBeUrZxq
qnVJILz1FIssAGzdjcmRLCLrd5SoFTdbEUn4xqkzM1GESpiw4R3zTAMV+5seqfJk
2lK9TaYFl+6ubuyFzYt5RFOPRndZnuXRz6nC7kLFEOkzl+v4dtFF88O4jXHlUQQn
nutYNREKFsHD7e3JCfs/KMeuZwRudIZx1xRqp8QqR4m52jS+FDiyrEJ7zPZRkibi
qR8Xlidfm4guL0DdOvrz6bLUabbPEfQxQBW7LWPkTBYugAzuF1ZgeGkbkYTAqRcl
78JtuZrxzVKDx5xK/yhsph/Upr+nmPsG7G/wzFrm+3EZQ1/OMG55s9clgM8/VD8g
oySDg83yu+BYqql+3rS0MpMowQR7celq5GpoV8JMe5cntXoHFxUuiqpAr/cWd7W4
+Ph3e9TAVmx2PO8scSpPR/DFZlwloxGEiDDsrUpso53i59jJN4IgHGxKTdS9KFek
sQrAdftK7V6pm6x9Muvs7E7/5ZEU8LFaBucME2Rt9Cprfo7/PsLKKHn0fXZhhSoK
qMa5UUJ/KD2FlNx7uyLj5Kiud8VhbVyTOlX610noTRQs881I2vLEi6BA6uRPL2Nv
2odkZ2oQ4vkIWDJRpoYsriTZdOv+0bi6cuvs8eQW3ZUR6KVk4O83yhyrRnzPhKQZ
eU+PYGYqznoSzngJUI8aYSQrGj+igfrgMdTNyzQkqzwqWoEPeyvco7xGv5MGb3Br
u3S7SnIsJLW2smqMBhttcOxtMjYiz0XEjCwMgZrXXfXnC6NyPZrN8ihqgz3J3mbE
cvOnysxP1Gk7vJYc1WJYFWx6UwdjjBDghJDpbsl2A6G5Ak5SSGMpVm/A0noKlvJ/
Xmw4c+wqwZQa5lXg7RvPbNCNzUJ/EuX82xqdXAkLfPHp5v1ljRQMvQQbRph/M3Gb
+2o5k6OBABvC61vW0jItdXmyzlGgBKf55clhhDamyGi60f5tEBiAS8U9OO9xdXFg
J/K8LsP6WGZ0TGP9SXVIIlb/D+XWriNUUhRYLT2N/L3skL13Iv0zs4TDZHjeoA2n
WfjiSJbtOm4AuwHhg2cEcjg6wwTFOgskNBWXIh6jxEnIHI/8FwhECo/+6sOKyo80
im181NTukQyA6o+30mNaBdSmMQVOyZRJSdCjf44IXa7Fo1ZYczSYfqoJBkAk8B9v
3UH6RlhkbQblB6xDkLodNefKqddosqo6iWU5rVe4UKcIlEZrP742I7yD+PhLxmoj
F2oHbvvKxY+VauusvSaMoecj49+QesaeliIAtYT16vYh3gEFgY68yp3o82Ua6EMw
hJCyPLJDlKLk42ywWIa/6CEV0KIIvuoMHj/SzXorw9chCSQ+udmE574nn3KrfPP/
y0ZvueBhGjcHI196VrKnbvRzVsoH7Iv8zM1jqlSlml859NHNUy6/2Qhsi67jTYep
dK6V7v/Ff7nrKJj2MrHb++JcdM2f4MJ8x9jxBDhb7GV1vQP9GPix1YpBRsnOkrby
XLIFqIRn2Ck3SRiFR0iblhfH8wOJeNM9+AKIKRXSeKqHTf3yPWtzhyQQ0DrCI29d
veoiGIMApwl10B33t3qxDAncKhdrbjb9ktyaJiP+KAatyFZtDuZ2kdAKvmxRJe7V
pabM0jjhrjzq6hNEgxG7hxTxU0J2xN/9D0LpNwzLKs7qNccyXPsG1dN74P5tVAwQ
z5EkpNGQZxrpIg0MWSpyQP99+A3MOeziJGPMTvWrL+fwQ4rvD5sHXsGttrlNTec/
MW09SmUiRYDo+6zwTRDu82kJDtBqPvUxXmJAX4qZ4uT1DkksPvcbcHbazDoEQpQL
Hm4cKPmA9kX7LLMfWSp4CTJywnqa3dVBIbkGVE7rIsSlXFaQG063sMG30H2D+Ght
Jzy6N3mr0ctVKQ5i6vrRDOXEjGGSYUg42LffC8TWy3ZSnmJCAk5S7KRTMPg3GqWD
bqIZg34HlrwKQzamt35pgo1jq44gZuKDELkAz/DiguTLwXP2ubVqJ1YeCCkItN+4
/T2qm6RPeS2E16egqYyoHhxCntA303JqnloWi5uqUCdajLTp14duvznNds6oB5N7
HMR3txjmeE3VuXNtqpF+e6Dq8U5ADD2FR+plPOIoVsmLN0+k6Qc9Pd1wQgLZWfIz
smPrFiG42sFLGVyFdSmmsA==
`protect END_PROTECTED
