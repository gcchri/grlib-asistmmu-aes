`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sHUtz0lTh2bk5CzAjqfx2n0aCkQ/WRo8h3B3ZOweKt+y4K2UhwExUYNelzBEKhGS
C2r3+fp5mlo62NPMcfYIyVOE4LB4WofqHBaBh1b7xYkiSVU+JDZ+OVSzE8nMpCzU
3x598KtEYP5vkwZ1bo+kOIPKMBVDXG0MGKQddyb/EK2fiDrSCaK2SVFhlfEs4ZfK
m9Lbj022jYgE/p8c9C/rGPg/+RV3AYj2CvLh7DN90AHAFIBED0R/ts6OWAX5uBx3
7Uk9c5t7Iwr/KAeV36SaGfzACv2MxtOJpZZcxNWgkY+U3Y69kTlY9sUnf0E2CKj3
4VGT5IKHo2yO5S/fHZ7CJrVKU7jzflsCPPlezBnAfkOqPJ68CGuNFT1WW5Rr6uV7
xwh9HyoIpDjziXEkJBvV6l3+UfbbKumWf6m/b2q/gunnrPcPM+Sa4kKhnibeDxB7
Xp/2HCeaqtk8iZzZ7mKvxmFhwrslqUx8VtH+qaXzIyNjyi1dcaDk+5OOtNJ2lB/H
VgEGJihNGkzV1K7XIueizN32PlRitfMNP58yA59L+xZCmccA4nfMBXpx4aIys99V
Hn+r8vpP25PK/Liyr9JOabbHfk9HoAhorCZI19bNJ/eigxY0fdKzGZdQDNAbZSmb
boQurLcLXtnnmJ57SPl14MjVKp+anJ5V/9j2k9naC7VM0OHzTQ21aT+8Dx+UL831
x8w3OY+TloiglC/oRywLDyYP7w6t7/qKkRjAgImEk0AfHyx7eyg4H+SPa1S0n0wA
gTzZlTEakBl64cEEuH5bOdpJYBKGIeIwTS/hsqoxC3iSrb+fGQLKhoA6i5k6eId6
N6dphUNYeitJShrVVupZt1/K8YLtgTHlrRLn9ZVHy+zTtN8lWDwqp2A5rMvcZAg1
HDiu4WSFJzdEyH7dHt//my9CjgdhFDqP/6x3UUFh1IjXIzm9l/CnkJAIh3D8Yuls
yxpNe3AtIZ7Syk3KaLpwiW2QfJvCsGsh6nRwohX+hec6dp7t0e/SO3C5r6+1oErk
HzplCw9HDy5R4SpDMN8Q3NgGEdh4arhOjHWBIbIwfDpOv/QuFwZKpzSaaVidKpsG
szUxIKJoToNj2VIUxotFC3kKZaGgxaE2BFCVUNtZbmv42Gm1+T71CIvm7Tyt/lh8
90kIWsHDJ4qz/dEuDnWLqYsMnhGR1WU8/hAb5qPLgfqnXrrFNbQrQcj7ol6zAuNf
TOR1N1+q+rxIposRFSCqHEy28WXzRTGBxCGOCAF+5fqrjGdMSuKezsQlFtBRr/Fw
fP+izYavjuYbsKCchKQA7DwHjbnINLZHuZihA6+TPGPKU2V9WTcFcgyx14tOuq29
g3NChHV9DvwmCH2PY/+SbouF2MpYvtiWGQ7CBW8MmM71ty37WArRXkSwo/kjlBBa
dFzbcgtaCR4cO3LQcnxm4e/5t0vBtrVtC6Ogdf/MOBYhXwEY9RAmfVAk2qeRk++q
bYbL8dD4XoTToYQ5sfaq0BHa8SlE6z5On4B5ET/cdXqdhf5zJeB4YiiFxmxPoTto
RFs4wnUsm6fvAYW4Zn2kIDMcBPuO2XJ85+RkKe2T+yjWrMPMrgf3ivmxEzzCpZsX
uO8QfnFlQ5Y3/47AMDzrNdz/ArlhBF2QU/YdkzbW7I9xZVaqAgzpHwbOqoM8bZ7m
IXzhfL2B5lH7cxx6pNlFzgk5hHOQTLBbVQwzvPI16uauQY1CaUTQ3YKndclSD4yW
Q7r+br0iDYYK8LsjDuSPf/VntZE0NseKIQG4aO4WggRaVePclftEVFT2KFFLCM46
RJe5shFNIIkDp494MzlPXJknqKamC06TaYb9QQ4e3jmKvVfhxHnDk9umqr5dYByo
0j71yE/fUAKEblyOncTg4oDzbVK/t7XW5HfeGtgL+QW1pjs5KD055zFRWlyJuo3U
ZoMW0dVx76ld27MK0Q0vB3WY/Zb1iUm3r4IwRETCXUlNoaVpp7b9EoHV3BkMpC8B
W1oKCmu31xnWcFY/XXUevp65QhET0loOXmGlP4NTlWXgwsiEGX9omKeNEeYBukym
OxTbUtncl0oKq2hyc1g4blCsOb5VxZZeSthS9IrklLqD2iffo8i5wBDMeLfcFYO2
nFRaOWyExm1jtTOhxpLXMs1LWcDP3x4NUsRyNYhOVQ45/xskk+qT6Af41pa+IKL5
3S/9uVgNPuBNCdtjO2Ixn9uE2jqEcQFjbfU39pwSW5so0AhZQSvnUCmC7NlOYcwJ
xVpkdpxH4TTnD09WzrE6nR7UXhDvZB7M9vocNFT4ZSJ+4SCvP1Riskj3maMLd2z9
IiV1vk9/BdzJdHE/zsu7SsM0mNX9G6synEpH0kerCHRUPSoHuhm3M5IcQRQDa8xL
If1dztfE/LX2SLtXTNvEFEFu5qx0axKSzaEbOTNn9LpMrXcZr3PwFzvNHgNuU4Xk
IzNXpxQihGVtc0odRmGfeJYFu7YipcRaaUzu5y24mswOO/K5aBoauDL392NE7Ict
YgH3qqUaYkvROt1yEJ23CBzPcyPtOCBSDxfD21TtgHP3jVMqBp9eW4n2chhqW2lG
8LPTKJz+/TXXV1qAjfvD8BWlVP9/ZQSPBR9KH49FDDta7GrcnLj/GKIPPoAmRTWw
RDQPf77uwO/zWB5q+yJv0L0N6uKIDVvLji9Lfa08ICr9O6rNVFJVEVKuTkACJCHz
ADNl6FkpjQOz8oS360ruuZAF2FF6eNBnepoB0KSGCAfUbyaex3vSsw98WjxtpmDe
fEFTyZv4/K/UBhwkcZmEjsuqv0Dt+qjZGQtGGOlFYWLPMYB8vcwriEea3Jbm4cRO
ZPxV8SA4Q07mF0HkevGJEYphKmqPryCwoR8VmWy16LC5c1kRfEysJd9D/E4JvDj8
1IdFWTSJGY8UY7VZ0cAXZj1H5Z1oM1mmhPW/kRcr76yCMSm/JHVlgrQjCtDh1fIs
/PLhnAIJ++uwcVF8r/d6r9bbDblUT5Wx9HgBsyOyAxrymSou+i2OkBfliFLk/55L
ngjd11z+dtmz06TITjmM90cMem52I4XRPJxTswi1GmeTAOitJYkd4OAqF7CBHMem
MSJloLSCC71Fsa8itcYK6dRsVLaXfj3LAEKC6niXu9/TcHgnyEonAYgYPJmfyTaK
UKEqYKaVb3JVee2GMkxsNBZBeZA2S5kIhAeVwwpau/8Us10E7DyNI1VRT3pa59YU
UBJkQ8HtCDD25juq7rKD2WwDNrcO60lO2yfdqCzt9cDy9YHt1hT/0dxam4aRNEwC
pN6qJgrC2PHqxy8pF1ozYAcH/wuF3ZKJ20jghunTmocksU6cqgkjgHUtFuH06e2A
Xa/9T4pt4InZtVyWtRemJkVImbohGdNPCagS5O2cVpPSJ/IGsLQGm5a4Gzk6FPg5
lYvsMObCdtguVev8y9Kxpa7QYV/d0n97GxKoPhQfN5vg3AbIQhpPOoZhNeL737+G
m9Y6mefG3XtbVqqgKwu5sycTTU74cCq9zHOUrvHovqeXgbx6WrJsGHk7pqYh+hmc
GamFz4CdFigRjLR1+Ji4VPh+mEKYBQcwHzdp1Ubs4ed+QZ814gy0pFylkjHgp6+j
7Rjfq03IUcDJTrC0fSQMZsyt9hvASzCx7qFx0pLc9N7Nh66Sab7CYo1BDQggoRim
QLQLxl6knWh/IMfwbdgM9rnmWFwO/VkXDdc/0c76Kf9PlSRXU0U92sYXCD5GfY+B
5U2VsZNzqZQETmRS4fFnGRmB8p/J/lKsT/YS1Iinpl/VGMqqCquq//tgoqrXsSna
kLYJuE59O/NDpFhbaT6/R318pr6AusFOyOHXMwVL70C1oGfyLxtd4VO8bOnyeCHo
owa0RlBtXsHoJC3gUqOtP3lda9BKv6yFdQh6gkv+PAmmkKwaYpwSjt6pIVuabNuA
1fRKfN5ggw6zzq+hmX32m7zpxwIHd/I9XN8wlqEPCrXgCfFqlaz/t25XvfEDiROn
EqoK+6Ga1qGh+o3OFeYh5bEXRiqmPxeICcLjkMYDYddDk8yf6Z3ERtsigZ3unI/C
4SADct7T5lsnSZnH4jBnw3ITYQYol1v3UVkyUhCvJDD9OKHRL79uf94VLqahlZKY
WiDwFuju0hLeHhqpwEihWmXf7pEVMJDJgcw0zWLtvuK1i1gB90WGlnRPGgZzcL0I
jp1VlyteLSPdiueOIZ3m0vVDst183NPtBofcdaaapOgJ4l6sQ6cc6pqtxtY0So+Y
Ay0wDH9qMiHi+kzpRdWC5iFGqmR3sEN9ryAY62PVxDilTLQi17+ZYfVmLBqoNNMH
hSbh8VNFeG1ga9agGI3kizevvLeT7phC7wGmpOk1EEGnl5B12QQg5+SqKN4vBhLR
rUVFWkeHxV679Iuw1LQ7wKGXXMR5fi08kcQFooSnV6wJo6qcqiqUbfUlXMVnF20g
4pC2rhcqgO98rDkBb0GJDLrSVAJPVN1mumG4i5sFHrzx0UjHYDJYEFCC1ZxKjGj0
ZFtnwX7zdNCDhKocak8I7I3CnjNPuDx4hveqtrCaLHkRZ+Dg7/EIxkCkjK9DFjsb
27S1G0pTnSXg0BXiBwSVBLUM9mGP3lSYrEcqskB6kF1MK7kCaK37JuAs/94wCrhc
FqoWsa0zdm/PYlpkRMMe+yiwyWZkbAH7h3S0MwvkGRkMRW27wIh6Dyz68fcHlMSg
WolQ+2TrOQ7W4KnaGpP8uZ3zGPRZGHK8YWndzK2dgly1vWMv1TBewvlK+t7M9Bi7
7J1uepIpcVjsfgtIKeRXPy+3MlczWLm8t1NUBpqeU2baRy0LPluxTPcgpOAv0BXp
PSwGBhSjkqW5jtwoSNB10onuvgwo3GObFRp/fwYqgFA7rr3XS9AVZnWmAMW0LZPI
H8sANqfhLjDUaYuZRDtBeXWMb5O8DlTzg/bKrvNtt7LW36bOMwoIz/O78azoUUJK
Zr7nt77TYMMboNxo6G1k/UoJexbmOBS3RVSaKSnc9XYvB4IYjIliGk8p5cGJ1oMl
FiVcD1tGV5n9cigDccDZt7xLdIDJB6rEhToCkZYPrik=
`protect END_PROTECTED
