`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1d+Ykk9sL7masEQoNNNM+RisH+rbvcpHyW4G0n0fVXpifOPkETaB1ry04QXgOfvg
AVhA9TWjAR27nPSPhUKSpSzneykTnuDgCT893xQBs3pTh/ferPAvwpHIcrCV3Mkm
dboc3QXH7Bp9QUKyUg7bwl9mCh7xuDVET6bkKw/Frh5tHIl1DZv+81XDZIB/dte3
WETUndM915ecFd1TyICAS5IKGP6EiWdfldpKLT7OdguyWTREZL4x7EFG1D986jAH
B0IyXaB54FNW1WBwMnk6rn3eQxPhubxut1ncPb4opDkjEnVCqzQjuwTcEwFQ9rTe
fhH/0w8Kv1kuf326FzYMAmlCJAlZHJDDqAZmzPtAvu89LTCGvaOd6jOR3q3vk9BM
xWzi144qETWuT+YOEJyvYqHL4uw2jFrAK52cQplE/xsnKp+rxOXSWBwOGsI7Wl1E
7iZ3D29vRAl1Wa/DXGoLOmtCupgux4qkXmIRPYhL1PhvoEJ9RLuu0FjML157PHeX
3w8hnG5RI5qbpiNSD7MD5EN1KKWocSAQXHOvesXpztGaMU7rkmxdcLahF/8Vl9Eg
36KlAvEvnEbWIJ9rUih2gS/6IWDv3viQFPukqDntM5N1v+hj7RqWMvivjAJanSvs
F3c7NowAuqdbBqbgoFYsJ+8MnskS7+Bt4vc5qyyXm1F8fNXMLUAFgAy9xOXc0QVE
qdb/UOkhdRaQH26IHX0p2fr+1u77Sj1m/oVhiGD4Og+iZ+XtD0rS35rhhbmc86vp
/5AjFLtH1R4Zom5IzyJnWOD4n1vLyVAcIcX6CBUxTWnBw1YgdbFkFr2B5HNdcWnb
Uytjvk6jOhWptoi8LOVIjcjEbiy/nfffEQXhVgjHmck004DAR+DD7CqI5RClaTho
IWrlJY31rF0aqp9gIeX6/1xu9/6HkttjHfEy0Oidyv9h2JySazbo8s1ZYtFedeG6
7ySo2HCEHrSrkJc4kjA7XtUps6O9kuooEfjWfYtKbMxGaunv8bmJqteExjCmHGch
ti+6JpupfbsfF0BUXC0EjQfF/C5iQ3GSXdit8H6+/sdRLGQYvCeqD/ZsJrhgzr9c
GoApw+3ROrBpMPFRWrDTaE46GUkym9aw0++zWTj4VwxItbgb3/Tkbjy89NSwDfGY
F/eG9mf/lInYVlstA/1U5K6zmeOnAySaE8hUsJjg3lyC3HW2tfqDTmT8E+H8hK3p
Av2dvsu+GYGr9bQjlvvQ34lzNMaa+PjkOSAyCCZHZXKvnYb/ssDYRwj74sktn/lG
b40Qgj3kvxIfQrQLjnyAE1wQ2r2eRAlhrYO+QbPf78ogC4m9m1q1xXSele0wYa7W
BTvD9Qj8vQOKgyF2AW673C5ZSm+FUFsVU5c2noeaqwuEGIEN2X7uVvBLN02v1Q3x
ydSEfIEq7rgmOvcfpgvp7ENftqhFrH4QC7HCu5jgPhEGMEtUwoGmjKevPujs7EM8
qItVcrptC78jyOfxivoy3/qsT+wmIOb2qpQoEPqo32h8efZxDCeKbAGAj3/2B0EK
4U+XKeXHHdl7pcHWbXWzlhlfVPy1WolGRh/XHb2Z20tgAAa2g4SCINy3S8G4gvaW
k8HmFZCvruD2HROeo9EOBXH+7XsTE5N8wjebm+O8shuVOHmsIW/TAGC8lamvQeIC
YkH4FInsrQtaG6+VRaLlI/yp72eeuMfa9IphKF5IVGnhdHBL2PIDtI4iGlUciBC9
WFsKm6AaVILCzeK178zNb3TDBLCAwt8AIZYRM0DH0xGJWSFvez6NA85+bRBcQv4p
g6wtVsprqkyOLWLIMRMqgrIZP8vPwI5+b5urlyy7GdSr+VVCOm7Di6o4w4tcWsEk
ylSRTHbBi/ZaDBXuOgGn1zeOMqJhqL/ACGb9UsG/7q61GHcde3q1Iwz5lNsbbMY4
pyBKbITY5I5xZDsPsT9uSx9N8zxVj+JAbupRU5s0WfVq3K7vUVrbm8842mgNxFtZ
hPaVc6TtXqGD1UTUfc0C5Q==
`protect END_PROTECTED
