`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B5b9w3xopbLyFFUSkJO9cK/cc15qHvFRcGFVopzO8akzsizZObc0mOutIplPUHAC
99GI6tihvjxqSJ2YoUerp4N3DqBSgXzhdOssO+mhBChAgHCB7cqdGnVLOC7SD86Y
JEACGnzZyRhAYUFvvclIHyZXyDdmOE+vFZPt5K5xCVREtmB/LhZlTJ9/9DhbtIpA
r0uCom1jqUOfVQVKMwRmkhsblrglwAMn4Bv6yXwGxFGtACWAtGT9vkWaeTPDENEp
lSzYIESb7XYrd+8TJ6Z1ZVtUMEmIwzUv8jx046ZeRaHfAkrKejI8tM70V3WjMpmu
JIhbPGUIpH246f9WTu7d0Ms/oSUIlCTxIUc28Zl1aYmIRzbjw2gALnfrkcGpaIxw
3X6j97iZbIwFCtCXDUvGzzboYekAS4GZfm+jSOLm+CpLIMEn0PW2auh0b5Glv1i6
+InlQ+lA2eTTy+eBnO0qWhRq97Dfj2ntyswDLf/LEPnp+3XHDNAriuHLecalnfkI
Mkm4yajfVPVKT5ZWS7HANoSF60BQjFL1vXK/ccqVFeUThUWRgOvWljL3od1HwTgJ
l94rv+OjyNgQR3CorNPrJiH5t+cJnKSWnC3bibVVlEv6Bzsy7qPBXxe6xNZ78ozA
U9pqkIOHGoe/FQV26i4LL02u8JuIfEE6dWbs5rY/K7r0tMj22cIAMSzyOsRjk11o
rEDhl4shIIB0qVhxdLnjunNAGHekAEmriS1dhy0sI73TwOHLpTEM42uwXAwx1C8L
IDfbluZn8r/Ho5TZ6SFl/A7WZPaS1pxfxvdUPLt7+ftl9eUV01v9UzcYRCaqGyIX
j57V2Eh/M8T7vguUNvSHntQSY488B84u4HBLNNCzgHf8/S27njUwilTbCoEmPMeQ
Qa+zOR8V5dAJOhvid6iQ8elrgJrBWDlQsAHZTp3hN4Ve3xOZk38W6e/NibXKyUVs
ue+3nyA0U6x93mhQq32watlqOIapvuZ28woN5L5F88B1FExZZlO1wj548dEfvdkG
nDDew4sCPPm8YIFUeji9HwGMuY11tni2u3pOAV7iUOn2EsyBZ/sbKcHchF0hjf/r
dCLLuyG8sMjDBqLONisPBdCTzB8GVNVu91wRSg0NR93RF3DzA4ERUUcpjJixpZct
UiEo7m2k/RdFJAuRuiWxkgWiJdO/YZbNJ4rnOt/XRN3aY8aZDj7JypfBUQDI7oSC
mDQS/g9toEFrzAgGwvo/T6pevZaXuETSfEjm4DKjn6yNmCQi9wujFi1NVkvFVEAM
huyirYJnFyy4fu2eyNiAH5+ABmGLyOp8ENEv5bPlG+QY6v0afPjVJ2SRQ9rRj+cb
ekCpxa5azq9oT6hH4ARgXM0hcNcRG843DtG5WmN3JAa/l0Eb0m/Z66D9Q4COSDJe
2WWGHjLzsJxDtWXFlrYi5rK6DQJZENo7IFtOUq/2Rp4EtU/5ES0i/b/yAQueSLoz
D3KztNES8QsbnPkV/ugAupaslSCrpcSbMS/U1J1HwWL2oKY3bo3w+g4785v9pTcC
y5kOw0XsAYAzLDhFPlqK6Tq+oWoTTUPxSRwAjqQK3qLsjdIzLDcP8aFTKRewDxwC
wlRLIfkfeg4pOsREuhPMqFEBsZWFjxCJ1fCooav4Gyy4ssCkeiGPOucsiaXolDvl
VLTlRfLBr8axoIzgR2J1XOfTxJINgm+t5gHidl0fNLwWOPcoV7dmJDxMOd/nqL+m
nZ7/UH1yzS4Zk0rj2crTfxZxvQV8u/5oWjNUGr7K1mxZ4QT1IOmRuWcUDchVvVPg
nxQTYBIbHlI2e5fwEwDSYwqYtKjNBBNy0xIUz/PD+eoPoyjJQCuLh/mTN5lY3d+r
JmiTb1WtLsqGX5BSXUQ6SFTqjziBGVSzLtlpd7i2V3lxQO0QJAZ9oIsQ/RCmla9G
dcZNRBljJSptGj1zmDiQvwaNAObrBw4vtPowXXpG/NnDdqPKno7iT3BiGh1RFYzQ
77ILh6LLZ3nKWh0CsfVOurBdRKDnHahzvmBE/uOIqfQrEjO0mKZVZFrVfMV+Kh9k
Mx846Oo2dD88DXMEF7IvuXhLqFFu5Sl0QEmm6mCMtpIIKnYYWhFGB9KfzQp6qjWh
yHhURCmn5zXGvy/hXVZzQG5YwoTkHcBJkWCuQtRYFSnDvPUrwUmmjELCL0O5Vq0T
PdKh1SH2qwWX84fdtRMIOI/9s5HBugaihV82NBw2g3KjcbJGF/5mppkywohaomLX
nOcF7959+tpcitlxT3JfoofjFelRTyiuVVfOM5gLLZUOG4PSruhySunRyrS+Z6eB
ZnKj70RFC285YupjVy24xY3EO5RS7zy9kn82I2Mpd/MXJPQE4YILkz5wf+cnkMLe
hskGcm71AOakXjn4+znST6w9Eei1m25xSSo2Pdb6uaTOYw9VDjaQ2okCoR7JHPGP
BLGefVRBrIIjMCRLN1+GfuI3CVTEoXP7PCbQs6GSRlMETSDf+fMeh2P8cySYTvsc
4F0cKkZhK3O8xTS2fX9rVVxC5izDffuDETEVEUqUoShhL9fqzsYYPVa+yO8QGcTY
EgnL2kOGkAOjs5Cukjw3Sv6YY6tMYmj4q4tmyMDOwQDoK4R0bKEBL5gx+vkNuE0I
BcT/s6MPf+8CnAaDK5POugWl91jSy8rST1ovGjnKQtwkQjYdnqiwt2VF/RVyMfqP
50XjOaoit1FnVVXLTUolqlMlQFzjk+r2DP2XeK4W6b4EyqCYSELIIzJf/xHtSAFn
tMndw/QLskHlk8p8fLMRtcEGRXdISKnIrbPF2z2AXkdpSMGdqXa1KV7j4QmLvEwk
unCMkh+TYNnNNCLfwJj8odPt1Fzv6qHylDErGfEJ9gakZTT427O6h6rKYZSHy36f
wXkdKo3c+7VUaCpjOJksVw6+eCQugywJGycby2PgcI9O7W+/2HkdYCiVagYMO7Av
5uME9t9gQokugqwZr7WsrDn2kcXG4gLdYxsnIn7MHzZ8c+vrosSmws7njR/t0bt4
IEAOGSoC0q+5taZ3K7UDKFQ0HdAy1759JNddZ8ERDo1l5peNC9xYQQGCks9M32/L
BiDpKXmRDw2/57E0mQYmqxYzn2hRz+yGj6T1R6rosjvDAGPfQxdkx+IG0H2PcYic
Or2Ko7gk1Fk4+2GhKVBKf1qfNbFUR++LJQkqPlGGWzqSoL7FG55Z7c8VwgUS4jG/
9+Kajp/N4Ck1+624afeXSBEI1ZItnn4l+6ul81wIAXykHQUwKEjBwTSuesCZBnI+
acKq1grPxZV33SF0Ihny70zWdppQx1H7edjBq10d7CMG6jRzILpGygzTApqhse0F
pYJFTqRBiTrJ0zwtUZ1Gbv6lVvKn4UGwakEV3+EiOugLOj53NRK7+AUMEKI+Glga
CQCX9lByn+hGz5wxF+Ui+36SUIZIlKzyltjlHMSFUrxbqcBoIcc5auOlHGS7salE
nynSjfJpQBP2p+S0k4YIGejHzXJ8NDArl2KFHMfI2OeUjyizeLd/Fn0c6FeoqFQF
U8El1jGoTl1W+lZoixPECmDmbZgfzZb1Ijl5zfeYwl1pxchjsbqAzJ4+OHijz/n+
Bwj71GsRlHG3m7FwlGeprzraYOx5QSjUzMpOErd6U3JJrY8aIOIPrFJaL+pkd667
riFbztr/FQcTj/8785ch0Sr3GtetzqpKbjNm/K2iibsWHs1ebK8lqJC51NAqaFJ3
jqjGVinKIVl+5/TH1qiy0f2gXwo0G2MBtvFZPfdngVVdjy5iv0sN1Z7CFh+3e3Gv
AnSAPtfOsxY8Q0Lqv9dT99hnlZ/iDptyaqdzmhRV5WjanfDbY3KbEMDyhjBxYQ1d
KuGWlbMGlTq6tBZF4rv+np6A7/6E61j6boiGPXQbRfsw5qEjeikEgj0HHgMS9TF1
EpsMwI/z+3gbjfCR42UIh67TNBV6eGH6UzgGkGLh8LgGHbCyV9Y9HGpKNlRLb6dV
DryJzK9XMWn5BzInjQRVEmcVRDVxAo9k7EjOm2MmtqLoP1NlW8zQ/7I4NIZqXoRq
tcuhg76N4/cpvnoI0fm+5c95+vx8BKpE03VerV15Bxv6h11eez9Gi3hh3DzVZWXf
h+9n6OA/06eGg0WDcHVeMrSowZ6zC3z2DStHt2gfDbNShZLb94eA7SGMbsARF2fS
7xD8Vvb4VD6JEHvlWxMRL8Bck4vV+NmpHz/b1HYLUaW4cEPRE0xCMFwvafrDpO/l
9whLHf5sbfYDaIksT9wyybW7+zl1QPXXOFThP7oFoSIDF6aF+TyeJsbDmkn4W3nx
AAfQYYoX7cmeI5KNJJ0wjYvYGnCRHbRDjAUR/62ubi71EMc+qcAO0uiS02MuHnIv
8Bd9w9IGud4y6obh7YzR2EAGejQh02ixJrVBHnP1ewblFoj2O68YJEfvLpMtfwcH
7GAUnPy22Qa2LgCxAaB1+/tLMAR6OpLtsnhy5A7guBs10RlnM+FPEFPwM12BIheJ
qJket+ul1Ay1YGcn3uEpbPc9K0oBkKqVHgyoNHeFvMlykWkS6qyJE5uiPll8OJ5O
gd57vew0NXAutZl3fCXfeE5xOWawJXUIPgsPdzr25lHuknRCHdWbTL2R2HBj1hW3
OSrKLadGlmN8yshcRsYgrTEeQhgVd1Bl+9ZGOzz6klJKXHqXgTiC+1V/IIt+D4sc
/RkhrnOocoDSOcYhMhoxcZbXxyO9SB4rwVIdOPq0p9xtCMIQqSabv7mfZwUKqJUK
Hxm7/VKbIPcSzfas9M58z6Y5T0B0Ixzbh/VcXQ/LCae/mrNlEM5tiYRunkRbXu67
M4nOuzolhla7EHgsCELj3eAvNJ2mK9JL1OTYT/LRb1xUbASjjpEJ4VjZpBCmYi0j
Zy2H8axLpDrQGB6NpTjTdQg6cyCEM3NJ8aiT+SAp6gVd5e94hTZOZI2C8N+n2YTO
23kkXOlz4aSLaRFZcnB6UDpOXsgurob3lzfeHGpysnIYgLa59q+V83Mbot+gv+B1
HIzEd1cARY/J2Vq+OK3awmqBMpaRe4ENu8YPhvTI1YxQMF4C/CMc8Yx2tZ8lUxcC
O0Xra8nxtZrjhWXMZoD3lZXz8MH0vz/BddDpm3QwG1l+Ie3aLBDD+ZXAW6zuXxWR
H2s/age6GzX/vEgc0qlhqzJbkeUCUb39fdVykkKJvoPse+lrDXxo3VXXNesjk13T
tCx46tNtrnHZFkTI4/b7G+hpP3B56cJitU6LaKsSUsj3d6SSCnc8VJBHJ8gUgeg0
xEiutI/4elv84eFJhG1MJHubJCGqNLN9uFnf94Ooqx+/53uE8RK/DzXELEG52GDQ
XKaFSiv5oc7dO7ecXEtU7bgygiU2rXJxy7Gh0zmwu27EIZZwX9CnmuiM9w/caCez
iEjAKrsfuTywbAgS+vZ4qC91Pv0srYVN95eKiF40qUvcuhwXXU7pEuef8eiqiG3t
z05kdbNQgtVUudjB9ICB3zY/W7f5UxNRw+rWnfIHHQ/a5IJgLRD/4HpxVQvV06Wm
101LiEe8abThR4JErd2OSQUtWvRuvrLlYdn/xgaYoPk0/e8Vz8VLZzM3btUaMSW5
N/2b3NgIn8MAoS+qp++IldB+HnsBPiC1tTI9PEudR9O/sULmP54PoCsAvSZV/3os
txXdgBsGo0meOpwQMvdMlXoFQ3lJqoFXZT7NNblo3qA7W7YLjfpnLAo46Ukp4kK2
blDgamLr+jd5s6d5a/2wecgok2pZ6RoPr6i5/dI2v4twQGjF+wT1aitje9aYpec1
7S1uWweo40q9F6Hk4BKb6HikQ03CaAUWeGtLJbYHppgd98SMMubKCKMR1jeXbswg
prIzrEbhlnWmtRQ0JCndnCBo5rqrOfuO7N2GRW3vq47FtKgZWEUhDldZ4AGebFEU
28TXF06f6QVf6nGSO5uVm2L1RxzXeiz2UuFPFmgYurTyiV9RKigrbvTpwNugHBzP
5e7JfxUCjvR23eptBHvZmpWEqLlxGvkrOd+ZUJHS2c/C9QVcpJJ9EhraqZn31Hw9
gDd+n8MbJfKZ+MtdLc15AW/TkDzwbwy3fqoZaMNutmdxmXgekYfwmP6SdQQ09t2h
yVcBOOTcx9YF8mM9UTmQswZmxrl7iEIiNtbvfL3w50Md3uXBkF7fY2UsaFcautcG
1FSXoD1rDAO9oJ0Z05R+GWAuAeg0Hld/zjzrMoaBH5zpniO/Syt1+T9gGR8/m2pk
gh66RBhoJ5a6OJiiqTUm5rtRaxj602QMF2HnrUThXGEYVeAkSfej/+PZdCSfHYBl
OB910BJlLmHa+75FG7zqTJx3QrCDeBcqlUE9QnTUvKUj0Db/XLTqjFnR5NygTwqF
YriKbZo2Y3X6Yq7GYqCVXHYDOaGzMdfrPTzojrVtIonYMMQRwJMBmAlm4g5/TG0E
LujDmAJSXtb6ID7OKg2jr0nAAvFps6yUWBljOdgFcYt5fUCxPes7gQAvyMMSJ0lF
h/w2jbL1jIEiWIMjIC4yHJ4R1LCYvQa77HZV2Lrqr6J1Q47XUMKyyeBxAWR8whbV
gMqtiOwTkmemANDWlKOo0bsWY0DvZZVkOOobwrfb8dbV2M2Q7r0QFtgIJaa6J0Tl
f87bzQqN5ICaLhW6vmjNBjD5vB+xaBda8oFDlui1nHQ3yn3rSwdhzpQyapv7gpoF
XxDccnjCwqmMYmxHciL/JOhTUI9DlHRZ5KHXT3+XxAs89shmLsUO8h1I5j7lyop0
vZbK/M5DlXl7FOIaJQN/6TR/n2rEy5eGXCtVrx3+/MbTubKXIHdacRMI8gBCFFRF
K9vIFvafpYtI2H8nSXVR7Fd1N7uAh4a8n/myjiMbX8tqqC2eQNE6Sa/edjawaHRJ
DOXUN2ruo9qzaNSpWF0afu21b/lElTCqZe1Kjxiqn59av5Luin/9EBfJhdETQ4yU
p7CA8cUDnLLqYQY2nf3MAHJCXe1askA35FXgy/qpkMu32XQp+wMwPZa60RHYcUCT
6SVSb3oJEn0wvTWUPlX9YgIh2hygqDBM6kAs6DODQQibvoxFdlifLQ1XqFpcdq8c
6u9SC3s3g6nH8JC+uVvicFDNOAtJ2Gqc+EkLHJEKOG8Tos0Pys79LZdfVoWWAvL/
zEsVpDtD47KPaYt6PyUI/HWeUKfwDUtKdTRF+XMQa4F80rfStCxa4rcGm4lsdeau
pQoHjZVbVtwWxm4rHtiOjw6411OHlV8fSQsXGw69f2v91SjBq0Hpg3UXv30lzX4H
4HdOfYWlgqugQDOXplZYXolWdEJonqM6E9FwBwIB4V/IG3tD7dKqx8iAXOGUcf4W
RgLv0Y22FMGTIyfIQSotma3XRpWZzyWiJrkEBeYwaVOd0/P/fXkYGfojQAWdhBjc
zD84pmni4rNef+5ysT0V8yd/5s82xZq+tk+jaKkOqDcsXmsFWQzlGe635vpwOHtV
u6lu6PcUUg2QnEC30Nu5T9yqbo1o1AFO6E5buG5lpuGq3f+OKAM9feHnQ5TsCgm7
GNI9ey2d3gcdJ1wf+yNRENu4ldwDFOh4/e/l9SvBcHe5OkVkveXKUjTt2pxT0uiA
i16m1zEoa5vjrOYp08OG3fYLuNZ+S0bUrXTszmtY7NW4dnaexhhMYZ04A7NhYbJ0
le2r1Ndo3px1XAuvbEPsycelqsydzMSU0UgU9RudFQwdEgMtERjYX9obTBuTjUv9
pL/ReNXiadW07RtPeHJjnVuvwZby8tC6F4PUBl/+Hv/Eg8KhKBTsq0LX/9wXPi3N
CaEwE7AwlVKyoh7eP++B6BkKQVRkXXXXleR5mXnhQXutyTh5vY0vJ7ST56QX96j+
BQZpM/3prEOtIM0u6GXW4ZFJSgRWQe+nuHbDDSObGQjW60B1u8qog8yr1HT6BAkl
YJsG27IPOIkQ0gj2afil8vWzI5+Ujkf/71GgP+r04YzdcWNSybnqIJyzwmMjJPUh
6yzSp4x9OdeGhdTRlRyQoUKpLyQ6GkMdVoS2jToKgAh+t6DN3rknLb8oCEL6ONPw
YMWAUwVCpqmGZDvHskosi0bNEfLeFzOHqdnLAHDJNZVgDDDVteEy5DrdewIq9VXh
q6wtyEf4dqcE2BnRN0gBnZZZRJViWrvRmCmyA+hzpwpQwCJBJc58uTjAGtSpJHYr
zd5OcAh8UWrRplzKTLy78iqSQPd+/YP0tS20o0IF+rK4bEUbqwnGjnDZw7t1JuOY
p1ujB6m3N/7KTTUYNlt/hJyjircf5hqD2HlQ1ZnIpu78Rbn/VO21Gpfczhx6caQa
iemk0SmzWe1SZ0AS6SB4HouOkAyqI0H5kEPmq0+JALOSliJwCc9YEq5XRJUbY0mm
bNIh+gi3BnHDoaXdgR8cAJNjKGQ6/7Fnqdzr9L0j6Wd5G87YZkksdcpBg4Z4TnvW
ytp9Oin3b8HNImLxpO0YCaXjzSKjyiDDI4Ltfya3TkELjXy8DVDg/kfSOqvjirdT
Ig5o+J7bFof4R88+cBS5T0FWkhKYE/b6WQKucyv2+YxAKWurzgHXdeLQ2mOU5QHM
KHm1m/Jt2yomv/cQo+RX7XZZgd3aRYgAlqbSN4jOQF+U8PVNemnTwnL8IymMaloQ
PXGnjQF8azz2QSx1dMvbII1MGHF6LOxSO2X7Ojs+jnUijogH9x2fJ01XJ9Axl2Jq
phA9Pa7qoBYPePSZZyhnscG0z057HauBM2ANaFIYP+ZMVBIn7/dlZzjaTqpspo3+
4Z7wkvBmUwxeCQC3ANcL/qlBNxC0c5wVSdaKUnRoStfuabbg1snzNZa46SY3gSaN
4KQSvqA10ibmZ7PoD9noYch80miEHkc4CQjkh6MzJceg955Qhc6A3Gvucmk3ZJyx
zZ8cqtbwePkMbmLS2wACqa/5AiiYUkwBZ3PSGYtxeo2M25cvlBAlqJuc4vo7XEA4
0ss69TaJL8r01d7yW5i0mhnIRi7Hije2J1m4h9ecwf/vc8xVKkSxGrxquzdsmB8n
3UrUCcxwGpvUqPP9mhMvq7/cBoJ3LSp2P66s7Mv+kAVz6ivKnmMFlWurFjZl4kU5
MpLBIS42/Bjy6xmrqWgE7ktcZoF5SveqLIR/5aV1ALdxr/G8ZIbUPEEsXSaMXfTZ
QW6AsFeKvLrQ3BhaSOqGbU3YruQMOCbR9Qr9uBUZv+iZ7CL+P+c4qt+2kSQnMPoX
WlRHxIF29FjnyquZvbO9KK/bdoRAzhNUqREPO6yTo1H2hVMwnUu2z0aD6GkokqA/
vfLQLx36DyKAAZ65f7IwDVGOfFi5Y6rOoquhoEtODVulTI74lijwBm+Tsn53QE6j
SjJ+W9UcdN/U7CV5sJY3cuOEuOcQMakd54DG5zahoYVpMvAkwKcvNp32v+gqO3PL
3DkB/WDsSeeLYClycJwLr+V6/bVKSqb7dwq+eZfIlo7PY1oI+bzasGcycD8RSfLS
rMShbrUFxYZu5qH3vV3AygLgybPJcTNQNezFkjcB8mCCYbiihn+bgWWqKcdmn94r
6x2NCePBcoHrbqBbCQKCg5rN0CyeeUzddzuJEI2Vd5Vk8WhJa6wEJf89zQgFaZHM
JbKH83JQ8vmSJu8lclX5Iw26C23EY+AHsLrjdltE+J8utL5+x96J/koArXo/DH+j
rj5D8dempnfhOfz/PzafSJatj8qrbL3e5X/3piJzkTRcRkF10dYTseUugypx+w/4
GkJPppf/RIKzfEaDMFFHajLdNY63qor0T/YedgE8XRhmOKtRzRfjYpG5pLpZZs3I
ye0pD1asPVVI2Fjouxc4l2FtgPGzpfTPVuUIpOqQfsD/3z771gr/DPUDNlDXyXQm
FiiCfzYR0/4a1KwNzp/Me+8tzSHv1O5jo1LnptPYc/VxErJmHSbV2xt2LfCJ9nGE
SAnbT+YWUHoUIKbxzMXoV7PsrhKblg7QTRglVD92rEEhCwuaxE3nmiPvsp3JnNfg
XN7rfQ5vW/RYRgpRybdNed6e2Miu9gQs85HbKTuTnGWQRYSBI97Q3IpC5kk/KCg4
Mu2Mf2AXZv/mjdwWkHGuQz29Pez8dBOiBnSivZ+zahAMAwvxOxqiWWeoBuF5xXE1
I9iOZicuHGOTM0ZAAH3Ny79gPjwvT2Tk4zRUOiPikzxZ9PsA033Jnh8oQ+13zWqw
dLePHS+y3V0l5k6uWnw6trBj5epu9Pi0cF4VrBpAc99fp0QJ4SVegLqI1Mix7DOJ
h8pu8wdQshjkv+BCD5OHogJTrbJ6gprRfsvq3nbUFRPVloZHZ3LM1N8VjtOpHSH5
SUlBcCPpGivvMgQjMt1YyKvMl04x6681yG75DTilcbyxGyOsrjZJ9ENRRlwnCwhz
jPbPUOfn/9kqwf5xBug4d5YnSo+kjbFK5Vdd7hbx8iUR+5pjeUFhfUUEbj6M71VX
kv6kLm/fLAEIlieiiAePZqCwROnHeRD1DzTvenas4vB0GX+UTpdbirFqKDvv9IX0
dMAbDja8bpoT5RHX/iCMorjJ44zNYO0YOnL9bEynGpZ+o48HfCYOFspmMxrm0gbT
aN/Q6qWDJxuc2j1qhgGvaGs7MvBLw32XOyKb7mG2uGLxBrPJcIXJBVdUUN4vXqip
vF6CQ4asy5QBDh0s3HvLicBUjXY2POweFjgsaudeNVx2zno1c3p4uM8aE+RBWERM
IgJWG8LE6Qt5Rxnd0cIxw1Ub0nX+51YB6byF1pwrfLwt7mfqQat07OfkhlFDy5x0
vtHJQktYuVTqSwLcOmhCPiwNABJPWAZVP9fczbFHBfdUnD5pKET0b8w2Z6ZR34Xh
nfm/VmIyujh7a4uS3k7ITWYv7tvPGMMrDcTqF2f3aSp2+Ea+T3v4ON4TgqoOfgnj
YTECnqhucc+MOilBmEa5bXjhDujCXETkOGQZ3/ixYqM1PRmyT4YRvnBtOMpCeREi
US1KSrbzyR4fg6twuFxUxtpmc+CUrE4EUvG6s4k6c2Q9wWOnz6OsDgpjprBb4kIB
G/81n6OjSxfH33oSakz/wwcJRpf6RsCCy6eJ1Sg0YFFd06pRTMjH6dXFNAtoXaOb
fyCyv6iqyQCcnWhbr18hCsviAmnGySxT0Lj4lhww86AQ9ud4+sF4Sp0WZrxuQ/Za
dUi7JPSEq+eXwkhhslGoenF/xhcjrnUSJUzpy6lEl9HqeGU8oV0mPKY4iHWkEPMr
kMBZKcTYR2/DRYqufvzh25n8DfQ01P3zSb1e0RKynXZo3E30dq23+10TLuySY4oK
9OdseDZYHyCXldC4wUYlfKxDCzmuuFVipcq7wYKplp8sJsZN2jHTTN+OVsYwTzXY
4V5XcmMq5UDk86Dmmo09Z1wBn6kXjU5CoRLYTurD6r8GJkjufZyAW7y68io4RGSA
XujBM/C/wl5Ch2S3dbAIPrCQSv1tgvQuNvBm/WfaOvu2GHsWj76M2VlHeV5a0w9e
zUNlf6TVnL4hASgfD8Q0f6goLkgZDP4IubMO+3GrngTLBMx6b86iUyiy8IbJqtWF
ChdLANUCBlassLtNy/E70sQGbejGRvt1NY3/XmYvA2EwySkLJl8RyhEOucMRW8rh
w9tYX/x0N7up70AmgsU9EqbggIR2NTS/ZxUG76uWzrDeukKb/uRZpPW0DQdfjSvY
nOjCjBfvYQjipyTHmVHhD5mLdaO0rzkjazSeV3rfJlnuIuy2sjXBPpCbErYFYz2w
gWpY85QaCBnnRZ93zTZ71bmg+8qXNNbv/TcNLBdBvpXH/YnZ+d+/BFyQQvcaORKq
PlMFok44iPQi9GY0rYzOZS414kfe9YQP32DoOv81JTtbicsOhWgiFIPyn7VcWiYI
j9mNw64dflXQe1b2KJeQbjT2xwRRjgOSvXW8oE3jtppVq6bCd+G8cP0sM606U0rX
O2K9fowUJlL8DA2NXN69oCIzM4in5pL1euob/HgczSec0yXhS58X+6XrsCp3iKPr
KQmjTafxW1Ov9T1szS3qFRQ5RDlqmm3unJ3ixW/Amop3p2DR0XqFVfNAkzT39ARl
drvjdgFhTvG9xyBZTsF/zMzcUTZ4YXjuNbiioTuvl1s7Ljm17nwnThusoWXxdbHj
A87SBfyj3jkNasuvi6fn+JPfBu42kWwr+AiU6E/3Jidsha/2F4AdXgVj3q9y2R93
sn9z3DlZOMoi7kO2HcYa/tiS3uaTDocTDvjym9OCBdjVyLhnr4VK5mTK0MMAUsYE
Dj/Sy3k2tOGG4wUdIn7M8ftrFgwp/D68HIf7x97LI1vHIQBrZp3eKG2UBRxSgd8j
I3M+Cq/7q8pyxaAk3vR1x/eVTfII9wwUoOowrlkJw2L7xkx5UWovJ+cVxIjuNaFA
UoTCieG0OICkZX5kemitPprVuXCTVmCV3aAF+1Pq0zXOawezFRmEMQTG27+f+MYF
GRXpwict92GokcefzOKoqWUBjb9GBGovkthhl9l0Dm5bmCoFIIfIFKakyoKejiSM
oLk5FqanTJab7NQKDVSA4V9H85R1PG+0jqqwceAfBVS5lrd7kr5xl6R29AqEEZ9H
cYXTsSVydCg6IMkwvXG+09kIUNR1MvXmrHc9lhcsmhDq1Qh5MUmqpyokp7OTiMJw
07zVmvwi/7kI6Zik6ucw024w/lXUSpb4sL/46i8pjj6P6NiXtPMwnNyKIoojZQVB
P9QmO4y3JjkSSU2zKwVB7WxHtNCMq2/S6lUkI5465xtkdTTWZv/nBKRcnSvx1wZm
S2RmRN2fmnY4HhxdlLn7EOA28IhUp7FJz2httaTiMIfIDc5UR0nScRJiFlHsJZSi
HN9SIJyadBku7EfsR4qTNcE077Z1xS0EXXkfn6u9yafzcFDJyEDcpGl9/1RPOVlv
ytW3TvVUiQLeurx5bazrODYEClOPLsHtACoJsXct+ZFfq+DYw5Mm8IcR8CDrjcuT
BthY5i8LXdqcGeAhg9Au/wKGD2awhiIAgXpwUyk0uYAN812hE3f0MwGSGbCX9iOM
LnUNRVWNQcm0s9kJzXL05T1CWucV+1YzuGCqbldtTapgPZ3WwZ/PIFNCjDrPe6vm
nrbpe6PZEubK7aTt9+zj7DMAyBOOOCEzwLGrwsgxUKzE0Z+qSAUvjrNhZpjqS0iS
iB18Ri4f1ieAnnnIdIKOUynZYp0Pwp7Nkj8A0z01+E7SxwicfhJAasFsjilhQAQ3
DFOeTHn+XEBHgidLphToSFaRYhQofKzWUKU0lWzP9dkUgB1Fn2DHT8Wxk0y1WPf5
I7du1XaC70AF+/KJztJqjdTFVg/pMw2/g4QfXKheHSH8Ydd06gcChfr8EuIFmpFc
8VZiNWSR2/j/IagzIzfLiHWsfaLu6qeB4GpnQsi76m15KvoeQgUxXY1F9raV9ESm
ZzJ15YjrhkmBO480N9pbip3NupPFvF90eZbW1DRZsj0vmlF1mM2eXCd2BNRaS13L
wjaL2P1dOKet+6kk+tATZOBZ3XUMIOhh6Kio+SDcXCxJ46/u7Jzd1D/5iY2+OLZS
KUvCr9Y9GCtG/zoi/1lyUfvPMsbLTe8EnT8OtVbxZlG/2dBcfF1LA5SZBTuDu9jS
sinYg4TTc0/ssLxinZSeOGpopkfvpIoH6Malt5wZCcogpeUT/TbueQzuO0KIKqXI
8hlJUqWa7FcF4HyIIAg6ryyN1Od3yKiJGrBh4ZBoPqVNaJmTWmIHdIm3dlF5isX/
eOvWdCSC7DAXwvD/luCUeJTOZ7fjsSCQNyPs1ySCIXWY5F6MZVofsTJ4cIOQNWCT
U0dOBrStWDLrH8JP8Zrg87lwMTVTm61kD3DkXc/dJGKj4zVZTOx5vdl6XOriQefF
9qhPBM1zGzW9kC1sIBMKiGnmOrClnN/PzksNTbiOeqfq8NgdTJSARKKY0gROQqXt
Ki3GnTHyMStAvhfddXknqsyNWl44wHpkXE/QIVJTisXno0PQKrsaDS/T1Qo7ox9O
1I3pKxUiyXEh/pDlE1qefy6Q47UMh8tZSs5W17+UaxKq7N8uqHPN/w7iHr1SiYXd
kPZNosiWtiizfmKBbTymN60mvv7zdB+C10+SwWxNF/Ws/x6pwLKMFKSVtR61V9P0
jJFr8twDxqQeWO/vHEKYhIPx5hd6D7k3iRjgzvG3xF9jtHKl670A9uHlcuLP4zo1
cZTQM4QTM0K3KbrCkQ/hLwNZqCVs67mCKBlyROZ6Eu/LZqQK9spGpyl6jLvU1Cx/
4nAmMGDcxqaBn3vBHQi4rxyBCJyEvgnFPxJgOOmoK3FQt1e2MC8sARn1I78l//6F
79s+6jloLuC4k7th5YZJxwFPxHiG07E+IssMS2kfmnQg2BTRl3iqbfdU5uquyqEF
Ft1Cn9DuKHXeDzTB1cZ79nkIsF/gIeKLzQ4DXUjioRFD46aBDgV1eZZ55X5eY/9G
T3MZy3aSxOuQ4AkjZXMY8vJXIL3LWlZhNnv4YH2QMD47rrTZ4sAFrtccnPnAWjtX
C1J0/3/QfddsD2lmTUQUIwxCghKmoY0Co+cKbVVaXyKjHgBQe9xyVfOVhYW8JydI
P5m6bvWlq1mL2Qc5pcPwjIp8Cfd7vjSSYRr7QkJNFr8K7vqR2DPcFRI0a8gufDH6
4pG3fZJ6fcf0tZUdhSki5XFOYCoVxvDDaGgTyVJ+Y7m6fdiuo24gvz+Kea8j9Lhm
fQwT87AN/1qcLZDk5T4iebeVkyw7ecIdVx4DH3HDHIypPzHGIwl0pVfldILGdXlS
MXQcqctwPmnHD85bhuWMtfX65eWTvxlZcsgu/pkuiz2hhg1dlKkoS9zPBpol8qOk
grzSL+HlG5b82knJBqcEKzpE/A7ZewA+5zFQRAJIuYUGhvSmfP7g/y97bgJ/v3Wz
ssHR7ydpVPKms9qMdO7dlVQZBFTB0Sm6tVIqvRitXArdn1NZnBmRr9qF+ARa2GlQ
5ec3TLG+QfLVytr7ea4r9CP/Lzlg+IOv9vQpgO4WbCfowbBOtuB91PSpApA+G6PK
HSYLt0oRSCPO96mSlFXfD4xSGY3MzWWg5EOKo28JDCpSe3VH8mMxYWNxLIm+GuNQ
N5QGHJh0u7G8gXN3WIwbti/tzk4QeFkqcy5eEuRiqyq9IOJ1F9Rlt++ueMbHOIcm
sZIXF/to/EaUTXAiT2/+P7lBfof74kF2UE2kQEO5sk5eqcI9dK9jTfldkNA0SH2g
R4a18ndlgjcRHh31mTSmJRqXNMur5NJy8bcFzIkUDmfnEnaBAGrWtTppIEtfmBF7
6GlozomWyjF81vZgMPDYf5tkRGX2ul5r/l9Y8MwuJfBOQRONyW7sHuLl72k3tAME
6swi1Llyza9WmJPIBNm07xAzaBG0XFnOKOy7teLUeVbyAS1H8g0+UuknNjtBWNC1
+hhmtgg2ANmrHJdv1Ercp+dj58IPMnkrB0aJLmzPM1cQq84tVVVOLOJqRwS2gZnR
PHGu1ydAvgSzTN//zUqLG/mrYZttDlMUtbTzQNrILbW3e4Y8DPhWDn0HUY4CnwXc
LD8JsY7KNoM+/d1LBO1wVVJQq+0HnENq1LBrdBTpuR6AK6CM4ynUzK9kDZEXBT7P
TzazqfpwzZGZq9EaLIAGpcK6pb8mIqhTloALhnf9neuJG6b2Ij6MgJ38zC8SEFoq
f0Hs0EoIuDZjI50LuZWjWT4cahwKQBRiUar7/9xA1+s7srgq7TFstE92SgK6SRDh
PG59L7oM2P6HqFh6yTbUNrv1KhO+R06wEZAZoy20R6GGRi1QHzCXXup5NbZTrK2X
3y5p9paJLJhJsUwcCldounx3qKan1wrbJyRwXhEn9Vk4M9Vhfht75vjFD9UgpV9G
KeqKuwUg1Po3EqRm2WLJ2meReD8YknECKkZoEn2XFvZuzgwKNcCfrYKTwGuTh31E
6KCVjFbeLgb6s7BqxmKlEDQm0NpRSUOCxTGIAeIBSMi4F4S2L0kpf9xwOpj4zHaY
VDeKulLrCAMkRJPeHHmgvgqChYLBSPjiMZZYgRsqvuIHRHqbDxt6FgO1ic6jhBTW
WJ8pVDEvywyWFn8q3w6Z3t0/uwJot/OHcV/4RvN8o4PEJvsdQAn6q4W5Qi9GvlT/
xcTsCfCyhTv6YKZNxaACveJv+GmSWHeUANEOKpBlx56ye1Po/xm3GOM7Sj9hvVMW
05MHCg177ZrTCbC7bgMqX1oJqXJ4vnWQsesGPVNzBMA5zNyoBuzlxFr07vGn7wwg
zs28OZkCY24jjPhKyjF/At9Dn7kqRANZsUHHLU7SnxbGE7gwunOKdo3EyAz+0n0w
lYFv1MDIDXNknvaHCOgCCm6DYgdcYKL83YQcqhX+CpS9Ui3pf9Cfecuvh2Gjp60s
bgYse622UtE6uIJtGJoFVq7RLZY2fhERnF7idZfoR/YukNtvwKEq6BRZjrqhgPaw
HXAN+FnyUdJ7FnBHyFu2aCSTChxztIUsoih4aBeL2rE6dFzsRgpiXw/xANrYlVcJ
AGHbxWr8gL1uAxWoTJzHzW6LEflagPHhzR/uY//KokYLD+wkgIl3Hpll74gZS8XD
Vlno9XS5a0osQBTQ9B+mGOtKD3waafkfrE4x5KyH0iE9za3Ex3sgvcj3CgZFgzu/
9T3IYQH73yoPjpGMBp1Z+gukjzhp65yLLJdxtQ3GZUroxe+Q+4YRa3vMWKa1FaWL
zdzaYssehEz3gM/j1V0XODuE3lY23YAjUeQQ7Q2HX1eKDkksg5SKZyo65nyIeiSE
YHKTGpK5bTj3OaLA8ClKdN/MKCVH60b0w2x8+2QbUrqXBZJBwn7ZIbXh+YxCCahI
QM0DHBDJuljZcCShW0Sx0sbmeJ8GDEH/hygsUVnNCFo6SCC4p70dtTC3TcbXqIRS
UbI4/GoRtrp1GJXReyp6HL6Ab1hEqXW+3Psc1ma7jirpvPzbkhmYLj/EKBoCdhTN
3D6c1ONIe1wc5beA+YSEcd1uMpJZPlN5LeReyowDxf54psDCL6i43SfjThMdKMdO
8bgc461F87IRUfksfj2yz/MBjLkJBPUSxMFRhTTNjxaM1gUnsJHOgOLmKAlmQhNr
r9JiRCOfhpGRQJeiG88rravXAe2Y+3N6D8pthwhtboBWPu5znu9dtiNG24gCOjIj
F7DNKuef5c/ztMA3YagDoD3NHNW/MvS6E35Tbjhmn5GNpjYlQey2CgMEWbh/pteR
Yh4u/3NDtnqBtIufprkqw0Ssjqrd6rdF4CxTDaHvlMwdG5dH7MisrhmSWFMcBM0q
dTAtZNJkVaN+C7kVGmn+2EIb7hVew82leebKLPCGRwy/m7TXvQaTAHsUv4Xq8fAb
jtOW9QYL1x4VYFlHMujqzaB4q3AjJGUVfc5vGVpHF9OWzHGuDDkBmjjC6zpeDtDp
ogW7SlCLmVweDFe5e2G10fT7rO82/5fcWooCc3bVwV1R3amf3YCGrX7x2awbtSZw
4EDm8iGHGOArjyCYsQ+RH0NSpu7P5HpBkNo3VwnSp7fCRRqK38hRCz+YnPx3Woer
MvlR/YsqosGDeVYZCOBrv9JZ0Jvmkm7cpdVHQLKw3ScwhFD3jx4p+6lJc70QkUPh
cNIZeZ8sVfg4mlgn60TqLV2n5gQ5UVIGnijk/43mI5XfnyB2pzvu1aStMJt7FQKO
oJgBeSF4X40GuEIHOYNs7oldNLKRuJN71LjLYd1CJZnaDlM/KQVObh1kpixK04PR
n3pjtmo0E0Ktt7PqLA6nmfVQW1NBwWMm/JQ0qRNGfnSJLyVB60nwYxYwSPwogPLo
hx9XM4eT67QR4jy8xcGKvOzvq9DFI62qJqh08GiFmzhms7f5S+eFXfyY/fMLblcA
jmdXF6pwLXIKamvUr+dyUk6wdZTMhZhN6W2S48geHEn6k6EDKeu1QKeeF7kHr1L+
rYWk9zpAvNk1gP04mkH4R2k0mZri8CgnhKECGl89BVAbT2w/uuzxWr/tbun23nik
h9k2s7el0hzgSMB2aW3QkwC8NK/wdS83VWoKNIv5xr5YECLAUBtUh3WZGJ5gNRjA
6543qsaGC6um5U9C7i+GAPhThICmfsdnF8NQtThtfCVt/CINhlUj1Z0zHoWMBcd3
mp67Ek+GAVX7duSWKTBj7V5q6mexkYNjrf34LwLDYHGkF/eRaVbfn434qbvLraSZ
fPHrI9+X4qyqJ4EgC90P1TMN5kYlO6FZH2hwHenVXl4arM0YudprImqvy/6Q8Tc/
JK82ceqZv/LCnjnCF5PbhLUzUpjR1a3IqB2bC0KBugPGl1gF9BwKztbYdKM/BhcH
AqGQTbsdiM/Z0u/lFKxpP8uteS7W7q7JdPqI1ou1+CYrzdrAHV+kT53lekPLOr/n
yI7M3WL6dUwE9zESXQSyKPQNcRTO0nFA9EaElvu5pHFlPoHyyZynmZl0CyNsj+Vl
PoUW8VrBSzDuHhkW+3oQ7QA64zQ0Zn9u7A0OdWoABPEZxCDQpVnbyMhgW0WIMzXC
2Ll1qQml8lH5JTvs/ct3TnqgwClfyWsOZ6be//s0yJYWMfqOSUVh1ltY+NVoUBU2
lIdnpxAX2BxXHzblSwVYm4LDkJjHI1qFVzeAAZhxl0P7tE6qD8LbBFKCcv8QwreK
S1J/e58bbOG7si3VsXt5cUerPjdtIxfuRaGWvk6ag+ITQp+OMFiVLyatuDcpHHxM
C9w2+bdXSwPfKG36SZ4Ep/WqBchaQ4Pn0wlsWH+DGbEGcaXt20ScycPl3vIuEYhF
/nYYsPM0HPWsVBIgSHgfSiT38lWrkuL07YFE5lJEVVgnORLuykaMWkTQEei8I2I9
2q005YYxnQrn1yzcXnJVPRcTbr7yhv+0vtSu33/bfPxizIHA5psG4u2jJl60yfup
/SB4ike/0/hTtgpzJNAVi6a0IPCM2gk5wqetW1M5iMJmtr4Cr87FgW391O7vYnRt
Xt1wCTFHaO6VpijHcMGk3f3br1b52e05cKmWA3jqmKTTowOUoK5sDnyNowk1jXHF
kJOF+/hFddCwBdcrUixTJMcm0pdHR8xVpvD93UEatXuwtzDQCKaoGIHrIWtM6eob
+EgNxEBEfyH8KfLy9OIax/BMwyQ+073SU2zQthNlAuSrjf4rzDJSZ0+TU2WErriV
ncfdsSSCnB5L5ewACxJlc3JP4/fcdBoX7jZSNbdTTc2iw3YjQzEEZZ+hw8AFB2eq
nZIT1ewmSjTgJeHJ+F6wqtj5V9uE+RQIsSZv6u7CHV0rrmZ2JGKI8vTDGujG75bp
pcOgIvhphRu3EhAeZOku9/+3X7Nniq6ALdT7+192BsATfEO1il/ijnAUpirxXdN3
pw9NwN2EhLZCCnxAsrjHVkgFuTAX71nzP2J+LD05n6Zg/OStnB5NC9nuJagpHDXT
7j5t5vPNyH7aNgq14m4x7Ksi7ysEw7Z1BBIqo8v9ouw7dFZuf2m1g4msbi4h6QOt
Vt/z0+5DKqNVhCdVqYZTeHRLnfOjzw4FvZSeXZYxU4cuBlja0LFDaMHTYnbHPXen
5BcV9QfF8Acd+9YLucterHsoVSh3ncsSHkjcmhOJQqlGO0SNbPXP7/LdKfcmNMJp
vSTnpyPL/2YyWKXTMVarrTWjAl6kaeeM1InVIqGjgpN9bBa46RU5u29sYex+sTOU
HrmZe3rS7WOG19Zt+kkVmpGaOZ+/Brc3S/eOyn8Qpe+RPgJ3aURXgUMS0liIDteO
+Jzc2H4odYrMTs05mQFbnAy7Qk6zi2VJiiT4xdJFoZ6ILgeHGUYcSN8JSfk8bCCc
bN6XpeJslWDsB1GgOJ/xYDrHczkujlKBj6IS3NOz3spA8UCxZL7A9SGoE5UyQCCg
IQpO8qXqeALUWfnGKgEe+BTKIrQoUAx/1QuK4idkQg74YwYLCeHwuHG1EO4RCS0M
M+AeSPBqddqUuhdUfEMZhqjsce4KgKK/tyHfjs2EYM+QXLbqhJnx7CAXe+iFFEYo
v1M3VhQrPENOKZhpjlXZLrvjbdru7zOEEkJT5WO5cGFqEisnY/s43uFzYYaf5Uy7
kdL4gV9lDFRu2pmVmrGHlEnLCJxYuodHMTIA7lSHkJICFkFUA8nfA+Gk2SlmA5sT
OkTvfpf/XViaW1WAlJIPtug2mhVLmOz95XQGls0gJncA+HfWMuoC2THoZmA/dymL
4ONYwbsJVvOWtcAkcSTenGYVjpbPODbq/NQ7el4xvIirtjbYCV/nTrbYAAxRnVfF
OznSr7ER6qawQ33g1y2G017EC/gbJPcSbLTqwnL6vTVqIMyDbid7RVKkm3wQXgKI
yRUv/tosKIncKoTwmy+XKPlTUTWoT5aHLpWRnWr2x8ybMdjdEJqCQd4OvBpnrBsN
Hcwt6ZlEPy1tM82yVks39Tj9Q9WBRvmnqjfbw40dm9MH4IE+xULnWiedoX5Q9lxD
wc7wiXsy7OVunWMeouNS05oKLNrKM4qWXoeY48ILINrjQpOvWggC7k5LRcvXaQWO
c/IIpedE/K7M+/j50BAfp/y4vtGmqxb3PoJeNjGMykZdvW5YsQCvCp8139I3ijOD
0V9v+Hb76OlTpcsvVK4us5JsypsugHhLmomVhSMya8ZyvlrcEw2P5MxpNGGeCN3R
wOkBv7XrmyswmEjeA/5gvgsPWRzm9SJcq66EBQndb24yJ9vkcijV1D5PmwP0ZFRp
Hf0HHrpj+SGkrK7pBUklGYrU7xliZ/61ASvhyuflziJ9l/D6qh/i3Hn8kw8R40Mr
It9DFRCcDZVYbzA9M6q4PJxnwwOSN/pBrhbrLmQRDTSVwkFteiUryFFgGrW2ruFc
WODuLQb7b/TUpbPnam1hr9skh+nrIoycCzOGy07uBQt52bwN2UdzHRzTBUMsgX6O
wn1twqqbmFbvJFt3CRYnpNle/QhO0dhbpV+xl4zwPSkWx228AFoF/1nG0A32z+lj
bXYwAFM+cJqhH9e2Jr9UtyXUHMaCFQHQMdQ0bW41fVXViSSpGiGT2Rbaefl/zIU3
jiHptg9E6Mx499Eq9oQKMImJbKq34RGWJNxGdMBl1BlsCtOekr6/njkf46V16ekQ
w7eISnn8iv5517S987lW1ff9QUsLpdfHd34RFmk4H9s/5fO/s8pD7ia16F7BfY+8
fIi/o3YoSzydQy0J74kA2ql8E0iIsc0u6LE49NV3OtvBOgJS/vHfR9fJ7mTVuPiF
W1Og851u0a1fhKp5DFw1DPVaBwORAsWdhzxuxUPg976qMbTpAm1//7a4gcc1+Lxt
uurEByDxag6WhTM7aYYI9AVPzIoFayg3DcatJhDANH6bG3StQvyOh4+TIDBTts2x
GKCJlUjaNMZE6UkO/2XwrKdgvoGCRe94OHTa5Dh/clfZL9UP88y33NmIrfNdd1fi
3am1Z7IrKbWVJOx4j6bxZzPF8z3SCP8Wj05sZAU40ttEwtlPv8VXYY5L52eXCIsz
wqCpjroOIsp8qvstSt7zPtBPDWkw37F9b491sDM/Kwdr+pzaj3cxnnXnZWFP30ha
TGdmCmoPbEdvzA33DNdqORVeIZ6MClL3tDgL4RV9fWSPNQ3RVQCSN96CYj1XExzt
JFH7wSEYb133E50Bv0gG5z/1IzpCV/sm5GLfkkPeDbo+6pzTqcz3fYTwyhjPpBps
vAGFI40imLX1UtCqwKkwSW+QnNNceVs3F/FPTvrGv2tG4J+iEnq4em6h6EHlFN/L
pJ+L2xJIxde/dfKF6Cw3/S6yGShR+sujgmIHKrZ/VaM5Pazx59U5e7gYeRzfyz2q
JjoCKTCnh2yyGjZODrm7M382w1B6XsBxYzECCUYvyewB+PQ4WovaT2HNI+huA2hd
HpdyxMmCbvQBk16u7a9m82Tntn32ALGHGa53W8uMxZcP9LSwGVpNkg67qZ57Prdl
8srs93p+luJjzby3RxjAxTlZVzl+Kxvzqohy31ryi5JdGbDKJqw/1aRGuwIZRz8X
lQIKtIi5sR7sLYxu5s+imbxYjC9Owl3ObiQjcp4EnY1dnfeOoGeA39Nn+hrPCaod
w9yMrNOZelA5qNbnyOtlTzMhL7LgwxLui5x1M93V5e0rvsDPNWCZdXhKIr35KRdD
rl3ymUC9gYlyAqns09TGqwelXmZMP6LHV4ce2lpUZS2XZU7/sQyW/v9wcY1E/uHJ
CVGrRUYWbBTSlN8PlPNYIyQ0VM3jmuPESGIsN12SMQ3CK47NATPU3YE4crw1z8N+
Xlnx+Scon9b8dWvXuoTRUj1BLr3xZ6PV8/44PZ017aY1/uGKkORtqee7oUJZmnRL
etMt8w9KA6q4zFZEnuhtU0HhiNIw6bTbDfvYA9hFdQuHLMbz7WiglMqnDNV4NC9M
MdwXwZnyrmaZwAPcRkPh3JGY5V+Nk4R/vlF6xw6ZUnu7YO2sVuzUBIsTCr1lA+IA
ZQ3OrcnOz9OVYaCdQ/b9x2F8LN27VU5fr7CPOElRGEt1tHTUV5xT3dp74lT4ZDIf
x05kiQCSO9XwmCBJVWjIGUtER+U+LjfTNAB/VF2fynoR5SBfQLB46Pez/RyhbyI8
T79GNYnYyej9R2VDf82/aXOtzwycEzWJJitjAbBTz0h3Hzy6v3quVU0l/V5h9uiy
gQSebkfxgBGeB71pFkpFUacakDxLIrHoSxdeMlRmKUNiTO7HqbeubxUpAWdWv6Zx
Ucy5RrXU/Hvd3FmrMKpSPBWMID91aGL1eMj+kzYn7d1gYA0OBh4C1Md7gQZ94nwz
LzidgdZNFbovBLj06afVpSOuU6WF4Ko853KfG6cIC+yJw73c32JCInp5BiJyI8Bp
jmEor8+eu2ljLM0rJP/Q8pWA5xg7THFq5Z5iMPbwdxRc+LdpJedJMGgBZY+JOlnc
bAA90LvGmCmL0PNzvFGUChwbXSdQlWimUcLjw7+gSEgljTemaUFn7+KqlrfnNGc7
N2vk92ekQY0uyGS5nv8jH8y06l+7C515Ck3jjeK9ij2yrMox4uY5d9hKuzBndkHJ
CmKtK8Y12DCsEqxH45jgnZUFPV8b/wk3z+uU52b9wM2zGvNF0skoMJXdYlG1v09O
ZNohXxZ794B8fw3/r+N0p/6XiLnja9BqZa5wQfn6YYi9AWeOzcdbWtQ83lwywlet
LuyQr7ymAKU2NQvUkiibvmmQkiq/VoyORN7lb7HWGL1+SzYxAWHs3rNpSnzIXcLc
fDG26XA2U6WgLXhujXLA0thjHfTqmv4Eir344jRBrGISnOnjo6wmQW9iqRbeLtza
I+/HzdK73Ss+Pwr7uDyYWvz25jbpYnLVykdUBoE3HHJ11CBNRRHJ7qa1msJQAruE
pCfLjeiJPh3BkRik9SL5NK6tVTUtuSIhvQz11m06+ibJTIjzuCqUBnVB8tM5jA5M
FRmno/h6eJ02hYBK3GxAx13eq7gvzHLL5Uqdz6JgHTKtSuUectC0v22IqFAqUoBU
At1KCQiX1hqwbFcv588b6c5lRionO9mtVL8ywR5KkkDX2v3a8L6M0xIeDxz0FvY/
Pi5TJGTZZ+g3+lRVhqRi8fp9YL5odOT2YaYibQY3FJMc/529ff6jJdNdnGv75mZU
bQcbt+3SWEnzyjM1ewibevUtKvTxqBYBUwrAfidAo5HWnJ6Fv2za4/86ThQpWA3G
pYkZt408UuWW6dm2omUN2n1316LWef5Y4KHYRP30Eph1GEXbezXnUaXeFWr+Z5Wy
VbLKWInRhfgF5oPlcF89xY/7vQWWR7YQWNKfwvuCdPs/fnjXJa9pbOrABge/crHc
K9OkXt/Vfk4LhFkMqKBMo/JTquI8k/FVhQjMTR5i50rtHOr3QApV2gS5H9GRy26+
7yscvHyjZXLwXuZNAMQDlQWKgi3+o1AWxpYRyxfuCNNmOg2fkcNKwjbQoB3xE0lj
Xky2QtEmkbqDqXB52+S5Mfsi8pmCnhPIW8xKivtLwvOetcry0Ej0IfjV6HfKk+9C
0dBt6RDWN4YLHjmOtUbyN6cL/NveoRyCD8iAWEdwAHRWsiylShTGLCFHAEwv+6Gc
t9YAvzf00FwsGKUfPLXEUtT34OK9IouG6hw3DpvRhuDGySr2jO1x/kn/6f05DmiJ
p7xuxcBARGQoRJiWdO0Y5yLR8iUV/cSzMsHqNoZPfVkHwbrJ/bXCcL1GNeRRMdAC
0NdoXLJUkfK7q2DI6I4fcEDvX8HbKz3CXCR3CRegotJcjHJaOV+ijOBmjYX59UCf
CB0Iasm0v5yWxoxWwSfJKvcASH1A2DaSjGGSnNVhwmeXAZvZVqcK2yDcLaC9YRt+
YJ9x4JFHB/3bO0tVu9KsotlnROBgSmbxuTPv+uoQhDx6cDLDydksTXVNsWlgGf79
nOTF1du/oL0yjqUozB9CsB28j9zrLfqrofLg3OzZV5MOQGEYyS1G2M1JjyNBLpF4
zKeRPjt0PtVOvG01ZYTuBjclEilzHgs3ngLexTOqTPcYEoUTUX5Odz1fZXdenzMb
CowEXcjWlQOrUatUrcY/kqviFjxtww0zho49Oo4ESewIfhA3cu7fmzxIaG/Vmz9h
Cc+PoBL1UdS54MK/izVKzG7Kmd4hy+gHP8QgWUOpJoeXzOG4jTGSRFxbgioRlkPh
wpvHv1EIbmriGoOS/2HaDFQULB1WdX53Oa4EBfrDRCvEfDZtIX9NcpRkaIobmLUt
WubyMGJzH9FfRAhTvU2qLKMR5K7cVgy9Zn6GJS+MKuYyEv45f4f8euijAMfbBGGM
STCYelMFlzHQu3Nyi3+3pYGO/7eKmzwl4hVYLUSZNYJInx2rHnEBoKbKDaMdrNMB
4u7PfHL5fwWVzY71yMmKueFEYlex8LobflBzAD01CvvWjnHabciZeeltoj40wo2Z
sh2APR3W9iT6QojH72hXUd1oUyEl8TWovp3E5HHSUhFvOdIFnNvHdv2psYuSBqh6
AuEgNZWREO8NsRIkqPrbvEUu5FuXqMR9Y31brZZY7sLIDPGGkBjfmz9VQooGC+mz
7dZLYQo05uhtCQ2C6RituBODR/fhQD4isbnZR2cgY7YZy390KayoViJ1INE61qIs
VL+ISzL05nMcXIFXcPVt3QqRbiv8MPn7mDE/2oN/OVam7J8vlATYkGtj34WoBXIb
szpcmnI7e8JiW09Hsqrz6CySw8fh2QYo59b1MZNEHCrbgWYiby6JyjtYlBtq85c+
a8MRJrT1HYi7ZKMcBy4hCCQfMjcOciqE6ftaCx2+vjKR9BNCe2lM1Y/vCvS8uVRd
0kIPU+m2Z3cRuqCkRZJqlo/AU/WMh2MyHQsLyZsEn+oA52xw/zgByyivpDp59lY9
cPcA9GqwLWifWPaSOH4RyfcwmxSCsy6BtMxk9sNeoFscxDaSp8rWT5oJp8bnUadr
C4D2I4YTmLqclFz8KkWrWmmboSK67I5mI4GhGJvNyRmoFWtGgixjLQLMKgYA37du
GNPfe3lRtgaclBIJkV7GHBqUJ4aR5ghgKwtKfihpg7TVZ4QoF5/s8drCSLqm5bgD
JiThb46Eirq0Rr+N9XJHaT5M/JNvyoPL8QfZ5ITHfu+XiAbMmI5J4k9MQNxD+lkC
NIy6L54DW4A5OujAFMGAmd3FmcR65Ep2L3+8pJwMFrjw1nF7qTitwk63zrmwaUFX
sPK86/SGlqalnF8WmjVpx4VrEsnmiIbgJiLQtDtUgicwXMcUvep3zOKtKwtUhN5q
Kv0vEkV8aWuhW4887N75oFTVQEvsFgi941W364wYZ5NUOa7cB0rL9nW9RPgWN9mE
abC4x6Mv7YqE2JdtfXoUQ5Eed9GllRaog0Lf9lJ6MkULj9TioqCh8rPtTHuLNr2U
JxppGqKH0OVCWYH7L0jOy5uHyHbL5l9ZJ76glsQ0f5jwv1JdrwecGyKHuydENCja
/VeDZAhsMLGCWC+w+dKudDpZWKH8L6TAcp1FgGpNnFC8CKKNgzfVRrJ2J1T7n7q8
fAAGtiXCr7Hgbwl2H5F1NDseTjGF3ypLO2ok8kVQz0uI9z5ffS7osOYZyz0fLMJC
dwcJTyxVokaUJ0Ls2EcdLwshGMkRDKU5p8Wg2EWlKAKsjtpmLf1xDG2csqM0EtAJ
ajmGrv8Z7ahturukiCMdK1cmV/wSW0WevSoIHHQnN2eNaw9REd8VrH/e8VaWg5pi
tIM9msr7y+GUSAzVI09soZQ/Dj5Ix0bi+JyRi/lrF/VFn387CBT0vw6IfeBn9xph
59WRZ9Iadq0X0XqMytMFkRwSBn8oyo7ohK1rmyX2g4sjWQ11RyHPe2MnLbmDtBVc
K9FqM4VVyrofxlJJ5+AYXoQs3dAuCskkElploeqPRdkU24zO0nro7klyeEnHJgz8
dZsOsYktYC1F4qWwX5jP4xindkPYRq2mNFbCzDGNGGFNwBguVqfMIiXKLZT3x5ev
v2wetJMivO7dGbA6fLOsb9YVrrCDf9XTXqZO4JqizTnwNwpr5KZ4/e+kufHoKl54
2Mor4hE9RUHTkBaR0d3gqHneNrbL01GoobMDjVl3NLTqshE+wgKYTwmGpTQkFYzz
08jyNVG/6TWlAuqMyT1MbbYE/gjIoqXQfjL2fpQvXo+QX7oGEvLDLj11NLad+JOE
ctBEHGSSBCsAzLl1hDgdNtt+xUrUjK2974G+UPqlBlEAoTt+snLSKJ4mqz9Q+Ion
GgVdA4FQD/6+YMwnffktgiMWXL78lCdmcs4Mq3UEs4ZRa1S0lm6+ivzVjdedEfxb
/EuTZMtsLSvYEJMeotX5dmYcdfm8r9tnndPKqFbcz0qhcpE8RtWFh778BLVoxs4g
j5EAPJssJcFDRv6lCn8npY/Gv5J0ohy/IUlRSruwYXHDaFlQdAtpJUOvivpRNHxj
4l1DJcfyGwT6bIB4WtN2H3+cbfyk8pDGMDwH3w5ZJ1Ebsuxsp4nD8jT4LDmwPItz
DZaig+i9yidBhzmfyIWI0lewCd+890T/CWGKPD1mYpdQtezqU6o8ZqqkhEHjSXe5
+bDiYxCiFxvniUNr95sFCNAxW9xGRUBzwq3pKL0RfqXUkjH0wocIFalKPiOLMvxl
yebGE179+1OCWzZoUxBbHvJ+ksHqfgpYjW2misVKqfagYveBl2QiIaxAver4WReF
yrECcE2m7bZRkgtXpYwVXodu+i2+KRIUyQbPzg0OobLdkFREkTB7fYk9EFqYB+pd
eOXLjYEYPmXfwiOTJRGdefAoT2sVGepLGugIFaVCzXl7U9IK9r6agJVkySID4lqN
b0cwevflMZMRxm0Gum8jo5UZrkal+v7FlFSAvX4FmpAaMFoHIkPHvpa4xwnptpJr
+qLhB5FtIS/qZKHMyNRYNZ8gpX1ocpUuEKs004n9zQepz8ED0ZS8WGI+lpH3QBj+
d59AaXwEnqdytRsdWwVw6DMM9MP5LzRYtoHkLX45u9MzmFye1dUMf5RkUoZ0EJd2
KVKmwavnDa5/RJUQBeKKny1CHDF8CFt3B66XgLPpG2KrTM/U8p3jhv8d2dg0JGIU
YzKunZxTtcmk16N5Lt7fk24J7DzCF0Ihqh8RuiFSCi7AwxVlLAP9NfSlnoybA4kF
uaCeaL4nK1RQKf/saoIKpfsZ/1IFmNxSEoLkrdyzfvhNu+appZPqzhXnpn85Rws6
Fqymjwba3A3LBbEpUd3JnqJXKqkKqwmRdJsY/56bGV76f+XAqSoYiwE2vb4a83JL
eAxBqWgkcjCbE+yuoiQ9fhRdt0ygcHZ2NsFLIxWP8g/sR3G+oHZaezOuojc2dHRU
KyOiJC/Qxe51g8cXMKGI9O7cY1wBKXMGZee+O3GvhauMGUwmEUtKriG8yl2quXpG
fTpOW5F7kxfk6ckZ+slYBMd45RnUThs5RdeOrc+g7L12d+Qz3er+0KgN5/rodppQ
qSZdfOz6ZGtXh1m0Pp4VDpUMzU9EI0v0189jYhEiJgJOcxGgMWtRqBV5hbrH/QX/
o96RgW6FC0DJ+BnpGHvgLtqOuEDLTWmOZlG5k68eiNmynLf+CDH6vc5ZIsn8kBt+
anC00DpvD+eiqYG/p5QZFp4s/q42tPtLSDzyJGsD6lJ7MsiuZVAGZOL3WPvul/od
Rd+h/CxRAA6sY83D0S/EbTWDgteLz/C+YNPOin9ly9ZREgopd1d/eHbId2+iqwAm
37T2VPotPCHyx/rbnBT3/pXsh2Fvw9IWpqKebUwBZ2PpbCO4MTyTBZyEqpSyIvgw
Nk4g6OWxsRQdp+hgGIRUoLrWl8bwfoJcZK+ld0psPOV1gk8bziTdng4vIrKsG6SF
tJh8lAKWloDmOTBMwGF/Db5HJfwcu8qdANPfZXphtjIR/dAg/L3lInCQ5sR1AeZD
n4lgxzO2W4RIV2E6B70fzq01h9wfPcH/3NOU8x2kPD8/9W57+mdonhX4KNCY8Xy1
UxXtGQ8eqjJA0OFHMw+RpDuUYNyM8MQDKgefl7VF0iEuI0vLPyzLik/Kf56VdQlk
nyQOE7t9Esf1lJ6rTW4fiL9XZF1zD3E6XgZAKNOvkfQcpgGU32czMLTxNlw8i8JR
1bhl8M0SCxlYrZefrVs9wPSjKiNsPds3miThZ97gkg2NVVOTYUo5DK3TZpW9mRNp
RWd7qkRuwIPXwPm6mvX23uDFG+cNAVV+OUXaaOGloBGoBJPr/LSoKvZdqIRApJHr
5b5eQj2yBc5gaDDzeLo5+KKe0V/BSFN2240h+1h49JnbFb/e03y2QhEYkmXUk8Ts
MkgDICEfAgpKx+HkM1zy8UVLQSFpynLcaX5COWkDLXQsB+9yh5fGavOUOcbmw+qD
T4OjvtlDJ4MK0rERy5uA76IBLzvmwyueNrydgv0wud6puGKBm0a2u8kFE8C5TmIB
3UsgP81ZcCJ8n+YbBs7e6sIke2vvToIoHp6KGq4W5AS1j/FWwiGzH8rZgNUS0L4e
ski6Z5W5sbzZWKPfWtETV5R4FwwO4PCoxe35FT+YLkFOXN7gbLTy7cDpiSiT20g2
Z/fmlweLQy8UWqkC/+unwuaacz+hH/P2WhWppsCdvpXsJWqLEFY40qsjnc4sNJNW
4mLW73lLDc6l7IkxMkXxtPtz3m+IaFbr+CpRQVOCP1nWiJZEkpYJrzHcmDOS0jVw
g1at3kONpxCElw/QgiWptTzzc5dmhQ6H9SbcXTLfxjCrckoZmVw3IHRmogryigZ5
IZ8vyLEg5Jc8zPCH4119eSzU+I0nZ32/Mj9554yChdBSZ4USY1//mpKvFqFsDVNH
56YViUEPQNG96aeba+6cTJt5v2go6XCgvr5xAaUl7PALRsuYESpjOtq5HdXi1VuY
xaBQe/uXLKakeUJzsSxMpk9Yr/uikBqDw8PZNJJyGcFbPGHdSpiXKqKyz93te7Qf
a+2SYz+Zcz7l8WF76lkA+f74roEGtDZZdAbkXnHgbDeffnLUpDuXArn6VqGvwwWk
peHFLeB6m4iB/Asf1/7KOYnT3uJEWZPD2nvd7AJ6Vhelr5pJrmmWwvfg6PuY9UOU
qlDawmx1/hiVWmJeiwS1fn+mXu/EjGiLJiBzT0VVd1buWwda/2IB+e+EVY4mo95a
Cuv7rfNUNdWwYI6cgecjmgzp7WKEpDdQsTjTl1XotXk0JKODSlgf3ffvVX7UyYHi
fIqBUa5Z4aH69NFa1l8yUFM3eHQgN2aCSDGy7rgBR18a3kvAhgIEJc70l0BOqGaY
Kz/w5ZC8z/m/xuM6HB3eHt4OAVjY+q65v54gy55l6PnjtuqWFc7BzFyT1bnzYNf7
YXdzVhaQ6y8gXhzvRLiem78hQTjYUoFzzQPPM4Muy30XhtZBJfnb0qMMlYJa7jgk
4/BuKr14t6dBwSiSrnTqIjl4Ia1iloKKk2roqu6EE6YaS0Ke9siNwEtLEcYVxgZ+
6bnhXRmuofbeSHB0M5dU6tRyaU2oFm4CQpmj95SUyxKahq49B5HRc2S8s7OGldr4
En48PEH4CNov9rn5NMiTHaMmR3l032qeMsmOo2pMjPiexTZu3q2lqQOyaxAnvjPA
VBqB46abECXMiqEGirlYMAS2ACscSUu9xCU872jrkVLg4N62Z83gZwAEoSkt6PWG
FjkOpeH2UhLWtHehj1SfHOygCa0B19TK//bonJm/fB5em7s4S84kDtCdwxPHte0d
g3CoJSd2r5dAK+v1Dfk7JT8xidchZ3X2FwI7qMi91AHYeJmOHLljUD9X6mYL/Q4s
YCWGK3+k64TuGEf02RYT8t/PCSmhPECPXDlkzNsQhiRXJYW/Oeu/47glYPcjUy8l
27IcSphiMRdhbXFPZ2hD24WCxcbDLwdpstbpGJvQT7QUYUSV+jL8lsoMVjy4o7e9
0GipdHhvr43q6lSizcQgwE1z2l3Tm0BT1GVpdefsTI7lo4J1AiVT5tChcL9DQe2H
s5V7dHt0oZikIJ/RS/s2C1E9Z16wPw+BFNx4oPjiF6GxPxDGm67Ww+4SbrgJrVxv
Gr/wiGyw02OfgpkbDE6jsxrq8iKaR74BG90dT/LenZUKf7LO2XG61pPbElR7fHRQ
JiwYvl8/hhTfujzKWhI7EvUl4fwCE6Erj4tvsdVrPpJq5OeNU75cCQr6CbXxccGG
dQZlN7p+r1qz/ooaiZgGxmGRiH/ybHG+hCGi8Dw0AoTahBm03+Ylcgzu7TQ6lQyt
zzRfz7AKmg23+fFWF8YyRUK18eJUwwie9ICvmwNO5bzAEsjS9Mx3Sqmj4DT9YW81
GQX4dL2Z6F8ZRbvR1/asmQO4s8CSyvusST41wUsxV/h2r8O2WUNdiiMy+gObhNzJ
r7GUirwjLb110i1GwYRJw2kF6E7J3xsI/cpv5xuoub1q/deeO3GX2s9qkpu3uLFq
jLmx2/aECL0TYdLHbG6iki7Bq3j2I8PiCY5vasdRS7HjmDQ+oLKSyiyNW2UDVaOG
DkztQBklNRO9e8kh/zQ5W4bJscLoTb5Jt8vBRdTySA53rPtKRkZYwCebv2vaJWvY
sb0fdNXJfeXCgjeLDavTK0IKOu2qlHHG+/dNuTu+LDDVsjOTjtdt+H5RMxmFgQGj
T48IXHuA0ZCGeHIdRLe8MvLLaN848nEh7jT1V5KgSZtEKXkf2YVQg5Z+c9fgh9D/
qYIPwbk5z4GGMQCf/aGn4OCWxWB91S5ZyAm4CCBrJhK/lMve5DKZRuAoUJqedz8J
+8ge0cuosyGjnA1FnVfkyL6LXynhvuC5tk4rsw8iHhkWWrgRL2PCFXJNqZiOvgkI
hbAOkP81AoN4/0+nx5DenFyAXe42+7P3PlOqanEvHALwSJo+v3J1ElDX7+n1qeOK
esNpT4RujAQL2MGRPAYmxecqsTN+9m8QK88vzXdvWwM4kS5S+PZG57R1moQJ2fKf
Q8ctaXcRA4vFTQM8Pxe4FgfXeTEVwdMb43rhnTphdzgPNGbuF1vFk7OrhWtuQWOh
BWZFvubg4f56t+trp6SZ3fRzZ1SsRRREHDR8yWCb7zrtV7HU+jUmRDsipKxM+MU1
saiP9TQq2otPQNpjR5Wt+PRBfg4dEuih2X7XlizBznDVfKFxlPA2LlUsPUziBimg
J9uxDFiYmG+ydOazV+AkHNW8vZ9QAokNm5eF+K2xXlB4jblwuHh7TGMFk5Zi4+/e
r9ObFkLPcW2M9YDKo9F+M8UKuYurp9rJrb9D20IR6Qg/HOcyFtShPmwOraAkGoHx
tIjG+cPEPKNm62oCrgUwuF+RLxJu01mkJJkaXLtuidJjvUTABKP5NJw0nOk5JgB9
+i4oIOTCaVqfVs58Z6vf46pwgGfR0Vi6znEmj8ZZeASwxB913/jyOcZuf62VtCJ/
WK50a6hOFfoleHBH+mPhZBGqwnEiCB+1VOhSIdy3KOEKa0lXJqXzrytSjYvjOTrQ
FGz86LJxGHNPdtXH6Hp58goFl8d+xShSdJV54UIkkL0T6Lgkc/tKOFUWGwRwA/e3
I0pzmowyrOxFVIJ89m2ifBMMqCn+L79y2Q1rcw50x+6W1JfsXTR9zTdqeNTTxlYz
VhAhnuJDfWeFBRK+9aBzt0rGZGoMtxZ1QwV64LF41Yv1UgTTc4TkfXumL+qAzZ3B
xdCXlP1C5l8UxrKNF3ZOnltn94k+yt/x5j1fKZxZgrfNqUOMpIn7lCQloB+4TgiW
8w6eJUCOTHZFNXT/w5djXOGwgm7KZG5zSrPg/5+L196PUjygWzTIhOZLa1L3UvYw
0qzC3SLvYLKaqO56oFWjKT31bMDtEyiboZxIUnLxNl4f46YYGprqN2fuUWacCROb
gy+0R3rBTVkebHZ9uBSo4zuB5ARG4PfgDOFn5UMfKinnec+7TVP/TTW3SNzsql4U
uOz4RMq6VH5WT9f0D72w/9qnJ4lLIKHWWX2SkH7v8AdoMp7BVUHujula4AwcpvxY
BGJAc7QoN0j5wfwTftASZNU/rtjScFxr8/wkqDB53PBPYNm6yVma8FwhHRnNNEp6
+khKrw3xqp+Kt7Ye78Cp/Ku74UnCGD5i0x5WBN/s9BzNmPWTCaZyFxvyVvnUBQ9c
R2CZt0VlT9xW5TeZiiXxEHczAN3PLggdCq3m7IJZuYrP2/M5x3xzqZS4uGXj+jTu
L8ZUTFq16r/Tyqq+caGw3lzTQTdO7HTAMvTKxK1o/H6xp1+CivdVi7PwpMpNCZNE
JJsQj+lHBig4DF+7kM4Fx25T8xHWgiWMZ4X17C0G7BbH9435lW9bh2JcTpuHnM2z
v2WtsSmAlxiEiCSb+m5diw2l0FDHwq5DY1frRLXiYm+W/olF51DhA0qQfVIBsaSK
jbw9foKsIovCpR4rFge3IIwa/zOciBxyUMzpxopYwyh4nbhOBVodPrVfAqf19MA8
0UhyemVN3umhaGeNJSc1RWb3nrn7++d7KxosE6kR6eVT8bOWl/frr90cFpkUcXpV
zJlR/xfLuL7+sl714BF/QjcMZN4q/CFiPG2PjLByIreORvk9tw1tIkbYshWhKXg6
gvOa5TENpKQ1gQNn0vYFCv4SH2lbwLTfikIJecQdKdxDgfIs8czAAEbbux5GFLOv
aCPJYHzkFwMg2cmT10xOAL72fkaO3e3ASYE7q6nCLhXypZGT+bqM+2QezKKCsobr
5UPedRizRSe+g8z+UxMMEjAxuisQPFb87DfI7CJK9S6+CGaXOFvDJghI1iWW5R4S
Bz+zkIevlCZ8cnhKEYo6eWO55MYxfNZoLecxl1SAQ5UmtVblWNHIqZ4sArDzRvC7
aBd1szSCtB8Na4j8096FzSgP9DrNvTK8mIcn3sLDj2hzxF8KqFdQ7WujwQNgmNYK
kr/iP6JxQ3pkdIYymov5VrNLTcCFO5eppAOB0UruRffCZ0xaQ8A5/ueM9V5odNtz
Wa9xYiUAwVepx3gKbyJ47es60f4kae0crvCxCNL3Axs37lz6Lr43hAP/rXnoeVaO
DFZKi9ciUptQ8lxTQ7Kjn8Ldr2VBXnoQVQqZ1b53Fv4PVb6WoHvwtTSPgn+8WACS
wD/7yf56u14npJ1D8C/Fx30qCrfTkldtbHHdBtGW4BgMk87gfXSBStjdCFU0ayL5
TMjEpyBFSXq9WhZZ7S24pxfmki+Dbe5LgpN5fbg7ODxzM5C//HqjjaPSez0Rn9+g
4ilb5UZ7Geptyf/RtJbpGChJDDgA2IRrnmYdqiw33vpjP44a1eL8aJ79AUxBtTUS
VF5Q/zovRb82QhJL2X1RPt7fO6JL6gYEOwxMVCumtPdPeo9XYL4PmPLeGg5P7OVe
u/qIBAJ5OpAeEeelgd4a6//gT+yyiKuu+nXzI+O7pxuQ7Dk8eUkffBnJXY9+81r5
yzg7zX48P/aH3tsa/iagu+cL1/JRiBQDM/NBuMSoEpduvGH8QDUjGid941kQf92H
NXkscF7yR8fJKgWTU3WqF01aPjbx3avsdQsxYuKqnOPIcBXRI49Z9SDRd8PBFEbh
mt4XpbgZseV2u90riEkfC9ZtZaxIXDNtXbJa1Nf0lZ2g1i4/jP11f46S/Uw3ol3u
TirFnnC70Xj8lSoeydbXRMouQeil5uYwBeBf5bM7bce3/8005YRs1RqecT6FPVG+
Z6eVgQt8tIopmGRXyB3Hh2HtdhXkigNF+iXcKWXdPUs7pV7c+2kj3CqgQkQ8LI27
PkQcfJgC8SiZY06o8yMgjNXVZf0HMUKASDgPfS+uI7o/mNXSjXqVqU13fwL5/Fb7
NE2OJ91n7CkVo9WBwRqW3SIF5UNG6Zn8KKeYGIDWfrE9TieL7+9Bwwo3D1EjOsC2
I0aw/tAGVisMDTz1axZw13QR7D21ksa22JI10FknYscnuEg16k0Wlb64e+3ebWmq
W1tHNhbAWfTTvMJzCBbDrpeEcb8bCHfr5famTG8gpcIAfJfbJGct4fbhpLe+PwXW
VwMr+oPyP9kqYdu7phX9supuIicyMDs3im10K9k+Tn3pgi7mttSFl7iG94U4Fenr
rpLa8TWyr9NFLVVMmMdg7IhH3ekg3qiRSewT18NA8+8dcjrffa8p0iVe1OfNHXV1
ern8Mqj2nzOkkJclWq66uwlKjPsATJiqPjAFXP/ghofe1BwPpBuLsFney715U5DJ
to/21+8BsPjxfoBV81eirmFLbQNKc2802ty5Q2wfecuWvIbGdT1GIdJSiqa1Oc7X
oF2c91YFMTMtz+bG2+TqA7/ri71qRBKsPip0yg/GS4ABaEutPyXkw2wD9vKnfgi1
SoTVayqpafZIYONbxSHZyHyEwS+87/DNnUYAXRLlxUmI8+bU7dGQw9qnZLJ3R/Ae
CaiHcHxmL5Oas03lK4pk6O2qNUtEyB7feAcA6fKd6T0SNq+ugPfaZVi+MiHey5tf
WiOug516Uu0GHvpt1vfcC0L0odJ99Q0T1AbGmgKPJwYmy+emTxVv4YZJfAINolQS
LXIgtZBqZVHWNnnnZz3uZv/desoatjcm5ty1v5nf8nyq8AdlCQRnOeVuK/6wJMH5
W91yV0hH+FZpz5piJ3IlEkEVnl4fyj9HurFszbpLI72NSdWmxxfApv6vk+1eFS+b
zjTpxN7LfohuWnFLk5Q0sw3UArGgj/fIto8C90O2YtkqVP7Thp4ZaQTDJcHc6krs
z0YwCwgHEAdMve5QrPIc4iGwiv8TSi2Mz5TWIkqXmFxX2+P32pPdN27pvfZ18bsV
U+6LqTHCyCQWI4oZSRCmcAV+OSrcUFvXtyyfBlwSAF8Pco+HVieVkvbOorGv9pp6
LQuco2kJ8LSqQOdXyYwJUJuDPknZKyX1QaiC3ux+3FCozlAmBx+1dPXlo091ysB1
9wMfiVMBWz4w+02w5WlX3s5li8b4SATU6kOvtqoDpg3yLaMkLHw/H8aCb+D4TG9R
CUZotTIsTuby8d/IRkOwbgjtidNXiI0xSgNOAomEfeXiS9HCux29jTkzRgavkNwl
x2fOAV6Hf+pUQMWOUV6O2k11JbgLB/+69pIiXfnztcITjZfA4FXLEForTQBPJqAs
RUR1VX5ZmErBw1jguuHE7msOUGjVEVxC5c+Es4ccsZDgrp9M/2PXJA97HvigcVTp
nn71yJd9OhGALhZMUwJ0+dZ7Bpzhli97vQSyJ2LmV4eDAAGWfGUy7Ff1F5tELPgK
xoJUQranH9ZnI09rN+Mksfs6MO5hBGr9EEox4QcOpqh9ZQvKdyaRHykb6NgZoKdD
N29l1KxeCf9pMHcvTiM5NtGact0PzkpeQl6A7Eh5MAFFiJXyAMPNpkMlDK0sUyG1
Ksug5pSyvm+iOkaSVPtomri5YLf6sRQjYKSqwxyxtduyil28pHSiMXDigA+dAQnU
AwWWlPYOlR8QmgAUjP1YAT7ZWnSJiuaaIRPu4TpC+51+fg/9HXL6WBROB/nR4XcF
w0hxuaWb9IudVXxQ8gK9Mlyndvk5xcFU3iPn7DAvyGlFtIMmLjHHA5/PKFlLu0Ot
uy2bh2JASx0oo7U0R+7hdmKpnNKOkM0mWfGIh5TDQwsTvdcHJQU9uIoO/lMddEC+
L89JT4Vi6NJKjYDnihBOWllR4FniPco1BKQCJp8jw7epddSxKvcFX2bMG6SWPKoe
Y30KrR8kwclBhYDJNkZO9GUoceehs/2RQPa8eXD0DOvJoXgB5y9pY/4nsvw5IZ5W
21DxixQV6s2Q0iAF5Z4goEQFiXYfHbXnOWEvwiajwHmAsQIPq3BKk4cls/crR46t
st1LD/VeFtxVlm4cdrOWkfbHuGr2PY6bpEBjyU8HaBYLDww18GN855VQFlncXMtC
IAS6n1bjTQ/afW3iiXzzWwsMcdf9D12HzYutmfUlvt++nybbThzsExK/r7grqKoc
3IfkQgKoqi1Q75J5v5B5fJhK2iCDYigBF+G8IApahvPOc/9dt8tH63n49+zD52pb
StW+P0LaAgRrRh0GYxy+7Rjjtva58uzecCj9b4YIG1vCcDrFxpP3byScBp+qAPH9
D0AVrWSaCSUPhx0M0X57R914sVreatpdo93Hm/+IL79OefBsp2u+dRaRRryVuH6b
U1LQ3M/dLsf5NjVK53yxMOx7XNB5yqK/r1kC5Pn7TGjWL46UFrbyo4r059TLgOs1
QWxu5ga5i8Xs29WAZLikIhIliYJVvepfnTWWeh0KcwDSe0Po2oelwVsN8oqACaY3
ViMkGTLpzHZ1WGQBIvKv8RmTUxP4lcQ+pyMcP7be+zekwkDmIlvstgVSLvV4r5W7
a/zDgU6+pEfUtbbDeYhxCkA0M3pGfQYvJww2ius9B+LxfG1vBogpQyCC1By3nFFx
jPfcdbM/X6/YZb/bczjgSTKZ1iIY04wsKtk8aNBvpV75PkyNSkmWZuLFcw2hu79H
NT2jQ5JKoMc+cN9z5Ge4Zcs6cJUS1ZhAqU5YBBd1eZVDp26fizSHlhqMCLmA4aM/
73KE4R70gRAUU2BCvu5DVHkJJiNgtV6tYo0cqlQvSBluLXcICGJIb52qqCCg4OHI
8vG4pRfshgL2w2hnMwFEzUbHRVy4sfw77y0Sy8h8DdRCloiWdalAzbIN8UJwUlFV
R6oK7QlvbIJ1IGxwot3Rhv4pIFihNWYr8wNBkffS/NqpbX7fJi1M/jseHwd+y7gL
Iy28UmjT+ZLqFCqslZXOjRTmaAXPlkPRY9RQnRANawba+Y2YZmYLUMNVDDcnWwSp
NVmWtuygk/XeqstpK4oZEgUdX5idZwOp5HRjEasKLhs56mOk6vNSg2ATpHoEI8zl
HjX1yvet/Qr7xbyPnIItwdpuu5sPB/oLSpbCSrnZaNu3d5R+eVpsb6P4aNh3JpDz
wUP519qleRIp2D1mKKOJmFjZLdIpfQxyLxW4yFCiKPnLXreyWAlMMIaLyX4OIFT+
QGIPp4uyp0444wBAJw7CSOYOzJ1VLWZvw7JuhlVZRbnZjsgg8Q88yVcd2Zp/5Wpn
qbkLRmA6EJlH5xL7+ZgUq8twOUTCeXcpaFpIV32qJ3qiOdXTa9VXaN1XJYTzfwTV
Ngsp5rCqRWHm92KYE/TxJBaCnBloFWQrGXKCnQjglGJ7KY3Y/bjM4UUSZR4rGSvf
6FKkmxy1Kl82wj4KGWB/KbaJh1Ckas7FLChr8vyqNEZZaRZ98fYDv2VV8b1Hzj0E
fb2fsaCIFiQ1f0Gf/DV1Bf56zrb0LSnRJc7KwGgmjN+AjO9aHHC8MyMG6sjt+cnM
AZ2XiX4MQ3HVUpOg3HgYFw+tVWjaD6Xa4XZS2n/b1yKbK2b5eX56genhfyDMkhce
577gqkkCFAHgtAim1B0/22IDCCnk0F/Mu89KI5y9xJzP6srjaPT0FE8jN08FWCa2
8A5+67BFVyz0A8HqWpfyUwuQnxgrrlkHYj8VgToOt8iNVF5nAJm6g0yY3fH9M9Ft
Igw+F/Z9xojVRXAJG604bPjy546UZh8xygb7CMSNltNywxgupsBvtW/diKuwi7KD
MwwVVvbxHbWsUAQ0+6xPmRtr4q3ZBVxuimmcYru2j0etKLTkKMbt3bU3OMoKFvpw
Q+qMqNC1teToHlahvXftrBJUFcFmv/kBUmioq+Qqus1esGMOnYGXZFbr1tQRrEvQ
6AefH66Cj5ko4z7dmCCMWiuGq0bCwjIHdTpbP13LRPYdpAvVNIHeGD2UUO0zbfU/
oFtvxpq84cyCz1qdX3wJ4+I+RzK3ZqmNp5pXanMgkfslipXdFA3PRbsUXWuHG3L7
gFCWnmOdyKyvLWFKObwHV9ieezvJAeG5ZFlJTvBE9O77sEHnQTXzSWmIAX9VHfGK
6oS2wM0yk1xGMxYbx6KrMEyOhWNN4wWnyZJQ2ANTOLV6lDcFL0L2VSC0PkFAaU9S
mQguCw/8tpMNH4xNC7WDtaFdo1WXri29uW6UMh2q9YxL9/V04JpFpsipwNL3MFWK
BVTt1WHq4baBAemanuSFHcDWhw0bTgCnmk2t172zTtaz9pGrvT8Ikb3opazdQwDs
JxhSVnischziBKEdAM6OCtcfTxnleBnXqDgS3NR2Zv3IpR2uABl70byEjQeNSrUI
SSIxmF9rieUK2FIe3IbssNb0hZtZMqyLgeac79WiNHG6cqfDY71otFDykFW1VONz
RbKUwXuTDxAvfWYSVwuqRFdNPxUqEEu3+zgtK39S4SZCrYyj0scPJkMSZEZpuo43
KsflpnEjyY+sZi2QMNZd6b2200WJDSQzvuKlsIH7gwH1Q4rXXkwxeFxKTmakYRaU
4ZFdhrB6UzqXp022SMZBsvU/X7y8AgMR1D0U1u6e0ldX9eT2omZWuMbD1BqRXpd/
ql8cwb22yCmS2psx9TTvyPnQ4zEvt77IuV4kMok8QXVbKUvmOS0q1blEz7gLG3LW
Y2nNuclCnZ+dnAxwE9abyncbsTnsgF0ZmGVGD0jDWeFjVmxhffWRgDWRlwLsM80K
+qmFucS6qFcXm6i4rOZtgWLd30gEInyZI60dy+ytOPVZbdcdX04+XnX1P9PEDat+
frK2giKUw4ZCUFy/eKRkBLW9eMywtAs2yUnUGHuzUIW6/INvYgl9N8qWIe+dlrcY
l0fm/AZunaip1MDXvDHgNWNS5Z6CYFzI//A0jzYYQcgx55XnPmrnxz1ZsWRVz3IF
r2yAIAu+xacGGLmOgXgGSSCBzKEaxVLo8lIdvxAd+qPSPJYR7pG16g1bf9DaKmjb
h56uZxwbkS7YBL93qT8JMVUcJNY5cwNoMZOyRsCyr2lbo3shnftOBWKISVkSpV2g
SPG/eyeqbQtDMoNLw+aFgmKQJsmNTI/iV2NyN+Tg2hRWN+srVUodjfc5EUxWOTj+
7CWjYSJQ2hkMoqBxkjOTNRbWd34aEh8mlrx1cSYlydxWwIgvq0HdAwOs54WTW7xI
X4UeiiNx1IkptBfZMUaJF6Y0W/df/NqTZ+nYuJrbVSfa88cLCx1KfLwthLzQnSht
BPFPnwieztbMdQ/xuLLdqXk1XzJu1CWh+Q7nt2MhEGgmATC3toxZAqswdBThCo0N
F3cAF24Pe8vflfm42gCnXkDBfKGuFvdhs6Lo70A9oyPpagOH9pYFapS/cZ4oHn59
pm/kzv3fo2hTEsJSTd3ZByPsqbrdN2qzwSNXZN/eQiTI3In0wWVtZJH13tXhm7iZ
LeLbahqy/4XvjKp+9Ub5S5EAI5FBlnqts3cByg94hxaUONM0WVCUvIYxjjpmGkcB
dBg+T4n29ursyCD3HUetGf8bRm1eyaeI0EFQLqKj6FfLXzFF+2seAOEYYySwy/Uq
L0tRhlmBU9XMxfb04OjpPeZNmJLm9JGE24Ld4ovYWtFUvKJzsjXKYFkmfue26gkd
2r1gIcMrX70dTVFMjiJmo/CAAQ/UMq7PYzc338WoFjUtxSjXqK7mncr+9F6g93eN
o+XONF41c8vHk0m0O/WUDJtwDCL5nUOdbaIFdVJrwjAf1Q9ZtI6xJ/UcJlkPbZYv
V0t0mfTNVZ9dRnELcV5DO8ILd+P5ON4Ve2hXWnXA2bowwnV/pg45iMiRmTtGz/nz
/GHrNYLXsT5x451qJdeh+FMTXjP/4wV9GHSOFZ4OjJYDabHnRizs4V7oAYUoiLxR
NsmDOJQkt0dUlbQQPutEt9+ICLvxFjb8MAkQYbuuO2N77wRRufgLtV5UgJUaTUSL
Gj28yNCYptwPoxtuBsKU7U/0GLA4i9Zu2uELRC5ryAVAcA3+DsJHpEg3973k72AE
yyzq/ofcJhfDb265C2RR0jvJbQBem28Q8imMba+8eDs/exIC+0W3g8UaXP7VSBTo
Na2qPZdD9JHSumVJVS/42XIks8sP7cb345YWRBd6566XR7jRU8WG0S3WxtqrIlX0
1USFWRdSRyNAVmeywGj7itzmOdKP2JfvF8PGcRefIbR7v2s9+d8II0criJvdRX7r
fXEHgiCY6isj2xwlwlEpXclO2dNwD9RGqliJXbNrmIp6rZja5glbDzRPLKuWqhB8
J5AFmZwyzXOr0U4tbvzSd2RBE/DsFs5KnKhHd9ODrDi1Ji3IEwkSuyXqaSbx5R/w
J0ydGhgGBfukScbj2dURmdF9hY2FcY1HdR1aaQmMmmbQmAbVCaO9MFOx4r7jDjkA
ANnHUbWP0frapPNDBFMDxaiCrGJO5Jyb1is9kWFbJqDxWKqteANkLUkNVrS5L7r4
cXPICM4FJ1JkkfCYDHaEeexMuHy2gsr1n/9zLxH55QO9W14XlZe2Zqto9/mBFfBr
QieNPwVscoGzAcLtL79j1ubFR3YqjoI9qh9cvkLlj2IefViEIPiSN88WPkEQWUJa
4gOtITLdNvuFlxjCziFTyAVJhHgeAmjCI5zPJ8qokyOV2qHnWb2y+LyzATZt4yPp
8xmIJVONo7m62wolI+UZvinmuVzCs/1MqqxrdyXCct1RogH08+iTY43Kq1NHrZbJ
FVGMxhCMpx++u8BT7r1XVCJv4kZINVypoyAq197YjFj43pFi+sATLk6NeYt45zro
1hEyyOExGZN8dReA3LmWkEx4hXq/TI7XlVN2FOYUxW8RgVm4fZXJqP2FWjEhtb3Y
8O2g2jEwules2aFzjMZLdjNafu173a+bF7sgTF4wE2dHSJmcNO6LeYnOWLDhl4py
lo7tcr4MyIVO/IswPX2PMkVl5v1Vk+LFiOa5iChvDexFzh6w9v0kK7QgExPkVIjk
QIpRf4iVWCvi1f7shx+YdWCIlyoDaUKhDiMsvQLUly9ji2smvmkD9LjmbYazfB3Q
0sydMQ76Gg+GaGx2TWLK/DDM72XMZn9zoCmNx9qGi6v32VKaSU+xDc2bK0Ps2qTw
uKpShyeN7yLtSQBpWMYI6ZZ4E9JT39qBKldKSZlEZHA1hdDD4XNXzHsRcneBCRHZ
BXKto8y2xvPLTwT3gjMcWZQiKpapBYKGC/SsMGcjxBQgC7zCm3y1EmTbPFr4cBzS
oJAZaJkYvXEQPr8DskPQ140Kn2JLklLhuLPD8ChERIYlMjn+uML63/kAi3XxoYGZ
CoBeuCWiRJo2v7a1VhLJt09oKT4J2t/+5HNZ0qpiOFhtTrGHGuypyrzBxSj0Cv7F
up/3b8D6t/L+g8I4rKCy5Oz+w5GqN89RnPlcTWTXVf4SU0nFheo5Nasj1gsTNI5F
3SatQV57oaky0MPTqT4XNBfmR8R2/1XUMP3YHn3b+svC3AmdLB6qr6CYtEX8u/q6
M9AcWgXT+9mxGyM+jnyw+OPo4qhQTHtWHtxFc+xmYCjLcRh4b445XktXQmUa1JNh
02XHpbhOBckkVNgGKnRCdwwDumAPcpgjDwgnxJRjYXJdYoZ02BjIaWv91/KG+Ypg
Ml8Bwqw0+t7nGasXDlOnG+9K+DS/u1nH0qhHr/UFQz2xw96dPmGEq1nx/IfAGW4K
XfuFJu7LCKYAdBS4B3XTZXyoRjcDM3v+4mkjHCNH4zRGwqUYQU0kjP6vT4YcF6ar
KAO0Zc4fljFzKZuDwZY11Bom3//ZOtrCltb5TqZ1VWamdyVAOs3xgl+uKlRZfeHp
y8Bs+FVIQ21Xl+kINI97CpGGf5GD8lerQKVT8JyQENO9vY1I8WRnVEZ3x0n2qxsL
+Q1xf1UUaa7zgCM/7Ia3SxuakWCzvIe8PdS3WmsN3FOFzI1pv6QqSLoo9lStp1D+
zicgk68lZ3pItx0eWwTH5ikPQQipqv3suDsqVmWjwvSGTm9lKFT6yictLspVKFB6
IO35ADO9HFpHM57P7cWAwBQslsBWuwhz+U9U83XGQug1yLegGtpCx3ugrarfizpB
VUTNiutYXddY31ND+pfhYQAsESvxvcL2fEOFF0Jd+ka/DcShJR6D1qli4BAQ5FVl
9IPX3GVOCJxlNGM9jJqvoIg7OydZZytamMzfz7Rp4wkZ6D+jOS1S0Cbgxa4PbM/B
KEnGxIfSz9oZ3Bqe9GNqfKd8fhpPbZuXNjGWpgKfGPe357RhP+Z68DL+GIQV2vIp
Egw53khrBb0d4GYtyCUT5UzdEU7+42lBF4d35GfVEcdvAKx3066ilZKTEc/hGKn1
EDE0HxPDxDMIaiZfrx2i5VvmKqqRVeQ37mzDgjvDLcnxu1+xsTUgrPe7NhzhK95w
Yy3iXiicpjjwLo3KCSTvn94k9uTbY7PClXFsLDLZRrSg3NJIClMWvFy2AhQqx9zJ
eTxNNxRWlsqIctwCrLIo1A3tlOnxdAaK2Fe4UxVqctU/RJCxvThWF/tgbF3R7lL9
jkRPbGvZI8TBfSXAf3aqtFMF/n+t/A9NTwwJmbJQ8mfcEUNXRF20rTOViHabR+wi
gpDF/fh7K64MLFpJ23LtMRxRBU9Mv7vSQ0wh3UejGRTsfibxoyhKvy5JsO4KtfTI
JmZkPmEIGPw3r11IY3B7dVMk4RNmyE9kWdgBL9YlcGDMlXRSnNCf7bzgEHKgvwyh
UrQIPKuYNy4WDHBN5xdihcwMZPD84MUV3QStfFKNWeZg0BRkc1hq4RQfKfKYR4gy
o+mIU+v0wKQYD/qREXEdFwWQY3vl7T4q/ZU8sOxPVgjxCO9RGhgt1vD8KgWg7tTH
N6grsEQG2cYVsqmtBLM52LK4E0olr1IojzH0gDlFq4Ei7GmDSRq2tJ/5TyMYH1dN
daFx8iF5CDydunMhsp9lpT90wRRhYzqRxSO5HiEBGIWj+yt7Arl0hceMRqkg5SsC
NrqtrXQCjvMINUcPfIBNW+fL8AL4Gc60/v+s7ztA+NeOIA7s7Z+mC4MTfluY59kr
KC+UJ/6Y/PUMqpv+q7UNJ7eyzANyYQa61Ioy7c2PYUqnT5Aa0MH/G81sezgJszpG
zKSApX5r7Tas9HZ6wQq9msHeGOoAxYhGNJzoTmYCOWPVdlbKPpXoR3c/WcJ7+EDF
qXHU2uRtkhVzOLVrLJows31mhlZKEWDh/RKlkANQqvzntcegfnHzUqEeziwwHuUg
F4t6in/HZGVl3gTPCS2rzIZvlOqdGzePG+ZVbCTfrNos3Fg2YWgRMtB8WIQWm2a1
W9r8soC0nPp/qAKrSCileEWm6MNwj+mfc+L43eOLTYd0mzVkEpQ7eX7+nslmxQvY
/BdikOooaFNaSjrxtdxXa+7Q84YQ19jVU+UelKMASL/0blHthL2inPAY//1biYLr
DSI3ZA2IJlha047q5ztTPS89ZopGydsQTCERDqCeZIfpLry1mPg1NC2WLxsRUPf4
A8dtfj7Q0NTLBDAdjmaPxyiZkzkE9GxjRLYtn7h5F1MB7qJM6pXkfjvZ2gNIWyH3
8CmkZ4XBDxgVd5Qn7ZoEFbl568G/JJmZVkkDtFMIqk+Btry5fZp5Jw1BoIpea88i
dBwp6yxUjRVz0hrz+zaI+l6nroPkQZAGeX0+kB0FxeQfnkARcu9XMJT+PRBmtQ24
+XhA5SEfduaj93Gq8smUq8oqBHwAsqDL9knaeABDhbAVJ2i+XWN6Its5wuzjfm2s
jHAATMldxwFSnAUmk4kOe2hcPeyQBaTztKtkPcZiH5Ng3MZHMPIYyNh7jWfivJw3
n3P2TCLpCuX9+hC0RrIpGVcMknw8la/Y6SL9LCOYM0bPrzoGFT+izjYENLHYQNW1
ZPu392lhjCRiokA5Z6w4asGlKC5DuxXqQypy75iXZ5sYIuGorimiu1svDgFGU6JU
aI219mVIlLxlvnSjeJ7jwmj+iSeDGRdGE+g6frUcsTgkdD6BTS0tyIsunr/R0jmm
U/SzZ8PDwQPD27o32UCqg9pHeb+eIhXbHlkenH1O+GWadZeORm2uil4I+/2qMyvp
badfu43D2jE8nMoFKaiXZiNyWXOvb7QWdkk2UlH4aHGvaZLJ5WlHHcsqJFb+Gb6a
bMpD7exKacbAk4YzBA3U2P0VHKfQ6YfnaLYNHahicEZbvVVpCPy/inmaoF7Of1P6
UhJYyAfO5mt5Hxgq5gsF93xIzTf/IV9sa2YokH27fT0/ZNlbAUp59Zjlx2H1hDNh
EVcOL/wyYaGpa+xmY0Uf0ZONrSHtKsZ5sy0Yz+9BVIZBwmQRvFLD26T0yrAjWNPs
GhHPeDM2HLAienV596Fc0fxW6HtdTu7qPMQP8JvEaQq0O0uhAM2M+foKSFDYy7VC
8KEXptdq7W7wafuZV2NFwf86ChKDWv5UeALHvw6vQxN2YYbXUuyHaywWZZ6WsZhH
PedA2s3OP9m8MBvMB4EB/1kyiltAum5kxLcn7c+6eiYEHVdTFux1ClUmkjIJVs7x
Rj1Y8rD4CKoGqoQkWd4dp/6YaR37TiIkFa119rgUtGpE8wkh/GwdCpKlnIw6KLbd
I+D1tN5mlTriJuHfgv1uvTbK2CbAxknJZvIBhX0v52Yj5QHY7vYawAImqhm2wB0r
0hjDrc8Xy9yMrpkGg+0tYsmPjKk1rbg5Jm5DyGSrTFdXydVbSrjSGpuEC6LPkkF8
Ht0gTh8O2mK0/f5K96E4GiFFKHQfePhCmJ5N4BG9SGbcm8Et9sDuQwepWVwzAEpp
4ySLKW45TQplB4pnF5OFyVqnZI9kpmQvhoHmdwwn7vkyjgkl2hdUX27XbWXsO2VE
gRKcx986ekbhjW4l9Ub1RckznTL0IhxzK52OQ/cU4ztc2pwPy5pNxYDqDsRv+7ao
VTsPpHvA1yN996KYJJh7Q6H93KjMoPd+UWaITMfte8+x5k+lHYsl0hWTdCaiL8A5
h1YBfMd4aEULEJ6ubX17ICuJDdKMHLZ9+/hTJ2qrcm9Cp7fCuen037aVJRY791dM
zSzZN7gpAlCN7+MDwai9t1vpoWAL+Kg7YkXJAIbBYWFHRRNAyJkVoJiZyPYDwJTR
ozChR1ItFez/gTGlUaTWhTClUNRe3P2PePKP8g0MrGpdRO1Jdf6skSwIFFSZx2Mw
s+2ESZvicv7wHZHWIi46tEcOaDXvX/3Jjt/HxsvGW24JgdMWwOYQTol9fViWCYMR
qYQzwf3OAElR26B8Bbn2ov2DeE47CCUE1uTmHzqP++HSiMPWtG+xnjY61fQx64kH
UzyPEWi1GMdhZU04Pk2vzMALZpau1t8JQqjv3+uKn16HKsccbD+yz6Ze+cG4D/GI
MFSBs4HAmEVfH8nQ3r522Skkr+PEJHj1EoQeniGVU7aDQQ3asYTAUVCaCveXnX+y
aUIm8tNrNd64g60+10WE5cFOevbZ74IT4ACDw+ljqHIJeCrVtqoOj1+OvzpHyQnY
xZyp4XwGMYQ0buj5G/ez3H4cCviANDaKvkgj3RlBmWlMiKy5VE8MAhIAogTLd9WH
0N8ncZE930FOhPQVF0YolgsUYk9AUJSnMOc5Xb+xMm7PMepC01vaz+MGe5QklQtI
8MtyXt45tXvmj99VP9qTGqIiEfk4tRjCy20Kq7yIp2HKE8/LJU21ulyQ19YmpE5z
tzbzHw33lHOaGMX/Hp1V9VzAeYybC1seHc+0Ub0whYti3dY9ZuuV/ns5TdQOOFiE
nRg3t0pTipk+URtXzU5394hYzWTshWj3vXgYaxPUqgv9F0NzO4ZO2qtAesXyjuAZ
VBpKTwCjT+9ErUrekg6L2cCmdwv0N/dnMTRekx4zuAj4E5bYUYMdyq3t5IGC/V3V
iraN8D2a5Mg7+OfOf/BFcNAkRnWZ3ty8R4lmkyAL/PKyNZg75haxYM52G4ZiQqeg
Z4dZDAA/ourN7Jg9qleFqkboBnrwSoktCerOAPWRGC9Dv3V6pHXax01Sn+arjSNA
KcCsj/1XCuAdFgLIYWk1eyL7n+2vkUIUsB8/ETpqR4df8lYwnyUzDeW7GSvIftTQ
Gnto5zeW7JBiVkIo4rX6PDgCOfoXrSrlksDtpjPWe2e8JLqzCqh9od7Yi6eoJAk6
QrN8COCDRHKrkVNKFnzAQUM4zYl/z4hdDB60gLkIUFfkcws35xHx0LFel2PP6tXD
JItPIRRQly1IFv1PFgT5wom24UwXiLlX0RlwO6JJEBmtzGjnC/CXq2kq6bAjwRBK
BNpokWhiH9HxUHnMStIWwpLIh4JlN3G60LPAoCQRTxxBEkrPF72yOx+NiXNmlksH
HOnJDWNPQpaQcWuT9ZEMNa4CR3HJRhD2fDnnmuqZJ3R1TzQyciG406C7XBOpzIDI
tuz9MSTdFHuLII1eh9nXjQTnAzrYtxQaMNoowtvK8kgRu0EtiTXgPX7OQjnLyDTE
T9EFEUdIHKh64UOttSwEM0QOrplacuL+wBQ+kRfEVwPwXbqLBekctybNFpGJbqTZ
Adiu0mb8gr1ttphyVB29q6LyhKSusuL+g/dLPTEWW6cP2tDxAW0yC0XI73kx/1he
AwJ0B7X6Dun7/U/qbfoRKrDQNIfb4glQgNeXwLdS8KBBdCFZPx1G+ULFdhjjY+ju
z4V9A/RuVffnIaCbPU7hc8W8s4H2kY7IssFUdd2xhBlTtonTXXfwl5MrGB7H73Dd
gPgEpAQJQ8+KITZKK0Ho5qjezKhTLcyyWwqod5Gb338qhJSLqCdVDOZWu3VRTGNv
7knjrEmmr/gRZHEXuSPPN9heeshWWx09VX4hNc6eMtpxDmlgzNA/9RUq4taLxA8m
AF6BqxzeKTbts6lQWsR81kD9sGXrjQ+evxPDQ9/in5TpaHhBB1zkSEXJAqjz2e6J
g90r7LRTz4mpIKW144HEfAsNpO5+1/zPRx2SGwG22/iGvgok2c4cTl0N7HKBnTED
V61qHj0y8b1tuwl9W5mvVPkWPLjkhOGO/9+q6RUebcbTpRl3U3lHfFDqo5Fyy3Uh
tMZrda6qgF0Sc37AAx9eyZ8kAIaFCs4MpwYqmGttmb7LmYeJ0Llelp2sjHkq4Kgs
QjsG+bBxZccLEaugW3EkB+PWoBu1nnxoyuTJ87wtzGbiiCtJLMoHA6e28QPtih0r
dNjFCymAR5BTI8lVLcTd50L8zh0ElMZmNbqqbh4FTR2usrMtx4TH6zqqcjAgchIC
8ISUDkS7jFWer8pyGDF3t3cl1d2m5/jCCYSpHDdG45r20xlolJ9VYMJenZRfHOq1
796gf+kPQYsJG92uMjNlg3scNIKofSiiY1VhfabEQGWuh5EcQchiKLtBviMomb5j
CPCnlfAeRm+UzcRzU/7LX5jB4PcHMDRF6Wc8jetqz1C/8AeYFVI/BJXFu1heVEjY
yi+owTeLWXKd4lhMIWiluJHPvDFDBnaQ+b+RTQwExm2yag62Kw14SBIDhNdyfqWQ
UlNiqGab/VAfWJVA8KNd0zx+vC9MVjQKJsFFWBuUdgXn3nCJAUi6Ox6xNOI6dU7W
S/H3XyTeUxgNLfU6MZX10H/mHrc7rcS1ADjT1pgbJd2SwenlvHGa3wrSMV0STzwK
uVRM6IWxRZGaqg4vnMQ52La4JMl8l7Cc3PZhxg2KDaUycknzbGyjQ7BXuzzD+vZk
K+oOHpZJGHI1AFJhUTFl4JPQD0lRHA7+stAq1qlH6FZqw+Sqa1BO+CQDdwN2Yphk
P+SEnZ3HO+9T5KU925U1OvoS9OHMolL0iaiWSr/CZLzpVssEeQ9VHmGcJrcrfg9l
H4Pj5ez/tgQXIm1PTRBrB0ode9JkZUq7pFFd3nIpcsLrRs0LkZGKadxzgVKLJ50q
09QJVmoy9OdPaIPCQV3nwsYdDdYKXZ4X2bmPzgDc/S1TVdXd118rfUtKoyz4w6od
X2UjJIIxh3JB3rDgbIt+jU6vmSaQ3eVa4suAt9lCMExZ1AIIdIzAsgRxcf9/7xNv
eG61huH2/IsrLifDJfHIGYQVa1m77ZivhCpsa6ZgrTGvm+ovxQeJCga+dZQg5T0+
QAUjPwXMRW3NDGnDAlb4PZWOua7WL68dKn1uyulytIurUeDToeausT7f4Yf2OtOA
JIkKvqjWLQcBDiO+oPtIBKp8dtp9i5jQcae6e43h9peLr+8y/mX8reYTSWjw4Ob6
eD+yQttin4MldnT/DSDDqQGcxG0CNynIFEahiAILhO56jqu3aNrBmTw2Y3/GFEkr
UtvzqDmSelp3LlgioEQkEeiEsSkTdYtCSONqy46NFzLMBU2erPvU3Flh1HdZBnZz
/tMtZxyRAWK0Npnpp6QEPycGqindMwoje1AiDTYFl+k7Boo3Oe3JbreX5FCKeb8e
`protect END_PROTECTED
