`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zqJb56vjj4k4euC/Hs6+bc4VIF2kukPaC80EvERedcq4RiAhx0JJs5tcj04C0J/Z
3N9WDZ5tpenctXmCySCtvmdeVO0BLuxad4/LsFoR2GIrEUWwYfAzOPcJeEh8E1W4
Swxt17XcXUow6agaIX+3M+xK57r3cAOENHfIRJitUljjE6oJvF4rCl36TxOoKRHs
DTz9QUjsXER3NXgypAhrE0dPy8HFKx5TQBzFWNpjA49DaZniSzoBrLvYzUZcgHVt
B3IkGLs9feVLQxa0J1Qa6tQDuBaWiwDoTC9eHm+goxdTn+LqwZSOb87w1oVuH9+X
PGcGIcV1nWDgBAsGMCLSeZCaiMha09qml2nIq65L+lXwDnFZJLcXsf6rDkMD4uZJ
o+/DLOA9qdEUYUkWLfgVsTjPxGoaQYhhzE6t8WIvZdtpMvIU8fdCNCzkd4QAVQzE
1YXLEF+bAcTQZl2W/3KfxDlB7sCWs684ix2KkZ6oVz9Exrh/ga7gJ7AuyXGAG55n
a+/mLSS0SUE7pkbantoMGJVOGF57TGFltHO/bQ9C9Ajv/dpVhvzH6JJM9l5QSmEL
`protect END_PROTECTED
