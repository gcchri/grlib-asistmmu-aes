`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1JHu9dvDlJvwVz9pm0XFr92fwpQj9lZFzydMQGc4fHc4VWA+xbzqQl8UP/PRx6+v
1WgtQQ14+jZuH5KIhjdiCyEUPo+ENScP9x/+Od8A8mFTA9Nwqgj+DxUf8DFDsnEP
1VZzXXFWp3va5RxhgUd2N2BtrnnU8bq3eMiaafoUTlVjXtPUKo6kryMU/+b/411H
GGMyTeSG3pF8/Ev2fLCNQxOm972r710godggEjeRoFM4gsHoNSOuxrRQuscvWcy8
QlpJz1MUvYudg55Hz69LOTfZDUgyFfXLQHWJ4/BOFcj+GuHdmf+FtavHlnEG5dJB
SvYVZ+OIz0O/zVXUgX4qlOolEJXhLVeggfoLxwbFdrjpGwUAr2HBOB2nFOKW1ItO
dN/fn34/KK9N087No7SS/FNuZyS+W5adf/p8bE4QBrBqUhpF9DQ3MDbmTn5s4srg
MAaGjeFd0TscYAG42JusLbQ3Wsa7yrmwrxz7GgjBcMa4C4fu/N/XzXtn94/pSZsB
Lnvi+pJIumhl3yZmLdy2U0uKW4r7GMblmjFGpYzcdH18MYALceD41blSYzTUxm4X
5/ttPyA8yH/QC0+tuwLp/RngH1qghZoWFOqpK5yJ6ECVRU4v4e5vfKngWj7H+Dr7
iTnVmZunPOFzItewqexdYMPN34zFyjTfqpnFVTRkoVIQBVG+yZmOK5KVWnVj8zkI
Qgk9RiOM17px2iebC4evioniRmJ7hI2cDj7Sr+hl6uocp6LwitIU92Wgw3RyC0fV
IVsSI8CFV56DtxIbEmYqhc/q/AYFBcUYFb5/7dSxIR9R1B5jrP0t9GObn2yZwm47
dedQ3MXv0pTukioNd3VRqmpvhhKISZh4z61hISzP9iG4/IKQUaV0AJtWKHGdBIz7
IQQqxyBYxAoPmYWBc06PZQevRonVs83bbHF/TvmbimJphrugpWF9bYwGb87ZXrev
A0tWuPta0rA+c4EgkuCPalZzSOnkr1U/cOXyTpXwHlc4nZwBuZ3M8ja9Pvwr2fTQ
8PqTkBR1EQ6eosKG/HpHg7YeY3cwMka6GSEZ2fUCIMV0QWzCvBPaNGPtk3JvJq1h
/xP+PrQ/aoHLcfuAPdkxLYjEP/kflpQXp43PaeANmkX4PzaUfF8liuhhgWx35Cgb
vKOGIolncpdivYW+LzS+97c9GWQVnSrsR2bFttYZoWy50MltJ02nVtndDfmyB5YY
EMaEBi5bDhqjvq521iRgQABTA+5rp3Hme3JSpQ6gDJg6S3vKFe/kgqD7IWdLVxIT
X/beVKf5YoGn2vCR/sma2oOUsQoMq/cUJAYarpyPtHaulRm1e1eaFfT/hoxjhYY2
i8XOZmUIqJyE1DqBAzNEky8vBJke2O8OWQQG8BhYGrvQPzdnvPITcJ4A0gcWdFxv
ifebaR02q6jUEMcCvkyhxk/v9aH80okYs1fWurhqrBXwMqdy5a/oLFE4Q5Vf1Ww1
jbZ9WXapkyoyba9zk7uuVwC57HbLs+b9XNuUGtapGtgf/W+uy2GMoJ2OWk3LNKEo
pDEXYv2eCe6BEyK8Nxq34ugf9IPMe5LqmC9AyKzThojeeLF1YdPust4cdUgv/fxi
5doraEmSV8FbbPKEpxKBr/BJ7cP4qmgI46QPEsPih96WA+Mpj5KJczAR9fdUBjKF
GkC2vqRlZLffCZkafEmh0g==
`protect END_PROTECTED
