`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GzZ3AVG3Jdz6iOKZnc1Pn3QcR11qLXe1nVcslC33h4WPleyaHpY5eqFDUpLSm/WX
h+UBj3YNQAivLUO7U7UXl724umpvpyYibNzDdTDkqYH+4W0XwfKvxCbxJeSunov6
PBGCmXGM7tt+5vjYOYyZL/hCbi1rYmbL03NRchKSwXbkxyWGxUjt2siElDSlb4Fz
pgPEe1xsAei03QIqELaiPTOxewolvt5cJQH9sV3uXAvjV6/Uh7eJqMNjqtvSYShZ
7SNmvvm7MBXte5l1M/pr+isO1ueJchjxrmTiUO3z7uDYFhD3z2EtxJ9In03sRDF/
5ZkX+25upCuV58O82myu/i5lufrbrDf4OvUZ3ssOqADxwB2KvJk6t/J6ZQHu0Cf9
//c/4fl/mFJimsISqBxfGHnpAR5lWnkeVDbUgHhLSh0=
`protect END_PROTECTED
