`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8HIXrHNovs0VbSmwlUsnjU5sHURfZp5dSG8mIDjbbb9TbExvEwX3cgojhFmxBc2k
NRUNmKM6jL8EKqfHysz89r4dK4YbHMinUMDPQQgyN/q9qKPmT0wSTQCrrsGJwemW
d4ugINkGZubFbNJ4YOOZI1XslZcvbkuF3a69H1iLd1YoXlXhdpYXz/76zZRo6yOZ
lknOQuV7gjlrMQdmMwp1N8EXpPLekXIef/YcXGdEddJzlGppyesEpQK1dI2wOQ4a
`protect END_PROTECTED
