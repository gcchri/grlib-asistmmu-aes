`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4dlWeeYoA7NEza5wds7OmAlwUkjJeFBrICvFT5d7k8GQ4Rsz6Yd6JLHAzylXSUEn
EOVlCNMvdYvcDbk+tKwFYAWE/c2iJru5/cxk+TXYpLt3gD8fN817LhoXsvgkI1kq
L1q+eV4IuGx1J47rhKQaKczrX1iY08gDdZeOsdBd/oogZrDlfm3vHFFjIHpg0MOT
BiyWhhQUSFBygVArnWIxiXLON4dXuVvZfGEbY+n4QjX8qjljyrcn1UrdvkRX72Q2
zw1AOAYg/f9yON05jZZMQIVgm91EG7oXMZxwHUghCsuYK+fE/EAmJ+eMzNLUHpG9
q3czBTQzKiIfHsQAJvHc7NpTkmoaRRPxw2rxlKeWoGLIE3fruzh8kztjcpLU2jha
`protect END_PROTECTED
