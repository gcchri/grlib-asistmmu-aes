`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JZXph3/utX7zfDqrsrOxE1eOaiC3BD+ZhcXurilJ8OSRl/AtGxi8064KdC8ToWzc
6qP/md8VYjQePzYx3i7sFz4v/cbz0VeKbLh3eCtxaUlSuYsLH//74UI/8iQNoxPM
QhbxcnXQvW45m2tMfKr4XVH+Tgsl2NSt24nlJ/l76eq29cBRP+TFF8zsZ4tnttkG
pT83t/iKqaHlnSyP4QUxMubQNJgu9th/NZ1SrTSKZxjTnO8Qqbf2bxj4OIr7riP0
lFNiPIVG7/28e47RT8PvR/8hoUoWnXfSN7XonEwTYXk9+KZKN/HrzC0ri8v7Yhyp
WoL1FSJEmk/bnpXK7trKH10PYCnlBy6nfakQqTvh0KWAQOBYGNWhnUkoOTivQ7Hl
RFogXdx+Xzn8Vcd9NUYBagoAVItGOjjQcpQredY6+GPhvb899LiSVkh7hV3rUbHU
V0XvV1UKymW/neU8plc2FdpuLA6I9l6F1g10QQxikNDoTH85Q9jS3nWzdm/4oVIs
fd3/QSXw7pAuSDiDUg/aFgZl8nsl3qB5uIFSIQ4SvkdmQDTs644dRvUVweUcwLwZ
1qTH6SkQynkxr3MFaE6mpyoi+m0tfUeEwyKN0kfFKPKHbROI2tXhW4RsZ5+byCNE
cDRiOJAiZ6qWDeL3Gw1B8c4zjqwe5+nJ4Yz5f1VUC5jfeysUIPHM8HxPVbpXCmw5
7QIcNh++pOo50W0nVR4Ra/GrRsHaYCWT+BfjQSADAPosUF5QCVMc7dZeYuxyz9OL
2EPY4Y/UFfowvVIN7DD3wzIihoLsN8cpNyZFLmP5CJxnnmHxcoc5ophqkiYn1qja
owkwXlPDcM14BJfvrmaxYvmHzDXVIl6c2KsFJdInvx+UrbTiYVPFehaIrzR4NwG3
NX55QZLGpDNYkYjesvxHF8VWNNJI/KUlJIBRdWAtaI+pE70ek6ZPPp8VsO16EfmX
7lBRKr3FTm2cXSQFy8IRwY+/idvmXF/tL7x9+YSYKANYQBC9O0U7Xno6qjOr7u0Z
KivfxbZhMFTo2myqeNMYY0ZObxY8ajwuldLTb4e4lhxmNHKK1QTSjPk+hSiX/yoA
xOU8AlZh4YL5mcgvLTSoixPFB4aaKHT5MioBPeT0xmz6J8KXQi3H8wqS6/dBQnpV
hvwW0lyQx/YIPFmie1A3IQgb153IVbVXtKFTnCjsFKr9a6dzewx6g9x/ODDH/gX9
H5mni8R+JS76Jw/VNcJLbJfWU0Ehp5BdUa13PyULkWSOlH1GvrlT+g/hxjXCCbab
6Wpop5buRaxz3ZrlV8SC/EYDBiL6NpvIbHm6cy3CCb/74y7QIa1+kB9TDEeHazeA
ya4bvKbefkf3VQLhE3k1XzO55idf+9rJSl/jl3o5B3x4Hv/I0sOHTcRxS2zWaD6z
bG6zcUAVGeWNceoUj+TJmnJHaPizc0JNLDRl8WKH3f8m3lz+U0SIOs6vQ3n8E6Xy
SesJYZtXA/IOSbk8QX9uwWIkSK27ILGJxfYfDBl6kDQ5PNfwJHa1rNuqvN8SbUhe
1Y1iC3LzXNfTtjspiHpYzYHE86UrROVisesWwFr9bHYFoAimQRwI9gnLkxyqMJ8Q
unCC9r8U3WdK3ZtPrK8v2PcwRKcPV4/H/vA7zwaLHvevx8YThMo2qKhIcrk6++rP
Kh9PvkuXtBvw6idjOUk4TWTxPRjq4hckPoqzOpB3RmDxdqWZvkhexrGkD1aIQuvq
Tue7NNQ7mc2/Bv82c+OcahvWj8OkgfvbgAg3LErsL3WMg+/AYZzOEuFsX8AOGpv0
F5APl/Mozch8Wmg3ADbJMeP8OsiXUxf+xKht2/d7eGyVqVHdCXvW9KDY7nKLHXSz
QxpT8SfAhDJ9Rj4442OkbYXI7H4KtW1gyPwGKRTNJLb8r6WgVjjf20g/DyNYmgTV
fp/A36IDMdA9YTn+hDqOROMPN66fO0sR04HQQdFGH6X3qoRQtuexrMqAtKmJb4g3
D2ormDo4BmteLOaw/YuMEBApNeeC1B7fIXccCkLPG5Hy5ktKK9BWSKCZKUKPLIDh
5qaHEzOAn/yOdGoo92fprrSgYZNQ82EhxeJsXTEURaxRYHhaYY/jo9N7iVq8TUbb
OSbvbVp/oWzls4nGffWcg32u+6a31sC+3ol922AS5fM=
`protect END_PROTECTED
