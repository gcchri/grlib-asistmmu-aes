`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vhcjFKNQ5f867EaF311An1Jt65OkAojqX8fLJqQ/FxA1LPKRC2tmAVAHPjuRYVBn
xfIImyb8uKooWFeWVt5kHF3NMNFKwM2zvZLbGu5N6gJKZoUTdXjaW7PlD9TNObon
iQKYlFTTtNtX2NlwAH5y42avareltHOjg2BN99nUN5Lfqkd9zx0nmoRCiWrl90v5
r28PUfzAsa01GkBqzbVf39+nXRP85Qn2bVx5pAQEiVX/8uW4/ge/p0/WLugEqpea
y4UB0B0Ukw8O9OK1zlKGbyU8m1OKu1JXEkFM6qYA8HoLY+XnYNSO6CwiVw6mcxKc
KzLsTNyV/okJG10PJ3EzH6ddd4eDhDb+xZ6Z6TNbBwcwnQz3EHXcVoS9CnFIMVzQ
pMAnsqzo8bFix929QROEJwb2mzpvW9oEIaflTxvygnOwTGoN+ncXZLvQAEng5xKJ
WWR1VajGedaz13Nm1RJN9w6XAyD++EYpqDohibk6ldw=
`protect END_PROTECTED
