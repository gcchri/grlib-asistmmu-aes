`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mNfHdJI8NnBFHWj4zpVb+/XVOsVEUdlG4ypkObe98uJQ+h2SYe10ebc4v8/MMdlQ
s8q4HVclTVJ4zr9tYD7jibpAJTEjTf+6NgoSodXLyK8+fy3QDN1yjH2J6r03IP2z
CET1LFwY6S4GdMcnjOC0TSX+KZWwsSEy28weJmwBbs4L7uEuWRyACx5DSXv8Nd77
OzJymMxGR9deiz8kLo/6jXygwlA5o2bX2oQlggvfSULm4JGrCSr6PmJnV+ph5WoT
tIFq97a12TSmKH4Bq7zh3T/LGw7vvSIAsTG2hlYDD+MRKdNFU1cod8oT77rEs32z
M/NfngrTxGJ9oUcNZoGuhkQDi2BZBLsKM2xlmEF5Imhh763JkWr2MPbbEQUFg4oY
D9CpqxfgKmNrjGyg+FuybA==
`protect END_PROTECTED
