`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MebYwAiyy2X8vmtOH1Eu6BTyurOSrLBWidrfIzWx/ZPOL2J529egnpxwqywPLGMW
2NVvDyQ3B4WArJnp+tavt2rWxcmg3K1vb2cftjmxefFEfjwjc/2kCHjbAoS9MbAH
yZCyWjh9qcH6YVrp76wTdOGGr3vy2qX6KhprXWcuvEYE7UWGrEG7vobwkg6n3Y2E
fi5zbiAgsfHtcVymE29NbjWZiYJmkHDEOmN9RO1C4vME0/9SvAU8GMFjFwWuBS4h
aGayHDcUm6vXaiXIRfid/k4ANoh36VXTWbvhxdykdE1SCPKqxJzwdbd44IG5H67q
v65DZRH9SFgH9KisZfMD8eYH3pGyNjJ55kzU1H9McA0O0UT9NLeBVB3BjN4iTGkW
fZNqse/jwlfB5HdwmiU2TS/Xei2v83b7cDVWic3aj+YCDcOR3j571mgegRg31zM3
nEXwXlTUC7PkYCkio3nDwo8l6E3/baoKUdREkrdREFjtfvXj28l458ZCpnBe04WW
fDtNOFZQuCdcmvTw2tW8Yfqp8YflquY3ulIWJ1gHGs6QlsSUu5LwTqxQNNAmjIvN
teFDlvIjla1b0jyoORn3vK6dzIcDm1L+SU2xEPWXidZfr3WU933c+lDEcueOFOs2
Rwhc5U39wTWi25k2I321+NIOVz5tFk8tCL+aru+lb4ly94yzqdGpPGiaDgTaTEF3
6xyzWF6NaRZ1il59eZ8LRnYZVSxMvjCG36T/2h4FuVK7M4LqeoDfRft3mC8RCgZs
ZrldTSMz8GXWE9y0MJwVJAtmu0fuZDtDNkGc5hQa4XGWNInLxwcTV9ykpgUiysao
yyqCtK/2NH7XOyPXeLf1mA76xZb1w6oNkQx+FIs4qgD5JsFXfHSGKgh+v5yLrdwi
PII6k6kIzicYd92n5KZaj9hbge8VgLDjUPLyaJiRhm4dHK2qlyp4WpnV3QsgbSjw
JN+mIqpjAkmCiFdPsscHww==
`protect END_PROTECTED
