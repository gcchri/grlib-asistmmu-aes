`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZvUuWiKN9C6mSa1x+pt3Jws/U7ckFpvfLjd0tnSOqDIuoOGM55tZYl2lp+Na0at7
RJEuQ+j2CjfGmaoIHboEuYdF9Rllk3lJct5ns10Bp0ktxHNuWePWcL/2bQjbijPT
tmaQADf9ypcVI8eZ0sfCPA4Uynn2o15smpAyRdqG3rwnNCTeWJVBwJv2hX5GvpR1
hu/no8Nr2dc189T4QleHq05jH+eXFMxK+CZxE+uuve140bMcZGprPzGzO4bdQd8c
ybHgwxRGa2aPiNK6+6pgJQ==
`protect END_PROTECTED
