`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hNvQBDOnCz/3wpnikl4vODaT0gADIpXsrohug20Y6r4feHEGkFfDRyNOC7P4M+xr
wMOGLmoaDzLXlWB8KHCZ0p/mhMjrGNR6RPcL98skxVCnaxyoYI0SdtaKdyYtQVOA
0qkfqU3kJOxGB4bi5SnfPp2okh6XeXkceuOKt1AByxy3t9UV1akGWEMaUVg76h/+
XiAhw/dEPpv+zadRZBoKF/L95jmKn9fEkFTthveGTtsB0ZllNs49J3UOW/EUKOfj
PidWnqTrvuxQqWfNgyNjRcW3eQvLxK/J8jXRjKgG01313PgOj+qGwUnWLVowckAH
KTGko36KaYRg5oll4UPj46GFNSzjaOjtH7V4os5ayGcYCxsBImpiG0onGDIctl9Q
B9lFs9Smrv0b/4W4WrS2FajpisPweJW7Vv8+St9xf9J/efAiGw+53PwQpitmZDKw
Ax8U83xNiDuvGWePtc5IRSzUz61fFD6M4UdKeh0YT6k=
`protect END_PROTECTED
