`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UJDPV94YiqqG6wEsJzcvxDXaxu0+9Zp3295yvccsOgRsElnzhMslkdqsk9Rg0faf
VmvPKrhW0CQhAs7Tjzkk+OuIREXc0XOSentOSi+HHHmZohCK0HsMrVZkgk3Y2s+p
PSPMQiPRHVB5sYCAoVGz/+24WMU4YQ9DQwBZE3OBdnEXDVEuzFhJBGanGlxxo7Zb
q/+SxqjG8EXpDaLmJfz12tV694eZ/pjnHmq/PYbDVS3348HCsjxdqOom/M1gg7uD
dSOfIzi7+isn/Ul9X/zJ2uVR7WhwvOmvsa8WWtXc543Mirx1Iz8a2kcugzoVOTf7
9ksLW+LFm5r60AhStzyfP2aOuIt3oxbmWRLuI75rLLTydJnPyzA9PaI4783wCCwX
P8hUpTLWPVN+H96fKIJlPhpwP1hAOWm/SjikOeOhPE47TmmVQOOZcQf1Fmh3F/nw
KHojLbUFCyt6lt5u4BG/vZ2bxBFb17zs8snPAwfx7lGs+yvl6591g9tJDRA02RJh
Xsej/CPXHHfbRgPo/3SXAZdfVSAub3xu0c95+lFXLsJNxJVyC22UyY6dTlUO1IB2
rLYry8PaL45RcCcnZWGRYpr8g374hH0CNPQxvTUg3slbAqTBmJcpFJxXGf3hluLQ
nRZwwy2X0lNEoucN4/IX82sEpMyIfcFXcOBjevHKCthCR5xKxE1V9Jy6BYHzPFfd
sGZhn0C41ziYArHs2Cm16jNY6aFLgb77KPFqp626dlVbTsWY8s44VIPGVMZKVwtp
uImBa03Yoi6E3UKXqxumlhaeF2YUBQuu7hAPDxlnMtzXtRgUjaayt3OY1+YTFy/1
KRFFyNp9bHLNlpPx39otK0PY7k8UJ9HPva/vgtC3V05zVGa34+JkIYjGpbT+QQB0
W2j2YmgbCfpvJIjSh+vDeWQz18cLES7XTeB2+tNptHYWRSWioY6XLJYsRa+hJc/k
ZHIRNd+nctlalaolUYU0kxpu8oeeme8AgVs53n/DdgblZLX6A1SHTe8SlbQBZXpr
QeWm9jVeIDJsCL3hv7KZu2WUk1eY3OW0ZUYQHQMZ67KOwYiTi4+HCg750LrOR1Kj
JGiaNmBNTF3f90AS0bxFviHZCBLxcRRuOWX46xVF86QFmRVZsJw3oGKcmaW8+XXp
g0Pm3pQzI0JP+PFf1ApnNPmQtxLxLrxPCtQPl/Fx92bGBG8wjhxOZOy5ATvbNaxP
XZf2BOc8Pj4sg4WZUJDThckVyILVjVlBUctpePq95zECWYn78ch/49+X3oVfw1PR
hzTbNcYks8WoJ/sP/DQ1SAccJD/AcSdRGqLDlezyacSi2LuaBzd77+az6VvBAQct
hUmqvZgQAiWnjOIhFT0hAiZfpVxWrkdz8RMVwTTBuj2YNyhmpIm3/pkArV6f/oQ+
dodO20OYHPNd+3dstpjGYxW5kGlETrW1mSUkI5QXIqyDleO8bDprHxu7T9QOsiRS
Z3/NhA6+j5jyQgiHuAHUBZIg3vZ3kB+W82+xbbff8V1MmnbS0egxocZsxh7QCsFh
Zk/gE/5hhcnSL46tpoIvNvSy2U4EadINKpmYAnCwl3VGrIrBPIfO89/JjwdDx+DF
Gik8YyAUci4GGQZIsUWjzptiQnDCJM9/JrsUNO2m1VhkRi88w3Bcy9OEZ8ChJx8Z
dAbLF83axLeMpYWxzNtYzAO4Uatw4dW6y2nlUfSnO8jwmuC/g8D9N9JjvJ8JO3V3
2Y7jA1DQuBHBdg1/Va1th8Fx2fatsWM1oymBze3t63NVWC43HrINeCbDmWdgwSAu
n/OWgJdgqiMFHnQPXov+MPGr2CSCDKA0Tv12yxAQolJGjephXWsntl9MWyMWppD4
iaHnzGUTIl/jdpniXjpUECNsDwUyPzJqVl9k6gVUu1/g/tF7prWzv76GpMkCQrSE
DhEBk9Ogm2R+dtIcSiYcpAYu1FC06dKAMcOnA5AETRpQosQ5XYsLS9tyPCLQJOF8
CKfg2HlWChEvdro0chePmx/Ciy+5FGZJQzsjsFVedC/O08VJKv9jNuH/Y/pTSNow
ve6L+q3RAjzQ95lUcC8niq2urqtUTlR9ObgyMmPKCFuyXXhceuImSQV06ltSWUO3
NJFI43PX/j8UskI8VR1Yud6F0DyWFCJt8SvFKAIMW9hBwLQRcf5LFuux8LoRIn7C
2Yp2oJbtxNGTN84t6aQAp8R6qdRQZ8TcQIC3lzBlZBy8Bjud4JoJExNt8ngq2Ddi
bHwDvB9uqDsPg+BoJu7avzbwse3/sM4j5WjrNUMshfvXJkGoZpMz73hBaMWKW6vN
zJdQWV85F4RPESeZ9uRZdw==
`protect END_PROTECTED
