`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m6KiFDczeY53VBfcy4kdbQVJ7ncgRiMi6rkRXIlqBmRIvY9ztZ+DMlo+Daj9bshe
CvFWzXi8iusVMszHGqbX6cn1ONcnJNcG+3LTBuzSV6hoywJRvhNkuDmYdmggfH3w
bshKGCv0x0Mp3FdsV4ixJ4TvZ9AVC9e2gv3y2HQRM7/3KCCPp8NvvEPWaiCLL/DK
D1nbg8D5KkYtrWX+aNXrQnonAwEotoAbF0bNwaCXdOu2GAh5iHY6EMjv4dkIFVei
9iT3IACJQk8h61qhn43Vzog4G0bKXR+d2m9r1VVDjIOb0+qrmwsjOtVSWtjo5uEQ
aKIJE2qBZY52pZa+oRrdaw==
`protect END_PROTECTED
