`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nz29KZRXxjW+gAiWiyi9L4WcLkyl2F4pqk3gjRnHDIZNeXI8UnLJLB+cI4x8qQ7q
1YUvTPXPfCmKhhxjbaKKCL9ZL4XZjpPgg02XpVW3PQIq5sU4xvFhG/oRHjAuh8ON
jKAtRjXPgDJGetzEgSLsxzox6XLF9NE+16CW3rR4anmGSz1Xxs3I9bWK+49O954t
U9qiMpcCtDeCrn83ZSMb7DT9fcQ0QpF4KWpWFSmfw5s1a+7+cvOlXBZQxSAy0FmP
CMj7k9Bln+cVObN85l1ZnnwVrxrbRSBIFbYl1bFlcnjgzGb4xU3Q3O/C/LFhe2xA
PJ5QiTZBi/rFNSvMS9NYTiz6bJv6SA5pWOugubm8KVMcWhdpR3iCBTReUINevIzt
kyEn9jFkRNxIs01nm2/VRYpNFWLBzFX21mZg1Y+IYIxDJ3XzCM+9fY1/uGPElU+x
1IHr6hFxqj8AOLKmMDhljTeyzpuEVIBdim78CFBM0pkcPl7uvDSe1eYUGREQiLT+
0IZlw6EnBv2A9P3Q+Ull3Y5FMlmSZsEqYEK/P/+6HIckmVwTe+HDpTFoNjlzPaw1
hHTFViSLm/bBg1itzHjfglwJGCg7QaGAHFnVCUO20qnwOJU5msuES77vuu9j8XAf
GpzVVSdqTpzw5xGichm3RtV4M/NzsHinnWTpq9YSiG5Z0nPQYxMtKxdTg99HV5Uj
0JS6etYK/BPc/xefvK5oMkKsXgEfHB91fX6IoNAiZO6cV7FDNPvBjFO3Ytm5QZ4J
tDYcMWdNYFoatXvP0KQd/9IPMU+wqxLiuKWWEu6+dvuRzmDOT7hNhIdtnbOjouXe
9HhllllC7JeC6j68EUHj3g==
`protect END_PROTECTED
