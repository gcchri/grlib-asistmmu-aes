`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XeU6hXcwDDnzuM0PzAE3+DfaybCRrmCunv5iADRoTavYTf0B4/xGhO+QgRBzD+FD
eAZVlZoDtqS+X6y3pPoMWrK0DMygK1XhZuJAHENA2cmRL7yvt9yCO1cnQLn654Rr
iLQfsguVXA78I8BQksjXFKBaUoaiRxAeyM2/RynzE1AnjseCdh69TOz6kMqV46x5
HrDSOdMrZVo/BzJ5EnuespowzYCLMqrJnbrY04znns2lPqVEAVV/DMdMdLIqRUKw
PLGVz741ZmDsYx59Z6wt7WFTT8vLJx32NkGgiEVITONRvhnPu+8vUI7igmAoYa0C
Tc9S7VppThB5s96d82HQSM9Z1TF74V5HQ28AVKfa2bOibovGD6YGPWnsRX7O353v
UVyL0Lh3szPVehgePaqDrD7wHTX/xq0+SzDUxFaA7xkINQ9FG2TSK0FB1YbiOJ9n
U1F9llFMeBZ60OKrIUH/HyZv8MDwEE8KejDgaRnOLldEtJqUcBVMPfk+fDAt+DkC
9HiLzUyR+O5LPXWFrn7T93p39fgLCz/bvNGkbVIuDaDhXANPXFkkVg4b0HEdKqaR
3YBkFRFcjU4rOfbVvWihTbLr4K8S3No+Ob28X//mo5vSP/mmGsj6Uli/0/fIv5Ur
SViWLH3EkayUAo3+4guLDS3XqvDPT/L/PCZ6qYsToz1pqVMQEl6LaoZ8RlTpYeuJ
PtHruT0zkdfzzslNG2ex1FewsfCx3on4MVbZCok12wQ1+sKmtfHmT5PtuQ6kJ6e4
NaQ5gNr/Zy4Vd+8jBc8HhLw+4banXtpC3YJmmh1DwwpBso3RvjFd/5H+cu5tWk1E
8fh8wM5XHgWK6Z+zxa+/H8j1xG0m1E1fBeXUoJO8TR+9y3PZtWRqVXxpuHWP2ysY
4B+2wZHVCB2YSHSgtMkrnveTC7ofxswo7CnrD7hOoK67FK04J7hm6D4hrVsdvrfq
tDMF9JmN+5/nWn0m1AJP3PWwSf1ZyftdEZ+UpUyQaWiaupjLQFHwSMUG7vbcu4Qn
uWAXTP2yCJVG14j7ByZdJHzlRPrq6ycD2RVxk0DNV1A0exNW6avWVx5KPkuzFwKw
zYOf7CzRjj0luIZOwjxxAe+/nq5o1fGfKnTx7m9AF8k4lhpArztkpe3ry73Zb7Ci
UckRRXuuy9pKEjAbe/cko1wHVYQPppLmtPzD+yhUb39C33Pg2NFm2ZqrXKIL3CLk
0KFZ1inlanK6v8mzgzmiBnXKksPR6OWQ3q1O/N0kfBlLOTPF4NqnZt9PwcSL0xAu
UXsh8S+0rPTSoMKX8TypElb/EmVcWC18gRDekK/YmnhSxv+3ynU74QmuBwYryWlh
II2pRgPdwy9AKHgxhOqt9JD2l84TUZVWlL+WIcb5+6fBtL7ndcP8uh0Y48Tg4PPl
IQrSY07cfrzsR824XqX8QYHaTXqpNYwx2ctIqiFyc1QX0Qc/wPhUWnYGBql+JFeE
M+jHKQbBYAmbwaXxe3Vgnj+CpqPUkJ9g+bb8nvnjDif2VCqcY0043s25xfS9nJYA
eIJFaDsSNBjSnqxuiwXwkrmzymMNdT7OGlYT9Fewc4B8Oh24jYLu83iA1YfAHrmo
DcgduY6WOWvVDShZK4H7GJ7/uqnGKfFAaOVaYVZ2YUJxGzE1yOJzSfASPMrK9Sv9
N/kiev2Gbns+o98ZeHaMS6tnQxkuki09LdJx4bCmdhg2w5Guyzbzr8peGC2zT0TX
W9QzN1iMBDJFCkHKdVRJB5gjZpq/qYpyHifW+3nWrRcIC2maL7khqQi814SCpYF2
g9Sgrcfr3WuaZQCE1KXf4k9oRsv71cgNXHoarkhVtKIrSHivzVEKhmH0IqF9iRTw
Yv1BkDGha+YMkcJRAk8EbRy0DckAUNOpdA1YTH4/B6wPeRJUDcNiWTSF4FnJNKj3
YrEm/Ccfkha39lbxezq59xzQY1oaazv1eKYHRWjQI9WCBhYuQUsokU8C2Ssx7kiQ
TqqDl6sr5Rw1P0AcEqZZr4PJcdaxv8RFxWz7dNvi+A8XehNDKAdB8B91ws60gYTF
DMMRdw4dL8IJhtYu85QjMj+M+pCKF0T/x/YR5rGd+2DOVPJ/1Ahyrmraqf013+yV
M4kTrvPos12zcoOcN46Dyy3xVRxWyT68mtb/1q/zAqeiW0OgSfh/52C/GvkAv7ti
Ax0b/mUvaI9c4Z/7fFql8ussBySVgpcx1+YGygkvsIeUM1pPDiB4pKe6PtdTJA+o
GNse4sSqMNxFaaMnoZQiKwqWFGYzUDz4M5bGHzpE7CVtr/GOO/JIsshMLvlwgTyG
YJY8eY3Tcn9iOmc4yvMP9vSysDzhcMan/LsnY60v+1m/uU3cgLrhE49iTN0kOpvt
EBiT8b0EFNBob2WCO9OjkUphh5u/RQ/u+Ns4ok1yYynDCAZUQ/Fr5MR+VSlJOCoQ
z2GjRCsGzNNIfylmYNiqL3d2MWELFcq7HzCFbx/Sf1xl9o/uATeGjMti7f0vag9O
7uq07Y3NHfL+hLGkGdxmTliqXSWSvgKUlLAg6eFIHd0D0U2Vgvc+2+slV9T70H+u
p6Y8I3cfD96WKNfyme5hGg5D1mb9+CKXvTL4SxVmKNLZrbgoANLefJg0Wh56EEj9
9dAC+Z8WNAKhhVuzR2CIcxwbWJ0v6mrbYtS3SlJPiIRS8pJ8SZlfKjnnhSFGQ3W/
cWvw5h50dhHhSKEGFC/pSu3/tWnsfoZERPxIeHURS1ma1IM6MNMM5w2aovlwmgAV
uQh5/muYGtk+uUmDvdVf4uWJP5fu/uVolGo1zLwwU76Uh10tNiQ2GTDpxiYlMcVX
SHzVvvMi5OwSjhW+Rg7p86SxyjTaGwQl4vTx1CWMCihoZaM7aqo4opk6LEWay/OE
E+xYVCphfkO23T2NaGhvciy1sdDnYrNiBCabWtzGUTgvRirPUyQJml8z1wfnuSH3
z4mFDgTDKAxWu/AdGLKT864K9C8te3rRKkc2dnUNcygmuNfXAO0ZMFxGD+bFGn+u
dq7sR1WrfrijPT5Co3UsUGhZ7ZlK5HaDiviMeI68SxmdK2QmRLm5vpAfnjefCASz
PqYNk0A9nDplA+Xbz6iRiDBUQp61Su28hVs/9nWLm3c=
`protect END_PROTECTED
