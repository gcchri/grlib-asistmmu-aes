`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EpSx7XxNFLCLV4+UasAs8I3l1/v9+5dX6MGdmdOxJG06fB4CfzRL2tL3f6it55fe
DYPIzbmSoNuhRrGqNnkzFyL5iMr2YOaKSrpU5Fasd2PANjVZYyBV8Y/mENnHN/U3
xsnJkeMZsp9LByaVXx3RKmHxsKnWtDZ9vgRC8aGyMt+zHwtq9jrXYimFLrde9uK/
YpaQXFSHQtGE1tNX/8E1LnYbkapAP+N7PeM6l/YikN4tIxComhS3q8pdpPKjrrZD
mV9VVCwm8dVOXkvMk3JixNl1bFrSJ17iseMdDZwvw2TPl10gb2GOvgtZd8ulDOkL
/TKKIfaumyy9q158GZf1FZUAT41djU8KIWug7u53HRE69/8YkND2DxIddjgx21Z9
gLHLFgXjcpNTYxA2mXZaRM3YPWnSBnSi/BOtEZ3D4XlBumH0UC/2Oc4a/oR2rH9E
3Odk7czxWK/HamRDEky4tAbfWTF2/yF0dyn10wKxBO8=
`protect END_PROTECTED
