`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0w81VqBs2ObuGYwQueE7UIhdNGrygZfAYvpdt39wyRxF1IBaAQa8vRCEFAi/2pkH
2XNq/+eRyztUfEB/zGp79KBh3L6o1O8S0ZMvaooV9BpaiaeiLun/z1ho3cDGnCji
ZgcnELObJDR4+9vEYfcy4Yi5t7K4fOrVqYfgactLmIrfp9iHoVYteIMiFVEQ1Vmu
kivdzmf/LTR8QDVmrG4g4M+w0umf1LLpclkSRD4tawox9zmakD4Xg1RdLT0YtCQn
QXCYvHPkwDPiKi+tR4ErpNbpb7o0DFo8ZxQX7zS/Fp0BGRXhdVSMPHcIDAJxKCFb
qMWJi6bNmxiFsKpCKfEDam0u2B0jbh0gQsf3HOdwkd4RJQLU95g21M9N1EFWQt0x
7WJ6UxrpWZaktCiWuAjjhtvZ+pygHU4qUZa33bbEug+9R+mGsp7h7pgYtR6GPf2r
PeHlyGtDJVuU4V2n/2SvsLKGdDwEjxSQGwtdGuBbb9zARsVcOE8cZDcMZctE7EHm
KKS4IO5tvv40c1GD5rpMkvy8B26hoEZBD2zKUh7KLpW/xsLNGTBBWFNE6eSZwOR8
KhJOpm+YSMJtD9SCAWfa8674JDbrHUM8EiMlpDyGzCPfJ6RcRufDy0u1hnrSe1yM
tZjwyG8JV3S7t6aUxY8EKl1Mwsii4T3+F4KwRiB07Mc69jHW1wUcPSOraMB8IYfB
IBY7566621jS4+3E4wRnSM37zioDAQTfASgWqALlWmswmMUBJ1Lus6amAugOdHX4
q454Us4De7J+vZmnjpf826I2ckiCU8g5O1/dSK/tiM6EKsodcps27p96yEUk1myJ
`protect END_PROTECTED
