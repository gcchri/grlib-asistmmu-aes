`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DkhBecsL4VG4kckGN0JBxY6Ny8wsLI0pQ6YGuR8A2mQov8bCmZcFMj4nOG1DvWP7
JNyGBBzPiyYgSoWX8Nbzn92FPmDg+LLOwRgYmSIJ2j8u7juHJuxwj60CLOns1QEd
ivbSj2MC8t7yLJqIKR1qZapC/3HcbXzX9dX0lm1gtVBwCRm9/ujpSBvzvmDbeovX
myW7EYOiqFozbtjeMN6J0bjdPJncucS9IZda64w8p0qzvq/yUehuWnZ62OaOcfW6
QEhGoROzG4vHLK1d0Y/Ez/iiYOiC6JzECz3wukV/gU5qaDErO0sX3FR7LlHyCELE
3bwodHlPhOx+/+vCzwTncQEOP764EP4JQPgvAiI6ZO/8Vo7KWxk4myPekVg/Qc3I
mjL5MsIWAJCw0veJE4oJqlgQZovP4FDReL5zQxP9LX8ZF/uN6GD7DlDDMZytVZe1
9G3j21Uq2uXc9skoPOgJ28maEKtl98QHwFsrcQpjgvxGwFnvQJLAJYpBB1fEOnVe
84gzUCglOsqDLR2Vgruxv9NME2VI7E8SgffBqhOhKBP/RDqpR4K5nvumUy+pPTWj
g4DMy4pgW4K1JWZ9ZwDjpg==
`protect END_PROTECTED
