`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S4itsdca8h7GeVXWnWBPBk1yh7geFcP/MhbvU6Pc7KoCy7ofyuKFYmqfrT5EWa7F
TXRXko1aMNN2RZpLeAS4JWe1g2qAcOfxXv1QzDRQK1o3XWxe+oWtbsBl6tuKj4UI
gUxiPx/T5BqQe9+x+obZ+rO9ON+7x/0CRC9P/jAZ8OxsN9SLTfRuDCWb1KibYAsZ
sQ2aFw2/54HWwJWRnBNt7whlWtKt3D4HXSs8AqTwMflMJLXcRWR1ceWPbRYOi4BU
5V/Dg4/5RUa8hvU3uzWAHsA8TGWadtXI6uVrqyMN5Ck6GEdDCSnbjFQVHOHWL8vY
vJtXWBz2yRp4u+DJQhruPwjBFdZ915DBivVEd+IBNhxG6V+77BJcAk0Huese7edg
PpVbweaEBul6e2UXJ3FEaw==
`protect END_PROTECTED
