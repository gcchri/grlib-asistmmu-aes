`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jve8UQlkZCYuqoMiaml0UI5BrQMo8F9i/kIH4bxNmT4c/pny3kg80Fff8F1fNw3T
75IgQq6ePS5TGzu9CrjumIZk45g6hipY0N79DAZVR40ycyYCBYJoAs9pMqT8N4vS
hNeBAXJD6yyx+QuH+ruTCNpDzC/u7JrZo/Te/Hz5nWQSZ8ALqHX1RJ8ws9tosRdG
HRfXmrmlAqLA6mZjQFKr7ORLmht1sOP3gc+oByJhTgAsF8ojYpFL7LxsmEO3F2/t
YsVxdwMa6bpvleCNvjHz9eb3QnEIg9SKSLp8KaaSdCzzrfAM0RlfHEpCeojsNHmm
0tTSq8Szx476tjHrMSY6Z/qYSZG2M8n/f0qSC4sMh9DZZQ7iis+ZuuoMI3RjrPkY
Wo8k8u8+dE/YTMZMAKgVYxYtYva1RXTTHrbDTevDkeY=
`protect END_PROTECTED
