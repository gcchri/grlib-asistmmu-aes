`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zNTYLLpeRCov+pPtUeWinVnzQCz3QRON/LJHY4KVoZGyLr9RdjFeZM3BfhNeM7C/
YHKpy0bIzExcHd/k8wTp/QmOfUOMoU32PBGgL4gT2TrGnvutYWcJoN2HbvCwMrjB
omJ/QJDK3TkhMeiblG7CPOfdnTnUn8LOj1jCL3f2Gt31+Kd2qr+RUIqoYy1n7PcI
b3WajkeWiYxTArzVA9TiAXKxzgeUCy66dhEg3sMXOf1useKWtO13VRymHNk9/Qi5
iUFXK7yuHflslBfCANr6yU+IHJ4MU2xIeDQvd8AnFmqgY7fAyL1l/UKBKbv4pnoO
g9YLsXN+5zusqhuluf6zV4mmPFRv4L9E8eH8FdDk9olCf+tPIJm2URPuQH7sTIqo
i+Clf6kLFZUb47oRC1A+FVG1kF+yjLD2OMS0fQKVVg2gSWGlAsYLjZ9tq6Zs3ngj
FLstTGWBmKEmvx2+PgdHZYPWqB/ePGS3wrSwQhuoTxcgdtFiiDKIv0QH0WkfD6+5
3R4GcgjUesYsfSPcHUFIcCPSRxSzyTEDDRTkZXdhu4tyuCr0wStcinZOWpkg7jeR
R/NUG+89uLhT6OLUH0vNfAXLLaCKD87JxNbCkZBfXo5n3GjDPGH8GM1SU72Jr7/C
Fo8FhnpROOOcg4XoQr8iEOCZV0WabEw7OGQveBymoZE=
`protect END_PROTECTED
