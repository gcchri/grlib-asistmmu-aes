`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0n4hkAO9c9khfAtJVyxbZ+MMfCFL+bYnVaEV4g9TuVjQLH38g54EFmxkNApy09NS
WybCzq98aRbGOEOUpPSnESD8XC/0iEZ1+3qngRu/TNmZSIE7zfth58dF6OluniLB
fvp8qeja4/0Fp1XDkzRXo1NT8eqKydtAT7uugwCjDut0veGlno1WkLSVit2CFSyj
4t4riDhrfFebx8QSkwYTrUry8AELYc2op7we7Ce3g7KLJrxLQmGSV0LlHgXyl5Va
uMs2fG90/4AYWzKWty0A8BWjf2yDZL10zqXWs5NGXpEJT+61gUYFxnQ2OIvWPPwE
3GVH221m8NcukjmUGKNeScwsNqgKGwn3qqxIPSz6DqkE6syNWzG0ldWm1V8979N9
wrIlMnKPxzTNNNSco8rpSg/a9wjxLDHxAKDVMEhAsM/oAl2Z88NArydwKwTfiUXp
6thxCUWagslg5Lr0oKt7tfxDDKveA9+U4tu1lwT1d0x9yK+6sY0DlS7TqJTVVYD+
za4O+gnsSv0GGuOPL24jCjqmMcN+84u1joSBgqbkyqHZoIB61v90m09TS1pIzlm/
Uoqq6koUnjEgSQclJ29qdIyRP8nMapDXZFdQH9CNyGV64t5a9Hid7zfCPdvqZlId
aoGsFDwPKF9K54iJ+vMuaagd9Swpb0ls8ESt6VYyFHOsJtMS5URPVe54mGPeAD07
`protect END_PROTECTED
