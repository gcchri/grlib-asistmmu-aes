`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g2YVZJYDFGUn+fq1NHHLgWsrnZmD8bOKZXkQOxC0RgIgyarfFwC+kzgKMJEUD+kX
4M6OTsArqEQfBRUU57M0RBP1Rr87oKyLHbtsjkdMBBtxvMs6NLhp8CFcpCczuq11
BcqUIQ+uQrkx42MoWQwfhk2PqdgPnFU0jaTnMXVcxztyi2uV/kUDLFV8q8tEXoGC
ucwI/scLLAfR1IZufG8BoZ0ZP3ubhWD9mSbEs9ZxVOpP2tcHEqPaugX/v9XqKSKb
bTSVCOsVRdILPle+5aUF9x27EfLNJdpmlm8ql8/RxwnUBQaBMU3XAxwR+3hOG/xq
nvuU+XKPBpsa1lv2oLbECTSqK+ft4mv+tjPMnnmT1HkWDSJGcHWj02fN/tx27vAK
GCwFne0r/9tfwGWHeSsvHh6rV/qUXED/GHQd6N4kIti2thK1W7PJgjuRfrCcj6bc
ZcDw0bYOCpD4rEzRr1L/QxRCisoolVbCzdcEzrcpW/1OaKpesKeFJKldlc2X1rPn
YpRbA4WzvKWyFkiie7zOvg==
`protect END_PROTECTED
