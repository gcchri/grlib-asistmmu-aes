`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PMyy55c3f4KmgM1HIs3mTmGDNgw/azIzqIZp/THniSNftFe/Vx3BQ1n/gLxz8cjm
mjEGbfyRdGVKVCv6/cMzUbGvvs7ORQxy0lKaF93TJr+D2GuoNcQCmwe82w7lh2fn
n2Lksom5OO2YT9AYxKv3c70xHjO98z9+0wp4K9ycCeKrvDlTE4eTjYO0lxJPh39/
T7NMoUpiKVfHyykU2cHaHz8BrBpvo5CLyiFk4fLuYhx3cEVBlUwApHMHj+XS43TN
GN5LY2bK/aXgVQ487/EkPRxjAQ2kUkfNRw54FBDvKuJ0ZJQW4M4dXz7Af6egMF87
LElJ3EEvAe3oIa48BXtUUhVcqgJmG5Ez72Zmh8EtNtWPl86uKlB5LUh2SMTlYg5a
/OrshnbhMA7mGhxMFA+12/JvJrs3049K/hjlxhQIcdvkRku3s8t7LIf3D/7RJ608
H9xKVLvZRbzFn+vM+dYDMNyVZNkyhco6iUw8A7S27u2NrF7hxSXaeDcuHKCiyJuD
ji6RfmQZn9qXBFuNPX4XveFQ0OehLv3QEp+2ysWm9537FXIuhbdGvOwYPN+MiNhD
BvWPLayrUBVLrlIJiM5yCP+16w36+iBsnlYvLi0nnlXOSh0vH4DKW87KS9/7NOXv
s9IAv5xtlkznDOuDXw8DRLdHqTA2riGUQfOvaDoXYFq3XKJxKVuhQW6xZ2I+ejOX
KOUByswGTxW36J9yk4MboeUV3h0uMAkW5iDYNB3xIp28/apYHOtVTD/b+C8POxJ3
+JJuAZUHCMKLVLwBf2WDOVpc9yHuSwRzSY7saRUP4xC40nhkgaov1dkLUTuHiVai
VHSp3jlOxRFVY8NWrjf5woRmTWcEQPnRtOSjOK8TaFga7vFCTxP5FfMRoSvkxGGq
5v0REZptoa+ACITTTLPmlT5duNAl01zoScadD8vaUj6GdYHIcr4ffGxph/UjC9AK
kz43aNjpXrKxS7NvUwwGfpWvBGKm+lucnXSOa7/1wU2dLUJGnXW12a52bttM7SSh
AuSENdBxkngVzw5qPlQgrEqtl/mxwfakgz7853cnj4fm+UASgHhueFCOwZLI8QGw
Alr4gHu0ZDmCg0MiXQX53Q==
`protect END_PROTECTED
