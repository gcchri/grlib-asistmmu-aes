`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tJN87TlU8Xnic2ExZSxT7UpcqIlp/mGGKNdMl3t/zpX4Kb05XR/si+Tk6ccOkc+r
g/gWc3Ad/Pr60bFmC61DXiTrwIls2BovWkMQwBunEBWzw76wtkpI+l/rRkgFjfVP
wjjoqKdEVUcqZiRh/G8A7QXnYicNm6562PG5uYA03H98sxGEunAtseMeUBLAkbFN
beAgQKl24QSzTmHL2QMQIBXGch8qF6cTCbCaCpIP3WN7K2Nb7e9EuH/VKvWjL1Eh
3axHbxJrYlDXhMnPBYdAJR+wxfQaPWmjN/s7HFp8MQanlG8Usng93e93XYCKxaye
zi5u1F1Bqh26uJTEg/WgMqzO0iLP13Qv7WZ4bOlzCIWaaP83VI//CQEVh0msyDoZ
KS/DeuBkVOGqI21lksEf/QnlN0KPSlkm/AklydayQiwnzNFKQ/KUwfMLxc4i6UJA
7Ksn+41HI00Ygymf4f5AESt0wpO55xps16/8yL7NV1L5OV3Pz88k7PwwkoljDan8
pp1F8usSOU6Ytkm6FLIgm9YxRsl2IBa4FodHx78wZsb9XOs2Wq7SLFHfRjs/hPYC
9xyh0O7k5GDbEcyDHQvBw+bCnnO6qx7wlsXvBwUrYAPMCWkDjVPn0L/ZOZlaBZh7
MQpbaE5+hX4RWHpdmozXw4RCU07vtQwQhkwZrYmI9kA=
`protect END_PROTECTED
