`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rlt5Q9QyhcYXe+FuwN0j3elxRYxy89OLRweF/l+hoO9U4XGdk0GCeOMsWCYQ0+87
cGnyu/I52JEjpbl9uDSIGCTkjy+S2yFV3y1zcJS2MpXwGHNeAgGftIK2u5lvZ8lM
e8qL0m+VCit5+hA8ONAsfnDiyDKL7P1BtW5S4fboCzu8pUlwgR8tnJbnHyZ7GbpG
PY2peb8kEduv+w66xLMnxSq7WI9g23zlEVKU54ZmbYH7Y2yc2c9Ins+lTLlhhqjD
RR5CJl/gBD/7iBo+ZMpgcSXwgV+J8HkPnTLWf8FZnq4rgehqiqqZtCFvYNEmp96C
SIpvTvyFXf+D0WzhzTii5XaJ94p1cNasA6KVdUwICe1uW2IttdmlDRgQyJmTAquU
FIvCbkA3YIpPcvfZFd1BufL1JY1hpRDMN+fSLobbZRyaVUvRkfnCdG0R3qcHZmjK
JIXFnVQ4KyuHBN5IJAIF2lhgtHrh3Ve8KSxakbfaFkVpQ0bsFZIyiYWfh8utyqLj
jHinP8QuJmjzZqlAOLQ0HYePLBnvRiLo72z7fk42wyWcgkWkudlM1YY8Ot6AX7qy
8zooYxhIhN2zUdttYBghnqDiGwcQ0cCD0dXBCEAHgVC9e1mlIGK8OQGN088aiC8r
wr/+Fw4pCBybncYubDHG9PksZ40ptECqUtCFJ7EvbWM5g3gLNsYD2j/XdlGV7Gwf
hrbTHHXwNsxkHiGk5Cg5Chw9TTU55voL428SsLcy0iMfpatT7RinJf5wWcSXFAHZ
LWWJobdleL8UwEOT/6t49eKCTCWSoDormaKfrWQn65TQixq3fK9FudtSOA75Cy1/
FqFnk+rRR2g8YsrbbApnPF1ER+4uRx8tQCEpmUg6uVGNsQPNdSKLis2Ijkcd3cr7
Tam/vHgWLfM6o6qVE/2u2h4zZXKr0QQDE/5TzvRPlqkaLa6DEIunLYhNEcRQpaSS
Fb2vCgGroUZHn+DscJ9pMXWfokXKEmHHHkkDTYFc+g8JWq5e2oPAwl+EKgkQC9xy
1oWjDs5BbYf5xWXGNq9UQr7oVOgPpb0A6+OE/Ud0B4uC0DazoAm/GKBRdqChhrTS
MWReGwGxWPy/pEhMPVat4JorlbQabpXI0uJKc+5jq09dbXKkmZBOmMcKcN5ak2zY
gvyaDmRHGXzqy0J3iSZIQyspZLb5Gl8D26MFM5WDhJYE7ebCymooF6mXe84IEnCw
VwKwQlFaRVkZenwI83JfOvPPqcD61+u8yPrQ/Dh6Ol9XpTJ57cd6Snucbov9oOHa
iO0m7Xre3kEh4uTppCc5PVkFId4l5ea3mXAkjbOIx8xZ8qapUPSbb24d2bsa6a+S
hQ5RM2atWuZ+dsE78uOw5HxFM3tgMA6X0KrvxnS8H0gjKLlmqYqjGUQq/3QBJHO4
viwH+deM0s2f+IgHvA6dZiEWKyWf+WypE1MA9GGEfPUs12heohi0kOcx77jiIjrM
U/IDoZlY3T4aZXSXfmyxhA==
`protect END_PROTECTED
