`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LIqjpZu/4UgcPtKGqFgV6gg2PPfaPJGH/jCzq/1AHTPrOoyqKwIh6PHHErrmw11d
k3wNjn8Knc++qp5ozgARQ3ioleDNWxV/UdgvADVgRKZ/pvXeligN1japFNK6WPE4
4Ijmx6w/lTqSjjbwmDC/pAmrQbRc+PFlVwptHYKVunPRyAsHDd0sWQFM5Obo+LEZ
PtkS8Luobk9u6URssuMDqQ==
`protect END_PROTECTED
