`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rh2KjpZkHi5IhC/2VptbVomyuFMi7MxDvI63y1zdDDetXXSJPuNY5MD2lZJ5Jmp+
ctMZPbNLQ1nVACv+CxYqwageN4cAuiRgvC8Uw9oAGm5iZWInv7tHECjIQpCAtnGp
p6Ig4EjMMpBthcxoVnOscKMA2GfnwuZ87I8jFM3deVq/55Nj7xe9kUcw+oDHSGaj
4YRUxASRFkrLzh4ivD1eMwuLOY6A6LmTvc0YzlMkbpY3W1zq9uGDbp3f2jAiWMzT
bmhweUhaS59Rm7sBoIAuajEwX+Xk3HJJt+4S5KVUoUstOtwp7UsGyQrA07ur5Pb2
oGyUWd58cnGBQ/ZZI+l9+ZO2oTHYEYG/a8ViAQI6s5Tkyt3i5daSkMZxa89v5IvZ
sqzxqMhklf9nMmFeIgVf7AowbCipS1oRyqn5kRRVfyFS+nSEJECp+KPoLQSfoZwi
Gtjq4M0/bU9wFb5ikfirgKuELNJvZsvE9ZR0pcMSeFw3ymASBscIBOu95MebtlVI
9ZEk3kWfCC+PPJOJBmoI6N1/slLeesb04AaMN/rEwCvcK7bTkTeJx2TMHpQawmw0
XWQdva62q2/BnlglxUODumfugeUvthbSkNQwP/eo+sEaS7rtK+8ah2+K1MAy/L2h
4/yi5wd1Kvfh+SkPiGSMmOr7z1YcyIxpP+6Pfbbfv8Va3wO93K05HvPKj8VY0rRn
GXAw818oUT9KYsZvF9l43KwY+eWDuiofnSNKZWg1KjWLr1k1PPipeA9HT3Z5WzXv
pZ5DCuwQBdI/nvLa1OmHhruXxujC+zn0L3WDHxEF9VE7goP6YkCbUUUS1ebkXSGb
LrfkbdSYRDxiQG82qISOJABnc7SBFLKZtaiu0kqITT4xCokJzhHgqjAzGjjjbBPy
gFaQBzDxlWU0ScfCJZqg5vLwk57ZlKLWjuigRMUWPXXVjiLvx2BmLZ07Asve6WOX
akHEPIQJw2apekpUQ+hC+YFSKZFezoUnmWVFwpbTuydySh0RETYmyyKwdSwUmDPF
KzezeiPaTmKOLaQkrersLFrGMJa6HwFsXuvPlmUaj+EaFm4UUueOvacxRtuoH87l
XRuGwutXzsINE31NS57ImT4BwhyyTyIh1vJnB+cpIWkMN3Wfa8hrjua7zqsRufM/
rUXntIwy0MVXFAx0irR2ICJIibOQOWqrUMcE3A2AQ29WsqrwSxhCLZ+sfPLD/2Hy
uMJydaiHji41Z4tKIv18xzUejmSZzlnSimtuDEla+5Me5+G/Pp0+IQrnCX6s0Cjy
xRRiS7Esyw1xkVbQAWR+qTpqO+X8dw0ned02l/2U6nO2USXSWDFG4HAPYiBdWafZ
76P1058/977hHZ2EEik7RW5cQqoBGMa2N55kxaqa5hItHmU2MmqiQqV1XqKlYLfR
XgBwy8oKgr8p6LRLKlWpfdKEtYBjb4ddzN0bzju0vofrOT5EjUXAlVnbm2v6JCl8
8Tu4y4kXc93+SOoCaZ52loIN+keR/7PnEybgZJGnahxqCIrl40hZdhjJ3s9I66uD
nTQqCTxrO7Ok8ModjJD134sZsQEVG3wVgLeZlFtQCK8yq4T0kBYosDI2h1LHOI1Q
awVyYoUTLJz/+CRICGA9LJJou7z5IIyfMx7BVG5SZHO8bkHgc1x94k0CpPd3eZ8p
EmbOVKs0517SEXU54FJA1cjk+7WPLWiMIKBC3vUB2UnyZdvoZ7oNGTyvC9fxwPzP
IkNaTUD0uOxs6v7zILkpF868y9+BtfyfdlX4qVEhQZd+RY3qugTluZCncJFQ3air
klMPMraJ2fUb7Hv9pkan0YChjev4/+1YWrycCuwe1crTZ9FehedvTYspmvKTkrHC
xlmV9LMa28lWEk0b6Kw9mxAFMsooaDBx8IWOxC5OZVy3en+NpSNh46uZELfz7fjM
TpL2yGFmUhkytc1utb70gQbpO5jHLLucNob8KDUnTY1bJefxN4om2DSF8WNEwajK
K7NPFxU8Br0PJAy83QNR58WgUJT9J0CgOkw+C278i8i7cCV9ddN9vuvOlW85wedZ
Uc6iCPCvGV8q72eIrMoSTHdOdUvE1c3AgVkcEUXHqa/5Ypu4CEf0bK+pa6SoWShi
9tFNRJDe926ZeGXSg0umrbmUAN8zC5S9ZP1D6mgjBpVGiOCa8Z5zZCPejAl9rIh/
xaEApw9rD50GWl2JvhFAwIqxDPu/714j+TwGg2fOSLZ26sFv478KymAPNqQxrHmG
BetNuJH3ZGKnW2kwhtwRQDq2axdaamUj3DCTnmF5Np5gUiczk4wgu+zgHhtV6Frp
FyUG76Ywx1Sl900KRw2NpEjc0hhBRbj5bumMAApShQeWt27/pPNTIivHUcYA4Q2x
P46g9d4+tM/AZ60hhJ5zp21gUE1WnYYjQe2u0pj6Wc23AEWfT0agu1LSCA8qhBGj
V1G41JZWfTjpEQkPVOzJxGBJPYOWUHH+uinWG4lhOVF2Dri/jXdutsgJ8wHmPHkn
LkWCSj5bEE5ANhQy9Y4ZQkYCmvWm35YBwC0qbVuklbX7RtzS1r657kHmh665ME42
5khc1WW3cLeLlDSrKGa6WsWvNEc//eMq+s/9UApDD01y4EYGfdiDsf5voA+URtO1
I8M/+CVgveDQXtfwKv3/U6skNimpNmVOQad1WOqXeSHXPJxLI4X8tXDc0TsmpQLk
Dco1L6wdzLH7ZUtKKN2sKYTR1hRle7bKlYnPK76GdLMsvf80/pTXA4MAA36FvuUK
OB5puuQ7U4ZwrX+tiq9AEQyMRphkkW6Idwg0x/6MRxa3jZ1XhbGbkk5gF45VLxjW
6tqVPcPR2AC3ouXVEREneUHv5nMfPc9GOrpfLAcRbxYERB1/wpMlZB8tKp2tAFk9
0e7mX2qq93jxC2QVkk1QghtrDYWF8YE6vZjmgAWqMuBMiTLBCbJNL0tnvNj+JNgL
e6CNo/ocZpuQlMLnZuGUbA/zDu7Zc3TXkopNbmWMLTC5kXeh7Z23OhaLv8XFHEPT
o+wF7ItBplFOyHB2FOqevoqT2vo9kjUMAW/Y3pZEFNLUBiZAPhMk3aiTXCMghCmO
AZczuO9m86LhaWpriHFQev/ctF6vdD1gO7RzQ2LYco26LsAyJS2Lz91ljJ6aBeEz
jiCtZbFvJyqvQKfNHu58NJBRYHl2qvbiIvLS+G/XdfSC77dMtW7em7J6uYW/XdAw
COTADC2h2HOPjjCj9IhZTvBFJavM+E69DybSPDdSUYMT9ZOPjFgQN9mRoSTly6Nb
WyIY2/o7bwFUkHr6wjwe1WtOkXSUpgIxrUmCzA7wivmw8TpTkg68DLlPFD+/bNzu
JaNtYpPgSyZBaQw4K8s9TPcXXPQC579YAYm5dW9BoVFFQvF3loxjzCdHNV22F7pg
gBZJF93M6Fcy+1tJZpuLpQCwK6YDzhz/amOGWu/IpLg1kBcxOdupRUCJa7zOYgzh
wKWEhnnC5Q9CvzBBkOpwOk8qud5QSfIg9bJ/nzuQmM7D1Grie3HU+hnrR/Nb0NNx
DKYCL4qmImP0Jn6480wfCb0YBvjc+92uR34JpEUtb9ChzjjoOC5eBh3dHsNc0CpV
MA5hpCqUJTb1NdcjJq4SVrOMPXVnfgS1UYUJQFCW0f2GtsMTGVanSwTchshIlXtS
M+6A8E8wLB6YhgfVOi18DqlSNBXMwZIqZiEvJbOXGMIF8Daxs/wQDg1XZm7JMWgt
OmRN9a597dykUpVEGdZj1qB8hdMWUPG6sCbVbFQiA/ca33ADLe5qvxbj14i4SHqn
ugVYuoBuvk3kUEfyT9lW5IeZb6gx5nkGPjCwWhNx4/Yv3E7XJ6wFhF3Wx/ocuYGY
zsf9bAZV3RThHn0uT8EdU8zHE+iUGVry5eXAKfoCA8RL/2J3ZiZAMicP+V8Tzirg
Id2Hylm5oWa4BOkXPJYKNgPF0dNCQaGSsFkCiomzMRrUJCklz108w+Sqj4U23IKx
uPxoGXBxBmZ19/qa9HGYhuI0UcbM9/N6HgOcuJN8gG/VpHVBFR2zb12fd4q0w1w0
rqYN7xivlL7/L/lKhaWGfkeqX9GajoGYzkEdVztqwYAUvqvDKd5nhzVkutea649O
gQ6/DDQxQWUCg44DhtlDKK7iE0RPcj/uZOzcS5/hlJuZPCLGCHCqT3sva5H0yyvr
6V/wZIshnroajTID+A1e0gNhB//VgsHW7sBPBfEFfA7JDvIe5SSOCwPa9/lbjAnd
MNRFoIwSCrkVf5pWJRctxIV0KWT4acyOAid7nx//2ZrWIAN3Q5IzTVAql05Jr1P0
PCCq7CaIeqnc20Pyp9kizqPSrtRaqjw2wHWicUQSl6m8iYEGrGlSdJ/Te52jM9bu
teQ6X8UcoXKMnsdMd0IpdMhXdOO4OuvIovM+XrK/AzynMUP79ofwQ7bcFKcEn6GW
olsSQbicYdThuEZSsCVnm6dDdmcFikvokqVlBgWEt1d42cyjTvfn7N2Vr3DtByLH
WfvTHWmOfCQtEJ46BXQgHj/TfNtTNtSSFrYyV7ukLKtN0mFOmCmF7Brmg60nj3og
m5xr5RKjJHdPDqBStZiwNeEaXdLyljLOeS+ZsqVfKNdwxe+cl2IP/OE9EnZY6Njr
CtS/3DWgR3acjrQcm4IpyNQc5SqzEhSGD1BGK2xhCL9MHWM0vLDiTERC1B4Kc7go
n1SmOfcNGecvYlWt+RZZYuzwfxW3BMJI02GZW8oM0NvozAY+Of9p/RK8pkT6jHcL
oWm+90P92ORpRv/hBbUmpKEa3qldbe6HXd5v7RETMp7QT2iCoEFjNE+JhaDZqgJf
WuT9kSGKAJni4QYk+rbqjw==
`protect END_PROTECTED
