`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oMwG87QlHMFxIikYZh72cB+v2eXz3oZxBMQscg305rUr/b6Q4Gcr7sS2Larf90b+
GESO2BP8PJ+vB3WD6v9zqaKAvPdLB87HoTK0HEQ9rVHzcVgRN5WyQIgLxYXlkKHI
tyUBm3qHA3q8pDINvmk0OJecZVUkXXGzFnfu1e/dC4RqS8q/ktnhrTh7dnaYl9kn
gBcCViLTYqG9OF9xabZ+hVZQ8YmqIQyhbMZ+5+TPCTUGnnmYAnJBR3/IN26poPmW
avnzVH8U9N5HPINJ1ToLrHDNcx9Il5pay1W6flP5tbzaHp3ttQO6rGOwpXlb+1zh
/sDHEPC5rVyH749chPflDjHnlCcxIBsJAsu1N+bPc2EF0ctwMjhVHWlPy2ZgyngL
9G2iQPc5TjTmd5YB393oqM0NFHFSz5EzAHUZpXVuzAG/IibcnK+iA89+XbZGy0cG
zbfG8OCqV0/wyXzAuZ4O8/F0nEwELV6OSulx8nNeKuXDuUAzZ2iYqGvX03jpfs1b
/0VAPJErPOuwqlC0hVy/3T+hn2Uc+EiP77OT0UbF+DMd+sKG9LLbFdTft4GK9MJp
2b5M40TorTzd1YaqlvvmUbiJ+EnzXO4RL6eMNssI6FhltKkw6Q2wDPHUO3lV9Cnq
XShF1Bcc+DviVCg+B8H+Dw==
`protect END_PROTECTED
