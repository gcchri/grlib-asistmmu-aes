`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h9LG6defbgX4Tmsg9ayi/qgtHJkzoTnkf4dTyoXBA5BQqLha0BX0OI28YiVyl8N9
kOdyOn8LV/rAFdUhgz8wqDlt5jLQSZe5Eh5J7hzL035uI9sZFdJwH7tW6MVXJ11v
VugAw2zqIYSyXggs7APWRcz/P+jIvPM7gXYF3XhMXrT/XCJp5w99Gk6WB2PG7xNC
e2nn6FYejpDfX+0qOgeyKVL9H2LFCmmjFHjMCtaKs4Zf0BLf6mEEihbmqihSsrpz
OrV32zyxaWiGX6wIpXRTBJ+Zyk7qisk9OzAReu07q0Q=
`protect END_PROTECTED
