`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mLVGM60BNH6G/kTxRjg/GB4f0Rp1Wt8Dh/TQvo82BPRZG0GHIIrIXKdrvm2fhDfo
jH0IVTI1W7ldoOP2tZivaG6uS6ju94ThkYTutyagX4sP0wjqUP3ai/8VjQsN3oAD
NTzP5xH9vK94+mJoLAIiLwhi8Fx/BjB94dGi8risUu9cxH4ipjwzL92kr5rhdoAY
8+3vZSSg3yTB1dCdwy/XxT3KboB0iDQGKD9bnrE/6TW4bxoP7PlfgKX4oBsDzK0S
3tW0s9vhJemzVioOxw0Y//JJ5sEAgyszdnYlG07n0zssADCSviTuYBktUtS6FY5A
xpz7Q6DKSkQtEwBD3zahmOWAZj4V78/GwrHCb1XlgcmBJvcUKNgYPE/QqbWlSzZC
fd8s/NU8IbeGURY1IQfOXaZ+8M9LvnW3LqN5NwvEkrIZ3qcW2pnHeBGUCWQvQ/dy
HSqZXxg+lDzBuHz+CK4qwdTgdQZa1XQlmhu8EgGE+VTIVLx6njrjr11NzkrglV/3
KJVCb0RkTyFvmxvShmN77yDwCEszj/+Yqv8uc9CGhAdpjjjm+4teZGy70G/vk6K9
b32uXinrUV7fWR2j+eOwC51cLD2BO3GlGmImWbVXaiM=
`protect END_PROTECTED
