`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dBjJF9qUmgXE7fQYE2xDkxtFgK+qktWFdtXYITIfIgGSw9jypY9pEE0x2UY5Qccn
10FWs4pDSbGnEi+E4OzTD8hvfkjpFRfRJp6LZV1lg7xSn8bnCabmw3D3HFSzhxwJ
bFGZO+A8ptv6VGHjAJBQ1o5M92NsSC/oxjdi/HkE4lYoXyrKk0Lj2Oe5pu/AUzQB
V3z+qpeuaAcmBwl2jhLR4yjnRd2Q0cQE0v62OVhq1vuYyGmKynfnAWhEsf8wQOmU
d5LcOguYBttIreHV4dGAkmkfua90NMamajTSmh41+9a21L2pCNB0d8W8Zvz57SiV
ThAlqe5J7jYpNeVmLvON2WYbHTDoLNzWvsRF+F6f1zcrD7sw2YzvvmX6MrufYyn6
rpSHAmOvh8XnWI8nOilcESP96SkNM50zB16kj1jrlWAMSUXXphfxPCT309+TpTA3
aX53OMFfTcbFyKq7+zwpcTBENJXJHO5iBOlqMUTB1/K//e24r3WFmAHP+za3BF1g
A6wV6pfgbqlFrJdvg1Usz8qMqpOexd+vwgFR1xffDCJ+X2O0+b3f/lS3tBvShbji
iwtev5g+pa4V+JUPWuvbuZuV2St9DPdSYr9LkAy3lW6RiR2b6lViLQgDt1cf3U2x
xpzoBE6b1kEaXFy4QoFfk5KSPSfryVQXTp9dLw65Cb1BKceYLw1CxNu8UCizZpoT
kktiYwLXhuM0aQftSBidXVawJ+yPHqeaJRqmAKoijEk8OA0mvs+AVBJ37NcGM4aa
B34BsR/+8jACNQX8OHs9fUiEA5auroX//IzQGwVs+Jl2+6SxVTnXYEFdKQtFqcWh
WZxQoDigzvXmQD2lFKW+FMl0mNmkD1zd+ExAEAC1tMUUf/GLCunvFDzNM+Ca3F1g
FvHz83aBYK/Zs+v2Oz9J+LjwbDWHzCLYapvH7RT5QzHXGi7h0ZBm8jXPLmt01HCl
x826UAwIThG+j2rOnkP5fdGpgmHYzfpCeXjpdlrZ0yH9N/Jazs0lOTQZG5h9NTjH
8pJHZNVE8qXsHasxAiUYwWw6oKnlb/7RPnXjgBVTTVSMCrOqjvM+V4LBXYFZKKyS
9UfDjQ1B9djA7nHcSNnnelhD2AyvQXkiBP51N92JSdDMiv9/P0HvLzNawuJJ32Yo
1UqCOlJcLus1Ttb8cnj7KlOjwRHFPYRoc0dqySSC0KxxgKz/tfkhWl6euzTSOiqt
lcW8Rkt2ypTWxdDi7/8A69slwA+984rXlmy8tg0vdPpMhoTo8Z/XCoYot54yCfoR
4GxiMuKzJp08BwwiDaeSAIFYquuaNzeAyRaVxKokQkHVwV2DQTpOSCml5AXuq0Fm
zc0CzNQCJbXE9R+4E/7CWkzVZSnwZM5/20paRzOu8EVe1PZ8JFOlKCGVIjXZ+kiU
uXAoCRyvVBg6LkLjURWVTtmQI86f4fn8IAmzhF+mWmqYEJMKKHpssrEtxyCVhjlg
GoPHjgslwYNJPKZgu1S4L9sJburDyqM/UMsfmGawXmvrsx+enwy69Ktvjwf9nJEX
qv/O3Z3wwOo1ONzV2ZLxnucMeA+GDezs2Y8EuB98YHLYejSyZOf7OjUmHh/1EPGq
5PDMRvyLWH1SDXgBhqPmJV2drgaKlXoxQk4CW32d9BL/wXPIK73XGhqaCu/kP5WJ
O7l0hZW/eie5x+v/xS8pT6KLJTqM7YaViYxvlAvaCS06e6fo+gLBkMWYXu+3qrVi
2eQhjNasEW1C6hoLzIiVuduXHM4kUIk1LrBbkLrCCVOyIbkqm674pl2mg3uBmrPR
Cr0MojsSrm1yuKvVySBNGtmbR5ar9yR6J/u5ypSCGkbnYglvDbL9GPZjFGMwI07F
2hV6vWSvEaekuVtxqG811CzFeTTvZr6vmZMUtRF6G1iGcuYP5Ad9OdUB4lVxn2a4
3kBLM99lW0Uw0+BcjS7htFuhtuotacwb3HKjCwkhU3SDHIQQRD2b1uaKtIvV4H4V
AFgcOe8tgSaZXgEWaqBt6ztVgyDGXVypCTWR2xHbom2An7OcRyULidjhvxu9govn
3VSUC8KI7kDy5iBfXnOvBvarJ2qdbESz2UG7ib8dVrRbEVMNpLS5K+LH+7VV0vFf
v+YIAVy/ytoZ4bRDehlbWX619r/CZjIHKxzPC8lYAqeKi5fHsT+yLlzsz4As2tHx
EsIGLhTU7Chmdg2btEWYxpkGxUiEEzniQNmNV8fhsNmmnhAbepYw20OwOupBg0xJ
ZddxPKEQnap9+kB0O2HHFchn8xxqLL+bs4QLHpLQ+EOuJW/tNxUVF4PJIUIDuoyP
sZ4r8NigPouJCr8d3+VvA5/uNB5r2GP1ZR9DfEir4t917qmgPGWQBWeaMLIbkjro
qmMIc0UxQIisplUCMLWuzp+Ik+j2XzOqGRm3O/TT6T9JXtagz1ws4mIplPHjvH3x
KN4IZW/l/uFTdlwtVeRCQiGq8F70qYaZ5Fcwsiyba4C+LGDwz/tBXMn0j+OCw3u5
m/baOLDK5Flc0YKc84geHIEdGDJGPq5etN35vMzn8a3PT9mQvd9M0ywhhSImwjXd
vqxQwTG9jxkvVHb5sDZOVHCwy8NKP6ZIEUtpy+i1qKIm5EM0DvajxIUVvkJNnp7f
g1zhLJ8yxthXrzD71t4Sc/ZbujTGhBGnoAAX8QvaWbQL3rROhvS7wQdiVlHvocUI
QpT3tGdD2W1GlqkLli3L3oDha7DgCPAu8pyTqad/q1udIlaBkVc7ZEzO/20Oa9RU
iwyfmVC4ZWdnEqc0/eNYaKZLgVwCL2ncVdKVb+FsxzYD+wRB2b630oDPN7EDiZbX
hgbY8wn8mVI79+891r1Sso8QxgLgx1mcmTGBNgBIkKxPVw7VS/XTE3CdNjADT4D9
Gsj7Qr14SXLHuIGYIAtxRoJVOmZwODWioXwNIc6XTo3IIMwXzM93cgN8TTGg/yss
FhHtkobo8pS/rZYL/PW4utGiW5b4wKmUkwWwqrDxn31H32ki7HT/+UllJtG2xYFR
e0t9K62pXIZiIHyNiFEMYQiDFo1ZRFzTibFR4EAvQqlcFDWjv3s1SXbJeCtpQnuF
4XYNFq45y1Bnpnpc/rXdp2pl1Yhjy82E4tIpTKOHXoP6nx6T8ZVMMb1zwpuBzhIo
Aw+7ZnTJ7z+N3ua8HFLCRSsbysYhOwyorAEsQXSUbn2EVH8c9OykQ+9v+VdgVtee
pLRKNwtSZ2ANZk6wyEZRqDUHa6MuuekAkWPZyoBqm8AlyukmdsmUclILDNZUpUxp
2j+l1z6e6nn3dqRsNoC875ivg3p84CDvOCWVRzMnFESAV9Js+x/giDYT2kFFagzl
u9S0q0T23kbd1y8xvqQJACY0AGZsyeHd9enbt3dihUVs6YN+RykzfDx9tDhx7YhN
YUhPOyjswflcjoZ7G/ZW5pPfNN3wWU/bVvijyaSITfsYklDATM3s7UzA20BRGc7M
WbDMxaz8xULPO7SJ9unyWhJ8n+aU8itpJ6JQzjJ1F7OmOWAiTbSk5EBoP2AKryzd
dOl66qEMIih22C3gZRPTBaceJ8rSqMNzDFgmzA5cTeSdDk1x3qP8nA9RlLlMJhsk
8Mi5prfWC5PEYrxhtVU6CwriE/d73ZKOzkL6SJk/KyYZF+76SLD8DPSiGkGgZ5Dd
R+5GTVxOYdnkPK+SUrhzI2/X9Bgy4LUdIKCAuK4Ms9/mWOt9ZZtl1ihrtAWC4MnA
Sc+Jc2q76498tC7HXTfotkjOdoqVsBZ0bdKToKAhWmmYGrImf4HdFKSPW3VJnpyf
oGK5C9KF58Sx6I/W8Iglu+9U76KEJsOtApXOye1XLPupzqrrM6c8LTd8ab3hmPEG
0/WhyFUi8BZjM2QVVeSbw3WJe/SMZU0HYAUqTsM6uhkNhkBtytk7NC4wILIr/DIY
zlUw+Ogi1Cek4rq/g+UsWCNNceftOvXIT3Jj+287qUjGuIv398/hWWzbQxgZmwfU
QSjkWrgwcKyjAQBkAL2n39Yb2OOmcESlae470Ptoz9H86EAzXIXYNBPxtTE8XaOA
C0mnkr0xUhGYVWJGLEWlFbacMGEXIUaO55Ui4ghhqSi7iy3GAXvedBb87+RfoQar
`protect END_PROTECTED
