`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L4E76cCEqYilFIRLmT/yoF9rGCPJXKybALt7yLqagDRZYy09sKSOH5BcmaJFMlbf
tNKz6F8GstcCD/YLeznG5piv2STXo08HFoi5wPznNOfbofF5m9WAwCByaNZQV6s5
M9VclUN+dU+YXEH0/d/S8fgmxXaR3a8gBivIIS65HIeisDq2EE/OhaktzXu8qx9X
/Ji8cEXEzkPr9SM6s43BAPdR5ERtUxVTNoaZcLYMwzPZujZdxetqSJGFFhaRAjx4
I3Wh3Sxwuy0S5pVYPBLSbUT8msnhKHCvvgWKB3KsOewDCAP+kSGt6r7forZIELGq
SoRYqK3idnuYDlMkj276EjmvG431ACx3EAUBylt76mv5yyJ6p+QHhZlGSFVA03GM
g+jeJ5hPQv6jrgLbi/E5ssfl6F2dEruby+puBaQ8fpOfJje1s76DE+akMwji+aXn
rT0fsBuDqKC0PIGihKwb2xLx6F7QNPnwTfdFSmuVaS5x6M0OAVAU7VnmJwKMhWrF
`protect END_PROTECTED
