`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sQ8PVKqcBgC8Lyy1bhQvO6xMU1hBWKRrh1eSnaj/JndXVIV+vhZUAQbyNIMqms0e
6skKhImmgORD6TKHipRM8PUt3ml27/OsCGGaMPV3uzfs1YC4vKHtrYqxFSwU100d
hI3uKy76rCwTSgZACtmGLR7EGonFnizsMCsCSBB4Mj8jrZ+XvyLgy8Yf+cfvXFpo
KQhXg2VaH+IufBzSDt6m7Ei0By1DG4ZRTDTfrFn6X30YYEOQ3lYAGPu+sUVBFw+T
ZQZ84jOpX1wcNZzkyX2g/sUBISZ1PYk5iRhkF/kqgFXfitycbQMWUWmmSimafp4a
YGhrdDAMklBFWVS403vlo24XZLauRB7DHWITr3c/xFw7fxZdhRxXxyIgns8noIyt
4iOdtTZEixaZ2BiJPZDf7XZzyRW/BCkYCSftFKoreRD7LohHfYfQiHzUbu26o9uY
nNgpbS3PksAS0xKPI48TQbIynsFyUTu8Bqp/A/qB5LVxZhhBBPMNRpz4mYJtH+XR
OtKRJEVxw+GjgRzRXWAmensYNalOh4XB9d0apRiaXVwBcHlfTVBB/9UHhxCadRsl
l7bbYTaSO160N41lDDYuISHnCaWQCzjj92derxF7PdHqQGoouFJkOgxQ16Sp2Sr4
M1zLd4fg5S5A5euLTed/AmVKuVH6T1Yzk0GuoUp/SCurB2X2+SPfDD+9oIS91d5w
VgxdXVn7m/SUeQdkfV8PRdFwFg79MuRU0AdXVxZs8ZLoYdfVKpt6f1vu+xRKgNWt
DK/zZ07PE3IwYTw2/MH/d4eS/0rQG5e5vOnjf2/3x/km1GynHJXX8ZPmeIYZ6ycB
OfMUMw7DkqtWq1S/aKAN6CayxmdoIHDMvWGDntwgC7Lm4MG13mhBDGz5NmpHkdjs
3pclVCvupxYBUOQvTZF+fkThyiTx9hXEY5gUFRxm0tL2Kay6WSx+o0+j74jnEr2c
mmbpS2woal/IfjwiR1LOSBPmhzpwc48rpze1CYyad1sUyWbk1bEpFS1FA/UOIiwJ
3lPvKUNhaiH/44R9xSgU5j5zG8GSmk/5wHdpVb5mFjIDrhsolgzIEDlNkAmDkMsb
GAOLNoa1eTc8Q/AT/FrpzK8Aqz3DyedMJXSplU2r0A57P4rQ1ocoZjy/YGp0798q
5QgZUoT65QDuObq/a/uQIPVUineb3zaRD9eyFMH8oRYTSe/1gcqQ9+A9dRsN5v42
Y9IyMOtoS0sDa37/Z0X96phJ1+F7WnsQIbpAu+kqvhcbuPHk1pANR5J2vBtZ2RT8
ajRsRkMAvK1dBDPSdNeXzpZR4+txN1yjdUou1LsPF+TQgyCtiq5c34+/R0OTpjre
Frqbt52tpuVIuxfPIQ391Uq+iyYgzdEHVUeCLO+ds3Rg01GwXfkdhANtOt2dWyvU
jZaU4FOOgT7oTLxBp8eUjNXeBnyusQaU16up5oFOKWPQ9seHoaM+TZsJcpKwyB7E
K8jauipy8Kf+XIbNj1Oh4S+dMAW6wQbtxFiqZE3E41iBYr6TLHdTujWNPKV/5ez5
CtSseyNfub8LOYZX2vWfASnkxgaVLKpS/5U1bhSCfivpATHxdjtVhwBV4kIR9jKG
qd99KxNg514lDjorMVop6xGQqi57HIju82lLybHFY+SaUl5wrzfiejk5FuMuuCp/
P8Y7gIPA9dwA7yp3++8ZV7GX0KzCmoGCOCXH0l/D++RjPQVeKIeIgpQnYCCvRnDc
7CW0xwdIuWajhjseq6EBvL1DVfn3ccVYq5x92hSNF7tjI7kZpvxMw9mPXql8eity
ZN30QAwZflhmNzxggff/DQ==
`protect END_PROTECTED
