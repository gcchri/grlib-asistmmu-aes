`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LQc6q0pyhRKymm1uvPhYic9Uvokx4vec64BeXuNJS54iCQCtul9DhFb+F44B5o02
HDd/gJTZoRhoUI33SKsbpd60On+2ZrxpR3FD6FB1N7F5nks+3/UGSxeEGuZa7Dsl
MFrps3kC5y4+IyMQP/8DuXwKl6KKtVHJ+h1BMewZpXir5fcFl+T42/trtkeBFEmp
s4gbj0enu5thKkuvzlFoATp9d7gUQIBVQ4k2DpEtuu0mlKUcoxDwBm+aNU38gDr9
gFied4t5ZFCSQ0axxblZH+K7cb6ATiN3r5TnJT1D16rdUHpX5za8tSEVYEGPys+G
qaWtu19/gTdtzLm2oAAu+B4aF6bxmrRq6kK/bJ4czT2IJGZZyGC3A/3khGPfIjgU
mmpzIac9ijmkM9McqGtzuYcvgRuJNw7bssWGDsJJvn5uSi07lQVgXsDrkCYjuFPR
mzglssfbaFpPIoXmOHIspyOkEZ8elbuA9k34FxUzJIhxw3ObG8nqtrGxAKIm/8sb
`protect END_PROTECTED
