`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NI9bTAHf4itCJhgIxGsJto8WZXzK7YC8O7COHniF5yvGqT7UtcY60io0UdfHd0r8
X10XMTh1DlaQD6uNFmsJtgDah3BatGVsAcr847U04N4l+4ANz34sMy/WWmDuswgz
TloNBc0WC55fP0Buz6XtwUuda8pdkslb7Oara/Bfbr+TEJAdOimmPDrnVDcOYS83
LMJOxvWuHY+QMUZt7zNeD6fD9WMnDPVkj42/VzWbD7HZHB5rJ6Ndsi00XGKhzn/z
Lbf5Ua1//+0Ini9hB7hroL55PSkWB8HxqB+4cTyks1PU0+eSw9sUPYddt3XTQobm
+HUOTYHnY8LBJCzMV662vQ==
`protect END_PROTECTED
