`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CGtlRQDEHw52S12fH5RbKn0uM764sTywGyKpq/fCp4TSrDhKFH7W+bk277lFpnLw
9hQlGLlM2WT2Qd2wyg1jLewRbcuonG0fTf/eFh9jfy3//Jxbmv1a3JwgFd5cEj/n
cGDNhBdKL6bj2x3S3ybC7XXgSu/EoLvRTeLufKSU/or+5C0W3jP3I6n81g032Zq0
iSKngcVp1zmw4+/0r/dCIoyXMXchceU4/xIEePoFZ6ab3NbdA8eHB87vAxcR8VG0
mzzRBybhQGZeLjJu83ZhFldsR1I2svhy/kJ23OBqqoJp8OIZPvanrjA7Wr9A83Hi
5qjeslhifbHPNgUnVZ+yV1modknF93I0RFcEv9rhj4i5kgtnGr2dm9Wup2gKo/Pj
gzeN3E9DVLUgRBJS5KSS+EXZEMrS8ZrxIccA0KJeNlnMEA4Vo1pr59EQ8R7vGTp5
12b1LTGUuTSHKNw8rdA0TMBx8LJOGsl7QHAnag/BuzI6+nL96iKLW1Es2ctfI40W
3l1gAHhh5pkmi/ZUJvRdcpwDsC2eaL9y+U2AfR7NtdIH+hoAZDn1rtEYxusXtmwN
eT9UEFiAK+Qx4UT3Fkw92GUZS3Y6ZhoMPCyu5m+W3eEwevtwiJawaMavD6zGkUWC
mdRQQ/gqb/3P8bdC830r/rG+Vu8+65VHdEUptUpX+CNKmwm9/fzrOHKmmm8Vd6JO
7d9tmxJ258zE8ZnprbSX8gegD+1hbiVKrISH/W4gcICf5kBEQ/USdc7gEa9pEqc2
de51MBuTP21ZcChuwLDJ2ooUbksISg5O/Z9jzh8jtyM+LCHGQ5+48ldHMHFJq4IG
7dzXPF3AUS9oiIhzlFMgiEm+405D44vef3rWpwittfwAxaSKkRIQ0pXt3re9AvBr
`protect END_PROTECTED
