`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pcL4E+Q92UA2Cn08rq8X71ifJ2xDvnGtrFr04Z2qTaHR00yHs4w4W81ScHKax2Ay
N5XIfKOJOg5K8y45N76nF3a1U93Qkm02VDji42uaDlT1T1ZUdVdWfkDRjj2Xroz4
xf2QG69fPbiOE5NvgpPNNcmEIbOBBZESg+TwsTRBUwbknlfcezscScKLyRRduqvH
j3O1XdW9EAuh/pHa017j6XLF7VTg0okE/ZRQ32Dcrn5gaXMDXojvMnxMVMYWjz4L
mMBfuHA7kxREElpA2ElRN6JNyqsQI8iOOpKJM6RxH5XS8A7ViF0uDmk+O8t2LaNk
1wzDnWl0vywey8ECVD5DOqYTAal8oNAhJUryaMGxIZ1QFrePmN1vcVghlJ23pC0E
fkmk+HeqsC3ok4qnbMINqg==
`protect END_PROTECTED
