`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ohGi7JdMI5w12tcOzi9/4LdZwm/JVbXAnXDLWctgjTcxBwTnwKoJQnGk1BAQiKPJ
rj0WWTQWQEItvXDQAxCbGzpeWQx3XQe5f9Q0Fsowl5Z0nNUxBMx9/ioR63pv82gT
PjrZEi0+kNDPZukS24xG0+2WXHV5rKsnLXP5gmZEJJoWgu6d1RZ9cJAFsOCWSf8C
S2DOm2ym+Ud5DWv04PaEpR0n+rwdXZgQiATijHnNxMzp2sRlRsH+9RqMiBUW9rHC
luqxl7m1bQMuQdh4a2rO7bxOwm7IrksC7BF20vTNe+wjCRb1BBeCVBXlKkiln/4o
fMXDgi7lsjfljOtIm+SPlVGsyrbUqKjUUKYH8UlP+AqC5DmsdMik8UuA0s7YOvK7
G+dLjPdLjydAcISjf+kqTw==
`protect END_PROTECTED
