`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
37AxyyPpiratXALawWFi2ahcohtd6H0+fIHpxqbh1NhoOE5cztNr5zzsKFOYuWZM
vUnQQN6iiqp6UmG4W8x0r3MA1FoH7ghVf3p0gU7vxnSTX3ZdJ5jEYJSFELDjaIeW
B1OkV/1KklKAzWs7TrjOBrlSe/7l3KB2S5zmil7B9ynzGSxGcr54FfNWyo83wGss
7ya/wmnyo71RcBFZCA4IXnPNntw5bfoBvpZJ8XB5dkjkBh39VgoM2ii33m2TEtGr
lDBrKn0fdE5ycE8bcOETV4yQ7bMhFH4vrTTAMCG1BbEjbiWLW0BsHTaRr6YX5M/V
YTYG/ihMZplj2rFziPf9AbHsy6mjgB83VA4Mbt8/chocZmitis2l/A48YqKfwTQt
MsSY6Zawao3WRyLZa4kCt36wFFSAhGJjLcZNaY8Peb5Prbp5Vik1rGNviFxl7ife
9bqMv47rsXopufKjDBKRHhKF8AOGcDqsp24VaNUZZStkWVitoofqM4MRxnTPRhEh
tmzNt1wsdylxr9spe5FObga11s5iI/vHpqmx0TlK+NQJEMbC/ni80c4tUewpxRrv
zM2mlspkhI12iVPyP/NTu2/Bn12nLvluKpqJMm0vWURtbuLSBKJ51lbNBE6SAMzB
0he5fxCcJud1JQu+dfoh/De8LM9emEgKnL7bCc5AbOQ+sZDOaYXU0Q4+iG8/I1UF
CndE5qS7F2x60GxnkbYkpmD9cVnP5C3MJiLbUzqHKJ9jHL7FWq2jhUyFqfqQk0Ge
k5cxN4hSZn7sGWqPMo95xwod+vFh7Jz30+cxS+AOJp0MxbysRP0KouZQZ0CQY6iU
QzdOrHOmKOs7INJGGdLznaH/biVkojOp/K4VqyE1Ad02AUlvKxMDI1xL0ux7jkk4
hu5rQ8yg3wocmZRfmi2i0of1Qs/JM+MT6iIQJthtYf+UgOP9VHmMRFiKAYd0JyuY
8XlRwF1wRDw47akRpSQVxhBhKe3tWqjTNFMSwQknuETHI9jSrox8s4L8Gw91ypar
sPP4yWNJcqrF8fC+W11R1nv95YtDq1tStOU7uO5Vei+ZYPTTXX7C9G0VU3EFqiz0
SUAq2bQf2in+agN3U3qxW7d1xrD97b7vh5fQyysHAfiXPe0atCjxr1huBVQNbTJI
Jkk9+bKWAYw+dWQGTkJyt6oQXGslbNlUX0byHpsBuQdDk7uNpQvf/2D2gp0o+2wq
XhDLhNW6gDrcyT+RsFABvSevUATsnILiTBh8i594OD3qx0ixQAxI/Oi9FnxsRPTM
5x11adufnbBH14HvQWrz9949LRcO/r4KAJ808eBATfKrHEN3VcyZt9RzOMadaWNT
vM85PUMYF78EPxneI1sqJgpxvPri4Hj9OqijeN/tnfWlksfLz5eYyd1YavVRwOdj
yyZ4LGFAIhRWkrcp9FPr2WzocM7DxlhqBWD9VdGsqdYh0q6gTq/oiHdUgypiv857
WiwCCQyUG8rc+Al/PbilO9FY4y0/TLOZtk4fH9LWgE4fmSHG2Igh9Q+pKbhpYxUp
BSSzUltziSU5s5m1Ymnx41b8IUGGa8Gzmfvgk1OyrK+FQ4QF9kWvajOOKgrEi4Vl
6AglwKYdKODthMy4107E5Rdd0ox58k/Dgks57W5RcITQirskBOyEsiD3TkesI2WB
sJ+FsugenBFRuKjOMj+lJZk2sPiKFE7cVOry2R4EGMSEi0JJilb/6cJygQvaD/Bg
FrTnWUQGigDCkMRtqYhQmhldixUSbN4cxjly94QalqXLdYNkeuGx9cAYs4iN7gWx
/zrR1qZnca/KaaFfcWam6vjOMQMDD6bEGAoWHOpij0Mkx6GrsKdrCQ1ohRGtfdUF
8ZHeEBgAAsiQ2x4AnTefVhanlCE3rTVmsnFZvYeK6gdvm6FR7lmQ10fHxucfs98u
RGOiRmUEmz3M1LuHzTOznWnL3U2wPTdzSklKOdBExprzypHhiUI+Av0gdo7i5Rin
umScYddzPXhHC6ox4tpEzD6gfsg53S3A4q9Q1+rtKinACBea72sdwAaTwGaDSRCC
ecOmUFow9xSwnI4NySFsKaRxZqvMVle8RU42JytZ/+jyxmcO3pLPnFiik3w4oYia
Z0Z48U5/6W1Dkrfj6z9VDAcv+2m1OaFkQE3WwILdoUxFE4dj6mx2q1GuD8p1pMj6
xz3HGJxFP5bqB8Hz3i7A++wc4BVXtJ9GT8j7/wrVriRFk3h/cye2k8PoL09PxKL+
8j1sAghd3BWMsbd9KmLAAK18yRQg1Nmmqf3b6o3qQ5rcs3jwW3uQabtirAfNceWT
OVLw8XspESkqjGSRfK1TopuhR3kVAZq2c6qG1us81mOy2OoxzXZOupkdMJ1xkbzU
TPolHdRRfEIQ1mk+QRzKT4dNyNLEPpGnr8t5BuTrppMHxY/wxD6ry8N9bJOSBcAV
F+0iOFclgNwd8YYha/vQv/H/1pcJKkjmRczj3/JMt/JeFYUoVaW50yH88S+xk9uH
uycuHpHmq89v2DM/dC+W00vGw87F4ry2QEz7qnMFttfSUEBTtLar+FenvcOrK4zX
b2Qrab6HvvBDBWD4cU1Ck7FF62nB33ui49VCt5nQJmMMrPG2/sANPZcASUmjUUxa
dDqrrCde5Wt467elirJa3kzgYDTYd0wOVDrKH+mKd35Zuh9BCkcWRepxRI8TYPGS
tml+eiT//02iNQyeUpOBYW04Fz8b3wMoEjZOMl5jsfDobyiHFFBb4m+BquST+Nrj
nPpRDgqFDHRAZxWINPgv7jMdjQCXdPYmgcoy+cHits38zURyw9M3krutKn6oJbKG
Be4H2luuv/xTheodjqHcHYuvT1JhFzl5Gx4NNrY7OgRx/WYXbJ3+SGN5rzfcnY0L
`protect END_PROTECTED
