`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y3DrTWOewNdt81WzP4vhzHRySb4suvzYghOOTIXqeo67Yd7V9qYmwk33Ga1Q1sRU
WZZOLZTguHywfYtPnUpjZm2e16l+h6yfSC86rOPDDam43yZY33PNY093/vD+PtUw
FSZUwDfP1ddAlhfbcyNDHxNtIGbPt39jl6EqVRhLtgw6LRfdD2IRVtXxx0/CM4qx
SCgBRefamvPTP9o1WNXsDaDXE+iJxfqw7gltYCsZXCeGmpUUsgoK3Dxq6oR17Vyt
v12c/B8W65Bp3+eWsDbb1r4+qkHPRkDuF7FuREyAw2s2EAsYarEpF7/kK61c4YS3
iCjTWIX3yZjoNtq6tT8v6a4W4za0D4Xf8rryQ4qIGVxIu+G4ZrVP2yGOd7D7kj2r
2bt+iirengvFp6rZeSdNmEOdWVUky5lnvBkie4Ce0+w=
`protect END_PROTECTED
