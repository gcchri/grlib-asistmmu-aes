`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pUhvQMjQOYhyVqe4TeJMezIXzj3+doPqNrHk8Y2bz9bmyp97GYMSccuE9rIU8M6y
dIhf+2Ys2flrvYh5Ws0LI2o2lUoGa7d6gyCcnxq3sBw0ngQcSETDnGjRBFp90yrl
KqZ7gtRPiue5HDYohofwc8SMZ23xJuO8w/duAASw1+fId1aJdYhLhxDL+jI5l0N+
E0klnlUK/7YHSYBc2gEUlKenA2AFQfmqauC6fXgInC8bVI7X0Er1aGCRJW0YReGv
9zof6LA2SBjXE7fvxXJ1O+CnOq+LlbhlgE+flbhqADHw/O7ePWhpEDWjy/6Xm9IZ
XjzuyPfMTezM7nwdS/bCAjdMquPH8WgalLFXbE5dYDS8ivGuxRlXCGsTC1aGv+WU
2UVv9COLbrAU8IlQJ9VxFNLJNggBaDqLhHG/1zQ8jrJalhq7KZSzjX3gua1wG+la
6KRlAZHIT7hT101QiYxTTNCwVAKqbSpgaKNfbPmgYx+VEM29qL++LK4uharYTZX2
U4qCJZV/Hqs3HCEsIgDoNe8LB6+XcQKgqnmy7ccX76+mjeZxSExXpqcaXSfmP2gN
E5MorPzmRqvmohsT1Q9RLQ==
`protect END_PROTECTED
