`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BMiVVr8xpMahqQ2fmkEnRlZKYLL6hNqBCTLs7UxkMVDuDJwdfZ95m/nZ7RYoEMzh
crnqR2rsC3rN3AjmutZnkM3LNSXLdAAYgQIQMph2+aWIDE85lclJCABPGTaX+C49
x6jtWerCkqZYHSgEVZXB0OuGQ3jZD6iasT0O5MkpoCe60NVyGxn7PtVuTPmuZ62M
ouf32x8OeOZnyHn3D+W2uLns4qzTcFR5WX+DwAQRh9FFxp72nAkTf8FJoAD7YA2n
klLZ+cJR6QyyxcdgHCYVmPnwa3Mq9KQiHJykXsumPY3h+htaSzWDJN54mdcy5Oob
RC1F8WPrYhya7fkNpsdiMiP0vV7lq/a7DynB0INED32FSzaPYfDmcruwgK24eVy4
6y2GjXj6VdxKdJefA47dEwCwN4hIw1ob1yTpia/HnNTMUBAq5uSYaCPCc4uEdrzf
9VV3reYa0cljPMJmLkbJvrz4Ht8GDfEaIuJyJ1asKnosi7UyjxFTuoi6MCSF69Fn
S8A37zv8CXzxWOtEIe+YeasQYthcfnygu1xXpUZkfK2lCMd0awkYgVQ7u8Lkuo5Y
gE2vEn9D4/3p9j2bY1lid40NbYqnZzERDDsHnExnBC5HPy794J1QocMBTCm5p0An
tzbW123iLRW8+vovHbLFa0obhI/YLjSwy6EwNi5vem9btPYIhGmFwS1rVcGBx2gf
ObURY2qDWoUEwwcoYvNwWkO7g1u2L/ynDvWSmE59sG3ksHQTe/eurzkNcYJNj8S1
LajrB+1VFFjs0OrlO+RFoXa5oWyKaO5OuwLALEs5BUR8e+y/v89b55aRDOx/fyuD
S1su3HBxqjwWdi6cnH9MPui2y2cVpTYHanjgNniQ9QasAwmoaxqwLsAkrsxiG8bL
bmz//oNeMU8GS0XCCUjl2F1hroUFECFApOdNEzDA+RKHGtynhERind+E6SF6KI8E
2lPqVGwEsg+VxGir1b2iHFgoWl4wXKWKUrj23Mtr5tFtaLaP3xvTHugUU7+rEiUZ
X+2vPFnuCjFidRsDBLUHzAIRs4Elx8gPrb+BKtHLzv4aj4T7o6QVZCSJkIoKcUS4
Cz9sHUSn+c4U9jTUd/1ozJIODZDtXJbSaxdsIWMrGyCQ2ydj8pmaGkDWWVmF0FVW
t5dfl1XwXZpjwXvk7z3QktNVxGWeDrNfloZ27wqJG6EQEhKQnCxjS+5csoTMfvWc
tOLIfCNm39ylBjZPQLOS8Ai8skgYC2AjtJ2JsGS9q2+fgJoM7MpMpvKUBZzVkMkM
qmNh0aq2EjNiTqkbG//yMA==
`protect END_PROTECTED
