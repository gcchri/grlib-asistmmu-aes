`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mRhlNB88s4nnFgqflS4lAVoZn/I7mOsmfOoRGGuEHzB8iGhrx7F0Wd7Wo/vupV3x
ZpiDhKyF3WdQKrgjfPG8Z1xzdK120DhvKEO++ARvKb5akGA3rk5xgcGtgDwTDQyH
QbFGy5+s5gthY+xRNBfNLHySoRSVQu0JHGPjETZebZDjekUi4c5hyy2D7Z31z99k
nAD2UtE8aL+1f0dk3naTuoUUuCodNC0EaaHIVZ6DZJ/iL230PyQygHrLZfuim5TJ
/Wh6VOpSN29hTIGlAGRKzUQAzq87bWy97CA5nP73pTtsqbfYNT4+/wPJpZmZyJeh
SOfWkrHX+BWdAPVy+2Rqxw==
`protect END_PROTECTED
