`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
888xFfYjY+lQs/iKH4MuAUARKOBDXNSAKj7Pk6CEe4yE7pvXkb9GeWx+ZWm03/JY
wmcwY1aDMpKBA3vmdzEua86uI1gfnS+WnVW/PJrCyiCV5d6sAwhGclADORkuCjiI
7brXZGyInOcYIlNNoqX+EEzqL62BgLfoICX7z/Wcavdlv9ro+7IZ66ot34NqZpTa
GOk7JJ5/2CZgWXTFg6TbMJMFuRKl7x1G6dH0JOGn94Bs90qHTXRZpkVsoQKaNJ4h
szrU1OwnuHzGDecjWyWxu8e0NIPChtHlwW6i8/OC8WQq5BYUaJ3Xrib7fm7ECp+Z
xCggzQX31nXLX4WAgHCRB0vlpTkww9v4MggSyKXLupjZiORbvnBKJn2Ww4MxWbsC
BngJG5c63kMB4bPNMWAVpAtvzpkLNEz7wAaH5FHPf9l5ab0rDigBpwibUf9otD7T
JZla5ueV24QUjnihPeGBUw0I/lZoupWVUC6Q9190adzgYvhs2gPU6IPJCejUf7aV
01yC9xVkzUvAZbzgdAdAcJI8u4TL0T1ECH8ORfUV39Ihm4sfEc6URSa3pTtG0nlu
BgmzaO62xYRmxoJEcIVqFH3FjmxqHWQHgb7PMy3cmg797d1Ik52jnLM5GiUiDHwd
T6fB6wigFen/YMxLYGjwGltWazKHxbtg0MVp8Y7Y3HOuy0DuT2R8Nfhmq8S/69BV
AAsQmHFFWxTZj+DyPscTVw==
`protect END_PROTECTED
