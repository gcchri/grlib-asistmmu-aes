`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wwGkoIEU5zKEf3rTcWGKY1tOsEspk0w5nuPc0nEAsMGQZwPr5rSYZ70q6dzkb21a
qJnFHvNPWt4k0Ow/2uqtJ2YXvoMaBHnaTChKu5118hVr375PBPRX6v4t6q1jYLCD
tkEcEd0b/cD7SHUciZ0ML+jdbibLBXKEflmbdym5NBK9YVBvGRQenCvmds/NZMEQ
fTe3mvr8jOvlXP+Hq1ZrXkcpQ/W4ucwOFXmyYJgsRMKkJT0Cr6TNoUD47N1PCVPs
vccMiptukD3dy0+/R9ZWv2gAba6XkThk+/K+nm9NHbgQBvUOMaKVsyl4yxXOlE7D
8avdfV6f5m8EL+ukiouGalX3elQfvjU4Bawpbs3QQFHBb1HG0gW4DU1ElqdBeZfq
aopSXn3Z336+kWq56MhNDzeAtNgQSIpZwk9rf9mtMedRaQTslQ6LafuSQZhef1vu
onQgNH7XDKKK5m6sI/6A/qGLdyJrlfkC4mAKLf0YXX+MKTkE3zzkommm8AJUf5sk
hWIu3L0eCXPQOBp1gv4/MqZ9lZC1/CytDJBZK/VF8gq60IR+OCLrVpAe996qqHEC
`protect END_PROTECTED
