`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fitVQyDwuhwoiqlpbAZ4icSCOHiRkw6g5h2pMAeEi/6PnGF5JF4wo3r8VQc9WQVF
QOWpKcoIJN+SztzitxETxGijteslVkIbJNCar4h3ebleySqsulRwlsYGul3Evfkh
v3fjfnnIohCpkTNYSG4a+MNNAKOyISzjjuoIkVBZwtxnPCxacBNDhPCwJixQuWus
7yefjqCbRsEKmUlGOFCWTwASy/YBQ6LFUqyj8Ahagqo9JuhuRtuIUbkDhEnc8lDf
CGGxNUPxcV6P5cqY2xe0n1e72LuwD2jZTIyE4gJYOTvbE8OTWPsthzn4OgoAuzUN
KF4CizVXTTUA/nrvZUky2DiY0cMp65P+GHPaxWICz+s+noiyyszG8XNiyr8ZaMb3
guP1P5Cekb4RCULfHEnMmzEHp/24MaGZ+K2ifVlhU1CzDeEU81Is6nX8AFyqzuSN
b8sYEZzHEzIeKBfk6gdVwE6hp8j8oU2rasd8TmodgOB+mGmvz1iPaX0MDtUaW16l
LmyDNhR9Eh4/WWgSR5ztxcJuG+fGUjURPDIM5op2+ZVJ1TS3sz6/Z/ceNDUQ8ctw
Mni4JICwr7qmc/VAQBMp8DAGUcmXnq0awqlRrVk9nl5CdIHusAOsy16ZnCSoMxsF
mg96XHJTBBVWq7n1UHZJgEqecAq0t7myteNbU0uDc4JPPO5WWnODAf9TeUfdUAql
ipTfv3876AcLAU9oOCsvuMqMkmcLt/A66Yqp7/6Opm0cv/o9ehp6mGj12DTyw4EG
LB6bKwrfixb+e6cdE4nwxabSCBtGXSbHYabfpqlpBZvXxvPZKdKeEQkstMv6W+ei
tcE6f8IvPGSn8KXZ3fo1kUoOv5+X6ia5WHBSZxILVv+AUf3wh+lM8hKlg9AMmJPY
G4j6F9wp4BK4zwxlE0470LzLHqLDW3gAQKFnSBfgenR3LD+KogzEHqeqKttmxZWz
wNBqVkJDVoqTMt55rTfQdUc4xO1/Tun+TtwvO1Eaw2Yjv+Vs80QnU+uGJ3rzxYIi
MoFeQOr0GgR4AVjmwf2mxuUpAQ0ts7XIMcu5AhcFIkiAhLZ+kB4UeHp+HGE8ZcXC
6UIFEqSpu3D90vzS55dul89Qy6dTrBGDtyg60k3o5WM2CvnqOTbi60c/t5nQfUDL
74Hg7WahmDN7FOBMiNpZtzfm0yriz87p4dZ9j4lz/InMY9YDDzBrdkywFHL4p1qH
ZXmaoq2eRZZBtH55LUJA9gpCXNtXQfiQlvoAHCl5f8kOmbgFJlDtD39uF7gGRdCZ
f1f1jlKjfw8yH1gYst7z+JtmK0bMV2h5wd08Vfpuuh+UQtrmPYHBgQikE0BralMq
8cjNYBlz7j9DU/hl7PfFDmSj+8hy3UhKN0tXuWxCLL34kwHgIr3KwNLWYHhMiAjI
olK5WoP4ycIaVvvIui8geCxc8r0bnmr+EIApTxmNv4BU/8ouTmUEup3USM2J5z0X
L6i9OkuDzJxamPHIF6Tefo/5l2d9C8dj5mOWPtf/RvuKZkavQgLMfDyS18mqQS4c
pKsKkZQS2/hH4xvy3XPx/lXoU4ETo9c4CQDUBOYsUcu/U+HbKfxFiMihw+fmRuG8
jkQpdn2H8VIjGrJLeYxbvFHUYdUyPFa0XlUXoU9uWs+TgPfAyP76VzPB/MSNfFlR
xzJ8g9h4sGs6FeViKdVlHZndx9EOGLJ0vGTUxoAWigCjA8aOJmPImDeuJ47McuEB
TizlrcN9AkkMUz5QavCjKOySRU1xbg4Xvj3YOuG+LZjtUxv+rfXeUA7xTU6/wWls
xhnaUxxIKfTH5whYS6ze0bZLGfauTdf2CNo0Fdh9pFzNX3wwiWMOL5gsyafaHXWi
/wWNHPjiLSTiGkf1V5Z9HH/Xd8UyXyNVNNGgKp2yWccylcjEQFJXJZfOuCTZwmcl
ulTB71xs82rHAKTJ70g9SkwI/8NmycXlt4rqflJrnnqsVzIxCvNrmNm8wtM53+4p
pL/V3W8pUXAQv4Nxr3X6mdFRpcsD5aL8Payu6AvBOswJGz0E65JbzonNARZY2iCY
CilOKMI8CByAS8qmhttQxdW+MLVmuX9NNCJCRAQz2aQ=
`protect END_PROTECTED
