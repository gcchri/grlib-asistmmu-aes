`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OoTT8HuL6MgibwxwTR19HgOkcqSoAkClchhMIKdCHqpyk70/DuL5D5w3zYoQAQuk
8I+RFbG+tKMSyBODqhK1eoNY0nCXlIs0MGPLocuhrLSRo1PchCdGfoW5V/oZHQ+X
FUbyLihWox7P8WB4TnNT7nQyUTr4pOdlRDnX0oXNJ8Kz1K8+VHlAw/mp9M1RSnum
mLusUklkvcN4s3gd7z88dCgAAio6CAJz10ooqrS5At10mpVBl3lSXN75VD2RkBDe
4i5AcoLMAhwuPq9lt/HMp5w3+if1KKeCRenE/OQq9tx/1QcfNTwJUdLgeU9N6VP/
mkc5Q6iTIt5qYrBX6sEhIECKqxAhqXx+ZbT8S8/9drdnh0UzZuSiWhhboC51MQoa
skYRgNoS+nnkMV7KEnGZCgpkRVRNHL1ZKocQRuP5T0UnMMvRLoRrlVeRntqEJLw6
0/39wrwtR0+E0/iyTpglciCAqFVXWy6KOdec6ntI/nc=
`protect END_PROTECTED
