`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z1paWInNoBAa0UcI9SESgVkZrXCRtqBcMWIzgiY9GnvhrDS59B3j3FY0WJOMXJwm
6VzyQSJevSDEUxwt9v3R2O2lZVXYnoiBMwMfXIVRUjSbU/plgwUvhaowC846dYLb
bS/ugqEWHAsoCYTfdyqWakzZP+Yepyyc0W8KboWnFFHSdiKQXv9PpVEUahZKefiv
No9LzrBHawr/+IaQPpt0NhEwesWVAPoA7OIxVaDhd8KD/QZA9l0U8FslFBofAVD5
d5xQwTZwP/PIo7VXcdsEpyOebQzIiA0HaM/dEjYrV8vuztDb1Yuw46E/ObRpbCQE
q7OQjSILZS/6eKKJr1AG7Mo7fld7Fgt5EDl6VwG99WcJsfJMF4c4CduYrLzQW0Oi
NfOBSFYDTeHQJuCS/Rrman+QcT1Gtnqx8rmBMoDtAqykmSqXoBOwRdv9BwHm4b/x
UTWyQGCnBLfLYcvQkLSKOezY961Jlq4/qSAu+1ZV69hZWufAuggFgUcxoCswl8sV
rc8yKeuRk31DruE1p1+HQpmJhpkuAECy3eR0w7+2k1GmZoycNPxTXUxKj0sihRaL
t89UXpmBAdIRas0cGDq6yDH/HnGW8yS9cXVt83FBiSmOcaQY7n7bOFpgUY9uP2oj
j9Mm1yx2pP1A+4u+e5qYtQ==
`protect END_PROTECTED
