`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7CXQmY1uh9kub0MOPRUEeMS6WfU0y0XXH0cthKN4TTm4x6om71f43a3+ZKO8tRDX
Q5Rq265UQSmTLsLJHsr1c2Klg813/STFmk8vERTZ9sB4rjW+Cd/3z+23ICFdjqAw
1H2Rn0Ex4HBn3oUsFYcSI6/j5H5sibRiR/FOwv2pzh7vx8lvyiZi3F2cO+cV82t4
4nLIiyJl6XkJhNIF+PdI+/ViaU0hpLA1aczS0H6CpcE9UnG/AK8r+hUgtW3LUEce
kA/vE/fDtCjSR2fx2vfQYvsA36Z8EJUMwEwmQHfnwng=
`protect END_PROTECTED
