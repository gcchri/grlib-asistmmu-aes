`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RaJR+4cTkDjBOd3uynEYGLEq0JNhjL1AGeBbKVx8a7WucQRi+UGnpFgk1AAalISU
fBxh/T6EqLIynwBkNWMQP/rwteNA+VzZAUae5KH5iwvCj2o8c10C6fUv0dxy5VSU
2nonICqbEWkIgJjPVEIb1iP9kdEhewCvQyFA9GEw/TD94hycwSpb51zxMhQ+YrFg
lVo0WgwoKKrywlpKjuPWL2+A6wsLj3JQm0axqS3e1a0b1A6DYGI/9fYaN2wYIU1T
+cnAUdQF83194CajomxLYRZYYY0Ekr5DtEj4hgVAt0w=
`protect END_PROTECTED
