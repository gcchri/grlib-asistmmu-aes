`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pXJfluBSkizbiWQ8kmb7bbaRblVH3GotE6ILM5tmTYIBmeS4YXGTWkv1iVnRnF+t
YzUCtFg8MOY2EkSfDZ2UVJxIFJ5tzOIbUSNXKyqlN0b2Jx5m+7VG0Fql8tcgb5Lg
iknjTivGxbV9PCP6rdgmA4gLfm9C4F3nvbWB11fuDowCtkarcS79Xzsi/2ADuC12
SklQgyapIOYjMZse6t+SEvUMuiQeqvgbyRMRFGjMNliPIEpXUD0PBjcqREXvAiT3
mCyVnx1cR+u5woIaCd+g7outbABUpPb/nNDSSuM9WsRzJZvrqftMhn8v7p33Dq8O
TG7C9TjQrkttDlPJ5OHIJw==
`protect END_PROTECTED
