`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N7oYOLWz8wal0Yru7va4SkwDrX3LlMLO/CConqcl5WAeoAIL+hhShXQ2hvTyIQp6
DUahUTtqRIBdnZY1/Nc1tkvrcKKmn/UBlqJJFAzA6fP1RihbmNjM8ett+Yb3539h
fGPRpLSR8UvKzo6JzzNKOmH/9/Gm1L4KZ60ydlCd4nbST34J2M21+kwj1ZysBkpb
XTDwpgqG5SnqDzW2k2038D/aWyuOBJeU5hZTB7BdK9o4+ANKe5R7OKGsCuFm/xDD
7c0RJjvxh9bRni++2q5x3Q0BUkpPVVePmA/h5Y/TJsZr5jcWAWG907T33FZeHJ0W
`protect END_PROTECTED
