`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ge91sBoQPyit5n7SG4ccoUdeBPjiJBaBtLOGcrNtr+owAAt6DJfzPHzWx0OM9a2F
G2irkR/jT4yhDi6OQv8/3eraHmz5rZtJIwMUEOeopOipYjpl1cbVWX49AUY9N9D0
ZBF7GjkADmJxlXr4zzpg8g3LOX7RqmyAhH5Abk1KeOKAYDKN6UFy21KbwO4yLEsv
YbjKm0F27Q0gK4KFpPNZEuzACXugDrimZWBHBpk1wOcfO9vgNZKPY46eFwAbYP1f
ScIbquZ5WkRt79f2A2RxpEydJ4sIo6GImQc7z95XsOoYtv0OrzIhG0Jd65DB20YS
/FibxApOapzOxZlJgroDs0FLCigwg8eTlVpFs5p8N7SvSZCqajqYDXstJzu52ukA
tKiAdnlvlmqUP85ID0G2HHTWyQSf3G7s6+PlNGLDD0V/jNn+1rnFiyYR0g2ox4Oa
xOROewbP9hrsML+jTXaSb/o/sH4wDDxmwGejiNgRtFALTGUqI4Chn4+q3J4eVMup
C6HgW7UmDTquesmRu4lDPOgVXLHvMuUqZHCgJnOZJQE2IkQ2hxQ231zLcKaagvI/
7STEv3Iq3bBWTyppAG169hUzjr8IQHc97s0UtjADsuS0VMeah4ns3JFIePgclaT5
hN/zK4t99VlEbS8u8YTs7zBoVLtOcD7fo+MykqePMuIiRb9ZQZAkt9IINSIbT7qI
exyLTHlXmt6orptF8nc82ua3NvNjGDNZm8eI0it75ACY8foV5qdNDHtQ4TVyLgTC
BD0sIOeDrWYIsPaMY6d0WwMLFH7fwNU4BbFz0O+6+AlZdp4mZAuVkN0fTfUIoxAU
7bhVudot96r9YnTOBOO1nQNEwMC8zl2IKE7eqHMx8xf33bZFyROJlwq7iyAY8L49
MdEIPUk0Jrg8ccQZY1M5XwhG+D/ORnVW4+SMWdp57dVtEW9lSP0rTaJJMVx641pO
0QQEGAoDv6Dyu6+wbGSWwqFqVC6rUhua1lWFCOeqxK0u7JXbdQbiRFlAUY+kRqwi
TBWPTh5poH5/dAT5oLrPa+eU/CHc3OQVT4LcdFCnS5WcIgfOzNDPZGNNZ2hAFPIA
qs1ZUXekx7qd55hQ3GDN18fNgbNkbIGdCCTJ8Vg1CpJTxrWsUFn1ltXhWChekANj
zJnZOECC8T8M1uFzLqgUPF04GmOhr0KjK+K/unsCQ0axLL9MgsPDLYrLz0s0lAnn
bw7K5rP0i/6ieLEuyx8xHegAxtPzAOAbLwzdowFmjQjt8hdOEeFQE8OK1cm5vOtu
Jgb0d/99GTXl2GrXId20qWQhO75YuB3O2gFgxfjgj8ltOEcytUJCu+zFJGomYGuP
GIdhB/ixMlvOhFKe9lmuM8SStkNR9prjR6tyVmLDO97eTdK2ng76H2i8gSEoO8cF
QykhXHOqcHUZvMLjSVhUh22ZIzPwIQgU5T2th5GWw2CKOw/n+qxwygsqthi5iXWM
zx6wq60E9AlknL8wsqBhfeH2G//h+V4UokdNxcdLBHWXwuZJ6KWSUhntMXOuPdWK
dVcvMifirT5nVKNFeplO217iw7ZO2zMwKPcD77Srb7MJMAgPpvHCjVJqpLiKNuGa
yvPhlk6EhIp5ghX2jAR58ev6orHJ99Wnat9ByWFbymQ2KGbFVGrfl+Sb9guwszT/
ESLg3RkfqtUU5nLYunjIVA==
`protect END_PROTECTED
