`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KBVqaljogDPc61VsEMTN1l/WxxVfLaJhYalz64YQqig+VxHt5DQOrRHKw9fWXhym
gVEvlTnTlyTqBuCmZpzCSYvf7l0CZVkWsiQyybScvCcPXmq/p9QcFJFNtJRR5Dtl
s6y9CYHqXbZ0AKfel2ewp8LcICAxgCjeIFz8Xh7b4tadeojJgPYZ7pWiSQFYtN+o
EKMhEVJowUMWukui5uwR7g/wAIsIOQxiifkare1Squ6ktBULerHEPT5cdTY7pcSB
zeU1eFfZKR+CKtGAtclE893uNfRqo0bHxH6bnDUup8gaU/rd/WaMrObn9LTMImcy
thv/3zrqfTwtZilcKA7+bGYcyO//QWc5/PSiASHQohSZoVmMCciSziU5OFzEW9+a
x69b9lNvc4Qy4wedKlHeU8JfW9GNtuncm7ZaMVtiXcEHWBgXJav703b5hB3TAD93
ohM8YaQZrQzcPsRwI+75wB9BhmDW4S+LiD4TZTtcrWdGuTz0NjQHZt4MgJ2wPm/e
gVsxnSMLldz1D9D+5BGRYkn7PY6yiTCVrridFiMIYYL4/PQTpf2I3JDbfCKuGE/Q
rhwNRaG7/aY8FFrb4U67fr31f4LuZMNyWokKBv2GUsF/6tkj3sTjP1+DjT+EEfKq
sGSIjALS54vciYwjVdhuX3qRx3P4SbqS9V3Jlvcosjvjl8WC92gE4rKhxVIqVHVF
f2X7AIbFKbZcTuY9GjWwPMRcmch24v9/PxjGQLIzkTTwNFmypb0OzrHkYnJx8WGa
u23ZMhqfGNqKWUkRNofLO1pkJ0aoP3a9zzrggcO1pbuUyejYuiIUENlA9NOrrZ1J
HhfS4ZL+xuCR3IBsIzVKJWy0KvJP0Qta7eh2PtRZiLhaE2zEv1BJ1gH1YLNw1N6L
luw2YQiu+DkU8u0PhFGfqGjWjle5MDnSTOeSBAaMLygAAWeuQp1DUpCPJolQpO05
JUePtJtISMqDRrAh8FzbIag7dVSO8ofGd/dq+FynXqt3HqBLlxKm8cdBFPQfIdZR
kEDtVm0pMaWrwGzZVCNeFFO/LbkRa0DYd+DL7lcHVPQrbSawmivne5pJGBq4j/D8
u/9rASTx8PAXpqK7k03kJJa3IU2zm0KD8vhmCgOEN3cb684fXRGvOfxbbWd22nFo
co/Kqxwrs/rrpnhTTKEiTeQh7Tur2op/tw5HfOoCTtXxBILm/qWE5CGMWziiZvNm
vf/2TQ4QwY3jeDXH2ol4LRwMjS8W7iKJjlRY6cSPBdYcf9aKMHAQFirwkdK/QCJZ
74qaJn5kMrU/IS9WyVgcg6+mF9y+kSzl2esOad+tQrlYyHQd0wD+ggwy5QhP76cp
QFj9He1Psv+x3OZJ0KT8V3vEM8cc0ac9PtOB2+PObxf2Lb2iwkkw08ihQxbKI9Mw
8hgIlKWuyYfOGnBrDXWnnt91hoOQ4im4dNh9pZBuMjY3tcABGD6wiwydK4pjah9s
w8ke2vHadc/2P33xH9hOdqLKX1sQeVI0KtVqT2+1gRX4rH9g8Y9g8ULa+6tRFLfK
dt1gQ/gjXOsyXgxE64GrwSB2Mya84rp6evjnBkj0rj4hYNF6GM+TL+hxXXbY0/2n
a50lDhmwnm+L1mvW6z8UaV8w1LjN5giHq957jqAU5AjHz6Wt3IDP3jc/7GeACBKU
2Dq/8vyvR9EKi/RMgpsq/jOvUss2QznEzsCL8wFkNQBUH+vtwcTHbntAvJ6vsnB+
`protect END_PROTECTED
