`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rchSu1srDZJcGmhO8Q+6YJm8lo9Cz5E/jggBybMKJnEfnVgbtXmmi4aV0JADZJr1
qGfrGZ/+GKxeOAXtJu9fNIzBJ5zGDV3aQT9/q6uFMrX9ipyTNJVtTKmTBbOD3GEO
cNHwRzUf6ccQ7zQor+NhSaVF6kU3KR/Efkn7lznl2oRgQmSOcnxONRIgNC9UteoP
3V7Mim3rltvj8aQw9NEhCXTK5YFhYqJt981Ph3jXP+OoUb3Mr4f0opCL2P44Q5pF
Sjl0cK64dsI9rW/JSGt2yUsnmvt13ivPmXvY6BqJHH07upg285huefemFtHTMlrj
m6hknJORqDu1ZyGWZo03wjho66mpgIigMC4BJwQvTofU/5YkzyevMsl4gHKkAjal
P0PnmwGwrmUsRkoXNwRCtz1+ofX33i1Nronwqftd9eBnctQvpTvVy5bS2yEkERp/
pMvqnBxLK9YOsjl7NZSa3YN8vxjlcjKem0j4WyFvQ5jx44bz3m/rrtltLYWjBeaz
hOx3hXbo6FPRNP6ZKmQspRop85Pgd/DXK9G2N2j0BCf1HIA3/YPuBwfxjxZWXrgl
RWU5xGCPh7U7ESHiffib1Rz8UNwu0K1PujfFhBJB3XsGwVOe1CPium7gm4umQgf1
++YMPcwdHs0yUOHWcbgqoTf6BVwiQoN5f8rdVdY4GaxEpL1HsTNHaKFf0ciivO3L
a3EumhdChjfkaIUpKJkeDzk1XrsA2hEtUUpg37+8zraNU3i/1swLolH8EpmzD0X6
rVnQbvLszFX6T/P0brpgc5+QDeenb8W3FaaRVHBkSxnTIrNS/DmSUXyMH9E2BEUt
f7N0BSyEfLxZnwf01iDxPuwuyQYm95XQRk0+l53jP8FpjW8YDX02a9OcIMv629zB
RvX538jvSOXTSxl3v0aGCzeb4UnTSddsM+25/durBCF7BCtm4pLP39SI5F2RnK31
vZn0j460yu6TX+xl/3uMIofqnyop9/LRta4PnmFuizE0uWQSQ9GYWHO1y5vJyapZ
KX5fNJ7m4hKzrlFFbW9xs4jE7BO+q155ea0hW945Ha8BYxASSTSAsLsE3CKw15ay
zfbSPflpPGM3P42I/dS6Jg==
`protect END_PROTECTED
