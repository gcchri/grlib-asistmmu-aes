`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dCmJGkXjgAJuSxwg08FZ7TBf8vA+VEVYG5rQ8wLOenFmkDGNPbbuiZMXh7sxRtfz
1a2kmqyJYvtu7ez2P3bcrio4iNHTjj2BWl9de3ScSIRtrUqXLxvSS02IYluieHto
TcmQ+fCeTpnVm0h8x1NzwRQultYu1ymcdRwSDzxMikXyzW4NT1Zh6jCe9Q66PT/w
OoM5hgLdLz2O7ixZsUSHJnjK8G8J3jIo1xT1LYZymcwRSfYh2kq61xicC793Z8js
dC4BjN/G6rra7lrCDClmZjeEjdR0jJ+rvWH3A4KVrWCTM2YRIfJ+1onTluY6yg56
linrJCRkpBG4p2iSEH0kBDS31L2Mv2gMfUEZAIfgaWkVMf4PqqVua9YXu9Uc+WkW
YMhNxqFYtA0K+P2J95trRdyIKLHjn/G2KiagNOoatfAdsgK3dKAEfGgu/Ww3UVTN
E2af1CvXcUm44qF91JJgaW/eXW6/zNk/qk+1/Doxne7ZMJ6CSXWONLjt94MParIG
cN56V19t24qTdVFWDhtaUVwd3r0N5Px/F/tyGpkD11Kim5aGKs62ZpHFi/Pre1SB
K1VE+uHOOrmJgmEjTp9mCbpKhu3b8d0FGZT0Zq+QtRl4ItvcYQJLzGVk6Wntcaee
d8l579GtHrgqYm5vsh/tfBN3JDXej244hNcfDq0GTZPwj6/Zd6AQkmJ2NwuSalWs
tMU9HRDyesrs1RAhk4eAo7XbEUthD6VrXmgW/uRYcV6bFbjcEjFP1HBETHeCimbC
wkVMm1FQCQkv1wCLInnbmCvhnJp9x+5wn+/akCquCXj+47vrM3B2QVEjsRimpn6h
SBgH3orHG8QQyOfHYoiYj40aojeWwSsuQB7lNAX2JeDoHMS9F5JGeAt6NzPN4X2Z
DbEDvcboAV3f5v+f2QW9i5nYV6bXKexod9pTAuUypCdRahhle/ny7irhOM2A0rCT
O/L62o0TCE6KYwp59L+gIFEgNGr5DD/6/5NOq23KMIdc4ndnW3SH0ciZVVh+aVOG
z8nseHgl57+m7alIlPobkzkj8gFWuneCY2+i2rBxHpjyyBrkh6V6i/YyI7DWBNWK
s/8tgZo67AQskVNfL+GiL/+TTweitteJ7nHxK0AzMGoVWgU985Fk71sCGPA0J4ab
daSh0otYimq07tJ9sTQZWOjIQq1OPTwrT2pZ6CwOLh4+Owu8HE8Vvl2Ma1rGHwVg
8l5NBfXdi4J63SqmIgARghEndtQCuFxDxhwr701JunXEp9A2o1aITxzOK8J+8Z33
`protect END_PROTECTED
