`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xfufwV4amFNevMsvs6yNYXIzRXFfVsJaDVKk8uJDkZCGTXYreQHwSMjM9kDhO9hS
HOykAF16kDIIOEmxs7tl+St22FV9APkdiLdmJ0LGwp0m41MaKOxGlQhv6tiLCgHe
aJMwI/9KNUOY6s4hf2sVhPyx+cqumfBa+POnnMYgT19CvGIsAYMYuXATtdPhGCz3
IUBZwpdvtAEEvLJx5Ou3JzGXEwKp3i19JUavTyXTPE8H68Nq5xx/JX5Oqd95kRP0
OQxvDQnUPkmakWxwuG8HQ4O4MdyOMzvK8RkfZFwVf2tKZKuWCX2kcULXVJ+BEdVS
JLRBkkpTbSHcgWGsl+XbKOa9yV652Wzd7sBOVVmWQFwMwO23f6zR8yiBCUUi/6kY
LwJ2aUNu5QsdujfqZYYRUEmM4kcGzOGnJWbjq3URCUB1KH0r41H50JCEwMCDhiEr
Gac+MbLA2ZVHVK0MY2pXkrZOPDEqTMckKnYjfgPZfI18nVu0NGPtoWdrXGPvYUpU
8oWhPOEhX2TRJWGj5xcTDhUvWv35/ke840Vnrsg9vhgMe1xrVDPkpTdo9PsiIFv6
BRHF/mkAvxYxtFbv4YnyEPwDK9bLQchyqrYopCO/tgREnPqMVljFbJKpZuYtbW6Q
WpWfrerESho/Ux+6GHd7uKLAHTC+qlefjm+BiuG4Do5kQnhtHxTBgqsJRpf4TUvX
bJZjld/I9Xe2TWa52PIzqKHq0KRdS+kU/h6P0nMTskte5tQ6Yx3dwyo1jzzgxTPX
b4+8dhzAeclPLTs84WOv3gVVzbaPqYKd92nE52rDDPCt378JbhqQvYxFhpUal2qa
VWq9xHekQMoYRKTvOnLB8FTY2RQMwdo3hCSxOun6Pv9SMiwbQoMllJKlp+Dvb2No
+k0ivTxPGTygprcOZzNQWCRCUMTYHWB7Pvw6oHAAU/qQ10DPvUos2ZnxLR3H1jKQ
9BRuAIoNbLl5SLrecSDPeamUhn78RkaGtbbY1BAFfLfbuUzeFQiPbRfa7XPFXoZE
CWIaY/SyhM5nZA7ZPsb6tQ==
`protect END_PROTECTED
