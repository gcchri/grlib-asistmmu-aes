`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0p2BFQbt07qcq1ymu/jBqTxbjaTiFbEX1tKhjNBmx14QmisDT49gPMV5ms9yv15d
Cw61r1P6zoubA6994uEYDWHf1/K8GAyDfVX2BABom/9l2iRRHxZjeBpUQN9P+Jiw
oGi8YQh+7TQ136pTKdSdnw2XWOQQ0fS1yAwyhNjhXZxS27iCxKCpf8Nh22wfZXF6
18zzpwhsDt17OMchMspeJN4pkw55NNap65Y02V6LMXOFLG2VPwzTlZwBY3L5GQ0u
uAKMDZ76W+jSbQyn350OgcrPXTnXfEIrGZskMiMmSncNa33bsrTCzAdtDh4BK9N+
BxL76+BF7M8pXnAIagUHHNEFsiiDQ6OBjp8Awjs14t+i64qsgmy9wuFbT5LztGpz
nl3Q631rvjw6xI6+K5ONMPa9EFZsoB+eyx1zfFcdt+KSQVJcx3GMIcdWL+dPRZo9
nML2LlYFgIZZ+69SuBBhUMMFtIIPfsMAfqwhCv4IOoU52aCRobDVUvwIQV+2KoZL
KI64DCK+DYmkwEF5KMF1puJ/ZlTAJIn3hkuIGE5A3F9kgf9cKLdRVTEO5Zg7anjX
U2lQYAmhlD2pUJUetu8Tx1rL/anvAeE/e98sQy7lQaWtFg7TbhjoLKMSAto/Rk8h
L7rxGWle4bKYagw0I04v9oAoRLdPPoanXdEuIbbwiW9Q5/6qQQmDfQKM5KSAMGtu
DU6b0qLaugaNQFn8bjcLVIHBkUzD3wNs29wjYth3k2w=
`protect END_PROTECTED
