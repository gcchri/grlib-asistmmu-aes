`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lmFcbGjO1GtiM1zBtSTb6SHINgsKl31eysU9OHULtnfDUoirJtLBpKqVSAeJqhGD
NMnS1VkYZohlOykbDfrXf6Q1p0G8I5ezN+oi0ayuCqH3eO65IpLtWgfPMwoUw9B1
6QulsM/x3Sk9keaDmV0dT47eAAVZ+Vo213qsJCJ6eSJTjdnWF9mEl3qxObDH+/lq
qHWTG1oa+5bF1fYVrjDH1Wjj76GnmHKZHuIhQL9+JYZGhG3rt5ArcOkFFyDjpHJj
MiFQ/0ninwQlh6WI0XjPAqZkaqGcTK1P7VTmV6t05NQNGoDVJnBSNI1LyqQfkYqW
pEsfsUlGTa2VL++L5TKKwU0ksHY5d7svphTlT1rZS2XzUXc+scm/hmudlIJ5kVWW
Sjrue+nzV+q/eviwoK5Rqik5dZTlFQ/v7B7VUuVOn+tBkCytVO9ohOlAs2ApN6Ar
4sFqf37vSFXBZJG9MfyEOish4fssneeH2ZgJrdLsrlk1EUW20pPem9X00I+4zglE
v1MtATfR59Pz7HIcj9Ct1b0RqNfoHYaPKtT8OWF1KIffbtWPe+JE6OpFcTDvyeTv
PQ5joh7G2ZUe+QyF2XWpUSDNVM40EzBf6Ng5sabUHQJM4l8YbDgO+LHr3cGatzZX
PixumGj6vNw2hTq5ubchSArPQwlYbOJ17sAaHjip9HrW4i3qcfKXnCuHnFoAiIMN
KrT7Z+0uKYa0sZvGqN4W2f3xBa2io60BPTZZwo6BpypOMWwsWSz/9xURiNnbbrXB
5UtEwwdMBg1CTYCFP6Dr/e7xGsLcCMWGcCJDc+HLMmADFbP7+3R48ATHD4ORZkHL
nr9jjiHcC00xzYndXM+bV1AnZaaln5iVV0FWAqULhlIUG2oCFl7Nr3MgELfITlqS
BEpBuyZKsJiuKT3VuDnKb75Ss2I/JNoRHdrSUwFJ80QiNtWkT/a9qZc3fCO/zUYG
fdcFY5GFYrg9R+v0RRyfFuseuxwCpvRXJWYXeZK5VNqRi3f6RwVijXz72e5Tadoh
Fz/Ccmsklb0QrmBBaM5tLLUCPjboa9i6IC0oS5gG+xdZM6a7q3cnBg8hrY/vcWEl
diEJLcqyq80GL3WK+fGIgGD2jZIaPosVyvzzcDTFO/xg7duRoCtBkY2ZbVVvroW5
DlMh8k7RTwVwFotV884WELisFpXZTr5ZjcRBSPSPn0e0Ilhw/33tXJd1WLXlgJjt
skMEuServbgzyYFH9uvgq/RxWybTxMYdk2K/gOcuCoEwDvbyt0rfuuV4ECqiV/sU
3rA11JA5Mb3JCzmtp7hyEDi/4m5+N0L71aaxELrWX9diZwzleHcQa1YiviRvpD+v
ArR0vwENu3ilCljIKicDrt9i97YZkUjTAYJ7oK6tNWNGSKKPuTz7ncBaXK+5f697
BA/Tn869vbVzBquwzFKjXphOYB2fRmS4D9Ki9+IBOop6Y+pJBcLJvGtMBj2ON+/N
jcRbK0V4JUXH13eWd87U3clx+QJSYwMhJHRqCwJXwdNENhR6D4ctBCUJeS6Xijzr
m87bWKRZjn80vCJS6oIdsyeDV8Mi+/hK6YtQ6sVwCaQGk5yuXI850N3fv3vhCtNM
zlW12Dkdyifi1FHA10BmcZbYcziE+AdKACdhn4UHTWLxKPVlIau3t4x2poCR2Z4j
nkoGDKHGDG4XIW0F6rY/QoPOV/8czb0dM7T+GtK1f51sLnVXaG72rV8I17nMhlZQ
fuAw7chU+1DFKW01ruVYQXjb5qloOUYE4V2gXtf4mvdcEsUhk4ppfcoFP+u8L2M9
/AVJpz0jQ3n8ZuHtfVner9tMqallKcAor30/2taLyHU3cNyNTaHjj67ZLcDF5aXM
oJlyB+9INW0v7NJVJ/iVcWaDBnb+a92/X5SgBAHmkbTNkIYmxSJ+oRoClPoY3AB7
Xtt5FV6z7HylI+9/8wK2g+HGytriaZ9gg4RMstnAtmShhME5CQvOUWVtLnu28gt9
wJ3Ttp+6+I0e77ZRcXBgpqjA5U8Z9n6agMMRpMG0LCgZ++ci3AcM1pZCDkQIthxJ
4Dg+hRuXiBWfpC9mb8ilSuFFlPRBhsELYXm9OhPWi6cHyhQLGDgKq07falAfmUTx
TFxlyDd/htfzbsAwxbqlVEM9av/LLvAu9mJH1DVKNehvkS+KoM4VepDxY/PEUIlg
rWLs9vH/ABLpqoeRuG5rV8qMxvVdTbDYUYc4wrc6mzHjMDUe7b+QSBrdmGD21WEn
zgBISFmkT76sL8SFj3W542UAI60znvaj5/ahKLSCjym2as0oaiGjQNyRsfRW74ac
cjs1ShazAbJn5erRMzr1MLJzNFy6ymcdu03/WBryVqKwdPmf8Agd18uj8JjLturz
7Z4lMtghXpbnvWBNhIjQxnFbfwB33ZDo5TFC7fGK+l/2a3E+B9Auf6k1Tq0U+lvz
x3RKrPyMZOsc44CTcF9h83xHQDv4Nb/2LXCR+/ermYhZ8mRMrRWEF/DJPy7zVoYe
k9R71AqHKuBXuaOxiAGNWLiadIm1PqE6lzZehu/agmJl4WHOlh4GVwYQb/d9N5P3
ku3BcuTvoVxrsjfBQlw/zee7VYag09fERxf2Ip+jD1Urnj8QuITB9jgI7yDAguH2
Ej9Ja3L/tSbKOFsCEN0L8TJxl00GKVrtjgXv4ZWpBgiexkyur35xm5o+Jf23vAI/
OIOEJrZMjay7w1CFEs5xWLoCB1qLIb+O6s6SKhLUw915RyXtF5tcJBBEmiPtuoHJ
M8XXJXzSvEFTfYIGb2pHXVMN4FOL7pCCH3zcGXpEeX5WGJK2qWAXyNzQarZljM2i
Bp8HVnQNDQc31TB90gw9GveW2NSXamZaeb3JJ3veNz9PCDmRqRb6JH2EMq9N8CDN
RtBjwdx2q0XvoVOYcjQJ9hb1UL+Lbn+heALcazMNwavlaPBITlAodfJ8sgjWa5Tx
g7XOGsQfUiukGgoG7ezz9gCEKw8Zf6zT36y3uFzyW7EpLCbPAEo8ahfvXxUwcuMg
0fqSrzvsuoLZsMJjBOckvlIODMH7moDT/zDo4vKYg5XGS7nSpGoKON/KlBx2arbN
GgifklFBk/ujCyaWWTaBn9QemiD9p2Eia8718Jt+ddbc8cFNMPF+j4ExOfrMq6/Y
Nfk5uRjbcXR+5/HZAvcF3GSiWSMirppWe45VG7+xRIHXGtLF19Kji+MFcHBPBcRx
il0hGZ6ABXeW0jiGTPRIJQ7zVzda7UaVVrSiNtDXQp8pN9ZcKQyFFjfWeh/YGMtu
5Uq6Ypm3Ot1nIfQxWbf+QBge1FPbXQh+/Bo6D8p1nRTbn9+SFAQDAtcFzsNsaML6
BxzdahfIXX5g5t9rwjmMUGm+OefDHbq5vIGT1b5bt8eiS8ZnyRg/oAeXvZdh4N+q
LqaqQizKUmGzJOZBqe6UWcb3e5R1rW3EOC+pxpjq5Isx3UHJ8Q+LaJZvpOV1rjjQ
2BJpEAi83X4ZSt6dCfME4XxXt7O/wLdBbR+D5+pw5Cmdovf1Weum+9EWD7ZBZ2yV
Fs/GI353tiNiYCmfDxwsJP9gL0vkrE0buerYf7BOZaofRIbUCQEB0qC/ZN+kll9E
x2vtwkd8lSjBDH3xUEGvT7fXbEbIZu/nq+G0tisWdcT6YcBapXgTwupvSz9tG8RT
ReF03nK5yQH94aCCJGnLM98324JjAZQjzmPUzYfk4BqQYhuaD6TN4C8G+Z8evKrm
vs5GXh3LfJp9iPLkR4sqrqxjVhNp5D0+meSbJ9TS5g/YYIVmQWEljnJtlgeqKKrX
JW8YsnYtUqq6fGBe0u5xigwrdRlIltjl75o/FOKunO8UM49ZpwJMH6Dts4a+tc0z
m2aTWB9yoNbQE9ZpaRAcrS0ISiditNjbSdSkzBvy+IYMWxlu3N3eoLum3aFZRL3g
t4YLBCHVpMFwbz4QFWlUQCBJI0spCyJq8qqem+eb+24WcgHhPGPB+r+hAu6ZGedz
x1l/0gyxUUwldpDMtNm9+lZOsBcsS2ibPi7UlXbm28TRXRT0dwTTNikMKi+GqJhB
IxQ7AXOwAf8ieocDfXAriWTJZkHBXHNZutCTq00Z5AJntU1OmwlIr928nwb5B00/
KHyq6AAtZcHFWP3+/46FaZFecuX9ktL2IzcJqRqF6y0hdKFAMqxSZF+LELB7eGcf
UBHxeA6ZvNcSDk+9Xudr7xIAAIPKNnPtqUgtihHRkWpRUdC8l4uqTS8D3lRFB6W4
WEWa85yP1tlCc+39z/DphJCFtdBTJDs7IrvTYAqWyMAN8lOJMYtczz4gjGONwK7A
gD98hZTD1hkSB2xP94XnXhS+wbFYI83OywNz7YQpF+X+er9b+c3Oa/z8khkMFWEu
Tgkqkb9QVQ4+1mLN7QetkGQ+mBAf9CPGU5xGVcncyCxmNqzZEffBX9UBRGuIw/sk
aYvVICBw8UIKs5TzqymZvVWPg7T6/zpMPiBHMrXJOBPee63nwNKJRJ2ArvcJUdyb
OMGUCLj9gf7IOHxmoSZ/XAJgVgw1Z2KJEFftXkmXXDX239+mo43R7u/ecoJFtAww
3aH19U5LCnUG/ttnc4A6V7ApPlGGJOhJohXxA3bSM0s0pJ8WH4/ARFMJ6ks2D0Li
lu27t6lyq/omiKwvial1C50j169s7NiGuwIn4WEy372RkMie3RKzppnPQnfA/+Rh
UNx2EoDUuUrDyd0mYGAyfpVTOV8TIXAOV7SVDMQHZRz2cCksM0WibxA8V/YbyHXu
fcP4wduyu6KlLpaMJsUf+NeHDKALxZ3OEpBcYzPVmSHIr2PR7dtuiyhyGn8RJ1Wd
Tl5uEWN9lwkbV9oyRH3CeXpsnLRVbb2tiab4IBuESRZ36aWvFelHyfj+q5RI0Qc8
ZVcSgvXgXCqzztPdIn+eqqKzuLK9rlTz6Du1EDLbQ+cNVkFoHxB9UVjU2rLri+Sv
QnS1g4F4d9hKDpBbm2xejCTRwOYeqMlK0ZSUaj9ztR6gd2qAffGaj3S2RkteVRvH
0zfUWyMaQIufvLMlglZj7xnkz7+73hBnWG0qj9CWsfsY5Hcdqg21vzb4I8sqFONC
NacshXqaDdrCT4Pgd6oYG93zlhjgqQZCK0M5FsSYYFUMDOnrAWlIBA2ZMDLSXNla
4G91Ph7SkFjs2n6kYJNL9CtmfkTCwmWRpP823vf/sMuhuK60+kPLBViT1tXuB6OJ
o89clvtg89evNjpE1IKtovORNLajo7I5twvBDtCAQW0DLcHaOD4SY9diVZS7R4af
zKg8aCxfOsgVw3CmXR4W8lp084a+UvVqv2IPQ6tLGRRzOSTMP8QBWVmPIkvR/jav
GOHoBz9GOJ5TuiYSxxQ/wamyzyFwEQfTEZF3eOy/AYs0SF77BsRyph9pxWqYrDjZ
siA5X24TeQjWI+S5jIo1A6AuM9MwA45V28DAnIaSAdXfeO5E7gfWZ5fBee1CNXPA
v9WpwPRr8nv6jcQMS5WCCkHqaHk4Ea/wJ7bYAcnwLGcX01My3GC8MdB4SGxvcwh4
xZcpWKzwB4mYE/GFX45J6wMX+t9CjJHHHWEYWWm+sJNJYfnNZqGAzo7HveO8EpOd
nYKcAB0RkuCkmSI11Ig1XA5ejr1YdUe1tMB3Fa1Biw5cZJdpUzv4InTV9fy1pU84
HJJz2MDYiMhoPITzsM9o58PcbejnimKnvkPJ5yHXDe+9WaN0xdjU48e6YNpfiUu+
2O5ptmyW37DLLNwyNky0tRtAaC+FUiVTLQg9cQJPN/Lr3DYnDohgz7cMS4FIGLOo
6MxnCOmASgbcbbZiki5EvPaeG3xoxisU75SjO10ywWUgCbunEpvLvqJ6JuMs1zzJ
qyUNZyMkpKm/nvk/kIN6oYACKotmu695gPxgWKmsjVWGVDkZyG0PCkhKP6k83W03
NJY2e1knPiolK7dqBONbMg/J6RD1ao5rYRTldPyjN3opgyF9LFcBypj5r3qGAZaz
46i7Pc/U95a1nGsjLGEiMRmoMzdcz3bV24CWPbNogpT0bbdyoB2pY3+J7ewwAjHy
SZcJaUoFzAtmQttFpsdcAKRb4XlL/4YwA/wt2zuiXg+DUC1TesofGTcTWrRShQFZ
uzaYvuGz1aeXaWMevLbbPu0VbWGhgKojMjXgPklfZ82KMG9H89OGuD/HYnrF3lVE
i6jIE9E+Ag2c06iKlDhW7rPsLFjKMtVlRNY8W4Jh4Vp/Ig20Z84xWRYeLIb7DuRE
xVIOJh1gAovzcPw/12VXmGyo4mkcfRUgKR8CHDcf4QS8wk95Iy0QNgugS3yaTE5V
RrmK14ZncZl44U1eeXPDoMrZXFma1ri6kM6IlSZH4JXlnl0HDDwu+cXF/cSMIfPP
XCeFLMBxWh1RniahZ2m24KlRBoB+cE7J15YZh8p1GTBGTT8n+glCwdzJ3ZvTPf18
z9xrL1t8/3RgVzdqdx7/MZH2tZxL0Kk0vh9BbS3oLLVOR9ciHm1eE33YKQobYovU
Sg6Vo0vdQ9pIexL5t5y1Gs3iYC6ProDtID29FGo1cFZOEZLCjFR1aHv0WjSq8/D1
g+UEgzqNVleuimwXRpYvMNKn1bg+VqLA7YT9tf0DeQSc1cX/TfZKAN3hmgn9I69s
RiDwfZXkiD9cRIqS3gwNiZXxlx2yBsAtBihxppDTHx761mlgAeH0LUyjYbBcXio6
NVpsrubTVID169xz+lx7JrYWZVEdwa4Vc8n3EOnD+/PJhdBJ1IqOw+jLbq7NS3Yu
IyiNsubYEPSlp0WIPpzf1FGitPgTFHmmX/i1wplUbUolZu35FxFQwMKjtUGTd1BB
ayd4p33V7GGgXLoCSkp+vrl/GfO72Wvn+ShZE2V1uSGBE0IVxZ3i5GsSPLih2Xl1
NSoDFdpVx/a4ALGIixHMm0wG6S8r6t+j5nHO+04DldNroXypoWB994lOMXcPrETO
gf7nsJDE8keUZv8+HoOQTMsq1PPjGBn4CNgmWNowAY07aURc0zALvJu5GQfJT56Y
BqSn8DHzqhFkyWfNGNpF4EVFZLsXeLtCgHX+NKpU3MOBeORqP5+0IYpmhpXQrNb3
nhInrwQ2rhlrPe+THBx2LQto3yFmK93xXeaVqyDud4pdnUa/z2N0VXhX5q2O6Csi
H+SMQUgP/qsdj84Kn+kMhYx7DwtDO91pbKfnTIfzaKpNZ4PMrv1nAf9sJnzuQVPC
Z4g6mgTNDvu2qkEu7SplYybX4f5sY/gojOm8C+5lK2pEOb8k2QzSVa26uioZ6+ej
uStteSRz9lHMWdUHnerj3XaBBa4bXROilREmssXN0aRDyZ2fYkvOuG7Rw9GGnINj
6/4xAbm590cP+zKZDmNoBOw9DAmFVsa9+am+q9LGUftRGkKvGBQqjR2cwmRmmek0
YlA4r+yE3JB3fiJrp5OXx98p+Gc/PGEwgOyaEnMFTiATV6iisVPp3MX/NiTGKs+N
YrTgUUD10Dq0RK8ewXTU4UOAExqXNvJOhlPF4w19iJhcNTBJ3ZhMP0AS8coq+HI3
uwuqERXipZY0y1i8U2JHWd3qbtAmPuVOXGNEPbUSeT5XqlZTRzmoxCclu/Hil9o4
aUcP2rAID29peaf7rB2SBzXUsyVW01U71n1Ss+DIYvPfr4CMnXzC6JzZg5dtDB70
5+t4iIMY8mFHoS97HoT4z6IiI5/a0+HkyQNSnrNX9UVetulzqct7knGyJedTrQCY
MCJx069h+PXNC3GBbEpuYBqCc+bCLmGILT/qKZMCa1FghrSCttYd1u/R61efiNpx
GJaGUYf59ed8XISBLtvIVIDnru13cBviq1bTkikB+j45oyfuOyDkfIj6OA2gHtaS
2/qPcuu6YT7uwuZx/eHr1Y8IXqXL2A2BqkAq0KZQgD08mdIXbw48bcbKuqEhkSde
mKJsWTyneIq89uTNuWtEtwQDJ1oM7RQDFkq8HW5/G6z0xomWasrtGstYEJMsOIkH
GggbyDTesjFLrqK8e/CCag2ozYgWy42WC3vSfK7eTH7XnF2PTaUovquJEqRMYmUI
ufaJBkVJxCrIhS84Crw4XDZon7lY+NtQ76xjs1dehoO1uPON5GoKo1OwHBoRT6HY
j1jQOEyBUbHK5xrONAfbsruxEpecmqoV2MBsUWDTdOgf27fNjCKvhJlX05RriArX
Ode32RL8AN4Y7OEEqmAVf0P7G9c3IuMnecDNBQTZgQxOgvvoYwoOh4CBsxiq7YU9
M1bRC6n1Sort8d231R5+wNF56TdThZbGjlMTXK5TQ4HsRm4jUKgzorZ9veN1Rgxc
J+ZUlm3VDi5wlu+piMF5r3pDRE512q8GOTJNtaKH2VF3WdUWU5SiiDWSEQVXbpNz
3GARn5JVo/ElHpN95w+gqb3R2+mRugM4kUUGmyJcYlofggLzqlJJBCt9t43+g/NK
Tb0KWLbJExJC9F1VENvj6tXgeyEOLm6DKnUQhmEJtjA8ZmOKXC2kyuhXgzjwSyiB
kWB4h435IDQCgaYfmIiYd0yUAWna/bszXgu74pziPxsSoUT7da1NbvZg4+3alWob
taly/ubahw3J5bfXOJumAxQA7rXjRdaGewtNDzySY7yXIjiLnh7uNGq4+uYArUGR
FrEL8whDxjm2q4LamuftTT0fEeseKUAvzYDe5ih7FWpxH1+vuvRRRRpIZk5ZVdTe
ho6KTQ+Qe30/zZQSTZ60ae3rUdqL7LZ9s2sHDfdARUcA1tVSacVJS88GepAxMDpR
UcjVFQpLLX/UblvmDHsFs8XgkAy5vHYNLS+W9uz6y68rlTaaJFAcUq4NmSAeavdR
cgeBdSAem1C7BedhN8+cqWQ/+uUthfFLgnd48CcpFc175ftDUcEtZRCghtlkM1R2
n2pbzG+aC0QGZTDnon2jrnrIj0bX4tAr5apV7ONZPAxlVx98xQXN84Q+d7XEo23m
/Y1nZJViBk7SAYoO0rwQ0QCi+rcvKwlJBd3AxpfFAXZRW+FVfT0S0zz8bOlt0mCX
54IB/mAM8GOQtc8XXg44GGx79RIeWT46ktSjgHsqRRlHVLla7iSB31FJYN1X3QBN
MZo+jsMQuANfCl7oPpz6iRVaUVFePYwDCKhLENboFpgNtBytLd4l8d6GUntBAHzI
LCR6EDCuxfG5KfmYZ/Joi8ntwibnsZOLIgVIflH54ezJzyccQJ4Viby/TpYaUrKN
1opPqmb6fbj9NpOeOuCyUaqpa0ipCHP4PEwEWdXJT5RSxI/HW/TGBxHvfFbKiCB+
F6rOPmpKikau1Bx70CuIuke9lexKUDzmngHKH5TGkXoSoLZS4YSMC4Y6Bz615CaZ
+TOyTY0Kk4dBrxLtcA4vUTNIwUiKryvvIFFfbMTk10wd0MDIpTuxTTvfjPnKraYS
b+5G1ZF7xYZk3BvuJy3lztqx5TU0MKxsfmK5G7tmCtGQwkj8uD5At8o9o9SYHC7T
zHf9X4QiWRd2Yr9ttZlORP5P4NDl3sxgtlWZ4be2XMcPfxwwSSJNNXM59WQzwxiA
5UPEPqEM0eJ2LBz1iysAd78cQBXo2vSZs7Wjyfv4fXXM4X2nlwr6dfhnqlKiW5RO
arOfr53ZWR492QBLv1b7Nd49fmk5a5I3Z+oeAoG6WpPLg3Ee/dYqx8e2YyF1GQQG
pUiNEk5RMBzEF+eVYvhINlqHY3WBknP7mS/P0IEHhwm45oAHrNqtLBXeXDuoO1GZ
ukF/6erlCbqccqgIK0OUVgozgw9NRvebGiML6/vNTBSNHXBFDiq4Gi+Nl16jt5hz
QR7TLKmfEcpOOIMw3JAfX5NsBxWunPZEp+dfGX0w365R+Cc/cWdn7hr9dCkppQ1M
F87HtC/RU6BMt0NSqUv0/YfaDjGwnjNQ7Dh6LzM9NbxjmMHiKJ22kb+loYiLJonE
JBrFtYlTZ55hr7BYk2PA9OB8Vs4vjVUwkdSi4obXnm4rvpnX6h4210neX5gc4reW
F8acD3QfqTy6Y6RmX74S96oXj8C/42+Puvil66X24r4onwbQuTksySxnj6vn5WeF
MWA4nwWlhCBFHmcwjw4N9gdd4ECLjZxojiRZremlnXDDSRk3FSbayU5TOseWXBEV
CDspSYmd3ltqbvvP/WY0kngPUsDZiNZbS/7ORefnGOErkhuzfGN2xQC4+pNmWQIx
fH1igga+yYPGD8FI1K/bhGlWJP4+4hI7HFXEeQUMwqA3Uxq8oAws9rVIXzC7fXpF
xb4FvaYkIzbmFAxFQ4PbNlexHawNPVNxM7Ivhw5XBSNAfW0GEyMZml4a3J4CUWNP
UZuWQmlrRVllwMZQN+nqP2RucybyfnYXxrtV07mnfxIpEWa0l5N9oTa+gnO/+kjK
ane0uWkQyVilGWV8TKYNudnmi/DxFcAQVrqdUIRoKkpz5kiIKi51UF+L52+zFrAd
LCD9UmfPI3crigg2IsBnS+NM7fAEFvduXMq0CsgA/y52zWVUe8a49vvX+jBCEBd1
ZNSh4z3VRzRbm8GLWc4FrS0OycRQTvvNP5C+Y+tICF+Qk7SU+gLfP25dp0z1zCZk
UUtdl5bcben/mwneXRcvCH/dsNsETJMD/I0Vbceb4JIVuu4qoZaOLrfe8vkSKeFR
Mllq8ZC0vMMxk977nOVXGXl8e/gxhrmKvdZxeTjNTb2pEzHo+BaQOQ3HQpiDZeD1
lof32bK7YiCpLG8WAl4r4flcth9nHqVRQTt+iZh/dUIT4WaeyS2ylkgdaWAhFdM6
0/VESBIYtD9iZhxVoYn6PSl851Rt0I+sJ6HFBj0JUEZ2WQ/mRiUFmaHD0urfZx1B
3LnRrAQORa2+oyFovtXnZwZC4hdxZVUo0XnQIpIzQff+zPu+PZCTY3aZHz+JpQ5x
zPMKx8n1D9fAYmm04EMVfBlPtjrgJ4Dfi2RuJ/ehHwQhFR1P0Sn3fSnOl57R9MJf
sA7jD68R16SqCNYKZJW4mX9z7WT9ZrQsk3qlgzAjLNCUZ7fSdYwb/Q37dfJRuPgD
nE7UE3MBABcheQLqVMwKZoRda+z/YAX40bSu0OVzt4FUMqCr1gnffzsVMLvkENmK
PAZ3pNzmUEQXVGh6zfVcRnRt4OLhisMXUUv278e3FYwY+XD/o+B8xqMosboCsVi6
kdTOpuKrdJVO50TYHIt3I3XWwYPW7bxSLvjgTLRTmf5tpozKuG31fSgCiqX/GY81
wFZTw9xcp8V4/JDWiMihuXzJNFO35wX7rsY+JjHU11PibGsTEXJIr88Sv5HXDZjk
u6LfRO31jW5UiPi9+RwNHAsbaP+yzR9fcFJpaep8EpeTn5r95gXnp6kjO3Bw7zZv
FqELhkPDIr9WNp84+yLSGP7vvYzrRpP1lOCig5Yw6I5hG4b38kRCsSHixt81Tduy
fM7kNvkH69ZthEgtDh8/2RtEHq7381ZvC7iE/p8FW2hVXUgF98wvuhTYHHYmNl5j
8v8BORtXpf2/rqZf9knxt4P1dHdVWblKvYFlj+M4peh4HctbxOcBwRfAFpPSKjuO
e8FlIkMJ55V9hQEsrRXlwlJNK1CK2wFQqHXl34h9/CKyw8mQw3hdrAxHT1ugje3k
rEglAoSKA/+q64zxHjMlQunmujHCWmETPalXMSmRi+8a0caiIHqiccjDMs/i0FmM
qeW4C3IS2r9Fb2MRwvODSJyxYce5cVDJIxMG7pJOwYMLlyn/AECJMQNyY4+PKgLm
92ts3FThvkxaYOSHR3greTQj+WEO+wBakCgmZlO1ZW7XNz/QCv7aZr09pk74ADQw
N1bLVYt937ImW7Wjd3enjv7U2lwZDNaPNWX6aw+yEjwjqM1MTPpwbbjWQSiL39Rt
P2Z5DMnjKUkZFIFli1O04moV4OobkG5IBJyqKbRc3JJuVu/uf/qAtALLpEGLFCje
SD1LCCy5adifyPv9vfzii7mKJ87E3cxhG4pwC83W1ufjiFyTHV8msH9/xSbHqhnJ
J+r2aKyko/vG25XB656129gIQEiAXTWLw/+a0+8pMWMzJ5i0mqWzp3VBn5Ep4ufx
62xmtOzsiNK64Pg2ncBnmv1gNYy4+CfVPgJp74IArlE6WJrbFOypeLyLalTGubUj
T5n+/cAy9CVNBuudKM+DEK83AEapjFIeyu7HPNaaEF/rpcyGWc+SPg60uqdpLZPx
69h3Vrku58F6B/vqHUTU5ue94Bj7VJe4ez6Dt2vjxcInEHzHyQL3OspFhn4lA+zc
F/ckCa29R8+tbtbs+SAr3/xe5iai4VGTOsV9462lyzcPwauDsAALn3lg7/7Vp/HZ
ZDPna9Pqn6AEMZC4IEsiHHwRCzTXi/YdbsSjumeJHeobW6hn0yh9IHBeMXEngaSS
9P36uS1pnBe9LhMONVJXLIu0qJpIre8CsEKXT4p2bGVKuB/1FGFYzlHdoiersec2
N86CZ5k0GCy+yFl1EKgv2CWthANNPhLt1ImiT6shVYM9dtCSF/zokpnPbUCulfyW
tT2cdAp1QdaX22Y/d090KBwFvHCwIMpRrxcKYBh9QkyDYtWubDGyhk4XqdlwG/gH
Wdk5d7aXCQrEn1QaMeh6vVCnA772OLQzbZEWjZzFiNYf/PyXhS7C/Aa9SLU1EqLB
wegwXc+1BDaKuZqDoBz0OpyRbTpTpb6jkUMDUzbo7e7bT+c2XwAlOCiqGM5OTCUg
ZSuqlPvxshi5C+QMsWmFEih5bxuE45gidLAQ0DgktuIVgt22oK6iCXa2dwk5se3k
ZHV4gj4UYDQqgegUKjyuHxM9lc2MrRsOGd1yjh2k7B4W07T1b1UZgL/2AMuQVou0
4UnzCtMspIAUDTSlQwzsPvug7btLpp/g3f43PVdWIHrMPE5XBnmXCoCqH3JpyVZ2
3wa18wz1tW/a/lJyyAXKjJGaqIEzeQobJa5uk8WerIXTTUyodVmKacRw6toT1uE+
VrbvtaZ+P87eDRhQLdgf9jI/ndw2m3DKzE8zyBxEHjYc53H/aKGCDBmcCuDlZMCQ
HAWZkpaMxPTvYBiFQuIPbV8T+38pZznPx3Ttc2eo+liPYSxl8AMu4Yl9v0Off/rs
YyszVoYuEudSqxY4jyyUc79rey0FwSBpBrZv9j/nWXPsQ5DypakXHCItPAcnxHcL
Aow3KT+txTnkIfBKeEMtM1jOgWkoUu7v303tUtSFqYGvsRKecfkzojwAcY6SAge9
nBNZRbDn9pIyst4OiocyCSL2br5Ee+muy6nVhPK5CVvJp8D+V6vfZnMsxQtsC/xd
tpyJCkH7evp4c+V41fjqy2RhVY18Tn3S2RdOEr4tvojIFXY5UD4F300mqUawRytC
jpa6h3UTw+xfG301ICePQNspeRgy7YqqAUn+LXOAA/PyOEPWI7hG6e2q+fPXjJxl
m8JmF7V809fp2Q4SM+WAwy0l1pK2esmEjuzbFysGk+zUBzLWOY67VbsY0ATXy+J5
zLymNfL4MAGhGHAl2vuWOHBrL9il3heLABAS98kEycauKNzrPN/4nbVR2exJtQRT
KZN94bUM3uq5gF7NLH+ytfqCmGEgh6l+jzj97+DqzeUb1xGIQxpqkJ3Tc2s169WE
+n1eZUyKtOJYfGH8Ikg9yypeUJZt2Bp4gtNKnejX0eweEgbnjLPIbxD2d82lNXGy
lgy0b0rlQfamj8r3FbaNEUaukKBsy8Fd/EBRoIHLa1qxlQG8mxgPZYbB/aD7ccVl
MEAIfnXhXU0iNP0VI6KsKT6PnVwIC369QHZNENO7dGTGQu0U/AwLBPFMCbCQk7Hf
s9plYvuUWyvm+ZJ1kKPkoAF3rDl+s/tkyMfuywZnA4q/grHFtSKJpufu5sJxHfM9
LpW9R2hw+iAOg8nljsNRI1/mYjts5bUPVw2spPDcyO/5Z23mTb7FQrrnDDQZIkBo
fY/Msi9UOCR2iYGXLMb8wTfDfQbb1n3MgWfBQfABsYHjXp589EQ2yZ72yq4XPHJZ
3tquVu8fCH0egXJ8htv0qCK64r00xW1fNIQAPS37/nbD00/XIYaSu/ssuu/Gv+Vw
ZvFVsjX+RhqsRQaoPPcYiYOEF7px0tiZ6EFZwjFDUoG7WfZuMxxlTOxKDa7gQrUL
nM49N0bQqFkSyLwOH/kYcznC+RkWRxpy5XqkbBva/Oka8ihzaUOOz5hD54HfenaR
IhLZlLXf2lbOMMPIjrv2wj5mC6HK09vLOTzlyBUTQY4PgmTtAjzujpQLsmTMjCKK
vzONYw850AS/aBPv74fxbw/6tWx1dkena7Nc10D/i5RoZOcDdyfiFDmDiRx377yt
hDeMN9nAe0lUNXRpVG0Gu4n2g/KWZ5BD/rfJDt4d+LM5prLFflS5rculjJmFIpVm
uLvRlQK3nBMzN7YM9k5A5wllPhA2NiwRFSQhRYGRlmY+xlbPiQ3C7nZZ3DNh9fQe
16XifRh95XCj5wcdG0yfynr7heg5aRRtlTDn3wmMsaIfIJoSDePC2+5BHUtllwbI
NPPrdNRhJmgcCQju770aTsDxss63wsszhmSxmDz8jiQIdOfqHnySZgESE7RrEZG2
1s2UqczrvClVOBsbU4wXXeDLFD7JTjo3ytAJTXzzRGK23+RzQvB9ClCUoQGG+MwI
dcIzpN3IghEvAiK9WbGCL+HOfi6tjosfXlSL3H+qrMjlFOreGr7wQrhjn+sJ++bk
AsefclWa3ZhVsJit6glS653N/vqAMteugoGFPvbKHHnYzYAOgDVbZsUmi18LrO9c
cpYJV8b9u6tufwqh9stQhGWuHmXkNBCsU0u3iMBUhzHTg/J3w2rf91XNRCw458WH
NsVEUOqoYqWenj6+g5u+ntYM8o8MraR8a1+L1Y+Xhv3LiDXXBropX8XAfxgaO3yO
L60FPz57DqlHFMMaBx0mS8DQM/5wtfAr85oZqOv5G1sU6AXZIQ7gNTcph9hO1sAM
3WnEqbRDsAnmJiodewydHYL2TOwS7IBclffGWy6nq55EwdSKl9UZiH0JIhtOSNxp
eUP6fPz3AaieIh6V6ZBA5Z2hBP4aDIfw44bd6YxGSU6jW7YIerxx8tHMBB+5gzZg
qxHiSoNb032IVd1dwQaHNdE3GhdGU+ED/yw9YOkjJQw9otoK3uqJ4xrKlsCnvZNz
D5CFcFYotuQwF6W5JECKy5ghkjh0BOYqlagEU3vnF7QYLgXy5QFdB/fyc3hFjPCe
5GfzCJLqdZDA5/p+zchGOdjhzEjMz5Oc2mTe5cKA6MWMN3+LQIfbDsSUuVAG/LyO
XHhy8EoDThZg7mlNfk9/rMQrh9rRWhcnh5RzfiDk1BHF8vGQQkTd5tTgd1YdwJoB
CZEod/q9+IHwhTKXmp1IPRD7PbAFpo0mwIPbfwQXmeLEXfD4/YrTdxrki0wefzpc
9ezU9XoPKbv7yUodr/T1rMlH0YixYwZ/e5OilOADKwEfJT3wgduis5Va2TPItutb
g7DfI8HqKiKTftRhiwSM2uLNFNdzkgjMVaePLUQyGV4oQnG27moiHPEO/c65lG5D
y2vRZ7ZJUTsWL1lICznRWoCaLnNKBUHhZ1aljTB4nUNBSr6C6o/8dcLDY+d3oJx1
i0Lz9cgTLzA9ni6OIcWYL4A7/KJ5LE8NC1mZTeadhTJrnHiur4J/ev7pzMCqweCq
2Zy1hOLpONBd/0FRYLlyJldYqEaBFevqRwMdO5ThL7LnMdsEopJ7uc16lPtCsk4Z
ESeYdwfRCWtZdkHW30/iRLO4EJpSujUh3RkURPOR3f5RbLwrknAEJhi1ajCxS2bj
g5sIBSaxcbKAKn4uDoKAYCRCWriMHt3GjbT5VNNYSYaxGDHKgL5j0nhMkCkfjHs9
MsV6gotcCOQKR3qcnQi7sUt5V71bP3/klF6TkaNMre1dGahZWVz3ynzwXsAowFXb
oRHsbsm+d6tTvHRFHjniQmsNRZKV9ilGGibqdJXdVf79GYY1rOFJHyxcOgiFflVx
e2Cgb5RQRwOAhsAE2ssNHLSL668lRCABFUF6U9STk1ykTL59rHVTUyPLQqb2/pKl
Ckcc4NTuZOkAISW8A7SN1aXC4fRtOCyZwiJ/31HPW6lj1tw7lAzLpCvs940WCjw1
AmuwxURr6AVCCivhl77NuwdrAa54KPTcMUMzkgPQBPhOqjYEBa1AJgT8PErwdLME
NN0Y0J0RXD8H2qjEu3hwAInVouKrNX/X8LnR4kdVn0GXpkCvJOOYgapRREV5xLeF
L3VPpEmFYO1m5tHtFnVrx3YNghaQBAV1hb2oYqj4Pu30rtpAkFb/I+0KMsLVhLJf
mzp9+xPCcD9L+LSSUJXgcdk2LcK25lu2GanESFIdzFUFdSnpTY4RqvD0YWOqFngk
0i4TsZ1HLzb+O+kD4lGl5y2h09/wCSxYU9qVUvLvxB7kZU37fqd7OpcW0R8c8RgO
fngQXsjf4dAdKq59Hmx/2viQjq/5egI03Rx0EPVqOA9lhvRhzoNOB8hR/EmpsWfq
YhzMNf/0CT7e7Bgqb7SJvJzbcy8FO04ARbOhVI8Ca5AY6prtCpHdUvycJkVw3E/N
LJr7G/D2JvRWcowhYUMVymC5oi+SpM5Bpnl0G1qv651O/9o81WM66HO/Q/UGE05w
mA+GGhIYPThGaUQGczu4XiaPHWJDrr5werBH14ysb3NAKlS+Ii20CaoaWY4qN1VH
RnsKqs2WmhMBDX6tilIXSYuoEm5mp78TszvUnBEYC/T1SkS+h0u7YL9sgmry4ZZJ
y1k0Xye3IkfbI+33OrFk8uwVOEasVn6TzZ+qh+gNpXPLWSbuBel53xTnVnH93sWg
8ARS048+W+GEpH5r03yILej59uEXFmtu6nohtuZu54Z+4Kv3L1CsIGGQOkfCeNSx
UYiWFbbl/8Dtef2rxToca7BuWU9qJo6n3DNjRa776y862XoqjXfS/9rWq8b4TcE+
W4nYyUOKn4ZJX4Tf176BVnlsGiMoqkQbosuGcCkc+4mDgSODTBySEvpQiue4hDuD
8UWa/bFXNQEu0t4q/tkzbn56S/3V9WTFCcysFPcCizWul+rkLiAFOJHg89/D9hgq
jJntAaL873+YndWKIdq6jbN0f2KJlo9omAdjtMMOm5azgzj+NnMyWjaR63mwO/4R
yW2dzM9OSIEcnSXM28Jbnfksdb/L0bar+E22qCMzoACrno/tj4Vg6HzRmBFup6xV
H9ygFmw9r9L57nlX6CA/zehU6Wt/77MNZwDCljWbSE/SQCwDtPwSG+aztrUNaIfj
ZLduaoQ/vch+kIm/KphjXo4iGlhygYVIH31XSJ1jNaKBvwXr/p5TuYV6T0clzDie
3i2mpSXj/av4HaVMoZequPT89XLcWsAzPR3PHUlrjOpu+ttb2pFDrVWJmXoS7yb4
4M7gw6j4bi4bntyO71KX58pc7ztJoOlcM13C/5oAJPhv+Imo1taROY2VP9e/iAlW
ftfhUeePe7C+MJGjSNid4lAsnHo/qc0SRUVNsXwDzvJBOeDmYG2ehPcxPEQdPMhd
QfTbjzziFw/awzoSusbgFu39zAyjD0rPS1wN/NE+pFa5RU7Waeg4iq0KUKx3VZUd
j4FvgLiYNrQBEm0sGIGo9F8B+x2iIue9tBnEwpkOkQzZmUGyzohzGPtBtWDeerLg
r5bQ003oal05kNIq8mvi6mapUWFzoM+dbXMXBiYZSyyKm2aiJGE5DlWV9R4NZvuv
lLjTiEaNXOOvS4XR8n48lvM9paXMkvqt+VwgUG8g0I+0R2VkMzkzuGxl66IL6t5g
mAVpR03sHxPhvt8ZG/n1ksONKvgN26zomvJ4zpSXIADytbLrWi0Q5ivcMX5urgP+
x2OsgLonuvLEMPvkvmYmX8vJXsTleMYt3HZo5q8J9/IsTxvgwcO5kXNOHRyg5MpF
kUZDip2Ex7afxnRH69NwEaxo1QBu9WKWYquiPVMSGDObXaPZN6ivwQtts02Kdvlw
3xjQMlRYFqus2532/gXfxarAL6vi+HRhGeNgHmq56GNjzTL2CHz1pD8jPItlxU9K
TP/rEHToa74leagMhF55/NTK4e5oe+3yUv8sJR84RH8v7LXGuCQzDel2/YIUluov
eM0iTHf4NVTqcgfpUYDJkXPt4C5zrsyml0ig89tDXedPKJa4zNE/6pVytuFoFVHk
LLfKAsz4SevMCcR7mJmCs4+GbKvnA3SDrL0PxGrJtjANZKxwcayiqM1kQE8QqIB0
E57XqaSpjA+WRqMCICsnd7ofoUWzvSz+RbTN5RJtiJNX3YxDat7UVRXDywXwqNFj
xWdVsDsUYxsvJXFrhb080el4ptFIpJDL8+uKuaUOcYx+itOplX3t83yPHs91FFoL
mn6xrSTTMEuLk43uGVVrQ6DXxXWRR2w6u3+OEjBFsoD88JRWyLkIpf3CCHiAAWtW
deL+CLJPqKzm+XkIYRypChBVCzNAHsd4uQyjaqqrHBwr9u4q/KzNie89/wSlW6QK
3g85s+GM08XDTGU2v/vKLKw6e1cW+2bLq2bxFXJ4TVf8HwdtkEFHXMEr2Os4IPIQ
WNlMrt7qn2MH/D8Lg22R7zC6DolBmCygPA0qzO3d5i5o8dkALe9b9qevSyYeuAuN
FpvV9xBsrovZxUyRTx/WRloA6LNp7hE2XXQ5GO5gvWOP4SmH6IPWXXU8ZnS6svAd
WwpRVLQhbj+RGcxkWWyiKqJzjkH2qe1lOtCh3q8OIy8NbeZDz2MNiqgEQWl98YRO
xoOV0UV6JMokL37wP+GHlaeoarM0/jhUcXoZAuhbuCnICrUGKTwm8MkEpA78PPMw
C+bFf1nEnPCb9JpzXV12fwJ/s/QzhiKK3ObxXv8mb1c2LGaoFQzEDA6Vi1WqVPWB
u/iADMO0lGmYlwJjkmhHM03JhgGYZ+CozRdeQCWhkEXs6HstIpkjT9PiXAGCN5mh
/o1awq6TIp26k3yl/feateKkuffY49ChvtK5Qvo3zlrPr80mdXZ4gDBmnHdnig/q
fuDnUuvAbrGgTQLIPGvMRUAgwADnnw2s8lAC0BF31MUtk9dYyzI/rQuZYZHSGWOj
YYkJxR/56z83r6S8AsEHkdc3gqnWB4FmKC00ahIaJSJ6h6aDdbKQG8k0AKutiV7L
lpiz8y00G/fjqb4wXYfoR3HHoArxDSRdoQI2Qwtpkl0/LazG7z/tJ86euzvuQJ/k
+1EAZXfE3qQZgptYKjGVJCBFbcMApNk3FKBVxndB0uqEoW7BzHSXESeq43A07VSH
RYt+1ilgWUCAorzUv19lgRHI0kQLSmJOVFKPDDvzgiiqd8GC6DS0TAGO/5PrBYt9
Dr4sn6xB8CHC9PB8nTQ9JR2MWE04rMoYUMvtqesMZJ3PcvZygNDZPhH2UzesNnrI
TqJO8Vq5OKDqS7hecN8LVZs34+0nCVcnRIJBLmQ9+72IE8Qt/vaCnz89FmQS7eQE
wDE3N7mImBZEapzzg4Fbfj16WZT96D4g2yT4ojAzRRi7u2Gnr6AYZkJEKUs0jzCV
jqtdAOwew8nZDP+TkjYTllk+oHGPprD5xmCujK4JbFbiSkfcjYwY1+KuGo0GkqGy
/5No6eItCOF9c/DrHy5Ma7pWcTGANU4zphwOJegX4lcIe7QOrDKXEaPS0QE+QInY
59hM3Bk45lvTDs8WF3v9/8VmBNEciEN0QsENa47zzeB8Tn1RWA9oVnP7PqUjJela
J6bz2KbGcQzHlBaPu+Nv7x9u7nxJsxJIge+tjPJmvIdkFlJowJAIQRizkJfx+nja
51lSzbWaIkmKWPIyTuejD1miCi+aYDTB+R5ZIxNyXsFJES96qrwVvPBfeyfTNzxo
PP4WDWfkdjUcmg2YQtqKX6MtG59CbHRLwlLhS8UVBh/Ey5ZdIcn7Ik+AZixI5dNP
iusvwgP2vU+Tzoo+q8tTuilOc7b9pZq6KAJedDvXL7Pw15Lpq+4btqdslqrvK5xm
leiaeBV304I6qLzBs9FjM7DveOacqg0F5+HrMBorNZc/g/88urGvyyUZT0gYAkz/
tCUBKuRPGcMar2HiXr6T8dsPK7GQfW3TmmtrPLpTCbKwlnWP9SKAhFP80PYg/2IL
BEVfgz0XSXDKsoLGME9HvKIzyiAe3L3bAZASjKFbB6p86fuy7LNbK/dpPfJ7VxJv
XGjeOQdnAhfjoo4+oYKGfBGsYvQg8VlUXzwKxRAuLLQVs/mqXlxknlAi1d5ps+q4
Q1Ffv6L3Y5FAOa9cv9bkQh4s8txJlkvQ4DVfBP5aW3mDYjx1BaaGJ58iYtDLk4No
YaNvx33X6pC2h5EOJbJ7hl5xWMXmOu0C+gpsimIAz9/jsaVL+YYNzPW8qD4JNpDT
aAT5xjAWofHwDQ6ukD9e6tiF/cNcJZKy0at0hGt0ubWOParG15n/TTY52I+2kcsx
OZEKMi+LSie8QXKD/9X6Blmh7IhnBSfpqIQNV6m6cJgQjaLBOzJ9NzxSX1iBwvEg
hm1m+ojjuyHdqJfUXvO7UXZGQVzGGQ63mtYUDL/DbBruTT7IlGquKyPy7CyZhQh0
qbyT2o6EZcuKZhefHjerrJrK4Xbt4RqIk+JoOs1UPPXJc/DiVYyjSia+iM+qCYKj
OLBIdEs5f4sJVzQkuxeZ997fMzNIpEec/VAmqQl908VFP1CKLcfB+uUgpwU/j01U
1H2VIIGrhLU6pGLMKkm0nVcemPQe/k456KDkjqnaB/+jS+aKBuaK5F3TDsP9kV2J
ltC8bDa8Bejqkr0M4n08FZMvLQsS3OOBfMIbPdskXcRCYIwGRObvOxG8FAalKNJ/
NzfbQcF9Nby/QwBaWUe7qvPG2d2QZ30ltMHobRqn4n/ZLCN1W2IXKarsGtP05nT/
ceTpxQk3CRuwhbhdiCA1qq4W2wHPgrauHs/aSJ3H03eslN6arDFzv45/VuD/mPcm
vVskr5rblhgjYuMdlsc+GDVUKKN+R8opDKeXvF2FEKwP0WzbE8u1ngpmLaMU6SjS
WHBA9kgb9d6gyZ24RzQkeUM4Ij8QbqhAVQ+yGK4Lp/ZdhM9bZ3i7i0FHaQyXejGx
MVvccV9AyRYY9FCYs7Jkd5i79ggyZwyD5lwts/aNyMi/r6XsmMx4sjL1kZ5Lr9xz
LctDqQ9qILCVbMZS/uVXrlPs3itzj+GNtJxH4X1YBdih8GDB/mY/8ZS0IeK/Z5fR
cr0gDHhjunDut/ktAG2Xbw1ePTrJA0InLvejr/i7kIv0Wt+zasZhIgsVvlSpGZiM
tmb7UsOEk5qg2uhikKFenfcbKUfKCG+ORiUvia6gO9/71qqglxD6uU4B8i0VULw+
PbuFjjEaBLt5ZSSvYcfaJG9Lv20GmH6Al2xw9pfer6p+h/9tvTVxuizI94JE6k/m
YcqNQhXaBOXN+tnKYcuBnCbU38NSpUpIvjISssw4Yb8DeHXkKkyUJxZpoasbH00l
9HF1FzoAKkMptnrsdYvFluJeU+tQC8USlmJdFB+0etFNUKyXT5W0JdiAsQIwScku
dgUTpjkCh32sc4niZUKk2PZmeaphr9gzoo77fZjjRN5zf9zv41vFLP3/agkYpqVP
raU0PbDmU1HD9gBa1IhEgug24Tbo1xiljdxn2CnpbfvLvF091srDCGTLURbrdnhH
VBTT4lprIe5qHZr8ahBSSSwftLy1kdcBlnyUt/Kf+CiKgJvxtBeGteXpNacoQU1s
Wl+ckDYoI9pjkUC7hN3Fg7INWND9CBWDMj1rM5Nj6v564mnkP6Olu6/6x0ScSxqv
2XMP5uMa+imbsnPfIJiP834+ZB26ruhuiJQimwA8NBbT6t05HN0zkyoadAQBmGyI
LnONwc27F4x0AKPjmwTw52Y+BfMslfz5opwwzgrRAmY4VSsV9H8MlSu8zQSKfy4i
vH/xMC2Pgfgi98dxIxUmjskejM3AXsgz5uFj/WQelL7EX4hviCQi6BbbozWR4j+9
Xo1peyZnTdxSN2jmkW1s74TKFo9afcJbHabbturDGGz9gJoaSLpSDFWp+VGDH3yH
sdlvpD6tyNbp1ayEXO2vCoBdYG/bfCiDFLe3SAWJYIBe1ZV7X0QZsuS7Q3F8WEeU
m5wClQ7iUAj65TgbfDDELES68RF7cdZ2V6x+y7J3kNsommTVgalID4V5SU9ws/wk
Y9FBiX9k/IB303+6jLAkSJCfRqi1mVt226bsUN3OZLWJLfd60HKgMhLxfd0/waxC
dQsBWPrFlXGZUKe75e6PQ/GMfgyGsWTbYzA6VHjHoTUUM2wTUjrfkZQV3M3VaTKW
0dbC3iJJWKPzVTqt8lFABJaKBVe+BjqN4tmO/BNdPH9ZRVK11RDwPok9ZjMqXu2h
tkPexh/MumSqCf4zwpyHEK3amAln7L5jPnUWNyLS5oz+k/IXoqg5t4nilMpNm3c/
ES+h/NY74/ae6ixcN/Zh4GMoGNQeSoaDHN2LfhBkuGHHyCsZOcVQZWrCiiEg5HSv
dPj6RovBAQdTDQCZ+U6nYllrP6FbCqwzKx4wVE/gl5EYxPyJ+77iXyICdZmwGEvM
WqmWf55uMtaDm+UaHDgEeJKCalR+PHvbTSVTEKj0/tFsAig/05pR/gquGofL5wqv
fLmvPjbZD7wVBCdEv7RP16QcYyGK7rXacTZyjXETIU1kOIhPxnnk8An1adu0nitr
8uealudPtz81DRD8o8sg9R0U6O8PyXyVkHy24Aom3Txs9+F9mEk888GrASVWE8cA
chh8R8u8JCeS3T9NLojObE2zDhruOWUQ9pAWFPdczq8jtGIry36EDMtSqwiz3iLp
lSBmGynwf/Qkg5a5NdM2MW9XpYbOnqxzgPMFqVr6LrSFngZFINEGqmfSP1x3lig/
oBSdWiZZ/jYgVuUlJGNVS8yqLfcX256ndIE71f+qkUgOY2Ic6ho5pZykhMryEhan
MVMWS1RiInMF502X3ICSUFh2Hmb/d8pxor/Ued0Z9Pj2O6hwr3mFwvnexepGJfRW
tVX+AYyo4SEL1GmJ4aF5xshoKL12vliSGvRIAS1k8R9fUULMQUaqKnTysgFkgCxE
0MMWC04y8ESzvXFnz8Ubrwq+lU8KqxHdD9K+522TWeJwlSpJO+nL49rsxGA8DCuu
eIRlJ4VH8zjudXLytHkbCKA1Qu2Erkn1VEHJuEWQqDsxwglK7lFQWILFS+tatxTk
k5gEFwfi5Hif4pzB5NcU89frxppucs+oKLAjHGfzdX1O07mnmizTcVUM2G/w6Efy
gnpWTYeNnW9myKwYOep4HO6VktiubY5h6ojLvkWrIqRqZwaNPs/19PYlrz83MrgV
B5r8afFrP2Z39HSpoR71Vi1G1W7U2UlR5MARmri1DOkBIrHTtN186PQYiAd+USgj
5/N0EhBidT3j11Gg57F3VFYbO4Y22fA0Nm/Px3rs3ErR+xHZDdatX0/I3xxR0fOQ
SlWhpmcn0gquazRzANCD6Zgdnk3KULs3dIGo3He/bI+IHjHxKaLaVikX9MsPY11V
lu3zSiUBHS0BwjZlNaeUAdizyRUineghwkCikv9opM+nJCdIIOiEju1nbGsa3bc/
LN9yXVFysjqbIAeQmnAIsKNDIM9e+nk459bZxKrrAARGPZ8fEiImybMpk+JQGLSw
0YphQmtpyeeyw84+2R4e5T+CGrCXuu0VmlbYvrabmcNbsGezgUD9tKnD/qRUDBJf
NEDyQB+72GKpQLyDadC/iJr75czPhTzXk1TeWCJuKH07/0Uvot5L3YK8CcjMarGv
5kxY4JrKU/5qRX4yFBjCx3jVfbCAlevvXJwrwXRSImg95hxid4nj6BH1UZbC/L1X
psUBMkzZil/ZR/vR7BMKw23700ifexC6fhG8sQoEKkB3vD8XbW+sGOcyJBXA0+aT
hYWZfxjGOfkRyWk0guWWA+c1INw8cgjSmchHjf7TJsN8Q1dHfrGJLNbi1CmVfDgF
icRBUTBDyUo7BLApacWDGmpbbPOVxkz37RTArb4kOhmGr8XyNxmZtvD4L0esFX6M
l5Y6kz45MJBM+XIBHfZJXe5uYEhrHaWubBT1S+xT+JLXsQPqFjfcKcwAETVCfWcJ
IMP/pVRhm5Wk76KgXpzVSRqmWxGJoqBv/LVZFX+aOLQU2N+sPsR0z8Q//B+HK2/+
3pS2OagW0sC1gGRR/4/j2/Htht129fCU6Mgs/ruZUI7VZgnkqE/TerB3ttUEmlbL
8AFEmA/Jz4HT8aIpDGKlTSVG+cnctq/i9bi8/oUy855SzXxKK/aKlqaObJbQuQO6
+3AXwH+nEcT9MwNHlG4dQAj6flBWliZlHB795l/090tnnKrppPBR73SMTlP0cCIa
kUwXoFFW6ODBT+cyFcnVbXH6XDfsB/l/Kg6IFUoVclTkoBcm42oUCkGMjIaorfjf
++FW/exSplZPMRH9DyPA0EzBMDx/oPsXJis9vMf1wmynkIihw9PJDaXjBUTu4nuE
9NLMBiXTHtbjpw08Nf6xQKPQnc8UFTe6FRum036C28fUisZ3VgReCHzENDRzN2AL
yrBdoP8pS2eLSd5L3FiZaQExh7JO67ZyIeiILR73GA91SidYOsPRtM5PTtBBcETd
DXKrZtztmyeAv9WbawBlgqssDwpmv62jhI9J3e1bi8razlNZA/TkVEzndfPCUOFz
4YlRUHrXRd5flRi9rRCssMeEKPs4a92LLyULfrOO+CxXFWez3BZUuPtP57JUlUOn
4O97/Ct+LOVVm6e97Xy8Qgn2GgtB8e5l1G5ZBn/m2c1v9CwmhjZuYqDRZTL3OTlo
vi2IL/CAu8U5dVPUxYul8H99oBVWbuReaCyXLJusYvUoREuX81QmVYf/Pdj+p7zu
chIHsCmO3y4hhWe2XmOF/2IQAX3MJ5aBMNQo+vsPGmYmhBsueS4UkYw1el50I7zQ
dMLEtRUTGDq0rskHaYHygALmouL5ekh52UUXyLU5EpwOgmGc14OpMINVBKCbBYpm
ub95Uh9/xhyyZfUQV2fvzKmO7q1np3YzFht6aTwDdoZG5Dbg9oZz97dByiS08ZXj
fxdRUmWB42x9AymGMgqJxgo8YiDKIa6RVweBkQ7VjKEZHKu5glNG/jYVJoOqcfn0
RtIX9T9zZQ3+1YJahQfanEsvU7RyUQzEHTktuIEKFpoj3phZkUXDR1mXX4h+msIN
Mxj1QXSHtFyalCScUBvkR9jAjvYHAu0zpGycPXuX3ksVEZo/veVtpYxurPb3j/5M
pVHJoTT6C/u/M4nAb1cBd459+0/pUmAad68ojGjrKNTjWTBbAxm+K/bBjou9TPz3
n/8AJi1hAMaZ2JI8hpyMXTwrgrQjBzLHBs2IrCfwB5lJd2HEBPfsvuGcOih2Li/R
lC6zNp9Yc9iq++8KPU1D64SIYofsk/z1OxpPnrG7IdYc/JMRB20kTYVjANgn1dVb
ov3BxudvbkUDUMn6THsE9BsfuuCmQFGtVrIZwnfI+B8k/i2wfSZ8Yq09wudhH+vt
/gCiQQrCcLKyrh8MDTAdfe9R9vP9yKrvN3wiEOeCEBsGM/WHrkUJKMw/NYNKmR4g
1X/mWWjnxPmCEij0McTMeWGdpI8xbQppWM3F4IsJ61ABBZXJmS2Y8QbBQZ5PUn/4
djZLZ58ECACfZ4KC8ZJsBKjahM7fBmJFAEl7rDE8xTsoLcyER7OoIhpN9CoAKQuO
DLid7FWKDbRnKBJEgfxXtXqtt06uFoM+SdCi5gqiOWGuhBVoE68bKUVNvxOIelWB
ybDmpqQHf3S17Ng+pl+Wtk4zRj4yZVH2m0EhVpgHqfBMTRto5p6+8jQwS+xgs9aA
3A/HpY3PE/9oVKfSewtBhSCmjhkAH9kCGhNexGE8RocdAi6RdPghdxoepqbTkvtj
gGBNHQb1oisTS9KetD+qWBXO9W/cYBHNluANKg3+tpSQDwvMh8NeSfrez/MeeE1m
UW8fcS9nUCpV1pG0obzI5GHM/hGynPV/JdeAwrkr2iiAaUx9supehDYEUY+BY6/A
PFpoqXTqljnDvlKrh8b5nr7AHzHKSstjTSK80LjGKgsnCrgtVpKqXksC0k5lMwwh
tn0BvLFGy3ccRCBgIOP8pjTFsQPI2jlVvcqA6wCrmtOzXcZMfJO3nKDqOSqgK5dW
jTS+XgF1HWJILrV0xjW/q2EoXIGgzG8TJuHlpBWlIFxRx+dKU4QG1EqbJx5XsRPo
w9Q42ImnIHT8WIImVHdDWcW43nDR+MiOrCMd+c+zphPb5Z1Vck+ZqSfkWHhMui5T
MAq8Q5eB9I6svOX64AdyuuFkQDHlei8k7ZP22KNmrKwnt6dDKi+OeNN2xubM7JYH
GLrqPAcfSmtMV396t6lT7ijWzGl/cKxLbBysNBzZ4Do3SxCsILArgDeBFFot5aEY
RninAmzGBgnMR6wp6JFcPv/54oVbqdXCXUXYWMKHfrY63tow4uebfLD9hQVNZ+8b
wiAK3/+tHaMAMXJpH/uIMzH+KPL70Dem+pj+TY7HoW8XhZwI8zHHt7zgpF29k2Xe
J2WjO3mPEY8wxa/AdMT4XMvstr3MZR406NGuL0TmTxl1mwtNn12mPpe9GzFG/yms
uPpcreeZMyWHjI6z7JU3BvNuq7t2BX1nAq6pGRd/LpXaVB+ktikF8QgMGmXwui3W
E7HhkpbyaEg1FoX6TVGQLS50yc+z3x9fnnauSXeVMf3x1a5BzzEWv1phs28HB9Fq
963BNdvU1qz5fZJzVz5YwI/BQqnnWiehA/KBha4uak4AFeDu7ojz4LZUsg8vaG2q
Yn69BG7LiyEooNzXFLenhUeG9IHatkMFIcJKbyY0C24Mi2fF+naPG7kt1tzkBRp8
GhmsWP97sMsrbuoDhrvlz+0Ak2hNUTTgiBhXAvegEjvNTm7iGVqY8f0ay7D/kTMY
gkFmviqC/JOb3PQ07jgXzt7ezPX6LhDbSL6tdv36J9SoqgtWYsjB7koKF3bjPW6K
ZaDHuO4T1lyru33D0MOX4SkzvANxhMswvzzTlk3RetOKTZHaLUWzE2R7moAicXyk
7pLlTjiPDnCoJ3uidq0/pSB8YYxmCGeh1dySemB1maZfXCV7EfHvSoFzZqorDRF9
5KLfZEDdZpYcgNI4fdc79a8059Axxr/7Vh0tE5HTNe7cHyMpQkRfdA8QTrhNx2/F
GC/WEPTg7EzI4BUL2HwovzXbGjDykkObqs7junwo1YAiAIednkm3QveH6vqrgKId
iJFBA7LUQ6L0Kg9AfXJaYuiP19lxcRuq9ptXanG5E1eAsxWPBOvgKNTNBde9RmGo
83JeOcBQjx18UC4m6nRx7Rb/grXghx2B5SqA+eHMq2L5KWrymHST1Q9aQkalL1ek
EXkksGW5kL5DqHdQbhX6OWRHu8/znOknJBNQPbmUgSsJVDZxGDlQBRepOxfzIOME
jYQz9f+bO2SzkzplYuqgdUqiIBpeJ5UQnkDHS2Q+YLSbUSLIJkFqTYSwRndSerlT
noD++phQnxUpcnWULeru8uldQpofGgemOvcODbOa7tvuvWoHGBQoQRTATx/nNtcY
GxpGG7tXfHTkkp9XSmYc+fwo9nXdMIXzQlYUm9sT1MoK+wxLkXjP0zyib9O7kFW3
YffoqqnDfrzH7uaFOBdg9su3N7G0uLr0u+l9Be+ObBwQjITXn7bN5MIsLuYPZ8xU
pEN82JJUWyUnLdCwK2PWQxIefJK56zUFFNr0c7oRl04leUhahLIcbnyZPxDNP7oj
oPxZObzPi4UmWuHCNQa94HZOpSDKB9qGwSzKz5wWq+NJBPD6v398/Ep72xRmV+0/
BndIeWwaMSGn5IMV0RIxu0WvKASvk2FWzsFhO3w2RSIxpEviKaJuz+Ma0JAIfQfK
mEX2tiWBksSWrgPD698i1vnslwKsGS5m0nBbVlEHTxfj/SgHctIpmZAyQWttFJt5
1gfpdr4xBIm38Df4TK4bo0hyWRj5zxA1gIvl5QHyx7mOYTGI+Ev8F9SticyJBToz
oVYN9YOp3ahs4rZcJNgHAqR24agx6lzGaHwBrnRR8qCwJLll3C/cjU3Ozr2wv27z
zvfxNvBL55Pfcg3xRBO2c7DY0gkCdDSNOjfORRhkdB9yUOZqpuoY+hlvz8VSmpxe
kEkIBk4C+tMf8msZ5WX6Mu21ZskCGxzx5Q8mB+4SSmDLYlC+OmR52K3dpj4n0Hj3
rUISY3v0GWtTloeEvIv4STIiC0L946SrTOGwfxMV5gI1JEuNn3iBvo9U3SXgigkF
NO+lub1Yh8plmiooYNU+z3msHhDm0PB2tMWW3qzX8Km4J9eC8W4Pid1wll/w/cOy
8SPzBM5lvplrWH4HVkMp97aOPE4ZcZ4B3SXxyMD9R+qAbXR3tpeMwoKrxoExwMgg
P3TjmnXOWhu3V041OH5FUCLMvVb0ZYSCVgb9aDkwT+FGhs8bPnKnrhD9DSiZ8ZIH
iCGI2/G8u/DW++H2PWDgrjvTv5KY/HPwDvwgxSUz+I4o9YXeq5c2EGX2vFXpfiST
iJqSUDShA1x3IJFD9+HoqyepF5SQwMcMtjGyOnaBP3Ezt7M9yFB74Eq56h50SsSm
ZtxX/j3OUiQCDBvTawCuGI0/1jx1a9rCclus2Kgit7s3qjZCqjrNUiFrcnHRxeM2
/+fKlGwb1X5oBFyJCEDsRFeyIJj0YSC5OYcgxzoZbxUE/7bs2YAtTLJBD0TByYUt
P4NmHpjXioj/6teqS8So0PPZWq6A6YWDFBx6xXMX29OypH/2n7afRoR86dV27MCc
cXVirRO7Pjfb37ZIAMnqNgd6zfq1OHCHtSZ0YKPU0wmqLBn1jqE4AQdIXuoBF1wK
4XrZUSSD17CoIHuB99GD7sHdhOEJGO2jmWTy1DdaennVi10iz8bpnk9N+/gX1xaL
Bvk4RXRawTrLBdO1aMPCemgPNY6Y51TbHzOdUmx+DvRCaxiN2OfqaSNACFS9J39E
jkOWO4f61eLHPr4dRwScjImg5AXSIfFB5fOTiIbAEMfPhPY834/5lMmM0klONWDU
Uv58Kxnpi8BdPozfZBptMovmX57LQL9/81xKSvdrhHuGPcXytOYlFZ7UbnxDoTAl
ExePPRCBQUb9Y4BVgNJmpXFCbNvVYUMh8Mea4BIkQcr16iVWbBZ4zERfvFIqYLjw
dbX0kVktryxSXazohHziFtgdj8ey0Rg67zowTURp7Zp/eolki7tcmeVyETKndBwH
hcsJP85/3/vaFLwK7JTF8Fn4v8wSfQrnHvN/6iRw0GIquj0+h1nHm9NpL2zeVyYq
YOIyaenthcxCuz8qDoh1NiFIsV2mWlbKqgZXmsIIbQWDqBL4+eVxToqLJ5ndI6BS
+5clScmCwE1gzwu3PNn+sGZhNAmFmmZo1szjolRiF277NS9rDaAtekE/B8bgTmvj
NMiL6P85QAMldMeZSRIzU+p1Q/DDQBORmN+Scc5POlMAmcRX8u3QiT/ofU082SF7
8TqwSyIwigGYHsdhGlCw2MwPkQo7z8lbqefin5JDofR0W3hz6gmaknqkxNV/q8G4
QIsDW5DFR+Ua/nt/glJUPiFB27nJURpQZoCavdLgHdN3cl376kD6V6q0yBUENojr
EZgUnQOAe6yBW+Ckkx3HhZ3PZT2aVQOljbtQZMHZ8YMfMiQhrEz7ZsN75w7hvXGG
YF3VjCb0lFUJMZCHExzU2TnCCcTpQryr2jvLO4JPTdnffbJyMB0H1lculkYfUgw2
Ar3yf2ZIppqjcc4q4zmoScqUwwaUmU/BP6NKiTxR07S10U3Tm9jLbz76LU2hCAop
i8uaLilf/FpIYffu1lcJl/xVzE5sFGq2VVKHtKrBiARIqYNiAcmWb0+8tnasVKi3
shlYFG4vtC8zBAZ6AxVgwrsJ51ge5MpxkA8MxEozoU83sapS6hHjeUg9Lxe218Bb
evnHsDywxyPbTVCYm6jCQl3rZKVsDIAormQJa7zZey5KvksixCx9DhgMch92wYUP
1VOePq24NTkpFJqTgE1zSwF5wJdwWgNW6EV0VxQjLV6TCheOpAZ7BNll4tTPPliK
vvDxaopq4RmmQykmyXBzpUpbnwyeFZLHzHC43RD4B/Vft21S9ya46Kk24wdEF7TX
q39mDQNVuj8aVajNxVsfHsKXgsL1uwnCpAYy6VgAmnfqZO50Akuq3P9RAB5eLmNQ
TIYxucwFehXfZBIiltpWhvY/GHpmsYruKfbAR1+5i0ioHS3d+eFZx4+D9bAnQc7g
5bv3VQXH8FxacZVpGsL+bnfA8LXc8i7wvKcBFp0iIQGT8z7KBbNl8d/jaseI8h8D
gLnVq83NZD66dkfLEsD9s9W66dbUD7SHSGYmgaykuJ6/mdVg7sPxYG/vyiD2KRRg
3ddIJ20fsJ+alijpNlaXwXG8ztUyUNUl3Ym07EL3epgznF34x44EdOdurTxu3r+4
QtnRKOWZGDZhVbNH4khzvcWKLvg0EQlQF+rzwZULAyFL3e5CeljGw7fe7UxqRDsf
4TjWJ9bBpooE7fvazDFatLFe/D6C3iBrI00nzNPwxj5iJ9f06uKOX7IcUMHjUrwO
Fzele7K6j/nmbZWZlHh9C9z0jEDPCSUmDWw1kT+6pWnxNw9pIb2YjMC5Gwu6VTNl
k9bubjvYO54rVhGt9JWRTppiIRxABITNw3M7lch+W8B6kefmcmQCVKy+dJ7y8L/y
qvPfiI/Nw1Mfr/K3WEY4wOHht8HBgkC1X/0R2/Qvi9jQBKTH9srRBkkbd/QZlK6s
c+ze622NQo3fqnbGyWtaRSbG45MbLYWFC/hGuZNRlukB4cEdIuaKQFLnU9fydBcL
Dz/7cF9RC9jhm7YtfR1TyQUbdtTYF2uKATfoYN+q4jQdq5uCwfmyVXbUkGzQBWr+
545gd5qVnPpXyTXdtMikyX3xaHyh9howpsMFbJtq7l3C2Zq1xtotx/EwU4z+mu2F
4SmN6Zld0KZxStWGld7RP4/NdiZhWlnJDI1k1r0hVnBKZ468+POxGJ22c+6nihTk
8h8jTSbqyYPRYWgZIQCUz8RTY2hJD9OQTvp4FCydBWDVu9H33mvh//nO3fZd+MFa
MN+3F8L45Xw/icPhjU8yMDaJCnV3CnSBKDOBYUToZFSKfe5RbstLZsYBXDE30sko
0sbarVvl8HvH/ZFKtI3yNKeZNTAEJKhFLi2ZkQ6igA+BiDE6IYVMOSB9UbK70giE
Jkx9INqOXtCTh+2yeqrFqdiin6NdAoea/1hkdgcsZEYN4WyRke0To2Yz+JoItIE/
YHCa7sSZZdDImozW/5CtkHLuEBlL61A0AlApu5JYgms/0qYhwvb2h35yVquPE1RD
AesHs1DpKzWWCDwpI9azIuqW6KFdyiqdYAcK/pzCfat8v7XlhVv03hFTmnBKSyjR
dVZQTzP+kyXmXCY82zGsOX/57rXaqvT7uT73VCDUCIBt4lbeEZCHO0vUWJePGn2O
1pGZ3V4ThEGGZE17IsP1ORiUMyVJtQPEhAOCJDSWMQe/CUTYm1kRDIpdBaYBaaO1
vxvawTG10tun4wCPYLLad34+1uSy9Og8vFp5GOGL3KN0vsxNtGtWOux+O8A4ywy1
YSiielIvzs0WCom+njgw3yLP1CVyGECynaGy4tfpd+9s+/F2ls+Rf5Jlb1yTywzj
ZzWN+Ocz3gou0f5bvdf4cJ7Kct1KXIfIyg5LXX0ptxRc7k2ZveUYtb77aLJusTEx
MaOYv8l4V0YBWmWs6KUWLVbFOslJHZWUCYd00oq0HqKoHofZvDDsvKgX44QmDRRl
wm80I4g668GJxfPkzTcCXemi0mZKU2UTYo+7rhyItUTiLRZnBo1eiSmLjbMW1LBy
hvD3gah5beQwMTp4/GqgvQApEFdwg3CHpdy4Rr+hu7/xX4zbHOsCv1VKwvGFUj5z
QIEi0P5N7QAe60eilGK7tGHbBG23gS5bOd01XXyiOfqjcnTgPn7aDE+GealMm8CJ
xSnEv2d4TvOU9BHHmoM8jKpcs0YJdAFF5UHd226q2Bi0Jb+Zzu/HnU+N8nyehA5r
+NxqWk+HweX6s9S0wqkl6rYs6EgWT/DC1pELgw9WHBGeZE86ApgtLyevU0C/8JI+
FGyUb5v+RCI1lNWg+7p6x/eRdqEoxCnZ2dc7L1XitJmu/E8wmUfM2B87XKybAkPw
MY0vJeKpCJrtdbqGaej0+ME4gwO9ZIDp1TonnlyUY9POjOFHS637EXXqp12K4gp3
O3IXPuApPL0VqHZfxxTPhWGK57qOPWiEKhoIZY196d4WpOe+lbX4juYRrBltO9Ei
y7kpPqOj8XHvMaCjLV9FD2tWCJuP4rmGIV/+w4ZLrc+S11vViVGJCFEJ01cGRvoQ
7MHx1kxtMUrl2ER0xwZfhudOnceho2mT9qIKXkPNHp8M6BoQBamfRaImVYePQ/h2
qwvSrhL1DCun6RJk46vgTbOLxE7KNaZ4dnnUxlE0eImd9vFPw5NafUDIoOvikXqQ
NcdA4HvfbIGcNj3LRowrl/MwYAly97Bjyg6FVnhIPiEw1hiDy+7kPj8H2Ekhqg8v
SvQ5Lshv7dP3xEVqrME/Y72ztiERBkIZwuezvfaKZCtN+mX4QIQ9O+DbCmXwr1Zz
qGmzqXcX9teMTMflFPSuzVzVkCgJcvECKumfusdmccSsLdEm/U7U6FNFxVfye5al
wNLoFHX1bNJj+J0tYRg25sYgzmy/ySezGb4GfMAKMRT6RUNXiXgObTVftd1nNAed
iETA0c/DOzBpu6AZY2M0IPhLx/AAuZtS0dR2YsaC+GlcWwGpXT25GlhsiT3jiImo
QoJ+cTV5UXH7FSQcIr3ndIcfIUd5vb/JzSu0FkQhkCOUqrY5Yuw+iiSKMFQ+R4L5
po0CvAVomoaXK/pyKMcHUfjqvxUlaRvjg5eeWUGpNwo0ho68i4cPVX0ConjPnMsk
qv5odK05yAQwZBEQFv7TIy3d/Qd6nEOZO6NkNVo3Q/f1TTD0e2SeGhBa4jdeAFxg
lkFE9OZ+q22r+iYcECAN9bhvfmDS/k8myDmriAHqFVx3FfgRsYcmMT+pFDetJFza
ND0BRx1BsBXTlTV2LZJpYZE7AxLwF/CT2Ahmkm0biKJa/x4xJuBg+9q2UKDFskC2
cTkylyGEMpFg4GTT5dyNNyGTC87eWSb4dFNAGTnwcdnoQQsoQFHC4eZqUlryVbfx
Ymnk1Y9/7+fCYJ0gXsosUgluW3FbQ6yLs42jz+MUVkeZ1rkDJ8NLa6N1WZpiaU3O
jOBz3S3t89p3wTQKNRLb4yZ8JM5r4Sw5ixer7YB4gp/zQaw62ST67eJETi9umovQ
dSbxe6fj3xSixKuJMGCIdvNj67/Wz7Epki9NEWOzGmXTp6FhOoDVLYXwkJj/RdhF
E+vkYjP96F3iqoFe2T0hiPwaAtBP+4xOsbZOsaly9IG+sqDa3Q74evjzAnx4qPoX
2ptq54qEqiZ53aUvGkx0ozf0kY63AKMYUSYu2afDVY2ILR21hBwDlb0+IKHrgptJ
VMWbDhFDn5omdSVbRDF4x0evAsdn9qux+/6ppB5NvbTohmgQrWGg/bQ3W+5wU/zZ
ukp0Rhz76wuME01PrNudaC+EH4xjniNy6PsuIwrw3scogUnu1tWJbkhrJsDtxY/l
KjPcdfncE1xRxGuRuZhz34lGyXIRcUlvcP7AxVWJJRA/ZQOPzqowbU2CGG97/mqx
2v6JxOi/pA3NOvrWmDn6ss1DSDiG4V3NbwoWu6ozyIS0qTHKlyuICOjKmJV6jgS1
7papBnWGtSTQC8IY2fzETp0bj9x5IUkaJ+0ZhlXkV1PlFCFMsBtZke5GEegUN60m
s8WyIULz0JmVwdrOKxoyBqqOpauhQ3Ydg5tSBsd+56rz45anuit4dAZnt+FLl0Xa
ZKKbKxlXo+pezlT5HcwhyaTmUKkl++JAdeROkGkmwh06N/9qqgaXyCR595M0ay+M
uYEEu4ibxZQQzHncBtIeW3PStVGDdvQH+TIrDa2rh7WmTQ8zF34j3+pHO8ybi4I8
CQlgAED7kKIBVkJAh9Ed+Wl32rNBIKBAWoRg8p/rhg+G5n7A+TdVfO8QxOBdzzHr
m7izUbI7usGUuQujs98tmH42WhQluTAQpnvX0WIMOMxhClYIRTrW2VdLTaPYLy1s
vAAxrXKt4XlspgPurdqubH3Yj6foOrtm1ZsncLRmWk2K5ZjK7oIG3bBwWBirD+f3
5ZcZNH7A+OZ+bexqOHGtVCKVfTaOhSZUnjvzQ+OMZz2uBCUo9yIaV0jI89XyOvS+
9LZ1RydCpXK/KnWKiztLvpG1gwKDKbceqs3fRk7nwUeEs21FSMk0JWk01nEmz69F
v1WfYEboShKutGSRqzfOu5HYm5Dez2xrrkC2zrOnAKh3cm3WE/dscPLXnioztOp8
T9ahVv8WkuloZ+w9Dg3AzFMthPbnnQNAwW94Q/9AhFwF2HkO7TbjEVhUBiSCLnVu
gDlD4pqBI0GQUq/u58CO85cCuxmKUtjCCj6utYfpQuPPyQIvV/uw5fa1xCkz5Pyx
8cy5+Gctyh3uzRtP/f6wYHIsFtjsa2LTmiR7mBUcOw5LLI+GxA/SAkpkYDeaHZfy
6sTMbzNd6fQrLBnhJolyM7Qwi1v3C/0G04eOH/0zMn9vv6ahRAMQuD+wrbAwthSt
2laaFBe5hxvkM7KRQ7U/CP365+t0m+o/XQ6Pfmsz7LVHrs/QuM6Ud2NrCY1RparW
Db/+P3xjMtkXQqA8JxfM0wpyVRePyTTUVRLJyJZF8pSpgrNRWbgU8C4Ca8LHVnBF
4XPDRtrbiSqAPf/b6wcyKbDOh1HzezxsvJXntu4jkqfLldUVflWC8plHpCdaIM27
tISVXVgOQ5fW+QYujPJ8CAW6stuLo41H4rBm+NqTYXDssaN5UjcEnfR5xz0nKyCC
0ZHd0qp44HHlMlUfCJuhaodcAaNnTXvREDwyiYzVtF/DAm0Utzt2q24DZ/g26vDZ
BuSHjY4aUGE56vWnjEthpNhg17lra1CyPztE08n1K0+zO9UFE0DO9liutp3gHUUQ
Zxz8h/RAHCi6Q02VgJt5+arWPXqvpcgZGTM57BAsVfE9FFuVqJ3WqxN1XQlcCRZo
zSdzSFtrYxQ6l0QGFuh4xwGCbyRiAJkzCkPN9cAwboYdOOJV7FEOeorUUgWc91y3
SpxGNnwIw4BZ787Zw+O2suelHKu2ZxL00Qo3PNnVScMVnsrDgTI3PvXT0jd8oWRr
b1hJ5oqcjvCmlOEmQeiVNTwTxkFPhvv5tc1i3IRCFxziAYen9RxS+Y7aWQ32Wsq0
wyUqBebLVJuY0YDeOCfZIG34q6/mQ+i8BKkmk6FXjYGJsL3EbwgPbGmB2d3bSuRo
Relx1TTRE4AYgcQjPLHY09H3UaVvxXPQSltzfSzKRzr3/OcVFqnmpR7vfGGecrl9
X/ydjQVZRXNudbNiRFuHcgwookJuIIRK3n/DWLCJcvQlsX9KRfzC3Va4ymLVUiXz
4MjBojc0LfQ7xH4cgVyfI+LXFZSqATK1creqOm86P6KQMi4LQUENf2LskBCBcrAN
D1X0n3G1XIRAj32eGRcoRBWzFPrvDIOQ6fxj4abfCKieR/lE7kbJ5WuR5Ka7RUD+
KD0n2mTYN2KqY55ZVWDdtkwGKFUNTiAD6STJ81vOrs/SBRNMwFDNkQaIxuhQQJnd
GG3TgjKGoVzPU8k0GWTUrFAWPRIgnl1lMgg+wxUsHfcS9QKKoq5ALW2q+KbrYfBm
Z4Bq3+hzsGUiGxuzSOLImUqVvJ+Jjutp+a2Fxi85N4WlpsBUsV1Er4FJc1qfcz9q
DPRyJjqeMnj7gYGdnn4v/4MweNkbqJLNx4dFwNvrHwTBeX/VryYMo/0VrswGXWyy
Tfl1bqnD9AIO9vFEGSybAQ5e7U89N+6/akDyT8z/vs9hzimBtv1HGcO9HOULg59G
/Ye7D1jO+Pa//pc96cO5ivocUT1IaG6IINM09qimISsc23EbhL/dDXl61Md8WlSz
WLg+84xMI/eE9S6zTZJgoleAHEYqkCGEQBOO+GW5v2zbv3YVsM0ahLtK+hBLqUlS
e3SsMXKfgEH8G689/35aTwD/HIXfTQvemsqMqI0lc00Td9NdnEmYy4QUSCzD1R6f
VhZmTR949oWu8tS/hWgPQQf6VwqBjhVlrhN8+UsOnXt6vQWXZz0VkZnpZH97lQVD
amnUtTxDGZNmyFlKgelHY4OlMmBojSq6WP3VHuc+GNcHzfV+Gx4yxEF7rkDGwWC3
A2+YcgTj4JT/WOqFDWWh/Ufrqmpmd5b/d8C7oOPTjL1gpTmJHUpgWyQDG90iYjlu
/ZnVHWcIihRD9cCLrqabgjm0GOuy/hjLDys5hfVmbGhzLvcQChFF4k46tSyQjMyz
5jX2JpbSvUqlRDnJG6BpX059d17/f5deKwbbM81mzjv6G5aM4QcdGWx7VusvO/Jn
vd6gn2YAd3HNzQPBpNgZlYz/jV8e+7W5CvCj63J01CezYno1ewRDvfdZLDbVZP9m
MSP3tVlnAqttO3q2TskwcxCil2oTtvbmksOX3ImsVrx4LTeZtXza6wjQ9amE9KtT
3qnDakDz4z6Mp10JVqffN3faiTgmXWLEpmraRs6o59rJLjnspY+6KaBfPzqsx8RE
siAO0zyghiGy8wxJ0Op5vxs4THE3EBErHk2auvSVV85gLk7uBq2tJxW1CxPbLLu/
HTtEqzp78zPNhp+cRiGGkgZtgDdP/6lsU6UTX+eZ5zBQJ9sFtwdpJQAXaKIi5uKM
gy/UtQOj9y64D2pmu0xlEZ+n3mGjzZr/2J89/xKl0JaCR7qVOD/gkKWWtHKpxUPW
0aYyZwQKD/8Kq8P6FcB53uCG2YGyPsJurywVIXq/0n/K+XfyX4iJCFMK/3P3ASPN
Ao9fCWA5FvcCW4B1VMFAOcagG1ZS68s/RpEH548eerN8NHsxtGxAdC+6kvkr+Jer
A9LWrcAh6+hw4yrou29VFc1Vg9Qw82KPkXPJGTQ4Is3G6NBGSeZaJfLdp6XGRkXl
koLbRF7tFdBJVpEDcF8A5GmJkbzsG6IxdMgQn0T/ujUajliPMWIOlcRhUmSBXwod
G+tohBJWPNkTHu3fyclMTvvdET/Jok6ZYlwtzMNDLVIgnj8Q8UuBQAYhJYGK4SrJ
6a+WvyAu+3kp9qIhJ9lSNRvTwBRJptEHLbVZSAdXjiAd8zHVzy5TqBmwuIoBJpR3
bQo1Hyf3iEAONzIRspN9DqTUTR+VVwyTDGTWg5n5U9NMBlALQ3kOG1tNveFt8dzh
+umGVPh+PHWTjH1bFgW5ZL8ktnHyH5ywfyC2xgY7W0nrRk5lRMHfXXL3A3zNzjSk
a0u/il9cPrfGgU8Uy4m8JtRwHVkcjZROJ5cEwu04IvyWSuMjuTS09MfwZgZmXA54
kJ8CBtBfNd93V98tzUpLyzUBjvmNDu035v7BzF+SNWxoeY6JlQBYlIgHeHNYcu/5
bAOm4HDLnQTC9peiMtj68jJ6jaClBWGnlQTk6VK2nW9d2OoARlvFs20Po7odiKoT
`protect END_PROTECTED
