`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
60i63mWWveDRymI58YoybczZElI6DpmGPos7O4s+c6newi2htfDcitBNu51mmrlF
/f8Md4UO6RLmXUJR7pUWw4tGbJBPHNjGF2rxKGQUDuKsc8SJDPb9GYMShfr7vwPm
QcPhBiJpcUWMCcvS+5Obc2LjlLlDFG2Bes6OGIa3uG/hWkWjfkhuJJ1o5o0eCPiR
T/8skrBfJsbAfkOjMbjfqkenk4eKL/V9Njb0uIMbvb0nRSKKfsJqYaHLDV96MhsH
5YKyYNCtduKmxrZ9LUlz/DzuzzfQnvrPPf+3TC8uX/PEsm/43EaY1QesRptYip1w
CqjyXBS7l/hCAbPFrKI4wnpx7lvqRZ+HCd5U4qfYt9UJsSSUC7LMJ4JJOLpEnmsZ
`protect END_PROTECTED
