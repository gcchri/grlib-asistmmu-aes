`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/WLMkaQ0txBrXRyoQ2Sp8q4XmoF9xGqNQQf3ESeBogPampSBGKQ4VSRsuX9ZVKoz
1tsmHP8O8Qs2fKWsmt5QRXzFtVlKDQhZALF82DDUWX9TjcWLrXet3bCUYw+6iy56
/Zyg6JKsWUi77/TLorzwbmHz0t7XrTs56rMs/FuU8wpAlXLG2wx1BnrN/AUp7UCz
sf/QcbRD25oyrTTOXDfOLdjNaCC00CYQannGD5OPRAX885eCzDpO/r4wlePxJyvc
z7sr/sugtzjFoWoYu/crzXMPHA/Ra6fL9BF5LnwNEnf3EuMwTHsAGxJgZd59RP7x
p+lNxJhoHl2hCJH2YOHXNXh6IZMzWob7u4dLatg+DIT94jR74qeR+0IsobAYmcUD
t0J6Qb/tMB+KhhxgE7yLa9d+MQcS+NAN1Hs6sjBmMDhfrBVa0kyMgWgpLyMgJ4KG
Zi8BXGlfI3mhfGgPV1x6z1gX3AOZGbOSJtpUkXwsU/cYAzOa/zwBI+xynbzMi27A
4EUgssZ84zbam6d7Q7qSfx6wvtjeUQI7EHGw4dypqI5HPn/0aARiwB/5c2Ac8rmg
bT5k49kdCbagj66070wrw/M1JawUNdOpSEw3T8rEAyt7lLi9YmQERA/FIyD9Ns5u
inNJZXQclHoIr1NT34Vd5Ko3ReWzI48tS6S/Q9DjdRAjPN0v8/46X7kcmTXrhhom
nt2ZNq07gIAUqhpOMgc6ZlxOj2hQ/omCFw2eCGVqDh2nv8ZtYnto0fTLZwz2STfQ
XqqBxtVgOoBZJcYmnksHTw==
`protect END_PROTECTED
