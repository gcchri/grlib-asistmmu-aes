`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KfgjhMEz9DvJHattg22La7fYjvuuG66ZdAC2vAsuVlHJuyqBKpYNm0SRWBu71ao6
DHteE4EzJ7679sDmNGw80Hf7D9tuIPVuRtYoI4WY243VH4rUuZZXBS5f25G7bE+t
uCS/5DUDi9wNE45e+SdLC/F25MtPg+xoABzV5TSEH+X0h0Fk9HHhcsEdFgtItUtD
qSkYyxHtITEASL43OpIci+M2gCDH6wAOx3BfHL7Ez5Iqm02BEzPVvs8IiAondybz
AtOO+2cJ2y2mv8lyBCQh5YAsWaEmfwZQI/FYx5yK/nf1akXJFomfvmpisUlNHspE
G/iMEvxiH5yMmeHh9fk1DfGbdVC8M/7Kd4an0qCKYGhTm76GX3t6AgEvps//i3ye
`protect END_PROTECTED
