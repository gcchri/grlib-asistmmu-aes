`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E3w6HOia0uPX3hLgtzUVercdSLoJJ1PX63Xcr/uao0inR8pksn9mpkjHNdzj1Yof
35RLaJnx8rVhNz00VGGV8BGyNRKbHUcMJNPZWLpij3bKPlmLwyDxIjZA2ZNKo4cn
lSp3elv6htZAQUa12B77fRd13mzLM025OAvfrxheivsl/J7Abx82td9rzWx7voRq
PhUAeAFbCWKapbP5K7LGqjGRHbCi+FMgmL9zUmgz7m81G/HjIRBL5x1wqtbhOYnS
JghLNxEIcXcVyTMXSC/IuHyCdDgw3FY3aM4M6iYRQDA=
`protect END_PROTECTED
