`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
evJqGzDlWucVqcM0y+xCinESg4zpPQvqRsUojJX7eYALX9zFhO7YNPe8Tsi9ei1I
rXN3qVCHvcUkjHlW/0s4FTKJlT7vLtFh/ObMkN5ooV3JNKE+sVL6Gv7qPjup+/bo
c/12ur+Q+awE6a8Wx4jvJcamtoNvsQtbGGrbV5PNlcuAux9dInPnc38mqnsCOFiP
b0BJ+TM8szfNqhJmZQQVsQZ1JIzUJ/Xy/UxhSt1Wokbgh3Zku/1GzV/JnbwZX735
qQbaAVuuNyPRZOkl8YXO4F2bQRP9Nm/sZHVEDJuXAWeovkZT3Y0Q/darCorC/s5Q
42upP+jzQI/pXg+R1vcpy8dLMNMkBZMgtDSbvVC1n+N6RhiaLuhTeqU0Kb3iydl/
nvRs7jBJ57eJmugS5nq8NDFUs0CLlzudHtVrky7YL/7B6vMvzUqm2aTsBMGJ31uk
IJyIHdiyDOhnDUrpTVhTwftOFmOJ6ZgehgkODJWd0fjaeBlxMIMDIjkR6FCrK1qK
TyUi194ZZV2R7YkTR5k4djNk/Gwm/VpN6WSXVWDlD9LReolwrtMkNZS/Se3BPtZl
R4q8yENdOMiBgLQ/MXG2vZJ/dHj5c6F29wfgVbYK5o+CB+Xnk0LjBYKmQ0l0lxT1
QlEBXJahN1WZiKSedM600A==
`protect END_PROTECTED
