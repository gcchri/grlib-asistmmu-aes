`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F/UVgc4W6IG0IXkKW3SwVHryLIc4S3WcudakY9CVKpj5ct+hmzcwfyvditHuGHpw
AnwnnXlkz7TR7AdGfodA5oJPa0czUItz+IqUVXPS5QHWnnjQJ2tjE3Oe2pVHCYgy
Pq5Ufo7gdWgF8QalbucTE01y3UgWmIBlk2ip7OdV1TJdGZlS2N70Bpq3ss4HOt6Q
trWiG9P+pGeyJ4ha0z/A88R9rs2FUxpItTFzyst2rgV3udRUcVXHoNKBsC5rHQOa
tWML62cLTPNiCoc6C5bUjCmhVPBjXmWxOqnfcyYsI3gG1qzCuXx3JdC97E6mMXxB
lIlmIxCd+G3X18zGf3hAzRS/ASxoLVsXJaCSGmLE1TfpgzRlqf021lI2ElZH1xk1
Za545WGbSjgw3JJ+vnI7ouRYWDRBAO+bKtcu4mib0htb0ZYT0Vvv2jTuTkWF3CJf
Xbq37REKdO33jWLdKkriJN29PeK2rFbEWwzUfPoi2bLn4N44rEp+UK7dBtitbVIz
UhE6vifZKuX5ViFu19KiVS+d4rHWGAPqnN+aEmf8777kw0wDzh3RaGo+//vq+6XE
v8uz9WJWJgG1nezdFaK+bixnKDBoOXZ0AS4xSD3y1nXVYH7s2MhUbaGZg498dgNN
ey9jc5zguYuOp/t4hw2YO7MNie7EncFFSDq+zdHcYxJxen3LZfd3vBzyVaOSanxX
LJB7eQ3h1Ix6xHD8rdPIRFEQzdHekb80ypMjYo9KRbAsxoSnZWgy1iV2rUMjmj93
IucGsFqgG+ewNCS7b10rzO/3l/xM5rmGavYaHpzIOlVBVBX7aVqkMMuFx5Cp9O2M
dVPq0lMh+E/jYdeKGgwxddITUwgznW6Y7vWewrevQD8U4qjGNUpIAEUZCOL1hJfV
wsUSaG2FFgwWWBokoTAcTDvPZaDldTYflJK+P/PLsPVvSAORRIKWQVmnUZ0Uk4O/
61AtwAABKeAyvq6eY3OPbHeG8lZtD7lvQ2/CE0P7ffXQ4YQVt3krz0cK30y5+eMU
i2Ol58/FqsT4+9+GXHkmiD98BPhFQ93kAew2EkYrkRP0e51+HZk7k4YmKT+xQ0aK
6WZWfFZf9gdTRRe9MNZWt6tbpua5Vf9A0Ynm2gV0B9L4WA86u/3oC4p7bdCGTvqL
YsNUuiRPhfIuHlgflIxgtN0VHnB6orWuSVgK50wCS67kkCZbvTDhzt7JEhX/65Bz
B2D79z605vQtndBWGhxNtJAXApObK6QQAEoN8THIIR5/YSJiWNeLczC5NY+sn9v1
iZy2xUJFuxIBggva9UwHdJ+Vsj2QYCY7y1j60yaZI1ui10ZBd/WExry25IknQcN+
F7gTVR6Xl8xF+Uo4RA1YF04Lzb03O4lkjf23SexcG2gY2Xbgs9yBagrWb/2wZV+8
b7eoOUPds1DqBF1p9YQrbF731WqUSIM7V4u4TPLPSFwng2I6wzyJMrz1LzZV7xmz
5uqYFJzSQmBX1aHpFy4NXaWa9YyQO7Q868yMi9CnqQYJv6pMBWJOMdwquhniyxeT
wyzW0s0bO/XVnDIW25fASRpkdG+ixgD8hWrU50d5JiOLSp6MpkcofrjNXa6SWcjC
LzBH7N/umtJWUDJqEwCaTF/Uk2Im58fC2/eQNX2dZ8woKtRHfrGpjJgwUoCM0oWK
V9n1KHv7rEy+KTrK9+A+xdrWOyRMqmJX+zbj8WszQ7Fam7cNOe+diXydOEl8t4rK
GeFJRbllh4BNJgFAHbdzdSvKKX8WUPcBya356kFp/QL/u88NpULKdMYj6WyTbtKk
JwU3f5j/2Nm4pKorlgc7gt79kq2tATBxyRpimSRoGy0=
`protect END_PROTECTED
