`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rgCfFnz2DnUpzeqrRnpeyKiptzaAh5TCs83RNBMHd0d3S+D6+kKMtjUs9mMUjhAs
sfakO5tqbVBO6R0Yu2pWQQarR8mW7CyIjupTABRe5L1+RgFoI3oNmTjop9fsdf1N
w2IpyrUcPq2NM34I4w4uS2iLlSDJ6mbp2shNaDHtyyYPzNaWh/ggnXnUptksM7cr
ZrzBMpj33f/G78RDHZ/EY55+LSwRADxyQdtL63EEBGV/wYZaDqNbNF6HdnUWhaaz
CviywmjUhK6HNr2K06sazC5B4pqgoiTXzXwi+EanHwXxblJ5Quo/Jc6TSQJtWhNA
hDrIz4krx8rnRxvdaXoth7gNmqluc+HMNQSGrpspygl7IzKjGkYkFF+13gK0MDZw
7S/GzPcpqSHkZEjkjt4VBKxcl7cIywhpBRMGbRbFqwXdJLnvTZE22TsoSkrPcsgP
dH2kIx2itaX+PZUXSZohwFxTf87BijqGJuBLwOY8SoFzybCW1btPZmxoLebIZ1nN
sOTV4yVFtZU1rPhBe4ZwdF23VTsTeq1szCzjysZWUy9DyMGvEEDAT9WtAM0GoOTk
WcrGIWJe9RMbhNm4+c5t35oyrv6MKnRzaul30sPZKn272fADP62cyz7IHxcgjaW8
3VVc6zvYbEgjhlR/7WLCKQF1VqGFWQo7FkVyJbbJTwEUpYFyPsjCviyutltz5lwy
7Sg1v9O40ELN28XbnSJ+TVa6qHypfYEapXKWxyy86CgoIBH/Mh/rzPymTPOIPvCk
kGB+RS0roxu5SqPwucJfRWZgDhzuFR0s20xz1/BhbvJcbeJPn8d49tu/TNjBdCiI
YI+PqC8eF4RcJGaSTEe3ER4Svwn+192i/SeesPjwfyAPpQa504j8SbEkB+srOZYs
Vo+lE7D8o14QJKOvXcvo+jxSNNZTMSIuDPfem4GmJmZogugPjoDVBUEHn4yvDkJR
CUj4BKqrK7+3IoRy2wWFD0OGhu0XrrTV9+/TqgfrtAmYCmTCYWfXduGBXHf0up3w
K1COplrpbZ5OAdVDI+SJ4dMRavRGGUx0R6WruwdEuirP+6Kf9sv8BN9HGIrKRe7u
2GwE3k8Ch3JiDFcGi/rteN8NifRwcQt21tZOdoIizhM4q9O8kayysq+0lxFIx5fP
/eOfbE9SH1Sqd4DUEjUZXQvnDRMQv6nIaWsU9XlycL1jCO5LTD6Zwq0XjSlNPmCy
yTquzf2tRSI3aopoyTdTxNZ4q9CqPOQcgL984GmGYRvVZGxyLWnb0sjXH/vyuMyG
zJGJDVv+xpZ/Yn93Ljh0HFweDPQJBXVQjB7VMMn1jUPUZvVnVSGj7M9Q0TbB6CJp
Up42z2+pntRaNvf3FqsJLjJslX2a9h852Pup8vP7fjQDZdZ6YdoEj74ixQZX3JZ1
L/EIT98d1DHMB6p8D8AEkPtB8LlO/6nh5hLiRJsfjqSBqxt7lQOffsiHjWCCC5hm
Bf1BAg6LAtdxdcNo56QnCp/cdlhmMEDFiYBV29KerggkVndqDVzi1dGE7azO06WQ
Tj8+joqzx6TFXWVTgddohdvNMvKjEecIapHkeK1OXEFgnT8FWSPow8+nhboSbG4+
JOfzz3ypqsY0lUl+cvHLS9Lfq2hohh6G3Wv8/oXDx14wHjYiz0zZ6i9MeYT5+gA3
3NaMxro6qUiCndMNuCpx2hk+3ERR/sDEO3o+29K9rRF625vBU0KITTybOwxjjq6I
RL9+JeE9LW3mPCaFvYdJmadqO3U4yQjGuScmk0IXno1gjeBpqjDpHF9uIoI2/97E
UzWIjBA6vOyJJQlEWOBwXK339gXAuhr+URbN7H4MULo=
`protect END_PROTECTED
