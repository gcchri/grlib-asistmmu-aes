`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iM+xKSDY/I3QVagGHyqd955FRMPzTZp8txEp+nxHvL7x2+4O1sWltFC8+wp1uXVS
1bxNaxQWWq7OuFDoUJCxVslndNKFfL+S+b6gQ2pGiwb9/QibXntcrCqUYnR25XRc
KneZHfEHn4zFwFhJTkQkYKtB3DZ0X59QN4w9GlHW1vXnnhzQNjfIf8kbGiTUE7Xh
1GPJE4z3fWZ437TdF3Y7hUmHEfx/9VQUDrRlP/oNekuJiEAKpUGhDdZOxyJt+uSj
tsLGSP7Gs4oAAroFI0IRpQ==
`protect END_PROTECTED
