`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D47BAgHm5zPU1Hd6MMTVwR3SDOqpmOgsI6tv/Qz3ftTs3WlOxQ8M3b5WnksOryxr
vCJdwnKfNmFQNWa1nCggpnYgATWPgURUVhDJYSYThmYLxC9X1u8zaQaX9fzEo6j/
KuMNr8snDYxU9eDbVDB34GsX8qyf7T9Lfq85phCJYrssdhtSNjlet2oToIaK3jGR
Spz7a6cGrghqGzIjVVjcFnjJ2XUx1sNEi007iC4Ns+rIsNzyZNJoQtyECIY4jKdB
w/EWyNtB3MgSJjXF09Bb0iPB6fzL/BIsTOvXURKWVDLVaiYEzVuTNU8hGMQueCSb
cMWpLg9DiRQspZntlaCA5QhWVHpLfIBn1HWtWRxq/gvF6GbV3ouMYoEpvwa0dgs9
`protect END_PROTECTED
