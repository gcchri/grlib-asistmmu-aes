`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LC+cD85Q+Ta+uNZEOal9bwS6VPFkz8kIMXbEZwFEOWXsLP5gEmuqyXsRkUZSGNje
oL7BBjel9Ax+gawQQiJIVBM1J0r6svhN4jjttLl90HoYZd5nnG2wgNGBI2LQSjVP
egvTQw0yFm9xa7pALsNHg0E+JmixwhPpdOlf6JDslPQh4U6QNGryps0og5XH57/F
rOrvogcVcgQZcVFZZIz/lVSfCHC8tccxyxS+Z0Y2IqL5zXNPqESIF7a0IDa/P2t6
U+ndNznXNLpLAoojEiBGYE80Tvcx0F7eDqK5r9JYFwTGPioDBbkWmSa+0tuJe62t
42z4iOql9BggF0UWlN2MUNWEuvYJQFP3/wN1YaoYzhRkf/Zabl5aE3aYV0rrdxqE
+Kt43AMeFFckAQ5vd4Rz5QJJl5tOMiL5BM2loPLHEYVp5VTO0L1XCbUEWB+rWIfD
qKF8BjGZXPIyBcwWmOjn+ln/b4VyfDBe7KBCvDlnFvPLdogoc7Sv/9/tazAqfo18
`protect END_PROTECTED
