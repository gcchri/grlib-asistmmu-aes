`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MFj4MUvg4zyzDAOL8gytXn0wAvkLu3RhgIpLpPwNPkcVws/TFd8PUysNpusaDda0
tG2Oe/e05RKlAjlJfQHu+QpGrGtOns/XVw2ewGd9Yi0pwKlV7npUoxHgWEJlW6Bx
eBWWvLAHWcOzbSeXHlPkhz3UVkM9vMq0Adxhv//D9br9Z9uW4BRXUvi/2p8VPYuB
e7+k/99v+YkhOZLqhWkuM0LKqZ8GehThVhgGdoUYEeH4d/wLF3bkmcRbLr2f8aap
2NHXEa++SsZwrTsGWYD8NkZ2RxuiWlym5UVLcEMuGQeb+urTTKwj7xVEgneivrj3
w1F49i1P/Cb/7JT/QpJmQbccBdW8CLTOc26Vy1u4ylnUjhqsyZCVvMPsdVdQevZx
ITOUiS1eZTBYgF3n5SVOJ1KsbOR2kX7wOhrRCUQK6Vuij+GMSSLhWXj2qLa8lwKH
40uZ7NC0CqcPAfUqnZmk0M65UGP4n1uds92e/XVBjnqwzAnZzwrG0oFffKffgZuU
I2TAuEQ9g3l0A8DCr1NDjMMnVg1Ww0HKY5ZfXg0Nbs50tLZUBOAHUVFNmyW/majk
eOM5uXjSpCVeU51Hap3v6CZwpBUjcGoO1MMeqRMVeA77+XQQR/jLkttLAG/K0tKC
eYxcnbXVSnFFuDaLHY9TurDHOlR4mUmgkP8ihpeO1eeHsQZTmYCtSIT+X1ZRaCR4
vwkXO39bSoZuT5Nai/KRMy+rFrBWradcPjLPShaxIJERk6Ho9zLtYBidDjEI33S2
/uXbnJ7nUk8ikb4kZ+oAAlM/0QOhXrlNaR/d4+/pOZhz5WgzielILrB+1zCiBhQL
1kr5DY1O6lY8771TqrKg7+msmssY0I38CwUzZsJNPpDvO5FaC1chMr/+/p9s3DmM
S2rtUgnCzuyH2KcwI7Lf5u5dOHp+vJtBsTrAIq2tZi7YCaiqvIl+DathKLLwxZtb
Tf162stnkBIrjI3qn80a5E2/tcO18UjabWy1uTu33UqxANECEyPZkMlQtTFihAGn
m1zx5TCTGatNR8pie9h8EmOaZC3HrivtUeTgQk28nitxQR1J0z0G6o0uE7vJlCrK
Mng4uwWriefCM8xquwUsi3rojsSgJuU68qWBD5ykwbBw6JjG56QUu+5217wO0Jcv
NckG2GLXqLy8ph1IxaAvnzGluLDhdYzy7shye+ctGZg6mJGEerl8+pZpGJBiYTF4
1g7w9lyX+IcZk7lHb3QxvjiL0OVzAsYeRUBogiDuAPheqfk6H0yfIx+G74ZxgOMZ
cvgxanwFyAONgzoPSkB99NJP8DT7jJAETve5P8GVaY+12pancdyH2fzhK9vfQ+LS
jZFpGbKQvstUFZ37kmaHvTPINQUhlGciSrE01BV5at3JVVJg7ntDfDnwpFsKeCS8
1U34oECYGX+MJRML/xYPVX6uutGmtkmLzM1ecXwoaVBbE3SQFKGjDSep8RW8g7PA
BQvA/5osuX/VWDR2HjvnXcoVMQOm7Wu7YGZjOK614Mub9tBFiIJRQeHtxR39DMXN
3TUFnH7diLjLCwBr5K4o1qnjMKQnEpSfB+yP9JaPyhOz2sQ01sm8IYKed2ZpeOeY
wjIHWl0LsBcel/GHsaKpSFxJhOzULzWmPk6HhtCuz/TBsuXdqYz9vsQT3jJkGdhU
811sVJqoSaMPu0XsTDMMMjNaggt5drGcBsKerH/8ni82gEZsIocUS0IGYXIN5tAP
cAATXJXdOKWO/YcIwUjW1yxSnBBDBnHVpMDAQjJJtU1oNA6OU5nzcJyAKWcAvrcq
W+Uh+zTEfBZA274AXqYbBu6xnOAMtdpdTqcrY8haxDfpm3owVjIOnLDbUvIkl2cA
vjxqiNm+gc1sYdMDUoYh9SalGgoCP9zzcZ/nQq4PUOZtsEjD+/5Cmd3OS3AOibJu
5p534Psvr6vi0ivuYf6e22ukIL59IGGZjQGeffkhm+0xCLW7VuOjvWFWhiLYGpBZ
Evp4lsO4vG7sVE7CGHrxLhIsZu2PKDJQa3mBlNeVVPcxQa/42pfTmQH2lX0FIrwW
4SPRjbstbFVjaB1M/iRoCPeve3gOJRPJmXMjb+9mqM4fRilP8qBL1oGBe55QY/qH
3xhJOAz6G2rCByxZwoFl+nUGownIwYapDQBi1BCJ5y0Kz0R6nWolNfqQFMMUJQI8
eZ6+zOqQdeT5InVvFbEFhqfdJMkO27leEvhDR7mMEYLp2ine/7sYPp3J/FepsaRa
HNdtWUpgRPaHI/sgQc5rNIUX1ilP/Dpf5v10qy9V5hZNjn+yI0br47beQTkljah1
v30uIpdv1zhJS4e6TEdnquYvmf1F3SqLGIuBC2NbaelyaeM4O3b0+zaccfErxSUS
2NgcqPDZxx3EPfCQrQcliJ25BRm7s25h6BDiDt7AeVOTKP6BXiGnsAYRDWljj9G2
aGYOKT0vodmFBEU8r3cb0n843/ab6UYljH4CHC+XEpMgOtpuSWiz6Ma+Z2ILgsnk
90BfNdNpdcKPC6aTvSC5ivCAvN36sd/YlYWWoDkRuSn4SYhBOV+RkON6NYV3HtiI
6dCIpFnPqh4tWvPGG3MrMhkFAGG4FF5IXPd1XRd6kNIimmNQTfr4byePyfyeeII0
WxJJdDzuO3ZHgXp/p9U62gb3fjMvmQSJ1ELVE1MFWh+bXPdEuaHDHMpQsEh8pY5P
3C3aWhAh3TIoK/jMKzgyIgxTaVhKlq2ONiEkq115eow8ZzsVQyBbzqh9LFrwwLl+
znjjEdYtc0cuElvrmiSjZGmsxJ45BLKV4X1FvZGK/Tr6PHIGHDK9ndcZUFGnAKfK
MSp94ExbZeElcA621/yzf4uWpwfWU3X4vUdKtkv5N43hQNelHYUCkYPiIAJmbDu/
53El0OFXAIMpN15jk3qsw/Q32MZSwn3mG0xlF7czWd4kzAyTwe0gTLYS2QeIwxyF
hvNmmlOiD6Cidm1ooJIFCBtFE5sLiYByaa4BRSvLe07sw4sSsEgyd8wEkaV80RsG
5HWDZo3V1i8DuRy87i+08GTuj8av0w7VoLQd+TGp+dQbx2qEXfpwLmmUwzZwGMx1
7KB/3Nbu1PSyv0+nP2MxwrHytygB9qCl1TYUYzYYa6x1dN6NZwHRV0NriCfcUmNf
2KvnsgJoAVYl3T1A8oyzzPSYkksEgvNjImIxGqPk4m+bNYInrauvawV6oT3Tv7dV
CUWp9LDsApkrc1ydepUMreC/iupjY+m4vsAT+CqDI3wlLU6VlYVGl3lZqp2SFugT
WOb8lle4oPeBRe0iM+ncQOGJlxj0QG2HTybHbVCV+o66nqRous7YpjAG4RVIP8Gu
UKR3SADypXGNuOMWJwdFzgVdfIj0k19vajlX2UZ5TBnRP3KCNQFeZllZ8DPfYDgu
8awV0tSMML/N1tIhR6fnCdDQaXo4CSLe/YAYSZ2Ii7aaIkvRhe46FMB4VEl2o6Or
+KtIgttpLhQguuhDssJffT2WmF8q9beggMXCFQdhyrX11jj2nQlLMFpYhieJW5MH
Uh9w3vgVIHMlW/TBAtjkQd3c1nid+cG+jIXAyhFC4CaTbmOssjVx1PgndonLSkfh
lB69x2+p+M+7x+BmL+4gw7cYOdYcEnwb9Ajd9aoErdGwlOLQWNesDaZzvyrC8Mqh
Z0xTeatTGlHe5s1bJKrxENEct6fV8FO5o7JNXEYwF5FX7LVqUKEdAecJqqSMIFB7
BV4N6i8rMxY6noeq+cGNNNdifiYzxg8Bq3TU2BZ5vT1zPPLr99qmNLVM5qDeNcdr
5E+K2IzIttw5u1r4gSA7TmHPGGm2YRpqzl3Qs3zYNEbGu9i4x818oUXzbZYNd4iB
588lOlH3hLEVtuDxuGFuWZ0zZYRTXSHB0AJfuz7y/hsFv9nzT6DVjjigLRFEDQu8
5zi+VXz1DT4zOjD0XMKT4VcHTE/eOV7cH/8cOooQoGPrLKEyqJaAygZchpw2FC0A
8mthCKrc8BP3f0EcpSB0vFOQl0py+XgEDsG0JmKo60csVI2y671D+fjEA0wwaoUA
d5ImDYT9iMafu41hmWt+SBmOXENepEoOHCbIC+9i8cpjAYVLYmBQCwwvZWqSNBA/
ZiD7Zu3loyYcBmzVRvikyHknVWXnD0iXZ0AlA6jhqBTNiHlhLe6IO2GDoPhPu9K9
WnXmZ3tGAxxWSOHVFbWUkX6PGIhsqRrillZjnkrL8HrrJcH7m8JRKtr2MgUN8/b2
sVAM/H9jtS9ElkrYC07RkmA1ENgg2MsV8ftUmcnYB3so4D7ZfYIkTSLccG5rMem5
JVD0d/ub1Jyw7DRNnY96kp8evMhcS6AUusHSbqXQHGhd4R3zAXxwi/BfM1qVc1gA
1kRMMrmM9A9V4OSc52o6PpmO2dRnBZa2l7UpZKIs0WIn100bU25pK1Ddio9Jg0Ix
ATtH5lKyIGJQO4PoaHk+ZKH9GUlLQ4I+ooAS3fn+gRs6W+1Jz21vbrmgCMIXP7O3
8iMJu6gKofdIQVXjQMZsxxkgBeSNJzuZ74iw/0FHN4mX6HGcIeEg1Ah3cPpE/owm
z3dgsEZkxhkJuZH/pzZJVg2xcZbO0a4qJNZ8cvOAHkp0ZJZNK1mXJmRbOxwgYLoH
uQzHnj8aNQFjsabbXqXZUItl4Cejz4JOIVrb6TenTnyKTm+r7s08sir9PUWBeBfw
kwfCVdBj7zWSsw1y5gOyS4zy/JR9lMw7WJ/YdOfStY/NlxerTkQW1748SZBxo2H8
vLBn6D+HO5zkZpl7uBLfl5ClU1rxm42e3UUCLWmN1fe9OMmeEgh4ADlNkKDW595w
EIEFcTcdtcGsDUG5JqIi7bpL0n949hqKf7LgH7hyspgsKybObAhLDeR+rsXBAlun
G2R9Ic7PAZSPaPAhN8qKNrCW1AP1kcl29dotVXg12fwJ+xlHVnwgHH9H8r4Slwxr
HvmiA/zbGzIJqaRkfTBCi/iUwCVDgIbrz2BvfFH1nVx2JKAxDnDpYLdsopJ/UZTA
obEsWXpEzjQRy//Ry1XXmxCOYcruV7M69dF64v7zTS2gsru/YKiWjKVaqsO7dNWK
5yRHgI8y2n6XrlGOV80+BAbA4MfAvdOhWoff3dJiewc3vv/+laHOvKclL06WxD8K
lUBu3qd8vpCf5Re1b1VBQ0fwF98H6oiCnb9g6V++JcuGhY9wiD4i5A6fxuVP4rsX
lzgFWTheMySRIj3y0dA8Wg+mjKADSfvjt5CN8XKnLp5Jab2y/ZmjpXopkMQh4VOK
r6fZMgZSBzSa+BFxKNwz5spjSdg9rrJ3RHoVjVVY+K6RNQ7ZK2270loWK/mpOeb3
YGS+XFCOXJOYh0Obt53cxxzbkUHGcKBm883n8e9J6t98cSYAgK/32dwmkslqjR0s
PErdFQHAgAHc2yR/02l02rD9PeLvCqsaoBNS4qrd4PB6T0AGn4UO8qXGLrMNzIwP
kBBrqGj+/PoUmp0B6xAmz+XNDRjSrdkH+TvdYNaGTN0WFv6qfasFuHCgRp6XlIEv
Z0xzvIv47NAG5svGOJH7PXohasEN33E9fS+nVWj+elojrmBXwt32Dnk9ov0R475F
os19HzH9DeayEPiIbPs0vbzF2BhNgIypYnAUYURqQiP6C+us4fmk+qxoPGc8KwaD
If65L43voHjO46jnVrAVHxjhSRQjsGats1OechA5FmeOA2L8udhLt1ZB6eP7eacC
gTmUHBb4O7/gcbULX+x6iYdgE92oW4X9ESViI4f94+Tcj2gSt+QN8xhDpRvYLhB3
fQx/+cPzrfW+cpG7pEM4nWz6OLvzxTqxnslI3QeycPB1XcYw2jW5PJYje8uBNw7K
otB956Xux1n/XvUCEzTpuGvgkFuyp28/gEL5pfK34N479yrQp8fGb//CbjtFE21X
UqQSLka2bC7UCELuPFnbAwpFR1Kcj43hxaQzDHwFcFddP69OkbIeCIKtJDpWu0ii
PtU/bLWUE5WkVd0ERENfRjwypI9G845Edrz7zUVh67YauhDICXFnBFqME+KuW7oW
72pFK9l9PvGTeRJ9dlYq8Ig4LJW+u/zGI+/2F045wcsTTKaffaVAD9kcsMWtwrfF
ybFAPHdk7RowtHLKzhhrTCZOjdOfpegcfpBxyiB8gb/PIXQn6hSBcLYZN/smJBnO
F+4sZEWqwct59FSKOkHgY64gxgk61Cd5LxG9otLTLv1Gz6+lvSVHk5g7BMMkoG7f
8X1ifbAFSZ7CPW7swZBkqJw3ibkIG4wCU54OJcCL+ipF2Xr8akRhVOrVximQAKn8
Aja7Rt+w4DmPdCpiQAvBnyam4GSjuaDuOFudCtsjRZCJaRU2ZjcxxCQGnxU1O5oK
mGxLyL6D6gsTKKHGK7yH0EyPLqkm8CCGTGy8+65nsvWL+QG3q/vQ9gnFTOFrDL6K
KGA5Y/HywFO081RKbOmE2p5D30I8KNk5UYEY2gZ4/Yl0GQbhvc5DHPxAqfM+VnrV
PQMwPfESoRl8ln6wWuzEgkkTbmmZM9BGqUgT6bLK2yzLR6p5c2jLu1PB3bPVjkOP
usfIhQy0uj2PJ955xSbVkIbxTPZ0TtTrb99vOuFzvqWX4b+GDLminQqRuXYuD8/l
px9CiLEbU+D7qG2Jm85q6/B6Y05URgI6s8slEyuMkWNdOuW0+TGMUXXKM9LP3lgi
+RRrKa0zib7xtGbkSNbFTtqnNAXJ7jia8iwMsNhU8w+qaDO/Vd8wbiO5uU379FMS
BED6g7iCSu91wlHKYT/9TsG7zdJ1bOpsgiYg5XmemUYLxdVSxFxhp82cWSEoLm/3
r5dEcqWFY6xzhASHZa8SKY594Lmx5zKY0S6nWZDdCUzyCDME+GReNide/pCzMSoQ
IoJmVLoz7MPAR4RliTdchB8RiWJnbNcqlRFzBP+EMKcoqC2yKd/HhLknyY7Nq+51
J2NCyHCNTXJ4/tZLGQiAXfLzZZJm3isvGMKJDXGutGpC9yLig/+xddpir+mc0Cjo
MxHn0SNkTdMCi4eZW4ilT67Wfg6I2iw9geWC0kueuFZenQz3eBEj4SViNiyTcT1i
zqHE/Nj2m/e9qVpZ33S87uJlPcer3mXpbdb5LxsJqW4qCNWorl/83NA7l5PdSTJA
gAwtaart8Tx9OXqQUR6M1JGSaASdik0+AOFzgBQtrOxF827tMxRyE5l9tpiegfmT
3BztaVw/sWXNpZ3Lq5j6kVPUx1kjCmltQTt1KthE+9aUkPzOJZkv7NfkpUjVSiHD
3IWaDBi4VvZtufm8tS2n+edTL3J8w0V5gkyylucvafgae78Tr5DqXa3Yzzglxx+F
c8XABbB+XRljdcWsLcx6MmnCiwQOa8re7n/qrO8QYsEAid+zLTuBEmm6NEAveRCl
V/aupw9QqpB7JXRpv6hPPcf3QoPiU2eOjd+0t02pp6ACCviMwnhoLJOKL/FZ1WIk
WBUO+sYoMibZwWmLBLbIfmhpebx+5+LXYCC90rGd0Sxardte0fJ1mnGb4CyTj1Tc
rRU4RU0QBHV43JpRgou/hgaODh7YtcL1cJsf0s2MRkzyVVuLpzpFPVNDbb1/+MBJ
ZX+C44lVvDmkvf2BRG9rJ3X9eWBww6GBS5lImttHhvcW9iVprKsp2pdYCLHZslD5
+UHc8x1JETMDgAfbgLgGDbHX87IqwQICzefdww1HcFw73EQhs0LZJCrikja7txtQ
YYsCxfig1Kk7oAUWuPBraBNQMy5vlHfXqKdDNw0JXkAsilrJMWq9u1Yx7gbBpf7L
7IwjjVoWVETEo+odL6xG60avjdZtTi4kf6MO9WiPrbBZBC1fL0fRgtt1mkbAHeL0
JKtsnBdLg3nLRkJ8pNozv7NZRp6+NZP79+ZtZQVzSYj2VJ9cpTMlDM2DHQIEor8O
pXRpoqrZ9s7Z6RxN6REmPwbn07ZWvpzZXjY4AJ2YvQiGbdUrLPd2uYJ+RSLJnTiG
HzSDEFjj8WT0JoIFgbmiI0tsVyrvO9szODqPYXD34ZAWpOclcmOxSQxmMMnrcZrk
+/2y88APD9PwErtZQzjtiLqwrfSzAquwwrSWT9nWOkKleiRos2wMT2uAi7g5pOJr
wU8RZRxU+Xsyfs5nDDYDk6Edp9G8tYc7JaaWYjVJaAcgsdEJ+NRvPXrP+LtS5FuU
VHBVoRKh9vjsMeK4ymh7e1mIVWgrqf/u8YiPeDbmztw3O4hi84T9e9eDj17aLq/p
VNBDBWfzqHHwX368ABDjEYQW8LhrSzDd+JMNbOj3lMFe1g5dzBvYkM/YU9O8j8+R
+c0V+HceLRXLPd+0wAslFN86fj6Jg+J0rHPY2FvZHT3zrcbdUuATeA1We/x8C8SR
75TczJD+l+vo+Z2zWEgRPkaaoTBmtU8Z0BavE/73rNVlym4ChwI8dd4v+W8cJ8oH
Rnw8lbhNWFpffa0yeIIHQX8NnvOC5t62rdPLFXPHZOWfAilvGCrH6qSTw08A+WL3
Adj5f6Dp5yryQXRrec5Nbuunhm/9nuvtJDzDcRmgSoVC+5m3ZQoBcEEoAe71vorS
42GQphIBBa90b7CmeaAZcvm4IF3gw3aq2JsKqHMB3/oZAkekO2Z4fkfWXalO0J/1
zKt3sJpEbSKArq7VyQIyN1hX3UfzWkh+B3PAOA3SBX/54q8WTHN8loXv7RM0P8B+
v6P5ndcEXvldPbNNShETJh7TqlxpEnAz2CZ2BUzU+0M68beKuZHOLi2aDkaynHUY
j0MQOOJfpginds0B8WHZhc8swaiRb7IgiWQ/PNG7jbejBm3p90M2361IPeHWoz8J
9txPRKR+PNf+yA0VoUFsRx68ge9lqW0E8usWDLsfDTv2eC5K5ew7xG3UYr1SNDmX
I9hRDOSPjsPYiP+xeS3LgxQ9YybyiTn9IMlyNtYuNLLMb8fZPxYIEdjZjbCP7ZNo
T2zwcNgfN8A045qXLknnnVzefEmhHZ9UH05V8bjV3uk0Q8VNHsUhqBEJpy1PS7rk
jwnnk6ZJz8ji2uHWV9JT0HUpxjiw8lLgpNfeaJazYjo4qVowLY0xYDsqQecsjw02
Lg27qoIbBxOjHazffzx9fNzHoHY1/7Ks/WUlmTJf5NZNge7hgySzWk/jZJj5Ojn5
RsmwTJBRQFNzOLrD9vcbQzheGa3utT7Ka5WmZCgq6NQBNn5mRYGegiEo2qC8XE8f
86xCefX+wmemXfp+X/Vyu4auAwHA4qRJsahbH3FJJ4INUYOsn+vX9HtrTudzZMTj
I2qTmL/eEHNea+u0QYJObV1WLyXo16MZSH0YmGQOUG8=
`protect END_PROTECTED
