`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SZK3xXSl2X1dOfYC043J4GEWd8TsWNWpojYFxhWWQ4b8NARtrSFfe3mNa7CWE7tG
bl7gU2i6izUOP/HE6FfnjRuLhJIhFaPhTAPC5vNpvNk3vJeDPBw+jxOT3RlI6smn
qvfPB/EmmN1HlqcjsnP+eSv7zanSGzypCrnypp+1RyuWxNIz2lfAjV+hj0cE8dWC
STvoy2X2GaJ2Cy00wFXGcRCddFME50wqeQ0n4hfvOuM5935rovstPqfY6wb4BtT5
oSSJyd20zzmxUGLOoRDegWI+YNfmkJVt4PE8vlHc8s2Yn5srwcxosfdjq9uYARxY
N95fxsllTzyZNpz/CZ8aVg9/1knvSnYUq7ScbArMqRrNGGygOP6DaQiY3DCsUv/7
WqBnfRhVrx2cI6/RbQ5XQ3t1YdbVLhOoVYO4F5FlvXaD/hTjlI3p77hGByn6s68I
+by57GgF3msJ43ORuR3kV7ppEH0JQyTymZrcbR6sRgH8oxE3+F/R9EDs7K+sDFSt
WmCpVB6YCo0lu4QQMjy/8e0bFkbeNmvVde2dFUyn2JVqwalVesygUD4l3gXha58t
3bPCww1TmxRgRuDqz/pbQiDfjLSjLmbqGDo+gIdu/CoJgRJic4CvYvMP9dy4QIxz
vBned1anMS6x91qjgEQjQGvi2fY1W8ZzhmvfTYaRWVWKZaxOt5cajw3inIzwmxD2
bHBiTxPIRyYXQAaPqHphUecENVvdY/58G0RnbLN66v0/W4AJfrkb3VPg/IU9XHqI
XwVMTPCyAFh7vvll5DWE1z5DAN/VRBYOClAQ/3AGU6LLln4RME1x/98ree2ghsK1
1l554Gkby0wkfNdGFFi0MvR7XDEz/ForXdlwHOVEn07e/SUV7Dy0hy5IueRgSKNx
JdofO1smSfua23i98xxAXXgsLXdMG68Rn8j7hqM7Z4xoYKU9077B4pdGb4gYWNF6
pX8rsPqHWqe4vcaTU71XLxvTBUnzIfj/WSMcdeGaA2Ijiy7xBwL/gt7KRySeNsa/
nA7CpKfrTpdUKnMmwWiotIfmHnevDcTT5m/zYXtsYbwASpq71KMw1/lYT/YG8ad0
Iz8ujdrFmD5pAMu2e+VYFMk5I1MQuRlOBtQRtJFrvJk1yxQ54+nWoC5ndw0WSYsF
Qu8j5lwblIUiGkMyQ63ejU27/Id5UFqW1ObFFTKj8AIQ2uGNAZFtTlnLt0TgCzVy
iHfqw1OHg14vVPAlN09+K4WRzjwDJ7f3eScAJNp6H54FK5POpGe0ca7Fx+w46hQz
3SdUaBwlwtkfD4284oeBHnKXnWnxGhPtf6hoiyj+VSAiCFxtaNjw056g/sEObJxU
KY/grGv8nYOco+9ok64mcSNK3ezgqpKqJa/VH3rorrYdgS+rxbqkZUTyT5zxQxqd
aal3GM+ErCnGwFcMpEXcPW8lu6M86DzNhb/cw85KO8XaskuahUmWzq9ztmf9cMZz
Z9/yUtpYiOtw8Q6NR9HgLR7sOGbrJxDctKeWgcYBjQuVrrJrb76wFFCWk0Pd1USV
pA0LcmDBklLvTglYbldD/m81TvAuadFDk9QAjASFACY=
`protect END_PROTECTED
