`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GHnDn/P+sYuUQzp9k2WghE76EEl+Y24waNAc9T4XctRJs2o2+0nSFnkk2ZlyIaGS
kVhOSUcj+GQyJ+A3WwJWOupk7lSTL51PaILs97q26ojOWMjkmz46j/lvaKppX3U1
egHi1pt0mRf9MjcI2erowxXKDLTF6EA7KXUzgXpjcT798C7wt5lwwI0xbVw2VRA1
e7QwZQOp+gBX3ir2AhyGq1O5CZiOLJpm2ShaPoPNbxJw2qk/nHSWsDyu2XBmCEBg
56he28S56Smhh405zgGSqfllaPpQie6xRcUADSvMiw4h7XBqZFfynW/ZYhYtiRh3
ABfATmUSisghHxy7BrLmbqpPlU6H3xt0lOiQReCHRbaPyl/IAVGwQgpi68D8xw+Z
DQme2vKuSpTOAbWBLUsTKyCeTK540F7kuKeAkukVJoALUxXicazei+QU6+kEh2Uu
pCG9ptSxoDxv0dyzxupSnQDgmiboBhmGqgJk90SKlpYkmYiQfFsMg89U7S8oiCPa
C4Dcyyqd0hUAAVJGbXy5yLsaDFXAcgBbes0ura9hu5hntP0hDjQ2oDoOPVEbhDtC
/bv1ARpSWPUKh3etkLb1u1OUK3ofZEcnv2EIj6p4jG19/zPpDV8lygG4B0ifbrKm
h+QbpvQSNBN/CBymlvzrGp0RZtSpB5+u6XA002YlqfB4P1LQW6ztgKI+W2Xeqtw+
CEQOyKGmsajIcgQoWdm4HZpQlGW8QmipTLtAAnryRTenUHHJghT5JUmYRvJJ7nNZ
A4Q7dI2F7aGXCKQ1pZjctw==
`protect END_PROTECTED
