`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3fARQ+cq6KHIMCbsQUSIUy9V5q34NV4oda3kkzw+VuksC86ZNbbGkAHKqvFZHMhw
7MpWTpmcUTKV9W3PHcVGnonE9/u7kcECjTTG9d+HCwZWEw5cTkicer69/fk1YIwN
hKxmtUxyDQ3fC9+mB9mIQMPH1YzsGuFdWqLfEH4XaC+s1YHRRhKiH9IqRwaCl+zI
h7vxXBW/h+nDxieoICeLPhj6s04WXXeDpbOPBUwOyUe8Qit0ABQtcWyVvGwlEe97
5ByhsHXH/C/LHKCze16gJfzr6YNbeXBWw+yV1bfcVjatpJX5SXngGWhD1XXwBbcN
zzLomKJ9pGDwaITlHtJX+GGCHw45IyyffKZ0Csses+e0wGwC16mKVVlFk1Pe+x9t
JG2uCR623vuEDYtAknRNpUQX3A87mJ05RpDSHxUbCvQ6O+g18ZUBTSsRiidkkm0t
46Tcjh/BIahPhtKctL2qDMemUOcwtTJPc3eJSwg4Jf2kAlVSq33spVpD+BIpL2Rv
I8VC/2ExmFt5TN1SQdlQR3owdYgrit70QpSpIyvRzk2LVD35VcnXUdBp8O48Iyve
oIkAl6X1e8sEWAiI833qlT6P14u2KXYlj2QCUR0IGfxzmiSJfdSR5DSiOHFX0FnN
YLJK2KhjpbGgp9HehdINJ8aStgIcy2WbqGDOSo4dWcOSDamZw5nSGHj3Y/jpSS6x
bvlcR3koDZI0BnAd3tt38/aYW5DasUaus1+YbbD5yE30BERmIWlt+1QwLvVgnGst
XG37jCtpfFfBsy4l6tD+R28VfCh8QZpOW5RCGRIPRUFoIPrrQdMV2qvg4a8kyI8A
FNahZfbpJER3yS/FPJalQJpv48XTHya8n9IVPra86vTyXjcm0cC61hK3bHE2BsWq
Igrkk7uJtWteX5LKocrhpTJ4WkTJNL6+iDnA+QZDstPMQ4emtLq85+ZewCfKsWNP
`protect END_PROTECTED
