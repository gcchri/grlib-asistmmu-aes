`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k3WctRPw4QCcP353qvG62OWbBaM9r8NRlLneCFEUNEmVp0D6ZniJLI+GtFE/BuP6
Etn++2TzAeMfgJGII6R3dVfYtx+ol4ACMBy8PDir7P0agGvmRmzGaWxljDR6Ma/A
bVnUGyJgSqDQUglfzN+PKe/oRwuh4aaQ1GcQ0p1TPrBg/UeFiNOu4y7RFUsJ3o7W
AD3qe5EhnPqld3i6AI5prvzoftgCI2ZEnXfEai4yP2/9QdipPFTiN7y4Px04mxKp
fh7WVxrIfEl/7zkI1rXczQaMrDaAC4GborBEM/4L6zLYHIEEWHEw979DAgHktD6J
0UVYt1sjuFU4fkY52cfo2Dwh8qNHrwRV78R7L3xCFnOM7YdouABOvaESDJFr/vzg
dVfTH9WZqPA3nHUAUycGtRCTbKebUb0sbwc+hIZsUKGNz4SYJqPcsHEW5d1nYQ2m
9nav7D6CsLvDWnFwHwbt7VDZvTq897CL7282IHBXyK8+E/DNMHXY4Bh0MU8eNTLB
CWsgJJNR8e7Nn4kGiXQMQBF7+jsjcbo+IW4soZ4UXfMAVTcWxww2E68jYQCyuRbs
WfwGaO03o8lSydq3sNP8/T1EYmPg864X7Pi6LQzCeWkPvlAwC9gcnJ8avH1cyLc9
Fb91Lg8gFbzb2qktemZevNkNaIaYOfsFnZOnCWIuYPDmwhpPkUuWjvxvrFJ8ZvtY
U9+aJIUzSirH/BXCi4AbsJ6sYwIcSAhw0UxVGwasrtMFZxbLKVjQyYUjQK4oPRjg
2ntmFqCsvY4lRAtJZMGasjuaHS8ziMge+fRyeFrB6ppdErM5w0/YJ6QCVi8p0YZx
Qasl+KacmQXT7skRoM27j0ZB6tbKc/y6PsFhObpBuzldkyJxjvwJ+C5XuY5dt0/y
7PmJe5f04JD9th+reSp2Sw==
`protect END_PROTECTED
