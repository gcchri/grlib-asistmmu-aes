`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PbF3HmkIYV4lqr5lNai2Ubh1v0iGfo5+yiTa4U9ZeVZH6EKhjo4x2sntyZXQRSBJ
IbIgZvI4BBATkSbKX/ZquM5zwroBmACOdXNPQfOgoLpSYnQE245wtm8JhtH/rNwx
TlVdXZFL6im4B9TAM02xXE9TjVmR5+rFblXzHufXFIlIrfQp8x0IXRxAJEM4AQq7
LEKH1AtnsdeiMX1FueVisshdSQpm+W3775WFJYRXf60TF1yz5vLZeJZazPd93EwR
+apnjEQSyvmJOQ3LXt7RjmZTY0RmC5nIRGgSPZCrXlEh1DR14ZpGoZPcYV5/RsUV
hU4LjdkCr2y6KTu8wgzHZxG51faTePVaTeYkUwnF9s8x1xxrkPK7VotNT1eEcovx
+7TiED1OOnoaaotrwamZQJjw7UrCh+jP3PFRPjwVFGL2rqQqePXTDVEl9Bn8K3To
`protect END_PROTECTED
