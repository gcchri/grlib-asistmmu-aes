`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OaIDdlD86tNFovn6gafdOcTuHvjQbOf3DHdVWhDdMqTW6er0OWNERIvsaLOEvS96
PsPY90LbMwh8tPUDKtAg7wScjOpgKR2SadVmhb+Uwm5kPKBLec+WDmm92mUohNew
apoku31Ormj3jAIQs9UnarXggcc+vXYC90+9DBKUC2I+LUETXGkEjUH43R73LyHn
UfGdsxuuDB+Z/L8a1loez2iEUR4Tyrmo93Ne/SxDbAXnAYoGXvZIXStx/lIZYoKC
CcBMj4o8xWIwSAbL+tUeV5s5qygsUuBnqjCEJwIhMcv8NjQHqKMa85wHu9E1n1RU
ZWVPKAwiqynTvFnK3n5620pLBsEORtZTTirJsMmqn3bHQGOLSBelBxmN2ksS/UTA
IkMtaMgKkw5eUpZxLEFkTjsKYTnv1MLyaTn4wzxD8mrOaPf1IJa6uUZaFEck0zq+
ONPdRbT7OubiIz6rUiTF4ZyjoRwo1rPX0tLo/Pa32/izAhngUTMHCe03gAV6qtH+
OXcjSX2sx2Rs/jQ5Vc1nOW938n0i1v4EKdn8khCEijvYJFMlOvw9UmUR0IiR4XIP
+eTnQMTrECSWSYhSfQNQJD+V8rivOWzF3YoUGM2ssgHSTSKSDRoBqWCuhvFIg5f+
z5OZDekvbWwLEMYVsHocpgz+o2xc4y7PVlf9ZwXztzSdP2MdM3VZJU4TEToSisCC
kArzvlv74I+fNumoNpOdo4G5h1Y96FrQ6cEwncnovSPTpH92T/qaUvBoFJEwH+qi
LqAyvPvJQwC2h4UWmU4eqJFukxbidE3mR4fKayBZ10SrhgIrVKzcpa9cvoxRPFlt
7ZD1gA8IO9+wLBoZjmAc0/p9OjtisNR7brcwc3Q9Y96O6iBme6Yt44gSacmBhS97
2vDRvljFHTPcsk9ujbkGYJ7yvOhYX0ryqoUj37ojxBanzTy5d+ztnRHM/CJtyaF6
pUDA1ztB5l6xNPCB2wn1aNw8NdLX2f8BajJs3ZD1e3Or4a3oOhnv3kaQ2TxzhTkD
1P5ViZqrcAT6lrhEOe7ykvu//doc8vLnti2YG7D4Hw8/VSffC5DK2wIVlxFNZUUB
DceK2yh1mMD8BDvYp/o4L/rOMAMXhjHZjX28wcaY+DoALK6YVLDo8H7GjzF1N4O+
SCd2sY19idhDEz6S4uUPcSo9i4+5/R3Ar2zOWmN/2h8zQhUaRoXSE1hUA0NUPbG4
JZYPh6WhOZ39KXw+oM/XyXsFKV7E7cz/cyvd7yL+Cx7OX3z6r0Ka7CPcGDrOKwil
X6WPx8jlZGUl1V8B3zPN+7s3EWPbCxTc5bXi/MMUMtObPZ/DDaPA1iQTpzUpGWW7
E2R2hxN72144jUh17/rk/ttndzLaI/hYL5o7KBkFKwsqqOw2OMnkruLouNMoSK3v
xIZSageveQuouLXSdganZ7j7QDs4J5MB7IaWpCVVnj8zr8ShoL50uxvdjvC+kkz6
vR8P5i2wLMwCzNc9UckSjpttdwHSuSdvM5I+T7RNhhwbqYofHOj1kHBAtvdnf1js
JbmNCnUROC8UFstwZyN8re9e0jW+HteYTyVJ+2XnJ8BARX2/FqM9ocLexFhB9hP7
UMzMlEFhBzEnLtTv9E1e0wqYpGepZ4XQbLl7dMxxZMI3z9umh3mRuRuFXAof53TI
P6Ib+vjZerj4UksHZ17on/qxXfEwmH3cMQ/dkbqZ5umxyDp2CqBQXnWMtLfPVktb
BSi8r82JFCCnp6QTvsOEguaNei2vkrsPe8t776cbByNJob6Uy4uqeJFV2ViFlOqb
VajKjC4Qcs13YgduNj0wNxbS+38FTtvhle+VOpFZiI6ilR3pBLecmOSZXJXun76X
wy9/qwf5ELxY26SQyF+laiD8AhTIcAR8l7xdAb3hDLRQ5T1rdYX/YGujKsSvOjwB
W9XGfwOX2+VNDBxU5gVDVOiJYMYkoT/8UIHndm+Hets=
`protect END_PROTECTED
