`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ez0v08CQ5swPyPybsDi2UrlyedTQq/w+4OKtf7hVWrfL57dWkBLXZCD1BrjQHSqe
2ginlu97IfMi4eoxBlAec6CUTRXe96D3NkrQYk6ECzaSOloThI33PkKOuFd6z4yR
Vi8tLnxrgEP8NJUDzNYk89gVUN8Ql0RTSR/wNkB8/UIzDfb2rywetImwuY7VnHD/
DICEL+73y4qGcfLEn2d9VZpsZH1+TQaOSCARtfcbmvmF6RyZeHfg00LxmfKWadqT
xJ5+3jIuHsENlG8LS0d22UT8dSsek9x4ZzEI2ce2X9G/SB77DeMZjBjT85SagoaS
tdEnu9sT3UFGyGSB7dPEbEKpDTjYyUwP+yvCa7U2XDPHdP34pwKWWG+SLr2u23Kx
wSvEKBNF1uoTI3hDiSQCFv6xyV0/TXDIeglFUxXbLnjIZxdzfomy5bE33aSVx5eq
+VrI0G4lzrAspUSforf1nMJynonPSOoctfd54xr2PXZQ8WaVcfSINusDsqIofeid
2eFvjQfv7AzlYae9+UfCiwld4Yx73pHnhxs7oy56zKrv59/ZtTJIk01u6iSIEQBq
GlKFKlvaKc1BTiw936xke+G7cVcBSMdOJZlmf6zMj5V6rTsIZXsBdHKG6Y6rb5Vh
x0vhc657d36jR1PH8gPXc6U+U9V9qiqcFXZnWZXqA2kRXtUxoefYiPQ6s0t6+tNd
0Um3oZVkaeMNgcp8uxneSg==
`protect END_PROTECTED
