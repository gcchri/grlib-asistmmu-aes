`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vdh8BglZbbODOC1FzVQOdTtBVHj30+F3wnU50g2/9c0ed5Quo0o2C8IH7xOnvGWs
Oc4O/p4I67rMGBmYzyfiK+aLrnP+wBeFmVsF/MkNrMEYD+cBysNiiBi6yurcN60G
wo5FEOuR4sPypmyLXEj0AG6vCacmFO+5mIH0Lxj7uWPRJV43unYnKkdedCUeMPF0
NArPGkf6B20tk4lViO765knjIZ4bc62gO1TzMZziCiJCMjnhnLbcGgGFIKBtJIo+
m2Jj3pjQJ9yqS9wRNjcAzr2e6FU/sWtKl9GZ2xoga+VawNyrzY0Q3QCiltPikMZ6
eK3M18mpcvEJjfg/Ktex39UNyzCf9lKy4GL7iruHzSN4BBy2fImYGBMuxc7o/ZgS
xqBQwarGeDj+4o2u7c81SXjUpezuXy+SkloG8NAvNuZ05o0/+zjvNI8DU4kjHvHz
u7sHESZVdfw5Xrav+du0pOu4BStjCXDOJIM8fH8OkFq1p/vg5PSNxzU5zIUQp+A2
8HlNqrOf5e6LwmnwFqSs2U2CzehhS72AHEs2d9jlwSzjN3usf0xGYgUXyHPBWwf9
TfFKSEoqNfFz9eR5Pekq236XyG/hl/p/ZzCSwznM/PTu4jMBHBJHYzhi19Ns6RJ/
KNUKZ368NODBclCy4yU3XqfaPCF5JocDe/hJPeZFraSVo1iqklonaPQTn7iMf6Yp
CehQV+V6YpyUJr8OCwvMpB43smk2qqhjskOmZw24LIBwJTNomy3TL+43hOvVWjUC
IvZzUJsGJ3BY5DAOzNEdhIWGgAypo/8uQiMoiP5FIFolWbJMoI2RSCctshNIO4id
JK2VcOy7VnhFsw0KZI0Qf8B/h1mRQOonCuihG7/Xr+xgX+u7fYuYeAovU2aBQ4gz
vX7Ir3fnS++TPCZ9yYxbRs5uelw4RgOlN4WRdwbnZbQ=
`protect END_PROTECTED
