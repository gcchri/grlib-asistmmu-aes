`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xXbX/FCloF/xD5+dr9yj+XEvEeZH6NVD4KucT/FlgKQAi6cWNVcOxY0CunVGY5Kq
CKBx72pc44GhRa1pI2cS6UsU3YlsE01h+9ArCWVjA9ufri0a1z7CWHyJtBQI52xA
96C20AdZox8iAOV8Sp1EYJUTm64OcEvyhirjXYfTP6aYTsDUxp7JoirLIXreIet0
H5cT+gLyOqaH3PBK+c1F9IhI3mctZUbkqCtPXXWI3BsT7GfEaewh9ItSZ7JBbyI+
nMrn/XuMauipuVuD3ec8oW5TVZtxepseQA0qplCuqEuH4tiyB86KqgWPK4tpLWxz
hAvRR1GCpGBdaF0hS5JW1r+HUGzSvuT65hMKXMkh6LczoTJd1fN/zmydx+VyKmet
F2IbFN+xoVUO7W0u3pie4lh7aetgSZyK0/Nkv+nUOgZP8e1J0GrN2aAe0ekUrGwk
1KLwWwS4V2effoUFTQSvArCNSJ+ODJwkJ9crdZEsHVD1R6dp2IDjmqEvfXYrtAvW
lhpDLclaJ20MaDsUuS7d/FkmODa4mfjcoWnajbXMHk8DL0oWAnAUYkMqzVmD2QLT
m2kWzl/eMKkYA76LNXp4RLgaAc9nD17N5rqp3HLidPGeCPNukpYLWtgpiBjJxELF
YY2btwdvy2LsaiIpPD9TUOkwzg1Lzj/x6myDU+TqolARuuzB50Z2J3RxDj2f5vgU
SnQBmzmarwiu7PA0exdo23l9QHjOKD8SFxLEIBW4c6/tbOZjzhrtQHYrS2lC303m
zLI0MN5jFpfH1H2DGLwqmqNB4Uzg0Z8IiB5f1sE30yJiVj36iTK8eWLeSzpwdnnu
usgGh71Ei9U4rzWIr/Ugcw==
`protect END_PROTECTED
