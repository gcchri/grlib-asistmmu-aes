`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pkcz0Oz3j2RxZ2WTgCB8SzIOBYAYHD2Fs/OWKZRWljjuI+itxWFET7hMu0396ZP5
GcbvlEDV0Ye3lmCNcknGNhOD6NDFnLriB6XoRHh/Fummxo3JA0Ol/h+nL2LCHqz5
MXQQ560oSfThAEs8Xk1obqxn+MwJG5ZQ635u+OiOZlRUoc6jVWRAx6ZuU2sJoIye
JFc7snZd4ZN/axeXMuntzxysi3daM9YNpsrJKgQypnJYWh9+Mw745xIixtWECu/y
AG6WCLJre+VWLFtwN3UxWC9YUfamNpxQyR8ZOxw/AFqiX3bglG+ODM1Y7toTfm/B
jXeSrwPzZw6fstEw+i0UD/DGnxK9btnvOIqfThsxuqyWTXMlRyk6mHtcPgg0rpJa
GAZyuFL6aR8XsO3FaSb71BE/8ZflSmp46/M+fwo5J/05RR5y5MCvl4+ppn0a9B8f
IgwtG+YwL97DZ+BHZzfb+1zlxM9Eeo3nbMTxOTJ5Vx8265fHWD00eomLB7SUjpiv
CCDYOzSTILLSvm7hXbPUDViNqmm+Rb/xFRjM/TZiPJSnGOZ7DR3M3PKdq1BqUlbx
ejKK/zhHeT4Z1/GcORFlxYz/5/0T9QRuSp/IYQQcd8UTQG9rH2h8SVKEJ+Bl69fK
xdv9lrPLxK0SDXNEeonT5DflAzdNGUCWkWxB2acG+OZQkucdsOwn0ayoZ0a/jKS6
BJiQNJK6F4pDPy2//uP+1evmxDN2JAFPtrywLUNw8uixJd+yqagOIJc/K5r3LVYW
YJEkis45mK/vEZpo9gbpWlEZjABe85xjdxvDad02Uu2Y4r0rO8YG29T0BdskLzYU
azHchwk8ISKQ1V8NVcSQuEXOV5k+SabU1ZSozAJE4OVBdOdt7AG19MofDKR0WGHC
BozaogtAm9F7Uf1FfA8pAEvOUTtXw6oV0hoEapSQEWqa5KtJbZaNbo+0gcBc2iMP
V5frDypxYLveLF+VdTmfDPzYo2w8nw/iCRfoskt70OPxBacqmpnGuQ4Bs+jCt9zJ
2ZyeMDVflp+yFt9Z2Kh9Q7mt1/IIOJKHcRXjNi3r32xxVDm3Dl8P9tJ/27haVMVI
8Cafk/E0bJOhWZJG+twR+g05sY/OlzOU1enSGDP1LpS/cbOSrgq4Cu1Bq+Vw3lwm
XwHowaE/zPutO9haY+pCUzu8Ak6xWmK4Zu17fDxlLYqf+o7kalcx6Zl1UhGzHf0m
Seo/+AU1EJeJEP7Sb6NdfPdOqEhn+eM76KO3slfzxoQKvuyrr+SFHlJfT8usZsKR
TSJV/VkWqhMhsQJGvoO7lB2tDZ1PEaoTQqK7EJfILTPQ++UmcIBl5udV6Zk0ikNN
Rj6tUuyXollDyEJNPkW2sDSKwhLPjRE9OGu/t0y34IEaJH1lUDMgya6N2jjCXtCG
0N0eeyb13ABPONXaAa9qWb7QFRBx7Sv6OTIQXsG2Q3yga3w+BPHxA1bN8EkywvOQ
nREnL6osgecEWzZtqC7rPAfzhRcMxGb+7MLE6RHGj1EHuaTdkxWfGRSSbUVu7BXj
24SfZj7rVibPyF8EwP7EKEVELb7L0SJF+yEXEcv8xLsC0ydRAw+SiiXbn/dp7CzH
HXrBtwXVZobqb/+jOV2KCFi3GLfx7DWts+G2jRA9v+Wysuk6WmYJ4KjsP/klWfLR
XfwkfkqvOZ04xLpLeFHhY/dZQ/BQjwSR9kSyrgZEn0DkeoB6ZkGd7zuIfCW5mHFJ
c6CJrhTOeIN02xuV95l1oXCDWoOvuOs0e05AqjILgU7bVZobwXHEs2B1ksF0C7/m
Khqa49yNNisZA7WtDEh4giOlbweaSlnw4eVVzyfuZMBW+7SeDJNzZRYK7yAeW5x4
iA9rRvRsyH4a9UUgoOTDjH+6lf/SlXwZ4E3UgC/r61YR9W1KnsiZ3ltcDjlZeoZQ
fe2grVymJnnCsXh/Oc6JpjZBSo0OMyFakRMJzYMIQL1Qz7das1MNc84TGJykMcKV
4TlYB9kZ3wZLN+IJD2CdMA+XdSti/aYNC1JNl67KDU0yJjb6a1DE3wVZVSl64Gfw
mWj4bAq+u8YynlkuERsWM7UlRKBP6Aw1VLHt34n7Al5/zoUkprAAb1FiUS5sXnYg
vitv57YUCOf7tFNhEKvNvs18MyWcg7DJhfgMI6Am/ra8K5On/T5y9Kafo2ey4STz
ssxu/w0ZUz0d8E4+8VeLmpA8nLO14FDR1foXcWqX5N/nBv6xd8VfpHW88Ryf11K2
WxRqk8pXyzr3Ir33H2Up2EOo4tYcSAlf4LuFZCa6SMQoNoZcqUnHjqtHgQCT6RLE
ZqX1lKdrOxpPreE6OR0rp3v8BlgtxnecNcWayxsIA8/0LWhFbVy1mCo9adnmoK8I
iosnwmdIA99stDdwuU/EzPUBqt//NGILfijIF/d+owlFxjEz3PP3LUQYSjPHq+dK
+rS88B/7EbEs4a0DyYWFTbFBY9FQYaGBkv9sjaTBtYIX3YRBy4rVgQwMH5jxCwB/
BJNflfvjJMXiWpNah7uYZua7MuQhYTFuKfSptiJLC9I3vTrzc/ZlZjxuy0q0M8Ha
JuuDTXZLyu7nUn7f0tgvhwGUJeBxVx3wRjOklBIoKSCLjNk6cPCKMyBl9mTzIwEp
COs9BIRLM9N+FoVB1kAgsFxWEWh0nFgjUzaY16+YUVr09eAPO41V3jpuFGnOn6iI
utKU4yj+Ty6lRwbXW50a/dMWUVPfEUS37nyJv27Kc213QdS9tJvk3pdK8TJLRILu
qRSUyIwILlQfpFlNP0nXFkYcXiOLVzMTc+UBqtV1OaV8pklvioXd7aVuUsufRQIU
8OuukSNa9/wwlVT7sGw91EjpplFD/QcOla7wcJB9DfGE+5D8sI7XbVLXA8aHSfwB
SVCa4pkgHSuzZ85HDy75EVjyirb+X70h72FdUB809WE+COjzwuDtii8FrgxUtegj
1QcX0N8blR3piEBB3WX/5IAuIiOxc4wDorth+9BQVkCARYYVsDWEW+V4ezxWgFzN
2KaUvP0s7DI2rQxRkfnKmEz9ZD5mTgLeXLOC/Zz/88rA7NFqeJUMappTR3B0aKGV
Z20VxZSF27N0WSLMFSf16SJjz5C//QB5OIzjZyxttdIK9SMBg47qDt3d4FpQ5g7l
bRJ3tat3aqryNCG5lwbhL8jAbEpGMky5H/dxxEd/ZTNriXSu8l2uWMJkV8JdOR8+
jtA/v8zVFSmGG/Jhz7kFAtLsIsB8L8DVzIrzsUKSVrryc7b0NY7cCz4YrEoIpcZo
EtU6BfETluA200g1J3Syc0s/KEJzFWYbQT28KLuRDeDw6J7/fFrhKDVD5Y2UmRhE
ejfjFAH396GNhkS4nMks+TCd0BwDodZph2lYzIhXq7rz3PnM2DV05t6hcBIpi9Q6
8MtWzmWCzgQPVnUmz/KuqH3/JyoC3sCWkKma5wkgRIw8ohRf56YFEyQQaJp5KIDG
L085G8wiQg5aibuemgmaf2z2WPy2eppSWRZiGxB4eEBcudzzBKkUloRxXqp98mi9
cGw7XUjIiISgYNQ2/oxNfSRYF+PnLSs2nyl/6N076utS/3SMfzy2RwiXNzWI+xqt
mxhOYwqCKNOUuqixYgO++L7a0akte6lp36buXKdhjx6I9DxDKoCxrVP/2wqDwUh1
h6If9mQkT0NuV2sWlYJuerLU6OYQLbSJX7NReLX9u8dWDPU0ciOr9FWwE20Rs1lD
ZQU3eaBE6/RkukryPGurPdx5uhdHgE41h6cikYQHjtdX3UF38cQN7sFfoPAChAz8
9vGlJ1iGtS7+U37r3m82G1Z4doQtSf13yV0TGg+9rU9m4+xB04zJ8lGWjQpmSgA1
Vnd38ll745nGNJkr1aq/6xzajbKSdUF8xJqQa2WV1wPwLPzGOPMzrPEIhcK+KNbr
mw+6hDRgNzgCv8FEjLyOCgl84/Bv2uaDEsHvNYiFb/Xoh+WItuSM+tH/qmJwmEt4
bjxkdtsXyvIAq2lJF0rVbu7EvvCRK+x6IRY9mFH24cFnPi5sOW3sE2g4kPAdSDXU
UueBtiW97wuRJNkpIic/AV7luiQzeknTpELomF2JElGjKP7YnfNifyQLktO9H/Vr
koLk2UKfZooALjSdkzRu5XFeTCGfaQSV/RDgK2ltXoHfJP5hhuSZYhKVsJX3PXtz
gkcq6EPAnOl6/zFqLLTQVH3uZM4GchSRGbBVnSpBNx8XLXMSvVnGqeOiVLvHP4qF
D7j60TDSnPhsfgxtVgyrmY8UN14CBoJST7IRQzr60NB2jDx2eLkeiJGiOm+4vnzu
8pgZCsDtPsLRLRcfy1PlGg==
`protect END_PROTECTED
