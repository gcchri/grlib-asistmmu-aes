`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YlwGLFFQwnf1q85JEZL86/dOtFKJlDEGOjuXUVj53SnG37z3/b/c95uv4dGdDnxo
rvkjwlz/xU4ZgQoXvUXB6oiuy1X9jJYhF0qbCFlBbKEcm+7GUrToHy/qdW7QrIhl
vDIrQwUOjaLllfOe++GuPP6KH4tK2UmHIJTFeDwf5L7xGiNwhdEzYHOt8LUaYnZX
D7r39ViLN3HdQ5j4utoWc7FxEWKZNz9QehawUSTkaVZ6mPW7w9I2eTUJ3qoMtpUD
bx6eA2LtVYRB5jRAwiM882zTkbDhQqcBnCbwRV3fCUvmMaphESbP0hHyEEZZeMFs
FqJ1mGKF8Q5+seJuZ/4UPsB7vzCpipE95S29K0OYgQUGkRFCP7y4be0XDaFTduYL
kucS+Jf79PsSDwrHZIXI4+DtfWAO3eZPb9j7+po3kmesCkEAZXyLZAU+mU8ti6JG
kEodH2I+cw2GBrIwV4aZIw6XaTjmPPO5Q7Jn3ngnqIbyebTnnmXlIyluqz9/+7as
fqlMhzRLZTSg5sacvtcDS96ykrNLVRMdPWSrSfBeod0FEsYMlrwQo8ozz4bB3AFy
tDnjNEJK8PKEqrDt7E5Nl2U3YNt1xz7cAsJhHW1DUiNyfvwqko/HWPMKMduu8A1O
HVPhmbWOxbkxK9p41NMgjqBjAqqpsyHuowqoQLz5qmQf2KWbmtoqA4YnjNgNvk0S
sc7TKFKf1NHAX2nLvPZ43PxSsCd1LbkGkub7FesW9Y/zGTxNNmsLS/G2lCxIuC/x
550ewcYYEMqKOUwyPTWs1POafWGEzGzOziWfwO3fBzjNLRksN234r79DPRHO5AbO
TXkE+/jvu2vEc8CvpA8gaQ==
`protect END_PROTECTED
