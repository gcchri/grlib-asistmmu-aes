`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yTf+CIUlGPenk7UvWpSCTNE8KJ+mBSYPaA8qXytntmoaf5NmPLbTXMtXKufxIGfr
Uvrs0qVLgmsASxiv/joObbyp1yPZsrp0DJf0Ol6rYsGV+KJjTAHot15Btmokrth6
x36B6v66VXGYO9weJx0FHWs4NwXU78wbw05Zov/MmGdK+pgM1RbtCVOlGmhFG925
IuX5juhR/6UWnljnD3fuSJK9VAT77NFZwxMF83A8zYWb4DsiToBmbg7VVnQnS45t
hormlUnBpo3N209IeB+nrP6VHKb7arQ/r/PwOLbJAM0a27FC56pEJjLRSSxWz5r0
0Si7Wggs803lS0iJoAA/g9gv//1lL+7l46hUUcmy3k3AzLPd/5Y+rsEQjJmVdheg
gSn3WIdAHdHykQqFGYgOnNkZ6ufwdLhmZKjEHQk8F7CZfyby7UjjSLxQUfY/Bmp/
Tk3CL3OjbAKPavcwhFPQVHRVkETHoWN3Hh+XnW5hW1qq8GF/UNvHOttV0zDGB1Cv
lsnfjBQ3d874B/RVQyeZYNwK4WjN1hpeV0xEWbkdp0yDwWU9fyuyFml1s4FSx3UG
DbZjOoNsJct9Mrhe5p2JDv69liNX2mEZPCLm0b+xfXWuuFDXlYxwPJtd3SNpQ8Ty
6DsSB8hMO4bQv6MmtdSHgJ6crmrRnqX4J6wA5ORxeWviC7cRwxdW3Rx8euEaqE5T
t5RQMfLoMICIldGPqOrhueNkWXDhAsWgXfs8Su3+xMFMUNlOAtWAlyI4levdQDO7
VTG3XSy32db6aBBPtACLZ3YadF99ZlDqegyv9LjJi76GlRnwd2uydhb9Sz+TJKTS
R6AcuwZv6PNXA/CSSa0oRvHy27rpu2TBFubVqS7TuKXYtCt8NDKCM01nIKbiK4fq
tiJ8Mz0A8vsaov9tnRIfYH0RMlyC7y8SDbEmsTC3eEGT8zU0Y3Vopr/7qHmbW+QD
a0sbg2jPgOC9gxw82hrajHg4eK/q+WNGPF6DjfOjOU4dpNWAfTncdAobbgAkQaM7
j1v3+4FzBk1GDIttV4WjseHYCfA8YzvY3RVjzQaUJ2lXDykSYXs/cyyWGBsK1VPC
1qq2iUcykoANHEpkK+zl2b3BotXhLLWB8MM5zMUwoCq9lZiPqgLKDKmPl0TOVh4m
09fwQHZhZUjz5AXokrz6fjHzdgTZBaliUJcjlnqto1Wwk5GKPLPFy21fzX2XpAH8
6Z1p1oQGMdBfXBJxKL2KkUDF8GFqsSUI+q0OhsN3d9eQ0P+ktAVOWw5Im7yb7h/b
hOng0gIFZ6OCZSmdIfaKlsDemEtIEbThzNr68IaDDm/73ntcjRnvzjKSIEKBEbJc
770ialApzc+10HIZ5Lpns6+42Px+V95ZLSnmCMFjtAMYWYcAvNWiLvv5hxh2apNE
BiV2P28882TZY+gy9nsk3ZxHCFtcFJQgqG0tA/jXvNf8ne6sIVlMCj39QwrQq93J
ZtGcNRf4psjj3ILcYgNRUh2szAzFXSI3UU68a7la23+JO2TMhL8bDpciHJg0hech
D7hfvTwBszSaIM5iJElEEmDBqNryPhNcI2gnKAYiHzdm6nmP0mzu1UV2rl3TfbR+
DDtG4mtOMnU7zQryluYtNfdP8MuRODCBQqfpF87L/YArnY/AqwsQpL6lJun++hVQ
r0+ES4QTgQ5tKPtX05BGp2l1rhe7VMGlt1+hmnW/KrLhzq5OYfuWUeaW3IVGAEsM
86W+4mEn/TSqw212D4CeZ7c36PIrawXopneR3gqqkLIKttZbaCpq6hE9ZAIs+m82
xP4QUElvaref0a6PNmO+OUM3neyus7OzgB/wGylzn5wSeRh3iy5KVfn5il4YT1uN
Lt3wNzITShyYiNjchWcTBQuJbIYlBt0mi3CjuPrrIU1ZWZ8UTkh3R5PkEkrRiO2E
AhYbVv4fwmRSJTWiGTDvdjFk/xER4zhemtfP7sd20xXmiYtMdSeCdJClWroe9Uq2
8snQkxfuGSEh3B2+NnRClzC85PYZ+e9JQdMQawZwdNynmyDAH8Ng804py64mGa0o
YaDyjEsrWd8VPHsFeb9WJV2Vc+gZnsKCYx6b8KL/NQ0=
`protect END_PROTECTED
