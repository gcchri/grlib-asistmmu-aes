`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dryiNFYFT3ILm1oCb+sGGFFVwafVHF+SvuUKz2+x7enOIezMddvm9EaMG9K2O9G5
hdTQdAfVMlRndc9qTFFnl+qeVGzDrHPgGmMfqcvtgDQINSp72kyHfhpSPJY+ldEF
OY9tOAGjKQTyAU1S2U9SHETgvI82d+vA4nnliNGBtTXC2zOhx3g0TfmOIfkPPNXp
7lJWR6emYN1okFBTIr4HoY0GgLb6svoAcAE0UiF7ZBNnCQPFuXD+Bbdp/2qB+3r3
3ZHiva2CPKBGOA8MRB3QqmILq2Qnt7nYPSq1za8/1I41/KjPRs7xE4Ism23bcGHv
21BUEDpbtWYVX6njaQgnH0HvGnTebTsV2WOE6u0xicBXD6DG7C8gIIAJZ6Ew7SuM
`protect END_PROTECTED
