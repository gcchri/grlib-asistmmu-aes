`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kGqz9BBdR3H9DQQY7P0mHH6w6hRoei+B5PymHceqppR4iwqUf5iDwIskYWGw4cpW
3B7Wd2DMk+uj8tP7oCCIcEiPVXNbyx7U60vEVrDB4D0kYrcWbEGEAJWiSTwi+MWv
sx5krexPu/ILS8ATJxxzuhBGwnAG1A1qmZv8k6TkeFsl5JZH8RX6IPvYRY9aVYDo
E2wz0Z0f4ak9WnxzEnPII6XwiADkpoUw+xtOkHZV1FPslgo7G0X5gPN41VHdNnLV
VTvTjN4MtmbwH3yE/kcnHiYT3dbC5MKPj49l5JlarLN8RoUVz8Mk0NtGSeSxfOPf
lQp7o6+VEuGRBN57phhQu1LlOe+PSsmJmHb0KuL1SeQmtDGuiplThA7D3VY1Z/9g
Nc5MSco5U2ZgtjUqmxN+AH0tV1iRhy8T9eDBnw3Le0J/W8aKDwBqTJS455uxB4El
fbGry9akOc0wZstXKobnPkOl5cWYvmQT0FD6s6STXgO/VDX1bSAj4n64u13r9buQ
lTQ8409XEfIe/KWXe4HTm1GH4FtqRJ/oqOKE170bRDORm/3rH1LO5ZpTtsRAqIuy
HiEM7uXGAr0HrqtRWlf/kqm+4fjO5mdFVMyd1LIBSGTXPue7frac4bvilBLKEDrT
GkTv6eBKm76LuN8Ih+ZEMwkYqL0w9VFHbhCauiNoelQD7pbXPbfdbnHkNz592pj3
GP/xShrqmFKBjZpHV7htFyn5qhCEoex7azHdhvPBmFQvRgjzYwqszOXjR2lNcjCE
6mdf35izKw4ZHZSfSUglYjVZUKVocR+UKt6LBBSpTc69y2T+84+suou8BVIjGqIC
x4RwwuoxxNHAe5/tuejfA380F6S3uUcBIJeAfP9FChcnwGk7BvCJtpVQoOzOB2FZ
3t9jWSj3YEw4kwkaPwVIay/1swZxyGnoY4Q2hhnhkBjrQLAZv09S/tMaHq7pqvWG
ejkVNxIpVRoNpOj5QqFUxCTBC0uvxQYXe6er/rf9jwk6s+Va8blHDJZYY2A/P0K8
N34NUlwm3zXcMzaVL4NwurHRd338PsuF1ttSWIlvIxSTiHWcv40UvZnzwX5mYEi6
FaM+94crPXwVHl9iFxjDk2AnjSr9/pBUwGhXLslAvS0XC2vo7wqiIUfff0XPESdn
ZjDUA4JcjZo2B4541JvnUEQN54aexe8ijqeEl+SV3Y14FOT6wvEsc7hGLk4uHgH/
S2gUrYxFzDzXD/VwiifaFD9RB1TZuM7HhmJ9/OY5reOS2Fu/m2cfRma1W75IHnHA
gkRnn9VWhzipMlyQaokTX3gx7iPmSnxLkUAaRcRcR2Z+esBUwjp2QyntGja8lqGG
Eme9VX7ECubo1ySqr+VMGkcHTfBbp1x7OPSkRKWaAz7QxBTPzU9UIqvxP8ImnVql
kbu9ivIKpguqcWSe6KOxmR3maREobd+N8nJhkmLWv0fZkzxdlozAWFXPTGIrkNZ5
a/2XcifWHX9Pcy2xhokmhWGneEBkbAxmgo8yy3gr63BtdsTL/u5m5xkcztSrT/cY
`protect END_PROTECTED
