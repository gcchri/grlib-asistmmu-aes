`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UJ9a0D1vedE7MbAnLMtWakFro7OYJKLNSQv4X5vVwrB0zNyqazk4LbAHCN43ALxq
8ZjM7sePjBZiEXoZJgAkAXOgRblGh6UKoD0em8FLA/Dq/SrgEVprjddfKZDQ+pAr
KUtVrX/a58OdtQjbs/JNLjsCqd25/HhFMf3dcm2Ji5vjp63832a9zFfewFT22enJ
AJjU1+Ph6kaophSEMo/MZBPf/tTaGMPiVYORC6fFWLQrW/DceOHgxHj05cXUuALQ
7sSqJPVLx1dvjdowDQbIaRgQ1LLxZV3YVLsRSCnV7hPn/oWrG4iK77GIcT+XGFv7
gCdYyENGF+xTSti4n7nBk5CKJ858Tr12hjc21vCy2Eg7Rcn3g9MhWZq3t/pziBcA
PhP1USVS63sZqQQ3Fb2HBE0d/i6BRql74/Hd1U4UAk5peJNRe6eMOzzCbmJTxtzH
tg8Vzi8jDw6+n6gvHsOsG95Es6d5vzOPnuNBy3xGwFIFhjYQB2imyxyYdYg7s200
mvpZe7RSh86wztRpUPgDb5G1imbOEBvFKo1UKq8jZjNcFlAym6fUi7AW23g0Upp4
8gmXP5iRZvUtq/Ze1+KwEgMQ1E80XDLOm6F9yXoV4LTnj02C18sksLoSk3RYHwz5
1VsVBsYkBp/LssA30Ow7/y1SL5WOT4xTnqIgnT5dP/Tn6zSQhAmY1uLuH2yEw07k
D0/DRZ/8IT7oi4zcr9BlAXsKqwdFeFLPoEMxJvJcjxlESNPmnohBEeEtvetcbi+T
Q5VeqyXcw8DgKK/87n8QRA==
`protect END_PROTECTED
