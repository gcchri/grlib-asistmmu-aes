`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UrgJhlreybzLPuHnRAQbBtFnOAHympI1hv2S/qpMVb7AyAoh/1RuO6kZD9+ohtIb
1riYvmAKqtADKaIiDHNNKRlZutuZDNknJjZcl/G9Vx2H4mMZboPBofiCV0f5OBiL
GXBpbqZtiRtVl8imz5wBvReKHTl3yONLjWVf+294sZ5h6jqSVlqAuxzOpEB6Jho0
2Cm9mNMBG8BhJvaXg2UzaAVZIMYL+9V56s43bEyZ0Cq4AeFVNMdOtFA4830a+AdL
TZKhwmq5wLfDxsszbje7bHhZMXHBGC+RkvZImB1haPuMomkyAq/fPARRXkAqjkOW
MztUoaT88D8oECfppk8MDVub/mfMcghmrG/xAMH5sLVRLR2+1mttbIEEm6vJSYxK
eAu0fCJ94gtOvMNsjcknfAVEbdo3eTPdYOfZDGypsICE7EwmAIJXQ6E/hI5d/YMy
nO9u5CRtx8H10XaJ0TMIRe75cWWdnY32F+N4OyBimMTARJswKnuumV6lYAPuQnHn
XHa1HKR/J/EQP2XtUbE6N2EG0TfNs49P9Y57qCek/D4ociFOoaqdn+nlM4xhtE75
wNvLTgsRnLmULRx1Q4sdjXkNRGFQPbybkABtbbLWMRoLW5a5AI9oZIyFxvVz1o9N
NnkUtBRC4BdFTPHbf8FvIIN99eh3zy61dXYL+3GAqwBlDWJwTAU9KdkeAxCwMF1N
n+tsbPFGLIOUdFfnqKHdWk/wIrWtEmP8SO1L8OfzUKR8Fhx5IExwJU/HEUDQdYtI
r7Ry5BNZnzkgHEBuHge0YeNJcV2F8+jjEbSNN8UmRvrdfQ4KQ/vGD+l5uPSsKCi/
`protect END_PROTECTED
