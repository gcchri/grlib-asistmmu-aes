`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VR9K+0r40OkNcnIxzmPb50DZvhoHmvvuB6bFT7RhHkmaySmMPLViI9uw5sokPcwb
Fp2dDimMa8e4iSYKx9ruWUBZfY1OMaTXiAQe78+19+J0Hn8KFt+i4d73OPoPSDOG
/r4TGrMBuDR1g1lRnntwSLW2AAvl3FNKr08BDUZmUiTE5mFLpt1R1QtOV4F0GksJ
jYYbXL+ajRWxXnXfySr9qqCh1q3P8iNi/qH5kLuSYc9XyYyvQmQhEyyesJaGtADA
dB/v4cfo/ONbRaHzJG5/lM3YfvL36xqQLbuGHE10pUIAEkG+whaGSoPZ/U1ywTrF
OGjg436AcjAIhYQ9c7DXYmQ24WG1jy+yHY/5rImmZ0JOK0Jmq1agP3Yxv4aUg+/9
WyZyTSGMKsMXU+lxwZt2Jrv7N81yB8Wqu8CzbFQ1Iax+EiHDVRqtvKdsK20Dhpa/
QA+PDLUlSK65lzFJ4omeMbSewEt7TI0iCN6dbrFz/gNJ4zrhOiJtT/YUsKqJLjIL
BpSD1sTtBEh02b0rJQri66v/q0X10X29rI88Tkfd4YG6XQ6yte1nt223kDxVrBS4
2F195e0H16cFwvV3IcMl2yYM9zFWz4bZ/k2bbP/0wPQNiPhus0ph6VamNu1ga2jQ
H8HG6/jU6pXXKycOoRtpX+6c0rvgUJEYWtdPHz++KAaFEwdF8UjhxKR3FyKBmhZh
z82WZ7WF3EMwQi8qdPMEeDnwWwDlId51oqmS/Ej0h7GgTmzr5h2EDb432eXzFnrr
NWtrmDqT14Z0mJPHsQ9b83KHbzwDwfKtPA5SyG1uxGzuJyFRvC92p6kksQ83GzaO
0xy91tFg8+xnRrlnD5g2TIxdKoh6rdsf6tBoFFwJu3v0mY4RYlSmNNKQIvX6L9/q
3Pc9MLOfJxjh6xXfCmZy3x0Tl5m9kFtQjMfydLS7aZHpju+IBJS+wIRrYzun52GF
rBGxgjozsdrOL9895QiBVakXlYmo62/71rJZfhu64hwB3267fdSdwap1PCiIvAOc
RjwKgU9DE0Q9KH/q7G97fH424QfMuzMavc9i3IrtNxiamuvjsW46ZGuDiRxL48Se
AKRuhDXUCYWrHvY+991udxE5VOKCND1M5n+iM0gT+tY=
`protect END_PROTECTED
