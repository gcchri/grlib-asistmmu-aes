`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wb90DnBRM14cPB/bA0OytuL6JLuu46Ro3fiSwzRT4G2GsfICL7T1DWxaiDSAnXTg
OQhnL6Z4eMnXBCbL/B34TBXbYMccHFeRGGhG6R5fgyPGjZpNHIC7WR5e9Hn2AXuS
jstMwpMrfaWNjU2z3y9WZ0Gtu84I0aTVr0g3FMYeU9Vcs0SwnQ7tY5gixkVP18r2
He4vg2ZktYhttemmoHD1g8SW1xppZCKbC0sHjItAV7ZJFgKYa12PHXEFDKLcY1rN
+LxK0owPeYZ5NepZg2LfgfV+gZrnSiXu2guIsDohDqZ0t8zSuctmxwTbCQi3O7B1
i43XwFMBCDC/HZGxzBf8Kf8qJ7XR3rzgWn16zqJQYuq0o3uBj1S7mDyKPaMnw0Px
eeG1LL9vlLozMcyBxCCYWcVNxNKst6dt8xr5yxsp7iALP5WDniWs5vH4LJCOsqsI
mUrbeZqFNNnTr8lMLve7tIYLmPHEBznXAaLEoHS8nfE=
`protect END_PROTECTED
