`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wWZ8z2vlyn1mJWWBpOtlUftE0xhwl+EaFzNzrEeWd2PjGt7jwKNCwzDipj/RwdoW
lNxfkA2tj0lka7ojqhT6uJomMLh4OPLmQBbU/ngelcqtvnbdmiYGV2UaE6YpgclP
tbtlZbYFsESQrup9Kze18TR2xwLS3TN3afsStTQ2vs3wXYHTi1KuHoMe8nFQeSdi
5GflH91DOpHZXcOPbzKi3sSiBgt7XKNbIBz+Ojn0Oo1dyU4fFOUdmAJKu2e5JRaj
8ORVh1fCxpr3yCckNTRtkCSZ47ui5a2rdzukcJfFfzu81db3sLfdfyJjAgNK9MYd
oIVh2UOExTbZScoa4bnUNOMQw6uWwci4CzYq25WBIgWO+vCoat+BhGSaB/dIXWir
d1FY/JZuOwpYUDmj74srt+SpmdJQj8eG0OXVv6m+9DGss9coBsUS47Mr3vsbx6cl
RXstQ8Wo65qlW5OOJUv8X6bDY5/oPz2V+EPBPgckLJM2aTM1tk0v8duzo7Ysvyr6
N9Qe+PjVPg8FZPuOr6Q4yBBmGPdW4aQCp0KsrH/J2/04TzpRj6o1KcT96BTgQbRM
lUPrXgoHSiM0Jf9E2DhFX1y6S//ZNpoTKw2MTjFgkFN7iT/mOGXCCm0O1gOhC3qB
Nkzuyym3Opqbdin9zfhQG9++eHR66kI9/XaiOeajx8F3c9GSVOzeERw79DsruJFn
NMgYIfsH27XIdYKM8VWH2wab1AiCZ/AcXWJI02kQsLX48G4oth+K9jbwrjVl/KNM
mk+yJNT+ABFWeTG1dFnNnmyU4qjlFxgrIWtLdXnT9ZgyA/IiWsJxxQZkf9Xc00Zp
+iHLiPImYXkdBY4Lw8uKa3rOuTNyxChj46HB1pX3ffKFBi8Omx746gMtSsUld8e4
6EYJwjqCPvFIFtzxE8Y1kB45s9F7iazedb9u/IbfdlicyjnYhzu2VS/QdPDkNSgk
olMWZKVYVXSYuuuWubw2tYRFahgjV/4OUNdKGXaGFDlKCMCOKBHX7BEcSo9Pcozy
mWd9q+95jvLQhOiCIWXDjixV7BlAihszUmQ5TMiUvrMSgaY8MPsSlPFtr5gmLxgC
JEHMQVpwjUhkgjyGB1eulOksIMdn6vg6QD5RqVHBIULXrY4JhOrOImQuFKLrU+g7
oefO/0NCtujp8sokvIGSIBtJPdLQF+jLTgYcsPEavgeMRThzPkTiwfg34PELfngW
x7CzjdxZRSvU9NfxL3C7RandUF0J0etb1Y8sTUXuL2mC2LlAfxKdFJxqC4BlAkGa
bRk5DutNcu6cZspImJs9uVuoNvzl5mz1FfejKOCSRygo+pOPOHA9K4U3AP2xYWhY
eV/ELexaQdg8MniJWFrXYmNzFT0L0Dbp6IEnnUZ1dOO+RhaRkdttXJl9RKULp44Z
CvX1HlrJcalQ/HOu1g4mi/zvRkBO6l6F1UK+LNWpiH10iGBYem6gDOQtW4Z2i74v
Xa0Ee2Um8EYuajfg5+u2SS1DOfZ1AJVdZWKAp5UCLouIShwJXu1SzXcNlaBPfOs2
35UTgItNxt2XiaeAI64dkaE/MGmFTSbRFdRYK04alnR1BM6jLnqY1/xCLijQzb+c
Wk4oIdVbZC1rYiT24z87lwcT8m/8AaKdAbsQcXqgJBqC+ma5PeSCu7+2wtk8j+jn
uaif5u+nYAHpnuH8nQjhtmz5B1f4sy2YHO8JZyKEfSJQGY+0oVubeUsOeVrQPtSS
A6HrJmtCqjoMtpl2i683z9vyjSulZXCCXEgNaKR6sLRIQW4Hee0TK8/ytW/uAazE
wyLZT5RbnXHA1NJ83j/FZAYnUXORz2+lzulC1v3EZalWOww7dMiDAzLq8+4GZ3Bp
CK/sEv6s3UodD5gD8UYnSZPbgjsDzGDIAI6Rnlk44MF4l1TgnIyOVXu4zp3jMo6+
poSZ1qx+4uxRKMxLiu2A3/U1MFGWVl72RcADaQJjuGGZznLtcaNl2S7G0mO9Rgkr
+V1/L1JZtHdq16W5EW/KqDe/2AbaLB2Pnq3IRrFGg5XiRwBmRW4K/1cuwz1n0yBw
aEd9H5LsbowRY3QbKoCdKai8um9bhP5S3FbLnFmxEsvJL/SeKHkYW/zN5n/WJsc4
QJOm7/aMnD0X439H/RZXQ01rhRFM7E0rnff3xmdXrAv8Iz4qQTQWaA8FVnbC8IHm
TnA3XaQSLNnWvSmcpQ+xcDmvxRB1N0r5K2C1BUPFFWcHvfjgOHXWsxWBPfe9/QxF
a2rNr+xjiuXjFF5mnKuLil/mNU0GgSJCU+WCLHGP6+kvmmPp82TPcRECCWUGwBo4
jTVluawK63MHA3NC7rovuRGrcpYBXeHsW96ZKw7PIUlXFJAW76zdgpptf8QR74Kv
jhZZYD7iwk/e3odgzEkrlXfPzek17xMl6/drSUgpqq8r8P3oiuZESCawAFi2nm+x
zt9hnxZlan42w/CwK2lZ5g1OnkZyZ80+YBRFJx0HNrSnxLdj0WGfEU8Lvw966wNP
714t+kXC47sjLMc78QPq2TIle6zDucp8m/6xczY9cLfPsCNJJd7Bt3Wxr/cfZE3T
c4SVFYYk5Ng0usB4G3AcSPEh9RsIAbvKXq0tCZ5ZQNmHfKJcj5tBFl+s0hA76oZg
B2NmhhKJcFi2LlbYo9TInoY44ZP3iBFw+ZY02lw9CHlHyfOLw90b+dqhSDcLdiH8
3nvu8iC4wK3ayHJMTyk+M/Rc/JzkU+J0o0WzS9NhzuDAGZhHBnSq+QREsA/3kDV+
fweigXD47Zcn4KRI2RdEsKae+1TlW6Oe3jd3k9g7QEtCwW6Ds6g7GXunvK/FWzD8
L8vzEWZth1AK1HDX8B1vsp7h7yNlSzjxo+MN5W9LbVqDtXWdi4SWvsJ7qhvNWWvZ
I/EZWTzfcPU5rG1E7iqiDrod/4Dlq905P/4rfFSfgsWg7FJDhk7UfBp7MN/XdOwu
IW+NwqPxlBQ1BF07jQ043gaxnO9muKhg8f8ofqXLRJU+4ORmnpM0BLalmLUiENvB
vGvhpI5tPgFioy0/Ms1Ho7lPewy3jS8TW9HAWc99O6m881uW4xeoh2vvJ2B7nMmF
rH+qUH6EN3odnKYlUW1pe5hI+NVb2KqZXDX0VMuFkhm/oT5e1o/bgDwiW8HVuoWe
oyHrRpuKvXysTme0UtxuFPbOCLL4III158MNsqgY8t3K+4yTQ5Rwjf3sxmUk0sbM
lSIuamX5zrfyXtGE8+hrt//RK6csSwCu5n/IRJFWR1LXIA9LYNDsnESBjkIKcn4L
LnOcgs1IzhLZQE6tazL04ukkkvWwQZPXbqpGIBWhnqvyCJBObZwRWbNsSj16X2I1
CBaBCHnLX+i9k4RNpnGJeBf9MFkuhXZGbnvFtmWrnHJKqT1FNx/qIlRNgszo9c1J
98FZiuKdLIurAsXKKkcGZkLWeuIDKfz2NUtVc6GAdLmCUsXRd2SJPSH2/BcjN/Nd
Ash1woBs/wJk/hCH6hZCg6zUNo5qc7+6+TOsBplXIweABdPYhv73uZ3a0GRCtXOr
BZABiwzBL4UCSeCwp6WdG5uGPuTUmLJH5g5nBy1YImPnto3UzN4lGV02Il98L4sf
CHoJTQRxZ3XYK+g1auosQYz+PmJapKODzTMdw/YN3kzcU1GoLmhMU7hg4yK3OPSl
CCMVlyjCqqTdMquKiktOIprkl0JKjkxLyD6B9UGa99r7rtkosmgNTpdEi4glVVbj
1UVq5Ve9Jb3WjB5SybUjnBUXE7BZ5/V01EPCIoDoKLJ0vNS/P33Xp/Fct4qjZWoQ
Di4NeWKElv0OaddOXIdrMjEMDfjdSXd7Iw4z+bdNEBaUlGcnQggsdlYTStVAx3FP
Q2JZ50MPziYpfd4rdTf6vjUME/vFcp/LnBCVylkhQLj+pyQbFgUkAHzkbqyZ7hFG
lOxKb8J0pRNQm2SfGA0GO1AbLnL8E2x2/zSdX+11/5rc80Pbl3scdywVqsgSUD8s
9f+vudjtttEgqfIU0FZoB5XWP3s6QXowejcofMGpjov83i0Y5e8RGv3Kmj8jS3Fh
kj1UCPV8cgMpWkdmhEUNUDKA/Ajn3LOyAvHEl5qZwvEqm/BXJrPM3FrtOEQaR8Zr
d2dRWkI+33wodf3KnVnua6NI+KLbJlwuf4ri+3YU3nvzXPIa4kz0gYO9zKLDGfRn
+il/NMMvVRzNeIJdGrtC6jtV1vdf5bUFSdey83sf8ImtGi6SzeWIrxT6L/mG/vuj
yncLj4Lg/brttvTKt+YS7NK7KskzK/spvVpoq82FYmk7lNdmz7M1fCTbPpY62UI4
pwv3pCDxHZVqAcqcCCdqurQvcZsVkxmes4uGfjFJHJIMXJtdJe6bit7PWB+wQUQ6
o32I8BZqrv+o8aqo1RmhJvobupFF39HuZEoIJpzuHjmkMF1vk2N7qUL48cV9ScMw
lIAmRd0iU9bl75qehbUdh+jwxm3VGARPBIIVfIw9Ki8IQFRKKBVQWInwQqYZOi9i
SlIeklcQFT3UwvLyUPxPsWpezSqPG0hUcSkFSoeiTCt4LIbyjQOnvurgbOEpkCkr
8ICsH9h02/aeu3ErGvTLRZZ+QT8wAmFACWBZqxCUS3WMqWnL1C+kPTasvW3oEYC2
GY9m+6lZuceY0h3pc98QcLhtowq2DnVlMpSnKl3ovJ1cbFufDUhoNglV5L7vjgaE
RgNHpd02GDdmqs1MiyOcvYfBdfqHIbSMcMwVF/OKDT/k54YKI4aS79KQw1pAeos9
5oSoZ/coi+929VSAnCEsdH9Mf6edFejatZW0NvjVIPQZ9hmDWmEM0JJ60d3JiSVF
ob48256L2MhGQloqHPg8QL+Dxu5kPvKzYrnSvkwRS36eHPDiYVHAcQPgbBaj9JEa
4S0XOqt1Pm6+wT3IzbmEGbzW8r1jCnqyDPlwE6gtLmtKkUCMz8VsfgzBJTV3hIBx
D7zTmOlJOwOz0U6IDxj8oYbDtp/omLB9+OgDrCqNmU5q232dkIz0YRkEYfUIw2Ru
pIz9gxolQFQYGc4k8XTO3+VWfo3AD9m83VMpZnj0v1QQrWzWw74B0qCoUkvpYUzm
Fu8sLkejzPXVXEzBl4nNYUqYqKhSTj2UYC7orhM5SEd8Jvjf7XgFvCfK3TQi98oE
c8CYzlrlL7ymjnSovgpG07SIikTiau3ybCtfUpkZ3btjxZNPUaGlOPZC2St+SkOS
5hzEkp96gjrfbfrihC+sUxFBBcpuZapG1CzQWGPUWn7t030nh8BsImhuvsm+Lh3/
99HXrs+zAZbSSm+xykmO0QMWR9Jp+/Nzh1pbB38LeZXpyQzTqqoQIosLHEZtEKfj
ubPWQsW7+RnlwFguI/cFDHB3RzcNAJ8CUnZoWppKboErWtYADi9eehtn2YMaMEaK
qWuhLI0bMQdnvnyPtkhVh6+i4MStjotvfo3DDZlQRyXXK0yTGA3YwZMXz77KKNOF
AUej1Vp+eVGoScglPG//aZRGJIrFYmcEzd9WBoXh1qy/+OhH205Ch3HyS1hD7k/u
mcrZhZMQOWiqhBeHv/xri9Obzdi2RsxJFWY7RxgypxXiyqH4vUO2QevnvysUdtue
f+/P3gBwz1smpYpi/42TEmWRtC0UTbTWI9+b4DRtIE/xDpjzDirLaBfPqYuO+OoY
BPfzIAjgfyRYc68+QSz23xUTXIZGns3CJQVu9Ve5QQ/v1amtxwBonW9gIKC8kKp9
8bG/Ip5q63n1ja8W7BPyAug+drnPGUdS3WlqKZl8rlaWRcIINFzuNYQc/CjmI3mw
83rU75zsksAQUJ23cY9KOmcur+D3bmR4f2C1IZnpvQ20WsffwEQMzets3OiuiQuA
xhtq4zyv+hubSYR1A9RvJTus0GWRO2x8roL1pW1Nblod1Pzxctb9lKf8kKGZAMib
5o2bk9tVp29Nq0KkizrrZktaywzjLki9ozpRTJsjGA53LqyGmvYlvbJSdEiJXC8/
aCUHuNH3EJ9Ece0XIOESck+YRDGDl79tZPQkUEsmeYpKUxwhlowhZ+q0xEhgLD9M
bXF62zdaOGqPs2mnIwdPz92Zi3iGQExP7WUaMUbFq1gc/WqqG+eFZGcCOIUVhe5U
6q6LOVLkvWxEwOrWPAH2koJauvfSypHipDiZcqlM76GcM4+sdjmw01wm9rUy7V4c
/Uf+Teg/KZ+XxkjAghm+6mlL+gYBe4/IHBM2AVU19w7AeVbwC3J1h/nEtdHYKmSV
2o6kq9CHn8mHlYnZQRDoXGAtGuJCQlfYeVHaoZZTvliMWLdGxF2ka2ArB3SCWEs3
mnrcfp7dGMixPG02xy7suLJRU70NJmiOI25rx7SAUeGpiv7rA9iW0Iv+zeM3qq8K
Fwd7JGCU/W3FH6zw8wHx7MyICoIn9RskVOB+5VXxN/oUnLSPzyJQhBY6lrhyoyLw
gfsDSPC1f08TJ8kKijuPWCtBdMTw1UQ6g4I8SoXKr8kpn+aFpD+Q3TCf6UzXPqHq
JnOMWPC6a+rPhHr5TI9bSrrUnbPgCWA7f7Avk4X9R1zf1mYeJCYSeeEgJt8BP5rv
1zZhe60Bvr1KLh1O1MXkO48ABhQ7sL+I14MIjhZrlsjzYO8umOsKEuwtRI/y/xgV
ZCPKHTWdp9eZwkjHFkNIcxx4OUyDIwJkV+hKINe9Jiz3snbaKpBVI/YD+cTJcZpU
Edq66j+YLcDLjWAKz3mZi3K0HNVQDjZp5FD81GerutqEz/OlNvfZlxwbHm/T9y5T
M5gaSH7EjSxXkUd0wfLUJIGF6Ni+Pu/b8BOoceyiGPSDf6n/h6pGlTwGh4YInc5b
wPxbbzXFvocAE0k7q4sXriTGgkSdjGlbxOUZQNX1liZvAci4IYm8bQsYcM/1RpdJ
sjAskNDQcoEMtCxJ9+v+yi/7jQVVNNGz+55bmZUKpOG7PfsindULPEQjVQbzMOto
f05NaE6a+eedtWWGspZd2YrQ5lCvi6JV1xUfJjTTtSJ57rdCYhFKswIMstW653FP
lunEukfcenxC89eAJzlGMiMgJN86nNZ6mZevR621fwSU67HX4F7QXbVR/aEThGq+
47y7JX2/AMqdnhrYB2+hnmsTC2MbADwHT+7nYQN9MpGU4k0hMYAsq3nWxc5gZ3UC
16vGkEhc0WYdQCUG4g5Y9SCM6jXhDpyV3CZm6ETZ83/GN2SFpsM3mcXweYFVg+Vr
wyhHAehywCYM8mtNIBZNKrXNJbIpBj737bkqvRZ2hlbCNQen6ve5DTtM/NavTULS
HZTroQrKOG2jxmQyMY/pUeudFVw6NY0NM3JkRZnJh+DE1MBhGjxJRucgKRyqt1Jd
UTAb1+cv2ddE0WqjTKY6ODTqY2NtqEM0lKw+QzhsZcLzqvq2G7ampADa0k7BgMg1
P8CiP04wSJfohXBB7ULQW5EN23eNVuVYOEKed8PPs53IFh8tZgoqh1ik/iguVjm3
p9AjVPl0HQL+uFv8KkkzVplvDhcc0LRbeTAKkNWOnQd1zugBdwRXzLUG2V9dStmK
EY9Hwqfk+xt7c5hiF/hoIsDO9hNm6SEV6eWlgPuCFLTNEtyJoDkhhWkoAwH9/6Gm
g7gW+x86Coq6W2kYo39kI+cHfKar7oRjtz9u927TIWvLzFMeJrICb7HFEJgNOtWL
GMPoFLlePuP5g/t4PNpAixitKvFPblObktlilHCQYVQsgw3MFeOO3f26TkZi09Mj
a95RxuLHzQb0tcpDdWfU/c4M3Us1IWTYO00ik31gqWpnymQX5WHVGCr6yXRBwmkk
uoWQwMytwzvY+nYQKWeoHLuZh1M9LzErJbAR7f3t4RTJAcK1DH/YpjQYEREotCR2
tqGDrQORSm07+T5GHm/8Nal56P55KIz5job9ZGFnOIjgvpBxI5dizM0c889ifZ2l
0sfSgUw9LmiRXf64dbn666Yc6H5X0crey8mLQzqws0OksLPYHJ95H78vsvAMHELj
vaBYrvamTrJmKJhbCli93+yOJ0FbS/x+FT9HGKuIR4hIEyQ/vX3fjFH9/I56KWcT
wztSJym+vVPdTcB9iOXCQyqeZwOvc3GbVAMLf2BZr5YQIrc0Sspcz0nKz0PblRAV
IWFWMK4N/66kMwhYv6BHiOhEMs9QiKvBWV8AnZ5RgMNwxhtIRak42wMrTSXZWgTT
E27IKGTMkq59bYZIlEHkAcvaFYIIVISwLm3JmPzWcWBnKnA2OGpITb64eVqTq3RH
O7NB+qkjvZxpgCRT8A+wBFb1JjJBEx/JTt97Yd+umQnhJjg5lVH/eN9Dv0EFAT8X
P57QFY6UWTas8XhkjERiapvJa1HPDR09nFCk7mi2Es8PuEF8Vw/EiXJhY5+J69d3
qLeG3Em2As03kIA+YkatF5VaV7XLhwz4RTtrVpdpJujr2kxBn5IVPSRCh8Vt2n2Y
L8Y1+wvFnnl00efFAxBQXirHe8DDDoK5arXEQ36wHjSGZCNAoXgspVtU9BctmSSu
FOH7zeSDQRxNO8GBZRIzFkUdVaii7l8VVeiL62tW4j2fNYAgMCLCpMivXxt8D3Xr
DZgD3TpvLWuLz+Yd8NY49d/blum9rHLzTOouoA5nQN/0UXaeyubw9njqfhdcW5bC
DebfewsOQnhEwWbVMP9JXzy932169y/pyN3kj4njwnxZFYq6+pIUrJoZK30m6kw3
m5jmOBw20ZIdqYHEHmKD7XqB5VOlvRNMK31XsaswiKS9M1ZIiPqSLewYX424KVf6
UDiG5rvXRDKdc/jVFPhbRcXd/64EfsJ3IOFCfnSsNK3P5RNLdPjn8RQUZL8ZNhuA
YULdlq1kp6LPCagYDSoZaQegxxgCK9BrLR8XFwTsAEDktnjMo9UGmqfe9QkDwSzo
iw+e2L0uPsOubN9bU9/k/o8BqARTRwoyAyu1sdqg6NZZIddWUY0yHMTKC+VHA8dH
0VPWGPUmFoq90Pym+5f67n8GvAzC/L2IGdmzqWHXSS64BTd+InmdI3yrBLko4PSA
DEhtWT43Ghto2fzYkm9vI4OAvu27Wg6FdXXSLmasWpA0LYPhKXJaS2nMfX1EEdgZ
+RX09v3NG1kkgQRg2FHVfhZBSFwxuIqsyu5oXPExk95W/KYbq9gBA5ArLWFvn6f+
XukpusqhXwrFU/o61UxvQADYUeFmm7Ng33JcEks5E2p1V/I4kLszkiU/OcHJiFpG
rL+15TpewoDtB0Uxr5T7PxDWR9TMO6aUwtuND7Gddt8aWf+djxcApvJeJne4xWRi
xINkg/h737La41V62IictD742Ex7OqkJ35Yp9zY2WTeil7EY+EdUC35syO08JWbs
RwTexvF9FlraxtDYmDVvH40azfyAsXd7YsFYMAK6mBE2QIovqm6x9r39yc+NfgoN
Kf68UHGGWGmtxYYDOVydpPuuxRpzrmU2a4T+yT/FsxBEWWEa0qNJL+8ePnKNCfpU
uvpIrZ7u8tBmKi1kAwey5qxdmtwY0dXeHJBu8FJ3E/x6re1L0eAhJn/yuXbXJZNC
GrxM8KqKPtS3UKD+bNHCyrBa77gcfzj5IWaGjvI6cPoQ+hcjSF2F/J3g2TVzNSb+
BCSv2XHeZ2ceWggjLhZQ1Xc79NUVwraReNVFYso/oFmTx5QQJHdI7B2r8FFmaUI8
FgS5P6bF6/7H3P+W+Ab8TW9dPmH8DS+dpVam51/oyZl09OZjYMe0/ebq3MXVICWq
Vuw9Tb5pLakK97sJo7fKXxwDNhgyYP7gR4dz1+2qqnsPcaCQimkmTzAC4150/oAa
fls0kXuxzHW+F+X2AB1ylfDIHW/SmFj1oBmQNP+iLWDy5zlZspHrXHL84O1rM51t
GsVWgcoxGcLFA0zFQKjMKglPZzN1bdg7nAD1nHGX2YA/k8ILJ/yC8KjFyE83/zBq
8ofreGnFhMZtE4a6AjHSya2qupozTw4vJVqSaBFixlv4TKtKhE90FaVSQ1nNO8IE
NKaOIPNFM06uz0zvbBM0q91pfPfZAn0DMgBgdKrKQuI8d7EnV5KdV3Oz0gYTcByD
eoBFM3uhY+elLpy+GKsfY7PLo5w7oG3ry/jheARabMLQyh0bOwtNEAdKvx/XC9wH
o+IyDRGXtzD6jTqGfizfqnkc7miVTj5OMD7qt/hItgxtphh2SrQa/I4iHBKrQozy
+Dgzd1h8redROw0WQYLIuFrnzcby4Mlh8kXWArEdxuVXdusO0wyWpTt3D2zu5Piy
0i+bAGhpRMdEkPeoswOSQJ+7gDxURgBf3kk8weyi6n/ssLM+7ehnM7HGG/0DtT4L
O4ZdEWOLkOX6nO9S5cJa5Z6AEP4B1d7IKRmvhcNCUAkQPjF3r1PW20DQ7TxeQzP3
IZyWuPWNDVcViX/nYTlyHcR66N4vWO4FzAvzfOwRbGl4koxSG8Bnfotu+9KMzzTZ
JSRGMva/83igZyJ+9Gstyr1Y3dvTPR61Ae27sJn1I3HB4X4jfl8Uwj5woBECVy0K
0P2yMp22/iqazqKaWLFIAcvhPMf1iY/xd/rKu4nCKQzILdfu6jaJmC5mHm0UCK8w
ccm7uuekVNFhXviF13yWffBH84YgbbT01AX0KdEjSM7qAVHz+Y8xl42T+mY1FyPd
4YEBngQxyfXsQXhjorg7wMq5aWznTHkPeAKWYzApxYnEe+wDj3+agHDbFTsLrzjy
hcSvZhU811zB6BUBPrWkdP53KdUvJTaJX5sMuSN4Y2VlV3WmHfYr7gHd28j40Pnv
2oVNTKwtQY7H8RAC3K8lhsE8DWWHqIYGU4j6i3umHoM/+xeruJ2CWQzGNNNEb2fc
7nOW/g52kH8vZN/uobbTd9LhwftAaB/r37iypX1+Ujk9Xag8t6yCeWKZuK5O/XRg
WAlipAwl9bkv9tvur6JfVQrfSuw8VL1N/cCI+9pZ+J57TW6wQzYByBGXIZTFxSAN
w7bQeHCouRpEGmrFtI6at4JW7QBz2CC53cy54DRhH4HTFDUxm/HIAgym4nUpwjsA
sHqmc3fDJb8jWh/VMgoVdjZjR8babuZQBhSOaVb15WvJAhYmC0pRfJ7Xfxmo1irx
36Pb7BSZUdz6WMJq5N+Fca+BkwJPtDdFW3w6PRc8hM/RZJfhJod7Y3lRMB1RRhAN
rOqCVNzH5EIZ2Ny5YpKCLHlBYnrNzl61aE9VLXN2tBpat/B+IgNfyQyejTrSDX5P
4Smt6iswj6RKgOOefbXvFswKA4vaWzwpBDMAXanJVnk1DJUN9BpWeJHrmlk3/vQK
BaJAH/lI+OAXlR4iZUh8n3uKvBYBBVYIex9sRPTAzmNmxs5hBVjc0fMAewM6+IxE
STfrpSqnd2rwETyN8tbGfDsRC2ndTcta5eSsFqj00VFObibBQPQPXc5ziqSwNo3L
GDff6Y8rXlwZyPPIRmzqjr23B18uawwEizNE+0QFZ11/xKYhLX8lKDizBiER6MfY
gWI4V6G1QQrddi4jxcf9ON+tSmscv6R44LRTW3B+XPUuhcCQKSljTusY1vpdKA5I
VJrBFs3m7wUc3ZiW7KBP7NRICfkxrkxifIVoHJ2MxBDgMEEbG2HYZt4LuYGg1jOq
5MHTy5FuPRf+9M0wwGL3AkFDfMxClL2EiNOVcRLe6za1TYLyOcUPglMtFzOUTl7X
QEXwBkrB+wLNfd0ZzjoPtxp7KMs8b2RsIKaR/B1EDvOIKJvc2UxLHpshAVjqvCDw
lFBMSwpAOFtUkWE0fAr/njch7mAPwm9XEgjY4SdhMvh2joyT3IOaLAThv+j/HZf1
xDSyPiIPewZserl8soHVuoNoC+0IOiJIood2U7azJk36VlFWqjUB48weTvusyC7D
9+QR33gkaKRjhFgoTtqQrz5qPB97BNlkmDhrLULVko65a7VD2nqY+6lPN9bncJHE
Y6DM1llLX2bwWUbURMS90ikIYk9+VDa5QuhdguYXWZGThIt7KNhzyucak8mw6M8J
EBEuj9qLUxcHNibvOX7CwXOuo6x4eRTP570VdWLLBJ1stFNxnlp3tgY3ihxEL5Np
M0iTNPGWauH+P+xxmB7UOxG9PHy+C5o+4ukTtmbyuwFmrETSr9Wc73mh78vywNgP
vtyYxYhUBAb2dW1ZFw/WF8eAq4IKz3cQjQoOl9Ix0kYiEEp6yxXVwHqqNen0Y3F4
1Jz8moEWnlWVtYc1MvSny2uyNjWnfFCAhDPaFy+fjOs3gFsy20bNJNWWqBJgH7p6
zE/LT6yH5188jK6DpAk1QhyKOLmNLINp7JFTZfX2MmOAuG3ZVdJGWYNKAyx0aZpN
k5VMPF7F7LL9U3dGbvWF5OA9ynCWOwv7v/Nbdf1emV9IE87/68dPyO2RaEak9oGe
NMLJbHf0mQl0nxNMcRTtdxP2Prps5lVjFv5tFHm7UeCUeLijxRYZnTHmZDO+kLHF
tq/XFxBnPxya+HFyKYSUHNgw/fYFx5axZF2/S9W5lJNpEILl/kFG2J5hYWJmK3/v
6z80k7Uj3hE7yjcse+Z47xKdkrkHMFEFvoB/06cBTrBtef7w/nsMVH/i00/ol8Y0
YDZyhgSGX+mk0S7z/36x86+86bl+Ahh16OnIMlOHCIXR1SkV2YY6I+XfjRG9FWSQ
oLN6V4TArgMA344339SGZYccpyGEq4dfXRSd+jLNMxDloK4jOJyqk7msUtt8wWNa
otBhGguNL+7izltyv1w6p8SrpC7Fzxpq5UjWixhW6jAQ02Rl32pkxDEQ0/jYVwcP
V0im1f2OcIYYFGwj9rY4u44Gnx8Usw6vO0xUHYW6Ai81b2eA4mSgVYtwRWlVzWr0
DQrBzf+k02RUYXvb/q2PsjQLq5muX/2W2cax5xouRriFHJ8rYS37/lzy/4dAAYiH
85A82IaCOG++kE2DfOv1syGq9b5IJ6BUe1uD3AexoJdMHCFajxrzkmMtpYJ+Tvkr
twKt5YPd7KUQOnF5+tgVWePyVQD5kX5vRvxOo+Y7JshtCpdXdpfectecFGdeUdw0
2ZvJIure4Z2+i2T2nJY+bOUgJwE9uu1uuZIdL5sjBjRZfQEcURk59H20e2ZaYDZc
JPckildIJwYL4w4giKzQ/dh6KVWekLaERSi8e9AEAnPb1Hnj6w8TqsY1Mit0kyIo
REXhZZDfNe247ET2yN3scozhaEK3dsrKKeHy2HuSa+bYf2ws1rqfw6bKmqp/uRxn
8/VOCMDEzuT/dqhHvBlZgBQJIidp6br6sY2Dz6eJ4w+cZxU5QZOBr3LUpejMVthv
WHzxjUmqmspjBtuzxCYSgg9Y2cmwx1qBdMhX82MuBa9NZ2xdoEI90Q0fxMyuG9XF
suqOQutCS9c6iDDVbFXb+Il+Yjqf2zhU3VKkc6be8Z9lS3fCQYyuf/SlvGX0K8bs
Qus+Mokl8nwKeXx0aBYALaiqqB/w/k7h542X6b441M53xtSU3Srne4GyQwcUHRLl
p82vxbKARRHRiZEx/l6s6RLo0f3xc4BEvXOmoYJi5EafPAmzasPfLExM4O7UtWHC
LssUjGpqTk4sXIPKy4NCsDvdLSQuFRND8gvLPqw44dpeoOQGydEWXAd/VlNDxILq
1Uap/8DbN/pV4enl7nVl1cD7Intm82STYKvZ4bW+FANHks6imGiVZdOB2vv8Ef3a
zD+6k8VBK+ppwCs7hH1hvNatS+6M2Iyvqgd9IiAT08Q4kbnr3Zx1xUFOeay9Lihl
1F7da42hb//7zv8lOXiqGskN78HNMXd+Fn3HfZ7ZZG24Wy8b9BAtHYw9bnWmTlO/
UT7Vp95a+bTAZ931fURbIkfFP6JBz5rxLt70QnFsSEkdlz5S8EC0xtMc9EFnqUBO
SZqh8owh37iKJYMVP4AO+wLJT7/HkgwuspFUSXJAXVFQWst7gR6TCvhRddnLYE/2
94FaPsZW/STRKe+opO7uSRMSSThG1GVRSHlwPl8zEiNIJK6wi6H+eAwpSZmI39tg
fAG8ebmh81ZAGa8inOQ8zeDXddO6pWnAextYNaAHBGP5kVGU+mgrgnibYOcyWtyc
3iup1i8X1V6jQ4cPvIhfy4JV1IrAE3b8fKoWyQDxL769UkDwy0lt5AvI4764z4tS
RYOCGH78sLKv0J0GOKshu/6oPzQroOLgF9G4ZTZOz0R+JWf/a2ArtcREUrrq6NJX
HL44p9PJsix4US5s/VBrhwLWyMOZQzIFqeGuZBkF/nisydglEDQw3h0mijXJ8JG/
adUJhUkNvKZfj+wu0j6RVqKfFkKjg9QyEnKzLyPvvVmkPE0OKHjIRK6ym+B4A69L
G1IChgUospT28KtaNh0xxOgR2OUQFfncZT5Lughm26hlcDJ+0lWsUx68q6ae5P90
d+v/u0Bx1xGC6ubkwcxx6m5qzMahmCHAALy9vNqH1rIqlA5LpBOZL+Iu4z0AMsQd
DeKoCaK+u51oEWGsEszPyEH79JEFam88Hg6ZDYbvSffIt1RfphU+O70ntwl3utae
6GTiYn6cFNSx+2CelcizJ4CWy4eKWBMn8UYSaDicgx2WvsK1Guefgjfg/CgAx+k+
wRnnZz8MA3hvpQ2kk6owcUb41NqZpamv/XJsx9YqX9bxBTSnNQQUd9uYl7vmumyk
yroRYYM94cqDWhbRoWnxi03lR+Jep6Vrwm0f3VZZVLsk49UGlXCLQ6hDLtTMpY0u
Kfui4MDIDP2/i2ln2aglcP8hpRpbb5fI7Jip0r7q9oZ211I/UVFbmMIj4Unsf1/h
lWCmMNW/uNaVQ3eKMD2h+fGv7pKewQ/puzjdNl/OMQMO10DTJ7o2QAmoRfCCmf4H
+lXuVyNBRIcfW7sQ57ryIemSOjgeZwLyV70Fnp+eSgiJkwvlR+USFTIomrNmvXI7
+DUmmL2YryjrB70YynHRcPPW6lQ5ueJwnShtTeMOrPQP+8S8kLaSCoOtD2pjuqkv
PWNsqi2N9fo6sie7pOmw+z6jL5TGwanSHkqPOFKknknExavY+cPcaSJyhTnNw6c1
ruj7fJV5uMGh3pImjfQmgNTtRUi2zxa/cyEkhMFkg++XxIJyX36sWoIvuC1K1Fvc
uPTzNu89QvaRONNQQ6RFrP/TJzK4lg2xnpGiPa9iWAVtnX3cob2Ke1/nTO2OI7z5
J7pjMSm2XQuCw9zh/nucOET+VqeU9dbZ7RIPwfmK8GERJ3oQdoECcN6l7G7lhEL/
32Xl9Ke3511uwek6FsV2CWwsVvUJhOAnT3GZVq61D6MZ/1gmxEdxgwbaQgndQa6a
A+aMiP+4SXBb9I9C/NXRWYZ1li42WIud2csINJ9UHOT5H1H+yl0goA/LxmympOaF
JuP5Lj81UBwvBhMNeFWTGgGbtzaanYcXO1KJU2fBbcR+NzHwEVEDQdEpH3e+6Jxs
wJ+2gDXiy7LPvnuTclxLlvRkWhV5cB+1xK7PLLoKyfYrkm/nx8RJKChlma56HbX+
16Ey1uxE8k3PCTah/IFvT47LumP5TEsS4vOamcZ9WJuqST3MNnGQx4bEmIGlKBJD
8+cS4PBbJ5h0X8jX2Nh7+j97uDOpqqQ+h8fkjxN1Zusf8+t8jghR9cmdOjkJh06i
4f7gSoBSzjyTGAgIpT5UYkbfnIGk9Cgeqybl3nO1+olBkedXwvgO1/489fm8Z7as
eNKcNYIVL3KC8lRk5cACm0viOw9Y1htm5h3sSMSb3cObmJFzXWCJ6FIObq5TQ41r
tmHs1Eg4k6r/r38fiN/9SYFM8PhRU8ZYzI+nS3MiLl5xlscxyMRQMyE7RxFkPyRG
YBzITjxX1gFJYKW0VZ4Ntex3gpYkYcse5xBBMgNBPPwI75FVxR4ghDCCK/CRcynK
22WFdvbX6ZdpGaaSkVcnEukAg46oxvDXebetg9BjkiLfSMacaR237qvwQRdaUw3E
wWaHoUo/54BmWVcDe6/6Ep1T07FBhfZTBoI+luoPxYprvYAlwmmf54AFL2L2mKac
SVG/8ek8YpRhuJl25xyXTk9zyzLmo68rZ1JV9Fi4kYdoDQafDK+VZ8lOZP1c0XI2
ovUatJB7nqPHOMvnZMTrjzfQzAHPZPTXl+D5m4wN9YzXJNlnqPhIE5fnIWvvW/a3
YcS0/2/ZPZMqhOo6nvfi2NdRvNHLG4+zOSHoaSv8VfLReHUqx1FL80WusSJZdX5X
RiOTDSFVkRP40vI7JoLc/+Vo75Kv+VM/tgow8WoMnj8oAj1qAFLu37RRLsNSqVhg
feEDrhkINQAIwsPK5c27ttucKfrhr2eQdYeTVf5umOlyO3J9oPgu4//7albRq/Rm
M/MSb04zs1GqbGuVqMwizIekGwe11PcWcNvxOu/etcc2yT7MMnO6XoKS7WxwmN5O
qqMSFDRIer8lLIFwjxow2hbWZATo2im8dR3fiRYGjgQY23+NHpU3h4StskPVC6z5
XnIhFjM70T3tcsYLzgrPuyXkkF99XEvyAREsRx5kIqI0wJWt+T5ozhnq89ANM0cK
RUP542PRTgFu/+xeWf7oTnnXT+IwemyFEn8vaKcCpa2+thuyYF9MfREGgXIXuYq2
8b/MkcG+LfFDOZDc/tIZd/7i5BonzgNazI7zSxLp8suZwltM+1H+9xqcHk0ZiF/5
lvYxk0prJa8kSYoKDUVGYOSYWrnO9xG5z/DOar7ayzpBHeHYgdpZD+UJp1asag9L
/2jhG0nhTjOUwwLr5tEgfiBhjOmag3gJDquQRIvPEhXsODiJvvOw8nrDh3jV7/cF
0cKviEySkaOlzkdhi+xyyTwr5FXgS/W4gDEbe28wGngWMxf0k2mdGZYxhlYh3H+6
0bTWwgqKBI8Nzs1tLGtUU69K5wmMKaZaCmTB8zd/z65pJTH7qWY1hFVZREROwJVB
4KB+M40ZSC0pifebmSknj3SAa22ilvUIC3g+qqy0Z4tdEPEvuyNFdsPh8C7X9Hal
5lKALJja7uYVoQ9EV6Vm9GSlfylmTZSO52/DjGQ5iPPWFIkA525jCrGvcyvjZ5UL
pSz5h2CtjDpdExMJ6+g2fVAkpXg41Pig6QPiPsJE7vhfnCgKmUXUIWLPCgSd6gVd
0aNIZ+A7bU4cmDW4iDKWVLmL8nzjWPI8uk/1pk6wERNZi7twPEr3r0+LzjfbPg/T
/1Pp5NKbPU4PEIHUcideBaI4NDdM18Sv1hXFsY0t9pS1S836Nu+tk/YKi+2agFw1
CuwwSs/U0K1QvRf8CVTI2fWxehvSwKH3A716pwMcCemycCPqK5+Q2KaH/AtF4uee
+0xK71+9lUHBo1WNnTTRCiTiYVvnkQVnr2+oaDufDGsNVzfvWcL2u4XVgbnnGKXa
tuUV+y4D98gRLb8RGCIUYUvujh3qrV70ZX1yO/hY02jgsa55QelmCMDcuCgZ3nuh
9eSaZOX3c+fka3QOfhMMOrp9d/um7t73w+VFpaeAKTRlxpDfX9Hm6xfze/fdUAuB
qAI30NmA9+Enbnc+3UGOKnUuSkHAV62rZ3UYwel9flQm/zFA3Z3K1FqiICCdLc7q
U1kChB4T5E6MAAENk502vWKiUOpaI8SxkgWRohxhyLb6Ys2KYjRb/Oz6HzQ4isOH
8w6nRhZPBKRYm8FNIihLsoAd9i7iGkyN3bOn/8JnCBdeRScn+H0j7XPVol0qDxBb
tGeepKV4tq8dfGZcJpbk9dGv09IMLbDM2szckbmncicE6bHg+V+k1mZRUEEutof0
MJx34UancO1uFRxfDKA2ksVluRvaHX5OG+XJ7ieJWhI9Jea4zmMAmkE5tvoKIc6y
BQHC3neKcoYBggkujKYc35XtUO1PH5rWZdtPlpkeZ+NofICfr4CDT8T926yq2VX9
rfeYTeEfuyPKPqROhCqyR6m9SW1NfVdZ2ysc954UVU6N17qvYonPjc/ka2f1yTD4
88Aj+aKjBD9lXteNsZ7YON6r7qaqLp0ZTooKuek5S4Hplu9ZF9YdwYhX7ooGa3IE
e48basnJu0uMSXDVKa2HUfJHkGeNbUfbBytx+j+/IghdpjAoinqTWOgk/FXsSggr
xziCqxnCTLYEhRHebrsmjXyjfpI/fTSeSLk8HAXi2iQGLhUtAALlo88PD3B2gjqw
29gZgOEnmTpoaSEM1bxRJSX3BclrBpHBbKy6LDJLuT3DwFlndYS9bt1qHj/MpOi9
c1kIoatAZ+N4v4TO15HUOLysk5XfQ7JOjKt530950BoGG7hcYDeIkLu7VRYiBItQ
6HMeV7kDNa221gQHjROE8EWDFJXlxflH9cG4LBz4d3hOxZoeRUeVFwr1xh/eKGd+
t60E/I3uOauv+gv/3AXUBrpkorQuO4Bf/njQFRQ1cjDqDFrwqqvRAycZvJI/wx2c
9phYaslAPotuGaf+lYZhgWwlwFiCDGwIVeabtgZguE+agDqvVfotmr19EtTGnO3U
vOLldEoeCtwJ+b6/91ON+i/I5D+NwqQxtMjYvhDC9n68bOy/WHgAptCsCEGx//7M
K98xxH2fMWa27HRdPUOUYtzXErMpsGBJdvvVfAv4++ZuKncubxR4NmOjxH+4QjpO
eBlNag8Kp5j3A5hV8ljUchPmC8Ggvca2Zl6WIsJUhaQtkoOvUMUUU/Uo5vX0KanX
UkHRCB0O8tmyoqi5QF80OhpAHfUXJtPWTA4RYiX6OrAxyd5UNVajyWSZn2QyTDMN
gUYafXCWfOjZZXy6zTyxAs1VfieEb2bqiXeTkjqIO5axn4Eb8JpE46Sth86YpDJb
k7NAa6R8c/hysriiCM/5LuZO9J+UgLMR7B/2dxTQsU4ayEjST2ICmCdlyM1tGQIf
cZklUwCjlwVXDxBeFu5qr+vmMgr7jQtV/uD8Km0Km14Qi1WyQyt5sfnsXdTYb5Fe
JuVCY5z0a1V9D6VdxUUxYd//u2CuXeXW2nrNL/z65tcZU5/Jd0uzydy/mrnYGV61
jTBUI9m09QBpeOgwGSQIn4UMsbQvTbgIiO3uVHuUtugmggSshboqhk508CSpGIk+
WlvlaLUXroZ46oLkcnL1hHM6AudxI8+9B0Z0En5uHNKULbvn4v6WzDjSOSSmawsF
a8SY+h5ycfoGhHLFBwjrZlizVjnbfwBk0tXlnk+FYyh0KTbszeagebe6BQDhqvlT
LjNEkN72bcYANbPsrpiZ0vyROWrb3NoH9PIAmejPQljOninumK4gPdb+XyJfTqG5
0dMWAO6T5yuChJue+fEf4OCZAFMwaKlNNBGpw+YWlETun6HxS9O91LoDzrVMt7e/
8nYmRwf95Er5nt95KAl/85NRXLQ1HCpmANv7yp2TbQSQ9tGbML4paLOSSmtxcbU0
e5MIdz0RwwS/Wd5bDo7mPpaNWyyLP5XticZRJvAQY5FwVB6Q2PmMs5NIvTbcBqsK
hE5Vq8mEee+zFreMn+6Yk2HWk0J7tkl5mcFr9abS/g/F+vedwgg7yxeIIfNjYUSP
YweNIxqANtU7zGy3xyfIY4PYKCuqho3AsiixhTJPjRD9GamDfc3UBzCS7jdYfLZY
7vcd4jDgnF3BMlgxV+Ex/vycJcMB0b77cR0kVyeo78FnJG5Du+g4pfQ2lpxZtPwg
oPPTJXu7ozvNy/vkY2/FcjGXOYYJO7E8DjBPBpPHhpac5znX2Y3qnlrmtynIBGRh
J9thKJRz2O7l7yp2EMf043TVbMqXHIhdGVqfw/SqmMi4dGpVt/+qTP8Y/JEQpF86
IfIY+FJo9ze7+z0jzneBQe/dE6fNXhTYYRg2hRcWEayAeCf5MC6/wNocWDUroEGM
nn4n1tuvV5dxZ6i0vdx2nsrGPNdf9HjVxw8VJ4LoztocFAVKqQaOnSUiTv2NEYID
774xJSATfwHN4u9u1b9sBCzEKmvj0aOvmlHXiabkPve6NIyAMVWhWmPg0phaMV8/
BSijI3DdpZaxudglTJbSbdLToGAJ5SrAlObl34Mb7aJKMViURx7XP1fE6xgDRCwO
NpbHlhrcK2G2dZaOAwnuhhfCpnAg5YcIGHGM41+/04xcsBj1jYWl1iU6R3RVr1OX
NC4n/U/cUxSOyvMriF75O4p2evkebSXbOzN4tslm0VNt7+4WrYRPVc+vXKUuRmcy
ay+edhUk3YLI3csrFV6vU6nOwRKdvuj9TzJkAjqKBRwT9lLv5VFQBkPrB45agCR4
WATBUUf25cuqfLqIZ6ivy5iYW2TAc3lqc5NulTIMWS/8UCtMmYkAM1ZA/i37j8jm
bUBaiqeIXKRSlIqlH+vwckdPdqNXgFUcWB48ab1UQESFXTjCZRiV32jlo9psPX0D
mapyvCQC74GMz4rdg/bPtxOHZlwxYaB3ZJ8KDkcuw2fjIBwMSrpKePczJXkO4KZ2
kB4HyfYx6vRYges6bPtOMwO3KoZKAHs/p5b/2T0qBKpgxuo/aW2e7yFAooF493A2
Pq7namlaDQoQnJA5yBUjjePuZza/qkb0nVZRbompD0Hf6LhaH4wjLLAdwgU0sj64
aMZJhhJzBbwFx66Cut/JQUjivDdY7bE/hJqOYMInA+Y0XHILadm2tz+0q0X0EyLo
CVKggrKhS/2J5/gUs22WSXHSaC3uYpx9d4X9bHlBO+sRnN/FMqvOlmeXoLeLPF9o
LS8Pmq+WcMiktfLm3T7gEl5AXCmQts4QIkIF16LeM3u7rFQFB2aJPMjMRcHqWjkt
zUcu7PSforBHE4d0gs+eCaGNoHFCSGYRVw8Hhy7gzaPdA62NVyFipjSmwM4rGbit
HuiMWwxdX/KASSKT3jyX91+2SeoKr6GIyOxxAogiMe50TQNsbEtAr417TXjPH4nk
TBr9kRHXpk/P6lac/GdGvpBiG6UY3oRlCnWHwFZd8dKEZOhxD5dLI/ntbgU9+Egw
koI152SXcMinvbMGGnp0L1pI3vVmOMagDN1Q7q8dJ6+W9O9kzAKXyn62hbr93gEA
IkhzONoP23MtwbCxQYEc8Y9ncdRg+cVyyvspTpcooQNcasSN9YnRDXXxnGXMD9nZ
pnWCP8W/9swYvaoS3FvliL1rDDi4oIpc7VgaKg62Eu5lVcjNbEYq8U0j8Tz3KhbV
Q8IVZsUfSWugJYd5hby4t7PaLwxaY44jDzOxclnePa/ARJuanarfiRHriOyD9FcI
2FURoSwF4k70+mdY1isLegEfRxPFpjmtVVHZv3EUSXewpcqFX1PItemPpMh3daoq
iKM2znfZhezjLS1UC9qa2kLnhVf+3ft1xTijS8rJh7yXJumRzei9WaU5QcSWsX8d
WODJ/Z3cF3b0Sa/ZRs009Rl2eAkRuzE+/rvww7WvjTNF817pJjrG4m0dS+q/Zcug
REYM7ewDjWyg2atU8I/fsRjpvKOu+xE9LI+lfgiPsh1NpOsv63SFg53gsFm7ToVH
iPm8GiT8vGljrVT4nDqIoozaPzWzzggmsAWdb43tBi3wIgA//v3J2bQP6FSx7y2R
xPRj+fZgwTraQtAzhKqOXLW6ku87I9t3S8yY2s4kj1Z5mBoXTuJgzamciEzH70Mo
TteAXE1SmogfbOwmDZD8+fEfbKB32EInb67ONmYNOiE81YxyXo9QqDmVzwgYCVGo
EEgVlwKnsqc4sASB7nDyCdflQzy0ckJpKMnoV4e9YDP1FYvBqWUE+pZ4/IThLej3
Q8jnSGm7Q5FMrzKwiN5ykzw3WShNFThHMDZMWSrZafkOU+KkdFzyvJzfm1RLLbfj
0lOVcZb3Q9ikej8JdyQ3xQbSt1tkrI5+DK1itDp5rrZYlcgM56Fv5kjFzwoHJfPm
h/bjLla8gZ2Dy69L15xoKF0VqchxJqM0P/KOfwoJV/a0FnvLXv1PiASD3zX9252J
fwGqgk429pYrAjIxRdfoG7n1JWZYz7AJwfCqsEAE1rzyYVSCdsw0JNgPcZcuenyf
V/mT6yh/tf27K2GdAHmFfLR48Z6hvwxwsc+OUdWAzYcF2+2THqias+zCxOaH8zVE
ZuLZILpZreXdyUn8XKsJX9U7FS/h1hpcl3L+0n6oMNfmYR53P/G8FNeptPsFCMAF
kedG24hc68TxQN+S7NGRX0sYx81ypA2kqZBHnU+9fKfifR4PUS/nFDVyzskI7eFW
nuIt5hL1dZLPvV4COGwQqcseuW7DzRk1LZbx3G6ewJ7MyzpzIzzb1ofTJYWunOKw
78t3j+yENHfpFUObRRt0mIUT/cq5oXhUKSXoDOpn1RU32ANZmRD7/QFd0fw9Pzfo
ZHHB/8DF0692x/BGnxOPwwaAVnEl/B/563lAWL+1GeMUa0wTGIGgvgZ3VTQbuq+g
Ef6zqMPMTvXR/NbCGbJrhILxpJDwDvKZXV5NhmnCTBvZnDNcSWge7Dq4Na4Zig68
nssOWavKL4b9aLuwJzTUNsSGe9oKUf0NzJq56IXRt6QCXJLvdJBdTsUpOX9wi5sy
biRvb2hAxEseu1WgqhW4Kx/pITCYt2rwzhupGFxa2+im/Mm4v7Ke6U7hXXRNeYla
/IH65rTiQIu2ch2vxlP7+RJ44fBt5PSaMfke2vi0Mevnlmtu6pd4fnGmLs5XpKFv
mqWQBpL7BKM3veq4hOPXC0elNzekZPy7W5RnNNPZEyMNTKJqXI7kLvKy6xFXCyj8
QzC8aPeVfxvThWE1RuSegqSAMWTa14pAmC3iSHZqTPeQ3pxaNoDDiooCjxzU2g2V
6gPMAGR06m5/4HsUlax/BNYrl/ZP2+tXhAW0aqclW635+49T94CnsiMrDzC3UGal
jwVdyzi03/OY+DizfuyKLZ0FDcRmGbpqsJjScv60kZE6c5HAp8V018v/aTK49hEw
MJFzl4AukOWGrrgBqkd+9NUlxxlmYnw21RzNYU6snd3IiOFiNu0LMCZdbb41tIu5
GneGnyo+6Ax+swSfQJiwifUfGHnyZZupJLUNCCY/vTzKM4Nfx5IU6gWp6aTOQCZw
gLBWPvnRsRDa6yMWOH6N0rtsSkYC8kmQoJVoNbzaK/VQ4P1ygHa983ayYtvKXDHr
B7LJhOmZ/CrMaxc2SaNplAIXfCL0GyggUhr8gRRUlRxdephqK27BlYF2IbboecTQ
HryW5z8KqSILQ+G/k2vEou6cbmh4v+BUy2HilPW37oLpZjCVSPoerMeuVyR2GhH5
Pd3oGO+VPwc9gbACIpIvQJPDyTXfn/EOfc48MT/tF501852jJkEJ9yq0yDCWs4wl
i62WGdLtzpNyYtp4xpDPMZCN2CMEzpFFSPug1egVF728DsxmheDOFf8kf0/1TZRc
92vTMd55fHzJNgAhcxFbkt4NBM6XsVo1qYAwUHB0KNp/VLwBydmWPqtLVp9QPIFg
FFlM6yuZDlzJc4cn8RO3iHQ8pOCLt0SJaGEZjSPUhvsTCctz6X0ro4lrGHHs4F1V
bMn49Qhx9TtRxLvvnCH/hii6onVtZqXIdxObbaoLvtYMHg2B0cTooimGUufekIEW
yJt2tYIQkV1IlV7xHo7FjdT2eEIsyIMh+l2AnJstAvjd2glVaGJXqnWDVwX7toOy
Iw6t2pzpB0UIJAu+iK5yloOct+YoPDf0DczJ8jlKsD/aNl4KWYVkoBM+vJY1qXie
f3gXBctoH1DdVIoica3KnwiQ/o8jbrgMIJ82SNJcTmWGmsy4CCNTN40FKug1AOx7
Trjh/x7x2RxOg/WyrX8NQI+ISAbrqRSbGxjkDyg6SaSDWeizFSCQJ9TeCwGR3D+9
ZGDXJo6eEGpLTmn7kROMAxA2rUzCYLN7ApCQCzfnjr8ZksNq9aCFW39eh/4fHngz
yGDEStijYex+ONAqgRkthon7pT7Jn6G5WFJSuc4XXTdoQkCbjEsB+Q9OoZDFVz8b
cNM88wgDcGyTnDc1fBND1S3wpQdD4h136fJejlp6CYQH35ExEByrcSm6z3TD22Xr
F0yTZ3Qbws4+uIKAECoAB2ghkn/oaz1+L03c4tmiBntKy9tir73M5vonEf7Z7M4z
r8hNVp8cSRQuagLa4gd3mefGSVGx7UHAW745fy3eFuQR1HD0KHlQ11mJvtTrm7xT
cpK5JpxHaFwDxh1fSOir4uheXyq1c8dHHIgTqyoN9KeWuFMIT4xxrBChI1ZgvIYU
SgHsVBoYR3QT1QBvvOjkmqEQ3MZVQiYTKHjG2atKlQ+kN3P2x1XNeNg8iLg9JgWk
`protect END_PROTECTED
