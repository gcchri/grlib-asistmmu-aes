`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7v94s7FIiDAQhOOJCM/U1f0yZRAPJfvcQHdezrubX5CU7Kv1qR1bA7965yY5wTQ8
q0pz2Axe0w4bN7QMrnk+mZZejwq8UI2402w9WMbuY8uTAtZUtieTsnQ+reKzT1kV
YP7TEzv3Bfe1AvSTV/RLulUTiEs5s1pdeb3FY+1jdX7C7q3KgBUrJ4NTAhY8eIOH
+G6gEdDscQfaohX9vftpdaXOwdcLhweWAwQdqtwsu98N4qBDN9zSlNlBbKg32wRy
U6sgefoFBlNVoZ+zND2+9BhK1hMJykt6bgMTbTo1hVBiCu+ypzrnuk3eCUJ3Vptd
3SuPZX0JKQgjehq7N1ebbVYjtjEYal5k3MUDGUe6to3IN/udjEy0brTt3nOE9U2I
mYyNXLtgQr2wLbJGQmtwrxqF+ToZtsYmwNw1R5aWT+lgsoKkK/oJWtwb5cQ6D4dR
eRBbwBWqt+cqo7+z4CYhywwEz28R5LGWsR10Gk6mm/sd9zpYq8hjh5ieRtEsOHKr
0C9rkZr7WV/SfTnzjO34hflhHEl0kuQHPguCXSYwd2EPHPahCu1m1OuSUbLR7Uqd
Hy6NipAN9LBckKFn9hKECQ==
`protect END_PROTECTED
