`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iWLWmxigN4QVxG5sgqfCo5tfO+FCM9LnWMTM5x7KTWx3+CgEplrHy8VTOVZwyqv9
0IS5rjbaYhjScuCesu9wQcLtCJ657OflGQpbCpCucZr8R5MVLTrN+MeWaLNB2tO8
iv2iQTAJteByzKW66SaMh/YMpinavzQO9e3+b7NzJ/ZAT5dLnexTAaGUS3bRQoLD
U1K1lHlAQbBJ2Gj9nz4BWm1f3B5Iv/mqwgecWligi/+jUHQcbJrp8zJm4ghZXXpY
p3ApQQLgLo/ibC7pGVYrw2Ec7YnTAwEncrYdcG4SMo7CHxVFZeIcVbWVQqEqfZyQ
O7vbkHN4NANhVhmdKnEETcWrLpjUaV6yI4wXbO47+SRGGAXy+dq2vSeYioRU34av
2J0BbjX+1Lj8kM2GkD8SKVJQT790JBahVUEBCOjtZ/9YO1XqHBzOE5znndsylbuZ
WR4Qc5B/fXrozkTlqSGR4g32xpVKo9njop8F8E7dLo460zXWR0sqYTWM3TcjT1o5
mkfDN7p6GfGhoQ6o2plh6L5ByVGmemx4C6lRd+aSEzQ=
`protect END_PROTECTED
