`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RJ04CxJrl8aeVUQtKJUClVATyHKheArBBL7tTa9peWUoFQwXUEhiz6O0vIRT7ZKr
HoRd1uFsLyTpbZ3RFtzIh7aBIXJbDKAtRbOsfhQMb0LFE1jMdyqgdCTY89IgSCDA
SDPdD0YNOYr3zi+nLtLJtm8JLZIvIcArVYW/I0d1x5gD/TfHnV3VmDh7n0tx4wpm
UMQOYhyjNyn3tD/w1n4f011acKpDxeJJbZjScaVksu9KqMALJ2ggXlFhpNxcjKFX
E2KdhL3xSIbKtbq+My+z6O4Pmn5ZzFBMSV4chdtIgS5E01wWQRwt4P2XEgKU85xP
NMYERTAjc2gJr0DBOj2BtgTBGCNkvW9nsfVKwAwIYcIRHw0kHdJEWiOgGCKTvf3t
rpiXmwV1O0ftN2Iv5eKmuZnqqG1SRWMDPxHExLJHRJH+E2/sdTuS5tiduqJy6FHt
kp2BW1silZNgTffTBP4nYqe4kZt7ZfpzKlI6XXeSYcZjrLQd6lInmDyedDbKiYoR
5rWu0ryqLdX2r/tJFZhsM3cXyxj1W1E4kbp435y5iZlUwM4SDiCIKjjcKu0XkwSg
wzr9oBo9QdWVrjchMLdkTZ/TCw7caSt6UIp4mluHMRM=
`protect END_PROTECTED
