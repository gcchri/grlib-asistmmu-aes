`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YkIDrtADlLKhbixgMO+c8TDeXqxf7No85F2T72Dgz3j8jgyzOR5EJWbupxsrFfQl
50AIYb+BTvl4t8sZMPKJCaAXEz1x+86WjXU+rcqeMF+Sn2BN5Qqne54EtB86Ls4o
tRJ4RrW2QLzZpYF8CKOtlwGAoYbO48cJvu6jv/pmQee7iRizuyF5mwlvtEnhAp3q
Z2UVqY39qAIcz/JwAEG1PM16h1NMasy2xxnDTJO51ZBc6ihxkhj1ICNiuIBzvfBP
mHbkN5j9A37XjkMLRqfn+eVFujKDfySeZdI4MTbFNh8olHZ6J6qeHRzREzKHssRw
xlwbYk0wH1AyLrvYk8PQrWoqSkf2EbCMl83GMmqRuuxMdKt9E4GeC3CSu/FanWNq
Ea9TDPz4IsJFH2wiKQRvvNlpJjggMJZfP1aSjXuEvjKH4hmC41hJa39iZggbl/CL
`protect END_PROTECTED
