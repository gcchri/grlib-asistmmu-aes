`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u/tW81NK+8bo7ouGcHOLhsO9LtSDHW4UKpMl1EtsttUZ/nR1akB6TJgSBrURHc7e
VpC6I1Fnlwf2udJf+Bu0ClfNY+drmn4m5aVTbKCqRQmfrApY+MqTZMvpJVY4ZOVU
N1hdwRk+Vlu86eX7Sg9LiJdLCRzeq5GaP2xzxVANA4+SUMbhMVsOpOOYGgfN09ar
yVmkk3dShRV2heETspbUB8L69UHb3w/ReA9eQ3DDqL0RqfSvbpptFklT+vxGFoZE
O6PXcHheknL/Yj6R9570r7dHqKeBMSodG+rZ3yRK4xZnDdytl8zZ4shMYQNIe6gE
Rxg0bZ5dE+m5pb6TVP3tvj+lHuRZL4j78g3CYsjNjNBFMJPiLH/rdaiyoo9z3E5b
uwUN79DdhLFxfqrTs0VHxnhbNosXssCeTIpaFZEJWMv09vlH1ItqGE6tNj6b1XIm
DVjRaFR8HUVbwdMMFEK39Q8utJTFPRpiMwKuNjWYu9Czdqtxn8Imm7u/QLZgOjbM
CN63TJm3z5t4e11gEiopCeJuG562VaIo6clhsvJYUSlzYu3w96nVYf6xJG4TjVcw
T7nG/PipMJGRqdqVX6rffYthAIkqTjqsnPUGq8KtL52sc1wxhzoptPj3E8tIegUP
p/0qNSaEnBUtaVKc8udIjg==
`protect END_PROTECTED
