`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kP5cfSWcM3r4XXVo3fSHG2B/Jh109iR6909J8phtcJ+NCzgI26qSdf/up4pkGCmG
cYMz25XkqfL9SNdw9ivWETu/LAb8FTw4liJOnQ/1s/nPWRJwH/YWoGb68Z6GmE2c
vTplqIyHAHUR0L6IkSEjLnHtZZZbQObA2K1MORICCy90gVw0gHsTxko78suMUiCK
0Y0ZUBLrBLZuVSrn/4hagID/Zc2GEMZsVQ/GXPvBpzx5ja+8zb/EyKykphDRhf/R
4zpsYRApP86N8Iix/7pTX8OxhtY9x8PK/gmH7Ve4X6AY9BACNogLIxLy039Uyt1A
bhmgD/mDy59cp1ho6rLJ7jD5Hx/N/CpPx2t+Kyqjjo75uZbcznrCAHLICLxJyWRA
wSRJ4YoCkgQYNZkwEZSJkSLqUAlFGaz4Dq/v9o04jdk=
`protect END_PROTECTED
