`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dU1TW6gY4lBJ0XgTEAMRukOEmkShjb/XOPn5hn1UzpvcZel4pVDfbx4fQf3EZwVw
hV16RO1Eq6DsiX4YL8U39Dezs+U9TT6hYWEbKM6vZzz0C189DPr3GbzHhXEbVPiR
UsOn4jxp77HhCZLbSqdwuAcyCPJf/HidYzex2CRhH+w7j+J8P3mwH37ES9VZ02i1
IknRRoox+cXgVULc6hg38D3Vgg6SaQ2nW5Mm2PveYhVqHBHLiHaN7fmrCewf/WCr
kb97wC6aEHKjPpCGM0YeezOGNy44nrHPvxZE61Jfo4Xbb11PHdO2WFAoj4+Laz/p
/TnVV1dQW2nwB6p93nwpvQuQiGBeb2+iPjROZX1p8tEpYm37dmswe1kIvALpRMzC
w8U7pRFZ64RwhZp2GLp5fguve6bNslUo+qFQ/39xMlM1faljCn0YaSSIsimdrjfK
`protect END_PROTECTED
