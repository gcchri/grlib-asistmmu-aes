`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wQtLYXwUDyrGm3zBQVn5R4S1InpBsmdyNKyKpd62R4maXTmwFSpl9F6lL/PwaER9
OcW6+RwncUxtF9CBIanTpZxNpCeqwCIBPWODgueJIO/p4oFLDtcL6OYp4UrNN113
35/7Rb8/wdWk2Zp7d5EmMZXSKi4YOM+iIhqJYtKpgl+LaoZ1eL9PuliHZgOh90Bu
Lx3YuaCTm3WF7MKi4ZEE3BmIcUEMmj3/pGUJJrscCDhL2uqMBkG5pBOjb/MZUVGc
lImD29/hYeFImKFqJDpJwncu9NmMUR0OlCHgxscAfQTrPteQXXzT0IIPQ7Cbr+eJ
L5e7N0/ksSGoxUIpElru6Ev1WNjeyHXV8oWmzeP+gDohACdPLyprAI++zXSKmO0o
TEJIf8jgpOH3DG00qRCYAWKf31nmg2YJ+z0VroD8xCn64X6NYT1gBsKC7+UwMcmY
+l5ZKnont3eOwbZ4U8S4pvxd9kXzW/C8z4enuMM1/wPmS4kXyPqjeC8ewID3p54B
THbgjca/7/Qt+tGiex+iTsgJ9/m81Txs7FFhwhVhsmn7IkoC5nt7k5/nQGMRMods
+drsONHeaTqsAoFoBVXkEpTN3HJ5UnXXId3H2DnA0Os=
`protect END_PROTECTED
