`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E6cmG5XRx+M3eRWQ2xLhcMkS2ZzS0SmDTwZz7H9eohD9D0pPfOjHXEnhjLT7pIiO
s9fB0CRIY7v9op9anNfj0w9JBSbnMyGgaA/PgNa0Z5ojRKkI+ywsK1vQT5x2HbWN
lzeaiJ9a29wLu9r7hWAfORv9ZlG+oIrz+Rq4WA4myaOxoi2Sli9cu1vEHD18Zbbl
PQ1jEh98+gnwpaT6Y3DyWONXiUhOPvaQF3rdJDxjQfXWxDPddpQ8EBZBYGqoVV8X
xrty9yTwlR4ZyzC7p2hGlu7ugHaCR6nRI4tURrauIf1KbWb9i6bdUR7lWPnXlxCF
WFYRisI4LPlcUs+3QZhwn1Jd0adxmOSpw4ki74WwVYUBzsIy5pYC3dwfIgVAvb3M
BIw/jYLhvDcQTJPdukDtmIqiMyCZKsFxff30iSRgXhlYbSOcTYWF9AOXpp9dPqmA
OI9evuLUIy7IFIXK7BhqFQSI/hQTrnCJWgIFJiZL91dbc0OkNgEt2u10XqI4V12P
DCQuZL9b3JzQlcs7gVb832CuXNjng+hTvZ4V3gt5Je4OGxvFLpzoob5EEWMvOLxa
ZK1psn9eBQfS66munzhBQeDMLjYw/mg+1IL9Nfk+23x0xm1a8SZcYgW8cEyO/yfS
euOWPXM2eYUlzK2o9047DLof2cM7WGYKvsJRTv2JjJuOFluV+RgNq4UstNI6KzJe
/DaVfXdJ9d2dvb2UYNXCNjoYP8W55ZeqdOznb4iHOSp/Sk4ipfqxYtNhi4DWZpzM
Xk5i+dt4HX4QZVG7X0ZzBKY7g+pxK3vSnbDAhHgEsLzRoSjDKHia8TkW8GWTQtsJ
gHAOBj9rksbQaWv7VXgtgigL5JvR/GzKpQVTHr6Jikg3NZwz9z7ihlfle/x5lYSx
NEmDDH4zABWYLtVbdW40GdhNxH4eWxRXRigeH7AokPIA9Dp3dR6N6F8fulTGgymK
Y91wCVhQfGtIEZrTPZ5Z8KMpXf9qZvg2iZZZS9XgSJ/A1KfvlcPATMAW0cmGq8sF
CV0nGhHAYojvXKuepVqz2naQbcnGtFkATCzvAOOcTbhs3SjAdS4FsGbWH52PA6BZ
1NwzaDwK/4RXCG/40GkTv+OJ5ZZUeHPDyIn3tYR+/TZdTMNUg0X7SBYZcNSknKvn
rSmjMYBaQ9k36QOYddBTlI7OXon9m234DaaHsatzFfE=
`protect END_PROTECTED
