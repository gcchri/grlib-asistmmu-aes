`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9zdd/JbqQMF/DF0tpwDxXMmDbF05l8QRzyMSQk6Z50D1G0+RrP1NxkQJJKcfTXL0
sz214G9vipbupWqoN10+BHxInyW2XCChjbThHC37PC8ZCCUm3hJXHHS3qr0/Eyu4
xy2lBC0rcSKE++kJ12+zHc/sZVEh6HBPruOgWF5UFxQ00WIM4gUJ02we485P4nY1
+aLBIbNguY3lEY+Or3LUnREDicHrEUki1oChdFm7jen0C2vzUvtNbkHhfZOVozv9
rv4t5JfZX8K9e1F3bGVFUxWL02j4nLWgt/i0hZNGAEjJhjwD258J2j+iJN4LoCxe
zp/iomQEaAeKhI6VX141q/NhdUBhObWh2BXfjWGOdmA+ZehCyllfKbUMnCM8OmNX
W6CZRuQuHhr70AVKV4SKirfPkmBXZ76lpX4VUdo5JqPg4wbtgDAObVMcnHb+r2G6
vlc1MiOLW74AQLtScCeQtBbnylWvMeebf7hanaqySdaYJIOeYBHLn2FtRjoXhFD6
OYGn+A5nFGRbFkLhLiNGi3ki8eX5zdL6DjquXVdBlVO7x47XexJyAULlZAPIsNlQ
IIeTshxqCnqfIYt2y5yp+b5Uwdq9r4r8QMhjj/qePyrjNVt6BgxkRScfULk8Xz/b
7CcC0ilnxzHEnyLhKgkAsR8YratL2wOQ6S9N2N92/ch1ecsyhQZ5Xi9SPclbOH2+
`protect END_PROTECTED
