`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
58ldUQTZb0yZeyjNz8DgAdrHvRaM8/X1pkLr10j9wYprAwvikt43zABSWdhij4Z6
1IUlERltduAyWw3/yOkhUqc1F//WBbwY1D17Nkw8QGUNDAPtxI26McbxBeVTqc+6
qnbyLof9JmfmjmqPpNPZvBs3GxMcFeBCy9mske+LAOTpnmW9hrStENliAWRXMGlO
hBb9XV9eTxyRPOkvDHDpRakJLGrg7ZiCrzJB/abK9sfA4atWqtg3wzhCGpFXpMct
r20ZnzgdXiFno70NSikwVHP7Z/HDCdIMOWTPFbeHZrFS+yg699AvqsDTdF7Ymdea
WskKM7z6sGa4M118k1FO+QT3jt/SJQfszNvufXpmZPY5awIMulHSUmx0ReSaob2l
VdBJkfO7fmzl9XO34ngbhZSpng3fsuRBSp2mHazFM/Qcd857MxfQm0kl+DyulHNn
8AdbrkgeFIqh/Vn1a3Y6zsNKMOB+BcAJDMlL93VNvJjee4TgzknBxPED8im/EA79
tPd0grwCPM8nhXX8KXL32I7ILEuoBJrh8JLDOvfrAH8cSDstBTBTboFAuZrI8Cel
Gf+Rh5BfROUkcKKsvH9hOPbCG2bErR9vIbplKfkoMhDpzcMd6CSc4IwEf2FuFItO
9aWgLHWRDeC81gxNeZ+swwIzbaMzu+GveOmaQGFDssSkoS2ET7vxzIkMsA+y5T+Z
cJoT6T+yH/CO3brcn7L3n9fplFop3VwGzhrd3Rj1Z4zxFgb5+r1W2U+AIzMVa+GC
yd3vq+raixKYhkf1JcIaciAFIeDr3slgrRkk9OzWX984rIGFLbQJ9G9KC/iSvxBt
A5FhS+j099TUBOJ9+DuM1gzsz34gJ0gb1HTSnpCrak1RNkGI7+5+Zd11D/BfZ8vI
SVPCkV/Kb+ch8UTjHTp+umudpnM0RP1NDwph037JuqFTmZu5ZPxpXxsFOZ3wOa0q
CIJIIvPkWQBrNpvXIBzWJjPp2sovH2zP+phpNAL6IIoUf26go1k1y+2SM80NO5Ye
ARrQXoyjjDpoKAHiP/xnheXnEMo06P1BFhrKLFbjmj7FxoLeifZoV1s3tZmu1Fd2
WOpcMp4a/m1OT+aB+Mf91hjOTerUKzbwAWtyAmnvmSUCqPnFdmTiECSfx097OaZ0
eiDPEXIO+xJ0w+V7ku77HagTUKxjsEMbcS7xTD/4b47Zam9kr8/XXbhh7PBFRPRk
UZ7/61my1VVFa22sL1KmHHL9/mOOwHQf+dz0V7aDnxqQCHTOt3Ndgw8iT2LCDVbP
IdwFVN47I6w66GuN7EJeb0wUThQ2kz17krBOdL6qFe6/Q90B1V0QMcTY4iuy34+6
UYDYs5TzD++o84ElHJJEzTd3SDDNwkhNglzd5VJi0WBxfpztgFWh8tRYTxztVhYw
cbS5zLVQjQJYxMHqozpROZA/3S+XmVZHXIs9itu9s4jPn6+gjhOnfqd8SoAHgUjH
wAXofZOf9LhSewN5vVKFE035lSbOmbePabDqTJIrcnF/QpL+VmAhJRfTKXZs2MiL
bRxIWoWxK72NZkG756Q9B7gJtMsxiRMwV6aP+C3/Z0mN1jER5JR9eTkBFJvSsoHK
5CJNnbImXpnINZyyGj36uiSzBz+ZMXmsoHR4iH9iIKKYGPlwpszoZKSoexUaJGBg
BvFeu9GaqKOpbPi5MN6mltUY0Wh8N7FIkFMTpACjbQ/zfipZugdJkRfdO/5KTUii
oY7RF5rnPFJZQYHrIqVruU2/QqJ62uZwcxqIxlXPyJabIgl55owvjNwz2WqPw+pe
NjfibGJVQNHbdHtwBOf66KxAwjgmuWwwgDfAGQNXz8XknJHR4+Wjxq+Ng7o4GlV7
O5+eAixQbSpcxN2NdX0oYfQ9XCGriuAp4wykV8Jzyhf77o3G7/vIcqiFIxTdU20e
`protect END_PROTECTED
