`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sz+ugjgusuH8xd1mRGpaYyshMTwRPU0KkXquu6qS8uEmKtRwcNMpTa+uO+OIpTjH
rraHY2tzakF5Y076OVcAk5dgaWFjSHTtwRTzaleEjaIuJYj2KHV6XA+V2LP/Zvpi
hg9VREBj7bPXGDWNDPm/GH3rn5pGcL/9odmObw3k5SHh5ktpIzIpYq13mwX4FCci
Ccc5VPvOaudbbz2nKB8F4bsWyCV46KUzUamL4e75dgABhU5VEoM9z/0tugKXp2vp
DsT85Hdlnbe6lhUZxUrnriwGp3Q5F+q+/bh/yTTK+yM3kfnOc61u1H7sxz7Y/7/C
/Jz3B9CmJASorRiAJh32Y/flt1ACMd2DBiNSFA3dOE1xOJO4KrzjWvFcZQ9GW/Vk
WjaZu/jJKn2R6jjBRFmo2iWF0bTS2Mf/A3PZ+Yk/pROchzqAmbNc/swGz0TwP9cI
1MPXyw/Ycdo/6gYat9LkTpA56m5jG0+G1RdWPMEgzRggP2/uezA8ducD7MQCORVi
+JB7K6KHJl3sLInYWf3MrNeHxqd2/na/eKJ2Zxksne3/B8APN0TB1kOSv0KWMfDz
UHPB1HVqlM01qkDDjrdrsY7/01FPXazch4Bei9ZkuQ5fTokWucdUBuZOQUfXtVFK
jGjRUGfFpLBurzts9q62xiriV2Q7dHR7g395N/5umNoRdSLJRibkibiO1kFIFTVn
5HUJa9NAaS/NCA9Pp++ISp1x9sJRqQ8e0SZQ91J2XvAqF+0+kyGM9wQ0yt2kgPvr
K2AyZ3VhMP9Fl/z410om8t3UzNehD75Ll9W2KBkYibjsDPrg84uUE2oF4K528DUD
SoB0b0UDzxhxFRNMopa0qWg6mg388siN+e8lPj0O3COoC7hqr+/HGFnXo2/u0mrp
Af8ZWJrF7Ymwq9v1cmXI1Y+xy4IAnV0W9UfpFIeEfc8Y4fJvRWqKaMAmH2YTOv0S
/gO1/nC9Zt4Fm3kgQ3VBL6Nd3nYHSxoLg9nEL+3M5JELjm89xVXhsrbAbr2QSTlO
W/YPJz6iWsTikb7yvhcWLE22OJ4iZfE4f77//EQfxQlT0hf9LtlTmghKaZoYWikO
62J0w5eLND+bh2xrxBcOBKoIkcBYFhxljpjOv+pG48k3Djqrv9bAA4VXGkvXiv2n
ejESXecSZr+l7lMOyj+bQ6ym0yRrClYHyfva4pycqL/ezwLh0s3mX512tFmLjxbe
Aq4vdfQpeI9z8vAIdc3SL9fKXPgjBTWkEsdBXA3diepf3YmKP0/DlJCqFHbfue7q
fxm8FkqscbwNjG1EHGfgHWm2UI8yBem2/mm8Q7ezUKD62HmDmdFt8Ik5Ck9Vcuie
bkXMS58aoFBaV5Wtvpe7Uo9/sIY5bhNQWUdzrzEzTtK7OJUmMEjARBqv6PB4Z1I/
f9OlQUFgq6ocwHvWHBCDgW7FwCZewcFwdH4ZRZNV+s/il7lQ20TMYm1YD0+mJRJf
+b7IIU8I7cMCYTB8K8jcDUjGmuSKi5HJ7ORoQPmXmPxfRPDCdG3D6nIYsp8ZsNHl
qC9uf9TSRIwyerOQXpXvzUSZ7svrIes9ul+/SKvlI8WAnCaCoWyeIwL5aP4y5b/e
9OU3X+aSmAzYU1VuY5/nbT3R2LE4Riuuzb5QWek9gRG5Oezbiq/kt2JCf6mqRWas
BrSzmEY+2uSzJdJJBkFFdg3iPuuG31O4TTyVcf2+xRURTN40uRqBXqdtrLieJ4x1
OmGsK1oGrUUcNIl9w6BhgWoxGbiYO1f1YSuefgqrKlMve+qG9m/y01XUJRa50Bnw
h2qTFMPub+Mx9QbkMIYeA0lGaCjlcOmIOppM9Bt2ePBnBzfWaCHmcvy/LuWbL6Up
9R68dBXmgGOq29JcSU3IVneQYpdiaDWhzQYY7DEhtk2UJskOn85j1rhU27eve+34
B8f4Y7R+ctcTZsGXupGGq/WteR+mtK7PRcvYxlpoulok5nBYbiosAW0o4UFJQvl9
XHtNwfDJYSMDn/+KTw5oKdNoHcOwsoB/d9aspERkVWdwPM6+uTFtLRHjaCdB7NgI
nBsh3p8QOHnLAil+G0vW/Gv2BAAvP4iJmqEtC4kl8MLXbqf581cd2V3Ulb/MuC1b
K4Nmc/z1Rlhts/Zy5e8wHE7OyOWn88hW0nskczPnrrgn//fobfjyxaMvGtX74FA/
1MR2oWnX1Jwu7t/kiGE3yoQbeH0OLPvM9I852bM0NP+m4+S0RG4GgRQ0caFvsY5m
f6P3G1Kac1vhDb3ZS1e53HAGU3tkq+GfbL67u3nQSUF4ZII1GaSeHo2/W3tmiFqf
Xm2yAeIJeG0LcV5ICerfkd1/581G4vKKHd2/BKBQ0DXA0Uw2jB7mRrPzkC0+8Laz
WBcLsbxovob4SS6lIH1iAs/MeWAlRPaIJHxcwTqqP5ujtolK5OxSghsVQBJu6kc4
0Wvu/QNF5tKwinqXDaB5Gty46If+eQ9t1uJJNMCHNtRm7arNYwKWu0aGC6DzfyHi
RD/XEccVQT2f1O//9L2GR8+xHfKRqazqSs9PE8d0zl9qvsNCxr2LvLu56AEvUyUL
rY7RN4El5YWu7L0uEVU2wA2LfNM3LtBUITdgXklHwTkzMjprm5k7SEHxx2YMzw4I
tCqE+165JPkQpH9B1myaPVHMoaoYeyi+doyzaO6Jwwxy0CRpRU7BvVX9bBgk1yUG
7DR5CJW6n3D63zRuESXOYHzrOrLeGEMM7FcHnfct66/G4PdI+RyCDTlX16YfOobP
CYz66J0ILCPMQN/vqwTZZ84hNE7jR+DEpfNF+bpE6K4VCXHAwmjBYtMZs+k4FDsF
XuyDu/upAC8/eGAbd6mJXMg2aHhx1A8GQ4D7S52oBd/b4UKvd7MRaAGIWKgT8ACN
vEt2KfX2lzLaJ7LxV4XI007MgZ05bOOtb9bBVNhVQ0hXFU2jtL3u1hUzIO3qPOvI
5yETVFAY4ljV/xb2fnWW03Wf67rEbxCmjsF6779Wy8jTHlx2Nb+Ki880xGCTSI6q
bOUh2Je9ZTJM440rCFnF5e0PcBa8wv6NVlZZh+vI5HXYKNAjgfhNoSEkh0VNGlKj
Lv7EFtvSFRvLdRL0umq/mHjrHMo9bSbvf27EHRADDsr49GDEDrDyOjCy77MG402u
cimztOVxHFdP4TTzyCCKNgCU23y96ND4jPbrB6/j8mCIWnbOCizXEGCDxyA8ZyvB
tbnKbjEBY00jbspYmi5NLCUtL6bpTp6+pLkRjJxIlo5eegs2ufYGbekoMUj0qFpd
75O3HZo/JFKMb0VLlV62padhjg+TuCa+qRbMfoJnPj1614kagjvNzCTh/l1Q/4Tb
1DTC42yL1Nj5eH9Jl1D9BSktUeWO54fd8ZqM9bLHbYoLoswJHXp3N7PIVUoh0mmc
GbmwnjhPbojbgGd4+Wjmr8z89hgJlonksZfHPAL3t/VcoRpoeqxDOhZCwQkkNBoO
LsjcufZM6xotLEZDqdY3cNbI/YDnSJTedzsPWFX+4IR53V3ngO1BBPi4RlcIYGF9
ZYiEw3Hxfw87GgegPOnb1H8ggM54/rvmfmamM+WVRSO0PRCl1X6UU9wquCHpMpTO
54sKsiDCTGkzny7lIC+fdeigq2nvDwVk9JaQS9T+/RjeLgF2Y06s/mH5faQlBIDK
`protect END_PROTECTED
