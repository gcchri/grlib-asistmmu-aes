`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ubnwrjhkaQNR7h/VD6LKEJ1PKHjYs6mNmcKOLlu/J1QP21l4ubQMMjwDPAOvxDrD
LQGF3FSnsZ9Fv+nZLuxq5o+tzi2xBVhTqDbylqpAgR9mi5d4JSJ8PIzp0oxfefPN
Qv5BhfsVbQwvKGNqDpWLqUaKtPzSpoDSenzy4zSOnCUH9dgDnmYXuTlwBRfDjZWQ
zYh3BYBFiM70xW29YgviL123uqgpxaRHK8Y49tXYjfb5vo5o5MP/B6Ce3Li3Jpg2
HO9rPbeTnm4n3jRwvvjfN3bR1QpwoZ4CEHRZNTqurJ+lrv1bGdiblVujhm6yIAD8
luvVg7ICdrH2W09zjJ4N497dNhc6SbC5VrXxdf6W/f0j7re63ZfVzq398m2/00DC
Bth9oBT6is3gcTrOX8Hx7WCxrGZ3MydOpQHkmQBxGphhuisLWWmUGM1aEEdqIw1k
i/vgqujYFCqKmGU26mQTcyWwuarcuWLVEXeUhB9h5F3OFJJntjFRcqr0ZOBL+YQ7
3OjzuKs1gpjrmy96QYH+8tdbQkzqafPITHwaXzNACscVOirRgLSMi7SC3/4WmfTt
dJXB++3bEvNaQXlxHcmDku6s5dempaVMbzLVwsRhSSZ8w6ndmoAZgI5ZM9xkMNX/
QhH0kamjHG4aZSXWX8UmNJoqMT4yIBPMqKRwlhEmIJfoplfPzrSGon90p2K9DZVc
djicKXqp+X7e4oX0IAc6w1/rjknqF+9Kyt8X972dfracnjqgk1i8DxUc6Ik0qZfn
UKq+g01kEjWEAvhwlozJZSTBYmcGo94WJpj5DQdU0Ya1EWe21OX9jkqEfe8kH3q4
DLL1DFCIEMduhrNjJgXaKcsqMpNDh3LDAYvw3MdSGDNrWZ7WA4YxebsV3R8nlrMo
v9eKdm+eGPyuSDORv6zPOlu8UnJB6lNm/1cj7/mGpgLfPUyqf6d1RbEBCwqugLqS
fJazgG/g8MgAAVv18JQJiIuDXbiQ+8PWwWwGxi3ceBReswqlVbNMJNu+sm/4355N
1oNEMyonLxIXpD+KTz8gpHqGQYB/mVJyogOa7YkoYxu+GCQEnc8sJhodhcPCSrrJ
`protect END_PROTECTED
