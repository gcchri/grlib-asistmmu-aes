`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uu6wItrPPzKxtjH55IoQyzyznZhZb0Ef2o9H2MCR0YfzvsiWNJx6PepHi3s+VjwN
6CVIQ4VVaChqQd0I3zmOPsEkmi0R6SiakVolXaalrTwxzXjoTFE/wqRKKsSZcdyS
YoceRAfBMX96DZaLeBQ+muC1H6dcafZSv7o9DkAXp7Upqj3NA7GkuzexrSKHOwNa
eQgJ8PYD1y1oVsaAmVMZFI7DMGAe1MKo4CLDODhB3p35k/sgCcQhyW//AuT3nlln
OajBnSHIdFFi0G9Nu9FkCP7QyugVp+HLfbtG+wGg4ZLP0qcc0+eR8LFo49g3F/3D
+Mfn4SsZG0c6Ei6xPaACAythH/zxE6y0Y3O1rDA+v1La1O3EObQWqLPTLe/7xyIC
SijeQKKG5uH2Iuzmf73HnUKe8UaypfMBiNdDp29dD2vJhfvgKALzDDLICBxbrsG4
zq10E2XF1X4g2rL/k5mL/K9peuG62iYSoV36j1UfSv9FihQTYLCm1UUT3jxmhT2D
EkkdS08WlXrWsrj6tXfhDjbPmEOYru+Jc+y+yu8DJBYOt2bpm/d1zop+Cq0LbcfS
NNJr0vpfS94PyG0T1LYAdwWUyWn7npabr3jJ7eJbUajStL3S3fhSr83vyebZcfWK
WoKc+liJlIAxWQm6Id9lwZFwjuME/6jQYmMei5mK6Z3cQeT1X6tgqpVivLYor4WC
I/3kc/N5J8PKS2dGPFKeiteg2SqhQatY40nF5IZGc7jukmpgGHs8HPnQPRU1UiI8
YD9Xp+E8GUXnbWj1x6eK2cwKFICwJ9EyEGCdhkc+qizSqkhCPQyJ2HzNnJDoJ0xF
1VYEnaWoMpacwMpETBY8hSg2oU+60TteozMtyckZry3DBJp5nQWLWAQt3fC41WrD
wx/KUTh5PS7D/9pAaUkoI2k2Z+QL4WTSocJ7JnmRjxVAJm/Hg9fVjOBDM4a0VJmy
gSdGWJL/lIiOnYy5ktcoTmNqE2NAbiNHPzWdtNfvYmABfB8TZm1xYOZ0G6X+l5DW
V8pNzD0NNOMhTSCG19Dz7SfIgUKGCXlEnUN++VgwuHDMynweivC/ocKhcZ/sZFIs
4vAa5RQK7wlDHGweVaDIbGrmWKDVq/+Qrb7HWjELuSj2XpPpukDBzLTpHyPJSPMU
imfF5GBAr+ZhyDNJIlvGmVuAzoYkSzd4/+8nmWqg5VAmPIaezmmL8ltMBVtofh6f
YvjCNNS/L1A85zcUnZSCbMvGoOYXs81BbfFdmbRGuILS/3uLFjZE4cauAk/wG06M
IXCmY5l9SDwFlueFNSTAHusGL9HEI4+iG6KbZg6yjZQr6B4A7s5WSszCPpId9dT0
h1uaIzVyHyOq70J15ibbMvoqk9Iiw1hf9trQB1/OuvS9G8EI25ubE36XUTzf8Z5r
tMHO7tpaLcLXimQexXYlrhHMJhmrAmwH0ma/CRYfJfBbknq1UY2R7ryX2m2B8TKc
anupmI+JtNJs+4DC3ebjV2iSoz+Z573O8Yq1rdBuUG16szyjZKoTPaDDrhu112Lu
RF8KVKY+V6mOE0CFjAuct2gzQ/GezHgp9a9Pm0gL0uau1wx23eUA1q2FJMRDjDdv
zC1uolOm93r3n8DT0uepm2mCx2Cr+SLcYVJuOBartsLzjBLaOf1fkH7JADGClqDk
+lia+bequWWpwFaGzOisXIB1nSxS38MMcy32sOjkBgiYjO/sbpl355h166gPs67v
Cu1xRBzUfClpuaHBMnMonjo0RKfM7fHDRrBCj4h07SyccjAj+aIfZ30xIUUi2ebt
bAGIDI/gHRayMCg89iI3emckP+NJFUJBcGmnQjH3aHx3L5WqKCgOLyXQDOZFXIE+
ycNspRmvxKs+dCOBhwO8fnS+YEVfu+oE3vy7G0vq2/Jj/y66hyiTNlRHqIoS1qdY
xrFERf25+Ncf1z7HUGa9laBeoCzvo/HOEuKNNXb5UFg01bFbQVOade8xbtSMoYtq
SshJxGVqcgO11KSYEHZrORr0yw7o0QOe1bD4XmJDzTQ/HX7PpZBe24TPDnEWoPOK
tA3IxwmV7w3GnRhU1UMcHO/iQSm/wRc2Xf6r+zXekxvCxSpt1JROTXfV/HWHatN6
m9pvNZexrxG7AJyYKLs4ASsqeHHCT9XKSiLcOUHYVFsHlu68MJrviD4DPcfw2H6f
d0Z7tgpWGtChPJzp+SwBjWD7JStEYRMQRl/8/ubds86Oym940Td2oAPxCaVF+EtE
iO3gA57S0nJZGOKPhbpqBZqx+Su1+3Az/1NXtYW0aor0R61CM6TS25rjwEx1jSqn
feWRfCFoXqrJSB5B3FMS3M2R7spHLFX3JJgLhC1DPTgpVm/+mkLd/0rNXUEtxqT6
MLi4sZij1ugqXSL5ER+/8i9gGlwGWX3D8zmXMzCwh3nKwJg4BXijSmFM3utYv+ZR
zbp5TCiFwO9DlxGkh9FBGp6pvlfAjkpuNyuSdtvGhtXKWvaMhKFUECnnIQ2jd6rS
zTGJ/r0GeorornYzTGBxQk+4rv2gF/dzeY8wgwwqlatOzVXvHI6edFZjPA1W4oVB
OvgK59U+EZqIcBJyYLKaqp+so/rZo5gI/8MUuSAIPjAA0VnGKY99hN7o5A9MU6fz
+bBjLaKW7x4bjG+81CHn1HJGEGguibllupmYiNUcseKgjDB6S8u1q7HyX8YA9T/c
4LtOnPT96uqz4m32gE/vkIxQ8jYmXyfe0UeBvQbfqTZYOZraxw/PtNroy3ycqGC4
PzMINkgwdhPhZljolgIo+HiX8WLB5B1p/5GUKJU9bMgrJfzwY9KT8m5+JSHQU9+i
gK2zo2A2jBTeNuo6vQLKDYgx0K5l/Z0K+XETzwMdAZ5KBGHGzQ+ifp42qVfoz3WA
fFg2ADmIecA9xIba4qd/CKRjD/GK+/Yg1THuwObogdgT8AxF+q+uWmtdQ4RvgLVV
p7/+vxmhuAq3Oic3N+0tMGS3b+M51B95DJPnlMU9yHFhEu+9oeTeegZ2TSWX3eiE
r5lSbqW2K2scI1yWAZXWbFLYR11znoTwrsyxTKDj4xjHAmhoTOw8VyzBlqErx35G
3HJsQy0dQpwrRny+iAV3VSJJOpDGdw6dslAEP9z6sUi/+C2oAXvZHrpOGPDowPX2
LlDoUyYQ3QCwIVv/fRM20erXOgl27D4bmGuFEVnSPiNZxaj5YYJ3fu/xSMBdknk5
IbKdf8byJXtpjOCxDFZlv8lKes2ss1PXaq/rfayw13rWZ80cfs7Xp21gQRwI5mr8
uBUE0qKWG5inWvSpM0wTG600onGFozWBUfLrSxifXErMO8Rte/mhkoke0wAUsLVI
EoC4zgLxNK76w5v15ojTytcWBv0CiSBWLvwwyZCmjbkI52AFCZXkWawvPi6N2Mel
7Hcq1mkrDZTF3wKZbR40wei2hOs0+942UYtIGHsCIYxEjRE0NZM3+WqUnZBqKiDq
/oHSqWcfre9WW6Zqm1wApn8Qyl/JRAf67UGXahMNpTmOUzOJOjJzuBhJFOobe8tQ
5WMTyTJXFQL4ohaZeYOscwmlG+Y1Xxq5+0dU2PDyLCOYDX60KAqMJc/wO9a0zrDQ
RCmdFORQhFQFr+To8rHT6umBE3/mxv+yvF7Ih4nEht2cmUdDKLEQp9r2i/AKqKUL
r1AlQY0ZSfci4nta5syNcIK9uAQFeaSPqjnAtpqARIUGHLYa1OgBLI1kkZ8SeWVr
Zv6K9h4ZdbCmpKkMj+A7fV+jksgGiraXh7B7FWN3UpFYoUz4DYOPTroNChxBjtm6
xwDaY7rXerm4RCls84EGS9FVLcxvMitVysKbRgt/4A8/5yEGzlMRLR0zY/ptaWAD
sj1hr/2JrwwZe2YJbxFm3MVMlkqnX7Ha8GlATLv6ST5FQUPIqzXDb2onoTQ544fi
g6sQR2xu84OSMLd6iclCg97TVMFG/1AFv2COxcnE7NbeL52SOjli5UrBu/vGdKlJ
1+KF/s4f5lMk7T0CRx4NtUsgVYurJkGMLPeEpUA3xBPDK14NfqsanFsnMohU/GY9
o+ug6aX00qvqbv63Zckt9+eDnxcmB2j9QbFUM1jvkw49Djea5Z1e+ZBikxl6AzGY
Ygj/qDl87eV+NY0emCL1mDvJSCXDCr+a/BiHu2zrc8HhJ1kh/Ci7j2C38xgb/com
9kS9NVnlcpHPBAoF3z5kyvS/UDFHpxq5c0wU7/Iz/5R512vbDAEJPnHb5LNKdGsS
zefzOR3p0hLN9g80fBOSnHn/H161ZjR5krdo9nTRjaxz2UhujVlAvc4FVkxc5c52
Y2SJC2mTHIfCPrmGPxmR+T+4+9VeRFOToH+ilpUGKccGqq/J5HLHxjsCD7/5WVJL
tXOqYcYCSX9ZrpL0SUmiVRY5qZwyDAqoffkyUJuRDKq/VJZTseO4AD8g4z76jZ9+
o0HNeyErwwru9wKvDAVMcRIGQak1taXC2geNSueUXsI2JN0d4oAv7v7sVlcD6D0x
wyP5H+CgWd5LJ+BNX/OF5RAe5dFV8RwLktTRduMB9xuB6VoTocbyf/KAIsdrRqSM
ZnCJ3/E8RAuExFOgzfG3iyJNbydYCm7UAbDCrttmQYVHJpSwRcoLgyku8yp+EOAl
rGErVxcBEut6NRKhU28Y1quI0+5k5sPMWSe8f7zljJ8cHRn38fEHdJmwJ+RlsdoM
3dmZyY+7ojZ62gv+5baXZVR87fZrpo3AzFCPzEWGI6wf+4sW5AANZrWiBJiC5E1c
n90nIo1sNED/rX5+5JVKDl6/qqOX1z4iSve1KT2lCPXE127eN6yGlLH3wBP8o/rf
XRPvawdhVJ5LRGKr64Qgb2IkQ5se7XFFFox92rgvL3P1jmWsOSdqRxR50GckFOfw
toYon7F05PQM0gFqR14m7MHUYSmktUCOIOBxAVWXMUM9LzKWgiv4rmtnUJC1cOVW
DxPgQ2AQnMzqFCtB8yGs57rA+3NNwdfS4qtaLatK5oFBtTHlpfV+rcQ8Uu/sAuBH
7G+mIuuTY0XH65ZHoTUkjzmyvQsqubOiUyX6IeLPT3Q0+8FJwQPix9GOPP3ir4TJ
JYm17dsp0p+Xu3RTxuXlHJRl7dBJ/uugcgzBYwgugKdDanHB7cXjQb+iLY9ic0I5
PoNGOCFoJnINWQpyijZ4yBM93lufJklalovvFhq+uAB1IFPtZbMvcMf8ZaSYmOrP
H/WqyOjBwaX167iYWiz7JzdL/MP+CNOg5NFNhzH9s39ANj8HcC/EZ+7rFZCnRtjA
llDe9llyok9pg7GRQl14pLoZmnu7ChtK1Tbdz5uXvxuHT9rjThrwylVe6kpOC5jG
ouUXQVtAvlTL4Lx90zJK8Q0lVC7cMJ3y9hdOTqMZwm0PvJSeUEa6NRVQyyvJWmjC
uJ5CnNa3PTnPtjQucyTzWjgFmVxYmxdw882QJPJFq03Wfdoja29eyeRxnqrdBrYv
jpqBY1/mS41Aq8TjnzKmxgXsMqKbCL8U8dJPOCEcwGzQ42jXzQ80GUQ6Te4lRLt8
R3aKtxMP7XgRfD9yBdCDTElD3qmq1hnJnf0jwgi+bDzEDn7LdyNGpPCkf/SbYB67
Lr6ahjvH3Fae1u6r4iDXl9PGKg90FyGuhW9/uTOOth/t4earw1Hg7Z1kxce3gUph
I3BN8EBDUb4yM7P3eswgJaeo3WBLbP/zF3eiB8CPTtj+h2EZWBhXx9t5+kTLK875
g6Qsz+5ZGfmqMDgm9yf6Ix8GU50oBRSSQyQ1AyuC4Pkjj4HMzWZDgQYd3GFA8hlz
03YcLp3VDwngXlH2ZClqmWZXVQ5ornf232ryFpuGfYNcFRsEWp1zpOsbuY613bW0
sz9PgByBQZtSujOLQ+LE/+h8lV3P4fBxeoct9bQQOQ4bpQJDP8wKfZg9T+hp5W/H
jUTVKcjNUFZJ7M0eI8pby93fTbp/RU97xYI6V7IB+vn2QcyontFzYDInb7fyXfd8
LUSDwQB6NP8Iks0oRWEmrNmL+1+DE8/VSDsCzSrCdM3uOROWaXUcKlWQMnkKzbSs
Qw7YBsRe1sYk8WsT34JWpXgzVE6LDSMaPiVLeyeRmo2Z9ffMFjRvKva/aakGbcuU
Ko7XxV+iVgx+proXsUs5qiDseCR2YJ5eoubfJxJX5NKlSnetuT4L9C6jh0KIeMcO
hjmERJesjcFGVuQxt/ArlqFpaNBWdEIJCOAO1fhJNwayk6DdWhZIOFINuGiyEK1g
lOM1/uyYH7SprTC+PnDBaJ8DLh4NJ3oJvBf5K8UIW9G1zHK3SHbr7Kn56D26NNg4
7eOEFId6EvbcKnDo28TbsrwF+B959E8lsWZH3/aVHa89ORahbTSrLbjjcJF476kO
bV4Bvu21eUY8f496ZqU1RpuCoZPVPBL4FIOrRVLbMm8VpNacK6rSCOpOtEbIIznh
smKcgfFx4JvwdnbBvW1He87mSy7vEWHLuN1a1GnHdUm5rIdZJtnudq4vxR6eXAYV
kZ1m5LzwBijXwywwh+31itRRWNSeuScKVjAUcXZF3mXp5dw0iNgHMYIKRtPfq9Qf
0gjymZ2eeNAv6ha0JLilSO+yp56NqqWxv6Ah/wBGgAbNYBMAqidufzUOyzcFtu5Z
qLvKxfSN6B24HYp4mdcS9sFKtNUdKFDUNtukrdASjTy0H5BYlaJwRVljTz+JE+Nb
iZvsiSovX4zlJQbF+BBGv+sr26+Z9XXHKe+9kpMSZnMfiusPc89WynyDZrJJhCsg
F8rCACGbWSe2Ap368H28A7Xylv//YFz2NVkgIeHkr5wXI7Yb3o2/O+WHUpufWFTI
q2aLpsOWeJuZCuP3eCtLLi/r6uU7Co2WRX0ndkNlML4eJrhV4QV5den45bpJNOYh
wWc2VHexKRHrhei7xv7oGSPHmMRwSMt7JbaapmU1/bI7MxgzIHZwX7SjyG9TO+Hj
Xsytwsv+hOyGT7FBj96e6c8FAPYSHC11FNF+8b+Y/nlOfsWLmY2b7F2Ullf9Ca1a
8LmjiqxmehMR7IRYZUcSwlXfdmvnKc5s5D7K/zieNlX5sxCAj/A4Kj1GhDUaZsgg
8EjjcgFF7P6hyC+4pHmb0n1qc+IVMje5edtX/qHLVaL+jFocKiJDM3HMdM/aZDS8
tBFnnDxgRZzj3VMd1++FEunJWdLn2z98gFLqjFyIrPbqLbMuwYi678hf+Frph4aC
m55X0CuApVhEseGLrX3IrMM5cTLu30xEJjgQG1+jNVmBc75ajNU1z+gWz7Pke39f
0ioLsw+ZLKJ+/BWsRYc+RG7Ie5g7l5fI1uPkPH5D7nJu4lmIh1ep+u8C3HAtD9Om
5839k7poDArfbRN5ThmGRSljFrvivRF7puxYWbNkeck0y2mJr2A5A+MD8EYu6RZP
kJn4QHEC3wlPGp1YuDOUjqR5BU3Wqsx+rzmwWEJtC1Z24wYu2VYvqpize993qytZ
w+ajBPAr5bumAXEjTZ4Vek2sD5l4d2DxCaJvpDYpq8MPEWbPc/9AK96V7cSLGSNT
BNX8ygHHCA5Q0EwaCzzkRKTC+SISd87PduEq1lz7oawGLmK4708zX+rVkO7tH9OS
NRuC3Iu5HP2c4Wo+e8rESc7ZkWlSm0zWu62laDOG+A5grajSgOy0vQ3hynOaVRGX
oY5GJSAWoFrh7ESlr/5yYk32bG5oY+fXW6VJyIWbDAjLNZpE7aHn8KRljGJM3ETQ
yPokBk4MMb4UfGj6JUGmHDpjFo0I1dzyXQCBQcasSTwDNhEZz8q8NdNr4VuDk+QZ
W1Sw3Vx+q0DAul/owrMcojm2W8NRKM3mz/KirNCBFtSJ7W1B3loPGCUItTX4uZtp
1wwUsP9ZyXH5MlCxHs3ejSA6mRG0uSdr4Ma9s9ScoPHPNBH9Kin3n5NSNOKHcVno
5V7yOIZ/3cP7a87bnZzYRiR0SJhuIuhauXj0m8qu4M687oOTLhz6Deb18vhYd+2y
oAxk6VQpASki5SuMnXloF1anfuk2lI5TrwGkiFr+ijh0eVDd0QA+pQ2JmlMndxRD
a9Bu3J2v8cswDO0XnXDvGt9gHrOibmwOfccMsTmWlg0juQqGh1xb18a3KjGYh7vz
ZCe8NhAQEFVfL1fO7HTGX+7wfBJDH9sVe6kjRM9j4F/P9Rea804LlHWROHq2reBI
TEJIsPJUmcM0j/8qCIZuX7rpbhrkY0BC+8TLIcT6kExWl1C/c/kyBQ/XRtrAWBOq
/EQBBou2pH6Z2I8/RpCYneCmjTvUgc73J7ECtla6mI/o3hsQh5D3mi3CKIdpIGDR
1sqAuqABnUjk1nJFh3vLjdGn/kdslQL2+iCwoUeXYdNtcxd+BI8HsaucyTJpOTc+
InPs8y1vjcHLL/hGkdhUoGLXReUnd4V/kudXEOlHwaFTFNc0+pSaH2cqjFSmTr4r
1NfkIEP1/hdE4A1TJ6gJZwtRjlWaiFoK2ELWfGJmXlhD2Py+++6OcyeoWiDlOKhf
dbnv/vJg1zEjvkwL//P4YGeNrykDZDH9/+Z2RSpt1e/j79XtJ8M4j8H9oREPduk7
VIW6PJPfnmx+9YFI3nGr25+PJuoraNXKPX/qvsyTHACBo7JrSQW5q0IPfclOJbf8
OTitrnJ/7ZBmFZ8YS4iCIcFr8Yuv8Nc9zXgNivi9AbsOz6CNy74ISchRtDaqo3HD
XHFnvVjGkzMbtyivQzb1JDcV0Oo3IdCdKjBdkZbqqIkcXFhFyf+4v7D34nWSBqb/
jjJfiQQ1axNkdjRbxlLumCLG5zTiepV9TFEmUjl+IrYbh0dYAKm1zhdjydHP/ZOV
2lyZHRtiroiqeEKkDa0Y0vWwl0Ofd6Q8rGNZAlKRGJ00+Wal6tH2d7kVSk+QHsr5
sGIoitSzWNfVkxkmqzJhP/RTd8poDH3p+DKG+kEbrWSpnLdY+3P4DVsUPugsUc/K
oDFAJGm6ENp/dsCjexl4hBt5t7e1WczGFjBkY43ZZ2wBq48iJXGOb18kESyqHM2b
C9U6dDtApwEOI6eE0FK4im1xxZ2le64yUGojDdQ+XMzYKpvfVoTLpMAddvN38Nzx
2EtVXP3clVqxhZsnA93qd4di/+Ek/CDM0p/yev0IdEsidcbCumi84mxYy+C+f0P/
FRaNlRf6MKpqD+o2F9gUVdJ4cz1r7TsF+5yHreq6/RKts0bghjWan6MH/7QpIj/8
CZoWBgoW4VL4RMjfWn5qdPLQDoeJ5exgNPM7kwl75l1R5W7DOYShtVfqkGzmlLne
mJQTLK3Qfxqd8eNe+RClTvwaQp7ZxmrzdxwAIUw/d6vSXkJr8CF0gkqZGLZFdewn
Zz4fg+5X6d5y43h3OmgMAkef9YQsl0sefEJWl3ZZxEgiEJWA3M9sADThtmdz9Vx+
rfohimVAiYIlUDZe1OBQz3ra61fUmj7Y/fddvg80gM+pUrSZSHOjXaBlXm+q2tz0
hN5nPeUFhatYqShPMBlssS1/wNDG++TprynXgs6cEESBHD3QC/dLE785wpAyRyAn
vFw05DYfb6ulTFSJdH14jrIil8dNRUxit9wtgEW7rzDbC1ltS/on7cCTXadzlcJ3
ONtLXkvLE/+rM8NqSJblhhKgFfZuTjgEkoDYkFg0o0CuejFARUGoJs9NNXEn37Xc
IvYmADCW/VCAAAYUcqYG8XPN3BWbdEuH+frvbyyHq6eelRNq7tI7UMmZBEbsAjdB
WlYh3srtW2pTLA17id7RFCYdm4RmHLBXBt7Ej1LXLRUDDTb8XOK6U2Kmd6ZDGEYh
MrabWzUXqef+DruZ88p+hxkUIIUaaxDlb1C/JDenEiwH3Kx8ST6kg0Srx+cCR3gv
D7Qzb/H7TQFjVibvGPvALN6MQRSWS1HREcegZc01AIqq7MZlAdWqthG0cjFx8+c7
fv5LWGtiURYXXybLlvpAM4t7RH0r2e/NKg+/8hD1gA17qYpVXS4Z/f15D3w+OOwE
56zF8iHbLilugDTrYJiGwwr4N/2fql0kBN9a5DOLTo163cen7yn++laBR6ya1s5i
aXjkkF2biaxCihmeGE5a8pXUCAOovNaNK5RQUry2wioKgcqG5AVmn8hraADs6LoD
0TCQsH1qPQEmuT5BqNvDsCDoHvrtlSSuXzH95HXppuAy9dYRxHsbSEnJhePDCr+T
fdKfu38+GFscQP+jZv3xRdc52NxUSPgxPnWqVbdQyssnlogoHUhhJMATLBrCq4wh
cLyb5MYvUCRXc8rQ96VOav5bhBIoQw+ylDrbnTP1V2y06fHVMF9buxkKw1PhAN6Z
1zq4WroGo3Tnw2kUXt+IJ7PDGXuXUfmNcQN2syc8T7A+I8fd/hn57MK8JK+XrGEb
HY1NoEJ3Mt6q8OEw4k5lnYczV3sOLxGvqETZka4AfRA+C1jI/kJxPh7xHPXXJR5c
dEls+8jkgHgyHNX0oDv9E4HzBqAMgegkyFWIMFQUFS8vz+ZBM9In9RP8r3a7QDTP
6+UzhZeb0KvJ4D2ibiRDlZxN9Sg4bBGvoEaNoa2pEG5lC4CCqIDrKFwpDuDXyC5z
NFRENY9ImX+tKgDehX9jOqRcUoGPM0BCp6CVrRGxfxz5w/NbRU02gCt+/pzhif1g
lR5ltxjtLzn0sKyrzqU1VZFOApuH23XVXO07GK4KksUCGfWrtfP3n/N+yVBiKaKW
D2qN/xn6g0qHK0CjQcqz+SL+04YnsvnG0sBpGd9WD6yn/d/ZQ4LgjNhqi/pDXJzP
eZI+QTp1QMrYAtPwHEinX27ZPszlIEbaTe5q7CSbOWzjME8OS2ZaDqyMqYBpNoUR
vmo3p7/LuYnkRy+S1Qum+qWWtOw7mvETaIAdCtm2ZhZTurm3pJ++uqJY870aqj0i
GGD+vQn4VReU3B9qo0fj3DsP+9BYcUgU9+S6qpPUJcS2QN+XJ9K7vmuYCZx5MnmW
4LpKBniekmcbvw+TI5tgDIaIOnc3Et/sA6JfLdjnbSRo2VD/M78wIvk2yMFhxnnn
Ue0OhImEnllxqZKcTJceW1ZkjxLns3UbztxBJSm7HiW4AOy/L0D09rEMEPBDsFdW
C4Vlre3dJEVsb2ZTodrCRyvLCgupdZh+UlLwU+Q62s76ZEYMFO48hi1KgWzF6+gW
x2H3nhBp40c7/dAHODDn0mYKnJmMV/xFeinmiY+dXfOSgrwzwOvTvD2s+f9JqS+W
qoe1op65KsnpBFbu2IV+/PVg4UUDBdgEBVTTd+mkR2p9rTo7QOKEas9vyiwRMW0+
gQUtObjY1U/IRTHGsY56NJUB/kOaBFWAZcQMEmR6PeEwxFbVZI6boJDFBqdMuiC2
ublLHq+Oue7IbnPCILJFzw+xgWwxJHg7DkJtDePuUDpK+gW0PZWH5pH5aOx/rqpC
s/CuIVV5YoAeP4Zy9ymsT2Hw/tYDQeBUTe2dvpypsLvwBNEHmD2FhKWpZvA0tS2+
WAjcK4nwTxmw6JzoNg54BSQ94e7HIbLWcSTYJwK82psWVwoSTtf9Ver5XtrB9det
8M+EpGNolVvcNvjArwsqdVjiIzhXbRYIGbopABvO6YVBC6jlaHwh/7Z+oo3wd/86
SdavfzMGXjcQHk9dCX5dQgx2xsC9c1Rv46cyWW2bN4GNPs/ssxmQ/l7UGT1I9l2j
u6SdjfyyGeYVF9p6X1ygAIguUmBZK5dQ32kzEsuHDhWyNblBMxVbzSynDecxsXEZ
PWgXNaXNfxeHpBjyIfpUjM4RsZUpOPWCQtihht5TZnNXtY2uZkb2F6scbTauAaM+
zlH94I30KODoffyGH04MUCz8YGwJak/NEqbq/8JNVEJVGunwU0poUs/VCW3BoJ9I
6ZmzebtFBeCmsmn1L6Bzv6L4UPA/aOgXhhmIovqX8Fbhvrj8DWi+v0CtUCGBwcXQ
wQA+yey52P7XOYBodEJg9M6hoZCp3T1cSZiA56/mQ2u/l5jgGH2OthFoMmBqAoct
MUwJs2/rXUXv1mGEhbelbTY3w1p46Js3g+J+qRi8HVxZT2sinrpEujNFe/g+6r40
Dt88wJuG9IpguuzB/RD92/QZQCNEv1OLGLRQzlakERA2uJCZ3XTUf0lFWKt3TuXD
QekcDl0ha5m2s5Ag13B49cTjyK58uVibzF0UkDhYEQdExobYoYHQSAJ6wrpAK7W4
ociISjnYmbjlIeBewwfrCUXDGXN8yAeEgdZHnOM8pQti0714csrl58cnsk6qU35+
cSLta/ZTH6Rtxwhiu4fClFDVZE89IJAXr/kDHzGmf8IbByY3weRHlJorBj8wvKA+
K0hwT/MB0Xhb3Hu0Cpwb6I8CTFTfqv8TvSEk1JnslhUyHu80PCjqi6Y0jnWxB4k/
qdcqIlbGpXs7JnaqQr5Fg0T0t7OfwBt4BEvcjXDEUdU7i9ub3IgyXZQR4fUUVuwZ
irdHhwL67AWBF1iKfjFu9uAEbfYC3rKNlYEST/PaaIuJ+1U1QXOmzt2f6k442L6N
RQdQDJLOQgQEY2YuPcp5jyZVdi0PODzFf/ceXeEbixpHPIv2LUw3GcHj3eEBfGQm
MxQ6eJ3E2+uexIQEAKTLVeJNXCDgiqnef57bVba/XZ8a7UMiZa05Iv8D1MzJ4Qvn
H9RgszUHYCyWIt06xo7znrqWGV9UgF3gyttb3sJNh97eDnhPEgP2MblGDgDuVlN+
gycaaB8b8HT/DkvOdo0VJK58cmvESVPZubEEl3JbDtKI3OpCW+N8TkNh3fTP7Q14
EXIPddZ+a6IL3G/LV3glD/4idVyQtWGSVxMpgdoYtH11kPYwt5Tdebz6Mq21VVoR
xOepNNZLbLlQtrTe8/Hs9X0hFXzdiOqv6a16hbgKO1WQI2jqwUQjf+RLEG7Fg2Fk
PNB/NPhBUmBw8tGyfD6EjLNcuG2ATYfDDCHr+EeL56tevVm1geZq0/XZ717josnt
/3CRY7yUy6qbX4CquINN/f+35BZQvWfGnNFkOe7lO9RBt3Q0DgWFd59aDSu/UfUg
MPQ2yxkPCi1Txq82cfZ8eqKnTro6Y/euBDGZ6Yoe+qAIn3PND4cRzNB3tE8ZpSrz
GlFSl1B8L9S5esXAxTMqjtSjoF9fqJB2cO6nvNdI8/WpsdttuvidK0fW1MRodoBf
d21vPgMZ/bSpold6aAhlg/3g98YcPUm7FxPUtaQu8bj2LAKlq47CDciN0RRKDurK
PKHtBHSQMDbQITfs5CJ3o3JMslWhD5KugZ2x0rMjnMsZlD99DjippTaAqMi8TfoU
SdwnHJnZecmGdrefvRiOYiDn4UfVLduBMoAVL945BmvZVvwoKSyp9VQp0vp0EyYX
H+S3mXhuxr/tn77fT4Jc5mmN8aF3g4tR7XaD2eaNMkNRTMpghrH0vODI4xPCsaAL
GyDe0zLq45RyWF8+Lz824eY3vBXKM7ZIXKG8CWkZqL4nQJC6JzTMjs+0WZo0JQnB
dNJnqvJ6XHPF7EiDSr9r929auUtYz57HxnQY3DOKeGSz+LQ8x9yKejg07R6JZ8Xi
qsxp9SRJ0awqgyURi1CC5y/cdqOBJ8MiQOm7AkcWsZSF2fKmbDXEHIFeOR+Hi2Au
InMfEkuM9VhPRwlXcEHU0IKSQ676JoFCl4R9Qiq2hz05LmCavJcmzOVh/6ixpcVe
n7SDVml073C6G8SGAzgTPvDE1I9rHcLMVpRT27g1Svg1WCinsTCMoVQhZOKIwaRt
kzLHTTmN7XVGPi7cK8rnjG75rGiPUDskI5/Qg8Usv4L1wUO2Oj7dd+IaS5IYp6FR
MV1dUjuHO7If7+OisbDi8b0wmXhEjpsZdkujwIZ/RCeMt7UilHui+Nw6V/g/QNEq
Pj4HRlE+UgoCArNtoEROixNgqY6w4f0JygbjLPK2DuKYufZdBEcRlUESuEwEjD2Q
vME9rnih67MkIMLpyTWjhy6h9O9nXE0jBlzjgGM3y21+ds2vlrUpwEo7vixvLDrR
uwlGpOblbCtsMAJtFT95CKawOQLl4foqE4wESGyo0lorsmIsLaPtu1ZEdSp7M3G6
ZFnWvYH/C8M4nyqO827XQfCME4WTggjPhYdmaKASr9Xwko7Mts3DF4RWehgtHtAA
utD0gkFHB/CYzpLbL3c8ONtJIRTeY7Ib1vxl2V9NN49uQjxKkc7RwQw6bV0fr84j
S9tE71Zgf6AuiMq/TXnSLsHMruN/zgPT766MSFr7GckQ1JcqiOv8XZen5TGRFCMM
L9l/IeS0GtBpfJCYsXGfidI5jRo6qr47mH4gnweXxX1SdrEy2yCHPeCkLpSoIw0t
Mre39bN6KgUqc8ZqAY5gyd3sQ6EfYnyYLn8Xugy0gr8xJyCm/RobBDmpGyWn2IPr
rzhuz717S/hbVKM4k3/GR3afzDuTOHn/Q+RWNQoTy55Nc3JIt0chAjFHIupGmYSU
vkIgrLXqdHtV4QozFNQ7Mvf2E08hFRJiXsKXI6LSTkhSCNHzrRZkowLogvkSHyTM
OsqI0EM9yKkBF8CwGUgCRAw+DylBH2FitO+yi9yC46Nqa8h9S1H2s1YMVP1fx6Bo
Hw/v/5+X/UTwEMVtcNEasQ==
`protect END_PROTECTED
