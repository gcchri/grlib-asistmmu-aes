`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Utln0n1joQ+z/iggt9oLqPyJZ62N+kMfh89siSbqj7Jee1EMaQBAoQiWSbP/Q+DR
O31Q1VTNhs19d6ix6L1L6Z+1E4DuhGoUdDPYi/7vnMmQiegzTX61B/ScO+8HxqH0
xXQ9uXcQHmuuKIFkdfgsNYom2lSVihCq+tmJKJjtNNMDaLcoImREPRyuL9XBOb/b
3u4t0vYXj07/5ZRGClygYBDcUK2qXJ2VqgxZGklFJX44ZFXNSzLotSnNBKRxfN5r
1qYDUHEUbl7XRcapjwt7zIdjWJA4LajqQOp7nT8BkaiMjT81BVRlG04170thKqNT
qmcnCmQC25q4+TdFj4IyD0vH+lGgxKG7sXTAvz+62sdUyQJtWmgpEL7NQh9kwbYC
+qgGzisz01nGmTWRmjkCPnYiDp72cBrYhp1rdaTHZdhsCUr1wcooBltHyYiIMlF0
omJU7/gPQWeJQMj7ccV4ziTzoDogdGw7hjEyf7gGHwrE45I98W6SdPER3hPFO97h
`protect END_PROTECTED
