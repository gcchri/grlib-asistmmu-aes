`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B1vjgRI16snAlKav77cnjAL4AUP10zHusCV0bIRhF1ojSpxTMFpAJ/XW2t9xBNVd
54YII6JOyGj5wmWUsHy4vOkmcRx6IF9HLt8lNDfGWQAqhWB91OUhTXSgfz1wqCL4
MKN6TC/JATTtN0P/0YGo86TLS28ljfJgSvSffeCKz5CdWQgKDKAw4nxe5iC1iPeK
KCD5MT3WBfiR1xJP1yAODycOqQ1VHOgKZnMylhz0Jq4mxTwEe4HH2ontjhvh0123
OgST+ui8YtAHr4AgxNEW2ymq9N74HUDpkwr3YXscbGpHMBDM+WIxjdADOhKWl4Ob
x8b7munDxNLE6Gg9BVXDbpPVAhtkiD+QBCPxMSQaprj4l9z05IB7dK954DPE7zwt
Y71b9OERY/iy40AmBrQL0jRkDmoh/+PVGIP6C+qMC7y+aExRncOtIBosEEqWFGn0
HW98flLyIhcuO1EbvRAEiumkhDrVar7sIT48vDHw/Bcu87KAQgipZPgWSju7tElR
IKcL2STtXSjDQB70uU3OqaMHcTsOeuGYN5kzSOn38ehJaBZzVLnIOk61WQsFbILa
vyNnaWS05QuPKPcN/uRK1Z1neLGzwYwD+eIVQYMR/K31dtUvE4y5/5f/AQXn98GP
evo3PqmEmqiAATy2rqAY143vzI8BeJfSDhNozdvwAquZLu23kY4tSlZHC0TDIYWO
GW9N1WRIp8EERRUas/fyACPICSnIYCPe0xEXNoFB6i10dRslgTiQ17gsdtP4EAUr
4a5GVg/z+tjqxoIJL9WordjdplGu1Dqp2Sa0iLmkpGtLjDw0GqaDkVbDfGjSEGsj
TPKS05P6d8x90cmS0JSdPFfNP4X7GDPcQDo2YZTkKsFpD7/dOa9qa4FFkENRngQA
z/9CQl2hpZ9vaBvZATwvGUNRky9H/2f4koTCmYmtK1Qh394nPTipdkjW0eYbJum2
sGPYcRSSVWN2voTIAw+T/NM9kXKVYnfa5Cib4qyPXINoRwUzbl7h7NGlCd/Rim6O
uOyGo78doEsgO6H8qASbhjwqGcThlYNmL0LkbKT/kVGXTQhPmr5dG5bxuEt9zphM
h/5p/vxbt+x/tEEyrqql+z00BPVR6htwKB3nD+o1BEvYOiEJkScQruKyvtemn4Uz
ubglRv/xM7fH+IVuF7WAMX+t12cjsykiy2mmrmQ3rPTrQ+V3ICO/RRx/cXh2NY5y
ypRMroTS/xwIRR+yIxgRvAJWgomnH3yFdkaT+IHDuUkIq8q4jckgnUFFaDZFsaXh
3BVGxkIxQ6mUXBPeqdi+vWK5Iir7xFs3d9oY1gj9miwZeKiFn7FEbbDzdzsBVV2A
RiSJlkJL2wIRF0oNax1S5y9VSTG4FRvTLL31vgL7JInGpVM+Ow8TjWCku5RuXBRN
q1nRbq9fAnG7Zlljcsp/Q13o+pCjQf4OoAW/dT0SKwefeZspgexdIUlWJeJ2FFQH
b8bBNHiyHfxDh7gY05H6gk4lh9cwbQQTbBEAjDbPf+phYON/5WNaNIRW6SGj/w5a
++QoPKsDvK1+rysUcTusEFXDb/QdkP1DVOFpt8cwzjG7UYHuIcx/a7kX/5GA3g4G
bGT0gjFiGt8rLKXF4jkNO0bFCbCmwvx2GETlQmACMC1XVmJPLfvlq4B5hqOY0VqZ
31AdAVbRw9QYfZlCuaVC5BFLW1rymXSlFjWrhqRHfmMGEYgO/Xfg+GimMp6IvsHh
vne6VwNGzegHW725GtJFla68LO6R4lcsLhRRMf3zVpZtHJTjk8FyjfhHItGEuohL
dQo8KfKFs13uCg3/MrAh2PzjK4IM30y0H+nW6yaCl0wcqsQTLs6aoetvFr+LoIAi
1NFiA1SB0MKON1f3hfjLFYCxFE12mwRgW45n++pepzj4LxqDZA6hVElo/A469+gY
hjIm0EGS93Sv4g6gFlInTJlBn+nlXBW4cf/Yd3ZS0ajoOZLVv8AZoc9s/I0zLjoC
GncV5j3wOKA29B3pXOl7b6qXDcEMInbzLHgb8J8amqTKPKAMnLgb3XkNp6nCTNom
miV10L6+xn4wGgrFF/WhwsjGuZTyLpFUfXeX5oC0m+w1Q3v/V4srAQxSeDV43Ty1
aTfjlS+9ddqAtQ6FxL/FNnynbrwYqgRX9IYPjoI5RE1NNhC+NpoyjuzomHLYylLC
XPwBe3sO1MZ11tcPoZTL9nGREBi6xUY9XGgFyKBeW1W9Q4i9JbZTJ8kLw/M+4bmp
MFrsKmfifoE9gDMLpCCNGGCZ4m+AIzpJ7psBwq5Fxu0dCd1gyCohzQoPYijW4l4A
xVChFRZ701g+mRGYtpLQlgn7m5JXQbJeAsVJkLLRjuSxDCbywNGWeiCoJFeQDBWo
86Tgkb5kt6HaUPUPslEbSvX7qJKxVgyN29efr3r9HhCczZXNmldEwVgwXqtVrsce
etccKxMSHXtg4NW9QQW4/PU75MCpb7ltBFxOMtk6JQJ6V3b5eC1JBOzY8aSsRKxp
r5ByGVrW8adQ62xPvjVVfzR9eXpXw4iEkZqxGy37DtsRmnhYlWXLr/gfcjjpIry+
dHJ8gwLOYdygNvWp73NsPJGxpLo5wFc/awAjVUpyaRlyvrYObPThw2Vvb3HOR2nl
i9P8sP2evyemUpiwNW71NWbvyvGRIxgve1GiU//U14C9I/p2WlA8TSLnNh2ylkr+
xc8r0oewp3xRfWJWCm4aFCiUXPq3ZugynkGL8dPYBHxi58heiJCCDrczAKcVMwoP
BgGA02jI3jkAbLCWyxA1L2CyDbcl2JgKWYwIkw9GYYJTpK6rNGEIyagmpDMqDdFl
y5p6WatcUkjhQZNhURcx0A==
`protect END_PROTECTED
