`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kB1cXSO+l7V0Dp6n1juQQmM196vTjWxPpjjAnJtk0rrmsSRnbb+ic1/eVG1IbcTE
Cc6oTmLuModA8uyvWu+ByYmBVD0m0SVxhLoPQYzUjx+y8prUOfCE+BIchN0qvRZP
1QfjQjxZ/AEwv/0m3hmS0ZmuoXNphUkCCD4JzA0cS4oxz4xJIOpgfm4Q1/ODe9g2
wNGqZiA+ugmee1EhG4svP9TsulvczxEvx4s5UK/AAlOne1zQSO4Ksz/0+7OS5/7i
hnMoc9qtzp48bxvyPW7AtUYoJLjUaDYXAN1IWo9sZqF1FedQnoaWZN2uI4YHjQar
77uLk++SUYmNYZRuzIQHR9IOQI9sXFlucOZlylKbXu1kAbuhBlRNCVLQSR1yoSqJ
8gjfz8WK35B6dUovPfnaPjTArPzOymqsWXny45ds3l2CBtYTtw7EbmCxdDsa0IZj
8MaPVZVhpIW9zkYJgRq2ZeIAJbzXWCuO548H4iIqdvBDkXM6ayNf4D8Br8Fx0vkR
oG8QmzgqFxyIYUfSJGEuJyLmCmtYRWLNiTaNiLBNf5VGiZTzxBygaov617fooqoc
/AXD73wyfTtOFPhiXDAN066lKev0ZFlb61LqwJuz4HtAta70mdcqIVxChmSQhqTV
rmpW0lujJ7AQ18VmEowPVIqF4gx2PDyqEAngvBeKHEsJn1/f+73DE99JTMnqB4U/
o2xAES4Cb68KvomGIPVfuEzk6FIp6r3XmO8OSlFDitT/gTrCreg9jEOKcQNoVqwJ
WojeiO7vElnt65j3h6TNOLIH3+AWAzppBb3qgFWS8tQ5XCufCfb+nykTfaYiHVHT
Tjj4ZAWVW16+QTnbf2DlFfOYYffRlJVEhmycfdgMF7Yf44hOrJIW6p4a240odzrR
V0no2PIXM6+4chjBtgF/cgiIhgz3bBMh4z6+x8ghYoi2UQqVdlFjfU4FH0fcz0/r
LbdQ3ZPDS1l2+2smNn91c/FodDSV1TA2OEWBY52clW0wCl2RaUY5g75iZwCrIGQ6
HBUQGR24Ng8+AxBNK5/PCI9OW25TdXJJVxzVZB7eQ3+mY3to1D2VBZWlYW7FiFaN
4kMgwhJez4uGa0Uk8lSFE5XxOOa8RYWirz5ixZ7w9ViMpRjDdGd5iP+rJKSDJRGb
iN58cQe1aExNo4zMh3p5vVTGe9WHHrTx0aqkV8ZIFqk1CyK3gBBG+0vR8Neh+PcU
lpk0xLWZ2uX4L3jcsmP+j/vg+ur22o87gVS8iCSPV4E/pWYpnPiQlFZT678g5vLI
ZpCICRAeT3cz8NttFFf/R7aKenvklEWRtpsrlJTV/WZmk9f6oCjtoKLOD0PCrrVE
85v7wHM+0WAVCKtifJLpNNTfNkekYNAyW7kTh+gFI6lreG2X5uuEKcSVVCofiSdB
unQD119OWd7JarG9nZxu/wf1/yJDErWVrPDmnLWWxEy0cGy8c4Kad2LYLepihdR7
+y6AzwR32ljGscOFYqfl370i6ef//ciL4jsFG7Y2kmOeDY7YAC71EZ4+HLqK+REJ
7Afcva748qBl/OcOeCmpJq9KvmRH4qaFEIZLeYMb3oyPTMCs6cUGHBCljH1p5O1A
enm5F/jKqlugnrh2JpCwA9jjRDryNrTEGMW0oUMULZ/MyTMnuAu5qLrPGRiaFfzl
icAOWik2nlGsyFlbVL28RhSKvbelRVWWuQuTzLhWhgN0s+xnFFVh3THu5qRqmE+F
ujcgWGOhtf9pRZBstzGcd416Vt3+4BNM3iIsEQO/dXJXuZOxYz4stII1zuCb6OUH
jjOI2KB0oBbH301JsPNd37uH4HdCXE+7qUecC/YmjGLhZ8q7gb31PE6Fzoyx20Sz
3MeewJXrmUva3KFUKe94F1IYA/C6TE8LjGM2MRyuvjcH9G9xZJ4v0LCbvdUn0puM
YPThO71bdIREF+aqiIW09e0OJMZNx+ZAyz1yyH8x9ve0AJTV/1G5ZhcFT+/iU+KL
PBhvCwuR0vhqrN07FUhkQSMnFZJt72+VGcnNJhAktuc6njqyN02/91V0q773otJW
4KLbCsx7mjcc73YZPHSTpalxKwhOGY2l43lzSmrq44OjjmpJVne49+eOpVFABzma
RJ235I4WYCAQ3BNzSXO+UGtH+hOGUTjBfjc0X4MgIevigO6jnplJr2aTsqVprwUE
w58VkXtBQE47RExe9Kc2JxkA2kE7E+zTm8cUYF3sOUvehdQA7XI220vwwU/Qc3iX
3Hn/UWCFKjNy8AY8KjqVex94fPpimFSGOFR35pUbTB/ekSFjpWR11FXWcNIT/j2p
gFoX51Az4/Smdim2nqZE1CmgeATEUajNPtzx4Qll36IDYol9eoFZ44ps2KdnY3dQ
cESNPjR2hAGp9kGm4czo2p1gh9e88aN0qza4QMx7JL96mTShtpX25CW84alT1TR3
FslHMP9gs0TDOiyJCQf6/lWM1FNaVGUDYISrVa8feHHiZwVcQjec0cZorIrqcQlp
Kt2gmg7KgQXhDhluIOLubjD628HByMfEgKRgHGND2HQx6C+kQvvPOg2RKIqa2COJ
mx2DAQE10YTI+pYcr5/ZtUDySHFCwIKVrasoOOiatdqFMmGsR4Jt+5ZIld+Ig03r
rKAdzbFQUie3iKMXnMvzvoKb5mqCloEOWBQNCMuHr5dKNb4LYOTSU2bCzC6Rvk+s
AzTdqnicn0ustmdDuyi4WNqjjnpNQFpogN4OjC9FlGrKekz3rbtf/+eMfH5JwK5j
Z0O5kKs4W0VQu5hABfJdI7r0I6TuxUxalRksvPxaVnwkodGdM4qs/a9Fda/WwQ2B
qPjQgJh52dgQvrZGcBDD8eVCYr1v+4OENCm0Czm+E5+42NWnpzPeQoKAr77q5Cd6
lva40zhiEO7ciQvi3s9JpJbKBbfeBd6yzpHJZem0IHg6kcMEiAbQrp0IErjgT7BB
AEUOsvIGhLDGPJlZLXKxR6/fF/1UE/3EyqxaLmu+wGw1LKBIJTi+MnCKL7x6Z/iQ
/84NuQfFR951BaRAT0ppCMWNCQz7odb6dPayErNaFsq2OVTfGVJUtEjA7MtQ20y5
kDfTKW4wd8boBIdQjm0Up8pqb8rARC8J4fAVsS/XOe6nn7AVsu/lkQCegcrxAHab
dox4MKOKl01M8rfS9VUJSGaEBekni7oJGGdvkFDiyAkGYvfXCBhRO9C5Uw7oPq11
zxVrqOqd/OVAVWeyjVuxu9hbAB1Wm0K1mnZ1VDGNelf7eBxritoCw1MJH9Q9EDvd
hSLmHHSyCFCImRU5cRQ1TK7JVFR5fXVNgfIr4Np+0BLk9YzF/q6A0kSl90cnNNvv
fL2BdpK+o37cWiV5bLQ+cP4WFGAP2hR1hfNE0763DZVNQIvMtmNK19BIkiO4VWgR
I8TeTRhsQPHTtPDLwSVfRe9KkkAomY/+Tt88ePZRcKBu3mr9VoTWGHdju5YxQlYr
atEIwCuCVLX2t7sHJRis4r2ddYTwTSEdem7EqIV1ne5NoOXRIL9pLpSy8YAZOnrP
DoAVInx/5UAllDPzKZVpL/EZmHxMa8AR2RffoaKCSDGRpT+Li6AX1/OUpsvGXGzk
5cyAU9Lz3+0nq4wvVN3UPw2HLakVB3Qu1wlWSnk+o+8d+HXA66f8Le2lnnGTgt8u
PSSw5rwFAdhk5jVIG6d6nGJBZ1HGjMck//RMpqzyG9tFFethyOU15RvOixuwghcZ
iawc/HYWR33UZcCLYGogEQytctZ/UYzJ7vkE+5d2baSbbzrdTUzw8Zqc3WBndaY+
eJybxFL8TbPUgrT4ws7QS/wMBzA5aenHpIQEutoM2FSiGVhSCsyqADJrqBqc9yy8
7bdqKwEKzXnlrveCr/spv5uty094bOC01V6c0agNFLbJg7wbgGBeFdF6t0y0tzTk
wbxNiWixkDpcq2hjphy9+btTe7tSIxSNKuzj93j11pNUScAmSLalZUh2CUOlrZlb
JdHZHQQaYCejV/zcjOx28JZgONnPmiaw1PPhpjeq5ulq0fzAYYWtFT7nGX3S/eYT
Jb2hyLx27nfGuI/GYFEbb/u7xCy6l8QTspf2raQ+ShRePwEmdbIUfv+UuIDNJEDV
ODgwNmByFqsiekhjrhJTBPTJLnF0EKGnlEjkEB8/RINT2uK0fwvACJLV7YngZu4a
nMhIDnuEvnm8wT9YFeNjOhUKXEvwSdbuvwL8rj8twUAxs8hxDYu83JgvmEVnOF8Z
KU4hpeNte7ZMeaQj2Dj1EoEXlzH+FKrTfstAVzkzkzEoFfTpTcc2jMMBpCcRkxg0
JZNeCGD1ker+jSjlqX0wi9cYIcRHf97P2KW1nSnVT2fJCTi50UzgtONFBuZYrNeg
CC1E8gz+euFH94JGSHRcKR5f3/rLvKvMPTCrM2oyjhTVaq4u3JF2+PdK7s25Ul07
IuL8s8jIJ/J6atR7QEQgBd4olmbzROu3OdN32dVs2E+5uwKvxGW7dXMnLxFiNSAH
ylyDQBdfpL/8b0rRZ5D75Q7fCPFqGxp1SFK++oOKEfXXwoTIhTPjUU+gYErwv+Z9
qhyIJHS0EZc+CgD9sYGKU+uoZN6napYYZohgGUK3Of/L/iilH5SMOWFtkRoWGD0S
FRYQ+tyItV1JbNledIWiC8XbWkYgNBT3xOtIm6qNFKoahrm57YcrpOn9jsGQdkwC
IoD4HoS+36a6f/yFGJky7u7DRc6Kl7WwOWD8/paFWTnagzwaXNPZ/hnlIQo+Qi4H
/LBSrl6vkOZivQmX0oiDTXfnX2sAmSSI2EZRANWiMTuPjvwXLopTlTlmzMp10C+5
zczxrP9msTCll5C0aO6kjrsEH9gU3hDrgtWoJ7sSbJGjTBzkiyOxwVoi3RRk3so5
HMf9ZJGypLrUBhbLRzdk0CVhCCURKVujtwbn5QXQlUXcKX3h9tHG+F2BHU2+atao
2DZmIdBJ1EYRsCE13YCE9NjIbGx0nmA/llQd2AJv7Xao18usnIWXMH1KOXTPJqbR
TBillX0Kk4c/J1X4JWBKgdO5MGPTwLWDQxW6q3T76y6pJtQ3wEJcrq0bjc+T5oiU
fD++9KG+Vwf93tUMgzxaBewJds2tDOjx7qRvCYKZ524XnrosdxDcW1d85Rn+yMcZ
32dBezeS7OMsKGqE5ddd64/9c+YaR/aUUhyqovh+m0mwFCz1lSEY+6Ixy70QQhcy
H2yXIzHl963Pbi0GXEpi5xy1pCMxBe3xgKKmg3Ve2hExHqRQ2FW2IyjkK9+PO3hG
/CZiMxnrI4zjmiFUykFz/lFWFHn/CLxmdRrKuI+pq4Z8uDOARd9C5cAWx1imulpu
P4xfEFBAPbfw7l3T9+kHxFsnl0jT54/Mqr33xDpCWewQ8woMFDqKal8MBsSAKy90
WQxI5TQD6m3s9HejtqQUXEJIYT3473IzvunatwlKkI65cSMRePKR/31MRD/J1hnj
ORBp/vTG0TA6qpUj/Qz8c6O2vk75+cPeBQULasgbfdDBep/7xbjlfBufqvKbSCIq
g1ZmBAF1PRndNTCmbXmnxlFo4kQVd7Kzloi2XeZzUQDtSIONh2pTH1pydOATMWKC
GETCv3lMaE/1EKiqkThABzuo4YCgeBEZw9L/J4UDBr5gzRzwrBdm9l9IRbcL+ZRD
YXrneoz86yvYJaJhcQZBgED1euhdIOz51mfzOXJQc7fONEtYfk4lN7kHDBJG+lhW
Y8LaP0ELScxwyyIIN21V4ee7HLetdI012LTXJNq72rvgjn+B744LCxyLX8iKnvQl
zA7cwbgyq4EVeAJq7+EowxXjA30u6lK3qOcQr/NpWnTSByVupSTstqOVNmuWT66a
6NiynRNc3BCK7r9I3CPDNPEYJuMxmcd7bOrt9Wn2cYFbK8h/S/grfGZmO4CMwYWL
bpIhc/Hj5ELf2TbNioHJ9K2D6UXzNzsRi4/UGmOoQ3VV+wrQWRtu+V+VXnvtnJYx
QuwtWSljValaiGRzdsJTGt7Sy+yl1HrWx262pNqHQCGkhhLtdlYKU9/AV7TybEmZ
pPHv7+GlxBpD0r0y29PvRB8myO1rCj0vKooxbUDcC4dE52zZ3/Zt2amok7fdlxTq
SzGB+NCnjDzao0yPGEjw/gNmPtjszhEGFtz2qUiDo6HCQETOXwBIqz9A7nCHHOaR
k+FsKEp6VU6cDrtUCSryzGRpocT/Qr4zzKZ4HrVwDKA2hfxrUYX3DUFPM8+H8tKo
mOLBIXTNo92YxzXaez7HlqkNClsOihE0YCWJ5oU0TSm+mBInPV8YL+SUiaS6ZzvH
BVc7w7esVlLRkXhSy9QMpWGEYO8o1QQf9fJPGpqku65GwrKqSh+oSV2bpsYByrzP
v8wH9gqxA5U69a1S9pHmWlvXdi16sh4+SRgK1+ouLRMAcLjl3YECOEVQXO/yD3vP
W5C09wZ8Q8lijaUlpcZVGJP2Vg1mNhPBWFPrjo3LlvfiAs0XdR8rR5fxOePAfpD9
jgQ4kc7nd7AEqHWiwGQyCY+ZV3aJD6KlRVqWCs3NQ50N6BZ/h7Cz0vH/mHukCZ8q
qT+Q6NHcCWU2RvHsTpb9r7MvDgiFz49ma5Y2XnlVbBzwi0usvsPJ83S0exkH7cVD
lPiIJiiWp8mlcVz17VmJ/CjatKapJzubF4fAQ7LdROkOOHkbD65S9yT3dFQlc00o
fAkexjsSxOoP2HzyaX/Qpsy9eVEZoi+ZmJ7nWB2C4s3T78we/cX2arI0XS03Cyt6
qQGRok73vUOKkzCNRtFYIKTtBWZZahnsnfUy5SBidLGr0JVDbeWVj3sLpr/IPpPw
XH27BmcNVGFKokB8FZyXuQEWT7+IYXY9cMQNFuPVt2xnm2f9eYB3yFq1XI6FG/T4
IjZyLMbKIwl3XpTyDZj4/BSg7/3lpd/O2XCrGEI1HPcWIjfQAJE7t4NwkBug8M7V
7l2O4gL0thMU2by+PA7FxlZTS7XELSHY1naTv3/RXQdhQ2KAGmiCi/isQYtQkpOr
XcIdDw4SYGaf0DO3AENeQNTT+kFDAnbAP3IMf1jFpz/X1j10sSsaRTW5qqnlQVRH
4P2O/SYDGaa2RpwW3ZMADk7CM/LdY3TZO4xtPGhIZSfNcRoEJs21AvcG62YDBX/c
BfQFxS4C8xWb9yF9jq64J/osJBWQBKlvgyUxvNga6bqARG+FRCtKAGyzNULWkYK6
MzBsKvT6gA82ZZKzKMnXsfU9N2nBENCx75ZrI2mzjbsFjNINUBTdqccEBVmwUJgN
WZjymGq1DwCkUPxByAmsb6TQAkIu+yF9uHNSWvduG990shyY2JOwj8bGjdE/DNsz
Y/CoLzgfIk4bjmmMPFN8+pAVjmNC2SRpyAYzThkDlkViTO7ku2VgUsAW+9BMWNON
Ig/xuwcsiBWIKTJA2+WpuHZoVqA9OlRbePAE8y1Z25LDeG1MRwu6LOIOyH7D9Yvf
J+ZDp1HYrdPywDlT1GHoRm9ijWHTFMhCIR0b1GgGOTaPRIW4TjetrSSikrBHH3CM
4xpwO7WEeAHRLLp9PbNdAh33SEH0YInDlaKcXSkDB0TsKcWLrniBR+6KNIUJcs1i
HQOig6wFShx4WB73iRKuqeh0kfjUvLkRW/Uc0Y/i2TGfGpn4wiJ6aJXSvVEvjEGE
JDUYMv+UoYb6PUkFpELljNof5rLfSEgUEtP2uK0JYeUxR0jdCmtienMolefrpuXX
HLdFIkDL3pG537xPze8tm2cg8zqEV+/WHFIzcPGI7S3mNDukaDH25LwldcW5NGkW
QjR1sZ5G4KU/V8Exc7bLBxRmbMAkGN7lXTo4/+Dc+bw9sMvjgb8vEkvG9mgrLLZY
YzzfZ1IyAHQ4uVpwnfWlAC6f0+9Sj8uAg410hdDz2xnFgnK7cb2V3xJBp5BI1ubn
AQoHGY4OpECj5oz4i2q9W4rKsBxz3WI+3xnXA18CRPN18VAP1oHe4rcCIm+XZeEJ
FWU11AD0BX98L3VVPLc18hJCtEiXTP4dhuF3Bx5lCbSarmQNAytjOEwkd8UwCyPx
XYsygD/i8O8ongD+mOAdK6IIMIoIeDU4zkzbJVKA9txM+VA0aGefiZEPUmQYGy9x
KNMIRtYFbcDkBrtLUZYUFsnPRqNPyUqDFN8ME0NIBveYfy5EMTZtheoBaFovbxeQ
nK1kdyjS2hp4Hu+FnpdOf6bj7v1fF34C25E6Iij42JGX0OyrNUtAmj7A8W9C2dsS
mlliXe2Z6sDtZSVpuqgKgFYX6rn3cGb2Q9Ux6gJjwaBhug2BqvYYYyUKH2796F7S
Su6qJlWFPJcSYjaGXHXmsm+Vy82HZLOpp+e635e6ZjhrQowsAZRfxIcKKlEfyQpN
2LsJzfw6OLDWZRZa12DrIIJVRhFTLDipGbShR9LOiEaoZNWX8ou2ztX7LH3SkNK2
vg8T3IBxRpzrhcXQcqGEMvzRpIMaT/meUYdTXLYg9+btzWMfqxvl1BTfke6URc1Z
jWZo3K8zhq1h1/AFyzGllev2wrejE62e2nPCPaywsNw5LiR0k7pbbqz33VZupX4E
w9PTu3k+Rku6Ac4gQ50No7owOT2606wMQgXVvzFXD7A2GfagHXICji1Zgns2+8B2
4g2HUQ0B8qV/eHJv1ZzBK+IOAaG85+0/7wHCw1t95ZRXstPRW0Rn6jDrkXJktFKn
YkXlR3lWOjL3A3xjb9aRcYmCS4ul9qiJKax2rZ7g1oQyUJ/EsCzjpd8cPqELGnWj
0lO1hLEmtqMotCjenx4E9w6VHcg7IslmkjzYHsCnxNFcQZr2i/WhXQcbdPEL4GxN
Jg/FIpXeeihJnFmbBLuenA3OOsK6Z0QbtzjjnX1qY53GDkax1SLGizhWb5XeFbUl
WJs9vRMaBjBXvk2OAtqyjWo+U/4kenxyBIz861FC2FNJ/PZDV3J+B8sPN9iSKAEE
nE5qp8trTWSVILcUyOvnfRxKzsy9qovCiMuJFRbTM/vW8FfdKRzGEAuJlE/F5QnB
0q65AVrfcQsUIGf+EFth5xIlWs+wuNSHvCRJjzMXm5FFZmwhkg3NcpT1mwhSoDot
b5x10oWe5ua757LTTP26brRWrPq4mlVuZc6L3cdgXunflQ0i9HcZJbD8rHHEe3mL
rRRJqPDtK2u1xeSfXFGHBasiFlf7ja4L3tLw2nD1Sm7HG0wqGk1aePD6bcxTIfvk
6YWJA/O67hHlUOluQPrUx1ZHgC0X98j4A0/RMlSZhd1BtrR5IveYMBL96+Sh7Ms0
k6Kop/42PXMiP9lxJxvalBgJCugoIAcjvBSfHyhZ2gf7Hg3FXJBoowfTUhWLxeQR
Ys1LF7TqBGN7crKFiRr+IuHSfY2qaq2mQUCLqviiOxZJPrl7uEG0YZOPBqBTU9w/
P4ahw26yZ90M7vkShqjj6wgykDTjbYygHd3duaNRvld1tt99sT3mN76cSUpmQAH2
nIjkJXC1OnEDHqGl/qEYlzQWwEz8xDrRKDANlGMtEXgplwY3DFmMW8AqKGAHmmPv
yz0anza7KcPi9IHvBISSm69L1SA6vqbI+z7DrGr4hqhCndbfBbmTdyEpNUtCEVEY
rrcSpiStLMkHKHePQ2bwYcXVJEa3Xu91sKKeb1fVPvmu0hvR03lh8NSadTJNKm0C
k5lwG9a2s2RAvVCfd3VpzmauFsfs+0JOcJRlDNWw//mAYHtvO/YCeR3rFi6//Eea
Q0zDUHrn3FNZmTnLlLCYDHoJGFuUNibx+tS2iHKbSDmxP7YiRacc/9sMKtNbFDf6
w4PY6hevTwAVRRHSqz5T667egaHyl/z9Q/N+HxNr+jrwq4gIFIFT47hP6GH1yi79
D0ZbGUdnPe4UAXqt5MfBjMbaOTrB2MygrF78kiME+aFvzlZI9CKkRvp5K+mpoTYw
AYI0V11QZtZ2bjDwQgoHayqD0zsa1dIFEAJYZooo5+5GE+WlR2IguzNe16YWsBeO
LkdZWhuca+71Iq2KVGRr48w1pEkKUakjroBEPQtsPjRhsMxTCy6c4CtQuG3JB4y7
U7nftELuXXWWE+4bFOD0c+EIOJ1IzSRrAzdWPtW1GpiL2RHgvy8eculVcfy2gaC8
c8daqRhgl4CmIiUbFcdUvV5dA7BT8Gq7DWtsg0b6Jkbn6NlsynBdo4h3u1O3grOr
cNDEw+ck9L3/QFwMlECwlSgEfpc1nqGDOZUVxMjmrlNyHiFYY02ej7+lqAmACpHI
4k4eDXLsKBbI+DbVZRZBYQJ2AFKDjrz0rwXszlimSRGQlQtL6wzgRWPWwUnIUcyq
gPNYvKwpyJScWRrWSWR1D334NBlW04yjtH2B3f5VBgAwMj5fZxUF2IP9SobA/wUg
F1+p3u3Rb5QRpSB9xVtWYS8DLSBXLrN7yoCRmh1FGIQxOXPO1Xo+yGYJSATeD2/L
gKBsPf4G6bsRo8usJ8owjZC/V/FKgLE0KD9gfjNgWlUXQLXbQevuqob17iWR34Oc
0n7qc50LZP0ZHGWUtx8zF0pTW8CtczH6aCs5huQOjVIymOlGO1PmlsUl+zyOWApS
K8YWpNVIi0pl2LJElcr/Pv3zOUaEbw6IIKTlJ+5CJgAqQ6QGT5l/L204ZaYctAWE
0oqyS67acjz6D/yAAeP85plioB70KzrCYaJrrwFWBrVf4ybvnBy+sspArosHrYwZ
ssgifvi+idwLHydXR7h931lFeR0LE22YyAqTN5ogqs/ljRPiJOihH5PTH8W0Kv92
YupVah398QjAnBG/dCLoj+402d8GebOrTt6boApXngOEraxKDDLcFPcLH//KsAEB
U4YVcLIck4DJktpa5bJEwaHdIohXuHq6SDxm1ksW6KGyXbVH/0XoaRyOSPaCKQn2
ksYvgFy7oPZ6iwjhzy/TF9xD+boEJw3C7x75rba1jYWiPvlNvB+Yk7VUN/NQ5GiZ
lBErt7F325UEparYwoCM088vf/ieHCZGbgus6Guy7XEjan8UQi/efskxqFQZWOQo
RuX9SHAWsLp198UMGZQ7jbrQRLZ/eddREaAHHfzKDumo9a7ZVykroY/opa4GVGJT
kmywOq3Hzd4Iv1bINczvQONbf8ZAA6jDDE1y+L9WIRZo51DudRA07wl2yUzl99p7
PMigz5Url5neXekQzHevkSAv+Jah43JqOsUYVlW5li6PqLfticb+07+eMwhk7LJ6
n1nnOPykAz5MXac/A0rgCWCvdDevsSKwfCi42vVgxwKE8DhZxcxZ4Cc4kbJTF5Fq
aMIDREZfCsDncDtGbbnHUxcBD/+4BDptIiOdW2kDV2YeKB5xj7Y3sIclZ/vAW89Z
Jn0HX3j2P81Jz0tyorPYvnABZjLbUv+b+1k+cUbi7TD9MVY2NcuAm0cBidpBNL7/
VsxddLGu1frBmh2LAQSKu2cEPeDpPOeXSxFTsINhhg9VXZ05XwiJUzZxei9HlTIA
FIxDGpZ6LSw66ctf973zCnazVZ0Gcp9Rf1QUhwirzT08IFvZkBuxmVKzReHUpz06
gmdID52StQOsuYWkh6nzMNqK0Xma9U5qqM54q45uuX/zdGhKpl1HOVOw9DVkOf87
pv0ZglZ5FU9VovaLVMn9qvMkFfRUmaVaY+FFTLsnQczpCvvOWEN5CqE+wnURaBDA
9L3JQVy4RLTN/OIvjK7L0z9Nl2Ry+VsIPS8Wla38jAo0+rufFFQeRliS8YcDXCT+
/sy4pJGEcSO3LfbSEa8K9+O/4pPfDQoKoIwf4L/oyC4C/z1Hq8JlgB8EkmnNSiAt
Snw7uuzar5NKJCEiuvp5sA+H6FIE/yw6SHLtUDYIDrkOSVYXd0FpKzgWcaNgnF3r
QFhzJQEARblfJA9rC3Dc+CcNAzBCSz2CwVkalSzdPVzOy4XTi7u08YGlr6vYj/hS
sXmBxHn6xeQ2yDpc8jd5h9Re9aIezZ2eA3Kvm7tyVQTtGh+YQN2otAzna1IK5Zre
31jIfCWjMuF1blt3pJdw//dBdJxOKCeb2kDmJMxsRbducAlS+euCDbRjOvmkxswk
nZpE+um78ltwVyMlXpsmWe5BwJz1s0XSnllBtsZ7B6sQrNaUKJWlflRAD10WbboC
nwmbyQ9v26Ms7OPaFXil3npCPEsIFQW+X1Xug7yyv0B1aYARaTxanC+6G9bWstXK
3xQ+C0+fPERS2pNlut3NACy96ni6IeCi9gJpY9M0b1iqmhxuMi3PT/CgP3CDo8g7
RsC40cfOdMsFqal90c6yLjRjhvJZ1wFjZILErUVDaSwuCsi7rBxUMGShryU35Gca
cnbUdx8Eys59/7POD4xD1gVFu0TVZxFkC6ZxPvY176qjgesTrvbGzfu7040enZjg
t037AxFx/dkP5aiZdKMQlrxcq7aDKQNpAk5Pinf1X5QXwCgljPyNvizI1aNWFgqu
+Zb9H91wLp00sEgg8sEsQ9oy2dXuTwM422bREWMJ2DAQpcXItK+p7abESJKGnJxF
g/JpFN/D6h6P9HoozFsHyYCQWHrU81nLOQ2cTiadNWQlXo31YdAbd1kLid7hA1mK
2kOlIlavOLofF44PCix5Tw4QmAADXxi9bKeHGwaGYVxRbwCr+usBUWW/t97c+wd1
H1tlHfsqbjNaM6jnb5Wix7xHOyO+7DuA3eX/hDbNlPTlreq5J3vakIGaKgs/gRMN
HQwWoSm4VUAg8tYF33O+XnlNDp2Jh8uvCdJ+cfyYxdDWu7cAXbx+EmMOMmcqGIr0
7Cb9E/NbA5pkoT23gd9JAgtbUnwSlSEPQ3IqEFZAv0xlNSewZ0ITBdEciu+TTE5b
8DY8dBJhZBs5wzCrJg7abKH8XnwTYlaJMXZZbO/BSMcFzEhIOvvl3a7BSH2+VlWC
vkzSM5lpLX4C2HC71TVtQLk0bKodnFIhOS3w+K96YyWHs/bABqGSQYByBzfvTmSt
pK8KhRth0D7pukqfhQ1WJMmRl6wUe3cuJVRE5noJK1zP0YHmI4oQsw+zSXvO5sRg
1ITMHAe9AhcqZD0dAaJSjpqTFz8gr8dfT8drg+N6+DYZMLScXlgKy4q54rdxwuNW
d7pjHOfuEguSOcesb3IGrl4YZljwSCkXo1+0x3ij7bZSppjrbVRY7h+dxJgLZOM6
YzUd3p/Cqg1gky1xDnTuU2rMwe2OPkYRCdqOnpLZT/oKoZ9v162mQUCPi19aIbC1
aPbefR7ahjI+e/5V5C+S2YNMpi5a3K0btw1j+UMdNuCa+bQAYQZiCzHhE/gd7cgQ
ZVhpZHUvr+bHgZ9vr2xSqrSP0fbV9AAPD+M3+qGg5uW6kA08hijnHAigvFeUW7Ae
FFVZhytge5DPsZoeH4shmp+XxqMW+PcR1GydLpUMVjhhRWBinS0hch8/zdREY9qW
UNfEYW0jrmdDm1EWHU9K+v1h2erJbD8d/vUROn9GXMnq1LtYLW5z51bW3BL3Xs7E
PakSfSCTixyOi/YvWj+DrsDBAtxlKOpcyGn02wSZPrM4CPaRe5IvxkP2z3SM9NP5
X5qZTjp6sABxfnf18X1WSoIcVCGWVHocSmldXvQahIp1HcC12mitEEoGBxkLtpj/
4v9Iz5eW0oNfV0ubbWnyUze8YX2qAqFyw8J+6q6ig06Q6TXkIYt8BB8Fo5NFlY/0
aSO1bMcnEfYL0s/geRKjnkR0D2PTot8GnAuMLbCeSHa3qt6sLfMY4O+nxHTw8YUU
gGNlz4sj+1QjxBmkWQMQRFCz8dMtMZoMIElyEZHPtA7OkXfZat1fpBV/OOOlQKnd
5ncgYuwelFoc2kVkEAl88O7OEW2IIfvUeV3e23/XbF5kCVmp3pmEnjPwO/J1gSfl
8Bkv+pkdW4mshLQcJUiVmjl0G68um7EdYOo4TX4H6ymzajtW9OeS6zJXyW0ezrE8
V5bRO/gyyckqAObV3Dw+kfsePfLO2d8XC39Yq5ejQeIhsYJOHOmrJXKwBO1NFBjJ
+DP6IG0gVerIqgb1e+HIzUexy5H/RTkoBMyWJSNqANc=
`protect END_PROTECTED
