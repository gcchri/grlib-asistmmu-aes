`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tol9fxD+IjSGI529uQNuS/CYJ5EoVwU73/87b9ClpLggB55rN0y9k2UYnB0AR2qn
0mbZv2W+Siy3rZuDG8LSIqrwVKnp3oISLtEu7kve8tLqw1FManXB+U5mwcmjMFoT
Mf3GEDUe8CPGX3pDm+C37DV4y5WHnY6c6iKpr3UO9QSz7vpiJj9Ehu3JN7SmsheW
HGWVlIubu8U7QRDdBJJCh5tVCFb+f1ZJN42o7mtk4pz2uN+Xz+2V7xA1/6N5gVB/
r2rbXzQQW2wELERy8boCIhMVI5uBJBEgjA2ISYW/SKEQfjnL1FRA5T3ZpOwSzbFZ
srmgnUtkJH93WqT5hCtW0+S/9HD93d7LVBxH/lEGn8x4p7duEWw0hq+2lRNelAa8
OBHqoVI4X3cfFDgLvSBbls8TTXGtQ2l2/29jTC7VWnuzSQhps3YbyRB00qsC+uJW
ilgs+kNseTCRNZ4Uy276980XXzyPymPcp+jtm1UDOIvA2RAbXaFnUxfznkuZ5IjE
mK/s92tyFcwjS5YjQ39Yxv9bqut+aFajARkDtkhVumbrTuI0Zki96dh2okh8yrhS
`protect END_PROTECTED
