`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CxKaPowxQvCi/b0BOOcZ4bYVWkzZoGhQEtZ/bJ6eRBY+jT9VrJaHqVrQTkIxm8zK
vDxH7ONyLB9E46li8igSMFRlQqZE/9LtxKyjmxgfRX5hhnh/RdxLgQGIUA0J+vZU
3VW68tfB/tsOFVjvPfKStuT2kN0rcZiZzjE8dCdFErpC4FMBK9Wnwae4MC5cdBlo
MIHNsCjc2L2Nuqq7rUvcbnkhkNa0GLSMdsMQbevpgoj4V5nFHOLKFyn0stLKrNV+
+O1fB3zjCo4+FGGY/5UzZwj3VrHalWUhE6vFtZt6aPnjbDswpAbsnG19uL6n0hDn
rdt5FZlSlCC3Ui+mpq7XOPnqDyLgqP5Lx2gul+sOqF3nSBg86RMGb2PhEJ7thPXM
rFnpOq+fj3uo1LDLIbAMIsFsrewi04HEl04NpnhoqLLFqpSVrsNDZLr+6kohdGvM
9nLlj+jYMQQIpZCcS7HVwElNczeZ6ao29GyMmHcmV+sbrIvxITttL1j8eThFFWVr
D+fkJrQjxjG1ahXAwm9bNSgUjDccZqbLgfn0h1ZWtGBXdBEB7+4wbnEZVVZmO0kK
/k//hHZKqBkD1SsputVHiQc+VxxhxapB2wgaA89aoVT/Q4uiX8yt013F9VMG8mQ3
km4+WsCzsqIloUNWnc8vyz0bb13lAS8t+S3i91Nv5BDHfe3MCX6gTMYY8M+e/CPn
TuQxUp9CIRokWzXw6nT2UeWs0sZAAE4pI3QoNJCPV3AXwZUSqNeiHX/Q2SO5Id6c
zyHragD0XMyrt9y//2OeJv3Pjl4+aPkT9DM2H3XiWhvsNm3gkVif/xGPwbo//Tmm
4RBvgpQ8HZRm0wlZBw7z6RJtBztBwYclHcLEa1kTuMaOrwCGnF5YoFo+Qah0/DnS
NTzQqmPXjyWoDsd4KxKzN7RXGhtblCn5VAc2gO0eiwmfqQdgkS2xQuOQVLmqsNTe
uOVhTd7YApBHSMDwcb4kf/MWo/VBG9fXHIUKwW38E7/I7lwefh7JBjVGOJAQrxEs
l/YTesNFkaA7vF9tozAGqGyIceBS1Y3A35D77WGqrVQZTRDTP9IqTjAamaVDzmVz
azC6isi7BtbU1cAgQ0X/ABP4ZewaSHzpONpX1z4M03rOYxn1lNqHANaXBTmJQ4iL
dArZGhzdMaG9seexPC7fKuHO6qa+dEgkpE1Nsqi8uqKHQzARPr4hH/nGb0n81JAo
k/4vQc8C/Lpm7WQ/L16cSGlVHNEGexCAUEirYW05WpgnXRZDNGkCI+75Wu4phXrM
i3jAg0G3goP9aXpYnFLJ59S3Heqsgn97HPC7quyreBqsIUiTBzxDlFAPekIctf1r
jVA4YtzgEBrGpZT4GCDOKF6cXdBpfDlh63s8jYfTl1KMWQOSKsbpfeiSvTd1HTDF
D09hDfpuyg5yBkSGgjUDIjpL/dkCspo2qxuGdW/eTTO/h9fxmpYxTN0abJI46lv9
O1s1CuBQcCyp97/zmbncQbLIhPK9v7gcxd/dlNyUzsDP4hbkku8yCzT391zleSWj
GSrWiTYF0nYUJSh7crWFVRVOjdm+6QmHN27GY5dDgACUlk7CQzMIBlK2NAHsbAlD
uGeM3kvPN/n1o0n/yAzX+Yaq5MJVufJKx/upKxDjIQy+NHoisTqK5y2Jztk2Qeog
KRIL82va4fjJwYxFa6+j0noDFth9iE8ueU8xoC4Dm9CFkW/CNs5FG8zz9LpLSNDL
0ELkoL+IIIeGTTHP2jn1YHBvUfLqTKiTgWwEds9J188=
`protect END_PROTECTED
