`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gWPo6WF+0JvzcngGgybi5PBi2GzrBS7QgVqXh+AqwG9Sx69MfHQSngeiLDZeqNiv
gOVJxVpe12usCU5XOUF2jzCqAwu99vfgf+G5BtLNu6yRzBOX7jkpsyf+vTeRoFM+
TSbuve+/Yvn1OLCnpmRHcoCKlRAYG/qGmvdDqU56PM+uvJ0tOPgColH+m2b2VfBB
aCPyfhN55eh0NaqT3//MOvABVGMKNiY/hw9+fKssrFwYo2vworQf+es5YlwgY1za
SCnzUsTzIVJykSduUtOQPG37/aJ/eXUzytTBJyen1ctNypWEw3osH0EIpONe8dLy
B9Ph5NYJVHFj2Ju3qxI7ME/gqHi6aTQbWopFYwqVwMQJVnSPzr7HxOpcX/hUOcRP
ZPumNoo+r0yqOKdCujiB7ssEU4yz+QzvtAAh4UbHIqIsvGZ6qwgR+DkrzPrrbjNp
DqGPgy7r4+uw7APynf4G4GmS1OFm2KWQgcN3QIWnHxbXQF2M4wZdraOFR1UwmFMK
ioxoZTOCjF1gom2KKiOiohhsdAkI6Y38DgQfEOtXLFGPm6WVPjUKWj+xnN3AOlbv
Y7NtU6nmz8iXaMVu6DJ/jqK7ypbSJcO5qPNGPn8pqoI=
`protect END_PROTECTED
