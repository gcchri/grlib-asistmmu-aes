`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gE1/LMk5DXvkdUgNxgOsH3KBHfnyqg8wXDIpXrFGOrCatQK7LW9WNzJSSDqKkqxb
HesJeVFs5tzIB07cAkXA/7SFqorzUKMU8PFdnwrpb84h5LaDmeYLffkfuYSxiJ1l
wulW9LfUWKMwBQtzXn0fQYPeODT9EAT9jycyNhZjSsKEfeWfCjg0shmb+pauFIea
FXhEG7zYKBuQK+lsXjtWPeet9dBdziLTt/WTPqavk4qOoUH9pqfnv2UHuskiXfu0
iNGAve2Muzn3xDrkJmZjYDxCM0Z3DHbm6bisH4VDGXfbN63gpw6rsu1Z4rIoqR+C
oTpMRTKetOWBKwmRyLATlqBPN1mbzsrcTf+OV6m/JovOGYXDmPaAFqntxPVDpEs/
QEyEzO5lcfrNx/oYz5lD25fYDPvfWgEzZmEDYf9GK/hG5c9HsXmxsRc7HxMljQXB
gommoHpphByYrGRUR/AYHMYU+9Sshyop3fo+Pr9SdxQczdTt3iQexcdJo+r6l+h7
IxyMp3Aeve7WriYgfH89cLJ5PqKXcntdqSqisYpCnYiccz0Jh1E0DchxJGedGl2j
YAT/uOMY0oEv45xNpsd7/RjEN3w3wn+qeUacHzwj0VdBdK8M4vt6v3pNlEWJ5Hu/
d8A+tCuu3I+5XD6ZM4OWg0/Jt1bCkz5afkmcWPT7y+4TulY3qOSGCu753m5HXdnn
BWyQ/qaC5SYYEBplzc/UwbCbYPPZAMxcCBFGHQX9xfUdCxZc1P4ZKSCZOhEv+t/G
Uu4XMmz7RJPM4hhJbYqA6XILfOym+jRZNn99vaY4mhHtJQ2pC+ttGqDs+4RWThUN
T3pC0/4HWcbJUsSNXEbsFWR8YpxTYBuxk7mPaOBPTYd+N6tZAjhEV83y4ReMWiMO
ZPdBMsAOZDnz4MjedfsBD9bHIxV0hkZZ2utPP28O/AEgA2Gtyu9v9/Bi5oEOkJ/r
`protect END_PROTECTED
