`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
586qc4EoGmZgGyOTkiUY15pI4vYemaBp52nsIjpie3qYyxREC8KxHNFtEAEm55eX
ZHbEWOU9qB2JWtpo853uvlMwv+k2YQrGR24G7stCe2ib4xByTNJHZIzQ14az9sM5
EBl2BHah3WWqtoHAIBRbnOpTC4ngBlyyh22xt9dHTkB07GKksKzIx8RwzK+zHHhU
VaIXYjfq9K/fr2K2HFpjK8h4Eeyi2ntO2i/S58S2prqpnwAgT8LZC3I/HQOHNzD4
CsWJ954qTeGfLY+gcuorTNTLn0hAAO2A0yH7VK2JhFKU9KYN2O0McLSv5S8bNEOi
DZ7AMqpLa5KKKoY8N+vdumCdeeRbqlhCcI3KZz8yTYRhUtbL3NhStQKYVHvu4Q23
GCj5jG5oDirF1bzVhZzagnu4Xn1Mzu43U02saMzdTK/IiirjCkypDWKfEu4giNCb
Ki33e31g2qAD7Yj7JlYxjkTxFNBa7fnA9SmbVVsW96pANZnnng9URmfjmRT5phiY
bIIvVhkteGEXi/TtK3v0xlA94n+S0F/FPYHLaf91lOXfRNb11CBNqfhp/zKk+aap
owJHz4IS9CQsW2Xzt4W6lb7DyBUKIIMTGK92yFp2nFmX0WfClTPqlu2b2gliv6Kl
uGV1Gux7cq+GJwcnBwGJzL2vmKY+jNkO7eS29nYV8Gb971rz49Cgdx3fNfCiPG1F
iDw9OnlmirOxqp0WFUr/VFjke9YCL80yyf6hpPSurt71+TIBPMKaz1oA1kxxQK5/
r6S6n7efz6UObW6rm/mmYSbEEeflbpkXtwpBlNlQA70bCPu8/UxgIQtydA4BxpXF
sdpIsA1NySIJUqOs4Vge3kQ2S87b16oInc22qaSPm6SBXS5m7VaKoOTY86WPK0aF
pI0qWx9U3+0vHt4HuxflAa1GNXYwcNcgGiCiAYbriIbwvCBbtFYUeGNQjj4MhRml
ZmKPMpAa1WmNfb4+k89BD3brKmeMHw8oBvuWN4nXoYF4pxGl032w2Y84IHMDYn/H
TIMZuzNlt4k58KPAHXIzPGQA017sHsdgddsO6Jzb/TcRfXrOt1RbwYWHCHUM+66/
5n3afNgM9dbommii4eBpA9eTYqnH8txtPp/szGUtvovp5aKA7AYuVvmvl3ux8oZm
RockU+U0mpao6e7wbF17E0UhqzT/9vjsxXnFPVuCfJ05LXd1qOCG8tmpWdztl3Nc
zcmvRdlPRs9dMraRm3LufJIRD62998XELwgi2lAMWQmEwAi1SYk2WCLj4B43eCKJ
12DNQkNqrH0HmJt1vw5ISfkGQ3o93zCIOOBsg7KVgm0FIgybA7qgdU8ZBskfS1mm
30Sh1fKKihxEPQMsY7QJPqHudFND7+jedk3qw34PozsEFoq2l2SYWIq4ydmNbv2E
yzQ7LFSUP6gtU7kmJlxc58mnbzZhkv7vWxPLiAniQA7E5ikt0rp511HRwj7LlKHU
/E7NE6Ma7c3UdThH2KjHxEVrcFgf5o1qtVaKCgMsRANtGeLEgdPFTXxIuL7crJyr
kJf1TKNBh/cUiTNKzo7kWPJdvuTcbgL7bXdD0G3Tac7P+nqXSuXyqvcbkvdOPP02
GoD3qBj+qXIwdneYTCkQjFhpPNdyrqn5BEnNNISu4WwDxM3TE05mmS0NzInX5cyV
LpcyozMOjTc8eIiA5t8zf232A6Hx7bwBiVygaJhZ1f0mAN99wdM7cSKyQ5zLn20V
9WVSKEz3P0d89exT51JP9HP8ZwF/ZBUh/1pIRrvhQt7PHm9ME7QGIbmW68YlHx24
cPkkcNKvVokj1qoCV2WBK4QN+KO2ybQ/WHpzoSA3j3U1oMQOxtqi0euG1Ch4s4ya
zCu5S8QlbEiktgZNfNRT6Sr8csimrGf5/bVxgrN1PAE7pJAQe5/jqbpmtsK7QGRZ
8tBInaKo7Ra5s9Cqdp/nmrnh+HUoCUuFG0a7RYqnkQ8feH0ikZrD2aLYsbDuaduS
4jFP2FHTl4yum4Hd2sDzlWEiExJbqfPESbutcdSYAkuwMtlEGbNuhCUQ97LYQ0cj
PB147SC+J2PvkDC5ygrMAHH/CBaZfQtmBwQJODGS56MgAgnb3ruQhgTF7YoSBYLN
fyNDBg9SIxYX9lcOPPv9/qI/4S6/Is8Mg7tNcGaBe5pFp7FRrsQmV+LsLP1BS4zB
yJ5wDsVv+36hSv/kOwHgWmuICz8aNxLV3q5l/eFCHRv4avaz/X1qiKFZrCdlRfON
nxPbLjFKr5iMQQRZ4zHW/w+iOc7mBfWGyZchrjgWXCkKcbMBnnKhxeY7HnotnLbz
5vzE0NPsFzfzA3C1WzNh2vmNAqbTnzS+VBe1pVkQCot9jiQ/gOIL6KefFTcpm3FE
FWsFYwD3K0ar1NyThN3T8G3T1TtU7+6qjm8q2/zSqvaMEkNYzeg0cnMd0mApQM0b
eCKz1+do2RmEAj5GE53TJAa/tCP4eS1aEWt1XMWoA1KKe9aVI9nPhtUyc4Ee5tXV
LeV3cKR3LeGgI0Rj4HQ1zI4OMeK5qs6C2Xxs7EH7hyyiPNObucdxSUgP1h8hNY3K
3T9iZ5A5kju60Bs0CwfEa1tHnSBitlUNtZo93y3BfiAm5caJhFUwcsqwXjSoF5h0
mdyUdKF7ETmTgfA4IaEQR/FCH01VXWoQ8VWbzGo0fclprDESk9mhc1kSt20cpANP
RzQyOpEmhN1NbonSQIJgDtanzobuk0JdwBmgHOTdWIj+XO7AltcB5FlTYGmf5dC4
pWp7HG6z6599wCaR36Bai7WUY4Bq6RHNxtq+zNF2SuLiBpgrcUGfWURIiEllNSXp
LyfPKdDSjp+Y7F3m+JbCWclgq2kPjjGGbWnrWDIbcZ2Ixw4d5k+CdRx9ekRrapIY
ikfQJkxBxYXjQZZyXZrAAzT/0Fmu/8jXkCwNzNS8vTXn6zyo75FPgyttf+ONocN2
96i3zeUJPpFB14wKh3+GmEriBiWqn0H/O/Hwf8GkqhJ6RwQ9bvptDPpiL8hDNqCQ
1tXRcvcMDLGhZOI+wlnuzDN1EAuhokuslGh+zuGFWmtHFgtWRRjyD2s4LQsuGRkl
ew7Php8kCmqzXPcYKUfB8hWdRvBmBy5Hk7tBwFSvH2IRt8Yx6nwgrwEpgIgHUPvr
IHZ+9wuYNaKA55RMqWiD9JQ4tLYqbi3DEeYKDOxitX5BDQbLcddWWwUAqZ3d3V0R
j9K+bt+ekNocr7/Vbi1d+5kNezekgK8ymRZUnjB9ZTNtHHPcLcUleiRHDoxNWDym
GrrFluKmrpvBP6CWtlNnCKRd/9FtAA+4R9s1gstB6/CKUawfMoje+iMPjG+JaPKz
8iCgdRcV18Qcs9gXByZ/vecOgP2yjwthTbZdF//Z8JuLW8/Iz+cTGvLA1dCDJ5ZT
`protect END_PROTECTED
