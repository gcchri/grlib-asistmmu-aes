`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JDvIk84QXTK2Aa3pQuntG//JrRusEdSC5FIYjZTxrOxRakAKcF4cRAI4xKFwXM/t
vyhe4n4pcLWz4zbwBaXL1SrbM7XK/nol5zWgCWtaav7plBlUM75syB2mjiOlEPLq
H0KscdO2jq7lzLKUKhDaM0pPf8LTNREiJYHEF6zZ0tIKUfVSSzkYuY8ZcH7iwNGY
U/UNH3n6EEkjCbvCJkTWuMYQsDWudskpGCEUD3WPzu1qt5tkLUFA1u/nePaVHqD0
SMbsYiMiKhcGOPHIiMGpUw==
`protect END_PROTECTED
