`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NGcL9AQ01qS/vhnLD8C6YTDKd8xcOMASARHr/nGNW9rJNHFl8gr3uwinMYYvQ1Uk
AZ7PFgqr+RzlFYHppYaPNF/p01kcC5V70U+sKVOYSKPZ7nuQdN5oR8g9L8awSV0b
pQKs640pPGfTd7lbYKx1FOKtfztrLl1ULJBZvu1W4dPZ+79uynn/j+CwLGWlCQkl
exDiBuxfXaelQCfa0g1pE5mAaMGeg9eIH67ZWZ1EcwldNjTerteXBa55w57UYKd9
7KFvgTCPyvRLVykmnkVmzTQgSEXafg8ypHk0xyO29KmcoxySoLSwBMgf0YLP5S7r
osX7tFoKNBgsQ79SJiDx8QbpPKB7G01SgrkDn9/nPL8LAOxYWPOYnzePa7jjufq8
4uv7XHYFKBdudCR52vV3Bo9zpqxBAzndgA/tB24j0AKpjW3qxbKD4rYln8vONfkA
`protect END_PROTECTED
