`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9JL1OLekUzTTDy33nXaxB6/7svOLLH391x7E6+VOoXH/cYz+iJ0uEjULwxamZve9
juV+8tAN9TMs32DwQj/ixyrJOMJodL7amZyVUdLfb6Xjuk/Wp1Vplvf3LREAdDMk
vGRPwyeQeIcXSlTe9Ktf5kzGrd770binVG4tj6I4XjYO74J9l5N1puS6j+TuGNXs
8Wkq+MZNM7S5pSDtMMUTHFYv/JW1eqqpzqpX6p05hTtVMhTVW0U04dS9vS+BSFZl
5Ep5yizGUlkYVwM+Kf9iyonV53DyT33LtPxDoun3AjIV2mZvMfd6tFA9t1EugmvV
PQqs55QQqGRlIHIwnZ6Xk4VAfDD5I2foI/JpSD0zrA4=
`protect END_PROTECTED
