`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IpZb4KfNkqr+k2wqXd3tVQLox7VtZVLwFNqs/mrf8hmhJtGcCOo8ynmSpO2TFgZc
+VPhTqfZpQObuS2G+Wsyj3zDx+gLIgll4xxDBKzbXo7wmBIOt3sJ3g3LSNFDp+QD
DCpiKhr27Jdf2VyR12jpS0Gn6HAmapgiAeB8fZ56KdAnXysT2ICTK93srBClObbH
zOcuR5lKcqbgMwURrahNDaugcevSYQLvvdIY8il6E64ZX8guV0wJPuVJ/Gnt67tP
olCfmidnklZFVCtSEkQby7tooIuz/DM4QDa8WA4KSPrAX+UBn2AhZ138oeK5YdMe
gIOxCjkScIDQPXeAC9iTSTZykVtWEaptlUOTuyrL5HtsXOyedwCP91UoaioMyYMX
pVzaPpya1jSgRX0gPqMdllOo7/TtWzpAjnAfD9sWYjQwSNHuIpYZZJqsfP/pa6KY
xyvl0qEsHwUMsHN4EDHUgaRmhCFlzkqn1ZeQFpNAbvnIrqXmhU9/vqY4uX4Vv1XQ
LfH0u83qzskNG6ldHoh96QbR9LMsBERz+89Elt+hZqceWpGq0Hgq4f3iikI4y0Xh
MiFhUQsz9piv4jzpL9OdZhRd3luUJUgtTdCJxfUMmH7oI0PngaDR9GTriXM+IzaZ
lr8zhaqkKCgOwqaPbCdRoDhMsWDyAnARc/gRXrSsbZJAoQsAIi0nW4AUN6nz7+Dn
aZ0f83iH0EKq2L4fUrTH8ze3WItWGUKWLaC+2BkJpiMybLcT9bAeuieFk9fYneLz
MAY7C8uWowNsgeP1CfH0gMjISHbCEc44jgdoIsudp8g3AUM5/fIYSZY6GpFyi4qJ
eG20+RVH2KTyUFR7Vel4WwvitkDzJUBVLuvjBlz7zuqKC9nxwIhtIwwwzj+7dOYY
Wym67msIjN5mut1wKledZ+lO/v5elhW3uRVp45lUzv0dmACC1cTQVUiuo17kXNSa
FsCZGCvgvYGjBH0CUqTkIYfU7jrMMz1+96s9ANdDb0DY1Ok+tTfTlfYV8Gp3T2NM
9hiHlZ4Otq8MGUKb4p6tCg==
`protect END_PROTECTED
