`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aoyCKlSaCMNW7xco8nRZ4+42azR7kDMmiTkDsdX2TJfN1h5e8KvS6HwnjWXWMn7y
kSWw2XZRMUu1++mBTVx9eTULjwDuZz5nXP1wzu0AwHBMJJLRT0jrlVICLtq6Zk0Y
Y9GoQMRZFjqcD4H4z7yyfI4rKBOZRL36EELse/IwOFVcUWWEAE3SStWAsZJqCqgw
wnuNoxYMgrH410riOur7fhlumVaeZp1j15jLFnPVXgeZAU5VVgx8+X8K1/nnmxaX
Mt+cGYnDfUUIf7a62h19tkA963Af4yN3lBVZPqW1InFhXeYcsjvFfPQIkd+fUweV
NJ+nfEhGE7RmEE9qUPAC8cvtb5U6cR8ROWwPrMLYaL5H4dLzBAFQM2Lwo4My3SaZ
uPgZEuS7Z71tTQRef6Vp7aBoJoFLGYg1bLb5vVg2A6mPQsF06zwPAuWUyQjtAm+q
rKuCtfR7VNKqjeHGHE+Y2/1BFPSCR2ecPNqPj/HLG2irNcVAi4rqfxDtorU0zaLf
5o4CI7N/NJhBwtshwZp2jYBsb8tdk+WyWZ9Ky4Crv1IZSueBnVgLcT7KRJY6XQCq
gcQUOgVRvs3IBp1gXS0QVdiH4HEwI/icHfX6hw0g1saP7lwHASI1h6S7eWseJL+s
in9ihnYjmMkphokZSd72JVvbZzC4Z2V6MRvgvhbGZnY9YdoP3iCk0F6KRcKbFgtb
7aR8Zza3fYFgv8qCSLL4/NyJJXNPOOhdk/V0jY1CU6k5oUk16q35r6qB1wn+R82u
5sguwQV7z1oFpPwcOaWIvT94efRNxsxBh+IYEycXW0bJM4FLYvBijqsw0+aMLIVo
iToKSiEPxziqfyF1KOvL6Blm3kn/DMM/mRfW0mP4mTMVXReROZ7t/LK2VeYjVfG6
gC4KSLlggPR3dMPsulTFGrXya6+rCa7EhTAh3aSRulJ0c1ZWGCSFYmkhU5/NkfZP
KT9PmuPMQu9xGMKR8uBsz4bRk+0s2xXEg5pzj4fc39pqi+8tsTEkxK/lRELiKyE8
J3OdUjJDsaaKHIfuMEXap+xj9nq8aJ2B+y+qVL45YWeytsIpwqczCVFwqki0LUhY
AUWA0WEA5Noe3RMTU+23xNf+CqbhVleTss43mMrTFFnafyWE0a/kKKosdG7fJWXa
2dkBg7ILz3ka6dER2mIhBIp4nbbbQqY3DBlAsvVyAy3SqWIWOdK2/IXK8kCEc/f4
zMeMtMegWt6W0tQuQhj3+wQF3WAn+VW1nhX1XgdyMTN9s5v0rkB39IFAK0CHu2HY
LcZlQicPx2kvFz9Gd005wq9fLQiBnWugyCbWtR5p0gBJzway0cwoUFD29fP/BIeT
zpxPkTEXYP/6Ej1NBmza1V1Wgz+TMNrZK8IQ6n2QLCJaOkBXjhoxs+lZ3qBRlUjS
CKj8+WnasVINKkVQ0hn72kDO9wBEHEhp8Gs6GQrAcXLcZuNqRfwBsC77431lLR/c
tRTRYYQiWhnsJtQj912b0dNZs/l54rI5GZ7lArW7gNv36dSB5UQsZCRKqYGJpY10
fSdRiah1gQselOwYciy6iLQGuTZ9eORJBrMPH+fioPNa+goPF0qnt4we9kMMZvzT
/yQ8KA+iVrHBBVUBFoVhKRp/jcpwgb3UPXhwW91/3zuF9lfa9PCpA0ausCYCYaq8
tEZ5aHeRbmQH0bhBi4R4YeuX4uPVJrhhKAktUuOmVSm5G8CR3EhBAOe9JfsU31T5
GcEFSvGuvXI45+WL1NE9/YSvIH3Bg4Uyg48EnXh+CXqx/8Luia6nmeNpBpCc9PYY
wE0FqB/NmHon+e78OTSdei6iaDZrjxOvKvS7UpXrLxz86z8E/2DPowd8Xb3YvZRb
FxuiswFD+TLObT+dR2CA7o0v/45FmgYvvhMOELsObDz6zSfMgwIQyJFgTy3rtIJf
BCrQuy6Zwg/jauqZFgS6b31Yuz824NTmyZOOvkPXmcuFZo4MnUQ6ALdoHQ405FoU
yppYa+uzfiWiUvmEvdIA8E6fPuUq6Jdv+PQxOotM72TNxeBwxahaLf4jWQ84M9FE
HLP94cObu+FjPgzkVN9HOOSQFL/NXkr4c5sG10Xx11fdB74SaYK20EXQseah2Way
q7MCDFYH/tEcFtMWRm+erT8nL/NI09BWptr8vAdnGQgVemr0HAvTLXdy4qq7oPon
0k/8/+l7MtTS4LHqRk7HCc2s61DnylY3pZVMELHyIzsF7jzZF7+5j/S4irrYsfkh
4gyeT0/cPh4AT5sEPaf7wc4hR0jRCiH4pLNOK/WtPz3T9et9HwLTQfpZHoTzlrP2
yptXSvz9d/hTJmDWKZRmPSHziXP0Fmvox4Il2zIQIDnYLiK2ZQoKkO9RGvxu1mlh
3mhlfMrxD9M1I27ANsejHeqs/hOfNa2MWNSqiI7+hG6nqarmdkcd6rP3wBd37W0U
aJSAQr44uyHwiVrRckPddXRM37PHUm476XR4A4kxRHDUoLiNCyq25RlPjxOnSeJR
5yB6ZiZKIRevnAC0GjJ1gA7d0XObxsqHEcbkukd62e4eunb/f58/6vL63A8LKqOM
miHoCdjU019rCZY+Nh6LT1lRX29DEY/kuGUSnYOXepeCKs3E+3+hm/C+1wEl4Cm3
k9YuwjymS5RrdFqj6pXw3KDJI0qcuvSixx25kKz1+BXMGIEO/09gWLr+0f9noHHM
ppDk+wS4JVvS41bvXyNH49PNOp8chMybqw37Och3Sa7tnteW4pEYwja9u56PEgzg
cyLElZMUXdSniLemgHGaM9e3vZoO/Se39R0xdvQi4TfegeWvD0/6OdowMKvin18t
ZRaFqO2+HXOycJ8kGO690jusvZvuSLJPqZKMcQzxtJFc+YtnIo8zYVM1hA71aGkY
OWIXZQReq8S29GntQOuZjHAajDDJYcwOCZkrEIac83jU5vWAh4YzH671Hb7/UFnY
kmCz8pqBeXQmPy1CLsJqrPmTeqZBrXIYjyrAHq8+O1CwK2KzqhxBlb71MYTaeU43
WNPcmXFCEcx2lcXXZ+6V/DGN6OzbiwLtnksWOkS9l24vJVwhAeguK6rwwn+NtrWX
5InoouUAQU6oqKOhX9IoYz2RD33hKI8oGnaEGStBayI/iUyp1bUCfPauEvsRkgfS
XfUuWIib5vy5XKj5kvONJFs4LZIfH9o2cxqa1wZJYaHTMmnj0njmzEpOsC83JQ1x
i7CiFQu+hage0ZVZLhssDsDyOa+cBjnG6JKE33dqmZG3q8ne/F7gVhsuvZViE9mE
UQcf0CFIueAju8xvI2f+Qo3VvE9zN2bVZyXZl5Tc199wP8E31VvceMCVUkdic7wo
J6Q+dBQ/gP/vSxqyWAYNRaDnTNvk0IInkn9atqzT0nbay3DrWKwrnDhXWvVv+sbm
acLymCAIgMWm8aNYlDFf0BzLuRPTRUWK7EmHZHZOt9bPlJ5Fjysls8LpLdANT++m
bIsyx7PW1cfV2BH3KbtLiCjxcwlKlzQlhs+bedBMOEuo06KNHurwoaq57Se/wG50
1Yuga7p62Cb2s7KRf/uLJl9tmFCVtt99HW5/pwb//L/UYay62jvVsG++wJT+2Baj
jqaeDT0px+paclTh2XAzFvQ46OkGO3JrEGxzr7OTq604MixqJzPxWKFFKJiEgwR5
3BjzqCb7FtQz8psvCfS921jumBOLIaMSSc7tXNJ8VfjVslLTD0er2yH6DD8edUr7
WTgL42Ix733IxBVluK8p8CXrTiS9nt4qUS+3lVwRTICTFiZmklnrTmodjroPX1pD
6TsnHPcvi1YWJ1Z1gNYA9nW/IWDJMsnS86Qd+OahWbh8keElBqkwMgkj8HG38RE6
KbYSwxqhxUG9JqJoCC7w1AuGaEZ2HfqFCHFm5MkRwFv5stIP+2b3f8FBtP466U7s
W/CuxFCcpypxeUDeJKaVab0i3x+HIojhhSJquzNCdErUepoodr506TDSaq5FoTW6
LTa6F7VFgOUY6ELO4e+My9vYg5hKGSxdEfBpQ6ZI9jm0QpN7w9g1x9ki1WhF8jL6
Tu7/9pehyKVTmgQdPC9Pfgp5g4+IgVr0NmjGh3eF9EHdaAplpNPrkkuYUt4MKfv+
H8AfwmAFiknNUiuscQr081rsCdm48WflVpwu4fPrwn+1cwr7uUgJNhv2pf4YM0oT
UUGjEGihk2LjZ/kTQhoV5f9U7tj9S1u/HMvVoNcCH6ib9TfNimIaxUpVpPd3RyxF
UgGolu6lAf5NmihxiNyteptLOEeqRvhr1cNwVfH4i3cexP7O+qUfJY03b/RD+D8H
Xpto5iexh+DIGX9dn0ZK5pd0ZLHBlJO5ZX+NHjqyS0jJz04fpPwkzFjeFdC0tqSc
YYk7AAzLINm7VpMRHn6jIJM0WJItFlBjydNMKhgKfotTB1gdJnavez+wQbAVyiAb
AbuRkBZB4T0z7gDP9ztF7GjBYUpvAzhFzqpJytUNsgKHiEVl5HwR/m1352xgu0BV
Aw9DVdQpGFsXXOMfSdc5xofI4ftOF2lgsQjVAfwWTmVtrtOktEhYBv4r42JqZGn7
WqPhviLbPomW1tVXzHpd3SefsEYYqwjqpPAg6oWBaSQSEi1tBdZt+mHKKwtF0yY0
f7cnqRjGIkRD8LRVToOMHgYyi3P2aeY57q/RiXPOJ5FQsgfffzzYHzka8cO4BMSW
z/o75/w3xYF8XkPLNctIjlQFLBc5mv6G6F5elWgjJRTMo8jNMA0vjLeyrDyaoWla
nlbtajIoOn99004v3KO10YFOjtdktk1Xs/5VZQNS9e4W36FwB0pvUGwfMbGVqL2V
DbDwmSkaclOuAqMGmHBhdqNWshl4MjQb4frU8MG1S88LaJvhlZIQfatIfMjwZAD1
Wjyph0nHOkd0d16sAYLBL3sE1baqtZUmQBSduEq/NMBw9C+Zs5IHgyT1Al17u6yq
/E4v6FMsDGNrK/Ji75iQrKCPte/4Lp0Kp15hx+vWaV/9zISG0hC7o95m02O9WWjs
a+bmUilEP1HC7tvokJRd1u1K07Z3psICIYgZIT+Fr0cy0fRITcZ3N8AMuJgpO4Jk
xeio2Y3e2dfOGnjHzwYxknHSryHjHSu2YNHNBn+ffHvN8vL0tOawh+SeVLwpTqN8
2OmXFmwc2qDfhTUeY8tilePYq5DeGgMlRJEyZdII6PiPgqONYauANR5Fc7c3R6uG
rZD3xP/474qKAqwoQiljw/1CoMZKkXi9ZTIcIzuUqmi6Vv4yeu/QIduMb0S0Q6GS
7w/L+YYdkQH7jClfI90FoeSuYAwc+9qeW3A1ItiBO4QjzkRWcLgSTnbJDE9rChx/
KIVIwQxZPAXwpEauNYpv59DEqgcUuoTL6NVJ/cDCLcnTkDbVrD6xBU+L/Akcl1Br
TBdKjmRVQEWY8OS9s6PGN0n6Va1gRaPF9pzkwIp9aBvDTQDtpzvSYBrcQBJdjcaK
+1tV3HsoMHGdnytwhOtLQa+apEJmtBgs/0D3C61dO3F+bxWcH9INGqJmOULR5nJs
5PZP7iSASooh2bqjvFKWvW/oS3yx+k2uynoqdG3QGLpR8+Z5aIjQupBP3X1O7f++
iX2y6T5UlAni50FUKI55+DGjMj5SsrQE7xMaRR/Docj+LlEz4ggsf7xvMksEMZcu
gAXE4fMDhBTqwlSpi2ax98wZ1fRjM2TUoB1BlJga3zSzrXs0fwCt8SR6cMzcAF/2
6HV/Rd5E9TJUnJQRisGCYzm9DetD8gaOHSNkAxBfKo8dezqlsU+v5p0ZR4pvBZYW
8qschIxp+F9+8vJuCgWF9SfZE8018qNlRnM+iQPkaKhVxiesq4qS/wVaWbWgSo8B
f5mkONUP5mdDJMxs+RKrshaQbLb9RRQDyHGL+K8oOt4=
`protect END_PROTECTED
