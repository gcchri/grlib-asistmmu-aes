`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8/Dubn2//KFtMtlzBC4AMyXyk9H4J0gl/7fQZd0Jm8eh9SXhNunovJ9gMsI2AFG1
Qcc3Y19FSReYlELmXGPhCtuGcqdKPObdzFmvBiPwMacWnyu6hcaflDu2oqR4ppwB
yJ35bz9iaIyoDNeTC8YAEzYs5elAZ/X2drhHtlnWFZYxHgv/0VCoCAbNUYLGyOjA
eiaAdJXarNDM6kjbFRC4hy+3KlnU+FrfYiVMj3tFBEKDikph6UgjDXO3AZwPLuY8
SuIrsPFn8b/Eu9hPFAGohVXY2Va9az3McyuEkeMYO6Y6UN+p5ubbTgTFz9jFYokb
cUxd8okgOdt+uJ963kleW4wYBNSLqAM6gg6OJgiGVKjl9ISc/6NuDCwNfAhlyIVk
+H3HVDI3eQjI7shfnHHwGDLwhHcQAcrzwXydqJSfGKNRj+oa9RDfB8pQcrNtwdh9
/uEquzMrcFfU2SHNOlas5ZVW/ZBLKDaypI5CESJBrlgBX6VPRh7bVVLsbRlAxNCa
MW5Ek0hWE15KiYrvdkesfq7ahP3sqk+N9MyWaTSYExIi2k9xtsQbQfceFP3cLj2J
H3qxnMlPd1TXM7cbRM2XCr2lvNWhj6TmZAsFtY2cDgcTcholr1dUzWqUN1zM9BJM
grjclhZJ9+M1OiPNIPqmlWR6Xepup2HKhXziuJjzPQCecOGcfhmHP0OpL9oR3glg
c+NGB1afpvglPLlmubYmg9kcxNtllPvKENxo8kLsShkbI35ATTExC7a1LcWD1c22
dJ9xm1jLIv0ETO2S43LE7dTerU2AhyBuETyWZgBjUC79HgvUPVHd9c0lnXofSV6n
KPgraLHXCYfWKLNrXKKt9wE8U41wsiHm3hG2Zvc+FKLQyNS/zT+8e4cX+I4f8fC7
Sfr6xDI4qjngNS7ONz6F0zovaxX26VmZnlag5yVc8aXVTGAEEpAKFOudbFij+Cv1
1dDsUbZCmLi1PYR3OGCTur8r6Qyn4YWChuK5p/v7HLw80Dhi1MDtBtvktcqZOOUk
NoFEkOJt7wjs3rFa3Xl7+jwmxt0RJOf6h7osE7fjjIQZvyl05HK1idKRc628QjvO
XgUZ12idp8FLi35dOYw50H42ZqWsg4shsDO+Yw8WPIIGc9X6toIrgMxOxfCC2yKJ
HAHlQoSZ6wCxq+LgI63cDQulrA3mdmZrtAvMwJxE0ZW5YT+TGiQFN7JbaPqbghAE
GNreUiFxDdRKjK2rQYLlrafzRByIG7huPUtnqgjFX+8l3jZa7a58PwYJAKyiNPgG
9IgU8BGbi+vhK5CcUhnUxmjwitrXWe2p9/AdeHTddiQtP4ebVlUAxgoL+87ZmmJC
HfbM4uI1moSyqUvJ+0o3smjjlm5QdGQRMGaAKFN+pBn91L/A2sftvLsKUFY+ikid
VAV1xmDi7eUwD7nLznfmPDURaO1N3aezqV/9dBF5tb1JgSCWh8MS+SXRmXCZkEAg
dE4QC2Yec9cajNQWvmCg0mspcfgUEkDmxbf7+UUBzJyj8SAwQtLEFE68fgwHnQFN
7WrE5LRGUD3SMxbJwj4PjbdKeRkwS9a2h+VxRp2PRaQgs+Y4X89YyMv7/MiEjgNJ
ItnYTbFhdKLQwNR/acXehZNve5HVfGguU5qxRyQOn0WdLjCJgDvpzBiLjwuwcpOF
K5Su9sIqKvhLrsTf1+fAUCAz89tqQYeV7DKaAm9mnjYcgsC60/3cAE92xi68Gk9H
8Ab4/OXRrfPL2iSjtAKiZhQsl6/cAtylwnHXTZt6nG9vrCvAz0aB/2gezv34husa
pD3g6u33g0oSr/hZS6rPPqmmlCXb6lx+rJpGhUbdyKBuWOPcsOMGOY6tCnUp5cLQ
biWRQUV+wTqBZVbnjs5j3X6netSHQDvrgXk3XsHHCFNwMThJX48HMolVaySbv0Bp
eiLh7aOR8n9y3yalG36tqfUqOm4G8RflEWh2xiTk09vOgnFMG1wrUGxWWV9c1xsJ
Io8YWLIX+k6ZREPQdr4FUMCiBWdeqjs42R5IIwfTBsgLTf93mfVcccgB52bVUw2C
uWEJSv5IbpwLO4pY5E/O4U4pNYG3QaA+iiAJ6XQ7UKfXecIF74R/WWFZ5+WqT7/j
33yn4+yMsJlgicxCNivTX/rb39QUjj16CcbCtA0HkOdFV9PmQogChqAvip6H3bL5
Q1bN6qPnC7qaIsYXxr/3o02M3NB81grpnc2WlyqKqPp6VtHqsWiI4Gx6Oa0a6Ibz
hBtIbgRJtXOD2lZgTrJjRwHW/PtwM8NOSH6W1ttdBDuAje7+LJf2txD/qqCZ6U0Q
EFXbrHO62IwYMSpW65HrSXk189ti2CqSjS2O9p+3aa5naqr4iSYrHkI8nkgS0lFA
jF7MazRh/Gm+j6I9X0U3Lt27sZUcGl97MgqZEU2W8aDSG1GEuO8D8nzkWfbhF3tV
lWITo4+w2bDpAuvedN/CjIxv71rkFqn6i5G6hyNnB2kaWpoyU5MdCglz9KkDHwgc
fWX1aI/vA54ilPv/FhoPYj6RpL2QUgFg7yhB8DNbs2LVtsKhdsrcpNqL30GcJXgz
7s1gaNYHsTQGsuRcJe5uVQo/yvnfMKzsWW38/MCNYiQF/ret6bcvSF/8RrshJ6aU
vZm2D2C7fkmxusQVD1S1emGch2duqHPkGNbDVnSEoqQ5pK+r2rBpJ3Ccc1Aose+S
CF+e8jPSyJTMfPlqoRw+mKtafCM4n/HRRq/UdC7+O0JltCysxAluVn4gi1q8op9Q
l5PZUFi71OOKUNSXY/cDBjacZOhoxWovqllQDEtlNdE0fkukjO+26MyIfn30SOR5
2YR+MTQOhdU5NDasLvFRErUkPJ80PCTMDOia26ZRHNuX3H7EpJiNkRyC9FgTH+aC
Hq8bXG0xDgWqtoNitvvdqtPEu8bxeDKpnRnw/qn46ZD1gi/+ay+gwTfw5Zrc7kHX
tCG1dbbBvQdw9NNz54nMEqoLvOWSpcZ8YaDDuRSVwJtM62yUoiF/qGjxGio0bJW/
jPgIcPd1RT5mqtRy3isDsfnn/zj4XQmATqxX3+hkwKANxtaSubApeoK8E9zjlmK9
EeZlg7QIoNDsm4q3Y2wHSgHzaNum0krjnRFTgB2rca20tRuNVH04j3ob5rx4Ta11
HXc8WrU+RNSN2w20+/2lacTFb1r6czLGNem63ZEM4XW1ekYfw7qYEJCF50uzuSV0
iJxWGHshQo5QGzAo61RE69J6Qrr+97giPWbyYSZIyt7hbYoi6EMHLkIBHsyGmtXW
tBfhhpAk0NlxgMC5Gp8Y/IuC4QPMAmlTm+bOC4y5o7wIgatjVn+ik4ITPPVIVZwg
78Cp3IPUO4Qc9eZBbc0SlMpfSowDStJefRHBxFVuEI4zgCk+h3VR4VDqZvqRu5Xb
zppvqhWHkkLYF+9WjLa/UNHstQNQsddYtIwisovOGHypv0kC/MSMS8LnsuoVwYqj
4lDw5B3IQFzgGcCFnr26E5aBfbPvLzB/Cjnc2eqZkJUQts1OuUm9nEYrB5cqy8gA
rfbxFeMN8ROYDIKXMvNz+AgPcnip2eie5K0JgCCF6/Ir6aBioPRUBL3L87cMx1Df
BWVMofuebti7CLghyrxRgsHZKf3nPIQ2VwU6m9ns+cObx/tbuq7x6fGDO8U3O4nM
aILI/tEQyYQPZh5KVm3/lqCghifYVu6gqVWoe1+bcA3xYAbUxs+mqTmxH0KQj1xV
ac8Zc3WQ4WK9ZCu/rRxLnapHtv0SYgy51dZK9Vc7TYBgzqR64bIGKYcO6GkxK5XK
zcSw+zJd4xJ/bFzyBBTgLVpWcHWUkqmtlfbkyQ1Pvvdfd6RQ1oXRRygrwZYaLuY/
rjJg2u0/laVydx4W6NAUyIM/fxy4wTPSkUenMu5gxxBS3vZramcmKQ0Z0JRkeKNm
KZyFFxgxHeLJ2K6oJ7kpaZgLlHupdbecxMQA0o+s26sKFQhhv+A86l0PuASsIXG7
ffRUxNR+EDyRdl+kufN/ac3PSKvgymhSX45HH1JvmVWA+CEt0Ud6rtRy8+ncqOsz
7bF+Bpej5Gqvx0sYxdLrgYRDpYmXUOMEK7nked9+O2VPP1r+gQ855alfDC1Rygu4
OCcnVxt1fuXsB7QmuhsU0LFX1nynQZxy2UTlOmAITV7uA27oBgeEWoAL4wNuPfv/
kAS5xIWLosrbBnqzg2sU0ICvrQcxFogjWshZk9pQwzLHva7UgdNlmeRKHEVOXZSZ
6DDRvT5lRtnpRDWF276LCgtftmfV4xfPz2PSgGxbcuDNywilbofmXPdvaoqUgSTe
e7Azh1Y4rU2w/rg1uJ/2W+QStGsgN3l1Z2VganEdTngcOUzcJXyx3KQbVRQuo1Vd
E8DVQmD2Nu3nZXv9PQkYgnkfNyzsdkHQe11DYnfObTwjb4tJQuX2G8w/Whz2CCAi
nCt6Fz0JnzmpCiNAaCL4MRWt+l3+rFVDyhj5j9XAMpmyov8ilTGRrDrNYyhuUUIK
PPO5Rpr1Ox4rkna1rz2Xp9Z8g9R8thMsW6ljeo8droyGF5zDbptkd+qM0q1a7gw7
KOSi61kU2deR+UTQSM1va+5xmJ+uyqWHlrTWDqiXRh60zG3X4QLahQSKJssnlvR7
HI/hStMj+V5bpBQEZ50K8JomG9OZJFWJnyxTsfxspk3Veh0AQ5MAyElZScwdVE2y
65a9/qU6LRtEkDf1Djx0H0yKmFA+m1C76ppzxcFgcQQtPFzSaj9REjxsaEvh2LFU
jL5OmdB9guUOnP4nSYWGECcgaNUYiY8wnRzvqlZGO8qULY/ctNXey5lOfwUYJFh7
clnm1qHNgiA6qiAzZmnoTAZp46cvp7kxW64aRgqgVbcHWe7JJv4Q7NO5HAsdbu+9
FubxnUdBV9t3BSo88fTOWfNx6471/LqXo0SBB4bdrpyS+A9lVClxBH+1CcBoJuBC
7n7o9c8DSPoEfpoVb831R/7xhZIASh/8xyYKrd5KzbGYCTUraxQD9+9xW1YucB1C
rlyU9j9j9rTXBvcdETaZakKCo2OagCkz8E6RWZlS7VHsv4JSq6TIjZy27cmB6A1c
T4UJ2PptJ9Zh7+8VUSF+5hVWuyKZErb0U4vhy11WDSrRlvNFgeRHZ3weSYMJsqmZ
mYShoAzR556UbRioRlh4qveobUwXvVJPdS/9gHbz14jqfIjkXOC33P8eyZMx8pKy
f88xR4EZJtpilQRpklwQ6xqI/nN2wcQ8HDHM3almzwXzhRkqPuepdssY1m5L69px
57PKj8bdrN/IfkIE2yvERvExcyCFHrCA3Aa6W4FI/tm9n0Z6PsRCyqauK/QL7Ra1
NkIftlQbkwPjWqBdU2KL+8sGOMbIT6aR/uWi1z7q3fUnctgRynm9wukXe+dfWej2
u45zc+sY/y0DpqMAuv2NiBKZ38lOuVZSckdmIV3ftuvSsvhFRERVK5jyC0nBdX0m
8ehBojR6sfTLpns7Eo8R9xRSQF668weLuPMmMseFaDSS4Ui32r09RMX8W8HUy/CC
/N9jIrlrsTV8QFOYRCxFo2EY6HsLCfxpKGM6XNKbqmCIGRtG1VEQkaK4smWppp5V
7SLAOJD54E0nj7pHek7eD5dKzLc+G2/aYNy6wHW64X28/Ibj63Su6dzQrVpr0/UQ
v4pHq2pj2XrdRvlJV2UFXWOQ9uiET93XJp+vsuYvrldgYuc6x/vIpJtFGY4QiAPV
lXrIfsPKTG7zDrESp808f10937mFGPnd+XhcNz+fGXc7Bs4UwfJWrC1Wx9glqLK2
4cZ+3usqBJGVkWh+Mnh0J7+E+493NRSbhF8o2Zld71yDWH/dEf4ZSbAoZB5Mqqaz
buoVpJQOF/8+MjiitVpyPBHDP0Q0TNsEEv40HJU7M1490WK8F0+FQWReVNr3kONN
gB59v9Kem8IHsGjYUV6GMgTke4lkSUdJFIf7/d9x6FYf0ApKTkrq6IC7/bhnbYm0
c6wHCR2nv31mMRLYtQyNGgMU5A80GXXqAE7DKm5ZMxXVguTiUegzRyCI6fREaTm5
EN0SKaGSjqfpI0aOdhX6kClcqU0pU//72TnMtUItY/mnpjyFMYpo1xVx9D7vbJBO
HKC7TkJHxRnii/SqZErX1gtIFGjzi/9oqcmMnJ34n5qtJvQPVBihN22pBL7PgNID
bH/093nhJ1NnMV7mmAehVNG6QUsr0Ffe56nE7a9hpyVThSRecKYVRr7PDQtj6VXY
A+w5+0KWD4oEG/yvkl8qsuHXUJ3pATOIxXAencoLD+SVo1u97rT0y6WHMpTStmn0
s3fNtXwkaI0Gi9sRHNt84VD0uHOM/3K+Ezo4ESaEvS4RMMw+VGOZbzjUcIH22k8T
3XhrpbCRTchEfuM8yoZ/fyXmqpe0aqa924H5324iG9ievUp9CQnKAnMq+Rlvb+i3
vuK55PZrE/DNjlizC4Z/7DUIeZr9BiBYFlp9uWCg219SeFk4pAG/BP54r5N48xtL
cyC39OBPY/SkdZHhxrlhUL9SZ7nojE68zgIXEOUA++2q5pmUqOkMKyn1DG68Ht9U
k7G7rd4STYPPR67GZU/VRBd7/Mfpohae/cnzSK9STj0vH+sLtKbTC+UvCkeJVBlA
qqU+W/dU7cEJaqVYTkx6cgPGE5siRqnNb5aJryWCFjefD1636ea2NJf2rkKlpaZL
EG0AXZuVNBMeD35PVF2kpo0goQgBRhFLbJjzusM6looA9HT/ekYdrD/cPCsGplDW
h3IW4kdIIGNhpratw7LTxtMEQEIbmQ5muCHFQaiv9iSbjw44A1Wu9qH9/PNmRNlm
m2I6n5B/frmlZeGAEW86VcvLanuhPMtPe3NnpunS8X+UG4ma+EPT+M2q6M2EHncr
je9+dzjzCEFuN/ey7ygfSgMs2ttkMdZauSu2Y+2s/nbCq74mW2PGQRkY37B7GxgN
Wv5vGifw4lxXN3GIncK9HYHu0r8YFNtxv7Q4z0EA94lWE8HHsnB/D3swWyjt9Die
mAtfoETw/Jl3Eqi7MzTh2sxS5rCThzdl9iO+1UljetLYpDdPU1+sejbFWNzhT/LY
m3BwYhpIVKM2BHhWmK6CaWIwCcvQ1A1xw5DJsQgqYmfHZLPGGznh2O6dP/kUkJPv
FghmewkJokXc3fW+hS+uQBadjbo1dYCDz3zFTCXXXxfkz/fd579uXf9Zh2zLtAJh
k7HOwOek1chcZ2AoUVUa4fh5FhrxHzBtzuA+a7efASURKsgQBB8I1mry9Ta1wNE4
jVI6ItuZit7hcE74Yem/w2lX21Eixpx8LF3xxQDc0usT6aqu4g7rYmwCEy1imMdT
/F9BdNMMbSgutbxfpwWEvSojR9Ng6JJX4kX2kCsdNszFycBhqefMzYrUjS/cq8kQ
dRIOYZb96ksdsl5FALNP41eYIhQP6UtuAXXwiD0ITOsC1U6Ft0uY0iG97EcjBxDr
Vy3Pq3Goa7K+hPEkxJzoDCXNIs27R+IZACPM9Xor+xKPFk1eFa1ayVDiz2EWfx8K
jaZBj1x2UYN1WK3j1g35NyaCl8cMFVvHYSVLGqf0OZJ1qx5cKpkNLa7AjNZdkskL
jwq9TqcqBoYzAh6zmlE7P3fFDaJudQKTMtmCEWk8mugcVWed/eCNU5n5Kw8hyrhp
NN253L1j9I/s0hYNXI46nP7xuMzxK7/ULCfHGYDuFMqjzPfXvtBewgwW8lu9Fx5C
8Z6FVz78rO1HNcWNx7mQfkW5c6GzcsmH4cYFK9fLluG7DktEQ6a7qqisu+aJu7tC
yCT+BaDI3Nkz1PqbRFR0+Sv7jMn1261SAM/bP+99/BG+4WSLuAdvO2SzFD/SLHHR
3aRwQ7Cz0qbmViL7G/76m41xiNWF2SJ+MluFio4xxato2r3eFRJTix3Pf2yIj/QI
KgeUW1rUPZuoq5i3zjMP8OxfsM42BidFwSXQgWc5xjVYV5d/RWmJS8sOaZKJ85I5
7FRMgbRRHAd5ebG2dOhZZdWP91jj/DVOG33pe5TNvZxBhr/ESMuSjmCRqjj1JSx8
BlEUfVhmCYr1deAmrAPnG8bc4Y7Q45TaN0ve9jfn6xPn2lTCP62XsPJTRMNjdQDz
kDbMOonEHzRXrY6R/coeNx+Ar4dri16EHbrKDcXH9Pnh8nGRsXMAH9nnk1jUU/Dn
X9PSwnp9iTUOpg+wVrTgspnqwBPxDBh8pdS7MaOwLOW2uOg7nb3vWyHJM8pngfgd
GN3f9DHKsRMDNep95YqTd07DJcZpXr00ofIA0E/f5MTnyCe02ASsp4spPEunZB5N
ZsM89NUQmKrRvfuZ+nqaWMwJyV6sYEjAT3FvoZQ3SbLtZRTiTHoHqik7oKmKsjk7
9B47LdtuMjMuvAsp5le93e+pYpeO4i5MGi6ekRjPTSkTyJSvzR829Whd/lfg4pku
KQYB23GDYEgMSIvV170uGqktnImUPdt/ryqxgErZmfJRTFZAicV6S7C4Ujlfv5Kg
lOCOZjspEjSNidPMCS4buqNwC0lQMLXQKGWrMBaIPGio/FIrjpsfnXlk6bD0tjqg
2lLzd0nN6PFup0da6pZGBBYtzVUMEoB9VGhNVRDEZ3O3G3S9kBxH8/E/WUw+C15j
rYYqfKa39VddSrJtHHC2ehFXWD/QfwfjyXtbOqOw6pejX6GHjQ31oudmFDVC7BW4
sb6tMUtyNfItL4o92H2VlAf9g+xLPcjwTrbUzvElOsrEcUhsWcx7ABVdmybHvAeA
uRY2kvYNT+BRkrSIpE3n9PakgNW15Wk8XOjbyiMfkr88LdsY6R1NoAThRFNZeWKZ
g0lqIyRxXFbtp8E4OpKXX4KXdgid7d6qd+5IMd05eh74c2FpU3n8W7zKeyhLaQUl
qwuMnSzYon0SmFdJxE2r/342Q8FGotm2/H4fW8LexECgCtQSgqLl1inb9eYUtuuP
2TtTlFGlInD5HQls/A6TOgowia9t0yxlCmtrCTCi5QV+A/Ye2O4gqoEfujL+X8Nz
r+UpQVec5wZwy/QVk9je72lkUHfrLfM/jTTd1qZoKNO7lR5RCIWWQIBSt6cezhn3
ytp3bPfB82In83AQk4oFObrV2JQNepfQYfAElTVVlX1frL7pgFmBwFh7gpMyo/BD
qRj2I+UFDv+bPddWEU3J03xbH2KgB/tl3p5LfNyHUpqSUsJYnTWR0EhvcGhkQWDR
mqH/zRp5QXe8Oy9swNjNthHNacJwqvVVEo8hTMdsW+kPdL1V1A93b0qsOn+5aqKB
ArtGjXpmjLDxGk/oeT5Yx/EIjo58iAgS6xPaOAW8CNh+sIQTdPv2Ij3XZY3Y016C
eXtL34lLu6WjWG0awToW6N+WwUJeM83ToOzo0eUatM0ShFmM3ggtxEHlhd2ZA0E3
PstN4/44avuLluQVjhfuJOIc58NxYxS5ocqnJ1/qZdDAaU1dDPk8Zz98ayi1eq8i
M7nmdJ5bi7m8/FYDLSF3B5h5EP8zaI7nnLIiBVN7yqAmW5wCv5tBox8Dbv6ZWbmi
3nmznqByUn8Q9bIvvA2XJTEFzPFNO9GfzAqy657ZGYH1LHot/Eetlf14p5/3/2Xq
aeYofy/6sf5KnEMqmiKA4W5qlSn0wCG0YlB7Z6FzYeBw6s1bREUEH6uHGQ3fOr3d
AXns0UxcgKhppw12veOyOQWLWRTB5dT94hFJDYpJyyHw16mV5dWC4TZN7oXvh8cW
Nirv3yiQaSiss4+FXLtGkjdJns+D1Xbvv8jbN2PQ1NXRpZifBkT0Xcu03v9JiEHW
seWpM3arnWtl9lCUmahshgTzB7mndhogbAEGgev6kv5bCDzglQ9agxE+gnFIJGC5
YtQnYQe52dLnhoC42/rAqdRuu6enJVuyzsoZsi8K4kec5btvrad99gnxiq9GeQlT
sMC4XWXHwc1UWcqcBWjJ2/m6kZ4MHTkOEPUFvQeITrlAdgKVWhKm6cZgniDqzAGi
Fq/DSTneSR8fAJGvY4zHADDlK/Q2X7Crl6Y+aXQGmdFJqQlmWtBfN+XhXTuGR1ny
EyLCj3Eaz8yJ8WFdbBQuoGFSrUjZuJExQEmBrtOT0iTEtmVLGsAvnS0xpNV+FAsJ
MPuYHk16RUAlJrDhnGhi5qPwpUqCscBdNNIpsJIkk3fEGaiiPVI0x972vZG00q3o
6G9On3PWx09oW46K/+Fk+/UoCDaZ+yG88NfvQa4REHLT5AQlHMLKeAs9qG6y5Rby
kd4gt273nV4iz/8kWthJrSr/R02X4g+G1F5csD5eJjsg6Iqb3U3ZQ6rrClJyo2Xw
e9EWyIb6ovYzZg7CevXRMOVRpyY0Xm7PFw/bQwMtiz/MUfIGRHqSOOox3rwnxiqB
3wz5/DqgvBS365yU1VwFCeDRxN31i+Gg8pSoA6zZpTXjvD1U55aDzbdTLarjd1dL
yDdGUmfoxJZaL1SN0hQAQNigTGjfsS0N74r1Pus16Q3BfnrQf+4UIhaaTgX8SvKG
8zGz6MXYuMCj0xCQC3WTQNsErrJxZ8NdORUu8+S1LeQVgCf57G7YTWL6iS8uAHti
AUBqlSBfcCaGfUDBn5d4w4jhsyIaKPWlgEzQlmG6ighEpXwpbR1NCAoRjC4SllP6
oFttSP3Zpg0rqaEnI/3v+lS7ljMqmo61x8fSNRvekz9F9RCCvGeT++w07CeLFPcK
AZVXCY5dHpzBd83l2lPswpttUwTxByRoh/dXT+QY3QD9uyq2Smnj+Kk2Uts3w6vc
lGgd2KNhnkVisIaBTU9NlV0FCiJXN8Sd8sr90fkN2Vdh1bxo6mwz/GM9FOcRcvnX
c/kI4xCHofQwiX+myk7wr/zkjpdhb0LbCN9dDOuemTQZVuyLHZymbLKk9B52UaGy
iyBE3uPRqLDiHCBClGgub2OeH5mArbCXym/75ja5q9ZHFMR609Qv+ZobaAP7KjaW
KOCL9Tjc0DN9z6jfnQKl1I6yr+5nkfd/7O0ML3kOOxqHMyl32lVACd2XJJ/X6Jb+
w6kY8WNYyEtjfiWBIyOhmPiItVL1q7dDfJZyd5dEjYoHqpjmDvx22P+DC92n/Qkz
FVGbtFG0GopUh2JgLYSzV3tA8FXuGlbCjPDMgZ5jTZXxggL9/u35im6y1Rulb2tE
CGkhQaF/YhjvKhHH0HMrfj265EmSekjiFXRGiTW2fZQkws/3E8iTahLnvoaVYB1X
oYBdnuGnIgUnml9E7YflRf8kNtLtxapPL/t0VMsuwYk5+37pCewqUuTPHX68EuPj
/AFHbAnRfq6y+/on0/c0CSMnJSBvp2nylzDFtMnzSu69fGKMshtmnyi4L4auA7zG
gUKl2m9nJbEvrV8PsZ7hAtX6fHwnJ1fNPdcVLvhh/YxOeOKU0KeAsgUlJc7JD46w
uAKX3bbm6Jt8qdMlKeY5/mbNYl5UzvDy8am4CHUyvqWKbeHPQKe9nDa1qDf/XAfC
Rn56M4bv+2ODCZZJ6miOB7CRQwPd/yGTD9Yu1RjwbgdQd4ExFviHs2yaW3BT+vIB
XJj9sf9c2x0r6RINvO8lSrVFRf5iflvLRBe4WsUfRqcrr7sDr9mEv67OGNfJblT/
NlibBMbPYeHdBYrRCpUEqU/SmNCjcKDOD+G99A3YQH3x64WyOK8EZaRNt+2mHG2O
bRPoSvB5nBJ6CFIjj4VdQoFIii6j5IWzKHgOeU/Zkfp1oxeObZ5fsALh2IJRf0l3
A1yTYjdJoPTWPWv5U+I9r2VJz+l3NUT5bf7DivVU/o3mD5KyZxN7mzPwwTBiJt69
KqfulCUdQTO2EHi4dSVyOle1COgT9+hbfKY6lZQZXF5fPjqFOpwQg6DQI3UG/JmR
99Q93dYXwnDv5CS3NlLiCfI8QgEbTSDIH4E4S7vCQMb1LKaMSBYaTOtUwXLdZSn9
25VFZChayXMbn1ay1AJ8s03H5CHaN4Zzq2zojtsgOVPSYG6kq/nHsRpmlYz5mL5R
XRyfLtzXy6G4QTOQI2/J+OQhjnpppIiJyqWlq1KWzdiPsyHcgmrjPrefTvYurx/s
bhQPIYTPQ9Qk+T3bUwYG7a4aH3jCaV2/vhwLkfQprr4db2JpOoNarHsZB0ZBSpq1
cQmlXjm51fUEMZ9Yt3okr3g973TDF86gKpgevx5e8VbNpBZHjC8wAriyKTfdJ6K4
GAtul+qsYJUkCnQSJVUp/wfjhYUx0YbqMI9DRJS2XuesFEZdXpfCM3UtSS3MZS93
IDLuaXkX9ZhRue9j6EYzwSlF7MHVAwuaZmOnB6iJmPu69RBxWzqSsU0SrwrPPcZ+
4IoyP0W+J5lYHaGciNQOIMhcgHZctrFDS8cCtVschXjdg7cZBKnxr5z3B8TvU0mO
DrbJBBrZ6ISBZ0ugMOvgv1jcsghBjZLGIUWzR9DNpJUZF606I4c9Nbnu7cGWdY6U
VASeoC+tALVwgalNQXqusfL++zJGiEL3vhxlHwKWn8esP/C9rUg/d8T2Hxsr9StL
obGFo9h9ZGf/wsSJZTDvmq2GQCT/P9Yik7xmoMZQsmlVZ2ebk5X/LM5ytgYcjN5p
c97jsf8ftnI6tyHpAGWRGOREVOCnnu9H1hD3JxcVIunAtD8NLQX3mf6wgT7tlbZI
1WRc1vfFRx7xAmO44RH3ilt89OuNdRrDNjQIQSQCnkpniM8BwUy61TJg6YCj3rY4
cyA1k0q0W5Ygksj14v1rdl2jRs1GeGH6S3PtuH181mUIalYPmWtE6nMGr5bbwl0A
e3bXRYcvYAXxA1DzwhyXUCLA2NXLPpQT5nFSVB4H9oYSF/xPQzC6vpsQb7UyvHvL
gtW3d57Hd8hlY82GJpSx7n5e8FwdVp4rNpKOjzKtAXxVFywe8S6HKn4OXAGAcM9q
aJihCpU1zPqWXP/40Fm9IRk7xqZQcWKRGihl2xvoQ0N8MAaKUy7KphyToFt+PzZC
UD+7CdBziSVqmx0iAr/cjHrlwNWGP1sCtS35PIiEwrn5nEcv3zlDEp9pa+MoRSXK
XAL97VQrVNmawDMur/25CxY3da+lz/aWu/X3UHc4BIMiLprt04b74HYMTK03b16h
q1B5/JRDrychusNDBlVF+HAlHJ75dyWbGldJHe0m/WiF1RWcflyY5A/TPFjTOAfo
MObwf/9mPjAXcy8O6qOobhHesYoKmL56nXw1yi8n0Xh4qDTh9xQrBE0dL0PFgT3v
UDjTw+Lpo9+SRa3KdKTLsbkyD/T5DHso96inuJqvVrixm1srC8WD6DajYESqqCSq
QfLGTKd+2Jt8X5052YaMx3NcC4u/kOJlPuMFh9FTZ+whUClsxkgZ/4c7+REbxiXj
/FWDDnqSaOCaDg6YSl6KUfY8SeoMMbDwv6d7u3c0h0qBIsSIPV/Iy0ei43kkx0sz
8JOJBk1NGJqokAGrqMX/W4XDdh4ujmk1MzJdvroDVnGb12sEY43wfKgb5qY5EWQd
JpbKl2wrg6soOjLHH/y/sDofGnSDSyI+V6hzznL8ZYmRSmoL02HJAqPAA7ZWK0Sf
JCJuVP37Kkw02QCqNORFQypoNXkzWoeSS6jex7S9nLPY2nGn1DFHqRJ3+nvjumai
p4Zdj85ZZwcC8mLIQK6mvBtdZ5uzxukfVsZemrd+Zy8J+1VbUvECO7VU9xcRGc+n
AKi0Ro+US7rfQi1VIsonwXGGV1ls0eTbxJoh9LOunCo/zlifNKQca54TyuQSoCwH
GaXA/qtGz9rO3lcmUqCoxW5sAWQfhrga04/z8iMQHihJnRif3hBGzPq6/ntBz9pF
HbzutbiB4FEu74GX5hbAqd606PV6nE2o69CnHOu9ss6J9SC4phBNqvhzMHXfjsqG
4uH5pWZNLoR6D0hPkAKSOOrmPij+cOcu9NX1CMmu2IsRkR/vab5J/TUaEDDPy0UJ
TH1MRa3/WCcM8Th1JXHN8cEDtQnxU3OQNwySLqZlOtHOC4zpTfGk0oKA9z0Hthpf
Y4c6z11zQYGM2X4AfeT4gFjXuzG0k0emiks1fXHOvDn0WUBpvLGqg7lRPh5C8N5K
xtRMfvv1788F/lGu54Nd5/2MV8PpPSxapk4omyR4/FQe0avAveGcSpRmcuiJjRZz
PpUwwlQ3yrRNYOWoSSgvowErpxglHh8db6Bs7dOQSMehPPok0naXAspeG/gRs426
M9GRZPsoZ4F1Jv5IanU2QHLMyUhskkRqzcPFw71JCjlvaJiJVnFP7GcF49KaTUbr
96+zLdRNssRGGVkiBwsV5OGmMyOTcxcUX1C9nBcMkmiO0zIln6lkCABBIfah5Tyy
X1TFjWASIGggetTSmqmXtsXokFFgR7SF8bOeCTE9I7NDS2n9+2hcFzsJViivVbcj
BRxeIoOftM4iAi/A7H2gY37g89rbmrmkAAPGie2nuF/Rv/eLPSCYzZGp3h2gwRxo
Iys9TY7jlyUMM10exwxqz9gQmVCmIx1febq7PoGOJvkqTu5GFLJ3x9OiEonQSbBU
ot3Sotuc442ixwnZssYRvTL3LKB/8s0O3/5VsbCwvSdh2bmLR9oKuNjumdjtO8lw
1L6l2Hyq7QeOerJa8uLp7SkXwrj6nt8XyJwl8SX/yhLI3wDIRCa0vET+zB4rTeet
k+GDIrO1QO9ig57TgmhgzXqVPj/TjQq7F2Ta4w8d2KE9MaHpVv70DPlPuPQODRV4
XocvL3u6gXtq+Yf2Iynljsg/Vd/BvblR9w8mwrnNlqtQn2YSBVuJWalD8ldpyxsP
anhx1rkOENFPzE4muOjdiLiLYrPj3S1lhXqyLesXk7eYLNV0laHGqbumebqROPGl
xzvPg5omVEC3X/dAJj3PENQjuWmc/NJpOwzRN4LD+5rY8GfcWv37gV0sVJkT3jnq
HOy1RwVyttqbxn/CvjUXrMAxNoXs24c/h+ncsPnjhgExtU+TLcwUJmV561dbckLP
VdvTzHUNCPSGbTsc7347weHGzY+0KJcz5cVdq9wexz4SQT7sHEAu/D/eXaG4fS88
J+84caBXNUQC2Kt5WJgD/V/435lbXK52Xh9liIY5CuNu5NCQ6yWkTT+ZmmmyIyvk
cOC5lftnBK/boBmVM4KJf16FPVToSd2G1erbWmausmg4NkN50Idw6/9FudRvnV1K
2fmJ6HIooxOtyY/wMvwjGFIL4IwYyGb3Ao/RR9lmA5ZSkJhJA1mx3PFJjq4lLP+u
K2yrMjvajuR5rdUFuYClHhqeW1MJluhhmMuWpaRsRkLHw4FoFpCu8EWFQ7i1WG+v
mcxZgiQFjmda9iCJy4NYy5QvxYb+R50a/yNRZ3XBhCcC6qOWqYTqB+DApbuW/mVh
msjnubwc3hO5nUok3S8gGLLmNFBQJxLX2YCb5M8Fyymb72XFwN3REUcCw09H8wGy
lAQ6jHVasyZmuF47AURlWrke4OHC5/RCv24Rw3+nwh3FnEmkSdri6jkidnWSqxxz
alTSe/9vdcNYMA4sbEv6VbWGJ4WOKfLvYIoEugNYUpoaU3GCxo6mAEaris4oVjHy
WQq86161XuaflJmwErBpj6YAtPhXkLZxtVvAermqmbNiAnCv2IGoHlBnvOCtDxEu
041jIDaMbbnypR7mVzk7CDU8nTaM3cPsfjg0N0naQdoD2BOdDY3EZpQPT9FeEiPW
H+16gmnN/DgYp7K6cipj0lZwBj3HlyxYoqz4mYu4zjIibrLbILpRBgcJ9Lh7zmiB
rL3bb12vASDY9OItUhfyzJxFq0BnDDGQ8RbgBRmVu0RV3PeKZ2tjp8XYB6eXL2sX
Ka6e4CYSzVPwjRBgyvJNrGu/WEUmpMoeZtWD4hMBSG7NM3HuNNuVDklVtDkMatSu
iJkmBkK4sP7yLIelBCQchnnh/z+ZnpitOhq4kvD0vWsPEKspUCrJAZ9D23DzVzfV
RFg4JNMGme0lme7c/u981ZsEERJ8EYtOHZ78Vk8a5Ez31OGx7pO0Jbwb/w/IBxOm
raLNR+XzKRnWkuGNerYZb6gC8LC1PotQcDhxzJijlNx9xtbl4I7/RqoQZBzGxWQQ
Y6mOUGjL7CUfbra8tdhmeZgffIzzJB2OVPl2ZFN1FIFAkG5vCFIJOy0A4G6+6DIo
q2EN9Jw3Dj3ZyVCsnv+RWpFozaT0P/zfJKWpt3puvDwGgQRXCy94DxsyDF2bLxRh
bI2dKka12q1RhCogikpOGzwNtWvzyUI8w2NcxG/BLw8waLXccVgNq4f/PQqawN6+
Zeca1KLrqdSN2nAH+AWHEfkKR8SBTVaeitX28U4EIFOrqCGc2gfEpfLul/L1Iycd
FpbchzfiOTYumKhQyNcHY+AVnEWlMaONpCQZl9PUoUZHrufmkaeP2Zdv0uGnjCZG
8tH3DPsZQo5bk/T3rnzlo5GuQFNj7PZE3jBCPW4WmCeiBVM9vxjqbXeyP7Gq/MM/
rB1/RbCEymVtrkfm7B7BoMYgZTipDo2RMyFLChm/RsJCWnTg+Eb6f+dL0gmrR3+i
r5aq8uEoCyY7lwSAd6qnWZGhLG/XcD8GS4J655oZfj/Yf2IBFWmqx7+64BNWqPi5
z7u5P/v8d0bC0nKVrz2lM/bhdyz6CKhinx+Qaf/c8AtC0PGaXaK1y1Gf0bHtiUSC
OWczDBhdD7Z5k0Dyg8jwEfPYKzDQM7e/j4eu2zCWrJV+h0asyzQb3gNHWnywnibw
rF08TJV6C0YP6UE7kQEkkV3un55ViW+tVo5m9uMAs53dSHvlBMee5jESYJ7sZ4Zp
PlUHcyFaUeq/u4tOW13mfdaRewKrjR4npMa25a8tTKlGm7ekYyzPb4sXEKbL6l/m
3tf0GEYSoPr4FF9Fq6ZbUgrNV1d344T4cAPW2ZmBV5JmBxa9AH8FSErXhUB5DdzA
bCRiIqY5KNjGExE2rXN4O7VYoCNaJ5QUjBJJDwRhYTuPh/omn1BpxMzUVg+BgkZj
vly01cvqoggrHdLOqmU/sUGNvIF1GDjFvTyjfLvcrpaM3rDylXdOwt2RRf4GPBII
RZortmS8d0vJ+j2dfQVj4K3hIsDu80ZdnmXKUfjpwIKYJzQXgPFxdgVdFvrbk6bh
95xqX5WwX2YvLn6bTSHve92dJyRirimpDylaZrEjBq3TCUc/lbpZIi1+mo2vc7QM
auKXhIzkb8kaVKRWA64mTigc2JJtP3Ij3PVHzkwFhfNKUOsGpdAvpEEb9Xj1u25Z
zjCL7HpzGO4MoIF7Av8Z3/o9xch9t5v+wBtUeAC6bXKbXxX2zQ3ezPmhh5aAFD9S
5q6xBjYm948f2Ffz7siRPW4jbFWq+w/8bNsvoxQ05nFCX82+1uxNEQzHaWEOLTmz
`protect END_PROTECTED
