`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z0JPm3yO3vc410aCps0ruyUoMf9QuEutElVmej3fw8EBi1IyXGd9+RNCIJ4fbHbo
JkF1jFkpmlR0dYrhUM55AAuG7/vEVEotlI1IAMG/XvQ5nIefBn8z1v7izZc8vqdN
Pr950NQGpPRxU0yCf8mfcGnChwMC/tTuBSNQ3Z0YM+nMCGb9SYAiP7wDDeIG6ZEC
zP4Y3s8o63+ZIx8+ohRdeR50BFOPp5Fd+vRm/yMGP2FA1LtI0cMg9uPpnJQNdEiT
/X24AARayz/nFP6s3a2MAQ==
`protect END_PROTECTED
