`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mMJOKmW8i8nrkz6oQSMlDR+yO1xfSCg0gW5+bYLl5aRe75lZ88jTgdMwwD9fSQN+
CGd5eWK+jumq1huVKoBxvEDjuQQoaoeUUoYZxrk6xuU8B4ySM3xCEi2PMqJEB5uz
ZmIrhbt1boLE5wWG1xhnkAoIN8IrZnO06ewRcidawyBIah6WSKp9MhYN3SoFeX9U
8tbu24LPpgZn5JPRexMRJrPwqcUf+ob7Ji3QyBCIhJHKomrTH2ydl172T9/NijIV
bROQCFrGEt0wnzNyyvnsINu570ErsYe0tERUmUlXaolf4QZUaKoEWPt+dGippRpD
mZn2GLUbUMw1wsy5q5ryFl9UclJUvMPkzx/vJL78Xyb77i2G2+bg4LpwBJLRCyIU
hplVQxgTYksoa2hplMX1NjZogQGRrx46CTsPa49Jl3AfMxdLVCsoQfWI/f2+WM7N
PvNUBMpQv//8JBtIWa/xzfFRgwjAqoMvMxovyFYeHCsOVzBb4TmST5gF/7UU31/d
z1KBXVlKAHTmMWSGJVWGyg==
`protect END_PROTECTED
