`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bLZGEdwv/xvreYYgRfiH4NFLJs81MwJg70S/w7xkOAe1vh6GdPxBMwMJgXwZWY3X
A8EGuqezRtJF7Vcie9xLXjq2mvD/Ut11wEL/LAwiKE9ecO76Nsu2WKvEz9lrvR6y
6TXYv8qZdEs7PZRlhK/PA68OgPqHsQoneKOxfOz9Smfu0IjuQTZel4NHne5rgM0A
X/IvVx97T4jTRB76Fe6JojTRPsC3DjsY7l+9SHz6VRJIKf9hIkFkxOl5gD+BxxU+
BKhec2ppXELQ9FuPj7KVUhfJ3xb4OrlTYJHmnR/Tm4EzdTWTqBgMG2K1M99CjMSU
VFLCpI9DtMDK4Yy10dbJU9/ZBk2irYZbfcg6kfMRPgQ4PmJ8LUJpBwxfmJXfqXVM
NHpCkOPwnUFHKdD37FgMDA==
`protect END_PROTECTED
