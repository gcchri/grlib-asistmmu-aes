`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ak5m9qSnApyASchpzLRYMuIxdTmdTj2JhodwTmO8w95PLQsqwfgxEfPFUxLxOH/g
/i2Is2sjuAgvCJPE6FVNQK169fBc180tCEeIrvnHr+VHWl0noU7C8dddYfKUJJ4F
bZEDiZlbn1Idw/lyzfZaKJ7hTQX687/WiCSDISFCPkL+lxxg3TEzWL5sJ2rcu2br
8RTa8Xdc9WlANvvYgPgK3u8Rwuu3j1KnU+0cX6Qqi+ij5A6CLyX+0u/mb7DWwSdn
djiIB29kqOLMkUt81kejXiYwKzoMBjsHcWLqscBaml5S6y2QfPLrlR0sYNrJUkJN
`protect END_PROTECTED
