`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NsVxlnLOafiQfGM5ZLjCswFXeD8OMwqxRfvVUd17ENZFNg0+zF08LFTObQSAM/sZ
Je1AIsNR2qjMp04i86PM7WX4XP/L334GbOX0EaaWOiVqzbPeyqVxKyOpkMmC6YE5
3UEApZlbJTF9npOyEOPMOca4/VQqEiKqN7+R0KYUj6JarY+SwCptbdlWfP1rBQMd
HItQmZKNqm1VDZTUxunkP+H1oPs/1ndfw76Hfc+YUXNl9XIlBSIn/VSLfeSwzD9D
TQ14bMLWHoF8pprwIDDI31MIir3cMQPSF744Qqy6TMkF2cX4TwwW350TLm1txe/p
uPAGGiuON60xye15qC8fGju6LmbwO2U+9ZRV8NX7wA5aIWd6NiGbty6VLcC78U6N
R9nZgImIN6k3hKCw1SxWM3Yk8HcjNj/tHzw7+iGtlv3dWPNh+rDMsQC/WlaL54rf
`protect END_PROTECTED
