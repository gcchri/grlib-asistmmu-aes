`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vzGXO/TseF0vnk+b/ZbjIvNZa4ng9S1D8Eufdw8DQnMO4zWkjY/k4418n8D2Fg9Y
QGyElhNEc+VQiuhImW9gLyLp8BwJzCJFP7A3dqYpDZvWki9v2+uP3W1/dEi55Pp7
feJzJiS0EpXCS3H4Iv72uN9AUkKJy+AnFDEwSVJleHRTZNmX32iUJX2IoMvBqHBq
jEhc+Tsm3VrZMCWn8LIgJwtNcnD0HxYBxygxTqEFfBPoP1CKTT2EP79P0eWv3T20
CXqmzmlQ3LQNgXZ7BMtk+fBqsd8GE1K3rjyeKMJuLH3B8nTzACtel7akF18x2p2L
m2oI/o1JeYIBbB9362xSl3kuGoU1WUYWrRGacgfhYFsaA1ds3EB2Am9jKIOkETXz
tB3wzJ5xttA9kCHYN/ntptj1jI4XdnAolz1OokEr3AxHVJTjO7lxkWmM0YTZwP1K
rqkz4axxovsIYtrvy7NY9w==
`protect END_PROTECTED
