`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZdEwi7anjBYDTnDSNk7oLDYTC3Q58CNB6u4TDa/lH4gsSjg8/NazaGCddMSmy4bE
E+vjAgXgq0awaTXgcJ42XjUqafPoTJOqM+Y1XW5h6sSPfm0j2rx+yiwQJIsL59c1
OdldH06FxAE4j2c7SA73m4sgI50N4G4FhApa+V6Im5dmISby0XOnlCZY8S6kFH/1
MFGNakTt7yHYEd5Lta4LfiqAWegqXY0cLVMMNTv/2CHTRQC5SqrrYtJPtYbWTmFn
4rDufe0OwrhvVc/mNYpg1UUH/jkgFmP2nBpEargCVSBqKqviVYEk1ZfEaPc5j1s4
vO3qY4S7hcahorVfnxVql6N/ArYSMhG2rpnvwaEeijCkJmBJcDoBWiQlQKKxL9Li
hyaIWJLi1NGhGj41UB5MbJsiu+osCpHqjAqbZCIrwKyWYT5wR39wrR5bO4kapM7Y
PxpD3e+u+p1VoTBrQ0/1Pf8MV67JcTKtM6Zu1N74MdMOsAKUbL2N7IEiaVO/Z78k
1g+ZWqNpbJZC868LrJyUxrujTYxgZdzIpylerp702mft9vXKw4UxeP+LxTGvPYkT
mig/Gjckz1Wi87FWFQ4PIVgbMIM7O6Rj7k/amDLXFtb3fKbZGNGhEaO58Ciw2MGo
sg1cBALyeqPWCa0Iyj8XzeckZ8laBHi0hNVTjxB7ZEwpW7znuEwb/77MeLZ5Joy1
v/2r1+58ZoNTVrZYxZY63fpxYl7m40fjvGb53wGVg0f2svt047usQwFdPTE7ZGu9
snrbU2EvIWmuhRrj51/7A6Te8lCDiQrWuD9pLRWjIGA53j6uu9OFe3+HN6EHBB4s
s2b63UO79MH60isa+FRAvvrJjXKLXseOOZpIT0NB4MNvtG/y/t6cN5YuXh59W4zJ
Gvx791AoeL4/arOq3edp1zb1SS8LiDtfH5ZBEbeOTnK/kiOEjo49MKMDlwzjc7rO
b4EwAk8zzXgNOopsf+8ttrOSPDK1buIkxV5kzuvv7xayR8sVpZ1yFaKgfdJbgXj7
HLkGFpsb9Qy0P5ie0v9qUJMRro/so8r2DvpNSgDNLyZI/q2Wyjub64upHCjACZlm
qeZsCAMUi8vzkS3624YVrG7Ds5Ms9TFpcoBEy+ZcTDkw7XVFV3azVF9JYrrV7qdt
eKBpY5W9bnDj0yHgy0FwacZDBZsbtu45oB5f6Ua0VoLwupIwU6qVKbsueB1avGa+
JRx46tHyNNZJndXGG/yy2bz6KG2H5Wodvi6sWDrSYlZYOvQA4NbJcPHwiuDRumYg
TwA6ijL8VbnnK2ZCYl8vPnsEmvEGs0gf2WfZFfvHRwQ4pWN6uIAjFnyqfsaWGYFL
f0auX/331R9si7YBKhQQ3RjpK6O6sHYDeIBBiSCJnKGRLFQBsFigryv5ueGpbBnn
bcnaf9yroR7ag73o4c8FT9ZuvHgWaMhVOQEh5Bdd3wuQZWrvg8PHyFkZ2BEDorfE
4RI7a/ocyMmR2/POrzXX8RwZd/f6oJXz5xs4c4gXRpRkDXsCm+jGe71F4KZFfiiU
NaGviCTon2MfUYs3R+UIDzh9g1zxt7ySvkhDEud3OAV1vTzfcHhrDKm2DkJwG/qn
MqT0G1G8F1kED+v3P6pw9ayM4Y/eCQ/r9ty388W7Oiy6o1T+s82RhPOccIMExmr0
+uJ1yEspVKiVMezHD/aRBIXLoqNISsd6fnFgi6Eda8EHnvOxWbuLQ3kxz3iqD/qA
39gzklLeHtQmUxclDsH95FEpFVngxc6hs1R0RWPnRR+lerWl+q+yg6MLKPVjNTXb
BeNYU5odY8Lpk1oMHYzpIzfY6FvQoEGlmXyTmIgmjnIQ6zuDIgY8AYshXX4V3Bz/
zhUg+SDjPXM/mx1SDEdy2jlUjIRSiFxnXMLLe17hjHNtYBC1FwRx7ISWuHgXvqLc
o6aHlvkyy3IAhh/fuIkNX9VtERmlyaf5UPedJLOWyDkLW/Y4YGChE0N7avS/kMQH
GdrPQm73xEM2TkkOqsvpt5hDTEQXErJB7K9WNYvLkYoIeBt/Re27pXYmP4KSeRGL
r5oi3Kn2Wbog7mLsUjLF6MiBx+4WzII7L+t7K2Fp85c=
`protect END_PROTECTED
