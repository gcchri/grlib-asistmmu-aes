`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0dfgor1BDO9UQ4UdGsbXfZ8ncJbDSt/c+XaSQmYfLhYW/BM1eJSs73BD8mmeEk70
AQiwCgJHXdB5IlKmWXBJKi1gLxBcp4qG6U70eUNIvkObI4qbtpXT+Ya8SghopIPT
hN7HtwWR/ZTZgiMMQQ7yl7Cis8IKGbndHpLBHBEjacxCumk3LlB/ShH+8vLvV/tE
OWyUC9pLmM649NzVtC/TjYUvYwGcEkwAkM7nhBqVocoZ/UbnXDuMkvAtG5wqeiHs
S66GlkTpGzOqgiFTOZiAXwk/itGG49mcbMSaWEUMBBOzL748ha6BXDRD1qBfCRSx
C/CvPV+ZL+qFjczzbTHCIheYfRmwc1W+7mEtlEI3Jx25MMMVUBt8UBgIcVVQswDP
x5JHyNbXIUX3YgUYL+p9FWgEJCBlCs8aE0Y5GJ5ihcT2H1dINEVPk4bCIyM7uu8J
sos9rz/GAmTZ0gEFL95RMU8OLCk1mvzbbVJPkCq5OIbVoyODjgQ7PjoVE3JD9NbJ
x6pVqP/Ew9axDnl1mK48WqZIBARLH/A+WLJBQq/1uueDYh0iGrXv8+2slb2znqkq
aVC1m9P0mCvTtdwwzia0KCnz5anZ8lcXS5ycaSaY0vN/pSlIhLB909moQw4fNRY0
m/ouYmlk1wrWXreBb5qUU6gIGtQhubPI3M7ZRo98exgLClLje8OHDLEBEbRXdwNI
IHyYjzjXuXT/+bguuGjjc7FP6RZ8wn+TMkbyUkRWwsDDDaU4Xds2AXxCE7WEDUj2
3TbCc1V2a1TyzJYqPboQJJfvjdfCgGG/3Jc7VCVkz00Tca9jPsI9JfxlEdX54afS
hRR4EqtgoOAMi7a48/c2rYagSuPuJrjYu7KZlkQfuALIsrWAoNeW3jmbJfI4NqnQ
lazz3k3erQdqeN4JS7utcCmK4vBtr2xHowC0Yl4nd6T13RTqOBlp28kSYfoLm0XP
HaRo85UQkkxib+dwqyDsPvkuIH8m7vK4q0xitWeDmFqdgkKmogKvZRCdN2zbnBCs
Jbic/iONK2fJHuR2Dub8rYQRAUQFWNUgcW/46078jKFmMP9Ik/7n6VZS/W7p61sJ
QobqObO7ND6qIrjyoO4hfG7qItnL5Jl3w6pJCZu3e/PzQG7TZKSckVcd5Yhn4lzT
TCA0b1DA/TkCDfR2NJWZTk6HfAwfvCkPAg5RO6Sy0yjLh9bGK+vSyJxrxT+owEGr
3RwnwyCKAV/wnIqsHklqHgd28yoN/wm2zeaB6prsgG4TcIuC1vdaggJHb/y+OTkQ
K2wro6eYxJMKF3VQFXyGkIPriaoyhiwP72Cwv6yM5fiv8Sn3uUn2IogWBrnEBPfz
vvzOw4KB4cK02cppgT8WIJ66Qp+EK9sYYbsDBwwGD1diHN7FDawdEWL5bQGjl43Z
H+mdtGDKazIowZhJN8rhZNgRBJzFp2nEaN8DqeG7Licv/Y3IT6RiZC4LKfGQIrbt
zmhDUCU09DHSl2VNs/XzuWQa36omrxqBDABH+2bYEyYmU/mXFlSPKauf2XAv9TuA
KilLLt270fjBTJme8TU7eY5Q3aPQMndZ6JS1Xjkt8Clj/pBnIwCXmCaSeU8FT6Mr
qkLt2i2Uso7GALpC0ynqUWCzMeQVLPcCOgHlROHlmVEJJxz2Sp/OheDE1rVatQ26
2i/7W9NU8kVvjMJ9tNZ6FtbXBIfL9toQL46e7E+5DNtj+1+EUdXOxrX4vgSaIIJZ
UdRdMhTS29LKo30bmSWE5nG9TBzyQbC3UVh6zOsuUa3eqcIZMr8wIMc7N0I3E0an
VMzMBtvFp6W5Xa2o3Oj9e0AFas9FIlcRUfeWCtiFX3AByrD12PwF0MxNnBrxXyby
as2wIsvBCUa3D4Epsg6C0ujR3nIC9HEiK+Bc14PQEbn1msLQRfRrhr3qAT8V2gCu
CRgMcxKKgz/vZQVqTpmpRpXzQNvbHPOZk7WsrBdtIWsYdngCxd+MYDt/I/PdR9Kb
MKPIjQNWrcSACpH1fg5ZJGLgXK/aSL7X7Uh5z7q3TzKuxsRDO2IET1Y/DA8Y/N+b
esmNQfnzQMcCWei2AMHo53Om2nqlc7MA3Lgb0KpTEbPUBkSCanqkbEjOe9sA8HwB
PvR7Ng5nPnh9vPRMT3YvxWE46Cje0G9SBxPOPSETaWCtytmrvUSFSzkMYut9590N
8Qr3zTlwPy4MECxEMtFuhfUA8EIjwIDV4sFxrFHEglePDA3vH0lWdKEZWRmibBLl
yjOzQHPc+rhAwhvv1UzuCJ5W8LJ2ie7zFTKzHjlduIPIYtU5JisVzkzsvhS9959j
MhFyo2zcqlvTCO0BxqbX81vUzEbJG3FvY+FKTX5YyE3tulwFCa6gVdq9mWK3a+e3
MQzjoUDL6kk22PCE7tlqPWcFwWKCJ27koX7n4T36FcVQS+Ezo1JAoyA0sZ0vMC6p
xXSATMAuiUL5TiC4PhFvWZOrHsyOr1Ih8WxHeyewm4BrMi5pBWYS/BBA2FVR8rq/
uFBsuLMfNA1HxnXVwwcngxR0ZoLUzXJ4GavemFTpEmKbmoLbSC5vvNKZvn+c8z8t
AsQxI9Km0KSfkJXrhWxRPe4v+DU7VVIlOQT2twG5yKmP/y84lqD+JyDf+Wh8msFa
qhb2LmqCFftxmXURV4trDyJCcvfDnIruVyZBB8k+NOhpsXRGFqxCNG9+E8JTFyTy
5Vv02Yxz+inCdrmlXbhoALpdjLxPA35EE8Nj+miEG4pEACEClnKJxKb+Ozxkvp5Z
voD0dw2/D8iwSmCkVFvdNUgRE2tCjHeShUImNJRMAk8cvro0l5ZXViZruMWhGTuz
iQVEyyiJ88yaE10ucSYIkap3FE9YL4qgnpz9JfMViJWKSv+v5MjUEq6X6I2qQZPI
+J49MW2LSzoLtFBqU1vKPQ1hOgtj7KOUFtXDEOGCqE/S9VrsLsBsQ+JW76o46oCG
CsycGsik1JynaNAtVPiplR3LE94F06xCAkMGpdy/hsC+gXnADYH6rc1fF5Tv1nA7
mU1Es6/4fZ7raLZN2/ixlDHgFmNp2mKNPIxzCcHRsDjOFEyOmH0Q/sMc+96CxI6i
Ooae1ykqwWhDg2aNIp9Puz+z02Y8VFUeCSsFFyjs3Z9CYLPwAf+PlpokD7pRNuuP
N/ImI2far/DsFPaJAHqiJe470H3RgFKJnQeUsKzBEulrP2NSe/C5NLyPCXl8OpTY
aRkPaVhBqH33PbtUgUVkcylrZTawvixdfxEHqKdLerRSiMxI1evgc1Fr9faN6D+o
1ezMCseYpV3ECNDIEGFtEjbjwt8T/BCAn4UpyERo4Z4Czth8v8EV3qy3oIn1HHDh
WkenslqkpEH13KC7ZGVbLMdQrzWVWGkMBjPdkwRz4n21098So4ukWoiyzX9EP3SN
IQEd/Ns854o3vmIxGAPrI0yB5Do6E/Mz72+iN2J6TOClH9IRxd4e0uEq43SiCalu
vzXBuRPnPmbcweWbxvYs+qbC+1ch0WLKd+r0tW/Q73woig34fkrm2jyLjurxaEtF
P1CEAgHNzShbYdhzAraaw2FXv1WPqUWqFjJVAK9NZcMP9ffJA21DMVYENjwVXzV/
hupHnjxdRLU/ebmA9rcD8FAMMZzNHXh0U6A61fHLsSPawIepAZzoyPQV8kwBBIDf
OO1jgJpzCJSqdhPRZgBcKPDM6XEuf3gMnXsTE/N7XzG7hi8s3nHcHEK57V1GfM+s
/8ujXXVDTlK0Qlg6s1p8NLdaLy+oImY3R4cP6f5ijwCo6GbzjPAd4hH/HaS5wrDQ
VkynGtCjehYW+hJ7FAoSEPN4MMAEga9gROSL2cVpKxeMKDdqrDcXr8987G9rN50x
DO3P/fLlhH695m8XOpabnAsXWX6bok9pFCKkyEI+TtkXmGZYIEDEgEpAw2D/agNf
V9hXfXdwVYb4SpNIMWhxVrSHgB8aazF1MdlGfkH4UTAg1xhS/KQT30c0vii51sTv
oMen11Ko6+uspUMY76fkFGXh0ToG0ndxU4v0n/BtMFkt+kHlhVwaUbOfHXLyRM1n
BMOxfMf3LWIhv1xQcWqrsS/Q0QsDLQPHaOyfWo1VygPHOrLESy5JqtyzRnipLvY0
Q66Ak4tkxe1lYfCyzidrgr9p0yZfhZkHXHvbrW/z8EgNAtzb1Q3Fe1F0nzfWomeB
E5a6sytCTD1h9E0C8WUVTqNlfoYAZdqL8zF+mteowfXOm/bLbJnSV/bFnpau77Cc
hUVk6eGFD5Yn9q/ABFdBQj3yoZMkdJ4lCavpDhU1b+tnotbuq2LfsGjHhFYv7wqn
dZy335HdkenHN3qIhFyODLumsS0m23/e5qC9xHjRFjROV0mRpVyR3gNF6LMx2qyG
czaFt9bFL51tDoTj/QHK3xBkG6KjAiihSD1johnQLpxzwbMT1wfoVV1gXVfMkhM/
X3H68pEFHMu34rtdMfLvbe7Bd0EIeo/v3r9x9+3JwCJuS6iO88lN5Kc9/xekF8CW
QL5Ye3foAUX1zXqRoDNJlDuReQIlP8kYrqimbgLM7bqMeUPVEU5TYS4rFzMBsSs2
FlcYSIeEulGjGzbBXjZtngO2XL/xEOZneQhUjSYMYWolB24e19OgAHqqZv1wBOTv
TheHJ+mh0tVMWtqBLGRfq6sWWVgufberjMvzdejGpj7FBoCYZz4a8f1OaeGPei9K
dGTNnx0HYlayRGdmMEf8BWVhDr2WVfySV40Nu77J3WNZzlVnpf05U/Dbxy8zQlpY
rP0ylz78wpWkWSjkAY2vn+jXzUvjC48o3vDCLgPlF8r6WMbyJshKAWfrGccIoRfp
woEAxQmcjsH/mMOB4LzddS+avy7B/N7i72XnQyWYYHYUM9FFY9WvFKv+sLoToqPm
ZyqV0KWKF9L9Wjll4LH0E4SWM1uHnJeR1l8OsPVhTuPyHzd/e0PqNc48aBbCldrY
2ma/I1/fXT+PUEkheGi2rPV27MCo074zq15nazMFGAkv6eRCfyhDb0/4NX5uZlqW
oXJXDi6r0rbo0YBy8AdMEgpsSS1mC2twTu3735aesTadf7gNnXhweiN+E/T/LIo4
J5EZesMrZq0HfD6WTloOjtBoZ47KYGmI3Ul7T4xxsfigRCNnpvxSbGh/z+JObnrR
LtnS8Ofq+psg+id9JiISBMfnoYOQWKrB8fGp1Mb3YFcIUpRZBQhVgsZ1Zcq/T5wU
pWutrj2hF5QrwjYcH+jspGLCNO23AL8tbvRaM6LsNnSJ6Km7WTV1gKUD/ADU1BcU
Vd1f75ezelFu6QJIsHwqKImBVA4JUHy1aEdwlbwGzdjQolOEMNSaiFS+I8PC+V46
tj6j3+vqKpaCMssc1X7qaJ7NrejH6itIUhcN0zwSjI4K9wv/YAAjw2Wbncim1JYf
i7BRrEY4/kdA5IqbQU5/0ikYMsZ6iVlQ3EIHQ7rzeD3IGjRaSlDHsG1JkCREeKUw
gUK/n6l4zQS8TPhlo16jMpG7shbQpWRaks22h+wZNhicsAX8n7R+OS/Dg+JoCNE1
JF90LbAPJ3bZNqamyknwfUYFUSc35pRr/aCivLIr/3VCTzC7N08yVLv5zE8H6CC1
Ytgw4vKnD8MByYOn/XBPjFfOyDagOMzyF2cJuZMCJ8KvjaT0rZ6vhgxE3M3lFW6e
zcefezNDaCdA95U0M2nyYB+C7cfzQEh6LyzWFHIPbSAHwF4SDjCZOaH4CK3EQ2xu
j5khqFG9duGSK45ogr3jCq6TFRJrxXQlrkriE/jgL/cWebq8xR9u0qvesNZTMT9o
EaNKv0MqMzkSuip1Ux6JO51fjY6VyPOjLsNdNAGGMB6mROMLgwanIHGXkHsAAQsz
8ZOEbyZSS/hVVka1MtoZt1/Tn8lsUTxMg8a4e8Dz6m6LbxTgFPlnhmc3HI2dT2kw
D1LL/3m5pJnICUO6lARjVHI+TmjXRiZB6jh7qGZmbLrTwdbVwf07HYJWZY8+dYyZ
hnpT9DwFhUgfABVMso+scafu9F0Kyw5x4TlfHQO+Zwt6riuzWseIxZ+NJRb4mEY2
zND5Ejb24HwZCRxj4sX3jO6N0XFzHZc/e83LjBJqt0c0+Tn7Xlo8FrKTGwjuuJk6
gwmq2k/5pH2FaH/PFBB+vOFoBetXZg09r3G1Sc3bvi6Xu38uVhe3BPca7dzgVAac
7ThM0MGMnNm/9YdKsKfAng4fMlbkx/1HQpwJbndWo2O0LsHBwswZjFFR6Peawmnx
rmNidM3HXJ41xFC7AyPZXdWEWt0QASmjalYLrF06b//fpvm9VF9/2zAvZuOoSEG0
b9iLW5o+MBBx2ClLi7issDdXJ4F2FmbYT/8imlaJ6jU3JTwMPM0pb+OJ73Y5/GQE
lv1IqLeBc75NAlfFsipLNA9PTqVoRFlr1JktHdn7EbdK63ggaqyASFBYwlPbDpY3
QeUGlX8DwByb+59o+DsGKC2pw931MCSDRGxpIVNgooMFTypO6xBjZ0s60zkYF2uu
cKHxcVp57s4WH3G2soM7h4PLOcDnPbj5ekmpQBnyvqcdZyV3aHX6+BnXrkPPaTpT
XgM4j1FAnQyffKmrm43w7uia5j9cTaJ5h1/0TlTkfum8mjCzYhnridyqBPsFj0Vt
m+6Qcbd4dehxgryopzWGPBcuqcLeX7n8CrCGwaBja+riQy0192jK2enQxYEUZttT
J+pgYVamxqrhsNpi9BkuoRKDQ8gU4QWjLGLfvgQ4AkyTo4W8t91gk/g4iud2+Z2g
Ti2kvuRCTlC93N/JJsQjICMcG9X9LXTqI4KwZLLNO1rE9trMxemhHpPMbnUdc3Dl
P4RJFiVQZJOnVNz2vDCH1urkOOKkNJuyVDyOilwVQv8qhG4Goyw/PyzOz7fkWuVB
gZ6h/vD+pK6ICivEwPm5vZOeSXl7rzEBq1cfg9t/xOpPjIG+UOlEXgr0/QIvDw0J
YjKsFY7bHS4wWc3ilZSJecg7wHGhttkWmyxyISG3B2aC5+kBM/xzQDbFTL3NWaFz
btcit0XL+Xa8wbO9FASF+6gV9FGcZ9p8bBVAuwZVrjaD3StRnhfEa6rDOhEFS7I8
lmwgiobUG6wFQSdb9P7qCFeAKeThLh94KrpoIbOjbtV79T50jByAOuEUmQlHVZZk
WQ1h9B3v8OjloWf0lhWVpw+8W9zCrNAPsSRjFbeDrEoYHWK/LOPwpNLLvHKJYAun
ndMUubFVnGC4+4Jz4lrXrDEBzONRKTM0goTq7RaQEFMNVXcPwlH4cSz7eEKe8HIy
XSa8xeECasLXYvJoxYBDPjVM1YN+iCmaJ7Is4SBLuRU1ntoL1eheZS7W9ctdl8SO
1PRZO2ae38/3AqjxDSANz/AOPKg+7+ph1ZLXVfr0rjVDyon8JxWKw3N9JrsL0rhz
o9rJl47hw74n6gb3fyeMCmMf1WScDEpCAoaLg/s7sW6JE+KsQVp1A8JTHi+lfOjD
48YTeWdjIFcU5+hrbUcjUYoGz/2fL2kNVpLYxFSDU3it9eAKQs6HWvSE4RbnUJSL
c5nkuP4EDf2r0sVmG7ytoarQjIvXq5M29pB1py/qBKMnzyU2GalFgUkBhJUDAxBW
QsK3i7fjJ1qoKwqSlpbHgOeY4lKkS0ANEEUbw22sr7fEtNaXJ6ZZ3MHFCWlCVxPC
vYx1xYNdm5jKcTtIiRZAv1OKQRGzs+3yFZcNakHi340ZNCFP3K5pmIhly5LzNPYs
x+jaVOc4wgwkx5SW1MN+YjYiCSjorUTJFGScqHXONXB+8Yts2qN0+wLquLN9K0cK
NFHfe+/npi2kodvMOxy6AaWYjGWa85eFh/dAs8JGZoww3ENoSmcqHya5sfPCi6Px
XoUP6MuYtMyZt4iwE1LfEHEwW3sDMqFbbj0n6WsEwaVpZtNlzO3o+Lql+U7Sj1VD
EX7hVlauRSAHWz9Rm7kOjUMsf8XEMRciT61EXFa4MHyxh36zdBb2ARMRaP8ogHoK
E1xPIhundeqxh0HQH3zYvaMcLSSJn7oCOQ1Utwx9cwwl7xKiNJh6cIxQGk7Vvh6G
yTHjBw7PG2uR81nKuC3HGapS7TdmY5Se/7S63kjdZx0+cI4mY9mORffEvGusBVEL
TzsBrTdCSf4FMtn/ODdAxexxO1FGz78zyeKkGd3Osr5kNByF4ZjnICLzY4IH05FV
VnzRVMEiWwAy81qw4Dc4BqbMxzYfP87Da3H7HM/Kxc9nZQRxe0v8cxboQlr/+F2Z
7i2ir5pJDKVNAmrLky+FBl4xljaEUx5Wm8S5txImdVFyPOkFCG2kItMI3a9rRtml
1nY3WonmeXra61P9Qf8Vra0t02HCmlChcIqaUjfy2RODU1VhnNB+VWHh9v/gRcT8
EcOk9Ywmu0JqZRObyo90R94Q1oXVKpdMFktovp1zCmmq4pf/sYnvAPSqWqZxCZGK
eQnRQSGfMN0m7rtg0pdARgNilcZDIMG/24lKy5Fo6Fdl4dlXC4ZVVr6kaAPaJ/3d
lB7Xo0vNyBx3p34TrBaCXHSmUbXlS+2/ek10Wj6D09NmTwYsyBo6Jdx4FwQ1PfDg
bfKQ5lQyWv4YCsqpHbGyZxxiJvvt6LKi6oATpqYgqar0iw7q79KkmsaT+ULCiOT5
Nku96gCFpokRhF/kqMaKmy8KKK++M7WXr3dB7u+ZWnrEmzI2fiTeWg4zSMsHCzA8
vMAOdJAkB69jz/QWNvPLcZazTBDAP0k4uNqK78tk6Zt3lTCm5h+KvX7V8F7VFzhl
xMwUyd5AknwvieYcSHOFwnOI/8O7h7lSj59Iu+WoYl7pVhyE9kviLio6KHwiWDjv
bigmXbDDfTmXpWoUGKfmNc3s/u0XntJb49eVww8dkA38id1SqwOdv5SQOIcV7b/P
SjENcN7CGFn0XkdqV+5yhE9qtFD97dLLj728Er/ReG4wLWRNkqTNt2Ka39+hMhVg
q1P+TGbekm0/SfGWn7wMf8exgQ8y4PErnMd3iZYmcubx8Rd+DB9NPhG+CSUEJztW
osSWE3em99z6cqyZh2olVFJjfIQCIjL+65ijBAwrzqTiFlfYxMbo4JuFsASdM/HI
VjoQWnvNTe499RNJhP5WLCbDJ0Dq8SVte4d44cjtDqFWS+o0qx4ITo2jyUpHZV52
6bqmHXKlZLNPQTMfjVTYCw3vHqLdwwEnQDe+3o4TAe5KHMXdDHXdfEQQaEdY+81n
/C8R9g7KqfkFghmSE7P6Ccziw3a54s11ESJmrEVwWnGGb/qvEZxDC69alvNcalvR
3Q65tX1MW+AZhgtKDow8XCG21Asf0YYc7/TPpQ2iHMWBb5PCE+xdKgcpvEAJv/2Y
0fuJlhr5Vni4jVm6jxEBV2TCjqaYItai7Q6Bh08RrpEzxmdKf7ILdlnPrg2lAy0B
3Jo4N70/c6FHT2kX6FpA0AkPUmt3ZLPzKDp783H/xi5emP7+lmkza9CeypeP5yLn
Q7WuUlnDOuK9Xr0DAIEOKXqsMRCE28oiGJH8eYmmVrDORpw6wgLwywJ7qUrvSMRt
7/3N7wbTtbILp3c7RHMlV4jqqVFiqIhHjmZkoNhH8sO5DTQnICD/77KHsZF41i6v
/B3u8MakqJ38k5JgRtqc9aCzqzlc4GnklUeUvmlaO42lSKBgM6B8m32emYLjhOEE
2wDyr/DPlF5vaAD69Ug0BXJ1olYOTSV4m7kCDkRw9Slyg/hSTF+3cXYy11TxC9NA
LuTrC196D5CrzQsf+ub9laaVmaHGvI8tLNwxd8MTl+ekmhygsfozGbNcNF7TJOzy
P9vU8UsNbLuzdlpDnW349tFlA3IhJ17MH719jpAM4yAej3MhJvNhYaJ59mIiXC4y
77gS5q7+R3LYWiMgytuf7bkIdhRPmSJ0bfVIRHbho3tCkWG6De/7tEoMuhgWA/Qy
7xAQvp4lN6sL63IC8xTrpxDF4QFGXmVMPByEywtFqfXJb2eSysvGI9+rQMqjT5TP
RAkgY0MqPmoMtEAUsoCFHeQjAcjCKMbOAcnxj+hWljVHT45TlFaMjS0VnkXwU5cl
zeJfsTYg6gRbgrplYTG7TSqi50f0CI3I8jGqNw3tHLMoMrIOOuAiBi2pBBrmqzca
fT6TGkvJeQdntQ/TKDAjZvkFnIWRhHjNpX4Vevaw5hLrSPmEUf1etoJxL7EcqhPB
NDNp82L1QpXQF/bHMzeOcQLiQLnfCR0Q/Tith+nRsnChPfU/jf2toRGL8mF/zszX
XAJsdJfJUVKkAdRAtE42vZc8d6EtLF22S5MaL7t/Z1HN8nVAmdh2liEWR9W8C6jU
CAMv8Oz1CggPjIyPidj1yZ8ujIzR6SZVjLyS5XT1a4MzrKsbvntrpjxXLsccvzEk
3mKLMw77w3BF3vTXTGafWDG04Jb2QRFG4CxhPvUHYcrBxUtVZG+JUXwIcfK2LUsa
WOgCUbkm9AmfAdugEtc2cnbvejhffbnbVfmmsP5/YZXrZg4n6dgCleg3j7g7rCqM
nr02QUB2cMUHYMkjDJBNooR9l9fhvHDQgCUS6FVMyXs0rxoqlI8YYjojkviKjy+j
i4xPSMG6wlXc+I4w3lNvdJwseys1Tgk+wA5V2NCuzBJ9emNYnTnZkaNr07oRgYK+
SPS94D6BjhP9jKnqffT/9+PoXw5Rm9vAq8Yddcdjjw83cSaDwBVdkJcD/LY5nWm6
M07MZHPVvHx/AAUWABBT4fvvXRFlWYupIIQSYqPEgoDSr4W6lehKfugLseOZYBGO
+RGNPgnMNG/wB5JSH4ljkLxiyTZobkcrVmxBlKeW5cqE638YYjuDeVOXWN3+oItw
dA6G1GB08iP7mEO9Eb9GmBZQhEwdkFcLb3BTlKooBKRBWpTEpRttM/dolSy+UPfz
GHJOc2leut6sHMAubPFTCqNpOsNvIwcDWr8VRJMcWspzl7nmFwrucTEJmmrNESQO
o5jG8elBp8isHgDSIIg4HeECUV+Rey2ZZQTaF6yue1PmJuJreMbFn1vghFQ5XwZ6
Gb/M2RmIUeu2/DWgX1DzpnC92sa7aHDHKMYzHMW2+WAMrx5KImDWnNuyveORheuG
Hdj9y2YT2jxyXgCPSm/RyjWfddkF8iQA8MrqXNwh9xaZvoBYtqeAh90GbcShBjf9
feADaa2K+okvVk9dVXFHQzErtDGCMlw56noEyyU/tzd/tVfNbGFTmXiOq92Qw8Jm
ITUN2alIlhbd9gXXpx3lU42qm+kC0LCFih9mr9wqS/ZFW21s56lOp1+iU+tp7tod
atFx/IhTSA7tsHBipJPhqKZoAFC+rU4tTIAdskXz8MxRvlStnRGc0Z/pgxNdiSJm
jTDoGRucUHGuBvOtuKUGf0fEq/TZQ9cOafOR9S9bTvljH9p9CRtXy6+7v8/xNz/U
+T2SxZfNmJQ1GJYwxaLT0IlWC6H2dKw+hwmi0zOCXY3//tOiR2gWQimCGTaM+WGU
37x+0noxErHurKCSx/8zLU+ZBpXN2JPfU9JdmFw7gr5Qfq/TsjVBbOZc2Er+K7/A
YbePNRbBhnGvWmR8/Ar+BxTYCto6BMmSDYHqWvGJke94GpSN7WIutdX9v4j20YO5
wK8e1kLVnTDGnv6VZtiaaEDFH3vzB/z1u58UaIbbIgj2U67tuLT+/6V/OuNuNkqk
cObIRYBDM4sxJrEgz9+R7HuEzBTUGJGqv8BGR/jjPFBNrCpoaZMEAJ3bO2btPUFf
gWUhsT30uLp2ClX3uYba4KYub3O5FIwwKnoIb8WRM6S5ripeKIXI1FUKnSNNTZ8k
QE9+++OaYJPqyALL8ymwftEsb33FfBMWtSjh9Z6Zt3f41B2vN3z7TAy3bgKFbxVH
YOfZ05fCQss8+Rg+Frmoh0j+GINtf3Blm4S9d5cFU7r9QbM51KQPYX/T8tTzYv8o
ghf4DmtpQ3WHTdPGVhf3/HO5WNycjDUimVMnKn1hJH29OCPyAYZWex/KNosxxt6E
KdRwQU8ytRWIx+0ARw50+tTEupJOGPd+Y+ACBX9NXM2rIJeoNhl6PKKINHU+nH4q
pSe8XcRDTZ3qxXfWtb7XZL+PDlq2RasBi0BQ+rojeQBsdSNCa8BszBtN27SXcAxq
IMSoUBKtb8g6trZEONCnJ5hYUELEWBxJWdVKAmWvSmLfm0fJACB4w1E1r0A3vxxw
Bu2qDtgPkW2+0YiVnxtUb/yo1T28zcd+CMYDvO3l6LnDiSps3qXXmr993adrCSgw
IUfSrCfK/7RaweeEG2Ve2s2wa8ddxsJrs9B9Sb054WMWhdsUkUQq3z8BQGGguqRe
aSUJZXdIEJMb0AD/24jJy3iwf5RaKkA1WCCCZbcb1f1QsBwZ173Y+2dnr1O5GDkI
U+/G479DKXwPGuqvDU06UHMeaY3Hn7nRhRCFUDxTD1KOCDMpm1wYantfG8cVco0k
J/QSo+gLz0EpjS+3Xm5fFbPYooVtiCxcO7yg+dx7+9z9RtZLTsJXtR5btrBaiMUo
uzcX+zaOhwvhuq8KM7rRDQK6VAp9MJYaDxkRtrT1JO6JbmTu7o96AB6COEqVLAjb
If7hiry4FjIjUsLAZehQqRsFsaK4A6AQsz7Hpyx8vLOQv460DSfwQCyosepJ8XzK
NrxuftCaPbJTctWkk1smgVVevct4WKbuP4R8MfAAmBY74l7UDgmGTpRsstOA+Oeu
z9TsEDbQvyGVXvXwTP5iiDf7n3eijyq40f8Q4swp2RTblkgbosyFoG0iRptMlo4j
De3BPqkq5WVAjtcoDyiB47ESpw6F+TS0m7ou6Ew0tUr7UVHyMxsubq24qVhC451R
9kGgBW3w1R5cEBaEJIovJC9mNzW8v3YhsVb86tmXN8SoxLSjmCO183b8FIRk1x/z
yaVh3LOoScI/d5uxYFwfIg0BOkJaYdGQm3gkPrUuUqDpXwAzyB7a6//SJNnV3ajZ
MV45Fdb616X8VA4GKTnYm83jp7mwp2H160Y5hDseG++vbHmwf0qO9T09UZ1+yKT1
HGy7VL7YKnazYE3e9X+afusrPgeEQzi6YQPQ55/0W9JsaEHs9TxPV1IFsZoO0Kkd
QT1Del8n3az0uSUFJqwE0aC1O1XclwkfBDURBUAapXuJWZTdKUn5fktZpDkBSgvf
cXT2ghyJBjGPLD77yH0gcebfrB7teRA284MEUXdfvl1UWb9au2OZIVeGmsivpwZd
+kQPg4ebBSdJ1QmSF8TyZGOMy1GQ+liXxqwa9FbqtFrsJCoyh/lM9Zrty/Hw4LCN
cWbaWe2XJkugGAAbXHrvS4ZFazUq69TWEYo6K0yr2MKwjB/dcvTTaPwy5vVf0cUZ
RlH+SMF4TWjEkBFxbseLOxyAr/F7dA46pTAyjyx+6ZR2Z923xrs5q8HNU5C1Came
PJTrAu2oNEjrFlNnilJ2gfiAqB1oWs8yYOk2/iiW980TMVu12y+wXqQuzuS2lc3L
qTweB1wgUz5LqgPD5BUM9VK+cEt0ubZd1OD+VBPynMC9gy+W412hrEtn3JVZxqbI
s/4z9EDO6fShsRxkMqhTgakmGkLqOBf/+qg95Ka3rqwnr3pQJ3QqY9hPVR67bxV0
Nft8ZuvxoUMLaHt2aJVBRbx3Ob9xaWX1Gzve4uDYuEfEE3bnI1VMbBOZEhTJH6mv
OLsZkNOhMtvjn6BAW8mIZhxgFTjeg5VaUK62g5c3CxMsYIC8MrdAWEULAVkIzmXr
oMF/OqUoml+KuksFkUtnHLPlddKFjWTRcJV70mXeGxGrYifSfi537/d2smmveqJs
HeHe7hZmVJYY2ORAhCy5L4PfTmVwbIRhtRC/BzKoAkVftpOf6PPs3AL9pL71hSzj
W19Mren1G55ePXDXbF5M9EfBieacFXSG4b7nGyjw9ExMOKuIKEORxCtOxeTjm1CC
rSL5JX4cZI2jg3X0ELU8FKiDu4+/hi8uUhjYgvsDkeF2NiOJ9c4nNe9eWfo7JnkO
c8vcCu8TrMr49G3pprFHpis7bNkOFxqFKxKxubsidygitdqXLwtznPl7yAO/2cPm
LKHpKDtthomois2kaXu1e/GP4anp1Ko0C5fQamciTJQvsaSLVaQ/TEVNYAHM5BAa
VoRleEkZcgjG95VuqA6o7zzaggLTjQalSLXLwde9ijPGSIwCjsqoYrb2er5XgRTN
72AdD9snNfEHNRSf2wwLisDmhVlZK6+XNexKr2DbV7YejDpwdfggCJaIt0yqlPjR
5v0PM1u3Tl1vEyBr2MZM8yHgn4brrdOwGVkNfqnEnHHGPF6xxzAcU1nlSv3r9+O3
U8rLeKRcyD3Eu5QvVYDgVsElhas5VLLRjG5Ww/mGFRACbZmHP+0h7kX0lGw/7x8Q
sgTdz1Mze6Z5rbcsE9rj91WfMWBFUj0nn78FWz9rNI1oAXjxHyDzjWFSmdJi2wHe
+ajcrmEiB7XNQP4wLqZ0CXONoOWtUpDJS0egwEgSpb8iQA1+dZriEvndRtq0gHs6
b/bbJsnIIpj3hPKdiYsgrihwh7lXsgVBhgfvzl7NAXpFhCnEt8q4SMTMtYqy4qzf
gNq9ZY3JBmX3+7sRoTuCdP4Rf8sANyTE6Lpv3IlrXKNCcZhh5HY6Vbzj+Trq3miN
DRlYYTnAOtojyA8xQPCp8dS35xFXf9Wy25d9StyKD2pS+l0I7q1D7yiE9eQyRUGj
d5V6SXZQ3OKFPihO/vPa/5elOe56AzGZVzQ3XKQ4hkBCR2auf66VgHAXLMH1YFDT
j4E/eo1Z7INO9C+xaQkfjUU+C0nRpqPqnQfvaxiF7ppveiFlL0kHtu9pHDwfUVB8
oGPeepYjMqoEx44+N5l6oNCMaD4DiOZ7C01FW+llekjl5Pm99wu4021RFGSrYW3n
4I2Ugv7BDO6TNolnROrwKM8x6ith0tquRbWD6XfnNzdwSOwJTyG1sXmS0oaDjx1d
20uINleYn9Lb65rBuwKOJDtOQHF+KuppdwkIKNUMs/qoxecREXy7hD+DPfahX0fs
ItA3y2VntfWWdxBVrosJOZmB3Q77ZtQ2kG96BRK4Drr2y/EpLZzzYQIw+VNvrdrK
XYIFIkL6NFqLemAtdqiLqTAY3m6rwztN88II+3v5j3I+s/A+qykzZl33ykqucyDg
b6yPfDOGsMEWe77G/2gtEf3OYafvsn/5rzktJfuNztecKzgKeLc2xz9qr6Bpz7Ro
K3hQskF2KETGtdyXf302FcJb0ksHFdYmXwgmgVp1dCbnS3NvLYJ1MXfhdjixC61T
AsaKSDfGeGkCtvU4x9Jn6Vnuqgr/I1lw9FbEjideNAX7S8P9XihOl1GcaRekNmvJ
yBtBmBF2pgotfM9eMemMB5Q5tnm+CluFXIywMjLNlpMpybRQYWdJgX1qWM0GYx8I
8Q2cJIRCaHpf5+I60sZ53+CImDDIS5q6nYGYT7qcz65HTiESlYltLFr7doc9EFGq
nciZLPiQwFY2e7bB8iqZjzVRz9zotl3r8qhQp7zYxH1sNGqS9Sgrk1sbCzup1AR9
QLXQ3BmBVktfe2w1PJ9dx1hYpQC4El2W4Ao4gHFvy26pe6ubTmnqf05EsvAm4rx/
VNk62JCuPj3k+RvZbfF44YdVf85hyCInpBYETVfqaPuR23XGvM4cK1TBPV8KiMmd
HtKRF5zYoU/hQImusLFvEUwpYWWMAnIUkje9bpgbCtReofyjczdniKN9mg90w1EN
R9K/QlDcc8cOXcYw1FSlbTQaxKHv3QpJd16d7TzsjXjX5RQRD3XaBVumC3c6slSP
zC/p0IDBpSvv1lAGy0QvQsWwFKAyDNWeCV1+XT7HfS86DQUSSD3E127hJBEdN3l6
9yhJBR6dln4wgUhiKuSSBRP8hPKdTCo052lHqkmRr6zkZ8Yco42GONDOOanFwU5O
PcPXi8CqSUpFI5/YFDnM87TthuryZQnXTfw54uqHd3kfyfisVBG2RnisRqfKy1bP
uyr4O1C/I3unxur8Ys2VtrDAdoOQs//pCkXb8Ip6UvIyA+BcGTTEFLYCXJ4D6rlt
NNxzndD90Lu8SP9ifnzsnSHAiAGUThv/p92o7zXEqMcL0xCtizWLJ5gShE/v6KLn
KrvBopxG11eAvaft+syqspBBzKZP6CgK3ptebtFmwy4uakUT3XSizJM+n0Skndtm
3SgGQl2fslZmwoLlc80FTP9sIUCy4Z4O6nQauUMS2XcU5f1ebNaTbF66e9LkTeck
7ToItRTegnv3uBnkfQVof/lzo26nsBuZXiE02CdeiGKM7juZrquEncUG9Wmikzqz
MYU4LSTh5i7Q6M6Ai6agSJjV800X1RFNcoavgpEJ7lXnphhBn9t3PcI6Q6Dyg+Sx
Xp8FTnz+dhlczl96GBBrZ1Blg4ASEskQeAnG5Zo63sHye5V1E/ZDFIxWOQLf2qEc
AeR03RDw2uKlbeKiEccTClT6uS2r/Cls74gG7LWxWR34+kGg83MhSS8sg5mHzLXP
P51o1BCG7JUFxDuCE6XfA4PtGGCebcbfWUIKkWbT9k3GWlSl1/F/DowRof7761Y9
OSXllNpRgucABaaEDcghk+VwEeX5TYi6t3YamQ5I5eKTuoziLekJ0JM8eASyVeN5
X3Bh+tDEnWoZG8cWLn2BTYEuEqlz1t832y4ob+eb58dEnV1uVxe2Zl5GqkI8fEaM
TsU6whKKiwisx6q6yBr1Q4QH+zB/o8REA1tBtFdcdKM2hZN5xAG5eDkgA0NpcEeX
l4jFPmJQxdk7ZL8ErQj0nuWmN7BK3TsYm0wzZ5x6KERcTSBpOxpBNMKVQZzkhUh/
Vtarj6M96clubkM8kUjGTpr3dSujGmkg7REC2KnzRWRtSGOtT8FqB3XbfRmmSpBX
txAZZ+gpupQOEs9WGkPE1gc7l6NLdW6ng9KS9nTYeHIyp8KwamdqC2Iv1LYse4KL
/kQa40wtrI1b+yMaiD0esWQJDMPp3kuK616RgG+5eITrYS1YPHWWyaq68Vfn5o1k
Na4zkcL3TA8tn5YFJdoLlcbPdE30P1NTuBjJY+o2AWqeeE2peVojXXQPorBR0eQ/
iMLRiu0Zz86zwkxbwYlHAiN8WWb/TWiUkzPShKk3/rM4Hi45DFEOsoxeUngAsTXs
fwhMbGUlhFGCbB0T3daRGRfGiPalYBW0WKQ//3bmN9AlZkczsItJgigyCPeiICZf
MSc6/V6ilYp9YUsnqUpiD5ut5uE8sazQPzq661YrvIzt4lMefzSaAfdkP7z+25UI
3Dm/DqKfFBaU+g9qKQKHrnKAn158nUGnrsAQOTIaE4iBme9JbrYsuXxs1+MVuDza
S1kvjJj4rTLb1cgyK1Jvs7pa2AsKNmgvBVNsnpTLHq8tYzty2REPkc1WWUZqayse
6u4zU2y77s33sDsjHGGhMGgWfe/ufd0L58Y/hI6Bzhmy5Xqm4tRnpNg30+cmDGrM
Ep8LD0oIUV0/Ms5CXH6m4Gcp7jilys2At4Ju2hR1aHtZo7FI64y7yeflWaGNZnpg
h9V/3iKS4cmMnYT5gIPVxgg5Ca5RENzO+esY40b7P9/laSYVnmlQygDDjQxas2D8
qOjhqKfdgpgqkQ/Wpyo2OMLbprWG/FqpBhGoIo/3VYCBerE3LDR7q1D6wFdssfAd
bTODovMS7SojhVZ93/RbYFwnT8y1Ih5NwDo2bxOqlT9ETQNZxvrBX4M1cRTAntxR
jkcuRsKvPev9xhBhUhGUuQAbJjkn953I60KDQcd6eH3Fq1IJpzKV6Eca48+Q7A+j
cRQMGSwCFpkvb9ge2ZVPl3tOJMDGLcB+a3gHEG1BBc0/0/Yc5ILwzekydxUkJCsx
m55YazkBwAaqNs3b9kDmf0GqDGJEsEujJ+eQbi/MSVWWvBnNb0SjRzrO4T6TQ3g5
oOR6SvpXaY/aVu6AF2wZjGoVUUtnmxi9B8eBnSpqiJjKEZD/tP4FD9LF9DSqwF3q
Ix5aTo1V8D7wymDdiVcHdvwvBqjGz1k9usp74I7wVIcab/cV7ptHMXdqhzDEF2rq
xT8y5sMQBlKo0VTn7isYH9pyua2IkfAywAYiE63n4y5F+TMO1yJJ76RVDYSmzjVQ
Jg22EzGG9+wjPN1JlZVHz8UD8EsWXVCsPNp1ItHHsagnatwiNcRBgt9gLPqWah5u
9IJHZ91v9vqZQ1ytMg/wSryMdNM87+mhDscCwXy4nUyqO8SDlyzr3cU1fCQCU5Ug
Oo9z5qkUJibBFdG2CuoTIPLrWnL/TZanYmxOSuqoBV/2I8AD0GhJ9PRmvfQ3Onp6
ScMpe262pDvcW7YhZCCTqyls3qJjqv8a49kFrBwuGAlToXaYab/GZkl6f35Lw5Vr
ToLRumRlsTUbQ/4TcfZHVx5GBALIFKG1AIa56G2L23xPnee6iMYZScYUvCoUmR9c
CMe9hmZtm3dCcpG05hakbLkEE662joWhg9D3nrXbn9/ETv/vH1yEwAzWHFXSrov8
O55bqYlNl6xZ16xRt3sctva4gIVDLizhul7WkNmpuVGbl7wuMk9+br+ysaVrTVDM
h8owUp5nUSVmldFW2V2GYQiSmA3SsmFKJuvm7mY/qcYF/otDUpuXZzPshAlW9QsX
EJI4R6zECm0hT4ZKcUpDh02yIaowxQUE4U/oboqpqRfmhtcrBKHU+jsJPZAya2u+
6rWc45XvcLvKLjSVcswYPS7Zz1K7F9cWZQLIQfTlwsMvInc46GLgKDM6Du2sqTQM
5aJgPooF6QCEW+1+y9L3Ny94i2qzp13qiszON5THkvwGbFoNmuJB5UVsPl58niv/
4mRgj7SPRpsM7uQtRsMVsnpHZ4kxdj7rE7bC1oBOBn5UulGRyYemxoHF0YWwgvjr
FvgbDD4e6vH5ZJGIk3xBNQrhzthLr9zNBaetWVi48p1vqoaKxZq7sEvpQ5bQuFpK
CFLa9+qVkZPES0asdtgl4YtszUv/XDPCon8T5Wnn4ynGt1Zn9UC87bSIn6Az1ZjO
MYNGOO2owgVL5ghnMLnlxPEsoCRLOIDYBMcKnHd2/B86F6zinv4rXver6Amy9I5U
k10c5Uf7ctLpqod6YIEqnBr/jZC34NIZD/hWbEuXutHluG+TR8qc+IHwcBj36ZWi
bbnshoScO/esjtBFtY7yv0MnFfVe4vScaNNdlxmLHUkbWebfawIEpobc/mwKoP9/
/sXJ9NZ1cjYH5e6OdmmfIyNYPicLp/Ep6TdkdXK3JwPg1AUVbd4YwvgWlUaNNrY5
tr4kkrYofemr2I40iVoZLbKUMhtJ5gEUkyUiqkOAsY9ZZ6zod4hFSbHFzpGUaHlv
syST6mgIJYU55/25zime0WymWBajDtJ04kEfP97XHrjWuzBeSE3q5dD+jdqdrWMO
XSpMmbelrS4GSMoAqpq6i9HzpNiKan1xPqzCTCmOQIPFfNpwK5h7rmAtux0Kun1w
2DEJF6IC1rT4OfQrNtbAZDgQA48j2va2cy596vrFKrlbo1mg4hjD75c37yLW49O1
zFWOw2D2awdu9Q7zYEPTuH+UtimiUPyR/IwyCB3ygeqsC+7Q0jQ+u9i4w+ZI7VAw
FEWLlK6vJd50TJ/hD3vfd+jHw63iptxetS5BFQHxEzjiGv2AQ56PCvmvG4+ewBRr
zIg2y35TXvnXJbwQQP6bqztc33VFjdlQgvaXqCwe4EXlgsVvF5pb7Kt7AXCPmilI
IwvUjfz3nCzdr8eK6EzF8Yhd3yhn3D5YMHBmt1pNx89dXoq567y6wAj5Occ+38ze
aG1eoSmqRsw+rfS5Nj3Fzb+qp+wexAI/2/4gCrJ0QgrnlzroeQNH1BMGCxpWgvcs
GXEM1GhmgYBrCU/7gzHE43Z8roRMXXgJVE46j6BTK1t2fr2NsqXz9vnqDmoewqC+
m6qdUhDiKK8DKSeVMdD+OJAme1gwAz6b/HXXWgD2DiwmKlX4LMU2IX49EItniLDy
JxRgkmOYw9IC0snJr0Il8IcBBP7D8y7sddJkZnNvTzJuW/4u67uK7tVtG5rMiI+U
1PctrE4ymzNK0KhhSYHxlOh0GTlkBBX0rX4bW+caAcYMKIc/kZpYo2MwWQIhQLKC
yKL3uA5tcUHJgWb+M1D2m98LIOeW63K7Qx0Bv1dTyliO4CcloFi43ItO7Dkq6buM
8aBVFKpnS9KHtmGMWhfXcnpSyQ9lb7RecUSGhTv1z5itLZhWe+Q9BO7dmSYyyvEj
3YH0llLIFG2fvH3usqUgz9KzVFTRvVZ3b0C0kM1J/cLS0S1jOquZ+TPPnxeL5jfP
nXekOTsxtfqXKanU0FHsGhqW2WAIQbeYKvsUOAAkqdIrDpS8eE9aMWdjgAJkDNU8
VfkK6KHmSEPIcDvZ5vG+YaqX+r4+3EJq57mnXQclGpKWNxbsOUJGQd4Rp2k37YMF
CnLqXdcU/yRC+4srPTHJ+dCpKm25O2Eoa5DDwMbPcM5IftPknkiLW+5Vtirzsj3y
py1uMQFouIOx6yF7YXAFXp8s5DLnXANOCladlvltzzusuVbbn7k8b7JhofAC6Avh
zAK6/4AjgQbgNouGJNcsuHgw4pUhYsecnOi2aPnZFPlkHBmJZ3AONUb4Sl8r1uff
ErUzl4sizUHNWTVT9qblWUpZFsJ+XBgqWjK6MQU3qZEM3kuHiS/ODKH1OmeITUgN
7/v+94QnWMLmZ59CtFJXUTvwfgG6Hwic/qUfxz5GxrB41LJ3E/c0JfVo2V78xIcF
q/gvxSf3BnKVlweQqL5dVR0To8j4DFIagSCBKRtRsLhZjjs4COuwd3SiKVkFGAEm
/AKjL863D0v3Fvsy5TX2FR2vVdscqprwb9LHZdlvQ6kJp0bZbFJT8H6Vw7NZNYJR
PLL1hCCTLRBo2eyRxNxEldaTZUivAs+6l0IijRKRsRgOSDWtRsHkUT+f4uNbtsHT
+dlSCfmSPUha58IBYiAgGUVa00671tiuZT504oEPvPFaYtAsbTJiUAl1AkzLJGZN
j1bOcWZMXf3kP0v01XCJ164XfvU01NWw59q4aFr1ByA3HJ+a7Nn0gH2lXVoondi8
0vgvYzBM1M/nqV973/soE/X+O7uUHFyfxApyoXB21AQ4ggiRMuw1WkR1ibMiknHQ
qp8Qgs/AXd2xfevaCFp1ZRoPY9xCxU2hXJ0/Q+kENFY92TW2vNWI7tzk5Yusebeb
+dPtj8oYQUzf41/GSbXV12WxblfDW5DQl9cDQXkAEIwH/GuVVpbm0nnzi99k6WrA
oqGMeywq44S1AIvwhZwFUp9c8q0UrgMna6cyAv/rx4cmwTBU0bjnT/kB+8UloGrG
rcn9FVV/5U1RKYrlkoZBCwzWsuaPN9bYOwAfWDEzGnq+CZRfkuSeIn5R5zMTH+CH
ER1MFf8H6BOoac9oDkR2h8RQx/6FI5+XPxdgKMgnEKYf/3ddHHbNGyWgFrr7Ht5Q
B2X1ilr6cmz8WKP1abbqF2UaeO68F726tBYYtL0TSDF9pKI/CQicb5aYHNqSxzft
cmS1IgFkimnRJlOumLXfIqULtyh5S++F+/A6IZ7X7NxqOhdWTUITii0Nc4DE0xsX
PunvdWThc3hlY58n5mcYLVAe5VK8Qsr0r+Vfir/zpEKE56/+jpNkWy80xZEsqDxe
GFKdAFmYyaY5y5oUXnwgXHTGFTqMr057vazNbT28g6JfngYKMu1EvkFuameDSpEg
o9BCfF7SkuFDVAb4RyKD+2Y1QVThnuJ/q7ogaIx/2Y5r37lOBPpJy6Gj65xBUU9B
z74OCfu0krQgt4hrcb6nJB9LO87KbFcfvbsVhurFKlsWeJgcq6zWde0l7rEqw8rB
9s7Cq6h+EPBbrFOAisonCMJsXJtM9e4T1K+KHdx3Z9BNTz8qCpDJP2umAwJOG5As
Y5/y8ejUKZlPapzFvWA362Wb/8Mmail9NLiyxdvi25wzRlJ78dP6wpI94SruTvn5
kSer1JRJPirpM88QCY8i6MNkL7Plpmr0pzqYIOwvDvHZcV0a734rzpY1NFRKG0vV
TmeMsQYjjkQfPLYqXYM4Q5zL16z+wkl7iSHSAfU6BP7nHUcB2q4jNLl8SGL9FMe4
ON2ec/VwDLGXtm8MKlfmK5LZh4nhn5/f5Q7Yeg7YmiT888kQk/ywV/1nNysUirFn
Xen+8S8i0LqbbNPso21cgKOa7W/bXT/TXp+j/1YcrkCEln/lnlUN/+1En9jbB8kX
AFitqeMB8s2rBpK6JfspI8OkEws55Z8umLtQIvWd7RCGAD7JmgIX+gWy/b1J2U7U
HTP9bhK4vFC/AFW1363pWblIBF1NM2jRMoDZOXfBbOY73PyJ433YeB2l/kVY7Euh
l5lTQt+FnJGdK7Uv+kSgekOsCWcdYwzkoAjVtfqSuhrGGUE13NzQFOkWsbun9XzM
sRMuvRbetQ0OtsUC++aUtfA0IueXYYpXsBSq5iiNtYrAzC1qbHl+4FxF1VA73yXV
V1WKGT6gsIjOwX/jtUtomFkfD8ulFob7eFLoboAaXK4W/zh8mcRlgPgyhZHRHOUS
uXMTSBy9cMX0rp/1o9bK46szmG0sbWiOBWyP+z7NDP+lx8UkzfRkFAhRCL6+TgWG
sCZ115r3hVh4LrAirWlywbmEebaLr3GlVQ+XBBZ/Js+o2iHG8BgZMFwd3OPrX3As
DqW8vX0HOaYj8y4qf006odxWKTbGm+2Nj393ZShRdKgBf4MmGAckpDIaRlgMnqfp
Uqj3KEL045IcRCQRN6OA8/t/BMRcqXww/dLi7Ko3nu+WeCWI9VzLm01UviBbenRz
HL/3IXHjV+2dDzLxKidPdy03ucJbqXmomibpY8BLXAEeKk0IWWyaOIZ83Zx5ZoAy
LyPoVozXE9VTwPwxxX71SJwrPqAJrnsOaDyBBpIKqCu0IL7/WJ5nI/DyOgPh3vN7
eYimZQUNekb0w6nkH1KSj7Ou64qOTOtsJzMyvNrWdjYlWHScYgcxsALmsAYt8ouL
1WIDszIcF/ssAK3aiRGONw==
`protect END_PROTECTED
