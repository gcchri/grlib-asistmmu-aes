`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uEIFTG4kEdz7QA8oPUcLYQL347hazq+msGtnq+47vXIBpHETt8rodvWliHvtmCTw
2+Mv1RXFLD3Gibrob5H3nP+1uEZYffQJiKwP0bqZNyLbEFPtmwcDgttGcCPLRAjL
u/pGf+UNInCNobb3qjNNboZpsj8SYUaRbmsZIq8QqJTqTpMhvcexKfdREOrWlFGt
wd2UrIdu9wud87Hs7Tjd87O1i8TDNkyl171bdFxU8/0MRWG5Fz+xrmtU6Yb9Y+12
Zkgrvreb83q5DsDBKZXV84jktgqJuvDSnPgIE1ihDyp88HCDqLZ+Z/leywFbLlQe
s/LtZczRAa6RWX0UJWGGWKX4qnlkMCQJQ4w6hY7Ryla66Kxbqj1va8g3iiBEgobg
9UHpFkMe9lguwl++YJxCnKGZQL7pa5FBFnpm2IPQT0gF7QvtlYoHPF7X5JLPcVna
uaUgnzNPhi2AbNCFm8KBng==
`protect END_PROTECTED
