`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dv/xgJDZNJ1FUSlTR/sVHVdEj2sIEVKa9UkHDVrFI41tFg8FtNdgFbi7ZiGbu8IU
fFDPHNRTOcQqBZHQWbuPY9dSXY0i9KBuMg7fcv3K+bJZjJvvGDKBhKcXdTrpdPhi
kXUnTRKHqTbchAt2kfXB5aaTi9iGYDWYamBVfk8RFh35FTWcUzbE5wRezMsASxsE
zj9e7O38dgFzzr4u0GjwVLZrKOdtgK25ZF05pR6ycL4hHmz/RaYXdckDgYkKkGTe
HCGZJW5bjTPA6greAwv/YQ==
`protect END_PROTECTED
