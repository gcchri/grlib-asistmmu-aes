`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6C7jXmVcuBKAgGcX8j/oXVffg/7+HCzQ3ZfAMdS09jn7WySd411L/Batv6QEWW3c
P6ikUN5Jwkq+lMXgIyYkcjU5c32+i7sjRFNDbjB7VWD3hvBkTBGJhLaKWkZXXSRo
FyUcQeiIjTJqB/fYs8f4bMyZPsfQWSScN7MbRmDlLZr5tkT9Zh/4GSUWlOl5joqd
TZz0X5THnmf0+xbBk7SvIizyNPFZFCHbpJYnZsO0XPz9bOuxuQAhfVk5dcgWnXOE
28DMIiyW7vb50B4wydX89PF4zidPk6iYqByLD0LZFAuqY1XUBpiimxFa8ZDfqApZ
mYkHFXraR1nLs2dEXGcYAQMdZaopTPVSyxbs82uQoKkKGd7cInaJbFDz9q8Dr6aE
mWv5T8tPDrDmEzap+NXMD4+MpgZCoh4/go0d7yT5oF//Ikmb2x/BF3Zbort3E8v/
`protect END_PROTECTED
