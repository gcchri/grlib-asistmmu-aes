`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TMP99fEZft0kR5QR7iAJurV+e66XoxzrkuPEh72mb6iB3Heki5EVV+M5J22kdeNL
UGDXIrZCahttwjyIyiURADG6n+j8nihTWvhutgcwMPwauTo/wBBaoyc2C4oCSkh2
8Z+i4INn8bmUNxs1nJ64si2SqarP3wHovQasR31dWhUgDw7N6MpgiR6WBKnIHB8K
TW5iP3aUbX5ecNYWvRwKqUX4exWxNA7AHCtGSBpKEebeNcvHDU6BCv0byME9z8ba
PecP46zPZsXQsVKM0RY5Tg==
`protect END_PROTECTED
