`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zhG7ZxcoabJgkllTi9+79cIYpWy6de2PaMwthrLbHYrdVHSC+1cDzCVd1DU2IjzD
dAj/cdBDDBjKkd2ZRJQQNJWijBp8zlSnKh7HM9UzS4yfnXQDI8mBzzai5pnhfhp3
IyZI9FjGyma9d6XoX10u8JvaduY1nFrvHM6Y7J8hpg8u495EddHKOixQf4YWvAZc
HrwpvnUHMcZrzAouEaUh4xZCRjNBTTDOvn5g/Ny08379pHKKs1AUBTt5mqZE29yl
k4jbSjXGMDc5JWDGuha89623dHqBL8Dk6QiRISkDLffjIfoaFWWEJAeHSKJdiD4z
qSFmEnI1KvuPeeS8gud/xPoqoXv/X2F1K2NvDLOgRux3ZdDAGpAity6R/EsFUIcz
9gbpGYitVP5C7yI1oSbKjTdOWqafG1mcaJzDdv2nZ9T7n2qTUzRxPGt6U3MYbqzk
C7JCQ+sFjtIUlJ3/q/yDjY7rUlGpKeKZEwhQonnQkKrf0JXLGrMXc2p7iU1KsBU9
RkRQXFtwCGxzWFJa6Qe0sbTVvoK9UGfOV/F7VY9uoGea8KxGBlfDCiLuBVQeQWjl
6XVKOPLuXuXIo22Cutan10aJlwPH3iqT2JsRxQfAuZWf4ZqHNC3R9l0JY7Ng6IXI
/+XOotCM28NmEoAAhgGmprJH55tk8NAjYtvfIswTVAzJFiK359kQfl7UFnCAJ+TQ
hJnUIaV92CxQLAcx8IvR7HP7C8csrn2Rdk2P0ughGYWPYzVXmgUkSYtnmEmVjXvm
6ZueO6G+w/R5cPlmdtwl/2QBKkVuVtD4EopRF/k0XSj6E7np7+zYH+NqYRDvhymJ
oly0JyH3QWWL0DE+uVSog2lU05w+rdiwEj3Ogd0zylXiDV5bsC5qfbIJO3WhuBOT
pgQeqDHIbityQcrll4+5s8qABKLp/G22m7B3wsfQ3Gxol/FhH+e49roV5rDzSerJ
XC7O5MuHuRU6LjWoxtlgd9RzBpPDAkXk+tLCZIAZfTplJXkq2NveorNpQpjxqbKN
8LUgp2WgwW0AOnDS5IxxxkKAOouh5/o3SFApAxmoJpkFcXeAFoWmSik1u5FedT/D
Xty7b9psUo0yI+2Amuk21OuuTWXXmQHbtx0HPcl2tv/3NNGJ+E5Di6PPvtHavRx+
n9FFzqcTg4zM5RaHmF55GicXjV03KKzNSs+bYAnw6b8Ztvk4ssmDkLGXJKw7SUF7
n6n0ra9VAd9uQgOWQTl0bEXUeW1bMkpJk5CqQ2GBMEkJ/ZDFzmB6FKU2uS4y+L+k
CEMP2L/PFSqgrwU0h+zJTnzXGdROWc4YnFCQqvqqIsbwvRF16HxeduZCVkkenrYJ
vOE27CNI3vAEnEWdtttMD662CaxEHC8CtovdLUe8VnDBsRXZnnL5Uk05uGK03mFH
HTlSfG9qZCPXSKPRZpa0V9S9UQJzbtKySX2MpnJ9WQLLHp/najVNRMwll73sGYV4
`protect END_PROTECTED
