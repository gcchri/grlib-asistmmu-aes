`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yny35ZCWZhlIeysmhSIraNJ4Q3yuSf7VKRIbuJkfrb6aQD6VlD6P3KR+hq5rCL/a
d7CAjG2+pVbjYlDb+XdyAiwfTln86nkBhDhDVYXG/KCXc1Nh0vOX8ueiE5v/ohSv
4j+9DgTZuKrsYYet94OqZE2pzr/gAwmcRtDvPjtiL+toxTgm9/rF32Xrme2uUxcE
sygTuzeuQuH279INYqhLrkFt/G8n9A60X7l9R1ox3+1I81ceCwetBUIInAYjEAQu
OxnmunzQ6+2TjB/zhXcPRzL3rTjpBN9QIRPYlK0Q+p5Y7ii28jV8zYIzBSjnAaCp
exkiepBeuX/I41bWcasHEDEMtmZJcUx8u27ThZShmWt6b7IrxMN7vDdadtbxjOoF
ad5z2n+KIE2v8ESuljKfWQ==
`protect END_PROTECTED
