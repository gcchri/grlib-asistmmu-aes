`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pIyFzaNMouxCIlhUzuio5oFE00ugKZhcQiK+u/qik7+4xproahgVLIDshIx2NNOE
k2DssfBdoeINH9ix/pSYkrMf6SfgimoLW1LBdQJg+xd+DJw7OGyAEBlIOJPGQclN
8Qyp+/tHji4CeAelk5GRGVpTT+OcTfVLLzHMQoCivAknao5SUv3StZ1PNgPBGLa3
2+ktpspqD3VwzuZAqyVsfoQuCCA0SrbBnC5C7iMMDu8e97s0BFD9GKT9VKMI/tfU
lKUZYIoXUp3de4b4H4ApLNaIXQlTpEGeGD4dNO2eWJnOKtC1mzFwK5gl/g8CZ0/F
PkSRnwCtOx/a8/iiViVAnHw3xXdGpJg/E3Xq2feoLOhEpnLHuwhwxQc4lrzCWXuA
5teWYChSRHlME/7KVYInIQ==
`protect END_PROTECTED
