`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CW0m8l9kKdgeFNPHXxu7h411doAjS+SMOUb045iOPW92wgMHow+y644YjW3kyar4
1VLA3nwrSqxN+ZzrxE9e2SEYSET5QSSc69Pl83krE5yiBQIFgH5wp0zpsEKmFHCH
9ahm311P7sPq2yoDS3ZnCLYgveUf6JrkzLjC4Jk0T83HD6xyRI0en/gwVdrrTaRD
Ri2b7se9AykdYvXMVfOoxef2DWGJ5bSBO9xm6o8jlzZmIRFrN1W0rZpwDCMtX7GV
mW/0uuBsioRlZu/ftKdGhDrDANYSm+6k2L3BHTwkDDa9H21HGk5Kw++b5X+OKgCI
QKWZfe9J7ZbFbGfuDrOIYkYxvW3bk+IF27wROu5tVzFCrGe3ZSHrfUQ/qq0Cojbb
0pm0sQ1YPLrF05zK6ce6XoZSLHqstRTj/9I10ohDn3XK6eGnfGyh4qts2eECBNq6
oL/YU7zEK7fR6BpyXM6iqr9k5JX97pdx2oyOchjXDX84nUWYkzqs1HUCpAHoZUK1
xJxnuyD+EZc/Oc6RM1jOTwC/ckjKOdeF8YSI/dXMe1o=
`protect END_PROTECTED
