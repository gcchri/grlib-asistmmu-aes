`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7XNnbis3u290KHXbaaN5vP3Jvsixqsean9XAU3LGqRk4prH/12Pc4NxStQ/q1Kn0
CtTaRnNhOzrAdC9OPjEhtJ3OC5FLioxra3WwSHJAX7l2TK7LKQ6gHdwZTl2GHZic
sLPS9lwg12Du6d4/MAggfh1wfA4xgwySIX1FHE8JuWbjjHio5OwqHQxfj1gkdB5w
BxkYp7htx32BSQGMZluTm9viGLauv03s0KYiZ6lIneb1CLIl3fvyna1BiN0cIJVL
7CtrTbKaujEI7c+rUB+NfDkIXN/NsNBdnefUWflf8PUCdsjDW/g9PssLhc0yp3uN
EF6pYZHfdQXeBxA/SIbii4E6hZJbOlp3T7Um+8pbB/5PjD6mgD/iZFRwXDxJ2DVx
`protect END_PROTECTED
