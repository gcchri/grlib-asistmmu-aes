`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vi/Q1kDaDUcKRj7ZQhu1y7YHs3PkmFSLd4dNnN4X18/z8c0KKxvZAxkICW/mOxyp
G3SDJTFWpJSYkQp1ylfINvit5W+vnd01Z7xKi4j8HaBo02dIVbl0++COv7tf/aje
A28b87cKnvvjca7sSwA3tF3iqCsZmZSsiQepQNyUDwgHFI9kklsHU2Khyi27x/Ox
rFXhZ68H5OFBADgU4jZ3MI/15d7PKtvnc0lZsUoQv7zbzjH7MpMqaKGsT5j/U+IK
WRQq7VtshmcTuXPSDPVRQYeuLSsoaFIxtAXejqmgeVaurSw6IGpD5rCvZLJMxi2j
ZtsdX7byz/6Lkvr+G1s1c5b1aCXj2XNERnOAfbFxSCLPi/Nofqn+J9FXAoYmhZ+y
`protect END_PROTECTED
