`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VXJ2l0Kr8kGV9RLbSrBIuc3Gy9RWCqSCUqqHXNCsdMNnfbXODwHpDen22OFTf/VA
Lgx729WSLORH/IYzwCTpfj17HLGwgNDL8Oy5UU13bGEQjGuc94xE+aKOwwtbfk9q
qxdkrpM0gRLJ8oM3PUHYGS91nn9oT95YO8j5ypI68xzzYgfArb31hzCZu+CHSriU
Tb7W6wqckpy3LmxK6+K4Dp+r3ltW0/gknUFI59ZsOHCLuZYMnWRvzMGsg1m/TuOS
8g14qzmXWfmb/14rzt9NuQ==
`protect END_PROTECTED
