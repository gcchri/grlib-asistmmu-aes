`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
De61OLIsDgXOMMKxNFznbuQbp/xuTEbRzWWrOeTj/14JbCZo/O31vJ0DZqVXGzPl
WV2jQLqm9Ua1byCgiKWUIHD5YwLE/IO+DD6ex6sQq4TNfB354pP9aKkfAdXvy0TV
kqTcDVJYq7L7xUp37SAO522dV0wJob2Y2RlFYl7IrapNA1mKxGKimIwg+Gv3+XkV
dfRpi8f+Nbz0lE7a1NIoSywlsJsqGCdVwT0p5zryH6X5ftwO+yGLu/96E4kqCPff
iyhx4KgX0pBWr+Qju8mq55oEr4tXpCOfe9B3Wok5aVAm/zVIj3n0Fw4Wt+gVv0he
WUuh2VQzNPoLw9+Wv8hQG4o7c80T3zeOxGFDf6cDRQCwJ2CiZGl5jGv+HYMZ0NCE
L+cQTn2zhzAAISHU4mCU0RrLjXIcs5kKiUW49palttDMqb3ED+o3vsaCGgeub/2B
XVJN7FCA/QqSYCdvvPH14B6G7n2aE4vM8OTs/C5h8EGryumU+ZSlQZrJ/apfbHGm
xBd9yvlmO1tsQ1kElX6TlH1suJzRjwm1HjsEv10wFotycjNAfyrPzYcbFdW96taP
YV0jd0zC+uIAAzt+RLMPhmGTkfPUNwQxJN52HEdcyrlQujvF9mWVnQD+MhfvvZ/X
nSgiBD7uqWzPCgF5jb4iXGZC1CIujeO0psb07eyJ5FM1t/jH7VFZph6c0Nrd1uWE
sLFuyMZdxwe2sQb5hqM3VU9TiWS3C5IxbfEJFJVd4/E9RcHvPiYE/vRF7U0caFUf
CSdmWgA0IHa8qgnf4Vwy1x4pFWcmP/1co9DemdW3IRTlewj21rmCkqcayXAc3QOp
WDfTBMu7/YRQ15pphOzQemprmI5EZCL9FkzRShZz00w6rIKt/2xCTg8RKf/Eaobv
vUTQS0tw7dpHae4BugzakZNbP1C5OCS3uJNFFa6w+FImXsk4ZXL9JoCn5VJa1QhA
HzsKXhB0BAoXoorBTdJnY6AKs0Jn5hIeTJ9So8USHBefVcENULn2PmzPazSSfn1A
dajxaFAmTdfjXniG42umXOgArIrJYU2rxWA7Ct2X+CwDF4m24poDW2x3fxcTmbie
tsNhQOd2kGzZslIs8TJ1Wv42zZWnBiKLf2vQ/tvFmCKZzOFDhUZjovjpQAmvggl3
j5j5+ZhkI0JdF4Sb2oYSHobIbvxxMlq/9WKeQLl43AGeJfhmuz/10AKMFJqPYBcC
cSqSlTGlSOWePZ8MczuUKoGUh8NfhKQb3d9BoqDsxlFv55vlaKdWGnZauzqAmK2B
8LoGAWhATMWU4+OKntBcH2YKTh82AbFjqNZhEiLwCoLfC/sn2yIyo2/rwvqcGffn
KJkb1Fi0RXv6Rm8dtreVI83V5o0ZxNPgGGFXFjXKYCtqVJqDzllynqCUIkpLCeoX
GD6E3Y0fnwGIRTurfpBx+RbhU2V0pcFqiVwi67jX2I0/bPnpBTVKns4qtlA7Ydqj
tnMZIoBF+HqxQOHt85FhaOc7kqptc1BTf3hv/nKe8RILmdlgxchzRyo6tcAYC+x4
zHn3gvl0SaA6F2Ow+uAHuVcMvpAQCMh0qeuczpzuL2QPvC9vIKU3NZ1PPHE2RWti
nIyVr7PpOmBgIniDh5XqPjGb/CPx3OkVod4/+skqP6hX3ehas/5nbA3YAVsrj4XG
mP1PPIw+/qZo48LBNwjunsZRy8I02KWTx5RZHBZDuLZdBd1sHXfAgNdLEJxk4YJY
sbZB52Ci4FFs3ZB8aXdh6XZRNUxfgBIkaz/MIrKefr7NZMj1M7xW92Q1z0RDkBWl
KATQ0a+Pkkr1PYKMEXkWWXyawGY5a66dw0ud17gn7GMYu1CV1oAC/vmywFTo/ELs
5f7A3Fpoa1Nk6D0gQwbEENtKqcLAUP6nuuvsroqOUSv1xKwsM07eGGk56nekqF6b
XNFbNhmiO8NWbAjJXl8TOGlrq4TkXTLDUTl+Z7oOGqp92ey9EyL3g73czmbIA7Tv
39Gbgh7O6njqZdRz+N3fJBoQOXGnCO3tQLgzxQi5pUqsN/5C4hXkkQSNp0kdb5oX
fqQcV5zq3U4Wi2jLIBdVcBKR8Y8QOaHMHpgU3Yb0kCxUq8ZhTF92l7UVF/VDcKu4
p4cLp3zHLPYb9L8k2GZWx/edDvVvkb+wNYrQv0gX15TPW+FPw0LKBoyyiOSjEjh2
Ng3m9fR6oYXi3sX3iz6uBqj4tm0tJm3i+cuXW6rtwpYK0W4kDotW3uesAaQ9yz9o
ZX7pJrMggdhhLA/sfKXFUHDvq7AZkH8A7zL3SKO7ueqWLh6ZCf1rIgoFkb91sSDp
7o+2i7YiOiGvu3J5by06QHZ/Yen9euguE/nFLSxivsObHrG8WVYqfczyJ3BHXrxE
3CduittwDm7sfthUiROWtXcH55jLiMkhdb1zr7vynLd/y0KIl4DKhZawaSoVdemX
u87Cw0KOCmIYfJki+yOC+PeoDC8q6565Xv87gqggSZMtNK3wNHqu1plEJcIEV73Q
wnhhrkgSg1F1t07SsBD/OqaoPt8T5It7IR/vGi+HdeYQghqGfYBS3sKCLJpxMwCh
t3njaaEmlyQJdgtbnWN3raKIFVxMh8FwCcbYekosmw+a0XQqC/dQINqW7Xe2KN4J
VXrsTaLI9iFLSebjGnVTmA5o+43xJFRlP0SlrWDsS+vsTVQrjvZqjbMY6w/1Rm/z
8TvG/0dMlGwR6R9J3Am1MGXAArQs7eLVQnM4gO4pk5baTDKW+xaAPj0xKpGMasgE
oZumiZX0YJduPLb2HKxDMS5u+6thoOMeaKOI2ocZPgnoqAE9FMxqRf1ldGDOn85M
mxAc986xh2RVUWjmSCCvtwASRlcpNyJfzotYmFd4ApZrLxoMuPM2V5FDMzmTHU8t
7f7Bhw7HJXBGC04+yE0k52/ifsmkUHp6y6pl6pFbMQWNMLAon4eNut8ApJ4FvNSd
aAW9pttIEf4WPfNExkOFRmgZ7yycLS9KsJaFV8zUop6C7PY8xWPNtZTWwfzOsKRQ
pycB5mbS2xB2jArnWxrJJ2kqc3/FGrEzzXntnaTRz/lo52Lsi4oITEAjtEMhqnno
jci58ra09Bqixu4Y41Tcxm389OBqhjZ1vZtxB6qDdlhSpSLZAjW5rj9Kdx8GYD6r
JgUrmZFjjYf4WdS3mzMXeJ2oYPUkIvoQiQ5AEveehGCwLgdUCnr6FO6jZ4+khqgA
YTGC5xMGkGC77E0+/XVzkbdIAP8x+M1BId9p5uJX8Q5EJwbUn+CQbOb7ADdEMhmG
dYQXvh29pyJcluOIrczNUd6+D93xpJYtUGo9+DhsgklYkLGo9rr5iT+jtC+Qi6nZ
NUORAWv1f9qtW3dxxuEZJWe6PvuLwHGN8fTUjnRDN7cgZ+9yj9P4L3Vd5prUqM29
svFRQV3TMMhGdpVw9LauESQnAY6nRrVutl4UpWSevFcNGpn30SF4J73NA8caDo7C
zENOFGkmduVi5nPnvrCukDBFl748PeB/mbsAupNWr0lUoaFZq4MNyX8fszuwLRCK
mSlXsYm/GHVv+IIb+jwD5zMl3nS5uETe5yT0dhWavbYFhWQKcBpPAEjGfnVXWR0C
iiArQF4In1ORmUF2CNeGXhqsrZnLjGBCZ5oAPZvcdy7vpoRGAI8vqQ0Tam9Z0KZc
PyzfjoXFME5GQ1wriSChdQFyELPt1YPBYn/a1GmT6Yi6qcXCdSJDYWnQrkaqltDY
DPM6HaaRCjLSCkLUBTwbS8uaGQK3/zTHAUZSP/sJg7EavdHaCr1wsE138W4AxOUF
ujv6CdEoM98bd4EjOjxuv9/xJJib5YcH5DyCPHmxweTb+zmcYjKu6Tatqt+RcF1P
A+ZebFXaVYMR6B92dCKMLLSvHUDKVazlVBEgmWf8pKoIxFZrazQMygVD/tIX7lzN
V9jq2QbFIYPMEmFu3hmmAsaR2Xsz7e+qklyJGqvJsIb/dCqBAdVymTrCDaOz6waC
oRmq0v+NiorVYVSeBC0jeIpE95HZGVROOgRLjyLopTiDnd90Yhv3V4zdUa4GLmJi
I40Qj7DwEWts0zvFCWgvBYzrPuNTkosAi9nnt2lPmN1czSCIij9/yhOi5wHDxklC
/oVDjjoA26cAX8uvoMyFg11nZcqe2yjFAiodww8wuYdLJ9q0iu5VMWaq9nI5Enad
FcuReM/IqVAKwDD1alCoL6/KR+298rrBi7NT44cjrVG2J346X0HMCQYfX1udIoNs
INwrLlVzvsGnnWva2GZiaKn7TnWPl7jFc96+cxAgzPF7qGhN1HAK7F3w5NM+PKqG
ytt7kfv+JZ9iXXNWxp9G/bUWaahp6MdM4fUt++Hq/SdK3YaN8rQQGuP9baIKjzj6
DHVD4/hlCBTdyLpdQMr76B+BXqeT0Qn2iKf4k41UFsAujsNiIASGhQ6cAcueErf6
BjkfH/1ZVXveQazSh4HRgiRHaGVMV5bPz1uAmYDN8+MCSmjsjgptYtoOVKe8HP5i
L8o+wWoibz1OM2dc3G97rStKc0vWcVwl33AywMWQHsKJvmXbFKzgrMmiZuClzf6E
PNx2M2gDaqTzSh6Zo5HNGUEcVQY+AKOzBSBi77Ryd4tVKgeQyjnmL8iqECfcvkOD
APee9P0b0RwD/Kxo2TcAN8Q5afQr6BDPnbOoZ0tu2jUXPKt0LehVLEKJ9UXFYkke
lMhNdyp5FBER7jNw+gVBnOoSMRItBNU74CHbWj/qFmz7jzZRfadqBAuXjcVurjoB
Eq8WhgQb9Pvd+CqlkYeGDlSUje8NML5v7qtYpZKM14LJBNGKu1OoE75IVa5srHLF
G/SbOunIQMqOj8iY9lZKIGG4UIpxmyFd0KeLC3Q40bfpuCUWlYbDpDGcYl1NODc8
IUz+/1yLEaYQyTCgNQ6D7pWkckyDUhSjQ+3BQ5EJNirmPAhk+2cSYSROKShLYt2q
SSMhZjHupKznGmVaO/IQuMHqE4fjVoI7vT+D5S0Qc8jtk1Ib3qoNi/2uX6oaIrqT
6vDbOWy1QRkH71mzLmSvJNoXGI5DJuVnW9qW5VbUhz+SFImaGaDo4gRkiuuAqOp/
rJ5hpkL+BNckMaYTRv1haDiUlZOc+UUowKWzGVox3K0r6g7DdHqbxd8S+ZUd0vOz
sGdlBqeHXGkxVqrlAp0Y0wToSmaKgjAUfI7TKhzdL87jV79cvYHouy5Iw1EP8lm1
p/B2wtrqknPSxMlS5XI4crmyYe6WumH6BbjvUh8mYwtHPQVjS+x1dS12lUuVhECc
eBYSM082Xxv9iJZR0gCiaJr8YWm3btMhjuR8TduhImPjWdaoAxFPVcCExxCNpX8W
Fo0ZEz5BoC4+4Z6yaxLUp5/dr1nfdxCs/R/5NnbdpzASW/iYmFlAq7v1ieETpc+N
6+6ui/RP1H6+VCOAqNLFoVRU5jJWXMXakmtfEY92s+e2i4D9N4S30QpvrfegZ5Rx
NNz5H0wb2hhnHUCnp1jH/1bHrjYH5Sce2lmxxv5q9kMtGanGcZ3tTqgSJJosfM15
RO3ALTUA57TmB4M47DmdrdNGTIgv+05Ow73fVdvkuPU0cVVM5yoMu7yL9y7eowoV
I2GNuFZUh965i3jlEJ8VU8NBkDyraPHIk15q+uKQTts4gzxeLF02asswkw0fYkum
WjA2GIv23XoGlh8GASBdbmu089npgf7AYUiAR6yabj8XYYCQUSpQ16K9BdoXR1Zo
Fw9NTkO2ndAgIgpd3m+SubC+T9MaPjromCUyTpyC52WFKm60UjUABa3MGsLTEG8J
xg7lBXuyb5sAix2Jfv+GJNjHs5glJPZyXj7yH9h13nnl5u4A0+JFg1o98QrnDtIW
t+1c41Rc7aO5RWgLdBB+rJiGUeTFtHoVG/P1ZxuQutPNB34E+LFa4fQDUAgqdnlk
oIQGGIgrXUBx2IZjcbxrU+IykomWUNWNSKCAPMH/m/Ij6dIL5GBX6TDjfUIIkK1Y
vGQTRsyTpK0Kiq4815QLF6PLp+YEC8LH3HI/7cNSCwwzFuy/MHhwnkwsAphMWrzb
6fLAL826+y4vYDnyPMkUMkpDwJhdnQE4W+U+ocqB+LNBWq+5Q2jjPuPTw3qoSMME
oerCPufvr/MY5GUQ86DW0waYBuBn5z8sB4PGZY+9ar2LewO7Fo6P6qy9eGxBWMwH
d4HfXNs4JIGtrEtguio8uJ3+ybephhISu/JXdFjRA9Mhk7Fz47JEypjpIg2dO/6s
n3POAtjLw77mW6Ub7WgGfJGU5QGg/pWdQnubszot0RG3QrOTpIdeXJF8qz41QKwO
9i3sSj60fC2G95PIve1VMZsBtOEr0wweaw3mfsIYNWHmUMjUwFvbMp6SwN/FaCAb
xtSb8lip7C3pES8pdd52fW48/b8e7CClTMBcmm42V8dgx5dDoGzFGdxSt8w+Gl9L
Phos/Ia6T21N4eURdZvx5enSH9EYWWEmjjNlZQ+FwxAHeusOQKSGTNfBRyoMwt4a
joEn0GBI1SatS01IwRkKJhaqM3i4/iPuZQ6oGdxz166WJMApvGlplhWAvZNRSPU1
Rds8WNx/uPgzUrfUi45CyF+WIMVosUltCQZBWPJf9KWSDB1KSIYpf1NgWBHpwUph
dgoJG8HPJJhz8U6Ce1K/Owo8NHylw3aTLw1vc2Ef1dDG9t5erAdwVJfzjFIV7Wg2
1+ZEDmbDwUmKzhk3vmI+RTHr8pMVlP9WLsQ+IJXtjm24W0WZCf2sXas355zFMmsx
ySy8Gs1j9GZxSkTlhNPPvpD29RHKYHEryqq7rd41EVUWCEfsnPo59V7jFujD/1ts
zasEJFgo1dYBnORN7Q3q/OFhINeE8RDgMMU0rKwxyDxwSHQkMZtjbCU5e5iHwxM4
2ufZqnC1UwSLjTiOgWNQWAKiMYVdo92drmJz6NoN3Itb80LN7/U2KzBurRCQLLZ6
NB/jYJhZIoE0w+d22/mMf0Bx0PjRciMwhxrNfL0nGfYTKE/7nAuGfx8NZtc+JZjx
mL02LWiYy4q7rWO0UW6XN04u9MLKtK32rT2ceN9twLJEaWuAJljdLx5z2qJL/Gq7
fRm83HXCk5ip0hto8+srrWzOCIoevChx3iEMmJV8YW8O5z3zfeaDMhSn+4ve3kHA
E8l+RtWNcJxZvLqtxzjFpcaQklcQYS3gO0yuXWMJ5MBWq76kIyjhF1aRPa5b5f9f
njcVL2l7p9hCQjqkYHumEoZ+GsBCueN43I/Tw3lW/rXClJlPRPBIjgHKcsBQrdR0
lqTN6jNv2dr2NqGcuRz5woWYj8A36lM6VCQMwVh7h7uBbP4agoO4gcUBDGdMU1yB
M249R+UD3af3PaaTnicsvxjKHDrxVBLkLgxu1F7RG37xY8sesbKEWtJTd6sjj70r
KSV/6g4U160qOAMnShM8Sn0ygtkehBu1VYhWvg8uVwUad6BuH9P0e7E3gAkwVifk
JlcQaE8CRDdmry7NFTFQmUFVUmLVOMZjkPrKDm8YSuCLuQW/o1kldtELZgQiQhYG
1Che4Q9PSdagGeNuLkfCaYpwXAsNQc4fCM1wX0vbfxjEKvCMFbksJSoWfF4wtbKw
fxbjno/Vm+MatjQTwR7eLijas9FAVL8EcGWioN3yRTI910zoEIwW/MDBK071DKcl
6GH3Sx7VFqJIjExDTxckmnuSdQd248RIrs0eZVM+ys7x+MiSsUiML+Zn/io0yo3X
q8sLB9y+6ngNXI867/UkHDxJo+T0Chd/cV9Ks1PMPUIXL1zFBqz7+r9HzSpNhvVN
nOMzeUQtouuQLrYB309lumI7k20bVb1C+sc4xlGp0xVFrk2H6XeXjHxNw5C26ofs
igIw5Vf/v9Q9HeunlVaDyjF6X2uSlwRIs4CPgms2RCgqDE6S7R92ve3vOKfKfHBg
oiphQaZIR9yKH4ZkvjAxCPAKCW9COkC/lLp1Hx3QRzIPA5M8TiwNMotCIx2P5zRb
nX7eVCzkl9uWVH4askJiziZmKi5Rpcn5KF+NxhfxSacaSBLg6qsNQii6s+vd40EH
XGRPKJzhf53qIpY+kbL/jq5L3eBGdKfHkjEP3NEkK8cTSLHPKtEtd6j17OscpF11
Dbp6cXtTfEXIyIbVOxZy7gEddjzwhLEFnMwHf8gQzGaThPpns9jtjPVjQXjJEpmR
6tBUfmZfodvhf32JOa/uXdp59qdA5scMie0NuMrqGvzm5HgPvKy39BPIt8Kg8gkU
nwmIEOeSX+zej6X1bGqI6gDdiiySTyDVaRh/CBt8VVIdsItvVTENSBPdVxgoHPOT
LNQfYaeNKmLQZYlfiH3CEoYGWlu9db0h6HwQrVB+ueGC3g0K1c6wIwSzoMrCdqkK
GGQRBfJR/YCWIS/gmjqGMpbH4cm9ZMH41Xl7covmdMVO9iBMuzHD2TVkLjFdmUBV
F+DmJiqCi6qdzv/WR5tDIHPEQFBWZnPeQZvC/+L+6TmGRrwWSVUieRRV1Pj7Aedj
qTqrm5ZDizMYw8R41fWXKBmVQdOYjrzEOlsYK/Gf/eMitOhDMY+Dqnkpq2qzJicr
LS3+DQshKngdMpLB3r43EPWlFWJK8udQbW7vpMAOePC5UAMoDTj6GokCbVoB+R/u
01Z4GpkSdq7zwOMlvzUO0AJCJC5ya0HOppk8Q+RxePpnyQOjpKCaZfGkRjuZowF0
LBelNbz7RdYj0YwE/W62ENjVIfa9vI4QxUHNiHX/DWYSzyBGTy2NHLeKVvFo/0HH
IGGhkDHOg3sWoCVu63CHu2dcGT+lei4PsjtnnH7kztItHOhgryGbaUQbSKsAMMQR
LwaDUNwtpuLoKOzCEqPQIoOcQEknT2qGHYdjrrCotuCZO+3L/3Rp2pajh2HIPQ2x
vBWAqKSw6+w+qVaB8I2zsES8SgoewQNc2jtFCoX4fauHB+rDyzRhmgWxOD3+QIEd
TqlAaB48wA7ywDuEyCyjGPyCQD6MVHrIexRjcBcYTQ0t2fu7LhlK5Ty8LdrNYQhW
h4dHeTrVPnU3xdcjQ26+z/y3xjbm7EZdvyyZ1t5pprn6VF/Ij2lkmzTiSVINrg+j
MiTcBVKmfFzAuROdKv35v/BwzqAnq3pHsF1vGMQ0g6iDCqgauCRMoXuUoVzpJCVM
g3qfdPc+Wuf2gvH/XO3Y8Q0v3TMOrLX0ITObmLkYDaqNoRP4pzcWdeFx6E74XtzY
t5vuZFBKu36lPZc45ORj1ZjaVINnT3EUJWaZrHR6Ykf+3IDqqFy8jPItCfzpoLpt
nAv7GRlDzNBU3ZPTnrHQ0T1SJOZ1ZT9LKM3llEZTOz65bXla7RqERYDoMjkuXt37
OR7+9oaKLkiKlfSGwHfRkw25HYNh5/HuJsr5tBUUfGNYysvyFurHMLGekk1KPIIi
fSFr6oTMsr07uyj6LSyObAJRg37beogYopnJi0+mo2rX/CK0B6bg4EjX5jAmDkRP
ywGPb6vF7KiDpL/jMmU7tiE/RjYiCytDuw8zc9v5Li0bwA8wmlvGiLZ+E3Qlar45
14MYfctpbHw8He3CIDcPn8oiO+BUJ2gUlH8ObHc9ByAb1Hym3k7s8scvCzYVTr7/
pvOvFMhFBy0rD6MuGWA3zHGr9E/4S1kLiwF2iJFNZPllMVYpxLdiHDV3U1Yoh4rR
GICI8TGC9euaW5MFPoNtHzMtOmIVkIYXTJSyxUyWEhILqhtm3Yt22ZTxwQ4lfXkr
xGP9H6om3eAw4nihGj9agrCa/fDInp9Q9YQePCXDh4sfRXN6J+GoMRXKTIraLpuV
6CNagOVICLDAM9SUGzHSxhAW16pYSk+9HwtZ4930s7mNckzIYNUW4ultTE3tcsVW
MEbl6vCVyHLNCKW1u/Af4GaM6ZwPR0j+hZCr70rbKTKw6EF1oDbbwQT2m8RaRcbW
pQ54eBJzzWo3JLrnzRzwHTPorc8+KBHHYVDySt9ggvTAu2MuPCTdlevl0bZZNWz6
seFd1u9rVXZgAYXpmhuCpt+CgcrkkVzA1+BeaeL6OPDdwt7oKie0InZyAmiTIRc+
mU0mrGZJvWadfxuVq9wb2mXW6qHrrmfQi9IG/PytmmuzB88c84iGZS/A7VO5rL+h
Njqs9MrWFoj6r4K8O83GDp04Ntd3eUwoCCS3IKYOdx2bM4bYJq8Kp19QcR2y7t1g
OeHAWB2LiKV6qHAlzJQSBy3pl4KPcreARvjyXxMsBPDWBAl7g8FPCnT1zcWYgEdz
cs4iCBujyNvmmkCMNP/REn144tIAz8RczLC71Yx0Yqj5ekC7WfZeYOf1eKkfv3f3
jQiVUHn6L2t+MixIqwj0SqAICXrsZnu3uAgWfFkwlIlU8f2hU/WnFP0VEsGiaE4X
AEup9zXwFWxO6yCBYZqav2d/qu/mN8D7SJsElpP5R1JcIs9NSqfp/I1GY1+HPDgf
RKS4SX9epBQPNaBP1aZ3BA==
`protect END_PROTECTED
