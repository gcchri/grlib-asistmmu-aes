`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZIr7SEClmbxRpOEQOnDqc8fPB2lUGdnCPcAINpjKukZ8F70pG6oL4cG2FZNqkf5/
7BCsuXZe30qD74Ci8meduJnLw+9i+nIrhvhs+RFwTUkMA+w6o+HX8K+YBeD+cPnn
PixRiAsf1kIpG3j72+7TqRp0y4untU8w9y2IWisW1wk7oIVIp4IYCOhuqpADaUsC
s0iISA+9nXZ/LeEXr6iEd/t0nJa427WCb2zAJMWhg/hzY84NWBHbfguz6ZSOyv6K
Xe3GCm/i4zL5wmCjfQel8FtTk8FpaC25NT47wWtlMmQ=
`protect END_PROTECTED
