`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rMgruAEuE4/dFPiqJAtQe6VtEuwMPFpZFYfcuiDoxLn2OBei6KJedXZdgiW1vWPk
eQtY7vtB4guzbMdgfv8SniDITKAEwZI1mxqUwffcHiSZwFd3b0ORo5mE/LAtL73R
mkG4hz+cnBOiW0vJFFqYOXoc1ecm6woCdlaCqf+KYdXmQMPOIIELt160KM9vLpfy
j3ciKr8pcBUJvOyl5Ply/WafftDvsjPKa+WA5aUeIXDOELSOFFpXBHDYySp5Rxeh
aN2PPbuBT8BJU2qjiWuDXfHCKorLJ/X2hRbXDu+MZy1UD7sYRB/3hyfjHDpDyyXm
3nwciesTTraXOBfoeIsvl9VgvLdjRBqFPXKc78pAm++2k+HEPf0Wx6hnEYd5ocxi
hnkqymzzg9i1CuH47dM3aJbnz51ePhVY9r5sAOczdej0U6pOjAssAhn7V45GGmlY
hRfFcUI45FGF8YDOX+maohI2SOj2LaksuufQ5oSpPnZxdPztSc022xcSlj1OfKQO
meeax1lnCgL7quBd4iiIhXi9234yeKFueO8CmbTfcqee21UDcIFhWv8CsGEuzNjN
Ngo0jtwA4YUlLJLT3Z1NyTH+thT3no1ExKPXTC7zpZPiC3bvglLpsgh7lcprp57R
KZgl/vuQmi7dpkqYeEl/zg==
`protect END_PROTECTED
