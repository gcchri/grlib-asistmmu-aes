`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8cZaUqbl5ImyehTOVPY09M3bvJiE3eLQvfFB7LV0fpxCxAl1pJyB1vrvHCkczn34
e6zo4BIiXmCMLeF/zRX9pk4W7jZ5UwOY7Fwbge9Ry6vYIDWjd5M4Zj2eCkED4CoC
CutJsxIPLBTUkTEs77GB3p3LE7STTP1fzs/VwLBHcEmf/x/sW71GTvpzrnBmSkdP
YA9s2sX4qj3q86O17WBGv2uDnzOgw5Llk5k1WYhaUOZ6FWJweSKrCQ710rm3lFLR
4TnX/1dP6d+ZhQJgSRcGPQ==
`protect END_PROTECTED
