`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yw3HppvK1r0NNy0CgKMH2gBFDL1KGCjWXnET2TtlN7HKVLXtYB+I0FinaFdnAWP9
w02yFRhPVQ7fK1r589JS+aUgen+NU+21O2Jm+8Z90N3feO/KkwtwoWWy6avF/sW+
E8pbMfumFwqWMI/ZQFn5crbwM+4mRmlm3rT8Yw10lFZ5I1r9ieAj+iFlfvjUu63L
1jylq5+sXqxJwb7Riv7nKgSjv0XVRxGakz5WYecjgnCCjEpIxz0xcyXh+k3qC9Yn
MOS2mjNAJ8/hKQoo9oZptYQP2khIzKsb+VOVYlmbbvrxfOeq18UQA0kl+1m/CuuD
zefYFK3DUX/4W40MTNw4p9YcW06nJNZwIIBhqoWaTOtdFRXJaVpO2yTxChTQR10/
lcoAqnjwVd01e0lBDym5KNqwl4OYcbp8h259cwv785egihy5k+m+0g6kYSfsNMIW
JzWpyFdRhIGjf5gGc7MefO9nAmAavspjzp5dYK1OivmtqyEZAIG33dJjiHGBmGrD
`protect END_PROTECTED
