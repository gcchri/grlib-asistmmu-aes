`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eOSNMmfdKIvmPQ5HCbc6RaXJuqwE1wKXVCBLRRNHxvrT5DQhTVkynDkWM7/sKDwK
Bv514wvOdOeREW+LX4FUPsVeUrU+Zy902InUCEYQ3Gt9j4XgUEXwRI8j6zsJTxHU
KSp1e8klNzceBKae0XxmdXcVcIz8JzTCedaidWk0TCgquEfPLxMihDnYjOcz17Zl
/NKKOa+qCZ9Te/voqOHOvfi5wNQWCayPu1LNi47bQdtW9UB0HdzeTFPSFj5+JDLu
cRxO8iF5YDL/Z6Tjb3UJzpSKnZNchfqlBjg/gbg9iVmYmafRxMaLLLnzj/Ery2Sk
K/1L1bglfPF9rFh9x3uUm+7nirmGTZCieekycRXgSQnjQbIuGcqx9JAi2CG3bYE5
QehsaBY9EIkmlVoee3kVlD2ldXUxAYe4B3ShFVQvAodRIv0lKnNNA0xlLctEb3Oq
FEaQR24z1I94wpJ7JDdIwMGsvXAQom54EyqFgavT/6csXZaDnbpVvnlNJHpIi7QM
QqAQ2vSh7srlcFRcwJkjbJdbZGGB7H9pqJYCkCEIe+L91LXorHeMTTZr/tXgHJjl
3yHuA1/v4s3SfcV41600jlllcaVSuU03TBozgb5rqk/AvO3pNOL0WyFFJJCEJbgz
`protect END_PROTECTED
