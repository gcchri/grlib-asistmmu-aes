`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J3QKu6+FDlhRZnOgLp8qtzZMkWMknsISm4rgNGaYCliU7d9zL9bukfzFt+1qTp/D
JCOQymmtTVkHZPL3ZBJQsolo4LlD15wbilZWyw3p/oMxF45wGnDhZmzTPbUI/FSy
HRrblpiGVt5SJQJTRnOsFyFupJyAIWNGssiGROuA0Kz8g17u3QjFIi+zUYnmRoAN
bv30J5ENkJEmHdp/fmQWaasCAYU/pe2+scEksR8NUPVjunWAbFytqpMTSPSm1CF7
PNc2QnawYno5BbdbZu5AxheRpVk7kMS4Ci3QlaDWidtwdgPY84VIBvgkpgJ58F5q
yyqZY1EKzyKl8FJPtAvd7QiREKb58Rp0hhyaOn3TtDIgkBld3n7OuRxM/G5CO/Tg
+NXpWaNiniW+5hG7Rz8NW3JDSwZ746hIhtdoQC6ggnDTpS0L4Pn3FzMbHYBtVoiE
9POxjlcgdOydafoW2Jy5ZSyGtnr4OSzSMY0g13jwDM9ItdgBpCkAnoB7HUXzF/+H
qbeBkmdfvwlSUvVbHAnnHCizAT2nu4HQYrMf4TCjYoshJKcHCDMTR/D4n20q+QrG
iIeo7zB/DbBl5Amszw9q1V7mNgjCGpqL2AXdYbWPXg1NQmEaxqAFmCPcpTu6svbN
/eeUywuWWDNbhoaqexnsN87icu2m8k1pbrg7TqU7niAQBzj0y+iH6atI+TDZXSkP
aUiPHIbVCqfxiKKZhBXprjEqIzdvc0gzIS6uNkHj+8tEdPElRLmpP2ohL8mC86jI
9FWOn5CV/jPQhe6AcU0w5nyKA3htyrqti6NY1in+eq9jtdHtYoLCxfGfaAkYfdke
H3wh5GmtZb1GrHNQdOPVCXK8SieDn4m8YGs6aiUAiAcVZLhu+Z4GCsHlCJsQ4whr
oeXRCFlsIY8+HdIaFOdNWXjuDTLM3EyOjbgZGthy60+AVpUL3Y6ntZR+ozRWlGgm
eB1Gki5FPtgjq9+MDkSqSao89uG3PbLKxZT5G4ztzUZXiz6hIXjmM+YXOFn5nkO2
UiegyeRY+3z8EvWzalv0r5PUo/FD/hqsvR6OI3DuzWyv0ZkzaLBqt4FB8jT1599K
`protect END_PROTECTED
