`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iaH8UwvK+8wLCp2YPdDguDG/9figibXZ/H36Fmddgs+o5ST7qQ059OTuegRg58F/
UYsF/TFZoGW5awu2sUpY2nki1z1+kK0S59xyJgk3Q+q7+BJm7n2oQjH6XWQ+PzRd
kI6C61A2ZAeU5iisGERMlBb4E+sbrcp1+yxY6252fGgWoYV/wP1FbLKuZP+wrhEj
uxBNLogpjAsObu/aEYU8KqsayyOSz+3j2QLKk3/tNorPPLoVZMc1OVHZl92dIaTE
293upfpyl2fPIklMX5sQga84Xl8WEul0uiT0R9pqU/awHdU3sNO4PirN5xfoVwbY
nd9VsoTalIMs/8YwcNkHnICL8M3J2SRckMxr8zB/ym/XPC4Hxyvl5LFVArCsIacD
JQH9C6oYjlU9iQxC0wWi6sR86k/AYxFxSiJc8TQWdJcsOTudlH9ZBEA3aOlrQQKK
W0S1ykv2UAel6H6Kak11Noe7ESvHM9xBcaOib3lyQebdX8EiXFyNRjNccmnu2yAF
p21tNvYpZy5V2FDz1+x2cxkmwIg9YapMHD2znnnQCrOfx2Q/YdIveOS7v2iB8ajy
Lx5/4vu96pXzENijIJTa0c/U1657SBKUKaInu8eGp+fzgxlDMdv6/0fZNkeKxv4W
CqlRuK6I4NPTw7TcGt4Q7xIPae7KcLAhkX/VhvoEHe/mLHIrmPfXRWgm3y6MHiA3
EgCo8c34GnCkwugk31aaF2VtJEgPv+1a5B2Fjytkog6BKsNRntK55Blx9K/hddgY
1nCXat2MvROswLZ9ImnOsVOXa0hUwsiRvd52g+VH9El+OpRsgKEKrAlmWy5putlS
VZCNSdNoc/KlzaoGQmLnx5e/jdcNwXTQVR0FVrKXy1cxISxRh4d+AXd4PjG+Fnsf
hZfssxRhRPyVOknPPb625BzheXuqK/IDF7FuO+2A/+ffI00ifNUMONEyc6sXCTcY
nTk/UD2/q8DMBCfaftAmTnaGKhlBu+pm1GXhWbKis20=
`protect END_PROTECTED
