`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xa0FtiqO6KPZHPvdTyJYeztjFv+/NXfXv6lTpbJ7DlJMUMYaXRPcWloRUvr0UIds
Ozq5J2TyWqyMMNpsgks0ScxMfFdRnrdZMhj/sYXLZjoQYKXCG/wJF6FSpNI6bjUz
qFs4XPxsN1HceJ4QCROVlwksas9bJlwJ/Ybwj5VYpA1y584Br/dTXkNAfyCLqT5/
1DlmVTCeLkHCPeRphC8KFP62mrf1MGGni+FrCVCCsGvbLvbzTVC4xsK2bvi5759e
XLohv9Cql8ovf6uPWQZ15609Socw2AcYf4V9P30OyVLBclQj5ivtUl/4eix/554v
PqgWqQgQGo5y9aTe3yU6Q8U/+e6YTcQ0NUch0c/kJLC8dXhSqNRE61S9jAh+RmfZ
ObEW1epze79tcdyFFjzLumzVU+gGkmbMJgbMXDX3mLGP0zgcGwI2k5JLAIDNyQpe
rGasWkdZmAeIJ8EMcsEn7JYj3H6Y1ay9bJBxFXw4Jg4GN9fz1827Wb7tEbVnMFb6
RllmqsfXHQg1Wuh6ctkUa5KiXVwanbMA9W7JqjRPhzK+Bc8QP6cCfeAzro9qxFt2
HFjHQ90WmyCd74iMS24ghKm6x21yquavneuVwhI2lftA6awyGEA9g0kLC+md6asR
bGO39iDOT90ESSPYPhnde16gIBCNOUm4/DPtiyBJqgkwC0tML1e/jMp+9tzppivg
34Ypki6dQcJBy09mMeCgOqXKnD7VgUaF53ip7lDEI96AgmDyrlg+E28DF+3px1hu
ZsbZTiXQWrrQ4MwMAElbbr4q3foi5YsK5Oo/geDNQZAmnm1H4mBjlvVblwPnn9t/
YP1Cq2Co1bb7YZF8MBSOb876jYB6WrbKvnoaRHdC8CAjQC7XoPF8SPQYz7TQ6Xjm
Lf+udCzSBzdQlqYieF0+JBLcPNZnAPN2JhJecziHfpI74pDkxZ78NZfZWpf/G+L7
h/Wnh3/gIeRdNI30AFGasiS3gGVfgHaUeWFNeivDX42SI4f+8+zUuHlv1h6uh2Ec
vQvcRkad7Rek3+eCDVWZYLG49Gi8qcXg+SwRjCQfOauqKkYxbI6c3FVgZqXrZxsz
8zpEK96vO5OQa2WqFkPArxfj2WaMAA+U9QpGLC3q/NgW9qZdCuEaiyWziTLFIX4K
z3cxEWzmo5CbYqpp2LxHGB+hOE7L6iIzrsDz2eJQsHl88I/XvAJlmx4tx7QZQGWi
J3EWksyiqvZsJcl2r9bmLVOKNs0gNYVai9+tIjhtBTlqZbx6TUUrn+Txr4g2CGsD
YI6Q8n3zlDSaGwkIv+QFnqyCXG67Jws2dUVuf8SlAQV0XCcjMrAaUzzUBFLdYTnx
sFKS/qyPIUBKUZMLNeQe6yGzFmd5r4Zgs7y7sf3IYAHwJP0DehINZ9BNc3ubiRBR
EteJCdf4wqbk6+w0myWxYlSuZeCSiqkwmFQ/T+kfJj8rqvDhaZlqHrOWhbPiUIRo
6PcZpyKDjO5QGr21Yb912WKH3CYAPP0a/YcAgelQhFFBbs4EvYNkQDWZwb7XIMKo
wZNajwIq2TNdPrWnbDEAo3f0Jpc078vYQVleDq4AUHA89hbafGEXxrUQnDy/JJxt
Rg7056obtY21B9Oz8iLtrA+R39pKC+5Dd/q8CYyspKPiWhRWfePgO+rdWV/Y4FUh
H1XQetLGqrJROa4E4M19KQhNNSIrsjxHhn4vvdp8Ad8CNjzJ4rRYrVaC1YZ46pyd
+DLl+4o094HzlzDqlbtr8sz2ZV886Jja+HcBInNMrpEggM8zcKEOqrIgKLcvsCcQ
rp2a5biN2yevHGA9UXrf+xxUYUOhLKixHwgyqvP2/xVp2SGVqYKUQ32JNB79Cs6J
9OcHQb47+SWSaMtVox1ue2frJ6/h1Az+glcscepquY82a7ccXCcY6RsW+w42/npE
XZu4YMKv0Xrj76oO561u3/bybGi/p/C5adOlfSLZ2/M+BixcotLd1xmSEzD9WS4M
16UelySPiIKueFUcYXf/Pf6g55m/RmY+5GMzCjYty7fNXkxnvd5yF486eiOQ+KAP
bvSP6AIOuxZLc5eGkLUxkcHEoGmzu3p4FL4VSGovzKDPXyVy/vEGX/5rmqLarJ+f
lRIsW8nPZtHmrM1W6gfajCGJ9U1b6LwB0S32qbuH/MQ=
`protect END_PROTECTED
