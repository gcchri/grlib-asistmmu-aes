`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
faQqayaI/SZWpQ/wKAKlCGG/wG2+OurLSmNkfOfL9F+1ESeDyD3t2kbzFlgByQeb
famAVp3AM2ReDVg0FHw7GTxU4IBni05z1p9flc36uL0mdzBO/5BnEgBHAfTOiH6J
3Q5QMtkFpJH1hA6ckqQtIRe633YP9hMmR9uIY8tLotDjuUsg6Ybo5z2o58coEVC+
DADWFnzc/3zqjpB1RyNnC1F8k2kHV8lt/mk+maTu4KFmzkik5nVfLslnMMXmrmkg
AczTsnBE+WPjNH2TLYMupZWVuAkaaN/TPJ/07kmM1y2BzYw5eDssT40B9yTKhC34
J2wjHwL5wC8jWrl6608FOoVNXRlL20YlCWwGa1ufyWv7kx82CVywSwqOw4TlgVEJ
LOkKjGQOi3v9NkWMuL9gSVeECAHPu0HRPdTsUfOVQ+WTWaHjAkA0xRdOefkq/UH/
a7cRqc6XTUubfpn+RcNdRe/TlpZNKUfW1cQ/dW3fIX7MjfYr1pMR4K4xoA2pwZGw
/Ix1qSw/HoDIrHJhE1b13+7qXtwLKa4aWGzw6lLOH8VdistWC93d9ku/y8Ae7tLA
YiTDiRE07z8pbqMhVXr4qtRaGaVlh6j6wxnjtSC3AuXAj8B0QorjpocStppxkOAE
DGVuzZ9fH5K+4eQje6dIXYg4rNAelg4y15xB7i7s+gmwRSp/o/rQ/TR7FBWzZLct
+CzH7UF0zDRhx5LUgbf3axWz60svMko9mxPAjE54k/SiBTjlnCSJERl1A0jOJ5J5
v2zINQavHAKcj0X8k9CYIPo2Ez20Oy9EZzOqhGF7xg7oF3uv70jGJMA+oUzcowPY
IKKQ2KXB0R5uNgu606jA8csTVjqlEOeSS/7rcT1XLqA=
`protect END_PROTECTED
