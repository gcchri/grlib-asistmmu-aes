`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DDb6976QznE++zAI7iybM1qLNSq3YF42qXZ3eEsJ2mAwgcFl97hGsrOAd+//G4yQ
WWyRNej5HURZg2JNsuslf9wNW1jBBRemB8/Y7/SKKCJ903p1Fhdl+gU9/IT+2bxR
TVmeh584DyCHbvWfwA4og3pdngg93/kx04DFWXWg/7bbZGa+MIm3Bq3rh1ohc4Qb
Y1ScrF/N2IKc2du+1twv4PhTsJjG3vj8qrXeGfMcbwlg7BkZmRrkRQ24QxIoOcWt
RP1jHswppYcecFwsZPLGW2QtWz6E6sA/Ulepn+fFD8TtNNTiid8iSckn6N9CSrJ7
FjgbhmuK/iHCi/NFJXnYeqpQt1KlNZDs35W3+GwElXidrhrC95zltEsdQn3PkoCW
RrNUZOugli40/5hDw47iz4BPZd3TQFbLKI3O3fRBABXybe4FwyRIlxOaqPUbsjFb
kjqogHw57R8o3JGIozZ7X24HoSxok9kryv1cCTKcXvNqAx4sqZCzrYE9PWZYsS0Q
+0lw/87bAEgdaXIoM51norlPpzxMuz0Eid72fNE1L72eh4V8KiM7SsThHwHTO38U
jCdV3RqbnecClno9vl5QIJz5AwsJoIJBeVG7ii6jsOpCNt6I4YlvOAovipBWsnQH
txDwjHJWNScBc7nERlTbiwuDcvOQCl+IrOxegmyXtmE=
`protect END_PROTECTED
