`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wTC05H0UX9QoS008mYWcJQdNZWe2w8JLkQz6ZtKpnKZXaCA+vHqXneeocAr+JTYv
xgypFQVDf0nNHE8TNRiGurPm0wpwLVyemWhNppZ64yWq47nHLrXRxiJBwpM/qjpi
7W8Wh32QxXR20j1jy9aOnHN7VrDllOenSYw1m8pOhA6tB3vY3SU1GxOr5TyfdrG0
+RBxOyHPZ3mSVXFZhYtsRyRhdLVnmBISa4B4mAEfZbF+x0oovz5d7pVxjnJmGBsc
8fj6ATF5BjRcK+Mm87jW1OeQF/5Te4hnqdyEG4jS+Z0JeuSVWBJ9okfwnv1XX0Yj
DiTvC4pg+48oYjen2licy8T4Ixq0Td8hbAcFJrrVoo3/vtWIC7IgvxgbLxgsfGa4
e2qyGqQl1Eh87mCim0BeUK9j1wBh1mOJ2iVgz/vTOfrf+pzz0GXE9wgB/BovtlwY
3Vfjjx7POu6C7dQO3hn9MaHkQcIJUHTOwE7ddpwOOCW66zlRIQsdu5OtMqZKl5hS
/191qRzsZQWFgYj6aL+s1dKPIJMDNxmZcAsLzlCh+hF9c031A2PhKuJxJGS/c5kL
nOQBSi62KIb57xQ/mfKAVORcFtTAuv0ZlEezY3iwluYFzMTb1cPbpWDay5yq7VEv
So9qoBxjPnqwjl5wH5ux/HJBaYS99SZKIDXGm0GijStsAwbOvoTrWSoLPDdmPw+e
x7i2TX6MY+Ov0yjVjRvdYhDljrV3URnGrjGtosFgOaIiH02RgBHua1wHCiL6UjKe
reNlbhxGpuMpOuvEEhu1+zJX/VeRE5usE09lASy0ezX/if0D+Zi0baMBJMiS/pD1
MZfCnjqVoUkd42+MS5rsYY3/+lqoe1UoNWZ9zjS+QCJ6xHC5x0YKWPWddjgFEQOx
zLJDV1oar86r1D9+7qQPF+J7CuUrAy+oviZYUG3BuGShRxORuzVFI7m24WxHo1vD
1FNcmZIjn1q2HB7Apw6eXAcNSuFuRwTzkRi9YWlBGylgCaH+c5nzLzVOcb6/KfU/
zp6lBCoq22eMhk0kmgubv9+s9rBd6GikwpYgSR0VxafziRw5ipRGoS2u8oW8HkEt
BZc41BxCsDqIjl0yR0f/2zvI/+tHAOb45QghHSIsT+NslK8KGb2YLP+TmrwjQ4/e
wuvvi6ExqRgJBw4yLtFhdcq1YYej7GNVlDAT5UuySgCNN8tpR31TQ2doavK9AaRo
b58gZ0hpV+afFagazJtJZD9iiT9nbDKbWInsgyohjp/qYEFll7ghpLOXwI9GNckw
MjfAFhjQ6aVczflg0xc2BisCw0NIRPR3lkXrplzzLB9Xbd2esXmOehfvgLeZa9l+
MaeF2ci0Q89vyujgWTxEQX05hlagjYtvPRtzBOV0Lfy03gy6ic0yWP41T35fWgDP
`protect END_PROTECTED
