`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XfuImI0QbsrjNo5UYV6Xh3lPYQuOJmEvYjoYWFjW+o5/s4jUquqTPCxAnWce6ldI
fwk6FO3+7n+zs6JpLoRDdHB+aPRZaBsbsgl3vhqs/QtYSRHUeyYp6AotM5CGo5JM
dRqS3MRoyU3BAgpNYGlRroZSZR+IlFn09J+2ZI6X+/ugpNMvwSGtUINo5idJxHRI
TWd9SCyrLfnYDLofaTV8eN1/VQ3He+JksuYa+F282jYHNvSiE9bl7lOL0pxT5qB3
NDKvBbEAGe+MS93iaVtLUCj8pZ3iAEgCQOzWw6cDTfOR8FI9QhWqsy+JgZoFKHNx
0n+05+6bbTCw2yIdObqkSJC5q7G3R54va7neo18rXDNw+c077B24i/WS25lI/aby
0a7AseoyU6l4betEReRurA==
`protect END_PROTECTED
