`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
crrmHjOYpFmXNedUp/+WjSl7qUE3/Ao7kpjRNUwFrTTxqrz/K/1JexOhGUim3VzZ
E2NFKv5UajUugbboc/kR3z5bdWLPL6El6aEPgmjoKkwl5/GxolQE0g23mg3ScISe
3+oS8xaI197mZZnurqn15HHU8Pb2soDGzUE9VujLMkLdOELIMtEYOz13Y/39JlMc
sCn6Z7N+E2b1oHwFe8Wk/bXXw+GyzPfrx5EyopGd/WDyEirrdZdCaQ/5lMraDeWg
9hCc32Spk0jQUYCfkGhxxkFs84Zb1zIeWcit5pM97mc=
`protect END_PROTECTED
