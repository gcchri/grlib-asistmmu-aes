`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+hrkhRvDgrjIowu/QpuKKoHpcb3hBufcmO9F/Lysb9sq+K9Pj67wZHZDb6/qnXA0
iTS4WjbQV3xmnW9lyT74lUqGVdUIwNzCMcIDQRSYH8Do6DVRR1Z+ieXIGl5ISpK+
voMCxzUlW5NeSN1+58veZgOSWtrL46pnzd9Sq7VliaCnl5kVig4/SOEQa6o1eSzZ
HZaoFYLclMT4uYroWttm8Q==
`protect END_PROTECTED
