`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jJHQK59iYiZqL2o5wopZHDsiPHRaanYEVZWW7AXXGYTyKnCsHx5dUMcFj70Fzs+r
ANBDAGNcbaFeq2NrBYDTVstgSnIKLOgxjQI73ILwLRUOjzVUA+eUB54hG2MzaPta
EcEP/cUxtRKkSpHgFPxPEI2STCL2ihtE1N6Aog9/iDFswIbkirPwe84t5JZTcDgF
iF2vTRayolqUEFiC1U3tylElynGcj9h01xIqhPcWnui2I3zi27mF3+01S5jldRvm
Rs2QDW2W10+Hz7nY4D36wLv12pyr5nK8xHiuZMYZLsM=
`protect END_PROTECTED
