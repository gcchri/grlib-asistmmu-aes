`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mKuA6tVJsbvKCD+E2Rw9HmGwiijGEGATLDeoYxppy972MvQZnPjAuK7zE52rPjWp
XUlv2Tfyk5cm7IhNozN3BjQmp48FUpDHvFjpOokO1D8gGMOx+IY1wYm0hxkOvMwN
iQK9kIaFOKWYtDTsN4m57RNOkqTY38dnab8uAVBhua0MqV0lAOWluor1rbIGFQsc
B97kTiWiPNw1nolF+BFGa2k4xH5p67eEzPmEaDoLeCJWecUKgr9sKpZg13f/m+P8
VhWQA7zsm98sMRC5PtBUH2kVsEXpz8ttpV/EwZ6eXy6v+XKc93xYIDGCAgLDb9bc
xew0Fgi8dNCF7CLUPnRqh15vuPLNTd4+YNRfRxrsFpyOLmXrYPaUIJ90zADOVS5p
0Qwx8TnahaSPW4RcU8eUH7LbiyvF76eSerHa55fwuxTofXuVV4nrKgPC0MsTaJV3
91ReA+ILpnjUHu1zRWGTUTThfysJDidQrpv/mbMujB5lnwW64jCOQJjJzQWMNjJ7
l9mmwLQsUlB0ypG2ZUBhkl7KmUcyBhTTp/4Ptw9mFV0sY012e7m+cilMYRT7vkEj
B6DaPhoQQxq0U4EoxckeGYvDMwkjs5R78JEzBe73OgTZZGMEZ3s9QRj2Gr7vyR/g
UOrczBumky/VsF0hz2l1bHJaZFfG0/IvN7KNXfDPZ2Kebf2W2j8EqfEKaVxz/xoK
1K0/uhC9EuyP9pJhoVDoZ5pkb4rhHd4+Mu66xwIXG5+1GDVha4Pi0XMNh5EWI9Sh
7ENl3UJfO2crbh8sUD9eIgB9AD2Nnj6OIVa1edD1215xOJY3j1eOLQ5W6lzo/vCa
hePFz3gVaFsUSu2J8SwB+rd6V4Q1Ybkgaxz+CNl+1jfqCdlahAfzD9sQFNutpfK3
Ioz5WcS3FROTHsW4etFN/p5zlxjE2+O0aq5570WNtVd0CGNK9c0r9PHEIiTjONij
Ng7/aRuliOAGxUuy9KJdnMRjUm0zIDu0WV413FmqkUa1vaNrWeI7kQj1xJcoS94r
fKrLYmNOqJjV8CR0M1uhhaguCVJjdMSL6kDYRMuibD9V3ZaIDdK44LDo+/MyPRo0
XQwzLzFL4XhBwfi8y8CYeiN7lgS3GZivTQe6QmFahdVcJnmO4GCmMnPw8Fi28Rr2
d8mE8C5NvKJKlSiPtB19WQMMi6XHHlVYf5g++LrRWYv6ylxxOdwev1wCIuGzO2Fa
p9e7CVzqf2ffZxmaFBSD/w9Igp+zwNtImOD5otABhOochCS3I2mbIoNP93cfs0Tk
Z5G+oei0AOFH2mhfWR2uUXyxMgunYcPBS7yY2tyZwT0Z7n7EbCaiu+MIXEBhfu+2
9pVJ3eHgihUmbc0gVL5eerxOAhSVpF0IFRK0pCcXo8jQ1JhUMVenwCza9mQ0xCaH
f+eDCjAZYEuu6vU3uNsGkw5gFtHjYznKs2JA/tDRucrYMz4B8OjhTj2WHS8EWyHZ
mx7Hq3j1aOAQXN+YS4wCzm6YCkr7ZyyUG01bvEq3x1c2eiX5l/wD4/8Xudph1XYZ
m1t6OlTUJWdlFyodg8wETCMHwKJPM06XCZLcXDPJmTrKTf0r/RzeZSPbK4Dfqi4D
8ie3Xuko66hdNA9xoIK/BIg6PUyCTuqy5TRKfYjDfxccalmWPuexmMJwTdwS93x0
KXgZfN7MgGDA/MVq9p81k4jK4F6T3HcPSq7rs70UkmR5JzJ2JYaabcKTdjESDcl3
XkUAU/j4oC3PBbz6vTaxObInhMtyqU+MT0rPNYzkr21AGsRAoovcpJjLnhFMgcnc
3taDSwMVp187gbR3Href2oR+MjISpZxdPkgo7FyCkrPwBLRUxatLnX0IUV4QH/RV
lre9NrOlGZbd9YzqpAmWwt2Ll4rm+UWkhDyvxd9gXSz/8/9aWJ3e6QhZkmYaPEIo
DdrGgG1z5sPX23CEMUibgG4I1EtM1QlqHDEblanOHh0IVXjWQmlqg5OGA+gSOHbR
oqLGUuVRct8eTmZbD1VEdC0K6zoJxddW53CeVCJ/fujUJByej1uZEUTtDmFA2KQJ
9PFXori+fEWvxKhDAJ9vtLq4pW9k2IF9RhcL/zlGq6AZ7qOnGDJh28jIb142Bf5f
QVyTgEKnH0MnxlAvjg9EQZg2FIzZNR8IMyOilxfWJG97yswxY1QnCYsHyaWt1t/x
HatXuhMZL3gbIGYcqjPMmA6rePGlApNYRPb14UEXKgKYbjNnE99iETnbrMlRn/3Z
EIK51q/lmTVK9vZP8ylnsVJViNi4RdcvWUz9C9KmMWukcxciSPJvomBZI1vpUeIy
Em32IE1q+NDeUiOr/xga6+5eu2UuQOsUQOcs4WEAbRa/Gd/cMAuo97mYZaYr55tl
TtjIHR0Y31O/NcqLIOH26VRHMNvmseWc9WCWQYkaYXUm0XUC+m5iaBWx8nkM7tdG
TBzqma98YW8/cFjokOkmLUmGuX7FNazjbf9XaTFx+tRaYTJRHrE7zMnenu9wnIEN
FNtK4AMCwlNuDuB8Vldpk3BB5LBMjiQrMZ07/bNUZyp3ApKcOIUSfUdCSroaQOy4
Zl+4y4WkxKEdCwRvwjfSmPyFVxgYBKa5eCwKRSBlmTTLYnSNaccKk+YFzEdUSHqJ
EQARFSsoMYRAwIQvwLpXyBGhVlMyxjUByP7Bmvr/XgZvIvuR/ZxqUNNQXxpLSq+u
0g1ICr2JBKAD/5FmhDckGPsarxWL3PgpnnbNxOoJPYUZxg6+DvXcLnBsLdSNC3o2
FJy5yQ3e/KoSVzyDl54VgRtj3rX3xmR2u1NMnWYCKRlU6ImOhMqO4HxfxYTTzETS
OzdbLVjYttvZ2+q9p62p3oZmdeqvHdo2iYVsY2/l/HgB2L4J4ImYCc3HwUb+4Wfc
D1Yi2726hbAAyFUqyzRCF5OmCy16yFgjn8/z4EHt/CsWngiuNaPrndU+qSfpF2zO
Y0mBbMR/Qcfg8AtMnxsC3d6iUSytkWEWUyM/btVpZu0ohVC0Kie6XPEWb1d8ugRW
jgVgWwVmh3eC8ooRETduWW4GuHDlcTjq4bIc40181y9osAa4tYn/Zsn7pLy5Dccy
fkQ0o/TjMgK9xs+RhDADq85q4ZhK6vbBmHvJ2I16/vVxERn/9ueIQc7uaWZPV4+/
ijQW6PeeeoEqlj7splDF0JMfkl67JdiVADEjsb5K2280vRPmkA8qC1eq40eIjSXg
yllSGvHfa7vSpxQsrOZRewYWMInS7jhc44sD9GxAGwxYhdZGfE7fxNDg4OgQ/d+t
LHY92diSmF3Yi56vgrFMPNdFpu1VUDMbpIiDacGBWDE1yOTUgJbGHWSP1NcBkuSE
3p9aqaIWKEju7iuuRMamFWw5ZWhvfMvTkEC1uje5aIbTpBBLsfk3JPaNc8h07Xa3
/C7gq4ui5q073GTbGwR3EyAawpf/vp8DWsXOfyoSPH8qlfCKau0B5WlHrSZivfHQ
IU5EsZDSSTmBncD3Xcl+wcqdryQR1+p1MVdjL/klBzAfqIuwxnzkUBJUlRprxNme
Mxwyuj3ljwR3ui8gSt5molQPwYsWtGznCbJROijelBNy7IzQGsHVQ+s+i1CUslgr
aGthU2gpnxuMQRzACGtr0bKxAUuvq5zRWXA4Ehv24Qfb0OfblqyikYMnwx3jtnpN
9uMvAAlTIpVbL2z/YccVTSYRyJSE40Tq6ZOWra67wL9jPMYOrTkUNMHKN8E4fsHs
SDU1IrwID1ccylD9PUvo0anDvf2K16ik4/S3A13HRclbgh4+EvS4wsp7ukvqIM3Y
l/nbZF7nTH1vWxD8PfcxmlEzHEIGF23gMlQbc8Ba+Q0gqE05S2uZbf8HZd53mZzK
GXiPqun4TdJlDFsVh3XWCWjD5sbaSVrXArdeddVAc6vTsoT/fyW5cUtwr0UwHbgT
kqZ7aQ66d3gryHxPuoZTNWmzM6uP9pdZMJqNtSJJHKR5vTslrowL2KB0mJGNbVo+
pfCPZODdOGBSzSzj1LupcQPVfS8WS7QVx1tGxTiN661KzDzH0GIJ8FI8DtRkrTOn
WlmV5J90DjZpnFfq76CSma0uf41OuXy5WOP8YO8/BBZSsn4lkE8quV049+1FEhNi
owhopmSJm0s7A12O+cdZP7ZShETMl2sWrb1aVGlt+5f/NfvmIXYvUqJP48JVEoTx
CBIQFm/H/mgGN+T7GtglP/7MCZSjvAPlTd3Z6D3UDfLiQOL50ay5mSzqkK/TJ1o7
AlP28WZSoOm+z+a0XUgPCe189lEwzp5quqzzDipmpuxrAPZiaqn8LmeH275oEgrY
f/qbPsLO5V4cKCUTnkjb1l6+F43XQfztiIxWpainRNpCqkEW5yrIOvTK3MbtL1T3
/+Q79thUylhJUWqMFDIwtFhuSt6PDYDQ4NXgLigg67TCVqOh0E0uXwME68GiEUCh
6wYIyjWDh016UYzYivunadc+BWSTLEu0MYnxM0gAdapYWa3kp22hKrIf2I6OzXT2
DpV6NTlPZjer/t5OrRMr4Kw0wtkahl/A2kx/k2VQWON5XxlFvJbXmTY4+uzqe9pa
+GTTJ5eh3Y2gHRdQ6cG4p2Piqyfyq5ghNNf+3pdfShAF8884PBz++FnBhPCclBPA
90WpuCP0nENAIJNORGWWoQhgLRXN8mq5PFI0hMQY8YWWnSo5irN4/Quoy46fLQe8
OeI7WTh8VdlA+Id4ZSRFBB02GpuCCjoljV2QltT9dlI/lLsYYFU92FQQ4P3YFnr9
UxZuRxBeqOoRQVBWH2pnkExnQn7aumiUU9SWTqIA8MJNDLHn7H8Rt1TdzfHBIOm6
2zBREdLuDzKcEeWcMGXJWKwi9MCeI8PuNiCLPahPw7TCKKcCrEDx5iGt/2ESbBwR
gSRLIz/VLm2CYNKBiUDDwIknT9JltxUJ47ONhFR/Soid3MIce3sy6fJ2Jkpy00E+
zjyEuIVXERdY4WyUoeVX8RvMci6zRMhpj3jfNxsl1KlxWsAL75Vy5GktCqATLHAZ
8B5CoUDP42aCC//Ux2hrRW5X5ntNnQzC3AofWX2MRcN+qgILL7xDTktkjvplG57u
9dphLrxfiIzNQuUZL3i8/uWWEugflGU855oNj8LlWIgNm5gB/A50miwobN4WQeqv
zU5Ypl522rPTKp7tUC33fNRIBbMzG+cn/g8oPIZ6pwLtDeA/nTF5805PypOUwgCQ
uFLLAC+1EjcgeQXscdNOQb1z1xnF8Vno3UNaUHMighcQ7AIncIGMs/5dpNOzpIDr
1Amia9bk6zrY2Sl78WMPr8iklxqD7s4uLTk9iXgk1YOdtHgMDkA/BCJdzA3N/EZ8
SFuFp/BJ2wM2fPnNtz4eXf3NoabypeUy3An2VRxZoy/dEB3ARk2JC26UO6YGPKjb
7zKZGYLZtdh55OGISDu/EN1G16DF9KwOs/RnRNgIZ6Q4AlkCG73dJvIYOJaDcE23
oL4jGff+nP+WUg+UsUhTv0OhHUOwEXrH8H1F8wbgbAwGX+yBWn/3LDWPQM47q85b
1uzc+wmgvCNGIso/UpUclmqgiesSPQFgU7IrczB/Hs3IqWraNWB9WMmz++7+ckZt
3Rz132yqPw3yu/NrVQwxX7oTFXkU02N5eivxI/Ao42P2D+YeM6lOODU3JPEnFR96
XFfncpEtzOTDjSfohczfS70UJdHwqCykYZbo0KodwAvRXqZEsXJlEyDHMtZoIeCl
U47WZp0MjxVx+PaYwIPb1rhB+uDnnGBRlNBl2UDOoaIlrDp5H9aeBKKc2ioGJ3fv
wS4ivSXeOw6/EyUNXnj65wLp0n7btGbH1YNB5YxfRb/cmz3ync/5CLpvtMIsB9AY
cKu8mReP5/ZbaDpv1ETg1ajSpqPAbiRu1FyYv3mLFlRsaZAS0BWcLOQq7P8TsV2O
zOYs0hFLc2iiQoGeYN60Ro8uRQx5bJKTdoGcMCOp2hXpN1EY4qHsPdJX4jTbMGfL
V+PkZBM+Zsf4DRc3D7RZMG9t6bbnylE24IZB+QABYqQoBFaAo3ith+naLIpOtADm
/ujpbY4tnrJaGC0EuKK0Q6OVG0Yxxyl9y8nnrEOnWUmXhD9vYvFarMaVi74I1UTo
NLOf/dwehb4WvYyuWl89sTRC4v5nny12B6I94ScCU2u7uDu5SETC3r6czgqFDp7+
I1xSMmyiZ+vOkr671nv8527vmWuHaeQh0B7Z4734/Hg10+kry7zZRiwYrGrdSqUZ
LG+0mjXU9Ksam7qcXbYna9EkIf5U725WCH+aiwfKnfrfLJCjtYDMMLdV8EmI/6Up
KJy/kTNM8aHIY9jxNPYVJ3ALPzLyv1wHNoO2S5VBEdfm4TMgNx0RI+uL2JZl8GV8
qBMkE/o7v5Q0y5qhJeJ6DGXFbYmYJjowA1OVPX0LeYJoIu3eXXZUM1gDVQtwhNRg
KztJTGu+LZ/XWP+G21qcb2svqQ7t+H5qihQeDQgwJvbRv5nBWSRvPgPtAwQGWF+A
CvQpRXw59Tre5J+LNbdDmDMs6BSiox13D1La+jzqgDy47XEJ/JeUWuSxkLXiQjUj
0dKGwxARrx7zgH8AMCKjX6Ui4aGCS0J9mZjKa4X6hcpHujpSyIrlD3FW1mYPBCiY
DdXV0sTyEQteiYg4x57c6KAuyGwhddxj8QfER1JQ387xHfQDnKYUdebS7pNASEes
6SrrHMqQ5JxKi4IL6SgizErxCk8/dN27DbmYaw21wQOo595HdsrWPV5MIwVNDFBa
iWJg0VL37msGCYSraEjBGTLEerZjwgit/XKumwBP9EFK5XSvFhSzxwdPiTj94Tr0
yPSagVbdEcvmVGSA1hkxyCl8bLtx1dWGins0Fqoc3mtov9Kg4NFhjo3m14hYxRfT
RYDqEwACnSR0PjFfvDPr8N0a7/rzF724OQoqkUZv+OLsC/kbxlFR7pgk5Zhr0yK5
DJ/7coz0nlRPSR6A28Vtq53qNeZU2Dp3vhp2Ex79p923+W5fytfm0d781NPKyGcR
1Vjt2+Jv2pIVcnRWxVZljvoIXQsOxv5hq+FA07+Y8jQry4hnNYB6Io0/k0MWOB0E
4VAJ5tye1WgFQ2/c3HU9L3cNAHhY95fgtpM+KfjPX5vCu5jvdIrBQ/E2gyQGEvLm
KtB4ISr6d0QpqTmp2eYrww9ZQkFkE3aWpXNDzI6OGS2t7N3Af6y5OziGiGsumYl7
Z8INIzmIyAkqRp/iFfEx32BLxG2VR3NKLj5B7RE4qSH4EBHvrtSh+QoB56u99+1H
jRtdNlsuF8QOqiVZ67flYljR6PPp9Wa91KoIB3KG9wKpixQxlfkizoCjFr8vnAMv
V2rXq59ZZqKr/yxkgwSHLxZbMWr1wAkgK3Cu9gB0vnyuLpY/2MrpyMSWKwBstBKI
hEQdThqfdpRQVIst0B4zVYUa/Kt0+J3c/cCpMMBMra8lsLuvny17a7P25f3nBqOb
4YaX5V7svzdBIGKTqJYxgG9KQl/K7y8fj8YiveRrCiyYRxmfack23UBrJpKFSVwB
unuMGPozHlDyta7syw/HPUoAbXZZRrCn8W9Oa2M0r0VmURhWK4R+ZMNQCyYjr+nF
V3ANfGBLDfe9r3P71ma7N02cz/E7cZ4dAWk2OyE/59RdnfdvPNUHW7vCvBqg8lEI
C4I6JYm0lBfO9XXzJ5QZcu3p95LekQupWKhSCNeOgq3V7OUDnq2DOfnAfwedgdh6
v3dPgebCFJnvwBqMZ9KCwMZbyG46cnraOWk8ffcXHX8q2ua2RlOOhXL3lIYm5DkG
0EI1WudasELalq/G9tJRgSx6rOcmoXvgf46sFOfRbBN8/Sc4IcKgS2rQlSqwKX1e
uQ/AoN7LtkYEKkmCFHugBwRUkzj3fpEaI64Ro44dlT6FKLPjScDxcLXXXPCX0wMc
2jDzMYo/W1ZmmaM0osj+wppfr1FtDn9qGL6kOmxD47sKK+a16ODNIZJiRULzPAnO
qAbKWMfwKKciMmqspDOjqSWP67WFNWMzNcYx5M+e6Q4U5sF6A6zOjICEJjrCLg/Y
zOOQgwT+m/SUN9GibcKPyUtMFBQcFbbzC28ZAlEA7pRGuSJliWs99hTruOvrwLNm
ll9ZtxMpkL/b1/63WG5WPlThcCp+flrNEjHgv1r+vEN04ObLrs1IVJ5xP9vUOgk1
iLP3mdckc3yrtlOvWy1zu1QWcFRilzqWGKW0H0bLbb2C/RXrXNJzWRutVYg4BGul
yikdqAIx5qPyBMTOBkDnNLEY9e8cWlFMXCHbpD92riQ6NQEcb9yALMnGvtzIhmVB
1mNsfn2drJrVEBToXidDSDJo/8bFLfpQtDxg4TNmo/ULf/CoMw9MRwc2DCyLPPRS
R1gKTmf24Jtc4rK7RT03F+vybpR+XWVYy8JyprEazlD/Yd9vBPqFeI1wWfETNsXl
iAAJgWXdkSiB5shSMwyy2lr4UovOXWJegKd1NtJPQsLeWw6XAbj+i6PvflWWlHlQ
6DdNHnuURrXIoBJ9emqbHZvvPqgqwjdCjsiFlU514Xvkq6WS7h6IQ0RdJBalLk+w
L1NespBpVk0tv9sWduAZDf96QjL1qbmfp+cxtxRGNvq78gTxxwN4BnfxKjkh04BG
qPK5Tx8cngarYbGUi9Fw1mfD/mosAg7a/i7UY/nBPUbNnJuk3sfcqwzhxAVOmR0r
b55e78j0wrxiwpHpYWgu/TijJMgvUrD3frKXCNzyChY86krDqPKbHUOdgrMHQgjI
XCkpFJGSNWXRAoRb9m7JxU9ObTXoTmY6aPymFrtEcOZww+YEoXBQxXj3sYp6vmiC
4A5shGoMAHS+NHhEVtxB1Cw/SRPilxS0Y+S4yAmL5YsGQlxk+clSdZnF4oWIEsOF
SZ/lr+WSSOmbPnBy3pM1CsdZKFfcr/1LJvv7c6WpgoV6/uvBqgyqqSAJIL5aDvYV
vHSDWCxyIgmtmTOcKlhJuDXRR/bo8wQ9sjlQFacF60bmenVXtt+AGMT1Oh7Jst4R
Y6dRk3/80+ksVv8RfLUQK7ph4QePzcG3ZOnGtXiy2EWCFSJ9++4vFN8abGUmoV3X
6eQs3f7ACUdssAVgYEvyIs5V+WqvQgVfCy35rpVuXTMURmn6Tt8kK80H9mEA3/vJ
8eHTIKW0LB32DuSmQ/sxnN5PZysNoth5nfNpEVLyF1nmMM/o1AZP6y+cYSZBpRUC
nDeUp716o3cs9Ao14+Pa87n7QhMWf9Wn9vDQZaHRFoPPoAEZPeHW2sDa79h3o+BY
NU6wLyeCL+ukC6SgXHUfPzFKClFQbXf20LldhyStzjKGAi7ZHLaZKnmVlhhsCypy
nXgL9Mb5cfFmxx4SwO0XDpDu0N3QMFWFy59I2aO3QNrXR8lWAHVde+X9MNuvwOk6
gNQeGIJZqirdgu1nT6/+FObeqdzzA5eRf0CRfMYXhZsksQLOR7IruiJJE3gDf9bQ
KH+Z2btzdIF1Kw5PzZyjt/j2ufaLf8KWuc6G5OrwiTqjJGOLn9N3ghdyNpU8Nxif
xoe9aig4bRBG1LG8nND3VCQ8IWJauHqSCGNhtMo5XisTy5XoFoL/01RAH0O+0f3+
soOJ01Hw5NqPThP1cyK68KVOVMri2bBZWfMnvBI1+YU6fjucsZGaB3fv7cT0O9Gt
2GQAmHaVpLyM9uiG3eHR5NahIdzssVPS7d/eyECeeDA+BPxxH/doHOantK2qT6XA
mimTRsskDulL4yycTpEOPRnyusBlm52Mz2JcIRcO2hZkpUXFO5DUNfySPoLGSr75
QUbLbLJBta78rX7M3fwbOih5hzemWZj7rKUWTYUih195yA2BInwt21AFh+igz0aZ
fUf98ubbMVUTPlEpVKC4cL0jtO7IOdPOx1mnB2SuCfpfmDm/+v7XNCSg8LgGASAR
1sTe9qV1QKyiXF5hE5jwhVXjow/OKeSAgos8zyuWSSaan/Hix5N7mw/N8VmdPb3V
RzibWWPGWNJnPYsdfZ2YtlBgdURVYYlvvV1CxjUL/ZDtwDVOJa+hsYB28ilna6C7
LZ4sNO2RJdswMvhg3opWMmQIvOPrtSbVImCKi1lJRwnmdrPwp5y0BCCDwfGLZpoN
+RufQB7HQGHzcordp23TRfVYJGTqNp/8EHiXMdF5pFevUKaN7MDmTr1ArE+QjpvY
OXuTIPO9oGw4R+ACLvzb2lgxFP9CtJetbTvlouPO28lcVB7ysS92FADkfKWxgF5E
1AxT0+eTmu6w5da5G3o2y3Lpnj/QK6G5XUYRNjRuS9g6LNmUalVuZmf9xdCe8ZgZ
`protect END_PROTECTED
