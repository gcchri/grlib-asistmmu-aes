`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AB19z08FYwDXbfhulm7gr4pWsCyDzYjaGXKEOCo9sdxU889No9/saV7JSl5JvNKU
vTW3PKO4wrdWLlx3vfY08k7UI4YeUvjY4k8p+4pA3Q6WNX5LX2Xf0q1El3J78267
8hksPzoq3errthpEbtS1HI6H76FH6Zp3uP12D3y2JyUv+VLgk/w3xZN/nXuoN/t8
3XAWGeripgYsKgzE1aRY6awPFICCt5LhnmxZu70/Kgcrnf8gwrQryT2WKMzRoLJn
FT+DIOPSlTomQi3Qts0baFFtPgjYPI7ARiMBNsC2jnFVP8ysdn8OKoXTYrrIqwf/
+uYIs6kX+3/wi+qdbTdFywS8tg3SKjVBJiqIojhR+1VQD683w7MQGtQdFi85kb7E
3xai/WOM7U+uS8Rg/+9tJLfQXwN0DdPBU5N9y4/f5RanEEtOgpHZrt2xiiKLxCmd
wqZAsB/WLPE7gjSyu2y5evgnkVDMhZqZJRAD2APTYLHroVTEoSXYgcGa8GESDenQ
`protect END_PROTECTED
