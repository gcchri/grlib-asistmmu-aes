`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+5edL1xM1j8nRsJlkNBRNOYrKxMRwlS7lpzNpYHuT12pdUcBjE37e3eaM+azHlY1
PQnfSeuxBQAk1c2FjnklRYyP+VWiJRvK7WMCNsuqNuNVSZSjC3P/LZJgwOnimItt
ZKuL8be+rEM9yd06lSvB+MXKoJ9KImTuvgTd+GgyUwkIjixSxy/gHEmnmWaG/8yj
osFWwit8V+SYbCgdk8OHq3KqCwFhXK+HeNFOBiinFlViADp0yRVtTtl7JyF0sfZq
5jjNEBJ+l2K5fWAzUHNrDzNZV2GwNgMGnIkdy8qixi8RYnb7C4sb3rXygwD2H5gl
Vw+/yAv6S+kJsEz9ThrwIBmC2uqfNVqRy2/HzXL3ReVkoyr9ejA0CpDXTmV9sQoI
XtG2l7/jFGQfuWe9m8UhxmN41eUAleYHeQXq10z2XfgTo5NlRaFmH1AuBy19E41s
P/voFAo96/TWPWwbIwBQcUDOrMMxfVgqxcxVQMeloNuVnGiTUzacNYmQomtEK9eC
l0GX41dPxh5kSUq3JinVR26iB1zLy7g7Y5CMzSJgNKwJRqjTOYt+sRzPmbl3zkZ6
kDeepbl+HTUaoUaGlyGRJXiCtll6DVXeSlEBINct9pwh5nJRRFT578PIp9+B34d6
XqHnsGGMmFoRJKixnZzKRg1IvW4yY9+A4Sy1j26uJ1EMwxilfZBq3W3KmI9FCgyW
2mePi5I9ECFmzu2r4eNRbFH9sRyFEKW5LiAd2c71MTQngXkVuToWpx3uckS1IWjt
jdXUKqyM5WN4Ag+arzFd1neuOg6HF3IdoEH1gK/2Icu1PmdJIOsIi6AX6BLmKCGq
YSZ0YE5Kife6NeWy/B0x/FsTNXG5O1r+d+qWj8+uh2jV6qqvqt+lpGz4oBOY7b+U
KbCat7wDYd3sFMMAx8X3MPBm7NfpBrug8nQo73ZXbSNx5gCYWzwxrS0khOX/pl0D
vjvOblUOOxe6UvsR1VHM/bgyU/fdc5q+RSlxM+/kDE9KBCPrtyRKMx9svTGjadJx
+9vVblxZUn4rEOi1/ZfkWQd8R7PfYRPghg7gcGtSsIMB4kQADfE/Y7uN/W+kd96c
SUCwvURZPg+bL7uMEDKYyDN88LRrHIokxPqgrTqKuZIBbUq3qwi4phdq001kQ58+
sGWkx9mAbCN1Ff2z8m/G3/9vkOpUBMGklAsyU3G+CWY3tOmI2LyWVcIxZuCDNlrC
uyXPQIhqHp1zP8aOHSBiiBr7OiWp8O+ur4t6zbKzug12DulRQgOVd1kdZJslg9hG
aBe1qRfIPf5weixMQzMfjnxiMgX3niVPP61fe4Wcn9+Z6dS4AQ5pzUUgJUSA6xkn
KTinnsMX6vE5rSBIQwgT5Up5G4Kb8cj13CEs/ebgqynOs813fKY4t4QC3PGMytfq
ZrKS8ZD7sp0UJ9cmaP+n0+Bfl090BatANigsyu3ZS30XkLx9oygwN2FutHXHJum4
N8q5WcSXBe3emU1U/IrZvVkonH4/IuLXxuZou5zUvSTHMsIM4l7ij0q7xUDG21uK
5liSGR8tyjHXAWbJw6oX2ZoYOhT0HTPWImbiQWYGouFw1Y59VPFK/h+Qf7+AI7tD
X4b+CInnXUmgjoXfzzbBpylSXV6mEhJOc55T77OOhmp+6Ypm4pUc3Fxp0IBFKS/v
Gd4vrS9xa356H1mtjLmDjKH5j4hDghcaSx0wvvzgDxLBMCNx+rV7rCuJP1WkXZlV
lKvezfmQa/MqXIekkE4QDsjrT39biopHoJBrF86+TkROTDBS1wUFeXk3Rni91FhH
0OwrhKFd/5g774KUlwJEZw6l5F7je4FvXNGiq7XCYIi8p11BBgJ+UvD/xKmOrijI
h5Yk5lINWWyXWP6ZvaU+03gWQlIP5jAEJvlrrD92zktAcO6G7sGpV+txVDAe8SUc
FM7lQ4cYrrluguk58tUu6wh/XPtEQVqGcDav+UfWHvgm9sppGh0NLoRC3uDWrHj/
RKleq2AophkNwfkoQhf0otpP76dMDv2VjRa6prNR8CjxgDzLdfCceOCTSkZbg9tA
BuQFm2mfx3YJYCG5oaB/ryQZi1osLwLy/LlRFkZEN5LNGZhAPWEZKfZMhKGQwJH7
5xupYwGIhphUr4iKlGcB2phfXLJ/zlzLfg1VtbEtONAid1+lgbmyTq51AJzTvcQD
tb6l8qOguoq0JninnD8zkCgOlCtOItfWBEYlIynaRhapEKKge4VIiQD2lvmRFxEU
NOMtRA4eB3EaCJURvXlbDoHatAc17+4dT6GEAq5NY5ZtNXNO0KZOnTNFQ39FnB6Y
wMaGubbiAfxhbjtEb19anDVTlGVTjO5cQyYToc+gpF0wllyRK7VeYL7AH9oZaaB7
MxvXLgOIhfnFjIF294rhHP9/jnYtPle/tEHfbgXFrlJWD/nj30mIXAZCd0Zsjj36
kQQhrjVlmDZxjwGsVkuWAtN7AjU/DS81HXJs9szOaILmCRJgHIVBI93w4+eaiHyB
aUKFwZCASBcfsFaO9Ad0awNp891v3mVHXA4e0F74MwZzpn/4YVN0YoEB861CRZLW
ALzw3Lbt1BhI0oDs8y9f/ZIWATY+eDk35m7sO2SbrcqPA2VQzQVPm/DWhr3KgwPH
KgQSJrQlihlX3pXB29DYZo6IjtHVXwPdxHUytpzXgKnpam8tgIfqDcubncv968tq
lYJJY+Bf/QJS3MhK5jnmOePxGArejBPS/UPxhsdkUy+m3y4TWWawKFWVsg52HRtx
ERvLA06UsqIC9r3CFsN+SUws9pToZUPjJyShTkSOMFW2rBk30AHW+mCA6ZTI8ixf
4E3z0MW8EBiXDm0K2hv3QQnY1+TOIRZ9TossCgFpiPFuXrpbabuUM3nI1S9K0Zwb
FAHMkZ7lkfQaev5Xz6zwycEdqN5IcHi33KYJAzt+o5Mnl6D4Htq5n/oso97pza2e
QicG9+dnjudZJVSOzO2kT0QqfAw92cS0chUOjc5vHK+VtjiE4pkvVHJ9atKwgv0L
WTmFplz+iHDx//HsYA5VtPd3ybERq8aksFDhSuW9j5dYtRZf2T/nBx+ibfDj5ZQn
CY285bKwJS8U/9r6o6IzeqHZMVL1h420bxCcvOeoXez6ZZH3BcSaO4QfZX7KpUp6
Ap4qvr6wpr5itVv3x1tUNj/Rr51H3m3m2fKMRYU7qTzpuGX8JOj8GN845xP7NFEO
ahRHWmvrk5QaYZN2B+qTtvGNlos1VcQwDbJOqT+SnZqV9eOqVfKVhL3HKYIeBVpo
EvUUUlAIUGZbauB0zTOwQHfEUmqgJ34MRXpTROykRHZ4D2dnvSCUo/mzSwhilnuA
+HgZLcrA7/3equ6uU+bapO7SaQNc3lDgnN/BvvSIAhbh1AB6kwHkAEUoxWGL270e
CSnebsGQvSYGGFYkYLIUrA==
`protect END_PROTECTED
