`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ph9/0P/f+M7kDmlhdNdDoxUAIr7jU0UwJg62mjwkAs4r3AaUn9thbz9yAIty/SfA
0rF0GRv4Q/E3kpH3nQo9jH7SWviiYx5I+t35s3wrZ21mLojg7fHKw9zseynLEhGq
irITyjrrfMWGUH0/UE/J3yGgdVsUUEqG1cluua9GfBwKPdNcK/umxOQFCyFi4WW/
f/A2m8JC2SrLWD3o4uPRen3pJh4NY/qAhMgfh1Pv/77HJfwyG9z01b+oSrYPthov
cDvyZkBcUT5+E08X7xhYWxG94Y6RJr08qUcEzvcO5vI7hmK8Yt7/h9lIT5pO5kMR
SY5qtN7EfMEi1hWqJCNdEB0fdj09sDqrurzHTK3+whAthd+tZPIMsGzi/s6y2KDs
r60XChrUJpmw21tW+PRDG0LXxwZF5nX+V6MhVDiHOXP1GoAcx4Qwrenv8Q776EUM
z8viJL/egI+ydFxPMLlYgSk59fNUHDDx47y/Ncrck60=
`protect END_PROTECTED
