library verilog;
use verilog.vl_types.all;
entity mobile_sdr is
    generic(
        tCK             : integer := 6000;
        tCK3_min        : integer := 6000;
        tCK2_min        : integer := 9600;
        tCK1_min        : integer := 0;
        tAC3            : integer := 5000;
        tAC2            : integer := 8000;
        tAC1            : integer := 0;
        tHZ3            : integer := 5000;
        tHZ2            : integer := 8000;
        tHZ1            : integer := 0;
        tOH             : integer := 2500;
        tMRD            : integer := 2;
        tRAS            : integer := 42000;
        tRC             : integer := 60000;
        tRFC            : integer := 97500;
        tRCD            : integer := 18000;
        tRP             : integer := 18000;
        tRRD            : integer := 2;
        tWRa            : integer := 7500;
        tWRm            : integer := 15000;
        tCH             : integer := 2600;
        tCL             : integer := 2600;
        tXSR            : integer := 120000;
        ADDR_BITS       : integer := 13;
        ROW_BITS        : integer := 13;
        DQ_BITS         : integer := 16;
        DM_BITS         : integer := 2;
        COL_BITS        : integer := 10;
        BA_BITS         : integer := 2;
        full_mem_bits   : vl_notype;
        part_mem_bits   : integer := 10;
        part_size       : integer := 256;
        NOP             : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi1, Hi1, Hi1);
        ACTIVATE        : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi1, Hi1);
        READ            : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi1, Hi0, Hi1);
        READ_AP         : vl_logic_vector(0 to 5) := (Hi1, Hi1, Hi0, Hi1, Hi0, Hi1);
        READ_SUSPEND    : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        READ_AP_SUSPEND : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi1);
        WRITE           : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        WRITE_AP        : vl_logic_vector(0 to 5) := (Hi1, Hi1, Hi0, Hi1, Hi0, Hi0);
        WRITE_SUSPEND   : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        WRITE_AP_SUSPEND: vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        BURST_TERMINATE : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi1, Hi1, Hi0);
        POWER_DOWN_CI   : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1);
        POWER_DOWN_NOP  : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        DEEP_POWER_DOWN : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        PRECHARGE       : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi1, Hi0);
        PRECHARGE_ALL   : vl_logic_vector(0 to 5) := (Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        AUTO_REFRESH    : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi1);
        SELF_REFRESH    : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        LOAD_MODE       : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        CKE_DISABLE     : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi1, Hi1, Hi1);
        DEBUG           : integer := 0;
        ERR_MAX_REPORTED: integer := -1;
        ERR_MAX         : integer := -1;
        MSGLENGTH       : integer := 256;
        ERR_CODES       : integer := 16;
        ERR_MISC        : integer := 1;
        ERR_CMD         : integer := 2;
        ERR_STATUS      : integer := 3;
        ERR_tMRD        : integer := 4;
        ERR_tRAS        : integer := 5;
        ERR_tRC         : integer := 6;
        ERR_tRFC        : integer := 7;
        ERR_tRCD        : integer := 8;
        ERR_tRP         : integer := 9;
        ERR_tRRD        : integer := 11;
        ERR_tWR         : integer := 12;
        ERR_tCH         : integer := 13;
        ERR_tCL         : integer := 14;
        ERR_tXSR        : integer := 15;
        ERR_tCK_MIN     : integer := 16
    );
    port(
        clk             : in     vl_logic;
        cke             : in     vl_logic;
        addr            : in     vl_logic_vector;
        ba              : in     vl_logic_vector;
        cs_n            : in     vl_logic;
        ras_n           : in     vl_logic;
        cas_n           : in     vl_logic;
        we_n            : in     vl_logic;
        dq              : inout  vl_logic_vector;
        dqm             : in     vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of tCK : constant is 1;
    attribute mti_svvh_generic_type of tCK3_min : constant is 1;
    attribute mti_svvh_generic_type of tCK2_min : constant is 1;
    attribute mti_svvh_generic_type of tCK1_min : constant is 1;
    attribute mti_svvh_generic_type of tAC3 : constant is 1;
    attribute mti_svvh_generic_type of tAC2 : constant is 1;
    attribute mti_svvh_generic_type of tAC1 : constant is 1;
    attribute mti_svvh_generic_type of tHZ3 : constant is 1;
    attribute mti_svvh_generic_type of tHZ2 : constant is 1;
    attribute mti_svvh_generic_type of tHZ1 : constant is 1;
    attribute mti_svvh_generic_type of tOH : constant is 1;
    attribute mti_svvh_generic_type of tMRD : constant is 1;
    attribute mti_svvh_generic_type of tRAS : constant is 1;
    attribute mti_svvh_generic_type of tRC : constant is 1;
    attribute mti_svvh_generic_type of tRFC : constant is 1;
    attribute mti_svvh_generic_type of tRCD : constant is 1;
    attribute mti_svvh_generic_type of tRP : constant is 1;
    attribute mti_svvh_generic_type of tRRD : constant is 1;
    attribute mti_svvh_generic_type of tWRa : constant is 1;
    attribute mti_svvh_generic_type of tWRm : constant is 1;
    attribute mti_svvh_generic_type of tCH : constant is 1;
    attribute mti_svvh_generic_type of tCL : constant is 1;
    attribute mti_svvh_generic_type of tXSR : constant is 1;
    attribute mti_svvh_generic_type of ADDR_BITS : constant is 1;
    attribute mti_svvh_generic_type of ROW_BITS : constant is 1;
    attribute mti_svvh_generic_type of DQ_BITS : constant is 1;
    attribute mti_svvh_generic_type of DM_BITS : constant is 1;
    attribute mti_svvh_generic_type of COL_BITS : constant is 1;
    attribute mti_svvh_generic_type of BA_BITS : constant is 1;
    attribute mti_svvh_generic_type of full_mem_bits : constant is 3;
    attribute mti_svvh_generic_type of part_mem_bits : constant is 1;
    attribute mti_svvh_generic_type of part_size : constant is 1;
    attribute mti_svvh_generic_type of NOP : constant is 1;
    attribute mti_svvh_generic_type of ACTIVATE : constant is 1;
    attribute mti_svvh_generic_type of READ : constant is 1;
    attribute mti_svvh_generic_type of READ_AP : constant is 1;
    attribute mti_svvh_generic_type of READ_SUSPEND : constant is 1;
    attribute mti_svvh_generic_type of READ_AP_SUSPEND : constant is 1;
    attribute mti_svvh_generic_type of WRITE : constant is 1;
    attribute mti_svvh_generic_type of WRITE_AP : constant is 1;
    attribute mti_svvh_generic_type of WRITE_SUSPEND : constant is 1;
    attribute mti_svvh_generic_type of WRITE_AP_SUSPEND : constant is 1;
    attribute mti_svvh_generic_type of BURST_TERMINATE : constant is 1;
    attribute mti_svvh_generic_type of POWER_DOWN_CI : constant is 1;
    attribute mti_svvh_generic_type of POWER_DOWN_NOP : constant is 1;
    attribute mti_svvh_generic_type of DEEP_POWER_DOWN : constant is 1;
    attribute mti_svvh_generic_type of PRECHARGE : constant is 1;
    attribute mti_svvh_generic_type of PRECHARGE_ALL : constant is 1;
    attribute mti_svvh_generic_type of AUTO_REFRESH : constant is 1;
    attribute mti_svvh_generic_type of SELF_REFRESH : constant is 1;
    attribute mti_svvh_generic_type of LOAD_MODE : constant is 1;
    attribute mti_svvh_generic_type of CKE_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of DEBUG : constant is 1;
    attribute mti_svvh_generic_type of ERR_MAX_REPORTED : constant is 1;
    attribute mti_svvh_generic_type of ERR_MAX : constant is 1;
    attribute mti_svvh_generic_type of MSGLENGTH : constant is 1;
    attribute mti_svvh_generic_type of ERR_CODES : constant is 1;
    attribute mti_svvh_generic_type of ERR_MISC : constant is 1;
    attribute mti_svvh_generic_type of ERR_CMD : constant is 1;
    attribute mti_svvh_generic_type of ERR_STATUS : constant is 1;
    attribute mti_svvh_generic_type of ERR_tMRD : constant is 1;
    attribute mti_svvh_generic_type of ERR_tRAS : constant is 1;
    attribute mti_svvh_generic_type of ERR_tRC : constant is 1;
    attribute mti_svvh_generic_type of ERR_tRFC : constant is 1;
    attribute mti_svvh_generic_type of ERR_tRCD : constant is 1;
    attribute mti_svvh_generic_type of ERR_tRP : constant is 1;
    attribute mti_svvh_generic_type of ERR_tRRD : constant is 1;
    attribute mti_svvh_generic_type of ERR_tWR : constant is 1;
    attribute mti_svvh_generic_type of ERR_tCH : constant is 1;
    attribute mti_svvh_generic_type of ERR_tCL : constant is 1;
    attribute mti_svvh_generic_type of ERR_tXSR : constant is 1;
    attribute mti_svvh_generic_type of ERR_tCK_MIN : constant is 1;
end mobile_sdr;
