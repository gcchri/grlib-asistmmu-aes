`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GssXd8WbrAMa5A7kEcGgtF+55Aw2Y8nm3WS/7Di9CrIaAQLbBFsKrAIU4Xdc6PZV
zJj27UC5TkEPEofPlG0bqZfDADBXcBXxxO89oYlKGzhvbeZVZrwM08jRfji8Dpmm
yqX+LWzE+2LGow4FHDCFSb7f+PU7OaXYd5pNryZTfM/K7tQqF+HCaObeBVDIoKso
LrRbWxYj6lKBZqTRQkr4vR47tzNO8la2hbfS0Y5ZsncXsDQnI6Hc5TAe7FYd4D75
pJ+3Ig8ENqOxGpfmGhifmL3hlmvqs4ul7kVscMyquxRcuk+rHFWRAPJONT8WXCF3
IPb2Y8rtiqQVFF0QHuDSM5i9RxylZudKe0BJPAvy6yQe7bfV97RZHcnKgpNpQp48
HslctTqZ9UNaQ8ERPYTDYdQNkdIzhPATCV0FY4cVSG7N4u1G3KoWP5HUSzOU5PRS
koJu6HHGK2ggyMrQfES0Y5yXfFl+irptdmFyAbbka7UJDhVxFnu/1nt0sEaSAffy
Udlz7sqjkCYmUscTWhXoUWP2lHantfEbPk1eZaHswzBiJbWr9HaDLifxL/OFSSB/
nG0QbyQjqdCkjCjYqBl+g9d+JwPt2UFBsBPDSZ9WMJBLirBWDfpPJzr1SGr3to6b
5FjqfLqK36AdrT5sdioZj8Y38uju0nsZ6lwPxz4E8+hDAeWV6ckasS1bKuOqAP6w
pNdr5pH07e7m1Zn4ChOUMoXZ0IbEX0uYnZyATtIuyyXpYnTfkViDeJlO3e4/ycQb
CKcvs/xJth9QYyo/5TVGRqqlXK4xwFkxQhriTFSkiN4Wb5ZFitfMm4Tc5qto9+IT
nisvJnw/CK4vxBK+kcfsP+lqmVYP6EqfqgZVAQta2vZUmt2A0q0pGlPYnjs1wFfu
G40ffuNSRT8HPA6gEtq7m2DihLZMHH/gBO80ekhKRCKTDIu2zYo0OcQwguqZuVQ1
yvaYGwSqApwGqHbRsZvF5q5/NeFFx30y5n/loKuWVZESJ/zu+glVsMD84r2cIccK
`protect END_PROTECTED
