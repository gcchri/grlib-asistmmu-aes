`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S2/XvEivvK9mmAeO4M+DvBKeazaZG914yz10YlVZkkl3s3TpHOdEaJa8oA06Yj7O
oW72uw5Kmh+o7SjTOD8VGWNrBOtHKWVtkSZHXBJ2sqbXpvYMl+SmzQt3svlS6LbE
DybLHCByo1Lb/J5VA0yEqlVox2qXzOyuyytqPciyIxztQmfexOfzttCSqJqzVskX
NVfCAv+5XvYElpGtlbYX/NDvgugEZD0MdBPoEGu14Lygy3SvIELWznoCUQmiDiMS
JVXEM4iASl4TtIirikWxkl0eXMLIk7zkW/0I6Oq9EbWKpg9irVmL/hAFngtFruU0
Y/OTA0wQj/1t1fb0+LxdAQIrTwegHZqj5Ca1cnfeSzljloGVVTBw+nTphk3JNfcR
u1HQ1ofxLVlP/zwhd9PwNsutqEZL8lYiR53wnU2rnOEgoIo1n8okfjuOAvmTSg10
emtblEhwY5cS9QbyXutq10ZML3od+VskkY34LOdto8slGhGNynO4gkxtKyam4Vj3
6kyACLRhoU8DIhaWr3Mu/fOqZlTk/1PLhZZpNBz8TzMq8Fj02VQEUMIVPTjv6pWw
YWymTdViaiC65BHJg8oEmU0pZCWQcLv16Vci+anf+r/3FmDV2iLbO5vwKlXjzWua
i9cVmkpFrjhbL/YDZDqYKZwZHlldNOwgiRj4t079bcaUpjP49uheKMyvS5DFJjhE
iGokZ/6qBFOJzyR+VIQpWQdpd0jLByz1LwMppBHC8hAIS8mIgFnxr3EpEwZdWNqo
+tGwsOIItCfocIoM9qCavuaKXzoVqE580haoqfOZeNIRjMjL7yGDRS+HgKwf8i0D
qIZlNWN00Td9G5JX4qSlH8jw5qGh00yf7NIfcN++2IN358AIaWVOPrzdePmaqD2y
s26zKgmB2atBKzGB6Rz2KbyH/9okq8CDwtMdXc+x5W/7bOOBzCeo2lFBBnYhiSs4
xNqD+WaqK04KU38opaiMenujQJCbmFtIpkAhRGZlCPXu+kAIbTMckMw3t9a+MAya
2l7/iYK8IG69uwtMXg18Z/xbUnvZzBFjaAHObV7QKfPhEBiW7UVCEuIrNSru2lC+
NyPJVcRprN6dX56Imk8i3wIdALBF1Xj2JG2bU20d+wISUK4qKpVQuQh1yycncQxI
Q7e56bIVT8dEbxLNgzNuRIZm6y0E++0UMlsXbUdocLtd0GU7ou52xtpEWHbZCX3D
Et4IDbbuyfDjEsjYKKqJX3t0+TXNVBZnRhP2MmY3eaN9Ph25QbMIP/fZ7SwJFpf8
/X//k9Ovq2kR8yG7t4U0BzExLxSRc05SS3JQcrRvURzDH0BMI1ZdKxWCBo3l4Uef
iRixO+cB+hIZLDlR6dEaMK2Zdr/+xaprG7prWRFO3HS2p7V+LHQdWfexXAGQPtbW
hQCki6G2zW5OLJCkOI41UFrFC7LA2A438HkyWf6sH/D+M92YxK2JRaB8Vd+LJ9uC
FsH8WDJXNoeD1SfC8vQppEWaaBlgVca7AVL9S0NmMgzLuOtK+JGXv9X9W0JYZfPM
jOs74h0lO41XjACBwl3IpYJcblOQ1IeR5ufgalYNF2oVS2gNxF8EAV6r0mpj1OfM
GWn1A0uHKTLfJ2yFAFwOZhQTPrmryDdidQLCoFLDeN1i0mEEjuj/oNAw6bC1pPyW
KgSB7CAxJhWCkrC+oBRAVyN0tUv4CnmI3uzfmc3EvYXFFxkv76IfARPTmuM8mCBc
ijayGb4Ew8LCu8y5rVkvZePzAdbujyLOzTIIqdf0D9ZOPjI1uP9zKXpPkVaG61gT
TMoef7jy1E405z//XspRcxyGl4xWMDe75AL5a17XK+f19hYToA3xZhXDIfI+LOvT
NlpUkdtA4PBEq3+3YXrUf3dwvGVhVR4XSbLyEHu5G2oeQ2CSJ2ovZvbKxx7QTVMx
9+wSfXYkQXU2CDP/me7xyxuFhYM2No6V1meK9cJe5Qal/i1mcssDhd+y2gdleAn6
y4XM8Gg4lZ4p/gvkKv1KvJb8/3XVyIFtvXPVILbrpO11Z1RAVkOE88Gx/1J19aFP
14PwZjvQnimXCq4xPhqDoq98lZJsCRmHhYfWHbuX8lsYFpss4uYv39Nz3Pi4En7N
v06QNoDny59D0oJfzOXGth5vVaZW2V07DPCplEfTwOh5TdR4E3hkz6gH3clt3X1d
EUKSnTWlLuqqYWkeII5rFVUM7yLDtuWGG+LyMKOgqon3hj3UTL/F4TIlJjxoBatf
JAzNe8xeveYt0tgzqA1y7R2KrUBIw/V96n8itXAQeN8ZwusVCM2fuPmids43yPRZ
Jhr4IeAtHd1zi+Jjhcdas1/fZxp4hxVEFX0T3Vgn0A2u/GUzylKwYc896Y2fBvy9
c4D44nhY8BVBKW8uIJ3+DJhJ4gQZWuXOsWnwOUPlkj9z5NT2YzpKbN/UTKsdsoF8
KHP4flkwREvT1yJH9lEXwTI7DOptjzTlgy8QUl1ulrw8GCEPg6DywB30yxA3HXv/
gHWMM3M6zrzCMmRTCJ1uqxvnaKElkxss7Hw/dVpJSsAYpJPtIzovXFf5wtH0rPR+
wQMMdgfp3HXz2LJX9ij7PjakPmK+AMC9ozmcX5r4PxlQ7a45G3s/EkQIe4EM4d9W
pLvfnSkmqn7J5wVIHamDIgU8iZLZJqfaboQT4dj55rloNi4GIWZe4Eiz6McTdUxA
7Hl8xxi467iq9jLAL2hK11dRTooOzxFf9vbFJKlw1tT8AhWZMBJuJ2xVboZF75jw
jX7jw+QbdcStyuyoBc32fMjFQqkghG5KEKAGO2GXbuaKj0+9d7j4yu4sqyF2mIMQ
m7rd/8TpY7njVaDaf+el62giFJhb+zETEl+aVizcJdeLNaiov6cOjJ8QicvtLKWp
4GGQhWcsFdtw7BuTF7jsRFPYf9l/9/0QEC4nXuhU40oJK0DR8xLEwWbOxPJWLjUx
+91uvecCX4lNsxu7UDJI8njJRS2JAt6+qlzv2zauGSUtu2e0it3tlzySYD9ni4Qx
exSJUwnN1mkQl4zlgMui1Mbmg6ME1X8oUS6R4k8H/Sizap8wqYKFr2FRgiJLA8zA
dwTuoTHle6sQfOnCHYIuc+9J/YgybYH0CKPcXogw8wYsxykQYttx4ybv7hUa8zZZ
Gd/grWClCq56sS7QoIV52ahRJP011EOCn8X0qqFKfkd7CIBaeaWrW5iZ8chivxdM
PmH+xY4fBZjSpeycnR4Y2GvwQ/G5b6h6DzQiMrT4tL0UU2/rI5rV37VtuRE4XEgA
//NEHkP0chW/bUh8YSbOxCpLiZXWf0/GMJZt1B2W3tWoXbMJDQ4zl/eQES+L2Bbe
kwcmYg41GlHK+Wuqq3cz1pienx52WGyxwcpokxDLxsClAv5TJ58ql2AhEYQnEN1g
2dtX6buOb79G7h8q45DP314maKzHdTXEeJ8Pr42NGyluXj0eaaT+e7F+N7wzktOc
8ZzgRaeqputqG/HFO2fsYrim7Z+N22MJpVnBpFYLD/0rtligtKVreGymlkTw7Ix9
BupNSTDKyGDk8jL9RRcrnzdqpUeK+2NtrrE0Fpwgv6LEN00EBzLHvi8hig+itSJa
ZamL/7ZVLaH5DYw9n3ny38aBZkTko6dsKnyA7/YI6s9p3pjG/n/Z4bl/OcF3Asqd
QBGZQb0McEZJO9wqgIt6HxW3mHPF/jQox306gBKadReBfZ+ECjwEMCzFzKJsOSKq
peHhsHPhiT7Pa33vOZhtvsNcZZj14MF0fWcpr7aNWcyig0xpmnZVBZKGiCThzcZ3
nKPHQpzEtKSmCQnZG0Ypsw/AymraxgEIv1VWtGWqaibwWGSYglcHrrKB+SGOtVWe
+M80v+Wqzi9vHovfl6Ri40XZAHB/kNuokof3QmN2R9zuimpQlc/aV52B3vRunHoN
CKA6SJ5K5q+iAxYHVDmpJEDdn7xTa7UwuGWjezW+RTeW7r569oZTZE83QDe6XpYj
mTXWPp/3sVtFJJD517F1liAnQalYexc+BxLBuB01x516e2PqRmrC2+ZWP0oYOxYL
bQ6gSQwvxbBMYh5Zaeca8qpkG/A1a8GSDb17n5JQ/RYbpKFvYz6YOQrCq4WNX4C3
yr4KrKjkhn7nqCGp0VueV+aF5uYkdjTWd5RwSBxtC4UNzS2PtIQcBM/uQelnDlZ6
FezPTEwtAtZ4o2OkBDPAhwZlNGCnMWvxTZPeseXcWMm3ie75BvcNQArdUwIC18l0
hTeZ9sNVCRzMrl2X9LHiiJaGe6DEuFGO2FJPNw1V0BJuVmjr8R7nITI52zl5kdBO
zofzTDTjHMCEWzmMiOfmjhN7T9t4diZ4eKveuvRoG0kbr2Mb/PkYczKNHiJvCD0q
T26fbPPFoK5HSXBiSmcC+Mp0DTh+qNintmcltFYYzUWPSEZv5iQZsHIpBwYIqmYY
AbDVnRI8DW7I18NuLg/+EmwcnEP3eRBF+pzYICpfAWJHvm9Jd5jkmVSDBn841Ksq
QoUKnF2P1GXWk4A/artOXMq1McB7HgMMj/QdCHkobChReh2U6+UTw1/Hy+5cPPzh
9RUIDqvfLrZNAQnbKfGOmZB6pIm4YboKYuaAD/0lfk5iE3NYKAwA27MMSCPcxPoD
Rzs2o5+i01/xF9g42b+jF8jMpJkp/DMUxSDGRXWvNFCZwMTV4eAgrNdPo4nvDwLL
sDpOlqIPj9ByBn6t2Yl/2Edrogr//c2iytxmnG/PfAHQNuAJU7Srw+pOHr/cP1qV
0Mkw43ZiQCiCXXHAVUuQau3n9dqqul8MG3b4Hk7PwSGfYu32NgEeHbNORRFaBzSr
swtOyIJdsGctPkcZ7Rm8ymdn0bK6dLJV+AB++ysfElySCVn3YaN0JbzaggRdmbUw
R3W5W+DnryW/xFhx4Gm0wyeuzi9YgkaZj+cEJcxLEtJW4PfWmOWbaC3sYi6BDOs3
6S/42H1Ufnd6Km2gsQ4/1gUWitFAdqglPDI7xyBVItaGra8JBwXZjiG0bMJCEt5C
eDAqisAmOwJlP+vUHq2sj1T+d5qlvWvQJUwPGCRyzeVKJoJos478j3QR/5zxRqam
lxX3zCTkZuLNLK2f9YtOLuDqYcp16rTlUbqqDNc6SzDgbynNzJ1oYfSmE313uArj
gpKH/2TizLobYcItlnS8byvxFe+unR6BbkipkHr5lsIsL9TFSBlT0mX03e1Tsd3g
dxVLRZ23chG5Byh9kfgoH42/eaja5ceaCfozNEpXlMF3fyn0leQ+zODVGZ1BaCmL
Jxm36Gmi97RBG9YLNiy9MAYGTE2xUzHFfGA2bCgCOsBk5Nb/qoZBv57GYuNxso7C
`protect END_PROTECTED
