`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Apqr2v3dgPpMwz/dnpMsvQOhSBCsh746J56HVlaBtf273aVM1ZXdJNsNSWKPP7eU
BWSBn+DahbmsWUXm2sHLwoTcwW+MJCfaOHoNFL/DtA1O/nnnqVDOXtfQ1sBhGnpE
m/OH2z+niHUuf72LS8Pog7aPd1qrVB1clNAxVwlQwSETN5HPUQyCHJQJN4vq4P2T
dy/QEuEa17KPiL0EIOGXIwFQVu2j+WGIM7BvqMepwl9W5gU4f9wQrWY14naPqcoH
wcXUYUhbaywmVBViiMdIX54orf4nL238vRbgRhW6lVuFVOhIE1FqarRpVlmzoyeY
3LbNLk6TjAZvXI09KwiIwutYI6eUjl6flYArkXh2zbTJtJw4DBY1wmDMOuAEJL5u
ZLeUKcmdi9uRLUAYJx5VVJBfSj2MD+gTgkBaVHbIdO+sjdMnuMFzuElVD/HzCvxZ
LnBZuqHdP3BbgyyB2YQPkoAEIxw5b4bEo/sIcJmbANxMc19T/kRXc1I260jv/4KB
`protect END_PROTECTED
