`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E1yutOcFHXrw3C3b59obiQNl61axsFs4UqmpDeJxQl2o2sFgGN5JE5TpN+sQgKCh
Kl/jU1gIYryIo/a9mF5khrp4VpzvLz5oKOZWIRfDQ2ZZLAMOg9tVIdLOP2pGNG2T
V3w0c3BYdm3YocLiroxYx9ALlFBflYSc/brCqs4bkkaf88iNYCpDRLBbOrATVKm6
cFpkuuiall2Ym46gtkHVjY3gCQS/DJzI61PyyCy4G6qxLwTMjNNL/XTRDP3A3Jp+
z7a0KQ4OvqDI3BLDOJOYpJfPgSAU6tp79lAo4nTfjOXjcWaB4KLu6WmmeQUv+DTB
kbXeJjS0pGMd+QG1/YIsMo894G5SrUZMPB4J9PWy8qMu9k5KDIm38EjTNAe/JnIo
zm6Ls9VII0KvvlMNLQynVziO8YgyupTsSuQbNJL3DFRaLIqlTnppSq63vY+BlkJC
cTsSbWqkMFe9RM2VmvdawQ8vdAyQZABUh3IJxB0ako5glFqdTr6fs0EPMJCt6liJ
i0jFbZrJECI1AHu77nui+JgEi7dYGnkUSPgARl5lmVlu+JMT6t8O41KnrmpzGUWs
fGcVt+P+ECZmL61dxVs4cjDjI+z3eBBt47mXp53kRCAdhmtwHuh4ILYfqWU/+hVN
/SRvNaBnVPENCWfSRjh5+xk/ZVVcNZKVQMHSdQWK0fEyu46ChGb6tZ4DjT2E9+pQ
s8u2Is3ti1SsGFa7qYGSi+qdwh5gb9eD/sY1vyI9NkAx9KHH2D4tMo6RiSosEgvO
s8j32JZLTu+UI/7CZEyDS+d7naFVRdaa6C7Ip8i0GmMKQ2wxAGoCYg2vvMLDmwqB
`protect END_PROTECTED
