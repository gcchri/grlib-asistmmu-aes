`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WJfjnBakXAudG4SNfQNyawdu81X93J7yqTYQWLKw43ipW1OFuoTV43jX0UUOe8Fb
I+MjOyDuG11kT+6nTkApEVSpKkBuwaW0I+OieexMGdfprDC1fM6OKI8Tw1LZOcFP
ghkNoH2w8jG4xqiea3oB5w2q7+y6zXkieIDcAFU5tMdayO5+FFu5Q1jCusYHsCV/
wQ14us7LiqS0oTP8sAdMUOdnmhmKIxyS+826QYzJ7fxqjM1/EI2/vY/hKzu3mKxl
EOqQ6nVcJMfOvwEY8vR34CA6Pvy2RaPM2g2NN6hzmFqHIwKAYJtdLjAjNId66PsK
38ItretwnRfkk+folCF825+kFGhly44s5FlouaQCK2VTSFaC7X7SwYnIRCvihJOw
x2MWH4Q0+grjj1+1baCZHEdJfYc6UcK8rnlJzHuYsgklJk5Kiku5/7FZKSLcDoV1
UtxWS/AppKclPaFTE+xznqunow5NqAipplEUuBL0Kh/C1xw1NmKejAT0mTwCBwrf
XIjAQxhWD4qE3ymh49oDweJnD5X64xaAai74PnA3aA29PVgGygbIMq6uKZeDE2Po
f7efZZijtOq+ec0R4gdpUXFSzZ0KN2Yvdi46lF4mDURU8QVdBvz4nkV9chMIYxh6
Ok5RAtwRq4YvO7nhUPLY2vPOA0cSsk7GCP5gqB9V1/RxJM0n8mMCLUjQkgxkEynP
9abV37dhrtrpiFTERS/CUZd5AThvAuqssS7Y8XYCMZERrQKhSgFPH4fx5TESf+bE
OANSNL9tjAycIXk9PXiozmQnGQ0I88O7e4w3Pkk9Bd0rG7IB0Sbg5yzB3JFERehT
Ewl9y8b41OsbGZl76TDAQxROYCJHO4E1fDiGOOeYK47UffPf7Kq6v8ID2uKwlMDv
MiId+SfRqa9RHYDMMlwO/WMuva37R9CRUkJ1kryBCJMcPQXFCMtdS5c/njv06MU/
7RYL8zfULLd9f584iVCJDe1DmJwKY/aECAgSvH4BTcQOSLDNNtCZwDYiL0W58GTW
`protect END_PROTECTED
