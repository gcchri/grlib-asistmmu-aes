`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2cFrZg6R6I7PPIwIDzdSRfC4JkmB9daul11x/EFfvhiLG/i2M8InUTLzie3pfGBE
T61syrL7hmsnlkQIZstI3runimhTAR9Lcuu68HtWlY8Rb9+Uv8bErL/elnINw71W
TLhkR9QnzSY6B1WSi72IdTNW7FBBWRv4r8GLf/KXlifqeyAaG3pcFiOIS0pQM0kI
3mS9zMv5Os6jHI5sZ1oUhFPBYWXVcwgmfVUrFtfJajTKD+wWj/FlOfB0QcZs87ra
ubZhGIRqcKmtUSQ2yuvD7HOWXCH54vEnqIuZuPTVFmLUxY4jTSdgRhEdpXgwqfno
GJJ7T6kApAAF2Q5+Ucs9OTobaEuD67J/qexfu3QvX1z3DV2fxJJjZ7T3S3kGtXRc
`protect END_PROTECTED
