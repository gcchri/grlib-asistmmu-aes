`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BcdU+7PtddIVu0/GSz1pXnqQHhAu0YwnQhS6wQu4vfcHWMabVY1eNXdXeKku5j84
926H5v1mFZlC5bSYj5m8Tendjk9BvxHGBQ6a//IuVCYvy4oSSAkXhc/vm9VNbgrc
kkb9j3CbF8J6RmeztY1+CWkS9KbaARZgQ0fFHozSES91akWEQrRN2UfWrYrWPmP5
JRWzhAd2+eO6FfU/3nGGgNE8YnUcnhSMJ83gPpXXHysU4ZZzzvzl4v3ViVtM8JTC
qcC1FOG5eKTmqQORkqOW/QFTEQqYHtidEu2Vv8KFr2RrM/VbHb5mwZQ58rmsX9gC
v3PXin/9nLIs0Rn3yfNzUoCEo5XmXDP7GzAN5V51AXQ=
`protect END_PROTECTED
