`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nY/MVck+sr+DMe6DOwGSiycyuRUX8+TRalQFI870H1LADGhf5wTvRcIPmbmjXajW
tZTQdY70KkLRt5gksH6T3PXG42kIlhhD4MXBpCPw9HkMD+AV+qPcqPnJIErmHcxq
f16YNDi9zN0l+0kxVo4zBQcOYacMDVDzmrJNmeN10aOO+wgC0OZVqC+xPhEUn0E0
Cqc0vyVlqkLy2Sz0Q0TwCB8cA6J6JGW53B/CnAXZcdVV/6Ub28HT4Hql3Wmp9grV
QT/3QY1zyiMHKvAw8KE4Dcv0P7O+Bnp+cfmm69+0uO15dLjBhz7bUJXV60INyuGv
g6A9BefGvsrDFqNql/sHhElIH4bwrpSQ0S2czok1O9i8fktGlb5zjeiEV9SWZFQa
`protect END_PROTECTED
