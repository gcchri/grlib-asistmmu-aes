`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6cBVRAtAQV1gjIZd1BhQs+kPqbDofGArjfFP0MrW6mnynhGuBEtAUKQlEjrnAMw+
/vOwmOctJ5CL9LaV8ES28yO3GD+kdbL6CZ/E717F89SMozupeuNnld52uNU0O8kh
mazBnGPB+nDrmEJsgCJ286aH3k1yNpo5Sn9+J92+2ESpdnVnRWKlZojIPMwWVTyB
PsBDlhdFSkmuzBdV+y/PiJQT2pP3UerZWIvCisl5BEadAF7QporNoxZ/VH1HOukL
i2p/FVnM9gSL3IBOs+P43SCpQIHBL/SidY1hEZp36cmMb4wyyOJQX65KLTmSsskm
n2PPx5R9pLB1l3PRD7SrcsSnLZUW0tiEIg5J73BOHZhFra9pTvRcfR/hTuSH1NvH
1ZFIsNb/NkweRk3KyZEJppJa9z83f4igNpHRjwbZ/O72afuv7cakqfdMyME0eIRN
mNEg43fgm/PhkurmqNe0khWTBYwWTcyQ7EppC1atpLP1dafZlEY1gmcTFOklsBIZ
Ip0wdLi8ec63dWZBx5vHdt0E3dbNfIZoUW8XTVS6dI1yp1ICTA0RxKb2JNM4EshZ
Gw26uiyftHIRSvgkdX0Q+g==
`protect END_PROTECTED
