`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
901PVOZCIcq2qT4g7PHJneumsmz2xegtf2+MaZCR9u1lqHk2q9zu4qm8+OZi2QW/
O8wGsvu/MJ98M8FzVO3ze812o4+Vu+K9K7dx6NQyaVjpoY0Xkpc54V3FRiZkfqvH
TC8j9/GdcJ7FFqGHnDUIM0uW9M5IOPXWHgZ+DYpIRVIzM6xCxNDTxLn+rWaWzI8C
4+49huv4yM0IZqjBchT1Ecxnt78Amp36oZodi/vfRrUtEifWMXOfD9oRLxmfetel
E5VfRiXRHuj+9P8E12dvtHmQSXEi3DFjlArxPeAZ1U0zTNz9NmoqYaGBTVvWDbSD
8iNaCcrfEy04bIlWp5tuzv7z5C6hrkc4BBjsKLvbuguhHqdQ+UAgx0v/Yq4GfMla
0pmRz16K3c2Xyku5YAFUOvUo8mElLBJJnIiCwe++Gd0PexA+GoqfM6Qor0e9s5pt
pfTKELKWQrlXet8KIrk2vMp8WgPp693bxFWzpC0MJo4Z0M/2/1Z94OFa+Uo2JqCi
m11IjnjZMPH8TiISfATfugDM4g8Yw1DORcOkuaa+tcxseIo2TldEcgbnoYwXJNwk
GhtQUxzyaRTJy5FVJJJS5JUB7Xup784GiwZFwTfdVeCgfZzMGHPxOCH5nm3cc0aV
8A+3lvsFwa79BSiry/NCnpKeFzfYVzRIiriqNRKh3JgVKj8IUO0GigGGOlhtTQLh
vGze2+ReMaEHM9BxMmsxgBhxxDS+eV+4XWRFY+u8G11HMseBEr7jNwkQPn3cKIx4
jEmMltKpLicwjo7XakmoM8AtiBLrBtlGJIK+UEuaOuAYJypbI9DEXSDC/nTRDaOe
hdn8P/UJ2mepHUP10qRIa56axE+Jd9sRUzewOvx3wdweBntfM6bxl1YnaLZ1KQUk
mtWStMsJHJnUz7dUet73aKb1ONphm90nIztWjquXvn7k3fieiMmVn2Fr0JSllsLO
5TRcDWMtdKvqpUjpW/nwrDKMaxGtJrX9VNIon6cFI0xn2F4SPrVQyCs3WtYkKKC3
g6EI3JRgfIDBg6mpnddP/zSO2WNWsEVVk5tum/hheNDT5xXYIlUAwAEBh3mE93Ot
g+ODRXagtvTXif09dcjtIL41K8KEe4eW064/NF5TIHaBEKQba0mYblot4LoWP4t6
1NELTajLz7NZaxMku06NnwQNShUGI/wgbVMalUdw7Dat2fAnXV9R633ri/ryqXqy
0Kp00bJ+yovgTEEXG/BGMnBcW8fmELu4q11eOCfjf2+sx+qCWcOUn3q2ROki9jTz
22EHxQEYxf2Ib0gIrHDGQ00IAdtq/MIaIejdwaCdMEwr0tCQzNdCuuu/sB78m/8G
tmZryuLaEeNziKeGMZqM5DfJZ9cRR2bkRGKk9GoD7tmnSywF3FREQCnX31zgwhKj
d/x65moWiYf8sGZrC0VfgyoRwrcK85lb6z2J9Y4tGXtLiA/CtOG51uRxoH7O8r6A
sz3uSbJoT45j6LEXVu4cTpqTAcHWp89QfwisdypUt6dlYnjB2tWb2vJLiLJOBGCQ
JSILeXL0/XS2itYdISmGz/4mXSMezv2d7gZSmEqnUtEZV89xL5eObHZ3/Njn4gSO
tHP+SNbupVa/2Dk+2r2YTo410P8VxgaU6wJkpkauuCYctBjPpZxEbgU6M6BL2DcC
tptCynLrUSocno03RGsp/Ipb2MmGM1rSqQ4zYDBdXZp2ziPKR1224Jh3bfPzQWsP
9+waxasGCWGQwgqlSaDnGhy4qzYi50cO/C5Mal1jxiAZPJW+MV3RSVmzGiuDRWXk
t05gDQ7AC5VcvSWnEadgsj2czEsRrAI0HPVkJLa3esNE88gRTjgnTMSe/dGUACWx
3u/P2YPjRzkwzv+00JMY137HynLVW2GEadBLe2tFvOrp7xPnQq7QFr6ScYvaTQkP
aHr2ssej+0hHD6PnX4EUMK2dcsEi50zr0byUMAG70pdFvsMXtEQ7C2IpgODO0grO
FUrS1giAy6W3lrVxZfqNSan5tF7dvEAptXQpmpxYb6EcmpQ2NINYWSsCfzTO0YUY
gU7LYCZ6cpq6mg5zTr/uXxFJhehDz/6R6exMFEO/ktN5xnxSftt/o89YpRmdoQzz
0MmWXFh/e9qTAW4cPy6xDTYZTqyEcnpH77nJ0zNH7uvuTwv9mi+QJAmjQUs/1V3N
kG3LEUTFRkdT3Z/56gf52xzxsSdNaeUiurkpBSydMeD0cz/LlIDg+tNltyxwJf5S
vnz8eWaZaMomy5flT/PDIMNZybz8OgHxwiRaEtIa/pq3bWeI4RVuGi//XYgMeYWI
JW8nmZDR9ocQAq9KWTEZxGhGRErw2/AwU6a1A0qtR45ZSl4Ya5NGR708bZpsB/Pb
fIxEm2uqyQ8hnuBdDROf4PvO35sfGI9AvZzhbvnQx4gwJIaRC6VAxeyqB6En5/ar
kzv0Dzp34UmSA6ZmZ3BDnR6LVWiyEdjSlvuvNxv1K7zEqfdL7b+xWEQJ1oJ1Ukw5
RFCg6bt1XQkOtv07Werx+b5chHZM3pB4BPshwwahMz3lt4oGOmPBoKT1Qnigfw7M
7uRFCaf5/H/mMXUeScMYfRFfnz8jE7zx0vBtxtsH+blWQ+HXo/+SghHunCzmYsmF
Dy17Y9ld0YPEqIKvfIGA0Mq+UXBbJv6jODlBz7t1F48zSQV2mAPAP/JgTYxIZ1ZT
IdZu+gEYTfPmZk5ebNH+BBOR5cU4ocfWyGkBSFHghFJKadCIjxb5lstuLHjfz/A/
6DZXXM0TufwNHij0xAgh5URD/k87UPg7d1gUls1RmGGMuHlpzUEDqI5MYZet6RCj
G5Jw5hmF0z5NoLMhEuzVxkuczcOYogLOQ3x/59NERZTKdlqG0WpfBf6tIO8kSMDn
c/rR+g2lVqyxEG6vWaEuHxhqE0crEGOw21Vr5nzJ4fFrVq1dKld3F6N1hEdg4WGV
N3fEkl3MbRRUSQl9Dym4aCY6IHwfWTc0Ize5AasaHV2Hnq1xNW9msE5OsJGIBJkp
omTHyCH3hGQEMhidhLTAKqdhhNj9GAiAE/B4/jTsltmuxXJ+5Rc/XX+GjlFRy/ui
Gb4Szr7BgAHxEdmq6KgZvL4GnskPo6kGalKEPWXQB72VoJFKifQIhUZEHi2LrSiw
/M7uSAJm/FOpP3ECDuYlbTYt1egCSUAAMngRuTMFHa0Gt45WPETEIlLhlQLh82oZ
xkPx6TA7oNgUYWvhNbQzTUU3iSIWLDIkMxlopfyreB+LXhpDSlInBqgwySStcBiO
lZtsSYhG0QiT6ZFZq5wsikoc7MyrePFeQhHdUyJCL3+RsacmbCb9SSYtrqQalyO1
bfXx0jVUl79gRHJInCJ5hv5baSvcmh1By4QlbOuxg2E4VZMVLQNugSlEn1bbQjvH
WsSjWkCG3CN+lkoCaHKt8R7MkE7QeIx0QthWkurl8jEYeensSfNvWV6AGKwe5c4i
aNUsM8RzhMPbg2vkPne+AaTZFx99crG3R3Y8OaFlKqkfXiF94qTDFh2eFjg6naD+
6LpQPPfdrW6xX/wJZ83EKnivoUNEyxabpT7KMZ7HUmYuzXg7KvZHhNrzpmNf0veB
786c3MkdXkmTUgZ6FcJvxnZ89QJggW8HdCkw3Cf4CYnL1zqK3USNj672+xfjQuRD
+jNG6u5/1fXW2lECHJGGclP3JnjleeviV5gAD5ADLb9EhEjWDPp0XEQoKmrOEbAc
F3610louvUL8jq6IultbWJY18+n59DCnYu16NtVbO2SJSPuBAKXTAd1lMGlWtnlz
gDRLxzhE9SwI+bIgjbU4kclnpBW03Yon0OMxpifwJo6NvlcBZek5UVzpcdUck97d
TMjeH0hLKCtnUlsIJO1uizYjKgExAjpI6l6bnndWxMc=
`protect END_PROTECTED
