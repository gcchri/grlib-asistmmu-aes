`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mt7NDN523n9lOPD18XCEChf5VaJvU3t0p7TLzzw4GlJi3V9tbVBiAPxf4uSgUGpp
g79NarWTFQ7PXBzJIhHj2B8vYfKCMeaY9GH9gg9Iec7a5ZFng0xutNgxRecOeYU2
fVMi3LeMc4Eto4SMmadWKTWHxf+wW4e0jv1GutxM3v/5dZVbw9nz6NJYrceR7KDF
1ndWtVIDab9fDT0VZ0dSPwDIp4pZ963KV6iH9ZNQlVolb6+yvCSdEv4GE8gx24XT
Mz2/01fxr4WC8x8vqxdJ2Xypx/O1NeOMxGkSQ/tRav0=
`protect END_PROTECTED
