`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TTWvurBd612hsUnNkme75UfMqRB0OnEq2Gh6Qb7muCQ/M9HTEedgYVSEZoGNGg44
a3s3+9JvXfzVL+2LR4hEDnyBWcGlgCHzvVO7d1M3dPxRlOp+hOM9jDkUaEWbvOo+
8walHVOEqpmiJYIlrNe8t7M6DJinlqe4CJmHW/itqCEcIUod+Hc7cREJYN3zDU7T
fGOA6KN/xPul8tdxwHh75HeQ7+9l/oWC9jSLAxmZ9Fa67sZmUpJaHPhjNxKEz6+m
0wY3fRT9aTZokNVZbyv/TuG4WedR0Xc5R30UwYKn7iQZdT+IdlJsA4JK5qzXdXeM
Jz3nftjp2/BOGVgUxJxXoaRTYl3RxPA1f5FfBjA/W9dDKtH7pPesrvI7aqxBm4Gj
EDFLCKfHUbX+SoGhN2CHzvxCEsuckfRos4fNWNtI3N15r04+yyuGIvX2dJtDvtSS
MBs8RcxmxXQ266O2gz9a/IqRkahrT3yjlFOFLUSn/rlN5akRFIXfu4xdsAlsc1ah
3WoOOlQ1kdH4IokfWFsCqg==
`protect END_PROTECTED
