`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jpw3zR1ZdVkEIcNWDbkJTOO8D/cNJwnI2i+iY1z2/Ia4yDE33qHZUOYqYFGmLAFD
KXKRmuYK7bQ9StQqMrBhdsFY4eNrAVuZCHDAsz04wmOSp7ns+bZlGmJtRSZ8juun
9+mTYd91wuRvxUg84Z81kYu5pGW528mS3mbbSzW4/r5d0HPgid6SaoWVdXEOpWKh
T2aJkCit45pehxz/XbEC+4v0PVziX+4yP1hZ4yx3rQiQhaDTr9hDhl32DF4tm5ti
jkt7i3w3roxH1BG9TIJnHBK4N1fg4hCcsuFCVLqSzCLxuBP/Otwfe6xWVKldmpgV
SdZwfXMGgxBBMgHAiKIdACVCpi/rHftLIvwMx3sMsWiu5KeD1GTlgld9WTFJSMNX
ty+8dwYfl4ZCJ1L6Mi4oEkkhDkdenKLKmHMB1iFs5rBUVljBNvk5ftIKxdGbcZmS
MueXpBg8h7KnnwXTh2M8J39NXC3gNh/OGlTsnHKlVOPKbzvUFdBrAMX3HoOTST1F
ABwzoKlXofvAux4WUvaILCKxOCyioqvYdcWQZ94W8tQt8LL7sfLqzcjj9/rgT2uW
nvSKaY/HJPibctWPFDO91BgIrVJCJgG1DnJKxipPlOnCRXBoQmwlaHUOsmYkRLed
AUT8TH4yHcFblH6/zbAFUcOTnYfEghlpBX5XmDzfWixGphUtJfgs093fhcWD6r1f
UPcZo74qCFzbQpHA5RHiEbBWrzZ6sU3HobDB/CE5AdnGQJwKYbW7a22RbemFi52I
cSq1ReaZ1iameZEcFdzdUPRKhzO9wSmNsYC3Xn9qFBT8Of7viHBd2wd9iFguP2hL
ie6M3d151Hq+4RMP9AI0CrfSBfDQaidGI6NqNNVlWevZbznDrvtbCTn5c3napCtN
F7Zl3USUjeOH8pOJylnhkvpYvDGDhCKN6gt8QxiqcTVzSC509eU/JN7rN15kR3Bf
q9OGfe+4OJlSo3Ofz6h7JaSt/1yuabQxnIgNm0KY9ex2XRGZrc4FdUV8OS9n2xO3
AiFRXKDFtYhunkuRPWla2T5mflALhNK0Scd18h6mO2NR29/wcn8qEW2sG7ht5rCJ
C//DXBLaLH6wuFMv95KkwUl0ZuCZIef/wj245YxIchJ1MBJW7Mrc1bBKrDeS87jn
+hm0fxwhP0AIXE+IV5acqFwwMJDZ0Xu4Lz30HTl/ZbOIa2gDQYisnsNy3WAe9HS1
vjHrWued9CN8XKRbS/OXxFKh8m5+K7vmWkGNXxhddv/AKAH7A3eWkcmS/dvwecGp
lrBe4WkM50HvkdSFQC9PgtiJpURWRflMcIZqGdxAargpVWacj41Z9NfreoAfCjvU
7NPsQdf8pUZfbPiTe8gPYFkFQK6M2SZK2ESXgbopR7wcmtf+wSzpMZcERTq/1fgU
kbUjVSJ7VAKiXsnqslZumZlez4gO/BfVoC1Fsy5kU0vaq5YU3gr/Q6641/XuZLxh
GiT613emftCNj7NOkyfVJiP/zTEyeMjBUYQuI8tLcBEV54NvZgJ6BaXARXlYPpx2
u1z3Vu/aweQ7QyE/Uvj0372xHfh2F5hrCKneA9jPSbZj25Q43V+Q9EYGg5Pi66OU
JYgzACJKZ1D3JpICi04XjSe15zoOJAkkWMKxQWMkZgzasVQ2y6X3hKp7J+yodRRa
0I+a0o4OIl1aNSEgdrzNz82/rfTuDDN6gF68THAuNsPoZP4OKUgrBfo+a8Xi6pKz
k8xeQ/EnxyxhFdTggWjm8UjpdwX+rwYpxQoBMLZExRtU7GmCfrtBOxLEzSKjQ5hN
v2WWGt9H0ZPn++E8ULifldsFGLkyTExr0u2pze0a/F0w6MKH2zvOyUIJzt5srmPN
mlxX4i3dU2LvVL4irMh1YDeKVzLvFD8BIsQYMZ+j46y5uiT0krrcigadGmxD7jMy
MmdkIjf2IfystnttZN/rbEePmHhReX9Y+sB4Hszmrc/j3mOG89rD6ZDFetqoUhT4
MV+bkah6CVTpwxMBNKlud6IoWnjwwgFfB2E3JZjhD+SrA+EGzZvSAWxiSlrvAgXs
BBeV4jGCLeUDHmr00kbtfvojdx7nP8KE4VvbZD+OBUHfbRfqdd/JaeGaLRUeHuDs
Bv5H/ZChg5U416E6vKiR2RMsZVRLfgbSpn7RhEu3Vsc7N5B5d0OIyBK8LCBqhWdR
H0jP83u2zVWAJcLIDn2tY1Au/+vZhBKMfl0n6Osm7n4E0MmhSi1vpHi0Lxunhioe
jKwOWxGKvNogL95Q2rAWxcSo7gNR4EVofOy1aeo1//szeX3MmYuLknrAV6z/6wDs
9ChTlWs+XJnrBWppXZ6z1pxNnylX8xQwZ3htNbe21T+KUO4Atl5CbRW+0GYrFO/9
SFa73JhZw9S/cN8o9trxSa/LpnOaw/Pk6Q7wgw2fr/4Eat1hs5Rs78fgfQfQOoDV
q15Ognn0LECR71XYQ0b4PO8Dj26lAqEZiiMz0lqqRMFgGK2bFKWrqPwwgQ1IfEwj
nNkkvjenvTWtPs0v9HSr0ufvWFFqyraOP9iX4CYJ2tjy6hKqBvHMPAfe8uN5jD9j
qh8q0Mc81sDQEGsVDOWi0LWLoUK8TQhjFF/QN3RuT96eBMgQHC6ojmx6nPhP6Lg/
i339vrM0lxQzOvWSOAZgx95nwCevb9K6Z/iorfupIAXaYKhNhk2/ocZjy3Xd/tTT
GHUj1QuREyRiwkgXcyUJ9H7XxHRrG1pFMKCQExpWVueNSdD1yPWhu1GMeBo9fTgG
/2ylBaKCeBKD6Tp1bx1bkAdYPCr4xAmZI7NREVAAfl6kfJ52+YtUHNayrLS2qNUM
Zta9R79qahH2OKoCOrORiZpvpCz3Ug4laPX466J26flt9aei7h0NpuZKwhDEhsvx
+LGQSpO89aOjqaUxcgfhTM4xCw6ndU7OrzujeJ8DFMUXQ1eZ4vQrmedoaiROT+Lh
nvploXZkItMGOa8RxKRtQX7aZDrFUP4BohVZKcqE6GyU2euC5BWpktBRdKnXSx6V
ecNQAgDA19abL4SvHCOlb0FRxvKy0SLNch/zrBTtnxa/rmloVk7NclPyW4qv+4ZW
YQ6MFjScqBp728zpXBsEQhGmwx4OzDeRRu3oRZVeA5UNT/uC2iNcveZ4603Uf22t
tEJr3cN0J/7fe9MdR7wsdqz3WtOVMicXHq1PTvRCC3QUg8aMAtYkcev1a2ZT9jg2
QH8HePorwcfdFQyeDqBGwTeIzudiwE9gMdyMRzS6RpaF2y7NL6G8qmv6lTDc/3pd
GPN1Dcjn6qQ7ABCSWPGup6ADkJv63OfJOkkC9VA/vsiGCtzMX00EPScOBAJJCRsG
Wdz0goGvUGdmS/GC0mCCjhArlmCrPJQla0BYtlMaFgR/pGqUzOmRZxG7DSb5lFTn
JHuSXftbwlY8DeW/rI18u13UDudTbVS5prpT3BHGtAMn9cxogfamhsXPT1EUXjT2
Oq6vrgAdD04t0XI9VsKVFGcgDn0PWko2QRw7ax33NF6JdnflzvBPLGP+ZDeVLqT2
ExB7GTWZtSlkrInkNERzeOCUgsCCfWgbXi2NkXyi86A89MlWy3ZtB/HZne5wek/J
ysji28Sbylz/hpJJeReOJezjD7LbU+5kKBC/UDRTUcX03rfy/a/v8xQsPdjbqjim
ndooaFjrj19B7J0tWs09mcXXisTbaB6UCH3MsAU0nUo/AeslBSbWuBk9HHEI6W0j
hRSv15uvVOZI4SWWH5lR629pF1cDEHNUViKZ7C193Ja8R2rMtJha93tWajZRwt2s
oCpzN9hsF3aasy+LlbOZvCWSKWXT0QxYn82dwFvjzLyAtxL/1cjBIb6KoE14SbvY
ZwVdzvtbe1MP8zWQRWIERZSKlBa5Nk9p7h4saBmjXp2xV4h9DmmLtuS3Wh6LMBXc
YvphzlokADrI0n6BJi10qolsK6x6snbV1gR7ERr1xNLCFOADJI+zQ+y95SwYqfqv
oSrqIifwKXUHc08olIwP0oGLhoY3X4AbCX+BYrDD45CMP1A1+PaS8mwraSelOsHd
X3WRKzkQs05RsVIJCTcAr7CnBZmLT7VTIAw5AXf8QbUDEd1ZsPb/++VSuUgcWdmX
lQgI91+gVig1hGCPBUbtbg+ImDKUeZQ78iq5hfCr/0ZBtxZR1iURCMoSwnS8bicb
gp64+3YWorUK0GZttS9hRrBhcWNp/iMfvzzu313pWrwbv3aH+r2JQpeZbPA61CoL
O3ndYazN4BFx1xLNePYXzsVo11QWHHb7YljspqzAv52o9EmHQXnoMaTJEmBkvukI
ruJ4/sIzHxFCuPOUN9aGGPP+B3N1MIB357V4QuZII2w7mt2nVlqKuHJl3jFeJj4m
+i5mpGDT2hWYlNVQLxRELkIsgz6I7R/CvasZRIDZJPTOltsAYQ5HasbqX3zT9ywC
GrYyMymrUfu2HPZxGYWeCVFEg8vRjz9JotnKiSgIqOtiC6NdBNVUxm7U5NXKlgGG
eYJ3I75J4Z+bBzF2PD+O3d0ZH4ivTR46wTGbVtfHfpOkOLVZM4V39x54owZMPiTd
2IDfVHVKMb4a/M+HDZhJwJ4xq9KnVoSxrGyNLkPTFqgg++wonjxvblu0YxSyVZQ2
8GASsMh/HWLKu5B5DBIqWHxUSHPzXEpwkXyZ5GcycVXcN/Bu+Yet7ZbhlT+G55Tx
SApbeiL3NdaOI5l8UVa7FlElekgs1fbU83rm1Zu9PKwQ+j+MVeHJmTUxHEzI8YSa
jGsnsxEvZ+2a9Lrhf1H4L2MDevBdbj+1b/WYiI8Rs8Y8hdKmlJHJfRA9idHF7rC3
rCgfrGdIuNMMg7DKJIX9OX9yaHhisbu/k559G+mviyvCr2WZ09zbxnUy09/8EJUj
6hgOLS269oO5V/coyfr9T2NFQggG8oGAkdfDw0YqmBhKaFxrESzMpz/vSxD/eDnW
CV79MRZryiHduHgCHJ1EFO5QqUzrm+o4XQz9pOOlQEpIxx0QqJUNwowbITO4VTF+
lH++3RE7Y6B+gEbQ5Tc8nyrFA86Iy835XCWLPFbLIheswIHDuopBfL54CxtrPIbH
+leoKYfieEkHMJt0cJFwb/eNtahS7tUJWoCAcWDNQYxNv8CqKrYblsB88XuaJziS
iXVp9Sh/ke5nOZ0e1ns490ATSrxHZ4qBTHmRF4FdEQeyB0AGY7o/m0LDAH+v7HJ9
u5SaGR8okDsbm8uIK0t1tg==
`protect END_PROTECTED
