`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PuQ1znqorJEwNfPxWBEJNavDMymLDrSVfmsxBWWXO8THCcjJjln6jA+1+gzKOOyQ
iXkpqoGG3CSe8seA54vQDTAfdG2j4/YVLhiKTr/1YeFesLLsbQirA9Ub/jVes51L
kLKVULISkHhDwScq/TnaeMoSzz6N0UyeDIIwAd+19NUFp+VmFzHnIVeAIXLIs8yw
lvep1/5E5Ht5efyiXBLRntAdHJnMRZ7uYv/OsCD0n7iiE8G73htyXYTLtTFwzM1c
1HOWqdJr5ZjKuBBraIWS6wwGgkmEugzQCWEsCiysdJhjOYSdcevWrIJDX1LOrqon
caH0Y9Icz6W37cdJ9XP76jzhIzqdiU7E9UWKgshGeZ8ln9xUgGpPZj6g3YY/7Bys
5xitnr6eol1RfqX8WQKx68kkxydMbYB11JU9dk8muQc0jhMtlJ6IWJozfPbT3sJo
OhFx38rk1HFXEroW4SmTVtlVbPkmAODms+K/LJJK25lcJBguDkpMM4OaNB3WRWEv
lkPiPjYPM+cFwyJCkqIlRsilAuaa79oYr/eGZbOJ3gqK8UdmI+F5cOvxy2wD5bTx
/CcH6iiZ2fEPTAyPPC7ednvZ4+bnA43yzz3QCiNCZbkjMISKbLbU32CfxEjkCzve
wRZeVz1nDqiHf+x3xwMhqQipqEz0eJpfJWxpvxm6Dppe/YWqahFIxwpoVAhDKB7G
sMcGjNzpvQOEWa5wAGYksyVIMGVmXQZ/Ujn0PYs5YueZV6XBD9Az1IfI68VGxkXX
G1aZk3ruVBa7YxmviF29fVSJxPwrb5UiXYfeiuzBeGc3KG+eBQrC3R3pkbaAO1WR
G2z3E0N5kRBAca7FkZsyfSX/c+/xYNL4uSM0lzKClUtHcideClmRAh3zQp47qa9k
YZ+VilLZSIqZSYhQP1+R7LhlgDqSxA57DkBEDwbAzJKehWtefcZBj1HTOovVmJ1U
cdf+PknffUHeM7oycHe1MtSOLkyNssRrF/PoJKabaow=
`protect END_PROTECTED
