`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z577J7biMqt2ZOnY3ME/yrxtGohUG2DPtqH7kdP1Uq0Ywx8oMaZF2cGcyWervHMv
vnT/Rh68maTEgFYqil67Swi6jnCBmvU7F5gpNHjcLd5auG187yJ7QNIiiWXKE4Jc
KQrAYcAFryuE7o7s3skBUd733r3krZ5T1+AhrNR6avCm1xxIgER1m+Mof/R7I4yU
2D1uGsOcyC54w1Mx19JP9KRM6MHzI4ucs5zfgSXx22i8LQ0s6VtHnvYoPPN1Fi8+
o7kIHX+IvYjxARa2ftxTE1VX6weZw5M4ipABWHSUbNV0edFW/PQS3V5xlqeg9F9J
ZnoC4mUe5FHdF8Y7Lq6ijtKQPAFnt8Qp9xCdSsuBMeQHAEn2OVPpaZWcYy+2GiYA
W1GDUr9vVPSyGtvIEplNrC9qFKlBF15CvBjHEfZI3R/FicPwB3I5PlSGYavmWdnw
fpWObdRF9of6TmC9NjO+nyUZVxQU2LR0jlxlaor9MZ1mTnFenVmjN3FZUXMDYUo3
DweOcDeskLRC1CP8iSYtGMx9g0Ub4EOUmRuJsu0BzkydrIzezFqaxLGu2PU+Sc60
7UDgHRi/O0c5aNxq2a85zbeZR5zU51PA5xldUrwFJq6WAQX4yrak3Skg+tpckCC3
QIObXBV49X49QNf+DZG7p+zt0E0L+YbIpRZ0nO+T8eMVW6gzYzCEhLubrK/dp06C
Ac0A9HlThTf1X9d3AxF3ClsyUHWf1fBstWz6bz0YDtO6YR9Q+7YKYO5YHXGg2bIv
YfdSZZ8xTaVsMNrH8vG4W8fwxk7wIP2Ad9xw1mRfi6eWwG3yMtz0lsOhdgbRnzIK
ToRGkh2juE2T/ByA7jM/2Eqbfhw6mk6FH/99BtPVN/iSv9dv17n+qO/1h8bJHHUF
RgySZ+dRFgprg902EnLjL/wcmoyMU9gKLoFE+xDi3sdMVseohhFJzyyMv6PXLOdd
`protect END_PROTECTED
