`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bU+G0VitQWImPsg82tNkddbZUQp+ytwcm24tChyFTLX+flKrTY0BknJXyK3anqGp
rQiLqwn/hkyXSpXATU/V/n2zI7HmCMnEjV73apBcGeZAriGWxJWqVj3QW2roXjnv
tMB8o4zsZ2qQ2Lb7vtDMAPs7XP+28vy2dSNq+NpvkqyYHFfaRLNtSGpIiTjDDF80
EEUPBfQBfUtmnlP4UnPrR1ySaJLiL3YWbj05YZVqvV7cbMmOF2icxvSk1N7SPelE
yyRDyW4+pm4YpCl/urWLbqiBCJHb4EpMdeMcUwOwT6j+m+GqtX/tAvvFtNhixvB3
OKNrUH58rJF2d2MIlKlBrO+jPuO87Gt/NYd15/nYCzja8x2L9GJTs9UMHAN1zm/n
tXNXY6ViC3tpMEVAar4ofj+Vr8DXDb+JHvD9GVW2ouP8REOenhH2JyGSghE9WaHS
fALWMIGQE5SYNEB0CN398saX3Q1LP9POlU9cUBgGOJiQ7XVPKw+daeZj/7VXJZHh
6IQ6fZ5afU0khJ5v3oeEYijE1tESal+fz/iQfdCig220PGYj+gDz/cJqhO+QJVdw
G4hfmaUbfc+IB+D1eck13/W9wf2T17K72eiChbBCrNW/y1ROZ18rhFG3czBPwSM1
3q4gRiDCQN8VtqcbAvCQqNst8Ryzgfc9TPI80qLaogox0cGx/ThQGTpxCIzVjLrC
re9vUK1ExXYoD0ZN7ZSsRtvkR9eFxQUumTYVS9SHXFabott8MVaUeGF8eAslo2mZ
l1HuaMkD8+8SCWrotHGrO4o2UObyTfz2CK52E6Eg3DSpGmCKBaP/pYbCcG44IkU5
c0gGAwG5ttLrknXiKaqjh4iN4Rtd1OmhvfkTUhxgiMkaoEuE5exdE2QcLeAfY1dt
z3q/huvDNZPROAIKYcniXGj9nNjgBD3CN1jXzpehj1zxj9mKmYX9i7QWd3A0imRS
gtH0IAPaQ0LA08S5OD7IH1dRBODAy9Lz6ELbblKWWr6BNhvus95y7A7vlMMjNc4r
Uco5hEGg+TcFy2O99DSWzn7uOKxYdfCe3wgS00rroTN2blR+RDo2As3XuKOVysxW
FYqYxnbXKaG+MvIQSKQ8IXHQk3zHisExr9TyaM21IJMqllWmjSRwF3+KgBwHGYGV
Zp7C5ul6yFsE5ivanYA6Sl4zczuJN523AqXH326YVr87h7ivIGRh1HSBPnbkOnwo
`protect END_PROTECTED
