`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LDxHkKrbkIDaU+6cYSk95QMnnLc0v/0FCYKajzFEHWiaTXpjfrxuoYL1fVR73Gcs
Z8pqisqERCU9PDb56eXnDTcTkC/zKpjqL6mqxOfbLx7l471HMki+Vg71biTCZfkZ
LpRQ1u0GVquwe1gpN0KIq9qUKAGzsHxf4KyoWN+INBJSmHQO1DFQqXFyrgBCCH6u
5UrlIWBQ+/hYOCxgs+5FSBc8w2GHfd8jEP4slibzLRxgg+JwUscXUPYvs+sMx7pW
pjtIhcJC1KxwNxVDnO/CERIDAs2g3b9ACL24ezUymyiYlwN28q6i1iVJDi4kvIhV
KxOnWtP4JvEUX/TjvDu0KQNK6Yj+kDOkdQBBlsD10/YPtgiuBXlCsTqup8E+FN4N
IXD7637SUGDDxiw81XdRq8wzzPKhLQTh4uxSH14LxQZBMs92LtJ4Ov/WVXE2vSQm
`protect END_PROTECTED
