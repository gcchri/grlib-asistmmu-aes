`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1jxdg+xakY5n0J2qQVzjYcIWkYZP6uOo5N1BW5IMdRcTGopSoVs8/h/1tiu5p8c9
AtSyMo9UUYBYCogQgP0MvSxSDdhhGsdqoFtuZaEJI5AUmYvVKz1HoD+vbjAKw9GY
83cOUJ++jdrqGunXxF36X/6gFtpnJnHbRF9A68T6CFtSmy7j+i+dRk1bjwDGb9o1
LTbbOpAFDOCBi1/EA9gTAgEpoLaNaKBOUGFH+voS0K4P2q9xTLQz5XRHkIyW9xt4
LQbTyFGsqJKRDfOqkmgynRO7TRmI1TXGdhDn90Dk9zNA9xNgVrzEs7VHiJI0X2V3
z4CYlWcAx25EQt++HnRYsh3IvLhZrIcox8UWFI1s+T0vjb9/IETL7f/pUq1t4dRb
9FgUrmjotdgVyA/OhACoPg==
`protect END_PROTECTED
