`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FlD+4j56VI2fouzeUPzhK+wstcbmLNI14ORJ+9NRjtcEwLZobpLNelKaa1j1iPf6
SQmAa72xR/sQLpvq4Ur66uVTK65bLctMqtxsK9uag4x0yvaUXgrNeXPgP7Y6GezD
f2FpJQIhEOE9g6amCwDQh1xoiw2wCCGJfBY7StmkIaC2HXbcuJo6DOZUTwtj+1D0
noETUpPiQvVnfdD1fwoyLvyaWc7WZ9BTlhorfirNomI8uyyYNv3kiPFN3k0lN8rc
v4bZyv8f8Ir9aIUZnl/pwPHxydQCmF7ns7SjAr1UPGlPx8Fnnk1+dbs/4vAR8is/
X7fiFujQTKJft0BSxqHkyu7SOXJqxFwm8aNzNDgBAV17pfcmW9fywvUsI+UM0/hv
Kbe0G2UEWnEWF43pmBXElGsclurkZ3rFECIlqOQ/ADc+9xd6x87BKVfLtgHFQICL
8oD5geRqYV4b2PvXBDgg2PkeomSc1wqK1UPdvK+0vwt6q0wl6H4TrcKoEXY/Q3u/
XrIhX7byxup6Yo9ttrJJj2bkA5l8AYuAS0lJ8NzcW1nvRH1UcDljxXg/OR2sdAr+
RRxIMXbzbEjzJLXZIE1RZIt0vm9MyNff+pwFKMLTQJj/3Ev7M481Aga/SHXFomPv
VfZK849Q+Jzt3Egw3gpf5sLvPWukAV/Mll/cwuRbqKXCh0BgNhp56rz1MB+rYnNg
6kBq9yuuGxqBt5kk0fFhyK5N6d/KBRdHQGWFenomKOTEegPiw6jmb1JdgFoKlXPB
WKuLNOCnG1va1skAXM7ya9DJMtCLxxh+Y8tHB5lg5d/K8BrBJMnEws4ON7J6BNo/
6oYMsbOkH8skDcr6zZR/rU10yIJ7ydRCLMnMacmrMDYLeRVuCf5su9i+jDaF0jvS
saQxFEZGXJ/xCahzoQsNYe5uU8ikz87k3SyfP/Ce53XXKrxKhsBXf68QU72zqA5d
wFkFYitonY0PAfw3bl1rhDrRIscGj5hPu0/7IAS5YWrMDQuJ4RTxjWHR28JXKULp
RJYSK4N/K28/aNVq2/IfI74cbnsJQkwP0aUkAC7H86YixbJXWnQg05QtFoxDofks
Ao9zHce0BxpWIu3oCYJR21gSJicYYig95rnXCX1OFK4lpnz0LRJzYgs69cuE5dr0
/q0znYnnLNddqJWKSZSaCKdQhmatL2miJ/zpyFCxjBf4FnC7ICiqQAD5PVoJtcUF
3yPR+Gsu17mdGNZsbQpgqRo/weDDJK5auAL37Rmcs+JobOKXza0sv0piMVM0mT9Y
IfrPlKiB+iARwcD/Oz2OaVNHHxeqi4coBN+VVQonhJyTA7MF21WJhVolc8pew3Kq
tagJMCEFjE8f1kG8Y5+fCyfdgZhn7BqKvYZG6u5WTBRPdIs1HF+bEKupvVswaNi/
9IeZvl6X6jfeuEXlr/B7iYqNZGx2v2PZ9p0ETrLLw2vSpAbvGmGCLPI9H2ObJb82
K9mDEacTGSB7L3Vt6IX2hfE58sLIK3EU4XbrWqBYfYXx02vb+rfd6w+QV9PI2SM6
gYVzPw2hPW1TjorcYQVWmoPsYMQlhWWQSUNRt0CLepEo1lARCKbfz3N47XDk9V3L
kshaa+IE5MUgFR0oaAvrn4wsbKhKE+DEG21CFa1T6GmDL1JssDgID5K986Cajz1n
NP1yhYorVWaoXMp6WdUqDMjAzCBjSu5XCdmVwbUEhdqkye/PguAOAUVic0efG0TN
O4gF9feK9RjILFEsVrngMS5JP4bQ7qx8ug+pahs8q7+zxtNMx32QkvcA8+E9nRcY
hG26FEHEqIo7UlHNV9zUzHE3SqjDZsAWryS0mUoapxtabviCOMjRLWUhuXsYf4t0
6hoz/rO4KNe2wZQElI75TtyrKQ+Iech8Bb1sU9hvgMLdBoFR34lpbJSDRFgx972c
UK05lnC6e7NKLBCUraHih0+Neew6ELEo0GW2dAKBZGTgd5egFiHtbXAlhfCN9nCJ
kwHGqWt5M946FLlomZaEoQUJMsSB6HJa32GSDaO885zWFlKO+kF3DLwi+ob7Pz8+
m3OSdH5j+V9GFN+KqE0BkNHOSevRGweY99MvezgCEqr5aQEZUicGStUflGedXFxA
MQ3ur1IEFNX7ccQJCRp7LgR2Thg2LBgXGRoKn/iyegHrlSHNq85j1s4IN//+J6E0
f6wtrPJeNqt65FboPNmemaLGJqZNdc3twhtZ7Si/oR8Q0wsoA9grFlRt3+JuQyZo
SZz+T6RBEXq7e3Dei2UXRB8XMFhR7mAdrM45VPZeD6VIogHfBBehlflBW4q66h5z
hllUTsxRSngNQAyKwDjarmg+XX2FUpzVZRIYHncy5QjH5ml0ZKc90IW8Ups7xKUo
BTDZ0aUg71LA/Y2ZJmODMuWMWmJjUos69DhPQkafU7ISChV5w6Eq8mpzLOx+oGLt
6dXq02U2aLQiL6TSX7xSZDc9jP7RCjTUowTYdtMpNi4yBqbPs+vK/kMzPWPZNJV7
jiFQAxPLfohobZn4qcs4kN+oscTyz7YSja4vTJxhei+9KBulP41kasgIqFH+dzSk
5236z0g2Cy/mbGUulVZZkV4pWVReR56FCZ80Iaz7hnlxOhZyH9nCHLflPi32NznG
Bjxy1/sx4mOwuohQF2D4O3HwNTmbyki+1gHU7jRFk4FJzyN4HB++k/WgoiTcew7w
ia8SfFFntVwSjhhRAi1MZtKLPd2pv3LJmmaar3u0FdLW7HgwvoPtPIAdA+t9g9NU
moyzXd8PINIwkgY/dZNoxnj3PMz0CJRA8lkh95xeB6kZZKsSGLappaEYCZzuJGHL
Dp5us2i2HPKX6/0H3WsWQaxPbPyAfNHB4EC18uML4f5zWTyemWkxBOG6L6aFQ36B
2oDiR5P+cyv/wRkfalrA7j2Kt3idqU2nySpjAytQK1AaK3fObnHqjDkRo5Q4vd67
gGhRhxK9ZfrNrr+q0Try2ykJT0AMu7psQ7yDOYfLGPU1plQz21RPv/t1lccVDxI9
yXZek7zIk5KJQK1tk5R43PZNy+QQoc5qkLTl+PcuHOZqCIwK2wy20bSCov1/Ixxv
SV20a9nvWicL6PDlptj1NztbNMil0ugsm5ax4eww2g1RWUXbGnVLk64zO2dPq6OL
4gs+A/FWJlTdpnIHnwfZh4nkEjaLoOEz1iJLaplwJbG2scPVPG7eWxycqVq5NrgQ
cgFG7foATTAVSH1phEBUrqBE9ozmq8+dXgW1CPMME/CsB3GOTImWexS/binx6NvS
yjQmwgwr9atr+u5JGo9XKAa0azpLEIn3eO3uA9AflYoteAfkHRqqzfxZWbCn04EQ
p5qCiuXWhmIsscU0qBWWlyPpdFOzBkEvDQxSZdNCs9C70zECmdZ2pL2bFNFRew7Z
VeOEjTOgsX3ewtnO9Kb1MD9GEcwBKsN0ETPZSvGL/LtKNPgvj3Yi4hfyTc7c+B5j
oyCmufskdj0liaXE4IDtUjtWXdynRB6HBV2g1g6xppjEW8VWET5jgDO6gpG/3/zT
+/SvIFBUOCfSeTODwtXMOyB++DA0FkBPI7Ps05JKttuj/XMVAllylAPActfPh9o8
RFv7gUSS5zeM9yMc6A3r5QIhAu4hl6RtVwr0M23N9Q5DHDwomx2+CCtKlkrpZhVZ
zxbfldVyat6PQZk2ANsQm1i61AmRRypEFB8W6v61a7G6gtcIMt3hz7Msnr7oSng6
xF5uGy/bPDd6MBALQG2+Ln5sFhpXadjMdwgjpQpOju8tDUU3EMCSgLuTajG9bUCp
FfGQ9ESTsh68+6b7yBtpImEJpoOLhsmRC4vUBWYqpdStmF0SmbjXPhss3dh0rqWt
PQRvALPqsV8o+U3m9ucHgfp2SXfj0DW8O09EHrXqJdHM3yiw4+XLnTu6lNkjwhXa
31FV7Wx+2v7aRTtC9UJGQqdmn0tg/861rDa6nr1wBhn0zaX3wgMVodDe2WgXo/EU
z3JtXn5pHZic58I2JN2CXqI/bxUe2vsBMPbXEQJ83Py+f99BpSc47qL1HFeDKErQ
efiBeaSy1/59b06M3zPlGRr5y40uSo6X9ixROlhFs6xxfa8XGrm8jDwzL0noGiyB
PWZo/WkxWkWpy//RlVeXPj9n8O4GZVYmNLK0zCRHGD98Zkv2Q3Mc1HBt16CrV+uS
qIH6h2UWcoc8QtPLaj+XF3MpZhFo9q1pctqDP7LQKNr4Iq3H4/O8lhwz8sp6kfM9
GAKug8sALaQvXDCg8tUwrzueNRs7lWoNV3d98yIH0pYOkjAdKGGyNmHPLNoyT0n6
IJ3n0HFozNAssL0OXmeSJEpws+kKzxUryqYS3hGMyDcdqJeHTPxJR3kec40iS0Mp
DvGd5CT5yC5UPQ+TEKCMCf9LItqeZ8BJf2acmcrtPgpnIyy7yk1lEx6aJpqi9Kq1
57QpU73w6KyzK0iss+UHRa7rTd7xidKsHiDPvmQNM8VFTjtJrtdf+GsYBDBfwp3h
83rV+aTMcSA/medIAAC3eS/d+ZBd6qvE0ejQ0UNDv/16K5PALKsNwvpU56RqfsKM
ur5qSPwX6NwT4ICOdP7Yu7Ijuj3PrEKmSRzMmfn34DgH6PoJmv1n1+QpdBKyPxD3
3wpgFcICu1D1BgqwA41Vi4+g1AXZUyG/XbrzvkfepPq5/aSUehsPI3Ect/qeK9IR
Rk2ewjPN8R/I37VDeS9nBLcP37pZs5jZsMC5YgELLBvyXJo+ET3cux6cZisATIsy
cWo6DhJTW3EzSTGph9lqBLu24vUVUx0xERYiGk1mLPNyr0RFkWp7ix9Ha//20pdo
gVtF1gmBRdL/+uIAPsEIsg7b0DMR8UwW0HNznIozW2yxdWCNLzhENYcSBduonzGR
viYn3Ckp/9LLho717osKuKO2XTBcDLDxsNXi/Gn1pLcZzoETG94HuV3XbGV4wYuV
ZB7xFNM5lXUKv6zrGysPffkcEerKKrSCJWFE5Pu1nnJGoE7AcS5RPqu2fsEQPU1+
C9PgOV/99O/e7zO+VjxA7fy24iIFmSHiJRr4JKBT8TcCHlrXrSjcP8T04508dqLh
tBtNcfrVLlXnsMfX5T+g+Oqq8iFak2ehWPOzJFh81pAHgp7GNFxQyb7mUtkyP/mB
CY8sWYbQmooQxkgdy8xcNlvOMVFarJl21wgwY1jWE+9GGW9m08ojCqA6rdzgSk1B
/5FllDrf72R6l5C7deBIlEWvJmFX6JHDjsBGZnn/EwJ9U9/eRWedDTuLIoIGs70a
oBqLGRpaMD03ebLWkQVJyLZ9oI5JogPnCoV5r+woG9g=
`protect END_PROTECTED
