`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ymZS4vjznDz5RFT17/ELylc7HkK67N1agh/fG4wCCUOLEr20b9pD6rHQ2/xkvnF
CHGQpHUZBsNYrEnzlmxorBe9EoOMbvaMIPq4fH3WWol6gKOeQ7zj9m2UHs5/l+e0
o1KrZZxyY3lOg4yHAZERtIiotN986am2XUalgqY9pMKeb13DzldJkAdLZUDfqWYZ
Hrwp14TSFdBnE0UZfSGMctYI1zDBWivXeonajMBtQ79QskzN/HnkyeCAjLox6J5h
IAoc+a17RQRI8mXVUto1l9zcnbelOg+DkXe7gn98OK4DhJiuFvJjlHXHPR3Dg4M8
QpZ3xnpRE+I/dpVCzqJBTKOV2WKHYQymyJmIGIESx8VdYi2c6mgYaJpT2EYKePMe
5O6dfMVGhPwfgPH6dSwjnVIYt+y340QtNJVr1d1B3YJOhXjLY6SSWl1zSiPUNxzZ
Z0OjfmHcEEOeR/gves6pxPA5aN4jw8u4YrXBSsyExliXzb+hq65EMVyJNv7BVZfm
vLcYnP/miecasRqA4VeIAKwrMnTdZ1hS/EzNs0GcO0WzP5iNrHkZt1nBL17XoL3c
TbMlNn+EORzA4DaOBOIq7LDZeA9g67NhJK6OCECp4LWzTfiGA55/rXfO98sls32r
7D1p4Kj/agR9wn7OZ7/VkPnNErMLBVxUNT09H6QxisQ=
`protect END_PROTECTED
