`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8V+4vKVS96AdajwmexAxity7GGE+tcDyPLVOoo1LUe8wh5Fwo2RjBHUraqNT+1cf
5637HUfxwtxGnEn48m5CrqTjZk2GAOUDNaqU1tnhzKCRLnz+C70y7iaAi6yaZ2kJ
ttvTQAOaUFG7ZlW5M8B/WMbdxu/gIHUFxMA7TZPvZ1/XOjtJ7Zn5jrUf52kAMLCs
mK1pNhPlyGeqw9UPailVNaFBfH4pmBYO/21a/U9dl1S2DWOGxKb/kUjXFDlgL9J3
hGBIVLuBGiWpBuRjTspuew==
`protect END_PROTECTED
