`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hk7aRampVwZ17yu5uDXVZgHvj10c4GhaDcHcyTdodyKCRyn3Ng/eYMiBMN7ew5d5
huBd9ojos0JPHrWYvGTExzNazDqkViYgD2g76TRW70EYvOs3D8M9goR4knPJQort
Q5Bhrkocu0fIi5u7HvM2ifXhma+n6b/QioySzMy8GmhmRUFIRWLcLhSg8Nq6Ifws
y9po9436GpGs2AJHxqy8srb39e3DV31P36QQnRfcs2UdjjnCXNp7WNx/I/s2tvNJ
kULu4vP/EM1q8QiyWtBhynC7NY1TdA5+DT4OJb0oLLEJhE+e0YQR3AO/jY9xhuhO
ifA5QlcPf06tVjakDBzh1+EAiC+6PN/ckS3IH5diyjhth9L9sEgsbalAegXLCiiE
msvCXpdJqJqEhtdK1KSJxw2JV+uvQDoG3Po/59/CuubOvlKlDtPw1FCk7cHmAO+C
Jtm3SlXQaElvc865RnYIV0L5sHtGJGnbfzve5D0sFAaoOOatej49SRe8qhNkiz/t
YAGuoTnNXB9PnWL3QarinGCg9QcSjbrnB2pZiN4Aib9l8GdhD0FLJ4b2iKSVBGxd
QsTAIdq8bzcYzpzX3chhNbamBoj6Q5d03ScWnVC+Ke0pt+X6dKeCBHV4cn4G3RLz
yky2bci54WCbS1T7Fi3FS0sUNqkE9pKzxkPfv6eY46jZff0spdEKQO6Qi4YJJ15T
1WiXNDGYLqjGs9Wt8VcDrjQiTsUDESZmqWpdpuZYOx5HFygQCF7vdt9KPjWmdz3g
X5zsRDGcMSKAo1nfOCBAQ+GKp1nhhso+vGMVS67oRcXPKOdPKPxt3sJsXj1wsnAu
+G74hJsYKzXfN1RH1XvswiTcpD8+60VMbs4StRTaqe7OhkXfHGxAaHVR6wowNkdy
3ATNQsEAmRv//8BLudQg6yYq4ZE6jp/9YeWwasfp0Wf3F2uEvhywLdF8wHEw3GOU
/D5igt8PyNzBpxVbDfVal8QUOX9UMNont0DkPclwCnUFMiKR7MCTjLYr4lSB2OU1
tpMTvnYbfdy6YmL9w5qKFLz9vArGH/VJnXr41zQ2nx6C2imOf15V5wpyFwD8cXD+
Zv8pf/5e/n1Fva85OvNaJHN4j11stRiQRZFPBqQqLNaiYNXrTstmRjm2+3kCZxUP
tue7X7n+SCoXMxOwgRfHBGMhYNajcvxOLP8Ee4FkYwZ2eo+ujIokAQH7VcfrLQtT
gspfsPaQi7owE1HLy3sCnjYHborpHUfZufnVZPX+p0NlvjCoJJZLOGKJAGa51aHX
MIIwPrqQshrMLWjW8gbzAka1+6QiQNXovrQCNHhWyBCQeNDbykD1TRaMAs89oM7p
UJFHX2vs6lfbOMNBmenYToSGLgH9q/U93LwFMYHr3LY/dHDx56w4nPMiflJB7SBW
UIs5W5ze8MN+wJ8xePjFoPLaK4hVYHohCpz8SJNWIih/5GIJZqT/oDa4HZeGtcfK
GRZiBdDXSm9lWg/92A02fOUYRDAcbrY6wRT5HoNIX6JiAOSSi3tYBrKd2ghEju39
DWWqB0+K8BzmxJVj2zKpnBuow4AlnmqKMA0rQ/2fPy2nSo7o11nyLwfuaAQH7aQU
5Ne+YFzMg4/q2/Ho7VwGYqlad9Fpnry07z+TtS6pRkgKMRKhrKr9WkJoqVvKzsJr
OygEGggQ/QcgKTlyYl4lVzKDsvQXtB4dtN29vgQ/+wcxMZwCFuXDd6jI5JK101bW
hD/VJpmQt66f5V5N47eTn6b+I1CjvK6FHQjY/v+g+aBj/jIFIYwpnHhU9dmrV4KE
ULW2egVLt+cWcxgsW0vtpqGMS78XlFteEKjYHmyDOY1LlaCJkTELTDhOtemMF8+A
7j+EgE8Mcn7EezYe7I9VmBekNzGqg8Ute61ENO4NtMiKjGazp6UEpbzNPoeFNppV
EMapDVIAQk1Xq+dGwvI6QelX4vqb10zR9dI4jtLStVv9RdN+Cq0CnM3ClFTD1LqF
IOYSoVhT+b/fCAa6fOpkRTz7f2PBvQChXlz2u8HYdrDlK/CM0DwKe6S+PI6Cld8Z
vjTiAh+RF4LICY/lC/0tnopgpbqhWQUIrgLrBCbN7Rl0AH6i1zZSWJrSFBV7zH8o
VthvsN/BVXbOM/8NUhUA8OZbW90Rs5rHue8j7m3OO/qI+rZrVp/aRDusCz+cCO00
mGWHdXS8jBhBPJv9MziRqbqZPJ2Gd3WlwaIa2DP1T64Duah+MLEayF6SQX1Z2Fba
k8ww2rCSkxnJGy8SooRs9fMX6Dz1l8da+n0aez+jH6B+gEYRrry7AjShYqyT3nAB
bYoDNgOPRTZwp2kHBxMVOKIGm3FpHaznRN0m4e3f7OyNoOTBDWhLCCc2eoRrG9xh
EEUbdeFJQKT+hKZYhvUMTdTpLg5aO5gjt2mbEohmqr+EMLEVPh42T/kxvBN2goHJ
JB8WdpIiF/H/SrmBp97daOEoXrvT/o0IVYGN0D5hJLRJpE7OvmYk41ejxbPlgl2a
Unof53ood6FOJTbhRIMkDzSsHQihCyRLDm/Vr5tXkXC2jP4HOOVGIjx0oe4K7YGS
5Y+iEcgpQXgiTwpt6dfK5kNyqzG6oFeqoq31oX0G6csJHTYQJgEjQryR4qAAVcgO
Hk6HwYa4vO9L8G6LwbilonLFZS0OpSVQ2H6k1SSRC3JU2z+QVmmNq9A1T3FrPkcp
M6LgcRPll5Zs6GjkZwDP/ADkOWAOV41o50GoAGQEeCknB81LEFaEZ1D3L/eiLoIz
2x35u7ZhD/FBYk/hi7Cu8oXdBlpckrZFhC9cID9AFiL5W58ZHVTdkswExMeAlDZn
ioANGoAXfFqA6tUReJmvc7sa2nTaS0pcUQEKqsqExqrXid6EyZHw9YPxURtAfnQu
95RjRDEnuRM3tJ9h1zwyH4QWDGm0kZWZJ5dZ9XHtvxe9otAtOgu7dZXEp2eHYgj2
eJOPtAWMbnH3ZYMTsFn2EtueBT+S4dSgPPJ7FqBkm/yXBw3X5N7XVku1RV1uqaPy
qjylzJaeQgZgULr6jr7/W8aJY9mhw0XAfyIsK9tH2W4+IzbxAX+DqBrGjAtqj8uz
JzCk+mAQ+mWd5HlzkzUuFrRNbQZZcuzBsJh905ll1PLnsVXcXhaXCd/Ni5dusGbb
4UMhMD89A9VejeSQFSV2+k9KRe9CX7j/o40F2EWSn7JRsYGkZe7nHBlkBArRvmss
5Cmi9c1rzMkxFK0kQwJ/JKQ5MD7jaMKqjBHw8Dg096awc2YgXufSVyqqV00v++Xq
mpW+gF0Vx1yQ+ysb6MygX59Sv8VnpjxNE1eVEly0b8AGMEciQJi5w3DoerVO7pmn
sI66lILXWPlrYXRVXnCTArTnzI1VQMWAyf28NxBgSFawo7hCZ6RzSZ+WZQZxAE4g
N39jb3gmJp3yTp1nZR55ChiEm/c7KgMR0P5atv41jNQ/DjuZxm75FunDTFrmh5S2
XWwnNAMzDY7Nl79Pe4lxKCOlqZ/gHXv/hJ1LjSQ7/hqmoY6CvtvgmHw4rSg+QSi6
0Okh5u6Iz57iE8l6tIbqLoO/MVolxk5FCoiIqe/OzHgTOEZ4MHN+uACQujyrcGho
fSjWsBBDEpZsWnXPneAIwIYJL8d3VmnSTH+l5yzREeoNLeBMtN/bWC1VBMBi17F6
NR5N7VhFMdkeSdZS7OueT2G7SgkBq08xjbtFlJWzYxaM8b9k3LmpMh0Tp1m3YmNS
uCj/ySOb5t8fV2vmyVgicfCxLyF+kkHyAZrdDFCXt3EZSVBQ/SEZEoDO36/bCpGH
3v/2lIfaz1ccOPtJE9zKpw==
`protect END_PROTECTED
