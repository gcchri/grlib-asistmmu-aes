`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VpsTmTfnFIHVF7nqxkiN6SJES4fJV4ZHF98LzX6viAtWIyAbI2HmWvNw6q5wwEd2
kVYGRFGFWQWKra3/NlOECGdpMWNEQXYQbn74ze9r2CgSS+fYELY3PE1ZQjcxW3zs
0ibqWA9ILQTo3wCZQg9IL2dg80AuAqEuoVTtFoje4P8yDd0BpO6q5tiMkMVQBWtv
nYwTHvgeGvsL1z8bOXBcubtL1AQzs6rzrf6DIy2e9r9Vp66CSXsPV94h+5KvB0RV
8kVpKcrXIBwX/aUYb42lxv+aqf9UphG0KCP8/wo4pdXz5F2ktzZR3Z4iMt6anbMP
gCXoryZQPlZ8zV/eF2k97LueIlNODquKy5rJVLBbPtf7PMTEN3OC6YSFbCozMe7F
qfxrKMHEYfDy8NTvJn/YCUgxr4AhwHz/CpmTPhmFnIYpKmCzhl+JjA7XWqyVg677
G6k4TsfLcvfQeRHqVZxQZm8b85bOD39k6MLc9f6h6+HENdDGHzAtB8KqXgCeGpZe
rkx2STjrQucF50QwzLrnMaEs7c2eDQ7DjW46VqqeaWczV0kuJXF1EDF3FEJsztWY
vU+w1FnlhuXBysGNqV36DYQBhRL8l+LD8hBW6n849hP356yLg5YAERbummb1kumD
tikqs6PqzWmN9u2WnKMB5H27oHafn/EITS7B6+L1H4Y+T3e2W5z5K/JG/dMThPUF
8DVwkc3vW56mTaXcSL0p6jZU6MB3VTEFj1XONkIbGfdpWuIUWtiP2mTvZ0rHhzt0
acBVSyNse1uYChnV3fgl2oWSF0Rf3U+Kc6RKAQObeMJNA2qQ6h5plghGEUO9Yn8W
7zoFLriI00YnkJhNYKPH9Q==
`protect END_PROTECTED
