`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G0T0oFtd8xrmanEfXd9ButGDxDhq73N5mp8T7nfsR222XGw6tcOHyFOxUuiNHcJf
pdOC27l6iedoA/eLhY8GGtxzTjY0cQ5/clVgCrCjAFl0URieUWdwY9Lkarz0m4RS
v0nyOcc/GwLsGg4hP6tqKpyqHVpLJSVORXR0GIQNANpgojs+TYcgk4PGXn4cPvAQ
Q1elN8MZsw8YZsLvmqVNdKxRHwlGBNR70LwVaV1WUzc5gRkvu9kuNiFln+7z+eWi
5AyDWjDnkWADjqPAOqgiE5WM52rxfN5ZSGExISjG3BqEY/rFQ3mwgr4D74WKsxWe
7B+hUwsLfk94ecPX7e3hkKbRoCIb5ClPmBN4OSySJ7WyT81WLkrYuOMqFVU2Q6wf
14dW85v/Ipkmqi+S+3dd///3obRMeLrEgYUKdz2BLeXFa4T7KAz6Y8XTOxwZ5sD1
lk7dZZ4cQkdIWKcqX1o0On1mAH7ZXucvtGd8BITX366/y8okc1T1wwkqNeR98C8M
Yl63GJ1nVWAXyBWT8C0ZhKOM6BtVB0ldAdvbtVMx30NnYLW3xFaCAW6sMWo2buR5
woVoNCCVP6L5vXeyuNGN6kXkDgcEOCHQwB1K54WiCqaQK5URxSLDJiwYDdy3pikq
8TLUEBj8Lzxz24Hx4NQkYg+87waaN73mOr0H8J6YaXddLnjCKMdyH6jbPkjExgKQ
xw8frZ+CssgMFMPvN4aZPDdM5g3e70bUBCSJfBmwEXH0ApT5znsbngVG4r/NzRgY
tW6hXr/n0hFItRZ2p5PiXFMT8y4bo96eIsZ+LkgbsgRH02dXuEpVMeLUdG9lEyw+
do5pr1zqgolgTlvWhtx+wEniV8cy3HetRroYWgYLPqB0EJO3tEXx8cFRVBH8JZ/o
vEsXi+OeBWcXx1f1ON+s1sRLXiEatdmxzrk8jnTZu85pqIvre/zNPm82hx4O2Xlq
yuiUdtSA9nKwYgYsQm4+GUuvfXH+1ifHAXqlLt6M6HRFu64g5+gKd7Hq0ifAwGLo
xR3j0azq0SjvcY56kF6XQRyayC+vqTlUeHhUrFxCyCm1oFaWtlJL16swLqEayoVK
yLxNLMEUQreB/DVOb7szl1w4WWx7fjRNU3plDeRs4jPNd4CUIgWExRJ9xU9FWuYX
jBT1ajwYqTtuYAEIm+9lYV8sJi8Oi0z0YI6ETnYoJM5HxJGYdmc1oCptQ5/INw+t
LyrAL7G8aHVVm1eZvmvTxxa8yHGhUX1A5yrLpmV17RUghty/BXJq+c24yaVEyFw3
6K+/QbmXz5LjyxuFgu5MolvQPD3u81+gZavuvPCMhTELClM11VSS6Z5B0qaIb92+
tF5HtKMWXaKAhGh8xUiOCrJZXplDnXqSI7F0B+UK3sDAWjmKquCm3vIVI/TxB4T9
JcHWD77dojS6WaskFzvaPJ605mMvFW2TDrwCaXdy508=
`protect END_PROTECTED
