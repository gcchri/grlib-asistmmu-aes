`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wVS6FXmoCSTJW2Zsbi/IWr/xwjznIjcCBAfa+6lYu2Wp4q06/gzYNf4I6sMAUxJa
uyfQSFPKOgfXqRHaZzdbnyjnusjdPgqcpy9soZGQqXP3YiSP9xBRiuGOplTKvDgA
6CdqADRsQ8kSE/vzwsMSKNZ3GsnD28XZu/BT+IyYUjNwhyta61Pnuug+RAnfvT8V
RMsKn+6+oskUiL40AU4NhvUlfh3o93tJ1Plltgj7smZe4Bw3EdK7BvoqU8tWkYCW
9ZKgqFhIRdPRlADqXbDhel1Q4qb3/e5K+kMLKrH6FRg1jlWZHiXHpFJibLbmNGT3
9UWpiFX7hw1FSrmbmany7vis4E50sTvPvxgTCiGYPsqme6G0ViC7H+D6rV4vNb3g
1FNnW2mWuJb23wzwA31tjcT+0lD8lHYHgk+uqdBtOtGAiwni842Y8DMyPpSIZyX6
LGgfchqhJoez5iDFV5xx41AWHgrLVE+bIEoezB9ejAfCA1fR632Stz8eR1UnZJX7
lpdl0bDEhLrpzNWdJEJ23gQmz6XpIPNz7YipMM37Q3zrkzE5ZECKN9ZQSwtmpDl8
HBhvYpsOgMXhK8JQYvtk3dv58aDAz7TzPNplK2Ril9Q5KFO8t6IXhXFELzLKIOsG
qHmhSA1QDFQioFZtp6/5LX6csW2jDhNDpDZUPR/SC3q8vMZGlY2FlqrsG8jb1p8x
6W3h/FDJK0+0zrmpHcHdqJuzG6p+2ZYzN6/h2JHQTiyYd2WVJWgF7XU3DcLDPWT2
howOahpJFFwHdi843Ls8GzW+ZMSptHIz4WdZGTfi2BIRPInsJFziPtDgLxQcntMT
Xa3JT3BIs3HcTS0zjExAYw9igjPL8STIfM9aB3y0FWkkJniMHUA89sREogJvPjxf
EkJ7Wd6gWAlI1TqE3bCkU4kpEjVWtueZ1yRT5SgGiPGsAZ7vD8Uvwwzu57vyvJCa
pNb0rJizdasKT3DjIhQwQydykhaHAK1j1v89ElUc2sAkuHczxLOcZXU1Gst9rqF/
Ijyg+pQn1W/cs5qZEB6OdTvaevKMw1y1hyGKc78R2z/GqspzMQVm8pWYd1q9YLYf
9pYCVjPHOXVQR/t2HgG5FVQLlkh5S2y3D2fEFVtaV4xzrhPtKBSUHNks+WvSk8yf
C6ycg9IXLNyjSG+q/Tzeftd9WXioI/dg8/emZbGbRM7LJAY0IlQMMAoT1rog0w4X
nuRy+ROwwdjQbc0uOX2tlFdlQkbu4WZZEpgyRnss+6NugITqzq+5GVvZwgmLXjg4
qroC4PBKkzSnCWvp7GIfyM3Cy4c9bO+Q2U3gxOEUsHdEKiPKr+qLVFMeIOj+bixc
6rfxhglKCX4ncp/TnVhrkuALuNNCbdeUVAJbA65tIAsSxSPFqp9ixjwO3yICYgSG
bxwTzNaLW9LoNCSgqooy7c4YCNuVj8Y5IoTUfFkCpMmOxuO+aVDkrICBRaxo6a5R
oYP2/VdCFK0E6j/J3A/E6r+UhCkVb30ebkVm63X66qjJLZBr8niHyLtzwwtJQ5OC
sBDtF++oTE/dMRI3U02I4eSQbLOGjokn06aSA6bniUivgj1Ktb7WGCoWyWksmRHi
`protect END_PROTECTED
