`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jHJxx7lafAsZmG26kbrjYhNEzkgERq/cTOA7gJ5s4iOsS5hp+b9TMLpnjFcCl10G
JKogjKvt4Eorwr9GA42fkuFz/aXbKDQ/e6wyrE/Pzz5BN/NJLpBqtOoY/hbNfNy7
fIwd6J03Q6UGCWPj6It8gxD/ZgxxQPopUfVbpIRsWNnxcTMfWduTdXHZW4u9fv7l
UJBdKMa6y449aghbDmyHDADzNRQ/co6XPo0fq4SIXOSzyAw/ODJOW9CvKLFVKLUD
dagRQl4NDgWMyge/9S18O2lPA/JqM2lXL5BNouSup2qmC6K2S+6Owp/hXx6qWZFb
tkaFN9aOWN6VDZKmm2adBW14W0qR+ypgWbmxuW13Y9i8/w8GpzqNpaw3dRNeJVPA
4SsTDCCSmlSDyucbyhyqTxND20Zl9km9PSGqa5MH3vA5hOGojHi+WptMcfp1ZklG
/MtuudaFSb5p5zfGT2noKdpI913leK+mWIX30bfKrEPEA8aZLiY0pDPlSQDwKJUc
aDIWN0MdysyqGTMxCYcHJ1mZmYp0SPRTAVuXwN1iGr+Xk2mtwamMDI+ENE7p8RFZ
COk98yz+yYY5CeermKTPMh6nAqDYCfqN5HbqW4/Be1dQHCnyt1YC+3qlHbY6is98
3hvvnY4PGt7+bhyDps3d4Sw46TKJr4lKOSqt0+IzInyr7G+B4CErB+85VPa5tIP7
lT+iM8TERQySchCtpJneDzmTuRtdo/2vYSQ3lTbdmL7NQfjjZ8TD/T9k7PU/vccm
vW23GF5M/qz8HdqflXbKSqm5XzNTTdB1MnKTkj4Trb5YNef54Kkoa+DMT1FCH+1n
wVBvhcSCMv/12G8tQdYouw==
`protect END_PROTECTED
