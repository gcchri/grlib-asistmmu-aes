`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q1p1RoAjrgVt0JIw4lJrkO2ArkYQKHuu394uIhF99esvpbXsPTPXLLYluPLLXQbU
fuXkBwPN4xATrLidvgLbEZjwjKLd/UDvc2XGL84uWLxzKkk+fvz8iARrD8qiljpD
LiMrz1EmWNiKVwRTvm7EY9JcANRYc0oxVyFNhaPwFjQklMC2xLxhIlOEEpVg06kR
TxBkXiQ/w00eR6nuOdcu06MvCyeAVEb88+ST8BH0T5fKv+ioqWslc/dawoRlFm+r
Jac48ytStj8eDBnWfGHCC1zMlOeF4CtkmmHhftucApXV2mVuqqP02Kxvdqkd9zlQ
DRodHAgQ1wioy6TytBhLQnAgaDeEE4M5VC5Xy7hopKToO3oDuhyEYG1CWO1Sl1Ev
6ysQf7U2RuKgNgpUYXVZhbNeWI3LTu4dwwVCbhRGcicYHMNBvtBcz87ssKhlOVkK
77QhBtU5jhVFriQrBu8HDwRspt52DR/eAyJMGYUy1g3gYxKUhp2khciopaIC1rzy
/fV/Yz90rA4EQy166Ku8fApfLQzrafb4cljcOrk/zBKIUKE51jSyFSN9oOClGjXS
4GxtBuUCjed9Adg9spqtF6D38nZoM9mpkrJDSTUnX7xfzsGYjO89Fx3lXgvCRaZQ
KsUr/m0gQ2tt11HuS3BAmERapc+2spAohD+JpSQyM//UGMSjgbEHGGPuy3KMMHA6
HooFs9v+8P46YCp4m8PpFr4HoVZuzEKV2w/3pRbnRjJ1DHZRj6jerxW/rbInmevF
xhDQTnE+klqgD0Bqc5YfzAGeaoMgbL/NnpYEcHVL4SvwdeOGRk/4csjg0hOrqInu
Uwv1xIqnKcdJMYDxSJiV2GFVmgPNuMwPNdLRHuJ2ltCAgn5KtiDHHN05ARKdfhbX
QsuR+rD6mQa9mzCmmgAoFFBo74Hy2NkmJMPv8W8ZMEPkhtIomPkYwIBda7g3145i
lgEftKMfxwyO38AIU3T1CsQ8ggUWvTJ8K3kfr0uIDGZWCqHZv72kpYa6VZx3Pzkz
T3TfmRNJcf1UPEYBgPUtHu4TzzsyeFQAuDx7FTnL35k8tuabkomsmCUcW8fRWwSh
I0Y+E0wQB6XpMg/ATPeIEC6ZVILPWeqZCfkBZWI+f7p3EAjLQ4T6KjTSDJOtSrMi
axPPjOFrVsYH2TCfBSyJGcoUVhSLy20yIlg+OA+MTRlgP6hU6llO49oURiqE8KPv
OAPORE8JEc5eADIWojxmXkwIAil39iLV7BzssJwkDKYBgyNRo9XsmLjwwWwM8qYm
k1bjnYJ87VLhgnp3aByxOtaVGGUjM3fkD+e9WtBX/z70fBO/ycM/vrlJde3EJQIz
0kI54QSt+fmHMuHwzBF5ZR+dWj2lcKpykIYQ1ZMz7VzdvfeYuoq6lkTVtQUHpq1k
SWLUXilwJ6D8prc2wck/TnKJganCm/WLQlm9EHB4ApmcB4r89mFRljrDiPB37kbP
S2gWyJEF2eA+t/s21bX6OqIxl4a/6AUgZwTHvqywS2Vfgu8+yAP4cwajOViajnsu
otBnx26t7WyEw2ALZ3weGw5Kltqth4IufDTRarlmv2nV1nyG8ODzdLiRPjAChf7o
FwynTygoMf1kVB84wPVSDZSQwq0ruB7MkTmI3ZiEeIN9sXNmmV6K/jdomVzLWuGa
6ZzRnHwqGE8DMuDIUrOxTjy71vYDzOR9XT8lbJS2oVTrZ++RdBRiBTeU5Ufu8iwC
ApNnfy5EcILZKZkpPk2PtqnlWeDpNsG2Oap5aeqzcOzfnhk7oL8yJBMXz5aF1TVB
cqBMdbPZchpLBfo01Vmenek7J56FY+sitZwu0mvsKl7AAb3sz+DnNShkpmTAKf6Z
01U7tKV+EMQqii+eSD3SLDnkoC3lCVJAL25+KN+/f4sUbirS8u2NlEORgDDo24Wp
Ix1XOUkVgsi42fE/ziwGJ9JXPSplDVZ5DsxU0FINHB7osRJ/nJ8T+5rUcfl/PGdJ
hpxt+4xaTXEE5iGY/BuvgtLkUIWP/i6d56XOMX7JeHBxurgaz/HDFPP7Pt5NezRC
ctNzMCBfuHvIpObCTYpgrbftiak+7IaqBe3c0CNZFlBm87gGr5FPk02rilsFoxld
Dj57m7AfnOjP6HK4nywufuUKKSL8XYhUgjh2w8A129ClcdrWeMR+BoFhhAjNPvvb
SYz+aWwZ3Kdhhfx8GJHD/W3ey3ylPDoB2trVZso0X0+Lx+HAWUwoztvYrSH6Om4f
QySuXHvWpS+iiB8vhONT9ZK0ksKTDC2wJapSikP8euEYO1nJ7tp+H/bYl48p6NSJ
SpouMKoMDg2lMdp/Ms9Nr7HGRTmw5PrZ0i3xYm2siPPlPEkxXqfYSHWXxw6TSf1S
KSajMfBvY/1YU0KizmXJMm35MF65D/E0xiqUklrFdgmr1X/tFvU5Xjbsl/cl4QQB
BGkbsXaH6aUhxuYG9MltmBuw4k9EyE4Bm6HNszRIWpUFiYSdaUtA5ASvGakjKc30
Hp7R0anLbuXyoGbUHRx8frPnHNcA5mUsK7C0/iaIEgVI/74nuN3kCCW0joonhJo5
4EJ8ItM5jWht7Y3XT/oQTvx52CJ8FpQEUnOhW+2ZCIeKeVyiKcyQg8Io3riEJ57s
f+52lFSYUCbpEi4+yenYVajIyrkkzlTtYIDNyD8ecpk=
`protect END_PROTECTED
