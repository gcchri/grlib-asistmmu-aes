`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GgTBK5t5M/PF/bE2Mw7LAOaCvaJJX97XU/RVkn7y6tmFr44kNviazOBMUA5iFJ5E
iknp/C12bOxBUMp30o3oQ1FWVoRcprcwNSoI27n/zwngy3h/p9ORfrkhZtYXyb/d
vUOpv0KWBwU038UAC2dTDaM3oZj8L5EqPP/NHZHRTWArX/U0djztD0+O75KPcubF
HtJhv0Ps/tGhugb1Gu6Lvw/+qnaWeqvzhksvK5Jowl9bfk/zJiYd/XSyl/PDdNJy
2TgO1aAM0ZbRojcRBbRKyp6BKOvfvhVbH5YFYFGq9lf2TmvuCvc4WdYKun7s1h6J
b2ir/w8POqOa+VgEueX05vznFaKFJapXoWj9M0PUqBLMNVaKsoQfsfaHnISxu5HI
lOzJCxc1o9VTAhWRs2mhbtkCTWfUSfAN0NDSw4LQ0XMpqTEaOzrJOqvTTh1j2S7n
i1X8kxCf4vWEKhlGcdLEAJ0hPirBljz71z271xFS3uTL2j+S0yU8cIedH2t/V/5v
TsdjrnDt+2j7kJgBBLr/sdTMG85tpAlh0k57NmZlQASw6Dq/7mSti8mYu0FFXji8
UA3/x1uJwMtGkNJTS9aS751ekWd4Ll9NSiL9TrVV0TEi4bQ4S5y5CmwtHwsnzXdY
5Fqg0QcjsBsllTMXg8F22Ki0nCcojKTUFKIrHJLSIBY=
`protect END_PROTECTED
