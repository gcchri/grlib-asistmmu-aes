`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LqarupFT3vuoXhYhtKFU4Aw3zxIX0JaIU0YjeAnMzh7kfnq9jI4COGEONr70qJW4
daxTwKU5Pq1D7Apb/fLoBBoU77kIn8Fb0ZrcA+y2Jq9EdKftzmP4RV57SjIU5EB0
QTvWVVROLlxT3WLSkAQpx7kzgANDue4+hvrp95hJ5XNSHA+ulrA690wDZgDnLHpB
yPC7YS3woRNlp4PEb6FM1RZGPVM1k+oNKB3P26K7FrJLm72Y2pu+Hp1lQvJ6NOJ/
darLm9UEsK07/A0urr57FSMir2yt7q+tMyGzJuZLTr6N3klQyaaXAo1swjwQwh+n
XZwRykZkf2pZHNmFzyYOt/CvoHN0m/v1Y+n/jRlO5hsJcqiPoh6uxWfu207kfINo
GGdtFU4X2zEzAfSq09mnxj6pDeCTpj3UaWyKFCpJsZFOrzuwKG2tzMXvyIkJLme6
xXD9syrsJzMNY3KCyNxvOlsoHWbTYsAId6oaNqpSTAR0GwkGsa+ABLfh31RcDhGL
JKlHcPDIeEvHkR5szEMsdqJAEkMz46i7Mg4zpJU+07KRVqlvKgsMYKzeRrX2QCFn
FcUDTAObAWFpnUyq0u3fnPAN/8XajdKfKQFkJ0GQKNmd0x13uqsEZcxlmSWUGq2O
lerhv5OtgzsZf2Xao2oLpNHrjmUcMinQ957TOqWBA+YeYaxXxTkU47FbZXBmDpn1
I2kGuJ4UKhiWXeY15qJ1GC1OPwlzN2qPcVzgRsmfof4kEcuORTJ0G3v/jFJfzPSB
ipMeEv6zPcpeu+bFVqcH61lj4hm6qOgUo3XpUJ2fEb8B0hjeChbrHxdI2aQK7RjN
xWydBbeVQUAs1xB4no1FT1NQRIfI6hXVWsdWMyR1eMaWQvDiS7UFFxJcuKNUgSFr
08wmS1kCZ7/gpRVmxn8JHLeuDY6biIbjhTjshOE9Zl93rIDqf7m7fLPEtJ//Y2bo
j5Z8Q2KMj0iEplQD0n6T9WQfAoMc7vv7lzOjCru+OmLSxsDVXKoGlX4O/srnAJ6H
kYIc5FsnMgddaK8V4imHtqxVIw26t7XX/LBG3NIy6tBzRZtcdr3q1lKig452jN+d
HVtI2bKEx0uraiLKaLrMXs2bzp5/UoDW0CEjs1mX3qhSy9JuMck3R5y07fNO+hwq
tqZ8F6iiWfhHyIzCQ75BZhi1XBibjQou4PbtBChZLvtQ9EGBuwjd06V21aU178+P
cDnz8pumjW9ixMPV2b40H4j01JWZKXeq1SuAXKiCidFrBzxSYarqXTM82FQkjHQH
Lw1g0XmEVcmgFH8DZnlaWGpJ6r9MjZ/MzA/UFEiYt6T6oK2CUB3UlwYmTpuCOfAo
uyumfBVOZWb8xJ6BMTuupmXmy5pRPK/JjaMY9Tb9zwTGeYacRIRgnpO6+tc4n8mH
rH1SQ4GBsxUq30vbHM/fztaLh00Sow6/8td9IXI+nIjXhEyYN3XNi3/oDTFGa/tF
2ZHAkuMMUhonodpbpDwjOnU2OmpY2dw7tIEaMF6WFkhvtbRL+XXm3E45K/Eh83Ed
MS/9eVbDQLJsw6OgGKQMxqn2Ojmp2+2TxHP+06VMR8PpehxeizzDZsgnNyXhPsUI
5ioxH2l7mGYXrjQ/AGO2DzN8oRAUGnI+ViBTGp+/4mNFXVOpU07ta+q/12Qq3WDR
xu079P2SJaiw1Z6NlJzkjE5eHALJE8J3QaMkNcDwHquYqMfUA5kBNuBMgZnxpiWH
2y6kRfrmQeh0Vl3UetKU7R3ebCVvC3m0GKApgymL9hTI9z1z2Q6aINcvQYIoI/R3
F1QDof57VEJal4zNM0dzHUdy4U8qNxX6N37weypTn8dpXdxDMKCAiE980hyptMY9
tdkDWUdoXCrSTPqLncPN5m3+bYgQJhRixGTg8xcaHMFAGd1b+VbgSJAjYnATsMPT
69VA9ZGb2uxvsrAEnsIjS4Mr9NC4immfpBerk3x3RSbfmQnWX8/d5ubG4IAb+Mv3
yskS80yPvBxdmYSUanNYBoDNr9QE3b7xHzudf+TFtTO1/DjJKGQ+8UGpkFb8iyLj
qTLGVai87wN3l9nU9wzucqwo44iKhBHMZBlsBr7Bg0/tfEpZ2WNWdtyAsbO1U3BR
6H1Uw9klZziYsIA0kAMj/DPj3/ZUVkofTASlh14eJ7jSf974MI7GdEB7IYxRPvPk
NpMS5rZcIwS/7VoEkdlMgYcciII2d70ImEJYvbo7g088iuqI3JtLYbSHeNvfyLY+
W7pPWzSwchRWuLcFAr6tPpV0B6W8dONlvkMGI1lMu5Kc7oJt8UBc4Z0AXxO4Y+c8
y74hY+vE11eE1gAYZTvePwWUVwfSK7HhWRyzLJgqu+Ceq6trGkeq5qcRUEq05Op/
r4mHHjL5bh4PQwNVmgbOAfa+reNYKjiOXAg6gpPgpWwN/UEwY8LkJvQRS9614r2T
5DaJwIYXzOoQaWQaVOKb73lF4mF3HaolXvM66Y/smWb8hU4Pz8tvOPQpipU+e74q
FJknDYuGpwTcKKk0V3+gylDVKHjAh/N6GLybVRanr+ZdviBeZ/W6jTXjjLArDKze
Vzn3qS13rys/iynUc4hkve+KrwcnQ4WfEUmcj0HkvbBcoRyxnERnZh1mIAq6uX20
iFM3+rnvOjS4d9dhXjUGlRglswiTrgc/+OxeKcBfGr2QWo5sIFKo2+r2Y7ba9K8V
Jpz2PoThd6HW2P8iNHeiy0lf8mNS4MqbeJctqfcWodt0wfqz3wSSWuV2/exDWLUu
2oiHX1YbZhpAmx92S/qUUAnMdgtWEi4CkUSR9BxvyfDOdyZITTOPqqQgvOHAqRYx
we2W520DrYqRbaDf2v1EEKgw28R8iy+lHIq7LV1jaZt4LaiJ//m1dC+9sUY0OjPv
FPHIPV2v9ffpEInQcJ9GUoSMAcJnm/5EI9cODFhdlLRwrEa/EQ1z2NmFnvQfgF0u
JrSKzkM2WFeYAERX0OCYVOj/xbvwUDVcxotdDEtg07eX7boH7b2wCdp5B2KEqAlU
j0iHmdt30ZGoNCM8BLP5jQ2Gq1T3BVAjkocHkqdiXQVrMmYBxhU25uMcsahPu/rn
jUKaCie+TAUMbW5DrA+TTJNkF3JWossUA/t1Kq1mXQHyq6yYk0yY5/cJmf77mcEn
8vk73a3eF2oNr72u1TTR0GDKPQihbgv4X2HK3WUlWqNoyHBKs3kPZP/YCHZ3n0lR
2jDt0NLvIi/28WDnOqElCnM+E1v1j2zfrO4/ozhv/iTzj2ipSvG3P6Xo2WSXMjps
YGLj6Qf82BqrOiiVcaOeb7wCjRMSB/bYPgs/dlAEXbiCtnaOcQOgQiCJt6fRDAqz
RCF4TdyVcy8Hdi5V1wtjARjJw6Lt4Ydg1hc4usuGMmVcJqTuwvGj/LY7FB+5qvKE
/aKAMKvM/j1VGOWCCzYk0iNiG2kJz9mXcFrXaUuQn6xhfRk5YevxN3FDuhxoUH7n
PS6Oq6FFh4d33Nv8xqXr10B6PhDu4TgecKZSu9fiVw6MBAMgevoX+xpRr2DaYP92
fM2FZg8bkcZBZSt2pWZS4wbcYLwePf/EbM5a325iqmoZRzlQM1tK9225PR6AAJEU
k/a8ZsIAKjBt9Ht1DQcyFZ9fGOmZ6z/lNVM8ZD/Wdfy2HQQkNLJt4uQwzs1IEij8
8Q5FyptU5bG3kVAaLfP88kTbYF3bAypcA6S8GBIJ9TYA1pm3EQdSdvhV563Uxz22
SR9tkyqn13lIWUV300if36DhKYD6svKFDPmRd57a3ibLCN6aO3QUbwzN+T/KusQu
LG3Nfo4uOJtyod9oZV2xrUxeJFagt9t5vOGjAORC0gatCIz15YGWoWdfa/TkdNmQ
vzy9CRQT+IuJOKr1k/BOP1QemSP9t39BTHMNQXCmOGpL8rxz0ycV4qP9PLKh53/C
1zB7xypuQ3mh9ACPTdZPDxE9jchGap9ZGlTHXSplpmlZocUiW5JOwaX6BntDn/w6
hzon9Xnt1wtSyPcdycivREKFbfAhe5HdFCZX03VoM0H5DspryE138Wab+OhQMF0w
A1YZNmWW2tVc/rTOb7qDoxz3r81T6hAP6bvPbp5iVERwAZIqQNqpDiCbXC9twhi/
UdGReNoVTeLigaZFXcQ6FsD8BAvKW4mtIWZ4i30Qc9iAdRQwlUuqwX/FT8SEVZE1
8JcbgaksLPRPhCX4Znk52J7/ijZ1xlktKF7JweVgPu8eayfJN2pjJIorX+2C675u
LHe9vYRKcAhSelj1K9geGMguEM8c5qECTHHGIPcqvY0+vG2XQnllhEy9OFF3rb+f
yMttS8yuHRaAbwwzVrlRVg+xKlaIuqrOqJtj86j7HfJavXlNqHEy2BgFaA/xlY++
1R3x76gFsU0O20oYhCwH4M/Ztft2NZta+6plmn+c4v98L0eQPQaagMvJp6iwcvsr
Jh8bG9D42EqtRWK6RdrMNeYm+YANy0w2Yq1fpVwj2AICVYOPMczkc+C4n5UFLIIL
MWfKVSn05yBxxZlYu6CgBhqcXBJKZ+qEXlrFJxhHqI06GgN1nHY6jnvD7yfcsdds
isrDLd5Fn0fKb4S4aADmWCVwIwWUxGaEz+bP8QmrogXLcf+nTing8f5RKo3ATEzR
d0b4kl/o6sw/0ooyyD0tW0buzrun8/Sx7jeodE6loyqH3wW1E7d0gKzVzlI2Oy0C
E0GAR4yJDtw1dhn1JB7cVvwwQ2/Wq6nOkvRmtfB5CHW+Q8sQKyq/SMJQ2qeNJ+7Q
sXIKbMmxJhuH9W/kEO8hOkoE93j1y/K4qhOjl2j0YmvELV8UC78sfWnAqiNn5CBr
N4kyX/BcnfPFGL16H9klDmVMPL2KIgX0+54d8iYwT2xQ27DZFQKjrG5oeqsB1ctj
5W5dMk2FgvUBk19pRu57FSVndnX+UFzfWBCcnbK6oobCYCVZsJTSJEQ0uV4g4Lxl
THrp2PjvNaSO11CpvPa9KkjJua1eXO5S52eVAEbUJuFqrtw+nN8etQR5erXLRfRD
CF9R88itky7DoyF+Bc+qvW35IoL4uKVPExJbPzqmlK1gOmZKoImM8kE+ehjZc1fP
CEdzGi8THgrydDY7O7FGnTDl9lVWWqvcl7Dxqt1znqv5x6vIZA5sQ3rDSt4Om4dI
R1sCWpS+nl/MFYfls9VrCSChzDH+VUnHtcXA4sHxNfRSIJf0lZZRgdUD3dKUeFnX
8H1kE+yJCIIP4/HbZSuTOX2yTXerAmQn7vs/emWSVmM/MHihjMcgrv4F8cWXyjw9
Ro6MmiSZ6OjyUlTkbxs/zkvcXeA9s93efp37YxgxiDcN9T97dfPvv0CmbYVg8veC
RndHlRwzENAROOKDJcJ29BCDj74enSlHbmHqCXXLVo+j3TXGmQCn8IA2ewc27biG
+27+IaA84Hh9Y97mkYTByKExZojwlvw28MpGDz8iVbxh2SG5RHit85EmxefeVt4C
86s7TbDVv1Irt/UqT9Ek8d8uI6XS2rcQ/VXWojYaC00gNiSebAgvgYRZi24xXmM2
FikJJrdzgq7rwofi+8yjWedEgGGqwbaluUkMxS/vFiukkkYNgjOPGg4mB3MYtpGs
g4+S8+opSjuLWXxwQQuWfkL2Rd5sslBv0zBlbve++j+oqj4HiTkUl+ohKDCgnljz
PRF5DFnW2t+7+8W8me3j6rPaVzQTI3A1gqH5o4rHr3PjRTuxcsi8sfATV06HN/o6
Q8u0mEGVm0/0dXsTqac9ua8JiWdTnPWgiW3MKvs/SeWInAjOmkNSvFIvm19zyl2o
O500PRJ3/w2zwehAJkhcaDADgoL5QjJ+uCb1V2OD8rjs8rId2t+HCVQ4hGn3hHpb
8lPJjH42qEoOFRTEM4l9P2pcH5xrceiykZjcgESyoAoPvPpdKK7ROQtu0QYJePrd
7jL3DQamz6eIQfOOcBF9fzpg+LKFbTBSwU/KBJ76ywaovfrIYhPmUtm1P9ZoP9Qc
mi5lPW0iA2Q7OcxVbZibx0srqUZbwB+PZgSvUpJTHwB1hpbXdHxYzSioCRd9V1Mk
seT1KG+ad6zelFaOWauJf16amNGjmtujn5jU2sD0bUi1YlgEJeR/arAhQHzTfP4x
zhcpkYRKrsCgMPJ5FXbzECk9qBx1vs3zKz2QfBdy+TIPVEMP6AHvwKcV0K7me/lH
xTs/wFTFU+voCp50Ksj89YefAPv5N/p2XhrvwV26kEZoYR6JeA3usLSRlUzSOI5S
ceHfNcDABR+29rquDysTlrVpWrh1ZNLrtyLEqEiOI6uGRDetaI2Rq6piUc1FWLrm
P6nxxd3kpm6DKG+wVBv6+T+cE3zdMJFNHlxZIUC32dHJZolK+mtPYyghqve3usVJ
LHHdMDuUR/ACAhrPNhX/+5kIkc8b6R4oHiCJU3nKLnITt3CKXewDgANSa0s96Vrg
Dfz+QJqhjhvjKcWERpw34kFsXUsi5W3CNaiYtL1W+PJkyJLrFMhoZaWQLIS+P8iR
dhAPPbLDKsqR0TMLPhYpyimb3lxhZj9jhCKKk0f1KMw8geDEXg7kwKDPQ901umjk
9PI0Kt7ZNGNARL9Xj55iOgw7bQgOWm6qcIc6RDKOBYgkt6HR+IH+G128jkIfzeVI
O1K4ORKpVoQOnDscpzQ12eqRiigTWphPfir/htD7Kzgq5kTjUXSUChH/pCpY81gz
UcrXYteCtQYzxIBKPqPeA1b8zDlJrY+32RNZvSHYpE2LSR2LBJS6fXGrGKwWP7In
RnJeNi/u7IZqnTY7yelNuaPTHj+eqehy8X2CO/3ukCBO5AqWuOpb9OYw46k/1mWQ
fmF5vPZDESxRjkOLARbciD4BANoRsiJ/xLWZc+N/BLFx/kZR4/ZoPTmkk/7FK2Qd
yHCekQ8Te/lCmyD6UFH2UJZOWdMWsmBAVUtWuK4jGRjCtTAA6DsKv6G4RP9v+lly
tIww1qpXLGVrNHCe2Z/Hv2s6TAimadLfgCBW1QBhWfDRWMMXpfGxlSr5dlcBU0JB
gmJPaWPIPzG6u6cSHbZE0tPp3QV2w1iPtwXNzmRjWxqzZgkuXde5JEHN7qu8IV7e
31miKSHM4eKEN1eGW6OkqjP0VSHANwebA8SsZ9DKrKLHd5WQJApQJZTA9dgb2r9j
3+9UXnQrX61/Z8MemA9MA2fTjnI7GMaymkLt9czYzqvJ1POosiCkg/oZIz+vHRhM
Wzyy9TKDwXLyfjp979MbYSzxtLcmlNz0yw9y7Ov5iZ7ejvDMLcQqZQbBJQG2ToSp
Czy+3Mllu4wiV51aLVR6Gw6ANJkgFoEF/z/XGl0Fhc+ha3uarNc1KC62MuJBoHUx
vcybuYjW0iEsYRQWHc88aM4l0KiPWVcUFq+slD8Vmjd3fROezPOgaXjJqt9TdUeg
7nORVeU5ajyTcCiynUQp6pTThVpDlQbT7yj82UYNRXBiYXfvNXozutBQDhkHRftK
AYo5hC/C0cUlIdOFtW6JSb/FZcHg6jdP0fwGgfrPAFLF5ZNEX1rcx0liO+xjh+79
/V6KGRRYH3YUPcTrT88JN5TQKh2dnsMJDI5YWWWCxYUOuw0Z/7j4JlnzzKcseXUD
sWp1/CkULKX6xaMwqyCQmjVd0MttQWogvioxNWHDfZRsTNpjNvU1RDIg71ELTI2m
scVpAnkd93BljoifHEhbaKpB/L4FXwAkT4HBbQiWL9R3G+ClMvAfNvtUjCa/747J
ntEVLgVyEop48qUa3g70xJea6I27Y5TFTtTJvQrhMybYJjDjxmbvyB4Ie74/pGmP
xxG9nh3wTW/T01A5xRa0wpopZlTUwm8i5yJ/43Kqxk4NDuDSv5jxslHL+VphOJLk
971m6XRA1gMWMupXy9vg53iEuooSu1WZJRLqNfDmPzFksNNvRQaoYN2KB5FoTvEU
3yCNWL+PKg1nycaoEli2bHDk0wU2KgFs6rUb0pdU8OoFbrx5WXQ9JmGHnGxYDkcw
auywv4Y9p7OU9G6tDXbcMe+ThCKLASTbAS5QskBApBox/PnmI+BvPcP+itJoX7Lt
5C7wxvnZIFYm4x5DXx0Ikv/zxHk46I3f0ysSWptYZq4bXPYneHh0J6B1m/7alN1f
ofczxY6DC7yebIXg1MErEws/AIIXQeKk44Yei0COQNp+7qvN/y9Tb7oJL4+GXlyj
wyOlvtK9HHhJS/nA6eDjRaILExdtTr+EQNhehWcKE8pQ4zctfRWBt7FanGJ7hmI7
ggKFpTODfRDK4hDU3xTduL+YTB26B1cWqJZdHo7vv9XYq4jPp7GwgkHqL9FRNnKb
3ZxKQri7uePIoq1yso6pGNLsjQ25PK5qo9WIk+UqLfNf92q4swJsTOWQBEc/3JcO
B4e8ZiWn4BU46bcc35zh+k+IFYnk++m5AP5nm+VaL1Q=
`protect END_PROTECTED
