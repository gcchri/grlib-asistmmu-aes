`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uHTEA0c2JuxgE9C4bAu5Paa0T3nnMq5CSEi7CW9WpH8GdbmdnDdugZ50qxh1O0mM
ORbYe+3WL1Er7Zrj1RoGzheF8Rc0C8SaKfUWcpM6gCm6ZcSgE3wyw0N8ZtoOP/DI
DvcjPVUQ+k70IzuTiqM4tFUuXLPWxUYuYkxg47DXMYJwNheKAmFM8v/5M4y7P4D2
BDzbJfVE0hhWCS1ILnE48UXjK2a8PwmTUUT7eZ0DrVmTjr8WHlhzL7WtchUPHoNJ
Gds0kCLf4ANIaSXH3hB0sPGawcynwj8pLTkFxdSkTbUQyJ2YaIyh3xl6cBwP1pAD
Hqdi7Uqce3CVwmRgQxDZgDljzNUFslTmhJHY6/NlhvBLb4PUkiNcizj0XRTKZe01
`protect END_PROTECTED
