`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FaInh+MPHPdogofFaDUZ/NNmDTsc8OLuxYKXj+BFV1LLS6yqSzdvs5picVY53dsG
2oyi1c+iHVKO0d40mEyUK0Peo9rHnKOfv6O9B0WCKxtbOlCR9XrpYKCRu6w9YjOz
CbiUIWXxSsTjoRu1H3uLjBr3zwR7vejm9UeNFuMg+ODKcBSIT3GckjvP+z+96uFh
Hx7+8dUqsgBt370Wgg+/jFXyqgS/dc9qnYAP3yMSlUkjGAT7nYp4wxluC0dBgEL8
KXdRqNCQhK86ZN00wzg7hxJNKjr39dv/oO6HrcGFJB8xvIWLYEKTRc0iUaiWr/x+
fE4sn1vpd7ax/Bcx3i17/EVodbe7U4E/X0CD1MOxCMgXkNjRLV/h3KAKHHCrahBp
MqmLM61M3d5o/puTq/t0Wsw7KrUE9r95wFr6rmyg86+IvTCXHTLwP1xH4w4ujzcM
go3i94/fmh5gxK0gwaE27A==
`protect END_PROTECTED
