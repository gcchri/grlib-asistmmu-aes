`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3tIEs6TVvMBi3+CaIcb6qylSSx7vWopJvFMYXWNvwuFhy0y2jqkZeHs/xTbtPumF
+BmV4yalEyKGU4Zt+ogCPbTGQlLDX069zisqUDAazYKeqowaX37HwffmtN9hy8Vo
d4qrV785nFTQl7hU2qOe/jlP3daJ3Kvzz8GDi6Y1bb0vZb8bTAjgb3cXU0VIfbLI
uIvJc1cf5xcfWDSMz8joxEwYXIk1SQqfGV8YazLykEDo09Bt2d6B2NPTkkvDcL4E
NuWZxsjR/vmGQLxQwO9F6w==
`protect END_PROTECTED
