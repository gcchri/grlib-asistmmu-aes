`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tEvdQ8EInaVyDVI3pHbLuYBhNIWX+lQSCeJFRD3gnOkY/TqEd2mUDp56UetKC4A7
tyemR9v4ykAgwokqWp6sv4YyMlC8M0j56NcuTTaWf/+Tw3KMRUR7HLbaAxNwzPGW
eE0uZ9dMHx/m7um04gyzC15FRgaDJ2fu0lUvJkrfYEa9KMVYgrqeUWS7VrZzW/1A
GgeoTG6mXl83vuoIuICQcsDfG2ntIniRW4ZzrN1fiBbZQyDqt7vT84RHtK2dOJuW
Lbme0nTzuGV/Nr0EcFvQI9ESqDmdFAunakIiHHQMekNYxjjzFCnefHUU3RxQ50I9
11IKirv+EMX4fNDlQvksi5SyRLZu+wdWbTLIDntzaxcu67SCLfsj2lSTZ5lz3Btt
XMIuB7UAkKm+Kouwj/UzXd5NOT+gxCmE9AB7JzXqDZFUBLMNS0mMgOyf45Ebsq3+
+l8ECdNJZRAYi/3xrQKT84N04/NmPWgBlXexKtOCrXRe1Zx54uF8Yr4qzvRuZCpZ
rfTB0RN/mRUoCkEVUiYudg==
`protect END_PROTECTED
