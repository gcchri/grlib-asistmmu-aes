`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9QeGAcBJOrMAuJ0j4DWNCen7E7xXY8OM7WjL8h0ixVoMpYI5i4w3CpJZY/d5CBQV
9inujEMtVkbUL0WnbVjRDJXOtzUJcjq7ULp3Pj1fIZFKUW5E19yMvh5ozz7m03UL
JaSHmL8Q3XWa2YVLav/uEapZJAM++qHzuc2wgRXyFcx74M4aGkHJKvyhn4FqPcZa
bfxn6HUX3Dzc/dRGe7JsBAZ5uUT1iL6Txj6YO7YZtPe4uejADpc1lXRYsmg3FXTK
zg85csJ2F8UovrHpaJNbXA==
`protect END_PROTECTED
