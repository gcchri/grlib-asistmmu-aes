`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JbjuAIVX5dreZquHFmdqyfYA95XdpIyOlPd4SxAHw+M8+pnAo1DXPWHF2SCeXOBG
9o0HGsVwNOaR3JU0gYyEbnuD83j48lErcy+OVOV2zYYx5Xkh4dud0dDc5pl+KKHw
2iRZSZm3HwMwzaMt/2BHJmWIBiXzVn7Ce4Rt9jQhEVoRMbo+xawwdrKGHximNfPF
aRLpCaLJTygMeNdWryOwiX9C79ruFXFP+ZVYlAT63hYRFrd+D/GjwZmMUQrvHKSz
qE4BWU4BUbuLe8IFT8xKAClmKgPu4ZE1XBKrxrs8jCovYIx5wB9q7rbgi0IyrjuN
GeiJ1nFHNRhh2V/hmMY+DXDocy7ERBlwh83mHIxiun7vw518xmlbFGOt0n9iO7hi
L+knZ6UK1LTD8OPFlyl+OPMvwVKtpg1JL0SRwHOT0GDk6l4cdFCNCIbsW8/zZHPJ
T7FaD73uFK3I8CSR5RqTFl5ggWCHGpSH868b6v3OGF6IwjwYqllvRA7wMf/AmpN4
r/Uhj9STNLw74i+mnAZbas0rHHvXyMOnQTkwsbILgfe0FiSJuYBYxedQ2DefAPNH
Fl/cpaUMFdZpgEZAANcLFkWBCJRt463OvvKzCcd0BAM3q96l3cicEg3zIix8Dq9k
IDfKCgIoHyFP2mLAVcPp1ity7pss7D8ECQ7Ai9tPa1/kRNFEl8NefsOuHVdx7EbK
a/91WAIgrD2wXKl3fsysAA==
`protect END_PROTECTED
