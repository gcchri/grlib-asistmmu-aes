`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0FA8pmb1biPtMxfWKm1IXeEb9oZbVXUPH8ohlAFj2pOm2fo1dKJxlMsCiBF0j9UI
5AX0580WYAgyF4CTF77vL1YVHSrQihJ4ephY2EFX/qaJqSfrSrAeMOZ+T0Z2sT7w
fkZ/0QrOqAV7e3OSVOeH783ghHJQqsOsE3BVjLOLmwEIlFROI3wSHsOYMUqmqO4I
UmHYzih+SrGYnx3HH/0t+9NLhRzffTAPpwMc+rnkhhJQp7n95ClSprSK2V11JmRK
ARBhajvCoGNE9Y+XaPf42QaoSBl2MEYUEcAy9xrOJZT9YeaDtdn7TF+NSjM7zNYM
8KhRrp4MHnVCX4RlGWUi08oWfxz8fsCSz2GUtltjZXt2mlY2rtnhrlanFFYo8eTd
LA53gA5QFMclGV3Bwig/ZZEUJmQQsT1CM3C52//9BHE=
`protect END_PROTECTED
