`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kdPKHPvmsQezRIj3Phc9E9m1LGKlYNq/fSnFEmWlKhhVukBlhruWKhaDjQnVH573
QhKscfNU3MfouvFdDDy3HAPr0PUdquKyqEZwPCduekWs784BdsvIXtIe5RVZht6P
9kzhd0nz2gx4ghLEFUFUI7tsWlnPPVSHl0GfDZwJLYcjR+7xoLeLzpRCApqDLpOC
dkTYYUy+jYbyAazoayYPb9PpnOahihI54mpBjueFOaZ1Hv6nJugl6LaGsm27GiMy
Sb9ViqllQooZzodaa9tSWzYzgsruJ33FTLHEZFvS5fwGIMDHQWBQR6enXOLqei3T
FIoOhlW/d5TEAkXFmjFtFSbGZaSLSimI7Fq4WgMSk895cJbhX7qbIZFVTzSYDEYR
HKVEw9mGLII1N2MBtETJp9fJp1bK9cgZQnSZs1+L3mGEBUmlJPRa4E8nB5oRXeVn
Krj1crIDHL018PQCK5td7RLVlWeodbV/EHsNtdSUxrdFNu4qjqp7i+rw8HRWocJW
QQR24eCDIdaenS2ASLYQ7V4DEsW0vLc4cf4WbAirwwE=
`protect END_PROTECTED
