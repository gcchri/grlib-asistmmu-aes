`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s9YmEUmHQgtJq716mO4NnCRjWQoCXpiNx+yA3BswaCLu3ig1sFIuGeC+PZM+fWSn
yHZwuxLx6z3bj+zLZAafyW1V0UceWkBusbbqNWKyIqPga9L5m6e709yV4rSf7VoL
TtPtGlPloXZ1fTBScmYA6AgeOabhmeNYJjimxfOWWxI2nUgfw+kmZAzzUsVuBMwk
9nYswJ3fSj9Rhg+cBEL7pMW//R2R9N4mlASW17eluNH3EyqidDYSKJJ1Wq9LBCWW
IRHh5XbABhdLQkpHuSvhIUQxp4HrOt6hEtCtBoSTUPfoGTa+n63+UrOWl9VnjaeF
+L3BhEUbJ1FPsdXKCrd1x8avNN1qeaT2JeXHE2gU/h+RaZNjIoLTNFYxqGKE/+rt
BcUeM0qPT+6Zf/bh5AQh4RzI9EJu6MErlSn9IUILqndHgLhjx+4ftjmghPZe3lO7
`protect END_PROTECTED
