`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2kDEEZLet+p4bBQNKjmTNH3FlueelXHQ4jp4NHp0qI7bu5fSWT3daAC0oOmBH7oU
MRdaykJa7tLlZFXlG0aWlriOU6QFfarPt48L9NtKouhYRG22OkW4xch3YUAV0mE6
hHa6PTH71b+do50ywTOzJp3ke4dk/30z0KXiPAoh9OAiJ88swMRZnrafhbQjYdHO
tIkfCAJTWcSfyXpUjUKePVxgH3xUCg4RcveITcEdThEkcdECxQ9864jLIOG7RmuK
+Q+Q6+pMpO/QyV/Ss653HPAsse4ftLfjn7Qe+4mT8MBSPP8sOD5B7yW0t4hV3d+h
Nm22FbxjFX3qo6tb1UWoq65/VoICpNwU4aGj5gshgRAj3w8aTHFKQ5WXk4ksEB4E
eG/8gXLMwoezDZeeLB0uqwbRIq22FMf/H+CfRuSkwW6u0aq2IuRyupRtU/YbatFT
2X2UPJd2C7Za7g++cqalr+b6u+8j+i6Xo39gpN5uYlyR/D2TSLZIGPIw1co7zRL2
1wekq5Nuk4pqdn34o0ADy31hn4g72DY/lZI+1QJ5BiXygXmyP17Wni1O/C6pGAvV
TRU2hTf9P5pL/IKRdpmzEUG67EAGWauRomgJBmQeQAZT45s2EwzE39EdgnSpfcIn
M/lx6TaMwAEiyk2bQshwqmgdJ/6xcGiwQJo2/iOu9Phhske5BxfWfvX6McujIR6X
B+muoFXeeHmzN/zI7GLjZV/ezy0equ4vspUgSgvRpcxZNsJq/i7+lkkcwx8QGEsL
fdUD4rSnR7oUkHRGsKyVUQ==
`protect END_PROTECTED
