`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XRTfOdulYUVAYFj5DJLEH9lWkC2/PtVNjZEz12c4hiFxw1q7uaEJnyfsHLKQJegg
qwuwbeWK45in/zA/6+ayudvx3xKLzl7W1aOHj//1kL9wKWUjc27NYDbIH+T6SxcH
Qia7YszfhQtTq8h4u1ZUlDQoNbbrhEmPtTescNpxFOEoz+8tn9g8PokPm1ODx+MH
FLbYGDGrGEfF2LdlHP+sgxQO4GkatX1QWmzhQjux8SYTXs/HY4lncIgdoYEy9iC3
EUID9CP7ErxxX7me5GkSdtr4M7/stzc0OXLbPMB7G4wO8b/bwVwLTiEne5OGMidx
GFEgJEVn7HpKaW8Zq9cO0Rv3o2EyRTWJd7yrL1RqP0prQK8VYz2eo71pPTR/zwSx
X0eqBn7qf1AlCY3DZuAGQctC7Yg0wk/8WAxlPPMkMpqBJSO29Wr67repWB+m94dJ
sA1dVuCc4qQ0WQ1UClXPGHFdVKqDKwDZ9v+J5kkkvop2gR4dUMiWnxrdVgS0bFMX
qchUdk2RBzMkTbMbm5tsryw6qbMvwWCYKG3yE0K/Ra1xXMeqAnRjJS7qFHasUr/8
9fMxzLDP+gnzyIQFWXN5+GjvIkRaQlzQ/au9kwuONkGMmXoZPvqqsd+FYu2sIvgr
U5HMHNJHfDzEhPcf23NsrQ4Xua5r+d1Nru6md9xdN1HHo4eEvu4sf2++fZ/upUDv
u/BuHyPEg4uzTK3iUEFfzrZRDXMThnyoALB/8hofVQBxUbx1bIACPnFXsYQcb0y+
XNu0cEs1CeQ7KTsSHC5TIqpLK8Z0BiBzQL7+1d8mashCTih7rpYdIlMpkchW500F
i7hxCNWF2CYD2pnCbEY4oPEQF2VHrVCqW2WKWeALvmvp2pc4ulSCi0xuqrGWQAOG
0tnG1Q2rVKisJQdiBXtFA8Zh7PEhKaxxMJuxokHaZsARIToi/nbg1vPLh9E66no5
hWW9esAV05HVwmgnpnMEwvBjP07w7ACAzNd9FUOPXyx7Vtrdm5kd/z5xgDCLmCqU
gOCE0ochGRw1gICmCzCZT3vmH+KQuRUjk0wzikDgKBPnF8cKXqxZEYAypwX0He0y
c9wqwzSz6dzEWcNislP3f2wZak1Tsvv3m91MVahdAWCji6w2NgFPOIjxA9jR+eqJ
yswyZRQqj4Y3pqh/gTSKHZWbeaItEVcQeSx4j16sjvE2O2ECFq9BFIgvSa0FN78J
tWSmfrVQaQoBW66hd12Xbdz2kbAylqF4k7mlp9n0okL3uW6hMVj5Nq2x4g5LXJhy
`protect END_PROTECTED
