`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BUq5sjBct10ctIzDdM0yzAU1qBiPRh2MyrKWLo/ApWFCAJs6/Oh6BsyggS7dBdtW
jlWd1kRglOWpfqiHmQZ1hLe/nSxvE4/cKwzuFMv9w5K5vbqbpYWEoqiJFSsEhKjC
oRm5YiFtLah/TuOUi4n7uGujqrVaS+08XaoYicNQD1XMvoHsgU0gl3LtExD6cEzv
kbBtUMnpQFgBZL4tytkmplMC0vQSh/4uRSrcdPfAKdncPh1BLjuL3wYwo2/C8ghb
/E9P7oDqWUyTdYxuzPEatAMbcaAq4hc/L9/0klik6War+X5QEoXoUeQXtow20HK/
MwCtj8qMvwcjyMj8lgSuRCj9kju4A6/ps2GeZ5giUZTJE2EPjp66iNKi9vKx9FoH
yE0JsFqDYAetSFkiQxpk1/o5+LNMkd0/GjG19fv81Hwd31mPeZWu0bIVNiM4aK8N
/6frH7LwmthapAZdo69FNk0u2w/PLVqbO8Q95Zb1grmm6q9a7+4v6JqFy9O66g40
u9I/x2QjTsa9I+ynutLWdQM1aXxW0TIG1E5bDzclrcZuFvjxXN3EZBbPpU0osQ33
ld2f+rwRZRUltByFjzPIFd3HTIMgHwg5ciJXwJ+PU5MS1raIZDQ4GMK82xlogqOk
TtNRyYKp59wcKcUITNp8Hg==
`protect END_PROTECTED
