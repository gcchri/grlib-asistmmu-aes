`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5bYuwGZHoM1lKIKw5fAauMzUcOINd3q6mbHKNxEm3WYU1Y5/9Oz0UTUj9Jbr4VsH
tcpH0i8ay52ST3t/AbX8sknlIl1UjRqdTfIqhG/kHpaf4WyETzyNyWVY9Dv0VaOt
jNYtiqQMiDoAGw+psUtB5WugjNM5IyNx427WOfPLHEX+TvW+mQNyzUWGXdf66xCN
+N9QaD0jxbGxmaczaR6UJy5Ut3g3v0UCTnj7j2ejo4FVj2D80+u8hDaSOy7qtoZC
gKEjwarSCZwq/1VoIIEO9wiaBgg5tN1idhbyOM/mMJgS6T+ZywpTep46dTy8DN7d
fBy1JvvAEuc4bHaPKKMKAEgQZTLb9tEfps49+oRHhWusrgLGfbgayCLnX5r57YOU
aUTzk6lX/nq8HUXiZj+Elw==
`protect END_PROTECTED
