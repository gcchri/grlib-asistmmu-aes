`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bn93B53UQVMxuL9DoxU3INdPYpbSZKEyheEsjh8oqVoAsXyllJu/N8CY4IqQYjDI
CcHN2wwmHrWKbUiA5iipmRT7hpowj7WuI4xlBKnsXhK2iAL37Obb3chvrEZ7gz1T
yP4EDGeJsIUvgCIiZU+BOgi6z6EwZf8Y8+lNLvQGD80HXrsBLGPRs9v673NS3WuS
aXnRWCPdc2YhQEhQmh5DlvlNUgV13Xoyes1GLybgNZV7ezLbXpn1UXgwVV8zKjFm
GGdbEZvwKHc2LYMaJeT6BDCL8uBT74ZweWS0/fFwTCM=
`protect END_PROTECTED
