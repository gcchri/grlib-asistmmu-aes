`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hn+a9s8DK92HjN26ApbnONoPRiCb5PJ3F4qEFxRqR2C8EoWlhn57Q3UCqFhT+x4N
6/M0muGJivHW5alKi/DU0rOrU1EOxqnE96aBt/rBpQjJQifTNbTGFQ5bqS+qf65D
6wPznAHvhuym7321O4avsRiUN52QfYelzOFvt6cBTazVVqaRpeu5I1HmpRhyBhwH
lQldGl3KmJyM3v9KB2NGnO3mKBL3slHnO6ic3hc/omZTwZuVzhK1Hszrv00VWXoQ
FS0oNbXTD1P2DwDIOFWH6OUmKk/Msw4D/L5RP3ExpCnGnJ7sanZtQroPheQb2TM6
4JF9nfz9GJBb2wjytIndhA==
`protect END_PROTECTED
