`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DWnaQH5rZh+DJ2Qpz9Hk3g9m05fp/zw/UOz0eSk6spbFCf8KrpBTVtnBK1aK1oo6
Kip/yd55SrUIBnrChR59FHAe/0s3YkuoQUznSLcj2aD1oZl3BxO+F9LmrwXTZkjJ
SzByCfgsEx6eZ/yTjzM9c7GKkCcOug7Mvw/r2ozShxCkVe12j8bZQnd+E+iRVvJ6
7Zd37THNzrHzkJmp5qWKwR4H8/hWrINMWthj7cfie5ndX50kzq1O5MYjditrh7pc
0ZcBTrbJ/tJvt7a6/i0T3LQy5odIdmHZEC9h6eh7Phk/ziT97cepdtycl+rDVKO5
NsHj0VF83162lHRFt4jkdxw38mAzIhNVsRiV2XvLV9V7H4W+V03PQme327tWirl0
VAuszf7rBQG/Bjw9DDs2jsukG1A+WL1uP0/gh2u+xCwt12VbsDmoye/aP4YpHVqs
cEBudEseRK7cMyGgo7za9rgaglxfobdEc0b8v0Bvc74CFimTxqQQliClsXYtalgL
gvLvO9D4Vn+UwyI3otNYPPE/ODuUsE3mQ9GpksbrV/+VatsMR/fMz1IXBp9L7ZYf
CCqqQv3ouYJZkzq02/NKHqI8KKyim0N7X0wlDTBrQ//9ptYn5u9J1mDjdpFbpJAv
T5a7fH3/YoQ7cWxMJ0G7jSpBLc8XaGVtH8GYnGAjSvXURx3XhLFkNVi0lsNmLV6a
bf3AWiRrVORIe7wA8Zq9ca4igwOQCszzaNVoblppjnU6kTvY2UjNgoptqQE8FyJy
z3Qiw3aaLan/VQqRHMqDMMKauajqV15tErdTRJXYcZ+6yim51OET3yRsMmeW6cbz
Doz1+lxvjju29ddTt+s7IhvtR8kcxvgEhK1L2NNgeqtUhZmRiS/cg0NED2nqxlNJ
Lr78UKDzPyGabeZHIEM4ZPGn/YvQvOqefTmSUTwO4uo32INto9u85/HFWVmZ/jkO
huyVCT4cT/oTZL9lvsTpcyagqSu2A2VY/jW05oTrJa8gi4TtgUbrzH6uOuUoARHG
5toLJDtVKcZq5XavbfddDLtlTDy0qPQPxDfiR1cZsy3F8+X5WMQi17c3lyr9ZnP4
0y+ze3L+O0fATjy5j4Li7g==
`protect END_PROTECTED
