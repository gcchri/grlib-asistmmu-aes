`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I6l0WuX45IC7chxB8Hn2ktgyA0PZUn6X6KPrFKhihYFXfDmsC0hgn2F8qXsEHt7o
7kLOOpYy6dUPKPYmRIhbrcYzWHn4x1CccsEZgDm6irAEYhofhwlalc0FrI1LA3ni
1DgeI7YfM7AcqqR8QMgOL9/9OdrQHzIr8LveGZnhn9Eez2Pb4WeLclDt+LiwCfK8
D5czanu0cs9CPUdS7Sq7nx8kzI7zS8+5Mx7knDUYgzl5NyH7O7fLCvgreLfNqAts
AVWbUeAcZm+e6/ujxsXGYfA3HowVkjgxrMOKhetOzYMruDqt8AMOjqwXWtc0RPp3
Z0wXx11jT5enCPsPJ41bUzkzNW8YWyDgpyPQDJGJRpDY2kH5dMQdahnXMcONCp8Z
Z45b5PHRK4nrZueVnJXrcjT9A0fGT9K74hkt6dXp0pzoJHNkV/iIMyVCFgJq24mv
sHAt3zQzMs6jkJ5iYMhL2YAyusL1uQ07KyRzr1OVQrhEVtjgwquK7+SjpwOpI2NX
/6MIsgEXF/GD3yytOFBnli48c+Cotr5cizmZq92SJbL7akMjyYfNSlTaCB7lWkOU
WYScj2mkkaXAc/Do86jC0UKDsmyed2Q8zwifnWAj5/s=
`protect END_PROTECTED
