`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
st3QLWMR8Udqu4ukwJhq70wma55dsd4SkYc5gbeoQ7MwVxMWY/5Ww8kETqQJG7LF
kJqzcbBQv0dU8b65y9xxSjiCvarDaOYTBp5SGV0HbYWPWdTpmdWYympACfj9oqG+
whumSGj9U3Q+vP5VMezrDNOQ6hBo8a8HfJoDUVKaTM9CadijEawdysCKdn0OiQOc
WEogiGSRr9SJQ8kpiiXBOcwTuXDUtU9efnb01+lq354b9HE2Mb2V3n8A/6fviysA
kCnYC3yAApI1CK2c/vxCeuRNZRJCQNcHm/z9B/Z8WKNlD4iG23fW4PmSdz50FBOJ
s6qQROsaoKaGU+mBqmU/WW4WSTs/QelLPagFhYYG4S3lhmih+Q7ixTLsBgnzFD8j
wvdORJJcyNhK1Tv953kfONl6LiBAaVckUpMNSVCMxruEajm5r92mSJx7SgB+m7mq
7Epej+QxnQUyYUtKDsV1EzJSPHY/Fc0ewZotdmrBkqb6tT8kRpnmffAFGhwTZl5Q
0uZBia4qV4hLi1e3E30eOkprsfpcVuDLuBgRIy/ZBAplBlxYigDKW7SS14itzS5S
ofyCWNpaWEyy0DjyIFObXhAq39L7WZ4SFNqGu6dtJqrmAywG+PAIhVlXIGwtpY41
xrV8D+0J0KHx3EQQQk8OSeMgKWTAFNLNrK7sUdgALDfOOHUI/LGfgCeY1BQi9Lkm
Vk5Esf5VMnXHyr7TuWHfry1w/QFzLYvQWI1zpVXKZuwJcN2/8P/MgP5siifDtpUr
meE8HDbWsGHtROEkPifoJxgebSbeThNOR1PehRBlhfTanEXz99rR/mvGI58gLoA/
KHlN9GPP9Dp6lETvYQ4uo2cW5fHbAHsTl29D7aTC83D1hP3j6RFtXKIVSFeJSuS2
Ptq+nekz2gVHA/qxw2dajpfT5IeURm4jaBf9gkjNE6sPhBOH/j61uY5Ulotu/sim
95o/mUW4v3c++lCrE3CTPwha+eM6wbLdyoMNaKZKzZmgYASMiA3SFCpP6Bbq/x5e
geJYjS17BE9oMGeXgWnhFFx7jSGMCWntGGYy0oUp3t15oyHTDwEyobvkBrLcwTQL
qjZCOBrhwtwfdvK9HimHitTjuUCZczl5aPDEPKviLJpBh3iB2CNfPhDHneNNTUKC
KI8ACYhUMB6A4m2mt2i+F4N0RijNtwkcumVcY72pqHlU0hQGmyXoaHWMZzKZFHSQ
ibv6NfXLcWVLCxiyo7RBiUrpQo7Jfkl6iqByiBsA0w/qD/gdEtA2rvx3SwW8ohMK
/VJpGhP1/TMPqoAs+8PFvnxJC6ZtNjlpQj61014xboAMA2+NfAo1t2eUfR3T6HzJ
wJazkMxDfpEL1FYSPQ77nxU5CGS5UyUYMJbwD2MadZ06xiyYXsJOnSRuNevI0Bwo
z2PbzOmQ3hOIowPihOE1u/XHjk+g+inF7SVu8+cpaj++sHcqRNxI+qk2Q5bOT84B
wlALC29ps03Z7DD9V3rymTSe5TVgO3WlbrgQUcjfYedSNiEmHAx2UwYBz0gy4IP2
SL2w92Bp14zlLtTxZTE25szt39KO73Iohrm17vndnse0TuLZKWY4UEICf3X+9TU3
f8C9lcEaVkiG8jTPGcUBLPlBf3lqsFbEg3zptSN9Kryw7Y2kRZpLdyt6zFxUh8ZY
n6iuo9rjNl0AnoERDlh9zSS95X49xDXz9O3nliPS6Gc7lawoRmC2JhC5dIbvue4P
oW4dZInhPIBZ6oIHvZA9CozDZ0U8/MSKNSVfQj8z9EoA8A0s+px4jy/W8o4hkIlb
JlevB/3DDfezA9U6F2WLZgzubIyE7aLLz85BHcgnsNhLajqBrmAVOX0o5IZQ99El
Q3OKXSCunh81rrK+qxBWeIdM62tYi1s10OgN/wGX6aeLT9eTUBPAfOABNxX3Xvmn
G+yB9Ab1DucZfcGTXbQtaNqTN5p5CcVDQj1a8YZ351Y670HVdfwLzBh2eMwEzOUq
JKJFS9S7sTLQx5dMj08jS7+A+yUcnmVhpbcpDP5wTTkt0xQNwwZOdBiJfz3vzLkx
xG86pMjo//jZSl7XuCYZ2HQL+k/zZkoh0zvAr/KvrTEg8I7W1/2kZY/UDR9WKQnt
JalAFeF5sYABaB1nEGPU+H50abiYDUhXbAtyel2TzeQyAD/H9gJUKrMo0V3sjonK
afcj9hIdJJk/vYJrZEuOhaozHNkre+2L05FkTs2QBf0J6r+cEIpdoTjdbsMFYJ5h
rAWwRhEVyGwT3yRdiovfIoXlXAeBIB3i6KrikdxwkZOmabZJ/6tXR90nzZp30oGG
nsVcgkNRXRDzm38/8myxFBGgJ2IFwT+FkXhB0QU9eFx3vpJyFrHqalmrNhZDRw64
+nylXjSdemmiW7O+QuabVR3Vf9n+nv0re8UXT/WCeEI=
`protect END_PROTECTED
