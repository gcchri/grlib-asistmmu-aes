`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yv8Hvp3PDPOS1wHlRnItl1qiWweL9wM/FXD38ZXd/KQcpy/4kcXW443qf00JPQrB
mTTQpeETObyoglxHmhfMxEBzPyv9bqYOhhUQCoJP+2hy2DVx3Zp1qtenPuscITTS
flrPZPML+Incc1La354ULBxeQ1vXGXLj87zCeX6wgNQphfhdiFSW4+9Kyw3D2RJG
3qmRIIH6hAeKZppYsptj92qjKcLnS6Zi9uqorqRwcGMmniCGvtWBhljnlHP2MSds
ZEyLDgWSshTvshA7RbbImRhkBNGK+JCLiZzhCEl8LqKFW8Ayz1LuMUUhCuYiI0ZN
K1d9nghDDpfgoWWaOB6aspmaH/WwH+1INAwJa8KLwTwwd6mBdMzZzlCRBFRmyynM
F78GbFGwezi1ZsfxwXkdmxYvjZPs2kw4SMEu3W7yb/Tkh2GzfysgW9kPAOLOmF3t
JrbgwumB324H4uQoCbGFkmQcIC7Vu4dPUj6kYTvaa8l+662OcRkitklBJKuO/pqo
rklcbb7tqsECbbGCbAybO54QdXu8BTK4/EqHwB89N4CbapRHaVGpVr2+6W2vvzsP
7P4P/1m/BYtoL/2HBK93ae+RChUEOIzYbxC5XNa9IiSQBas6XYToSQxUmgMzSN/L
zJAHRCBM1jCs3CKgvjwc2lrCwKKpn/I8XAoKvog9Uuc=
`protect END_PROTECTED
