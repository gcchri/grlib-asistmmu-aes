`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iplKLwC6ZPwyR8Shp6TTvhS2SyqDA0B9INYWJVeOMFOfHKqu0jwdu0UjMueNhb+z
/frb//cUH1E36zhwqt+9KLaZ6tGFDhUpSw27oiRSNQT/6xPbVJWfkrY7rn16fpn4
9avD/CjVbO+3TeS97ddAK/ZidYCBLIakpF06vCdZ9O9qeZ1PYM1tK7iUpwk1jxBc
sABF1rceNx2h/SO6unpzQ6ElZAkvjEK5mAqNO3J/autzyJwtclMBp8ocPsJZU3Pg
NIb7ZW2S4qRI0zN5GMGP6KcU0Ct88wJ61m5RSnYI4H3Y+rhoFECgUkQN61mjfRDq
AQWtZ7dXbkr6+yqao2KUNFRbc7asIi+vnyXYPa9NnFLvNsN5xQkn4r1lmgF9WHk8
isz2XxljDRx/vFTlBnYkZRUF73FslAMtp52/qRfnMoeQD5lFdtyVT0BP1g5rNI1U
kDS9b54tG32zqM561FAyk2yVHSUOpfrawIkbSjxhaMSfUwNLA93mYwnMlu4tlGFQ
w0f2N29J7nM9fZbLfC7EKKW1D6lB5erCAoVJsLCla7KFxjvZgKe7HuZbMpNGZV9C
8ihb6jFGfv5H4FTaoQ3RQNdhUYqEb83F9oxJ+sMv/SL9SRHwJfZr8+cfcGqxlejy
LclG4Y5WgP2kDPr3a+E3cEt/NIGNRX3ksjbRiLfLNWC4dHIKiFJzXE7q6ZFmEREa
wtThb/C6Swh3OWHfl26gULnpJJPBy+1Umqj2XmsftxU7KAAqYTWKVSeF6Bxc6gLJ
gDXu7w9yIU50ZZHwLty0XDMiHLwqaEeKwY6ZqGfjSRb02XubToMZXOAOEU/LdN1A
ciYnjdvPWNFoX6siwqB1zKc6Tw4B0Ed7VzitN0HcOjKgPyutueRJPZOJ+BFm11Su
i/M+V8/WliEGveq7bsir0ai/t7wwQF6A9/1U8bgS8DJESzbX0mU9R5LWQjfo85hL
QjSswf70I+2CT6eOKF8uC7EnTvdGCyNFtdeN+uM82l/6ESbpZ4LsqNshfwwQPUsy
OS/8base/MgTLYGpeDINivgoiwSTrWgHL1SsIem0ZEiLqlZAK+gNN6OQfuSBOv3g
k5mGBsgBNTex/ppZhqZRf1Q5CWtBX7LC+Vw7MiU5S7QVujoXaCRp/AvPfY7n90G4
zIk7WRqK0+FtDjhqn4Sk14x8dF1awXtIkifI0PM0FLc+oxD0oJpilJZqWn72dnFZ
Frg4f+tJPfps0dEybp7SyQ2y1WgL89W7yGFKxta/haa5rkazwVeCGd1RPnP4gEav
hrr3WBSIgzk+jRdioD0uDekZfzfeTfAwJttg7U33MIwwkAbmU3wHDST53P9mcxGu
aQEKKzvjcmFbv4bWYE1U3fbF6Hp+0rLgRmZO8jGNbOVHjH7Gg1OCY+/HAjfguG7y
TQpiyHk7mnxC9zq27CbeIVk9AL4FeTu+8vxdS+Ud2mFCIGdSxL+Cmv3qw+MiQ1cI
1hiCjRr9I1eGPTjYURQFyYzTtInVgt33S74KYMqkdKOhJLf3vPA9QVaCu1lyzxms
AtHcC5AMbHzwu+rW9JBj6H5bmT5svnUCAA/Bo1tFY5sb1jShtHTf8HvlIwYN5iXU
AleB5fgD5Q9gedMc6u/RQIy9bD+UmCBLCq/h9wee7ykt7aGj9/wLQx9WoOzDks2X
hu0qaSDoH7WRkjx2o9M5+B4nRqqFUOZ9ktFEZ/BtS1CjPE8k0GmTF9OFocKsoFAJ
sFytMgDXHK9nfDemykYLTHaC4c+BNwhtevd+eiEbmtTBBZJLGNENxD12cm4preer
xHmpSjxmEdXLfqKYvoXc8v3CYhOALg850asixFyY+xExxOsfJkiEfAxIQLhU/HOa
wyv/HunHi0hYjfV0RwPG/VY+MDSDJus2Q7wfaJnqkRRp+UuVTA6QwI07IWFdPRR+
/JRe6N8b5OsVRoZA4FS59sJfmXBQRjhA1zqjmj+emefkRl8AWOw2ZdwuCewxW3nm
BhaVFR3vWdtBMKv6EmOeXauPquQTEPaNsmb/OjUWXl9RGA37GNj9RzqY2+Tp944R
RBdfmXKddFduR3t/TrEAxPUQIUPzKV0aVlsGGQy/D2BdJZ0ewtNUyeQoltqI14aw
HH5/cMxHZr6gLL+NHF3l0KlHxVhy3DjAkxRYdyR9gaJSlIZZcwkCQr6IJHFeZTV/
vS0PR1hly77hGG9h4BIuUvPJ9J2ImuycaA2+DRqKDMTqGz9FcgnrLbShw7js1uqM
LYRNEMM2UZ5VxPsxWa7glF+0a9WZAVIZt7w1Y4Ct764QfiwuEeJG9lYrdkM3rzBE
vRkol8kmrhPyZFMLk3ioEEgrx9sNALoizrUon7OZBgGTkPm8TguXAASf6y92kOx3
zIUJSFrZ524J87Q7wbaatGDlPAOZLZ9I/BEcybb4rMfCGrJKLfKLYiV1gdnOKgMQ
8436fYj9jpHmOYOEBw+K8t53gMwwbFQA0sbifXohvaZwSJKB7zzV8Tastw67jZsf
9rWBVZxNoMB5KE2+ANjJT7lyE875qZASU8f8xYFPnkHDezQhGFWb2Owse3KTDpUa
PYsj/Bj1lbVwSPap3SdOKWSzLyFvF/u8tKsnvHcfuaOoB/B7EtRkztrh0VpPQiQB
VIjZkrQzK+Qz9qBtKhG82+JkhI1xhv6xFNa+QgPjwHg9vVhFf0Rk6+e0HRxYS6VF
bv7pzBYe5Yo1m4Mv395so0mKmI2F2cc6Chc9HfmF6dF/UMF5e4TukclJoDMU0g3j
lQqvEVvZAffV8ZUH+Js/GUqCxQ1byvEowVJWqi0zcrenqWpGjatXO4bT3Oja77X+
ymk7iwPNMkL/1NFmgq8NirRzfTJDqgenYjYftSgDkJU=
`protect END_PROTECTED
