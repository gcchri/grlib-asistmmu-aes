`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GbTYqw824lHEy6psu87mciJy7RFcO/ag1f/iEC4oynRZKhbo2dByFL0jqTLIdDx7
pHtPH6STqeZeWKCLcnI54/ek6oB+6Mu+L+MTuYjiNMggT61fw/6aUkdtifZncpuu
GnfSl8SMI28rGYq6eB626p9H5a2N+hMDTHOPMcTcAxWH3LmDIHOsJzIn03mgS09A
9pqk2h/CHSuJK/E6WiP0vBbGczFUNWUJHGWHwndx96es4n0bZtM4aOaIgPpkWsz9
0qOqGpvYfBGm6loExEwzi/dmkKataR61O1XLsiitt6J+tyJ1OSesUFflPAjhtP6J
SG1dwP7e7jjRDiKhuAhQD/sCEJ30vtg7w+8o3Nh9iNIzNMPCHy8QjzRTtLeyyNBw
Viay/iqfv6IgYMKgeKOCc0AnKcaAY9t54sKQMydFO9fdYp5ozfOaK3nK+xlLO3WP
usm1I4Ne7VZpRZG5kmQYJVPxr2bjk6jY7f8fZ9Gql2Ay24B/KIzOVbQPD3oUA9PW
`protect END_PROTECTED
