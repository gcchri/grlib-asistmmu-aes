`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pV+DWK6EV4L1NWBAerbPTK8RZJerTb8o3cfvfOLzcTb4AOiFKvXuQ+xsL1OtRzWl
oJuKe3u+aK+9HtdZMrpgKkuNi4QgaXTii1Et2diVJJPNHlUgj3b2GI6ZljYVoykK
WyLjkaxIT1L40v0r9IoiKKNCoiHDhWujovUo03jmDreMUc9RO23FftmecZY3H1kI
x6/NjbZgeThcVLoy/GcE3VOUw+jIAo3JPkjUgsvmKXwsTmlwqItMITdV3mIM+zhA
BD4ETJSrQQwEZ7aOhz/yOsB1Xmvq3+ZIswN/Wiv1dnbckn3xdUNL0nULG3sSiaoz
XlpLAMLYpQsm2X0Gp6VNMky9/9OaQeDHRE9f7TtBxXYap1iCpQEWN0gIjfpU2Teo
za3tD0OoBNtG7qVgcFH8nVY8PcW+2mqJ4gaqubecCCWYWKCK/06CzQ+9jYjPFmxG
Z/whb8Fc1ki9dG+ZuT7kdVCeARWe9CqCfonRA6ABVN4fwzwMUgjxZVMmoZbIDaRY
pdCEgUmQ0ZPc9wMa/irr6RnwKJgNPYCyY2QRV4ioNlpHdqsPFGsx+dQ4o6iQ+jZ4
i9pz4XHbAOElN8gS3CrSne0E4JqaNuHQDDWwSmwhAuwXI5Ehmfh0t+iIVvgcUF5i
d++C9XWqtEadgcjjEaJI6iuEddok5q3/BWxbb2Pc5o8WLY0K6BKiOTL78dsVQjth
izx+qHAF0tOXvgQmNqoG5PsHY6i0UypmgOUdAmMbyzvC6/OkfHSzjoEc1nN6ef/Z
Z+1DrMXF02DYsWnRcMiFzQ5vgVdW99dHtHGGlE64cofzfq1pAkW7PbEM/4LT1hyq
fnlGRifCkXBXlohEne5mbe/sol9NyzpzAJeimK1wXPAXhoD9Zi/vArvxeKsJo0GZ
vrDD+IE+EG8R9x7IoWMWY1MQw6XdUANeGPupcVNYO/hTvJgk9n2HW//XlPZAlQRU
/hUQVlRRcMXkfUCjMGUsvxQWrLTwjaj+uQKW82L5zb5FUcdbfPy5kSUUh9eU22qe
w1sSwtRs/gPN7sR1Q0dkc4bBzNe4orpBDibEIckqli12rrrn2sRFPMolpBCYHiUV
B+cTu/hBSP/A/WrHr6jMaTlCmc2xSXEsR1qnu1S20cPeRBeaem4lRfv1G5W3eawe
7LF6U3cluD0Ke/OUyRDKWsC2LnYgftBHooR+WJPhI5hDiwA2KvEglTqleePx6C3u
uKPNE/OBTrQNEJdWNkh8pFehxuFFV/FXkXtqBexSG0K7hNTMmjRRru1SVzMUpVl8
VB0eHmEHR8BfGobgorsQwyD6WP47pTnbvej9mINx8q1noXQK3L62gT28RvKDAcxM
91HNL5gFvkom0EHLVwbgNzYiOQeBC2FCai9nLMukTD6XP0F4pHbXa7ofVZK3G0jL
YaedexbHpAuLDoU0DTHHochxthsZ9mEHpH92bdLQZRIhk2WY0dgkW2WzloMV3QeN
SF+xTrPOTm1/q2a+vD+7N+K4OYNnVrXLLChwKp9ssA5MnSqPhHoRZZqReIhO8MNF
afvltcYlfuJSvbTDYge0E4DBqvAHM6KShgXeADA7R16MbRuPLWpLfEC+6B8zPazx
KelOC6vH+8vpcrUp+P7PeM5s0C4C/+R0zuRuaBAzuPsBjAR7sGglMRPotOeGiOnl
cqm8jWsCqfY8yyFQWb5FaXP0Z0oXjAtQ6iuT44WRuS7gJ8YokKXo9qRoqVko1OnZ
0rQqjzo9Rvose3TPAugokPBZfxlqQvOaN/7SNBJImkuRJV/o4xFkDcnymMWQWnQV
aMC5sEyWRlG3wonqik5Sj5zxEpIYyMuckEwZFrZ/HZRlYbueuDHzdeMn1aHh6twr
3stvk3JrDKDzk10UFC6NZ1ym7fhWe2e+KzFM0mn1TvJPpLumSfV6c7UxK/3tMRRp
IISGtz1nt60WDBZB4sNpPFCXD1n1vUenJL8UOjg5vc1Jr8Z2PPu0tjFm4v+B/KCt
v4G1ZUOLVBataxxCmP35lWHDVXHuflqjK/FXRSEblrDNFullPuHCe5VfkB0dendh
IGHXnzcZXEv2tETCeD7OkaaMyd44XWLqT7my1gt3s+OJTi7uJVz+fdwfaYJHukhC
/oJ/H4Fk+fa6FqKNhGkn0ZOui7+k6uKOsfdgLJy89OpxJvkFVYqqrlTePI3i4EAl
2tk5MP5G0SiLayg2ID8Ok5lUBZyHvYiMz+63cVZqMkk75kj+U7zzU1Q61mytYUI3
K2doSRz8eaQ/yFVba9ZImmMmJ9HIuTE9558OSicLwpRq5win0hpvN1XoJnw4h3zm
am+WcfrGB9aaHCyJboUS/kgceYEaAlk/1w5CZqsYx3JrytmWy40HSfj5ppoqaMgr
Z9HE6mV6JbKBVXxWN4qEom9tG//jJtOAEwLrp88hIN4vs3bnUleGiuiVJoxBHttQ
IrvKB+vrITB0cf/iXdUcRHeYZvdByO0jxuJPW6CXpJNx0f+2ukytu8ppUQH/s3Km
1hZ5ATRPNBPQe04Fy0r8kI74tikEvddTEBt9nzdjOtilMcXP9Mbt6n8vgmqQ/GqS
MSmPPtxLFRe0RmLJrM9gdH+/DkX84pNfNNVcNxABUdIMRCtsI9ktU6AYOBFHHHoc
bJXzkLzNEuGXYWJiKi/Ro8Nl5auwl5Wp6VJ8x0K0NfJh5TSRWFiujWTaloD32Z4+
BRuac+nCgNK/3xMMdpGNXvVBY7zI3Fp0+WzSi34qtytfac5y1ulOwfxjVxhko3Qd
qmkTrsS5JCFnzuAGLbyHA77j6q68iOPMJIsxGy/BIVPJ4/pO9cctWbyKA5uEb0eY
66g12yuSucvCYF6mPqSXoLGNn94j6T+UAuRHNYXYsxNBUzeuoXUOD+ID1oq0G2Cu
vBJ7kHgqBh38pninAxSshdoTDREEYWY7Tk+ywsPzMBrDlg7p4uuRIOpBSE3vfPpO
0NqP6WqvpR86c+hnLeByQIyUL0R0q7iRdaMgJ6pxYdsDSWcmD6SJlZcXZnPu0iIH
qNKBduLGMs2GR7yPjrySdiiLL4DuKQVCASa5mUEREPFShjrT3HGen+FVeUj4SxKk
+NdoCOGbVkeyPd2D+1qFT9FAHafSCb78umAdx3HZjdAVuCATt3sG8IoJiSpeUjai
/ZV/NwEp8sf/tA7a7EG6JQkIvEUaNmb6c+08wS3bqL1qio7CP7RRz8GbhlfwsADO
qxWapzPjar7bTfoWWNV/r+RkRMrm2G3+XH6FijKdikTykSw9lGen4VhJXaEqADod
oDLVYFCHtts+IOB9ep/w+6j3GWWtOe/vrAiLO93DSOznODJFCAtIq+JzXAvIE0eM
XmDeQSd44qBO5e7Wt3u1OMLDqXwuBEfPht6GFXbCumoyHM3ojOL2g5KIJ9t5DOqk
AvwbbzWKW3v6SEoMEWmoSSZ/CJdEE0td2szMbZuaDLtZb5gz1zchRX3D1x+oS9IA
4dsJfork29w7DBFhqZipIKTOo6z2o6jl3jDOPog6KDx75wltRwx84gmRgBIedS2+
nWz9AhCXP+b8zRZNSbUQD04pQjRB7MNPSJEQFRa+D+Jfkz8jID53HS96fA0MAQla
FSVZmZQeZQlAOMXU6DLfr8PidIf6nUVWXjdnzW6tpzcs8hX41JdsHDvgEJz8tddU
nwSKCswlkND7yRhS4PXFoMJor+7/HcNiaCCqQCj/FmLQSyuVtzmcSRY4rxTq0gis
uIPQ7wG35DxhmHvSgdJSg1mLVRqB1/plFZEKMT1dLYNKwtuLyqOqLr+M241Otrko
vh4t3X32ugp3x+mJFI+proIlDEi30nmjz+B0/OIgKL0nK9QY0/3B946LWj/fWrii
v0uqeD6yKq9rt0emhyEZSPvyB9tDlAW16tskxpWKchVLtjnysDRh4ys0Q/CVWUjO
pVfMJB/lUp498xDUrwbQY8KsCBFHyKKJ67e2cmz0Mm0O+6KuKFRy/7SMgBo1cQFE
xlbEIxWizD3sIv8UXQwqIHbNqy5IIUDPqUFp8zf/q1z7450SAjUV7K88atsaEK44
aBBZ6u/56uxY4OD4rRbgzK9/LqFpNxt3wJIDdZcM0yh/JzhBhBR04eSnpxZ/MkBR
4q5KRYbs0p5vdsB/VUj7SuhaLHcs1epsbqlBov7npMMgrttsK0JFQtcTf4kTIvTR
ba9CNQyCEpJj7ykQEtgLK9/qr6Ei1nbiykP68E+MBK9eQVB+3x42sZk/BtRT2Jyn
nyaXiCN3069OP+gTrc2K1DAOqpqLet0akQGkChHrPGcizcDCNXP81Fd284qme34x
QfsSINiW4hY9YvstOXshvaFFJ3CLPck1tyu7jW/jRUK6gjlrMSle4GxLXsWa49tJ
6L/UEhkL4gSov7s1e3etk5NEPlw3VWEHuS8ZDaGeVKl9DYBwn1Ygtl+7SO/E0yfH
SakaqH4ZDhe5uHCFgqwocwdmoLliq2ab5NM5SGfuVvxt+RwDNEYGXiCFK83eRxZQ
dHtfPVsuqvUA5Y1aQJlIFz6QYXSA6FG81D/yUXuq/LoQ4pu5fEC2Ur2uzeIC/v3v
y9ofGZ2t4EzqRiEf6XAr2AqBaa7UxUIt8Q8rMfn4+OltY35tYygrffhWt62WaofP
/6KkgeMpze6v+qCR2I+zt9unRJP5PzI1KbAKyD2wbEW2K1ugZ3barqYRvWQTGOeP
C/Zr7fB5PVXdLSIzKlvQZwmsrlzAvNe2Bub0v0XFBq0=
`protect END_PROTECTED
