`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rrzVFIVO6w9jQ2ScUt2aNn32Vn33yCv3JduyMbjl/DJAC7eRUsMIEnprrDNulNaA
vT/B4l+LuXIn72Vxc3YK1b9Ab78NdWQp7vTqiHVQ1CJajpEkTI+KQYnTP63OPvgB
+BcU36Zs2VZedbhHl459spAAeh1y8T1Tt6iAIqpWqeHSf+xkhuKWlQj1eRx+qSCv
BMdWE0x4QOkrU/18JujXdoDCyJ9yF8q39p5CqhtsPOoHXa0uXPNknnGDUK7Gkue9
LpiBnkTRyzu/yNifqkgufqkLzlBafK78SGdne5JhRq+lvorR3YddinC5lycKCJ3o
Q6lncSjaUubC+qK5d9nnUQ==
`protect END_PROTECTED
