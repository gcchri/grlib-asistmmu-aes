`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2QvU+1IFh7M/mrDW0xuvQ5kqOOQFzdGtN8Xw15PX2eeiqL7EXYx9ueldZKM6Wssf
HLry3Ih31hfa4pMfqra784McjVJKUE6dTti4tZ1pPghXdy4e8GoKA59P1p7YSVu5
GfJPnuuqZIBmKNQYlYmrB+nVtaEy5cFoFLkT+pWhAaR48jpMjDJciAZGAZiGbbRj
6WwZ6uX3ZWS3GJL83lgeaEL7u2jAmdzGG1dU7Deq0o9e3b52i9ivdoxVB4+iSEeG
zc8jHd4LPTgJlpyjeDt0pNgT7DtI9X9ZgxuM7P3oQa5IFHu99aulzTxvUSsTPcUY
kRiJdyOkVhqDeMWh5FV5LMdekLthV2ssYxG+zF/ImrphQP2AO6TYcEqTZEo/UA2C
zVOwgCYMPN34f6W0xhCqEtQyMLYCo9i7hpsBEzOlCJrgMMa593fnbXYmGIUSXWtp
DvqCwdfWR/X1zAqKtXdGzRhKTrmJQjoTBMZEThO3wG6BQYlW5bGnj8/8AUxXWXtu
fpXxH+2BWi4i51NdRfLXSlHbd37wS0Me5jzh8q7S+Q0+EbjCw9Vex/1Ps3uFy56o
Ih5v1MmR74yOxKsrGNQ3DB6VhjKAkIv01HWYglgieYM=
`protect END_PROTECTED
