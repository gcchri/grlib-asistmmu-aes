`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HGErmBOUZ00asMKu/WZaaPGHrJ1ysoQqYQt3PlMu2PmwLHU6fI/m5pAo+fVJPJJp
ysVSGefMXaK5TfVPi7w51cdu1wm0sWWkWj8H4M22AmLjyIduC0YxhMGYqrBI32zS
p907CdxbXvrSO1skY32O731zbmJzMyPaF7gTi9W0AJHK1KW43PbEAVZ/Cs+Q3XiC
mVv+QJJ/BfPPLDCEwZCVMzWBLNkLuiTOz82rZ9TKn25SaHao6vcLUjNfmEygRo/8
NiQs19uTMn0AaA6ZLKbZmevbpXJKFh/TKv5BLZtfN9LorotujSw80RcKriq5ZP43
6i3BZafBGXin0yyPvpbwzQnBsvKepDgfoJjP0GEAFTMmnKy4zzpIEk/M8zj0SWXJ
EgYuol+10foK0SuctWie6B6VXCEod6zvdma05Hd4WhaXxoUmXBJqSThr+HJJwRDz
pGayQL4WaFUJzfYKfOBK5LXBwSgW2PnKnu+AGXXcFEB1f2Rtz1jS10xIDyEC2MSm
giMhqC5t+d7YHtYH2HiX76grL44Vhk4cxeC8egBTK4wCWrZ9VDjIDaGZWgG8h6SZ
zPViuIQscB5KUHNgCz7qnxW65QO1UOwD/9Ep3YVH59+me8M3dK6JHh501xkMCWdr
KzkGqb1+DWv5PYtGRcPrNP8cdc86+A1O6oaigJmACa8=
`protect END_PROTECTED
