`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ODT/+9zVlY1YEPstyktnws6QsHXEsmu1GQ4T24Fgp36DFWxk1U6uwhGuRSjorZCn
YHelrPWGM1nqJoxasBq2d8oSgHHMLbzR2ol7kMwd4Cx7Tgo11OwmkDosljJIeEOn
Or2uu78o0c2QJG8fLDISe8UzvLAfq4WrpcBVwsU/glWMc1EUsOVovSpyyD+ngu3g
f/Ga2CX1JhqT6r/dqY6O+Q3YCT2HchBzXE/1BkYcCGB6o1smNezuzE9hDX4EXfD7
rStGD7PioAB4GtTlotQQ3E1GqnlqZZ8m6OBAQc0iOOXXySLZa2iqRVj1xr2OSiZb
0QYF6Rm+4VS1Z4qbG/q6ZHtaiHZF9ZkdL2Y0vPe+hK1K8nUFr+dc4RcQb30Rt3uQ
b2E1J8w0w57FT76XZOtDhL6PC8sF8TpRirsk0Wk47vrvxXGuJ3AvLZoMHpWFTt6D
YA+3HpWgF40Fth6YXVgoX1skoJMC/wTBPxo2bQfnhH+MWZXfONwOj0z9qertQolw
nVvsdveufre+y/DQgh0J7COcADaQ1TSdaYHeQIdJ6bnD782c1lKld+nLuTomD9DA
5qfSsgHsHUlVqRntAQWDC9ax2uQ8YPzneYCq0XHVCpP8u3S0QsnkuJcornoMQxsw
+uEFvm1VCTTLJMoHw5KDkEVsAVdxq2SnySi5HLItwEpURswjuTZeW+OjGKUS5lVu
s3LuZAwSW46BvGU3kkjr7XSu7irOVwzRV+M7XCVopV/8Hun7BEIWa8CpoM1kPIy3
S+DeXFw0Khc8mS0cqdoonA==
`protect END_PROTECTED
