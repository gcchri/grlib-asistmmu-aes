`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mZ2s1BqvMhrmd/RZp/wwvHLR7ZcKZJIlsinj8FS/O1qVlrevnztdxTy+3zgghvH/
dxouOAI6SxslVZXDZ+G+td78A6PM/hx+hJCr1B7hKuetJUDDqbVyFbNRPzOB4P+k
e/N3JSnwGL8gvP2CYozYXnOeWSRkEMsxSwJ6DMpGOExC8560Rb8Niy62bJlLUJGq
7psDsBDOVVLLSw5rCXT6MXvReEepKbcaS6j14JN723fufF62e1AnmwA6Gw8UHu1W
Pii1UuptJb5uCZcXmfji2e/ghiLjX1AFd1bVJGFtZ5EuQ8wkn/n3U9Zax1IIVlZP
DaL3Gy3hyt2+jXsJkW3s0fUivIx8f2pYWN0NeE60i+F/ktbMxVyHyzlgalEaAvDt
KeILXGlc5La7+zXS0iWvmwPOm0N2i+igqioA5lfnAVm6MB1esHl7XxqsHh7Lkn22
9aPKShBLo7Lf8YNxYL8xI33tjm95bjI/HuQlFwPI2VyLTOGoOCA3BplOS2y4X1QP
`protect END_PROTECTED
