`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HiJ6j6dQCZUL9fe+WN/Ugxz4T4OK5S5eqscr+wTU1DjXAT+W+yNkA060gusrj1mn
THO7FOG9t2VcZyPI8P5la6E/LFSVZxLInomEslS7xAP4iRJgaJAWKfg4BELHRguq
zYSxtpwKY6AMiyGFix/0l4cPbsz4WMk9tMJ011KlhNHoxvSd0mZZQr5M1o9oIRJl
iQeCI2jYFtfZMiiqdJpKRwybqzRKbmVNhs5OiBQGCHY6Sn+l/9shwgKSPOAo2P/v
qwYnoIdJywpHtDv88YfUQvrmWRtVMO0ehUOlx6jWq6RIrGsxbexUYRES5OEotAQq
quY08aU3v6bZmU+oLcWTHi2kC1LDGuPeyfBqswdpr5foEdKS4ZOynDo8KhwfgcVG
NCrwaED4vIiQ3fRTTP+bfJfTNf4ABrI4jbJpeuAUDOMwwSqnDUb6MPTO578canR4
jOzLZU7LC5gKRa25btoJoQpEIIcI35GrjmuHeomtVEiSw7D+VClyRNILQGv6f8d3
0xuTikVYPkuIkJC/1TGujzguFDsxSVk5k10opem6qrjHWB3NfxlsZbiBUZTvWo8p
3Zs8JG5HXh2cZupByO/dPzeIh7RyMPL3YS93QK++Bc0nZ4hlI7zkj/pjto0YIxO7
Rj0edNAxPdf+kydoP/j/rvy75dOXV3bOpBpEqi7p67/La9dgcOkUOZpBMLCcZswe
z4u92TXprokCoT+6Q+GkR9rUgklnD6Avmwy719LUUBva0yyjTf7hexjZsFFJtl4N
ueE+4Vv+2vz2bPE8IOiM9sW9VcEj+frBXDx9z7IXbhXMnOi2joLSF9iM2Zdn0LSB
ZQYZ3lzbR2E1rge9Kl4Koh1T9jJs6IqhRcBPfUCX+vtSkOhPffdjCiArbl9PHGnk
sx+LzAzJz2xqalmAfF4pFAc21C4UqJwmStAJeGV1Z6Cp4HUwsogmsPGB7w4ZXESQ
zJNUcw7evk2ySf/OkfhZp2VsegK1DmufrMKOSkEsjQIROPMyIiJoRCn3hPwRG7ze
0Y/0qyo933e81AArhcBeVf6qgU9KQdtFZXHBhmkjv33fKKPQtSnbyCkeDo5+QtdS
5ilyRHIU+QVH6HrNs0OQJ+ziRLkqcC2J4upi1pN/NSy6EzPGjvDkKcla6t0it5CK
A/xyc/colgumpnxwc2HDE070yD1i+e+Bv8pa2qHVQIv69n38c2WdAS+1vUUfwjCM
P5TdiR6ESdu1e2+6BC6akAajIn5UY6m88qRGhbsivw4jNyK7aRbfH1xALHCLNZuX
t2pS8+tgQn3e9oIz1EnMBfDCrZvmiCwOVTGzL5Jbyk0XVuBlhZjkNBW4nurtXqZ7
Q8NUKBrvaBtPMk+EjCgWHj8oelwByy/iWWc5komVn51U+Tp+Y9L4KHZUNCy6HP3e
NaMZLstb2x6IIIhvfbgTlHxZAOObbFXCkfA+klDc+/7W2ScZyz5rA3jQzcnB7/v6
aTWgSGnfAaFxdRhIr43KmlvwzkyDi4bqGKqgjjI9KJWvDNpGsWjKphHprJPdNz8m
n4EmmfAbQZe5Yhm9DoHwTWdxbZbLrdSCoqnrUCFi/kuHaYIb6iu1hwUaz7Ui3C8D
ThY4Yi/AXzRM2eRtRSX92UtblgmDRcF/RYJcbOwRjakNkm3JWadURQOD8rCFyvq2
8sCDuZfKcQ+0tGg0+fNHtmfGKkdEpnX5QUKyeAI3KqHxr/gm3i872N7J6Y/7sgwT
nK/uBupDHJVrWQRL3ZhLv5BoL1eu88rj/QKLh/I4L2MhxD8vFXMgSPfHe6Y5zXoF
VXBAJSY3RSo0IGhFfUY4qlvcuhvWu0NaQwLo8bCYZqctXS+AkKVScTFYvuJA19cP
2HGfBJmZSezZLcPJoRS1JyVuKGIWMzZNPkmeZkDoikOwqvEC/z5otSvFySGdOaIf
bCNdFLGtJCxY9dgYtORhKtNz1U3a3aDewiCgPdsSFGweAfYBM7flkRmIY4GZCkyU
TFj015MTW/Bjp1R5EN1xw8vdUkjFV+KdwHZzpZQPRfvw3vtsYM8Bc4bwamBYsuP8
9gEYDcyIbBWCnRDJMGZgR3OL3r6tRl8xSYSgayiGwk0e0UzRbUirDR2W5VuTSQYs
I6sIRblXCiloeJ8vWDHT8QRCde01zNvXFQI6L8s43yl9cstY2/Q5QvWzi6lRagn+
fv5XIwfiN/KkeN4brzXkRL73+6h5j8JEFyhspnsln4/7aoxaeC+EExQRk3NArZX0
qrzBiNXo5LZ5gRjN8Lc1zspLdOxP7toDJ8SCb6lh4/Jr/Pv4rovkE4W0lD+FWlr7
o8r8FNQcmAm9FfyMH99+yU2BKDB75neehga2J54fk8y09KXbetF9erEncM4SWDfd
RpHfs5BxNRjDp8VguOxJqotEbjSMtBq3SUnSuliBqIbFn1qt20oTckbwnqs23Rm/
/EN42qScIHQ3UL9DQoKkmux/q1O/6Wze7KbUTXNlxOOOlp0jz2i0+RO7tmG3odBQ
VFkqwu5GZFhFeDVsYu9764adEQbiPjWh+HxTHvN6tRpgNRxK/jPGtRX439Eu7RWz
Jx/YeqO7tTs0cAUtNGPbA+h9NdIRUyb5VCvU7pMPaSyCNXMncLzulljdtn0rixhd
aa2vprhEqkbxmn+1bTShdzEM281yJ3yQ2w4i0jdyhEnijELeVVxa/oocsNLzTwNK
NnmCnHQICOMVEVXYoFB6xP7eWye1aAjZxTNyaTe+TpzW8eyR3WLbbWHmgvpvV1uB
zNuD99lvz5JQ/z/EjqWV8WDSIMIuNJ/Y2z38+O11OhZdy+shMvSCez5KSJ8lmj8N
90gcwHlZqEWrm9i3jqd7j/NIuHjQ3Z+5QQ0l8oN3Ps68Y/jpeMrYJ8L0hNDsGl6p
eV2W5S1YUJZWqki7TA8vJjarF7XOhJP5TVb1/5PlJr58/brb3aRfHTeJ9jc5i4v5
dZeqa7sKfvu008TGwWc7RIY6NE/8JXn2KFlr6ILbFEKQNbXrrfT4Ozc0OAvM9cas
OTprfanYsgG/gZL7LTUDIlpRTEVJc2tQiRb1vXHtnwbLd0doIrpplLIiKhoqpcuR
0Gq2FtEJwItAA21IlkOVBkEcwyzwiwlYt34ssH+QhZgrxK8/SK4A4iOijfcaP5Gr
rEjeWukV7h+/Cxj2QulvzxD7hd0K1/cp3kJwTxg77VbhEr0VAwNve4ttKGdqnETE
W6OId0v97Xjw967U/BHPKAVNtc3brGNNf0QUpxaxIaBUOOpt1kA4j+cqOU11pHYL
cND5y06OQhZcmgGRJlLwoyjyfXK3Kk1Ix8J2/YOgEmJTeYN8m70/Dpj2rLXTdbMA
EWWSuJaFF448wIjJ8ykNIw1z+ltHXBM0yHDxHRbqpyIZMFN2mSutXIkJI1dQq9H4
NK2zY4E+IbKQGirbtWwbOoX3tPiMih+tFW6HSJWlM0f6ipFk+fweZYMiX7/48TnA
i4dEPhJIuhdu5LEdk5o9px3jRgFSn7uhY3VnvS0LM/ETk8r5HCdH1Dlp1TI3+PG8
/hwAH1HIvPZBQl/u6R44FRsZxOPOl8eQEDDIL7/b3DyJaAo2fmUfTkQenODa5hXf
SJpHzfbiUGTbCJaIsvNP4RHVqADJ16ZtaCKDTMSbDag8NAwBJffUJTp3avoQJSEx
cQkd1EgST4CyYrd1iLV90Y2JUhEqBzqt4FDF/CtWJdLkSu5hamF9heUxhTJsmOYD
AIo85OSZfUaB37J78TtXuPZCOjX9vVPs3aIbTFlyorFZrhBzlyXvn4ZWcb5/bRmX
GhRPCKQmTtMTRgL8FEnjeuogz67orDgaVSdr5QGdSgeGW6H3vVFW2L0Z24RjJdUG
l6uN1uDULH5YRstCtflJgkIYOTHgksnLZe0QBJHcZoBynV3YqXaVcuNIgc4JqlpA
hGqqietco1i6h8VTyAQ6rE4hvDEir6Q7mV+3V3O29cOeEfzWFozKlewmO007QM8n
dZo3jjerZxIVMxnFWNqKrqRAYhzc4pbcjWavtR9seeXqkbkxbM94Czt3uWp4pVsM
FiboLbq+SuTur94L8U9Gwy7pnjCBc2DLWY8VdELJNj6whmEhz3cEHSkwQRfA7MSm
DD6NByHIQsPYG5jqSm9e0oMTPrc9bmjSNiwnWRJHf1aSVZ1hd5CziL+G4QyYdv1u
FkIRNQaLPvUYcM8v2ciaasIDUlKMnsvupmV96XQeFSpLz+DzSzvKbo5GzYnndLwS
oe1gHDWLCClBeuXYovMzCtlt0an/eQuNnrRcEe1wwuPNaCjcBTjGgfH5dUxxtaVd
oDcinam2oGjxw1/Ge1m4HP1e/cSVDNpwTcNjrq0i3gNDa4UJSGKF+3FD2LUXde+u
+aFh8h2NCjsb1Pwz9glu2dmp55md/8bECwpclARUt1xEir4f68o9ch6vb13VLVLx
zo50B5HKomRhevEv9d4ZBCocNCJo5nNhGZoEfLOJU3OKpSHw/aTgcpqhsrGe22RZ
p0jboljBz1EUJKw8umc9wSvg+kdF+1ixGOsfZiLftkbTVoT4A02AnR5iK8Th3IDU
UsTLakVOT55YHJ4QNkkZ7DpMBMm1I99feZayvveuetQ=
`protect END_PROTECTED
