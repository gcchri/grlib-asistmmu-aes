`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OygOycXkAEwgJOkgOkaYUiJez2Y1zGa/B8I9u2CzIa7w6uMDvkVbnLud0IRoIbJs
R22NjOqYwuRpDSkh6Yn+PyL+WXQTZCp1y5U2fShKiKFC5EkCOJyPPdQNi0VLm9bo
5xDH6GduZ2dloTReJ8UOdOGwcorOT72HT4APz8mpEjQb69ssjt8P4TEHtJapXKH8
7kWNVPXt8S35blFuje4BJ2DgaI5XM7f2BAnipB22ty+X0TMy3Dcfrt3Jc11oxpw2
bMF/geaj76pe4/3f52hIFXLLKQYma7JLFMbyf+/6N1EOhTKScuSgNjeQcXYN7m6z
c7FK82eqeDmKHbaoRw4MUZMuzreys4MG05hqSjw+IIqV7hg9+MBMtGANgb121gRc
+Qt4POd/zSWFkz3xuT7hzbC4XgX+4oY0EHD1RGxrnRt62Z88kw+nGcRkUP8k8QEM
`protect END_PROTECTED
