`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OOGJOxg+4bq59TzHTPNtB//jnAeroDuomyK6NOPPTgyUHvG4VP+i5E+aWcYTpiQt
cnOuekk8K11ITSLamTBYWpaa3H6daQwHleHJtXdWrM2gZWIJoMtrBBubdsiOMVFG
4ue/jLVRMAlu4fO1aouTb5OWIK0WSlrvrzj9eIJRar33cBRe4aya7rCoqeBCfTVp
8EkTyZINSdsXvQs0tqhKoooKl1OERbF/2qIxsqFEi3qGPPSoXxMz8tmF5fCzdJT6
HXje8E96LJgTZOt4MxIlg36UnywzqO0GPPDIloba57K1lzW0CYS1C9xWB09zD2KO
O+KoA4dk6TW2s4CYvAGk1XRf6qDmseNcj30ccWJC5k/PN+uDVomMwZRsZ/s4/UCV
w2WAiF/KsT10Ei7r3HL5wqRS8f/ii7gVoX65DxivcHkzNNx6uQFNt+5WrJ/l6meK
Q0b88nhSG6cJYRIOof3ATAd0fZQlWwwc/Fz5iquwm/CHsFqQICbYAzvfybxeW7NP
niurUo9WmYc5lji1wmlSddjLaFJjllAlScdabkABUZh91u5y+mEJHouLLSy1OsvG
q1BFW44p90lBvtJKlHS1PJ/Xnz/GfNMuSG+cTcCtyG8=
`protect END_PROTECTED
