`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/i6oRKxxyGKvAOHqP+z3gFTaAkR3++KlC8vm0NKb+8I1p09lAdq+PgncPENtxU3c
lg7dOxgdYhEpj4g+Z3rxfYR+qk8muXBBNRR4vkmTeJcoqWsLirlYTas+PdfFE1u1
eK+rU2HcNvQDjNa+7YQyZS+X/5sKHJctty7MmRm4ac1vXFW6DGbYDOKUej3cVZfQ
uTIw3gNteBITYk5hoB+Bba7uRWDbDiyRyMZzKA652PE9bZFXY0w9D+nTfo52r+1W
U1A7KFo4tNoQn5ziP44eDIathruRvpZAKMb4RnWF/3b5rRVs3YHFM1aS1dYoCQwB
bV7O/gH1hGxoNEhbxYN/eFUgp2rm+D6oTCIMUbRHh2cB9PKjs6R7si2MhBs0p424
ddqlTXayIqfQtbq3QDK07wQ5np5arjMSMqYwjuWfdaSSK5gpLjSkieatkH14CNnh
1w6qhvGYnvyT8KlJO/J4D7HbRjHsFo3SBIibrzbZdd/EbvCBvzCTpjsLE6CO6uV3
zt89o6LBjBBJ3bT05y6oBee6Q9rBxKsnpNnDDB8zwqAadez2ZXdK3EdjOs6dVfSp
StbkQvWydk5Jk2Beoq1iTrvkJik7UEs+gBkX1E8cwzdK7aomta/zVXJf89JG0tTM
OXW1YtYa/GmZ7qVpMHQRQt98PNJAzv8zRVap3eJxfGc=
`protect END_PROTECTED
