`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O74ZWtGHkwfu4M8xx+nFTbexdNX81jdBpQSqxg3ERzcD10KavK+uPqSmmAu0EA8t
q/AM9LKr2bKwF1G0/tfs03WNCeDWYl7Cl6hdIwc57p6pvviUXcg6Z6StZufyG2Qx
TmMRrYjFpCMak29R8UFoOkZ67Z5hkitGyP93Yui8JRaBHODM/bmsYIWwhlUrs4Vx
D1UZ/ao9ZHRxLOsthkxu0RaKg55B/1j10Q+L0FxGd11WypO0PPYWdvhDeLx6Ukk7
/rDexNir7j8DljRUs1KWUzG2wdwTpZk28Wkz0fobTBEjM50/RX4verLsxUarr2eE
/kMlZ1noYfFFrB/8M28iR4UWKJyaSTd4+mKfnv4XZXdt5XFbCPu3lnZaaguyQzaV
VQCuIkidlXaB/r2Uz5XrC5TsMAGgxBoXBAmLal+mFT+280pdF5/GYEkGziztLtpw
unyBVdHRvKIsoR2B3jHPa0XE54nRra+DORLgjiM1rMidf3NMSK2gobkEqYVrTeem
FfJpc1RlMSsKu9SB7Tk4mdDstnRChTeHDZCCEL43BIqDwuy3V/JRa/Mrrj7D7ZBc
7GeOVQXFTer4goGKbGeL5KO9Opi+wuCrruUB04GKpnFiQ4Zo90Yz7FNiCK4BcaJz
ZMyXq2izCAQFfi1hgkHMXDt+n4FIOEe/tij0jiRl9AxT+wSJFx6RrXpn9BjTiDp3
Ksq/De61LWmNbojS+Kkdyw38fquNtt5CT2ygCA69U8x9vSQcJh4ja8bqG7l9HNfa
lrZclOEVAOwbHN0NIYfSJmJMKjdn9GVf62VgGeD6BxDJJZSRHKACTxzgRvnV7C8V
z+FPQJIFdDUmvz/W7JTJGbI8zRp9+Ufp0XC7orKIKBQ=
`protect END_PROTECTED
