`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4IchAQLG4ul2Uia/6JNjIwPK1y9oHy07oQBbvvEhQ7aWE4rYvlAHI2bbffmr4tyF
wRGAgT0KnwYXdKKOQN94b9BVwz5F0o3lxMgdYTDsHPkR6ViqvYz5merKYOPNjhxN
rjQb6BeOXkAw5ibP+onFuX953t+x0PCLW9ddqNNEB2X0fFaeeX04T9vKIlzM4duc
3Gbgr0If5bLInhL7H44vitqpg71unl0hZaCzTDGG5ParbVArStyThULo60Gd+SmL
yP9F+c4WLb9sQPPn7DCmVMBZ7QtsMFtk3qutdXYt2UY/dEszurgq0gAG+WgJmwne
U7eR0PCNDw6m4DB4JhvNOobNkPLHcVEGe3u2h3C16EaCr6dRkJ8GHpBe06ypo+cY
Dyz13LoR4Sx/jNLzsGxLy/kW8pkgrkOYqz7icEZZMukVumvapKfUxjTO8vd4rxGo
7odijkaQxFOnq3lnoncdR4ygMgoHo+srMtnrZgctJzgE9i8sa7apca2j7Wo94kGR
HNtNvDgpxMI/QBs6V7DNOGkXQDRnE9KumWbpw+FCopFnQSrsmlNXHyB+H+mWO8RJ
CryyjIGa4oXeI76EtlrDmDe/2KCqn1idZwiG/lTiDD0ONYG/m6FrhajgxAkxqtBz
4CgYg9LoQ4kboTFD73DN3AIiQ3B7SGdTqm+BZ3+5aC6ZDeavP4OrrZbLul/e2b0H
+6v4lkFpIigVQWnGyvB+Op7K3cNz4s/68jdvkY3VJtQYVw54EfemWAzsmpG4UzIr
wQ1oBGijqoJTWeq2Rh6x87SkCgekBT+qA+RfgsjXNnFt323t2RjWWK0iptBhvXJ3
CTa4eRecyuHGt720KJcm6EMSWHTS501ngVAzy1kPv+rOwGGXCFwPJ8FK46CVCuSY
+UeEQAHyPG+AOFhNIWEGD829sfVysKtLvWoJNm1YYHsZ/ECaGqfIkS7j8IqTbP2I
/GYKlKzoMAkevdpsfJu2FcBHxnxPw3xoF4+L134KXK5AgsTRgCmm5PD2KDFXJGrk
Ab8RxY04prGizfZZf0RJHKGzhX5KJagP1bWj3HnFUmDzni3xHL8vRWLPw/ga2Oxs
BjWDYJlhBna8asNLulT6oUMKHwMoXu6QXjOkS7XD5XlW0G0g3ifkvM2o0oyO7knC
xvM2RI4yZyNsJ2M4g7kGVRyCKat0O6UPF6ry8VsDqFxrsH9YsY63NWLBcqmqoWND
EWdvccpCT3jtQ4cOVZ9rFAyB3i9FDTFTDJXaljG2m+GCsZL8WDmpRUWbszA5i1/a
fDNKIQGawJ3Gd1tCU/CgzWut3dqM6QhXrTRiY4vIW/u6BTK8j4CzKvkJnQoOBl1u
fIV7ztCjWT5Gcs9XTHMFsWA6bpryRaDRyxUfjALTmP0vR5jp/sRpWX1LTRW4J9bb
5gGm8yALDx2Ah/FXirjZ/zBOQsucW4rlMULChobc912ty23N2nBREk2SCk8qeCQG
cdDl9RD/FB5pxvXW1+2g1CViJ6QShoZNGeIr6b1Hvpzb0Hqc94Tz56GZNJqvvEku
gyJ0Cd324fwXBsBSWCA2rGsY5FTZL9ew1YL8+M/2ZXA8+pcPFHvzB6g7BDEeV0qy
NXgfuzpWlC88JGq/py0uT8pVhUoeWtXRyNVJ+LeoTsXGGsnr94PLV9QLGxO2QWzT
/2zvV2Fg7hdYYJugBu/3oQpZmGvy3USdRYniUkHqwRss8JiwGR5KrSbkZgXpS0UI
nTUxw5jjH4F4VoIp8TgygDh2y9KR+kaX89Zuznu7yMFVxyEuUxAlsZDGCi2m+2Xc
SLa36uDLMssqoKOdehE6BtiXJTGqmcom1l/xgUObkoGYClM9eUm6Ep8zZvDSZF0j
FtSPEUY0KQXRdXashdluz8vphMgTFcOpe0ZBbsqhQIItvgolqAspRz9bpCY+kRkw
OJqQPbzovKfUqMkPGJekqEgvgTulbDkKj+m1eZVvVJBQsfWuiw9tf4e1IKrvZkt4
KadcFZrcD3otlbP6YamGFqbdgFES+RsPhaN+LYiAA+FWIqhCkPUH2S9nM977x4/v
l7MgBnytAYohA0WJwpednCt3z4UpElt0Xms/1wDLM5UV0ObOOpZzVzzmOX3KCU88
8mI8IHuZNoxPZgoRbS425xc+21clBWjs8xkC1XtK74oT5JFfrhQ5LMariq+xJ3qS
74mTT7sCBJCkCLTCvqehcOqmobcraSFIv+6u9lMmyPtTrsc3Y8IFj5pTXvA7dFUA
RWzFLdZx/pMVKr1ktnWoDyu8jSdmZG2HMdGOKoGYPpqlGlOhU3GEIpxRR3vu/LWF
xaPZFwKNfwBN+XQTRcsK9hmQJwJCq/o+0XW+Aij5f/P5a26LIXK7zpFKZBpzBUEw
u7llReJ68zJLKtMtPOOyLTdpgRB2f0wNpGFB3qMLGU0375Pbf8N4ujzgGiA1PFky
XlVw0E57JdeidhpShZa7TcLoWtV1LaZsk7m8J7iR873pGHjAxu9RXsKmbyBRtnYa
wPYx4qIua29gANNfYtP1/ROckMLahWrCGveRi/VcXMxv206xBTBm3xqNo21t6e9z
ShLz2bcBcHuuDtGt4GbLERjLkAEMSzlMIKWYSOe3I1xwJN57nvYfeMSDW+ge4MRa
T3a67kcLwpmcQdbROPvKSCpW8P1swSTczuBgiLRcwfNYkNvnl968q0uzkv2Rh19f
9tHSd5UmBq6YClkrmp7JYKNyqnTBBSuyRQc+O5RQ2whq5YKcz3SVpF7mBO3cVspS
QSaD/fpKWq1/Ctl8FPUNPc2MGo0oDcJWoraK9N+Cy4kpkEWKVdUt3WyrqsMmH15i
8KL73w8ULt0d4sLYdZQXoL3gRSRIC8I3F8lCeqEA6uFA6vkGYSMazbvLjqV/tsMP
G25Gut3Hvo/SP3SxEl9OVhCyT/2lvYwhhtFNHDFxTiyy0X7AA/jyeLX7pVogHF0p
58LXXl57zcENsdiKEbzVdKbjJ0CoTUfo6wPCSAJr2O6Sc+NW52zIHCQyUvyqVbb3
P+/TaFnKec/cYo9USq60fyETmAT9qj5JK7pzgTC/gDgg4yRDFXnV/Wj/eGYMmyn9
m67+x8ALGiOSXKVO0AVm6bz6l3IqVZUiwAwtQhPHCJxEyossnh/A1AxKLmECw7N2
by5J/H6JD3QJcQXP079y9QXWI0E6eC4c5usTlH2d7Mo/9xfAZNHs/eYI4jgz3BGl
wpoQgXpdakcj2hQoOMjARkD636tKCIEx/dJDsd/9Abx3ovgnVcKgiWIVwle4kUBx
DTDlrkP79SprlMXHuiNl0oY6b2DlTyJxFg0Qs/g1ARu5fQTPBk1/7wYOBTBGY8pM
k4nXsvUsLUSvQxnU1eRtFU0wgnVO8iK7qZyb180w8qA0v9Zth46kozJFCySQ4Zfq
ruRcLoHh5m0ZkkrM2NEHmc52MfOK1J/fodjVeioNE8PoYgJDQo07l1CP+wzzP5Hf
Iq83KKDaDTCvQjOjGxiKRjLCJJd/rLMMIrc+iNl26b1w09eO/+HbQnH9kOnimH02
SMHuO/IY0JPy++CdQ1GeSlRU66WCOB399iPATpIz8dKbbZv9OWK4J5dAgBBw0KqP
iduWrnpaLYHpnFyYIHq46In8QiZo1uAOhILlH7I4wEECi9DtvZzAkVDEQRA1xDLG
7pNxgdalbjr3wh6vMrPGvHupITBEP2SgCT/LsZOl0TvvPqYCmt0DAIKdQBlR6MG1
oqQzk0wu5Z2g0JblKJXt9AYWbNQ7GVMbc0f0gWQiuix6+VZ+jQJ56SH8oUeOzVoC
lBya24YwKjiyQDvwVcaUbVSpoOQI8dKDkgH72xNZ3KuH8mnWzC8OPnJHYCE22dqi
dy86Xd8ADaLAPcGeMUMj6J+lD1DGFxh1TF2bFXxwb7vaxLSqg4RMGa7YyK0F9Dsh
V18Hy/m01uA8icCxavRCvVRqKWsUWgF/ul9eaRPcy66ooEpBBZg5zHXxVud4DEYJ
07MqF3Nkxdj6nzKlkkKy4dfnxOOB+YZD5Qyl/mTuMG7p4EMCsL61BTm3n02JpZ8C
5P6GRU2/L4MOSPuORICj4QW0LMWpEXQZuJb/PhTq1oJJM3yIxufiJ0zw79fTaB0d
A7S3a05N4/r8ZHllx1r1Mfie/BM1X8nrD2XJDhJhoXdEnypUkd7tl2NiY9O+5JmR
kX245+tavrOxnIACLIzgnA8e2pGRrJ3a5+/poK8q/L/zp29SGjvzyOcISJYZN0da
3uiR6X/3Wg7rEzUtX1U6GV00LycIThRv4lJhWubSiybSD5vkFvtMNZp1SHulna+i
rakJk4I7zQbjsCjApO4xgRwwg8lSsF6kRsz9G4CpJFuM+dVgmN4OiYcsywjfnJs6
avXMmPt/V3i90NCMw1o0Ig8fKdOO5jt3qUJfAX72kuyn974jx/9ozXC1ehQ11wXo
lLfl4PrGkBz0zbGhQ7DjWK+4jNhgS68ndylEWn8pidrOKtlLFGLb7m/UWjZL2uPJ
RolkvOuIrrXUon4EixyY+Z8PbA8k/a8vFuA64XlcHbYLd8EMi1SLX7cNBoE5MXuu
Q/1rGnQ/zympasJBKTK/eIHtH8d1OU1XWyLFbaaCVRkQ019EOO3aQGVDIvH717HF
/Wl9IfClQDGenNhXXm17k9R0JI8PuHppKtk4cpJB6obXdVzT8PGQ0cOeW595fT6k
ttndbFgxoPEI2zVH55b5owjIOh1yZEkKXZ6jdPltCg0mp0gH/J/f2e0Q3y+AHckh
Tod3QMSB6hTdCAPNCTNBLZgwxigZjGkSJIvhgwjVammlZpLvvcKjxFI36x5ZGBic
Oup7vdjMdR4ePIPe0bivep9tPgn9OX0RN3Azi75J59qJ6bWaSbGZzDDSxKqRGjWD
qekmIRsTCMDbhd1SsA3clRU3nVD4ajR1rD9DqXLfJoIjGiUlZ0q9p5rUXkTKOlJU
2YC6y/5s/JCjMYregqYyBq7lY3OMG63giLCOIsMDwg+dUW2QVzZN7FkKCyZywUvz
ctClXowTFkVdzGMwUG8rzea852tcrOz+4Y+nhBzQOwW4Mh3zfoHdEMPq0dZjUsja
GRgYfRH+nWZu49ACjeUZ4mFlmFaAazoG5OGYsKeihr3y2LsvpWbxxQmAsiTZzPlO
vwovW+wumrVWKvx7S21JTxNaSemRIDLHvoOhYiUhZ75fEs754UeZEF/AzK7FZDih
U1TEJqbGyEtbF9XGtX/j2sbGrhkkkUQrMc2r1ETDxY0AfiwgBIfgeVds0QtawbKP
HjeFTWtsKRTZBkAtBpoflI+QelhH0ldyoC46Yuku1e1eQnlZBj8rrLNIAYwOQMrC
x2vF8q4bs+K+9P+Z6k4v6bFKpIg9rtNFzvPT4hk9VukW5qGNKN1Kw2MOKf0wZIVt
Le83UMedjj+iteJl7Pbzr+OKCSZwiYk/d42knv+siYDt+voV/pFNELrZw+TtyZul
2uFw/Ibn5BPijHh60AzDzJQL+AQZfh9+4fwG34FhYdlqyGg0wjYj+7dj2ajQq/xl
Dmgc3SLxsrGYeFRpJoneEOhGlZHt/mRVF6wWa3vx7adpgwV8S3DW22PuWdbnqKtP
NAIQNEBCz4lLuvGQzSdf5lUPoR+5KQmh0huqRgerIaomKH+ILseYolRFQO+NHgXW
TC9sLFt4rp1Tq9ySJTOwoh+1U/MwtEjQPfyFPyK1r+wKu8cDyZmSRoMtt8m7Y8z7
t06/W0XYZkJISChcjANg55eGBRErs7pshxd31fUccgMaJhu18RCgnnoBLaZJjSdl
J4NmGc0O79WMVxOFRQ3i8G3JLxJKf2faKXJIL7jEZxWyeBXvkd1k3XVfxftdkM3c
uJ371G4Nxw6WN8CX8L4/6mDzCbTzQxi+HcLwU2ePNZZdbEW4OkYMT5U3eCuuTwJQ
uVSXAWscrS8Clf2F45qM9mbU7zQQ/oZWNC4t8rjxeIIkDh3ExVUKdRTcT+6Y37wU
LRwgEJdkzO7Dk2jU48+q2uBBRrdv2rqM0Q838julm52wBn039/f2DhLvaT6MfSVZ
8bO2gCQvA16pUaMbgs/6cyDh2fY4qLwVenSEFaeMHfRdRgLlcb/DLoT6RhMQ3Woi
+LxBuLQMuyN0ibyTPEQXq7Yp42NXjWKqkv20Qt4AcmptLDHkrFqSpxWGdmxAvbRc
seH96jSS0BAK8DpXY/Vq+U7zJxhRX/RL7J1Z8XuaePKjU5hYYi7ryWLiHGlICuQa
H1lqe9cQ3wJNbwovD4yZ3ojXSaFIHDdqLkmgz6LBqbIPTevc0PCl7iOO1qLkLGHy
6mBifywfeFgwOQ0Bg6bqAuHSTRUFP6dtiVpYq6j6Vqz8IHPu6XNu8L3C87/dWMPr
fjlgaIEs4C0nxvIXBACPNivNNoVZX536APrsRm7tx6RvpzUnTM2lAbLfAyHAGFoA
gDUC3DtkqINWMT7Lgg7dlJmMG7zNXn1UBezrn6OryfM6qEoFg90cqkr1JKXpfpLr
oz25g158vRg9hsL2Bq+j+fei+IUEgrEYa2QwIjvZ0Qhe+3ADU/NEHOYQdfZKoPIo
DAib1XOWr0g3kmcosKCyEOBmPynvCpBtfzP54ki8n0mnf7whtEumvKuwH+HTt/JV
4JphqMXLNjbeREbXXV5R3NgErVbHayPM7/bFQyjDv8mg89HkRirIB4BR6CfsHAME
fu7fJ65end5RfAuksDzE3HShqNrz07GXIyjf3YzjrO0GzYmYvJyDYvBlz/BKFYZ8
omAT5SBtBJ7KFUax6Qj/r9zVlnkSN/1rt3e30teJOHupkpZaFLZuSNkK4zbsAcqt
+FZjkUmzeYZZ6zZMQuXQ6YjFmJT5HGx9SUTCgjCSfAgHqRVZ8IJOiNh/TZzPHhvd
l3LUPKmY9BizbzUhcifOgACT1OUXhEyKs9K8bK2K2Gt+N7rq5aor+QKrdo+rHvCo
MD3Rnu7DbljMhukues33j57T8YMvYbyOM3oQG1shCpzkQm9bn3C7t15cEmUYmh3P
10zsjWVTKBFx5F9YM+T8kvqpgbw7iq7B4VD+ioPK+9X5yIAZt7uYVKctcXLqHQlF
hQNACc52VOEK2mD9pHr89UfScl90D3rastaVeN2tz52K0+N2kXTCrQJbQ7UqtCSB
/4OyWr6GNyRtD+casQbRtjL3X51qfRaM9tbkDQnRbdFNm1jarlIyC09hnZ0bF7jR
Qca8w8urMruJCZHulaGGccz63EpFT0r+btK8tFmaUA0mIvpPDa9hFRWSKt0WVWmf
R0VgwN/1+/Haz61xzbXwmGnNvn+wGeX4rxAw/TqEpWchwrkedVHr7/Ipuby21GxA
P66379a83buD069pFfKAemUtofC8A081/xcogTTCUhnQjoayzPNkeeiBGBlIAyUi
o2af2h4Z6kQDYYgf+hBZg1/HMYi6KoXQJjL0bXmDVvRfynOvBqsidwFw557sEwlD
weIZJZlpsLpVZR35ByLX9e93fXGTVWpX9Z8yykqZI6HQg9b1LdaVCbu3c8Qa8EPc
bMfYUUYwkwqtq+yvbeVMCBdZbsRcH71cjApDG26G5D1ceywH0nFbxB85A7zXL3Ro
M0NGuZTaMK7HarkZ4WPpefWpJCjpVKwdFbGzy1qeJkgYV33QW6PzfSgDKaU6Lq2v
2RaYpUw6sh1LmygNE7x4uOwfae3HfbzZ4nJ7QeWrL24TamIYieOb2l4qCY4zyTBh
6z2dcc1pgjqy6jj8jmlWYxSjUZVSDQd2oBLUzb2J73mNELgblr199zDDQLz2FZD5
lUfcrrw0lfGJtacPIUVPOBmonbWdDP3vbKogMI/c66qUfiAs5eEXzE7iKgpLQoCn
+RLqAfiCwpzN5lMwrj0Rvyre2buNw1mQLib6Nqg9VA3O1DRcem5CSwrIsraoTdli
ijujOFozt8wiVJ5ZZDMXhQxwHYk39uPGBv1GQSHuHEq8Ld35/GOLdUseZ5ImuZMc
AKM/vsr4WdXDtkz66RFYJyGEOEAa6iJD77jOw9x6vBuxpf84oqmrCvIYbxR7nO+Q
oHjynJU2zOgztohSaMErvYyPTRXyZeEB/AsV/IrDAH4Jojpr9YAeX1SMbJ3C0h9f
FHMf0MO8/EF3h1TySuK4hwq7mbAy4/TiDRm57Mung2C33zJp70HgBI35G7y+C4yw
+gH2gB6H6IFpu4ZP3+18JkCcG3Gb4LlmfjZiSFUYAGatp05K/6z4FAPI33C49MD4
5iQBGB64IGWF5h1itnAyhM8aAXWbzTgYMWb23sI2iYX0a1gt5J9s1feXWCle6Xd9
kngUwBxtgTmrHGw7SSginFQPt+esKkkxKInrapdEpYMD3v/XXCW0ieinRUQUPehX
9mYV6ZvHcqxsX065Iayza+g2k55INqvPfr1HY6LRKoJPyXltce0I9U+T8Ni8YK5U
BbUB84UjfYtYZc0E+Fc0YeUL6L44PvdYkSPEcgkcKZRZpyiw4lAi993sGwE3uLVB
yHFk6zLW/tCGXVehXh+6HhHXhNGbU924ik7wEMlQ3C0=
`protect END_PROTECTED
