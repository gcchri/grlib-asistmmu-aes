`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
blWHX37CE5DAKgc9ms3G+J4IlA9Eizr8TdBJhxSKi8hm24Lz4qDjZOKXdYF87XRI
gZ8I6Z+6YeE4+8RNrL71Pk/1CuFy4tLrCa2dMrmjZSahsYOJwoz4XgXcz8QC3T41
K444Frc74VG5JoH+30/43fElh1PeV2jZrTJgQBeAVOZFxCqBXRhlvCQdraL9I9kR
+bqddudGbSb0m8fM2GP+JL9Cl2NYN/KRDTlbYo2YMBtVZl+597cyZSPmujYHNHKV
GpMn5E2SgqPBYGaKWVk6q0zb/Y/2AIjna3Vwdjp3231+YWPwZPYGhQ6SdWj4C4+7
9jHVgtKs6f6JIFyDnnq2eYxz1aEkcDK+tAaBTXXGXuEn6MvQqZkGvS2Lfv/MVxVK
r7ZvDjta7CGkYCVBrQIozA==
`protect END_PROTECTED
