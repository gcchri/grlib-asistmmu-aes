`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
impQd4YIuXIydZ7+LKh7iCCIoiJuNNbRvOQ1joZeGlQJHugHx6eNeJHwHDWPVQcr
hLS62NXW4Vt/wNjRZayDqnD7bzvAF8oLiVbsoD1ZHf9I5lMg/5mvUaTvdWlj3XFt
EgbTgky7dCwnizdj9n9tn1pmp3pik65InoqCF4cK5FrZDw82n9rTo09FOBLdtPO0
DVQcIr80jwrXd7Gc+qU5deivDTV1A2zvRquzcSiFqugbCcCABr54y0yUEpzuwibY
ajYZCtYOif0IpSQrXbwpJun3DJdKCjTCQhFcat+OkGVhgcmm1eVl8g1YWza9pLg0
6krh/rbS69VIeNam4ZoxRXppk4ni4D1uRTZzAYn+EpJWmDl3sPEVbu5sVAORn2cG
gu4DeecOvlD95ZlIDSE9HUr8LaCwrLN5N+vO5OzIoUuREx4ZcwyBV+5bPTz8ZPgz
c0Eu2DwmfaqE4ZuRx5oYCnAdZLIKkCJKC4gq26iT6+nqAB83hhGtujE9LUI75Mdv
7rl28OIInWbClRVqmNyL7SgUjfLly6mqAibk0PP1jcUaHQ3HcwryA1kx/AYiMcaB
e2trFG7H7yKqQb1LjNssNMoJX6VgivTildEu0i4+TJkjT6KmN5ENzARL3sDAc20o
nDxUe54aTal5A2YRZSgZIBgfF+Jlr2Jsb9CMAMsKoWqG2SKkD69/RmcvxO+0JvQC
kC7SFLowvAi2ZiUEtilS2yR4mO+XxFA+SNRXCbbgslAcQ+qN9/51bU+mE5G97Y1l
uNUO0PhA25dtutJoDto0y/h7dn/ew0WOqbu72JBwEGA7P/31nlMzDrp01MUHmufA
GvtQgBNFKu9K2RG58XBxpvifUbVE3+KIOS2TRdqmfEO0/cwAOQZ6vmVtuD4i4rLZ
f1F/2C6oxJVf0nwzQmIUd/xNZExKZHJkr/mkhvpBq7p7N1+xakI73QHNZ4ELYju6
S0BRL/ZtkDlj7IUXKiZM74Qhx1twgYuz30+hSXJx7b+Ko9Sd7QYBNDDOqx9ZaEf+
dHdIi+9oGhQl+fyikCEuo9TFlWgb8tWLUjgtlFe/0e/iUgeoE2F31gwL9h7dbEWt
aQkgmzITIDUIxLqF6rJ55fbl7tKE2wUXR3GY9YrLOZ7JRw6JerOJWQJUrP+bpgBH
3y3CUVdUk+Ggm9LStaL1Aynr4/ewh9JLzDMxTb0P/wImHBMf1e8IodKLayY7oX1b
VTBctjdTXoxD0sxCLEfIWbctvWlpBeX2ePXvNb8+t5IfQ8F+VAXAFIquTnAn3Alj
x2QG6gEdS88D3mf3YL+0TmnPG8yX7SliUJGC5Uxc2c9bXbEU8qx8iu6VeyAljQVt
flG9DsNU6kXykz7ATY6ID5iK/JBALyUlg1t1qGPNdsdYnRLrrlL5/R1OURF9F2wC
E4TLFGRYaBLkqIOBZHjKfR3nAj5PYKXlfPFW6X2O4H3qM+VhwXcH0lqPWtzIUgbL
+SBXkXlvkix5/MTTYJrDzJY3yoN1S/Jg0u5ZewLvdMV8BxrvEHQoo+z7NsTE5TD2
eSNA6xTULzuigZRU+bVyDmsV6pJJQ7tnZD34U4S56SW3Ljr87queL3lOPq3MlTXm
ZECJlWBBOfvgJdtdQFeg4qYGfm0C3mW6TWcMZBhjoEzUgmQPSH75fzrZxSWeKydn
fQZFAcc7v0rnpQJXbcBEmRqRlr9SEuFy096uqZUbn0lJ/pwyoxy+c/4Y9POrliTS
jeT0voahmL7FVlpTGGOHxaj46E/lbKOmm9co/zIU1YOeYVH36PyQivX3pILGGlmT
YYI6NnBRkbww8boIA6q7aJy2yYS91z0JjWzjnK2WvATadDW1UHcSWvqg6tiqFQw6
S2VHonfyTo1QLiZEMmwQZXOMITK1t522FSJl3CM2j7jyx0p62q0L0VlyEMKr/TWE
BXVcUrx5V5EgByUP+vwsyV6HcVcNdvggEGebF/WyNdu400mpsW3H6x58aXmpTsVu
1tBOa6i3gBV3PvMwXKVUgew80FSLc9r0ZvNEK/BznN8=
`protect END_PROTECTED
