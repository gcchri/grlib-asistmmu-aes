`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KRI9rJH0JhgSRHBuodb8/Jbm3x3UwdhrZYOuj6tO1HALJwQzzBdeITNK3+6iP5xi
j1CTVGSjJ/fycqLjZS1JjlKVah6j5W+M8xCW5u324wUa7DsrYSVWzLqCa/5miRUa
Ci+QqBHSH8wn9oFrZ+KxVF4RWaPWMr3E5+obgG+tLdi9A7OSU/eAG5ZIwpes6R/c
L1yPemHif1MDhIQY4SIBxztqUONCc2JbAmIwBVLvfAhXY9Kg/0UoJ7bJhaekPKOC
ARa9x9HkE10k4f0VMrNmqYxIfRUW01t/Lkt6R6pFCbPQMpDTqZhf0Z9Rd0tgfxaD
ttMb9yIJUJBluyGjBFsW1gs+Hk0K5AlZORwE0KZh3VU=
`protect END_PROTECTED
