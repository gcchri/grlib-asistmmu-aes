`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jde4eK0FcNEee3z9ICbp2OVB0bBOXxrTGBUD4RllE4muH2pYEsevVO9jP4qcnwrY
wdV/5V9m8qbbg8/ld6eRYNiVvT+5sv7ceXvSECnA4Br9v+4od8gCRsY3X10+GSFo
GGN99uUxUVNviTEB1SPT4vW1olCVTmx+Gx+CjjZ+RmPx7E0hXV9k2dDIGGO43j+0
8xuac13Tql/bSSicyfEHgcO7gIfmxjIZ/VDFJKOY9aswbwRVdam0vua8BE1NnOcO
N7HmjliQfbhCp1nBXp+0NIt+zTVzoQEQpkB3qG9xcSY45RB2vulRLrKVrA4mL0Ue
xzxjNRuT5Kvs215zfRMCXLMmTJhX+aGM49lOc7LN9HqWY7N1YYTj4ztH1ReAlEPD
PlUDVozlix8Kk7DqBsY8PQ==
`protect END_PROTECTED
