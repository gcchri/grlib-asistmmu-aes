`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xnszVBlTlR7TyGVj824dfM+jDuDJZ1cvAWMzZIfE2dBCKs7zrYWGYJDk9B73g4GV
9wEL/0fDkC8cZIkRRQeL/1TIsd13B0lgl2gQUMTNDNZAGgKQr4qlQSMu1QeevMcx
djEYTi948RDU70lilt8RwlAdOasWFQorIpQ5HHBUqJ5xyOf9UnhdnAwOPp41oSeD
TQ0tVtaLbA+3h2chOyKx/G8LXa9BJXFypQjfLXPpbA0AI1zcwboMwQYikYU5sMkc
ff66K5r4l0+AK0aDjIXOiSpuL+CossZmEyKVeK6E6JA=
`protect END_PROTECTED
