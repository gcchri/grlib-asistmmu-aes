`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qn4XQWnJ5gahl5ujLVyxi+uZyXKaXzhNgYd2v1EvYnoOQ9bK7h58BUUIEzY1NIUx
46K54OYfMqFbWpVKW3Ak922KCy1Lh2MazhOWT7g3PvReFTxUO6HeXqMvPpYHeT9L
Zdg1oj+iKbsDlZRf31y5bLlZOU8s1RJASuLrYEp9PXnpVyma2Jt3Q2cjcW32Dp4b
hFGC6yOyiMNQRVxSg6D/fsowgEFfqy2cljtKOnKYcreN9RWkTnSAySShIAxOp2qT
CQ5ZdCAQ6Cu5n6957e5/innsCnA5Db8J9R0CINfp4IaCfBFolhDkWibBXJrjEg1G
Aoqd2ravjN4pT8thTFw7WXVjf0Ij01t9MwvcihY9EFBhLP+dCA5KsQQZHn5jUMpK
wZApueeSsXzox6S7JN8ZG7a5tYhGBHQGDw4g2k+VY6fCfX/mmw1gGe3N2i0HyYsH
esP6aQ8tZPaHdBjQw55yjSoSw8OpzmiBx04FxdpLcRuKj6iUpIhZoEEWCuhk92Fw
GOwwt9KPOgXjXNDdhh4SbdHnta0dD5Y0+6T1iNt9pa8o/lyPK59XtO2sg/rQGpzn
8atmUbEcylxYRVvT+xtaUQUgTjOi6Y6zsWlnKWWfFSSKemJYDXogUXBG8qdKKJBH
hOMg5LQKfIu0268bYngTNJlcSt+ppZGBxVTf7tRPkB0ZUPGeD6Rac63EWc1M5LeZ
oNcTXvrRI8nZh7VGui+1iyHM25WgkXPZIYGT4Eqp06Bx1ZpHxZ3penxuNfLDB+5i
icF6rWzYgbsiQbnIAEh5Ynxx59rhidDuKdowQsIzg0E=
`protect END_PROTECTED
