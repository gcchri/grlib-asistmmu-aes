`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K6vymxlxJo0sHyj4+XTHsTh+a7yy/65YkyuTac98WdHdAkSYIbKaoDMdX0+cxgQF
8AlAAazci+z2ZCw95xwbeRamf+P+yXwt+RSwYDU6JaEf7TUo79bXxFYlqudICXVv
VBAbzR3qdPLYnId7vrKKtXSUv6QMz4QYKTxWLEBLdAeOGYP9cm29GaYbhcSPo/c4
itzIvllRTBkzXK27QxENcv/mj3ommxv3Vv+BxBxKqW1h5DIrX0HmbAMGI3+P5iSy
tTvOEX9qbLCUGQhjAYMrHkN8l9eGeyl/cWwZgaPJzwW37nHlmlHVek2MtNbxAzRE
ib8jvBsfClHuXSOBBONKhqqk8nD22mlRrxnAtxoBitLTsmcVmQkbtKtY8ja0xQuj
YhI0pCD7o2MQEShOfYF6RQ==
`protect END_PROTECTED
