`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
juOO9V38/AUePsbt2BmJAfQKRRu9c7XgCih0R9OYnvXYNUguTuxM6uuaya9KAv00
NFnot7DoyXbe1ri5lgjkSOGeEXGB4fQFhTlryxWS41m4hf8DEWzgN76rEPP4ZWrH
AwpAyoehiMtY6XPnLYp6P9VL1go9lPuy9hPkqHu088aooEt9NIWe7+iWa53UovOh
ewey1Nni74J/pKVb2ttOVaXPXV1Y3+o0gPIAUBLcnJY68V/3rXigDjHJLKCTr3OL
VGyQbKd82uK/rUciaV2I/frQrQYpLwm9aDFUYbhJFy1ryHCha1iZx+olr3QkT3yd
X2LPb9rO3N5XZY4879DQMHd1Giv0stUME32IL64+lGH4v5NhUw1wade74cWX4v/E
jEYEDLyKOlsXb6b3M/mW5n8833LyhX1GoihbbyRJ1ndYMXLG2mjIPZYSbWJKtR9B
QF48xQ8tmcfl6btwhH9ESxBFM8j/jsssqE41N23SL0ZFu6xfcNHNYBsusKOZXBHa
o3CA8Oi0+kCf3Jmw8PkYQ8tlmCQ+C3S5bDi8pfJW8KkSgRNPtJr0Zz85upIpq6Nb
0d2EaPfkNvrYcLr43VCXJQOFkWZsMCerZrGdMZzpbS6auhivGdzhYDOH+DOdcjR2
6DwiFakyCqOLyMr26hVtp5rPHI52pyVpCN2PP/BgxkREDZtmZEo/fcNRhv3iSWev
ff30S9JV+Bi0R6x1gfaBebmUaBgsS2e2KuxmwkOIlUZSTRy1zAzLD9j/NMWWoTjq
LLMmvD8sIdOnKDYJI4HagQ==
`protect END_PROTECTED
