`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oBXnes/zDidzk9GmBpA3O55LQ08jDxXzMwgNdk3xvObWoj1e0vz9X/1QLBvPdPKn
BidcxHPTGsaNXx6pWjGJZlGEnH5F9EDFJAzowUGeLPkq3D/pWhB/wVR7rX7RE9Qg
SteZO/iH4XelXbaX2Mkrsu4CiN5YEX9KPpqHLHlcvMnjKEV9HWsmHUB4ENKn5461
3IhkbMOXs4HFv9bfbJowYLiVl4XL/tagTDsg81lVmHfQg69U81ymvkA7rLmnIk51
3CBYMco2EQVFx4oVk8wv6QWB2kuEVkOuJqXISTiIjXV1ytBWTmL1kNb1pzO3AQgC
UA9PgSIj9LgHxM3X3NEVFrcMO2T7PE5e4KzuFNWehQDWOnl8Xz+4zn3ZaqHRYPxJ
MckY8n8VdrAewk98vSmE0CFyy1L2U4ytbmZPOPniYspmSyK6ESAdV69WvbZGocIa
crfJRJGzG0ZMwE5tTinnnXOVxFVpqivtCyajd4h3BRWWpo+ACsWuRiDOSBraIZif
+yZhAqh8DtnSsGDKUYCseiTQv5BmA8v1ur6HAXkGdhTgfydbDotpMpX+82G7fpKI
fItcy+HS50C+RVuJZLl3laWGgSB9qkAcxXSF1UiQvVWO8b+dtAW2ih0DPwOgG1iB
4YIrTb8QPzvzW/PvQouDMOd/PRjLWnb5aN11h1WIzZlYgk3PAI9nJ/dxkZm804kH
lZLMz4bjiCU0VMIi8IRq4fC5GF16ClvO7LYvLEIALl7u9JF/bScNCnlq5c1VmOEL
lKoP5dcGV4od08wgAxVEvg==
`protect END_PROTECTED
