`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rugqKkDToGyk2BKfmxwFC4l83LtCXFdvOJ8TRHAevs+nLhbnffBiEmOqzuC1//Cr
vzgyWl7rpPuoUsjZ60kZNyiojPWcMIhLhwm+Ypuh5lhe/hA5tD3tTUZ1T0uo6I0J
e339aFvz7A7tdZ+4QMBk/IrEzu9n2ylqdg14ILbycBMfRD36ijuDzoitaQ6izVkI
8k6+dKaFbts/tnjyRe4s0xVYeq3CTxnz/UvKp1ThH9ooDKg+W64ndQKKe0uCx8ZP
+LVIlz8VN/+EQsF3WB6uOAyL2j8a0F01Qlw80Y0bMVdl8asJXJQScTkp3FKesw5f
EJkRDsWJH3VhYsXvZCEEcTilfnQZmVFo1MxIpJab0KHn+pClrDOH6584eWoCMeiM
OnhwP1pYJbP0IPqrW8c1CA==
`protect END_PROTECTED
