`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EHo08CNQEOrp8BMZ1wn08zyCMIyF4XVcOatriEm8sraTHh45IM7tH4pNov0vzYf/
yv0LFkIhpgZ4QwN+bg88zAtmQgNWRskH6KcTzz2tzuT8/r8bg7i1UdQmw7FWBloK
CU1Nf0B1Sk6tDLoxS6bqlelIUY99oCVsnyrhiAmNdGmYQnSKp90COS08NCqzcMui
OjcXxEsmzVjkoZjh1Kosd51sju4hIo5MeqDMY7Wny7ZFd603JWR7t/DFcuLCPC7k
0X7WJM9yf2fCXz1CVE/kqifZavdLjNCOI20xmFCgxcbAUWVHqQ7dUldiUwXbm53K
`protect END_PROTECTED
