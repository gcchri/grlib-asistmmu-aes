`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
60U1XCjoAvq0skpXWeU8vo50riHes1+yyo2HENZir0gRsD+0RScBrlhd8yQyVkPK
DjUrwgQnmMSpjtfco+uXDtyrSlZnrCzj9biyHAMwjOznZI1VWoxgT/+15jChLXgD
MEmmSBwbOTVC4WNFQiShoJNAHQDJ5kdd4FHTbGs2GthAPeMYjZZfx/lJyWy4e105
FaZEW73hi0yNCW4aICjnP0gW+YZ1wZeSrwgmg5tfitizCVnnT5krXNV8TFW1Dlr5
9tP+YKCKNp7guYDUtdzfIr2wRINlca9Ao6/6SvDnrB70lbZ253V7MyQVxyoe1PLN
WZ47458DVyVG+7KjX8jIsQQFxSqHpkLCVAEeTWO2eFr2oN4xvUWdwwJPFQ0oXX76
JYA7Ze2xEpf/6jxFq3xbkwoyZQFPXz2P+48MQAcO/FU53UkPjZe3kQcS2Q0216QJ
PZU8jd9aSKjC1eQN6a2lqs913vyjLSUjTN0ADD9lL/Eknpz9ovOgSYGz2zrMqbpb
AcT//PWjL+TtPrxF+LimveC/uHgcdEwbkdRD65VWRuYos3Bs7oibAO6fF7TlPdmS
p8uDqsW2ruE7k8oUMkdGx3VQkJGm1/L9hkLLpI5M+tX3snabH+EXjla3MDTUroJ9
k/XVCNpM4Zqg05AFim4MheySgE4xPUjKlEXC1ostX0JagY8EvEKjmGfuINrjaFyw
FtY4vNDuLyA1+XgDn1+VuoQmXi1mQbjxH54sKV3s4alcONESc43ip3arOav3gxhU
nFiFdjchGNm1vWE9/xeU2OEs+LgsbQgQ8eXKuzO+VopQVWB78K+4Qs2sT7Wu4gta
4hM51G74H48SQwClM1O1xt5ZHDC5W7l0b7AXkWmNSd3HTDnIvb8iWIYqTgEP5GvP
HYZZxnQgoHnwiH7ahzdc3qXhbvP8eiNlLj40xenI9HlLPRlPAkrDAm3cEGc9Wuop
STIf8IQ9aI5PdWw/WCmCQdZQ9YrNsk/Fr5axaU6ape++F7RcLdMwxRSVWU13DxU+
7AcKVEIynct+e3aQW5kjWKKRpb2JAkgotk7wnsalKOqiMJ/q7hc8mRJQ4Rb6qncc
b1avlSycQ5uYJv1pAcbgPa6cWKddhKedF9ekzoW7fCcouuMro2R4T9XPzthkF1iF
UtTDbCKa4noEMhpBYExogfaOpY6Qje6JblhmjBYiguXjU6uoSOudrUvaWV0N+gkZ
tM0cR+OykDOVjqyp+oIIKP5eOMdIc1syZyFIHOd1DkebD0pwV61vwDg1JVqBwupc
kfLUizfgjcWYQoeUZYQzjPFBTZ1Crds+5OJwzY7E21Phcf6le5Fd4IjJj5IbzK4a
5ENsLRxvbCyGiUEU+3acemWJXeD52w6wkoFePKPIcIrpSIXW+ZCf3eWQz7B7ap22
RiS93DfU/5tGoBM6n2QLW9LH417FFk8mkKhs7GFrGYxpDGslqbF884aXcgiRP78u
AX73q/NERxA+uwhKqYUzU0847nXQrAraeHNg+B2AAsHOiLEioi8lMMrah/tpYrf5
CvbGTBM8CPte11wMwvNCrRYr1/F0ZLseqBbFhGZ9NKbI4PB+GMQ6/wYPLyVN7O0o
gKuUUE3RDInH7hb/5vI+9RgEm+8VtRp6g61Rd95w4J2Bsh6vwjT6fsPP8Mqbk4t6
Ck0GbdeK9ZZYH9Z+ciGkPt6iIlkTW7GYLAjzV64IRV/XGAQ9ShYVopdcgUBQ/E8e
T8M/Fajh0uqdo+QLjegnTCXEMY3D1iXMUqEnN80ZQ4j+oUS5Db7N3BbYV1L3rHUR
kanUqzOUTGU5cllYFUUhiOpsMpA7GwulQtP5EKvgLQiOBZppmNTS89Q46srdcU8n
7mIKSBj2DmAT8Kj3UR6C1BFFA4XiYfcbxIH9m986yUuUW28I1lk4XdPrqzuc7hKd
+uRv6MjxnWsqT3CJMExaOYUuaoDAbyOBZoNI+S05czbLlelcIrZQhD08wb2MR5Mx
2iQ9vhn7rsypOLpYK8r21g==
`protect END_PROTECTED
