`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
08t/c1Kpa1fTz6gDrMCp9YNf59I815bQ7TfWqhixgz05kWAqTgriD8Zg7L9/As0V
2WIo/T7+wAQw4MPybCGWQdhCry5D/Y/iHCk8dx8CgmUyqqYzsOtuN27RKE5VH71h
qBrvofGk8Ui3PdSRWECZ/pSYKsp0hIiz/bduWk9OxTIfroGMnpLzE/UnFCLQvBBf
ZdPgI3FK4VMOY50q3mnWQxRvTr15Ua9agUKwbV3mSyu+SzfqvVXjHj6+H97GgjdM
d8tikNXYAvNldpEoZdlCEyS/e+kCsjmucfhAugd8r3Q1FD7Aj9HYOnH5oUbJP8et
Spn13dEa5HlzW0Yil2q09DsAkintUvLziMbN3GiBGxiBpuoGhzNDJwqr09WWtunl
EcC7LC9+Oq6dVduGTcKH4CyryC9gw+KLQH9iPw2zQHylOMOUkcvgAaF6SLxKVZd3
5igkw+TDucQYeIjHZTU46b9rKDpKeWxEq9zhbBRqtN3/jMxR/XBtIhPGjV3fXG7g
iv/V719K7Hk2qzEHh+qr7u14j9Dhu2Q8hhD9XVBpTvhUUERvl7a4MeaZbP8QbDiy
L/XvmrKvQrqeYVn4IFg/KrpNboomgWErroqkuml37G3j/M2lbOTMFo8dHFFLEXq5
jDnxbpts3coClwQk82LUJcchprfedNjB1tr5SQgivbOAe9xLo6YzG3bBJBHzgtmY
OD/8OVbvYc4bsHuwMkuIwpowPBzEbWvr7DhW9MH4NSwJOXkDMk7U+rE2nZoiFL/+
w3MWCNh3jHFpCHeThjVbu1u3dFDkQI5InMkEOcMATg9CcZGXg7v/GP1jfDWfhmUU
m5mjpZmIXlHVnz54TqwvD5KMaUmqb3RUdOnpvz4DC3o=
`protect END_PROTECTED
