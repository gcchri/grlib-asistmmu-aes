`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gtxTrqwfbNXC5snVN8tL2O5XZvvALnY1zVvQUa8HBOEVALohlNZ6lcuxwUNW50sn
PO1t6SpDLME/vl7H33Fgu+bpMR7wSkAHxg1zQVVEM2Kzdbpt7IKFAAnXD8voBH8P
hUt8q2Pg2JSEoKMU6mYVq2rhBX3nJ7ssVyQb6y7KxVlUTukrWKgnSTfpPCxtxykx
rVTdTKaSIvO1l7ROMLISyKwQkcNXV4HjxiMr4fPoCxbM1gnNITeLHw4v/ZwCcuXt
XLPQyXZVP49/iMlJH0KwZzomNDeWtKwDB3+GcTxY0ZpuaL6WM0+Kyzrd2kGXqlnB
`protect END_PROTECTED
