`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MjF8uxWSOIu0McdgsoZnoxzQb2OqYNJdYWQBnC5d/AJKw1UzZzjPJv3lYur7tMp2
3oqFcqeqPIR3R0V6JqX0lltf2eLJCeR/zBFg4jy2I+4lNKCqpwt4GU86pJ7t0wYp
JFkVp5k9OT40IHOs1gpQ1c8tHphEgseqNhYXmziqdKKmDgUFA6wTtxS+OC9NlADb
DEO55iw3cBRWLIiuAcyT6Cxl9qO/LvmPSWQVdrYScIOW5kRfH65CdeRnRTD9bWFe
HG99fCIBoezH3LX1z0gb/CP1TTppJ6xnUmexxqdZdvaCqmyVFBOVGJGzm89wnkA7
FhESd5IAEw6QNmh1LhZ6zpXBbf6gWX6LHJO++gZCOhRw+HH369cHLV7etqjhxkkb
st0PBXqwcULTWnSJRNpgEw==
`protect END_PROTECTED
