`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SI8Pxsommmb0tJk7t7LAWHenwYQUJjLqySEx6KQbyTC/JfpkRbPCP1Tau5+rLDF+
e8vNF2M6Szshk7p/OqGS9YkbTalHR0/ryjVkYHbphr1OodO4vj8edbtdSe5HZNCq
LGE3i1s9IqzQza3b5eJThcl6n3ZAb+cYCwuxfwfmnbTBqstOiheK2Cgrw0MMcbNa
yOlFbeo99DNjQljNhquTLpEOkmZ+fBDZM/AYsC5LSfk7RnAMo10iM1cQqhzIddjD
5plvr6wqupzKFohYPm6Ezp4PqOXMSE1Jduujkxow0dvq93iDEGtKfqJG6/kVg5Ub
pXuMxFaVj+dqZEAhQom3kvxB+kpJEWnmrLiIMbgNbxr5zh4d/mk3GvZnTHSYNBAH
E0EU0Q+eeyWOcbn+gHTQS26Ji0BcfYrjeAbtIrMmDxYbJdLop/4ALS0OFlwpcaIm
xu6SOpE/7aciQ0hG5Oqp/yQN2ID+DwkiCB/Eem+IQ43jxMcRLHYgQvzgwkgVWLif
ngoLaEYK9P0ByA8gGeqJ8sqPK3vye9eKhSmJz1gqCWdwTioX0I3rJ33laoOoivGO
xdCtAt2x3ZBan91hKW8aeQ==
`protect END_PROTECTED
