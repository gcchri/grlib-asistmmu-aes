`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YTyGqv7kaBKhKH2G1FSs4vBoROd4SL1iuPkkXAtRKXwItFeoVUI2BjcSw0a64aYV
ISK6HRtHB7GEHHsU3vC7QPhWjZLqZ4IG62BtKz04SEwEjLs/SxgacY4upO/csAFu
Hp+tAv2TO6tHpYd/Npp2vZ1I7Wpt2hlr0RD/Rq0yUxC1jsKQUEGDFSt4a3OuDIaR
7movOVzZPt69Zhg/3xC0giOMyx5PwUWtXSKUa6K8lA0G3JP8KFaixslDCVNVbW1C
QjNjMJc7n5iv7hvzzLJzMXoXYc3vOB4ZDNCXOazZx/JtzJLtmtKU6k+jnrvRHLN+
2g0Ij9AfSCPWvXvZDSOtJGf/pz7wvi0xX+ccHvz1f0ozXMEk2AR6XaBLipQjfYW6
nuGaEmu+sM6np3yR8oWbhp/pd8Rw3tsQAdsum4+ShL042rDstff5GQyTmVa54sbe
CR1uX3BqPIdvO6Xr0Sx4JQJrZ88dC728D+b0CZ93UDDPc2hayh33ymxzDvvpV0Fc
exYDylTgijqDiz+rozo1HXrRuC8O1LVZ86gqY+jj7Q30WE2JnSRUh+vQFNsPiFFf
`protect END_PROTECTED
