`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
niMRBwfZG7wkzKSp+DdCB5aUL7WzSOohJEGCGJeInw9exJvpyVCAkp9U8Yd7QSbq
JZ0CeZ3c9Ol26b5CzuoXAFhAOTy0rsraVE28WOxBBo02XJoS0v/4JyEsEr9TFHe0
RP0zU9vtmIZL/IpK/76M+7/3avZqnXeqLmO07escbxjhukPPNXH1rb9fMYm66w5d
XX9aaxdEN1kPP6bp0VC2KLI0x+Ra6w0pcKBkP0MjMwAXRMmusfu9IHUKeSB/oUsY
GMsiaK+bRsursxTEz7NrsZ/VXEvO/aAyhMODn8FLj/XY0RoBvl8psh/cm8Ux9i6K
mQL06j4NK1Pgl6In3398Vt1h4XTswL+C/PY/RBiFdMAMbSpZ0glmOz6DwJs+wIE9
lqVYEAMmyFpGNyR30jbF+2yf/I0aZ25hdck8460RkKQ+dHoMnahjRwzBtvIqrGtN
/mvXeZbHfI/t88eIzef7Fi3onjFmV7stz2n5pjovH7QpLF9SDe+IERuDHD6tRfxj
j8tkZVQ029tTxi6UZrIjNJCpcd2kYopJVjV6G4O0JPDeKZBe7VgPhGOmzODe8Ev9
1kHrjsLnrvd11fUQvZEabQ==
`protect END_PROTECTED
