`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/8kH2wm0oHvGldmQXpLaFmv/4vhXtgbn8rIRs9Ns+fZN9hLYh+L9CXSPFCa2ZG86
xWgfXRvxDTfP74XYzR2EoWl3oAp0giEXrH/OlWRymdchZYsKfyYiLZ5rL2MWVKIG
KcIu9xzYV1kYNy6wywSsLBTFNv9E+6xP1sPFpcMTiE28KcdjzXCJbggtxM6/SMxp
Znw9sFtgffHZuBu15gYtmxmJDEbSxjyb42mPLF8gE/j+SpU90Rq8d2IM4S85Uaby
`protect END_PROTECTED
