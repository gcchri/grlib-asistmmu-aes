`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fvPNd6shJDAGnfqUcajBeQgLYZoIUnWkSTI7KR12bFlhxsM3kAbn6jfrqCHcHOYY
JW+J4Zcd/bqKhpqeKvKzgaPXfp1y7JTg+QWRSVTtr7z1v8hL6ikyE3QtPBscXvdz
eZp8VLUtC+eAh+pxPf45Fu7o1fBBMRfQ7+dLzC/lBpEY1CnaPAmrLeB18sOdCBiQ
tMnfh8urLBGQWxHRF9Z3D2qh0DMK2Mlvr6L0qGH51ZOMSUpESFMfAQyqVWp5CV3L
Rbs1njvvhmwqpQ1W904GobKvHEbqS7+/z6cvMhdMjjt1s8IlrG5sW8TcQLyZlTkd
vI8ux5VwDz3l8turI0tVsXBrqeoFdC+poHOi2UmX5RNs3JdrU7HF90LqOqwsiEN9
1H7Weoal+g8WA2Xwjz7RLtmRRc3oCk6QaVcqzb5TsOrsYNUM89lC59L6vwArZlIm
YDeXJMGGdUM41BdyISTZP/WGG1I6N2XJNt4iGwYkNnmuAG8LcbpXlNVtObiz0g74
nAIpGb1IRGWDzbbdTpMJZLyY6aFNNKjleTcVruRAbprXwdsLjr/N6mjOnhPIQyy8
ixDGNihX3n/FlN9UyweNiA==
`protect END_PROTECTED
