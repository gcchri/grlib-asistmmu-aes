`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KqfyG0GQ7ahWPzhupgAkpCtd5O9wsIeavjRQVQVeoVsbEI2MgppkHDMAKDPH58o9
Tg6Y2iA6Cd3cCHhGqwYY35wMGcOASKejrU2TU+oor1PU0+VadYoX8Dqcu5anzrMD
8p+tca7AeVE9NHEKXo2g+EysHzb0i11CA4YenpFtGmSkj0A3NZvi5cWHJhkHrO1j
ExbXd/YtfQuVsQ/Jlrlv4eGr0I7Q276mi1vkc51W2xgot94Nzv1hr5isbiex5DJz
scsmZYTNfR1hFPgF5l9XX7Gf5yNKgTFaRDnf8mcx4S+Gn+HMYMAQ+EoUH1/++c2M
Y+U3e9+oLBvZm21Cp92pp5oxXiYxa6u/muAA19aNaUcEbTjEoKuF14Dow4aEE7mp
OmC/+8e+M5hpAd+ujclSL4jfkiPux9O/eT47RpHPrHvgvaL/QiSz2TY/z29dVBWh
4BlOtbQ2dbyDN1E6nS3sxNtCnbg1mu3XQH5LmxuhjfI=
`protect END_PROTECTED
