`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TkKL10CDZS7WTzM/zD79qvgSP9qNjAfMzptUn2MByYoJm2CRScdz8z7Kp1tCLi4J
xZZuGPpO7rNRiHgPrmoyl50nMcf51AksHR86CHFANxu8D+FyZQMfuNtDozb6oyz1
hfRGbgkD/ZQQn6cuJ9jkqBADAjUk4qHnEm24PaBk3r0stMZyD7ToWPDQ0eWXJD34
NCxRz8zjl5FieckvnMt/AsfkDAH4pKoF0sBLhuCB+LLvnWlROVbsuHJ+LIX9qBET
eHi9v3dN+N/L8xPIrDORaj5SjgObwrq/9d4K0LqURhrC8cgJL/q7EfidU578V7x2
D2R9cw9f5GYBCJYzWiIldNhCbtfSvJyBqMOLnrkz0u5KqU8c2DoeM0DekDVybhEf
x/b1hebUia+mxlWV5YMZzgwWmbpHa8C+xNPJGlm3GktlKqBrveBV7N8/6dt5AyLy
qG623Zn7dns6kfdwQCXYbVcfr4XF4HmfPYfONDOMppmmAR3XVu/TMRH9T9Fym4Mc
BhfWmGcNkzN8gUEZ3Yvacw2Mc6omALeoa+jViP1FsDXyXMk8nIGaa7cpCRlONuIA
eWCjmBFjpXJYLLKFiTwLD640uKozu598hQ5my163DE/t5ojqdRCCcVdKKcg8k0OI
l5wLaJ9DN4k3z0e52m6llSzkn6mbGDy5Tmzor+8KE7onFyUqM8aSTLiX5XUzf+5u
MXfLrne6uh/aDbsgX2Ic/6iEgZ+mis4YgveiZ53Sbsxh/Bw0XcZbzZgnUvtF2sSk
0cb7V8Rl4fsN7KDQzDXp5Jo8tUydfluqtzuOuJ06SYRxASHkhXg+pLAJXsaKHtFp
35Kgl2msVkWclDrkfBt4mP6jDYl8spt5YBimkVB8qTFt1DfJBoBXtpIvDgKUgcMJ
wD3gR+0D+C9epSsIYZ2r+4kWRM3a7wd5a8gL8GNflNnO1IscIBxw94vmLxp9VHiz
BMoWwRsKczJ3WjrqkzHS5a40mejc7/Q4hwtPCMcj9Zs=
`protect END_PROTECTED
