`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S5CfgdUpEDhfKodntSh9fgTM8ZzzN6KtZmew0dnILNjNwTlWalgK4lPqA1hpXNQY
pU5x8R34oxTQovpq3/yySmCx9v3dubm/kLoeKGKRh+2CoTyu91AELSkmZpcztEX/
7iWX/rohzWUorM0jXoauG4uYoDCLGWfq9FMBiSBh5gqAHSPlPOwQMl2Bt6qz6VjS
NRPg968QkQ8UXVX+8uGMTq5t6To7iCO/FratXiwKHzpuqgSIu5+vchelQ9BgA3BU
Q0hPwNAI5ujrvs0YzXYcZg==
`protect END_PROTECTED
