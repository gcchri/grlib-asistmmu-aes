`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P+nCIZPybzGnCOw7gaNEAgDcxZKbg6GGBRMTy1o7sOxYTVcFEN5r6UwS3DZzfCKv
3VE0T34+fVWgTTfx6dQHeLySZkkiHqbwMcm2E9YvgxYvj3OBjZZvHyYOA3SMIDNO
cS3OUUMA3uzs4CHRBmPobGo/DXUd6WJKSSTJjR0+XK6vEvU+v+3YQ2HyFLbslO3o
Nn0AshwURkl8FFhTToiHwOYKyZaP9C7QwVFhPC1Mb0tXoDafRQtbyy3jLrqJ3VEp
8J8dxehc+IbYy0r3p2WqtFiPZ6Pl2AwrxBjcqGsiU6DbpNY/JrwhWRQOVoUj4oOV
1CMRh7SOiEz+bt0j7H8ZfGCqC33O1QWy+5i7afVCzTVPY3N9gHtOSAKek0Fz/Bbv
ebfRUS8JEEsuQsmL7VfZWzilzoEJ77jNcyKA7ExCm4ToPQzBqiXtFVxIjhl/0YTc
LcU/oRFX6sHsQHzPC/RMfB2SW2Fmnv6PHQlDG9+91b5VcKAlNqG6+CxgybUODxLx
nvFJGwTvXN8+Y0DK6ba+1njBK1iEO5VQu36ecN+pS+Uhn0SlZ7zfxAJ8eN2MxQ4m
9a3xFLaE/Ck1A1j8GHSC9wbXqvgnotWOh5UPaXzAnEOY+hz52Wc8kDx6Z06GfxJs
ToDe84tth4aAl+xOLg3Nh2t4t48OFMumxBPbDE/J9ViqZgTGF3+gfdXEWTckSs3p
UBF5jNir5J/HiGwfbVeESV3zc07Vm7ygOqsTAEzaY7+6GcV2gZDT8PfTjRM8q/NI
mQmRRtKT1kmxspMGq53gUOB7lBQO278s5v8TV+c+ws4vawn3m3QfoTTP2qdfi8hS
F/eh4eBiji6DaIYfFUpFGJMn6YnTkTCrCpQFgu18KnDxxPMRaqKzNCNLKksNK79y
VBeowGcpBVgEqPl+yIr/KTXLbbzabi2kL/GH66+/4v+3VdR/L6/69KOAYFSk6xoe
3+u1X8H4o3D+sAeNSc+oEg+HSdtodXJECWBFBqDF3fmHSj4LDBZpYk1ZNVD2Xl98
e3yKAO5vtwTrLd4Wb/CG7ID4Olsik08z6Xb0Y3riN8P3lOkwmxwkmnNKGGU8ehvo
bYe29jIY2+beR0PGXDBjfQtWl8gUOvlhZm+SOyZHyZq8OgIlqvP0Ap8Rtp8KzSW/
qyfIVJjrmBh8gQPB9ZRE8dKeI/LxaWKMK+vfSpOWfwCyRKo+Hwj2kJYGoyvv7yms
nc+oNkthhQ3l7rtyNuTehvrg5YZEEFesE0UNh9clhWOfGcSli7irfGr60vd48Iy1
HaQo+itP1wmlBBwVZDbHv9tqYm9hvyCeFV/2tN1BS1DllbtZxGNHb35SYB1/3m61
E5wHq8/AN96kQpmaUaljDkB4bNaZJCra05r9X8ZBtZREvXa2i5vgFJjd9xrvyo89
Kt8vKTwDvDm+/SYhi/5lYy6NIDqvIZxSsimyo9Z3keNMnAX1NyOBxniSCUoJWzts
3Jg2IXVAmDi5qFIR/Wc+6MHFdGT1jrmXdbd72/jKgqc/J2w9++1u0nhIagJaoq24
Bn2ZH7b0TXGAe95tCI/HnDsmSdf7fLyUa1NNmdYJ3t6pPoykUoRxUWJmGHN4/Fmm
IFMMxz48ahFV9cTSV1yxZZyXquLW5Xw9DQL0NYf7r/mE3kXFZkWgtVrTGwxuyIT0
B2x3fNEa3WwCSoYW30vqfMxOjGu0PY4xxjQUynWdetXM7Xutg27a+d7ioUEfmQ5I
DK9cFaopAw/JKXw+TWvgbkO3A0EThL6Eut99XAXXOijiS6kTG0T5heWXkNdu1VCx
bCSoRO/WtIlNx25+Ks4Cl6PP6oeLnsA+boW9+0Zs+f5ctXEP3pA3G95RW5MwLgoH
lJBNnzhFFoh+1KJES1NQNxiJQRIW5YmTSHWVvZyFkFS0SM+oKFsRYjl0lVHBjlte
gy4Wawg8r4n0pIaU6h1/ILebu038FBDDIDwq1CKRqrNecwK3+n1vVIRwRRoUnAle
xgtcAnKwx0xxNo4M1xoKmyFI7z7VEI2ROs7dwlc58zZ79tx4BULVzWTteTN6R9PI
DcawfL3410v+XmwBlnrEkM0R+ku5VYwwI7Rfu8oXYYC1OPAX601QRs1dQynlkvCn
C16q7ssuFTxbJ0PKGleHA6T0zfEskmQO4xzl4jmteSmIsHxbSOAy4Wp562lr9GS+
8pGT1Qz5GecxIm9NmGXj5ONLHDPPGSSrhoS3L+8wmwXtM259IGCwddqNAS357jNy
pucn27wY+nYE1b0xUGwUNNJBpW6BxMuvyDIydwLm8A5HrwlP7I3UUu9jvZ9TL1qJ
aO2jIBEyGUSE3ShxVUHhoCZ1/bcQf/LdwjwPqdzpeXhvUQBoWbkRZnN+CCph8fJd
YjfXYJZP3W1MHtdA8il8N30tyzG4tg3rfNNBibuslKCHkfaBAZv6PL+FFzb5QRp9
hIcIJn5gSiR7UXTcNT6ivNYvGP/l5ezhvHysnUjcw5lBMoSrJ8rzgfZEXHuxu2z+
b2HJ14+dlWZEc4CdDXhBsuWodrmeUlOypPvgqQ1etSfiDXZFOyhfV3FeE32fgFsM
Fj5MJZetTzlTSLOKLRZNzCmmvGxUPPIZkTQseSJMVS0SmldxCuHJ7/5jUaLit/A7
8tg6jH77IwqTOyEBugoNR4Opj15+tuA+4DCZvbb6Ni7QQeFDleunhzQ5J0IbVHvV
gkFOKx7nY9HgKWuOYSOEaIP6GbEI/YeNFr0FimS77RjzXnk1t4lSmVgNzqlNtZMC
JABi0063KxW2ZpjmtICiSls4eYvhBbN0EKM7h9LB8GspbPWJV1Huv6cX9nXjQpGw
39ZXmTO9gO5EtXOxP86X0b8ONGvEkR2b4C5F7FpZ7qKvsunb/GFNPzyQXeBemIeY
OFwjJfeTVyPNctijieg9qcehSSt7VRU9UkmEXkr4ATs4Z6wBLmNXtORCpZh966hj
FjTiuXJNcTwP7eI/7jIJdWrqDs0CQazj9dHt7sGNXnq1y+GV7RBOGS1jMH6+ECcx
pIZoqkYjxl6s6RqhjhVwf/ja1axKRAQvIFa3PP+j1oPkHraxT8elSV+rjKCSI7Ok
TuoMystbYe12j6/96J7ViLBnmv8r0XK69/LsD2Tx+0wUpB7iv6YdHPiBPnk/1jUB
f17/4r9HPLbNYXrypg0vsI+D3ysPEpv3d9mSYfuEQkLRfGnxyZJDla6cSxBeMbU4
gGRnZyDQEyESitO/YjA8310kZndxBPx9dEoZsGNTKwdKveXLy5RAvOt1zf0LX4V7
TsVi9E33INa1pS/iyyoqle73nfuvTbiFAFi1u5P1D/9vPadtvGKPYyOuMFKhkNz2
Opfdc71aDJnVI1YXFhyXkflp7FCDM3BB0QZU9NlwsXAU3Jw30vSpsw6QFjeTV/Fj
7R042MnpmCByo3FnYGFAcXGtPuPRsj9XYYzyr7YBlJ2Fsox7X6KMcLCtCyZPgm4+
ogyv2Kt24MahTIYCJPGgEVehoE3iANNrDMRc0S0UG+pBdwfxlwsZ50kWpaydEEMG
KlUqYM68YovqjbzGkcHLC6iErQy4DJa2kvS/1HbeeQeVdrjy1phbtbaXGOmhfgzE
RUaMswqosaD/nrahPFFHMJJ9A5UsfNXZ+euun8WkEczu844pZnzm+MMO3/qOhfgK
gLIkZTKxFNPm+4+fPKADFzEmjjMsG+DgWCq57hvtGpLS8H1g4D77ISQCoKQyWZi+
eq+WTt+A59ybZBs1AckNY1rawcZro3aPiAdRDXxG4cRgWzG7KKNliCRspgwXO4mk
TUEzTnYHSVE6ZGnuSqQXLmq4Tz5Nph6Q00u7xq2SoUVli0MLp7vOncCe0Kz6cAKx
CBM4rAPrS5yZ/JbD/aZSEzNizMUOs+MT5B13HLd2QyF8AKDPEQbxfibmawo0N1GT
Pr7hYV8m3zSZ8FIFlzFYd15jlQ4Tw3y7ogGgHWwCrzbU1cxfb3YedGm0C2Y5Bz7G
8CrK+F+pnfEo0biDbgSPe6kgTJS8Z9CKSRVvUX2y9Zs9bxm3JrHOcL6UEm10gKCM
LCHD8FR7ILQzpmZPUQ3hf/UwtZ3DKc4GwBo/tK69GMFfAfPLzfbUur64LPyJMpH7
8qLVSg+BTGYfs8nXtSfMB8l0FtQ/PoQ4QYk0SDVaPuES17QtHd7hTEUY9RuQBXoL
3tOrh2XwUBjwUrSz/azhAz4cHkvXRH9rCp8+U9lMcm/nbgUmE4PDlh3wVH5V5oFB
1+98TY4RQL8Eztzj4cZUUGlWzVsOf7z6kis2FVrc/qYoGx2vesHgcOjqzCV3p892
+EZq6BgwhDfqBeojJxT56+tSkPogWmc807ciENNzllr/PI7ClLMgQv6PjPfOF4Q8
IvUNwY25dvfXxQcanZHlSLMFp2yHgHK41eX+H2pjIp+WlYE0UXugiBDoxNMhRDGp
qYxTA9M6+eiqfInDRsj67Y+GOp29Eb7bARLKiujwMeghNxinDXxPLl9gNseWw2IK
sR7f1RyzemmADQfoa8b/zBHYBcZyp6KhPeARcJ7ZGKg1uPlRvvze8CLNNtzHYVaI
MNzc4u2uw2gZGgG6yT5b3yris/taGu1TWCCWxxTz7jqo/IO1J87zX12xx+PK3LO9
VBZWFwSl9T0h21ibofEBrCy2ArPeBBgStqoOShSD4cf99YQj+6vsX1Ypi/RjGpvJ
J1BMs56HZFRGokyF5SVHKGXFGbDRUFi3qaCsT0w3VeReSBzSTcWR014HnOsDBLGg
ZwNdV6EBbRuBMRCkSgrMUUMF2ycaGXC+Pdun5tHiVAmDNAxrsDYUVMGqofhgzOCI
m3+MdiyAqyS3dPjxdq7oWL00kvZ9lFmu3VhtrUuJxjzkZrhL6ebKzWsXg+36Rc8p
7kHmjwrAVqzPP2/ca8d+msxLZKk9YhE+dN0tUyA5jfh2a1sLcFNfCjJUKX6bbRLj
tx1tBRg0MaEcReeE+YE2VueD9pSxTrgQLCX+opJ+vdxwiJGyW3QdpafhikmiHYh1
yl1TG9VfT8HGSh0ukRbExEBJLlPGudPOtBGSfjCJrqAuyNPxaTswXnbLh5c9JJjt
riKCZamO9mp9FG3IDDq/6T5VtcAVbzl7QwFKovUzdOJlmleKTtf0IwmvNnqGw7yB
nhC+lm0STsDqwKR6NKR05lTdnMJ7e5YfMtsemYBMU7gTCFZZW7LVhxZqM1D0xfjP
D6QYvdg/MTAICKmtfuvgqG/yVWQcJs7Bl09Qtsv3MVxTS6iO4sjuLmiqJAuHTK9P
tbnH+NCv+BYmdFkZUIHmzScBu5xFNUui+1Bd6AJa0lvukjqH1gIfVJ/Vx7hBhsAP
owH2GcA3azcfMRCaK0xUlqrKlokX7VIcBD05kGGp3pJkHklqOaorBKmEbn3S9oHK
IjMfd/71OHDv77RbJzDJHWsHdWgpVntmOAvHMdWZD+SuUr//+7hOefWvsKQgroH6
nMWaVZnK06nhA9WJ5xQu/D8hpqwsU77FJBUzMdyX3qY87u4czVtV3sYRUx5asBTV
YNB38sQOj/rfhWxwITo4ffuLdlxoawv0tFNp9u4Djygv5UeFOdUYoVWZzaY3wXER
6a3cd63VDWhVfnNep0lK5TwneVkaWQlX7GK3OuaoojgirCRyKymdilOeWzRPUI22
/pP5GdinYqdXzkuyVRKtPFiuF9pD1N3Mx3H/FmyzrOxLjdFOPO66671G6cdvLA12
AXF+F2TDLKZRtJHb05GhQp6uBB8AHs7m0vBOGivCOQ44+oQSkfMjen+xWcdedE7v
fTICMcBlpkngacxXKZieZ01ldxgTFtrJkFoU+cFsJTOu/qwx1EfJnUQlF+Nvw4U5
BjSXJOLurlelcx2LBaZ0H2le3Epb+ja4vg/Sr/eTQzoYHxs534AaK+oKneG6SfrF
DSOOtPoV3fKzf1WfhLwYcgbayrPz+B4q3Cl0MAzaxZ76Y5IAPlChqb5Ai8a3/Q2x
zAKy1bckpLVrbDY39QH0O2NvIMwZrsplvhqGh5wH3vPkpC7/2hhx5mD7GMsQf78N
N0EEJaCpMrSRq8cDGeOR5CMt1CwjX/3ZWr4iozEnZeYUn74d/C8U6gV+GUNdiGao
M4XtrD5ChrT55coiKhDsUrCFBgv1qmC2PUFquwpT4//LzDTt6e90sdFBtm2iIpf5
gPBaGIeUeEcg3RxWG74Vf3rHbVRaC9FMlIlbhWi9tVNEBWVJuUmoe4kiw5BEK6Id
LX5UJVgmewvf83OVJ9uSPYlUgSOHd0sJn+zNVn+6OxDZFXgT6zLnwg0ERQ2bSt59
PUXEhbG73BUWjPzkjl/oYQsuBJ3XO+eYjquvSz0bcDBje3c8g6BIQSZkVtT57DA3
/gPHcvfSvip2pTBxNApHKq+M4zeO0uNYlk1DW5NJ5tJZ16vVyIqidL2tfjY5LqTL
u30oHBof8ZVlLbvAbOCL/Jdf6ZhYiVSusK+nCOpElukpTwGA5T2o+j27rO0LooXl
eSGOSWioZTjYYhcday64qm3f2Smj9YL+H0BRofVfd75XnzjUU732ipWCF6nP882/
vEMsOmAXvBfjeqJF2Pf5E62OL0Eo1Wsa8USjMo9gm4nLDIDmy1Kv1rgfTOV/aY9V
ApiqNJS4iO/Hq5lTGQyH226b4es/1RCAnINGDjdBU6PUUJwmQT67VmPPGKVdcyfU
Rk1HSsjGYipROGLYQPxckzI9wYKwzHvmAyVjDRDK0is=
`protect END_PROTECTED
