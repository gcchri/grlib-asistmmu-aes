`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d0/plAqPYyhJkqzQ68Q75RBSEzJaGyBALiaFaxru00Dqx6kw1dJV78Hm5Fs5QMhs
tb5yAg2Tteva9TGa1ik1HBfxTKYkEKV6in6WoYcIHMOdLMU5facvyEDaq5QRpq76
hj3TYn9PdjzFcYVGOlC4zks0eQxmNApAyb0e8rCKOMyLuHd2KHEVQ6ocIUFfnrZE
R4E7ik2cqZj7ppiL4WAZMvDo9aqI+dPM9bFZXJK6DyJRMYwepqFJa8rPDmxcJmDs
RL2swVtFjqcwc4EXmSdYq3wB5RsIn/fLU6xAGxepEXNNH5fCHW2iTcpxOD9wIhxu
`protect END_PROTECTED
