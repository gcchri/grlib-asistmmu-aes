`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A8YpnCynnqQ6ddqiVufgRlns9ZNexB4t6FAxmKWDxql2JEs4yt0Ufx+JShaAyQnE
Nir1+kDiW54U5WlE+KG7HH6hgeeqQGvwGi6oK6xuigeao/e0c8sy+plphC6/Xw3r
i/W8wIv+CTEWh3BCoBcAvn5uD5XroUNa7VE9LWEU5TSalNOIfYsuM6LOI1bQrNsA
/vzn8wzD9Rpg6U2CQL7udsBHloTlgs22W2Fz98EojYe8RySCYA7hFx2rfYC4oHpP
C0s7gSuoO5WXequ8pWz7uPJBbPLuR1s8rTCgAhXwVbpX2v3gCjQ0KmguxbY11Dmq
kZ069H0QTIU5AxiVnBTlLcnSjavENDqqqg3LOjI0602lqQ7dRXZD61mOaqYa2c2p
lHBOLLXtUI3ZW5VNx+LE3cY/8t98PjsJ2rgBOM/R1d+c1REG2yhpKKO7PP1q2bnq
IoROMUywd8zOrk3wYUgyjwHJqffpfesiI8xGJ+s8f1Gnd9DjHymkUDuE2UK6jwBr
SwNV7rc/NQLLtZU0I6d8XA0OHvW+RN86o/t2DPrVXbIxKUEp6pj4LZP667m5iKvl
9O9wC9f6BCR6F1/WVUlcMg==
`protect END_PROTECTED
