`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fTmx5u2ChQFqxIOwdtAFYClgwmcaqCNqmKYjrImeAlqLuOYOXuWi1U8JG1VGxtuK
Dj/rTcmMcKnw6v7uG+KdL/MZhVTznagMi06I4tmKOalwE79iqjLZccYh3BfKlsRf
tNArqk9m783BQ1SsaJBcEbg2urG1vJTFmmvUHAtmS7/h8sFHLGc/3NHCXU4jAEvn
XXBBarg/odgC8O4MFGHU3jLW3Rz45Ut8yJgcGDiGHxYNp8p2/iAKp69wluHKWqKk
RKJ52IUxlzs1XfC+PerHr1GNoT1PzKEZ37H9pY4sEP1nZjeSruOXOelnh1BFNTIc
MrbwVioKpIi6qiZ4jjb3VOdLvWTVpMZDzOK1i4d5Iu4SVgiFcZ06/aJUy0aXRiZK
sJF+yavAvKMc3PTcx1xxjpvAgYUbd2zGV7qEbfaYzuKEw/MDVTGS5lIIz/nRlXL2
XL7KcoX5p6DpNwR1631kX52Fxrdv68ztnz58FjFkHhRmhGvJfQmsXfAxS7hLjdk6
sV7HF960BUmXrfE9izDE5awmlOAoB+yHFJI1M+Jld1J3PaRqa29svJVi4sX565D8
abImgLTQxmfTk1Aff8ZkbA+ghsvHEuCvcrjF22z5DnQ5rEsVJZeDcJpxu4epR5TB
UfkejcpL8jyIAjzmV7lm0LjQQ7rg9EzgTObPFqFEMeY=
`protect END_PROTECTED
