`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PUYu39k3vjCd/EKZTSlUkWii4ObSW3FpqOpPKZ1y+/fi9TQKOnnwhjdqxzlrBbhz
7dddUpopJBjFBbnz0Fgiz0aBY4TiGrqEYGp20p1hEjxpilipM1Jm+Ve642W/4Qmo
KBQYVjpKYx2uV4siLjtiKr01TgRl9uCDXVVIIeVwu/8YCzrJwOt2yRjNiQd9VGWl
rG0fh7zvF4KYEdSMGgIPF+Mt2RoIw1PM8N6s/Lx/1wQEVrEUn9a+TUCYhSgjD2kr
57VxdaTX+rDRQ6B0UIjHpPVITae9tr3t/ildWfFtpXLAWWoOqN19UTxqFGzO2pW2
10uQN4wkBNMjBinZ/R8rhg6tA1WYN66TBVH9qZtMDxbYX6psxuj168ANZY/pk4Rk
9jJlg/w9pxa8vnmsRzZdrlz5J0yb3l47uWVKQgK+WLGRHqXwsGEbI8oyxX2YQ7H0
syOX5CgS6mlwz59NWSCc7g3mnK88rM3wlp/mpYc/ed0XW71x66nlOBJDSMdjPvmH
uoAWm07FvVLDV6YoRDUooZotF9B2Un9tciMWNY7PHEjBSpBBUyKIm+8xycwzXQtI
l1mDvR9OQlhWKSm5dpZ/DVgP9reKeVpkgl3sfmJEPKOjcPBf7uJbwEofTGDVGz81
nQmK6GktjtW66HJB7LWzUOFBzbR+hcZLE70ohT8b4h7l8hTuVaAJHQGthGBLEZYF
p/SmD0XZkMw0by7LIsFrsl7JXWcSDMgaqKgMXllKXBs=
`protect END_PROTECTED
