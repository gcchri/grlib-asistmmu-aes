`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nF92IsW2NbDEHVVCfk5JyAfo2JTnKD0i6EyCfWdBlE/0GKu205IAv4aWCzFiOj4A
QEW6K/SXbXH9OfdRrmVWDfdsGMdf7y1Qklcjg7DsyMRDVz4VMDXRepNC15DL3yS0
ATktiNW+2CPuNEEPXDCgnxzNfbCt0YfkfNDOGR0DEXw7vF/1x1EuOVKq8OkknLhB
xNB0hFvWHSTYq3ORYGdjKkKUT+9eSzvb56Stq+Z8i5GJ1oIjOdvZhM8MLDrCqfnV
YKmdSfT141rNCZ73WEzJevWOlunImYuZqekRNOJrMhkK7tei0bA3zmmNuK6xk3Yi
0OcKbZgnFyAbtMJX35dgH7moEkBRqSBVUiQy6GEseLn8PmgQM7ogt58Xmb+BVru4
0O867LLsDkQLcejhcZQHe2+ZiaMxLNM+/CEWIseiDa2xEzn1FW5FL8InrmMJFxcm
SlIsXhPj5+BpGSnYaVyi5TEzjpiJQg/rpGMAicfLX8kVNG//Uhh7jra9GPzjhhyM
IcCo3KD8cR0m0h1t0lCHPu2mQ65+LG3QbaFCwYVRzYLmyf/5TostlZ8lu+YjaO7s
oj2MSffRTNZwaH6SM1mGIa4SzxvO81zPJU+x0uprYDbxNum3k6WpOHn8YrN+c4Vt
2N1pxG+nuJmI/Q+vZredSsHn8TD393Woj7yLvZkRC7eM9BZU/+S9IMJsTLPKTlh7
Gss94YaXM1dUOMvxacgdMCjtBitMolKTBZ1r3UD+G4I2OtnMxNEyXWqL7A/i/g1c
1NkmZzacC8MSTXXO8Ug+Vj9vBFL5BXvXtIBYq64yrJK7sUz5taHninXdQq/5l3/3
fpauK7ShAwPvC+cn11vWt8Lr0wITRQpa6bAxlhzV5OK5LIu5tZ7YvOzP2HKzNVhq
M3N2MWOxSEYr9PTj2uso5mc05pOgwCKEih4LZ4K0r1owNTVu61x3pfT4DJX/LZ0C
dXH0YC0uizmDq+7n3ACUnKL8tpLJXG1r5guqzM9Rmp19h5uTYB5SOrxDFKIZiJmB
`protect END_PROTECTED
