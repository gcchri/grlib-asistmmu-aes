`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oyUqRSMyPnrxKSAZNiqqr89GNE5aM1EkqKsMYO6GTLyMAabwVs0HMp3wETDmqcbx
nJwYzuZGTP26+Bm/xMzemocfNg07vM4QXREwq0IRRa2A8RvoikOlD2jPN2ab3rz/
fYbAtWunlCt2v9iMwPqF7uaY9jI6eIe/RGq917tKGiZICY/YvlcYf3KifJebq32r
XczRTDYBjt/3b5bh/Pbs3BGMTK/bG04jDrVeeONvXCoMbytTN4JPU028PrzyXWqp
Opkj/AambUJucpRKc8mq2BE47NBP+hp3IIjC14XsFTDDI8Ev7jiJwidlwf0EJ43d
C+h06kXrIaw1F9B/EichxiUWVI6WKk4/VNZxFvnl78r9cpiVUOuyGco880WAj5hU
yHbDcCenJrfFFst6TKGbuWKBFoCsHi63Qmfct4ZuiOe7N161BBkS573U6BoJBfGv
VqC2UI9pnrmIpj7inns+YqqRDcQcy8uu33YBliKpMhP/XNwr5ad3hcahghXSOhhw
6E+CLZIJL1f8J/iaNnxb+LN0PkLmugFZqhdVD8FBETrw2oJqnMVC1pGJM0Hd+Ah2
TrzKsiVu29bS1v78TOKdAexD1C3ki3yVjj1HCJPlg884TkB9kgAP6Rujp8EtY6hI
DlOsJEE6Aq73CihESyImNPdgSPeYzfI6vPbxV1MMB596N923QW7U2htmNVcRrObh
mJj9Z7tR/ayzW+j5dny9DlFuzuyrxFoIF7e8RIWqjDuIVMIuPbjv+psv+KhsE4rq
pZkfn8nioQ4lx+YoxO0HHyq/FQy0IRP0yrpJRcQTUA0zfOD1ODM4W0v0raaI5xMq
YEkbXqo5KuqjiYZHRYSWEbiJPKTDdm0XIdO2m2/mmErWfB+mQS7qQq5o6rFjsiAN
XXO/1Cmy1cPCk8+baCxsMwrlmp+pyb1oW3KDeUFIrXBoXOTdXiPOeznNmxbs3uY8
/EwRVzhkVh7Zgn0HTIoBASO4TEvDziAuSQSEkizBgmFd/DHcQyk3+YLdaNpp9LbS
qqXmvupEamrRr0H42ePTEXfSDMSFdoi5tbhw3wptL5itG+fgRCAHUiyOgAlDkImU
+9o16Yii/jIBJVbnQoP+GjGG+k4pyhMjZmnTG96VT9EI+mBNhns+/TBymGUpBF7D
9iKceCIaO4rJmmsDT1EAFB5iyijtG/Iydw59DV4fUM/NnWPU/s1vRluuWrx/cIuM
0bn9cTxukY+SiKikI0cU52sDfTVkfl+N8tnXchjzbOmjw4/jXqOaywVG3hWlzBU8
wvDQ3yB9744i1zS2J5gAdu+1XAzLfzl4kSgPNHbdMIbbugXI//DcTfDoHcGBLJ0b
B9YGFHKV2Oqr0c18eclV9pgx8jLnzJk9/l5VPH9/3zcwrzqEMTA/ef4XcuxynGmI
Hpo9Qs3pQ5AvAcDkJnZDIi3DRaDoPhh9EM5EVvwfflm+qYfv7ENJZyR3g+Xl6YtA
HHj9loZkzV0bjB/trxzHtjyu41ZdP8iav7QXg5NcbEM=
`protect END_PROTECTED
