`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NKLwOxu5C4HQmZEN2JEtCsChjvdmNYOxH5GXfZxOwzM5OVElfMSHMRTKETZWOH26
itWafrzn0Gsk+fSUoKNs3PKJodTVSTAD5uzYH49fcjj1TXe84uvkKrA16/KWHnTb
W28H+TUEpdD9nEe8eCkcy3rKYAHmgibCMQKynD9HK1H7pQVAhyadIgJ4NEu1D53c
l5jdnWE3T6/ZOspcdbd+E2qIkLJCaetrc5g9/k329OQnoLKaHPiqx2ofJhOZ9BGE
9JA1GuKlUFcG1FKG/swcJQ==
`protect END_PROTECTED
