`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SIs6/8dldyhVUtWTKADmscIHD4gwnxI+kqoV10fBBN05ZBUVqWKUGD2WBZwWFuVh
Kq707NRjGSrHI9qU56CeAJOJzOT63KGra9so3ggYiRqcq5pz5Ug3U+R5hJQQ7Osq
1wDPnpaQYGoxfCIFet0NylBbvf9KjUyaL2TVaMQsP66bJGAx+mE++XNwNUue0pdf
gLSrP03mDeM1aV0cDrg6tPkxL9XmkgcwggyF5fYhCUQfUrfgzskLqbvgI1M98EWF
WtTW+rfcwxo7biBYM8+ig61at1miBqLLA6AsdJWSh5dzUaaes1GdOtThUU1StTaP
IuDY9bv0SsUK53AdqrOMb0Ry3OF+0mmjYVsm/bqTK77DxhpLGc0kiwH/BG8l9VXt
U+seh43XqW2lRmI/vFX2mufubHqVzJZFyhHNFShma7jN3ObY4hXEnm52GQn5nUMt
SpojZCMmMnCM6LCpjdglwop28HtM8rs82cEL/LU/KB+ugZKE1EwqUWBuLugxv7nO
`protect END_PROTECTED
