`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pKcCxSeWrYvHi7r+FBdGHoc4Ibscrmp03jRl+a1uLm5yYp/OPSdEC4Fd1Ril+DTD
3I3VLbl8WmqeJJG3ansgUZvt6n+j1VjgXRIy+WG5tw5csvCSspCbvWroTH9h5w1W
KOjoWyuFCHOIWFnI8lF+mgHvQhqD9j5ugL+uB0FgIOg2W9utN5hfxDArDmOYe53x
rjE/2W1LEv12Ke4r+UBHTixvj8PTSb3BO416t0ghYzbkKAb06ZfxU1saEkmsCmqD
3x+Lvnex4j4Hh1e8KCvb2Pa0kTY8WAbcqcJ1sAKs0YZQW7jKftXySW/+96AaXvK6
SZFTC0ASgaNw/cllwQ3jMPP1DNeZT+sNo8xcl0C6cFvqz21zAYdWby/KZEZkG/8Q
VqnjoYo1Onj+h0J5+r8mhtrUDvuiPMlhIahbFGEacf5pIQIOMj1iEaekAgPuc9xX
N6Ub9eZx8gCTaZ8tPGyyORmrnBr6y+0f97izJkrhK68oK7sdXGunpfUiLdz1JtqT
/bEiMR9f7L5ZGKRgcN5gFuHfVfmZRNnt5inhhs9ehcBk3ElKckXJcYor4TS88GZf
lHYFVhlzno3bjNeiO7HVnTmPqdJjK057o1pg5XVrKzFYY+3SIwa3XgyNCyVTqKpZ
bjQLYW4nCIBnBgCv4M7cGyu+EXcS4x17Ewhk6cvTYfVK/ezcSGZQROs5+8vzmx+P
`protect END_PROTECTED
