`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HCMQ752TW9DrXdlE95NOZFuDcTGog0cPx/00duYCLGotP5XzZzsn48XndGpK/atf
dPO5Rw6CLSd3aEzS3Gp+szHtfQihsR3rb7TTd+d6Et8GhcjtT190jt7s+SLNPLmY
IEKTSnF/C5XUA/moRpWzHxLG2h7lumOoi6lp/w1Szo6yfWbmttBqZ/tH4Axfl/Um
rhgp+6XB511SCT8kQScfvD81wFrSeV244D5MFT/PTcxp0IonnvLFzciThirEf8zh
YdA72lSuUgysFhA5TWqqU/pAIoT44bJ7ylFVr13Nye6Zjqy8GWaqi2CbsRJQF4z5
Pk8P9SX01F3UoXRvC4Dd4WNT9k4Ip2MRWqRnJ5KYgRZ7bl+SHAwqy5BlVZEaT8Jz
gaIIjfbxORYWZsvPxFuMV5Bxl/GTjqUCdWp/8Vx8DH0HVVQN0+QkdwQiJNQr5zFC
ZMjtG0TF+PWrL4knYUGCVqYq6xsxtZZWHX/EYe44X7PDuoCZtSbIunSc4K0IxZbg
S/POLbSN8Dml1EQyRZLKxLxXKKqCjmRtMCBGWK05xUhhuEMX+2YY8efPZYp9kbDp
Z1eprg+tSTZx5XJpSBK3Ag==
`protect END_PROTECTED
