`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
65gd4n87QzZ1blxTVzPLGJmTCz7nBbW3qhLqAHTEy+toMVA3lY27UbokaHlMDTE5
t2EK326ljKfaP2+HAhe3BKt8Fe0VwcoTjRQqm8tB/KFzvG62A8Xs0b8tjmfWDCga
NzfJM5JdiycHrxIvnCjs4hyickbJkUjnxfdoEGP2HDWG7nuQjS1liU5qyb2xlyFR
w+LJGHt487+qDQ3IHHTboLpgrn7Y/M1Nt1Y0RnEuBn/XgnDluZ11dJeeQ232iGWX
zbdfzNUcyKE7H4AvFuknbafwCoAui5SqNpnyqjiATiBqsimxpy01/fxRXU0dvFDD
z8/6axij8zTzbOK41k8zPA==
`protect END_PROTECTED
