`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xrI8wSPytN6Mw4/mjWgEdACiTfyo3LBtKosD+kRaMwt5QQPdGau/0QAP4LQmhXjy
TCGfLbDpOGNPxaH20tY94O6fJsNk0SCXO/M29ThLNlF6Pcc7zKkcaniSCFsPwIBq
bnd8CGnmr4Z+5YHVhOO+ca4LUjN/gvmNlHe9g2SqFVrGXeFfjoFzKmIiUMRhwT9P
8RdBzjs8qG1tfpD7HVTQ6Jo2sFT/3AAzvepkOecGLN+n9tiWwPkPCbq4EP5iILg+
R+20t2stP1jCeyhMW9nOIS3VpEpZv9SY87no9Dx1Vme+sc2qyP73wbOcBGGMPNul
I+ptnEStuqGJyX6Y/Hu1o/4jx0eRbPr0l/+0fu2FfSnCCUP7NAn3ScIfeUCd9001
CgmkpfFdiZ8mW2dDLAR/SGpk7O7y7JeFC+ZtOpGYzmEG0ezGjQIvwqFTZVaKEyol
ft66n3teuz+KCOKfGs3sPh6zSv5z0Opg+dmdlG5uwNKNi4l23t6wteCjeYrwQJj+
suqrW6crLsLvush/tv0wNUYcLiM/Uq9XpslwaIvcGw93pqxx1/sU23Wh2cw9jKPu
HnF2MW27WmmrvBeLsALJ9E3KD5YBfog02xT622PryVPUkOQZDVdlfrTJVXPvOHQq
Z/fyVEIZy3Fha1h1NhWZ7qAIjYRsIeEvh9M8mmrZfnBWLTS6MWEklUwl5bbRZHLe
v+Sa8hYHy2sJc5BYgFqSbe0wrL4SV3fQI/qXKnyt4Rplku1pccmAQuNPMwyt9u4C
4Aew6Va/2Knijbm+RcKxPakMY2+6qLi8vhjeCQpU3O4CqdBsndfG2Xs6zkEr5W8y
AuFFbm1f3xX+l+sUmJIAEpAKIYv3UG7QMAZY4jYXKbzXEAJHrFAgJR3/KSiseXA4
ncxF5zISlJnTH5HwP/LpMJMQLeGhYhLZKFQ5Yd4n+yg99nq/jZM3L0TH1JZM1mGE
TomWHX2TUrSTj568a3UsRU/Rn4yZp7qc6SLF/IWnwNNc3RXyg66djjg4d/C+l3M1
2hFOrn/D2gYM20V8KgVaLihyJz24NFs8bkU6tvttkTMws6KUgBpsV7IXNW3Xx2XB
YInR7Oe2KM1UMS+LMf64HwyJp1ds1diNqCn9x8Q6/6fO/U6aO/igNDqk+0Pnxyd3
r9O7Qc+22OK9KnCESngFrOw4tu/udpHM4p3KR3Yh6pZS1JZ/mDbfJSRfGpHmhGeL
zzKUhCRHHDX/23UXBSJg9apb9qYAqe4nIaG29YmnkG9723POS+BqWuXnclrkKh6W
QqCPP7OE6ErOFtn9rRPpQc7YhsMZMybgfw4vuxlkae1Up85pBwymHPNGPzOSIxKH
S66PJQP1F+zI1xONRlaPDEOeE3WDsrC0HmIDt/8C+71mrB22ut+92/u+zPvABySi
c+wU9Ljk8rYJiCSMj5GLJujGSd5w7/41iF2ooJBmuVWGoODQzF8GQoYa7N6kRH2M
hIpK2Dmr5mkuhUF7Nn8zqbSAm4mP/m/EQhtSesF0PajoDsnGa9M+llndAcYnovuz
6LA6clwYLbHGXsURWdNrhw8WaLFmPgMg92Whicoel3qvzIfM1b2Gd9j8ZY+9TS0k
pk0Qw/rBGJ/hWn9BxvulR9tIN5RANsyGVaC6SdzNCtyjvB8xM+FfTe4OWkurL4r7
ueTgpFNgUUzAVCtnkNeTfXJkNh28hlNuvUkVWJg8D4mJHReettTS4vjQzyTajNPB
wa5hE8MVGpAkVi5ZowS5YCONfiO/dU7izhhv2Ubmkxfvu/U9RrNBWNLbpUbc0G27
gp3jIL9Qxxw+tLhgRGllZ7ZR2+DUvvcj8wHZBfBVbQFNjRmfVMv7yFmgZX5a6TWw
r17lnk0Xp6p3khutxZ0BiaWrXmF0vFAeZ6XdEiDKnoWh2qgpSqD7JKdOIDtMzuJH
FkTJ0P/Ji9TrxGZz4JrmQDElxBZEBoLCn+LqBUT52NoSvRgcnRnC2DEkLuS70Zl1
KjSduxQLNWON/IIISpeob+oIiJFLyvtYevheDW1wVCD1KJ4hkLxyjpeEWBrqxYzZ
hwgEAheNBDPL9Wt3vg1qCC3bjNWI3CAFG2A/uqGNwV+LRYAk7IKNnS2NqvHC3yFz
WgVMCzdERPgFIxr8dIU+M9yqL6D+5YQjrAlynfrhFdNbiaGzfACD57HUuezYWddH
RRD9xx5UzohuJstnn4u37zMorrJJk8k8U8zJYrMood+wT/fDDzLLn17Wh11U61sL
aTxPWna4RwieAoNmw6EOuehiErHqJiiwV549/EStRVIIGSLR2rsiBbNJeImbBEnE
atfuIEHFKZXLnf20CpUjbI9pp0BVmMW5QlDFMSgFUSS9xXYiCd8vOzgaHqqyL2wr
JiDH4hATaP/EGS2dh8G8+4mgh9fu6151OuK7ZD1fo4Z5SzkPI0aMkZGBiudkQ7Xe
vmHnORao2R+miQBZau+tPeyigOrJfKqK/br7XLQFp3s/fe6PLxrTNoiGvv+45TSi
+beQt0NrtYcCn+iPv0HF8ODt0RVaJedrE/5Fv7LKfqZmp98YeG+D183TWjBf294D
A820XJE9nVIpMplzdO3xeIYWBR+OOc6JtR7am8of07pvPSYWewfxWfi13yEfDJHI
sIr8DDdyoTE8JsKAnvpqI66Vq73Yhcw7MZpqtCgEY9eCd1b/CMW0Qx6HT87SBNbd
bUjEPRcma6PKLxq17GVYWsiDmzeai3WwkqMOPdPWVMn7/GI1+6wIKGY6mk8zIrYn
5/7k6wkeiDQNfStWfNQ/K5sDRSiWDcK8kkokeL/mSgi5bl3po5/BiXBET/C9YT9h
2T2PJeQPOR3OQRAQTwvwBEwC+cGoIYHphVOWx606P4EA0DWMQINGqlzUhrxuQbCJ
SuisXUAFvzW/7x7wSk/KJ3Y8nz1UC1Pgr/+/3niuKdxrSLyNXVDl4WfVwvZiNo/H
4S2kXuFf6uBKRW/EfPsTZup8nbN7gB0RebDJxw6d1sHmi0HqGXbI39zhu2Z3etCY
n0h+g747BE6DXt4TPUXw+PFxuZXgYz6fpWTfylUAixdRbQ9QQ5+GsATenNNvq9RP
ypgC/NdxpOd+jNTs63Y1XvZc68fscPpX/fzc/Gxd3h4/68Ra+Lv+8S6iZ1iPTh4x
oTgf47ay+fCp+Zj1OVylnIk5Ayy18bcPt0iO4K/6Ml4cicYaGliNkcapkNwlRxsa
HZBlPWcHrY2aB/3MT+x65ruppWk7W6/GkgQYqGciLUHXJcjpAk9xf9ok5UEGA1D1
PYnNiZIoJG+wxswETSIS7TGHIMMR3YzN3Oi2CGitd1zxDWfKmR610mtKkoqW7rLV
k3JrCF2MRYstR3U8ngcWc7kOw49yjoq1LC4sBPfh5O84P7nHzJffsp0cJsMJ9pI2
J4BqiMdU4U8dlV33jldDqpjOkbFBewOxyshAF5xm9JtoBo9z+cnSc9TNrsHGUciS
Ma0lzvXlNL9U+LWx/1Z7RISeULTe4ROfC7EVAbBgYXKM/T0HfSbaCym07BoKjrl7
z33t6HApbbKRsy42pqU9aXNyVxyCI5MhZ9HsVeS/mihWb74nE21IGIlJSMehRwx3
PySy0a7fyUx9CM2/Gp42WsPi22f4zQf4mj0zflccBv+5lIVRPnz4FkqObnz+r9/y
3tE5G8wKeB84VLMpiCPmADYpLcnjZ5tzFuR5p/URZ/K9yGc7yWOSwlY79WPuXhdB
+TDH2zdDN75PQBTeavYhH0EmIsMvd9HFcXsYJcsaXW3W47pCKXQ7LS0rEJqmp6/6
4gCgBEFxddt+sFP6LS2LkxrTnudq+nC81EJ/e4asvTbpswS4mLKpGYU13vxZ89k3
xwFSXrfa1XVWJnRfDrO/Q1YUsGhZgNHiBJ16YSM/RLvY3iSkLkOC68JtYc0C9u2l
EsKEP4Yo0PIiw96wg6JvFTWuUx/trXEqGZMVKcZBnYrA1SoP/DO2xoMjqRoae4AF
iBXL6LhdlkESUxMmtwk7j0dVEGEdIw2Ln8sS5DMY7lgPEDq7TD0ep6VAchnFYdnK
sK29VCj/j627PdcAxgokHpaI0Bv4oAD1N7KafIrwFGOVwYxGorOmYCVXzpwCfi7S
kikkoBST63sPTdUez9DLX6vKWovEZ020KV7JzzRF4XMuZ8e4WMuj7sTV/ZWr400/
suxealeA4CNBpHSPLRC/h475jZQtg03U7ZLpODz7x0Cf8PJs8bZ9+qK6nBfW32+g
xmQTkywi+V2MVoPgX16+vzCsKBFmv2RL3HGV37FAKJ4fQvrqaHZE7jwdn+fRP8nd
KfyG9hoRiZ++oabDsQkYV+TyHoWZqVxLkqK/62Ua6iqf/bfUsxNRa9258KJjkGwF
DsfuZupoxW6aPySKMrrTL5zfC9RH8scDznrmCvGFs/hQApHNkkOOOvSAol/fmxlK
vtaYiqpLp9d19GLcX04yqYTsgQc6k8ifgdlXZLKeboOpZHpcUEY+UDXICqDI6D2V
S1nW2IWvU6s40wx1/nJ3dRhVCMGfl7bEFuIk1ipXAjOPA31RTjRui1D3mmuabd4r
QDmiYT0n0xL0v2Nx9+8+2qh4yA+opurX7ZMX0uc139+bAGgDjyWQvk9YPDw7gNqf
EX352DPMqTM3RxeLt+isiToZ7pGz3V5MJ4EIF+gcpbRcC/aU+Fgxzw7A8uMco3sI
Jw3zjDryhb0DIvbxcXDtc2BThLzsm9o+v6YMzdReSK3fnhg3zrUhuXvDEREU8RF4
1xPYs75/DscA8sXyivSfhE4hhGH/EAIycCEElAgTHDlCAGEL8zyJeK2+7fNGKdDy
0pPVlFk+Yw8KN5DOlZacovdhDL/OkvDwXPZKZDCKsOPf+nO1r72fs0G6z/j5luWZ
2UMFctiKG4KHvMgSIf8+ePED/BXtegg4mI/IUZfObVaUW49f+Ujm8Oe+XzBAJ5Z6
a4pQWbWliPVuxzaodYb1/P6610Xf/4G/UMlL4B3Vq6LTBlUxIIJjaf1mjyQ2x9AX
6Zg0BDhoDHEryyIT9ABg2dqQcrJNsk9JMtNuxJ9j/IAHf64YrO0B9aF6ih+kb/5q
zOnlT+LR4XG/HRYwxn33K2+ohsQ0QtXz1ui/0ITOUxFxN47bygWzpop4tFotrCp4
/hEAP5XXb7N8yeTBZ1gV2OcYp25wIjPleasqOVCSMryTadMmyul9x1p8w0E/iCi9
nnQJr7fL7Bs7Gv7HWkkv9hmNpDS77uMf4O5lKi6vmnnlY0yR5emPfL7Cw3ri3F2M
AwFxfcnILJuYxKEqcBn4DD6q8PFr7vdKmEOfxLc4rrUFLH8VMwuag+NnxAzFfCkm
pGDY3iEn8i3eZMysMKs5drgQc3DEqHx3fT34ZYxmtz0Q6uc6gI6oOYZaEvJD/tVv
0djV6ilLVUcq0I26DoECr0w4Ozfu+ImXqabWpbQI1UCYTAZW9aiJPS1J6TzBNlEy
1M8qazlnOPkNJUFei1xs5OV1/zpmlxv+BIhrarJdvd/sa/lRqLD2uFaZhQieVPE/
xAe5SG8loWQYSklOPpH/89N/iSeroR7R2CzpCuLvCFuJ2QgZY+W73oPuhr+czV11
aTA/gl7BAc6E/anG0X4HfW44LFo5+GySrRGnWbnS87XGte9HEtsPAnAftiaug99x
QG3yGIiN+Z3T/svoB8Vz4nYB02Y5/KXjIxhDJ/sN9esCQ77u8jjjmxPR4lVdvI56
su7IzaaBAqu533vfJTm5TNk1lMfCI89CtkiKSiPnVUghhyDTBmaSrIOTOpV2SNId
E+Gzbtn6e6qzV+ekHPRGqA==
`protect END_PROTECTED
