`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wUflalFIbZMVw2gyd4x9gyCrCWtwV3V1M/eQq+YrfKvQLowx/aiA65JkdkckRbRI
ebmIOvdcnvsHgtfYJeXbDnVIHG8WIo+paoxU3Zq1WnU+fEYtjji2itZhEzB3x8nB
bR1aeO/7jniTLTlGdcGBhyV60ftLQAJGY9hoys6P9DyiL75O3PGuaa+SjYDIs28L
362981+bZmUIwc3gAA5G4adGAEM0lG8ydPKMUiAPO0Qc1uuDF17sRw2f8QMgJO1+
Es8v628T202TnWFJAk/GG4AWk6VS0uIH26lGlOtO7rU15bRo/1ulxekGnyPelw0V
`protect END_PROTECTED
