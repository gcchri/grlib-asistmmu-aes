`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9ct1hhFr9O6FU+PyhOHz/yK7LlwlnNLg6RfXotn4B6J5/n2mOdt395swS0qCaU0W
kPFI9mihcgwrU9d+4c6JPxF5V8wV4DRzRn8ILOxp79nvJ9vJ1XQnbUQfRMdzzMr5
FM5tRHLJ9a5M2c+Ieta7i8bgPy+t4nUuDhlqt+hC9pDy3OnwPCXwY1CaEpSdNd/V
XWBynTbdCHmVdwmsWaTsc5VRyIxaPkeugcJSDfTpB/CJckr1APSLl/E4fmxRQ2H9
`protect END_PROTECTED
