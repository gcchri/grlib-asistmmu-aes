`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
etLqssqj40FI0wR7j5iq+wH8Z9yGPcb4HEyzEeWqElXVBNSf+a4hrJ+799+F6k0Y
97Ufzyhf/mKrEC4sRJWVb2OhVQls+nwhQmcv4ASkPlqBbmVZKYKosUyW+owGVXKo
FKeCT+S4GA+ILH9SvRZFWWVnw0B0wPK6AgvIFWFY6FrD+7gUMMuH0b3SG2Grodu1
jxJL2jdG4+7xZ6xvAdfnzX+Zm7MS4Ia4q0Wttw1zwxpI01/ZxMfrKl99msLGPgLD
qz9KK1n8U47Qr2rFpaqP5Mda2Y67D7Dn6P0oXOD/CNgO85w7an3kTIqzlcbsvmbT
XKmMm/p46HMc5kN/lPufmU8prIg+XbfJXGq2TjuOBRWK74J7xaOp8aMgRi77C12O
LFK/ZE4NGBhLGVNpF5ZzU6NSFB6RJo6MpDdh1IE/iuk7PYfjXnxWKWLayVIXcmW3
5/ZgIITF4Y0QBnALBjBKhlypK1oj975HKs/IPxzYFwEi5DThMpEwOR2GszjFU4lY
RwSataR53/c0y956Y4dfxyuS4zqTuKOMpfiHjBITgwVM5F6TKbVb3dYjyaFg2Leq
lloqTYTA8hZwa/YdkhYc62MX9MoUYItEu5D/2ZQ4DrP7Of+29l7kOzqV1T65pSEt
EI29QYZky/ItILTq0yl+ECM/P3tBKe0V/oKRZlXW4d1MFppam5rawljYKnow7Plg
dQyLEbYHxizJY7BYr/AR+IU36rN5Ez8YRz6cTVh4WI/WWc5UrS6/3BOwS6aTU9w4
E7pBit6uNZ0kjMq9HlKrxK4G417TcifOUev1+5UGXRnH1ttjp4RKuCPC4l68mWGR
1wrQ0Nwl3UWJE2tV8+KRaRiIbxtS9gmcnPumRMMU7Ex7L/ag7wZiLVozRKvGcl0E
xsXYxUba8y58W+CaJihdgEEv+3k7kFvqQvgFyQH4d8tUBKubUqBUqagR/BthzyaX
`protect END_PROTECTED
