`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wp7X1BLZ90XSgaNTXEgyK5vC0IjvCcrdjnMdGGnEhYJ1tcPSQG+0CCm8/9PJz/2K
G8PqbMgZnTSo0+JhqPkGnYZ4F81TZ0NODhtWSNlcApNDrboz03xIkp13rmeEEJbc
TypiZVO44BVXPhhAwgW1SmlPViwvRDxFpMzYAVspe4LKjDlbOs8jqkbBkamhzhDP
CVR373awBCkPSDY9KhVWJB+ni05DJra5gIC+AhIlkCqabCAtwxpY8Hk6fQgYm4WX
JNpSPiTaKxjgow2BenOMxtobWvzvkK9FWobeTNHWDCIfGBScRTpeTCeXFfTzdbv1
JwFexeXKQczYR3IGkaCdd9rnzfz6eGdF7I9E+A09BXZt99K9/idfjk8SAc5KgPaL
`protect END_PROTECTED
