`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NQLFDlMbJVom2klhZIdg6WzCkuzgH/BhRiJ454BVGTb/aiJzPqZCinuJXHt0Z0Ut
N/KmFn/UqKBhTf8eOZZWWFsK8XYwA4pxaULde7Shi9RTqHGaM3rl597FRKEJjOC0
RWaA+VTd1BxLSIEr/IDYfAhbmtzYIO09wYv+cfH92NJ68ebA35SVJZAnUHNMILms
Qyfx4OUpOf4jzesFveMogvMGLzxjnG2RwPijSNlSA7uEwlZ0kLjtjEdD2sw+2FM/
Ly/7nr72k5NENaKfK6cCt25Vz8v2gy6MIYM0nHLo59zwR0qmKTYSV8j2wynDNL52
iOgFLBySZtJ8LRO1nb9l9+jLO0TpEElIwUvW5Y9C6NzgX1zw8Fc23aAQ/3FAx4RX
NQKr9EnR/VuRZJy5paVdSyqznrod8e7ExmyRkDLtpkP5YIMjRo+cjjYFM4I5LiFT
8ZJJd02UqwjRDihHywIt3I605SUP1478l7ATzukNxDUZYcZNtKx3mUIui7ldcoVS
7I272HXPwxya72TY9m+RHiRSsBiN/3fOUXj7WwgwxzQEMStJWSWtHkKKlCRTa6rm
gat0NWZb91TocAdeZkZbqqqdGOJAkI/eVHLa4JX2mI5HgRWVjQ1K00saNqM5IJFI
fJua1OdTkGnYuwtSBI6hrZnwJWm4halRgn07nw4R/uJYOu/vuRTfyBOP5Sjoo7BL
4Hl3uPQDg8AOqae/V9xbT2ADmEIXWICUbR2l49Fkf0fi4fh5GVtt2htSEKzqeWGb
Cw+gTOYYgwStkRB7qKcyFoE1DFntnsc/g5KBJC2BGEe4JDbEyjhbSn4He1t7hLMf
iqIwXHej9tPp93oSvu2KXUw1DwioKYK7tvdDpuKG0iaj8ds43c33rbU3CgddLPSW
ba9dmke+nx0saFbm/0cJEkFSUgTQtQn5PH5hIoBBjOjTXr+jeQoRYroyrC1lEbsy
S1/QHJmRzC9GTvy6jGbHM5sQ2+hzwXn5B7i6F1gJUgZ2M+lJa1m9AwSj5hIbMudb
AOtkzrLk60oLmrQoWiEfK5fFx/EI0U8nATW5q3arhvNi7CZaJGzTboJKjGhidZEV
RIN/4dwNFH8FosoWzF+VErCnXD0BWZ8rNIuH74kA+P+DnkBnjxaX9j/zftrmlJpX
REAkpjbGYvxrNndD+P+52saNL7No1kYe4mr5xk1kW5HICPbIguKO+8GuXui2OhPx
lpfVW349qADDglh70lfehPpRu/X8j4KIGGtkV8giGtk+aG4mtzrJC8b3SNEzE4MT
UHPa7UqVBRHeS2/haN793+VYr1iP7urQfUqgBDRmF75JzdnovzcXUvD9toKW4vxh
k6bVzsw78K1cqfV6qhrMwEWhhMGsHopTiyEssDc1o07tFWUMFtVwcirOUrNCQj2j
70s0vfDKh/hbGo9wIIe846BD3OCncWHR9ZH8e7KzM4wTvnY1HSyuQhnEIgfvM5sj
M93fMNPJlpXqD+aocuEE4NNLajWbkjjpK8GKJ6OJ7I7WStmMkBG2qEc8k+H3MXcJ
wL8DoSPXAURoLSRXBGXkAxrZsgk6eXmYDOTrIfRJr/HZ4Gb9Y9YbElSymEU5h6rw
t6GJeR5kzbF2CvSXpddjYCKR8rmJ70eO3qWKMJxp/sYioEIyDJmxFz/i2t2acyWW
4F+SBXQfGCH+bJzX+BVRypkxM0rgCQhF4dfjzHdsqzWHxJJTLcUfAO1dhle4BS4A
fR6fvZt11pbAIll03HlObfAiXQBgAnCCkVfR2EduFuEXIbdOlO7aeC6OA8sTWAit
8rNrv1Rq1hQMqPp+tonZ2X6bwvJlzeHFuxaKnbfV3mmu593zJ02itIJQInydAOGj
BVLdtjS6jEFeut0PPpmUHYlL1SXVUJDzLBpeaaaMdJQTzMG/KWonaVahPf1RYi3s
SxGMa7RmmKLPHBBuSOtG5ItjtllwVCCp63Vzv5SYb8ofPCFTdngelOqxEQIATbM3
C/A6eyDsutMpvbYJdTxrazqOOXzRU7jL46+T/JBNETOh7ugxhL4XAk1+sic1tgah
8qZC5qzyjhcILNOscbPhhSq1hiA5Ov+vxslk2LgPgIaQ5Z8poCn+3vBMpSLkTBSH
Kl5ZeCJQHJjhNFpxVQmHfNHwCuzx8PKGE+u6ANIQtV+/JgRS9q12zcntQGgFcz8U
taC/ln4VLl5bHd6NA4ZlO5d+0hI/EIZdz2tp6c+Zb8F7MFpYP1cshWpdjbevT9aN
BWxmwTNrfj/JAqdQR3IuaLv2BJ0y8Yglnzi+L3Z9FBJjUM0dH4uR2AJppc3WvDh0
HqSe9OqehOXcu44S27hzuGFm4Ikpvzv0RTeEUKa/nRCBJei1o2JV+Kdr7naDt8ca
LzZ8CELUolgkI7bcwUi6UYHttktVekOxKeFWkHjFh1w0ti424JTgoxlutoqfMO05
8D7Sb6iIP9DmY0Sta84v7j3RlZgucvNu0hJ+g+7kJJGe3aP1wjWwtHwio+Cy2bOc
wPQw0vpwaAmDp8psHV1ts4fZjkZke84rsNUFkDGa4k99txuo38gbbhmxMsfAySVn
PmT5bwGFbkFHG1FmmfSZyYeeq/BDXjgM2+7/cD/dbSJrch0u8FXK6U4/cVQxbEbd
akmzGEPeXNlqBpoWwp3TBcXPMWoQ6Te2/BRAFlIO/YYPz0b8bw7LAce1nq15QQpu
i9VZQt5l3KFMHjBBHt/Kb+CNQjFxeQtjTEFuQrreAdcBHSrBpdU8sVqlU1pjF5Tv
E+1WeBN+eoqDlUSZ2NCK2QpOTvL/q3nZIPF9fwHPPLqmUdBQcwF+Kl3aVUb48eTU
oDVNmBva7Z/y55KU5Af6PDor5s4tnZ7fbFYaQO3Fsi2Dcb/RRYKeUtoQ2PFau512
kGNnC69LcsheL3Kckzvg+ucnXAM2iQQfOci85mCCd9nlC3z5NzX9ANkN1wESx6yH
Ck9d1jCzdHdUafUo/fvtz6teRQ+4iEhIVVivO4j7ET4r3bqYEOX866BNLypaM4YP
h+Sk+fZBofC06S5WSFXaVmeifQ8hERP/mWcRLxUW73CT5XHMmvTcTDt6QXdIGipf
y1ApuIElBWCPiO/HPfA3zoCE1o4M7es+gQBTD51R2gMz++Sr2c+4QVAE9mScDDeo
UmhDPmwJh6zwoPYpmY6Eh7h7cxXLUcQ66SkayG7g6psL4/KzAlfuRlKPF7vtuqZw
7q5rM3tkM6Yg8UGBfSHC5RviM03rpgMN5++A+XADQOh78PtIFyTr6wylJBHQnMfh
SOAkjGA1cN3QDuJq0cBZuEfp14Ocl90xuBNJ8zHj0aWMuwiJkGwahOJLGnYgOHvy
X1Gf/z1rroolteNzqnzSyH/SqmrBlQMqQLXq4FJWuwNmu5y3U1xn2+Ygb8mCkXcD
BFUabi04sHF2hyZ7aKyDS5esoPgXkTorV6Mpxelamv2RPniGG14tu7/Q1bajbQW8
ZhbRv+uDpmEU3QzE+qLHVPw8V64pwUfyIeNqC0RnpU/a4O070wUOkSws/gVr45xs
3bcMe2BdD4d83m6FmEgja5zTQo+r3Mu8xAAE1VQhe1BNkzJirif8dxFxHGTrgrbj
WyGe3AGv5RxLMWWiUngkH4sQQr+KGX42gF9szElnO0y7J93mGWlcKVLXoecF/KKm
zpiJtnjZ52UW4U5HKFeNMSeHIC71oSRxV3W4QwNtFixc4ufPz0wjLHiqzcuHF8rF
dznpv3GO3U12z+LN1DaSe/kr12/2O2EpKKxIyRDe7BSc/lQOBCB9B6x1fj6XoEfm
oIGfew6G5ZmQOvUdrTzjDJxl8q3YadY1yU+TUIGIvCCp/0oWw8UcNcfXMKaY4+sG
5xFzBSqUyZsmnnGNjR7CZ5aYzJGB7yjDrYoJPvfqqCDjJ/GTz7zHYXPbUlz+cpXv
/z4kbXrGiK7Q0qKS9e8Gvz//grGlX9JE8OptStU+sUEQ9R6HOLDCzv1KRQiWJt2d
j3syscRyw0YjkVQ36TEDNFiNCPql7VjwsFFTHBebYp53J6T725JomCi+2H7kzohS
Mx7xPSG24y+0yg8/QdzJv3L3f+ZeEFLXUuX1wvNt2wmjAc7abXrvJwnFdAaFNa3B
C5oPmoo88NiT/lsU9MhqCquMSb/6UC4th3TC4ABGSVwyjO1K8y93LKE2rXUeh+wQ
C3WVoS7rcwqoDNWptIYzsdUvzhiNudJryBt20H53rMAYJ3E1w0RWRY6earTKXlzS
XBkoYs/nPjjBpt9oG6joPzicFQg+6nGyHbmiIi5u6ELyfw3Nw65BcMAElzyRCzYK
Qjnl664+Mlzxn9SPKvXPLvjxjGLv4xd4RSPTdCJxuLICxn3iupUL2n8fNiS7c5Qy
Q0uirALwSqnU0B4wa5+Xw2iCOaeyPlFyk2xwPA4liPfAdb+/TTdkS+oHxdCrb8vx
YLA5RLG5lozfO9fsbnD3p2bxWeXRKmVRmH0M4NJRYF9vvkWNEblX9KzojVkZxBRC
xrMLHwlw/trbjkECNrsDXQMdFSha3q97T+2leUBOyKNNe2UhbPetNUvdrE4hptCD
hj0HNA/9bszdQac+qca1X13qJvp+4SKSbVuz79UYF4SkvtQN/o0LjlVUBi70qXtR
gbSYOQ87d6CJ6ekxuCDi0jLur6s7yHIGtHpvL0UHCeuP5xVGqAKqpoD7N/ue87+Z
96jhxYC4kjr6hTmyA05nD5FFCqrczuwfNVZP60Y61ePCjC/AUeXlI2JqlDxbjgwq
G8BsV2m8lQk4STKuz4IA3SnlX9cOBL4cfh20zajxyLZpXOfq67Sa6MhckwVdJpRD
C8LLih+u5ZmPFawZpa4GmHDm+tGR2ftgtfAoStZGsBDFupN808d3g06vZJxA6tvW
7hxHVl5kPnc33Q7ICH8ZA42qtcaD+XwhWYDKvj4vbGxsZWIzW61RiZ8Uytbw5Cjx
Dy8IIPZFJVMx5dK4y3gL3bkt6+3oO2LV/hkhvzzmYkxi8DACU7VykyWlXAPBEj5x
XBpSu03HLAr/u/2AkeUr5yjSdr5NxTAhxk2v5w6EBIsyL1RltZOQcLtFEoQIa4Fu
Z6PHqJLPFX9rBvY01Syl1DjmVurRg6KzLpAaeVdTy1rQvY4xL3HNNr8n8/V9FX0u
ezt+7gBqtfp26rbxxwMItg==
`protect END_PROTECTED
