`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CMX+P7olNn5c0JEQKtRgb0CDru2qHmaXPey44THVOykStFqAvwQg/7Gkaqfweelp
9TR7JEJ6RugqjVeZ8DQ3MMwdFi0Q+74kp1HkVqRcWZN98fcqh+LSWWWU8vbov1Ja
+krVtz9KwQmrLRShLY8Ku6OTjFkZWG9qyOGlFcc0hptXnhXL2ZB+29avfxMCU3YA
1mUy7WGuwGEw0EUDDz2a6jP2VHNWPI6CVs+c1N5N0HHdMrMcFSl7B8QhnsFonuA5
fKEy9DpfG14SKUBIDNJAWeaDhqfvnUzR10PzaNTOcyfMS1tdOg6Rw9L7kX2mznn0
6GM6lGCQ1EARExCnX5OXLPA1ahkCs6UsxzPQEOss7lD3LqK+JYVNEIHHPuTY+Ok6
`protect END_PROTECTED
