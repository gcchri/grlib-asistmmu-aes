`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wdqCrADkpxU6mBOdAZxUG3Get5IHDhhB7+i7r9LMHiymTmiAphBUJIw3cIg+a/OJ
T68HC1GXWROYLLxm9Ce5x3Gn+ND58zT96CkAPNp3o+iUKYvDDA39iE044SJC/FIX
XhvWIqPauENNB2bhy7OkTTkUvV9euncel1D6tT9mTtEyIPhbhpYVieEV7FD7iCF8
keJC/DF/38wgZVGtg8YEtnJs6DaepzULelfjIxews/LZWdoJhy8BjXEIxsyBbkYV
2mKropCm89ymIHLa9U7+7iIucI4VolsUZ4oO/F3lKE8O2ZwbTyC0fcyOG9VYQc/w
r4k9Kbnd6cASjZJSRIh3KHpWivvVHwREWvXYEqtdBSsai1GO+aYi3vo8sWnP3H+T
Uk3FAI1ks/0y3bSp9eo/b9pWO/CkGL6axso+Ie99sLdUL8PNcpTcGzKYxmQDn5OM
o2w4N1ICGPH2JPoNzDZm5NBD2wOuyq3D3GhIma03EmW4NkXbyk7hIinsOSarscss
w+Kk2UUYXy1dMdJaOT+tKhUImNrU5iTk0oSpQGpFfL2rmdbB6vtGDkgHxwrUJnKy
bhxPUPWFsNTXGkeSGcoFrUpfpRkz9tteBtNKLX0dlyFZqLHTaHzO0RI3D1P9YqVz
7qtwtonnayvdv+WuPDAzgOoKuTB1QqA8RgGccxB4FFvsxrMd6FVW8mrSjwUGnOhi
eI1P2HIhRgTxVSKKKBeQWpmtu610ELmmuwDkYRNrtJI=
`protect END_PROTECTED
