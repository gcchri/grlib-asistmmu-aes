`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RT30rx2/zgtLdHgCYzmZaQF47MmALt/3ty7DxNNN15kEGe4diMM1veOT/Ejdxjgi
TOkvCTKr3B+i6I9Lb8XYCXRl5WM3ps86KHPf82Jlg02GN5Z+nX2KHkGkQtd5xUN/
41QIWQidXIIF2n5NYURlIj7COtMNxCy3WNOheDFaU0R3ByLKD9K6X8TPxreYwgLq
y3IVwekytVJskchWLO0gyHaXSK/4QaUZc2IWtnS9jXtdWbzmSP9zLFqTVFnOv0O1
vhXpOSXkwGz6+Feje8/0vNng70kGcHsMh6+zqTl3LlQ/ftLAFCOu2TVw4L8LCsP/
f7D5I4BcTITmsoLyfMYlIGeIhLC5oTtHLKE1ojwcmXdDTvi4/r2ZU1pgyQMXUA4J
adWJWtiSCWeqp2xQdYKawN37F9r/J6nk8/VUt7OPooODldcJ+TAiOhjnsim1XUFT
+1dC8W4RyzH3lo/L1TwSxixH6aQC8yc12u9ZFLtA8spnNKxKe83DxKpQsJ1V4IS4
Kp24ebVkcB7pV1dvqVqcKzM2qpz4/QNjFTKApEHz13V0J7mb8MKW8esLCBK/2atH
4UNrOcw+Q+qwvhdNsGU1BNUE2TEQdqFGnuAuGQO/5njHUtDfuZCvSRMso/BujcRr
YaTFGuqlk9iGE5bkvUPxf5Q7L0RJEf7CbaO44z5rsyExp99eQGwGvvKBqfurgj6O
lNvu26lo6EbuzjG6A6EIQtXSGPR/oFBMPlnTh9L6NGj45tnABKcOXBwDZZ43Di+z
BgVDtWTlK8qzSlAmQ7NNhLwF9/XcOZZD8m903eNOBN7cL7pBWAC+gjz7KwpeoBSy
JIQGJAQuDI98yosi+0OV7KhudQxDaOMIC7FHQq1ifFVSNKwydAIbY1zCfC4bQxLK
UGoTWfVnkDx+2O6PaeqhQai0kTitAMc9FeU+gg2ZkuA3IOUPMo1aelRI95f0VCYJ
4oA/zuReBKJaNr4e+m0mKb9PsWZmb8wdKTirz2OaDyUZr0ImPzQfvlgUGNK/paFI
xYdmXUVLwNNPnfD/CHMPE9dhDNnqPne5aVWYERm6f1QBZSN5osdj01/wVFXswZd9
Od0e9qhl+7qy5SGrKy82C7dxlQjPDBt8LMfvpknmB0CIL28XDD2OFTqVwhf9TbCO
b67u3lX4+XW5STa5CBnGIoIzzja9ncEuirY5bk6dDauEe7T6kDECXUplhKKsZ0zB
wSIjripyEplRfz67mZo7k3y8CtOGHrR4AA7tP3SaU+eBAjdM4sU4DuLiv6WRSc+3
0OD9NF9NA9egacB5JezFGxbuSTlkHrwYd5WPe3SVdEBIVBeRmj3vCBwL4Y74O2+8
RhGB7fhjgEzgQGpOss3nyMQSWeupluvDRQARHyFppOUZSpU96Klv01RhjrbxSoW1
967aOotER/+/yvUZvbbX/bEcLqC4DiT0YdNAyeRvHphg+DTfUF5zpyq9+db4Qdw7
kkPlf2noiLi8X5PgjeyBLilk3MrDU8a77kxav5MzGGaMUsY44cY+/S4sXJu0rvcu
CJluVioWpszdX37sIlbP3W5fCvahlM6E/rJG853Ezi0MEbFIK+Q2WpcvTtVmrJVG
BD1YE2iRKue4fWarzLzM+sxHMO8SuuG0UtkTZH4L6OD9/kpfNY68KE/T8qzZeYZJ
yZbF4wrPEZoMraG8nxYT6L8hu2thh3KLRUH0npkgjmrfpm+UzR0Bpkncfabd0EXr
ynQlxb9R3NuCEIenlMeSYOqa4abzhMKdnhjZt2khm50=
`protect END_PROTECTED
