`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Ghso8meGiiPs3ui+dCS38QB2m8Ym2xxRonLCHAm/4Ya8aidCwFnX3NwdVEsG7NZ
lyT+DQrce02juWv1FH8WixCqbEEfMqUvwyN08TuN32g0sfUezuE5a50yExNHP2TS
rhx5I231K9ni17XdYBW+dm0r70wLl0FyaRY0lJHyzDKiYdzOeRSBl20wa6cV9PYt
wbvyGpYbGvmQO5BDFVODJVrXeOhHcnTQC4utyTzSSDb6HMVTK92fsf2B3QmjaBIS
+Lo4YdvW4oLuVFCYONe5o81Q2wSOyVafp2j2BsTIcdg=
`protect END_PROTECTED
