`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZkMg3pV+fhpNkkfBtoLuanrdRyYrlQUpWDNmYFN27Eb45mD7dYYrpmmEcJi93qrG
kWbUBKm1xIvZzRlGhKteNJ/KGNI5bNqhBXbAbw2S63gUMnEOY3ikW1aYoGiiDlc7
jUgcx1bFK94ooPfCAIqLncV13S7vWh+GtBiws5Qr5k+O1334VZODdNfK25XxLib5
QlnfRj3uiJ9fGzC3LR9PRyfE3eGI2LeJUwvGmtBIBHluc6mlpPZJ4f4n3AZOz2Rs
qgsyQxiT/hgiudJHlYmKeQiTw6adrsbypJPs01r08KTsJMK/zvoAiTNDP6pUASUG
X5ohfx3D5zULYtjQmMhRNMj3lCR+LdhLSCDU5PivhqohMOGmizAMOwER1bjWRhHi
qo5iDCyV5TDzuxRWWfv4sFFo3H9RWWS9dHU/Xrr7o0jsqzCXm4nDLG1JpIsujEcH
o7c4qr5PyV2Jzrq+czJN74R4ce066lS0uwT6X5yAdPEF6SwD7dyDoDXZQxOa80hA
2BOwAxgxhHFiO0W5j2K6GIS2X6iz35cZZF8xk1L4EkvL2dp0yWRrqayss60VEKmF
kz4v/hjD/1ZXg9+a28TgKtOOabbO/5VFoQQlu6zRhr0YqiBEfRTFNpMnWv1Kf7Ot
SRWqeOvOKAmDjx4EwHyjpZ1OST9XXze9a4jM+NiAf6Z6d3QqTRtzI3nmg4NCnBO1
+k08xzbqUZA2pVrZ/BcsyQwBWxsZQ+baTwaKnE7Enwis045xTDXFXJaGmpulxC77
PBkWdaP8g9i0PnkrTuceuN7+P83MXnC4bzY8MV2ZLXI0jPNBtX5656uaxrdxvJ1P
smFKZFfFiGdeRXnW4gYz4soCcJy28z+UDRNTLYx7kjfJ+hkzV/Esz2beF8O2dbFy
3LYnA64p+5Lyb/De1CmtB/f91/wLWsMPUCiW9/x8J6A=
`protect END_PROTECTED
