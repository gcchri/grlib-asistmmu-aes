`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fYmGsZYoFll9608/m42J81fr4BmBDYp2lmy1P0AbTVSioj5mkRJTE77i860LLy51
CVFL487k+8ACBp2m9SHytDG1q6DmsQvclV9yrPQiKXj+hSSwuyRj9VhlSeWAR1Xb
lafAFHM3LfzdCjRn9AT4xkR3nW0WEEVBPIo9wdThqU7mQwlMuemA731Tx9GLbVBM
04lh5ZO8XgM5D8UelD2Bvg==
`protect END_PROTECTED
