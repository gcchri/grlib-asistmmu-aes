`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EUxovpOuS1+jRkuRodaiANvPvCjVzB7MYNQ5HSJfmw8gryPDVusVqwq+PgP+KoPo
k3i53j9OZFEOqCEG+Iq+3Z4P3q1RZrJrfzz0T+becc8J2/jeYTHdtPrsP5GJ4qCS
hrflCOwRdWL5FN5hkaXh5SdwL/1skkyH8SKJpB1nuDrhpG9Rwyabu259WYgZbdWd
e1F8miVZ96ViUARVR1b884isop1ZNnucaKtMuiOJ24VithsFXbHI4IZcnxjgyDyz
s/5SXazQia7cM4gp5+h2AuZ1KTAvcdZFlL1GMndbYqOYla7ittEhTmvnl8Sa6yLV
UAtfFBkQuyawC+7lFk3LYxFmu2hl4MFG/v0mJV0N3F9cVutX7owFsCeKzegdTQ6Z
4NJqNyQA2bMRMI0NpGZ6arhtT1Ff1rKkB2uVhhEoDCnGKYX3VYXKZKt9uYsbS5mC
gY3yJcEUJuf8fn2PjLD6WO3Xwr71pxsBnl7VqQ4wLiARCEFT5QDkKgn2TwVOitvq
5rHsyZGjmQ3WQwhQ75rUjklKFSjY3h44JJhJUZdGXSQOhg0YWMS10yr0aomM5oKV
uXTJsiFTizTWdJ/qeKLrUVOfAsQ1m12+aCvUgmswgYrDeWFi/+TCfuFq/0qx0s32
/sD3gRVqSogRxlLBAtcHjDXVFu03aNTiX2094sHd6iE6Ri/xPiw+a/cmqVviurGV
rmEyxYhB3drA6uBnQ0SBiEM8drEHNwN1iczuA/e+lwgIHSVzf9/CgTaKKKzkE59P
OUlt8S6ZMLOooVrz2/qETQWS44fycan9pBvKSdkG+kiqxAoCITwOZ3aRrf5dHJCk
4bVYUN5qsIF/1D9RBbgdOsT8WYv8nDeGWkF6wN1ViUaXrH9F8HpL50wni/mG9QXw
4y8bWNmXxVCtGtCWYw9UQw==
`protect END_PROTECTED
