`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZIDw2dPLpeOJZOQpzC8wOsftHwzcNHsEFXH3iazotuAWR37pmQkni2YmRhn2uFmK
/iita7Y/6uu3Ti2sS0ogDHbvfiNoeJui/wZnMR14xiCoJeU6VjdQYQqPkJ6tVvFA
rHObafBNZoRGlFBanBHcstkFVGeJUEkVQaf45vCKsd+P6uc3J7wnyhIW0IEMWYs8
LPTiaacGdC1sONu6RCVOGUL+JQLCkvd1tvkgjf9mqgSnX7qyc8+MnOxDgeABerR0
QSSOH1VaGoLyT3oeYizaKCHM+OHLXDcvMm5qzMRHq1tvijcvoAgyQyi40yE1RpMu
eMz08xOmNsavSGWviq8vGTJXRyx9q2ZFJb7GINDnXO0GwfCNImHwij/0/0VWFXSM
GtLpRyx12+1guvFiWg0CCxPsfBUVobRk4Lxb5gzowaFznA1cnqGQqb6SwyAj8jT2
1luG+PpXmr9LwZdZY2cnqtfyg91iPV2Q0ugASYpSmzcn4HFLSyvL0qb+pTy1ZufE
UiZeun3N7ThzQnxsrVBuB2s58TiANUZ5+DNl3+gRuD78BFP2VS7V5loSyBrbiPJ/
3fiQmUoFneNfSgb0mVk3nO4XDCer9LUfZ7EnAhHjBBXnexBxQapgT3XMhjmhs+zk
CzYUa0GILh57rJZ+OUKvkCrlO86uuj38gDY8twe0svRWmp4uBHHDmaIDAE6/QNGT
b9/EvlAKGze5ut1tpIi4JIWsWqZnfL8v4kPwgU3pc4eF7LT4viVQl6Rd5YLSLBcO
eMLccWLN2J686ko/dpSKKapUvtD4tLYNYOYdZTKOhiLRyQKFI/RnzII1UD9mDAL2
yG01MML0QG34wo79U2g2vHAGeJiSvUy1F4mtVbPn2lq3+b+ZuHnvazPbxeyHWMZM
qFO6ZK+Voqg3Nu4gIEecfz40l2swwpL4OuQMKr6NsckrIOF0TnAKMXpYASTeqhKk
`protect END_PROTECTED
