`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GWqulEGE+KrmwlM14RGki3bSQAZDr+671frBpg6Hp/htsueWGFMpBp1ML7UcF83z
DDbhEe1VLxA4N7nnumceHwSfWxagOhFX4GlVO1VzihkVr/vAd6fwyLIDGunrGoum
+IGx+cPgT0eFOfMNIp+LB/TnjQkuD1YYYwDzHX7D7odT2ZDxL7a0CLDQtspH4VvY
mVPee564esbMPknOJJumTAY/UFezza7nWaegO1dJUGpHBX7iYIttW/QSgx2Y8slD
1HDmhCm844+BrYfVDXmscMqvt6zfSyQU87dAE3DQP/Y/7xpRowrkaZXhjzMRDCEA
WUjP8qWKZu4S00sRBFYm4soqAOSg7+fq+MTqsQfNIYf3cKMNtMG1EMRuur5wNScE
Ihd/vyhCcp1oaWg/upgXeKu8FcQavIuGSQ78jv0VUmUtM5ZKpoOMKfnmYRPH/0G6
F8tKOVOwWOgbo/LSO8Hn7oHv+3hw3dAZdmHrU59HQdMHZbM6EHViz7SlPytEIU16
UpC04sPpwjMStFG6iyiRYBa0auMX6fvowqmC+DNbdEmq8cUp680oZbvY44BLIDD0
HOLrm9nRebzhLKO3l7zpiA==
`protect END_PROTECTED
