`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xVMMCd/3hFh2fOhofV9hTWdGfdmegHK1+0ukecbNZzJxD/MOxODIYQ5qEOtjkN4M
HB6GZ+pvAuFzy+WzOR4j0bT/IsVyakLis+B2rjtySbL1fYvdJSZl68wbuskc4t9x
X6lMSqwnVNxPzpyZT2dJt4KQiLq4e2WZ1zyXosIb9bcIB0fkreTnOh0Vslsighbi
3DBV2LYaFa0EZQcdSC/w9j7dOCN6w1Rfcca7cjgRb0adgLhchxT+pxoFWKq/CHps
aF9PshqzPSKu8TRLSZfctgPUQZDe2ki84R/yrIgOpZPBrRLvCOVUm6A9nI74Orqo
JcoY6Egh8OCuzoyHTDftRHB3vNxj/0KFiFmIvnCIMf5w06dbPBNgXXMVwEV5NNsO
22lvTYWC9jaYFgTGkzWnFxxzBdj4ByHSILC9IGNLh2vad9BGzjb+iDswX58vbwXq
NzQCwcelS1rWVpnOzxJOHaQ71qTvC09YIaRBAyc5nJ/fGdsQS8fzr9mANhf6njkc
`protect END_PROTECTED
