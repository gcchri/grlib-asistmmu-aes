`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HHlvWoO0RIf3yBbLWIxPqQK5aKQUEV8wBt0AlsqphZnamqkahx5bOymV6IQ5UFeX
p7PVMYnl3uox0dDblqaEADp0pmZL3HLb2BhQ2za3Jp6rGd4vtFFOKgocwXKLu0iP
mbgSP2Sq+b3vSaYdC2fdTzxBtNVWo4s0MZPNpiSVs9VxjuGqd38kcbop8a2LmTHt
eVSQbdTwu9nzlJeo/bUXxv4nVIs3mCYzkjlDGdq6kj0Bp0QQjUO7DVSsWFq/Zy5J
1wAvDvv3w4Rqs+npQktftXoyDd8C1U/6f/0PdaoKaEfScUs92Elkw429/WayVqzk
1F2dTw+2SzBmclO9DqUbcA0v/qysRyUcyL996HkQueN5c/as+MfrKWUP4KvwjAeJ
nCfnCEJpCCdVgrxeHzRjFrLy2iCfiNRV2R1u9GFsUnS+0xmMkR1xpqkbcyZpX39O
6DqcDYt8B4ZsAVfzlL4CXo0BKHcE6nuA9CcdB0Iq9v/KAcNG2ltUQ36M4gLcLhN1
aDqHmS/Fj3CWyUknPFR8bX5hoY1GTt5Qipd4eIzvwLVRNtlcD4a3cRnR15pHU8MC
f3Lg3DTKW/JH9MIYDGgAPTULXALRNVjZZrehzx0msBWYqYfzDcsaupL8fzohDf6Q
gqbLYGELzvb9uhh6Fo8t1DpOhx/dTrAQRS1bJx7rlxKyi8CLVyFc34SisKw5tLIp
`protect END_PROTECTED
