`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
do0Xjv4Qw7CwTyaAhzMde5lcGEVBwZ2mjumNJoIETT2nKXMf8MNn3tmd5ocbGUbe
oibJgvUWGpkY6Yyk0VA6cXDLrFLsHa7hP3+EhD5XzdWZfq6F07yGBb8vHwu9NV3B
1MBmSnmyT9Ql64rSZLhldC1ODNh4XAi5ujNnSmlb1QE54Kg/rGHia9SUyPrD89Kg
LfXsQlX80eqtDntSgpT5PeiJhv8MTlfrBjgKb7h7O/Ht4TZCEWfZrMd02T9DCoAu
cnhncz0pgo4aUaEc0G6sw1ftcj/fUlyAeWeuz2IU+AmwTzIxpxZgEN6ScezZHxp1
7cudXjlQ1EwZjzPjhmeNrpvSE+xPajQ/zQGdD1rYzFaJSH/mtH3u0ErlvINwqjlS
p7uhxX3FLL/3SRlmqMszNNRLdhEPsBRzh6+uXa4kBCWU/e1z/Qe/1GJ+mmylvs1g
eXTLuRhgPQWLaLmfqUiHgkg+wq9CA49CjwnAPwiAl2AGI6Mf7k5fVD4LAr9MXlUH
Vr763TQ+19Fl7RxS4iIPoK0HVMcyeezQupiB1EIx5lE160c8bNAU1yd7Zw0xTIRx
aJA+OdffTOJPBBX+PTb5q29TxGlF1K0+5M+A0fj3ewsMdWldmZmA4aiHxIGYLF6i
w7HiVQF45Vdya81Te+EEf4By0CGqk4gZt++yG9wCG8fk+CmawryNH3WduqMcL2g6
+R4/PF7RwXML6SirX9Udtix3wBtVbym8XqC6LdGZuz+aefJaYSAWByT5OPoWZWVd
QfM5M9nD/T+1lpjllBGX/6he7w872+Klw/hlQ6RCruPVvcobASyP+m4VuqNmbdJ4
WMKLYiunCHOuOjVwAgtLGyVoV5wQoKahKbGU9h4VuPYtltLvQ+Q115qXkIs+graT
ZFwAD8UJsgOiOGVxHiYMdwl4XKnuGJDeupfRE1LQYjDP7OEp+P2caeet8Og6W3qu
9/ydJ1NJKQb72tm90mJCCT0yrRRYD6H7UCK15KcCuQpQdir+yH5dJ+vKXHyyV+Nw
bz/9BYTRDS04gxTh8oe0+v39cCMUgW8bK4d9gO9XoXH1WyE87b514dJBzw17Mk4G
H7vXd8fnl/1lThTdafL1UEzlA9vy8UmCfZczvHVyoBuC+T2vvCDBKpDPYMhzZCFj
0GFYXLevHail1ItDmMHGzRee6u/x6bOYdBNVa4Q2PzIf97yphuWhyTb0cZuvva8k
nPIDLJcxyOyopHXgcNvkcJXTYVikXVZoImJ58Y8H1C0HVXUlrtp4fqdFm67XQVfi
Ctc+38KWaJdWg/M381aZ+meCe62FhPGpYiZia+1MDExUg3jzBATpTsceKe/L0zaM
t8mwq2nVZXPBi/VuKWNZ+dHq93ZRmj0bS9lrq0rpL8mf2yFYeXhLHbuY9Zzu2LOk
zNeQp0IbAA8LrBL0VX0fcKmugnwMD/hXWzb2qd/9yKTQFb5niOvKPDZZdH1TFk8f
9Swxm1PBa0AnHnqya2uUD2LfY1QOzekYYQR7kwJ4i40=
`protect END_PROTECTED
