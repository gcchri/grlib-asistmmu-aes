`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mUO8M+nRPdEWbJPAnVjrzrHmxisqosXgp+lp2GNKjBoXWSPJP+PNLKXoxDmilqiA
YLPM7eEwerqDj6Me1yztPi5cz73hTT+IRtcztNmUDSfEJWR35sIIgB6+zbvMKhRj
YlD1qHAahiqaUwsrR87eXIXYI8LeUSn2IeBkSHySvzvyly/QNHm5KKsKkbrBtp+c
r3Az6pmHbxo9WTZjpCymDha6FUy8a5JGtD+PcFXnhM15FwcjXARefSlLXgQqlpnO
c37GCzb51UE7mlfrMCwcedLTJd2wcr3/sDsO8AcYEA16Gg6X4wIjJhd78Yy4roWX
eWksdH7AkiMUS/YvS/6UMGrPImADX1HJimHZanbEj2Q=
`protect END_PROTECTED
