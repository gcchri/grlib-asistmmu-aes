`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XucDm9nl+c7jBNCdAvRueIkXHMXz2wKk0HxnXHy/jEzBU4WZg8ZCUl9CQtLSiN8i
Nv8rQ590qLXp5CL1+ROpibPqlyKIEfxUd36Fzc5xpvCIwtlp/okZiA1ToJvlXNRY
Uc/RRAFq7btoeV8VThKNQymPx3I3YQisOiHJfc6Hw66IdJqcZj+IeKZzA6EI2n3t
VnNTSl6OEjTeu2TlUtnfCistTqJpiyWTnqvGDT4Z/TxR4I4HKN3wRDxgLmDCPCvz
w+SGKhryVr2gONuJCP0zI6Wx5B2i6X9zXC2JlgZSx2ZlfoS8dv6UhTd1XC+y7UQU
wwqredZ3SXduIBCcHLWkphr4xsB9xS5OPtTrbBkrx4dY/oP31TaValXIvshbcyGn
+Mg95AWF5HFnU02qW0rrU8rtOTOOGdls0bSVTRBqIBsf1eaIK5usXY+l1ogCpbI2
`protect END_PROTECTED
