`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YVM7l/5Ka54UB6ZvuS5oy2JyU+78NlLJwgN6sbRi04eEU/nHvU5qp3fKanHlIZov
e10Q6zFLjjapNWrUiX/Lx8zAMfLKDy2dRJu8MSUYE46k9Gj5+hLA46C1ONFrYoPc
IeOpUjFzvdp8VujpdOrpN0dmz6tvUUQvq/Jd9s3/JqHrAHO0ObapBgViUy1pjVXR
zgxI1pE5SFyF73Raomw5U56aj8DcZhAg4JkUqnnaCU4cyMcxsaGc4olKvsLL6aeX
51dS0cP6DiiYos4vESNZ961w4c0cZ+jd7bIQJXiLPFXQki6QL+sgd29tNPE56zEr
6CcC0fLNDmrXaBwmDB/8zJoPgygNEKwa96Kga98ljkq0h0sTxtNClcjWMn3kIq8y
+Vc+PSb53kHtyWfNWuk6RGUC+P59TUGE3SV8+FRx55sTx4/i1vYKbUyme6sOxvMe
5QfF5TQYARxl9cOXS7NtocSKFD83mATolM58JEzAUrm963ukowZQmVxBfBz09swJ
tw6HnfyBjS3oVF6IRInbG5cVLe6ZkyN0G4juDzeTkkTzW35e7CNyiNhuywzHT2ns
uGk1iFk6PWvqsCvSTOrC5XvIxnjzyhdK8L/FKpc8tp1f3OT6m1Dtd//zC58ZxizQ
EpNkZmTfzP9xxUazUmnIQuoJ5cbJuoGXYWVtUeJTeok=
`protect END_PROTECTED
