`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Y1Dj0jcsWiosvD0s6w2PAT5oV7vunjqupwKHqRhwPXLk4HREQmkUBWfHwmrInWk
fdPFxegr1cKjs7XQKdl2xOLbwdgNi8S6RJb+LqFm6t798C5MoiM48g76uFRzdVbk
wbyLQW7U76T4/6nbNbWJCCvnMPvt0lRLuWPITg6XAJcEvQCZFp5z1cbVWJFeJgBz
KonnixHcTlIRBlpxQy2suLaxmWf7pOyJ+1n8jvWfoq8heknBvtB4sCa7wPbo2OMi
e2eEFPmmN2Eeiamep5mYxHnOwVWGLRIFbHLCrFs1Mav3VDyDuvvHqkSFeIk5DWKI
0pL3fAkzqB7SuLIHifI0TzcVczI9EUO55ln2520XD5+xAIvvrZ2MYqIbu3CyosP8
Wdhq2+Ax/hvTnrigXiIGs1Ya0gam1/dgxs2ehY8OhIYFWfnktq7Nmdhn9wJJeBVn
2/ppJCN+b/qblGFrq30qB5SXNNMsDplI9Byi/QIFWzeAvwuC8DhL3//1+Fj8jg2a
sYZjveqsKF1qNLc0fJwo/JDV90hwi4HOqo+bxmc/Jj12ILCWxLKz3RYnbN4e0Kv7
UmN7S8a3Sa75Pfyels8vyOU0a3C9obCUMWO2Mo5Ghq478vhuf//LCWPzUTl50X6v
IDtF/nE/1hA4ON5X3e83U1SH4OVlFgD0gFBjFQujpqNVNog/Bs6BIINBpboY1KjI
S3s1CrzaGa/1EZ7/MAAmG3VF7mim/SY8qvWDS1Hmx7VWQzk2GUUU/Q5/RCnbhFTl
4aihiLbpvF+amZI0qkJOVviMgD3RKnE7hHo8GlGGJQhBg0QGiK/I8zE3iD3obpcR
izshy355yBUmqdXvS/gQhx/kDYeL/vQs3oVLiUuO5ce8vZLObKLy8RVj1FV3dYpm
T+ufr651TUhx2zk/vpg/PsHx7NKkQ4FiZV4gdjru/Lgcywp5KfTwa7tPGiYdAW49
1j1TD+lkHrzxR0blxm3ky1Yc3Zs6QPc7ELEcshvDZduq7JpLNP++QcyB0XEURrIb
EDFi1F7uP7LX7cppcWLHUGFIjJ4KhjkD593OlxdFyGBEjvL5r0KsThXUIWxRwyMm
+7Y/OI3dF2QhZtegSHls70l9fnBH+i/zXn5KRPulxv7D+RvS8j8WC1CotgHnIC+4
tdDZbzAhkkkxIK68VicH90KqsNQPJt9Y2NQdU3bFShWwmkgZEfcDmGAmCQWbCrOA
mMwf8WfsTYMwatZ/JXQeHiyB2Sp6ad/AjB/T6nLyybsiCe38okoAL1mZJgb+glks
`protect END_PROTECTED
