`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kiYzsNwRb6JIjVS0sdxxrqJUlF62oBYImKGfLWLV/zArk9h9ZRpSItWDMl52HyOJ
YGIxW9eZUyEuyUNmTNTP3TGdCMR8xWMYRiCdNPxfsPz4OgyXGhIoj80E52WlbyXG
/jVT83ELyBP47E3Usm2oMn03AgIdwybRU4ONI0Xo0O7F+wU3QOF6s67YU+2SwgkG
IpvR55gAbFX2Qa400vFZKx8HhMejTwpPAYGds1g9aniHChwg6U/uf8DQSGLAB0JE
aQ5HItTHQq1031wGNFefdAcSCUz8KjlTYMoHiqnQl5S6DKNnyKpii+aSh9E7wLdr
UzHD+bh+JgWPBQBWlVh8UdQrQ21gPOKLJ0EwCu510uhhwqh6CXDxPStIv//s7uhw
L+CSP9nqXfOBGtXRl+C4PTAvkJGGB1EPOseECovaKSGtyZ7B0AHsF+xpo6Rp/T8Y
Ts/S5/Jrc0zQ8wrqnEvQUVpqAxk9Z7nWtvCKijSJwwQu9X3cdmUnisE2V/Nx2izf
VAPbgiYhyiDGQwVAgM6srZfInYJper0+G6L5V56YAL/MyC4X46Aar7dIjcS/lZmS
`protect END_PROTECTED
