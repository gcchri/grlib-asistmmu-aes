`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+pkAE1ic728lzfwT9enuuYWFUiXGVLiiouC/L5mmeRZhKbS55fiRSIRjWl2b22Ql
HWReIbnpZfzB0DcunapyugB4j4fuAFKs9FjeuUs+QYxkPtGdZl1ixLYb/1Hi/jk9
7fChDr9KfVOTOi7Y62+jXfcdPPNn65ol9JjI/unckQBd9tRhaehyhA5Z1aslhyvY
a4Um/FzWdsMzmdIjm+xJenbyi6N49KpwkLB7lQPgns3ylyw9mMl/WWnLVdCtAIFm
wt4WZGVysD6xSFRmiUlHX0H0uejRLpjjzAIvmfWLXnLpbKjNRubSA+S4tssJHyIX
QtTUd8ufrOscEVnyNZIV964G6OCMwSr8VIJ9F+U+kmTHt3N/gnfC15axXnRJdk3b
JA578SBw/6yve/PC3PrHCO0FC3CDh14EICKj1ajfVhuxz/QSOflDHHm2mzApqKsJ
XB4hLgVL29vCMHeneEj7mPQl5rqJbea3dRmB1/VOy6CwUAf6bxlKyfL5pgW9FYZ0
qFnqrz5Ef4oNMItr+WXKiKWfEzztqHP46p2wXhNc9L168M8+x+rQk9NEXv//KDYx
O8ilB44oDfI+sV9b0okXMQiJMFZUm0tk5VwPVqcszEE=
`protect END_PROTECTED
