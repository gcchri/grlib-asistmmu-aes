`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
//rBdvPc0jXzQYuUrpNgY1q9fZ7NIY5rwkA3om0aJxgY2ubIb4n+r4Ol4kqyKFv4
iCSfUqg6xzYDlWmcPn7FCDXEEXIyTpFi9hBQrfErL44hh1X+NcE8Q9/OvWo5bM7i
8pHHncBt6hxqm3S/OEEpnr6Z4jLVg7/UdeQcPZ9UhDzuASUrfKXn1io/C/rj1Yan
vlfaqPHNtZaD1ggN+B+C/+2of0vX+ZpWMKp7PI31IQvmtQtS7QPLWb33MN7IYeez
p54cimlDlhCtsskci7tsXS6ORtwl9HnUrLCTsFiZV1qaUlWjQVZpHAIKpPrfhQPU
piXopR+HDOzcIh79kfqYrZM9HzASlE+76z83Yt6iCkgWCzBxUl4Me9BIw8JhsMis
lR9Ri4IF6Nfi3hELVKX9sA==
`protect END_PROTECTED
