`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FnM2qWUcEmNFKmtzGdHDZ6D/A90ycWu1qWl3ZdrM10ASEH0airUP5GWphLKlrUyb
2qhqyWe4i8hJvBt5TuHLRJyPx/H19l4uJ8aEaFHDYVQ2CDxbUC4J45Bm8OoH2dGV
uiZn/d/QI9gIaTyUpayyPCl1oNyL4zkJTfe+JTjp8aELmfIR31xfho7dKbsNer+9
hrd+ZoYPeOlyUxjUQ59W0ZU1Grj2XupHx4bh4eTZm6F599cywOWUqZQkwQuESqxs
xWKRUZF0jXiDFbuvHVS3muMkGBwgq9gpDB70l6CdPoEGTiS8473JiyeiRwO9Oy9+
BTGSTLW6NGfFxW9ogxFGknxiWUY+Mm75iKZVruexkL3MgzRcq6z9EhHCtXYTeQVC
`protect END_PROTECTED
