`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ggnKOlE7cdiPYuJEO4LhGhNKuMMrOfYavRk1QuSYo8G9fKIl6LGWRgfXevlL7diZ
KjyrAJbRrXzSfHjD96EtlXBA56iP8BYAHTFR7Umc4CcwNFmxhkKu/PXJmJ+DM8Xx
KaQUVN893+vIuRQAx4f9On6Zi8uLPRzaamNx227rWbRGTpUkLJd4RtX5eG5V4kTK
quaA+lia+a4iRg12WB5PfMB9lIq7fNTNiLJ62J2+DYMQAXcctScloB1CWlUTChuf
viSUmFKPN6W4Xdlv6vVdiFQwhONrrPOhWCuPIKPAO6t7F5XWHyzvpOZ7olElE93l
Xk+9SxqnBYn/zjnSx7ikoG6Sp7TJCqXTCFoWufoI8EnrZdRsl563x3+YAg1pI2Ni
wCvpkIgplqIL07XcF8PUzxwS4FOenH/rPMe40mCMcuyAPY1fMpmgHSYxSHJiIpHv
bLQmbEIJNrketq2wTt6mZz47T2oH+cmAN/+2vQmuWLCgpbNu7+SNbra6JPTcYR8p
zfINjQubIooWPO/o+nj+TfuYp7Gf3m/+igDCpWMEYTjUfoveskFyevnoi07bKrjU
HDFC41DdU6ESlxrRExiuJLSqvtyj8j+45gFQdGf15NJQ7GzAJ5Ofb8CMHUmxI2cu
ou7spY72XMPxVjndPHF58k92bEtTKLXUw5m1Fcs3Wzr1GbcfcAcWARBndVDNQFg+
Rq8czaLl1BAzb0/PbRptvTDOQ7R7fP7CfmGSnFztiUfoUZRi+rAOT6HqDbf1enDf
EcwempEwDXnqnR9+pkTvQ3mnc8zDrZH8j9zdtJHHTwnvy+rBkGTAShlJP5+Yv7Ve
EPfVjb5l2JDev9vImEK4d3U6WtvEmTrMW7yFTucjQQy0cp/WV6M1OhEv9cAlXFNC
h3DQFaSGY7z+r3gIhWDlfAAAmlXMkC0qKOQ+TG898N4XRYoTN6roBPnINh8lHBE6
r94uFlkq/PMzcvCXQuFMWrSuR9sB2iUQvSXe2k/R4p3EwAmq/Z7qguj6rHFrgL6Y
PuKLOcRy0/aF/kZ0aR6bhf8angCioPNi35cJTIfWhNjn3zz0TRzfh6EOVnpJiiak
H8lqYJ6Oer9Jz5wsRCZ7Nv+sIO9gfffrizc7dKxFclQnsxZXTmLT877ydn0+B9tN
7PWwoeI06e8iAauXrC+iGEuJZd+JrtHalKv5ZnHcDB2JbY1P0kFAZ9g5KNeeFoFd
LthcKCzmu/VlK5kBCpHZ9BA4yKW186Y1+Red8EumKAF+M0DbGycJgSXmxG1wQBSD
3cUfv1dTy9zexyDBFQcGl4iBJT1aX2oWEZ5OIYiSzRZwrSC3NclX8LjbMwAYCsTG
xgHUJ2vC664E6hc2pblfVh9lO9enreJDDG70TNsNbyzxTtl9fZ4a+xiXcZavd05+
nee5FitWmy3Js7knZoRaohzj5eX2ljrzRn8VdA4u1rPhC1X6Ilmxg5zqglJrDtWp
sIO5VDMfpHnyl5H94vL4ydvVqS5D6bSEGy6cpW5+2Vj19eL9ua0V5T2KIGesFwYb
10gvn0qgBEr/63wT3px6xYzNFn2h+Zs8ZrPBnYqCPGc9aAdX4uRxiDvxBEI1axr5
BUJYG7j81pyfe+pf5MSuLBqyJidlFBh6eJuXPEMrtfOJ1H0v7Aumvtb2nF2lL3nv
8kxqE3APZWr7ZkuaqIY6KCg5fsPaVrnGCrugwKS1Pvkj27+nTboZxCr9QsN8Acgd
d0KAIDNvrYtQPBvsjlVe+TR3Fj8viQt7UqZcsbVMNh513i714Rb7oXuBcRJSeANS
EmgCFFqbmUO/rqJJ0ryO+WgFq/m0BBgxJhLqzPJEfWHZmHcWUEDZNdWQJRZ8wZrU
uP3dAE6MSeoXyBwy3c7nYzKt3sjZSBcf9JtN4Jpx0HnAzXM5zQokdd9Ypu6NCvMI
zfnxfoJNtqXfErxDHlHDBwvBmmdBg6FRZxy75WWGrAk2S/GbSzPBHgHbrZFJJoVi
GhM7kUMWAD42iMGEr0nxXl7be8bFWGo8rVBG07x3ZqGB4qobjmty2YGNMt89JQkJ
PG21grnRGxwif71GMONKe6WTvANMcKc8bb9gQoH+L+zcCkvpWRUumH0A5u1Q/BXU
Jtdynd2+n7UEuVvYqqGpddCVEye3t5P4390uDYZ47qlvyg2m2+3pztykNjMwEDwp
5zLYL0LvVXciJWcIZVdgIkfV1Aq9utOIHnkQqDxJx9vAnMZ2s6i78MQ7boDVOZYv
kLwJKwGAPn4r3cTBd0oz/0QsOSLr97+JYfhuCbHPgkJez8GK+MPgEgyiDw7ScyFP
2/8qY8gWs6FzWhhZ8kp1fgImXXTGckRPrs4gbQ4g4641oXIOi70G/LK+DoGKW6OG
JxPqQTTMPpzsnJXBo23ECYlblxe2zoWTdo54PfGD4HP1xEzOQUfQ5hEFl7tYOsF+
dBS2TKh7nEBa+qkgAxFsqbTp6HwqsmrVYLh4QOTQwb2r6qaTpSTZpqBTf5Ue6dr0
VLYGosStVBOTBVkipeWbikgaysw/qGLhiUAi2DEoKDvnjKF05KkQHkqXe7Ppsbur
L4YUZ7KXOGCd65F5IREGHDEs7BU7HzhSPkOoJsjh0eY8Vyh8aP8DkUzpWXV5Vwo5
wStVz+4YVhTUVK+77zOi8oB2xwnzbO9BkH1kj+U8wLd0DcgPJx2htIt+k5wdqwKq
jUTL+ezcIrtiGuTx8qEFTkzRtWI7RAlKKIxagXMyZVF/ZkYef8I78ZyakfVTkXuE
KnQNZfckGhsGo3QIoGkz3Tf7I+dOwXt8OZT/Q+Wt+2GBkXT30aVA7AxK7Rrq/s8r
EQC46oq91dDEEQNM0Q/UDBnKqgnciZxJkqmVPOVepzWoPOLc8TltejZ5Yin0VJ0K
uhgLigATu2Xw0lpm98noWnzE+IYREi7c2zjlEE83pUqOiV3RoTNlEmhGASoe7D+I
qw23z+5e+csL/65M2TNIeLoENCSV/Wro28T+T5oM42ecfWBSIB2iKrOXAunAsqFQ
BqK+e9x1+l5oBT0ioK8m4lWP5RsEwXtETYKqRUAjf92tHM5ryn5JPVKqdfsz4kAv
9d1Ku5rHcEqPwZr2BuhRYWT8BVt/mF8O3rLBmR9HDnpXTa0Ng0vxyuP3o4jm4tZ2
VESNQM0OvaitinEK7OUKdhSHyOK5J0kB5bGSli+XdGE=
`protect END_PROTECTED
