`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+tLg9g3X/NQ7bu3MVPLui7Cdv+J4z1FMSrofib+y3B9hSZdFVj5kFCWgzVXB1Jrc
qFTXbkip5qF4j5P3f5kqhopp/mDbe7crA0haMoxwPCb2tvXzDaPKlpflQRAC0WMm
oJOZpUxrpMd2Q0yB7qDXvcszdv4tB7Uxora3v6jRCPUleklb0GfSdk9f+jcudjFS
gUwUNufh2TXYQOkwe2lOCQkxhefurKugoZ5KEXJV+MAu6LeBOQvLZc4ijjVlaqRk
wLaYYpY+mPEVtnz0jTLFr+XwTjbURODwSl809Wg4isnTNiPGHW6AQkIQX6ecZQQy
4zX2WasJhEGnhKfxg6HJuSgpKStvzYo7eJJrpH+62izitUdHKPYajPOQWdJx7OoL
it3gPj68lmPv8z9E0MtqmnHaXhtWvCYrtXbeTvONxKxa+zMeK9mhaAZgj4oCCi2/
q08l0SvIu6I6KFpucvKJJRimxdbdI+M0hfUt/MvQNCGcqreJVn62umDKR9m2MiYZ
WTmKO2Bw66WLXVKRPh9d8tAKSGzcMQfpbUI4ckB5ussG52nTK3Jab4FZOWBsLsba
Oh4I2Yf+RyWbBeTOi9VHLw==
`protect END_PROTECTED
