`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yg1ODZkptea3DUqoZZH/EEchoa175RRDxdLUhAGPxjFlnBHeuyMrvWkHvz+Pkjlv
FI0xUjZ1rYgRKgbBaq1JFBMf9aUgu/jB/iUA4OMN7LOM1r6q1+bvNSAA6iqHbmJn
UrI9c3HEbPQI1ulqG3q1+Rfiia0Vg+s6d6f9qOVyXlZFOLbqVS6yEW9PISZJSO8O
XpycMtsq4O2tquzGCg/YwLvqHjnSezrxnvqJKRA7q308NORJ2uCJcMCJEuYhhnHj
fYmVPpzYyrBWr6PfJTkUrgrAjFhEBj/XTzfj3QD/pxLISZP/sWRogJTwsDWNeK3v
y7GLc8TOONCK0IxkBfK4KRqUefCPYZW7n+tyvkLVfima2MDTby2cbleTPt2EX0YU
O/iow2C69LeORZMSHjjNokgOI7oEXDKbuwewpLSf8ly1kYdk4LZ6eSTnNVfZXoEo
8BkRMISK8TbQF4/fSK8+pdAD5kU9cZPHsS7cNcfc3zclXPFbjk1j2anuc/DGA+dT
gqFiGs89Gjtv3ExcdofUureEC8YcsUWHGfJdoZhhT7teCEwalJTaUjHLEWtWCCEV
21jT0gUSnW1MjttEOlQwXGiVdLAedzuF2E6qUG6qPDM2ihKje36J4AILPWnzWHTB
KyQXYC34TV5fAxDnx3vNa1ciMcWGCRa98O/3TjOVC4wnU+8YV93OGvlCBSWZd9VC
ogVXz4umrcHBdF1ztEKDUrsyHkaZr7Nq2Im51Si0TBHYg5BxsqLUvEvtYKC2AiRv
kL8zSY3iMhdU24g46FCuzX4vcAvd0iQpHuHmlTrP0biL/s2pQh6tmTdm/mSXlH1H
vzSprluVTKhcvBONT0feZYvFvcdHzFjWJdEmSWIik2st3o5YK1ecR3lquNkzsrtN
s4QUi5rY/F+Bpj5VLkE4jQ1G+SxNO7wgIyZpyfegwQX5+zoplGrAYe+UxpwdOJCs
Entdbfx/gA+T9WiU8IodldHP2DUG3dED/qv5CDpj1EOvuQ25hieObGCc6YAwweoe
WakhFuznQcYRj4CTLDA/33/h3pqjDdYvXerpFAG0AQTBnLCsS290g/qXfKu9nsnx
3HVNMFCU+g62MYzB3bumM/aWon0qQ/bdt/cw9BGqaLufvsUmmFqRMUJbtrbbNFCr
v18XdQeP/LmpcEcBGM08quUvdjpXc+OKC2Gf7f9K5q4jfqb3optMcnpAutSbfiQX
dqwOm0od1auz9Sp0uoHCvA==
`protect END_PROTECTED
