`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NkZIVsnHABMwr9nbPffD4GOsB+BiJ7hmgBTG3mPIJqU0bfgZPyoqoY5K56hWZFgq
mzK5dBeywc6mzXLZeQgmUYbWimkhY2eveUGB4OrnpByyiLKdwArVNwjyjY9Ye0HP
Wa323pegKjGiaoX3i88je7AmKBxpTnR7cveBYx5INC5uuGkLCBOHHYAc6jWhL6ey
tFEWDQfJ4N8efIqqK2TOxpvE0p64vaDS6ZD41jsdexy3FwJ/imtMdu08Z1v32/2p
1WGsIKJ0XJIUF/LTxTP0TWPKMIZzXsJ+LLBZ24waLwEgJi3edIktFwJDtQLzzlJ3
Mf2uBq1UJQ0uwTAA7W0+w2EZYIEVTzN7O0npvvBvRGZ97AK3GEGAnagDN589urxb
5FbN4yon8WDBdpg1+7cZb7SVCnaMg2DmdYPQ8Mxci60Z7yV0sDmsI96qnH7qz1QK
NgdeyYxkIx69ixw6QPUrWamZ2QHTgq34xKyxIw6zcJaVqgo6Hq9RYq8AhMvEcuU0
TnMJAxj2u5Fve9GO1A95xMeWeFzNzNHR0HlzTGR5DUWBCHXfFWCbR5/8VsvA7x3K
SXmZPBDZ5NQd7gHyL6jWJ91YHgU2cjF4a45YUeti4GnOqAYsWFKmH+TbS39ezrFz
bSDUG3dgwA9zy6OXuUv64kQl8CZCqQ4wrP9BAhntV3/I/meaUChnTzMC+w3qjvFs
NfV/2AbWLSYxJuZ2xGVuixYCl3iNtoyR3Plpq+oisgocDVym54UfdlW2LlOb1Ze/
kYqIKtO9IPYeFoEr9+lY1z0GP02fQMhSprrp8Sc3iw+vh8Gv98O5DKVczkzSUJLe
1ILXrdlC9z5daS/E5mCYSdUrGlhXm9i/Vj4KTjuBGrzHrjnVz4LF1z1mzfRhcyLa
82fy6n1vBo2oLW+5IcYLVSCwB/nXOu+GU5275LpXebt3gGuu0ZpZoZILTHPq/Ggn
vQNUrECTnZzFkGfGHr9DODlY8JNXeBxtm/NmyfmhfcZdCnYHjbf+qmpUHWTzv2NS
hFBbZ1rk9ER4YVWTvDM5Uu/PBsM21/e8fJCbSg375sssEwat2SurxvmOtHAMIFYG
enDB1AAqsuv3hvA+epm746Fismw6wb58OJEwaboDQ9Q4XhhiNNBfQy/d5/U8n4Dx
M2rmOwURO7Rj1aVVi1fdYUKFT9CQNUrnzKx50RWo6qy+J7hyor5vilkG3tn/ChmJ
W5IvWU4Vv0owrvQflBOLUXxmo+YZE+WBh8aOSlksIUwJSARGQiicizA7t0w1GRKW
7jL2lEgevNvtzB47cMPcEGrYDeRgMUJ6lt0UCVSTaeSkDc5wL2VzfpUXcHwmh7zy
KtdGDE6VEaNhZpbJPahTi9alZATn1wWspvV1DYNYR7OwyHrdMpRJjx8y/3kA3UU4
dOGh62LUVwNEVpaQo7Md90YK9sLWkG4xeUgCFeeCDuYmYUKCA6hNfAEY+xWd4n51
1uKgtRzTXf34TkmSTII24W8G8gqfwxEwgW9JV9Tt7OqY6kYD5Y9Ufd9SRxAbtEY/
t7IjN8e8vVs8IzUbSdedTi693X7ZvoIQthamgz6w1jl+0eQBj0REPIBK0fjmwD+A
+s56Kii7OJwF9xPc9342k+1lmiX9XzrbIjjsX2UVao9vtPhX6RqCE/YpeiGK5zGd
kbKDudObvrIZ82JZUzS3wnyuYtsTAB1GpyVDDlS4KriQb3Cl/TLLkXR2B2pZy40n
2WoT6M8YIXZ0qZN05h/0iNCRkLHaOeUGcwJ5pvalRLU7y48UuTGXV107R3/3jgUs
u6t1FZRLWhvUbMc064B3f7LRi9RD9QV0srrbQxbK+/XT5e6+kwfG+kie1RL8fdjo
AM9QLE/S2jI3XK6wMhxamaDSYkr1UWernur6SoONdxwphOCjCdsJiRbp1PPW1tF7
caSjgh2rQ+0a7OLYtPjdsw+5YPPb/exdbv5OO7DJy0LWT8Q58m2IYoRIyNz23ZMd
uU4FbzrsATwumbDGvoOj1aXekyUVfqaxcIwlQzTF+GAJu5NCCGifT7gVM0OUPzPr
jtS7/zOdveoR5XarhQM0AsKAuYTIIycqs4wHgR7mUn7cYmlUVU/YpLRKu0FpGrGC
PAnpCgRLrAHy8Ul0QxzT5Te0cxpaw6MD2ylWyfM+lJkwwo1xXy7Qb2NZOQnWhkWv
ieCn9BLKv8actfVB6EXx/LQ/9JhFGV9j//FitJtgGI3BFwDj0Ifsk0kYUfjzMEW9
zTsKm0wF6uPFOvLqoJmDa6jxkelq43WzYgQSOgi/8H/idEaN4clmc1NTsQu5HSBW
63NlnHiQW4lY6aO3Qbg9C/jZEC6SQvMIgeiMajv+jcwn8Z0I0U0qbtDHRkdAb501
IPldI3y3yFbTgxGjeSAfB1bdSm6aYA8ISPzZHMddva+M2M8FOjul1ST2s5Fm0SIl
vGTXL8fOSpqsf28yfaJ89rZe+gdpyDZYyYXiqqmLe91fNJnxHZDhdy3UZ+N+PHCH
gnEaByRYn6ZI0ZMO+4+XMUiJg2Gvx8DBh2mU64zwRZM=
`protect END_PROTECTED
