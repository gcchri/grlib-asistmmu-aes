`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fd8d+bpPNbfRDlhPiPrm670luPetXEAGwg7RHDPLcr7E4hvnR+VvskD4UcpXzn2f
MX99v2dF+/lguDOI9w2qMyB8aR7kN1ebC5+2CV9FutYEe5HikD+29vkSz5eZXVnr
7cug+sq3jMfH7FVi7Zkg1eJkUAr7MJEAIdPOJMtyslTEWGwGsF55fQYmTDm/WT7O
VCwF5mHMEev4gG0GJD119NHA9snK5+1VtvHEmHcppDZ2zf8h6zsJhye4srRtw2iA
Vw9kgN9gq5Gtf7JDr5GJhEd0EHgnAApzdxge67Egi/olFSFnjpaCc2QLYWabf3Gf
H5u830NPYV0E+AeWbXs2N8rersJK/FEH5oQqNAvpuP2661jruY+0UjQkuV8zhddS
OGLsul+QvuJxBlUpmvORYmrdlAwJ9jzxPtmjCC7+1UWS0+mwYCJGSxUsFTbRuMqd
B7HKYbxxInLPno4pFIEvgriDCjocUFnKRfTawkqlVCbQ/RlWThwecCphOiwvoZVB
VYv71sBqJ87VzjruSDhMtfBfU3ePrT8dAhCYNPPRNLgzp1fjjFUDxzxATAaIqozR
7NDUAzZxwdLr2uVCz6VJ2otGaiQBx6O6BqTddGZzlzbY6ykamLE0yfEAhW27zNL/
Pz0QLe2Qud302kzkvNb1KbmtNAl6nRd67/9PK3bUipIjpXIznBWED6ZR82dAmJpD
UrpGoiqgg8wsAG01K0qeAFALGBWkOndI37lvR7D1zUllUJiPwZaCe1JpJAcx4Ujm
zkFQSEx2Ehes84+jiKVJVQRd3IvqxVQfxiKYaIDQglS/e373A5m8KSSKegWmCfmn
1RVa+0gt9q7y29F2mjVGCnj2iM7bD8wKjDaRSdevq81/rg6VxM1468l36wCN07jr
rpBx9hyMuuTzFq+F0y05Vt4FOTY4whPBBUO327DxAASwQ4jKNVxmir2hRfkKprZP
IVFZDNaXaprPDYib1L85Baytef8ppqdXt7cm48CD5VwFSpDNFls474emfmabUzkF
AQ21eymIKsvqMe7opMAxZiLQvzyc62hJcTgsP2G9XXRMZJJsEI2d26vfP2Q4u0H/
4+eVTS3v/wtyodMXQfjWfU5wfYreA+Vj+WOHq69WGxvjG6b38wx6N9eKqT/WangW
TevYnR6sukCpp1wQK7mltvGiyV93f7HLd9Amka7rzDL8D6jw2UsbvqQoOp7vkQww
Bt7nwUfVGSETgwk+GL8c/gairSGLcVCDcW6QK3SGrd7JXAy5cJlueH4KZjp93vL2
OWwA6/uygcDxQVk9E5+yuowUDZzLsp1urV3JC3kvQTPHEZWEefvEB/mMaUC+Ch1u
dlx6rr3gdNmALZY4pHz5sSkxNr7huZT9XDyjpCBt/6/0fPd9uenLAevCr2bSw1f7
rZ92qDz//nAzUtCPvAjLph/0u6EBPFaCgihSYLtMPgzS6JKG8s39E1jeEeyW4Y6l
A6VM7U/3a1TPXRrG9LAXSdDHqc+Ug4JawQP6XwwtnHx+svH+MS+W9ZIqrJ/lXWkF
xQE+MKxY/Wxk9ZgqZMbTs9y9Pm608lvpUh96RgIhih9/itwyTqMOAtOyFLzquhN7
EoLmPWBzQJmlKolPxsP0HfV//i/iCuyky6D1wyADZwe/j7rDIgWyZxUYe2od9VYE
AsbwdH6zpWJk+irv4YeyiECMYiJE3IL9DR9BmMqSDB9eAS00BlRsnph7heblg4F/
4ToUX56Hl9XzWQXkxnX80jxkHNcO79WVONtZkKOV3V+7zpA9qrRNXqOq7VpXsIVz
0N1icU08Rn6RwzsIbe0gBgi7QorNw+qvkMXfoqwKW8VGRIdEm4miMPy3/QxOs09n
NA3++gM2gi4hRpSRS6NeaCLM2phJY/o3isfuK4szhg4yK3c80qxS5bt7u8bj2m3Y
TXtyxnzWaexTxVW6sVwVIuisnqvteO0S8yRZQQyv4zAUlntbchUmgrf/64+u+b4n
AE3GczMPx0aFzKTwfY21t1q6JKe5yg0nXJXMbvP0kX6VUEMBk/JlQaUKVXNs1d9l
bYcOBWAmzoCyx+C8T/8jrRWoS79HDdTJTaxHbCW/5Tx6z8voVpLVXBcYqZ2a7vg8
BgKL+pQeypjQbXmxxm3WoWrzF/9hidRTzNeuYL09qF1j7Fa2bk76/JCAsQ1e1kPG
iMw8bzr7vD+wz3CLxV+ndwyfA+6UgtkhR1b8U9Elvr1rJj550VAsqGKWdW9vG7Cj
WlsXsEmR5c1D3z5Hxu6fHXNu/FVMhmzH086XMj0v74dVK9HsXK43x9Ba/YiMJ73q
0YE5QoV+RDWf+Z2/YmNgJr9NM1Wm3SYc136T/49Pj87yuKJ+p1SW+NbXie9QpHmE
ryrkPG2HxptWcHpx2UAya9C9ut2Flxs3DtXj405xDxeyJDSCrtFf/adIaEMY9yHG
WhZorZ6VlizUMxKME1Cm3g/ALbj7JNOCMh64p6LVRRAwiu8x0hj3GAgBZir+e/Ci
ZlCGVSTrf0VzXMhDyC2VOmFJi4cBpfZDg5DFBKi+bAN/2jNpVNa+e53aHHS57hZS
rb9Pk5F0nYu4+eranzgzKJrPs6+yTkiEUbV8w6Lvb/Guu/Oz6nvmR9JLueZszLyO
f4I1hQM3wYKVarWKPQv4oohGDPMaQYiUz7J5f2IKc+gckDaNjpB1MW6cA9dQocbt
G/MUyxhInMny80GuObbN1BNpYcwIXf1XHStDbOTHNE8sl7e5+r0l7KUId4+IlN2f
RuvZ5cazrw23IJbh7i8Z9twA4iXqNIdHdkXzoy46uNLbnlc1wtjDExajyv1TS9W+
LHuQ/mDL5fWM6qLOX9h4krz3dk7L4tNS26CGpmW7NFFD+7spcjleHJygrqDBtEmx
FSRAMpUiIp8xlBxsgi65J/DSoibR9hAltc9Y0FWewgCnvKiijpLBi8V6QNLDf5hz
EAB9gFYuIvslZZbePoJnNulMWdShC10qDt+rT0MGtP3bWV1nCgTKTESez/qfesv1
Pky7ys+6qvywpk9UwF7RBQessjrIX2E1tVjx7FlwM3U9dR2TLAxwZ2VJXHcDOZCo
kj829mI70t/EGawncxcysVgybeT7i86PtJk4vrdXRC95UDNOqXR8f23xUByWyTer
sUNqu0G0ZMUeqWJri7/O9R7nkvAGjNbFNaCYIbiWHxKODLlt0luSsNb//a++JqJN
mwCZS5oxVr1Kl3KKtP1Pq8TUG8NNJYsKWjKS9EwH9sXe6D//X+xG+V9B/TGWgKYr
JZXnh6WaAc3znVFdMDRi3ntMz/gdoFVU+aEZeCLFuLHrtQSKklMmJPQ149UeJI4a
Y+g5LlMLKuxbJaw0Jz9Ob0PbGLNhWELNq16dr507MCV5ZSZM9D6zSIrqDnmxJr97
5AsBRryLxb/gGPgBloRdDyp1l98XcGyU0awRR/HLp+KXW47pjhY2sydx2HeJ2+fZ
uF35lOUnlDkTct/rFrrox1tVfFZbW6bi7w+mjAztoaTUQ7cRDcK4TsT6Lw+DM/Uv
puHdteD+O6IG/GNyCmCeI7+2HIOMA14CVFdi0bBv0mIW/Y0SDvGmAbZiOsSHpFiT
hIJVJ07Bta+OKeVOqIifIqrNAmVJFU2IIuWfAWYTVs+CKDvmSjPe4wFgjbl/u+7p
p+0kS7HcPO+HFttpIlGnMoWG8eh7gA9f/l8EdL/5SZUyRUEjb4GFeJnNIT6wBdGT
F45b0isbQJUI1MPDt1wlSyZDjkUC1BWhAoN54Y+gVgQO8PR5T9CJoltO73xJTh+K
DOjmcMOReGoSKAOX7Vtq63oYtU644navbM4ytCoFyP+jGkFaes0m15m740+8C/DW
lDPcqUbZF+oWMv2LoW8BbowPctD/HIdatWxJESh8UCEJAeH8YbHE2umdY4ZHQ/Md
AaMuxkU8j67MzqIuMworq5tjRC9TU5IPVNSmdlJe74TifuQuexPWxj5tQFaRKv9h
+Sz8bKrwM2ZzxPMnIgsT4u8e9yxJVFI+dgjW0hUI11yq1zaXvaWibXrSfIvIpzgz
NgrIx6TCusXNXIgOW33O5PD8srmNKBGNCSOYDm77HO0wEiYvE9Td4G+CdecLbtCS
Cn/UJrvLG/g0EMisnSHmVMMcPuz8n9uX8T8BHnvShvFVnfNZlE9lhl49aubgTBqH
zTek34sVwO/OwrfrpTiD+qtkxBjmfD6Ma8pcsmSnea3bwiJfp+UzFvCc18iSRJ52
H4icHkFIA5K7j2czSDNhXQ55+/mEKq0LcncY+WdU+CndoU1cWp94dXq8k9vnPUq7
YNOr1fwETfcVUQT7c5lHpVrG1pBGcuXpMBEtDGQBV+tzVHPglqvLAa4inMaP622u
3Iqe095iAVGdNcM7iGpKQn+W5sgRP+fKfAkFymOAWY7Ka+88YLGRxevRhHoK0dBM
+VUyCGsvkk0kH0sBsd3WiCO8NcZ82I3uyy29KQ8uSUaskrbKjogUJGS4gN4deF68
wijwHgCoNbNXxMV8AavZJADfb8U3kRNDsaXW95aHFKUvPFe2S2YDITOesu0zLfWu
cM8myELi9r3KuOqOdCv+q63fDBZO68EfpG5Z5NNjiKNv4YW1WZd1Lmu9tTsMvOXR
qT+mzT59eP7igAiPJo6xwzfMsIZIcItXI9GbFHN6ailQ9VlYRrEId0KuOXry4ceO
CFPpAcGMmW1gt2npqXNUb0woXTR474hDNINB59oUym7zH5qRxXz5XXpEwmsh/5Fk
x3unrSkUEIwI+73xKh0IZvaAmUEKPZvb24/uwYyGjNUpWk8HWx5pY6PrommhYnTk
Wg97QNxzJURPne8S/QPz77Qp/bhJJNmwIoWO9Vk0oecNFyTMkgo9jB1OZ5BoYCpz
fnwrd0hv/naVJATBAABdnlz7CqQ/GzRT77lDk13JIMFOZ+QIAYTWc3ZPq007Wpte
eVLBK+SgT1mZUupAk710+e2vcn22buRYDczJkx01kvnrwwqvz4i/ZaWXN7KwfkIn
DiQwfZ80xlgT5UWAjCEf6hP7wf7ZmCPjU0E2+HItCZn6xEohc6DuNRpqVB7FNaF0
q3za3n04tQE0QTL7IDcA6l0V1hHhMILaO57YQoNM72rM9I0itNnoj6qavm8wioup
yPWXQ//Un6FW0xCZPrq767eYDfdX++LIIRgtamKtsLdwa4IK90Kwcqd2+j4KezmH
BHKtg+6Ml3XVlCYQEUqNt+55WZK57Bpt9jjh9wa6EAZZ3/Q82fLpun2J2xZX6i82
Pb2kdS40+X5bI6OIFbYlQCuHAHGIddYl/WehvhYCKxbAkJojqWof+ESlMXbLiJxq
KQI8GzwVLbGsGTSCYIELGRKzcnR3H2H2amT6KbKRyCj1CwL3+Qj1Ep0y6AmcbNqJ
o8sXZme4U/iTM5E1CsYRlN+ZRHNNdlp/Z6IECcaUAt4cdtDp9xjdV1uQs4+h1rgW
LmmwpIwprUyqzl/w1kc6lyDvNT9gBd8z84ESdcQDgggKn1ajmPmfcBhZTIfSKRWw
k+37sanq7J2vhjjk0a6R9RsGlJFbb/qu4z9mr+vc2GRG9XMKktzFlQAM2LVI8xmQ
1bEjHR4Z+P0ewWGduGRcDPMmM8I+xv5YUrAlhq7FUhz27BRJPRU8WGmvt65bcWwZ
Ljs3cMrd6eLJ1F7XBiT/5h54enA8URKNaDGU37BsFwQJq92noySNQ/5QqKHjfTTT
wa57a1cnFV2oeR5ESA+jK2/zSckv2UEFGDwif+/fWXWMVktV7tuR5KzSBsQlzV0R
0EGCOwSPymSozo78UVleivS3BmQRHCfASf4QRl1JHs1yQxIe3jlcDna8cwZztt3K
xLUmbX3qCfcO05kUk7bIULdu9dNl4LQLyKj7KQ09qoUfqRIbgG4FoEdxvJGMhe93
Aj4hdr0kAhQCCrkEvV/uUXyZvy7qk3Irksi311QZVprfstBT901CIW7jA70pZz7u
WUmg0vQ+icrFhzypFId/+0Io3+LqruonZgiq0XOkmfrsAbGj+v93tlR7mAQWF7m7
x63bnAcaeahJ69x5nURaW1rESWr2nEndktkPs80k7JR06L8blpewuyWdniVRrkEO
JNYBE+1Shdi7uX7Q/OIk+R34T8RKEmITdJhAMeWRMNfcw6oDENzzwoqX373JLzwc
H3PQqLg2YIah4g88wmb1TFkfl8K92nnQP/PUxNufRBPxa+O08jzWKPF4LsL2N4tv
NMKcl/BKgIk/GePd4XAs4UOhK/rMQERQp7OhS6Z0TG/WdLdLjU+nGIN4H4ZlSnyI
AsmTbqtPpNsR2FBJov3EQ0Gp5EDmKOY6996GW54WU4dWzcORmusLX9WeLYw6lj8r
M/PvdGbQz2oA0bxYAU69Z02PuvyZG4r8q6VtXol4ReF+m8mI/ZnN3eY1zF0HylAG
1lOb+NLh++8RlTyYabeV9a+dGyOjolbS9qluN4QQu6woaaBrY0eW0P/a1CNLtYS5
niJmyDy3HEsLdVphGl9MJotYdsCheB+zIdYXPLCE5ZArfPNm4aganJlcg4bi7ww9
OYo9YQL0R7ShRD9Yjvm2JXHUd3ZUwDgJ5QJdrA9WCTkCqx0i7VZ5vSsQUSs/RPmB
jbnDySVLUjQFB5635ROUTwo1FDcgnKcQdM72H8HnC54sY4wxlRichT3P60vIP/qD
CfUAZjKaBZS8E8BWQMhHNa+9ypUluzNEheZc4gjhbdD0KBexy3jdVMhUVm7tbyMq
By4D0O4SfkGXr8Sxu9rKttxbhsO+/Z2V7QeeSX7Qc7hNWFMdTuAwRxxETm98ePZs
+YmPmN5y80Sx2M7M57D9H/YKb4i39gxdUCTGvi5TQrI2Jk+/nZuhUmdMW3+3uD7E
vjdQQrSeiJIVdaclRu5BAEXlPb9zjrGGsptCY4YH6gPO8cH5pdLbZlR1+34Qah0E
9HYjXCTlEftsPc5P+4fnh/IILqah8RROrxFGhfi1ERMNV5r5STJqjuisCK+Q2OQ2
SEsWMh0ounpCR9XrQEUFs1W0DYcWv8uG80MbcLGEYV7YdA/z5XB09S4GOUaTcBCd
ErpBTma2HwzE9M/0JT8yC1/LQJVnZUHFwkuvNbzN4d+ZPn7P57KhZNvnWuRnazfZ
4sDlLJpeyY/BsilPHuvS2Hx/Wha3RUZmI+ZWEkqJyzpsAXErtYDQRi7w3pC0DVDx
zFqVLvFag6SryCrT1iXYDkHsojEnHLqzLZads35USOct60Zwn2hDNZjE6otizUQ1
tudJKGUaFYhyZ//JlDlY2MWMxvpgP4GRpV8KNKA6uxbyuJ7gRqSjOcFiIZOnDZ2B
q1l6VENqIscZawL8yyjmO2GJMr9GwjOv0/Rox8YfkB+8MAF2PjSEx9cZs7iRtA84
TBBVxlPHO1CLmT4unehY7q6ScDQ4BeyCcPg1XNc8wMWOtTCPKMT6KdX4I+qJUXyp
tJvhY0R0s2xxFSD7gqAlfQQ9k4hmZZAW2vt8BaDp7WHsASowvfpIrTtN+D3ZT6iy
RbSi8+bZsxhwlV0dbRQ0vMEx/7ONBGWake43d44CP5n7Rlc890tFNl8MQvmABmfG
zANdLHfc8Avipw0kW3iLSWjoqu/EMlDK3mzEYzg9hY7S7WkaHSXiEzDcfke00fpA
kcePKr6CRraIgfBhkwkGqwgrsluHui6Jt3K58Ts5KYKH+I5QEISgguBMIE9Ox07Q
IggVcUDKGrGsAYBhX2jdJni92kEllIIYszz8ZRi+JQtWZCaRaLVsiCTTKkz0PjjR
i3pfBaNSFHgWYmLJ3n4vg2xJsEEJzXCUF64ZehlvWfIq5vN59qrXGbsYqme4O9Dq
VPzKfCfr3rbB9Cqt2JWdCkOJtHrlOFaWCKlE4diCbCU=
`protect END_PROTECTED
