`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JnHqi9sKaJeqFAFSOERxmpy+sxyXXtEvQBcSkYJ6R4mBWMYz5JMIuvauvs4smdAw
gm3WPQ0Szc79s4YOdZ3sFH7T+wgK25INdTLWAGANaIRSDP/ABUuRHsIGhJVKJAXT
jEq3MjVN5G+QqjXdZhydglPEjC6Y83YYF5WqfDmxdKYluqRouNBYYWzDHI6e45n6
ODkoNEYivG18hYQh63fRM43IE1KRc5/LOMWVdp2fj7Iqcs1eq5uyVKe1KMh830Z+
8ns5MMDcdXX9PkMGKfhP1PghyWm5bmnRr0EbYpIegimg+L0ytDqfX9KrlzNZnTQW
Num8flWpLf6F4PSd6YK4HiaPTFuql21zrX4i5ynSAP0q6ftBFuVIb1/BM4Nvf/tA
DevxUpp2ZJ4+Re3TSQ9CyGAQE+QI/9pX3QCnvHqEnLU=
`protect END_PROTECTED
