`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/2Tn8wG00esFmnvU6EMhTvD3AlEFssQFHNU+FtcZ3z07+AvBFkXkMKajjzUf3oLi
durjXbel17jFSBGl0AoeLyULNhyLekbxRP7ZDRlAKCw10SJVO6ZOjfKY2kqyGR50
2DSAGfF8HipPrfi3oiGuU3JWOTZY84myhGOu0l09dpCp0YS+GCZEleKo9wSALIgo
mTNzhb+Pgl900L7brdb4AOLUcZQr/1fnQCYrLAhqCaLJ8kjw6by99zF01CKY5w6t
uHFQ34rJQXMkYJiCs6BNtA==
`protect END_PROTECTED
