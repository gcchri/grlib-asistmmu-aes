`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+H9XlXC9DjbvCRWVUo+vGvjzQT5ncDqVK0P24KXhG+/01RplQzR7tWRR3uk+q2ir
VZFIZ7gRSy9RzO1c6dREAJFg0FyjpO/DdkNSxgAolprZRfgiorXzUdnBSLU3wHW1
nC+7aeVxMsc9AqIENYtPLnzegMT4fMgWWmcqKomYJfV2omftxFD8bSHl8Pjatk2i
TtGGbwbycIMvbA4ndGigKmimS2eKaFcPvL9g/mft8ds1ga9y9lkBVw9OIPqUjGL5
WEQTmIVioAoRVRYvIxiXW6cLrXhPedoZXp3sohLaxipB1sBGCEe6bEb2ANn8C8hK
5Gz+5b4oPbcfQcfD6TQBPQQUWhTe4Usf2Ahf0pR2RJWkcmdQ4i4GKogCtr/W6nCw
pFNQCamB7jmOAYwm8nLVCg==
`protect END_PROTECTED
