`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dJixw2lLSTlZlVszJnTcIbufVXgYPAQwVyZTQG4VichikOvof0jeHnQu7ehzeflT
PqLpITnFOzsYFEkWqbFvXUlRkNgR5+yLoydKICpGqhhfBCFaVdyDxqzx147G31k2
0hJs7etKa0FfmcKPZcGtlawY5NbtmFzdnFHfoAJdzwzdBNeesp4of/f5+rT+8h2D
JrUXqoHyf6s9Rhr/4G/dzzAkCI+xVof6rS6JTTbMrjh+lziEr1mJ2ji5SqhSA1rj
Of89QBqCr/I4NBs81us8R6u0vjISFzkzgeNW4khsjO6ehQ66kYsycMFi6LkXSWTK
thhw2ViIW/rDw8ukS5WLiCUpq4OMsF63VaQVgcUYdQNEHl9XJDRnrAoWdY4llA1t
Di4DgICyMLCiwGlfkuuPDX0IJCxLCTDObfyCsx3ccc7HEieJL2TnMzc2Cm43MHm/
lcJz+sQbe0asyXIervd6+ZYbSXHm0ap/HGlxqi2V/O6IOwa/EvFf3LQenNymteUD
h4fP9b+aVh9RxB21982kQ74Y31NCS7BP8UTXI2VTNlS8smKUuqXoeUE/kdGZukeY
LOt/w7CgFnsUGliSF6xGDAqTLkzd8aBf84YCyMvm2dDorZvytIe4FLLqTF+dycpM
/xAAYLQ/iEkpYQ6cb2F1J1zzbSZFV9MB9q1gV+QVej3xSSE2pQedKH1oOozAynlA
Uz6+IfOzkcdZQy2hIgrIopz20gEefSpUXZZIoSjRDpK9JHD3wGiVrIE5cJRNv1jW
fF2MtmwR+ty/vu83ywReMXJWjoRI0sv4sgxNANRp7HMKfV4TqmkBRi6Duat1hTl0
SFoheFrCcMzcjTdYCdFWbbMFgNtBttOE+gYhams+SgIeii5zZ8jlxbqMO0gHFK6k
uhHpPFVOjBa3CJDrGtcue8wOgBMPoItyyGaekIeJW6KPZ4qXPkpjS0yUxaoHaMoK
3gpqnVWmumIYn53er7Jg8cyfDV5gqTqZmfWCeps/TFy7h3JjEaoCmHYhY98k/rwZ
fSF/MT5/cUXeABiL/GHJWzyG7FKE80NF69ZPcU1UmddIJxcryVHhYdrsF43jN8AO
TgpgoNXWDAMfG1Fh7qa3wQ==
`protect END_PROTECTED
