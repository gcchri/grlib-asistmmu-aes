`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SQjQEsoxC39v3EDTCjNHCTmkscsaOmk2NaxmOVmb5hwFWu6Rr2opnKlDsjhzayZj
IQTUt++gcFj9X4BbMEKKyShSGfLBwhPBDu2h2pTsoc2qhbeGtc9lf/mmlWResLP4
Z6gBD4+VMvfUGxuKjL/kf6pR1j93Uxp2JhZsTVVRiE2U0cRkw63yGqaihD1cFPsL
fHLPCqoYh4jEMVlFFTH1xcOdLMi/otVW42of6Pxo1StuZ1sAfACZUgYMZ83MzJAs
6IRJka6TopsZezfEfXBITn+Q8I0uKtMCM7XLIwiwEz/qTQQpXw3pJIZdC+UdRjFb
5qa4pYkwSPwM0UrxuuSXuf/IHevRG5X6vHmrme3Bm4JVWgCe2PtrWT2w1yw+g3tL
2gYI1nbBHFSrkNuwuSRb4ZV7OOdLy86IxV5NftKiKg4HCaFK9jYEihrw5IGRO2J2
fwAMm68vBQDEYQHrqhyTE1xDD3Ydfdo3hHiKl42v2Dcsgo8Mg7aORWPx2TXZrFcq
lFBekw40SyS/Go+aJIJn0LIJudOofTRjFT2Rg1hNp2SkAg/BQ7QcDsTCny2DsGg8
1V7iEK7LT3NsNiPhJaO1HuBTRji9tIrp37au4sSR9hEH2YVZuB9WjpwKgVfOeC1w
agPSvsF96YO7/jE3JL7fPz+9lsRWQRFIzZFN6og42jgcjFhRlqBvfc121HSuGkgG
keNdhK79MnS0MoYojRbxfayqxW2eM+uHvWSRm1NzjdhW7Pvi5Pf0RpP+o4On65L8
Hcva5M80/HHq9472yZTM4Ym8k37iZt8anOZ6w0QwPYrheefEd9mNvjXvT7IlCg/D
`protect END_PROTECTED
