`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hWHmSScUlaYAqHBOB8nXWLnPZlQswv0JZKbAD/5NAd/qRZMJI/cJd/n9mnmh2pof
gCaKOkpXauAGZLtlcJfuSHoDV2svJ/DkM6mEsK2qlz3OVPA+JFyxkZA+bnsYSnu5
s53vwKbT1kUMPGmI5rldd9OOWinEuEOlckXfXMQVF+Pe6uyLoWCpmO+UahXJdLb3
3J1Ur4pgqFFuwk5qUYC20DOEHWoEZRt5JsMb6rVmnz6fCG0wz3gDkA7484PjxFl1
wbIrJ5XjmZRDYpvCR3xvjuF3YH3JtsQ2QQ5nofEZjzMwzSShDlcRlxh5GK2wdR9M
0jnTihbVKI7rm9jcGpsGrJfAT20XB0D6Eu/d7KPHh/ayOsdna4PFdGppdf/9TAEG
Zs5ro0jeyfJGvEkyz0KG+ygbxEIx3EXbeQruvxAJ6dBLeesIhyappCJiOUWRaLpa
yDs1iM60P46+70dM4BFoDjryipDCjytiVC1Q9BVI3LQ3u3b7zRyVD4AgGzyXNVId
v//CHAzavAOIXU3KW39eNjEy0uv02aOfsQ1alXPSsHV3sJy8fVKq7sB5mTz8A3T4
k1oQyLiCf5TruqxDhUC5zhXxi2U43Q73e0QOxPhC3iwIHh9VCvcjaWddnXrcCshb
xJOxfPrwh19u83K/LdI7Ie2BrF4r+Hvtd2XLdc6eNdv+c6sf378ataadfThF9jea
dJxAAHfIv9+6jm51ILBsVlLj4qK/gF4jrsgnXXjjR2Gd7gFJrVXac0ra1b3r+MeE
QkrFswNPy9216ha/SFkw/A239xHTRp7goOjjh0kOHoV2D8L/hdQ/iTrNpldCPG6i
sdKoaGaZIQG8xSjUPZBnXMw5Hg3vyeSbVzhUVkzc27sqwEe/lNqaDP19ngVBhhRn
9b73LS2AaZLFeBI36kpk/s1LowqWc4cL/aMyr5mgIT4=
`protect END_PROTECTED
