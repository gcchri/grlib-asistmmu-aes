`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BQkiLitriEAkpZQGoj8IKv2GTHyn0B1sBIHO8SsRQRrOuhd7JJyklN2ZEVr2dO9t
9zV4etLo2s/iu/of9Gy0KHEk/S8H6eGPE5OQysDl1GxJlS5P6lKVRxP1QT1Y2Zbh
Wv+oJ729TWDyOCRC1WAUkGM52b/npGUrnlBuN4gewSpxunheD6KuwRzOz6RLEmeB
TE+BpWR4tCYfsyWljiBo1ozkMhmf1rvgCuCii9XtteabtyvE6OD5WjTaN7ndSGBH
zISDq6I7Vz2h3jyqloRyOeCjBo/OPpSvWl2y+KlzWXVKHwJN308arxqoKJmwUL+/
JpPngqtdcY3Y0BgPoMoiN8cNpn/HFcgBp3MLkZorOo+UvbEoJXDPPZdoSxEG/zqS
kQrbfVfJtiwpCtk6Nzt2ODTVQl4+n1mDkTB/h+0hcmKDOTk3JoYnCB8BWTdrCyHD
THHsJqfUH9vo+yDsVth2i7oTn9BMIlZ4ujgY6c+n0OI=
`protect END_PROTECTED
