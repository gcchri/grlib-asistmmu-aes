`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PWpwfdbQ4kQaxUGepKFPB3Yzg/Wew5+y9c/sarFIk2sPKexx3bWxN+quMWu5GjG/
ozS1V1YKlOr3Bky413FAjLSd/Ahs/wxv5BF9aBzCAQinMLt6airopfQFqA4z05qQ
mCI4kFLeyQbHD17NcpZdE/RDnhlvO0Lj0niMVniiVG5RA49zjXtrTztEHplTb5y2
ksyNdd4i/1LAJCCk8m+NzW0LXZk1tKwzi7zHfPE0OiLbETJhPaGmr77RZLdbslcm
87LAedj73T57IHcfnnXsWTh6tq76FHPtTiQaSdvqAxnyrhQxxJzOKql43oj/rM3x
H4mPgtSG4ZEEL51KHkfbA0SP/C7vwT/P5SrIRqCzuxt7u7AuaXPjcmwOGrJAjx8i
NJ8eSxYg6t7QcDY6pXvW6BZzuuZ4nTVUrUg3YH9yZY7dCbWfPe602ZkDelf2lP39
ZCvjvjw3TQkfRpZcPX5V3OQVLqQ/Sn4rtjekX+QfboXlOWgWPiCH9m+DaZOh/uqR
`protect END_PROTECTED
