`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZIH6k4nuAC/3+Q6zZVk3Lx417Ng6Dc7Ee0eWhnni28ow0cSkugXBoHR56+DTy0vs
vvODr/JiZj1Rz7+oB0p/8+nNsrDeuY4sxpUKtUMOlb4aZtbMqWd8kZ052C68RczA
/D9h4hLJtb39+uXZ2N6MTm92hLPLdI4sVjgCfDwwoF8bY6wuNr7rDl7HTcYjuR1/
xT/IzMhB639sLVXnLA/RU7oofSDQur9hTz5GFnppyuA8tXoLoTZPJt4+KDi1gBsO
BTzoAUyWvwq58cn/pyQ9J1iBus/VuR0pYeeut6CX7cJ/OgXRESJFjHeP1Wm6InPU
jBwoQ5exIhQjg0RaZDgsCNjumINqiIctky1466L1Vcj0gzlsxMmJlnEhKkN/yXFg
ZUkLmrskf+GlYjnP3UuiqHAPoAsCVws2d2i0c6x9gj1w8e3zYKPKiiQGSA3KV8o/
b04+YNDayXq+geY94TGRP8oQNdXMVjBykf4bht85ZdClthf7Vzgi5A1kRm3D4yNo
8wBMwQbmO/CP5YwDxiWgho+Lj/o0wXSG5ChtBhaciAU=
`protect END_PROTECTED
