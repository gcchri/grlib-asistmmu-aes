`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
piChRqCj2Gq2Qr3wh/Fqodqt+5VZmSNhYsnkdcqjqbmKQFgGeQY5JMQqp4V0hftP
KdCRWztbm7xxPLeec/T32Op94MDo9ebtzNpNZ1CCB+puiItL1zBoUMin61Ax1aqE
5Ivkz9Wfj+t484Ej3tsgdkiz3UdszNhrj9MmpVtlOqBeIoTheqegZOswVo6PZjzd
QrHRdlPQXEjyWqeVccIsy73yMLn2lK1/yQG4AqU4KGpU6LHsmg3xXYufW+d62KIj
uS15c3AIQ5q9IU5tOSh08gljuHA9y4eV7bAk/ZX4iZ6Q2zmxs+NEsO+Rm9NioSY/
Yn7VLKp2WojXAhFqNj1WwsZUnd9xXUuBpbBFVYstt0/PVq2tXoUQKYkcrDcDc03z
0AhjCGS3FUtby3u9XhUBsq1WBOa5x2b0blLPmmcja8FQ3aNSSwc84lHcVdaGULRD
y0qTrWLc6w90c2Y0/J2J/oDaw9AyOeEWvSnaNxWbco0PKMz2tIsf5wooKM2sQUE9
DM4/ZYwqOXB8dEGPOni5f/mz9DednR+h5vpkFnolwqkpDJnmMhmx0tQUvfje/sDX
eF1MZq3x1hVt5YlBGSfVtzxmaUTDLe6EY8O58CLmpR3kbEQNsRqenKNtF2As2Qix
Ku5MdZoXQZt3siKjxbjSS2RqPvIuV5W441kg4IVSYQiix6+iSSVcZT1TqHjdgXta
J8pUbBS5AtldHCEYLBRi9YfhSBExmCHNJ5X3gi8K8y8DVNflDcc1PK28ySl4gnTR
LEVIGS6OkZ9GwFuTRRW2vw==
`protect END_PROTECTED
