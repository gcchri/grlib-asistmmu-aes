`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zDnpun5vhvW+PsvG+gCJvs6KSIqjn0a0BVX/28DmwzyQibxc0/SO1CHgerhxHMxv
5OWcrNucZYZk+S8NcZzs9YBMPyfci09ep8O+AvwjLrsudi5awQ0J8ZkWkhZLWJhT
fdp3qarcNYQtLEDBr7Zz/+PUUpHhC5H34lcznbNdN+0Hc5JIVojVrRq1INJqfVL0
a2ZOuPrqYQvLu8ucd5LMckA0IvjCWy5dbhuzcrkDEIGt17kcXss7bJDnK4eE03he
w3EaUIpchvakoSg7PtIpPT+E2GjSX6JHATwjwr2P5UY=
`protect END_PROTECTED
