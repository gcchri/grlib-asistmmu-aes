`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vgc8Et1qtZQH2HYA7lTC6ZdBYbjJkd1Za1F8gFUVpiXsGKYcUb41q+U38FMcQGyt
xQkMtvx+TOuxjFWzjoOynsMMmeSZXGQzvAnXeaKAPTITQBda784PW0ZXGmXshn5C
5RilKRBWD3dyQqCXlG4akliB3NHDL7GQc6YvspqW+eoscz203WhZemQQhZKwhU09
88KJjJiZvwOYLt3bXsxnTMO8poPhhz75WI7YoGWjdCNi/QyGs7Zzuks72to/jZ+a
f1HWnugqW4PzWXs+na6r/+wg5ZDmxmFKnmdFJKdFx2dk9FhjMDBjnZGBaopARHjN
PwXdINFvYDSvfzNjZLcnVlxrYgkD2TXHjdkdpDUsM2tV1ijOEDZvJmEMKdMvt/dh
GkoCAK8quHygWykwuq+44W1M33Y5pb02ruqYx/zpwRQ+tk4llKoqMvcxP1OOJ+sZ
FznbLLuV+gJpKb/saqMytCu+wfNQ2HKAhAhV+yTqzRCfAXjz7zgBsgd/JMyty1EQ
NBOA1NW+/Tjf6ypxdb32Rf8troSl8ZMntceF/nu5uZVxqv1Dprjb3RoqS3qYP0rL
jNeYv86K9Hd8B+7juxiMMBU9neyspGVH0DyB8hnpWThShDWu66UbTPC8g8CLKSjG
KKdyvZyvTv9QBnOrT0p9Ng4Pp9L17yg4TvX2vYjDIdfENKRL6LEMCnfUaqIzGn0P
+bd3ejnHzclMG1io55WvHE5M3BYvGPn+eJvqg71L2QoXkzOYDx9PHlXp3WeHB2NI
X00jHHOUwaTfjXT3eUdB9r/PCNVLbCQhAoWUL+qVootFD+o9w2gy+/pbUCaINPrw
CD99MsYjKpy6D5pqivSCisAANCgjCa+iaxMEO4SAamiFad9KospMJvrn9Eo7u5NE
tqiAJbOLSUbFQd7FzlUwrpsY1lGIVcqw3LES1xl7kiaT1ofd8w1TTPxQC1ZyWFAV
tlrDx4lyAa6d6FRfomUI1XEq/3/8LEfxVIMFVnAjVPlwq4Z6ns1GrWiMnyLP7Bs/
yE4fhAraKr4S09M2eaf/R7h2GIA7woo1h+RGVdf4TyChrQdgVLeFQVIMKBqQJ8Lh
3p2RZSt8O7lzJFVm/2HTmoi1sltyE1F4lFvVTtEcu38NThKyR3+9v+mfsmXUef0Z
bY0cHF6WY+r92H1dyjB2KrT/MIHejAZhmgva5mhrPEDOl1i0VxXA1rBweh9k573E
vve50/uY3fIC2yB3LakCA4j7nz7Ii5AsSQXhmKExereSxox1lMfxmnbYn4/zMiVn
lrA3cQBX2wRj8rPt5HXffL1wX5fPNUktamKc2vLGyeJutu8na0uKRHgpNadsKn+f
WSIHWR2vhC62xUQQwHI66VmEjNW1+PLmSgm7m89UqIq5wruhWoqx/k2AlfFsxfli
AvtLc30tYSvndFr73HXJS8rOmXhNrRK2cj5U9R+0dBh3WV4Ik7/w6MGxFH82DM/x
zK0rSS53PKtaeYB0xmF25oBFXjlrFt71MYrJ7MDuHKnklABxwVOiP0A/xzs5StbT
YMxBkKhphBz2bTu0Z315gDmNCgDoBa/AYku/mqVLrIJu2hwQTHWclHUFFcXGGrfL
anjfJ+j+yghqrDzj1ea9a4ksgPDSE78Af0BK5RLzuxwD0RUmKzo9CsFD5U4b8sv2
F6LuZ3dkuV6VRUQ7iMwTtoKGmYUL206WaejWen5LaL77pW0N7acLMLvdGDKokUL3
4lgi3C6SxHp66/phvThewETZyZ1PR19WcSP9xW0MV1X50DKka+R082ctIo32gLaS
ssSWBDWrIOa9W2gO7YGFaqNCdpftkNyd6wqzT/kbJCODplBJRQd/UV1mtmO4+SJG
eG47ke3INSZOxUU0/dJ5/JbswHDst8ZA1GryMhtVdl8dIph6lVgBlqzA66O6KbCy
O7xDrixUzNXkTaYebNyI8R/xQ48SYoReqJqDGaqZVCuuRhnBTebBVHJFOXlZXuB9
Of4vezp10vuN7eYh85EuW2DoiRnzNfqavhmI/cPCABPdxrBJuu5oSP2tWr9i0u7m
xFi3CoP2BKWHmYxdzHerOekkXECH02OY5ZZicdI5kydlrKGIXZn1+Ec0iBEMD9V6
3ZJpqG5v9mjW/40xmxklSLRSo3FzqDGF2THolDKgqtW39zsiXgOOAoAM9XyZu7e5
juctD5E5CPDgB5GECq4MqB12ugkssdC9r39kAX7KJsw9qG2is53ADAor4o2sracp
PkJ44Z2JnhnJRsBNEPmEZix2Cn56IQ4k6ZBiQQZ67/SnDzrQbRxTpLpwFiz4Y1CF
T0bVEqeH7Ejhxasie351T+qjWcAOPOAYWcF1jU9ORFBLGSWBer2vTnZqN5JN5uX2
2PA+947iE/HFPQ7lbq/9nYZ7oCUHHOmRbvWJl14V52a2lcAWTLmjzxwDX7jRe57+
bz4Yf1OArqucToJ0gWRanEjvzIXKdqgOP0TF7KmH3gKbtR0Me4Frl40s6AaF90ca
rVeW2Wyia6zLzGd9OUhd/F0d/v+ZU7HGB11WnvrT/ShKdGzXLHBdWGpuKcdf+EyC
XcQuCmMciF/Fad4+aNoD41nnmANG/JopNCBufcHdRGIKOX2kWhXfsNwFtDQJdyrP
4F9iuOsFKemdu0GWyUrZdUlqDV0+YETsrp4Wx22ge181XQ1olxHi8D7Rzxwul3IX
lTiS/CJgJM5FyBloLAn0IJ+rbUnugSR8Xx/jXUHoCM/yAxdQvvz0UMBrMFajRlEm
rBmBHSFB2Aal72lpKLnl0Bw8YlOrrseVayWZQXDWuCwYDFZ8DEDIw6r3AS9VqgR+
DhkakmBRq8rXJTOkjhMJXJPMOmXGacEtJO7qTBIvrms=
`protect END_PROTECTED
