`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a+9Tw0cZJ4DJzo7sD/di4V8/FaDld+HmyWhSDv3Gkj14wcctBTfAlrWPortCevon
LkyqySnrCtMZ48y/MktR0kF9Mk6nPVr1GkugXidfgAfp/7+nsg/7RqQ0d+oC3WEx
93Ua43auoxeJoAAptRWIJf350nxpDf+Nk+Gi0Dj4bNSW6ZQ7i9FG+oEqlt2ZSIrY
UNPaQNrb2Tec3OGAwc2af/TISoEbGQLw0BCZqyhtwITs4sGWmAEdknjr+U9vLqNx
g8lPupBHRwFrAmAj4U+qMVP7U4A9gD0nfILfR5n033djE9lyzwHiRgpJ3HmwmhTa
Fkv9hEQFEqEXk2GlqkTu93FWxAKO4UxFkpOJ1K8FeUaz4/z9wxHMzgC2ZXLN4w9A
fcTOhHNA1tu2B4T4vVovg03F/1+nfrU2cfcJHCHH54IqWsxtoow74fM/j8qY+K3z
jepMKNn+8Nd0ejZhQVUk0RfSHVIdJWE9tZt/HrgIzA2YK7NqrsDFGeJTmX8Lo3Pr
OhPxQ+/3D69RM3tPN66jlMM+hgsq64tIfvUj6MQIPEiXd/mzjv8v/hNcLDG1ezN6
tc9w/+TP5c0guCu8nCDN+TE9S9kRMl5+OXPWmyPwjMEXw6VIyCdulnEFSwfm66P3
66VM7bFRumcgWnZ3hcPajA==
`protect END_PROTECTED
