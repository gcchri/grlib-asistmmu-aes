`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9jSso+9zve/q0A13Vh4crqx9j4yvV+8ZLgThOyTrmHCl8shXEXb4UbO/HO6gLgRJ
BbrUjUTAdGz3zIvNffLVaRCCd8LC+6hGLlVCFD/W1af0MDOwVt1eKrZFpaoN64Yz
BaVGWs0VrWcLxEpx/rzwIoWSMR9V4/fYLl9O+kKqxAKeVMEYkEDAmCvj4rU0uVya
qIFy3qyahAZhUawHeHq/0RHW42+zT9TeqMdFKWSUpDcXDCGDwAe4TqeSDsScsPdi
CIpDL8i1HHqCiNZMPcM1xULCwiAoOzr71CkD3h9M+9ytv5RSHFEpoAdEd2LBF0MX
uW/HRklUy2bvj+cdXpzpPGRJd411FbjCz3polB33nt4GviLyJ8yx4rJK5NLUTzNN
asny3z4dvYHH5yNQd6JG3JNBGjqdB5ggDEBgQE7BE+em2JrA+KYFHK9/aDMwRE81
29oj7b66pzEfCSyD5OQ/aOY6uPalDXCkoKMefJeGyVCrjAtI+mVzvmeI+Hn3aXov
/nLT0hHQ1IR5JEuyhAM9mRKOUF3QuBk7cP3VO+E8W9CcGZngO2D/tFBJxEIEPNmI
edE1Y0coDS49IQKL7UW0jLU2n8I8ellWOjXkYMFL5k6e56Bo3j/hAUGKFCrfJctY
+3f1/1FZS5eBxc9NHz0EVjmuuc8apQAlYEK7fa/z0+qdYVoniCH924OSrZ3Qfz0C
TXw+Ezdhy/G7loVNVyNzlewAxudy4cGk1vK2dtdnmkaOgRInni8EvMUueriB6ibl
`protect END_PROTECTED
