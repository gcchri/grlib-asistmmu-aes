`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iuCGDsAxfmMYEx4o2o5Jj2KCQRok41tsBY5JI3LZHX4/xNXMQEeYMxMi8MXE6fKd
S/iNbCkqBtlxY0JI/c85uR8L4iB4gJ7onMRTah0jq1wE8OLvu/fEZm1/DcwBiDhT
+fm3d9nNuhMMhr1+765HlBRkfjqYm5asAq9oGxhIP8ArFOFd8qC5pvnYH19mbgYp
zazt61eRT3IelAIduEHjg4hc/xX15fuGNAvVKFZwQtbvaSuO5rFpDuNrANqI7T/N
rPLBgmXLZ749aObFXhjpxRguS3xA+SC3nAE162onWWJSDOyHjzGmcFPrDpGq0PTp
z7Ebi9mvFcH/ZwxmJ/g958RwSzOxawBBPTMNvXe7SCHr8QFeJ3oX6yrsDEkTWBoQ
XetUfhbcq6VcoQTua7OW3RjWRljJ9kYvggW2NBFLWGq7Y6YQYr39RNzIcNjRAW3j
NBuLx5odDAS7k58JA/mgtJzx+0Wq4JAfsdMED7t43pygIoB9Btn9TRbcWF1EqXrc
0Exs10FEfhIZCQMMneXYjPslWKBBX7T+r3dGGKQoRLaHf6BLlGyJZDS5MZSXTjnH
IuuC3BKv9mWviM2Er9N4WNd/rOh8j9+be7jX9dKKsdm1u6UC6wxBxr36MkMS9OXP
ET7h/Fp8CuC/4btuGFkQM27eJ+ntU/3L3swXXEjAET5j5ZemWbJWSmSTXTHwJzIM
GEOJ+tI/X7oquZN/4qNGPYhFlWjbFn3qJ69SiVmdiRlpsJqZcgv3tWtuLRliyt0F
5ARKJjGpizIhb7zHdGWYiiyWkQJaub7xzDCGzjVL+bvSqZudnEUaKzJv9qPIWC/5
ZlPweoKplikaJA18MTak5nyWSyvKVV4Z+B3Mo1iPTZLlIpLsR9OxcdwxTT8MB7rm
7uHtc57Cr/sG5fMgWFNc9o6IkonYuklYgy06zn1t5vVFY5sxPHjuDSS/3uDZq4R+
4bVi0NFPvQB/AnPMg0eM8YUm7xab+iW8qhlVACG5XThaXU6An1afxA/OmE8Lj8VW
rue0br1VsBKDAGPhq67zCAdIaSaiLIoBNX6NoNQ23raz5Iaug+7Nua3nvaV5r9jb
86bHryWIZ6wOzZnscv/fQ3P7FXSRnj90Hk485hAgTadXI0IqJCgFR3T8bjDKug6x
UeWeSfu9EgQGOCjzRUeUSf3zr1QL6qDfepWFCgOojna2NGDWlED8+31LJ5KePXra
sQNUqP6I0KkqYmZ1a+dftQJDOhdRNnuclA97BN+SzfH4TsKJ9mJ6cV5gFzaM1T96
ey6BP24hecDnDc6/6bZAGzDK55ZkNYu+MoO555EIW0DwY2s1u+S9pb40i8+dh9IU
`protect END_PROTECTED
