`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gHzvv9tGVxVU+yUPgQA9sZCcoJNDnhPWVEVqnJfzaPfWR6RI8syew/0ULjXTlOCo
Fdh7sNOJEhNsuMPsEX6+y8vfuFrWqt+KP9gGaqz5fgMtlx4otnFX5nSMo6+xKv80
h8pDrPlyoAXglh1g1Ahyd/Pfb5C3jkO31Wu5loV10AXY9woR8JhEiyQyKdLw1Kuh
aM+11HBsOKo3gn+Qui488c+tzFrICi9hSxAuwrGm6is03dqlYXYaavRez3Fx2XvA
Xtejdn2MmoMCRqbEHmmyoCOch7qir4nxjPgfYF8D7ZwYt830sqBs1A0aldGfZZ1f
8hHGoGvwD4vvHPGx1kKUzK765mytZWV3BqqcoKTQF4Qt70N/Q+bEfD34ha32Oydw
9zsJaCLrREORaRI4LU8Ayl6xcwaE/zCAkqKrbRnUJ6Gl4ENBPcfUIy5GZMUI2EqN
qZGSMD1iiOKFjr8NvqWiUv6100jhJVVklQkkd1Qq0wRv/VNaO6c7sFf+tlxc7SeT
Ky3zpzSH1INm9lJeMJ8EIDCvee8QI/KrQnsvajiOLXkdUhJNtTrr65ElJY12LyVA
CDUIZrX5gNwjDyA8LHLa7/+FCP+OBXsY2psoRxh7aHv3npV8NelvBPAxu/QbCvnV
3KVpvArX/G07IRgfzu0E0g==
`protect END_PROTECTED
