`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZKTW7nSES6EIdSkEIGYlKmz9aAG9oVpb/VErEjNKzmYwBrY6Zd0UjJJNxwfUHZON
3w2XN0B8WWfz2mw1LmV95S7WuXqaYKDI/E/sNEufiiMVg5CFH0yJno/BBJTla2qR
CiWKMXrxZmc4z8pYMVoq/wcGKt0JRcJb1fOxRUwB2T4TG1+btLww5AQgwONov1+z
0CHYTjeiOx1Z1qv6gA9cXC+V6af83KCNJFh3IdtWa0fAYoJdB4TkI3nBs2CwdoMp
I8T4lGy2mxO6zl0WgUAFBe2j+QOdjiPwInOJkZZ26nV1hzxiOWASSqS9CeJ4HHJ5
l6ITA2GNHrQEWhXG8P11iILYJKgveVeCuG3LLRfGwU0PDt2W0a6LgeSrCPS1OOQB
9HwQ3OmZjuUJRnxRhIScqFlHy208BTxIweuugSnR6po=
`protect END_PROTECTED
