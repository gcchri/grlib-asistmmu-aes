`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OkvbZBPVBrc6c36UJwa7gZkyN2slg7N4XNZxdr4YgBXXVH6dRjZY1ANxxeUdFTzo
43pzmVqhwGtNmLvTFvwYRqTcGZgT7CbgQeJze3vKTuMWNzh6CG99S6J0W7CeOpGc
sd7iz9dnxjrGWj/gQe+1GE+EtbmuNQyEFsSQr144fccZpCw3rp3dNJUv2a9WZqwD
lY/JcCQ70iIsbGqSlCQ5bB9gSbOgT2E4NcNIyQzB9xAYvW9HeFmnLX/Xn9nazCiE
tBkPCDuiFEbVShJw7wz2ydVMqewgp43Pe+nowzPNiQgoeSuFv8Llz+P+Rjzqe7og
XMrFMix/WfP4lHhmM1IdLZSkNAorIMd6huOEZI7BnuTs06UdH55ZnGuS94YvywOd
QZuWlHa6YZCo7ICqx8ie29dPnjEsm0WsSo/5Uo0cPlbZj8RmgMHbeSYnVX9gXCe6
ADjLMvHREnNqDxJWoNIavbT6cHfeBuqaZ+Lx8EwwibKfq/Anj8IJM4AaLmKuAcsu
Vxvv3ATHM58LEjmW0PV/v7y/iE5dHGZaRl/M8cSwS22WroV9DNT4O2bZ/DxCEe8H
`protect END_PROTECTED
