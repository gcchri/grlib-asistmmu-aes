`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MqOm0xOiVjPmYttWZV/Ae6sMHhVttlph2hbiOKrvWn4Ohe9Lqfj+Mkyox7DORNi0
NOUvpCWb0SXen4D5yKZ23FosA2HF973EFuL+z21d79jsTV4aWrqatJ7cWaJ648Pn
oIbfG3C6KXTgcDlYoJM1QJ3V7MsHMK1r2/+tok/46bqK6sH/tGMNEIfzbzmYFdiF
HkAYSAldvRiVFz7O05QlSw7P1/FhhP5qnwbMu7k+UsoLY3uGQ6jc4fFgKXdMACj0
Hd2rd3wfxDuVoHqfN/Iq79NLbqtNad0Qk/bVZ0CGDBvONHumACi+gRqewwRyKO3l
IcQjQ9QkN2X7NUYXHuF7H2tlXj4SKRsRWXE7zOr4uOnjUfe4blODSqzWU7BkfdPg
YkCIQVIbOVQHFnCe7Sh4imfs0UyMtEX6QwxVIZyd0tGSzsWwClJpxUOOZP3/GhVs
q9cfOyuMh543B9xP4D4LnY9/uHA9SaNYi6gVPzXMLyZxPyhMOqY3oiPwXiJTrIK4
iMaJ0DHhmR7DYDcT4gag56pMH0+VcItZVWq//TtM2mOR2TZpVixMalSxTnqlgYBK
TKxnORqmCuHR81zeAzLSeoa/9Aj3o9wiGhJQBrqfm0l3PvZXf7ufG9gbi9BnORrt
8521bSFBGFZRQEeGyy1jTlkK58IyhiuRLqDByqYAdWxhfjhv75KvIBbs0BquAlhO
qHn7ryojUm3mRKdftHR4sauALwQvyCE3Tb4H8sNgjcr7mEuPyjUq0WF2T3vqdDzR
Vj9ODMRpF+7uKpFq7ML/l/CpYiVVz2zZt2ATGCqq1Bzhfd4VPy1NuvY9b/GaWMpC
alqUzxV5T2NB9ca7w+5mBkjSk6GoShYKaB3npy5sS6NnttaFeg0fXNMMBBlX+UN9
4P/hUpEtINT4ckxXAG0cCT01NyA4O362PK0/r+rXPMfcBgYv6mJLZp624clfGXA8
MfjsAZyXEtdHSkoshFEEUr90S1dReScH82eXBt+/cxMVC5P6tg2fX4SZxKznEgzD
RWuGXZpaYi65KC4YdnJVgmLdQ8W9SxX2hX4XYzOYnhelpl0hq9JLzwdVDfw274+A
mPBViIxAJnhuRNolMLPKEz823shegaghqoTjD4lo+DLQOsZgkyFtlyNtRXWrSarz
iqxqo96E7CCf/zqSQ9I4kkDFXyZ7bpwqzqe1RYYehdbOkybXuKKzczhDjDVUCxIl
HiJOymg9c7UNkMx2oKz8GD2aD+RhjO6Fo1W7didPxz/iVLg3EK+w8mbCX4x6s/2/
vzB2yukg8hapOUQ/NSihTLLBDjiCYGwwMcaJttIGDxlbUbJqXSpk1fEavKSzc4L2
hvCZPXCh6ptRDmoEHxpFtLk9dEM8+41jDpXleJlAcnRgult9phZz9QMOO/JUO+to
B1hy6AiykiC8iw+UHdl4n7ex9W9+Ew1aYFab+vqxLduE0yfAokhV+0AIJfzT7pC7
Q8XcWHJOFuDaLhWagrBOMQF/pS7dqTOyJ+0/HoMxiJVaik4v8lB/FWD6l5+O0G69
5htzILoslVYp0Xqxfxmzyj3Ga7sPRdRDEYbxK+kAN8q+1RHqg/77ImM+l1EjsQNN
LWkd0XJ6EY8dQ6k5o0/4PzSo6DKxbr9LHIB3BytciW1ZwjE96fvnpw9Rgj8oOgG/
9QPC+Fu3MsEd81ONPSj4NwNExUs7/kAGkUK58sgXmBFelEJlklL1fUdYsaJK6Lh6
Z+b908wPRSTTKVmc0Cyu78LUgMBV9kTBw3TB4o94/qbc32pycZQVrQM77T3CG9zJ
o1uEnLP1GvEhNuo8LLphszJsaeSOLsNvj8TUynRdST/Wp7TCliq3GRJ1Qwv/cf6o
/lsSmfK+9tyvczbobhRXwN8Hq/IcxPJakP3zkzFae6gcrQPbXf9w2VcOIlAwsnLr
GzKUPPaQqzqRkRwzho/74Hpa2bPHiLoEocWKXrSvlTQW5mabPXknrZ0GD53ms9BR
YJxmp7VHSP/oa8AbalCK6rxxkvQMTIchAfV2vNhjQy7YcI9OLmGafFu7jqDfTI8+
iZ/l1CfjGBQR2eEsLD7TQfPb0ycuW723Q1Fsg5Gm1WPvdyM/ZE4L0Vo3AgBHfUHC
2yuPtfhr0kvmiGJZc0ZasVceQBIDs1bCsm8f19iVTp91ELxBdo1SgokS1YLeZnRi
mrS/X7heWTAhG5c87iYa6PL+H8TU+utWpIgAfn1IF65hzd+JRCO3FenVJD/k7Vgm
JO1eClaX/gryIYHSc0EbL4ITOyIkJVoDUPXDM1YTkiWIUHyMLA/vGffLuLurYNur
Aa7WBp4TTGl4lmqZbAdICGwpZg7n/36dmNnDTZpPKs185ZvrS0F+pceKoEYIkBcL
mLG/BYIP4BSuKZykDmiB1KWte/ipgeqdCTJu+J2lNpFjRqFQhaoZyA2IpugeiwUe
Ojj5Gt/OLe4ajRfXJwYG/N6YRjYmQrgJErUgHOgQPWIv2JDtqbRxxF8gsJqEurFw
RB11lMAfBKNbfgD84SXIGZzZyyMMEpVEuXZdauIENLl/VS0gNND7ycQ/b+n2L+Yn
hPU0cfDUMy5tCAGR7oIajojmEsBzKybld+nwGneSQX4oAgcEZD6T+aWoid2zf225
weSNWrLiLndz7g9N7G7tHC1gthXTFPCkXDxKxyashJnuTK24Uwqh+5Ci7iJETicw
AvTAcyRL8Rl3rm1N81NIiwjvmFI9RYYhuGIz3Ik8OQ7BdrHyNX2EWF0x0BdQLYZ+
85tgSTYmuENVUoBd72dPuhHCVrZl08vky9L07e0Q+Vol7KWOKXtnrRO0CoVm8Q86
`protect END_PROTECTED
