`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yck8AqMLb/wDLxS4BlGSKlLAbgjtGytWOdR/LeRlGH8nd4HFox5mWcN8PpCEL5A5
dwSuO2ZgNzCsq66FWcR6di7fFFoLU7hOd0LnA+l6xzHnstOLXJAx7353mSFLm6DP
qqieYWwjy0uBsAHzNFNgftM3joAlfw+ScbKWi+4z8nwN1/n9CL/XCI8qxfgyySAd
OMhL6A1zVVjcZuuoodSwZ6iLy4+VrY8QZelVmn4oCwN58uTgkMOtVZL1QtwsIn9n
yRmNLcwWnbQ2GXsq+lQLBAVf5k3UI3buUMHCMPfat3HRUiLo4cQGkscURKJppEA/
KZo9Ur0MsODkuDJ/E/tb++D98K3FoAYlO9/GYdF0geFzIL1+7sAQU0ax3Q6h2uL5
V457a+jsumOKmM76yRBY+wx7rzaWjg75u2nUCB1K9uOM2Q78A/hwO13NGdfMlCS8
iZyPP6L0J41roocSykYiTIsk7O9wWVsMiXqs5D73FvF2XPzblwioLjCtFtAwuR+u
XG0MDj9ZdmqwrMYKAD82b2jRR1CmFlr6/QOxt98bO5ZzBxs5+6mLQQQVkdy+vPtO
PdEgJiFAlj1jpxspxRLsgeFmXb44Ueprha7pQHDaJTjLySzDPXzE8KrK+6pU1Ezf
Hm+NQRgwvsmKsDJFr5kbzRZ4bdnQ5LmQAn6RT9Z1BrQ4vUSMF7aCzQNZXRXKwNIP
U/jdPRIuP+WYXFGk94CF1sajWvD7KWCm0lDUaHVPNB00jjuGZAbX+woaB/2q/7Bn
gd4NZ6eeagqOxd6UOQ8ckjlTeSjXL5oYBjlXTjg7BaH0gQvmcjGlJbuObgXxsc52
i/v+KxPg15bBP2vymMU1pkXBImvAt0hKAhicMg6F/NuK0/8EvvPNhGUAeoMxeD3P
HwDhM8nDfNBdjqy60ztClrFHIAc9luV5vtcHGrvnyH0Zu1GDaOw9NBqh2Jibbvkl
Jwki6P4Q/dcGLxn4iu2DdA==
`protect END_PROTECTED
