`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+jnf2DsznPSL8m8ODkAbYEGzgZtf/szkls8KF6NFDurQtqkw87L3Z5JT2FLiqaSz
/GB1Ulg8GHOHD8Kg25FPbS+wZ54RWGNEpzJHzAntQPTM9y/1MnBDH7Djv13lKkm+
JP3iTHtTuRC/Al4/aswbclvL2IVGBzMyfuL/C/5LOCPABTfgFt9jOvyxqKVvLpRY
rTKYID3CkrZDD71ocYRWtz4QHrRcSI4ZpPjiOiSheYFYAGfbX7UPalfwN+lRZJd2
Kt3PAKX7HTP9TVq9z1Mag4qLkf8WER5UNuiLDU0E0vnZQs9HGVBOvaqdyFOy7Nw5
wbjM1fUdMC6h2d4NGHpg6kWqS1C+fS76l6qM8QHPxHOmPwWL/tz+KiEJQfQ1KWpH
GXx1u2q3LBsWpRLD/8rILzRrSvwJ/DuJxh/ZC9h9PTDPmHVRKiA8qdJa96g9ygNw
64DaEmfJ9Rq7x9A+ZHahY6dCipKR3A5hqsp/hEq17Iy/gfjO2udmwTTb38YTUq9V
WTWMYda4uDvVECOd3NfV8zDB6dgRGuFYW8OS0SvG/34lXswB9JRmm+WxLavzhFiV
B6NlUJD22EXZYY9Bxi9dJWOyugFhuysbwRq1VZYWqZq0zE41lKvE+KaDbPU0HTP1
fRB1sSDOGcgPOfQTOrwB/YXldTBveoboqFzJbnjAz7gMwXT5RgABykT8alqDFpuG
rndjqvBwWi2mQjsVOPqS/6GfwRShakXKJXjmwLGhhiRiVSAIydbg2KvQnaMRuy/J
DATTrjbbwiZYftGut8yLefHWs1ORU9rG72C3rXHyg7MQUmaSZaFve7vyQbNVQwtg
zDCSkvME1HwmhoRNNdz/giz11r70ji7i4xC/vTGEgaHkA8Gie6K+D1Mmgt5avE2z
I7gvApdKmtozxCGe5dKOWyj+tkUZhqk5KE2wSAaBYV9kxMr2B7BETD2nOTuKpQt0
ZdyvuiS2OhnevgztGGM3qb+zRwyTU/UPBWZT+Wm1znUNB8O+aJixrmOVz0gGUuuT
NWcFIIxwwFITwKhskyNrGChBwzLpmo2SOHGOC0F8Ec3EltnjevGYdNU+NZXt5KFT
ex+OcUTAv9aKGXKHdQE0xT10SZZOgqGYngQ5yQD5tyns4eoSz3hjUiP4RjFhpS89
SZNt6e1M01EPCXJZ6uOujoYGglqoQr5iO3mCDo/NwusWddLg9rW2+RJpo+LROJWy
tqLAiMAUVsb6Hq1fQEsa7Cf/Cii+roDoe62sEwSawXBeqQQwxXEY/fIECqHm0YKD
cRZbV5A7UJ/V3rV7mxAaBV7uvdxo5IcYZ+GNz+GYiN0fH/RiiKpXmX3AYbd+JIPW
DCHlILKPeIavw0j8z88/LYwDRWO+jgpSudlqZkro4klWSF6n6Y6AtauBxuVFeXiX
s/XfEd4y9XaFnl0dj8MHojvKTYnVuq4a6HZhgUdEEWtqv6btYO9d5cQ1VJj5VpJb
1/l9tiTKNoRUJ+0NxnsEbLgluk1gKQmq166ii9fAlTnRJOIe1wRvWQrbehx/Roms
T28xP4Lrd3nWHb/A8sfkzdm6CG2/SYBVT2EtCoopzkwZbXGQZ9n9yQVjYeRqPfc0
cogKWG1I88ME00g4gDNLaMDlnIpeZxjeiVEnNNPrXKH1hayMc0dDRGlTm0WxuTOx
QIJXN7ARs7YpeSSnj7rB3VlZp6T3Va9ge+2phS86JctqTEddAo2PBcxx6imoEZ7R
jfA+dEe1pz3CMTQ8gO7gaGAh/61nCaKoQx3IW6YEc/P038KWw2Q5Qnk419/yJBUM
uZHB/UD0G8Wk9iK3GMiITn7gp7XgnSUdtIHZHaL9w55a1P3yQQr6qzBgHXkJVV63
ngMftdTJU81KkQBqvKDUmMpBOtGto6YQ6FdmSupNghOqLR8g8dd1evPNIa8Hfmgw
s+K4bsVi32YzzhiOrlNJNVyVsyOfYrWRbBVA1hLai2GE0xInkgGCpCxdsk6v0D2B
DY63Sp0fyYRoAvmk22WCB+P0LNl7pcQuyz90WCFTXC/IAuZrF5gw8EUCeyWHHHcv
WOQKKzJaxHOggwGAMhy9vg==
`protect END_PROTECTED
