`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qVVF6D+Bd3EygyCQ4OeHb6SlWAh5c/gbpafqSb3B5iHgA5YYgHaKX9wIeDM4W/k0
P798vUgFO723vc9OO0+F9OleXDCm1VgqIzmFWcJkxT1vgD2YTOszcjEkwtqDML9u
BN6+1KqxAr/DKY5TWpXUmRKTfCoS3oSNvUBN+LEK5g3etRX2b6pUt7kb0lVpoJ0L
rIQIY+dzU+R4j19HYUtfXD0gvdKd1LEdKnWUkyZFhDPN9NxoLJmf9REMgOOqdyII
xXPT6gctmvJsLuoqA59OHOJaoc338JDNB979U9y+HN/r0tAshDa1+0zjt/tEJS6O
ZgervLzrizFZEKkKt8XtW4Fm5vTcR6RdEalFbeMH6e8O/mA9X5Djx+nt7/HAqjUN
`protect END_PROTECTED
