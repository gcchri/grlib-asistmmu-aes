`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pmDTVqQHLDMu6VUrIeNf5fKnSWZbRxVGDw+ew4/2ggSMP1ltqT2d0YfMaKZjexaM
jl1CJ9h/S+HNq1YMY3OQpllqhWyCk4ozm1h53Ce4PYdwk9c8Q0dYbxtTbo2yXLU5
oFf9WeJs3XF0Sl5lkPxcBuz2WFSUrNVn7tVuvW6/4hpZfUM+wziA+XXpBH4aM6yo
whTGv5bMFxpsGfrttXvupl66FZwXosF4Uy1ms5igeUFolQcATTheS5Jgu2pso7iu
X89h61s9bnZiqoCew14TM/mku2BUEPdOxWKh4QG/VTGHTFJFfXux4fV4ZwmcjhQy
Um5avwexELjkxFjcAzyb/Us0I9fDKYHE2BY9+6RvW/CSHp1iyQ+XuacTSYJhzmjk
l7HmgTBy0RPl8h0z15CP27jkxF/uD0VLD2xsPfnDVCTwad9anPDW/j70l9j80xMR
X2p/n0SHUojg8TBtmPodkoGcwWKxMgsJFnZ0uahqKVP4JDzQY9hIpgNdImv6HHeA
iO9bufCDt2vtVHFs21V1fHdIntWitokU1aq5E3wk1pWS/v6AqPU/aPICQu9luY+B
iUOpe6hEZBkC406O4R+snE7G1PDcT/b3c/+2htdudJ0GFmDxfSSLxvIPEDOkrKoY
zREaW9CBfrgWc4GRQcKbVYHwTRWaVK71wnIdXhzYiW8=
`protect END_PROTECTED
