`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HTo4DlP0MOTFe4ildCy1hvJHRFWnrpErzKKf0Q+hjM07jPmUb1AgxCz/wXoo+H0w
BT5sa43lnAOMJzA9xCvxBpAE0i9qtsK+0g4hMyKBi1H8Axhsygl8LKLXjTllMdFm
1/58IhlLfPfDSStDjRWuQONNeEwUmHRxo9uq/qR7rc24dXLGRzDioHOZAkdU03lV
G4gBkzmY+sjEYZWhNOEjUYX/tuyWdzzvWmvPApACy3vKoUE5D0boCyNTcmQ/hPPA
JLJcPQzLieJfW4bOrPRZkbnFH/TasWZDm0Gvgme1ZMBO4dq61vRMhrv9aVvOvGOW
OFrYpFloM80UGtWHR4ZEdmxIIcdon7w5I9Ot7YoW24aWfjWeXud6oolZlVTgic2X
RuTSzeypHg1WEBdf/raMYDYO/77HZsNLeiRf1dF1CZbZf6xYFmZnKXg7vq75jbd6
a6p21+twHWYuR58QyHi13rmbl/SwDWMBesFvuyaTsBwg1ivJUqPzskrUS2a1Cw9M
qemZsD+s48/O/PM37DYMtnVLaEea0XhmXFn6RRtbZVvtRE7E+wSAKMTaPNm5LLaA
vkS08FmFZClWDn9C2neUi0LkFDOC/pS3kfuzcVcuZgR3SM5lyYbTAZrnpmfabVSm
ohLSIAkcgMllPb0aaMoysx+IXEz194a1L4AqJIeMOpzs9C6IZFMyKdjgV0mLDSZq
ltc/xZjJ+Br+WPCeIR0+97fvjLbVSwZqtbHvGvVFYltJsUlAgCxCdtN+FkMoX20i
9XGZ5hUvyWtHXOyvTb/ZF+X+P65OFGHqr7/1Hiun4BpO5hxApCFdSNtKPAa8zSqm
ySHKaL0IWCWiqHH6VxSC0A==
`protect END_PROTECTED
