`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1c4/MdfjUYTZ6dJ19cvJXp2cW7JkXYX4faJDTmGQNGgAlp0wFeYAHfeLwffoZYSA
rzsxEpIOcut8KGkxoAH7GXWVizcPoy471b7pK1FMhrmF6EBlUMp+wQo8lguzPMR1
KzqK/OoXXrUuXQsNVWkvn0G7KR5//h9DPRR98paFhyOUZIWhYRRMqEcm9Fe1o6xF
9gp4pveXzDIQZn1rPLQDvB2fKFTerZZGvoqNkmt+RSQgQGrZVrXczgHwHaUAgONj
dZmr6fuwsCg0mZ6Ua3c0oWi8Bsq2ZCMXL5e5OERdjB43YYA6EBa+FKI9AbpomxTm
XGnjDdnPTgjXwMsMbFPuPzgQa7AV4bRKW3soxCq1URj1+BvpEPYAdOWsEOTwTZHD
z1oTiZuAqmpjB5/pfOEQdOQG6gbQFAdtKanbma0MTmyOIATv1ZmW0JLqOJG2s4yg
4QbyAyjAXoH/cQ0CzN4VAtZ1JQOn+ocCFkUJCzf2u4G1kJS+GDZcg511F4pssf0e
hUYLOYhFA+05Pb3stojl57nXJAFYtXRlf+8Qn4r8IHEYlw1CwY2ywU58czOpMp/V
T8Q2UC2ExHSneaigjtCU8WbCnlWo4XzTDeTYY1ZRGmDNw2HJWxnQmwmHYFtDYowJ
tW3uvt/ZF9iarOrdMJu6Ll/TqyZrDPjyw8EawrEDrSC0lTmaEGKxcb+1nlGpnI41
fbaTi/7SddF1g2WI4S9LHCFxFDjSavNTdpwbnnwOsi/SKx1aLB2Qh2LFqLI7jj1g
HrMYiIoFIk38LAnYeyZZNmOGryzEvzJ9eBg10saWJeoHOXv9fX4JhUyDOzFOAJLf
oRFyZ0Nuh1NIdPWuBLNlKgwrdUye+yOXs+N0Wpr/PyG9QEhdmsjYyYItLYkKwJTf
Ujf7w1BZ0KC9aj/7gl/T6xFLrUTFgKJaiZeXoYOBOrGb5gsmOWVOT0ZeselHPVjb
g+mGuR5LDM7QTUNI9l282ZiSTseXpmakPiEP3wNbTRx9WykuTZ9SdNgpGr1iTGKE
gmHKHjknliixe8zWC9fqArGXdhLbeugdOPuRfqzJTzORDJ2WYPgkGmRjHhnsr9ab
VUFRUeciwf2BDCYwzLT3naXf5rctai0zc0sI5gcQSK5JiL66jdd41nj/7qVS3bKP
EE3+VAgcLpXBfMO2OYM3Ed85Y0BCT+B8lRrx2eVNFmnZipnorm0lzyVlrNAj8Hw+
6LOOmRtG/ataQf6w95hz7jK3tGO8DJ9OP41jePV6jKJz8IAATRMYm1VDDbFeJVrs
rc4AQIK+DtMArjmb7AvQDOXJZiuMZHudAmfRWHB464uYug7wqi1q8hJLrjYuEJ3a
xK0b1iUQSn0c8mOBbcKfSuWW6q0tf5MGQtsl/qQdRVFtc+NcDQxlrKR35kQKaHxZ
CxJe1Yw9ta8CZ8Yky1IzRrpW5doHGUSeNRc4bSJAfzNBId3YrBjCeT8gDThuDmr3
wG6UnoRvJzXMXPqCOzGlCTzQGJmNIb2BNtHDAMk7g2pT+Wzn/lmq8vR4vxTI67I3
dipdHP06A7IefcZftRC3lmQ4L04tGhpMF5euQqUdu9TV2AkNwLtGgnuKpSUtTGbY
4iHsIk+2a7eRSsYknJDfsZfHxU3D1ExOQpe5NUyM0LPwIFOD4nZEClWctUKg1py9
Gm1DmxQSgLWDd6LJZUQB1tDGdEd51SlD5DRmNz3ciWMSGHUNlQuwnUai8NoMt+wH
ECdfoJv/3ja4GEQSh6FouFosRscGEe6dSaO0W7kO2916kbdHxpEp2FVz7J5zddPR
7xP0vN4cysjbcVEBFjgrutT7rvXR/JEojgB/58Uio0wMgoLXw66SFJTtxfU6YwwP
VkorpghXj/jkASJHezg1f2+AiW/bM1JUZ5Zw+QqPcIi87h1zJkQzv712oJ6iLanm
DrGKlkx7vvUbv1U1lVKXNZIUTKhO1f0VM4MOECbThtdMjwv/OIlpD4BccVLWd+55
Ju+UAj1oXGAUi+rdfxr11ypVfY5hIxnipS7IYhzP42XbEz/TgQpACwMnAIUA9Fzx
o8hCgkEspNmU4kVvXQVtWoAwxwKZOme5Yip3nJuRgSM94IWtdAUKgf48mN/QOphK
cVK6ubRi6cX+AOLo/8Hq7KMzobXplQ/m2wiA8lDpn2uoY7pndJFtRFTe61VKq6kK
/a3Q62albkmcVDzYqX+Uwy8DdKVE9aBtk+0EM74D2bb3VxggD5GvUXo9ApEQeFxw
e77iy0i01Uu9xP00+i7g8GZgmKx5gNcmbTL8unkCbKytN8pKJYHn1q2mEKryhWd+
x9pQwqZ6zIKWzSsExEEEffk0XKDY8UDnBW6GAFFrzF1o8TO+l5tAJqgjudKiHiRN
gEAigYT4plqHfCuKy07xoGD4GbTRSmnOgwR/ZNzljdh96sfz0fFd8O65EBNyvfE9
KF+8mc41bL5paU5DGZMireh8pWOF1r+7XxstYcnrvW3orKZvVR2CGM9szDbwNlbP
urMGbe6u2XQTH3Wwlvu7lQvaGmdaZ98fGgNbFQZYJIZ28aPVmXsfEtkXYKghsyld
K3GoPYFwrQge0CNEPXVg6fxnbCN/r72g6pgBR0w67GcMI7Lomn3OOsM+GXs9t6x+
+jGck1DzONpgh6uio7B7EPSIfYWo44FGcegV1szltdWWx2T6jmTLBd2B8jhUkTaS
x87Zxydp6mmt1FDQ/5YrNiRfHuA0AGm7IISb3ZO6RfxETFVIOm66A4JisDi6Qgu7
WxAEOkrS5DINRx+OVtB92IXH+qC0v6F4uUyWlQaOWIeazD163ORJd5Deqe+gk5HD
gCSHSOhF3vb7lwVn2AYN6Ct0b51VvUA/rJdgqfJ/6vc5aNBEwCUFj+B1xOi3tFHN
nxmL/n/jXLfejwk4gKci3alAWzuhjo3y92H7z9vWhhbH53aM/Es4Xo+Ho2PzV9+l
Eb5ONUqYgg/0HJ8nP5dCWhJHEVhUWwy15OtTby9jA0xZTYfQpAgz5/RRaq/hFwWD
WGhTaHNpUaCUu6tIs7DisPOgAg+MkQO6lKNnLIl0O5C9lY0Mm5e8KNQ6hBW0fET4
7G8xBQzNvQXntR72EZOgoUYE349MyBavRfK+SC2JQXOxj/A+Dq0Wr7KqrhwBgKHd
dRcMwjQxs9gSJFwwdlpRR7FZgVUjL/9kn0jnlW1bel3bAxc6/IcEQNDSPVgPOhu1
oZKlHl67+p4nDtWe/kFJObAFm9UF71g7TdnxTpD64ZqNJUUYUzAjzmgYzJsVjI45
ktR13d+6RI8rfHrvHafxgaSpvd8UUP1rjvAXcFjpDdIR4qnomtUtMLp4z+sSC90R
NB5IX3J4ZxxdQkInLRuzHsUX5mp3Vd1PgeD37y5oM7GDxKIsHZTfpfvhniazPAp2
trMZ0ZywnnnCYLuEjd4JmsvzYuQiXRcSy2Kil3myEjzdrpkm57wHk3c1R5Lkb3ak
lZFC+b/S0VgUfTbJ5r0jks95CYvyzsdSUyGf6tLo8CiVaBc5Wz0XyF/lmiiaopWb
ffKw4GBfoOlNom48g9yL7N6wvFr/kejxyuyerDHC2TTxM6Gvn14/YWh365b7P5tU
zrVuuytMdw05XadOMDK9wo1nSiyww1SZBeJggB8ejSAeTDCleVyoNlUaC3+6ZzG6
3YTteLFw2kESua1Q5anTd0+ZkpHBnMDnxqCXGqEUUnyDuMjRBeHilO6gwLYV4+pa
JZ25eJx4AwStHW13K2MoVR+Mwmb8XdeLVfdsOmQPqLClGN4JPgdIGVk1w5+RBY23
srS+GxN5zUT1qfpc6HNLmO5xFlmWSHmcP0MgYY7KzZAq7gR0pb/DW31q8okY/frm
Ov4w41asRtQSyR3EgCHMscTpEzz1K3TzmWngsBIrbbcSWKPgzn5Qc8SkVD0EsyhI
u0qQ36W9+94+Xqhqx0qf1NrwGqbxZ1FTr7gN/j9CGv3vH3aJtKZKIxk0nAVAdPyr
H0sSSDfAsL+8EU2BclLBZRM8pofQ58TJ9Fo4+f9R+8vXXJ+1ZVEhMMTnVHKm6iOv
IgTBz1hoJOBv6jq5d02qsBRsG7PbVy6PuZdOmntLyXTGOOU4OO7DrOheThukTmGG
EpHAB9qjpy8PR+OxjzAIq+YfB30MxiY/YM5Ar3qiWxHUMUIvm+bvHdhaj4ATZRSL
Fnfs9ywYks3Y5upchLySWgKa+PGpZfx9eoqe5cLhqIOf+WugxfWt937e7sidGhy6
Tu3ScV68MNrRCRIOyXAnuPkwAMVLMGj3TtyryG1KDIJNoHoXsIGskZNpc2wPXSgO
Vjr6yl/ezpy+tbOm4W+euKvnaXHwE3w2FpX/3bpVZoeggyed4ZT1BJAHg2XtmB3d
yjeq9Pt9HtqX/sifqoOfejMlmZZeoFnjC1fX8zS5no416ROA0tkss7r3+PDAVW1t
QE5P/mOlAq66OE3FrXARC9vZZQInf+Pcb3BnGZTuYdIfu5XpKEApDro1XIyGAotJ
aVJ1xMJDB92ExmwX2A+7j6RLhZGqkfwuytIYMxRJNUjUA/598Hw46ll+JNy+nJju
32N7fepjjL2t6geCiZmajIJ8hAgh5cZDb++PEPw+aLwXkGrK6Md33pZvEp+Muldf
/CpM2CVjdnqZE3hcgE5uZTPNTXfShQ0AbrMHogi7Ek7HzYGUqrFh57RKcOANivO6
XCP1kkmvdyYKvSXsNNnCtQ==
`protect END_PROTECTED
