`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5R/GqwLFlNYvGQd66z9gAyTl8GHuaXJQ5gp2wrWgTGJ0kmFy05RhpBwI9ZDP442U
bf5rqFzvl822x9R+7ieMG+1SfpiocJN8cCehgM6VC3kgVZAfs1SY72vY/rpdTxg8
Upb4+fwAxHPV9q8ZOmtYyFGr6pqyMlZh7goXf3qtkw1ee6mSvEHJqo3KTcHCeFMD
55xZtQwcBFb6k+dmjx54n3J0J2t3STNaK0m3B60HQ1vQ7P7z9BUQsXG1fHPJk5vt
sGseoI9wT3w2cf3nb4rGWIF0L/fd38xxVhpnqQXbkL5tAmeEBbN9qey+Fo5KNUCI
05vRi9FRHg4a2vRi6oOAoSDLIvF5HPlSKo54vY3Vj5siw40f7YmGaewR1Y9PKWRe
u5T6nQu0r4mf/LRKkbpSVz3yDR6iTI0qj5GVvwpr89jjqT0ckfbGXPW/ylrtF7Vb
h5+FU0vUS1Hi6LcGxQ9d5s8Pnr26Gvb8D2HHFdpl+PqHe4QTFaduXoPvjGtyiA/t
n4fDBuLJNCBoNM/cyCRragXEDjviV+2/GFawDW5skxpuDzHIVo6XuCYu+oIMtkYW
pHkjol14HGp/5BfT2vXi7E1H8KY4eHZGTNPE3pv7zeE=
`protect END_PROTECTED
