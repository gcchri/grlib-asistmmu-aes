`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DTxcMGCBkn2LCm6VtCK+faHa/yjcQkGa0mstxNBL4SIHlLy1nTcKMqVwSqprZ1y2
0HSivbNBM/smqWUxFT2YPBYnwPSZwKwHKhJzfYcuctCx/M/xMtObzqA+kVrqi2ZR
eZwC3wKLPZWnrg7zMRLv9DQwbQUeymiWH3P2Xcqs/PeKD7vkoDjD/uwqxzMqRiHL
1+QTP2kiMDAN/STfVQEJ05yMDBM7lbwKlROIguMdkd2solt6Vv3E4cm+q13rmAym
QKe9fBdpccP1Wi8U/bHzeGdorIBBcyHelvi/NjEUtsjoBy66614SrxhlZKdr1C+7
g+mVZZr2gyzK4e7+HcPywDf4wzgdFix9FeYkUYcGo3bf1EbZnl3jupjaG7cxqmUj
EdvF+EhWogeLs4GXNkSQtBb40M2xI+x7VXlJfCjrdEU=
`protect END_PROTECTED
