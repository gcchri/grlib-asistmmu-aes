`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KacVsarMsD16jvfH2dd8YDqgnFNfdma5VQ9BYNNUdkUnlSjxD+t0LZZta14M9l+T
35AqM6PHmgzeodrYujkr+ro26VYkikhKdJKABc9ceiKLMEKJWTN5wS8u7I9MpLce
mrWJa9VX9z2j8TowlRr+ocGweV4YijtgmG1Llubq0qzsARdRvdJgyKrNq46KBScb
NNozudUos5plXhvZ8rBcAYXAFt+9gVQiGQwTA37wB2cHSqHocJ1r/VDo5V0U+760
jsrSho390YSveZOecvx9LSabwhg1C0QJLo2ADZ/6mDOfk3T96IcKodSHTCBxNFV/
2aQpDq+B/lpCYltahdpOYsHS7sDulK25KHAZwWLGXPl+xWdlGUPRYsnOnUnYxAeP
yTW7FPCt0hwNXiIk4ge598ht/npbGdln04P3nnkUKK9emyqHzTLB599ABeexCURV
tsumUPSqwhIbcGr4BuIjxtQlJ7yz/UqqfgzWGN/UQV8GZkG1mI9LvVpXObO2udK5
C3ztBQTrnaLe1JJ7LX7TpcyjOdbbYQdhpOpNl99/gVBih2q58hJh4BH8bGby8GwR
0lihR6hn4fkPGGC2uNjyqNCH1IvlwP6+AC90ukPZPr52eNDd0yhMTdnfCEPnTVCw
DCMDlmHmNIpncQWxqnvDbfuoEAG8HJRwhL6eHNNA7hdeNrqeDuPXfkk789OaBu93
Oj0I2d7CguYOWiDxDzR8IH8rSr+tY6RT49CK8wBIKXNlcoIc6kFotVYwAErvDEY0
sjxOpVzP7Ldeq07A8f/qOFJoW/NMR7K5YCp4gR1asDUQkc4oXXJquXFcKL6puO3w
9WcC+K7dt3Zfo0HOXdETI6EGoZYBWDyMf2BUapZTK6R1RDouIUEG3zKx3wkdDsdk
pBjCShV36fXbyDsxw8EiIHrxN9dWyjusHb142yBUUwouUg2hQy9KPgWgRZt/5pEY
HrDIT/rkgs07KgJCQk19zp7urdHhRocyLMJ28m7aZv2vNlc4QGXe4GeHwMruD5lR
2SSoAYWk9Y6hYmjosjs7XXovx/AkiVMj61Qck5XlG7wr7HUlsZcL6k1vXH+XbzTF
biLYv3L0+MjwLqECWMUzjb9iCmlwU/JOL5iqrhaDJTtM947bx2pBE0m+AFFg8kc0
E/aeWNSB4ZTzeUj4lseVGBUvBmEqZITnvAf3Kpt836vijyxXHq0RmTjgYJ+h9uW2
FSjvTY3yPjCrxHpP7rFYTogWe4X+nuiu77rpOVoqrdxPQHop32QRuVLxyK37yQpJ
WLgxs8TqRyKEqFMKYjP+05v9mreBC2bIwHvEsO0qtzqtvPad4kNlXHdpV1rrORhD
vf5qRjJ2qjVgGNzYR1/9iiJ/lV2zKyVUsM/rmm8TenYQ3iPaIzn5nAt7bwFZgmXu
sphr8d8QoF5e3kfsr+ouaWi3rSB/u3vzDD1ZtQyf4v0A+xfz4tcGS2umGFYKGS4B
ku0k0w8Ij2qRhVPyZzZUpO1igUhJgwAKsLRUug9w8UGy1VPetWR4rNaY7PQTDnQZ
cP4iSx6L4QWQXkb7oAJrNK3V/4KhUlf7itx7Y2TF/6CIkzVoJV7jatprXINdjZzN
YwqOPPaYfwEZ57eDm89NVwfK1RcTvQ7KcA6QwPTJe/peXjkRhFSRaUN0+9g6Cytj
DJm3Oa4JKYX3e9hhjkB2eZPNNXpBfatKJg6sYIlpR4kpynIJ57Jw/azWLuU69Szb
JQ9oYlHBVtyymGnOGDRlCtC3Q7JaO1IMSarvVlLXT4yzGVIDkNIqlSYMeUEflCLB
cZPp2ii93t2m81jPZ3y301TXrJjc6GMKPhUM5x0sNBY4lAnVdtMN4+KV3cIs3yoB
iYS1HTcAfpNqUk3t5MseHg5Ra5QJLCOP/zr31hYKmPRFRB87VDNXXM/rqQKpdkjC
5J55oHF28Y0Nq8LF9wn+Ic2Uk6f6I7Es9GkpEwDnTkLiXQfe9qKwL2Bzd56YFomB
sYS/IYrt0xXeJ1xLpeNI+29qpiMLeNeEZMANvZ1t/mUY55zCCisEyg0C7WOIOjuC
bhPrGfXhbnxCES9BONDG5KR2rSBoRl+2m7DKTKb/ZhnlG3LhIx+V+M+qzphxCozY
o7HtkIIC7o+sk4xnI5UAvgjOa4aYSgKuG6ioIGMle0LYKWsLMXSXaNLbA5K/EPtn
nk2R1zIBl8xG3w3rJK4x8ixusWaJK3MLUD0B/I7+TABgK3bg/5ue2oZHd8lA+jYL
xhJUQfzrBveBklWjhlDMGdbpRiM/I/Kz9J0VOrhf75vT+euZuPY2dyWSWPQBXUTo
eFwSIYw0sl625Gg0MzCjZzrU5uBFqcMFqMGyNXGURWcK6yHLARSM0W7OnsczzseM
EA5oVx/XhrJIsca2ScCGThXfpF3/CnwMUHeQnbvNP3Brm0uwp3ulEbadXZhkQaFG
fgXIobCSYuJ16GLt1Sk3BMNrhmk6ewIDlsaimmFChBg5/VopoKQ3t9z940yXrK6V
2XEetaaofMHs/icTBpUGNxhTwRPjrGVAP6chr9UxemdcYhhSHBtSJE3vE2xoPoKa
YPU4GTMuX0ZpGBvUehbigTs9arfipskavwceIVORSiO8EiG03oqo1pyPazjMfC/x
pER7/Z0ysjIQ7KUuf0T+wGC7IPI/vt/NiwLCjcrQJ+QQ/jEpMoslBcpyqnuaoPQR
jReoKWLn7ODd410roCSDEmekcOUL/CO709cPLrUbsOpGOWmOD0daqaGT45MyS6BH
Cr9wQSFeUG4Tvq8t2cKZMd/J7Ju6SPeFOI1s2dLdSrWLgR+DyrdpghZg+xfpcMxd
h7R1MdtxJW6IRGVrj1uqaINh8zIL3yn1lZ2A2t4BVQGYxiRisza0TOykNWDBgZaQ
noXdpQHTad2btfM0/wls1NgJV3e/KrSeMGUE2ETm2vl5M0dA60bA0OX+KDrIZ/7n
6xL/48NoDF0M3OJp4jvCePRo5rjXPE7SijiTozZ1qeZL4gaYvhxblUfLI707GP0y
fvdH1pnC9LrjWWZf63MNPEnzFnLrvJ3lVC3cZFt3svMgY7dfCaMJFvD61/p+f9Lf
TrcKe4M+hgEOvibsq2JaH/NhiF0WxNAH/RqyZ72x9+UTEkyFa38doZzrZs5bbfiD
EeKT1mHhgTl5N/RdL09WS0kv1ehT6z8i35iPq1EhAQTcu0bxcNY8hl12b00O4tZh
yguUvPqMkKY1drke9FW/Yl8lg98u0VLErJK7INL2zV0hkBp4bo2WwYBqcqrUC956
zUETzsljBTlQoJ5Ph+3pdsFpx2wCqDzrApIlU6SLgQAHkuvmhy/Po4RggICg45T9
e3cFye6iEzi0XWojdT5jlv6mvnFq1JBjNiEnwdEmTYQlQHm/0s6PclaL6csXG2Kb
9cJF7s5r8HnL1t1YnSOAPuI750Lz8364+kaQu+3iSmlOIhLciyKSNVSWbxyw+EHs
+S30I07/fjJrdyl07DuuZakWT+qMYVK95m9oDTFBt1VAgu5cpPuwsyhJGRJyP4Ob
e60CCO8HVFCqxLt9291emuQbzhEXCRRNj0xFuIPi4IcCFXjfk8iHyz6J855ks2c1
US+ubELNU0ebm13C0LkaVfx3P/E7zoYOAGtsWCPY9ThiwpRUMMfv1mObApxW3OpA
riUtEgPlQWekdZEjP25FLZycD9GFwuPvhl9NLf6wcXamKPtI0A85jx4zmlUOT6KP
ai9UGjcYOuqOLSs8CHbXK14Y1IeqU49ghrKXF4/83IDZZMv13jf3RSNGHTuVzVBz
gTXzlTyOe17Q04fYo2JK8lDlx57DxPrgQ0HLOPoa/6ldF48pO5xNn51Z9mnPFH5V
mflTC9QWbQuYxnlLohkaNXvB2u4qEZBaBgmn08MkOwP/msTa38TXhinmZFh41Ilg
djVTDYpXBlSmAbN778Mb5oez2uIj8Jg+ejdoCUfOb21PKXYbr7iQ5v8TJy2OLHhE
taOggHa6fnWIUWtVd9HMJI9iAMJ4KMVfcVe++kopG6uUIjctcbOmOq59T9zgFHqd
rccBCj+Ec3GtqoAirJwhnvUmLp047tpnHJsqiYiD7B+5uGWGb/6JFQNHAtCvpqbG
eShc0/DRWDiXNHTj3Qhj0fXXiFPkpktL54oEQ0RgF0qSQTt5iItFwYa4U84qLiBr
KgD3UJVEc1sjv10zdWywR8vYlaDiPJMtCpJdGzQ3AGk62f1wnpGI26eZITqhpxvv
Olgy9QwPLv62HXz5og1X5SJUEY0bSeRCmEcht+n0FEFdEZBLC8Rv8/6O8Qf61r4M
e/rff/t/recZUWzdS7qGizbR61/cSG5gImF4u3wr3tO5bF4efo0jPuKRsKO1LCeC
luWRaXI44MtavFZuMn9qiSKTIONR1kXKcqhYri+pmK+GqtfolOnmVQ1jabNYrXeX
eId8hZvxBhnUPkAaN7XQ0dW5WA471QQobb0wwB9KTSZkPzQ87fbKXTs2z/j2sc+W
kUq7yCb8X/vT5RuwrAL+0LBbAN0HV+18efbW3CmZoR7DdTjuuBu2tv5cCLH+IJXa
dtjwTjD53Nu8mDaTVYZ1hiuTJQbjewL4swB5QtVRFXpfehUXglMf+oGML65843Ei
sYuNNf9XbBJ+vkGGdPtI7kqba9kKJ6upubkKkekuoPyaWaIGIXlZNzWjuCBuR62D
XwG5O42zOBUSLgs6rSRH2Nj7U9M+fPz5bqa4YD5AxPlzpLwi/KW77l0m1v/dXckG
8yhrYVgnGCenTp7QMDni8GPwhMYlsRmeAsmUvYePFZZSL5hWQlvGJ2dO+BZ0X4re
IWqzKY9I2E/nJNKHQ2embb9mZWkcKxGXfAYlJ2i1EBnnLAdrzphh819X5b1VHoBA
nq1lNm0H7wRi6eQbCwKog9GB1jW6I6PPPFNaYaSz03GYgFWAnXkrk26vuAigon89
pjPiZP7gdmyNAGI59lo3CPbEBqQ/jYplUCTXkhM0el6aT9gzQOLOIkBpKUM3175e
EMx3OMUE7DtIEdv/HZPgsCUjY7C4gIF2bEpgiygOdRf2aGxGTDQ+YjAyd2wQ5KHj
XP6aCAWB8RLQJelhtPDLDzosNMW0foj90LH8iDpsPNQpteKcMyCyWuaREJnX5zwT
9hfpIHVbawYkBEWQqcHOqT8FNVfp68FER3tN9eW2HYkpjlTd7QHIpCcCkksuRjr0
JO2my7r+2m5odryGq4v+dBxl4A8PpPEP/0NdEGP39ys4BW/TqFZ7Ha5+2+oxeL7K
/iVyKxVN9KdHJSPS5Y68Ft4GvcKtYpv8W1/jWvwn9hZFysbO67xY+56Ry63r4I6n
Z+NR7N1OA5XrtpkdRKrjoqoBvJtFL8rrpRrky/QZNYrMND8XjI5Z0KB8uArz/dJx
+5UmcUFKEcGMropCEPxaT/HiMnj5MshZ0x779rsw/J83wsU5RbJDwwVNH+f9Uja0
FAfQO3+rkI1n0Vte20k3O7BdY3A7U8AwTLUI+Xjh55uHmaHZDDCFZKnmqeMUldBU
PDTu8ruv2EacXQAF+sg5I34xM7Pn4MHEIm1OQ7olT1iJSEyBNfvhMpfvNGids99d
ho+E9SZIosjhiQShEGAdXxOYEcvW5nAqXvA9PcGgK4xf8oqMsiq31R9AOl43T0Dd
g6XoH/7hEf0bOeyBDDRnb3M1NzIiezEvW3UoCupAKWzc+LcRD0QZIjIjbxkBWdtg
wiuxDI558+uSvAAniw1A+gvO+s72Ua3TvN4G9myMCelGVjucS5c/JL1pAg4+wAwR
GvhpIkEaF0MpedyBawHwm3HIPJX6z9B+HlIB1zMijTzwTy6LVz2inNzVPG2Tc4lV
FXI4kDN/khIcXDYF/b6jx9mQaDrOj//+KFolMyXShlraHWxFDRdFX5C0Eo7JGF7N
QtUNCyZnDgMwcCVzpJ5YOPnW493OgE0h404hikqsVi+pPTGoPjCJJ+BQwgj+/zmW
d5AzsqTmLCuLAtqJpJtZej0up5pU4dQ8gs0e7pVHq/vY158NfSDQOz/mJ/cvHqFB
vGfv5fq+YB2oWE6X0VZUZembU6EPg+FRF2qWbdBBBh1Altc94jhc6NpVHQLhTFQR
j3l2B8pocEfPCs1HNNjjVa3qet2EfwK5LsZAqH7KAKi2ZYExrMM03Ueq7Ps5Di+w
F6yNsoMZgF3HVlCyaHJilipBodrCyWRtCZ2SNTMqTdF8FGIBrqVjBEATiKKS5rOW
3x3GnuB0aILsXeeZbzGlFD3M2+w3H/b8e9nphBId5iERJlPds/PfUQ/QDIfwneqA
eyxmHIJz0KNoSL1C7pJnQ3iA0IOjMKrnZDboOzH4VFef37BzMKW+PHaErAq6+oIr
whNfuFn2VF6pKRBqs8UAcrcR6ApoLf+UZLgzVJn0oGi5sFrxU1R+vOedDQKUrLm6
/MIJjhWZ2Mr18zB8SIw1itS0Fp5WiroVcbRm8t9BtRPZQ2169pJ/dGbXsITk+BcA
qFKcyD7RppwbrQnH/DBBgeH5cdKCukoY2TnTzLfYWHvSdnOa1AHPKUrmUSAAjJnp
9uOnR0XQQ/7PGssaTEbY8a5xRm/oSFA74asF1jkAJ7+PZmZttwS3k8dw8AU9YshI
GL3hm1iqPms9FBb1Rnx0taWVpr+ZbQal4Kh/RpxFdpWmw+o4K8kkFfM4d7Vh3Cjz
v93TIYpy2Yt1pzYJKb12oe6YKfu9G1DsAF22uFH8M/mUiuRy54ouVao2zuutSsao
F2aXi1aWorF9FWhY/qOdmAVj23LNL6yrrLABFR6mDvLKHhfJ21+Jj85XfZIISuPh
e966/qUpK4IHk4MTNKgZd0G5VnVDd65CQqB5WPT8MzUs7qUCfxIL0ENT5t2AvZTk
0ddxt1e0e5AzlWKnPCqJ9LXKUoGTpZFVUQTM0b0ZT1qSWNg2Hw8Vv3q2NynkuEkT
fkwl2rZZWiYOU+0fr42aL8qQXjbdF7kwPmKN4S5e3Wmjli0HebIXRgcvl3Q7fNgg
9oqdAaoziQlzs8QvUwXIH5b2MZzCbjunkrddOoBFw3odyZjLLjDsQaDRSXhhlJfc
GvP7o2+3FRjqbhNoQoEt8scuDd2ZNPUP6Ad7KGrwTphZK4UvrS7j/d70LICCt2wH
2OYXp2zNdoCgWP3zL/uGaHK85rlxXpTv19TVTLHQIoZWwB+iVQW7bQ6gPS8ZxL+W
HZhswVj17GK/khaVOcwa/TKgZgP242ND9JhjdwbsLSqfIRDwkF6XhfH8JyY4iSxU
6nEaEJjgzvzp/upLIUB5IX/7jxGGzLyql7nW3GpwGjICLPJASA9Gbi4xe/6ECVlp
OSUrjm6PMqtx++bwuJ4lgqDzzhTLym73Sy3akKLhXHlHzwr7cT4n5jvLqbV14Aby
KoCUXGAld1+JAU4luhAngghIKEj1PLbzfyqY9GA1ld3/V45co40lLCFf5iUi1yog
Wy4bSccaDToB96QjI4IgQcYu+v5dnst6FXSHURW8DfFLOllj7IhcNVDbv1ywgCom
RempCNUbbq2+U4c9GEvxLeC6oW2nhkl0rbxTuRqQ0wfxA+VUX04z92oRue/3zq0O
E++0b+dOe0AzM0B87fc/Gg8AXv0a3b4GNgr/NJLJCWjUT0i24Sdt91DcTersr8Gb
8XU8Lodlv0K5Nj7cb8GC5spCLWkcSwxYIJMGwoAVsxJoUq4WNfxEaakafFfkoA0v
/tR1gZoNSNLR5ENnhZL8dL6XgJuQaCvjPZVFC3RcHCV93Xkx7Hlw6SmWZu+vWm7c
tuRxpBUHRd0yTI+G1eox3c+Bu7VgEIr4RKqc6sVFxv4G1FvHd9YW9rRJsZzV2evi
x04V0G3xgKc/ISWvEunDMfKpLuQ1wPvdWaSULuPSqCHAGXz5OBbT4S7X0OHUaPu7
JONL2becWzGqn7YQsxG09txy9hJCuflZyBltdaog3a7EW0aJi4jJATcEQhGs4Icl
HeWjCtnljSnH9erFkYN4crBXczSTp0zBZj5vf7+pz+niPZ5uTfX7rBG3P3cKAC4Y
6jq17mjpDlTuJy0OW0Iq1ecltasQPJn+a33sRS6+I2WXz2dT4+8GB3zEjq1Wy9YK
atQgvOK6Qi2YoFUaDuDQUz6GV0Nx/A9JnrSqjuFP+97GyL5PJGqv1jtDzCin3wfg
sIz4Zyp0NLqi34i2Z8HR3zWAewKQzdj8xLr5dhqj4NsIiy6F9eXCBHXq6yLiFlRs
zQjvInMaFrpl0Iyhe4I6+QKCswvwk/ZF6flPaSF0CfKvd4FqQTl+s9lKxFbRrouT
TwzCyuF5scMBDEVKG3OBEvykom+dzVv1wP4cDHN2yhGgQauO6SDwZz2oGeQ8Oz3l
7XsWldr6tJoO2BpBMX4vIeU8QyjPdO3u3SNKi/KNcfiZQsj8MAu01qe97BkHHZZ2
8HDaA1o3yQyUT+nDR1DtuWprKB+d3y/YjAh3P7KAvwZbcT+RBTjEsn2y4/swByMz
yetktc4E9sCb8AYULMNYzWZIHnrKZfT1N/ZG8VsIZfj55oerfG0wsUN1vzt+0lxG
9Qyd45otF1N7a7sHHCnyk6SDtcJh5fEyBnhCpTr4HfEeX9omvy10pYoDjTnGYouj
F20L6PqyuDAE83OjG3JLvCx7IoE5aeSBdwzQEvuD6Z2qZCBVlGcEqBEI90pTK7KV
1H3yf9pPKNSiWNzeejBvU4ZLNEzVw2/x37UohqBsD8V97KA86LrgGPN9yjnvmjCP
SqmQgCvX4IqAzh6lx0WC44GuEFMdhfOngkVq6+Ba9sBvxwxIGfHFSiau7+lwR1OD
ZbK+TmNl3i7blH5zfQvlQJYZ4jVrwSKmqaRuND/H24/Lp6x78QIGh8ofr8cjNyd/
F6oHzIYOV/oFy35Sl5ipqbGeYmx9MaFQj6iEuk6h0gsYOUOaFIDNcz15KqRp7nQJ
l/9YV32UE+f9jUOkFsnCjCC/zGLoPTTdVN0A8PkcC/ywTzIhpInXDAKfQPLH0uwI
6f94txqX8glQVaKuLtsSVylmtOderZvKUffVoPExabIQ9S0vtVKFKLq6DVy9y6Va
w4NDjniwmnXOy/JHdbMbEVIDoCtFi1z7HsT1qD5aZ5SGEix8rtHK7y4pRnF7+fO8
W/xe2h9YZ23zhY97gxnFgDK6FHN6xMs7gFMHI5f5iBH38DrVBXaVRY0faGRDjQqX
4hUkmUGDam3ScTfVJOUBrJyunJ3XVW5TVvUAV9u4kFXyrXNYJPEE8SAZU3/kUCzI
ZU+HdClmBBaQ86zs9LOcq48hem8f3C7tgIcqpStsvAeW02tXVlqHNnoQZUCeQbRo
CC3ZeaujLrguttTrRrSlpagWANYEV7PboSsGDFuOszUwgnVdxRNhJ7FEiZflU21F
BvUyCClRKlDJBfRbRvnT0AsWxwk0UxD/PBL3QGeACXTvnk20Wn2Uo2U3xLQ2nNjK
qjICbUSVWPlB3EMpj+0PWfWBonq7XWOUhRU1emTxzqXzO4ybNqEcS6fV5UQCEtPd
hGZj+c1EPU8IS7LSbegMtyZumFmG4hLmsc2xrzbeGdtkzh8PPCto6ZssYqdIJOUi
kTBgN90FG/8HWvKUapzdLH091kcbzazMuXpYqnrXKE40AIUTJXjFgkbQMtsLA9QK
rQgc031XAhfFqSoT9vzwSISkFo4L2PgqUmrbW3eGBby1qUbFx2kR4HVdKUF3gjbB
1KuIvqvrWiG7wrGedC/wzUNAtntqPC29EOCXTcued/Q97fTZCuVPXA1wrYD4YUPp
l7dTieXl4pS17VdERwxtYVjcpIAI4bk627UlkbJUTU/xEUbrcKrPCghmrjEJbiD4
gJ4BwaLY8Nu7ePzhaLmRTHaZk3+vYLY2eh57KgFfJdUhaKdEd97VrZ18n7Se7pwh
6Z+9Bd1eHvAEur613jwO5BUJyTUw8SFYbq0bTNTRBA3c/dKUmyoRClhx6FjfVgAf
/HTTT1ca06/EIg9CgwGEGGlS4uj9z/CooA3m9WYfK9748BfLA3ywPIDjXhtiPg6t
ULqMfB3kR9xnInRydpU7kPP9wmonoxuTgDCv97PHBrcpXnB1FLx1Bz9PANYlCl/7
fC2K+2DjrBHvGo4xmtlQwGsdBeX6e3LrK5SMV0KJaviuqT+TnLTKEyWBO+VRcvLf
gmOcsiF/GXS6bvyNm3E73hAvKwMZ7pyUlXEOJX0YZ8bmiDp/MYXn2+fDZ5VAFF8m
9utRrmFgZdonv/f0A2RJ1Pqveq4tS5hAW4bngyVAewXxj37W4hHM2rVDvtUXUUrG
NxJU9rxr2Wu4sVjLk1TlXZaK22rnrZG/1oA9tO0UNwRL3frqF2Yre+HHSZ0PiD1X
XVDKpKyFDXSHoOzqnXSSX37jsN6WrBX3CDWlFIkA9nWv/zSTMAu27tTLMgdd4Nfb
TPrFGogwCdUo7dpyWA5A01CL2+BTRCMj77pW2eUl27HJ0FX1zOZzgElrydGjpRIz
Wq8Ix5HnUUCpMDibhD92seOXsGh9AxoFOmSduq+1lbUFocEsswskeQC/taHVaSBK
m4YyC8QxplZTXAM1Jo9Mib1qZvtoe9zqRHZI0+pMFqt3Us2UtOjIJrK/ypDhkVCR
t+xUd2IcFode+uRh9N7lJ5JFT7RdyI78Wl7GA6TdgOwYWy1pqzynCt/YQtaxaZJL
dNh/8xKQxrEomDThc340wxBTMVltBjw0UbcDAVrUYCm6ptDT0zhvRsTvl28swJcK
vSsI0GkS8Qxfio5fGRjdCL7NyPa+9G0oXibG1Bihim5uvroj5/TDeKYx1IlrBWQi
sM0tWJC2YrWHmd42Qzlf3ca75vNbK1usQwofqCE6acmUf+rwevP1kFKzOz91X83S
gWgxrENsVoe0NvOZXQbKnfcmD8mRoQZq2pen72rWrnrQpeDT5Ba3b9je9j66MvMs
EPenqMXk0Hv9GCPbzSqC7WqdFWyNcujm+BEdKZMQhbuLVkNX9d9Pz9Ije2OU9D/k
SkJKelthAZt3kWNUItuLs+TGZ1u8i/zZRXRBg8WUK95ZypHTlenks0iqK2Dwjxwf
5GnU8YLP1VAU8tVf7PEojHJxRjLHaNBxR16mcx2ivHM+ms1x2q+91AmIxEFJrpnn
8YJplhEGYGiyJTah9kk1QM7dpKN6AGlffj4gIEktcJB5KWcXqxp6MT7lrXijZZTu
jXq97j70Qzb3GdKVb84aUyqchpSVXXqIx7Y04f3De3G5cJ5WA9ao1UUVQlOkJoGU
zhxL/bvfzrEMJ9pP+jKKzKLWZTE3b1nlnYDyz4kzYYCHZK5Pj02QuXNXgqoqdVE+
klZ+hhOE+pnoWzGTzETUF9RcdJZ6yPpuJHLMJ3nobsA5FFzoK7D8ZiSVa+o4jCSD
EaS+hVlq/ysuq+CAiyQ9Ij1QNXqGRgGJlkoM+dLl3Sm+89IpSDTCtJnMvdm1Oa61
J497dVhL/xLp5wm44uqov4Lk7PD6CGOm1wolq9tqurkVliepJJicRClKeFLuEgEh
XYZYazkyt3x6DWGtgdPyrmzXK8biEtXerRYvWGB/klk7yLM38DFagbqldHxyNrij
ltLiLSw8fRcr/efEcTeqvFOigkH2CBA66T2TAjlZPPPJhEkBuS2agpKbuX9ae03b
sZmWuk5JQUUkKmgpoMvcYHFgAhj9lU819iDA6TGIJdub5dC/B9ysWttT928dxM6Y
gefobTYG4+kwCHg1tjtmvXo6/LLivrWhZjZJgrtRSVkEu9/9UPdo3Bl+K+QvpEKf
D0Qpf+qjxy1C/z7rOr6wCmcl1B2OZdFG6imn1NZWTr7I8vt1bbOuR+5nyhdomoas
ugVEG0g/QoiPoMgqKst7MXG+F6PvAtT/5S7ZkikQ5BILDchVJKJQq8Za6rHOjMph
KWRDx1dvIfdbv+zpwVzZpWOE76A87ITorxP5jfOFMSGzPM6cWkPFCvFKZdUDZae7
BtqCIxRK9PeTMW/BYisGbAEsyad0oFCDzT6zg9O2CBWMtzQlxlso6YZrVmeeoB0o
6iriuaP2jmILCFKkHBIoStUgzSMH3iVOY5OmqiSbw/X3cWKGT0s3IeAQOkZDUZCv
6B4Hml+oVURS1YM8679mDUO/vvPS4YGNugstUJ0LbbTJsMqE1SPXRHNC8+V1j5jj
wn73on7qSimbRT8vahvu8SYJuRO9b3+Y/gkCRfiCQl8St0ONwFLmwoOodoA4KEyG
9qPS41HbgyC2/UuqD2Mmy6K0FlCb9i4LxU6NKCc8jupuZ1aNMsUFG7iQvXn9ZwN4
7nptrvAgTNPH/vUd6uNm/cI8t0c1TMYW/CjfuZey58dkqtKK8dcX7aOrJnoDzVGo
hrwMayTMxR6U8OH1flhXqiaeP4tt1b/Hub2c9dTvJFQkV7uFhf2zI4z0fP6DOA+F
oczTteCtTmOPGJ4OLLHlUnM22IjyYS+EmnFq4bGqmMtzSZ95U9J0AjYaNKa6r1FA
mZjJOLZyst/bLuGi9oqtLVuMop3VRbGmd8pYQd7Kpry3EzHJXlWms5cal85oIYhh
uSPbrPFwx0izjDUgr44/d6phGX/ReBKt8jrWBQOLfNPIraUoTAEZXi4GX0WMoYE9
wU8kfv9vQG8LeAmWfCVkZIXMKPNVV+d0PRAAIBhhwOY4V2H7UcdiyVokdqnECTNd
cyZWmVwxCSUPY+At6utCeujGUVnxuuPpmOb4UekSqXz00NFqu/XI9+109cxv6WEZ
g8NRy36J/7Co2EL5DVTQIOU/hr4OT+2XRyjFEsE72Bn4CNkT9tv35YiEyeyD7mTP
YUjQAPadXtsxirUtBZxAMemuSF0XtBQ1VGBSRdy57bPxewhfRETGyFkHHAa2OTbs
n73i47fmC5XyfEMjx1UZ2gtXlWTGxldrBkrUv2xhawANaC3LVu/LBOu3F/eaI8J2
rcL4DB4ZjIwkkv+TfnU0xIUsE16Yc3cHdkqH89QU7Zhs1u5+pS0vZm4EK4lsPF2T
tuBiHA7CVXCfjR7VlmT9dFOxG5o8HEz/JbU59/m29l5ZB4CTXpMarzwKujEn7EJt
2XHWsfcReIBKAZTbVeIkqT+u0AFJx37ZC9EIm3mm6csZuQ6IefszrCHqd3sx7jdQ
31OjMKqcoCuqgvN6yc5bnXsOTwz8gsCWbUTdMbEuOHtoNUBtUC6XphRJ3XVKkvXs
yiFjirlVHKq53v2w1BqzJg1IUobt0QYIT1SWxY06LP6beie3GceREMKjoKPsfD2l
nzlv36h/A3XIe6EdduZktAcssWooc5a7wp1f9T98ygYltlqNaqFZN3PSgdIAgYyc
siNsQkuMbExuMP1kR4OgImgVfcgft90GDUOYGLd4A9xhdHHb5bhMzT8LNWVDu9j3
Rllyb/h096Nhi9QCFHWUC9/M9t38Fr8qPZK+JU/xABZCbZ0rouGvwEXfo1XTDmtN
mJQJk8qlPkdp5hCgmfh8sI/P2jwJeR2+tF1BEogsSuIeCnVfB/Lx0+NDGHDGbG56
roMTK3dKtTUeh5fDDP5huk8hStdRsR3L1xddsIGPCl1oN83x3DVWEl5hS9ZLxUx4
WHhcXygF3miFJrWRsFSxbxueevhcFeDCIO17l2V6glge7PZeSKg8kNpf5WBlB6Cr
I9oFl3crVJ8P2TMQ605nqxKixt5yEaiqtayZ7uwqCUoUu+v66YTkjsXq6xoEJArR
gXOMjXA/VEaAX4W2aFqEmn7IwwU9u2drzA1amQNsSMU5wyo0T7PVmBu1QlSwEOXH
Oz9o6VSat1RR7zgFROs9T0py3BwPSK8au7VW8gHCdOYrHg5ct9gEUYpwwoKvLR71
sSkM2NXy17sZqP/awswEDWtH0w5FF0UlCoswyyCkeae35nJQlkXEi7JmdIhuaIr4
ncyegm2TZv2XbO//RVp4eLjcFxEBnWevjaTf054UI0RxsMeSPcDZ0kLPm5C020A2
koMBXuCV4ehFr4z/7/OYykROgsDT/iSVOIIyjoFA0J8Y+JSFYKzmxoMG96fEU0Ha
qXv2syFMhBFoL1W4P89vRE/Vs1AgihbXYjgOndZfqfycbYx/37PGS8QY28xBWQUk
i8P0e4WZNmzpqICiZ9dBDIyZqQU4PL3RjhN92MKoam6wr2bD32WCFIWTSt8FDIsV
afyuPXHGJImGCJSiPSG/6mduCN0fBrFoE3uS4LVQLXm8l2pD42eFPbbxGZzUh1+V
fZqHxlHPWBJW3BHrRjIoN+YyC0APhuKs1nTKmJDJmdy+oopK/fdT6e6hkLZ8d21M
Riuz0hY2IxGTgcrXlP8ps5+LuHF+U78i7KsSYt4o5DU9jp20KfRgdoe19hNJNddc
2AGUotBDKOH7/TTJOKkTjDjGjaQbCUBs643/EnyCvc/fzWOor6JmKtkpvGABl+th
lsf9nCkS3k5rooLC0Labp2qT9spxjQlOP7R/baLq4LaswPX63alxeP6cKpo91Ra7
Ayew+Lpouf2bTno3KEgRT/IBsSOijge7OTzhqhBIXFXd/OZXIwmK+6FmnsjcolSa
G79qTsvpR4HQvd2c/Y5iMyd5HpcFagyDJZkzLcaEIBXi7JwAZq6lZwgMfZXvc05h
f71QttLWvOdmaU+khCot/UOnYFMNCWUpE3sGqvMgza1QIwWZrocZa/xEU5vnDTFR
7Zw5j2kNfII+iMO3QBP3auDIFpD9iWBNQApNuKzISR0Ktr2Lk86u+YKI79Y2mJXq
WR618MdzBMggB29x5P9c6el40ie10fLodCYOpiQeD4jZJcK8JqLKthgxqbjs2Qvt
5j/kPMsxtqd9HtYfTPfgeWaLYPdCDxEA1DyD613iAVqHIuMDSK9qD6L2ITM1vrwF
PHfNbnPavHiHub5SqGb5fDyfe95JhdR6yDGPj1DMGxhlitWz/NmxhzetyrhOo/fv
vIa2BBevxcHN1MEObBFjI8awMBBVXFjgIJMNkC2ZghfbB+XLdNkHNQcwxOPukNyt
Tl9FBc5Oi1I9GI9uxgYQxqtV3SVw9fHYMVEeEMATzdcERjzS15PtnsGH8lGtXsp3
gw6f84Li8WLkS7OB9bglfdeIel8HqY5HIZIVM+W8JuBf7kdmUxx7It8DnzIJSYVN
ZP1xCbezKuORN2tRSkwuvW4jMm8iFftUzvXUvoASRHH/o3mlDLKNnCSq8k15H9qn
KkCziLpGlYYYbS0VRWiXEsEsQ8ZZKUAcrwq07GNGFrj6eFxCw0KqoKAc/wsTFjG8
AvHAsS6C4Uy+8JkDDh01EQaNX5ZQPOsROF1pFgRNAX+AR51LBizEF01phoJgYNYS
EJRfeQEqf+PwhU/YccfXZ9hXmzSUCSVAgvXu/H87hONlbRmLqzjcyLEa1XKStdG+
MI8b2JHhM5tbhVOccLhJvwBTCY64PsIwmPEGADZTdA/jkW7w96qWZv7cRpvw/jr1
1wGRQC5D+dwzaiGlzTAptL9oTzzsIuQkYQaK1xMokekMGivPEXuJ23EQQRFkwpMs
biQP/Rn2kx7arD7T3p8PEb5pyhOEMpFd1LvfnLdbTd709QXnX8ryFF29uv1Kbp5o
r2XvoTmugyt9IOFMSsq4ZCUfbTdAYHS7JrsY8NSRwUuFdKt5VbAl5TFYAVIbP438
gE7v3jZqK/soBBPoXsTNJe8hDN5t1Oay4cetww2G7pSAAVzHpxvg9zoluuWJz+KY
vMe++IOozu/d+VCpuHA5SBg+LaGRCUoXmy1nPx+qiOTIYNEevY0YxIMG0Fuzwk5m
/1yEzxIQDntg09gbOBqIVcR8J0Xl3Xen4f3a39iuBLFW7Ag6Efx0xDu5obO7mfr/
g+sJjO+HLsEQsITRrWIgniej+JUAtsHWuBhowLLvzXQP7Pm5qUyaoLuCXpsbgbcn
5XcE1/TOVLJRVMal3nxsKd+zzOk7YwWrTLdUWZt2OHUwJJE6fsueRX4sE8Bgxdpw
EvUQUs5qpLjklezyb+WRLJa6LAqyvCkNAPm0MfGpgT/3BXL+VoUy68SpYWpsvqKD
3MHN0zJp5cwjnQSOHNJQPzoSOEY+0YR0yucHXXzlLr68/mf1cXvW7P12x5qmlADI
IoejY7jG/7kBelT8SW7FDziVANcbgaAqTsgavSV1WvIFa6q6mxaD87d100y1wIYA
38N4+QBK1o51lGPp5P/1tIWCFeBkteGq3bzDoKuEXI/PWA8d2Bmcx0VHvZ8PZCA3
EU7hbgKKWn+PRWj2i3RLHIZSqs0Rp8MYIvcXT8b3SXufm4eb+d1y1UQqkeC7lDDt
Yauz2KsRb1U8zlwzjdVv2Y6J2/gimORyF40Y9oeafyubgxdjJaI2OVWaBzdlSkKg
Uzg4MrsagotpeHXjOlqweFkzYEQUZsA2V2ADnaPszOfIqMJu3PDX6qe+H+rdp3VR
IdNg+WbLdiJ26UiOdTJoF+j7rdE+vjXS0AepGtl1sVbUw8b1eTYYz81u4EtVbspI
WOyTbr4tgB85jmTQx8dk/0i3OKOkMEgI0loLXPkTjIP0tE5UItqI/cnzM38gdqWz
uDbpJusxpRt25qHtolKkmeqVHE9C1L4i+585pgOryDDowuwYaUqttqSgMqyp3Ooc
VcCuzmsBusdyiSHyi4To4VqoH5kj1DiCzssPTXioEb4ngoXJMz8zLnfjMcmPXzuo
/Q7izNxMtK+lBIxJJLQvzQA9Ft2ZmyeLZmwTBmPb7xIXnyv6qKbAjsEQECGq1ZeJ
CNhKCQaVs4ZLc4/uKwtKq6TgKBmiCG+55hP0tthXhqra6dWtsHFQiDE7XePHVgNp
skiAgjOSLWS6/pny+eky8tGWa4ZVISslSYGmGGNxl3zmfajz+xhY1WAv9DfK1xsu
VAWoI7Tv/e3/plogazLllRaC7pFyOxH/8bZE+Ozof140IKZs0bPd4Snya6oFFoVF
IQzoYtaNPil9QAYJL4bnqKKt2I26MfeyF0ijdeZn2c1RfAgpE+2pY8O6Qyh/TAn7
7g3+eJM0yoWKqPaipX+daH0GUhlilszUFbOsWxyrDMVCfRxFAE5zDw489/gqxYWz
hHF8ymv6aNu5G4PmISAh94cn/0wCOs1tnunFnk6MW6etK4cK/JllSPsgRj4twBLG
tvXx6BQ7SIE2+aMh3o6JsCzvjMvc9TB0PJ69e2h9PiystHyrp9o+j5jHkleFXBlE
ZNm5Vy+IzVsBAlxEi+r3SXCRcqNeTKSUKkKEeobbPQrZI6jG6Zw95cbzts5lMnRP
YAn6tUAIBtKlODf0W1tmRpO8SYJEN6IHUY3octK2D7TnWrBUAWTApiqZNvXp+TKX
CLHODLjf53TmtxD06d5Ij/eCDgCn0KX4cDFEF+0lyUsBNzJO1oAAl+i+qZSikwAj
+VPzo/+NZHt9k7wI+H1cMITmYp4itCaO1/ISAu37m0ejph9pUSx2LK1gDhs8KvV/
oBxBQAFGGgBIZosgLTiKX/SqSOtr7uDG+6Fhq+VjuiSreuTffwxwgqjH1oOvmLaK
hu8L9zstb/FLZnBaWSs3ey79IyaUZ644o5sUISylgCmlSc5dbfyHXN981QJ5rlCU
XqroEEHMtnZ66jQcFhgrb2BSIykW3lkVyTgHHsXQzX12edjgHbe3Ya8JQyCuKpJk
AoShwdioKj23WiixJJybGMuWnR9UkZQY5kjwF3KHJJ170lfMal/1NwT2IG7f2NjM
9LdtDQtwbUBCnD1NBJtLVBTmOMloAknVtD9NLvAxMr71PZf9dGz1QHi5OeStQMNT
+0LFM3QHxwVzAyKZ8cP1ItCYa5YHUKNY6xi5dsTosZXEA7p3RJrLPmwf5/xXtbTO
9FZSeEgu9W75KCvkDXJ4laEPqxgzCGUY+i0xgG3bS81i2DwxKEcX4Xq1vuwlak3z
iNHWGrdgNlUCRr6FII/Wi4wqWb9Gmc4g9WH9P6QAudV5cK02OlPpKOT3T7FiVBwr
ak7moobn9dbAxF0jF506nuY9563s7zKnI0yGUUF0kYvhtwRzJ76SU08Q7pqLRVat
dS6J+Xc7ww8kB+3Vufm8EJrDEZ7sgHe20d3sgQ+2mbBsfLmmb1lGB1PJ6ENowSWa
hxjCX27luH7RmoAYQgqzDLf5iwZrOeRCjwphoMqkz4jWYfy3Zm4y41Z76MFhJdi9
A6anKIoZkDXxTde9lTSTNy63xxHRe3MMv4DF/e1srjg4qN5CuGHrIVe6IC8MOhwJ
X5b+/K0dHq+MGCMBaUQjPVlmRE3SyEcldK59y/f31ffbm75esQ3cUu7V13J31ak0
jHOWycbfCWy71Oj655qkCr56OvhpbYD8Wi6IAt9XDI1fpGOT2kv0JyWlIuUXKXA2
MdxJn5bSOThSyRMBWqL6y0pz6IXNqb8ENyBXmeC8MdM9Ut58xb8PEXmio2y6P7uM
PTOqf/cXdpVlkNfEp3JPnTGl5Q34+IShfQfszHhXgxBU0znOdUsoqwep9Rk5yebZ
HLPNUSTPQHger1A7Z8A0YQbZqKVif1AcfEeDb2COQJw4HYOanLstXpRX6Rkyq+o+
CFgSCAkC/HFeQO/VGF39ZwmFfcYE51CRN4SAih+ZQZGwfoizWM9fLPlD/P/EBC1p
5AVNLoB60I0b/+NBvL5xtnpiR4O1oNZXxy7vw+yAxScqCEyaTpAErnHB8SK4859g
mz3ikp5JaPuTF+a61ghjy7BBsN2NSXJcX9msy0Zr50eLvh2lZ0RjJr6WajRqWfhZ
ypeUuFx5jsmrmhuQlF6WSiOERamG5bdyCMun6VP/S9mcDnuICW5PvptYhsizAwFK
hV9X1/DvPSwhiy0/m3Ra+OdMaW03HG9wM17BVCyT9KLnKPolaPDZoYu/kUh9/Drp
IARVPlwlXiHQ6sSutRgJxQVuGVYr20XNHTbbtdK4xuD5zI7BWUO4M1O2h2tesjMr
C7aMZvYGdCMzBNs7iW/O5h8lHCvKnlVhegRuJC9hhiXVigtAC/5zb6rBHpFPt59a
4zuc7+tyc+yVMXdaNy1y12HvCv+UaahQsxytsGResRlDoTRCGF4DXZRcrgF+F7G4
jnp8W0/ZZ9ix6xYsE92U+5R7U4cXr8oouDe3lyjoCBfm3jtZ+t5c5dBlTruTxhEq
MPh9fZpZ6ZmH4TkJchlw1SLLo1Jaf8R2xXOgdZBXd1NOS8ipU/OplA+Rf4NFJWbA
5F15EnbRH44FwuxpGOI2FkLutblmFztxKIZVlN/YBFNQF6jBVMFRV/I4Cuv4lkzM
1pedqPtUYUjYVTRz45upsA0Ufw1FJWwMDNUnTZgfK1q22fQoYJnsAne36fm6sIQh
UqrZ/i0vn9yi2vHghOdlc/jX7ElL7uqEw05mxJzGiKXK5xvXayaGfU3GVeWWairy
bdsH89scjhZHCV1rLPRjygKscV2ibF+8Jl9OJ30Uqc9VAJFERBSMcVvPaqf4qui3
lAf7Sd7ByNHoBGdYH2HrSPAhmbZaAW7clWbOZLw2g9ieYYc3WCe7LepbRAsMPvDO
w1KGq08j6MwpT7M06MBAj5zzTfBNp/PpD1/uDObFnWWNfHGqgi/+CZGonpuUf1s3
NdkfLypAmXXrY6JJ1Y+uaS7RPslwCqPzMjwq4Vr4nFQvcRApDg5+2dwGPtriDaPE
7+sqQvrOD7Lm+GkXjT1up44xrWOiFQ38SGSyQCsenniEkofrkFk4amyjGWmoDRyh
adux+KdTDaXXdG6dKT2kBYRFJXNPSc8PwKGT/q5a5RWLnzBInTb/JzvVld8pQfBZ
3r/Z7uwFqJ/yq+D6Y5mrsgikQysa35wxFQ/X19+eL5ilvRYMWp6LznqEarvGoBA2
fFxlI/j5cS8aTKDD7HhXpAbnaMpsEf6fOLt+LUt8RQRaG8+OvDWj6kPUcL/jMN9I
X9GUeTvsKdBOVWm4OedCmMd+0d87UoOX9DxbNGDk1rEgfVyLgSexEzULKLAY5qFR
jyAzlPJN08a4+sVeoiuZDykhCPKvor8s8aUXg1d3dhQwSGYn17GY50vUEcW7arN9
/IJAzdqPBFLODlrvVcGClbKU0LmUhplIC/gpOkTZQcRHqWhSIRaF/z3cjRVIJEJq
l0JeI1FyMUNZwJ12ulctfI82T4opazEidAk2kgk0RS3bo0c/kszAfD90efI3cB5l
kF3Aij75dL4P8zQt/24wmd3HtmVQaLgr2HfUs29KSGjR0vwt/fSy6ERkCOXOuLw6
j583a1xRIpikCF9uGFEd9NIBziUWCY4PHDDlr5+h3oQUThJxi2JY4nAdHjWBE4Hf
Vtm4zcqwuq+7S3NXKcpD8yST9rntGbKtbB41DLa0pwVkDx/8ra9Kb+KW82uwhV+M
fQLqC88MZvutWDNpdqMFgPkL1INSkVyjFQ41rBUtv7vkgYjbhts4/qk6yRnuTZeG
ugSp0nbJrrPN1A+SOFwXwyZvG9b/qp8jmC8yv9IL2jFitsQUXhF+MZENfnTH1IJM
6VDqZyA5kDFUS1E2Jm7MopYwTJyORSqohMjVJY50NOJK2IpCWDvlXUqTxje/a7t6
5iIPrItGPDR43qVtSX8/GdYo2y0OCOCUoAq/d01K19U57vBq0Fst6rP/jGnhORjG
stmGtsOn7dpFprnP/PWQ10qbHRS8UwFyM4CVOn0KV9aaH2ttu0LVRAVh1kGNJ4rH
5vtXns49Kyfft1DVCIm4UBL4tCtO84A/ctQsdqiNeh0I56htFaqVsSX1EWXNPJTj
2O4MhNy7INWSv2SSpXVDIbZq2+VrMeTWP5t/WVnWe8OsdoCewjD8LkLTx0to9KRd
MfJsvHmmAZo67Yjr2VKwZH9pE+6c3a5zXbYLdU6tsR9V9Qa05L36Kl7SeDXg4T0a
48Vlz+za5g6q+D2KQ5qa/YDj3LTfQIsNO+tXAUH1WN7urM4pof/hIFALZ9V+NZ8s
xTqoEksl586l6+GUZS+p7UkmbsEa61TJdvkEteU85RCHD7jIFZr9E6uqNGb8tQv7
+yjmvQd3D07WwWiD6VLufDz0fg4kLhjqP626hrQbF0d4IfQRUnjMDqA3iIMFejdj
NirXsLsJtRiVyqK4R3qq1HnhTVARfVaaqy6J1LXH5akqMZV4aBUeegoCs7JIgJ+y
o+dt8+J/v4rixIqwl+Ks8R82fDpuvvuFE482NfKgILvmcS2WXLMBxXQjWwSNPW+9
kH60j3vLuX34r/2gad4I/kEceR9j9a5lwJ3RTuwldWpPWVfvzyuK5AODmG6BUQ+R
+j2Ri2ihvK/Gc/CxfG/wpJwrmlW0N7xminTz54JfmRB8YksmkE+5jzzmfj/2wQUQ
k7iqnYQtRrckZOeti80z4wHxbkCIjfcRtWA8REYvQ/egE0nJ3mcGfylE7FVw1bZ3
Z8u9XReXkgK+fV/ohA6/bGR2YVT+/beJsbnF7Jb/1NdmACNSVbFLOj8gYpixWfCX
HEc/dzc0CA6NjMHAZdjbVpMQqg5AngiI9gPJ2srWUxp+CNhx9LQ4bcGUlVk8cFIC
CFNO4gpw4zGOraJ75taQ3JJGcjBldmg6AyVv4KCHUJOJFRkJF4e1hnrCZ6OYaZbI
WTtG0gOcNITEaSdBwKfVJ2OAQ2Bi5HJpVnfE7LVbBGu32wbdeM4eNP8haLeWsqWp
PW0cuqscF4iQvuvWW3jOU75lIJXHkaUju/Y69KwofyV1JRr2OIwoQwKEmG9xA29F
TjOBTKJ54QsGRP6YLq2FCxYzK1XhczcWatuks+I2amXYSALMrR+JWemJbzmNoUcq
O0qZ4ihTHaOXVOE5V4PlJ32zYlN7DVT2KUbH2j4PA+an+/R5FmFz/L6xzVMn6fSS
nhNew8aTf5HKXxQ68s+lYsFdNF5YcFuTr2p7sW8gt5ssP61Q8qx5V/LbP8UqADjR
Kmzj+Zuw+zJ8T0prkbqGz16vmLqM9Qi9BXdCdp1ykhYJ5wJt7YfadMkU9p+YFckM
OrxIiJ5mf6sWThH2yRKohfm9GJC5VlBp9hUCKKnhqRy5D5iAu3OmyRnMygt73HIT
UpbcESTe8RcL2w9thFk/rwvB3ePvP6FHxDSdR4WpA+smJGu0w5lbX+oARNdFaESh
Q/JpgGVWtlX4/tduK4gHLsiESHxMx9mZK619IJ17/erGJHehcmmNj2pBMpfVRTSH
+cLs26Gba+aK45kQFQ3TZX9k6M1X0/ah2A0oX7MDb7PeZMGIrnq5xVaynwjNt5fx
E5Z3W+Jx3TVBWIHV8lH5+Ca9WPxVS5zzTnz9Phetnf+Yx9kIqJcaQyX2QVY+qKV+
ibe1GPDSorBIVcNtFfI2ebF2yk9A5XV4VWCZUhZk4Jdeb3g4ZXZmuFzl6EMMjM9q
XDVXkKBzXX1zKhuRf7N0xL7Fh8w14eBsWWTbUSQ6psuDc1+M87F1j+eWbEYmMdPa
8wCOX6306jBs3NCM+tx+wSZpBkNN8fiDx+PkMJv2c6mc7Jn4LjZXNoyHHrSr2ZN2
fxHR4pexs7xpr8pw2Z5EweO0SgTYvTbj0ZTiG/tB6ZH6jAWkXFiiQ48LhYs50zl1
sjrYmLDEaJASl54sgnuMgtI/kqmBx5jFsopdBUrJLUdR/OApWVQ3iHZDn7EsC0aC
y95yflyGF8zG4O6UnuJhdpcIFHBTOERYjrdzC5rTMa4tvvFrF/O/c8JKd9XNWv2E
PKLr4OFGdI1w97S1vBCsW5m1MWD8vxQD23vA8q7OhMQAh+3FillBcy2upoLr1xi+
zfsZdEbG1fMh6IJgHnCvNBJw6jz0lRTFo22Idasy1tEhQYEim7med11DMuA0sGoB
6euCTzee7cTAurx3jn+kH+7QBrZdVlA1m6bwZ9t6oegaarMXu6JFL+PtLtACt47c
Yp4iVoLMVFCnQHCw9VdaQoJb+WN4bYeelVK7AymkD6fEuCxJm3A84E56V/10MDBk
mvTJYdT7g6vI7CibZIHLtQZYx5+am0cFQecyX7/uTpudDiPnZClSa+1lxjZbbdbt
5LlxCfDSYj3GlCwSkQw0cVc4gK3sLBfE63zT8/T027M6VyVPktMeGmBGv7ync9ZS
HHj1m/7PfForbFGAj2/zgCSRWRvibczLT9B/WargouxIVR6TmYw0cc17L8xpdUKJ
5UWZOkK+txaXbzgXNPxvvG/1Q4j2LMXmeTm6cFwZ2oOCSqa4v4V5CiPg7/ZJMtKC
sGiqsIwnfVufcpypB/1975UmVSL2YRLL3pDHYBYGZOv/0zribCdWKsCygRcrauMg
USRHbqYCWyqOdZFmr/sw4q/z4MujKb4PmK/k6TyY3cMqANRZkJcpbQF1ue1HicsM
q0mQOsKTPPIsmyiSmU+m3JXprX1vwckkczZeU1u7G4womkfcFyUI47O68IYRoT/j
FSqRKGf12z7hNdWeGmkvJwQCWwNEUM7zvqPm+R1RsYN8kFnAvsMD0jL06Kp0tI7W
vmV32L3KdL1YJFr1TxdST16uptiMvsxZ54AEPLh5aptkuxMLDuL+lCk7/srKlb8y
+sQ2LWO7gq7KBgnEqGnGH7FrKi4UpRbFOp/ZWnSvBxob2fvU/G6zcMqti6Lh6H4n
/OMwQFAXZSzWvGF1V8edXjR9R5D+WhXrKDnFa5T9DKOEzgYcDhx2b3Gp7PpSifHA
V365yC1/baA1ULAlEXW+UY7/oEJG8PaxO/TzgDXFXPXKyGHlAexTfwTp7jKzWuit
esaZPtekNAkmeQfVrdTMJ0jb5Wu+gTH9x/Wzf9an1ybs9sTdLP3ySMRM3oOFjnJU
DqquTgS5wkDdaoggh+XaS++y1UDvPCzTUPwyHTLX9slN5cGf5mrArfLw8iOaOfkt
rBOjn3dUfJqy3gYU0a9k/wMqxMXh6Aft4tMUD5s02rQVmKIYMkeeptqKIShri9jF
vFMQ18M2TrK1stkoaI3DTo82vM/4IYCVAByyX66OPs0gU6EF3eP2U6oPNyVFo3wu
AIl2wlePRJ1Nzf21qKFfNYxmWWK8xuDDk5UckNgEssYovUEyI36+uvPkV5bN2O5O
1BkKjLUkIgOUxVOw1/PcIEfKf+Ua/ehOALnAv+uA74pfuM4A5IvGsmwDdxRMdrms
zfkXfxEbJyH0vBkwt+EfSeTvGhkWBsy8HtF4GuCLyz0Igiq/KgY2JTQOAc923EhU
/zMQaSx85UuGEpKfmcyKPDJ0ouiFBrP4IbljvArBKwxTnvAItj+q8ggxbrMaFMgZ
dV/BJDYzADOs5OoZ4D7OwN+/4n2xCBoJX2RRcZW5rL5Q9hNuqfyZPNPnyhVdcUD8
yhY1Erg79H+xqk2mkp8yqVb6PZqusoLhS/KYY9dKTJBUwwOHeaP64Qtg0hRUc75g
1PGt5BE3+cagrpAO4sW7PqJizbEfKr3x7zMc7Qk3zFm6dBnWvr0E15zm9m0pxyEY
h1tA6QDHoGAmBwC9OnxIeAR4djJ/CeIpc/ThRzZYaZ2C9dF85Fr1IfXgJ/UV4hPU
yxBz7W0jSJf6es+UsOQRC6uexgCL3ZE5/LWnK9aoFrkvG9uCsx9UxngNYk57Ing2
C8LJ/02N+VkPLTlajP15eX5LV62Wk2B5on67DGzown9YlGYmCZ9RSIKSG0wiBzPw
5KPjD/SjIZBqey3BO7+ktEV2K49FTW4K3UYLbiHLVO1fmCmOSGHVpNGG9yVHTQEW
E8jc9xCifU6sderQ4ibk86NRuqHr2Wo+YxVUAeMgpVWwkMajmWFa2JLzX0upXIuL
UKSiYEtGZb5Gx8E/0Gka5Tg0FH0dyFpbE9EQT4eg4dyvdjpKx9VPuJP5ocwAmysf
yDXRsinnPP/58bwqQDSHCs7ZEQ1uNP3VczNAiCP7ZbwkR1RRXcWZhvRC+4sDD+bi
JMdB6RETW8tVs6P0kUaz3HT9OQf5U8Xj41wGGLPqcs19tnvB8oUVRl0AtVoV9QmQ
cyjQtI8vMLwgNBzXbbZvJ6BojZGKZHXIQ+IODPgAUXuVrfJ8vrKoIQgfcBJkf475
HUEiItQ8gybzmUflCckmAQcOik6Sor8IX080047CjpV7Oxa3cNY01aH0WkUWmlXP
TnXmytP6jQJI27XFcQIweSFWBMrKdwXE1bDqEBhBfGuQ5j31gIOmGWgM+qEvJaqZ
ffesCJWxUx2sdEN3KhYwDzkPn4dM3y/iKpoafYuNbyRgjnEnwFWJZgqj8j8MVv0l
Ei6Bd5MWP9HwtdJqS+zbqJkSQRd3oicc+6hMBzNthEi7bnETzH2n5oxoEhPgFna8
yMYYLsuoMlwvtbuj/dPoEEtdsuCaer53OnfcvKls2G7UmRjm3rIiiaZrOxpXILrY
arpwVcREWr+JJjBE0H2jq6KputIgWCoeFGoMKE9J3NYHcgr9Baxez1YiIJbF8nQT
469NieV1723qV9GacJu9rQHLcpNNuoSe/HSTzRgF/+9KD1L7ixvyz8gn02ZT7N2b
BJL60e9iIzbw5LiO8sH4oGXGT82WJ6iekZl3yLoweRq+wgHypi/oMvAvGBw0GjD8
mQ0OKpruonj/HKlvnzdCqaNqBkBbLLLJZMhjQpAt6PH3W9ZX3bvYO0FmJuUU407/
TGTAP1GlgcZzjUDl2bGbC9ZxNs8NFF6ftCg6X6fseAAl4MvsoOOuk3qJ2prCPda/
+2pX6Kaqc5jErkvCgdRMW1Hbm2BM92VjtA26Z3PbFFlLCt+dEFxDtRZKCrvnPtYg
/qkpfGqXW9JxrJD2zRWDw/9o/3e5Wox9rZxGl7RKnmsVrFgHzZdiMU3zpBbrVcPe
v17I4b+ZBcLhHMWMhGp4ZSwquTf9MFtbog4yga8JiJXFNUs3OJTL3P1r6lgcxuqI
asKPFGsZYfZnXDK594e6jRUayMFBGAuiQgSCy+QLGSnMFWd5wD+9E39b0dLkrF2t
0aPcOj4uGV/KsLR55iyiAQSjeMvmgmE2zLeaEW2DV96byXTWo6LMViJJH8sLEqVp
lXiUePCu34HsscnWH58vywbuCj/SXD52taXupQUVw+gNN4DOLlClXzE8TQPvAfry
+XAmS4vnaDu8Z4nxkH+ZMTy1bjSAvNYlY+daEY8dqcZqGM/dguojlqbWS/GUGp1L
LkqBEw+7zc3MgBilhbrphQQYYslfttBpdRvFgCCXcc0hNZojnpSmIUYLrStVlYxL
Dg/YJ0ppaMUOLSG1gxQ2+Tnqq6De9M31qV26vDXJevi2J/GodjIDpQScDszijfvM
yJAEewfipp5TSlEYMvJwn+tdn4ygadXu686DPz0RzxsSr4brcmZ/4sfAdgomvX9N
npjUl8oDfmSI/MgfJOFt+7ZY8EaIoQgKsFzyO/gEN1F7iysIUNRCa4LFHqna9YVH
8G5buDKl4mzFGICxYj2lNa5A6cI2iozfDm9Phju6jxD54XoBBwrKuHwGxtMm+ykP
4LQwPZldUZKjp9ZWkFDY2LR5g8YOJjcaCa/uut1JuL3pYTN4nzNtLNvydt2FTuoJ
hamfvYtrYXirIHpkmhcIUvFLo+RlqMJQSSBmv4BZLiQ+xbTJ2truTfYWhwsJubQF
XPIsAWwrmUrkOX93Pud649elreG7jvYThAFCfRNZO0jsoSpItYqHnS0rugaimCJ8
EwP7P4GBAA7zzsive18reVv1Uog4iKZzQS+9TvBcY3ZtyRMyxk3oBYaqOOm4ZUIV
unbIQoaWSrvo9Y1AnrXqugYOhLcGNqP9ZJ2m2zDMzW/J4kGdHZJmBysU/IjGdhdB
rT6yzTgA1rFHLYeuplTdBNGG6q9LmNUk3dgvPwAz1Z1JiGqP6rx7hfGPrJBn44EO
X5r1ka1Q2w4q2jQqcdMLRfBGyxtilKEEDLf2kneL7zravTLVSYcTftIVY/tYTS3/
Uynelf8RXlY4YGCBaHYpRZaHPhdPxnU9tGpAw37I0ji65g4Rzwo+qY23a8cr0Fz+
kpDbiXPYiIumH7gjHgwxsUuiFs2aXhcj84u2ilhVrepiyWRcIoJzP91EUGv/yS6A
zJgnBIzYqk/fQmzwW6n4Olm+ugpHim+uooaK7cQl0lLBAvJSRFR34qY2fGQOkOtZ
9NfQOfyBZNbl8tip5bG87g8DYUHaqYXR/tfXMJJLik7lOL35wsXP85yG5fQ77Qwp
ewvoHuMEe6/o8O5gqTpOHGEGqrHJqf1CTZFlA3VQuQ4VV4sHquwe+s2zA6MGzpH2
c+2WzbQO9BQ6DC14FUEJ3CQgDSm9X0/nuPl+gvZxCdNo4HhA6lGWRvGABO3PWPnD
cuyh9NnzCObHEJzAUX+0dxasomb2cvelJqDD7geWZGEHQ5HlXzuI8hmc9jhzQsxn
wk+Js/VR/qDXhnDHKisPCkKPU3Mp5QF6RB6gOKTzhu1m4oA8FIu0u2DM1VtP3z7O
EJsVbV3/OUexXv9UWwojuAf7KfQUQN+IHR/47UMjlcKEVh3A+DtmVW6Rb0AHA82X
s7WIJLMOeaktkAvsBvjoD7XQOdwnyfdZy95IfJXVjYPmxC7nlRSfcl5i4qahk09S
ksvHRksjfCQmrZ14XkboM51GUkD+bsQJ8hfYcYdlwyE4+Y1+wAWNz2RN7seIaxwk
uDZrPL/azSkC9bqPvT6eHgyhjBNXJMb5U9c5wOeBFNaCi/0RQGhKZOh4GRUqmSTK
mof0oL8KYiqvBmwSRqA8OM3fYhqq3wOnBpzXT8TAFMib89gRis1NJNOwxlIBsleG
W7jgJf66NB2C2Dz/9QDBDmowyusr4vV60zS1VoZLVQJiZWqspHJcJDWRnntKl1x4
TNEP7UxoEyvSx2xZbesToC0r7cuh1vKxr83FxPGLKqiNunlMLCPrqt1pmzSpqRrP
V6KgSAJ+739PGY6++kK/JxIKOhA1pVa/kAitp7PNY9GG8ZJEQ24FtvP1uPwuTlTJ
EDYkWIdZNUBJNc6+upggTHOWN7/mE4gf0mJTR4B69sKYz+qxfCTmFfRPlRt7rvtr
u6TfaBAGRANPl6HDueGLPAULtPb8DN/iPlNMdQLVykK/Mt/O6sedXuTpvhSndhf5
jgB60pXMcDc3PLjG06wi5ThMQfUWFNCRYoUSMbg6qqmpneIrXbuY2DV8fjYBjNKM
c2RZFYQgbumS729O9ZO57gJIR80kuqFl1ORh09GXAzSMnuM+dFxHM+F411GgY8Yw
P2kOmlI+doQ9Xw68gbRxw3umtDto9bQ4q0Xo9fUWqSVqhbqkCWCaerCI7aIh384X
vEl+D+H4QU5Mwmi/LJd0phMO5m1CrwKaKMqfAV+0dUpLX+UwSoBSW1Bw1pNjRTED
gkjYLIQYhDOKJKcWGsmNS+GVZsIrXhLYsyS5K0ZVGEgYYdTjuxPGUcMiXcHKTaHi
XF6aqyREDiuC5gatjc+N20t/+VChC+tm5PQ6l1HX5Fd6/NgPxxO/I5Mt8a7nsBPZ
i7kgQZsGyxORxu+gRZpE3m96EVHZIeCwIWRFgAs7e0TfIdUmzMIONBxsK+TQ5Ggm
Im+qRzb80BBBOJCR3w6++N4wrlnxX7LP6Cs+zQo74aQ0uJtZVobMKfCITIeQhTLO
thQ4LW7zn41DcdPduCNxDw/JB8wiqp0dZ2xuQcEJv7ylWY+satQ8LWPBNrn45olj
FRy4ak9fyr+/FFReQAwYYb2XeD5C4GdDh5ZU2u/w3nUv4TSU2HdEVyiZ48a9ueHo
SEI4reyk30piYNJlDoZCafjjWrs8g5HTFmeiwExYG0UVWTuQzKnfpenqjRSn0HbQ
pYvfnd7NvHEJWsd9MqU5EgZtSfaKgUyHA8klUF/Jkd8cD/6y0Rpg1s3fIwpj9FGz
3zMPcLfYJ1TScLYeHdlbhzTeFGq3eJqctWBnawgtInYMijuVhymwGGNMa7SxQcCy
wcsGyi9Hs/HCam25noFT3sw1/864SyAuIT2GmxBw9sJ/3wTs+8sGe665YkDL6tIV
IySKAnaOtZHmBt+IYHtRt2Mri22JsyJuFgJ65vHstC5bM1hthSFHikzqMbLFb3fy
eQlf6fRZ2fiecRklqgNRc1TRqAeU+In6rwIiOFJrnFPuo0BTcTVIAivKnlPywSxf
kmKcE2ZWLN75eMItgTUMZsPCnLD/7xR85vhuAo0EBJJqtpFRUoD5Yr56nAy/gCfQ
/u55c2+sEIuFHbf8YWOZ/dWGVrQ/bz9ve2JlrtYFp60T4Ay8z+CJM/cVuqKrfZTz
3mDfTJOX/y9bp2tz4qeyn1IdyjMLrpRb6oipY0zE4mNqLRxPLMZOTvItC3zbG3qO
Cg+52frm8Hw/hRCveZa6IQqPFt3Nznw4W6apbEWFZV9BuCeTxUuK/DiYGzHjZR+7
nQYt2lRqsKFCPfTaqcel/4y+EM7W86EeX5Oss8zabPm4XTVP64bD5bvtBD5XAA4A
wp7inB/w/oYUr9mtjwLBiFTy1GYbWp/7szWhenKHTWWR6ap+hrv+SWdQ51B7yMK3
UpWfE1rbuybJKTUgS6/BfleqbKidb0DfdomWo0Dc03vxz8G316sXiwXxYBWivAtV
MwlokNZj24+o/u06yAqplX0pn6RK+Ln5L2OhJkAFCelwWBiZNXnV5+JIEcxRp2Jf
Ouu+WSkmVS2uYNnWjIR8EQsXAPAP4Di47vYcjS7dIaOvbZGKtzvsFlYSAVNpty0a
5ii5WOZKqkNVeF6ME/Dv6a7OoBphtV0OvVTlFBCVEOn7Qw5l2OIgJSDJi7tSOV/O
Y3O1H192ZCj1nsJy92f/3N3rXoX0W62iQB4XW0S/6jaOWLKCMiBsx7S33hmiKU+Z
X6f2XgwDOpJ+ok6Gn9wB0A3BcZniylR0sdHJhEdqCNcMVe9eyUBdp1eThPJwNtlz
vSroylpdX5Q+C8OXFcttAWXw3V5iThE7UCRxwNmfVa5fa+UkWadO8lrePfhQKkYu
WTDNFIDytuHrcaTSS6vNNZRs/gKYGMpLMfylT3c4UCvgCkZrm9EVbHi07L0+WkkO
IBEccrNZVaEeIN611IhiXsP8jbOgfY/ASxpM9UAFvoW0fmxJbvL15TEJ0l5gLe20
thLjWLW/xKRRpOxgVnN+fYwTEX2vrgmVzUs8SuTBrZ0OcLMaZ6WiyXbz58af32Yu
qMCcY3ilQdvjzLqtXT6lUT5jdug5LtYjl1+NnnZxo1Iom02n/qaTRFyILmUlebMw
wCc87Qri0YviFpTciyRwJgCHDXNRpX15eZwPz84pWiGyGeBPZUMTMqInBaZi/rgm
6/WoDW4r6Pi7YtJY2b2db4G3uOKg5zygQLut7g+lQhpFebcwTfusEM9ZPbxUsmDn
aONaOZLNj334A2QVRvhDXuL3PRrxq0HIn7OKdNV5skx1U6fjS+GwHumrvZRDwVXJ
SKvf0ZqxP/68+pJTGFdBOL5tf2ca7MU/D0g3HL1YZSS+Zlykm8MXh3Er42EEuRgi
mAloPaQ4ep5eGxZN2M/DVTn/qxOKXo+bckdbX1CHd7xPvangPwuTp4FFfWlc+RGA
3jE4s+U1iD+oHgcaAJ9F2m8trAfX30fDEPUpHmQuaX17RTnY5XjEfIW3O2VH7HRn
41w3V6gE+F4Y8jUf7KV3zkCBuLDMC7Ye3hqtLiwbSVIAtQOVVJQofe5Q639P70F/
ZeT7J5GbdCJU/HKfL2tSwJEv7L07DIdSDQGGIG/GNkXaBPnysgXXvK4QIeAu82+v
ngUB3k3596aExdpV86/WYQX29LYaiKthF40NLNOFXzHJb5mICS+ck2c5hYUH3HsD
fwVaBO3kdrOn35+l+G8kqDNl5quLusIbp088mosFP5vJ5yvf2EeoNJ+eCqcQlVDk
RrLDQyZBUEap4TrUDboBPpaltjsSH5XyYoLxRBcChDF2iyeAiemQBzeFmVSRAanH
GIdTWrqR18ayC4BPZIwMWfFb7FyicNuLni2dNTZ9a2DiHOg4+ZphAqqHLTylq+p+
MNwou42xyXvQ6W3Fok9NsVuQ/ZN9UWTlKw1Fumybm2vlSD1TsFxuW3sAKCSch2ZQ
RfPEdPZ2RUril2Qbc6bt3UwcAVIUTIX6LbwqrG0yDN6AQW/GX78nkMJQrr/o7X8R
kJ5Fu3Zs69m3Rs88JHLDpemj6bhw5e60glRaHIm9SyKWk3MnxRcmvBDLMsBO2Rj+
6jW/gZdyS+1fCOyTxq7o0JtL4JPixA2X3ou08UisL5XISYe0a567PeGGwFRK9s9+
fjjg4cjNXt8yZfpiNLYxKdvf0LoUax3CMQh9ZyxAtJj8Ba1VB8wOr6460CGhsEut
ZDjOM5Rag0ew6fJs1OrkNq9MGsl39YAnwDkKPX2+7CKdKCxQknjNDKydgJ2n+r6H
/LkCc5rBr/ddix0BLFoTJyk6/hyEQWEsCeKjkqAYmIh6usiMJwuJUxMgTHxwdMc3
jKbk5WJ3+i8EMnQNSQs50FrEoi766YcmErf8KhTkeEPs4mRWMsCNuOtATJO8kypD
mjvczZUPyHSbzBRiro/aBPsEHVwgRuZqQV7/OFIScUTHLuPOUctZ1sQNKpYxMvrg
3j9rGSUB759DeuZfAHTL/ruSBtHeYEoNpikEfiKWsFWZKnszruq909TUzmIUl8su
PlKGwx0BrSo/wg0h6G7b29dj2fJxafA6a+eibDG6j80sf1ttcO01B2ZPJAPyaeFj
MN4GoE/Z2wjqKsViVCAvwEb/VUk0Lc3GtGwMZNT7f1y6W/dq7MXEb2n5bnX3HjAk
uXYH0PSHHWeNdI1khxa28qITYFMA2WGp3XOeumIg2M4zuXiCtiYNPEm59h4wWChm
XuhwbzMlMAUUvm6ZfN7dcR5TOegDvQXKkXpg5fE5DHrINhlBzoBFjhtyLpho+tim
ptavuNoNNf/nraS1I/8/mHiPaOD3JYfqX2t+TGb2wHpA/B0+anFcNIrjDtxsnFwR
`protect END_PROTECTED
