`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xm+HSoFb65qmx9rfXUpe57GBxKbf8/kLqfeV3im+/48IHFpIfmgwno90zbxUvMFs
O3MWINhU8bI9thBLrJnwZPGpxH/8IKnt/hHI13PKoAtDx52hsxsvGehD2TLdpK2Y
hrRXLSxxpoE3HooYZjYraHxbpUvZ08t/JpaVrNYjJVJ55Q/29J5bHxYpnzMgGkWR
Y5SrouYYANsyk2EqM90WyuyESOF934dzJ9GhTfgki2yYR49ar+VU4WLLFCdFhN3Z
O13eqmWPNRhO7VY13irTjVYGsHBiUuS0/j7C5qFNbTdhZ6OajbJ9jocEJnDIWQhY
0wI7rge9xiWI6+b8AT8kOomBG9jhNbYjwneCQpWJt7SyDNEq9nLvlsT2HheXdacS
`protect END_PROTECTED
