`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AaKf3z3Yz8TWPuB0tnVz3BCHCwAWDOfIPN9fKLwhjJyFkcAcc4StAGosrx6/cjrt
h2unhgvYMV+PJ4iX4zzMd8Ce6N0I6DzPFs8J6WUHHNqxnyyOn9Tnb/peV1hjzWaa
LgvMZOim7fw5Zg1fT6mE8yRa5b2kNyXKy3WZd2UXFonAZzN6BjJCnR/9Sb6I3ima
tEecImMlPazZAx9P7Wkc3E5+VQoTaU8LfcJmA3Cp7q3eq9KAdPW9wVCQm5/HUcmd
SDxcNOjQPp2pq1sXYy7Nl0iyQuG0CtG9+uGd9j1F62i8aq3oQ65GPAokDMdXEbUZ
WPGKXpaMzQDDwU4RF+l6jQ316+CsybH9JQNYcm864xFx4kX/Wvn6HYcJvLXf6rxf
s5ZAyd4d7FGzZD5+YU1TN9LaKiQ/6g/q7I/Ee1kORkRrlzzVOLORBEYdsTant+aF
Cnnkr2tT63f+q1K20BBZa+/sRaJB0O6vfyKlBkdcb72s6N5C1C5p+ziUuht9mlEN
`protect END_PROTECTED
