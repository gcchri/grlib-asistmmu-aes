`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RzxEFjoH38pE/anDviyhgFZP+3VKP+lMbu8QBNcHEptOUTrQBhkmHDi33/rZZksS
dwS9QMl7OS3mBg9nxMDNu636Sf0G+X7sjxqCMKwr9Ij8/vmqR+bi3g1rlJYGqm+/
uTNp3Gmr3IB1GrsQs9T4pwPOz45Uingmj2mzWy/p6wJLFNH4fQNFS+I70NqRbiaY
ZhIgnilD3WRnrmHuN3l9Ey6XuEsHjjCAW7OhGWyXzwoxxLIpDSNcOR+kpJY/qJ1f
wrVgBlpj4KMvyWSqGk1AJu++ev12lh6Ddczt8ukQq8tfwhHYDkd3VabnNgV6a+OP
hb+A8Pxi++AGPxkgQtQGqIcwZjUVH9CGcT7Nrdf6EVG7jNwdj1uVnwwgjKA9bA55
52U6Tt06H91BTUxdbKIupHeKj2TobSMQn22uUquDpxd0hyi1FruIE7A8XBRp3KIx
nP/kUspFhlpGzUJ+QknZLNgP2kobqJhxAxZFM+Tw321wVjHoTq4RdR7dGYijCXfa
GH+EkfdNfCSLuPUuvBVA8GC4NUi8qdytR+i4223adawIqQBQzeGcEoGpeWQbBO55
/1HvHd8Bnn3RH4Kx5DZq3Ures2/MEXDD+BhgZ7lu/k398d6SSm/LmHqxb0jfSAOb
VP3WYvMMWgTqe1chkewiyzK6mcbwnB/mL5JkUEk1bO/iQ/TzwRDr7vfpw82UWMO3
FL9Jnjuc+uB+Wfr0ZwK7LESv5fQBqmTygSj5i1nniAWr/gVczeNN8Td3yKjvPmtZ
kauUkLAZE27Ba/axstVvnK7/L/OTMvPljQGHvrJW2Eg=
`protect END_PROTECTED
