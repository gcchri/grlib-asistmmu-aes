`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6q8QSztvgTswZhd8W9X9p/T9/en3E0kbdi8E8eWtpxuEJxhQObOUyU0OQFTE1Bpm
XleIsyiCwr29pC36UoAwymWe2KaG0IYtCswbLmyuvfrMHv9XRhNptVALEs2S1HY8
iT827fGl/Vg57VzXjpWoJ5tCJFsCTeTrH+Lv/kOako6fYEL/Uika1IgMMlzlEtF9
KqPASNw6gS6gQREsLvUVh5XB3z9CAZ0Ph9SNmbRQpJIuXGdUje8eCTa/Y0+VL/hE
qORISlnw1x4o2D6WY/MfkI+Vp9MV1U1EaQjjIfrlrQ9sHrNSVlyoNiLtcmdBOpU1
RxAmwDczEghMCpvouQEgSGVPaRMzIbuhwSLybddq5rxuKOdmh6kZpg07nKM2SWyM
k1asEuHq1cyi80c1tOaS3BPuGRf55/AtTjxxr3nJ963aXmC7SaYSCZ36mAjjrQ2y
Jo1xYiKlxWkazaz1eu1xs/uwbBIlvVnUuP/wMLnDz8U=
`protect END_PROTECTED
