`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Y45h+o9pjHUM8UE8rVLKoAoxh1qxMned5zyRPsHQeoBYqcvELnrF0g7aEWra8Qb
uLVClJp5iFLm4yNsgpBj4CovOXj60ZzMQEezESLmyoOYHOOaFh1rQ0gQt3gQ2rmT
aivZH1wc+UFWlyEezWutTVhj1EEwWLzrLsvtd4VQ28fuklH7VfNQ+uQw/8ROOwJh
+oCZRqsxbfaCcLXeYv72DuPhx0RploeOcw4raeIMPUiwttekZDxbifU7Eg1oF25z
6euefObAPX21BXMfCxI0F0NEuSSG/zfZtAFAdrFeIQmFUG0MaRvauIAIf5VaRwnj
b9wRigRxlC1SexieiV7dU6v6YOC1FaeLbe4mJDTkrnrtQgdrCoUJhvLvnKiZRGoa
A7tgbbKz8Tz29eIFnEQbSP7PigYHlA1VbAA9GBMyi6CZ1jMt4OaJpwCEIwxIjUwG
BUxrR4KEGSZEf6ezqFtpzVvGnHjtLIAflLYR5w9VCY0=
`protect END_PROTECTED
