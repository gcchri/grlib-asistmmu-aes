`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
owq23l5rusanqEOB5XpWdrQrSxtn5UkVH/pOB3ZPvzdAj9hxp+rkAenEGPVSRXsS
EJSdugf2qWeym8krDnQqiaYGEgvAvZx46zn2jangsFXSHrMHhBx8bV2DCK+6B7w4
W4SE6J1iC8tSB5xXqGXksvJU0pBJ7CFt0qDToLqp2HSwQ+xF59GV6FLfvdckow2K
q7/26lyEB32IQdsQTc4Q12BK6Yc6nIcPG3dwL0L63/EDZ9FPZoxeRXqUnrwKsMR5
vqSkIonPgh4BfDxasLkAaBDQEcGovd7szgcmRz+RkOUeZUVs41tYm4oHncZcNlHL
3AJfeCkG4TUpfaMY5B4SGjFc/+iIn8p/nIBd9VohAbofkf1r+YZPsQwCLu2ngEol
Js7hDBFZW2q7g0NgCbUG+QHkuwFaWuOQR0hgKnuOlHgypv2+pN0qsgrKpcQKxlkl
ypva/QqHC/T24xsNFRl2dTcWheUptJQn3JleITR5gV24WlDp8AAjzq3DYc35lHf3
UM97r7t5s/CmyCgTn+557Dhu2W6VMGo7DP2FzYnSpdLng5CL6tG2aSUjDBvBAc4q
X8BjBeGZ8Of4DHPA2iD4tU1pZ0eHeX00vfwrUtWPVKADUnZBc4+cnrCkpSIzA+TU
OaS5EHJU7jMQzpbEDKhUKTHDs98uY+r/YCXVGtuupsWSP5JBrmoqT/CmMwD8Kjdh
2XVAf1ezg1Ga/MVMb/XBvPbttnlmOHqJhUsMFRG/CaGrqNWE7hsi36gjNKkHeD+Z
MjUVhcPaD8IjPIg89/FgWWzMrmwxU8xLR1Hg4CbK47S+eU/SkqVYc1npMO/HREg1
jf9SEP3T8PZbCIoLvKtz44B0F99xZojoBPlr7yJdfAL11RZFOKp83Rk/dCP4FNdg
qHl19sS0CVQS3yPIFWmlo9zKUjzdkYMEa8lklSss1HGDesuUtBpoVvaEb0acJpNY
dUw347QWdM6fCVzT6uZF4UDKWoxtc1OYC3D0foRcm8iz74JFAGd1oczYMaseDmzq
h9tSJK4BJC/QgsNijdVq8RQZJlHHKA4Ycje35jyFOcOPlNZXf5+OqJUyKpqtekoD
fOW+RYxg0VuE8wK0aDQLUQ9SPqnUCDu8qHb/r/Tfx4ozeUkj+RcECiOiOP+Oh7PE
4VpzKEvHITXbP4i/CpYNb4/s8Pfr+SVha4urzkro0a09Qluy9Dcbb2c8F0vKt0yU
aFqj75f+jlxORPKRGznOe0nFyAB19AowRU32SUhm1VICO89yHy5n2I5BEiCwXD/n
RLuDI6Vbrpno1/Q33r7z2oRHiBwQ84C6pUiQVPCuQGpb2w9kUjm3hT4I8Z+jiTiB
dNO9eScNqMW9UD9Ls+AXdoR8X+o193JcFA4U/W24i++0lnnXHRVyWy6GuWD5SA6e
6ZT63wlaYZrR05gZQ+XQ4dOZM6xLAu+XoWw1+TCxJa+kfkZBeZC7S0TtrkH8q6gl
AYNSsvzw44WKzYGYklRHhqFuTi5tCfxwyoph1xcGJTsRd2wrlcApWXxXAJzndhDP
ToFJ+cYF7urtVamjawOkAUps5CHSGP4aB+iQGnEeikD0IzmztkYg0Jlbz5w33G82
7YiXlzg3NT+iK45vRfdF7mn09agnZ7PY+6PBPdIF8mEsxAyd+NuNqQjzMWErhHfe
ysnwiegxEtnAMnk3aAVVykXf56fH/mze3FWV0UUaRPVNQmZrURJSOx5Rq3KemRAp
mqX/y8H9ShmFZ01QKh42BzD5fTUo8PfQsJD355pv0anEA1UVW4Sjlwv0ErAy6RXp
QLY+OcTkej62LUvo6fAl3J195QrRc5ju8iK0KkyKnI4dJWW+78vlicBQIJbOYvD/
bQL+3gvryIaj6PUkg6ltyfKWU8zVve5MWCWJCiXQzEiXQ24VR1pIYl9HqXi6hyti
wILME5hpiL2/4FWWJiqwRpCloE7Eb9E4zEKxgUF4DX1thJOdAtOG1rGdgd8HSJ22
sQBi/Nq2Hsas+siAGoZ7SOB3tp7gon2KiMhZGpQQkajY3g1pLIGu06u/KSFtFimG
6jAlJEbQgSgO1lx0LxavFntcQW/zZmbiSVCeRM9444x2FK7ObKZ7oIt3Gm5sH/Dl
IuCq3O0v/TXQIQQEZwt5bCD1wtjWJHlDMQ+3j9br9VAzbzi9zLfDnDugno2Zh7Yg
y7td5cmHr/UsjqF5OJdgSdFLZ7QfSEyDX1tgqlYpJc9S24UBGDywMFKkOI/TUn3n
z+5Sjh/qVqZMoMPp9MpZe3LM+FSWi9TXCe+Au4gC+KoZZylfeZpq5al0CyXyDfwA
RTSfOsytkY8+ZozWpbSQv+AvxUDmjRsqx89tYr4WT9WdoQVhKzdrsFbrPHmR/ENI
zqL3fBT7oINlvS9gtaJSWd0ThlvKAFTNV2DaDcDEawtuXVcKLqyVM7RyNMOg7h8Q
n5Q5JRfy4p4Xd/rQLOE9E15d+QlxIKh86CbS7WwH/6TaTwCtuOrnCfE2nC4GWxwS
z4SN3J00Pd3wuU1Lb/0eIYtz2b224MFmJVwJd1C4fWc=
`protect END_PROTECTED
