`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DseDO1atVTqGqA3e4OjkA9OUWhXYgS5efbxlmq3zIJ6X5lIUG5olnXrINgOAGSxH
EvfYZR5nAVBWqX1aC6QwIqg0cr3ZWPQ3rvwWMhbGqbvTCwe1U/bb5DB5WvtWSx8A
KlqwXoU8Wcg2ihWHw1+ohDEBgNDDfLkfx0cawl6QeLfxt6ZmR7lFusLQ0X73EH76
rQz639/x6SyCZYZtcTZzIATa/wq5O1teoH51h7FEok2hDfV681pLOj+Z/z6A5mNe
cnfAT66apE4XqXtQE4rDOT9jq1Nw+lBNRFNodehu+PZn2fB2gXtYmAZ6s4GBvXZw
ZWqhgoGDj0ER3rVy0g8CDOfm/LKYsfInkSaMPGRJ9BzGzeOF8YRgX5k8aJL5902D
83mOrFvQAwosDPL6DeJaDPHCSUXbb1M1LryPaiPLLGG/CVeHgzoVrSjNE9DXUfIn
orNwkRWY1oQo9ZhHxUCsROQKBK4Y72uiwSkk+QBIPaAvh2Ac41QG8M+14dWzWoxG
pI50d5BWFnYZA7htSCYPD6131cL8j9CN7nmDGYwGN2LKp52CbeFOOnB5Y3tZzCkS
HMwr4CGZoEymKvGb4MImK4zCqwvea+KTd6cnfNjKWixUDUcQYMJ8K+5DnCAUHk+F
CpWZQckmPAVbn3q7tsfHHnld+5Lgtn1lHUdz+VTT+Ogfeg2GE1j8nSx8B1CbjIe0
fGH1qF6H+mHhB7WQLyKW4fOXiU14tY9nR9EO6qsdWQXuOUAf4k9rtPkvytelP1lG
QQiF9fB+DlQ//YhO/6+RAdzezS41yJ/Dj0tyqVcwRP2vXtNqCEIO0WjQtbAWjgQJ
KLS/hF5Vt6iSCfIvPv89xSUF4ldAsody4O1H8/AVTEeU/3ChkgDbm7ThPwzE3f6q
qNXIZIF8fk5PQth9jt5zokfgp62CATJzmiAP9PQH9ywlxXtvbqRRcrlCL0g1fHgk
qieAF3t5GJ61NUpAkHFFuO+abLS4Y37V/al0+qOCH0ThjKZP9Sbq/cC6bJRcxwKK
6gipKVxLIQi8hFIOFgIxUC91Qj15e5XynwJS7TQwc7BiiijYRb8/BTuYgY8Uaxrb
QISOOMqogozLp54IbQfh8gJ0JLOqRDm6JzHH7n38FT9/4WvlF/hYZQx7j02CZ2UC
rZwZP7FHw0JjGD6/+gTlnYSDbkbZ0pQnEsgUnAF1uSolbgK8WlB8EzZoACsKmdk3
lI01vtHkMIpNJg74SWYqmnE/L6y3lpMPQvgq6QxUSquhMFxitTtz/7gLkgaoLACf
iOdS0BOCzo/IYjM8X0Mje0jF8AlqOsHodg0s/jn/ozJyXafsT/3e0A12cCrhwvlY
tU42t6V7GI6k1SCmQhDwxQ==
`protect END_PROTECTED
