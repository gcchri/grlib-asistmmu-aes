`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cVnlEGO0a2qLYIDjT6rLbTVlVWA7YDDAVxgdCIJPtYbcm2Kaa5gjGOVaF/66jvYL
0epo8GSWaQEBCgsUl9fH/meGMw+NZ+05WUQg2B13UCdrsqYoQunJ8yseTpdXYe8/
zePveQy9E6ATWqnXUL3AwRZQHZHohaIND2v7MZY+nrRF1YD33W3yxVWmKzlTBxX1
p5/VV0e2NQ0cw3uu8bofkH6Y8GS4u6qiNRUISrHKN/Vjd0udm9gI2Zl/iZsra8YE
i1qu1H0mqfzFByafoOS2dtefmTIu6yYuh+nJlkjKId3DV+CblxbHH3RLap4qgxhh
`protect END_PROTECTED
