`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MqzLWkk06zHhj+LfoRvCEj7wu3e/WlHgIWTZa5MqfsgCuSKyVrOWtgDHNFpvy6qn
LXhLnoF8weYbOUCBPWXkuq2WUg6rEDIKmeFHoX4K3cd9Gl69RZH42D9M7+ldhm7h
kBIQqrfsNovDk6yeLkeEIqzzRcAKpXe+yVnS39Ji21L71LdxQ6eUNB2PIz/cku+B
+/zCFCboIgKdC9MU2NawNl5dSr16YtThq6234cepL2EvPhh2lXOIZBcBXYwWbqs4
EEIaDyC31qP3uA4HCyz2VSrbeChFLPsb+Xc83G+p37ItjvsrH3+XbKVJbYE8MZpV
j2/K9PdoLIhVwK6jlZS0Q1Ngjm9MTPOlL2Sfv/YuUq0yzIhUC6gR0V2iIVptK1wo
6AudwkTX7LztwGH26sF5li3hzk3e0TUKET1FpZfb+YxJLsjpve05bYV8icRMXeBe
4m7/lQcMPAak+k/KV3o7Uznn0GwYoZRjnLrjwOgZWdE9yLKB/lYyb25V4eSlQtXK
LhwokFCgvPe+fLsPQYLteF9FibKPebf/VFvABHkg9niLNQgo8XFcwYklJLzj4gie
g+EoGefLSgIQMy0eEZQj6w==
`protect END_PROTECTED
