`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H5oxil/gSKueB4uFW39rblw5jbCaTGEpRGzZo7uWi272shr+1H11GceF7FOSVwXL
u7qlr0yAd74K95TiWzQp1iVrCTn4GqotVv7Vq//6cXLaogeZyMHeC3FmsZlRuvAr
LaP+4/CbI5awVHdvwk2UG9p+8kOsTD1/gmdoBpu4cq9cdzjZXLUGF9cXpYLxmKOt
58LCBIOisi353jeVlJgL0XvgCDHaQ0/eJ7hXcexy9083Bl7gXcEUm7qTXVH14dCy
O5op/eHlpDXUDQ1WEEgegDe4r8kQmF4gzdCtqjcHcxn70asFA9n9nF51dIz8fwT+
JDrzas83kxSUMZ1rI4MXaqZPSgXbtyAhV+CkV/Kon3jFbGzRN0N5jVPNbhP8E6Zr
1jmYrSpWCo9MHU5Eca3h1kURlctdCFdXSTiTcnoiRhY+EP1JwItYtvjzZNVDIgYa
RLnyhyv0QOCB+THMzFwR93OkqHxBUJk6yvJRz6fOWsK6rlUoAleDGHRmzUN+EXvu
9fDCCRcSyvT/NLK96YRw+85ZFuCbROSeZYh4hywZcu1KlHYGEWcseF/eatQkKZNc
/1yNO67Bm11trk4FWtYratUqCpS3hwLzDDyXQn1jzk+RVDPwu2DqoYwmRaRc2IPn
R7vOWUk//pp30dptN25Fn6NgvYdRsb+HrJ0JbdEcVIP6fU9MO6eMS6s9UH/laLeP
XHqDR0ahd+mgBO2YtCpUhOc2dpMvpApjHI/+QtEn8mFnSsx2JeiI91fPIpUYjFhJ
SxrTqvqDq7z0KrKoXIOZWU7U/rk+QJLy5FOJk0lbLDCrgAPg8l2t7kLSAfbhcd/V
DWvVcVuwJBMAW4Y64HqOSJJg8Gn/CM9equIJu+iZOo1far5fRLgljddmCMPu/BCM
ned1tKXp+QmoCSCP4gGDqLIlMmgF0jhz9xR1ObgJZ6BvL/mh3cO8viI/PBs5m7pp
AmGQdUG7nL20yRi6nQwogyfwJgkBsgayKQiKsyGlekikx1y8h2+JQ/q2qtgbsvc3
tz1/uwIaB4u83/FK0cJyIeawwdosZPpSrF4v/eac9xWJ+LIy7mS+xhzkUohk+hHW
9JRk7Uz7bPxFOfLbpuXlEL180+w3qo7Ed1jhbpl4sVsofC9LCiGtUI8JTdivmPez
kmzqFBubAUyhHo6lD6cA81KjyGyOmtwwYV2itB4DLD7pbixX2fxb2yb3ZgBEanD0
70+PHZleZ3P/3mpVjI6Zm388N4GGfQz4MIg/MH0JL7EBLiCEPBiUZFMRtFBrrrrC
aC9A7bqhjxfRbN4XfpmKz8KiSNsL9CUc+8/S3VVrYReyei7k9sCvWZtXM/LAYCHR
O+drN68Jk1bH1fFZdaICGJvAYVqfLmPye+HXJXZjUPdI3TDeIJ4Vl7Uk6ZyHdvYF
WcWy23t2eZUN5IihDURqwQz+/d9K7sCnM5r4crrFTUiqYCqzWXVm95HJ11G9ewsB
Yo8XHzmrqUNv+4WNCoxfA7oc5zswpYSfsQldoGY3SI2q03tZPn74xzJneHtkoYof
wn/HO6SM204PpghQwI7dstKRTXLfdi6UPZAr6aUvvKAg5X6/6u1KUgHUTpCTvqPA
coP4NmqygUK8YBS7WuKulRWlKSjlFBEV3Bu3IwSnDExbtCxBKR3HVhe/5u07TTmD
0gHyx4D72Dk/8cmm7udGMezTG4N8djOhlvetQM+VDgOWYqygZt0TiwIC1D7Z4Vuu
CEvLCKbPYQkjMJy7AZIRbsWzKQHrjRl5FgxXjSqWd1iVyOFYerrRWw3fnLZrwcc4
L7ad2FV838GQ+QRkn2L8tg5B9XqFI5F6uKgI/9EEZ16nu/v5c8Nubmj6H6G7GYXT
D1FaCRJRLmk5xElg0yyH0iH/leiLmeS64Mo7svoAtiOVxhO2lUH6OXWR5QtIBRYK
3QrgNjLCvzJlPh67Hg57XgNoxXRsjItMqzOcOuhCmv6OW1sBBQf3/ukB5I8LhWjB
MU9eIPZrbjeJmVFovE/E+Gf0itgKsD3bZjSV5Npnk9iem86fmICLkoW2aSdWkPLC
P3gTIdmD5G1AidVL13CRWWA1aMA41lFz93e4YkEMnAi9C43kPtaEt6xivbly+qrU
ukHauXozVJNR9B8ZztcgeRV6Ja8eGWDPU4epZex8CMQ6V8flP2dPxqJezWi1RLoG
Pod3W0xzx7o0He32vBGWpiACOhRwdf6MBEPCVItI4/kfeZo2Qs0gGyrrmqNDcO0M
qvfS0c9F+mLVMz6JoQm5sbEox8ZngveSy3AsdNXihfhdU4OaNQq69lBmjSb9zfsD
fLoqlnzFoWJ3F2b+ZV5JfEHHyv7yk/46vZFcWxHaa5ZOqUEFob372rRdWlOOY+LU
D4dHFf1rfP63jml/SeBHoTm+fITGkhUU6fvZ10hcwtimD08NkUsRz37oEHDryv5V
ZOrwoEg/RuW03ntJbPYjBjra+Afjp2knzh0ed3HYhYZ3hLSYVkPOCHoSqnSWw4zL
esRfosLFtioC/RNrt/aLAsuI0Ziz1EuYMQ52JP8QqqgHx4dr9HRtoIGutYvm6nbq
+rw9pT2+LqfHY9LqadESNtEp6NdOe8OljSOwMIynPsUf3gkVWpWfbNpRSYG2FOAK
35cmJNoLIrMZTK5GG6lSFLqaRbE35sKtPCo0qKguNJDPAgHwYwwcX5+D265ELDSc
H/Ea2gZ6R3jESp0nmSTh7hdn1Kg/oF90t9g5BlgYhMMg2/D2J3xs8IDA5s/zvdOF
dRzX5fLXOKCQ0Z4mTd2R0Jnvut3RmiPq8qlm1Rxz5gMDOv7awBdNU9NYS3c7nxvB
QA8pGFDbpdDgWmVV9KZJzzjT+KIZR/zau3WqBxTS95j6/hZCuSMx1s+ZvAnGjuOS
dS7LyKgTrM4l9WXDPz91YvH3FI5F+BwgWSbO3eRrtDoeX57tI1s1IO8jSTE9Lxso
/Bb2skfuMa2pMD0qrqw2PaDUNauxZh8YJhCLhCO2UQyihiIbVU493WtV1ByBTc6M
jSt5tSxs45AisoQdg0fQKUA5CaLBSlp00VmZnvz30eRvOYXivs4+vjKlh91FpLIk
TcA4b9uNPghCuiFf6K4wQeNkNOzLuLebp7RJrOuInfZKOl+nEsnNXjcapkW2pYT4
ICtE6VsGlerJpJAMAOIfvKWII0Uk3s4nrZjklNv+oqh6+0t6+V8NxLsl2cxsNwvi
peUb3C45qRuMMZPbwyS/0qxz+mEDy+cPD6DVOYaA6gpHU/BqWERcLvFyNqSETqEu
M6qMSJeiiOZ3Mxka7flHCcQzcDXd2dBXd+e+pavSC554RTOhFFUH3iiHcQQ6svtf
K6DDJvTvBSWLFjEmY1DfWOkv5hfJJVart7+JNmI5XcEcrJ4AW0PkH8T2WU2SY5DX
Zc4FC4puk3Qvsgf3LpIijHA8LomX4NUb5UibWGMsDe/ZzWnbfNoHhVumuIZ0SSWx
R6p4SgiAobN22TtrFVbrHXbGcZPf5ecVwz1iObzwOfI6DTxXyuvqn1aJCZ8xhw12
W9cXzyJbQbINaQLJxOfbyUxMKwRb0/7DpcpS9yvwEef5tKn2fdjxFA296zHAUGSq
Emekiabx1GAIpNs3Qwk6Ju+ZP41xtIWh+hpq+ZA1ILKi5bv/gTSJ41GnvhUPoeMk
v5G44pMcP/Ux1qTomyhMr2aIBGYQ/UEz7WhdB2qhPsClwHXEuy/2mm7K/5IAhulf
Qccrvvbc2ffwGAMTW9FEES1i0gf8HZL2o2fNCcsCw97FqHdkcjLG9tOk/btbYD7g
eA1HbY0xtnj72F0zjkXjdZzvRS2t18+dOY1muquXQ+bO4GKdR9YRHEhlFdaZM3xY
8tAwwLV1FPV8OdIEZmfCB1AX5N0m+6PbiqbCmz3ytt/2bwebTjCvweXIh+HvzCu3
fsEZ47g72opnS6UueW/B4H+sdLR3TrHoUoJ9N1ffuIVWPHH/xATkUpQsBEqkz0uH
N2Ut6snCmqsZ/1BofeUNmc6nzpBqx89wTKRNDjHek/8DFMj+c4zDBeCLHYLkH6Qb
QGGNYWCu2J3Sj9hGa20n0bSUb3cj/3nbDZ6mvhdfSAqcCyttC6eB7E296dTMHn6T
BmoqhvMVxva81rtFb/WBvhwSNOm/esH1ag9mUuF4pgB9m6ZMbEGOd1o3t3qt5EwF
f9B0FqayASKBO4leQ/Mq98UTqOLp/JBPS0n6pOXoO3Vh5RV7GemIiJB5of5AeivF
b1jTdt7LYOmgYvzQrfvziYJsKdwCSeKpVgdSQBuVA8e0V0DdU9F4YIa5B1Gy1CFh
B2iR7nx1Ii7HZaYEPW0wvCSE3ixVctVLeGDoV2R7Oc0OUbcVLKDgR5XJJJxi7HTm
gUzakVuNIa/m/DNe5LOcROwxiO20UxNFvF8jcVRu/sFyiKX68G5iu9jjAfc3Vv2H
2zVM191JRFhpqs5TKST43regMBux2klfVn7UCdXBXOf2F91neiD2iT+h21ij7KiL
XZ6iehOJutQepqfdx81kyoobR9dGgIL+1+jNsQ/aulKL7ST03Z3hJiK68hzriGZW
kkqh09qtTzpRWNHt6v9MLT9ylKrvYYdW1So4IoWDfQr9NqPVxWX2L85ESj9NfUSj
jFLyQIcnf/HN/VSb3OqD+R8sVJNOontT0y+JyK1qkpQZY6/cVAPuLC6ytSh45icJ
qMSC0akmBOxyBwpNkZlidsuuSvwG3LjKbtyoN8FO2tPLfAJ7AaASoZHzDEDKWqzP
8XBTV3YKTWv6FZqqpLvHv6l2iBDFin3JR6zj6/7vaqnUwlqvZ/3WLSm6UsFhP0Tt
e71ENMnChPl8JLKd3ccKziejXaBfm10DqlZNhQBdJ2jqzUEQRQYnAAXxkI8iHCW6
ASf45wEBe7PITr9fBC323UyTSPnh+ZabLrodi/6mz6M3vR9Rs1Q7yfAUhCcmlDRV
k2rocCOVO2R5WL1kVyoQMjDnuG91ATdCJ9//zro7BPscweQuawJbJP7dk1Ut8F3V
kpx38Mhm11PC7eO2NjsT/HfJSILFZ6OMm76TveorfPa/+7RXyhfJwElCrSnM4qnj
W45G53Z6xnNy4Ul6rCGB5KMg57krBElBLwDSKUt9Enm4nWn7ZJKiGbj9oBciq9Ha
Xf4WA8y0PsxoOcNREc6S7QggJEBXDeLu6T4Scib7YDvO9lMhNnJ3rV/AYTv9jzYb
yodOp45yHKiqF5qPVAMa6micNIkS2hTufckLyqDsBM3PAIRbpK06PDqYVicrAsFI
vixzMRCz83Fa+6POBYowICOffPGWrZTfvvRtmuDAJPPT90Z4+Ed/cJPsA4cCnr+M
MuiemCajn23t4BdoeaRbllnMimktcdFp1wahOAff+Pc2g5FIo3GL6PBXHLue+Oib
g+eUZIRvUuS906C5X277QH3C5UVqrMrWvZHdYPTUdRqR6nTLDFAYv95JIiQvbYXs
pRZ0zfgrs4C0gKM8bq/6sKDCwOReBjrUqof+gPNVt/QU5hq1bW0HxHRZj0mXvtNo
tXOj0woufoYr4CKIKKFVeiqFQozZ57mJPozXZCvc53RZwL3LfdFEY9hvfri6W3WN
eW+5fNX/F9TM0iHrPCEFcEYu7uMv5t/Y/S/UQ1fkP7GAmN8fygyr7OTndyru69yw
4yyliR/OfNqCZH0Q03H1Qi+lYH59GxSHy/8kp8xQvyt41yJiALsYH27nElokMD91
vRV+ZMMoPKttjR2sIcEjpWg9B3+86SHVZxrz7KwrJtnYLEiAkm2N6YWb3TP2ufe/
VWPRL7w7DKR+MUENZaxBLifXclhlAVXTynMQKc2F4ToJJPwkJyz/Q7ySQZHtZFgl
HPs/14y3Bx8FZ0sEi3v3CNL3owbt669uzNrOvjpAs7w08/XicwKzPOm+p/kk24W9
K9oR2f9mTuk5RkWEOi9K1N1cNJf6BV8hvY02PdZfPOaKn5goTaKQq0wTOxuEd4Cv
zFN34b7alCYut1ZR6cnlrdWY+2hfaxyw9m9PY133Jz52EkjGdnXXgjS2L4U0igBY
wENExSFL9WW1v4Ovr8zd12mwJXdw/i84DA2XrYyxA9OGwd58/80+cp/ACHFKES2A
cP8E2oxDpwZncv/VrcpRhjdaFYi03S/m6ZQeiNSw5rRVsCIFYEl8sp3ekxmTrLW/
cc56m9tG6Zx4W9GP8Q6s0Qrsw6XLgQQ4dnwl4C2YhnB3EEaWjAbhDgia8d8iXcqG
btEeeefumzK0IF6rOasB3PWUE9y082Gz1fQZnUASBN9cSHrYDsgn9Gz19Eirxzwt
2+WaqmC4AeNm7opgUOAhkmmXWr+xL8xh5VwQC7bWEl0ZDk7Er79ViYg9OrmO6XHp
GQt2ifahUsojZy0mOeFwTDAzEVSRyDiDrzYIOyEank6tzRIXoJItVN7ll6AS7+T8
g1sz0HOrNz1v7s2rB7Lx6Z6vM3o8BJVvZUnNquyoy9fcRNVg5/RnB3pS/4qUU2g6
m6zmeJmT5+saXIQhpRsomo+VW+H9qRJix5WVo9XsERu6RFk9Q4RLmZhDy4SlcS8v
qxFussxEMFIIowhd896hEJ/brUESvbpMlD8x+IP0T0pM3ElQj1Ze1+BkBrtf2AXM
icNUy71eNGsgcyz+IhuKqHYgzI+p0pTGtMMARY+t/ujrt2P03gtqsFcJQIzOsro+
VQcPqHuAttbdRAe2yCRId9C+Op04+pdv3uv2FgBfLPlGWbLNuCRd8CiMM2qtPcca
RVu+dRVXkIoiJnKGX7vH8A==
`protect END_PROTECTED
