`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Er6gD0CLT27hc/wsRteNNtYADEIP9WhQi61GnA2bXFiYSWZy2c+ZVNVqCoUEwQAd
X4aKcgQBoPu4FtS5hGCE/9T48Be4Ii3+GnS+cLpc+I/ecQb7mX4YyuOERaquDdSe
ZZLIIP0dkA0Nk8+1fZNve4vWg38cIW+3BzQ44U/0+e7kkplX7mGg8VdWJzWsYYOQ
zoLMQ/ELnDWICb67ZSb0l9y9eMlfJY80DHv20itQjYbdXMsY5RBDgfsv0qGuD8y0
8fMP27vH15aHMldiq/8DlIOaGYPX2hFfJ6FXVQZXbtNeTePrcswK922OHR64zkdA
zaXSszE75epUlIaRteuCsyc5vTREzivztNDj6vySLGDEEMT3MazxFfeRgwxuxjTY
VaLpoycOroO8dfA8DAn7PA==
`protect END_PROTECTED
