`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XKJrj0novwVzWd2tKBOanl8Gf6YqISbWR81ClAP+9/v9Hab7xC/Wsc5dMfF0cAZ1
Nx2spQ4nsJl0hTs+wlaTY4OkbJUyQfTjy6uy9FuSZJeAGtm9X8xzrbznI2Tvd+Zu
3WTaVLusscK2cii04BZm8G7RLn2M2Vd6YvbO/NRQ+n4=
`protect END_PROTECTED
