`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g/bYACA2YuYPZp/B6U+6/zfAT1lLGWjQiD5w2Wk0g6ls2JtytxQOMRYYAr5RvRHP
q1NWIhQsRSXg0bOXu2J2mzlx+uLQQILdKLvzhF5N1vLvoI/zP3UcV+dFtA7+D97Y
GuhFjvlzo9s8zg5hR2f6JolcN6r+S5SBc6NKjH16D2U0Kd/tKwTL9StNT2tkC83o
xLSdi5wu5V2WLwcCBuQ/O9kWxvBNhZKnEM5QuqHOsx4NgJ4i6VnMFxzs88FPMLvg
3Xe4+1Nch55AHjkRaHDrFZ9hAno46YCchp0FXozRnYP/plzb7z5X8j7IYNHq0dpx
PGWEdb7UVKLAaZs+V741rBF6HPQUC+hY7faYW1QZyu6q+kmvKUGbQ4HW7gcn+FWZ
UeZXM4k8hKNitLvnvY+teCnOrW5jNTMwllMoD8RmfZSiqNFuqHwI3E6H+WrpokAf
gnJx5M5kwHztG+UTVNc1Q3CAUJ00sxqjHYUpOAITvlz/XVERortvjsTl+S4GJxth
TnxZ79nupcDW5XULOz2t0bgmBLYQqofZME24cPL1NSmP2wIX3uT+ni78qj6I5Kpj
ps4Pbb72od0yk9Wy6zbYiCr07SYPDjx+WOUUlCDCyxivVsEWRGkYoQWEypkP5Zhu
UcxoPGdzZK6GLS+FQbYOMZMTlScXz1WnnIyNPKDJjUyHPcUqYKVUB10V9VAoXtG0
U1Oj+vlG8ktqX7iE7XOMe1LKWxOdQY2buIDvZ4EsqnGfyDtAnZBwZkA2H78gM7q0
JxddpY6dAlNRR6NkiYLSDVt/l+et9sf4R5wJquawREAERprZYFPqdh/51Bio76f2
sCcwfPjetRRJcWFipsjMKgP5d77ewN9G25zYZAHoQvJK/cbabkEJzBRCoPrqXDrP
e/6rPubge123ZVmizcDmsK3wrxVOxKjUrvBwYoKNZ10=
`protect END_PROTECTED
