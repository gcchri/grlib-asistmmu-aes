`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DTSBLbgXa3pDHlZRNEna5e8/Frva8CkTzLkTdkFrmhKrhiK+vPgkUTXoZLQ1mqZX
TK4MabEnABl09YBVdLGyOGGCS0Fnv5byBqs/w2c+ij7gEsmOUnXHgT6RRuCimeWC
DXgA1baw2tRwQWfI1CXF6Ifghsa9FyvMVmZxlxZegi4MkNzA6CmzhzXB0IImbZvS
vaD2vXtqRNkIjh+un0u6IAmFfyvHqWRWAoSMcqqs+I0YE3j/Cm3mXkF5c2OlRqJa
eEoKC/cmtp2AGeaPejo6WxyQ0+RloQUkpgJf/6uhJl5GtFh0R9HoYyoGNa60XmAu
uopf7IoWdOhQNLFSE9RTRLNXHBqJ4sQDizxVOGDAq8MR1xiRmeOrHrosQu+dOMBL
PHyomYzT0vE5CN0pre3zfhdSkdd+EO/vAMi7qg0qGqgRZ9NH+M+RW+a0ayjbH/y+
xVeIUAi2w+Yf6Tf7iIlb3dqNbN98GqfdO7LAUyRy0haeHXFqexy5SuRRfjibuIM7
kCCJT8kZYLVfGI+68L6xnXkj42CmnpN3CO3VwSgtzhm1VdIRtX99nEPrAeqketRw
`protect END_PROTECTED
