`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VKlIaH84s+iZB8Y5mGMeH4T1bSuoog9FqQwY/8xQHVvC0FG32FeygnHWoFrsl8ko
7szXJJ2LgX4y+cGgmy6h3my+oC0eKAmbDz1xBlNh4z1wCMg5rs3oQuCUufUznQYv
TXOHqth70mh0pylZXXhkxul+lo8vUW2fYd/GGT2b2xIUYir5k/dFYcNuN3ssl1mf
PxE2Nox37P5DZIzHUVws9DG4i7/aByAU0GjSlG9A3cDgo8eJ26cF0SiSgwP0/Cti
+2Q3biF3+lvP63OQuJqtws19Q5lS/qLn2pPX3yXJjzYrx9/8hjzwzFqmA5VPkkAB
U8IpCaTJpbRP82xyBv4EX9uCOxeApvUZrSNlN/2X2VK//aSTR0vhxmM+fs8anM92
H4wG4gKxHoO5/VZwmKV+3CLljoUJcEpiluJlz+Ll51Vgbm/IP0b4lY20EvfYtQcl
1RIrGDA0j5crfQ09uqAVXXDdynW1EVe39pYVe56aRlrmnxef0ELEsYMnhU4eL699
jD03k8Byy7zZSymEMYWWb24AGn7V3E9cJ8rKMW2NBZf3ffr/QmMSggUaBGl+RzIr
9tD4aaKdI5x+KIQ6NCwncqJfLYim3IjZZ2/JVKWHnQXAM6FC18vJvQhEmd1A5CJJ
l7dyh3QNHeyojEexEO17Vw==
`protect END_PROTECTED
