`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qdarZmMgptOq9RlrkSA7D6Pd9GkLur6sdmJ0UCZKFgSVIVKmNysPJ1Bt7wmDDtoE
KoKo0bCpfkkx7ipg72nOvKXsppURx12vKzfOd1odc5rKQ2RZIbKN/x83BbPwF6ZO
RN4e7YbAnMHlemItmMdorVZNlhUn48w0VtOGwdnEwdHnMj8cTGGBvmbwn0zv4KPL
BhreXUwBGKjA43gGwf8OZuu1r0yKhtXFSMX/o6LaAKEZ12wcrh+kFju2TAGgAKaU
YJYYj6yB1SBq4Gl3xRKhaQ==
`protect END_PROTECTED
