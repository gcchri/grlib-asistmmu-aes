`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9fAIS/19Nsd/K6lgncJ28lReCxX0Uq8z+zBCTUr/fXoWJe93qx5DQ8zCS7vaC6CS
/HRGC9KlMYO7Mg33SHQwW4A3xizmDOE9E9Tsxob3M+UT17XnUbqGz1MVh0ij0dvk
wcpSc0XMEJpB4rkIAuU6f+JWqV8IiiQdR2UQO+7zbdMTl/2LkXVRxpVIrRO0ipHn
/dKcnPndTxdlstcW5EZ8WKYq+8iYY+/tFl9EfM3SVVEi9UIf6W6REXPAzPUGlt1v
9hyO7I6wdqniVbVwERkTKc7CKWFG2dX0uZTvSU+jzZWC/WQvQR/2T5X251mMkx+L
BOf/c1HzmE/abMLRKpyzdT3SLOHIHmuJ1EvrVcDSk67BGmyP+V0mwSXJsuzgBPab
xBpNIrxRQjYXRfNsBC7KeO0MBOm/1SMIx4IAjPrHX/ITeIrXWimU7w02qCja3Vxr
JY97Hz9AYYklzQGv1C2GakM1TojdAolPUaECB51XCMAwibwb5cI2FrgKB954nXy3
E0ZttVcV2fWgTs3yHJQcpw==
`protect END_PROTECTED
