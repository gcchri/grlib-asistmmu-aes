`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SCcHEWn8aRg+VeEum6DKWp338rhp+MUMndzdT6xLX/mMfTocuaD2EXiM0t35kQ6O
UA6z0Rk44uV6xeK08HHvhq8+RwOgmPWiAhJBH4Fz83iOe8rc6uxF4Q0oQDwECmiQ
frLo+nnmInuJOY4lzD/AcJ01e7XHJ7Yld/LNAa98dh5Uvm7FGVSe2KEZ6Lylu5np
O11PrhxoJ3IyinMSfsQiEvZyiQq0w49hOBRVaYesLpTTiuIFTHVYj8tvW+c8i0K1
iX3zJ1HXcqae7mnWgUaGNDFvYnkQtaZIFme1hnUiiSeSeuOsOGa7KsGHvupVkw1V
y4nVYVmX3pDsFlGRtdnecQyu5VPFFrdQA4QM4U8KGleMwZLiyrYzYbvwWWChBAek
FL8B0Jq+Wo0n7rYVWgvvTRON86GYAxHNwuV2O0e6sv4lSIiWEzaKFHTHu7xVwoED
5YgiYULIIJ2wrq/YzrLmIXdWySzQA1xjziaZL2A2Wkg57pdA/S86LlwW2kR/aw14
OHcCDteGCHImxQpon5BcSURCjSUFrHBnib1m9ZTrAOgJpm/Vmw9cbW73I90we1SO
EXapplynSL3TyHm+HioKPENJv2Nas5/1iqH5UcNGP+TMMIwvradfU6JTtoHVokUw
tAlVpxWdJtCP58QPPp3uvtXafJ5Nsw/XT6E0cXTSweaEHt9kllQkwvT37aRj8fKd
haGvp1uJuuWxuT5NS0n7F9B6W3OecYv+4lUu3GzMVIjcYJygvI6QUVMY9cdweEGA
mzaXacUoszf8QMh5H8r50LD4zxou5xQj78weL0l6fw8jrHJ0KHFjXcuNdkzdLkRr
HIn03QHo4CkGZXLh9BUAKCs90qGoPqX9cdi0Av2qfuiR1lGg4PQMBh9pjq2mKGFx
5PgA8HUABqm1/irvhqwhOnWtVM6okoRuGvh5nVSEllBeSrcjBftC6WUtmchRfFft
0Ur3iAlg1dxYIv0i4vi4ptRTH4QJbZ4NCFlvmtPZhM/Bd0KhYFaaH9gkDentzZPK
E4x44rtowPD3Ks0rAb1AB/f+BvU/pFew5FJNrxpvtiMviytyf/PNjIdar66UljyZ
7dmsBDLYeZwAbPGvvAJHqE++4oiJVDhQnL3P9AuEXw0opmbbPwVG4kzFzzkDPKvC
3UTKYqsEWtFJgtONtoDd9aZO47JwxHqVDN0uD/fMiMM+rugoXx/FVBGXzx3ksp7U
AC5VdAv4eH1dDL5rpX51VPbqT93ETPF48diTv3wKnTmI/flGJZj5AbmpkS/KweOu
hQkpMihemsdxKQnwrzr+MdfUg6p7J3MJ3rc1Y3l3d2xurbWr0sDQtS+xLTuV5ImQ
SBDFW8iZhebBaNGREt6nJoN5lLZriktFSC4h5EbkoZCh9UvfrBybmZBGCPPFO5tN
r2ZFIYb1yHTXa7g5cGBR6qjXEKXEyYlBLRXZLfsObPvPPDB0grxrkTep2a2aXdzt
cgiT3kbggRSc4xdRXst0VmCJPUUHK/CcuZ4TQBoaupSzPyDIHI/VBRphQdIXEk1+
IOIXLCnN/kQflWg8KiE4GKHuTo9zxo6JdRgzI8spuCGBHhhjaDVHzd4w+pJwOB9d
Rdk/tG6ZdJnUjHVhOlok7FjmYJIa9H7Jq7bXMSYOSELRb2BtVRDeWeAVGX77XUtH
XZpCZKp310xWoUvXDKqaukev1X3+jXHLzVsc7bwUTQLbAjVreyy/55kAmLyw+Erg
bOxaUneFlSB9rCrKmr16UEFRihUERtwXKPIAQcDrcI5mh6pVZzGq5TRugFgDGvYz
MGasHreejz3sgV003IKILEd19ZXf82JaXLjWBV5Gs2VdCFvwkRYmeaDWr3sHFWES
6QXa7m5ye4aZ+nJlEgaQ2Aca+jEbhbVwKw9lN3dSaPCxOUpZGb0ylQwKOA9SGokA
VFg3L0FTclAidV1gRLgVVsqVJjGUwMUrgtq3RqC0BDJZ+a7yqUig9xd7gc1hP5rC
+h1HwvN+YlGl1LGzE8x75jvJd3+8IFv5ZZ5wsd6hOGgRrO+7dxjFvboOwet3WJMo
6FqvtOwOYdm8dWM2GGvjFLmibXK+TR65di9+Qy85YcUwJI+nvV78NLZjeTdds2fJ
Aa+qJWeCwICpMM6lP9Rary/xeqiNeTa/b6N1Dx0EoHSvOCWKr90D7az4RJRQ37R6
CcOclDoH7EK71ew4RwzzqhGSSTfsIQ2LBTr5AEbgGkgN6DtT1XHcndt6w8cMX54u
GwgWL575lVrxjsG0twpIrMK9QDcGaetSkxavRAlOF5KECNXimYo+wYDmgHH0NOJ7
CKXym/rKjWVA37TkUXxzEoY5dYYvtGp7bBAK1Vhp48/Jgpw455k2I0eOTOXHEJsG
dtqvadiFnwOvWIT5mLF+t2wfRe7p/LlvggSYAza4xmTXYqwXGLt0N6A990Qpjyyq
8txkCDILegtKJekX5vx+fnJc7ml1Uep4i+9gtgwNve11RTctRmUiPL56mv5a+cZh
6HtBgEphghLIoN0avnlj3tR39i8nsC/4FQ6ie4dnasTLKcyjnzou4s2wjOCFcsKh
Dylza1do7VcxZ71h8h1VOnW9iBJlPw8HqngvzbnhXkuxk/vtZkHubJSNkvbTPVyt
eoldoww1TU33M7Cxr4L587Vy8nKhmJD2hEmjMIXQyP850GbrJPZn1mv+MBiMxgx/
Kj7Ot80lFWIbPz6m4MUixKSjdqvsaOlSy1TTwdqUOU8Pch6vz+s4o5znwrw7TYRU
ytscYIhrP2A34MQOpnsYVCb46SQFJjDkLkzYLDy2Igfclea7oEJL8M89AiHz5ILW
ePgAfk5Y67BePrP1YMugMtQbPWGigLD5j5FAzxszgDaAAfcn6aRmXiKaLroEuRPd
qfDmVi3aQTMhvTGewqr1oxRfk80ad0xSgNCOOeZWuCck0jxWFIgwiiTPl9mHV0NL
WYg2JNuT5sGktQw7zidNNGEuX+OomCIl8e8t35R7+dpJ0JQFg7o1FAr4oCANHt+r
PDG9AfIIDv3CLKbCN1bstYYp0Dw8IO8FkX2Yx1Z5aRD1EYm9IHkuC/ilHv0DbLOc
yYq5Hpe/go5TduwKAWgcmloHduQ6N70faivxcwgZfQ9RkkSeBzRbcdwYmFa8i4la
52xDaiNIZCDsB+v1prgIbRtLpOWauSWDCgMBGwpekBaIbrYBiM7lP5xoD6lUl0Wo
GFnZwIoXq0AcsVIySBFbFN5tjt531u04aIFq0JlTPGEzKjiNCqL+OmsCrgzDRIIH
Aj2QWb30aPTIeU3CExx5dEVTw2EaKCd+AjTQDCmlHAEgIqKQzOMNMrNOIviHe5HF
mQnMb96eiUkOkb+kJBv/mBNccX0c6IJL0euefVL44sr1/M1qLR8K0d2ybi+31vJq
FmZbLZm5MfJH31FtpGHdWrf4X/5OdHllCMBiLgMBOXfgO2RHxnuwXk/wVYxinDZy
C/VRAfRMElz/B+mMIHSnsZmv6qUV4YZZrmGiskYxcFvl9o+sF7qoFVnCd2bcI423
EW5qAduHxUt7u4qGngwt6ZE4d0nwDucSVXX4B8foC0diZ6Guqf34q+BjIUhDAoJB
JOUM+JGpafQOQUiwZSdBIqIdM6KTbF1IlogjNKCJQHBnmEMFZYJrjm5LHeRwdDvG
yz3jrtMg+aEm6mSFDIUBgifa6niwRuTM4vKzl1LbVy13p5ufPdm8WGtooHMQA6iJ
5ouDiyu3gzGmj7GxnC7zrhxarWnZY5zkkbi2E8wtHZ/h5JshzxuqGgZQMlcsL+Em
zoedPYUs0xO1uzW90heHpVeY7sAk/7NPWGKYoXwgIspXSHvKWjMYpE8eXDWvujC5
bkefkggJeZyuhK6+v2cw5/gRhndhHOEZCTTf5W38nwrS7Lk3KOMOIHk6rukbr35x
/gou8FDxlbA0Dy4Tz/UT9uMI8tNcpQ8eODK8AA4npIFWzqv0QF8uuJfQf6gfFpLB
m4yAeYfmvKT6Z2Vqpa48OXcgHm/cKhxO5bbQeBSfMQvLLV00dO+1Egz3uVfayQ+A
aJkALmAipEBBpQClVJtpV3TmRbfp/SxsIOj/EvLYDMaAeWdC/qb9JwBqFgVRHkal
wffMlREeQErdKAIQ2A0nvjBaeVkJvH9udEpSbvsFEXImhkwkpvoRzKj7HnZNtw+C
JPUbZLACzboOAa3t/jCYF4GQC8kWiEaqqut42oRNL+9BpxZm20mgECbsDJ4R92i0
ebZVJGNzBy1as13z1pabmPREMAiiCUc6rLO6T0LrM4t5HD0uyY+oVsF6Ptcc3h9x
MwQwZaxD7IaBZrfbx57QLzW6yJrvtOx9EziUn6QxIK+OXNDm/hHHwNyooTV1vyXI
22n00epQA+GFlh2qTqSYkmWV9JRaC6xq6gNzwf0UlPw6IxpylmzD6CSILW1hRu6z
PqCZ11pj/t23RaM6849FyxpT8XZvokD5T0IVL4nwlzTO8QD6DPudGBOCBuq+Hx9M
nh9Q8GTHeJXqlxJBdt1EjyvxswCMNudt9rAgnoA5MLmL7uFAyl/F7uRAHejzsF4L
6hTUrACMMe7wRkEC7hKdBueKnzvU4cJzB5w9aIM8VTAQiupiy7KV0QhRoWIXl+o3
352CBv0fUBgZQoQpdcDo3u2ERrUIJmJ+WhgIzejgMAIS2TxdXdMYjM0AK8KcZf6b
gTGdSFrI12FgH1oFD2RCxNwEDZwvGYbA08s5Q+caqMdkxd+OXRUco28SVRfxtWLg
WmO5ICsKU+IjBQqRWHC1983gp5jAvJFiBYc1P1YofBKOktLXtCSl1qg+QrHwQjsI
SA6faSqbGKh1+dNp1g3I119j1VsovSCcfHrqgn3WngmY1Bogh6RJeRx4KaRHM5NX
PkpJMg1dI7K5m71llF9Wv1B20gsYWzTYcrhaKjhPgrbXvzxuy0ireXzPEirIuyzH
F8gyQRtXiHj2VBsl9RrRewvp4SOprEn7Ci2JEyuf+Hhmxx6XdR/QazM14dMLqQG8
uK//Y+7hESNSLDelflXj/JpT66WFLaY6vIU0Ol0FOdWLc4v1cL0hHBLphW0HaKKe
0SfEO5OG/mCreHRNGO6Je9nYjQxNYGYWuVo701xQy8ApOIHocMI3Z1hT9N0St9L4
8NziPcUkaK5eisa6wjTkh8txAnleT3UMNG2UiycRx/QiUpxycFhdMS+G2p++/tQb
o8BqFjQildvHwBcB2D5dFtnKKBleq9NsNdCpfr8WaA0v+aT1s54tviM/E4CC0XbG
AAWunn2IvFf+oHyBY8U9xf0gmaYRo/m7JHOw/cmlql51498WAfjyZau9O3t+kxVA
ET8KDsI3S2V9I1fWAKizZM4adkt6YbsLZKeFG1lJvo208Atr1+mk1qVHd34cP+4t
2CgXvU1vTSzJ1B9OBXrn/+2PcAfd0bkU0VAewjGbo6S6j8ilPWQLVUS3zASEa0JI
V2vQmtLQUUUqraA5YIX7I1sGgCszyU3QopysbZZ2WvAYxfcTi7OfeP4QCq8sRduM
q3Q8grL7iB1DYdi3i6kcepdDwMZpNA2V9ySTohrqGqaoRKME2jWW0m5yVh4iUkwN
8nNnMMERb5oknIUCqLcGng6fiIiuu6vw9e8siMjbeuSQA//7aH3+2R7aC0L0wcFZ
gYQcRWkS4PW6ZAo0CyIwFtebj8N0W3vbg/jUfWW7srKitRZBYgkOzW6pi92pbIPF
L83l+PDzkSxzvvjQOSbzHcsbCSEGUrnauiQfU4WcybTy+wkOIUAj3bS30NEH2ZcT
6SnZ3s51lwQEb9LPaWTIPWifB95EyID3DubD105xdRklcZKjMKdUyXxJP4KwEBCo
g/z3jRKdWTOzPyG9V33bFk5oDq675ROkIV59XYUR68gMMq+TO8N4RALuvNxmgToz
Adcj82Faez3dgY2xwiyqB+FQywUcsSJBkarSfWQlMMa9QeOyVmNfkg29lMYil9ll
c3cYU0oIak8UxzZiOObzqklPYiXe5KQJ9vzUggNFE31UdPscjPrwTHG/MfjCOft0
e6YaNBXGS9r3nA4j1dymuUHw4lCGf+8BtKb435BQ7RY+cssQ61Fx8s8Iaonb8bwf
s3xxiZVoIKS3f31hgzAHMLgyLtIcl3yT+pCE2WaMOCPOngP4Y9VYHyIK7LBLXdTL
w/zKejwQZ58Rc5EpmeBh4zAE5fCTe6KXodNVQdoCmjp62nsyZMxWlLh11ktIeBdu
cqOAj7DWjsQPEGPGXYurzcx3D1pS1fWzU9WuzInYYz10dLwqGeXp3NwVsG1B2klg
s/4F5WCyrbWPFERJeNjv5+SpFQaEnjtfhBZoAVyKkiy4wSV8kBHo0U11WNZjE9zG
3QcII089fmZYzRL2ecPoJVLALfDlQmwHiEJoutLQecci49AIhWTH2XI3b2ISyrd2
d8O1Tv+BRvrwmpZvOjlKXzijaFhgqqgh8JkyhqpsC+S/HfOyOHfd72giaGWsLRQj
ivqfC58xG4Wt+ElYIADJfpA5JJTXdyEua6CroH8AA2BfZ+74n2K0V/fBy+wZQFMI
RILoR/IiDzAXodx8ESWhE5WVb7dhqZRpSIUON2ddyNjYWvdnNO/3T0bOC4HUAjwP
SuoJDZi0yuHOW5X0HIu9PV3/8YtNM9b61MZbx462q5gd4283Kx64OUKVMobpuljf
y2h0pOjM9ptphIkdSwekNAzyPmFXHdudLVYY65ALDqaZwGzxVCQkQtlU6eluCkA/
P5kxth0Xw16r9wDej6ALzQHlkUK/EAIUhIMsYjSn3GzVf27dKlSFQxaLQns1H/6J
G7QfkSMgHeZhGlmf0WCpugG9IJXTmEB5S1V6goRRXwVtdVp+M6WAWVVZNnm3fIJa
SLu7YJ0XgUh1UtSCE+EBa9rIl5k7AD11Q7ZFQ0H3w7iuTNZZMzxIwOo0yZMVAYgq
LFYdK6fwAbK2bYp5eC4ZLsvIZXb+IRp1NGLaBlOzCzoo2itIgv+my4lMl/adOj2o
+kNGmNJzvkdTwRH7HW2cfe83prKnu6lkcjG6Kr3AQlxy+xQvWmjsm89I2FyM1c/L
jnRnnKJLZ19zR0sMB+80YZpP/+kXvfBkOgkkOT9PvQWXTft5k+9CZhW+3sGsx64q
6dTZyYejFjBLkissnw+XTzhLrY4sYbehYzy4hkYk2GRYsdSn9o+NnoRMFTbEYozP
UtvWoE7oUhlQILlXKTy+jbydq9/Buzg5V1jAbZx1j+UhJyyks3ZaCFAQYcCa/hGi
7ECDME8E6fIa3KCcdnGfOqS4n1U3fAUMa6ccnctUZcylQy123h4m+v8UxnNZ4M/S
BLCmfVHbZQMZP/DqoFfYwBqOZCLPiahJF9pBY0Wd8meftnqpCrP/8c/dE6Cmby1Q
rS1tZ0TJiWEbCJMPMF/8cDSdND4YluMIwZODzcZt+Mzx6RQclH1T8ikAu37PP1zy
F/8x9yRKmy2fk4HIkPH9puBQMOkjfinenBPSiD03EhlITIvbgGCDfHav98MYw/Sf
xxyUkVbxUVdC98j20V0iUptQMGNbmvByhvHLfBdH9LohzZWlSrPOZHO0s1EhbwWt
6zcY1eua3U7eySREbcoJytrQ7XGWo9NaVLlkvtjQniAtzjjoooHX7oFoCVNgG6QS
44mU8QDLUYRhNsPu3OXh+0v1nSaO7O96kuBjulRmK1dg6EP6elMS23eUIoXi01/R
58nZDpd79Gm/BETtYQiwIyX5c4ydgbjGjC/H/EE8i0tCwrN7OhKAUCGLwV29Vy3n
049bUkC3kjPXhz3SKF2iV5xCbemuHL3BMVBbJrnc3XZ35TLhvlklymvScOdMekF4
51m8r4qcV6rlPrtcvvt4RbQsYnvGGbZUvVC4xEH17nAIP/IvagJ4gM+fQ8N30g5y
UqJAFuoak2GXDidyIvF3LITNY3ptcDpt9GxNVQ52m02hKZBoTk+mSlPPO6y/3Fdb
PpLsXp/fztetoQBTvn4laTu860c35hkVYEGczmd07PboS/OB0FbBxrHNCNswFdEQ
Wj/dpMqHCgGrAhtGZDWjWf0Ml7/w5bCXgP9US4Teixtnfb9Ybb66wt/DLgtuYupS
YX0ANhMTfgYkhxerG2w7thrJ8dG+5K/abw1Pk7Lq+z6FYEh8gGofQahK1dHRMdig
kdZoWOjXdFdcL2gCUPEIUISzp5WY1yskGiByuFVENCSnaH9TAmzylVWQA+Hp/e/F
NyWcoGXI0OxaAXXLjDmf69EqlGY5sRWj3U8fAqruX0cD9ygiAZt3n81h6P2dVmKN
VlkAUOfw5QZQcKZ9X42mnTqtQOggBGHOf1jCwfMvLr/GylUvDIKcCzqH9OIX+Vb6
NUahbWI62eHq8sQrrOKM7SgDnRtEzsK7VmP+ysfxxWCGHeWy5wD2omT46kxPEAKI
4L0J2Hy0fkh4UR12uSlQGNFqBD5z86Z0SiKqw8DDOmWs2a6QI7T4HCMzEvSqb0uw
xxD5Am8PidykLoc1NhieJdVxBQKROJHhXy+76H/taLWWwH1twUl7uORAqnbkukku
uKRUU/bbAr0fSMiJ470Miq+/ORLjt0uZ/rOGvl3Qa80c1lq5n3tJNoNNYkjjYbRZ
Dmtk7Sk7Bu3CrGA0iCaGHgMEwW7XCLem27y/3uAf4yTDMkG6w1sE03cmcskZjxhV
784qIrJUhHqap22XwxlqppMLTkklXsNA6w+U2AAUpwaZyi+dWAoONP/adrEowCMM
IzAiVRhJ6E695l4hPPL9RKW72dU39BOi+boX5OcVC5ixrWwP+3/vcUWrY4JUbifi
+sLEV3XQfnEm6olM7xhp0jKiZ7Qaw3I3XssibwqjHlNkGNAEBXB4jTkSnONGVLHR
G7fq9Fiyiuj292Qo3dOFHjcs6xsSLU9s3L2kTcqfrEqGxRRcPzfQi9uUbNB4zDuF
QVsZ4RnE3Y5G9wInG3PHS+qtDbFmZaAMUXcdMygaDhyL0zFPjeE+hjXB1itdkGs6
kg+jbl/cg/DuZ4D+J7I0xwYWMiz+B+1cIm1vmrfiGRKlY2PuCDW18InBHKjc1C6C
IrGhwyvqlAzrA4Jf3bTHf282NkMRJwn4rn+5+smw9gxsfgeSJWS9/tdw4Ig0r/za
aJ7SzggWPUCU+QdvBumvhAKmefKJyAeT4brrTwzszOwumjUnwjiLHLHsbcMBKBzV
KOUN6j42crXSUnzcmYiFsiZGP10BxFRBzVSKejRhCuwt7L0cRdUzXZWRu2Kvhj2X
TfrXbgRnynNzstrc4zw2y6b0LaD+8Pl7VCYkrhU/w+kH1d9srGcYgmS8RSsbBRRE
pthdqgu9Fq7BOlh/hwxea3e860v0OO8YqY3ZUdtxAsOwJ2xml9U4oqFwqtHxFT+m
ZlOm0sDgxcsOFmq2T5GCMeKXSb0DJB8jJGDG8H8NXFvivLIsjzkFQcB5TjpRllne
JKj6t5Ti54L0oFF7X9GngQER5Hq6MiwF7iA+Iz0e3LT+cnxpwpIHeWc+qYKeeAtz
KMvuJFunGDwavxY/2ThV53p3h+0nvs4Mefsy3EqiuxNg36qH1bh0DQZJiemMQBNm
EFg/JUDFEHI/zEsCvUwN67EfHCv3wbOR74ZgYolMalc3lHVW7jdhA3ZsxoxqMmRR
n+ICWQAJbcmjqqSjPQJYjPcJ17/OFlBoj1/xEfghrAh9EhKTt96Xbt7eIyE72aUW
CqT3tJ6uba7HGdzE/rOsvF9qn/BLi88KCqQA3pClAKKPvafognbr7qh7dYfYz6sU
pgeti4WVDa6UwYem+P5nd7Y2+BHv8VgST0fNF0LX0tEbuMSyvQZTwhG3E11PPUS1
QoHKQD/SX0uvHKgadc1kvZD+RCqg1UVSA/F+Kn/2m4hfgiRAJGH7pfXsBXLJ390o
Nae1sr6YoANwDDUsghLhlM/b96q0oWVpnqyXrYrloorFw/1IfA6HwzlzHlcZOorE
TIHXIrjJo3vysb1gRK/ZdSv6DMhHUqWtGMlrbYINs40aqZy57NVSKyqPeulxpnRF
iUNEizI/ahr8xHW9+iSrLfiMejmWYlmibHujrVnZUNk+JSUC9Ms8E38mEdrBxQW3
k5rfTz4Fdb/0jqCQZy46urhHriXMvBol1r+eLC0gbGOCxLDQbR1tMZtkKttyriGJ
6O4eWrWQTf71l24Bw/gL4y1xbp+6i6TE2hiZwUfXdgjvgzaIhqQwpBG2wr6UtHDS
k9HkRf84VMOZQJbBODu/vagglK4JFLz4tpDOr9ACHufHXUP2nxOCXzNt3Me0COMh
NIoB2wgtNzGKVt/I4JfKzH6ZCDjUXyMhDfzEiN7x+3IubWNQQtp7T2yTZnGrCnh3
BOiCGgQxx85GJHeLZfLvl/U8VMe7YX45xTI8owgee5E/+CT5Rgm2kyGciyJFj5Yi
2Dcn5QEQXI+l18EidnadntAcCmbQg81bGqazKmeXVPD6dXyioI7XknJqCa8WyU+y
0jGkbq9SpuhJnpC+D0xO1my1dL/7iry5gyci+61UBYAUpB1vDcHTg5yXZZYfP+Uc
leCz3dvQTON1UnmURWRsps+HUaLYQ8dp4A4MS/vng1vCOi6xppZSoVZ4o9SsizTS
AE9YgyK4QWNWIUBLUX4ULMVJfrZf/ykV0OFYIuzXp7AOl5JCKu6ra033enPC2DRd
f+FtxevcHOZfegdxzEpLiLnwzjdQLDIKOYZioZ/puE8TpAi8TuPmmU0QRmRRFAD5
IHwnRsM5cYCpaPB0znddnThpaaC3qtp4Wi63bI2p5mIT2FYyv45P+SF6zJU4kF32
AT/os5G0ZmOX9MquCOyNcM4zqg8cZNQYJVvrB2GPZMukuQCD1CrAbZm27v4T1vHu
8V18/em1PGlDoE5s1wFt/ow0O3L3wEkpgX89/kVszOApcQ3uSzntorjjFHQX3gXW
dOlWR+dSqplmzUxz3SbZ7jrj71KnyHshhZ0lK8wjl32xzTiXzRdLx+arNeSSjhT5
5S7cNlB1x49oiSDVKYYo0JIB7h0KmLq1ZN/TW4gRTLU1b7SpK6gcXpc/M1DZgy1m
TYrDXtqqaD6laT/vejRSgdmdffQdtjKuIIDIIqCflwM/WMT+Z+NCLssIl/7d8qkP
W1cMl5Fa3E7vOjcsTKittNtChKNU+1OxP85EIoVsY/jlWy5ChTsvb2ieRLZgFmay
aOm/y0pvRtaQ9wYcjAw7Q96YdzuO9TWBgzAA5fmnnj3GtV303VS+iOS5Sj+HlFvX
Oc+3nM1v3Q3BVjHguEi4hdC2TqkQSZ/o5v+6o8gbqlmuOFzEEFfYsI9dx9L/7IRJ
BTKKJ0S4tgmKBW28yyzlIGF9V2sD4kR7Pr3s597kWRPHiPoyZu7jCEMHBQWPp7wd
ZSA21nTGhb1pRdx9CyyWnSJCfr4uRmCZ6oMI3gXNuHdSDfT8dQdJn3GEMt3R/z9K
92OZu1m3btRz7aYrVL+l64ZFHCAPVlEwLuVrvfyzWsWbGYtCRfbTqJVfTNqaGH2i
xRHOLvarxR63qJXxMkate9/uw2TWvlS0+XcQQqB3L+j3HoOE1VNk8CSXqYbCl99e
bo01sSYcwvAyf2VJR4GinVQ7z4jkkccnnkYYSZav23QdYh7yeAXkBTWeAeLaWeAb
Nwrdmgd1ZWse2tRClyV97Wu1/xETIEe+AHT4UBy9zNOfDPs+ZXCBHFQd9QE20s0I
CtgLATYqjDbJQB075xhFAO0ZiWytd4m1KcKfQWekJWyL8BcETIp1KpX4U8WiwG2c
uc9ycm3+uees3wKjA2u9MygfDz260wTBAVZW5UXUBCwsIH16ZKBvPhqRTnaBNIsh
QfX00UoRpNGNW4jCDiLSlwuyRT/BLbY4A7tYfleunxNmJdBezc6/IDV2ktcqgKug
0n7Dxr8oG7hsestsKIDu+0xHd/dWS2WRvBIBoOQU+sTZm0jWOmLw1Er28xS0eEJV
WxWMRSGols8TUk3VeM5fM9SNijf3jItx7jG7WUKb3sUzBUZt2fyfU2hzsEKJr1V6
boMT5gVdsHXMZz3FTxic48/WlmScKWipI4OQyLg/MrT6SkRR3dLTIulOsWvKNjgc
pIz9joJXgiFHpEphKYKpXnsIjAFGp0nGyEldgpZAarOMpDxn6JqhUPAHf1eteUI+
CtWk2mjd5PpW+POYf10NGOvJX1lnblwujK5i5z5WsRho/be3ojvfCrF3TDCK4KcE
mE1ohruOs+xWaMUakaxugO2rlPqUR+Jm6MwXcxKtf020tTDKzGvA2CnDURz6kSHh
fCpo3FlZ/DDQPbEPZCkdZqcKfXIOlVAhyZI8XFa4dMyLX0e2D7v/LWQILyB25w6p
xlNLbJvBPPl9o9QKuUpehfk2Sq84Fcz+3kkaDZ+yCK8tQsU/hmASOJJNK2w+OVZ7
1XaG95Zy/RZweE2zpMbOKCRjOaNqMeP3DQRSBXOkap/tJCeRBqRBRreBJjO3L3+u
z1ojAkxmGxTPsIICmxUrmgo0/nEuMaiWV6kEvyh+jc52KPQQulhwyKCoKS27uHi1
cONwsYF8DChk0/pTBJBKlgjr37NbrT9BP0si84rJNbR5KgAOIaoswvw2/m+FWO64
+r+Rtd6HGns8ryp7LOx2bDOVaLjIdTi8CgMeWeYkdM7EeAg7AtLPfdnbdM4LOyWm
3GVOqu5YqG3HCaMCMdge6Rlx60SUBCGGTwlKAExbwtFHQLGFKY+yAHSgHmlhGAmO
nRsIZSg+zFHdNuNT0nQfANI5upX5vaQ0N3NXEdtzc7paRtrR28muSttbyAL+fDeZ
JULqHCAp2SX5ImFXozI0Ym6bfgDaN3IM7RP8nAA1v+Htv7r8GNVzdd68FVZZKbLD
B1tpBjKjpYiendj/MofSlBhZIFqVsItyryKxhlTmLUA9GshQ0UmQg0CcMMvyqTUV
w4/VnzWmelNrNuLnEcrm3Mj9PS3/UvOwf1tnQ8BD/AeG23bd7Kv4l+DyPDB3+g1b
39ew3krnvMesblRyNwhWUwSLRMhNiO7pIlaURrqW7n0eEA7Vp63IE2K87RxLZG6/
aq4ZrM+R9i8w3lNuXE5EsZBTsEEjjVlyuIv10TpZX04GUZn/ktTGk7S0ZsGXtpDC
ehZUGVdovRlwVDaGhGrcp579QWZ+EWScFzZ5RKA+p7SJkOyhXqTudxoO/bwd1sAQ
BqgeXW3khxyJvJ2Eh+KLc8qFWSOI2ZjmXrLgFnYrZHvkod0pU3OapL6VDwv7szKO
83LVBgc82CPYT90OaOvz80VMuISRB8oXYu7c+Mw5tkGQPBJ2xjxhcxYR4n45lA+n
XYfSmc5p3kFUDruRAitmlMVHPV30m946GMgbMyzzxK/Cud3Vx226v8W+OxnBegRw
oNZxoCmOX4F9nwQpYPDzOK08CfsDErnBT045FpIIF8B5/rMacn7k1bupl3LnFSy4
8savLfope3k5RElImgdl1iNgg97ORfhHLwGbuEOl7GP7284kFZgsJU8nv1SSEZwW
hWHFpXDiiwz9YAQMeqQ2p1bazrpjj3Ehdobw+0xJpMFAmhmTXlHHq6J4H34Z3Xnj
nIQQUA/hqmxqhcMBqL/P+9RdJrk/13ez3aQgliPmHYwCUvJak1tG83Cogc3WbhMh
HjqKWQ2GkvRz0mgghGxMqywzJhm5Kp0/1B+g+hEoJnpN5z+TZDnX/i/bO1XG7J0H
r6NOwk480bhRIffN0AZnq7PQbFIyE9gZsMI5vQB0CKh88gaimF5m7/5oPGIF92hd
3y3aaHKUsaJN/gaU3i2/dqPRSndaDS9BuBH2LVwc2wPSwCKLDwZ1BK04dM19Ldw0
oRFs1zmcMwgbb/om3DdkRAzPbBlaXZdUaJrQfm+sSR3xWZQ8TSgY6QnImc/pcJ0E
2oaCZ3JB3CbaQjZGmYNf04r0brp6JhpHdoW0TVDZrJiilhij41k0ZGxWh65k7vfE
phRlk75DWTvSxW+1B5RMY2+zLEHGnukwV9fDnnYEAVCwAi5Vav1oHqpktnJ0h75A
Xk95yiCc98u8fQi8y8WdhvSY8kKZI68SvXp+7hj2D++BmDZXswgHxnHl/vBrn7PZ
HkBcerUQ6KZWYlz3zUL0kbYMy6gOEhlaQeG5uFrjkQ9i4SipiFAH2h2cVEwl8hiZ
Ga0ZUZf8/LtG8nq39oBDFZs4G7yLpOrlgU8NKBp5q8mGfRafkgr5u1xa/E9ZUmJQ
oySXQWihED7RqoCgJrqjFU/SV3+ifxLf6UPWzBR6XrIdSLEy4Un91PaWPC0216wT
WWUkx1WW8SI07zrpEnhlFCGL3bIbf7KVlrhb29r2EL4fllnu27JckzFSyPFnn+Tf
wj66skPM3aNGm19fGDaIHjdhS/skk+FJz+QMvgZrCtFBDSuxuh8wb03Xr7P4S749
zYWwlNL3pj6xq/mjKYDVujHCSIngasgl/EK5OD2p9MyEkifyw1eSPs+AdcuU+xei
6jd4trxHH9rw4NsjVtZftN977mIZv/yme4QATLDguxl5eAVnrDzcN8zrLu3nuvFr
9VStzX4TgGrcUktV194duKPbOZOakhqxGTsZdaMcqietRK/8ZtBIuoP21P8dqQcg
Bq0a9wHZGOyIcNKU+jCqcOOJGlNGR9IK+4+MPpfK+fMR5XcRSIo7q/TQl5s654un
QLCnizfajgbv239pGdOufpj10QVBf69k6j1DAOIMRjn4uczKUuI7K3T4xAk3xMh0
1Dgq8szHXBa8c6d4pYB5rpGQolBLoSpHnrQ85DTNrLBjQcLjPG02W3knGpZjKzLt
PD9mdJlBWHjleSa6D0iVWqVISh/3AIm5TMVFARapnTq0yclRxMZwdsLNt804npHd
2CxkxSl3hK4t0VWc+BzirZ7g2JVnMOt5704MmcoZmJSXUjo6Pa9FW7u0Qav3kmmg
jQZ5sOGXo0pzKR4GJADUi3JRRbL/IOn8GFE0WZI38JYQ1AndqeV+xfNarNNgEr+c
U4BB7k2v3oZqcUPtO1c4Y03+q6ecjtJNXxyqcaql5+59ci+Sn6vZWgQlzuFvLlu4
qwgSIEvWvYjFIBEXAzT2r7Asz3NGjavpyWt7rUGPA0oieDeDUsVylLSKL6bvmYLb
2J5uBATM55xEZ+ZhhRv8r10jzTe1t5CIWW8SvPlZZY+lhxrWylX040XIbhJbfuWq
pM5TgeyxVOEJN2XHwCpqyeCvHpQYFEGvBdeNkhcBjoAz75jmmwhzJZascASDwVX/
hoHOM+DDB4/LMolyGJsyoTkYfMuVj8neuOUN2SPlFfZJayKVttM+udR641BKLPKN
gpSCfrREAiGkSRcgm7/s4+rCiQihSQ+Q1EqQx45yWkZQY/FvT/sF87iQLFUz1vzW
nyU5hGNBy1nlKDmKUnR67MX2ZyWkvU2z0XsBp81QtZZsm8KykJ15oqlWog/+pCWO
rc0kNwhhbIwtsuEDHu3XD/En/rAk45J3e6zVu9BvG0EuKiRVVvz33r/k4ChuQIme
nLGHJzEJYBRQ9DIMxv2dqNoIFsC7F9vOyjzcqX96XL2G9GkbPRtU9YOCyuFj5oUK
0YFYN2t9mFchu5tbLyXTGE9xP8Pi3N66G2elhHGI0zA0J0yi3hZ9f1eBppWXAUHQ
0f5AcBLUlIulxR+G1+Ao9hLt6f/e9cIwAKxGZpyZQ98I5ZNa4KADOOF82HWvcoJH
ag+IyratZCX13M54en6eS5r0ZS6XGCON1VirsWMXJhe4eKPYzFFb8C3WrgB0FCEq
hc8+9sCJ/N5p+eklePm47ye/ArB2eBBZ7XGhcCKxHj6xhRFuy7FaWcXdCzHWCrBK
30+oragvGdpM+/8XpbjKLzZu/YACDeJJaX4XYIldnJ+kxoFfPEbaSnobZmjESozB
G9AWL4B4ed2c62IslyViBCGPeASQiN6rSnFmX5YLEG3yLV5aKIMDsmIgEHMq+WKn
nXW7thXj5AWb4TuGdvVaG+Drvt4llgNTV7puEKpDNhJPE7dnH7vEVA/o19ZFdp82
q1lmfvobXP0dxuAZiFmj4O2vJGlXjtdFHS4e4E+N38jAadRSa/chrk6VJZ67G3+R
Neud0nSi6bum24D56xHdUHMZskEGoQHHtn4hYAPNF0YveCiCZ/anepI+zHRq2gmW
fXwBhaUUy5Erfyy4OeVbg9POPtS2rGxFKwrZ5CujogbN7We2TBchYoxE2S3WZZ1Q
HokHk8TfvtKFqTcGrv/FtBZMTZsDbLRlvi5tkDDgqI8aPF+BA6slYxmJXIiQ2VYY
fufw7QYYTClDdS1TFQR0Goc7saBfz0wfd4fNhWnAXyKVKlxSIf7k8B/y/r171RMr
JLDEbInHztm1fTvgCPYBFkyEMJUrvR6tkHHwGfxsQWeuQoGm+HYzdb5Xnbtu9H/y
F4ziRNN9oAz0PU0j46rHced7xMtSXb/kbKtDUZxw+FES3g2dEMkMSJh3IE1u9fWh
f4DdLjYgejtMFVTO15rWnCPEe9szFlMlCPZdA4Ww7vo1gHPqVMlNi5+JX4vHh8oS
pErJEDcEAzlPnp10j5NFUjLH0vAkH4wkhPR5sKq6NpMAjqMZ+8ou0iWR8N2H3SyU
rSOIV3yF9sHyUsb5Wde5kynsQ/AI7Ey2hYEtfyc35j5Y/TbZzID1AcrMDT0hpaq/
BZctrQBymDmGCkU0Cnm1SEO2AeZq5sBrk0ePjF0P8HJv+aOGfsmP8l4Dfu1AD9G2
5n7PwGajk5LxEBXp64iYCidDzrf5PefwH4EbC2jjdSTuIKLfyYXhm/BoUP6CwQpG
XScyCIF7zRfrKUEBZ9QcGos8GC0X0JRZ5wG89YvIJixUMXJH3aQi0+iiacT0NYWE
0GIPl+XR4AAuGLIvWi8troAIvGdXT83lbS4IVx3wzuAhqYvw3VZO3uVL2eBzxP6X
8cDrW6uZmwThYHepXzEEegVh8ex8+0asABaS0IoukVwK2vD075zmBg4cIF/HXKSV
4dQBWYrE2zd9b6EfwBM8GbAdDyYkzfA6nh9Wh4fBbSw0imYMNY49+L92wvD6KhLp
PGjd60iIZ3Rb+8ER15caihM4AC77iygbUs37EwZyVbt7/LgYub/93xGkg6WBpD2E
uue60gFSBvqXQvWLk3S2jj+G77IGVc7uTxEEKvXxGmSTjGQ0VOBWouq2hDs6Vjdo
XK7PtRbMvzKdBnjGoG1WCOlJixxV9Eyohrz4D+XrTrQnqUB7sH48Z8nDeIgWBRk8
XOc2c1/vAYn/7/zpS5Avleea0+FctjsSVZWJBo3YAiF0rG28jxjoe/3wVaCRt/Nl
x9xI3dF4sHzO4oGZ/vV+37HeXyytTE4BCB76hhARIuW/FTYwMvqodGZ8029LKbiI
u3hKdcdnHm9E25O/ht2szEZbaT8L5+xCWdnUSbOl3wcISWQVcYsFpmnK19VdRS5K
TY7JZiP7sBEw4kwto/1Y7wzhddTcqTqfxc79asqwN8RNyCB5+6NEbAMbM2PAlW74
5PrY0L+8dQHkdp5REAPnaoskNwp+iyGLrSuA4dHBU4h2tIP4zdu+oD3Dq0kT4HnA
JxoY33hGjNr2k8wLssIvz02tN2SueKKjxlVO3hFmODMFZmLhE6UHGaDj25qP/VkN
yQOik49d5VWNZQz9eo6H+bKqZ98+ZAhyotw0R6EDlswIT7/f/YslXdBnS1cy+QoR
Z1if2COTY/Nqgphrsa993LZKciTzrEX8YU84H1JfioJI3nM/1gNJeC4zy7Ab/Z4+
XuHcU8ysC3xIi5MmWQKe8hAhboZhpXkyRBXcSQVODsZ/GylUN10X48eKwrr4+o6B
HPO3rD2pBYWD6uvzWChTpKEKj1r2v58KqVZV/Ap8kzkys0ZW1flPh8zSfarK0iyS
WWkDDBNuAB/4sQSg2KUNVfGKLv77QzP5VsBwCIpacIVtW1znY1Bd49EKsaYIRfrZ
wAc3bWEfHYN0ioOSARYfp9zZeoq89Gp7BeQ7gdjoL8i0KGGDJyAP203GyT8Bj45a
k7nJll8HD9Fg4A6GocOCiR81fRwjtCyCXqJX9X8/W/2JQT7Ik1S4rVYF81mH82lb
HGJ/T5+GwbvGrwqbGYQvBPSLtMncyeCQgl5xnuTXQbj8XHOaI9/81tGDUHVMT9mm
YALt1Hku48aC1RQHICgyRDLG/3ZTPgCUQVsNB6dFOPuHkNfq/hXWqD/aJEqRrRcA
YcsfFwMb6z7pYWly/Pfrsqi2w9HvLSXQHpDVREBt3bRDcwwxi1zXc5lTPyytX4vR
W8BjFkRMBw6F5OA0oNFGbIvztw/32BvrYqgypbJxT5pYhSOW5xDBS8iLlrF454oq
83N8DcV6hcenp73MmYQVoEeYe1E0AwTExWeMCcrDCeuXk08p8fV5BQ4nJ/tX3cjJ
K8M7XgJNMMWGtn8KDuT5Uq+ZNvq3ERQqnL4BnfL5f8MtxjskZvJwLhuvXMB+njeX
kOR/flLXNtORGl4I7KuUGJnvn88YFoU2uURZxUpPMqfuwn2uhBeRQHt3k2zOOayQ
5d4zW6m7sFGoCd6wWcHjwllD5hPayUvXy8kf4NXjpJeg6Os3t0bVX17PpKzQobLq
wGT3+5hSnz4qr0TmL2/50eSwNAzwFlSZ85iTrkdLlTUyzrH/t3CQw3M+Xjf3VPmm
sDdQhFoAQnaF2DqbM2xul0q+QTFOT9d2VwqWqTWpRoPX8HsrkqZjXXzxuarMzKsZ
uJFFiFC3M3mYmAPLRanP5BXNvzotfP9mXev8a6oLEekkCxkvRZaTyMgmupFdfcK5
ep3Hliu3qoHPffPrsAjMTC5jKBExvGnrgSRsTOc/YrF4SQ9lCe9B7K3+g4zEGq8t
b5cQSKswyMAXvgNnbSPPGpBAah+ccdjrwDlcOhmmh2vArLu+7KhtP5YttGjBchQ2
H3wRjMe2A5udcxkoWf5G3hxOsbsWrhDoPVp4BbLZvSLG7T9C2l9rFATB4oJn+TmX
QqvD2J3sS1ACUNJALT6+05ax0l355AiRjl9fMSjOj5/UjoUQMCu5tt8IM7HQb/LT
7sVIMgdBMgc499rmBad2WM+Nn3YgRn2z4cmeYn9Kqj218UgobulZS91A1/BjBfic
Dzz3XFfCIOQq2iAJlA0e6R1uRqMHzdWADP59rSdo+SMiceNqVg5D0/MZLYU5cpOo
311Lj7+Y+rL9tGO7wRaCMEoLDFett48wSEGfoKrveDiuezvmqz2WWKYwEy+oDMjx
kgWAtR006i0sI8pUltYSH5O6v2MqJnzda3YS6FLTb1lo8tmtQPsVCyB3IHNt5fr3
Zy+NI7Tt5Ni/MgYdfgnKI5FaMiQy/T2asNFoN3squOLrEoepeUs47ueJS6HJa7oT
gZ3Zf1J06Ojrgr5w4Gm9rPRQz+RJlbD2o9ZF1tFAweJp5wZ+IH0ETFhrJ03JzOg5
5wL8p8wAQIclDF+JgoiBsV6T+lIN/6o9gaMko4qFo9LgGQaPsj/9HX/WHyuD+ZKi
Tm1sFMFEtO4ErrrdHgOn0mY41ltSccrbAMAnfjq48eazDRTg36J18D7ChtZHi2uE
4iLCV2RoWlmqFVMS/WJLjq+dkNHgSdzz6ljTtHuul1jsx6/1sJLvQX46fgZTg66U
l/aW6D1Pu4iYRYcWewqyERM4H5k1fWI6FC/2TViEFDM61fcWPi/J/FyoqnzP8IDR
zvpOuiyATrCNpTF/9dxfR+6ScXl1SD4oRBCLYogHT3QFX9asdlAL0ZMg9U0ysBdL
TynmwQ518Eoi6SOVZ11EBKh5uwX+ldziIKhHTN4ICh0bjSvw2fE+wAg2hs74SHJA
iXuVsX3JgibU6OfL5J14PWMATY9Bv/aFcG3bdCuMw+A6wD+lZbDxakIVGYQj5sE2
MiOW/S974oAu0k9v95Hdib6svvhiEVETnl6rszw/ADyyJRaotli7/oGtGF827xxl
z74KwCarljd5Ts7t6SB04/lJcJOUp6k0SXF4ulrtQMXSRsH7MIHR7Rb6eXWV0DWW
u+m/QFjankHUs8nBrgLuwhBj+INArfjDUAI9tccgdDzd65J1u4xV5qDlaNCFOzPK
s3lutSSeoja9q7ruA8NAjqHg3m9cy06txuQrryNGHkmsD2vSAgjFJ/xE4O0BiisF
0HKgji/scKgNFxaHSCjSYl2qq6GPg9vvTCanxw/zZTL6SbHsJxHfTXq3NaC3L2oL
LODkz8vKxJq9AKzq0/+GQEZ/F/YAI7gOdT56tDHwVPk/V2ecAShL1SgT+z+x1ec0
exX6AtqzvMaE8kRbe6aiC43o6+4tcLB63sOXgtx4nm0BTsmCFtqJa4j2el+/4FQO
1TKYubD9CQ8KVRlzAVX9tZG9vplXpKhHTJ+D6UpQH9J7/gerFAN6yw0TTe0IRU5w
izq2gaWHgoXPxh+Pda1cZtPJijWg+oOtwiuUBzYIZFaJ4Tda78/XaQgPy6azsWp4
myNzn+r9kLiphm8Ix/bl5CRYMwxA1sZYpjz6u70VpuaX1GbhyUnIQyayH/0biloc
i/+yC/tqqjS1VNuCVVZIw5qmRNtArf42nuKUXIit0VZTcU+YadRj0QU7Mudz2qjo
GN0iO2+6QsAMvDFvL5SK0sc3HiAdjrW716nt65d6tENWM4k3AxvDTM7OavlWPvlP
eK/uGSqWGife0jICmNdC4vDwei58UdttJysTB5bMACa7hmGJCjc7OONBZ/6D/Cpy
lMbqQMf/UwhMBsl4i6+c1zBnp1yZWEvQNZXtH2pTkfvcTW8vBq/7UUh7ajOzOryy
0NeJRoL9LCpkMpLqrvobJVsxPltwPb7LKubEwJpxibt9VD95vPffEMcQh/skaiWJ
BATqGVdoBr+78wd4eCdEvghwagg+RZst/MMIlpKKgoRub7l/wzMUnfW7qstneAgX
N/BHeIg98S8ezIRA+bwOWR3VRW6HeY38pT2iwbMOhJLv1Z76BIhQcaHaatzsbKmc
AdzpdvzGyiGsb4Vap7jNR4l6UMZrumzXsXxzDtJ91toTQsKXut2dEO+HUi7BfqjM
dxLaH1MJterXEMr9Qeu05EbAZDj4ibkGnOaDiaisMsWoC2r4j3Vb6kDOI/KLohNS
ZfvLuBLEWiIM67VyvXaMIOm73yEeqEAdOOLnVkgS7K44Tzee7qSQh9vgTq5tv96L
dJA/16nzgz9mF8znzLvB9UU+FaGswPVAR1pOJO6lrFXwzN5xdEhZ4Ix17d+r+tLT
LWhCOOPRCyJIXw1nDT3fUVXqx1C9VPNoaHJEXfMPszA5Wz3OVnR/PiTYner7lQ6Z
b8+IseLA5ecG1Ak4jb5P9UWW74QNlKqk8xngsxnkLNovzOhzagFT3U9M1MYW2RUT
u1elOQeqllVLf4wSXus3KiAyG4ag1/5kEj5VwLhRwMk80waOQgiQAr52YgBHZh6m
gARt2vx8cmCVAVuH4VJp531G99QhB9zFQ/eTld7gNLR+uuiKK9r75Sbu9PKibU2i
OQVGqgjzNj81rg7/ISQKoI2KJ3GeL+4RJxQQMR4EA57qzik+Ba3uDLKV47bWyEDL
8X/O4t3BW82JEDJ8TMoFWoocPJ0bbPyLjnOJeLSsKnAM5B286HSDvNgPxhmx7UIJ
R2EHVEdLTHxQe55K/RQ0d9JZTauvmaGbdUvEyINTntva9kybAr9hhwjIIXUDvASc
WCFRoFvF09rAr3Fe7WSpuf9s3DLTU9oRzUPN1DauaTLgXrrQKSl9yYXA8+IewVpv
HZKBLc+hS2tpa3GGkJX7rlsnAt2oWMqV8fdYHYK4rLRSVIsi4SUpODOT7suZiGbf
1EkACi0ugWWuy5/mpCqxI3YGJhemkBZUyozaQ6mtPiyo+liMXdJZgCVBEM8k7XaV
pQsijFM6fwbq0L6AsJW7dz16/5/ToNslneeNlkKoT+DcYeRMGMBPa4FXXLfXd7lW
RbE/3n2YceTlDEZzse0RaR7DXw2ODgBKXUqUMIkqQNqCXR9ztFuXUvJQlq3Kl8Iv
mq6briWPzZPYgBp5WU/OKeq31IITFCUphyUSvt93e3Vu1QGFemSA5cYR9bTczbOP
9l/c3JDKQL9IRua1Jq5PwHZY2wkj3d6mRJ+YoYDgt+ipw+ky+YVB6AN9heWhD6b6
+Ou4tGAxcaRhElVry8zkNVMjN7ijsrh8B9xgoM8oqFosMdx+Rx/yBgXhRhuRM3yq
ESzMbZyaD6ThaXlUzaOYN9SNry0SnlnhO2hob4guORbi2md+s/fSmbVRoEwIaxBN
TVuRiKE1lKMhej6us3JUVh6b4aqFECBFgguUMX8gThOnh1INzKdPVY9Nw6cL21H9
WTiVbk/2BVqhxGSc0VivNshElw/ym2jbWNvXNscLF7BcXJ1rJvJEvtpKGpeuvmmA
9VxIN/eqksbij8UQD/EAeFK0r3W0fIBL+xH2CEllZETgvQ1WqIKTN1ZNEBefjRag
qcRhb5KH72q2HinycN2kWDPdGWplxXAqREUyQc2PFkmiuVRFRx9ezolgLOuKt58M
DJNCVp04ph8IavXYtiv6q0LjpTG9E5eEEO+MAwH5/66oqbLmZ+TGmt2Emn19rsz6
kn8Ueo0yBheCOg5YTuRK3lEys3TqvNPqaEFTFvE0r9XtTrfO++KnZpWAiuiphhRD
GfLS0EL6gFY5t9rTA4Xl2Y3++gyHHlTF6bCmp86q+cbDOmQNkwgo3IH5HAUzKM46
Gs0KAGj670s+yHVP53AjFeBc0bXJNlbqSF+MWB1xiPdaGaH8I74MBHPiTxg1Jz7C
vsoF90Ivk5sn483cOn8hnyl3/44XpdK+9X3g9crhRM3HJJrnkAu2BB+DZ6mmhpjv
X88eQfk6c7xHXtK+Kgw0Yo+R3AYRDmkHcMJcS3Iys5XX933ALf1CUa/b4K0WXYNC
X0RLznD2jNs4kQx/XIeTXyjTZAZ6bcyhzuOfdFjPpdYscMCkvDri5EDRWmsgBwXc
0ZAGoc5/+AdQhORAJKHXAPCZJPqAgDfOkUUU++HyBYnSpqiTMhZy6+ZZyTl2o6yE
tzou5aXTXgcj5RbaMFz/+P7VC+Wko9J55KK8bby0mk7CRP9eNXDZ1t2JO41+OjNN
VoXCBH0EwRIRIgX3/NOvEOFCIEnH/WPSgWS6H/pXWqYlhrmnOy0yDEVfD42bSkfv
gJmRm9D6ieGtKFw5QXF49VAsQCP8kP+4f/jT5C1Bme104AgAq+h0zvcFEHs939z2
ErZaKqkkdFw7c+tay3/GeHWjwMxdC0avQcCwvZsiSt5z5A4JK7J/74dYwv9G5nry
S85GblOczaK3pZyxNyDx0mg1oAGd9Dsv3A26CP7dIK57dxWP949QWvVUs6JsN3Tf
TgL5bBN3fvPBQs06Rhqoy7NegTWoEFhfP9YknbX2ALkBXSdFTr5aMZ7kfdnc+9dt
4MHEfyaRcjoGe3jL9LXV9/fmz7/fvXxbs6axyiff+nULk7ou+fi1QLfoqSqeBWfz
SNDrF2Yv9wRaqskGys6cbe+BTf4aovbsRtK+TzfTN2fkbdmf9WYEdUGGJlqq5NMM
VR2IjNCt+1HB5vGUkNB+CVLAu994BERxZD02PHQ1KGaKh2QqZdP9xsBPJLqh5Oel
kdWbcaB3FI3OZnBNT2qVyD+R7SoMpJG+sr8wazXmFbk/ap3iXGnNLoKH1DWN6hl9
XNjdp1DG025LvZfk0ulVUtRLiLKzhSDf7mJlHm1rEfcg8AWdady0wftzww3EpyMy
DkUZ4kMCMzpaIX4+2BfV3eABl6rbHxlsyHvl9F3tJx+5ZTuBO1s5O7JR+HJiK95y
FhREbLou8XbmwzvDePmqmfs07JrScsCJQhWw/QN7SN37qMlIJZ2oo8jZl9XF51GT
teDT81Dl/Gp8ZqOy+IXhAL0WVwP4JJb5iprsj702VXpMfGYODQkXKI7S0u5zEyjk
YvbA4RA8e9+7NP2CqByyg/NSrcX+/CKBn5ILky1M1YO/9RLn1y6fbI2rsrUFWGYb
oHZqScFRvxkS1Wb7egDrbWITkYXT1p3ZNR7P8Jh8+oPbfzdsC4NlavwJXXFVjv5+
TSjAigaB0tztSxlCTB7Gv6SXP9iWuTl8ve3iv62ouB/NC7D5kByxTgN3yvdP4fWp
vmIyi+9yKNU0hDEYyFR4UjN0+U2W76JRsNyobHg5vMcLbl/AO/46xa/gFdMW1HEe
J+TQEyUVIOdHw0lanieaVzgb5NFuJLs9s+Jh8hXJ/XMLH6YwJiqlW/k9dB6pkIid
KjBpmPVjwbRh22P/kbwEhSxG53tzE7O/lg8GwSlgsCmltzjxHdWZcoawEN4XszaK
anfgrZUs95G2mDkzZAx2pW5LtGioyBcv6jUcjezrmDhUU+viYb0fK8BMSwj1zSCB
yyHo/zz2eeoNC2pNff2WGBRY6BwZ2I6ZDW3LpA7uGKNVUcMu2+Qn+AuqFU2B5f4P
0F/ghpPyLfCwU2uDXI3KA2+0E5QXJphACNRoWIKIhI72gbJ3Siky6Hk+hclnVfSi
RNWtgUKV0EJEc0iNnNcUw0whwjeILivo8g9qUGBOKb3I0LgQXA8UZeu64Hhl+5uY
gZYlOneyx7jgeg79QVD2CMv6fW44D20rng5b48A2IZf1xITCd1Kk3QfE72cb9Uhl
DvTbewwGbqSa2MR7cS3QnPfogoQsqaGTNEJQ/xm588Su/E8ywe8r7gSYTgjN6Ddq
1HbjPffvXs9+7hWvP4Ge3ixc3uPfEyyyNIt/bSbVho48ssZ2C+pdwrlixck8hVbp
STMCG9rlRmmywa8EDH6FckZMGTs1ttDK6Xp3K+U47vn4mdTfd/MKu8YAMeCR2rCr
Xs1IXqcax37PaA2h3AOYyq8Ca4+qMokDUpj17ZlBriMWXgiklPSkxo5HPZSj/9pi
fxFQ2UOY6JRN38Ighxym0apMtIFf6e/X2ykCvcdSQ2PFfeVs5aOXpX6Fkr1aEwrE
l9quUr0sBOs0X5blsIlOcJiojsecVncyjNJ3mUhkZyTeGNrmWUAGhxKeZrSX3VRH
6OlWzgwL8B0DtwMQxPGs659w4zNn1FfTnZzXP+AZBbSKkPrp9Skpdk4Y/fW36KWD
8pvMfWEhwPwTufNmZg1xRvmE85RQJO6tMUTK9G/pHPhYsjYNN6vCcAYkuxjyqSWr
ZLZ/1jWuaSUChO3psRLjcFieFh2tuqsbpNFeTGivfkP74VdXyDlRkJ0jT7ShJMYB
hoLAHCnT+qbAwnWHgeaqFFUgZMFeqdtBHmC0oksqD4Qa/7L5pLFaVWgDdBmPkeSv
Mk1Giyyl41qBA01Rzw9RVQw0cDj1yX4JwzbAFx5fQ8y9iBB+HQxr3DHLvt4EPLMv
Pger5FkXkxpNHJU9WE10ZvQ1uXJqkso9uESFAbNe+Xgk+cTgpj4rmA47MXav2hke
6zhRDxDgv8jnc/rt4pzP4tVvwa+NBu7/UM4Lb7NzQ8o5niafRddTJliE04tA7WHD
yMJjofpa3XXnUwr6ti669PSWTFx4467v23YLEWI363cpglOEWSo2PLr3SToL8pGb
HzJIxJSY4JG0hXEs6vZ0fcyTTImUW0qHJeMOPyjKZ3nL4zsp+hM398dmdYR7aaBu
ypOv32X4Rji7eZNbiaTPQSAO0e95hRmTOxB8Zb83fUL8EIWWWa2m0okWF9X25u+/
Je9YGwqiaJrotbMUgzo6O6pN4aS1A/vcqor4z9UsFW7/1VpBCcorWyZrRiCZ5D8u
Nxyam43uLa+tnt5kFQp5F9E0q1aZbhMZlXuMuGy3X6YiTRS9PfuIZoy43QHa7Zoa
TPWqmjTOCVWjuGvFzl1pD/2LqPOMDRqZZhTNdBwz+0VY2cT0ai9aFr3tqbIo0Pf3
Ljb8iquSXvOaz7VD43AjLcICkvhNuyqnH+9VWA5guW0opPWaOXFEffPQwt0W/DKU
DeCpQDxSF2x/H5+BlftkBe/JHAnSv190OkKoFJsBSh950Iy8UL1uoaqApr6N7lgH
yvudl1Objg6x3+cQ691yjq2HtGrJ+/E9Cfmm9DOy8wQjEVxeCfR3NbZGyMsWMSqc
dYHMQibbEvYikzsZCLDGizjC9tecKTFOM6F1ySCwkFYQ55ECLgHeO4w6aoHT69n+
03SS/xBZ09wL12KcyUE4kacsP80Tjk2TD6Df+fMI50bZXZ3gE5VcsxdRQgvGxbCt
WOSOUICMzFTrBCkI/g7N081UUE3JMaW7/Ii25HJjgZI3+3j0PJkRlyuavyWed99p
Q3PAC5trtwK2tZ6A1uIsLsSXVzcDLaAPxcrq9XxBumyk2Fi8XLowAAWCB/br1BVD
9VgE996UpImBjem1kjigfCwyCte3rpo1ZZ3egUxG4abgrvaYvQ01138ACjrV5rCZ
c6mX43cVwlBz2baZ6W25Yzli70ddsxf16ZV3KNUOA/PqCTIC1RYfMo3eY/ZCDYV7
HHTZRYGYbbhWW+77E2T3juDzruDIyqjhl+Frt/f2OY5QhLtPuTKkrBdD4b3YZYQR
hw0LL58SRfYoMyOUZyHTjs+Wj7+VK2cwPWgANz6Rg8UIWjiy75u5GXHjmtsyTITx
1LZ4urZNu8vyeNrzp/b3q8WEl6262t2pnTwJQDpb+n8Tfqrzzhn4QkPoHG6EzcaU
KQ1buMtsU8xUqOMOlsodQfNOtzh4NaF8zbYEaXxE3LprGckMiI45dbBNTyb7P/Dk
XSRDT9ojzmE4jVrnAPZngXhrmF+2zbRG1vu50gK4Vyj5OhP9FVYvH+vynSRm4Da2
6fdjt3ClW6pWmxK2WPf1EKroR5j0WzZ/Epc8WbCzMuDwRuA4m0A0kkPoBS/8+tds
Z95kT0+RRQpXVkZaoNRAAUj8An2xuJYbo+jayCQBEfbm0+5WkpbA4k6Sw/bbvA5y
Zj4626YX2txjJOVbwfaaVi3jwEi12ZuWCiEMsEyvQpQkIFfYdCLZg3wKegvOh2nj
P7+1vqcZrt68qWVUOEsa/99wGsMBFCQk/2ThrPNcNMZzX423HU+bWNx6IJbD/nzd
AnmsJLjCpgUNhYjcEvQzPtzVBaXd3YSZJOhZuIRyHTHWvx0hNxlGKYvez0FyWUr6
OH+5gES9w3JZ2JNu0yHu8D5cUKR7BWfLoI7oVJxBXzV5UJ4qAxwELUcCG6OHHHSl
jBS0MsXetR3mw/SbRDFb5D3OLhoPm0E9zdqn+l6/t4mTnXG2UQfA2r1tfr5NtTOm
Cf1jFUQk/crJEwbhn/YPH+OObbfTzpQqfBJF3ksU16nzYzX6GZVC3FFZa+tdHf+D
1GQp8qMVN2pGc0PSuyaVd8zoukTOtb6QIfmi9sPQq0iBvny3dRnPWUeieKC+HnxS
rcagVUdoHJMJh1IVoE0s1bOX6TzKHyQrH6dOMmT3/Tdyu4aYzYnmeMKQlZU2nq73
OGkHp+5QvUVu0VChdmyAPmNEdURe8esXYHgpKX58/Vshera+1f9KmMnZUdh33TkM
ZsAFPpxBQDsKOXap4DlDmitZe9NziwXWv4X9c1J7GoMRAWWlL2GEqcXunosKLa9q
c01Th4BezVElupJBram5EwizvN44u6OYjA3ROYqJAs6JnS4wCRrfvLH78v6WNsTQ
PjTdQ+D4lCMHSxHmmTTT08L6SnTyJbGZ4bKrMmec4jejtcGEyBTTtEANbewDnPR/
ZMMjM2HMn+pFQ3bo4r0GcuvQVqIf/SxUjr9JULjzCMFWKKew7GkR7SpQ57pBeKIH
NFUSwjF1+K7wyYOuPIthB4D0ACieuJfNQ3QfgbBSg9CJEq1OpiGGGPxRoQ0Taxz9
RjpGYqYc0FKKCOogyAotZr3HZ8L4bAms5EiyTyxPGBo0J5S6G2fsKeq3UCYOfuHr
DRc9jUeHZu1YTdzhqsXZwpIn9Zty/V4yIjJrxtyssa/SbEt++w37DR0vLMupngYg
QKGmCjYFLFoKc0fje65EY1Vp36ARMBnbR5XRck+rrLRgezZa/cXnubkfBWHQTaad
mAnG4uy1GaP/4tJNAkLbDAtmDhvsLpytMtxgKlZOFTGHqfU/KQ8C+Fo888CZfJ5n
NDIMIRqyxHUQS0HLESCYEBIaDqwYIqv/rMjySGcaXCf5qZ5mv1TDtmMJ8HGkB8RF
YpLMCVyc17KIGPv3fh/Qj8otughQgAy0EIEJn99As4Ut/ku3jUzhzmLLE1f8uLY8
WHntIFtHsjvENGiWqoBQqwDEh1zL+u8RNNG29lNjnRGwjuTqGsxCtRwj+YrEqHCJ
Xev7gfavxAPHpcVZO5xwAnAb4NoYXVRLvYnGG2f0MHuyENGQPIHGaBD7Ok/tuGIB
oNvwOalMWFgXVlEQxHAqxi4ga6trDOPWcnAHW3E4LguT30brePT675qzl69rNCjM
r1yk7F5BNaPTZhl1JeCLnLgWX1HNLFKClmSgcVq7i3i+mB8UJSY0aMKuBbszCQY9
eonXbNmzItLagndTpwepGnig+21YZ/sS5VcLkuJyFCo8z7CvCLIge0YRPjXbA4m4
k/MDiBoBUloiEtn+BK2JKY9FGlmF+SdE9xeAzW+O61FAY3JDxT3XlB5WBYZQOzFD
U591VAXTWnQaFnhzhoya+phDVfQGX9y/WL+aDDcXOljScF3nOeW3B06btyJ1OgpE
fEp6rUfJEQP7KZQkcja3PR83bAwTAaC6rWdQ8kZ6k3CkQaOwLao+S9OBkRBPYcO7
FgdKmoPpYoEjNHk6WCVWASbTWP0bct8dVHBHOvZG5C8ZfkmdgCy1nD4jsPM10eoH
LqnXU/R1gRWw/jOZDI94wScv3/9JzmWPsJz7wHarfC76kwi7qRJzhzBKmxlJ1d++
JhzTew2aRTYcePmflPmV9XL5I+jzl2ix88ZyhCvXQTGvBp1LnsT1nocvomRyWS1N
k7K14yWh5dArKxhiCCA/BNeOOpQdGMIMjbGNu3wqYT6jTV+huCrnS3OuLA/KFGVH
//LzEeAUKDgEy7+OfbwkNYhpJd0KJd3+nahW+4mtLXK+aG89gQuNBpUVJlzp4T/u
nd6L4tygmWDaPKywnldHsFZ2ZfFMXeB2vVkdO+ZRW9GbRauV+pldUvQsjSUAE7zo
3iw0X0cSD4xaQsTD3yMbWm4hYI2aohJ1BkecW8ptPsVE/+j2HrZ+/HTjjJECXgTK
wRtE5nihzATLCY+jfMWK4l/vAq6XAE6E9qE30vZunuH2wrjXIU4wWsTaDbQSrIAc
0kDCcq7UXJ2SubV23vPhu7BLkG+ejoZlfyRno2FQLmVB2KTHfZsOiznJvN/9p04Y
vThpUgU+T67C3BjVrK+cAU5aw2d7V6HE27VEolJNgRsC+QjI5yfPYal/1O7++zem
b51oJnd9wjoKlhPoIvQBAEhRMEBVPOHUJJcAud4XppYSVZOH8t8U0LCLBCFBuiZA
Cdb1IqZkx4h8g4oDUQqZZl3nD71Y4LLC6bXylv3HrD1b+2OALoTlf4TvkvkjrnNi
3MQz5QrDTOw0bY25aGMYFvsQxWBjfWNkfgZp3H/j41M/CbDYsxkyiMy3Ked6hlwN
2wKx7lKYhoE7aljCsDP+VRDZAFP40zrn37aMmfSmiYWAkg/i9kjU9B2EBLjFrTEJ
y5ahovdGfw3wy7s6NhQS0ukuVtytf5h1aJjHniwryiATcgZEyFGw313Y9LexXcYR
pRPr74sWi9atmHCxmaviOcERcnOp6ITCRNVMKN+YN5AMUZ2BfhSE3JAy6p2YoZHR
YICPh2cRUtBm+9XL5fYfEunVs4IwYQVQ+Q7mtmC96wnxY5QP/w8q9J2iGv49Isha
NL6YvBfN49HVJK6J1raT0qFpQlw6zGU8cvmaudrLy7ZomCoyRJ++BfTi9z2LkQH8
TMjAhGy9cI3YWqFKa3GSLGINcCP/VQUOjD4TxjadCU8ay7I9yCQEmTNZdtuhwBaj
ViVbCeT8yW6vE1aBLtkos54Loj1lCmFQeHt3eTLb2a7FNmMYJxOryuPuY8W2PFFC
mgAwzQDjXpot7RSVNZnHUUJufu21j4c2CRm67lYFBfnW8Z1GI0lGf0QsbjpzdgTm
5vVNuSGCJFDGP/XWI/M4kAkVAwitPabqshoBSoYPItN3JhexYyZusyn6nW6a9/cE
Jv+oZSWj6amwBs1BqeoCVnJqkfJBVy3YiUVgneZoImoNdok7IM4BXZptoxJUzYGd
rspZInKzowAyZnjXDaLcfJ1bPyFruiP+CuGRtItdiWxPU2sk6EcL+onP//nmQKLi
ZjYIgi+DEslNNsykxvAVC6J4hwMjo4KbpvUiHIWh0jL8MFYlmZiCBVXaNHr2loOi
1jNmI2TVf1cLjFdVJnOzHZI7ni+eoCcSU2DVCqC4x26RTJelGbqCPxJkg2wHLyUo
rcLIwGVyqmPGu6oQQ471PnYxf3SAHRbQZnoegNz6M6DjMOJ/15ubaSR+t7E9p3R7
smPcKyMjZKiVxgqTxdwZr9eJCqySNZgVzOcb1rv85fPzr4GYJr90AyYtXBEVfJpY
t29eSxvr0c3Yr0piSbo5hUaGXTDLkHgcaJF0eZFls73/H9h3cq5058IV17N+PTCq
9clghdCc1ZwBogvzYAliufhZRhH22NVlF5u4ARjI/lFngO5TFENE7oys2cidP39Q
sHfmCiIp8oJ7l/ZFSTWacsBmihnDpzgT7b4lb5tqkEc9Dxbkxi7UMFlhVeisgOeq
OitQRQy/rmpN6ylTAdhh3LqgROMqO8zusjpNZiCOm9pnbYjOmkoAN1qWw2ENHpBu
4l2e10i5XQ5EbwGMa+GV6tscEYz6j9F1sh2PUUbgsP1fPTUhhbMcnoAmcybpzn6y
UGb7XpPxGsYxMyuGC8PNvNYJI8yYw/DMNedl5QTiGgzPCrmKMnDcoP2VMvXN2/AH
QMsEY+rXJte6y+lda7R2iZF3nEqezT8pwOCeRFu4xMxodYsgej2F3j/sIHMR1GSK
ZakLJmpqXFCpzt01jo1f2QBTZa1K4ammtR0ki7oGxStdsWOATcKyc4DDsKOChYSK
/qH1GJ2rqGDxmUXI2u6NwImKt4PNvPiUT1x2weFG6bpypwzZqFtfWT2QwXIMOfZl
bdfjmk+zuBh9KozCJckkh0gdPq6Fq/ORtKleOAp8joF80eaj8pAyXvAGQJIr/5+D
Zsg8EjfxrdVpEZGZK0aQ6ldcz3hua1JuraJBVxBj+6rHhwXFlB4OuVVgFtPspvzT
oZVFAkoOSq5dTrH7pCaZCI1Qd5YvvoCxUPkfGe0Z5gZq36uCT4viKa3yGhDAzzgo
YNSUfyf3/T6ejfg7wxHmrEx6xsqfmmXLimjbq8RO1us0jMFUHUyhD3L7U6LwGF1p
x7iVJzU26TCfMieLxWnmR3nH8yEL9lfWsYAxXo+coAWfQs6n/GSGvEpW6dH/j4cw
w/fOWfLzkijmmXapfK7yjy6WeRjdQ3qt6kT/qiTY29b2ZorSiA9YEvczQcgARekK
vdf8PWvnp1EQZjpKpv6O9WDWxH41gs6pNY8tZZXlClCQf5n8FUkJbMd1korJwase
4wYa9ILCGLPaLHmFWifrMuO+06R/u6EVw8ygXX9D2BQ5Pg+pH5xEHj5M3uD7gkdB
XKMWHatfChw7Z4QRQs9/Fw7fiy/vIb+YnEtlMbfzbkYS3HwnWfRJDBGZQerbXBFY
gy195IzKq7E3Ivz8xUaNHezVeczFubB4B02lPKBCOUV+A3W74ANUXn5WcJ2hQ3yQ
URU0ieZ6BWREh7Q4vw1MYULM2ubfq529beoLYrCzEkrpfw/QRSnRpiAmzQ4/HT1Y
ymQU20aVz0QUafbZo7Kmbv1RK6zgdLChzs0/8Rch1apnYEnQd+UAvCCD/hCQnPWl
6HTnYm0LMuvrZxo+dENHGhliOFn+QcpYS0Jl2gRatSpE6kxhEfTvLBZxHm9RQSoH
xXERsADWicpH6AJ0XBTUyfQyxdm5uW0zp/FFXaUjhOIxZpARnyPQwc7DARZFg0ut
wTvwP+t1WUq57GjG15dFfrNaOSW7no7VXIqpvTmcu6ErNWQPWKuRED1zhb+zHDuC
UY3sCJQHhv27mrtmK7++7QdatarOSUG0ry9N7kjUdEwNDavekwxLnM6xVbbbDGSe
LY5T+q4fCjF2k7FYRM95h5z5ygTFzFa2WjS2FbzLR8Y7fvK4KX1vzjseMqABQ0Iy
JzCFEJuluni29UnKdNP5If4tubxsy84IxlRFOQp/XqjhJugIO7ycTW9OdaGNw7s/
Ga8ArK7tlAPQuc+bCtQLZpKq6zGFDYvngQr3rQK65WFYhye6cqA5GPmsacUU49j1
nStw4j/MHfmVrvaF8eeEAZeflyPGBLV9JkGarGhv1XU8dfrDsjUcn1+vAIzqzTAr
bJjYIvkPTPha3smCHzG//Z4aSXRcBiyQPUsxE6F0B32VNf11TGTKRF9UkglS7tXv
Lp33M0ZC636qKqXp4rVvlKeqDFJfmujzSRSmA5HP5Gp5JTRDB96/QyrJ8to3pLQV
KBUkkip08u181EcIEaWT7g1i0HqC59Z9pIByhMKyrptdoPgp2cQDR2Oo77ghYbdP
qPXe1TKeA60O4FpKErimfsou3VsCCYu1bK3crnfdsyyN1+GXa8mFtAeNTK6tx7bN
1L5QEw4m7G3nVNZA3EhfuI4cpKFI3uDF2FUsWpGFc7xQ72t8HfvAxGY/5jDSjwsF
fvIfsRPq5xIVtfGM4AJXRlQop7NZkt/NKKcMfENROYsKMneLaxmMdaQc1tzFaySY
D7L5wxf0bLcAF9655YgmQiwb2D3jmsV3hYlr0oexFDUZCBpyBYXRM1BpylC2nYmD
DPXTVlttH1IvvZY0NeDFMaNonoDAO0/hVVp5CgFQbNJa9yUlMyTfHrRSzX+GLS5O
8pp8ItCOJj6LXfYPYp3k1GS1ZEVKaECnpmbnnOX5pNLq6aWts8PZwhzY5ZCUl2Yj
PHbB4H4dDmEVwTYuej0vENQK2pqWA1MypdAHggO501FYQdZAPl1v7uUidNEHRCR6
b0uUr2o7234AiS54ts+W5WVN75AcNCPHkjkix44Jou5bOi90rnXcRZ0tc3mzlG0y
QgxMMCEHC4YFPKzHBXcU41zxjqwSsWbYtHpIHZvlRvKd45DhRBd0wuZw8n3zdqPN
SKkqEBIsQdgR1f3wVkcwbwkdLqxDyz9LVRQuz2zZuGtFzZQeIl5DUcX6NPgaFkGA
fAhzOypwUDRhwSUEZHZtKI2ZJlXBwYKtVXMuB9AzzJ9WUYw7zEe6PXvNMwwQQnn8
kqWx1rga6+Hpt0U3tWK6Npmlsq4oMgit9e42Al0qaO7Fff6VkOF1h5hpQJghElSd
czmMjNuGk95gq914CP/wwHmMtIQ+ke3ubAUwqDtUzu0leG3VP4nX6D1fUzRuYHdA
in5RjrkpfINNNtzmx2xLpHfhtT5yTiT2wEOvwXMtqwXKQ0pBj4pH88RlPzYdHl56
vFfaEBVXwEHYvOiLzgdfmlqViCgHbP8x8pNgNespsyUanaLj48dywFdsE1a/i05S
DkMoY/2rg3EnmRYPrTCAQRnRtFghOcNjExWsleBGnUFt6AHApSCCNruRcR+gTEMh
ru+Ir+oO7XjRg28FIXOyUNHlQF3Ev9mROojKyE2rGHn4l+mrmoI4GTcdPcnCHHna
3SHCXbcQ0U5nCtOYKRieomW8TOTdenW44I6vlcqBfOrDQmqxFLW62bEtBTwplw2P
M+9m9Xxm8Ebu8P6Q7NF5Apm6KC6Z3uCIE1L6h5IVhk06YkhFZDhzuePhc3LGM3Vj
JdrQngrMsqB9VbDMNV1cG8Zzi+ph/8Vb/EnGiWdgtpfYctJSS1gdXsG5lHkjXf+P
5i911Fx7IwhZekpOn4tXBBFcw6FjEynF42K5ob7s458NhZRcaUlRZ+c5Ra4ozkIR
PeP+vhIY1GISYIJWwltoeXLgK6XzNrzORNxLYvS3CVlgclB9AnhWEkKPAFDL6Zn8
3Txxh56OXtoNbXyXqAsbjyZvcp4ZgzhbJiBGpn91Fy6LibIysqN9Ju/HKxSkbC1a
KEGK/M4FoPA3Y3CuUDQJ/GGn79Lwd6GAZ6z2sUOr9wYsW7YY4NyizIirVgdR0sm7
gbxrJRJNgWOvo3V9GigTe/suwfAu2S1C8Y8MuIJDrsHd1xrYrk2TMujinKq7hG31
yRlZ0h1ls++xZEV+DfEIxU+a84T2E7psRgk3kXYOw1pKlqMwt7toEetlajk896U3
+6XK0DtluAgKwntJhnBrKUO3DfgkrCjuc+YAeQEFluuXnloTbWYanJGplQSIUCoY
YPEc8aKzYuP5P8WGH02I5X7wT2X+qaSF0bNP5iJjppFhFdy49CWO40kuUAF3FFHF
ErPx+UC5t+YgVYmG4krj7p3uD8wGy49MGQyxl7FMUINsqyCMxpZEtCeWIxzpGakR
zO8OQngV//qkIx42dj7/7hVpUSadbKmKlAuAdc0z8qwVCSJDQQHU7TsAqiadXcsL
O/zahlhfpajHAKT6WxylzCmHOuzhZ2t+WdctWmai+FbRPgzd5O8wGraBFpREipDb
/3GoBz8J4GhxqlGIJzu4rz8m9poemMUVSsrY19lpWzN13cITRTMd5d4GLmycYNzj
mBz5vUFResaiZkKfIAORqFcoKbH94VcjIyx3SCtG4fYZwk2IARIauGxeuuXfa69o
iSMBmDwkBmCqc3SxUWjamBv63knMzVNXyizalBLm53Hiqu00aG8UZLFbOvQR+yjp
KPDWzPP02CqIeVJm7cL+wKrkC6cM6dOxJxSDaKLsrPpuVN+DzeMtp2IojZ/DUijO
H2OlZh4RvL85+tGMAniwS2KmGt22u4WrJFUA0HiZRP8mUTogHNBNdXNFsTG4oHVF
L4gjl3kfQ7+Ehh2jHa93qXCPv1drRRiBlBPdcrH3gjRIpfcgvYIcE3T9zb3k6ujt
x+xfYVCicFsNc3lECkgby2mH48Lm0gAF1VTXEhCPWsbqlB+u7s10/tzIRDxygtGi
cQnX57brXEgN8trsp2veg5ggJrjg1nUkFEnNSHW/HBivBfUXmQ911ToEJO1YD65N
1Uhi5onPuIMFT7vOWau3+FTrzzfzWFfm6oO7QINNmJAqcZOj1PoBr1GSflcQPSSa
N/6IKmIAgXYRb5LDIgur9q74ccAx3lrJO5a3Gj9Hvnqzlx0wPgL8vv3hNsAi0zi3
XLnUGAOsG6G5ho6FGOdw2TZpLMVT58kXSFfC3pHI4+XS4h9RVDkgcQYutq8lGkfe
9nqV/WTmw7YRfknc0FkV+QXUnx4L793Ve/ZAQgF/EKsdKUWwTCu85y0zHSoGPwEn
gq6x8RJudS1vI6gbUw0gaEP0B0WY+zCsEkXbRd/fkGTbRiy+ml8P58oMKYyG6cnh
c3QwHZkK+4ACKOWJNysG51eYQnzzZQLS4ZbjdiLL5N6iNxzVtyZWSFfGfXKCPi4r
JTRAm+OTIXXMa8H8fFslXytlG81t55KfoeCMRZOw8tuU0J1P/VcvRCGzSRRRvdBF
dgbdyIpYqRTbi/QJQ2GzWaArQ4FcVaKg2OAuRrZ9FKaNBV51ouU1qgsiGi0WSW6Y
LFnHc4o4Vu6K4QLYvB29QDQdfpRFNoZLxmNLK52aBH3CmJXrgi8/WoJfUnPrYCuR
WY3LM+8XSNNmn1MnA3KOsVSaP55X+IUwOnZI6iGuS73mcsRGQp6mFusexfsvYnWI
fs5H3mHPuanyT7T6AVfkQ0q1amnDfrxvwMDqa/PZdukSwYBqpsjgNvSNhyAQolEO
dRAEiWmB9nK1/pJtFKoSh0ZDld4CmHiSahGzo+F7XCMrZwdjLIPo0h7to/SMz4hX
RwJGEeX0U/T2vTCcScQQuyFTX5Uz7wI+5urm3jGZeqjMH2/JN+V33N+fATUCptMo
/jsck2vmL129gcqCqq4jgDDLFgl7Sf8o48hT9dB2ymCY5dl1LvZc+yrE3eAPNhIr
piv3l0cMqDRQf3NQTTFb2XyDcjyNSK5UeyQ2PGRPUg1K8LqwaldizCG5ncGwU3IX
/fNfsCzG2KNwxjk3QjpSxD60s9C4pYPLmBu29dfaswMAaCaFMGANAa59qNqrqbp9
MKykILgQScxP+dt2sHY3P8dTDOnrSLcTrN8vr1PLv6dZSp6X6kN/zPCh+yTB9WtH
6ZHOUZtvEu/4pOTCQrrkfOblEEFvudZ0sMPGlKloCsZUE0/26hqSfHorBivPisPc
CihozCe+otykptSe+pERihji53ApDGwmfTlxfKkc/H2qF7pB4uAN/RPuwwkQoKLD
uqJUCIYYCfjy1fzDRbDbPbhcV5dbTcS9JzDQgjSK7+vt1VgXaulxlqIGrYHDhtfi
yLuD3EIsGxlkYEIP1LXtX01p1t4qnyiARjyDaQZdzjRGVJ3kplkeSv+co87ADxTn
9TkZY3Pu1Tf7xmw24Zg9/c9e/czn5iXCinIiooAFQMXaXLOgHC6fIp5ATq/p45NM
nq53oRXMqTXzPic8ndE9go2OcGMq8p9rBJ8EcgkWi+e7lERscgUyMDK08HQSOOxn
4xja5LsyGJtfwOx1kIcDvk0L95uLhcC9tA3ZTGmVTOy6tLcgQvLRuzziWSkSPlfy
02Zh8lH/eB46EevGFhovh1PJEidqG4clpwKDC7+A35eDBB57vXfyOBzi+ONAazw/
Hd1s5PK22JEYMDTkv8IjjD9yZZf57krILUvjNyVbocMLcBjwTOxP1MHWh1wUUPWA
66XvAg6G4kCW1IYS3gdv07puOcDW38EZFzZs7vcRqkUE3CKSkLCAS/h4vCGdt8DL
pzpOR3LOBPvFNky/hn80+7W0S9ovc/tI+PTTmuIyldMMygRs3i2LfpNueWJ9lsgz
1PojUKRQRFPNUmLaxRKaOf91vJIMSID40yN8r+mOwrGXp1qN4iVIBZLuXxOWut3T
MYSCUTxTkiC7bPN9/qoHcVPwDGOrb+GQT6E/9wn56NrEuvvKlTQISNiPbX4AT1xm
70OW15NkKS1bU81bnNaHP/wqozba/jSMI7VpEUr2RX8iePxqje35emMGHBK5NkES
EPhsYIE/Gasf+OeuGvwe+XAES+f3bM3pdE2vqc7dFy5JxA+KaYbgYgX4cWTs7ujJ
eQX1EF1iAllfkc29opKoWfd32k5cTtCwhkPRGVv5qeleCxOxt6ryrIRq2Pvs6PFm
muEYz7MrKQVZfDY4Yi3pPXDAOaCVMzSL8W/yW1lwXf6HBg8MXy/SIONGzvt5Ii+S
5FXhhsso5wWPMlbhf7fkmyj1PpOye/fBSeohKZ7xadOxYiMUrfOSPuj9HyIPjhQH
tD7LWf0wDeZBsxIJLHzgrOL1UWYWap/Od4mlSpofSHnddVAhYTFU8rFGFZID6g6q
S3JOP3rFIMGz+z7OBjJIIWb1dZzTX7OhjaADvGIP0dwNF1O4b/pjSdqt1Vaij2LD
WxEYeJOxKSFDa/RB21PXpWO4H5iHFiMLMn2wToW+KK9olDeN6pKPofoyNWXtr7HZ
ZwWZ6fPJPDkn7IiYzCGdkGpTwmoCG7Ij5TaTwaieYpwBQEkd5P9KdcJ3fdo4qRjj
5XBhWnlnhzJtoBW2+SdTU0QnbzZ99a6yxkHUlu6A9Am0GkVJ2APEp7djE0NwPnC6
ZsX1CR7P+mObW/38pei5HqVVLVOqtiPtxy5gFnMlM7yDvxkfR1ZKP9OjGMhKe49I
zfJgFWRNJlr4Pd2tb3S5T+xlMMb2uWqCB9sB1CiTSFplUkcknBjIK4xcjybbtndT
goZhT9fbVQ0AjiGlXJ7QhqvIfYUBkH6HZ/fe53tq0RsR40lJqunNZekyV14z8dUF
NPqTE1h8NLM+UrBmfHdjOdPJl1ePo5UGzR131YPb8WI/pqxkjoa/HiRxwjY0i47O
6t86UXMpaent8oB2O0Z9g05NMcxvEFQoDSB4mETrUNF6PtvAjoDSTso0XNATiuA/
CDEDf/0an+SFvYlW2gkiUmwQYwHvUxCpDpgrwvvA1kNz87MY8u2vpCAMrWd9ITBn
kpYbrqnI4QvB7t9zvbMREdeLOTkD5AxXjDSuSLKeb0uMA3z9m3DPvemJ4nAUMt+h
xNyIfImy/W3VeGyGIG6oaOj6x3I9GWz0SCrOqPrfe3Qaj04cs7rMKOZ6rsdmftHF
CvbEwf3ohShnONeTUJMqQPEwIlq6xAzlpbFqgh8nOtAKFKAsEefT+Uxx+oE+hZNi
S3CaApfbmT2wZulNWUwmtLcuUb+u+y0Vze+159i5YKVvRr57uopJEYC8X4fu5CAk
QU3l+N0UwFMRsUA/VNRRiPeg8p3Nu5s9/rrXk0zEPyz/7i06x0a+FTGDBcA8ObuZ
8VjlfCSKqLpXgZxIuOp9d76kfwlrqbiIyTue+Fn3tkoHd1cCypNPC+LheA9BpPLt
/3PoZcCaxb0yqqI1gWpS1jXQn7qWEGBwLiAb42g68hKbttPonX+24dsniK/C8Tw1
mrfE3ik/HWOMj7AvOWQZbqhBR4lxtJkLg/KZO5iuc1arYrSUdn+7NPAD2X6fHoZB
deSDBscW7ujND4QzuLwkzSxh9qvN2pvoyghZvmVg2i5Mmq4utMQeRcGGOUlY5DbO
k4JLSk9uykPuTeswP0KlAh4kmv1XtzfMEsgyfwei2cUpzsQRZAK2vuEJ8XP3p8xZ
jAL9VBlk55SEz7N6Mr/1Xu9QpKf94kSP9zogetQgXGoVbOmcB9jMaqSKWzwa8xYm
mksixMwOs2utVmwRPHEANaV6webLpxIdkUyYauheMkVXk4dtxfVc8+95NXMBL5Db
VRda/M2ePYZbwBE0nOKosQRDTMddHGZ072O7UsEIa/CT4hGL9GDpPNwJRMjfIlUw
4VsGsQpRL/y94+d7i1Su95cBcLjSXSEC28aTyvIOdg5cYp8QfRgaiPGpf9rnUtb3
dsEsv6AcXiFPRrVREdQ3/fWEFx17ug38VrsRsopBFmwTrPwdbJmoFn60305ZoI/P
CDHOMjtvTTVsWo3ai6etqzPbjyFvPn8Fj3LrSBQEKrfE0a1Rv4QvezHas6p22FA2
DPvAQDbMyLZN9e8MLNldRNOX39ijh6bTdig6C+6RF/0srOClV/2e6DcELutEO5xT
e7Lx87NoyfCz+43pK9z7MJvUjAaABinPUdCVML27haCfmtocGFsxRZocY4a+tWtH
1uos0uxAhI84VQy9EK/nuQlz8xqlLcqV0tJYcof8ycghA1ljYCp6tbZ0T3DaCI5m
lJGBC7sSLO7YBr+Oh5tlSqttjDUrIfpxAkhUONYbznXRXj1uGHMjfNFb02bshVRH
3/HcJNaDDbqRB8bXq0R1bUd7xRCwW9Zmep7EqKw8O2KAkqi6/dH55pDrv2tsl+CN
ucX4lz4eqo4+Jb6eEuP/tkT2o+7rCAd1ow/W5w8t4QilXszKLBfXx6xGB5l3ixRe
rizcdf1W+mtJzIhvNvzzducWUGfsYPJ5TdhYS7ETxFnNRWtHaiHNWptr5EZxdG4A
f1vITdCDkqXxgeZjIuPd6PRWbB80e5RwpTrPtqfX35sCawrtRBIqVw2hnu1bm59u
Txyxno3wWfFOrv0rNWW5LxX83vX0AoKGSGX5ezSAqyWjf3/xoRMk5ydNTsmZfvUM
gjVqR1YJiO27LO3wCypf/Y2BwwfFkTHdiKvS5QLd3uUpYrw/hiWPFsQEd6+e0RC0
wFe6ZFBQSCjp8RrvRn/kUCrVbX4Fo+hkY0fJwdyQeYee4yYtpE2JadVYCapk/Sjv
3Kf+yLZYSLIXRbNJvZiaYluTf5cpd26+5eQiSMYnf4dv7jWIKkGm/JAT4IhvQtKT
rzAcEKWbcDKWfxSNr0g9vfZuS+lBK9X6GWrtV5G/ollf/3vCyjz7XvD3d/Tr0nnG
llm29c33Fbs9Q1Qj+oinE1Sj3z2jJ+eT0xQP0oTbaa4A/fALYKK1/p6tu32pnyiU
lR8p/oqOTbAu2dRygE2RypOoPj1skqHXvomEFmnkqAxEFNghS+pFQ6yG7lWPu7Cp
Y5w8gz+zMqhmR+GPjxpsPidlI0o0gtsSYWsjrudt3TVB71lqX0ekv7jesDnhNCQZ
YicPjlknSd//qb3J5X2+6p+f8EfZrn5+m0z7OAkEny3Dd52rh9yW98e6cl4ecTj0
gZKlypJG9ig/k+P9wNC3tScslsLItiidA+97BL+V1H1hfNayW6gsLKCglM6/Qb7Y
rQs6E1jhuNCE99dVss4MR137CxmBmBUTjSg2Tj2j728wgorQ9cT3TVf+0vfJ0vYi
gtDaj9AdC4C2KOVraAhfSg798dpBVqPIe+SuGUOR8ZO0i6zYrzse6P/FpikGKUqs
au6NNvtubwfrkmSlIKs6iCFhziLTnVkRaZf+pp/lZV76hb8KHi//tjzvd50qLT9G
ucucEtkQWBr2cYOaGx8xXEeR/PmTHJ9PPvvNjezAFwMAWPdXcobWmAn5vj9XV2k8
MpM5u99hVLM+3uSuh04Y9M8yF6/hcm1jCRsh4AdU1eIt6pJzeD7vIUiqUYVIEUNA
RyzGJkmuaAY0czY4Jq01wo42TdPvIiOHec6X+HZj5bJVhf1trMO0KDahtWtqU+p1
TyTVGWvaQOeBoP4nAlQSWYM6olUpHU0hmL8XW+M8i+q5+2cKstlWUiwnBBK3FJbj
lbODt5nXCm5G1GNP5lRttcahief0eV4eUpCvSGsUR6iVNKzjHigbd1k32Mz2Xg73
NKQZqZtKDXShLtsMhQMPTSaOdzI0/tPJhRVhg7kAbnfcH5nuLRN+wbnQ0MZaEoxF
XW/Yg4D5rIBPqOIogiHGA9s9FYbEvkGy1gNGFuda74DjsAIJM+C1I89UD2kE3CnX
HjuaquIeokqC3hrYDd8jqkBowGmzrG7lC9MvDUBVTBF/1lQ+2Fv6RBdpi1G7f4ut
b4jgdeEkvboCbqg2lWvEh4QyXzibLVzVk6iC5Ak5s6LW0xJkms6i2n5a4pXLAOBX
PGl+Dj3JGNQk/+QET8md/AQ//ETHdwVL72B8zqxcHlWrR0LFrewmU8q/hl32Boc9
HgBFV5I4Tud7msQZVyz4bML+Wp+vNv7SWWoex91kbV7dbL9xxiieLraeSJWoJhzl
hMEH5INHyl5F8Ukd+9IXhc0DyPKqskobKnjmcfys9qgS+PitVENUUYTpIl0rP93J
Y3gAkkm0p/gJlS01+t/vqQKhem+TMFg1KXiVUPhVCofFc0vJ4pCo8RrZuDxldEdk
0Wr6+WGVBmJLmD0oGCeI4U0hlshkhHrDAC8FHkll1rpvL6uzGXJl7mM/s90gQTmk
tfzJKiJxqqkgrIMZPd5mN5S1Cb/KGPb8bGNV1k2CMVJOga9rKaT7MdKGzEe5W5fc
KTez0u6SZ1vXqcSVUAE2uFqqAqZTbfVvWQbKxGgXfBcQGsD82gW6RtMichr+C2Vi
3ggcPkkwaM5IL5rkJjyHw30g0MqVHlh09mMqixoJMtkc/Iayh8nJ0HaOXpTUCGZm
hBIFFUl+s2Sir/hnkfBfo+GUONaNNXezqvvj6ThMesy5AAhL+zmXJTcDRtgU8u2q
WiTaSwJeOgIohL2alojLf1X1eRbL1dtv+EaTVWADBjYYBd8OkFzYWJOIaql/VanE
CYpAX1dfL38XjgcmsvdMVvWtyZ4HS4l71lNHvhgUvkpA/lmvn2NLY+SiVvue2X18
RXDTHb8rhGavsq/lEM3uWs444EQkEXA0vnK0ibX5CUjiXO1jLsmSNbqoDWGkXMYm
V0Te0gE+63Acjhw7oN2qZgWZywaJAXTUwH7T9s8rtAz7mg5knVLGxs/HNYjwrxHM
/JaRZd+HzwfJMliszrbJOgVqbUBhdBgJLVoAYzP9HsxpgjlyOvE0aFE4mzvT/yj6
RkuO3UYZ1jHOXMquJqsGAB1aTDSyDh4trT7Niznti3NCUfeyUU1SPW5rFp+tTXy2
Z8kXktx8uShu8JFZ31YNGocLZe41/PCqgvbRWV8WVufAxOz6YHvP88bcQsaDs8kz
hw+Y7s0mDMwtPbiA0N6Ix9CF8JfRFUgLeE5gsTJ2mBJ/5X2JhHML2YxpYbK3v8Bl
c/6CSQdXYoRdz4O7t+/lahXmg6aM3L/UM6nf9pRhKVHijuuxQ8VDPfjTZ77F7Vuo
vv+oEbLZcoPvz7MPOnzZBKRSPgbgmYRnDqe6pik2DMloEbDtyuP7k3RMoj0MgqFN
y/8eCd3R9MtXIpWirIBjBbHMgelbaHs5YClGj2PF8gjzXWferOyYEp6zL/cxR9F9
J10kN0FhKFg0KqFESNdY85yAOlpxL8cqxP12nPqaw+sG1yAy6Qx317qPtgDwE7IL
5GdyTpNDDivhdFeo9GEkd9sPeXvs/Y7TLCsY8j18D56OPXjYQmz+KgSH3s+EPvBQ
YuCjPf9KwHzsWeWqxqV3aKpsfC1yHedDxFXW9OBwoEQxk9b6APT/gwBEYBhx2MAh
LgwfY351/bUNx8U5uNYuDCuvxgi4s0cIpxGMHMgqSKp+CksWWBoA6QfA9oGfRzEB
LYiiFk/Ry0nVh//o1OD5clEL/z3zEtLz1h7wJuPBt5NiZaQdgnP3hyzVs6cGssUa
V5BHC5adxT4m0zB45IQV9RcWIOyZjosigY7B6/JEOQxXRn1sUgl017kqjoGFhdBz
hr/ilvpZagOMmOf2Ysle232hqIOW28UEhd/NsgOQFaXjfevV0WSsmhvzosqoI0iw
87Zk/SO3sH7Q+UDrQmW+BF92nMTqTGy5KGjCB4Imw7t3u/nUYSJ12q02KnXsK6Xa
VCJtijApU5PdYR2gQEtNkc10xFAQXIKeBOqvD3mzVviRZGM4chyJ0valoShz6jxD
o46v0N2ZGXPHpwpJVwN5dfZxAIeWk1UFcXCB10K4EG/TVzvO3N42Az5KCkIR8pOt
IDM/O20/eKk4Hn/sexysIbybBYNb2/a1lAAt3JRnefl+HTaU/FYERg9dF+7D6/Yg
86LJ5VBa9Omzsy0pPQCxMUFycJ2EhTUZo35QZjYvLKml8gmEz+5tAWirPKDMG/e1
5+TYn9l/lnyHVzV6DogpLVRIZ3I+Z2U5ZBfvebGntydB1L8QPkCgdzhOzxlQN16t
3ArIoTKeEIPTPmgz6U3/33U46Tvfa7TfmYsRpyLpY4EBubUczgbUmU9fIl1h+VPC
GOy+mpXwUhSYlTD9HmdgdDPFvUME7SFFiRYXEr2+j0Q3w2YL4d790bgZnNvlnkmw
CXcgS33A39pk5VQ9RtNGSfckQtr4I0lOwg1xJv8DlCkpuFuMvdjFrNz1xOkzJbcg
J4BaYm34nenI1mbthm+kvedvVorDRtZ5ks3rDWRi/Y5K3BBdUUNCA+d+ei0T+1YE
Xka173gT6xCoKWFCU7YZGt/+qtstmPZZDALprpnvCkbLuu/Xa28ODRy7n+xmv3e1
cr8t/jBjl2alhODPSx5oU69KKyfMyJL0cntjDYVN1HFmlR+cnrOh0eNeyZ4RvDFa
ZwHmH5t31uewM6NPH7NXfqo8hqoKYeYSmwIDqiitnPJvOS+uNyMtiqY+GdBKco4K
HwC7KPaEow52K9mv5BqCjgfZnONnMM6xkMTyb6lcCjQX89QVoBmY5XNLYZqB9Z/y
Cx+ZZnHZyQfFhqReOrK8+cKEvHkYiEFF0TDibSkUsnLhQZVNPdh45xB97YxFJr/q
ajT8NNK9s3MBLtRSNitMOu8BssRSyuHZnLQn9Rre8GJIzzCAAKmnpLhHCP87xC2I
HYIvSFkRIVHaoyGL0d9iBge9OG24rqKLfCEXc9MzjPhdF5QJN1Cf5/coHyCJs3tW
C2G9YAf+YNg32LWUd0wG2J0/ejJ6g9MxcuqL0ZoZWFiqlIYXljY+i5fDygHjJMU3
6+WTXCB/sdjkeshIauzmwQrk5E4aHVr9qFiH+BRGtZnQecGWtKpNMXVhngsqllHS
ozW5FVPENjHJVNumAHCAXClMOQGzEgwNf2cTmG77GGJyftzZCDPcNUMlpHf5tepD
XWCO9Ny0bCNv7fl7Zs8NtKqQ3rchJMV91A3H7UZWmwSUVQ5G2WjmsE9HyPfzva7w
Gluu8kLQU3bOsdog5DLQglPQ08hfUJzanRgMUhscNUNGjcDg+umWUamMmN6OpLof
o6JmgaaHbCc58bN57EA9lqeUGK5V+AT3qAQ89xUHhUEbPt7yZz1QTDv94gQEXlLI
o9smJiV7Ig7f0XHw0Wrcva1eF9yrfgzzmAyqarazEMEXV3EzkVn4UPZwgRVCaHsB
euSZqeIwq71hYKjJJbT1lB2vYYznpR8fj8szu8pNZxiHX62EKTTcRjN/wmo90y+x
b1gKGMLmrT2J6BghdgWtWPBbIDCOFXKx2YrA5EPHwgGQSZ4IBDL7uya3ozoVFJmi
UwmiSjC0fiEv+RFOpSB4weXFRctTtEsnNc79vn7dASaJ49WEVm0/pWMBjhI8PZIw
XFBdyK7TLSUKazT97BTqphD73xlBe2GT4P+S7iPACbe2my+bsMA02GVKU4onsNMX
HE0hVmJB3bNEf02ZT4xLhcjClMBGzem3pXJjHghHthX2ZnOi7+03MbjYy/BLRLSL
hmOw7Vx5p8MfF2nMLJrrDIpIp4o273RC2RurLCyLF/moaNx3MbKz6HipNvSKjc/+
bPdUPiZ4FlLkIcOWfeg46t3b/HUjzHxM4usVg26M7jgZRyIwTKQg8MpEhdj5n9dQ
L57vJhkm8S2sI13HIWzDycCvyN0/Xz9Onyh/fFBD2IGkRoagV34Vo0KeNaMhpKiI
iIjeCgWQ8lgZD5T2Bh+JCLZhSF63jMVLzcQEZ64nKVLzjubnhoZXBz1wSd15s3Uo
3uRnTQXHVQYR/vMOf1L3wlUz6cF9hjtzzK/CQSnQ5MbqBNLEr4pAuOR1A5y7VcnE
7FZtno23VgRVo1F/+q1lk949+bSR+njDBi8S4hs9hv6N9uVGUf0AISWlw1uP2mMM
QTsect4papYaDzRTEvIdCeKXip+HCdjvg/ZZ6g6TVH4ODPMcahArO3cEvEnCaMLF
QSHTIyjTaYTMquRJ/PAM1RpPN4U4NtQR/I6UPudQV8DN3qzNooYTybE1bTpy85Oh
EJDVTcE9pZTTgdkFF5qNM//ue3zwUZdop2XMFixg7nhyhzFOq12dqgjBGMAV3xuO
u8h5zBY2ixFcWsDfo4PJgek/36ceCSxgWkdOX86fPsUMyRJzzBhYJCns/KftxO03
5Syq7PjN0DH+QHoftU3BgxfKSA8hDjZ49G4AX0/4Y30sy9UiwEz6gaYK7R762txJ
bOu+Y5gVJO8CnF24iUJgq2iIJTYpcylreW5QkugpEaIaSMBn9gBM7JVfRDLfwr2S
kz83cjUdYccScjuJf94VP3WWYuWIjgomYkkjdv29u+VNUG+d001JkdilRKSaSKLS
pa3pnrwIu/zvQr3jypIj6FtWcAFHACtQ2rXD24gnlG6SwdfbTqMkl54sMdCh7tem
8oItnoRDBCqvu2olweb0Q36ppTeLW2aWENJvE/IGqD9FqdKZxHaqryzeVnRgxGoz
MDGKGAOdiUHY7xp3z9+wxYkrvF5ujD6TrqJLriLPSXP7aR+aXVPomsyjE/FDGfq1
MsoDvAsGSFUN1jRcV57qhAdH5VLkPlSmI7b4gBaT3fGs0olgMy3cZlxE7Xg5WEKo
7mfjGXRTvVOOPHtl8oIjHGlUTPGqGGukPiucFmx49spiwsx2bNohc0O87cEASOIN
3IASdU2RBkDQbaBKRF2xW9xM7f0XPlFNq/b4wYm0BY5BSMj0PUsX4H9+JBhIc6AN
HRn20MSQL8q5ZOArRs1tzxotzE2FqQhX8+WNuJVKhsgzUBYL5Z6E6yK6ecjb+i4Q
MD0aQzUI6r1PQeXErpv0Yizm/9M9pxmEnU0hAXjGwJRAsFHa2uxNcVp0bgv64xHE
L6J3wCNOmZg7l/kWzI8ARazKXUfvA/PPY5YPYH92DJA9WRjh4PoqLaPD5V9SHkRs
sDBPkI1o+wPFVHfl/6Ur+eIz1EvamdXB64qNXmV4hUGHXP8PWpYZLoETYbXNr2GQ
QHRvqDf86IL5UgholF6UuGOLEzi/Lbem1pl5qEbBHZKE9EiECc9HbQaMLwuLBzk/
DwJlzIRlVL4Y9x6U7mBC5nPFKhYEosMV7caDiFfUS0YYRYizoTEuiXqwcpg1Pd5q
jYoaZNy/5T120I5FU2a4aN3QoX4HKhu32H8+J+CCxFF4mq1aUhZoKGjV8h0hBn/9
GL46ZMuF4bIPSDq9nNo1S334r/ENIoU9KiEt83fvAXr1yDQ6K6nXLbceBQ1bmSam
clGMvoTBhcpuYx5aMmmLXZKHwgNWlR/SQPy0/aQ26fbbuVD+uCF50mM4v8AcAfWQ
m4cSRtvTSpz0fSmM3g6iOHP7FERDa9/yg0cz78EB3E/4L0/57vylWoul9HnVV5+J
dSJbmLKMLGJqCteNdrQKHjYV+e8ndfAhrwODMqqRCDl3jbNkEQVXml5uSNRIi/7Q
f1g2suR7213O5IJpITy7u4jHwIA1za0e6npuy+7KyKt+2VUblx6AcVk/aGp9C3we
oKimeGTX7fdXiwRf8pQJxyC0Epk3B6rIEz3h4k42R+DxaR2cuBawmjUvtetoPcxy
rh7Y4yfL7DLVqux1zLyZREUTYHtYGKHPlbSA2YSTsA0aXi4xjMd2K7+qms1xbzae
BBRgGmsf6V8oSnSJ5lL21kxWe1Wp3BtWi9+9EboHqwQPHG2Y0D8+01EK02YVNXPk
S4GrXmrAONqjQM8douuQJY0XFSCjz+Lt+aYm5jOPhBl7JPmQC72AbMWzbRmnnb1s
6lwn+FvBS9M3uTTCgO2ZRRbZgv4ACFQYyMW9KFIgruXoJWTCnZHvQhpXOVm+QxSF
UIDeErVxawlPK+iNHQgCNUyV0+0rW2FE2Y0xZ6fS0OJ6z7e3RPutJQHQ+HL3RNCd
J+t2dX8Tcph/Elwy+I6UbgbfvQSCjIoEruwj7SMhPXX/nbEEyMdDTfiEksAi80el
9CVfTr3gEEGlVekMcIf18V9bVHtdGbXqZ7TaCeY3LA0twlbNEU14xuv1864t3r1A
N/0juJ5tXwCnMvDPEeZhKyJ8Ivi6MIn8H6RDa/wBW9k/MdMAlZl1KZIOV9RaWZWW
v/lJn0AdoQZmzh+42njOyF3oPSzxpswlrM4gUd/Qy2uhy61P1X7C6orjK+kDdVGi
QmxJ0kOL8jsWhCvl5W4yTTJ94ue8DX6MyaW4jexAV6uMAepsJcCCzd3qUuIMWY9y
B99AUdh5w09nGvdTs/NgsEGmZZGw41kst3XG3GlBcnNMgQdZdGAP30GNhCBnQtS0
m8eWNQld9yjpYIFv4UW4XIN1QKvMy9DuqzZeJuyFIH0Upx+qSSb5pPRjttBLKEtK
X8bHalmC3H4JMDMW/gIGcoiGxj2pxqqy4lSLgPWJ7unn5DYgAOUduDgCpSGGvA2h
cFBUgCcFb9HpQiISq283hl0usJe3y76Y9YsxpTrUESSBF61g4+CtR46LLg5UesJB
xwR72jJqdPmIe21ym9lAlftFJ//6QKf1oTFxeKl+6qJHga+de7dC+6WsNoV6f7LZ
1+ffZaI069p4aWy/00JFFHKB8bfvg6RzOLKzpMrix1HfFjW/nkedwVPQLdpQrNqk
aeJqs6rjpFWX8NheqBNG+pn/tPiOFG51TAhFm/5tmGWQ6+4iBeBIFKHVVIARqLuY
ZfwPgnQsWqnJEDsY4LIpM92SWRHkDQMd0ujjxpBQIcKjjIbz3AU/xGuIW7kBBykd
Rd90Txt7EtLX81xU2mS4fWp5w2VCDJ6uKu/5+gTvd+5rPFB2hEgCxw0LJIdhvCwx
lGR+sygGX6ZbFBmH1hgbZ+NOqT1QSCbPi63bAggKBXqRMzy1F/b6bpJfMhhwrwHc
c1PeMEZj+FSQVRUvmOG26oZdVY8eKkiCI9Z/sd5GQZRiVShhriCGyGOnK0R/x4uH
U5+u/xXkpv8NpqXvNZiivW9B2J6mLBUOGp79GtWVofikZoc3Wsa8Qzx/grmri5WZ
Y/iMWz+GydgxHey0FmYIZ4FI1JZDl39Rqo8JL7kmikm9O7jkvIG+P1Fb4q8KiLek
kuwqBwr0wTJt6O/TNhuecGFU43rsuNxyFkPY++wsQNx/7AxXgaEDSHHJDhu6c9GE
TPJhch93USty/1TV4rTVo/kTaGHPQ0/848HRfvoJWV2BWnwoQEua3H6DBjx7v+ty
3DsgW/wupY72c4D4VuSW3TMwqIMWfzaTbOrJYXkCU56EL6ImBhUIiUYjACaTW0uC
H/Hp/xWe7R0hJN6324iteZAfFEULSEwsgpP4CJWTDEDUsGTtSQr5Pq87zDZ+DUME
1bYLLVk5JAisbUkr6EzrU0gMpIeiedCyoNzO6vd9viHlbWJ1y4g1ATJk/3fkP9YW
WewGd92Le2beDMaClXnaSeaTV/0eMaikZoJO+kQv6rdfCQj7cQx4Ap9X4zH4JPHg
egKJtoBvbDAjilj8tkq5Z6Gf1LiFlozMAAsWyY6cQXRr/oxJpxLnnO2CQ1Cqn2wD
AOxQP/FJL7nUp0KuyPB5793tiMaG9g0s5//yRcoWpX4IFyDVvmmoJ2QJAvUoTBap
g51qHXyu/iYkSmIINAzYagK7nkpRCFU6rD4mnygUxbGvPW8SjgBVGNOEQTMporoj
LxpCjMgsFfDMkoLER+0XH22259J8jgfBihoHaEh8pnnCmMu3S6QwI0WN+08J6Hc9
KGZiohr4z6d1Z1jxVlG945LqG6ROoCVox8bRNAj0XVzGGGa7YGlK7VRZAtlAmljQ
GlXeAsytZakM9yjG4ksCFBKicTbLxLlEZzHb9ChiOytY2GJlIg+E9e+drOn7yX61
HvX2YwoS7w4KPA+dOffClO8HUzn0k4hADOCd9zPKjYs+tnqbrN+1otofu4a5Uwqn
YldKL1COxdKzfVt3MrPU0zt/aFg03lfCkWVPiWRkuavhkTNadyRyVBO2WJ5v3jU0
fyn9DLnIC9MLJQeIx2q9gySzlpHkeWB4FBwZEFO8dQIjO3xXB9kDmVVcqiZpooJb
teapf+YYoemwFPrKQP42a24rx685SdC26p3sVKu6WkTsWM9T115SKR6kKHOukF5J
2V/1MbTSbsgoWOjXwT2lg725tsqTxzM2dK++MaobiS6BXwBneR1P4KweK9UPEAs3
xNdDJaUl4tKrmdBjxpMCzksS/RAcEhwIL2XrvPL/fQdTBfuPNeYClr2kth7u88aK
EsJmfIicgc5oppH3ckFXx7X1DLBaVL7U+7/2ezy43iOiiKk0e3D+/EsCu/E88q3y
EACGwcq3n/wPa98PiRB0L1YNoSWe457a+YP622adN2vJXGjbYNYQVGDwROtdFoe+
sMl3mKmbfy+P5Ek6vrJJnbpNqULnSW8camw4GAF1KpT0ue0tn+wZrXXs4gbKc+8e
iCBEoqe2OSi4O7WqjzSR5XeRRCFECL5b4u+nWaSP5ejhe/bfgzQ4/aZMv+TYzl3f
S91BOwDvmJISe1Kafx0W4q0bD/MZhv0muWRJ9Q+FHHybG9VoDWOgxLrFcscMj39i
JOuAlb4V9jtsWRT6kfAorO9mCVDd8Q8KWlZpmiquu0Ws/pE02mCNPakgCnKypV4G
/mdQNXeWwfRNj/KUUqosg26vqh9KCjqoKJgehbztoe+v7HxIVDu8/FyjwiVkgHt/
o42XUk+fbzqNg1JY8OqiM8En0MWcIANzACAWgSJ0hxeD4eRtU2LXcPWrpZqFb72q
zp6CprN1Ei9MYIXd66Ic4o/t7elzeTlFmwLa9L5oT43TJ9P8IlM1kQwIxth0sM6s
pO3yyITzz+fU0SiSxPxr9b0JR7Jgk2N2bgDiNJ9gqULGfyVq+HY8Qv7x9Qsi3q+e
/ziKRVLZQWZVwGten9c3rpw89+Q3TT/PtsW8CIK9yjutCzG6Vg8VGaamq1iw4YLM
Ak10V7+fg0H8XDtGBZrMGQSFodpPUF5mt6NrE7re2QhN9SBRylMG+aSgeJPrV7Fj
E5NwaTo4SyxTmRSd1wCfSrj7lZW8PtdAu1XzZxA40HF9G46PjRd9Z+RZVppjqRaa
+ZUSpqQREKpg0+aoBjsVsUMFPi25WrFWbwRgSd+ioj5qfC9F4+tHfnxiImjWErXI
xYDsiANkijaReciRNod9TkG0fYWln5XYNQeolTvGSxT9nQmr7czcLed9kYNjlcjt
LBWWBijJDvdVsy/Br+QCTD3au2vgismQSK97qrtKVEXsVA7narmENxE13CHWEs2d
MmX2WWjMcmEPslbynMI4PfW+lYJc6La82VcJqVAyal24bxXYA4x5o2ax+wGfnP31
hsxgadbD7EoJREeYGkWoG72DOctHqq87lvSJqYwo2/+dy9ErvGr+GY7yHQYNbAAd
RgvChGlq3cTO++lK0u/2MQ1n+hCdXqAj5/eq29cJVXyyh3udFVU/ZUh970qEMNL2
8dn0bDWQHFu2WkiTdEa5REjIwqoPeJvK+ELLDO+q2GrYq20q23N7w2yH0z89+oqb
tnG/3+nWq+TPARKjFDYaGCoya4obQTU5MkYOSOX9C08bmBwSzZBjqBMiXWJvh0SN
AjjRrJhWjSNOTvLUJ4LAfvXfZ4czbZJ9RdqUAlX+GuhVpSKyWapJa/YWoHHBmuYN
Nd1KZU+lD38E44CJTy4QWACiR3dshnDASuNjlzYM36vkrDJ4MEosXx54osDwpCBg
q2C8BsrLZGvtFM2qQFGc8RwA20KJAiT4DaxELWTNfcZue9e9Yv3MiQEuNQ8PS1iL
qs81ZksWjUdLqa9/ScBPKqaALeXPJijRUrIEcyrrVvpM490L0kHd394pU73phV5y
DOKCnX+apLS7V8amHVDOmfZTid4EDiYHwuTs072S74A/rE4Ctf1YLn66dN/EJncB
N78wI2xMzqTBxWQtWm5vZ1ujUxhhSYpsMgVG73fG97zd0g5usKpZlqgt9QfQnclA
ecLRD3izVkVkoiqppmQ6df36x3koVOjk1cEKeqWJhm2MXKbUFdHqSQ6sfJGDXKEM
ucbxC8X9cQfmorOw9LRPIHH7HluOPrpKyhe45M3c5fNboy17TQT09ydrmVjmR1Uq
IGQKD+iOz69KXsGgAgGAOquyrRNV/IMB7ngofRUisq//zKX14QI/XpDibBOVxpcz
hTWnPs2wk35mhDB2oQjiTIvBiEtggVtx/jbV+6QsBYNErPEjU8G8f631Flqydxqk
CeCJS9p/tkYaxAol0GVdNoj+4u5VNOAZPHdHPmakMfzA3Ca805qLd08bf7fZHfRm
6KvGd+rcm4dnvOOzGioTks6JZZ+nvC+rPgAWadzkO0bjULvlrq7KrBHcPb3EmwK9
RbjDOqMFxCsaHxvdEtK+UPOivoD2PCvrzq8ZSpjo59rnLBw57aelXWlEXP763n6i
lHYOwkzwHyFZC4Mcl+lljBGIEPfh7ZdSU3ijLsToO8sD7SQG74VzVmz8wK8aIcPz
3j1Oj4xBEJvGtBhM6lWG0eg4JFcqTshh8n/NF+Y2VhBGSKJZ34X7Znt8RqqjKIjR
dgMpWafddnp3SM9Xr3x6bJA154+1KrUMpWTGdd2E9NJxKGbmAmg/91ZZAYQXF72f
KQfX0zQcBkdpFFQbZO6cKNtlkcrC6IR3SX7rX5o5APe0/U5KhoG0XtJ06iQ6VX/e
+zhwhmZCxJK5rSqMJdMwFW4bliC0mVYlx2PtqGvsy5PrUwS7/FC0s0obbOp4QHcw
dvVgKxMWkRZMCkHjY8PE0T1bBidoJ2i5Dt4twaF96cFDQ+Va0oaacDxzTU2xzXiL
sFXUyXCYsLc1I3DKJNp+vD4PJ8ex5bi2nj0ohGCmKa7rNS83O2NS3HaMunum+cHr
UPyIHgvC7jZ7619XKKmD8/De5J/Y2ceNfJOuaWHJNQYp7sVkYpca2XL6DsCwpxLR
m9hweqGlWGwk3wvWIOlmh8tZ/mksai7DDltdZDY1/41GDj7G0ZYNL2koYuDA4kOS
G6HOeHcNlPGMIh8JzOZJpofOPisAnlw6uOluZERXSXM8eCxY6mtgMxv3oK3thiij
79l0BKMmn2Qb7VZsMRSXMWrovWaW5ooJGizPTcDt1mdWxJVx+u33fv4x84epdDop
mFbaOj/zinkd93vIwQLppzhZ5HEdx8lUqNgrXdjBcS5KVVJ/X8D7/NfbcC5DTKPO
sEBKS6RhS4rT/eV1ccxNj19qOazrzhbeJS/xemnKvUmhNqTVZcqDGUwpPCn82qXl
YgFsWtWIkdNjG3yO/mVpYi1IkgbaK7vHMzWhoDQmrcOq/8Nvl9uvjCsRFCkk5C9h
9Gw2O3NPXHC3rL/AauBVxPQT/r8QOspwI+IlZzJs7anFUt9N0Gap0erRMZNSKJM3
E2oRLLEvjtvfFBSe9wNuZVwgiHDJ1kRmqS/DL9PfE+SZXdM5Ut8huhKSmzOtC9B3
cPcRvjM1QGOPu47TCMO1Q35VHhqF0G5Vepr7B4KzHx+dgAbVx0ANL5bGRHZdCBCn
rea7QD1U9LQfrcuW/zkehTZIJhodLyKqxw51yVdy/4QlvyZR6oWWg5XzKcK1IvLB
UbnxSwcuRuKu4IpFwYVBc0mdp8ggoNpL+8qF9Ta6ByePZR0FDLtWuuf8DNKJFmTK
D5B2YShuGYmlvfq4q47dHyMEMLN5CC1ZbEYZYD04ToU+naeuT30agCO+8cpK9nJF
0G1EdlNCULVZRz2d1Q/kyd1iKWT0wgw1SYoEkw4sc3Q6NLVQgxRarSS+utah2zqn
KOaUcRtqazX7mVIOe0MKg7TKo405MjYWYi5ISZ5jBTUCQMUzQsjtr800iw21V1B1
p7ClzqLL4eMUqdDO/VNLFqxGkuxYWOyyITzno1CcJCPFU/pnWp0RviVe8NRvZYmB
k1lpXD+OqG28zDwihcrk3//sDgac829FIaDBblZW+k97t1BVZb6SvWleu4S/Sbg5
OiuMBgRCZ/P6jt89I9SerYhFxryvpl01E69eiqYacBzJ6Ye7Uj3z6i6oBi6A1BmA
UpGbMLWfQcDBH6eOqH8pLvwCPl03MltbicdYVAw8RiK6DFM2E0SfckO7fcVbN+tn
zx+Rt152xAYxlKiFoamjqP0Puoqx+eoGPEwTiXIHlFqdLuASCnWiNIQd7VmEncBk
rxRGPxX1QE1lHgScZoAjQs95JJW4YO/BVtJ2bDcmcwccC7TX1DuvC2pL7Wlm68dE
zGhzvudzLxiPY1471aTN6kWWaTnCFHhjLS6twJYnMHTLf0hgW0hAwuMfOe96sdB2
Q9bK+oqOEhalz+xmlFFYESddpqBgm0QN/CzucZqDa4YOFrtRbNeCLkFcfYriN6CJ
zOLqvra7cUaolKo6UHRtO3/9toreAybAW8i5No1nmutDFVtcaMWqC0SeFeXe3wqz
EIwnGkFq0jVmov+zEULZ7g0r20rl0100QB5ffg7OJAtBzZv/+R/WOLTTqmnmlDEA
M5ewTxsRSzMkFEuriv9fB5e0xbi0JsgqIhxc/eeDcNM8Oaueq6lokmHiIYvm+ukL
n1d6pPNvURAmjUz4hnFTuL9IKrVpPcFa7vIAtPQacYZsTkaIUwsOteIp0+M/A6WV
4svaDQ/MXIb5RZPhw9iz50GBnZwa3ani1wnGzuAQRGbwKUpZI6s1FMwXck+ib3/h
w8cVqNTrDAFSxJXy93Du2PrUgsa31F5cmCDt1I8nEJwAJetCI/aj7XOWLnJ34M8z
69gOChIQ7Y1N/wiRrFOgsnXf+V/CMMrhJWeEqQ/FWJNcjWDarXL2YTPm/9EBLLUt
PiF+pGqHrzbVHoWeQJAyamK02iGC36U1CEvDbHBTeFj2msa5RNuHyhjhvreoyWoA
0uECgNHMUZ8hqZM5b5EFSxO0MDscK/mNyBgCjKAsZOnBBLv8+YUzp4t5rUb4uWZ0
t0XcJaa4eX0Km27X/Ut/L1SQx+mCRMaNCfU28vhXK8hPEqE8WWjZuRCV9dgsQcC7
OqXXol5M/nQsFsarPWDUVHzp5m1b/b58VBnjXhboL1QJ/i9XU/1rlJCK0cbZXcKT
Y+q9FU26sX9wWUpjb/CnSg/J/t5kXroym+TazoSP+QUcz51zCs5UZUfSmHcbOvfR
bnOaPTfdazfG31g3NG2W8rmNUSxFYUh6nb13PT54XSnNyA9bQcML5WyhJFbTHdo0
sBbl2fBJX1PUKJp+XGAhuVLAqWwPx8gzFHG22xnumn76QlIkH5tApYyOKgLnfm6C
1jjdLOP6K6ugLSecrE0S1Au2urJCZq+YLHaVKf5CsDqG4L+xwUhEWUaT0V/es/DC
EXp9zfXqtgZ9LDwQ5Rxa2P+S5gKnHwVOssocGo7gFvTJbbVT0Bd203yjkI2oxek0
PGBTneUkyOHkL1VxPEL/7d5Ipk63QZ1b0SESxpNfiBkgUDIm6N1QuN4M5iIALy9r
c6xvXp2rB3I8zi+XKaea7BI2va6vwpbojC6RSqXosRoMXBa6vmffy6t86MRsrl6q
Ok2wDJYStnpiGO20yqcN9HRwU6nbewtucl+N7s75FFev3742lN78UZ0GVNp09uFb
cmiZf2zIIF8Ti5Vqb8YfJuiF1TbBYH+BZBeygo88ThXNgDXyDXQ6e4wL0rSZzeLm
Bmy2+7NcOneazz7Oqu5IY4HUSk0j9ffNlelHIuFZ4h5gwLHQCD7qwC9Jrs+BMFG4
8EzMqjfG5Xtp2KhMJ97C0E4VCDI+J04F6LuL5liL02xuaIFVhHUXcLCvvcPMHYn0
n/4NwLpF5fo4MNuIkn2t5ZXUgYfij28lJ4cTvsCFekxEGusKumKFy0V/9FNnc8vF
cXdUl3Atq/4FPfgHqx44WvXuC34TeD7CO0SkbCxAxonJjflypo0C23nuf619yS+C
0rjX1UsmbyP821ms1M1Fvpvx0LftfjzsuhZH3mkYLvC3+gSZDArjCEWbBEErO6fT
lNPFsjlfXeGrwr2H7rO4y4IQG25dCmWuRTUcXF0XIR3Y0qmh/G6583H+JxGhtuz7
CbLeNnpHI1g0DhvcM2tX0sqJIBXHA/YjLe1StXoX7kFaogHzntBN8fLWcEcV0d7h
Saa6bLTciAyreeCzIPhjxcAGOqb0TXoGZbTT4RL7Tc33zYatnjJ5lB3PJGIow4TG
AptM4kmn6hUuQzrCDoXBFR3vro/KXMLWiHW4odwshWrJFC8kwNbDdDnACwQTkYr3
eEDadeJAmavjYJAVFEyM5vjZMeh1ENMxVCLjKb+tBGOXPAtOIQlOUrjum+9SvnHt
El/a84uDDg9/9GNrmmTfAsCyyrxUj8WoxYszU4Y2M03Doqfl+J70DnwBYpLsVuGy
VAMuk2HwzTmSwQGCf+wzWZzLI5XuPCitg6I1oNV4+HfSdT7h1OjW3QMsJ4v7Gioz
r5BwBOGfn0gm0SLb1YXkjKtoe9iqF6fya7XclKgID8OSyiAnw3WBpdBRYYKTcBtk
sLGXnSEBbVQyUwmftpeZ/8VJLsj3Aj5MIO5dMQdjvvyt54dGavWhCyOQNwsDwjEW
GomziZYW382Aq/cOKjHFmACuCVjfvRy4XlLmMUi8CLxeQac0jg3bl5ngUqn1Ymol
HrZOWDfCv0C3pMfyBveXezxXv0L15J11NnIQfrqOBaMGoOBhXY3BZn6e/opPjcLZ
YmNDPdHaunmUx0z//4+9NegtfPgQtZkOltJqUsRlcqlRqEAZowF8nyA+zpLLg4dt
miqzI1erXDZfD/rEQyIEvwpWS51i4jsQQx9tUOw/lLVtUaBJoct8d11pJMyOz+2H
OPeUF0rDs2YXtVFen/s7FEa3Fj24b2I93QS95WPeFb2EDg/kfj9YkGglIIx3a860
CAzTSOAwP4VggD9h8qeS4Vrq8RrS5Ep7MQ77terLY/2Kz45LujtqiD115O2XAwcq
0deLrLDguEqX+heLApCM6Ty3tOVj+m1i7n8ezmeYADce2f7nxv5SAbyIGYbqQXCC
iAI2tMMUX9VXNQ+7Ds+m33AQJZJGdRB7Lb0TWwpOdC3ereGthcTj6DJn2jpBmPK8
rXFwhaOuDRFhLEsQTqtdLq4FeanqSwZdnzTIGMYK3YyGlkl0rBeh4rj7o+46DOae
ZocmvlRr0rqthqgLaoBdVHWu0+P3zDTmAw3NS9XJHfU+hXoDWiF3TNZ5LB76fRbp
Aaimd6bJO4vP4fCCKBEfcS5YnhiZpsdNZxZtU/PEq5/GabM2ySQHQVnX2FF+RSkH
7vUw/rVvSguyDwm5gMpNqg+SrN+mG0FY75pFaXHVrY+LPeEzFnlnQUVzOYhAL+hP
ckxSOp69cxK3GAMthyfT9lWwDPhCsIOQSklcqj5CIcsP5vUIeRT//9yZHzitMBLM
DdRxA2gUELiO039SSvVz9TT3ojZhdBlH6BNXr0Gx2J5POMpcPVSDj3Hsk23pmE1h
LGjIC1CVW8SBrRUH7NslN9/YSgyWogpwVUl3Ylg6CE/pJYHdjcakqysN1gxxP7RA
R7UfDuEZioDC2zRT38+4ul3fwW1VKFAKjou0JyhaoXw31Jgp0pqQyMjKfRjG+MIb
6O6uvUX66KQpmihs/MZSYkIgFy2H6axbfjk0s3TC5/NskZ+AZi+2b6gCMZmLX68t
Xz9KfLQ0YJNVZKkhPQrqX6xMWbKgV1AhaE+zPF124JVK3f6/okEl0l6DFS0duEs2
Xc7TzlBg3pt6yAxg6EVWVJE5RYNtHzzgL0gbfgYYpMEU4Qe0qXfoqRcKfMpxiGfF
bkxd3rzZ95KjQiAIlBOw9NVr5y4HK1b1k0sMerzHd+E3IbvhOukASGw0b+f43ID1
TUnpcwWVeKcbj/JG4V2yl2XJyNLouSR7GnDX5iLREHI5UGDBrMhDzly0F5qmq3oB
we+hLg8V2Em38xz7lreM9GfM/de3OyFxSdmPlMRIO5MZrBVL2N6/hxM1bDw+AI53
uBt+J9efWGJO0JFVKK1Sh0rpaXhibqPhuPCCMMzW8JpLaskdxdFUn1FK7iL9igRW
R4pklL4iNkTk2or9JOsie840Qo4xIxSpFcb2CVoISfzjUKzI6rlqhsUWyh2FPqZf
nFj0LRpQtwaqyqqUeT9MfymAfk2ng6Vvi0lk2NUWPGGfig2zzJ1RDA9IPgafClLX
k0aW78s0JMGS8ylGpYUQTu5i7aT5na4bV/yxzZeDJKbnKiQ6X3zm228ho9F7DoGZ
iEDmQ7RHBtKualX8HZyXIaY6FIl4J05RSocf/fkSiHvy1NE6J1RsMXgpsjmYtYou
Dj73gqc59+NSL8ddLXvk4+o09qeTIW2L3VZc6oaZJamwxBPx7r9TN0kkA9beWWp7
ahqdNVeLng9wH4ta4vJ6jLt5F5oXnYf0VzD2Tavg4QIOPTYOF93vUMOBPqmQp/WK
DlHt5v1dBdVVFQnH0TuDuxSsNsL4rzytH0acsJ1K3rlWb8vJlqWSqNTmgJFQ/36Z
BDsinW6Fu41zCqBeNQRiP7ZTEPUUP6nhZPEFN2bgb6K6X+Y1JVjxhHYs3WB7lLGo
SHsf7/mI1TL/ARakY60kO7W12KN0Dnj3PCC9s/QpxJ6NmFRdzBZZBfgCMHvIzEuf
Ax6ovnAaarM+0eTg3/ofwvApYUQDWWhVpYD9l64wM6YRzoqjLq3pRJXLFuC1aT9B
mR/WjAwuWVOFkxwG3NcHR79vV64MmvNXbwF+X3FExH94I/RrqQQQ82yJaPzxs7S4
WKUjaFaumuN0bhrW1uDEE3zlP+HX29wBEBBA5wi4dKM1e5PgpaZnlk/p8Q+SMvqq
k34sf7nDZLAm0PYIDLrDMDBUaiALsEkm7zDXjPFw9V75AC/cObRS9RdBQbUbypAm
+7yFtMzO56VKUpGy3hRNRHXUM+xzD6XohY1VP+tf4GvVfB799tZgsQqyXWvwIMOd
t/z8NkQSHqOjwsykBDRNxaYuDquE3JcRJRYhHVa0qAq62coSIkCpzayaZ7q+45KD
jyPg/zKU6+ko/tRhe4uoKyO50Awi/DX86InVCCF1n1jKEujNVEn/X3gHCv3Suxvx
xYD9KgwuRAicM5szc0qVswe+JvWkgQLeh8PtYYbCPkCblkboDDwjguca7+nrlRW5
BBgLEFaxA6x4dHLcElwU3XMzyQV3yNe5+EJFL6E2BYZxqX5fNjjJ5hZR3kosFp+V
fFUJnDd/N00mqdNNKFulfNkmB+fr9RqwMRxbFP0ilRhAR68SserKQYOV+oCvHW7Y
q266K48uKuJTJgeZtjrQKFDO0N/jqIRWW6B4QzASE8sI3mxgpQqCoArbY7S2UD4t
3+w6lKlwQA7LPQMnNJ/7sD6/UGvQ8CYlfAXxSoN+TkW06Jrr1rV92mT/M1pJOLnR
CJf/qNO717s6/Z217nQ+0YI+MH2rzXp5XG56u/TAkXGrdmxwIe/5QJV67jwDucua
duNsWk7yMczmRsyu4ivSxBEjWWTNg+zGci3cGgm5vS6fxNGcGQIf4kgRIIBuACoF
Y0bgmIrceSitayQXYCahYbVX3CMH9V+7op+V+3Ti5hjH/sDF2Vrvha9jWuZwqVAO
5NpgIiRDqGJdlfVn/9l1ucYL+tvSYZCru406qyG38hUBPfDdsdHTM8CV5HaOQ436
SaGzOnklojAJgTEeX+Td+yVAQTJZaEGX2tpGBv4HAxjG+B308uwVSEAXjypUIs4r
Be5IUbcbNUbXValv2pJe8QDIxlupvUHXd0mVKxNn5+uNOr511igeX6uDUHN6Y2Wf
Uoig8U6Aq2nKvcSAb1YlZW2dfCYMW8DCheVPbxH9cNP2mvMUs6j92om7TdcdVthC
jY5nrtO5aOykNirJx4LAygveCh98eH/OmA4fXbMRG50qrFlofvXdWQ6XKRtYmemu
c49XkQ2g7XyuvAPFuFAEK2zYoR2PFdhOxLdBSvo87F/rdGmu/atRk60QZFOiqGF2
2rhbyMsKR5y5yvdyVVZqzCMmvT5Jo4JJI/OWNJj0HAf4DRaZ1UoOLTW+bMjpT9Rk
TEsL9oN+f+rzblsaI6Yto6ePyq/v/5M0jzkH65vMXHeJvhzCnStRsoeIKrTBVjbU
V5lnVZLFKFDk+TMUCYhli5dnELP7zNJD5I6e9Norcf8knlD0LG7K+NSlI2XEc1Me
2vOVXYhpvp1EFv/Ibe/e8vlMq+s5EfkiJhDBPgERoBFUSU9AJTor3i94X+8oQ9SH
mC82mfn3sejh5yG9oevMekOC/vqubF86CdG+He6BQUgHoWhrvJNR8J4Dtybve7Ca
d6RPVBZPQ5ASFVOtJejJD0DOrOYHEBUnkVNF9pXChzJfuqeR0wV0rdoIkM3TvUGr
PVBIkxrp2Z9UKui44CxXXd/aQSDmgIaTL5sE0Tdo9p4+fgzTFIWeX8M7f1itx3xQ
bKgI/pf5TgooyZ+tJUQVkcrUUnzBB4gSfSRjcbFmwnJhWhGYke0c/2An2iwphvgm
XTH4ucNt6YjJZ0rT7L1Z0MlUBXtV8SzmmqlV/fbsDEdaMC/DB/lDSyH9FEvYwI6s
pCs5vEc/DvXhVAddliEpk7/il0Mouw0PpqldFR9bBtZdw49wecdwsHi2L3xLljO3
W0ZD7VFDnJmUqlMDANfJvb5oZCcUZgto6hUirdvxCUm1atF16+DSEJpQ3lHhKxCa
TMNLOxAcxwwXRL4zbygYty4I0Va4NgELvYRggWFK/pKIj1gNnzBwfHP0FrwwnoWN
+gk0Ci/aAYNJEDB70QHyrUB2HTDhOnUG3qrxWkRB1RggfY8UmxHUMW3YirvmKeXm
etkFsP2x+WHywXv5bmZSMDgeTX4NMHurqUF2NuHXB9+HlLtf1uBvHHNjxDbgPcZg
7TlI0LMzhY8hJ8RWK5fHkfvktcQQ+gKI1Cq+XQRE59NjIWmfcZSStiTzFdPyQMMB
ETrIhVzRwTualKSYQvllrKceZGjdTcXK1Zy65ZgxXNXv0qptPJsveiHhhXmNHFsF
mtW48xkEqXvHVdjKVILLZrI7XdOUVDzIA+1jUhRbOzm2WGLP/kk4QoxgHFrfiguF
KAUSFQR9H8cnuzVN2FuMRDpowg2nZVeXMCev+uQ6vl+0VWPqxY+4ubknff7jRcpT
cbMwetUgb41hDX9Nf1prI0CL5kHGJOyyTxdeYzVGDTDVWLM6JIsutXjCe424oWie
XI5NltitFrMoD7oQJRS/3aB+xR+0zMbpj8TvlfNXCP5H37quVFOA8QFJ/uV8ch+Q
CHjWVjRRBH+cWZ9QrxSl12VQg29PQkQ2OS+H96j61gsXClVYV5dWQNocIpHPaW3V
erS84SGuI5VjUKKeNOf2YLXA478gIMACH0homKotzSP5yRMhEtujl9MduuST9+hK
05YTZWaAFtcEa+3XsAchgo/F9trufp6e/e91a1oIOeoFl4qXA60BO+RRLcoSV+HD
z1/m8bczKfv+Y8uHnyDx+i2ejxhWlzp3UF/7nVdDFixibthRDk+J/93vgFV6Yn/y
ie+tO1JIhMo2ilaFcFvimSh9GeuijZp4T0uNOGp6rld7hqvoINIrChX0axj7cl0g
EzpufMzztFjABexf9R5rGKm8MkYlnFZ4IlA1iqtyC3DhcxlRy8vWfe/Rl7Rr4G+8
Ss2VzPlVnhO0QRXYspb0cXPILyzwn0ICyB8GxQFiseQKWrWto7bAXmV7+UnJ0HWW
pQm8xnNn57rs/jCW20exvv2KH4c99POdiesV40y5VLZC9YGUpLJzOZH4WLF4R2KP
1aB+xn5kd5gBzqvmk4TImJqDVjIqF1pOQpT2VNn9DkcQWyUQY2E3jYTrtSRYHq7/
X8tTSMCw7NmXDIcLDwZgXMFTYO4kjSptFcEg+6fnE1jqjKdB7IBqXz49e52IaW3H
eqaKtGx1JGTXokQgCITwos16KBk/pj+hIILeJ/FS8sV1q0wkUkmVi6W3e7u9ItXx
N3X7CV6FnAtk6JpbNog3pOT0HIEpYs10AHjTdQ7Pcj/12ELTAfcZToGgzHS6MHp6
7Q4gHAncKxqDAJeur1kdijZrXqYL16jqfeLdqtXMjTSbR9QxDJ6RKV7UsqBzaVzd
3wgxROsqklHA/OYMhJyCP7XYTYXfRree+IRaMtcXyDgvzFsq7qqdQ1sBWfR7LY7z
ocXV30q+vbWx7aChEIfLsD/Jb0THU3sUMPCtamS3yY+KXGX9kkb4Ciz9HgEJXfEI
F06gDFhEOT6K7tOvrvyszHpdeBL42L4IRICWOiMutceCTO8wlcc36XgwzDfh0Q7T
3/ot0XMw/xu17VQ7J+Ps64z4/n4A6T2MjX54U5Errw28AAFP0s3S8Ojkx0fpRLev
fpOPJF9jXXXS/RXCn3Nt+m830HsZdmOADHeQ+O6Bh5PhMWy7GIdgujLhsJpOF8sw
x4XF67NeRpBTVELbUCelWU86BId06t+36pZiKprZyZZAPCOpULRZP6lRBtaPwGbF
sXVjOGspwXfpXdhzo43wPEslgf0DRNmUvHsToVL5p1aJCQF6buvjGcjGDegztBNM
RCtNzfcuztS+P7QTIp5ydCtQ5zZT/i+/4/1sN3hRTzgOkemFLE8np92R2D7Iv58A
u84KawfnVcPp/FQTIDbX6V/SZjxaKrAF4taeu/a/k4WPWApcp467FthFtxVVyMXC
9mX0EtFRo4LRHt5KelC/9naR5Xr/qfwk6a2L+Qk2xLwijx0KgPuJjk4n6CVZ0Num
xT3+WfciXg4sc4Eq/Q2skx5boZYQ6hJRiCEax2jcx0mMJ9E5+RoEqTC222l/3UM5
unIoJp34l7iNxCrzJE412KZ3pKI+A1W1AkvY/ztZH4fBVDIByPL6EoAtLttQ6Um2
HgXK9OTVYPSLFn8zAWHN62lC7u/tnhD+S1P9pjwanCWW7Q3m7hTLsoZwBubpIeaJ
vqXEKkjT/uzvcXf7eHw98fQDOoAB8+nKhHwKDbqkDu01LHau9n2ZfjCdhjLCx6Vm
uiExYy2ruB3c+yoHXoQeHNiAljOdGjEjLV6AszcoszKhmUPR3xWLIaVotzWODEqd
2ljQ6TY7gJ2baRJVEIfL1yCL6f3iI2YqXSoNzkZwP2WeB0h1Pu7Swfvr2ZcvfiB1
MAs032gB/lI/j8CBmfYAzforFIlM3FN/t9wSsekOVxycWgcwqIPGwf/rpA0NZpm9
AebObWd7s4DqaLLtLa5dVt8PaRYg6bF3GbIYCndfQfLCiL2gHkRXQiDdNIjQOEBz
O4+kWJowfgYkEUVpFN2qs8QkKtJwzT7zz8nhx/AK6680Qk4hteFD2Xs0M77otS9w
zOWylNlQSToI/37YzN0vhFOF4+6FZj0f1j0O3puIPS8e7EtP1MpXsbiwDJU3L+HZ
r1kzXrk5thL0QA6wqHHG4r6bhfG2WGbCe0vkUbeo2h4QCGaMfWc9zxu9Zj04wBhq
5q5Nr6ywyfmF4cHzAOELSIwPqhRFQ83OAfAKuOQcOMmBkBHMcK/i/H4wUeOX95pG
HYiIsdCfnc1reQrng1G0QgF1VbPQsnLPEIA6XTLyNjfw9wqu2Tn8G205YFiZHVgF
/foxjNx6TacIUfhINyii4bRJxTbmekqlSYR3kTrHGp3w3HduPrK1WlGnU04QgKHb
d+pbL6nkif4QSizBB8+UV2ZbfvAmZgYQzKFUKaVlWDPyeWo55IW5MHGCFYbwynko
X6LbTu9er/cv9WnUgqNU7GE2AZ0gR0gctD0ogA+0a3Hm5piVJ5kGBwcR81yaoGcH
mio8Ld/syxegN+qUsqwjJQ+GxWUcwuVOajOseIQz9m7Wq9Je7HRYQcdJpwwGOXF1
2K9n0dNTgSOz+Ho3nxOW8blUnuEXqxXg2w3FeUcXJ+8zWxPtKSA0kD2zasmmgK2j
VwVhh5Tsw5CwrYkVhltlG+WIq6JuaABM96v9Z7Q6R+b/Jd/9qFPluladq/6vMOmX
Ak6z3zGFWbxFnhKwJDjw3ADzcju2EDBudo6kfxzDcurE/QQ/lPxCh0d4I1iwGGHN
POv2KS0l5Xwr9GcN9+KDAxzpFfLANEj2BwaZ/ax4v0hRbRx5AM+uPCy2onyP8xam
NHKsQESMGN1TZq/YTH5FE+3f0txAk1XIaANgm9cyna6+0/31C+vifEpzhQhEZrCn
BsoAyut4V6h8woTiLlLPmX5G0lSjWPqPUCeVlfOiHxlISRAqIsVAhQRSU940MuQx
/2M0NaXScOmdRoYrcjGBwrO/yU0L6q7bpJSYx+xfcXty+JDQv+cQMmuVji46bDuQ
++gtl6J8Dfn0ytr0qnB6i9G6+khk+vK4aDZOBF4cfwIFZknwuJqerjOkGl1kSP1u
sgfHjR/nUdlvjR4GGti91RGb7gvKB6XNdajfczmnIw3mm7INO7JMTcjCOZC8X1jN
SVZv40cQjbO1GXcCr2fl7JuDxgUN3n9yk15CcaHty7jeRJ6EBBGHXfDVJwxEU6co
c9i3RozjDUp9fLpIUrgyrTSsignvbKChtKH0YhDW+VsN9xoSS1A89bK3srNbHG/B
UVmMDDQOQGRDA0IplLDs6ck9LjFrVHui8WaVakdhPA1THkVjzJJD2MVuW7r4MuDk
UxtukN9vua7e5bkd4bt60vngoW7KvYeHVH+YwZCKUTl0BXWWufEoiJM/tZ3OpKo7
wqF07v+srUh6DzTY3HcU5X6MrZ8oXkTP2i8OFgNzkDufC36T/246FhJMr5PO3/fk
5aN9DGey8cSR0uvq3RCgfNUmMOONuAvwcyx3++Djc1yi2B6A3Oozp4oOfPKvKgfo
IKr9dsim+fl6yRr8PbnFJtBefA9gS7fLPDgCFE/tlQtu5BufXtALFe/TvvsbQ8/R
RQF9yKc+CU9BDQeCORnWkE/jfW+GiDeA8g3Sgt4/ud2WxHLdk33ND2n+EUPYTG7V
+u6104SKyKBwsSguRsTcmqH09MUrIGNIdPxcJ13+LAt5mOg6m2QxA211wEIhBHi7
uEHy2reH7dBeH1TveVp3B/vhXcF29vNvkuUBUp58d0snPiI883/0OfhlbAYoQZHK
Z4BSax37ncMQhsPQ7W/RogiYrD4voi6zaiBJgw1oYcRp/Hru7cQQ/TuRJ864AihB
GxsojPLfRUNRlNU9EX7AUVOUzHt5SIvdRo5IYfx5/Zspw9z2HcNnquN9+cS5m33L
z1Y2Q9ibzQfT0BHiQFSFBTk+PNLjIY6+6i45yfE182VnYkpJopmAIN/eJsF/K5qt
7ERi0SVoXR2qXGspQTAHgZaPXHikJzI/9msc7mlx4todMq0Jr78tmPFmnyhug4Tk
SZHs6Umdt/c4eBkXKdIOBX+ZmcorJcJGQK8nSk5i3gt/gXKzfdzxYLwRAYO1lfQY
bSFibknxx+/3pn5BO3ORayWwWmjKsmYvQruk9tZ86Ytd2RRnIYYFr6N1SAzisNnO
RTDuJ9YM+D1/4ZhVhJinV0gJl0ouJPmwo8Z0L8j/SmQtYQM7z/xYrDX/7lhc3oMh
G1+D/XQqKgz8Pt2xeHWLkRBVn0b3CnWrJ2NCknuGLTH4FtPu0BIyrQsSfyjuAngD
NI1YDkxU4CXfpB3dYA96fyDa7TAgonWa0+5A4MXdyOi4cmLzPz4HuFod2Jwx4317
8WoHvfjwPjgk+V8vK6v72o70RvcZuGVLjrlv6KRo9mvwIHBcTMhxjWh5ElQVJg2i
gPDIHB5wlBNna8cC6Nj0uDGQDLbMd8xEGnRaiUTqgxaObAuXJkY0sJrk3u46Rl+K
5ds4k5dGO3tpHdqvJRjklR4SZjupBCRkD23RvfuyPRUUal8PJidtFdnkNzQzT5Yi
DKDMjs/gdHXoVW64VI1p3Y5w1MbmDF0jTxZ9tNsbrd0rjPackcvAJ3ImCeKD3YOh
cKB2BXOsnctNuqZhyj3xDGgbz2BlQbuQhNhzu5ZFdx/X+Y0xR04Hg766Xv/8+59d
GR4hAVUoE1c5wmRqRkzHlAwmjiHcOrpFePQIrdpuUjIIROk4JuFZFN3KTFL+0+RE
4J6rrynPnr1GU/LCSJHGmiCJcvTM9YoCtVR+I6QnQCF8M/pdfQFo4ZPQM9zgGwnD
EKx0Qv6SreLf0OMnlQSK5rdOocCUavwq2IttEJA9sUaqGyhk5mdTsn+j++Mcgjdq
fD47s1RtyBV1YBDeD8bQMTrLLyip2xQsbrkLRfLG3HkgmduXY8Y2yEisCJmQqfYJ
337dZSsFlB6clWaNKR2i2wnYfSIiPtYku0JdRmSerDAuKrCrE6DUaEQv8HV7IwdS
A/3IrjKoSed6vcpyUxT1vQXUMwmshFbReIlPO8KDSwyzZSDrzncvim8KfVIoHDiK
lrZN1HEJ1Ds35MU4giuSyBs0HsFeJjlmub56miI0T+j0pecwOr9qsMwu9pvmrSMO
kMU9JgB9IX7hagqoul2LvRhBTA102pRKxwFDOJwZIE6589ZaESlziZ5b4Kztqyy9
S5VSTU8FCnqK3GkWH9vYW8etDegyzcFBXjgVsp82x80OdAO6pvtAE8Et9Eh6RS7B
+VUQQ/jN6Ig8BK/htk0YmSubJ5dkQLB2X9rTziyFJj4+0ChJXF5tQvq/Au1A+GJ5
Y+rTNvYtBhWsd0vzOIZmZ+C95hMLjf53lyfIfud6Bom5n9MPasaai02O57ia5rbK
umbfLmj9FzMvcrmrgZrTW95pkNBHBOWJvZqZGG/OxKveXl5iq3ACVEeAwKneZzhm
rTx2eD4UOjLc4m9Ke5EAXcqk8Un09Kt2jGzRGHnohVVSpGEjubSxEJO6dgqN71uH
A2bJ0FwhNP+r0Cx0BSS1uszpTJLn90nD0XHr6QtDjJGhVAygxCdxlrUEnukq/aGr
GVyR51Fh4jsS9kQ7zkTR0Beg/zjDcBVk/QNiBc7CAEOgHMZ08qzn7PBXcBlCQd/i
EYL73CQj926q4Arl6GZTSRVLLE2ScjDWSG7950kMuS9b/9HziNu2XGzO6mM3IIAQ
09r+Sza0YcqyAv4/FG9iipKwKTeob9fXAikzmPdxBWqRpY+LWJ3sqtwjxZIfHB8q
yAofeCa1Na+7qJUcedoniksUIDumL5hGcfVp9nV0atsJPgfAODRtEKot2RPk+EXH
aBqkxco8P22AZ2Q4b3qfDpOdgZoa0/yQ+ZQEag2MgN9pysZE0vVikzybhelE9KSD
k7cxQf0REDk5ORMPc9rb6eYE3YqbjCKL4Y/ymOvZo2qo5TqX7N3AO7y/7ZLyT46w
YWxozUP/9d2D4QW1t12sDsMYe4nHQAjWUjEn4hfK2fTDlr31CTjIt4ZYmDkR6Vpi
ECZJCCDWBuKdOe0RHWnMmGwjPYCpWV3Aih5zGgRhNaBu0FAQAsZzDjeP5pZ1CaFJ
mHRD3VtxL7P5eiVzH3LGlgqmMUxv4cujPty6gsmJlgPziEFSfsFq6I2cwaPMcKWz
8GLjcwln6AYxwWkpyDLtrjbYNpDWbDB/i0An41iXzXk6/m0MptJXHn4sdVUb3PAm
Z+nx5HIuz6Z11o+b40MZhgKC50pUozo88XorSKizlSvscWRORo7n4y1I9FTTO9xS
AS7E4qHmXj6Nibkg49MD5onQHMTehI3zT70P3HUmmKrG8G271Dvk8SxozcFx3mX5
HSz7X0mBDu2va2PuK7u5sfKcjuLhsxDDIeRUaKaojB2NFSOmzGdntAdjQ8EyFPVS
0or+avWi1pqvOo3kafQUbjvAyy0NmVjDc3ApDu0WvNsidybmDJvw1/3gx/8n8Yvi
XRnbc9FUyHclJDX0phYyn2p1NSDaKEHev6OuqNQXUXTS3/4PiOHPGM3dlQEPWB5W
21utG+ctyDZb2tg3RnnwCVodLH5sgf1UvVYfuLe8H59TXYtW1KZK9HqBMHFLY412
+lkVxEZQQ5pR89xXI5ycKN3NWQDBnbYRi2N9PV374muoZOpGQddpV0ljmuDcbLsP
nZoBckubx9WHnxwOKYecQa78VlnApUSUAMuOyfMQzodSleaQMjIokhcHOw+IVMG6
H825LNOk99B9bKDBcTI7Ktg4exGVdj4kJ63XgMqtPHyEnGpCgXNf+swkgyJ6dcVP
+3kFd2g9SD6Q85Kwph1j1Tk4cJ24ipxO3bgnV8wuZeRYZ1t2HuHKITZvgD9skAKS
4hgcBojTVB7xZSVyrB6dmWZmRpabKbtINXiWI6MmEO0i8H3JHUQazvOJ7+Z4DFDq
vPIh/Ywhf1JYbeQ0HWWTcex+cOoN0YrijdSkobUMWI7uCUAAc3VPMyUSj86c8nff
KOAjh36/ApGfwn9/bQXXVcSuwKgPbYrN8mrp1pukN73GxOmZP+B2FKpTSHPfd8UI
CrSo89zt4vSjtXrSDpqMJK2mqT3yYZGQlkrS27EX9JYG/OPTbljynH/VAfnycFIS
H+3+tXduwR8U9VfaR3cn1OoYfIwdNXe+bcOZVWR21YGECtrODRGeZv50A/0ZTIsK
vhLPD6K/b4ZtHyTOlKcLt2E4NF9va2Go7ebssojKuXTbf8h5NX1vaZPf8EBG0Vhj
8jVSud+OQrceG6XAIsQZdlqkk0Nm4T21D3UorhFXvItaguoOPQksih6aFP0/YnwW
SDU6IYtfo+08GR2alSy4XX3Y8NQGHYbbLvQgpHDPk4SucNoMTR443mKh5Koj7+uu
vyI40NiqkIsdUuFQIGIQGhexRjQJt+B7yctPQCw5TONnYGuobf5P7o/1sv8LSq+B
EimIc5DD3GjbxnENjNOnbBmW8bsfSU92AM4yQR0B6HvhL3s6jgNF2WEewKCQTnkG
wHDuNNO7dpf0d/Ew4raJIN9JjppYW992m6WpBgYKmJ7jHer5R6bepBK8v3Ilw+yN
AFeRONaWhFh8Y5nKf1M1mnTtntX4Inlw+P4FmsSaCyk1R0/ldvqR0oMunq1eQrvN
iGSvrq4gIge0cZx9L0dL6hV76zySjbhBLppXXTPgj00PcmiyUiszXz9pu++U40j0
9tPrYLSrN7xUxAHhGgnPmuBPu1kYiIPa9hRR2DsUbiMEWq5BLE0EUiGcfeVhh+BT
nBhYbXQKUon6WzO45zx9LF/peienC5lyJn3g97d/oz4UFdsbFnO0vVkbFWEHXEZs
0ietshv8y5bsQRywEE2GyJZuhqfLo4Jf37aWBd/+4AYVpDaSsRlaxB1w75j8VZxQ
3s7jNSotr7bO7A/A+OIrh5x7RCXIsNG7zyCXUdyzMYGnFZSavrAoscPAt56luPJU
1P+YS9eufqni+LEHJkhjFmaLrfD94YzssO0NqTs1OCjgRIOBdagDEpoO1pYoFLoE
b+XqwS/Ui7nKnA+YlvWZ1Wft8mpDa1hGaNQSadr+FChrYnLhZKfi1Or96FmAGfNX
ZXLX9eF1p6WarQAP5jEn9jUhJ/L7kG0u9CrHKty8KcGR6HRMQlvNNCsz6CB+/l7Q
8wMWxfBsoVSXrAl18SiuOW0Ia4nS5+i0QLJJ1eBs/EJXhC2piAPjtXmmo3NIyG23
8RcYgQ993IdqghtqwOg8ByDtSySXv0MasP4GZwSUpTF6yZGobyI9OZzG3VboWY8o
d/3DCXZ82ho7UL+KFyDkH9n4fgOCWRJxlQ3rFOUSDGMLf+XlzQlTvLhoBtVzaGqX
7OZWLP3ei9O17+UGqpJMMq5DTOxezkt6ckwP3RDBSVUJHuvSS2QgWZCmUpCSUquc
hNal+XZ+hRD+Zxd/xhVuvIhhBwfadksYeLdSaWKvOeEVFuTltjLXagwD5i1oPnl+
gAQ3SvMvWESLbP+GgSwmfcFlh8f/Q89aSy55MPk/Vw1Rnm/3W/HRoqY9AwoqJDup
gxEMF/C7dnARuVrkZ0Z16alQWNicjTfSXH6cpHSnjPUf7I2OarNi0eir+DOlI5KN
AyM69m5MmXnVKq0MH/yaqAUUAt+lSqvvVH/xV9Ql7wgMDugHQ5AA0IpSfAV+3Osb
j/Fcc1qQRQP6Lg0dW3R9e8FHzn6mIauyCtqqTPJ+vcS5LPnk8AnvVrE+ZP+jTrob
SqMGeppKjGo/6RyZdm6N47spJgV4MfEe+jcpmyUttOrWf7KBTm41S8dDd116fpAI
BkLaLTTjL4/HIZZ4cxKjezT+2IFNkt55SxO0/G0Ny7or2GUIny6U24TDNy8hWZlm
Z9ZI1XWD2D9Vd8qLCQ+uFTMuXUPSydzNYQU0ewaSWvEaGEDvqBYUY/KIjNmnSnO/
Dje+wjQCmpVbzL9cFEQ4asiZ5Su5VErDHGaLCdcUmWiKSqMSv1d4TXfI2PYqVhZq
ZA5u0zdCn7jJkioF62rfLkrMTuv7qmk4UHIij3prRR0PH9bPFEaHW/oBgo/z6jz3
9cfLBHgQFWFikPzz2JGkX7Op7KwpYb9MYDsk3Cx4bbX1egpfFAaAhTAmyq9+vY8/
4af3c1RX0RpLZ4/tS6rjzqjaXmetSTEBtUOhM+dlXjMS1BtLIatTv9cc4PmlqWjp
lUqF37qSDy3eRothH7LQc2muVLj7UQewEYCCMwX3iIlWkAMmhCYb28D69WQ14KRx
mCIHrRGupDo2KZnnWf8BU6Rq5XMYQVmWnysmKBvWZT7W/YYETA3GSxhXfbclF80N
P5IdNufRUBGbj7B9ClVTebrRr6TYO7pfgXcpcISirykeP+bYxJVe1v7p0twuiffn
nBun0uIo+VbEI6a9sHYQdXYzXiGquwwtRyWM1p3OQJLgqm726oUhMQyJtEgT3J1D
iGwQ2PDkHzFRk2jCcWowDyXDpPvmUmtm7MkKf64Vxvdk12S/Mc8+yDUmn01Na9Q9
syETZ2sBWcYb7XfDanY6JxjkhJyN8bjN0GWj2Qoejw3kuYFQMogsTTtmECyJLcs1
caDEj4ZBYO79jTPcuBMPbUSFT/tfW4aeZB9MfQqhXIqEPzyT7b4PES8j0euQrspy
J7lBpIQSyfvpKZcYkl4sqiQbFkP8KtT/odFOj8Vv4a7g2EwrmIHzmBziqgM9rRhd
qqPV8hNN1mPmUNXNizLC/pwjnUAjGsQpiR8Bt0cKAUIJ39Z/uKlyO9iy3LeAj4BO
FDEW716g74stIIws4yzoyoQ58CkE/I/9+5ppz3hw2dWrxtQodv7yNY8I0WA2URdi
5UhPsnPcLef/0e3XDqftBy53Evwl5E2zEh8W2h5qRM3Icjgs72uIhdfDnhc0xwlG
vXNa8lMT4W+6G+HRzGUr2Ojyi69D2/Vs/mk8pF46JAUrbn6fwyxjL/uGJ/GHjMpg
j+8nxQV8RfNn3dKfFMDvcCip8eUrS4u9XJpTHqOUw97XPQEIs6JuVG2mwXgaajl7
Uckc/Hi0kW0sapi7ESq+0uhDDo3XnZnaQ75ArHdTGzteXmD2acJE4QcqKlH3ajSd
bZkirt3TVkN3udxaJ6FgyVv8oZmufKJ52mnEE01e0rVCH1i9Gs58iancXJRj7thx
NgRVis1VWTehkqGXsAUAoSLzQFN9R2ZpVdFJRFjkbhxrRGkmXaN1DnM7/cfAwZvd
Oj125zYFKI0MTCyLCqRj8U2kNi9UmGi6qucvC8YyYnGLOBT3YZV2hrmRIlqPKMQ5
hUa0UJVz45pJJvIzKNCL8+CPpgzNErsmXP1ajbUnjI3Qu4aqnisY4MnXQ8GPxjTt
R6VlRyqSfsuhUlduDNRL+Fd4owPEjoLKSlnBKmg5sCyVpWFYWkIeu6+daOykLbxH
rxObg2MOhmLmjVamgz8tYobQsjfKcSW1qkYeo7T2KIapeoLojWJTp6uqVI46FDfi
Q1IgHly6cHIxYRk87GEi855CoxAmRXV9HYNrrkaErZMTMuKAMQcYjld7Wj78UdtB
fvX8lTneGGMA+aQY15cmSJiF98tN2seLbAYWgNKucivB2DEQX8BgsDNltCO5xO15
QyT0lad6CM8uBMRmfQSOFDflzGk1iksrMplV4Jrc4eDJR2jddG4nkljn3Gm68TgI
fTXzKmF0WICpD0Z1kn12q9Gp6yAVfV0qtoJwAVjWa5kMOfBzQkncdz6l0U2HOorD
9OkSTSlnvkXOP6qOfgnFvr9JFT4eVz9tYRf1GJKi+GyLaanCwk4udFf6VznJuX3c
p7YUt+2Nwdn69ZMjWUkZxt6qDCtrTMiQ36if5St9Onuz8Hh/NJkrO4+Yh8hIkGF3
xE9rfkQtdSMuH8Y9N04/UF7ZcRqV8abQTwyFriCDHsSPJ5zcKVwZJ5MKa6/JvF4I
Olkm3BCU3livPUVyectazr8LTTOk4NFsutD20k0F4l3mM8GajwooKEcCiZqCzaEn
BEYbrksQO/SFawBSsNVSbCS4s3NcksKFjOSy03/PhbXcWwUEQKq+1DRUswz0gv8N
DmLssiawkEAhhOesvmS/pTxq/Po2WFaHOaW1JpfcxYgqrNgmuR26IcZ4xIVHLtEW
8qzWOCBHBoe1+ZBpa28Gzd/rVRydCtaaGrnogU1kyWW1nuywG4mXkHWBWjMyUn6d
bBl5/rWz0GUq0ZfJ7hWjEnWwCNxOcFeFt0a7DPbNBxatGSD6phL9iR/qTzrpsZT5
EMKdU1HzfRJ1FsAzSfgWu94X2ZUsvdzyAGcmUYAhlfqNpv9Xm07wrnlc+Ry7f2mt
vGvlwQKp+KSgZ2RxjaH0mJ42S1HXsuxDP7aR2+laciGgqJtBTXoCjAJcfUseT7dD
8FmG/wI+0JPMfLGcb+Qlvi46nMgZY2COz7iBsDIrYWz0KDQBYVva7LyAffYTZTdK
UfmXvPQgNatu+k3sY0Jjv5972duacIX7B77RmhXrtCGivetD4f/RRo8HF/HYuLZE
Dc6ZkfKklVU2ZAz74bv9E0wcZqg4uog+p5veur2Q42G61w3j2rFvfYqhHsS0oaxI
ICfpsZTXeEAUFttisu9fJbjTw38cQhek0gwC5LNgEfl0qzA1aUAepI9of2vUukEw
e+KoDv3K6yxlJgzWFDM6yTgSwFCnL3OuYrLIxWijIAJzoyCbIrn54zaaMrLshXvx
PdbxIzwOffZo25DZ6yUeDL+PTMxu0TKGaeJQi+zPckwu+ou1QFg/WoE4+ysofaSp
SETYU4wPwTxHaiIOuPsuhyHno7GVhzq4w2QIBmIb78ZUAJtIguFMxrg6PD2ADQjw
5WI0o3IeR6SmDbawMb73usO1WLEAV59I5xepcts0cvPlK3fMxG/NBcyAOt0w2GQo
AcZ9uiC9szaYR6CbzJQBBWCYbN9j4J2F8JW1tQwWvqjgc7MUY2T5v6+qbXpdqncr
c6MUI3HeBVoyuTTjZ4B1NO9sSypmzDNru0hZy6Fb5RR4qeoqbVbYcEeTVmCtSGP+
kbFAX39UZEYxvrlXtMuD2VvnY8sGZ+th0Q70SIfb52FYURqMnPRMrHpsc40yd3cr
6YfsOsjYTWnvbBIFDL0Y8h+KkDRZkjtKzVYHQu4S6bmdol818pP5qVh8+tWmwPvg
CmDUhi4BhwWIH1EiETo0hqNgPT7pDBDVUUdraMJW+O7kzZWt3k1fApm2oxTAjtw5
gz3kXFP2vskN+M+Et917+48r1UpgFzLSKk9FeqFTZPIo0PMNohKJcpxJufG28ui5
FxBHfTrBlKXWClFstf6zrv8oAJh+G8Kf4QmPdVY0xYs/Ie9NQ9vmrt2o6MBCaXoI
znmfYxWJfN+174M320dm0V0jaRcHUBAGHtgmclNGJ/YI+luiTEohnYAtq5nm+ELh
SXsLlXz7yUn1q6wWgKl6SphfyCgZF9vnsJ7kRSAe+vhlllrtoAOQEDdtsrP1sfWi
95LqBYdBjkxtfNR/HIumWCMfNf6nN0EQnzTjPMdOZL+Iwflexj7H08SNyKmHc7zR
P+/F0VeXqFAZCTv4oT1KwfEDw+QKaoAvfHycVqxb8maM1vy05nFGY55kyfdbW7w/
w/oRQYewH6xoj3pY+aFkVUGgWD3/vjhJNhLMSIdDfRzUAXz2hPobs9niPDtJ0aOP
R1ckdL9w8ycbnjZX6z3es/38v5Op3ziAnEw3FEKWcWpwf/I4hicsYc7AmWkyZNHQ
oO4yTLNwNjMO0FfpUGt5ivQOsAWOtlZBE7z2QkZBHVUcS1jNzGm08G7u5m+u9wy7
gwG9nm/O3aU1QmQ3/Ep+ppsciEeMVbhMXM0/asoTlTOrv0kLnNk1Yx0LNrUa+wq0
DyIKgDl7kvjcUVMw/5G7WyGmKBUewp2W38ik8h8R6tYJbbF4TBPcGQywfEGVR16X
5om34Mgitm9Vp9nNyeTGa1djB6Y619R+1zFm26yP9tl14PAOKRmmT7ogM6bSHo6N
ktVexFdBIUAc9NbpoxrOgNboGqmDg7+TQXqfQ+tluIX3MwLj5L1dRKDyIu3RrDjl
6ROEJyvybVbQrSZgX5MWMhZCkYBHcoQJuCEPUbuLfujMxURI/folHwAaw1fj3xL6
APnwEVe4cNovipXot+aCxsTshMV9jyOxHM9zC+til9csNODysRX/EYD8e05lhOPB
HllA+sgN1WIiOUQ99PnKZ7pJGaXKa5DaS/ya3+eLPLkKZOAqp8lwEN5rjEj4RwqZ
QV4j/unTWcB2+dT2L1btrP12giffCX56aungYCMRoKwVynu8CHPgH8L+6iXFnlp2
YamNtQk/4BrxYkXZImXby7acoUkGVq5CN02zogHb0qmfdKhSEak+cHigi9drztlu
1ku/GY7MQHnmpCZ0VA3/goAw5eM3eRFHxbSBpi0tvPaJypi1H1TJhcYytE2xza9F
/yDulH63pg9OpRO6AvepXFHABKUpFFvxl8d0teSHlgjMRYPnJ0Hgkp0Bt5EGXEhZ
nq/tV5cRmfxU0WWI6QO31E4RYNdyyQDsxngcfVZkKVXu9AsS7KNy0D9+dyChcmRa
T4ZXEUeFiTtLtcO3ewdH+BMJ8ECey6+cf+ILjIrKXeP96b7xl5BMBMdq1xDW32iZ
susHVVzJFpIKIWc7jiReuASeQcnpBdjX0fcrOeO0UeWmTesRXOd4+ryH4ZMrJFFv
THIGyYIRqzRHovsmq2XECj18yF7oW+zMnzSPS6ElIsIfWylY5FUDE1tyWS3lgqzu
l1t2c+fckt0PuQ3lXshM/6ROnN7in9tViybdz/y5iB8YvseFEcnztwxCmbTY/prG
fmGrR74C+XoginyUECETrm3BDU75u3e13p2Lb1UXyxiTeQin37s56ia1TNHgr672
+PtadWsoO0A6XbGWPuS7NeIWvql6lDTvhG4cyHNjsFtJbgteB18xDgiuEjSYn5R2
JCjwNtKkhaGCULRSLZzb2ZfobEy+JNLxgtkqX81gD7sKGMVtgxYBgAnU3QNksfXH
xVAwtH4wCpOFPG5I/vrWwzBJ2RsaIOIjudBLmVevIdJh2ucwovysqV2UO6Xc2b+I
0/kx9j43U1n5QUbfM/9hY1re5sJVePJIDOsibm4ZDqJHzH1G0sp0Pp2d/jLCmlR/
MwlxUgIpIaP3dH/KjXY/oWFQ72nSi3GlNlhU3SHeysUWG+ZOzTF4BPAnXY4XSEvy
p3/7J4E76LHC0TTSURbtf3AeEbEvNqwzq9nIuOqsIJVgk8epmUKJo+6GrN32VzRT
fiJ388S68lHsyQw1FzxWAeZvjCHJfhOL+WnViaWl8cDMZFr/3Fc3hYg0cMzhdoYO
5HzpcasYijLpDMLncHCBOXDeClDJ/KcmkCS5viKcGG9uuF6znXKbBdrGGKFKbbvv
L1sMelPzDMUxk+nR1h84St5nQluLi1X+FPcf24tx0VzOU5IQu6J8NGf2Vlg+o7y8
CJFQ3HB+vTbaCBjYI261FoT9DoZXx8AKKty+ogzKRqWtdbduIxwBEDlFgVj7tMkf
HSn1fCgp0e4CwIpiqY1AkzxqcKsCQDvArBqBTONjwh1Ag//ctuBIGDL9irRyF1bW
hDuVIzHfATNcRXbBKGcVcP7bi3Q4SKfO2P5c3VVccQM7NstP9kAA7ME5Q6/Z9isz
CqWuhqT8e25+gOE1RMu1LSVzRRMb2CFDsdd3j7c5b+IGK1tyExJE4KuF2TR2cPpG
wOQWS1sDff8otQx4ykLvnYB2Q/oi4Rxs4iPsta7mebiWpZRW02jQc+GDmRbWVY1W
v/pRtdhwIAqFjjUFxE91lQROgwz4Saj0VPgy1LCFYHa3EcIdQFLFp+T8+la33vzQ
/WV7E6RyWY9wmZuVkP8wljKdwXFE2GjOpYR3GgDVFR0LC5i/tqvLxSonwxC5cArv
f/ryQ6s2NqAj0au4s0XOTCshTtzDXDjzmv1ltjOZmNWdr6xZAMv6Cwea2014VNWd
PcIhQAVLrKDKskB6AMiXVx5uGu28BBhW6t3nVtDx7dVgbzogz+1yX0t0iHevrPWf
KfVsJ8mLC+0IVr5+yOMoPWWs1qTwHDxp5X4YECjJqnaKXqvOEnAWSLbA/aZDlOhg
vkr+ZlbFVHyv4wSyr8VUtTiMHv7orI54b8+6fsW0IKumhIQDXHwOHOBbhhyIGz8B
ThTZKzijeCZkOe0S5YIORi1dO4Fe8malhqn7C62Uj2rquVdtKQNqQPAukAQGvcCz
bePATypz7CdRCKsPd2/5HfoTpBC9j/go/Iw2gUBtKJRiwf2t7OusNs8zGUl2v9Rg
u43jbeG4WB4upVzRgKKh06t9LVcOKzlMw3sRO9jiVsqzIbj63Wgc+6h+/+9OorJg
irnj7ZUQRySHdUNYkRO8u8iQFmkAkHRzY65rqUwQsQz+IgQtpJUnUbIdn8vnH8FV
jea7O2zQIjJzikTz7N2V8cqzbqeccfIvitWB+W/OyDfvtftG1aP1W2GHDWJNm0Db
5LVpzScHVE0HZig1HvgZLM+syA/GyrkL157dx7RYf4XQ7+cWQIkkXsqAWtsQMcOA
va9j0PvbeoqXKgZsaxTlMdYgoDOdOKeHsYdxui862I1HVXF75r632eBTxQghijlW
MIuu56XioU7f9yD1k5d8+wnDXGo4qksAUJDjxISRSkdXfjArldA2pQ/F9rJTzy3c
e+a4HQCF9m3HuehXsy9uwemlvxC6SKqxglWXwcZBB2zI3h7aZwMeZcNwcw7K4mnZ
AgPehuwotT4yBuIc/qbtpXsZpCkH3QLXpr94/tAF+5/nDelmgCCZLI4qMylPwtGL
z+6DfdmJJlim9OK/yZBeYbYNmnRcMCdndSGOMy80Hytu+2dWV/e4dG0ENWnwTTGf
RxpU5j3fUPstpsNjU//syDfEIET+J0+FPAZbHqcYffq6LL9sQfExEEPqHyRffWoC
u0nuFZbORZu4pklpMw8PfF0o/qJbfZSu3CQBzZd8ZIv1/weMERph79K4sVsowFRB
8WdBETiPg9AOGhkQvrCKHIfPhIOsltSdT2JMgcJYgo8BppX8e3R/pCc4pLiocQiY
zjj2EjEhnwSOG8Xbp3GJ3bFZYrcrBAhHqJj6TX7vpHYxlY5SJfkR8Qdc59wKZzxb
aSVVjUF+sMl1MUUI7+rKkj2WzMxoVEgjTE0zwVQmkK75nTY7PHlaV7/uZEBx6ovp
Lwxa8vB6atMYtRadsSGcbPgXC01yXAOkmpKF48BCFs26S2iDIoAj8fSWzP9QcY16
9ds/vJ7ZH5rK0ioLkYFkJiEqkdB8KrUlJgfBnMPUXXXOBCagUnqkfDULxv6J4DaF
baY8uyqDUrTCgxaSMEJZ59cVAsnqj9BfO4KixorYRxerxTFPeVc8ytU9htaQp0P3
vvgyi/IC2l0aM1XzuYRjavxzTfZpLqreqaMhmJwYt30+LcA6COeHEyVEBXbqEv6F
5c2eRsZEJk4mLdvT9UMRMPNTdNH2MONL/0doZSAN7AH5OEK3Qdnz7kCFAqXdsuCh
fd/I9uASc51wFf5SdoYKf4epphQ6KK/7ESIZae+MNMZpKtzGRJJY33112orwUrHa
igNT3pM3syg1c5LR7q2ufubMoPoZAkI7L7JZr4T5Ndcnd+hFz8dpNBHBXK0C2I6/
d9erALTgrmQ+b8hBCaJ9Ky7gKbMxbnWLDVuPI5G0Tt3sh6lz5fPU5Rgxtbd2NqQJ
CEIo2MeDcfUjqRwwHXpP35PiUrzPiA8EK5c+CsKGb/eBw7nyJWKBsrjttN8IKnJk
Z9YnrGJ33/kWeJCwFBub5zC4cojAhbsRn+WAq/e8ULgDoFuuqYeKXh0rcOHOu4QK
x443U/3lXvqqLSBUWhLMa397FstIv7cgL9LsmL8H6hr3P5r47Nx6tt98HxObr98r
JkSVyqrPgv/hD0dpLMV7DkqKhD8V5hTtP25TOnFMQiB5OJ6/E3lU23wfs+xUNknM
ERa5g12nLTXSfahrpcQ1UEzWVNjVSBKHNjT/LG4ibXxut9ZJkMtrEzptQGdogbu/
uVz+JVjEzhxDz75wh7+AHRKk7n2ZbXNls82sFT5v2fBcVkAZDogtH4h8cObhOyeV
8fUmYm6WMeZzJx4Pqa9OxqYJ9Qwo+e0c3sDIzuT8NsAARnIN3FA5BsL2uAgvz7wG
EdCQs0UiAFz+NfM4VsvwX7qwLkZ4u38bJZCG2bGVFzjcndoXGCG/SIk3d+yKV8FJ
KV+tFthGUsV8qvPNAo5i+pvJslSNQYpCbXq5DZ6nvFVFC3iURn6M/c1QIGa16ypx
haELyLo1r+eMrJDroZNqUN7EOxphN17JAYaIf/ERkYpjlryQCwS0d9b+XN5HkHXk
oCw887TiGhPhx0SofED3nsdrk5ZQ8d6bxmcXEBGWwAMpXCMijT1x0LxlGoHsX/q6
hW3WiCuUW+cvh2tqXeKAhuZRjSdix5li2z4eNuygogSUFj/FKxD5rHZz3MBGTawM
MDoi8B4rANJ3PjXT6L0Yc0whTxbZBaI9OAs/Nm3SwOgRVzDsX6jKjkYV4trvmgUu
NOc0cMy0gR6hrSNVF+G3BCIvQ+PnSAJsyaI7MNJ4jMvC5BwMXpmNUKZgbQk/qQo0
ATHH8bRjifeJNSn9daS8b03wPyfp1Yqvvd443uJAixWb3264TsjTi95KeCHVStgz
fWPNle49tB//KS4ZiYyjck6UzWOjQjm21VDIZZ2MolHK4qClzJrCWbqxOyEOdBoM
Lyi6C43td0UEiJtdb9D4m8utySYOIcjQGGCcmkAf06I0Iq5x7Ud3NDK8HeeoN4l3
swmPRvKgTZw+MlzmLckP9U6lJpR3AIQf+mfqNs44MQF+g3IoVfdYmGqsIRPADlg3
lwa891LU/SE1MEF7XSpL909k0m3YrFwyRHh3pZWMSrLtl8eF6wueFKWTGimJhdez
/zbls7+PIdUtJERr7OQ/hk+bvqZ0pMBEkRMECRra8NJIbckAR0zq6w7ofjc900/U
LHnNbFwXBxBHlUC+/KnO2cRkvgZ8czSdciMiNIltHkWbzzgb+gnR1X0ShSGP8vtn
LEz5gUgeuFub5oKFjNVi7CaCYnYrb0UzJ9Bry5pG3SNMcuKg8aC0/tRf4YAPRxPu
mFapmqUcmkbdVBPbShNnt90yRVZd51FFKSfry/Nwp6qNt4D/+Q7p/Mb/0usYKJdA
iXQRlHcjv3JmsLZARM7YqyQnaxAcTSlhYMtDZVk2zGiOZQM2vKn4Hpep8qJ/xvIo
CZyX7EQArGEjt1NRgmssjZ1STlthBAPa4RCtxQcvtxi+qVwuaFQg2+qgLqoYacZ6
Vv39v23uW5e8fnC6XZWiAvObk0L7nfImdQ6wWOGpUyZwbvcex7zm3cJST8qM0mDc
n8hL4um1FZH40gQhsaiGfhKHVHkC8Yl3mRvrdgsKLEtCfo5Buv94CJXXoSEY7Ow3
nsTTONiEt2AbWUACKPlfbaXyra4lhLggxarP73PD8j4tzCgAQb2qsZGTDAuZKMgo
gfpVItq6R7KBj1uWkg16GH7gMulsoOdTqJAW+K8GooT+SKemIHRmaY3/qbYuDq8a
qR3PkRQhazgGt0iHevVKkuzAxsAYlL332SjBnK2rjFjd+JoIP8prPNlk8T4RaFRi
V+xFrXVtj8traFsdbZBZPetvRHIULenyfdYF8DoVRtjwnG0FaoA5CSpEf/PPu6AZ
Z1NkS9ONaggItqSD9oZcMsg8dODED+0n03J65uQXncb3cQl4lgWlVYq+45DIkt6B
vs0CuMQumsjz8PaiHHjZtyD6FZKq1s8VzCjUmXYroiYhMIQ+8m2FY1+8YwRIrEGL
LJSi3e1Zddj16gqKLz0ZICH8/DV5l9ngTiSncBjZ4O7tLunir0AhL8GcNa/TXOsp
bEaltUEs7JVf+4mtKIFgnsrq5MGCoDD2LdXL3mMChVptpHr008oRdTZ09+oXzFxs
SPuOZxukounCp1qGRZB8pcTqUGakb36uXWUegTrtSGH6YnzNMMTtQU6soSBlC9LE
ESPUXnKE5baE67Vc6fjSneQ7XXBJZLtrO0ibIewDVhqwI/bJH8T/Q/UqvFe6maMY
etoqaxcxousi32Jf+dih8Q==
`protect END_PROTECTED
