`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gbSJgcFHU0WmB+vvgFG1mYM1NZY8ncI9QpLwU8UUy3MuhN6unwwHjcpMIPMnDSAg
kfyewF7w6pl/vC+RjYKJXMkcktzzYTm3Y4NJ8BwYrth70GgLFPS/z6LR9Rh9o8Oc
SBskGoXgcRCpy87xD1M8GHBsqiTLkpa762tLyfY+T72rz+gCTrKVSMoiB4IC2B3q
/egGA2dYTSf5HxV/8+i7Z7k0RxqdDdYgWi6stpcN4QD7ZSNbUEHz4+6K2Jj1KTO0
U+3DsKoFe9OATSNLmeop31IT++ekqKvwzxgIhwQbhp/e3GxGYGA0WXXXOD2lxZs8
cMyQicoqV6XVJ+RcsV9fBGAWUgG1+1Yy6kauE2wPaoujeT9ZasMoJ6/OWpM+wH71
oeFmtpM/AMOaeAuurh6AEw6zkV9H9MzGAprnimo1WXJ9IpNPR7fzs3yROOrPIzBo
ALFXSYuFptDILz+qI4HUR/pRvtVnM0F1PVgZGfulRJyIs9fN9TgRYHghznJdovo6
o+TtvHGHog9Bd2Q20D6Ji54mUvCCTObOraa/oDXGBaYDvTyr+yJyllVtiAKZ0yJT
0G9UPC2YY0WRuOUhHycbcj+FMNPvQBvo7eqzJqOObWVyzHs7bedXSkkU3Nckrzkr
euYsr/tFhDElqPa8ZeJnoA==
`protect END_PROTECTED
