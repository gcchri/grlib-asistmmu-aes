`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O/X29mvJva0EmmwXpSrqhM/qfTOk1JFQCfSL3MyrMcIyBoaqUfdXnx/YABylt2nR
H73+2+AwWRa0M52uK1rZiT7qshq30oN6OQTPnz7+lYWi5BgMlGxWQexY/+hD6R7e
aQJ0ywVQUTiED1L36er4OSqkvQowov5nUNhCU4OD/TBNh652zWKd/36O3CKWPfcz
8mag2MjpI8/1itT1wegoh1t3YqNa5x/pyaZGVeIhMJdMUysRuqTEQ2DRqoSQ/ea9
`protect END_PROTECTED
