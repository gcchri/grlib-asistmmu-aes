`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pvhL/tqr34/l5v4M6dY88gXAW9bFVabv730ZVP79W3OnwXaJUz7u2vWLLgYi1K4x
sK0s+fpRnPKZ+UUgMFUkxUUrnAXl8az35txisy6pjEUSXo79nzzYnIkzOKz0XLOy
1fSNwtiea9QN+wyxHMt1+EfbSmsbvB3i//SFAY0RE+6zukeynQlnac7mn/AmgzaV
OyDIixjTBax9yXCbpjDxY25kxCJSGlrDbl/pkNYioLQ38eq9fhJcgA2i483ENBQH
vmMs78vT5uOo3vBjuHDBSPPBQP/PCeJ+CVvG+HsdJHW4Y8JJD353iRWk6qgEwuWy
BmLMphwBYjtFMeh2i4Sq04JnJODO8scLmzGvFCrG2pWEZXpIMkv9t2aSF14XMkeS
8AnJIHJwEibSWGdsC8v9spOLLmsB/awHzCYCi+VlwGY=
`protect END_PROTECTED
