`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/nFS5nF2mb3+9HaZWwY6L/ZU6nwFqzvEyKoisZRLPmZ0evV2ePLiZXIVSgDPo8DV
3GYI5Yl4SyDR+VjY5OBsEZdqDvcCQIYZC6VEhclW2VV/piqddjXUYcRp31qt1r83
xFAY9E6r8rjh5HiB0aR6ufNnJd50owVAhb3ITxmRH3Q48inUKDFa1o3sJJ6WVIUY
3c/QkYo+waXr1Dr0ltwmiXUvFtsG5j3Odw4JTG91vSLuB3kRN4lmcC4xsSoovpZ4
k+ckDDKRqf2sL1I9XkU2zfMY50e/Gpcwb1gh/DwJC7raM7tCH53n0hoSuDiKY7AU
a3dv0Zk8iCKwL7aLVwviaruVrD6gejnEgYlT7fG3qZA5zFMGQ/VLHRI6zhHNqOAM
uJ/fiyH20jO5woXA1LgJlc4gqk5qA+z+cYZieK8hvSYYsFFvKj+YCw4ggm5ckYC2
Pmd1Fpyy3lYHRQMAPNcAwg==
`protect END_PROTECTED
