`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
faBfEBQwRZLVlj/gZsKb2iHQDtgUHhoTftsx9P0YqSDzXFqozlqEbqw+q+vsAFTB
OEdHjoltS3igmJhqNTXIkslhIVMSFnnKKtdRKsaf/jopAEpfH3B99qoOQBozaaTf
J6bZzc87aYyz8fSQv1jRhYhlUlwyq+XAIZZFPX0MvtV1iMGVlSdskYAX2xl5zkKg
wD61FhPWDyBAH/wPUoEZZRIgi3F8Pjd5MREJF3NuXm4pRH24vC5ncPYdQcnsLDx7
XHdXjXXuYtTHxju61fZDMIIBu5aV7rbamL3NakOlLp+ifllxdc9dqqMKAjEVcdBK
SpKYyVXy+MYrVzA4J1IXAT+Kk6ZSfeXBxeKeBtYBl6h/hSmI+JGR7z8dHDQ0iRJS
DSayWlP+IqTNB2QwvTVWbg==
`protect END_PROTECTED
