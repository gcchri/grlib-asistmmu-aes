`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bqh5ezu31qLS9SkzWC/1aVwXXWKZDBeVP57C5pnJ5KsGHcrfgh49d67ltRDC2NsM
HDU7hwi7YbHl+5KdEU/fIwEW4JdSYZTTWNYripJXobVdiDUS6GZaRiubu7R++Gl5
MxszziBdyNYf1rjqAOhV0rCQ41JSQH+SPwVcvTzJLNqbmOlMmjpJ4WO2ZepHB3uA
qoAQSnukxrgArEnX1g3YL6FCca7EF4d9fTQkyau9Nur4rUuspthqrANRvB93bdI4
WnXyjo0eVYgXnj3l/ZAuyevb13SX7hcgYSbMhE2OG8WJgWYehREE2sy4JHyTi16L
4TNkPbyEWY6mr58wVUZKnDux4SbXUeDlye3ipjXcFGEtigBNxwdRUHdOouqIzbPC
sWoZrXGRw7q3cZpJkLDtnHrWX5SsDI1jR5iuKQdUJfxEH69C+8HZNk0eVUy/C6KF
oIkKN3lbxjF1pcuGU3k0lXFk9hJS8uLHwVwguEyWpSLVHzvOPCIKkIaPQ0hmDK1y
tVKSiQr1wiubTMfenw9ez3fG+pakg+8uZauFb4o6jOj64FyVYa7+Q0GZq6S9zANW
c3kMO7IU0ZR1bMuXfKqqskh82CyLCtkIpEoQ5Dae/rE=
`protect END_PROTECTED
