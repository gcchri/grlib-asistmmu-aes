`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EkqEzRJ+lpthAIJs4R3YANeoZKykjVZ9/PPqC0i+cNsy6I6/vVGA4dEh2ypgZXnx
FHW5XJ7dwDI6sJEjQ2CYp/BRmov7w7fdvQ3v1ZKJgIsN9qVYqKO5XtoFrEqp/oyn
0bnN+ypCI/Jy5CmqK5ZzCTELq6RLDGsKayOtjqOHsBsT/fw+ld4GLZEMbSViTnAd
c5kEPSf3HmafviTpKlpRHi6EV0vtNe2TNTLXTA1uWEwsSKxntNJthzJatPWsThsZ
veKMAtFEATfo+TLEsxDWr8w4FCXVy1Jix/0uLS87IyL6k+USINrgW4Vp1yLTDAbv
t3E1W8Nuin6Yna/AnKPPEUf9tijHy6eZXmeqtHADcbsoZH/cetjdiJ9EWxA2hB+k
2GFFvb0qhn0VRgHeQmcmU+ZsK0BLT/c0t8iMbMTsDbRBip2NPe2L2cm/01vnRheD
anhW5oHX7GHHPBrjoG/tFhNrRt7TlqvqPvj0HHsDvAJO6Ip1ngd+sIaOQEKrtHeN
M2HPEkQMt7ZHzLXKxADSpf9QWiFzEXRPZir5mhSAA9eTgM2u93IKQpPVmNsAiGRx
BuWjVdWLvrNb3Pn3ixIC7FqjAxxI7RB7wa2g8Or0/fM2EsK3MxGAvQpQh1X8dW0M
AbtXFeIjgfzglSje7yxIX5LKOVrxFAmWzvK8v967X6PStgJAcGFw0mf28RRuYX5w
AMYknL7Zn97e4biJfeXyqXW29qVkZPCkMVqII4j9P6k9AbH7lf0kCC7E6Jqn6bVW
xbKBag1KWcTGHfgwEUSvY1UGxznVIGwhYnlA/HXveq8MRl9A7C48oWuv/E70NrFi
JWigDRM32DrT7xdJeYtubEwBR7NWlpNrEoTNBSDs163Yvi/SEhVyL4GAxhQLyWbU
wIgYScCghooxPs3nJF0WdYRo5hQZSWJBq2RELS/JiHcaiH8oHdX5n00O1b7547uK
LcusZB3dbzmmhN93cbdpEQri1T0/N7mD33Qv41gOz2dwSkxgkZhbNyojjLiKsVRV
xEQ3Wsomh7gEL4P0QNJ4TZ/o7d3DhT7C894WngicGv5hQ+FAdGbZ28aMAiFeOc4y
66EcTZkIBjTLBY+qaoPavWtSFcssS7KMQ1L6o09bDLDfvj9SZlbktbnDJEPpnHN3
uEh26gys4FuhRAMHXQJaTdsqLOb7KAtA+AueFcteS8WSc5uriMftogAqpFOl+GQr
9ULcHl7MychK6CP+2jkkXkeOmbuEUTQcgwHYvzbIm7aQmkW/iTRoE1S4xmMeL5kZ
wEb39Ok5kQVmvY8Bq7bclZUFx1c/LOsjjSmHfMBgJFdC67+VcDpHrwjrNWCcrJV5
OSR8foYCwlX6YVTK9fkjBsvZUGlvRsP7CeEPZ1sxUEc83b2rt1TNZ2uEHBKNvmii
YD0LAw6Jdr5DOJH6jsOo4j2ygyPrG86zMW32ZFEwpHBY2qUkjOf5F+uT9W5iEiK9
CMTIzh7u2AcJISHUP78JpZWdErLsU80pu1vKdTYz+725eBw56wG0cSGGRRwqET35
xt1rreyGliOC+eV+MPaXYfasse9OLHUlv9MfsC1ug9uzFleED7f7EWYaqBsZbxmC
c4/m6IorDq0vDVIIcDgisHbF3cGJ4gImKRrW7kiWQzjJJA3WZ64HokrekD7KYQRe
dW50NVdfN+ixOmiGn+NjtZfHqCodJ/J8R9Z3o/5jYBPGJVbuQSH3wn2rtccB5W3M
Al5kOBFhLHvIL6m5GBAM1Da843mGFAPYQ7vK7VfIknhPKTUFhEBKl5q/w7kjdQy6
e4rBsgryht1MBCTY1qEvlF/zlm7wjvMNK+Qdh/6FgNImxk5aThp0064ot8H5NeFN
mg5dtWp4QCMNUkJWdvSOW9869vnKb2Bl21/6r4Z06uWiyqK15tt0R5nW7TXp3EG9
z63A1SegqzUgKyT9+LlvrGgcX5SiVw98OGk3AJHZMfbKuiWWlmLekvKmCADNK362
CAEszvW8Z+7oBQTJq0CmEn3dCmEBzF1saqOYsYO8S7cx1qsjrh9COSjkZO8LcOAu
/fw7glrmjnhem06Jy94jyKfg0Gim3RS1XKGkLb2SkPhR/Y9b2dyomMS/XwuOikqP
ZN8GX1K3YOXeCABegVXfStjo0m51lFpRCBC9c3ESflxhGjrFLe8adGGOjUO4Mv8m
UHLWx0/KYL5GytLoQ/Zlb3mM2r1ZG+0c/3N8/kmwISe/gTkhgeZ0a7kdVc0DDsw9
jv+a+3fMS1iooj07VYfWRPdAtGZHXlGtDCwpSbOgh5CxFndVN5iq6Vf+4fgsl7rn
7Fiprbgk6FW0V9P+Prer/XLoVWaxO0s6/JAwydeZ3GP7jKunNY9G73CsKcFbOCX7
dFpA4zqwKN9RH5+71BtEVP1YB6iC4LGqsbJggJCbOTcyE6ukGJ6oWHbls2EbXy4M
xoo1IoIfkSvqeMbK+kLEsQcDWTIhUWGQVVFJHHdp9GFB3MhNjRv02rYWVHkSTN1I
wqtS4H8EWCyCv8+0q7AYROq8Cie2YH4qLKkD2BUeG49liRzkdFBRm/ZVQRNg7aGN
MaiCk1+2QszTUxr6LR9yJwt1+FH4jpEIOo5YGmwcUSP7WhExZNSCzPGsvBk21JH7
tO6BieNXfViZY/e+fGu6kTwNqVd8lS5GWqpxlaJoOkH2g6VY+EmHvfuwIQ1pdavQ
B0k48GZTGN9pq9La4Lz8kB94NFxUk7HtxegtrEnlfbP9HuHrejX9Pv2OAo1d50/M
2j1Iue7r898iFLZjZkaf0mM2Y6jCYub8HXgWrbVWHlkyqDWRy7OyDe2MLYolnMyy
c4heSaLSqX/oT0AHNDfY/JyZ4JzWmwJRkXv/f61wdp9arPzpTeSjDqZpLL9f+D4R
xupfGVkXXXQiBke3yJ9Ux07ihuc+Pwq3vEBaFbYZ+5TLPpoobeoAXxyAp/P5Yl+5
Xzhumrhypag3ZW/cSwwogg+nt+4VZ1ru1JQBZYdwZrgN2PrJqiL25JdHWa0t/0Hx
OpDbH/R9TEiyCy0gM/bNHbVyHSxjWxdzs6KAhwnTK52wTvyGBz8e/p1I2A/mYHkW
m0fIaH5LTLmVR7GklgrcafFL25YggSErGGIhPFtIgl0IwV77WJaCAFPUMbUY4vv0
6qD0EVSwgKEe2z51VSoJINzjcKa0If4pZUQSz2JWweJ8ADH36vAkZfx6MZEZ0uKe
EyYQv+tggBWwZEXfQju9EAC+A/J7wRdngshUdVrqKifGHwWUbFB9MBP7IvTWZqKW
XbP2M7JMIVHqx6X2iC55VspF4rKgo1+oZv1Nn4AOczs1haQVXE6zOfU/BQI2ruVf
B1WhLz3oTH6BRVisJ2dhQ2GsSPIUAsmDw2HfsykfNhfmNv4rjUkRHrMlAOf4OuE+
hNJ26FHPbvcJ0wG0InlLMKUYUUQzg84/7j1au2LegLFJeWURJCDaQd8IYuPORfET
mayi0plnZ9YykJOZypg2q21sZeFuGY2kViM08z6k5z8sG1EJE+RQcSkohOCvo4yd
T+27zJtOTV1vWAjVKNOSeqrAV+mPWcy2/zc8wE25XuoP27nf/I2mDAWl11x+KuFN
2+5Rw2bIRM9hYYneCtIkN66pwLDqMRP5PqoFWoxtMMSDTOFJ1Aukc9cSaCLwL4C6
uJtXYl4kiuCZEIiaoVHzaaC2KxVYNqb+DzTrSaJ8pHpZBMXpgrLY8/qWUighXDcF
IONosOULHMMN3as95s1z3YaFLDnTwoaufVqYUOiM/jbEFkstQNLB1e8yfRJGQqMM
8vpWtqgfRSykyeE2FPCE11rbGByzncmczFO+GYVvvR3HXU83oT3qm1uHaQorVkQ1
0Ol0qS0eSScWZOpAJtgKEgL+O0CQeWGqXXue47B+PA5lk4mZQbKGFXZksmQpjC2f
1gw7COhcM+K0nPs0x+pYifVYeudzQPs0ukOgwAp6aEFea8rCWwByW2RdQM3XFZIK
OuWLfh++cISaX/z1btWan8rt/VwwZkU8hKNYmeeNGPCDrBecW1tv+Qj2OQxIhnJA
7Gtsq8awuFa+9kaUVGONw587/TufEgqSV2mqW3bMNjPCo807uveM2tx6af4QseLs
0FxzaZLSSJnlcwI1zbjwkMZf4hQemaioakT6yZ24NeV04DMAH7fLR377wkNxfsMk
W562pPy3MP/UcYALOS+QFNCGvi2whHmDzrd5jWJexfdG9jse/ElrKi3zNk+7nxKX
3ln/zH3KHW7MT4mFX5kiKuAOH2d0CUUYC5t2MSngGszrZ7QnnF09miQiU0Ok0DRw
SaDsOtzTin0v7bNKNrjgDsbIL6sWBKoSmSkBGUdUdq29ezKQIhYiiISk429xZs2e
2UiAdqBX1s8zw6hwOm6Bnlrlg7WQmhAVQP3pV0nBAP340Z81fXcHnYoaAw8ttRlK
3x+mLfd6001e2yPWeED6ej6NqAKT95iQ+z4iMdf0qbHRepKLUdZ+sNKhPzSRcuf5
jqIdtu73uGrwwLvH91jmI4xNDcTnirjbugSWG9uQsF6IJ9tqUuoUnLSuz2skCVls
hvd+GfE1V/H1v2CVhnt6nQxnv1V4n3GqMWT7OfqRBXVdxB2eVA62tdlhaJQQSiMs
FyuS/BecTTg4pp0JBJo2wrX0iAwNnv/tMIPdGbzVsd57Xq658FZHBjVopfFirvOT
+LGxcXy2TmuJsoc7tBd7bJoqwFH0mEQ9akwhskWIPCrAZKzBRD+yeKWmaHg3Cc5B
VaqCEra16uxg1Z8LbX3DFBEY8EfM2Ze+TwGl3mEQQo5BinRHa7KtaITMKv7/AuNx
PztZzPUlOzQzh1vCkhSd6q3WD0oPGZ/Lg9hDerRXixjGqoI4fA9840y7IF8riqyV
XSvGocvVD5OUt2KUqx96lCCpMLMKbvsRKS5X1r2tGW3qvbx+b9ijNoqrAO+e3qrj
WuUnkc8gHDgvi7SQ07BsB36BUKyvIiojzO5WM3cNVXwPAMQlKPzmp1stGw57O3jV
XzHfjIjxtxFFrwUTMqW88wTNzK8oaQNfFNNPlzXX1jN2FYhwm9ff7//Fe5UOuKKx
Q3Xbb3VpdM8ssOJCtH9Tha3YzzT10CZIQUPQ2YGUdRCKipnir0hU+x6EuR/FYaEI
JDepgijA4BGPBLcmcYf5fgZ+/rwoX4ucYwiYLO+xanaQ/QwHf1PXzWPWZD++ybfN
SmhH6Nv1pnMAslP/plVMhY+BmgRnr3NMtAYnltkv97RnltTqtzmHQW8RbQFcbqHo
np9Pwggjili771rCdqY6dsfREmJ8A8LWZeWlFy5jYZJRW4t/qtEJzC4/HBJJLBks
4V1ZLGstDAcYgPsKUdki97Rx2ipRINQft7Aa6AJlEXlGx6N+OL0EbzU/J0bsmTvU
K0T+0LNW1J466NCmhHtIgi5J9WdZrKDJXN5s1Ao5g6lD2kTVP0LNcCG+LhSzJ880
mQJsL2AvLnGeKhLT0gdalmqKZsxFkrcn5ybmGr0mIHQ6IgTVQT8p9L6ume1xDkG3
2WgZlnTLtk+mYQFJleUYRKOVMYLUGWrOm8ZFrobkIhkpjwD02zol2sdAz2aLIMsL
KzsHfeFMHKIy1RiA72Rmqcs4A8uUOey+aTOUFA954ngmqkY97NcpK0Z2UfbyC1oU
5Xt7KrDwvTjXtGoQqdjGrYR1A47pp7a6TGBycrW7CeepfTffMcKgw09tA3kD/wHh
8VEyJGV6y274woc4FhFTJSyT9n7m4Z35EAr/kyyBvzIb1J+URV4/oPcLz1HB3mGf
NzfN6U4Av40daSuTuLqgTGRCPadrNidKDQIlztPvjiFTb3Lv2ecJjfX1jBFbf0OB
NDcQi6BhA0UgUwhBkIBs1QJr+PmEygr+Mm0shLTgqaSyHYxqXVSi1AT6U4G1i3VU
5jCXLswxqB5ozoq882+MxgjQxKkN8SNERyuvk+Lyk/yA4l9OyJ41rxXO0/FHoC2Y
wp1FlUjmXgiHIhh0YVRG2jfyVDS0qdu2XtTUcrObGQP1wjnebjRjwJGbjpl9XVsE
I9lWtTMxhobBNCzxWxictweWNj9DNSKaENsImmugmHG8KNKiMZd2BFM3TVLQRzWe
C0gLNDuVaxX3Rap/5Fy8NtHOcrWft4PdPnbHt4aMb14YEOtiu6Q7KZjma1VdVFDi
UCNlLIWOBoly5KhJ4R/K489jTwoPdbBxa13GWKExM6r62aBfd77k3e5G78o493L2
nqmU2YUTiuq54Yz8cd5kdgDd4EnZcK33BYFGrT1FJ2mzSfAiylVksimcYH1SopPV
7cBkfdLF3K1lS1zM/8SOXVKSQqXJIkLEFvSMzhdIIPYMj36qyF64y0dyo/HwhOeC
K7qN+wb0OAL2pCqLRsizGm9GC4RDZdO/Zi4S0RFR6N16CSaN/DNBrry7RjEwCGux
+MvpUCpHhCRx+2uWE6JfVolI2XFRiLAuXSBW/vPzNn4rrVogZ4d/udwSbB1H7tIW
CqqSy/gUKYT96cmYCL/W6HRRrHLOCZOwNwUBfKR0Not6ZfnFq5bT85ugldARbJ09
V29lNWgFO9LDZkakJfhBftv0h0VAItha7IWn31P7YAKcwVsbKfwjFUnqkSntZ2tA
l2ndfe9wob7bWZfkKVZ2fEFKdH1F2zURWgBb5o3hrnDUtWqEr8ZsOb2t7iuE6Wng
zD7ak6oPG6Wj8NfgLibaiNFFHXasHZ9Cvhx4mB2zylCTcig8jPwC69nuBqN/qc8w
W81qevpuGf5MeZYHPnoQOTjzIRQ2WhWxwvSv4wLyvyqLco2AtJYbPBrWeap9z77S
L/P2Qe1Rt2FQSncwUzjgpfyWRqZzaELn3XElAr832t5tpgB5eAkVrheMhUs2vHjW
9ejy3SOMjn9rQab7d9//ILe8aT/DTR5GK4pkbgtTaymSErN4rpL+wYmoiROffqWP
3b3STf6+qt6AWFfnYe8bbFOFnHqzyAQB2QwrYr9dAHxkWtnzRQllqBulTAMaPblR
qIScu6WkWHPsvUD7jYkypswZg6WWIX2EdrUCn6uLaIr0b5WYddmM/ftw15DZla+u
37WBGw2QJVkBi7f4+o7bMllreVRKvQ0Qox62Dok1Vjk8819uh7QSF3LX5lU182Bc
YaCgniZ5UTyib3m2LiWmDu8YX1k3wKUUc9QDfJSscjtt/hDSg3oa7O27/WNptc0F
HLfEbrcPLUFq2t4OTgZPFAJlEljjcyTsC8XskcAVFY7fHj5M6/nLCO7vvhPN88/p
a9KI1oQg2GYgRI085AvqjOp8bbOvv1nI82gXdGOnS4ikhRUYypIogHftjOCRZMcp
WL3J0JEC+ydBdTlk6uEDS4mHQ49fdxiAgO90nNYfDRTalHvvxln1w4nqPqQ84U9R
jvQD2GTJaMqpeKtpJCPyFRQKhJlwyCT5yXXqCfggang+8kWTlzYoW5YabA7DYWIW
U0d6vpcsP9pLSA4G4VBt8LbWEGsvsd2DSR6J0U6oGKlrWSDoUr46i8eWQTtRz5QI
bW3+yCUIB9NBNOwkmTKgMcySqya0Wq0D4A0xx+HgTKhnkDGsomBhmY7y+QUgp3wn
EZUxF44RXkTU8Jjf/QIjR68d5Y1GzhFTEb9OL6zpCqjPscu7QvzCnePMuSlJNPA7
PuiqVAd3Yc86ra/gzn2pdHtK2EkXO9LMvtXPHpQnbjR0yQtypcuDfVS9Q7QbyIHP
k5cVpliex5JbE48Wi6eH5fnvcdB7drrfv0TTMLfZxXu8Y3ZwvItlTCLFMLErqx0R
hBHunvSBD9GhwPmCZ5mcHLjzHor5HuizmZ8hbgqtsnmbc7lBF5+egVtfKWY/ze2H
VqWVDo+DOpK+ZJrW9HR/aNnw43fdvofj7LucIc+pM1DCSFiD9FMQC2z3PUGizHwb
OTJxhYo2JkSp+spB5FA4uXbM79JRNcJV4fss5w3JqbqfG6SKp1I4iQ1OsSfK3CZ8
/p7HVBHJtVvZ+Q0le7X9fTSZFJrbf54/jnhC/YpBzmRa7fzr8S01ajIppPDHM79O
OO3DWB+ENRsykrD3ofR040bazfFigxdSJTLb7jtGWkX8slFkgq4VZMPyA2gvjr5E
zK96BJ3NN/uyfqqThAQaPeAb/10QNzV7hFyYaLnvrnEU7UYJ4Qtpt/6XWA+ty7wF
KXVB35op0bfqKPuNJwwA2SSKcHajFR+LZnUdjT+qCBx8DmYSgycIwU4KsydDe34Z
+0edlA8wFdmPDqM4FFkvXnNAoYAIb7zzGD2imnKRqsxQqg4YDS9ycMt4tbNR8GVe
jb3bkjunQfYtHEjXdN37+jMQ4pBX+/qFlPr/cLnGrogmkTo0A+PYniEkXLN4OpQ3
/+CEi/PEgJllMoK+FjvGs0rdbU9cYBSJvJZyyIj+VxdEBoT8e1QX2FSD7BpgnR9w
s3cnMYAVHY2x1JE80keiH+LcNCJXxFruVpIL3kVyZ62hgJBu16eZoP6KmKtpdlwt
CvIosjk22q8mr3cxVl+0iu5450LtIddhSI2JIxH0Ua4nDAqRWMytPkt2+9I6taiu
LnrfhIJbLUGEDQ9aGIBYEAQvN5Y76WtU6CFkRMfaA8pgbTVigKqLYaySr2w2p8Mz
VoE23oEyTDmKBbPvJW4N0Q4oT5YSa4yFt5Zr90juYSxkR/KQgB9CAtKEwxGpgFv9
LL/ZTQQIsYPMDttZ6iIoBid0Cz5FAHS+utVAc6rWFPkkLnyG4ALYkl6jUxgpAwuh
uZitqd4O3igvygipNPmH/aZ48ImIKmeWLm8hp5bmMrWbm7njUveIxg8CBGy2uYbs
zsQxoFKv/fbJjecJVwO81/BcKr7v+0cdqfeBO77mCCd+SLXK6jG9rV92yW4W7pMX
mP4Nv+TwTww1fxhRjVbGyRzGMQaV+zfSWoQj3b9V49pTk0bnttnctaWyaR/S5jFU
TEv2B2f4mLBQlxI96y+TMO/e0dfxFVsNhSm+mvCozvwipIpBHhuGgHZwJe6ZEKBu
1H2Ybaie79VbNppwAZDTSsPiFU7mqcJ/jKCjnRPGcJElX5kpET5O2GsWtErgzEni
eZWrz5kNQsC68bTDcpJ0okVhDqf7q/Fx7FlHIVX2PCuwSt5o554lnXMeDLQ6YRwD
F9vq9ldzX/jSqozGIOt76M70lfJRK5Vaf3zVTho3PPWr0CFAygMxm0egbm41HVcy
OCCpQNCHVGc8gyhvTC1lWkrKlLcICt8sKe1Skjnyu+e7aA+jr1s1EKnVo69sQhqd
4Jp5XMjogg9PjJFo+VxNtzLMz1zZyWgv+qNsk8qBFlFmK0+2CQ4anI+2Lr+3DFUY
6a6zR+8NyDyVHt14i/OeU6A7wY7rmPo+Hw4bwghXhD8XroM2BuPJF1jVf5C2dKOX
oqZzj+qBRY+a511Uzg0PoeXFrJULpV2jpRQJArm5YM9L9zfjxj+kTMtG8oCnIj9F
fbNrHiYYq4X10TI1PDdGwpz3qTL+LH/KYjJH2W7aS/WL5JiljDQsSGeU4jZCl11D
KrAPP0W5/Kf5QPcWmlVG8sDwsFFEH99I1qdKuVFjfrZEoJ2WOFg8xEre3223AmxM
FMf9NDAvF7CkcHScdfmUMACZXuEObDZOSEwgkSQRNZmHpITKJ5Jiuy7y9mMDgYDu
iV9dHe0//ezCHeDHBzalGd2HcZlCMA0TLb5Zgc4d5prF4lupMhvHnesNgUFixXAh
3elVnXh0L8FMY+eGQF47iqqF2gXfewP/2sfHy4dIVHzfJSbaY9oVZx7FUiaMFBzR
KFEUf2ObemeFc8ASmLaZvuM541a+40T2IYUVfwfkDBxmxIsoikXMSy4JoV4EL8aC
AXSu35MG/irqzOQpVAynFtZE9wtwGGkT9SiIp780p7CsXKgjrcOlZudOx5vQw1UT
p8rV1iQrzJHjIP7KOT2xtl44O0pGY+538E6eS2p6WykXmz/Hr8xhvutHNn+mQgGi
BfEeIddixG2ilVKTXy6lmMbHo9CA/Q+/yqjtUn9ELJ3ef4m4OIumQFw1RjXQOhOB
QjVGmYiziLQ29WHeywyf8cUHVGh1jtfhll1zzvnvmfowJVQqJKjcqUyXrCjBDuoK
p4CbElTjTIdAMqi8NMKeHGA5VrRPsRr4UHQgs71cfy85Q/QWOgLCnFCDr/W43Z+l
rvyhlvypETqCJfAPg3UI3jGQkjsmjaHTHJtbhuau2+ae2XtUbelur/BYp4SaF2wY
jIZfpYx2ghOqs3euYjLbCnf1SwsWgwO3FOI/KSPd7J9OPS4B/udTcXwxDs469zZt
hCUIesyxA3CEKb8Cd/Eizbt0bP63YyII4U0y9hpb49ZpdhSy36bsM0yFIXpDTXe+
MQrSsNA1N6SItxgBGZph0KBukZ7VsboF5fMC1yAWbbGXOlbhUNePX80W8SQgmMdv
/5CRL7IHFHZtMo9rnAIsLVwANUsQsb/PmbiCywH3wX79T6zgMciy32156NFbMrd9
V80h3S4JBnanIHd0wmG75SnpP63+clKuuYpumyEAWTxlJNi7DfqN5ktbGgK16Y14
n69q74oACrfr/tRIJfq3bDtTXYasIjSIBhP0ycxyK+rkSxJBKCXu2eBhBi4RjXdQ
AxH3YXAdYdQdSkvFofk1jTrfPUgbp2/8OxbiKT+aYZdvybyNN4J4vVDfDfyancpX
Lw1Y0fAQQ2J32cNQeCfyU3LnNp15ldOShUgnTDxFEuyIWhw9HWi2X7u8JBAPRNZh
QgbnF+dCFrg/gprqh1m9GIpZJZ5qN4pEH70qb1Ckk46Ssod7mot+1B7PVZHcjLv7
qbu9YtVuZvi7m5lC0WCqjuqBsZsMpQuyV35Cy13p6ODeRCvLDdsGwPfs0cSzqYsq
zEnSj7NwFYtYIhbpqgfS+RzCEKlOqyiRC5s/xQsIVa/DdTv7wK8hpnx9PKzDk691
nVbb1U42B4oNAh1effHfSr/HyKDlDTRkvYDl/dJXAyRITL4NIQ9Cql/Nzt4CmWzW
8D4lMAyhx3Q+386BrWVl5Uwo2XxEk4ySuEbZAJWB8IPFvRkcUnRrATrTKasgNS9I
ZzpV4dufBPusdqksLR+kJx85Q3/tF+QUlEUZibypsasXwfEVi0DfIVi2N51vZm0Q
dZaJu/WkOCo5Jg158WX3YH/hkUcDWQNKsPrmTCBBpFNncgRUXEGnfcF3k3Cxpe7I
/owc8EXcW9bHe3feXRm0d3RiSmGNm+HR42Qg43lhbIeZrGh4vr1fXolRraFe08Ul
oWafPNfOKLRDDr8tiI82KFHVG1Ejv11BcdUaGOTX4NK0oihMYGtttu2ZyRA1iryX
UbxJR91PuEQpRoXlfU2xdONKJ2HzgkzhlCHB8W/Hq2OOzTDk0mYpSTpy5jTTOmJ1
MCKVlsdIFh4MwZs5Vbxu5OwtnFEodyWUGKND3uy0Alz75xTTMwouoJNUJ4Oe62GE
kRwsBG1nIqbi0SYf/XWFqvrRc6UdeGK6gG81e4VxNUN3aSFApcE7ehu/hEAVVitS
zid5/G3Pq5fz4VK/c54HGQjueQc0kw5eMwXn15GU2eLDtKqxge3yDn3MSm+dIrLn
yEgEmwtnvRi1cGCpiJTzg90dLkOzjdzVLyV4xiCdk0asSjytkH84Vz6W9QmG2C6I
8iQX7EvASZDGbj/RlcFtxbg8QUXvZq6fsTSnUsQMABrgQvLb8g6GKrys8E5RBoqR
uVoOoRCPJ3+yczcvEtOJDm5CAN61yEYYeS5lrjSTdpI=
`protect END_PROTECTED
