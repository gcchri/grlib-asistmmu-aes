`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6KB6gd8xt2udht0P0eAA9zL6ErVEi7aLi+iriIXsKeC9HyD848Jv4Zr+knq9R0Tv
mZkC5VywxLTthagOgU84iIWIiPq1agXmk6/crAibsweA6lsHyWzb8N6AwtDxcCSZ
TOpzpjnPZhT66MNpecG6sOsChwwdr1e6sJcWX8LbNDA61KHUbBfyiRVZ+KVlMKX9
NsNRIjNMpbPXmp7KIqiFgHEeyj8x6MnaSP+fJUVBDz/6px/3CWNsQovQH6TBq4Bb
cTRXM4IILaYWHINlIQrYoT8IEnJlPEmHZeBPM7SXh4vEax6NbyKkztpHQt4MJ+Z3
Tn7KQL/owvRfHs3Yeqfc2g==
`protect END_PROTECTED
