`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/+mX/+0dH8ZZG5h9wpBEfr8B6SqiQdd2KSuHBB6Zye7e47UfNYW+qYT1e0h3ZzcC
duTKiRQk1TTV2c2VrbJZwoky0hfnCNZXQL+4wQM8KS84APoSH0R57nLLcxxURrZV
4oQwz8i1XLzn5zR0dPMR5d0k3k7PckVRuQcVUdxUYwk2LXnWXWN93MCgvlLrkImD
daKHqswwUGla9fAX8OPiOR/ZKslEmGywNCYTkvnRS34uMGjHIhY/zjvGo4iUB9SP
sL4TK/T+4T4xikaatvU0KCGHZZX59ga+bM5/eIafwjYS0jSrUdLo6OG46QAS3aB+
qubmDoUKXs5LoN4kalURTftuNS6v+jwzZ9nw5P5WMo/iZS1CuqZ3Dit9Z5Tqu7As
q0LGccUx4ALVcog9BMpzFZJs69JmBlNeH4jPNxctCq+sfBfpztyye3lJekWkUOGo
+mP7I/IkL+wm9lSMgP8Vfm5sWS17YWJf6YTY0OKv9I7ZeDF2bhJsMGlafvLymj0X
5KWLgoHnveSafpTRhP+3FsyANm3ukHxQL3amYGaD7ujkaDVmRpetNu01PhE5ty3h
TBWZaCAJvUqtZHGc54lahUGbZRdmk7KkOYadNmdKmh8zLkqm5skqDacMqwPf/REr
UbxIaCTvjfaOZNKoDaTwXKeh6dfGXKqZ0cLNPi4HFdPErZL0pPk8WARS2z/X28N4
sBB30l2YZnLoeXANoDdaNDz2xvUQPml9j5TCHHkmTa3ENb9dnkLFSJDwYwJ5m/86
d44lc3G5SfBV2/qmfees9dY8US4Zyd5HCg+AnQ4rW7n9i7iom8/I3wQ6ecNz7q3O
mm4rtUSi9EnX3ZWD2S9agnv1W7D1PRI5KJlT+xIfZmQzruaqgSK4ShlM5MQALlmS
tRggCf9QXS2AsP7VULSecNuicxPbMb+8LRP3Zs/cAjM=
`protect END_PROTECTED
