`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3vBZxKJuki9ImxtzBqPe9Kj1M6qRO4J7sdjutdRw6tUeUg4H5GuCAQouI0tJ1vQY
oaBBl50MM+cuMQzPQb9myLRc/NYWtF1O+4ksMtcL34G1BZRm0SGNh7APl3TTt4RP
7dc4nrfCuVWfXSLnXfxiWrqreF2K8TD6qN8Aii/67SFld/UHat7YHQpaW3WtI0Ut
Szj6C6ZtFsOtQ3Cyq/s3TgbXFKR55VwrSJsQ3PAGJHJB66vMpE7ypyriTvW8GYRP
m5Pp+QRba6rqzZ2jFpDSRjMxW/j8CsRFU9iP4uNkeDI5Nink4rMaL6fokBbH5FsO
HMCIHrHdDb2pbtbbynHEJjGsYXl0DoGPBRFW9UTAUdGUzWYvSwF84qa9UHpWU+NW
b/ZLTQfZzcRSWAv8YN6CNDOvRmg6PeZXGhurapj/G+X9RVjPdcnc8z/laj5O8zGP
4//+rOdFNTkBNiFwU5wjHqicDFIUmoz1b66sNrH+uw7kXDdtptU71o5GMgSCpmdn
kycseMfotLLEJf8E7wrGojNDQxp2DAhUY441bs2dfd8jbhTqfEZzNxqHzi8yAfEG
dA2sZECyk0+ih9gNoQh+5GjL3rM6LQOp6waWGCgggIW9TYPTqulSWJuyGMrJ4tkT
bHmBWzgh3nM7++3NAvNLXX7p8/mmUWKVxZ7AWnBu9RWO8CoFluwh3nTlQFJhr/C2
DAgkmtnXXfJpENuVkKO2zAv52Zb6BY8gECXBEL59i84iJr6NVGQKpWlgV5esoMEh
`protect END_PROTECTED
