`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U8ojCvgkazjFuUxjQ/LTtmDe51bpqMayIHa87YncM6SbftWWD2hn1C8GJYkHuZ4u
JQEfrrvrIBkqBu4SjzO7bKxx96wQfH+fWsMBoEJeO2SfGUlJhCOIXlFKwbV9W2/Z
mvPXmto/H5G8R7OnO12tjWkq6f88tWYgUdErehBnqRI784shCf77zaCkN8Oe392S
6RKyqQCX5QsN+Oghrd187Kd81GK87xh1153+Ge9jUsSwg3SXq8E5DsdKBId2USC0
MVnzXpbWNS2GRBNWOXl+lYJfEEoYNY7CyxitUm8U/XoKm6D+fxstDFMEm4mdOu8+
Agc9elHEmCrbw62Q/QLktTYuo8GcxJ619Zs9vgKbkIjtfA05pQRv8yziQfiib9LW
TVwJgiEIMHEWchDn8Cf770QH7cr/+8OFzITEHpqTxXIn7hZqT+D+yME8qw1eOjMX
qNw0+V1slOvNVcBOJU4W1QLken/Sk41ixVwJJmiXytkvdw7Z97q9LzZr/710QLmz
x1q6djAQ+ewxmjlNv+N56O4BAFnIp+nj0YoM7eFMisJSe5USxSSJwtkFRwqc03zg
E1rkHnGjwPG0JlfaGULWRMkl/9qy4T2v5jVoRlirbNxXv9Y4YRaK3xX4IvihzOc/
v0c+f0ndxHn5JMYXCo3Awt9XSQfmgWq1yJEpMZklJJo=
`protect END_PROTECTED
