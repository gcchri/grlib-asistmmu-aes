`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z5PJou5EnG1/hxH5WIXCe2lJ7A/LQM0b5QKlO7k6xO1TsXBhBXZtk9L633oGmifo
tVDzQxIKJNr8oZ+chTBz44mBT107jhosNmlfnK5BQsg1jRSQehD0zd9cLRjHL0K+
jtYXmP0FiXv0vNak/4tNfIVPt7lI/Ujl+2gOMbIap6R5jDi8Ds43gGEVsKmKy20h
Ar6UXqJ5HaqOrSG4wyvpC0nTgDHJCMTGroOfsLFZmXytmK9q9rZ4FVn/PVX1u6ve
vcuhJza4BVIykPQSiLSLeIF85b2P8i+4LD74Y7WsLZjygC2BMutx9e/FjqqdwObe
BBj/as+VCvcadRpqsAo0uiH1dSN+9D95r+DQ2IDxBExd7mnTpgIWeFhX/yy37QGk
IadC4HpkieubsxtInc4buLHhkhHZypDo6IX3SxssDA5oUNjTjp3G6BWaez0LPKPE
QYF3DKHxZvStKV6F7lTy28jp5nanxMCA2VeRyRD5/sLuMb+m+cKE7ug/foXt8Zwr
`protect END_PROTECTED
