`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/2I/vXZIR8kyKPCqO6hJHG8q+8Ps1ewsF6aQQfoKSGo8agEkaQwVPjVpaOqdjzt0
ShuEzy2mkcRtq8fAXTkCxS9wrwdaG/KES6YnzfJaALdd1CKLE4Fu/h+BYTDQ1cG6
q/WMsR1ts83Q14TLzdh9SytbM6xWbIQLuLYiLh2pVy5t9ut4T+yKJ/78GACLvtpa
x9TOJqEo01JhNNFbLjlJTaDliAoQmDXsoFZ4n9nMsWOelD2rnG5d2kIXi3GHylFO
iHl+SjryPiswJoKtD0QuTyNwQrN300wNmnCOuym/jw56mvIKUdbDeMerczPODsM7
l98QrrvgHS+k9M7gXtl2tUlNdhjJqSVHVT0+vNvoiIhSuPqPwyW9DiitSoXyxPZq
3ABGsjFSGVrCGLkc/3yKQ4h2zIn9PsOPqoUjYTISjLIYCMoaAlT1XJ55hCdPw3lR
jOCsZtwzHY8dJDHLj9cLeXXeq37zpOWlrMuwILQwHfQJJMibt43RPkAdJwLMLnp+
TNwFJyn8Tf221iZsE4PcYepWH8GKGTJ6nqWMpa0uDtfAzklKH8K0VAZtP5jVgn3e
tYEBQCK2pmHYhEu9ThQFoTjhNmTz6qX/0siRxeF7a0JNHmvOqB1FxdULPa4B6125
HxzSOwBFBAvok2haftyTYiitqYI+H9stVLgqOVZIXiuyUlgEafS2Ib/G4TUSqzNu
GOJxmWCFGZdT+ORWnbsuO22P643Fnd/jprY90Z/UndSYpXU2vw+K7IwntYLy5B5c
n5HJYoNUMQtA5366kzPzC/dbttMKY97PRweMkFDZTkMCJmVRL8jZUaAwpR7/bu7E
hAxYmboLeXGzbYYJIB2sJRmZgu59/YG6WCrFMq9GkeK4nX/txUefQ+wVmrHq4TDV
xMdizih8rvvz7TXv/7+TPr+9OKkbp6sAtPArlg+JtVWcNUK6rpW2EHEvBUnb0yJk
J0h7BcdCLLoucAbj6RCKRLhKGdAnDYa7ziCJJq5vsn3/aXi87QfmzZIXq28cFx41
`protect END_PROTECTED
