`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WMlN1h0nob+8wxfRWkeSQ/K+owFibRllDt5YDRE1Mqy2BIxxjGHVY3XfvkA2deIf
jd7/8Ug5nZDxfF7x+2ke1ShEGh+vJIni8qnXdGULly+TQm7yowuCvqHBst1gEOFK
sR0LmidW1Ivkrx2JGKZz+OkeXZTjFSJLfV5ptEt2CCZu1bDpwEBcDlEzPoVfqz+d
MWijor5hJbI7WW1AGHZ+S3QJ1GmAKrj01Rdk4n23iTenKSojivYUbZWV+4gctOd8
51llw7Vbat2Tv8WFwh4McqXAKPwKb3+z7fGybTUspXnFljWZCPTC3tyDXecfUqKT
duVVWOYGve9TF3HLj9CssVqDXw/3aeofdcWNLkSYf7+x+L6vu8PzR52LxFLHK0L2
VGrRdh0kkdA+x6t/pEJhphyEadXdnfoI+J8L+G5gzdLrr6WoHKmnPDxwmhdAN/ir
uS8Pn9TKnmtwilpJJTYtgvzq9vKVqjrPFabGUum8HcprG5M91EbPpnGnUxKsghGu
xSVVbmoRFGr6K00iUMtD4IK3gOtKR8buOyJz3KGT9Wd1DOm0J9CV8kdRaCNS4EGy
1ThUqsFwOQn00ohgACVQdf/SqWV8eWuHAOB1CkO0GOlm1kcCq8fvigpB/ynW+F89
jAJZCnTA6Qh4ipDcrWucf9urgHDMhv5cQsycE9ujWrToahho4Y900wPwyOWK8m13
w4NxaqZHRSdxFQDfJl4g2zC4Rxspc0uCIRJhBTYllGM=
`protect END_PROTECTED
