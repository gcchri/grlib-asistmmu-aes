`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xi+9A9AAWLLCJWs6yX/QtTqt6zYLz1fM/ZXfRc69+oPf+BEkoZJ47AEKpd1lgwGw
pWXOGrY4agi46eKQqbEZqmRpZsq0WjzC+SJ6p2QZY4jVppo6CxY/7xFxG5QP1HNs
M9pgucvnGB4qys7I5hkMTAblpjMbtDLKKasxWh3IiIRr0SbLHECX1YiyetXeEsMS
TiEvhaRPdJgmET0qRw7ufcGtB51yrBnnkCl+TdK+GUMj4jInLI9CzBkBAVclV0f5
LhXLjza2jb9+1A4vBpdmwruNN0gF4Bo5pxYoVKrOXs4fT4YNDQwFV3/C6o0Cx8DY
4KMqj0ueMDmsHQvWnaZqP/++wNqVOpeuXLlg5DMjGuNiRhS/qXPJI66RfbRN7P1x
Q5i/BcDXj0qBkQVGyusRM/mPb5sE6CKC9j1haaAZUtlTGSau3O1v3Z+zjo8BCaCu
Fy4FWsTLjBKC/m9QS9U5Na1YpV18Jgsdkm7SEHcGgjVJdulfSTfn4CaYFPBqugAE
7VLSU7xg/ZWZ9EcLj8lqtNBMm4KCNNKNdiOs43qxb4Ep+cwWBX0z3nb3syJjSgls
6/68nFV9jbs4+rxYajXiULpYzOaFPZyg/QZpm17RVvKKNJ44oeOPXulubZBVZFcT
Skz2Ce2qkTw2K68mL+/9Bjm+6K4aJv4IlU44n8mlkJ0LCoNDc1Is4n58KNr8wVyO
iP2E2ZWBvI5iFxUaHH9gRH3k7FHgBZpSRAH3vYU7GvuZ5I1KbvBvKNqjcHxkshpR
MzkfYvbVLszOtK9ehbj6MmeLfGTSUTfTqCxLjoaYoGbrYrmi+q3WlZ3sBLs32cPV
bLGPdsRV9xCp+OUwbfSmvvEjWUM0jjKf1HCi9A6VBFm959pxUljdDwdG2BzmExys
TzwRebLO9rO7CEj8u2kTIw==
`protect END_PROTECTED
