`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EV1YlTo8+U9/PIO4yXAy3k3KmYSK0Kun3MTR5nzxVb/0tUfzl16IB3I6V777afFZ
KqUxKO9hb65FarCVas2qFyLGlURIyGFZXeIv+yU8qOuUpb0It3CG132xXjB3tqf7
mGXrImk6O5w192YL5yd65sva+5MCD1lRyOVil4wX6lwVaB/1qRDjIHphDh1OkqjB
r7vcsPegDbKiK8S2Ez6Of94VjkFrEuZLS04J084tLO9j0thcOMtzNMxoUwiAkEnj
GSaar0f240A08lq9QcPbjExv9IBFEWtSK5WmrhLCItJR6kRtmzRCGp7FnYb2sSGm
dpKcAirb/N2msr/3yIPw+A==
`protect END_PROTECTED
