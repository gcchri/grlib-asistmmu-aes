`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eWNqhu0TlpvnHMzWmyXGcNacFj8dVfNvqtnp/E+5iAmu8uRi/O2Pf+iOoFW9Swpq
TF45NEwRLG2znNSwJbVJjqDgljG3npGqvqTW8mHWex/C7sO1DVmT2bznnjU9tMqk
A9hDSyg9KU8yCBagX2/o4PkJYSqQmfl4a9u/LDVvqk5HXlrpBa0mUulyQe92Rrer
CqTYjjfSt5O+XkbdrMIc3gEQ0oacaWh+bEmSuCxxAYRjCUvIYZR5bz5BT9kiUlRi
55inBn8uF9r4eVa8QEvCZoXB5oBvwKJLBsaytsWgWAaaFPGBl1L7rnTsAcWO2MU9
nbIPOC2moTHvNmEg9B3jVdBLT42qV7lTSKuiCajD0l6snUpVUJEDtQhS3jr9NFqk
+iA4BzWZ8T/ElJj24bzaa6BhZB4ZZqOD7BeXtO7pD8GhHL/yl9jKD3vHC3Kc0DCw
xnUHd3KcgTT0sHH3MrpWoGG5ygongPEdCBDP9uNJ+d5HX56mx8JdVzpXkwcTisuG
aBiHzSp7m7xtxHXHe67l5mjzypI/ixYCO6w2fGlmFQqcTzWWHqq5O7FoJIA+oRzl
j6otFWW+3R0ysQKHbcp4RTPBI8yzTjZvliiYni0GZq7ZZ/m54Dymrxq+IR62dyyB
fCWnMvcpi+Y54VwP2auL0oXVQ3UR6QHdePawZG+/T/2BMJ4dJi/7T75Mhwudus8m
7ckxyibCa0oScYT5B3Sb0TSvu9omJnpPky/1aDqCK1SHe6wdxVKzt41pQZU0aG4O
BTOsTxW1mDQ7iOfUEy1AtDwefw4kvdgxTUErUwXjE3MNYlxf7KLT3hT0KYYzKb1U
KCmLbVzfnNtEcaVqCHXjXg4huq4iIcM2vFGCUtpjNTxSKRGFGLx2eeBDzOQDkGnM
7Ou2WScIe6uvIr5xOBDg+c/vxdARokRPER+snK5N6mt1Q/7tyZaP4Wpr6f8ku26E
Qm+eImExhBPrjeNpc4suu2ubJkMK7F/X+59bWnMVE2LBQrJDIOw/Egfyb6rHK8H6
AFobkVeG+YY80JSfHLy1PAvGm8W9MYvmt7H0i8tLQLj+fl07yoChQp78yqC6VvdD
0qXM8l2+K6PVD/FfHfhAV8RJM3iODRHvnNSB08qFScOTbzk+3nTpM0+r1gWqAY+v
VTq7n64sWGRsVixfgftN8kf1vxrDOjk/RW+dBMF/HWNe3/53q52f/eYhG/93U0Yk
QB0ukKYyiJxcFAkqiUHEqbXAz3+Do4qe3nGRwaTu5HnHvImAX/odY866Vwqu4Thf
Es7Xq/UwYc1bL9trDKtmgJ0XS6HCRVncQkLkuTqrFc02aIdt0L6OhR+diui5tQ3X
kzPlrCBuYZL6QvU6JsiqFsA3Lb385eHDqlFdGWY3zdbsklccmcRkzmapv1qvZ0u0
kSaNE2L+vXUjIyW61dO8jANWNMNWpAEkuZsI0MuwUiQ=
`protect END_PROTECTED
