`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7WUT59vih2jaWu6r8tNvvh2zLM3EhH/E1WWRVdGhrq0hUXeSDZycFQZsgMFwi8Nk
oIRhPLjgszgcEWWGyh1nMvDjgqjwTF+8rZxDUS3ndHThww/19C+63P9RZ+TAD9z5
2i3ZL5v6L6prF9VNYTT+Sap49WbmOiWg1Dzly94+4U0cFuXUJ2vZ4XZ+NuX7IVPK
dcmE16WS8/cqkFgPmO3qae4xutPo+iTnj7bwARdXmLejFxuPfcOtANoGim5RtSIX
D03oirRjIoTeeQzikkB896eEsW/YwnQYZmwU+shKEL3XEH5fBIn9GCsoAiD2SUVc
+vKOc7yPe5MOxCse/ZVhaubeAjeoV7vKvmeBwa9np9H21ICBvF+IJAYMsShXfms4
8fa09nxRcjcXWSOPu2pPQu1uYZiaOizDdLK3NIFa8PE1/K9ePre1rh5QZzq/A8H/
W0lQLwP9xAb1Desw0BvAnFLf01pM2StUY475ToRB4acKbIZg+JyR/taBmBX8RR2i
CzIy+tpGRhU/zV5wGiz8p/TQt7blultiBdlKKcGX/eCyqhEyV4rVW/J2dDRyyv4A
`protect END_PROTECTED
