`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AQDMZYo9d9qgoJBVGO06Di3tL1/QUYdpH4sHex8TtCXfBno1DIQAhcQWnbinif4U
N8DGan+J/RNfW67VDaD2b4d0gL7xZSAXVe4unBOYbRdteex3BbOqsgddh0FeSlZr
KcZSQWrOmaEi8tzJjPsTiVPxuBcETpJLkIpLE+FAhGSYp1L4LYDwR41CSiddX6m4
UDwV+yHb4a3i0d5iAaF3mLzPRqP8jNmBVRPU8BtaL7oqW//Zn4IfAVskH3rMts5b
PwKR+dq+8Yho79AZR6ISvL7Z5gQZvJSnPs9/TZar1o6W9uQY4F0VsaESLjhDA7ov
7ehsRUFzSKtzFuFK01ev4Zp/7q+BSY9T+oylFjEFFM1O0Dv6y7P1azyYE3ozjvwQ
r/yrsbki/gPpr9PzMzaayg==
`protect END_PROTECTED
