`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rDOe6QfaJ0FJ4VAnJTQ8d5NvJD1SsceevdPmWXLJiiGlCWPzSX6DDuGq0UUCFDX0
ZZrHTZ2KwRVbV7Y/kPnh7R12X8utKcLfIF1jk6Ib0UHt9XMTJwwHPsmBN4dD+TSP
T7LadlZ8qj+vT92NIxndSfUCuUdAuuaNYjrnLXZQKEtZ8AxFsKWNSGxR81Czy1Kj
53txmRREwNWjPeBO5bZzbM1TdrEHTgSny/P0cUtmnmBuMASPkLN/Vh3LKqnmajYS
c5HLfmfSbEVxBARXowrXd5TXevh9WjuW1CKYg/jFHLYQ8h3HZHhFxhDXvk/RBxkF
mLh04kmUVg+C8BOTemd4pNarhADwfxyTx4fDHyNkjfD+PebquMNrCO+txk64QsPn
GGus0uVn37OEefv/W9wgPfHYFLdgXcO1pe4lXJXXvAs=
`protect END_PROTECTED
