`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tbmmW9Z9bbe9dkosMA4F/IL0FkBYRJ/tJSrBoW/p2eBK3Y+lw2yZ7nnwiiLEzp7f
jETY23D3hCIbGSbrYqF0RHUw+cwDeIvwuc2EHteO2S0RtP4PD7GfeZS+cS+YFKb3
Y3Mip2aH0L4QtA99jHju1A17x2hM1i6iwh/skbw6abADPgJEprHey8KaSJOLQj7D
xZJ2eBurrZmNlnmxTcHjxD6HshLulaHFWWCkf7SqHSeWeyiGNEy08fUaC2eSYJBk
JTdxaWlt7NCbBXN+LGKX5F6vzIZQOoQ5FYFH0LQxYRdNnSbAP7KNdqgOK0+2FVu3
t3/WZiRT5ljv6rVzC12HVFJUs5Sa8JWn1F++xG+QXUP00zFPg/rcvgjn5h6xdfEO
`protect END_PROTECTED
