`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kgp+wSfY+4Mm/M2wbmElNdnOdYYB1Gnouew/US/+qjN/RahDx0K09GPAVoOIxIEh
km0PrUpDUOySQdmMIUqFuCDV5nHRykcOcPK3slDFDt7TNa69qau6CR4v8UfJC/pR
xOf2KmqGRP578c6RrHnRf2wWCl1LeKTNQ+6zJW5aJIGST6xqcCFbbDB9VhkQWFVQ
FWidNmuzdrPtXK8nUjKOXL/CVlkCz1KDhx8zcQgXP/o5Yf01I7kh/fYzUBj9GIIe
TDWIw1XzSzsxF615mBXJmDv+52BKjUI9UO+Zgal+RMHX/1WJW4GjzIyZEKpWg3Vs
GCheyqqdc8zIkw+zYcYe+Q==
`protect END_PROTECTED
