`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7QLOJ0cNYlbBSVe2cwbTIfa0AsTHNIBqqs2pMMni+wNj4CqPep8qK8n9dhYeW33b
W8s9spgnIyWWgvOTKa2pe6GxcrPTbglr68yEUHfyvuRtQb5wvaBHg9sl1J+cnGoc
/1KeUIdat5oE3lL3k+yYSw6Bg2Evd2+ATuznU7P2RE+jZlZclsa7hrh0Ma1NygIx
NJpYLPkofI7PpcwdMoZMw+IaNd3zIQ5DMOFUugDZsbpwbef/C2QAMafXtYbEnohN
qJxcmFdytCLf5N1+ZTaPQQD8WBLo67ivl/eonMe3nByT4B3QXiXoqv+ZHHLYJTNF
35U8WOtzTb3JilkYfpamqsMmb0Umq9aSSR2kegMW36HNsxba2mTF/P/nJypSeC0r
oataVLPq/mJSnvaHvPR/Vg==
`protect END_PROTECTED
