`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mkLg/vZLk/VxwmbFa/7KCVzRiMEHKRY+LUdkKGb+gjCSSz+yDE6NoetKeSo8AIwF
AJ8Pgrq2JdHFbLCdJ3PAgvE03fTKBO/Ov3ypp+d/+DVlM2D1TfEpUkTQlZUig4ZB
Kg6GKU9AtJVEbHScmy5L35+U5MVcd7BHnQNCBMl63PiLZRGwXrMU1t7BDWBNwSLM
lZGO61b0K+13fCKzmFHvz9YgG701xw7fJP1z3hlges7O7+K4Y2Um/ucafX1Da4yN
KYiCUyUuKP+dysx7At65DnCU9tov4JjTrQnSjgig89M+ilwQf6yGUqC2m1sNxWkE
XEccAYjIKjZoYeXkzh3oWDzCnN1b/pUdYvRIGymrVG1ApoAC92sz++re98mFV+5F
fanOzbC8v5LHnGr867GAOJffKjNUp6IrI8dqWNcAowVGfiz59xNPYQHfI8f2kb7N
e12A/cJwdowoa91gdJEPx6NsQ5xoRiPDASTPr9AhXew3RWdi6zK+a3vw6zFC+bMR
Nh5BTRkG33xWTuYaTJXg5UH14P8XRDahDLUvW2ZOwv6zGs8NTz3vLRTQl7P00scU
/WO6EgvLtgOozdMuTNF0haC5ry7JKVx9FU8nCCkBIpwyQKTJiGBinV6vOXunBFdu
VC9jHCYRlDeI7rf1npHb0XlG7oHhE7jbEuI1QY4L1ezeqOeK8+4A4K9xXsdNyymF
vY6B5q1MZtJtS+zoEBOSQD5rbTfBf6TTJK+a9E/NxVSCGUOyb9PlH3T26qJRQVq2
pWJeA4kTgWk9QHAvv9aWmFpQWMa5kAhZeiZ0JdQgg2S5uf0K1J18AzjoEnujDEj/
NjabZ+yJnQMoq103Ye520fvZvtvG9vWehQSsGYn8IocUvNa9hD4S3w5EN0L9GzYs
JZtS44irRQdLuq8eurak2B13rXhg4SQ1LIMwPTqZhubYCcC7Npekr4OB3YU5hQtQ
8v+nwDcvCRLlbp7mna8Hj1RS4DNAWevM5z8sCXC9qUd7+gWoJShsdXwsIczVf/XF
kxTI2zy1ZlXgNy67YWBW7fiwceXNohcjeVmwV4XcOX18GdL7IbA8qNOoxJr3jPKu
jtlZwC9W4KxjfpWbCDY0GF3SyfmtnNH+4Doarie6nUqdHEVfcO42yjgTJfDUWkhS
FJKdkbz11WIal1BvwqkcuyegCZkvx3Hiw51Lh8+xILfZEHO0kauuB2a0fNI1wJzO
f2sUIlqIqggeEH5DrP6PmnkBtQH8ImEt3o3awezfU959POuUaVbwXEr/P31q+4RG
psk9sYAjjvkWSAjay4w6DU4L2ffXfMgltAnrpoopNopg98LCosjRs0pAC/pmlUV3
5BvbTGwNidPZCabINNzVUwAPYuvWqVttz5yjRfSBi3EwZ8cCPt5h/Ia7U/nzxe3T
1v0aDCPYKbZlVSfRIitKjkNQJERqXHUUKOH2v5MwI3w+sWB77ytNhHhEEdZpFpN8
NbwHt7fx7CFhT1kyxkSKbRgOtx4xVeUYyiH39mPX+bI+yo9Ulip3zP69w4GrHlJp
I9BMlrC846/c8yRXlYJYg/4dgS2TZV1oxzyZJHt8s7f058apwFRKWHRhx25bfyzC
gnR7qNNyyCIM1lWX8PEnklGWlnufrdOTo8PQ+xEaMh0m/PS/zH4Wo5v9Vf+xuttY
7oE3NgGMR4WC4ua8yyGh4bz2FVRmOR9ehv56ZaktWGDq9WngzCmWYDmnKbVkPbNX
v+kjtvWinQm4QI20wNR7yE/9Uhu4U1H6ETmYzG2G4j7JXrO+FjIDCbcro+3WWw9i
XXadbxieFoin9NtKWhs/Sqh5Wbs3t0w4b8sQXziRLEk1RkboTqzSbC6mMZ//wq7V
AtTEkOvDvZ8f6kekdFuRHYJ+T9LfH9+kycgAqw4MP5ZkGjufIz6zPntULSPFli4P
gyRMexaceM0Ga8l611BX8Vj2pjAolt36emu6//780+uxOru3+Xt1f/EFRomQ8nK3
SfgRMmWA8zYy9noJ7sHchNz1S73GEDH80pcDflq+/h7i9o5LCIMuCO2ggFsSkThM
lvdpBRssbOfAN11deb9c0Qk4Racz3RFENYxoijYcdqcaScl7rfKArvHaGocEQXt0
Xi4/qBsacSXR+KSw7/o9PJ/64+PbA1lF0nbPTU+nE5kwsQaIZZxU0Uw9KI8PVKHq
BRzEwX32UJ8PV0qTg9mGrLLpdvnFVPAV5/cHrOUHuGw1Qjqhf1BvtOO06p3VAP4R
fiWdgpr3J9sBRk7sIfc14Ai4LM5d1HfQWAuTBsQ7lma+KJaks3RcIo0nBxQih+rL
kFAQK8HIJmdhogWg4u/P7gDA9irpnlUwjAR1P0H9OybSmPvZgyjlAsvi0yuVkXZm
UVv3QepfrdaWrv1Cl78SCVJfgKlaIPc6XS50nW2T/bKeKCH/8/koi90gNUilz+xy
y3CYjXvAHzED4dY8TKmcLqZWRMC1RbeQcRkhsYAtV4Kw/bqBYd9eVljIAUvk/o08
NNKE76l25QkKohDLwl9mQh5KSWkRAEpeRre73A8vClfzNudejRuPphOaP1KvsQyh
oQBr7UJiI4QzwAHNQj1U+q2QggGUr6Kn7UQa4EVLztP/9kMmKuC3/UZrA7iNlTXz
aFH9F33sQCw124ec3Yq3KY16nyAzdR7HdiISzpoYl1PJaPMDOM1rjDumuPaWVH7B
vJ6IXE30mUBTQJobrcOFmzqloDkNTFggLQHyJuI8U8dkMzzpRVoZRlCrYMfcsBZw
9F/TcCXphUmSTdxnz17F4WtB3V+JCZB8ok8JBphN2o+StUKqV3i8Xzrb1oqA070x
AD0PPbLLpZ6wqFVAQx/ABPdeqpaVV7yqTCuhA/nXCBr1zsFGyIirURcf6myKWi+A
S4Y8UoeOw3/vGHMyIZg91nmy5mqaUolWfs5jQLsb246Pu2e7eZH72GnSNT8NEiRT
nEFKoEfF5HkbabBCFQEmE28NG6stBv8NB1h3hCfLSQUo5tkQRbCHfXS7M7v3K8am
rcx7zd72IIYv4jCqegBDryRXFQIPGhUyu4K8HWrtaTkVb6sjR14jY01A/EVdGvVJ
05EaN1za6SlFd6PVIoMDP86kwMKg6jiDVZ2DSuJdnttqmUvUsSQiTXba9J7g4R7p
kcfRpl4jWLHXQQN0K3e2IsFhYvkf9aKaimughzYu6fZ/YxpxVzTaSdaRG8RxBC/r
uhHGUWmws1br0FavIm5q9i+6zYEF1smsut847SMkwTD/VlbhseIQUlfQ8v0Rfnif
VkMuI8fqryaEasvL+YmHXu9c0JfyL8u8Gzwu0n/btqy76ECxN4zUS6ReYXhaEe1l
h5h1ertwnapfHxCymMqdqLItYk5AUP0/VfaLwCwlfDXWCLDQNEFVHlOdCyGi38z0
0qPNV0Hwm0n73IhQSwBIETPNfoZPJ7+r4BaMU9ekiHdYOIvVUItYUZuwGItV1ZtB
FPXVjS4FpM2NPQZ786mCv/T3lZUZyJ6t2UvVA3qojjLkDpS6bRZeBQYKfJHMxejr
dNB9VC8xLBUNBljN/XABk3ulilt1m6EUW1UW83fvqPWQjv9Q0yFy18Kq9gp6QlVd
WVskd80xnzqv5+4fHRUjtLsarPRRTcgtMJsNs96w4XHjQq+WAH+/bq0OO/iP4Ig1
PwGQQjnOBVY1OAKoMD2GsN67mZqgFW4xBmGscqDNb7Ux68ZEOy8ThOH+gtazY6XO
EWCRVxVyOYFVxMMn6tlqdJKdPDXFKtGtVS7MdWl7oNuAzFc6vtrQDddytDZhHQzg
EFO8EP8RMGzl5dmQ/mCbBbJWeHuRpxQkYX4qiK2kDk8GOJ3bBKjv0MuMLFG5h+/X
4i/ykZLaxzObMt49o08LhTB4B/6F4MlgbkSZcp2q64RGrVXfYdMV4hIbi65CIrzd
LTFyuQz2ztl4CQEhbNo8grUGoVSLgIP7DrFgH03lOGZNIaiiBopTvcR0KeLmaOCo
5X8zGps52RtYgNPDI/Tk91K8KB+nRSgJWQn4nOLibS9XTxSWS0skOiIDizr4Tyt3
i8GsmpReWCv2bpzAXdK7+e9dCLxTj1m3OWHOb88QtvSKqrXl7LQf+xfGmjHtlJ0f
xjfjOCHatXYZbrKt5/BN/9tTNpZPABOk02gfdDXyXQdU7iJoJokxPXu7m/DF4EZc
Dw9bfM34TSU6kleTvxuV1ZoSOYfgjiRVAHTAzzlNQdfLJf1Oxiaf+ADzWg67d6Sy
un0g91fIMJbW4eRbOwGfllxVHQsAhqFFlumTBAH47ClwIbUF0swdz1281oobARBU
DxUddLEG1hudeI3g8CMoYA+6/8P98RS2bY69gbjv52fMsbVftkarwaR1Yaz0U0ej
OaRvIEpHaKXUFnmbVjh0aUu+C24ONC7iPzbPzluKbi1U8N2be9/bJJZYX018MjFh
OucrS66P9jnvsgDJU9qRYVdqwucCs5gG4kDFZlDfkDRUI8zpaxPk5RR4X506pWa2
kuSr433c9cOGPzE09CwAu8k3XUmqrgwKP1mA6jnT3hrR7TjLT6TOnVgXTxvRLb7r
CqNUq9E6inRQxH6jqwMRD+O/aXMoauTuBfFOf+pbksW21SatSevG5V82GFAw0DB1
VHJlJk3vYDkhrBLcryeFTYACb0nAumK49zY7GHSA2sOLKkUkYBR8YEHxSa7KotdL
rfwK4Ag0ZfozQ+vQxk7KAsK2opIRyvfFiT7+saZetElU8lgGRmgSNEA2bEbMhQKT
wk4AjhYKsjSbjglek2k0B8D1g5sAwyFcTPyUA8IxkhEpxYsE51GcYxMZtrXRQT3g
I4zh9Huf6JLdNp4mwh3ApqQKWsLYcOadLTGwE3LnCXu2y/WYqanZ/KWUnn2Waa0W
Np8kZqfhSTDQvsvitcjD1uRy5WLU/LvpRPl47jGBrjuKi12cOvWofd0aZrM+ZTmH
lAIEVvW8toe6tg4QxXu98VfrZhtmwcX3vFSF16mzldT8pVP3H6ygflkuRHMuz4/P
wLPsOIitC+ax8nDtqnJGWStG430R1SIHXzDSwSQ3EK2O0uLyxHjXrSJRVRziMgMV
d8RoCRosUQVG7VaIpytXkwxVPVK9JJqCEkWyAwXJpySYs9Tu5unWWsxoDuKxA+cD
1XBRZI0DQ9waaMZI3riHeDCkZuB3Lk7qfXC3OF9FUzt3DAK9leSxDl2gPH2YxfRO
39pS4e9bQupk9o07wP7QiLtFxSoySaKgOJAtv1UiLp37Hr3Cp8Rb1NreOxBBbX1T
BF/kUIaZ84tgfFF9xi7d90E9XVRZjW9p+YHrK8n7uyxsbXuvSf3xtP/rIFBDgzwt
eToMLkZLt0zNfqk/kWTKfxfOhVJBGlGPj+S9ja4KP+2BRv2KTeXueDcchH+7jcwh
URZ+txz19nm75hyWLgFtP6B4xzTjptXs6WsCQqLb1BhzubCQHhjtZrUh58NyUzj0
B29L1uAwtLoqSKjoeGG0Ojm/rwhV4IgytcFy5x2Y7l+BTSY3gccdaxBUOZ7hT1Bg
M0J2DXBc2zu4LqovuLzmtFNu+9HoBHdtiDhs6oVRfUL54jHh+TPQ2P2LZSeiutjv
ZAAfq7CKmeE3vjliHHAvRVUuiWB+t4MByoiIMX4vsQ19Tm718RdYejyDqbwAVfnP
xsffr+1LeQZT4eEurcpLmZMTTflsBjce7FcR7Pl7fHm86toPw62aZsx45eGuTXib
OL4wt5PG1EF5Q1O8v1Q9yJmxdb+oVE8OjnpQqOrDz3qTSUlHNtYGJ8uN8oYoi1S1
u+ieJkggkDjvkgRFNXBJOyExUf5a3kXDlv2u2PTKcP99qOA+1LVLagQXNvvelgic
0fDMvGOElo27q/ClGYy34JtEEjBk/4Zrea1x+k36tXOcF65y1wVtyb5byDjmfe6s
6aXXKGwAV4X7FvDJq2K4v8zHiDYi7i+Iz3NsMfOZBnazfQTGmaYjaf4VUkRNexd/
Nb0ro1VUiwUIMIxNwE/oMP2yT7WJOoY+D9GNgn7VQp2n+5h0GdXeoFVCD/Pis/4T
0TbVeX8Xtm4mZGNiEFX9mDAWHrLEqVvi3i55vQJyxWwAH8lY+5E1Q8I73hGLyoCQ
0Ctimi1sMQDLkvhXkoVuSAWiRvTdNq6ayXi2t9Er5Wbgb/D9fsNlk3ExIXxrm9x5
ShK6U6pa/2PmVQzoYwQv2DKaFEct2Gu4BceHhfxPfxwliHZd5MwQ8Q6zvQj69cbp
33/NOzFsSnZiHxTDelM/sUCJd987AGfbAGQUqLD4sZTjyn3WamzAvwvn5Ob+MYo1
7NWe3/CIEAofISdJ6tsb7XoxulhT8quebM7zMg744ArOmd1Qvq+mv21CMm1a1HYc
31/ERhxH3MtLy+ol7HtKo/UF6nGqYJRObXWYKbTVb+91s2cwgfX7OrP1JEXKDo2W
8BSsF8Wt7Fkic+Rq5sF7ABqufrOpFuSRsmBLKSudQP6fqsmhJP+wuiEGooMrS/5x
F1yxO+nesTXP7aBRfnRfkqyYpjJ0xQ5/qEafzIACKSnbrWfjs79VF3ujvMsjpV9F
dtiDxAef/zosQQTl4U2x+0THwYydt3ZqfFHbUnL23oWMDyE5Sx3CawVoJXiRl1j0
kt8E6i+8G9bQ27H3cnOtH7C/ulvckpAcynwjOn+p2wTKD7CE1h0dTKo+/8iQfg++
ORa4tbBl/Av2ghnD7b7dAmB63hHewSIjb1lPi+NvKgywF4I7JmDRTKyjwD6pfhLt
sTGKfkEQyYzjsclO/YX2zm2ZKrXU1dCatcOUUGEu6S6d0/E51m3As738rH2Ow5KR
ZVLu/WaSjQ/+1unoMTCkoLtrbqvWsBJrsDayl9jLBAj6WdmQtfw6BwF2ozIeKBsV
/UH1uw/5VJSPLFBZVejaXz4CxhfQRLKO/Gdy/UHwmMwhIUqkD6Lg8/M4awUfUwzo
tDgMbBaje6duwKvXJTxv2M/ad5OErmm33s10ufc8cDnlqa1iFF6HEVZuwBsNYG2x
fUcHwocMGpne/64/zSy+Fn+AC06Ud/n5JpBc843ARwCEe9CkmT9E0ha8AlfQToyq
bebzdyyaQES78XutgOtnKs3z8V87aBirz87CVRL6phcRM/EzE2wSn+4XtOB0QP7l
unJS+sdJFIB5kMAlLXwOKF4kGREBvJ5H/vAUquXqk7GODYhR+u2YRhm6HqTr8p1o
G8EKKpr7g/Lfx0vmprJke8RL2nEUakjMchLo+P9dYSjmaCuUz4u8bwsr+Tz/mB6X
RquqwKhE4+qOs2IKaCt1RJNeJsBy24w0qLUtqZ4QCvnOdmYfHLwTpK4XeBXKimJL
eLeXZxMYD08TQglmpnlkZDCH4oMJloDr1+g0lKwppBtWp3WoR5q/W+Ie/biTU24J
3CJ28bCSCA1yetTIOXwhf+RYKR0tGLI8aPH34241CKx2U1ZVXut4oeV6ID/387ZX
GBZ1mjKSrJ/t6pE6qSkXci9DW98mw5A2wziIZ+LTbratbJR8cOmJwivwhB1Uz5lT
K3Doz2iiKhrusnH2H5yNPacWseXhXPWJZ4KVtyovDFTNPRmMmjefQ9WUBps8JqKl
cVUBgSw9NyxkgQd1o6c7vb5303TKgRwtjZgeCKE6fCzZh9S9gTHVYiyqx8Qfnlzx
ge7+E0DLLMxe3u3N/OsCSt6wvoHujZGNWg57Q1gEpT6tbmf3E/jyN6qbbDlC5htU
ptRPTZdmXttc/tNd2W8jZ7nc2tkXqgafsMq5CHt5GEdyUgnMc5bwxrpgBm6peRAf
kroyA1VKtytIpcnsGZ6uhcDQhRA1/A0G5sXi6hiT6m8/jml63qgnleov0LhaHl4b
EnLQ7jr7USNz7UFCkkVWIEvPZvNAXejMX+L7q65RbYXesTKAYXfjiyeuEMhxBUlb
0jbCq1/6PfWycfKEMvcjHrVfjUUFsA9j6/E6FuIBTc67T4bqn3iFa041ssuRpqpi
dYaaU4RzFLLcJxleQLwA/Rv6K3RmSN29ybNg0wK3KAjbyfUoPd3Ivq03FAtHH7hD
YCy+yE+3fqJhhBFGKBnhZBv3fhadodIAqVeBk514+XEZIUi5amIgHvbnag30rdvF
62L+1SMtKXm46fw0ybi86N2MV0AOBfKTFsF2K4AAaVvX9GPXggkgos6rsEQbBm4q
7vPv7KMwRgEP8Zq4lus0/3CNqV73g5aaukisk+tSJxrGq/IK/QDCrHM4hKmkdjnG
BVQiao7XgAXrDHv89M0ClLvExtHGihHb5pUP4coXXlLoiRurxh24hkS0IFlwroGH
9KC0pDY/3/DxP7Zt17uoevNT1SXBWVe6AUjips80wvdvd98ZsZHsVm36W8dyy4SB
eVWEhsLvhkYcFMbp2UJ7+Kts//H7W5g880B4txdcPjCIHjQaH4oN8gd5mXVajCpa
N0MSNO1mdgP4478WEkMnLeHzXa8nPzGU7+hgbGT5HhUywaxVxgnIoF1E/JdTtlO5
UJVoO/4jc7YJFbSoQUBlxwgfhOo+nwzoN9yrTbYnwDP7y2jOaCl5cEWoJdfHD5xb
M1PtKfGfl92TWUEg/cHtWGLLYe3GM78EAQMCfSLNSQJemZrf1IQYqv4YIzgCbm0e
AkNBno56Vvxgtq2GFhDHoWXrryP3kFgJJnqZ7bucB4geVmr53rMuAkfdhpDMa3W8
iycwjLywCJtv7DjoHJyxxGEZh6qw5cdpKPvsmd0d3vHhPI7SNKGGmO+Nv9AQbu7W
yaIcRJpL+SNP9jFl2pxkqqWLpYMIuSA3sK/z37vYOd+wufcfi9QLTA12GMaqRRwD
btYNS4iGJG7T6wfzi9VbHYLQTVOUclg4DaqXXx9feTy3RSLvZNP+EpumVfx8vL85
3hngnFHtgkDJ02oWqPxyEwsv6UuT8QsqlMuJr4mSXsbN/0KrhqiccXyDNYSXaPvb
xhr4nJFDzol2qLefqQuJMzm2Ao8biEpuwsXjIadSURfPCQuWpDzbNj/yJrMxXzFe
GQt0aUGumihRodvG+9mXKKq0LC3qakHjSPUUv/UcMpnxHE2HULijGxTHzUsLftOc
6y4cEDPIvERAAHn+LSW2blKuc38yC286dL0SPBe07ceNscwvDkzOSN95QeE77Y0x
rJiFGQHAd8mZj7MUlzVSeApUigJkTK5AgAnSV0r6keCsPD8CwpHI5FicDM5poVJy
wcf22SjoUo2VirAW8IlIQfGktzLDbnMe2fl/iChnNaNSBxOXhGiajlBnOpDGE7Ey
C7mq6SmToXbnZP5rH3SHhcoallFmUvZxHkneDIOPtICHegUDyZq0DZtx1Xf+O+se
Nt8DVGx7RN6yw1tnGwNL3oiP9sxgar/t2WfEhExlzxJZHhAERzXe43yKzs0DIxeQ
GoI8kkOMa2yzr33mte9UHe0daSBMHgVL1LxGZZag01buuwYzvlqiIpBkWCqyckvh
u/TWNCb1Tyn5VIYKCMNWfL5twAR1OuE4f4GSekk8HG1luqslI/KTs3ZKU77uRYr8
ME6u7ZebybVfAcJSryZTJrxwHOjy5kPvFsq9HTEVMOTaociZ41O0GozZm5+4oPIM
xv73vIEB4YqNOBDhCVr0Lvr6iDbqTRWWTNiqSFh+EIyb/J6XogzrL27eugBevfsM
iHvZ92e9ELu4vXE8fnZFIL9LdmNJBiyAkXF08d59elgibN7akRzkEBM3XOUVtUth
RzAaShfPHHznlhNMBC/6HOrcDS3WLEuBHKml3SfRkcQKQs0+6OZZWwKMyVfkTYWk
GFKH+aluj7wWRfePorEwdd6zW1UfMbLQswcT+5SJTGl6bMzjHjm4eRjMivJoHB7W
QQ35KjbRVh5YLEQ+qC9a9qShJP2pJgKM4ZC6A/qLvVF76wgLBH5rnmjDsrrQDvmt
I//lDfKN42+YKye3Sil0NbpceixrnEfvLltkfii8XNDa6lYlISPFnKJt+18St5IO
MoD1wvYBDC/ajECPWHHz0f/cOetDQsW6z0CF62ajLyvNnlO733DWYWYKQEuqe1l1
+9EItoBLcu11SLJN2E3nBJoNi8hdJsGWqzGzn6Za0JrJrIQCN0C5PzemeuwP+WOx
MbdA3OFzmXVRnyrASTunnycIjK4Qy1fAPu36y5M6wbWfzViU6o5JQy8NWTLmpZ2x
kJDSjg+bwl2kPTpW18miDaqQxSJzITtJK0q6yVzg5b/MgUhd501xECim59haUVpJ
EWOIdgpuvvBYv6uTsmvpVvYtvQ9UBirviooAcOeyH0mfXXR8OEob7IW4+n3zU9Lp
rDpuzmxWCtiQdyo1sdbuyiDcVh7Xa9RM9MwbFws2bUgMj0uCUfw47OWr0l/yv2T5
A8hTpjOKVeSY/j3YCOA3+o8BZh7DgJ8IgWAjrjQEGwl15ApnlrA5UmxT22chB039
0quO4sibOsnTRd8nQRpK08RdlxNF7HJmTsuyZ0qdkrQxORpU6eNSdD3HjiwUiPJd
Uu+zwcI9gmP8ZJTk8+qIsxnDrQcxpexuNZhXxohLrcvZPwnm6JGvSXEQ6mw+k1we
a054F6UjEVJtZjl1oZBbCrwzYPb0lUmsGbTEQOuBy4Y+5Y/rM0zVQEeYocN7a+8n
rl97e5K96bYeLhvdG1CjI4On1nq8AMRwWhJLgE3hG+PHM6/yGtS24ht9xAVsFEio
6AqwCmtwpG8SDXmIhMI1d3s92UbUzXSQUgLxQ5Thyo0b6I5i313+MrSQGoOXhFzM
NbEWrnUZGWw8ewZCeN6lAZmnr3pRBMLwWLaqK205L1k0vL+tGF6oQMUb3kVved6b
7VpoClnFKA51An/vlN4EeT8b1X0MLQSCH/UBqVXTWQd559IguKQBogkdZy5vA33P
BMUpZ56ioXV6l9jOdZBGzM75RXVNOtJ12rlVTjr7Ro1ILZGxNpJQ17YBfxWw1UT6
v/aF1HRM4UlHPcgYSUVYqTiwPZ9rMoTOiNsq9XwGXI/kpSL93OSlFxkXZwGrFL+v
w0zjf6ciY7/eBdSHLAsAXdyTOnVrGmJA/DwqjvU7drPlbqAD/L01szBU+qe/0LVE
8BXnxTmpLMSgEx9u2L0erFbd9Y0p1EK7K9eiJ8RZdg2tU5HH6iJpajCTRdzQDwjN
FEuPa8zljAsUfTn6NI2U1Yu+uRYHMaD/Bb0tFPj6tepul51ojUarLEb4yxMXh4Y0
aR4T88XWMPEeYM6hHo3/G/G0d9J54DTwgRJI5Amloc7BE9chuisi1Eggeo30l49Z
CdEreiEngpewsWFohToHZ3L+57Vnhm96PRTc+WpZ6hFxuPoAOAt29J/BPjlswlse
m3KIBJ7vTSgbyVSdDtn4/V3HsHwAa04lP9Tg/E0i6TtcUPOWOoamP6qy+IBnhfEF
UAHZXAc46BFxg9x/8oM3bTbeHRF/31WgpVjyOzqzNXnMSy58DEh69GNl8SGP0MJn
JpLV48kJ/xu/yRCqRs7cu3FjvOX5LWS/s0y6G781LhC4vLr9B3sHjz1f57iZt+yZ
5pq89W8AXo0CAF5LczOr5kXPorA5EaSx9Ciyz0oQEIXIl+vGqeFhVeaVPHGAnKHT
jTMoIQ2Sm6RE2LlCAN5WjN563ZHok89t7DIllhaM3tqjVgZ7PweKFsxmGpZtRPE4
xOAI2aJluYpkbjCYDm2jQpYmBKJnNiqdy9hQhTg1tkvSVmVHtaLY76j33XDIt85j
jX+0v8GC/UYfuJdeTALqhw4IMyCJOlVzMlyUZl9JRZeMAqfE6YtV3+LCtLAGhnn9
w73jCDDvjctjeYr/hhjYzpa3G0a40a0slZIiYZPTrAJ8TH+oASoDTOoRU0HNSsvX
5mMsGHdrZjlRMLfwKCjIUDhGE0/KjLV7GiaEpPg6MZBoRsKL5sEePtUpoV1dGxhE
j6yEXdzzXNA8EB1hxVJlp4LrpFDpIXdZNjudHR//UfXytJXA8C2PCq9TdhnjtseN
NZLiAtmS4JL5Apc88+KMwgOdsWcwJM6rd+oRdldS9tyDxTcWSP3Unyy1Hl/hm2wo
Y1rRGeAp/TYBTqZjLCiVCKSY7CMYeRxtIW7DhvKGo3wBwmcr9FltyLoRF1Axcu8S
vcdFlwRkVY2gzBzqwyk/gsUzeCDImvXgorZG8uFubGOvZb7DuQg6S9hhMFUU88Of
3FKmrDVRCs0uPLaIKk+tKE5Ps+/sBfZhlYH0zaAf8SidKHSNcq0hAW/Ii6kM0Ql1
Bw5RNlFmRtdxG0A8c6D06sCG7mad9so9T12ItxdOcMM3Cnxh8RL3CviaDAom+3jY
jCB+0SYnxDDArub/MVNGM2ZiYSZJgc/aocvyEEfBZFfMfv6WaNAxTlxF4jQHkv/K
SlglKM7KsaYmcfSnlLJG7+Scxs6k2HtISFuGrE0bPxViNIVN2r364c7sxN+1uVnr
T1Do4w4csGRv366TmG7o9zZ+mYBIg/+TBAv79lOMFVYErkjeAcO5l+FqRbHzjfRF
t+PynpNi02ry+50ZxASI7KK7C8TNH9BLrWOPB1tblOEOTSYBLSzOPdpu3PFGqpMC
XK0GSRqkPTuTchjAUvYRwifhQpUKe4ngAzG8ZOaG4NVlLcFPJFxcnMWBYxEvu+2P
0C6s4e/3e7TDsGTuJsFeIxR16kLWNCVPSQdkqZGaa//E/N+aA0istJBHbtAe+221
UMbldJ2l2Wu8Mn/ZnYFQjuYd58NUqShMKCT27Z1klulBDT/hulQwbPNjCzgBRSNK
t3cg0LwBJ16coHi8jsfFXm8FsWm1BxS9PqisjruSLFBpBcv18K5Pf4YwDDz0QTA2
N85ngI63k32UzFMKlAJ/PqN0dXrlfNhspgHMzmVrOoFO7DQ7WNEhvvsx/R1RLhQU
0y6ius7E/PEb7maPNZx2J/zIcYfo9qinPrNNEsz2qtV7lMsrSMqQpF+XFEvOqdx4
ahYBIcD5dmOPVH+ZmB0UbuPI8wt6KTKWZunF0blXTYCctjVvhEFB63zvaPSejfFO
WJSoqkKniFLMaBja9KC2EU8sdqjG+0sJXRI1OA6ajIZF1Tsb+eDdomBuGh9KKKw/
+B1eCWMu3qHqwpfDWKIGKGISVb7pZiwN95Wfq1MRlJ4KViElK1JJXecT+bnyu6Al
m3nofOlBRRF1/LBZaLVOBRWNWBMOoqMYPXQPCFTI+LhXM7pgATQ/hIsKIkAtMqxs
Udr94ni337MrLTIiHRqYjJ268AKAv6nxQiv1DmL23Ejqwcke7ln+jS+GEO2/DHmP
ZaP6RlQlyPc8BN3f21YWwd3jLmohU/YDePp7uTvtSwXbAiVeA1f6yoQ54lN9C7/N
KMD0GDd1EWRIwMl/BudaqMbfcbetDnYBxPMId7162dWNdJnc4w8Gzphj0VWRx3Pi
FO97ri2A+e6EUIgg+6TVUZBR0QKesz0Kvd4S4QXjSbdAhejrE1tXcaElAqvNLxqP
6eLPxqPba0oAi39xZOqAVnxFci+sZ7CLpsn5QcyT7S6BVSQaA9H0YN01nvGuhrEL
Wx+NIXKEWdO7YzYThBxvFvVeXzWuklw+o7xabz/jlBYUWnYMwitcfE5v5tvzKo1L
Ld6PU4jsfh23MX5pMnuUIQn6qt7/dU/plKynmnHmQoPLfrUc4ge0sYodnp4Yf69M
HFUeYs/pHYH4J8a62vdanGtuR6YXbzPCcAMLHTDf0aJjHdVdt9Hr5PSvZoWNKh75
Gj6xc4X21pXL1/KzZ3DuWeOhP4jw/DPQMIAYFleP75f2/PHc7c6WPmYkyKvvEhZu
eCiT/6oKKtWcwTGXreRpqBgJ7g57IzER4dQ/4JZBAfkDo+GSbZSjH0vKlw0DoKX4
e+LRH/qwYA7XNvwvwC52vQ0qNoEci6PrDOjeauIOJDViALTT4W0jEhmoz2Tt4LaS
qCsIuDjV3JYvOq/4SD+y6BTERrPSEvbuJdEUS23qHEznzzeHG4Xbauy4cnrTIITh
LW9Lc8sL4enmvYyUrSRk4tqd41YYtwkQaHMZS2nODEhpTHlo4pQriO137TZAZfYe
W524rnOK33vcL3FiqMcCLzNZsEJpFCKkMz/8nRX3I3x077n8vErTmgHiw0XNRk4/
NAdPXPHEhHS43v25UOVqcwS2KK8m+lPVQgPtQAq+14QBMT8hHCEvSWMhctnXQXxR
kuJbhc3dq08fT8c5kqkfVZtUPOriNk7woy71Sd52oqsx4Q0XxwGFSzQX8rlFQETy
T9xscoamOWEMNT1fMoZnw8W0MrBsAQZhvJVJVBjwq8PC3QA993UGCxj4ip9n+IvA
MaqM7wpNZqM9wl8phpRA7l4BpWZcTQ8w1klIVHANbuKj6627yJmtug0iwCwc5Rdv
MGHWksgK26Yu2Zr6lC/NLu3A/yGXBhOAAfBqLyCmjTL6l4aw68hYgKNOgPqYNDNk
p1WDP1fwlxKX8fdF1+I8mA788AQparrTyzF6RswWnaZdx8hMfCuZ5qiAcodXF1oE
uSR13uA4o5nHIWAyi1LKn0609LBUn9mXCl2J1st3f4w3wVdBY28EQf/aiO2KdfdB
9oY1mmhPQABKhr4atYVwrWvbkdp4ZlJrgGmnPQ8mmSCmx6tCxvme1XVWLFkAioSc
9DQdgrDkzxXxYi0kreIuat3T+sYe9ovHJSJ1rMoVDVjpzXiXc7nR9CLR8JroV75b
HB6o5CEykcmwFGQdKnjt6U9DkeMychc9kDGi1QQnwOaxcwPSPKxWjPVoGjIOWARl
k3mwjHstRKi7BlCKRrr/ThrDTsHnMBBRRDQncMHLWK/nztdfZGR2qpixnSEmdD1I
nESxXD9vFMuyZHZhCs8xqwGnmU9wTBxmrfX2goc9TdePAg5oVHtTEJ3NQzHEoVcU
L1MbOVhxXHSihnvOdQ+yfMSWwUk5lGHnPSno+JgVjsZG/fG9OPBISW35FZIxxsJu
Yw9Z8Ckm7wHdcCjQn0lJsNZ4esIKsIiILnwzt3sgUYDyFS/bgdmFl9PLcc1TY+9h
1wDFYBGmR3GzAY6W3wPgGLh7ZPq15RfXky4zumKmjCtlAm+8ARDKgIoJ2F4YtxKW
qeM203dPb4REi1gyIBRgp+g+YZ47Q+FGQvGbs8o1sNZxdQgTmUeOEGb4ka/eTIjO
ZlvExU2YaKp6S8uxEbteUUsh7+2syAn0JuezIcdR6JZGU/9VnNAFm4ZQCpsDvr11
ilgiHfG+g3cYxnFDG4m8ZWqSF3u7uCkqlfeMV82W9G+pcbCVM6l3aBiBovVnf7vH
0QTqYCT2hn4lo4jpbKv/xEuxd0czcg4CpsezwJaB60UOniRIeWSAYIr/Cq/AlR1x
EBZpnyx93p7eeJGHcmrAxcJmQf/DqJCQqA5+NbpHL8CVsEy94J3j/Zn/UulqH4vh
lmUC0ELXeVYIxntc14zmKa9LYzCvAou7dFfsnCcnYVTGfh87HHTTrXtZypin1Uhj
Od4HhwKVACx3YprufFj7+o90tVWA85IBRkXmIlDhSGZ4qgPoqpsBb6c0PmndEGI6
kyl1lJdzJUiheYj0mbSiQhswEZtiN7Qn2o1onnqIURq2OQvYaXzh/foXpVarE1NP
ZV6OqJaKIw7JHvJEyJbHP8H8LDueBsyvSTiTxxK/su+Epc8t2pJ3nfAzLMyOxBJ5
i+ceWtZZzByFjguJF8+aDe1cToxumCwPNAXtQIzurceRye9BmTcO7KUuVOwooSDM
AwJjq2XXKDhgrE9l3SYeAOlunO8Ker9wLkCGYif6HD23wh59tG8ijngVRv2xdirV
N7cZ3MNExA5CocqFZeQD5issvdI6euoNY38wYq2oYekN/ch6keB1BfPPpQFF5yk2
fcSfxN770i/jpfEIhWZ08Un2t5sVeQT27wU8xjnxS8bQWmUNZRRvS9ah/cF+SHp/
DBHEBrszofyk3kjgXlPBuwwFnCrd9ZlO+oyll/nmBne+d0sXPzRLJuSyn3Nhnqqh
Q1hG58u7bCFcXYlW26mdRcNqXjGdYeF6hT6BsJ6m7njLDxRAiyL5kBb7Wd6u5uTu
OVsPaESA0nZ/Zgh5CH6ounvwblAaAPUDdIl+dQUQ2jnrt86uVU8XaUs6q9fanIx2
68CPGBBfDiF06Pev/4hR6HeKHjs8qAedine15I2nxrgK7OHuLivtu6It/lPvmHZe
qSYx6Y6ptW3hm5AyUqJXTK7VTjhoX/noeJ5mfW2inFo0XsXKDPX0o9QjB3ouKLQo
4rjzWERZhZMyLidGAPbHvB/m6bzYciGqP4BLbzT9HrQc/KQBt43bpiHgHrTyE3Jq
Kdcq2Pr8peJEHE1NVpnWT8fNTH31l8sF6am+ajD3YUG1InSjT9g7jHhyVf8ITPNC
o/WokD/NCfY2dlmP3yF52pjrdxj92VhecQvMm+g0oCJHO92PWJX9tl1Re1vSm7ma
hZHdYRykFMNJesXG3igS1PwUgyR1axTxxbLXi5Ej5B3Utlsy71VnmAo4gQZc0yPN
bJTOIjIo+G9iPdLV/cUEBplQzvn0IEExsJQquYima6mPWF+8pB2Tj2kT4SGG9Kyl
RK2970dqvsAMaRqDDXRq8fQ86WL6i1l3xq23OtLxREIu6JntCkl3RrM5a5kwONk6
pc9pM83rruoB3R0YdejQz0zjcnL98eFag9lpEV6iROpvoEGhGUYGs4YbQxDUekEV
PR2FJSW9iDDtwr6CXewgGp2Y+gAOqEio8PR8PIPF6r/HanVvX2hIEL7SAjYolEO8
tCDkEJoicdD1qHzOSjKMVQStbOuWeuwvxlVSSpdaPNX37hJI54+UiU0mRash9moU
eI+u/bP/HdbJyo2SmDUlcP1rDythwMy+pZkwQN9XFGA3nQP9JqGo80lJfS1fQM/H
6H2wuKD+4C0mK3WZt2C8AqgU1vM5LC28yd+KeTGVOEjoDVFqznx7rd60uNGvUUiG
kzHBjgKntXhLX6NT1wNV9H8QV84cOA3+xN0s0LbOyRpycV9FlfgMg0jQ7QYG5g97
xpr0EC52a6AOam5FJYqJuEQNzNb+mTC//gNdkWjpqe2OFes0ScdfDzuTsudyZUO7
RqiD9SdMSYa7HTX0U8RaDQVJ8BEKmlvLvHTah9YVqujzM2pH/F23VvSv7mWoceJ4
LH5VQT+05FdcJBp2O3jAfv7vZ4sVIJUiTqMWYtjH3R/r2++Uwwr+fjfQx8xJZI8W
0tRo3sNnyHDOCv7WlBKcF6hkKlWpAicGVZBJl2j5i7k4GAA8WDH33PBxA7jHpk/9
9YYKdvirWwfozcJmvoW45RqEL0ZNfLUz3DyusWyq+OUzfreGihCkwTybj7Tlr1IJ
c5zZXxfC78m7kep6bLFvyVGoRw4ka3VhrZlJ8WCHpPZ+H3aQq54/Gd4ueue15f/p
5ipATGt2SDG7EwgYlHoYnbl7iT+cQe+lEZCc3z66AS0txLEh3JbQ7rB1vQl9t+TM
CCgUTQGrPpHacxftUSOmfqrdcSga6ej/HpOhUPdDLJHd3EW/f9Ef1/GcT8FEMtTr
+ABllOmj7Uz/1MYHoNta+jPDBrHIpnke6NVE9O4uKJrVC3laq6d1UyFfaUYpSmp3
gDtr6XmMM3M7RtfH1D+qSDpXPxnIGThJddnijTGxGGuxs7Y3dRMZ5AxSQyg+94dU
1JV0DoBM9DPgp1Q41VoCq2c8cpe03DLQOYy+wBTHulokFb0e3Frnj6/1KdFQtd0S
isJ2ZZJYtFWHkQWq5sM7nPEOMDo/dJaJaGoZgLetFdZTb/GQ4Apq4RgC8yD75fs9
4yi04/xPivxnytB4H5CmbT8Y3i+ixQ7ih3u2t9W4++VyMg7f56uy/2CX432kM7Bd
6yscixkicrZGliyldhElpaRp7xV2RED4mszesJtJs74PIp3xi65W9TFjOOnRjGed
BpIbPmN5fQoiePqrRmLWN1EyF63MWeqmANlR7B0Qs15qmiIprJfOkhNha5Z62Emd
6HEmnLhXH3gwzCuTTiXdTQxZFrLNdBKUGaQa4rfuAStzIqBmZNAkePMSJ9a9wpj4
skKDgiL0PaY+RDBEjwcT60/fyeMRcAivQ+bgBJ68MXg42sQbjB+FE7XhXpSaOeJ4
MPmbIEjJCZ/jp//9ME7ZjHJw1xovt2TzGzTTXUbhpBoox7nmy1mngeKIxN575hae
SZmQQ0o8yM7yGTcgt9Me1UPTCtsi41H7Uuu6pSqEyCS1RJKFfZ0962itQXusGvPU
+fFaIoiF05dewpMfb0mvakopwLShux3aokZ0rYejiysq65TtfBBPHiMmjJDxb6VR
z8D6Fm91k3gKSQnR4xR5FevhlwsSgyEseXVl+SAzGJczoFqvcKjuKW6GLDg4V3A1
MvddOMqnqWUeDAMoVpaNBtlY+Shmrwb/bdW5lbOAlbJ5gU/p+whWutVSV56yotUG
7S37pgKsrWcFdZwoj1MoHinQczL9AJwJF+XVVZ/cqyeWkgglL91SXh21f8l4IUVJ
XGvnnnOA0Urquw3/UY40AdXYTnGlEKD4VTKYHmqvFyvvlsgpb9aubXNNqWyu6S3O
5ZMpX0iSglIm/adsjM3aitbuBx/ufHERiKnVGdHDfSgm9ks3yE5FUchhkb2yqsPn
mHnP0b/uqie/9GUaFHfDSVD502XbYXHoqrXnXzJ6mMwMch9VsN1kQLaflTFuqciH
jCsO9vlcTUdn5NoelXzXngQl5rY1M7ntxXFg/lDsmZ9BMdYAM8+S5vlEZZHTEQ1W
uyHNmHJI5f0tA7xXOYL+36GnV0PaxfthiZCDiV5uw6YpLqPMIFQpFdu3t2Dw0qoN
McKKU5WqqXVPq+TcU6PbPJIQSa8BPmQRickEsyr6tJjyoTOCXjSEgN1HCqHeD5E1
hNGgoTh2VT6cmoSnDzFE/4fLdTtab/XiSrCnI+rTfcd7DH1ZqIsgX5EYZbnCl42g
9Ca0EfUsruHfmAVORrrFu1EiIEisbJzlL+grryuFEj6LXN0eRuMJCs7C1NZm7BtD
SVNGr9JXxYyKfvO1dA4txlw+ODYM3hlWdrIYoQfmemyo6U3AW2u31TbXmXf0yWzW
44OhRQ4Cr3utgszXy/IwXWyc5IasNfN3cvH2mqeeXGFVSsPAkesyboNQXlG17Rl/
ygs8ZnDGWAfh+bWbf6O1tDJ/KznuAUTVNkF6H3zQFQBc/tAVpQN+CPTSShx8bByH
2hRWw6iu5yKxGP9apw9gJbd9wA4cJPhhtwQv2mjneuPqYhtszHrZNQpot1RbOyaJ
8C20K3DD9hnsrmkyfM6SrCQ8XwxCp8eulFYrlZpznbvfpXk4/j3N4VYrNZIUD8p/
wNUotaj1b6wvqpX/KLxqvMONx//huxUnqnLIMlaAYqkLJRN5kxDquCv9QFzCxlT1
3u7UpWgdJ0VotLnuAMHQtCEtrAzXJyJu+//tXUErOfa3AfNAOwGFFYJ1+dJyCNNs
sDrf7gKl3FofZxrJG8PGGU29KihQ99agBEFqrNIK5ErovpR15UrmndTnt5cNg7uR
W0t3IEUWtYUzQs+GqVB1tVJ0ijn68m8/HdPgKtzoK4yevPudezOBk3Z+QltSiqns
W3c5JG5u5d1D5fnHKw8e97QjBKpo7HnN0Xs9k9JcPtIKs1hZlW7iGgP5vQjmNZ7d
p6WnFnUT/hSrzE1O5LKliwXZcs3nKWMnYTVPO4NsNQT7cPTf4tzC8TdUfXUuGPwN
MrnNjNo/Wr3GxbNUTIRX9AhWaXj9daryKcA9DTmlFUZuVWBEaYBx9AtQO4wi97av
SD3riOkueBiodiKi85istyWSOTQYlb/O+LeDASOiS7+T7s1zsWdg4QxypD4C8Z4N
QN9lCJg2thG0/sKX9CopdUq/ffTd9nFhJdHEw8ivJcPM0kuRsvIPvG1mS4PUGvxD
Gc44Mc8TCWGNGXj0uYunx1kSoVuby46KW23evfeyeQXGx8AJUIpPjwMKvOyM9VKO
xKPSFB0x297vT5Kp2qOfN91IaCmv7x0uihoM4YQ322pQFiEjWk5dfX+V37ejkbNl
Ua3rZRJJcUjmGQvhHDz79g3xrznBly78HOhyL1Ck1euuJ/W+Azsc+D3O2DLRRMK0
CiDVs/JXcqmd4EiXhGJeK33RCQRsoozzuOYj9Cn667X3ESDoxGamqSUvthYr2wI0
85zrtUZZAqfBhcTUcWateNeFNFlQilSyURSCOX4vpYf/X61pOBAMWas44Viyf3zG
Sq+Oi4mWL+P+TrFOTJYMTmrPDv8g1hl/SQPItr8hRrCmfkuwDh9mXQIOGSnzLiiz
h01T+eBe3mS53T5p+xEuoIUWgtadHfPzklRWSJlC6L+BCgzD4Z3ZvhiLIx+j3WWd
wxz9zx8OkCO+NFVFNvJimnWQxSYvzQnNnOzy3Mf1Dt5cBkTpxZFHojuhtoo7UFY7
uNhlD2j5yz4o3mYlZjQE+3PrqkGl0wO7WfFCNELgnk5lE6rzYj5s0nVos6mTKp1d
d3DBsKZ7fc7VRiD6Ue/Pm/luflLmQXOhj4WBh0dfEnIinlzl2rX/CDTBintbZx/Z
jX5Mw14zjWMGlwm2W4bL06uZpSbUtDfg4P4RRWXiT0XjSHf0/amoAXADDeoVoboc
PxP8jAWlEQwzwGY+dym+1mCStBOIiX//sF5KrOiI0Z158irj5eQx8UD5ajKPphgE
sUPqKkYHDRABT4Lbk/DnAkezgWB6Ym/AleQmlWcKB+HfE8yj9rblNN5Xcwzan0Zz
hfH7Rv0WopFOHveCK88mvWmGc42qPfhBnKLcBd7I+pjYVbqkeuzWb0MtLbIttmNA
XjZrXSKcWcH+ECv7IU8y0IT7D5dKvS50ZWa8SIHRvJ176LX/q9JXkzT+zOEiJkta
7YF8gwGmgfiZTbMVfrJY3kaWTYwj1b45OxS8rGC3E2Ppz8F5QD0dPo+jDdgELJ0J
YWeXyir9wMRyMQ3WoVd+zqI9PWTJppjtFb90ZC38KCb8Qb91f80h4OQons24gMra
I48jhIDtpVM14wnkIDghWrlweoLYp4SnzZ4DIj6xChw7J5O594D63EMIbk1LN0uf
8Etpg/crP+CnClZ8+Psa+7T68+B2lSgBu4ctzYjYSf13M6eFn3IPCB0wPyuMYdR3
+ZXJjUSqPrTO60CVaQCEKxh4E9FL5gRB7nSeMbH4KF4jyhfb52u3scKnLL8bXjfY
Cl3LrTQrEBBDvsCPJqlJmzRq9NsAPulKgHIQqUf+IgkVLtZYYJ42t8clY+7VatZ2
9nCjHhRKmChcd8X4sYve0moMMpstY6x+9VFAF6liJSG4leJXZjsCGSXrVlWEQjZG
h8XiSVuByONGTdzKCeJNv5R1pulW62Y4kFX1qvv9CgYSsUTTKiJgbb2Kfhq3QK4p
Q9Zf2HrKFdQoQIFC3mtImA/hO/h+3r7XtCVfqLQGFQb3O0RlUrltK1u0espMgLw0
lGeWuPZe2V7pXOqbuiyZ8qNJiGDDvE6m/Sem6Grb53lmN+MisdEoNUpzg+eSyDFj
lO+13lpBHhSW4fB+zKkAiInxb3yaMLLavjDxKZFlLuua7zj4CkSa5kEdIfpUwqFk
qukbOl/Puc6L7sfuDKwCmtONX63gg7f8ybE+0IB60yGS9mY5GFpgSbXQLm4k2AFY
rvRgKZiKuV3Fza2SA7n2aKuFzN2alZrGuXfF8XNdPCjeFdLSNNMtAkpPZWOwJXy7
nQXbkyJI6/0vacKHHJdAHaK5QHuFKMT1jd/bIglR0i81bVhzX0PyfILTbr1MKk2j
K3z79jPbwkGoCTZmzlHnXemDDHuj99B6PDpMH8bAZnIZjA7KlErAKQY/TbDA7DAf
Cij2Kn5o2DnSV7VGLxeBovKm1D1KSUCKfZjDjCLEeSWBmEza6VJAIDdFij3E3E3E
MMWGPGGokr5ZDxBmxPvuxJ2wSwfdGPw+Akm024c9cQIXgWg11vUh2QsNu1d+uJVp
sp2Et7s16O4G1NYxNlAj5ZIyIEp5eTMwZ6wF4G7boUru7y2Xni23yCQTKt/4bUzH
f1I1UJrx+6yHTT22X5SeZzoEBgN8Vi6ds1/Az1fYVlpv3wMQdVdtov0E4Rj8tvdO
yiljQWSPC6O4n5wFV478PX+JjIWzQUSQgRfQxWyUoH24/27emw+xF6v/oblviN9v
f0kXwOJ4kezsncpgIrzn2qVbkc6c9sd8F1p77R/Uz+w2Lzt/UPxJTti3F/xcep8m
7RD0EjS6NvKLE2duvNy/Xj5LhRaLjsRZPpAu8GuTP3xjZwBFeOs3RTNRe/MtGUB/
pfdboAu+oAyrU85xO86xjnfGGmHzvnSndCyPv1/OYfPljMYMJAEeaGu9mOi4V1Ch
VcihG4bLPec4MwOMqVZYyhLnFWXCuVvEdu633/7gbZx3/ewf9xmxzDqKM9W8GkMj
J+BqaQ4Q+QD8YJenkcLl0V3zbLMch+7B6mWFYcpyR8UWRq0K5UdwvnTarQOdD62h
2R9CowHXigeV0LkYBcRwpPZ1hE/rd0/B6wyeFutGOBE+Rritzw3BIJuE8WhcnFxq
eechgIhMNJG4YlDlsa9c212FSWYnIEwo6/1O6zVGZuB2mX0xF+BmeX3rG6V8Ffej
RovQwbs/Fy2FKLUfS8OLeivahZJUKtu6yoWK7Z3psDwImMiV/Zcv+bPtEFc1Mnsk
D25vQ5Pg3ZHNzKZOclPkWZd4C1vrYL6umQ4dyf16vbAZlXe9q3+Y6/L18x6prAvQ
PRXwFKVk8uoOSMhmwEM5Hj6Z0vbNhtEiEgfMcG3/aabYxmHnFfnzuZwLxQoYt5AE
SBrknGnCfCT0zvi4Dr+oHIls+ZJGxnn4edtQgksMgudR1xyV3VbN3txHwGU0upFx
ZB/xGAEVGvEdfcddQ0gCktn0Q2Ihalrpd/lDFTi7kiM+rr1z9juPSihiNevX7egi
X+AQnHZXfbKiCt+GOChmJ/DtwGhuqBLNEh8dBbLo8iLg9iIlHGsWu/FjIFfWnFQa
1xfDSrlny5mj5o5LxYGVJriq5NPipzmKYOv4bf6xuTTzVpvjN6YgAz/a+6B46Br4
Z0kgI9B9wBWGA+tfpFnF88V1J/45Xht3qGhAM+PXL3J2au+h8oDoSSWwKUlffBgM
uczbfQuGJqpAocN0zXEq0YqqDC1X5NzSrvq1ZecaXfGNJginKdoWFC23K9aQtve5
YpVAwcbbtJEPsJtSP2PbdHqGxH9GCDZO5nPNVcmAT8jHmkToeC8m7jKkIEayM5rE
EODXBKcjqJ86x1AZ5WIMFEcKIoKZshorXI4CTwjV2tSedE1VmTeqV6TMUEsqPHuL
WjXKfaK8MagM1PnKHaLiwjYzpZLplOhyiFV473GdzdpCv12+8TeIXKeldjFmBkwP
bTssZwoXsYFDLyfrdd5mGZa0b3IQs1eW3nFB33bit5J4pUxkARa20w7Qwn7fkrDP
XDzuI1WRYFIYd0sPQ3o/Z5CbLv5OJBk7cKbWhiZzcmrIdEY1vURln7IDs42OnuO0
uTJBn8UUkkbHP2gbzwHbkxCdZole8lrAE2j//3aYgZWg7FNrYc5YtusgMvZXokZe
fg4Mh6ot8IZUSJBy2SMMiw6mtxiQ7vME+Qlt3AOtGprnCDGkYpzQArBkrhrFwcEG
uy5tWwQXyXbFjiMzZY/LR8V5Z8HxqTRkMPi3+pIDtAYVNcYp8/TsBqkPsPMgGY/t
2lwr6hFux0z1/9c0Us/Gl9zjmF2O5bWbO9qLQgpsifvrncPjs8YLvmjtLPaF5IIJ
kb3/o4dqydNZPrrHXnxIYTKLMpvR9YO9ED2hIa747J9Zuyhd9pS/2rsX3ZC1fizO
5gLAP9ZHQvgy9Xk78H2ZOA==
`protect END_PROTECTED
