`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IUlcXL3WMbjhJqjL6QYw8HIsu8OPAt1kyXVDxIicfoe+u9andrs79ClYvOgwMNv3
u6SRmSGb8j/XC6sS/taw8wdBnFmM3w7MQ/U8GVdR1GTHscPWzGlmEyt6l5HypNe2
01a9W+JLuRIA4rewUmXIOGrSbZYskB2BFXmLmLjCI0BLsFQcnhVQ7UClQi7BAZ9b
37eDtInPVSA4O19IkTlsNO1y9uEq7WCGW1Kc6swHhLfiZXlQj3hG3OEKBc+Od39m
DLfBiSkLTcbmpmAczO+uW7XUebBc8MF6eKXXjrIZvMaUJW2GW9yMs/Ll8oct/Tt3
PAbYtJx11yPTgVjjBikIUAaF6RAx2WC1q/zL39XCYgl0WJcWue8dvQl5RKbXauvk
Wh4LKOkCZqcB0VFUTHwF5HENstUe4wOheuu/tQg+1pLpBxNF7znTwBiDneSmZM1x
lxTXFb1lUtAOyrz+bIKFSDKha8l7vsW0LXRTe9Lr/17vlaCSYnPTPmzBtEQ5g0to
`protect END_PROTECTED
