`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7FOSwI2iapy1cpVzSZsmVFnbRP+piCFaMJx7gxkiXtDMmVfsw9V44uthLVTOWEDQ
serA4QMINrD8/n5DyiVnctTS4f5VHCBYhF7CTxdb37iiCWOnU4fuBE2pwWhIRa4s
8LwOXqNlQucHCOfLbkmfMH0xfAalzfKDCmitFxyDjbHkY1/r925zwiHP1WEFHXtD
H5iF/phOo6XXoQTQNd8dbIWAHoHxTqqC/QwEvAZ4flp87e5v8hMZJ1jj+V7SJYj/
J2kJzwA5qB3vDd3kod2O2XVN5x4A98Z/eTo1AEuf+sg=
`protect END_PROTECTED
