`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
54fKDuhGpG+KnPwAHCrER5VvImr7ipkqpZYDkkxvdVXrjnk8MzbijPgjmEKWaAm9
4CG/MC0n8v3h4zgeWDrvTTLYWyyJCVRPDNM4KF466awsJaIQhx3rzCzFn1gR7gvC
03yvuJoNIMvNpd39jcAw1wZvsWBK/TB8w5MnQitbUXlIpXkep6P3UrYIQhZeeEI0
IFsgYgG4L4Z/2PoqTkB/wW8sbhIwGQl5lFvmldlG54r22J/DcXnK5dbdOW+W3xJk
l1v00on1kMsg1vJbnjmpmovXbypQfzc4ta/L9k/6OPyLyK6h+C+UvI4iGVPfjFpH
4ttwrgH3X+vjq1vhUjQjrRB8CSI6b35uk3132jd27RF3eWS9sOiTfDnb28v+USnT
klIJPhS7wkO4Ds5I9Jhj5QEHdlk6KLKB5j4fvsVZskI=
`protect END_PROTECTED
