`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GRxa8ecxA02HOsyFb2oFs6FwEQnTThi46XZ7KCTmTvwaW1QdzSKNPQPg9VzxTF3I
rGIZazGAuxUsbJURRl67BOZKK/6dxunt+mJlt8juJS25rOXr8YDHwi7qpu+AOO5r
q5/IU4sSi/PeaPcjDhgWoPlVrP8ElfcZgUvqqmzDmVC45A6Uoz3VPk0wG0suOhfc
66KwQuLqSIrJDcmie/xFQlvYw7DZlgOa9b9+WSwAw+Inc0AIie1BUgxeWeLDNkb4
scY9HgLFE85xX3QrSXqrwGHzs03t8j4GNgfx8MvRQ7/vWWGHooOTZIY5KQ2yLjxC
RBem/yaF2ybyc8Cmib2R4WCK3LkCIyZAQF5ln8pIgGDt7sbR4GEpUzA+LiW2IYqR
iphDTW2XRxmP0Gmv7shH4YeWJz7+3uLeYSN7mMiklXxlCeOyQlmTmHmVh8gjPBus
4GIvc5D60clpCu2UmOMcjXyOk47E5Z7kjeZQEL5UGFZPmpMIXBYbjsZrQDNS4Eyx
`protect END_PROTECTED
