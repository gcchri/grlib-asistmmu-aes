`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SKBIlYiWalEJx25rvTGrIRdKgMN5FGol7fTCveM/gV2ATYmsLINxpFuRNparQg4y
DpCp8hLUjS/RDUFd0G6jWMAfjrXGJF81cskDMbRqkH13omuoNB46WcrnN3xRhRPB
24Q9xMoOh2wJZoAxGxu+Y/gZxI7vBkwClilEKJ8WIHzz8Iz+OkjktvpDpyE4kWvO
0zABjE99Qx2xWVINwqzkhVdWMfwvLDFYTJ9p6cCZV1dhBXJIt1rkpkcD4lKMGwAs
LeDGHSFV6fno6269n+SHX8GTBroZfJ9Cuk0wQGSsvtqH8Ix1vspq8a5LWr9VQup9
zSTkQ223bk7PQTR5XlvJPFhxZ7H72ZN9MWEwNNjEd2GCN5gZFGAFJeIli3WH9wNP
rsnypOoMDFcISf1MyTCAzfpiaFJcSsJIUSV/OjxU6aQ=
`protect END_PROTECTED
