`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
94P9ySeZXkp5KYfDppXd3rGU9L1LPXLmhsebGfXhZh+cwVBDh4W4n6/CKmBVVhx1
bTdsRrD0yLYth9G3zaBXJ1Qdlkxq/sdX6CfhW8nRfBqy9fgYDmG4XGW0LM3FjgPW
kU4/j4B5aeHsGxOjN8P7OkaiHDjbhvrIgCeogUHbLlTcx2jT8ALhtlixaZluArdM
Eb8CFe96Tfl9qSYWnzqEyw0FEiFGzjYlUwnPB7G71UcA0cqqOLnnJ/z8P6krqyGu
NtPIAxPD6rmT5DdIhFiMV4dubO1uCWshOFcqBTbiQYjEs666+6TG2t/Dg6fuFNip
U7yoQCRBzCoCd74q8YD4LA==
`protect END_PROTECTED
