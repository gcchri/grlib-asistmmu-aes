`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CYiCe+f7FFQYNLQKes3a2tpTuHumjHODFoqC5YyNIgOZFEo0tuurPGBU0yaeynN1
i7IKBe59R4lVvG1hKVaSwdIHR5OXR7lZZ2SJJUYa0UMTE+ETqZvTcdMaaBQ0AL7Y
VVN2D0Jhee9Wly5GMhabCbQ9FMF139Pb2uD67PCNZaIqw3KdyJpSwtN+ng3MXH9d
yYwQ7pUZaNoDDjUr9rv7lhNcmpVWLoErym/9JumHtWiAq2juezlfc4w4tzQpK8xD
rv83SPXGYVpA/1+5psiUCVViM47XSpOoj0oMZiUyEyUyxjY8YaeGtf8WVEjJAE/x
DzuL34AM/hiNeLhYNtNBiflGoGzepdLx4UFa/eK/3u4qIe4ortlY4dxPmft0jQOe
ySKL5LNodPTt4/1W9nEXWGyxIAjfTR/P3D//octsHNB/Nld4XCs5LbQYU59UHPWM
kE/UUDK7bR95kYaplpjAGR4upBkSH8NaMuvUpfu099F33Wh41gIpIdJjxNKjJDAC
2w547ofJdAvTig0NpWF34OP09e45w/dfdqTrysn8Mx/42cyROJWRIPdT+oh2gRqk
LkoFB69jRX34VecZsemkaxBkUU9DrAsCVcj4I18XjUQs5T+ePRIbCymY0L0DAqv7
eJZsKOyQnnCIiHEFN8DgZwYZqBWG3/NBQOXqTlKQL2kJrTpRWR0JxCmBOxYlx6d/
tnuI3P1W7oeh0IMGgJRxsZG4SGN7J3eLBmNxLGb1I2Rh2/2tvfQg5wGvxTif7hHo
qQSnJurnM+WKYedkytDpDiHXAFgp/G4vU8h/N1VSoQ+zMSFLLpiLLpppB+eU+pcX
zfBKQUUfdvdS7uEOdf5wnMdbErUuiiw0dQC5h50YKsJd0fE1lMhL5DH04gaBSxCY
e34elw4M4MMPrCQLzke71XH+sQCGoqFHLzA0MLJznzELMCTl9/PW/0ryCsZoJVdB
ygou1rs3Dw/uG9lbz6rTVmhAtu7mSq0ZaXi9XdPVmvWtKythZJ6qromm+UinIIxg
qiJ5KBpTT8ZoMioR5tjU/z/VcTH1W24qFMePj6LAGtrcjP8Ukv6fRuhb8AS81Ml5
pSNyDUXris8xCSyGU85IXIs6KJOGlQtSQ1Bo2L+yp1K86ceGocm/izYRuHInD8Ql
H8NSl/JpQZGt+VRc0s7q7eab+qReogBTpXWBsAzUS6/Ha0F24QDn51DQsMSO9/AZ
30BXZ4gX9mR1vRWTDrGi+79BAJPZqjWhXmerg4PtnZoljVgTcWeoGTlpLTGXE0C7
/FGvPugeS4OO2IYJugcQF9ygLpKDqD3ynOnmoxjNtljozq4pOJG3TcKApQQPLMZT
lzh0Y/s/Z3McBE5ltqJFDgKg4pA6u6PC9XVelpQNgJsjK67HBt2oeTPLEYOQSnI7
U3RvR8L6msUaB65lK4L2SpV3NSAxP1ZpEkvRUpt9VhgnmYsCtkvcAXiOIxQpq5jd
XsADmB+QmbfubI91qmITrcyjWUr6OmgkwqyORxjEwoiw5/B/dkX/s1SzcFuWE2N6
7RFRHPvWQaH+AajbjoaRadrjZNs5rcAS/VpDswiBsnnTmF0Wno8ma9nokzUM4YfM
097Jas79I36sIeYd8NOIaORvB5yRuYY9J5YSURezVyRhQX/xopOKemS4s+iEzPwL
L5YEVoYlbY0+BOeNYMRedxb2i4S/AgIqkXu7IfSGZNavINI/ES0juOthws+OrppT
WPLDIeaQ5ZtVmuUES1Tf1mimYNmxVqjbtmzpMyJklqfPoM/xycvIDErgCn60kuvf
I28BP+VaaF267pl5PtsURbFaCif4JxiPT7TIx7/cJ3XSlPU4zNMHV42mRUa29S6t
OpjOi/b2XbH71G00TO2b7URdCvlMiJ3cHCVVxUTtdAcQ64TM8h0/oIrSOPjVEHPv
Xu055SyKxNTgQB/S05koxXa5ZIXlRFRMCtAzgjyIVUWvp/+bfbhU/dMYGBCB1hZy
KRcw8HfcuMi8torgylSlBlcYK5cHPdkxcDKJ1ZVdvNV6oMHD8Tonb/pJtpBAWTL5
txkdklNEUX4gnUBjjD1v5+iPFffeNxKLWdWnz8ZBiagv5wCtwTdV53OMZJksJDcq
1Xma044VikpO2yHjmMvzxRz20zMHZyM/aovoCmMs60zxwLihtDTvGlt5UFDY9rIr
hfTojnV3Lz+EO+tMyocoeoYOMoXh0obMu0hBApOEALY7u7Bg4ussjjudeQ1hoSz+
qGU9l1natfGbrD/Qzb1falGM8F8RuIBKvai6j9kLEJCjo4o5S6Xo1UX48AvmzEs0
i0/m6p8JIZSQszpf7Mzt19zFRacWfsI0iS1BoAETKMiThtdW5gdLxf4KN71ovXpH
IQR5ISIfhySngLTbnJu8vLIXG30WCeLEEV0cYzTvd+DQgXvGZ79ZGlt8+wb8JqqH
GsOXDUcg6pCZcvDZbwJNIUoJqY0c19wFSjRNJ1lZCyGCj52pLzyrTuUO+YWQFCCX
1ufYV+NZ8TlS9WNKRLG8gVI9G3zuu7CKmdeR/kr93i+s8r4A1937G6PmyBGwOnZ3
3x9iZB5OZejjogOyFrwlBSpFNApU49jGOkBGJ9MgEKIhq+B2/zzNBytZzjWMj8hO
/L9sABqt+U8OxF+DPTTjK9WYCZ930XgxT+g/kJF51HZOFf5ifnxJB5LkXaGDA/2P
U5LPR71Vd0YwKScHGhp7bI2TSfDEiV8e5bwv7yD6jlHBDN2CiZW7xSaHHDfNDWL8
+VfIQGT7f0JuzJQ6SAfKx19CAbsOKv+VUzEAcHIluVSEJXr43hIDKgM4tkQm8ukz
jU/yWCvYgQEtriRs3dg0iPFim3ebs2rzX5c4ebP6fkJff9l2ycuGD7zT66NkgZD+
7prsDK1kbXNyhLvXcdLWUzUTSL3DcDln6oNxBiXr2ZChOV0cSAOguyPI2ZbQ1KdE
LSOXkFN3kYYS9ZVPwH/C2f0LINWZeKilW/pkY9U1eGMytKDeLOJQFSnUgxehs8HM
vpw7c5LuiKJgo1vyQbxgRRI/0h1tNmx4ymkfWE8aX7MJ/AkVJ3EmkTuZnbAGHlD0
EluxVnRes/9TT0Kj+gJMxJ5pXq1aFwLJh8Yj3aTX2T3fFe9GrF+vzLEy3A31DOeu
5gcsdbNFKydXkcSiuJ7oPpT8X+HDAm1yer4zLG5QKOw2HRBHwRkpODZo0hy0nmBW
H8JO+RAyiq7XmIYDDuejDlj+XzKUUiQfku5L7hjb7k33dU9sUyOBMZ6rDKixYPmS
ISyK754vgpRcZDf0OXVSVlFmz7dcJftb5n0gFIY+Lw+Nlcldbrfr5cscUAoiLPWh
Ebjg6d0kbdNRNfJyPX3HkJ9KdWlLPAy6y7BpNLzOgb+ZzOZEiBQtnckirgu6LXYO
qUvPHCo5iypCF34jrw6LwiOcaVzsEJbo8JcXH7R6u9cqMF+16XYnC/2qmZocTwta
sYoRKLbsZK4ODuoxeoTYoHoGmD6nKZuwliXZMhG38lP6LXxZ2T1PcL1V0NFPCayC
iQVNCNGBICkXoukF55dF2969qzzQLU/DZ61IuVhpb/ElpHiUz93IWIrtVYpvOsNm
Q8erFe9zTxj4q9D3mGpeR3VVMv9HDaoYGIEkdBmFVVwPebPrWJNO7bXIhnBFnq4f
SaZisXcKYcpxxIZTMe/tXRnaxGDritnThscE1SLy5fGfNg7vOUlGWWM1fBLoXxZ6
0OXlHztogfScKM50v+p+tnVvCSeckNQ9A4zf7n97F8LA6j4Pg4h9VfMnLV6CewAg
S9vHkbv/YBmODs6fZLn2RTtq9eiyOW4U+sOsplB/qMi0K1lI50+987V/5Kth7kNe
5Dve7tw2QJw2fqI2NDE5sfqcSLEY4rcGJRxJ6fN0TtUGG8I2DJODJW8r79qSkUV1
4Di7JdLQrxMcEip1rC86TUP5X1N+nRe1JL14F92KEHtQaTe0QT0U/nA3bzfdCSeT
54dG11FxhUN7JBuD0JJHzwXLpe1i2r1KbunHjov+7GHOugOCtIIp9dpOEi/Qftcj
V6cPzKWr7aVUtuE/DAAmrw9pirAtyAy7ppslO/4HheLn41xTFZsBVZnE7n4Mh3kJ
HmKjo3Z0NOWfjiUg6qU+1nMNWXp8ICVSOaupCYYJlUCCB5iJshRWLCpp5FKC3DQ+
QnZRBvzfpyNdpcHJ82CG/wkwnG+Msdwjq3O1iC/2Jw3AV5KmO8AxOIeybqPOSUp1
iKiIfiWZVIvJ1QN/rF6apR9v2T4ciLA1JTqEMMiXgvHIiNZjVAiVS8J2vekvi2Aw
Ag7+7j1LEvbH/0tPDHZdz4o5RcfxqMa6xIHa0jzOiS0GB+2IAomXAwwlH8ErS9zA
6WJnqg/pI/VHI9KxMOeZIduI1LqzAN+blLO2amWqYNxanHiyPvzcup6Q5dsSSnVO
`protect END_PROTECTED
