`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zpnGrMXN9LYGpUqm4UZeQ1yYeXJYZbMB+3d/q3PwYRU4yAU/otak1sxLplyUz1zU
U3kZi6y4gqC/3I5mLC96SbSATvDpow1AJWG4Ls5bp9PbKhCin7ybDz4X9gtebCHh
OKjrn47CsHQtJ1dlFE2OWAlO/1MFmN5DxDMYjs8Bs/+oApIF6acTAjm2sGwtUyZP
SPUOeba3AuDxWY04FH6Ms5ag5MrNN6KAbQSjRIiS27ct4Ui1lnKjlXeklFXJyeQj
g+m5bGqz6lgtwzR26YY3pxAC4aqtUCdl5TmCvaM3hnZJ29euiERdjDJTS0Ulde1d
auItkrTIR6hOYlMccFSG0fbdbGgeSG6RVdXns4weU4MUCYzK+ntJICHlsv2gPGYV
J9u8ZzGvQNGUCYP3YJBetcOmLuaMfgiWKr+b27Z8oXc=
`protect END_PROTECTED
