`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TMXTW/i2/0+YuXi2Ac/KLPGjkmfc1KPDoGJChk3Lj/MQdrpm+t72RH6gGmd+38Cv
D+ELpNzXbXbg+t91P3gUs2QFErSyNr3mBc1po+9DRKMFCBqGiB4VAmbR3SHVp0SN
xXgF2Q3rawsUjadZlGq2viLN3zeO90j5ygLEhUtNNv4ihD5GngX+W+jcVmUnIlPd
q4+ih+AYUOqZQXY+LwsdHzCr1/OJ9OTwMN75KhhOUNRUb6eXxmv/6ea6OMJSyeRL
PHiVwX1DBcdV9W8vCk13zcLVb8WAdsHhpYnf7QhLdWiCD+c7j2qUxwRMCscQy0TH
IZi7H3X7dlw2P6Da6RIgjiaA16Ccg9S0pUCN6ZS6O4JQN3Vms01pDea/myZ9k6Hw
x/tIBQYUH0HXD2Xj7b8aKDK5k1eGkg01W6KpvHXIxLur+iiYX/VtqEZAb4CnwC+O
j5EhTFKm/FcR6qxKe01JCwSdr86V1EqNmBXgYJf1+NgeMOqcHkVcPmpaf025aWTh
ocPiWiGILj8y9bdbPi29j+dVyNi+ghEtrr/UWJVf1ZCHglh5USoCngFBDKsBfssp
NKTcBL2hqV4pEnsghTg16aMUhZPN/Jkm8y963JbM8Nz4+s9NCIsmA7sI3GHiZvkX
MaZBVenwnDJQU0fWzAuaJeS1npp5l1uZ62s7BOZjC7q73fCOz5tzSq4Ciu+8xmRV
mUAXJXwi8JQc5J29eHIzkjJkxgNvzJQ0/pLvU6nm5rrsInO8oSaY0I5I6PN0z1sE
OvcJS9vPE3N41fbvYcnQAxNKbX/g6hEdzdJERePQClIw6QoWar+jk4DiHZd4SoZD
Pl9GaE6qwegBjcwCyoqIPKlZ5H7eu3L9KjO2EEo+sBYwOlQcq7HdbtGEsXGr/P3D
xiMOkVTAAhWjdfuFBdp0coDuvc3GlMSu4pLMc/dz/VittoVc8lyteIJCccLTFiIq
rnV243KV4xwmjKqjPHuBMCqzM4HaOzkZEguJUF19XT50gX0DdBChfdqLpWZsI5qr
/Lk1kxpqhU9n7LCEi5rodOW2B70ou88aeLJc67s8zyAyCpmOozNrwh+QXAiiR1jy
X4Mufi/GOjfm1qYJdfijz7EYWiFRkeU/AOM/xNJs9CDAydxZYhLmQp2/kXPDBzce
3qBKdzZDmEakQcq700G+ctekkKcq9DECc4ZoQDW10X+nEtlhsbQ2WQsZqqjlhgHm
hQ01X0+D7Moqy7hrNrxEUdxij/Sye7bcykKPt5r15hjIgnWm84oDcqiODa26YBdt
cXVFsEpzIO9t8w0BxoTbQeGsCYDkLiIcQvUbGXEOh0wbvnKpHBNiWQuXph3WsMJi
aXcQnbJhT7bi2Q7+wXSYQA5r0UxvQYsjLnKiW6I6aSfYh5IGqhdyD6sFGMA7Z/Nd
TQkbNrAxMvF/hEvGFdC7vYK2g/IGQFgK0sahxkMAm3Vva0FRjVId3/tedlvEsWEH
1/XUxkZyVdqcbfnZU7D+YGDk/i/S73BOgfdOhinPNPnsdwEl8+pKpc1bouRfWqMm
dMYC+sZQ6TfFf0EqUYJBQLbVqZS/HT2Qr461FSmz0SBYpngJGyHMp2bS6N9WkEcT
rD5pxQdVFdKcgtE5147Jzyj+0yK3tC6m+I84pGcslfXW7h3UAgnyB5GSrQ94J/5E
MlxapTpDjYwqnfl+ADcJ5iv/wX0Ytqjdtrz7IHJHWOtyci6nZBboEiMWkqRsf5J8
3WoZAmsI4Pp7u9gIeON7v7QcpAEbJz6cLaTzO0nsjnrX1O1LNznMbAkCkJrczseV
+bbUE05udpUV+RXsZ3Fr6jvV0f7/5kV/N+LxIDGztBiyb1ZHyWxjFg2Af7mOn8+5
LZhoMVfTz6YQ2bMojwilfalYv9sAgl1bd75ej2VoXMLFuSGhhESeZ9KmZVEroLWT
e8wZ6W0foBE01CmbJweb03ppxkJqyJNLugr/lXOaQCmevbZCEOld2RE3FlNevrj9
28Vbp7aHjZ51crwbBsXGWWuJyqzHfeO618qP3vvKKJdkn75pjte3lVCqiqIYUHSW
MaIF8TGftMvr55fXYymb2Q+2y0Y1Dd/Wwr+CUyVIGyawvAB4wDMPNw7rOhg8PGz9
5+QPnT89XI/I8FvEoFzZXpeVjj5ioxONRf5+7oA/YpO7K8VbeB4SYKemD7B/stGC
fx++8NCnAhuQsVuzQQETLtUw9TxBszcr6ALIAKIi27kHdKSVjYJyzSZxgRQtvUGr
wnKSP06Hk31kRO8RUzRitNu56fd0A61sdxe7baC0jURNA1nmaOlHrSH+k3uKwaO4
edN01YNwqAhBcX6PDuYAlSZIgQce+e/u9pufMIFeoGUbA283Lpq4uwbRRh5siw4r
oOCSYic/T/c0tUf5bDScIKrpWvXhAHGuEMEeiNERGg4Dp6wCShEcULev1fbGwRhL
yJkTkPyrk6tG/P2tx+jHUhxLz9BhTm7uqiaTywra0dalpppKNdn/BNi0CoP979bt
NHW7kBaZeZlJ8pxR1hmQQ/hjgWMfnmlko8XfSEBjFU9bzIvgz1g7x2hpIK7c4FiK
`protect END_PROTECTED
