`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WlzzPN1ja6PQaeJdO5OlcsdwZu2S56lp+nbMWnOEJYvb0nUwvo9isncEosPLttyq
TR57Cdkjh2kq19uJhmCPeaBetC1DfCeSL1kU9soC7GJZkLDwG83RXFDea7H/pTC6
VQK8qJv7WIJ2NoD6lgZj5+nV12LXDVjk2m7hEEtKdBVZWaCOlskBX9Ak0ObDKNOR
wLqYrcKR/cQ1NF3iOJbVcyib0NItti68PRtOhJ/U9fpxdo+nukIcf+eDms2OqvsJ
OMzUGfPOKcEnE9H+5IyIBo4QGEKTZf+I2iu358V4P5pC3jS+99qkLpSgf264CgGU
LxF0E5/85Toa3EvDp0muVGccHShK64b5oZhdDBic2GqJU6cdjDPVWg0Y4VMmBkHB
afcaMkt0d1P016bPONk1derx0xxc/Tf/FMHj59mEEy40OVxYJVClG7PhxyE2o7VT
85Q147CCMselPGZc+XjbtXYarpkzYBBQhFg+SdiwcAWFFow4YoRc8tnay+joAtvW
U4Za92Oyv4F6ZQscn1/3PkmknfBrVqvQA06fciWVnYduGpwyr7fBOD2wMSu9tFLe
KgcuPqBoOiiSQUb0Vgj8IyM9fb84yb9ZFKNhT0nek+JcA9VL0uDPsPqe2FhWqiXD
VQi2tC/4xYefhBGeuqWre/HjYKBA+6DB3gaCi39D7u2BsxTGFHm2oQ6V3issxJCF
UZJBfya6gK/HoiqTCMuJiD1T6kyoDNTDNuNp18p4oMbhhZhhhUP4j6aHv0/o9S9x
Zgt3WbVhtFEkISBDiaG+7gqcdOXfCPAWJgYtaYIg+96YO6U+6ur9iDMQbhRqaskt
b5I7hMUOU2ELxdLpDKjWhB4E3xZL0WxwJyNYp7uLnjp4l2vZ4Mhx8+Zi7G43ae7x
AXXusYSUNiH0ZZGobKXazmVXQuDHgkV62+G8ylKPPijcUobGmTY1V5bl7/kl4QrB
cofO7XwjnYG+wvrtThucvXoz/+f4PVRgBUx338uorW6aF1M0bynQJEcF7BK6SdYP
24bAxobGX+Wt7vP9mjerjKSr+f0+fqEn97C8zEbe2SsPAqbWS0Gc8u4FXjyw4jTj
n85d8j+dImn4jnGBu/7bAK30pt4KiV3Udmt8jfBPg9ZKVlpnPSmnoJUXCXTv1Z3e
zW01uGAFMdhdWOA0uyvd4Q9OoITh4bNrfk1UZ4Rpy3lFYpp0ZmWI209fhNMS/gN6
S2Yk8r8SQlcwlSBaandyLSJpltgyuzVPfDMx2dxLV66W0LRV53P016Z7O+pBfuYV
92cJh3LtuhAD+A7NkvOUGLKeT4nSulhA8ayu7kp6nfX28dTbPTp3dI0IF1DTCLM2
`protect END_PROTECTED
