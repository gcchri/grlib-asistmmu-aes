`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wL65KdNnb1G/D1Cd3+6kIBTUPsOCT1BsxdShOaJHtaycbwCSGmoqlZylRPzQX5Nf
twDAx/SFiIfeIHqd4pTO00mrWtrkyUEWXO9GvBgXXp1H5AHL028/L2rYFTWVifkN
HgowZu50PQJc6DC1ETqwHfyrOql+8hy8/ZncvrGqeAeXDeNd3/J/YRAKPmdowIoG
bG5gl3MN9I1E1dycBUbhJ1NgbM90hxs0RnjTSBfIry5DMakzjfoqXSKYPOw/fhCP
Eu5sb2FYY/kQi3tDF0pc6gQm3WfcSCtghNslZWIuF2bZ5XjfLWjRFQZV8gJUS3Dg
IyauPKuciLhsRI9JayuwwguFGDI1L40mk8XidjMNo5IrKsfNDQxiBpNsU9M8kday
2CDtPlCtRz5NejipNpoUcTDinJQ31q7g0m4jiceWmOqtPH86hevo7xqkofIkKTBF
IMvzOkesgSqcSSC4UFOxf5wBdqQaaytX4GRjCCrlEgWFYr78OArl+L9RTQIB88F+
1lQ3vA19r4UULpieyCdnTKXd4MshUU+rb0tdti2JD4SMNFQVDJhnrzDschhk9cIb
r537vtI5+G1Iva8p4qmmnBg5uRwHjvIqdA4KgLJjTVA=
`protect END_PROTECTED
