`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DELM1jQ+zLx/B5za+eBbPjqt3iqulZbJUgrQlq5RT4a2m6f9sK4+n62OeZvIxV/e
kwMmZLQZCxi7piMUjQY9rElMpSLdN59+Y+NqLAx7dLtW3KHaF7tCE+nSJ+jvH7tV
1cMFmUyt8CeWu1xDbvpP5aH2nvadzoCSI/m1Yp60sAWHCgo1nzC7V0cv+qtOBXzq
uZoTpZsOhaXYMqiwQpneW/lM31+o90pN7+DktLsZhe/TudpOOBJ4YjeXCYz5bAJO
mhm4IYLBVpIT0ZVsvo98uRf+YQFYojhEhz2By9kAJwUxcPEHF8hHbTQEV9vUl7+J
PEgqeuaRrZJe9iuKRtbArO/+EZUUk0WBB8BeqMFoPeoO0iHHtkJHt4qb8fqMl5Pd
MSbgGfoefWmmfDnQPQWshDnkiWfFi0ynjlahztkmbaM2+TCDGTlmQS1Aq/q3c7zD
Nw18dJWpLNKxnmKmkELOjw==
`protect END_PROTECTED
