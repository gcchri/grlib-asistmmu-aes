`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DlL/yUEakv7tfsUVLTzh/mbYrqk/xEIAQca5zzz6jbhqwMT1ttzeghJ5ySwzfLya
Hc/R2VprL+ajeI4XCHlk5nB5GINt75BZUojw5GwCsK8ischj7zcO2c76SLe/y/R8
ElNCU7+uxhID8wurmFKK4qLCGjvTOezDqdlX7mlVqJ6IdkN6KidMbAuZ6iExPP/M
fOwK+4MDffHusXX+jeCt/yoOp8ormLLqU6wE8K31c/iisHCasKVHgXvXlLtd1PGH
6MN7Pk4G9r/0gKhkMewQxbeTnYWW1+m6Fcr8/QwVVe7FS3osamdaU1LX14STdPre
WWoglRxL9x9+ALy8yYGWTEn2ZO8MNCJj/o+gJoyXyQqMdN35wF1HdxF5OeL/XDV/
coeL4POsYYHIePuS+DXSjTsSvvkC+4f+DZBg5weT9oCidNHIkRm5P+w7tbYQrDBi
tZQypTL4BvPzSOokgVxtA+fhf8SgLXM13FumyZt6BPuQquvc7RSLVeCC+VyyOSBH
yZG8HyBdxtIvEbEnP9V7xKqkIqDEDbhm3D7iAkn7yQuZRN5onzrU53xvGSVncyAq
lQ589W0W9PNRbbx9Zvp4YLX5P0j9Co894vej+U5sHon0PzXfG8sXIiG9pcslm2nS
3btsl3aiTbz+o0ma7OroqVn+JkpzlVFVL7/ViBsZCM0AI28/xxNMHTohmiH/RSka
/XRgR1aucP/3pRDxnx7MhNj2hgclW56SYntuC/P/orYCTuFlj+/esChiimpzjt3S
07+JKhLIW4VIj0Ukn43pgvGB3cioO0TalJVCMHwgVw6RE+91Q13KAcHPZzXvSIV+
Se/ow9TC8kC2BSZ3Ei72lcECLiw70BANrCpiPRjmtTp7G/zRGfFbCc1n/voAs1wl
lmV0Ieim4dMKm5m/5WlL5j8UAx8SD0fDjXJtPc7Tl39knP4/xTgN5VFny+dF5dB/
pLqvJzJaYcr6XayzUVk/Ow+799FJOBVbwnQ82gHQ/fBucmeFVwdrpmsdjQ7j53GQ
3fLdL+5htVfMVkB9sZjhGLEroUupUFeRyjpWJCzOlGKBt9WCdlqmrAeu3dJQwvq1
t9ZD95WqhbohbOcdxL6WD3HPzseEoZW6arpGuyidAvQsQN1Lq2lF45zPKPEyPw7t
sv3fP9VbK/uXnBxpK940P0kQKTzm6B8uTqQdSzBbMw+R9pnAE64qzKi+Khn8uwB2
GhD3LIUeN8//zY7DHFjUiCkN7NI4TymRxwrebTWQt9KmPtLCe9ZvQjZZ7rbDsItc
`protect END_PROTECTED
