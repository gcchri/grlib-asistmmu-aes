`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HEkHYUV1RB9VxNooMDdX9ped4jSzsJ6baHsy/vXO2Od6Sj6kaLJdliq30Eu8xHW0
/VOUqUhj1ZZkcO+RmwwrYYztEfhpxXcQ+fBIUgJngwGSOLNd5kR0Je8FmIUiLd+p
URrZRfwkgxZGbWO1YN0soAJXWjyLHUQzyAhnV6OZiSJO63lEdfvo0cXtadngo5fH
FDdksFDRaE3mQA2iRcx1DebuL8ctaapyupYmW8OrT0MA0Nz2upOQHkBdPH4ed73q
SqYKFxlenFq+AvCyi9YZNhqNr7fMxgZJo6b7jGR9+68du5uvFKokIrmhDP5/XMz3
9cxBMos/T21Ww2FZpYTkibbSTbMl5qEjJuh769K8u7ZmXc/K0w89Uobginb4b3a1
Q1Smbz1M2BnXKYZmuFTIEFvq+/snrzekAL2gEp2BUzueHYdm7RJAXcb8CqCnPTcA
EfI2/2LcY3x0MOZ5Idd2lHhRQfzrQ/T1wW1LiY+7/cMCfAdWnjsCzz4SqlIuClcy
slaqDBWJA4YRe2igEOBz4yAj75kXazSkZRHsR7NOs6Cp/N4uKSjec8Mdq67Ktye3
lhdgRXYW/65NmARxSEybbutOl5od0sCrvn2ODxSw/u4=
`protect END_PROTECTED
