`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DY+zpsKEi7KgJyFhMGx9sWG0WNGY+erjg09BfNO/VME/MRBLD+CbNz+s50tua8d/
UyFk+oYu4C3nEdLUHO0uYYp5LMfrR+3qOSFy/uxl/ep0EofgdZl2fd0L1krES+D8
y+nBych3YKEOrI8+nc+P1Mb5b1FEonUcbAdw/cnSAyYKrtKNY/3bkNS/ueD812bj
neVAzQppnD+NfrG6r7Fks/2+UVg0g++vaNWynBYQzIm66CNwBB9p5XXQML7NAXD9
/4JB7Kiz6wqlfYLhLRo2E103AhqkwqL6j6In+VPZUN7jU6mg6QoxU4/ojJnpVWHu
BDVwaJO6DVo7Kop3F1R0eMvzhK2UcDII2ipoAcyZPJhRjLxi6e3udDUaLXVkjOvG
ddmVU9plmXzQxdX5NAEkge++3H62bQyCtam1rn3FjEAwLpKS1MBDX98XpTW3OR9P
`protect END_PROTECTED
