`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p11xK0dpK4HLfMrpX9hppIujMElDt7bTfknmrLQ4r5H9i5paEcrSlPeswpnUrlNG
EpUMda6RF0zL4hf5NhIPmd8cJLAHZXtp/QKYgb04eIu0OyaryhktjBHaHaZw3xVJ
7eSqpnDe37Puk2cjnRjHbZx/3LVf/Wo/Serz9hMwh8PprovyfFEaxBBiEkEMSmwE
Qb34PZIHVB+6azlEf2lrGH492Rzc97eSN2h6dUzkcVHrs2fN5VVlyqPj4VMNKJ6O
IPHAOK5t7CMRXxEqJIVnLXOD4X5RQTY8LhtP3TLI7KvwogPEUSWNWooBcrqywEV7
C+aCbhscNNpU9/ExpU2WGi2LkiHFhGNrVNU3kW8BUaCJaNGmbb/lTtKfK2KWUxej
fInVnRSrKDL8reYaNXieSEnOVBliXgOF8wtZRpT9rgP/IOir+dU1I+jetRSIg+yF
TBjUAh2JB9kNfeAEAUAqt5O9t+q7sXkpveZTpPE8nYmO2f+2qzwNbGgfyigHxMQb
6n5JkUXlfpDd6FeMj4iOMyvCWn3QMTPVPBJn3gW6w8orehOlmevPZBrCRmv2jHs6
3hBNmfO5CDyJ1YEeB/SnJ2VOvgvm/di8Pqty4FSGOF+QCSYQcMEY4yDpgnMV1FgS
KoaPJauPBUSP5e7RwJHHsKvXQj6MkdO4n+6rXv+wjZT74sel1kon5NbEayMqRIOM
UGXyMLe0ZBJJwkbjGHSJ8LRbwkLUcQIWkNbHqSqy8EaVO00ZRERBoLh3lOf4jdOy
akH6rRJ35TUP9pEMQ9544g==
`protect END_PROTECTED
