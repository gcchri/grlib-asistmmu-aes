`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
79ZZTkq3SWFscg1wGZG2elnd9UomxKux6uZVK4flTT3cE59uLbfASRAClSphQ+3f
GWJt+mBebSvSCdMsLiCIXAKPDAaUq+q37Wt+0MiL9FDnV0v1D06eUSVwaflkPHiJ
D5SEwm3IogHWY5VotBjeZUbvQGpaIrZEs8kqOoGliIQFY+k/lV2FdSijrTMTNbU6
1p3449HE/9NUVCZtkxNN+q8kI7xYXEa/9at3ouLJru1Kw3LUokkChe4SvL/JDco4
d2bow6EgUoU2UM7tX5ncaxDdllXZCvccyR1tYUIOMEnM5wSW3x7DADfoCWy49EmM
yAe7mHGUyeJVFoj19ii9BCZew7S8iWw6sEPVath2BdSMmHgmM+8DxAOwzGrxlh+S
UN6/1fP3RCxkMPskFXPxqXP/u2uuhLpheaIT2GoTilsGD2Zq9Fle+4aosbrCKhog
Up99QI8Y+UfBmpAveQwTfBZuJywbHQAIdqqzUIubVmxQ8tf+0I9vwR95+HU9Fzhu
MeO5/zr7MYlrMZX7V8i/sUvmQfwy3Zt0sHAr44+jIBJkH+f/bSCx9RG4KqHHeztV
5C5Aopj7i2OPgneKepIg/8W9oibeEar+AgEtMjQLHZA=
`protect END_PROTECTED
