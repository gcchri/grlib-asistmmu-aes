`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XV1WuT49sJzlSrEhG+X9YIm9vuiREJ9FtE1lfhfUHJ/lxKAXX6pVC7VrlCif1YWv
77fdBt8twQNG3hfRgS5R3VIpieI3aHVeufjeaGGGSZzrZnWf8cPr76K2ZUm8P+1C
arkuo/h3LrGGDTUH7qKKJFeovjmyGQ0XnR6y9CFNMPfPjR6B/qc7C8oKjyhojrlo
IBCZtKbsQH0+jJXyi96LAi8oQeUWZU65usS2+YBEV4XMrJ7SVG9HHjkB5R5Os16F
pA59nfA8G6+K3BS4SiZfGzZaeSkCsV+ZBX7krSUH1iagG8ipdPlAMCPv1xX/bCR2
Ouv66jnab2SxhP9SyAm3GQkt+jKx/a63AOe8fIuxIr35AryzMMoMIifAxyHL546c
0CyMGfJgc/YDnNjuFB4jHzp/lmMP7xTg9azV+Ai6uTPfwuAXxEK04hv27f9fWOjS
GhvXniKFUrAd7nestZy8wKi0HNGxPxvNcCW203cka3w=
`protect END_PROTECTED
