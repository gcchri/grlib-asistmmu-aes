`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nxSokZnp1/hMp7wWGJN1OLRux5Smk7UYZwgCq/+N9oBRwJ7M9GwAe2CSrN8W2nhK
+sDcX5m9g/kEiax8VmxKXJp5s8dUFnclmwUZEr+mV/S86GvUArP0QTa36tvPCo+P
Ln52FfE44E541t7e8miFRm+8W4LY1nqS4EU3t4ndcQrS7kWi3GWSr/IL0jiRgbVg
8R1xKVblHLsjLyb4xAGj0rMAXgTe+wDSsN0knRnbDzyWw9SHCVT/6rwD7FvFULr2
biqb7agAt3CTZa6OhL3lAQcJ56xqSkKKeEhNA/k6Fu4KN4vQLCwhgnV5zJ5ZJP0d
+CWONNHe+YApZFb1FDwDbIIPVvEVU0kI//Ba1ySpNmKpVqlS4BUOHHUQh1mP8mTe
OaYREo06bD5HySAKOY10rb9kgxfT30LqrC9TEEMD288XQyrUOSaGLyVSPWgvudiO
PY83YBODxbY1ENFleZULwec1UcBSdBntkiePmOTTPq5KjQRkvu3SrBoGIK/CTH/3
TCF1siXd0fZ5I7UIuTBPM0uZbakC17RjnX+MFh9BLJtkZVWMFHLQBelorfnYftAt
wqTRtr9po50eT6abgFK7BfHw/VJWIFJ09JHwwleTzcBPJ2vggOvd4Wklu5orjhqT
5YG2YvaeVUgBensjQVXjei81qYPD31tlCN5PbDHI72wHcMkoIdqebGuT0bZOyQbT
9mTbXHBtkoSF+o5Uld6vY7Yh8V43Aqfem711NLF9eSpX4XNrN+ekLoy1Ng2fzQXK
ZuycokPnNCqFaYvgHlc5rBa+LwYTGx5boUV+lsYaqBwYLoi3qupTCdn6+ycbUWBR
4bNPbzWknTNTrejAJAlpQ31qq0H0ICsuW4uCm+YCVvsi3P0xDnemv3OYdW8FYhLX
Xw35MZanAbHkmhV6ArXf8U2fwDWPoog1sKXofl7ep7zVULT/PxwRRpNhXdk8q4q9
xCuOZQmIrvaH3Pu5uCewyVwYs+E+eqARB8ThXyfINnt/EmxnGXe/U7LsUjemz2ih
smI17SNM5rjNd5yeFXb94nq9GGka6ogtHGrl50wrKY7PAkjJrTEgUzRmd8HTXaRw
5U8Z5ox7ZbnJgPKSp+qj+NPMwhF0eSaFKU6/20bmGk9satfnWEpIwefOGqUIQqaV
6DwJqB0H64grNnPO1YwF/PT6ThzAuMQGqtQ/Bgf7H1MVWwW4yoF2ZVH2wT0qREFX
Y1VF77AYzJtcjI0/L5hgWaSsMYKXrEWrakesSGKgPfuTQazdBMdRtD/FO/Eqoi/p
lPih7J7HDUoInMX8xY0OOxVorZ3SnPn5dlAZpknp8vEBLVvKmxqDqdGPy65pK51y
N4p2MJ5wjqUXGILTIVQzQQw/upWXeppN+Hy7FoGCAfP+QHM5zrvSOFOU+sjTn44M
vVi8CN6y1UHKPFf3XX9XaZlC5/QF7vl73sxBinez+D+g9gNcjzukkQ8ZK9TEirAc
9k6lWuyLvBtUDIOVJKherQtfyvs/SBz3AWNvfjzAmdIxm5sIb8GEp0ljq1O0rC8v
g/BwDw/SbNg7iYMyvLHYIQCgb6H8bMgTs/+otCytL6ouZTAR08P4JFPIXCz3AwqX
z2PbbgUijEoUhFBHMzxE+0Exa4aV6F9H50RM8rdzLOdqu1in1wB0ivGd2GlNKRZN
Rdd00Io+k5VZhah+unrP9s3lNJRToORNXOtKIsYQrQwDesvRvFJl6GC/mlyC7vSv
dvnsnebtWTDITb7Nd6euqNGkw4L3CcgJzUQ1ShjyYtv8C2YFfKZhS6bA9LdP05KX
dONpt/oK23ZD1uZjGI7B20bHCf3C6RK/woqiJjb0D8ZoFreBd3QsVzBKkTfwDZkT
lNBUuxPn49T8G/rWT1veuYLdUkLxs6NsGP7xBkIBcdg+If3TACG+q3RHlO36nSwb
CByqXDZ8nmtOw6C+H1M5UG6tKm9QHAx2sfz0HlBMtF0m2DowgNIYibB1fjhu8wxd
H/0b3DhYsDoqht7o70OLJjy9IKRNMscpdNmEeATTq3lM6pUIMLrM+qfvnXE+8GmJ
AEF683N6znicaR9owupbh//RztZaXUulxNvKWXlgEZjijnMca8B8FwEa0Oho189O
7I6dgXjBwwdSWFlFv89oCjfBjnxUZMzYDiaI4BtiZxI/GsDLCo6hJATA3gsS7RW+
gythpTZ1WbjlT+CnlztGGhBV0nSZ4e1FpWDla+ivf+ce2MKrIbSg5RdIqDX8bBYp
+G2x1cRLrgIU+A1THZtErIjiYNl3GkQ0GNgHm5gAAmlZQkuoMRG0jnG4MF6yWJeJ
qZ0lKbO7unynStWZBia/pvXH5JmwN0mnRQub7H3aalwlfPxx0fWS8RaX5UTKzvdm
2Rp1Tbwd6WSD4Tic0RqAtsEdbYGlzJo2sYJLpC1cYH4rZVxubltoj6PrljnPRCQS
q1xr/mpPHVXcGujRfowLJS2j6iG0s/ygvBk03II5UeDo8grIq7oHXEb/f9AuCAR9
fVRmucpoMy6rWsUaDAkAtGP+TAaRfVWBOiv1hx23/tdI/b0a/ICmq0XtnMNbO2jj
NsOBEojsV5yIslwT6AJqqgsBkiXiATrtMovF7Xmav788g54pgIxW3OHgZjZeiKzr
Xrelhtx9Ohu6kNG6cD+VVMrpev4AcqNKdhvuizx2m0uZlDOjwsYzJXrfu7FkBtM7
5VFYvaBC0A1kuKqB6r8B/PtxSidWWZVt4i2hTDvBWefMxOizcsh3sU9T4LaU/MKu
h8ZLJd+GUdq/VMpTv7BvS+NwgSDTd92A9rJIWVpjcCh41aDZF8vhZuJ1qvHxbJSN
QeJlcjins/lTvdBRU0Qq9mJygjzOYUvsqlvcISV2bwdzgyU/enuxDddrzR9bFF4z
JZi4xLFwhbcXvXb4EKXx1LZtppRYmsnjjqhBxd+mwgtgOxr+NQOAUArBqse6Gc0B
ILkSav/k6/X+CVYk/ybgqaqgTeynWxrEPeOxj69DNuMchO9nkq3OX4NnlFmDHp/H
sVJCgPNFXprxJEftLNSZhd+cDDs/e3rGvZpQfT8eap3WqHpVl3Q4+MujiWqRvW9t
xqSE5Uya3NdH1AqyD2LvGxgsyhXBrPAqEvdQLMRljRhypVvFJYB8BEYsm+cDsBnC
BtNUQbrLMjt2fSlg6Wndl1R8bssnH9Gzf6Hbf6/QXFmBrVDNBEBSZHsJSGYeh+XI
Ei6uB6VsRSGzOP7xMl/HaLlB7+avppCzbN4SJcPzjIiLwtZj/e9B0FZ4D8urYEij
NX+UJvTaUHCyKGEI/5Tkq+/ls9/WgBHWw+hgbDZ7RFO6n43PTaT4cGY+otA6kAyw
j5X9mnNrQsCLB16dAh2R4ZxWAF1VE8rjUMHeI9hoN2ptM8h3sbXx0YXRlRhfRU8I
XD2Kxybifr+6/BhfXK1WUPf/vYnM4MvxiW4aJ91sV6mFYkszuwBIRRQdFy0mSfzQ
pUCqxYJqYRKTFY4CnjHqLF5nA07howNnsh5eOGAsup4Vg4gjDvK7cOZh0e9ZPMFB
rNYymscIDLbVMbNGjXl7JT0VebpnrQKqjmKog0mvoHYe9/cvXenaNBPYyRw6UE2+
gP41gicxGjcO/XSan7LrlJmjaCEoPy6lSUgDKM6+dCJgpVp37A9XZ7nIM81MNZZY
1Zv3PKJTB/Nm0m1iiwRG8Kr6Z9wzRl7fKLq8Pq7rPrpcmR+C6p6jCuflFo9AayCv
qDdG7OET5nLrJbtsLYpCyfCvVZI15rp2QMe7NchDeVXKsugxgjgi29qT6GV5eHgp
WTAUA0RtcvaSv1CB/R94Qy/qNxSScIpa1tEXHzxgwzE9+7SRoQMuoosKPMdBo4xk
obHWn3Fi0h4nAzVH0+vwKtzWQJ1J8GcD6XRKA19yeGEdzotzVC1TIu5CfRFldHR/
eKEvU7t60A2KMFnhJ097EDtte7Srhgra6XYq61LQwI/Wc1Gy9Hen0xVIWknDEkD8
9qKRD3fAJdir0Hdfc2zJd/HCcFHoyY6vOoj1O8/CwEPEv9MUKvJhiy6+lQQV2qA5
Rw7Q6mWh1+x5zTNJLWjZsBKRTezhkWCjgEvuWpEONjIdiLYu3IgzH5mKyqMegDW4
KtJTimhr4uKa9iXDeYoue5AvGrFfaLL8iYpdW1HuYP8evIWFytd7nAETJehOSpil
Khbw3t7R0eRejNih0y3ef25eTV0iKnV96WtmE1bLtfKO3gEsQwyQ5i3R+73xT88z
CGdRpIYxFEhZJRbtxxm160EsLOWkeUp3GAdWhoP/1GlvapQcktLnCXq5tqfitE57
hPWCmy2Es39V7krs0eOIEF5UlsQzPpjAeOFF30gECE6iBpUGaoN8iFDgitkoFLaA
EY2dKTRsHcCgcg0gTzqaDBiDX7VTqk4zVrMoTZyE0rkWHzQ1TKnlD/p3kvmTzRUi
yUlNs6ky4OmHADFaH01Bgt5d3TZUYtwXbtjl/XUylXyd6ZUklbioi5eEI51/LJIc
d9qKLPF7LlYRlJU/+w05JV80f3LR7K6FFySoAJuBeO7+iBs3nFs4x3W4eNWXJGwr
KHTznzmMNuSj6HABkagrSxd6o5Fzf54z4mL/VvEGy7aR4eRfFNFkr6dDs2t++d6e
19mt1sRan3kK+kBrAzrkYRZqCM5sC2y9M7HCBidSTMoubaPcfif18fLnlOGITU5F
AF3s3SiY2Qhxezz65Uj6hoN08eFezWLB5KCl6SzbUl9g2lw8G47huadEYSpbC7BS
YzZtjlBnOzhBnpOjuDzDthMXNP4DE70lxbEhwlDAZHkcx8T0Al66kVC2AD9YpMUc
Qbdg7dlj4ynQSOI0BuxS28jam0f5dKDUs4f6I8e/v5Ul65cOAldXT1SxHbQvyIwn
fTFuJeWWfnnvOjKesFeqA0+nCHWGrqDkzn5QWdF4908dnXWFjXajII+gF5JthCb2
iKmyb869UOaB25AP5bMcoua0lgOeV9E5CZ6dguZd8r4ykPm8WLLE6hnCi8KxEHuU
EAS7Xq4RaO3K+0dcRSHuImEgCZwf8zA3OJHMxiFwiWYZbSCWwkCfPQ/uozpw1oMS
RZeEEj1pSn0G/glbSgKwsUeSt/QqoL6UaoXhdN/+42crYxWMBDYSD0C+Zyhowecy
whDKVhtaJWL0rTczBwcJ7CLZ8GNr7UGAyiXqei8R4fLYYKdAah+dFt0i4Lt7AIJR
xsOWpbj+vrCUyo/kbdL0IVnJXv0RoGMvYbAhiFHjGdBZxb743mkHtf4j2a/pjiE9
2nyogmX4/AvdEetGSu+YuMMFHLLIFeYn6wXbMgiEWe4f1yFdPbJseNs9xngw/ZEz
LuZGp91723Ne7SYga/frq48DTeF4X/Ys+HGaZHd7jJmNKL5kcAS63tbd7cnsxzia
APMfchy9+ZKN0pHxHcJm+C/GICxDNdgBfVM1P5VnzSfCUW2t61feqlOLsehVckPh
NbOQvjytHf0VsN+twJC5E20sZYipbFEQCr37He+PF13MQhUOszmbaG6XP75i5kNk
CvgrIMnCRcE96vbUp/lJ7cLMZXRlAR/QOMaZ6LoIDAFmgTstGjX29FYYYmtbiyWr
u64ThrvIxINf47uqZ3NEyK1uf/gK9npFc1pstSCMODpDblyBSFkpKs5XkTCSBJRP
l2PQdKDkvT+gB5Xv7LMu7EFNiHqd26OxcOjca3fTYjb5ooFzvkyUUyk8Mkv42KHQ
L80Y/YVirf32yw4RE+0uo2JZjmFoJVxYjguupVB7PNBKR4xbWoRe8BqsBsCLL6B0
+SscsLISjOgf6xenYeQgW4/nMyumKEQj8AZYgAZ0st0aXjOz1uz71YPKkOxj52Qp
CuWP1YJ4GGJ0gEsuK7Ot9T7w8dJTjEqH9G0LAP67L5hXp9J65jgfPPUKIrFaxbpJ
r/HAXvRsnSEYMW5diBanFjQdrjxkjvZN/r+yhw+55B/YcTzg5nuWMguccmBzgkuv
eSReZmTUACQnDAMnnr5xN/SGNGwg4tVIQoY7IVKEmZKdz/5+TufC1eWN9H4pScug
HvJceLmBDapB2MhJ+AL6T+KRqnuYeQ6mr9S0BUPvM7vYk9sI07rtquKUSN+A4zvJ
RSwok1P3HVfi5cBkaVz2GdyEZGVUe6Wjw54ykNYHRpk4luum12vESXs5lFhK2ty7
Lqys0/Hzc6pNrgOJLCF9b3tGJjIeOmloULVYChqT95/hzucquK4bxW2flEL+ZzPI
T8urmiFQ7w+P8GzOLFQ5oi+NAGAY4xkE28KqmqriO9fHjoYzJ2Wsl0tyF30WZE5+
cl2P/Djo/oJ9MHiWYzLGg7P3i84Rx0Vk92usANkBBhOuQyIu7a4Zvw3JworEg/gM
ItHkYUFdul/6tp8aALJl/WdH3caCSjOZFWb3ZLoLDLnQWetUKquo2vB4cIbK/veb
k0/zLdsMclqxUzBDnosFd/WTWqsHuYorVzrzQ9DRysnydYXBUuMioATaEhg+6ptJ
a9AoQ79FWlEgcflKCVmwK/98sqe7YhkBJMu6zrTbjEj5nmFFYDV85N0sYoTI7PJX
NSfHB9moVZtmQQ/BCGp+O7dnen7tuzM4slWUErAovU+tSxxLwrDwfj4yQVF23zoH
7js4yNlAG1/NWtC4qdRAHcvNIivto4PosWgMSo/N5RqbHYoTzpJnqE86vWa+N1mB
uhwqlyLu9idVNQNZbi91dNX4denFrXtf8tE1J7CYlBRjULJjDS2Z+fHmtAkYbIxo
RrhVxcs4GUVbZdRd4M4pCWur+kgOdPSSiK5oBIBsnIBzhurHYBSYtGE7H4HGYYwo
SdaS9N4AOTee9n5wibaH9GDYh3H0iSuxVCPNiU6bmLdLxRukeoM804m9lZAnHyXU
pXG8iyB4FknXP/iyfMueqWfs1E5GDYrGo7Sr2UKZb01kW1gsPcF5U8MBYPKi/fHr
C1guMTBZFwBqKsqEeBBac5nuqH2xAB8mVn76O3H487A/ucqq+7G7KX9+GS0fPs3q
By43lozPq+NEUuYgUiEYbGsnV19fSAnaLCc9xz3zR+EUK01Fajlu/mSDKuLvan7L
T0bJbYvbI7Iltj61ij9WwA4uKiZ7Hv5SK9pYPqxcYzXczHuBq+SOWWM9484PLSCS
h+abpJuCm2Z8CCUsGtSoR0Hg3AQF7u+hRIeXGgHBZYbok23n3UWImR5/hUNlSSOi
2ur3DmgwPB+wUuOrWoF8yW1t9rKlC7vCMcN9AlDSFrq9qUjS8B8vR5gx9tGwYI6Q
7shn7bIsXQ0wgoWdRlkaprISSdi4eADRmJpwdEElW5wCGqOdImYB3DOCU0nYnKpK
TicornXVOv+zoNDiIdRbrvXU1I6RWymZ8Lwp7mAumkbgTPCiSnaQ+lO44KaI2LpU
DHGl/e4Z69S6gFe5/7Mz9CbcaL334/IPBL8i4yed+QQ11c2dnnHn8mCt4f7i0pdg
lAlFQJfaCsGRvxXV0RPnLhHMw6RZ/xR8Jl9lTrFvolL+DzRAidrkUk3FDECeanIa
y7nLXRnm7yBsxiGe/AqFv+AeLDN0+M7b+lSydcf0Mo8hOYNJoubsvSnqyco16arN
uWe2ByJwL+firp4A5LbHmdtEU8JxqDHHFdfVEQI9gv7eXBRv9ji/9vpnsYca7wAO
Zf/NdkGUvKz04pFxIrqVhS692wwG7cdxFTqPVa3ygbmqyQYGzFbnMgbBUWCK+2hx
J/YMnaAMzQpARQ3d9Gr546+vnoWYIIYqnnd6wuIWpjuqBgrCKsY2oXE17w05ndB2
qa7vuloeRcY6wY0pY2I0LS1uVFmZS0PyCerejVLFhqMNNqg8ym1BOr6oSZoKVuHe
x562KKXbF9R2KO9qQ1Rpu2Kq9Zi+pBJHWFGjYw8xzq7VvukOSnAxKVoQs5Wj1/1a
4gNcgy2m9Or+Ott/F3BFTbvwhlbVvZ4Ll5eWdpasHTXh+jgATWi5rQeT0YESieqA
SM2AXTBSVSQV39s/2WEVt2158dF8Vy5665eM9yE3NJURRGvLn1TSFkRv6wMAmoeo
8fbm7M1RRIBbalKNyi58pNFH0wQkPOrD+N+i6lnHuCYnLqvY2lvBaIwzzWgNQGgX
73+w4IKk8WTTOeSPJBFn4hAAqZjsiqdE/tp+tIwncTltGb2bWehlV7TqZU4PI0JG
WOwNM8sWxZPmwQPpQbF+isuLq6cbR+LLk6jX0dzrHZzYp9jtWaNUbZ+B3T85aL1s
48zJ9c/69gXpxHlWleHSa8DTEFqwGKxZNXmDUlHTM6sSm+rzzEG2WfW8u1WrEZ6O
8IYaLtywVfuxAfLfWeeVFKwQrW2CDyP+b7/cNRpA6hdA8QDbDwLzy0xcyYwd3Xwz
com1VvNp5DgbiZUmK974V8rwb0/ajGh75zwxak/BbOEQn1il2EKf57NtXvonrFlr
zPfwPv2skdIUL1XKiqtq169zxZvXrdngq3g6+bwUkmG1HJcDQ8Xb7OoX52WICLdp
q6cKOvDOrIIhIK4VrRhCNwjyJcEZYQvvS7wgcePNuo6szqWdo20ls6wBhktpoUBX
ZVdBb0j84QfoINgpL0NgclT9mv5HouWv6GFug7UsxVSEOceI5hD2WhNKAQF2OFf8
YQ/7pmnY9TTlvua5cwPlctcCm9N84eZVGjYk8sw60NU23UaQMo1RUJIy0CdcV8ZH
xLyNcZv9bkuFilErHMQcXXZ+rqYbDji4OWqyDtcCO3EC+XVYzNfQnuETW11Mnwwa
KjyxAUES69d4chwP8DhTnstJLWFP6fESHk/+BqI29bfEJ9+5eLGHZ/H84aHK+vmi
aGQm6/+1xEmtXftyiqDXC3WBO0FwjfBqY73sMZSlMvOzavBqHJHLscLiZK43ZnDU
VyyHc/WT/Kt3977QZEyFu0z5t4pnwXcgItG0AxB2PGixwNdpSbdlhmV6J+4IJ3ek
c+SPHsU1ZGiz7Vlu2R1DHBPnIvt2s4iRzDk2tLTBRRPGb4InoZZkOx9wGvFo03AC
gUwCQuduquYg5uP3B04VdIg2t9zhZAw6mSmsRLkuAMQUjRCWP3OMyNlY6qHZ4iDF
rchSOYXzFrb2euQ+d3xAY2HDsG3a6ajWAWNu+msDh+zGwZ6LL5gQDRXzFbh3fKXp
ocwjSLO20Lq8nEjZmv2QwcWNnuAPVndcCr8EAy8Bw1xMMY7hDVZJbZ/hJ+1MVzEZ
WoyTFkcEXfVEtI4eL9cHHBBv7rIod9O0cEIjR++Qu1NzHQc8AN2UN2BsYOVDN+vS
hJkIKAzbfQC2Sga5OmQ0RC+PLrz3Em8dDAxQ1C+HDgxtBFRRK8qvCxqwlvhJx9M/
P8aZIFAel41fI+6J3rJdQg9PVxMRRE/m7/TZtYTYjWDbu3iv4RvckfL8tLvCs/Pe
eM5o8RA6PSRz4kNvluQ7dJUMBTPJmxyhtoHz0Y04PyBJkvTHST5KoQ+QVmrkWVSa
H7oJT27SWCDloB1PHA8txMmbpZut0gwOqlUH/vm0UeYOzpI07E2kNccSMY/ht5we
2oX+V9dmjoP9NmE2EBnqFK2ILtZQwascZU9bpj1oN/G0PFecvIGBpZCpQU+XAPAn
qCfKK5zmUUnMieewPAN7WIC3Md6bfqxWiHRrV9ISTBobJFRhe58UC/IIrs5H+YOF
1ax5X9Gv+eU1S877+oWN3N94jWshZhbeiqEUPsBwS9RrTF307SoZFB9MJk5dBVv4
rFYGb316WthH5yP+704vCpqZArf7udAGIfqE04XcpqUBhSQ+v8GDeQoUSb5EwXLt
77dtSAPUzE0A1dGhIkqkL/mmlQbiqh7+H9pS6SU7tF1b78wWR6xMKNz64GBfIIe+
XXMIhUIgFy2GCsklp6K7NqT8hFexkfYHAcEID9Mg6NZt+JAabrVMr5qxv3sM05hF
K8CR4IH/cM7cQjebozGppEOcQ9kphAl+71e39Vr77VmSeroRiDDg1rQSbOrgHa0H
tqO4qNPqNMjW1MTYST+JTPZAJWa2QaKzO9aSZs4MiqNJgmvI5C0J2hpeIczfU2VZ
JNNYAYugt/9r1N7X2yBTJdz5F6xnzXXClgGAVs1hz4v4AFQLyF6HGMv911juxVEu
R5wWMN1L3/LyoFNePSGbvIOpR+HHHqiZFfERVgZIoJ9axrMy6N0XB6KAW5cQqCAs
VEeyBlJGzg8UdGukXE8MGzVrH79mNmv8ztiqkpGlI2Bov/8gYxeSkvB/jNltHXPI
kHdJZvyd8l0NaANUqH2UmeWIpm8rPC87KUmx+S1kvid4gEhGeKtGSDrD0VVXXazf
NjG74Wnxad1Boq26l1uKfjsnY0fNkhCQeYwpuFN1li0=
`protect END_PROTECTED
