`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MYlr3Wb1af43W73QR1c34KoulMPKpuTfhYKtJNoPKUvfCA75RzpfVy3CHx5IklQy
fRnk7PDBxFzSDBg6RlWhfn5xK5CT9dB73zXZUm+WwZ3i66zVauCghs/PQfonojj1
Qb0LOiN/0knX0z42tw8/t0IqaEsBk5kNM+cjzRURKRJ/3tRMqCL2fgIlEnYWl0ls
FbyITFxxg0N6SQJV5Omms2Ns1JYIBSr2emjuoKyF2caL+bgDM9F69aQRwoRnEoMg
uJqF/bC6qRiYrx1bYl1cfuG3etydl/jkBUSSFuRZfyjecvw049Y7VGgyJkF71usN
2t/5SKYvaToK5X11sBmi1e9z1b3fOeGi+mTJs7lCOSfdoWdR63ncuWOSB6y++iLT
EztWycCAnRSohwzkI+DbJ6o0oc1aP3tqMrLCI1gn0BKbH0MG33zxIllxxe6+2yXN
wns7MabZAmAIDixc074s9pI0zNAUOJLENFFJY0w2tFfdwQC++czGu5SDkgoE3V56
qIokzDgf++yLCcO7Sc1An9UfwgtzyOqxonj9M6haWifrbp4zz5sukOt8SivFvPss
bNMViVh7jrmhkqmL9i8kJSJJ0vlwVuReHfZs2LqcVNGGl744bHNmGRylRW28plpe
Wfc6eKLTLB+xqJsmhOa9DQbb4mMf/OcI6Oe/tE8z7/RcFTelCkcNtlHGMBFn4hUi
FYyKO8o18/QSRIarU5gYiO31mBpd4Q7miIG3/xQUVXgoJvc+Ag2r6mklWvgtqB7d
dD15u5fUECugb5aa9XoADwjLH6VITTryHqeN8SHoiT1xlwFfTXFAAGdMDGoMBMN5
dfBqhW/o7jxBkZ9+nbQ9roABEdPC7atWbbJ4LRuCloLyyrjFahJMdwm2IN0XdEKg
ArGoicY92ZKf5WykW0O55PfmahGee5iW3nK20hliLxoh0zUolUN/94Q9z7hBpq4b
pYMt6GZIXavYDBEHgP5QgcshHEFHHW5VMH8/Ai5AwO0BqLDb3YCeqKgjSQ3eRes6
V3wIKWggP1gjtOMde/p93CXpr8xL2KGdlSkVDcwFDzEmR6PMKeCVHsTfRyrjd+m8
ITYXGqyufYJzH3/cc4Kw9j23/hYj09LgprZdtrV89SpolDVNkir9UWR9HXhsNil7
zJLCRr1f051WZb2dJUsBGj3IkGzk/bWIRXdg867Jhw9mzUSUeMf2Tujn/lZCJ//M
x3K3l1T9hAke5++YWddOzvN+PeN/4V4dKn7IQCukIikbw+grToJh9eGiX8n/FduG
3W0b0ZrVJDcluS3OC8G9QvSeWB8Aujo3qc3+1EiVks7rGCBpQlCuNiz4avBxSJo5
UAB9X6q7vVlZ9Y+7oJPM0q658H5HdwrY3iIZPyg0HYs=
`protect END_PROTECTED
