`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o/5z53WOtJ3qPSlmHqemIFxHt48RKCx9Nhqdz/WV5g2pzwHz3q2OVyzQQ0Lqgzbd
jsQZH3lWxvonJzSaUPhY3iKlTj4sHkjV4HJEzIuDm3VlYAIYxWTcpPL+SxUH7Z07
nhG7liA4nfSeKskg+Ms/49d2lTUFbXuIMEvhb0ZT0XI9ZwKLe7vwEbiaRCTUNyT0
WUOS5KTxOKT+sQ+8uA5ujVY6INKc4e8bxE8J3zDX6wtBM2DwkQzioa0jfcyM1X/r
n+CpwGP1Vmw8nwWMMWiceIdDsGWC2z+9gkAee/8zXebCfpjnina6jC6cQcGJvbPY
7/Y1gBedwYtt6bIBkg6Esw==
`protect END_PROTECTED
