`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q8/SH53IoU96c6yndUNMMxhVRtY6RXVZcQ84hWhRO7S0MZw6sfeel2mlW2StkM3k
Hr1WJhv1xcn/NxZVah5uvD6/zWUVrOtT4/LQESjKln2C1dAsBRCFecvVT6T+bGug
lGKgQWP93GAv1bHWAIHZeOoJs7XwU/Lvo+ifynMt0vjtwCrY2P8FGtcoWEg5Uo7T
pOSA4OKVcU6kjZ3sxsTdzhEV/+7Z+9/DeaCvdawClqEHJ311JdrUo5bkebTqIbXU
3GC5axFYo+4uJGZIb9sfbcLWDgotovvcBKEvO3haHzmkc8axumU8dwpD/K5mJzUE
zNU/CjcGO6T89RUddYI4IjQnP5m36wORW+N4s3lS7AcwaMR/WNG3XtRs8hNXdGGn
l/bDnrhNf5Se5Ow4KlBqfmrTEFLMph3T6FaIbeYywlRYVGvN/GjzmUvKzejvPPFY
bPMVILi71bVOXRWugFOZJEf+dGbDTy50VcI+1gklOBYyUB1V5LXLWRNgASn5FQ4D
/bXB9gz7PLH5hkJqsvUYow==
`protect END_PROTECTED
