`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Bm0NugP0ygWJ6NXuls/HxHR/z7IUGMK0AneekOe6uESDETJSdSOBCs7XNwKqZOa
Ef05+gqcAIq9oH7ia5Hk77w8uQ+umJ1ro0QfQE2hY9G86QWDLOIuw3ljWGIF1CIr
jeJBSZaH+yT7/O8a4hs7+u6elI2VMU1gIDVrJYEsXYoPfUpeRzZ8/dmloyzt1WHe
t0V/xDXExp/mwNWF/b2KZqpXLmoJaM6P2051Qt3SYnF3sJdVgYQs93zUyNbi4NwG
1/D0fBdz9Eit545R30Kvua/iiiUfPpMqJlaGVnmwJKe0l9k/kYafOAqXRNtv59SB
ieasYxfkBG0RAKfOGRIhrVVWXcja5dx3CZimCh99tZt10k/CApqCdTnYVyQAXdzs
YEnaMtVEctJ+Jq+ZfaQowMBWGra6iiiKEo9YJtZdiaReN4UeJX4Rwba1h/AlRBE5
eOBQ2dXG8ub24ZN5PU9yOu2IUeZGOLHhEvPCVc/9WWUeOjl2umkcXN4p1t5fn6sP
nsEQl1y+FLQNOIJTYh+z3laK/NGtsYOBuvd3ajX+LDjmRd1j81a+l/lhyvLk+f7l
sUAasQ5yTzsUJEz1tIwJksEtfg4SttP7d4goYj/8/sqolxU/tPXnNs81Bka8iFiL
+M7piq5pAcyixOszzu01eSS/aOIWg1aZ9xWq0uA8GyVcAr4+s9lhHk4jztj1PsXP
WrHrbFU79w2AjcVv91CIWBhd8670+dogV+7Yu4Nwrp9qpPGC3hJ7IxvCCDRvsGuq
gryRCmAXWNtf4NXifMxeLswawcAQS95AqvXeOBTZlxtrC+izSd4qc4oH0H+P6sIA
H1vCcPPmr2J50xNr/HNsY3l9mHTEEe4DiIqSB+JZI5jQkMlip7jr44SbamcIvHV+
MYGQNYaSRKusjAQ9TVxISoZJLvJ5XX3Q66HsibL26uncKvS0ROf46MpBBafiKHj5
hxyJQMo5uYI4NXIYgEIs4EA+H0GlZmHCUDX7+gAWNHj/ldbiCK0BsDRKuRcXKlG+
nr2qgDf8jJs7g51XCW/H1dvnM1iOnZLR7Nb1jejFpHUNDt7kTJNrR3WIR/LuUV+a
h7qX934UTRkcbvSsDxla2KVCEI2LYnxx01jQIEY2dHDfaWtr6CzzdK/vLIIfocwY
`protect END_PROTECTED
