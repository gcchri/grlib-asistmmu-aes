`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MZeBAwqi3HkMAGhbOIy8HyafkqFMXMv68Uo1ABgfg4xnzLQxYMgWIWBaUR5YQmjZ
eymZCMqtcN6K4BYsbCGgtC/xFEcSOPAgcPZqGvKj5ItvnKlqhgMg8DhuMdTcUyfd
mRIXvowKBzVsW/ETJipLDoCG8NZPMLAQL2FVBjd0pfNnb0JBK0ciSikEP7SL2zPq
IqZiXimlYqUsErrZBaz5eYBXGmWClJLrzi68aL3iwfCpggCSslqhj1XFq9YKh/kL
2NRA39ITBQxx9/1pb4A9GN0tn2UAz0inG+N6l2BNEySV/FXBqCVAAxOS+theG043
XbLvxrtElSu+hcvJ9STCbBN/MeDaN8Tz72ZyQHE9NtAIH/PPUYcXMKX6bXLIt0V/
63/9zGV9xn6X+XX4dgBZ11zel38FZBOxdFRlIuq7k6KlJA8Rfklnz+OXKpYPZ2jC
`protect END_PROTECTED
