`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OT1AVZb1io5FZL0xCQtumuWSYQPbuLWJXnoOSQvS3wTqiOkqxUTG1S5WObjdupOV
IjaXjW9taaig+FCU82wNUlMEo9UcMMvtn4X60y+gyO10SlEHrIslhpJKYj9+RZMk
HGorbrgnEebQfkRVtYOKuRlW4lZQCm5RrJLjRV3dlMf/O6CCZNSL6ar1EZL/GFvi
DiF7WBwJj2Euc6y22N7KQYOtLOMiPN4s7omWRiAJ++XMzTmVFApYSkhHhndWz/Dx
su6z+ZaRLMDcB7GXZrBb7s1MWUPjsdhzJrs+v+ec5V97+jQTVpn+pK6bbYnhUEkF
F+oNS0KB1KJNVRHcRn1vveNtqj+rHwb/PtR1Y+U+UpvUkMq2CmNmi1pARgd5ESrD
1v8YpYTRd1HeMVAE72dCLrveiENIIkGzFrVllOjFC6o=
`protect END_PROTECTED
