`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cxo+qsYvqxxA9ag3TKWB+dOG+fU44lR23BI1ys+/sHNceV1JckjP9V7LM7Y34+sc
9LLddwXEJjsj1YdWzzwkN216ocNaO7ex10tLBwKQzPgvFEsa4zU+KzNWpVLgDGrL
RbilkasE5Aq4uODZvPpddp89im0Pec6q3+Vt+Vratwc1tMmRDioJqOd7cxCT3yVk
ONWXocGbz6FlYzA1RVNYXDDcKSdblyfPD5QaoBf78+cOvLYlWAabWKyj/1VEMxzC
oy4qIXGA+J+o2FMUHr0DHhhmKwdMNHRCOo0LXZSlk8SVRK8CNkNrKxYBNqMvORFn
LRu4cZmTyIJe0sVJPynR/rp/dNrOOoTKuoLFfVqRcU0mrcuvEEyr5rBhnAtMtlmQ
Njl8jhppWXhsAbteiZASEGQX7w4MJfJwQJFVsRxFUbGiLkOLT3ZCq2EW99zgNNS4
G5ylEPEQ/cuQ9KHPtLCygEksUEyiCGenWvAm//bFPm0TyyqGemhp2I1nDsdGEgiG
etdgtIVF5PPBlkPT5dJLVu+SrjsVdg3a8TVj/xyt7vidqy/ojy44G+D/B6ZwGaHE
nzrfKXZ5y8GrUnYLhuks+BUYtFTxa165IcVDQ0vgHC7Kiao2yP4DlatIbAhcwOrh
TOo3krJ58JWT5Hq519+p3QuMvAa8CrA6zYsvr7njdvYyEX0vXDbyAoHL9lvjRiio
4C19PP98d/q2Xt5yIYUz6pkEewk43prpBg9Zmzmmzc4pPfLufPDv4D5B7jd7oFFC
zaLiFPHgv9jjOK70Hr/gnM+QakzTwhNdZ9di6grDn5AITXaFVa+H7eVQAcHsghKU
77yMQp4QwM3ypjUVc+BBU2bKb0AwfA/PyjC8nCp+S8X6r8URgM4s9YlRs5KTgQw0
3iteffWwoRY4i2RKF+CBzBtolr8YzrCLx7x8V6LVdr/veNqPfJ1x/ZKRP2MUt+/D
pORHZ3TTc7AOptkLROge6qCi2Mo37yxJVBMWxh703T3ftgLv71um31IMyH7MuXGl
emfhepRQkRiTsT0b+LE3ZFjpMOQ8QHNYlejhYiq3psLqThecZ1m9HJqMh0x2Wpoj
Oq3hRSczi6tzQcrVXFlx26X8jz8Z9rNx4K7m5EB7TPzdH6Vz3nwWkHmWEJaIU4j7
`protect END_PROTECTED
