`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KVGAnc22QrTo8SQ0N0OjoP+WUo8yMRCIePo4c3n9Vo+ZCfylBBoX6yODbrF1+vRk
q/In7c8IU32EwrtyyrpqrOI65rHTgbScbmmssAUnYiAOJTrOhjvETWd77DKA30Gx
g71hbML7sJep0WhJC2Ts69lpaOb2oJD6h+y08eSYEQ5woCvzEdBgd95gGlD/Hn8D
JbnbM/5U5y9ImdNuSg/S2BFFf7xVAg6s9oM7C1b0GFYbjr//lFnhI/lmxkPCniet
bicf92gd9FJwkr2cHV+0EPih1sAWbimaooRru54HQsS9mgatozf4AKD8t49RxcgN
SdYtK4twElb09XbGRYei60Bpakkow825LNsEdzBOro1OTwLRA4nphwGvL+Kpt8Qc
lzVaKUY1B8gH5NuPKT9/wGgk0j3IsZJGJ+it+JfdC0uEqUeMF4fcK2NppJZZH9TF
SOlFeVC7odO8i4UGVE09ouevqz7GHyEGKq97PRkyJb9y+mZn3TInexbF59NlVP5v
fO+CxOpsWlFJio7REl7L5/ykxLhvR0craYs3RqBkpIA7FV0iiZPTJORz4ghzJ0eS
OPxUSM0YiDM5/l6G466lKA==
`protect END_PROTECTED
