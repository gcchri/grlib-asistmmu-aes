`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DAL05nOdkBcoSqjAlJIhQYfjyQNNwwbPgwxL7AX2LjxP8lb4/eKUtR5W7wr1eDCA
AM8/2NvVlZFvvZBm3WWwuviWAzX8B3ggLOdSCEM/Pv4M6xIt4S/skFsNsL8Kxy24
NO+gbRRVdmbbXqlF5Jf79COqIFRmZjrdt1XneB4nNUxCT8DxcouhIsHRoh6tYelS
B5pDErlcleZoqNP7fsgTENT5dQH4+R+RCYEzW9qJpMSg3UKalLeWai4JqANMQSUk
Qd3Is4H3mdbcuV4/1Q8XqiFImLApkKC/bIQHGhfxW19J/IK8K0zAsWS+P1UGl0Lj
oLTO86D82PMCcsFwBnssoVKjlMxxLEBTecRJn+bOnfcWTAxjPft9sqWtT0W03r+C
qllIYT63dx326F+fbOpLJWIav5stCtk6zTW4xSC4TRY=
`protect END_PROTECTED
