`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wKSyXa5CnTX12y6Gl27Vm/pc8vIvADSpxpNj5f5/2w0Ww9n2UgJUWjGcSbrq6OCA
Zqqnmg8q9NOC26saf4GTqO5sHqfxOiwntK43b7HNvkGVNJhJ583lVRj+D/gBQhzD
RgCZoNvXYF1Z8fGemSsqc4U3dhZcJEp9bp/PRQRUZxDxvoi8vC/eyiWm0cI0ka6V
BLx/zJju9jgfu5bvg5sDlWYJvZwmQ3HFI2rMgYb7zljpkgwGlO04zWCQ0gfkG0BE
hviE7B4SRFwzQhxzQnxiDGy73EP7L6e1DydaEovCigZmBsUEMphpn7k6WFcVqhWP
uPEtmOZzGTNYGWBxUWIlZg==
`protect END_PROTECTED
