`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XhD1fdbE5iP/DSrTJBDsCBbtZQCfv2r7iz6d8w/TEOorpwOdePrA4dYAxqjayaLz
38fNC1ho24N/vk9Eym7ITqVCLwsAQ+GMX0zAjPVymZ0F0jJXGTaKirORObnJdmCf
lTF020i2Du9JENanYPw85ekXa65FChN3PYlak2YeeJ4B3VsYU+SAtk+S+bgkQ1kb
H03Qjct9LkPJKxEEkTqET4RX9LFK5UuA6xEY71/SS+QYoI+FaKqwQ5uIANF5xuTv
SMJc2uGQTp5ut1eYE2OB5Ae/USQ45/40PkQF2le2bV1GGiGSWMQBXlk6Qt/9yzvL
amZnhiDPgHmovd2dihtXUqxaXr6nk+7Xwk4IOCD8EJQ5bXZ/JAWyEPWIy3+R8KWy
UzvqyqCu9GJS8WEjIuiQl3EscKy4a/DdaxPtPpXcTWc1ezDbEbMmDlkvSznTdnIl
4zoVH7f7hVhlYMGkM6SU7fHR43VagSfzxZELc2iLljYwRrEHIvTqfxB/pXeClahf
KWlQmWcQ3+tU1yekGrwdYiS1076Di6BzED22Y1cl/olzYQS0jEyRoj4wxtuVor+K
TdcEfkE84WDSGba/JFLwifwK1SDaXsx0xM7ic80v3dqSWnpdvlkoG7TwKqBB2qjD
qj4xNxYyRiVOhF3xrGoIKSYAuMZaxAS7NdQsA++P5numDNC2WOlzKxydL2dfAxVv
D3qz0w2j8J7xkRJeckVjipjivIPwWhDtRNsT632Ad4qPyH4SgVrO2/xTkxppnXUk
HH8PRbtJ1fYeiZLEfJX3HeWZYSjJ3ODvb7jJ4ywC8RdPtIOtTy4ihnl8+bIwVAL8
XbWvzqEKGjNVeRONMO0WbwSISll9uCn7xuc4+vW6B/6tfZ4WX7ZQ9Z7ySlrN2IUc
UG8Yr2jIEBkY7gPfCubmRo+6dRyGvXF5JKywC+tC1rATT9XO0Mip6Zh7tM7r4TQF
6WRu+8nQrHZP1AAMWc8bretUqPgvLRz0bEhnSdOZF4M/aupj2C8UOWcgJq3j8g29
qPNati5KB7fAzaHkg7+ypEf9lnKf8n1zE1m/da67mVmtepVbDtA9vSqcEdNWk5xH
RMVsh+f9gjeO570C9q6vvcL9Eb2ZbMSUQkoGKU3QwQWJi/stD4vudQp0vuUQYOwj
YE9uNx3houOHH0QdChwsgu4gXhQ3sDKCw5Si9hkeNOqnhKc10adrh5GMA8rdt5n+
CLA8StEPdnx0G+TTEaX5Ld0CIkgrbrdHyDgfQPmXna6pR+gssWg4D05k/ntMbAEp
FbaJ/702y0FYFB1mKYpHnMxElXYf9HcOYXMkQ+/nT6xRyj9oYBnk/h6jV9+5oWpx
/w1Rjzi8Wrk3pdFkH3/V3xNrlAZWHOIRXe6S3PGi4gWWTeveAsShjWT5r6jDKAWR
LJ+MWFOZg8suvFU2Ch5R85acvGkEi2AyZvcM4cM9UaB4RIU8vluwj4lFqKDKuRzE
Tt/7ubq1lRnbBvRQVOk7S70AoqSyKGgbJa+zCMrAYeyOf/fDmYUANKiS3rQCJRE5
n9/ew2AkQXi2oZo5WSmN9iXxxb4BUWi9snaKApJSCgZpXtMgYpabXCrqC7m1OH6F
npOugkFfuu/Njg5XQhsF3FdpPvhS6Nk2gfZvMCLparoeuyu6EWSYS2Xipz3z3Z8U
1YFX5Z6lPhBWL6zE17jxJTMdVLdJI8D1JUtdsP4WsBv8E3QMxDCCbkMqwi9Nc8EF
4MG6W8l6Q5xMaGR97MCLk3a2+JO3qbNje/zrtZytSoT9hbwARNWw9cCSfp69ziYq
uQbP9xWbpkOQ9u1FSXAEGT1KKmmpq9bMv2czTKVuvrg=
`protect END_PROTECTED
