`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MJVlX6lV7hLoHdV5R8nYZyMJVTvam1BL29tf1k+zK3n9ggcsZ9m6J/3bO17xqwiY
dpw/XtbuxoRv9mAhOB1cqhj7ZsoetvpllwrH/RDJkFnAyir06g87x34UcdZEkqsP
7IllmIgYKNtMke116LdG1/ejervs4R2a4+Vfcv+I5N3gLr1dwq5wd6gJBSaGdhH1
IM9+zAdJvvLhqv/Em0pmIoeT5ofDpdofJUBdeCaEyahjKl5SL/8C8icstepEfoJu
QPEXRnptCouKWuCcfmWHGYyx/5CFrZ2sZUw6YgIEewCOpMSpOy9B/PIS4GFKWNPZ
4j8+sXPrh9zRU3WVtR6lwtu1rXiW3Dta/JR63MVrQvNsfoERdmsIYP73b1QBu9Ss
V+2zhEg8UiwYk0Rb7L8F0g==
`protect END_PROTECTED
