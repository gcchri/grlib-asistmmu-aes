`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
agvrVQehMvPRJpq1mifFkXTeAfGUylujEZNaLtUB9U9v6151onx/rLjcDrdG967L
MVL0pgck1e+9MZbWMBjmgiHx37Sxo7goJJXfuLdAoAObpj7YLM5aeRHLBaQDJF3s
bFENJxsocioZv1/nn9VxmlgDxHoAY6ZsKPlJi6G37dJt+Vn/Adnx/gHgfoqXQ74e
rkCXvxq0lBGcVbJV8nHxaN3U3HkE1XrkuhhqLNhI7ZilxeklLaOgobWlNGrhls2x
VsqUYBf671WP4YMFYPsnFSY3d1WkbltnhWkxcQHHOYHaoBOVGO3iwZUUHy2UzE/a
Djf5ssOzdkq6OOF9/jt6S3yWb+5FLwhaqFNV58KMGILuQQw0J5mAPe0OWOFj8HvF
hFY3JXxJjn24mNpBJDAcjV6wOJlA+nXcV1kiRW6kgyY=
`protect END_PROTECTED
