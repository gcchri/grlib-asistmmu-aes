`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kS2U2cTbSiDuSZNlzMMiHTlotI+/B6hHqBYmFHTuF75qXWkDNtaPHfZgoRvy7RUn
Ze4o5I6tZ+vDnCwRnjmjpQGrmtSPHF+Hgotap7GsDWnhSIqjQv7TOmf4Sj9U69cy
wxB2SYbDBSNJx0sDA4enmE21ntY0Mb45aNGb4rwVTIXMakMjZIiKmg75ZXiokDKh
J0ZIctu01qdeTR3ebr+g/CD5SW/NmDwXUmsjkJyCWomwkcF3r9byInNS0Pa9AESH
D9vu+SA5qussHwCCV52e7WifYmdKRD0AKpmbCFuWWJh5mHNPb9AJLL3HCyk2o9nm
mgWUbHtvNLA6U6K0UMQX2Me5lx0WSSjDyu91SHlk2JXrvm0EExxHwyyKhWeroYvQ
6XzhdlsRw7p92lPMw1gt6Abv24bAPKFIGEDbYo4+x5Ly86jIrYpjcOtoOT+DqX3D
V4Gx9dAXnkTtDrmq/x1xe3RHcYioeO2FcAsn+r2qHcDQIG7DgBL8zIHkw9idfVo0
K6X9RquA32Q8yZ6/3vrlavt5YaWzhI8ryx2luJHUMVDXxgJGyvqxKAgqGJGKOE0y
AkHhb1i9bZ7boeGvYh7TJXHyL/ukDucazZVtpFXPDE/9uMOTdfvh3QpiuAMJpECk
g8ypUCLCJhrlfOebDm/Jq0fnEGWkltvopHEJXVvsv4WngmADbxGCoJ6eGpGI/YSU
WSOKL6B7aQFMmpC70VWeyQUmgul5SnjDwolZEcwtPEmGIsh4rTsisWs+V0nBxeHX
9ClBUc0tgMP106IpTzb3K7gPbQwmH1uEgdEosmtJLjy54TrGGo5ApgnBuCkOdPII
u5Scn+YTq9rgV04XjpcUKQAUVKy5qa9xzNZSX6YLrsQSuLUbXmr9MYn2k3ocW/bD
yTGazOhHgNhyVLbFfEIBEaQ2FZ66ou6koojIHw7ib7KUIFiIc3nabTPZUo6iKpqo
FYejDEAN4otTYoydxy/uNssjGCnyIPdLcaGmbUbssADoSNnY0qz2ZCocldKCDFgA
9WXyMYJ/jtanxGPIYEGwGQ==
`protect END_PROTECTED
