`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K1ToPrJvoBNjySe+t5ak9OmgwDeRNaV6gHwffZUeWl0AWouWsm1sSJStN+2LogHw
sOr7fzr+YhRpoJuTml3aCXEKkBJGM5owdSg0ZOYK+7216YzcyiKMkJYEldUb4bGa
bxzz6nsCt2s20bOoQerYVHmlYZBKltxirru3CkGHL2dy0UTRBT9p3QvdHQp3VaN0
1b2Xo2i0gNWd1/FYSIS1DMJFGjgTyoI+9xYw3Bwg6ZmaKzUFU3JlHXnFVZQyIIVI
cFf13GEx0dGYwEEFmddXEMJ0XYlb3QpwgXRndnTzzCxS14ydEn+J1H/sn8b3Ao4h
kWY9gbGUikKdGndMNEAN0cL/uO6z4AwHQd9kEL9Ra6zy44gQIOOCbl/F4UCFBIHB
4rfms5Nvw7XDrNLHcAEvCDvxIOXj9KhpAwzkYlh6k/ay8bBPc+zAZSpVRaMof/fC
Z93Wj8E7GEW+fSCdvVOilyKIVwKPt4DLYjTDVg5UGTpzHjdraVA6ZnFFSAQuCd/Y
is6fp1uRYXCHtJ5AHWKNsnI7NGhEc1PMmukzAOmxzwA9qCR9Jq5p5LPw0a/JJwQm
`protect END_PROTECTED
