`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KGjuhxuqY+bw9NWLo6z/DaecobRP0g0YqtBAeq4ZEqSmQgkMhdUlVncIzxHDuv1f
ZT7QPTMx4uksujRsOEM5aGLuFRZRn0QXLJksyEkfYeQXKA8S2OxydSQOszYgwdmY
HO0/9ihtnAVJ1a5l634nZyGaXBfgGaHKpOla44WFGSTpesbrPIZhyXFd9xSrxdIr
F4iR+Xqe/Y/mYuJDa4hwtRrnlEBwDUZ6gRR4OIWspeXgt1k0Q9ei5lJOwb4hr/7o
h4YC1z57Zrdd0MJQuR2DDJr0Gq93aun8n3VJZlPrYtCMCcRKXYLbvXTjf1V7GldN
`protect END_PROTECTED
