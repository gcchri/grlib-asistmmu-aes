`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kJtxYVQZ+tu1qnTwsU5yeAuLbeZ/ce/bBPr4La1vRcbECT8EJcxqVeIgXSF6qimA
69QW5hfuUM7STxQMUuDpubOaNCAqBGPSelVy5oD5R6PzIhbublfxs16fMaMY4za2
qH51EnVdYfszMEZADf+09iznLc2UGTsq0y7e8XU9ldY8wTtuPzJOKNhebbCVU38z
q+sy1WjS4+c/ibLVSEgX2+BDRqKa1hKgD5846+cMq63U7i1Cs6kh7ZnnPpYwlDVV
OOHZNv5Pk4cKw60K51SuyheJbJfVMENC67EwqwsGyvavZAiDl+ohzu+qAKCnwUC/
Ez9sW5Ohv9Rzp/jq82NLU2h6mWapK0IfkGudy0OL6mgrS+BThjgAoWLfJROgoT39
sRF7I4oKvnNi974Vj9mD0iIJtMNyvkJQs01MqHOtreMksFOl4TtdfzX25KPYH2og
ZY94SHCJw2bPVxf5mowEMcNOLLUAzXsnbzCo82oqwuOW3b2Ox6c6Ltw4fN//48+v
9hMk2gAQxMQorbFCiaIrhNaXPjjYwUZVpVLVnQxFAI8/1M1iClhWqeS2SghKDDW8
FoSI3qoIyhPfs7cHperbG5reY+/MCRUBDI4cnOap4KY96tTf9jSmusHrkovNr6fI
jxHyWI8NhpMJavgUrFQ2mzbQhpS5+K5aTb7rvdjkxLwnK2FqiBMdHgWGrWsms9ba
8pQUJuaA2tNxsH4xL9ufau+gGKjRCWWms6GewPURyuNNoGp6fEFIEUmNZdokH/Jr
9a2cIV9FcdotP2v6R7JLka6C5Q/IM6jQse/xhtZGHWNuJes1R2k9sQGX1yyjAWwu
zyHGTdYEsC0I9a/m+q3sVZoYLum7bsNLcX5hWDd4xjQm3gnMjkkKVnm0zqiGHwj/
DiwTs4kOjfqDWD1PLw400UaqfJVYMTXdpcxAcVoQd0kKnIq/coc2HZWHIXgw0NWf
LYP1iXP/Q+JBHsAoGMS1HjLo65IyoohbcOxRvTr/ioS7DBS8+BKJVhAUrUFiQNmy
BQIkDIqVwBNDjp2JbGIYRU0ql35rwcmUthSeTKgGzzTTuY6O6Hl2lt0hI0/SrJXw
9vsHEIdtTsLXuXB6m53gAOfE/DjJ/MIMspUQOouxHSusfxeyAZrqk+QkyEv2aWfn
ussOh6QTYFHqwFHUV6w77y/REkQPRkZjaW8HJS12KrAv9zsph6RyfMXQgxbh/DXt
21fkEOiDEKnZb6co3+F9dPgDBcGNIaPVyWBPS3ioxieKiUxzLgao7P6kt08FQNMq
aAoyaB2UuFoAI/Vn24XG2ztJIxK6hkrkcbAU0KUInxC7Nt/v7k07ML+RfDE+W/9i
j2oqB79Iht3DggU2cuxw/oIUDNkbyK5RFtfUMO7E3FCCQ8Ik3bFdJaJ+yfeB+mUm
D/hQXJgt8eimTAck3TQuZl+HJAe1wTwabCA2kt8eB5ECBI2hGThve/SjP19zpIlo
DC1CGQWApoU5OnSYk+CghKBbBqsErrDvIIFjG2k5uiPbSJmpzw4R0/bf+qWPQnK5
+oX9m+uVFuePICL0xHMEXYWwzu57lDMIcF9EeDu5ym7oYqhmWz1cErfPyf5/+znl
`protect END_PROTECTED
