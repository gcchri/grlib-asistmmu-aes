`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jiN6XakJuxo/K1X/oBghq0DPr7RoKg9NecZ3hbPlfRECBWx3Xtuimblw6ybNowsA
2DXP1pGrBpeMYCfhvhQTT1tn7uaRl7UiSjFvi6k9FtXe18oyj7qJz57ReHFiWrel
46JVceZ7H7zob83/1JdvpkwmyJY/g02YwBJB+5fHleluPwR5gdHZXDRSih+TOFEn
JHkGvGZ2Ds6zWe8s1u6/x8KR1UpcOsikj6VvcRfLBZM/s9eG0M7pmKsoGJtEGuya
6UOVSMTEFzOyVnQVZWNHivZp9aH6bkLvds+CmGm/7WRNMe/kmZxbxTkomSJ6gVDZ
kxV7UdzX3f1NwYvF8lheQrBqHAqmKzapUHRMHCbEnpFSkG5Vmwmf302t3427N3el
ffk3vGFuSnq7A9KhQdk08Frp20zZT7yidvDbi+1vRHn9A9DaaHSL3xTwnuqDBe5Z
ipCDwm+DvdPlE8P98A1jmCqr5hB+hTv1WmwgS7/PydiESCLv8KmlgeBwqrZX+SBy
AmXIznhqKQrFy/zAEJ6nE7bbUaky1Z1FHBEp8virrm2me2WtFpu22dN3tEJsCcDd
WqZj0Z7Jl2neCdKDGYcWTOXW1VI7U/vq7m7SDmSK3xUT6c91IMlO6DgTtRl7sPwl
ZVu93TgNpaLaFL8TWq3o4Mkw3swV2bqgtq/EcuSHW4/auez8myF4pJrMXSfF6zI3
no1o2M+pj72ExbkiZ/d9zRDAVCy7TD2iMpwYv/YESKh0fmBfONyD6kbXTnqidMXC
QfWMwa7yxvUEklW6sClD1nddKgUTgj/vH2uXU5/EICQNGIvD/Sgwty7TRPEARFTT
HAN6jDRhr3pdnvKmyp4wz7n9XEXQ3UpuMPvrdQVGP1j702Zk9dU4/1jdXoRJSlgw
/kKefeAyaNZEK/q4FtuZ5ZhWlnSPqS/f/cIz6K+qL5imi+VdGk5NgtHqi+MFwnCk
6kzlSitgUUUcO34Osuu6DUEU/KoIIVPm25kSO8kHHpggGO9oUBYE/fo4efTFrrN5
sdnoHjsSZWt9ANrKTQoVG8gGwWDmDS4Tbw6skSIEzWeYtzx57g8zSv0g0/IOqrwZ
5ZaorSnKdHOgSHp/qz1gPP5vVB4fV254q4UuTQ9yDpY4n0RAF8xif57JSakoohED
WPx52IwuNudpVIRGUdb91Q0r8pPkUxpl9owyF2GxXKFGkht1+hnFL63cbavePyb1
3vrz5qfQR3kyJxH7P+X/s3TolbYijwV08meC8n5Mlr6UOg4IR9a9BXNPUqYjfP3F
IRWzl1ElTiKqPs7TaeFT0RQYoUXRD+viA0sg+XKs4KEuYFxIXjjgMte28cXNwETJ
2enL3SR5xTL+9kSc6+ke4eRhFGHtv1V8heFBjrtdC6JrHHCEta+gx6p97WrBo2gU
SWo1xth/1g13yAAdE421aDLS/fCvrwtggRLY1c4k/1A6+DxvKk1JIOisGJBG9rNx
OW5OKOFaNW8APNpWIoJGbN7OoyAef8/zE2Zd0Y4X9GkFrA3UkMO0kcVNkFJjSMY/
ceTNF/c6HD8iiw+KChzsuBQFV7q4XGQqVdGarkSSu8NmYcNpMh3mO62zb+B4dXUV
8mmS4JcWrCWgmZXyatUSdhdcTE1hZ0PgvEf7XrgRS3n2UAcrGXKU/UlTWEcjau+I
IVkZxyOLzUmYsHv1diw+aJu26ABynR3DBdRcMgiuNgPaqbNqjSS01nE/h/ubEtbO
/gkRBotOzFZ90yO9jFyXxh7UTbVLh5GCS4zEeec+sGAmV/pk5vVjhzKOmF08fvVv
gUN5leCHF/WVQq91VOVAXIg0A9VCPHHFM0x0nsTi8Z+ugSgZosQqkPSvAyd8vC1y
c5jmc+ehX+FoIkkJF5y4kukc57Nq1sirZv09Ofus76RY4tR/0SS/xGmCTfxK5RzM
6s4ccEyd+DlgQ3HqzukkEZ+MUXnGIpOufydau8YlsweDZ9Zo0dDwFcurLp5dPm7l
ON783GRCxJDcRauN1MjabZTodrdRxPZYHfrpTyO0TkUknUfZ1+e3QD7aXbX10x4G
EhonPr8OQ41+XFFj0UkYX8fo41KzjfYWjEfMUMNGWNDkBR2aYRc33YYasgM7L3DQ
zwDp3jwXuQ1o8YcIecyXTwUJLh2FpJm9FGo0Z/GX/DAM744DdrBxkBKMsW6Br42n
AuEuUEfJZpzbyRsoBURlGbCzPVgmW8gtfRLFiyqa8vwf53OaLJSpRiRNZ/wkmnZZ
aDGLMOOMDb0SdCuXTNTW/xIZ1a7Ju9BlTajB0xAdS0c25dkivK9JxxgyeIUe1Wsx
Oybazf7NWC+ks90OLqpGYRC858TnUasKO5iUtIktMQG+97LbGF0AxiKnPVtfab7/
tg5nMDHYapnhLNq+GbQMCIZ4qQlKnKq48bK3P8VpbGhTxt4poUvt2z+XDZIekWr1
xH3rvh9TITQK02GHkGESdkCHqWblkCQP0hLWoDTAjqAW1uk/5xIczV4nenAIgd8f
IbjsK8o8ueexAI6ccCyThT1IU/aB7MOYzLXLacUEO48ak/r4vXR6+5BAxrV5fOcg
wmjIJR8ikm+6AiWTbNGV6LTLcpaSca1FDDCamGaF+bFQpmu6ymk7j6Tn3XdZxwDt
KcLtw+piOqLBYTAHkUOuJt+3/i0bGMCTCyYOL/tjKzfq6JR9KCnoKSFlMqJnjWKm
Aq0O8W9Faah7dvh7UwzOAzk7yV0geeCD4Vz5GkFLo6UgcDganRidB7wwXSI4TaUl
Oafzdb0UKedP1LsAYnn9Vaeg1iSWBt+f7vhWt4Bg+uuH4kzYi1JF3olTj8Ujk1Oy
QoqIWKlXadtfltmm3VwoamtJDdxamao76XQlCx926qJaaamGzujfvxJqd0cOeCYR
1DNGedNtiG6tJnzwpPG7ugBbC6VTw41/Ar+8CDixcnvLcFFacWqiztQ4HBFcEYmb
6hoGbnsDatFp1fKWccZsEUAT7ULI7n0rCXs7ecCg0dMog9/3sE5VuYCqBNNOMrKI
IWIazM2kEeRY90c6MUZ/1k1HNHr5U2kMb8Ss5c+Gu8ULcbtrtDpCr7f8t3aGIZ4z
TXgmFUl+roO8YVitzk6vixwzqiPgqw/nL0NGjI8mWmNo4lIsI++kmG5NtrSHzXI7
mwZgZr35QY7FZmK+JxnKp0Q/YZx6nRNiJWb3xN/4pAMzqmkFeWWUvH1K1UY+B8ve
JSvUkN0M5XBkMfQxdnL/zq5e/iQq0gIxqfxB8JXMgARmJ4exbRCb4uafmJjUmTqM
ejUBX0TtNrf8NOPTk2s7JmbZZ8JmavAOZr87r/FstyuVj2Tq8t5D1g5sdSLi6Wv0
1E9ZGWLrbrnATQlrfCwM/5rrQ95bs6x4edXa2vWGNQZTx+IIjchUWVQBtoK3KFNT
Zcy3SutNWFSynV8rGoDE+mfOuNCycZPU8F6sQMiSId38JBksAmGkGv9iqAs0EdaF
zahH12MCMn5BYiWh1Mu69JSQ5ODh+7OqITnfmfxMvXusHmxZqY4VHwFsN2woSACs
z9G0uQRB9ymgcE0vozcnxk5Vh8Exsbu4sa86n1Hw2uWhVcxkj0hRwJNOV3dqeKlU
gLw9CWpfexEoZKNnAZlZYSIMi8Girx9IF+9kX0B++vBH+9mBmUpKrzuI0T59mFuY
XZ0AMQzwaCL5JeC4Zb/sZGgQlN7nKVCbuvzbbB1W5tYeYIm0fEvYqnyjPfprRlAo
iCcfE3DyBYgj/Lxdy9dHA1T6fXks2PkDJJPZanFZmSr8pIeqDclz/9TfmB5Pmiy6
ouMdgAJ4KqXKnVdYTRzTUw5cLNclsqEeS63CwdOtoRtSSDEIyz2YWaDNH9c616Jv
qI3Q068i432nDpaw/Jtsi6bCTeXeQanTRBzHV4onLsCd/9KtHc2zIrdjSmMENxn9
znvDEU8F58ULIeuX80oCJNX9faLWnaPukR0612Ngz4M3zUUEO+4MyCde6tnVgSj0
sr5Bz667rl6FlSXzoLPJoQuXR7KkZv5MR+W55yD7cMzI0DZxf1tIqv1ovY5UBwpA
FshrNwvH2Au4Q6zM/owJrbEFanDCq+Pk1bINYKMm4TAQPHpKOmifwhdBtuuzX0Zm
UDOTfwwjcvBHMLrw+ZracXZ6gSEV7VlNOcHeLbDsmjKvZfsrKR4b/ARZ+jhqYbk+
gjdL7QD54alN2mhvxTZarqnuFVvDGgBdRTqpRgs1Quzx6alaCCNzWIeeeo200F2u
usx52orE9Wbluld3ECvTnFB7qp3csYWKs8QdEG+puc1q6fhfr5DgIWuWZOXYPzLD
hGy15jwzHzrE/u5I/zYNEXIWIa0H11bABKtE+Rz75DxvUfJA7yy9TrQbBDySt3Ej
ILfd7awAxxPcIlyql5X9Ahhvofa9d37eVV8w9pb/U4+DVD5HD8+oXfGm62Vi/845
V8/GC2DMXmIHFXRmX6RXyk0KJQ3HYcxNxNpdQY/Pw77ggYWLntlp5MuYxfrBktW5
5aGOXzzVSGgdK7iW4uSwkvIFMRTaw4qazkncwiQKwruEf9n4towXFgfkbQMaM6Eo
ppfbXkrx9P/dbJu7IF7l8veXkSj52qLDReF+XZ2ijBKCVo9LtBs/+F9PCa/aceOL
isOpp1jc7u8fcBLRUGqUz/FEo8qEFEykMOCKKisT2cWmHU2xqzt/fwaeFwgNWZII
ZVr3GWyu+2mVrfmw3LH8KlYygr6mGUNqso1kC/GMAHc/aUKLURXQsk8Xx6PpucIV
EoS7/2eUYJ4p2M0xUGE2+SB018MifHKhBqdgS9aGgjYL1FjqzYwOSmVUeKEZfK51
5ntLgu1xFYazIAvPc7YrbniJOuR8RuaUEginHG5zrdXxw+sbU1S+eNdHQnEiaTyp
MFC7nmJQDmC3hA0MFh/IuuSc7GvVlg3fwsaV6LCwqNov/QRE1MeFZq71ooqwLVl4
hNkjb/voSREbHh6QJ7jwPjM+ilY3j+ow4BYldcR/4xMWqD6FJLRbEDRJ0UCRreZp
6ZnjoAISk/xpv2WXUN6GR00TDILd5LziFncbOo842E/vUtF4bPmlqcgKRQnm8nif
R66aNRTzQMAH7H3Dohn5CpOMQodoOIMWjGySliCtL/bHLiRvPDhlSl/bcO0Z55J1
VYO96A2/ilFanLlJk3FWDVmzmTrMk/rERcXZ93Tr04VqcCwEx1p5umAATA02+f/r
ysmjB+FAkbfj7B4w+0fvj9aWIfCS1r5VxI0pexUH6QKkIp9fLaQjPmz9qXNPFjES
niUjdILlOyw3LCWCLaxhn0kqmTVrTHyVhqaaMBiQ7jBfhorSr7asw9E/SIcEe2IJ
OpLCxxvD2ACQyoiwyO2T5DS/5bvDX1g4Oo4jP9hkBtclSmg2CNceh/1KpROwwAlR
1EmTG+fJjhY0yxy0pWl8K5ghnG2Z1bK3s8bWh8vQqG/xohLHKN4iFJH0Hj9V7Rfu
E2+3oYlOEEDGGWPvfHOlxiwCcUA9hssVlF+dyX00MsM8rw5DogqckqEn149/Ohcj
Xfr51u4zjiUFxwyYLnbEvyvaJ253zF0kTKUqUNmy4gsiU4lQAzRzL39wifmXdZi7
s30ImIidjQ5OIKk/O4bBrxTB+rmpAmTG7T0JQe4j0vC4PfNO+GTLYmomlg8GNpQS
mxzfemgsxAPtMDHNicwj16uTaVYTESnOvMsM8tg0xJj5vExjIe2oMKbTpFratHrT
H0EyJ9FwyB+FCglPODLHfw5t7yDXHDPc8QreFM7HblP8yKzXbeK1nVySFfiwfiHw
gNuGmwSvgTLfr0KnRgnZdvcUVtvZKgT3/6A5ISXh1UI8bfGQKMfXi3xNBFO0TKGu
j9AHy3hvOflZ2P0sa7MUp6+rPynwXI3hwnwSMXZqI1emhSWsP2E21H5Qe0QM0zMH
xK9MLrtdvQUA+PwBzGtt/6GehkPT8WOSrIdtHf9Uzw3863X4qM+zJPQpfcxqdrWb
6AIVJzb0Mt43oRZaXe3etsePf9GPbro5uR1CagHK1NRdGUbZ0MMqxFlYLhLbN5W1
J3lcYKmqeF0gFeIArC3PT5CaeWZnITbs0qmM4T3yB6O3ePlm58IUEohQY8cWuAfj
6dVxtJj+43w6T2nXi04VNxLjaGd8RCQXXes2Wtjx3ty5gotQxDqVvoovH84u0PQU
4yXpUq2pw+8k5Ww9BJJr8afDPGao/9dz+BdsUMSQlv0Fq8f/5r9UcpRxRJ6hVjT6
QjcmKGvZg/E+mF7c3uyx3gocURQ73OKsOBp9Xhe6SThI6MhOs7KKW0Df+ggvn/l+
eB183YEtu/381eGpN/WbsHdynoKdeBfYn3dNPJWxkbb/+hbpz2zNE2xqvuMiFZ7r
mxmRdKLovENnIIZ9my/T0adk5REBL6wUxf0M5TJsLpucV5msjAno0e30VxgA53Z2
fqKf8rvmjIKvKi4K5VDjDnFDro0hGSlhdE3qZDkY8qjQKWfms8hzYE3NtNPXhJeI
l2dIyxetvAyn8ghndiEXvWzaqTuQ11vLz2lcMYX+vH+UJnTfIK/43MtZfMMkHSnS
7LNIC6quVSXU0zp+3Snf5dRVHVID2kIv/BPrmxq27VK53q7KuatOKNJvTmuWICps
6BNie/VquK9j2WrGgncJAA+yjV39KyPznqjrUrsttdTpCrZbC9dxMcpOOp+ZlBp3
5FiVpCCiCFVzc1y26/PpH55jz/fVUdqXossfM+NF8fE0A9hvQ3vCUu55LUiSlxkw
CjO3OlctD2PG6bBJJOvnMIoCSHDoLm8Y8BrlWCIVw4nTUlfTQQptlUQzN3DHznEM
L0BPl+wY1RZF2xD0NvO0mbQKrrqJbmfqHpEJjeg6OQWLkUQOPdRrH0HKJ9LqkHWR
zIBTsEa1meQfHZuXOyVaIkh8ehZZVKmbfFANz/hbCGG1NXG+kxvP13PgBY4u/Wsd
ggBBD1GnBBG4ACkLdm07aTSboFIuwRjl08ovyzd2NCPcgJV026rx09QI1U9beNiz
sUA3bQGWetUwJhhB/pJSyyXRi1NcEqT+7CeyHYCvIxbjrjjuwLna5Qh2qNBfVptP
3qdrsXSnnn5Th5pVDy5W0qovGvdB6ozCYGtYpPZuJMCXJR0eGKyWqbNR3LxC4oCR
5J1DL0xa7pLWG6yOd3AzJnFGOENCsRK/WvuCS1YeeNCxqrni3YCIci70wCsgYsnd
KHxZwud869aH8j/E8GpRcYe54lAhluJ6KnZl/GVuhCNKCXRYW/zmib1J4l6IMtHi
fCtdQflLP9jZOUASSaUJl2SYLBBpB5mFkU/6TCz3ICCpevFXSAP9KsMltubZeYtk
w19ko3t5u1guluu30PbKuPdeyN+egU+22+bun0Ao2Q/zpkXeFCanTUfw7P/1LPpi
dm1QANiUCkAGNgZ4Fz62Sh5GgmTkr4K0ai0BXFhJkGkwhyv/8uwtbyjcZ2SUMViK
xdCCykL5t4DF0WzIJ/jcDPQc3U+xjRklp9yMD9l8f2E1GZrxSDS4hv4gfKuKNCww
Hpd/wM6C7qqJ8JjfV5qd7qSuyyS86izBgvCseoVdJen/PxQ9KYu1GpMeaHZlVgQx
MNvIlQ6b3hrIUnH982S9bTiie9eeWTV50URnxATnyDbdXOC6yjrBEFHOWICXLg8B
qraliA2QnxFayri/8R8Etgy3F/P9YYCz9txSkrjwHBSjqnAeicTTKSSyDN8mNa2d
1jdR4Q3VkHhV5QuJOXIaT4KNpPsXEGyI/F2QLOIMn1I1u/9E9tjomH5lPGvwGzQH
SnB/MVHjOFgE89/cv4if7KkXPTCqN/yAJW8/8m3Egmu2cIpojQmOoGGi+EMirSrg
fBvRs6BK8YL/yb/LwPS7FWpZBujkyhVN0KQJYG4Q9yN1a8s7RsQdr4VOI2c9UvkO
JVHRpGScMkarDzGZFBWW8V9m3CyvGlGfEyeK5HE4aEOL8+hPUIrCcyu/zBymWFkr
bS9GuSL+BEJCpGdtX8sIwmjrUVz4efngforq+M/UrPTlb8mBi7yUeoxMAEujgkgF
63kVRH6CMR5Sd7g3ydB5fAFnQzjxXo/00HXYawJqZ5R6z1riXnv9hpJK4ko7jHLw
0Vu4Mv5fK+Gj7Rh/c9nF2JK1lPwpril8GvdzvNUusqocsYT2ulJM0hVN5HMyZd+e
v/dWIDn3lv7pzLCFS70Y7bqrAHuaNmK63gTQT+/9yt/T5vCetu6WDmLOvPQBaVro
gDXmQl84fdLPA0yCvNKkI8PvWnggh9I1UGvBKBWNX170s7xfIoUPKHYwRS6KPOLu
GawDvzb2MwhyzKLsIIC6BO7nCD/AYyD2B/X763KcMQ6j5zocHXuyHu5DEcTd3Ove
P41PJhYJK/jKSllWPo1rHBSD2wl1H/klTM5bbLZjTuZ2qJ89Y9J14U3uoU4x1v+w
01uHHma9zVoguHQOuY3Wp0duiZvSLPp8zGaMxdDjE876OYw6xoKpy7p3EbO3gOav
I3fug53gnEqtroUxQEmHp3XU4DBKiTJh+DaLgJy4THkK2xM56PKp8v6+BP9rpKlE
0/sOebmCEkvlxl8ynYnRSpzSrgz53F+RA5alQOufKNiayA2CYMtCHkPwkTwYx6lu
CzkTGMIXD7SFjbcaaaaF21M9WmRtsyy90uJ1uKgELqTkXyI2DIBjSf2Mf37BHAfc
5kbOhdLgDk5zcAM/qnZGa/QniCLm2QO9tZhHneB43P0Fadgg7532pEzcsURQTH1a
XW/9C/ZX68GSN2KOMdHZ9Flmjs0IwUHvWCQ+kvLXJo/twmtVXV9AX1cYcTkPGgwr
4CJWP9oKArIC+44OhzLtV93K7bjPlQavE174NVTRn1J5wWMxr6bAstr1bFPPdNFp
3uwVZQ7L+FkmEKNUUGoYl3u9dGNyMCRti+epyeLXipeGk+xHR38WsIqmd9HuGOS6
fcLmqE7/MBz+gucINtbEm+xU2lkNNhhi0x0tz4oLwLl/tuVj7lrTscKr317w7D4P
eA+n8trj2bR2wpRImmoCb/i+F28CIoh7eNXcN/umNPuVfq+7GlVv8MOJKnr0fDkO
waQhODw34oW0gPpN91H8NoJS1mWgE533GI7QABpLBJa/SY3uIBM+PvwABpvgUmxg
Il6op/vPw0E6KZPfkksGHDLvznSUF5q50zac3NvF6pl1XeFRi5NiPNa0RsUkHxEk
6hlEloQKkqBuY7P/BxhI2ItGVpDnU+zCaog1U1hDkoXnC4BUnlM7AWGNzgUuBz22
nNn7PFyLWrEPI7aLXBtYVRMfJQY4ZgL61yvHTVhZ6P7NGR5GkcmUrp7LcHPriVbW
zBeXbkhx/MLlZaGUG3vYIFPGqPBjGUAZlt9G4ZfrzTQ0J7wii5E3sDD3hC8/dx2s
4elVapeNpjArD2CLCOBKGdJos7CBATGRFiPRoIsx+NfuI8cBfcaJVWkuayDynLkl
NTJeoRZeYs5DGfK8ie/i6JPuW7Y0IxW3xjFocVzsWpNNRCyfLKJ/P13gz9vRB/cD
yj6XH4SBYvGqEb4u0yfr+HgDT5kE00J0HurH3Nr1RAUrq5JAI3G5cq6qSgJqahbz
c599Tw1BJ1JjHcZRASpp0lBQyGxNf4O+0RXD9PUITViFS9A8CtPdnDKN/XECYgxp
Ryuw0wQLvEt1r+4BgegTrjJ4wZ6f4Wiz7hvCCrBC2MmhmRUnvym2RUUM3Ki/r4gl
AfPTieB+LPdafOxRD2WhReVVal/MQ8x2wbezTA9uBxbi2vYbOAr0CUljz0M71nqI
JAcf9r0lP0weKZ4wy7I1tydzwZHgxcwwKG3bsLeyJZp66bqG59qcqq0J7G1KyvhL
ijBqu93Jj7OG446tkaHHNKvKCB+e4PZRIeRGSHvF/pM90vubHnjwddF/Vlwxhc7k
y7lzev/ml1sFVZS1MAAgCpKBpN8N0+Z0CGY2ziDMAvm2LtAeHzV7cmnlaDG3PS0f
mc2TYQGjiMGaelst4DJVJkEoFyUBLJc1C6FllSQedDgKnTksNuv/1iy1fL4+vpYg
khCzyZ5bRohtlhHXOUd0UfpSBmtOUXppI8kDQ70IR9ALQjxwgAuJKKaIWde3otbw
uc1LZChoeHrfRf6MYpOFfCuDOOth9I4Hj+5M6QaqJdIeGcoY/Zi11N1OG9XKTgIH
GIo2sxfKJWVJIld5fNMV57zNqSJwLnctktkzFF4BQlO+jEyy6t0nNbvyLo40MWOa
QiQEfQD8g6u85Q5QUIU4IpUKoSFpZ8UoZdpBHv9fC7bTwmFC3+pXvwQtuzatoAgD
D3vvW4P4YwH3qTTv1BEBmoL4QuIj2dk6PADD6AdRlRXAfPU9vE8fP8VjBJhVxURT
p3e4EYWnG5KNj3QPVY28W5JUb4GJ/9xpwHThSCtcKdSP5LfdvmbZ0WVOJWtnrsOJ
OqmDzUDau4GDy+ZKQz5JCC7ESuxvSx6OrJ5cTxhzznmcLJLOm4ZDcf8VzKkKRiaD
0FzuLRAVsLKGnw3dnM8YnjJvq8l16exnqtCawZ7pOdVNLGzW9RK06Hi3h0mdF3EE
BbH3iA3CLUVhZgjul2YmLIeWegTD/WIX442TwK/j1L49FhNKQbZHG9F6VRyOLRt5
wcqjMEoB1AU2nUYDC8h4QP9rqmfNng03EaLbuWrYphyUx1AostJP5oZBD0ki84x8
KbeuEQixTq3ziuc/1yGGgbWasjHIGQ2VaY4Dk5YMrH02fcoLTnvmGoRrhGdqJZP+
t160eG9sHdgKQTL3jpqcVLkcA+/IxM3SfoP6WPq7EaLFhcXoDNFEhUqllFFYtSqk
N42txZBMmWeyH4Lj/sbO00L0bN28ag2579R1v7GIhC/rOln6u1d3ZsQXYNSH9StR
9Hn6Ipd3aC67w/ovgl2XhvLX24Giuja1PzeNl1tw00X0W71DmJ+57dRQrTmCe2vp
KEFFx+hOdN7zm3O559U0+S1Dir6h8HSeQv7vzvselh9oJP7fuzCGrIzijdKQdNic
vxsMNR3KxLIqUbFldj+HtTUyaiumYijXfv34JBc8i9wxMWbm0iomioYOJTLTcJUD
KgApdnCv6gCKi5AA6tVQE4P9GVD8AnfQu29Mf+Hnm62NGS/AIH+Wg+zICxkQVXFv
SvOs+iCOvVk2ykW5bWMx9/cOlxQetFqjsrfkHZ0SSiWswzQTujZqMs4GCMwWTKs8
AK2aPh0yzT132HqKeSZBTbIFaQFBYWItLaAh2PkAxspZosEHhJMt9GuIzEr/Qlrm
t4yv3aEJGIBwtSdHtQUBi+WXXMdQiWMcp4iYuSAW+tFDnhmY5S44bNSBXbnOBiws
HmuQ9tvC8VvfFlMRLHl8XPxPSQWmeDsj7qXDIV2q6FCWzW2tcH0Tizfb73CGn6v9
l+3xgVbXlBVk6OeAwmrIg4ZiQ7J24h4w3y323iow0ItVyvxb1bXHuiBGpXy58z24
y+2g+Rba7fuxyY66HqglsuD9K1SzmUEFLMYXhrpMs43AU9dX70AuxPsicjdk+RvD
0KD16eautbpaRx4sTNJY45uuPtHc9Zjn3svRD9sV0m9+jgtagIOr0sB8hWIFWM2N
aSrbL/KTm2/oSDufxMq9lILuHHybdKru/MtXZh37fPqP0jt3jSq7g+8p+H1EEoM6
nLmwCUrf0/apO8MMPWlOGmZmGBtnVX0/VediZ/HCtiz3ygh40mlEb0KNcAdJ7TtN
P2vslelgbl4akEKc3337r5dvUBHYc8H7SUBcuTeNyEcCS0jZhJMUyGCi1L+x2cES
ZIHLOcq6RXfPluoAtkV8gQKKJJh9bik+39tpgpSnoEj8oHDFHbEj5I8sYrM8wzUy
ZYU8WP+PdthLc3i4v5P0S+SuTrvbiFjyT1jbWH67CUW0R/ml3hkG1CGXDcPEdFsG
ccytnVaaFYK9qG4CbsCjHsch2Q3HV1cX5Gpmk1oCfO10qZJpanvR4PznFhU0RnpI
AShHXkIoXMvBO3vHj13AKCrjwRitkAiNytapudegGFwnzW4KCZKQeKuRTQNVq36P
83KKz66bMMhHzTZFTDv3jO6EbmvNwJNgPAPFxq2CYKlUzicvVIfwIxiNNnGubgwm
NW4OTGv3NTvh89yQsiC7n3AFUkqRpsoS/v8xfHqrB5Rp8yJLX4SVG8mLO4B/AU3C
wJpWvLsayJRjPM85Fkn5HIznNmgmufimOmWQd/RfDyQdwHYmMCyx+eHVOL3CXXIf
Dxt7AkXbNKD6EuA6e1Jjp/mAv6M38CKunit2NuTJPZTGEC/1ERooY7DrUVT+xi5H
2ocfSI/Mokk8Q76fQUXQd6WOh+NEcQOuczINKuvraMvNzCJbdVE9haJWCJJMcg28
shlqrQgzynVH1dyQb5SKyvjM/pZLQoYuxFNHfjoh/s50coUJWgeRrX7d911gwltt
1g0q0yEJJi+QSduqNzsnzUenZA0kyC6XIYgPE/ahlN3nWzRnJcNZcKNM7dz1ujpH
5KbMZp+If7dWw/xg62aW6yIbdr+EkH84jcNcGi3jhg1JFBiu2DXMEYP0uEdp+NMu
kt5oWMrF7R2O0sYAO4M0B/C8yMmxDsIQwHUGftbdHfWuwAsK7dnvpYNoy+V4dVp1
saLQbkjaGZMWdC6GtDA4wfodlotwLbFOCRsogn0Kd3Q22+VFaL+cC2/kbpe42j3+
EQzHEct4WtPO/drob/eFbO3+6P2aH8rZcO5jyRXmp2rUjxp0wMUvOhaPQp2vQga3
4M7a7U0VJ3+2HBylV0mMPNUnHD7EoVz7Y4kZq/aJ2D1obUF5zoxbIDfg0oH+rUh3
PTBfP7xmhh+dKPHO+wVuRrPQeFI37/GUybKg5ViVD7IO+qMqkdTYvNFQ6vDm4IXd
roQzHq4HrMbb318lfdRSuQX+8jPfNZTPeUXcNGanUckPXBBzhjayl1mEMwauHsXS
3VB+8HIxC+NgSBN/3ZQyZRAJI3X9rXjwwBgcYkdyu7mPtnCqMjHyH+mPq9D6WmoK
dR8CvNiYswXfM6ht8U6TI0PRz0vZSd/Rhn25u/hkjZczH2msG3FlAT7RQjsjjtED
mTL6IUxM8Mps2n+pVE5AfFJ73CprsJ/BPSFfIuNiy59YzXjAPY8hfVZnt5h1IbYp
mltBgOL5zN4Tt66lxzn71QVnZnlH8Q5cCx7qZozZYJc/rLBsGDAykzjHJtSll+8X
wmWaH8SWXbm28AujIzcu0JN/UhBhxQ6DGBlbA80DwPVDvCsTY3EB02tFOrkfmsky
FUvefyXHQkbAWPfR6rw/M5kl5Gd5isrTB3LEqqIlJYQqqqQHIfVy0MGbzTe48EUt
4BvomIzzbe2BOcA8b0uzpXBe0jK7yp4ghV1P66E0Z3JQ4RFvwb49IXzsDOssXEst
9k1r679U0abvWf9PHmfQKJspHhjUUyCpKYVQ9xFk/mC5621nUh60a92O0Ynz8ny9
MQ+xlT/C8oXUA2rY/0i+9WICPVXzwaNw81cpTsUUcHfLUhQVquk3Imcm8tFqxjhR
ze4ezZA3MaTj1b19+ANLB4iZNdi++wHme6TEK2Yd164dhxeI5+IARfVtttjah/DA
fhqzhKBK04DN5GU9Z3b5wM9ZYuKcVCd+8WTnPn0vAD1rD7WRWW7uW8bzHiL10OMH
C1M7q7Kx5dcUmrILQfFZkFgZPOSqXX9az+DWwcqJQoBNlXzVNkRMt89zX2gRbWNk
qvg6FUZ3pq5h+x76pImhZDwX6BQuYJ8AwLfc2Sddqao2QyDFRBkGAIcdJQkiiN2J
AIn6YlHMrbqH8goesKBnkNqTEzk/9kltU4/DofTPAo+iC4st/i/fx1c1bzDwgnR+
8PU6UEhN7Bh23TKmtqm0IO2mmlhwQyrjCD0d4qywQ3x+8C8wnMqpc9vdNqQozajC
YoO4L0ay14ZiikgVu604Xsi0hSpskrtseqVF/d5Fxqs3PF0RiVzpsR49ixUhRIJk
0nh8EQZTRcPpQxthrnctvxcn7f67QPU0S2wMeX2op7IZgf0M/n30t0IHVWiIGF2/
f842tH98OJ4/8P43z9dU9sDK9agWeUYEfJm9FVy6cKKJ9Bhap2Pt2FSGuu/g082y
75FWUqD3Wv08R4BSZikApYozZ8/NIFSr2vjjLW+9Y+7rPWFh6OH2ajd4z63TlpFK
JHMgtOBa9fBQk55zV8ZA9X10vfNr02gNaf3MfRIEkxqVL1Z1qWVxKj0sKa2uOaL4
JdOnxq7iAPi9BNDXIzNtkSRGAJJCWbZnsclrIFGTK8ZEUug/AskP/7hvc4neMCwW
4oqPA6ulRiBkObtwyvsI5zaKqonFekZRBFdzGqSeoDfosSw3TlZVod5lN/6pBd0Q
t1DH++eZDkSPO2FU1500ZYMiXMmjQ//x7ttD9sCczvF21ZLVOJtnMR619cCTX/iF
8WeGiQ5c//h4wsaxVFbj6WM6acKcb4M1cDF94xtvu5ylSzdApjIqy977YdEq9UZ4
n8k8DJDzVMdhUwMJITrFlAGnClKW3u3Cw+NGFWefMMdmJ0zKmZ8XT3j3uFnCX6ls
UY+uHzm4KnHUw3NcWgY4KGI/wix+wTIMLAfobTFPbbyoazUcG5RQS8yGQvt06HhD
bTJvc0gEfeeycqkbSvkNaRExyNcGkUzsUP/X4CByv1NrdbBOYzs4i0fo7xLKp9N7
JKBCsgACARH93QzWNB7veeBK0YYSerNPyQ4+5GTGEUCrlO5HD30p2BRtsbaG2Q5m
4CIKvgJPP12zLko/NVQPXysbqO70lcUZWnoxQxq30Xm+1P3HLzzEQcN4ezswTfCh
sdExb7BkYM5Js2RkL9q3a2eKrfuCWHlBPZ6JRtBnTG8mHMwe96ajUb3kuavXFRW1
hALPFjm26fMcF41cBIct3007oup3kTyZJ0mwN5lYkL1gBow8up+XK6T81EBgI4PM
5SXswZ3yaEDI6789nF9fafb4h9T5ChbYl6Ce2AF2kOU48uVmIU7ze5MhBmAmFN5h
UCbYxEOr0JHYQQtKIEYlz1bVaLu7VpI7J9e78RN42Hovlx1jYt/ZmrMe+r+jN9xC
TJ26qq7asMMC2E57u2ac9NNAO++HGJo4ppfnSiJBTgZOsi4coEJO7GUn4pWxNujp
BTNJXAquOrr79zFx6kSQGhgICAG9WEL9TTpACdw5xhbllPYUEqGOloMt9IYA48M/
H5ceWlyTBQDj6CyB8mDUM1PLPNMlASQK4rnTB5+Mts4ifGCV04t0Sg8+PmZ0IPWf
HThHJ7XsNP5v0GPiyIi6BpKlr9D6wmHucpw2BjkdP9iL6IGKbsknyqO/JoED8LBf
BKd/FRI1mXkBj4NkzWZCc/lG+g7lJCUSQNkPG8kwebVkVSuxKbLaaxCJ652gcuOa
qajoWlPjs+2tCCNTSiKI+FBYByEfapjDVAXF2cxOnPDMEVZ9c0IayeSkaIlivJgg
jfiE7dKVFOBbHjWcmNl551PgD87S6eu5MaHxupr4UcuVTGqNIVm4odWhgEq6r3Hh
+1EuBAK2SjBSAZw51cOwkYfEr2nCnxa2vEHbTcpzcCYUpA+QfNGsokMAw/W7CGI+
JZJ1IQKRkXkcMTCqCM6LXtJ5/wTEVcFPQVTXiZCDWKrLIkklDNx5hz7IlmZDgC8b
OxkoZ+tywmBAz4vLhV4TzZQt3h8inlITV4jIt57bR6lAP82pV1mRwWSYjUVzXCac
wjFslKXcqkClLOY5kBKmD8ZpHa6FcUtf8FIOY8bWHj4l3oA4DDL2mKNKJF821FHi
O1od1YJLjNUMmgZkgfrp9z/mULl8jGts4HCT8sFEFUZhVmqZo1Som4sCLVc3wOXq
B3dFeaXmcsSTgcoVXZRDiqhuJ1ses/DL5ZyhEbixvTR6qXuM5J3ANXwvAUE726Wa
ziBJwiB6mtAFeBJ2teZGNnNpw/0lrmlc027vE5LiFEz5K7G23xe17OlZUrz69FIl
I5Gjw8Qk50Y+0/sLgi8RRZ+NEsSkZlzCH61YflraXJ50KJKneRI46/NBfrjS56QY
dVV4/G94OIyCDbkXU0kppNZ0sv/1W31c6iMnr4N+ysTCUNe6IO6eH0zy7s+PJzVY
/+/iHH//n31uuffiwLNixbkmIjs8QdWkIL7DHx1GG4ZpsRRWc0KvOEHoJswsYQqL
o/gWqkey7rymJUFzC9qHdAnR9EKblwqkUx2kWwaLGaXAMxD8/OnTKazKCD8yIPvw
zUenHI4kXBvwEAA5e/WOHxakFLBmvq7QswNtXMfYsiv7bLh8y5gF5cGldF6TIHZ8
i9OKd5PJZX3ioYcnBP+R7Crbq/zCKP069HVbzq8mj+H3g3yagzffe8TFPVTdKtCM
JUVh3rJiPTrRA/ShkIhzwDThbsLOny32k3n/wE+eQpW3R4/O/OL9/do970nftcDB
PYTf1Jw42pRYqlN2J1Wg+Uj2f4ffUC0nMrtyHNrkhyr9BY/UjsOdMV9cClB8I1Lu
kRSj6Vzy1x6mvJbFu8tsTvvmIzZgYwXzIdY10223QInJzzIwsE/oIB1E7NsCvNrt
wmKcoNydgIr8ZIisUYopH5mqj//aaqnpHR1+9VwGB8mc3JZ4uL9ZKeHWixQqZWDD
d4ivCSdcv7IrO8rlo0Z53PqR95+9ega7fkliV4cuxDvGRniwZJ5Mn9eFJ/vs98eS
sVHUsfHSkOMwGcnsk98XHd/qeO/10BJIJpXRoAMvJ/aFasgf4M6j1tMgo5CO9rpR
QlF5tExjIfgzR8wIiRXoHma9j0ZLKgFSqF5h532Hc5lBUmhgwLb9UKi14dyEHH9h
fkdqqUD2k0NoumrBDlVALRV05aiFHgopalJ/pz8tsbwECXFkZj59ieL4yVGPJGmX
ODSxdDOYXMXEcdmhynH+AO3Pm2aMjnKtBon99ym9twLjFCc9iciIEtx7DyJrd07L
U0ipWC9TJzqy1VrcH6tykarrG+uOV6V+FVj/85aWjV2GSSa/rqMp7/TEFjBrhijo
rHBcgh+NuV57nI5uncZAZjOQuQhoUg5JIP8GphaW9GpngYtuSnlb6+gKi4psXQ8l
BlUQmH9PJfJpPvJWJwysaCOgaFxcaoeTxhqrsB3D+WrIdYCbS8iDvqP289ZxGEfC
l0HaKZ8PYVO1FKcdpQvDtCMxeqDUurjihPygpoOFegAWnuLhFD2sdjgOc5hTkPRc
VSv8HoNwtuJN2Om70QZJrb3LZjtF8oO3rs/kAmS85kn/mbPgeNKvdOpnschbQl1n
5o5XFbHKJhB/BgQbu+mgp7UT1eKphgJC8lf7FeAoiEJCBLmDTozwY244tXnXtBuK
ruu5LyQuZ/qRqLOXws9CUF56Qg+n1IxyxYjK8zcogNnYPy4sLSJ45m6uOk4nj3g1
Kdm0rzqdwqRFt9mzc7zwKEMPdobEXRO1ekTR1f1dcfEGjQCQPRbzPyy8/sUioKxz
AGmDszQcnrMhhN+v3yLM2+iFHmk/ZKj5N0fy1w1oIAnWuWVtZKD0wZwKchthc2Qm
2lNXav2GyGR6A4qWkEoIv56lXdv7PY+mhfoE0H+XpoIt5QejX/lZeY1wNly3AAlF
5f8BAGf9bRAUh4xogLeimH67gbhFzTkFJNVPgAcLB/ile+5usIWcfJmwWtOe9bUc
oAuS76eSSp/sw4Df/lk8oE5UBYpGtP0RMvuouAAelmPPFXgbjEGcac3DLQJLVUnf
wAZUFkssbEUiMhjCZVVzC+lPlnsI1BetXAhWKg59NfuUG3p1YYTxeCOfvnRv6iF3
+jB/70LzL24doOLD3eoqyJndFZiMWGajssZ8QqnlmC+rKBZNe6JpC0YvSvSA1L/X
09lX7s3aP5r10ShVMgJPRqYRAL0As+iT7iexPLrQD2ursETsXBxGyyDadqKzAJqd
ij8Z4FBNRKnjQkgK/GehKjdSoK8dPLuzHa7d9JVrq3JocNfHQ/aoPieRDfgZMwdp
e2s+Q/apj8ikkiGq0Ogaxq2/Amp9r2qVHsEA7tEcttAfPRpZCqL5nutxVh7LN43P
cAEVuXIpc15Sx3jMPIxjsjFQUOLftt7WxSZc4exUcwIoavh8tuoL590aIRoqiyKp
wxTEJMgYDEvHV9b6an0/eb3yDZ8Bqfctm/cMNZPFdxEg25iLet1hqBHGi94SB1TC
bZdmzIbJiCvnvOHwXZN8TmhGRuy0h8DPNcMUXMZyly4gF2k3dEYd8F1BJeYp/M77
gTWz8e0/eABXpybsW8HZbxvoCc8KzBaGV+gZH9Zgru6kBpxR2mju/AEayjY9YlUl
d88q0zhApScaBxQTl46rH1CGQXGteCEVrwLe8lxuREdtM4z755ziK5RqY716CDZF
dnoZdYrqsBPAv+OBjaRbM5Dumpx6nDcXlvfOwnHEixxQ48F7PECLnhjPYHEOGvpW
MoFAuoaurmmr5tfUBnBta2KPeDnpJLi7x3WYE7ZwuZ+ouDDEdYG9Zf2QOvmiwEpk
O6/mVg3vgV2mDrCiTCc4k8hJItQSuMQR2nuLXsCBq1ppQ6kFjjC2ipWoyVTDyGyy
IEQImOpUzy8Y+gU77HAD1rdsZU3NE0jajIkNywoSjuRE1q0Da43iFXLhvMaTQgAv
sEtqsspsqsygAVsxhhX/YJcLeL/vDpR3kuLirnIEsv8FhF5gfFmFyMm92x+nlQW1
KeeNqhJ4P590lKu81uv8MvxhMaEI7KTrb5yU6kgbGzZ7W7pjj6w3lBJ89qo9dbBx
p0yMNvuAUX6FwjQCVLFXeyNWolNRk03RbLu0HTC7RaA6uJvGECj5iFSM82cBOMWP
FFucf1numHFEhX4AVRokEhO0eKgW0LQy+rpv9gDDaobt2K2zG/UM3/ms+1uc8D9C
oz+XWOJzhCO7Pnb7E/Oyib4AcbhUbIMWB+20PM2o1POQBqavd8ILQCN/SQIBAvWr
ibF1ATcUYSriKmizx5w1xZQqX0AHnhhNcD6c0xtn77EzhoqKqLZAxgIrb5Nl7Ft1
ErMdjeVdRLgEFO9XE5bp+JP6t7HA5XN5xeI/p+Ees0HAKa4OSA0/5s/iZ3Ebl7d9
lCpZu7rpZU+XdBBmnK0r4ZDAukNnrL84Jq9gknh33y8yAO2o4CkX+fpha3mmPNU2
VOFG8oD6gQVvYUOaGjQrLMLq07KRSM70w+xpGVgYZ2nVqyZGBLjIRlI0t2cxP2HW
jiZmaFWjNVn4RBaSi93vjUCCoA43fguSBroPPbih/Knck34L8+wYPMpIBZRHuZkB
8kcG6ebzGuJc6k/iOMQvB0zm9Z5aRCdKKX/OQgdLxiyyDT4oHVzA/vf/ouzC69R2
9fFmWCqCQHCMAyQxxyyTi91tucyBqRUCO4ACT1fY6CTiGtDyB2MNoczoBpVl7N1E
CWeyF88co02CI7gfkOYbO3EEnrpRBAtpPGibIighIlraSDmOixyzkR1cwbtoeGuN
vGi6Is5R3WYiQV90vCp1HQf81htB4eS1eH6uBaNM/aDjKCH4xbBLAu+J0MivbGbc
OI03K4WcGijoZbSJjq829G4ZFOgxomSzGYyjPtBlV0L2SVpwqxFafaYVxc3OyeVP
eUdDpEdrUHcXUQcZBQCagQXMGarWWEBMnBdEiYkUdobid+JNXuNf6S/9W3ooMAQx
Zpril+S07i2pcISuyWRwz1PcrNFx5cUMoAjeReuLbGDwxn7flmPyXRdNAOgUU9Gv
PGIp/hTixM07rUCDSoU0KdudFrQq9CqHn2mlckuAUMCNeufDXZefq2BHuEifNT5B
PVHFiEBvUaEV19dWk3kpCwBpDbDGYvOfpq8h/tJgmSTYZodnBW7sH9wAzNH2izGa
UlkymomuymuO47C1BrgDXW9/bwOuwb5vMUK9sUj9K53tgPbK8+HuFJOHPaJla6jW
YAzstKojnupKN9XABCSu3dqpIDKBOI+dYpVTxGUObZ2tvW00122Xk9rj5LfKHt9c
AP3Xjvp13niXFM6NULnDyrL9u0V+hOgQ65nsuEDBSaKb46bLFhEbKaFNcGpITonO
SOQgJFqnmeybdr1bD+SU2VLzU4arjVxNt9PCP476o6/+nLS+6Dvyam2oyG20tEau
dDLsezxR+EjdayrJskJffB/7KcqKt5aiPTAUl0C6Un9gyosMibMU4rvy3N4GzqyA
s5aOCPZcSY/1HIWk+saQin8RwBZ+2VqODOPvNb0pqdQMSub/a7XaXjNMLbb4/wtQ
a1ie/ZgQfcvWsNq+5/3TMF0f/XgdtgvkDLRHD+HRKLZOk4HS1HF1y9QcwWcWSsI9
Gvdfk+m0bxADA0Spl/T7sjuq/0itRt+Z086vNLtDphQY4C7D39PmOrWR1bdHdI7j
Vv3fwBdODqKjCpVqJpEFuRuLhd1vBUzapDz8K1JGHmQQVm+IJ/OPx8GuCumPd+u6
nmGTPofZGEbsbFSD+I1IF6Mecvl8byWlR/TrV903ABfEk5WAj7ZwJDkVnURo9MVY
Zm60MsvVyMaIWxq00PBPjdPyMG1mULL7pvhGOod6z+gpBOP1SRKrRjBfpSsr93B4
52yM1fA2Z5+zpt65kco1AK11+uV47zWfvW+pQzB5gOHt9vAz8lhJhIBJJwEvuIeo
o25zzxMlwP8YJ4Zk7keL9bC8Mh0iJKCTZy6tPYIKsy4coxfwganDuLBrtwEJzWE3
p1LF9b284XukQRipo4uY8bdyW+tMyE4tWuKvAggXD5K8LLSpD2QQiDSYwtSlU5+u
l1qG4fqIboUmao41yI8v3yrXyFrA8SzKV47ubsGC/xDdnvFPCxEjc1WwiCfb5WnP
j+OYWeBnBhPkZ6nrHRN15Qm5OLcqUfDTU65YJWTPuPdo+/H4s59cBy6Hm89fmVXN
BzmMDJNeCKT3vDpD32Ua8acvXbt8LUE6jq3V7ASUpXpUotlo3Ler7X5jO56zcGnA
+6QZFWK7fDWqprMS27FrpKCPT2Z55dFYnEX+DfBIoW3z6v9dsxHDlaqEI9ngSYTd
w2pKfNJOd7HobjAV3VuIdv/VasgexM+IW35e7AZr4GKhzfLWdwgjET1+B2JY0u5E
iq4YrNp6WEdTrVjl3wOPP1ltzrApoFcQznWy+EYeQVMjK18X1t2AxxaaochDWoBn
t9R3ubSXMqGYjOKJuO+A6OnDam723V4WcXIGHUCjRHUZG0bcA28GLSZbQbYDMJEn
uM0ZY3pJePPqBjafnKCg+EGxJE8XipI4mGmwHWHYe/Ci7EzaANmoii0v/Y9duTgt
H7vamwzkzRcxn7maGn6NirMAgM6BY3UXIeOaj/v1CQTLM1HCWIw3HKWsVS48v10v
VsodE50y2pg41pOByyeqDQFdjneD3U4Ix51v7dnD2TcDsFBs1sifaxp8dVSH/2Po
b+KMuUKosthP2zbNUsPJm+WsnJaBOBB6FEsJDBmegHIi7A/a+/c2mRchrxSQcwvC
xWw3E08Pe66YXBULQRzNIR7WrtDpfMkPjVe/9cAORHwDxhYXP9RYp83UrUGqVBNJ
A4q5uXGlWl2mscz9WGnCaNdIVUcoB3aodra9ROCtv+vF6oanR1fBxc6ZiwKhEDCt
22UGnc86+QWR0NKgsTfyl3PTK9i7XlvrCrOvkxUVQKeMzTWsthGacOKR+qfBttFI
Dv5Bv3t32BzAknUGgFnRlNhuGVsgbb1X+nIRBnT4vxwjZWwCIHZhKR/vZltODqdY
Z/R1jKgeM1BRjVmwa8lHPjnouAgEAYgskTAnntiL1kZGP3TrMqIfrG0ZSCtrclrP
YPCFdP79Hc4RysPYWM9MOb5OVwlrbDGVrdLNwEtT587i4NyqxvIqthkggZp8GMTf
3TCmo9+hr0yH4su7+xcMV/fZ2tXipQ0Y90fpHmgK5HBz3b2iWGlcxl6ANAEF2FQ6
pdCxnUgoziQtm/qX7u9z9OWyxNR+DHvylUlTnbXXnZkQUtp4yyQHfAtTGvM+Tiqd
l4QD2P8SMuUe+UOoBOv/mqOLw8SfNT1cHOCH0F6DvD5EQ07yrkhUp64Akc2yX4QK
I2Sygnsv9AjvvHSwjx5XGwEdOYG8tTquRF43VLUjqVlmNYuZryp+xhNNyXIwM6yp
/QKHLR3s0mLK4J0VjwqI7Sta5tkHhdKzKqIuEloWZSm9kyE7lv7zMF3kEbnTxW7B
hIrphtbg5xSp6FIdq4AEHhQdwnI1C74uj/ORDor2M1B9dL+IFVxxTrn+FwJos7vQ
zJxXz1H+3JvGR+BGKIxzuKtMAepfCoiSplv/QY4DdU4PoiU6atpjpN3N03M5Ap3P
gzbkzFChCdiiu+yxfSuYcqlKiJ4+oCADs2Cuv20vfU2NDHr8eHGMlRapIdc7N0tu
uHxkOt2W63iM4cnDycHXUYlTMLUALQz37rp+gM8PaxADn2Yj676oNHc12Z9L6lB/
5BCJD3EMPXBHKeA5TvjP4Ak4KlLun/A9YeynfdP7PPAf3hjOp+7Z8bK4U37pDIds
d3tTYki7fSi33GSdBZ9hXQqy6oSV2n4NvKWpHH1zGHdxYv2V5qOq0PoUkqtecx8r
/Pb98W+tFyTp88ILi0hhvfPTVSe0QyvqF3P6CSCSSru21bMeQaDDEgBDvrqHlUpS
C3dIe2w+omO2ceG6ldifYshikeujtHwl54bM3DD9sGpRsBypzOLN3oO8uK61TVDt
raFh0SPx3iVwZUHr2YPSIh/4v7R4S3t5vWYdthOYyK5MWKvNjBmGiNwm0whHMlbP
qBZX3sINK+npGuQig60oRbYMK12udLw1dJJL3Ak8f1EButBj4NcBA+R6DDULARdD
TOfsYkoq+zw2ou192T7pTvgRgmJSEqcUdfXqb6Qa1ecUJwQ5mu+mH9Z4lokM2sjY
fLT2eyJ7evoDLzhrQYOeJ6uF4A68W5PMbOHs36/PjHaIXhgf8z83meWbUJPdVBe4
dCjI1virrNnkAxfzZNo+xgdpH4fJgHV5WfP9fP+LW1HaHnr0OCl86HmgSLyv9vQU
UOCtuttWsppgkw6UQKhN+t4p9hHyP6Umvw5Ull44DiPYLfBKUVkv0cWGQa12Z8S0
+5MrwFakCDU1U1mQ+9i1EncJwZi6RPC0HmO1HNf50mt2HDgeJq8vcwVCoBM7Md6+
ZBUEnBp+tTd0hJ3NSNFdxgJDEpR4/CMHCQUliNI9DDmMDErDpejd18KLyEalhQOv
y4ZTOOdDdujA9gkTQL6nwLw6h7yxucCn2j2RRGS/YVe90VebiAtaKPFqYW1b1Qyw
l5lHNHrrFHoUjVBp55Fs5ISXmhqZvsszjhHQVmGuD/OKf4InTuWFmy6+PnKfSJas
IN77Og/lwzwGEm4zOBczCtmeTDoTBoMG7NeVjZHH5kRZEmS0Gpe3UhjwbboymoHk
XNGl/Z7rALQO1RZ7MqpaXxEkpk7Q2Ut4sMFpY50JEHRnhGBLgqvffRDvVH0POD9U
tV91YzouECl44wpNaoDCFC4Jns9hPw0AtYGXaaJdQ12ShtRuLUkcLVN5nNkIsVgg
XwG+5YCfV8Sj87qFIUEpqsXdTbcHnT/yIiyaxVZPGShvJWPX4LLCfzsTiBhWsgnf
QHlpf2F0lK4nxvUK7B9SsradCQQxod2GfrcDuzI35J3duua1uYw9Chao1cqMuV1q
AY6S2OocaILZyA5lke4eGtAxqxzZOHFQfp+5To7slc5UaXbVI/5XXv62LTprzX45
FYNiP8tyc5NjYPHW1Cr6oDdRo9kDoM6/7CdWt+QFIYvXcE9Rg1VeYOag0v3rqxu+
rSLb6kWBTGRl3SrGC//Gn+dYhHqOOS50S4x70uBFeEGOF2vGRXwGvP3W8OpaNJkO
q7fROfUOfgEucHOmPu+xUNpudSw7KiY++6g9lqPze/oVhGb1VjjwHy0zQhyJEscW
MO0pJVoWLC7AyQ9dA+EIt4nWJku+WP9PVkfx0m8noowoc1fE2CRmvR9vmP/7j1G5
mawZ/IfYTueD8tVoxMaJpKMERnmZeAWu3X0h/qi1x57owUxxmP6EX7MRLN1zN6On
Z87aEgkKmn9tFqcxYpEZ//i3PaOvAZb30lE2CxzCjOKYy+bogdVh3KkowX71liPq
T+RWVItIJzVxZYj/SBbUwfaoKx5t79jUPIRclUh6HRVeiM2px3nYpSPPSyOeb2Ju
hoDKM9PjB6nMVVnJgQQA+zCn5p9daryia87vE+kTXZGIK38HryVHszGiEPvlDNF1
Rw+i3bUPUmAPmMqQsqC2Z5aBsRf8t6PwT9i/1O5Db6pX14P+/8uI0tN52QZneoho
8WakZGPVu1dPjj/avWZz+gB1strXZ6jlBDi8kbCjKFGWdbvsdrnY4N/oBvs+gjP8
9CnMNzXYjHy1EaSzJ/ElKMp8BQ3hsxFgh3Zegs1yA84vCQ4dGVG52bXk6pMsqiSm
ZgKU9El03Lx4uM+AZhvVV6xk+5QzOzzNN4FlYLA3LJexSj/FU+A0UdJ2m3j17nSZ
97IDKmGEuL/mqdLfHbyKvYFbuKZ7EfE8uEz0d80VjuVOMw/SmW1Lo9S0xZNyOXpn
KyhqdE15qngAGpOh9NHSKg+bnxSwoybuPvnRB4fA6s+zrMW1CY98p0VU0UFWqObK
ubY03iR/XaNj1heOuoWxNIFZmwk8Hrg8AglFNNuUEuDtXA29ZvrV96mHLanSqi4E
w48E9pv1qltVoiub6uy9YGs7N9RspSnZggmfjKcXVxY4i2yUOxK4odV+fmEkJ3Md
4kZuLq0AeLomHdPjhObQV0nQiTzo/3C6VNndLfrMy//fsUgCI+94zoyYiLPz7KPb
j0qJoA+gSeZ0T4NJuOTNbnDLfT3T8EXy6qdbz5dezZ6+VjA72/hoMsFfkLoD6rST
50yENT7w2hwFKE2xguvEBmuYyMz2y1XLDofoh2rT80a8MxB7cHFEbCvk72EniQYG
C/6GcWSwSsXUd2+zjCQoamkEgyaI7GwoPcYtYPgTX2sitl/+K/lXfGvNIvQ1KnIy
6GgDbz6Md+Wj4zyzgBsC+87yBpzdvWb5Lq5OIrKhxea3i+wITTXslW4h8JeMCUQg
jxBWsGOuMhKSREQv2C1cO/xBl6+GQmRMU/9W5PfrfGFZK/6rWZlwKHjnwggYjISO
q1sfDjPyLckPiefCMMne/2TWmX+TMIkFRvqMbQ9+yIWlcyw3qchISsefa0ZlqkzY
dcLL6eL8sIfr6rtD69aG2bIU4FI2UrBaG/HlPMfp/+AoCR6HjHX7g8YG7IKmBIQB
WFEPJe+tLi5jy96HVjKRjx5yBGhrPOIwiRrtHJZ8mdsGaM5vnbj6a/TgqLeCuXlI
WSPlt95mPOFhSFFiH64kAxVYX9WE2WhX+YikFCLLZdm0Ex4SLwQY/IBACSsNupbb
UdGgEO0nscVAp/wsaifXKIq2NTrlVb7OwXnw3kveOtg9TqE+Cx/o0bIGzLnFOZBE
gg91Qe49PnjM5itKMVIWS0+23OZCkFQO0P+o9D953F/YS98DbU05oLct5QIfEwVJ
Zp6idjse/60oRARVWpjYjQqEZJB6O3rfI9bcQBxZw1UtuJDXs+iOOt3ukie5CBZK
YRfdAN06vceABcoEskbIh37EhITQlDn40s5H+yIl7eb21Jixssl8E/YVfqewEDQd
wXucYzCnb9XmUutt5udmLmoc2E33PAH81u+cNZmU/DPM0v9afRJ7tTgo/fSwizv/
89Q9a57GgnqT9hVinpqjcULBE09UtnM933nwDRcqr3gdFx0c7blSYzK7kjLEhktS
qscUIoXUgpFJeY/add9/QVIiEUkKdaWXyWGj5NPYhD9JTa6E525LYekDmnbLS36s
O52Cp6EbHk+R9gUagWiV8M3YSEYXyt6xGau5gT9dLOHFbq+w585pOfhsWZ6N8ltH
d+ioCjysuZQuQXKwSwo1hmQQVa4FcrgP+miSAoV/bHRqIZM24c9+BiNGYfQ++kHM
IQTNW6vKUhlUaYqUyci2ONi9ehIWZxhYLAb2jXLXqu0PjRKByBgpgOvsWXnBP6q6
1dtxouZeoxhTMvBFPcKuTBc1mdIaCnkNhnSdWdQpzyZ1tEvmKiuvEnIFkDUA1jTn
5JozD8nYIlfmde4LIZpYQcKqh/Jmg7UDozVrqErn8LcPUXG+P0quZ+fzz+V9HfAt
jUfFn/CdXee5/faqweqOu9RBTFPqwOyk7NDxFbUaIXGPuBBHCZZYW8bcoZE6RVTQ
DPmLMEF1zsoB1sG+a8mK/IEyQGJSRL8ioWXI9L7cdnkXNp3GemDr8L34yd37AAMy
ifiKVaMfBHiNXpR0QUPuaeu1gE57QuxAxspQStnJRFSl773yP8gpAwF/aCdb0nqa
wmAmpEjg6CJnDp8x6GMoy3pIRgR9LjmdTqeK2AKu4NBSaYOXStVX6n2TpnxGudWv
Eprb7ymqJB6pNbwCpxO+I9NTVsrkUFft3I7nuOcWwcbmHxCPKYnZ+ZRQBF9Wx51C
Wr1a7GHHuDtnRGVf6uDNDUrmV4Gjp410FWYZ4i2HlrOJrUuNpwvUPcunEMN7r0j+
Zz4vVfQmJneqXE7LM2vu36R3HD3jeDUMtPJVR4p+afX95tU5aiav9FDM9qnI55/l
K51DpBHiuDFhbwVK+elp7kJa3C0cO+sMlFO4VBPTqPXyVDD9rQwDaLy18ZbR8BFN
4UUIVMWrB0a9v9n9zj+LEUOPgZ3QiQKgG9Sn09N/3p9Iaxw+1Y+buVGqxgqZmIqj
8qLRPLyKM7S/UwtFLQFCA/J+kXQ4nGOWGiyvARl0B+mVI0YhZBXnwHXXBMlIZ0EF
pzShE5rzxp+ndG1a+zdZsByWb33IjWfSlEOfgKefyuTMCKAHiwAjYzNHmhxOEfoI
qGrmqMVnAEYRfuSCQO8OAReERaMh4cdFtH6CYU9LTMWdaIHGZDfamsnooIKI8YzM
iu41F6TUwRl4765X4NOfbF0AUp+ppMerimgN0P1olsP0ruDdo4AnSVvJCCIbQT48
emNAXRc67Z2Yf81z8cOuob9g/8wUuQa21M8+UrH6SN8sO1zFz1npvZPuk546vv1Y
UZHgyCNetnVSvKeBCdYZVbTbrGy37zu6ph5VEVyaQe3z23LkD6z36AlB0/SCOK4j
z96Wt0oG1zhY8ziTgPJN5NNrBWsUAbY1wxWcIwyk19gwCaOr/Ic0a1fItUuQ6gey
WwYWcpmRMSc69sIHpeODcXTR7IX2bGQ6Umld1vGdvb/BYD0InFuNoPykYlm0PnIJ
g/FqkHjb7EcaEb+sVsyeWalMfIAct5lW3RpiDsoKR+nu6Egh0qizvBGS15LUpygm
ExM8NlhzWZmac14y3DNamUMqJgZSdLAmAy/1J9QpRWui6rNJhert5KJ4DGRYjSEV
H2dLVEiYH2VdmxFr4SqrF8uU5Ry8JXTDyEbfqgAQhIpFpORtYY5lAFtTwsNa6SvC
UeIRpdVgA49R8cbuOA424Nmn24U+czQ1Ej3Is+H5qYKs/GfkOev9pVbOaI5F2OlR
Jwowc2Ecw4Nzm5CI6xnPuYeCcEgC5IOlPqdN13Hc1N8HYEuTq3NGS7mgyCiLo8DB
t8nNCOW9mz4pFwgKmrZNcX+mWVeFX7YF0iMNPWUXDSwE1ec5erio2nZjWjOvgeW7
U9BE2mfxER3ZezH1QGshFSB5GTc3+hu6nEavAc3UL555jOokmeKKNLAgXNzA4sTl
2WGpaFQkfvlKw8CQyofYsLG70EkPDxHMNCup3RwnzugVT5ACFdYWBQflP29au2Gj
IjvKf7ltORpv5NAGqLej55mBX7JH9sF07yO0hHsZjSs5G6m2fk099GN0EjGCrC1y
e4ILzHCTc9JTczKKipmGi2Ki/7koKUoqqQc1CHnTaM1sPUSfbR81MrDJIwnJgDNz
mVoq1tc7ETjTlkkQtW930T+f0+j9t/BW3YRW/vz4OjtRfd4r4xWsBzQJgqYXYJn9
WRTtbpvvo3rC12V3omKmNWd5CSEpHkUIC12c6nE4hZdt1lIQLa8wDJ0/JPENbIr3
EyKERpU2tGaZLkifaRmun5ufg3f7vZmX0SOhpWgilCjhUiUuX4b20SH8QIslMrrB
d8Jj72Fvopu4hC0KwF9noCfAXencFmtFwMdIkwg+1ZfReRYsN0JMS7ZoAQd84QWJ
hHA7EbpMxu0qJRWMONNYrShAKzn8KzbvoxsGWfHatiNjnGfTA4xJG1SU2+PHnb1F
5799sXhGGtu8Txz94YP5bB2Kh3DPWT8Q6PZpevsW857ocXD1xpKT7KwjK1vJxHjB
IpP2cZODPhQgeJAtgoFL9TzyxvhomeNV5+7qmzO4Y940Pc5mFHkyVrT5lg8h8ZSu
GiZVogzfrTdwYf0AABjcV/YSkZ3H/dABI9CaR2jSt84g79cZyFRo61jcXBRXve2s
o2X0Lgujxq9ApKHzmzGmNXIyByNq45fuTASultY/9oUvxTkwrxkMEiJs4IkBbKmR
Z8r1TUU1icsSu9SjbE3rghSP7/DyzBWtZqHlWuWHxsGx6CZ5bIC+oTQqVgWs0Igc
U+F4SfhnkcDtT/c3P+ED4Gcqv/sNOvmpleO8SzcG6BT9uPvB2x1cCu0O/saKfDd2
aNhGf3Rk39AkGYmwQeNIkjOGur6DHDgTTGkf1QsDgkBWbeUG2JHPEk42nZXVGnnG
p6dVNoHEYi01qbEd8hNAyRqTf7MQ1lbp8BJVFsgwEvq6W9/3pmz7XUNdT+32jozm
geqt0Q5aN456EYZ6SZqmnlX0b3tSn1vd8uj0xVpO+hAVftSX1XWKoH/MHQiSL5q9
TG7rKw2mhTinIs2s1eJ8xEuQZCJMiYhzm4fIROfP5Rvht3nOF4Co12vtOdpZjLHT
FfpC0xF8XjR1IPXIUzR2RDMp3iBsqw82flJ6Ic2eWmmIDlNz1OFryUG69JA43qjY
FZZpbafVU/tmHFGvxZz9hmVdFspa+0Gkpvr+EE2k9UmW8VxdWee7ES+9nGRVoTsb
h2YuBNNXLdzMVPHB2fqUqCYh6wyOClOnCke2MZm5uWyXJP4jr5ygYUm+elA5+4TU
i31Zq5OUcrdlQkszSA22rWqchNeuV3uj+3r6iVX8Vuq3MIrRMZIzZt9MplyDotnG
9Hv+DPTZRqZBw4Tp5UnD4CVGspNall7sSpso5aTLXrax1op1sIdIfVor/8Hiup6s
QyqshcNp94QAXoEfN3wYoFs24ncjCMPFOGbX3GNaMVxy2Drk2F/ON6B8yDtsJMAY
YQdZdZIwQ4m2Fax/pvqateCjGbIZTuUga09OtfLcpqpSUlareNm9ymy24aS4GxNB
jihg0rA6VFv3/kBPqOUhv31LV7QLsu4C+f0tleMsxzfgYp9zn3zVFqJqtybb0hpu
ZA3/543aaHPQTTFurPh2RMISYUrLKiAi0SQfPrDxbJN0EcnNQg//uYENqzrz4iye
PCqnbYfhljaQ7Keqj6Vu9Xh0z9A5mVeUGLIWJQKsx27YvMeoAV85Az5OuT8Y3dnP
+vKPlplbXpts0Ny2KIKyJZYqb1eaGlswlKsLXf5LUZdWu/q3501RD+sSWR5hoIli
uGNJbgxSk6bitbAWOMvlycHACp/gvfFz9YvIxVNgBplAl4s3quntv2lG8HiqNs0k
tWcYK3gt00m93hsuNFJJqvsHlSo40Ax4BgrYm8ebKpcvheIqBhnboyFx4vSrCWgL
VO29R2iilKpgH3oLEkZ5hYZqhEhY98CBK8aV7u6qF6HQVL+PbaL0Ng6V2K4257SO
/zEAq0L6LjXEl3ej6EXc/vNk8JrQjJkXLabEiA4mh0vRXST5ckKtbPPk2mhdg8/s
EWpmomZefGpe4qyp0b4YXO0EYF9tcApDQ1hTX6vnnF+BjaFFgcT+2u7XlJQQx18T
kid8MTBkfjQRBhIUoXYReUbMoZDydvdy7xMqFJ03UkvBY9Mgixc7G0/7dAOJ7USL
Wy67ypT8Lg6LorMEHEa50duxSvpfgMAWLHeSVFJrMBWFwgdjHMyn31Ut2RxJ1FfT
AoMmgUqbyx12TrfGdbYOYiync+7VMgwt3w76U2tFoZPBeSJln5yUiR1Vr2lNE10o
4u6KG5ouhMMIBMux/3jzlomWfRn1UnDP/ZNQnYnikkfIY/C0BT1X30POdbCgEa5x
39/UN+QBKUdWUO/H2KphGD099sMQwMvAl21GCsweWvjjyDMlD0luBBXCTEAHyZ9H
mbWhgb9lt76ZgKC/EDZqkvyFEiTSAY4MNhnRN8VzzcRUL6x5CpQOpE61625xyBFC
PpJEFORI8Axe0CdU5aJNWLcTbIxGEksvyppc/7RFGRAgQp5RSaW+7QKka2EnSaFG
rTEYhQ0ys2d1aetFFo9W1QFOzpnWurquC7lGDBtU5p8Qs6UC9YlTgrMpO61geHGp
wuON+3LBScbYY9f1R2HdE7ltkNZLfh74DND+SFxb8xM2lPhL++dna1XbfiX+9x7B
x1ho/k4UU0Ls1jKA3NseEXfQeSSxW3yw5PI4A9UW1Jjq0ICLFmaITeBw+c3uBEUo
dXQRPsJMn/6VGh0s19FJ9MO2Q1El52Q47d4kkGMrjL8SOJkuy1byEGe4wZIUOv9I
UwCV0QuY6iaHSNIWbsDEna5x4PjjR/Czr12As40M3kr2MR8pc+B8z4FrXVz0Fyah
oNbQq3NI8ZaGHVwfqSu4ok5e5wW4gtb+DxH+NOFTc6HNH0//l5WLBfl58zRixMBo
Jyxh0M4mZjINOPYB4JSo9WHVKordy4oYd0wSTi7WiyoSmykH4+qEi+artZuOc43A
3AQy689PRrCXwADq9gb/ExBX/9RQnwhR8ftkMN0C1OZcJJljn+QY2KrnP2fOiJX7
UHZg979jQbkhC+s66hl7+VjLNpfTGnCSKqYoyLyTRLMsqJuY0p+OFBqvY9DGRSug
dROICt4PM1k6yxBWg+rwzDfDLLUlDPxDPtC0TRCRxG9DYTGldGyOEmxyqb0SSioM
31eJEwO9VilQFY2Gcqijgg/8jfZZqOhNGxb67aIr2oyt7hfOojuedqC8vn5b++Wr
3YcvfNTIa/Lfrmq1OwoDS5hv5Rge/R+NhCS67mC5IW4YxsjlHGlHJS8ug9+Es0KF
tpZ1Byo1Gk3IBKfRiyZTjp4DPoVyAkaSkUsAEuzrB8mcm2k1t3Z9q/39V//hkF2l
xoZ5W2z7KL4j7YxbYSsOaa1VVqiTh1z3yCWXezB/L4JcQ2bLH+IZnYhdXV3/i7qt
uiZoREtMQ2E2m6UxzkBUFrxaMn/FHNtpyzW+UR6vmCQ3K8Lda93M6k/xs8lTWN5I
hI3mdEGIqgDTFnHrgTUZjlLPFtZi4cszNlmoeadWynim2GNxdU+Bl/s0ixq2xrjU
Pl910NNkb/x9Ew4enpBb5Ln1m9z//VZIQzt7pwBrpchCjxBooNOC8Ow+Fyt63Xzy
PxYHmqLaH+7aQYyREJEDCRRzzl4w/mjzahZOG/O8/tY+tf685yuhNq+LLgssuPjM
FxpS6DX5l10IIlz0NRUve8DC28v865AaB+Y11DuqhxCpehEZi7E+EryiXhCJIjy2
rK2X5u1mMyRo/2Y079RdMJr34lHoFoVz4dmU7xHRzTXcqF3A7R0HFEEO841AA84i
H7GRYk3oa7SbX3+9Y+6WH9qVvGezU2TzXT6v1+oocVscJvv6COhA0TMyLzcPPAJN
4hMLdMYIRlJ834ei4KiF07U8UlmWs0JJJnbryps088htuDlYZJnEKmY4Qsw4M/7t
qm21GDdz4V2H57exUqbywYsz9TH2W/zzKUlTqraZramkWWCPn8Mny2BotXu+UbeL
uUbQ2APVY5qGJhO/auBti7LFbPcDbeECRxMe+UYgATsgHU+tRwsjezCLbPcExSw2
Ump36Xvq9lC0grEhtjtj1gSeZgkMTfeGmhVX0+GwecIS4RwEV0AKmO6QAUictN+q
ouAWGoJ1hUUBfR/rU634/e8g7FbTYrQ54rKpqDpU4q28R1uaEv6ncpLt/NjLNS22
cjHEr/Y65Q6JFzK1SKTyxD5wS54td4SBQGCn9xjHcnBnHMeaEoU5yFRFTwo9sdnA
RWDJbsoAQE7stHVrtWAGJiORGyB2PeG4/wa+NHHQOCwsSEp9PIz1Wli+RxHfRz9H
bIcGGb95urhQYhEw9t3aP9UYNq7NvfVC8KrslwhaGMlESUSaK4AGzZKupnKO4TEs
+gEdu4DEYxpsW8LZ9Wx2p7Zgq0Kn4m6GlHGhQjFGxLcpOB8P6UiRUbCKcE7Lgrms
UC9JpzocmKY5cLCuKJAJFWI0/C3qaFoEigzedzqa0neUzMxTzKI8lwnMEUG7uOIV
ZPQ2vT/Zq69rd7rfLLmWQgRL6NtJXkY5s9SvI2FKKAmdasZuZXfZP/l9VXewd/s/
HLPfMnEeAJK3IujU9uK8jYYzUtciLhxnaiJpl6MV2mQkzpvElgVYL4jnn8PcPiYz
6BtBYBArvq9MiDE6r7j3Pu4HLwjOlMcd4nJ3P8Ofm2yjKroP2ogAzymx0aS8VwmW
JgfNgwFHjBknLdM9t0BZyVOS5e8P+PQ5xc75oqsVYH3LAq2EVaySpODMQaBx3geY
MoCpE2ESCez3RsauyMU0+59jzzAZKO49OLbfuSAdPh9CzuoDhrIaUBGL9jVdx7Pm
qoxzZ7gm0H/eqTJPbpHD9TLxW46xPpD+BlceAYhZBe72/HolvTJw7uwY9Z5xAERv
z9IdnTociRM9JmDzr0w6dXN4dPkGmsAiqxVaNW5HApGvBdAW5Z311OYHIwAmhvzk
DXOrzOs2qcNFL/2DNq8QcNC4seFSNZOnTLhRHLuXdS9IGjayOC/3pnaeL/cnRkLV
Q8L5xtn+HP5kdEe9VEDnNJgbG3G2r1j3dFOJPxRkOBPSAm9RG0fHbCBhcOqu+qKd
vn987c/A8RVAzESCMGReg8f5mAYSjDk5NshFMIuNjmluMrmv5MAueGk/mG6EvnqS
5C6OraKH1uMHhzyR1Pt6W61W2dDfJHBV4z+0vp8NNYwfdvf12jVT1a7r+XJAiRoQ
2l1hOhuacl78ec8n+LIrUZMa0TA1ZEwrFT2OJPrg2x9jXn8G5O1wD9eKQivtDc0N
UItbs8DRuWZ7jHljJFZQyQHinP9Lpa2zosGeGs4Zq0FIgAmKBFqrWzxMwOCBN0+0
VsjCg5aXT6XJD5HnpaCjdkLVY32G5qwVLqssUggay48PbWx3Cr0HmC100MYyczzM
NR5FojgqwfuE2hwuyBhGmJGkAA20kGy1+NQU9bX4v7TzdoOKiO5G2Y2+/GyIFwEV
QWqBTps6tODCLnZGYOW+wdm0+7BA9njxkQoP0vf+kCqr3F3GXs9svJRlmSON/YM6
YRavTwN+cBtVQH5u3UerTYEMoZVJ4evy3GEZ3WttZRbCFZsYiG0yg06O4nuyHPYU
fNm7CX/9PRT8nVsu2SOC4nEJnEY390aqNHv9BqqHea78TCOI0npldlU+HMThrCwH
HGimh3mS+TSooIS8lVXQs79N473DAJkrUJ7PoRzCRmwUCYByE4PZOhKMEzwSV7Q7
kM5JtHXiEnYHsGHoJFyqHH6T9skLgWgg/JvX6nD4KExVnBuYC3jYWwvS4j2dZAwt
vtWAdAv10xC9fNrCGBJW8manLxGgKH0/XGp1l7yCibJvZPYrp1PeRdfKRF0SdUxg
IR7q/1YHmrMpRyNzJaQgPGciqiiyE5r8h6GtasIKBbr8EFvF9Z5e/ZSDpMCaIpwq
xxMEcvAMLumrboCpe9XOzkdW0k1gOOnXbnr7HMVbbrjM1/ZrdjcXZdc0EG0leei/
ACW1fyreKHGXlePq3av7Trv7QdgZosJk7PLPgtT2HRMNEx72L12tqkRqEqsK7Q59
Mq6oDFKAYfslD1K67rwaxmWMd5ZehkaeMnwXJfLeQQy+RM3qoaGQHKP3bs9tT9qO
vCGXQqR7EnwZXzWwt7OMvcyFl52Xtn1+VwlDfw6U7oJyly53bNMggmBaK8I9Sg1B
Xb8pB+bhnQoWZO13OmDiUeCdzyrw0XTfZaXFt5fTUIqxkCUck0wR1O+56DjUiVvN
YSaywlPXCoqFvpNCwFtVrB41ctw19MG2dicPjdw8SCF+Gp5xV1Aoh0KkGFhgQmW0
KArCPnlrPRlhSsXCdMmVcIVoTldCkp/a2o9IgoZ3xiulls0UUUK/37Ybro+CfKKr
TivpLUOuhkc3rXtDyqnQa06Uao/2c/OqLukIFZ8ZKgf+MZyPKUsbywM/upYRbVqs
DVL+UVm8jzucH+bTkQlHXl5fBHmm78NrhvPcaZ8kNjz6h9rCs2qVnHwR1m1ghAeD
MirEpxkvJIRdLp940Apqc/MKEdsF4NnQpgiJR0RJPGFNb7RI4WXScDTEQKFWy1eu
6Kvv+Nxz1w5ox7YtunGpa0kBJR6yb/FbnbaADofB9QjdKow0Sz04LTM/Z6Ng3FCq
ipaDoPHilBvX4QsL4Z9J1tQvEjsMMAhCaCq/F0dyLmofHZ/agKzhDEJv/b9k5dhG
btZUb7O4gE1smHK639IKKfClnQJqJS03zmbb16Bvu36nrlOsaRVYdAvVPzLeVJIu
s7rK0ZP95XHvyfvUEEx68DYEKztu7cmiEaMcnOwnEau0VZLkuOMYVebwMRfxoGww
aOP528RRBBdCxng+qrzrETx24jp+l/tEvIyPoj4dp9qzP/atlRlE9VFqWL3R2iBw
ApBXE8ww1NWpa+VpxSm9BanE4ie9TKLYWVhtvtogXNWMJm6Xr0cWiy0yWJ5hoHla
23gXqoFKmaAEnGfy4lbyItDonCeu+AKLOwixnWjnfhpPdJx19bUY2YThcFiEcsaI
d2PZ+2iIcYI8ckLSp8MuVRuP5Ia8KubLbCv09El+eC6qoxW3iF/gAJ8dVnaKMBoX
v1A50FechHabPQnvBGmMjec1KvxpkZmwJmCUBThnFS/Ji3dJI9NfU7M0hqjYP76H
dUiHt4CHYfajYIX3QrBOrPLDEqG37XvkRoNeH/rxvT1TYn1v5c3HLCJnZFztbjST
LpF5FG6UJVCHohjIoyEqEHRby4A7yqC15sP7u8cNSXz9EYZ0n238dIVkga0TSxS+
EXm8y/hf9UKTLZQx/KrVVm57CP7sgMBVa3JJy5+2TSU0uqaiXGZph2xgZ4r5nAmq
oMHm2NU2rGxF2EN35apSbrmeZeIsFPAn8nAf1Tv4tYZF10qhxTUMyeHkIg6rVCbb
Vg45n03oK6BmuMzkTF+wMDzI42/bGgsC/imO++SVFVFFGV8axzrCm1lSr4VQO6cQ
K5HS58JGMhm8253IqsWWEDnNPCX/HbWiYg1obXCnC48+iEE3Ziq1w5ntjeHGXgP2
hElKPWkY2wyX0sxZZYqs8FUFQoiXrGakeexSlJywgc22rul3trWWX9AaG/5HD0V5
HyeF47m1j+laivss50+KTfE8UEAPPHxOqEYrYOeWSCxbNChnQ5WEHzI1CykL5IHB
4gioHk3jRGD9tGIwqn7Bv75WTsRqzZDeGK1azN0pMoYoYrI+DCzhpkdpHxnBU4+D
kFAfqstyhFSCPYvNb9xghNVY5KYZGsAtMO5DuVI1R7IEBjhA+gJjGX/diTLLE4Hg
0UzR5pRTdKYfih9rWyVoc91Vt6WzgKC1pBbuOESkcTrbJNhDRL6IdBSWqLyJ1UNP
lZ1amZjUvPDSOxWHSw3lajDnwzkb2vZ1s3E2+tFdcWXgbkXIb1dBfqOGprHeU6/A
t5sxorjA0miJ30jzHM+w083pvRARJQQQoLck76NGzJfcK0v7EfiYx373A7pk7hsv
SaDwfL+obhMvYvrex6/pfCal1meUJW9DWxUjEEEz3wXsSbgX1Wj/qtpQR5coPayn
r45kTbcUeEx7ufiY1nnFfgIh/vbHSPNZUVq+xkwZ/PPjSTa02+RJMiI5w1MvK7zF
vJfmxGhN7Xsg+5ai6nHHn2JBVugW9WSfY6kguEfhh41r7/HUDrUFatyeWTYHpVRP
/WIWRwJb/ZinFXsMt/n4vLMseM1g+pZmkXQlz+haybGh14TarNp8I6ZvLRLXFlsx
Gx/yk9xKs3ClLxGPNxcYEkU/H6fDOSDZ2yY8xYYCukzDmqRcayAyrh+Si0eIkOAT
xoVTa3//z6Mzj8xV2fyY1oBv9GHmANuokFQWKAJ2F/HmPdq94380CQR50xAy9Gaq
y9zo5wysj4g2C3agbaWGxCjbIrXm6Jqm5ptGtzLtmwDw6c5D7hjobK5UPg9QfBYf
RE3z3mZD4oSYB6w3n/ru80LmwUeUryzidUNkKAA9/b1+daW+qbnj0xA/vxBxxR5K
Sleyh/+iDCGFe26LCUueY3jIveIiux+f7u1mx6HLnq27wHiNghypoxf25PpdBQtp
SIY8etNIVkFU8giNVCXr6fQ2fBcQr6SN9Offp5wyLZcGbMDqqS4E60EhLa7Cw9/S
lXGqUcF8lXUiACPnh6YYrqqiU0j/ZyDB25vN9VUC47Hu4bIVcPX7hMg54YNR955q
GMKUt6Ad0xuM2axA0ODWz6RGkPIZAakqEcW2Ijae5LE/AQ4NBao3KWgZDDCHzceq
Fq9vavjwy4UBD16munNHRiBQHet/KNQUQBLOL+aQT2/T9++WSVib81Wdpqjj6z0p
zihZPxdSFiFt24qG89Ozfgoq5wEs9jpAu+RVz32xeBIQ+dVHwtSKXTrSRZFhF2FX
39go4+dQfH9d8AzkrzPENcdyeb5snbBD+rfg+tp5i3U174WCQ60RW6ZJeffoDHXH
+7G1fyBKvb/zJUmSOyqX9nB7t7B/5e5AxXCwz6PCEKBZxWcP+xi72+/oI45+5neG
0xDpBWfhZQd+BmXTvbiWBV3bn3rMucMoGAafNDj/GFI9Y4dkWrTnaBARMlfsPTQf
tAqKH5qVXfe1vu4GqGt14WwIxE8wHqCHvmMDD4sx7el69LwiPKFbqrJgL4ecYT/P
Zb1apIBoHmGNG3yhbIbufv+KfoHDjPLQfiy9IoWUQwI4ZVn2WIW3WSZ1AGAYsRk+
MwqOZDVgRuutX4/TT/jnqobuN7dJdeRld2I3qLVocBGSVuU3pUnYu3ycxKFQ2bL0
hxtU2xRe79kuSDERYVVF0tA8OFpaTzXAOTxb4yTZw9/gi86pkx8BuvCT7tOTrPaR
UwDla72FKMDbknfbreucuA+C3NoMGmWKueqeaK04xiVvXJgob5QzD8BAxhM5TbnI
Ffdnjo4HnLBwoMt2zK5Nm5wH37XWIX+PAkwypJo+d6VYC589G2tQotwJZKMDkHeb
mHjUPFC2C2XWkK7/zImsiOD6t80NWHyrdiWfpG+zAFRWk3SbuLhvu0GQTiuF9gJO
b01Sukw44xaUeocirPUZMJk0JCi2ig99tITesdTEXs1gjZSuYEozTglNH7XkVzrB
eIlwZVS6WJ0o3DOeuC2dxil3FNF8qPcdxmBmVr9CxOtF29G2HszMv4BPltofVQfM
N3OgWDlWEttQz82/tpcqgJsMDPliZF8jHTCFrAERxvmWuEBrZXv2YukC3k0CXNyX
wxya353Iu7IY18miNUU8YGKQqk8nAMktXxt6eVhR6o5gKBl+65pwOL7Mucs9U1Ab
pJjSknyNwN6uEao1n68sti9po1kLtEk3HmLA534+uGpTsBWLoTWtfLdaF1HSKv9T
lusK6vrNz9ZJ371Frd4k5OYzSJgN3NDOaepM+qey0uymQAh3WVZAdXkQxpprlMGu
JOuaBjBHGxw/JDeC7S3YbRmr/FMoBZuHMat3p8RID1njz/31H+Y69vY2UY8E3EIK
uw1sY9PW30UeQWedkzXC++UEDtOUwvmSkrR61GAuF7LxSv/NlfAUmtMRGIijsvQQ
QGjL4JVy01UvNMxjoY8PW604dNDJSDk544xq79gBekf+H3zSIAWT1mZL6pxzOWPC
Vdcpdtr2xXlZ81v+JkntRvuN5NcNfsgoQhCU9+lZqlqsKCZiB8J9vg+lKxnk5WLi
+2Q2NP75YqlGQHJK01qCFb3s4VAvolGi/r9nY4HNvDbWG7/BKN5LrJOT7CvI+Mno
xWCpv1xikR0oS9q/b+zG3PJigzV/aPAqfNhgBXB56tARIbDz0/t7AToo7/UM2ceV
Rc4jKpOAW+P9G2flp/EridawDuOGXseSrZFKDHEOuTTMbwa0OA77aDzrk7K+ucKP
nP3HcuW7QfDqqRsECENVqSWa6twnmXuen6FjP3ZZ1POH8SP8bJRxe560W+kb31iY
h6e6FGNZuYYUTb8i8eLcicOFcPKR2pV545dzuItanYymQhD80x3NxncOX97u88d4
57220ioo+F0ZIxHksRjUeLiXMn2yQixWk4OiiKnnmNRSYRRayQj8VZHOiHtaVH6x
0w5OG0kxTR5zwINNG1+/cYDg4ejYtWuUX78vR5aZyRmWBFzbraXWtXXhAYTBWVNV
so9ZoVHSyB16yz/WX6weayNxH6sgw9T65x7aZjXoEjFM29nS0bp3WHvKCzb7pDaw
i7cYC9f0s8FAG3QWw5Dga+LvX1MxgGUtfUJL7nAIg+0zoFNZ+yU6EFbwmNBkqLjs
+bimMqlgCgoSX0yHBVDBxu8wc3koe/vjh8S38iJoxZ3hv+Pil4BLkirV09SM/7e5
JXlzi4of8uPjXIMwLxJxlQFqbC8rOHER3lcmeuIO8uwb1nfhM7x4XInrvAr/nT3s
+aVZQSZnuKbXQDS3O+NC+4u80AEZRvvOsQgJNCijNzxuLICel1gbrjSL03ZH7s3W
4Dx7ZQBJHB8IAWaV5zqoZIXhZ7Kp1Z5BJO1kEyKpvrh3ud0sXcz6I1vJo750Q9tw
04siHf8EAkBNLeJ4IXnRd1DmV88I7AZrPTP0rQ2llURcjtKJC66Hc8RVHyFtR3yf
YNMFbrQR82teTddQO8CLhqghtGlEMqHjYTjHvnPy3EpxZcgB0BcKscJijNGm0l/5
+x0sOisaShlRbMIVtbtGrD+KL7dilTuChWhvYPjwN7eoNumwhIeWyyOO/cBYo/Ct
7oEYVgxAMXlm7SQ54QnpI4y+PoNmT6YugH0QkEt5kBbyYQcl0L+6tCKm8XX/SiCK
NTsxu4m3uM9vsUafK/T1UEagW4x5xFIgF/roXdMvL8vScG04Umwn/C/dJNDzZLez
b+s9o92UK5Z7G2jnVB2cJcYpqtU/PFWC+Qpq4nMjorEhKgB8l/5dsSl3Gaz7s9Ek
vmOW4lNIc6HvsL9COJFf2O+FsGaNF0/W9Fzkefazm6zMoaGAFucTXfTTjoMhE/P8
3znhKL9cGYg3eHbN1vSjNHsR61ugKvZ0oyvlMtoa24LHtrA+Xw83ZJai3Zeu99+i
yQtgkXIYzJ3oohkVXXqmFCwMuVV7zYo316ltcd03stdhDGKFjaumoeKNRfi7U+B9
dlZ7wI6ghnXt7aB2hAX1LYRCO5OrnTJFQOlyogWXnnXsHhv2YJl0vcPwdjJ7mGXM
DdjnqcU4hwRrps1or7e1k9Qikpj6qr+Dq1swVsHcYY6H6ck6PoUkB8DyguLJ6pFJ
vwZ3fMXg0eSpfKz//r9qX3myZ/4c6sQXHY8eesRpcrNaRDjv6k7wCdG1Za4N1JA0
/ItGzBytzcswyEAbu+8+aYZZJJN9q+YrKR7AERmWSn/JxP/gCX3bE6f7n7P8URLL
UbA10R7/ayHTYIUBsb1ESgnj1fR+Uyh6tPKL5e7tMyhABZQhcv45AFfu/MEc5CFf
42Z+U5OzyjlIs7dk7IrVoWFy5b6dg0PjQUIZiPWK9pyDRqE/PBVK9SPlqXmkiV2D
vle+NifpqCx3w26J/7Pca2W2hS7eJY1qTtS04Az494XBFWTh1+dVF2d4HGgQ5+U9
u9+2Fr4cpoef2xpns3OOl2fPj96Cm19/uKmVtkX0hBE9QGt2yWdOYKd9R9zoOZOl
nEKYkt+KMHL2xdPDKEZoSYAZpM/krP7cjp3tabKpW+zQYWPRIQNsdSMWpKH0kLrg
2vxxzUTUXZopvRBZl8gJyEV4PQjRkCU01M+r5Ugmj7+VUGav7Crtxek5+bu53SVw
4OfxKBCVHnnzPCqedkEwBLm+aAT0R5pWVcMnxfYLfJ3QOLvML4ihL1M3jlDFFkcr
xupbIk3FmwKCrGb0S76Fls0HqDJlitovQriWcUlbbskCPO9nCi/L83RezQyzSZ/H
mvOLAgU4ll0ZCbPqnNtsHExWAQsdc2kVcdgr6BYu0WhEHzXfd1UUUZehB2fUMLlh
adYdho0Rrvnex64v2q0AOmpYkM4vPlNI+wK+06GjpmtvTtSW+buD3lQAHBySBPOp
HOwyU4jAfhtZ+fSChiDoOPwNC/h9Rxz179rpOYZUvXvwf4mD/q+KX8X2GkgcA4Vr
1F3v+gJihF/VwrTtJ6pvEjtkTjcsmKcsDX9YBptYhtaPFEgHRKOR6QvJemAgR0Bo
mNob8RVy7tIsK7/RP+SXcKmaOP/7p/LTZDKuCENfej37FSTmZtqE4Fcw7wlV6Bh6
6AI91NjFhQOB7Sqc5xu6aF1cpB2Ff7RPAzciVpARZ4OEtGwWnchTt2O8zeaWg9If
pR5tJzOY2NKAF7Z+HjZTQWI7c+S0T79bG2StIGQcyDlMNJxwz/I0GYUYPfq/7rNZ
nd9PcxFnTpGom+EhLQR9G26n/syngAsqs+9/aovvNUMNqsTfDC+cSa0LIngfaPgD
skGRcsvgHoqy5KkvTgiHyMuuXh2C7NAqCXqgArzLLoJnMEPhsELvcPGevz27KaWr
DXSgZu98pvLM157Ws1r/EzlkxJXDzDqY2LTiff4BLzX9lENqFVOSbsqTEfFjSS6z
yC7krplZ7bhvLx2BoxUPmhR1gS47nU6WIbeerSOyNkvaCxj7xpw49o3jDxcYzoII
DDBuMMSMKYmF05GWcbKuBuiYlUfk/putY8+imh6pFmcOGrVoFJo5WuHb7dz3pau0
6UZpl9azB9r/LB9v6cN706bVShZDwDiKMV+O58vm3BXLkkVBTdHz+R7atHiY9Gja
tTJpaopQAYTi1kUaUayRcVZZPHUQJZR5Naeg/9iSJT/OBXwFSQ5NaiyYE1Ok9C8e
lk84BogE1Ko3cKoNep4mkI1TesCY/jpuzJAE2VTDgtOQFNqzDOldD1d29gM/+e8o
8Jd+Df3YNb1Pg/QVoHZ2AR0CJOvO/XD+6VJX3EXagkTyD/7B5P0aX11r5gqjuGOk
t8cZP6RcatXzaRgjUqRzJWCUonsghI79mTlUxpqD+H7mf2MnHA9BDwoZboWeqmvu
8g1RUTpVhyfum1A5ZlDonGBxZUJO9vTuj+huV/Cvgzjck9W8zlGzlv8Uy3ZM3jes
O/iedjR2SiexNvp95dO9gHundg8PAIds6SSKob0mvZBdZ3yeTbGAiJDmYiWR3Ajd
vSQz0zNUuKwu9LcS10hVFLBxIKR5d4DQ6YfTKEemWsY5QdT2sIbA+UFRi0duVYJ/
8N4gUuZPGgYd0vvdeAupFjtrSqzMCX7YbYjRJcBJWZ/qbcY9MgszNX7uvFNIiI/K
iyWw+LjmJfdm/InoxHiLz55VftYSEghCd5wJvfsPdjrP8wTS64SiZmDA8rWrn0HH
tI32OzNmSLc0mrKh5a2i8irVqqiWiLPEyYQSXwHrZacDGwxu/QCun9g4At5LVjwM
DLdvEwMaA5ZPhxHf1hXuyUtWN8nKk6XBCTDE96KLCR8Dg2hoKMNSCp9rPN3wEap1
SleWZ26Y7bFtj/NPmB/XAQVtiQ7a5Yfr+vSVpzNcEl/cnHZem6ytDll1sYeJRQ8N
r7cHj3pdj3tpaPTjjEi6849UsnFY7prMnyRPubFKj2GuJVx6wgpc8m0qAhM64haT
puI8CGfg2Zs3/8LaPn6aq1zcKIG8OwMEHL4N1zNdfOYGShapuHLr7BTKpmTbjoEz
3xwdAD9vT7C8jE8LnojCmFB4SOzzzyIkvRVqriN7Ehfot8TjC61+gzMB/gv3Kliv
l8/czbfiLwylocKLfGa932KHRtCsVlnGQY4spnAzxOm4NePrY6b94igCQJsNJZvv
nmm6RajbutXut/qNKB2aDSTYY+VZ89oK9OSvCnkHzHtZPv4mNconLmYi2nKikDQc
rJd3th1iVw7yh6/hAU2PJc6i3EVpOIJQd4raeInaJ4wj58Jilu3oanzXz1Mk/9S4
9oFauAuwi4VbGOd1+dEhD5oTfa9XZyaLytrsWNcclB8OBGVDBpiCFlj/eYqhVodt
Ip/LDzELX7D6ht3mvsUxECBPniG8attQ1VhvJ6B4gz5fEdum65VR2JJSQEeN7yqS
BZ+FC71GOwfLjpu5H0s0F2VXgr7AtCdjIh+Z0rUYXJoZUZ+fI7x5oHnd/+RI0Xfk
eYo7CvIacHdOARCHl9/20VyiYSYVRINPauY93/l5FT1cCLFicRuM58UZGGJHAWNm
aYU58Z+z65hP96meJOhP319fewqfxRgkaeH+5iIdjoIPj+4U2cs5RnywWaR4dajz
BKK1Dj8LvGPMKx0SfJyPwoWRJ4KiU5tIlSqqpvcPa8cbDdQSkdC+Dm5tLXaNzQ98
JnelOahn0GsSG9P8CUHxfN6BioHQ6EHGlCOhLOI4M52UrZk6iPFilFgZ5CKOIawx
4J1gBnjiUNd39mmLLpe2FE0LsSNFZKK7iHndBuP25zaAIQxZSLJplrKBOCJUaqcB
rsM8nmDNXLl3jrQyE0+y/IIDyz/DbVMXZFzXCo5UBflvVhIMY1QXUpqq58GTN4Sy
BQB2i0F+ErdyZ80s5djLeUXxvAuuErlzkBttTO5fQlXgIur9R8yotT/v/XaLil6m
BDBzw1/19X0S0NnAzmxUBk7VpKM02NB5hXZJIfQee4pV4zFyhYFpKsYGfEW5Skqo
2CWjzI3gX8ctLLXDGCkO1Z3MqWSm4dmZDwodY4B4Iszol1PsqxTtfLQIYRfQ4dDq
0BUADE6l6i43f9bQoLH0x/UAS+nD5u9ZxUMAEbbX+d1thFArdfut1iGfgn4Gn20s
+SUG7N3ocso8+H0sAjymS/WuLfbk/MlcrDmWtc2c2obgonanrgRgzPUhz/aWY5gJ
BfehrN2w3kCWFL+731sjCzcyyvI+Kd5B5+4qTcHDSNeabs689RCDQW3G3MTHfMnc
kU4fDAA1J/vGxcPKprFa8ebzr1ygKr76WM8apfrviKyeq3TGNpei1BQbvoW6Zibh
v53LU1W5ml1AFVvG4/7yJxyTcCM/4mRdrx5Qdilok1NthNCR1QbobHIht7ZQPaUM
CKkcql5f+2vyXlSdFHqF6ql+yovtoZiJ+orcidaMZplc4loAv5ZvtY2JclqxmiPQ
sANAb4Kw3TMFI648mAZqUMZMByw0Dx9t9BSU0fT5qItUHuSQT+HWvJRexeivzZe8
mwSozAwBh09qeBErHgW871adDhTwzHVvYS0/KAm2fRE6vFzeDNQGXyUSLM3m8T23
AeCnN51KKnHc3OiiwlrR+ZjxRMGlIs6PeOsUdMdU1mg8BWHKf6w/5M5g92q4ufi3
`protect END_PROTECTED
