`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ks9qKKPQVaPYc/mssXvmxi9WxWseKVll7WrotNXJ8rwIo+CA5k6ASm4i25emCrMK
N+p3EGPBS8CWo0yjRBruXvxbuf5jNYF2Uh6+L4YSo6N/PNW2i/pR9IBi2riGlqLF
JVZE2AiYqGC1QtFlmfALD/fWQIB9uZS0/rTqnZdnl1XTlcXAuvXqpkWb7vSm249X
TGTiPsYKDXLvWHar+804hFidq7Oasg84kK0y7gMDRrSjffG/mca3Xl/ztyxozilF
l/tZs8KluNzgBOwPbqjtQGnnyw/UU2ciE6DXJ93Ie3vF2lBn8uSdqkgY0R8Sxq7C
TD410pELY6I8CRQ02St4P4GwrVtzMQhnD0wMpJ39IEgarRHrkAXCs4H1i+opuSld
dCa+vuxglLLs9IhgSaN6WHjdJjw3TaKonDfrgjnfhDVZJXCrd4KiNhuWJTllFYG3
FMg4oo63YSuaO4XboZ5FXpcOCS+RkwgKEvThwznRcIc5XGhjbZ0WXBNb1JKD9gTX
LFU5Sopgb3BafSXLlqNuvWVBQg1V+stab1KnvoV1a0Ls5mgFlbS1a7xygx5VqctU
4GewXlyachAkeUba003+K+EMOv4U0x7T8YT6mIP3iLPjgRHlfquZqHdUXjiI3cso
2We3lBJ3uoIlBnl1nONzVhSLqV33CbraabYwwtesKZX4gSoIAQ6gAZp7QIyLHDEy
iTaobZuUuAvY2G4Ho5fwTHSfDf2In+SkdvKMNqURiJc=
`protect END_PROTECTED
