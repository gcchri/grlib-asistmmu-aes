`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vMCBcm6iNPwTyFa1tsu6O/xLULLqHbI6W7fqnmaBF9Hx+92F6nrwikkp4R5IrPpq
2y1n5Ni73iG2x4HXhjWmPhxJWFqCTMjHTVFVwacimlzwvy1dN9qzrRnyYHg+5GUC
JgUKtSJQ1cTcRPNv1X9ymyyp7d0984ctcjHII1MRH2jJQbZ7Fr2YwJNUMB1pTOKL
0ljjR5TZ6NFS1TgnPW++JW4QJfVZxJ3ZM1BJcnw0Y4bW4SvQqXCQwohBn0Mvj40q
eNKNuQhtTXDL8CNG/wjYg4c9cLLSKlCLkCDQE1EPmnD8sJsmx0pznnIyPsuJDEdH
jLBcjZLJaebIO6//VTyS6nXQBVq6tq6yx2VtNZ9i26zukIKlpK9/uk96RsY3IUt2
cVUY86SySh7fTWcmEpR5Cw==
`protect END_PROTECTED
