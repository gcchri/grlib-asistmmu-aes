`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KwjISwiHNuiaqJjrELZYYF8MBWMCTOd0fdBK73TtMog5Y0WUmj88HZkgzr3pWOv/
aTgHJ4EW7QtHBRisqndnQoP/8dBeud0W4Zz57I2moyVuNyK7EaGe6SmcbiTAo6Q2
NsIMeI7vq4uP+vMswcz7DMGIjiOS6VMIbDeLdxUHeA/fRUeHEz9DgeXJ/898VPbA
vaZv1TdoGWGyJMZW67sWis64+CFYx4BvnQ5MOKS587GS3O61RBo7w2+h3EbcJBdq
nb4O7iV/Ku/k3ifJvDX3ga+Hsim/KX9Tnmgb1GoHAi0AIyTeWR+POsX9gg4EdJem
61xptmgN8TU/qzee0sxctUWf7B7RP8d1ggW4J55ubK6Li2DdBL36QqpNDkj1x18R
BixPJ/ugN+HVbBKK47+PQ8A5ujw+S5U+olZFbqPfNuHB//XKVRm28YShaLNblnU3
CRocnm3eh8S45+zZUrDNvsC3bq5ydCivDXBsHrWA+EU/s/8WLYATAOlNqe4W3S6J
WP8NlhoAiMl0vmYfoUKHDMzySSEA99kz+cTcpFYcM6ynSVXa3RX73IZghBce0H/D
rpfIXomDjrJsnbTGti72lhfdY2upq+su7UGVrZIU6Uc6pb71skMfr8jFsysT99br
dydjPiHS4RLrW5rh1ve7fiyNbPg4Als3lNARj+8A++uIAI3KwuPO7ZQb+nS4/r7/
wiZOzhAx2U+URIDz7lWROw==
`protect END_PROTECTED
