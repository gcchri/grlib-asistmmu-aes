`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bpq52l3UGYkpZiy0s3TVAYgkqL7zpwe0my8dMwSDooTqbiG30TTZWuKej3zvue9t
Hwj9lDC5NeWNVXKTUvvRwRoV8Yv6bTYWM/JpMt+LTjaCzbYcNHtyYY7ZgsOHXdfd
7NhfsK+P/L7flL2mjfNxi3HmSGaGPykvKcWQtl30qOqcPEM9fx96lM4HtIJ27YZZ
HPYbN5IEQ31++d8ftc3tdriAw2MyhSJmb18KleAfqoLHfNeeYZvRKGyjDI48tUhb
maoD3s/MeUbU4cMSejoNhsgQjUpQj1o+bXhtfB0rb3Fk8bhIjb3tFj6MOId3+kQ2
BvMaWPMEJ3AG+9RAqhU+j7Yj/te4tagPytnkntgeURdVQ9aXUf3Hg3wQSsZvjTX2
Yx/OAYRXFiNbTAqyxSGcWgl9TeJHaHCyY2Ggli/yRokxrYOL25VKLPhtqJ4HML+1
GwjKDSFfHmFfYaVjC7bXoolGYk8AW4eOAQ33LWIpFh8=
`protect END_PROTECTED
