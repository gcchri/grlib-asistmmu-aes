`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q2DNu4w0ozUrHqF5OE9povuta1tGzZohlN/Kqs8gDy8hrFC03t6XjrFECo+OJ8PE
7Wh8rPLNAQlEl61ADxm6QWTPbr9ZfIZxO4f6xYGoU2sQT2yh9FLV2tDP3+mgWt7D
oxFQ2Z8yVf1VGBlxGm0htA8zPakZhJ/0XPRcYzOD3tM30CimnShMJP6nTqipdB+j
K0hjRRGBSM9fseesc/hRn90s0wXnZNjA0kAhejmpHi+BKmRe/9L/wvLV8DqpuG+d
TeBKNgch8XyRJVRNRMp2hcf3IFF2kqIkHCVlRCUF0O0VYppJyPV7o47iTDD61TBA
qRFW3oimctBZoymYq6oTy4TWBl21Es2gnvz1gvfGJF8=
`protect END_PROTECTED
