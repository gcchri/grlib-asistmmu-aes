`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mhAD6Zl70FVyzVyLWpcN3rqiK6XEe4BX4WYc5LeZJIcMuSn3ZUopY6rcDBdFLcWA
LNQ3dm+fvb+AAay2ueWuOAr9Z76BaxvFfXiUdUl2Ei+iLCxCJpxudFPMtjkmrqXB
KIQEH6iBERHNePQJ0YpI3PJ38R7yLP9BcnhLORcv9VjSPEJveKNCeD93WP7HeoAb
LU61MeEsheIHCenJyc5hv/gyvjDk0b6EFAttpnVuO3z4P4IgMDymTENriMckyJSv
KrafN1Dv773xKkVecjljw5Vw3Xm2KFJMemLMDERo71wq67zhdezvS9YhZ/pSu8AL
920ljbfKu2PYvvW/sqnJsNV1MhtB+ict7GSb5NohQzkjcoT5lYRCUMHSQ9pgsEvu
xE5PLAo9v1CNe3iNUsl+nxQ5ELOPRCyJLUjuPzDR7nA=
`protect END_PROTECTED
