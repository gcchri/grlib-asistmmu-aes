`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
54tvRjvyydNT+v7fgx31FuXNkWXTJQ1nbxXBnj3bHPQvMZbasfXs66yw7GvOl53R
s+0f3BC7OIB403GsY8qaDR4UUonxmDl7hn3w8BRbCMKHHtOc3qn2vOHKMOJkgK6q
DetjwQjtUzBjxleZa3TXyGme+6KLWDYSqW+YWIbtsmwv4s/u8XHUdKOrzBCMC6Vs
6qSO7D7R8YIHsO1r2hvsuOicRyBzSFkOqmvvh6REyyvN1Oj/F9HpDcXCD586jbAE
mMtC1R85703rip6BGFvs+Ky5pxJRWNQxflgvE3yBi0kJTIinMACjYg4qfV81NFlP
3zyxxmqHlOctFAjoWAwC/VpIv/eYDRiS2rfgRb1XPwjB8Jl6IahvTiWTlUQdDcdM
4jx4GbFg/m7zEO8QD9CAt6wlc2tHny/RKEwYFQfe85ha2oOGAsNWRv2WZ2LbB/z5
0Wzb8P4i+t1cD3cdQyuip+MGVvCC0xxn47ZDifZBU3AoHx+BsMid04yQswbSadYr
`protect END_PROTECTED
