`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jgJ6/k0vqXbpiLEF/q+2xrqDKdWCuux3w4EufKu80OfNOaZKrtekXnB1JEhY/qwW
3i0x+idYHp6ol3FO2OJAD0j5tR1qDhQ6nXWBwFt0BwhQIeucHE1u7Qv3HOcWRwIW
XEx7Hv7rjTjXcUZo1e+37GXWVf1b+28w7cWW3C4OHR+I9JShVRXeDMBpaPRdI6iJ
5675shsrG28NCjZwAKhsAGECdKC0iVHYOkofs4ks9iGdEnVI00LNv1qqslQpUrm3
I6QBcXBZZO+phagixOVk7FeO/exxKnCDzDVJVqOS6deq2nkF8lm8oV0UuAVE51qn
m5ok7FPfg70zeG+t1WZSHHPA7nYwQCTeJ1NXZ7ZTtiuJHUGwVMWjD4fWCKsffRm2
wKoF2OJJgU7VI0RoA6xHdKkbv3qj5ZAUOgw2a0oFOwH7b5TPNDX3MSt85MHSRbMt
L9hZKXKpF0WyALHesH5dLKOWGGuPQg05QbDZVmBXdnkj/XF2W9tIBl93T/bKi+t+
awpZsgf5beN5hoO0p02PqnvcIBiNk9ln5uz4MWv998F7H5onglRibN7IsUtczUPG
`protect END_PROTECTED
