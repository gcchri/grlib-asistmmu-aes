`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U6ITIjdo0fOf9/PFyJ76NVH3jnQxM04KvWuY5ds0f7/sWwq9MV0dP39BFlrebLMP
V6Xl2webuP33x2WZ/JLLBayvOy/acypCKXGGH6cV3K2Uw5gTGJS3izaj7jkAA6U6
B0KS/tSGumhpZfjt/PmyQUE/ET3/PCHERbY7gGGC1OJmszKMIeDgpVpDzp0GMbZE
W81nQNcbUt0EIbvCUznoD9puHq5hfDkmAbAlgOvC2aRzQji8GQ0PeivGP0Fr4qfX
R93NcLcnaJ94Eynj/YitLXCDs2tRu7Rhl+FLxHf6ZaAtmQlwJzoAuiM+8xIQoxrH
X1L7vHnCjfcHwV7Ytfc1i10hpz0dAjdq/0ak/EUcGe5VEeXz52jo5lec5n+Hk6lx
ylTMFebCrK2GEg4/qCbf0aYRHqihA8qC6Qs0U1LiOK2W/JQJuERsaGWv4a1M5rRP
Cwv+gv9BVutuWQpHXM9Bku+1ESn16rbkA1AXDYfpcJ21nL8Zqrleup4/A7sqxs23
uvmMisVJ1VqwdxO/kMiCkUEslJ88BribUXd8UtHm5pfOIWiXc6tVL1GqK542TuMI
lJS7WS3ZWvss9W/vyyZl0hPCvt293Y3LHDZNLVbtDWeWzV3kuE8rL3AOmHaMZ6gp
CwcABPx+O7sQeJ+wVhHDn8q3o6Tc1IRQxPAfFdtGJyhfBj7fCD4yGfAq7h/8+UHF
as9zgOr47U9EELQMJFI3k+2dU+9NsA0ODy2nF9DwnRjy7UVZADBqYPhKiwZrfgXd
BvHo3VzYLUW2SefFJEGCm4fiZTRFDLP3m7UOg5h8m673P/xkT5tHVlPpN365b1OK
2PgaYCrg2HTLAnMLwm+sIqsLRiiQLd0aEZc+yzQXXRlsJV2gzdms0LMf574mV3QC
S/cOVTDxeZAXoL3b0MhoD9CA1Jooo3momhXA/T/GRAsUMBpv3Hcc67PZUh5tiLow
wzevKfw43RbRd92de60fl5P07FIVDWlQ2wHKh1CBc7912CFoD2Hj4/5v/YtkcfEy
ZaSYCsJuN9fUsOErAzB7+WRQFOBwLmrxKf32/Jm0vJOuVXKDejX+fCAC8MVSzCFN
uSUtLwOjMkydeSmbHTd2DA==
`protect END_PROTECTED
