`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U5EBi/2DSjR2v3SxRMtmuMKhVcyby5EiuvoxaL2SFWBnn/A9pS0QRcXFxmoEO88/
oyX5HTWtJqJzTcsCPtriibqGpBY/NPSk9givB9RW/BS8CCULCTlOX+wcVB6kU3i9
D23jSe+1g5Eg6YxxwZn22G6lJ1fBWeC8cIrdTVfGMEmia+Cx5MXkZyz149UTyoTf
UxTu6cTXnRCghZYcfsDfVEgF0HDHzSqObtszIMm6UVqryKAIxZ6J+CcUghMOYufs
ScRwsf+hV2jxijNHjYD8vb0GkXFYYrHGrobw2PLCE1O90BugPGH+d602QpUawShO
Uqvu2NTFwOJN+qswcjGWiveTY4/FN+TQuHnIvq5i3detOw2bmdU+T9jMYW69n3jz
GpHLcIJZjqUeZKgPZ7tax94n1Z0mJezMb2d2Tz9okAaTIXA3iFwnrSZobIaQmeYG
287hOgBn2sxYu4ZU3U2KciGA9sO27jCW6H0oSbgN5IfIoLqYMiV+eDtioqzub5Yn
Q973TDarKkh9RpkhzuQyqooBdlvyDxaYadoj3HJ+C0D1MgWvivnTUz3AZETK0scx
6DzKlr2moYE4hCp4grHTABcLrfrI0gnSGFWBKKzAjv1Z+cDKZ9NG4kc8cQkMYNRC
FGIu/wH0DH+00Q2NNaJBsLF1adlyBKfCoHfhynvzTV+bKfAosYwLIuRgDHWuK6mJ
GrUmRJDMIHn+HzDM6ZeCQYIYSa4q5fXGozUC58/HprbmCwQZtvrgBwXZw+viCRKI
qqqO7aXrLzy1AlPZ9NrbXWmSlU2kHuk3UrRbowxTAtIFlqlI2xa0k5paXSSSXD/t
6b1WkrAsZ17bp66B+KO68Glont0htCoX4j3yWRaxY+O3D+tFKvFy1fCYFwEFTiHw
4SK1ZAuinrsRDjKAsvyhbCspi9NJ0iZwUjebYR+97JrEyP44S39Wvrw7q+0byV8G
amXBrfA3yTN50F5H063lYcgWm8ttkpAg1MfqlUEEsGRdc5sjPNW01mApVHDobn/d
+tCwXwpMeogskJ19eNBIpEbYoxfGJp240RMiPh2HcCI=
`protect END_PROTECTED
