`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cBz1WoFyWiQyW0fwEFNH4Y6qrEMU6s1fDux6iyt5gdrkq7TsjM8Xl1nOYRZOkvaQ
st1hoCqH/FAcL9YEBjPvlgQ3fvh56HoKDBrqiVtOz1c1WBt+I5h9lMtgyajEHPAi
Uli4b3oGlHJvKDSAXacB4cqiNB4Gnys9OIdy3hbAxHjtHMlyQfm7de9bFfDkmJE0
b7Tc9zganKkMfkPD8hEHZG6yxe2nvxPeQs4sAqFigCN2sHpA1/aI2fbsSnesqHtw
9ULeeySnvlvAsAnBlTOx42zzWa5/tLKpNAvhYRRtYrHaWCVhJziKCZ7BjnCLHlqS
W/debTFiIXRDIVUY+oAQ3YanL0rLgaqJ+Q85z5D2hbCA6R4icVsu8P3ciwZQS1Sm
iVa0pv6O+ILq5uvF1yEwQAepwM3RA+zZVTYF2Lfcjc3XDcDJxE8j44hEc1Kd+kBw
RXC5nQ3TZEvJcb8rudTF+8TAlTtLohDy93fNHTQbhHQzBqv3hzI6J1dQsV+PWLWr
rrrG//3JqDsgwTEoj1C1wyfR59GX/lF/g3sWdCmQjkfKPI8n4jesdWp8SMGimOHg
1kfoiAjVICBDwKIYirsY8g==
`protect END_PROTECTED
