`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o9RBfqAmbmGath8h3LrLEpgVMPAw6nfv448GQ2z3u7UclloIXM80RzFz6UGxoHT2
wb5IHXJkcpdqv1msrHanjCp6IOqE4JciKxT+VKtLV6isSS1qK1NN/3mp7hMzX9Uq
iO+b+MCcdUZturi39FaC36bCCezmDFlsgRk2Fb7WjAz32rsdsoOcyavtozRHv8+4
jpME/mSoxPDstAY12vmNVk+px1MlX4YPEjyuu36v7Stb+s7DDXS5to3GsjN2IbpR
FJ5CU0zycjMzka6V8ENB3jM+1kCsUhW0DsnRwMenpHvGV6ekJmZDh/m6xQWZ62XH
Fr1+RX8nevMi8DK0oCmFq2MMTXLWY+VnNRPgizrQxYEaOON0qqRs02XrGhvAAR5m
tsNP3ivzum4pTLPYqX92++Mr1LFFq1y0dsB/I4zsuKi0iBtTSXhaln36c9KyiiC0
`protect END_PROTECTED
