`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iDKy1Kmctxc4KYlkoXUiBpOCu6gJIn+sgZUMf/9x2D4yaVZPFh0fROqjlRujKd51
P/ONO2VV4zrJaoKo40wFY42u4tHRpAeOoc8+l31PQzSSeTIRcPGJ6rJaLFqjGt8R
hAxJJnhYqu/wfXG2QY5CQUQAP+L9LSqVn1Txbgrzs6b1bN9AZbX26wpAj2m/WZA6
qBsqrMqxy4ZxLLwi2AfwJNTnj6db8SFZCJsrV6FatyPCSZtX1xNvH4TamZtZn1Z3
m/5LXvPX+s3P7M67WZzxrMxOa9i5LgnVKJmpMi+G0qKsQCftDGat6V2NLzgq7iRr
YH/CuZ9YFllXvmB0uA2+QGYUnL/Kbw2PQrWHu+Yo5AjtadmcHgmzQYDCXqxidbo8
TF/772TIR0a3adXhDlBhcNSKuGRPN09Dqq2PtO10ML70O0WN6XHMxqxq0qxKbTKl
iuhX5WKdsHLo20ra12BaMp4rX915cE2npnZbiloEJZ+pqNWWtdE5jlUnav6IWF7g
QTqFXC5kMoCJPEDyvTJzsNj7HaVMZNvTBbIlZr7n8ZAIIWi08dIJMxHULUE6S0gM
5ZAgeAjyUvKL+KqQ2wT2AoNlsN45CNXz5Gs6nfP1duGcCymE7RlLYFRcYyuJpZV6
3CqgSkYICQn93GYhuYgY+9BvWQk/kJr6B8dpvGlvM31OpwsZXecxvCnKQrF7pPu6
gjtDIOoFkB4hy5i6FoOeiDIpZG3D9LqfVpJrBTRovuYaXkOuASr7V0baf8rfIAZH
/sG9/yFWqUZHPZgzszw+5Z/g3zymkL0czMPuY1nGDbzID6Xf2A0iGBwH9jIbHo0J
iasSkaM+BtMthxmdYY+ehVtc6DnPXq0VKph59qpQ0/d4SGs3J7J5EFVMCzz+y/TV
DMRTHj89lKzg9rPO2d0BPZrWzdCecareJs56h3zbKEfqZW4iMfb+KfFujhua0Fjw
bbjNoACo8FXuyIOsU4WqgWKol40KZDkXhEprc487GbtVZb8rer0S7jRy/sQgNCg1
NZKImi49KvQgRx1ZM7szLjK5/6vxu31BltOljmi8a2DQvZedOSedn00nHQuimA3R
lwCgFIc4YYvokjx05ezsAmxDVsAJvI7Xa3YVQB9FJWnNd1OSBI4afOq3nM0/imZd
14A3rAnetKqsufOIVhEuOnf7loAOErX2YUWZUFhKRh+eEjTB3pjyVeRb+IlOIKwp
FAhYUdQrbFtxoWmF3N2KD20B36TbvoC+1YYqPLN/sZUS/FHt3mynKSpzX7YXMbGq
KRNNorR8VOodrEl6tN1JZONvib5iCZ/tXIYgPPGOIzeWMaBL8WJ/UGM6X58f1yX2
9E4X3YiOVvsmwCQynBm/CQ==
`protect END_PROTECTED
