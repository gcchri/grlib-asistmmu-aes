`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fuc3DebnVXci/xFbJlNrUu3cQ6fmx9yKgWRcdCy+FQf0fQilsckElb6wXbORBn6I
Ux/4C5lxRwt+/pMIn9iJmSyUeQCCRw4O4wvAP4kQ5GCXgt5tdBD4PooZLjTR2pIB
H0GKuK/9rXa35dwm+EDPMHMVKz4zB3BPgPl+4w1F6E7MwHLKQH6xIBJo6u67EGhA
yaS6w1EgBbMBi3/x6cbZt4V4u62EUzorEDfOJqhwhgsG82YwCOB4fDBH7S7iymAS
uL3jHNdX3uFodlZgX+9hwQU0JwDzmWkgg1ReXBd1aPxkGqnDDWKScyTpBGGNcugI
g2EJ3XZ9oZqwK7ku5CBlbxhkpyUTJiFmr6Y9/Gnzl2DeefrlWWT3Dj6ADGrSeVVL
sS/B3SgdtovWUKwkP3Ipzwy2+MfFwy8jAXrHGjOg+5My2N3w/pX1Ebmrksel1yHw
TngIoFHKKjdGBzjAxP5MFQ+pEG+a76bbNJoen/AuAdK7eDHlYCYpvlOW1FI+yiGc
mMMeGleKLqoZpyBOgJT5ewnspf8XBLshGiBJWBZiLMppA/z5QpPZ7jUkpDTUXpXJ
VqZDlTNikN/+ucEH4qhQ6+HhgAfN6V6Yunp2dzGnz2HHUFo2WLETF0cOQ5psUXn1
dmTmoIrpmrrX/OWo/d/C09n7vlD/BNaUmDUgysr15rFSJLXqlCzRV46Sf+eggRGL
kjHTTVTDP/xkS4pDMEl/mwxATw4iDSl5Gg7Rgai0r8LMo5EJVjhfs1KyR09CoZM2
lmBAZPO5aErtSLny3B3FyqQ4/ytZKt3KX53BHjCoCzsGC17X9q/53YW6m7QTrHTu
mes7NVGtY1axJdSCBOxIWamR5MzAU+5C0oPuph4My8KVI3KnJweEoHTk9wvxsY9f
V0FBfJkWIBMOjkbcxC9iaY66B+82ejoFygmwHUS0cbQZSIiTbTRz75ZnwbPKzPj7
Pt9auvfDt7AGkZtL3+qELnVBMv5YepYUseuSdHEKm+PQMvZkZnOW2qASTrAES7lP
cRHQcS+47uYPIaO6K0ysXgakIYTbdlWld4XHYL8uFCwKvxLjfdEpigGcyWCnio6T
d6kcIn++tF2ajhNdSWo7290dcdYc7vLPegc+lSBJ9hawcNFdLu14xn6NjcvLn7lL
GdzLolhCnvkM98sjJ+OMnL4qdsb5jNrqd3VqIfYbfsIfsm/vRr7Mk4GlD0Hlj0LF
HepPTkwC0/LXdY6RfjQfKNBfXPK+JCRlPtuegr9ajQfWHfaqhiTx8RiwTcycAqQB
sfX0OJfX8JfO8W2NEQNws5ijAxLRHSPKz8cZD0LCCT1NTw0EQOdg7FjiT/9tA85y
1Lkuc3bMwZD/f5YYBfk8co3m9Bt+WuyyhF1ntb6XZUNpvJ/imkb1auMXcUSMAYyz
vMyQsZYZ5KIRUXxvINohahftswGfccmIhVCpwp0Xrvzx8Wv0KTpfoLbo655G4pCr
GbsMwrlfxrrMKZHho+ixoPQxDITPJwU4BIj4FczZ68r8o9w6h8kAVqDRKPtyb5bD
9dRXNMG6j+vSjBcfUClxhjA2QBvav9cE9Add2Y7hppNKSviewl2OB/gOn2bllRFy
JvXB6Jkobs304V63BK+JrCE75hon0g2h0wAPArzfxDuuqCFMGn0tNz2k1O2p2MWg
B75OjL2l4qs8iBAqZtw8VmsfWfQSAURcYNZaUJxOUKwpovQTU2qfxI3rN2BgEEct
gH4tyfBymWPbyq7AYEv+1lg8LhzCWSZ4mHJIImQkSwyqFCHO6H+tw+ZfdxImR48g
2INjphzCwpExyGhGQnVeTYNYkHpma3kRwkbHjFB34gDWwe+W8yFKCj0//i0MzVU7
iX7xkn1Dg++nt13ufiaVMN6RDHBzTB73TIpbdv3Q4GocPePuC2KSN0iMq8/IW+XV
8H/pqp9XA8bm8sxqwPmLvtxm67497zzxFzKHkFi2yKSVSpd4bz7zZWKAcj8McxQ9
XRHPfhQ+MVBGpPS2ns5z6CQWHXO/3MuyvRB7I26jEf7ivrKTJVvSWnqnQ5fahYK2
BNPnWkAyxZT+O47VrrHqTN02hXO0Ko55spYAioQJeLY=
`protect END_PROTECTED
