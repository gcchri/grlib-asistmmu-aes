`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZAj3INdHJmenp20aofWJTEW0IXuKGjtN5//E50dfkXsWp+qqenBGJ572OqrMvm9a
WKwMNHb08t/aGp6Ef7Qll6Xxf4OFq6n6/ZTwgKK8LmQngxCm7fjecp1pTqI22DCR
Heh/JpXlQAz+sPJeIKknCdlP8ZaEm/BDuHVGfm7WED3YmRYOGnXddBCN92NPpzit
nWO8yGW84WLRMbVvNoq0pDjJdmbgDR71eHSUkKCWHj6FcitEXmkGJkkI+Og8eW5N
DXhtd0eMWxOULHoDeRasWVJvdC7blIGuj7HUdVcZTGjdR416lrvIn+fsXWjs/M6r
NiO/ixgQVKaOMMCvrX0C+A==
`protect END_PROTECTED
