`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dn5pM8PkR0znNe69sJXMyFE/0A5ejr52+7u7MucTJqqEJxpEoTK1+5xkE90WTNg1
wInZ/6g/87Z9Hc1n9mcnqYtJMbhpyMmDM/OW0upHFUn3phQBUPFE+WfIgmhJV7eE
xVGTxQbAZr5QqKhqjwdhXf6TgsbqxqCJ35va8RCqIiNYv0/rJBlRWaSC+zbzaMwt
WGMYxtsivYfp/kE2/7yvw6x42Q0uqbfuJacfUsV1bN5Z/3YCAdVclHwnhsY8jTqa
KMPdJSbqqRvCUl7Mz4lGSeN6yFhEJF9WBDTq7k0YJSPJo9gtVrya4hcobedo5xRZ
5El+4GFAEoCXYV5SjSCnsDaOtMP4QoQGKlwcR17Xw/xfbDs2k3DcNK4Zwz+Su7hp
l1DU5jnx+FZjIU3bxsIj00IYGB8M2UeRKGiz5vP9Cz0=
`protect END_PROTECTED
