`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t8hFIIz1uSpygl9D6aAI/U6sFJ/TnVVcL3Htmo+kRGH8kxPMQIu1mr6I2i0ruVS1
yCxv0nXktv+9HVOY5QWGQsh0/qhDEL2lLOLNXXwclCZ4m6vOlhMb6qcPF9aFhAc/
22EAbzOv1OPPXSLXFKSoSj6Tu3oodJmKHtzmGth/x5938Jj44H8JPl0UTcvfrfol
1IrvvMNbf/nztGqWuKqJ55JtDdctXFfxFE/mIhJOin6jebaACNH3j8YgnxOVGT5U
On8CHtoQRsXdxa03aC9CfIbE4dzjsUbCJB2U/ORHH9AXtdf9PWV/sh/3vE/K/JiB
KTF4jEhfHD9FnLDZvwfi9amUad90/7IiSL2VwI+V63rh4/d290ClUKm07FW+/jkY
qaq37qxqGuCiy2rf8VPBIhbOmvy51/9yDKWyuLlsc2E=
`protect END_PROTECTED
