`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5SvL9p8UnlPShX7m1Ag8YZ7UMIMyrmNgluZ7mP6MqCw8nMHWiuUL9zxGjyxLiIz1
nuvddDrLipEH6497QYLstYNOPY6/gW/0tjyjinERdoJbQIEpEZQV+kscmY18VtYs
vyjcCzBz/v6bgsZ8XvI11XfWGcOLp7jECNCZrGnK6UaqPBZVA6CTGow8dqz3eixD
4uk4Bb7FApPNquKjUaj3OlPvzdSHanuLJSmcGOBnsSnMyEKzN39tyXDjFWdEexfP
YhF7iBzrAYXQK8GhZi+7bj0sDr5D9i7ansrrZgm5wjG3SKSVQobLYlEQsY/gC8DF
o6//K1CRvEFoDHfJ+2FL33Ie3M1uiQ+Q/OTpheWTDMIRM3lmryzeWdsY/S16TSBl
1zW9KMplxLtvk+ki1odrQeCMQWaC/pZh4mYX2L68R3yR10eW++crEKp4+M3wzQ8H
XDXGmNXv6t5zanFCpHEwpnliBz+9w1rmJZKL9f58n4O61jY1jq9+4P6uC9zwJCJ4
Su64ZW/K691ILF48EBPGwB80WwwXP265KYfM3hNVJwcNU+dSJoh9Nk0D1dXMqJd2
`protect END_PROTECTED
