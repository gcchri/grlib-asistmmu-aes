`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4hwFVqVhKDpi7oMUGqZU3vUHSUm+cgnZsD29QoB05jZX5f+nHwn+dV/WJXZKwjAf
IZ9KjGFdnz6Z3EyjRel+y1YjSoV/8H2i1uaMfn6eLUVi+FMXrCs0lt71NRqo8dTW
qsOGMuofjEBPQrkC3it4VohEk/tLT9CL/MNu77wEN3EtqxlGspwcUivknqX5XyvQ
pyimsAU/PcFM5IOpebyZ2EIo0lhdkTm0tSy/C03PKcSozv9HbllN2kuMrma4I/RB
yyCWI3V8PNjliqm/HGS2rh0I21uc4dLBY/ga6JiQBjdnT4KydcJXvKaEqpkaGu3t
5Gppm38ehsjc7ksUoq+M9HH8YNHNBs1B6e65VzACA+vPz42VCPgsiTIXAN6XqVE9
DfBGOOvHtWQOIQYqKD439xaZKNGRaCn1S6+tXZdOAou5kVypDubWXVe3UMYwio5m
MYdItFpDkmEUzvj+syDu+mv+0ZfrMT6K1+QGPQRC+rbRkpeX3BaUsDfdlCK9NjvD
7vZOX88uCLJz2YF0LK8DWGvw2PE8xGnI5QWade1hWPEMxPrngF8yocfjyhgTDz+O
bR3J9nHu9FDnvm2hGa9i1ucqnsP7Yz+DAgT5Ql3ffPMSQ5xYfWV946dgxClGH1sy
PF+fdrIOsnJ2/GbapeQ0s4snFgk1Kk0oDTbFG/u/IuXThdIrYwAx8NbJGd5xuKOI
GuktA2BBidRDIBQh8wwFacOsJQRC132HZXoc7OBJj9nm5TSPvT7gnhTjIUtw38eO
UyHlvZbaovaFJXST+axr1MBD4TDpzIgdRt8M4pqwA171XF+E6+fgD1U3dpYYtEC/
R90hpI9UGLbjOGx+VtIWi6xZ4/QiX0TAFXQcT72Q0Hmbd9gSPBhBHf2+GA1uXXT8
qxQyRO9q26rVGIXmsvpfygKgr98A7c/P0F3cy3SEhmd5bLl3jAVt5stBYjzEW3+r
hqcjcPWE3BlmXlOKB43yFh4DpvamSTThlSlkkp+qqe2Hd/FYSJ04C7L6+rpInvZk
`protect END_PROTECTED
