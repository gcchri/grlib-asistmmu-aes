`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vDmzyR6VzLbW+OXSnisgU4e3J2WXqgB8iYiTrAwq+v2/YP4SEhAIdEvsq/6vwr1V
A4dL0P+1+qngBt71G6TZTSuOlFcOLwe2ZVR5JGEkeSu/HjAiNlOL/kXPiIAWea4q
sC6tZU+DOvJfFz+kD/Jou4R8wrJ2p9fHY5nb2Y8a3RpIDER4KMHPWsSYbOYpD7uM
TjK3i8ANcAsSforeTJouBAyqp1GCP0qyvqXbzGMV2drcORX0EPdaUYxY4IvMog5L
b98GP+QrJp+OnrJM/AJangnP/CIJ/Mu5t+Zk6IZD1Mn6srxuSwdq/fUE0gv0Y30L
QWICnFpVmyS5LtY/HUWb6NN+E6oV2yLJj5dYfrez2h5FkwHfDU3sMrvG2ptvrZyI
`protect END_PROTECTED
