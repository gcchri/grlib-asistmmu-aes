`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CGR7IddJTytV4LZ9sZ7bGJK24+aqJ+6uY/eS2zPBds8moF7IZXBsvCoogb6wSkY5
eLyBzH5jqkwZs6uBIgotiel4XZ2EbecNbVseGS4j4UnWW2OWgZ+gZaz0xj4ayx9M
C7fxFHnQ/eW9JtWjONxysXWtfo7wAW/gat50u1B6Aztz/0clkxHTr8iviFflddVy
YE6hciY06O4YsdlzYViT14MNN2HgGWH/W8PoHrtSxtgeildU9uvPhZd0DHuaU6Pv
28niB+uaMcZDPnHM/qVYbvvNnPIcbX1I6XjJUiy67OEAe2iZpXj/Q5pgrInaPi9A
t9watZlXOB6cdvHV3fDtI3TiHYObbX/GHgtIhI6rDlYjg/Wr6CxzZBrEcQ1UF9yA
hUlOarrrx2wmlPRcHT5hJAAPi4pvVd+wE/PouwxKnuI=
`protect END_PROTECTED
