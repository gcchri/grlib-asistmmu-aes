`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wDchkanVd7R3Bf+cljIackzwbT5v3kjAzrhQ4wxWUba8M2nIvIBHPAMACmwkzhjG
fWMcg75hIFCu4s4IcVkxI4+i9odYXSXGSMgfD9fC8I0UQEDo1TU3dFLsURxMYTT6
BV/98GeZBJ4EY0VtuPpFFyNPt+iANTxI8YjA9XqL7jnitFgaZBRok1QeVWSpSdQH
12+/XG+c3TGbn7vWhDJqZbCeVB1k/j+ryMgJpAKI+OxBq2ZGjUUUdpxy/t1g690v
UCxUFKpj3eZ/l+cYhEFfv+hHgtQvnZIWAx3r93OkVcTYllICzSHsq3Ww5npxzaMJ
VUIxbKBoDgEmxOaHmkYyf1OhHAF0CTjiCmq/q8kahGRBCXZ3nDA+VwJ72pWnJk0c
TM4WfdIa9y2X6ybwZ/TYPEfNsl5HWURAeKj42vMwvwwPSE2iLgqL5N+nwOJVGIVK
j2UW4cVnB+2s7RxlDMAsTkugrgFkG/EqoFrZEl86BXcvK41aghPsi6ngFkt74Ka9
vC0IOY63IpewqbZZtrugV7UupqbzfJxpvyOlLDG57NjNRdM80SX540iuIzJfnNdL
AjKVdIrICRzSNE0uhIEPOvuRCY6BSFgEilMhWvTr538OgL5FQB8alDUvV1NBVn/L
+f4saa7zr9mgeqfxrxFD9NWJeiqptdMmDCQnnS0YGskVoG7IGLeuVEmjwyhKi1sB
NeOctl0lxyCQNc35mU3J4X+yBhQXA2Ry76zLuAhIAYKRXrDsibHMc9sQIW/t5X79
D4BVDYHjYvF7Pn28bEq3IA==
`protect END_PROTECTED
