`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KZ6fnEwUKisynAgCtDKOGyShMGPX9CdKXw7JQFbFDC/9zv7lqZpq/xAkkqXT/cX2
NMS7M53KcrFCcWqQwEzOJacvCF55INNuQPYczJrZLK026/tt+zrUMcWuKBOR79On
rdidjRh5on9LBE9sgpbYyMJ6HZuo7kkee4BiHT05dJ/TO8cVN3ycZ6R87TaMtyZv
PbF/BRJ3AOwsTkvz7N8IjTDcUB3YznX1ipciN4FmXJV4+nWtXqmMQNvGfQ+px9pD
VDCacqeFj9lYVnJLezBF6iT48ugo+1tUPbir12zC2Ay6XT6JbkzbEX1BVEsqUCGi
QyIVKm7QP+d31R/z9Qfww9iCd0UV6WiT3MhNOtc58gVp+d3pXGZnq9uZvkxkRAyp
ucpnb4i5j9A0HurZdkkOkDQVoUeoTmF6rrS9npdTGd1bnFifnJwoRBJjrvXcY9cF
rHmjFIsEvzlfdpImy6irfzRQeyFsxoZ7S1cnNtFN4BXL94fX80R0SAdqWe7SyF39
Bpp82lcxrBWqyCZ/hBq6kcbVZImcaZ3rzP61VVavyzZgEcMlOwqnYEhJenzIv6D/
FhsEvTGUcW7J28swqHoMAj9Ln/C480pDAe0FQdSZPlEXLJHGFvd0IKL0QiTKnFe3
ATHIAY6viaGMNdVLt0Htv4PEUjbVHCeCzt2N94Ic8Cq9xi0/cIk95YK/pOQsm+kc
XLw5I3yRDTJJr63KM4t/F4H+Zdl4wKWYXr4ZKfX7wTzoxcSzjcs0EXL6UHvOIKe6
xdQuOOGjkcQ9TAjTPmLRdzBCD58BZi2NZ56I/MwafNKHS7cEDM1f0TeCIJLR1z0V
iM9eJcZSkfiVincUsoIqaTT44RMgHV/h96oPwUZAuRyfsNcjYAdWM10ps7QZLzDg
7FPcQv04xjYQgZTNyIZuzuuSFpQA36BY7wcaYzzCjDAE2GslSzhD7lP599HIbUBh
OM7oSQiRaq46GZJK8MwxssMSoNesHxibdvPq7Q2k/TgiLgiQVJLzU5KRvj7vHql3
VOl75CY2T3ZyRwle/xm5P3fV6vhcKMQmSnOVfeAGT2yhq9Mx0/fiEOxjKoOBudGi
Hn0OWycjVr0lcnTs4bw5m2ZpK2pcD2nbRWZfeItyUBOxRSrIXEw9J9zOcTL/Xs6V
/NuRsDmDWQ+dOJH12vUJFnBuPI3EA0yN7lyy8B3+CiTRn62G/UAdjLXvS9gQ7ZBA
0zvOJXXAtds9bJ2mF5wGLRwhfbzUgazicQHKbwFyy66dRIKm6oloTwF20LdPyMuU
+yOMS59cl2myS/IppUOHhzualWZVmXYWtjZBQup9asalG3fbHffsSl+ndJsgL25c
qC7CeecyLZA9P2UOha6Mg/hcvmiNSpWp4EHIxfLQ5MxJpw7fBgTVGOS6kNiCSHUl
fsowr9ezvDFsDTYxBSsgmYF2bq/ZQ2zGEVyKpr8UJVzRPcJ6o+qFnyaAnIy6WFJ8
IgIRbNAcYO0DovXPXlwBYeJ9nOb7QdzeKNGMpZnm5Wi9XiuRLKhxnGcsey7lNsHk
M1hW7E+aY4PJ2jCoTXNwdPlMqL5kbY3YABXi0Oo/Wx1pbnsRbN1kV9nZYT5MAgvs
zIr6blV+qZCUFgmPxAHC81x6appoHIeSUY4I0kwqTX8BgO6AuRojY4lf0WPj9FQs
CAfriBzrU8L3EL4esz70UN0v/3GNe8aYjSAC4KZxdBiDFussauxQOP4vD9G9TVM8
P6HCWH0/NMi0jCWzzbF1RsRMaCNvTQoXXPvSrJz/1pLjKXk36ZYHsLVkOa8EKClb
3yUIjVQzV0l0QALHCgxMLkCdf4FzkkjPvfCXhb6t8EdbqG7MOWNy5uR8YEf396wC
WMgcMOZKl6J2sM5kP+ZK0xL27w6xMxLuaQMCzptqO7DIfX7RYROs/p4KiDHmnu6T
eFcmnvvciPddhEgGoUMKl6Gvr9cOtaR95nPyxTLuP4kmZ9p2dxeIr/O1J+eArKxt
FKS6dC86OwKwf9Q04Wwv9zYu4e+uflRZ5LrGLGVIDHmvQrHtHFyKkZlKkKMhaOZE
g/aROiyjE0G8193y1ayzPsfJuKyogm2iFfXyrvJYKWxAXEeG+OhgplZkCXb/OEU+
t9wQw9AlbcMkzicOtrLBi00DujGMo2GRaSwBf3tWtSouijvUCXMMms9jqtOZ9zRr
bKwA9XEl19uCn0JLQrPiZkeKlWPavJ0yhDDkd8UGd4CTrV5KiLVncwuHpeZabTdJ
ycmPd3YN8mw+Wbziy3QMcgFbIOuuMejvFCGX9zjG0PF6PAzuNawGgbabET0HgGuW
jX2my89As+EoYOkr7u60bfmCfENw2j9hPVR0vz1CrO+fHfepzd7dbQptL6x9mqgX
DLo0RyWDlFlfzBUYESkbJoeXWBAfYDjV156Gt5pKrA1oOrr4Bae5nKbJs7if89fS
Buzg6dSJYcaum0Uu/udngsKBhnzHimlryDCqL8ic8peWfOMVXw4OXeRTkwNubYx2
KkYxH2GEUkdVo0qTGL+Ix+M7u373h88PVA1JZIx3lQNRF71I+Lj8WzQ3qzq3gCW9
uhO6504gPUiUXQVDpRw6btMMUREkVZvoRA4EABpdZEuVsYFN1GIWGK9t7aA7gf8R
pzIFIyT8OgRTyZGgVZqrb2jzOLj/AcDrTP5OVQ3oTk58D1LpqAGI8lHbOtelgmQG
sWQf6NvdiMo3vGg+K+xX7ahYg42xE5+a2qIaqLxw/+MIAyJQrid4f2h4xp/fQoVC
bsPwLq3ZCTTLIN1wNAr4oIhkR6w56A4tJbfVuN99aLZcXcbMm6EruJdU0fJdo9zx
KsJBZpimkCGPvzw7vU7Cis1dEscYLydopF58T4iUtraM4aukmF0xYrnbGnj2s2eZ
mKmiY3ITRhL4/aSvS/RUqOLHeepGicrU2pNOT5cT79FlXSHrjqi5mUX2b8JNNgnx
3p4f4crQGbkgJKk7dUzUzgD13FwJyqnulhQoDYq+Evhorcoxz5iyS1Iaq0rDTZt1
HENO3fk9ssJUwrJopoXFIvXZAkYwcJG8GYmPTN8eJo1mnA88cg3tlJfwTIQgclcH
4s0xsebMI8OavCOhN/jl7E9MHBPm151LT6J9+AFgntFNf0q9YM6kFMM6n3Q7gNI9
b5N6FizgR6ptCxOpUnsX3gduaQ/BlYhDSngc/dG+DSNPyGsJrIpJDpvgxfN0KTK/
0Az6MXIO1w38tbNW52AM5u1OclBPaF9OfSz+OGfzz/JWM7lHLwOonjEILwc9dMWP
mH6FUcxl1Ba9jM1uMzUPTiskhke6ueV6kyPgD+duCXNeoNCYac/tgjISrZAr8sfY
rAnyB48ltxdchNXHf4DD3mYD2gAza5dB/4U7Bvj1GnOhfj9IZP+tw1dFt3dMW+D9
sRi/aO3zN78MP4Wj6pZ0CW2Z0VAoCFFZstDUD1lrcdxVQsx79d1VvoxOmo42eAnh
2l7CSO2EJ83lhUzNJAgBH0N3UBB9iJWcbJNi6W5W2O4IZvsVefSyzclvDfHYVS/t
hzu+kCFg8CRqi3OhNfx7knkETQuhBQBcwyUipL27ZkWky8DRID5YWfHeiWx042XH
97uVJqqOeLcUIe3WB3xzWNjl6KNBoXhUikAjkE7aeXGwNoDjjPngD9WlQ2a6PzOo
hjH0qLGPkAKRuMtnNAtYTj6oiH/Rtk4hIgwQUbdfiEjk6lB6b2ZLw1ljE6SnLuLm
uaRBv9qmu8lO9XW5nkXqlnt1+A3mKsILZ/Paz0Zg33Eoo+xCnTs6C7fq68khh7lM
gWIXVxOF2JKEMw+JXlmYROONBeQFI+lu+h5VaOXn0GHAHTq/pN1W5VcQvbovqQTz
WtsLAOPVd10i2bK+QRzp3/ypD+VmvgxyU9exgt8L8nOP1RK6Kp/QvIsMJ61bZtxS
QOxUEWTPU+loBDeIoguNRJAmNUidmJnejnoxtMpIKTd99uD+WS2T4UOBKIEAUxU7
ndFtmSLXgJs4xqT/q/V+e7UCdtni83oBgWOMYhZ/JK38jmedXItbd1ROFq3U9iGZ
y2AwvpmVlZP1kzn5Vdn2wI+Np98Afba9PSITiSxRnVLNc3LEJGWUZUDf5NCCRfAf
BaYMzg9dykZaFO1hp8yq1AouAwqft/e8Xw1CAfwO+f/YgneY17qcyl4fWjpN6XtE
xKZJ95BVD7jbFdgL14aBa9Ro0gMvweWrM85L51S5nfmrpAEthEkGMdfZZnAzR7mR
9T+L2t+AGkZx5sMeXTqIJKlV2L8za+2eLtdZKTLJvnA90XH/TKiR3b3EEPC9PhIp
GWywsJqN2KUpvd/cy+nC0jf5aFUi/ZJ5zjpDptL9BfZXbqai4X90jWNbJ/YvXUvj
JyoIJEmhw8eJ0oVDWgzCeBdOPLx38yJ6w3HoL7AmUvRNnC3wYsqsPPJtAhH/IW85
CcYnfIx6tfa5mxVM7As1sErxaQjDBk8KW3ju6rvI1xvZ7xikjWE8lzn6RZ7JfGMy
OMXUiyM7+U0jqbaWj/7DZZ71A6t7kllCUpEkJd2wxHmvK9UUFujt+43Ndmers+DF
yjw+4Alc+s/Dj/BrVBcbCrIFPJT4Ml9gWqOLZmBzz/Ff69ymFcTKoomACWxO3r5v
DYqIl5oRIIvTiQi7ZPJz/ytkFh0KeyJ6tdb27l/OcCkHrPxtjmgSGGo+BpKHnryh
jahXmpLSrhPiDziNiYrudaa40WWXLJfCPbAMVu0y0HC0/AExy42e4VjMLwQTL1BG
dgIIfIvtW44lBll+G+yZVA==
`protect END_PROTECTED
