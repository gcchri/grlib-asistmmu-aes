`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pD8hfw+RXWo7FzucmgX/aAwSbeYENtnxIJoNnVuhaXyGQkymGLcg3Ojig6S6L+er
VPY/Y/Rrgjz2AHLilEm/Pzxo6Ab45zdI2lKxgSrwf6dbOoi+jFdkxJv1HItMTGgU
Di29Kba8oQqBZzC5ChLvZW+vYZv2HbwsvbphQvk/kr3qN8GCUf6mjqmddljBJpA1
25/IbzUlxrpY3o2pM8o1LHuGAieH1WXH2vtLcUJxXJv52Xz0u+It5K+9nugCYvaM
+AtmTw1bPIpuozpelCBF5e4Ri+xegidtjjhGZA1Ck6PAeHPlr5Ao3aH9Nc1cvlnY
Nbg2w7QONBe3dpTfKQCn4h7OQgSUQhxujOZrYWrwNcUO5wG2oAifvZKLJunQD+my
mjVOO6Qp4joJahUX77Y0o3vjA5MEvNRqa8qWSVrWAKXB1JbnXYj7YW17jP6b2fPT
v5mHTEJqGmizjbozYHN6fJqMRLQcQ2FyZZY6RBBabwKDKN9wVtl7/8Bzlvv7i3+y
sqygg9e82KD2+98GwoR/10G1wcIMw5e9EWu8OrbjZ07npDtlh6Bft02pN299SDD4
EEVGMwbJDCCtXPk3iHUzzJ2G2Ih32cSskMCdXSgFz2cvsEPCm66dlNzGJvYjO1pc
xOI4602WYHSi/QWhHAhPSlNWlo7ObPHBvsa8okTN4FDhA7VcKHH9NIRNQURsMFOn
RqT/v1kL9toBQTWGmZvM/vr15NPjWGEV5ncO0H/YxlxauXd/kJhBgE0Etr/aTxkS
Bo6FwI+Z3GxHGk8EgogJU3eOFZ0fM6IZeg3RzC2F4OdxWHGkSs/tQ1h/8FKdILc5
FyHP43reSE5EXviSh6RXRUXhDsuvAwzRWK7PPIuc5oG2V4vxaTwPHz/0k4t6C5Vk
8UxLNXNJfJEEAj8XZePwum/4AN4GGszIhb54i7DH+6hMlep0stWMWAgfW8vRWNBs
Lk6ajQEIKSuZ4qaNhSeXTasoR7D54M5uQ4ek377sMlQ0d8+f749TXhPO3MkShntd
FA9T7QrxcgcdAVKAsMkUmP7j06nhTJTZDqqAA6mSPHRM1XEn0iplpB/JHs6P3z1b
KvLRw0kyiR2Jl2cxXd/zTQ==
`protect END_PROTECTED
