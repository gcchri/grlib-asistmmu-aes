`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
730SJYWUTPyAQtUeACC0BtIi8qCJ0+EpAmGyh0pvcXbkhZnzmuJCPD+XOsMg+qcI
dp/cU5xlzXmXvrwXPd55ckHaeHexlKVhW5hLT4lmSXa9jijKCZ/MlmK9f5h1/AWu
9a0GIyL0YIdGDcgIxW69w3xoyKBBQDDxpvlt37Z7RdM5kN46Nl1v7YpQ+rZKiBkq
B97IYMJuthkkkLFl1RzdqKHHddSIyz/0k2puPFdVnvme074yvPMknAC8tZPurYMj
xM/c5KKQZQ08+5wNkgLVTYkmmZV2g5g012QCgtB7HoM1EXI6Wad1d/6aor4gvs9Z
/J5f8qkCq8PjiKhJYg3YLdw5gA3Zbzt6wnQ2A3ST6YWpvnVyOpb1IgJhG5MG1nF5
9SuNpMaTw2QIumLVbEdXL05KzCmkDg8rljEsDari8dw=
`protect END_PROTECTED
