`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kHVBjzKLlO0g1GvHph/IGvVTbTHsKqFe7EwtTHdQRsamyq2JTIg59cursSmaGFov
R1CPLcKkVxK/SUAgQfnENORPxZnOzE4Vjs8VpvT0nY5s/pjvEEcZq8ymXUDsirU+
x5oiTRCriJwCNk6DxzJ/ahIi65S4tWEYKC3pzSO2L89Vi+t+DuG66FmD4au4f10z
Gc9uClUPUd5NoKloW4gG3XGKuVhRl0Z5B2GFkg1eymCqCA2sRKGZiw1BN5GYtW8X
cf7+SQ5fytBW/Xh0TJaeNpz1P5wBaeSHEj3N+CK2uCTP7IBSGEUig2uJHf7T0WIq
ZxszTtqH659MwoHzs/1aPpbdIBXEDG/o+tiUu8dQIFDHFNABOrW4A1wNUlFShnwd
j47a4CwyHJEZKgY/+DXVxaURzF9Glc6ZXSQZWFeO2TtPj8OP9/rLn6zOw1/4h//B
`protect END_PROTECTED
