`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QO6MV9BRNVfFIVMKHGcZ9gBuvdHcMmA+lgEC4LNKRiFmgfe3xECZkBOvsSS9ZRWN
rh8YHJgfanrwZpsqzf9bN0ujCYE3xfewuKG5rHoQ2wOM5qVhvEJcnMPBV+wb4Qrh
l78Rm/6xB4TLObiGf7EiR1NVZz3xJQ/vpUmJ901slahnO0dWUBJK82dBrOaZ7kLO
sVdVytu8U2xD5zu0PNidZvfUSnh7MIOj/VZKJcQzboczxj2Wikq/flKM99RdBbQn
pMACGrEBvLXZ8lYDoqpZGeP/v1b/mCh2pWVyHIjEOsSQYZX4b9P/HqG6pYHfXUdX
f+xibT5+MqRL18MLYdklAfyKdOg3vxsfRSDVt8ezQUoGQCiZfX4EYqr/0ZwPkdgp
9jgE5h7waMZ4STFvvtQDA2QPdZpkYzC/tgJQ6gB/WSK/ZBpfuJZp6s9u87c2a2lG
VcfJFdGRAbTMuVxRJiedgHm/fhbHctXp1sHBozYCBKYzTSvKkWTq0t7JyjWHde+n
jQ9CijAUJE25PBfMkP1vVABNst+dZcw4D9BlOVLsCvgTMgb1VNEPEHrI6Je0Pyel
DDEuIbZBSX0t0hWbtsIDTja244roCXwzSN3/MtAxK6nzXBCbpwGiSelkW2hBWnXo
3eqDNmTYWMFIqet1TSIBPnEiapUlTXt1nyZ4/GSLFsDiYTnBzO02U4qcWVybfi4L
poiYePvXH8SJ6jAzk82lISKl7ILj176r9dKkIHCxBnEpS9SU8IDS+dsoyvtylxFF
Jnsx347/aRD6LpBVEW1wDg1d/nmMRZypwuEjmNLUdylOL8SxC4ArSpmpUj8LJuYa
SIPxgpcdIgc7mD2PwL1YS96efR+xzNPfX47+mbS4tTIj/5Wjj+LU9NVHJAoftnuX
D2QCtFwc+Ui18s5drHGZfqWbD6eligW5M2y5NjIh5BrPJP5jVliNqU7jljRGw2Vv
3jgsV3Yk+Qroc/Vi7SUUjW41zFBfsTJ8CiipNpPRqAsGRmlSVGp0BwnadG5lpnxd
chbUH3WGAmt5qLaCc+MrcdW6Bb6xE9lMpMFHrfu4AQq1TMP/XLTS0fsAzwsaRKUY
jFEVi8oUTgm5vbrjZzOE5Yc61e270+wnKyZj3HpTOOOIEyqZfVphWJWs+AtKrRbs
DTozdRzCEKEgC8ugGbyqlbTNYrVEy3QofGfDZyfXVlrNh38GTaShv29njrgMlUR5
WZlyVl15vWa5YVxl/l8sX/Rx8J71FN7zznwg/nC7/adVXfokTadMMWblLTvLnn5t
hSvFTmX0SCWjXEFS/GuNx0c1+JNrXmdK4py+9dT4bGdbdgNWv4aVsXOPdlgcVrVf
`protect END_PROTECTED
