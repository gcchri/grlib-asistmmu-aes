`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HejGS52OiOV2PjWyqY9HidlxCHBRKf5hZCyvDBhHutKyN7J6KvQjhavXXqyjs02l
4E08dAzX+siH0JIO3GHuOvasEZ4dKcxm/2ZXLGhvEa2eZVYbXVFOluUpOY2p+If5
qTJsDI01X920rG5WO4rVUB2dmdhcjkC8saMteJAhBThYjIdV+AXhxjjAtDkyddxW
yIauSZp+Nnj33k6Lzpr/7+iuXPYFGo2USZYoq03dpR/uXSlwbRzdmcJR8umQF0ra
3QremQ5i4TRS9dP554hR/9vgFWOCJhJErPYpic/0qyj1l54k/JtsLUKA6JyI2iDv
S7sIl8toCHugZ+9ZVZQL4yQawA50/AFlIB71a1zLWiaLGt6BPsCH2oLhH3sGczwX
uB2GoLROVHTM2Y7A6jTvxHhHN58BhAA8lmIqkrkkIm/gYBPXjoADnHrEGdtlbGut
T4YqWaVwC0RjfsSPJlB0D7vmDrYtfKN6JeX9p/hBAGSwyTT7AHA3tSlEDt8WNO+n
QYkgHXpnCnjDCuPhpe7xYYVZ3q97bjpalRJIEiLX7rU=
`protect END_PROTECTED
