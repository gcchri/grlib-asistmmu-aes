`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aA+pM5DaHTcKRY9t6FhFratSD+5VuOTJC37p4rSpGOq45d4atuY1xMx41HA5JWcg
Aw7BOLCt5b+WRcyCj8wibn0raChwh28fzH9XtNQn2ybW16VoISALLAHo5/DYLP9V
EU71KdJZCKjVLm+XWop7L0SgJ4z3IhEsrd9SK4otiJnQKTbGmqJ54TPX0JpXoEe3
rcTQsw75s4CwNju5nwSm//GvSteUVnQ92XO/D1bj9AfMwGL9PYwFaSpOdThbZjCJ
Iq7wyQ4VBUgDulqbQ57ION2AL3rnCfW/Frg7QGKwajwhr3U760EeKu8jm6xD8RmT
+d4+C5wPHS0Vi393RuA+B12cHYzBtoy2VVLmUW/FCRWEalquK8GqA5jlP2ZdMsHY
Fytzb5ae4Y7fILMkwuz+B2Pp63eSH3XxWy0hf/pQUgqvMQChgS4y8tZ2p0ysPR0n
IkIUDpoGBPbV8HzXe8ojJBI8G2KANccZklpDqTr+vK7Amb1zMvoxqy+4iqa3ChYS
K55aX2gUEk02hPkAZ/zJrVjhdjPJeVKGizu6b461MorjQw9aW7LfrwaseFPJrflF
EghA/G2nIAkDKw4NiyHK5T5WUe4vn5bo5dgsy5GpxmFn90jg5aDbQ0PmBnSHvb2D
u5bIEPNyBywaPmXsU9PmNZpynY5obZSSy2Mdqlc5plaK3LvnwDfxR1Y5j7bodnzz
NHyODlAh8uooG6qYsmMSMKOeJtBDUcL+Qqu1vTQY9mU+2+IEFMZUk6Ipdtz3Q9+f
bryMjPA+VYwr6WO6uBCyU01ute85/evsO0y5Ag5+Udcg81koRKAMoK2sm+900QHU
1n6/+xm34gvUmgojCTuvK/d7ywY7VIoQNJQ5uAnTH4Pi3xUC1srZAEBMPnm7MDVT
rMnfKTOy65ED3FfwK9vN7Zh6EXv/8yAhg42eIY875ZCSU46Slr4J4C7cBjHK/nSP
cmw0sfg1GEPlFHHUK0VD/5JdhnUzdNZDu084BfIr8fAf0i7fnpxC1VH+WwT3QYb/
9uwNJ+ESr1QTh4oVcYpJl9VxBWy0i0tFz+1opVIz5KvTsKxDcFUAzoyNikEwPAQ9
d+IXvXsRTtS1SlQHg1HJgpgkrB3rCV3Qwb03vgalCO/L6pNlm57JQUQdoHwWFoVx
TIflyV22sZ6nTbPqZueTlfcCbGO0y+aK9laU5BIBZ+S94Y4smNWFHXsMzRMjYS8D
x4XRkzM3VSGqh4CvHOPYv4hQeKCwBdVw3YViEfsSex3CZum5y4YUpOAIs7xzOCam
yx1Jn9Xv3EyIFQhRL1/Eqo5V618zh4KgA5OoYNtvJ4OTkXLNmSYFjQRhRp/7s8DX
tjAOGk1il9hIrRZk18D93pJY5mBDeapwDa6F93OB8XXvD1I2kw4fBiv1CTw9cerW
YDNalPTHi5/etSsdMPIAD6tkjXZK3dAOLIStQPZIrmKtw3nBBoflPdT3BjAFdz9c
XIUmy3DQVvD4Nsoi5t+ZeoWc+CjaTUPYDuVGf56JMnZWjirgLahvNnctZToviSwO
7nugI75+ntc3XSJTrCsYdBYmDwGUZT1o6zzDcusxkRDCA2r4Ysqf/gf1wog6AuKO
/XgtsacZ0t6kyA53/YIa2uS56IGZj9jaOgcyX+5AD4mQ4d3Pw/VRu54bQAoMWdJc
jktYaMAH8B52qvX39F7o1kv3wHZp5JrMQCIQoJzDOUwu4tnXBtZAcUKopa9ooHv8
r5xscAukP/WQfEGkvy361mRD03oPzsNu5MxVHuKufNVZ7ePdfpnP45WK39P/qlzN
P7Q6s8mgT+EjIbRLzFlVCzBNsPyE1Z1I8HxZwXVMjFVIZ31+bg/TA4oMTmR9N1EB
alrhuE/CTQn16PVBqWKyoL9d/ejjR+ZNn6u1ml6q7X5dnny8c0mMsswXqCJz3wyn
SggkoGritJLn7C/EVsuY1yTyEnO1WHlumf7bixStLXxN8hUIlgSeLlpGCmHSbsVD
+b2ivPAlCzQILe9ByhE3dfwYUl1oXKq79R423QnSd737lOfO2DnPfYFygfCYhFqQ
J9GYAHyRNB395Qn8Wm5ZcD1n+Nc0ZDxceKlkxNx14X+Sjh0f/L4OBDFHA1whfojV
JzlrtHV9rG6wHrHtycmYcCrPdGH1vwQ7T92k3P6RtTe0Yo0tQx1B/+wOLkAp4hRq
3KFP+U1tD3Q8I0JJNnhPtzGX77SanReKtDV9dSWo90Fjm1cMn/URx+wjzNnWG6Ai
s+mQBY38C2GmxaFNcc2g2aFtpR/uLh1QfHuRFrCed3S3BWUIyiuquoS7mv9PiVfk
aB5ySkKxMy5dikTZlO6hXl9rup34fZY3Q5u3Qni3fphhnYx6y6JPIfrkOqHdZRba
8Q+Emu7+r8VSq5GPvVC4DqgkoiEidU8tDF/KqPgojaJNFRygpkklDDxEQsEaI6tg
Og8oxsQXgreYkej/HPuCd9I5xPzXn0sIS2mEprmW85DrJOvg6bM2kMtb3Jj2gUq0
qzgzfslIfoJJGImCametI0O3Lv0xpT16eVDLNHRRPsJqgfhCd1vaBTXaRL1CjzTm
yFZjZcUaUM6qjrV9iWStBvU9NhUnYY0I4iKUf1WhfryXf9We0vZVkkEQC46YHkB2
fFho2th0mYtOoszq3XLX6DEVKqYpDHLPCPqOczArH+k1CFkjYl3F3dZQUaI71CTH
BtwnYiyxhgGSstu960fuCzX9Nm8kEw1Qony66q9QKDIFsGwcpSwponCMRHu8LF1Y
Cc/vmLKeybTt+cdBSU0r4yrS6L16l4EdaJtiOms+GTEVMvEcKYwcLM0FmnAviDAP
+jVW3rJEjtJvSBUwNOHDUj7EWSep7mXjgcSmBAph3ytZRUl1sytXTyDA0u6TBOE9
tL0KFfIt4JvVk0O6S8CSTLyPCXIe1Vv85Cr4E9Q52xzc+UJwaYalQO0S3uBaDpSY
qS+gMr586VCsviYWfVoAUUd3bs4LclBxp4YSCeXoLnuHML2Dg+zqZGoho9HgySR/
z0xTJt3q1pPFJic1q3XfGlpbYIeKYb6/XR9aqF4WcGBcK7j8LxiSvf8CmC1VCdZi
4b4nVL4Oz+OOwKRnH+aDHvqzNCxbFkDukTeTv+AzYmRcLagRX/QYrI6Y7jfwsNYx
H7wgAGW6M4I6KBGzHUDPNGKKPJDTars1eSqdemaBiieTPUQ6UChBlo4Jd/+aIA+S
L7sdAH9EVB/U0X2nXpPP4/f9fXhVZKlsv781/S8b5DUzMz0C/oeT0pdWUhuz5bxC
0Hl4NxrsqXA3ypjWiat4kvDjYnLjIDYmkp0fJviDPYlKcDsD/NHZcOFGISJrdlYY
cN9FSzBj1WIGF+koZGte2vjcqr3fWyuXRIP8r0OhrK3LcmT83Pd+5cRkkziqN61m
9T5rpJ4CAO9MgXfK+NP8RfJ8aDg6UYCyZtbN9HpJ3zMvV3PnDeFQm1KCHcUqHij/
U7fBHv5VfEEyUWDBl2PWehIQn5WJ31OurcrEkkcPrbIg+pozl0Z1t++jVeJsQTNY
50+WSdidvIZ3RKEg/PVGLQ69ix1wzocB51/QJpdC/ZIrdviAP2PRAgnexj9SI7Jj
q9cvvYX77xSWX+U442oxN8gTbweWLrmrjX6q0ocP2NZEy9EtFT9Yrf933X5RvSbN
WCFATVQoyRLWJJzsleMa/vm0HRewX7qUnMo+9pQ2/qDaoLTjn74ombjq91SXebK2
JAGMPz7XXb9N0Hsff4IxAMFAviWJ7rQFV2RYahiTmNS2iHAvgklqDp0rOSbe2uVC
kEWaJRcM3MGvPwOsIG+7Dzt1tNWBqAqFF3FfB1eYCxurPO546ygM1O+t09U535ya
ZvfUXmXZmsrFFx3y4EMGs5Tx/E707a6OfthJ5qM5G/4MbrtKm/xLR6YarEu+IWds
tXpOrHUs9/hJEUsg2XZyx6cDlD674Eu6yVLT/OSPt/vJ4lvmwTPJywueF0pJ2yrk
AJMsMLP7k7ba2OMm0KpHgxYiteAgDyT/d2Aw9vohV2eV2+IPZQ+OUWuus3n31104
rXz0t+txf7k/Caj6D+1HeVLD7/v/Th51VhJ75ABlaZ6HqcGDEAqmsWdn0pfzck87
iSt5w2q3KhBMN9Jkky5sPEMFmR1ePaD4LLcPZ1kqy3ZqVI+SaqS8KUWRlK8Ug5tc
JhdojvBEeuZylIUmtjMwF9hMyHRNtNxMq3OmN8wKXDN0dqTF6OpnC8O+rLVfiGfB
MyGg83TfbE36txxNUxRUEoEct6lk/Eoe1h6XcOs0vt44gjWOhX9aoZPDvEwF5chd
YBJKGrwgFJds4P3j9K1us6KZ0klHboeOpxjBIz5J3Yc6/gFvlojrx5yWtWDuozKC
Wdn6OznZNqY1Fdn0xKz6EL2VziOl6s9z9/yP6DJYUsD5cJO6Kvg43YGas3Fpvd/R
Jj1MsCq8iC4KiXtAofHhcyDXg1y6mh2XMJtVmZoU0KW4UGQ2G0ptPCMbIXA5hHHV
CjxtfxPBX6YN1pmjfA6bSab4NueolI1bXiNKlyvh7cWcEEBrSgbBOgOwxz2rfCXn
y7zUp8ZLgh0CREBAFyONznFNWGMyfxKAETgU3FgzQyLkIInnFKy/hYRCykHRz2Pb
DZJkgYLjwU2nV+Kcg1qMb76GqlWIsCObIvQ8rFp74i+pDkMQfI8Pl6DCAYxIIBkb
NU4w9/iqiS1amWsAK+b7nmcGIUI9mZhMDR0+jzFK8oaNwpC0xlLdnis1yRrPq4DS
s2j81zFhLT2oJMe/7BlvsP87TuoDBMMiOGD8JYtXO1vAzMMP+TcNbmIc3xPpP0A/
SY24nXcyTT2KYqKI25D5dOkyk4sxHs6pOQD+G24KpCapFG7LpShIJBsNDcqNpptA
2GZ2SadDU83rFvugEz7dQOFelq/4h+5ZZ0TUfWR4X+St++bpzHfvAgIMzALsBhb5
jjpckjKRz2YJMsbJHmuIDb3FxpA8zBpEA27kU6Sz4cO3BAsjth/w6hHPfjj2jCi8
sl5vrcH4z33uVvuAU+AGcEeU6xpEaKxRj88eD0R9dczCowgHwb23ESLBij7dOXxJ
e9Vdju329iRCHvfztMJ8cS4yCHaCR1q2GVw4CVlcz5HfnIMj1RI9/QkJWZZ7rCxZ
rWoa4zW0wYBCHx4ODRa99cKWgrIAkjI0CsrraQJ04cCAxPOtVKfx7AJkRp5AOOuJ
yBdteAkl44AifZD5m1FFWOSWcuT3TibEpAHxmY1A7zpFMnSMe0vbAjOSDF2ReJ53
DZSi8dL8X6HF+VM3gTVu0YthPwMUtXjRvs4nBrICuWadWMoUZtTXCRmEoC6VrNvx
Nh7TPxLxsOlqUooSk2QJSmH4OlFgPtME++F1TtNaGUg0O8RmR4/hIegHL72yr/CY
kGATa2FzKh7IGvK5KeGfi1Mt9Lx1/Jv6f8C8iiKPkZCtMF0DQ1oVoQya1oz9ea0v
bGh6FyJxk5Uvu/o0iuHdxnNRc2F4CqF+KkxYVslMJoIthCSjSsIYnbXvgxQgtBrk
pwasRENVlPYCt0mjWViSHiTXp2bLlfcvYjnyWuMiu3L12xK86kTSFKeH5EYUCxuU
RobxyyE7PkTE3muTHoRRoneDyzDsI93UGWpmvYLpW1Kjl1tbtQ27bb7tIQoQ6ipb
90RvaVugFhM5/oBlNsWgzhI1IY/6IDRfXvxyOjp5vMDVOnQSpuMs1v/yJ75/ElPC
kQJjs+orNNJL48tSNPwlWj2oLn8Xtjz2Fw874KCMb6pQckRcS+Az4+Nzt5ijMel3
mGHesNLJzcDFVHP6tpZutzQwbVyjwA9P9GKpDa6Z/ni5qd4/JCehlAQ0Sa8kXmkV
U0/TCEh+XIyG3nJr+FJ7XY6rtar4Wj6Et/EOq9MPKKut+JVG5nPUnTZnUKBYQxDJ
PT8WSarTTFUfGQnCwvqHzdgGgVA2cPCAITnupBJtPZeLKdv30q4EmNJxTk4CLBMO
7c5jdzw25IlimlL4jMHIw95SDB4IR36JCc9aLn5F84Se0i8VJEho5kJlQVfaIkBA
H2oq5Ro7bpdkwj75jjzhKeHEEQuas/whFDTGOKCyutg8nAxBbIGyCEa95EK7QdSN
41u7NuM5yt7SneZdvGb5hiaIHu2bwtSN8T8HWUG1s1T7CRfLT7UpNYva+RMcsy8a
pyJaWeCdzffXfuRadI1vZiqwusQJAgYhnLfA4Y2KH+Ycxu25gXeHapbXOpwsZZ0T
d5XBuJlfdFJqCtLyN+TFgH3iYrocHBLLFjIYEqUQ5xYhuV57bM4tDuK+SRQMymcf
VOhlLFwCZtoJBC0Cs62oWg/sL5I0RvcBHiYZDOujUaLQhR5tke/Yg4z4qDoDt5ss
YUZ9GguGyoW3CqML7+mcf4GpLkcCZ12c51Mga/YWOquTLCkiR8EXQeUqDPNzm/Y5
kPDkRO3cTZv1hZc6dxu/TzifLINEZ3BYm44aRlzDNFOSc80AyjOhwJOrGTXvWzPV
nA4jjBTtimc90rGHPI+kahSZeBwlwSOVNiQtFKA3FnuzOh5tTJZvBcKXR+/tWjpE
P/McsAQJh+Xik5o7Z8rzKtsMR6zEXjUBLe6pEcbIVu62oQW4k4jB5YXlB5A0qYxF
CFbzIAMTZC4hJQ2tOJmpoicmUz88u1lqTXK7uBPtN2geQeN/wnzumbE9U9041qPl
G/sqB5frRDlAJgrQF0bpZNgrSrjoHCBQPSxZOLY3VKBR8v/TMYs01kxj3hJwWcJD
aNV75IE1+wde6827ptBVe7W9hYQgYSXrwYhK7D/iW+ngkJJgIzJJjdYzG8AQpmKh
GkFhgMHgWjnLPdspWH4olPxtz/3T5MIIUORQK121mvW+ZlmTCqr2huA+tdlIDPRa
SeEdfXQoW4JhGhM2ftxkTlOrBtuCLV09a/1te1r6ZmQXVjyVF8PEwIgPyjiYegoy
K3LXLSqFVq0Fxw0tQlFwMGJo81pUrvHPceeP7Aa8a2aOWR7o4A0+rmad+AnSgble
2KGVpA9non3GsnZR7dNLCIuIytKlmZfr/nVZXrldLr5K4OzTuzxsn31EMH59CKMv
Mo+ez/XI8/BCPulqulPHLVDAqRrMCx3+DqpzOYZa7FEzIfn38ESkvy1leonRMwCz
V5ienmbfeCxDkaSGSm0OvNIzGSJJSb5wHJWFJtEBOvP/bVe6+b3Y6OHVVflnwGcw
iBOTU7IdZFtIzXa5XPlPybpXz/6puUpG6MCm0RoEq1Goqmo7zDT0d9/ORrAt+xKF
aT7eo/W2wFZUoV8ItgxsUqfH0j1xzA0hK/IaXQhmpqoT1SIZWMcUXlH1MInHfBqo
8SuXEu3i0N6JhPfb4QKJb4voGA3FyGY5m8YEy/wmW/UdvaOQcGQ/BQwLLuQT3Hew
IT7+RXQQPljgXosU6ilRL0G/GvDOIZkjxyMEGo86p+OEfVvxTXNUdeGRDoB6lsc2
/uWWrKWluctz6IRm6/xEYmNTynQdNXI8TQIp8LBlR67eRgZNsbObP3JJ6m+haqOl
qT3ZunOg/htfupsvodmVKxyN7DmzPi8U+OEqVvhSlpPI65tFQzTO8xej4CaiQpc4
hTFFNzdxzyXY0RWvPtlGWNwLJ9p3G1mgEiqkdOoLT6GepYQ0tsI3njHE8WMF/Zc7
fWMGMIBHoCy5QqtyKxoDukPxjo+Fxj0H3Av1jF8ySHLaHh5+1kMCy8Bb13lUmv7E
rWZtcDso1QeGcyhTVhdmpH1Y8e3riArM0U934b5XAVm5RhpZEqKZqNIrNsSAKePG
URw6K2FweTeGaG8QnQDuIaXqGIjoQzjbgnuica9OGEUGRfQXfzd3nSVHYdy8bc/D
NcGR7k5AYrTPAQ8KYsAIV5UEVjty6IJ29Ms6l4CLnCdFBTcpG921qttXPUdIbaJ8
BtSf+DPrXr9x+X83IjLpEARjXQvpz4W9U0+pyyhoDdMLXv6Dlq6IjHWluDbj5I3F
UOA2IJfgvwS0zuK91uOdup5E9WyT2TGalA9XdGDPjQkOijuQBezV6EqguIy1vOVv
kmP+aaLtsxGSiGU9gf5JgwM4r5hNLxX5UgLDAVk1jT91P4BGgCF0Xh5vReXhWS+G
00Zf0kCATxJMAu3uzi6g3c6J1ldIEYoAt8VriQeH13ooTHuP6GOAr8MLKz4j6R0k
re9foq1lU19w33AiiS4af9Rk9Ax3JlzTNY+TRYWGGxXFNT3QHP0BsmBJw/5TNiVY
Fqc2fYrGBq/PuYkmos4KNhlCGiuenx59CYJaNde5TE9ls+ViphHquWgbxfhAY0U0
ZKrV5jt9Gjlw5fndW658zBzkbgW8LI07r4Fn2wrIuVpDSBdWosxtEwMXrFaw4leS
Jk1YZlxbisuJgzAuXFjtj/mMBKJ5UGtNzUHu6aEMIiFf9OkiLarBkYqQLeievvNC
iC+c2kZneHmGjK8ci8uZhMrYLLd/r9nl3v9C/f6JLvcjtVhYztL4RQMJty4jNeqD
R/Ud4ul+w55U/SPfTYpZUsjvPzsp8gvWbRdW1q1ULH5fvTPhbT0lGEnA5QCoBnaB
p7LRL8poflVUfA3hkNPAnDVXrEIMQ9VFLi+4CNSnFRlMqPSeUFqGUcAISS2roTW0
mgeaHxG0QnHqYZqIOPNpqVnd+o9Il5seAkmq6U3zQT25nKDi2RBY67HVHB4O90hx
/ZBKhW4mukDcPvEk7MQyVzSLKX0EyiiPzRyRFMddKXWOM8n/1XZZrnzEDMr/itKL
Wuy+MK2Xnnb0pBIo1ha7sdmY20JCzkNWsgRj9yzxpqytsxCVpqQnZ/tQN4Hfhjob
ZE52dqUCLEL9dhziW5fcsmFZaVCcT0mnhLBGgLwgqdnbIjHHPAfbgkdy5BHKE9x3
LQgv0YPIyDBOlJHtCn7nttB3l8Pyb8bJQQVTLvjVrsC6gq2mdm2sglBBKXndI9BL
FQIvnC3H06uOdrGs59o1W5AuFmGPOn3n42gD1RWChJyafx4SqnO/Ycc7LstKoQFS
Or0kFtKeFeVZpS9vwzyuOfRBqKulNCXHd+AXQbrJeOaNeIE4LuUfb4aBL+KToXEp
4Oj0ml5257fqffzfh7diLVK5jpaIS5dKjkxOEIdN1jxG7F1NBEyTvzg5N594aIgA
6277vThCQ57D2UpYsSz3DXVMV8hFbT8C3PLDqi33qIOMby67nX5WYjgdmbWksckC
GxlIpiLXXIJgx/mvICnzMfEGHyfQ9+DUsCVAlh85VEflUk+Gupaz/yV3cZzmRlEH
a68z6aH6zTWQ1gg16Nm12zSn6rJLJbf1BAyW9wtfak5eJWlIZHyfzub38WFi+Lez
35UJu3K/gEJmFNdV5T1rQVJ0Koz+CwvGiLE7Xd5tV9jUKUzytB6mKFyn5JiQYPxE
6jXMEjmdcm1i1v/QmNbAMXPotaVRDTSL1geZNeiHKodRrE+hhYFbzBSwJiIfqqy0
3jLm6e9MyeJ+8g8E0bLVczEieOQuo2NTPSYdTYzz2HljTWTYvSIWQ5uyQcSEfeT6
fXoqo+2RGZMiZfRJsAPJdhZV6Lo7ZusjpID/wz0UwAEO8x9RKESYE7Eisq1HID+n
v2d0pb46K/cY9dtPFJ/gq6qOa9Se0LIMnPGHhTexGuaf+Har8lggG2s2gcO/k/OK
VgiGP7x18L8vNYd3BfInA0dR36qVJxim1R+RQvMVxg0n9RJNcPbjewwk+Ky3IcUG
fNQ68JvWXaPSI0R3iYKOuATzkQ8RHkYCVO0/lTTYCS8xSSulKU5Kx8iShK5JWWeG
pCTRRKJICukmi2E/DMLGeuvSYzV3hzOAGQwyFT1r4Cp1rKqM2GFHUbNSiVhVz15b
QhjaDbA4wYa61hL6Vzwjefw3tFlKegnELcMd5b09GIYrNsR7tJJ6Zr9d6fw4FOi3
UmwTkD1l8N5gLRyLHxCbuPCeiaRuMArjJX2W4y3IQSpp2hu2nzXupU6mGogRlJpv
MwEJ9XAIOXf0OsmLhmXoNHHt4TumEYzXMpMU3ZYz+gTIK0Ydu2Pf8bPjtO0YxTzh
hcoFodom5gc5d3ctL8LA7ITzv7PJ4S7OTTlWpx2IGEmibKN+ttwabd1636WRBAPq
C42yMcNsgTDSkyyBxoA1SlhgmqlBygm6tDMWA2+goiGbm5LYPjVnYJJ8FOlcDA76
OeiqsH3cBp5WfYy3WP+10DHLh3i/2bQ0Q3j1R+FpjO7kQLE/Wd+pWZ49Hgz1wXit
TyyBzQgJMIYz9bQ1sJuD11Kt3IDsbSsFdDGhDnYonJhA5cgGDEdzi9Ofa8CfIRD6
1Hs4JNxcZekjtU8cncM0SSBe8xaYhY99uIsPlpPb1klrVLVIYcxWqw0t/6vaPQsh
O8GJaN6UrzqFraEV4VArgMhwYAndrMdW/9vNGu36ej6B3Ch/6J5zycUuJ+3Gjneg
Hxu6Zt8k8xE/0Y4mNKkvHVwLnlVmJjJ4KqPMismM6G5wYZ3TPCco631932U0yyj2
oHcDwtZWOJ3Di1BuQ/0wvRmnWJeSafdBx6LvU6r4hp76mNXU0mSP3reZNbgi7OBU
YyFwsRZIB33FJUzLhqtwT8/nTLtVMKdVGM6W2K/l2LwQToAs27egUdo0Lk6+CE0Z
R6VZcQzOlibRykcovEJ1FlKOE6EEhu+lIl6h0zqE/fmKqavyUB0+XnSLmT/xgdGe
YeA2DF2tyGOdaKzhiP11BvY8lQpQKYNB7ExsSKrhnLowkdaBZG7vdxSSktyd0BSQ
DoJEH8gVGjE5CfnqhJZ3ikMYvtUWjk+X8T0d5kJwhuOlEn81EoTZ2ErPSRafeoeq
++khW4V2zD1+m5re5EnocjQD5d9HxaD85bt9Gkpoj9FXW4jfiPVoyYGE8KKqK/z4
nHry731oIH+MyfNMuvysx0EHX3CXy3JiVnhQW5vwr0AuBFbjqhIkCdXomEjWy6WG
uA6uNCFQ56vD5A0UUBVGFng+LApF70gx60ueS5aL0/t+ZTiauW1lHYLwKaX1HACb
yGmbT68WqsOs0B00H8bu3v7JrR5JcYXoLy1qMIIHGO2ZT1qJP1N4/13ZkPsCh3Iq
qhTynMeE2yqSMfsKy/o5ucp68HdX30nO/xHUL4GmsKWQNfmnrZTtcQPTTP0JU3c8
Ct5WkPSPASGtBLaIHv83eRI5QEtGhVpdaHDCVnc7EkUx6EJ017kOGECGaArAGuBB
xCBvquKUl0CZVZpLCqYAoz8ifYBN6sUz8BzYN/1IaaJON0F+6ThJS+4ExRrrG1oi
W2iogSP5hp734bKi6k6J7J43wXzVbUYcFm12JHm51qFh/2/bTIJbr5yRgCttRO4R
/hD0EFiQMVKSDsD+I/k/d5Hqho6DSn2r4FepvO8+e47YP+Ko57flS1XNrd0oHUc7
cko/OvIYIRvUOxe6dn3Npgz6c2YkXElhXK8NM/PJBBxuc1TkEafaaWZqGWi04ZH0
jfwev/aFyT7vwr+5kRKDkZbUdkrW/fQx1FyVYEvknctb72X7vwZkSPXb2hIizDDe
DmJwh6imqQsdfH1UCO5EuBbHjqIVGXikG0bqd2ZKuw1f6PrYGVy04pXyNNTwdTdU
4REvmRDeeKaOAaR9e7YymUhVLcloIKfbBm1nMk5cdg3NA6WlKxrSMUZVPP4tYVT6
9Q6umV94ssDSpUJQOnxujug3CdjI/RY1kJi5ymPC15TVBZoT04lSTlMbvMF2dUAc
M6iZXbIfmVtSluieQ3EV4Pw6Eozbl9I09maybnKXf0KRXIXvKoJI4Ur3PB3Obvbv
S2iOJwigOuk5XRHp419pJUQWWKliPeTYKtJ1uibKmT1vA0FvxbzVb4eIs5LrBaO3
6XyAKVWMYZeYE+AWOz72+SNpd66FlgZALQkgKSj3QxUspQ7I3ESQbqZRKg6V8K9M
q2p7xB0CRnDmsajc9zceEKYnrNjYfNy8wETpToG3vRqvwLdIzp4il7FeXnCR1l4L
ORDA6f/yakle4ndaGH7tr5nyksiLKAUyZ35VrdJ3kO6t0O6YKEA9IubiaWI3sUDC
njdB+6eMGmcZBnCQTNcNgqN4yxcAmKUGsIYZH7ExNFT9fPaGS9orUwdk+UPtuWhp
YF0guqdADktnjnq7DplfmqU5l0dvyEEhyr24mAqTf7BTPGhRqB/8mYx/VYIW6deP
Y2yhRO44GhbCB7w64OTAMzNpFpHuZJ7TX34YAMIbqj4ndWd+FKXIwx4oyasZ5gwg
JSaWcsYQOn4yrM8Hn1WUmSn9rzwZhaDCVIJ8j9JawLztx11e+hNDQoY14PFLpEBc
L4x2Xvl3DHcWTQveomG6AftkK/N57C+mXwoxtC/fakfTHQBstrxHAYsaHESUwFw4
5kbRyW3mCBihFtx3UrKh1M7mH2IJ95UFv4HcOLC5oSBg39Srkdw+7fbz0zjQlfyB
vmBKPZUvatWNLXSEI/EmbZ/m4Lldy0dbBSos3ApAfPCwx4jQJcZ6vUykCcPbxeFp
1L1XnjENpnSqMkHEsaK4wUiZa4SpMKZ1tfBlBzj0NQYgl7LagGgrSL5srjcTCldK
7vSoXQvOXGdFJTLjf67OoCHtJwaXxzKYKtGg37/DMuphGGLtiTS5Gp2WkV7kozvQ
SuqsweSG2Tf+wVPQ12dEUTia0G7NPdyLhL9f9gScXwELM0sQ+dGJ8k409jXzDmC1
DX8TqcGd/CqByykSEH+Oj46FmICY3yfSbssCqKqMn1FVzMuzQBrU5L0mfDDNK1w7
Gy0BQOIlqYdk/xlwWn31oYC6GtifOzcKoGqjAv3l2Ku8+NewwHmCt6NNs55W1EA3
DSt5+XT+Wh12yNJEiWE+C9/TjGZQli3YRouJcPQ+bsl2QibN0RAGFtj6vEGr8CK5
Jl3STsFaFnJOg/HMm5cdiPpklPCDaeRoCFyYkZC4qfwJYm+jQSIB+8/JGKONEZPl
q/JACltjgRl48lmmCw93e5XPnHXbeZNA8QDdpCuUO+63RHL/3oTLiGr5rBsLjwAa
/TjJNCZUEE+tSOEuTW8reh4FyFYr7gQpN2hb9nzs2TCvCpHgP86J5PYS0iet/wGg
qhbvF7rIbp4f5SHBsrqD84JoA0NVTqj24wyPcte+92nfPDrhzVND+kNm4aoK20PO
OGLU+SRwc+272tdjDbXOLItcmmeK7g6CMniZepIVzoONk0pXIpStZBmHUbOKTUIO
XEC5nCQlE98h5rgzufbtSVlPR19325Nw0KSlPKHd3pxcluGxUL5uAszwYs4hVk3Y
VSkK8nP94uIBOZT7tyIC0oX7q9rHqHAvVpmypLrPN7NdMMyl35Yk1p6fAEakECJd
C3phKZWqOgGS1+oXSKCrxP0OKYsffn1ip3O8MIMuRMAgXZYGYzJiD7MPgk1AvJzK
Xe7okkXWYnIdTejzW2M5cACp/SYOV1KCOYEwrE2pwturHFysHkrvVNrpc0oxmXrm
h5ufxwcvUVHbUHgOdrbjJjJReXqdbv8OtBBbgYGl8avbnB7tO5h8VQVx3wOCofa7
S/QPWyGijnWbsdSMUvMyxc1LvMrqHFE6ei5rTsAtEOCLJQzI+W5xgV9gdF6sd2dw
K2JygS52ff0PVL3PoZA7D8JTjcFVJD8liJfHBAhPrtVJNvmKxT8Sq/XcoDnIWwX7
k+4WrQ5Lz1k3h4zmx5EpiISMvfDhxkzp5Zixb5A0dSB4UNuBGxtdYppxZCZokXOj
RgkxCjtmdt+SIYs5Jrg4S2yYoRv4pWaU4Z04qwfOWSRc2WAxLKukfj6LHuNG4nPD
MpIIe5SwYirVcSTNBqUktXoCRisFvwXRTBaE1KCK4UyMzV32VxTWGy7vHeV0ZgLF
Wb2R68WaRR+qtRMo2lRw7Ehc/twkTyRcit6CN4ZXJa6rAjku8vCn9Er4KG8RM/Ku
TzL337ncZL+MmODpLzF1FPNkr05RXUHAGLDAJE8YAVnYrp0Y91U+A1CJ5OvlHxhr
1yj2DR4mLqnc+8M5HYXpm6XZLw48wDRBybpRtdg8Bg4HNNXFKTKu2dAwMhXT29EY
0rAXzB67FRd8nvhY2LYobmc/0CVq+xpecHNnEiHfxZRqNzlPp0sZXSzqqDXnnijA
EFCHwXDcVB/Xu9ucCmDwDlIoK7AZgYjQo6ag7IRxeBonbAxmgB/ayycC1FEB6fY6
LQdYMAIVZr/imqbPSvzcG1mdht7ld//i0RVYn3wOog+haBGt//Hg/dtEcrM2YmUv
rGOJo3S83gHSmKP7uibUmsIq2l46L32EL5FyDkzl1XU=
`protect END_PROTECTED
