`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v7SPKSzVlr5Ydr1FukKmmZSaRPmKIK2sDteaMt456gm+HOpJ52BaGnk1F+msQd0o
CT17tOmIctNIhPkojaKomsl1tD5wkVS12Shv2DupIfMkBARQAxzoP79i5dD2rO0W
nKqpn6EZ/7sWMhCH5dgIA82LZfB3+X5TTu/lGA7dy1m4rmik6LpFmJmrnaaqDbtg
q96BcfuxQ8cn1JSO/ULudzWVXNBgbrsc996R3MOPKRHAL+YgMKnb/5SL/JOXYQnW
HYQ5UJmN87vFHFzfKXeAyLe6l10vl6egSzkQJ2rOmWC0y34OT03j0W94EM7zjofd
6L1b/jgy10cL6971W3kZ6MoaNN53HyPGCyLA6QnDdaRlKCOS40E13NqWWsf8XvJm
wnVSnSScMpTxIuhio1Uddnmo+Js+W+uLPSuiTxsdJypigDGp7l2pHsKfAI1cdDP2
6w7qMRsm4D/kDvwiUE20VXE4/uwywE2WWUxFcRPDzCKqHc6r0bcZy9hTvr/YusG2
PV9r0S72jI4YwW8UNo0dqXsz69hdoYPCT8Z/dLZHtSdX8imaWjdnO3Kk4LH/ITj0
7f/HLS+L4uZtsgu7V+80vg==
`protect END_PROTECTED
