`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/8D43dkaoKIeETbyv2mPdjwKHmlsr/e+v3b2fgNovvo+eXdbeF3DiKQk+wHG9FpG
026NIxlP7EYHbGpo1VOT6QLpUInRvRHJs7IyRNorlxEF5pzoihkAaT8kfG6ZaS8u
n5GqWEqOp0zNB7HyEI2PcrpS2j+2oeTHzXmPGTlXPdh4YzDLVd7CCV7qe36k59FP
9K/W+mCNpgzeEe3ZfhmHW/fAuYshEmw80T0Z9mIbiCHGCQ2QDwwegW3DVJZj/EsH
JcY3gv/YA4eb+Pi272pJYJdviEC9Sk2oa+kFkQP2/YU2qnxz1c+GOFimjeNW0wT8
ROQoC17hQOf/luaV9h8QHA==
`protect END_PROTECTED
