`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+cNxFrEP5I7c5PJDHy7KGKv4CSB9Kv1XdCx4qDIK4+mtwhFj912GO1AU1u82Kj4C
UYCslVidp3MEFZ+uvPztZ+QWZ/YTIm0eLHEwlyWBrtj90S+dH8YS4kBW6HMc/xg4
gjo7BmdVQG3PJ/cvXwSr6hChSBmqYKOcS9v7PVLGp5+PpGQ2dGNw1mjJAmF4+8zb
4whT6f3SToAPzNEiIns92Z4yoxJ9fR2y5AkkcJ5BpCjWnaOwtJbIgpPanAXhpic1
05w3E0UohLpoaQwILy3cCe76gzYYRZnF+4ncK542Jtaxgk43qA3ZjkDR8HL4zXyi
v1bFQSZQXIcF8fCR5liRnGcpWh7hjpIxRXOtCFMOyn2Ayr8z1ag+HqWsfYQ8rswP
b6CGiVhe29mgHcLfiF6f0kXUyvxjxjZ6EJH4lpTcZzMfSvULulQgZGuegPMcjQHZ
Ml6BX0vFpgV7BlQ6skJW4K9HpQCnrkUCicBzBc1jo7ptvhdP8Q2z/9U5wy4Z2Mes
cEo7gDwJAQjGa/Ut61s3TysMOnTccEueIuRQ+uGrfVUgv1m+CJ7rle5GFhNRP/1c
++l1Z1+uOLWHLmkkYdXjgArv1WwXHzU/qexb603/xftWNCK5UzBfdCsXXYePYxDm
`protect END_PROTECTED
