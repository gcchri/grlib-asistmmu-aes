`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xtJca5uUZ4t35jfAvpMLPClNoARUQj8RAX6VYHASQ9EwskRaz5pp7cb4pQI7H3zd
J9NWK5wJIcu+ZxWVrWg1o3PdVbaefGWStpspC+EZPV9mxbi5k3JOW6//ty7nZWmp
7tepuLnah20fa6vaW2At3R/iw7jFnU3BUUrcEgEYJ7gJySSZF8IejPXZQo+Ew4sO
DRNBrXSPrxxosxb1LKDjdIDIfsLaPw8By8xGWfmAq9PfbdHNVxFmAZApIPkHnC66
9MjiCCZbVx7xElgsGqKAt5ta/BPT/mNZJLOHqAaR2NL43quDzvXgV1AbLzrDEXYi
Sy9v/vY0DgY2pp9i9gD3Zw5oOGnWdFd4oNX+g88Kl14H6TXf75UMsHBCi7t7Q6lz
GwELflNMZRT/7cHDIZNTFw==
`protect END_PROTECTED
