`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XBDegAtY1K/74gPsDEcI8gEtsnVIh/q7jR7V9duBThZk45f3eX8tT72dtMh4oeOq
vj02yBEkmFmGkSJx+AxyInmyr53Aj1qCQIJUiNsyd5XByDENPGH/KIItEvknMB+v
W1T43MeRpo3q5hqe3VLJeELh3OTy1a1rZX8YufCpbYdsw3BRRjdUEU+d+RtK8Bdh
hjoWjzzAj/UItnUcWCAS9Ylzv4em53gLA/ZsN29ddxEmmn9q0YDAQveT4Th4dlfi
QGEUu3mmbqAlP/8VkvMB162UjkWG3Tab5biHyuvmA2s2jK3lU1nS+LoBnfKWWyyB
v/rEuAk7X1tpmZOh/rroa9iTbxY/hdiXq1o4qgnsNJD+qCoWmlmcD+BPJbI3SuuQ
7BspNuqVngf/REqvh6MrlCRO+9QJJubCw4+L4Wg51jk4oyCSgJ4sjJEWgNra2eIQ
sWtr6yN8ZkpMG/srrYZ2GXM0mJI2fBKSPb9jNDOEA7ULpcEx5Lj6AH35mgcm8S8k
+80GoWwxcppWQ6GfyfJ0KISQy2ERzIYoZmn2eCencK3wRung6XClNAC2dN7FYn9D
SXlUQ/B0NUNI1tcVuPJOiSK0TvPhxULWYTGYSAZqrB3LffTtWJ8gZRq+kHfsECrr
t3IAt+GR8pshg2cTX1PP6uhry4etAQfPK83Ke/f4U13/WmNYgf4iQfU4CKrsDKgX
S9rfA2IPeKWurennwg9HzgiG+22AlfEx76OQAsK/EsROqd+i29AQWnV52jwnuxDd
IO7kVXJv7m8u6sCzHOvQuCIJu+21w7fO1r4PZHzZ7curDrwAL8jjPbS+AfpO96UQ
Fju5x49pbE0MsK+klupbwHi30L/bSvT0yqhNrmWAzZNaGuCtBCvzxy0BOx2tjRCb
24ANzARg2tkpJv4fHGIAYiKM5tGf/+o3jwQQXoLQGIzL948xl5JQb/IRzKsfrSSI
RlIOk/BWfpiIgfDUbTcCu6PwYpEp5xaW77oKwJl0IipTwkL9PLlLPtvW9JdnMSnA
EDSC6W0OwDIrwoXPg8wcMfwCc0FaqGGghIHhtY0MGK26whtYu6y6tad2TWkbua/m
+fJ26SZsJxQBOGgJ7DuZsMpuR09Ojq4DGHdbUghiXbEswx9oy7KQC6ZtKNZhN/8K
Y2mWMDl5IsHtAqqZwU9z5QxHCfOOczwza029TU2Nkqe4MQecbNxGuKK79L6D1BWh
204ZpDFIcxSSBzL1uRI+O4EBwh5xsF0Ik2+0QEI85U+/YE/gp+M8kkoq0PTTqVjU
+Cap9ZhiJud63Lc9tcY0Jrb4GOXPj4dH2JvauT8sRTHdUrLsh9OMA1D1w7jd9FQ+
ZpLy4EiJJXDmAdqhbaKcTRSaE1Ahmab32xqw6Bi98xFtVIhG7+kGKlNjpAgI5OdV
beMyudGNj12KOWpBpGOwjJmYteI5Fq4BFnZ6HM1j8vbr2Ar59UoTGEFRWlCSd4/0
udQXIvyBab04u6s3mSOdK05iNh6S5BVVuvr7CcJOfKsovs20yn14vQw7e+scidS1
sfV7Ku7anYo4kEefn2pbmbyWWd1wSa91S/RGWxOy4bnqz6ioLmkfLcm4GHMcA71B
g/dK8kH7xhYBhfOr0/bkb6F+jo9BOdifbQJpjSfOSuNwy5r0Tom4n47Xoke3qfFp
qI/JMO+nZfOzlXkMHV2rsgV+oieF1dEZoiCAK4XefygdTrEKltYqY3vD7kJrxtRq
OxFza5uYY1wsenbKeY66dzl6vISkkjx9udfWpIeW20RdERNq1PmGiTxsiBd5R7Pg
HrBc210/uhkFJos02P0TMApbvjGkaGSvZjmqPgJ0TM0PsXXQ/XPrxE9H+0ANViuS
3pmd3Rx+hEZ1hqv0+KFydpVenS8C/UuCkOKahHPk2bKRJxy1zHtLZfbP324t3a1N
PgOcC+lqr6AUfjnpkOywIAS/GFCtH/hOD5lc/hOmZVtO+8plK39TdxB6ErTtIcFU
cnbTQvcGwlcet2YOdj+57dXmOas/a8TEiXjrSVaAd8TrSM/SnxJw+YG7qES9SFJj
18VsPdaG7nien+qgI5UP4rphZbq/MGTbQ1OWPzb0rNEIVQkOeRxeDn0ZqNnnGrbV
JTbMWRMHJd55igYTVO3V+5I7G3seKk+B7l0VDWT17ytVwRJFf00GeuQvZxP5BaPu
LxkdiwVG4/n3kROOxK80NfZbcUkh/7I7Dq7/sz6Eqikv9qshAPXwpdvtnGXi545a
BnV+Tx4bgxlq3Pp0I59wUtY/Se9Iun3c8VjsrSGQ23IVuIp9Mb3ttr3BQ3MODPnK
Kz5e2JIp0GjTJMQaBoig0+7/T4HwUCzSswefLDVAbXlZdSHXVvQTcndWlPz5rRsO
ioNBQBsS2nLlC5s1SdC/NmiXo8pCgCqTLAQwL087CTyvgOcw8JOfjwAe6PLYMyA0
YAED5OzOEY6Jrm5i7bc8/E+ox9mGb2KENcLr6ubpWDxhtCfysWjSIkSX4yKV2vkT
izFwbSfaOnQAmBeTZEBahE3B/HIqzajvoFdQk8gFD9R5Oaeo+IqXT5v52MzD4RIU
eDSRgvnG58fBkzJRMxmZ7gsTm8/oT7kVHNGj9WPExl/XgeVUuLz9Q5rTU1JqZ7E2
8mm4WKvwHORbhCQ4IrzV/QC7cV/oxTJzJrQpqdeEvDVh1LzuWhFrlLj14SGUkJNA
xVmtKIxUJGkaoe1lMZpJwPbBVNwIy+z1WcHDuyLSqcBlf6xIbuTfSrqh0lxDwWI9
bj9wvbFtBw68EonUC8IX1yY3uWXQWrYNruusbyugf3/EUPnsEnHTMe9JtDCzcW5H
AnK4QCHUihWqe9xiARYeKjTG4xKeAabTMK8Xtm6Wb3r4WQ6ALfVMjBMj/0Zv820P
e6OwSRQcGee8BVpLliBkC8K3OsloABA2GLlvqXFtJw3tStEVuVBNPHN+Gelm6i2n
G+FY4mQIRz/RXfJV9gdFCq20tqBakbarFlU8ds3W6d8pjzTRsUO97I/MF2nyYwFf
0cWp7DMrixFLAo16YoF7qStDBcVkDZsW6TQAXweApvbAnoByHZXtE0SmDMI9cpFn
6fgpysscEpjStm8HACfx/tj8IRWpCKL6kA2rgDyHQfU/MXkErnrNqKhMpgZJ6EIV
M+BqGY6Wahbr8nlGzPvqWkE3FRxNiV0UZl+muHynMsPdvjuD4l1qpH3egFb5N8DT
9ZV4kURehXRCb689YGCDHiJmLHWTUPRltJcGnd2XpfDpEkDIVVoRsgOHolnzfYLP
uKUHRyTV+9CbpIhvydLmvZwhg773aBr/0R5n1uYP6JICy07Tf8gIaIb9gfB0RC+M
eVum7uEfCsO4w2W4jmukhR6lFXOgK0Xz0ceV2hLqA9o=
`protect END_PROTECTED
