`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hxPKEq3tI6h+gWnE8I616GXCNnP8xXe0H7preqitBrxUvneMyOUadypeSVj9vc2U
bWmva/KUftA8A3lm+2YHj5Zn2pvEmkBcnNAE7mkmMKkyieoUKhVkMvn1YFHdcGli
IDWcXxESB+mUaE68AnmQ0St5+Dajx5EONrTaQ7W+HyJYdhj0YjZ7pgsTWLVRzbcH
10nQeIJcwetlNAji6opp/JL+161yxOXAV7EUuRItqHAs5PHihRT0bMvNrSYnLJY2
at9zvwS0JUaJX2sZy8Y3dw==
`protect END_PROTECTED
