`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lhAWbf/rVqohBy4IsRuh6DBHWI1YR4a0Bh21HBnaGz4VD60rA1JbN04m4VXFgRWV
6MXT4K4CjYYx7ytTgpik6v/ZzEco5dayLFIrEu4ft28IC8iduJ2cAqln2Q5tB9Mp
DByFw847lnNA4pt1R+kEiEuPRKm5bUlv1RdiLuBgx64JpFW5pLNg3qcfALxIDrXI
P8ZLHMgC4Y2wwKhIUUSd0LJ4zWkoYeDY9CqXXa5QSL17zYAy6y5/QiFAEhaJrIBk
1E2xKjXD0Dbe/+bW1k6PPGawEqzGv+krlOFSOWHz95mgjorK6NYGcVsPlNRixzQi
GSGjdxzxrPG4diMfLr0nDBlRv4GJok9wG0i6GGnLLA5XSFVgVC56gfDySZQyUa5g
eKl96cGrA6py1o/pcfPR5WfQenMqJzKASU2LI94rpYEjqftpotrRZVjKxtTnx1iu
lo1IFIdPk6apeFjSHpQSm8Db5+O9DMSll5S29EKXXzeV6rpMslaV3C6SgdCBL4Oc
`protect END_PROTECTED
