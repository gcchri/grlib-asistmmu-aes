`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+GXY18VT9dsStUlzYtAnQBnXOXf1g+YyNCshVBT1qfxyodCtu4yJYp8VO7gM+O+Z
iZbwcLLdPCIfW25hzPtEwiOo/FEXR9j8k7cBDFUjAsbjKmPacZGDcq8buMXKDnaQ
BYOCNp5luCOpeJ0BcqTvy3dc05D98P3/WQ7kSJ8/t1Pv0hhCWbdd2krYvYj43Gg3
tjz6cMrGuRBWSsYMb4Ta+1+0oR4eGGgDIgJgBRqbJ+imVCUiyjJnoIfSQbZyAepp
7RHFHpdD4NAM1pVhIOcNWuTj5wC0H+augye/0C7etmsf1l5vyEp3WF0xYvWMyaCj
LfrlNxUdAju39yIEdZOsdw==
`protect END_PROTECTED
