`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jaL7zlMzkE/1P4ET/6MuYveX47eGttupi8Hr/OaktTHeebns55sO0zyv1hTK862x
BwetuxRWFA9Bo2CVRtLlLDD/zJTgQx6Usbn6tpEgo1VvZQOYOR+IsilleuSY7fQ2
RDQAahO5iXtzmMk4DEbbfC2VWJ81Z+cS6XJRiu8ea2CSAAyzatQt/5vENWyXevYM
PswVMqB94zyqLozoOEDbNQh93mPc2YRCSUs2EScZulNHCBz4fhS2D8mUiqG5G/gI
1Rq78KmiyY5anu3HTkqCrEEes7mIa/APknM3t5BLDA6iWmsvzMwnhtX7BzV2mIhu
iRfR5JRcP/iGC2DvcGW6C5xFiLvnfOv8IYcLC7LXYCNf+gEk8+8URncEuFurZzsY
nMXke/Td9XZaAJWt8dCAh09JyiIlSgCsU+okB/2vZ9Egoh6O93M5zfHb+8w+ezB8
GYXXw1HdDUGxhKRLPVp8e1F+wXujI3E4mhX5LrTgPx1m7UNAfh/+7wv6MlbrBFlE
+WRfUofm75Q7+nj83oTWfbieNgEcz1+tFLBsmK+VLrrGZhf3t14sdQo0ScwQufHB
StHfxbh9L6a+qmeE81bHsl7ZD3KlE6ZnDuGhuUyCTr+keskIKKo2981IfRupy8PC
SMWv2gUKLf19n5xLRyKQMR05E2Il9RNePmiWY8tMvLYq72nII+vpmeIazQ+V965r
/wcGObg9jnsjufVTUBo8gXLJeAPiYegGU473lxtCw7Iw820UzJCzKGdZd0GA5FdQ
6r/CA7AEU0N6dnONpkc1dRrCNbsxatm3gMGXLRujfAIgYr428lERVySKrfVAmz2h
4UXuok5qZBffknyluYZjbE2BH7Vi1nMDza9NHPhfoq2m7fLUvMJaLhVV9VXI7QQP
6NLWxc5D/F0l9LVGOi/FMDN9U3hOjqR+Ue7YZ5SQBMyhEKl5xqFtuQpX1mnfCMki
O3JETp4UCOi5NZFzFWbasP76pHjxwj9LocMRwNmpVmp6S3ClVcdU0Xiq2pEoxEMS
`protect END_PROTECTED
