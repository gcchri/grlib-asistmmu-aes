`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o+sJd82MmqoQ9IuJNcHPSN+87UauCPSmY878Dwxu7Jj81RwASNq1CYtiMmIMHQoM
mHhQmptm4v0nvKVoQ5tWdcX5ACozayyOGqa0GBhAxCcdTndViFRk3XqTW9SakKFg
U1aGdu6YLHZ2wMCUw+eg+uYW1n5It/sjcs6h7sY4eCYNKmeuRa6iEegT/rV8SNi9
cdFP63wXpxR3PiTCkkQBJOrZyqqS8TGfGb17er5bBae9EIJBVHc6Z0aRKoGNBq3n
eMMh/pMRfgF/ArXpVw35RZmf5stkZAom6acbiA7Usrdjq0H9hDrnnLo/xAlRWXUT
M1h3vSdM34qBP85IZVmUF0IAX0gbl3j5bWxPmQfi7TtY3X3GmYczPC4iO5G+825W
9gstRsjjHgJ6M+uq0rqp9zxd8ct02lwc2mf56qaVIKVHB8R8pXiiCVd1lPyBOnj3
g9BFzJn1WJX0Smn4owxCXBbvvYIknuli/xsRjNhdCDCxgAOAMEBdMkVBCXeYHjSa
dfmTI9dSMaAPJ+Ust7fIPec+mejdyqYReKQtMdGsfowZEeqSRVj0xFnOclb5ZxkE
zbxAaEBPrkYeoZMb/M2EJtt9b4xOFosp2Jpe7Db6k2ShD3CoaT/L5spxo1mQ53Jf
AjlrTytb8dxJugII6yhEv/vmCGtAizqsCTNmRE5zEnF41d/IDRTkkrb9Rp2YobRT
nsmv8lbogHdKMSf9Dmy7f0pNaO4VLRQby9FXoYc7UfurFqSBCOWx+muxFxcn76US
QnweB14CaYChLNPlRkb7vdevWJb/SwfuMmRWTK8FWp4HvK+jCQMUoM1GeoNhf6Aa
96SRoIX1kPvDGQt4P6/5wqaoNmP/eglGTtwIj0ft+yga0Ib099SO+aV+tOzzYMWp
6W2aW9qYzuX8pkPPg65A235b26/JcjG8CkqBZcfvCeOvT1I5ESbYQJ0kVHgviTsM
GiwDZXuj+FHo/Fz18pDdvbHK3m9pkKzEwDBlLj1fPp8+2gNxNXxFIOLe2OkTgklf
NXekZEmY1sRM+2dHFoRWhmRFlytVsNYw5szdVrcHjOYxKXIA/nDf3Dk4l+U6Xlu7
oXZofMWUfOfrz/2ygV3pjo7hqgxWTbmQrY1Xzl+sZe77GcKHru64F1ib7JBHFHqc
2t3eoSMYnpUFilVlRQSe4OnRKMcXRPgMgJsCAtFl5oTEIOoiFHsicmxJbYnCtRYW
RUvEX0rHMbWau0CIvEXw9AVn5yIdG5gT5m0uLoJsq7C62dJPyyFZ8XQF7ewQBgYe
ykeDLJ3NroJ1YwlGM4hOV3W0iCbzx7CPiv592vE892U=
`protect END_PROTECTED
