`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
68bSkOqfGCgqiBU4zkJhi3vX80YrpZS3BHjgeaXx+AQblz0hD76tJqbc6xD6j40R
OJIAGm7HFjDI2KMbkKYEtJfOcAoH1h2YmxjPy/Kw6I5DSCvzapR76V6ecFysdZoV
WYj1TNNqc0IWXG4QbA7HJKk43jnHpu6TMlCVJBqGM+JlkQuJkaAZS/jQze7BxSFR
F5defNaEu2QJ8A6dw1vQj8Xy9exYyDXJloZet/MiZX3uSsen3V6/rRJehXFEYO0l
f3Ebk/XcJqPVY7fdQ6YvbVviFMIV+VVOQLkLvbdTuWzBUmLxWV9Y0M1jmuk1cF/a
sGKLwEHtKkAC1ZIcxBDQe/81k0G3lU1gtQqWMUOY6rhGQ7xjpZOjyqut+oaR+8jW
sRUT3TdCc69yCNmzfK7A34uumfjeLEnIJU4yqem+nwQdqJHbQFBi959WFVCmUpZo
JT1FTotOoXY/1k8Tovc1oNMGIOqBfEFSnO57NkPxpcpKCXCRhY2hD8Klx64lc4qz
9rMZo+8W4ZZGG4ukWiXlc393JbCXudNiz9jFKWbVXfdftqpIbQyjAxm1N+fHsNyk
J7+uN0j2A6DL07OZqtesDvex0UMZjc5I48yDaDIJ3o4=
`protect END_PROTECTED
