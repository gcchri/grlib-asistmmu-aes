`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jU4CTy/zWTDR6eSTI95b4vc8UzhOyCXY/iYsjD2SZok7z87zYm/BZ8OSxTAp4xKp
pI54xUYg4lSNhX1e1aYfD0Whew54b/UqWiNJsHPqqeeIZJRM7Fhgfqye+LZyzEE4
zvgz7dW8mRUPUpq9VF+bRa8pC16AkrkGnvSSWT1InAQ/yHElbbJ9Kt+FCZvk/kWE
ZwfqCNlIxzJbA5xnwgb2S8T49DwcBTVlQkRTYZpDjGIwRq+MehD7PWRxETbBUlCm
UrVSyZhAwSyjd5OdyxPONba1sVAvjYn85ptyfDVEgdK45inZ/XrH+8mzni7J4etA
AzA6hiv3lWp+Pg3PQpAVKg==
`protect END_PROTECTED
