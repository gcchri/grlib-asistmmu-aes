`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vsFzD6fFX6DY/aEdCEGkyFhCX/T9aWKAVTrbtro9a4I/hE4h8l1ZQMt5k0lpXXxV
9m0X+pFwMWU2BGuw3EGHHgNsFqXJh35dS9+AZ5lvpZeQpinshxId+1SfYHS29Ly9
9q7Cdhz3HaaDnqwMuOjYGepse7WmQ+SbiLYXFJes+BSCUsdIX83UkiF99TW83bVV
WCyLQnvsSeGre1HG2cCWmyt8ZfumifADFDwOAdLjWflYR5AOcifd/Eww3EV9hf5q
UL5GLrGYOlQzBhKavwgfVp2P0YQZT+QC07fGpqsTA9trWaSrAfvtzerVNFDIXy/V
K1fkpHmenng171iNlBzDKuwVYQNcyQV+CQDpA3dkHtZGBWCDll2yWOX8lyzNJiE2
bK973ltL/9QnreIPTLxDlAsCVXK9IclNIYqu0c0UGynFJ5IBi+B3dPUJ0wJqRBqk
7UKNgZglKL/aCPmJ9ONKBYikDjj3XCxqFMcdHO1inYuTWAbTLElpVyf90CQ/9OtV
k0Tc3A3C05C39NiAnpUj5ThIp+6QyDa7oeAQXlUBym+eRJnvgcstN0wcgTR2cuEz
k/KTSzyJ2/s3x25HVBoYhwoz85NuRXDXVF/MJxN1pQYPBpctGxWxyIhEr7WU2Nce
PNLktzpWIEgNxwpS6dM8eJGaGuqQohh7t4hHEpkJpyjkaAj0dhZnfm3wttyuiFGj
KPS1VE8Du+UPUrAZ3X1qr3D6Ng3wopl9bDaCz1V5ctiHnCn0wYRE1SJ3aP84DWUC
ch9AwRVJgLwmP/+IRH6fUrHgfb5MmyuxBCJ1SgTp7ePORoX1PQOpDksFbqAPRsZt
T3N9f3GVlHikkZrLHcCDcqB0MQee+P6jVvkCsiz4pTktYCXLZ00XTxb/igCYmsOT
viDkLCGjtGE4rEouuLVG339n+qyZpvNS3nkfgJTjrRLv1/FwaigTldrFhHX9OHm7
1UUQdMEkX8PF5UpR3hjlDhvctxC948UbQU/h15fDw870GDnqVTB9xMmeEBs7sx92
D+OsPQAgnU1RBV2i9bKVzM1Rvbs3K+lY0+NExYfcS/BuZpKAVjFWkXZlCEY4oq/n
lWlxhgYmlcHJ9TcVPH96o4l7EzdTaOHbgf5nZO2TF9SeK29gW7IMNOjq6AE5nn/I
3nuFx6M/tI/LHFcWTs8J37r8glu5gtDyAGhqkI21KyYmFwZ8omV3Z5mQwjs+CUNk
AIcv+Rv8uB7yqN2CnrIFw81eRzkmo7V4XnbWX/wU9js=
`protect END_PROTECTED
