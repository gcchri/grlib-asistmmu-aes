`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vdH8iWsrYdby3fUMA3vzv+jjt2ZvAJNKIF8DoPZmg8JlpdQvVw+A/GHYSqQTAPu1
4ESmFZYll1R4y59D626tXSMBvTP0pPhDq91AYkUIoCllPdU6TJO2YZMbgZ9kjlBU
O4AXxysuwAwfanzbDBwqB8JezdFbRpuo9ocY3OHL+D7TumT1hlGZ5QhwTLZgmZrL
LanQZhVkNQNYw/o0/QIDcAESSTUdzLmT8he6TzOynjm3wDMjKsA0gvtsGUZGUOyY
Ky7yUBpRkQQ+nY8d0jyj4WQiE5UR6nBQwDs/pOpwG+0+by+qcuS5o4XJHHmKoCgl
59J//rvg9aoEdc+BfU5pkUSb7YYfGtzx4VrlsJburlUk/4Tmxj0eBcGgs+ixTwn4
3NrwrAb+W4rFMWjxxKSUeh/WiuYkUj7BtI4nAwZVvkbBf/maR2wrRtTS6p7qI27V
J9fVQpEjJVMoZKDnFrIbaII4cEDfAreBd9tzgT1mp8qE8UxaK689fbPhwN+OD98y
c7psp4rTdsQVnKOlDS3n6jg7cHAUcgSnu/pAm51wtGb6+WVXXnANjWwq1RBRzQPD
zAJMqYOGi/KzfnaiJD7l72qo+qnNVc7ZMY7erFqcc0Vi5Ai57RFUKYYNDtAqex0Q
gUrihvPaoL9TEmHro+B+BMzVWSTvH5PFKznICzfn8jXGVxh9+uFEHNmJL+bNjaNT
YG54VqUq+YojDAm5r1GPoFeRBP9tkAvqzst5muWjYUHBdk8cZsXa6IoxJDtUsMT6
WarbYU3YEgQOWZSm4irJuVo05vkRGKzYaxO1ZzeSNGYpH84p/4hqGBvTdyrODiRO
+/vSeyk/YOLIBpFH4dP9eUdBhaRK6j4RgT6TVNHk90PJNZLXbmbc3ntpBTxXWHXt
ZwXqPX0ErvsN/d3fTCYp7g==
`protect END_PROTECTED
