`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WJx8oBg2g7uW8s8o6npBIfb7bNC/Knkx1eBO6MzT41Ci6CopCgCA+Tb+Bt5Ni/9k
0RC7sdD4sysBZJ2za2JDIgfPVs07guQxsUb9AS4gU9+yXW/zrBs7cgaybXGqdU2j
1hQQpco8e9v/WQmlXFAFtxxGXtQwO4Jc8R/qYkCIyRU0Xq72GAXsSsTjuWTPABLX
C8v6/StbdvGX77Yr4SaqJvwLrI8lycyE/h9+By/aI6fSsTWthLJc4D/pDW6DQ3q9
AexY3UvG+B91RT7WcQaGMMsr8t2G6hCNxyEJR8xldNquvMBH8QMrJIgf9XCBUB/r
DLywsW/ZSl8n1rHJFidzAx9rL7iLt2bB8ajWP2spqHInFLtAN+NFSJv41CdNrm4j
d3U6rthiFbdaoqjbSvp2bJNfxnbJHHfUdPUsg+vEeUpAoJsxQjkd7kcP79bWgBYa
B82tva89mB7RHiDIS7KrAaJQYeDePDeDsHZpfSD85rxxpLyFia1nYsdX+qP0EbM4
nd+roBxXutEe5R5ndcLpmN9LiThYIneXgLZWklA/p2c6QpDUA8nyz3SQxn5BHiC3
A36N7JcgzKaP3KHgtZdqmO32TMxvw6WZc9ISHZ5h5M/YQVFLIsAjHW0mf/PdJwHF
biupNCx7+MfEZPMMsulrcQ==
`protect END_PROTECTED
