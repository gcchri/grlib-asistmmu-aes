`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S6ggTIuzkNdxILlsCM0XM2ISe0W7775dS4vRwxHjqrrkSGcGiVcce0BxGBtxDsPL
SgA9YjIHhg1ZxNxpPjFS1SETtntq3XClFAr0ERIpqFNBhs7F41GZWXSE9koTe6kT
FCzi1TiINbh257/omlrOoNCS+3pHjtvlGqw5zei7iURZ73l57wQR22ztoD5uhJSW
o0TuZxUPRLjzRVDWPDIWxaf9GHLZzGPsO4AKw0qCIJ6fz95562uXn6gDShxctgNk
LF8dco/fKvMJDxAftqZEc7pQG4fO3zMy7GKoKYXli7vbMd8Mangg0NIG/P497dw3
WCkQhtOBmre2JrLuEptqvZtjsJR6gika8YmSvhY2CIYRjHknB3htPetJ0ZOnj28n
6cB+G/8nm1qAEtwS07e1YxtnrSXENHKQDc7ElWbilx9kji6GLsOG5EkMJUHv2+KS
3LVuX1itsgpZTqaKYwqim0Iux1OCzhvrcFcYqr0Id6BsQmdidKh0AgzIBZXd9C3+
ZvV8MBUdTRAyiZ7SEKkhHMVZwar2e0JOz1IiuwuCMK6hWCLKzDzG1McsXlqAr2V6
gzUZA4TEuVHdBMzvmqvgmGVJPSuQ8qyBOe3QbU5PnqnznzscMQY0FvQud62Wy5dN
yVA64ngoJmq5LGRWriynJadZ8PVlxQt3x00E/FgJyyU=
`protect END_PROTECTED
