`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4VxK2Lo7q64SMri/UoDQqs1+P9C7EWrwMkDxlnaWPVET7tiWEZLc+nAoyAsRmxvS
2WjWyOmFSRa3unb9Odt7xcIXb8XzzJ2ikpYKv6o0EhVeA+weMqscJovXHJvML0gA
YCYjJu6r56JXJVIVmYvUYbJm70HagUkEXhgHYpHQaOOHVgvwUXeMXcUMN2SE5P1l
/gKHnlUj4MuWsqW33O+HoOiUsAhdzjEZtAsyAMxMqo3hFetO7JuJFTVVwDvifDmQ
fUxMYUWMsHPKyB8WK0kU9b2igDNgW7x9Gmu72I5OL9OwxX/viZiV0/ciwfpZrUil
zPh2NTmqf3PWER8NUnKdj7+f8TOMaGvHQq9Nq0ufJxk=
`protect END_PROTECTED
