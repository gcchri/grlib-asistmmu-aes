`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dv6btVht29iKl8RYSTSBBv0SA4FvYrSS9B0LLibA6i0Z5lIhBsq3ToqqKK+8UQhS
sKPsSNxCc86Yn4dWsJWabTKEfCiMm12W5oPIc05LsSDZDRUL6Exbw1GH3vOzxjec
BeR7gJLMvCBpnLsEL/Tx9F7RNlZXZ96wvmlOYFdahspQdKoLTfknnn2ubRY7opWh
O9PWigYwqOqs7gVumCa45HL59W41GAoUCBdUNHyWnAvhmIAt0BH3aFpXC001KtRY
VN3gwaIWGY4qBg6VS/KRKn5jbTVS7sNXatDGsGT9QgFwXkjRjZLvdF8dlzMQ5duC
nJqy6L9P9Y0l+FiqFMqek6zsA3pg65PWFPHKRnPb/8MGXni+QGIxKyBPgk27mLBG
bPzpVoII8dHBVzXoahib9vZZyxBRuGN1W/gsDFBXrqOXiynLcL5lClILEU/nDqFo
FKNULO2XW2/YXmOXYs6Zeeo/koy6Pwwoktlu6qbAtiALQXOKJxfSEwGzhcny8kRB
OrM7TvMhsRocNL4GLjEW7dFY9dj7PRv8wbJTfFIouBCReEkBnEh23Atv/bOCI4DC
q+qM8ipFzEvPJkkwPheJgoaWCKXOD6KnknZ7axQakhPi1BEArcKD2sCiG3dZkrME
r+WlcoiY92F+cJ1sFEyP7SeMNSqz+JK+6slzCWb8ip3oJlNkjvH5/B2airyLrOEe
fAOpNMCC8l5diSEt3YDhsjxLkTAZ5d7W4FUpoB4+LLfMiw9sp0mWOS8O68dpT1E3
t+tOCRlulLHOJBUcQLAclPxVPT+1hPP+srqGiF59Gvr4Mf21M4asiJytRR5zoF5I
MKx5ZTUBK1PmWUuDraRuLEmj2mEbDYue/CbjgboRPIebVbOwVn9HZzC2+E9f6br7
ocFTrd1hr5sOGXwCWYciYUqYyXSc9n5ltAck9J1lPquFY/aL8KxbiVJD/5UjAhL/
Punj0dJCeLZAJ1aqHYyl8uVg2YZUILKpm0/fKof0dAdQqEY79pc1DqgTwAhweIPe
2u1gDZJvIYW64oWfrlxlPwfRyBgwLJmVVH8MjgYq8yE2pubTYLchl/R4aYDjgIOl
YUBwbRRwmXNi/OUU8LVezftofFmkjEoUtjT0/375QjP21w4zcouBU1Qwrrj9nlcJ
ki/vuzaCziyFwF57JnMSUYp8lB8OTCH5WomfLMmKpE8Tbm7KRzceJueIFVruSACn
9h5NYD7fZzpUcIUXNk+y0ECFnkbMK9YcC18LkzthvuQC/L5GsnAl5vbO4Pwa9e2r
7/9tTX5m2T2bUNpdhLA4cg8Z5GdSb/uPJBGiAs7HsetUJjQsCdqHRfJiWZkF2ZhO
XoVsSI4WNgnP2Au36ID6eQ7sUtUmWwM+Jy0T3Ff3G2QRVnJHLTb1TuYFgKxcspak
wiBgvkqyZ9hPfEqQScR5u9innsQH3LOosDEncRCfb1n5ftrYZDS7owkRwgUnksQD
Ski81drE1NgxD/G+FmIg+DzjO/m5+oj8Esl0rCu5CfVh8tW6cg1Svo7Gi0lbblYo
6sQ7dIfdapYXQ1X3eLuL1FamsxviFKx0eKuUPFHWye3b95Hpwmef5AWp15pihIO7
v1OKLGiZYK5rKzKwzy/lXyBzL/4KRRsju/bru9nW5q4C0ov4RojKqEVezQF0Kcx1
4N11bsIWOg08nfOEYzhfVlAyU5Kf9bhj+XfERXefTL9qyYF6XQ5uo3L+GFG9c7yf
e3NTKVPQQjys6vE2tm2rGtaUsJK/LrqsIvUfCe4Jn/Z+FdOglxv1LBpzpdnwuGiy
Nk4Qyy9DZwayOIhGCghJY7MH46+cS3wSbs1/5he/8Repl3cHjDJ4gIlOA5vrM+Jp
1PjsUTqT2qTkGcq7xseGtmWUmAfg/GNQBoraO+a0eWUEDI4SM6HnmbmO+AsTgAFq
WH4aspph0pZtmu/bkzhOPugBW+goNjDux/F8URafGHrpiJ+hqFrxrcMtsp2BmAKt
Fg++FC6V7lcIi8S4Q2oC0glVCRKQQ3uzcqzKW7vrj9QrIniFiAuxS+NGQYyUVcaa
0Q8w/E4/U9CF2AgPYpGGa8VsbKjR1C772XUZpp+SaNLpfJsBFNhOlrLGDJ2QHm05
t564GSKEiU8a9+g1VLN+nVbEluYc5gR/ulau9j1QD9nXV4cZufaHv4uNJU/jIYFH
810hdRZn7pebs08kB9Qbptu+v62enYtpA+BxLfhtVZjQs/9xqsrbnPvfkn609G+y
RymT8yX1lEmUJniHCHNeMJw0OyxIKQko2yXSDP3XtTGc98Fnqs40PFuactfpJGGt
v7TOK/Jyeq4EPp0rzD/3cRsLRVOXS+rZnZ2DcyLMowRoLTXOrQqEhG5FXr6ZyQzC
C+WAt2ySPl4+Ojih2KJ3kmptrKylZFDCRm5yaqY01UZ9kaR/BINEetn/wRVhAKtJ
1MH8yEWSAzK7oTNpVMfqW0XqglAo4mkQ13pfi/+y/JurHSCedlN+WCKXK8JQGo8Z
gaUm+sWiMxXw1kMvG1TC2aklWhe/5MVAxUP7HKnwy5AQ8AVdY4vd3M1eReZ061Jb
RHjY3DIU67BZ5yQwUZZ2bJX8di/LRj2gKMaDb+3WHwiK1JhgcOp3W3PW+xbMBy4Q
A67m279Ciy23FG0Vwv8TE/NYii3E3Ibs38plQpuKi9jQTPgji1jgGAzfVg/G/1/A
taL3DQ3UCnzbMH7Xw3+NATI/BJ7DXJeAe53a0hmcFQOuAUjGTqkiUdbg5eGQBXW7
XUn30KrC+PctNiQ6u8PbP0aXZF1ObJdfE7ojmaUXlq0k+n//TY73cN6296gTfwpX
6VDTtbdQZMSCjGsmfz7h/8h+nOc4038glxf80aX86dDbyGRzdj/S+eufqpCdBOYe
3BXmViOYsrf6bKK5C1obYDM1w3cuW1zQ9gr7xkzY5ch06si+Qfc3DNwUu24HAP5l
hqiei+SJQegIH44+w/wLdnV4bwcXz/zNFsLh9fyft9R5nbjenjFtH+zrmmabEicR
g10i9WBxU1I3BBzwA39di7gpwwofd824YM3zVDNnWyldFfsXCdP5ORE9VuUKbsIH
t80WkJhURLe2nFONljYsLd9aar6Okp9NeJ7GxJiD34tXdxO9P5pgTNBI4OIH33jw
w8cfTNPPYOhh2KMCgHO7CjvCUCSIWyu0oYzetOViJ/gSujyLGAiehyUI0y+4ftvq
t6Gss7RXxGNtvsTvVH3DGvmJ48xmVh5+pAe9MkbKsm0AruvnIvsLI+PaHoDZE+Xs
IVSN6+Pk8n5SNPpC4vA70REJly2iQctYbqb5RRYg9Qrlh8dpTme47ArsdZIfgt0v
5uUNG2DaDIlnSP6vjbUJs29gjTiCARepkYtZ1X1gZaHaUKeMh7CXE4WgjW6m2i0d
/WzQc5MsYsAiyco5bsTcbB7W6sUowc6J22WDQlquV35jjjBHR6Y7bBnps2hbgaqm
/KXbS1z47BPiRzcpINWOlZvJhNIv9EUNxIUzqS2+Bmb+99EfgJJNIvjNsFkpQZAb
IAtjXt2jGfgGBhRUJeoZuAwfcn3kb57+LIDZ8MYCD3/zAfCGbFARN65mNpPqK8Bf
KOEFHAxDTzJqva3T8UlvvZkgUVju7c98eHcdNfOHX/XrF9lZk6H1z20iIBZ1u1lN
v+gkQUI2xNG/kViZmZ2Kr7qv90ha2Hd8Kord6+IUB385yruTxQLOrpds1FC0YZ0G
rzzHj3b4j7kMqF8JeuU7laHPKFxt1K0cnAHeuhkyzImHVRp/mxsIsGG4oGFJm8+J
37tRXyIo/ePZfB1llX87dO4/8cfdMIZrZWeqo+q9ag1q91lv2ABjoO/4oSH67A+8
8Mk1Ibvx26xSMjXTLSjAfEa1yX71A90/j3sWe3zqSI/Ao0XHLuceCidQ6O3i830E
Pjetc70BhkmwerG6BSGE+0pwccetwSv79jEsy8dEJYRBLa+q98885i3MBnENRZyr
hlA0n7NJCxxYsxLL2UBWaAKAk2gx3n6KlIjJmxSWffAXqQIXB8ShrZXBw3L7rNbH
a6GuvRzim90Bf2Z7CJZm/QDVKtDopTOBudXNxvWs2q+GTNbDpYRzxtvHgcZHmxsz
GvxgX8YB9T0gXh+PvrseatXL0oV0rC6Z7bCM9BAM8atLz+VTfTSAd7omg/PvUn6o
6hDYiiNb1R0SsVBlWTWJtJt6GhTDbWBBWpGjHDwFEQFD8ePxZ20NUs6na4NjB82y
VyQ4cVkU1vnEgJ53C5aBbJSV1cjZXWkE1nd5ql4ZUYgqN1NpQi8PtC8JPl6Dhgoh
18z2MHg55UoVkGCAoUC7MMyMMVnGaj502XRMj2ozlhAVKxTN1k1z1NtBcSblhGDE
PWkZAKDkE5E51JnFMUjs2LMF5WdJRAAVVXLNGOFSUwI9yMK6pkXbVrxxpDvxqBwc
UNYxVj5gjwhlKRsqeKEweNeLmOyyxPgB5YKIuiXTCrvsGpBIqCiotmMsjYjyHrS0
vYNrKouoiU2GoJGF7OIxD7psVYx6Pal97ebGImSW8DR6OtE3Nno20Tga+eivjQ75
6SyzbtLp+4oCDKvASSBt91HWcMufgau403LcO7og863GUOFs5w/LxwJOs2ii2bFG
PvwD2FOsT1fiQFAEiNpOpGbMB8Dc3KCYtFf/sdBCHbQhjYglRq3mZSdEmv3rPPcm
3WR2G4RBVnvOnpEdMliHDIdFmGN0bRqtdSLMKdD0PJtMnPBl3Fb90rx8eOkVdSC4
e1nlZU33n/hnPnbmM7SpQM0oPyPk1LJPOyhbw0KGoRgPIOiuw1dmaF49lE7Iq61J
XafILjN9Pgt38Tds9eAlzFCe1iY+H1ofS8zWoNxalV2+ntX7O4UEu/yV1tj1UO3C
jn6OcA9qXc+z7yOQHLMEbwDE2i8fWwqYXwue6SfLz/15CZsOkTQQPEmxJc1mCkBb
bCTbH+Nu6XXX6W5DGFT40/hY6PNAdYxBrl+jgwEsYWCbP+wnMDE/hAHq+yS5Xj3H
NlZN2ZqTaCLB7AQ9t5alHU0riMM7oiqzH8FbTxobc5limv37XyhzKY/f7oee0pyS
HJ+a8YnzeSud+M/p8Of2MZni9EOMgjptJQV1Y6x+BWESLxidue/qrfIQ/nUqBgTU
PPRsccXPkgd215d0fCfnN1jAiSiiPkP01GONFLBvNPItwe7mcZUZl/znOCLGeWUv
J+Mmi7nMZumFVe5Xhh0L7RTl825nveI8n9zr64gTGIy0GaRpJk5AH/cKKGGH9xy3
umN5GNv1Z3z3MbV92sYr5/pxIBIZvimodSLUq4RdjW4d0x1C3S8KS0+uMa/Qs0OB
uKrO2btiRP6iWFrjogqeS8VNY7wJ78i0MC+Y3L90EgReESuqGq9AsuE2flHt8yO+
Kebc2aKd7Gdd5xeI255Fpm9qCDxQYiA5Vl158EbA5ee+mC6pQqGjCcJPTzHjm/Py
KyN4Ovw9BwPbM+SC6tpRNfOJ/ySexguiLGVFEA4EaWkIiVA+eaTJ6jQhAQVF/Iij
+Pfik/qXSwkSSucJ/+6josUja0KjDTYIxTqgm9+Y4Y7+jCw7nvbF6nipm6dv4I9S
W8fGE68AFvSLMFLl08Rwd0fVS8c8Eo75bWOQ3KFiTFPvcm3JFd3Nb8PHMNiN45Qc
Abe4OkvR8mf3Sh2YDFFGLXauBg0g8YmAJsitOdsp2qPWIZMt+kSe+Hslcn7PEXK0
p6ZOJJ86uu2RHRLriH947SQ2lPVg7uXfOrIEXxvXFzn53qZTHNZENeSPg6qW+ho9
hxk/w7INQ+Hb8rkEf1S5FZa3nYA0wK89CJf8W6yorCIVlW4LSV46Bcw6xClZm57o
BPgnDa2i7EIjkSw+PfRaBV/vdFLUbwmSfuNNl1YST9aSwWqbzqdsWIFrGQjfMyef
Z788n+hPEG9JkyMOFFwTQhMA4ion0EE93vN9+AyLw6vRzKXaSE2PrEFC1QJe39eo
WTpHdflmfdXaMr+esv3Cy+gTnEDgabPKcuhfE47umF7BQ7ps2Rx4BCEqPGsF0SHy
Z+GWQGIJs2gQecoF/64kEKn8LcTietkG5Je0K7Y1iw8028CNxOPZBcT4Dic4oFM8
l//9apxTlOdSw9wrpu11l3zXXTX+A2ZNHhUtQiTRBf4Klq8luiXtXP2qa/sEDxly
cjAgzfnsjhjQE/uPC8VT4FDXqxp3V6Ms8t33DksCjZ6K9qTR5wKrxr8oCIFKdsvB
EI4xwvKb9v4NHB8oRNzOUdKO69rHsQEBSX5qU/sID/dGyo2KcrfLEs6fLZv9PRlJ
rDhL3CWRo2pV6HuDUNC3j80GGJWyXCBjTTUlY6VxjU8oFPFQqvGhm0lnjPBiN3tv
nwT8Bh4eSTPekbEs9o1GUY0ccPxGq25VpiWFmx4s1srGIiqKL1ZTEBboLyjn36/P
5AfnDkXZl8GvfB8fzivFxlvNQixsVzF2L+LevHPr3HjjGodTD21OAnALVstJ+r4n
jw5PoX00rPi6xvxIUXx71ih6Y1vVZSN9lsi1J88Pgf9c60XW1tH/p0uCxcgfNlMU
m/67CrHkO26yUrbZULXVF4f/MNPYGi7fx54i6pSoa1Xeo271OQ0d3kxdGZByLbTt
dWCDnBYt0uPOBpD+8ixLnpxVWPPyRpbFFHr7FMaBEbvTzzh3IM3scw684YQkODub
9WZdBhgFLPQ60oNL4GrDLKGGnIOesegIqHXP7aAgZ+ToddA4uwTm8Bl1/0eHqg3v
zNiAXbiDdJJcppVcd+cF2cbN3a1aTyVysuq0cOiB1FyJr40IkrOVgTd5nFvrDVKX
sloxqH63I0tA9inVk8oEyP2HRJa7Q1LL65XqZ2M7+WquNAGsvoTnMckqXLhaNHxX
IudniJCfJbg/Ya+H9Yi9JkCoB7BHE8O3zhfI8SiPbVsg8x1AstLRTW3IwoNShKtK
/IFiD1ZDNv4yxte0XftFUnCtOJdThtJFDEgV2Sfld87QAtOdBfv1S+Hoo6382Vhb
SjmOVAOLDhsyEn5KTxdrzA8L7BcoU71VHCZePdQ2nQRuyc+IEGglXztX5u1gInPO
zAQjvAyhh3PPyGmwd12BOuc3zlIcydpRtVcZgWbMI3Wit7imRjzJXt+aYK6ODdbN
GC0PNEKpR5RFHAJx2FPWKqjmSUERJ1g64NuP1fMU/8mYcg3RXXWCOnzE2DT3Qan9
p7ePFo9lfCpGQmdlGUAtgAKeep5KxR4JLFCjWDnZXYw/xQltMoJdigEV01i3jkj9
W9Hq20u1v98DlLQyPnuI1+Hq8ohSAb8FciSQaWkPojFegbSqaeTOegVnNykAn89w
xOIIwZJx1CGOugaxd51h686mmmw/DWFVLeaECoSRewr8YWisgcwQKi0IFEbZuXFh
JyAQvK+Kqe34IkzAJWhCKZjOdJPEWry8Vpm2SU2xAkgmfKbyLgwqY8G0O1dWouRL
wIwz93eyiCr0QdVET0DLt1RwM7w7UCDE+27EeImh1keaoogZz86I3XA/WlDoi83R
lHvXodvMeu5iTnprvAx0lS6ijLxAd0a4GS8MqhMHshcFxmKOapRMT50pusvyRYEO
BDuwhwzuhb5bnCjkRdrgIpJW9J+6EZw9yx2x7azhdxDBcN+oeU+jkAcIq9PoDZ1v
XDLv/je1pGm8E8/iNQ9j6ZpPxuqrCgK58RQB1gG49NrrmUxnB54MXlgie7kLCV2D
C0raTBqhbFeA1liCihrNgoByISr+hjB/MnfvAt8s3VHEm05XCkzPzgsOkBq/+zVJ
UAxIdoHfOU5RLUuBIYQk+kvtI3owoSPUnwDjOdlBfHk2WafBcHfgglypkD7og12o
53WDIaBkMbIZJT5X8TxQbkJir+hTB+7IcXt8raDtJgt4/vyk2WF3OpiTAGUnGIfJ
T9t2f8yeaHZ57ZuNXAYoAMYdlWL2KTg1AYKL+xTtj1WBA9jO5rqOFmd/cQ59IWgr
1mE8SFMUGX/qb8kSBM8UC8Ni3UANlOq05M7KGeNgB0mBVd+W4Ht/tXJ1SpFHF3Y8
pEd4NYsyUdNxhyYmRcIaiDhLak0glXpnGhoFWtEao17SrW57Ojl1MxJ+XIGgvtJt
qJlu9doitr4Xxb8+v2QqNiMUsYWv2xli3tDvP7Uf5avSfwgNZrsFbs2mTrfJX27I
3O/NhVv/G2K1MPTwGB83cjrAwfRApersq+uz4X7elpUcG9GdU01r3+ZHjcWvojgY
KF58zIUxx90yNtArd7L6zV26iQTQPXKDyNdt2BbXq6GeaLhbLu9Y0V+AZrVjZKvU
4cPw8D3ldTCREfFVjJlG1NO/tBiyVODKkISaTQq2krJRdMDZ5sjjPbB/n+8AUejn
lVHPqlZ4ca93DMqXPW/swns7MI3WlYlElKefTDWk6wUQM/Ceea8L8tFlSir+dVGU
85ozLa2N+jANdnBEShxn4VGwQemOTk+Vct8JbwjPOVxJBNfxeHq/I7UGCbGJyVYr
6rjdbr/8wZ1UKQ14i6fQqIgZ/us+1hwpobrNRK61TTRTO1nuXCaHJ2h6+BoLp+w4
i6y//Ghj1iQ37IdGMIDEmmqkEf+w6y27prQMb7abc5TL86Rt9vBiqTXR3THMqlIS
xDl+aeWR/XYSFAgz6s0yguGrQhsFG6I/VjKlUUl73Q9crw2VsOhlxQPxH4aJAhLa
lnNTIgrLUv+cdPSDIjzFQvulSVy6xwBMt0qU64Pd/NUoqzjJUPfsP+Nj5R2S5+Nx
JliRnYCZQ9T9YfsDknnVP92HiqUHZHYaci5gvhugDNt0e3l66zNRAAgSb78/tFu8
rQV+83k4aAhbYm/GoAQGIzBJppXz2WxEV8BQxViiyoMpUfEUDTeOwXhmq6pI9npL
dLdWjfRFsBu6WZQU6Q0gC8ogVw2sjRh5TuzvYmbhVzCMkWveH/u8clYcghwum+Pl
86fpotvnZuvChKGJJMRRZSpX9ThH5/dgtHMUFgQ4plyu2rEFo7MByBJMuZyyKX1n
HmJkG9kfwAI4OmyS14wdQ233FHzHqW6eG5w2XZMaHcZVxqUzmYG7i2+w/Cnn7Kqe
gSgcIqiUTbPUHyuKws2igf251a2U5hq0lnz4JrKlujf2pBoPsWbmd9Fi4Es7PwL7
CW9tiK9RJOwjXURXzXTNdTgGriodRSZbj4E8P1NF5gPZfbsCAHM6e0HxEBRsQAki
rhKwNBQc6jZ1qGHb8PfJnYsQhxVmghZMvzcdXMOC6F0K4m1JSsHL2CPu7+nIDJWa
EH5ti9+SUMm01fBXbtCuAPqD9ill+b2mQlI7DZs/ejuEXWgXY/AT9XxYAvK16iKc
GkGAY3o80ta7gFrRVULwVa9veikLL/EyhauDkUjoSkqR1YS7l1CuaBHJednCfxXK
j9SWQ+qCdiDsYc8L5+usUWXkTNQkg+6UUvNBnETrXuKybSTWp93HZBjTY+JIGx5f
Q0JfMzznvnGGvKr0EIlzwCHW9jDOMTGeRGz9oHmT5V2x/4Hw8kiSGf3tJfpfdOUr
QZEpQ2gQLNZ50Bg8DLoVdL4XVCSC71/WP8LNlwNpH7xxRn1KFOSKltERjew2KeKA
u4L6eD3HuJUDMLmDFDQz0UJRY8Cgd7j9CMEbZs46yBtciObGD795iJeTRXKBdLRx
jNk4XaLLkeUhOHjB/oA2vaRvCYOwnUdDmi5vQdH4k6cgfD5wfhz5A/yE+VMX7XNG
O2FkuIzWmlWPAjga2eyTnGu7XtmohCDHS5YRBFqEFj3bvWVcj4baNSPA1ou8nGHP
J9D3Rg29jHdyEXg042tq5NQvV0fPrizStXwOUzffAKHSiIocvlbwY5XyDagQU7jg
CO/6+NhALmcqbdv8TEJWUXfQj+VLGc2QGMvGrNTZ1RWEpBD4stRJMEm9en1inxXm
aVNrgj/ikRF7WW1jK1X/LaEco9LrFD4BjNHNN+e/dfkny1l7CmOHLLSKo4xbtX/3
sFgG+B7AJaAS9awQ5hpysr002k21jNHAG1Jn3RBHTWxFzujt1FXCnqDDuRVWLWl8
1ROFM7QOfBlqkanod10531F4G7sXnncSUr2pWejn00HklyEB/xuu2mD2wVKpcv0Q
lw4r24IBqP2YiddabLf9MqDDEYf3pR3YcRLp1XJsbpLRnY/4v90jWlHmWAzVWZBb
jCUDhAPt435DalQ7f6TKMyvFkIASz7nTX6/6LXO6F24FyH/xcmycdB9DrEcEEUZK
2tU+VkxJBUId9XEKnx3Hu4wDKWoZEjQs+qA75RGtShfxA5uIcpiYrPlAMU1RlroZ
WAU1jBCrb0W/vzc5Wg+utOVGO4n9zKHrAgX48TN2X1B5ISiDjuFL0qbpzSSbcDgG
UlhamsIROTzu8xKRYpKm1hGC8NC29TKCcpgrgfeA64Lae6NUwkBJCN1C4JE/Kpot
TPBc9uMOIHLcIi3r/LDL4QljJsZfo+OFQvgTOZ0chv8zi45lwIinpYfzBQ/b2bSb
F9onTHfvcH615w4gFAOA+2u6MHr+RDF+ObHUpNZWVJNo8jWhwvmwvQDGKszjdm60
8nNWk78D6HMhLI3Rm8s+O+qO1DI/VAqRgh0IIY1jtjckgMp/DTsr+VBmFKATgapB
ZebCQOA73UMzqurOqUbEkGWGsSrk5+usmg4ioInfD+AlHBsTY56ROXhq6a+iXFrs
Sx3X2LD3AuBrSL+7Ga4rSv8fk4jZrr8OQkvXVEiNKkeYBWQdW6EecEQXO+autyH5
jyRQAF56p/XpFX8naDh3ias+1p/Erukad0aiQ9BC/+jgA+KzBvIIW2p0GgIFpNPy
NySnMp7ZORzkeTJ9NpywLXDcoRVDTsHtYsLmUC16av+1/9lYcAw+DojmOShwDWpG
7zeUJ/Gl5laOWLxh/KXUyMKA0JsETeUmHsYn+GDEcRUtC5UsLJrmScvmW8odnhVy
xCDZqnTtXG9s2P6GgEDVSukYQTiVyAibJglTXzEWysb06FgFH6coXb0IguwWy788
TNpKsebN0rQ4kP8QIM4tK0dYZ1TEPbApMnP//IxsNbJF+RISwoYjia7GJhx2kFKe
mCrQWkgkGw3r7AtOnwGQLfcO8HYstawwyoU8g8FAcw0++aX3Df0IKA1l/BkZMD0E
T+q8DnLLntkSNUInzBdzyDMtWR8HOuCecIJqfH7eA8UXfkEsyGYONa8rXOm71ueW
FZz6X80oKHKdg1n7gG1fteo1Io2cAqv+9VbqXMqA1XfWHH36FxRPjcLJ5sTh0SsX
3a4eF6K27hLQqAn7vtvGZULeu2bbPmWo4F6x9b7evkSuA3eFlLuhRB42jUkwt658
uprd71EuYCznsC82L3SQXyFYdraq9UUKuNffs3v0zvcFMJKXfrN6vVoTIIn8vKDc
WNSLTY2Xd5SlnKIpQZsWEl0txcfeDuUe6v17gmsKCdFKPxqI/shB1aTrQGGGMHHD
iX1aIhF4WLFxuXNX5gpNq3tCzeFO1sM+zuosx7JdobNRSyk/Ym1q2p0UcHyy1RIG
pYQ5UkzoWcZkZfmSmtziyfueiloAYys+ns9KbVHUKrMSLLRon7/Hub/Pes+tP3u5
lEHZXTdFhWic0YuIxmPi8ZtZdopZGZ7BIAd8mdBisk12ROjHcEhEICtyVCHFBLuR
G6lIbhSgzeE4jXdyaxvix1ikUyGlohq3gGRnJResmLE1z+x71XZFCJGv3Gq7ohQd
A4l0fUXTKNbCe0+98AyRNrk1Y2b20Cb1JumN5y1eFGkNKjgc12nZDnUMDnzviUyr
LTlyQXfTECzTQaax55ScU2RSxiXTH8ODPWS3naoPe8cQKaQIqelWZ0B2iu16IDEM
a7h4XoG/9BtngUIW45iRzuevgbA+X+GBu8PbjVgVm0ujHG9VLcdNUFilfrP+nzdA
hJprikXMFEKOVIDHHwineCx9VHXXxGP2ce0xuZXnDmVHbaqXscX10fJJuuaRzUrc
U31MiVxqjEV853oHeGgNKv6qZxsna8cFkve5mfEXOggNzosh42MhYW7ds0mnXtfp
QgVWThMQbnfQKBi0ad9KrfSLgY6Z6rFwQQIPowPHN8F/IvTzKHyJd34EFEwXLefp
rCfpv0OpRws32e6S/kijSXFjKpeESV6p5XEAldqFI4qtL48zA0YcM6CuaHV+p9NM
QZQB3R8h6QfINXAAHsRHSZ64xo/NbOeK+Z9e045iqspyBA+p8tbCyTR4d4IRcSxJ
3mjnII+5VjNBdxdQoP9574nPtUxVchb30h2cB6r+qaAnP0tS6FBq1ri5c41fgCvw
YjZxO4Soz0Y/kLVMOKt290Sqwf+Q7zzRtNS/aCO+kpQLDJiF4EllFjKaYAE/UhRa
KwBuKUC6JHePz+DMhzuFMZVU1mYu0s02CFXqFwz4K2zfHlF2FGpiYt2L0cMVHU6p
ERthbdrGuoslGiZuaPhVvZdHNbftIRXqElANzAufb+2dzeAymkR8a5M+j9PyC/73
mcOwzphYZ0EAac6vOxJpY6YXZGqrbDpnvMZNmRa/5jYHMVXsmMp1kEus4yZgOm13
eOrZayKK9OKi9q1x+WoJznGMjdLMm/Wb3K3pFjF8FoE/eL6QIiOl2lQTEdyUCmEQ
bxr/Na3r/hUZSVvLtJbjoNL4d0a01T6BRTqvDbgRrL4JOxjWh8iPmrFDef/Qp/0y
sx+0RGsZ6FFQjU9GQQ6L/mE5V40VFrZ3CJW5ui4udLKl0CtXdjyTRZ6C8giNzfGa
tW3zbSBkWnVzCZM8I9Mu3vgg0VJAVVtB6ZOEO4SgyvLqEFcMLjV9ocA+1/XJEqy1
jrhTfyHLQ2wYtmlxwNYF5bc1pnAytXHY4+OfxbevGrP1OrR/bhVwkhFvuUpc0Xp4
fLkgabqnN+/RLiYZgT3ks0IY6q44p+jYfKyHYWPHzs9eOVQekTWWT3Ztt4GP1/rW
bY1kawKTuWTEXp8LPCZ+YdT7N7840673Q0E3IV0rvSPironIt4JovdWF4t3pJCFj
wv+Q/4+sj36WFS/welf0xcCvywPCJsrqE0v7Xoy0WwdMkD6iyI1KNGucR/E7V2de
iBFVzhQ33l8iMFR4PyTVqJllk3owFjBLNS961y+e0FQQowFQ5AIiWjfWze6iGJ2Z
IOVG8/8WFNCdeSHpZmFg+EHi8WaM/rjLIxbe/2FuVoYs5Yatc7e5+HG5eRcNPdGG
kf4Xe09HUIN1gmLbX8qU1okjmWzLRHf5JT80lZedngqLHeBuOMXysbuQRtotEvL0
QRwj/S21BGcYwkcFKRgM9aEYG3xNIbPyCnv6LK1Bvud7SsRAMy0T4korRtkvoXw7
FfLEmnpts+Cv7UHPt8wzMeWh5pKIFGE+JIOmrQejf0Y1SchHmLRakc3LdBZru2sf
RCv7joRbaFis6jDu6mgWytU2+cfweUb1nrwlIMoUis5uvS3ZOwQulI/kKb2lg1S+
vQ7HWkLeU6cM/8fGKX0EDHQ8gU7UKfd79ilukivK4XUwOk/rd7Pn+REAnaipyo0Q
gNSsJlEQ/XYLHD1/aCRuW0/F9t3sqzGrUNi1Qz9yF+qdR/j7TaCtgfMjzfz942XY
VYZTo5aKphNw0KzHVIRyAssreJ7wfkiXBvm8UwxmRU2FAXvWrv3jEDU7nAGGwboR
BfwgaF0NLD+YVPyE9q7TrCabV8SUHKFuj2GAA6BxhElvB6ssuS+8y8c6SOx3U6cg
6yhjMqEkoGU3gpPUlcXp57fK6ArqNYi/wKtD0tFpiT8YF6mc9opMOiQOFy5+Yaft
8sTSCQag63xIrn49nm50lJsHvoeM8TIMwLlTBI3phG6t3lHv3p1DUwBYPdDIZlyM
D8zK6qaFKbhBXOCNHY33pty4dlZhR/n8/ugHuZsk1jn45hYceKxnvkqOpc0kx1dR
85FvDAYXWRYtI/A1CrCYJJrf7VblG6BPBxPZ0KFUht1u6eanNj69f1SzdVgWzaAS
T+1PQlFzpBepLf2zXCR+xLO9ULFmwFCJmLuEpbYmLb0S8GgPe/JMXHxUHpGnDNaZ
IQSV9Ziv8caOY3FfpvzuAEruquJzNbHLS/eAlozNaPsPOFPCrRIrq5Rl0WqwLAbv
srwgIEEMRKttosEPJJnHIdMSz7bZSJSYmfcUb2jEZwGEGFJw52tefW+3BMos1HNJ
KMPBpLvRTBKhvmZYiIvUw5Va2hd6pogV4rDiUaQyKJ6ubgpQW0Fg/JQiJQJ6cBFZ
n7N8kFQlUYVkdCh5gZ31gaDv1KouYMojJj+wv9q2agZp7WfNTZ9rJKEjViPlEJbI
8d2FNnObVKrEGsrtlx/93o4w5H5JBA2ztdltORbABCnZajOTghB2UPghibd5wmKb
K0u4eTrxn6HIjmtIPIOhkz7/YxSMNUarf1QJ4yT7e3mzu+8aiDoQO/OXnKamghfZ
Db+7ZjyTU5hSR0wtsoz6llmR3B9wHWeXV6vNaF3XhCKOaWK47ib2RSh+pUc82Okn
Tinxuyl744bAu28ozW5Dwr9rBnOwvvqlN/1I7CRSg1lYH1Foc4oQy22Fwu43UdZI
1A3WGqCa6laxeV0N5RsKPWFtLPIT9/7N+XAaYqhCOtG8Iqp7TPeu+gyWvUfDx0Cl
tYCibe6kmf82jo9Cf+vaGGS2Sa5ZpRDj62bCakuM1vaLsbQh9KrOY3idhzC793ya
ndx4u7hgerDO1mvikNaCDP8zpMNjlehCtZh63a3v1h6JMBkz/48D5ZlEUB3gcbdQ
IPMgKXbbHKiP68wdltU2j7wd7WJqr1VNEBi9rqAoOkRd6yet0/QZ3y53UBbr7oxW
DjtDyw9KAnE8Be/LaNTfOSTDSwyuSV5IszIpjEngmXmDRFSF/ySZKZMjUea3DHu5
HpPvZCP1/eQbRGc2kLjkerIakLQbV/S2OQugSwhFjxVno52zNVHtQ7adaPYJPKpX
WJKZTE/7PDh1uWq73w30NWq9VpBq3PV2u8U6bQZbv5Zo44jw7b7gpAFRxLckNA2Q
XgsUjXmCUq+AvD7ueeXzfkK4e+T92yeQFGNi53gmZXKUTZNCaM5aSExhqpZJXojI
re2AW/+bUsjlt1TJZz2WOeLjqb5jzja8opMpNKvhynDqvJA4LjjwwHm5NtXMTPpF
mToVw00FQrK4NP2/cGcuydUejRgVHUqJ4CRx+6noMM5agP4nGfVVTJesC6K43fzn
2p2lNR/iUE3HOCyAwJprgBbzo1TdpzcHR1+OCgqIjtbkjw6VMcUm+LijwJT7TAU4
VwNfXx75oKpfiJ14J8HsdqgSqj6K6KuJoVdUlcAU6JIxbHjCsG6Tjz0GQ4fGQkxu
351mssAZOHrU7ZPgXkcR63KwltuuexX8S3R6Hb7YOS6r2fgw+w9H+4v3BEYfBQEa
R7tXrsj0ilfTg3WV0POW8N2EqudfCW119RwR0/1THFGCcPFV6d3D1Kk1ODvXLiDJ
zaSRDT6xDss+CZ+13ViZoKvMoYMA2xENqXRfvGORUug6Q5IyrI2+l1+NE8MiMxBH
2GVUf1Q4ECnAhvRdxNpe1FRCewcL8FP7d5kDXMcwi7imcOsbNIfB0fk4cMqcHAns
1BPWFuZS79RreqIOfhj51UEbCONaBE77RmVfpKaaj9zZ7Wz/yjLtSxrDIuwxzB9b
`protect END_PROTECTED
