`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yFSW2oOV4Uc91EILlqIDeFVDihYOMKqvFnu+6UgXYlwWq8OFAetu92q7pLb28pq0
Jxp0T5JY1/y7W9qS9SPybX4I29c1RBIyWJ8fUz8G6UUcu5uE2Cpr5ZM5Sq6bkeJp
mr3cQn3z5a5wlY8SoEQlCkD+eBZ++30Dz7qytxe4vxHHHTMKcjVgz2d+asQB/HuN
rybZnC3HKv3QJO0COxgveG6NZoRyXFQ2jUyarUO1TE+OUQeSdz95/NJEeLSwo7Mf
gwG+urZ+gPNYRpUj2IwuKx+5B8wHH0QC2h5mMGTM9rH6FXgZdNyC0n4XjS9vBUxM
oIkpqFd1Wz72okPzXoiV+5H3ys0+iqY2B/xM+dvHXSB16qAAdd4caIgORJjll77T
vFc5J6r2eucuSatXlyV2+7Oz09m0G6hXiVsVxpGhZ/pn+NF2JKD3WgdZvpDcFA3z
LlCzgP2TyBVavCOIRG1Ty545umqklicQM9fGZLM7uBD2jTGDAU7hkVjmvOi2pgvG
V5JR2gJKTtc72ntnK7NUDpXYoiMgQXXR0O03T5Hxblg9QTDI8sD8jamoJQdqNFXO
FZQ3sERCn5+WNDLrgUMH3Q==
`protect END_PROTECTED
