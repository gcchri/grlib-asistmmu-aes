`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
arbxC0hhLoDNj43NkfsD1XANSuSM7Qm4TitucUmeGaR6n2iuVdR50cyPQbBu1oWd
OnrH2PCd1/1BNKkYOjfNRtwg+yNB1bQmikg6BGQQa1wEwIoHAkTMSBqf7nyou082
lNz9rWbTSfbfucf3Qkq3Cy6+hZmhxy8/9f15YnfyTOrB/1sAUJmoXk7nY4rbvERD
TrgSayFopfGM49R5j5Ytx6NdD0Rn0FNQ7mbq+u3cciMcD7bGDi9a4BFWoZ73YRhI
h/i7hCc1oxvRLF9MZKaK5+BzVaOQUsNiJgolFz1sgFsaEvtbr46IYZYc1M7zfKMF
`protect END_PROTECTED
