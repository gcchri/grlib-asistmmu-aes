`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o+xSQOgn0qFg6rQJB5eTab/9y/gzdQ2mw4+bBysuVAP0BWBnrxIKYeszaKU4s6B5
Z8XPgr3sC1zyjSaGDrsDEleCnQWGMAFjvzMTBzmhZYxBgBoaIrUxglJ/3Qy3ETa7
zsgth3I+Yrm6BRDm8AnUQBCsVvwoZd+mP2xs64I0tK+0J9xjCp+Yjv/VnxvIYKuk
ttUv22HhimGs8bP8l8WoPJBpwncEhld7D86HDiNeEuNt6m88/jGF2cMRyGD0zBI0
KDfRmjaOm+aW3EUmIqQ7sMyXR0xFMMBpy3+gOCMvO3FBB8wEAHR2M3p2LtW8Y8aJ
CgtS+J3fExL0xD2BRMQ/JpmiziBhPwu/GJpou6hzkwhqcIwIV5t411UNCJdVbATb
oLQDz8HZa8WiAUSqRXxTYBGsicIBR/rhrDrxyVZXtl7Muo8PrOEj8m9c35gCJrqk
QdXp/rFrcZwLuRaBiXVaRFzb5DTkBgxLoee0F0sDWN8TSnCX0o3K82fdUmVG9Cot
v0V3m97yJ7UzHuYsWUAbww==
`protect END_PROTECTED
