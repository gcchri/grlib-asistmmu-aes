`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p2PfYVEj2rrnI9joFj9W4qOGCosvf7cePHKevAaVbLj0lTes0YLI2CMmg8hs0XKa
pPbwl68D5qh+suK5NXEJRoXCFuYlsOUFpuy1dbfq6ajr49ItfgJzILcAlEGGbwnz
cUBd4pyKjAZcKFOuuYdnZiLkLANxO2Ctv85wHHrF2jmOygl/UjPtr1mPuUDbMo/C
DpyRLvT2J56hugix/XwBEAuonQShLtlmzu7ZcoGhliSoUf/Zankj6gd7xc51wS+N
P+U7pT97KCvvszCvPTyuz260IuK1kb5j2eQAn8aSYbPLLglPoz6epUV/hbJ4wmAZ
IKtm0C4eqNfDZiF7mjAFHKZVhmlnln+qR8hcL35fXHHjmDJIfohF35btnXfmfGlg
8zE6PiErwmRR7ixUTm7znNJGKHV+Kl40OSdwIbWajuxsJeMYBzLmqBG1JkbH+0Ud
CscDhBM/96wYOjqY9ohzTLZwuJS5toiSYzS1xfqsRETIOZXaqLHxfytcLMVLoDV6
GkgzPoE0y9dXW8Fm2m97/WHCEDBHOge8eS2Ua2MZRMDUngMkKKOD1ZcNgaYeyFiM
arxsn7Xr8wQzeyubEjPQ8al4cqH+L5LvS6gIIMT2euDYvIYEY1zlLvMWAiDbU0/I
G4ddzs2tMnwNJrADw3N8BrA1nMdXNcuMaUyL8WZe15u2FA/41fOg7cA3zLMx8WKz
Jrp0a1ABAEhE2xh3X65QoE8alq7/Ob0xOcFzwjqu/TYiVRTQF2c0RYln0BmrxGfL
oXvXh4BwOEk/HeUFcGhXZP+bnfWYMAqYbHRgHMELKAQqPlWNvLPoSpFbr17Tep6M
ze2ByADGq9wiUhM/kAw3RUypzaCh//AhIVeSco02spvmG7akNvjkfbmPsnkoDAc3
/ObPGwwEkclE/n1t84E7tfM3Kn9RZh49leLHjG8gEA/aNZ1g+dC+5+DSebZ8X1xV
LwI9ZdnAigjuX7oaMhJDt4+bWlLQBlXp5Xswb9yzWM549pfwe8AkPQCc75Ul/0F6
VRp9D+l3GojYV2IIEJe3TgnQM5DZtaMViLrrvrke4Yy1zGvmTgXTFjdPa1MktDcW
QXUT8TMWKUl31dj53qFgd+dFm1ovSBWov65nDxMqhjndWqx5BpV9YuGyzvirh9Re
hF0uOOWmQk01RP8g0PWkoUmNloq0BtfZQLRuMkUuabyf09EOtdUVugTaWKuiFdgl
mUVycz+jFEsbZRtN1MIc8aYpReujaQiSrsiNWjNaam9r74Whl1N9w8+7Ra3ZDhP5
6Qzx+0yr9zsjPus8eJkn8G9ZYGzAkHT45aPPsYpzIhNuct1oBqtJSwFyQEOaAJ6a
xyJISvKtbuUmcV6xo7UCgvM1t8zJMX62l8qWNntlFaMhmDxmQE3GRpiTyOtiabji
f/TVMuDVVYOcocAoch6OTwfrZ6CkamOOup4kRkInz8QgolI6xMwwH0EE9yXeklNZ
KRK0sIWBKfFbuXiOsOrmQJUUeYeN60r6Zj4rJBgvVZSh8NYancvFWcdbBadebG4N
u8ITn6Z8nRm1f+IaRxMarBe/q8b8T0p4kyI12murdPrDQXCfX2J1vS6kQQlvcrps
YGOZS7dUndZ+EXEb71pQ73/PAHj+PhB8O0Y5Hyeq4k7ZkQ3peuoDXa9VTtwGMkG3
fCtTL6mQFepS7tiFHRkjRH0W0Z+FSMNaN8YUmNg44XiOR6seUU4IFazf/JXmAa44
9JnH2tamFxAiruAEQTl4Ptt8ai9wrQPffiMDBIjQy5ghzUVEe0s5Yy5VnD/dhY+8
CwkupeVNsNRdulq3Xc5qBVdmia8PrHyk0CwqEWXUBEDeVYO8sBw73lNHzPv2f3RN
XNTNO9rKyKGltPKYuEyTabgTYqiT8q03egkT4mcVMH6aI/p8HlqZ2VeS5lAU4r2r
cyciv+FuF4JAaeKJooOTjl3tdazMmTUdda6g3ZiunuewCQ4htWAe3YXSwUF3ElDM
rcaDJ4+W+kQucxGPTxbSVVgEk/vQAL8GKuhHpjXcCb70W7m/EiWENMG44XkQsldg
yOiZ92QQ/JDUJzAmFPbOU/a1iQvq4q8iwBcVB2znUBF07ueUAUOHwVn0szKwj5rY
ulGUJ2Q3Rl12SEPu2pM4mrBHYT9enOOy8eiAx2BXBCqUXXRXiJX8A1nMISBxfJE+
0hx7W0BoPoPiD0XqI9d+fM5VpAU4cmgDNVOSXZAp9JGk904uuqx9XtMoSxxcLnT9
RVTC3m5SW7JLWVG4qdG40gfGO0aQS35sv2yoAW8QIPbap3e3+2oEd9+oHT9ScBxK
3ZjLeqsHXRSOgIreeZoEqkLAduu4d57YgsYPU8sK3WZA1nbNzNLk9MfeBSTD8o5R
6Ia0DqJ0m164p7q0PpqQG8YVs9IRaa4asbhTQMAG0KZ+965CaArInsVYdl9GLC/F
EjDWZ55O3cwOtAi1j4Ky4H2fixAJa4PMMCyXtbYImPByMQikJS97nLgedrG0Zl/6
9ChZ8MBVxH1nloXxhptk1PSIpmiZll7ODbCxJcNLDTzJiHUXAErNr2fAd5bTQVG9
tvFnm8GRZUcxDDUTlhyxmC5Fmsx3yrsRz8jNlkE4Aq6noqR9yxyKWidSx/lDyWD5
ztsmD4fXjtTtthafNfhx8EwfK7QvbwtaAdPF8q9wg3hDypKLv/oFeGRuoz8qcVjt
8r3pzSocbE0aAY8vGih1dt1QzPXB4gByHzn8rqaFnDvqNv1QcneABUcONF0JPTYq
f6A6lhCngsiTK9gUgC0yn7iDwI1CYF863L0W9ka/1tPQfGDD0kVeEgb0/3+F+Wfk
TN/XPoBjgCj/KRWlw6mjVw+pW3JP3rhC85YC/oEZfKqQqr0ZPTr7NKESN/wGJRC8
1/kxiGl0IeXMd5gADhguYMwhfU6x+fbFeRkT8Is/AvdGaY2mykj1RFymRnlNI2tS
gyq+etXo8/7w+EKeuCWG6gQ9oNtNVqbAlbroSz1ZfUphDj2tANBln0iK+C/ne4di
DV37QRuOwe4EyIcat2RV382+l/ahh3+nM97q8VbguGvCUKHnIKNf1VuDxXivbqgs
I0QbYzsHDUVDcpAfNj6qGaOWtcJC7NKVS3R7bacK/o232tI/zCkXBIiBECDmHA2Y
xXuV03H5uCwU4lQn3uEMdFluilAh/f1/RSCQDU8wXh1yPsoahWj9HTRUGS+pdiQF
aNv8kk7Iis2FQ+T3sdrSb18qvFpiun4+GJQ7sZvmN/8FCKyxqIMARaHN8mDY53Rx
J/D1+qOP8YN8llwIBC6YSIxR/9mk6+l/rkT8UH2R0RjK1QaRZewJtcSXHip87lx3
5Iq+wHACq54GNUKxpNl/M5pm+eqYYnkptDTzhPo4t1QQO4iQRgzHTpxVyM8Pr3XK
A0wPXmaYw5Wth6Kv/gZELulEraLazv06iHWxanhXxcTaZvoALrCq5ld4rtu+hTdk
vXsAwIJToMFBKrQslQjTj2bdyAhdl045X3lgCHLVQdFn3EHImEzSb0qn1u8sIsvZ
0R+WMzWb1oKOFCKNvEeEgX6NEcWl9itcdnweXU6R99Oe3NXknT0ttsamVyZ0s4bX
xALzxDFStgLBJLE6hjDPYjaRq19pF9vs1P59t2WYLAtoWizS/+oO2ZipwyLKGH16
nk0yho5xciZ24pKzNunD4+GRWetNiVogmEndPivyNe4=
`protect END_PROTECTED
