`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FjR4ogfUg8vI8JmbPAHesGXa1yzZpMqaL5EO+dQN9goQOcIgjd0uQyquvTC5hJJZ
9Xa04vl7XLTPIdcuTanCHclFdhFpN10vKk1ZRw8+gJOCW3IDpa0FIAtgv21Mxs9o
ykEcUpWY/evxhHLl42dL5cD7688p6ad8Y2+34HRHyErgbro/EcWt1JRO646+/DpS
YBmlXQh8L2Ou62AOvXV19tjwsthwu8AS1qYD8DPeRzBfrB0Py1pI6mkKnKwmvY0S
FaUhDwGRi8V9qFF/68YHP+CaxZZJbUQFqvPsJBLWWGACsYmD4AFkG9gdxYZ86eUi
PvK/5/9NS7TtskK8hDr5ydphiXJ30Oo2ziZHCMTfoqtf9lp0RlzZwU1Fr//gNNGi
rNI/s6ov53g6hetHB9IpYvnAvPJa8nbFQKagtwAjDez6j+oBlf4goZ6yWCGQxKah
CkuVZ59etHiqGmKL0cUwVAsib+gNuT1+nHmmh6aikBZrdaOzgVk6bkEvEk3j6DcJ
hOJgg6TWj7ioEfoBzrFOEjOq/wt3khUIHZBKbnVaA34ztdkRzBVfGI031FGdxMIE
zXIzWeYonmMFiZibtDt6dVDUrTCqK4z8e54Bo8E3qxG/d2/sqNpapSgveyuuxXmp
H4nlMdkmvBmFBsyDUE3BHnrNsY1L1d7ErP8pFJUdquiPkyy8jBmz6VzXZTnLtMRm
lCVz0i+rJZWNuLCn9+LDpL+CzmkmYxCX2IuSO6oPgRQ=
`protect END_PROTECTED
