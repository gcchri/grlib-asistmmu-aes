`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rObXkek0cNcB3kz+qc+T4yMlqcyKLlcs78ced6CJwJPavT0iOJUfqiCLgOUd1aYV
H/Hwd/oXcXNEIlITo8VIsW1JdgNPwB7XBKAUgBtsDrYEVnrVm1/sGoXBanaIUSw4
omPoVziPs9vR7ckfWdJpZjj6+p/boyuq7GRW+rZwb7x068sT5F2N5qRyVAQxUh8g
p7wJFHP3pGr/e5Q+f2dleMghfZt2+GdsFW69jAeiFegbH/NJAJ0ftkv4UlxzNbsl
ZycTlpyj5Tlu6q7fZ/86tRt01zjxDs2J18XFEViwt0i0xV27h5BSKhmR7lc3vrVE
pzPnUu5r/0wTmB5q5GMa5PXzDSGAHw6tdGLPsd0yWlX10wSqXiJGKr9kPYhxNQJY
3/4+MRwp3pmOU4+ZqGWmvMqfIMJFfML5/PysQCCpTTGm6ZJCFDHMFHgmejNGD6X8
WzTJIbNRz0cQbX9vsxVD3B3qrEKjj0/SVjX1vrw+FpZj5opiKhyldjZTptvspDZT
QzCZfDwdjFSC4TADd5X4B3TXj4jf5gA48dN0rS71EHF6NYYe6j41UwjpdF6AXZEs
mw0oWmkpftX62W/vQInlXVwWfcAHsS+mZ+0OL0sV1ekHl2NMVAwUf5vp49zWBF+9
JVyXPXt9EDM5zbPJYLkE6K2a+fWyOPXH5Xlnxb4+liExTw3VHkxDHhutdfoxrOVr
jJ6AD+1I6WL2lNAslEaBO20nI67uXJYhoN4cs5PTeS9umuJzwS6J/jT/YZ62YpKe
hFmbts7UD9mDiw63Mr11+E8t3VlobJrdoMssDtqN6oK994R5Q4PL3A0QkIT6cW/P
9zyCA9/NRd5FchdfThuJ4IJ1xc7AAjdQ+5++vT0TQh697rVOYB/A7zbGgz9OGi5Z
4IIb+ZdUmdeOdYTUcHCEuRGyKXGvDQoMwnPdjAFzQczlUEDPZGZbTli9p5IruY5Z
DdrJdOd4Douazrcj5gLDAnsEQcfnt13TwqEbC9rrr9yvFeRlPliiJhgg9fSYNQcr
ioIQDLf9lC7AiOW22i/RWRq+UNyhTBJRxGHYyCLL6/Qn2krzGpMqT922hXvPYmb+
lZCP5S2KVYtBLylSVj/Sz/aAxzc/zmNuFvPOmtNJz6JJ2iKfKinooOVV8lx8TITt
8ujB1jSZY+2iRGMa7yqMwp+lv5OvtP/mQuihARd7vMorh45jAhVwPjyOO4r2yPZA
psKpuSbjbvzT5L6ecIwF7boftiQWAHuqbfLg6PZxbKhjliJeuk/L6luGNUmFFhiS
37eeypctsVvC/jSHTZMA9XE0t74KzwHC6urWr3kN7NM9ET7bgsKSMUNTaowDfsqv
iVvW3WhQiOLtRwEUlbKpqwIf37TlafZeQmbELnLDlfckurUmcSRhHQXSjwpGegON
rM2fUQxikl9wBwXZic4XeDif0jqR8Cx1Pd9mPD9HGrXSSTYw3Xufh0esdTkfRVTb
6U+OgiZ/x7Nz0DeD7qWQHEQIEzbP9m/4tTII54UQfr99XFsRT3qwXBen2xRsqtl7
OLYsd2QCxcB7KwPb1oNMdBM7vR2a0/HM2LybkVNFWyTOPul3OVPxKL22mIPgZ95s
2EjnLshFCEDt8PJH/B9fuWxoP9ZibBMUWduP2An7qkCUzqvHMEgjlL4AWrPrc0ic
hGA8XZ3E810mEl4lFbJbo4RZrZ2e4HAEx5qSvdKHaWcjGHIJdSWiqPC/q/+33KiB
4+Zr4pOSwig//pRbZkK/hWWj6shU8DB0ZD3YDvZXbM/TuUhFuyakmWKPuPH3QeFR
M+eq04EMMs0s5ZAKurisSOPWPjJPHsEDewKQaCOJK7iBIyf2XPGZAxt3axxNTdUU
mXAMv8e2UTODww/4Z22QApxR5wP2WIBLrKDhRGXjxqq0SrU4T7ZH9GnH2Q3FDeo/
pB2Hj0NUWa6khQX9bdAMAq6KrA6pSBOhNCibV4TB6QarTxaxg0PviQJZb1FO+8oP
38QJo40nkBkEFwmZaZVnJwLbGOuJZ400IEwfyECMlcfdVG3Uo8XP9kNpJCNxBKiC
kOKn5zg5JiDYouTb2NSeiPqt9naTjPu/LAqSCjPR/v6eBSGv3lqKBFnpFflcWghX
Q7G27gmVkNvs44PjkH9NmHiGSj7GQkgyCDffojD8kxDs0bcCuCkXA4xpE5SfFPHx
s8/KW+eKWh03SOjn+jYr5vKoU9SVClb5EsYJRhp1qPEGt1m69Ak2C62ARXqDAo2z
PeLIwFR1bugqzuqO9HznzW1xeDpwZMAhY6O/N6zvcTyo2wCIeUBv90NDUtGSLJut
xs/1Fa0ksVGA8gSSgAp9bX1p2URZya6uzKZlKpokL2QYxQ0YBMy24MInjE/fFFOG
oDj4Tkj1ZliTXEh2AqwZse7IDfLTvkTrzyt4fFptwxgFPWE7CzmhWvynKyxUll/y
SIY12tN3g5OmfGePCbkupsrv+yZY8KtrpcVyQrTTtyNOIPrRYxLCtuzHlmdxGXFN
Z3053FYE8X1qB8MJwrfLWe3UBDVqlf2r0zBVg67OSWfRpLPCoZR4oF/wsCsWPL0Z
c4+o1Tdmb1oeXT2DV5kbIAa56yVcQL/iLWmeavY2K/UKTVzzOUVAdnSSw3NlWa4h
MOI8wK6bvj4LhZ031wr6PdCeghFU2FadeYpMVngSdqQFVk+vmyP+5w6yCjcMecUj
Qmwh8Z9ysmjLjUlBQUqERmN7MI8x4oAtjiKxslz/NlLhJHGLMZNl3lKdpcRJHBM/
RS3ydn+1ulKhZXpjFCXtvMFjs88YAwtODqWGcRgO1QuNDcBeckjP+YAbEyggByyR
6gTkPLHQHcVCZjvE/W1wxXRyLfcHcZX94GT6JZHKw3mCduRmhj2qtIp3RTKVa2r6
3caaKcKWad8cE9bYbNgcgXhePjqFeo9frmZGYRw+v+LWHWA4BUBd0FBr6FCm9qnp
Aa2W8FjANVyvdlRtoAkPXHwiV4BuOmCy2JQbLGNxk9+o8dT3BYkto7qFTmR4B9pz
w1hGWj3aTOFkm+OE6PHV5ZLxlFPH8GZdfWK9381VZ1o=
`protect END_PROTECTED
