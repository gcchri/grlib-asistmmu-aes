`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zVwXuVZDx2kmGgqjrHgsTy/uS86CGUnWcxgQewlBrFPxHagqK1Y05hD8lGoT6v4A
dmAKGEmQfKNko9Zqyg90dj+JXG7V3kDXeQzZezfPjAuO4byiqg7ni0aR6CFeWT7a
tZHXS1mbQqz2JgSQvedQdzB6swt44gy6X7jEvg8RAKVw2kclpgC8BII4YsMZA25D
g6iTw0QEhmA9blOGwQCDH2DM9XjRZlzSjj9O0kvdQUU+3WcHDdvXyxqAbmrzbfi+
7cz30SrLpklsX8xc+Rk+hGPuKoP5hmEafldMIlsr/6FPPxQlbS+80l/xC+jj+orD
iE4FHUBfj0Ml+Vy+ejDj2/n0n6aytqPmN7BCjeCjmYS5TAg0H6gr6o8GM+JKzupS
+MEcgFWoPrkFoNJuoc6fZ/dYQg2jAjJ3VsL54YPTzoGN9oHVIt/cr1R7QemEWTgh
gCijuLHeg3hWIMGVUfpnSwvaekvTd5ra3spNU8rdVBhRtYGO+uzMH+mRLohKYY9a
2DPGHWyE/JZvsNajXpmCO3zjEsMCZ0+usaAfNAqaHO5cdU8mpqpMf5krkFmuYpoT
lHoBsXtucQ3nLPwWu60lghfYfj91TRrYat0P8I4C2v/UfIHdyqmbqASH7FY/3j50
NALA/XWpcHjZTv039ZNXUi5+6VDggZI8Efe/xrGfwsZoFSdTdLjzm9CfXgGVntoZ
Lgw8zMcKmmyCJ5jo9s0NBA==
`protect END_PROTECTED
