`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/lqBwFhVxYChz0F3pblFkHTDg+RKiNs+WJbWujWCJQC+mpFkcjPSkpJbE3Qpg2WX
pEWe6gVOVwAD0mnZdj5hTxSVgWu32PlaVTazeD+onrtbTQcg1uJaBo4f/n9EBYt7
Eaq63YQHAosDDn1SCx4+1YDsnXUJjUuiOfyhIhHSitaVRtJZxf2ZGSsa2m6zzHAr
Hn1JxhM3cJ3lfGZmUetejDt3sXND7Rdnlix2R08sxnOolbB9VfD5vCs8C5Z19nOi
KnkLXgMnjSUI/woQMmuIrJY6YLM7r40v1HmxNfWCkusonqySv4LuP3bHaCTz59tA
OolFFU1AoI4EvrxNmHkrkH3SHcRaHURNIVLgNWERxbvk3IbxVKyE3FtGFsRssg1u
6gTHfbr5BdkWaZ2Gray3Dct9twCGmpyc02GFD2o4v2DIQeTu3Q2QHlwS/NoDDMBN
V+M47QvdJIcV5rDbD+trFHHcxvsR6kq0+9Mvidpt9u8=
`protect END_PROTECTED
