`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9ScPyVWncly5F9j0LL1kKJo0FUkMhpXSVz4ejvVJIsb4N3I56zhN9AWt96QJQXd+
xBjJKX5gPp54sqq4zUVoUq6PD+2WZVTIXp72/YzhsaCH8xM1g+3xwy85roPp/gKF
+LJlkF4oy1+VpWL2DPTniHgqokmOs5wDaLGweqetiRmRSCfD9GdaMK8bye9+2uQJ
BhmlDONQBrbQ1seildgoD5PX4u5C8PhTq6ILmXpswMcw0N1xB/ObxKVkgJCdKNB2
t37QIuxwI27Hp58QPk+SpGHnxl27le7mpi2QleIhwW7QHsRUqhxJkIwp1g0x2ctp
+QJdiGw7KQJfp7ftt6ypHV17+vGK+ZEZ7fmhBGKRr2W8x9+h9PGDOApl9XKMInaY
D3Qc4+CQh7D1K5T6h7DqlQCl/e517e91XOY75Z4FUmVwsLvbtzqVon7SzlJBwyDw
wvkYaYCCE35z8BJqf5ZHqIWfHYTMV1AMYnVpMtngo7pmY3k2qo9n5qvxMKgbs9fA
03YHITwF1kQwIHIPqMKC/QysgXmPFHB0DlgOmGZ3Ye5LtWV4ZBTFC7I7wInui92s
/TrTJCOPDQ9vjbekOGHwqnxTxabykAxP+SaeMVxiETD0ZXgk2df/6LJ9RtaSfWfe
bh0vAg8DR7u4y2HhTN6yEZ/wTZ51Bol3zeA3WPiciHWNxgxzNYPQRI8mAlyT6Prb
2gmAvmeZYOcKLD6kjZ9IEXSmOoW39hUgq4JtkR8AsOjTLa18fXZ7v6cJn3Bty3Oj
mGJ9OtrlpZD27MEEZfY4Uv4ISWyTGm9ZipIGXVW1f+HZCcs/sdmmxXHY1/ALOtit
mmHnILXFVsvoknOiGL0AbnR9E8p9udsEKI5daPkRwLBItN3VVKtWK33+DxXrmkDo
CouuucNQctzCgmbj+uTh/poXeM1tMTbdOxq6A5E0YQsSAWkb1fX/v3vi4nXMeZEO
djr9h3YLVFRTFFCYs20BZgGYwn9OvgQmxYy72IQbK4nm4b7iA8Sh1/ZMi2os95Wu
VFMw9FMQJ5ZGgQMREV7hIPc3BwUuRViSBXkUUF8HR7SAwYunavKqL54/Z/JA9gdK
fQxKStwC9OzjT09+0dNlE1VahVTF8yTmRmYZlstxpeLcn3W6XbHoQbUFraVKmddm
TS34hi8bd3XC8PqS3GzH8equ3430c7jAY6pGwTI6erjLRzCBzgjE5dc5x4tNyLFf
4xoVM+qWJnYdJFfT773j7Ho3JLlzmsCj3GxX1QMhcucpFEnJURF2E0CppMwcRxG8
n9W6LmxKZs8C2sYyZymNyuQlIbrA9QN5x7yc9z9dOlAycZMOK5r8e9MyMJUfNLcD
ixJyQVmH/GOkH1UqXc9ExoRf91JH0nN2oCqkKMfJJnc=
`protect END_PROTECTED
