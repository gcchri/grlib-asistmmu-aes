`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5qnSjguVEluNpcqc0qQLNRM+Tci8lVZVZ10nfjoT9way03duWEXBrtPICGE/Dq0y
tIQht+QCiy4POVtSh+yIgSEHt5liq89rcPpAaF9cr6ConPyrhR7XpeNdjOVEVPGT
sPw4E4Pha2YY8atNBlAMs5wdAr+7cwfbnAC7ty0PmdLJPYOZiwhqv9ZgNHgzEOhl
3MRDrSdlguohwbH+qnpRgPUMZxpled8hFjZJoJVbMDiW/Lz0uLEn7rN+tzO/7wjT
TOSITocOdlYErESJ6nSb0FiO3sn+pTCXDrgpT1kiZK4=
`protect END_PROTECTED
