`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PX/TX7trDZV9pAI6cH9JG5TLx0Dd6iKiok003x6bocvjKmpyLkbD2au4RhczRUvr
/pVNeWlRTfpnDNVbTsw6x5tNbZHWwCtsM9oA0JOvh7mMvYp/MbVb/JiPt7onNwoH
rqIEbZbjpRAfY+Th5fGrYfz1cBsYqIXvUkPXX9CgULdv2XMSJj0RB/oB3mwqLxwC
mFqunNaugkv7xT4uACO0zvomwDz5FEdMezjm7LLnbjV2MsFYOcHxEAcQqOp+suUI
Pt2KTWoWHniOKB7AvQyf9OY8pkqzhQ3Y2mXkCnxPT+IMTAyP7E+Kpx3w1G7VGYSu
uzPYnn53OdvrwKlO1L2/sXHSb6Qk1fCstnq0/BFlOhVOhzeyXqoNcdtWRfI8fLmM
zCom7OFNARqTEkcZ1h1AVjZ/zsUXSgGbKP21Ju6zxDxRRSad7Faug3DrBMzC7R4U
GY75t6YGbXHS/IDN4heyHY7K56NkbSgF4WjBoP4Y6XzQGpCnNNhgDAWxobC8PrxD
q2oI1eVY3iftK1VQ9Kf1eDo/oZRAX11aMBGz+FW8IhHE+DxwCZjM65G4j7m3vD6t
hw1hW/iHTTwL9m0uui9Yb4oWj3bFR0g63QRIuqqEB1828VIzNSshsloX7+04aI8Y
Lh0Pg4cRE8SzTI3m9ZVsIVu6tWC1oOn/tZQPUM1bfrw=
`protect END_PROTECTED
