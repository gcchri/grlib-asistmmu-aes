`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vcz3bg4u7uYNqhnWucYvjkEuxrBTFaKzFUV5nl3YvMxP2+I/ACTovXS+ukvuAOwO
/xRNPHWCHdsCHE8cidoN3dqTk2AZwzO/eKs5Pbsx3FPY8GXHZPwtb5odvOfcCSBl
Qu1q1Z8rPHRxUslctDdxWyWY5QJ5bjcPZztbrfxzUVvqShCPGLtjequNINE3BpC8
MsHLv5EYVVH/r0OHXRizFTsfoxTKEo27y9fro9IZrlKsCwXcm7bC9lrl9/3kF+H+
JG9rT/YvseuxMifKNwHCI8+IZiNShMgLLXVzaGtK3verkEwiDKxHpAiykohr5oFP
I9ePelvIHw+N+WAbqdLarJScYsOc5KNmRZmM+2GeDfiEM5fIV41PlvjgGJtqLOR2
QG0gDzJ26d6r/cICpzTiBwi8Gbqjo9pDZFuOTRKqTCJM/V8nflOAHkc8fHVw1Jwn
uYtOlJkv/vGEkgwbGjjpTQ==
`protect END_PROTECTED
