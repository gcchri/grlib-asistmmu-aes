`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8qncJC7Gb+xIFloTESFTlr7RakwuNk1/okkQporul8g4m/QhVbXBDFNK5PG0Acsa
ideDb0z+J4qfsEZZ9AZnlVFIsEBJeM4xdzXLXykBPP5/RVx62RIvDTbgYhQzsR9t
jHIQokaFm5vHJ9UrsLlNbIHEPVOnoKBf2vjrNOzbg+FAfoRUHWOrQq+tfz4h1fEi
4fj8yRICjV/pHAkJ5JRzoE5H0Z/+z1d/npeZ28htHoE2Gclme/ZU/2dpfcGL4YUu
exMAzs4VC3RhUZ4caNmNTAihxDyI/+td9s1ZkXGiS5SY6Jr5/GIroCjZLT1NxNwn
SB4tpi6PUnOhAcXQ1oH9B0NW8xapnd9r0ygE3RI0tIzLzqQotzhWutmhV7Rnn+CT
hIA0z6xwulbDUegYdyhn2/g4WYnd3Q6Q7QVRNZ6Ouz5a+bri+MK8u0g3T00bMkjV
iTyTIwnadE5oezuVBnFUZeX3lLtVuoQigYVC+8x+KgwA/p2G3ibpbkq3O3oa+pnb
RVVKvK+DGcaNcIogpPZ3y+a0lDnJPB725eWt5AejU78mih+08169NZ5fQfMaXUEe
c/h/yxJQJ4jaRTvBYCJ2fr9LxlT+9Wf/D6hweGX6LLqcIdOUqyJ2+HoyX7bmx4gW
IYMnfDbEHjSGgadqfWQciQ6lF1jBYMnBlcXZUQ30HZ4mA601K05sswRKk3+Auexm
4EhLiI7FmthHpdysL+8c1Fx8w753i9JB9dXZYYmkxQhqTWUfrAl89+4NrND4psns
n4psWybWxfU0Fv4xa6K7VYqsD13vFDJ+CqQDcX1It92om9iQVywZcDYvtlowv+3R
F6FMYjdC/efA6P5vJ/ldR+u0QCuZ2ZxW/2Xbg9T7gLueeClgQA2rAPE9EWhdEn1/
SUgfD/ZVXYK8AWRTAY2Y6uNnqZXHrEYXZk2CBnje4CV+TKE4VzZlFsN36PkAZzdP
VxAED+aEoXAcMk/Mi5Hdhe29hjbhVfvhiQHkTNU0/3v6SZrtvWTyKpF1MPQh4p4l
tasRIG+xnGREjv9bsj+9R6Q/9NXpgyx6IBCiBIIBJ5w=
`protect END_PROTECTED
