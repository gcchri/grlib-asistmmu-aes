`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ntNlfe6aB+L7TDSDei2NCW6IZBTYsjZZiB2jI7w36WfgdHesFjvPDv8ircpnQLvx
pgKm2EKk8211l6KxCW6uiLK8v8oWXLrqFfEvNx6JqG8ju+39mTlZG9AFd7vXDs8J
hfqeX5sq1IT0ihbOg74hv77/Nipz6NgkDIYPogFFDqOoVF8RTGf6340cF7j63qca
CFpNhDtvo6w4yBlffr8gz7KMXHnNLPQcykL7BmnGHYG9t4kd7bdxug4KNFfpIomT
3g2Xd88S3cPeUHYlEUrPFReOJesGOTmVtRAzCGTYsqZoZLrZCvbxBvFK8popPnIL
KnPfp872UVMPb7jWw9bYcZ82+qHGXPBgxUoDPY6DxHE5/vG0cwroqF/5awjeJuCq
VUByg6MItm/99hQuBnkgHFc//KyLqEhtkeV40mHnQYPOjJTaTbdTs0s42l9IiC10
cxlqJhGOi3qrM6DxSL76t0I0e6cTEyiw9Q/Weffoy9RzP6VrQGh76P+fK02eD3mj
`protect END_PROTECTED
