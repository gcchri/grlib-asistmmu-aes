`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vD1rYw2gaqlROCwwOfTcRLypEGIDzwLle3ZmlWBlt51xWdDED5Vpj5Vhj3hRXSmd
7LxevgLtYC7VlOwF0iHEx+Ra0t+JOHs4aMJr5gvI7pA4hZW15WwcfLODLKQYXoY7
3CWkgilPbY7ww9Z6CiJEgsrOLxKsiQyCQ91lBPvwTvmjNTt8u+haqHHCezT5EBpk
+M+ESg1Hi78fUVYTaJhNO4HS8yfE/R+HhuHA1mI9xV3TsY1YjRAYHPW8CZJeUlPU
PgYLK5g0wWrzgXRcZ0I8LI9GbKcknBKSL17PdLSPhyF+1mRgTL5K4IlQscMEz3tN
oMNjF9XRTBZbJhsKrmW+qmhL0d/xDlUyZDAiKbPYxtrzVtAYOCK5mIPipwrafPEp
/VxjeeV8XWN1h6jmhHHRdGYyTTJBXxzCf9qe+CmG9nSSaMQI5AIeb+LBBVVUQscA
ZQLUiebLWPfqC0jwsQw7gTeYafDQn0Lvi5kyxr3SHMNr5NZI46mLN3upkOUyQuvJ
wRVGeiUAv0yN0yZrSKP4VO7t5KwiyCEZcB3QGkC31FeiYs5s8m82bY6jwksKFVZR
0XrQCD0rgr944e5HVWuLnluIscV8wv64ejt+PFbUYECdmbpn1jsFxTY9jcpJF7tG
2QGf0gHZVjT9vKWeHRI35+thVCeFGo9x6g07DdhAYVVF04ce9y6wFe61Ilnfsswu
8KyvEt16JBAr1s64XdhU/qLnKZ6Hdgd4ntkzwzlyJEhAFJXTrUDKJPIlNojESCIN
V0WYV+Fp58fhxDte7UHRzkKO6M/RNAfjYlG2woUDema+783HBuAICa9uzMouslxf
+L/proVCx+poZGwpxs0pW28Hn5gpfRya1K38CNUL34pYsCiTjYhJ8x7RR1dJw/SR
/VvyETKcuGJj5bzLJpdZa4MjD+gOlHdpLOrb+/ydI5C9cis6D085dEdTzwCqmAs+
Oizu5HylfV9aJiJX+rpG126BkZL7eepB64vStUeZW2Mp9eVwRv1uqQkW4LW44oA9
Mw7OmlqkieMpwGtiYOBKj6bBNUOfSxCnYsjU/6FKcJ3Nq0vtZ3NPJuc5Mtz+BAEX
azPNyUKhhS/hP8r/13yolsYcyK1ijRtQ3MXQDP1Odol1UOzd0NjCTMmNXcCuzPBk
h1wbWxkX3gsmfV0617A+7tePwggG4Szb8NHGOE2FW7ftGAdRIgIZ4WnhJjz0qf29
cnS4XHEBGBUMN7QuhP2dIb/xSlNY7yZH0ISmg2PDbVP2JQcy5eLRPFTDwS+7tihV
RQV4MSbdTo3CUeCp/Vyct871Kqy1qpwk3pob/BYwb62qm1lfILZqHN8as1bOOrkA
I4r0aijI8m3zrdobltfyl4fTtMm1SlkODybuj9kRpKn9I5fMZGGOFVBiaqPOV93w
4eEqZN0Xw4Z0R2ZyTOBeAqteZFJfHWk7OJgl7Bvw54cjO0KsmT7xVkClpUDttrLu
BVPKTy4y/Kuw4zjqFMSHjHK82UdEYXAkHnkmSX/Nbrl4fI/xX0IM5kkOBOVXzwCy
cYhBWuyzdLZWJK4yLT0cwDSPpMCpmnX2cm2kCYyHNtkAQb7WoA3oUilQ5h1cMrB9
czaJdZXAToFVNk7IX2kqulMbdbi13Gzj5DrgLUbC/+0xs9ppVitFAfvVd25/Qf7/
1Gl6U999W+Yosjp4QE1XcGo5xc07WkW1EYFtgAX19/YB2AsAkz325UdPEz09dZKP
euNA4mJ/CWfrpbcvooX5zv1LS0mHrx8567Y5FKpO4WLcGPHvrzzbIEt2SZ1HDg4q
tS0SUJSdQebYHzktJoVGb/Qd9AoDlorqylvaf73RNUOZqx9BQAPF944hwFuSTndB
PqhNOqmg/xMBNaxxOu2El+vfDzxEDuyFM2T2ddSqu6CKqs90F67WPFkxVcOn0aIz
QZPe3z7+XVm5bYeE/UbojXezPJvk6/mQf/d7GgXApws5wLO1hhrS/yLYT5Lkq1po
6Yzj6mZ1EsOlrAYiugWrQq9/aygYnocGfXRiAQ8vB6aP/K3GbF4UD+mcjgaYpTga
zknouGHjTIZpOshfJ8d1oiXj1PTm6TSRf3mZt6TOBM4Abjto30IUU2PgMs0oKjiE
sdISkxzQ3r4XYqKH6nQLxcuf9xdme5fw2Htkvzqsi9ffacKYkLOXq/UNSrt+dXJd
aaCDPuAN3+bzoF1N2ZzfL7dNWPtjNl1INZWxhnAbdJbTc3GtQSo/ksRzR7AVLyFG
iF7sZ+VGAhPz8C/Gh/SjOH3ZGRODAUw/ul8vCRv5J1GOjsf4YYyTg4+qm+BY73mV
V7sj5HIRi29T8+ssKKdtQkby1pyRxg4JXE3neLazIWJNKiKcu90w0dyrwl9790uV
PQm0JtpmRwqE7jPUCTE7+Qfr3suRyeHL6NVz3C73JOtzCmc95zl1a8cqJKWjttAn
KVJb25CO2LVdAwFyMYbTmgDPxnfN/4pJ2kNakfZiBIE659GDMnBcf+bbmFs3qNzh
uhsd4s7TDPc6bju17rZMm3VTw1/z282nvlayhGnuLu2Y6UypuP9PQirnJ1rAO139
DpjiRWyVeDKM37CewlzCxdYFJuyca5PWTuGpTmkI842dFcQEVKYle/2K1sI7BcE6
V1dlNcRGcTbVWC8YcfhaxG+Bgsn8qrHmJBe1s7t5LisEpOR3xO28VzCiGBniTZ7A
8ku8fOHViEZiNj/r2LvlxSH8w4orXV89BJsDK+olT0USwXMbfpkyiHaKkjC/oaEr
a7holZ1N8AganGmG62tr+WFQYwGCfM1XFk686LGQjdbb4LRdjA24mT7y9Z6cl173
EwOS5z352lNfZNY97FUhrZM9PqduBzrN+DHqWe8hsbrNORANFBuWYlhAPk4a19Ym
aacUU/FVsGlw8gTRCpspJ3NBWTyDpW6wjoKj2Ntk4j88OvbIDBfcmX6BlaFQmJNC
BCoL4dqBl8cntJJv5Y9e8ImEa+MErQv2yOcgJJyLhsnTNSzXRmtqkC5qMmiUPUfO
leP9H6IwPCmnzyyU2/QfjZpjVe+CrcIpMFldCatNlLCOxiNja3SJPBFmQUGgBWID
BmlBT3vVlwl2Hc45ubaR+CiRJ/XDpca3+fkktQ8u6p0TD99iKp/E0EratK2GCKOy
fshDEFeow6OBud7A7DuDGJWvI5QZrh7Ceysw1fahc+pC/g4e4LrfOzkOhigK7Ha0
j4AzIhAyevN2v6DK0uLubT2hJy6Jv9xG5+p++dPK3oUHicoPkOG2hSu7SECzR6aY
+b6hiTvs6ZugAu4Y0fiAeeyVHVKXBH6cVBGUds1dEW7WpOq3FRIkg8sMVfI9uKAp
HI5LaTo832UuBpfWtgUggHpytm5tdtPwRzM54mizZS0lHXJWyuerPqJmlx5HqMHT
FCDHwfdZ76+LCEKfkN/qc4j40A+owc1NSRW1tr/iVKwmNqcvlqLHNSfKu+5P6TVw
pX8ckQI0j1Ne4pYlhS9OVpeFNNYnbV9m2R+0p4yZANFB6f9XzZme57PvpU6XOtIT
S7/igbqAgkDjgu2moUi8HbOv8EKZEM5XKXymI17YyJKeDBIk0X8ERY33XP0wKT9b
2D7WJT4wAqDaZPd+haNv1C7igywDsbBZTghrbbgMdoLWvxRtGznQeZztpwmrKBvF
HlWeZH2GM1Sj+C8z5tPJIA==
`protect END_PROTECTED
