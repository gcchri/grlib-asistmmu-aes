`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FfN8ir8QwkIAWcRh+knKQKY3g+vbA20d0tO8SXZjjIMmq4qDMAi7IxB03dmv6yCn
nJ88sPd8J4MP4g39Jb1LgyTRh4yWJ1SZyt+A0OoEURj0GdrMTLsyr1WkhPnrL6Mw
8dGQw3+aer/xvsSpegL1duxiXn3fhXyHe5YqHpr2aWtvPSSCVC0ztbtbJlduFovT
coYyR8tl6ka2pzP8ko7ImGzb1RrIa5qkDdKLKlEsOiC80fiW03/mk4xiLdOfaiy0
mCQrX67WjDtMJLRwAmKmzKg1liGJppbyCK/BmcrPFdfOpDXtAR8Xq2eeylHrGChq
3irJPvpTgZs7xNxjNbU8Ds6GYLB0Y0ZyLCeGnXfWeMODjc+DR+0kVZVbzyAD4IKp
v8uD22Nl8ijHR9mg1QXEmIWDnB2E0f6DPuvpLF9m+srIAsm6TOV/VLVHUbIH5Ws1
Gmz1EviRBIQs8bZJaxnn7cC1MTqMBCj5thuo7IMYMs4EAkv6VylVFZJHtgjPS1BU
wMKW2v4wBRo9kavWLZMDVTuyLR+EBGt27Yir69ah2cz1ZGyZAs/Zqlnno89HX84O
5Z5imSsx5/AP/Pb0z3o64454Fb5xfSfslHlc/WjKEvY=
`protect END_PROTECTED
