`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bZnjwMN2pziFlsId8jZwU/Sfmac/jy9JbyVZSMd8sxqbC+2uZZxXkkZ2jAT0qI9u
Bi+jti0+tLtbkXg4Mle8BSgXS6rdGg0oKI83+HpqEDyfN4DEV+hArS0qNbb5aZlZ
H4xMcBXfBFA7/gyyWls8M/dbSB6fZdPvLLuGd3WNVAEmm+6S2ueKQCIH7tby+zLh
0hGfmZ17b0VvgfUHbSaFFO4bXzf9SN6IWBmbr/CGYQnkFeL/3bVjmU8dWkXdlv0K
qixBtH519n61v7LeXN2avSGdOfvX7/F+ULUMUkyXDnN8n9EGt4zbMSsq0e7AuqXR
ZFCMGk8BdIs8nHvj1M3+v68ODHfYZwRhz42slqwczDed1IpIy4/ePQops50D2nVK
alCYZrGi+sadtvMaHlP5aBfiBi4sc4yKKm6DxxEIBmyaUPETsWWIlM8a1LwcwBvD
56DTuFYPKc2n621UrMVCKZ6S6EKpncneK8uv7zbUYxM3n4UEQPQa0ibKAaybGRDH
AvsQsqGas68KgROH5gjg+5COfxoZ4Iu1weI5pAizbqewO4jm6/hhn/IZCr8YBVQ6
`protect END_PROTECTED
