`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hu0b4KVQKI8bqOaZY42kkLWYwO0F6yfB0kYfF4H8QJVUcHEA6HHWtfZkgl0i0aO2
zQFKsDWmUUty5AYyynAPWvsHZTzZ39AqgJ7mfYFdsOwodF8O/ckvTMlAOBhg9i9B
A5u2teDFtaiWafWUYyrxQD3g/AZNpDVfo5MNqcIOd+PK2HyIjmrRYK8Y+kC1MhRE
jlL58lt+uwscRZQg54f72EXTaPnIW1SQxnm31p6mrSm/6G7kjs1J7MJQ+sT4RFpF
YhQ11UwBlqzzmGXuLYZ4Xy3pYBfBRnzt5dYjnZJWUT9pNinJbbLPEKp9ULX4nqmA
EX4Y0efe6ngM7zWjn1tP5xDESoTi5fwufEvC8UsYb2SLbBFn5cgdRolEBvuozxx0
vAK/NmHHLpO8Ux1oo5GJqOE9Z8V4RFVM+/6tBHdhNhMWU4a3vAv7ee19UypsxfeC
hlhH7/5TpAXmOvsBi+Xh4ove1QUU8RDrccoC5aHlUVt9u3rToHF7B0zy+jkBH7oD
eb5DOM4g6aU2HvX515dsb22Yrl0Pgp4slV7FoMSqgOpVNTbgxIMHeyoIzm0Eu4Ke
7hc83Az8ISVc1XHjO1DCrpkVuQUzC8UPcYMgIamtJSnWkwlpP7MRT4JZ/4OQtQb/
u7zfkzCZotxswfH4PWSVaZVN0p70xjKR51fZALmpcKoJyU6OxGdq84TE8v0Icv38
spCAqiHngdXMBOh4bfBrA5R47if9GSFvCIRQ5TM9PX4ImqwxMwizFd/X3kxjynI7
qp7CzKRF3DncJojkU7FWJQUtKcWnPH5SjFsaAwxl3WYlJ2Lmg3OUk+rH4wSfBGaW
VvYczZ/2bzrfeI2SWHD/gGZnsgNMsz1OfUbVm9M1l28MqZ/aj9QB0/NOnyUwIYIP
99dgLiX8NdDP5k7IHG6dyIwF49TwooP4qvZMZ3LYwBcC5YjfSZIlzGxuq1UTnbQJ
Ucf27D2DseCKVi6gp37gq9LSKm+FMRkTtRoFb1LfphGss3aFNq8ohTELEWC/THdf
/1b/2PEuJXrqXrzJQYME/Q==
`protect END_PROTECTED
