`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J+UqDlL/Br1q1HwU/sji7RvQVqfvsMn9yS+1XoUsTNey7PdtUpsjgWB3NKWEAxId
Z3aqyPHsPa/VJ/nBHlpdfTj4AIZeA4bF1yAIjPHTeRoAexlDk94+PV2CqPEReUni
DM7BmL8YLuXlo5BRL8MIOBKwi6ICoCk166RLg/oLJ+3Rh63Lmqyf+ntpraRYl5Lh
p5dq8h44YozhhAXuqM/VXMRHYbaKa3ubTa94mwaUye79PnD4IQr73VOWp+2ENF2I
OXG4Btb+NBRNTuol8uP+y5MUBKD7kAekXRAglLKB0qv0bhSrgImtm1Rqakx7hyX0
LapKvP4QckQkMwuAXJjFzfYGmjbjFd2QDdsvwFNJWUoHw9J2MlrmCd1OCE6u4wus
3zD6cyO+KLp70bxNjPh7zb66vVcMAQhfu7Hl4hEzwEPx0dqqfdmqqbJXJlF4D1SM
5UY+gVHnKCI/W6qnRa09vbl+luwbFIlM88cW6aWQ2v8QPNSq/RF8DBWx8mQ7SN4h
bvEuZ1L3g3YasUmGP70Xl22IfBChjIvuw+QuxWViilwMAqoO+PPzpHyGST4AcP9d
x3biv8lyJMR8xN15XM4Rk+crZ2OdbpAKKaFE5twxn82SYM0XU9Q541iH7ly1FiPe
owXftRlI5ISqwNdLIwCqU9q01xb+d3QbmzENa//qnCuaCwo0J5bCgL3+LleJWzWE
jjm1kBFTe6Qa2BOoxabpUewCho12U2PTt0yv3fnuDoQnitLmXNq+PEi4kH51Co7a
JHpidr7lR93TxuC4hxF3ofTVamUlEZkiOcepLkN5p73GUukQPJguaNcUbz5UBAMo
DtIFunvtBvxEbfJF0UYKnPfEbQmwT3jcRD2rJssR0BB+z1qOX1S3MjbsMt/R2pn1
7dtSgddUoyAPCmRg+dWMsS/3fpdS0lQ8DrQjeB+w2G7pL+jcMf449wAzNfq6Nnkd
aadE76TeHcT/j+KhTmcKY50CxcIYVD4Ij9GO/5HGa/2tZ43QdpCZZgXKaIG8Y/LV
RE+RevEtY2fc7JvgwE/scr5iU9bngGatdT66oBizSPTm0XSjlCWwOD8L3q9tDroc
Lxi3FRk53DiYrzv0Yewtz7MdPNjqeqFLVibJHrcI8j7FEe4wlI6Gr2xvFuVcs+By
F29k0cOLp1mZQ/a0G/zJTgqQqt28UKhQSlgnfXZ7v/gO46Jz/9YNTkoYnScF1tG+
NoSKQlrgkKw1U0HvhHU93lN4qBZaPHhH8Y3zowFz41bzsM1z7UkKm1WUFIGJYyjY
Cij3SjEeVmFnoNNzpK5lbtiJZmzxKu7e+FDQJW4Isi/NN/VgQTe3ul6Zt27OMF3f
xaruyIJKactITmYcC83UcKMsNeCbDRVXLUwqFTGzAoTUJDwq1VBeJMJGwGWONdJR
AnGqRx6GCtRCFwhtm8i851IDQTBGFRx8nqtu+hAcxDErdgqYsKyNefPH2o68NTcp
5FbryrAi0nt1wpJDB0hGovL4/AmNMZUGiyc2+7CAajX/iipZ2sSaa1ipKlPbCKVV
aAo28ZbpTfn8pTWamWIZnenL2v004s15d3c33LnHWCkcIdnPtuQKTNqsIVSIIIpo
i26qlv0dilcnQVP623KmCJnrdLUwinNBGU7Uuf7O41uE7gZEzP+VxVrDPIPRcCGQ
Ux1TKFNBr3bWZgNInhEECX8mQjb3rliZEcQ73Cal7t0AbIfUpMBPYfomYOX8rZXq
sml3iFmLQoP45mmbWvxbp36nYUCv8RTCosQxpgeh53s7FxUGO2q9uj0ug9np7NFU
chaFHmd6TlAZIzV5/CZI5PrOaABZefyFsFiBBPdWcWSyYxvslhQZwcf7vdfCNZS9
qQIWg+QQs8MPe+FrgpoIA3cmwbhdjKXU7FPidzW/8RHm7iXsRaGz3fl1dTtr23u0
J2v7clb/Jz7zGdHJ//brwSaWdCnvI+5IItcBZsezdvoCkedUqXs7+BTp7FpKGs8M
iXe8vULnp9x1ECaBh5WSEEtqrZQPnFEp7KHzu2MeCXxOjfHMBWdlJFqKvuTuR4Jj
0npdm3J4kjuT/8rhksYBAc866ThdPB/NGd3zYWieQm/7vlCuwLKFqeX/JooogNnk
t2L73pDb3gaWhWrsS06pRMXfOS9wY4gycD1pHnOn0lSQp8+qpG81EiQS5K38CEHQ
9AJJG7zDVlU/2IAtViw9/Qu7qOpoJY3GQnsRU0bmLAt46rKK258vx9DQpQVb+Bqr
XVC9XESr5gl0QCfgcnZeyoJ7ZiPTUfSkcVaddvL6gDQwW/zblG8RmUDD0UJWG6Cu
DdV5ZBHoEMF4q0DK0xAmiSDQhTQpECt6Jfy/6T9bqO1un/MihA02pMv9am4ao3pA
wO79l68BJN+6GHfsQLJim4FuldnUg3XqbB10CDcxkcNqSaSPt0IcMrWich2uw3SD
GmeId6JkGr+pfpNuXXML4lIz/x76HB73XpUiv/UKLVvsCwiCrs6Sk6BEVkjhHRnx
EvX8el5WUTBjqyN2CuMf2C6ltOWBAsi61F98QjEvJp3liCBbLgHO0bNwi+Uwe6ZY
dt0n0W8b6Inc18Ee3Y/4LLLtTXvt2PtPVrv7HXPePIdyH/UQ8g5k8o6EC1wMaEJh
ab7Ehs+u5ml0X7jiHRyHDxIgfk69yFhk7Cp7PlTdXqkSEzDcJ3boZb/Bl7mYRjpn
PoDkP3Xblqj/9VYL0/C7Hm+6pZOTtG0vWIQIHHmq0evjS646+v4h+w1Hl92luEJN
vmLDk1pGFkBsZ4Snrh3aZd5M0EOQR5bGkw25jlZrBb3p1kd9K9Pc+U/TtfyjKJ56
aTrxvcsFNGLM3vWWDrGXBamPBjINIBVr2tONwPJC+RoDrsfPemoP+7pJKcQCAfyZ
pPLoTDuP4vkwiSK8AUzCVjMUPg25KCWoI/HTw30UgfwMMevIpQCxVZxliT9iVT7W
lncOjh3kXUNdA9oimsgjpV0GvVcpIwOXiHhVd6r+n8joKdGwY+9xAKh9Rq/I1eIb
dXG9DnFjvItH4bWN70RW3VdjDM5D48P7/NfbNryf+icPL7UI4VTDdwmQk5wujb7H
Rb+tjnEC/2ZnyQKV9Tlg/CIyAGBelwGTlQZ3iI/49D6nfXnzrQ5XZQgRBb1Bvodu
Nh1hJXsL8M2XRutV/ivAjutCUjMm+t4tYAEgw0qQ1QBefTK5wWlaCPPQHc+geKab
8S0DQCaWQuSRcDE4S/CfaOpAKwmuDtH2Bfww+PLMPRRG+Ee5y2IBi6s2CGYbvpE0
+XmaVBYXWR1d0f6oxGiy+7zqU/JAgQHjiX+FHb0uZbGtXJ7JpvAhQYG0o0KfXlwo
fJq5p69MYEFLczAWt/rElnNG92d6yamzLUebfKiWxJseftGlCBqD0nJLmDB0d1mY
WZWpIiVPwmJvLvUJzxVczLBx0K8RGVwkYkkjeBPZMCdrT0IU9d/K81kk+Shpq52Z
JUmdNbBrPSjMD9WvDtQ+z3kxVsIY4H4Z3+DopkNgL05bgGz2WByhHIMQ1FGDuXjx
deKYaW7dZljoZxMfEKyvDAW+rkwAVa/hYDnFaKzGjsfYp9+lJ0R+jZDHMo7YIGkz
Sbz5QujVs5kOv1Aeg9hGrkeKHU+ojrYdmkhOT/2gNnHuOOarPPiJD2OluZWrQHJn
x3FGfUJzXA5hFxX0/1DlXqnPn+eAz9J+aRanSCy9jzhwhhlwEh2+RawD0vXgUF3f
WbAAq5StwhMnhwGB6il2wA8W5XqBMJJ2/lm9rJLKjW1MU1GLOOAauTcSFUWJTIkt
d08wmGRqG62Rei9MR6wzHSrCezrO/0rzawtPYuObcngVUUvxNZ3mrcJXsJ4jw0AV
Lyv3IS/J4t5UabKJnUy70TlyIPEqlWQo41+63eyE3LE32zpYobIk9ah9Dl6Z5Duy
IHajCycLZgC5XS73E0Wld6QTqFVbjBplbfxG1MBWuCIneS8W8RnY2Ufu/8oXc0Jq
zPbB6MNG6pWGkrx0684bYvhRlGTBH73U7FTkgCM607Q/NmqnP/QPbzputB8jDHlE
i4sTuRhKyUGtSQjy1cBdqTmDV93Gupc0OAYsC4E1YQ9vc/QN/gGd/YfCFe1YLCMb
2XrVgPwyTZ1HCafyoFcD46OjcEJNQpHBw619Ot/RaIUN+cteQKJp1fPTHI0sFQmL
ioV896R9DejvW0SCP4Rie+ZWGgsa18oqEYNdrWxI2wILUP890fLPtkDtHOJu0Yus
tCZ9Wk6jV5pG3UG8xxHdh90i3FZ4GXT4adiihmOJqUc6/SEbwnsUZ3jZ+AahmM0y
DKnaA5L0FY3tocc260TxhW/ClII2SgIvG0fbzmi6gvQH86jBgnwodgEkdxW4FLue
m40iW/b3ReJu1fWmBvY+2Y5Sv1t8z3J66X956H2eFfEP60t/AZ0hqX0+SB4VNyKg
yA31+ZITiV/ojLyoGyOUybUrzIOenryGU54O9WaCWwI6JKDxiaVT+pVceKeqgihh
F0GRIaZoArhZBWle1K9sly9hlRLHQeKFxH5tcMMZZRlMW0aXRGhXD+ysnyYvq7e9
/GJNkhtc39x+h0z8zGwD+XFJXXF40FpxaYpCnGQJriUM0iGyzqKXPpGkhzePlCvn
Z6ahkNOejt8AesFyoEy/mJyx56xJFRhvZVvtOp9L4lVPxA2Fjtapk5XoWp4vN3oX
ZpgyskPuJvdEr9J0QdZ8C8JubFDKC+LXlBGCnWSGEbrt+/kUdSetK87DP/Lil+LS
xRS10/qHU14HctGXhBHhyjyIdYvf8511XA7Cmy2tvNmBcbOT8M9I4Qw0GbZqZEhI
7eKFQuGLLRrtksYY+u/+xAAypTouQno18o90YDtZFn7yAuMgLTRBNE7R4DkLKMzc
zuz3p6YmlmVKqf9X7ECnW4c17/EX2pQhdRLdhaNikAJxhHKZoM8YHabvsEXVZgvt
7gOPKxX/L6jRh8A+7ecskWABVb46Y10ZPqVrEACFhkqG57C6EVppwl0gTNsnEKo6
AUfv4X9sxsuvQAhB0xY5x2QebKsTt/J61KKT8y+qslr5o/+ARuqn27rh7sE90zMt
EIz5LniuG8yEh/lzQkDQbbnhOo6tFz/LYmktoHIPcz92DBLlNqmm2h0k17hi2lHs
4nNdGKI0wn5kHxOhZibAi3F0coIR/702X0yoS7fHojK8hPBPkriq6ODPaUIWg+EW
kB53dRmiS+VrIRwbSa8sSPMO8L7IQqjmVFhooU0Nqtps4+u62raQg9ERj+imM5RN
n+gerH6SkYcKDtwx5I3TH2updvbBFbKgyw1i9DwUTD2C5c1Eo3Ecq2eBN4yNbHAi
a6lIVNJzXyJr/5UxvT5EFtSDvEhq0+JlOg7xyP3hdCowb8cTZyyRp/XYF1qtHLGH
UB9hkhMeRPM0ro31d4mlAwBBDVSshEBTP5XQE6OFZ8Mn6+Ln+htJCZ7NDO3+YEq7
wyOEcQDSMM6hGDQIEWYOyMo36NScNJs5Udm0Ipsg9SN2Le0yQ3vgnLXVlLKh1QLI
r/AVpJCXHK46ye5mWFjJpvDHRvOj9x2f7NUmZItO824PQdx1ChFqm56cy1mwnZLO
O1OLx77vEQmw6azOAO2MBAJZ98B3GQLNLtZpSA/mED1lTymq0PXaM9U5B+wc+ZWC
qkhvhudEKqqkYcARzM2y2Zwwpkj1KQkmmQ6/FMQDgYrV2QzOq62RdZx/04KE8YO2
HZtxgVgHchbSnnHJtlCQr5wDzBNMoI1hzm76lI+UE18ZSBYi3oPE6l87fc+SRlfA
Ci6SJWhJwRjbNYF2cRavwcUvEOG1hZSHcbyJrEqjr1DKKSXM5pGjL21/qT7272jD
V47wsuU9xZMB2PZvIQudWQWDjjg3HR0TsG5F0+BbZFdbVDt4a7Wdktg9wutOlVhk
Rtnfgj51y1iDZsQ9SizTdqji9TPgUgIDmq9Oy9PXO+RnX6Bz2WQF3q+zNpzfXmUW
nFfQ1oue7VBdsdnNqiZQuQl9UwEKsPDXNC5MyJlY8zIKnWjdX9ittquY0l9+0k2w
oRygKM7s/VQc+aot1KUbxv7BpS2RBFwOEcslKS3SMd4F/GJrvqsbSuzuc71ZdudU
8xjgY8G51TNgdym/XHpNI3BU/mETXJ7ZY2fjG8vZossmNZAY29FhpldCU75IbHmv
aUqGeR4b61tmMV1QX9n6MRX9IrknxL1rrB/zfRpbAh7T2+cEvsIM3+929EIFDUSa
apU0Gs+DHA/BsN9UYhfvMruXtQWXGny83m96Wbpk09L0vIV+P5ayyvGSDkwfLYlX
E0mVfVbveF4IAh484BQ/1AJKsPHJpu9uvlMfUhcq2rCg06bARrx9RvvCnw5vF6ED
BBPdTPAbne1QSqcwat+vkAQjW3vs0S9YsP2z+0oRjZ6U64ShwAnxocQ9si6MXdHP
Ju4SNLr2WQ7PF2xlJPqHeJYqskY21FOraU5Kk1+gHJx0pjUeiH9jKSCTFAZQyWMO
CMStbceS7HKFr+Trwv4zZ65qNzHaoiM3EMtpJBqCcGrw8CH8AMTlwdm74XHe4jLV
KlzBA4cQn0LZQUYFSbggx6uqCEsiRuS5EeCBirzWHfmBc1F721RJCzFAckft+DcL
DoEkh3LCwF1Lo+seIA3wjcKZ8aCyy1XagwXV1jQd3OnJvyL4qTaTzf9vMabkJkt9
wEe8ubHFi77fiXILcbNutiM7UcTABhaim68l5SCsE4TOCc1f4M1AZjP2AXBGcMth
/EKbDHJtvbtFSLsJdFn+okc1C17faBSRAekyNeumAIe1c4vtjqPH7SIypqlXFl4g
/Xs/NGI/oUgKvJcx3WldEjmGi4l0QE5vVbwKKxPDH0e9IfEG4w+kHjsEPki4CG/o
ORLoP69xTOZ8xsMmuDsiQ0qcHk2DqG/ycPQjYr4wRlSwI46JWddxM0YlaT//z3cu
vISSITwqI7nZde7yihvoF4XrN4SfO8aQDGj2aLVv43YSng7G8E2aF9qTUcSceHfh
eAbRslItyMfh1pRGSXzLsnO7JiWFRVO65QXYtstR+DN92WY4pp+J7Q2k7y/VZmVF
g5EU8yd2r4TADcWDjgu6flllKzTRkqfS2BtFr7B77ni1UFzixOvhn4JPdszDheny
Did3/ZKpCUKoBA0j96J1CWHFQ63djMzze5lbnZvExzI21dqGVPNWTQo69qKtDw/Y
HVgwJlcBWGT51JXSLLwsqTIu4hQfXVP3FRT52ZZ/d0UpRsvhuTi/zo4KVAohvq6u
ReZ4Rh4y3VNgGRhRkKm18iERiuvPd8hafBxGpuCuE7bcwCCmpfrocN/JWeKdLPUP
GdOW0PwhwOYVxtlbfGdy7HHYg2En7xibRVUTSZsx7cE=
`protect END_PROTECTED
