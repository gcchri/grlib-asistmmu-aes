`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
adwxGXnRNSM/mhnwk1pFUhLDauwNvkSgQ63wp2UVpwpPJVe/xOZ0eCvVRt/d9wE3
npNLtrVWXPgZLYrt1Ay3unibj+NE+m7QFWRi6SOBoWXeXMbCbrAawiRB/efoLNZl
ieTdRS92CyW4/WtfaoYtlCmbMog7OgvnVqPovYUvn+8G/ik3XVXlI2acPx/a3Hlb
Seqt3sF8Ndy3C4gkPqVFWIlXrOqNSx3pvObW4MDezkv2NRDllQuMojwpBqrURUxE
Oo1cW6u5zsO4lfXdUElNBRQ+Od1gmOQqepo3+KFNh+eLlomx4J4v8d5bxeRgEL7h
nHyHIR0zDzHKezEghls1sQ==
`protect END_PROTECTED
