`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CPcVqUw6i+IIimXZUEVWh8FPr737HTBNECd+5YsCaPurAveQq28o3wcqPhpKf4EU
tFTl1w5EU5gMdhhB8ifRl7t62It1Q2TScfU6aR0u/aTpgC9Vk5EOyGfK8+WVSDFK
mCYfUFU6/+qMafxHVg/2Y3H0vyEbobWng6yQUmgmViv2VHyBKZLcrHuV31SozUkS
NT9mrEnvtzi5/90aY/vUUpPS3RuPNUQdOsY114SvhJiSlvFAs9kXK4U2yptjUtmW
6pXSvdz5w2TQuJbacxEKEpRv4bOn3/GPldSXmZXeM8UTwnoeXutSuoSTOf/N8az0
CdLnvGM+CCRDkACe70KT/5PGWTfv9mvkOO0493w/1sthRUabobNqhzV38IpNIwMN
qkpO1cy2agJymCODzi/4nDdjvQ/NFwZXeNabpkmRxd8yHfP73RqRANhGAEyQE1m/
fu7d+mkHmKq8is4LzUZo+4zRQPyrrtRFuwYKGRQlRzRRN0oLCejgNPW5jsynnC+E
wNgPJsvHXdyHrTr/a7neTF88wKgjwMEOe38xy+Ps7qj+sNRRHpa5BzjN7ht6pqOt
wf/XYxpRY38qlYk70bdTk17CpkPvAu+xA/L7ne/h2rq8xLdeKrrV+IE9ynizJDYz
G6TeNLNbm4pQPdq1kEPuKUiLWVqtFwq/Xe6w+39rpZ5ZiDf5IxbMigx1WVy3H8Z3
+pVbv6jnfFATovXD5toldQwWbezMJ0hHuWU7FrtpU7BsIDO66cjEsOnFiRVBPNdU
+eCB6eI3Bj/w4LJeUcensyAR45aV9lTw/zkVVyu1uoVSJpV6Mqsp500GhXhBqLH5
f4Pnd9TBXRKXoTNPnGVanxDA9W0iyIKcSYXgq/3WTIW/lRCnWgZNNqrnSUZB+JMq
vB3ZFjuSEED50HXVLcst/jGhvrtBIYoUfOjt/M++zSfhzJCRnE8F/VPstwiRbG1h
4j+t6/5LIXzCw3gG31VgPgufkMxg2NVZopDdLI1at05231fyn547oG6SoiisOiwj
thza1mJTWX7wLri5YtvoO1AndYoML0pvFSOh+yLQ/wJX74ycS4kSV1/j++nlegB9
pd6lRyVcpp3L4Mm6AW0MkcD0ItDMYsy5zMzqACf83afOPVo0+gvEGxN/JJLyojx4
Pr8jWWOKCkEY/klsPHT/IpCzS0+h3YdmlhZOV5msNUYktXhvq1+Mwxx96JE+oT1l
c5hVvsUai9I3K07BJ+JTGT24RQB9rEVVfUDKfAicYmyCt6V/6igNAnTDdb0krsHx
vN4hljDu/nLwjPG6BTjftyzFmxQzerlJpiBORknhq4AsqIijErcq8VT/CZwhOQso
0V9wyKWt9FTpLKYRJ/9VS/D9cN3F0cPtJatPUvKvxYVZr4V56MSdLeVy8W1Vc9Ra
YQw3riAVU8pr/odRCnv1qiQaTycNymMGWFWCVOI3Q6aswZ1+0XyuaycADhXYE89/
XAymLF5MicLM1YwXd8gajhXtHWuS3rylpmTEumWHrr/xzy8+9wY1jaZ4idmO66tN
eNezacxL2BQgK6RB95ovNqtNOuMPyf8aJbXvpfFX19o=
`protect END_PROTECTED
