`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K3stgqGDUZd7QT729VHLeUkVLUkCDt0ilBBxrZKNV3g1Q+MSqdfJ8+mIAk6yjMJf
W/PhIQfKGWbKHLhzjy9zaEb128II7bHow7avnqLOmmg4Am02r9Pz3Fn5+8uSzE43
j+S5VgBsCnqv/hEJ66zg6zGRS6s503hE49oGH25dI7ZJutt4dCMUCv6Ln5dSKlC4
7NwFncHEibMPAVJ/Fy5D/TQSrSQXxGhN30gSPC52D6alSeZDAY3GMyIGNq0gtjTV
hiJnzD+ZzjUxS8Z0undPZMFn1EKnULW49Haq8bQrEr9/RmYNH9vZNOPGBwGnFPWw
IMgfcMwvwCKiC90WfrJ4F+XvRHRxfSsEwlmDkF8+LfGHUcmBwOL/CCFTd3G0p4mo
oHIFyPV5lNNYMCSp4tmSfCwz2b3wpf+2r5bXXVQe6NUiQSi6hJonqda77mTR3Nkh
WdksBb8py31Ckf+r6y6rJ9tGuDGeSJneHvIeQW8Y5lLz2AE+HBn1MUP1MOaOsA/W
RMTEyCXaLO+JzOrY6hMAXGRAUQBIQjhzixze2oP9B9TEz1PD58LXz7XoKf9kU6IX
VTlioMEwFxR02WkEmCqkEKcKUrC5x1nzYPzUKxESQdnjzyK498T6FKtvDPLKo9FC
fF61PRx37w311aGmFnwImBlFwWxjlkELyIqS7ZxBInEK+QoaBWBBGUz8LOmOXHiI
jcR6zfWUqdRG3nJ22rrb3iSEdqhY8Ddsk5+4YplzJJhy+Ow9W8ElAfrS3FsZv4Ny
v12G15KLNIDyjKSNTOmFWArV2eoTDEnaZixekWWXZijNm7A4pjFegew8O4Avu3Wq
9cmB4ah2NhJH5QvknH3AWHOh2p/DNemdiw+F1pTz/XsXpjmbvbyj+sbIed2bXGbK
Uhgw0t37sF01bcGtU1F3r93NJiYYZbP7k26cdO036hhm1iuiIZmARolYn/vayYHG
`protect END_PROTECTED
