`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jZogxqJdtylEAwuFmO5hAburmTKO1a61Uvjb7L1gz0YqtbFW2UG7JtHjWuO7hr6v
71jYg8FnkKEXL/NRxE2AEOO8W1NqsXQfpb5SM5ZjqrAvepGv3iYNzsaRKOzlXgB/
wXWEjbbXu2AuH/lPGy4rAvX5/jUkpkJiEjM6nXZJRDLtXnrhyACzVGKDjCX6L1+J
5abBLFCJ9nj3vwodEszhYJiIUC4x5UU4OmYRLG0IedlIqiPGEZhv7H/s+222EkWY
WM3n94Gj3HZ403g8ZAKdrigX74OqXIVA4W3SOUXo8pOgw8eC1vBjRrlAqi+nize5
BzUCv8EWg6J2kAtYfI/TvAmvYoBiky4T2Gg+8z+TzWntey9w1nXTGjimRVt+uZtn
/pogfOPtZ08Dxa8025M/a+uDZgfH9VmndQB7J7Uz9ufLKedJsTtuzjs0p2xKodEI
Mez1CPMIu6PAgne2XhUUw0h/PYAt5KwJz/x2cGgi5S6FwKqHF5PkyD9KBi4/38R6
Goj5bX0YUU7S7zdSidtO/4b1jtXOq63BPO1DiOUYjVXJHCyDyG8SNPkWvkN/nzY2
uwUY7X4GXvM+DA5R2YRqKrXWPVTGb1fVDoUCf/0NDfA40XEsqglFPb7WuZL3jd5t
XUxuHGIZj0dy8w/Y3kU6ypEZFlKtzAIJ4wG8CMRMB/JqhCT/BTxtDMbTlgu0PPR9
cNqzKjeCt5YI4nQsanv8swsbTQZ6KU2MyKJ+Gd/ktcb+pbV5Gv5iPnuk4lV6x4Fi
jt/RmldKt0v9hN+9AQhchkuao6n++dpwpuDYIwBf7t2fqucmKGVT5nt55KsNFnH3
mvfChrHA2+T2/+7+v9hRXqojH/A0sTfILrKb9BMqYRkRa7udYJJHvap79gxkT4Lu
`protect END_PROTECTED
