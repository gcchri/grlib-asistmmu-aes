`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C5fze7xI0SrXQSk37zo8MKKyB1xdbjw9g/yxw0VTFJHBWQHHULAbYTehvT1ns4kx
lQZn+izY+y6IsXxDyfdVQ7q0rFcQs5DyHvuh768NCBnMMUM7pA70e5zM2fWI02RO
9QBA1pPI/mVOpVKk6FtA4KE7alhg4a7bWD4UHgOXzgRSeQsDvhhXiBk+pks6N841
ulsJyqYLahtL3pPaAQYVxyjn6qsKVyriCapFabC8FU6jE23zBLDzDbVuMt6e7JDF
8gyXMto8awyI3qwxN2pbcL0uPLj46hUh9hnYVNBkW+2xX22DXkD7MfFPzaeq81RE
UiIYiKjd8TSm+/9JkemdYpWtgl8ojxiH/0aC+J2H92M0bvvGhfkQdG+iDgvNf1cN
a+PuIGOuWnXymlHbldwJfqOcvMB8ZluMXNfxi8lwHdAspIhswBmUJlOq7z3I9zlQ
YnmmffIN+qq7uyOizXbcvVEtz/RhsPT/gNVCUNmNb/63j6aY6lLo1LlP0O/ukBfg
CxDlEEldluSovUBxV9qO1hxRIzbC5slnzCA+zia2kYqR6XmmY8F1Px4sGvdm9neu
M6VH08Jk01Q9NWp2SEgZsD34/Ant2MJBoSvl8UppSyl8jYv+C1OT4sOWSRHeYNj3
cxefQJF+D7sE2CHSwqUqQcVuh5pfg+NmBoBr6h73Ez1U4RZpph49ViowvbJwhERd
vFW6XsxHBpJZlmpnHHN3VFmvqd01tlZJ/UHYyUBMCbmr+P7keIF5/lnezhqFlhS9
A77hiuYPYgFf5j1x3H7BKRELPq408GT0Oqe/48AOqA6Y/a93/gMIA7FDyWpc6Smz
6kwlay2lKuqKF6ixOj4sKpsqkGrYRAy6pX9j9Ov2jnuUJhw0KcEme0G13AF3Jzhd
hn97UI6GX0I9/DGe5aVTdezo+bMWAYu1JbGEA8E+DP5HGCXYJhN9EtbP8wGAo8Qc
sc9oqsWh8JJvOhKfZgrS7QXglMZGH6L4+ax19E8Ii2bOeQHNyZ/SGQfMTzp+nmhw
dFdn4dv+ZUmt5XsrgL1TTDHl6GhHTaPuH5HoFA3y0dpz7GyKYfqFq+KvSV5Xg4c7
mkY1EwG1p/zOzPgMk1YUEI8Z7sFOx9caQO5k9E9JpTCLkF/dpr0SwCB4on5ZxgFh
szqeiB2XejmG8i4iu5eHdbIZYkSvDTZLX/AEyofZmUzqkn2M28AGzKGcO13kEj1T
HAOT+guqouWCV8nT3G1YzKNx1lNeYzSfii7LK/tYjTzHIWc5HsAt2Ir5tvGylrEX
dHj/mmal4TYC5jXIYwTWSkXRvFeXJ4lX+pZs1jCYDtaO1AJoqg75f//u9t9sdk84
mhHixT82wrRzr9jTtxVflr1yPgvthKM+JKLFem6jxrPhOuzCTmnqlK/pmhK5hT8m
jmRIjxWrQgwaSrK8dwobZdTsBEGVe2b4AbFV7fnmn0yqn7xv5QSnjXvOTOz565KA
S/fpt9qmjxJf74BKWY/N25bRoO/MK35vjyOaCJ21q90kK3j58RF6jp5S/AFm6VoL
ac0vOeBqum7yvrsVTSNq/32SmdmYgYaWXCFO6Sfso3wVPOep4WjypIbBXH1V1w1K
CcHY99bn4a8u8aa0wqPk/4jifrJuMbX7H2hNOt9SxlUwpWUJ9boYNqQJ6RLt+Poh
RgvNzqwkpaGyQe8DFDqzB9A1LpZKQizwDhyJDCqv1HFXD3+ueh1A3E2fuPO3KMcW
cBy0foSuOqcED2iAu8U9CV7MpDUz2nZq8fbv1Zc7L/Td+l+x/R4+Ti2WGQ4quSD+
UfzFi3Zd4BFHUgKr5+nH50eZvKi6FgtADVPPl60QM0N4WGafPZhq2kxqsYR+mevM
5LS2yKZ5ArE79AresQP5lO7kl9Mv5ZbxRnJu8lCEEOMT/7TyyqoK1a3DgUPvekOO
o/D2zy8fYDN2Pd0BjkSjVpAgO8fH8OQ27nmzDHP55aFXtOE7uBBE1A6C80wnN0+b
eN15+o5CedDx0euCLpnBUeSFuRQkd2M/HFdSm3xjPYy4xrzJoolAdGCheR+QB3D/
WY6AqlGtKX4XmfGQhT3cpLr89U7EFW1dFG0evqKCHJAgRop0RFx40b9YOjxOSyvB
y2d7KJyiDZTPs5Suyp6P5qQ1uqKw75Z7NHqVXMpSqlfr/4Ngm0HJI3AQfCNTFa1G
RMlIsq7KtM2/ZHAu1F/hDuODegL2M/gwt01+BG7yL71mt9cfSFsJCjntNYV30UsB
zf8X+n0wg+irtogojlzzpONpGkmMKP7k3f4E1I5fCS6vA+kn/3tdF51D5bKxBp8w
CvDo/wBUWVOtdLAR+qsqcDYMqHME1FCIkEBYfcHn9CcvvfAu0m+4Iv3/jjkI4it+
Y1k1ca9IEd2ntC0+LNxXVZ7iJP+6ML3//HofKjShM1qCVYXs+emKIpFbB3FwCzEz
FTxKoARvc3HxcBQay0mEsouaUHTzfBJ0yz4BB5+04hEk3/1l7/roqKL1yVqeCGHH
tWubZ4wvkloGe1kEKXkXRHW7RcknvjVWb6I7OeWfZDd0laORpR1GGLEA/J0PGYCI
EaNZfAV8N9+gLB/+c1qTrk6tSdt9o+jsz7ZtOyMTbqeX7ozunGMcy01AcPfuHWzJ
xai1ND2BwwtiZ3LZBI0kr+vzw+m4ukLW22Zkf6FanZr+SUrDHxH6NdVfAA0L1QKT
RSzxOu5lJWeI2ZQlOHM5TIVsN9Yex9lf18XrOjfHKBLqfzBuBP2uxtO8tQaVythC
tEnYONLS/PIS+tkHyihe0f9Ob/pPBAh2hgoz5bWFDrD8ssoNijYU6T2qVQkePCwp
n7ZnF8gVyxel8fF8Xn3ucMXtAZb07iCEJY+yGf41FL4R1LULRvvXzpYaBknw/M9l
ajpolCbhRLnkgSzW5QKTYRKSzoDAVc5iPI9gh+7JUrBEggFcEngPkonZaQzwDgXp
6Ec8ggMPpBcaYE8opdyyIJ4yQYgqmisYqhQf7y4noaSxy9N8I0lyjGC49AYihrIS
GvbDDzp2YwqY6SV0MEXWjwZ2/CP/JtXn+0mVYP8LyvBc6cFbOx4OnPTUeMUI+Oqt
TQ0ro8rr0Msk+iA84Xe8NiDS6Tm2vTy6WTj6UWBTj1uCwQ+a44RCOiLJjPNAgwfd
6rgITg3VWS/6F6bN9vwS2aSTf+xePoIBxRp5iCnbp9CY0X8ehpAQUwT1xij4E7Sn
SZHjnh3L+BOw8bRRySO24evv527Jfah9/uI5wiNP6BgnfpYl7FtGeMnf+/VbE+OF
Qf8wsVb/PADGwE1KBTyj3Ys6oOXX1VmBTHGOGLDBffuJRRifELXLzwChPvCmIPFV
XWIxj750YstlvM+Im++GA4MpuUWWLZ1OlFrVQHdP7jYNVRF+UU3iS/uj2C7z5nG4
3rdhpRyGmiaa6I21/HF3VymFn+qn7MJInzSLNby2rVO4Pl6dbdO2F5MI4yLsA8pq
p/IpmEyalU4ErTGVlLmyVK/8Zr0yW/HN+9d3+U2IgKAlpVK1XlF5+Cg8oKjXLfpK
zTC21IKCiwLSFiErVQBBxeIms4xcRO86r/zwGMn6ciCQJN94VIHtYlrR+70KmoXu
jx8EnwHXlY78RhvkIEt6+1XaSoc+s1YoHnTyiUfbyjPZ9ADPFSNQRmXei8QE/OKb
AOj49FBM8xPHup0v1MX15NfF4xoyd2Hn7BND5CPZwRwbOJUvS22w/KzynwvOX4ge
ORLYdiuWL9xh9RKi5s53ID8h8Qk2NP5TDIbHjFfiRa9F8A9RZt8syKGSTV9rGDAG
3kF5a86jH7f/SenvvtD663reShMp5LFmoYatogsGemYn/3ZgfOS9z6HlwSQN2an7
QwcL+hM112yqXcTsBf7a16jtkHNCxOpU0lzW3oBHkwA1aNiZ+dgB5hPOzb4dtq2R
JRTTskqsTtcDoSP+HIfwDIO/pXUwwB2xlQtw4jJ7AbmqfRDxLZBH7QQ8/02B2KEc
RsncC2wxtVd24X+PtE40/DvuDAul4vnSJy6+X+yU8HNKLOYzdGcwBth80TodOkb2
bXtiMmJmfgeSENsRRduS7ZLwpVbjGYVJzphIRWXvHhjVbe/6U5VIOibyK7Z/eJTK
tR0RZAqA1FINZjQGhlnCG8ppNqbdBVqWYkQg5wglfASlOzC8qr3xtwkITQWWoIGQ
3Rx99epAEvdTTcEvUl0/pl3C699AfzFOX8NZNj27eXkI+qzm/X0fxNPTb4pWa2dd
Mw0N8CdMXY5artZX5PTvY7aDMr3ecYnuinyRGsdx7/5A41yvD+k+Sq4ZFRu6VvA5
AplexIrmIbvC/r9Fi0SWRWi2a3pYPOs5xSCHCAwsViADkaPKk3wYozVuxvZ/HgoT
qquic7nNTjAv7zQG615E5GACUZne2zduP18c5WCC58+5m2oeK9RCcNjdq6cS7RS6
4RgN+St+xCs7IY0ZSYyCpRv514pqP3/VNofUTlzmJ2FiGQbl4nLbOjzdgGBGuCrJ
SSe9x7KnrlJJSxIRaVmkIz6O8EGOe0hQBwe1uGkFpDlvGOaS5KJL1UCVDEe9RExV
1vR5JkrR91mhVGp9t0rNCeII11ra6x59HqP+0Neo3ZsGTYuFx88C1RRSdw3YgQ75
qdXjOv9IDKb/A4aeva8ug+hZCzwTjFxUpRc/atInDV/Iq4osXJ18gCxS7sYSOkUt
EonOPQCHs/lKYXQz++bL4SkVGsGbqiJJsQxnDT4wCUEC3a9bZhrMUFV4vrTFMLdh
fzH92A5bvy1IKKYV0ItcF/w6DSBJimFLGZHEnshlvAsbAjF9g8N59l9qlFHmPVo0
i8fMo+vb4mN9d6/Wtprhn72fV3lpBYQw/c4daBEgyJR/Z+6qM6bgF4PWcAbEAhk7
ivp59qUyJMm6yt6jWUr9sNd/XMglQ5Q25nN/1u/EzIacND+ixindBqMZTzO9TNC+
f3d5eaFO+3i6Ro9Mp2va0HM3WWjU+HVH2jk+gv6E9IeeLbYFxKgNJFpS6INIpW8y
owR6FTMKDJC/cvta6MzO3i0SeEwpwCgwK+lzpQkVpeQBhMWKEuMuGoJbiXjGotZv
PrdUOrSYAP8PdIOET1phRW1F/FDMbQuO1A5wdg+fN98rb+aPggTPIv17YLbLLqlp
uITZpOnkLfEvMvnm5X1CIYPL6tNeh6RSMxP568zAARlhamMXBVBfhG2LD+qjpwEg
agIwU13ZOaT4ZC9W2d4bYULHB2k1Jbh4PrrAgGbHg3Gdekm7pUDANCHm3m5FtJib
wU5Y9NiDH2lc/bB5+oNVjQFh55SE7/WZK4W1ExOz0Xk81KszsySkxCL0iuO2D22z
iMX/eZN4TAtUQIVA2qo5RiGtgFPIoLs0ltnnzdGmIXs44JE3O8X8euWwiV1c7CYp
+AuhIjivY2rFYcPUMaVPEIlkHxdIzl40yLsmD5IKm5GEWXmKWB2v0ISAsQiR4oQ7
cBWSYlVndgTG9HF3OE+HjX9ts3AW6K3gttwKzw/4TvsA1yYN3WDz944T5JqQQYXg
qgBxyy3fxQO2rPpk21uU+arNvjZp2Ycb3x2NU1SrDl56OZa+AV6MmNBWhrKldeDa
UMhP6xLygNdpFRA2iSlAXlvCl3i173GhXze/IPUOZGrGVKpBpez50z5QQQmQrnlx
wcRPx9Uz10xRjLtSQ9bKWjg+iUjx1fcJIh/qFzaxE2wiMM8FwPZosPRUp2lNZ2bg
xoLq5gpxD/gaUYCKRrlVyVkS9Ep1VEhWKPIlORnbU8FLX4IM5gxiMgHZ291GmRhp
hNQsLnv89cGUcSK3Cs60wN5J0tUzMq1ZJIn/7n98ge+6JIkxkh4Skdad7Nzk8VPU
l2DIzumMIu6vH0jR91QuvlOermyZWMo5+NRhBqwK4Z+CRG1BjangpCJMUmvwYJFr
ULYoaI8yChkkGu/l4k57qwvWFRK131lO4MFJ537tbpqIlRCqEBCqQw0Rhyxq3VxV
/G4isS54Kh4L5Qa7TO/SCTrZAxPX7LCQXk5oTf7MxHhxjPnYQNctXN5R+HFim+1J
M761nukJGYECVDolunNj2AyODL1EsJmV0gu4FTkNb4Demi6DB80lw+qr6IA+zGQD
Y9lkODqVIbhErdkCVyOn7le44e3BdLP6ibHCALtVTbZuwzMjPVrg8YwnJVwhPm0I
ijj6aj6t++J+bXO2h5UlYmJV9DOMP8PLs8XpN15ZOjKNKLQZi5zJ+KCsIBvwjndW
4zl8vT2sPAw62vOcnrTohcBu2cgL0CVR5VkfkMXEQadJSK8JvEwubuLbVdevDqLy
4jqgDoPugSrngiNkwifYV2vhXIKLMUka0pH+/Bxp04yuLhbE2cGlwyu4pWS9hz1J
6M1hKD+40BjYls4GEVBIVbGolctpx8vmv3gO4I04PicVGF5dGFaFn+n7TlH3ViLK
R/idfrfWAYdquEqaXEK/avPgO1QspYDXD0zORT1JvqBFlJiei5irc9PjFwA8H5kC
teT6KQFyNqlZhqnJmznySOMwOoVVxIFgX4SFrqPegypwZ3SW/y0O8htEbgsjXQSY
pfPEmxEWEtC0YSqWSX0+rSkKojmnDE1C4MwhvSL4CKg5+akgssLZ6Ug6buGukPDb
v4YEY6ZCk5mjltLnmv0PufYabBJhIohULoW7uDfAhE1irEue04Vp/HJ/DEnStMRn
NGOWmhQ/DZ3a6IDns2WrelVntamPECmrinWZXKt21BztYOxfZLHuGaq0zz6lWOru
WzoxLBq7fGK55IFiYbiBpLZDNOiDJx56+nzd1opc5CTdVsYydpCPuupZ+JJfAMbr
5M3drQc51R/LsO5tP9bcMMT+Ph+VGkZ73zhh1EAjacLUx1rqWdCcdHiZJwjVeIb3
abhBfnbPGGmc3B9noCOq4v3TUcdA5NlYtGkTjoEgRZ0jrU1USL0POYPQazohT9KI
RDvTdtzBQQGTmopsR1vLd584Toc8HsNbB8e+6fwRPqvG7w1ikxhSG6B57+4IxygZ
OIIQsspWSFnubfFgfg7hjWQxNZf30JEzYhrYOH7RrSc8PypH35cW6CVfzGa1mSU1
yIaSjK9gjKh7L8dqvkwA2kkCRydHNx5OZoj9xOZh7eMJe+jZYXTsS4Wpc26BguJ/
VPhazz8zlG24nq08xXccPha8wWIfLIGbVH7udY2vBY7Pn1JPYjGy1YUvt8252r3G
VHhuWNUEUZi/2KEQvyqTjUmmWgQt2P5qk59/TUGH3p+1gRxVBh+luIaD/etRsB9u
17l0UQXuPBK5AFNxvveBnsyizObIKOwZJs7S7RDp7/87sPUqtA840pBNj95ScSzT
/9t9TanOBaSUqGy4xJuYNrdzUmGTn02GUeiwibxHK5Zx53JFA0DP2MwX6ml1FmIG
P3G7gPeXEcpGppzbZAygvWAx0v96oHw9qmt7m/RKCpKIkR7s+lcsoD8GhBH4yGds
QxtXQLtJzIi987/nP8HH8nUqSKpNiUU/Q3H9S7OulcB+89zxG6nsipOmPoVmuSOr
XXEsczvh//MsXQV7qvKf3unLD+cUU81vEdPSdir4tIVOTRy2pQfEUW481/C0K30X
bcBPGB1ruGUKvSjlzowS+7HGKFDaIS0V8FNX5+2homgmyP7BD1oYRhIh5XU5Up8Z
Q4BFKzp+nMSCLfdjJ7HoqRp7YqskYK3xRgs4dxgk4eEfnMeqEgerohY+0ozwcDO9
qQqaHQ8ePZqL3tCIdYjSE+qkpgzPY2qjnfFWB2BeEPeWOUI8xUwXyHXgQ6QRSct+
APzfCPAaXr9KgYc6YId3cWcvkc2bE0OiPn1420JOpjH7BXhRdkNH0L/qrbKqs7Mo
T16GrYO5LcCwCim+C1GKiGhojkIACo1x3Hmbu2uOVHwEZLPBxTTM08eLGE8JZ0/i
MwuE4otP4IeT28SkTHDjL7eBoU+38MgUD/eMZN8IXyc4uHOLZ6a8pmbBAuUv2Vg/
wVlGN5eUO6KkJ6Kx9YPXYlSKdOM3N2h5rL2I39hmmCxP8kSCOTAHiITg5n6rNq1q
RNG+hos1fb1b46Alb3XD+53kPJYMk8ziqTRg4aDXLlXXahkwJnViFStLT2n+ZywA
zjgWvxNZ+JYbRR65mdrhpKQlKWrgBG1nvVjDjuY6Biv383/8m2XSBn+pjr8C3lCD
jxnQ4N/MJx354HVA/gh6zrN3/kikeI39KRJNxut11zmr9ye/fQZkyE3YZFAGCoCN
QinrCcTs3BsgA/C+g+pHwa2iIecYp+w/gRXNGNwiZJ4IFH8W6FxUDO4FluYTdE91
DbSNR1XWkPwfYxlQpmEULmH8BFdXnN+Lx0XESn8Uf2FbbSx/svutFgLt7V3fo3oZ
Sb0rICGQadOvdZKHb7OSMJNetvTSbuQx/xedc5nhBzR8cr0DuKgb0QaIwJ55ArtX
9lnS4n8HHw0+fa+0dSQcP2OGB3uHIko1/bc/ZJD6UaRGrHLLdMWtC2Va+WFPt6Z9
YvxxxvRePcTuAoqJ6MOOZcLuK2rZV3WZL0d6M/aFxNgPpSa9hjk7f4k6kZVwhz3m
Kz9r/VDifePEUfoTQ34/WpHzcuz7YKdC23h1QJr9DWJJoKOiRp74asTPqbYDNQEH
5zn8YzEXcelByR3vYmOIlqHccNdWR3Cj9xdKclw1uInfaB+WgSnygVHAD6S4Beoq
6snV0eG3EDr+GgyxSrY3ozSACbOZoTXSzr3hCEwv2ZwOaZIlqfqKBNxoB7yacGcM
J0ZMaOb5KO4J4xuI5KTAGR8pii9iNkhzUe2qfdBMDHcqwi8UIM2ofjgsLElIzb0x
GzVU012NvUEz2yYP/gRvYfiHDQ5iPPLHvDicdZ+HECUQwmtxla90RcvzTomNsWeL
mFVvzHYi2jHc6u6VZQR2Tj2zltLVn4RvIu8RMdLQfQ/SKFD2aKEcsZV6LvoY2aA4
/32g6OlxbSVV+lQaG8MtfMceFMDfHDHc6eR3lDthVnvPDmOyUoy2yCMDfIaBQa+j
HG1En6VdbcU3vJkyua+7CVO8c1UsJF/yznvGzndUskAMRUaefgF1iwyvcYCJqGip
LH6CaDTLTuFCPkcyNTzjhLLlMyyv9+QRFXAlU1ruacPLKu+SSFywl5b+8/dV+kYY
qxiDblarxX0mT/iHo2qGEyFUUco9cXRDtDDYWtljtrjwe5nspiYOu6AoAxNrnWBP
Vq7wGQ4/epYXWnqTyeUyAu8bx5qPl1NLqtRQfagQtG5cDiIB7/MpC8AWE4dsj2cS
cpdzXSb+J46DLW6k/J3lWKguQZ15ieAOazf713/vQ7K/ZlLJecEVD4X7tQyhNivy
7hapQS0h2Uq0dCVTjjtD82uBLR5vYsjC3O3hHCM+i2y5RIvC9aQ94ZVoKfahSvxS
VNCQ2Nb1b/BwtkoO0lOnIh5BcKJgOBbHAhNzVFk9XCig16BOHLQ3jPgs2hPTp2LI
EviFCzuGCcyCYGK8iRXAiQmqQFAfSjsmDwtJuYes2HAjqBjqiM8FxybAup62S4hX
+W0zo+QyTK47shNtlaOSocY3Rp3RPP3WGoU7sPMtupkxkUCNj4uKDL0Sujt+3D+s
q9Fp27x8lCRKaXSn5cFN0/+5opINkcXzYYj0p4Fq+rZGga5/+GjhMwcXtx9CVzLF
REukzaxFyIxkdQgDxn76kBeJi6nzfW7ZHyK9TukrVd0URmBavJdX6nGJ2U8vgn6o
eXr2040pE6v75QOM9oE8ViWBO7WwgIxt/kjyc7b1fYNlqf2GgPV7iSH8E2xcJt9w
WpCKWKA0R4/+NJ94Z+FHlBOUqhjm4RVh5BB8u6Cx5/IzpUgXV7ljiDWPaWoeokpK
npyt1VykaJFcnqOmNMz3LkiNBPzdHEbWATaj6PHtpypXDp39ltqbedUDoBy0ox2g
Dr+mLDIOYo1BH/1c655RTYwNQKgsEMBFAL7Yxed/l//UOnbBY3PfVbXMf7mJs8nU
MKaQRhxN497HkK1e4FF18TxWvvTMppdNOBZ+0S56Y7u/wAffKtSFxfbfD15Q2oGx
wohmt/QQbndX4NnDWUBp5vvgthobUbJCc0qMsjj0nrfHOluT4L5cemD+eGHkQ3d0
6Fs43Mx4C02qlH9SMMjA+pVGUtJigKuJeWvsjRxJEJuG77QdJP0b7JMAuAdjyixP
qP/32yv1iCEzD3GGtVrox8oHkY4a+QT/xuXciB738iiZnxGYxfKAsnaQzvTjgiaI
rp65yOcxZb8HTKtdLgnAJHPLr2nUc7FLZQM4fat2nLOe9fAExMxHDN2hKMyuZRlD
HNb2J/BBx6DHI7jJRlGSvoOWP9FPe0L+tvSPxox4b3lIpGdcHDHMsaaQQRAKaS1N
ajAEtfM3SQqQ0/ey6GSog+mjSkz/39jhDUWblBUacK7l7rWGQIiJdWLoRNBU2DKj
1ORX0xHAlVfa7g/ArFDjR4ljNOkBHH8dcfmr6uaC65s+y+SK32tVoaCxFeed4E1H
UYUxzNnqPmudu+6A0TWcFCDMJY9k1DQOmfmLME6Mhs9dbufePgfoAEljyt9VyPKr
4wmLH+lmYEFGXpAQJNbnfOGl291N9ISOwP7XqTx8+MJLg/EFiNa2c3lAw+I6A6F3
JZUe4KS01meb+vM/+3X/7BC2x4FwQ0wbpLJz/b4rsV2ngQCeof6hXhJD3ME7eqrG
06nEKySdf3Bky/y+2aCL7x6gftCCaF6+719MX3UWvn6FPt5VDY+mnQCv+kr9WGSR
D1XSvTaOMkO7tZnl4fCeMDVoTmklSx1zk2nfMKeGjiXHJvbPH5jMHdTQ2IwnAbuc
q+rqYHpa5kV8LWSWT6u2gtTFL0bJGse/8qSGeCAKh+yThhxIgSMn8cdx4KAtZ4aF
gugFU73uFc1kSOtsmJs7PGr83oCA22ZWWQkebJAAbjlaxqprhR1K5/28OikO+clG
elwfzIhDKbGnPiw0UKiDezaLvKn+bGQoacYlWJTOs2OzMutUBcc92aREIi6pwCzp
FZxApZ88VolCMmwrCD+arpB00gHpWOLcZ5xhByUkzlu9LSWaPEc1dbbtQ7jOI6BJ
a5YPtaQUportsOtZTbDyZdM4IlkU/4TtwFQgbWtlLoTzgl6l76mrkRpJ+nJE4c3l
1dmF6S0qWhzR4huZejXnCTOWHMVbJ30V0ppZHEYN+s76/LWlJm8RySz4Pafvx/WZ
fKLGMdgkGARoPC1yWezakDlbxFr3uEOYRhu3lcwAeV3yVT/NYAHm4KnTP3kWN+m4
uFkYZSNqA4N4b02HGWB9s7+IcJu3NxublWux6qnn4zpolXnxzsjq/FKQ/SY0PbNT
Etn3P86BItFrqWaLKA0YiJZjYW9qsTouhzU5i+YcYfBHbSo/sJqyOnqjWjnLF7Fk
vFq9sjTWSz4UkNsQRM78HGBG+eE7bpqCiND5QeTwWivTq5rFdd3S/Hzi91lf+MlF
Ob1P7Rsg6w2E8748lo3dFiWG/s7dfewKQ422+3uMDZ7pxBtHGxexsahK7nkvWEWL
P8rpt7DB4tm0kBy7plZMtcocsLdliKGAA3n7Q5Qo+SvQoenefkoc078iMza6A0Cs
QKB+tlB+x2cg/nD3vWdo9ujSZKOGB2OjhD1AfiELsHU3bCx/HOhfosZ+u8Kz0iTJ
tZeGhmILS7/dJEUf9sVBwWVxEO3tT1Nkr7xbWyfsJ9WruJm5EF1uuUwP6UrlaA+T
WdPZdpaODMhOXWLZHPIPY/QIAltWVLFLa2htB4CFWJ7h3ZJ1qcSiOaDShIzKuiym
lKYbHeUKFzFn5wd7A8sz9K1O5wgl0cpeLecVjPz0ldxChMBbq05ZodqwzLMxVkyD
5bqQha8FL3FiBv8ki28mfIQWJHJQaJgnxLURcHDiK/JnpbL79H7jQq2HUFidIaZy
2N4LyyJMnhfwbQCDc+ycXfWXrDlJJMuY45itVUXrThE/cYOT4YPOhMAuEvhe5jF2
2f9dab6A837ZKahFqOlVGyX3CtuZeJeLvl45Chu/SIPoexECayOvyNTCynb8Lj8U
qM5HqBnH9JGf52IWqfL4X+VBpX39jYCEA9TCYyWJZNsuNMZyBXk9Od4t6Pvj6Uyb
q5NLe8yJE/Q+Y/q8bMeeXsK5Zj9DPeiKEOUJB7wcyed6faiqKzsku785VCHFEc0b
FYZoSLpny+W4rcOOPiPar31xVSGBQfnrOMTu5pfOw1xa6j5WYDG8juJmHMp+6+TR
+Xkwp0QP0wUZ7cu8luNn8Mh1QfiGHctwHgzidtVObKCroTo9Q5PXFRFcg3arV4B5
Xs0jUgaI8SVqs2cgFQaRlIEW1bGO0fn8WtbIFvwUX7OkkNYhhlvoLMaY/zxHjxtN
1NfyqisTsgD9mVdLQrfd5TQQxfIZ67HpUpeQdjdjWI6DrUB3dFV8dcCw/g4aXqiY
st71Z+QuEn/Z8iwKUeVVGlLP4qB4m09kuOHvBFapDVrJjjl9aqV4sgvjyKPZvWWB
MQr6i2PR/PLiX7iCxL+n0BfcEG+TAadaYXYJJ0Ud7x3Ou7xzKDvm4eSVn4Y2s1Kn
5gFCIk2KSmw+qyoZvYOKoLb8AAwifJv385f3/pWTTG0MGwiWvHnPETNVDAjH0bpc
cTlf1DYGH5qL0XqKf9bGGL/aEbLkN5q91o1o1T9Ia5KkPRy1c5IOFocz6eXTc+rz
Se9hmH7JSgfsuMHOkiPGjYQo4/IYQfLpoWWuaxh/9d+tCJ7Ams/oPHv4Nchim5cJ
O7wmDtdlOOQs4r0orqaLymJI7og5+pgOzjGw11uA9CjUDF09s8K0kfnBvhTFhtQ3
OagNVp+G4xMl34Fsoj8BnB7hoEfCRd6HFeMuvZpwFmFsTuednOL6dszrNCf6KH+A
1TZlnijKUTQgXLtraWcBzzp21nlpFGwjPm1NYrf8iHVrzIviXNJgthUGfKcmpE9Z
/KqwrdvahOEteQABjnymV3sWV78AkJ6w+1JE0tlMaYvL7JltjqIX8b6YEPYHN+4x
H6tBi4RDmk3TUACWPWt4fdLKcm2SZFZg4EqK1zi+EH6hX5UG3eJqWb0cQ69qQTy5
ThOaGdZR0A+Xo1qU0+tugvYp3lADUa4am0/4kDfCa+rehuH1ODpjRjtihxob94Lj
u20M9xxmy7QUxquF0LN2D1hqYdhCc4U/tjrmpVRvggdJlJnX2BGZJ8+hdQ0QGpTa
LY5dwuhVWhvN+3oQ4rseKOPRtc7cpW5cM7z7gY6OQH8J+dOxs5Lt5Al0uxsQO53/
ehS3hP7nos8XGK9j5zVLfU6P77Dn4w7+rjlZHXYz9BohWB/mKBYYvsFGy4SGedQE
Ek7iau5EUDOOQ8zN4j/tXFUaGBX/WT+F/uOswb2bWK2w1yYebZXkUfMZLA/vhAxN
fQ4lYnd5z4CS/flZb5xWFCQtZi3vKddGJZtoQTW28RrW+9/8waACxr6SmZEBmXHm
`protect END_PROTECTED
