`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
whEWggjz6xhz9vtfTiH4fLlpvwl8cx/pReE27BpBTbdT8ml38RlivAFZwQdtNhRc
aDvRxssN2eY8yNTwvHf+Xo0aDxEi0JWsKM/nfuwh8sQ7ZQ2glgDjm2UVCBGz9FIG
qNF6viEPjJb2Z3J4uw5zvQPtmKKpPMvfzow3csBQW2vGeI4i1w4EOuC8eO+OThFC
MI1D5YRPIx0ZU6MbOAPpW3jMxyLvdg6FAmhODu/k+2uqllP2krD8nQcHXHJKmMPD
w4fg1Zt6/yob0ssHOSisG0RsEXuQ0HPuAPCIpTBsfK+R3IegY55ynP9x150VUKHF
TCnhlz6YOyuDZc1e6YS7ngKDzQPpAHhwPvfRDEM7zXI=
`protect END_PROTECTED
