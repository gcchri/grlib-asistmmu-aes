`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FMVFkYptROtsebmF6RGgOp9gUnzi8m22JJgefxGHpFgMrfaSvew8g+3Equ+FyxdG
bM/YTt1dqkRZB6dylHFLRB6mIP0UkCWMyxTOb9jLBXJ6DtHrOJLa8ONXgjaFyQ3B
AB+WjiwRotLYmuJ1s74EdS+18q8W49OZvShw094r4XOl7KhhXMT544UK2sHLeMU7
8rw4MfRcBN6NxlUffgpnapx+Zyb2H7NxQIt6W2Vf6eWVbzFP5hdxC4rr3DU0WtQS
dRqR1g4rNuhsgeKppbxidwT9CePRn2QRm/KuhRk7LBN9LdUzeG+chHPYS+gL/u9f
3WOM1tanA+QevZNuwFPJe9MoYEcmOxP6PejUSluPO/Z/HE4XTH+TeVYPpw5PVJAb
7umLew0UxFUYxVyyLtBywQ==
`protect END_PROTECTED
