`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JKlJvrbIfEASmFD8CaHVO/99yKz42e6sO7Pr3cIooHgGNg/3l3ym9eNp9on3R+E8
bRzmrZuVfOwXo4xpiHkRvPg3c8Nbu4MODEAc02joUmANVbxio7Q0Lzba/B6770db
r4GWrtGFY7KdEjt6Fha6iaeKSMssShwbvCUii41iGlWmNhXsHV5efh/mLFc6xCT6
+V8QgDRZknyWuNvVQ0WPUXv9lssEPUz0gtvGtDqSQ6whjjmzzewDEqtmzIs6lTMN
xiOTiGelNiJ6dVH9A9l+93aG2xjRjy9QuJoWCNjJOAt29XUaav2hdhTRPO9CCg2q
N1FzC/KsPzxvaLWoPC9GLwB2xcqGQlI8cVFxH+txV/R2yGSBksK7Frz/efAdT5N9
0iqC311yQa7RVEimxj8Ucz06HNUDfO85oacVAb09uDeWYMt4yb0dehcZw3pCsfAv
qd4w19TztO9blha/GnYw2NEUApOPT284V6uZ+aW2K3S4vQ5kekl1kscOEk4STVQF
D2To5g5Yh37dSfxLmbpZNpcepFKD10F8ttZuDDI5jKZS5VzxGyXHvbUw0gWCBz/j
CsSGuSl77rp4jVkRi/yWuQJGBUHqCasKO+jckg98yGEwR7KDoj8sukFjnUO2+cSx
cf27qvEUTELAELlDs9njB/bLTjkNK6GTWNPdofS++47nqCNIQ+VSzpDrdErVZVlo
D4DUWBOSn9CBNlFaT21jshGM8aky8mZ4t/3wWAsObd2242N0i7CLNBbFACOLZ/So
I8yuvzDfS4Lqpya1PZ6l6O+85qsXEOwWJj6CrJHrVoJvilvA8KWIh07KMfjsOttk
`protect END_PROTECTED
