`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LgFCD0pi8i96kMhbO/DcdWZHFn3006tfWoMrQgTEt2aPv2+SdGYmbNzwfbnGiKah
jL20sS+eA4gmiv2KeU36oGlNlm+tFLMKHpxFIJVtBcOzwkzIgZ+0yvgK6xPFrAzF
J3aMInOiQmyx2jz41vsYyrhIuJkiuQvlWOn85vKUJhZ/3OFY1bC0wnm8J+yU0GCa
vPyE2T9HeqEoGEf5hQ8MA0LrTn3IhP3yycqCqqQmwHfzpdjiEgfGxtXY4xR/LqHw
bevniWc9JHXx1aK3pmTfy9WZK42AjtGUGIU3GSWcTnOMsAvCvKHYfzTMiSaDWG+t
dX9s3CfGHRoDg3e+IV0iaqJIXLoW5VbV1g/BGRzJb6acS7z3t+KFj+MujHfruFHA
fPoy8ApOTf2TYhcSieR65h1kkAQaF10KrYHiXiMUHvVjQiWeQ/FaN8X9BwfEJFhu
1Xiq7ndCQRSiXPm05TSDb2Hnz5F+Lng0zr7uBm4ciwI=
`protect END_PROTECTED
