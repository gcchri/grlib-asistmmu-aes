`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uE4jqrtxuePQnBROUbHfWk1imqg7lLt1sefcI94S4euCQUST7c1mvPkJKmLKcXPl
zROSPn/Rt91FZ1gZM7QPFV9OKsCqmiTeCFcApeqJB7BPKPrAnKe09DIRE6bxycW8
A1QHAxcavEJ1RTfpncpa8cjqqJ+9i6y0G2gMScdkjJzjRN/fmtEymypKVSynG9LG
68ZLR1TEnr9TNc9eptOqIK+VCfbpl7FTpZz4e+9MJbwZq2FUl0I2q66qng0gLcaj
aD0sEru+gnq1kHPg+i9yPin0Fxjh5TVhDq/iHdeBYwNsoHgUSkDQUSnS3XSbW1G0
BllKdrQzaJnasZRuM81sdil01odFgWWVBAPgbHcKne/F2vyd4fpC+pT+FXUq7mGd
RdvcC+YXwLO/HGB2gywItxKh48Q5IJBUxkP7KK+HsJkO28s4kABimu4yGmjp6d02
Msnv/0PP0urRV7TgqpqI+BpvS8UrgFBnY0efIjJvUiEoonyv+0H4Q3ZhTK/x12YQ
lNeUU634UJBxw5LI9enF+K7e7gHX3ciqLqxh/9e9GhLXKGHlNLQTc96zlEBavcUi
eiwO2RBGABbOGIQDQPUSMTxswX2I+2qofrGHzYFu6N4x9fyaDRZO81v7YftBEbVb
FgXoEzw/++WvD9jrb5lkQEctmHBHrk1vzNAjk4iCMVkV/osYk4yYz+hoc2A1U2qX
rCS3xMCZ8v3RaBc1jD+EDxuwieTHrg4PGzTw3OP4cbT5cWGeEpz3PfDAT3mi6GJ/
4mVuKtS/ckCDCrpjMZGUTe+FYv8jnnJ0xpKFPSYRmrULjjCEmPtNmzVmt0oEswVl
poSffemwUPj3EhFt8qp+cQkSgCYsKdEiOEkPofGIsXfkXbKF5f7dPYsEn5W2bEVd
62N0p11QhV1QXO5+GWrpj+kkem9YcOJ2E66v/8HHKaA=
`protect END_PROTECTED
