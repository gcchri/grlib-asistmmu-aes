`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8VPDhSGyeaG6xxt9pZ7aQpyI66SM9Bs6QC3nBGWOrYQ2PFrdWwDiTdY7Ug8rQm8l
QCgV1XCICRjQwhll2esNajT/re1n3FpAIropQcb2dIY/abxKg/4Xq4gWRXLEXmVc
bFZVIVNY73LPL5+nfOEQ26WlG4oVCpH3YeVea35gndZyAxG800jmh7RIPdltvY9/
yjXGLhNeEBQuShpuH1lak4aCqMzpnaoEn5dRvfKD8TDTFVPavCRAFX0zo6uW81fA
3IodpZTuxxT71J3VxAQmwwTFT7FZrnQ1eQv1FsKugm7932ywUywY5J62PY4qaO5L
W7p/zx6LLPDk1mQp/JCIBZhhr0Xk59xCPtzdmM5WMGxEbXoe4CmhkKClNT+02ei0
IONJMRC4k5ZGqvXntWX4Q8QktlFhK26zoz1TgtnADUIzZHvKkZapJQ0U2X1ZV5ft
V5vOCG3XyQPpXwYcSS+kAJHpm6kKKJvcRWMNg/0TIyFvBEDnp26Fb3igMkOizNM/
+6OPmyzlA94BSzINBbLOrwgCY6Futka6krl9bjfLTgJHwELbkOEAexMoWbbKG+/Q
sXF5UHMy1sbnShXZPKN56a+/YGxCneWpYAl46MKcU+dTb22bCvepKwgnW9TmidNI
3bazG86rMzUdEov0LDk5D8v3pzPPYxwoklI/hiSmQwjvFhvnlZrL6TMFfHIurWnv
5ZiI1lnNzBKkwAwGuuqOTpCKavSsUzDhpcUodYE+ZN4qMBGPJUdv6CjPHvyo2syz
+JBOXDxFf4fvlZlw6WnR/OuDVFpVzYeS2LbfnV/Py/tOGgsZG1zK6wiUcKqqoI3s
4/+EPD/XSA527WuaQbYiLJI8WNuC0fExASuqFtXu3eEBEa1XYMK8mn4+16kX8rz5
c8xKmu8OnawClIP1D7LuIViYcELf+gQF5je1FVnq/HmYRyvAv9anE8n4NQQYwKtV
XsPkCpA5FQahRHmKIg1zu5+uJpXGrgYrXv0BspRUluYLjtADw2KwiBfHk/tgsfqN
Ui6qo40JF4QAsrKf3FA1gItwpSSKyciW+GASRz3Pb5Y=
`protect END_PROTECTED
