`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LxVjrTlKDIbKrjjaYiEanVCJhIZFu32c95iGiU3mE5Z+qk6i07qptk8mK+k7ana7
HL4Rg8PowNIbtxCYN7QI4w87ovCZGAV1W+lVTk8bjo7aKBUetGEexxCwWmlvGcrM
CQANyJonE0TtWcLRIAhxx/icJEt/lhJ83+sEQ41a73iwSAz46y8ONvMhBZHvSB7I
psGA8IC7MyTqRSOoKkq1gQvBPsUoMRNjNrsZW8eFOJeL8NgTrtdlgpHTwPL0zNp1
MOhtMte4BF9N3b+6pYCL8rqNR6aF1N/22O2gTehls1rZ9xLwDtATN8lD/usvq71H
EKG0RH0OGy36H1VfMOG4tCKSSWgq3bRfthfWnmxJKT02oXT/bTjv2nQ3vvW7hGPz
9X5eCpGTq2z12mKaQsdwO2/YPr5soFSLVPAMdhCmLO5Zhp1ZVAUB9C+0Wkqfg9BQ
JztKwsD06uJtxpBPEsw+Iw==
`protect END_PROTECTED
