`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tPon8+kEnQIyNNUbSDO1u5oJ45+Z5SX/oMfoYNFVhpR3D7SewQcfIGB+a6uN9BIY
/JVp8/wsTlFGzuBVT7oGXR3VE2gDmNnQx2VijIfWVi1p2sKswWAfhIfZ5L0dQBcN
hveWYttfXCRM7hKV+Bvy7Z42s42I5F8Rh2RTdCH4UxZLnNgWelI5w55RFHryRLqC
Re1ONDmfoixqBQdI7pUc7Ht7MK4fjfUQukcQzXh9G3Amlz/FuwbSjnC2aruMFcEu
zU7rAyHZpiChHx8h9KqRnuzi+KIjGS6vxSCreb15d5vdzJYGvpO9ylNjxZdCpWDK
8r4g5fkBb8rWtCPih2bHOLH2qdMhaOLQEZV9pP3dqtihMVorTDDYRtwc3Cz/nBa8
6c1mYvjPRQK2tei0Ks5qzdyp/cHL/Jh9VQI7YZ7sB/A/BQ/bEwbll8Vm3i9F7HSE
JZQ9IxPW2RTFMOvmuGohIKzLmqCtQYA7Nt51qZFPzSWTlURgjC7/IUg+Dfi4E8Qg
`protect END_PROTECTED
