`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5lUJs5hx89aWO6sUldO+elenqvs3rvB5C+pdPf9TPtz+hTiL+bE1hS5GDctUf5oh
pXvumwA8Rtsu/z7EkweMbCuwzTZClb2AKWMJxdcfuAyeh/lXej9kkPQ0toxSYWD6
SUcnEAFv0yl7EyLdTA0zfHayTa+DHODYxWLLpXu/VALvYAx3CaZqtACNeL4Vy1rq
v+fNZ6h9wT2whfDdkyQ4+BSd4jrqFIUjwUy9t1GNLl6AUcoshX1COM1PdYvxdu02
IKBXuYr7EDHzGjnv4cH0hVT3smBeHXufaruaWZZ/WS7W1Tr2tTnSUSN7LODMqx5M
yt33sZck7sJDtSWvi8mpSE2YGNO+BCQf1pl3u+zcHaZWz4GNJmbkpIsehJ6u9jUL
sat5fBIXwvOg7aKAoQXZmuFdfeOfIgBdY99ITKfq6uWOVpr27UwilGTzUFAJfsRH
LWE6b4U+zkXTFbzEO4SIeds8fo4V3YnQST14cjHdrTS0Y4Ap0Dxa2lYvdjYYp5m/
r/5t63La8urKDbS1mQ+Aj0ZAiLmMlNRQAn1s1vcu205szy06IsrjCff1udR4/3Z7
L/FdO3hEOQb6iXF2KE3VDIQePftgLiZAUDGFoGCTmGaUxBpHPTQPbmhI2vSdobem
/NaocBkVmPYkcJlCI0FSJnEwq2pXfFuHK8MYaAUxIAWu8L0prgix2/kTRqfcfDup
AJ/26y0ULNcSiEK5fM6CXQlrs+55qbk+yCoZOGncEBOJg9nEv/+Sa+An9Lb35ulT
vhLVvtKJ4+hFtNPQk0VaLsaPRuCc+hYAkZVuvLSC8asjZSaevuxjdnn0XNNj32oz
EqVWMK52nIUOHTB0WUpwYJPvLmL+Wlif68RJvZPxH9A0ysZxzuiv1az0WBa0FYDA
VEPGOFM6Hsf1+r4sHKv97P90Uw/BPXv3RCT/se+SAcU=
`protect END_PROTECTED
