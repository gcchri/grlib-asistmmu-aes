`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1EbpLZQ8wnJtf/vwDuWbhS5c6MoaKzeDNlBFKZr663YmDdfeMfJolzEzPVEuoGtZ
f3J5utMhOOcKmrJh7SqORMY1GRw1LknjBNuwGNtXQvI48IVAz7IbwiyH59uRV9oD
wFVR1B8m5MmGbIc0Z325mzgRLqpKw4ZjqyQNJHQUMmaAvd1wasfZwLnj9u7KWLr0
F2Rkg5Yx/+K5/1iFRpGOZh+yiiDze8fUjBWqJ27vBdTee8T/OW/BkgJUPj3nh5o/
asKlNzmfoNTDbBCYkoMmm9YZgNlNFrDkBC7DNTi5UP1obRH1NvuxhSbiMllOMbg1
kvoH4vR5BE6bNuIKYVQqP237RwPPvLSGQAMq4HESAuyDW0c+lX7FNaGbhhOutuNv
PN+ZzQ7ttl1e110QZKvLNIpnxHgu9RVlN6N7r3GOs6T6TE2XrQY+ae045+a2Cn+U
CcjFdRQAPcvvwzhO3m6nbkDCyBXqjt4ex8xoDXzSn2tGR12Pt6LnltnHrkPsEDkZ
uc2/TKjS6u79IDhoq9NyRfMSS+KINK7ONikgqrnzDKs+EB2hEqb7WKp4zkZ1usvo
s3lX9w47ih3UI1OskcbJ1CSgdumkzFYjzAXQIxsBTnGL3TDyOdr+sqEy88rJ0fL3
y/PK1eYHNeteKEk2qsN00QZDuz/Jy68ehN2wEoIgVWoAuAf2EDKORFZCuwCFCb4j
zQ+yTl5Q8/sGr8qgcXwf/ZtcfgXSoQYKhNq451rssHPJKCeLrE69ANlanExX6UHE
zLAXvSUeOszXyjKLPJT3tT4mYcu7/LEjaV7Wr5AH5yY3fQuVfqQzY6MorzxcG8gr
ioEQ8ZZVog3rjS278mMihTmOJUwhr677REr9juynLMVCpPGWxlJ8KGUDVFQaN/o6
u9JIVG83uM+/AXFKO45AX3dVc54W9PaB4rhosi+vCZHmO2aDm+YGd2NBAK6YGAkn
XIMz9iglTHfJtlMK6HwX5V4kH5jB6jlT5O2OoDw48LCviypZfwRISjIhYJ0PAVWh
lKR8yeCYeLp2etwmBrlsRYJEhvG0mzSuFx+RRypL/oS+wd/HGy6RXEdxx+oTAfPy
o8yaTi+5JZ/D526VsOxNc7Ibz1B/e0szthBokQ4P0GxTT3yQmmZZqBS7NPVAOaov
LTA/X18f4MnTSseu9re+GAreDonCv7uPt3FltJObRlBJgXhj64+2GY4LkRJxzySp
RKQyxQTjN5vWEPf5SaRrMrOsOiIvFayOp2yKdPCmhrEdsLMyKmjclXdPfbiMh+Bw
`protect END_PROTECTED
