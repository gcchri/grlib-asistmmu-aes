`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D5R5nJn/VTVDCq7pPm9kjGWR6+m0mT7JstXKUahsNNXzUOMH3sIyZWv7HulZqU6n
vUaVLa3impVNY42N/fYSl4Wc6l3khY6fFg471m3xW6Yc/zj7U6Bml7ONHM+hD3O5
WUk420NzK3Oa2IPoyzxBJM+GNvlsbGQkMRGoz8c7w3tCNsT9K9+Y2EUjnhzm1keI
xfJp3iWL6c0pJbV+ebQs08i9HrYOOe7nV6LoMqgUD42OfVCKjw5Huc1F1GZ9dr5F
oYgF/XLGCz9v8VS/VAIExJzEeImoWu+dDYVTikwHnQFLAmks/ccqcilM18hhmGs+
DHu+QXcAFkfCGnwS8dL//TaoZVqZCdqlTTfycIE4+IF7t8mOxgS1cQcCjrJYU6rS
/Mx6VRLR2BVJsntmPJSnTnPmTC4sh24wSV7xFDmWGf5DOlj5yjG1UqodJe5Bd3mt
6CgE56bonPuJthg9nebbidKQt9CKb3vqnkoZCkF5GsSIxJPtZ0OrSwgOzhm5pDQ9
vvlhYj7fFcu6lEPdfISIEvJvrmx0wSm8bwT/05Ia4AVvLDyTp1MrBOo3bCoD/P6T
mrlPnHwEn/JS0iZQ0KHnF/VuYRFQu1oqlUKiAObvvBQ2RFdXPUEJWlL/RvFxA2R5
EUkaeSnBN2aCOx3RGZD4XCuwDb8woRQg/empdbGXF2h7ExEh8+iXeskInNI1scmc
4V/uUb5h2WYkxOgSDbxlJyWws5i3mQr9Gsn+OMpKJhC4G2obB1QDOjFwNY2OkAai
2pSTVtf74tGj/wrMTO9hZRngxv4pzb3GcBg5Ty6/OrzkbhuMDzVjmzFMXtsrTF5x
0+4f7OUAJqLW5oc9Ct96vqDX84zZK2/pl/RPR4mNzsDARKkdpbPspvO8kz5BOxIp
ZJD0Y873o1HqO6k1av/ALjG6mDCiQ9DZjbehi6+MfUaKvVvJF+l9G7wvRdfK7PQj
+GmefPOFIUfyFyl8aTpZPIEsWGI4gLxl3L5bfq0iSP3HDdX8e8mC50Fgzx+R1jHT
ejXO7oAIiOkEnkX40xKlrw==
`protect END_PROTECTED
