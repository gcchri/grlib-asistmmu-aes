`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+roUv70j6iIB+QtxdcjY0Tps69/UYceB8yhY+EsSWSA+8Uw4r8qgHNgY6SaDKJS6
my1A3UxvsDcL5vAWWNW71bup3dMr5qbw9OfyLMSVyfOlliXsizS3gkiz+Kcd5wXi
tEr8KKYGAGPm3QV+pLikpN2bVgTDJefYeWxaUFOSwgDdLJdVdyh1AF8D2NgG1z+F
VJMyW2YhB5kWzZHACA+SmR9KNS2ARlEFtvvZ1jZBxivF3hGlPBU+d+dvUCassRif
dyrKKB9HC9yVQl8jtO4lPQ==
`protect END_PROTECTED
