`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+gwtaRem6yj5+lRYOdIKV9i/5nD35pXAdHYj6wAbZxOZxejdXoU3BBjtgcrq2YNj
+x6DMcZNtDxz9OWoAajNKlxbcmFMq8O0Ua4yIGwl4Uy1N5xkMLi6JI8VBMe+OfH8
TWZtWOEbPuG3sHKMHIWfOfIklcT4nB2KL+87H7SxKPyze0RZm21X7SOH/xq+yvdr
EQN2PtRIgKF/0BSEy1gNYmGcLDLlsMnNh+VhuVYxF8BJDUf07jso3cXIGY9ZBC+H
x5fyGeM1MzuRDR4kAsgd/DbE4RdvJz6fGbV+Y3dRccM6LVp8Ojm+39GCxCTU8psV
3lSZC9j5+QqMQc70wTUN9NwaS9f7uNXAHFJHef+QSyPhcW9w0YcU8olRz5j9qHQG
zaYU8tgRGo0V1VLrtD5wHQ/Q/GrgR66arJYh+CFhxUButPSsL4ZPam0QPpRANaUW
uNSzLRpHFgfK+mh3yGWYQdJYkjSQHTlVC+tPCypFadIRJFzhlBALg6LnmYWcDNoa
+LLaZS0JmRG54z7yVS3Pcv18EMA+NZWYZDxgpoWKpQ2iJA2fAiQBBSerhKLLLmy1
mKh11Fpgju4RqMZYbJIqkYRoY8Lq5Bh3IIDCzyzfEDvYmd8EhO/bMT6g+YYcPo43
k0XFWcy6U/V8BaVxziAWpPX19g7H5ZLF37+d5b8VvRfBhekVTATFWDM2qqJVNjw6
ECqZtrdX5O6Qcgn63Km+nEQGrcxi37+ZjQMk2TI/ojq48iERPPRR8uEiRmCGRDRs
KJq0O3mLAq1bf5f4DCpiHRsGdIZqDGc0xK8QNlqTdjrFmv9ljy9+cQx3QVpVHO7N
SfPLvpcgUUN7i6+XTjgNDxk1UkV5f/IlJtBNCPHAOkTAaMNCSemJ6eVlPhsIwtbY
cerFo/OKmTGViY9+sVirpw==
`protect END_PROTECTED
