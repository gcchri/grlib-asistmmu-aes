`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sgcMCTHqw8jScI1SUmzrr3EfVsGOl4bnv7v3EHjHJe5r6zWnd+6u6dSKsatdb/jA
AzAOhShgU98/LH+2qFw9IBOGpYTM6KDY9KuViyF7JsKINwQax8SRBjPDHVkfUxkp
MIAVso/gJo5sI5SppHOhJzzPrCL0h+VnVTb5EU2jApYKTFnlsWuyA2WYWmNXNNlg
6lIXIZDg8Dv2MbXxRMqlBLo29sNh9YHjkqXU3guLcz4sfc6FpbjIGr8fNJn+gJiK
qZdFzpnSidKjMrMfd3Dbkv3dBiQuxM/5CbcJFdZhzTe3ouJgyDa+mpwMySQAMnzh
348be8FBtSVvOY1f/hJJrrOMijLTELgATIuFFcLyrVYrIhDACs70elgAwJN54sC6
ipYjs87mWh6MaxX6HnmsA/DuZu90DKgXW7GQObuzUVQ5aYCUk/g44re9hBU3J7pa
cXshyzep9llESu0kdDdtjHyIVKgSYf6btK12riZuBvVG2wnYptVafYj6nvdS8Eof
r+rKsxTd4BrhqrE8spSIK8vLLPtOYOs+qL2c7UmqxWAj3Md+I/NorCcRppRvk751
PwBBbMRtJbmRfcH+1XP3vaiqJFN5XmyaWHc0Q97bjKjsFuFSobnuHNfLh5I3cKUs
DXCLv30QCnVYUtRO/l0ct9db0XqNZVr0MkVeUFWq1WES+GKU9SBsIZalLcJAfvnX
Ty5UkMGpm33nBbUICLOl4iuZhSBPkLawnRdc8ZbEJwfllSnMKo2OzfwI/0PNEuYB
C7knhPCQPOgSNzKZ4vmMCg==
`protect END_PROTECTED
