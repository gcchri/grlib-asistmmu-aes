`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1p2M6jCW97HVfOCclkiAJIbp6C1IYRr94IgiHbn9SK/jNAVHdaneKo01wbs4uaKC
gxPtJcLh4DbIbzmgdf9U9wWgWvjQNcT6lG03/OMBMBSvIZoIeLVKSoX2aEkqNhaa
P27TWvCkqy7WADjxkJfVqK0T9+OJWzBO96FDyDMJLXTRddi9kxUFSFVcqHlyEJr1
jw9fJdEdKPMSTnx+bc1kKknHoAk9YhC+YhK06Dsjh1zdh42ydKJpZ74m1g8KxjFj
vOrVJ0MttuiuvGc0t5uLGsO6NalOL6qT5JGBUmnMr0XWZBUgPgbHWSIKXsnkhrqa
mCBlBqxOEyRBFtVN0+XgBtc2Ujf4ngl3uY0kostCXF77q7JY07lZ4SkA9vdyvCkJ
ajF2nEyUYiQvOeLmCsH0bc28t74iJbpNVJ/BS+gKzDzhQiCHxL7oxy+01JN8ARtP
0nbRkP6tcV6fsvWgc2KHrxjWu4iCCteKYhvE2a/LvDJbppxlB55UcE0w4aEETRNQ
1P+X5RieE0tQvwO0y5R908X6lcp1C/3x7zQlAB5e0tuWWbmNcxwI4b3VnYXs56Ue
OxtNiDxpoqyD6KxXd1rqMWkIZnhwWWxQtkuHgcc5f0fY4WQKetcsRDmhubVPK4CF
Ee8HcrmE0tveqYqsKfv/CWgRLQbtSs5Nl45+8HkAxD8=
`protect END_PROTECTED
