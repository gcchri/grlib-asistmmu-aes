`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BMB0kCAbN5WBMYX1X4xkRtsb0qnvK2gVs03/aGAhuOWwiHmMwuVi3rvKoOOFSdLl
D2DDeUe+GM/4D/Pl9V1L6oCl0ROpdngEv7i07Jj06R1SKPf5jp5G9KC3xjutqk5E
R80LQ4hEe8+PSjPjA1XLSzAcYM9zWzZFXf2UbwhSHIVSSsMNv9+JXngwNKd9R1OG
9RnnMont8gxY5qVDROhLVF9KEoFXx7RcoNAu+au5jdwo4MitNePh3x2TB+ftV8Pa
lNibZ5WHG4oSjYqE+ZXWZ8XmpqZmuYTPbfflFq4JH8C9iAIl347mbztZV5Eqie/m
L+aG/Eji3XbBss29UAQYYP+xmG0jxDGsbWoEWMndJBTSFnv17E7oMPeID0IGpI/O
3d9yeKp9mYsOhVJFTcIxp0GPM7vqVoaBu1l3Ni7KkYaR6VWx/MV9cwUM7IsnbVkV
`protect END_PROTECTED
