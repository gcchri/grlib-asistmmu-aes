`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FzaS9/74qtvlFRhrw7zAa2FSSbGQf0Ak+u5Y/k2KwZPq0PYWRqSOpifrjvDDRwBN
UdHaM/BhYnnJas+e0EhYTXDfdIlGpDQ9czZfv6hIPlFCfFhUXWCkiJ433zMwgCHP
rvE3RPp42w7JJ4crAmlMZt4f0WGxrvUa00Qw6m17UdlocvYXwFBaVw2XEIu22UQN
9f66CfrOhi4QAWkwxqwCrbyxFoYjhgH+pNPw7rp/IxLq3V5KnZNk+9xUqakSpPs9
JWXFM7a4x2FLiowzq9LRAcOdFoeir183zYEoWz+rY2C0RVyCMJydichvvbmBNaS2
wHeRuU9I7zfCJ7gQkM1qfuT7Fwl+a1yo9lDvhXPxMSCjg+sXBucl60wa9t/mQDeq
xWJPlna8w6m2X4+B2yB85r2jhwxPY5IVg2GJ4TEoahuowGxaJQK2MEDvHFR4reQZ
N7vOjK6+ETdtciH7jmzIjQ==
`protect END_PROTECTED
