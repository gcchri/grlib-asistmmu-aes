`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OBbqttBV2WM6RUxjlCi5tPty7xOVMxXUBjC0LYtoC3NhllDDlGfd/IKG5eMbas+D
aBOxCLzmJVc2HDEHFqP6NIwv1aXY30CHVMjLaUgf/dWxcNzBCprxCvPAonvwPIST
1EGG67filisTyiFPh4plBojMY+4QYa3s9feVC8kfkxYoRn9A1BxrW3n1A78XqjgJ
GLl/zL2ACgaCxfkaYomwEa+lrm6r28w1SNGPucSBtKaGQRY7f8vVkVAXtjaw4DqX
ob9wSpvARGWLDZgjYK8YhgIIb8oZjSEJRbkYFya+XTTEQVXWOUT88DPHVAB4q7JG
kyMnAC7CMru2jBjxOM1EMLuW9B5Xus0EoEYnuyKb+9oNdHJuPfkTOkjnfl7Qd1wp
NFeADCPpqfqGldxqfy/+E5ofZa4VQGAH7WM70I7ZjgDFR9E8mmsjFoBDFQs77DJe
`protect END_PROTECTED
