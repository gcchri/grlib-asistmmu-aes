`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d2BdLrJiFZ/lNxP7dbWAEe7Uniso7hs/jHzMr9Zg7kNaQKPWQ4sg42LjEKi5iiBP
RBA9zYp9B+esOyVXzg0mbVD1AGz7zo56zfwwmR9RacErhP9ZQHdoPMS+1Pdko6Fs
kGVQvDLSqEHjjhV6v018Ijh3qGatTEuZRiSrpNphdZW5NkCRQESRYYqeTXdNY5u5
lUb40QVKeM+yz5UWa0r6sj+0wrJtFx5ksn5Se+K93jZ68Cyjpch3Et0fxo9j85/r
G4riRoityagUvS6ePccvLx4MU4OARLCZ18TxG6sQsuVKDGPJTI2vIOIi+IceQajT
E6P0zfw1fzEAETDQChKwL0pH5jqp11kYliuKvAFTDTRlmqZCM7jfj8gVZQFnYtPB
M6ojVrXmxZ4GfptIS4RTqOUnLeg1zIunLjm636foyPWZ11dgtBtSAOic7Cd0PK+6
aD3Vss2KqbV/5bOfxjLLydi8by9VoD5ZzBL/xEBGHXk=
`protect END_PROTECTED
