`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2iwGYzh55ZCkY1zf1TsdmghtCT/UIvohPZ8HtkscTY1sn8cMPYM61Z4mfczV2wZo
DgaHRBxoTxP9FZXt9uRyIC0z/Mu4vFGFF4ff2S/aqCKUAv7JaWD6ygZxW8vpcyeX
YAsfPVGABYSFL0zA1i+7VJzlB7iF/BQXtny9eioS+Ky9tYjgezPxG0KeCx1SCxgK
n87BX897YyBcqrUT2MVuhNu8Y4B/5A84z6Z1hSvRW7dSwQ1Q/nHGc0aHbmqRt1wA
a3Xv1Cc8I2S7rtGtL5FcoPdvY9hBe63Qt4vEwVzMchEfhPtSAJXxwdmTBMCHvKM7
lwxqiQD7sty2XbxceXhIShNGkgqsdMrCfkJTuT4tqg2vaLI1BZB9PXZ1MipBt+Ng
l1GlwEfVPhGmdc5cH0w0GCVzHkS5/R0WN5apfx39N8uyVQ51KrrRR34wzx/BYnWw
H63c90WoAeamR2imx2KE2S3PBFPpKTYLUTWm8N2MMlpdo6J3eZ42F6b7yYkKt2m1
XHmmqGpmSVpIuzSsHJTVxjq6TminphYSuA3lFXGuQ0R1TE+pSocy1/xfz65Y/+H8
ilVbfEbiSfAfR8nD2VstdmWfef8IzxYafBLM5ryL9HprRkG6wsQecF4x3fZHeWHJ
RINjkQs72CEGnjKHgQlxVxx7l+rOwbBCmMQFH6i1Mxt5ReUj2Q1+LD6+4otinJzC
SE2g86Na9qoSZV4NfSJgancYUNPc41wDVxZFT4rNgK/DcrMLEyykckQxbods50uN
3R9cHTJcWfheNZ/aq0t/q+7qV5nn9yxe1+9Lfb29Wuk+Irb7RulcwuYBBn1LsnMu
ahwTkT8ueq8oVqxtnxr2R8NPRxHwtXWQCKV3q07tGKdMfDvV/LHFC4HxgKQH2Yp7
E3LhwATpFnyuXF+R6qgotP+w11nfNjDk5WRy9ONOnlUfrTDyllFWZSb6nS1b6nAK
AcdcBb22ALMi41W9Pgeme8Tq7npgjslxdx4l6cacfIMmcxqBUemgy3c9Z8Bx0QSd
KgzDVaVIm/YDj+WUijtwkoro3+F9TuK/TqSi0qevO4tZb05xa9lBF6zKmtyxLvwH
hsjiFgMsm9eSzJpl3NSpIrHpfEeDZ3W/ag0iCuQd6lRMLNW+2esEjXpONXFSu/cE
zWdMFs4RAHH5EMKCgtm5orYPn5flm/wCVwXoUGjdjvqXfE132scbpg9zUeBvCLgs
kprDj1I5u3IYK4nk4dOv9afhk/7AC+Yc0V+rGwbzzrtf5svq5kEwjzQ0PUG6iHBW
Y2VfmT2VMYBlIAQoj2p/akRe2ZQ5HrNJBgpuHB5a/f/zH0vANI1FPdpxCnqrMPtn
Rgo8bmhIaWCI8rB5s4TPxGPpFezaLl6Sm3hD6rkEMjy8GmPXLBJkK2ZrAElDyED6
cJ5Z04Mv+r8HVAhiTQxIt0ChvoPl/G9y8/2iwKM11Zb3CuES7PsA8+1hFS0lYvY5
OZftj/rcinPisX3VrcHnhBXTYL7YcH6awq8nbWmdW//z8JWPL8B5QsVmrSRALQRQ
HVPTJznWszu7kP/ytMX44VZuBS4bxtdN4TzYp0UY0kCMoZ71MY8BIT8C0VG1/sEs
K6iWZhXTGeTdW2ut1P83v97VubOKzcx7c/UKie5w86odZ8NPKDGQLo6u2KTdjpOw
wSeoTMT6Luty2+NItLt91MbHjET2qhXYnF3PMg9JJn/NDqNm6BFPIKzy2SI3jvAY
AFENtUZEGjPztVwtuPPFnkAVPKKMpiVf719gsZOwsyw6s2zlfZ+plcdaKbIxnBNi
IfHaLkOHBIFFR1XZwVNys5Jp57o6LVRSMcKOtLWqtxC+0q5qD+xpcicfteoje+Pn
aAnVMPF2LnmBbIoLVn8TRqSv3pF/0rplc3f1ISeLmVYiwJgmrDz8crBXCkGpjLJh
1pAdJTzuvLapVwxLcIUWLxGmf73piZwQz8zXucLp9GfZWwWxYcy/P+7j9ReIc+SO
HRWCXIH9z/jmDT5BzpZGG+cZGmi1AeKMbWUcAAqkGyB3KaN1xvyTBQUH3TbkFK3Y
/edxerNHXn/m/+JdoRR/oJA/F3zeETWSNiwye1IjVYCFG0NCtWr80RUxqlzvWrDs
mxoJgf232dAKxi8sRm4TyCL6RKUtJkb+tzZpucb/QJY=
`protect END_PROTECTED
