`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OjQxoogSKBrh7op98J6Ohm6DYdgp6ESPYQEfw2CtmlovaZfdQVq0v3R2pMwaTvGD
rcAWUBj9cSyvfrZtJWvFSJ3eGjsMloRsXnIPKxr5y3AM/n/V50OoC9THWcv9DREp
uXYP3iWjrKM67Sed8qE/MuoEKztIv3AVhcPGRDOHKhvNKLj0wuDt0RoDtzmkZIP6
weUQmOYNd3hjpYGCJvyFAf4b9n6ohSZnLUX4z8H5maV6WHEJaEiyX0CqCUm9Tzsn
TP60XorhyEC4y/7mtjpujk/v4NzO9F4XdbHf6MxWRLwbo1Q0WM2Lwd4FPNWpHXR8
zo6n07Pg67pghRHlgIzU2t4s0X7QeZz/Bi/kxpjQ7ERQLgIl8kKuVXoyPVSyAEh1
iQnwEniqPNyjCVMyxjCaQftJC06F5wpw77HMgaIivrqThido4sJJ+yfAc/MuZnor
ZuRUmO/fDj+j5YCXs7v7+sdUfCfW1Zjug4vfhNA7mnjIBmQ8w2tMyIsJ+ubJFvGg
bbNrUcXDzlDsKMsbDR/Tm1Bw95UZbDrPEFyRsVyXuwX+JNkoFpPVmUFpHwkZio39
VNNmz3fsSb9GAwbxYNHSVAjVbBDLO/+tz7haY/EFupe58OVzXiliVnf9mPovs/ER
cFfZt5hHPHYmJor+s1ESXYOfnQmauEciTLnD4LhUyTjLRSeaRsAhqzJHNxyQrqCb
eEJw1knF1X4Y2/dexv8fLhWsfym3OkMDlPoapx6foSpMfiP+sUlRW4NdxGAOmcp5
U3RymlXabj0ZDzAj5VgAq9lFSmelsu0RIC0WoPT6K7102OlYgcgGPfkZnDfiH2Iq
oioAuR1LxLLC5PHmjpaD8zL3r9GfInoJNGY1MYaDoAGGeIB3j2OQPM8e41JLeCER
ECds+R7xwswzRwkYkLoaqkVLJ9eNN6Umh/XhWQdWt65Qusg1/dkEhfOKMH8+YGU/
Il0SlVIC6UuYPyPIrP3Ufg2SvgpdESFhqCZrta8Cs/R3ScbUHCOlzoQ9SZhcXpEC
OQHEDICknXv82BqO4yh7zVjNqRD/FfGNy6e7KnF5UabcmXGAMGfv6qj9c6OGKasW
sfyn/X4L5okqhqYWgHTIONVBW0ewz8vfxdsYCNXrmkywPThUpg4ipFWPjpnX7oWV
HQcMikAlM4KMXHaM18Zuda8gNcSaqr7qJMBYyWsGhVpSujFHO9aZG7cMLjG11ysy
WWCal/UsAptUfjxfNA1+hREBaYQO+oHB+XN+mjR0E8vEVsTGhqE3PfYvTFNaS+HT
XObTtR3rl+Njq+uPww01qEkUSncuskO0mx2wMX+3/1dHl8OUEjS7FqLAze3WpJHi
7jYUns/3umK4NeFa0pQKPWTebL8Iilmtwe2R1cX+ULohQhodgXK2mgoyr+cIj+ea
7zZPUnUBVWlDcC8vczudjSTydbgSv3PLSgJUKmnv7xPcxHG0T5g7wq5plrOMjgM5
jvi4YoIbielLE/Vj3Xi1vweLSg+a8M0NYbNkc1ytBFI7L22AptXgvSZtdkeGfL4A
odJUkrfV5IpOCsHbz2lvRsGk0IlBlDUjwaFuunC1jc8wyF+6LiogTtdE1900CfPs
01JVfHN4nZbJj/VKmwSsi7oTIAQUQsMjJRaYpJrEwoTUBWqR/AQthEpzQOZqJWn4
BtJY7Yj2G+BcH0qy8dPUW7ffvCPSsAkuGjw3yiojhc56rlGpXtUXJjyRT6LnPHjQ
D/xjTgs3lj2rz0LCjzDf6251g1gVDD0QLrRKmlKY8Lqi2SPFu/8RKezdLoNMQjvB
2cWqZlYIoQVPtJAv9izroYMAIXEwuva9d+eT20qLa67HHbcUana2niRyU8af3l7U
mMafPsx7syfFebkeY3F5aBru+TXiEIx44+ynmdQwFYF7dWkSUOwbqsjdvQd14faJ
WehD7GgFE4bAaRAURdVWvzIaLThZ/ETddpefjevPqkOewTDpU0+Hxh2uXueqRG9v
6iqhpeer6HTtlB1JsFriAbrYOLCiWLOh5yx/1SZvbgJSt0LEYHoHa8A1D9bDx3NT
aFE2RhU4gPLzw/WPNr1RMH8i3LCD04r6iHsqV7s2F8myO9GPr11I7Y14sVtCFKIi
5d+77P77YzyJIZl3CRRFOHEC2Zyqfz6klC24rIl3cVnRlJVkhJoEPagnmU56m3rR
A40cKoS09YGdc1E/Lx1OCYmcn5yVAyziypAQXnrcOTcXAU7W0V0dhQz03MDPJH4e
zrgWu1E+GHxSMLj2lkJhkxKVnRE9+YjUodl0bdFy+PPMpaH2Ww3e8hYgpsGNgsfH
1SRA4yGsosckVpfJuZ7yI/t9iWL7cggJv9VElheIwCjdMKJOz3p4gbVjVg6TfDve
nygCvEZS/EBZ4UCTa1RowFbIRPC0tQGdP/WTgRA3ZE5Fx+NpX2GPy6Va6moiXZIX
oUw7ZZPMmmi3b1KHHVjz1EBTe93tjezJjEJHyYAlCbwJQDBqShb/qytkBqCct2hk
NrTjlR/n7uaW9m6o0uDSPeMkPCF8fEC8sVLfux3lzxg7ZNcgjXmI9Jpz8QCqXe42
qQvdZQvHcgYfPVYfbgenylUa3qY1hS3PFmd22PNBOHQkySvuDDcKwAvkVBR5Y7qv
qEkOzPttlyrt58xWomYS+d9oZEh2KktxM9Dq0bsdJyr2UKbXt/XOp4XbaCvCcKM5
w/8B8BTneyq0G2lEq7ZFggaKCeWpr4PImvTktSV3jy0dfhQXdHqNVftie4cgIVDO
GBEDL1l6xpo4TxRLdiVNG+5ATVTEKY+7k/PG1BTRJDbRR0bpABHTQf6oX4ijIgZt
aBpLO5mJJoCxdaMxvyauzNK39OgWkpARRDpqEj93XIrs5uWdZsEbRoa4MAmgDqTi
WBq8JgTcRpxtGt9XZtoyOynwI/yqxFBKvcdo+lhEpfMZ00HBz0OodRAoiaCL57kX
jP7xpA10SW5n0n9y+cWiA92ZPYfqbqk3vrFlLsVfQaa8EPoI6iZ505731PzEdiCZ
0d2Qxaqpxuc83WwpbZcDtvQw/J5Ftg8RbvawrpIGgf6Tx69LIw5jNkMfTBsLOJvW
X3rE4PKwmOAsqL0kWzUeDA0oxjncAE+1OO2OFH2UO+lgHmCL0pOY/kKBJuem8uxU
mnfWD9vs+MLLrhQo6WtTdEaI8eG3JnxQEAA1/vskEYXxllpkafeKKr4AlttgRLYC
3n80txcDPca1cb9Py7b+7/YSkd3b0xfNmB+7SkhPo5DXvYPaHf8d7KbxruoogL2s
6JwIxIFbEdm5qjpFgr6ss3AeqRTFbRHw8jx57lmo9y9DT21eA0OUmTWofBVLXaVb
cZuhmDpHbmVOk/xIyaXzlj5+Xq5VcSneWvGc2r/2tQ+Iv54HxfET/dafiHoRJXSF
Qty5OsfnmqG7cBNrQmlu+VG/3XDcE6Zlw3GLD9Dbi2ZUSXJxebrxQTsaELRc5Uvy
T4s488dckdIOT/IVIeh/5V5SC5xrvC6q177BAGsyFw8VgtfaRRuZYJ3T6Y2/JZ8l
LcCa18yjhiLIGPED5SJ9QKLLETcy7TY1GoCXfHS5HL5wv6dh22By4nLdQOsMfs4P
aO7MkPyIf6+yNYibmqu2Tdz0Xu75SZpmIdigqgNT3RgCH0/3rqcq8n2ZGggUbe8b
8jdXm7NcWz6JkJuy419Br4Eq+LW4EBxeGSM+je//+iSs++Kxktv2eW19ijGXBtlV
if2NPqTZ05zy9DN0nNnSWhQR3ZJqgoJQkb5NCmYutntlFtoMMr962TNOc+/d0Nn9
PTmVWkZD761NuqZ0ayumJdyw4G9yYhRMfbeIKUPAm56pg9HlCg3IA/nD8xZDTvgW
3ohLTgIgfZltV6oLlT9lBwezX6uqgldjn5DqfhIF1RbnDsDBvxYCK9jd1epFZ5YZ
83jZa/xlSCkv6OQD7BxagACplJZowaAvfExpEGrvzAuihMcIjVEvKdlY/LKuiOnp
gfrPKFraB3wG1tmAVG8t4ne7b2+5f42kj+zYhWdus1qoflnT4TRiAC/zw6haTp1b
nemwmmZwnbNiB7OcVVrVIljYonCqH0wwBUJwtlMvOouupbcaBs4D3J/MQ4QZwjrC
t3PdwQ6LggpbBjUSUduNBv4JW5Yt18SDNdRNcmRAonBipfAITpl3jQDvt2tCnd1D
umdmhM7w3NjxaoutN+PNrghiyDMx0pIqseTU34VmEb0NZ7z+MDYaVLBwJG1Dbjsa
SUZRGVK+6Jks7v5PXyrC7ZVLpd1UHw1keAUfdkJvIABgJJDpUGUjUwiE0sUfObxe
9LAoFja+nDYviXJC5Bz71bD+BR1/u4qRVgDp2Ow0TSOsqOj4kmRX7kbVy9dHwpyL
N0Vr/9HAaW7tSjmnbvNPbooE5+Wun1M45q1TZpsmlEo8nAk3QFjJjqBiXpu+ogAt
M3BCKRd01sE16g6Q64VwBFEvuSzzP312tPTeu4AbtWIrLEgwMGOQXL3g1bp+eRJq
OW5aF3j6ueqmVbB0SIqJxHmtFKz9SXN1XnwrKl/MBiisZLnXnemPOJLrt1qYgagO
qGgeWGRwI81xvJnr6YwJ5/8DRnlRsOsG/mqvbfkl9XKfe0b9Xew59//h9Hidn0fS
zPzuLDDdD7fmgReyLGbLLrBxeIE2TAHldCz/yM8uD7yee1uunsVpb5cyAHHUtvcP
Hus6lQqVsil+vMHn2gN7aB3QmteHl30UTWZMyVz2JwBm3CeC+v0M3h2sAmcxlRN6
8ay8AnwO0lury0ZF1gstjcP2AvR9X0dTdKGZBNNVt1P1ua2E4qZkVvwbR1C5/EGo
EMrKahETbsIDgAMtc7L30U3nFN93iQrujihvGj6MNo3jQKmDk1qe4GNJdIEhdtXu
RF/bXiUa4MFJTuk7KY5JZ6okDG8sBeWHzggWb9biY2CsaUCRNkdriUkuzWMKgW3t
B1JVxy/ahtMQPfNcXONPSP7FnyCqj9stByXnNP8rVkYEaeDMmOVhnjlBTpk525Nk
ENZZZahT91cq+eMNg3I75fJm79BEi7HcbOS7T5+w0LUVmbQh/3m3v8tv+GO65RqF
I26Qlc7nUoNmhJN49Z1eYUkcHeu0CiHN+65a5U6j9J7iCmzPNKaSpW+W0k7fP9ar
+Lkx0ABXrz8aMuxXHGULAdUh7wa0cfRbDjbb8lZ7m6y2XnzWPjQdYCxtc4ZF4f/O
dCiCHWCnYp5h41N9LrLAbi9KSkXVnHVnD0fjRLk8REilNgBKG2vuNcH+ekYjF5E2
zEt26lA9LVL40yYtnu/KMzpPmSnAgeKwvEbjwGL481Tn9AQN8q+vApezoD7e/yqx
zmhmsGHuf5SlXIpzD3sCkHuAiYdF0TQ/GM602eSPH320/buC+kpEQMerZ3fNFUVp
a1r7X5DX0aqmimSDmGTv+H5t+V7bYCGQ1RNO0Kpe7I89pfCu+1JhweeBsOfM/xPe
wG8HkYonzGjx9i8M8e1oeTaHOaWpLn3DvlW/U7bKwU/EDlmEk0UhfPhAl1VETjGa
Q2WBhiJOGP6CVTMYoT0BM0niP5XwAabI4uJTdTJnWOEe7llJUoNFGDwAkZrHAf3j
AkqdFs0UZqZz0mt9ZgIk7z1GNJ2IeYAu/DdOaq+tVtqZaL2CCJX3ybx0k/G1uGRu
m6hEv90xX2Dv/SbixrLtXeWUbhgx8HN349XIVuw0Yc5miHG0D3MgR2HasVYOisPn
DszWEV+xKeU34k35+v4wz/Ed6e5GnfrnKw/AiF/fmRSq1GMuMz0k1NBAOLPyK5z9
CUtSa10S4bOytzun6F9ykAjdW2UaS2Ga6glAZNvOWZSfGjn1CkjZF4fLlbhmA5Si
HI7+mLWXTfX8qSLeEWpae27IpvCfYJ1d1Cs59zCj2Sfz7z5fEoPrP2L8w93S8tMt
TiWBZ6hMkITLpODorVvLOtnAnf1csN3TYwjOeJQ0+WEPuxF+W2mdKGiINkITPpcw
rOjJ7EpFYyqibtlXJn+kAhJYaBROfKTkNuWn4fXxjAel2fTrUNEjOXtYD4h7NXEN
2xmwDOisJtuLi5EvsHI7kobO+qE2sU8Y/TYBJPILklnXhd7mupkbQJFS11fSIPhz
VomdGvSkS1YwxrbPuqRCN6/zBq2niMTCATxyhcyiZww2/skSGKjjjIqbJkNM2p6J
67dSxQdo6x6URKmHFCM+rOCseeERwRyEhCKSI0HDv4O+qKrvJk+UGRJPQdUyCLfi
hWN2hUKageVdGl62pehvDEhzE7W4vSvHpo4ocW3ANBm/yprwPemw6qLuZJXKRI8R
PAEL5+IeOexije9q8/ktSEVsJ55jMkL/hBQziHb2cCFttSphBFOx5sOkYYJw+nuM
mdQpXqagwjeuiKw0BXWTFzb3ytCLfSR0JylbmC7glszfBdeRVUx+07MqQP+LNNpF
iPHFJ5uhN3k0eU2R5C92bLlLEoC/lWMbzAg3P5u2Vbt2UedumZdrhnMfyxEYsY8+
REZh0qbBLvGNHJvMP+PJMI18XaEnh5AsS9yZraIwmYfelX86mJz4vdf1KH3TTCFZ
5j5d7bIAW/YpX6OtJJlLZreBP6tdBXx0CisIGA0Z9mXXPHGsjdspFjxp1qNKCQ0a
bTHnNbHiwhr7u3YgMsbKpXl047qC3o5n3WKh8OftzWId43iXseDE4gThM4Kh7/DQ
e+YL04VdsW+pptQ/94WA+GVaFGsOop96eeFTKPlqZo7rmS5LCWnuPaTfwGDvWV6f
Q1zoxgTz8CpPViSOWR012259WCa9Iw6tsoZypkzIvbDBXpcXhelsX0KsjGqCBNmj
uwW+TS1NoN40cay1yahjZu1XZtjB5YxpBdX2hm0xsW5oKPQSYE46Y04weYwI5oHu
wG87vY20EDgGepwM5Ooz++KPqO+xq0rPlITQ394Yq7iRFBsYJpUc3uZpDbXh5yBk
sARJIANQTKDChriHi3hk4eXzcP+L4HKvziU3oJ5wi7cbBLV58VYyID8LinCeLkTZ
KIkCd8T9Zm4CnnH7P1EtgtFrzX3aXNm90hKWxXbEgcia480AZEPtEwpS8lhpllK9
H6oN8xT8ndfdlFTmY1RW8c2O5eSN+harWfPHrNbepIeYldt8dfiaajlyzBDGqH4M
mBbVo0L3j86Lpj7Aru67JF9OKEqvIyt2G1QsVSuQIWXsGI0i+a3r1y8K50pNrhxg
Xmpq2a6AeZnOlENfAFbXi19kuQuvEJb+TH6DoDdZzAOeyBNBSLilRPnZDMOU7+8N
0VsjxXkMUmgg3383lA3M/hSc4RdsSoAecMgeZbWHKpSWX/0qP18w9AJHdeNB/MHJ
QVrgoF7OJg5340SPek0EuSRqlrtPmfvDzD3g+TfyB9UAMiB7dkyRNWVWjlmS2+j8
a4T7UOSKPWKG1C/XWDXG2Z/0/fm9TrAwN1kLisN1KSPL10mfMhRnesPuN//BWXXD
/o3jvGd1JD9x9vMe7zJomtv742YQ4kLK4Drc7+uI6Y+yve++uDOVj17vybcWR2nQ
ijFCTveaP/1xLvs2gWvfBSEjXCXWz0DaqV+knrw3bZ3HuiVBGceLGLVGktIL86rA
dKoTH6iJeUEGdFHWmseAmp5WYS03IqWz6BmmTe4Rla1/VCvDKsSeBmD0I/UeTczc
ldl9V/r6WYLI7vy99jJKcVhJy/wvYcgdhvC5VzMyfavq8ReheeGZfM3sv6j7z8ku
UoXJ+Q0SRG0Cc5MRW4SXv5u1Lfx7jDPp7yLnSeYk4By2cBxPiEqyWxrbinZi+iJz
ZgAkKdhm1ZpW6RKnND7opDBXU7q+yVQRRPpWsVyKCMEROWykcvwrW3zCHkP7ows5
TB0lUaX4eifvTc67bEscZ4qMYu0HPxaPg6eIjKgch1esFegiA2fjgwlGHKgR3h2T
t9lc/xoUtE9enhKPbLnt1m0630ptlycXmqXjoQgWkVk1uf2wWec8vkseSOV9kBYn
PkFhUmnFLO1IrIkCYa+R87tq/kUI7mp7uBi5wr/X3FNEY4qpJuPrPpTVKH3gkhwN
PbuWCjK2rkGadp4bknyJEjNLI1VwIsrONdZlpnsZoi0jhuxQS+PbBy0CbvMAC1Eq
FnSyyLwi4FiA+Hp7x+4WekDbGn1bXzKWT/t7R8kSlWiLHNJfIrEIYd9hrVcyugYY
CQP9vro8fjrO475rPI1swS8V64cIRwbBtNiJwtI3+mNutJ0AUa/RfwC2qhDc0/zC
ejj7ZVgRUPzzb1w4ymt4oL1czaOwnIfnwdWlPQhXkOuj/WSyzxBuPONnyZK9IJCY
BOTB5L1LQZb/yDjxRF6bxGbF29NQB3k5oPRwDlZsqy3vfbusfewLq6JvW+U4fuSk
yPx1Vmx+TnCe8oqzR4s97VQgnbR/b4J7vhxoZg+nqxXVsGGae+Ef8kRhC1NskgcK
SsKPXntVQ4kK/rZvw2B2rWaDX6LkLJ0RCGjgVhgY5r10sNK7NiH1qHkQq8bGh3mo
p+TR5zIMMB82w67LtaX+V7YaY9oEiZ7KT/tZ+OlULKbDdFMxes/AMu/+mMbRwlf4
yKB29r7ovL/s87kQF0BtOhGTuUPLvLAj6tv2ANxu7vPzYPd5hoFVwx72Z3vQxOXY
myz+i1Rs2m1dEoJ4XoGOLM/3rJMh8y3hYjL5fZJyB0zKeP/N9/iUvJ8ZR8j4DuRM
W/qoToeOcyADehEKRhmB4srIKNkzAv2f6VQ+ABnv750zFhU1yq7ojtfHg6UpoNkU
7ZLOs31epzykJuabTMCvuKwx6JkO2Jgw8zCaQUaQyXZwWTLaLNQRyC2HMQ0YeiBi
mM33WJh/9eFfsDC695QjkdQxINLZDmIQtfcPWcH+heFGOR4yf3Wr6GSsbkPOcuvl
/WlyktPDh+QKI4vzQjJHL9NJZ05SqBp6/LlyebKf878N8Zv++yXz7osIZnuv6KB6
2qg16C/cDaozM+Uh36nl05cfVgdWFhJGMu/WdgSym0bd04/DLLZEL8y085FF63Hx
oHpctYv2xSEBwrnQbDmZVWPcmaZPZ8Arblt+V8+CtzQXg50Yd+2RqOpL7eOUwe8o
i3pgVyBAieueL6txp34c2i/lhg/HzZqX4kpLNF34Sy3+8CeMGLgIU1tlMXERMxdE
3dNTsoZGlyDTG9rUuq77ZV/iwSxeKVMs0aDXpv2zRf4ccyhFPYe1tWeQlgjn04uk
51mZn63fOWN+KV05PO9PG5yfO1um2imeh5/4/SEoPD0LiG1bz2vwNWcE3K/2KbuK
ocaF3LaDh5KniCtbUqEnWZQmYQncSEKbpiGB2wEbSM34oiMjjXAIlsSregBKSRdv
6Qyr+CfaiCT0x/zC+mw169TEOweypVpgICPcwNR/A2SSzp521eoMNfHR0qk5jR63
KKIiJvKzMJqyTXblNrMO9xWDHuBPBiouzizkDM6Kc335gcTCU3Su+Nz/qVMJNwx8
XlMopNAz2nwOceAhCIs+9f8GprlvsZe1UcJJzNUu1xfCdN9VWLHHhmYA3KDDlVuf
tk08MiQoMaVrpWsO6XKkH/D32AsBBwOtqd0ohAVPEEI2uAwMBabDJ5uue+CWPghQ
a8DApa84/97HLVmHQnkXmyiTtYFxurKjTwpsmti5oApJ8qaDhzk+pQh/ap5i7/qF
RM99zqUrvS69silDYPXhM57hpnEoTFgv1X93jWewS2S6JSJkPwEBYzrShuHvN61n
ATFPmvGygvWaM/EmgIWPibECQzFpiu3UHUx05gv+TQMAbeSP1bnvGICmEjxJPir3
dyIb/1508lxUJyqka886N5NB0WQQv2yCVevQ9SubSBm5nKOytfV/iaLXRDSL6OAq
DSrSOsTQ9+GjXDu1OyqOjrOK/gL6BiJkw8R8x+ZnBSZJwVw7V9JnwMzp8XRKVCZn
Mfy7kLZSMIWgd35b+feDpktqBjJaRFjYPQKlUl5TRgKsxzE/07lzQnnTTy/WtCDi
1NLS1JwWxEVA0WK69IFsbmznix+Desl1E06US3WPM0JZFl8kXAnJsWAj0W3XppSH
MUR1TfstUSIojUclZlPqS0iIbzcZaui3qlvm6yIMXIM34G+NCX1ZYYl0Uz4TLuAt
TWlru80F3Vv7ZfP7ILN7q2o8BqVYzQ6J/G8yb2NwUvUE1U+AqEuDn0s5XBU3bjns
W7YcUzTALH3/PfHKJk2L0QBzcPJXepHq7uxHQIOtxxftkBA0T5nNkqXMmvrFhf+E
1Fgt6lgOaPCL4yf2jjSvnMMzF2m49ODAY89oUO9in5m26sUIvPwpWO5gL54Y2jEZ
1UGNC5Q8fJH2so5wPfWLzIXfjDcQlW+9N7UaP85gR91wWMpWOpdJxei64Rn754aC
61slBfpRtTIsTiqUgjhBvagCFpCMFQxO8iP9TmpoZ8DmG1vz1vibxzQBk4H88XE7
KuCNc5TIfKWwXYd8xubEW4W1wBvYh3F+jAJDj5vz9rnq465/QdG185u72ycGK6wR
/U33kfZMCrBFHShRvrnkBDTxFMUMr0ji31Kn9PtTMX9QTm9uzF/971ijWqVQk/yL
5bOfLsv2d5UQXxlpI8q2oQ2DD8DbXgwXZI7JWZa7vxpOho54Z1WrzO/j7g9/APOU
Q5icyJrUYBTyXIGSiMi4D9XAYy8eXKgLgnLKwaeQvmUbRy0alIhxpKxsKEo05K/u
P7qLNLafgwNf4xOkfTzQOCYQpPTOPBJ5VkxCcEhcT9kh3JT5xHC7/eUqzuDn21Fl
M5nGmDmCwcKhQz/TvXloJMwvUt0M6BhmHTAaqPSQmpIEpyF+kkvzfVVX6f2x5EE2
OGAWT7Gt+f8EUJGk3abxzI/13x9eFQug9ayYhNstrwGGBxfjXpuZhJMelGTnnqay
+nug4dH3PwEyEswqqEf+lOzy4qdzuvS4hNfFADr5dPgX7OTFrnjx+YZp0/1S0pKg
hAps2BTqSNY1Pmxo1a2YUSM90wRbEvAXgBIiA+7Q5ZJz+q6fZb1aoQU3c/4pDQWE
qqH3aZaT+UBSc4kKECYajvLcY0s7uPHh5i4aEfz+QFT8vxlpwYODle1jK14mif78
DhPF3jIUzWFT9deTEgTDX6XHvyytRfDLsu7fm5pvlQoIJ7QLVrsn5M4q/SG2k4a5
8nu+/dPQdaLWgXuRM/B4DbaVICmkWeWJEU401Dvp4JzJjeh/p79TYUdNoJE/ZjRx
7brtApNZCCwpOiGxSohTwBFNBuKG3p/J46dfw5t5toe5bayr4N2d71Z50lTNU4Pw
7PsE83mp9RM3tZ0NMHrNc6rvSHQB94/mD8QS1rSgjgeJ7R3M5A/8n+Ur04bYVtwG
cC/OzF3SwmFW7XvpC0uKUlnhirakJk9s05/r4W4rXQJ6qijwiH9J9/Sy48FKvhKj
6zNizn4cUrfJ++I7Jue0Zk043aH5OsxjOYDKibJkWR7GP9utGzr2t14jwWg2QBf+
8kDRVVUJBsd3qa0y0aVrBIBW/NNqDpiM5sb39GKHka+y9k+0LFrzJVFqhsrVZdOm
qMWJzrej/hYsHoE8OhmHKiApqy4G1OQ8CD1ewRrVU1kz2YZiBW7+yflsuacid6dv
QFaAMzKVtIjbdShC2m7z3O9WaDou+RK3IsqVc+S+yLYELYlmnvzE+DwSJJHvULiC
jdLnobosNSxOYS9rVTf+CzlwoYVkufrq+ElQyQqkNK3Cvh2TIQsT3vibjr/tqWzz
NUB/p+kFCNbasQiuRELQqZVARG1vY7MHhkAXyMT58J9cR7ld0yf+4CzBbz2CBsXF
a7sIeGCvqQzsf4LKfoup1p3QukZbwEb3mRoTi9QAckbDv+GxcsbpLLuQDYS8P6X6
Hm82sTENi/xWL1+hilGoHEUH8TbL+HUGH2HSNcI0tztDdbqiu3xJnOd1LQKmu5P1
7tLepmPzyqqy7658JwBli1O18PmBIh0QxwEO/EWO5PNAbqWozxGfBeOnoENR2g30
RjSv3RkpB6slxYE7MqivjGELSbS4WLQRmOgZV0FhFvR/FRlVaBNrVbgQjQ/r8XJk
MvV59KwcUOi7EMr7GQBB9lHF8CfToExSSRFIIpM4k9IdZPvAIVWo7iH+QizoMyOF
8FB3vA+B5Xd7j7uHOQa8ZiXmeRvZc5I/Eeav0LG8ASowTc3UiYrpI+iFUQDOUtFv
5kj7vROfpgIKduizT55HktXhKPQV7VWdiVOAb5ZgG9D9zhE3QqRZHyyIlBCDnlPe
3yqD63MdhGjFxxeVL3YvTKGi2veL6dnJ0wIstJBMG/a5irYtB/ydFP0Mt9Gwg5Jk
aeJHAFrE7JgnQV0B22O2rabMMFGSBD6EQO4tSQx4ig5e2BaT0rEqO5jPYy1kMLPK
qnKII65c0PL84wqr2qp0u/wmp9GqZxSQ+Yq2lsiSt/BodT9oBt+0i0wI6dMENy3m
5Z3hg6ag5bQ1FBSBo/bcKKjtJkOape/YXDTSnpRXoaxsdkzKueufSG6gbE3QC1JD
C2J9qccVj0wBhQ5XvA2efOm1F9ybix9y6BMCqrLbI3zqYohtD0LrHB40uSidg3Nk
D4rZJLuTHqDaXcMjU/G6mrbDXjsLe6loeTN53JSRTVrUhHuil1CzfmHrkwOMBr4q
2/48bATyHdpnmQyxABV4bHyi9e/v6PDiycMN8pTK+NVDmyPGxgJnp9caDYLrj1Gf
ugEvad1GguO/vLtAiI5IXssFPsKMqDJLOom7+OEsXDUMbxNL+BupOPjFC0v4zlkK
/pQJDuSWL7NKZ6w+UNj+/dFc1uB5jkOW2069/N8/ieJlK0xz2OlW7Syl2uPzXCY7
vpSdHjjqbrlw2mfFZEusjhw1E1Qf1ZWymvOXCgzo3wYnPumx31h02oedZdrpt9+S
9yXpYVVMVgBtCPuEjmuu7KXAXJ06AM0dzbwJGlcTm7DkiK2Mw74sKBQnXZTa2SG/
MlKijVLZEr2Uef2dJz9/NBHrQn2CPHVR7X7S0CAHBVYIMEzyKpZZlK7jHh4VnMoF
HIww388yKY9iHc/lXNnOF2Sm1O+vAgUEygqKabDEmQ8BVqOLjNx1U4dufjXxAiuq
mR1ADnS7ziL9S/WSO7kaldITio0dQkCudxfxQMDkZvAfsOHQ7S836zGxyYgcSTqB
MJBjASZe/wmuKvWtMwzQ4D/jZo+Sm7GGTqwhrixzGiI1xHw9EHmaIbUmNLt6Xok/
AGqyxCoDRFsearu+umc7n7imCIay21cfFgjH4MFjB0kyimMsaV+/+2uE5RD43sU1
jOZFZt19JDyau1kOUlJwRzHBKHmcuUNIoHQNmvIwjdjBk5szAxo9KIQVuVNnOyO0
zcqhkoiHs52A+fnnLAQoKLivhok2e6H/orK7ma9hVadxMz7TwZny0fTIvDORUNks
9fgQEvhr/mkSglkfo1dBpuBEx5sDSBPApghKsszkcP1Nu3TTWB6aB/B5uRBVcT6/
qiN1cDL7lmAh3WlB0TqBxSUKK4wsaUNTR/GQw5GQ54xkXrCqKxvw4XbV5+N+YBxz
ENyy/AAXPwB/hEZaMfqrAACFqYN7Iqaqs53vCzQYBpkQhNZpvt0yjlB5qAQv0nSs
93PCfygx20ijdDKu29jWaZrOQ8VZkmBwYP0z/h3/IauGI12Kr6HIENlJRtjwrzyF
7b+wpAot6Or7WVJ7AFqwlLq4SmAh+6kEG6er02Q7UkUopq9GOVBczpNWJqnQJM25
W1UshuqORtBOtBi8HyMJh7DwhYIy5UQaBGObVIg7WObmYErOq8840tNjEsweB1sh
yCWq9Kbun5+agxeT2zGXsWz/jCXmrWUjp9spuzkJYjv0fz8ZcPNFVN1NfstDkOKu
ub/efxBeDAYNbLJZjlTFRd5t1KiZ6AneY17JhTiwVcw9a+SxDVJUi2IGokKUsJ03
wmPOOHEcn4Ti146KdhRvfGsNqQ6Xkv/nEeqJda7tGBrbPFtYFQ0IcFEQ1jSJuCPd
KECNrmEspz1cce8qQKJ27KGDyxp5z+qa6xVQyfYxS3AvC8bmmaEyzQwFBSF9aezS
yvXTHPpYKzUeWmF6JEituWe8Jtu9OX/X26saZoYeNhQCy99nVO+cIH/B8y3x3sfB
5sSyPiBNJ36izS17nX8jsQdoX1r/+demAcfU7WbP5tQbzqbSdpFYOOM0UYNXEH3w
cIHABIrrfUWxQVFtXiW9mXTs1HK5gbBae3A2hzJ7l014rn0znm7CjpfMthn65IiM
iNkHAT3Aoys0+AxsQ9m0rNh/DXgf8NmOxlXS119i+oArEgYYqAn1AKiD3+mdio4U
PukMfbUuR7D0q5vLsNN3ZObiYwHbDyrjEy1xYXRhWmmLPzGcTqo5s6t71WXJgEvu
LHZjMhh1+bmt5leTKF/GZ8efWgDZRU9untZseCTlss/SfddZpae6zX0n6hN6oWR9
Jww6N3due/oe522LmDZJNkDM40M9TM9Zf161lrfRc08+BxQLFyjWV3m28vNzbj0+
9nAyURLvLqbDhu7FrNHBu9UfBKZ5VpdBG+O7FUKGTyCjtCXELnt6B7PBpQHTk7ks
QgiIsZAaIqDy9vJ6k1sGBLT+XGMDchgdk6foqfNdg6vfeIfXW030HM1XB3y3T2D+
6C2HrBn5pigom2Jdtf0OoOvJXYuczeh1x+LXZ/u8BHnUNYr8GZ75m2PkO0C+4srm
0C0YwRmxy5v4wa4+mliAO9YIAcdBAQ7v+r3QXNfQ8U9rFx2aj35/PL+XCRyWqanG
K23d9d6RQd0g1fZ7aV+Z4F/tfq2/UT2YdNYv2RXpUOk0gb4msGO2lyNWSw/VOwWx
ZNNL5QV6d0nGMMxeacFE7SxaoMLkluH0+EIQHFTZxtSHR/ghFvBfUqMbOB6LkO5I
CQBnEG6eL/VaSZtJhYFjf1s8rrs6dtr8OAXkU2LUY5157+eTVqEc0cPRLB1FmBlJ
Sre/xebMiBzf+9/v7weLuA0YNhxXSYBY4EVxmu6Kmn7VwJhA/cuRhfDzsfOQ2HmB
BOnVDxMB0/HtT6nrGKEVx+APGHHm/+Tpm+TmJ+cRA3hm/OL3dIlNIj3fNg5LJqPi
jWWoAEwp4cpiemD7/Hfx88UJUCATXZn4Lokeu9oi6jVopkfkexCix47mTYpSV43P
Uw6NdGt4oQMCJ9rU2x5ktHr1uDI3QMUR/58yvTrqCiJndoKoadYES5Pgyki/S0Fa
eyrZMf04n4Hd42C6FK2VcR/r9iUltnbsw9IwcNMwSVbNkF+l/TBefsTzCOV4EVNW
4tmqcPSNPLT2i8N0vsLtvI71Rj+mhqOpO6e8cqBKc3H2OzWz/N7OZaxq6lZ3wSYw
yk+YhtmLq+oiMudip5mqBjfqxy7RBlCphrd5e4Ki7AMGfvZlnsqw6VjHilwAafqd
3AXvG49jbopGbXJM2l2BmypDk24+zSjL6lqO8gSC7aalgWjmZYWo8MXEHK4A0ZKV
1paXyPGtzXCeBeyLbJtPWY2bqLKXfmvulK1rYD1/lvVCVbDON5bBD7eyqKATcv3B
q+9hyj3SPIElp+NOZ+3wyZyF5t2dNe4kAs/91XHH/uNup7ecTLKimJIdx9rh7aUf
GqZXhBdw7qAB1hPOJfj/myFzh5SNl68HdH9tItSeh1HooSEqmwaVaFCvIZgiQHH2
3ckJP8SVaI927YTKB/lma0w+3udIkBoHKRIpWETSZ9Rua6aa6ZgNluR06yproUSW
4phhIiQU9xvcHlLvuMKWxuYn0zy+xwvpTzOHAfgvXQ51ACywG/a8r93gm4i3xTf5
QkStjG5uST1lMwbaktXNpr8m0hwEzIGR42Ke3qScwI41sJVlR4DO2fHGAzkk2Hvn
pSNSQGgr4Rnyj5TPXIFVoYEZymtIdRnOTgJs/sdlUTlm7J8i9GLMY57n6gODnd65
pLqTD+e6makZVaKm6Ihh8K7T1Nb8eLKWxhwbEvdVNW1Bjgldcv62E22aGeGKoE0k
fKgK43J44CpCvgu4FmqEPXUgAb/CkXJbf6vwhSWWoEh3xX+Rd+59NgE8h9a8PKay
cRzeK+xOT3NYkpDAhtvZXqeD2J+ywb43SkfyWxm38y0G/epO9eeBiQ8f24QxeKnd
r9F9ukIEozhud9cIHbTXqWaj2ibpAbNNRtrPbbqXvRPwSwnFLOSuR7LltiPzxG9+
RjxHLmIhJAqwr8Wkz7mBlMr3jc+riTONhArJSm6QAYIpphJir+5deNvj+XMQ95ao
O1/P54FRW80lc1GMtnhlodKmTSrimWa8pXxapNBbHtIH9mgHO8p0R2N5hUIPKNGU
h4o/mXqCC2Bd8bCTaI2KzmnxPXrjN/SYdW709xrfI3wzOdO3ftLyDfaFBisDsFAP
zeJp095IVVtgVScdlynkCE9xtjv5cg5DlOm8wf5VxVnOJJM10NhGuc4Dxn20Tt3u
JMdrzSKhsUEcBPaenvI/ipxv+KHeu8aRZVfX8fssjoQ4w0s+yx9M0JjnkH/Ovcft
b53jBl8Q9LrPr8ERmHX1x8Kb4XqvwbXRwvLmIeYqVH35wS2SmFLN2HCHzfHDcU9R
8rOUhq+bwm0qQ7GhcwLd79b1F8eDVZAH8BcgyO35//NU5XeK6EhtNdZzo0c0cg5W
Xl9v/FdG3qoGpCWZd4l8hWuy8XgSypmm6OaJm/VGLS5rN+3WFi2Ds633DVP6emjL
1H8ghDNhFbH1IglhP0Fd19pwI2UxKCZiIvSYKvvV29elS6HrCZRc2J0n0SOgLNCP
qVnFkIJBejwinaLmCaPxKCzmUvbDwXWjEVQlzKwGtVv01QM9k2WyKpAR8mRbPK3v
wU3qkLgXB+0IZ+GCbNBuRZJyJ6c4hQvgZl/+9+I8xcxRYULiMzODTvcTp5Zg58Uv
Ek7XhSQsLyMRxN1gpfkft+fScdzvrng0bOoHQ5ut/erBAuTfjMaO0FWl61MUcWZH
FBXKh57Stab93ddXVEhbUPdXdDZA5f7ts3d7UFBh5pl2B9BnxjuXd6YSf8rHdVbM
A56rR9o+M4fYGxuig7OO2IGg7fGLf93oeuBdANFZvP9sVdzadGNYaoJ5vZtSZ0tc
rJydMdlKxEITaculBI+HyqYkLOkN7xO4CJDZWduW83AhK0IfHtF649gbxJ08OXXx
xmndP2crpn582rMGI5iN5fYQ4pYC/D5S2lU8QK1+2ReTcCkKX527BcQDFwMjKrT8
JiXV5842OtPmnBPcOAzA6sZCMf/fBjJbXpQgfrvvxgpU/vnhHxyrMER9ZtxXw80e
8Y4EkxaaH0CTFC0Fj4UsrJPW+DY+eWwJdhQz8mwWUOtF+lnMpjGg/G4/KDyc89M9
VY76rBMImjt55W+pyyTCmyOVon2/37hcxyDn8vqe22bM/5FhgyVOx/ztiPNTVovJ
IrOVjAonn80wMISgzbDHMn/MO5nTyz1zJ7ABeGqtC5Z6Qi/WL4EzZNprmPotvpZw
vZTSh2wSw+G4zlenMh5hfGbf53gMeYvhOYZrgkxKtnBIHhFx7ag/92qyphJjUDeL
Axz+OfwO/AH2YBQk8UrM8NzJCF1z/52eO0EEMauzkz3cn8kJQ6uwNjadnjKiirTd
h8U7g3QlVRut5Ff2G3zHJ7L65h0ebsV/0tv7SrsG0aXs8/SMJE1eHZWm7fvEcFaa
e4d42xdH5V572RgP/lHMASwtZaoO/IJGqoN2B1FBL7n8nT4NQQRjuRWy755fHT1I
nftOel6qDGt5V5scvZ9LRNzggUzkixRsS/+6qX19z2m4AHdCR/qju9ixdqq3qrWb
1yAMYygn9+PM28Ivlbqmn89MQGRVsGVqKsoJvUIIVf9O4s52Rha7lYTD7ZHdaM5p
7s+75z9VNWMQifLECBrIArHTf+eJ1O7EXHRQpwHzxDeoAwjFZqD/S57CLF6wuRK0
eIb/Hv3Di7ls7gogR7AFW0WPmDmrXdmhmvgBB1JWWA9I3aZIWEig9piclGtpu+0w
nXbyDMIoTZaPZkDVMMy4GKxn5ABGJ41Bc7mDViA656tnXM6zdRT6hmnylts6WGqa
jfINHWzY5/YYTC9egwDzviXFq31PxuVcj6Enzdo2oM2RwJ/PwKm9unZQ+W+lG8+r
GINjFOxTnmhPh0Jay4VFzIHPJOpR9uuB2w+8a9hgjPhm/Ahbhq8Lm7hXvKIiygCq
40/aVDsbkoD5xajx5sys90Udp0L2aP4sWqXnwCUFKIqoR//Wq/r/2puXzCnh6aVx
oxKZwVRZBI6lpKN7P6pHhnf9v8S7fWenEaE1LCpsJc84ZcH6K+ppOyaJhwyj2ThE
VGLYlgwt4LC5Y3SjXc/mAizSj0t2sjwnvCJfS+HfTTE=
`protect END_PROTECTED
