`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cbNob0DZC7awBLgxNimnNuNyylZeZ3w+Bs49A9zPV4PnHGRmFyJS8q5CeHoCA/Mv
9K92q7ecaHaNx/eQ4re0ITnUw/IrbEFAegnBeIp/DY7t+7As/0yUzMmLoRO59uog
iBOmI3aZD+8YwmSIhwMo58c9MZx/0JCZd4rq0eefYbAfFOIKeehTq3nflsGNsrbr
aC3CI402pI6ub8ZQscMq10MiCdn0K3fo1w2B2+xDNEG/x4bDoISAIGC3GUKkcb+Z
uay2Ci5vy7EwoZdWP5Zd7r9iXD6skc8IPyxjbIyZuwdfQHgtyV2ipTTRlCPfiNlQ
pU2S75zUunEUCjv873bPT5vUH4cg2Xd2BugWnVLA3Sac6dUXvT5f/T3SZGBb5tN7
a9mm1E+ZU11cVH3r9bKNaZd+wHfAVckTmOBL0+T7suhTjdO1Kk1phuFsEYLB0jY9
A/7FZvir6dOUq5zCEHl9IgFpKhsSaS4BTrBQS3Hlw/l5ZG9G5+c+wKJxmLHBFF4E
VzGuMztHkJTCbMA+rHWkARK2cC0HiqlBw3y7itvus18Nx8FxrHHmF9UBb4AVt3Vy
6eS41lqj+zzNOo9ZD8YMUd6nzUtHf0EximRsgMLNkE4=
`protect END_PROTECTED
