`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dS/JjSzzbjuhjYZuzRpnxZ7nnswvwgrg7ghr5R/iyyTMyJBf/GhPZhfNhjHFAmS1
wG+paWgyvM9cI6xhEUkIf/6OFnZcX1aoGb8TX3Qdly+UjNJUU3fauMnETFvqZAPO
oQ+KLVVuoAl75qFswhPrm90KRyOEzpl+hFf6/rkdK4mkiadbT6IL6yJxnRkn9KRE
u3U1YLGeQ8gZ56DBadbpntUlQ64DtrFM9lepIJDtaBpWkkqD/Cd0kRaToMywkJIE
ONgGkE4kVjqvP40DsP0GN0uPXJ4SchEisbpsCBgZNAyPS6PjA3voUI6swYMg5Qyb
9s4YiSYOVYbVlkamV4wAR83slb+yuXIro7AoD3jYkDwUAmIGuu4qiGDTmo7L5e2Y
ZCwiiJSESS5i32+GZJiT5siB4crc0qBF8sJV+3dxgn2J44nV1aswFMgBJFrtDMH5
yerqV0Os4+v8if65AefgYg554zpAjNh9H00Ley3YSJlfADfo9BUeTdeym9tioheu
n8+U17yxqRZ8bhQH/fRyo8nlWKSsDEAwvV3BSEJKt6LXEn/a6zFnIvKNxC+yB2+l
OoOjm1jvh6SoeI636AimJI1NxYK3ZIlppaiPc/r/HTsOIQeyQfZqjXG9G1Ipcp/F
9kcpO8ZkTkfneGyizuA2VFUE0T8vsyDUzPf+tD4QhKusy2G46d63kuH/zMKC7ZVb
lrPrVJtt+RKRwv0IBY4bgQTXh/VwHgzUCuEzKnfMrsInH7puX2286Vef+IjIH2fE
1AqAxmnze0mvmNWuiLbpT+uVj6puhg9eAJGdf5jDQkCNosPSKuGkElZfrz6nvsyQ
25YaDYr4A8NDDbqsKZ6Xdi1+B9bVv7DhTzpJ5nUyLpZVWyp/3i9LqkUz67V+3qEg
8aH9G9X21v46uW/QCmS4LKWhFvId0TGiIy6DQMkuzYHacebqoHo6LVz9dseXfaX5
6dHJ2eRptMrFpdrNgx+J2Qtd59z1/qDdHCP6sD/oYjhQBtqMzx0AYwiRarHrJKpS
NLQE+iO8IlHmOQC+ZEOBx5noPO++2UaFCgeVutNLzCFzRIWoeqr+E0zKhOf4merk
`protect END_PROTECTED
