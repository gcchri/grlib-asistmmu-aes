`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kq6a6Im40eU3Ffgh5j51KowU3y9V42f6jiFVWH6mnue21dZd9USu1ciMUOrWSeG6
irPOz+RIantR0TculyqAWL+BoPsgBCQ5TeaSYTH/QxHXZc8NL7tMdC0hxeEmKYuO
qjQNWWiFFWVSCPa0iI6NF3D1SmadnoX4Z1DmR3+f66virsO0AWGOirHpVRQaSk6h
fkzchIMTZixPJpkpQRWGJjKzhg9tYwwJulGB19bAA7YW4H8JQE1fnjLpdCqh0rgM
EMbJsW8nQw4n+SFN6pMGYY3lBAPn2vTjAVZZ0zlmTW9gBJC09Ge+bL1/wkzcDqkE
94UECvxxLPrlr8w5cPvCM4Yw9lEe2beXtULpfeLVQSrd8pwn/++A+KHv59ciJ3Je
O8AU1dXuFGNWcFs3ZOi7wh5YCgEXMm4FAiOzv8bT5z0gv6AUkU87QkvQEDcbslLp
PF2mcAOxkf+iqEksoOBUEV1XRy33PvgBZo5d2Hl1NfBkNV92Dm2IdY/FMaMr23oy
Wgx1vjkSfLac2EHZ091xek2ku5XiXpctiwAWXQzZ110LgizIz0ZrI2Mx25anmoLL
ikXLNRyWzLt0AE5gWauVVDqsyIr039KzQ7QNVUM8LWaf0sWKu31+F0ezClVVXn7/
TECHVN3ownSTvzw/znnP8oFl4zCpd2zzue6amnyZsK6IiFh1sARKTbYmK8lsd4lb
GJkR9JlCg0A2lpXNAWyvifRiyLGRBjbUoquv8awG1Jt1Gf3WSMVnknJmnYUHhX/x
awVQzLW7lRFM4lK4rfb4PYipL861+opus1iQodxUfS/ZnGnIfLPE/mA/lOY7rGD1
GBiZaW2JNhim6PcqJqRix39iA1zIDQQS3wzDTicVXvq/33Kn7y+GSR5hsT16YprE
qp/VChiQJg3YYLXKKddaKS00n8v77onQWDEH8GahQcYFy+2OZcGSDHR8mWKCjpGk
KvsF7GAh0CdhxHvdmjDW0rPnaD8IMu7WbkHPdImetK0eiRc0NDXo1O8h0zstbTlS
TOd0r+SbH3kf4KDBHwiQLjthZe2TvY/sej5nnQcJmY2XI6w0yvW8sLkRZ1XNv+u4
nA3uwoU6PE58BJiradu5nyxCKodnsrrLvJ5AK+3fnAkApZ4rpFULRQ+IbqT09vPU
05+8OB07vYkUIM1TvJLyZtP7lWKAWmWaswqDYJJTHPrHN7GI3pYrFQ38frDrnMY5
Ua042/GSulHf1dbTjilKM35483Bz9FCGxM61Y6Ga5djgM0hjSDFZnnV38aczb9aq
wJFSyPlibQFGLnYTPtQeCI8U1TjG72H1YO8AQ5ovNFqOvE60xEv2TGuQwudZsfw7
O0ItgOCKMUmu1lN4pk4aUublxNIs6YOfzxK9dFAsRMQbJw1fDA+wtxmq0hFHk3X3
rH75WyoXXjsGQS4dHlo2TCvsFYlyG51RgieNc8N6qyy0r83SSMFz1jPmhNIWJCyW
xWvdI3tupo3lx9eK3mTUYDjrdCM26A9eqrRif7dpPL2k4cmpjjgBhTvANHp/0o6D
O6CvVNe13KZN+pKNCcsaays7V3V0Ei277Uzx67oG3YPozEiZOqlMOeL21JkjUBkK
dbt3GtkPA1JwNs0ahwaAKG0IM8XEL2l06eOtWbOIZE7FhDBkNEhTIwgz+cpQZ2Z9
6R9qCiBYqJ32oO0JE8iZATFG6+SpKX/jsoi4FMlzPaFOlIJMrrtw7AbYhFfqBojN
NFTSXNE/WX5wqODcQFurvw==
`protect END_PROTECTED
