`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TBVfOMKNGt3eeq5SCSHEsPjI1Ba3+lsXrzyRuCWMzcUJQnygndaJUkaSJQv+p+dV
rGDLvZvSGGER21wam0FFkoCEIDFR9LK61AlEJfrthoaMw+2phGmwvjgKrUYTGqTL
gjfp6Sfea1hdkJ5qR6oMyfcgfZwEaCerxK2V5+5Ll5z0ZW7FLtNAViGlLVFx5hl5
o7wdqaLw8OuoDiW+mfukCyJnvOJ182y1ax7FHs+1lhTPiUnlnxDse/F4QZMXSROt
IV9JssGupgXTSbiRJ6bXyMGd5+/pUXDzrJcJT9sAL1WBD0P27uAarNqpL3sXVZWV
8/QHtTUkpn9WkwueeBzrWrIB/ugPdeo4jV63ZrgSGyFiwM4l7io9Xwj0trRWAc6f
8f7RgMR324sgYWBKqGoI+AFgD0UFRhJFZfAnjXEkqdJMAlEbl+4vbi32VITNHf1+
JuHG3xOPplxzcYaWcJ3x8Gttv01Ck9vVKjvgiP26sgLBbtDUsfgHDdCwMg66NaJQ
chlSRtPLmlUABApcTtvUnaAUuqqGX/TLekdfYUpiPXOKeGmaJfdsHZMbXo3SjD/r
DzsFFyXNLFKwotuaFbkvAes+kNrWdns4+zaIHXA5Drq8r1cN8ZG1OAtAqCdFXrck
i83/5zNKeSsbAw7v6Nj7pgsPz36TJIXxyP2WSzrYw8Afdk8P9EnkFyXGYW8U+rTP
IRRZn0dEyvBs8qVdUrDAtRmAx0xUkq26yEqNeS1u0vIqnKa+0Tw2+WSrCltf3SFi
2mFN/AnyhIoQrKjZNwBhgawC/R7VbqYqGROAXlZd7NruLdkhAPRWenDDT+wrzYob
f4IxPaw+AGNeIMGNGAu9sqvBERnGGZzN6a0Iiw4NFeKe9Z8zbPemJz9tknYCvkrA
TaKGIGiSPTU9mXLZs3H5Mov+eijp6phd/X1PGxFNr1Fv83Vt8WDAfhTqv+4+ixK4
`protect END_PROTECTED
