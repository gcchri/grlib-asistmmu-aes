`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EuNDwtJjNZjFUPD5whmQvAq98MxE7Eed4n66Pg+PIbILKJS4vU57Fk2ps7kilY+M
spdX/pl9YJ+enN+MvHZQ+hYFuZkDe0TC7HIXkNSO5Z3JnvVk1E47wXry1lkfw1UH
+l54AxX7erRr6KWfJYIK+96PtG+01Dw5ZQV/y9/D//rAaUmQ+vdbHKhb/lRXSuBS
lb8yWd+sX4l+6Z/O1HVsGVmqAUkX1GaFlYKg82P0Z9OPu4JjKsvHbTHdzOugLByE
R9I24QeIrlJgVKerbp0g4gLIVarkXYl2WFZAx3avcOuaduowsGzMdOcEBbka0piQ
NZQTgmvETM/R8gAWqGwLSiu1bP8ZxTNoT88+buqa5LYD/CUuxb1cWMH7/ZZZTZH1
hj3c7afoOuglW86ZD9z6vlIxW0hhTEvWfk82lislhmFUHVKTWjB+jHWv5BeqH0AJ
Zj92zrXNjUgnLgysIG7LwVG1rQqpPb3v6E+H0hWY6E7pEoZZm3Gf8yDB9ws6qG+P
7BjPK1YfMThJCVQ4vKBRHGlwb/Ry8jZrgWCzREdi2QXMdGU7Cv/A25zoWnhYIQXl
LCXrH8SCCpqQik/MEF3VsLPIietB8RrzInt8Vd2GRh2OFY+LSQm50mNMkgF8H+zm
o9w9l3XhHCFdXSDaicVauMGzj/sSGFA2xylINYLcxQnYAT6vsru/fX0aMEaNB/dY
vwIxEC2DBOC84ZwYV+Fv0ryBwVF+/r89eDAoQUGjYqSYpJdeDOfiQWqsM26Kauyz
0PEWNrXHXiVS3G+CY1NREv1T3wWflxWejFCcad1XwvolrQWzr0q1oheFAvHLaapX
rAv6Ops1MCg5zkx0u83v7cy/XmF73ymsF7/rwhMc1RwnMwVZWp/U9tYYWYuugQQA
EMybbAkGvspTzSqeJHDuG0W+zBrFJOLJUcnAoa59wNufif7mjDk+zHX0Wsz9ke3C
wsYmHTHP5HBGDzApNpErv36/VFB0ow534P3Vthc37UlP8n41pZpqcabM+N7hT+rO
sLXV7h4Bqfsesn/ByYSxIX9ZkmKN9qHyDUtv8AUId9Wwo2UZVdlX7r4vG1N+2wEn
NbeiDGfIwckacwyaXkJ3pjznNGzNAGUPEslJzcpkcQYn5Jydzkm5r6rBKz1FTbtM
70czcD+EFm9JIpEvcNexSJqGwtvG9THD/bIAu6nkC3EsQ1bMUPPfiujuf5iVxXFb
HpdE3cp0vTG6cWo9i7IrEihTa4bmzPYhXiBBG/oogigikHC4Ol5S0nzvQlEOljQO
Wkl6aGJk+IhFoeRDKr2XMnAcROuaKd0djKy3WYqYLjh33Z615cMbnsCE9xiumr1t
7plPt6OT7otN6xxIJC82kadN23KFTbjNJB0IzXxtSohw4wvnp9LyoK9yQKq1ZG63
LYe2373mwxCrOVXaJAvPfcbmG5cPN5xt4+aIijdyVvJEmodOtFTtuTbMlecg2nM6
ESprUOb0Mr+NV9QGFBIxGSJjQtxSpdWKCMlUxgYJ+JJ5iXo9a7v8wI+eW4kopXyT
Lj0Oz/d5jLj/lo6VR16EdyaBgEfudpmb+ko5BlY6gHcdhEz9eniDXkPas+EUAwEI
Z9uVob0Fdx1E8BA0WCi410ai7H/5RaQ8NU7/X2zf8DXo8sk3OyWPkcHyiIle7wl7
RRmUbF3mVL9wCBjyUHkH5kdZJpvQje4nmPord8KlVbuiOmt4T+TrYGVT9lkCFi/4
qJckkp1UIE5FdpFXY8rKDQTV3Z/TzUk5YdzIwY+2/ojahv61TSi9TXLcBX5ob0OT
NeSU7E2HGRUtbQ/v7s4uuSuJy5YDBjDOaM/2Q4W07qBSDASUEIgMgiM7s6jeuFx3
LKDAyQpNwxxm1TKmN6h8XbMe6h5Z0f5BzgT+vp82LgyMWJwvZmbmpxXcpyxGi5i1
T3V04592PR0jbEQ8jfoTu7qLRl/hM2uAeKcUn/iU1t0EnCfKREuobV4HdbuWEDPK
MngUuo4ihSe96XlMSA9c0ioyggGZp14EueStJm1/qpwm6+iW2Mq5o2j9SxhrnMFq
T4Vqydqva1xMjfLdPWw1LIYDopchxD5k9+E05Ikirh8tW0+nkUgZAcDZGjPkPyBM
dBZs6zrranabt4PSxu9C83xR7kSLfPJPKaBo5aaVEt+VIIxiMem3DrRL6AmMLv2N
sS01+UEd2EF9c3fXxzr0Vz1oWZIN0XkOqv7c+qxWO4tjMhbZgHpcsyyYeBxL5476
SJtx94N/7iDO4pYWSX9wfTfZVlbS57WnGxQk0oEU5uqeWSyD1lZuVvVPOFHju0yS
kO40EIiK8qLWx5l96ATfgWMEqI8MeXPGAfb67LaUKKMGeig1j1Mfh4zxfIhiOtBK
`protect END_PROTECTED
