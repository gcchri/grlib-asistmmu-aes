`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hsJyo6KcQvHLV7+HiWf2YdbANME5n2YLdRAJwBIzwM3TPhAWavvk3hfpxUzZzgUc
iMsW9nuD5nvRuo1KXJUloMykz188pWmpUi7v1VnazFW7+BSMy7tbv92G99VVj5UZ
wk8Gm8pOpWMVSSpN4J/IfQkKwZ5Ye+c5GZoJos3/h/b3+6i3iwrDF5skYZg0FNK4
f3s8NprbemZAw8Ie8QsQfBApe/dg08DaRKWn8HD7Rs7DTzYT03w38IDX9YUSxe2M
c/ajarzK6Tx0MyEDCHTKY3un16e8ZeXgnt6X6V+VZmXkRUBLHdQhdYPdli3UC1uY
zO8I/pyOTpO8tpZuh4v7MQ==
`protect END_PROTECTED
