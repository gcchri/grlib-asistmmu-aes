`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ulFVRMWXhZcnfHAMDC/b4BLtwCFjngKweT8lUcbmwcMJ101sxUEWBslFdES9iUEf
D4MMm1u05X6s5yz2GVm8yMRhuijidI78twN5WqV36X2LLdJfo5+Ew+in/xdDvr9Q
IeWXTczUB6hnRCfc74XhR/sXdWKObMHDnbjV03Urj2BEtPU4D8oKepFGz5K1wQKC
63X9PDgaFtoMsB+4wiIUQQeAesuCxWI7r8m1qFUv/Oevq/cWDH68n6YQg07OE7CS
P9sP2ndOInaP3cUO81otHk+cBnOJWOrHi8uT8ClX5nJhZ28jH/lN7F5z4e85es8m
OE0JLUVWV2hDwgsQdnYH2zE+3AG1fZcoSjXsi2t9QAbLv2LpR3XPoUxCPjSbsriV
fy6dfDsphZRGCi4kMXq1zPQ94e4UcHa9kKSBpaHm6lAM6mFghfJSs8XA84mxYeZ4
+bV8KQYuBKRYEKIuZ9AZd7cN/C9v9suHQ7cmAuUY7k07tI5AnDZuv1FvjuyDOxF8
K1JagQ/TGNN1k9i1tflHM7+fF4pN8FZ/KM+u3jPIzUHCfnTxzMH3zwbGysPJcNRN
pFv9a8PzpNud5PrLP26LqD11Uj3WL23S43OoBGC1Sxhe/yZCRiX3iXt8G9SBSwmY
OmKEBlzNRpKL8U15b09zQZ5+6FATqkPwalrqCQYrVqAwVjoFx0LSFM9/ZvgCQhIn
oC4l2Aiyav5s7vdw956eD4+BrQgS1CEmNjOxyT3hdlcSNv7QM3NRy6RKCMxDRIR2
vjCubc8lV4ga9fv1bJon1XCfkeJpLwvJcKehMjetFu5/m0/quRVKn2fc8ca/2MhM
U7Lis7fGWbDmDLx7q+ECM/caac0OxkIIpFLw1WibnN4UptNmaneF9/ZGut1R5+fJ
6oWivO1GO5fqaRbNGRISOyiHiHwjbHvljtSq65YsGl3gsP4FXeGMMM7zY5Idqp0V
KvQ8Ar9TiGcJ4ugpV3isGrLTxSOdcYX3XVlsIMnfZ7tLkbXwQY2PHpXCdwQZcpM3
M19EdwXkpYl0eAr6wP8sNLYefTbwTWNmi5KJ2fRSdwFmaQCKwCNBdNoQlxHkN4Z7
MZbUJKORj8fkUQJpbHGPxAtfw6NqtQa+pNg3BujQU79hJ+4lpLhGJojBdYJIIqo5
ffcjNHQUSgqL4hDoC1vouMV/DJPSH8FYlSAtPSzVXM8xVlaZ62lZRcyXj2/QZNWY
L2Rao3gaB7Gv1a6sCs7L6JD4hoAH8qByVOohXG71xufEMZc57vTRrOMUUU6khrJ/
kcCVjqm8K8uTwBtCElSEQR9Qm5UPBcrobHdM2pHDwa5QvHb2yDfVKYpKA+6OKOTI
eVBzh3FCGXDSM1XWV4K4iL/gn8j6ivUJfdL46+nr5lwrJUC+MHPPvJowu2jgDDtN
lC46uo20I2RIGvVI4DOo18LNf48JUnzek7ucrqQkABNKTq/4wsojYELHS6wSaehx
AhQc9S4suH1CVR0HjT+Emen3RklrUYooXWHI6El8hMJyXpj7kIipN6LCFsUxn1zV
57AIcnJXUYkw+iFCgrM93Wtg039fAQ9cCVnjMLAFxJUKTYiFuZIfiNB8lmETlZd0
7mk5vk8/kU3NV9Djzcb31QkYbnSUJVpiB9PiPf/JRiD/VqulJh7R/ddwft971Lb3
ocr8JqANuT3yAbXSIrzVvJJPY+mFDscDXwwCUfOoWAHugAyApwWGyNffSep4o/g6
nd8HIBKuu70uqu/jt08aGYYJk6yNq6nw5dEOxUfHOT1TI3sOIuyTjv9u6cw+BdGH
WkbrkQU68WXc9upNEt3l9TVl69OSysgGe+EBK6H1Q2gmjuKbnWdyiX+xoj9EvUKJ
N3DWC5NkqGQC2EJyzvsovuNKc3kwdKBX1CnNyxC5rsAKHXhOav+ciOTWf1BaQVJG
qKkwyM+yXnZR92msfYeOS1HhCubBevq0XilJTN06Bg6Z+kzOET9jO32OjIOgEp+p
TmCFOJttaq/MsjIbD0y9en7+LW4i7w/FpnDUOjSbk0c0Uzb606qDCu8UsF6FNeOR
/XeHmb9NxW55FF7iDSzJMt05MKGZ4FkYCFpYmdqy5vHz6eZEAJAlrwncKNPMLRp5
FnxDLPqL8asjXOyfjTMyRtDVSVkYNIlPCsAddatoydqqNwHQXr2X6ZVm3drAdH5X
ixxaYingEuOC+llb8lUVDWOULes73M/ub5mycyRsYL4aXituxypXvqi+thhIfDb4
5bW+BiXVu3DJbbZRaDOybW0UcLijb9XwIaHZlJp5yCrBusjJxWAUpY78teNd9s+q
yLK56g8TLh73ErhqK3UHJ3h8AqRbj04HrubwcOvghVCLsdmbVhwRQn3HDyItl1/c
80qix7gOhPqaZOeeSETF2SPwSgdjHnFlzi2k+STKMtdJORR+bb3jlnts70LZ09vu
akQ/ReCoFiujvQAWxTWn+Vvok2kzflRZihKOAw/RvtTXz4uY9TBnVhl5IVtIfm4v
yKS3qq90ji9SPDIRlPILwwRoWkFtV3fC2TSPgNy64lbMLsJ+Jl9z+rUx9g5XM7Yd
TSuD/AFLZgl2anZw/leUPDlXd8un3dnm1gOfF8QmUdvGa8C4ud/hxQm50FXG6fXS
e85OfD4ojbjgo44ddDXJrCAbiM1a1sneUm0piZ4YgrQfcxsF4MzYUmNcDvfJb8PI
bXYQN0AOXTaX1+pJFMxqAD1iDDwI/ruC/DfF2BXMjwj6mlSMuIJfEV9vE5YpRbQD
MNArLgoAuZI2QSWO4dAWwUXa8pSWc0lCnJgn3JMNFHLuK9nKko0kOabBlg9hv1LT
Hm0TUogVyuMLivzfFFybEIPhfwO499/xmn/UvK65w8B/49StQExDUwz3F1cjC5lp
wUBX2miwUdT/Gvp9nucBBBfdmyzWVuGU9hT3H6nHlTHQj2qwSTBiTZPgfkWpHlPY
xJzll/GGixWOT+WHjt3wu47z/99oEy4gkW0hnXjoHBB9bLaQbWQwnQxRf+EK2R0Z
Aa1V0Mdm0MbqLhUfGfEK4534PukymSk1rwGcSnWPXwp6O3d+8oJPCSqDmdDxVtfj
ghqFYZZaZ3ybvZ76+qiLYP55xHu/JLFXo6oVrCQHBB5hlBoBGV3+yiy1rToPHaZy
X2PPHEjP+0mW7/xEP5sgckGuO+jpPDt/7pgG+EWsN9x/unz2ur2cGo3Pe5GpC7RL
UOzB+iwa99QgNZ0ZJMsA6dFe+cjEwP+jEzYdfQLd4oItxSxEis+lzUgZyz23ar9S
Qrk0fXKk8Bbe+dxaJUMTlzAXJJcVkMi6jAKs8aD/PzR8e/wugskQkCAxiu6xTwa0
NuKtxP3u/jrmnJy/mz0zx0fsDkIlhzr+9GUF0lLe41kdnkFSGLVmWbrcYuSrANdV
ozwms8UPPCtg0IMNe0mv+57L8vgPaAmXenN4fnRuy2Ch/LoSP9uda2Njr9dnjRqz
nOeCzklorGu6b87yfd3/T/Yaga/II0exoZPaV7Awq6gCTjJeuZUgFuJP/7m/x7Be
hjkK5E2TJAhXnhG/RpNEenw4dnpUS8n5rMB8ZYPqKowXMikkOCK7Pp4tkRIW05l0
rfZDVGzMO18MSEIwoptRe5Vb/ynqgVUYLqqJKF+L5A7JKJwLyzm8AMv0FTGBdXi0
Z6jWcWy44+YFLggIRO78lQ==
`protect END_PROTECTED
