`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ErYcvI0mXoqTw0ZEJhGreVL7IojD7MIxSHQKrfvusJZPpC9d/1ddiYRlLnQ1GAHy
AMhR9yOyQ+kCSb59DeaaquIUJ0tilVDOME7zZnDVBD/PKr8UgVBOCB0NO5gNOG8k
b9TEzY+EimEglMF0LbolIqjs2dXWfdWAf8Xr9PJmhz/5aIeJ/L1M/Gl9PPOffyZB
Kd1ol7xkJyVp3TF/LMCcVEc+13sHSbxpGfTDgTaSkAYuQV9OngAynsWBkLl33pKU
NIktp3ipliecqIhEcmQXy5WqqePDox9jyjBMW7XY4FgfiyUbLgZDm/LYyZTGBmeD
`protect END_PROTECTED
