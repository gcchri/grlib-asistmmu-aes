`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FDx35QYppVLKtBzSQjHTNnPgtPzGEMdZuvDYMu980GikzJbNPMKjGeuq/5zC9B17
fs0IfLgQ0/fezM765bKF0ULZojEdtXwlZ+ZAXqhsgMt2cDqzCsS2PgMngpFUt17v
75hRtPcy/Khr/X62YVgdD3omtPT7c8DJ0wdLyiqB6/KRKdXprEGk4A2mKu6I2ssK
+fb3snXJ+RhEd1v4+wh4vSdkVwl1TNdT92DUPfztGpiPPDxKY3HIP7vYrWw69dAT
yPbTvYIjnXeNAFu6b5D3iCQ2kKzunBapON9KW2IJnC/TiGf03llK0TH2rcpU2Yit
AoDGR9uPeL1bTJtLHkHMXeqAr0gGRSd3XkNTByddeAuVcv3RYP/P4IZyYTj812ed
e+IGGg/TEJJ4mxUHpP/vQw==
`protect END_PROTECTED
