`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M7fwr7i820Z0O4C6cYFHFeIgIWVrJiMXjRDcBBskK/KTg1pRd0RMtWid1y44VKdD
cncZirTar895IY+GNXdN6o1WMhtrv+SWv+xxGDLju7NT/o5wsDEPXrTp4JOSoATM
Hc3cLqGaVjLFdW+giiY8qnaXTFoCTR6gXohtb/tx1dMLz1ahziE9lQOpwtFlR9ap
Hxec5PIHvhRpuErP/Yt8Gc3y+FrJR/Xs4YE088eRvLPExX9NAiJG9ckzQOn1rNPj
dS/H6K2hCxaooELNz3i7IcZGrzcyrNfMwAkcMK798CmTnGunLRkns3T5q6WTzV98
/rMYPgAgRxHdyGkfllafQSAVmIcGcDR159RWTa8QK/bBB6zCopKPSbdQlLpjcz1s
y9060KaTPPQ0ipiuuqwoEd+svcF4Ys7ANIp/XwefFDzMkRcQEFb8LY+zoSBK8SxT
QiO2lifR/RXYYOMV7bY9neJm3o08815ZviDQJeh0oBhxGHKuik53/RhzKhirAI5L
TK/3psN9I9Qr4QSQx0u8IA==
`protect END_PROTECTED
