`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
38/IePC6yEFeJPREAg6TNwdtjioiMZ70POm19SQ8RGO8eDNgmJEeG+UrsEotQVlu
FK/6cCr8ttoXacAfWtu7Hv4CAbbLY3/XR4cqqSChpniqNIUloyQ0M6gworfQJcPc
HigPQc8fZMcM6lFXIr4EId9M54N0gLKMzxOgESeHJOms468FEO6hk9WG+YWhifF3
DxLfkfHrR7pvHD3Ih97qEBnwFgNh1ZVXwf0pgmpE5HBzzcuNw7NUGReFPcMvFU98
0PbaLD6bBYCpb52sNSitE+ZCsjfUl9zo2HAQi15lr7umGvF8bC6EZQs69DIMnEPc
3hjAVv7Kgu+t7WSJnHXNiAT7JTsPhDBXZfnvBPtGU8T5xzwaFDX8Rka4+Jhm2obV
wzyMcSv9Yq3EFaxGO64DNPyRsLjLTTildYbvs45W4xFG6hK0G3Nz+I1DTo4QXxmr
`protect END_PROTECTED
