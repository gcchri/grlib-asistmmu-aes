`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EgXeas1zHhiM7rivR46fUUd2Lp9hS2KBE05f7vi0gdm1fb+HXi2BG0Imz4wNu65o
EnFyZkARTXnQYcNQVW8PD7+ObN0NjbLhMBaobtO/82Fn/YAQTk+N5AHcLwb3xaKV
jfFhzAEbWjBlXYtMEp2mO8ZJnNcrBpHj0uK/mT0PA/agBu1HrjuBXMjYKQ6/ybKA
Tj9cM97pjwQBeEswnOQ0Fvi9xu1gkLGD7afstBcy954Kv+M62GUws/1wgRL8EJ+B
oqGQdS9WCXLrcGKsP6iPAZOw1gsmw/hu0ApokwrzN5f6RGX/Rf0xnz5Sd3ZHEYAz
lFyW6uDCw2czC2H+CtdRb8/BtZzYozx5+LRNti9yjTMuqbcp6+2XU7nUYMfRRVoM
ACjPBEeNRCkoplMSbrUQuNWMpXEUwifIy1+cMbfQaVKBWO9eG8W5LcKjdEHaZlun
/rZ/fNbEvg8eRspU/6FY0MDicNp5tGy9HX4LSWAWIo4CqbZ1sTRLa37go+JGFkYR
Y+sjmdh3rVDKhiyNOyUqNrYRQZ8UT88d0fwmIx7CYPrwIMjfpUIZAI4XYiumOPEZ
38rG83do1jcPA8GCDSUjJbW7yL5TedJjE9NhylGO6yDs8DN4i1GHmaXM1hvbbuHv
SQ9HlI6ZPfuY3ahKZD1WgiSjrEVzqgtBJIiA8BXO9BBivbu5tZY/8viGTUif8Tar
pURAVkzOYobx7qCu2ND0U51NYrMMYBXmkcnarO8gIRYjnIBjf2jFI+1iIYiDSXhR
ymUGB/ljJZsGGbx2Zpsbezt+6aHBENtZicksb/yD1G1zUffA2jfkL0NHeQZHCmpo
OwkV+BsCDF2SR1xznKTZ5Fa7BsGpm0GDzEIdGCfa+tFBCR9xlINu4qhq+7if7rUz
Pruml21Bt5pD697hF5eQFcur/kZyhu5uXQCxgWkQ+b2CeaeNZTk/6wr67++vV98S
i6GJ9m3ySoXpQS5nQaa0QpzBbvuY4wM1Yrtp8d4pXtTHBic4AUnRCB/FxFqUOwDO
Nw/tRaNuEYB16zEVNCAsSgjro4sfBiSQInEN/sWsnS3Mei36Adf/OKP/4qnNmqYC
aZBy2LLGCGVm9DCpPIiADaHwTPgTeJqqzIiUk4Avl+L+Web3QoQZKnWWexBY8fV4
WoOBBWdAi5V2G5ZagZhiGYP5Z6w8iajYGqJN8VdUdjJF1gFkoOKHSBpQHF4nD2MF
dt1fERkWB7fOFc66GUBp2MKSxrzbYTf0GjOK7Usf2VNg4ZoqXPqHLa7N9F7AUBao
/gp8uqZ6imxbnX5HwYhP/eQAcWDkbVxTDSLNsePQizPBDQcconQJCmXrD02D2BLa
SiY/j3w48IYbG2GK1EwrOIocJAZYheO2s/QSpnt5sQS+4lK1CVYv5u75VTWFvNjI
JsQbiqKlACzVJ9xuqEkHhW3g54Qse5cn5Sz2mUonstIPfuSkhMs2d/hwRq6Hl3EU
eqixrQTFTnJff2vlEAuXRionTA/etrs+5FKEO2Xue1oAwZ9NBjKxOMhmchvulpJa
qxe3tqckRvt1C3vmy5gHfng7rJlw8DgPNwvLZ6qsZK92Bi+rr3FMl7dNOoMjsd2a
O+NqZaeWgEhVgkHDCPNeqfau+omUB60osEZfap5SRdIvceuT33940FR0HIXvh1py
CpCYAGsxOCJ2nMVc1QdoUhkx49C7f85YcABsn6+9SCBKx/sqfMtmTiHQT1/onGh3
i/i1lZMipjPhEjc30QoWIP5HET4qZGAH0SLdpN3E4uN44mslUEeq4D6MkT068Clo
2I8AqgC7gYokIDV0EZ0lF1r7Q37aTd51hCVSfkhAx1NcFLgkGiIJh+qln/p/uMU5
pLEypME1l2R6N29rYIyDXHInbcM36n+D3JW+M9xAowqkymyRCMIPt7fWeKgiq/P6
zSWgtiOq/nLES7j6PMyKyOFHmcmttSYlOAfmf1G5Sc7PaMTzwN7ErAK8wUz5lT9Q
bbsMoKZanPp2NNPCVgEIjVjyqCsNQxb6fsNLMsd/QFRfVF1eD13l7zfgRjfc/Qvx
pXvPSGZNKj+poBwDbnyKGpRgwQIoVy0E/FnR8+0/Fqm3n2lkaEXo00SDw4GWjmar
zkKsEsDjbLq2pldNr+Vq7Bnk8HQCFLEPu1ZKnTir6eAP2VDPOYiA9PWNPjYH0fNG
8JsyWtW76eYxVK8Lesh6eLC2Ynsn1JWRgHZJVmVlwXTmHu8VwPuEUAbMaZH9Od6D
GyLT80zJeRBVm2urPmLFL+6xGotSCSqvzw+2d87zCAe9CST9xN89FVajlPgcICtq
8aeZc8rGArXfb0Lzxq0VdPLKJxmHsAJ3lmmVztfxQcEzEHWRhM5t0kpG5jUsmzhF
aVQoHvsTfYFQ/JBgcCM4orlb4og05wfk9v27jIioNl8FYSJ5t0R0q0KbwNfbnPJb
sx4Ec/+OpgPoEHb0C5auOCSg8KsCzOLFwg19a3IVQW30whw/Phffa3BfhaU1tnpO
xFylS1BU3j2nOrIW1rIwnNSb0z6znixu2RtQojcC3yz7UUNIdg5jacEV+3gb02QM
ZBLhrFkS2fJfW8s47BtsmL8qkwhrzY9QTQbxeIo0CVlaG5n+tulWG5vfpRpZbA4V
XbG/wd9Ej3Xzhvvwfnr/MzeVDAy1hSVE1n0X3sNFG1Ak2SpZ+7nwqFt1noR4cfya
IiQOFCDvS1zgdpEb3vncGeLTYpLeYwoxAU9YiaAXSmKautWdcY/JwZSDPHyyQ/fO
qhgxpTciBmNrrIXqThMzIJLPQSXQERhnNzDoQ+Mo9i3QzqtuDzRY6Y3bXnw489rm
EJOAmzOOYNRS5IiprK88AmqpKCOQefCtItsPGyywzC3X6oXR+J+7SRnmLfrD/Bvh
eGArKHapKhEq7H914rYxgYt096+lUg2/2OEfzD/U2BP3LsE2PFeauEhR71asdU25
QMaVUsE8afkjhoBMq03XuJK1+0wEhdrQb369esdndPyVpM5HUzsIyNGpiN3kF20Q
9jSWtC86jxe2u2EzYQOKKQaLpHQIq4EG5wwwvLbKQwsJ0IL2kud2t0IMIIxY3rkC
qYT8ko1JL/YZivsbgBsawD1zxteUKeSuuccc5mqBYVSO+aMQmPUGOPHJ8LdBr72z
N/RAmmdckD5NaGyNtI3YsFPHxNpJCvTqb4RRBp7n+2yyyIjZEYGiwUP2vqw9cPf7
oq2201CwwwF7QSOAEeydFq3T0QpZOQfL4hxmGStatxkx2eKwRnEdZ8euDC/2JMHs
+zq8AzFEFutBYA6+lj9zZmcyDlXaNzKxQue1irRkA7oX6lbNQBP1IMnQD+G247NJ
qrwLHXfh0fOqjF7HENeHGctwMwpGSfOs6fkQ9j2AT1W07UKPO7l9V3IvdkuQL3+3
ucK62y9o00ZVfskP4uTIBKcU5FJGAITRASYIqCMShbnMZaV5DCVuOsq/xDhQn1lz
m5Os99lIWSjJ90/Rbvmz64EGE7DSytSCrTm9P/SNt//sYotX3THO3KjPyArpl/C8
QO4JwBW6NNrJILCr1CUAUwMvcU2g6mYYYQXJW3o6GWTARSjJLJm/jCvItoSJq91c
adZJretZ5gj6Obrot2yhenmjAOcZ37+gQHiHdd9bzJU7alc1fWGftgzdoMmJHCkG
21ZOO9+jnxFGGx0WfmOawEQKHdAwjBlkSDSKX97pw+A0dLfoganixDeBPVUquLj/
IKhBNVJ2DtmNBjl63+W2LLKPsAPQBP7l7EQLf1cVC/qkywDcmAtm/Be9U/xyTxv0
4RO0e0qJcB5q0Pv063cN5hnO9E5YJ1lx7bhTpR3nCIiSuLUDH4Ig8LSeziGgHyql
pBhmULmGEWX75f56H8w3Re1XHP2GAx8uXS5C5IL2oEqkG7uxmtgXQb5PPq2Puk7h
jbrlk8mjvw0qJMu4GkoqIq8+uFeJeZfv529sWxFFJvhPZtprsIf9FsRa2jebdqEu
xt7SEdSBJRxWPS93OXfEsUm0d57OIrVO/iJyZRpDQTHsX1uEcuCl3v1qEd1DoA87
Hbfl2HP31k2GviNfH3wX1FWXC2MnWNWzbSKKFZL+SpVcb6XpvBzSfKY5tsO2sSv3
F7adgHlyvaPre8Dsld0I/TnbZmh0KUwpXFvOcE9EjlH8voNaZaReadyIvWncrwsH
6muVaZWU06b3nr4eKGm0YocRA9iDGWR6CWQz/RSI8OK4FtUwcsIIS1Up+Wk2sXIa
bwgCuBpU8g1IQUWCjkySvKWLIOz4eUOOr2E8Z0Z3joQpRDIQFB/TAf6BI82dUeEh
Jd8Dpat8cXklcm/uEFpKLpTvyasjaSf4QYT+26K8Nzzw5LWBrbJwsTQAiOiEMux/
gSyb/H/Q/PXUbhas3JvIbRaUilvnWK3++vSXBhWxs1JRSGLMOMS+BkvMVvtGFSnc
+mN4kjr+d3F++T8OTIgwKwFc30LyjGLLEznyk1NruW417BMMCJUPlwuB+8uDk0FP
U5N2ajCzINCbfbgJrt9Wu0MCvmjC0vNWLuNmarQvT0No1IMx06wdut6W66+vH8jk
wMYPgDlSi7TmhtBNq9Yr/bsibTA1LcbFCG7d6csqzQ7OhTr9CbXD5tvh5Cv+YKvI
qXgA0PkoTGRekhyEbr9h9Evl9FxXjtY+XLHD+bNlF19OQrl3kqIHUUB4DTyPF9yj
TaTn4CP7T01/hWMkxSSwEAOML3G1/Xl8/DsBB1sAHf5TGFM0bWX3lhbDmEz+qIfS
b2JG1eAzFYZuzfM/clzMp0wsdu8Ffia0ZwKYiweRxNbp3CN2yNl47aJcWIRGrTxp
LbzNGZMoV2d/fj2nOSeISeohpGbCgOAfdZ6sgrCkC2RdK8JHi9AlxvTBNO4empC7
gNymPiY8ZxqHuvGriZp3skmE6i97Alt57ObXyOQkypHivfkjyxB0BjZGFWym2GkN
QRUyqf8iSps7D1GxPzPOG/OoyEnCF3EVonqXdaWXDPaxzJUozX0O2eUB0GiO8TQh
YLFVOW6KbKgppXIoIQR+csMpHu5Q7FriWTal1aJcQkyUXWHDHNKL2iyzehAG5LOT
IxLrPGZVpEVgDNRBk09uHsaaUH26/kIRgPPK5FkB2w9jHyv8u+6nZGtCJCVyNeXA
mF46T/xclS1sMY0k5+JfyrbvXdWLsTORO5jsPQ/9rl/uHjoOBoUG29UNj1qvJw5z
/xdhAZZ+bBMXCBoaez48fjKmeea8hQoOPlocfVDBgZ/of5TT7AWpWTQTYA85J7YN
m+E7PPJD6hNvHudqwp2MfeWNpMav13sNVOzUDAyvlCVRcBf5VkVJwF2K6L+KJeGw
QQYoyyTmZHX2fIGDao47xDj0zAkScFG64PU0nW9wG3Kz5p28lG2Iw1kCssCzv4yo
pEbX1oVwNcTUlEXsATCSM+QsiWR7RyJdmK5wTdDZY4L19PCY8d3bb9wZ+8VGUX5G
DT7/wH9u/va3LbcRzBPaLAUwZK2BVfKi4BkP/Mn2HqxTAmcubQvKmgHsnt3Pi3C1
e6reXFCIO5X0LkhhLeo4rlsQWdquxApY9aR5wdwC+K3fBBWRf66i+j54YI/C89X/
ouk1KCwmfMBG2rMh+HrL4k6I0y8OTeQfqIBT7sCr1r2BajBLoCuGRI13vTRqPGRX
rEHm0IDtOanyIexzh72LRz5M96qjHR5V/WMZgmEuyEaKWlpU4eNGze8flAqZSu35
pnIUySi3JaI/QU7/uX8QM08I1ShbwU5TnJ66gDEXPAF5ePqVBEvXJ/J8eTRtYsNE
KGuUG/H3zLr9autIPQt8uTdCHMRwlS2IneKdI2OTFdSMG00AaRH0iYy9BMJSMq8u
j9Uik/dlbb1JFJkClK2SuM7wJP6WVE4qgNkybVI+vQhfl4OHItyOsKmt4zzjCaKp
lm62d9u64x3Ua5/nMkMJM9R733h+7EP1lv+uf8GG+SNnC59Ar6YsN3UMLBkGbb0Y
c5dTCu2yVxnzihuXUP69eGLkVHdtEkBas9tevemLLNr9q22+BO3PybURmK7BMf5X
XCjerKAumLOcqS7jsUYG1IWtw5zmys8UbZjpp4Umu0DLvSp8URjbWRoZUQrDk7Rp
QhneCPkV3c08qiOK1tCtjFxiUVY/s/bQ0492sfuOvqovg2co/7whCyyUgVskbAaV
/jnkQpRyQgJRmefx04H4xtVxYI8H2QJ6zj6NL4rdHOot966nveYfcTc+qDaVip7V
WMmpkS5gEoz0iA6YzVpOEpWGaxOGMzGwcKEFvwRzoG56VoOz229sxn0pH/uFV6o2
DAZJQ7SgouxSARdRk2vuUgK6Hza7Wa7F771fGesPaQmDPzxuclrmo5ine4E7SEjq
dri0P+26/eQ3jy++TbNKyskmET37KaYaFJf2T1PLBrSXcv6FAPzY4rCL7QnKpNks
i59EH9ngxeSNhAw0fvMkn1h67DMvQXaiUHooR1680WWSwgxhe0DZdZaJLNckiPLf
FT+iOUC1UzmfI8vGzzfLhLASH7qW/hD0nfu7MrO3G2hJc21SgWNZodLzbgkUR1td
N2m9N81acxfpmsYdLKS0PhcSB9HzRZtAEm3NYMhplOWnuSq4lay2XP9X2n9fXoFI
YwAPDpDSjac1VBAD5AfU0ATqcUiDR4SiBtVaVgVF2dZrbEY71Kdi2sx9KW+jv5g5
zlUJGxZ64LgPGjuOZTX1Yp2aB/bq4aWFqkxLD12l02OvuHgwRLu3l+njoK5VROL2
aMC0em51PK5TK9eZ32qzpMVEOE5c4v+gBthF9V2+U+d3dk/RSXGqKyxyC5GXNjYY
+bBXSqxZuJvMGrjtW41ErR+rt1i4adUAr5QA5Asbiiz4C7RS96SdU8hp8a8TAcJq
M99Irs6t5/kOYOCT7XVQ49sn1Oy4vKK0zCQJiM7l5jHB7ViLB/Vq+3UQ4QBI5Dsw
qdpmjWIXaw59ZEfFRsjktwf2GRi4I6yBdie6tihN2a4MneuwncvwsHSx68QxQ39I
2RjrngpSXrI3bFEJilcUXzQ96y/kRYKprFjWdA7/dAPUq2PWBVgubi+Cn2q5L+GJ
2DdeTSYC+QOtb5iVqePPAoK/jm86BL32Mrt1+UDYJYgIi2o46Z1CpX9PrQh+TG4H
o4xZYj2gFYTW11Ej85q4hqmScgjBh7eHdhc3Dr2DmEKRbnEZd3v0U7y2wwKY+Qib
JnEkfzfFEwPTtIH3fvpdxQ55QEhCfE8w5IdJqYZrjOSonIIvEG/c4yu8b45NARNk
cRL1saBImpQ+eR1df7WTt3lMKV41UuggtvntROsWoZnE48UyONBaKXHLGDbYMBDF
pIr23PIRLea+Lmzd+Q4XZkY7a4uj0cbEdFjz8saJmkKL2xq+LJiDACLo/jJtwr6b
ooV/7RdMRqRe0KtWZpZNrd6rBcsU7aT4peZhpAWrZlBqNWXd88X0F7SzlFGyY61K
WtiWqIiwtVEh8XFuscTXyADU5O/jFdsXI2x9d/ETJhPfgoMWUPKCDgG15IqM1GES
IFnQKP/FtsJKGloVa8qosuIkbJ4ZVRdzhMZLkUNQXe1bSEfJ7mvaxgf2cCg96QTF
8oFqKLZQRz1c3Qp44pKX0L2JtBgqHRqICbwCwO6rSuKHGzNiSck/IDbWtHlWEZ3H
AH4XO1rhgY90+BjcQt2eugnY6J9RcTVRiCG8XzCGjRVaddCPw+RYXJLCgIfarArY
V06Is9FrJQtKF8lk00KeKXgtftO/P5mrXtR4d0Xyj9EglMCuL13dm0aTRpmvvXIL
NKqVqTUZPRsP9Tc5RdaBeG22qPQ7kTMbNzUUeD2qtWBxjSfH6oEAahuz0YpyTili
jiJxYkAId4QlN2Jtp1YPcxva131oPAolOKn9oLRo2pwDNii0uEqHh5jk4xSigzsw
6aWgXrnCKTcrG7DeW+PhhVXW7u4nLZNADkE+OCGei5omI5fWt2lCBqE6zCZvsvhV
FcqDLehhjnzp6H+7nNVC7EhX8GofraM5RMnl6G4stTsKWYbtITgvs9hyklq6DTuf
25b4x4GBs4R3sb7DKk2p8O3zSWYv4bsoarWNzv/wpo92WqTqqVNyT3FCVNixljGH
E9tp/4fegBbCMJUYglQkdrVHA74pEqMaxMm0z69ponmKIrx6zV11XcLVrS1jm1sr
tELKd2eujtqFAwU5kXOujM6zJ9jfcBLnq1muMPKCopENsf05FDB0dExaDDscPTvo
UAJ1yzM+kxZlRa2V0drh5FZ3N485DnbyBMZxIGp0MTqtGSOjrWLd2fB57B8pr475
IcLCgNn4Xidn1bXdjO0OjxgqweYRcQ+9Uk7Uc76ljPEuOW8Bw2WUylcI2hD5fC3v
xwI5yLVX1YrgjRLotL7A/yA0Z4EhKswRx1dlBg3PJBssXHN1QoXmeNQgwBB+WcrT
bWoZcZRIp5PpXh+6h1fje5Xs2RNqUBs7KJ6UKug0mYE2QXgwbfVrZmyyO3gvqhN7
EuZecMPr3Fi63rqHBddvpl68dc3hWMh1lpeVvoZuNaa+Hcyz8WG+TixRiaF6eXDT
6UIu6O/8Gh3duCuwFo4XQQHW5GcJZ+kDtPxcAuDdGqAvApDAqRA23tC8GkHtOflD
Ndb2PA5UxgykepxGU61jeAnhlsrIb6bHy924aAnxL8+hLMhuu010xEIUwx9MGC0K
fyiqNibZ9ZCYI9q3L15oIvI7X92lWIth29pwOVzYhA+m/JRVrN7TVF4QFn9mYpv5
c51WmeGjEFKMtddyWmU2Kb2bE0trY/35ctDpYw3hJYUNiMmtIZIyYCaX/8UXoOa8
WA5HCeFLb+PuxNblnuE6Ia9W4akRE9ZuWqh8xNclKpwLOULWUersI5D6i/0mbCRR
d7nt29Z4+x5D2ZkRY33okdqSQm5N8iYv/tQFGZUvJGJDT2EqIxNy8tKRNYzPUzoO
NCgOm/4ceLf5+WoxUhfREFpQOYHnFKoykGLFK9Nx02KJUMEG+enOKHyJsNKjHKZF
znSB3jT+G2oyBrfPFGGsJhKXXEUHXszpedqbOVAz2A65PTu1djNTmiwWuwLn/S7P
Bjekvw569TQEIC4EOC63UV/tkjWX7T12y0qA5DYbU+wku6lexMyw5Kl+aOYh/INU
LswTNy+AVvkm4A7XyR4vULWE+ObErwmdd26j5/9+KFVcBl/LbAt8RK4r3SP3Usr5
0vIt4jIuupChJeMYmlJzPQ==
`protect END_PROTECTED
