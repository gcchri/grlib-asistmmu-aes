`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vD75rj3UY6w59ZpOl+4dP2+YS1iYVWAntjL/mnPLD+7yt2QHqMbZsSwrPIVoSC/Q
0sGvaIm8kM/Lb9TJDbHWqUol0gZ8u5kgY7XVOOFhm2+zcJy0F920PUebKID60LUR
SShCXkWdBvUufxaxBD4QF/CT3nA6Gnxj7CEuC3kPi/eICZ3SrHDDp+l8urgjB6pO
trIqgcgKY6uZyqca65fOrOMf9I8X+H9mdwozFiCNTRwRqNUtYvIvyVZ560slSGIB
r7o8YlKhUfSNeSLEFXtohVUE/hTxl+BiSDCp6chIbFu1RwvX3Ryk9x/NTWKQMngl
NTD4erbxelUqQEhjWAMOZl/bRlUhf5Ncs2gYnbVijxfhao2M1+gjjf65/3SVs1m/
WGt4JZlisjcpOrM4p27gcdxrVvLhGNI3uCIQV64NJkEaI375BM3Es97K7NiWxU1k
Bot4+tRxuOMUc6eg/GvRYDYPhoYYIk+BcHfE4D2MaA0oFg1TDHoiOz6HzUbEp5rJ
DNTgUqcC2TbAgjhEoVj6Ptwibure21Cf3NosjzcA6Ly0bO2gLvT3wwWgoKYgFLhw
j3UDBlnsLjlrYlgEkRfkm+WQa/8rRUUtCUwnr0jlJontGPAmE8aqncI6TL+gYKQV
07bQh+5551poMnyTWsDxgAsRH3mkSzjsD1Ijkg193SsfUK8SNRC10oc4nFYQGR2U
lWm5PsDaW26Jx/E3XXLRmfA7WQyc5Ut00t0TLg9eI+Ic6bpkr1jjJCq74wirNQeA
2RQxZDGMKQz8JLuy7zBXHcBb4kzwaGymqntCTRWwm+RuKoi7ZTZbcl9rmuFl5zBu
5AM0NESHJ+zPug8pxi1p+g3R3UcPE7QLbUzNLTMeObHpEnildLKYNYtldqEabf96
6cnhDlrHj2eTnut07LrIJGB9RygSuuIayKPugT0z95IkDDqeQiJvfscp2qhwABIq
XpqGwCWdTMVxw2RRRxeTEq5exAfcyUnZSnxZhGAA60TfKq75gIqREqziNNK9bmdC
dVrDD9cwLnpBfoX0qdqvs9fEUYhxHznJ54iVgHA/xskwKcUPiItOevUVi8Fwmkc+
ZmeBKmF6a6m+rJrHVzXuXbakQgxtH5U7ybOlM2MhtM+ewSXdRrifx+YBzXck2Kpc
YPoCDOLiIqDv1s257c3Q+pILyHbepWybrtvcboTmthaovHgBB7qY+UD/1N5JYuAe
lETYf16yc6yHMjScHfUhDYAUyictZOKZmrYia5Uk62cRKLfXB4qP3ZhbowUIXKsB
nlfjepyZwnP8nY91ruN+lX+L29desMQW8puNkTTBZoOUxk3KMlMbyOSNKm/sdScx
IBdtEWCCLiE36mCAdUAr1aDX+qh2AC9pJ80h36kuauSg5rl9nxD0JxaRUX9wq5SC
jfggEWSuWEVlVnsge96MDwQnazehf6bSBO2Z9KfCCiIAw+D+HojOVxoO8aJLmdvD
3ZuztJaW9G4WLERPxXSAze1+x77JXFXKJzFt52EHBxlZKhy1JxVUqIfQxajX9c+s
9C+Pgld+7k/HAgHP9kgWuJj9Pj3+tTkc5uwFjUuZ6qhX/ERX7kviQZSB4dCq6D6e
vMiFtzk0Qs4oeFq+JHj2I5hdvEQgw5MOATelFfjZsZ4T6nz0QysLsn/D2oTB7Ow+
M9OB/p4RQMP2IuRy4IBGFV/LknorOhMcg0pjWv0hH/s36R9AeRMJfkT+znocKygH
QRNj9qoumIkn+3vl9sKuEaRbIe4phEOkSr1wgGA59t1X00lTeHhiO8UhwDvM1EYb
fYHIia3YFztfrHV+mYYCdHlVRfkeJUpfGS53oOsv6BB6x5ZXkCrfuy3pJLzHuaHP
ifccNDeza/mmZg0sg49J+dyFPKhSFhiqd+1rkyliQ6xzsNLcG+BGga0ERHVZAXbB
l3dtyrQsUGPCzsQeOzxivCFRXPUYm5CLGNDWKt+g9Q20p2NpO2UCjQbi86VwdY4S
eqMo5ZVpuJ33/c5HBY7Vx+JJeC8TQHSGYTaK24CQjuDKHE7xeVBPN3FyNEIuLbev
9u9+vHMpojaqrpPCuN+VJms3ih8JEcigIViWIByGevSxrobNIPiWWaUKN29wzFUM
VRjxBdF1ndlkQX8m9NQqpLL/lLTknMbklZwUNGXUTVNM7by/lK7rPCwZwaOk8Jcb
CEcWIUiwJyvkZadcXKOvafctbTgbxRXQCBhFYZAnL778irxA3qH1eMdr+9wQj+CE
YqmAXpp8Upvpc71oywFEl21mpW/ywMZm8a6aS1JTbJ5piwDwbFe3s8IMvHUcDGLM
Xt0acA8POYKFOYZchv+DnirEr3V3dJ+ymt+XVFncIhC29tCxJ7tkKr8E35H9cfRf
mqCPWY9lD3BKMWBv7nwfBmm73wnVFLG8R6eDxzunN6L5uBYGPrU4yLCww579YmtJ
OxImvN8koXJ09LtLY68E+CYcsKcoisnB1Y4oSwie0IQANmim1hJMLbaJuGgszP8m
c6yxoXJFbP6NA+DU6KMO2j/mtERYF6JzO+PYvNzOeKz8FnOB20b0Ng7svIVAcDld
abpFI89k7q2qLMerzRo8YuaGmFBKK+uXFnrcqAA9fvODSlzsDTRS+40wAjk5PeKc
Jk2J+RIz9xfISpVIe2Vg4W+h8+l3yNJTE9N386Ja71H9pu7xY9YbnQa+BqTFiYXd
2KLuMzIVQ+c3LWJT3uMXbHgnVxFlYFxtm2uGHnLMdu1jZVrAL3EZCi+a0zgp/0C0
FmK+GKmU7ZHVpmAddKMHluXUGw7xn+ifwxGOXOWP7haEWojt33UXsoKpqmLuZng3
TERLlqbFg0WwWlGxFdqOQOfmitZuolzPxLj8ZR0BlS1gPSbkXEttIDFvy3YlqpVY
+uZbb3ainekxRw3di1GPPMs4sggerKq96gIXD4vKvC5iM3A0h//NfzR6TPx72b63
OrnnVNELw7jDUpAHLpakHLFVyvjZzOW8+jQ7w1uphRCFosABx2cT2CRF7zKBwyzv
B2nti2bpIwGdLg+J2iHZQAbZAc9r23J+T+ny8w4fXu8=
`protect END_PROTECTED
