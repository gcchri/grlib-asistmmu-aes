`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XiL+A8+8Y/1rAjP2HWJwyd2vgc/YrN1swUtrcrA15uhwzYUsCdBFYK+xvG+wJz/Q
QZdzdDpdRrhegaLqvNgW4w7EkYvqjCuJSQsXHMVP6qTpFQMavilw3rl20bcWLpUK
Alh0htJLp8YpyAM6qBneTvRNlVgWOAp3mVUm8U7vJMVxSGENz/Fym/7UWJGO9lKx
yc9Boc6WPVL73RDSYabIg7rQobQr1GfmYPC6uzbjojx2m+jhFj98BAyVjjLxsIK+
C3DaGdeY5h8j/u7XejLvsXvt48D9VQcqCq/QhN1YW0zhxBPz4znB6m+0g32RQwHH
xPEUldOUWvBysNw60ozhfCKMvNegK5wyTDsh0F3Sf4mK4o1PlCJgEPyGf4pky8ta
SJy3GnpEVmLao3XFhvXIdArD8HUSw2lfRV/Do6TO+Nb39rtSUtGHOw5Tezc754sQ
`protect END_PROTECTED
