`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s4JTarxT+oHp4OVzc7amOlTKRRFxBa0lwvQeFW+zcfzwtXdYbBZRIWKcBWCucSFH
BIF1LI2prYP5hQuhOnFr1assup52Y5//zbqSzI1XpXpKLLMwDcjDFuXZiBLPQySp
uMgY4MEf6zJ3I7VZyfDhwvJszzprG8TL/Y2D+pmbIiyBCu1UaDbm2ttS/z1BocwG
HhsMRItjQOcWv9VR2vj6dXhXe51wE6qPR/hlMB6gdDZVP3ZYrK/0EQ/Vx1v4K0yB
Q+VM7t0IsJjfxSiu83vqAQ==
`protect END_PROTECTED
