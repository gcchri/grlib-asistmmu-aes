`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
swlxZ6t0eLZzUgI0wFws1h9JX/X6NeGL0IsOQXE0mYOY1d4wjAo6cD8iEWneGe56
GbKD4V/OFomonQbyNvBxo+YJKB16z1qW2cKcS79Q33tBi90y+R0HzBUi+O+q49Xh
aj6MtskqlmCEvYTpzkk6zbePXLn3Mye9VrYMG/gg6hCwvvmRFiIANAlV3rmj3NBB
XDdxRvIiD/ZS77YzncPxC/nElsaO261GeLzpbP9R6PwkSOYuRb6JZuKlvaAH/1UN
OXYLT1AHvSobvyv8nf5Shp8L2SdoTTQuUVIChBRUxjv4eWdFkBabZqNZXMOKxynI
4rY2Hp8uQVCh7rJPzEf97x7Wdxmj3t4lje4JjDU6ujSSqZJMoAT+ulS5UB0aztRC
Jhlh53AGkQMotWENMAc4KAOyCJnBLLgUlsJrgJmVzso8GGPFt+2LMbVIiWfYZR92
Ya3QVdVpbcjQ1ewwIubXk9H6aH0o6MMirfqyi0LTNUKB9Lv8IAQYLy99hVCPp5Bz
7+BswhTNfvzeMhqrDBudAA+o7vBeLeypu282d3oCnWLWjXh7ExHAdd9kOub3Fr1A
fCUKCUnrgwivAdIals5BV92FkmRPqRlDH/9xoZ/TIT1u1ErLk2EMQ1bcSK6RhyFD
rNe7DlsXEUWiabqPK4enTbWuw7ooa0T2EoTuEKQtJfjJuu+g2r+HFDR3rw7zuYK0
O1syTrQuRYcg1aIXX45CEUVHU2/ubdNkxbD/5qpjBJz9bFCHPG/o6X6gWyYcx3TY
EbMhpzKCD/iBiwOv/HlYY5/4E7mT3cAu24dmOpJX0RZr1rckv64zZ4gWlev7D3tB
K1HOcblLX2zsUeE4yVs+CqgUKZUVRUfbBz3mVqPux0Nvqw0gcddu4UwX/n8f1HEi
vYSwrMVWHnFjLbHdrWYGYYTabsHblBgCz9HCcjyUQMM9AE5hLlmhtl6RnKcNRXux
NS/EllQUuuJg9omRIHbkdVB2Vxz82p4c04xfkXUOzEF1ckmG0cwxPxo4WBkwpC4E
VwXbki53vmWY+PVknuUnV53fSxr/Wqdw/2wMBvGAwEBONz35dGonVpwDSzwXInPI
UtwGyhmfy7oN9K/1mEakr7jiy0gTJqf260+kxeGvGm8bMtdCf1k8xDZinGqWFPW+
S4BNXHoiAb2EZn/qcgaXznqBwnFaESymENPqMM6u5F+7/kzMHanL1lmIwEf46F/I
fAzwJfjPoHQ+KrdfidtKa9SF51CqigC7MQGAeFBpo6KwIp1qEp4KhgKgFBFi4wSG
WGQI3hQXsGYEot2LSf2Ffbg5sDrgsk9uWZ/1srFrL5U=
`protect END_PROTECTED
