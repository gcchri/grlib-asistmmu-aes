`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
70fn4xHckz8If7y9VLtw2FXZSua0gTk/H9vXy7aN19+iN5411VTQZk225edf0smi
wCcOn6TYfEh9w8aeCLeZqaazOpDcbg0gMpBm2otk5HnwpV+JEA1wk46wis0z+iWG
zIPgs5oUoQC3YaEu7uCDKMe2Ws/raoia0IBSJoJhTzWMBB7H4larHi2O/L1PE+se
ygaaD9S49MhAYHYESNnjgvfkvrZ6zkJUOJwl9DWTTWfvKaoU526EtoNb41uE0Wm9
87Qm7dBhNyjNkkoLjEvabLtljUfG+PEnHuM367KH1ft2ItE1xPI463x1o/GvTkR3
iyHlTJtYhDxZ6ccEgIqytz5a+HqMIhW8VU5TDQPAL0EJj48ldb7s/vG4bpvTMJfn
qi8IGp7SRr8ydjxRTbJwCQUf/TnPHR5aMeJMucmBn9GzWQcgvAfuSmp+oDzl2AKD
+WqRI1XrmtxZ+NplYOCtKNAKyiFVkLIGt7+7DYP1Tk2ZdzMI0mHLzUomO9tu5g0B
DaB6saZV2HC530B3tdb4yE3FjzrDoKRHXRFOIBCpQLtIeIAd5ZtT7lp//oTHz+AM
P8+fYURcYcM9PV/8rw2bvizzLL8lD3BjqWDkNzr3fVWHXth2p24P1uvUypiF5HHb
BNYI9dVoJzAc1VbmhjaZiBJn1TBLRUPFl7FBTX+tCBX5sTNY+JDn4eup5dzhJGTm
14pFeWGPtRFvMruxj7o5kq7KzLE7MzMs98SpQZ3xegIwpiiA9F1z4GfOpLia0ToX
qZiuszU0eNkgs7ew4zPFOCCv2D3VHPM56NxLZOhqFlEu5c8QMiT8f2dRWHbrtgiU
UMUE990YsREwKUxx/PF5Xy5tjd57WdO6IlWwmPSEHaqR6EY0bHup5knWTkCFQ+3z
XHdABP8Go2yEgMtCT9qZNPE6IgjRgu9VHoRMNeHdYkqi0tOKGVi+7dhx1ds8LiIy
CvoROFJhvampxH56POCZOpJDqXYt25DNSSkQt1vftjZ4tFGZozMZAL3y8k8yemyB
b1fezgu0Dyu9i7YgOpNJQThgjNxcYYp21JWRGwLWtli2GUBVvvQD9Y+8PrLrk3Bh
Y5REhYKIWVkphWmMDwKq9DEbj+TRodxmAJdMmRIdAl+z2ilVMvYLJlLX9Lz8Phr9
eMJ95IugR0/jxwxDrUO/FtqVxCUejGWYED+vaB4hXTQJBfqFmzaJRRYElwU/7sLf
Imr+8ful/AWpg6RmROuVhAIYXUZ25J+k8bqqFyy+F3juXJCA/jBdhId6yM1s9Yua
LjWbtZQKluONkppWExcBgwyP22i+6iW5nz/usIuZYj0=
`protect END_PROTECTED
