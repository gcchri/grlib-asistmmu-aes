`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HZNB05SOuLVpN2bNclW2WuumIGtCcfHYQC1lhmjoWQDdAIVX00BzbXLRYhjfHavi
rbYdHvLyjgPs+1iNGxQpdNfl0iM9RQAe44F7d+porFCBv9qq1muPHqQqYrWuwFIp
kGQ9s9Z7Y6Ja1R7VpocqwPQRu02VVJHwXzr7RLboGhLaJRQ7A1H/wuauqbNwQfFr
o4afmtBjJDNaexndZ3zPEVbiIXpHp8OKeHqEAUj2cFgZMppVnPP9nUsCvgYTkAYh
tI9ZbmgNrXn7d8woE8N3sCm34eB6+bv9j0My4PZgQ5yyzEv3sKAr4o3pMreyZuWZ
8GUgWqBY0N8i9h9wgxu2FKTAC4XahElwN8z18t16Zz9+FnssRJM4g3GUY2/j6hFo
gN8iZ3+49M2iqtQILlKL2HUy7SGE/213WLk5uiGpjo3X986GYI2hw76PQH2uUzUg
m9bwfprCKQHi6oZj0ayCTUfgJ9p4Ky/rcxVQ/1GvUZ6M5/KnuXBgJ9hflGH+CNhy
q2s2Yu4y+nVarNfoWCrM0i75T5PK8AsdA6VyFde/KhAPaakQo5h04AuQXkL1DjtW
+DFsNMBodg4mPVndfGist12KjLKMMolsNhNhJi+26tBpM9969gu5wvyvB4+7CkLF
4qFOqlBihGH/GQyx32UIqzzFIOTblcGjKCCb7fSrwREN87BvhKzOb3T2huBFRGwd
REPH6Z/vG52rqoGkmjcc28R460NbtuZMq/CKvrOYMa9skh3O/4hx6wdTtz6u73I9
5oO+x+auzK4np1S7iOE7xeebE+Cxb3ulgtxlU0ZJNHmkMpkr0NtweiPDFMvLkXGD
o6ggpRmYOB7lhdsF5A4LDTMCCU5CLbLH155GGOuacjRK2Wk4AhvGV5vUGVw44Alh
Xlzqu7H1HmB9WZPMyP+ibmJSHBP01vPEoNQLH6Rodfnuo8QJiQx5Wte1JB25Kutg
omVrsKg39T+XVKcR0f9j43YpUAQHrgRR3Tc0MtCD2QQHlKFG2QU1+tRas/DgANs0
4qwerLbtYieHo44bF9ftEoEU/xkhrd0JJtpzdt5s5Qo=
`protect END_PROTECTED
