`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ED7U4QhbaXEn0+qJ8W7DgObIa+sr+MnNJl97ah5XeiyBbSkZut8uz4ORQhTIFeg4
wkBkZZ7pMPFzkRkFzsXLlpPoELcAVN4MiGcP7ovsXAiCyGnvvCYbNANZvqSVqx6z
OPdcGqZBbgzdld1gxzPD1eVwWLMsb95CmK+jGStu95cu7AFFCFZeft79eFUwoVbv
2jWtkg68e9+QIRWdWrG+gwgFpg5Zm4JPyEL8wB+ALBYzD/GxgmmP85P+kAUDXt2k
ANVLh1UkLbYk3JdGROM4UK+ah1On3VR5utSAsa3UmOeoBavQKH1rojIxWCeGO3CL
2xhupH9HHdy/9s5tixCGXg==
`protect END_PROTECTED
