`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S3W3Y2y7DkNtsHvkpvg85TWM0y85ZkfmZVU6dVH6Lo1QFrvncxDb+subuwx5jsvU
Z+LKBzOpSrfQsJP+8abegRAFHU6/dIjE6KKU5Mg5lhkfDvaXzUk42Rt8vovn+7W7
H3/uR2U7k7qERRjCrqk9u5c4FejMK6KoKrGh2SPfe9GSTUsXw4mZG83MjZbfWNWM
Mgh81RPteLD8nImDVMjKwCjwRaP4ZJh8lyVSrOMT4xyk1Ud9gKMRgzf0ydPEuEkG
wKrwNowX2MmplsAPwvsCCL05vpsbKiykOkD/bLJ8+tQLzb5oMo8Qz6CGElKOB4/n
mFwFe9cr+6RUAf0aAt7SkroEKRVb6FapLwbTBKrMDOuxP0J9UMUxZQgEBCArU5Gm
DVr4jgI4L82MB2jbpsjue+Z3RFiCM8ISo3/upqC2OJy//4WYUiAEPAHr/yxx26OQ
fy0uG92a5Fz991QXD5cy43Q/B8Tu0cUHMLeEgXph3kQssMtGky2LCue7brlZ6gkK
ArL2G87lF5JDVp8NLI8MZVkge1mMlhMzO0Fk928ErgW/PtMLpfQZcR5G1Sr3D+F3
3RAHp6LpmaZM9VbZwDKZgcv5Ewtu06fNEoFQBITPt+Vhqprue0lZfjt3D/Dh1cff
fj5lSzK6bQTmcPbAzjalFzbsNAtmvqd49giaqSqEX/cXKGOtDV3uyQZO18Ua2xFW
VgEBwUQsXnEpEygh8cmisoV+8zk9jp6aTpjpkGpcxtPRsblf0bRCXehiEf25h26q
N819mJ4SVd8Vf18aIY2w27yuPDyecu46AATzbwgqOlY=
`protect END_PROTECTED
