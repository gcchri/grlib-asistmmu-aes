`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wdCvcByqL5EOwXKrFqvmF8jnco6Agdd9UAOLqrHFvnh5n41LPHf3Glm6SCRZ4WC5
YH1IJRm3ZM3JjEhefb+h7q4ApH6Nyx3e8+G9zVy536Gra219W9bx0wAazYYczCGA
e++PfYgRU1rFUMUXA0pjtPXEDM3+V3BL4Edr+7vhPC9YP6V8fYbynkyjKVGOwIBz
je4kpOITVkB+xaF+Gddn3qAGxq4vNQHZXp1tp5cscUZOjaAFi/dnrLyibHU9Xtd5
YOScveqvAVETwCvwfT33U7FAjVcMQ8pFjxFSacuq5IusLfY04HxmY0PZM/aie7ix
7YHnJBxvHl9Rl6vGLaO8tPIAFuJKHI+tXjyZ6jfaQ19Gzlq6y9Jz/cZyjttfqkmh
tddPPWFGVSTV15xHbTBnM7FL0j5UtB+BhMK1wDnt/L0y1DnW883NRPnhgS8dT7mU
QXCHjrZXAO4Y92EBr+aWWGXv8r+t8kPWLfiydDNfCLANeFDSRlO/CdZMhgAs7dBj
6bXWMNy4/xLq1OeB/IfCOIFFofnp84HVEd2C5FnAuil3s0WGrwcAIOk1NpQwHzcf
3Y/iSQxrr9BxbiVQ3s05XlINpwMt4huWxUSeRtBI2df7z8N0SYoBNw7AFyj6uJxU
Q+7PsF1ALzobBYpJiq92RRh0GwnnOvvKnI7LI5ggPZqtnMTo3tES8AtPphHt6xkt
aW1SaWI5PyOZw16I907w1DWhR5UnRdJy6UASTLVW939hy9oUa4P9NgmETf5faCSq
w+CpKtyK0u3bY2+sPN/7dQMuC96Rw4Pl19mRwGrEOeItBL8Qo2JqfxX+u/ZgKWtK
ZJR7f8ohyaQzBUeqHg3z+d2HLewGFU3Je7ml1CGgQ8vHjtial9sPvvOva6lrBUhY
CxgtAfuxZ8mFlK9MoIhPGHcvcTB252Ku5HG/4w4JRROiGp07GLhImPTSqMAYdXz6
5zE8BGWuKgdPIzBAJVGhCWpPeZfxztD7HJpcjF9lDChxx3ZLEhtlHAKsgRpi2PKA
Ik/VohOSkY2DgX0VmLrWzbzGXlw1LI8cPqfnxG1qoyJRISKiaROOqaAaszarzO8E
E0X/6q0cyZ3Oi0DJe0AIlPRU3usPipjxKy0FYv+8xjY6ZO5pk0921GUc2kVv5JuE
f3soF1xVZ2/V/ZySPLtKBDCXYusz9tKcoaMSBa6WLkIONtMHmFtwi4rmSQ3lB3XA
cWbzc5HviKEvq8giJmUzZziaqPyTM4DCJLY4SW0MzZqaZzzpwntHXJJaP9g277iV
N6hn7sDpBxZhgM9zla+oa0HPpv7m1C7JeEzI1z+C+foS39FV4FLYrfyFHmspeRJ7
5XvhaAuoJuJjTHobgbLzztNjH+Eyv9DRMh4dOF2R/T15qVDeXT0ej18IpRwBMvIo
HMKkhS6S9WB1U/WyITN34I541qIJ98p89haaDLC9EXmhpYgVrNaKy7RsMVCWObV8
gMKLIcYvvYFT3aymF6eb1GRKCFMoWoRyHPdo5wUrXp4=
`protect END_PROTECTED
