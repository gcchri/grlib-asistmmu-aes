`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JwzTcHMnMF0LCvzLCCT/hHzisDua08g6I1C59ux+PibQu15VFsXD4XnBwQdnTWMH
IDSnou63YOPe1P4oNbA/W0gBNtst7Z/FLNmKZLbNIp+CzIVD3tYKOGk6S1VRXTOr
S7CAuEZk/uFHTXdqIv6K91Wsdpe94njzN25r0od+50wgRDUIQOIRc4oG7rqidozA
2EhXEQx2AJ4T/oJQCQiJIEYwx93vkWL57pt55YBYM4XmJCz/+/GmfFrZNZccMh8/
m5YpJXkr/3HC5MGJ/c/UAFJQ1bo/agYmVOdMH8jsK0nhI4tw6FHORUjkigkDYUIE
mM40n/48orcuDah7RftrSg3G0c5dv4jGV0mwslImU7P1pGkI4RJFPpxvL0A5zx79
`protect END_PROTECTED
