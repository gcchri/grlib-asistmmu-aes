`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k6bkbhEgHioEC2z8eRbg+hpTDywC7yoCiNg+B/1T6SM4/K5qnG1Py0GqPgu+lcMM
cinhKxGEY++zB+sKOTRZWSixAhqxP4c+O828xTzT4oCwXxEmTheEjBURNgijpEYB
OysJZ9wYoAoA17DLTb2u6xYq1GDeG3qg3uGSk8hAMSTMkquAURkKeQ0AptLq4BHR
lPmSnxX6qVafd3XawDGhCVBvGcAYDO4dsukVCo2u+61fK77+7LR2q2cGLFiY41WU
as3Vq1PNnkJV8g5e4/2lfdln0ntwf9k3377WFnu9gVEIDq8C2H6XviGx/tcJVulO
2K5CCbpF0zwS5yRc/L0zuLSv3PY3A8vy94i+Jxiau+vO2ITeqNpgWKGyWPC0agER
edMppxE20hPwNuijRhAEhIVaXtfQZW79cXIwsigN3Kg=
`protect END_PROTECTED
