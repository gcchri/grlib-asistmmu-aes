`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f/mCraj1d6KMK74VMxus99PCLQrXC7JYs03lak6kX0Cj9oMGEasgF+mH5IpbMsKo
0us1g2Ct7KknfxIDrixthqy73IKcrfKGPXF/hi5E0Xg/Vp2BhkZZk06z9WI72/a0
pK5krrms0jtTfRF4n7q+Ryax/a3atkzQB/epKsF2KLW7SCHi9ynmHWBu1wQENuPh
eIPYOm+HO5bQ8UVfm4hX0O8E82DDFetd8+hzgjnpmvIsODAUziFBO85Q8pKSikV4
lsyQyJDpdyS9aBgal28m6KXVt5rrsMh2TTl37qPG1sju7Vm1mkYbfX/q8BmfJqzS
1Dny7tQE6bXsTE9wjF6fDyt34l5MJZU+6svywy92mMxppDRsvg5qf6H8+4QB2udF
leZ29OIzHm1nspR9tN7j38Q90dLwSQrDTmuUr1XmXvCwbLbJBBJLV2SbLEwCidEC
DnnZXMQfatSRTTUFOuvaKdfO2OnuRPlM1m8pMm12kuWFt/XqlQvpJBj7zSWN/cXh
PF92BwAdYT1oOMBix+9THptgbkJfkn2d8Gy+b9kvkOAa5/GuKCRCZlNtT4eEIqs/
ewUugnrMIRcqvkyrERhUbUu2o3TMhOTUiiO6fvOrH4bQxlghaG/iFgN9lK9h/Xx2
TaQ83FehBYC1d6aKJ4ayqlK0/1jSMKmW4piX87afy1P6ZhfYDX6tEdWHy6AeCV3z
XYYGLKQmYwU9U8wNFiyQTx4YoBdRJ8yo8bHzr3xbFvG892pIxc9HbmyCUqk5fRDU
126XhWKzotSYew9YYBJHeQ==
`protect END_PROTECTED
