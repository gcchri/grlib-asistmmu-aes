`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LbyYpElZYizUTME6mDxyOGwqmiM6KSt4e1UR/bqHIEax1hslkTTtXBwmW3CYg+YD
1RRt/Ky2eOkDzy8M53A2H7Mu1R/kupofbRVLjY2w1p4/JJ6kI9n8XxTPQKsLRhGV
sfk2zm+/HkfxsGUdUfWJY5bXRSxKfLZzwOn6ij+tK7Z9ctoCQx6QnRHRgKrkHFB+
yV3ea4ZURL7GiAR2V9m3DHs+S44acau8v0Xy6K5Q7QBZi2TYd0Lt+P1iM8xolm8k
aq5nARldrppMOwwgtXXva4WRrG2MTgvCn06jKDVX4E2MaVF6QbbU6HKY44rV9qK1
WiPKy39BsxDSofs5SIsQuELFisrGM55gZMjlgJx0tcecG++guD+NBPpumkVmdxOt
tMxDqmQ9hw9X/ikDn9PPjqibNqYhQjnUjEZWrGsvLrM=
`protect END_PROTECTED
