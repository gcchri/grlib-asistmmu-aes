`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A4FaDYcDFuv1KfwDOHG1WCgd3eppKnGgyIBDileW7Ag0Vz1Lgu7ICOPQHeCnCIN5
fk39hXMrnIYAez4bkMudFnjVa8CrWpcubXwOopg+fWIOprywH9/kf32dEXij059I
zKOiDiodOgLwRHHtfkt2pdW2oqzwD+KyhjiPg0woBNNO6caeidWOTZgdv5iqdBhk
JFiT0Trv8bcrYZfamMcGDZKXscRJy1Nw4kmktdUqo2OQg1/M+guiBUIICixBg0z4
9OpKbHqMnzQfV6boXNGZwjynZ6epRapdcctLHX3Ue1lngHy7cwrGa10UcBf/BOmJ
HLpPU5lg4mBPsjCej2/9Xglgj7uvvP57laSgzj0GPF2F6NeZsXyrSlBkxXhxDQhf
T7h1GFpqZx3x1ygLxgvVxBN75WU/k3SFw8hRIj9EKK93SMf2tzxhOEpPAT2jQPVk
x4CLZQ7LKkmK64dSXHk7YpT9fAEtVmUO1Pqdama1y5NC3tKT5lrHC/2fPNc+QZnn
Pzv6ajoFdDfKauCQi/maXNp7M3+ZvIF4CbXoVB4DpOx9yfMN+lIg9khjU4Y4KRm4
MLAc1+ztmLh77jAAioPCiSnWhpH3b490krP3IQ6X7H8iVVZ3BiZavCkFDGkrUUek
vfk6xG0U185cN85eTXKY+t0hAmf/uuigPGJjOtjibk/9F+JnTtbcJOHBm+g71yVX
fb1O3g+KgORUDSsc9PajmLBZsYQsZTbr/4B+k31oztkOMLrnj374/FeAQruXzb2y
Mz5CC1NiMu99A/yuROPmBynxxI1QJ/vQiDLcr6U2k39t11zFbxOQMUJeN8UAh0pL
1XssSWmZJ2OMIKDwqoHfMeY6gcCdFb4oZeN3n9duXFR8mmqPIYiqz00kObGO8qOF
TDfWNkErot/3RCCZPLsAv8U9gPWcmR0qpT5ROUEJvqAD3GvDXS0l+fp4UzGxA3J4
npyI5hyOaYAtt+e23mKadkyN636xyqmbnsc7BmZv1s2hWGTNmeN1d0ML81WDiRaH
qqfUd7GMH717sqNAVlj/WtsPyVRIJJW+x2fB9TtQbyF6uYf1NHNWuioGnVzIdGF6
4qYPZ3bGdPtj1m47BQdHD7vVMs521AcLdouJq6zwuaaWebvsKNxq5gHXXGwc0KPg
NDQxhD5MoCfVeZEM4wxrc+UtasYPbzD+Mz7ZsXhKfJS9pIr+4IiET6UWGP1Hj5b5
wQBjKg9EDz5uaAC9ElgcQA9n5BtF8BVXy5B8n9GsGt1nz8Xbl4p+tXhePtSL0o+8
Od25cyvAOz4NSrwO9KeBwt3V2iyfYdrwxLG+Ll7cEm7VgBDqU1nFBm6pdSzGvqFX
07CFm/ajBj0tI7LgeAH4oXD20rxOZUk1I4R2qZUENIGpaRAznDg1+6yuip8uWDg/
gy0l64U/B1aT6+ZvL12HXt00mrbEQqPgLgrMcRRxy1VP7H7EEY/FSJWi4T9IDjO+
O1UgX7qdRw1SnxTWRlfEb0gZ680y5oBQ6fheo8JKbrR3K6lLtMSgyEXG17eGa3o7
SQvWDUpsHLQ2Hi8z3niK+M/hcEbVM8r1LoSwCXMWqqjjp2NS/uNvrGaWgLaVQgYt
26XYX36YvVruc766FGQvrZF2eIxjJRKSSYO+LmLDmPNr2h9DOTUwwQnXQN5PRI/Q
cDE/E+a9KfROg4nVYA/5jLFiheQ1G1QNWxqFT04I2heIsgDwdgbi5bqPoQELLgPi
vYUI2ri92I2aK0+fCavHHqs/C4uFFcd2BbVrayszh/XV4vSArzb1HHdS+9J9Fenb
qVJssVku4bw3NSlnWh8fvAbATcTzUTFf8z/UI68qsDtgU7XVH635zuORUv+4fvmT
+kDeTg2E5gr+ZNNsvVlwMqg8uPDwn1V2B/fzqyMAnQceGFU/irzaC48A3g6Nh2jN
1/78kjnFl7/6hAzYpvSXxhwLBc5piJBF8PsJ0lhOu/0AXicQgYzDWCNgzHZtp469
ft05oUTAX3fOUrnUOozEMFjmw0NbMOsu3x/9Jjrp7FVl7smB9Ho7vd/yJEVfaH/P
MP3omzbBbbn98EO549KcZfynCv64BxK/AyAj6zAFf8yS3Z2ZBVWI4Oa2WGtMjtKA
lm7pFVg1P0FgnaSK/TVzglXYU5HP2Z96Pl7wWBRDfNEPLcd6lHylJSTefONSsLvt
M9tCqCmKrhpCzP23mG/WTqrCcEntQquUf8514t237Z8kb+a0nwVNLV5lXkkmFfeb
QQ3lCNcizoXUEgY6nF0qyQgQ0x1gH79+dTRwFKSN2E0Uk8G0wqxUTv8Gzl6Qm6QD
tTrZGXW8f/1j205yn91hvfTFxx9OPqCvWic64R00q7930xfXIPYq933iX4y5jpUG
jXjXY1u9V0sjIDjWLaRi0973UOKYhdutGoGa3wRdoAk94TuvpzHp6H7u0XHKBFCV
S36PfRGr8XbXMFfUFtRs7tO/empBTc+UIbYcSv1DrlHUAH8j9nShBLD8IGuSU2nC
3sn9fMYnFiSQo7rxVDtATAdwGo3BTkUtN8+TXAWK7IzCEaMdsXA/uI5R9HGHHoZK
aYLimwlTXHu+MAz5kTVEyidmTrhBynIUK4/hmY/2PqOdol0f58W6WlIX0FkQiTAs
uLwuY5J01+OkQSMHKL3/TH7Sr3bw56t/xXjobiDeUXMybI2qUA6K/syobTqzK5ok
GQRs9gfE25K+2ER1S1wfWCtRscrGrwIRYAtkacny7GRLFoHz84ALXUoct5qoIomZ
fUhEsClymOGCNRzhhLrdy9iwdjHOzQHW32ccyY8sAGzCbxyqDHYzu/u5LVhYxAaj
zU00jXEFHHFC3yyuWpC4gvVxLZ1MBIAa/xD5W3kcau9MHECVXHfLui0A9/YTAUNA
CeDydP7hN83t4ZoZQ+UYUny8C0WvxV79DjV4oJPsGnWfdVxLMg6VUs1BT/aktrrC
NdfJPy2yR1dxgMv5lTtW11rarpwg7TszzHrgCbyB38VX5FxY2fJYNHvyAm+LvICx
HcD1SYwO6RhKWo0qX+iyfTCFxAgCyGI+refQMaVg7HlEEqMjBoAG5yo/Y5bMjhh/
haSHDVUF9ugyOB3L/zS/wio+GMvnHsJYzgRVDFv2veXwVZhqsQoZDr/IXoM7Q+tE
8ycjMha7OYLI/rE2VhjtWqU8xbNHE13AiXRRCNhJI3Sci+qrVIZBdtbnCKrSyBV/
770NYbXXpL6DYnhNUL3iqbIi1LotQ+BCHYTbZVsg5DZ9wvTykKvS1eRS7XScOVgX
StYglm53MziNXFcrpOYWxnuyOEiLOhOm/VRteE52Qga8K7gdBpWfIp3m651VTQlP
g2PAnUW0DjIJ2Wnz3r71bYMN2ybBdgezPSlSlKT33oA32L7z3KFClN6zejBfTPcG
pKikyksmcEMcy9l7dKEBTDAHNfUn4v12wKS0A3ZHoGvWgcazx21aduv0BGhC89qc
URxlLDlNVH3jjSnzQwqDPOXfuTSTqNzrOHfxPGoa4SRK1m8/CmDt1w/sc9IkT+M3
hakugtG/vfPiAZ7YftsUclkMC8brBa2YigeLDRjmtDmOhMPvIlq3nqkiZjWvzJAI
cDnnLrwZqFSdS1Zw7oVhbeuJydKwbmOL6vK3vWlz0SdKjEFM13vrrivn37cv/aKp
tPlmmYhrtnkCfCwk4LCAaO7cyLLT8H7DvghE6SeIJHP3XTJB6TMELNf+tqDaqN0j
YYA2roF9/h2sJxwhDFLVzF+iqD7J6eDnYYbiFNWJMrXk4yefwiJi9NEZMDiZpv+M
qaFsOypvP44MZIGFKcdeYq9QQOJUOc+Uhsf24ZhFBeNyNRdvisL2uPmK/qHN/Mc4
TGZxnOm104FxZQn3ZFp4gssV2s4b/Uc4rpk30Frl8UWhJd09DgU6GA50A1v3kKUV
BhjyZJy7hr+xUSZjBmkacGWHay7XU51Ui8QpayospwC7FcXS+HsFPc5XkNDrel9b
+WOxLwirCW/kGQJVjF7MbEa5ru8LMYBiyxEoiMkvoe4nZHA8NxqUp00yCpHKXaHb
8dB0xr6TL3Gfgexm209MGy6bHaxEIks2Nq4gtoL3OPO4QBxR7eopKRHrGxDUg7rV
KRhsb6HzyRhbWUorXrx8FPYvF2rQ+Sx/kMOEsbFRONdwl1AOcQBPB/NQVeeX2lkV
pAwm8Hj1QxAhzgCKWSCzdtHdubmyi+CokoJ91wm9D7d3UV3q2tzbcWtiGZHR8YFp
xneP7/wNq7Y5ZgRN9RlrpvoR3/qpYsF/WJcrc6IKT/0PpuIDWZyLtzWMwfEndT2r
YIA4IDEHSPlkEZpmQUylSgWooOlA2ga9T3yFGs4xt2CdUv6o5SM+9cRI/TJVDIb4
9t9Cqye89QCcIYKqJn3SzXCBYnP2Crn1SFoxLk4f57m6BQFzOpdTHWtzhzPEmI8b
VI8aoqtSZTNDekzfUofkS3K4poR2+QMoBT0qH5kLUNtEaSqlugzP8TJttVFucCPx
c5N713zy/4fyJjU418WXqqQ/1KDVwg7pEerE1ohqlVtl1/TdKZPoPkbQ7cLvbChd
pa6qAudz+EcvfnMZuxldtgbeDIMl2iquE8yL+tW2YcpbDrXHwCbFKoTkBnGKAG+X
1aDaVzxy0rDIsxA+3as31OWeKRzw36DZRdbTzPUBen/kHuUlAz/AOj9Tfh+7HM/S
jsExviTPiQo4VY1XylxCEwCunKsM9Ii5rBgt5TAENzFj3McYg2ASE7QIZAi4oHDp
ZLTY4P/bFWp8leb7VmQf1N3yapMncWy7hsyJTXkYRqA/QNO5XrGfH1ls0aBBDp0a
2aFni9CjXlMSWzrSa/5XozEMP+0SVVO6mZEDBaNCbvdxtrXL2XRmCeEr24+8p91D
ZqPF33HEEgUodZjQBysxoRXqoTICQ77CsXflObtZDviPZ8fMGxuYd3zVomv6Txn1
Gl2lTq0D4PATzKSwPpQ+G7b6yglDeSfi8Vvl4kf5Pr3fIn+Q8A6IuWunFkzso+nR
WMdfH8Cvnl0njfTqTC2s33hosYjPtZ2CjtyKyGQvyiQtj/TBfwbhFGtVlbt2d74v
1EfQaCqAVbk+dMEKdlnwwgqCyH+2PHaIqX5S1Tdugfj42LWaj5zlB+YRiQjAa+aM
5/Es8xl47JQ59Xfca+iQdKikjP6IHkJmeFnI+x3cK7WtFEBW/0t39Y+PNsfzljpj
zxkSsfu3L6fpNNBnAyx1N8ZtfUCEUqjUz1AiGExsEEysECJBgfx7O1bdxmok8BQP
UtqG7yE8BJw9T/jDux8CCrpK4S68512scUNtA4A0wL4DQtaGjoWcFeL4kvp3txbI
rLytaaeeijjtZLx1cmkRyeT/FtjqjV7oqrECeiDG+tnxAGpZ3dgTVjyURvAx9yXB
1DcbUOlLwq/iT74bKLahneiCuZGrNXxYc78B1ZJm0BfGL4Y2T10i2HP3NBjqYE6f
bgAXep/0dTv4AqJZdslVk5QJlL7gQW5gK9Ghka9AgfX4dsXhonov1fcQi2rE9TSG
z3nUliub4DRS0zv7dwCDW0wOzNdpt6+1NIYpgIz4UIMG5SdRUrf2TqOIas4uXWH0
TtsJLupe9EKs4D08IC3yofVq/qGpETKydr4sFz81L6ybduKOac/uVOa6cIf9Loqn
0PhbGfEYd1V/UTAflOLwbAg3aXTKxqLOxVC/YamJ3MsMEB2NRrUHEqxmhX6I3VlF
9dS3W2oK2cc8aEDCJydpLfBbHQfZebvITs24KjXpKP9xxaaAVwYHLh5pG2a5eLev
2ilUnFZd1fZ1XhedbDXjtA==
`protect END_PROTECTED
