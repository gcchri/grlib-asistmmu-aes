`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NGWmmahoBWU+hZy+9hRfpG5bma44v819roV17bXD4lYKFulEhtSVndM9yRZLdloc
wZdtrnTSUjwNu3jdtY283al1ajU49KotIfut9Jao1js41cA0RbmMvLs/bpqsXNkR
hRg9b5nG6x2qsqV22DPVi0+e2jUKUdxoRyk6XyBqoZOR4fOhPofK8Rn9gcTo37/u
PnN1tvstqlIDVKYoNf5X8rRKoIxEx3nDiBv80jSWwuMCmejHmt8HVOi2p1Ej6vyw
nhzXybFSd6cYi3jjNxdTSw==
`protect END_PROTECTED
