`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mMtyzjPheT2doFJycyRDhcrhtAyhiML/gXllIewuukhrvy+enV3fAxM16ykMH301
ORMZaXeddT6f93agCMHS/VmcoIe+sUgS+KhB+eOoOuU4iyKEbQ7HzN3iXL0Sz67L
RDlEkAStdsghV46B7Zd+52K/5TEiyJuuieyp8tlxaVsD2wFLdYKVkfXAN/QvZRCE
WhJC98I9cdFWUgwCwHgju+J5853XmphbFt0MrPDgmXk3KRIfdTUy3pkLIUKL77hQ
2BiIOGPW+YZch+K9VeRu/y6XLBZ2xMeQfLBvqQVQmvpvq9z680xQdY/7r+//y/iL
EyquDQhMg2BX+ZrLldIUwFpzWR/DY47+PxddZOg23934pQrIfRIOMlLdOIb0UWkN
czIQHGp0EEGZX064xq/lI9jtAVWfC2SmYlk5D7AnhlNPWzsFpwrLj5D0y4tKNiLw
/7TlLZho5vrtGyhqh5pSPphQEsp7aaC03Bjw9QkWX80=
`protect END_PROTECTED
