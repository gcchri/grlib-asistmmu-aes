`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6hgVipgQyABobQ24TxWzql6wdEC9n8jSmbibziuR6sUuOZmaql4Gh3SfI1z4Tq8C
0IRHM255798lKI9qnTxhqFD0KvaHUpo3B0N3SQ91IIqZJ2n39CkFuOx/GsEPcDRc
lbLIhfFjoaVH2PMOjmsiIPNV9gvOoIn2OEcCmpB4rRP+KY9Ccpko+fBv5XYZNoiD
vmFBJoAIdq5bXnX+KVvESemq2UMFrcdb2p4tLEuR+rI+kBDo1a0PHXxknsSeGYpE
ecd74CsddBCrG0KrOcxJLWFk732eHuw0i1ve2FhKIWuhs/vZoyWgr9C4kaCJvLKp
uXXeFw0eK8jQhf4uue13ypxld+co33S3tJI3ibNb8AGxVo5SS/G3qOy9k5JEH9d6
iRg6W+ilt/x8XuclRwjkaRQf6FIR/Artqwt5sNFwt4tzKPLD8E3Cbq/DV2CqyNjz
6/Q1pfFcOcqBSPK/r9BqzXIUvoxuxXc8TJo56cH3ehFeFYloknTfz6ENekFGOsDd
pYc0dHqATvoiOcXjmuownXBZUivreC1wbbezFl8jm/AWRPLJi2uV+v0U+4525M+W
6zhUf4jGL+5e1phaNdha0qFSis6esx/TAhQH1c8IZ5PYChIHebjfik3/5qymbzfc
ScCt2dJ9q//MY56MsrPq5bFn0cRvRWp7KrtG0rDjqLci5jv1DHPzp2KRGxjV8DQl
2UUD6BezKCtmv+x9NmmRnq6UpbCqU2HKp4d4PUxJUdZenaQsnByvTCydDO6UJnhM
Byn6efZTlsa4Ly8X6J5gcHsEsjmT9pQPxK1pA8M0rwJNLPU67jTurhqcHqKRGck7
`protect END_PROTECTED
