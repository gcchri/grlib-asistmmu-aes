`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cHs07tlDyHhiBaWrJKZLVNKOIotJnLDcbiKsdrdjdFqOjtuc0xM7h/JdlQ3lQgPh
pMGfrasABG4MT4A1h7rVsRn3D/BY4WV08tpy0MwLsuNG9j2avhNdNNO+NMpMZv2z
iVHV5W7Xr/1OHi7WY6hZMiTMrbVuKnjMXUz2pNh+WfwizG5ydykMdhASVQQea0i1
cMnTUT/qOKcy52tqpKhisKq5kVHLi3sa5YzFUs1Gh9h2QJ4pz+u2+u9S9PGpzlOj
ZgcJj/dLsTqStuKUuZo19Gi/v9/LKaGsdB2LWEttHbx7ihdaLhTRdTTn7e70qclT
C9gUetEG8EBX9Mj+XN01TH9U83MXS3n88efnovPhF78MK1H5Whs1akJ2aGcXsw42
USDdVCKCzHX1Nx+PwVCU5GBM+URuLmKsLsx1Cr/PGQSg3ZgfnC7Km2hY/y9v1tyq
pxBOIgwg19pxpW9kY7in2hZ4iNgP1Duo6iCQ9ub8uCpGgo6jUyZjGK6NAZwuSolQ
VCqfRF2z2171NRgMH3qZJBZwaftVcTp8FFQkUcL1+4c=
`protect END_PROTECTED
