`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jMnyQy8MYNz1J+1WkeK9ov/2SYOoBidHQIZO6GEVY2cZ+91vvysS3lOZni+YTTLs
wwEvMAgXsL9xnLqIHSwfNAp9XMBluQmC9PiGnH4SexYBmRL3hnwcSZpJ3JC0K4jN
vj2Kd55K+Q6FH378mXzyNWp5Op/P1GWae5MGFq8MWDs6bnHEqdmY14Tj+5dVTCI2
VRAiUJVvy3pSscpouvrQ1kEiO1T2bQLDui9ihD/qcJ6hyBbHqfi/l74IjZ6HQqo3
9BVdtCfCkwXetysB4ehBdg2Q4tlfCY5qVk4vqedUX7V8v7Wu1iDNS+ByU/fZvPzO
4AQCSWvUJnSr/4xBwpVktQ==
`protect END_PROTECTED
