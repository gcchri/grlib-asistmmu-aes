`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6d7C0t/pt/Sx9DViCqy7ecOM8cg9H64utMwHOuoK/KhsNB24rpKPIICFQMK79mO0
3LT8HO/+KZvEH/mmTyuAsPgtUcBYZHr3t720MnkIpNzOj7OJkCvmXF5PCgRK0sly
J+Ha6C/s693zQUgsak5YwHgaLbnsplM8mTFS5E+FcyAkkNjoGkv5B/HZ7SeJ0sWZ
zSemWyg9Ays3iVUG9y5NpnmCkBFp1Kxumqad8bC5oPWr4B+2mXx9ldt5Bs653XT/
Ose2C60sckwwPRU++4AqA2NB5S+tZHx3zB+aVVDe7akVj1RvmJDeBmbXiPxvHVnv
JM/o/18FCU2Jx1/IBlDmCLHAaBfSyMj1Q8HBs1N7FR8/ME99H/Pco88GDxKxHl8c
vpah93UbZ9wZzppeK7r6U6sy3HKPi/xGbX5q4amfu2KIaMF0t5DRpG2qBk1cqNCa
yWDC1O38felteIt4ROvEPA==
`protect END_PROTECTED
