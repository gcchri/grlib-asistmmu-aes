`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+MwYedaXoxhjKggOuxow1yjQF2kJNdw0IUm7lOVraACQIdD1K5GtWbIuYWdxe5uH
s8u18q7fXHh/uD0MsoPBV5zsdCVXdIQCg8IGjOMpdoSgSIm4/8BfU0Ms46XNbSZY
1OnhBbYUqHGRKg3WGc5G1CHLmFxAfUlSwD/9/LkR8FEcRokEiIlb7dRDgxGBqAqe
iR47h90Yk23mYAyeoVabXdCDL3MlpOMy+3aHgwksqaGg+sjd6Pfjbw7F/qw/eYYL
jIY6MX9gwpfgHFa4OBfRYc72KqEPb4SHK1KkYw8UkIXRKzmCIp7yBzweT1WMr7BB
ypP1Y3JID9You06lkxPM4SM7kYjzHlAUPC+E6wwJ/ctHttA5tanaeWwwrftFCo39
aKavswzDZlT1CC6HKi+PvQcW90Qcr97Jl7T5ZicULyvljIh3XCvc/2iRmX7khNX3
VEOH7+f+4KfZ0LBfX0KJJyZQHqJSbafw44iYYVcseUboRtWcR1J57a2v7eQkHlJ9
/AlLwvKJegzy/hpc71Cs0HOfjvY8wAUH2YJVM9IHSw7ibjlGjSiJXpkxCtt/e3ct
bwsANe6wIbM6LDBm8dFCjQHeD9ukw0IdfSHWxrOtkSWfYmQDnSoOK22v07jFl9Hc
ylEq92r3BWzYrhoJE/5WJduHoq5IdOEPuCQffdzOdGeZY7EOjAgtuZ4MKmzHYT+t
fzacGHnK9WCYCFg309wA+JgEC0mrcVfnygSiMHD0R3DWyd+vQ8tDwShDWsW082qj
ec2c2xBSrTjUkoSzwYuh5KSE+LyTkmBiYDk1UGa6a6pDNJpcvZ6bfxtAKWfFA5QN
6wRKKLsRP/EgipRDtLD196pIHG1clFnWfC3heKhTYIQYlVSbrAIzQS1PyeweeSRk
hyXaH66iZdwp5AkUq/LCXJWHIRF4unBOmpTkesN3Zd0TXRvve05+NEm646jKZYww
Q8IK6L3q/viqslevCH3qQhcRdZDIGMPryEyxPj7Lf+gmN6PuNNP2o/ijK52PCPvF
4hSTlZDseoR17DQRVNd7/259ZAo2j8/ap2obEP0MdlAuz1podkBn7MLj0GJHPLTT
UvRU62CHgxKaaRPDGT4GlBwIAFLu/iGf91H+mddF/1eqqwxc5gPBioFRRDDAQYP0
XXys4iDFdV3s1zKFEbky2Mnh52qd28OG+2Nw+cPiQ+4tt1Orn7ojJTJ7oob353Hp
Pl7406pJpd6s/H4dtEOZmeEEv2U8tjA4iZHpybiOSrNTnjT/nexP6R9ejvogMv/x
48ffxe8eAR6lCgr1Lk3zIaBIPIDVcOdxadt2GVDfmLS1vTZnkpSXVNPo8mMt8jw6
PFI1Tq4+e0e8h6qL3EkV4/I5oAiEKc5y6mNnBhSbGm1Bethyl8EEY85zqbM+27tc
mcwl7lP1IyIhoC3HioUyrF92xuhXVavgKNgVnc3SXkVd3vdQeWZTS0++Foe3C9cv
HUDSb40+aUqWRfxfKFY4pv0rfFTJy5zcOg210xPO22S/xIIleyjgoY2xAUJBUyUe
NE9hwCKwUuqZcVCckiPkNpAU4m/57BMavk3F3jo64YdbORz2LhGZ06iJU8yECWrX
7dWJ+SHvf88SnuEG/IdnVsrqS/3TWpV247mKMpZlRUBjTWbaTdzwerJ9BkGzuDsJ
222V7HrCDZ0p5oCUCGOS2poBvwTaii3Sk1M5gcpWTBGpgEopNNpscVs+aH9tmGyM
3KjU7vfrsIdz1p4QydLWkR0fBhKsAm7j+73JkGDn84TaZ/4Ed0LKAKtkeIsABgoJ
To/tASCPEDiLQ6Ty6ielr5KvE9Rl4ha/ttHEgia8hnGuObXAeOR/mvthmwF2BGGx
ZL+ct/DM8uoLEPVarObU626npvnMF3gb3INKbFM72pCEeGlDvGn2YlCVqb26rP4b
WyoQijQ4w5ch3g9qsS2QJpgCipyuXOJ8sZdnowsc6lDtlpNHBFOZd8hxI/060hS/
pVwcBQr/K438ysbXNDnJab6YYltKoQbf7GpkQ38u1s0rBRA2B5mBZcfmQ8ml9YtQ
p45vgQ4/4L+zl+wzR1dZVkQxXJEmc6bRMUFS5NAlzzqf5a4IjZnc8M4RW8/ZRfOo
qRqUSwI1kCMjo9FMFQS09xxsdbvFMyT4BjPDxKzHFXV7v4Pc7nLwNJdXpijSXlJK
eGMxQzypkIPifR1alNCsOTPQR+szVlPV+FJfN5TmROOwcHWQBdj7ik3y/TPNcXyr
XkitYU6ifRJDvn92d0DbuL27KQdo8xJ1IFWwaMVQNFY=
`protect END_PROTECTED
