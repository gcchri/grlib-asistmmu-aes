`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/YugNgIO2ihQVNrXpRNe3TPagt+bjwR1P1chTnsyPnlEWylA1ynE0WojCOn32/26
I576Mlx5T0izfovoCimzxgF2LNCzY+pNZmp5JaON8lAs9UBo3JExYRZPVePHERrt
+MUU6Yfw48jBmDBESdqxX2TDrCucndC6uzaxh6HXHEJJfu1MONtpH1o8IJQvklq9
b6WX1mYB29V+JWLW8P5iBisV0RBVlu+vkuK7JqHiWQxbAZMviM6OXZGymsAXVUz2
nxGNHbP+I1hE9Gqt4PtmA8lx96hamJqUdAx7KlwCfXFGx64SPibFD6NTNLPxMPsC
varCwTgGMv8EhAsx9FkA1suLQay9YHgBXzl8Gl+LBJCkm2d1RUunJeWoIsOWE757
EI1rRqHTEI7C5xgfNVwld8WmhXBPFEgGwRaHKmR4lsyT1vjf3yG8hRKFoD9LNfil
3AcT7scB3aYWHlwmIzBOf0NjJck/9QhUQDI5UNMFsXfcAXeJwYIemKpE/RB1WTlK
gTz0OX0xIH8crZnlhGLj4quHIuPNwjUFDRctXOJqW0tVuORBUrJmLYGmWFixxHCn
Ho/vWp6SNvrsP1ibToICtth8pSbnqNDgVIvx8elYjDAvMFTTE9hM38WITp/6mjgM
xJkKxFn+Q3QZR8RRAy3ZYgm0B8yBqCMtJCBon/7AvubrkTQtFRQur9r4wnwbXDju
hEYQ1g1YlESKxjeAAL3/f1aacMwfKt++Tme0kcO+X3eON10TyHvo9u9L14WTUUWm
qO5FRYZTIBdFPmtIjmvZtzOWiKHNjrlVj2E0l3tDTGEIhZI54tUZRrJMFL+hUw/R
qfckMEjLeY7cYEwX0KMbtz9VElCeUq7sAFbos/Lb206ltBgXPKHxBW5JfLuCVBeN
1ZnLBiqyUIqwQoJuiCndWO5Z+4bAWW8o/gtauMvetiyDY2lo0yhesrHpAXi9tc9K
RJ+m6xAaiJgAiIwm0oBOznVT2vul72yxHlamGsheAnPClm7uh9PB6G/QaWw/R/ES
KCCorbCAPmqDbUroyjTlbSr7pXWJqFTxCiYjQAOzIhso0aKzzAMNkntd2CtlHyNn
bVdKiEm5+fSH7kY7G6B9fYJZQbIV46HWdpiEzapHxjI+vX7kahS7R7ExF7d1aKLR
IJ8fGRMhPYMGO7v5KbpLbortvmyT73AqF8za9AQaxcTqhf3NuhS4sBgqOghQUnT7
a5+/6kJ0XHTY9VHFZI8uo8zpZKqLhp9U13dZ+23f27hmtrtphe3tMqkR+DV6cokP
xSt7/0X8JYjIZE4Ok101r7yI3dzChKtbomTrshTDAUxZH0pjwW/XkLPwSWTsvsSf
Ae2p5byzanbgcJn81pE2UPIqbONqSi/3d+Qj14BpjAwMVWJms3R5+nMS47sNY43h
PPvJF1Nb1WiVZOXtg2wNuNuMGasSy0nvRP2wvEr5YABUcW8XHh6/bYnI2/pZuA6H
Br6oSaDM2gAq0k7cYSwM92ashVdKDMKgJHmKLN3w3xwsT3H9qGzGuVDsudTo4d0t
XFz4hIvMHI+Ai58KsrWUHMJ8cHKGnJVp2Ehopfz0dOQcmZMBF+REnTArx170oC0B
rvW9mT2/GGnjdfbTSW0afK3xigal2warreklsjDk1H4YOzTLrYDR5c7CYuPG9V59
N11WT/6PB8rsj6enhaZKAq53JzmxdwkvexRqRPyWaf+JbTPGGctvD/xkhxPmTBQV
81xxlmkDPw8r/WphEsuJJNEsDLtbDJjHS0QepL+W8IzYoCsuxApKjLSVl4r22at3
8m6UurwD2yFJ6Fci75/a7HGsjU+yWkWpPoge/Wtjm60pjy8ljPt5fs61kmVdyBMC
nfn7Bs2Zpnk+DAfaaKCS15cYROoG+Rv2nsYRhwvS3pcKB4zW8SQaunPyeyV7cKRS
MV3pMDzrgzrvjVHdogczHS624CB4couM4TPaLGl+32+fvWOdv74xXGiFt5yZXKgS
OMsQRXFgW0cTpMzHlk75OPueDxNF5UimgYLQ9NkuTgGQN4k7EGmj6iMp3VZZOkOP
aqUHPcv1r78d7fpYwNj4qVYSemzEwrlj52UchR3aqvK7i/Ryvx6wRgdWHY1TnLEn
UH5qvYAz46RL1vvi+/dsVqYo8df5Rf/5PWOzSmMqBsm7YAfu+Hv9oligVqmLHYXg
H99B+Mke9sgKPJoFB7lJQ+7n0KdRotweqH7MAIzT3WX+oMIP2GRcb3ATGMunDvCi
ewRofD7FRK4zdKWbyVcHjN6oz7GVzghFmwCObOaBFK4HUnncb1e/JSF+6Xrcw98P
3gOUQ215QIXFNQlIkVIGUxdOlDWl1kuJNHYH8Z6DsrE2/3Km5zXNGlVoElHUXUxU
XXhx74SQrtQBgFduSw2XPif+dRbijDBVRX3ER2M6qttMiJu5PTXU8aeopjj+wmxL
Pz99vWUsdFuH9ZkNaszeCQ1l7BlOSbAW7KlIfMFb1ObSe1VwHRrIes7CtdcFACDe
gs69vbzznEmAu1AwXs9b+iBlmQIHF8Tspppd9yBf76gEzm6lmz2z2Dus0qkSFa7h
OJtnosLFzxqyEzUouxESC3tb5KfkqyydKfc5kR1Rj0MW+QUY52mFkAVJwA+DtMkT
kfxxvaG/OfwWN6lW9GwZq+3gIRvex/VKww2ewjiTHOtUowPnrMyFoh5FDDX8ArCj
/Fe5vRpj1vxqRTuyl6Pf2y+d9ePZw+46Px5TjuIlf6cne/+/TnQz5T4OtgD4p5RC
Az2l5d56nh1DGBB8Lh3LAKFn+cGPX9i43yAFD3Rg352swcTc/61Yys60W6f3lEug
fob7t5LM5K4ov7HnkafaUCtc+3GhYXFAzZLTgMGd3FpIIr9ONKpr2wzfbiFoRTlZ
wKJKQs300un29UYdo2Eu9RerztHzs0pzSxYPSkTGGAZyDUg323nl7Bmv8NYdIGdD
fsSWmhRFsIZQ0TvotF2/4mHMqC1xtBj2jE02RC6yO60wWrbKVVAcBiEko8UJOvYK
vxnfV4emCPD4AYc1h2ANC4LCaZ6zwJL3xL5HUmZfZw2OwU05JD7oZZ8CyIoWGvHF
ysQcCH0Dy8NYweUwaSZ0WjwAWFPoU39b5Ms9yQvrbK1N+Jdssqzx34YXQjVByOpM
fmyrl+IoPmAxrownvqh+WcQVU23vcNx4iJ3UmnsxBUMzXOa4CgTpfajsXPfBBtdt
vb7MtdlAVdBz93sv1OTBeplVp8hIHWBOlF9kUxlYCQu13W3a9BMPN2LXsOKJCG0w
reQyhCvymEfsLNCE76kjn7B4W4Tr+voIiHOFRF4hHClPyTMvkd6UG4D90GX3xVR/
1roiQzPbzca2v9ucm/LMPAMxoXUK/dK+BPHIm4P2SN8bLsgMGsSJLKrfpo7dlqlw
22KNBC3/qrWzaMqz4YTGVfBb+H1K3eMrLG1+dSQcsz7vixi2rcZNrCU2avnqtYMN
TK31KtRKbJIJ93k6tIP5eblEh9T8EKXqIOdaUDWbcyN0SVziEiXU+KFcefMVUwUJ
m1DwarFT+1cMpcIc1yVdFsFdwV0xFHZnBAwh88M4c8QmNHw2hAnlUSUURIEwWgD3
bydC7ZUyj64AZm8f3YLOcmXn6BI8PFxwnjcC5Efmn+8OBTj2kTeKtZ9j/7w3BCYV
nYao05JqOonMDRKNeqUtqpUYBee1KZA2xIcHxgqrwQfzrRQpZ/Fcfv2biNpjZBqF
EwaTEdSDxCrz+T3b53d1kjcwJYaX5EodhL+7IEt5jTHUa8gVsq/KTeD05oClwvLq
f/TvDDR46HNTHuMoFuk47AcqAXtJW5dsy2rsg08i2vMelqbuEPy4eygCflsR8moy
kIvJQbs7zZZj9ChX7C1OyQiU93921CvPlKhTFuuvFRF+lcZ4Hby6w8MzZqBhP1h8
++rfXytdHrC1oNgXl1TBREF24BWeuI/Hpqky4s/Sy7WgEGg3dLuAcmffdLXmM753
mTisvG4toReeUhdPqM7G9gRWK6MGmPVUDVCZadSJO7WFOe3dVvVFsFXuFG4TGx1i
+uCDkFjT3aEM5ahI9ACZMjjKo0szg9pOEqFrwEfiDAqnO3aXcSphsRqxsWndPE0N
5F/TCGzmDeZIDzd4+JBeQwv55ZbhiDz8lspS/dyz7mkZMEeUmSnwWiCDeI152YdG
A64DB8ZtYtmQJw7dL+I7AsV4zAcUebQvwJPEdplZwxq6moa5Rl3adcyt3lWgWEhJ
lyZ0nxhlftUM6U3ioVk0aSsGHRPvx868yvJCt3gPTqe7T3K1yjbQAzSF1Zd0qK41
rApPIi1peMpzIqf4Mp3Ot+wHyS/nyj1RFDUKE556vJuTx7BBI3C3oQIV0HYT/B7E
aMqSJmJwg8dHUvXgfGW5r6n49HDI0/ztpVwi1m3XwM9XFZRF5qrBc0O6ui4lGILb
1RWHtv3/N1MeCLjz40klere0VYJTyfunFx5z4qf2wA3QKzI/vqCQ737B6a491f62
7YPNHBVpIcDG02wyrYXKOc/lB4n1v9dRHuOa2DUzZd9EVDarR46Gr1LfOu0Oju2P
mhCChnclf9vlrFsC2Qcm9Bm1rCbwEvnSY0D8D3NrNMUCx7yePequCwme4rDOTEcV
4TTDKRbMOY5KZ+0H5RsbJaDvR1E73YN6/f21ImwVktTsWYFrumD9ou6Jnfofysck
9WRvEaouHLTQKjwirnAn9Auj/1iM32FQen+S3Gb7zcVtpjgYC0X9pq+f1ENzQwwc
Bkw1qCjiT9Svwqm6gon4bJPj7gT3yY7oRbEFudixGkkvNUGAwAQ8R93x/AnJwN4X
NI4DnNmYBea3pUgQJ/5BNTjS/ENu8w3VFX0slfizioUARDm7o7qrtI5Fmhrbdln1
2SQA4eZoZKvnnIK5ltFJmY3CnymHRQt7Ae1FmFRWM527w8odOvTqMycNpvifFhau
IT7LD7uze8ZsAcI17Au052vAzaKCkdP7xczVIhtlFXsu4TM9hfqeHVDuuLiOt++O
R6+n5duQrrSi9a8yYUBytoncehzJ1Y/LSZ5q4fKgM1NpKIkqZQwoMLGGmDlBBnZG
MyVWRGPmIjKIdTtUAmv+xAfhynprgW+Nj8/hwjkN/ydhppu405gY1b5eW+mStoTY
uHIhqVdyuB+F8wC0ckTmw5D5wIPryqqniA0pBLszqlbRp/O0sr+N22nCKNBVqHXV
5VZxF1RwySO8ngmcVjm/rA==
`protect END_PROTECTED
