`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qHi0paD0JSUrvNj6i5bf1RkQxr9dSfc8EmPhayG9dVPEqMQVMUH8/sl2wNUJsvvN
k16+yGlWLvDgoNVIZsaXPI955so0eVv5VXMHu+EGpzg0JZBTOYyvsYlanHLypjyN
vOh88GxfOdWpkFoYpCD++t2VCu5F2xr7Brh7Rz4swk5lmzfVpVufONFNf9DE3JDM
wwcj43hGeKEob1XWZuc2Lkb0/A6RMycWyrtfSEcn/65FOQMN54oIHytmNf+HEhdL
AV0HzmDlr5oF8G8JLXBolFUpreNzXcV77Xo8OQrUfr95/wmh0e7iAgGjCjxlJeM1
4h7KwHG5ygyI59O208xbdWHQTTeMMg/Hz8sr95ONl17pxmzkAWaTsnoHjvmaBzmf
eDgS0L9Q6FzjKEVWyn0EzYBLdti5ZqT4YqOyxc86WP21YWxl4XdKEBcoAbdM4mSD
XWE5hRZ+37DAb666QHPibqOEGWhL8kfJYeyCCWRB0Xs0DLiuVTHDncQXpRLcIoJ3
amwxcUvnLL98GFEFQGqDp1hQ1O65RMVSkD0VQ3N4YTMMEeAbenbWXzUOgsVKEsMr
WjDirvKG0mxmInp/4gWagBRBFu+HSuJxM/SVLRLBSLEwE2ZPeW1neltUQlvxt2UZ
NIwj48eun+eUWJj4vzvVpVOCQ7+fz07Xf47dc+weAVRBtyRfP3A0TZy8e9wRonGz
Fyy8bFlzohg/sSQ9NOcKmlX/8ix4UfjxaYy95fAisfWtkScFk6VjdNMs8IBwkTmW
E0KriZBjVGEhiXLBw1e1ni22bSR13UPF/FcU18Vygrg8l1HHtAa6/2pyVBHEJY1t
IL7EPh6bBWBEl+Xh5rNZ1jQUvA9H4wreEPv8FXB64HX9ynKVkE7FSwnt6/H6oTmN
4QMYso/FLdDhyR45F+GGTO3RYqGRlz1E9pdpOsGMEs7RxeTvkV10AbgY6eiDEBPo
8tr+S/eHVpZqTJz3jWHKQq25k4dQnQFzxSppz7e+Tcu/Vxi6dr72YsTyleIIOVzx
ciCKxzn2rQEMWuyT4J3D238qZbfUVHZcb93/NhaL/y7J24cQj0qF3/Aig++avyjS
+Fo+Sgg6ShW9+Gz0SnHJN43A5D9bD26c8lbJLXt1e9ILcmKtvlkZhyBEgjEVTTon
7ye/k7WXZrs1N61O0R/IkvKFAx+0vWfoJvlMw3I+/gnMm6KIvM0UwRfPhP4ltYO1
Ar2VwFogV9crJzFjuVcnIaS1k5MjXNGI4eblvHMsOc7IdF07CdiT/oiTi5qmvjnk
AD2fQra97waWA+YrNivjmjM64NvYC7M1TVG2n7wWoqAhrZRA2B2Vljk8fuwlbN+4
`protect END_PROTECTED
