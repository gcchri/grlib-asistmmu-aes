`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jlGDMtdq8li7090/8EGjjmBJpl0WvcqZ+FVRpO222y0BaVU0wDvCQULg94dRM7pE
5EdfUkD5a2P6zlimJgyLdfu/xjjTNqDVvXShTjQ1o0IwdD0P4hEBRblU6MZ99DLG
S2whu3quyEBDD9QkS7yZeD/yWa1Is0ZvhqA+jFKM/ZWpa5lCaDEkMGp/ygBDOhbL
I/TXa6utD/KKkj+ywBKvOVXhNpBbi4cPtU27LPBkcKvD8pDZ/KTcsOdnK9S/RyTC
8JpjcjkGfHqJTVjbGBdcWDZdf60W7JMzeF/v3eiGUKd3T1/vYJ5ONEjH0+3xOD7g
JyKRcqmYZVYhta39VYx9F2FUiheCCHR1k3JEBZQwes3KwbZLpIiP2WTFNtLVSIMw
0aluyv7Lk++2htDvbqUSymrtjWzkBoZMjQsZxu62E+A=
`protect END_PROTECTED
