`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MjzmBArm27zqKRdQm+KZOQ2Mh+r0loJpSRDCcBd9HriY/SxjjbBABv6vIAjzMbBV
KVk8IhmFSo+lbevSk/TPObYJfeATItPwS4GIsCTjEK0f8kBS+tMkWz0AHCuyPTui
gWXzg1Ah+KoqOUo200bjFsyqAeb3n9G8C621BG/zY0Ko3VhsvJsC+I3wF7F+6f0V
UN0MheG52JcGiIB+eifGG9xmr/fZ7WkhLrbhSyGYxx0bPWN31WAfer38cvfnH/Uu
`protect END_PROTECTED
