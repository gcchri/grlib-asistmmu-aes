`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fXGb2VU9J4HbKyqEDDyVgIFRtdu9ugfim3t+oAv0sklWPiXbO97EC3/oOKkNe0RC
/oycwNTRzP8q7f3Zol8UIHf+Ugvf3+7BvcyyM+5f9ndZrE2J6vA5cf7sHUGVyHyK
xvXONLK2dMGd4hiHnfq5W84gXpZnOjxCVhQVMBUrC7CzDVLVib0GYLtFrwBk/qAd
DkYy+tM39RJ/L/7QW8SRWqTnq1dRf5785R9CNnN3a3uVcPFEkzo3CllKUfcjXpmP
py502auIXaxsbc+9OuOaW/M1hkvhYYPhtzj735GxcnzRX66+UrLY4onFRzJmK5c2
jcdUtwiYohC/n5Eis99FuUYxXdJyAnmyiFT56RTcDGZ/z+OxGvma8JO+W7AfEHiW
mJhmuAttkAwB3FLxmqxDbDGVKcFebLt1wlwC2YsqVKrn/IyRy7c91+qLh96Fo6kZ
RpH6UUNTPBD56dGOmuz7/HLbMevrMPL88M85CTUtSzAoMtGtxSMnbJFp2zMezJNU
lX6WjZqG3kTuOkUGgQgjBSEQ4cbVrQIHFh1X7YNIe48dEwB+z1qFtKAMeKkCoJr1
Fl4DZQH9sRQXvec+BDcoMLHWoruFTeG+C2N5+42k0yDuVS0WB2vy6t1RvKaPub42
9KDRypVbZMi1RVVB94CdTpnoRyyFVUnzvFN5MXhm+0jiy8JM2+xX3f2Na3ZYk4DD
rimqXkHslf75CaUmWCx4Jk1PCmZtFmXxi+kCzQDOTGX3vUW8pM5eF1NwYHEktGNF
wODLC3M4wBWMCmQlDEvZNLnQVNvrAeD3u5byDpprNBNV0oZDAtC9igxRCwkdRLa+
VkPDBPHfhX7aJiMgPqHxI1fJiQFXN5sI/TAf1sclvYY9js0S4RJp5QM/J9W5fEEt
AJ8rliKYkyiUBNSjYHPHIIxElGhpAA0a97RdO9tqrf9FCr/+qmjEcAEApQRlspdK
`protect END_PROTECTED
