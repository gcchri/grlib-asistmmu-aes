`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eOrm49YW+K1De/3u+O2cGSc7g09xnQ7OT9phubR27i9FlwBCe+pD8dxsLxM6lt3Z
8vV1wxnaPAsDatKURsJh/KmaS9+q6Xu4MGSsALzvfQorzHkgZ1wPfqE/PEm0VYmT
74oimVvsu5O+d+tewVSfxklR8CviDI6as22EWHTQK8Y2qr5jXctBoRigoYIB47CT
JYw02bX/VdxNvPoyXuIcsW4N3ZimoC0978YZ1QdscD/o7CIqmK+dXkMfEqhkvflm
+IWu8+yNo+Eb9FSGT0P+pTdgJ08rf0/HperbCBkhJIAirJbU80PmaDCrqUVcImrz
8/gVr3RMLppNY7KXrGWr7YqUxmycy45xBE9KBJX5+OtOfe8A26x1N3eep/MW5Dpm
2ZmkC3MHjbx71ZnQuq6oNiCVpryi2hIfI6JZ77CzX+r/2s0JqRo0r8da/3fZww4r
/1m9cj3A+I9dwmyPmUVvsFp91OqOPIaKr5q83W/L0cHRAUl6kQB8lFZ/5jGumEm8
VNoi4+zFPtDQeb6Wvlc9uRFnIipslE39a4HsiMHZbqbxehFGsAJJKlTAOghbHMJ3
AA9V/3H7B05IzEGhSc4UQPFsAeF1I5dVDyLiwti2yh26tlOVlRrmczYpgbJSKcOE
`protect END_PROTECTED
