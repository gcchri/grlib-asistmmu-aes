`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kcyu09IaP0AWQsf3EibBEa+xMfHuxlYwJYxQQywTNEwpdM5+fbOV5OnS4CZS3QPw
leI3egvNq6ppj7eHdLxgGQMBDgCBGogkXOrSSPf25dbfW5QDL5lyVaHjX+caTLcp
XRa+SK5W1z/xC+UuSWI6pTqrybl7pIUPlizyjiG/hq8IMwjmlLOlaTsZDot+asGH
fMdaMDHLem7CNliHp+3nGHI8B7WN9OnIKgyHP8F5YxCTn2fmrnDqukYPil1qRdMG
kZqK11DcSC4EyA4GRIEHv014T3ZEu6pnLKnt+ZOZd/4=
`protect END_PROTECTED
