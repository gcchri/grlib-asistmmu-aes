`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DUwH9j3mdfVp/RvLnHLPPEExmYqUtD0OnzAK9/pBnr0NU8BHb6kevnhCcJ2axom5
seZKFuncvcOZLnbkCRSCSSDdKql9egbjatNL8QZ26PRT4VeKATZIs0MCRhtyJZSP
0miKcNO2DdXR7lRevr4HEknqrKnUwExzNAC7gyo4+z/bPKMeAxGWwB5yTXsJlp8n
puu2NmpCHAPyL4b6QtxthpQ/CUqeIZB3ydDHfRBXMifiXLtI45D2oUh+5gyXl5y1
4hnDEjuOPj6SXVc4D/HSd3/nX4BRUfW40rUAvmjJcZTxScbaiZJKriOAbZgMS++W
8OK3lxHdMH9CaEdCIJ6kcroPGRzMhcqg5qTl8vPggQpCgw15PKnSlKPcS/XdMcWA
L9xyWOOQRVlvakzf8krKm1SHRCntGlwXv50nMKaVXm+yFGl+bFzMWZBrs7G4JxlG
BMr7eInXeeFeXbI6qxAvRMjih3hzYz3fUJrJA2IeN9YJAT/rk4Kj+00HQuZsjZA1
3wtuYdsAzTR5nzSAGwczFyyBIsQxXF2fEFHOP4acykwQ2RF8ts8QIdQoDGp3KBSI
6oFyesTOqyHiLLgKOoyXbWGCyd4R1IGuwEKgoovIKnoO6n5jmtlXipOqhRfl3kUa
7HpusNaWnk7YQZN5jVUNWZohF2iuIOpiaZqcWWqCoE7A5gUNR2yys3SgLI009+kX
kXorOiITn1F/Ix+GI5CoasPom8bFXJZehByXl2WBygZo/PWbE3pp2xp3yw8SkCGb
GqaCSWUbvkNTYhDNHS/g99/TZGb/Evdx4SgmaEurFGRMlDf0MIEiIvg5rwKYSghX
WnTn0rx2NxEmwdY1gF6R0dSvdPr8baMn/krHJ0FhakPnH2yTgDW7W/3dXHOuR83d
PIneBSUGla32WBnWKWVRxHRy6aR+m4fC9vZQI3+IkV91kauRBEZNdW17PcEFgXrE
52+z4fYRLSWN6+VoluPcopvBg5dIzIEIYqLqCeB65tliNWSZvmgx6BYNeugmVl5e
Sf8I/KGYJa4FfOtMgIMv2HXNk8nzf21OaTGHo+DxtjR277yanIMrXZvIEoQQ1KLF
8OATWu/1N1+POPVlXnRkOEkKOGhSLJJcnVGqwRisW5/2ukn49bCGqfiHAlq65Ugg
BGXPmM2C2rphvsR3ZmXMsxKinKEIbjMmirW3ROLCh9/u+s7hKvmKH6eDLnAoHQDI
gws/JbLbbEE+pT5Oune6cQpXzerdgivyS78EQl31tpre3++D56KKAJscOHO3IGbV
83uJnpkAbWPX5oSsN8q3C62MGJa7DxB9VN1hSfvS520KMdb30picjB4qtNlGajMv
RI8YgaYeL0IjhR01dep7n87o6S0RdNAwtuwIJ+oL0i7pNlv4Qm5y1JLxcIevdUVV
ZgsT1emorQPVcUWfi/S5p8Abd2bRNC3xcsQtelTBUdVrZzkZmS/JvQIOXJ2mBMGY
SGdPzWz3ILS2Xa3EBKzdihnOTAOpczqvVNfjqEfBLoJwz2gJ3LATAfVdFO43syBb
FOGNbuHTh3vzQuHz711MQ5nPqDDOFtxQ//CwbrJu7yypy+qJ9qlFP70VrNRtR526
hPXFYXkVpcEPjcuCLut9+BPMhksHHawFV1fdvWX/wN3qBWrs+H/ueTCaMtuhld/V
+jvIJCm+Q32zhA5og+GQEN4L2+x5x0IboMLuBXoGhREzwKalqtcM5crzym5uRjRb
7l8ZqzfRWqjNXuGuJQD86u1iLJtFh411cnDF2V9J3R7Wed3BVt+4egeWNqBV9SAP
Pl7aDUVnijjzyOk2JDG0pw7uiYb4NMTgRIXdVONui5KZXJcFexa2lC0Wusj6L6Dw
9xTGchpmV1ksX9KJDRQ6MMN6oe6rfs0N2oadtJtxRHhq0eH64eIZbD3NmeAxvhpD
zelJ+ik52N5k6P/APXFo/lislkBHbK7fEp9+vxtcP/RUq2VMlOYEh3C/S4APYdvW
QmBJfgBf+ppp8QU5F5vG+LQGXWat7DuN0pl0yUaaDOMEre5IEnwDcGTzbbc0v1zk
kcMJNBHwI3RvLUG0QS5Dw/aXljaDaSZUVIe3ahcg1BjjuMLZmdLZIT8GXVVAe9c/
Wy7clJvWfU9M5GP463ZirMLeJbfqd6N82HtFD3c0E/j9XT3vdZ8nsmk0hKDRGxgR
cXULrOn8QCkcQTUMXY52WVjPoUbE3YV7r/7AkV4pe4QrN9ObCneHw0IdcHp+17cD
ylfmfhR+PB8PDN30QGacomiomiPGGEAnw9KfoVWFh9RvabWI8aolhJhtl7/4A+2n
AJt8J+e94ATiM0+cH+DU5hPo+7QCbxbeEvfeEDIVA9+qeIIhdo4OijkrZF/U7WzK
k+PnZjphQ0Gb7oVVVGjzrVOSaOiUcb4XH184zSSP3GzwXL/354I+PJWNR1A8SaX+
HkAvuDafiPCunnegx/Vke6hVmkh4b00/Xzr1SevJvfhbxuNT1ofNs/4bzR3YwFOG
W6CV+faK9TT3Gxsw//PNHQ74ukbOo1kk1dLQwMLW+pkE7Nn26lT/5sqNFk+abk6l
erCD2P4mi+rt4mTQ+ebyPEYzCF4M7TrjMORwQO2Ke4iRpFVwW/GonPNnJIFWWm6f
O0yz5eYYXsLy3Z12Z/oQGXFflUZBd2Wce/kytUAL/fy4s4FI9N8rdlAatusFYEr9
OjgnGP+LFuklwWmwpEgiNEQJWNVB1BYryynfegM/p8LsJq2c9PmRHg69n8P5onnR
W0uiIAK0UhQxQzgZM+mnLpWx1dI2XNUbuAkA+G2jpztqMOvsZSKFDZGO39gcaBhZ
+yeQolMLygXhHZaacKss73A9eDl6J7v0+20fYlR+HbsyBOPaS81LNnR0TLq29h24
4BFykLKli0FDh1/Le0/rZBrcq7Tehg7yxPdRf4NwGs9P4zfhBVyyQnXnndANx5bv
jvrY2uoW2fHlN9hat/zvPDDZuXq2CYJCE3mL0qU/VvZBesWDX/K/V/vNek3RBh7f
jvzXV1u7ltqsnsDJjtfPauPVYqBWq2YPIAv++ZP53/ZXP43Vy/M17+gl8L/9M61h
C/rfmd7XwpHKXSoGepDbNGPD3shgbhKXm86ezkYXkfCbtdpAOZIKDS1RwiO2223m
7yUCM7i4gvStMFSLncr/DnXqShbT7j5ml9K9ougwfcz5qQeYD3Mf/ceepzH6BBie
`protect END_PROTECTED
