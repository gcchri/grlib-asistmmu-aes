`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UZhfq6zfrF9DDwm++wOGcb20ncmEbCYwOFMjiCFATGxJ+0Z7AZ1YVDEJsinQoaC1
ji58UrZvARDLbp37GAuAhVCeOB9pc5WdyzyriBByD/HM0wfT95zBv+PWfuDM4E0/
IFxCh+oVDvlGN5psjX+aTf70Be7QwkcinLqzltIsizVS7W/D9lKSc/w4AyAMbf16
zKUimpyULfLeCrI3bp31kmlv121MVRALi0KOWM6GUHgKDX0I3ZxjXS98LXs3CU1q
`protect END_PROTECTED
