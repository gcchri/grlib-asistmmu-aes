`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eLJx5Iqka3WTpQ2lyMKh7RhfiF8nMHRCz3gj/GTr5OaxEFCMkiRFek0WUrl7U0/I
wMa3/xdBK06T/Q19v1oHIUUT9JVSlTm30h/A1B9n2bBo6eo/u+dS70LBZgIDYzOj
n4Ju3390Gl58RcIh5nSiLl5ug9nmeBDxT1CqVeCCdEdWWnW0yFeSchKKcdq3aaz8
prKWQBWu0CGWFUpsoD2Rhxgm/DxUdx6XZAW7bMMFaHBnmnNwoOUdcIvgN24J7Yze
+z6uwQwnD98eV8NPwezUgncfCDkXfzpJmV53pLP1oKx8a22axKkYlQy/wr4Sg/DU
PTlK0BIURgUNYai5KXRV0DKs8+6Kesrb1hw552nLxXeDf6JESfoQ5pvEcwYyJGrL
tM8DVDlydGUNCoDGuuJT//zWVGJOYm94hZsaulOXP0ryFwZBH1yISBWuc9zH2gq2
XohxWY23FGL26CVpjE5m2en0yfNXjlYXk54nuqAeJUhonU95xci8pHM+p62BWR1q
j/Syow98ExAcFS9T+qD26r7/5XcQsiWQD0EhsWgcn6WV7xF1tTnztDDatYqgY6Is
JJtVXewRxTKc7A0K2s4ss6smKUzuAeK6ECpkZJ83M8so0VRh4N0N/8YUHppiKPxA
aJJDugC19kzdT134Y2itRX298Dt9/9D655tBQqh0rwFzG/TMlOgF6W+8eWrau2SV
b9edpHmLrs6P59LakiY41MzH69Q8dbcjsGWHd2kd8AHubi4wCojDcHr5rQdifH1n
AU9ZS0IKyc4n9yMfypLIL1wx0Z2AjUILK2Zn+ky0gS8unE/Vtp5A2331ck0ebC7x
zj5zk1rZyizrP8W0TRkKCgTAoaWz2D54mQycD4OOtDkJYGAVmFe1soH9dLJdG7kc
QsV3ULNCxSADIKsmdCrKB81koSrB8BE9frlcBK+vachm55SA3k3EfSL7iCCoxJRz
37zI4ZE+XXdDOB0R7khtB1ApUraHo4G/bR0RVz/TYRfPb6YtwRGXMWPtYOgjlknN
9g/5WRXkNbxkoJ/j9oL4Jhd63ah3styGTEZ37hZyfmC+Y7GU+tIobAZLsRgxrviU
+dK03UjLmoO31znLWKW7gmLqYsgWFzP7qY1ea5QfMTmRsBEobjwtgXPaTtmpbVzZ
5QiorWI5OWJ4B3YE2lmyb13VLap4IpzSAXXLofhHQIvJ8WhgZT7LaXFyro1VR9GR
Nm9MlpQjJmbyPo9gnBBEZqeLO+u4S/4PWcs/o0nPwcmSwoS289AGMOwlPG4FHd4f
mAl7lnxlvxWLXu5N0gG0HPC9s/0ZwQKi3Imx0wJ00rTwoElETSCbinlbBO4oeRnO
RksDf5hBgN14zAnSDeVladj11qxVmLnHWaijm5JV0hOitIQYgKtb7lcGTnrK0MVN
Ibr7SZpqCzHTTBC4QCtR+0zjYeGPBd5QUWaCYqhNpd2op5m/pSbV5ZW0OvMS6Cf9
qttnwTnmdY+A0+2Uxe7mb6cUyiru11+8PsR7X2L3flKDKYvZckD84/UhTo6FsiGX
G447WlD2ApdBKKS1ZtUdpGC8rLniee1jXz3O05tGxUJ/ZPU5PI8k7If9SZUWCQN4
KYuxQgmaXwUl1XQadJH501MlKl8lfPPZW+lrIIHYuJp6Mr5hRQ64FaMqYG9+s3eD
oPpcVEqN0qDT1SfHMG/KSZR8wwRGYRnwj7BW32PrTQM0+q5r4T96UZFHA6ioUG5K
3MgCCnkUzPTDwVK4hvfclg3ciDpX+fO1aNMvipkPfEfvVUP6STnJcqwE+i59T0eK
clGeqOKpKzUiFUpztGRCpZ91KowPZiMnwNWW+m6gG+edoBGb2+lPG4jsB6KPMkAW
3J7ivmlGcqBRlZyc0DHD6R3Y86C/r6Z8JRsOFBslIOvlC0oQpxoMnjvY4Xu3idx/
fwxwCuhh3kpMw1bR3HZFiltlHR6VovbH9tERuro5p+gi/TrbzWyf7ABb1fYgNfyM
caYwy4RSaaEWYk8Mo+kYMKqYrr0Nj7LKp3+JQJPoEgr4/mEWoKVKB89x2bGIn5/G
ec7RYUs/FSukPEjSTEJ9RUloALQDehNWAZGmgJThgmxDs0/QEvpXnqfWT+T8s6QG
JhPJUAQr2i4V9FAF9eqawl8qSQ71ysfo1CLpENWdRSXU+KPEs1P09N7bDF46CsgC
71J2dWrPQwT9mSX5DEPH9+OrslPm++rIJkpox1evfecPUh3nmjoj/8UduO1wF9X+
6/GxM3kA0A3qQSR87i4hjQUveNsBjT3AzEqjpaxLSS57Lo+9Vb/Gvynecy2McX8G
GjzFWIv0k/EUz3MwIwokMhputWpGX8dZXDX+86Lhr/V1cbk0wVOS78w4HMG8KDZT
HU6ThF0dE59eKbJpowQKJjxOqGuvLZyWiaH2oFW3BMRTn5rKtxBHO4mW3+F7ZZFE
ckOhwsDrEtXqdnr6gc87gBNsMvelrTQGYz4tBpAudey2se1gio1jZj9wVC+rWfTF
7ToAmyQY2WNVi13jQpl/b+gYBeIBcsYiYUqNShIXfpTHwTcfsSdJu1ppnuZHTOVX
YudGJfHAU0GPqVvloJVGh/W8SHoxE2gFrEe2wHfqBciHhZx9SUvMMxhaC81z1Msd
GMvHMlfOmbaMVLER98V4C1VdES9OOVClbabtOmRw4ijBVkpy5cZ4JpgZb5jf67Vs
DqWPb+tOezQw4zOkZpWmUOvIJG8jUj27mP2pvLdTA0D5eEG5MMXsLnKccIqFd0cr
aQhU+abQK8NWE7+UbvRrKSo69J+sw4K4mpsy0627gSUWdMhzQqkmTeJUlW8ZXfCV
YzFUMAda/wAfrAqVQKkG1RFJ/wYacZ91dtMIbovOnnNq8kMasEpyx57g6MDaxSt5
tdZExLGP/p4eAnzr7yhJoKvdQKok2O4YnZuMgxIrN7kO+TrnXasN396oECZtEHLw
XoK85bLiZ0/SGmdSnjZQogJI52IWtLs8Q8QisdAyzNAGOctcJS/EMAUAetCVR7zl
oDrW4q30JOiLI6bAQQCH66hmabp7ixNDLoDPCjtqYXCey1XR5HyVSHLnTpLvhuHs
tSrdQ8c41EdMZGpSo5ojzb7UXGuEpN6Jss+irQ9uV+YaRRiiqzr1lFSPYN9YV7gd
MucDV/kR3kuNJZUakpC0bMfJXe52ujGl+PcHRhggfnnpkVlKm/Yh4usCH39hXHOP
hUtJLvHOy9EoBGXmvyv6Y4ii8vLPw86MTeR6HeqNNoYskpxfk4dHqGLmmgM+FBPC
/RQjG2NkQ5TL+RYJ93KNio02Agl9lYqqVsfMvGeQbFKBWciBae3ZMhAY7Qc16iSg
kjKqcUQ2ZHF80aBgUjK9pO5xuTU2fwFxHxo4PipiPOzN1R3z+sVI1wNLt4RHwxtS
952YMGagQioXb7ADdec1d3vw28tKF3U4pJdX6OvxiW0C1MvQVtYbsmputuGhIqFR
61dKBSv5eArQkF7zaMBj9M9aKw3XF/MxtBHmOHWJG3y4E6cW/qMqadNYN/xvndCj
gR+QhystHvUw6QHNPU1gjQkxclzLSXjsXmSUR6Wj49JUwJlOWdxGoWFIILa/+clb
/rXzGDelco9Ms1aN3iU7N7F6OtowPJu16lWb6lsEh2a5dp48HGV5code+KCFlcSb
rjWDf3FnkB7BvbS5XFG6sfCSqgtFlGjrxREO4C1i96S9kNFbF2y8hkCkgoDXr70a
B6KGhk4vX25lW54Fudre7hX+75cpEoaOnzM6EqprW53vfC4krm1iOmQwnGXyebDg
RLel3XA8muRsVKHYEfFC4T7eGNnXVMXKZs+ovpVTBfRV0xNJtDyiODOeLM472E5g
sadvFLDqx+nX78dFLiOOjD17WZgFl82JvQn3273m7fL0Cv4TkAAilPk+HtEFhoaT
loCubSiOZ3izYwUbsv8KyPqE4ZJyVYtU4dzGKK8j8wvKJqL2ubM7S6UIPk1yJPJW
fjKKwcDb40/2no9/c6erp6NytGjglmqCZkRgCdZeyLPqqtBAKuxXf2ZZRTIGoCtZ
6n5wbz8qdJDwEyaRwgqfR6xdXk5Ak+pUtJD9PQ78q/IvtHWjNNPYMH3Sr67pFzOT
/RNFJgOjFOK/IDmV7XpsAQ60utu0MdWUk/LcEWU/gUTLyd6TVdb1HvvgkL/jKWZc
bBtJFepNpXCnY+BAkbKLc66smy4be1C273QllKFP3Bx3TPzNMSr6wewariEHrjnS
pFYbk9zrvt7ay+I2XD9JbmL1Pn0vfTBz3R5+IQ3ROyajoHmL7FcHcgDyUYnDlj/E
mEFId/ypiQ+MMw1oybd9hGZJNIGqEq4/s9FZJMiRPGx9fFErm0dXqN7EQ6s3tmRn
tXaB5/9a0bMQZE3mMWQOVqLMVv25LKepdfY3vEuGCEV8TbvX/UN3cy5MECLOlcAR
zfB1hJ+4RFqb08VIa/gcORKQ143/GiFiXzfTvRMRHo+EBiCYInvqG38Gekn8mcam
dtAnSZIgPsfmge87tU93RdCl+3F22ZWSsBR4ObQ8HuambpQzkvEz/lZOqbnJkc6E
SF7tFXrdpW5A7ORfcnpdRxvx3IYeQzAOrzk0UdIkAozvE8N2b9UJRRbqDGTZrR7g
X8o8/zdgDnzkgEOH9/Qruzs5PSR/l9nCKzz/cH3oP6mhUwEMF2fVG5h/jL2gH8Ln
ZmyNSZ4/lsXI54BPv9RtZ/vRVVHzSJqKTEm5XOlaBi6s9PI8XxcYkM5X2xGzX+ZI
rXlHRZ99ZZ2r5npiZzNnFNvSEzkOq51e1BR+aOBLFTuZEGyrAi1lYR9uLeUGTUWL
S2StvSbdlmdIYh2ZFiaRXwLMgO/TUMg/3Tw8SHfFOp0ctj/ahpoQAx477lNrovuc
R2wIbLNetYA9Cwm26zIbU5fFCVdqv0NXUoklG+zRph+BUFI2TqGHY2BSqWmSJmXa
sC2fGAzdjB9diV/Y9xjC85NtxEqJyXCjMTbFr07prRCAO8iBsmWzPr3TMha8bo3H
yiomM2jZFrNYOUxHsI6oi+iLYmy7w5lWubP0rrmGvA01qgQP5YF7AhTnrA1bDBvN
rat/pf2dV6KVfvrSj7gRLSYEw8j1Q66e89r4biR0otUlT88nITtb1KPlzdCcrGrX
gj/mDiblZXW5oEAeb5DvugZXjmMDxeSCENIEnJPo3QhOzPMKa1qAq1KQDMSXtah2
pHB2UMiA8rvMTv7uIvQJmaFUlnwMEoX/+ttUU/SKM7iB2v5JvhF0KmX3gaqnKcqU
nf+umaCGpxatt5kYQ72ypID5ZVDcEsfn3M25DuaQtizH4BIE+q/UvguGC0eBGiZD
80//E3inxxUzO5gEISMG79HYVqywIZoZ4USiy3g3x3/3jFQc8O8fm79SVc3PNuJX
RZuMyztW8jmPEcPWXsSoCQS9TtA5NDsXrESZSukkYNhrZSRblu7+tJP+ADtbm+ZU
SS4OOit4NMh1N/7G7qN/MhMRtxaMCNTsMnJ4q+Sqza89XW9Gy7YjXss+2xU5RyGc
ao6OU582uwCPJSqv+7B1MVh20zwIzZtNIGViJQJoEerhfxah+k6tSCumtQJzwI+F
VcAyo2fKBv8F8m6G56fEMQZHv5r94JwGMbH4KLUo7b2nopNAyidHVYHQlczsSL0b
ga10p1rB+MOI+VNWJ3/mxi0IR9/mfYP179nphsgjqIEadgC8R6QVa2NvqKYtuJrN
IQJIg6ywN09fUwb1RLtmsRWSgvUXDxBdb6nC22OjMzgxqcPERfSjLWl/kG3AoE8V
McKPih1/tGMvw5DrgzagPfWTKtz3ODSs8hHt+jKEvdtgvmvk8xRVrZwwSLqGXp/Y
HMWsIeV+n+uWRwlisS7/6/THhLcWwFRdQqy6IpcuSHFqLhbgIz6vV8GEp+0HUC2R
YlXh0gswBNhGJsswcKdq+eFxlqjKvG676h7TGZa3NzgLkd+DBu0a4Gil2adLzLIU
pvxohbyLgdjzUy5/FYdrW+wJRorpzmVS2s93HrJLGIbrBgFC2o71wGY7Jsn4lHJe
C/tnJSKB4MrzO6C4AZnEld6edUUxjs5/yift8Ao50ZUOHqhIoEzfKS02IZgwaZsj
KnTJaTtMAvODa72CA9pBxo4xAz+dOyPliAovsQ1fHcDXK1jnsmuB8Hd8U58qTNtj
Ed0/WmNStGsXLzF0ysW9cP8aa40da6ANL14TOVEs2QXEYo/7SgNh+Ve6eA7HTCxv
2hoWdnLlu9m3L22e46Q1UHrPcm+knygR7MWCCdcnYQIUcLpCJOUy47wvivx/0PWC
DGNUNSMAagmthRZuDjUAG7fuVLPObRJZcoZ8jZTdE3Xm75mlB+sWBDZcUAeMN6+y
1tPKLx2diDQFJ2D2y8eUhpLVUcagY/YiOnHXOAchdIafgPXQ6ciXtAUATFGFelCz
YUCXHExpXtXKrRn8gYftvLKFDPZA/+Axw1ijGxLgpXDr0ZIpIwLBamwW4vac0rc7
N6phnOQuunHbBivYfrAAWriqLYXLtWKxKrfapf5/rps8N0qs1itqBPkT/MEgVQRg
QCerM8QPA0pum4Kz7C/5X2x3/DfgPsjuFVCwnX2wT6sFKU5y6KmAHQ0JKO6FZhMG
anXjvoVOryW8Uh5mwyzfNaNruMiEvwUOm6Re3K80L6cLkwISX3a2qBX5gNsaeYdo
gwpFSUgQOKcrDmyq8nkYE18lhRhqStmOI0To5c5olvMr8rAmQiqaKJvdqd9EZe4h
bYCQSzV3lLzsD2CEJftmbUBK8JDsf/qKD3saXuncQT3ZN5WJaYQNpWiY7zQfWTgl
cfO9wSik1THbO5cC1o32vpZwUjeORqbPyrHG5MtL+dzH17UIlP+WeYyxvc81LGtF
CrwFD/mLnlinoxy1kio7qxD0LoUCo9bOH/EKoM04snrGQSbgndackRVEXEgmapPL
dM1CHYIjvDyIeM1/cm5AwfwTizy1pZQVYdIRUkXorBySd9yLxLbkAogTVmGLrr6u
RlEe+50tCrf9gdV8QXCaujOOA4dQ9W5B3Ma/HBEhY8s5ULhGD0OFi5SEaU6xJTmj
Ei/nH7yWW6d5hAIyvBEghzTUjZ8Cm756guHgwpEIjreOU/WK5wb2bvVjCloW3IbM
goEv96ksMECbRdTjLWiB2Y0GZSFFMfeWXbl69MMZwsYzzo5TMopgYpdZshGOK/fY
UHfSoQ+7XW1UDK8JmiMaQI/HMTbR9NKaz3MhrD/c/jH6GNyBn9+a2KY3OjEOn5OW
3iziCaRM/u+IoXveC2Hr8UvJFEbnu96ChoN33fh5OvpWTDDBk74cbObONlclqjCZ
CK5VEUzrooSmOStSEJ0TYldXHBOoYRT7k2RDqj9F7IPz7wQ3Fkc3Azg/LweObJOW
cDzwd+FSwHIbZNn4rjEvsImRqxUvLZUzuHHPtPvaJzvvxlWBO1LmY/5aSIj8fynL
pu24tvy4R+e9OPzozdwBSOigJKsoDPeewBZDOAAImOo2dYEoX4otL855qG4AsDfU
7h1x9YLm/dED9XDd6JdjRJxsDwBKQ8CUum+E2skbI8fnyWQp9cmEHypNcfTqQvRZ
+9fhF6nYqeVYWsfJvNeDqKNKkgbspmB6MCYJWmN7FxOy1IY+9dJpz++go3NokNm5
TD4EKAOW4cOQTt6KQGDwwF0XkPzsTVfZDRgdEzzvzyD/KuwjsdlrDG/dyFJL3tOg
n+WKS5uvW47qGyej2vXpGeWdVhxmDlbBZypSQPHaPScEp/MqYHCNG5DbBLU+GGEm
dx+DikcZamUfPodzzkMDkN0kQxAVkTQBu/dJxgQ+KuspKS7BbeCi8cV9ZfH8hFTm
XcsNW8k5cQqRMrfW0h7X6frsxi1SrJOEJWydglCOJp3xYbKbGWPeQ1jyboDtEH8W
LuS5L0zdXeGLasnl8KU3OdT77GE6cOU8ld8057viWNDAqIEgXujY2qiVS+bBbs8n
p/s0vOtqUiDUOXxkZbsTAY7txYJ3lVEzvY+Y+W2tDPMOerU71LhhNbCSSafxfR3u
81UYIHLuBcw/XyPLKDPTmG0I5FLrWxQ2DjtQQqxY2PJY8aLpkuAEtrursSNMOMdB
VMmaLPUsaaxspynKyN8Ezs9mb1QP0Ra9Rlfqr33wosoQDMrEK6vUhpYMWSeJeXVz
QvTyL2dZ1j9hXkbm44rRgrffm0ZgaC+a7XydoO8Fj3YLqH6Oxtif+TF0XW86Puk8
VSRmgPYf2L2UQGPab9XX/ydV1qSI5fNSyCyaHI7zWUpCM5LCkiwLGfVErlpj1IrS
dNZhGkj0NF2EQ1ben1b3zaJ/1bB/dMQeLoTpG55KmdkdZ+0Fsx/Twje/YGK6h0Zk
YjRM0w/YLue7gYBVKLvezirB7KX3dTC1Pij6P6hHslo1+WYREeidogG66dunUGl7
M5dPyvkJ9C+zhhooKmF4+Byrx5v+Wbnunkx3ymG+QRwK5wRGwfpfFd3DYxGT2E5v
s03ozwhYrU/U0sZcRJt6tJQDUu1D2c5UY0wk7JIUr1V0XklgQLYEWNCeOsYcf436
kvFm2engIXnMSUqBBTwOKwGBkJbv2BentZZKD8iPQkc266gZTV7bEP/04JiWWdds
0leBbv21eLd+2r/735Ga1hxqXgRdLWzyPgc1IBawQEELDHbt8jJPOBvmBhmEP8j+
VoNW13dh1HQJK3ftNbwap+rVa8VSNoc4QpF7JgIJs7So+aa0H4mE/kMBjAYhAgRY
GBQuf+JqcxGHn1QAa1ZrTU00lMgz5OFo43XMgVFn56aikYbCxyHr1yKmdbUxeXE3
PBeA7eQDysiHllKIzsiGvPkdzZvnWQJwZtK7mz4HbilvYjrBu6h0nnX1x2ycwn0T
y57Mq0dl9IZAL5LNUMzbqmVMFF+ioGGnlUOPw4MVBgVnrj8Y/AxxvVAJI+MzwT23
R8Lz0pT/thAuALeu9IhNE+eduhMMTAzlCJOGCw6f1elff62fJKw2b7QG0eooZ+w/
uEW+ln5FCzdGWcVPrlYzVUViY015z5FJVjnWTYLHjRxByOUuholK1FBKAJKp0YpZ
XakMxYga477rOoAC66eXwu8HQqrXXH8VgZPmvQb8FNASGrWWd7dWi2IsQI6MVpEj
nREW7eklXlSO2cB436tPtrJP5DKO1iOKs83LFba1UzmWr0ihl0ReDJEm65hvi7Wy
RPcN1xGCu/YteGRx4A3j4LVXs8XypC5+QijENt6LEiNXQTAma/gs2Y+OdHaDEYiV
YVkb6Kv6hNKXx9clyONZ7typCbW3mGN1a+++vTXrLtHZisvRLShlSNA15g8rvBVG
5/vT6VRrdtpfbeTOvK0jK/Y6BzRZ9Glufyc7ZOVS49gUoO/3HjJnDexD/DidGqXE
4HdPrf78vjUXjDg2O/6WvSw+Fk5Uf7v8s63QnXGfJypQE2TS3g51kUS8AVQ3gYfI
C4ECu4dl2yKvO9LnnK8jEYANXf1P/Kwhm75zku4N5lhfezIWoMWAA4qNHmFAx8Yb
3tubH4vyiqYjSml1DdpW5cfy/k26XH0I4qw+830t4EBfH/2ikdWFbgpxC5Z+8W2w
mH+75ixylxVk3ugiZi8RJRIQiF4jrmz5CWm0yRok4/0K5L7smSGenojKcfTULui0
hdNclxI7Xt+8vUgK6KR1vMNc0/x3KvU8YI5GalBIwmdME4vtfJXymUpya0uSebUC
fDYGE+Uad7feSXV5q73lv3mtjlReRWKkffR/0iExJfFfk0FMcZntV0dYc7T+aTJW
c778ExL0lGRrb3+x046dxyAGC8b7A6Nnq1T3upWCOrfZcf6+jwF7MEJq2vrGhdwX
QLMMl+C/bLtzXRT1EqvOfSIJI4QCjotmU5PV8ZtGDPIEh90sP+nAqDn8zZRlJdM7
CpwdSP+S5/+yAwiaSWdOxZQ47u8MhJ7Iwu5FXdc6eAIFHLS9pv08biuVL3ry4BC4
wJ3Jqd/zlLUiUaO2O3sHeN7RVIWePR92JrBqc23mvRxSLcWgWYc0XjdnNMmssw4h
iGWjukFg6UxkFzVFUEqN3TapcMtSTnETa4d8J0guxcfnqreHs4XzXCCKnMl+HAgr
JbkHHN55A3FfMybvlw0heJLPB4E25yqQ5Pbwgztr4fXCTY1GIuxNJczHISnSj1jf
XxdFCIY5pzdS2tRbvUD/BtQ3LIgz3pNFmPZxk/moAbwLBpBZhVE2k67VwrmR7gYj
VGfvdCUTgx3+4aHjtbySAnWHfv6V44F8QzQAQr+nV5A69zKEN8dVKFSjgBTXcM6p
Vzhd4Y5gpwUZeaRalUl16/eCnVGVbede7vZhpneTwkAQByA5rZq/hWkq6whCA7Zp
mQALPmziQNIXrWkGpTbLE894HokKBVsnIxHXSHH/1ec4Rki67bX94D94/NHaeeyu
aMWORJdRW2gdKGTBhVvgcjlCoGNBBk2OzLdtq7TouvQvLA1mhf8m0O8rb6dS2rZP
rfi1Uo1fBXr5JYoe7eYk8hEYGLpIWvsz46QKoOQWp2LO6JN4wqhoBpSkt1nEijAg
pUBwzHwbd98udk3mkLKpsU5sS/hpVtw1yNBdrWqjtQ/FUafdyEJ7ImiyOZl4YtYV
m3o3U01VCzFpzMwZs08BTFwALGVmlIw6L5846QaFFT4qA8+H+59X/0ijzuMQDzjs
/faA8tkk+d9Ld9aiyKU2MPPev/E/u0XISFwR+bHYFsJa7tMmJpu7abg52jumuSXJ
/WAY6WhEM24VhzTC1BYOEerMW8y33cMJvdAPJ0rZoUFuYXQPV/qplkZolgmPufjr
jz4PtzZI13ZdlY8ponL6SB5B4qi66SQmy4yqFb5hfNK06nwlSQLBxUH0o9JQrhPA
B0YgsIf+BfX5C7s9fK2it7tBS6fzVN8vBQr7HYJD6cfRqztU0EVOf2ADysZkEtRo
9G+RYzJeUYVHoY9jUeeFTVgfJeMFrf68teAfmZwOu9x63oHd1jwIGrUmN0rpdJs0
vPFksJMmgO2QMKy8Cx9qcB8hj+4z2jJkXX+leCd9RTuQDofPSxPW4FiyBavRuKA/
qhXGLNiF3aCiGoqRC0yMhBo2mpx5VO6D5e588eDJ+pEiCnXgRSB+g2RZ5Jo/HD/z
qd3dDxwBYp9qZ/mtBtXXiDXbGIsnMQZsw4AtV8y5XF0wT1ICDJMKtByMpG/9yV0w
GxBL808zrPSACvoEecsuY8EsEB50o7B5Qb1j089sU91sXDurXawr+0qdWxJPjOaE
D4qU6T8LcCrJtdj+KU6hZiBJNI05uRTTLVtK1yibo1MeCdWX+2TTBSXgqUWoP+ob
+zuwdlJcSIzLQ613qgLi0q7TFxtzja0q1prEfa0MNTRhtU+Sy51is4n/M2pUOqRE
BHASUlz2GqPdsLpCbQImVLxNiY33yxynfcujFW2n1Etq6INf33SU9y0+/1xvdYc+
z04ZbAZpv3ItaJQD1wrKelZBxLLf8j6uLIUofIO/PlOB8PKBgTCd2kpLprIx5xPI
uL8o/VDlAU5MjcU+fkv+F6uDt3Ghs6K81mCX9++WFjrOytaJ0IzD/1PzZWNrhX/1
TySQivx2JQQIz6kmXS1xWL2tyg71u+pnNtBegmMpXG2aLy61RtMnsaUyOfo9sa99
8zcL7IVsWakQz6E7dw+HQtNgfuBsyk+kXzY1qOaqbzJOirvNhzMMy7nXYAhGz8r7
Hp/pFOp2oRdLxfibg74U0plfZj+ABEpy6mIzdN/3YuF7xFyg6ZPvzMl+gwVHPmRc
1eOEeRIv7gBmbGOlCMGZemLDawSeYqqgkTmgzXYrljDDY6JoGbh6g5XCuNdctRWW
4vJmAQA8WF+JMBtahRD+kZepY+THkwrDdzh7l9MyA4JHc3wOFahHpX7tkSkP5W6n
aVLkrCrUQTiFKhclhnPQKzXKeUb9F7IVGg+NQejRit2gxMTGPo1A7yhH9TqOsh1v
glsJXeCd7iTmzg+UI39CVAljuUHoDj+QPpUlpB1vs/AZNbWZJO+NB7wp1zJA3EAH
/6NsZtpvK92n0C/8/pjytk4Sc0wV8U/xT1jBF60y8hUbHgBOTFmem6jD80vkc8Hn
uHA91VPUcgVszd5+0n0jmqdTz4gQ3lHJQNXnq1GOzasLbwArHguR7c5fN0FW3PJM
sPYXQ2gKYNxRYRxDkGRRiB8ybl4xtG9P3hfxtDb4rJF/Jak6jJLlVhgVRiyAA+z7
vuqMwVDNJBjEPzKogR7YTx0h06BpNI9OPXjGvQDnw3a9SOMATiv0sl34sWth4BSz
SA9PwFYx8/1HE5J3lBhH2WSCXUGPbj8t55yCXubX/oHEqNLuy3Sn50g7S9qVva4j
mX0tUG8FKo5koqjvi30LBvlFpGWCIcR6vJ76rgbqcJyTOOE26hlEXB8JkKQ05DHY
NeP6ApOoLoQTZabVgeMi6BRmJ/ilI3ucD4QvcJK25scdQq0n9+763ghi9zZGlUYe
z/fgmILXpAMuPQRa+8L+hxN6rwAJb8fqbZsrUfNLctQF59mUyruMxxNbEwNMuApB
dHmITRGanN/RWh3HYwz1gNtM/OicAjpW4X30GYwikcul6I54zTJfVJg1bTsvjxNK
FCiex7Fyd+k+edn/H6qLPoBoXZYda+5y3FEHd7yY+FcqQBm4wq7l7erlIjpPUzBS
yNFJ8FDKX+bfqAGI8OPlqvJs2eZDC1D3yTyQGFCjDOp8IoDC7TugmIIc2BxT/lnO
lOCL0L/fDyzWc0aB5yKtaI/idZ2tERahcvA/ukFpsiel0NoT0K7m0B3FKipPWLzI
LsvDNDNMZEO9Zw8Pu9DXTw99P/hPIeRcuuaKjqhKNrzQztPSnAj8s4A/v9CeK0Tq
tF0Dw+KTWxuwYd7MRwaI9Br3j0RWzS9J0kxPbNg+LwIYoY2eRMuk+DXaBww17/TK
DvYhMJT3tG7VtKcBpwCm/6rbC5Hmkg+KAAqlLRZ0wQl4c5pNeAaGPK90C/IryMhA
prqmmC5aEXL8rB69jqABzPiPZoLomDjw3FpGv55JhUW1/Mkon1gfUckeqfz/gTHQ
lmudQ7yh+kZ70f0oKR1c+x/K27/GpTCTUuD/x4D1KFKZ2bNIlx/kDYJDDoRXiQWO
9L6/Hx28E4VCYY9veBRELM2dQfMU5dLyoDT4yvmMoNiISvgtH/GAYLCUdr9XfnDj
KuVYmGQEPw01CxShV4kL+C2L3ckRMAK0BMTT6FE4cNWlz7E/DxtspS2DSi70Wl9t
xNn0BPWnvId8RP2N0sDETYpqPemViLyUEMePc37s5HL2qKqClxZqzSY4M34sky3f
xPfYy04gxgP8m1Y+DMaWiKmcnkHFQfXkQdEKaTVMGV/B/qz6qVM0rAlhNWitB2pb
I95SzXViRBno9K2OVzkxOe9xpvH4c7fvE4p4bH5gTGm8UryirivDqnLzciGwmKL/
1Ox5Il+1x29ZePDx0ZDY8huVYucguYd7PLdLMnWo4fDxYeIG7t8uulEGw+qpSp1K
xMEiqKUyqPKBKZy3jlX3BX2E3BpGWMpcBX6Ixf0JHdO0Bvzo5DL4BxvHVshszynU
Y1Ptby+GvMvKzRtvOabPCrwjmHc7H/3UYRDl8EdAUvCgFeZslM7WQY4XBM+fnY/t
hjElHh7tfzPePfZHRqm21XXbk0Y1XYI24RYEs8vmh2/h20KuTifHjpKrvOkXWxu/
shkkyPxHKXJJUo0RqEabrIORU5f4nxQEPjCpk3lnemBAkFM+7o8CD7Ery1t/Di/o
ib1Owm9nCHY6GrKLwS4hsaj7F3jBA7K1yBjrwtNNz1OBXFx8bJ1WibZWvxtPIoij
3gRZPAvhe9A0MSIkFMCvjx1a9FZRKhWedRF10VJmK1s6tcXylCESDKIQi468Ch9a
NbPL73KLyHDzU6FvkmUl31vvTfJlwv6Zuk5adNgs6cuLQF1EXQRufJZxTw158rho
yoQnKIhTCR8RVTtxSuSi+GQ15VcHsYKZyCXb6/E99aUtTA2Yx9oyl6sjxTYfRMAZ
HLUdwJSM3L6Wy5hww4MSF8zzvlgMVk6nSkKjWTFVzdVyMI//F/lZTRITndy8V7bV
MDyw9kq4yXeuMF/SmNEf1l+9T3n0YiZ8brpqYsPmwZ3mjLhaHhX47UXLc4grb00L
9jVSilRX00iHMWDnXdh928eDd09IteI+Re6MnBZwKA9p0lGo77TE2MP8YufYb4bi
KsHjvRLhkIKagzA6vodrE1ao+3v9p6b4N530oEvfFFweKm7zaK7buNi0pL7tutiH
WdIPZ1uO02Q6UJoi1qsGcHJhKCgnH5Q5FMVmRVCiXIzAIdhaMk9g6o2lNuTYoPuh
RPTfLfMzqH2q8c2k6HBwu/wQNZb/lrkxE8+0fCy9xMpJzxaRtCoUs2kRvSp7KlpH
6Us+bnbksUnQkNINlNtQFtYfCId+03zXjYC2UkLdlf437/Sb8fXkfrlVhN1J6Xeq
BtA2QzYVSxGoxDrWDgZTICzNsQoOBqaAqakFhF7hpB2E8kD1qcX5BaVczrxox3Gy
7WGtM+tX4o6o2aQdeS3gsZKlhx7MnJPIwr/IzrLEwvLeR9oeZJZbFK+n6jBzm8t2
wEzzE5cAQj/reYs+Cp3VB/PS4g1aMzg6YYFxuBYj1SqnM0yLDY9410z5tJ2euOzY
tVbXv+FTyjk0Nq0xKSxQ2Qhdn5DPA3IL7tRU7xvK2GvCgpijSSGNtQu5oqWqWQMw
pHsrXrpkiwKNnygSmfRcta9VbiqnoYV5+mR05QLAgFxbmtBdV+QiBwatvxCgAYIQ
pk1NfLpQfZyGkV2nz285/PVfIlhlrQyKCaEu0V8omNtkrbpI7igBgXzqoZ8uVY7u
kEM9pjUMSe3KALmnlGp9l642g17/N/eAU0eGl0bqHW6nRNkagEmL8AlTibt5fqm/
3q6vZCBxnkM/wt70kTZS8FOox4FN2qcT50DA6b8FRGxjKJy/Ua3fokoYMgi6vfOI
JKFs0F1kdA8EhO2lVkvDFz1nlYq0ObPcy81mmuaPODa+gv/5xPEzaqgwn2tepivj
8xO+NaX0qk2oZhG7nciJhdmhIKTUSdpDGRkJypPENBFzKjWqE0NSIqBnYibrZhhU
YhTrNrdL0839kT21HT8vMdo8Xtb1ryICTdV/t427o1A5VZZY3gQkUdvI3wdL+PJ8
o86WYbOrLpDVXdFj27XtRXUliABjG+v4CJ+tnEyJ/UjWOs6xUgkeQjMDdU8/0Fwp
dgfAk6bW5C1PFGvjCYv1F4AsuupqGEDBtRR7F9wQgnU0C9BYAA0IRhZ/EdCj5DCf
S1B+4Car0zlKjCFNjLDsbiJ0dpRNHmjSI38JH97o1SwcS0pKJE4hUV3iTMxCxKMW
FlR8tBkkZ/i6JpoEZ5IabYzDP5bAFEUeB2zNFloyLhQuJwdSRG311TsmMyPOzB6A
V0bvDrO7/RCFW84fqC8UvwU4QDgsGc+MEX4Ao8/PrrPz0EXDQRSLsAmXzsLxg0yF
LrjWVU4XN2u+rO80+381CxDIcr9AyCtJF1yXctWqoDKafcax2fHGpzh+W9oGTGx0
X0mf5Z5XSRI6fX4qkr94+5OMsP7zeVski4QQ+GTgqlWdCYDIdkPdCXns80ZgUy4s
vT05x1K8OnnZ5CCHNSRpfacVS6+UE0cWmeYzgNI6fhEk22VQ8yiKcmRRHrO5lJ9q
HdxUtJGm2z6H0DTU13rrvJGerJ3mr4NMK4B/mwLqzl/8e0qzuXu9L+yMl6xfvs9L
GxmylEwtt1+H8Ra9CymAXXjYZfiaR5z5CoQy5kWZZdhsqk7j2gjRdtzVetkwqgzY
zIN88bvnuZVJJGE3Q4iwWbNbtNyxYDev3bpEc/EPadQKCgNnqqXUpsvN9xgDe3+3
6xYBf5FKzfABkteAVyin0pg12guDry7tBt+HXp89xpTUMNJ5AQ2QQ6H5ZLVJRhH+
+gA2hYzOsBU5OBaCdzuVET1zl5r3y/PsVOTJZSotvvbba9QF046/PddwySjZ7+h8
ebC2bW98gML+brOmnFwlont3HFoF9IRceMnPBoT4FQwobfkeEb3oM4imAlHuzYaB
XtLpwcbFpFCXNEZvizA/T3j7FysTCZ5Oy6zHcnN8ZPHlkIH5e7lbk0fG4zCgsPuL
l9kFJeyNwIcsEbCzFQn3xNgiVA2N1MTvAnQlkVp928yA1AyzaPLlvxyjwPNKofCZ
2nmuSsUEHpnyQMMP41ZGabqRe6d4NFvNb0PMQs4qTWGdD0nVMZIQuSHxq1MbyLSe
y3WPFSveVsOUhRdmiPdjJ8KYs5htlnS0vKbW1dUy1B/DxlzdFCZdMi03/QlHRsLT
dyQoemWr+Wq2qLMur1hzbP65V3EjPqsX+PAF1+KrDRYGPYsC0jlflrG7yWxDMtiy
bGrXDl4/QE+TxexdVeUOf09zX/ekFQa046AhhocKOvTkji6GUte3yKavjAj0f4L+
6Fa8/D5h/YI0697OimoVsNsklS2nTrmqRBeoRCkDKfacyIEIHK8YOzr4swdiwqDA
cV0jT569oEfShqdbREdz/1PGX87H6He0T5jIId78woA2flOHL9nbAtsoscu/qNVR
14EGxqSj/sk9i83JtUpdBoQu+I8cpQHqG7Vej0qfSj3C+QhLb5BHuVHMo5geT4Yw
QfXKlJiH8kCfJzGTouOq5P+tyXGzxSOz9AJ3Tgu/Cneo/Te7wEle8iWkrROs8Mh8
9u3rPlCvIDdWElPhI1Vz3FefpTfaE8uNzhNulEgy88Gl+i1UH5r9I024Dx1uCLCb
Gg9l5wrbQu1PIdCDUY6hO5g0j17oRZ1YHcHFCCv7JdL91UHMCg6iXw4PWqxLcK3H
ga1HIoQoAF4hhcQtKHMHyG0w9S5e9+W53cUkl3DzwesZHPUJPYq62LCPQZXO/IGi
ucsENgA8nJHWw1/Q1PFceZy6cQtGdmjStKOmdCxqDS7LZZ6PHfPYhl929KBcTYxL
9wv+23NBogELk0LD5vAIc9YKCEzHGeExBLT9CB1opV58gWiCWY6T1jc4JCwCUf8I
4qK46Of0geR9s/SfS6bRkDnys+xSjXxAphJvXRvdIYkPtdm4yuZ8HR8uvuP0GnhW
LXpkNZweYFlROHHt6sQ1bSqZr0w01A6Fl3HRtW11A+LYqUs/PEdjTgRfJHus36xq
8zYJGx6lddrnSweYYScAfQoZqRY/s7GtR64TihUYJ1vyA7amdnv+ExV2E+m6frGD
hiPl7tto6ccYGPFQgvEjYpP2wYqfp5ADDJVAx/Og0Va3ZJg6QQ2MvSZyAEVGCDRC
Omgp0B+gUrQFVr65XIBXPcwh9OxwLTP/h3uO7r9jtTje2E0cJGylD+fGPl6qRC6n
ZJzXcaJU1I9zQOenL6KQVeubHBYEnJb8HNLNBGROG44zvS6clCqYECBfXgOAE9vL
fvn6QvKu1fw31cJtG0wRK7J+1JVkX1x2gbnvmt+B0MZMrPzeH+EjqrbM+Su1kmit
MHZeU7aYipZB8d7dr1zNOVFexJYw6lF6qghOBobWco4/laCiBV48WxetQmxygKuc
aiJGv79rS7vfPIv8Bk6Egsr60mB9+w+DpgdhGjXUqHGazIClada81b4E9pomA01w
S6o96lunpElANINOm2FcS94JpLU5oTZmrOcR4D3tUjGFsRszXQkZI/d2XcvoYZS4
19loHHf9zj3az09Qs9sdFlLhc4gZcr7QiYIeAPn0mGo8O1wFWz6LqiSqy/O3kXMY
/ElSHPyMsomxS756ul8S03u+7wcPKJzCMvT8JA5RFaDt8FJEJKXgIwBuKajXq5X2
p1epe1++3dCbtIc2nDVlxhtxPGWRJQPLiOLALWMVX3MovmMjwiaVBLJvzurSuhVL
vLhK5X47nPa/8++zCPeTye3FKUbsNe4zxxRq3liw9tSMf6yPfmlJdVehmlwb1FFF
/JauNP6+KH71V1/cUZY7yBe/y/m1Uvpf4HjssxW4b3UvftWxBC41S8MjSzYqffS4
ovzt2u4JCyTWAwsx9Le/aBi6JO/cjFlXqyVQTKNa7rekrW49G0Q1xv8sz1ZjS6AW
rrvcvo1dHTqa75yzFPWGw2dEjYtTdYpxXpX2O74x+9dMTU0xKeqJiZpzXw76MgNl
2/veeK1PjSZzsF1Qb/8in+ivWwxS0evILv5FuZvi2fgqUO0GQ9BGuKBu2twNVU3u
RRN3B9n5PMAi6hZJhAHSWGogWTi77oFexcG4SBzYBASN3OWEhQEpeHJ3CRctYqEw
50OFwa1C93pBGFifmWWe8GfrgnWQUya3SCN4H73/fPC+tWBu2hjN7FkXPSSxw8CT
bFWgM5r4UHV1E1Wd8ZgLt8eYMLcanCfflkAE5Uh0+m02iswj2mvd3WNK6/Q5hrKA
fPnhBDxAH+B7ldwRr0cp//uKzy61nRfJZMjCfyi0fhZHuo9/SQOxj+bX4JafJNmT
QWfOzXbsq1PzJUshyz+0xaZr/SxrSEx5Bphn2mflCT28JZKN2BGJH6CpMrAKjJpz
vQsbFeHqdbxV3ueDyza+uz8GdgCbU8DF3oXNftf/0yzxhGYk8+7jLP9k4XH0W6K3
zvpTK/kUI8jiyabcJ0vEgksmkNr24jMmx1YpuHdyl9l++yelpO+LJP14I3xsrJq6
j77bkuDaSE9+UvdQXpE1c+HKaMCddBIpEO5vD8wdBP9/fT+BHfOD/Z6Egmab4Z8N
/KFZJIdawfxz5PTguDr4fs1Fv4ihTCuyT2qhzxocS9r9/HswfgRwU23xSZK0x+L7
dxs274tIkZOHo5g9KsFa8jQDhtObBYcQlHp676xGjgsiOYgMfiorjTY7BdSif4m8
g5hfjwkMy0gXAuXoLs/Vc2i9dQA7P8zzsQOvtCytKEUkyIK3lPI85CLhACZyebOA
XtnWsbQdMl4dUDBsAL7J6imd52PJZcm6XQ/j98xURb8tU8lgrI7s02PI81SfInCO
XI8IK2X+jE3V7Li+dJ1EkySPlDVwq0IMnNbDFGTi1Bno9rSCyg9Rp8ew2KHLUqAQ
RpU8CkOQfnTv2oLs7sI7NSbr57ECULcfCsuQVcfPDTg48NRXI42m0uar62ylGonM
Go8H+BuM+euWwOGymDzNhxLBc/gnwFmTjfVg4Tucgh44+zB80crKeuSOWVfkmY8y
VVFZjUh+5E/7ZKKoSraLf2sfwLflxbxWvbSRBr0ELYBRdwNjXqp7vow36KaeNWo4
pouqxthegRowR3e2qOQvy7pB6dbnq7J85wa/aSv8SMkkMb4Qx5DwXdosL1hiSmIG
JAPD3Hw/1YdunhJA9c7cnQolzcPDZxMtlNxWBlnr615kWbchqnLNIN5Rz1669dWb
YuirleYo80EYUQF7ULA5l9HaBYv4JD3LMYQfXFNix0dZJvFi9/en1Tz0YTaowry/
167PcrUY1SXb4rvdA661SVT71KWiQPeuW5WOho6CEXPUpqfQSIPjmbLoORS0ruJ6
FeYW0HVXw6cNNj5F7rh/Fsvs5+0xLyyGgn+hBXG8uH9PbzyiiD1Drg41ize75MU6
hcgixFVbOZKmgfyZ0lAtxqapXPSpm24DacEGBBf2MAGqYLuXggaQ3Xsnv/Z74fL8
Q4eQEWznJyohtY9QojGuXmPc5VNBAvzyQdeVqYBHyLzXKXjNYltkGRSVzESQ1h9T
Lhbvtd9gkx1rOQXno3tqH5Mmz4Cty6/wgqw2Zmuhhy3066mThiKOmS1AWUVw0DQT
7hD+ygkzd0Rvm4caQuVTDwL7Ms479/iEoQYBj/wPrlJ/t3XXQDHNk+l7fTN+mUyH
VPp+UvfixJrJp+ctaMLx7RK6NefiUF4GReLK30GaAgbXvZbdOHNEs+gVJYOKLiVb
S54MRI6KOC7TerdsJE0jVlDKUW2t/jLHFXprPvDgERggIZ4JZYFY+6caUYDhaPUv
/+Y9dFFv/lHoaKKQPTfssVMliTWFgIrAZt7IAKb63ODvXjm0Igjqiikmb8ixgFKN
gTaoSQdu6u/Ed3KIrVa6AUBQzk8ef4ykw9sYBve18mOwv4hQe5Isdyf//uFyJ++f
6JEWf87vzMTExJYcmgxaJ+ovQ0+ymffCKw18gLtZhdMlD6aj7JgpEp7YQoMYMJs/
zywLuOJbPZPcJJg8dPgQbrFJ6vPMc5d/sAoj75pODwn9ivr94EilmD4WYhyh89mg
pzQXnpazy46ujpfq7P95D+EUAbzjmbzwDCywGGo3GO9+G4yhwwF2g7RJNt5LGkQ2
/jLfeifiUux/wxDu+VNzS+H7n5wyTnBvgaSgAAeBGCSa36R++Bkwf1rH7CE9Drrq
l0ZQ2AoAyPt5b0xK1dJEOPwP2gCFdeVQW6z8L+SBQOz8mKEg1i3ndgFF8aHsgv3P
M5oJwgwHSzQdzxxbXlYf+eCyQCpagZxvtV3TLYP8oPsGq3AY0n4r/Dah+z/ORBGF
s8o3CuP/E98gM7AbHgZfQIv08XMTAeCYboeOt+ULuEgq68J+RZU2wzfUb5SvXB90
pHfh9DhxHb/qTy3q9g7TNZi5rv9cCysrzKtD+rFYWA6G08ZI7X0VZnMyTugFNX9l
HLuCozeD0U3u+JpHBtoDkEiaiaM8ajKvpBwYOtKGXG8ccI3WTqBEc3HP5UYQ1EpS
xysWSX20Bq6rP1Bjw5/Cvzdj1deOAnF5heZiYcFLNIHtMU2kYz0zT6wLdLiG7vEt
21ichXAcLQg5MD9TwM6j8dCkBdOil/8dQqGnSmnb59fz0FH8ePky6xT3D2rIqUn9
JaF1deSbMJ4r6CTRZq3toR6qnNWkFCIg/1J2GTCcrGMeFhYhDQBPKCsfDjabFhkd
XlQJ3E9HJ+qv5VAybTqsSzwq2U2CVHIVwWtadD0ELJag9ETyq0d6myTliAyJJfv1
FyJKTi1suWy6ZXRyCKgoWxXk/8hbSuZDCjBeFLCssaDTGoMDlJFfAUG8qgx2GfOm
TIERtDOr86kY7JG48m3++DO01+taWVY85mn2j1+dTwrgCaTFNGkWx5V3n0gw0coD
h30VENjKgzGaJ4nSnoNDYRtP6TkiIk/VeEBLiDD5qLkC/Wjh608QZRUmkwIXM6wj
AV0uwaP7sJXQ4MbfD4BLc3nrxRyQLL61P6eLX9LrxSNLIdf4ArkClYNPHoBs91WT
0ZfQcs4rFdn/Isx+IatTyRHZ9qHbvtqj5OB6Gpru37BdBA/2OzrZbUS/hdaywQG6
C9TmOcv3JvGqybYzdvj9NbMj30FgSV9oJlyrIsBTDLq9wEYF7yfxyXHMCWnW/V6J
8eDohf6mf6jEzQB7YEsQn8bulOUrDmNgoapxlfvmHy29D5qIsb+Tq4/518Mqh/Dt
5oxBcsdepfv7YdYP3jSuAtwbLVtKMVdgOj+G2LksHKoCxx1gVuix6z18q/UmMSdc
OWeSLVQHZ5dFb+Kcp07XMLI9HUQAinzNDscBnIwdIfvyDKozaPRcPPek0dv4JnK3
IQPJPphDzihtAEcGKQd8VPzngHnaw0AS76IuYJ+LHRnAMrxbjN/CT5I4MXP68aVc
+oKRv+5EjUfJhKr+5Q0E83Y8tKIL5zM6HQuwx3LoGt2XrnTo2S4Wp0rc5vzsGzhK
QIZOazOYEJ5ZKy0d6AvQ+RZ6bC4S1a1N8S+yG9SnR0mE6saPaRyusQM7tIAlHatj
dTAbqdJ+9FUmz2QTr+e3J4gIDFde6e8ADC5DQCP4EtFw1hRPb/rN2YvhZa+78iAA
ZFLbsMiB47gysbsPRtWEuhKce3Bbinhn3n0aoMPYtcOdKQd6zbff2GCgo93qV4SG
92pdo5+X2puiU5WCqcVoq/TAqSfbET5Rr+zobbfKyiIGR5Rv/eAzFY+jkDOajNDy
ueNsy7pJspYJXc1vSW1MPuFVEax4JJ3RaiAaJICDaVr/qCw65igcTLVqkVygvxia
Y5PYqZNoPgwovUfS4rxXN2Ka4xwrOCvE487GIX3i7L1I4kQzToE7fqjpannqjNvZ
7tj9dnTpMAxCmc0Z1T9anZtQXyv7hdQ5iKTRxnkDo7R+7b6brwiXs2ykvygpcObV
9z9e8WfUZkLiU7pyYCChgiHngEQCm0M8/5GkC+NQ6hS6QEE+AHpmrTBqqjq0Ugy+
fSWW/KSPypX5TpBWhLSYtuQwxpVeVMFQ3N0Vcog05Ky3F6iQgwtXfHHvasLMPCGG
JcAiV9SReIPbynqqW6Ri53g369S5RLMYOlQP26UG70baI08aO2t/1f/L2CNzkkJR
+8nWGFUZlX8qpZ2ufcLIzToYkfHPhH8xDEZiBYTHQKPr49zwKgug/qwdfaQLUcW1
1zvg4AAPYmNXq/FjVtcGu3RCPFr46IsGDiuDIH/ON8HFjdmimfY6XMERHw+8SJOB
gmv2afgVYWdjD6A4grmrOUMXs7y3KtQfU/7j634rqQfd+dqz2niCuAmq/9Zm3Rox
cN3zBkrTunfn+7UptaR/0Lc0oCjgjiQu/5uHPAle/RZPULb7SzxxLtJzVX42mz+M
HcsO5aeLGAwcsVBHQ+MNr4BXiihORRw0pkYUDDD7OdbdWtP+x25Lhfajr/DOWC3n
F2wNY6QqvQW64xE/tjobsp5u8zncsWDvFiHUljRjLvUZH9UY0bmaKmSiXJjr8S9c
baEpstCIk4aa8v292ZDIvpguveDj2KbWOANQAO4V7s5wCVrD+f2/fZMLoemNFLQZ
gAeH7rguzCwY+Q3LWofSF13uf/kof4RAlSShnO5aNpdAe/IAeYoK8ajZ/TQ2ADFK
hTJ0smR8uBh4KeSEt40Gd24ScMn22tGyf5YimQyD/6cwNLnXaz4C3eZrnH2HCkDb
2kUFn/tZYOmLp7ah6n1mpo4t/YnztOz9ssDqCUgVqIboRx+iO7qCXnxS7JwStk4W
Qb1SCTZFalLqnENcY1gtxg+AnTQ1jTXCqs0Ta/5qCyIqIPhE+4PQp342d597m0hl
EMC8dvx1H59NiCFqS+miTpM2SS9y6QHUf6pHpqOqGI3Ka13El1pLvzNYanbosQ/U
xsVwGG5U9ighl8XOZbMELGVevS/B9lTg0pDWWAWiAdydSnKVqzGFJW9i2qALCZll
q1hQtCXwRVvF5Ykz+HQlR3UbhB3anNH5DHzQXBMVjRHmZbOFv81wmMhkQjV536jI
wvXfwmIge85lIBgrDmCF/4T2mGrAhALXHSsjyjOjbvZpmia5tuqVg+kN457nXbbM
nbOZAQWAzvAg0bYKrYuo44ShQhvxFolZrGm8xU7sPnz+aKRDGsnQyQgxqt5gQB6r
bnAfFd7FolkjxQkJjT6oGJnPQh7iBy1JTKNVge3UiJms1zQMBQeiOASpj4yG5yU+
0UbpAn3GVb/SSQJE9D3bTfa8W9OaFmPLCkziJYloC3nTiLYRtjsXZCCdmMNHJkBy
W26dUpqhvZq3EwOpGKUIxdhAJur+di8mxOUMZdjteRBcmJ/Qe48ebVOLv3qb9Pmd
RhdXZd8DZ2nbvCozlqPwHUihtPzv+OaReM3yYyRdHuNgjhkG9zG1SVsZTxxVbXCH
16g+86Nt3hwYzuu2Yc5aHRmyW6tBfd0w+5325lTNIJvaG6nfOHkw/sM29MYBqcJL
GGg1NjXqpzFT2eUcYKZlJcvcVSVHNfPkPcIBGY+7LY6GdWJp30ZJcgHmQ/mZcweJ
PcUPeQOXUGG0htUjnNVW9nzpQD/XiZ0VV/5LPH3p6dFG7ZYaIQDy0itP7+svco0D
ruCb2n7HVgBM5fXSVl3JmnxJqUxeuSoFY7hvBvjfcCpPlUm58MDorqydjaVMf8xv
Y0TlhMbkjiwmMMelROXA5CcPmZaNXzS2UzAuXmRPGDUFnpt0I8HRP5iAAORf2Tf1
N4J55hoT2Q5s2a/NRwcbAnnRXcPZg65AWBPFGSdTEBBuGLMBMRI6JKVl1M8AoYVF
T75dvZ6IuLH+1mCpOBds5MoeMzY+K1YciQw4XKzRfKuUuAxzAAP8XW2BkF9QAOkZ
vMhJsAovO70ZaG7CvSiD3eBjTPOU3e4FFGXknm2rH2PEuBNszHH7B6A1kOmp+yee
Hba9D8V9C9rR1FPa5NXbYrKDkwfoXSpV0S3fa4In89Vw0BnZwbGBaweFwPvbChq8
fC9doNd6Ko7hYRbF0ZEwffM7DRzOyAvnJuUEUR/YWekIuwue7gVARZObZ9ebNC2h
2RQX/H+JzdkIzyHbhiIMXCACeQ4GAB2R7berASbqfwborsyhKTd1AtIqxju5KW1L
57Flf2fGuCeC1hqxxkpNyEnI0tgiRgbAAqK+m+DtO6dpuY+y/ZvnS0/JXBr8ZTW0
ZeXTYViXOWTLjBaGGfzj5TgyNfbxDBLe3kUKwxRcoulxYXdydmfU//cbfg8Gi4cB
k3Abh96vHPX/2uWnnAX0M4i1HCZ12j2sz3gD6t8LcfpW0Feie9dZ0FvNAYAlCVz0
/VBEW1rqQ80mPsOrgzB5lAUr4B9nRMEAgNuxMvWRV9Bq5hjwRYee83ReKxbS6TzR
LdfYb/f/Ug7fX/6eNuqq1BlIy/HXJYTd1V7aixzdgQAYU4B4kga2YP33fJ19nKBx
uE3OVyx7lpkCPUZjjGBU4TGRENZ3mpEma56hH8uUacNQtdSuNxKyiCNNbKP8aOCd
VQpfjJpTOXweudEtg6dwIwGM80TtWrRs2J0vtKVtiI6MOc9oGpAhnV3VO+gS1tk2
GMw9XpgQt2LBU0NbAUobauNVwV/m57njs52EeTO27XKaV90iUByic6OojsqWSFE4
t/D54Nf6vsU7U1o+aryhvQwDJo0LIzSGN7zLDGYy4KmiWNUi1w/xDZrPG8MS0m6v
MJOg9l/skL8vbEQIHNZ1/zHj0zFc6AmVAKeG444qG576D3AqGsWNJYk3ml44irw1
B0sEVZR1fZ2bLzX04LoTKsq3d2yThVeNI6p+v2wRMjsoFk3T2CbjNMia6LMIyi2B
BWG95750UzQe9tnijbKx5ldOYFia97KMDeJb6MaIIPq7iMpFCX5HN47OxrDv+e4G
ADPmfzHSuzVNk2udmldvN8hGmzuQYXhNt/7fS0/pmIx3CJdmwX8W6/v3yn23r+uh
gpcj3IrHIFKIDq4WpdKRX7i/jX6sSzC5MmubJxtX6OxLXYYN0uR5/iaENNocUAeW
FWA+rC09x1l0W4HfX+9aimFW2IfSxi0q/lPH9azJYgqNYE08UOZffxlh9H9KliNk
s4STlv0GlI4W6V4Sf0Z5S8aHZNk+t7ZNwDuvo12nF7qYOD1nHMxyRmPibOnsaeAY
bBITQbuuB9GUVMt/kBGut1TWMirOeMKefcSODzelpIdV7hca7zJz1qcH9ySvPFIq
yBkftHmE9w79eP0N/rZNwK/8qnZYEXzlGBOe15GEnLpq2S1abDfNkf8wdi1k8Mrm
dWkVA8eLtdg8eyLAcwbiWyTNu8IrrjyNp4gtVCF11hYoXcGdF8Ux2S9bMBI1sn3C
Qp4eOtgbMimOTYjo++aWhmCjSCN4PPhoRVM/LXvtEdiiow5VZn6Vr6tUVImPHHGj
gsKPIPhtYYVfOg1TRx+TH7VIDWDXq/sKubst4GPseEGloXOfGjMs4/jhN0bYLVt6
CfCfDRK9Tu+vOAJg0SCNyrY7PQTWaLgr1VsRjSqxGnasw7IDOo/gDU5dGXv4G5Ok
QXBed94UkdFS2uQZM27dhRNCPJQYbqZPYYJOCleHgtoDkASP/l9e8hrm5/uar8Cc
hjyvIvIj/ZcbzxF5NlIckqeF/w5THwaI1tOaSVFB+stAHayB4mc2Re0J+agfUQjK
CMqWGFKLXH9f0U5ghGtMWi8QUlylDUvnX1WeP+WA5dDlmGunMhYFoLmLXWzBmVuk
x4sQbIj2zzh9c9psyl5ZB//o4E4hfdEOd+DVxE0P+/XNLFZvXIcJ6O7a596gUF2i
2rM2N/0fvNXm+umZsjS/HnzUxpB5F5rc+e8F9/Bd/lcranXKO/Wfdt9wuxHkLfvR
tHunhRmbC/ZXJboFSy4ufQ5vzKdi5vlyqdGlWZFemrQe3ZYVnYDwF9pvWcV2uu8q
L1R2ZzmmAkxndBbpwBdMEDPCcwBc82oSgtK5pcB+Q5YmunEhckC7afwZcJtdmySO
DKWGuZynbe7fDPTOJIuNsqUpXGLuzTHKZTdjKj66fS4NRjxwjNzC3HbNynDkMrWt
8gOVY/dXlx8nK6PS+6H+fWehEJ49uSYU3+wfa5BTOBaGhe0vpJs7sS+3HsFND8br
fylUU+fetLZomOSJb8Q+mLJzb0M6CA1PcOdf2Y46ItEcVnzmFqgSa/v8v9o/L3uu
Y1+bLFDL5wop+nBKO2mlvX+KxOKU5jKZEC0WEGkgQzMEsgB9weUyGQGtJXTFvqui
eqK8POd+l9J+4lznL3y7BzTh1cAz+kQ3J9XK2ERdoeucbWcXK6nY+MmaHtqz1Dbr
A29dWnBuhOvK+7sngMsdWxgU6xDrUPh7yUE+6MidTfmp0KShTcvt/RELt6FyEKGp
ZsmeKJxm9+F2YKdBSA/UVkmhKKlgpykTk0dg7/M2DplAEH1HQIG6J8tCmjHCXo27
n+HsazivgYRXRdsMJtYDA9gM5m4BZqEfRR/0GeCpIOF/sKptGM5SpucCH76LSH4a
m9d13fnVkGhTc1nhAJYwih+geUo1HXwfGn+eItIPeqQTB/ZmDhVKc5yi2bU3fMMu
CGb7Fc6UqenjLQjtpAd/tJXPhmTA8p3aZ11XDpLLyO2+rMei5xzN4NnhHovcl0/h
NJ8hEFTUgKLhUpLVK8HcG4Kss27OSfmdYiAiNgUaVoMDOh8K83wwQq5oXmBvJ+ln
AVyn/cLgVlQCogRJoAo6rsy5kvcvOF6UzIE9sCaKCKG/XgjLKWuGmoMVSwMy2Z4L
jjGGIg4/5CATxoQ5OG0X8UpS+KQ3TiGwg0Vi3PkabLkilOS4b+takiGgyG0209wz
60j8nNBxQmGshC60k4IjoSABbRqO3VASxkO4Z7/I+apE8I5C10zoQBb0bvcrS/J8
rEMZThTgBAZOqWUQo61uTYrzVy1kU4Nbc8TtEeSxBSl0L2lH+tWHm6l+dSinffG5
2IAQna7AXKGIv4ZI7GtuZzw4hIhpPGbETyFUNzV4hDBRmulGcWgrj8ZIP+CkcREi
gbD74ms5ZI/Q6sNwvG2OD/W0ikGfhYabtt8KMqSKw7PHJCaljjISxtGNEW0ApOmK
iMtZkkaYbuVXWAUMbj0XnPB5VG7OsCD/FrlHCpLrXlgXPJ2OMn+YXvXUV8AXCCyh
sFOBJOZonmxb4/wO5Y+tWClrJSxoK98H24XGg8pqAhYi7ZkJW/todAR/I69N5LYL
dOAXuoo9jh0r5kR1bpVg7a/EU2Lc8yjHpXfnCS+TdkqE8O6teSV9awzvTEK7ZQ9u
i1GM9tMePqTkBOjXE3yG0WgERJC8Dld9RBmUmAgH+jdSFUqNzN+8cKwVloi4x1uu
Rh0t1gsEXZFQZLhaX4o/lMMMrvL6xaRdvoFB6iME73uXU0DXiG3ip+AT3DMHGjaI
9EfsDL5m0CDKxcuDcXBIRlQ+eWLpJsyWOz0Bw5Q/T4Z1Yd4lHsS9kNjXZ2EiEHnv
+ciRljbDtJ8w+y9g1YhDTotAbkF1KZXwPPjQts0ZgINcUFjyp6lpO2eGA9CDEcOj
0xfgsk+prsnp0BXKtCLcu6uJfth4Eh8T2Yob7klMgw2AymlE6wyTjrj3BvOdrGUk
twoXTnQrJEq1tFdWrZLb1g==
`protect END_PROTECTED
