`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0c8iuNtsGmn1Pu6dfvG1Qh3MonzuOHsq1j49fXE1Y6KBFEVM9meqEbOWX2qa7dkx
yLkRIfdudHiNFEseKv+30HrJg5a1VVEdLUMuVdHNQT/8+eLoXfd9vUXSsR8eHfzt
RWdH8aB+7PNccUvP585XbcoNHfNtZFNyZL1rSX7N499rLhY3POl//ELdp9EVt6ww
tNO8CPGfYvYdmcPfX5O2s3+nR1hMKchvaotKZIqohrlBg7/22KwK/PkA3z9TWCAA
Gl3nt6vw+97vVwFjcW56jV5qh58ubK9Qsdjyl5zBZOmq/Lf1o43qztyn0AtvVwhB
oe7PErsczb03YDD2YN91VA==
`protect END_PROTECTED
