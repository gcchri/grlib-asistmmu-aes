`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NPlr0BCwzzCJFZnBIjCIMfeTCA6WSXhdOEth9JfePZz2MG6uzjvcFIARF5dzyCXN
T+TECPZ9Kc/Hs2w92z7VQ9CxvrLPCc8b9Qd7+JOsC2oHLHWAF9RlYQ47HwBHf+br
WW7QvBNgVVhIAjZagRxy4uzStQ8+pjCqfT/9bf8A3p17LuN5SbBDYAQnPw6KPfL1
a42/OS+DhFLBaQbZPTUK4WXSrDB35f1fEQFwwWR1eSSN9mK1m+tQeDMPXSHoh4d2
ozvYntNAiUHSt135MbpliEkX4KdlEyVt2ur7PUTxOIsMw6TnVPflrdnGpnhUrEZt
BRHbob28anEl3xCJ6nEdN/9uXfw6fWK5nbNBgiIRD0ok42kcL8lfv7zPMwvIrof6
56Nuhd4qsuMEDbFZpNcPOeHzXjP9sz3ZSLkVNwLu5nTkNlnjZ0GKFEZD2tihIKPp
SvbAw53fqgl3ljKoluB6qG05athIx+MjnRJbkC5HHDP+4bhxUUTFGQLCAnmAPxr0
vhP6vlW60LyDl3jG4eIaKcvJdNGQPSg4rHLu+iWLCj2+jBipfTrACQ/iDJPvfy5Y
0Kvrg7S9Qc4rBzjYtu35F+t05HCck4g7wGmTOqxrRNgA1lHBsXLYj3piK5xpeFaU
S/sSWNwMim80asZEGImKbH2UvR2rRLoKw0AWZ45u2CiETgeWuvepLas5YCc4pmZh
e5kcFWTwXqs1HJtBqBsfeTvaP9VLlu87sDbPdK5bd+0gpEqbk9qVfDkH6qdwGoGK
hUD/PN+YM4KHAC6PHWD83Qi14o92D5BsgVCvsM+HJPJJuB/XxLdlxWt3i6Udts/x
l/U5J8fNZG0skqVMzrSpxw==
`protect END_PROTECTED
