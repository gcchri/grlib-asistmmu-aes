`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jxulPFzCkeQX4rf0Er3gylpMR7NCu5iycBAf255ANamSjxWbpbTXRVPxFJ+sPfkq
zk9WTQQt+kOuOVvRiT16WgwUZwC1H9R8X+LFqhF4t2TAwNYuJJVvhQPdGWbzpQ0s
4Z9wJ3Rlw5YVidcdVT1ZTTqejlwMQiyiiQI5znQNCsIsW0qQ0g/l1eIPVChqpg09
J+w4nMqrn7DcsvNmRtM+bMM68wwoTh0EbqoS+JXf/eOIfs/6F8c96wMKZOIHHOdk
LhzttcCYD/yXWjvYwoxT+SE/DUe+7U6e1oPZJFKyXEsx/qOgDKI/mL4GR95QpyN4
ZMBE/LLCTYIAAhDaE4hF2BW7gn9AJklB7hJ36WWwaLHPXza+7DjTiypGe9M70vKr
lvTz+eo6BX2dGkeMof1TwyzvP4R1Z8E8VF78PVu2wyXVOHT66g2TH628WOwdCrna
f69bXf97dXtA1GNUhVXh1oIxPLW44PsXhHKy/W08Tbmyns3lWT9iwxz0qcPbLxYo
`protect END_PROTECTED
