`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RflV+vhvhvq2/XTxYP4SE4/3S5GuauSIulzpGxq8oHLb9nnX5dDDoDeoWuEdGAnv
vxBIxuVzv+yzr15HIIqM748FHHcmYxvHG0GsJtzTXyyRI7vECeS6bI2hy/kWST16
pOnjOou/0bzaVjCieMt3eBJavxmCIpL7mI/9QrHrbELcNVFPFvjU0bQS2+rDBxH8
UrME+MBb6q6MPvPlbAm+i7p7k8SWtxHJpa4RtcATGB28JFqFrNZN4LsWTrRvThu4
s123QPbWPU3YCaivd0Fd6hfLvUiKRfNZ7PQI5bMnDYNqFoYqWXLHH8pztroZpNes
Uwk7jHN45xWL1yOEod3speJm7ec9fAw+8j++oMrXVxlnFSFRTsrI46G3AZIylbvx
r7Nbk6DdX6SxONbe/0EhxQ==
`protect END_PROTECTED
