`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LZfj8K5+TEJDeiGEko+/IZde04ylOeYcgl90a+fkaKkdyOVUm7VxnBVIaSSUk+P/
AAk3otxgI81DeFRbEGIlRPt2vAuDYD6U/l9fsfTJA+zXD5DoAYbmzL/0T1zjtQ9X
dn7t8R1xQcpoNerw6Mp+1zSp/7yssc3t5lX7TaYxtPF3/B4fBVqQhedVPDB+I+bE
VyjpbUHAODXjKXjqEJgjOa56JLU7n/Nij4mAKLHjcilhVCwaRgbadVk9SbTfhkqm
xiCACao22ijkJt9ECALRqu6E8DMEPGsXZm7yOd9OpNU09y+PXlKFMzi/v9phK7og
Z7owNYKcAXncyW/Ao4WbVBXMKCfrYjL8cYjT/PTBDuxrcxbmaLUZQ86Duy2SdJu8
hSahRxJz6p4G45WUfOxje2G+91vrBQfVUWTTBfLQnDp3cTdy8mo4qA3Oxao1EVII
1BQreHp0+2PMMV6e87YcGd3UuuTawlDJnqPsv5YyjV8=
`protect END_PROTECTED
