`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ukoooUBfPrR0FdB6VGKq0BbZAk38/4Iw9vuN9kXTGFK2zNyx8HEDFgx0pZ9Z6R6c
yHgmhmwm6NAlrMob17txl+PtQM2gAB7iY2okQUGKxN49JJpl/V/fvpcVXEs9ndBi
GnqUmJ+EZ/N+NGMwphisoarXHMsN9vVC//yyTZ+uX3GTGCtrIt8zsiUSWnY3Un9G
54QsoEI3CEtG+fItdJnuz89MN6K0av02uKxotnkLN6PebOUPqCZkMxO6DndPF9gq
`protect END_PROTECTED
