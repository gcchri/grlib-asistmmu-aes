`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WYwIbPIcvHOpzC3rM4/kO1wrUxJqLERoXUaxkOaK8Rt+lmDZQkpjLBrI3StJsxF8
m7B5RwFW4Y37W0Lj8C2o6wlrCN0Pu7Qn3saLWf0lEI5ZtaEBsSnyAeXGkMM2MhFW
a5xFhBQGBR+fZsqhyRl0qn7oiKsJ3WRppne5idOEcNTKGdjchZfoPKAWvr1z90no
au+Id1jtlmL+ILTMeCPdjiTT4Xo60GtTOa3slZuvzcWQveT1ZDZvFFomm2xw72Ym
KmTRa8yHfk0/rMJtBbRMpONZpZglSIbwm0ko9LH+LBS8ZXh/jm3gMHu9itbarE8/
hfaiO27DJybhRqmYdpDq3BPvnJkqBX3T5tkkDfSWGqybkQOIxmpanfhQt74JuOmW
z1BtAUyA6NSrcLBMQvLFoy8MUO3NxRbLIBXvaNt6KgQaBFZudiOYDrzQmblwU1AK
GOWnonVCCZJmZD9uVFCy3Ip+n+xC7P//km+8hxJfaoPB5FCRWtSa6i7UHQgAt9OO
aX1nA+m1R+eipD9stxtHuQDECkXEv9o3NoG0cGDry94DcPiTZucQwuyQzh6M5d13
607TwgI/UWTnJsWK2Ml9Jw==
`protect END_PROTECTED
