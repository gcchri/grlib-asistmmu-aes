`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GQSAZG8skQ78d6sfvLVZkgCTSkrCy6aflxOad4KDKCURwK39xn+lYhgnuYYnCaVS
oABAYFRP4Rr/YD2HtX1oaF/jJgY53fMjXSBm3GfUYTJDtMVUIZmrqP7ZF39rSj8G
ZkK0ygtHg7ii0BFyP40qgzJFWkCuIsayhFLR1GUYH8D0QHfSUU6Bsk9S0osDLUwg
u3HSWbtVDvej9+u59B+DLExnsqc8lt0yJzbDTCkMMdGfZ7+i3/Qz5ZGZrEJiNtKh
TjWPalyhk2iO2U5GbofI3VNorVEA5+T265M0Zd4ecv9uvANA495r0KWZuoFKrWY5
94CaEgNyaiUzTp0WAYSW/5xFEmRTAdNhljwIWoGLGwKyq+PDMjyBBj+1Ssij8Lln
hGDQg5AJyJ4N7QufU3v8KzA61Gc8uRTgLtkMwOcPfepWiH3HwYEdo0BdHcWvI6zp
w4lj+w+/EmZpqiKpxX8RtuBX8e7NGY1gU5n78EECG5kPjRMXTqNe0M6m9NdK9PzA
kdJkxRu1PY1nYCy9dtvmVICNw+xxT1QMNmbQUBryufCOM3J+gyfrQNkhdSOzyJEB
JDvgzdugNaxASIZGps+sPtA4odMG6Tv5kRVbnZCFrSADtjc03VD1s1pmJd6ItZRL
JZznnndqCDyf/ycfpiOkxNnbrANT40jGJ4HbgBN6W2QhEyky3FOOEvn1U3Ofypqv
9nHV53gLhVnLGE9nqSrzfnhNRh/7dE69HIopTVRgEW7h3Yo3wdmlj+dstNnkJ5d7
DCDFXhVntBpSY7k9d2O6EVtWdUJP1cdrypxouvSaaF78BxtVbOmPsPsmSWX4IK5D
jdMRpSawAMFg0KrExGAzWhGV/ukhpHaAoEBTfpYSiIN5udHd3zxvoahchiLratE6
ZaK8Ax97cpkvGW8XXGSbupmSkaGfDhxkZ8EuFzROPzRgEvbErPA4qspkwsWNowIa
yxq+YjpH4PFypiMVWF+su0E2L6ttOoDOlZBarZiUsoeaoZRhNtQuhuX5FgKr5bmJ
K+o9NOsENyjxEBNvnEhfFD+76JedhVLBW8iJgnjPBVL9dDDMv6+FXQNWbT2WovKX
G5Ds6j0C5q0LsC94VTLNyqfe3D3uC8QQD+P7gIjqnPwJYxaWoirjPcG4zLd8+6H4
1rQ0EexYiPhYEodEPwGCveWXzZ6kouDeF00lYE/Pw7sxxwy8iTL+fqA1fFYDk5XI
Jr3gsU+ov7TsnvAnS8GjawBnxV9l2v6Mgp2JDM0Ln292Qqi41gKCMEZZD+5ocN1/
Hx4eoc9+AeNLR1a+ZawOZcYJfh2qG+L86HxMLaLDNoiaHzdTm2a9w906VhyXHMtQ
qStRZjeLUrBwME8q9/TJUavXokvIAcS/MWVwzjKpn8TPWDKpGEdSMG0ZI+v/nBMZ
f+5iLNKOl3/90mB/BcZSUqlJYnSbCIDxIom0Gg2G9XeTG8ZN9AuAGfYVbp0HzENU
EdDrzHKYkSJqmJOpy5FoTK16JMYptpRwyJJg3srJL2QMpipzzo2vut5eudcMNy7R
f5r/kv4Nz129XUOIHGINeh4cFOrl38IXz6EDQQ2SBnoOO9ZZRWJdTmi0dPW1HjKb
PrpqM5WrIdvKarS4xQjM8U4VPsN+vbU+G7FBhDXLybPJnsANV/5c4VBLftoEuXsK
CbPhiusAwMNhJkbb0NWHlq/zgXAmP6bG4LjygPuTJnaCjIqFoESsBj51d9yUeAef
hQDeJ1VosWEhVkAFDeqDSQLbw1b/w0BD3L9Texrxem8+ZJJ5HZSFAsYMv7TFxggk
f1nY0EWXfzd1LBkCKVpPckt9lpCc1tQi1zpvoAnLurZiqMseD9JjMcOyB+5relei
xjgaocMy63JYG62iAbe29w9RSRLB3nY5P4aHBj5V4Qxw5aAlHiK+Lxije66D/2f5
GPDB+1waykrCtHR3WXi5aaNiBch1jqJ0f5xq5C1VHE9uB2UVFjyUwj+22nrpqyLZ
YjXrhSH9PLiq/wpC3TUpkBDXg8RXYQegw3QI+fkortawNrJaZSUbZ29bDW6mAvlu
t0W044P0yU8T8LkdG4unRH1/OyHQmuXra/hRiwbDoCIdF2vgv9yzosGm+qIez4e6
9yWvwOwlxWKhGDwdd2RTRnl4tNMvh+LzLnZ/31PXT3EbR2VWSn/8ewUFVxuXe3fm
ZTRp/j7l5x1oaYRKDYoz8HC0jW3hH0NRj6A/drFitjJqUi7lUqX9lJPTjY8/Ukil
ma08l6Yd3sAp4iiaLurro5gXWFNg8wb93ta72N8r6OKdE15R6L3xxD7swTj5b7fD
KySkeE0nOFbLE3tJeP0oMR55DUDGZGyajAaPNT4UJD7iOgvG8lwHrvAcnE6bOx74
vUlbwBYPuQzLR+yZYaVlhhmRnDTJlqXUuh03b9Cun0GpCja+iEmugHszwsCHSmhU
Ni7Vi+WMh1cKKDiSztcxoi5KtGI+iUSXoK0fpHe/XhMenR35/99XcZ4Am4McfBbp
O8l2j2lHNeXvkRcNFL+ubMH4h2cvIpDim+yKn603u4Vl/1JXzPP6GZVJ+wjP3rg+
UcQzSWnL1xmndLWZyvi7+J7Jta8B6t2VivHQD1gUxxs+kbTHWVewn1bCeyvgy9+I
Ibn9cTiTes8+nq+Hp36GQQegUtXlYsrO4A/jYQVIzCY0Hx6bduEDRlNczF/WlocK
Si8FgTLuEpbnVqtsz6Crkql6nbDvQESXxZukU56KGy/LCaqAYH4uHhZrkFtJnPXz
IZVgYITFUqHfegGMMW+38Lpqi55ZJXH+yv7I+CQDYyORy/mky3zirfu9kxrmBiUX
swlb4Q0nsUflRVRgEbinLKbMVcGY2Bzw5Fosxb7Q4hHlBAOVo+Wll2qQKiHbqNS5
22Op/wIIxVTPMn6hHS0y1UP8kkdO1jzjvjQCiljc5QK+vaflwcEyK0DJnNzu2LCF
kGBApcBRXWz2vZEhjLCVDYRcijRcmVzNldJJOKIpW5sd6KOMVtrggNqiWoKQWvIM
F1TaWIRfUbIjOc2Md8TaR6uIBfjDGn4SA9ngowyaDkY+NFNmxcfdmKdvrihnxwS5
09lhGpBQmn7efK//XY0OstEKvs8+g9ClxjsQXBGjGzYWtJysOYyu4gcJl8HhsV/3
pJ73RauViBk8vUrzu3JsaBO5TAJhGV4O7IQqDw9a5OkdrvVADgUi84P18zbm8zaM
hzYUoSd9jLdH2bK5x1mRKC0YWZEB8r1tiwneE7O1L56ga8V5JvQclDWxNl0qmFe/
APOcpZ+Fmv2MtoI6DxyY8qwTPdpG7t2ovFeEpVcZiMc8YbfwJXTwuuR4FOgb0+5Y
/Usotctb/ELcAMDny6wWkQ+LvRgGGb6it6vVEG/qpiDpD6FvLs2HRPOH04XoLZ4l
NxQoFMBlryLzOAuAW0pyYhMdvS8m/YubZYzs8bPcQgXYBAV7MeewF3IPQD1afZQw
8KuWLzN0qnU7MkDbXL8GiKySTJMtpV1k65k59VbZ4bpORbkRGdnV6Kn1uwkbPLbf
sbrXCIkDiOMP4GPQlzx5twSNVe2dSSxSGiYInJNa+kbbbK+Se73Zao3XJ5KhKfZs
28ZpJ9ARlrX+H07C97Hl5AgwCUv8yo8uqPpkFrlSTAgzFjw23G5IvlrD6mT4kq2/
T1DaSCz1UiAS3fVrH6qhSQw7JtckDb51WnowgjsYtb9EZiSQr0WtH/ngOcE8BIA9
LHt0G6J+xSYJz0nGT7UWM27AkBXHn+L/resKsbZbk/NKf8EG2sbZ5pBmU1yG0F/L
/aXqsekueONUK9B0UZy7CqjW+fIki88bw73gOYOjNUuf3odFeq2AxQebgjNq+E7E
HDJs4CIddXbWaTzvtxd/pi8NJcJBbB6ppN3iNrbpCoBC/eWeW45793GT0usI8h8q
afyVWPlrHoYn63XrhXDj3fhI1EnX6lhWy0GlDxuo6zSb76vEWDNOXEKPRuW561V2
LOk9+a2dMaSm0KZW+j+7arzruY8IMFQbtiA3AOcAfplTVIfPuGd3w1nJd+A3K4n/
Gh6TeJf/vuc+M89mDiXlp9FIP1po7CMak96LBYLEphCnS+4RE+X6Zr5p6IJfDrbX
AHV88HNI+QlzgsqrmEuU34Mno+oGl757Bwo4zj6Zr21rN7BBmQT3U/IoNGx0LT5T
9ExS8U6XVp61u81XJaCoTKHgykwxj4I/weiPqcRaxkpXW9N+FBP/gx19RA80Lzth
uD0C0DJidebBhP8tGFsnBU+JxFyYcEd8S8b47NXFznohpevwMPs56B9Qv/wy2ViK
GR150jjdPF4AQlaOGJQaacEerdMjuvZVFGa5H7F1LvYXLw/CdKRK/4vIfnDQL7SW
ctaOpucMXt73g3ouRdhbpTCpIoJNWMAzOHnqrvSTcSd60bveA+kYE/qg0EQFOcXH
2pfamAaeRyclf+y13Du2XOta2wXZrlcmmod1VO65Ew8nnd9WfqIFOF1exktzy19G
b1lQlqGDhLlKD4SX6655i/5566N/bK//FoY433CloBwvQKxiXkifRKHO7u9s8sZ2
bKPXuHYm1najowq8V4MXkqGZmDEOWwCtXAQFt3XiydDRLinJMi1Wm/ZEWcJGYBnx
D+/+lqRZQPLhplwkfQivD4wHnEE6p8V+y2pxvuFSwpCpAJcK681a8Q/BvG0y7rUF
SgEg4U29hEOPpwX/o5B4Qiu43Xrhr82Hp9O3mnPsBcOlloiIRRq6Hmib+jd3+f7O
jQns/tYfxylaA6vDzXAeqxyhw1wQOKY08CEFJVWYxIv/q6qX/E/a/6iCoOQJjJVs
XIKUybmTqXYMJ3fxdyYrbi5TASqW0UYtRRU712KhGMY465bv+vSwGYApHNYr3CJh
f6aQjV86hITZyHH4wSgxz+0gbSX+fM0QB5uR5E49LsW6t/0ZEVBt+rQHEenxEWl9
YmezWnZ9WALsoAKkMl+h5dq9tsCWWByKTSL+g8OsvC4roUPZtmorl9Ba84Pp4x4K
STAJNGfL3uw4NsfkiHGt3THIoql9lbKo7loEJ+SD+k0lFB8bo6UoUDuxEgCOEeM1
Vwc4XhDyqACnx6F5/PK33gcfP3tJ/ql9vxcZTflg2c5TINE41Gu3yHaojKdRX3Xy
lTh6F/d/mSPrzshmvn/qB23rNJREHgyR1G8JnmrpWTY3rp4L0f2cXMypLg1NLDVD
cms8kE0pq0PJlZy5T4Cxrd9EBGgOOJS2ckPqmakyL+RvfdZ5F3+WRpjZLsw2HUS3
wKULv6iC8y39edfGzCN/UN/yoNUWqdoOB+vmoXAHNgO7d9ZABl2TTFfhij6At0Na
Angz/O7ZNmD16sZUrbclwx0BpMUD99YHrFi0vKoXHIfdC9t0b3f36r8U+3/XVYnR
OIkcpVhbQwobrVsJbJ9fDIWMZT8nH0XTQbhLOjTBrwiqPSLbla1rkC3o3FxTmZrD
l6XcwzWuEt5YsBicV8nqvLrEZzN6W4HSa5mLRKshPMf9mWAIvQGXFyRvJOLaCCxo
nXdLiLgXFfaxnFVQ0wJkUFnMoCIki8Nisr+21xiG4i57op666BlFBGac5fyHNjG8
vW9hdjrohjG9C2rcLGXTsfG8/k4EpNwJkWG2KE+qtiNVSJ3BvIKobIeRyB42F7F7
3dHhR0fdt/LoRpf97nrVcwE94F4Htf7cOFJymIFYrH9DsnD1g9xz3mvjVuofMRwV
WnAXsaMRjI4grE4sucZJtwDDQViZfVWP/pogMVNagxpATLb7PgGYFFzxjMRAN4rG
1bMA1Ng6mOvj29boTOkO6cxokQTAP2OzqYxwgIC62liHexEjlzVplBYr7lK6XMrx
U4FbMN4U+qHCw8kveQmyNcX495sReZ5lLbs98L8obr5CjFCJR/w3SyoM74cnjDBZ
dtVs9+eYpt/HPyJjeU9GevuzDjTfHTAkq7YborlEReOdy4kCs6inDiKfCGm1wiQa
Vvf6HW0zbuxDaRBaep+AdtgQC/cFAWQG7sACwznE+sErCiz2/0ejkg2z7ljVG4wd
A/+t3nxp+ChKjP4olGS26YJ95u3Js3vw66WhXuwUgtIpY9i42mSOZXXLi9posOyT
POdPZMVWkjTsUJuHgP0nbUk8L59JwRPR901vJpDYc3xucKctHN2RyaVc/8RuF5FW
ybpTIFVFyXovRwintmQg1Irr5Wy4XIt28w5ZYG9CDYjm17TjgBOdvJpI0EtxCJ95
KER59yPa7GusehkF2WthXessU4B5pPPXI7+sz0OO7zS96ILE0ArsHTg0Y1kdbZdB
jRw3QiCGDiAisJE6w4IoohXaRp3RRgMr06lLZObyJRTCYMz8wxaSGOtg1gvC8rBJ
RriyTsqlBvaothh/48aKZWkMEWiEdWF7lsTopXYBbsAIRprfLxBBKMLuVQywHL3k
hI/r9A4WCSZ9QEGxhoikoCVGB0k15VUNegoyxWGWygUA4ebTqsph+uADsleVCMkL
ZDgbDmqC2f1U7lkLRxsfPFtxtXQhOvMG+LMwqPwdQwpej7mkNJjf1jXCCY8ePKgJ
hrFHeJ+wpP0WncmZ2nyv7YX+Mj8oGcatuyCc0kpGR+2OqntPXr91FDJATKJFdMPa
5OnGwNAi3K0lHXo/hEVUGHzaZ2xf2B/aF9ub05ZlLSmBh9UuhQsJuIRZFDSChIJ2
I0Mmvz1ojlQWcPJFaa4TpkySaGWnTBNUuC3i/hhcriKhvNS+DksMX1JQTuZVeKuH
jkRXpn9US7nOvsSuPwIvCRBKe4R/nWxInEfwX41S0ZBgFLg5JnNp2ukWHqQTgrhV
hYsioDvLj9Gg2ePNgrwHj48vPo8KfDQD6NdMDrz29f8ugZghnDkDyazxbTrq6ORy
I0EO6Xxdv2u7OwLiBPDBaZ2ryWcDw80D7S9TbUoA5m85fabK/Jet5uIwi7afGW9d
dJHvDp6bsESidTb3YlAd6m4syOGeErvOlUgTSzrFi0y79HY3Tx8a9LYgK1czn74d
SYDRFsGbyP95H4ogKnpxHhzdyfS5D4OkBhx4BDTcoIbpVnxYyVce4sEscLRkvnAj
KJgLJWqFSQi2peobALWwrdgyx0I2M7n1SBTEErmDONhTMQgKu89F1uLlXQ395aUJ
jyjNcHx40+CXyuGeouYbQSE0HE7pb7EKe1Izzan3GZ9gfsv0AvHxit5KIb9PwZqn
4fLN21XnPX4kcrnh8q78GFlJ++RQcHhCdHgqxp1oTndQtmR2XtIdbJBXE3jnBjoQ
26KINydNv+vlqWz6GNU66MO1AgFHpvYCc46Nu0oXs+YqtkysDIVRwMwu3xu12K90
5a67HPeuwWTeMgTSXuMUEpbRNVpDe+oRWU7HDTuX1bR+j1on8KVmXGZTo4jCXqjF
8yxNENyJnCZdsqZdeuigNWdy8xc2AbdRr5HvPntjYfeDMyAKTn2FEjw7JpNhSVbl
pxiKA7EWpbYVyRDn4iUKezVjexeBlps2HPPNRCJRbJ5GExnQ9qGsdka8plOlPHqe
TvzG45XxOVW02HPEy4WLDiG30eAnCk4mKObeXFds2GCUN1n/oGOXlLU1jbHwn1x5
98pVr8AqxvOvhPnGU88xk5QFKH5kL03hxQwwYi4zPC/AO1kK29fd6crwkPY5PkZn
1fgJkLF/ByW1ECd4bU48UrlLQLO2OtxLzFY8gN2e8aXuy0zMGEn8GZ0H28x0tgHR
2ZxTcp/7TaiThDZx2HbhV6W5LIcxLIfcMOy16X8KLltoFrFDMm33pQebRLNR8ohU
1kiazzmtAJrLv4Fq1ad6DO7mDP2ta+YE/AH+DBUnZ1kdg/P4gAhtOG9U4sr7ps6/
KE+P1bRThSshlctCwTaSP8Ebv2Dx/Apl31fm1lt14xA9jUsdVcIq9qxp9IrwmZ7R
WtIOqKP3ixW6wAohsTUvk9f3I3HMecV+tsDQfORdsIBpX99OF9dFmSeREHpUby8E
kKTKBeM9DbHX07QZFuC3HkKSbJKZ4Q89H9oZd97V9s/sW01uz8s7+E8UUVR8vhR4
iqiTTH0CWOeSipml8WFpzWuN0VNvRWtbNfYD/zX92PUlL/Hr8yLVRqNCbQgP5ynx
AO+b9Vzi1nCKLZzDq3PvwNb56GkxclC+ezuKcwjdcrg2VPgRVW5nn1s6moU9SczP
N7wA8bkiOmKuVyHo7a5tZJKz6cFNpkXGKAmQsmyGCRApzHTcGh8KsHyHw8dC/Uyr
UVg0cGbya8zJewa4YROhEnWamvA5e/jHtIwwmNg9qyVIgWAzKA86VAr5xTeR8pV/
aRV8EcMTlc4zicVMk4yjjMDJhhUIewznGyHB3GfCnao0WXuvDhsU9AHJXpvKzNq5
aAhGqA9irZrV4CN53uzYov072Ai6g+qn3X7He9t5MFhTn3KXRgwuPfxIYh75B86u
Z3O7V3hLBk+f5IaWp5pED6ft6qXgIA21WgmgJ633q4oddUoiCI4ZXBwX8+ODoIA+
DvL5+YU8xery1E4j3bDjr5uqW/BOT2TBNmurJXlmgco75KHoKwwm0o6LI1YsnwlT
lGVmNGpFIuXtC/g9OCF5p0A5SD1FxHesgnBaAtOmoBFwaPyozPTEqY5ENS1nQGxH
4G379SoQW1XM+NsEQ4mU+sy62ExokbNjP2J/IHfUA2jpCWUQLOo3REjovW0yZvEe
+Jboc+M8++hoQZK8JyKYJeB4VqTkRfPW6TF7DgkRxw9sQYAGitqkaI59QJ/WutSm
B3nqpFIwZNuZ1aYMxhxKoaSBTVG5Q0oSqWQAVJwbylfzA74OEFuD/LlPqmBa4BHn
ckkkaSaiDhfpJn580JbezCFhB9JyQwK3hQdbW9iqmr0ZUezFLv4ameTmwTuVyy0V
5WL3tEcbySlMR66z5w+5JFy/Fo1zaHJdjy533d24KhlPvDCqQ5m4j1MRbbNjV+Er
wESd7vYnOJ4poRKFYym3w2R6osL/uQGulWnBVnOLiXCR988faM5fWPz9VYJLvq0s
HFgoi4uYVyoEnG8X/VzSxENzYXSWfXNbQg/HaxTxNsohW9UBoEqlODN/oNrYbj5M
puDm2DztOy4P4HUM5MEonYMxjL2aaUHeM3SsKyb2BA12ztWXQ1Hc7cgJfhEFiaiU
is+53ddt1bUI41wGuH7nvDbKvKwUXri0MRPD5Kq6Nb8MFa8BQIZCU19QvsieBK9A
Daeo0oEVAHQVdURj3QI8eo2xOTr58NbzeEmh32QcQwnDqjJltptOn4gGn3Huy3Qc
9BAkxHmwA3Cy+PH2qro2h1xE5hY+EdKRHgDCJ16ZQfPLNxVZSjcxsYi9xqx68Tbw
jfcFKugx0r9kYm9iF2TkBE5ApYD854wV+gKuxvWCd/f2DWaoaAF5HW+sk203r6na
iYpw5gO0Njr6xFblWLKNXF50UQmPzMujMoRvBbHV8uKDM5XtvjZGnuYZ9pXdKscp
PDcMAhlB+tGNDVD1TSDfsEk33dKGHvsJmFOpEPP3PtcPhze8RjBzfbkD4/vvmbp6
Fr1J6ZsgW4vYtAnl1u163dUnNZIouccWhc1L0tLPEj2e8KKP2hX3xazMiAiwsC22
tC0z1NAKtS8lLzhOi0bweKgy3TykipuS1LSY3W0poZMq1QY144/Jx8ud8eXh7YnT
/449Dnn7G1yj/VWlpDZl9yl7r9d/gSObW6kNrbzIS6cpYsBoaMTKRRiQakq56kJ0
ZzwozhiaX8aRzCpy4DotexWiwHqnX2MkXGIu5FB4lWNzIhOuABIZKrdEz0tP3MwY
KPbg/fhK1JMkFiGxBGRpYn0Rs9Ygr1M/CCaReVYNFTcjWYnCbuZaOOPn++ZhTT7f
t+ewLJzmxTXNSA0hYuidN/yXlacVuOUoXdKI2gJ5wvMUgUELj10ATWCGnko5UQDg
UvUr2PL4yPvlXqHfu+tVtxIMna1/wDpF7XGKLL6XDuD1vtfFuhM+YN2UX6b+m/Dn
fpC4ENI3+RixPnpGjqJynSsA5oFZfrrJbT6w66nTBrqCdIOQW3evU/hY4yEvDuIN
932ldHoOZ0+HqssqupwPIICM7twPfcCRiOBsVnhvW5qownISHZInzjfnctnhFl3E
bSB7NIL2GNS8kWkYTmI6jBS+aV7Ex4aSzX/YGeBX3XMPwInLXFiaiPHY2guGFMJs
t5ADyLNEjcLtVPRMsPZYDfiHrPrtfbcp+pV89BTKK1eTd01JOBvggCg76qCoXZXe
VDd9zrVRL0sLrxgcQOR2/ur/AoVLHPOv7qlO+NdO0VGyntA04bdJ/E4Y73I2WoB7
rYZJWRntW7CqQeF5LFyp9V25735G3+GQ62ppVKfQyeDCU8BwS7Fm+RU5ydA5WMi2
d1Ar3WGGl3e5jlFXf8K7gAo/gbJcM6SwFLMKC58Mn02O1rTlRsn3+VUalDAtf49J
4G1igIzXTtzlfmmETrP76LIDi+JckTCWZwCz4qQYUS7HPRMKdx2ZmfePF6PiHSUz
D6LKJE2K8dU7yi1OsAkjNnRBpazDamDns9wc0UNGDTIAmhFN85LN65DCRnpormdO
f71Z55EXa15Kk6T2V6hWRpFcS/32t5+k7pIzAkeV3tpgxrrOc2mQXXjFNpoCg5Y8
3MNInjT1oRwmNGriV4KzszBKkXYr/Uz1/8fWeSkT/ec0P0gbHWihP1eAZ5x35yF6
DBXeA8HBEgasrU2f5b2t9iWhYFg7qmpdVAM7GZ324XR1gEh+H8Xrg1n8CW1EgjAP
EN1KvKus612hiNqjq+qedo8RRh196iD3ybC4jTBKK5UN6/a5KWwyv/8puTzKQpWi
Iwc/MWQnDqNdJOy4ouAevaXqrWKYW8tIu7dAE4MLOhtHsHo6huSBUcIiyJFlDpiK
p7EXKqnIhclm45OEkEYqLvw0NS0CKTYlXYCsUIMl15WtTnNFvBce6x8Tog+WNZsb
bEjJkJUyurxeLbdTqQ/ZNf9plA+RyKbfI+8Tq1K+DNWpjRWvqlipSibbZkN/Yx0r
EOc+yRZEqk4+d3VpnLWFeA2A1YPwSR1y0Q2yzsMjzBkQWjYMABS0auULg1UgTZia
W9i5a/OuOWA114xL1BOoFpD266UpThu0MD6YHoRy0qKSwOhvdr7FmUakt3zyxzna
Yr6zrksg5gCjwM56ud5ohKlzUAHzIPvx1OOlvVjA0qzCuqWz+6oPy+yvXF8dI3JU
iViGs36TFoxZipCPhCJNgQPaYQWK3cugqlXRckVCoqvRgAPtpErYL9669HJ680Px
F9YdYMAH1OOMlHlXKUTmXclrbRPW6qNjusa+UMMevSG6GkrLeNgRSEdcrfjXLxj9
JPrXJ/Xh70mL6cg3HreK0rpqhpTr5htsOPR1RTD0mVSpq0/AJ4e4rxFfS6uoXief
9X573VhUDjd0jDuunc33tIyOIX1305/6hC6ljJW93FxuqYnKFORPg7hiFHMm3ABH
YuNgt4tjI8XW8O63ELt33XUds+rR3uK90FqizNBuMaoLohEtI/zjpv96B7h5BJ4M
LTfTZKlX15uQoGOjVkewxv2CoTRVaRO/tyrmeUVashqZzrFJJ/Semer05pw/NzwS
Cog+Zi5MmwlUr5WujvhboA6uuQd0tOtmo4REdcP5A6hjXJ8nfKUOIWGS9z9L0wNq
UVYMo1+eyo30M43U8S1QS2y+cPIthhvKVoSSnEwA75HbHQ7HV9f4mc7Ozti+QbP7
ExeHLOKvQmuXyk2arXvdFj3siJP4t0DMeHXazR+vkIPUVTsN+LWoroG1WRaEWCIq
C0F275Fxf9Z/NVCahVPZOx5z61Z9KtMHv5nXv8zManBC3gMFN2m8UeWXTz9snthh
XwJQSdcKJ6nLW4L73RjqfW2MnT+QFe/sEovNYQXZfmmdUrqD7pXo9NBsjTGTIMad
XI7eBb9FyZN/nzZuYszSd98eVtlsZWBzaAnTxVW1gmBDu3/PxYIBBuCcjCbtOlhl
RCPCjQPy+003FJGvNxJwkGPV/z5jA9IVE2NMKYsZi0OZVMG1LgCJVAD5gQghFoZG
MMW4+Z3dCFfCcaUiG2dUmA/pOma6mq9KBpLxrB3Y/QJMF1tQFdI72L5PZbd6RXCU
7uEzO7dy6bPYyxnoHVOxZU/h+dsdYuyKNnqqTYj8Zxv9AvzgMAu7VrsVUikAcP00
Cnoq9iARCh6t//iGJ5VuI2cqKeJlPHDvL27oTdCHhrAezopFzUNAUzAB8gWInldw
0+KIn52EIuH9BoYId2Wu8nqxhaYyYSpEn98I2HUYSRiyzypQJRW725tju3moiZLN
mPHE7hVTTG3HiJ3ueyRGyxB0A94xFPyteMscMP1h6E2/m9s0AFlHNmNLZvjdVwai
lDoSCxGOJ9gwUJ3ehGm9IJ9ZUcp9UcSR3ukpHVMNxYC0mGQRnP7GH8juzsinmus1
VwdUc5oMmRUZLyZ07gB3OIk9wiuU51MVVnEMTPXwstFzogZg6fM1XioIGelzyT3s
AatqMchwI3I/BB4F+HVdbP0KSHudC/YeX1Cor5hOAmxefLUiRxW9JQIzEShzSMPY
5UtcgxDEJoxwFiu0Nm9GdaLX8LnlmLg9+3ODF8k8rCJK9SZ5KJ+64LjhRK/PdkgE
nHsSVX2ONili53l0da9fgWU+lPenQNuJ1SnL3foN7KwidMhgjg/gkLavOgCrOlCR
NJBMsmn0AOrB9ZtSy4P3bb2LY3QZWeZf+Zyd6QiEaID2dPZwhOqHOp3D5AdQIDXg
P3pHaUkj/cus1JHHjSCvy4vFwGrQebUbrMDB4jdyZrxOHCRTGZEgTg2wAY5Oqkjl
HDi8E5rAsYbMewqRL6galgnf/1o37TCGKcCfcf21HKI3sqvmEHBZUI+36O8fnc+C
2iIZeNGoCz3qVB+PWamDc9stPF+Uw5ARu6T9bA2NcvBn59toC1qy+Y9FGBeoO9E4
Td7j8JcqMYjUGMMLfDC1PztPVIp3AB+nbc+GDlU2ZarHycRorX04JLIPGDwij8+v
flK2TNMoUDmdIoIE0NcYcuTfy+OwfM0achRUNnkwZxOTbWByf/wcgd1fR8PNj5ZD
+crmEvAVefkPBXTaZ9Jpm1cwWQ4cW/y6lYQtm4FOPck5lImRfgozE7Ky37mX/eFt
Q9sm1iCvZ5HHzRVODIwhECuweJDhlyPyJCWaIr0gy9MWrMHYz7Z16Is9/AU3nJua
Fpduf1/fYk9Z+5Wmwb5OtNEvEbMScmMEH3pFs8HI+w2ckwKHNGKEDsJimE29ZgA5
urWRTq4QHUA9KeXj6lymvZW02s7WCrJNw8fG1llk3fQ1m22U4EG/SMuvX2EPLBJe
lFkGcM71qWqlatNqCsbUSQ9N20TMlwhCpHzQA0g1OtmhpOWY7YzUOvHiH1JM3q7R
izGgRDU0k0y0v+G6LDkF9WL7wdHkcFZ2BTAgb/a/GbdJqeHuglVvvARs8gf2+dlY
0qw6g0pfzm5ku0SOozGTvHtJTkJ2gy18IzEu1acF7uFmR5lN7mA+IktPB8aFTGEt
YMwWEHh+DXkTGF6cqX9E9lZuSbch0g5NEnZpcb3KskHgnawQpW+7VAHUmwNTq8iP
RPpHvX+xusp2bq2NVBGr7WMHIBbxLy35CD8YO+Wtp6IYgcOx+AH0U7zAks/nlSGg
HZwaEWDeAyOEWnfY7jP12bBpXPjXInoSrJ6wIvenoyN2fKAfKmibsGcvPHU8PC6F
PJJgkeNzlz9HK/6j4naRHGCw90fe1RU2feEU7kNSZ2odA9vS415JOKhZ3mx0dNND
XmpYtkCB2Q6psHmkcSC2VykkaN3BDQakHpQxZu44lkFzXN4uVkIdhNdgYAH/nwYD
8wLtmDlcFWeTcgk8/B9IwpxmlI0EcwqgL8bSdiwwtTBtPR4Lt9Hk21NUPSxkh9k2
yoz7lPHG/hpHgDWtPowMh7Vxyu6YQQ85omOug1+cTQ5dSXe8ZNrNrBlE+TJbq7nq
jD6p57RV5A8VBeQpjsts9N5hObJ+MkrLdgxQcMPuf95v9Vp5to7B1Aa5+DiqyJ1c
ARqGWbAR3cHWTzGjby9tHrPV26M+zBTT53PVCUI9Z4zNhVsI+9qmx9NIVqu4LfvZ
FLUYH7BKMqvENfkzjT+rxLC5IrnOFjKHfGFfZghFq9N9eeuXNtqdwy9qZcwgzY9r
UyxG2w7aSdewNptHeZc7Tvw0JEsh2wawzKyC5+Tf6hXbCTdTxmMMEszLh7tobzIz
w7HBzAnAGXT57Y0XHd+rnmMl/pRwuALSh0MqEIDj9fa6DeH+Vmcnt4l6aLku22af
BBbw4Pkc5qjHr58Y7sSpY3o2BVAMZtSrYM69W9jzuBDZ2FKPGB02ii0u0upGtJcJ
qWJSSar/odzNnOw31i2mLPqU0Ulmmou6dkStHwKG5Z0l7LVEQwSlOAbKWE90Q+yk
WRCb4Ogv0fhBfLpCHx9hBdbdcAlD2cwoRpqf4GY1NOiEC29medGtbV7g0xACCK8C
FXtnbobvRBvA6tJUVta0s9tdei3VL9khaXa/tEn/emZLLkByrG/+IkG0OQd/fAz6
v4sf68JaMoFIfOTmTwAlALEqQsRHPrE3WGY/YHblqNzwFvU9eJ4/UXUu2aJOGSkq
P/082fn68fn7VLLTriybZuIOjYHheD16F63+RKI0H6nnXoyDXh+eHOxETnqZ2p++
rM35J2/20m8XY9PIDAQppo8k8IAzDgnqh4WfQ74nJ4J9PuwFq4TBudCByVMzjL7n
Fs8cjwPAnKCFHM9RlRgGJqKhservUzwy655NCKVWcn1e0DMRKCIxaCNnLoPEkljy
Kg5voNYC3o4wthqMlx72k1qM6EYoj7/QGnBqnNLXie892KWlfMiZQmaqGTfsBRDp
hqjsCgjP+Xk8RMl2N5ad/4jsA1SmJTB0MMiezytgx6Vg/kLQdAKEWm/0tK9VM2cJ
AuuCkQHLfFnhByawYSkBsS1g0bS0tlzLvgCkecYU7zsmbXh8/uqAFxmlUwIZlqKl
DJilk02s30DAoD8kfHzfwq12ti7JN0R5PAUd5uPJyq1RHx6Oo4rfLz7Q6ZtA3YrW
PNsWdT4chwS3gB8+9QoKUrCZhjNONL69c9o3Vni37PJIY30YzyZFGaho6vHRpDH4
LZ5qpuavrC0SmNM49Wg1zdB5a/z5p8rRTOas9Ohk8027LQc1s3+0XpNts7u8ZDUX
Z/jabSs9bPiL7nuKaxUd1Mk98yqo0lX4cOMmnV9kkYIuvV7dsMDLPKNWpWL033Mj
YYvVVEf1mVXE45XirPGNyQppFrjgRMa0/VbXbT8gynCs3zWTy5bVhZjS7ULd25V6
ixDjNlIk3QjGfrflKWXcVlYHK4H5AS3WNLTZZsZS0tgpY8rUkYIyrXcfYjF+ED0Y
NPG34OxTp6ibh/T3u+5wk2Ax9/Dg3/uUPAX+I+1NIz83CZ+TkOkp61YFBmYHUNRr
AxA7DPje9GUxKf5gAHBv0hitmVr5nYPFZep2FvO7qDFWGzasspQA1U5JDNnDW1gn
kfayIR+3QxPr9Z+wHXP4YBOM6atq87y7VM4U3/w4y2cJ9OPe0gSDFe3XydyBlrfM
JlMVgBsxJUvtT3onJoEBzV7bB6D2+Npf/IKYKsimJA3+JCcNF8zt1bJUdOhN2WXU
WMYHrkue5bej2TYg6nerSlggKNkV3WZNFXf0ZpV1ED7sUNec7tiRdFdtX1y8fkM6
okMsI8JgwaNbVk5YNz00WnJ0ff6+3v17OqW8ogf6ZobQ6rQs52SP1OcvvPY0MBu4
64eNRRjP83QTvoYmd0xfwCBuFpdjTqNLiE1d0j67FmUoxZ1BpgCpZJkog3rjCbom
N19P0qQACUE0UDufv/3I4h3MzVbb1WjM4eiFNJj0EZOfC3wMTYEstyHCHAqy/Ad+
Xz72WkZM5tPBKbKGEUTCokQguelIyJcJhdr10LiSd+1D8+q6DR6kvgjhhe9IVT08
6sXAIYUJGP3p9xdmDOgjQJztuM9tZDC3ixoM04AJTJx1kAsNPiwrA/Ytd2EZBfPK
KJM9M0Qpi6pJdh+BhjNV0Wkp9tpfC5KTmw7kFTmR+okNaMlpYkID0tVjkikzjb26
NGJcqjU2wtaxhP0R/fkSPekqtq48TSBP1YOEgMK35y9ygOIdLZ16HbU2WFQrW+p3
kJURcrbi6Nue7i6Nc+NO9/epzJiE2OCS4kqYoZSOnZmIyyEyZmLVK2XXVGcettdj
UfWn4ph+4oZo4RRX1wPRjDDuD4yQM8lA264avk8RvfcoPTi2wa6CCJnBlQeMH3ez
wBdxoWhbptoHZdwad1pcH9xFi4q/QOx4P/YOHt8FWNpiSZmV9liURtGcjlN86pLT
LTU7cN9KgHwWSIJPxpBZWSgCm6Wxbpteq+lgjAErS2UHXmwUqCZnlTKQB0i/+Svn
6kEiIQ1Dwsq0lDTPuiz+iuOwB5QaGyaQ2lkmx14fU2dGcq8uX74lxPKX9s5j4HuH
Zj3CpzWENMrQTI6zmZPo44jTjR6e3J3Z2nclS8AD4ZTZmNfm7jGxvlt94ddrP97z
BUFGFx3cTTd6K/j99VOI0AkSAo8V9j3n4ys9SqVRCq5j+wUM5xb+kmaDvk7JXlD1
+yjsZfRPYHHHCX89r0mThAgQseN0HJuVxb7DthxGNdXrdUjWBo5OFMWSIcTJlQYB
bE1G6Sd/2GMt/H1WmRxOj3k+fisMgHw7zr5Xd8GWZ3xZmewr2uIJ10KGEjQV+8tO
x4NFcGdJdEGjEbSMh6zfRM2LNnmzGVP43cuUPBQxZsHBlxxcKpWhOBDyY14m1JL/
0hSCSHKVIrCoJouEuS6wAL8zPik8+fsnykbxBB0A20EBJzxQIkgkFtb66Fw4gac+
B4wPCQkYml80vS9FEEcAMc38ndownnWnuM7PVQkBBo+JLro9ezJTLTRXRYo2Fj0v
hH+YyAONZR71u/j34ENmre+SRUmZu+TAjECqFAtKab9Ysd6b45/b2Q5Lw55tM+df
9Nl6zs6JuGnHPl8/bBrHUr2KxYtjKmJDP5gJc1K7r0C2dB7b5pFeMZd00tRtgp41
2nRHOf6C4lGj7CI0zMqv/Oyx9B+h89jIAuAdWG2tJcvehvVUz5Aerq27PpgX9nyZ
HdDAa1YeHNJokThXW/fp6oC2D6QmSe6K82Cb1iLnb7+A5buparO2phkb8o7FOhfz
7NMqEY/VbbEugllWlUwAzFsgtRaxK7xjE2D9lMRUKN202YNV208KubWmZ5E8ihW4
ur3kL8PVF77bWCuyvFACJT8fAW3uF0nE9NRlySnhn1l5fQNI96tAxjZlt3vDuV0q
ebTM7hGc0djlvnM/lIMD225eOKD1HsCG7cyH5YsrSdk1LCD4CQdEbB8UTiCNQOrN
WOCs2QuGMUSiebDjjQwIQ4YjzUxsbif8/4M6esAX9gsjONr/AYL0G3bfyWBC/QiT
1l7Q0NTb0gV/SidE+so+s/won0UfE3XEMs795j8s03oqF8gK1BhpxAZOkYNNUcSi
FT6bui1sWMAkXBe5uXz0PZSzU4/QPrZRCAzpkIhnBurljBS9XNeOsHLef2jD9jY9
uqVZz0gpoy+pqsZ0y/5d6Xi3A9S/ICfs0ZJY5r4aSKAuq3NQaQ8e/jk5BgGiLcbe
33PZdigboMWkB/EsBSLTn9j8liiNtjIcUDd+lSO9Jvdu+AtpfQQ0C5IhqCsKSX+v
vuFDtNydRI9E2h7viI5e4dmXh6Jgm95IfDq+5pCiSvf8ukXh4r3dNaFD1UftHqM8
iPGy2tHz8H2WuFWcJ6oEO9kaJsLJnjgZKAABJWwSHH2/pzKP6MA7iYdzcg2CmJYu
j+kTmZI8+JO30Cnx3273g2Z/WDmWXENf49BExZOKOi2j4wK8OCfS2tHb44iG7VRy
gkYlmL3PihUwl9fADMLQlIz9jWt2hKkHiwaPI6/QUOmzXgSktu+Z944JMN6ayi2m
kD3tg/uzGR9319cBuHVPm6e9bILozNt11nUsWXMs1ARvXRUoO3ymCUngrbnqlK4n
VcxfnHmJpjKy1hW0+GJGcEPcbMSVX9NbdAI9dCUgkom+gtVHMV0kNnaWRE5CELIK
u5Oe4JbqdaIThMTCwwnmMVJHxXrseseF1zTW1945Z+auv0o4Mczp/tuKKDvCtJGG
mUI9Myz9VifaNIeweT0YGiH62eDa02iIGfhi4Ur6WwvonujkvLJM4fjEIUJF9iRx
eSguvhBSp1sz7IJB+Nan7qpm1G2ztil5Ohv6lDnySvH7Zqp1s0GUGImJqM4Uv8lt
WNDlY/xPG8KUDAvZZcJA4vuLi1dq6Ou9xubNeCzyQgojGQHt5Avq5bQk0V9PEr27
5BNbQUsmRmRXP2Tdqyl32C0KWdFmz4UyFbJGhh5uqFIwvlE50gfQ5+7tP4iMDkLr
vDdB/BVvd1DnmVBVboOqyKmsGZZLZCfRVnDzkJ+kmmBaDblyCdqOD2zUdgQNNYRq
NZ9zIe1BgF/X4CRXdbLVrStt73TTX80yyw5ddkm1ht7RoO8+yUf2F+dBquRl4FOq
UfaLGSR45qTZkNOVzvC/apfa6A2G6XrUyeDCMDimDXZcf/mnSl6QFmyXq3U4KF0u
I1O1JJAXxzijnz1RMoQdtDc8KM9ZOSWkMI6sZJvRcfiy6cck9UMs9mayCR7CQxXo
IpqBhCN2hLoUp6L3gGzhDNlX9TtiEUyu4F+4zSy7OgOpYdQAvZ+/OYn5dar5kfPj
6lLj07ERXF2Of55YzPI9hBi/fOLoWBi/7eh1uD1N72KjHYZ85bn/dZT4iECK9jPs
8/PyQDm6TkBq0eCllPjDxZwytFI2+ccpMAXTWH2j/t4fCepvjGqmd2Qkd4Tl1U0D
VHR0iyq0/wd99GvY1PUkbbaA+yuSvhWbYH/LdsoLdGRXwve5x0z43Dop8yWjk0sv
57m6ZPSvaCP3GynYwjDpF16APOq4/JqVaOmNAF17WMXWlgPZ8+PGPia7rKonD7nU
0koL7sI79P+91luTbpaWFiHlVpJVq/ugFuSKk4s2Keg1zkD+QqMO4Y1j84SiuGJR
040isrIMWGbLeWmtxo2Gn1Yx1P2C6Lelh2YoZ26dVflxwH4Dz9wR3jbEsUXTxwYh
bGydL3UTxO0AGEkdS+sB+MqrKxRmV1FjqzZ6ZW9hEuHZCaO9lOXksjKN7uETHQO7
xmBkKJtF5nbxfUfehJn8xplyfuSDoT8M04VIgGVoVG/p2/vkn92an0aaUC+lCCP9
SQG09I50Th1WJ7bTzssZRZqUs4DuL841p6FCgRS4zW2u+TfEdJsygjjPnyecLHD2
D3TnXOGLLz2lkItwuaXeeYAgI3VUKuHko5k3o9TWXc6VLVbb02AlWfnEZ9+TdUX3
Mm8h9ZeWkL/3d+3yP9+StAkGlpNu1YW+4JMQcJSkmSc7vV3UxNg5X/df9QXqV9ii
Vdul1nmCMyqv+xyeK1H4HyNVb6TMe7vc8km9zYhcPBFqOrThhRNrsSgFY4M9wil1
nfUrSnMj2WMVGWEHdDZdfk0S+sRaRFTtF+G28ok7J5cpqQZPw9vmLnKFyM5O/8Nb
UJbhVAplgzf9nmMw7x20xC4RRVl7OCuw2hxYgJXArEBA+XImpOcIcR/x21Kewv+S
Mz9Pu0CMIqZzxvK/HZoXVZKM4eeE7rEgne3xnKlxMD3ZcygbF27FTO7IXLlfKsl+
ja6RnGpi07TG7XX/1mz9xCYLdsya6M8mYWycH7U8oM80SCeG0wTlNu6v6cmxylGP
Je+CDaD4/ZdxfkjvmJsFF3Dh/xALswguzs+m+95arVyyDMi3RyDShnk+Bs720hVi
FQmQOIPFFFgco3/wVC09UGB2Y9orXJwGL9NxFn8TPtOzrKvjGMfVFBepbze9zwRZ
uFEnOes4kR2ihr4ofqN0VJbi6dzZWrrl4+07YPkcLJR650wWDkbu+QXl8oCgosiA
r+EtUSJxXsYbNbGhkDn15ARpN2op6B+Q2qHo3PUG1y8BzCP4VQwoWgnB+OYA2bQI
wgRun+YnRjqExt9/VumIE8JCwhNQHCnczy06674yKKAAQq8D8mJUoGIPcrCtYMS+
eGCUqkq7Ziyol+HPT5DHm7dmhkXJsbTIDYUD2mfIf/eqV1NjO52FP78GCR5nzAS9
LVb0ZJsT9570VabxvyIXnAHFkaylMjvFpqMRZ6FEOdoAbV9tMtiMIKD1rAFwu2n3
mFNTmgH/vT9cP1bOqo6VjktlLEa2i4fVtfzujh79uVu+6klbLUUXYxVJUWbnfzdx
qpkszK1qRY+eG/4QJhL1oG+X85e4Zx0IQW9nVG7NDE6tjd8OjTbp7ARBaf18D0bp
L5S/Zd2hHz363uE8iro1TWhiMBxcVGTQuv0X1HdfPA+wr97OUGFWu1YNbzu8o4OY
sMqcAfmgsVLjfs+cxZ0p3XIWLYpwKHBRJbuTyp8bZKxfdo+7dCBvHrBN9FSVJnmp
CNfsrsqYvi+r/ayNLME0pBwaNkuKBXmf0y64USB/PANP7kaLnCj4dqLcxidc9xVb
EYD3o4CWK3oINR2uOcUPO5B0qLIqcbF4VKXKFd+PNtrMAeucWC9A7gqVIZGtzhzk
+Dyx/UgSviA7ag2onOfqoO2pSufKdBqsOmH23JpDpvvWj29AGTwFOP8cQ/9+fCWt
uVi1Uh9Z0HLeRZq3TnY9MNWz720XPjPddzGteAF78Sp97Z5LSz3LRfTC2GYgNetU
k9FlrLbQuw7DAht6PFjX2VwvL1myqZXO1BewKaU/QVSU35jiuoCgVfJQfUFZgf/h
cFp21eFJWN8sVVizkfyvllv7Vdu7Bcl0YnagCth7ybBV9Hv457OML7o2v9MhgMFc
XvrsWhBM7s2hJOsrEyTePQOi7zxUx/mBDQYDA5OI9skQDzWDD+pxBPBwb/DY5VcX
jxm0z0hj98HowFXIvBtEZE4RIHlYLP6lFY0pgzM4u1bt+quYEBq63toAVIDiLiep
LiCSjVa6c/gxci6rSn8KhSAf5e6dy2wuT9Vl6LJ2z5QytIJ7v2JUlxYIm7ObAF+P
5lkz2+zR1C4T3O5caZnfSxwEF11WiYDQ7oXJGZdHQab+9QQem0ZTN/N8NbyKDcRl
03Pqy0P7jRUSDrMUvrMYg8kDnScH7x7tEWFKeWd1hp8vszCZgwIeIY4rlrWftAqQ
UksQL2rnCeiqHb8Ubh3JWqQqnacDJQ2F45f5z471H2NWA7/WBJvcYfZdop/e0cJr
BEMadMcv4+X/acDG0rsrrl4O7cMGeQeXkRTe6htuMJ14GL9Mw0HzsIdW0e5WRJzS
zBxFpY5qlG4n6BQV0XE2G1PiL2aaYaJWxMfYxNQiLD1MX4A19/976JJiVMgZ3gRS
3fXpzs2HLpxakJ1EKOaUB7cOV7pTeEWMa/IX7oev4D3A3bkHl0NtHtPLy2ZNbrL3
iQrf2e+aQBkvwmop0h4nFZ9BM19C7GMcs9npkgmMGNAEkLpOWviPE0xwTP5MC5ml
0wpXagyVCFE9SXcv3NH6gxV/CbNsc+jJi7hWMPJBJi+ytjb0dAHcdY5AKQmrddkc
7u0Kow9iaLIutCdW18L+sAkrWtm4mYUefOuQMV9J2QNKlb7OyCQ+5lYgSGJxL6ug
3YwZZ7uRc0JWNeuan2ZGp00WPwX3blkDzEdlfaQ4FRUNABkLGmgVtXWzWP+/cItj
Uykwj3bsDIn0iJt7KYqTcHM6//uNeWIVSK7BM6gPtHQHVB/b61Eeer+hAKcM1DB8
J2sKubr3q1aVk7ofoBs8gp8a188VLMuTlFCA0qgAHLAy8IhOZ//TdbEGrqAPXg35
a5820duwa8IEgYzjxzT8295O42FD+fku7OXdmjHLVg0z4m2KIOn2iO2SntOKWVRe
NfHIT7VzFdaQ4AAOqz0M8Bmg/hOZfVu/pqQPTUMM5DxiN6katg5UBFCRM2Zy6FGm
yi5gmUz2a4jtypr83Tc5LndPXWZFiDXjZ7JQsBkisqJ4qxr6xR8rCi9K0hbeKbJU
4+95mw9RiHRLaX8hGeTvz+QbHAkfqZEFjVF5Ynf9kP6UlPjt02d7HX9uAKKbcBmA
eHk6yqHdy/BkDSMZv9Gb2SVxaqmwMpM8DbM+Nvpg7o4dD5B+Ox+JxsrjDBoiY3Gz
GOD1ui0m/iOPNHu5qBLaUimFYqgInaEHwz9nl8onz30zKjdvZo/T2GebVzKi3LS6
+VyGQaPK0pASdLLAULWWMY8l9EqHqog61jUBzxxr5jCrG06tGIEKgLMYZyf4OyXo
driKgO+6eO0uxUxtE1P/UkYLL3quch9i8k0//X+k3ep+5hZ7mixE5MbRYsBJBsL0
OEBhvk7Jvaj6vw5q7aS5IHdeDoVhMhBuM3a1cbMw2psCEkPZ7W2SQrVtw7D59LOb
KsogLTAN5zPooDonq1EeHQw/HenCICw0enYYJearHPvtVbl0Dz1Cy0D0u6bTNqyz
1MpvmbSGNEc9tmm3uvbaT0jb0oCzOUFs7gzwkGFu8NLu8neVcmoM2v72DWp9LdiY
7iPlx7+fZpMTA5CBMHU56ybsFlSU/b0Fj9lSgd1QtRr79QJm+W0Pt2ZDP32NCN87
5GTfXH0Y6IUmn2VpHszBDk8b6sKVeOOKeBo9FX+72NzwNSza3zeQ5QQ/uQ/wXsCl
NFzHSAnbT1OJLHH600ORVZmRLUE1QXYHvSi3tXKsTl+wPqYORG9fD1jCSwxJFWjm
0QwfTNe6ROISrOj/Nk2nKPoUzvBl2Yee1V7F2zpj+xqaS50euCq9raGmLYZFeIEh
5zNsWL/CBqeGwLyDpHhSsRjOCbJ6wnP2u8Cp323Eqx1zxLf8Oerlmr4Etf9SQYjy
O4YgF8BR9gYo8IDzyrPgQoV8r06aWYZuZ91by6GJ3T5FA8CSrSqB34Sx7pMdvYCx
MftKuwU171ae1uuRN4al4vN/67AUL8ytwyH/1XopsaZofdWgh9Pvrqzsl423i1ix
3xASxDtHPp36mTT2hOzmLQpZEucKkAc03dRYPg3EjZu02ZIuRONVagbUCjYjNH5g
4yg8WqdRDwOYTqwlCZw0vh1qMTB7HrH9LB24U9BGs2+9p69B4VQFRA+3Yx8GHD8x
RADst9iZI0hB23SasdZ4R3pWnqNQ3k/xK15xe6swKYyLxp6oBkDeV12Ll4N7Su6t
qQ5GvnS80JoqFJuB0dmWJM5EtStQVeP0hg5fp4LK/U4SWVDTCsKwIVe+Sn734qCC
q1t6ZtN8h8+Av1eDJ9eJPt19CB2r59xlHYdXiQe/QikhlTOHgltKlWrpu0s1/FMw
`protect END_PROTECTED
