`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1bJgosmJBEhsfBJ2dDKQmdmvSohq1LPgSV5m8d37GkQnDQK0SOIOH8PslxTBCyIJ
taw2aEjcSIyY6CnEtg78V4pH4yMfSFwswIx067dsaYu88zHwA8VheCnvUjVRNEdY
D1Gn8I3yKvXELLQkhl4pG5uGqo5Nelm/q9pClLOUslno64eTAx5wYQdoggIVx0B7
+AD+8s1T91TxO0s9kFy9ltKvcyAykAvSnGzuxy5mQaCgEzGa6Nj+cg5fLTof4f9A
Rzfteo8KO9/t1czHvw8Z62WaL/XiEfUiqKeG1JUbGFJ6Px9kZcqdVQaMtDYbVZUk
QFTYHNmtFd/aCBlh82RMpbLqIHA7t7WtWeRWeGEyBMm7HFoJmEDoRgvuiOhP6R05
fzPniuJf+kXU+PddhALizBZMoHdpD/2R9aCjc7un/4nVgR8doEdboCOPDO3WS3zk
TbqxOQaYIoB5wNuY2W3JS0WlVcWhgCg0y7+Pdgjz1d9BTN/ciEFT9W30VhyDcE/F
pxW+jl3NWmN4HPeMRzG0+TiqzYpjiLzJ+15Zcv104EMCYGxnM+tDH1Ko0xqYUd2D
VZmZDd6+S++GC+7Sdbn2hQ7L/kbr6nadruQXIkVZsPc=
`protect END_PROTECTED
