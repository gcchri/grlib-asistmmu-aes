`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dPgy0vjWIjtY/ZlHWVHliTiEwGBbQRugUAJSgIi3gX3aUkQYX694cGeC/tCKhT/+
Sl9ETcIbwImkXy8Kyg1osNoxHrqbB+Kor1iMIDySOU7HmQ22aLRmTy2qaS72RZOV
buUlYmgaXokmcrMwW70Pb5sJPjs/NA/V8qltXtDhL08dpkGdojY29OYJvq5eD96E
IIRIvpKK4eaEjT/cBFiF9tAfmEXxzPeSVu/Td1eas5uGsHjjy5L8iw2+LJdrqd39
7b4iFpXzaQy9Ypkg8NzkSH8+XNCpbbmupwX/eDRtMhVYxKHilziMxxyjwr4gJpdD
YRVOhu0+TWPsVw/sd9UMPLSjeyjHkTSnq4BZKBJgMv2UMJtKTynFAGkMpWG5vgJE
MbDwp9wZsYbeF5AV8m0wBw==
`protect END_PROTECTED
