`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gjnglx2koN0QcBx+hQOTpPgzFmaln+7h2Is+HSQ6Iq84/LcGK/YH9mL2gcqG/R8D
8rWITCVpczPCjJDqs9+H92a7K/lKPZT1PMxigx3ZiAErgPXk/nOQFOdWM/nCO7eO
EbOc+ropyFAJRc0pKW3LZSCpZEbk/l7cury/UOPw4QaRTEqHN3tWMtVYjNf20/Yl
BZ+unibyqxCAzWe1MAdKP0vGIU1mp2RtuikZfi3AjG9ZmNHk2NfuJwyPnkjrmsDc
UeC1kwi+Vqf1wugqdjZL+k3WvB+DVQNXuovzKKGErtIwv8Hg7PWASaubyypEMpFc
jEgnoqH7oUft5ZRlHxdN5hJMiqsuXMAbZVf4RkNPJMGQSSXHXf6FBZfHhptwt6Se
3K6fyKhQi89+xVVDZ0RkimD4OrpF0iKPUfWmkxTMLRZXrCXSsk1hP1Sj0ENt1X4J
O7xMPHuma+6bHqmx4+jg9GKGbOotA8A2paEvmMBXanex1AocOcQMNYY2S9dRpQLB
fAFCK0TUA+NU9eT5iG9KKYIKG23Kv6IywiQ9pXuTRYMInBrgsHI5cGNmgcQHWqV/
/TSyji2tSXy2PcjUNnrndBHWMTmSyEr+wI45VjYPSOI=
`protect END_PROTECTED
