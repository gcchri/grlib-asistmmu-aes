`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KxSTR68ex8VFoc3uM2xgVbLq4Uuxm3YBHQC0/tbaUgG/8iey6jAvevCk6cGaWxuQ
YXJTEOoxscKYV+GOfEsxT+juSsQhfXAd1ZG4Joio4eEl8ZD1WGBxmbswp1l+rFX6
VJgmH7WqUkObZwC9zm/tr3qm/Z+zO+cLDxpD+x/n3eoEgrcPL1zyMrDmmgRW6d7x
aKXjq2YJDJ0zT0Oj5N42yNdtrkrSCdG/XnA/8ymm2W4q+JjxKOY5OrRe512NsHQq
ZB8I8nfcn17MxpxDTp2JLqmSZd3Iak8Hl6G7raBzFBcu2DNk135ZjdjBXi62DPbA
xNDPcYkGvAnCJJQqm86iEdNq/9k8S401SyZIrusTeBZJgAZtQGZUBL2ChoUZwhtX
m2+/quNEhG8GkcTc0jb5KX9ZxBr5ZrMMQPr+lCu38MqPF0yJZp9FCgTAz9j32b+z
57Xv78nY0nQM3Lp/HbZmTVGsSSHovzHY9nG7JSgOwSzDBDtzFQflYD9WpM3DaPmn
UdrRGYT9d+BGYf5Fo7bCHpd2SEUJVGEoomyedUJ+BBuyV6q0pZxqtlZ7KfBZUBqf
2Fo22WNBJ8r3km3rXLu8DA==
`protect END_PROTECTED
