`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qGnfbsXvX7JiAIv04LPVrSYnMcn1d8gbHxDqECOt6K4aq1lByFij6NGc8BTvnF3Y
W5EwXBcfMkmYegc+vLfkOM7uCT+tbF3J36INj4J1LahQSPEljHyAH1V2/2zofmZ3
qE7JWGB6sebeFodQdvC4HdTtVxbUb5y70kVpGkEYZ28il67b/ysFyzJ6ylPKpopZ
aqTbsTFf5EJqFUhQAomSZryDO84/Pb8iD8VTj48ccmwwifci3T8nQYlv6pPG0N8I
3H5mtNcJXQ3F1eEQCAnSkf+pe0Pf6WpkpaXrNZ88Ob+hzKnjWp5+qDbKuvIx1d6v
GluQCFZO6Ua1d+4rQVq0/3KEobDMSJcBC13uNbxCBUiUFf4fqFmCDrmm3/OslIU2
7xGYshx8zETBh5tYyN2qP09lASi1fVfhVWg7HJelkQ5RHMY3UMuZC41389OVoHUv
xSwa1W/DYP2grS4rkraVNRCu3xcmv19w4y2XQypsFXMlY5Wm8O+6Cqkx6nWmMLeb
6rUKQvtz3vgLvsWEkZTiXHoctcwYpTr541QTocKVU6C0eEtCJPDyRkzlwlGgJoUa
PjxgItc8kjuyZX4pZFtfUw2FP87NIRnPhckYlHX5OL0=
`protect END_PROTECTED
