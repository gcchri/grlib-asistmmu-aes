`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kcbmbRMOxX6jgPZShYmNf41L2LMt0/K26GY4M5M+h3DwaqDHmLn+Xyd7tOsJrucW
Ht8OAQ5jL1x+pmMCVCZ4TIvik2IU1JhfTxZoh2M3nbOEAOgvh3Pej/Rgz8JS5zRC
Zo/Q6uOMpzISEQJ1aK/y0mD1+mShN6CadynH+FQQg8nLhoFSYvxz3Jx0ZrgHBQkj
Vj90fjvLmhDg0+vBM/kGc70KPB4BONQKDOOJZR0Vmm8mBVvrloFSufBnS7KccwOJ
bTgd+YR36sOc6QLrPuNvaLQV7ASubcrwB16Em9SKYntri76zXSken4Q3BjBzAem0
x9GESNsQxee7olWhIPvkfO6pM4fYu/amX+Yhr1bqMLJ23Ai4h5od+ZTqsvB9oG+E
RK+Y/rE1iCecJCytNk++G7zI2VDoJ8abBHaEdx4Lmnw74xTkX4nNZ75oLE7+dsqg
ta3a3D0eN5rET/cfmJ0A9fyOaPX5yDGL2NPmf6hYRBTU4DwNPDoQIyhioQ62gcze
sV9T2PXlExndRAleedbE/N08oJVPm00PkG+nzUhty/yaKQsj6KfUuGEAFI4g6y3E
akBNh6ob43AbJqFejyPvJS2QVGxquDrsFAeq7HZroXgXWSzE+UF2FHb8jLgFp+UT
PePLteIjUSpRm7KgBqFCVr2ymSgTtMjWf1MAS1oTHk0NS5nK0qTvTUonomQZi8jd
aZFPo4TwlGjaAYU/izQuF/y4ys8kFT2O3LXGtwVNpXmFSZflxtWKVkmiYo+NzoRL
OGhrBvFbdQLAheDF8YNCxHuJT4bt09NrQnJW3xF5IpBqTmewJ+KTk7wB+6jsBI31
oCvi/8aBHP9ecF4jnkTljH9Yoz30SDuppI1qox1/FRHct4fyUFr6ekqACmMNMdSn
Ow4EmPAZrD+DAIaLrRyfSYvhtDVcOFKejol7Q9ypqeCDyo7UJXOjHE3OZN6Cd4pT
K0TZ8QFeVOBnYtubIux4aKgodal2djS+8dzofaxwmeaCBxB2YpRKsPKEGiBwtroh
JArP7PLamgUYso6uxGgbRmPF/s48GcC6xQ8u3G698a76P3nkXYjeCl7ClkeVEzXb
aNvnulAoBFINyU6mddHzLijGVzPo9XGEDjA98STV298MqB/UVjC0lTy1AMDcUZXY
G2M9bwqFQO3YGnwwcTLRBhG9K+bWH4PEWzQqdpzv9yUI1MDK6KgD832tt559OUW0
eZUA2Wkw1bwErj7D1xu3q8B4cw5LfU2aFxRldE+Qa6tU58mTldHwQvnuil7Ty76/
y2D+s10UffjdM3BR0NQ5XT8VCg1B6YygXkFtpkRUNhE=
`protect END_PROTECTED
