`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1r4wvBhOFe3491rPheo65cSRbyH7h/i+XA6PQMWN5wkfZo7R/+Aj5bgexE7ygS0G
+/cuiGVo7z6Zbi0gcpvLgpSmuQVexoeLETqSJEnnYBISWD4P3D8wWvkLIVmT4+Jf
O6IkKsK24QyWLlqpfk6TKqBqs0Z5pJwqJMMfyCPxH1WKK8BGXht9ABjMMdP7NoAk
zMfTXwJprhctO9TLhD7Xxm5NnW4XsQPPlsUwhjTrehzA/D2csGE6dXbhnefhpYk5
MrNF+mVRvlS0hbOaLZxFMDdy57id0I3h013l+izZfqyvyZJi6haecECb1rZUmqtg
5gY85kK7CtYf3RsTOqliFSNTRaqC5xL0IxuyVvR6VgLZxy/KdbgygkK4t81PVqq/
2IViaLMqTgxAkSdw0F7FEq01zw2Z/G7NUKXTUN9AnpudOQUOUS9tIB+U7wqUzQDi
FS6dNqlfMfNCXu8AVa6FP8Hl78Rhw9i6xYsrIhsLCAESM27MgFp1d6A2zkiwD6g/
hTNp3Czpl5W7G7wTwa4Q8Vq+rJcESWqpqyp/LhliYsvtUdn55MY7hXcGW9fQPDJh
Bt4HIQGyVdTr3fvRAvlmuKn5Qs/nBVAXjiJRuTGVTA+i+zPcjE6Iw9gA8mCj+5cd
nKQhGov83/DHoPJyaCX/U9yagUzt+nlB8+G2DKDfZ4Cl+fshSBFEgbohAfq8IwXW
8GNNV7r6Rhx88LsBxhIZzkEBqFSMMARxlgb6IMUfJyKZoDJ1fDCqYLWZ4NWYKfyq
CEVk3ieKh1o/9ctvAqsS82CvAjH40fRbEMWBjh1jju4LbP8bRGSpEtUemG0jqrmT
5Lp1QHqLEJ43a8u2jgiOvLVKrKoAj0cnO3aOUFpRIBciWDQnpxKMqxaVOxoL+el7
URqClBereZQd0bfrwK6TUKkEDPJsFhMSl2Z2Ai5Zr5MrNwIgw5UbWj49lHaOlOfG
TeMvJckIOW3HNRTXUC8ZgpRuCFhGKZqPopJsq134VBUPNO++7WLU8KtZcrvn7Wxb
gLr/ZHtmXEuMCI2evasF0StbP9s3qJEFiy7d068TAsrw2TUPUvdXU5XrMVfgX7g1
7E6NXltMd49GxDujnBV4X2KuY+tzw+3EFfsD20iQt+NxJpL8uovjfabpt3sA51na
V5de2HIyOSiGlZV1PnPgdxRYMXOSA53OkO/JapvHF2P6029U5dRLTrS+dkT4T+3X
b7I0ayIluDzBsza0coc2gN3sGOQJC8r/ZhZeoAq5SD3RhT6dHLWLU/TtWu3/QtlT
hL39IWws+aV7tiUAgAMWgqKAijyKcosj5I8BmoCOecJNEhamhvHxqiFZ5LmCrfbF
P8AGsAWCzWw7TJFjBNmQKh2PmTzPW48bkN4q/cVarSbU9Lr5oTEncxKFthjOKHwe
JviryNu3XCXc9qfbUGrhkL2RTMbtnCfEw4R0fJJI2PcYI3tg3ZC3S46q72NNLFOa
/UxgZQtso/5LXBgN7UIysex6C04jGfLyQsQ5zMHG1g5YJDK52YnkoYPK9/TmGU05
MbIx9jIN9LTB6AJGe+u3doGk4ZN7RzOHk2zFvX9QrekZhFqpGFqGbGYB7Iy7NyG/
lUaQlmvONkbjvu2Z1x1OL3bhol32QMce5d/Lz4YwFtvuDIZHhcX6tw4Q4qCmqzqY
Gb9vD3c8MdJ5Rsai+d90x4CdraLr7FT2JxJwp1DhrbTAKwjwDQEkOrsurOXndAkD
cIt1jSaTG4DPhX272SzcExZEKEWDCiFsmuPkA0IpldmtlsXrzuxLyCKAT1TmTCI9
UivQhlrd4ylYb8IQEYODOUw05CixHZGJjXDhb0DYC6EfyWG0pGi9mcC6naGwKzTI
ur1RJWO21+DP9/9u4yrIqhRrxtvweQdCPfCjV3AVNATgFWQBN87PHnjHYKEQVCkA
TF05TAkGr84gd5dq7AiV5VkIYXxIVVWbTESp8buesuMTfE9IkuFy22Sv+Dp+iw2M
zd/h95blSzxhHDFJGEsbQfPBMCdxT/hPb9cycGyeVA6VZCvwB0ZJa6qEyZ1+VLng
UMIpJLO0hJhqwmE/K/Q9f5CKv44RL8peoO1YzJLPvGxOTbhUyDUuifWhsVv0DaCT
ExJrMVrk0nRZkZhak8Jk/lEfzOqpmNCT67GuEvUdU0/aREJf9s5enI+8BxHBbrB/
YOr3BTENUuUx6JQLGC9JtVBKNwUCd3NeSjrkOlzArfVG6fr03gppWiyax3GxaiXo
8HSuz2yafhYqCOQgmMxmrZ7eKZhxlrnl1cm+IxJMN1FKPrJWGLog4usxknnr8Qcp
zqeceUDZA1u+xLn576jXUadEW3dcSFNhpJfzVyuBU1hFnhgrVi3IlXDT7HhLoMAI
AR8ZrGPUk55iFEz3dTvvkoz2gDYdmgJ/xzGAOv6/ZMRLgZwcLzNBeMINDh3sv/Du
LCGL43Vd0jllWzT3URkMUM63GPSPkSeZQ4ZbPWjhBmr4BTTZJjvPgnXWq+fIyGxu
C63dZCBiKgp68R2eN0sXTJRLi50IkLF6nJnlQH1IP/UO/S/zUiViwbI5Fh/c+8aw
peH0ghStiwvZQdAmDf4uF/isP25UsBOhnOKA/SZirM+AY0zXgFSIkfiERf/fy6dx
30mC+HxHEIFNFEoaVrwDfiPD8pVfmCi5tDkNYO+GcPnpLeyqtZ5fvRiNBtFB1/qR
SIyKVBB8qaae579sPXiBvLGwFmPaxwWle/ug2tsN64j16yN7TXLKeYtJ7Bv2mi+/
wQqcNlP9PXFBfS/wFU3JXtbvWuepLfCns0XkkRPOpAwcGSK5JEdbbjr43tUpwMu+
GkY7g27BbMwNeNBfWnsjJpOKOfxbpAJVbByfgCCAcZU12sa05HFwwL5Skz9kBDSV
UaODL64CO0RckIP0afBN9dE0i/DcXtV3Hqy0QunfYx2A7DDTAqIyKx615qkX9qCn
VAmXbd3ottBl4mwc1zOLVNPRCmHBqnn58ICETtMbsIMYHWVx7SQy3NkXKC16a3DJ
qaSwpxsp9lcP4Oq3a2OJdG4KpK5ObRPPS76l93BofivMmeDapU2mILkdw6a8I5Xr
oLS87sSAK1hjlvljIS2xZH7X+wEUeN4y6TZjxcOmih7izvfXJWddTDb3CXpnstCy
PEfCZEvqme5XG4bp5wN2+SQbFIDULzG6FAxgMfOY0d8D6/c8K8e5nUcByuNiMVWG
EuW4krVkdC8CkgKSsBxSKPQwxepD2jssMXWJI64kA6wUqlsvriDgKZESQGdrLsln
06/5OCckVXWWZQMrg+2fah6GRLGxmomkalrNSuIhXUr5m4PODXdIruur5B+VmfV5
HnR4VQWVcTuj8doMMVTbybD5e8WS/1q6AZhuvsZc3+kHl+LYmLKBuWKwiNhWTxpj
VjHfEg63+usMb8vxnXHKEnySwrQ1ymEqNOv/IOzHglNHb1+PzhIFWrDEZ1pER5jN
Ddmf0PyFdG/n3Fz3Lg7Le6bBhB2HUANVy22VGRjnlMfL2sSQ6axX0rSzykM5IPD2
nGv8QkpsJ9v62HCY9oU7Skq+TTso/9BH8d+smSrZjdI/eFOjVDVzUExuDoNQrTVX
js5Y/xQ25dVS74qeKqdyZYUpiGmVlrq846HNd4KaSylfggxxILriq6yD4JZqeU8f
51YPw5WDfTjuURCWgztH6K+qobph/S8VZbUrFUa+YU/Z9ciHS0P8VCzrJcC1nb3B
4IwWXT4uP3aiR0ytUicjmmiDLIT9X0I0syGhmOM6wS1lPXLKh4lN3p/KO+FEyKhK
pdrEZepY+f2V+4PiF8lHbA9+e7DoMmT11I35R3HxsThoJ48gIbxkLhNlyRRObefd
8+fu/llNTysl9HlIM89rsvEu9AwfbrI+cZWxbZF28QmyT6FDBaSrVMMyA9vNx21w
qJb53hPdkuSBTRW0KXbApzva6YU/hKQecV5GM1v1R0/Y8XIIACb0GP1+/pi7Rb5t
9BWrau1QU5gslI4OLZkxTPw/DjFqJapPYKSt57vIbMVdvI0wx7F782rWTfiJnvwx
`protect END_PROTECTED
