`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZZ5REJOfsHQoCCVCVlonlG3QYpT9maqW5yo6NE8bl6n3eqjlr4aGNQhXZeHUCqN+
btQ3CfI39BcYdePcZWo4C32dSXNS4YxAhSlFnfWyAVUXtAdVn0PfTFknq3AGV7oQ
ZKrSQI9jBz+3vIhBTu0O1HqStVEwCvocJ5FHTx9K1P8RbVvEW95ziLWVAJZnbzGu
EXRVMzgLvll9z7gCVDw0P1HhpPpw9YjzpJMnSfYvi0V+SgUaD0BM2N+bRnw7ZMYn
MsdEehTIkWitpJ9XL0XoHS2/29Y3WyZp4rp0Lx4GS+fv0fR8ivdr/eOE0Pnu1UO1
UdnIZvdWuRzO3cUEVRqzaV4Rrpm1/3mVX6WV+nLxLrfjqOUgV8nLtnwr9BQzgKnk
PrYb87jWSTDTIVh3cyWEF3YNglTe4dVbOaOc387mzlkuWMDfmzOhMxqZY0y/+z+8
uATta9PkFMXbG/P6Ma+1uA==
`protect END_PROTECTED
