`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8dkTMgpyhINSizgUpcSNCOf2eXHtz/gmYGWbgCDanVf/reGy+mdws7WqpkIsrBSL
5gtpRodlU+VhZ7wehLz9o1gx63YbhQWW0sF92BmsWT7tplSRk64m2wlThAkUwSfS
AvIJQzRZICxaLSSlppq2oXnDKJjXzuH2Pa7G0DTGTtU36dkHVC6hzaDgsjMal7eh
+0jRsQ2G2sgNOiocr67nApvOcbrM5G9mDLB9t/8JGSYUez+y4kkOizOe4PE2NKuO
pqX5rBYOToIlHJjJGQmMe4ZGU74zMpsQFQOiArXALQIMl17f74wMAKiED9VEm85L
fBsP/INAE5FRbrhJje7N7eKo42u90NksN1Ia52chs8TbxyMVNuSfmgDGb0YObvhk
PA4KiaF3bjgoTxQOyjI+gzqMjyRwJR2ADfqMovLA9HUu1oVXhqTUrYWlZpINmecO
Bx5J/lu+ygP+6gIz29apeM5OdVlUOJWWDMWmg2ttDkhEdzxpgDRs6sHbP1lY1ysR
YTFyFKSwkdQzbdvxTZLKX4bJEcwXF2iW9GOvnfnPWFfSLkPJoNH43ZSifsNdtA0y
PKAYjiQBFuxeMbCFDsUV1gxRcj5fXjBesGKHOHpL5A7jLO+D+Wxf+Od2MHjiktvf
O1OtNpRyNlUzlGh6sJKBrOVtwtudWgLFt8EcEdauThUw6c/TUrK8Z4GZG7LBORbj
FBglDuP3Yns/dUR3ICVQ2mnqO9eB3f8szyA7ecSJh+ipuPzVcDIx4j/CXsCmL0IP
ZA5eDhPm4y6plwDqU8VaQBgKAZy/Avso9j/mQOK0EM0OCrTrjYY7ceSMJLNB9C8D
F5SnpX3jb9v0giGmrS6kg/kFoPI7OdCitRn1BPfgWdjrQiCZFxkLG/p3AO3YS4k6
G3cD1QbmDl8K4P4KF8XUjReZTUNOg9NoZhKr0GVASaQzzSKRX2p4BeB3LArm3V4i
d7fnBdCtUg+7K8I3HbXh/93OU9pYO1GpoTIKTI6BBW4=
`protect END_PROTECTED
