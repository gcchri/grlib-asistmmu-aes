`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h43sVwMe7hrM7PAicnByvQeJdIQxwES5tgJb82KtAj2JkNU+xm7WS9EQTbsIankT
O2GsdkuJBTK3kjwK/KpcQ2DtdmJDA7l9HSv1rqJW7bIzYGkiNUgLCBdcQ/R/KX6C
2G9xmAysw1F6EF+fAn1wMu96GQU6Mee5f0yKwCGsoY2jssCsIPLWS9BO2qmwttE0
nGXXqAr57mP3Lasb2OalTSo6moLLEc4UQXE8RPrNFkqnIGuMqaaizAzs6wm9kgny
B+b6Lc8vTbbb549/bfsdhV2YPYYsl2GVVRUi3ueRNt02eT3pYxrfRYKecPKaNfkO
Fj0gYA8vTFk3Vzk1o+8sqKBVa0DNdfpLabEjyNEOX0gJjrDhbz6TTOuM6rZG6U7V
TwE+K3X69Kg1tQPqU0XSV1frLWMNcxzc+tzs22VJjLH2Q9oRv3VRbGJHU0sDo5ck
zRH0jZnZjs0G8Zhtr9iFOT9pn73OQnAtgvHkES5xv39IFaexckyenpvzc5wJ0kWu
AFGLFwMk4OCqR9no5yRumtFtsnJKTwkXxCJLaEGpcqMQ9n5Nw40Bh/HBN3wEgXZp
CDJbjUOVZxLP/naZz87SoCMAYhJ2uK4l290aVaqUpcBOPhmhJ6dzeNuZLbTa/cwR
e48SmDHd5hgo2rIu07Xtqrcg2m64YGAI3KcY1x4UL0t5eJkr+ETzHkmz2o9UZHbK
MlQNBg0L438C2pCyEwfglyAZOqtGjjXxqkWOW1DFsGmRom2+ohQiiltM92iUKXy5
Qz45fD/77snBTtoDbbK8TvnxuUd1/0lEW8zlhSle7rvNUuToGn7JZ7HrUrZydWe1
x3y4DC91TBXtgbScXyWjN/EDGJQrk4pahb6IqZRu1TSwvFnqMdNWGAlM+4ma1OJL
O8f+3dsr1R/nEzbjMrr1XSb/iwUOD9QMY9Tib2V1mgdIk7tZjiTR9XeKic/ggbU1
U2dIB/ZzqDJY/sPzVnneghIv0bcwLP3ZWghg7F3qxF58+J4VHXUuCyQ2XU8k9jrj
vCM5edxpcdlKmWO6a+xBzmj2M/GF3Lr9hRNxTyGc9j+FXhDbwW8HYNcIbR6uooZ8
ecff9RKVWexLP2fWil8k3hIJJGn793KQEjf1ZpPDWJthEOo1YtTW0HbXsO8+vn5p
1tH9jqbibwnw0A161nQk7p//Np+60m/UNRoy9oKpnuaoRCld4YBqVViJqUTbHRg9
S/DQaWzwvnwlsENJpxyhFxheTss76O9FdXwFsBBfb+4kLcALAnkekKInN8e/mMQV
wP87kUY5of2S4fduvlKUsnXHvjnWJE5yNBT2IxfcmCKb3iokxO5M+503dEJJAmLr
lvdZYNSYXVbs+0LHcq1u1uBQmPBscoEfUeNbf3t7yl+MpMPsdhPAFFFLKFeEMTdJ
EzIggzyrQXXcjScTCckTgL+MqCcOUHkPigmejc7rxjoBbnMwP67ZWz4wP2S7+W6m
uso+dE/NEsdtOyEPRFvYIVorJ1DVAcdyVBLCswe0RVY3O70IgtYj4K41r9m5NWsS
ydPnlz46PgDSnQDQS13nKcmaYnLKBwGlFz+SYZtorZQ=
`protect END_PROTECTED
