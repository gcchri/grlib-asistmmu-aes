`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gXzDsXrKdOU8LSVIrGELM81m5Br9Uw0JfQUbvMOPd8mBWpqe9COXRaP8so3nhDHM
Aio4TCZ9lXIFeFPZN3AmX9Uk/qoBwbwYniCEfoOCZtAAJIg8Iwafk3Kyn+FeQVma
Gd3KSY1EoC1UsnSwq9oBTzydZpmCUCa1L4DVt7sC50jfsyKY+MUTgmXs0lGQxm9y
f4ORB286BW5z0spSCN7UWCamtYaofcDiAHDO1My2FPOolWJyxUaXplCWLM6btKp8
ppgqzju65G9ZTbQSoL0F+6HhssBuK0ov9D1Gy7O437xwPfQ0SnE5DCB08qL2f99G
5ZC80XU3TKUwtPRfq0xOBdoCZ8UB64xbc5TUIxfjUxtEnWjSqQEffR9RqLXPW57y
m4atXf52PAym7afiGJoGbKZATtg7DyoUi37kz2SZaoEpMzt6ehSufT9hPSrr7c8X
4zlHdCI4he1H+Q1pih7CA4xqkQT+iQDFZ1Emid8qjpoiY3m7hS2MfdJu+C7fyCR/
JqErhEOUoGB/HrcArKK4wTIYOJijYH5fDVpK9iVUjtVYS/Do6kf5HRsU7aEa8E2h
YdxiKSDzyXb0UD18l0xFPvL6qq/SmE6frZzMUT+kqGq3HtwHgFTQV+37nGUMihil
5xB5bUpShgT8wkLbl7CyMA==
`protect END_PROTECTED
