`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
31qhDs/Tu+/6kAXZzaIqHENh6Bmu9jDH7VyR74tYSqr/gQqleCzo8xyWeNHPFWBn
M/G/mcVNBsEwBrrpz5BP8EDeXBOo48vE0noDnW/aWu1/Kop9hb/bjkLiZc2TzGqy
qV6TJiEBmmjeVEdHEiuEI3wcxLbGeJQlElAHXUF7N9Gn5sVPo+HRJ6bHeihZk6i9
Qy/B284KfHsFsnEWD+fH7mWm8k2larnef18O8PSYA4JJIUyWcaZeObUxO6FSMyKe
wPn3T1tzq2Y1ar3kIHTKluw+XOIKRSbI+96i8FXMmnbO4unpDkxrhTTNr1PpxVmy
Z5pRi8fgxgRx/ZFBvb5sVzxNrAEJKHmSrEBCWZyntPMyjgfhgc9auqop1k2xVoUg
2g5/AfyFmEUgFSHVjYAqdkQYlp5EBpoYMnKbXh5azmCZw7yEe1nh3fH4zF8CSvWR
7+8YGqqiMIvqaWBid5AalamIqx+M5rs38CKaiHyVLo/IER92bk9rb7x9NxPINEE3
5w2YizTeCkk68TJyYKFmMt9PmS9sJBApi7fBpzo7r4YRDC4GReoR9en3nbetsUqO
Bkn78I3TkWfRYbIvXw6/Ga0I3muvp1TJIf6BJ092+HWUBCPU90mqJCvs4AfB5sF8
DVwwUkV7/B9/b8OkRTmsUNo9kWhLgPv9Nt8oRJ9Yqqoim2vhs6+O78UpsyJSrR5H
nSPGruA0/vMsdekdtAP5zOJLRSjID1BaFgr8mXJqmiDZzWxJlg0u0qCrNyBzFktw
A4VG1hsbnRilRQmx4Nwg4jd01472XfwewiCvmls45Y0Vr2kFGFqUyeXJDiep4NyU
ufysw6gUBHBoyMcverNHn+z0HbJCPAv+43qmyUtvBDQrVK/29xDzNRCau7RGX2hK
ZhUNK55NNrt6vc9IGCsw5ujCQ7b8Xj644104azQuuw+9l70N5zN/5OJ19WcFYAAq
fhLb4Ps+b0kqS8CKtGC5Gm2S5S6s6jrIX/m4Ol1+A5SQw+kYmZQfsomS8wxjyXtG
RlwahRo0sOGZt6sLpJgFafUal8BN8gjFyfXpO64Stwlq7DlwmRHcm1mgl+bSm68L
lHsn+jcl9/y3nmy6WX0TItBdtXzqfYl1vgGLpXGhnokT8r2Fiq2U1fA6kxrz4OY2
9cRRLlq8GghNNcQOdpCAS9TGHhuHUOo+acJZb8aUEe9Nd8s83bye7fQgIEkVf/mT
4SbOOXpdu8roT3N4BaerWYuDaHnEV/DX3RsxaO4vOGf3nX2s+tyS57nTID+Mnl7f
zwoxEtdiosYKGnldXhech01rQ2NNxBOKI9/yb0F/ZC32DuUxBvgAqRCy78U/cNXo
qTsLurC/pkb8c2mxIuozU8jjd0BnYenYah3p7bgMw7iW43zrjBTpXKwzZysOdHbl
Xd54vu80hEzQKsHpDzeVwhFPKOYKlcSw8CKVWVOJ0w+egNK5MgR5sS5i8irmVmB0
RgLc8fvovW8ojFsiVA1HsRxropFbX+Y6RFcHWtWuL6TmK/gd7eBeS0HgWSaPRjue
fGsba02853S/ZBEWaD6kd2HeLPaXb1mCfV69golsCzf4xKpsddoZMiqfsROndMv1
cbI9W+H5QZpfFoswtgIA34eWp9wsbkrAqY/qvkX34egwWSRM+lEMdIyu1RtX5Ujg
O//n9cg2edURZNya3QiQ9m0Mark6czayVDggYC213s2UbCYOgb9ARUOm6o7f7MjY
Bb4AyFUEsiwIWwZoOX+2dpiOCIoAY+KJuFTC3esptvebYeRKmmLlmn2P7R+kJdnY
PN575kJhLcagMD+HzfXJ6F+YV61U3Ed6H93WqycvNi6mPz3q2SSZ5vxz/I/2goZs
IQKkmnqg7pvO7Y86sMcw59NwDrOLOsNBOGmENvVpKPHL5lc1t9X9Cy3XdrQqzoa4
1BuX9lCfaKx/rvjxAfxmGyV3fYP4ktvB19EU3jIya/4syKIIr1BUunBaFQo9NdnS
VOhtv2z7x7i2j03nkx/rbKSp2guM8VysbFOB94Q7sB7C3NRg5wnAv670JMbTZI9S
3y3Oe8IeFnCIDY06dIZiy238UxtUSl30+NW+iPwGAI2tVAmI1PttNYiPKqjkeVqO
Eu9ZDgBaz1jTmDymLiK+hDg1Ou8HgVKDy0KRMJ1A5WF1TFhInphMQgoh0bG/YUBP
fGEeD5kKZF9fKg0SSBPaF4FxxF5TfgmvfqJx3Pt1IUhM5XJjDA95ZYVVW2A9wJ1T
8MxPagMbGosDWc+pYaTdD4/BVTRHD7aOrXCQLi7inZkje5o0AfzWb7jxreWAy7Hr
53b2C8vdHwIbKhhrgnEvZ0sY8bjlxgVyIjSh/iHHkHn0/3npW91J/jsle20GYkNr
ZgmsCZPYOTSewgopSM3CuNR4JftNPbcuLvi4KLsg2D8Qcnts9QCdH2ZlGFfJcZpc
1j8DRgxsRnM3um+8xRuCG1u1ReZ8RBM9/BplnyO8TBUAkk1zjb+n07KN7vxOuI5I
OUDfsMnUGPDUWrt9Cl5/ATn8tJIF8Z42EcSv5Fa/7hdBFlFmvRpKdFXFxJOCV1Cy
FxGMF5LRJ6ZPtOElKDGwZHe6J05YZ2LPNRkNtVDw2vAp+BqwS7JDqfFl276fHSUq
aUnlNY0yhwMXyc8j/7Ag1hHkkoePI+rNA+Z93w42hx7prBVeDnfzcByLuMLfmgvs
gm10880qZ+rhzOa9jfu8f8rwJg1gUMRmfGQ0pXgqzx1X0HiwdRLQ0g1J1Xf10vvy
oDF1x3PTW3p8rheRCWcWtqaPHh4YJGegmEk0D8I9LOAk6f4S576X2W00VC94JaWu
vKGDNZ9O5eHNP4B/5smIwA9ef/RrspecCF30rZzNOQvjZ62lGxsASCE0a+kzsOK5
nlb+xDGhfRxzxBYtmtoRT9mXkCpZ9hOugI2nkTGLWBf8LsWBe8wVdrlhrcx3Nrty
iQGoa5/k44lsfQtfNkba9IJGoehRuMVLOP1hn+vOjbPGp23iMbrOpES+KcTPwdfy
pagfrbp9YYGKEkz/VZ/cgvonVt4zuGURkYqvBs8sYCfSDQo6HrAJIUIgctHCecsf
SZqeuoqnMD7i+BqU/KvbTpS+vEa0lMnyqb1nsJoRmZdDxx5CTbnOu/LLqT8/wqGI
h8Wq6/pFV9JkDWcZQU99rcv8V34iAyV1DaKrCcd8u5nwqrsRpT3hqV9adLl+fp9g
rmfFPOOlec6njIpxDZVIQlizT9edF8i7DjL/k8xS0N/eqY2g+9BBP+syLbX1ewas
L30ZrZsapY9bbLWtQEqoJZHFdtJYK2yvvX5rf5rAZLIIl0CECxCT/BeOVHU7WybJ
PqN5PahmrP1QeLmVpz3QC9c7H9KKQOg1QojVVvL1ZqWbCz+HwznHLSuOcSl91FIA
i8S/YVuoXfCIlrNp+wmPG0tK6KWD+fOsQMI/0dV0OcQC1zM9jDVER+nuGWypZf+V
xUg5Cf4dcFVeNDOcNnZToErDMwj7VTdO/tO0RpvJlMmvR80L4rMawgVdL0l0QIZn
stiORRUtWkJcpFiHHl03U9mueWkhvzbbb4DgEzJBOgbjQwL2/R7LIA5OxhBjuzaB
QtoFU7uB8P647PFQWtazVPXZBQTSY1Tvxl1R/zZ8ptr6ly5hyzFRnJLf2GLC4oJO
8MuGHcFvD2vfx8m/I+cjtORqGSvJNnUPdCEckCKa4SEs0fifbagiD7S4PpmoVt68
5EbsaLC+B9FIMyYXiRG0+6jQ+MQ9j0ltMM7QY6GXlF4nDKmtjSS65OvpVYPslJ9f
2OoCkV1yVOXvSiFxpNO2/wVfkbNjCYdoNWKWZDpwhedWRWrL5ng0YWdVAcwcKKlg
O0gXmpkMytUowlUyX4nid7L6UufEXmFi2vAM+4EAC10SzNKSecMOKyrlICHRqRMo
R1taLceX09tzca9sse5EC75y8+F6eqHkzK0PLMlrmicknLfvaKd61C3IhJ1GgGn0
Mq5EkqAKRJU/uoZ3+4uJiruUIgBfVWSGYwP/j8OKfFtqBcUww4PadLhJs4faNzKZ
VPn6LY4wTDa+3EHuPM+FW722/ZDOEQ/ftIssqdteo3XuIhv9W5j02ATzypqlOTfc
41jOG8+ckTWTPSczdSjb4Olf5vVh7mkTvdIcnUV+XKTzuDSr8woqkD9XfDjtK6Wh
4oyxTXoAlRmeiTRvh208Q+9TDCthTqxbnxt4IouwbL8adHjpjZ0z9EO28W5KkTQg
veWiZoPXTOpBuYUapUaGE7gCbeep44HZiM7md+cUsz7+VNusPBz/AZfNa1IlrXfA
exlXSsI409Z+vPgekx5xaNSsIS9qdGmDeEDhQzWPuQrd5VZJxe+Lm45RWShfEHAt
EDd2CH1E+PtkwTlb4GxSgDOmsTMJnWOLJq51OHmcVWDXQikCOnWu9hd48sGwWLDI
4TZUnqw1yARku63stCqI0Pg3egNdCfX4gNoz4aS3omMFGU8Mi47AE1EsX2c//Tfh
Ct4P4iQX2b4EtDS87STk86f00yBr8N55EJdsxzMkDEB0OtZmWPf/V1YBo2wW4q3n
Gn/AiFwGChAofA+kNhnaa5yhEJ1h04UZv5PZlvQBqW3RuXVw90n9CCMVv+7EDKwl
JjYTNbxrys+1gCfR8nUGXutb7/iIHwHhAyRe6G2i94kKN339IQZe6xA3DxR3W2Sd
0pUIhLfjWVaHF7Qoc7WlKitsykx6WtUD3jj+SMSO2I8dwOGuRjH1nvu48zasHpP4
GS8yyTMJ4aqYe8+GcQ3Ds0SME8unHy+ZWHe9uv/99a6GjNNkhZ1Pf1+WpTEweSnE
InxBfDTh3DfmGEj36uhGdo7eLJFSJavXY/DexAZ1YJrlyAs8/5R+y/mM8+Ip+zvZ
eOJwPXq0bTZIY+4es56jghBNu8Wlh0WyUbJfU5hP8Rl75iFYMfprt/rAvw4xWiSB
svV4qAEJQH9ZIu4ekVMbYxx5OIFM3+QTMrd9Ts0SyLxYg5CQpE6oM0B1n359Up3K
4j9Mztv+7bdihyGpdzLELAwPHNnfqlDXSNMN4zxz9MIbs/umrXGPkh9jR+sO6pxB
aHXfOguDYAbk1unBIXF7PCvUc336yFOKYEV7JnWXhqVcF07DWldzrbm/9QiuhCMJ
gHXz+LJiNPl2IFO0J0pi0f8phMj3Z5CSJ0Cud7hRjrgA1qD78NlEcGhPtjWwejGh
XiwG8pJWR5YdEdqZt/hhJP3oR59tJ/akQ+J0PHH7eqDakOP52xluiLT36zCbAZvD
59ZPYL8YtNMhuizXLIqz0WGYdGooK8jHZ3htXD/F3yzpH4EGK21h30knIVPgGX9E
Wo/dCU/IE+E1+ivumd5N2QGYg6Y9ZpnYNDbz/7WT3pQljgmRSgoD8CJDUK4GVYJY
kXf4Xwjt2oFXq1+0CTTIn9HgG+7IcFwiJWRjfAnrD9TTSkA3I8LZ75NvclzluqsD
B26laBip/mI/0WpNdUItYjKnPY7byAP+Urz8i8vB0rJEq7GfoKg+QFbLfo0B84s3
qb35Ol6jgcUXi+m8va5qzEIFIqabLwo85q+VdTmeGhqrO9uqUO9SyEMjMbdYAbOM
Bagsh/4Pdlc0ISqAF4lZbItn3PopSTU+UlII+64K/FulD0fM4Gsyia/NJkjbpJgR
tyl5wjTZ3QFTcrYgILSEIXSMLhNBPPk0A1A/d0VVq8pM02c8goPNmpyBY1TJo0Sf
aYAyTzYqYv28zPCA2TWi9F0Rr246NhmUeW2IFFDB8cfYgLkIQ9vcOAZXGl01y1VB
OgGn26EbGNl7iGtqCvl3yqjPwpvGiN3FW34Yp5guuiBwIhVzRjk9Vbkbp/zX84bP
LQEyuSoE/IOTQ26bN1zox1xchYpjpCLTPmFoF8c5/Wau87/m0gif93NcfYMK1rS7
aOIGZd9XTblG3gFK6oX4lOdTYAx5p0m0JRo4lFG5UD+GbN5uLTu76eYgdeWlMawg
s7A7mbXLzkNE+Sc/L1xstlAEX0rgcZ6xECgY7srWG/kssiwvqVHaS1hL0sku9uCD
x8V8Gd8fP1IolZINTCBr3IZIVQ4yl8VYhKoqq3rE5HdzYcwTJQZo3XKnLcibjegU
y38V5Ez0+0COA0rfdaIKeFskTy+wcTlJi4dthdGr45NjIIe6m81gQVE4uMHdUfxW
fUojq9oGS+V2RUewiUVP48SeVe77IjxN03wC8IXhkhQaGkkdmHmXobzv8K77PDM8
kF5T1rgbwUDNOmDuI7nbtwv49tq2WoCExQ0eRv9LjL+AWTMu4Ub90R2AFXjzCpB0
zUMpukPSdXbcXEKjpHaQprLszSzIBiBd+gdQlZRs6qhd2kfBVIhPikl52pLoXn1Y
r0BTO+QZ6ljgv2yKSknmJoSBl+zoSjIK4++lWmC2RN+Vei5oveH2aGXgBSQEH/mz
GyAOomn/LYnMt6M/GTSML8VxxObJ+/y1/0lAPf78ef3jr7noleMGaBqLAc9SjOfP
wLGQtthiFP8dGSuI7GK63DtmxUcx6Z7wJlFRUOFoQNTnBSnT+NPkirX6mYZYQuMF
/XQycuXjCKQ9d4h9sU/KNtZePw0a4p6qf0cxUNP0oSVVldjlWIejYe7PNa7xuXMd
L3+Mgu/PoFEb1EbzDv0gSc0rf2TAUk7HPfM0QMXiVBgbPVxYqy/cuJJrELvR6jtN
DCwoX9bDzDkAWmUoBY7q0hlCQ3c4xdqCXvyoFgPfoHoDl1QV8OS5rsjs1R6NKyMA
Z0Nuoj6rfSZo3QLvmFgLVPukq6A4SNR2KCZ+JcST5cDxQBUpj6FHoOhPLhFQBE5V
2UlWqK7pCOqU7psSj6Qbe/oMPkbhrchm1r2Cc7IYopEcbvTDqmuJasSsXWnI7ij+
gJLaec7A8WHcm+bkFU6yzFhQje316nrzUTEQcBU+sYNnRcKSY6AZBBBqh6s0RR5C
ojn8H2rMR85PzyUiLUhXhhQh7V9ZF5TaXhnqWFJwBTPlQ1kJuhNRyemH1bC1hSZf
MmTNpAqRLaYT0G5b629h9ZDNLmmzptclrHiv5Kmt+KlrES3Oozm58yReeylg9qU2
xgi+NCbuG9Wdhq3ch75Q3n+vZvx6pcXYRoaidfXpxxHuXJsRT7G42IwHZUsAMJOU
Egd9kkAJuQi1xuQJ7h/lWvlVcaHTKyeJlIMLGR2gLWCPLHBTKixnpfcfmmxVbmNV
cE+UcNbR34t2uHXpyviOVjBd37asJdakl3ZKwEPT5ICN4oydH+Uac5GjIS2Zlhla
4wFE4z/QqVR4cDvCwAJ2B9Gru+YiLlrrIiw+7R1+9V3daJ1A+UcpEE/L8Vx9kVu4
qv+Ola6oQetBNrju7fQialftI+OW+zBFW+/pRG49g1+Mfpe5IPyYPxyCglsLL0QI
0lWf1YPDVwA76QQMChpqrkDqWi9gh24A/SRa5mWuknAar3Qrj/YXN30YOgox+BsV
n/3WKmx31pYhJkKzJ5zrpgGJaugAHFg75FKui0mIsWEgIRVYRvhU7pMrPxK9MEDp
FGW4O9UFIWuS7V//pcNnTy0kgz1MxqzatAO6VwaDMTGdnKrnwpr1/aCgG3mnChnu
jgTdejmC5MTtKwg5Sqb3d2AwnEVw9ZwvNCtaNVX73H4lS5rOFdRiMq0BjPRPgCZL
UlrEUtvAbiQTM1ykF11AcrSu0W2sAf8ZvLRe5S1XVgdfUmLshfhtBWAim35U3Gzc
n88r+bUEv1BYHXiaSokucJQxx+dMmwzl+s5rzD4kYFWLMa1TU2v2QP1XNWZGNK7C
m7JYJsg+FiCIHQnclTpbPoXoT84GOymzkRKqeNVrmXvcMQ3yH7/dOkV6vEQ1Gf7B
2CWXUmSNF0A8HUxjbtShj6lAizLcYRSSiNSvrxl6gwt111ZPQlwDRACm8oYtDBOM
yoj88ghRYCXTKYx/eGruZn5s/WwL7SnEsVg885OHNo0dgw5EAWzRP0UuZOApxQYh
Si5SQA+nSNhPEQHg8N5Uqgbms/Ceutb5r8WfsWZRoJXEp207LqNSnbW4uPOAltDp
cZsRE+UA9YsL6F9JClmH/YobLzfSzcx2INfGtxa6yvE6a2zAtL+oZO6M0yZ7LWip
zkoVjRSbHp6wKvJs3xLPMY9gyt2NcGfYUtXDfqbUJiPTDpDKwOyexxl88TyDAU+w
PFhV2GcV11//KmowxKVnE/2eEhPT2KQVSP8WacGb4+6Hd/QZBDQIu50/N1BbwppA
I4nqoFlZd35lsbfD27Npf6m6Wx6745c8LEv+uvTB9DnuRyYCwflwfO+HFfp/Xtr9
80L/DOVEf2aRc1aGn8He3VyljVAWTyjuh5ftbg2iFIKu54Dbl7EeUuaJzWgPKJQ1
CLbcmJ329z1SlKEr20uD/Yc7XUJ5btwdSkyyERRaQt/n7Z7EMTeSh9YBbu/1/bKR
lQ99BoqD+uu2+BitIA/5/ISvkPk4s9Fh/NlwjhaRcXGQF90HOvLiApCiamBEsWil
M2F6ae/5FsHJzUa6dtbAGCkehX55CtUC/JLYWJhIO59sUKTd+AdBva2nBbNvC+Fp
C8pDpLWkt3MDe4vosC8XWzdSw62cnBVOQD6yQYJdIh29oxQmntWBfPy+EIzEJnZU
BY5eTyCwEbANzaePntnpKaRXukRw7603Z7R8iluo6AhjVowhQvTbIkkwr3OYH6Hz
2MXAtm1pz6CPOjOZuF4yWee22jbyWgrsGGk4+ik69chx5vis2XpapaIDNpP91vT/
B2Gy0KZmyqhGzHAeQ99AsKlbJ+R4xgccn3yeSTxUVwQwt1NdZtJzwGsylP6MfRmy
lvAsExT4EroT3Es0qdc16gGdDvHFFVoD6kTaO1CvUYgckVFByzn6e/f8Al5JTyMC
RnHMA+t2p4zeftbQnH8p1AU+CSu6iID8P23P/mS0pn9zQxLaFnAYZ2ilngfUXOHk
bH84FYpE8+TdyLxSGU33V9JBa8GpA8VuK22VFmWSb3QvwTt5vabemhR54cpjP7US
6MEXbzZ63KaWQTowIMTTFQ60033m/8iID/MiJ+JhzO+OzeSHP5a/IzOe75mLmpSa
E5z3Vtu3TEc192pH1ycn/YNZ2wi3UadEtAqO9egPot8q/zDVfYPQ4sfngjBp2onF
5UgE/iy8VJIC/myj0UKZQ5MdAcSagCNpNwt0IPfrz5UEtd1+1BUrBRewslA7IApE
ImKka2uxqr+L4bxoQJMURu9+JeaIak2seOyZO8GtugFxTErlE7ivO/+HQALWI4uC
m9wuBzUd7MWq3gRZL9HXpdmIe1lCJOF1m1p+erfWo64ag8jociPmbx7niUomgEzh
KM8RwCO64rQ5y9qkMQ8AMWiS4X27pEawwwy4wXzwBm1MgWdweu5A9jx6AgU4hWOP
Iq8fJd/kwWMKXpZttzmhT96ZEi7xFGkxg2VJh9qyKchzSFBvsrYLIwihLjmZpDMK
Ph1G/zeoC3uUaoAxtaDa0qawYlEgVV0pzADM/wssu9XAFnLO0aLuMOqjEekoqmE8
FuAmf4ii0QfehYLD94uP1DoBOX5LZHeI33gO0F2yedEWQNYJEykl3cYYHxxruLe7
ur6idQu0ySIW/kup/+UCkVoM0n+xxx5tk2OkDXG01k8y1KFjciCq7PoOPQvKuqv1
yQLrdBsJ5QpkhogYo2I6s/a89sJyCUqClY7TrT5F0VLeyWO8UI3XIEVSwqOE5m5M
XAZ4+fx0boE0UAUkHsZrW/TjcZdMbVntw8WrTfbopKutQJR5koQJN9YkLgngKwDY
mJvK1ZUMtHxV8s5C8qQllz1Q7jze4LUqeI0Ig6fNEHowSLHc+jzcVFN5R9/zInF0
7mPJbe/ixI3CfQ2mhVXVxGU8Qs4d667op6d0kUnacNIH4Kk3xMsaAfffPiuajvJu
QhzATdLMY8qexjL0km+Lwrt4KHd5+sBI9eg+vZ019MW/9/fbs1g2VVFQpdPTph3e
TxXttJqWp5GYJKFYg15ELjYX9PzVBjRGFZZ07Rc3Glyn6HjzCxsCCwijYVJnMW1Z
3JMRc81i7y2U7JS8xI2XboR+gMRFSRIHfD0p7AskGspDLVscOiWs5KyzQ0KgXxY0
hVfVWyESg4oYb+PFx+ho9bX08zm1EwXg51lAv9pcwFIHulGCt7rf/Clnfuniy+LR
/y99E2+M1F403bNgzu6t+/UyVxTDBYbpKIWa9wjvRy1XBm2OjYuwaPgclK9tyrYY
SONUlHD+JMJT+RpY5yBHcb8oMXZF4PgI5shf+bTwcjqnst2JwNleHJ1riQoJPk8c
M+0dHnltdgAyUTNRuvGARoUTtyViB2qRO3f9FR8AOoOqRsRw2fBkP36QFfnfXxQt
aaJI2iZdxYUNnUUkQnmQrLtAbrnzocNRIFF286vCBaAbOCEQ/0z89N8t13+ZXJx2
j/SrslekevxCDYDDqxrEuq9987rJd42kibUsK1weVuByH4zRSrx1o1zovMNz+MtW
V44QMvhG6WMXtQAYuvT/n2XR/ciEDeGQ5QZlWyDIwB6eOrbM+LRm1qeE2bzdgmff
mr2BXTO+PSUWFjW8RkeR4/cxIgB5g1C9QgXp/uAkbfIKcHZAVoohc7N9dkPvtnvZ
q1GELDryuK31mYzR5EzEViaYT6NAWWN7H/E2hN7Kb+l3p6KMXhB9jH/uE32mPa84
Mcgmv+i9iy2h0+26dlsx9eRLRFjuUBhrRyyrhZRiC3yAN4JYQzBpeW6HiRy5h7bu
hNTx2SfsqteUzXFQFMfkjiE2eJbwvH9V4WPDswsI0VX3KM2zaObjSJv9vZGhGy4P
WrITrrx2CJowPjyNBXe9mTnto9mVou0I4yrtIGDXjE5jiTqeld2qNg2/4nyvCAE2
Sr9uSViKzn2MtcUshjVFZwr4I7k1CxKcWKBcEfIE+1KfML11F0SLt6dP+XFAwwxu
MHIInNgIZZs2CqsliIdxuszqOfECYDbQJJmR1VKunTt+21PuU3Xna3qAgGX3jVpg
UavqERTeJi6TWL4+eEC5+tA8hDuumEJmEQeRevxaqRL5CwfoQqoIzss0Az96Ew4x
YXP6YqGoQUjrJKt/FPYnw7f2CXbDWYnBlBsZiFNEurbPoLxyNWesXqxXl1vw/5ps
Wi+gI0nkPexe3VrokFFIKj4NRX63BdnLH/6/HUmPlYEik+GxW2JtsKMl8kHSVo5g
rw9ZUsXpAgfNMSIZcCPTq3EliZ5OLsD/0mnoL4WOyllsU+eLnB/2SC/4cdv8sTxr
HuHle//I8DB1dkT/CPj13a89ozzTSpNpKmZS3F9ZjzPOFQ8m2GcSb19iZRhJQ00i
BBAk8dijfJDFzxv8KCwGqbernREEt6nNuz1SDL6lTGygrAZL4Eg98QcqwSicPwnD
gDqaprTQqZhF+Ict2d4HDStYL+i2jeV0/ccVhVljrnsgUD4ksSAiEg9E1AHg/MbJ
8cgmB8xflmZecaHDwV9cURSnWpRoCYi5J76L7Y7LEryOoZ5MwqNw3X7BHL6QFPHR
AM52ISHOQVrxZPnE2UvngI3fkKOjbiTn3Pfc5kSYkHexBseK5NnQdk5eNzh11rTx
wTxRAAqq2nRnezgph7evl5R1l50YS0BX61dR7q77yBjQZiPwdflhjFoOHAaDbmhw
b2gO0GMKxJJqZHJ0gvDI9vFEVcN4684BvWHup2q9tCN5CYucm3GXspPSvqjETveA
tGSEgoH9O2skbqRrSUJxCIQsqJtIittTBuS8JAD7k78CSKO6LuDvhZbdZXsQZKaT
39u2y4kO3hVxSaCA4yxZwIxWFDhWvcawS0kaEd0/K7/y8YPfmdhUu5GTYHDa5oz1
2biyyMoW0a0QYgQgiw9lpIuAVgC6bCWP3ppdoc8gL2DgLAPB8RiEhA78QhOz7V61
PWEmXuhp46+P+YzJjdoCz8PofZfuF0wAWMWjcBOQtl0ZJBajOWOzHsKttwFvQa7d
YdCYtofz+vRcgHaczGtxVUQ+aNmPmvsGZpbhOF5kC+GCJrocrm+gvDjVAfIiEkCn
/tOqPMJD0gY+oO9/BfSWC6GfQD7Yv7vwGcJeNpFiPZcHWAyLhiBje994ixGnTOyT
ilqKsnLS3asJOZIVeA/EHfJIw+7daqXZUmeVGwEdr9cLRU8yvDYtkqEf23UX9gOS
aWh56Im4+hiR6RMVdQdHpF7ioABLMTLIdtLzb+A+M1YqW4w6aTOkeRG1/ADn7k+w
6aAGlX4Y+sZs6zy+aEx/S4uvqu0CaVJoBgMflasmzdw3w9/U79Q/CiVlsU2sntKj
lzwYiu316ru5xKDTyVHtyRjcH9SVX3i9SL4I3z/PHhXrH2G3v4qChjQ48RUGHTuM
jRmPGHDhNwNdMS6YBCe3Fuhr17Zl/Mb5zxRfycvybOBPSLSWvQxMBYJFcVJe0soj
BWAE/Q74/M5xphAjCOzluK7y2ADAIzPFRIXdiezNSw3B5pgcRGmd30opUVd7Y0ix
CoQF1KQRcohD/JCqY1r3/PnCX6l8yru1HjzWEueh56tcLHFFYm7hTIEDJQEOf1lP
KeYiq9Yn+YHjcl/NJgRCEdXj6X57hDiqWwmf1si95bW7dBbhpxsuTo1tmfCUeCR6
+ixOOWCbNfokO5ZdfxfvfoQkQGKIxK1UQYnGKhmM9fAyQOml7i70aMeXSSyn+zJu
F6JqPx4hgCG3iVaso3VMGrJYMPziY3nsWQ5s3I4JSBj7qSTukTZuCXON1smiUC7W
qXRODWcCkgGlNYdguEippWv+LiGulZxyKz9keGaONAFVaC6MVq1pGpxbkX1wb5E7
RU/JzkyrWL8Sg2fZswXaHxVVGev/pRFwSrNHFn07bpSCctfSN7xjnrdqTOtZPVYv
d15WUNnsx6ZiDZ3Sk6OOx3TYB8byfPXkE9m+1ojrscNSRES5UrEwCAjyQDijQWiA
u0r1liHRl3xSuYyVsLU1iUghLxmpVfwgKMndladGPMOYQYEaW7ON2WDRPxkfn09U
NEwLsu9yNZPTUB5Hw3IY9mB7dNcG+f2wLPk4VMhRUnzCVUYG2m5/UySnK+Y2cM8S
qslMQsxhsAIYf4aHyV7C8juIBtJcXnvRJ71DqcpewMNOs+oxHtS9nyMfnm3QIU09
Wk80+NOK/y/Ro6BHgIklBsQDDDEybjTBEIZSVGOvgOlkyE2Yj0EsUkAXiCQI7+ZM
AR/Bdq/sULAi9KnBmhyl9CRJr/qUw6cMsDUHvZFt7iESQEEIKkVfEl085Pep/D7y
pTSS0j9tQEALlp7ZRJe/gRbGlc+cglGge7IVH1CZPufbYWztzAlWiqxhimT1PBh6
mODgJ6P507tHOkhPyVu/4pS1BG/H8qAWhITS/SvXbjYA67RJUwPifRcAePHsTp4c
mp/FQatFykBS+BiE1MBU7nP8svcDypw5ORXWwSs6jRJoKp743JMr07gYtQTXlYle
oZjKc6jMa6Px6uEKF6lEDyDsuMFreIfRI+gmYhMh3u901TRGh8IV2fzCpa0WysKb
O+3sBW7TYSwt9/cnScfvT5S7HVksPnw95AAmB+E1OWLuAwXAcuofrGBhN5WT4uDw
H+zoLW89Y5xBNrAdmNB6/AtfGGCqxiyWWKpdzrdYC5H4RB8RyvYLeIGYVvX28Wte
9hmGYiYMnULemW9wx5T3+w8NSbGzCXQ/DF34kR2+RGJVqfjXNFff7KLwubxcs3pd
JrJa5uv86qDv6S9qNW2NV2Z9u3wqkgsVXZGRrZic6mkBwi5F3PhcWP6qnpBXdpHR
CXBw3+zHr8fEUkpRObR/8PfZbr4366PpCmzziJKKnuQ1UIO3FPLg5GlMILLBRa3d
ikZJNwmm5IhAyZ0OCElRNoHcnZIjFYLikXz/HFML3Xqbs4JcrSR6dm3lBwzP0qL3
8IHPLH2MVI3k3AXBqidZdBw8fzuDuPx6m+iE/ihs8/5fFiQnCkmd1h4dhXPJ1C2S
vrtgilLLbBIUtOHte2jc2Exl9pZRbYRmDV8FbG2uuebTwmjXLVpNl/BXM00ir20w
scjLoNyd5WCNFx1Ia4npYuuw1w0fJjOf7Q/oLyjLfnuQnmNKvVZM1MTmjJY95GPv
cXPG4E/m/Wx3QTzUFL4rqCSPnnfnNyPid3lV2bSTgf9BXdPgkZM6E3u5FRSfNd0H
uA+FRh7wsNv59oF2t2l07QCdpRyxoMGvvGnZVXBRWqbAwQcUmMH9eUymj0eTAjw/
DAABA93PbFeg3/4vboaOK8Mpsi4MTZ4U6F+MT78PW4+Hz5BSvCBd0C7naKq1OqMY
bPJoi5fx/r9qz4SLOeXtkh0oBIZXfrS7Khy+fKzWuq9vDEoUfuPSHhk9duB2dndC
syObFljvxdlIrkLsX3nQ3qI+PTnjOm2pxntk6oBp8MmKjD6/HfegKj+exVraOw3O
hacHkfGs+/4AyOje+SAwoInazmI2YskGufIEPvtwiEWx/tpZwwZBqBiFHuiVIISW
/V53JJDx9UnEX24MtvNvH5e1jM1osATm6t8ciJEEDkfZEvE3z07Cf1Xi08VXkq56
NyEBQkQSUmGIOAvktCzSJ+hcVO5Cz/xtg1H3znY9DIyw/xi9EQzvN3b4PBwycuVA
beNCwCDphgSZIavE//+MLpmp1ZIxmb1EFdzysulT03f2EJDquNrHlOmLW76uv7OV
i395zB5b0M1wxKpVPOPK95/polW83GwaR/9LmaBacRAa0iCPIpfJfWgRaVDxF/nn
2/YtyCSkB9rXqKCnLaRI8Sh6dvdfMw5lNQjyHtX6L3/Zezna3bl4qq/Gao1Fq7n0
1JybO7UTBfGP+hQwILNffNq6QQ8lIa3OIIj/DAxJMuCQw9pFp8LXwzEZWZWcvOPI
rVAVp001tIRpKqnp/EviY2es0DMWnushPhF2xifWWCLWB3YcUT6Wwk6+2ez0x+z8
eTiPnzuQKf3bztoKJMEbrkdLoJC8jNkyqE/BNFSwyFxsJSDX8vhOlpktvsK18ljk
Wp/OfKbKt/kEAlT9AtP7HnVrIzfpxgPUAi3UrcjKXiArq/xXNuBWGoCNdmzZKJIG
fRyz7V41q1bScx+KWfYu/AAMUn885WtIMkfwpBUJVtl+Rw3lewJOwSzUU2snjzXn
dkP/PgQzaapvX2RnpHHaH3Dqa643F6+ff30iKaH/IALvmlQrQo+8t1BIczRr5iDN
HktGviMAG/DkUvMMS7XaPnT7cNbJc8gXMP0UnCSr0m2iOqzpTKXxTLS2mMdi7jre
j2xpmBmTAa2DguGF+jQxhH7/MA65hr1ff9H8ETK2J5wQq+qGNH4xxDZJoRj5HzR2
n2FCfJ46aF4mlqMBuVECkLuPDNl9vhsPEgm+iQ5Q1jNbMNMw/VvRGfbMPo81J30b
ucnB9yLHosd/yLMKtJ01Ad04A4oLxOXG4PX03bxCJ5M/jGOR28kRV9+OUQ6qLrnr
Jo4nwNi6v/GrY7gNXKPjW5Kbp1MKmVVmmQMYG6Dzq4Cpr+zE6XGftiPzMpyLd2Us
AS0MydMmKRTG/DcDHlUcsemNKKedwpI+UUY4hhS+sQ9DqkufQsW/Ycmdi3thZCBi
/MUsZQJtziEB9+pV+HZDHmQ/HicMULOoyGYptK1HxkKB9vNtqoBKVDuzaLNnYCO5
j7AH0hq0Vj2YARyiEe53BSBEf86sDhiAsx76A9tRVLyUVB3Dfw5qIHdwNKZVJ+Ks
6I1sVkiCfObmcGapEEv40AkpvZPlsOc5iXu780X9IxorZtHTAhGknHR1XrsiCDes
A/pIit9dT/PcLF0d/IitdZbZAgTSs4+AaFmypD9/wmPlKe3rOJx5KCAUoTa2wHDN
gEJdvr899fNf5uAs/EcK31mVugEJqUQ8b36fwAPOyKzyZPHJHEO/WyuriyAae4ow
nFUqC7JP7mJMI++rN8/YCXMwj72v7jVxTNfRef+aObynjP5XTEk/LwScAIsTQDu7
kCYpJfPtZngOlFBLXprEsjJyuspEGH7EhLnkcbwRRo+nL1zL1YApA/RE1WO3RJLq
ALtr8SbbtppR+Hj3E+zQfTTUqHKa6vbLtp4C1CELq/io2caCbl6d8wJ294MX7ec1
rybBWeDpL9AmNNcMUZt18RvbZvTEiztIkQMHTBOB1J+SoOOi0tW4qBAvEeCjY02d
tqCJOlg/4NKoJcbmRrxtdEZii7ZiA82lC49iD3BR+xxPehVVd+CSef9nSiIJF11c
nzaLoaqyk/n8LkPbZdqnYJRfArZxrTV21K1V7OMhZHDkTKauX8sizEfhKOh/p7q0
eAPKTk0Y974APmH7e5GIKd0Ly+uBh1eAE8yho02bGB9s9RkhFSvlBUM2uqMTgPub
bcSoqTYYtZzTCSpitnqdM0uaxl6nqsaPTz7D2ZYE/ZI7bqGXmyp6T96OPkerckdI
bLjLhPt1koYelDiRk+j+G4VCLGlPJ2klAkSFVfSe6hnbcvaP1sCMGqnKu4c5kXw6
CIONjXZXtxC4eagOekkpsgcBU3+jBGLXODPC88RcYRAXJ+ZgBeKqKFQAbdHdgWlo
7S/OoQKRUp0zbATs1n+aZLE1Lfx7CnS2a9kfu9sdOV7pe5rwdhD3naK0ke/SojeD
WY4RtkccsOD7LD7ibk07Qub5osXL8wIEcGOPh8x5B9gm/HPpNfI/ukBHopA26pro
WdsPQX0wDRW5ZfBho1x2AX3P+VLSlTu5/1tkr7lXJgQrEWaumXyLYyO+CNcISTRC
slijaSHml4Nl9x4TJRRktCkMSJfcCu88J9o6yWC13Nn8THVEh1XTWkO9tWm6pH4m
ztDZCCDfGSeFtb+NUXTTDYWbKvsPArSY6k/qIimg6fD0CNHedW5gQweiiBRaDUk7
TvIQnQ3jG04L2z434Yt40Cdh2fZFJ2wgFOGWYwiw2UoyKQ0ujBJmqDG0Wh3wbi73
yvzGHjYRulD4GdmbyZ/E/TEVm5G/k0bVTh8AWFlswtHUL1zwOmS9Or0zF+/PFlYN
xr1459dUV8Bn8sb4Ii2PmlwGXzbFHqnq4Q1+RDrOjwaWH+NsC9zbq9hqj7aFFTAi
U8waIpgwumZuh7sw4H0yL1ynGbeh8HsTawk+5qtKd+L6laoZ90o/ay5NFKCdwd3o
huWXwjk/snJr8y4uHYhenI/ZAF4rVXfU/MZ5YuhQYI+oWFqKR1bU6b9h3EQlmSHA
NYb5eZHE7RGl9Lr8j0x9aDDmBQHIAbmiQdnFfr6LiySZWnpo4sEwsznCrUifkXXj
OtkIvvsfSK7+Ee16dEcsQ+lObpfiyKxOOdg8vmvCJ51cpnyUTXt1tCVH+7IYfPXV
N2oGeIwH94JeIVjcYsvDaPCdEaYfMWoHPmJWcfTZJRj7ZInHVFcbIVkaRjNgBdUU
q3TJhSTNFwAcGpvTuB3AulA/XxvZbQKGKqgxzj4lV5S+nE37trNXycbrEYmU71pN
ZSo8Tngctc9XIy8MJZ3e9UBrqpuNtX+Aasrk9Y/GcCB5YVSaeOfdQHOcx0aWydTg
EwYl5dcOQeV/2t8HYs0WxpomII7C9kQOzQVvlwd2U9ZqUPJGY1tL3pDmjMmwhLkc
AiMFsgecfi292Qg/6JJyrGBe6E/GRsDcLQiJQVdfOP3HqaTC2ykUCnBloLHiCvVj
U2j9kuY1ZfRIrcAisbmuxy7aKyb+4SrZ8SbzH9PjXbwUZOweJFIimf9u7gZCCj0q
YEiLTLzMQQbcBQUAWgHGoymgeOvBoqNdMYaGwxfQMSB0VvWoQ/qS52rSNYlBZZ9C
hjxoQ2Fp2kTqBFbqr8a1iFIx76f9IKmwy4Qf+Y3BNaSaevaMHMfEgOeZ4K0xummT
6+3xjmcG9XfM/NtdJBjyww8qcnRGzJmbvNYZnl514pIMqR4fd7836YAEG4yvhWbA
iil/K6e7xotwUB68zXXy+n6lyvm9kRv85gRc1H5220IGkWF+IYI+ce9Q/aC8KMZx
g1c8+AFlTcptPlj1ETdCRvZ53OKjzudM2Zh5Bs30n79cNV7aHzIDCodj8Wy75MpO
Gy9dQNfmq6h9Bk0jven9mr1YfKT/hAsnOLtaL6OBTDootKHaQN/+SOvSygFgLjHP
EDNLcQ9vVXj/5mTDv5BsqsTNV5u5Iud7yRE2HAXV/rWbO/C3MaSLevCXVzppuPpJ
OrPOydXGNcPIxf4XSNAH4J7qcPEKgYFF/jE1Zp2xjCbjr2pluRk897kb8lA/8oZ0
TgNZfGy0AQhcAfD/3gGdFOPvWyOynjyBHyY1GmUO7mJcCjd4KG4zfM3Y5xsNGsyX
87Qryl2CEGxFSD7WrFD4Ni7d3+DQ3IijE4dwa+zjFvWa4U2KAkYagyt9Hm7s4NU0
wS92g/qTILQnDoA7LL0mTNGwXbnQBXl0IZMN2l//+0ON6fzWXA8Py7azH5TVRLRU
WL9zZ4/KoNiYxcpQ7sgrLLg1WCMMkOl93izXmtA0BP2iyj68ixPlRjzK82Xn9Sw+
7JKH01nwdXq1HkKjtaCFvZQryIWWqadObDwvpAxDIOEDFvyBW0wf9FGrrmzflB8F
lLGK+6ORUe8jESOKfexdKmJ9VSfSOr9XMF24Nqp0VKLEIHe3wUBxsjmpmWdq84Cq
0iwPsGEBNSB+bwVduuOHGQhEQpfv3mNk37xP6agN+LI3W34uxNtVsHrxLuL458ro
VrTmcMHiexrhtFx+FG71NYKSlsEcKBWrihMyFtZ8BivyOT39ekMYYk6ezUZ85xsZ
H7gSUga8fTFyTNwMOlsiQHRjoLn0Pt/ruB8YnKgREsWgSRXDpOPbwVUfVIRGXNXv
vj3/2HNY1h5noJXTfM5190RtYe57jH8bYz4/Kxqnto/7m9RooSQNpzuU1avScf2P
g4UJKxqmuOmpBd/oHfZj35RBHZBM8lyvUgGeyc7XKBSbKPuwucx0Y9OtViuG/L0P
HjnX+tUPDdxjeC43qyfwCiBMsHqIE9UMISJKYIC9bd3Bc6ji+JBTmIf6+NY2fNuB
9gmdxr1ZLrZWINhylnALL5nqZNiqkYCdXC7UgJmSW+VyCurzSMzz5DuwmmqDYjnF
956QH+gwTkNSp8oKNs/5AHREXklRumg5p8Aulnruw0LtcY6vCMv0wABSetF6uktp
lg0JhZUm1hWM3fW2qdL9OBXjgohWpTt4D6tsSNkhAcs6hdO8sUCQOGN6F/G524ax
p8P/S2zU0cdlLNhTBWg7Q1yl3XBMrPzFmUVyeBiOY2qVo2k8sJFSPTZ3wdP4OPkZ
4LKzecDzTBXsfGT+ynqZ7nNsgZxTjdfx/uk4BitfedO6OJdofEYrjb938OWFlWRl
pT/Pxx0UtEKcvat2FrfNiQ==
`protect END_PROTECTED
