`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N1XoZ8fpOe6jLWQQMe3se3j5Pt4xZitMU7eZNuuiz7d7nWMIFyONIAAScEvdeEqZ
AFrwakYx5t3dzX+b5vAuMLQqcqY67BDKH+u17LIS/11MqkxJsYbIrMSYpa9J77R9
j92jSy3IrTSgl80S+0U/pc8OApn63LWV/PMRh1CrxjlEYnFObrJcv0Q28LzeVPfq
ZAV0B4YeuYUCcTzdi8xLRNwjJ6WS5rYqz1S0SLnhOl0wgbm6KW4ulwwRxxOqk8PI
TtthD5hcPxqAE5wEbmm6d+Jx1xD/cUSsrdkzYbmjH2S56lMtjXN5G+IUudPJ8kLQ
hysI+4ZCkpBrJEtwudOy5g6k2aHCBry+0MwubUb6+4yF2OVrEc8xikxJ8Qo1p2JW
jNifBXI6IHqksakTsL4TBVrrRUmOdG8Wz1MgDm/ra1+xrztOe3TiroVtroI32Uxk
OgKtYtVBmeKBE04bsOpn0pPwngU0LQqtIrXgPIVM/IHQ3SIurLxdpxjgcV+Pg6Dr
xGNPP3UTnqEJUSGJqEyEj8N/UR/AdO5PLjnEsb+ROI9CdZEtKzPzhDoA8wuUkp9S
9DzK7PNIVGR16lj+/VUDVmLhc8NEmyMYlWUOHE+eVWw+tDdPl8RW/1zJjWd3Ppci
qiWHM9OIyp13NQyleu8G7llhWaHnPv7VFQNQWczrwSU=
`protect END_PROTECTED
