`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KmQO2HLirTwejmKMO3LwPnnQd4X+BJh0O95xnGdKWRSIC/hN4fE6EPVovV0HVPmw
ejAZrQHqOHHcM1bQ05EPZ43QgNPKN/W+78wPrFDc/SZQLpZEV43Z42u9hxEWF7gP
4oSKxVw/bliopOE5UOiqJvx3IiftnIegkN/dIRAwtI0t1oVRLsO9IhbC6ydzW9pN
SsW1oGxyJ1I+JvfPqbbx6icss/UiSSxJsB5pA1Nd+JUO4RZ1mRW6h3eQ8dQNaSBV
uDhhT2XqcnmbdCDdxO8jWw==
`protect END_PROTECTED
