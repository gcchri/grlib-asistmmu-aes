`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p4uXp7Z3jO6n/+Hmwd7CPWk/oEZhDoMxT69p77rzaCKh2QX15y+iXph8MyTgrTuP
VfFsGg5+IuUS8N79F/1l59aDBeuNIt9LOwCXMBtTl7B7LJVtmR8HLmYg6R5p11rt
bdYWFO8QVNn2IeE9TD4aR9nD4ay7GdQDXlzI60O+tWbcsWtT08vRe2GiiDejTAy5
DPpS+4/e1vB2D16x4qG9eSsNMIZ0AaAXEwo1aXcn4PQYhSz2dWOQUknQjZxdLPwy
Q2zqCi26iqrONmzqTsMkvCtezj3b5i5sj9Bu1vsSn9Rg+OXUHpUF5fgDnZE9+V1y
m84mSmhWIXxa9Zv6lGe14XDFge+HZPkgcRV0j/D2tTU4zY07bSJ8RJbUL+rgidq8
K/AqQnlLm+q6dHi8sDCzJTH2A8vBLmATfFhZ3EpprQY0dwXE9I2zJZHr7JDvKjfL
d31fgv6U6sPkEZE4uGmaaQ==
`protect END_PROTECTED
