`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6kkutCSo3ly8dm3Tj1PfTTwgnNTyMUaSlK0yFm4cKzxpf6xjI61Wp+f6EPS+5UL/
IpUmBOoaN2RgWCkeEv8iMBhUVamBt9zJGSl4E28pY0B+XqDeeQl63L2M+OS0FtWE
2vDvLUpEDF+CtGw9H/584ytmHT1jlbO9ts89N2BG8IDyN2jHKUNx2jCFr5AcwhIa
ofuR/dQ8JsZ2whKqanDXxDPaA7S+xYvoMC+QermlWm9BMt22wSVbPRjsyThN4pGO
dpkEMUVVbFFkfehbyDEkm9x27rALF7y9WYZZqU88TusfqE0SHrevVVOebsTNW9Lc
Wjz5O2oBTUdv7CvNKGCiZBrFRfjIDeo+dbbjZSzhKE+SeIqzJfJbYZEH7cLuWlU9
1FIQeE0XblFC7jMdAfITMr2SbcS8jxZCjacGdTEqWYfD105LZqooa7v0Si/JfD9y
nkABNCPiizI97g25agtytMjw5MtxfCWt163DoDLXluA=
`protect END_PROTECTED
