`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HrMyQV9pwHiLho83s9uafjSiNC01ZYHEhZ9ZVVxj+Q2NpjRAtM6WoP9AQ5CIeDTj
azgyaT0rJzxQGsi+TYOG2841ZX15glE2lmjjUEtxMdEILBe1m3dRJvpNj9DiRJvi
BCzqydZOz9HfFpjNm2voQVxrftjHbeFMc9MYZueMjpWmcirTsZjPY49qDy9GEOMG
h//KslwJgYyFvGDYesx2VFQMy8iEXwJMB35cvHSo93Op4idLCod/RKWf9aSHLe2o
vDT4jy/vxiBxm26MIZF8IJhnvY5W5mvzKVqdImFEhru+zGfBTJ0fILj5c+yz4L5V
hHNl6wmCTN2FWnIiIun8A7VWaUO3LsKCdxMbwxkcEMX9nY2L1myeKtfstI4BigfB
IhioB6JRdAG/FDn/5obZhEzy2sxHF5yx8ELb6Jt9ixxwWyWJJUYvjmknL1qlHpSZ
tPctendivicmmOwFzp0Wowj8nQU+5tEEzidilhfwLdPnyGchdDZzc1DNfkFb1Ifs
DMrrrtpXhnMJiqFEVh8hCQrEAi4Htf8C01bECJcJ7QOb3MRXoYkEyBkNKr23rfiw
EcyHJ5e8c7FWbQlajWtr6MQSS1uM/GmPZSyDe5Q4+tCL2Df2uGWKBSskysdXq4J1
Tn1jkf6F8q9EBmB/8E3dmF/Sd3Nku6S2y0MxGyyvN0l8JhwXy6ufWWv8I2CwTms1
l9QlaDIriCi5HaHgwmmdbGEGAiE8PshnYEeUtRW40DDzhEZiINobb4L0jQlyitPy
JXAo5IZp4pvZjnl735d8MFVdxuQ1L3VmWJ3nJGoO/jRVDi0sFgzul9Y2o1sv9zKB
6YmeZLshrId31sejE+PAouoOuGRrj1Y9p6eZNuK+fv3v1le8BUO4CPTyZlLvt2ZX
SpXXfXjyN+aIbvqZG5e4/TeBlL1VMrosyUwFagkcAKOlga5DeO9152fwbMBhH6Nh
muYT7Fza6YZ5/hLFlGn0IJx+QoSu0HvfABmeY832hGqFBeR92/g9PBNA9sWPaYIY
djoxz5EjYti+7LbXLD8o+I7QtZ1+U4YfEB4m4Z8nZjqS3B7LEzwhiZqN68dMHROd
UNqBiwWagI7M2HZJb1bgH2QcBh0KVJvYqM3vZj05apfS5wD779qMprTD5HHyToqW
HIU3rF/2L/haD5swV+EVpB2ehcOaCqtqOfrQFgv2BAn0QPoKvqhv6fCmjuxVNvVU
zi/eikRdNKg0frAOavWUo1kmxkQPHo0He1J03hMbhybvplVfpojInyyEkmv0GE7D
XcWNHxqGlGfCbe2ihcuAmLLbxSXGnGB4Rl5RbyEekDcXrqgEaJ5ULXVZaIw9ZDAr
TbznvFQRtv3U0wqblFtJtY/TRCjxA9GDUIzfWM3qgkV0jMQ2l6oEufA1XNe2rCD9
rx4yM6OMuRw32SN56t8qOUz2DYBfDaLImFHMZnMl+nRUFinlogioUSLDmdcralnE
+tszHBQZvx0S6jUW9d44olSxOEVB5bsD4oJ/lhyRohal6+IwlqbjSBfSbXza030j
ocyuJBhIf+ZP/vkx3LWT0d5X4PPZOt3X+PJkjsw82bN2EdMkfAfIXt2bGdKqMFB8
5J9tl6TCt03Yo+6YB1vYzNYzeX41rX1bkJIT/mknscKgNvjbf6kCcgspfbBAX+i2
YRHSNvfYaEY8PyIHh3AnCTth3BPexxOHuwRehDKuKzACseNC9vhvldtsc6SZiJVp
Ye/o4aq7vCrf69sgpme8NybuE2LmtcaYnlxyhexWoVU0FTFm/Y0NQ4/FYdd70gRs
0bxiYwR5lAh/FYNGpCum+MO1PdOAuOHznwtjO3GVM5pz57Q3NHGdlhju0Gfv815K
bvd+0B2gUtx/fTQbC9pGlhDTsR2+4RKIxCoAPVfFDAnzIR2FrXzSEDLw9gFAks6T
/AZ3q1NgDjkoUkVpHryUkrYNrGDkzQsi3uuigJ+rkiEyfqlpq9ZlUqXfCOBhAjyY
s7qURGkO39luX6THLwrIEtcscDA+Ok1Nt1rqtN4cDXrrBomRsOmB5O3TZIbfWR7K
K9cH9EDSfwT928pWaZJUwDupfkYRGzsvzjQN4uxaOsSv+OrbqMPb0OE2FWdvaXc2
hbjDs/Ui6xr8SpN2VoFVj7INTHYCuiTM92nunjzL0IuMOy7075eIWctIjSRWR6vp
LXdVtQqkJPXlyh9uqcRXuWu9nDGAZohGqRUzsbhUj+/Yp4LiAVCK9w/akV0qTi/K
gZfgZWv5q8N/1T2G7QDa/+HuhjkU6FwBMmlWF+Ez3kV2AjsO/FLeE0sqRI++V4hI
PYoGY0J3PMeLIARA/RSc+k8LgGGfCk3o6/9lS4SDLRxWqSlrhbKXYpA4kMXOsWTu
B/mNXpv9HxLMsuly5VBZptgQEarCvjvsUM/xq+H3xuQCvVrNYAaXrPXoEahXiUHy
Jfg4XZx3PhTWsD3fIeUXkbWAc5z74K/N8JLb37cKv8+msmKzX5r+vQWXXP3ffDHV
XRjechQZVeXYhiv3joV2kUu/DRKGfNaulHH+MAhSSZU900pCtDrJiFN69/jAMqiz
+AyF4iX39zOfiJgcsQTXexhv69Gg5un1gw9mW1cJTuWM1rOHJf/ZdaLdJAYVrQv/
V2RxEgWT3UNmlu+HOpMlwnNYjgmrSjSLCK/0olMu+hOzOOh/mWyvRUiiRKChnu//
Qkmuc6ybXNB4ZWePgsRDHpg+ODaYwBDJIR23YtWqyP6rJS6qjIUVAI1Olu7GN9T8
CdFa8J08XtAxCEPy9l3DN3xRBe2TH8In4TSOqUBo448NldxySnyRn0j1Ekj4W65Z
rdL91BqNe2XWuayhCk7QbWEpB2Obp9LfpuRZ9WB2seAvjRE+lUHSurePb7Hm7YR5
8UhbRxw8KArLpHD5jGR/Tmgn7aeSORabcMn+a1r+z0fKj7hqGLqSYjapqdiNbOLo
570QqXERPl1Iurv/Q++UV3Y7uabrmyLG+LGcy4cBlwqeSHBKFktdAiIA47Mfm2WM
TrY2onx8NKbed1QiiJjIV7nNfqwiDC99n61z5SyW81rdjZh7l+TnZGfoyu9l1vec
v8zykbQfcZaUmnoe+L6B6x5nXnuzDybqcnfEuIGMMR9Q6ve9JAJ7ixo8AZ4qJNwo
n1ZS9y057MRpOGWpCoJxVjxzr6YnspBnfY+0OHkUV6xXPGIC5Zzy/85BvfXXqHN1
Pat+jfdXZrDhmHRGYK4wlbN70PHcBCWKybM1Qm4oJ/vTPlGSgcN9jZCRLmTHMciP
CwD6QxmDmSDX1DV7XfM3plL0Uavv4qHefSMomeesVxRw2WT+DSW8W6JU1mjxLCRQ
iqU2VHpJ/mMC/0lxG5WRb22Cvhv1LNFkg2g8J3WWwbUoeZ4hDQk7/YYcJNfyth4A
pHUgKgHMnbCZ5I+Myp9BnY2XDKzd9X/511JUFIOQTNYHarZg3RCv8u+Bz6A4GpnP
uDWHDim0xRuVvydAJfpZ5SUiJMdV55u2J01vP85Ai9HRZtvVCFgVJhMLw3gMIlY2
cQLwIc13i4YYCvf2xh9ePxUwFdhylF6oUlrZxLTXDRZrTAz8TzwCWEXY/PMG/xaB
bwpVOGDwk3+0XgNrqUlWu+m9Dzp4tUi9t5ubgtDSnzFTQ9G11aoj6eWfI1I9Ntaz
RqIFxKNcUWEbpLvfDUtuyrPYp6qH++KtfsutkJW6ibd0AD2bPfrl0AEmNno/5nx0
0F4sJ2R83M6eMAHLV4PA/ghG6RJE5P8UqjSmsnixGJrfAE8eDATyI/h4lGU7oK5c
okAF+cAxH6lqOtHCimpygCF+0EYEMeoeaET/6TNpQ7SFc78yP+Tk5Tmu6fsTS3zl
LYHVRHQLAWq48GMtyNjbc9HE2GbSuB1uNQQMtyw3mq5E6LQWHatSMwrNfSQIG+8D
QK7BL65kW+1o34d9kgOSw7zO4z/uBa6yIS/ZnEwrI6Nj4WXfmBn/A9st9ngDfoqs
aqEzksPlaipkWvyWghm2KQFCSpoP+t9pR749sDUz4gKV6cA0wvYKKYOSNaeT2xdr
Y3X286NCgkkc6oD4Bk+3AfwU1gPV1qwMhcO0bht0sljkzrIg9udD0KZVXpZSEp/6
UyYTP/FdQmy+E3lvVeskBuNukA3XYCpBrJjAtfxPsPMzo/F7eSouvCWXPYRqevPp
BxV/XRvxW77c2yuIWgAIsBRjxDSznCDPlUxFE3a9pLW8w7xqkaPUczV1IDnyyp1d
Vi7SZNftuGEFvCY+oLfXpjlqU8U/RbPrl6D28+LlJYc3yEOKGF/3mmjltaCiKTdc
qIR7Cc2Si2HN13RaslUACDRBdn+/cZnY1os36Y7IR2TsISm3nOnVDFOokGslUyBG
J4LC8Su+UwjdSM6H8FlSarLgDa7jEWdkVmsmiOXlC3PHrh6MI1Op6cNoED+AKBO6
1DduP2IaYT4BrBUqT7IBaVupyujxKRvT9xGtKijE+TFBPy8C4kFgdwWXeTlMT8p1
f4c8YPYcONwpLQ43QAi5eVPK5tbaVO62ooiYok1Czngo6X+TpGWBunTdFyAiY6ym
6bOAzVn3zKZqbD122yE9Eqx/IhSS+4M0nGGCD0oPC8gI1Q1L4Nz0IkXni0MaAjs/
bjGtpzfQN2btCBluOmfSImLJceHTlFcZVZW0lwgGwE9Lx5V89AbtaBmHi7BeQVOB
qLpUmxYW57P1u3TDIsuD9ciZUOaq1y8U6/o4Vi9QKsQwVfu3nHpFff19WWT8IJmt
19sVMRQxvisxebOJaND0yiynE9QVhZ/WG6rkV0dnSK9vqKAOa/oEj/2nG97wIFqV
rOW+0FnuvWVRBlJpWxmr6+wHpXzqBLokk4ZTEAxOJ3ncKz/Sw7BgdljWcMd/9Aqf
D4orSh+BfRZwTg148fd33ul2s3s6Q4lkiqyzLoR7h6lxyMVvT4C5nrAm6UZ38mBD
DN3LDIjLpsypAZDDrb0td++LggZQLu9Z/0Tx7WyqEu7fEc6NjW9pYtV85Cof5/bW
arCW10RDb8MKp2o1nO6SlTLUmk1WkDbjKpNusf1mo06W8QvQtngyZok3n8eQJKNH
62x1iI5WKTDayp8TtQ25QmxtmIdDzW5HOW8C7kRtLq3CL5PlGSXT/22rhpRpgtn+
QxUdcIpgyaaPOX+m7LwfXGQUNhm3yxMgZyLouolfMrR0I0iQ0b3N3oMnEm3T83AO
avrKQW5VAbX2VjzndTt7Hbjc7icstFZU0rzNmb7NT1Y6xRulFwc6uzFVFGUYVzR+
JhUFzbvrQ9e8JKNiM0x4p/lMzYjca3iAQCDQ1S3hjspB/f6lclXxvZ2w1TUD5xoa
3ZmSAeOg4zQC2FywD7+2Nv63LUY+pBO22gMSZ4qSpXikVBhJ8vkyQ2QS0ZOz0aWm
m+cbztjQiOKe1JGXzToMEtzMF7F36eWQAGuRGN5phTZzcnoO2U+aq3rg2AmdZU0M
J4UJ1LJqtep7edule7ZUpHLO3tVjNBaZK8S/KfW3eGJNyKMUaV7mmUzFMS5oVfA1
37XgJ9TyvNOb+2Pmf5Vm5hUlaJXCA7Xnq0l/ziJH6zWMu787Q/O63LW04qdz9L14
t1kqhhm8Pjp+ieJ/VkB8/Sb4v8QJ5lOq9Dn+OzB2SvIJUAEELKh8jFbUvjlvvDwN
paSobg7eMKZQ9h6NiJIjCymub1S34NxzcjANPKmLX9PIlif+HymNuC1I7pDQLtLG
AFcWEzmnAwG9bEGxCUw+5y1K+H1qlpA4Jj+ZG9qHjSpqMNtbImjJd86hb9ARzTF8
YCITII0dnNlqJPaJZqJxsFaSaMXvm6wpgj2ww/OGW/8=
`protect END_PROTECTED
