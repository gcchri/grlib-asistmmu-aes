`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RTxkgnjN8YGiesKcCniTYUf5JmLrDw6wKajYv4k5jnhqzI25ctRpqanKKTwrjsPT
MYQRcR3eGm7ga6Syq5mozajh9Pwp21Q8cn3aNugsBch7JCsV2kewP4pK1qaoQ6Ho
JJsjvF43LxdrTtN9Cqkz+VFndIDgwMEvuv8iwyXE0bkIr5/G3iT8b4j4YeEx3+aO
POMpEiOz/j6SDVXyRvXLahksVLP5k5o9LVeDgzjfIHvCb7yuN4SHr2/CcPFGANQH
LB/peGZU2d/Wi/yCRlgDyX5MSoZapHhUdbB/fk2Xdfiv8/gKOK3JtQHbq4BigjgY
91wt6KZ3+CL/yhGmZ1DPNA==
`protect END_PROTECTED
