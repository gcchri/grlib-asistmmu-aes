`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/wE8ADyvaqguZgPtwM6ix4gt2B4CazFb+XhdHkctRnltCqiWUuQKWAZ9GdKfvzda
63m25IJNNv6m7f04bCZuTdS2QrxB6kQlOOv4hCwkx0QgbJVVsfXr+AYbmItqdZML
PP3djUfXuRTVE6rsnZl17TuckF59aN5tJXysV+dIb2aSdcEG4a8ViDyfg27DySEE
9qOKa5Bn1riwXKQMG1Dwk4QMw6RSUMKMEsSAgP0ZQrEMqEL+sLt3wd7iRijJscy3
aPomzIshk9vc8zvOOQNVEeDNoqfbdT4SDtv264vBaNio16eOc1dM92I3fju+sMdN
zlpU2seQF+Oa/T5BqanbF2mWh57k8AO7vWgmMXLXRDyj3ndIWBoLQnic0OTw/C5+
ZaF5Qbm7th2U4urSRYYMrTbocpQnDeUR7zNy/LqcbQX+6I+q07B+VtFVUQoft9F8
5A/jO1xZO03lDKFJlPdHkb3fiQkyWaKpRYxHdowrT4dl+DYR1ruo+qwSTsyyAnwH
HCBiAHBjx2mmftibbv4J+BNCtLfkky0d/CvSmvvA0SBaIry8vWrrPnnyeCUBBKQh
HRalAT5muSu1U5RFlGgQhvUEmhMzzQAbuop2rXMJqEw=
`protect END_PROTECTED
