`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pjFAJfq6WgFcYmlHMaB+5SVZ5BRdfGh7IMTbkvPCJ4AY+fqLDpgLcInEuRfiR938
maC0mzRW7+Q+OEZTUx/4GxpPZgJhpoCyNcMG+l3e7M1UuSgduQ7uqDfmHjZq5+OX
wTSrUy4u8WaBqLPclZrD3EQlBM9jPXgzdqVWRp1gKBzirHrx9u2q1JRrKmvDEfyn
U1TSavg6HFICf1+qNkaZCXcAGkT2ivb165t66x0elbmPC6X0R9VVTgek5J+2zuzz
LpJ60fVOcSpvdISMVuEmmB7OhkAqhaCc5MFCax0hbWpMYEJfNxC1NtxBlpqofURa
3VIA1F53ogNjBSaYKPt3fFQgdIK+WE9lwczXpSglJsrdknS7cXj30m/HsJ+Vclos
zL+hg2oWUzmEGxyBb41hY+3nZ/nrwzZYRmN1tvrpXMI=
`protect END_PROTECTED
