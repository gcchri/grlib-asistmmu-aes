`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i0j74JYdXxXXck9ceEQlZ65RHUaW9RLz5d2dsydGMQcYsStCSC9vNL7z1eh1iaQv
spPva3/AMOCyV2z5P1Xi1GCMPkZVIKbC2bl1ZUb+Ay8kbPuep7jfywLNa5xrayhS
Q12sFrJXQ4wp8mZBrHLEMD0+mrgAxrw+d1fcKJpVpR8Bv8qFHQLL5TAswiNz3EGI
kYm5c1QdGdSEh2F5JTj9gjiBsr59/E5bFhcfxTC3n/d9aYloyWvaqY1NGm/j4Zt3
rwMW6JjqFIOiZ6rj0wyTYQ==
`protect END_PROTECTED
