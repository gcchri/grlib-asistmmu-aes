`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IDWyHVh1eGaFAT4ehFhx1MQCIaw5eKIG6uw5XlA6Jy9RlNLqBMLoLI2m2PzOiZZZ
27HjXuE6IHedWdxf/CFsK4tMYU4P+TX1iVz4PhjdErb68Kq3PlKua4R+dMK5/0cC
TKJke91/3msA6GpQEKBSAbRhvMZbarmdsdD5F1icmtTwrwQcZyUcorelspV4w//k
3dvtemP2bw80nKKzwbp3Cua4Enkawo4cG6RAeIA7fvRz0jRBTvwpE4ZuFZxr/16v
pfNL5I7+xnQgF9dolT870oxuOufMTJkyXd4RFo0Igt4H282WI+43ysQE310rHwbb
db5LTvbuLjUXvFBHdkuGQxqLl2+7VC10udfsA3PNxgALZv/pRBFgDwzVGLpS5ZYo
pyk3Kn5B3u7sYU0s/59AF7mZaIjPLsd0Km4aC0GiHvTntI3tdbYFVvF9eyNBLvrl
+y5CejB9//w//SQp1D2W90dMmfTuwsM22ZUbd69JkkoaMNuQc5JxwHvz+mA1zxvS
WPQkjBCQtXUMd+sp5Rf7SjFtUovi31auOa9ci60b7ZZz1Jq17wJAP5AQtdtgirjZ
Yy4xZbznORb0y+TXOYtVG1f7yZmwUwbpvZqwLWskfctMuFs6eqSDuPtzSM3WP2bu
o4nPGpqBX/OB9ofxSkRMQMNCwVvLGo03N6eEa6zI7O1W0VltHFwgUV37AtukC+88
3em6Gc8b4nffR0xuyyn69KrAUtKkHJ6TiW+yYG/d3KmGwSl0J73npJ8BEeRNnjat
Q+RsKFwVGqWW2V0zcytw6MXExwEKydbMvZ97f2O4DaGbYkAzMP7jujAeDW48+fyP
lvJGfzVlv1JUUAZ5VpXTDStDTHiSg2iw87MkB3b9n8Q+os0CCRmG4LC1eD53/Zrx
N5hl0IJJA9QQdeQpxkboMruxdgB9QZEUQZrTSSjI5A2X9nLkANVnGxrvDvIYP52L
`protect END_PROTECTED
