`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tsbv4rIhEoHYmjxna/9I54DMihCYI9Nb2Qd3Ib9O/o+nMEd/34BlsnzYlLZ3XVOv
VE+SWvCIDZ8opdY8j2FzxGlz7KORl+NhbGXKLa/CfnlA4Sgw8iNo2p97jvh3pcI+
Iu7hWMdErO5bGyYxJ0ODqgW5MhVN/dL5+NqEmTP1SWYoD7Ek2cZS/gkDWYwPSDYZ
yFQj+9sWU418u/3BfmLkx1FQVYp7zmJ9oDTSAkHQDbuGWnuSJf2Xa4CDv3bfJMQw
yF7rtQfR/Z1u+I8jaeVL979RJ8kYjRqu5BmdKbpwsbNG9YVFkmLWoMvuuVns1992
O6lZoyMQh59rotVEy7lKvg==
`protect END_PROTECTED
