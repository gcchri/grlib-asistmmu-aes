`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hb2dGQR2q3U6B4pcPhPFUNNzQJ5DkgdxEZdRo25joFFsOpLQ1tzk3nLmwXIxhFDw
xAGEp8TsPYCWxmuae/1tyR1y8OSao2R0R8CwaNWtl/h7WxygfL7hdUfSW/R1gN/6
AVZIEf/B5it7m2BqhzfU29cVl1Teww/DwlpVOH4btGrgc4GtalC1F//dnpU8VZiR
/UBN5F+zCufxQPEBeRkgvT4uLsRuIs11B0SNFJlcjPcK2mtybZirfYknFtZcyq1s
w6JBr00GXcvDZCC+wiVOHI2nxjUsf3ZH3dLRJOUMQhn6zcibtRDqat0pK6NjlXdv
gSeRrrCQ3Ussz8AMxww6NPYEZekWeVByekCOBCBaMqddephNGd7Cl4piaTEEdFAb
my9Pzas4Likfc3tJ5veGIA==
`protect END_PROTECTED
