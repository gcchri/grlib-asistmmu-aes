`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
35HlKwdx/6LrKUtWT6VWyfW/3ACrARuKlkZAmaued9nD/V2s+mbwZgbR3+fNGgnm
RyEtzilseWZ81ZkXCDDvHKujizcsmg2r+U7NT++djrj3c9oZEpQx75Sb/0Z7vRii
6sFYMEMybEgotgu8uPi8Beak305koE2R1xXYwSAyeI/FE6zt0mqdBqn5Y97uK1k8
A0yAGkd0kaot4l8NQnmoMcPqOkKAMDGFy0SFKj+7ZBFJJ7gTaLij/9h8MN9rNl6h
VNYvSo1JJ/w3kr7xIIFHtUUxkLF8Q3hiNhTxrzBYB9ac+nnEU9RS2L/oWqXGy6v2
qk5Ma9QSGFrIxUhXiLXEL4me45rYV1/AhBI+0hOglx96pw7J6zILGx3Piy9odUtj
BJ57+tjyjNFXyzZzYmMTMEUO99qkuGw30xgbBGsiu8LN3zKEDdAmLoLXP8aFvgeR
yEe5A8KV2funvR2eGKGLgxL6lz78OPsOj0zNmewfIvlukrAHxtlHw6YyvC8Pi0f2
thhcrwUvGtXGiFntjD9hmYgjHB+zcS6lVH7RDa4uFyjBs9/7cgdVcJ3gZaVg7/14
/JTrdWWzgl2Mi6Nnlr4dTLnH0AyOmNHKpqonZBBtR1p440rOk8dZShHEFzXArdfL
pXyG57ou3Al2vUAP/2r4cQ/RMso/G/rO4VZDiiplXzY/mW9MTL6N8ja3P+TzH9pM
eDNiBK65rLfi7i33YKNjpCYNAvD6oa6PSgn9t+yGwAAfOcK2Eqi5G8JtgXMh7Ggb
c8gRc+0pHiFbfavLC8S/PKH4BXmcLM2xRlGZ76J/wt/wRdDGdv2YixBEYoYx1BJZ
fheJOvUJG8r8d1nCTly0v/QmZNeYq1wTSmvSraIsUhyE6gAOKFLT8JVnoY7UM1/h
cqM2uaF6GvTToJcLgI8rMh7QzL8A8PAjPsj9GjWRT1oCBg2L7kSnQuWTrNTHgiFQ
Gji78aTXpMDgRrDISwuNsJJt6wrqTu3oLOd8BRXq1ChhpmNKPqJ3df7BJk8oNmOf
Afdc2hcKq0xXNxBP+At4Dprcq4bhvpnp7f3J2IpkrL+mNXeY5+S5XHVK63nZc6Na
y24r48FRxJ4Wy9qreNn31lx+rkvpRZcWUQclksfX3UYkcwPMWA4pSRpwOelmyw30
Omi/GeUnfiPboq5Ew0Gd3CPo577JhfX32vcqDSBayOVMvlzV3G3A5JLxO25/tkrp
PrhQSZ5Mx2pum/RZia9/AzcgAIc5HvPXBcGEszKmOU6LD1rN6jpKbG7ozTnWOyYN
11YhCMPCdUzplY43pnFhAdk7oR9PX30WUJGJC5lVVoLSFPzBJrKrJ2/C8AM3UUkA
MJxcEa2qdyEBI050Xcy/zcJjbCGfqAV2U9q8lT1Ot7xbKRP/eRLOFxcpK74sQCJc
GdgU0+cf6n5vv7VINJL0H8HslqBsoeADAo4dBc9Mk4a+k4KZOYuA4BZwhrDDcXGx
5UTq1KJ+OkNKxtu02htoD5jBvovtWfnTpcz8dfjfs1lZ6dyopo+45v2eX8CiAXBz
U07NJ99zVgOkmVwNvwSUuu5iiSDGt7GngrDdY4EC7dFwTBcKcvrk6IX3hzFPQXWJ
xwHoFneJaO0CODUPIPivUwIufV2b8xskrAdkn6LxgviU8/bgE71OQExVcCEOnSB6
+zR3vKxZic2CQ2D7qm0/A9C1rLJrGmN48njS9N16zjH1dcpkq6hjow7zzKz9SLsz
cCVLhI1kvLO3kg/HLV3wCoYGH5ECbG00imO6ZgpaiFijnB37ol5JYNHBw0R9AN0H
xaszMxg6KR+M/G6E2mNqQ7mrqb6ZxKp1469tPSwbsA0ZCTk85YzHZTraBhhszo/H
x3gGbNocoapRluPVE3cBG3tPeHwfpQ/o30xSkNQ5w45cBb4RhsuMbcjpYrcGal93
idPfrj/kQY/E4EfwcLtjAbhbGdOO2u6IQ81dRuz+5RATrQAnSEk5iHcBpEeeLr55
slAZnMl2Bz7OsBG5PmsOy3Q+MteaEq+6nLsoe/GOF/qL6h1/tbSUOl9cXMwDV726
22Bcm3jcTglCYab/aoLJp5xrQse9m8lpXp+FMILTmZLKgx4dUIAS5+cCKI/h6rrr
xHWxOGG/lEw7bFQEGWe4UQ==
`protect END_PROTECTED
