`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BTsQWjycFTA6inUZsBBeNDWPoISZSoz8h+X7LCoaHKdC/jaAfJk190ZvCDx9jWnh
/8XHiRk6/IowKSX0NQP4HxTxoBwwAPPJqnTFI011fnAR4SIC/dEg5LRCwtCnYI38
/upPuu7bTw2iEuPFQWulGvLxxfQjVTnH1shVTxtdlxlvuiqyAOPyPlpMsDojzXaA
ssMv0VXF88Tykre0rBzT+2OXjudrjfU7CPb6ZdExY7pmao7dr7eCW8/r+3PCQVnZ
vacX1SwOd7p1Cb+NyVaDs9KIq0PwymgW+W9GwzMlBnDUltzrgkAgfBNwMz4cKR03
mZi1xFtiLkWGNvlLkW+tJpTnCpgDmaFLFW1A5/6TLd2h/+Zr0FTKAkhHuzWldtCy
uAiU4O/uA7ncv6Il6V5tRr/hzRq1TtTlJXW4tELFs/OSjLz9lIsPyzAcCko26YGv
ZCaHBjOWBGakiYYZNbz8h3zo7RdV/vSlWKHTT3p1+9LNCPe++iOYXP5hyLcm2r4+
3AwAxQJZWWVOi+YcpOrpMnQNBxasM09rSxhVR2B/QFLFN10XGHmSve89/1RFfr3N
hyR5Q5IK7y9eq0kUZZPjHTruqRaSMSdViGIzIhmpWCA=
`protect END_PROTECTED
