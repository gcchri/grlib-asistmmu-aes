`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mZ3FORzcA8ogTPwIUlCsYks+4eB93P+f5hOBeYKO2KqOTPJb+SlnuWZcGcwIL4jw
2BgAuDnHumWGzauhyyGARSK4HoKLFX5nWs1PEn9GDXf8GAg3tO7lZZdBcnoIH4zs
ILdRWrrPXv2+MwKi9EX9688jdz1mkw06Lso9tQNgOUWRPxKi/3VCvMx8YEALGmXM
Mhr2Npr6BjD/xOmMOOAx0xNSOjccKi7GN+Ttwaz/rVMfV6zt4iZPallZynKnBiJN
lqtsHqne+B/YF+MYzx0D4o5a21AILt8RZDmUy4DJcx4bCkRXloI9U5LRGqTOAsza
jsCxjzB9xJL91DFKXtREaLK0loF//dicPtfds/E3RjX9GpU+YIMu7Vixb6M5xerM
qcS2rJFze0M/vM9DPRvgpxxTS9gBEsIlpddkHiNk0lQ=
`protect END_PROTECTED
