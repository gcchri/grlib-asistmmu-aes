`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dj7dQXtZ15U/wohkR9YFUTBgX4DmXyfk6CMN5y2rX6z6iikxrLzKSYWU5nGEX/mf
pF5VQZPRvlEIeb4L80JVPOwLt6x7zQorSidQD4mD0gmeSq34fgBMuodP753c7or7
nLFaKz5/zpxZi1gsYJBi404H2O5XG4FJEHuq98Q9jp0vbBzmI7JNRPKHQDbGnsHB
4SA+amxYmLIW08WtyVx+ycbQyB+IZLJ0CQO5J9xaK7v15qFwLKxs9SMy+sPejeHn
sOVAwNl9QZKrpm7nF5bwGZpV3jNMdAG5+zWV9s+T/YJXt11UK6jPGJeqIW8tISS0
Gumw5qinXa7byTn2/R+5OBMasgP9hQWzvUYyOiP5CL/DeMSgWaK8ZUOZM6AvGKim
JECrbxKf41NgKzDgCm5YnJDIwGjxr8/Si9dDaQC7PaQ=
`protect END_PROTECTED
