`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MzSJtNiBIi0zvqcSjMQICfGi6yBEbD/Q4h46CJsxWSWoRhrqLbEjoFpPdiP65sIe
kWPUUdHIO12ZIL2zbWW7/j5aDhEnl87PEY0Tk2wHmWIVvmauD9B2kIXTKLGQc9lQ
Orx4MkbXaM94V91MUAhe/Ecz7wVjKxACDLAASBq/RDymOwNNZN/rqdhbkEm3ZONL
6cWRNaa6NxycPkfGZlmIHnP5yQ6iAFX0zzehEzgt4DKJLW0tJaXASq5iA4KOAii9
2eObzLfqFT0NThjyOPbpnaEyZCgMDTqSRGIwXjAqFw/yNw+H7XKeEGoI9HJoHzcg
Zy0iXu7cZv93uo0V67YdeZddf4aJxwrf1c+1RGS6ujphnsHV6DFnK+7yzeUynDV+
vP1EcKV5ErTt9T68jcpy1zCvFuewrOTaCcALqKX1q/9W0VZvK7lMBnjq6VAZwvkW
Ufy4QYjq7X3b5zRF3PgcAhSQm2ojkm6TL9vvu4USzmXXlQa6ks8PTLcb1ghroTcF
dxsss/J2pU0zwavs8BT8gR89Na/zdDzrid4zeB7HDpX40kG818/rMQqnOIaP0n/u
QvF5RGo1SlPq+asfp9DHZ0yVu2CzC0TCeYo+JpnuE9grvg2FlzEjwQgbTLoTBeG+
`protect END_PROTECTED
