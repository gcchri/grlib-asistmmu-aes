`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XiNn3cH9WcvV6ImpZjnSFNFZXc/zMzlAwGlw+bfVaj7CLrQYyqL3F3eRG9LmNUXc
W5E06REyWznwDZqnwjSoGQ+mEB+jH97j2KSgbe/8mPH4DR1aDbxK6osRPnomDKI0
Da/ctoSVnFmwNjXBHsMkBY61YytuV+0DFnPjfn6rd1lGo6vF30WL/CyLkFAaeTbE
e8NEcxE/vEnhmiP+DzyVm2+BZSgB++aJWcwvl6HxIL+jjlvf1cWBeUGbLIIwfQjK
imONhOOxdpNU4a7ShGeOpTlQnILtOvopRVfftRPp5/8d9GnPjJFPFPPEqks/h9Dq
iNUYBKiACWW88rV7K3cSHRdKglDGq5Mv5O+xSVRRvnhORuGSwQ7VF1k40VLHTOcF
6yvFYkzKSxLYHfXcenCv6Bjy3vy5Hkm7gAL+shXRREJIyfj9jdvjsllBdot+HPNb
ujM40jyXo0RopRC8zKL7MyG8LhQbhia0zlJVyJNxvHHpyP3LMlVwfoZSyUHCRFjT
AWy5NEQBEs5QM4IY04ZiNEhAlxxJI4o/saDkSnk5gqnrzhm+N5x9fEPRP3WYsisK
BgitbznigrWlSkXUfxZbzR82MpWF4uDl+dkRcMPa0RbQi5ZqQq7WF5yytrz6aukH
sjU7lJEw1mr4QOBC7OTzHDAi0A4rqZOr1BznIm3mJNmPigbYX3jSGUjDqYlxKiBG
zNJ7ql/Ucoj4B/fQm+ZSEz6Do4XJNJdAYZaOD1Ex6oHZWPkmaUQYUMLZyMIqqcvK
PJ3hYE9blf2xxtcNrB89afmLKdoP4bA3fVQOeh9G0UgkL5scm6phjzml6oO4amFJ
8nlfz4/8poq/yEzLAihrpJ9p/EPGsmGozCTBWlev16BF4uG0b5uBL8rMxJ0v5O2J
oT3a4evyTtirsji10420db57bpR5UzWvCWWTxpybNCbgfMoYVcP/tbw8qcfklxp9
7jAgFLpNH1/eByyPd+EwQvvg2bt3UHvlFQ1gMoyF6dEHGGUD4cZUq66AM2nHLDqT
RQZaT16fqgJCPq4ltS3iRAFJifJKV5b7MwyLUKDB/4xeV9kK0Z/9tPgTmchmlPVV
9iPa3niR/4XQ3TFNHzZ0BGesewzBAKCZaMcQSYiILoK/ERKSHEFJw9gqpokHA+wA
CS+ZkiVEvn9soU0ge/GtwbxYJbVtnPQd5iRyQAiHGg66zuGP0ZQAFXVKNB0h7Cy7
C71X/j7jxS6sbYFKQ3uSkq3cbEM7nr7q9zFRkL9+I9OLE7PXFclXTj19Kj4ifW7k
0GQNOAWvD3K1mPBnQ37h/PwlAXMBOa1684tGcE2xCHhVVMK3IM6aVI3hh3teaMtk
d5ZA6xb6w7HlZ6kXwADGjQfKFqNcCpOGjZqwHw0JkwJT3to184kg7z3JLei323AG
lEGJUar1olKQdhjGDg/Ma79KyLnbjtr4RxAQEPPKZ7q8t4lYBlFnPe3c86ixQddM
6rIO8eNFaxw/8zdXuEDAi51Oe/Ln42qvkGbkNHxVGD55xZO0a9VjSmA3XBIv8raj
5diYM1IQ3uhZUwklRcebOjNhG5S0nq93q59f43eI6ZQXWyT/1E6YqU0CRmiEZYu6
QOksKtQVYMgcOpk1JyauV01IQj5XQRNlqLyJC2aMJCs8yC1U4tD7ZLc1dWcshODK
a0gVANfXw1PkwA+kEUkGydHywyYWXW2zH43wRzpX9/20u7tsVHxFOkwTZ/gke1LS
jAq7YWmv/MNsA7JmMbcrhomjKRmRl2SFm9aU+bXWGKZq8NEJjtcrvl8zyyTo5yip
GbYfQfsWUHwNcSt1atmy7gKQrxLO+5CgNesu1fTlUkK744pfBexJ8gtt04bC8eDl
V/oaWLh91TLlwqVutiwYvtRi5EqwUPlZ33kCqvwo9R4QbkEw/0z+/eTd5neYIoBH
`protect END_PROTECTED
