`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qqOL0mL6u2dRVZXMIQv05PMVgpzicj7CKzfdODrNwZ0inWH4H2lWy4eawWqjVxSx
wcb2JYmR5QcWdy3jv2/oEViKe+1aXdJgNamWBk/uI8uvzgspvVzHxrnPAZ0EuUkn
AHIpedWs3CtIV7Foh3m+wXTZI0HTYqOz5gatoVSRVit6lm5IYfVADg91S0ntg+XF
hHtKLIrA6jUDujGhRp7OJmEO9gGdjpi4k5olAf0JcSatgxNfxXbSvL3D6Ib2/WMf
vhZqdxiOevi1+lp4Og49ur9qkgOvU5C021kcKlYyU9NV21JLyenEnZKADWpjU+oX
PpIjIOjP7rE65pR8bK8DmfMvtLIpZGny3fsXWjPIZPgNmK8PLAjjPhWpemT1WFae
fHWva3vIslIgMegs4MnyIpYFXSJf4vsmJKfH/vZjQ2hGYOk5w0xitrkJzr+3IYO8
fm9VhXjlEB3aGtVXFgh6MIItXOMFYFc6UoA7jMo/0W7O1NSv9h6eBe1hvZCqPKCC
Ks6PYuhJaCjO81r8dfUwlp1lLF8564/SEu1kw3ivYF6xDaNg6vMt3lft03ydIHhS
hQLUfcqrTEVOApmeZbbFPQs8yGW2SYZFXGhtKOLScd0Q6RkLmnZJPWpJJTmYdRgb
d5Ma9m805E+WPdgRox6r5CVNSFY40/KxcKl9GoU0UwmdYRbZKvGw2PHfUb9cIK5o
xWNKdpGgyOZEAr4xyn7KLrofXMumu2F4igSL1gcYh5Fa9ILnDAqtQVBLGwZ40rtP
ZO4jQWF+J0vemTX0w05to5ceBoWDfJAs0+5DOMPNJuco9jfGTVuB25e6esuROZ3e
hROBNZ2r7tmmWgfDYkKaBlvcZvoMR3uzD/YE/I+wLQigde2f2P7cF8e5HRGBbfBL
iNQl9ZVRDFMhCBjZ7aTqUIfd6e7xeK6tCYCdu6WVJzMYSQbTTfSiod6d6DZ6vMbF
I33mUhg4OIz/6tRPtNtNPFQqnrNMZtq4pghXYyYv5HDs3K51RO/LK+O8kz+QFMuN
gyf82QVS4fX0+Cq1a5WJhUpI6M94Hbbv4so8JEj8XK6BJOAPQh9G/IqffyyUbKRn
fOHScphcAKRJ9itSGsnpwZwvImBxXWkQ/lbwSe73uql4nuuDxfAq0GIpXxmIJsvl
HMy7Qf62u3eZkA6YMMvI8vaIv5gYxFZmtmCatQHPIGoalSKhpMy2qBHiuJlEoUAF
aCX8XXDwr/VE3YFdtEYgfUs2fpOmThKeM+yZJ2tK2iDMcRG2WccL5rsrK4x7d2jW
2wwI0NnYF9Deu4kFLmGOBY/kASc1lCiP3hrLpi9bjRPEGKKZDXDNcDmpcSeFxJuz
jHs/tPP3wymqSzq9qgLJ9GseoDas72zfisalzUG/Ide9nQ0QkYTZUecJ5S09Hubk
689vn+HXn7/I1KYXurBjUeHqEBXpMfoOuuoWT/GEtQTOjoRp1vVD15u0WBZwFADs
fG5laQfZbwiPoD3OWQCXVkm2+QQdSelRWAK0DV5IKv1Dn9py6yZ9D5NmAk7PBKxh
ZYrGL8ahdCnaat5b4NUXJtJElVq5e6MOzncMKZ8SghuZ1yErm36daup4StenqNER
8W0Pe6iqFVqDflcrVNLMyijPndKPEYJ+iTnDTk2R1NVCuzR4zuFNsXDL3jOEss6H
oflbcGuDgEfzklDkA8COew==
`protect END_PROTECTED
