`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4xSLszBuagT6zDWnZ+tUOiuA+IAexWXx3JUuLrcXQ4nJzQlrfkWKQqQxOHXi7iGy
gFDqGe+Fk5m1cd5ncy4P1u71+Pwwvn0QAEicmLUHs3LNKMgQ4SIYIjGu4PT777Mk
ctCNMTnX3nnXeMy+NN/hNQjvRaGFjKIi3sXkk1mXz9DugRDvxdfHbsCwxTMj7kvr
DOg0t7aqPYsSC2ZG3tObsni194i38FwHCzn+LthIPL1rgf4gnxkOOKdEU6kKX105
Hn/Qg0X/sktdakFv45eahcjjOo6gG97O0Efzt0GhxGbvbwmCsK/bmT17rTUy8o7j
IAT4KJKC9fJ5FpupBSc61LxgywPVViXfchuwEcceHqSQrQg6KPT1veNUrdTCikFz
p04TVqQByV8BB0JbIq/CzlJsWW5Hao8YzJQrwWeWvHE2LrPjrb8cDsHu0eIzDwvE
UvYWyo8VUoIQHTAUVVeehGkEM2iDTJpTVHMNmStm71H060LbKaYKRlPHcGv/nCYh
lHHI4lS8Eb15zYSPAaChPjNUKbDoWiSyK9GAoap0ZOWvIicoaR1RUKXtzctsJ3QY
aXojXHKFbyGNlkX2kDc57bhn1MOCPjSfU1DsXfweT7YFGqHYD/TN3yCToAHaETcP
ThdU37lRB7j+EYiguSeGmIzVhzpMwKmjPNqyvI8XE5VKY0qv02VwWUQ7urkiQqNz
dCMUhgAZWeiXMbFR9lMuc+Pjh2rMC6VpN4hnGrx/a38zoBVkH66uCF/GqEwkkPE2
4wLIOZuxm+odYuN8FBr4oIf1Qi3+vbaT9NRyAJgknV0qmpHBJ8egeQpuxPs65uTQ
Htzcvb6jjXy4YIRqOB85x9g1NvBLTrBJLE4XS6TRlnU9Z6chaBMJX1BwEwqg17so
yn7f8yoXVzjI6jMc/NgYWy7vCWIO5tfedpJ+kSaDY1LTVX0S0lWnu4wLkP5vecrQ
/EUCqBzwjbzPwIHHEt92NoXDe8EWO0gxeZ8MpQO8QtRZd/Zf9XY39eR/SikAILPj
GcTnyYufowKOU6M3CaejMxmRfjqck/v9S0SmoRzgBokiRKgnE6pIyJnzVY62ZmGm
BnIoV0THHMelLEqfVBRNQ0tfooO9mEVJqnRHbCKzsD/P8444DB1o+yBTqWO9/30n
1htNfFopaH0pykYz5bfvlaKG313ubSEhJlZ/nrhXQ/N0YMtyxl4SjOMdz8HB/35f
oiRqwV8oSzwolzgqj8ZoJFOTwt7yUyekUTgqIIpibVSXgUZb9xgmFN8rSOtUYk7S
zDsQ4ulNUDcl0JFhpC0XC/ums0ojWs627zB0fKix7TrN3lcR2A0IGmRLNB2rufjL
9MoZpejt0USx5MZld0xV27kAB2R17xAmF+DUKYo8lcJ2u4wEWG6aRQZxeBkHQWyV
3UIdwSKi8vdZKW9UX7vdQiFDozxfwdslOJI51gSe57t7BePxQL4BwarFh6eAqfvD
33nHgXAMPvAU7KyCLUUfDsLJLPPog4n8Q9qHWFtwGxxQBR00dXyoFvMzRF3XRrJU
kHNmNPH7yPMhjQThlBrVuK9acjvQdQYSVzFWDkezHwYDdHXo+3AI6QRuEw9Pz7BB
wSP2Pr5KGSZ+jgYTO8FZaXk7FCKkP/WjXY9njcgw4Sp6fKj0NVI/MuX3+p7IcUnf
+qm8Dc/JzNSlbJ4J+thEZZRRVrQkg3mn9/8Lia/K7qxF5A3eS2HsKWFXh9koVqpt
yecn6Hu/0CawplKRqTe0Zrn4i72K7FEtX5YO06xMEp0VzSnuISvlUNLa3rZgUNep
V0K1hwG7GHBiCTlbiD26TfME8NYYd6wXdA9LELuzupVqKnYgYbBzcH8gdrhnBR2W
bp9qi8T/fp8Jds5GjaWSJFbPmxVZdmrBZnq9Ylhi/1MGzjyYwhmKfmeQ32IeyxpI
jBBRPJLHoCTPVLnYC4XnRBU3o6hkNhi3Y5nbwXH8kc8TeUfN1y3fcm67hXRMCG3p
DaFOgLDVawkIliUt8tY3UyN7aPXA5WsfWocoW0jgW72gGTXN6ziooa/A34XyYQIn
bie6iGG2cUQyHp6b8zUXaXNcBoonq3r/MuFhKAV0i+/pPVo08kX7+dqmF5AZ+tkL
SQP0naNnERHxedtVty8GhIveDYDXuKnyum41lrrdTQiami1FEnMEc9cv8Xh1C0ux
DEqiJXXqwPg5yk+rpgoRcul2mmOgm+fr1Bvcd0RfVpDmCE1GZwsa9S9NXG8AId4Z
3W3GxFsraFyPf5Mieg174AlWfHSLU2lO8GmrV3fokNPKoKvGvUoMvJASDOH1zmZS
D8NkCoZAhj1cvG2uMm9vhPaC89N7x4dar7AD0rNzQ6ElX/6PBbsHzWvI2cz+fYAI
jJ6sRXrYP8CIRXLcS05DZnMVs8vI1BxbSvSyAlnr1MNHBJdNFye3GUQYfo9PxzCD
MI3R6DGCMI6c5SdcAel+7qy2XBV12fx8Or0OCCjWd2HWZqb8IqZUxIjgmk3lt1Py
1rs2uw5PAhmY8IZjbL/uEKlJm8XlQOv/1Bs1OaPog/sJM2OU5lU45ew0WWqp3skx
FOOfhcEs38I3ByKeZeDooqMPCBwPqooU3ZpFmpBx47t8Iv2c3VpD2Xl36pn7Kx3D
cmQOfqULaPBEhK6RAnfL3CzNbYLZwrP41yjZpJDmfQquNj7bpGYeZeyglj7JShi1
yyzUBmaeawme+o/fhJxoIsZaEME3vm9tTLw2oCKiwTO1u/td5ec4c0B/0E4qklwl
4/LtOfOYc7gwJvRjkwsolBJwK2acCTd5y57sa0yiWedQeXm0QTbi2iHQcwPKdk6C
MhbB5GtAj7svm32iMnicgg1yJR4aG9+Axev9I5JbzPAwlyfYXIlM4WhnWKv/JtAm
tUIh33K4pwLT+sJiaV5j1WaEzWeu0B8oUPrG5BqsxZa0958UZRx2idYphRZhCo16
ZiVODigJ6jROP1AR/yKw1sHGmMNs3r/QHlYMVNA5fWbSQeGIWNKdhcviTiIj3ZlC
8pK1Iuod38qO/UJyolBjqYdf0RvlWaV3DPWzCfcR9vETudEJKS+Ume3iTF+MtYLz
L+YDkPy0oOc4R3b9PPtIFcsDeoUoisk7eITSoFupVc4rzZtHSoKlSWN4etl9FuTs
mgU3j94bOTWB9+UZdcxHZYmj//niJNsPX/2JCQYpqjQKD6t6o8ilqBaAK3xz4obP
KjAEjxq15fwRThYPZBu6XX4KwHFK9hE7TkKNsE93+hiz/mLKkYS0Qq90inApSihi
v1Gd9Np1AxQJBwM5sOhC8h4cCDFWJFNnbjBN+Iv1uMGBtvlBP2jVOj5ckPvWdTMO
kzwdmEBB+G9SMymX3Mx5OGZYqq+VwXT+WKNEWCWvDIHivpvwFej1E39j8ZyTFR6o
jKE5EdE8jOivUS8RCk/ROBUnAQNnA46LCX1eSAIHXkLQeRoih2ntC0yO6sjjsULF
W6ooltBdTNduHOw/7kKpWRCgFyiLuFuHja3+II/8y/HmWB80U+XibyEOkEYtkeTZ
HZDq1ItzFuyntq8Nhsbxx3eUAoPjQzFzJaN5qEf+3YaBjdPQJ65rOc/Be72coL6l
FJL6Yff9ownt8ldrijidW3IYt3Om89SKVTpaoTbZ3s19qTuhU7YZzsWwTPbH39+c
ThSbT4Nxc8UznVCRH53rIyFHrznO/bYjjtyyN/cH4G8cPaNji2iRClXdGDMvc2Xs
hoYyAmkTebwEq/B/KBaKPA3ZeXQ7f8MfaSDRWANRWDFeT4PMtypTIb2vfXswow2l
oNuyFCCnpYAeybLXansVtiQk3c1DI2vkUfsMyTeUM7EWs5V7rSAk2CxKo/o4Xn+q
5FPM/EnztyyVAwGFiDB9tcmgwITcmZsfhpeCFE2+g6zXZBWJgImcvqaDu/UWeP4z
J4sQTyY3IEGXWz4yyfOZE2Z1nb2t6RmTtRbZdVP/3YtkJ+HNzdNVHz8S2Z/dhGkP
XQWd5IUe/ZtyZQy8GuHnF9060BkeGFJof2r8hef5elhth90tETSe7t/9bxPTjd65
P80WiNXL6FSw5vlPsKuFD/2Oq6Edvfmp/fi9uj+PEjgyywoCsDwtDoOojNsee0Uj
wXZVgkfd5mxAGJSeisC10VkMVlUJmtLpmLi8flw2yPIrKslYtolc17DsUW61nnNk
OceYcyfZVlZD1IwTPwGIuiiQUW9/+jG/Lj9U6KBgirC90QpgLKESICDwAKODNtTV
DypH3v162mKzidaqndFlyvNrE66ueonZQ/RnaDnhkwJep8w/47CYQpsBh+TnmMTF
N6uy86uYJV9aWjQIEQsQO8BwnWJNamoI5CpXV3EHVPGhdmLh+uBl3u11sikZW3Ru
DpXyt32UYFpIjsy89xeMD4g70MjTfhwE9JsJYcvnHCTCW0lYxsVfjfUpG6zcNt67
eF2zY+gFViovxOyM0fg9DL5TLsdQK0kl8U/wTLilWBRfw/EhwCWEe755l4HxPvBp
+tk+j5vYAouCz9spQpAUqdN/xm0z9EcZJ8pTTZN+gYTezTVQqwuAr20QDISh3xmi
hLrGG/flfui3D/4atKskRfREt6+ojJGoqsjlk8XOJvDixVllkUAkbWKT6hK/0keS
8CxDLY2X+VLJFp0L6DRQDGwsQBZXAvn1j2XjxyJrRld5hwcLxQp3iGGzW+J7aEQ+
iL3Tgd7Lo4t7R2yyQRtLyUiYJlVJikFQiLsp1EnZxrAvBcxGPfIdXA5JAN2GU7eb
Q+uIR/6CwICDGXglQouesH39r/MKIX5csvwbCFX23/VGJQRCRVJDiXAQ+KgrQHRW
N0j/ud3svtepcwPTPFtg6nrw204XqzKsz3AX15cgyD/W7q8wKEUbqzL1SPe9rnoH
fcuqct6T5Q2nB0LHZaOAhsodCC83yho+fJBawx/p4GfV3EYb9QwrUsUnKypm0bwY
pGskcQsBi4hSg5COBQV9nSg1BKUBMXPdq9TgCOV4C2KyIo/c6L8c2fR9sLm6OT+c
luDtpr2cFzQAItC/P6eqTJ8UCYx6fGejXRWfq3nJ9CRNwh1QISIg6BY2L0lhy34C
eycrkfaXiV4c7zLg6QFyXP1WNwsplohyjfMf6xR+T36yUM2tkR5a6QNQH+ITuMdB
spegf7UN7IWJjulbIGu63Sz4anm9QOl0z3WJhSx8cYpnH1oQF021cTStTsjY0u2D
a3tj+WnapRt/P5tU6YETrSq21IXksNKYaQl1lTDHCPmu2loJS4kPOS2P9lo67R0K
VZEAR1/PBPh5LowefH4IOT6EH0YxuMCi8AzU7E84vyCc/6C0WTdmfsfsXpC8Sneq
ZCh1rFF99YAD9dfDgF8tzu3TtWb32BBxenr15oCtWVwUha3zt3LblOlabFCNO1n0
lh+iaw5P3+xoDdX7AzeTZsPvnwHAxGgxHl2gkbQSBMw4ckmg8xQqEkPP3vAOBUW6
rUbjsx+zlCnhfyrPpuC7vtNDSdwK5zViO/yqwluB8XvkQMFfnKtPbZt/9mBi7qL4
UfpE70CHdcuozbpfXMJfB+XAWk2d33zNNZa2w8Rz8/X/YquEipZUtjjjpSSb7GpC
/EIfo3s5stJkqgTba0acThSdZfJNlgFqIoA8Xjb7quiHk7540pSTfIWP4J3tfV/o
79ItXPagGn6Ll0iu/3pjIM2sDnHozulpzKrhJ4FlZl9tKKlyHkdl4isMygadq3Jf
L2wVaV2OstRCAuY8/KL80kXRmCFNnZhdaq3kLsIMp9rWR2axPahtlEL6i9tDJ3Rq
iPZasNSSQjHzQxunAPqa25fJn5YEb0R/dZK8psiAHJSfUDbkGvnlzBUnWbm/GqoG
wCskg59WSgzdhgzsGKkdUVuPlvBhElVRwl1d4t33r1bkj12e2PQmvNq6+5myNQJT
RyZorAhOFwwmtXIIA8EJio+7Bvov5A00ekwnefrhI86HFzQWyJMkFwinHjz+XbW+
fN/uRMQ/p5XNBQ08GQMlMQsZrOZE8eziVQGKH6Tdfyl7zRPHiSvMcPnZwzFOrVaj
5RXHyMrsp6R3qea4W0MyYbxTwGY7koxhp9F13a7LoXzryYsW1/vFv0hN1bth3cdi
g8JTyoM9NqqrPewP98aW0sRea2jN/8RNtH2jzZSfbSvsYjNxxg8dDfVyrS9+2u/g
pEFZMKg8J1Q8eQpZdexQKKh0ymsieKUHbQr9sEhausX36N6r0N4F8c6aE8LDCxVy
tBDacyYXCzF3V8xLOj0vPHX+CnlI+Fwq3TfBkIveF5AeaacIFnlz8Qy+tgH+XDCq
uRwaX+58iyzb4WwbU7BcqJTIwUKkZ+7botwoExjMTGgr12le29Zzgs20DJBdJ0b7
AhUA1IrUW6L6KcpqCg4AzbkfPJka49CmBjjWvvQVZ/1IzjIDGs+CPs8HYsDoHZFr
oMzvHg/7xxDr1Wue3Z6iwHTDltSdkGvGNDLJwchP7FT+hLIyayqxbtg2fJLBx47P
ozdNkuE8DYYhL593po0r/hpRdS2U9t9Gb51b5rf22q2Z+sO4cGpXq/oNfr0KtIWm
+4vQW2AISY47nUVfpBHVA9bLYHDgiEA15CsbDB2EeNr1VilmyMyFA5ACN3p1qR+r
2kqRGMAbxLBJmL3C1shd2CkpEofA7SXhpgUPQ/1TCqQYgJ5ATXS+MKt1INcyGXGF
Ie/7H+NKQ/YRBDjrtx8fIcUzEaoAMz/r8Ulh6fgDAnvYE8K0QDAktgyqL7VJe99D
N9WqtG+1J6mscF0MtkY6mLhUtFmzuX3RsOBbLeI2RKe14B5l8OICB4x3wpbeaNul
kQ0E3mz6xnTBurUlpb0OBbnxRbp61oy/+OH+LIOPqTwot7kA534s/C67xplUmdVV
GOlJFyo0RLKEa1hUwdjC0uKkCxH0SN6QP0F7J+nfvrht4lAxt8kWdYINodsnfe6X
/xAlPGK8DzQZ9ko682LGIzmP0FfKFUeL8+GPH4GUKGaB1yH+LCe1BYBxblTqngGl
Y4K/lJInoB0USGalMTuKCppIlLmjLGkXyK4GH9rs+kblPCLNF4ZpxMVEdhpUHa3V
bg6cIyJ61wBejl/P/gsqqD5hsTjQg6oBedIBv97UwqDT83pSb6V9FJ2e/4IcAsSV
pBXlBDHWsyxDlEmPYk/UQNq5hFCnZ0tvf9HGfxJlRXXbCgiK13BdansWNj/6nxzW
WIxfjXzxm8OlSyw4GnMzFf9441Jt/0hu3xbUyI9lo9Bah5/NAqwk4OHy8gezYA6C
5ZVFyspINRPGoOmqSCqBWWt5mdA+Ap5xWXcZmdLqBrgwGvYhKVq2TmzPslVPnBwr
ZzJhiUNd1S9EK4fenCC6VmyQuzWD87LF6Zw3QZXbu/psNc9ji4rZnj9rgr5hFODk
pV268TkTdMvTRTskVi/hd26z3Mc6rBcpMBSj5f1BV3VoOqbIfXVdqYsBomwjrtPt
2sPlbSjxNeCL+PQ8I6BR74EAipFcIorzfxbOhRGb+A3TAx3bDA3mGc4y8NA9pq5L
ocwDB0mcWD0V3TKxfn203Ww4YGjzDvqB3OKMHBmJftGapDIVLonkiJ2Vx30x9zAB
RoWbZNtTuFVy1v+AVOs51tcsmQ6JOH62o3RM6gQJmGuI07Wy3jCAU5ha0y0YqZ5a
rIfGJjzijHfMOoUTUAeV7Qz7G4tRVgcBrJiMcygGJgyEIb5G+sBvJL197lXhNO8Q
r2ezThIhWi4AMrMd3bRbRkeQ0pdEqQfPjOXwPVAO5KmepzfscVN/9Uxcuqudct9W
fOvFN0tWZcyVSNM5c8KFIK/+fqSu5ArFHi1G8dNeaWE69pfL1VxjZMVb2G4Td0zS
Ef0pL8SFQ8F0Y069nGEQE6XeIiKM4BotU5XosFsudFUrlTbKzJQUrPoWv+Bpllw0
+JVbsRNQbTB0OkiFr6t/eGjGJ/alONptCrVv5e7Zxcq30wu6VHnfs0olhmgiZ7dk
Yvuq1YwiSZKWyefkHaWNAO6N9MzThTBI0/nc0Qfsub5NWWPZlwv6MvRDB/zVGH+6
QSbug0JJ8F08mTx0wS0qNhMrA3fOyslbv0dmkpw6uFGIF+Dgn9wmrqDWamDE0SZi
ODSwMEpNKh4n7+nsh8KrG0KlZBA8G+yvN2eo9KLNUoni42VnQgf840TFQVMRGM++
uYUgTnrS0T8/3uBxGZOZRlMaXTGP+3YyFwvWeuE6ZcKWWsdipQjShfL/WDoiEufJ
pWU7uyUYwb3T2cU0Fr4AX17wLcDtgIovzJfrwFVlRWcDz80THvHj3N/Dbddzrb/v
dYoOMjOywD6lRuG5OYNxRtWK+GPuSuWCQ5hp1DZh8Dsw75FDvDDEGkJ1qbDH1+hZ
6FZeqhmOAMoOuUzrJ5GiR/0SWx1wLtOMh0qB6r6AU0WjQavD780wtqT5ELvCP4Q4
FlfoyqXPgoEoJKx6JtX7MnRpw6zf5dSvAgKPAi57gqK2UZtNGWdUQt22T6dcqFEG
EBcqQuY0ldgw/M0P9FWy1poJ07Ny9vZA9uIi32N0gHjYWpjU4qv60ukW8FN5klFj
LysZNFz/fZlkzfpraBqC7NQGVxDYXfGuL46ymqrNvRBN6PK8C5b/B1MJVMpfXcCg
HtrhVBYSfL2MN5gwV/f/FdK2PGWews3mRe0gjHsmYv0vucn56ICJT8Yvsmph8HP6
fFISSwZkm/uYc7ftT9h3wNR9oaBz+dy+Iw/SWYd/laHE8SVIdTxDnGtxkpJ0SVge
fh5C2kHk8sioOo57G9HNkVWlGNeqpVNKaP8CAJG6reZ0RLiQQhT4gNkPyYK/JcQK
0/r+6DjHzFifVaGyQ0f7hKqweN2m1TYKKWAqY79mNZMI2mecMune09hEi0Yhlmsr
f6Ql9twwVt35pVZjkjlEhNLvCYrxL2pL4+5mSKH0DNz/bavIPcQaK0W6H/+0CHG+
PRXhpM1A03YVAhzGDq4O+7fLBgRhAPb/3qaltNpah99xBTM7STHo6OllM12JtJsC
0/+4O/qiECTVg8DQbhAOAVxKjGXhzWjIcDTUSXUOnhrgErcHM+uCbY6buHrAATZ7
QlJN40hZeuo0iFTFqMA3AmBl9OhT8DFHdV9WWVcd8Xf5n3pqJJHwWEkgwzetmfdJ
Tn4a9t/g0fOHycn4Sx/XvQATUEumxruk7Q1FjDx+E2BQIiruUygf974/b8hEeUzT
Kp7VhTa3UMLthztquAFSYUdIJW3O8jhf+C6gezfWC/n80lqYxrWyGE+DeolwGvjA
WhFDBpgngNF5DE1vxfgZFVW6vqmUoxvKdv3hjayvZKaaRJbNeg6zF3N248vzetJJ
WUB14Zt6MR1VdZrwqM44/7QY0gPtoH0wMpBRA3GUaLlsgJxKoEi9AvXWeeM9K52X
zJs8oq7EXC//7xV1KR9vnYHckvCj/6OAT2uI8K4Z8tgKwFj2JE4iItPV31zuSYQi
KvBUOpQFw9njloVOp22cudzJY34/nBR7LSblh6ArM6sA6S75CQ0H0w2/98MH7/m4
D9lV6ggL6XYY3E4hbLnSDaq5+g9qofEoWOjUvMf5KdhZviJgN/S8e/b71+jR0tya
/mDqIymSZjP5y0MG+E/vhTOYdbxqM2ZaUc2tONeucxx8eQjJztpf5LHbHp7NBW/X
HkUcmvQV0jKRRyJmbVciRJ2qA3XllmHMwWBDnZKxjeiwPsvX7lKdZft6xQk7MARx
nX2MkQirIvQ9NnVsnA+qfw83ira9NzUWZzM8zEC8vrDtqmYGfVBA5YPfFL7cFsF3
iSjUFjZiF7nkq9X9TUeisgB7J8gl7Z5C9gf17rCnOZWcV+M9zthrtxHeHtta0hVY
cqn3akSkUAFz8yHAOmrlo1d/D7ERzrsowrOmt0O5aJNpgW7eSGFnMHS54pGzkIMc
TO/IjqUTcC7rTl7jymIT4NUKoGWPiorOkn1Z6MlfYBEfVy+WtBfEAOSa0p9HxFV4
T4jW2Nj8h99F4WeONKEWLoaYKTH3lNu+pI/AHTx+kLuNU3Ee9BjRccTXESJxW0ou
P25wHxnjmEwJC/DwYOUlPKAklplGdLs7oLKyKy1jfo0A/cDLRfg4M3YYNI3E30lG
SAwqYk2VBMXvltqAoUBPFq/nZGDGkLtnfYEOVFjcysiEos5DbvpkSjfNPCrfXBjf
DGmCjrQwn8xFGbo1nV0JUAh2t8wpgEphlECZtRgqXq8sG00zHAiExrl68miC9GB4
uGx4HWFTxQcOPaG/yiVsg+BWw2J7/OQ7ag+e2uxR+6TZGYKMqMwr3i62OEU2SFjS
bkIVgn0/zKy/6Uy/AyAdMdNdgmQ8nUsJhxiUqbAENkhEoWi6dZSIlHxOQnK1QNWm
q+LLUvQnCgWnYLcEcOSV5oju5Q2gzl03uOMRJJTET0eF3QCvJjsNRJZF4G3xJEZR
AI5aZn3dSTewcMI9+kvsEZnOOzUK0c4BoIno03XqW5+KPSWrs0Djir8IOdgPRXrS
8lJSHgwyYld1f9cFqmr6f1Oy71j4zRzPDog6bKs4JKxTSZon6d/uGyN4IHvxkCuh
nzJVrwDT5MbhWTLGtHQps4Zx0AOBtxh7OyCJJGhRghcEo4qn0e3UuaKyMaCcxIlF
nt17rY6A+bSFirOuiQiCFtgcEnjH6bZBdX5CqULcEkAvZ1lYCXQyZ86gxyGZaBEs
UcMsq3GK2Nkxkj2AnSsiuqnkqtXK0wXjxedTlsxBvhYDopa5h4OK2vykU5BQZnaU
iGFb1Ozp+mdiREnfJeG7tZqO/g6H/sSfFUGfbHH//1rcFpg3NToh3PxB8KWGL8GZ
mux4wGCCBIn5LlTG3tD/9p8WyWcqMmkkHs49mdtCavElvJDGJ1rIRTEJK0WNaNaC
+Y2RM+7YxvvP2OF6at0JA3eijrCNFYTrP03tyQegBvSFaplHNaRW7RvOeOLARGYB
aSk/xoMDdmvsk4aATR/tNmjmshoWypYOmq4K7oR9XICNuSWxmBSwD+X3KiTAv0DU
moAvDCRfkm8ciUWWgOT3pW+mjuowrUsr2tAALeXMb7fbdFgy9g+LeivMaNHlYTBc
TMJiRz7aV4HnafVUzAMH2votqMWJWg62BgtDyUMVa5kfu/kwGILKJQXOJDxpseLC
ZyXh5LCgr7zFwJEbQdE5h0zObYrAcgSFxal01y2cdiyEULWgksAPWICGI1gaDOVJ
Jvdy4b/GHc+fugyP8f9E3/E5KQUCYJayusxqMRLGbQeOHpC9KiM0IfDVT07IHuKJ
usGm2YbMfdBlbK1f1VbUgBPdUeuc3n/QY4W3BInF2qT4BF5nwC9W+/ONINh3upMX
UvrZ3EZLPN5DJhTczE8VrzLWbuQFkF+z/UsEjFBLSRIEuxpaS2aUUId73i/sqO+3
wpMqNe1DuLaX9zbdke1rZYePrSeCx0a3QCNw56XgLy8CSinuv2sER/K1YXAsOU/w
oQTME77l1EuHjBUM0IT5YNAC/g2cilyEaU7moRdlVko9loBkZOnT2B6mvSF849Qd
GxQ91vNasq5oZTgVakQEcRwwPajeOCL5bpa/t6ISCNLJgWC6UKvgp/g9LCbLVNuT
eiyeUGAaKz/hP9bicm+n64vX1sEws8rmjeWzqm75xQRiPbAN/dl3MR0POOopFNz4
vvLCtzoJJz5zgA7+SrWqpNYS1w/OmMGZjHV678g8wMMsxPBE0B9/TOqkZndLmAyc
nipasWJlvZTC1TdZRCUfG7zpneF9vHJCsVmLloZ8ULCOiczZVbmQxcG0N1DjCOE7
XVa8K1MQS6CvOyhRh7yKZGJWJmIt1eVrxGBQJeC8fHz2ZBXqA08/UkjONTKo2q+0
6awlmN7daJOf15tFtz1AhnkMKOYG/aU8kSYrTvM+HkIpIcprefNHecQfVxr6H68c
f+LLziyD+EI9vRwYqyKzkuWHBQPZxbQdSAAS9uJ2lhTFDJETNwjawoQVrYC/OWrF
K7swmHFfKCvgdXIlTP5R/OZITJGg3NwftEEoMowejwe4yXR9tcW+zW3TKvcGPAL9
/x/pNmjcdjMzLO2LjaDDDXZIQyi3ml+PVaUzQaiwhMIPqX03LiZL4RUW3/ekAv7X
rsrJ6cTV+ZouRxU1mh3VsSRNMWrE+b7RTbWMtkVfkkaDJlDTyackSkgFBto+UP2z
TybIDfsh3cB/D1jLGJUlXMmqiMX9EE5GzyuVr8vTfwT/OLVvmnLZgZ0LcIJVK468
HKfFcs5ZB98mxJ4UNXwnUpLgy41RgjY/r1B/OKz9hLU0TSjnnCZ2laT7FBIgxjZL
3ib6xONfVGmMEYauICfSiJCgF0R5Kio+qFLLep6UUv/Z8Fm//ECX/jfoen4dBFdm
4J2kudVWVXr+9pIw4FqVfVg1+pdVhZEIR2mifFHT5gT4yx2bowvsQWUESIm7tPO5
raEg1MO5xGw6xK3T5ALvcoA47lAdFbLpJTyC3/8LKLmv6SMxlmYbROv4bbhvwHGp
3PYGRUbcSQbe8dKsSQjJ9rn/5njknBxu764p6e02spdgu0jfaDSiGQ4XS3tScDye
fugv8L+mwwI8brOtV8mbBkWyZJXLUk3hG1/ENRiiBSroWrn6YZLhDe3pK+CY0FkQ
whZtmoWDU3dnX0ej/pw4rv5g6wcv+8bx0Qi/SHo8gwmGDMMb58yQq8GyYEuVoFzh
USM+aX50Xvda0KFlOqUu28Sem0lAuRNLqwPSanOdMAP12Cf5C/7M5cyPOxv0GMBn
N0jMagn0klg2GN/5uT1Krd0VGWPeu5q6bOVYo7Vk52eul8Kp8Fq705xQupkNtrqu
FdFvRMuGpSd0b6ruhIBa4ngLqnGkKMiiTXE56GfKZjU1QKl2sKuOAosKYwwd1gze
x5iO5WMG9GqllPZOwHuHJpo84/hj9jHL/2fcmyXiiwYmgkdu/f8gTfWDOHPUV6xT
5aSG1/xlRNBPmUE7XVCp50P6XWGP2yyvYzt1ug83Ll9N5R3YrtXD74/frfezsjqb
`protect END_PROTECTED
