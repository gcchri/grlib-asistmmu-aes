`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UCcxoRzPYx7PV0zRQkLuVjc+TJri4rwkdICq/gxwH7SPz+ixzkBBDHW0WvyA7/6W
l+GgvTw2LfNGidPanVlIx8NCtHABCWKmk+cLSzAgOdHCNSWenNZnko1gDLmZNtlN
uXMe4EMoiBe41JMKCn+Pr1/4Yw6ncUJA9AAMGwqX7ivekHeobu+azZPB9g6EXb7D
7NHTQeMRY3hDEk1w67sNbyvkbuZbDi4b7Mmo5ma6mTd7ZYFU9scN0RxCVqxCH1jt
h+LA3Xb+CTwwsYD8Bebh/r6Vf5v4CDtQM9N05KDkBr0cQq07yCBpb2DFrLEp/0i9
dKw2vQsoKGkzyE1VdQPAQ6CNbZDb0uxWJ5WKUHIF4lXWm6CB9iMRe+fQqnzkZj9J
Js+ch8jluUFJ71MK8Z1+gQ==
`protect END_PROTECTED
