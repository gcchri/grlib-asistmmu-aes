`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gzYFJv1vfw2IbWfC+yv6PnkmwpdDj90d0wFMkZVAIrZNWVqtrPfuRsGrM5Z/4EZq
k9jzKEsCgsHTyR4GWxA9ap/QVSYOpcRmrahqPFBDpK+8b/8K5q5NjVOVJMHEb8YF
JNJLJo2WXqCYN7gngeCzu+M4C+fIgYrEhLdi3XzbLVXsGi2X4QR7PrqJTQagNr0i
1DsYBTJUIBOqPnIyg5u7WvSedamubrNDiRZrXLi7cLdEZyfmyAnUvGOkoMGy1AG6
Ry4uJsWGYF9B1RzD93SC1YkrKpF96v/Y4bUSYB8iAAUq+1L3Vgm6MYVC5PKQ/6uW
y11ZpEPUiGSPRyZj/AKac2nl+VZx5cP1zT+xLq9+TXJF4IpzDkZtz3E3JUK9AcSk
oNpxAWz9judmF6WvUD0r6Q==
`protect END_PROTECTED
