`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
idb76vvqLG/Zj1P/p45KWVf7gJiuRm15myfWHOE8d/GubLQVSPRoIqKq3A7RNaqM
ngMHSL8a87zLsIAKpiQMoY9SjCWZWdSet98JDm1hvzNwf9zFF1LdUfTXtTwwGsQz
PaVuJzpa/Cc17cOvmMQlN4iCyefxTGUOGmep3gL4VbmfiSZH7SVMva5Kbrb7ICWI
9LWrR6WkU0T4icGlz8LrtxznI/4mUDKBN+QZH8GY8cvYLLtoU0Ay3WSmStF1rulE
RZTp2+cc0fUESucNOn7J0ghyfFPY+hK+3QuyqXmA9jistgBSZXbyJ61ryAhbJiBp
xNGA/VzPUZm5xzwn48b8lNPQSq0iQdg7OCKnf9bsx1CKCoezvgzjk8iZ73gEtByc
gSRT1cQ0pqfjGD26ZRb8+Va/9cXbXmivPAzbumRetivtKBL0eh5AyflsyLZTZy/Y
SWbTn5tdG50lj5aI3DOs24nm8cEP7B64EGNDOM4gY7VaGWJoNW6KK6HDc0ovtJyf
cOmhLY3OC2ZhVl7G/0xmbr8Vj832X4BwzVuYqxSYScCZvu2OCRTqyKEOskPbFxwg
t1MEpqKwwAtkkMl94r11erXgOo6+C4kIwla70lTKBr0F2YoJQvV6mNEz7ZTEqMlx
NHdRjVDA/5MoJUmlCrewgA==
`protect END_PROTECTED
