`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZqzlXHMhUahlmf2Z4NziV0jytxYoP2ZfEvql5BoavK4Y7noUz0yR8/5oeXgBKvRo
bOk9D3nyhC5wf+SOH2LVkC/JyxzQmr9m6YmNQ8EUaJKv+epFQRVhNH7PlW0Ma3tE
TDgUpWQ1VJ187GRtCqnLpY7UDLEbi9ESXddBvTU98bJUwY1FAnBmlQzd3NEUfidv
ktHNP+TUSnBqeOLnn1fMkG9ipslacmqQ+p104R4yvHeXKSmlcql+oylLU0FQamfE
BnRt3v0Eixttlkg2WFZKiDb9kOsRlNUcf0uxgd4Ejmz9J0UjHhsqOPHIPFBxD1IY
lbvqrMZHHi8YaxDYASnlKd3/3yquJEwgsnLyUtVQljIOg0Ql04CNlHqGZNvUsUpR
TdVwzKOb90UZA6Jib9Q8hRtn1+r1rRiuCGPK4vSp7ivcCIMfEHhRF8n4ZBxmSMv7
O/7+xeXrhbS3Ps9y2IHgr4/B8zBKRWBLT4BNuDLCEItO0RZKsUEk6T60kGQyfEu8
aNtjCj3lpa1Zi5Dxk6dCIcG2FGVY7ofHqxaaExgJHgg=
`protect END_PROTECTED
