`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bQ0qBHqsbiN4B5JGyGo5Cc1UBbD+RJLApnksWhESm0n0xheOc5YcmFUenYjbWeMN
modOoi07Qx26Ce5aLInVMAHk4qKAftL9nWywHE118NK6vcbsJ6ydSvzrZVNBD/rw
7/P7hhvabI4G8zI2DINMUFT82h3gJEL5IOpDdhlf8+UjimboVoIml0gHJXf7SrQX
CsGhR7NX+8Bq1gC167OFbfZ0BTIhbXTjCbNVP9EahbckGrwwkSn0f8S3qVRdXJfP
0VrqcRtaFiRjn0R7dJ6UQTncGd/oYjpwR++yU3VDXzl2lLx1FaWKwHW90S884WPi
GwMfTWcj9InbBr8t0hHl0wRUegJxXz14D6rNKBUvzrc5O4qiF/DqaPyoGMaFeWiA
opBNsuwwU27k+/6PvvM2JiLkPfjfDTTLuSQkUKPO4w6cTL7uY3H/kK+Q25M9WFRa
qz5oAMwAMjFI+SpruI5r7L7/wIjrSMLLsz9xRxsTmH3MncyjfU3jFx9hUsArei9u
4RJ4CSPYnggSSUKQHdR07iiycJ5QocGTt3fH0+MYCAmp6Vwo1avws3CtFr7+138W
`protect END_PROTECTED
