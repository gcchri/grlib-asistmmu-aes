`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b/gWWcIKC3HigcrbDldc+mkDFrE7rElt3L5SLpacWNi24h3IH9+c/HvFlUZ/7rss
bWZriuzrg78bg3qfVHc8J/bRl1PLOLCFS/UL+b09IVA2o0alxu6blXkHDVYfgJAf
RWWmSREGsIC72Qu5WXiVT0UJe1mj9ApLxoYJpzTTg5jDiBp9AH3vZzUU8CW/FGBI
Y755F5WLMcdWGvwUnc8XrrxyG6MCERH7MiZMq+7JUAsoHH32XZSQdXjRDKcFHFqd
TTEZkSXuWwChdW8S8PeH3dphaxorl4t/dz2+/FCbK4a0S9Rze8WvkuggYfrEbNly
QMjFgOtArxolfuqaCFSdH0qA6sQRF/DaIlBSay6yemutHt8xUAel3mVv6x6Aw5gq
a/MUh693bgZGKuNFFTVPP5y/Nnnaro0hmBHqOXzKb+0W2iAH9m9l37XBc+ZzRPE+
EGHBtNxp0R5oGxpd6rKeGNbci6Dhk8yNVbYkhUOSBvjzAiuXe3sRDjUn4IECL/e9
rOFTaj6v5EFlIu5hdiMXpYKQ81dOKyNewvoHyu8clYKY08V4Z7XGrvfremfUGhtK
KqNmTfkOg+BsmCcxMv93CsPA3ckr5Q6GwyuV7krQJtvA/xgO/U4zaODXrO/mf3e3
YMC5isPE5gvnmHId6qFi15pbxDppmflzA374ft6Ez9+GS/Oqql5d35rF4UUf+4BR
7yOU03o3vG0H4dtXs3vxXzl5e58kDgc+e/O4DUXLh+S+AbbnLrT8fwguUkGp1PeC
0fS7breETBGrEettKQx+nFa5jHlI3G8k/9Ao9bgWOKjWZboB5xflpjjx9R3hwqtu
7TUnCXC/hDK3nEVUs974s1RSKciqCxQklGAusL2jGck4OsfELVOgSdypFzt13wUE
grCvPMsHKyOdP35m1/mfC6ohxG8jjRVgjuF7CKYmI5QbfcGB6Vtc0gbSEESkgMLr
92aNxARUIGdygYoGLKUOkWNKdKyGkPmEuvd2etfD9hTm6lc6NjjL+zwdaAmfDIDa
K+fHnWaOHCjpK4EIhbVacpkyCob/OzJH8bv4FH7XiHm9UVBLcBHzmN8j+pMunPPa
obpxnlMH14ZlDWgpDwpd41o6lrtvE4loSaPtrBaFJmYZCsaKnrly+tvnO6eJMoPB
`protect END_PROTECTED
