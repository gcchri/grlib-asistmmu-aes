`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5y5khm8AUHx4g9z4kDbXJC3og9L8TZAQCAmEtulSUgMqB2doHg++5bvznHnoXMZS
vuUDpKP+gKvjq/Fmp8zTxqjD2qrq6JPGe68fFn12J/sx4U8WVF1DLxtCz5s2tg5k
B7K7T+0nK+7YUfsBdna8MkB0tvr92v8WdmiGBLD1LB93YQgQgMYWhH9QysAMHkZs
EqybUaWfwxW0F8RRduTguzqYlOov5q86KOQIlx9+NQfMVABhf/eUe7/Rt43WXXw3
MOYVLEiEBOtCQfXjSVmt94ntNozqSPHOTnQ6LSlcpY4F3cuFRNpvOFKPKuZ8W5g1
1ox+EYQ8V7FrOLmmaW6iErx3+V32DQAH8qMG8hv5bYeiPrz/zmOueFhhidT3xtd7
DL2ZIcKeiJvaIQa31UepwRoQMRBakZRBHUYaLGaamiOXQ/nNLl1TP5hmDzggiXT1
5d7ag7X9MNc/HGQKADrCQj+qkqxwT0VwBumVcW5TcZu3JR2LqAzAnOfa4IG1QZFW
ACLXNiCJwMhRxYnA4owWH0Q6UgT3nEbkGyWMpLvBKtd8LkaOZiHfPbbRqsg7Z6M0
kiQkI5TiWbdjbCHeD3XtU6orjzSpecO/pr/Qp2GJKFVs9xN545La0HoueLySpJqt
qpVjdjciPRrI3iWnmC4MFg==
`protect END_PROTECTED
