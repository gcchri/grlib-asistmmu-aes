`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JiBjXZsJSCXw7HAB2yioiF5pKmN5RwR+GXFIwoL/+j4zQVlMf2xEUXbLXlCjKcT2
0SsmnjOyo5ASvSmMy0YU0+booKNKq5HMExrSGYI01EBRvEv0cPTHv4QPwn+/zlWE
R8+a7u2DJUK0vcRpFE6lg4e7Gh7AnTLt0IZKvO6O6c9K5YisB9mCEHjoL7WjQKPn
fc4WpmFnW4ni0zeUbBVqDE7MismICrfTzN/l54zhC4femqCWx/pfsd86ZAJBaReE
4CrNL0o8cXMCgN1/kH6uzAlGxOhRll8lnDuIPdfKVMbgj1QH2Sdnp4meo3KI0tT9
XxzfFAdh1lQpSDhSUdnRGP6D2kC/6QdVk4Yp+WB7ZsORq6ZQaG0q68G+0eZgKDLM
QW/DM2EB8GEQBbXgklwPBg==
`protect END_PROTECTED
