`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p4yGzzlo7yBxnlbhfrgGXVhMUFHkjpy95xIUb7NbbfIw1kifFWDlJhfKpCagHhng
08BlqenRQRQrhfBwKOgkiZN/ySH1JMUTjbedmaIE5fD5yfPczcnTWz90T664qAmx
UwQQ+uNOaXVjgusMms4ofiKIysdel1StSpk21KpmktyV9WEmBcLmEW2GYZn8V33J
cHVfSLcS5+qG6f4nafXuZctY2FGAMKZiHN5vm0gtvL1Hk0ovWbT1Fqfor5/w8B2s
nxzODH9muapn5fn1Jk0n34jGE5SvVnbjLVyYgPAUyVLfhtQgyjMnNfSDr3GBkI69
semz2Uz0tfoyw38UNO22QNrN9JXVS3T2eX4i8GWEV9mCpTBBMCZxgzSlFXE21N0i
aVovPTrMdfwV34QFggV9DCW9m3fW+w4XZt/54WMnwLtGrfWGfFqylRkqAm5Pkcbe
Jx9N4EwDEbuIV2D1Iv1A8jewmR6roh6/K507WyhQUKX9Bn486YKXOxd6vC1L5Wa2
1lgjLUv6H64nMTyD7cZs7isisZtVkb/yE9tMgV0y/b3CxPRmiFg67e3UkJRKVy13
O6BxdJs/TbLYZ9gr6bLd+g==
`protect END_PROTECTED
