`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zWVV8huypni7x8cBfYvkzoflgWc4HxGmoG0ogqG+YnnvKwjBKzfE7w5QNEreL0ZI
b5LamBVe9rhNGlRb5fWBmlYqY2PbiPBcUI5MsnapGsyKVToZeRPzV2PuD6jSHnto
+Xw9uR/075E7XDcsNBNBgaGego3yImT+NHsC7bzyyjp2xn5BTY2lMMjs+htwTDLc
Z2fE2fF+4NAhnokzmocvHSrR2asLciygY02ZFDPUVuGDaYXxUaDsJ6TSof24oMJ0
tiVgCFSeep1RBV7Ubx3e6+5X9xjRzgfIOr2hjIDFbItWkb6ojyKQuYaMfExoF9BF
XV1OwJGusstlIAeZtfYEMWszhNZco6TU2TpQPEGTy4YGKUiU5zQ3bOgFhzgUP7ui
VUhZSk2Deh2Fq/XsxyMOeCSHP39BLnN9sH9BvWU2y12raY5SN3SkOE+jZWbJBeOn
VfztnYO0XRibK0bFdcmXrmuJz436lyQfflj3NToiDNN47s1uVYX8OF17b/wtOaSk
7c442zWpNIsnLtMFwEOr2CYDCoE3b/vhRrSrDPuMdjRM/b/l52ncjLZJK9QZHKSc
JXDziw3fKhPJFGJKQCJ5X1eQ4t03y9oiY5PjLYoFKo0OQzA94K0g+i7rDzND0i1/
4U51TXwqwJ73x2FrvhZQt5GIF4BiXU9L23Yt9Q6Q/x3owlU2hRnRFXjzyq9o0l62
`protect END_PROTECTED
