`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
csiiKR32Kvhb3E6jNhDu4r+Rf5FlnU+3iffv8Co3BsLPm+nuwEe/6lbLKr4SfWc3
HJe7VEbtF6z590Yv9pETgBAwJrLvsQegW58M9h3A5WbGsn9bT/SiDDeLHiDhTtzt
+2jHANBu+Wkc0MwlN4TqY873qqPav9+bcfXCYBHiKTdjOvu3FMsXc+HVKFgQgTy0
0+2KYZrSx4ajzB1XjnIpiIEfWn9C3lSbkhgEnxrijA+zKdA6/40ksSV4r/jEPnEY
7vKnPNlCc2edDOg+k4AdNkvZLb0YR3mDzKRwvG//LQWwJCheTv/kLiEbWwFBpXky
9RjxAsYO/B7xe4Vl4pYpkytPaugq/MXflriMQqDa1aatqCUvMQ2bV/GcROQXVhHY
NKWs4gN3FstoVTSco6Rw855DgEf7MZylSQsvFJ08JtGgV5dHVNXEmclb7KU8AR0N
+PS46lcam6cCDwTkrVFvIoBf+6Nuc32E62OVLJPL2vT4PChnMv0A5RxpgTT1IfZH
TZgGrXXnxx/q8fPlw5YTD3nhccMSf+QbimSjbf2yZe2xhkYwdAJaf/0QKsDTucG+
0+A2nk/B1vMT3PFYv/O/Ra/tbsom9BOw9PLshq/UKX9pp9ILhDaZtMZ4zTBSM5Fm
`protect END_PROTECTED
