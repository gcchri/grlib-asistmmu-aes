`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pXLGS+y6Q66ckx3jkYTw7CP4z84DxuEEWaeJ8NMERjJ1KU2/GMXlDnuoOIY+4AIp
lxdfYCvFqimTPgpt+e6Yq33UiXnmAPCFecGYA2NC0HnFHjvpnDS0KbdFT5mMr6mc
Y23B955EtD+ts50Qn/zgsVyjr+RUX3q2B10Z/nZBC4fDnREBAuROZNjdqKX0mI49
0gGMzhF5kOXJejrkq/y5P17Rr16NJ8MIzft3ixSpBfPG20bnzV9GeK9ckmg6UEu+
/kM6LwSYypX0CBTgSwkwU8Jo571s0S/JfM2EnZMNvGxaMVNYaq45sICpvPhnxqfK
5iv4OqcXqE0wJs7rlbYdgxLN8h1oh4Mr/Vxo+lSg9LfndqEki7hEFLOmDq3AF/4O
iN4J7ZI868JKkhAFxC7VbbCSZcqXY9thBLsW51ZIVGI/0t/neMi07Pm2oiYAkI0s
cfYGkQs9Yr+sSHk016hWwG42ZjzH+96BNIFzkGHMP9KMjifXE68/wPLE/T9s4y0x
9A2TOa7QUxoNw7XM/ddaLcKTx1wOMYyGaukdXHHOt94R2rg73M0TaUjMevzUYz3g
ipEkbV6bIFvGeyI7SB/7vW+5oenRSmIvS8rrIHsyO8AivXGCqR/CYoqzgyL/U09W
qTn/L9ZDF0x8W2BdrJM/MP/nzfK6x9JwMSE7iZ+I9HOlhWmVIpp6FeI68bSBbvKF
MdK9HgoyYl+TQiZUqQnNDcaOvt/lo+RjJ1pX9s8TZpK4Qnj+jBdVcF5jH/gFBVzD
SIsPXfYuh1oAbX8PffduNYJgcv0zWGZkvsCuHSnEPfxuL+XOrYBdy/Nr5zpmCHU8
y6tUGpfVU+ZE/bOVk5vv/ozN9rwt4QL+i8cfwgwUxDOLisekuB9gCuTzbrqdE43w
IgJg9pt71xYmT5FQnc8hfvYDbuSfS19DajovnpVKOjjm8iPIUX7R0MV8vpnIo4H4
00D9Ubbq0tDhVraVfNBZ+zUae1NcoU0f+VZ9vKee4LvzhOuEiDpND2nf0x2JLPMz
JWCAmXiGBRXppksBpvN5Vd34VwGV6f0Zy7Kjq4Fiwl/l+Dsd/iGTpP7qpcNjB0bl
r0gen5T1WKiYYEyeUsxjSF4hZTC26QmnDjnOhk6B3mHVa9WImCS3Ir65/7rgltRF
ygrB7invYvBaYM/GoNI+AmIF3Kn5UqOeV//MTZRVF1gOacrPNXvMt6yPI7yNl6hg
TZa5ziQ5BzvqAJxSMbMuRS+vmKl/a2GITo2Dz30cdiYHCgR6ik43Wlyr++lg70sX
4eUQ+mlyv9CmfqwxFvu6n0Et+sbSOJrNmfzl8MVBhFVCG+iAGrELJrMXLgTdBYzs
UYA+VaIq7Qguvbil42hRvvd+NOrE5mvLff0Gs5iOOlcUrRVvHfe0zNLIeDD109ta
GRn/cWBUPSTFVsRHFQp+yoY22A7mE2ObnUa1mSKay/tg4sK7SU1HJDWjD9GA2r7C
NC+NUfJbEfs2XH/7BdoAdllpw11obxX10iWeVnfNZ79bQo1w7CRg0ieU5BDVAGK1
BzhF43R0uuXRmNzeGwp700ccpQWPOOYIHhIkyA+kXB0Xr8UdkTF5jIWQRBwZid/h
KLdAHwXb4ey2Kq1WVSWveBFP++elmREWnjCso66ZAvyITpB71ij1VzT6DxQlCwmW
E+82yVc3M1VIDiNCmvF8KceI3brGaztY0Vax+RMpRB4kDZyFCic5LUZMUlf6XwbJ
ifMQbGwPWbguG9D9IVCRLje+fnwM/Bqo45+qId5/hdINnlY2GMCo43V1E4vjsM+i
RxH3DdCgdFVscNlUdUAiWGj73QwsfgqBXrIYutYthEyo0iUzxSzYuvJRjK6gl0qm
slwnjdE41ts0h7EgKArJaeGXlC8IEzSV298y7lHMFXgGgMPj/wMyW+YZzjhj2FzT
9PT/oTxU9deDqrmRxwQ8+x2nuG6Trzn2GULku7X7efA0dAKw9AZ8RmnvHkp1fFth
qQksnGpVR6nbCizRV/GUuPHw2Hi6poTZkck2Qs8fSQsIxVJ2yOfZQnSVnts1Zdc0
QIQ5ilEN9mbBwMT1y8P5LA4fzUutBulG9Bn6N2bY3OW8LBGksz9Oo/Fh8BbakBy1
6BmqC7P++6Q0CjeRzaXa5kC11dqhb0k3VEY8oLyAMBtYLGI9s+LOc2qPJbHFsKIK
RuLSmxPGamgWsVslkh7xdF3GevQgR4yvssOhyLhZWh2F64fbIDeeSra6cJ4u5koK
Ic6PfHa7jdY5wKd3cgTa7C+uI9xIAm9ZUkcUpHbIGG1d7hh2Hw/30UWfZjcJRVZe
SQk23y2Wy4/iQjjKfSQBN5rkWfCB/lZmDqsWpiAqsOQAGAGllVWE1F7F5PhtBecq
pif65hDvLtB1pwSGz+f7KgDO0pJTxpEfbUC6d1Kjsx+3qvAjsSs4RLXsaVgH+Ff3
GR/KWFOPwOKh/Qi+pHRGFajdshcATBQJJQ9uOLYq9WCvongPBaMoYy3rPJUoVP1u
erN37hPJ47ZJbzJypP28dIIBp7R5Dv819mPddMvU+0UV9l2cnyxkt+FnQVJ/kfJP
V3vXi2knJmYh470fCquNdkfCEruTNB/BO4o7Ye5rtzJv26UIiA+sfPY1WR7gpVdy
oS9Y6ijUyCUMaVYX94J86+z7ed+bClR1USsYAZmWUz5UVkZcrkj6LcLpADaqlNjt
sXORvNEr0KhKZRTWnjVsxe+s6lblgEHEvLm5BpE0rQX4bC7EoEQe2yICpkH9dR1e
lMo70fvawraMYjUrPayfboyhmDwtwTDHxXhr0OQua5w3j6M6X8aQTQB2CTZwcjdi
n2vAn230W+42HYavP+4JTCwrfEq4Y1071yrxo+IZ+km8fwh/CJhC9NlrH0EnoIi3
qgnUllcZvRSv8zqRx2viLLkcetDuIKrsZmB+nP+vZFmIU+bor3+AnQbTVLPUu/af
oLmvy6evtkxB3eyjczOtVr5CXgRXICpKin18BlLTlJ9ccefMmyUD6FqmOufFoNzb
NKAVAt8t0o4jDx4zJJhTUawEheJcG4U8zBH3To6me592M514RGstn3ilFj8qp38V
47NPcehLm88ok4i0/XiHT94dJ8WepMOTWVN04wpiOK2jKUhwDynLDBUP9E1jTjiO
nCYwPTPgrFS4o8STIil6vuvLk4uZ8mr1LQ/lZ3OHjA63unr4HRSVRYdWuezDGkmf
JSWJ6wswrEhmNYOhQGHq8Ca50AaLnYKFMDiUhbXx8nJBuSageSMM4LEFbVkFNKYD
pTLZavNxSDWQ/opc0b2+g4HrU68q4ZETy/UtOoTJ5pi4qHwNj/LbNmJEwvhyPzVa
y08xn+uqKa9qNeElyKAS1eiClzn9CAy1fuoiMLjiXxn0Cl4fbl1ilyn7Bimc3mop
e2lfy0Ua/ykHciEnA5e7Z0KW1M44VU5v3idMxirSDfmdEfYeDSk4LOcneFksHiXS
YxKYpxo04EMHMYpgIz+pDEVKXI4liG3r/XEzX0LeQJS/GSMsMPA+sBC0TtpitDmG
KPe5iODw1jLS1mn/XrMPXi/URYxqOdDc/y0lTlbtM7JMZ98tk+1rfDX/6g+KIWbL
UyRmtpSkuJgcnnYPaRnT/baHYBgm1YeYxPhdXLDiuNYJK4vM3oSaMq3G1FLX9Nxr
QQfL1uxCPFWN3Jre8eZlqF0uJbeLocXamEQ+yuo6VRiFGreLGKOdqeyIoSIDNP84
RYiEYWPc69bvIUikhVo4IPvnkd/Du1/RWFSt62iNQ3eQrnhVVVww32diOgBwWfX5
ZpGF1X9Asbz2XbHadQ5F/5Uev8kttcBOYqcPCvH1W0WTruIhe+/5N9GtvpPS1hKm
mPrz6Zd6bRnJMUpAg61u6AsmEgKHTJQ+Db0ALdQd5ocqhupYz2c784HJZ/0PXh+G
AyBzsmwa8UxroEiJFnm1kopSqlA4lO9K+k5A4eztZkvqtoFucM/6TeLekjcSYjkS
Wag8MQUyjwMk7vAS2JFenLQOvFGUFLyQXpX7ni/2GuYmebjQNqLtrMZj57qCg0pO
EWq6p3jL/LZxLvt2HYGLBeggyqTu+Ydi4GNROVwyvZjVk/3EtXJHhlI3EKbqGqJM
HHQcuheIhZvRFRHWBJpYSIxqTnM0ZHTcUtxJ37qagg0GGbgrPCiOg0et9RDWVe3+
FYnT31y6Zvk9BTb26ThMS/udiYjdfh9IPzJguiDN8fJm+qLYFrV0z87SbuIEjLKv
KQzKE521M3Ja9DzVGZiF3S3jySr33/Cr5SxzlJYAzlh5ZRpcei8EHB7mT8jGbwju
h07sfyeIvky9jnZzeSv2b3P8/nk1Zz124A5+ld/NeLYu+Vskws6tM9mkGS+k/Q6c
cDJMAz8s8i5hstBVYXomfd9mEdv2N/nbGHr/jxv9LmXhUZzfbp7bXbnUN5TGXhWH
yhP60CIc2+w/YlZueTffTm5HizaEdMc7TNSsLo+YHySj/qakAeOBNOycZx4wRBXm
ljMFwsU2HDY1T0aexkAlV9wa45DhjNCxi9FmvMhYtlpK1Y58/AarR/EcPRXohgKG
Fh8Wr6E8/xeYlLZB8/IKUDCK9/ZgF8CYw/qhOnG24KQ3fsYw2nln5Ks55A9mg8Q6
I3TfUVLaHdEyt6NSlpKT8jQpf5D9SzSSu5GB1XABcWkoTQDdAvjYq/D8LsPhU1Mt
cF7K7AEy3xKcCT7JzJ4fpO2olPu5ObpA8VrSGU4sJPQ1Zns6ht6BofX3/0N3iGMX
mexIFTu/5jDIjuex5trf6bri9g97+90QZAHK+32LkBvK2JCvz8ETkh61hX7B26t/
SzZ3PL6Fqx6GMZVL7c2rXe21mXOUTlJZ9N4izvLi4atGIary2/cYzNGFjhc4uv3E
41YyLRYEM4voKG7rK0aHTlsBhg1AqAvRrL8IkZeV28oq3EnUHEQX4nMPPqxduQnM
lf4mcFinWpO+3q/qR2/3/FV/y1zR5GAdjiqB2jqyhxwgqsoZ13Kix678ObQSRm18
Q69C6MCCmUPMTCn1E+LeR8X6/twDTTMCBunZo2WKfWocOPc4lh8xVY9yckLgROg8
DmRRCFBJExAvz6KVx5kMisvRkZmf0KtSLdROno9F3XgHCL0X+v/w/boosl7KLamf
LFWWrEngVVMPu8th82cINQcKyC2Sx+rsjk32Jy/rxv6WQmCkqYoGC7b6JpkMZhpW
1B2eAsM2h6faGwD09gCquWj6xiOv4fr3DfRTkzhrqUj/KRC6HATh53aTcDv8z+Ps
qhiJZP/Jf5I9cYszHyuIm7qgXkoGnNpEDbW8uMbnd+AnFqZjguJHc8NW42efBc+1
/uF4JFzZYQftQpSYfo+6WhXSWVoMp6JSS/kBVvANkvwaSfnTBn6mb2rSWRvWPlmi
VgLyUiSj6fBVXcNHRO0M1/aTpEDZalIfNQ1XlX7Ts3KypCBudPFoF+CBicgRl+UU
JBy/YSxLanjfyWKSs/6jPhY62eaCa1FtH07VfDU9ticcHCQIknZmpWm0ZGq58tG1
N5L28aF9Fa/6fC0k7s1sKp3auOquWoSx1wbiaMW9kjymMB+s+wpmYyWSjw7wP4CP
w/4maTP1M2GGJg3tXxuQzTLgwZB9dhOh7ibUAhMQAJQX4cSQocUud7+hJJCYwpab
fOAgyaXK1aAKYdB8/0MsuKXPMJlMqRPBzxOvZBAVlVOtsrwo8kD/y5xLJ3AlPk2l
iWqTYL0u2gfs0VgCylrRg9U9fkWGTtUo4VipDfI58wqrtM95aFg9c4FxAQ0EDBoL
PJ1oKLnL58VGxqSLbzHNYi89iIax6Xu57tLeCSLOqyXzpqhlyUWvmibVmbSMKHy8
XXDW+J4uor04ZRGK5iHUMhCu/HY5U8Qf5tq1mEwBjOQ0NYl0Z9vxsz78EMGC2bq2
lK48pzCWsU0Zb8dhRoB69edS8pWK2JRjhNSN8fKZsMnDrnDJN4OQa/VhYYLH6VC5
xJSLKnDbUmT93RI8zizmlwtObIElp9AnUNN9y32t1wyXSh2SA7XLvBpCKP7MrInk
w/dcWKpMnTPQsWZZRrP9gB8idy0YPPB8W0T55peglWBXpNzKJpL1m1u+dXneCRRw
xdbMpDe6pMH69osO9dHAgNuo9iEimB9XPsgXa8szYHz/Su/hK2fbWSxbgrh7uaq3
T9ZTfGaRxqTRu2gi/369d5DW5Ahs9hmBbLU7yWefz9OqWtSNeuyiCEWhNC8cHHE9
JeZJ12C5fd1XPe2fXslGYirYfIi/AoGcs9PU1qQOAnGYoU9Q+AOMUAYQ5OnBk1VO
NZbsN3wFWee08cTsfBRz4dPWnOu+Un/lvp4bxyb9u52K9aq0h271ZNutiBtWBs1s
4JooZ5wp4avuY8rqVLE8qZhAvkSWHAHb/dbz1dRJSmxYCyt8U21PU9YWrpbnNc+3
dxmBhTGvP/tIBcRygwQoFP0KJ67AEPq81APV4Inz/b1svTTrlif5nysx+PqtKnw3
u51sYvnfq29ItRWFdSZe0GjNrLNdqOZtpTQiSWY1hixQG7ZBBw+A97uvb1EwIb5Y
vhEUdGujGLk/w0rDVlBATmCHxblB7nOXRDji9tSmt0yOr5yAocDM0491+eCfbJk3
/K/jv4vfl8srNZMZxxv2Hh7u0jdUxzLG2wKwt28ho2UjHwxJUgA20/vquGyXIixn
Qkrc6YnpXm4btiBA2bYIPQCvxuMk7Cvl2mp2d4U9/y6aLbDsk2ACLmRCHkGorZ6l
JxMr6hysBsldvYjNo3mSjug/64TVC/WLimmzy5U2wt2bodLeC1JrtI3Gf96Nr4zU
9s09lHnqTV6IxbCmHREOeXwq57gpIyyR6LaGNFK2dkvjwzeQCmonxNoV77li/suc
0IhAvB0xinZnc1FrBjwXJ1QDlghD2/IDsGw9q3jOrwUIFwapw8+yRQu06bxJhbDn
OdWQ73XSxJL8oCh7F151ijvnmeeo8T14apXvIPFWxfF4pZ19LM4LtvQ7fS12bi7+
9+W0JTsXt0UodvWUV+bMlL6BeTDPrSEgpgA6RLUqsxnatWBSVIgxvG4Td7ZQ3mNI
a5tbqtNcQscRIWodZ6uu9dkDVZpTRkfhMbGwoMWF35e1LZlVs6QRxVEfBkXJh3fD
jR/fkmE+qyiZi41Wr8UB+wbffd1N8PEAgOb4GLobExbXXfvXLCfS7JlNdFLYXVGu
2WGGSHtGhAHZWIbZ8WAib0Pgt2CLhyg576hvDJMLLvwM+Lp5h2Ak/zNKUgJMq5LT
Fgov5XXeuDyT3SEn5tmx9mLrGmYUcwi/zCtCmOq1O4kraZuWUjVloMWHR08DkG3U
mWa/3CIhOME3mJ4rdBduibxVneRnNQQwQuWkK/IbnR9wK86Ukw1TpXRpszVEy+z+
Afmp2ux5dmuxwaTfuTYnmp90cZ6s7fWzsxcildq7QUy15LztZEaJYFy8+EuhXGz6
CTu/NPKZjgE9QKX6vLZ7BiNET+H0CPuFPFozqYq7bqHh58TjXmio4u4ANJr4jDvb
`protect END_PROTECTED
