`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
um9xnM28gsPjuGCSlBqgYwxfRvUUqQSsoLLkCoIf7FQJJO/cqHYcWlYarj5y8HzN
cviuP0LBqp/E/ukkbGryxBXj6h7030hELY7/jkOmH5bqiUIVciOWHDwEkkAY/KyZ
pgcgUkOBL4MZnoJzhwqgkuPValuDZNojUqfGpAtwPaUvbua5X3dItIoJKFmy2aad
CuYl7FLXbo5vM+c7NicNyTLSWh3XK5U53Wt5Op5LtgrduUlNxtQIyD67FSTpyDHA
RUorC3F74FH7EFt7980EDKuPFAc4Bjeey2UsryRPAOV9SDnk7nmuMDLmm3ql6UU+
TEOrf7pmKA8BSV/ukOuLVSGFYEw/4LfUqh5sVuqHFM8zBlHQTKHh++HSFRtktQOI
HFsX40WIYJRsD6vjjgOe+wIyV2FVx7cpAQyIrRBx4aXkkmzMFAKlENaa5+dflP1p
Zf4NrvyRAMi4WScSFY7JUhkhvwHn2FGi4C/RKacd9RafrmJmAXOf37GitjMSfIfi
VefTwW8zelUymU3zs3vuVfeZy1uRyHxw3XQlopnTRrL91aZZj+Dh3H5Occ90BSVP
nuDY15mIFCKyDHrp2SBdoOx2hdw/6u70ra+oF02pHSGp3d8TBXjAjKpRy+p9zCLG
vid4fLGfdhu8FDyXLus3U1BmsRjaVSBNrCzXeEfg6AL2ACtyJNp9jmCeMXUAmIAj
s0txq8zra81EJEJlLy+8vkbc04doiJXe7g2DGI0WMds6jFnlOAY0r4HjqPRoBNn0
TRbA6ZupROWLDksZ8FKa8NW5U++p3rnRav8EKLmbo/8uG62EeLr2ifcyxP5s5o6u
LIJMeuNhO6QRc5TBgZAdeUw2bT6+2PMB1MaI0iee34gEhY6Sk9dqdUFb5MrWWh0V
zLUlps2Qorg/AjcW0NGf32NSZK1k3okHTBnUxt6zLh8=
`protect END_PROTECTED
