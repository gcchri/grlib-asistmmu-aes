`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3UBZv17F8zreQQln3OcAdVCrCjm0kguYGXW7gN5z0yjOp5jXJ71+DTUo1Ymp8hDp
1bO0lKadp7NB60hml8gvMFksY5SexXm7pb1DQ6L0g0zFZ3L5X62htNl37/54ORGb
TpCcliRKRX0qV2wTfhLW9uGmV3Wwz+VFdM3bKxANpw+WXCKL2NJcHIhttKNkLiU+
V1RI10ze9GAAhPqj5uoaOPgF7dAA08mLdPDvyrfhWa/45NwY704d8cKB/oXZkToM
1s+MRoCQx9SjuyxCRx/eFUvS8daBws6f+eFKL424bVKGhBUmjSlO6a90C8JIAsow
6V1uv1ZgaM2EGAI6fNsU4D7JvYNY6PViCvWbLlchCsE4l5Bn6Vya5DJThmWrJJzX
d5slBOGsk55ugJpFMvRIBI40oWghlyLkmZyUEPo5JdTls87RajCH11riagN2wycj
Ku4ScqCPLaKUiAWt1p/McQNsx0XMY/hZZmx2NRDbbaw=
`protect END_PROTECTED
