`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1BJzKPA8VGiZLOBZUNXmKYtdSbKDVqTpCI2xNa7nKICyEgrZAJ7iAUk3IOirWaub
Rii4NwxUj9j6YrMovOk5Liw4imghQzmuCeR1FJM7TWmHwRUVy99YFcguY6Kz4afz
7Md7Hufi2WzznMkIi2LDtfIgpnT85OVOUDPrMQLuYpgRCVKl2hiQR0bOEAsdGncw
z9mISfT96Wkxn40jbw0gjyp90V60wgzG6SGjXiioYjzjDk/zBqnOzJZGM2bwPB0K
ftN6DoU1+fHMPLDClcjZ3iPp9lVldT2ApicSOSL3WPXzgPBfZnUnyfXlOZsbww/w
Gb0v+pltBPe1lWvy4IL+ZLvKAQw3Ec2pKSGN/pUJBktqEs1lf2UMsRn8kzQ3mJrZ
2mXQ3jrTQ2hynaH4UIjDZySzu4t0dSfpZQOvrcTs+Dc=
`protect END_PROTECTED
