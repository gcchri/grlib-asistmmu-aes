`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bw58GWCc7DEHRMiBJuMDxqSgaDxhgFTgwfKga27wyCHTzfkvEjB0lgfLMFn1IkXW
58q19+ZOn1koJZQMMBfFkYBP+hvnMtMYhEHyNaFtSZdr/aLivyVmuZggOjL8Gld2
2AUGowdfohpjjM8nljbKSCeeMYWl0AXO27pjkQFKy1GmleM6UZn9v+8DP9bsAzds
JeEnQZWqOYDMIuyIjT+ju3ihZ741CpHQ+uGKWcQPr0UaVTsyJOQp9PvrZMFcEN5W
FrojardXAprYjG7oVuaAX80gWgPcueFB79C6UsXWsL9uaB3H4YFTgJYaQ5ipBvSG
qCvgVHvHVklxxKiHgmu/Kx1Ak2ZvagqyKixL+FB6CgqARc9wTFiM2yU8YYibcxq/
qlQny0nHFlqt7e5c3W5mNQ==
`protect END_PROTECTED
