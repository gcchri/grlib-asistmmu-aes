`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Oc332wjb5SOH+R4f5CAtUuvwX/H7vt2StNGMlV6pMsL6zxyW81X3Qz139pu5myq
JN8PVGa3c+tZ/Qx3WyfPIJbtLj1+TFNjWU/ELkQidi94QLIpLxOe0sGYh2Y5uSxm
mzVUIl/1XO8iVOm5uaX3uEnm/mlLgcfIO+wfaX7NOyE8yDo0Z6Koepl2TniX4Fzz
6VHud2pVt58QfvyfkLMegVhQFhBgtGdWRu4QPPSFU/mYfOYPuP4eShC0zRdgpmAD
egCei+7gh9mbYE/4ASp6j90wd7/sLz4En1rbKcxZ5lvobjRqYjwlnwu6Iqj9Ix3q
k9BCrlUgewDG8xHQ2jL+Ry6mgQtLutB0EquIdLkyDNRlV+u3MzA9Alc+LF/dDa5B
b0eNRpYPgKukupwDq+AnzOgMQE4UUoz23ceTl9MiikxH/m/MVylZu70glw4Ab3oK
GuZv9i7f0KlaYjAF/ACpWh0r3x37zzBbNmtusESDrg/70kGoBq1PoJD6vIR/yREN
3bsd2ViMo0nqz1uuON10y6zxj0VVuNOLKPhPE9wpxm+qwPYslzQWEsI6fDdPC0e4
dyhkKUKd3v0SPXHgQdMNcgfE8VTnra8S6ozfV8Yekahdn0XCFUB26nsPFXIuGUOs
XMGQDxx42pdfG/jDhlrMWuSwQLP1n4Z+7mmtlces+TOY06Jls/js+fJUfKw6dLQy
J4W9xXvUgEywD+KzX0LUJ8F6YJkQuYPytCRTfXZGlilCkN5puVyClk87EIQzyVFs
Ez0m4HgXKGoXkY4d6dmEoUxt0oTjdYPxkpgWB3hqX4CBaagCfTznGAfn9did8iKD
+LU1rOK4R6yv5+/y0yQh0ymgqteR2Bj6BV08uCJMv5ubFaWxYb+/Z5ozPWG9IgDE
TRuoNbmYnB3C1/aqFjsGLpFWa54foLM9EoQDkIPF1ohrAFE4EdzxUYpVdzp4rS2K
VD/jg+J9huwfFW2upegg3MM0dZVFvkbhfxEv/EiCEG2oNNnEZqZ9DjX2ya1ckGVc
V2lxHf3xHHE+ZsFyG+zUXklfL62bzOyjpHAWwH7i7SoSqfbrFjFlkYJ78zvOqxFc
Jk7FW5/yanVkXZt6seaMb9NUVIMGmtfufPfFwLrVZfmLh12lYQ269i3GMZkpC/oB
la2/tXLqfxUWGfoaG+QAQ16elVIQXX4zCInAMqoJA45xqHsT6YKjSGiy3MNQ8idJ
82jda5kz37tDTNPIutCXmJmd3ze0WHQaUyT/J3qaZMBvOeiAhSaCjFmt6A9/k4Bl
9Llw3j+Bpv/Q59D5s6jQRphpLJClWO4I3qIU8Sv1D/XIHzn40swX+lSGhByCFSIH
eQqmKO4+SE5LCggOCgv3oE8/idiZyslojoUkl5IL/wTkovw9UAKY5FldmBmWoKTV
Mprub6XcL0FrjsoSHYXktZfCcGHasxG6j0FbHSFEMiNnDb+8oqmxzvtouJOBd7A2
H14hlkFu9qfqH3fckllaedzpo07iJnGVgprRNRB7AubyUG4RVURfKMTtmZ+bclzN
l9pyMjOxKHgeO4VruQMBePJuDO9HIOpHJ8XV8iVhOCFx1RXhHOGrLN4ivR5LIr8O
+PiQ2/cKxwL2fDm1pdExZsLNAC0zEr4JLCBPl+MLSKHCAtjve8j3ubm9gkpJqNm7
T5JxQz5QHizA4ODS877fICd30Y4cXUIPg8Hz9wCtzb5IBwPz2xBXXtK69rbX222f
BnBrJUvtkYD9AS8usoainee+Ko6goDq80K32N/8yT57nC/n5RBV0tV68J3P4lI7I
QjuzmmK7Ex3+dHDPDSiq+dH5C/5oln9vMNVCR4LrLlYe6mM/AjEESlQ/HMJMTkki
MpnoT72Pv5cLEMqMYGGmu68DEOnd09NbffwTEyVHBV7JRhzGL6VHJgnWcBnQvub/
BfdOsRrFlAW+1TRgi+3/lRUxbFHI6UST2u92Hc4RlhMDLxOgHXpfViJEDBePV1NA
yAJ9CvLkU+cXHC9ZcqGFlYEwwt+Pf7AKBclpkPU33A24ppBM7pVBounVI2aAygYO
F1kHrfJspdXLJKIxY2QqqwrfoRv03oDxpAdyqPy5l4fGlGIkd2lPgpXKk6JnPs9o
+m01MiCYnDXWs5Zuo9bXSkzVWkSliBKXj+G6bkui+4PSoi+P/ngiOPfjCQw2mI6c
WbCwy6FciHj7Wl/7W6pyDFXPaN2hM6D/bgG+b6J6P27NN+h/nYMBgcGiDAxfOPmr
pNCGCYd4EK3OUSOha87qh/Ta1T4yCKrZaeN1WfKsU8P9a7l1uM7182Ejizi/8iev
WThg5Evs9G4jSzficDXuNMI5z2FTUyjdRUkHcqroYO0HfrAq5QVCJE3Ukm4phfNy
6bfwPpgnEYJ6bDjjUDMfU3yQDix79KOtuC3F+NRxe0MVJO+aoBGvroTshccJjJN7
lekD+PtlqtrXvYZx28V9o+9pUdOU54MFJkePO3m1OHK0B4IpyX+/wwMQjibX0KqT
MSpPeRaGuU6v5QTRO/9LCDt9efkPW2RedJozWo/fw+SnEJ6o9CHByctz3dcTM+qa
iBZMiNW6f8tQoMjdYGdYz5wISXWNHy6a0tGd+0VSo9Oj5Fvz41FDHS/jKp9KD2/Y
Hk7ypGVh0gEd0SPtlXl1pAd4945Puq1yymaXzWfClr7eaL9gaCCWggey11HgODR+
W9eAxUxWgq+S/dCh+2PYMPIaWFq/LciDX0QM72rQhvXzFvuJaq3AEyP/BDU45XOb
zR/kOznvG3O/fWY67mX/oSUeMPWVSRPbaVeQqpekfUS0EKL5+MwlnWbNaQWWuLIe
6i7KzGvxN0PDqWiref74C1/UL63sT3k2lER3VEar9WmSPoxtPn52J5Ber7VQLNTH
3IKdcb2F8k08tfYrOoJJ4Q6r4UwSgb0plwESl2jSTswj8/f7XRu4pqX36TdgI1NB
cgvUQf32MQhAMUam0GErMbEcZ90J+ifFKlEO+MJSyIiXWZUkBvXLtwFcEbNJio8r
CUxo+GarfMdH8vpUWnRmB8c2s8y/iD5ZxIDKBp+XsZvqvBU7cdsGCH1iTRkKbdiO
jPQswoxHysVdfGaHHO2N3Ko4tU9UtjOXtnod1kd7yE8WvhMpjz2baOGRe8p3PvOK
TrvZO8Ncfb9M1S+buibPzbPf4Mwzt6LZTS03VpRO8el00vSq29mScOoiYzgRixNa
in6lHcN0LNOVqxqxWXTZ8aVbMJd9OFFZiGY9BkOe0G2bVZNA6bGXfB90dIAl0Ldf
nPtr0Dsmla7d1PjqFmvtjoM/cPb4qHGKoK99Z8Oh/nPOXE+VDVNpaGlkGBygSQ+0
DZFLeJUR513mhOJ/NMYDW+8Bra0nPGKugZh1cnzmbkd/32JGZsI/NRDsJInEOYH0
d9KXtL9JnP09eJPlL2FFzsslK/OKz/DpwgNoGYfmU/2IviAHpB9R2EKL9Z4FiRM2
NNQ+N996QLHvGj7HI30k7DNsHOnT6nzvMpIFzXgB2jkRVUblhMqN3F2AODJ3iImT
fZYrPN7j9MKX9kHuIMP0zo3osJRUFePx0mXaR4n4DVkC9yMFjkMOgcLvPpXMnICe
2ssEytD3Nzk4krcEEASfI9rw2awSzoIWzqt/JEdXJZiJpMIKRW6sR5fCUwWT5hZD
9IcaIuVbQ9SaJpEmJPt4fPCVKCG5sWRh3eUNihxeNmelQjkU4aRruT3fNEiSpv33
9o5YcwS9XGXA7V2xrIv71CuxOYA1gOS03EpRl8bQaeL0HUkbovrxFn2El6//NcH5
z/WJyozYWbmnNAkxDkY9gQOTUjpmzzCzeVyWu7oI6tg5CDtIg1O1R+fO/KET2eY9
vWqYfytvj/F3nItliO372ompawSgFj3z3ySzexyf3QaImlZeOSMiqjghPJ14coRf
0+lUgXxCBMwOMqi2mlk5NaJdHYv/oKZulnfWkjKlq7TzD3y6UXN3gLzCjpy0TX1y
ySwylHPO/5wPoVW+eBkQLUTtXWewMskSOtcqJFcOLBklJDGhF85OrPran0vyE48P
rMgFYpGrwNb6W6Amw6hgDetWEKRZ/snlDALf2s9Hk+re9EGa4CbkOADn2bwunMki
TKxbd9Y4Zo6kJiTOMAj9zfAIt/GRXD39kSuNlY+SFGnpVVJIUioXKrT2dkzAAdPd
Bu35U/2l/8vW6mOyn5nXr7uoUQlHAwRnOBd1vDstpZWSLyA5N8qRhJtvSYFJcJzV
HZmz1cIUJV/dhkkLYF+exZh93pUCC4x8gGBPraFo4TUH/iA8vfvatdOzfbaFniVT
xF4aCDeFKqOWff+ncbH5htBH1ZNpYsStmqImZVLjArrv28F5x5T6ogIw8q9FwH5+
xqGKkJpr5RR1SZNdXl/DRatbDvodyk+vKpMclvyperUzaUb+Tr6jMIS167w0Q4q/
n0oT3qNHuYRxG4yk75TBCCrOdmwRsW7DqBpxbYGCW50xEfdJi2mC6KEdHHbo5njy
rIw12BEuRX08UN0To6xzJIN+BsNjFF4wbgiQ+mpYf4Ki1AAartOUkEPmdHNFoWgU
4F215wqPYFgFgwTDay8dVQXxzlvBpm++wg+8cfbNY6mxyYVCXAynbe01U1DyDfyR
eso3SAlp5CoVRRUyIda5C0sPpkWDWCHJ6J970IH5tFkn1DB4hTKdb+LrcSnbNwm7
u8AXX0fkI4hRoJljOVIRBehlwqoWI6ps7nOuUY/3kIDGSP5vCT1jD45jvxnPvPCl
3KOVJ+cJVeAINz2HDqWp5bd80n4txIJpmuflfWDrpgBhKnJg2lparGA8EKzkZiyJ
Z4O/XlryVjaiyg5owt91I86Hfply14BPR0qaIBIdpwWUL8ORqdSrdWqGIKYmXGpH
VqBqzO5oFx1xTB1lI1v3zemxpCwuB+U3PGyHSJneZSEzclApOI6TFBp2I8fsKjFF
ccwMCVUvWC8Lar7t1zBy9XsZjdfTmTfGZvVtEJyTnhivRRuHoZ9lHEdjxSmSvRqu
XWAsWzEKUZgUqwwE0rXqd7dsYzkML786inviS6v4BdM+ZvoCm6CerVIHF2p4ZKbl
b6l4/dSg9R1HFV0ZKA8Wgx3U5tYNam0QbgA96HoDZUaujJ7uc0tpuHjlpRbJ6USS
hflK0j0nzCBJpm5S7WHXwH3EUmzvkRPsu4glomMeESdXwgbVaGW3ngqj+y8eXI6A
aGieNa6NksLEcEx/yMwBKx8LbLqMNYaBAfYSHqOvwxYkdrU9CycUg2slwopsYqd8
j7Wq+00HNAF2aRyEFpC73VZavDPPhNtAhC5KH64cyg5vxPuhH5brh5cKoV5iFKU5
KvelVomx6tiwq+ECtBLmMepTAYP1W6EeH7okVqWdQM4MuXk3UAIM1NL216niBAZN
suF7K90RB8SPVEncwZOpiRD6Mx4EiGMHGSD2dnDJDuPd49SqvldYwS4HK08jaU4y
8VLIV+ftL9jH1RJS5tfwo0PZhOulHAmT6y8M7x/hp5W9uhiIiBG9zwxf49EJCJWG
2VSwBMGrwEfrXuyeiNHmKpTyZ6OYQHA0JllFDtO9vPXDipaUh9b9lHKfOd4e8GNn
OnqiafZ6Lon+wvWOU8xKaJ8G82rDh+2wtCyPvc8hipJFcSq4P9izTW9uRyY5mQB7
5o+79RwPidYImLfSB8o8hVKItuFZosACObz3NLJl4Q6/At3iQC8aYmMXcIACuKpu
T8Sparfdwe52O2uf6xoFkrC8YZX/4fiIpykiNDm4ChiCDEqsz2RAwCk0VPv6uTV9
DxSvyK1Y6KwGicgpf/x35yWfYGbC9L6IYLmcaKq/P0/LKuJ0ypWFT1su+OBE5u8j
MDH38OHnU1b4VCpsrrcvjLa3VI+AMk9dMEGDCb38FLf9Qsx/Nlf6HgFenPxh1upV
FDjKUGV9MER0ZySZ3bqX94v8iWeDibqJznwFJSXa+mt9VGY6ThOE7dBdTWkGxFqq
ICoQZdOVZ4EYasD0+syzN+wqRfv0lk41L7k7RLE8eYzlm/VZPCdGhRPRj/IEKLVW
4OthA/RNHr0vKEDoUb4/xG3c5kWUHNLdgLjmYIimxmHKDAewJYn1vQQosypjDLDm
ggTZ7cwF0ukNketBqxkN9xohcSC7O8dC0Nv18jpcAAj59+IWytQEvE8jZeFXgvEM
d4rbGqghxhowzF84ekKYrSo3y35EyvYGZD261eaM464hjT6SXZH+sTYMaFt5jUjp
6pLUJatnvf/t4cpLoAcjazU9U3cdZ7CxHwgnkf1dKoqR2cW1SIIhzxkQ0Qtj2qcJ
ORx0f2TQdRxy4/NDynYQlcxz2PuHD7z7RVsJByC00zevFAjInLneJ31tYDuTNEFf
PiqB4cUe7L7y5bLekAcd0auJC7h6SJR8wBDk3N2jJ02syGmOiMX1BlJnd6cncz8w
CWBonXn6N8yPJywnchusz9+PMSHw/nE5wXmpPBaq/YPIhQ8ziD2pQCGFV0RIJbeL
QoAMW0YDaIcgoaDmuOsSEXFusY07lTdlsblHrPWsiuKkK+JRtkIIRdt2mjeuRpR+
Wp0vmwdpNb5zb15IzPuzXANQzuHYA9eh3JqtePXvnqgQEbBNLbOvdb61cpKELbsK
DuN1H4iMHWhfsgxfEAoY1XU2T3jYrN3Hyg6Gekb16o66lnGE+KDWJGdU2RFPe1Dr
m5MsAhoCAN4xt7hWLnPEev6X1wUN8bUgrpK7Qgj1gFDr/dGUu21gMBnBpovkWX0f
8fI98I/jJetbRP1JH+lFf5tficSr+WsqPoUbvLgwlk69EJRTyW6MqOGhswNJaGeM
SBi1J1syUSKIBoIBMgQXJYUcMoYV8/v2ma/hU8dBcjSAF9tPZJ4Got0iMcGwwsKw
u3n2xnpNhb1TfJD7C4gR1HQs0Wsls6474nVX/A8Yakj2su0q3NmvFxVIoy43jk++
Y1V7sI7bEpW+b0pV9QjH600kzgnbLFiLSihZWOJS/QKo8SnSV1cHmf552p9/k4wm
raydGkLgL4lsja+B016owm6wy2ySufAEq157OrnyL/rC4uD5FNAFBMS/nYxfhnMN
zRigp0+OJexA8LnkQeu7OlsPv/Gbh+vR6KWRFt3WQQsY3WkYa0D6TZTYamzry5hd
rdvvMtETBWmcF5/F/5jqtr2v2MNffv3j/SDektc3ey/2e8JtMyIYsr/Iu90wKIMO
XGvn+g9qaWCXfW0c6Vd2I6c32y/tHVKzkJpBvbVL0AhF6SYl9wJTVGkAP4LixjQs
PF0j33R9v6gkRhxE188MqX39094rSJi6QtnEf+NCS7B+WSg1vJKUkQxgO/ixhD0s
jAjT18JUW4C8N4ht6My25V+kSALhJ60w9FRV4EC48awdGqBK7Koy3VsNc6QzGIO0
CierLoCyl3WZh4NnvcMH2XelJo5T4zjfZmRr5iwm3gQ70nnehIjnRp3lDRJ2eHKb
4YeMin6fgQ+VcogPYBIkUDf9mgOm0LStpzZ+mrPfAI8W87yEQ2z85dIh9vjCBycd
Ooaqxl0cfx/FEzGFEiMIuisC5wR4UHyJcem/ZZvkuVsFeFXuDBGAlbBL0STScg/o
fti2TfFPFt3UQIUf34uHga5D/rO0yLCjQRy510s7Uj8EPrRVd4qmYpQ1YTaUFBxB
WosEFIuUR19kVvMhHBaj25JzBYixdmp8JHZCuEG+HurcDr0XH28lQyptJrxONDFQ
GVbXMZeQ2sU6bOxUNqZpVUXYQWABjWL8CZp1IBOGQtq7MM333oHlaFkoep7+rukG
jKtPfYQA/UNPuqWDH1JJtDrvEoRAuTRc17T9s2h5JtPB6fN9hWFBmRgrGNVHuIng
TqJEeK5V3Zy+E7qT6FxFATV6WcLd6YtRJrmCdR2dAUBn5YIPWDzSDXWlFn9kD52n
flbJKCs2P9HEMedLrVBs8lfJ9h2OaiqUABlpW8LcHP4KeHI1PhMAmBHTse8Ddskx
soNbytCbfJnIubI4HYVE+6dnH4L8VGCvT8cPB5U+1RdhR2Z6HLQQm9S5h0BFp9/i
nTQDqJLPuWmKxQ3XWUsLZprMWg5+xmfL2+D1U8Bthw7k/Xyh59H3XL4XCirkucxJ
N1ZcbJW0NtYVBjeqs2nJI2185DWntceuc2OVSX9hUxe/GSLtIkz5V2J1ZiBa6nLM
1b03ukWzyXnZkialAeO9hyE/zZYliPLe67SUQ2Opv0OwWLsHMU/0V9h7Uod3yoPq
+RPPBwtmb424dxzkfVnWgWksnaMSXfogZoflPfp1sveVrNfZdW8qXONGq1F4BNE5
kx6PgpuCRVMs7qJWiLhD81PvGTD1DZONkkBCZyJFAeu8r8mpVgrZmyH3SNHTkerb
hR8GPvjUphK3qdEhqxlpUpO0lTmEz/fwkCCTHRZw2yLjW6Pqm5n83Jwm9jTZhwwO
aQ5QNLw9TFapCOCsJwzqd5unsAtCrVzy+O9Wp3/h7qHyU+eykogtWdd3otSMDw4o
qFhXVmA3JuS2mqIicrLDGjtlbV6QDb459E6/0EhuWU1ZkBlJ85zFD+ldQzXVfgP5
dNBe1JWiMvday6J0wYCOP+v84vDN9w4vEWcQMiyRLmjwL0L0PNNK/WbcvnU9r5/V
FpB7Ol1NdC+StHRTMZB2ltiNyXkMiKvPvGMsF7SXZVYbAth1MsSpM5ph8uhnTWlg
FnDyZBr7NeZFpRw2fWA2j5w+O/3uxLggrz6UI1Jc/G2qJzZgUlTo310WZIswTzUS
lHZJs7kqgtH5u1cbRwzAv24EU30JXthB6zG2bMihjtbIwdnmXlwQEQLIuTyO4DdD
nfJBRK6Nit5YJF32wjeldR/81CDMNzHrtn/xv8j1tljztEkM7ivGes80CK/cUxSn
LB3i5Ttep1idQt0GQLcOa5bEAR7Ws9rnOJUND1E4Ohmp/sSZeZXvSQaEBzRAcACe
0vzNoygdcD97MvUwFnZp4ks0zbVu45RNy9CKsefCcpvENlCOUXqu8+KWVkr4AO71
eHWgVzfBT+QWD3ucf2Ah4ybkDmNxRG2LGLmXNdvbE3KCPsHgLTEZGdZlJn6L/4Ou
u3WGONpmyxDFzXV0xllyGHPiTBxx3lhToUXStDhgkaKnd4Eg1jso2sqObAgsb68Z
aQMKEqmiXDP4wW4YHjUAUbXXa2f/o99zsqhSYzBowfZDeKi0wnbqV0FLSce+lByt
mQ+5W5aHwQ4tHQmDvZPB5m4VsP0jFN9QNfDmVYxEgezxrzba/QxoXc/6oCNqkAsT
bLMsSVc4UNS9h7R0jz+MvI4H+JceYe6QLb01ARnfWFO1e3sOAoG/4i//W5Y3MHeg
FEA81VlOe8qE4G21GCUeBC00Y+fDRU+Ob49LyiBk2xBokdlUUqmefHpa6j+jGKZa
9KkPxI1YKj76qqTpNtgn7I8prBqV42axu+kVfUZhd5npupQDUXevMNYT7tXRUGIs
q6+uedEelED5Fzq/SE6Rcq+ooZz4QCnYzxMLVwVzOq4+XI+q4liThb3TzXdTW4ks
R+SUV+YUrXfrds0lHkwKfBiWLTlN8ORZ2bcwL+s2lMKZAyon6Dmhd3+kBGVfa05z
F1dRZQ2PxK83OfHNR9EGSjH8G8AefrgVZX4v2J3PTuJE3rjcM6+XBQKULM0HPweg
C2hfI0qfQIbciHH2rbfYiISgJbEmHrSFp90e+97BAA/x4U8zRv5Pk4ASjqXHl99v
yiCrXcbINiQFLtZecEAAUokeokM/4148MVEIignSX/WRJRFUuGECvtTR5VnmzOAV
mPWI7qV6rHOr2pLLFwTFm5vFZmfo/sPtGTJbOoQaA2PBUDrFFEAoCY+lF+zZCnKo
epUSqqf9LZOAFFaBLQif9jxyc3VMLD1A7BjlNX0EllKSYJKswvoLIXcjq6kGt6G7
CH3rQs9XJsoqdihvx1CtbfHjoGpWkbux3voSzx8sVCVgyjtOgseFuPPuPe9jo7JO
KzF3/blYZDZLpY34cW5UUAB3m905T9bXWW4IPmod/NRU1IT6pgfgXZcK2jA0irh7
BR824nhdTb8Yj/aR9kLLKvTbPjzOPnJRGDV+/XKgIDceDgPCYSn4xYuA4GmjXMYa
NO78bGAdnlfEq919cGd8ivfG1IkyXNfeZCfNMp8lG2TuOCMwSYsq026yuDnJzz9S
18adtZYbEZnSNUupaB0+bWGN6vql/6oAbsHjjso8tvl8WA2pwZ5jH40vh2XBm29/
/x92SKbKQ/ewNVuOHuDPgUTuXhN9POWQQfDFjU1n8nsvu4Xl2hvHhZW/l2Nhreby
Jv79LJ2WnSKFFT7yEcLMQJmScDyovT98ndum5FrTliWpLabBgzroWSDuPMyIPkRR
5Ppx9++bBD0JaMd83ShxFprWsAMWKX0eXqXugtFGmwty9+ncEi56rSyJyDHNvJWY
vfQbr/w9M3IOZag6gB9pq8GFL6efkQIWrgeHB0ZtUia0lOUDqh53KN+Euobf8ynj
EN379FDwi4/nS+MZi8HoBhI2s8X7GRw1biQzSKV9IEjhZprzYLscEzYkXLZE3Jfg
k+q3MLjesCkY3VKi5xojQKir42XJNEKr/f1oEycrJRlcCezpcA+o1r+O3bh0YoVE
JSQAlFbX7nQofM2XaXfLwiyk8udmCuRmENk3k1qOUgPGj+ZRCWUT27B6DW3uiOrm
+JGM7W+OjuE8oK81xrarfW6OCXFg+M8q0ru+6VAI2N8mEw4tycEeMxJ9MnFZcfHR
4A5MmMcSflJwzjFpFm9fu5eCIsCCkSZytTqPVZ7jf6gPrOdmzWQ9oppXhM1qmsYz
sd6EkQuz5dkQhswHV8MPCbySeTQQtzTUE4dmg9pjUdm/BelTG8M7fh2IxudLxBJQ
OUdd4ZF9BuFMY+lBNVG6VpG3l/jdLolJK8NuROOY6iTIrdB/XGKfbZz5reShRLYb
9vZjqmPSN2r5Ob9QyxzLmLsdsxqwLNeiXeR/IpuXs2MGm0E7fzFRyGUs+VhdVJEZ
pH6XBIV/AcgdgxCFitZi9QC9KuOM9k7wYyJTD4XGIMawtyUqg7kpivYkYGuMlPJ5
Zy/P795WiYE58wftc2v/tn0EJt5MDwEK+5AMT12oUr15Q7G842HXcthdXgffB4SZ
9C4g8Sj5yN3dAmkD/MwprY5ADgdnKfZvky1358rqDLRXx4SJyiEDul88nmNQs4BY
cFW24b1JC6Wc4NzZviY6HnqFSoJqHvKY1oewpUlTBvR6oAK1AvhOLA2x87CBQQFF
qLvXtNAq4Tt0XxN2TGqINHwi9k6w1xrMrCDLfa8tjhwGy+V77rBNBaoiiebCRixl
b8pzfPG0EsRwlZiI7/Z0mTz4UMtkOyErQVZbFq0gW9ZGTHe8lgs9UavkI9j4XiHX
HDbMCVPAZAnu08wbvu5f1LwXgZmnptuJNqdUY2z+QsB/Bpf031Yg0ZIDGD7y6zcl
MGrzk8eY06O64k9GAvV+A0YZ7sRPv9X3w4tgm7LrSrABp2faHer9xoVXcqV1pZm0
bIChq0NfDP1FDxsMatxa7a9xUMGPJOHHLoCJXhLmEVfcf/BEMZGnlAmA+nGOLV+h
QpGOwc+VRrnLDn/Ckk/IscoLTJXhld7LW27Lu2TiutaKbL2HxK8ikwD1JnVesRHV
Cfw0we9pAL/KndzbxmL0Q4kwq4axfSYyp2DddmkJBCkF6bpxw0EMo38fwyX83fMj
nLUyrXqIgQUnxWjINf1lKbPYWF+LS5U/suwZ0tZArD8R59nccpvKPTcTzna8gmvS
o+2Hxk/YuroMx/MEcP2WEYnQtypHfTc+DrRwhLgvRhht5n1/Q+yf1HVoNowvi3Q9
YgM0xfdt2KDdxz1bskTg03dAuM+7hwbFZfI1Qt6FiOduQqUR4H/Zc2yBtMsqnJrJ
bJ5U7asBRGZt78wAVA2HWLDmbOx0IaCxJvvGiv13jLmfPurt91WHF60ZLmTCkRea
EaQnJlzZkfXenv+pYyLDAFjIhkHskriFEvY/3UYWwIXnFxDo9Bjz/udrPIErO6bo
QKFuwDPSr/DqCQovSSNKHaY/MOrK/BSG2ppKE8YAMckxDsI8ydDeAlATnKehEfru
MAt+pGXzvpWRvEuMK2bZJV4Ej1t9tWIquGdBfLmE1y97XiW/pKKPZgDG69AMquLy
3M/Fsu1vyYp1mYUj6sDHD9pvwilW3DjJWrOQZYt6JvzaT6/bccbwYorv+qQUphEx
gfvFS+HOwT3WyjdPXsRi6X2V8N+nzKk8Ur/jU9QR7GWi1PxPYz8l20zDgr0Prb5O
0gfNMout5e2grExxnynrr3iqswg+IPEPykc9Q/Mchxt23x5G/hSsPsLr8y1EY3qK
ZRlRffjPrGmiXQX/zvhipRTetWeP8NSli61oNvxq41jQ3vUFtw6MCaWGGMNOFAzc
3x5kJIBEEp0OfqrskPJAsQLLxM+AeD/W/wiXD/MNZyVTm0PcYkqzesXZ/E/ivwCS
vHSgtgGygAHJtkVjbN+VnKR+TKSjJmlPJEko2m2675sPlxnOVMMQTZ1s7NZ3o5QU
5ELtoeMDMrOmNyZHDXLDyOOXFm+maPPVoHNuk+5Sb+pajhc2aKN+4gF5UkBXSPZv
cmkjgBFwRM55DGFSI9aDlz4seV177iDBBIhcmIRqYInX8nFnQiMD+Epb+eZW+mja
3RcyHDkOKwp7P7qctMHqa13I0FV6UmYtNB+O8Y0+Y/vEOAVWHfQaKNtUirSOM9ef
NDBw6oEbuCKo9W9oZ0Ta4p+0C7L71rtrk4c7bmcA4nUemWe9cn/ZTxfY4+14F+vM
wfmrJc3qMPS417+Vxjtou8CMkl0s4I018RBTEuWuiidZAF+i8vFMS4IK007rbcYz
lqeJKwsBc+rCz3jkyBb0DFZO0yVltSKS07v/4JjX0eCxtP+L5s6TyQ7dKPu+0PvT
9XMzjqfRmkZTBoJNuxZzvdODvVF5fDQOL5eF46lIxG5qPV4WFDD5WxQOtlCvOoKJ
7FTGWDztu+qR7RzpQgf+j5qmLyk1HcGHsm5MOh5LlGuFE8jAN/8gfE1QXrv4nNX6
wF/w2YsE876uxBILaSpY00/x1AFOk1D93n2L2vg2bWSnTrC7wn8l+7pFB8Vlm9Pw
yE4c7QOGxJPScsAgeViaH10nfQQCzpqCrQTsdyO8D0pFFGuPFn46cPFT8deF0ugk
ukXKAC1lIHbulsyd9gicEVCLelBHggQ92C0FIJMqz3PgPGbTm+hzzQALNiXR2jgO
IusPfsepEUyKf8BZ2zL10KTnf8aOEzqdO4+nLpBdGgTSbCGu+oM/KL/2wj9JDj5P
zdie2tPyx7L1jNAamk4biy2hhJPuH3wJN0HKAYLH9+rga9n7riNQpB9CnI5pY00d
33xyU0F0jT4SBthTxgLuLQ==
`protect END_PROTECTED
