`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4ztrSw1OE0tqlmoajVExlUXtcTm0zW03YY7YCfSfaz6GPhKEpvVe3H+W5v5mG9t6
MVmMHEVVPmHttXbtQjqRab5H/BX+8TuigyvnsHpEzBGTWYbk9C8riQHspby/dsJc
d76c7/xYRcJ51ECWZUg+Le9/TdX2wK4Cwl63lAKhSuIcfxKnRfKRa2s8BaOsKSVN
g7kCztdK6zjY28EvZExAJ12UQAQW0LF+qcuTcgA+rdCPJJjcpr74eMbQJzGrWHg7
QMhfabBN8ornip9ah6hAx4BwhXu05zLJpJrQz+ZlHNQsmD0UKATLimoT00Uww9Th
aeUlDOY06XyiDyClaey2eb1TC2qrBgE/J8i5XORgCx+zJq7vxE7KhQVcZmkk0xT2
St6looBkawI+YJybT61D7Zn6RgcEylox+BfijbnA7472ot74SHZwCdTSP1Ta8Mcr
OjY9OvIGuIpjzfkh6ZpkM36IeUGLJ+SFO5b60JCGz76eG8HirLcSuP9j1Us7+SYh
KVUU+zFe4I9HB9Xqx10SeVlAe2t3IaJpi/Ro7YVx4HQzgUTa4NCspkIHYOODGvJL
XniHQEj5ezLKBCTTzCKjfTLsA8O3Db8YOv3tnanPjNaOsHE2r7feOm9X8725dxPD
kW3/18kzT9srZGJDagyRE1LzVklujLxs+4bCNfZdOvL5yZ3Os3taU7IkLe6I94kB
8Koxzj5r5nBl+uBESYSgxf8qPpTJO5MIMSCJ+jZxEn0jXaqIKj8XYZF+n39yE9Ym
9h8MD6oviLWJGoTA3/7+5eOiLAhBMySF7QsDyjKUFGlSO4gVQewBd0MgLHWyVEGJ
Ovml65zjH6fGR2akZxKd3vBT2tgwTzRDBaMFD+UopKDtHHSCY5xM90xD4WJZOsq3
mOYvUhJk02PKXqxGIWoupe3N1984x28ysBAfOdbjsv4Dh+v+i4fw9c7DmOTtcREa
fv0XKBhr2NItEHBVxE23vlPlUYG2y+fGwb0ZsUhNrkWiTloQHYLfgofotPQ0j9LR
+nRLHkcQSTG+3jvMDqi61K++FMQXkJQD7V4L/HD8VwncFydKugTuEsy8vLA887JL
rG/gvoAhPDgUg3DfVche1GoCwLpuDLeszzhb8ZfGxsvd1F7SrSbTxSR/dMfkOGOg
DxOI1WJD0QjP2lteSLl4hxdIV6zaK2zmZC6q0TyIOEciE7P2bZW/38Gqt1tCJSAq
rOhcqF/praY56Kb9zpUsj0onYjAm/wf2umnCy0SkL8KP3elHnu47RtKuLDeH+E49
wH6P27A4F35hQMffdYCC5oOQGdbEdZLVlj563eHsBnRx4ePT99Z21kDMCzT8pzan
tOXQwSWv05Dp/kfvDhP8UPhYfzcTUNs86Tz0A1tqgZRpOznIeb3dfK/WQZZKskqX
sTJGRkzuIg1rVVZjjvOsTe70f74xjRYdsmg67Me0a40qHXeSkTgQHa9Z3vnOWSCD
nZBh3hV5+wN1lKLfCrpHN95WWlZOBu9eQYnSPQ2bCzWBi2xAHqg3ZE2B5bAlTu5v
dUhjiT+gwnNCqZGDq1YriUIYPjx9RCuoqtzeIh7gKvEzs6yNyrx/F9w82vJbi0Wb
XbO55H1AnNm9z6AGkh0Mt2B+gp09ob1UC0lMfxZkYqw/s5FZPDN1J45yVuTfmDAO
PyX32XgzAmXMUrYuHAaaVvdsJoHioP+6kZLV6eNu9o8RcNPvFo28X/qDPPXfSeOR
A+zePH5kBu6GKp8/rRR2Bb61174WIvRp3n2uEZW+IaIK8HLIVg1GydDMCc+D45I1
P7CoM8l+TNblFHSWgtMZE+PIdxLx8RLBYup0jE8Yul4gFj2KzTBCmkze14mTkV3F
0inR5ge1bhcJ/4GYLLfiuPhTZY9eha2OPwzHUgIusRc0yYbbWSbY6N6dCwHj/9zt
++S15iogvZSQso8onoCFDwlRkYQ18SR/YsuHs7hUt+/blD/ljkXC0Q3oRZkTS+gK
5jumUGqINJj4eYI6NOT82mE6XdKvW5sIgIWSPwbkXQmt4NPWpeQYK39iXHWnzvsf
Vlhn2VRe6HiNruEORO6mMWz+Xp36KRIi1v1qc7NwnKsNlsxlt6lT+/cfmTbByn1t
dpKJCvA104pXgz8lXr9BWBSvxcmbIPlNJVUCsYGF1HU0hvUrka6gYkpvG+AKd+W1
KRSxFjCCHmidikl8/hFF1LB94Prqpam6ocUDw+FFGH/0G621XaPv+IDKKPmdDE1c
PQ/PmMX+sVRdXGMIHLi2P3HpSY8gg9pxeY/Kwf1wm/Ls3aYvoaq4dZGOiQ9AMp0w
T0SJI7OEF0sTJa11QxMAPh7iZVhggcICmLq2gHknVCklilALFONMIJFW2yM135cl
qpCr447e49TsR3p3KDtKuIdkDxia4r0qbW1P0klkTB5btAWfJRh/FkjU0Mau0R03
U6c/+YRsj9J9aWoFDJYqwW3zn0xao8oO+AIZHo/HP1lQbXA9UqH1QWTcvq2aVKgU
gE9sVhWlfDT4PALROwvgd0SCbairnTVdlmqSygic5G6sTJYW8zs4UQ5BEFoLRx7O
1gG76uOr/2MPJkN4tYXS7yOU7QNMJ9/qaLUSdn9m3F7XctGk/+PioVT3UqbZMLhI
FyEVxMoNl7HkmxR4Xg4C/VevcBYKMN/609xnV6csbiXQjEI8+m39zyu/6pnyyzFU
MWyn9bNRUGe24hJf0NXSoplyCPy/LyJQsn8FSd3ThFflDc/gNzS3TPuU6auN/sim
wdCPyHXCjBZAxwpMxJ/u8KOoTkYRfALNfejlYNEz4SRUVhRtEgjHcn3Wh+kHddF9
MiepIrCiegwhyjokLFfYho0+psm7Qh6uxwkQab+Zr0frPzwMgNzNLobgH+Bj5zWo
weR4jfWIBPU/ILXnWDhLprzULaHw7Z6ZxSr55kVqmgFamQtmuFCOs6qWiirar+7h
tAQiBDREWf37wmouvrstCJokjn4Qs8Zm+A7xYPKZSr2FXj9kon3hU++6FF72WNUW
a8vSLXHWSOXuO1LTOd/nsbohPdxCTW1pAyBShaY4wbLnjJlWm8G67nxUqUuJPu3h
BpqILv8Cr8HWH0BQnZJr8zqOjZ6+Q6Xh+R2tcbsr/agCWsQMvGE//xa/jbYRRI5Y
P8rJFudRafM1dqBfWwtefVa7evM21adEuughEwg8Y7Td6wm5qSR9QyTgCdvd+GdU
zRVMVxIpexdL80TYsR5och7MOi3gCJi7Ns4lk29PUWPTlCEpDX/aIVG9g8UvZ4NM
yLmnDsQm3zOocn//8iAsVw/AucjzIxqfwLNkqIQXNxGWUeGwAdtw104k9Xfmng+o
EvqUSFYiiNz3J2EZ3U/dHZYJmgdpgeAc3hwDg21Z8TqnL3oni+ZUttkn+9Y9KgZQ
j7a5YwrgjiRQOvPZMeY49g1BtEcDzmHHqBtjm6Cwy2OEY8Fv79dtQaIQf65VMrq9
bGRSM9eszyJHlVGwL/qn1uZ2rHwKDxtUMq/XaZbT58GzXdYQheJB2GjRCXH9q5CZ
wadbguvvam2swJnR77pyP3Nxuk2tpg3DLPUddToMIH/24lFOwhL79c7fwDQAZ702
crOU0PqYBabw3udKaRdl5O2VMRIAs/Y29R9uqOSXhxB5Klm6ijgZNSMOxGKkQPjo
PzrOCxKREKjSiquoV5tsRypb8KqtU/mskxW5Yl7UXuYLFBrgV/HL5jFC9gW8LClU
k7eeQSvrdGb3r8EEaIRqvrl+IzJ2RGEPPyf5EfYjWMwWQRL+4DUQVzxj2h8j2LCD
XE4qXILsJuJAWXkznk+Uip6PN1uT039MLMi9VNh13FHz16wfaK0qsdhYmAqr0Xvs
9xbgx583TyjMbd6/JsdKyesp5kUb06ND/m7Y/nygErZKj8rbuiy3/dA6eXHJ7yPJ
ws/M01xNNXtqYwejya/CkVS8UXarB5hy71yrQy5Q3ep+N2DehxmP7omXUa2rYvlY
wknPeclgxL6t7nUAsPE2/Hq6w8Tnr1uKU2NLOL6Kxjf8wvTqcFGL+1v/06gJSDu+
AdldaD4+ZG8KNSX4px3/5CCoCevFkJGN91rdzIWxwFsKRWTeF9GXTbvOKNWc+0Mz
XCrJDnYXUc1MN3tbv1gN0n3hzXBeTGm4w1ACKN3qhBNS4t/NWQg9/mpIjx+e+pit
S6BW+tJvGmXLzNNjvSbdqE5H40PguKSaUsLryxLblROgk5hoAsRvynR/mOXmciiG
urKp4X7Kzv0KP0qLS13puc+Tf67l6Yr7GfAnG+jRctNU2Cenx+iOgGi/pBtRiiTE
xgRU2vSXUJyq11dVRsq7me6BGKxaJW3m6rpP40ExLpgAh29wJYAoWUhf5TwzEauf
sbeNaiURoQmbaaCY7OHba7Zbz/WqoRB6+Jlbo5VsFg5fePNao1n53pLkpWbbk8d4
x31xuBB1/pXqWSVoSzo4LJpOM38F+i0foQ5FsJYW7o4N7Xku/1q4Y3v7f5ijUzfk
5Xn3WE/WPia99CAWz2dsMCQifRs/KEHuvqpzcuDDAn76s5Ja7AfCM4iUsY+ND5OY
hjQLZ2TEkL4iTFtZEe+6ZYxi5BtTprkZ8Tkmn2i80MRdGTd24KSy/aSskv0S2ia+
ec6E1jxs0lJFrb/xVf0z3Fu3mz9il1sJE4uSylpbuH540xPyAT8UFVEKnQ8FMDOE
mTipWYakj5vupBV0iLeoYA==
`protect END_PROTECTED
