`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4uvcQPepsim+9RQ0S+gFj6DSZCBodX07iUdg5HLKcRabjAfeyA2/a5cBKjwzxkze
X+7De6EponaKmVb8wnGNILw/UCYrV0P7LfT7IEvfD+piQnBPKZIMfokFgVnLC1l6
/9CjKZ4mU4XWMZNW97bVikUCoUZYob6wsTGdZVc7+9J2eyCcDOZqskyCIyc377Pa
6U9M4Ieeg49x+3KYy0JS6o1rHzwujyAdJZl2MUsGC+3fyeOS3fbK2xwutXj0GoSe
b1Fi9sXePfmz9Jc6u81PTXY7X0G0Sb01vgcL0z+jFqgtYT1y+5ji+/ahLoY9ShRu
TiQUP59YFYPsi3s4Mxg0nVzmI43k3KmJLEGnGrFYE1t08vducj/jAnggKpXa9no6
7TiqCpdBU+jsZn2dFyxOS8mCSgtkycJD7JPR90J/6dy4amRkYd+HBBJfNH50P0+G
sBEH9ol/7V/wRztu4Y3ubA==
`protect END_PROTECTED
