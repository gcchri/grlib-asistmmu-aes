`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FUhLqTtKbcHeNsn88knEa5nLPIge7ub0+EogA6lzs66GJPwbCwJBC2tw4sUQk149
LpZ0X8/HzhQs3+X1AihezFmJrq1/mGpjodSq4yXIouKAK6h+5OpWuRtTXJ42luTF
PbkKdBD33RJ8Dxsz18KFucRtGJ3nf6A9NmvYPFNTbNmKWK04reO1uFrq8wQjHdvp
dhxKKsV5Sgcw0ksRFRxDtxVQNJZ+MRQb41LkjROFLaAJqcqvWfB3aPMt3vruhA+D
XykWxiquSjmDGVHM2SymJ5oGu+avZSSgLfbwIfvytj2wS3Jr3/XDT6unXfK9d3RZ
skoSsGG1NN7YbLIKoTKQ98nx6DX3F99gNDn4xOEduhmzzKZT3dUCCAND6mNJbr/2
kOzo0JjuXv6kN874EwFT0OW5BjS/nskAxM91RlPTPiC0V4jgip5v19jyWHkQNSt/
HbvOarb9JKZCMsfNmacbKBhfjCShb4CywmbkrKyxSZ6drUp5d3XsSVutlUGpRIw/
zAFVKwajM8yYEckCGDriEcbvn2WL/379q9Ov1XoK6mglGSM8bBlw2YZ0yB5JiG6w
sHgdihG0IdKiLxzj8HC7tQ==
`protect END_PROTECTED
