`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QHAbDTyTwzKfOnvThkxiKbFocV2/KFUkkEz9PIQR/YNuqWr76pz7OPV9NxdR3rXo
4KOiAHYWVEc36DZ4oWLoXAexTdjsLuGyvusSMkdm6szYo//vuexhIxFPRcVF/ZNN
sfI1mBtRBJnWd2GPqNmQWEcq/diuR0d4v5ioSj7Zp4fANFvW7XTlNLJPg71lxG3L
YXSpZ+g167gm8AAQS8NT0uXkdxkUePjU2pygQwCyXBo4x/VifhTO61sJIGlptCwF
XWvvXdaRudbcIGalAkgv0J3t+nM67+Hw8VmKlh1QmU3hG4bLTpTSXX8ZPN5RI9L3
4ru6sHVkOR2BbgT9ufk/YyyWzZh1XaFKvLYPZ28hVdQuLcHB5UHg2EkfwoY3cvU/
KBrU3H0AqUOtqyY8EpfvaOvicQqorj95Z/5FZGpWv8mQKrqu82nMHxNHxIJVeg7V
Knm5c9xqKiFO3NeUmwDZBXNI0HJSSA0t6xpOm4JOQXuNgRhkPKriTpsRrtTqzzYB
Le7EjnRV9IOPKez8Bhaz5vQ4CCAk2OlVl+h6z+OqpbqGQ1XMmvz4CVo89Qk8yYRz
SlN3FK/Ck051Kw1Hx4UIog==
`protect END_PROTECTED
