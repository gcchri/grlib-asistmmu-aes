`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AH2p61lkpHQM+HPBLuTWGnvqA8/8XygVGQPaRq6Ld7jJRdlj4pJfaBpIDELhLuz4
hgS5QUGPPQh4Bx28O2zqgtefV2OR/TG6kirQW/z03SpoaDmWlvlcocFuDIV5fR7W
33Rke28oPOekEsZlY52ALd+fgcyNzNLI3M2roDLHxZMKuqmUkuMoOniw9RIvVFAP
cPKs93s7N5YnzyUVfKpdE8WrohDSt95WUQN27V7WvS1W/fMt08gr7N+CLSlTer/M
BI9M3Fr2akPhTOC9SGdhOOXkyr5YNauN5JRkm/zI1kN0h23ZyaxtTm2E2qQsAam7
mz+oquABpVrHPxDF6bq2WV2itO3N0aZeZcaCoy6//nnHjet7uyecAlQf1hG4Qk+N
+dbqkepUZ6oh608S9LlFFvqk5W1niWWRAJQ0SBLrjbfz1z/I+a4P/oUF4G27KrTS
FhsQrBl0e3Hu2xNOtHS5Cmeh5QA45qGKLUHmviEedn35fPzpe+D+RZYVQKQDi0o6
`protect END_PROTECTED
