`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/j0DXrkTO9B2pcTci7dy8oikS7d6TerzwCt9UFh7upYN4MBGvxuiahBUr8BaoF0J
ea8nFqZXCOof9bgbKvgpgQSdSVlU+NmKo3v1UKHiG1CgCVG9dbsYp5A/IHXbEGeW
4gIV4ymhZEAcqsJbqMlVjJyedAzIIHzeQT92+ztGwppG2nBTUbWS3FQYGuxXtplb
vH+RRSM3ySbtHr9gGBr6Yoaygjw7hPzzVzSqxUdv8qfEj8XIOa7SBK1DlcXFq2n7
yQAjWyI9s86mu+aVXpzg06ww9t8nL6kX2gwLkLlmBlw5S1/E3h1lDNG9L96B+dUX
vWdyEXRb2+3ZLtGAlWE+04+wlvdGdekfzvdSNKhuJ3dVNEK75I2/nhkyHyPW1y7T
IWvCd6/G8L7AZWMmOasrqiLl6z6GoHKqPafxuh7954UEwWUL8TvikvveoxlvKxhY
MFE8s6JiGBXKyMgu9WgXisc9wAW9T0sEbT3GXVgq4dkk5JXc2vxQnLeIKi1RbHrf
WXcqzWZYrIBkJQl4+Jt3DsQJG8xaVqeOvUFkd2ecA7yvXxLqucAYY/0u9WkDufvQ
a7N6gQgDMbsEzUrwAlPBAwLzvg2iXScM04nojxIYjYCMT4O1STfZmEv9sa+81YEC
UGiOcWnm+ECvEuvCo+WM+T/h+KQUISgpac+p+UvdB7eMbFasetouEWA+BMQowCps
+xEcDjW07/5e3oCL96lrZJu+2wbYryK0jqFOVgkzAj3VzCBxjBiqyn6LuDK27gbS
Z1gBExad8SxG6qA2hagmCnMTtJ6GsmoOB1zY2v1DorNYk3pzdkLLIQkp/uKLHdj7
aiE6xYKva6PU6Iq3KhrpjDLprq3crLRfeiuIHSci3OtGMHN4OpqXEZVsNAQMm3mU
WCgz3jhRYQSkohCnErFfh86x9+lK/KHlDQ4WC4PyIhTLlOfWhj7BGwmd7/4ZDA/S
WhSrSkEb8T+YmugLPTD1PRRmInon7L34+JxMEnhxAtrH6f1m+fCo20LTUSjVsDbs
EtvtL70viovlpZpyZMVlMUnTc+K/DKNnbCIzGVI7CYSSAhdKVOQeNOYqO9LadFuU
qHjQ626Em6ea/rgbBMerHR++60CcWBi4N8KUm1FgAZ5sEX6OnOnwyVCw1r7flp5N
n3auF0MivgSAD6OoLyLxCUN2LXFXpPpkm82PanfHd9rLQIeKNPiYsyCehrgxS6/Q
ORcCJ8mUmq7CUz30i9zAHnx2D3S5bnAloppp3OBKzdZkrcle3+JyzhcI25qFGSyi
scSKX4vK2uAejbD8dpPy2S008Xsq5LLVkDG2MqNxnKBpI4S1Np3QK8qI4p80pRoD
JBLSCUabe5kxsKczkU3yyebtz+rQsreqnTmp1cyVr+N7xBiY/1ub/JMzCtVbylB3
Q7wsVzrNHkRmYffOLpZaQzjRpvsP3v/hl5XRQVyR12J/ZgkBrlAKqUyncTw+HWzh
kJSHWteKX8mlLXM55gVm0ps01iP+DZEcJU+eQV4TW/RMv98T9Mny/alEyiSn8FaK
ouDFv0Q44wGVHoqX+Ak6K5gtOKSTOxuGm25vLB/E3WkLMPdaMbaJqQuxsYzt8qp1
QPqNCXPJ4RYGzITvjDXe7LHiJjAoVy1pNGDGg71HmG/DbEbWF3Nrh4UetFyvAhgh
FJ84oBaVyJfO9nhoOoDCZBmcNRz61bcjYSutJ7aNxTpGqdmJJBd2dejxOB/oGg/U
DS/JmX5p5I2j7BCtGeRi/WPm01u+y5IkyJtPNcyoLLNmOS4O6tQJhckvSZ1ZXvqf
V2PMILBcNRKbM6EYbRhwDWPL7z4TRiV31YIcc0H2RK+JVNBQiYxjJmBXI29csxCN
X8Q3fTOPe6qGzcljiULqCZpBDncTgqmxOLHBvDr9iX5SYIBUFcK+giyCWkherQeM
67RYy0dJvYo78yVJm96YKplpTNAUBBGiuUssMSYPxasiIZ+wM1yBC4F64iKt+da3
ytuqLA6wS2hlFOteeELDEiyis0xHPuLr6u67RrCBmY5gKUKPu3OBwWeAr+vArVXw
U3zfDGZWtxldTAOpZZGQjz9ZaSEH74oZz9qNOSTT3M196av3ZQNc91HE3uq0Aby9
DlyQOaoAC9bnNBQLwmiPpD+r4XPhC+uBCClMaSwlO4LT/YS0S90zg6R0XV6aqBOM
+7Y9w9ByxkMRGN/AS0DP/9w7OdFeV1FzGCItlClQkzS9qKyVQOh9u7b0Qf4QPyqc
got1Duuf/f6CvEzhKJfg0j2yx9bPZ79f2uRaPTCAkyw9QVvgLnBsGTTWmkkedmYx
ECb4sEiBSzINYVRL9UC+vLADj6WOQxfmzdlu3ZQMdouILXZRRPwvwt+8ml7d0kHM
UNH63g5P3xt8DFjjGGyD8/UwmiXKLvJrgi3y7xqVtDD3OxLwPLcL3tNC/cPzkGCR
KwDCARU17d/HM4YK30FXb7Lnor27c92+GBxMc9vH5ld6jJ44cC52WufVSiILhJKe
iqjZO4Xk8C5Bs8HcdiIYURGaueTchPROE76NJLfAcorUjNDLPdTIluTObMRDReny
YOGK93YTGkojeuoTOiGQo4zolbtvAwzycjFDkgo1FwhCFqABw9wwb6lPwIR7flQy
EFmnT6cxzLWgw6H3UOPcdFZG6UsGEK8rCx7wnfSE+hBOniS7HT4Tf1Y4Cd6/szpe
WfMIB3Dd0kgxFsmwyTa/tHcYNHz50SaX03TtbFr3yQ+HXge/X0l/QjD6SYkPykM5
kpBjw+M6UiuIOeuGjbAarIsr0l1s0tfpSKIYyleFjUl3PXo3pbCWLjEsilK33xKQ
PbJbelOBnhKbcJSHr1z8DfOF2sWZX8oDLKkFSsV/Ta5UOuQfgdGapbp05zTEb1Ce
Q+tU8bEJ1aQvt97PqbMKeAoZfBNPki4cacSlB3uI+kFPPymWUDMp7yaTYHTgPEPi
3Csg32V+Wcae6Goz3LrqmbLkpBXhRYAiQHSPeUwRbzexrlg6iHa6HqYidPC4dV4V
w+aYUExUB49DVaurAyAJZpp4bGHn+6XtVcPnOuWWKVhgniAL275YZGeWpYn17hYt
cjk1N6WUUNaM2LSRF4HH/rW18akrCs9RqzbdefOIoCPR6gY3YTiN0hJ8PZfin6jG
9JfWGutP261MWB4GsfzpPgyo5wXowM8UpuXcmLdLVjiePaAOqnkn8D/3V/FMj3Ft
/ln7feaU9B2/q3fxrTWiow7u70aibS8p/Yh/CmCnSsaaI3yyFrICA/YZGqhGn8/s
xQt0dw1qm6gEEo5FAwm5MME76zuy9A177kqTWH9r/+8fIBx+1j9CBiVchTeyGxVz
3fZQt8i7j96D9wwfQVuNQCs73pceD19hAf/XL/aOgVb1a/qE2FBJs2Aalh9lZMTP
Z+BWb7wado6LH4kKkEr6KQFvXKbLeuK+dZjxoXDpx1pGKkAnYFWJHK/Yj15Mf64d
D+zAQUAVy56dYqtB61SD4PJoHejo99uruFFcHzu8v+0byhpCz1X3Ky5SO4NWZiK9
oGHYxt0dBPwjWzIQQyimPKSZgUNq/lhdk+Z51KGU1pS8g9VygEA7EIEyvPlVsP/5
kzXk21a81i6DZP5OT4yhsjbkAukNCKwgVy8sQAWAEpdFacv7DZo4tk4rVL4yLByK
A3IixlDdBmOiaZHBvZKVVDADyY1pIvCbkA+9xNn3gmGd+q1C5c1UaRvTKtEZPkOP
RLZFrYN+uP6+SjtzztvGqIuuJtV0zlOFI63XdPjF2E0P1fzEBZxbFI9MY7J6mRvg
7zYK0PRbqEvJbhFB473JVjl6gcY7ECjdCHkxZZOeUe+d2+ZpHPDw5FNSS2kO807c
Bau04mRVkhW0mm+gZXW4hr2CqFokwsr6PyMX9c0zdNfjUX+vex+UJfBBiMsCuOFo
mt4ndhP9FgpzCsGvDl02peXMncSXDNbl2SDqVdxadRU=
`protect END_PROTECTED
