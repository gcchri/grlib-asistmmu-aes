`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cjX+jVow0wLC88j3ISWzVmp1bhrcVqir9tB5tadCmXn4aY6dsHxdaAwp0xpXv3x0
JD+CQwb+8dZvLMHeHdkANhBBvikY70DgiYLIUBcENTGkf1MIAbkNW5eJ2ee0XS/4
c7QTcPw03CHLGAorOiBCx7sZGdAGTEQdnPCD7pqsg27iQwnyhkp0YQmo6T3Mk9PX
yycbXcs5MJ+mc3FT6cNria5CgK4M4C1t4As3Lj/gjUK0GmpvHITQWIf9xQ+MqoHh
kyEfC8y4+1QfKphYBWnCrCQya18buVrQbNfZtJ3tH/sT6pKsaUyKubdzyu5lhfca
+mYcgcLmwMurWRD9Anh2zfkQ5iHq87vcQUe71ApdFZCMwzW0goaskBfhMwmc0yIm
/aEzZ9mjqUmTjpYwTbT6TYdghxZQMWgdfTZdaMR/lPN7nsHBVIlE/cuK0FYzkZI/
kT+XVZJTXKrrR0g0ZJCy5YxoIkDQDPHHSS71j1iiy7x+OvEwbAzyANzuKXextDV8
xbO3MGq/9gNwnca84HxpVsRidFbsys1Q5gkoPT6iZwnTvHkAo9Jz2n0E2y4WvnO3
L0dMRmam1rZJZz7EdCL7Q9b7wrf00yu3qlcldasZpLrSibA9xuDFKC/oxv11gu4n
vxmk27sJnX33lLTTgmOKwW2BPnxSbpdIn+Py6u0HuVjjNzlbiqs8ZqCrRayUOm2V
tcLq1JpOYOfD0ngF2wFdXKxa/sFZ/EFzAGmOedI4prbEGErHNVNBZdd9r1vPuwHH
j7VjNUtU1d2YIT+yunW0cw==
`protect END_PROTECTED
