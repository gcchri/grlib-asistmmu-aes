`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F7ujA9tmUdpMHMwtrqluUKnQjc1cq329hjH7WitoNiW1b/bKa6RCqJXeQoX3wSbk
g7h/Hq4dQL/o82WcpFNSEUOOeE3VBrN6Cr3JMppADrgDibT8SZxfc/eJg56IcR/U
t4YQ3qNMQmvs3JrbsW9/rTOmodkf4THWdEwBbXXKc1UYORmH1vY5Awxc9dQ+Hg3u
sKRWOsMEGO+z/DnxFFE/zLbT8zUbcyzmCmFaPKlIordZEo7arGIxJws+EApMUJQV
TpoNJi+HwwC8D46iUE9t83zOvn+ii8Qjl0Kjhy5JtUe/QsgOKqSfMSqp5Bsw0+PI
gOe3RtUl7/+fpLwSd3BI2TBuF7K+gX0CIUOoMXuGMlIw7Uy1+FAfRRp6aFFqaTdq
yNrqG3arI18vNRDTVuoUWw==
`protect END_PROTECTED
