`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TxUp913D7DdkHeCgR0eu4SHI4f4kETUXJD4tuf43uwvZQZhX5CtFPROLI7KanT3U
pGwjksw8CqwHfmhuB8VWXuQh/Zt5Tg49pIACuHAlsskczPBbTiE09xQ4o5nntJbx
wBgwF9ujm1P4UKMb3Mzp5iUEpNEorJyyQAQtcpj/VFGN9sFbiHD5H3fSxBFixXKi
/DyvT+7rYMlAm7aMpTf9MlCy1bMBVTQErlqvyJ2O604Cc3/Afo5ojk17vOwq/DHs
/DpXNCzCNYkeT4GN9/OB4XisBwMzW5olUODOKIHhN557jwhfPDsS0RG27fC5hdai
E2Byn6Inj5bxriZpOXvA5nt1cLYBy0g8MywT+9OLbUITXKAOuZ4jQOKeCYXhuMKk
iv1ee3sOKLqTS4PnKEaDK2PR6kyMcEX1hboa9k02G+rhiwzTr2f9AjpVF8C2BxXn
yVYpz1xJEk9OUPLQvElcRLd/EcCIw7PN/d1H8xKvEUAUiaDFQqnfNaDyvtf9Jdv+
474tOuF1Jf4ly8JxqdymlVvuh8tCY+XEOVs6+Zbi/5UxHYJpBTirYYQwB0qBXZgd
aK3hwUT59OE3cZFWkjWabw==
`protect END_PROTECTED
