`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hRh+TUKZVF8HGTVRiRrK6xu9ehcgMp0m/KS7nJth0TQUL0Vkw6pQdOmCf+8VNOur
WCWRVcUh+o6nHUf2bjkNLH8lvMIQ1zAXpefKrOPyolwDhQXNq5pYbroUV8zmw6/H
aMMKv6IAhvoOhvWAMnv264I+vtwr4o8EL2mlCFxuXlPSfnXXQTSFhpLQwK15DY8f
jDQsgHL15DXb7y25TUC6Kf+DKnUikYQLXF1gDLl6YTi3RijknXwdP2eNg+mqvh5Q
oSWCW1I0XrPwxxCj3PWuJopQC67uJzrYyQS2a9vo5ITyIQqfJlCQd1aNFbSG0x/j
LEFf49srNDKf1tESTHR6xGDK5DF/j5oIgJdSgzikt/w17g4dqePlFvBtOijHqy0v
eTjdpX0a5K8TlULUQrn5xIZHGF/89Zc/0nMzVp9hYAhlD0+hqA3CqnVheLtIY460
2dzXf7xcuxPwaGeb0Hw6NFEpFSI7noUJzdoeFMeHqRNZUFgNPGPKB7qEpLKpaw4F
41cP2btnyNnQll17swged6I6jsMsCK2VJdwZy+0ktXNRlEfWe4Ice5jy1982v2Wv
VdRMPNvkeQ4sf5BQ5jQzYA==
`protect END_PROTECTED
