`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bT387BpZysFEDiQsxWSzp2OFHzFEtE80g99Ihsx14CFZuaWN4ZH4Kf7jEj0jSmwY
5Atn5vsQwa5u4gU8OyG7OlK9d8L9RrEBgNJyjxPFYOvn2qryQwkGNpb9R3q/LJcW
tYo9nyijnM4da1ZzVE5hUto/Hkyv39nyU2sXpInwqaBAtHKmuBdadzLDT3m0Bsat
PSSVe+DqUGHa8A+AR5QTueBwo4YceGTw+NLLLuaoZkG1DCOkVfwc2AWMfSwsEnpB
NFDfdxD8QFRRfj48mDcX7k3ThxqN0IsMszqjcVsIKprRHHRRt3XSaqcBenipwsdQ
oVCgJEWRkc6sK941Tb3nFjnrJjzgR8dLRkmZ5LpXV2g3RqWekKji2QQOvPg7Bhww
0UCWt+F0Na47iBTUje+TDq6maqsaJhLRcBBC5wsDOX3YTQrCGH6M8B92L/bv3d7d
Z/u/fgf9cUShUjNI3oH2ZiGbIIbl7lCB9ebDjCUCJQpTPxo2Ollc87NtyVmCMSNy
cY5Ujx0T34o6nQX8ux/i/ihzWomsF5uDHswKL6yMGv0fWubAoEAdRPpISRNiXQsM
lWQPxXQA7EmJ7V6GuY9Uqn4ibv5NfFIAAwyMgFXa0gKBcEF8pTuG4KzUfibUtF3s
fDOqv/VeoAO2aOT8ifeR94wRvKHtQaeH6/jaNmhGjLh0FdjapeTCMhFUfU01Bs/O
sk0Yi+ahb6qmRmtf1C3+VF89bfuzSulcHuynQl7JPXnkY80kw/cR2fW449R+FgZM
BOe7xCTtfYn5HQ9Rszc8bl6lphvc3FYaqubFyW9QItF3ZWySribquLQ/nn7KplVm
KsNNBwRkxjm1Mi7d4BUS9ErLlzRpP3Mfv0XO1mcqJu/WxMlxNC8TG3xkxSKyNqQ4
6ZwdMIFhb0EDpvnVSNrEIIUoGvm53DFCykmFQO3XHlU/hRVb8O3MikSP4wmoD5xO
`protect END_PROTECTED
