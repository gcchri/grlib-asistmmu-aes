`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
asWVKjJZfVvjOX9ghkS4P+/5pcOa8qjwKoVVOMZUzvOlKEacPU1syDoCYALsB50R
+UwfCiZCTbEtj3y0AglkKP6w0Y0Qwbb+kwYdsufj/LIdDHUrOM9y7CxD1lps+asR
v7SMzx3WVLpd0C4O2udZ7AhrDZEscekOly5P0DE7xpVoDM2HO+rkXuIWs+pGjjwW
1A3bdN3l45BRCTouG+pbXLGhuSdi9EY50zPNqG1FKrOGO4F7FEn3jl4bf/gFHMaC
veD4xUGsTRX5WCdpXtOW3CtV7SXGtwt6t/VR4Pywn6tQVPaoecAVd/kXZ27bdnvu
DmwH3QWGsgntYZTsip+NlqsogwN57UTOkmrMSwikHu4A+nZi8jbMCqz6lT9G8VU8
iBzyta12RgbYhDozDFjfpOX4cU/QPYwI2awXDSDgYvIJZM5KjcMxxx/7V4nhUC7l
0H9o9MxcAkcP6Z0LVJlRE14NkvTh00Wl2Y7GNCjtZvLOIaeyO2gEdBuC1zr9NIeF
Xw6VBQytSaFoTgSBqAk2KDGadrC8rbvYjWNQULE5sh6gilCu4dNoomArYXkAh/Pm
OFaSQA0TLnTT/6WlZUfdjShodEbG3cx6+4u6ltRKCYAk64cdJjaK4ZhsNS/0onLj
PdTsHQLXgwv6pZ8mmIyzQWy3v0/5ucFyfgR9JDYMGg/+VO62PR4G/C5unZZww1vk
lUJeuWm/zW5ouU1mTHfUq81rwYPmv7slUAFSCn5l/4g=
`protect END_PROTECTED
