`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ysMy83HT65w/oQJq8P2Kg2BZ+dB9THwFTM21zTsTaiwKXhyIAoCr5Qj4BsOREOP0
0Lwp844NNz+dlbRNcoF3uC10fFAt4c9qi3f+ECWY+lQoKH9+vQg1rJ4hRvmJGSJp
ZxQP34d07Wa6FSODG0Ml0b7HIG1w0QOhcOm/yApnmMX/F/JjgUZbpyMl7e3jgh9f
8Jx3ZPYj6TWk6pCngq50rv8s/ywwd3QyuUuY5zw3s3MjAH8vY+AdVEgUCXyvx7+M
hTMTiWY2Fw2+HXzjlmDDpncw8qiwZOANShGRtrwBrnbtTuYiG8nAPSUMPDNCqRC5
Y8gDPEn7eAomoFTJ5Vsg2DytV5Uqvtj+UWl9hMJlJLRfhgVTaGrfRsSc9wky2Cvx
ojn9HhfREZDG6IxCGhIp8lq77guPzyDxC3cjMKarIIk=
`protect END_PROTECTED
