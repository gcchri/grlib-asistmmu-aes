`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yiCsErFjFuTpmQjltCsqI30T/HImEd/kgj73vQq/QKzYMNyppn3hrWkJMNINcjTk
+9WPLvqOByGjzg2xLfG40WPaGxkErejTfby3eX6JD9+y9dCekKTU4xVlibeRHGs3
JlBE7e190qJJdTaiIeO5aOmSRiUSSvNRf0zuSzAWFLLY5eoOXRgqaFaUBbEzV6o1
71iQ7FTfhWhPu3fM+Oiw3VJBqtl8JpWdTJoo2ZJD5rmRd0D1BUCx2XW5Nt4wA8vT
j5lj4XVRtGK+7Q7e+fRUH+b1DhM7tRIoXJqUrR0EhRw=
`protect END_PROTECTED
