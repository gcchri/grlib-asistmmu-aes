`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zlJ8Cby5ksBub//VM4/ShSLmusQuFXQceL4qLfeEKbnnbEI5C6krNZKh26AfCuL6
Bbz/C56s+ZjaroP/Ih3sPzcadfXll4qIwepsY8HPFPGzPcaovjMEu6rvyDJ4CHmU
tJF9Txrim5x68eZf5aS3i4xYoUDxGZJ/FYTp+DUoDpH1DhIcUvlliwC9TxYCjgzf
Ckwh2QDLJiHty2kFoFvT6nStM+6Nk37Yb58RoYlNN7+d2QZ4T06SaAOh9YZ4a/ty
JGF3cxxbPpPiwQb9z42z2262POo+uKxfNdNTSIfcNkETfPsY+185YZt3Y0vSW38k
DUO9YcRDcX5OfYi9znqfhj+UP3uDp5U3iGbSswzcdbmzqlvELmHkbduNdH6JtNVQ
ClUb4pDKqXSfe42M5rZ5biZfq8aaPIjdB/oRQfCk2poqU5XEPCYHmOjeWYPCMbSJ
cmaJ8xfnHkfldmG48jIYuf9jK1S2R13/VjLX7TxyFDd8A233tpma9rDSDaZRZXgH
W4zw1gJ3ncLiD351F4N5zcMUudWzmTr9UzZUMUJEw1BsYfRUQMJVi5xuTWQJbd5j
1gn6ibkD7o7VrID5p4DElQ==
`protect END_PROTECTED
