`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vPRWgWp/Hf4hgNRAvFjyGWPEAwD5VDwk7l9vvtm+j1JgBbh5IVTWTvyHdgP1/2Ov
+abp5/3/eX49uLUYFoC2MsPChqIU7PILNXINE1Qpi7ie20HQ/mxsayvOm4z056ik
dhWYkSkDbt5AcZLQKPH19uRlDvW8OsvKPDBoFMZvcuyOOQtoi+T6fBRtpl9lVwUY
4nSl8Q2zL/FUpzCp1p+rs/XTq4T2L4ErRrZUB4keFGFwh0/CSCDD7ScMU9LgGD09
kE6WB8hVz9wM2OBID+klOkSkQqqMjXRLJuh2jbf675aYd2ija6DpKMe3ep3X97YN
GtJp9t4ovD81wFB7SuqBaAfIeyUwhOqeBOelpgMgAM7MZMjRdeALj54DhV8MuCT/
k5t52wTEX6GRjCzlgT5Ch5o96pyH+YDMztOx5wm7ariEC0o2Yl68Gk3ddy0mK66r
eztSpJX3DGUyhBBtJS5JXr0hrrvcsucRPGKiSoLY8me2vNtsWQB2AcZTJ5E/xc3O
arsiW0xO7AboEhbR8vUo0kn42/SX3IhN0KuISCRJp+NkRe6nqyGzmuk16189B5Al
Z13Irdw5s5Q2XjLG2iXeuOMgFfwsO3xxg589KcHEyNp9UL3w33MNDabWqbmBNiDs
hasH5gjoYyD/m11InMaltHhXI9qn+9OIEdtgkvvfyBmkKGLE3sIpejsvmpKwbC4Y
wGOu3DKbSuxLmeb2yTdQf+j1Y99o7bS1+pUs/A1HPLEOgFuzrJJsg10+/zWGt1YE
ZGvckpwCTkHplLl4AAcZD0OiMq4/hQlnCfnQBIUDQfk=
`protect END_PROTECTED
