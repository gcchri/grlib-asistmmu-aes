`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wpg6Js5drOJ91RRff6OhGkS28038HGDL+6DYqZMu8K7YVHrGXfBCcSEbmx4IGWKS
piwo5qLqqFn9P+jPoAzLV/dj8tyuSRrMx3sue0JVYK7CaCMXFBxBMblbGFZsL/dX
LZNavhXzLyz3bC/QPGpIo2R6u4pxpFXIvng7iJMsz5VPW30HdnwOC2sPp8EQngo4
XyVH+yGe1GAEat2fdxN4MUuVt7+ZKCYZXaGN9sf/iTfKm2r69ynkZyZ4JNusPpdb
P83Xq4SQ8oWoW7oAhZn46CsYkj+3l+dyrFScnFMX+rhkmHp0e3VnYrVkDHTeecdA
gSA3ixwKo0NpJkSY6hShSf7Eb/ftSro9wK5uX3Sf+JCuzmJd/3HgBwZery6kR1+M
9N2Eu4Wzv1DZmoSiCOB9K4xm2GmpmGCrE0XKw5gtgwg=
`protect END_PROTECTED
