`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3+Rfoht1secry14RcQGOrHdnmwOBWh/p8U5mYiPQ60xxaDAi2TZchS2S3hVOryLO
iAv7bQ7ktsAF+AVn2rlIqxBx35J9BoFftoNs0UMzcaHcIvvNGoObQSimGmD+Ve3e
DpzSg/QHyZRwkYFcR+zpveaXJyAPeHSi/CL8rOkKsqgLDQocmvRxhH1+y0t0OXzo
HQT21uz53ZOXXPlwg2+SzYtbyb8B9mgm+vezvwl5OuyrrF4/itgXhHUUk26Na4CL
M8ZbWssO3i36TxT1W9Ioy1SZ3REN8wafOCCDdmdfuD5Rks0z7tF9k69kSl6qyuS0
ghK2Vh/nrkrYR3H3yeVqoUX6J0uEtQB63NOS2MJXI7fXRzAd3uYQSjDJUyy10HHf
ZUYTDkKwqQL/srvU2WFhhFh0orInXC6z40T7FvIOxxQ9eRSw3YwWniPNLbBzD8yn
`protect END_PROTECTED
