`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pFmRgXh5zLtj+gfPdNjZpWUusITM3kXLly9uekoo7pAtAAReyOWz6FJoqv4DiR6D
kaMzqsok+AEiYo6Dy/MLsY2j4WBv7sojpW6Yo/eo0OeLYg6HdYlPpCMHPunNppfm
IHhgsj9AA8poNU7yuKheYkF9BVG3E1rIPU2UhOdrEGVH2JlUkrRd1DWhnkfgWsmY
O2obHvmEOLXH6T7LYda/HHHeeTy8w326IXbgoHTRRLiH4MeHuN+HjO6StxsWcdLO
akhQBqb69mPw64cDDMko7KBEk/DSLThga4TUPo/Bd8E=
`protect END_PROTECTED
