`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4VcKeCQeCOa/4BPBBGxyN6NyilEYlAKbWD/+FzqIeTKlu6GrkUMJcH/9BUaiYuW0
8u4pAbgemMm0HBexqz6lOA7MGrG3W903FCo00RuI4FcxiEMIjX9+XuSElvH+4CRO
kWuzEj/g7U0fnK/iuw3Hg5wpMUt7MLU4rSb7fwdMXq59he7WZPKQ3Vs7AYTWJTJm
9ACFE58P0clZuXITU87vMBncjP0uAaPNPa7i2S7sLPqrLYtTrZMZpvB2RRHli8sG
VZVultqNMSfxD++wVLM4cC6WFfpXFkMbOUll8AumwTk=
`protect END_PROTECTED
