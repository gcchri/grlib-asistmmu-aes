`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZC+NI5riVdSnwbzDXmSOQILDMXdwmF/7J0UKKq+CNwXQ9epiI/6I2ZkMb3/pyJ0L
Za22V7x02y7rfdSi0aNhnPAf1ZXowQOI2FvNDDQ7oKg4XtFAVZnapsB7JELocS0s
xMDGfQ9tEOdOzMYuIHHFQ/qWnBMt4IytPmRZVtMciOk5D9wRHyeSFFsBb4YS1bFI
AtYpVlJ0jD6mpJtsnFbZBI8t8LF9LATo4Ya2NUPDnaukiBGc3+/R26ULiV0VCme8
tc668Vvr7SGzk1m2JZPQTTCvrUejgqg+7KUidkm8xn8ZZFENS6pz3bqi3OBjk6DI
I2u95wgvuUrNAzytHXA+DEgMTTpRPr0ju7y0YPITo3qKIWh4DAgCf6Wmqardcri6
YwXxGTA0E86uHsApazV1pGxR8Qe6CicdpoWnXOhIcg/NezsWKa/to+FGXaAm9Qtl
J6hOdsAeOtsjaPvSvZ2EjJ9Gjq6JB8P6Aa6tPaL8zkVpVj/pjYXD27pBuVp8Uy60
E9ANAcutWzExkECxDmxLDA==
`protect END_PROTECTED
