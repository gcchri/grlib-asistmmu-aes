`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ef5O9Fw8rQHlSGTO5B06xjv+BzFlr5jGDPXT+ayyAEgLsjujMpNTx+uZl4lLyzkT
4U9o1eXzvK789cBGw8QkqAX8zy7RgsHiyLHNwTxNDOvYebFK5N83Xi25YDLm6YCK
Rb7XvD1pAwJGCG3ehxxI083HV+Vx7bRPZUzNoCWtXvIJsUNXxjQm4zTgYMKPC/aF
atKV0BF2T7P6b2j1h5zkisEtVuG79e0MVaYu2w+yyHcm7g5SGknZm08um/7p5c5A
FDIy9Kg7MTE/qF/dikpZqAL4zNrk/SBR6Qpqa3YFUcxgF45frOvDIeqyPI3QdHGm
HUu2k1tZvzjwAWTKlpssJX9Wbkv/gUvPp4QC1pnKztE=
`protect END_PROTECTED
