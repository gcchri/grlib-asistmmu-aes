`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z0uv7Z198b2KokialrHacRbc5xRwW3/0aN7GBsrduGv29YkvRtvNAbOUX7pK00Ep
dMoFgeghWpgpkFNF69WPgefM52U/YEeFqr9lvMmfpVevkQi2V2yZTnQlk4Ph8MME
MGt+xocxmDD8pgv9J7UWMrunCG6G+8A0UuXF4RJQPc09ceJy+NdA4uVypatNjoDW
5eeFnpQlMeaSY8IkeUStAVsfVFmRDKDH+670qXEPchS9k+QPHbHJfVopK9rL8TGg
`protect END_PROTECTED
