`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0hrHy7tOU5NlUuturC/MUzCyf57tN7WhEWxE+oqGUiw4FTsasmGUG4oPHukyzApO
r2nIn80Ourdh6IKLUDT8TJTYWmRMNN1O6+L2lK3Wh+Oje9BgaugSQ/Zl4qASpGxU
I3eXQ65EVb3zdgHPXDYRtxn0A1ypWY5JDfupFv798a6fuhSjo+H0Pc7Wt9vAUbsm
bU+vFjwxHvH0QG2igLRZ+C1ffCxMoqZO64R5thHt8MjZyH7A7CFVRnoY/nErSMWo
/1XAfPA/DhSfdlluT//3897+r/bndUuccYx9Uc9DdZvsx1p6pG+6oOOVILu5d6mJ
VVxUxrxsZm8D7b8S0s1L5tf27Vgd7us13moOyg6sBcXhfuyJFDlbQgx2mqvU99wM
BV42MhzZHrWWgQPpwF5GrQ==
`protect END_PROTECTED
