`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tNV0+vrvdiyxH3XloCG4oiK4u/ajfuEQrG640JbcTO6mmfIH3L/IUUMkEdsVICwH
JsL6A0Q376gG/q3Mdiy5ik6+JHLnQK0VvICrjO/atryXYctLqv/M9ud2RxetyMz3
AYCwUotazFxQMC/1XHWsKUKowV756rNmvlOz2b7GdbgTMOmiHx+CZi0hNSIZPfoD
IkXXATlmcA7Th9z/dbiYh8S0CA8k1Tc7t+576qy7hWpYsEy3E1qEqUD6be1OXBnX
TWtEyO0WPoFF/5tj2jLaUUGNvj1xDKryOMF/bxx4k/88Q9eTiPLiA8zlv2CQ21HW
6CaV41X/ann22B5dUi8t1m2sGTjm2eqsXfCKTFSxfPuujVR3VnhlYSKN+BmsjPLL
`protect END_PROTECTED
