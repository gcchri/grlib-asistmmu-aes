`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+j1b/7Gz1nQjaKI1FBwE4OQvpGkpR03W6Ch8Wd5/8H9qyZCNoVHP/gPSJT7Kk8Tj
y8Fu/jmfaHjTvxKDNZXADG6obhljgZ7C+wMhG0YOp5T35kIsZaQ+eLBrqhhBR1a8
Po9C7QWL5TVg6oZ4t7s85YWG5stUiOUS+vBdbOObpNQAMjp1InfoNNZYJBG9QeX0
wuz9WMAL6+/hernM2UC5xqDahh1n/gcJ00/pFDdd30nRmnQ0QxCsP6B6nwFX3g3U
eRM2NOmn0r7RbQ5Y6tMue0K0inqyqW0yYI/ZyeDGeZl3yxnDDjEMDa3Ijx+L8cs6
UhKaQN4uXqh6Jcp/Ra4gLDPGac7cxIXfc1/wQocnOUCRaAKWWUgj6Olz2lRr4Vkg
enNHOuiYCDWbQOdV5/VwZWpuZrz5BfI8OjAKLVsHYu3uC7wMl2DOnJ0UeB7KwgfC
qF5UU+N/FHVFSIpZwqEJrP/Pu4ZTOCtMvQ1LvroJpcPTsuXz1+pQCYYtaUAPJG+c
/43/enFFOaCoASS0/XnszHeBxEYuGBmqRkfFmcUe5i5uuUEoaj52k0Wm7cG6+Cod
ZPqPI4odxdtzFBLPnz6rTCXI/L7Z83Nxa1IvP7xjpXjcWzkBR1fRqCxYd8lRAabG
0CYem8e+j6LNsoFsGFAIhBrnWS/vmeQ/0o8qnK8q76RLMWWbEBTxfeLSdZ4fJ+kg
688vrZWx47Y0u97AgqO5dBQnGmIGuIsoCdhGKN8Utmge4qP3dTthexhHpbWDEZmV
ZwaYZVVewimT6q0Si6CC7dPIjf2P6GKjnBiny9WOBuMMJLJboLPuDIRWDfV5tgA0
mP7YP4h7lkl9jubp+ikRjVLfaX2+Bm+kUTpSMS7qtecVxdnCOSZPPzR7YOUBXHCy
slmxvVyPItResnpxRzfI0tcaFeRorX38KuDQ/wE2Hpj6nF2Kez+UTUok7kqD6wY9
cEEP6CpY5cdgkzIFX8g+4RekhUfcsUKvbXxOq/CQUYgEow9bNoMaCit7E0WYBPUa
z2k20Nc3WB3DlI0qJocF4xQ5g2HxXdSXUWhtBu6HeeIDDmZsHREEf2SN5FMqalfj
YTQqBwwY+Y59V5JJGs/RRrVKBXSdH/VbE0vlNcJhW9MFPXuJkDiUnpzc3BOvesYV
9ufy/g1xqxTYNYoiHKkHnbyWFgQzxZt8FcibhzcSl1ZbGWHXfVrlGSdsndccTX0n
+rmvp8YaFyQLBM2eosnir/DVtxho+x+zKQIFqrYGdQD2ixaiKZ0GJSC4VGg5Jxon
/lI2a7gxehqNhyvp7WxQtIIcFw/1jnI+D1t/8YKOLZSQi02aepNltxHuIpSQ7jjA
4VU+9EPkluznEGhqWs/AJpggI6RdReVMK/OvpZjtRfvaZyEAslnmFrhpRd/DkBxu
8hrZdspb2dsH1m5EzLmtMDe2SIu9nCfIAk5y8EprOJSaQny0MFfzm/5OVjDDpueW
d6w5By3F/ZHdETydj6viY/zSiZIaadaw/zi117sII2VBaiJg/pdpSonyE+bs8U/i
JvBQDUeu5Fy6K/MBSCBX3fF8/dAz0JSJ4cFmDPnAi2e4jfAwB7sE30FIuq/Z4jfw
DuWj/e92/KZbRJkbgwY6e65O7PxA5o1uR3q1SZQlgFa4gmjJ+f+f0VDdIY73uaLz
91+0uJGtT6vfRfILPnDatdiCbyNAjcTYFi4COZAsbfDu72qNxRxHEtMBoS2GcG4X
4sW6n8VncOLLWbT9/PoVfi5gp+KxuabzxX7bAXkwsdwq1d7/UTKFYoiJ00T55gCe
RAETbd1Ca+1W6qpXqfKlokUhECGdsv9pw0uUaOiBs34a+yGgOSkFzNUCqJMl9Db4
tXvJjT9oSRZoe7oLbcTc428WYFb6iP+tCTThzptsL/11wQHQzzjND5MVUnlwqIf+
dzxhgWxgIglOcIOnXWx+drQ/LSAXauMfTpHD00bhBZ+KOZHia6QiMW6805WKZ/Gm
HBrt+Q6csiAVSu2mC1XhcUE59Df0VZwstEPU/HwkYEYmZRQ6NgWFIQL04yTXByef
KJSxJDL2zH2GUT4G1/KAQAjCOOu4kBxye3Cy1D4lP0cYOMFtgK8dbcM64m9rYexj
0cxhJcY2YRytWLgAa8UjSHY7nH7F8Ybt7CpL/qeiVFrn5MMid3CqyZ99qWlRaQWg
uy0M8S4PhJUhZsmU8po3V8VNS8MwxnHnWy1vM2Oyh7V3T81o/yKkMAzXbAQCDVAv
DzULC73fnKFU+u33L4IAsPIu4U2SpH+Mqzo0oFOf02jG9HXdr2Y55xyxnsc+EehF
UE+TX4PXcdpH0ckK6jLwLrnemB4fqM1vJrXs3h9KMF5F0sNbv8uEZqiK11Vco41i
PwcpeK9wvUuO+SGLvK+F4xXgJwL1WH0rQ76NmnSJXeNypBjzpMvxwT6dXkpW14ZA
oG4PWcxSi95TH14YMOoalAMfpf0WZS3Y8MR8G+BzTN2HKmrCNbAFsl6InMdMlzn2
7DkHE4OpTMI4RCfUIc0c6BmA+S7jeVLgkOyLZKpONxpkWvPBrQ0c8Y4GOsrag9Qm
UWZTv+4+V6DuN8IPYfx9pilS+NALcCKvxg2aTDq6DWMVMYfwfEVCO2qQfsj+Brsl
alh/0EZUEpgraGY+br1TLuDBkdacJHdIsnpStIU5n69r3nq0II5LNFmSUvdsuuuA
/6OfFQluqDb2/MsDkZOvTEKX1Oh2tUunHhzMj/7kzXGVeQW8vv6kRrhKDk5zBPbW
drybqH14Nb2Gz1RT2MtMhCsu6VAdLQgmquBrziuslz/nhY2bXIGR6zsg+h9eYIcI
afyk/4iEdK81/AVMG6UJKter5hxKLqTGU0j3YEww+9qTLYSQKzCVo2l5YIe9kXVr
zmc92lZ/5y2OTB5yBlYriTm1mbAXYz28muF9c5lpzPNZLW87ZmTi+k6f00Of2PY3
Z1do5+ww0a7iY3rHm9gx3Y7w7ibMBQlkvins6IgFyk2+lUeZMIanhR4ACbs6jyeQ
ioeWoIaqp8nNGgdq6ty1J1LBEfHZwsJIVOB/51vnoU+UzI0CuWYF8jjZdg7VtR13
tH+D2VU0nEoFNbmV57UUTsuKHcKhgKfVO48C5pZF52+3EwCdhLeBRO5oN5LsTg+J
xEMtf3JK/gvRUkgQPDIUB7HWw5VkIjRV3oe+wg/d5nmeip5MWtiNMGY0xn0mWaUN
mgl9J9xRuubohhKm1LPuXnLh+JtYGRnnSwK15oGL4AgmSOLoo/Q7ehb2GJBOb2Y5
aFu332zeLYCsnE1KA2w0z1OsI98JhIXyZ3WqKapLgvhi5/E/KGPe21CehamCAxj4
VpsmOaloOR8To489hm/oruIYftu0EUFdc8iJtlNbmY+gqeVPEU1YHPYZYnHrFaSa
00jyg7qeELQWjACtrGph4nAMlVkTkvIePBh0r23f8nidA95hyLG6ClI7VMdy8y7i
bCmQBEVZdsmPf/THq+TC7zjN8BMyCw0Xgatt8eGkUAtcO9CTrA8XP0+GQkUzrv2g
BDtFw4F8C341qk53OIoTnGgE0AUoWccBlOD9p3c6rFRviQ01Uf2/vmFnY7QiKEAI
D+86DxxaqJ7ep7atsN1UDl6GQqn2z/VKhsRacjYvP7h+IrX5A4MQUAowranCss0d
aU3OO5rvGfAPk/wNYGobhZ74kbPfyk3jIW18BpwmcH8jVcSglmVlR/enUADyTKyS
sdM2TXl+lEK0I6ubvSWmjBE9cTisaYMCvTP7qb62D/N7PCvUK9iZjm+I82aOIep+
bFYbNaGNAeRhM2KoNTIQbjafwZejDAm8xPjv1vfwPX+N9C1UR8TvEiavCnc4Sjxw
yNTsm+WR6FhoD02BlHvl+dXxi0XuFIoVpBFLSghZG04=
`protect END_PROTECTED
