`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ugpY9OxUQn538JNzCIg5sx5mXDS0Arn1j9wy7qFw2kx5iNTekgBQPAEamTdS07S
K7rqztSp7exytUIUv2bJGPgiWMjWVBZmsYsDZdR5uYz+JtXTMSpfUrdE0+J3WzTm
blgQXMbONUqW/E0eRIKD4xqjs4yKgXq+to8lnDzbRe88C3ybvaYavUg2gNEmvD9v
Yvz586hHXVr2tjfGDHchNzxzveF9DLgCbxisDEblCu8qpBSpACMNFLjRS92XRVM5
2n4L/WWmj2sf5zxuZYLxtXa2tQAiXi4nyoc8l5MkTh1IC8WeLWB3+TdwwiARaOJ6
Alqn+vDQS6TzbNWn3nx5dH4YRpSvkQ18X2PIwo7qh5HEPlI/L52KrFBIrylBl+L+
yf8Ar8iyekhSzteY+XfIYepn0AGqEFeyOQoYEQR0ton/HWv9Am/DnU5m1mQGCdqZ
uck5sjlWGzWU3Y+N2N+oHPuDaFtkPSW4qFjK/vUrgWSX9U2i44Z1bpOGmzrZZM4q
4Y2Xd9okYFPrSK18kXmRvX56FpE2fPeFcgZrIjbQJWY0OrfvCmo3mu72GAnOEpHW
7qwcfCJcGsjL5rlAc3lNrsU6zHe0MiXPWBeCcD8yQIFobWYnI8qfjlY8ZJ8U4vOH
zlhhV6yNCpVqLZOadMY7sIGcjxq0jM6d2lZLemWRrbApznrXhiGp4rwaOfDgt1FE
hROSrTCsQFbhQIMVYO1E9fDaJtnQfAavxl6356X4dDLJOCbvwk+JK00fEB7eYEJ7
VnFC6bvzpBUACijNkTW9PWIWjbt0Nnb9OOfVLiRyukSKEXYMuomlGpJ7U+DnboJK
cBw+lwrehThFUzDfB4YymnZXkvCjP9sj4HB3iXN/I+owZb1jIsSvjmhyrQFBEwVK
bY6Qu762oEJCpsTYDaGHaiXKIiwPwD9xmpabduGs26FvgPMIM+ZmHRN1Ulae0IB5
az3jr6G9/tp0REo+RQ3M1rDhFQP9bSJ4/W5edrWnmluwIl4dbGAF/6x2XW3cNqUL
u6BtEvTWKw5kjp56YAeQKWh195e5wBMC0GSAFTcMBDR3y5EIDgOk+Ta1aRwBNwAu
B83GRkSrB1u7uaeQIHIKcOB6l2kTpo5vnTsj6dQE/uo4Y5FimLcF9WIpl6mstPcs
Ssk+7Gqw7ibRUkcNTR6aDXdIoPIvw9/EwjewA5iovy7eGHti3uZ5/yUWX2aKXNKf
/D+5QXm0byb6OHw7DsIFA6CMby0kMrd/d+nZRy1DQXMpRfZLZm0e3hlNBVkd2pUB
3go3EhUZb3/R8fPeg1qAc0tk78GU9ITRsKKgtDCHcHAwFjpkrpibFbkqaYtATH/5
wpLPhz6UY2j27LmLAMRuqkRJTYNcWL13Wk0yXel8jXS16zHOWxlBMVb8iZ9/nZwp
yCDgZwrrbAi+tUSqR17175B9QRnfZwbiJZ6lQNmmarZFWG6KwMLkWWLOXCdLEvJn
0WX+WmBFBNn5QyfVbE0ng/uhLVvzwGLoglTwgzU9hqgcg9wjS+cCXD2SsU4llf4y
4gu+YcUZlMWrorFPrSXsODgaJSI6somnOG695WDJanwXO8ZYrsFSQgNFf6ViWWK3
wsd9rRNfVcI+CuATIvtKYQgOQf/33criVOS3Si1CH4hzFM/iVkF3mNFhye9uR3Ha
`protect END_PROTECTED
