`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CXAdIvwTw4tmv7DeAuHYtt9oe+Zx/9s68nuO6a7r25sVWeE7tkjgIHE1sDwkaUyG
j6q0kFtU4RfaCbwlyVfFJ0fAmfX/SF6CJzUxD5AtqC/WpEf4IO5R5YerYsgGefyx
e10RhJoNThJQsV8xiiEn4R2Ag43Uc3M2p2Wmk1l6NS83uYb1+B8KM/JXIn4+WrAC
VjDLXc4FMEhTXSOtKdUW+qzoAOybB4C6hMTtNYv5Ox9+QPy6R6wan11V7BBEZVuv
PpdpwnJAXbrrWLbWJNVw8kLqyn2bJaD6/swH6phUU5Uhf4JqyavhPZ1uB0WlJYpI
NpiBWnqKmEehucof4CKfl7nSThkCkxfwJMpFE7aN2f6vZJ1t1yR2cjuDBedFjuZz
1W55G+PRPmGED9bNOv3H7/fWSuY+zTrBNg5CoNWkTlhNyb1oHOMJOxBn14W0GSTW
VKdulPa5/4Ny6rwidaJ1FiEBaWpAcD/YogFmbdU1ofQGbiU9zunftU9tGnsRdgMe
Xy5WEFtlJxfHrvKGJqf6en4eWHctamHSNnXwV6bxzkqyxovierTnAEGcLdTZkvy0
F6u82IxziQZ35V1W7M4QutGueHyAXpTBw+B/uy/3AqDXaxckl2UyzOEVmEmXqmbb
4rXz89uzmA4/u+537rlOTg==
`protect END_PROTECTED
