`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BLxexfZ/tOwN+SdbmRyYzNTkVxB41A0paCSs1IjcFlV+wWi8DwJJS2lgTXLqehJI
5drnoSzYWI4zF1BG/U+fhqDMADs7iHYXY358lBgiXa6XzXONalrqRS0210a7QyLt
Icp9pI30v/xcPtt7LMKODajzAYbRDfHfhWwq+cQJYGHAT6HhtYe77Wtj7UPHMapj
TOfaIm7b+xV79dbOdAzjEVa9ipwCte+I9rCovEyO5WqisO0pztRtiZTj1s+x52ZK
+0fCCO4q1cSNpQH5Lj0oeKARvqwUiRv/UxeY+C9mY4743v+Y/YNRtr0N7FYvzu6R
iRqiBYfS3HuNIFOclIIUJVnZ9sK//sa0B8slhCPRb0w8Sa1sZn64ECVk9nFSgQmM
FpGlSBohzkgDaWI/k9VFO36THvMvx1dNCu3p2egKY9yZb3mO8rAQ36TQzIbuo3ID
f8Fi3ry6Yvjh0z2vVsCosN+COMyC2aO+vIo5vtJ6YS36G25lAW/qIQnMEFIGgrpv
5oKlZAnWaBbx/8gwCjjjNDWt5pE33W/DaNaVd2sZZcrHqkP4xfWtUthEm+15wRS9
l/JK6L5DG/IKKMDkHs6wUzrA4hIorL9435bTwIs1oQAOZXE7LJI7roRkNy1cwOke
HcY7KbzGCY2vxU1pVSS1+K98cfHtMGag1mX3nLu5JURFTS33qHrQiryYBlSA9bMI
`protect END_PROTECTED
