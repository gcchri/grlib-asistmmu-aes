library verilog;
use verilog.vl_types.all;
entity PCIE_2_1_WRAP is
    generic(
        AER_BASE_PTR    : string  := "140";
        AER_CAP_ECRC_CHECK_CAPABLE: string  := "FALSE";
        AER_CAP_ECRC_GEN_CAPABLE: string  := "FALSE";
        AER_CAP_ID      : string  := "0001";
        AER_CAP_MULTIHEADER: string  := "FALSE";
        AER_CAP_NEXTPTR : string  := "178";
        AER_CAP_ON      : string  := "FALSE";
        AER_CAP_OPTIONAL_ERR_SUPPORT: string  := "000000";
        AER_CAP_PERMIT_ROOTERR_UPDATE: string  := "TRUE";
        AER_CAP_VERSION : string  := "2";
        ALLOW_X8_GEN2   : string  := "FALSE";
        BAR0            : string  := "FFFFFF00";
        BAR1            : string  := "FFFF0000";
        BAR2            : string  := "FFFF000C";
        BAR3            : string  := "FFFFFFFF";
        BAR4            : string  := "00000000";
        BAR5            : string  := "00000000";
        CAPABILITIES_PTR: string  := "40";
        CARDBUS_CIS_POINTER: string  := "00000000";
        CFG_ECRC_ERR_CPLSTAT: integer := 0;
        CLASS_CODE      : string  := "000000";
        CMD_INTX_IMPLEMENTED: string  := "TRUE";
        CPL_TIMEOUT_DISABLE_SUPPORTED: string  := "FALSE";
        CPL_TIMEOUT_RANGES_SUPPORTED: string  := "0";
        CRM_MODULE_RSTS : string  := "00";
        DEV_CAP2_ARI_FORWARDING_SUPPORTED: string  := "FALSE";
        DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED: string  := "FALSE";
        DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED: string  := "FALSE";
        DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED: string  := "FALSE";
        DEV_CAP2_CAS128_COMPLETER_SUPPORTED: string  := "FALSE";
        DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED: string  := "FALSE";
        DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED: string  := "FALSE";
        DEV_CAP2_LTR_MECHANISM_SUPPORTED: string  := "FALSE";
        DEV_CAP2_MAX_ENDEND_TLP_PREFIXES: string  := "0";
        DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING: string  := "FALSE";
        DEV_CAP2_TPH_COMPLETER_SUPPORTED: string  := "0";
        DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE: string  := "TRUE";
        DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE: string  := "TRUE";
        DEV_CAP_ENDPOINT_L0S_LATENCY: integer := 0;
        DEV_CAP_ENDPOINT_L1_LATENCY: integer := 0;
        DEV_CAP_EXT_TAG_SUPPORTED: string  := "TRUE";
        DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE: string  := "FALSE";
        DEV_CAP_MAX_PAYLOAD_SUPPORTED: integer := 2;
        DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT: integer := 0;
        DEV_CAP_ROLE_BASED_ERROR: string  := "TRUE";
        DEV_CAP_RSVD_14_12: integer := 0;
        DEV_CAP_RSVD_17_16: integer := 0;
        DEV_CAP_RSVD_31_29: integer := 0;
        DEV_CONTROL_AUX_POWER_SUPPORTED: string  := "FALSE";
        DEV_CONTROL_EXT_TAG_DEFAULT: string  := "FALSE";
        DISABLE_ASPM_L1_TIMER: string  := "FALSE";
        DISABLE_BAR_FILTERING: string  := "FALSE";
        DISABLE_ERR_MSG : string  := "FALSE";
        DISABLE_ID_CHECK: string  := "FALSE";
        DISABLE_LANE_REVERSAL: string  := "FALSE";
        DISABLE_LOCKED_FILTER: string  := "FALSE";
        DISABLE_PPM_FILTER: string  := "FALSE";
        DISABLE_RX_POISONED_RESP: string  := "FALSE";
        DISABLE_RX_TC_FILTER: string  := "FALSE";
        DISABLE_SCRAMBLING: string  := "FALSE";
        DNSTREAM_LINK_NUM: string  := "00";
        DSN_BASE_PTR    : string  := "100";
        DSN_CAP_ID      : string  := "0003";
        DSN_CAP_NEXTPTR : string  := "10C";
        DSN_CAP_ON      : string  := "TRUE";
        DSN_CAP_VERSION : string  := "1";
        ENABLE_MSG_ROUTE: string  := "000";
        ENABLE_RX_TD_ECRC_TRIM: string  := "FALSE";
        ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED: string  := "FALSE";
        ENTER_RVRY_EI_L0: string  := "TRUE";
        EXIT_LOOPBACK_ON_EI: string  := "TRUE";
        EXPANSION_ROM   : string  := "FFFFF001";
        EXT_CFG_CAP_PTR : string  := "3F";
        EXT_CFG_XP_CAP_PTR: string  := "3FF";
        HEADER_TYPE     : string  := "00";
        INFER_EI        : string  := "00";
        INTERRUPT_PIN   : string  := "01";
        INTERRUPT_STAT_AUTO: string  := "TRUE";
        IS_SWITCH       : string  := "FALSE";
        LAST_CONFIG_DWORD: string  := "3FF";
        LINK_CAP_ASPM_OPTIONALITY: string  := "TRUE";
        LINK_CAP_ASPM_SUPPORT: integer := 1;
        LINK_CAP_CLOCK_POWER_MANAGEMENT: string  := "FALSE";
        LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP: string  := "FALSE";
        LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1: integer := 7;
        LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2: integer := 7;
        LINK_CAP_L0S_EXIT_LATENCY_GEN1: integer := 7;
        LINK_CAP_L0S_EXIT_LATENCY_GEN2: integer := 7;
        LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1: integer := 7;
        LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2: integer := 7;
        LINK_CAP_L1_EXIT_LATENCY_GEN1: integer := 7;
        LINK_CAP_L1_EXIT_LATENCY_GEN2: integer := 7;
        LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP: string  := "FALSE";
        LINK_CAP_MAX_LINK_SPEED: string  := "1";
        LINK_CAP_MAX_LINK_WIDTH: string  := "08";
        LINK_CAP_RSVD_23: integer := 0;
        LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE: string  := "FALSE";
        LINK_CONTROL_RCB: integer := 0;
        LINK_CTRL2_DEEMPHASIS: string  := "FALSE";
        LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE: string  := "FALSE";
        LINK_CTRL2_TARGET_LINK_SPEED: string  := "2";
        LINK_STATUS_SLOT_CLOCK_CONFIG: string  := "TRUE";
        LL_ACK_TIMEOUT  : string  := "0000";
        LL_ACK_TIMEOUT_EN: string  := "FALSE";
        LL_ACK_TIMEOUT_FUNC: integer := 0;
        LL_REPLAY_TIMEOUT: string  := "0000";
        LL_REPLAY_TIMEOUT_EN: string  := "FALSE";
        LL_REPLAY_TIMEOUT_FUNC: integer := 0;
        LTSSM_MAX_LINK_WIDTH: string  := "01";
        MPS_FORCE       : string  := "FALSE";
        MSIX_BASE_PTR   : string  := "9C";
        MSIX_CAP_ID     : string  := "11";
        MSIX_CAP_NEXTPTR: string  := "00";
        MSIX_CAP_ON     : string  := "FALSE";
        MSIX_CAP_PBA_BIR: integer := 0;
        MSIX_CAP_PBA_OFFSET: string  := "00000050";
        MSIX_CAP_TABLE_BIR: integer := 0;
        MSIX_CAP_TABLE_OFFSET: string  := "00000040";
        MSIX_CAP_TABLE_SIZE: string  := "000";
        MSI_BASE_PTR    : string  := "48";
        MSI_CAP_64_BIT_ADDR_CAPABLE: string  := "TRUE";
        MSI_CAP_ID      : string  := "05";
        MSI_CAP_MULTIMSGCAP: integer := 0;
        MSI_CAP_MULTIMSG_EXTENSION: integer := 0;
        MSI_CAP_NEXTPTR : string  := "60";
        MSI_CAP_ON      : string  := "FALSE";
        MSI_CAP_PER_VECTOR_MASKING_CAPABLE: string  := "TRUE";
        N_FTS_COMCLK_GEN1: integer := 255;
        N_FTS_COMCLK_GEN2: integer := 255;
        N_FTS_GEN1      : integer := 255;
        N_FTS_GEN2      : integer := 255;
        PCIE_BASE_PTR   : string  := "60";
        PCIE_CAP_CAPABILITY_ID: string  := "10";
        PCIE_CAP_CAPABILITY_VERSION: string  := "2";
        PCIE_CAP_DEVICE_PORT_TYPE: string  := "0";
        PCIE_CAP_NEXTPTR: string  := "9C";
        PCIE_CAP_ON     : string  := "TRUE";
        PCIE_CAP_RSVD_15_14: integer := 0;
        PCIE_CAP_SLOT_IMPLEMENTED: string  := "FALSE";
        PCIE_REVISION   : integer := 2;
        PL_AUTO_CONFIG  : integer := 0;
        PL_FAST_TRAIN   : string  := "FALSE";
        PM_ASPML0S_TIMEOUT: string  := "0000";
        PM_ASPML0S_TIMEOUT_EN: string  := "FALSE";
        PM_ASPML0S_TIMEOUT_FUNC: integer := 0;
        PM_ASPM_FASTEXIT: string  := "FALSE";
        PM_BASE_PTR     : string  := "40";
        PM_CAP_AUXCURRENT: integer := 0;
        PM_CAP_D1SUPPORT: string  := "TRUE";
        PM_CAP_D2SUPPORT: string  := "TRUE";
        PM_CAP_DSI      : string  := "FALSE";
        PM_CAP_ID       : string  := "01";
        PM_CAP_NEXTPTR  : string  := "48";
        PM_CAP_ON       : string  := "TRUE";
        PM_CAP_PMESUPPORT: string  := "0F";
        PM_CAP_PME_CLOCK: string  := "FALSE";
        PM_CAP_RSVD_04  : integer := 0;
        PM_CAP_VERSION  : integer := 3;
        PM_CSR_B2B3     : string  := "FALSE";
        PM_CSR_BPCCEN   : string  := "FALSE";
        PM_CSR_NOSOFTRST: string  := "TRUE";
        PM_DATA0        : string  := "01";
        PM_DATA1        : string  := "01";
        PM_DATA2        : string  := "01";
        PM_DATA3        : string  := "01";
        PM_DATA4        : string  := "01";
        PM_DATA5        : string  := "01";
        PM_DATA6        : string  := "01";
        PM_DATA7        : string  := "01";
        PM_DATA_SCALE0  : string  := "1";
        PM_DATA_SCALE1  : string  := "1";
        PM_DATA_SCALE2  : string  := "1";
        PM_DATA_SCALE3  : string  := "1";
        PM_DATA_SCALE4  : string  := "1";
        PM_DATA_SCALE5  : string  := "1";
        PM_DATA_SCALE6  : string  := "1";
        PM_DATA_SCALE7  : string  := "1";
        PM_MF           : string  := "FALSE";
        RBAR_BASE_PTR   : string  := "178";
        RBAR_CAP_CONTROL_ENCODEDBAR0: string  := "00";
        RBAR_CAP_CONTROL_ENCODEDBAR1: string  := "00";
        RBAR_CAP_CONTROL_ENCODEDBAR2: string  := "00";
        RBAR_CAP_CONTROL_ENCODEDBAR3: string  := "00";
        RBAR_CAP_CONTROL_ENCODEDBAR4: string  := "00";
        RBAR_CAP_CONTROL_ENCODEDBAR5: string  := "00";
        RBAR_CAP_ID     : string  := "0015";
        RBAR_CAP_INDEX0 : string  := "0";
        RBAR_CAP_INDEX1 : string  := "0";
        RBAR_CAP_INDEX2 : string  := "0";
        RBAR_CAP_INDEX3 : string  := "0";
        RBAR_CAP_INDEX4 : string  := "0";
        RBAR_CAP_INDEX5 : string  := "0";
        RBAR_CAP_NEXTPTR: string  := "000";
        RBAR_CAP_ON     : string  := "FALSE";
        RBAR_CAP_SUP0   : string  := "00000000";
        RBAR_CAP_SUP1   : string  := "00000000";
        RBAR_CAP_SUP2   : string  := "00000000";
        RBAR_CAP_SUP3   : string  := "00000000";
        RBAR_CAP_SUP4   : string  := "00000000";
        RBAR_CAP_SUP5   : string  := "00000000";
        RBAR_CAP_VERSION: string  := "1";
        RBAR_NUM        : string  := "1";
        RECRC_CHK       : integer := 0;
        RECRC_CHK_TRIM  : string  := "FALSE";
        ROOT_CAP_CRS_SW_VISIBILITY: string  := "FALSE";
        RP_AUTO_SPD     : string  := "1";
        RP_AUTO_SPD_LOOPCNT: string  := "1F";
        SELECT_DLL_IF   : string  := "FALSE";
        SIM_VERSION     : string  := "1.0";
        SLOT_CAP_ATT_BUTTON_PRESENT: string  := "FALSE";
        SLOT_CAP_ATT_INDICATOR_PRESENT: string  := "FALSE";
        SLOT_CAP_ELEC_INTERLOCK_PRESENT: string  := "FALSE";
        SLOT_CAP_HOTPLUG_CAPABLE: string  := "FALSE";
        SLOT_CAP_HOTPLUG_SURPRISE: string  := "FALSE";
        SLOT_CAP_MRL_SENSOR_PRESENT: string  := "FALSE";
        SLOT_CAP_NO_CMD_COMPLETED_SUPPORT: string  := "FALSE";
        SLOT_CAP_PHYSICAL_SLOT_NUM: string  := "0000";
        SLOT_CAP_POWER_CONTROLLER_PRESENT: string  := "FALSE";
        SLOT_CAP_POWER_INDICATOR_PRESENT: string  := "FALSE";
        SLOT_CAP_SLOT_POWER_LIMIT_SCALE: integer := 0;
        SLOT_CAP_SLOT_POWER_LIMIT_VALUE: string  := "00";
        SPARE_BIT0      : integer := 0;
        SPARE_BIT1      : integer := 0;
        SPARE_BIT2      : integer := 0;
        SPARE_BIT3      : integer := 0;
        SPARE_BIT4      : integer := 0;
        SPARE_BIT5      : integer := 0;
        SPARE_BIT6      : integer := 0;
        SPARE_BIT7      : integer := 0;
        SPARE_BIT8      : integer := 0;
        SPARE_BYTE0     : string  := "00";
        SPARE_BYTE1     : string  := "00";
        SPARE_BYTE2     : string  := "00";
        SPARE_BYTE3     : string  := "00";
        SPARE_WORD0     : string  := "00000000";
        SPARE_WORD1     : string  := "00000000";
        SPARE_WORD2     : string  := "00000000";
        SPARE_WORD3     : string  := "00000000";
        SSL_MESSAGE_AUTO: string  := "FALSE";
        TECRC_EP_INV    : string  := "FALSE";
        TL_RBYPASS      : string  := "FALSE";
        TL_RX_RAM_RADDR_LATENCY: integer := 0;
        TL_RX_RAM_RDATA_LATENCY: integer := 2;
        TL_RX_RAM_WRITE_LATENCY: integer := 0;
        TL_TFC_DISABLE  : string  := "FALSE";
        TL_TX_CHECKS_DISABLE: string  := "FALSE";
        TL_TX_RAM_RADDR_LATENCY: integer := 0;
        TL_TX_RAM_RDATA_LATENCY: integer := 2;
        TL_TX_RAM_WRITE_LATENCY: integer := 0;
        TRN_DW          : string  := "FALSE";
        TRN_NP_FC       : string  := "FALSE";
        UPCONFIG_CAPABLE: string  := "TRUE";
        UPSTREAM_FACING : string  := "TRUE";
        UR_ATOMIC       : string  := "TRUE";
        UR_CFG1         : string  := "TRUE";
        UR_INV_REQ      : string  := "TRUE";
        UR_PRS_RESPONSE : string  := "TRUE";
        USER_CLK2_DIV2  : string  := "FALSE";
        USER_CLK_FREQ   : integer := 3;
        USE_RID_PINS    : string  := "FALSE";
        VC0_CPL_INFINITE: string  := "TRUE";
        VC0_RX_RAM_LIMIT: string  := "03FF";
        VC0_TOTAL_CREDITS_CD: integer := 127;
        VC0_TOTAL_CREDITS_CH: integer := 31;
        VC0_TOTAL_CREDITS_NPD: integer := 24;
        VC0_TOTAL_CREDITS_NPH: integer := 12;
        VC0_TOTAL_CREDITS_PD: integer := 288;
        VC0_TOTAL_CREDITS_PH: integer := 32;
        VC0_TX_LASTPACKET: integer := 31;
        VC_BASE_PTR     : string  := "10C";
        VC_CAP_ID       : string  := "0002";
        VC_CAP_NEXTPTR  : string  := "000";
        VC_CAP_ON       : string  := "FALSE";
        VC_CAP_REJECT_SNOOP_TRANSACTIONS: string  := "FALSE";
        VC_CAP_VERSION  : string  := "1";
        VSEC_BASE_PTR   : string  := "128";
        VSEC_CAP_HDR_ID : string  := "1234";
        VSEC_CAP_HDR_LENGTH: string  := "018";
        VSEC_CAP_HDR_REVISION: string  := "1";
        VSEC_CAP_ID     : string  := "000B";
        VSEC_CAP_IS_LINK_VISIBLE: string  := "TRUE";
        VSEC_CAP_NEXTPTR: string  := "140";
        VSEC_CAP_ON     : string  := "FALSE";
        VSEC_CAP_VERSION: string  := "1"
    );
    port(
        CFGAERECRCCHECKEN: out    vl_logic;
        CFGAERECRCGENEN : out    vl_logic;
        CFGAERROOTERRCORRERRRECEIVED: out    vl_logic;
        CFGAERROOTERRCORRERRREPORTINGEN: out    vl_logic;
        CFGAERROOTERRFATALERRRECEIVED: out    vl_logic;
        CFGAERROOTERRFATALERRREPORTINGEN: out    vl_logic;
        CFGAERROOTERRNONFATALERRRECEIVED: out    vl_logic;
        CFGAERROOTERRNONFATALERRREPORTINGEN: out    vl_logic;
        CFGBRIDGESERREN : out    vl_logic;
        CFGCOMMANDBUSMASTERENABLE: out    vl_logic;
        CFGCOMMANDINTERRUPTDISABLE: out    vl_logic;
        CFGCOMMANDIOENABLE: out    vl_logic;
        CFGCOMMANDMEMENABLE: out    vl_logic;
        CFGCOMMANDSERREN: out    vl_logic;
        CFGDEVCONTROL2ARIFORWARDEN: out    vl_logic;
        CFGDEVCONTROL2ATOMICEGRESSBLOCK: out    vl_logic;
        CFGDEVCONTROL2ATOMICREQUESTEREN: out    vl_logic;
        CFGDEVCONTROL2CPLTIMEOUTDIS: out    vl_logic;
        CFGDEVCONTROL2CPLTIMEOUTVAL: out    vl_logic_vector(3 downto 0);
        CFGDEVCONTROL2IDOCPLEN: out    vl_logic;
        CFGDEVCONTROL2IDOREQEN: out    vl_logic;
        CFGDEVCONTROL2LTREN: out    vl_logic;
        CFGDEVCONTROL2TLPPREFIXBLOCK: out    vl_logic;
        CFGDEVCONTROLAUXPOWEREN: out    vl_logic;
        CFGDEVCONTROLCORRERRREPORTINGEN: out    vl_logic;
        CFGDEVCONTROLENABLERO: out    vl_logic;
        CFGDEVCONTROLEXTTAGEN: out    vl_logic;
        CFGDEVCONTROLFATALERRREPORTINGEN: out    vl_logic;
        CFGDEVCONTROLMAXPAYLOAD: out    vl_logic_vector(2 downto 0);
        CFGDEVCONTROLMAXREADREQ: out    vl_logic_vector(2 downto 0);
        CFGDEVCONTROLNONFATALREPORTINGEN: out    vl_logic;
        CFGDEVCONTROLNOSNOOPEN: out    vl_logic;
        CFGDEVCONTROLPHANTOMEN: out    vl_logic;
        CFGDEVCONTROLURERRREPORTINGEN: out    vl_logic;
        CFGDEVSTATUSCORRERRDETECTED: out    vl_logic;
        CFGDEVSTATUSFATALERRDETECTED: out    vl_logic;
        CFGDEVSTATUSNONFATALERRDETECTED: out    vl_logic;
        CFGDEVSTATUSURDETECTED: out    vl_logic;
        CFGERRAERHEADERLOGSETN: out    vl_logic;
        CFGERRCPLRDYN   : out    vl_logic;
        CFGINTERRUPTDO  : out    vl_logic_vector(7 downto 0);
        CFGINTERRUPTMMENABLE: out    vl_logic_vector(2 downto 0);
        CFGINTERRUPTMSIENABLE: out    vl_logic;
        CFGINTERRUPTMSIXENABLE: out    vl_logic;
        CFGINTERRUPTMSIXFM: out    vl_logic;
        CFGINTERRUPTRDYN: out    vl_logic;
        CFGLINKCONTROLASPMCONTROL: out    vl_logic_vector(1 downto 0);
        CFGLINKCONTROLAUTOBANDWIDTHINTEN: out    vl_logic;
        CFGLINKCONTROLBANDWIDTHINTEN: out    vl_logic;
        CFGLINKCONTROLCLOCKPMEN: out    vl_logic;
        CFGLINKCONTROLCOMMONCLOCK: out    vl_logic;
        CFGLINKCONTROLEXTENDEDSYNC: out    vl_logic;
        CFGLINKCONTROLHWAUTOWIDTHDIS: out    vl_logic;
        CFGLINKCONTROLLINKDISABLE: out    vl_logic;
        CFGLINKCONTROLRCB: out    vl_logic;
        CFGLINKCONTROLRETRAINLINK: out    vl_logic;
        CFGLINKSTATUSAUTOBANDWIDTHSTATUS: out    vl_logic;
        CFGLINKSTATUSBANDWIDTHSTATUS: out    vl_logic;
        CFGLINKSTATUSCURRENTSPEED: out    vl_logic_vector(1 downto 0);
        CFGLINKSTATUSDLLACTIVE: out    vl_logic;
        CFGLINKSTATUSLINKTRAINING: out    vl_logic;
        CFGLINKSTATUSNEGOTIATEDWIDTH: out    vl_logic_vector(3 downto 0);
        CFGMGMTDO       : out    vl_logic_vector(31 downto 0);
        CFGMGMTRDWRDONEN: out    vl_logic;
        CFGMSGDATA      : out    vl_logic_vector(15 downto 0);
        CFGMSGRECEIVED  : out    vl_logic;
        CFGMSGRECEIVEDASSERTINTA: out    vl_logic;
        CFGMSGRECEIVEDASSERTINTB: out    vl_logic;
        CFGMSGRECEIVEDASSERTINTC: out    vl_logic;
        CFGMSGRECEIVEDASSERTINTD: out    vl_logic;
        CFGMSGRECEIVEDDEASSERTINTA: out    vl_logic;
        CFGMSGRECEIVEDDEASSERTINTB: out    vl_logic;
        CFGMSGRECEIVEDDEASSERTINTC: out    vl_logic;
        CFGMSGRECEIVEDDEASSERTINTD: out    vl_logic;
        CFGMSGRECEIVEDERRCOR: out    vl_logic;
        CFGMSGRECEIVEDERRFATAL: out    vl_logic;
        CFGMSGRECEIVEDERRNONFATAL: out    vl_logic;
        CFGMSGRECEIVEDPMASNAK: out    vl_logic;
        CFGMSGRECEIVEDPMETO: out    vl_logic;
        CFGMSGRECEIVEDPMETOACK: out    vl_logic;
        CFGMSGRECEIVEDPMPME: out    vl_logic;
        CFGMSGRECEIVEDSETSLOTPOWERLIMIT: out    vl_logic;
        CFGMSGRECEIVEDUNLOCK: out    vl_logic;
        CFGPCIELINKSTATE: out    vl_logic_vector(2 downto 0);
        CFGPMCSRPMEEN   : out    vl_logic;
        CFGPMCSRPMESTATUS: out    vl_logic;
        CFGPMCSRPOWERSTATE: out    vl_logic_vector(1 downto 0);
        CFGPMRCVASREQL1N: out    vl_logic;
        CFGPMRCVENTERL1N: out    vl_logic;
        CFGPMRCVENTERL23N: out    vl_logic;
        CFGPMRCVREQACKN : out    vl_logic;
        CFGROOTCONTROLPMEINTEN: out    vl_logic;
        CFGROOTCONTROLSYSERRCORRERREN: out    vl_logic;
        CFGROOTCONTROLSYSERRFATALERREN: out    vl_logic;
        CFGROOTCONTROLSYSERRNONFATALERREN: out    vl_logic;
        CFGSLOTCONTROLELECTROMECHILCTLPULSE: out    vl_logic;
        CFGTRANSACTION  : out    vl_logic;
        CFGTRANSACTIONADDR: out    vl_logic_vector(6 downto 0);
        CFGTRANSACTIONTYPE: out    vl_logic;
        CFGVCTCVCMAP    : out    vl_logic_vector(6 downto 0);
        DBGSCLRA        : out    vl_logic;
        DBGSCLRB        : out    vl_logic;
        DBGSCLRC        : out    vl_logic;
        DBGSCLRD        : out    vl_logic;
        DBGSCLRE        : out    vl_logic;
        DBGSCLRF        : out    vl_logic;
        DBGSCLRG        : out    vl_logic;
        DBGSCLRH        : out    vl_logic;
        DBGSCLRI        : out    vl_logic;
        DBGSCLRJ        : out    vl_logic;
        DBGSCLRK        : out    vl_logic;
        DBGVECA         : out    vl_logic_vector(63 downto 0);
        DBGVECB         : out    vl_logic_vector(63 downto 0);
        DBGVECC         : out    vl_logic_vector(11 downto 0);
        DRPDO           : out    vl_logic_vector(15 downto 0);
        DRPRDY          : out    vl_logic;
        LL2BADDLLPERR   : out    vl_logic;
        LL2BADTLPERR    : out    vl_logic;
        LL2LINKSTATUS   : out    vl_logic_vector(4 downto 0);
        LL2PROTOCOLERR  : out    vl_logic;
        LL2RECEIVERERR  : out    vl_logic;
        LL2REPLAYROERR  : out    vl_logic;
        LL2REPLAYTOERR  : out    vl_logic;
        LL2SUSPENDOK    : out    vl_logic;
        LL2TFCINIT1SEQ  : out    vl_logic;
        LL2TFCINIT2SEQ  : out    vl_logic;
        LL2TXIDLE       : out    vl_logic;
        LNKCLKEN        : out    vl_logic;
        MIMRXRADDR      : out    vl_logic_vector(12 downto 0);
        MIMRXREN        : out    vl_logic;
        MIMRXWADDR      : out    vl_logic_vector(12 downto 0);
        MIMRXWDATA      : out    vl_logic_vector(67 downto 0);
        MIMRXWEN        : out    vl_logic;
        MIMTXRADDR      : out    vl_logic_vector(12 downto 0);
        MIMTXREN        : out    vl_logic;
        MIMTXWADDR      : out    vl_logic_vector(12 downto 0);
        MIMTXWDATA      : out    vl_logic_vector(68 downto 0);
        MIMTXWEN        : out    vl_logic;
        PIPERX0POLARITY : out    vl_logic;
        PIPERX1POLARITY : out    vl_logic;
        PIPERX2POLARITY : out    vl_logic;
        PIPERX3POLARITY : out    vl_logic;
        PIPERX4POLARITY : out    vl_logic;
        PIPERX5POLARITY : out    vl_logic;
        PIPERX6POLARITY : out    vl_logic;
        PIPERX7POLARITY : out    vl_logic;
        PIPETX0CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX0COMPLIANCE: out    vl_logic;
        PIPETX0DATA     : out    vl_logic_vector(15 downto 0);
        PIPETX0ELECIDLE : out    vl_logic;
        PIPETX0POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETX1CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX1COMPLIANCE: out    vl_logic;
        PIPETX1DATA     : out    vl_logic_vector(15 downto 0);
        PIPETX1ELECIDLE : out    vl_logic;
        PIPETX1POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETX2CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX2COMPLIANCE: out    vl_logic;
        PIPETX2DATA     : out    vl_logic_vector(15 downto 0);
        PIPETX2ELECIDLE : out    vl_logic;
        PIPETX2POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETX3CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX3COMPLIANCE: out    vl_logic;
        PIPETX3DATA     : out    vl_logic_vector(15 downto 0);
        PIPETX3ELECIDLE : out    vl_logic;
        PIPETX3POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETX4CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX4COMPLIANCE: out    vl_logic;
        PIPETX4DATA     : out    vl_logic_vector(15 downto 0);
        PIPETX4ELECIDLE : out    vl_logic;
        PIPETX4POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETX5CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX5COMPLIANCE: out    vl_logic;
        PIPETX5DATA     : out    vl_logic_vector(15 downto 0);
        PIPETX5ELECIDLE : out    vl_logic;
        PIPETX5POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETX6CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX6COMPLIANCE: out    vl_logic;
        PIPETX6DATA     : out    vl_logic_vector(15 downto 0);
        PIPETX6ELECIDLE : out    vl_logic;
        PIPETX6POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETX7CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX7COMPLIANCE: out    vl_logic;
        PIPETX7DATA     : out    vl_logic_vector(15 downto 0);
        PIPETX7ELECIDLE : out    vl_logic;
        PIPETX7POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETXDEEMPH    : out    vl_logic;
        PIPETXMARGIN    : out    vl_logic_vector(2 downto 0);
        PIPETXRATE      : out    vl_logic;
        PIPETXRCVRDET   : out    vl_logic;
        PIPETXRESET     : out    vl_logic;
        PL2L0REQ        : out    vl_logic;
        PL2LINKUP       : out    vl_logic;
        PL2RECEIVERERR  : out    vl_logic;
        PL2RECOVERY     : out    vl_logic;
        PL2RXELECIDLE   : out    vl_logic;
        PL2RXPMSTATE    : out    vl_logic_vector(1 downto 0);
        PL2SUSPENDOK    : out    vl_logic;
        PLDBGVEC        : out    vl_logic_vector(11 downto 0);
        PLDIRECTEDCHANGEDONE: out    vl_logic;
        PLINITIALLINKWIDTH: out    vl_logic_vector(2 downto 0);
        PLLANEREVERSALMODE: out    vl_logic_vector(1 downto 0);
        PLLINKGEN2CAP   : out    vl_logic;
        PLLINKPARTNERGEN2SUPPORTED: out    vl_logic;
        PLLINKUPCFGCAP  : out    vl_logic;
        PLLTSSMSTATE    : out    vl_logic_vector(5 downto 0);
        PLPHYLNKUPN     : out    vl_logic;
        PLRECEIVEDHOTRST: out    vl_logic;
        PLRXPMSTATE     : out    vl_logic_vector(1 downto 0);
        PLSELLNKRATE    : out    vl_logic;
        PLSELLNKWIDTH   : out    vl_logic_vector(1 downto 0);
        PLTXPMSTATE     : out    vl_logic_vector(2 downto 0);
        RECEIVEDFUNCLVLRSTN: out    vl_logic;
        TL2ASPMSUSPENDCREDITCHECKOK: out    vl_logic;
        TL2ASPMSUSPENDREQ: out    vl_logic;
        TL2ERRFCPE      : out    vl_logic;
        TL2ERRHDR       : out    vl_logic_vector(63 downto 0);
        TL2ERRMALFORMED : out    vl_logic;
        TL2ERRRXOVERFLOW: out    vl_logic;
        TL2PPMSUSPENDOK : out    vl_logic;
        TRNFCCPLD       : out    vl_logic_vector(11 downto 0);
        TRNFCCPLH       : out    vl_logic_vector(7 downto 0);
        TRNFCNPD        : out    vl_logic_vector(11 downto 0);
        TRNFCNPH        : out    vl_logic_vector(7 downto 0);
        TRNFCPD         : out    vl_logic_vector(11 downto 0);
        TRNFCPH         : out    vl_logic_vector(7 downto 0);
        TRNLNKUP        : out    vl_logic;
        TRNRBARHIT      : out    vl_logic_vector(7 downto 0);
        TRNRD           : out    vl_logic_vector(127 downto 0);
        TRNRDLLPDATA    : out    vl_logic_vector(63 downto 0);
        TRNRDLLPSRCRDY  : out    vl_logic_vector(1 downto 0);
        TRNRECRCERR     : out    vl_logic;
        TRNREOF         : out    vl_logic;
        TRNRERRFWD      : out    vl_logic;
        TRNRREM         : out    vl_logic_vector(1 downto 0);
        TRNRSOF         : out    vl_logic;
        TRNRSRCDSC      : out    vl_logic;
        TRNRSRCRDY      : out    vl_logic;
        TRNTBUFAV       : out    vl_logic_vector(5 downto 0);
        TRNTCFGREQ      : out    vl_logic;
        TRNTDLLPDSTRDY  : out    vl_logic;
        TRNTDSTRDY      : out    vl_logic_vector(3 downto 0);
        TRNTERRDROP     : out    vl_logic;
        USERRSTN        : out    vl_logic;
        CFGAERINTERRUPTMSGNUM: in     vl_logic_vector(4 downto 0);
        CFGDEVID        : in     vl_logic_vector(15 downto 0);
        CFGDSBUSNUMBER  : in     vl_logic_vector(7 downto 0);
        CFGDSDEVICENUMBER: in     vl_logic_vector(4 downto 0);
        CFGDSFUNCTIONNUMBER: in     vl_logic_vector(2 downto 0);
        CFGDSN          : in     vl_logic_vector(63 downto 0);
        CFGERRACSN      : in     vl_logic;
        CFGERRAERHEADERLOG: in     vl_logic_vector(127 downto 0);
        CFGERRATOMICEGRESSBLOCKEDN: in     vl_logic;
        CFGERRCORN      : in     vl_logic;
        CFGERRCPLABORTN : in     vl_logic;
        CFGERRCPLTIMEOUTN: in     vl_logic;
        CFGERRCPLUNEXPECTN: in     vl_logic;
        CFGERRECRCN     : in     vl_logic;
        CFGERRINTERNALCORN: in     vl_logic;
        CFGERRINTERNALUNCORN: in     vl_logic;
        CFGERRLOCKEDN   : in     vl_logic;
        CFGERRMALFORMEDN: in     vl_logic;
        CFGERRMCBLOCKEDN: in     vl_logic;
        CFGERRNORECOVERYN: in     vl_logic;
        CFGERRPOISONEDN : in     vl_logic;
        CFGERRPOSTEDN   : in     vl_logic;
        CFGERRTLPCPLHEADER: in     vl_logic_vector(47 downto 0);
        CFGERRURN       : in     vl_logic;
        CFGFORCECOMMONCLOCKOFF: in     vl_logic;
        CFGFORCEEXTENDEDSYNCON: in     vl_logic;
        CFGFORCEMPS     : in     vl_logic_vector(2 downto 0);
        CFGINTERRUPTASSERTN: in     vl_logic;
        CFGINTERRUPTDI  : in     vl_logic_vector(7 downto 0);
        CFGINTERRUPTN   : in     vl_logic;
        CFGINTERRUPTSTATN: in     vl_logic;
        CFGMGMTBYTEENN  : in     vl_logic_vector(3 downto 0);
        CFGMGMTDI       : in     vl_logic_vector(31 downto 0);
        CFGMGMTDWADDR   : in     vl_logic_vector(9 downto 0);
        CFGMGMTRDENN    : in     vl_logic;
        CFGMGMTWRENN    : in     vl_logic;
        CFGMGMTWRREADONLYN: in     vl_logic;
        CFGMGMTWRRW1CASRWN: in     vl_logic;
        CFGPCIECAPINTERRUPTMSGNUM: in     vl_logic_vector(4 downto 0);
        CFGPMFORCESTATE : in     vl_logic_vector(1 downto 0);
        CFGPMFORCESTATEENN: in     vl_logic;
        CFGPMHALTASPML0SN: in     vl_logic;
        CFGPMHALTASPML1N: in     vl_logic;
        CFGPMSENDPMETON : in     vl_logic;
        CFGPMTURNOFFOKN : in     vl_logic;
        CFGPMWAKEN      : in     vl_logic;
        CFGPORTNUMBER   : in     vl_logic_vector(7 downto 0);
        CFGREVID        : in     vl_logic_vector(7 downto 0);
        CFGSUBSYSID     : in     vl_logic_vector(15 downto 0);
        CFGSUBSYSVENDID : in     vl_logic_vector(15 downto 0);
        CFGTRNPENDINGN  : in     vl_logic;
        CFGVENDID       : in     vl_logic_vector(15 downto 0);
        CMRSTN          : in     vl_logic;
        CMSTICKYRSTN    : in     vl_logic;
        DBGMODE         : in     vl_logic_vector(1 downto 0);
        DBGSUBMODE      : in     vl_logic;
        DLRSTN          : in     vl_logic;
        DRPADDR         : in     vl_logic_vector(8 downto 0);
        DRPCLK          : in     vl_logic;
        DRPDI           : in     vl_logic_vector(15 downto 0);
        DRPEN           : in     vl_logic;
        DRPWE           : in     vl_logic;
        FUNCLVLRSTN     : in     vl_logic;
        LL2SENDASREQL1  : in     vl_logic;
        LL2SENDENTERL1  : in     vl_logic;
        LL2SENDENTERL23 : in     vl_logic;
        LL2SENDPMACK    : in     vl_logic;
        LL2SUSPENDNOW   : in     vl_logic;
        LL2TLPRCV       : in     vl_logic;
        MIMRXRDATA      : in     vl_logic_vector(67 downto 0);
        MIMTXRDATA      : in     vl_logic_vector(68 downto 0);
        PIPECLK         : in     vl_logic;
        PIPERX0CHANISALIGNED: in     vl_logic;
        PIPERX0CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX0DATA     : in     vl_logic_vector(15 downto 0);
        PIPERX0ELECIDLE : in     vl_logic;
        PIPERX0PHYSTATUS: in     vl_logic;
        PIPERX0STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX0VALID    : in     vl_logic;
        PIPERX1CHANISALIGNED: in     vl_logic;
        PIPERX1CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX1DATA     : in     vl_logic_vector(15 downto 0);
        PIPERX1ELECIDLE : in     vl_logic;
        PIPERX1PHYSTATUS: in     vl_logic;
        PIPERX1STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX1VALID    : in     vl_logic;
        PIPERX2CHANISALIGNED: in     vl_logic;
        PIPERX2CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX2DATA     : in     vl_logic_vector(15 downto 0);
        PIPERX2ELECIDLE : in     vl_logic;
        PIPERX2PHYSTATUS: in     vl_logic;
        PIPERX2STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX2VALID    : in     vl_logic;
        PIPERX3CHANISALIGNED: in     vl_logic;
        PIPERX3CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX3DATA     : in     vl_logic_vector(15 downto 0);
        PIPERX3ELECIDLE : in     vl_logic;
        PIPERX3PHYSTATUS: in     vl_logic;
        PIPERX3STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX3VALID    : in     vl_logic;
        PIPERX4CHANISALIGNED: in     vl_logic;
        PIPERX4CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX4DATA     : in     vl_logic_vector(15 downto 0);
        PIPERX4ELECIDLE : in     vl_logic;
        PIPERX4PHYSTATUS: in     vl_logic;
        PIPERX4STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX4VALID    : in     vl_logic;
        PIPERX5CHANISALIGNED: in     vl_logic;
        PIPERX5CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX5DATA     : in     vl_logic_vector(15 downto 0);
        PIPERX5ELECIDLE : in     vl_logic;
        PIPERX5PHYSTATUS: in     vl_logic;
        PIPERX5STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX5VALID    : in     vl_logic;
        PIPERX6CHANISALIGNED: in     vl_logic;
        PIPERX6CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX6DATA     : in     vl_logic_vector(15 downto 0);
        PIPERX6ELECIDLE : in     vl_logic;
        PIPERX6PHYSTATUS: in     vl_logic;
        PIPERX6STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX6VALID    : in     vl_logic;
        PIPERX7CHANISALIGNED: in     vl_logic;
        PIPERX7CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX7DATA     : in     vl_logic_vector(15 downto 0);
        PIPERX7ELECIDLE : in     vl_logic;
        PIPERX7PHYSTATUS: in     vl_logic;
        PIPERX7STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX7VALID    : in     vl_logic;
        PL2DIRECTEDLSTATE: in     vl_logic_vector(4 downto 0);
        PLDBGMODE       : in     vl_logic_vector(2 downto 0);
        PLDIRECTEDLINKAUTON: in     vl_logic;
        PLDIRECTEDLINKCHANGE: in     vl_logic_vector(1 downto 0);
        PLDIRECTEDLINKSPEED: in     vl_logic;
        PLDIRECTEDLINKWIDTH: in     vl_logic_vector(1 downto 0);
        PLDIRECTEDLTSSMNEW: in     vl_logic_vector(5 downto 0);
        PLDIRECTEDLTSSMNEWVLD: in     vl_logic;
        PLDIRECTEDLTSSMSTALL: in     vl_logic;
        PLDOWNSTREAMDEEMPHSOURCE: in     vl_logic;
        PLRSTN          : in     vl_logic;
        PLTRANSMITHOTRST: in     vl_logic;
        PLUPSTREAMPREFERDEEMPH: in     vl_logic;
        SYSRSTN         : in     vl_logic;
        TL2ASPMSUSPENDCREDITCHECK: in     vl_logic;
        TL2PPMSUSPENDREQ: in     vl_logic;
        TLRSTN          : in     vl_logic;
        TRNFCSEL        : in     vl_logic_vector(2 downto 0);
        TRNRDSTRDY      : in     vl_logic;
        TRNRFCPRET      : in     vl_logic;
        TRNRNPOK        : in     vl_logic;
        TRNRNPREQ       : in     vl_logic;
        TRNTCFGGNT      : in     vl_logic;
        TRNTD           : in     vl_logic_vector(127 downto 0);
        TRNTDLLPDATA    : in     vl_logic_vector(31 downto 0);
        TRNTDLLPSRCRDY  : in     vl_logic;
        TRNTECRCGEN     : in     vl_logic;
        TRNTEOF         : in     vl_logic;
        TRNTERRFWD      : in     vl_logic;
        TRNTREM         : in     vl_logic_vector(1 downto 0);
        TRNTSOF         : in     vl_logic;
        TRNTSRCDSC      : in     vl_logic;
        TRNTSRCRDY      : in     vl_logic;
        TRNTSTR         : in     vl_logic;
        USERCLK         : in     vl_logic;
        USERCLK2        : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of AER_BASE_PTR : constant is 1;
    attribute mti_svvh_generic_type of AER_CAP_ECRC_CHECK_CAPABLE : constant is 1;
    attribute mti_svvh_generic_type of AER_CAP_ECRC_GEN_CAPABLE : constant is 1;
    attribute mti_svvh_generic_type of AER_CAP_ID : constant is 1;
    attribute mti_svvh_generic_type of AER_CAP_MULTIHEADER : constant is 1;
    attribute mti_svvh_generic_type of AER_CAP_NEXTPTR : constant is 1;
    attribute mti_svvh_generic_type of AER_CAP_ON : constant is 1;
    attribute mti_svvh_generic_type of AER_CAP_OPTIONAL_ERR_SUPPORT : constant is 1;
    attribute mti_svvh_generic_type of AER_CAP_PERMIT_ROOTERR_UPDATE : constant is 1;
    attribute mti_svvh_generic_type of AER_CAP_VERSION : constant is 1;
    attribute mti_svvh_generic_type of ALLOW_X8_GEN2 : constant is 1;
    attribute mti_svvh_generic_type of BAR0 : constant is 1;
    attribute mti_svvh_generic_type of BAR1 : constant is 1;
    attribute mti_svvh_generic_type of BAR2 : constant is 1;
    attribute mti_svvh_generic_type of BAR3 : constant is 1;
    attribute mti_svvh_generic_type of BAR4 : constant is 1;
    attribute mti_svvh_generic_type of BAR5 : constant is 1;
    attribute mti_svvh_generic_type of CAPABILITIES_PTR : constant is 1;
    attribute mti_svvh_generic_type of CARDBUS_CIS_POINTER : constant is 1;
    attribute mti_svvh_generic_type of CFG_ECRC_ERR_CPLSTAT : constant is 2;
    attribute mti_svvh_generic_type of CLASS_CODE : constant is 1;
    attribute mti_svvh_generic_type of CMD_INTX_IMPLEMENTED : constant is 1;
    attribute mti_svvh_generic_type of CPL_TIMEOUT_DISABLE_SUPPORTED : constant is 1;
    attribute mti_svvh_generic_type of CPL_TIMEOUT_RANGES_SUPPORTED : constant is 1;
    attribute mti_svvh_generic_type of CRM_MODULE_RSTS : constant is 1;
    attribute mti_svvh_generic_type of DEV_CAP2_ARI_FORWARDING_SUPPORTED : constant is 1;
    attribute mti_svvh_generic_type of DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED : constant is 1;
    attribute mti_svvh_generic_type of DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED : constant is 1;
    attribute mti_svvh_generic_type of DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED : constant is 1;
    attribute mti_svvh_generic_type of DEV_CAP2_CAS128_COMPLETER_SUPPORTED : constant is 1;
    attribute mti_svvh_generic_type of DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED : constant is 1;
    attribute mti_svvh_generic_type of DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED : constant is 1;
    attribute mti_svvh_generic_type of DEV_CAP2_LTR_MECHANISM_SUPPORTED : constant is 1;
    attribute mti_svvh_generic_type of DEV_CAP2_MAX_ENDEND_TLP_PREFIXES : constant is 1;
    attribute mti_svvh_generic_type of DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING : constant is 1;
    attribute mti_svvh_generic_type of DEV_CAP2_TPH_COMPLETER_SUPPORTED : constant is 1;
    attribute mti_svvh_generic_type of DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE : constant is 1;
    attribute mti_svvh_generic_type of DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE : constant is 1;
    attribute mti_svvh_generic_type of DEV_CAP_ENDPOINT_L0S_LATENCY : constant is 2;
    attribute mti_svvh_generic_type of DEV_CAP_ENDPOINT_L1_LATENCY : constant is 2;
    attribute mti_svvh_generic_type of DEV_CAP_EXT_TAG_SUPPORTED : constant is 1;
    attribute mti_svvh_generic_type of DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE : constant is 1;
    attribute mti_svvh_generic_type of DEV_CAP_MAX_PAYLOAD_SUPPORTED : constant is 2;
    attribute mti_svvh_generic_type of DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT : constant is 2;
    attribute mti_svvh_generic_type of DEV_CAP_ROLE_BASED_ERROR : constant is 1;
    attribute mti_svvh_generic_type of DEV_CAP_RSVD_14_12 : constant is 2;
    attribute mti_svvh_generic_type of DEV_CAP_RSVD_17_16 : constant is 2;
    attribute mti_svvh_generic_type of DEV_CAP_RSVD_31_29 : constant is 2;
    attribute mti_svvh_generic_type of DEV_CONTROL_AUX_POWER_SUPPORTED : constant is 1;
    attribute mti_svvh_generic_type of DEV_CONTROL_EXT_TAG_DEFAULT : constant is 1;
    attribute mti_svvh_generic_type of DISABLE_ASPM_L1_TIMER : constant is 1;
    attribute mti_svvh_generic_type of DISABLE_BAR_FILTERING : constant is 1;
    attribute mti_svvh_generic_type of DISABLE_ERR_MSG : constant is 1;
    attribute mti_svvh_generic_type of DISABLE_ID_CHECK : constant is 1;
    attribute mti_svvh_generic_type of DISABLE_LANE_REVERSAL : constant is 1;
    attribute mti_svvh_generic_type of DISABLE_LOCKED_FILTER : constant is 1;
    attribute mti_svvh_generic_type of DISABLE_PPM_FILTER : constant is 1;
    attribute mti_svvh_generic_type of DISABLE_RX_POISONED_RESP : constant is 1;
    attribute mti_svvh_generic_type of DISABLE_RX_TC_FILTER : constant is 1;
    attribute mti_svvh_generic_type of DISABLE_SCRAMBLING : constant is 1;
    attribute mti_svvh_generic_type of DNSTREAM_LINK_NUM : constant is 1;
    attribute mti_svvh_generic_type of DSN_BASE_PTR : constant is 1;
    attribute mti_svvh_generic_type of DSN_CAP_ID : constant is 1;
    attribute mti_svvh_generic_type of DSN_CAP_NEXTPTR : constant is 1;
    attribute mti_svvh_generic_type of DSN_CAP_ON : constant is 1;
    attribute mti_svvh_generic_type of DSN_CAP_VERSION : constant is 1;
    attribute mti_svvh_generic_type of ENABLE_MSG_ROUTE : constant is 1;
    attribute mti_svvh_generic_type of ENABLE_RX_TD_ECRC_TRIM : constant is 1;
    attribute mti_svvh_generic_type of ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED : constant is 1;
    attribute mti_svvh_generic_type of ENTER_RVRY_EI_L0 : constant is 1;
    attribute mti_svvh_generic_type of EXIT_LOOPBACK_ON_EI : constant is 1;
    attribute mti_svvh_generic_type of EXPANSION_ROM : constant is 1;
    attribute mti_svvh_generic_type of EXT_CFG_CAP_PTR : constant is 1;
    attribute mti_svvh_generic_type of EXT_CFG_XP_CAP_PTR : constant is 1;
    attribute mti_svvh_generic_type of HEADER_TYPE : constant is 1;
    attribute mti_svvh_generic_type of INFER_EI : constant is 1;
    attribute mti_svvh_generic_type of INTERRUPT_PIN : constant is 1;
    attribute mti_svvh_generic_type of INTERRUPT_STAT_AUTO : constant is 1;
    attribute mti_svvh_generic_type of IS_SWITCH : constant is 1;
    attribute mti_svvh_generic_type of LAST_CONFIG_DWORD : constant is 1;
    attribute mti_svvh_generic_type of LINK_CAP_ASPM_OPTIONALITY : constant is 1;
    attribute mti_svvh_generic_type of LINK_CAP_ASPM_SUPPORT : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_CLOCK_POWER_MANAGEMENT : constant is 1;
    attribute mti_svvh_generic_type of LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP : constant is 1;
    attribute mti_svvh_generic_type of LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_L0S_EXIT_LATENCY_GEN1 : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_L0S_EXIT_LATENCY_GEN2 : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_L1_EXIT_LATENCY_GEN1 : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_L1_EXIT_LATENCY_GEN2 : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP : constant is 1;
    attribute mti_svvh_generic_type of LINK_CAP_MAX_LINK_SPEED : constant is 1;
    attribute mti_svvh_generic_type of LINK_CAP_MAX_LINK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of LINK_CAP_RSVD_23 : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE : constant is 1;
    attribute mti_svvh_generic_type of LINK_CONTROL_RCB : constant is 2;
    attribute mti_svvh_generic_type of LINK_CTRL2_DEEMPHASIS : constant is 1;
    attribute mti_svvh_generic_type of LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of LINK_CTRL2_TARGET_LINK_SPEED : constant is 1;
    attribute mti_svvh_generic_type of LINK_STATUS_SLOT_CLOCK_CONFIG : constant is 1;
    attribute mti_svvh_generic_type of LL_ACK_TIMEOUT : constant is 1;
    attribute mti_svvh_generic_type of LL_ACK_TIMEOUT_EN : constant is 1;
    attribute mti_svvh_generic_type of LL_ACK_TIMEOUT_FUNC : constant is 2;
    attribute mti_svvh_generic_type of LL_REPLAY_TIMEOUT : constant is 1;
    attribute mti_svvh_generic_type of LL_REPLAY_TIMEOUT_EN : constant is 1;
    attribute mti_svvh_generic_type of LL_REPLAY_TIMEOUT_FUNC : constant is 2;
    attribute mti_svvh_generic_type of LTSSM_MAX_LINK_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of MPS_FORCE : constant is 1;
    attribute mti_svvh_generic_type of MSIX_BASE_PTR : constant is 1;
    attribute mti_svvh_generic_type of MSIX_CAP_ID : constant is 1;
    attribute mti_svvh_generic_type of MSIX_CAP_NEXTPTR : constant is 1;
    attribute mti_svvh_generic_type of MSIX_CAP_ON : constant is 1;
    attribute mti_svvh_generic_type of MSIX_CAP_PBA_BIR : constant is 2;
    attribute mti_svvh_generic_type of MSIX_CAP_PBA_OFFSET : constant is 1;
    attribute mti_svvh_generic_type of MSIX_CAP_TABLE_BIR : constant is 2;
    attribute mti_svvh_generic_type of MSIX_CAP_TABLE_OFFSET : constant is 1;
    attribute mti_svvh_generic_type of MSIX_CAP_TABLE_SIZE : constant is 1;
    attribute mti_svvh_generic_type of MSI_BASE_PTR : constant is 1;
    attribute mti_svvh_generic_type of MSI_CAP_64_BIT_ADDR_CAPABLE : constant is 1;
    attribute mti_svvh_generic_type of MSI_CAP_ID : constant is 1;
    attribute mti_svvh_generic_type of MSI_CAP_MULTIMSGCAP : constant is 2;
    attribute mti_svvh_generic_type of MSI_CAP_MULTIMSG_EXTENSION : constant is 2;
    attribute mti_svvh_generic_type of MSI_CAP_NEXTPTR : constant is 1;
    attribute mti_svvh_generic_type of MSI_CAP_ON : constant is 1;
    attribute mti_svvh_generic_type of MSI_CAP_PER_VECTOR_MASKING_CAPABLE : constant is 1;
    attribute mti_svvh_generic_type of N_FTS_COMCLK_GEN1 : constant is 2;
    attribute mti_svvh_generic_type of N_FTS_COMCLK_GEN2 : constant is 2;
    attribute mti_svvh_generic_type of N_FTS_GEN1 : constant is 2;
    attribute mti_svvh_generic_type of N_FTS_GEN2 : constant is 2;
    attribute mti_svvh_generic_type of PCIE_BASE_PTR : constant is 1;
    attribute mti_svvh_generic_type of PCIE_CAP_CAPABILITY_ID : constant is 1;
    attribute mti_svvh_generic_type of PCIE_CAP_CAPABILITY_VERSION : constant is 1;
    attribute mti_svvh_generic_type of PCIE_CAP_DEVICE_PORT_TYPE : constant is 1;
    attribute mti_svvh_generic_type of PCIE_CAP_NEXTPTR : constant is 1;
    attribute mti_svvh_generic_type of PCIE_CAP_ON : constant is 1;
    attribute mti_svvh_generic_type of PCIE_CAP_RSVD_15_14 : constant is 2;
    attribute mti_svvh_generic_type of PCIE_CAP_SLOT_IMPLEMENTED : constant is 1;
    attribute mti_svvh_generic_type of PCIE_REVISION : constant is 2;
    attribute mti_svvh_generic_type of PL_AUTO_CONFIG : constant is 2;
    attribute mti_svvh_generic_type of PL_FAST_TRAIN : constant is 1;
    attribute mti_svvh_generic_type of PM_ASPML0S_TIMEOUT : constant is 1;
    attribute mti_svvh_generic_type of PM_ASPML0S_TIMEOUT_EN : constant is 1;
    attribute mti_svvh_generic_type of PM_ASPML0S_TIMEOUT_FUNC : constant is 2;
    attribute mti_svvh_generic_type of PM_ASPM_FASTEXIT : constant is 1;
    attribute mti_svvh_generic_type of PM_BASE_PTR : constant is 1;
    attribute mti_svvh_generic_type of PM_CAP_AUXCURRENT : constant is 2;
    attribute mti_svvh_generic_type of PM_CAP_D1SUPPORT : constant is 1;
    attribute mti_svvh_generic_type of PM_CAP_D2SUPPORT : constant is 1;
    attribute mti_svvh_generic_type of PM_CAP_DSI : constant is 1;
    attribute mti_svvh_generic_type of PM_CAP_ID : constant is 1;
    attribute mti_svvh_generic_type of PM_CAP_NEXTPTR : constant is 1;
    attribute mti_svvh_generic_type of PM_CAP_ON : constant is 1;
    attribute mti_svvh_generic_type of PM_CAP_PMESUPPORT : constant is 1;
    attribute mti_svvh_generic_type of PM_CAP_PME_CLOCK : constant is 1;
    attribute mti_svvh_generic_type of PM_CAP_RSVD_04 : constant is 2;
    attribute mti_svvh_generic_type of PM_CAP_VERSION : constant is 2;
    attribute mti_svvh_generic_type of PM_CSR_B2B3 : constant is 1;
    attribute mti_svvh_generic_type of PM_CSR_BPCCEN : constant is 1;
    attribute mti_svvh_generic_type of PM_CSR_NOSOFTRST : constant is 1;
    attribute mti_svvh_generic_type of PM_DATA0 : constant is 1;
    attribute mti_svvh_generic_type of PM_DATA1 : constant is 1;
    attribute mti_svvh_generic_type of PM_DATA2 : constant is 1;
    attribute mti_svvh_generic_type of PM_DATA3 : constant is 1;
    attribute mti_svvh_generic_type of PM_DATA4 : constant is 1;
    attribute mti_svvh_generic_type of PM_DATA5 : constant is 1;
    attribute mti_svvh_generic_type of PM_DATA6 : constant is 1;
    attribute mti_svvh_generic_type of PM_DATA7 : constant is 1;
    attribute mti_svvh_generic_type of PM_DATA_SCALE0 : constant is 1;
    attribute mti_svvh_generic_type of PM_DATA_SCALE1 : constant is 1;
    attribute mti_svvh_generic_type of PM_DATA_SCALE2 : constant is 1;
    attribute mti_svvh_generic_type of PM_DATA_SCALE3 : constant is 1;
    attribute mti_svvh_generic_type of PM_DATA_SCALE4 : constant is 1;
    attribute mti_svvh_generic_type of PM_DATA_SCALE5 : constant is 1;
    attribute mti_svvh_generic_type of PM_DATA_SCALE6 : constant is 1;
    attribute mti_svvh_generic_type of PM_DATA_SCALE7 : constant is 1;
    attribute mti_svvh_generic_type of PM_MF : constant is 1;
    attribute mti_svvh_generic_type of RBAR_BASE_PTR : constant is 1;
    attribute mti_svvh_generic_type of RBAR_CAP_CONTROL_ENCODEDBAR0 : constant is 1;
    attribute mti_svvh_generic_type of RBAR_CAP_CONTROL_ENCODEDBAR1 : constant is 1;
    attribute mti_svvh_generic_type of RBAR_CAP_CONTROL_ENCODEDBAR2 : constant is 1;
    attribute mti_svvh_generic_type of RBAR_CAP_CONTROL_ENCODEDBAR3 : constant is 1;
    attribute mti_svvh_generic_type of RBAR_CAP_CONTROL_ENCODEDBAR4 : constant is 1;
    attribute mti_svvh_generic_type of RBAR_CAP_CONTROL_ENCODEDBAR5 : constant is 1;
    attribute mti_svvh_generic_type of RBAR_CAP_ID : constant is 1;
    attribute mti_svvh_generic_type of RBAR_CAP_INDEX0 : constant is 1;
    attribute mti_svvh_generic_type of RBAR_CAP_INDEX1 : constant is 1;
    attribute mti_svvh_generic_type of RBAR_CAP_INDEX2 : constant is 1;
    attribute mti_svvh_generic_type of RBAR_CAP_INDEX3 : constant is 1;
    attribute mti_svvh_generic_type of RBAR_CAP_INDEX4 : constant is 1;
    attribute mti_svvh_generic_type of RBAR_CAP_INDEX5 : constant is 1;
    attribute mti_svvh_generic_type of RBAR_CAP_NEXTPTR : constant is 1;
    attribute mti_svvh_generic_type of RBAR_CAP_ON : constant is 1;
    attribute mti_svvh_generic_type of RBAR_CAP_SUP0 : constant is 1;
    attribute mti_svvh_generic_type of RBAR_CAP_SUP1 : constant is 1;
    attribute mti_svvh_generic_type of RBAR_CAP_SUP2 : constant is 1;
    attribute mti_svvh_generic_type of RBAR_CAP_SUP3 : constant is 1;
    attribute mti_svvh_generic_type of RBAR_CAP_SUP4 : constant is 1;
    attribute mti_svvh_generic_type of RBAR_CAP_SUP5 : constant is 1;
    attribute mti_svvh_generic_type of RBAR_CAP_VERSION : constant is 1;
    attribute mti_svvh_generic_type of RBAR_NUM : constant is 1;
    attribute mti_svvh_generic_type of RECRC_CHK : constant is 2;
    attribute mti_svvh_generic_type of RECRC_CHK_TRIM : constant is 1;
    attribute mti_svvh_generic_type of ROOT_CAP_CRS_SW_VISIBILITY : constant is 1;
    attribute mti_svvh_generic_type of RP_AUTO_SPD : constant is 1;
    attribute mti_svvh_generic_type of RP_AUTO_SPD_LOOPCNT : constant is 1;
    attribute mti_svvh_generic_type of SELECT_DLL_IF : constant is 1;
    attribute mti_svvh_generic_type of SIM_VERSION : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CAP_ATT_BUTTON_PRESENT : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CAP_ATT_INDICATOR_PRESENT : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CAP_ELEC_INTERLOCK_PRESENT : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CAP_HOTPLUG_CAPABLE : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CAP_HOTPLUG_SURPRISE : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CAP_MRL_SENSOR_PRESENT : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CAP_NO_CMD_COMPLETED_SUPPORT : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CAP_PHYSICAL_SLOT_NUM : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CAP_POWER_CONTROLLER_PRESENT : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CAP_POWER_INDICATOR_PRESENT : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CAP_SLOT_POWER_LIMIT_SCALE : constant is 2;
    attribute mti_svvh_generic_type of SLOT_CAP_SLOT_POWER_LIMIT_VALUE : constant is 1;
    attribute mti_svvh_generic_type of SPARE_BIT0 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT1 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT2 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT3 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT4 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT5 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT6 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT7 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT8 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BYTE0 : constant is 1;
    attribute mti_svvh_generic_type of SPARE_BYTE1 : constant is 1;
    attribute mti_svvh_generic_type of SPARE_BYTE2 : constant is 1;
    attribute mti_svvh_generic_type of SPARE_BYTE3 : constant is 1;
    attribute mti_svvh_generic_type of SPARE_WORD0 : constant is 1;
    attribute mti_svvh_generic_type of SPARE_WORD1 : constant is 1;
    attribute mti_svvh_generic_type of SPARE_WORD2 : constant is 1;
    attribute mti_svvh_generic_type of SPARE_WORD3 : constant is 1;
    attribute mti_svvh_generic_type of SSL_MESSAGE_AUTO : constant is 1;
    attribute mti_svvh_generic_type of TECRC_EP_INV : constant is 1;
    attribute mti_svvh_generic_type of TL_RBYPASS : constant is 1;
    attribute mti_svvh_generic_type of TL_RX_RAM_RADDR_LATENCY : constant is 2;
    attribute mti_svvh_generic_type of TL_RX_RAM_RDATA_LATENCY : constant is 2;
    attribute mti_svvh_generic_type of TL_RX_RAM_WRITE_LATENCY : constant is 2;
    attribute mti_svvh_generic_type of TL_TFC_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of TL_TX_CHECKS_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of TL_TX_RAM_RADDR_LATENCY : constant is 2;
    attribute mti_svvh_generic_type of TL_TX_RAM_RDATA_LATENCY : constant is 2;
    attribute mti_svvh_generic_type of TL_TX_RAM_WRITE_LATENCY : constant is 2;
    attribute mti_svvh_generic_type of TRN_DW : constant is 1;
    attribute mti_svvh_generic_type of TRN_NP_FC : constant is 1;
    attribute mti_svvh_generic_type of UPCONFIG_CAPABLE : constant is 1;
    attribute mti_svvh_generic_type of UPSTREAM_FACING : constant is 1;
    attribute mti_svvh_generic_type of UR_ATOMIC : constant is 1;
    attribute mti_svvh_generic_type of UR_CFG1 : constant is 1;
    attribute mti_svvh_generic_type of UR_INV_REQ : constant is 1;
    attribute mti_svvh_generic_type of UR_PRS_RESPONSE : constant is 1;
    attribute mti_svvh_generic_type of USER_CLK2_DIV2 : constant is 1;
    attribute mti_svvh_generic_type of USER_CLK_FREQ : constant is 2;
    attribute mti_svvh_generic_type of USE_RID_PINS : constant is 1;
    attribute mti_svvh_generic_type of VC0_CPL_INFINITE : constant is 1;
    attribute mti_svvh_generic_type of VC0_RX_RAM_LIMIT : constant is 1;
    attribute mti_svvh_generic_type of VC0_TOTAL_CREDITS_CD : constant is 2;
    attribute mti_svvh_generic_type of VC0_TOTAL_CREDITS_CH : constant is 2;
    attribute mti_svvh_generic_type of VC0_TOTAL_CREDITS_NPD : constant is 2;
    attribute mti_svvh_generic_type of VC0_TOTAL_CREDITS_NPH : constant is 2;
    attribute mti_svvh_generic_type of VC0_TOTAL_CREDITS_PD : constant is 2;
    attribute mti_svvh_generic_type of VC0_TOTAL_CREDITS_PH : constant is 2;
    attribute mti_svvh_generic_type of VC0_TX_LASTPACKET : constant is 2;
    attribute mti_svvh_generic_type of VC_BASE_PTR : constant is 1;
    attribute mti_svvh_generic_type of VC_CAP_ID : constant is 1;
    attribute mti_svvh_generic_type of VC_CAP_NEXTPTR : constant is 1;
    attribute mti_svvh_generic_type of VC_CAP_ON : constant is 1;
    attribute mti_svvh_generic_type of VC_CAP_REJECT_SNOOP_TRANSACTIONS : constant is 1;
    attribute mti_svvh_generic_type of VC_CAP_VERSION : constant is 1;
    attribute mti_svvh_generic_type of VSEC_BASE_PTR : constant is 1;
    attribute mti_svvh_generic_type of VSEC_CAP_HDR_ID : constant is 1;
    attribute mti_svvh_generic_type of VSEC_CAP_HDR_LENGTH : constant is 1;
    attribute mti_svvh_generic_type of VSEC_CAP_HDR_REVISION : constant is 1;
    attribute mti_svvh_generic_type of VSEC_CAP_ID : constant is 1;
    attribute mti_svvh_generic_type of VSEC_CAP_IS_LINK_VISIBLE : constant is 1;
    attribute mti_svvh_generic_type of VSEC_CAP_NEXTPTR : constant is 1;
    attribute mti_svvh_generic_type of VSEC_CAP_ON : constant is 1;
    attribute mti_svvh_generic_type of VSEC_CAP_VERSION : constant is 1;
end PCIE_2_1_WRAP;
