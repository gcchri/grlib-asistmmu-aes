`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wp0MZwO7K+UJzUHGFasTHw28Ie8IOhLBDc+6PNNjcZc9iHPW2HnFL6lLMsFIToiY
Uzl3VuFnrt6OFGLaysmJuXvB1Jw78CD8oH30rpfEZ+1ok6MGT6L1vn64f/x/jmrL
S+08v/FdK9SXjO0p266rM4o/jiebcS0W3qez8vSZM5YLddqpuvkZyrEwyO7UkRiR
p93g6en5/LLyUyyKq2cCLwyBz7InCBLeZWG36oIo0R11J5z46oorAh1A0ykn52pg
cGNXNeNcRS5IVOVedSb1y/zW3lPeWARD8eTucsLzuJj7UklYMxPd7DDp1dITlyYn
4hR3NQtrX6bjWQNaBBUnNfu5bYcu2ICJ9KhnrUNu1ZUusU5EdBoPv59gEBRNbbqX
/AiNPrVkxRzPcy8lxB0Qxg==
`protect END_PROTECTED
