`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xyaDb+Nfae/k3zLxPA6UIVtshvNq6LxQjBRBk4eQcLqOC97ho9+c6VmW7/nv5fFo
nC7CeiKfKoOuHqKA6WE1JaVv5xMJqZ1mUF1ss/Qm1us9kuDRvcKF+R4tPZ47RIk6
NUtEz0MfU+Z7Nx8BQ+95J1jH6bGVVO/OFSn8zf7kTduOuCzSILl08juKo3DiFmju
OuCHkpBdnvN2H69Xvt4WFD5xg8d2fDStIe9+S/xKQbtKBSOfu5tOov19fDI+8e6K
SoiPD8nCWLpv6i8kxIfUxMzg8NGwDkjp2lJuppZh6xu8RYQgArpSVf9SsakeND74
IJuIKiNqHVtfOp3kIppkRg==
`protect END_PROTECTED
