`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2xXC9aQ4Yv/v2M9qaSx87ODAbXJyoqdHJzOlks/bPp/OiYTEPpO87Y0tGqG9Olai
fxYM2DHDMJJzRI9Cr+788Y1N2AMC0IjEojHWPu8UD7DJuGqNxA170yPGxqaidVqH
6wY8YuGuhbyPjbKUW4FXvjTzKEcKxN0JPTnwbfPDH4OIV6Io+X2Mqn+uzWDh1BMg
toIZfZghNDkNiIBIUnUQYxBJdAIjNub3i620RiOYqKhOlTIx/Dx8bJWzDqaCPsyl
/aw3uHbpebJCaBYWv6AVAhn05KPS9kGS6Kombqy0kHAMTZKi5bvbxm8Bu7pCjwFP
cCN17ql8p8LLlvP3hVZYs1KkHb4TuDc44oPa6f9YI3lJ5xQKtgAFgCr4+ZLTqgds
ehsf6yF+ug96ByjbB5ikV61+k4RMmtkDpsyPJJB2DfFHvFeWrHw6wtyo/scuGdz+
fVXv6UVgDVaZk0E26Mo9nWWra2vJ0kRtOWwpav5ySEeC3kL+zqmxo5SEgpFiyYKQ
3Oj4MW+B82UOfRyqeixiSadP2OmaCW+uXG0pQTDdJXWkDrX4NCR70MIgWu3vtnOU
IfHo523S0XnfyZVqWlwVW5gz/C75wC0ohdC3Gv62DPUVdprcrs1G1/WXisBHQ4CW
frpW8o4xm4KP6tf0vC17819IPeRnSK4Mnku1ezcScmUPuoaE2KqKNpwwSp61BuwJ
Kqn5WYByNbXkSlt8FDyI1pAgpBVgIvTwSZnD2jAR/gh/zgtweuPm5Bg+C+aoaYW5
9pm+Xpy7DwixFbUblOqOwHQohabOfg7T4CVID4T7Z1WkXlmKVPvCFnfZl0BLc8KI
8mcv0fXTAz83jW8ZZXGb1n7wSx/cbNKtKDt0EfEDGxNS1jnDH+GpNtc6mJXXr1Rf
ggkvVfS/rmoGNLD0CcUK44wI6aqSal4nY2a5QxCSQSePiiixSU8A5dixAHntyEfu
dLbDuKzxiXHMtJ8wusuLEztjSJiUCGc3ZhRfl19qUM28DrsrnNpy5Y/cMGXveBBO
`protect END_PROTECTED
