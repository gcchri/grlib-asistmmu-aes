`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8xZJmI6NGlZg1wlsIRb32vkySocWU8SmbS4e2WZjMTWQZkoqpSunEY/AZRNFXQcZ
UnPCmm8PKTZJxQyiURScp47bnoHKMHu1Wv1Cs508t6xXIg/RGU0qwrfoMUcKuzRO
IbEaU4VlLEmauIUZ12NT0NZ3DzeBwFvAydlu0j94ubw8n+aSqcaxILGI2H+idMT9
2FFYJkGoogjYCmywn5HhX2ByeW4hJBqckoQLejprnqxJnPBrmzFgqTFxeZtpt7cw
VatQ644AhRD+Tr0HjGQtwjBmWAxRnR3VO1F/m/46roeeG5TVMJ3Qq+j9N2lFtrZ/
CyoknZC0Wp+By7AlUssKS8nPyey4lpACUdn77QP7VVsyuJq8EL+tmDc5vCfscHYJ
`protect END_PROTECTED
