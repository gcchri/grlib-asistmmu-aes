`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WjiKkQzUic3MSnUQUeOWIiGasmANu2qcjA9mnN0QXtXdn/MxfdMyimuf9KVrEe9m
9hKSnnDmHcAKOiyhjPDG/0B/gyhggJDK/VrVJlO64Xd61gSbEJBHxm9BvUIWGQ1E
ZFuyI68iJ9F6PlIz/Xah8hn9Yr1aERxAgRrp7THed/20ZBPHwUtcudf5BHTHXmlt
IcXZebvVqUcDQJ5mu8YnQNsHYNMRTGF305h8kzmsAcMiOQCMhNfXKlueyvlvfhs1
5F3AIlMfylj5/QTZyVn8sA8F7Bsug/uBBugLEl3kOGl6DgkvfwYhXTRNM4T61r7X
p6vUcT+o43PUrvkULKG1+Vt4oWu4HztrPPoKuRUkyIggPY5JIFV55gg778AtoDYW
rIxKNTjlPz2S3r27Zo6Q63402haVU/a3mQWB5ns3yM5jRbw6ACsWFSvUdw0o9ybl
o4pDHh34eQuyBxKLpJWBqEfWd3Hi1udRyrkJgn0sWq3MP1bc6CxYuWnyh/ozniRI
RjVCsqU/OLTQOJKw7FSiOshNAi4Kff3Cjh+ep1g9ZGRpsgT9f426WCkHMZ9wFS+a
C/b5z/01dgDSQuAc8+KzP1B1Kb+hzXy5wcba+9rtmEIhDvLO8L1v6Djv4VjfdKXs
A5i0F7kY5z198KGX+zNm8qANIBYek17Yvb4z76E7TzmfB61A5Jkf51k54VUB1CSZ
L5D5QQGCsOH2BQ0MrIDUt3IuhBYU/2QndArxUOKKVhCyoOb67eIzMDSyJzQZOsq5
rg3QCvp7YRKZAh+e/rUXxg==
`protect END_PROTECTED
