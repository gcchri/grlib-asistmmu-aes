`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G7nDEBqMBNxXJAtBuzbDzDQGQjYmKFwlYN+jCNTzOOiOYpRwWBM2k0gaqje6XPk0
jPuaedhpE3jxVGNBue45HVfyPy7OAokjer05CwQIsBFJ5Lr3zocpiaujsnwEIXAf
SRSVX+WeTvdw5C0p7yOB2UA7ezo/DEXKtd1tMbhVvLzNMWNL3LeoGwazGzB95yTs
sb0tgjYH5kZ0yVgX48HhSwojpaxY6yMaxxuaMXd04HVVQSvmJkNZlQxc7I6oHk37
c3c3H7Q7ccspOniKflJljIICKA54m5Mjr5MDlVeAwxFDSNRTSCh7IDLZNtNS5gG9
yaQE4TcRlI5N8o5Lcr7WbrPN6uUyla1atUNE/TDGJaLms9RRLvWJ6NqybC/tiLi+
yJcr3ipLMsaDI0/1VmTM6wm2WAIs3j19qa6MGGYY4iXUmQ/t6nkpAdSl63nZU2r7
arj+ZwEFX2MUcljKL1Kag409RY57Zn5p6OnI5hXbULdkDCY8ojIXY2NjL+TuTss+
DO8ukOCBSHYnow6up9q8tw==
`protect END_PROTECTED
