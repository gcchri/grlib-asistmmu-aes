`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I/EIGnSiZ2xBe92XHAj1q5vAhzHZjookrnNJVxZ6kClG2FCfdmk8pP1nUeFFdPVT
L/1Ih4gjDCfithYtAqLX1mE6V77Qhxr4OIgLv/viAC1sBSWeXc8dtUEY22ShmTyC
EMzDWPitiwuZtgrYFG5TDyLq+berN5mu7uOG3qu87sdeUxKilFsg7GAbWLShbmEo
mSIPtbtPcyJ3sP9DgI+pGNLH24aQbGEhqXvcnqQ9n1FSI4I2GxIgSmTaGx4zRAgj
+yenMRpK9zUVsXoe+/718MRFgZz0NzXhwggAy9AqYM/5I0z+YnP2MHcwhisyy+ZR
dmHqQmGJ8NRzsfmFOnZWC72J2jTpKk0OxEaUhYdAkwE3gG0B6L+hv5yUhqoiy89j
51lK7H5Y3TeZotyenGuYm5a7xEb4Zp+9ZsmSKmynVr1mfj1/TNuKJUj4tizeXUa1
7C2KCpsHsWPsE0Gf5zRhCTwYPvlVj+oSrlj52zr/ATFcqhOFilS9jRuQ/YdbRplF
/Wuegxv26Cb8sgTaqG1PZ1DLcglw5CeFR978EM5eeD5Mn7aBd5j1J9S3K39M7AkU
tYHE5c+EQizZv106jZIw4tNoIfTeA0URtZEKseHRk2EhbgDhChRBUvDR7fG99B2M
wV8M8bMnxqQOXFRM0Nqo+uVRXT2BoCOZdMv04NyUZuk+gSWZa+68xY5w3STISBNh
JiCwrMHjN+srk9u8mwZakciJddQFHF9mKyvFLpWpe3tQSe5KjMAKhLs9EfNUT+Lz
w7eApkpbEkyMUQen/+mNaMZFocv6NxEUP9tZt/3KRbvznyOmcMSCpqPp69BKwOfU
fw5VCGV9HnLmBkF4eDmfzbxN2PjD+nQvZni7ZVGsK7v/l08Y07PQXTc4+CaKSJXw
YvXYloN1w/Z4gnvAVD9lEx/rSzfChz08XsiKs6cwHgsancJXm0zkqxyJd/2swcuZ
zZkHq1eGb+VtE1eMK+4HXUu3yUniIa/2jE9X0zFl8XO1axYEodPRX/oJLjA/q3Im
af7yJReD8cYdOatwqNRf4rS6iYJzhg7oKoO/yZQJlHmO2/DK8/6pld/zBG7/N9cK
CRvU4QDZxrmjqEkfSvzTC0edOgiHbO0dZUVd2M7Xvkec2Pdwao7tqG1gDMGqGdSZ
Bhgvsss0kUIoMOdVC2PoVoOffcqpiIlA2gMT3S630/qc9WvXe4qdyNCx5HYrqv9K
2ipxAUpabEdflyQDxvE/Npc3+EVixhI0IQ99HJxmO/NU42BQgsdW78o1XHuqMil5
0p30WsHVThZ9imwUN0njqD9H4qBIsU4/aaZAl6ID4jFgzL+Ygxd4yQW67sUlZOCT
gMQMn6LltcOAvt8WbzcQGgbxkQ1pAAgK/JIQXtpfvOCMMSW7xN7bMaJZmA/KNP8Q
OP4FIOxH/2Yn6SG++DnS+OuUOxxxwXlxsStoA5X7i39eW5PqQNi2Q2E8DpW8sIZG
T0rykbCAB5heuDlLQtA076RLmDU9uzqwifHuyPpwIRgAV9M3+rCk8msbQflz/bBX
Ov2e0yEsYlFxP4ROhFKkfMIBwx++yR85YcXNpDPx0GFRjLQxBdSFKar9Y3LQk5ah
BjLG33gsdv/h2ljw2Lnwz0lm9BPMsWScBFWBi10ue5gai72qTOh94DCE7KuHH3nQ
dDlo5dpsbmJa8pDtwHhBCJPSL2JQz0SrxJ0hqVfEeqcbQQzFDPawFTdZYPHAuCYG
xMEPSv7+TNhco5QCnK8e6uRhvVkHQwwC/TvBtYvNogFCT3VSPc32CdUajHKmQE8i
yFU3aiyIri/57/QVupmBQDCkyxR6wSNt4Hue5wIOGb5Awbw4T6Iw5zoEnzERUUyb
e7s49rWjN/9ouiAHm2aOsRGQMR8EgGwnRwCBCpvJfrKHGOXCnBptqZlJT9NK6kOX
Uz4FbjaoeRJWYP5xHW8b3RwiiN7Wqsq8LqNFSDc4QxvB4q8R+aStSc7UAwhcxI/B
BokMgeKi8wlMhyiCEhoUEoBp6ijhCVDIFOExndrhjU7gHImpJNSuk+9WYGpp0Iwz
7M3h4gnmnFbSC1ruZ5kxlvvlo9mBGf7h8eW+D3LVQjVokOSuj+cXJ+9USSJPp2uI
PcMFLCPZYdvGuUDzMficixWs3Lqc21t8rMJ5wDQuJpDc5hVv/5stsUjxttmZQtTu
OQF4WOQjg3afeX/zJ/905VKLFAFZmUBVOmA+Tb3NUX6BSOStsq0tMbC08zps17zC
N0nQ1ALaB6mYrv73ltuSzX0A9Bx7UPyLsUrEeMK5zJW0Lr93Xhjr1E4jYySO3FOx
YazDEwVFU1l0kRPE05oKntXvBo1JB8/PWTkGta5mowMGVHhQD0iFf3ZeRWFCoT0d
BlIQUqXdo6eTwDb8tL5VDEZG8fKmlwMhY299AA4/L/FmH3nJv0jlDmaL/4HDYEVM
l3xUMXywgHw9o9Yaa+KNgP9l0tX0bfehZNIwsvIxpzptseIFKyHQEq0ak2dTE7AU
qZyULqL9x9OWBAUH1yd7iZOR3kAHn8zTjG2IIr5cCtZVSWgiPkVEf8BloxoPoqSd
sMddr2XPc6pz2ZFhC0swcKrshvmAbrzia6wICCyi8cBQBixXsy3DwWEPWRu9vdC8
R/Wn9q6lcYaDcmoOfoTml0JbeS0EpToOBkjg/gZOGL0uy+9M/ZInMr28A6ulUwWG
sz68mE0RoWcKBHDFca09AZJnR1rmXewjPblCcKPjC2MOvyd/2OD14dvqbNkopnfB
MUlM7zMv3scSQcV/RlyRZxYIacDVPRUK3hNq1rGaap86locO/Ro924+VRyUUzjDx
IWbPHvLevGVCXwqfBXsJT2ob9pErpHCtDaZp8oqH1CQV5tm+uBSbQMxHGp6vQwAG
+9jTpVgRRtQXbted276i7YFqWYhsPuVlJr85ktEXrN3S3spi4hZDuDpXSXyjM2JD
yDFulAcReny2GWOx2P7oA5csgwMoXkb+4Cct47kmx79Sq8i3T9B2gPbfO9B5Veif
+HwTSZuMIOxRZEo2DsHQoa50goTF+EQAW2+VR/qEyXXlcQePs4vjpcxJoNXx0MGq
wKGbYGKv8/h/JNYrdDVGzaGNGKxWc1b7oJlBdU+N/UZ0Y/5q8hIyXR9Sd4aVNNzd
EgvviUCCy1qrASgDmFG7sEHK9lKLBxyHuPN4o1V/2TZQHy0DQnj7jVu/1hSqq/7A
Ksu7caIIr80PiV1CjgEaUMSmwfV7VYq1o3SUVxa3PQphiJnB0857CjBdk61/RjMc
oeKsCqkJz2IH1j4J0n0uw6x+OjYYBLt5gmDsNpqlrsR/JFwUFufiN7MeYhfu2sQ6
aIvA5E934+h8+YhHMpQl5TbPV0oT4mYLdzBmZXH22m6MyoEhJSputqFBeNf275Hb
BtH7LoZpQdyp6Jq41e00ZPHcFBQ1gkvawd4xpfV00IFjl+a2iE5GVBdZlcVKT2sV
yXG/6g+mDav8MXhw7A0OLYl2Wj8vu4WwXeCZdflbRFyTOMuew/5xxoF/zF9AHU2q
egXnhqCYfTbyw6HTC8z4KDebGGGGQKXFF+1v9CuX4scGeyLw1+tBN2tZ0X9dKGgQ
SSOq5oIyL02PRu3oKBtxwrbpXMu/RNTAlbUdzrKTDkUxZfrHtR+VUjYmz389a7kk
IG2P9ouL9d3/7aXuykOsLD0hL1zWTYtAx1QudOC1L06YvtrlwwtLH96XfRIP6IC6
lwz1PYN7USeCiBqOBHkerwcLgXhjMtNasJutXCo+bcwV/AgXaS2p04TYILlHtrYW
DLHoEiFJEbSJKwnjhATH9oJl0Qwc54a0BRPKicOHLINSU8MgTo1U3RLnGmvlHT95
RgGvKch47vV136Px0QN+PdjBJc2AXL3RDsnlERM7+YvgLcby2Htk1VUYNDwsdL+W
WIiFESXpnM6pZPF/ogRVF15wca6nNAVbcdzeaReG6U/xWwHIsEyaszO/h/6AeqJ2
vXQYfmQDQq77B9fDDZg7co1TDUOJCxc2wFoiPTIEegM58pzBICMZCQ07G69p/JZG
mOdOquQsIRfgj29evxdCOb7pin8Aisy42AsX2EJdzBRDncD5sNiM4rtpuXni167i
A/0t8VVflITZJD8A0Vwnc9ABVbrMqenhjruYiRJzPufEYaQ7S+1IA6k0af6gQTx7
1miJmLbgkmdlQpIXuVUhietupNaPoXMfTsExU730WzsaNT1IPdbh5y/FENwnXJuF
K27fetbxxe2Ew98KRF7WqqcFAW2EhC7pmdxzeq2RIJO1jQDQxDbJ/KmtKn2J5JXA
XsA/qhhDkSAObE3mniozTnKjdqdr0gQ56GLcPqcOi4GKmAaHd49R5aQcoJidftRw
chLtrJSMTZbOS1NbtXX8Gln2x0T8aWGDfr9jWdGrZEZjS4VXxBuqIpXIFgn38h7n
XulAsTDSTHRQ/aNC0dCXEfSoo8UyLmhGXw0oSh0l2J/lx8fSwM3Phf5cswAEuFVe
ERDBjRvQj7Xwn4/M4kPwepgNAj41labdwgpZkNH20PbEV9z3KP49cDmQ+HGpApVo
iX1rblxMuWxGZWrtyuzi5fRP0FcABALXlhiFdhYZ72Gmo+jasIoQKYMzRaQNTfT0
41DXwBk/QR4/z89YVp8hlSJnEpaNiSeE5qSefLtdun9FE3+ZtM0xW8LqOPoLS4L2
N06k6Nda9wg9gkMCMqS64IzaIXjhfruRCgguSF4/whKypaLzDWtrlV5R+0hCgFfX
LYkzIfOtwczbLIWqCJa/gYFmvVZ1D6Z1pQb8eQ2DFrFg/okqnivbHUMEZ8DZtB1i
31k9bC18qJZQnu+XnrSI8GjapUQQ2d/8h7xjpBbAUrhIQ/L+He+SkRfe/X+Kohg6
kLW1/vuqx+iBChgXaFUl/pfJGhAIz+qq1yHAv6pvLkBU9x9uVEQhCgWS4rbzi8jM
b9M4cXJhLYP+n9oKdxG4bpW3uE6LbdQvlRBpCfUTpgmtUgapAs+Kvw6HGfuURfZ5
RbmX0eQlBs9XdlEo7fEjurZJUHZZFUadLETHaauBRYTloXCLdW2Nu6vqe01Jj6tC
4ZiId0JkhzBKkzGe5kkprLnvc43jCLjJx34Zk2a8BG0nHnEyAvlt2chNS5pS2L9d
PtT+EfDxGcteZqwy3kODIZEPYl0zir4YZArPEk1AoxTX2E4rTUjk/O4G468F2Lwp
WE28NcUrChFKyl33gKBhIAUvJyts0J0o5gBSzt5ao2irhXlDJY9vAhxmxCjH6ws4
gl/ECFAI8ZbUO3WvsDLJ+Xk5ejY2mEI103t1UJn01AU=
`protect END_PROTECTED
