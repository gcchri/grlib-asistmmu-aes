`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sfLPgo0wihsRmJK72ec93JjkY6V8+0TDXUgAWxE9qLXRtPnFBkPxu87GFmPkhTJS
dpjTSbnOEYldi9BA9LDCttSqM6PLFjlWBakrlnVNdDyzkpfRUeqKAOtLosn57CzS
21edZ3rOq2+mNIdeFndz+6HjjZR35M68kGka7U8n9JSWOQSAuhFzV2MieD/X/CeP
sV0iyKafTzwmk2qY5SGAY5yRJFxLJpHMaiC8fkcKV9bBfrM6m9O1Y8PMK/cX9T3D
IE01inu5p/j3GlJWc9m06fr0gD/+KfzK/jB9XFgTeXOvkkCcXsAJCQ/xwj0oeBbT
A0oQ/+aTgmNwavEkxT9JfnSOfw/nKaKSUZ2G2tcxCMQFVqJb1EV0EviHQBDulbR+
j51JLRhxYuV5J9TNo/2kiOtSVvj7ZIug0je9TOWyfv1dCBo/fYyd/F1VFr/izrzy
S11/qhJOnkDjqhGOsKZ6P8lV+SXMAjWc0x2YpUNX/YWNd6+orVwUmXHva54AOJTk
5KF0PoTYFswpL9RUEt8x9Q==
`protect END_PROTECTED
