`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s+kMunssrXZ/l5dbrINV19TQBgZwKRewmzMRlotth0b/meDhgiHJqpI5LuwXMEaC
E2+jbZnE48pyxIGJSEFrZQ0OuvQY/y6Q+QYaMuZd8M9c/8l7zsrbRXBqCWNfRcFL
Q1ETYtAT5ZihHM+gcwmACSPDICQ0xReMkY2hSz8j211bGyhmJ8pOgRjaG7PCjSHy
v2aHPIQfSJcvnUE4qkkqatRGrLqJtvF6L1SrxTJpWsvRTkw5tdbe/CHkyYQ3ZhH1
XnxslTxk1owJps8bPCTP/zpbqHiKX+KDvAiu4y02hsPvmEjIJQYfNPLWXSAHm26h
XpoOVEBqVMz3QL6z+ceD8Edg1Xa8QsKCupx+EHYHwnuxp0gKDcI9M4FzjFrgog7y
cRELgVsYqn8cE/c+tDHFUN/uCOwS3frV6xdAlHVZJB84Z4iXm5Ox/uYD0oEVZ1Kl
dHCmhaVkKVjdRJ6vmmj8cw==
`protect END_PROTECTED
