`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8a6dJlxRRYwLEqJV6K3oDCDlhuBj+Y93272hUCi4NkPBv7zfOZ8EHbk/0d2Rrtns
lVzekf7No/n7ZvxQ3ccfrkNY3mwlqYNPocHvtyuRlDjapseBsLOhH/qEPkyriGHZ
SCCnGF9GuTiJRer1izQHwpQLJ1jFd1G0dfX7tI6nxDK/1VssPB1mIoQMajO69Ez1
5jBGfRFvWYN2ZENOvGX2VvaMvSYpUJ/EEWgzWpjJzYPndQrS1xq42Nj/ACS3Lawt
0IL8ktqK9NTOhUZf+0SZ6csFBM7aZheq5Do3YBc6T/mu/dDNkHDVdnrqmJ4kpreO
M5FsZrrETa5+1jfe/XRWiL0cScbgS9NFLl4Iq47B74TV660bH2gzET2g9NUXONZr
VUrXimOQZYXj42V3xXtHBQ8xrKBl48DEtke8MXB1O/zDb03o3ejA6cSE9QAKtjNV
l4KLG/KaLCjC35UMNqItqiAbadJuXEz/WNv1FVslDvg84ThBUqINfre/OP9ML8tG
XmbPz7MrZeUpabEX5/oU3Jz+tkeD4L5gwhIO2vf1Bzv/ifEqh6UOY72d63V3hyN+
A+tsA95QUvKb+EFsWh4ICX3JhfeWEftNrJNp5vQqPuh1mTaG/z2A6dtUe+xdwFc1
0TTVqXjIZNkBTZro0/5yKA9jxOzTz0iOcQHjBI9fBUcp9uRvoEwMK57nFTKpGLae
45Hm28M1xMy7AjOzZJrxeLFO3y6nHS07IpRdIKmZ6Ak=
`protect END_PROTECTED
