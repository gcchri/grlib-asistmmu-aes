`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dFE6cA3xJafDSLFhJr8MKDSgY/ceFyE4kofMBhRRfo1d3jbR3lHgLFE6vxwK9Dcs
H5hBup7QBJWbW2yL8mKNC/sVNjUHQZNnMDeWVUMJd+SDYGxytvBiAmJj3ApKuSBv
INN5K/f3OphFBkuixyAcwz/mKAWY0a81FyGXwbnmpexOJkBWTFMaxdQHlWqGBTy/
DcCTlYu9fBmnKIHnxCgJsRAx72y65cXZ+wRzRDtklFTRK9hZi1ceKu3Uli7CrEO1
+xeD0LzK9vr65oAqTbR49rm9rPyahl/LJ9FW2obwySXVCcuHBz5/17TvyG5bipAp
hjlVL7Zkc4dve0V12HfgtLhHnmFJ9WfWegOTmHeJy/1mOp2eNdvXe3vSQjrxxvqn
CWK/AvsPB4ISR1Km4CoJPanghC602PWTLozHB+cXbp4=
`protect END_PROTECTED
