`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YOmQmivnZ/7xG5qTPw5aIkERr53sFAE5ogWjWWlNBlupehU2Ja6ayohzxkXlug/M
TrB5zlX9YBx4TZ4g4KmaBy8/GhEF1xEv64cIZRXMzT9i9gkiqgt6y0stfAcWMTkF
eRuR/06Idd3WA7RW+S795spep7D41a3CgxefbgMLWfMPRtHkxp4FoLmMVU8/taSy
Gd1MHAs6yGTV1PmvBv9X/fP0otoO2t6N4/rxtUKbRJI4d1DTsNARcCIo0n+BOoXO
wJA0qIX/kF2OmOrcdgzdiq1SbpDHAqV3LEbn0Jg1EN2UpkREITUwypH/VQsQdY0b
Esxg9/3lrmqBk+KiGKG9gA9oUKZ45T+LN3Y+04qnZHSMFw3srwd0o9X6mIPhvADA
O0sW3izTfZa0+izJqJSV8w==
`protect END_PROTECTED
