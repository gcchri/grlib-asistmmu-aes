`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bQ+6W6JX36hA+AnWHHtlcFNx04XAEISqlKJjhH62K1HFOrWgA6ikn2tnGbsJVJNB
45weu8MW2ZpGiUw9EbXGkYIpoG+gRGjATW0fGkk7pUtTNV1AOyCTEnYDWrLf0Vph
7bYawjsiWjjvxCBWqTW6LdjDdHDrGVuJG6Vheo3WaCy0ljxatbROwrSN54lGQFyx
OqJliq+rIA+iYhrNUlAfiyl8QQ4+vr+CBWYbow/rOcXiCOPymzx6zvxlR76ecdEP
sqKrzvwI4wrVfktY9uzDy1TdmdzuY6/kwj3/Ao8nL/aMjUcuyf+g+51Hi7cy9t0M
VxIzwYyF5+2zYiF2jNgvBJsa9cRvm0zjTodab6yc9W0mk/92SlEs38dX1iluHee2
sreUBI85aXfwA23fb59i4w1M5LS+wtUstNfuD69hXcCOgHemmGUlIQymDKqevoVT
jjFTLYNp4R3SDDHpIAKSseVNwEilJJfoIyk8u5td+cgJDqUOFrFM+8CIkyjrATl+
PmTszcbFvVcovRDhoW+BQG3SiSWQdT4d8yxY+WmQQvfcIjc87jRE8ir7J/tAoGjq
dCMIoBi6wirialIwi0zWhtq24YVsLfITB1fy7bGRjCdDYHdNCsEgzD5yBuaS1uzo
uE/cHteeQogF2cfRPGWrA1INDzC/nbmSRjnZqJjxaxEX0Rn/YgXahWB+WgzGf8w+
l0GmHMtvaUmpx7jMq8t47Hf73qK7sbq/sAWvpav8RJh2VCa0VpAj9A7Yq3okSt62
o0nqlqGTnOn+sx4z0i+p97NiXrAgkdKNvaogt7pGNQCCYo5jYb7rCOxZGln9C8BR
qkvwiWMnsajivYNG9kwi2qPdQo8Yq1LOn5MWoNlMFxE0BS6i5JtkfDvk4JO7xkxL
jo69iI/BLhjvVPY5Vu3kKriBvLBGj77ol9Ii83himkp+a96Sd3zfWnxACsKaINlq
7oDpkPl/ej/yOS2rDBcOBSi3MThS3Gpy1kRJJZ9ogkseSK+XsMkR1jA1T8cWDQQo
Rm8p5DieQ46nWmVqS1mlL3k6v6GNGXj+bLz2g5/Pj8BZXQXGudrYaeryljAxMgrP
Va+GCIXwvBTS1QD8ki4m4ODZ7T8KCwCrrnxwr1wCn42XWRl+6zufshjhWeSfIcs4
BBTgTr8gnf6h8dFsJRm5NrsQ0fXb9niscvBFSn9+QdBnbPkSrwvB1dDc+rogoRTI
JCuS0GcXHA+BpDy54DyDEZyckTRcu/jKx3QBPYhB2iZYV/SJQlkKHD+13x1nl8Gt
qjRhCLBtxvT5Jai+smxBXISCnpF82BALjaogst3cJu/0eRVV2Ybyp9B2FdmwC8fL
cIXDM3glPlJxxfwbzpzm28CI1ECv6t7F49ok3z2mS7gPqIA13rJRJlYPQb7QXBtt
wUv3kEeNKsTw2mkhvJFgAWTq1k3RY9/EzvXOXThvorNAOCjHbXEMS919lOCJdM93
uVXVpk46Ioy2jS/nCEMPSHWYgq7Ln8x7oaMbH5aC4OWx8uZabEgFNCBcJFDO2ymT
USyFnwp62Zx9J0tS4DZp5DlY7Ash0RpZczW/jMAxaypp3rHe09g6AhrzwLRmF0ZV
I2Fhzonwjf/lIE7ju6z3o6mMDTrzw3kRdL+LoFqRxiFLmP8r4OTi6MvFgbbztvZl
4loNxZVaOD98+2JwqItEFMj+MnRoirQOH8im77Yz9lzhDPJPaIwUy0ejia3+Umv4
u3eBblQJjY30m7xknBxWs1zfDf5BTYK7R6cCy4BNzwd9Tvhm5qIzEGXBbyCwLHzc
Q6kiIgwgxuVHUA72BsIiD4ibfi/nYq6Y+sgg9T9KOJEvzIaBGw3YO4K6nOQu8u1v
QNOVeOwjMLSdVXOdZqmhx2sx4iNL8A//qvRoCBEgCuTxNGBADpMLv/3FgDdsK3bS
Pq2Rb5Ujk2VwVfTA8HnDeyo1e9sDpq6gk5c1hntYXqP50xw20OoDRrLOLKQYAwym
GRO06V6Xr+y32LXCWhS2ZuoUo9Ig+Q4Qxm4GsJOrPDWI5B5SvwPgAQRLS7SJVFqf
VN62vL6PrW94mgQgh3vVB/xBqnZAhU7JkopDrrmHyeq6Tygw1G6yLuh4RLuQybCr
Z4m/ANZM0ueIsp1dyWRa1nPnra6avVEA50LQl9urpICse1AqizEml/fnlYWzEygX
zFU/cSTmDYsfdWzC9b/TC5aTurVLCt+alX5svN71iY+2lTuPc5HDbzlwvaqOyLRV
tKNIRjIZuLpQAlzDl3DyBI4nGEe4Q5In0aRvacWhIKl02NGHGGY3DTbAtMq5Ry7q
S7pkg2OClrLN2XCyMUuSPuxlgvYXlOcp8TLB6u4sILyPPG+8uhpfiwkYru8m1wfI
F8jISCkXwAwVw9+XoW9nhCURc+brN8O7eygCjEgj0Fj5m4ruhXdli9TznZx4SAKh
SoWIB5492N091KbFpNSuHBUuvOt4FviCKN0yiS/rtkU10OokIG3hMHroEE999iLh
k97VzHK0GioNSnTe7HKdWUi2rzJSN2UfF135A+jmjfFSm8iQYxVPDMPSTZ87WlK4
lcGAaAyH9PqYwip47Z9/8QCVY5SMkfrU7MTcl0KIPDVt2qO/Q5rkCMUttUTmJixx
tXamCcgA0hVb/l4UUY78hhjZcw8oP/t5aVDkrPl3c1WUHKJiWWkqExsCq0lLDFIs
TsaUlBM+fXwYmr+rCB4eu2hmHIgbPYdkxG5d8avfbxA2ji2ugHjzRfpeGIBztbbB
cMebHTGqtmfwFKVdZd46hW/LTLmYbCx1q/wfeg69uRj4iCBSd1ksr0LZeO2skmBW
t4GT+vfm71iV+bhw3JmVnCuOucll7YWMnGD3uhNvSWF2dtNKNybpu93zE5vXbJAX
VS5CXTE4w7LMDVCVFnxEMUK/Cx5kyz8RFUg/gCLhuePsYV60WRNnTIqKFmQ/6eju
rvoFzLz9z4POY4Rnq2YvrPBHaQ4livXon5IcHPRymkkVPCmjRxEDFIJSHmT0Q4sR
Yr+iLCiqSoZXxf4cnr2KQda4s0a73WRG+s3e6s2u7sz+3Uf/vZ+9f5cR2+t4OKOL
MB1QsrviQVXS2c1Wo7BUu13AyezVTdgCpdLsWgXiTWmQfJb+QrwkYVZ6W9s3FaBI
OOVvujeh3IWlfcsTB1NqIl28Lxnlevvpi5ZgmQzuYpUn+76v9ifM8qPQv7d0mKjV
SEKUNP8EQ4hZPv3TPmUcobcYhrzXJM0Kz6DLPynRSwZ1f26LgDFRKXv7DkbUmIn/
grWBLEx5qE0fTp7lkM4qOvhJc/UB7wXrz3BCrefo0aiukig5LhARVPyvEZ31PBw1
YwtGX6ubOkQQTMuOZScIdWxip8xA6KUzTmd00EhSyXQWGewaaIgpvWXvqLlDwWwe
za8rRpAexTMRh96yiHccxZ220BIFe4K7fmiHVDSW/jVak0J5+5NkvD+mItkA3x+F
Fj6sciiydPmMVs8cgjqy/mY/jc/49Wbeu5YYEob74+lfwkv+/fLk6iYRA5VJN35r
sHvnT3PKEma/tJtwEA7aU7bHoc1wccxfsofmZSHn7BgYhM6+8U0vGsbK5eohy91C
Z84wxeJRaot3Ea7yHCE8gQikT/QoenMC+j+9cqo4l+wCMs9OQknMv3qfOLCTw1n8
zSFPGjMj4e1rlOUqdNiDPTm/3Mx/MSi1Rv2k7PGP+CCJ6Yfd7pcOUJepehx7F3sp
eNzlpamtQ+sfSAwnJQ9OHRYogYKumyBIET89WdfdBd56Or0XQU5Ni3KEMl10CkHz
gzSuflFJ3/1GlVw+6kViuyEpsXQ18mkznWopVvieXrdtyxbmcjR1fWbwN1RqibO/
g3OMbYj9vxMLIxM/CGeGjNtf7BpZwLPeY0kJIE17IGcl9loaVCvgttrRUO2kGolU
STr150NcnyN09hpvIzVW5hCDGTd2W8aNKK9vUkgFvFZNciWyALmDP07ZFkPBZvBf
Ow/m/xS3jxuvA0lc74q1XWAk4yCA5dVNC0ugBhRNfr1a0wh5xYTmqtE49K24Pcj3
U7LhCsRhOpdJ8RYCnzayIXwOt4BEKqk3KB7JA54fj8QmslNrGkSCR65GmdLubCle
/3LVriVTNzKrmvJ/DpaEfU8U5S3WfYwVwJGhHehZC8BmUKErGNPt0NOKbHzmfM+B
WOua/ws3ICf9MNcKvWSGJCFdTs5GEhX04HHXCwmO5K0c+1adYw8qM/NcExY+rXVA
ASaqtJ41zpqJdgvgqbpahusJrBBeEuRtrUNrvd+2v7RZr9EY9cHL37CLrhdcSEl4
ifO9miHZcBOSM6qIW674qmTiH2nbgaqlIj+2lJ0ZjFbYhqBkQz6nE6MPOiTESaTA
I6mbXxZ/aUQG9EsHjshLpORlGcyuvSVliKM6V/gjk8E2pJkfgHDDfP2vSqJ1/Ier
mEEasBPLch+oJ15tovQ5i6x7EyPPN6ffkwWWTiA+S0pFAR8TAtHXeaM4bnZmZh1Z
k0tveh6JK5P6U9nCwk43BcgwUxwtguUuIF5qg+jxUbBjBvRVq5RIF082qU/pegSN
RtN1mxObum60FVXcttTYWA/F0EK2TVxhM+jLV27ei0gZ+eMxsJEtn5Dfujxm3ycr
PcFBW5ZINZ/R9XF4cJxu+RjUjQ9xfJgGO8ysW3GLBXyedbCVX2Q0X67coyWCGvZV
vKR97id/BPPAGKHjVX3o6+ot3A02mwh1mLUYNpJvptSmH8l2eLj3Bs7e17pxSUZO
zzfq2ZhBsr1g88TsXcUeVHIzUFgbpcb529jp9ZedmkethlTjPlJx/9arUq3ydeTe
SGVRMrWN1LqUA2pOiTJng4jCrXkoqZUTIyYX0Fg7YFjGOD0k3JyhYIM1A+246PCE
F89rdZvwoGpt+MXoSYtJXDSXY1hAuq/1DUv64hIiSEiRvWC3KOKW4r1DFfd0E/Q9
EpwxBf6K1kuHyjYLOMcnNZaUr/NUkgsM1Ut+rgSaMB1ViMmnKtl6Iwf7HPKMKmfG
Dk/qQW7kEKugE/4zZz6JSkARnnO8icT9/sXI4StpSrlNKNSFuX2s9LxfjtQzzg+B
vveuH9YGWW2D5TH3uoBW+p0YnaO9+XDmzWiVRqDN7yHM19za/UEyruaPGY3QVVMb
z0c6bCSD2IqMTifDDBuZ70jfTYbbeTz8LWpScBcXDlzxsmxqK723JmKBk3OlFnt9
OS2YnWSAQpLdBqVZhlTU+A3wSf1M4EULKN9c2E5CUGcuI1IDmASpHfqronp6+WFM
KYA9fibUttkCsvnxHn81bprV27APT/4lB70gBIwyoyhqkMk1MKm0NStp5qgscumV
EV7pOweCA35Bh54h3+xI+AxfYKfX3f1XcVv9hkwrwmpFOHMZqZSZmDLJs8gt1KkI
KHcvhAobhlj+0BdDwwSCjvsj5Z5ybG458yOotR+8jJVroxRM0OTvXTfEUJClyZZS
pHE/s8A3iYXXx/z0I4zWHbydHg6ntI9bzwa6+TgpNy7au2nsrTzCRtIVVakLQK8u
EXEmLLTmQmjeG2yv9BKu7/9KnMnea8zmChoF/34eaJw/VXici4ccdx37JNd8TKXf
LUQGEqhwHdzkan1U6yCzWNtXtKmNeYFx9hL2J3SDaI3IFPmrTrCoSvzYgtRO1wtQ
izaMT2MzKXXyG5UkDM57Noc89Eb1sTgkquEjwbxNNmn0FpdfqR349OM17LfcOTAf
dCpQ9kXYGzogcLIh5U9/mSntzzgt9H+p97zO8I0KsQ34xXDIwT6OH6V5tYTbI5dM
Ogm05+mIgSZC4/WjFYmWV8nIIvi+Rop3Li5fbnU7cvmMqW68u0xjcQktdtZyKPe+
hKW6vLDqebdgVqOlB9Ezq4jfPydsi9cz0xcbbHtuOwP3IznQ7Z05rdpknnBwYTq1
iUhiYok77fhMEo61hu/r+VDCH0ZB6qHnHkcz+eRg5qXUXSoZDeA3R2MkK1+iJcRC
irb5XOwRi1FdOX7aGQF1JMvOPVz2qd5karmzbEyJTP4geNHXuwbSl4yaj8gHWENq
7yIqtxmiOtv0gg7FRHYhfDDoDpIT2TfPBc/LJWz382XtBIeKdlnnAfLA4eqOKc8n
UL4jd4orfE0zkrJ/2DQ0QJr6iAAo0ai2jHkJO7MohvwpvGuHQr/P6fDdce+buXWb
2V+PB2RbV9ihqtZkqcOj/iMrNFLMqSUvHizSyAP4ut1KOgn7ZnEeRwbAfjw3Vi2R
TkS79UmUogHx+wCG/KvkQUSSYbXDdEQ02bgPLktMdi6VSUto3S2bhFmc5nS28rNC
u5tPCgQfws1MdPX5FaoaCnILz6/Vto3vr3jgZJcpyuSYuMEfzvoMZehBYiBT7BdZ
vkdWEbqQY2C+RtWKn7fcJyqmBZrAIMlH5c1Mz9hUxmUZcbVHY3CihBJgMTdRm8Vb
H5Z57t7YAluP0RhPdHBH+e7HZgwYTQTuD3QR6CtWwSEW4FX6wO0A6zwBvTjGaZo5
7qAjnqKGDN2ioH2CQ2jOxezn9BwxZVPf8/kPeLDOgzHnGxPO4MhPV83ivdIYScRT
cfNJYFNTvR4OIAAt4qodoOM3umKAjF10oyStlhov7SbOhI0cbEDhhMF0xns/KDEo
tnVYOC5IIlpY2L9+0K58uZpKFT2evSGvuroaY2a4qPzd73dwFPuFNLvS7tkWPPnf
9X+CBViCeiedw16O/DbSZws3XovjTuimcu5ZHR7koLDUjMB7fysqUjn0vggI225M
ex+jTMljNfazKKz5wHx2vIu1RzP+r2dYhRhaX2AT/m/6oAaYk9amFTIx5isHrKO1
Nk+meJ1J+wQA7xc8TMuWRyYHcEjLqXCFOXT6k96fWjuCredyn+Khkdzy25uEgoyD
rR5pt7YvlV66Lbn4WzNnf0BH1ofwCrpr5cRQ8Mevdt+2124hlT4i/v7kHSOJFSzQ
/QeXORkseVHML54iCCLdecz4fq2dBoQ7U2gvSN9PGdtTfeonfwID0JvAwJBNTxCU
zOa4KotvxTsVKMQnBKP6DckxxAokTUDDlZRzd8ErM2FHOnvQ23eIlcpfkDTWnXg/
RYSfSqVxcWEm8siUr2ZTq1xiLut2AuKJTMvW8toTHg9xWQpBLIMx8xCP/KLxocRJ
7J+HY3Znzafx1OW/4udSQOydjr2Er0YnaWUlZq9SegtM7bqmlThfc5nxyCxPlKvh
HJ6T/ZJMRI04mQDUxPjRH7gEtL6d0R1BwDBXfhD21S8eAXYkwlj8IGJWjHJX7W7e
GqAGI2P6PZozD+GgpYIn2vKfv9cmdkdRvg4LIa/s1UFoQtbhhS4vHX/tPWODN+Se
KgB5IdBLST0g08VwTYg/lZibX/YTZ/0c/DSWoJw2+1WUab3oywf0OXqiV4E5SBdL
aRS3HLshnz6V7Jfm2ht46VapdgSu3dulxnJe+va9RBLVdcpk/luJumbBc4fuf0pk
Z49R8jOzoQsJu4ZDn8G6XebiCr7dOfSTAKzCcEtTDNU4LwBatnKjQ1q5NrwxUYWb
cvm0axQr/3aA+pw0owbfUQzmJ+N9zTTmd09mNTT/KjWW2q93qroW5AmWInZQ9qFw
prYyyjLAkXwHoiDdi8TCw3v+cDZGejoDvEqF8YSfSwq5qp+FWpSRajWJeHylATQ2
rpvvh6TDS2KQGQWeq30qaIU0zWRg3M9lzB+WBUpH2cMnmM93kAgOmdKsmzIStgrh
WroajWtMOkiqD7ep2/5CLnFa51HUgrURdKOOh+R6kTDrqrv5384Vq0kdnhpIsfEx
HbouCiejUuRab42m7Iq1JwiSkInWDS03xfRVTpjjjMeFcCDvWn8mMJImIeQTBPor
1Kfu2x5mF5Pe2YtB9GW9eR8/SC41vkbrvw3Ckuyvy0sS20NC8bC99Xp5Lz2S1gES
p3MeT9K6YEEXvyPgcu13BaatBJhVCSXWjwiHsirwarqJYgIKNXrvUklsPd6meRFK
pfyTLd6dhpfSwXfkL7oxzg3uoJemBH7gBRLiORSy0Jz2T/yF8APyYSVXQ+6dssmc
juN8uUR9mJNNDZgtVklVfpcw8bNRMzd8Wq8hPgvEkaw5kfEr8Ft4M+h9xB9MTsWI
9eR0IEy/U7lEyDPFsEl0M3uRhbKHLpJWNbpkOR50GTmgkZoda6m5+gEUvqxCqgMI
x+4lgc11rKh+LWDgDXQs36UZ1f4lq9066XA0StjumsioMtaWLB1yhWe2EXSGqY+h
nuUF7YUdlxkM1owgl7GjbZ6bKQnYnQIx/FLWkFxAtpapqGs7Dz4TVP1dh4Nuoxtk
mVZPFn6dXinpyvu77+TIEbNRfKGqQJQWiIXyx0dmFG4Q+oUotSImaT33ha6AV1Lr
0Mb/CzdzN8fFQwZ0w1ttVHRsZ3y5+6yOXffF9Xk7v/P0go8FFBpv71tGVxmDmLO+
/qi0qlrxUeP6uGwsrlVDMokyMWT71RYHA9h6xicuWFEzzhBdc5HWq1G2juP1/Jkw
+0gQ+PefVseHoWnWsYRRdl3u5ppKRgwE1s5dtjaD2/TS9eDyjG1SC3GafxcRhHsQ
FI2oSqbDj/1lONqsLaxXjpWk+gjVL2sAugGfNbfuN/0MchrpzQ1FjABwqQFTPJYA
XL4firspPfHwtv7OLxfgCQQF1AeNykkoZDHFpiyXbdFQaQeOAxn/lqWcPH7mFlHu
taejtxxRCRxECiNeDBJZu+QfeirYKC15RHp1/HH2mFzhyhg71G09tyHSzBnYGorL
lyDBTaRUhSyFvoZ7Ec/qcL+FkI2wf14QMpRDHgGhWE0pLSwPDHCOB8EDnwElMmDl
iDlns0Y610vVpTnLg96zSBxtQnBUujFrnSapdV3j2JvO5Zi1WgKzrUmfkzpWwfro
p9nIztZVE5hZwIUokD7NoGI6jla9X/QmBk3wheHTfFffacvGI6NI2E5c12FBvTT4
9M0sBxEPolnH0X/JlRGIX/q38zndnTe4Ic9H2P7C13k1Kqpmu5I56/GzOad0wfW7
h+gZHN5MoIP/V5mW4Uxceu0QnCwqfWtMN3AaQTwwFmYhUU3lvrTCbHss7B8NzKAx
Dz4VFyQeimWKQq2ty+/ZiLM6SaVt8b+prz/P9OOLOYBKOSxqEfLAC0QhJE3XZDMn
qNxanVXoT9UF2ONlPI1xSQCo2fi0+JtSAVDU+epZVNJ+tcZtK5X0+2uC3nmYztKy
zXiajVhJkep0+sFCTlhe8+jtpQopN8rI7hgzdvJ3IW7paHdnEQw/zKzM6lOLOFv/
KettPF7BWdmtr28T7qZ4Ga1JC8cNJhOW1L7Jqn7rWx1JNYtQvvlARPWs9iQ/GmtY
wBJMqAE3+Jp8k2pilckYazO54htflywOiHrOqjX+abCCDgIir0si+KZhpyyOwj8w
nFdlCtpvvP7xDh0iPfeee+N7ZMm2f4ZAoldwtqmMKWn6FSQhwcvqM4itjl7cMx2N
QzS8dfgkw/MnAVZsDY725YXP1e6RcA3pk2xbv9dmdk1WDCmkRd8KJo9DqR3/oyEz
z5rj740GkrX1+xnxFRdMZZU5md1S0I4eik+3tpdnuTa+iF4GNKuSmDARG/idlFAq
lIKsQjjAWh0kmieBncmWmkKcXr3cSKek2uu1noLve8FGl0w2DMmdu+FyWXktME9m
9SwQ+yanHBR95FzjlInpZFQnkydcJSgy4Z4gAa2xTAKn8iU0KM38GP0RlLtDhGfr
zMVeP3CUkiNozCz/RCRD8VlYEgD71Lm/NtfgkCuCBgfMQ6b2MOBAIIU8DFY6Jj3A
hSH9utjZXtrvW65okMg4hTdKEC/kzwK9H/sfB0QxoTNae/ZmkEe11zisCHkou9ru
3OMrPshZABCu5vSvkmQMSqH/gQg37l+AcHhzegBU8/kN7lP03T2dJyRUcf9TA2hI
PaTiF4eNek+Kj50XuBkyezydvwU8NvHVbYK+NVX+dX+RxZe1w1Gbq/5lCueJ4TWp
zxvIdZL9aFgbSvHbRc3HPSgcTf1ad0U5pVaB3H5QkfJib0L6fhZjFceIwXg+Rlqz
5B8gJ6HhQ13/JPdQ99aJ9iWhHRRvyUdKeT3hRbMl9evLxWLQcjbNrAoY8Whft7Bx
MpCEFNNtoGB/LcH60htUMwN2q59mgKl7MfUdypXhXB+Cf7ki9/UJ8xZoaUj0jKO4
BazHonvWyWvDb6nlPdwFHS4ZAPDuSejNq+xYy5Jd/tIaKep1lvegWYB6zFcyHPVU
Qo6deE9vZ+IqaZUJX7vQWdvK4Vllw35O/Jo/S76j0wGziJRZlm3ZR+ShIOLDGA/M
WU77r+uug8hO79p/ZhNGDt+Cbs153epYvBrQoVRZxvaeuKFgYQgSzVYrvj7tjoeY
E5nsHwb72mdtyyS/SdPJevXfH7Z7YfCGJf4bEfVoMuSCd/Rsc9FbZhj98QJ66LbB
RlwqZPV2we6r+NoeDA7t2fvk8siFUulos2zE9jU8aTP0f55n591SvxkQVPAHQhXR
N9Fj29Ft763HWbSf3FJ/4Y8qbU3093Lr5zLcVXDfa0xuEIVTPlztXuACgoUvuiRO
PsvT1YR+zvyPK7pEoVwSE1Oa20HJUaYTlsYrdrGOajnGLCO1LgwnXepbwcfJIQcc
Pjt+8jBpjkt/Mx7U4NvA8Q==
`protect END_PROTECTED
