`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8JHHayC8bdA+l+OscOZg2U89fLTC6cKWvwwnDq8YlMtldZHGdGRgVT67mqMtKBt5
UGKzkRz4/lxpoGu8jRp/X1wdAarlm4Q4VEaMBQeglOHUifCB9y3rPsfXc/S3cSTN
K3xU3BCIcr2tLMQTeGG/cEZwUH2dFltnL90RVJYhiK7numaRYUvDf/Njtc6z0obw
0WdLWoz+G699KHHgKJ/p46yOTJ79dncqnVN7getILg7//SNqFgBwSnh9uP/dyCGj
Gr7E4XRUkmfuzf9HP+HniZgoy5WgfvwdcXFDZBtiOIn22DdupdENyHFUo2MsF+Ns
WPBgvq8V+uUVRe92pRPRNONWPPJ26iz6vZWe/isny2lxVc3pYtiIPzLDAHsgXZY9
Ya/X0ikv08vGpJAwttpDwvoPt+cQpoY/UTAGBrJBsjcOH6aX2i5AYGsY75nlBARB
W8GH7fMcXfQWnmIOu+zeYponb58qhEWyB7zjg27eAPVTyDjx1ZNj8WqwuJMronTP
gguI+1yZrv+mLDUL4cLa/VQ0A4yVfXEtTIOyeU2FYGbrtNG9lzBKocLpQL0I+UFk
m/wGdqYh0s+gxN4DfwHxBLyp8Ze1QN/JZf9nx/iP4WZ3g+gVIj5zkaRAeX+VJT2H
vnRvPY9o1p6Um0rFeym+zlVnDKH9eTPXqL8/EKkhpLCw7UU4WegtTVhHd8F7+9tu
1rjg0vtkgVl4EIRXEVfn3ikIcDw5KFwBDS+6IpIlrZHsvTXXbA9Heegj56FOf+5h
JCccWwCN7yMFQIonK5g2RFVZCQWNNXNawVHhD6m/bVpakwCB+feGHjWT3kQI5xKx
bgW0aoGCfOAuw30FtcJ/pmhFX7PRvMusIK8nOzk4KUj/LNAnAbWVbj6+GkkLcOGL
HRpVrwBjbukg1mbOEp21VXUuZNF55jp/HwQF2uoKP1gWkKfkCpy1JKhzdTJBB5JN
Ps22XE4l7FB1t/vnS/m2lflOUvTuftquIHEBNA3kGx7RcQ+9JyjVyEtcbAgcaLXt
1Kiuh9izrtL3/TMM987XsCFX3olMBYrdTRvy2HjPhVp4uulpqUalyOJoTBTIwE11
wmWFJVsMWyFzI1r9/XHx4m0989Ru6do1F7kf5dPBajHJIr9zslWoLBg8AhC4bVOK
mFQAWWMfVtyP/5v6Y6yXWDbAivFnWczjBEtkgOgH68n9BsKh1tgPPfMJXF1fVQ/5
stIY79ZSGL6+Sz8ec0Ze+EU7RH+zFdj64H8zaOaGsisDGQ/aZDsDMdqAZNk+nEHk
+RuBxmF2djpKv0DgqogmvZiGQzAkLXv4wipTRgtSZpI=
`protect END_PROTECTED
