`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zl1B35TaP8i/YwkgXGfdSQ2e33K7B48keD8F/Jgm7hWQXf9vIhHk8zP4QEn8zG/Y
kBnkgL6VBU8tR3sB7V6NvOE1KhpJJQsoPKgv68HWsfx9lZ7wbi5tmu0FBEern05F
XtZpCnDlFDkwSzQhfpKD0veB5OVMK4FbHH0blLvn+G6ota3nyFbIHkD3Ynct7DVN
35Hq6Gf/l2Ox/QOzdghNRW7/IqgPXv94gjzhmuaytThNCYsYuS1a2o2c+hC1h4m6
sM/Szzf8XmSyj4CkdpNzN4Yu+KARLSzDV45jD0Yr3c5ctqQ5UC4MwvoWfSNYjTiU
sE7uNXFZ3mmxagkRH+tg7js1i1WIL76O+5cGA9Fbo+s5bLvarJxHWUhvKS6Anmh8
Q8nZI1hx+4ULhsyAluhqZnzkyCN3S0ACPGL7AR6XWs+D0R1GFykAnYJwZ2ktiw8W
iaeM8aB4lwnIaT9U5cK6u6j/ETDuZlih7xKIVy6+t+sAfHDJu+dx+OZ58GaMK28p
`protect END_PROTECTED
