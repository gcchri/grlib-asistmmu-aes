`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4NwWvvC4GSjDDkxAizAublt5QNkpOa8B8ARYN3tSYPDheLP0lDcT8f4yHpxRcjRe
VcLyHOeHgrwmj9o8M5i6kZTE+i8SI6i9xM5Z9Prpb43wwXPvmv8jekWR73w5d/BC
AJYHCqGi9JItH/qw2wcibjLtCL0gPFIQS4F+oG1Ij0NYnx5+jkY4cJvX4xVz2e6t
Tc9rQHiku2rEEYOiMj0gY+KU+5i5c7pi8/qld03e28Gz7Q0/tDT6erXxiBXflpQ3
EJ+mjVbwinMozaz1GMF4qfXhT9RyWbblSIeYOlUMFRhBMs9xuWTrHQO/knGbxWYx
UqwXZuzDuOskjikcERdWijsstqASmS7Q3wS+m2TbHU4iu7AVdfp/w5feh8/7TnLq
Inz4iArZoXVe25TBKufviwrpc071QwHZHyrjiDF3H7QTsVyj5w0PJi+jETtBk4dM
Y6YHpskAsHTuJcJlek3k8SKNE4VGr4GRvdqx2GNHumJkH/Ess/bCXwJZdDi2H3h8
`protect END_PROTECTED
