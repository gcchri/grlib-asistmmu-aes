`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w9EoJcBrFDVPPqGMhXjly2m4tUdzxPbTLfQKUcqy0mg01dbalS+NO8b07AN2ZFlK
KetomK9gv97qSQ3z4geWKZaaUrHTJy2jok9wivYolYE8pl/RAoZyquS/a1s8Y9Ym
b/W1tfeeA9NcTdojirS4qYsZkd9kJaAarCp/rNE04NKYM4NK76aAf54widqBurG3
ZHgk2obZwzXVl4Hihy9snOUY8j7BPpN+RnS4LrNYhccIwNSzwJIXVA9wr5TpfzjL
wPTVi3eWCiBYngafoml55w5TJLO9yJJQRhFL+5Lmnla0OvarahANCKhYbLmx3MYT
FcTizd40bKtM10UJaNKNOet+U+xB48IDM+5zKp2buFzlADdMabRwqz9ao3GCA9/0
KTQbBgiRBLtMXJmhUDU5ndGOlpcoITeNhz9Gl03idls/5V/e5RadaTASysYlBhvl
sQ/aMZH870SeSFuSUn0FGp9hf0iZPJSSwI9Q9/+6h4ov3t6y+1smr8WXai2UVncZ
RYL0/cHfdj4TomvGhm4VpeMDsAbAFTeGwST4DoOCi6oPGVlWHBzru4K+3nMsv2t9
QLxy1rVqchPDOJMwJXhZyPchSPObghdh81R4jZqiDgFK/UkpNIrzVs7Jm467qikp
pAzj9uUzrQiYrSYkwi3h6qRMxjNZIzRHVsmw+E0L0gs2UEIqoj1Oo7ssRPLmKJnp
ye3ukn5UC/K8slvpl7YqJE9RbTLd2ScHtgmXbcDpPom9/VHUiT4FvPktc2OtDlFk
X25X+0T0SwOCzbgBSRwo/5tedgDNb/7+Doo9vzk5wse7r2t7BDasTNtFBeVYJLrE
Y2W9FYDuCLRAfFahTS0/5UxagCyOKgaXi37c6GW8hNU9myan1tcsoruQszNgR2Dn
yX/zy4yWOONdgMRWOSA2eDPPry4tFe6Guj6RIhmay6HtJWNAL0WN66vmAmvcZwxy
3K/V6dwv9dphXynSfQpkkc8qtkPRPkeb9qzPSEXVatUkxZaK0/A4Ra3ZdP7iEFv2
mtUyY/osBTKquFAluW3fPQolArraNvpjTJ2p2ZS8+6GfxtKfh/13hcntxX7OZCML
T4+T5gR5q6pdC9aFh8uLWDUfNDgJ9KhpI0udgF2/3oZyYk68jFIqfvmsoq/74IHO
7hBnuRKTWOwc5Phqba05jnx8yeSX1odU1CogXRY9KFmRVYen0A8XPGv/XHXkqM+M
ceBDJ/hKAYtMkXSjdAWow49mjtnTGFTBJTuVYcG04TauNP2xyhM05mR3GMXe2c/T
XllU8UEb1pn+0BoIVCbCCZcUwdn9umyaNuu7URmg9m8ARYcJ/uNiQBrZWOjjXV6v
GlIQLHVAxBpzf3ja1/SYfVkMvvmf98aG3bSDFwR8eWnI5HK7QWFDaFI7E1ysjXwU
xd6oZxSVWIAWzkfepO+J3VIoGPMiD+5ZO1XgGgmNZXrzsgEQw28d15EnyNiImjWh
dWSvhB/EcIN48Oak3H46g7DPZ9DPVHDbGAs25ECHBTzgii9G5vlUuhQqM/fohSqB
Pu2+oWYW1txtagC+qaWhEhGYwTJY8/YHgSJ6ecj/30FcxhZu8W0Wqk2x65Kn7sSA
Eaoe3+UqdFqHxj7WuAVgTM91o+yNkaYVyCe9l9GKPyA9PorLzsPedM6PkvV/LPlv
+YpO5FHRT4d5l8R5n5Pi4ynMELQNaV47Hz9WXLrWcnbW7bfcCts0TnPT9zaYYV6V
kRGacMn0uhDkBG9J+tMfe2ANWL/4xQzVphM7YtT4JhCToH1sDAasuRtP/eMk9xcC
O594WlAf07hPRN1hiITbVR2qgT3aW1+/5CcwEuynMcUkMmnnQ0Wrb1MygXN11akP
pI3iiGOyHfcRkDo9+Y9gEktM7anuwkoc3KZrgQPQltn356ZH4tIMGcADbZsjy0zB
TbuHOGI+udgNx2iPVU5bmZ80SMu3BEXhTuXczhwPjtN33t3rN2mUu5NpmKjDwLJ4
9Q3wzbv1uSVOhwK5Atn2sxKALalCfsq7OwIeEeztuYGX183UwbqDQFfi09JPBErq
ucI4gnkiRY2dGAsTUvhtqK9MtpLBQpqQsmNbIf/t170f32g0/rA2HOXaQKo4kYEE
7AFBlinV+XoVeqHjFAibEsfxIgSPYh7u4HMob2vKB3EycRHrYSZXAvWuuB6HSwJ+
8cTYGNr6KN4KgGAatrFTAUVw7GIV7+754tTTWBtQwdPLNhXTpfDo67xmapkQPJmr
ibvAMql+u+4hT5T2rxHo4tyxkAUyF8gdmrfVpMdMlro8YP9wa+MSl/EjnFtmw0D8
GP0pdCcOC97ovLbkzwTuQzRxsVuSbFLAANd1MqxvwIPSQ6c4FvUNaIJb3MI6woF9
z1cztEmeu0fcu3rpiocNdWD13pfaWL/x1cddTCSfNMLA4x1vReJdq/cUrzYb9ELi
X4PkuZrsxwvww5ohLiI6TfLRoIyJSfGaUGoNHH/lAJWT6P+G3igTm7CHPxn3dwMQ
g7ENlxcU60ejR0IRHKG13PZGIty13c1mSL2bO6wjDST/ykwE1zn1PW2t8HF4p3y1
tZ+kGorVnnf8f9mFruFRPAxuybkoMwbdbvh5SZpmom5OE36K1eL+Sr+v26a25v1u
c+d0vfclylX0d+E397Jm8E106rtAo3xdvwXnww2EJSqR+YTanSLnyvIQUMq8SXuW
Jzdl2rKcvTpJjEV7mbrYUngmNXVx4Sfl+PCbM8T/NBk7V9KP0iHzFAhvV4Z9Zj+Y
0mbCxkjrPAYzL9Lw+FNCdIyqOhZDqpLn+b3Q00BblV3XmUVBPCGTQ7t20Y+H2Ypu
cgrYD61Ez4SEU335FSH4zcoyu0B8TmtogmNvgh0zuMRA5/qpN3nelhgj5lSwscjJ
DA5AgA2eCIJWM5tabZuq5JtImge49yeCUVIKgTNc4YSYntOjE5/M4TzMKXqM3A0T
FFQQR/5qp4E3AKliNXN7AImTeKXssANtb76OcAn/E4VjihFMJzJkKyQ8cpI1BRJp
EZMHFMUEzWJUaVTnFm5IEeFb62t6X2nYNsPZ/8OTxS19A+rRohNPGdqx2kJrWrcG
k6HkxkNVFKEN1YanVK/lOI6YesG5g0S6JdzwXKrLpl1Uz0YGHh/kTlnDTsS5g4iR
dR/SSxrY/qX6sIY6CYsyzhez4YRSoh3RuNEY7x87Tmex6fno1RXS+v9GduNlGkpz
7IPK0PEGGjIlmkVAth3vA3HFEDk7ggFEDs0LTCQPCnwT8VOOk/8c3AWOrTGEFVZL
W57bX1NlUamV70IS8WCS67vJqWM0sxYiN/UOeKpA5QqDXdF4EHSS+ijSDKZASxVS
hv77deO2GB1MkFooztpj5EGMUcyILKRGzK1Vuc7a8gaX01iGlmzks/al372Csru7
xOjF166yyrty2YrbKPQP37uUbUTa+gUt/ww1cMzmXFoh7sMwtn6ArZ4Vu7Y9O7zw
r+rugaArSMJwDOuKZ4AYTSKGWOX/ZGojYcXDDTvywkc01pbhF6shIR1GiLDsz1hm
o4HirHnY3I3amFtM0wnpW0x2RcxQ1JCTAIyLWQJAXQCElpbhqSiBGErOUyddfa7e
/UWNDOHwpbfce7YsYwAZ/50QpvBj5L5KxaAEdi98prGyb1GIlMzPz4w80YqOwQRz
HqPLiVIII4rhUNBJYkZE6AdeuGpXkdweivs1RdEvoJqsnozW6d4Z5TsDQkuZQAk1
4X5LiKZfyd5SNwxIdikHOTcnonILzd0wSxqnSBlFpO56tMp9AGT94b/5YQ/IEJ7M
Pwb14XRju78EnikfP2Za0y4mVatu5p7Z7BdMq1Rsak2vZzf0hIJB++QSXserE147
6S9v8FlWqqsTn15J9Ab5t9Rq79sxpdiCkvDbaNFZvzKUloMh1ay5Tz7GeJHHorlv
7iNhGqqknQN6rlb3BWEsHWY1tKWHYFj+9aTly/OhdJc=
`protect END_PROTECTED
