`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IPU2XTwlQc9oruoZl2oBuLf1b1bLKnXv2TcBjwruldAneEkaO6xt0gwPtHiUAX0o
UH14T3ont2eZjkMHeLDcKQnozIBtdbPEajeIKetjIX4ZPa4adGkQmhTVxplE3luO
sizZiUR8MIKs3DApbO7mkt070fsMLon/W0QxdE7T216dsGKM85kSm989KYgfNJDH
r99eEkE2LvsuYA49ec+wTR5ZLUO//m2fCNGTUoQK/musp5b3Beq3rfBIQpJ82YZg
LQXFOUAmLXViuuFdVCgvdJHF88VvxkVGWmUZF4CDpmnVDOIpNhtLAIZckQSzX/m1
RRlnXzz+D2AKmFud6KA3xzKCTSMGhIHBhUfrkFPXTHku3/Fto1ydcMnSInqTyGQu
9oQ2RVj276scsjnOd3o7454DENsDz2bsggv5xWG4nHfqNRSs3ia3fgDb1la5oxcV
0sikEGpNXgdMb1EVbCBL/+XSCKxcAVRoKBKKNGphxNr4LoQOAQPycAzSexHfTpBK
AwjOir6//G9yMghYR9vdWW8/gOcabf+iHU9+qNFeGLGvhaKrcZyTyDh5MnOgQvDP
xXbc0+v6zpAsKQdRLhrw98X+7IReGPAJG8SOd/lwBizAv9eWBA4BBz4VxoRDJkNm
/cTM5shfytk25ZTh1P48KTAU0iVAmjx+aCr8n7zhSkE50QdWv3CwBeKIEztm+CXf
tONfDOPH/P7qjZk8rc/fCuICKYXwl+BEhj5sYYgoNVMsM1SxCfDuqwb/JtgePDRX
p7QRE9I5nfDx86jeSZAJdjRq2k1SQhq0UVTBCmJBWvxiubuLdyly43z1nZdxfpfB
`protect END_PROTECTED
