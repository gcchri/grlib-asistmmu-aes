`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7k7xS5CXESRPaYdwe/8O0ALo3KWaSWTsc5p6LYxWJTWK5l1rvPP3b0hPutT96LnB
UyGtFuxxN/Xkqz9MxxQXg0yovOePWE1PpuwAasfJtH8MZBCyrgMdGffnF37DCIzu
yq48vbsu2EjBvPAPesw7e0x3JfiAVGwm9xTyfiPIL1dui1mxiJB70Qme9XH2tizD
l20OsxfboK2f+0xoaF/sD+c67mq++J8UYHmgyo/jTSz/vjCyARMzt8L6d7Sne0Np
D+bmign6SduPu5jGGPfyayciUXUXecxAjsH4cFWUBBNv218ePu2phZsJTful8K4z
9soBB9tgtuYFT9uIjdOBYejr/RMy3cB8ayYewtX6ppryb5F7mtTCWweqjdmxmUBZ
FlJ19dhmDm19EXCzlS+w8mpY8JFToWKGYwPBOTZtiUnzvTZLeY1C9UMqPhpI41QR
jmTjllenB2PLjwy4JepD1eyigKYo31hl5N9EQ4WfJWo+6HY06YWm7KRXHr6hyhfc
wLk94NSJGUFPgowhNkeoPn1hNSXdCyqPxjn6GvB1qz/6lWyHBJQIOdxt+HRreeE9
0AnhOOQFMdLfcxoI1WsU1qVb/Jndd4W00GaX8VMjVP3IkvBz5zJh72O7rQyNVFiG
Lzmm7/6aazXYofv7+pyBSLOSWSoSiCbivz0ZmEw/dnGDkcw5igSSkKDVHikpGDRj
0FDuFPy7J489fihSr/opIzAW0c0yTbTH8cidw+9JeSBqUdk9nco7KNeZ7kpup1jq
VXV2GtOyUS96cKsFVNB1z6rv5UFC1iYpbvXwO8nitfMpy4Mj2oSL3SU5pnQT7nau
zZF4TGwyGSfoaFbmd5oOerPGJ04wrsWCkfKK8cXta7pNlF/8UHYtPvcVGBM6qvtG
GOUfaiP78O1M2hib207KpNsQGHcviblWT3LwhcnPjndOCTlkO/rJ4TKVl+QMo+Gf
ElRP1FWS2IfIBo8RaTLEOydgAMpab0F79NtoGvgiAJ1WT9pwLGKTWKlGJwkHYUwb
/nKRJeMA/c7GWuITBhvMHbvRO9YAaJZ3btmLb1JWXk6n4kdKEmeQdh6nhUMhwjIU
BDNx9HCBGarb2LIN3YBP97zatlwVzrBQfl9GK1HLA6iu0NVbiog8VpnASyB+AWiP
WiCyLT5fze1SLYWw3sE3EEYg2sHEnQdyzDIX9e34XTSwsCdjkjg8EjJtGPfyH6YJ
WRH5A+E501DI3zXpW6L+Siv3bQuz+/FlhpuAQ/UM+HvFoV9MB/RD42w7EXlpouMI
0kIZpnnRbN0aGUwGwvhOcF7T4CV52M1HUWpl8jVrrjMOWF6NW2d+vPS2Tr0/E0nq
Hj4u7Bz1a9bs+OCvTpPHEqdChisGJpey4qJEhrjvAq3yADRKiIXbhf5GM6DFjjg0
w6lnOnnwdf+mmfQeXi3fY0/Y+YpUYz/v3ljYAlH2F7zZQgIWxy6oeBesmFgMRl49
nl5hdk1MNbhMJk54gAUeiKzPpnLvh864sj7mm6Dt3srNt0LqMKpZhACSwr97oa+w
FgcrKQ+sV59QrCauDfwsYDh7T/U5Zlc1c7EOQpYGj3b4ZIUJ6CoOkzqEtjwPqhan
SMppUaMcJO4JW77VwvReVZ9cU0xOS/HAFFwSLG8EBrdHtClHSEp1XFkI3YkngjC2
795UobsaRIvr5Tq14NBaS99CRS4AHSuJeO4QY0ZDMYd5EebhLpiaejSUgMqteBgc
CA2ckITB9Z0h4p+VVQDizVo0SQshGwEfLt5ZG3YSonDu4yhiFtJUAzdXmPKpOJBX
BaifrvYzYo8KtJLc3O1Hluc2ytEB6hKFFgXJeXntocYuaPcvZrw8UZo9rtqUsJrf
r9szjAVw8Bw9265O6L4yOn5ShRPlEGp5cr4zuRrMbhXrrJWri4juCsEPPq1MBTVK
TAI0SPIY4zI+Hd+xLwIMQo73GFZ2w4ohCvF3OMpFXQemIQXSoEmXcOEqF3wUpAR2
B4YQ2v+ZTMRCTZo0BuHnn3E0lmTyz0PlLiJUDEP7rwF71kUHqvn0wjFX0kyb9BC0
n6jXJCepP21pMFlWbKlq2QXbRmI6pycLFjrjL8D1PZvbdahtjam2ZB+XshbhjAEQ
RLLbdhFzacWM6825a4lVXFC75NjUD62TBAPn8hbWKGoy9rNCtxIn94Sw9MB93Vt+
Ii9D6tttscVyTDp4rK+NxTumqWT8O23dyo1Z5fyoDXajBXp9Qin0kDYseZxRvith
ABhpbeyUYZGando2w2yqlHSEKqKJNFfSb8MpR43m9CiUtrhX43gNNqo922ockDwl
vTu8/5YMT9Vb1ONZGMTrNTiWgC6CO2d1eZaB6dHX1y5j10hQ9vmnIg9BpKqe7HGP
dUHdMdMi8AZqNYM9Lw9f0hWIQP7vJhrpKQiOjCKgx7SJdysGoQvZocokKroXVwxx
51fH+mrCDolklTkpUT9/0M1itp9V6GPyadDJAYHshjDMYijBLSiZLr7zJ8+PdrT1
yOKze3NjjV2HdvQ1rYO5iqK8oTCN0U5MDXns7zuc7UznpP0+EtQeJomFvGJsWOFx
MKpwLLd5ej+ARXRp5l9Lp0V833txsb7UkWBWwXqgkpC/PTC9vngUEArEVPsZ3Pqh
RlTTxzoba4HAHouMwzPFW7TofL817+D2lDAjIBO5kqrO9PWNMXiRauDEgv9Te5A+
q9xeo/wBJnGYX1aJF4SIx9DO8kgzaaRYDnkAvxLD0ei+OEvW3Ef5PzjvnV617HMx
ldrOVC4AiDjaJ5LWjgbB5sywGJLX8SBjkHvaqUbzV7LdZ2ZtzY8Z0mIczxTp6LvA
6onLfImKtjib0rYkXwePjLxw70BOxsfdsfJd0UHyUU1nNvo9th/ARw51oAWMpjPj
AZ246G61iISGJLceyvYV2n5nI/3YwWuPx0d7p+pSYbVRGAzI8ikwcMt0faLJQoRa
vM2XMLMeQpeNpGhexlHGY2Z5uPTB2WDU2rg6At8EE3sOSHZj1U36g41WZy2CTAt7
aG7IEYeDD4Hb87YnnMKBpfcTxl2ubg37IWlynuQSVZhGxq2ixzPXBYc+rERoZqDc
1jIgJsu+bjkQMQXmKUHicrwDcMViP79kiM7q6mU7fFQASWfICZ4uZJROfwPmhj50
rR8KJjmYWOSoG3Wcxt8rEUY7dm9B2h9CYZ5af1EfJiQNVXK+Cm2fxpFrKWq1RBfu
UqloeJ+w3TfJAk2uOm+E8HdmgGuljJI7qSlMLWvqfeuh92GA1fSX3L6MqD68j2oz
R3mEGPf4/sY/liOB6vswugkgYPkEq1F70scB8h/sUx9eqLJVJQJmaXV9EXPXfTAP
uzhyjbSH283XaiDWjYbwH4H6wq4ErWdzuI4tmbfz5ta6fbhrh+K0P1Ao3+tMTmul
D3aezRT0nSJPjaiSm595gP+KxVuuqYTDViF/EfOcXKOVgvLA4X03F2LwKL25O4Rr
EFavky6i/NWt3RN55Hl7DsLZGrmxCQodQ8sRR4UroY7EkjVJVrxnrHR5UU3K1iJ5
bsF9pJV1L2SGqXTuYykt5abVaS40V2vKdCMY73jf10WjObBLsPvjPcRkMz5gdewR
b2buM00xLRJ9IU3Glh5RUl7nmvdY39+t30y1XHNAqa6z2p3ckWO0WRmmUvjf+Md8
JviMne31rhF80CE2Y6G7Ncc+VQLHlNsIAf5TscSvAGrpGaaizIE479YPxJeSOozG
skKZYmGFTKk2CkQfz12vlkZGBf0eR/Bv7EvzSUP+GmNVUSlnz34MN1yGLwDmPgk2
p/yeNq2dbKO21z2ixMtdAUuTL5vt/pZzToKvEnOBNo62f3k69UT1SMCi7wnqiYHl
cgGp1BC9pDqIdKUmgw47+xomMNwcjnveP5FT4IsrapEVK+LpTe0rhwOpSi/jd1C/
0JmHxxhiI8OkzL83Yzz9ccRpiRUlh1AuPvo/5n4+rrO2QIDjxr8E3GzC1Bd4Wsmm
yC3f294hYWL36ysklqoqPa/zNGbaKQhmT0yjo/5Ffh4NaRNBfnvxRhLwJRuJTVKW
tmepqycE4vcTrIUoUQkkhmwbsKJZgPItvb7IlV8FZt41L8z+1sOzX5aWA7QYtgdY
MV4Mdx+xAhEWR9RhvLT/V+jxBFeFaUOpK0s+mgeANOZyGj5kisKVh50PSxssIncG
F3T2NqM8AzU6jeYy+L/J8py6a215xZyy9kJyZE/c+nKfse/RWr9TXfFgL2gHMiv4
ZFttbzwvYTUYwNB3IHhHjd9ZzhDXfepXNnmf4Wjri4HaDhDDPA7kPEMtRkw+nNRE
3MPyk/jXZ4xvxCAVwbY9bxG10fxMW9vuZNUpYzEZOOl4EkIQOpbBtMf2hcVAhSpC
5F+PfnAvTVvR0hKpX+RQbL+8T6LRtDwUYMMBzcGKgYH8sj0qjCftbxGkXRM6SWIP
`protect END_PROTECTED
