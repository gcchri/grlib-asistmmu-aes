`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iq+7zX4MWC/hid6shJu3tlkIaV2vJQzRvWTQBOV2WXaoTC8N+QzY84Ln+W5er6Ar
hTgDtr4iRTScV7nsSJu8vdtizksBsvvaBHGNsqDsc+9VgXckZ4aWlULCw3C4Bo8r
hKqPkiGYNfDykEjRhU801xuUeEhdWWECFo4UH7rA9jhnkSjnvJBkNpiF+rMEGFlA
DouuJ6zdwv8FeE1sRmUchYxIdTHl54b0uJskFBL6LAyictObDRo7v+m3502xwZTj
6BcQf85OYZHtsiju6NAQdfPK4OlMIDSQrjQcT03g/xSQT6vh3PV0JkbIdwXoPL8f
Tc+704WFQUbPFbl6W2/7mX40oYUJcB91KYH7kjt8iYFX03yURt8yHz8gV1i7VpxS
yUq8E+7ubwmprZ9QAvYGOTSQbpGl2BwzsN8zJ18uAMKRzZ3NncOvLL15n7XredLI
LHV+Cec1+5Vio5BO9gPZsHpojZhzZBObO090h3SVwZf5TtVy2zVo9Vjx13aoVt+B
verJr4abNZJ1BdF1lZhxLqMrqKbtANX4LL6FOq1OykhBzoHXLavDzrm8Ha5sPyD6
d8TWETWDZdHXo8+f+7zWUxg7KRHQ5itg5VD4UZSU1oylu2teoOfh2UUY9LQUI4B+
nOmxaQMbbnMBxbrdkdIMcIemFEJLMlZZQhL8+x4R85gWL2E18eXe4Xcda5fdcBvO
8aAF8hGjUPAf2uBUDLTg651mvexfeetNZiovhM+d3QenWrTjSXKEgyytgsEEYayC
RfKAt9q9MyBx8v8uFeE0UUhympyotYtwN2DOgLP39ZqKpuL0Z8mslTAdWCrl2nmR
ZFVt1TOIv0Qfb3Lz94VfzwzhJnM1QiaRYr4F2Q5S2Q9MXLMWhzHqwQAgLwotY66L
1YxTJlkv4VrafgTEuqPIlm8K7IipWbvK+SwK/yQDf7Z+sLHyOYOVkvgJDA0FAL52
6qc7rxL/B188gawRkNa+3+ddMslEGq0yZQvhQSMSkzzhhzDW4SpGR3z6NgxbKCOu
V989m6bIcjrw3gHRKHZ9/2FW9xkDD2L5FAoLU0gOPssf9syM0uID94WcF4rIPo0p
EMGQSYLsmc9m02rFwuE21PBvFjlTo1rM5PKGUWIbdDHh+T1Gbjx8PeDszGvj5+36
3d7400F+fiazr1hue3/MpG7mnDQk5UOmzaVtDV3e+5y0fZmAkkQE3V7gvK7Jjwde
`protect END_PROTECTED
