`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dqa7ScP2Wqsy0wFxsUsLJf828Hafl/WpFN/a4REW3gkrClKJ0FZa2Mi+y14kYC41
gLJihKOWpE7ZXQ4fWVbKTO+oorFAK0UAyTVeQJ/jPLEPW1Z3YKc/AX6OLppeHkJk
qDfv37rqTJcPIwxWDy31GV6SEUEzOuINzfEqrlfB7jFo8I6J2rRgXzG5hBGDZiw4
KdurWecig1LjkpJh8n3r7n0vGz+lRy4LNRu+4fdJrKDv3ZZlHKp0Pd7kQIqtxxHV
fBqWI52lkJmXJM306gpLVIFSQmoXMKNNnB91hd8J3Gsh4SaH+zFpuKkBLS84gsmj
9mVt9tKatI1xpBE7MwlkIvwB2E07Rkcyi5fd2pFX8ebc0F5pe6EqQndZ1Vlg09DJ
lm880ObYEZHeX4GZ/zi4fT2SYXAn9tYsAOCXR+XYrERmAWbxwMncBrOsT0+CNe8E
Y93pSaC2SvLw5ovR33fUG5nAq6ZdPsuo8Jza188n/B8a3D+3+KYAidTW3VRkbJuo
8Mzzu4DGLWqLflyIQMyoLWeZYLgn86pC8nFfrWWvHvQwJaeYO5og+iMjdGspRdsy
ryzz44esiACBSa/8ipO/VbIvQR3lOwGrqsjsyVi1v/WKXK3PSzJr4/uNxL0gxHIH
6RNOcudn7oooz3l8fYbRjycnGnV4EgqJCdxsZTezjVvH9hdAq7uN0Jd25fn8fiF+
2G6xMEqR6fNdyE+4Uk+IiSsJBpZOGk7XUjVU4LFi8nSZhoTGtYrSqLjcPA4rwIB5
CsOs3YGyKEV/z5u8n9d37/22emgQbhnhFwB1RMhYWMa5vbM4oL0VUL/Vmmr6sHlW
EwQEKSuZ0w9UbSHqjxJsCWcBjxGGo9aloY45TPo5opmsX7spIcihc7iN0SW1hIjZ
JA2Lur6U5i7GeIRBlizkhDtswDW/mdOeDv5XgOtwCcgxOteYGanoPxBLqPmFeHRV
DHG2x+V+4wGUqo3dzu6BldwhlIsYw8R8GLrkLjEu6wTQQK1gz8zMsFo2pYdaefOe
b+o7qtOqYeOHEi4HpJuR1KpRjEwsdJPfVyxTLH0gzwMCVDQi69Ihmlt3GMcI9B8g
k1KfqGsv1OsGqush0lNe6EpEcp/5A+QRRYglfk+GgjxUEnHmxaDykJDNtN6vkL9t
Yfo2mtEqhS0bD6oZQLxa2zsHYzyxtgH+Gqc1ZfD3jVTVW6m2EBdSiv/70C+1E+Zn
vstYQz8IFxLt8BWJ9dMAYw0GLH+UGYMjNaRfzbnGyzNuXLI6cGEq+Tm/3opLoYnv
fs0FzAWYXnM/3IiPEyICqLID9Scr4IHh2BpNWLaEFSSQ9xIumecgEqzsEeHfoKOl
Wq19A8T2pTELyHmJPIKW3JXwjTlDg02GbRsNoh3xdl7MbZnQZ2naYFN/tjhV2CzB
FUgluX4/Q/cLAkYWLDZdk4Ucd+7gpAPNjuRBfr5kgILID4OfRZXzgK3f4Kc/ChYM
uUNhGLXQcb58QwgUvYUHcXymbZLjVY2MOMn8G4IiUFCznvNmL4Z7f8A0sAe5TNzT
sIbxEIMmQT7H5PIhC1TFUwG+6tH/WHZRz6XP3psfd5wqwtOp8frHpOMgPW3DZUkU
wJhQwu66aiuw3dLQLNy5aQhn+aTrREEacPZ+IwyNVrdRuxSJ/7TjFqR7/LKd3hPy
6+5/IIpGgvtjnj+FerRYqPdEQHd/Jd/zvGOlomzoieiw4VUWDH7b67k/ZMo3jGi5
iDOkFIzjmtoHfB6rwtta7s9N8VxxP7EzLy+wEkwVvjA=
`protect END_PROTECTED
