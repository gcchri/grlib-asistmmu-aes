`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ArILaUFhsQOQFsgbtRKPaVHjU2kdgA7ad5BGJKkdikssbJQoIyLnb20Uk0gyt1E
o3W+0vrg+72/bOADYlh6C4m8Q1jg78SbZd3PAEv2kUI2H3ktweZWf9/0BSFiCcYU
z78h6XBefdq/lIX6yEuhrLjHqiDHoAvkaZtfCd0A6tlcEneg5aA3UkfHz8d1XspN
Vnu2dxWyWMmOVeQDV8BfDHR5SktxwD6HeEBKkHEmbknNRT+ZTjo3pXfZRGg9g/r9
ZTPBwTWAnW9gjVVvqc6UN+2cUzhl+LHexlhr23U/lFayQXppjTwtx+vpYuDXSEaT
tJxKAuy8DelZaEOlHr2y3n0Mm1+9sXvTcIkhD3MZ/it787DD7Adesz6AgU/Q3Huy
mFE3ODNjK+1IBsnAwKgor/OJcU59oOs8rBjiEcJHgH/PyACAzglU22dS668IaiVn
fXL6qTjc5CbeI58NYyy3Nvn26WWx12paiQEux2fmUuKyZ8TcuyD2C6XAUwXPdQ/a
`protect END_PROTECTED
