`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2hwNbMvV0A/O4ID2OdJ4wQMUorSMPc9lNWCK0z8GefqzDJZXcUtkq/KboLFEw43b
cjgD3BNuoF86tGEdxQtLT3EUZZuBjh1GDpgiOQcVStN98wICf74aK448NO7jrvs7
Ze4iQohghPNOxwGPl2ZrD5plTzdLR76LL8LiwMBkw4vIMiGZcvSkhUkA5zpqlyjg
NYIJC4d07BZyogRq7a6Yx71oyGHD47IvbAWW5a5pURLr3BPq2WYJkFzxo9mXRf7Z
5jzJL7+p9O3lLnkWF6fJQZ45enRX1wMJXjTuCrtqz4XvzoG45JH7nPzGljQ5Gz5i
cV9YvIIm8ljDjVKxmVzdaINeJlprWPn+uAOKGq5bZUCkB3tM1s6P1lCXkC+30kX4
tdqrEpNZ/qk2BntaKG1Pw9fKxNPvmTqbo8NKaA2tq0E+9TNLrjglElbKENiRnhkb
`protect END_PROTECTED
