`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V1njwIMOk5iG8x6/Q7dqNXp5RXSpbkvegzZAu9Kkm1mhnn1KQCnpU5Kh5u0klVvk
A2u778LOr41A9e0UcMuHdDkSQc5Y1BNh6LysA4RJOk6BOAaaSIVQOwjHaUeRzlBW
zmLQUsh9f1oH/JqHy/VkF/esW81rdTHiiM7zIfUPG5NQIZrsfT4wWRAWWWu/dtn2
MSOIlt+Ydo5mGZrbOOMyQBImxN7iYUv+ujYYgvWD+vPuIODEAbazciDMs8tIEb8R
arLpJKDFE9a12JCwO6jsBJInqyTkMoTwWnbHEcrarvgH4KKElURaEv6VoCnUiMxe
09FMmURJK++MyvxrYnospg==
`protect END_PROTECTED
