`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0EgviOOZY80vJw4yWezdXFryz4I+OcHOUybyOT2yy7uwWx1krq7kCOHJv8I4NxIp
EqMFmS9uV3GdXIG113WNDQIbgHFTOwKfutuzK0hazN4b/ZVnGDa6bkq/GmaXxzAH
6e0NQ/KRK5VFnAbp/6CIC1zHTA+0MxkDkorM3GOr6ugdvp7rJaPeWEfBCENhT6wS
IgKISI0UPiSZV3jqDgObq78rliNNmVp3LUbipYUYwxVRZbB4FR/nZRyKcSKIQ1pm
sWI3qRhxVr64Z9pErxUZ/hO/QnkgbpYYnYzrZVOkxjo4e2fFjlINTScKuxs+z5N+
p6B++ke0sHyLwuEaRqlNkQexAw7j9pYFx1acZo59keZdVB713n7xSxlw8YE8lPRc
EL2QwtemXllS7CcAtzxf8SQ4nV7eMsifHy4vu90JyHN7x/6vy+VX3iLU18D2tdC3
bB9iQOQTxiL6/8AjTB0f57wbWEUOwk6IP3Yr7gM9CMOB+AFjMLa8gmwulIc6cThw
s3WnYdJScRRNv93RurZ4VFplPMKC5qW7GLwxmGP6Fok89ae3ey300eYHOA4VUAL1
QsWIZr55cKTdqeBDdkiUlAHNtq7m4ji35jfC6rY73wfnFH//pze8gloRu6yv6EPe
A2qqvJh64zaUmQkQHm2236uIH8tsRTLkzL/9MRvwCCPwcyZMv5nbtmwRlkfobCLR
JysnEaZX8h8oJpgmARX8xQ==
`protect END_PROTECTED
