`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ftZFxiXbB+uX7DW+g6m1ZaTqQnDbt80Y3Gr8+UM0zy9KnGa8PrSvMJ12Bo4+8Fh/
lyhF7x2qaaPjhHilPufUA8rqRR/R8kxl16ahhEm0Y5BsFhslOHeNjQUhZVWnNoC/
bN4kZn+G8bPzawx6wBm7Xm6xe8k1hANXzhUabaeyKXIugEEUpCw84jWEzziCDvtQ
SR9A9fBydmCfNP/FXogFByC1WKJB2nqMaW3Fn3KXGLullB26VL9xyOLqSmKUoq/c
wVW3lFfg+4a2JluAuz+tNTlmA3BJ6weLEP4y2C3+jLGxn+x9u7IEoRrGVMEA4r3H
sqIWi4eP6R/ElFRBkliXYQ==
`protect END_PROTECTED
