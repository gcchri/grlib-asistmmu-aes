`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+x1o0OLywZHdyNVLgFNesb+D71h6nKQCnEwPoAFk9Ook1ytMZRz6nasTymCi37ha
s/uFJprlNo++zU4S9BvR/gJg/zt606Eq85dm+IbI4+mUlqeEdh7UicGHFNKGLR+v
z59a9wKTSDiJeF506Z/A2yd7/9qaUh4IFWeNpMDgAu528hJQyezoqMzgJV6S42KC
Qns0InDLR4n0NekzWHJ/Ojhe6/CqZVQVQPTn+VwCe4dYus4pb3FpsP04ycc2UNkE
/coJlGEb2esMoMoPM7grDPRUMUg+83vGN6EXotSculaJavtRCa2ry2YUwQo2z45V
Pg04VG9AqemhoNKDuT3QBpTPN7Zkv6k1sCWst2xAYKVyLQpjdHkv6hNpEOL3UjR0
5kKcYcMwcOFUSixJ2BdNzRM1ZLh5YmEt0k1zQdTv8mwnBYN1fdP2g0Gfmbo/rsTv
hqaziRJtTWQ79ONfJPWqXMSbV1CyaaqH4baQAZlEdYo=
`protect END_PROTECTED
