`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ljGSq0ziGi+6yeh02hTxMoOmwaeW0fxaug+xYpSUFFmLQMQzLQvcI4RitChHNLad
EqmsvQcw10XXyKEB3LjMHDDgbqYIHHhKxeLPkOvWIAqbkUAuVlyhyuJX/I8k8v+C
JyO5XRCsX02Spm/RuETjzgB1yhshFoS2YXu2HPu9NHhtNL/Y+g8iII3XaNXmbR7W
j2BAvfDjSib/mnUWd82FzP8XrS4xPd6UYglKtXWe3kKQ0xfq0/0DL7ZVBu6qeO8t
Ee0v2rwMvUG6JqKAD2qBcQ==
`protect END_PROTECTED
