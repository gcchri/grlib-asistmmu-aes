`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0ov89r+t6A7kvdZOm8ckpBzE+bmjuBpmI0NZvL2+OUYXQ/N+t+Oac5xv0kEY4yVb
bldfADgsaoRS+0uvOFOIyXAFvAGkvgVayw11LSARTyQztMRt9h5WtDJCEXLkm/Fa
RNWK8LMi4y2DWDLvfqKR04Rr7F5DfSB/bNQiNPmEi2mGc8KAYT688vqDMGgK46hz
Lz9m5AOErWLEY85+WyaRAe6673QMfj3m8q7qmPZ+RZtRJ1B3i4YyJfGgfnkkzHEo
U4Vgtdf2muh67Hh9sb+kROT054erS0wB5oOFGvpK01cBJKWiOo+T0a1xygHlczcQ
xVQQ2cVm2IOklMMINfUNma4usMLBPfRKR4lVptBvxUKa57Mab5N2Q/X22U2H3Xkc
wAcJ+5qd3opjh5v+qAZde1SoIHZ7IeDu34o2Wh9KJizirpAwdpboZqJfv0GuqBOL
jSbvNeNf2Rk8vz4b7kwgNyNqKe7mou9iiBxX4t0B4yJkVLkL/Vu+9eLHU9fyL+se
VTOLLb6PJzMqZwBakribu6rj4pqxHU+JSsdiFs5r5/bF8i2gqcJrO359kv8sbk2P
LEe1iNb9UlJuci14IKa/P9Eu2yBGDdv51nY85V3pBp9JrERZCApkdKD5Qzj02Tjk
qH8l7w7ahD8MbhQaQauH7tiLnLqSnv3HDXoVfmQvumY959p6o63PpQawQKiBP8s9
2GwLr4BAJNU+coxi+UAJ1J4k8hosRZARL7K2fz0O2+n9LRoqWW4TtqDofnXQ70QE
6g05JfLJpjG29QNd+G9kDnLVkvqadAGjFYoDdVkmF5LyiUvUDH8gkx9E8S/9okDY
1Hjrl0KJ4lb3/FPAOKZ/yjls9Zqvi6GG4S6KS8pf4Vz37jtPKUWXetwJbSZIEb0L
TxFczIuUrkDZx0wazVUyzA==
`protect END_PROTECTED
