`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C/9Br9a0NjpmG/iyjWZh9d/630luRRTpS7nsLFBIlD4+y3pZVxswfYzD5ao3JRog
/YuSBGIrIH/23u8MPrNSl0XHRrNwe8WH3dYkvJn+I/9c5mpuVoXSpzEabP5kmiWg
4n2w0H9HVdsfIshcmi9FrGITTph9hvVYafbLBSr0SJweKdoDMMNv92oFo/OVdZ0E
wQh828vkiWfbngePlk1eoJp0qjtPx2InWQaaB3QQvaRDx5RyylYn3N0uqXfueqW0
wfutMWpQIAIdUNHEl8EwT9YsH+pnAuc8b7TetvPm0lzO4OCJTPAah/nR577QnhyF
C+JWD+awY6i3bOhc2Ravu2WjXwVUMXph8m6eplp7vEKCFPj2b56PfDETO8pCmJZC
MQrCPVcJJNSbUoZcs9mCWkn7OuOFFdK4g3W3GGWOw/bpN2SrkKMVMYgHsJS0LaHg
kg4cGzenQF1otTlCFKemuOb3zaGW+JzQbgSkfB74wcb+mVbBoMxNrX8aPlOWthcK
ZnIlrJyF/JAl8JPFz++zulfhfPiizPT7CZ6hjrhZp0H3ZyyF2DhYsuGQ+YLJ9sbZ
g9JNXzP07bPqpDn90Qh3wOjj2iCjq61FxJhtFq0tcUEVIlIgBgyL1o5G7/RfvSlK
zcSXFARkEqaft34radMy5xT1Jk3RhJKS5MsvO9RqKbE=
`protect END_PROTECTED
