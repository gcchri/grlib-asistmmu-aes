`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GWR2fFq5y/VqWEWrCVlvEe1cyzM901atxLWmogJh9hF8QUQ4B/wSl4jPRp5RAM/P
lpuFCthT11v8UQEstRJOJsV8Js1SqpCz5rHArvH14dRL99QfiXhgyrxTr3hXplsp
h1tJQ8w6jqMM2fZ8de3yhkKtfng5qzvol2CdxddznLyE3VUNKj0xtwPpoIbSsmnG
BS9eXe9RvIcslUbHH3XwHYVm6R+8aci+DSsNObTgixDoNF7eGle2YI/DJAHE0Qu4
UHPiLf8WL7pw796BSsQ2mKLcqWKBobDKJwisG6dX2Fapw2WMrk3j2L9ZBjoDteBi
HnnVS/zNARx5C3/PY2yEnEUf/0s8mIKNYdySEg06CKs=
`protect END_PROTECTED
