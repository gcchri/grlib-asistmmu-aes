`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zc185JpHnxPDBr+/c1sLStE9128mWheVveqqAnrDTbgfBmuT3cNl3tO2do4WeyLP
FdhdVkIJl5mn7uHfqNTKy5yD+UoOHvszC9RJVhyiCEz187oEyPoikKnQ8syofsxi
NOqcV2ZbCNpKT3KWbAIdY/E1srJTlyegmUkMMzW6VoPGF6QkMx7M8KKFZ2SpwHI+
dWOvt3mYNPCBWv/Viz72KY5ThrdA6i3FGO7Fp9gWe5ZOeVDTZhHZHGRCtsxwTVyE
SegGFmEzfnCatQG0ZRgbbaCyG0dkhRpxqyVCJKX3RSaJSSjnFu563l5NfBVTMw93
U4uwKksslKfLoFX6/kJ1AVeo0ZsD2iKtvYJ4+CC17qEzMkFIc5+9ML+7MkH0wW5u
LfZKjL0/deKstg5xN65cAw==
`protect END_PROTECTED
