`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RO3Xy4Tfv9n0H3GF9sTXBL8c+ojzvxzxAPyD/mCsXpfD1N+omS9ayZ6jh+c3nlRv
nrbR3LTRPH0s0jWtPhzA1mkhzZxewv6efJ4mEoXxdIgb2fFZd4iBHi2dFBAiAGka
GF9xKkE779rWTt4u/6qWmOS879jqgTWqLi55wdB10SInefN2iI02SWQCpIOWV8eU
NEeDulNrXRmqBfO8RvopOHZQs4+rkwasoAgZo/gN9t32aB4xI+mR6DujZNxQ7x34
4M70u/Mkoe1DSgZY7p993v44bdoxZ+KG4fwDLkXu52N2+JNADgEZVPNGn0Ip7QRI
Ief0mo+OXlzBSTDrgc8WMtKmt52plkB7Hc5A14l5oXEyYmS6BLbY2mPJ4wec16yV
plDUcEbQg4iRXHrvzrlf1CdKmsmLDR3knmoEBvMmD4HvDcJzFEzJ8De5UvoaKKuZ
HcQuuZqtys/peyUITeF+lUcE9uIdC0nyN7D+kOsYk7QCqr/1oAc+NvXUBAUGwz3g
lohBIoLkcOM7yZNxFOrKcyrXb6OEqff0jSINGdzruUljqgSrwpwOhCy8nHdSQdeW
8ssH2mRVqT2CHUYLx1yFOSsdZOKVnrYskQU/48wdzCOsVljIRVMzBwgr/sPM5M++
Z3PBkBWnz4ZhqgOStS9z9r/9c71OCgFKajMbBKMZZO4HXkQLVCuXXmTOOmJuuVya
qBvXID/ji1dvPl0tr7jTeOQ9kPrGwvyMSDH3zJFcuLxMGu5buZPpQ/Nla6ndMqWt
f9Fq1inGKFybXZkATtJrCZUcE9aKZMFfNfOMYQnYVrtabonguyfj0HiVvBYOsZIp
3F9DzDn4bfh4PbWGiJe8XErF7Q0DRRix6SOjQx8Aq4XUSchoQI3yoxkic8zXzp3K
Af3Xg+EEduztTPVFgufvJmXr3EMKxpt4asL3Kk3ugWMX8yOtyEjbgBzn0XaMy6qS
a0KlmuHdMnleoLxZrT01PVIe1icZAqERy7Di9WKKAC4IeMydH9pkU4udeaGgZ3uP
0yjU2JRj6Cm5+OMucnV3kSsC7xXaq8SK5DI5mUbXt6q9jBBZYdwmJQ/+FRRoiVoC
Dvq5ELGwI4Vr1OLkf7fuApPp5pAeahxkfmafva+dV7lxPPVt3o1nrNyg+3JSzOib
sHzbi1ymoTg+KkDOeY3t6Uv+589DzAsL6i4ircvECBXupx42mZXt+JfcTmpQKJ6c
hBEcGQG5DP/fkNaNrjemZ+lzClofccBYs7cV39Z//qJu5hfae3VvnfKqNyuPH3r/
FWWlGYCF1EMcdU26IonXQDYeBjA2veg7eE+c1xjbqBB4vzUCjU7TMJFQ64zuv/ae
Q1RVNg6CJjRjBW6/V6HhbJLI7nnOeZ5jByEOmMSIdmxr6zNEzuODt8FxbP5J85fk
Tq3SOuxYBARFylM+uy4bRwZot7BNPlMIxtdY2l8pkhkv5S4SkyDF6IfdZCkB0Bsd
NHeLWUrtiu/iFpnb6H8SstEWfS0Ky08ri4M6deoYzQ6thR/0KJg6kRMBMBeQpKGj
3g4RJyOkjezw6lhiNyzvojcowZ4ihBjVxnlVSO1IJ0hY6S3XG8aIMiLvPnZhlIp4
MXHscYIlSJYTaS0SCwxkSqLo5SF7yMtGIFusqK3dg7BU9t3/DIzhPIV/J/xh5+DO
b4ctbhQNSRX8UufDKHU5lkJliQgmvp4MEpdWcbwblcw/xCH/bJx9QrhjRaY8IU0f
P8SU/S4RXHrrzFsleX/RNBeihyHeWEmWnT9IbnzAVKf/tRPb5nvZVXrWVkoZBDOp
OEDcqA8Rvb/QpdBe31tG3OuhNAtKgVbMnrsGlneaM4FeVBcps1FS6LNQrcRONn+Z
5CvBd2CjP61CPK2EJE8Wb22aij06oaK8W5idCfkxVxt4f9/ZSG+IGWxJjv+2Qvad
vOb/p8+mPgpwVjCPNDGePntKx8AKK6O4U4OE68hP2K/ydjzIezbsoOSfST/N0JXe
ix0YDK89b30k349Rh5eX4++obh9CR8RgPj45SZXIrdlfAHZ7oiZkpv+0Ca59kDtW
V2DElpbE9T6Ar7BjrdqUOye6/U1m1ps3de57kNItzBAW9OtAUouwBoikgTPLc7sS
G39eDmwgUB+WHv262le0AVDAstQpvTSvsydSwWCqKcShlQ1YEWGBJrTjZBQ/RzdB
105/pAfBqQx4BoMsL8y7HMT256su3F03PlQSHG0pheHtuLZqAVwmr6QYfoqxF2Rc
UVRAWdvff+4ueUbp45fI3+Pdiyk5HRTV9F9qspapEuhjvXzNrjHT+pqNHWLh6G9s
qmf84Q7KUeVELs5pwewOtP1vB3KQWUGs253qtEwUo5qe827jPz7gl6D/u7fPO7i4
X1zGERGr41JxOp0ZtKvellU8sVR7iDIMDBJ6B9H/t2sGlxbzgUI6199zuvA7MXPW
qHGEGHkKSK6rq4gADII72IVb7Upi/Zpiwi8Q80dCI1eioOclOx0PlT8S9VxQEP55
VewwhfyukuVUqlhSbt/H+lSYepIVt9BUeCbDvnwLFZ+S4cmf0JQvQiQpPKPQSkhS
sikuoMNoQMXfVM7Y531wM0lRylaKcw/7dCjBxw0Sht9+laTmkUaotNENh6wyMJD+
tlN+ZkOY3rjaL+2Q9fKJqid/X5GzeURjOfeDU8lgcV26Fv9a42p3TUkZrX96z8UC
1PL07XEyc1VrMgPrTaLvydl3pZgRaknlW/XCPU26VtrekQDeJyPiBXY1AWDFII4g
FKlDSCXwICb4kHwxM+Jtc0B/BWVxAoO+ekh5/b5WBL0i9H18I85p8UJYJcATyyQE
JHCE2YSEcHnA7Dvign1CrWZsm3LtC87979t3rwmu1QHvOEgFkQCjA77ZuMY31pxz
sINgVoVHzll1z/sEKHu7WpnFgtjeGn4TjT8I8X4+Xn+j9kRJ6daP0hgE/kLGLHX7
vNUVY5nAhQ5YRODhxy/qsSHB4OtF4KJHQilJjduUb4ABlqTrx4OEN0NGU/84l1Z4
9M5lSc2KYTV5478Gx9BlH1VCcJcgUhnhFnqIqJt2kpsAVoISWLel8W3zYS4rVrQ0
PJdtFBFT79DaYfb7Tk9qvF0mmjhxAd0H9AG1qKduFdvtJztuiVf7QepvLyPOA1oj
4nTIR5bosMqUJTkPpmVVNuPILdYuCUqDhIRRc/92bBphvLadIGTP4Y+xxZpMQAXh
iNi+Glfk3IAxew2KrGt0gLlQjV9IckBlrmLd5M7zKRb1emn7Na48N5wD0O7IbcQe
W//QzhAqf0LsE3wiYYWrLwoXyQwWmkpW1R7bRbuhqwAa3NUfFc2hZxPjmT7XCG67
BK2NrffFnX7tyMWl+OVGd5L95LAcX0yz3ZvBY1Ijfnqj7kqPFrZtLVF6dztS7Zs7
CA/8AOE4xwzMlBMSQasm15IKb4pj//vxxHTygwETWKnBrliDvVov5ekkegYpMOIc
5UWOLurHRMh5Y5fFclwMvC3oOipd6PDZ9yA9WLHeDztCJUyP5AwP6H47/zCyb+CR
yAAZgwazA+Qibel0aq2fZSKnruDpstXpuJxXprzJBm8s5zXftY7apWKitMbsuYIa
lyevhG5qRFiXCMIyc2C7ONTFd1uHkHRdZr0a/GSt402AcCROFoPsBOU91cqxGnvs
Q2uBF3tLb2wxwU++NnM/J5/cXmpNGoPDkrmOqysc5anV6KeOwbRfHPZqAzQDwHf2
bzJK+c4BMdCN4bZKLWOuucaN9SeEjpW762oven2gEMx9APiY98tNEjfnf5QJjhXC
aiU+NojXWY8sThK2Ha4FItGeV+EwvTVD1iDP2pyfQzCEbIcndfGzh7MOBvnMZ+p3
YyNq98wCDun41dxXRLYFyeOehxlEVy+3+hR24rg6llo4Ehm2UE5tbwJDMwOdcFZ1
fdCHR2Mo+rtPObUKfOmqNI+kRPVGJaYE6YLWytcKT36Fta3B0XmRy7H0Pd4qCF48
2sS8ReQk79zAmrFUIaoh1a1jyNZ5cBtoyvvYY3tvFjRyv8lkKKx41adK28ujSyHx
VwFQynjdH4zxjQUFeC8G7DialR0f9HzB6GY7GBW6ka3LvR4GQlA+gfK82DaUqgli
/kFdbFhiebxDeC2ZaIZMFs7jy5t+fkwUsy72kH69R+MLXhe8M9TW2P7bBBzMn1aD
AQHMYCOQMQL5T4hfgpbuf1w6ksHucoTIAvqo42VKlreVAuqYN/GekfBElk378eCK
/bGbo4o6WpqIM2ZQy9H+haMRbWQp5fBuxS8FN117L4z/e7pZQta12U7/f3d1Hx3D
1CxOa0SlJmCQQU/Qw3iYH+JiNgSss4LcPmfblCG2xJFaVoxZCipP0Z9s0kh6TNZE
9z9tCWfrHQN6ECzwqv2bpG0M5I9j1yRwByeIu5c7QQogQs0KQEhDNYoRIdfa4sX1
a5BOazqgmQTmMAX5ao8vda6s13yPU/sDL9AZMv/nkPhB4SMxOr9U9V/PmEA+YsCW
QIUGqrdco8KvVd1yLhJd5Q1f0l5H2B8YoYfNGQ/UpoIRHwSrOFDVGalsqrKFkx0z
9kd7ARHokJM7N+xUW31Vp7/VLEoZ6EErPrUFyidldf323jBLV5DsQR+QRf9nBcUk
ZjCB1OV4LdQwAueuUhGUwOkAe/+d1cQpBg50CjXk6jzivg/mQq7bI3dbuCFYi6h+
RxbQGqvU/l+B13mt5p9CE1pRdHeC5xjAtkKxRzR8kvuV8vXQB8b/VIuoRh06uMYZ
kXg3nIxRW5nsR2THp1H34pf3Cdt8r/qQzYjkwDFc63U02CEyGi37ZczjOsnz4ZyE
Zb2x/gCP+9HJnaApC4ps7FwYaHGbgk9Nmn6vmoZwdd3phWjbCpQRO+atojG36p7a
f9aZRtbVDhx9TAyL8FjbB/aBPT8aS6Plbz8zUCHGFqdewGYRN3Nxr7m2yLW/LVce
DC6AMNmPNQD2b49ycEFyh48O7f0jYcsP/5aJuB25U03lBfwUpS2pcMjRM6hdELhW
a0jqYmzRcDXdM1dw+Ufx+lDa1VnUmr++83RenBZMhGNt/MFn5YFAouG8h14wLCeh
m0tNy9Tsz8HlXlxyd9OzpQwLh8t+0z1nrZVB+dLuZfvk6jcnLN5ttnSTyz/Q6JYI
9keyqdXxH86LDD5B+H/L08UsQmNNaPcrEmq1/ywk4wJeoXsh0lh8AJVLuLXys4qE
rPiIMW+adY/+RT9GQ6plW0/BL7VnUpi9ljXHFfBr1buLrNWj4tuIjLpXANP16FuK
S6gdFzPLg9Acmi03WFAhTrXT/mt191265r5ij4mRggLEP0nqB9wHxgYLRBE40jTq
cte4ofROQ82GYE/gQgUsgwPai7e5mgaUJvkQeG77XVNUf72VVNmeTPTkgzTE6RYB
19tqrafA3SMRF6LCRQmwDGxucJAcESICGyvjtZ2z3OTBVFhyVgEyYCH2wMd9gWWB
AUqb5z4P9HTj1e985uBayc3cWLu4YzXZFpEXo1tB0rCZo632bAP5UEsk+BiYdkVe
9JVWwMS/egf5KK7bslsNNOSM7VGEApnj4P7hEVwVZBrz7vrfw5V1UQJEbzjJBXQf
jec8wU2t8EhuIW3rdCI/rDXN+02HWWQNxi8PYS4x/RTvLSy8kpkCcC6JdFOT7+nA
L10E4s0qoqhSjGDR8mzLN/FSzSfCKfMIcJlP0RMVD47i7kmervyK74Iwie7N2mRy
kmf3Uvw5VxFvJK/mqS3ly90IIC/rCUYNBmWJvfieW6dNGaZvBrw5d9880PPIdS6c
Tei8++cRfulkOrr4gLPmZjSrIwAEu/sHo95IgtXMKDVWhfVHZe149NkPh6CV1pmB
XqrxrstNEcAVZg37iGqcAkZKyiBD4YretcJUuYxU2inGlvAm1H3KYsX5LSfS6vNH
5C0N/Ct1EZbOOaiD5dG5gCMNLoyGovBPPM/UdgELHJVuNRA+sjA8V4vDEvMxvEu9
EaRdhJ4gDg7fJffgMHFB8++EQFjRyMmXsjer76JN06w1LjlQNFoS3oN9Vbg/eUTH
UB+6HWCncjeB7JMxjcKnzahSDKdmJec6RvCxDHnFcGnVY9Vtv2oPG3dOBh1KO/kt
+0RVM8psTKY+WiC223XPf0RSxjZlF1Ir8+rtyzBXI77OGhXDcbueiYDg+NgL9GvX
3HRdSj47dK+H8JIEnW4gtf6U9jdhlrz8yMACmAnvte9bIfdu2e6QnMzaPcLv0qvv
gNvfPWHjODfz4yjj6j2MXgWBwVIEI9Sesxsj68VvUsGUrij+QdQvpXcZS/pDH/e4
cNdhu2LDEgX0Z+5AfViDAtXZC7BB+XKHxhHsHNf4KIw6UB2CKOPL3wEJmYhaS4xU
dcYSH5REcPMP4w5G6swb5jIejmo8pHyMRfPDvV7FICEJB8uUdLrBkOBnpQPA75kj
z8C2HR4zJ2M3mmlkrjwGVej3L6bZZXg3/BBZblJKvr/SoD2cDG8gklDksoNsOuaC
hyc09DzoNLLUOU2Eh+gfFinzt9zJIGTmUteHkZwPCGA56RSNSiX0VhSDQFNqPKl3
QzyVEDyizDtOXJDC9GRUAjx/DjFFuIZbtYpuNR3ziBgmcy3PArNOHaqD4YEuwiFf
pB61Ihg3RhAdQ9Wijci57LF+QYo8zrwHE4DCe/eJ4M9pduo/VlK9hFgzI4g+I7Y+
7TUeRv2wgYrCm8bIGWEaXOSsdRIwmJjMwK6Nj/18M4N3TQYBmQUWMQxvjnnNCtPJ
R2cd3su4uQK728cmRyTkpqIfiYFyQAityGVuvrcQuR40bCVCbOl1trVyO9gfpy0y
i52rZ/9h5m/NfxhcIdpTayn7RkHj9+/w7uWBwovjTnYpXenHuZlANj/vLoMp61v9
EGDM0U3a49A1SUYBdCrkOZQNLr16NA0i2i/kD7ZbeKbMyZ9dnIBTFgbN/f5jOCz1
x6bOIeBpYMENAezSoypC7UNoJXMg4Mu2O3x5I2ZAZWX7pf642i6Afm757Z7i3fXb
n9zJ5qPXNB4/HCriQLcZY7PCl1yTEkx6NRoeUZ5IsFB78o6+wL3fw7ec8m+iuek3
FA7/trgpO88UV7VmgACMU9HwgnbG4MlLQt9Tm8ioVqU+Y06TLEnNqDo4xu8hyMGr
RlKoTDG4G9IOH0rBmvr1hsz8mHBZkmWE4EqbyO+c3M41mtVqj5m+a2ZDgkmS5Oee
X5u6AhJvqQT/M3r7VBn6/Be9bLns+5OHaY9gzDhRMgYQBqwaXMGS0Wi/UfiJkcEu
7A8yeXcFHMLmaoRJTys+XNqL8kUXrXlW8Px8uxEM53sEXaSXBYXqghkHt7+dpfoU
NY03foRgDUwQJjfOsHxo/jIbuNFy3NkBARYMYcxmGd2H6k1E/6TOSzcKvan7NIdt
ePGEhelrjitcImada5kDGHXVMXW4pSrCgwD+8DuljYDFh0LkPBXfybTwzh+tqH41
qEJlPJnMCtB7S01SBDIOU+yq6iyJbICr+TFWhCUnYJaHmkkEnUbcwKlX13mXM/Iy
ebZ4oRDWmaEEv/2ww3la1lUWj6SAIebppvi+sTVQecYCbWIB+7L+WKegnVRcjd6k
EyUIxJhQAIRiZNnUDNpkxMulnk7NzwLoV2AwFIq391TFAKWsShe6ITPZDAZnqmZt
Cty7wA6C51R0VdyZnPfrdoFyw/u0+QLfHp3sN+GpvXs/MHnL2xiuAOnwKCay0iET
nBIz+grS6fiMWSyh0KFipbbFphplN2jKxBPkOdVlhMET2gbSn9a3K6rCPwAaNERP
IXDDbtGPX8kNuYKFIL0/OM8elj5psZDg9U5xixRGfYaIitgHiV22w1QIG8hxKgI0
UlUglNtEZrnRUU40vMxcRo4Y+OZUwHWJ3W97o2rISgnIZDX07OJHKBfHMSddqeFp
DgtGZXE84BwpUZvbusHWaCipMCTD3A2zKK67q+j4vqbNPfi0C1QlrzRayLjXLXoX
JkaoyS9FC5ZGG0qLoLFaj73AjVvO1YOrucFtKsGB0v7hCOzn2sAP7gR9gU6jP2f0
vNV5ESDnr8JuyNA9LZCsoaLQDJ1ZuE84TaTC9bOqnC1Lj9g5ttxiOBiZvOxDMCy+
pYhT2KYjAmm3qV084DEf9C0VrZKPoTV6vaFIepy8RHIHN/0iffx6AyktKYBRFZ7W
i7400IMbVtSEeG4vGFmWn9y+VYLoYlAox26S7IXAbaGz5eWz1KGgK/G1ck0AgfAO
rHeZotx4a2fGLKRA/qYiGcqOBmngQtQJ84/fl1WCbLvwjIi+LzIO6fvkXad0AMi3
yq3lZtqgAtROkVHEAnpDyM6rW2hhlQHpixOz31vTXQd47O6i6RKZqo9ocg3VDrim
E8ag6wqLYM2f8hdWbzY1sMLTHBAPvofcPJwsknZdb8hiPHPlYhV0bcg3Ae5I8rjR
BrxsU2K71PGbeCrcoVSj2wjupLJPDN08KgDvTVLsUA/Rjef2nBTb32jmzM+RYsGz
0mDpaZNC0yDEAw+PXzrBmfHSTmW3lM1qDRPkaJ9O6dxksRqUwm737dHpVO62H1Tp
7oZx9NBLv9Af7fLKSUb+FFlkb9QU3r6g7yKvp62aBBSZHXssO8SxwdHesZZ+FXgz
HS0G9894DOgT3R60JACaMa6BDLrJ2vSWlyyIjbkJFJ6JPEGCJYR0kP8oBZeLFgq5
EdJC9FEu3IuePCYLMK3Gb6SctDCqNBIXxdhkuvTQYrA9vWTgvcx7fpq9LJaaIGfw
hUA2WWI8XwEz25OGyor4vpRlVuotQwg2fSbOuTlc/83D13CybI2BZgJlCNuOk7o9
jDoLuEyu4jgOwm8RPlobyJsIa7G4POe1lJpvY3sG3ESv24maeMzv4PgigscXPhkn
PeKWq+kIRiH9GT8HuDq3aBrMQpTcxrjSolpxCM3DgxcHEd35cTfAeCAW5HZVy9/u
zKRh6q3WGY1Ct5gye8BLbk/oHZ9uZ7fTElNJX2GqyUvJfTUQIPCO5/DDC8LUluP7
8Mm13iu5NO/pIuojjORdtQxEDKsOi91Vg7ofOt+uKFcIohe6LY5hpbYcf4IqS+ON
v+QJ0SfiFiMO5oQTrgYNXiD5F26hHqoNtF4zl6TlzXtzsTjaLv8DSFQj/rpzDKhL
4UWn7U8fujhiucJbRCwauzBQW0VDhDHm6aU/JarUGMNZD9AYlF78OCj8MdTshF1j
AT83vpY8uD86hpf6vvf9/8oOP8vs9oaAibLec2hBkBy+8NYFVPtEWTVGmu6UVUqn
wK5AVm0eIrs441zDLY8xOtTp6nkwFXVGMFMKKKv5NpLEor3oq3O/zjptm6iBkv0F
D4ung6IZiPK72QO9qdFKqXG4zLVSxxTPwS/MY3SsESFkQhtqgfYjH/bkiyfxonEt
5R+pd0EjPPFFO+fVYQ+r6eQGzwVIDQtQsrWiFKbdw23hKFjORl6ave8IO/SRrQdm
Dj+VrrZ17HWwmpnrsfiWcLCe0noTRs9Yd3ROy+1JylLvVaaf8SXRWFL7ltFVHqNP
7H44cY+OdQcSVXmQqXeaNgANsvO/h3WJg9Y7IgsSgPtZwQdRNb1COuHLANDVry/s
P39zXlbFPu7TYvqa5GLUC3ZxfpC3R0oJGeD2rQ967s5o1cUnAbUdR9Ww0N6qomBE
Oux7RuPoECMZP6vhFOtpATGSqwrdQzQ9vYoSR51eo8aYz9ZJQJdxUBmR8DoFUb85
tLdFCVVesTWnSHD1DCPMI2dPRZFyExk099YbUFh/1vE=
`protect END_PROTECTED
