`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
orMPSt7HAP5ailzfL/9Jv2hysT7QVkIEBMJMXaYlo8ExoI8UNgleWPn/t4e/0iod
B9LZthXHeo+on6VPSeBEVmy/XrOThIbh+DlESJipaUfif3D2ONmlTS1WJ9zML90w
rqnSGMhP6nDN8eYEhzgMBM9+TzZWhNSf+WOqKKYWSCiYLWWfpOYUFU1RHjluZ75W
PJ1eamcSK0vAbRXSbLlWS0QR+ydJPaPL7uTVsna6geCDWM/mwX3diwl5fEWH/P/3
53xDWiUGi7VkYQvBWsbJuA==
`protect END_PROTECTED
