`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uoJ7TAcuMvFqBNlU5s5+B+/7TBk+VMQRP1Qb/3Jr5XGv4WZo1eEmSxyGXqUosA+h
5BWTpVz1+8y1hFHcgYA58xno54iyn4nf+fwXhp6CqGUsFnmptZ25EIjrzRvoenQ8
waGLgpAvhOJos6M6hqIM/wuwKoxga5W6GyqyQ+OBH29hvr5E/2uRXDvAsnn8TJC8
YO9LJeALI5OwXIPMPdIB/A8tPunriCIsUGufnK+R9x8lhxyTeJSkJ8exHnd0m6QD
COYJRbPS8NPFkbYDUrikHP6A9+znvfiHQlXCOeTIFBK4rjDgdKdk1YxjKVL1LIZv
si8nI8MUFslfenEK8HFiIo91ikhfFcIVhsEPkYhLl7k+f4fly/h2GiQA7hv4wcn7
Ct0QExeHiwNV1quLruiSZrO8qFXa68rk5qSSRtTEA40Ghl7fB0YyEbIAL6Nm4SI0
5/BvdF4v+WD34jVcNGocleMRBNI1pPtCm+wE5ZrcBHhXyT/tWMfv84E2Xh5NAd3g
mgRNnIRTmVHb8feIM+4WcoVLrq8jquuahG4aoXi5Nxfrf40a0N0f6q9ZZrO/H4xa
vQ03Clg78jEwlBgAj3oKyhp56axNiuh0liIk4Kx4waxt3YqPI2aeF644lKL+T9rk
9BBU6kl7sUy291kcdOnR++HT6D7eQF3w2jRvYAA3g0Ly5RftZiDE2bWkHd7gswLx
lyV4rcVaQlhdDzXJTMY/AlLcKRC8w/eH1NWCFnFAiSrNmRvLmTh/2Y8PWmKmcoLh
k55GSOdVZTzbbEcoWyvPkyldizJkXnASsL8lEoAGKdsfroX+pqeC0MnGj3BSV1wF
VpEk0KYM684Uc/bCsuFYXLuqee8eInxxplGlSrDh9FY=
`protect END_PROTECTED
