`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
52xyj6lJLJiGqcJwP1m1e1rGQ2hDELpispDlQRBm2YR4PbPS0RpNeb2ukklqmERB
3hxuKwbjMCjYL3oXfXGhfiGT4+N9btzrFoZ/ksG3VoUjV33kflUGKmZMVrKsCicC
W/ng8AxxXhUTPh+CEAcOCl8l9IQkjcwNsJpOcMIC9cax4vXFHHwtIafmzRruTaAe
IDFBPGNo/MMV9LDfdfyAhmnCyNdlFLh0sEAYbgCXMupDsh2uJChMGoNnCMjbdpGx
ycHBmlSyGs8SL6jf4vSZBuwFg/i3ApjGh2pShoCaPctCWqBkwQzOF47cGVa0gXTU
uiaib/yyb8gectyvei04Z8CiDY/wufRaWlx/Rq0KCYbjdvfPiZinMUiOGO9nhOry
0JqypXNovVSCH9aP/+qQOLYQi8Ydj0iM4i3E6dYMIAc=
`protect END_PROTECTED
