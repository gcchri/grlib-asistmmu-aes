`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B9cztoygxmticOI1Xd1+hn7q9rR0Vm66aVwyu8HnvEFtPqRcsRT3WFURbgrt6Qo5
z3nV3rKMzpQbWZue/jP7liyVFtRFyno3xNDEN2nlJHf+ggFAAe6dx28K6+gqYDAp
2KuJkOqY+BrBwuCp+l9T+IRWjT9U+9t9n3x5WRtMIqH7B9wdCweVQFavACSzW3uH
7odauW9Kq0jyuWY9VUQz5D9oHO/W/Q5v2aJF84kPxCmBQNCiY2WmEd7pLRwG8hru
bKUtN2G4Ci01VMsIzJhomEXkrEtKGlJTIzfpEZNyPn3pc5BSQzwN8+UONeMEcmot
uvB7ynccDW7xgAoZVW5j+7ijRom5bPm56dXnZEM8onIdbNVx/QV2w18BSxfb/BwK
TjEuL40INRCIynMQfOhhhwqQItVcAe27FeDPay7VlWNtNz97Goo7NFw5BaSVtlYu
qUSD/5Ft4HerLuFXwqzbEe8vnswTTgwoRLNd6PSYLpERmXyvRqcCMv59yMT+AogM
GgTZgjONGH/TfoGpkaqrJosOufE55PFuVUdjuUpIW/FDrXBc0cFwtDXBcq9PHUMo
08l9WGxMLw7Lq8Uf7AqNj/s6fRtOB/HSl0mzMxrJvS1fJxbBoUZ1okRlU9DZa0dF
DkyfhArH3ISW2iOiyqUhmfaEfQceJgGGrkexS8G9ruNGLIJINb9O/ztfYqkZfjMs
l67urB869lky2hgQZGXKLgjO2KfAgQV0kVgsxJAIaKj/xiArGyHF5NFs5xI5J9Db
a/IU2NRHcdVTPsFctUXXY+gwIBj0jRz1W8J6d6qNV5UtItIWelGwyMtuL1owbhCA
friFPl95ZIKql5YOTC/EOX76bxNaGYhCttAFLwIvL+Ls+pFPyKcfMamvf0YznMjs
135Bhj/ylLyNV2fmehro79pxcmJfEtE2gxQokCjhYtZZpRwnOatMHKBCmnHFFgS/
9vBxdcm1Q5MT1lkQ2CMxayvsg7r4aHm4J0e90Lkkp9Scpcfy6K38LsPEqkzqg8ZF
bmNYBfnMtKmTgxV+s8RFSRKR91JZ7utnRzLRtOjkAOs95HrE12HQ64hGtVYAL9SC
jGnkaIQlddm0KPQ992m0B3zg3SY0qYsuEJNJmxu1BT8fqhAdxFzMSLQ8fMRq44cK
yN61RkU6YE1kO8WWAOxUSEFqX2vPeLosly4ZVBuVOFSMVfvyIKZzoQtawOUq1lJM
zLyHG8fLyRVXSVxWdMLQWZAZV06ycOma0850yKkyJip2EnQjzDz/efR8qrGT75Oi
bd5lsFK7z0vriloGXLD7rAOnUfD6GY0troqeSCMidkor/kZyT+WZZfGEmQRjTYjf
MBcnKueFQXYgKmZQQ6q3AQ8GkPOplOTd+q/Ga1WN3StI8me4I5tj0jSJN8erwyBX
Z7HnVG9QqKaZeVZqbMsUUD/DI2NgUpBTFK7mu+yanifwjwt7DWTWv9Iq+4RdrxAA
Pkg+5JdytMTw+UtujDwjHXLuckppIOiBpNzWWMP1dIBW7T37v8QWRBlaGLcUBUEh
/zRvY2Y51LppvveDvWTeTS7SLStOq3676LAKv75q1hIcAFgs6W4ow4BRy69kJ78X
0IbwNFNYcF4QoIjOT3whD8Pwmc5lYJRJimcObVAc0N/mKOMpWFi5g8PRDo8qfCAk
+vtLX9Aosk33UJBfOOiELyDjpVGHmaD1ryy79FSq9gxI6CmYXXXjpHBmeXbrfYnw
FaJa4lppt8hC0Btm4JUN4VKteQ2yg8CQOub7hDHfyq665ZAV5Cr7Hmct939i3GSX
rZpnejRaofi5lpDtMsk0A91RgW1yRKNJUQPHqLBDoEFE+9O4JIEYGnYhRzG3kFqg
qwuRlCe54xNRKX+58HhsxHmAjPNL+xccQ+ZZ4S6M4l+h0BkL/kTaCTk2n2DT0jr6
gVlWoVrCimhVN5jtjfflKbwO+Iri4bsi8bWK0Xk/CBNGOwbUJWALwOlM7EXCpE02
mxNaLdeDtsgdfVj/pxZdNGBb8NpeJ9hvu6NJetwxGp/cF2DFRieb5yevK4qWoLja
UmLBLeAxooJ1wvWLa7wolltQVpdxLzu21FIfWDejnypSR0Jfm5AhMSAIVGUeiu1E
Oh+7+b3HVmTv2/6DpZuxOuWsLX1fe2Gh8FijY6eKV7ngwwMBjl1mNQLiAHUQTuJa
AFZoklg+aazmfUnUX7zbzU1W8D0asBTDC9CObqkHdycNRXQ3qy4jUazHXy7kl6tr
W/MWGREuuq8RmeeEFQNnvH/SpLWBP5ViJFjd26D85C9v+99GTXxMGsAc7nIIghux
AWaHXzO1Eaj8XZ3KeprgDpO+3WLoTGLM8EvWMCdQXh4U5BXSZXVw4cHV2JNQK5Va
RHIYUjBkZ5X2R3qAfRuGbnbt7lKJ9yqy0NIz6j1DJTHxtpMXm0g6V7H5MjQ9/QL7
Ao/TZSTUW4EL4TxUjEEQGcKAvi85Rt3Z+hLHFuiNEyNhNvgNkZNheN8fwZf1YLKQ
eQW+BzUgdef2sSQdRmzEH+TS1tzE9Rz4xckzRSF0lBtq6XpfK5qk/zcXRRjUOMZQ
kn22Uflk2yqEjonEwQEP1Vey+a2+795Zj26u/NsgNzJhQysOC8OIn7610NF1aTXf
JF7YWlK9doZSUpjuC5wSZe/fnP2qaLQYf+S14APYpfvdYiAc6YsxitaqEJ2jP5cZ
odpfcZx48Bpm687Nk/+P4ye8q8XofoQmOLN0SOzUiKrzfN0Sigqf7D+R0Kz32rCO
RtWRkiBVb6s6Wof7Ekrx8QidFB1pPbnXBLntmLS6c52i56VMSRbPMHISEZXKjgc0
2F827gFSPZXqkyfrXokYLeG0gVliN5vGkD1Ulj3JwItvPMAxwb5EG2RpLsDzlj2i
maafJ0/b656b8euGQBW9oubXWgt4YBvZj298jtZlcRSVjA7+avBMznSB/SbwKLq0
B69FPshhn24bm+RJprOEljK+VQ2wxyoQuCQfQ2ApARS0h7AW2FEJmc0+50nQAAvR
GhvEbLQsHIq0M6YPslP2EcN2yhezWZ8RWOl2VG55JMCdZ5svYM0hIEIh6vTau692
SU81zuR/k/F8goPfPnd+454RKEpa4Lmj6Y7deVFd6rjbNDSonI9e47aOFGrpqcBR
KvpeMhG6SoAgBusLBuHZ8cBQaW6d8WJfAPj3Q2JRSwmbJS0AVx44W2omi3uXy1HC
Zj2ZA8iFBQvLX+y8aJczOpU+xgnmZaO8uEcdXpu1oloWnRaF2lsFtTaNRbyx3NZw
LkbuV3ffKefTsp8OO7wDP4aAt9b0S/58p2gRy5fTyLkiYThsT5tDEZHrDzzKMRj5
4qHtI1H992Kasvi+OCCTM/9WycrL+TUJEzuWXxxx2E2PorxEeMBXisUD8YeweBwZ
/uSL2SEDVsQVyLpFhM5J86RDNuG0PWSX1hSr+gfqMUirn58NEskF9EJLfCuiWmQo
6Lemqf51DCnf06BFL6iROKj3IMiF8JwyyPsttADHKSfRAwmnf+HvRAtHJKDUUs4u
kIV1IF0iQLjvn4ZSpFtZ2eIfWbzTtOmBPRRBjFtIZut5aRVMQDKN9qjPTUL7SGXG
wxSzQZiDBfOr7O/Bkn7eb8kQOO1XhevcegQTOY5ZXO9SiySt8GpiE7rERpHhB96y
gco1gsWPDKkVdlyWSrNl59g2CQBeXhx+L3gbeIhNnlIlwcmae3TjBB9Nolg+Dp6+
BZzZge2gSdcgkRfirtPnNN52z+C0CLqlMyUYxGhPoW4G9MPy/g6ATQnj9MiyuYhw
q7oqIb+/FjJSZDVM8LrJDldyj/YbPkR+xhN0YAh85aKC+5r+9e2StnkD7ZOmQjtA
udldunaxB6G4+hPOysZUgakqm25PaWrBTkuj9O0kY3jZhlP4SDtV4wjWiJpqQCku
RvI8CEQhUv8iUWreUuL4ezKqrxrpnMLicGCy/7F+sOooJcqPdVJEtK90rcLtAVHM
EGHJzvzvszsSxxWZWKnoB10am58l+3K+PsFTlDZfk9xsxqiglNb0qf0QhWIZ0lvM
kY0oLas5iBzKnhMBylCPt5KjBjiUY50tbE89WD0JIW0d++uN+TbeRZlUj3t2UqCn
HWZuiSf6EDbUa3W29vOh3Zq0PjxyoM4MP8OhughURh9j+gdNe65OcNEJMqYtXiAk
yZaphHhUIfFqwv9aYx7gkqBiufvfxm+RJybSj7pHTIgO2zQpa/yxIwQG4SQhVE75
riQTOuVu3i/SavL8HplrWiunvRnFSZET80MP9IGwynXkvDl0gIUSK3fA9fJx7qOV
u/80EXejMwlSXksmtWQiQynlp3lE66jxRtwXNxjW05pmsiU7tE6zuKh83nwxEiK8
bf0/W5M9WnIId4wGiCnam223KKgvASTwf1mXU0ErvGAPZjIGczQVbOfyMtbYa/q6
vnckIOOvQe3A1V1HzkHruLgr5j1ro/9oIIL+UxNEIbhwNTejF7XrwphbV59MuC24
JVC+DstUUFLaoGa6mSwL9Lg0Gfyiw14MewiKuFhL3+LKwC31veAdiSbdHcz8L/ZI
b5MMt9axAxin8Z/Mv2QFVKnsMikwlBNkUBTVY4ZfmpQ5nN0kzso18VHU63ErU5GX
hju1dS1/bBET9ztmCoL1jnAGhLjSOCWA3h8EXIZcNFFZ6FvxnX5+8+pIZrxpmUqy
nWHpYpSh5diBaFT7hXX+k9k3nWztdlyikEZxlFnbc95eGDwuRLvv7szH1420E4XD
6XhFj+UkDyiufWGYclO5+uId/kZSyTB6dvt3gUd2RHg46PWO/rS8NYg1L7BdMIu9
cBHKS92ZvfLDWMH+ZiBHho/UI8QqkZWOq2OYzB4fcJxKc0Sb2P7syRSPP7gKxR2u
cnesyCagItlzVpXQhO/Lin0pVPAMd5D71VQW+koNdfExmlWaRrMQIcR/WVMrdA5h
PnEkwRFlHHXeWjwOQZUxW1ssWloJeQYjjMOMQ+4QmiGKsZOYDeVW6SGjIgDKTtvw
q5NVVBjxHojdWolQYC49OmMDkqF2Hn/iRR+oUQ4hRyDDCb67DfjJl9F3suO7L4+0
MVfQ5/NFrGHQPxs3/IGN5J+EHWLde78mralK/fw+6OQAcdSf7Udy3tRbqJhk3aQZ
87GwkZEZOeVXagSKVXOUneFuPIdqmdKBYkKZKNh0jbgStNeU5gG9MCiGedlT1g9/
oMwL7qUplPq6E9G8lG2BVZdh7gNB38BLyerSh1iIYav4gtbGnm1xEE8uteRjZvU2
vi79smrXnLE7Kx9UZU+TGt7joeUbveGkUQou2zPLVMnC9HWdC0q6x+iT/AHD5zAh
YsgIs5M0f7EryumDFiEJ9EA0E2E3JrWoLNS8EZVxelV44ibeaKNHyZ4uaZUKjIb5
3yJLMYYEmLkXcZE0cGEGI4p/KkflHgY9RGmcB26XfeMVtdfejWWKJOqLvRaY0OGX
2L+VyKOg0lAScvENlYIGQeXYzy++gh+a8pwPaZE4xi4QqsTX0lWTzLWFdGzDhger
tGbWiKWr4w5EYLFN8AD4jkCC+NgjxfRrHsRaQXS2UJxbcFs9QjWuFpc+TIai+ExS
H85tDkb2Es8H2RgKq5Z14n8UujMlHHhOl5Sy/8fSDy3ecgXOC31uJpDpvOWNElzp
oshKonaiNav16npzXeNgwHCmSZOruEWlkAi30MekA3WA4H2YibeuznrUjboveq2a
UNifyWJ8j0CLPRhu9s9k52YoS8qKLTm6d9gFhvL7VzYNpZIp9rHVI1u6hMw5oaZD
dwHhSFs8Ztg8Oeqs/BzOGOB9OLuI3IWmwp+PF91sgFGcnUEguZ9tMAQ5/bxZ1Yyp
3kF+iQAsw54IlQ3FKUHQYU3bScxbMYkyGCOAUqMYpstBhYiaEvf6vS3E94QMjBn9
TI1afzysFfSgx/oMyrlQzZcBtc5+ZbRYX2M9KYNVen76n3NQxIGqpa0xrFTyGmKo
OwPsLy2FxDjIm89DZ39+lyInelj6bwJ9w/e/I2oIYVp5uwg0+Cdx4IEhDwXT8Dxq
je93v4aSGi9WtoTlqo46gxNI0DE1j9pajj6tBepkyVOXbzP0m/L7/0kFLcqZNO66
Qfv3fLidfqSp8NT8hAR6a09hFTUwvFuvWUPrfRPrr65L09JlQmai1Pm3f1Yqnku0
gj5/VM4K2X8+rOA9KwaN106qyjPAXM9irJaVqoqtYj89n6CYJMDUnFVeyFgxKdl9
styLYCIxrMJmL9UXvo5QxJK4d253do8a6Af9gpGyuzBOtUMchYl9OwxmnAHq3tYa
ZYlwR3tbSXfTZjwT2RbqtL67nTFwWCh8RFfsbKD7SJ3PS99dQXe3RfZzzOu3kp93
VuQzddIXEkEowyZpXveXrfxm9GhxezQyPvk7v86RxU99T6ot8++xzjdUY8sTqTwk
PHo0lou36xgflM9f01jq1x7UcLMYwTjr6BAHadfYnjTXRh1lZIAkBNzD4qat3+PN
+AFq//kBokq0/TJPN8oik4Xz/1MJ9Url/m0Dmc7qEU843nxY6dYH5Sb5SsEVclSJ
q+Z/K9z3fnUA3u5MYCQdMYVuT9Uth7QmqNZ9xqiv4M7gH4xeu29XwNszhoHCzucH
OiCzRWyXO6yUp++4Dfmr++eBlag9JHUOiEZfIlviZE4yd0C6lBH0u90NBe+VOdKm
oJqLTJNPEnSdgtBZGYq+/UIXRi6ymMyuwkhA2PnacQDybThCi8kGUM2Uojvx4t92
G1OX19GSZtUIQbd6UInqamP174i2EwQYAm9aEKECVArmk4Rc+ViByNkddO+j93eJ
fldXJnlSvQCPVoXPRfSg36OW0Cc3ZEMDdXG7d7NYaPmzR5C09q2iWeWlzm0mrs8X
U6Jm5betHRZJ5gb5xGSgRikR5ZoShUAdxPM0YU8QGSwI6mhHoY5EEoG5w7lRdzKE
noXywn+oejoqxRVGUe9ZulHd+tRhInmas3V6uH/52+U/EV9DBK4kxdsyyqmYON6g
ar3RgqZ7De+6abmsEMthkMQVnHWwKXzf2c0Tlp0zXa41dlio6GCHPQGvGxHcGops
wrprPiU98PT60jCgwbvbaiu1rShuSTjqvTgZYStgQtKxJZTFW483JYVzskGfUkYD
0IR6Zqp7IZ5GcJcKFTR4arTN+v8V9Lo44/T/GySnhPVORy+raJyH5jmu+ZOOPek+
STwaKVrpFMGprRUlVelb4Nx7AP8+5OaNS3Hgb/iSQWeVDrV45E77ce+wu1VQn1Mh
VtlzO/STmr0X9dqiQw9wrVuPIIOxwhe3qYqRbzMCDtxFQzZRCA/aOIPo00tsPn3I
Ar2BTwBFLotIayNOe9OD8oLBORmO96mU0Rc8SI4y3drnVReM88s0l8LnnpASnqdu
sEHIn6sYyJ58w+ohj5jb8NSBgt5u8qn7dvN2NjrXwbSZ/7V2FODZWqCiAjUNgJYN
kRjDuzFMD2539uSGcdTEbole/CL8WNENYHtIZ2u2b9TgrJ58oJ+Z6xJGpNbaIbcU
kDA6923eLbA19Emh3kB3wedY71+ToZPvmki7uf5fzwKIaF11n4xjySPARRNzKoQa
brgcS9WFdteR4v1+4IZy94j3KPg43IKdGMnEq5r/D+omLU3hJ1Vkggqnvnwkp2pm
QgC5/G9a0zjoy0K8JorVWSMR9LUUBHF3S41+ZY4BJ2DbPheIYK4rtTZcHApbYawE
QStUbya53NNqyT1g3iotHzImDuvHzBGoO4c6sWlSvdT6Gq3uHA5KLq3X+AKpoLAb
BJwgIj2N0kfQb9iaKAsn/wPLzfVqMAL5ojO4N+7ohK2alxNQCUNVETneU4Ty5pUw
W/9IjO9hKuI6cnUXwFEiuuYsX88JUzTuWMp30a7DVgkOEmQwkkWCdbEbYUPyDdq9
3DFofJFvDxXZT/LdDW/hnBT/uNjodpAI76pyeukTp9uANgaIP4mPOKkRNMy0spvz
E8MdT+33dmOxnFbZ/lGfkVsEdGyfYzTjsROOaGaOEMVSE8RutzvmqepgSI6BTRKs
Ywz481GNQdddWGgVi5h+XkweRTfl5n0yD2zvYg9mYIepjFJWM/GFMvtsrrIdr7HQ
dL8s94iiECF+Xi/VyaGAwctXsc0Z2XHviC6jFFuedffteRadETtu4n8iVjyizvTS
/SJ3Q30FjNwhmyseeI3RSKT9f3wdYEDS7vBGsGfH+cMCnHCB8PJRJIWV9tSzrxJQ
LI+orU4tLkjj35asjLSwHehx9GpbfYJwkTmlzfplw/Kk39Z6hdJeXgTLYvwGHM4T
Zz03QqY+sCf7mQIv/nusYeGY6Wqd+jNAoPLQGMggOoYDxjNye669Ih9zcdeDNow7
ZGNmIzLXXSuFaadEQPgOBupsY+AqM6nUlBq//K+sfTIqyH0Dv9ll1iq/o49c5a/O
nwyU0qHLLNF+02/J/3ac2TSnYFEtibILEmFQGEtiB386pWebePrXP+Jdt6JAGLoQ
nIHr4pxF8hBG6OIf/pL2MRiR4Q3amDwgmvWhNSZMaY+vITvWovxlNz0AlXk43Toe
dn8dRWKy/ZfruVOFQz4pzOYJU48GKgv/5df+drwXC4KtnBX1prEdirn7zW4j2E/P
hXHQKu53mqC/8AQDS9SK/sVGSnziBXPZXBHhMA0o2FBl06BDMBKneJ9JL61TmKV1
Rgd/hW+DrjQWhSTRZKjB8SJFlIZHhsiuOv/Lq91oPToV9Uo+Sx64+DllytL3fU9R
BWFjcYtDOFZh0YNONL7cU88arSY2bIHrZ4LYZL2etOkqq1CYQgbIwjOwudzqFacQ
Y/CkIgONS+jvFny08q3gW4jPXH38wLJnUtfXekEhqHURskQqWU4XnxEy5MPvclGA
M3POC0nYgbZnFz6/5jUlX+Oo3+ubuKXJSWtaVx0Kz2L14ja/nkAu4GNv1wEwrX0M
6x0m3NTfsaw/bPhelcqIAcTImWaAGOUZKRCiEdrCAwVveyB1/b9n0BnTVXl1Sl20
tQygvqpy4kLrwi5qOh+leNZLbJ/HK76bxyRQWmW+Cro2KIyRHH5Q12c75PEtL3N2
ktFnSB/tzNb6ROOt/dwWBkiyob0At0Uy3Z1Dk433BzjiGJu2qfArxA0y7fi3H36O
zOnDLaT5Myazh4ErBQkZXMAvglOcX5x8BXlwhl0p5z0HFUIGc74oVOZDd+FKADO8
UTYjuBvP2ubnxPpBFnm66Fcs+NenXMmCPID/AWl04sD/Ap5qzQB/c5jvjaypJAT0
mzpwU0mOkcDSWRqSA9L6RfvQ2hiZFNC1INrIdFbg2SqqXpz8we9SSzDEonSm8Ixh
Zv03hra/Fq172OUM9oRoz7yWUstkC914ftUdS4T2VbaGG/v4rWzL1xRloAeWSC/O
lZ16W5MBJfAsj84k3L25ctl1ASNHDiGQVXVmPjTfWxsaNvoIj7Ywdz7dIlI94rew
kR4+SMkc2iD5oRh+vfk5JBRqGd9bJze24VuqxzpHdp814pwb3tvGxNM5JR4dDN7A
DUSJoukThhLXibclglFiB4Gex7qk8PJUQaDULTy3PZjtuId8bVms0tB49DyqmV71
L42B/A8CFcox1AJIjQpRvNvl3e2pP86+BpnHdh12unMm/Hvn2tkrkQW9l7djkbUw
+/woj+MDrNPunE3Q/DDMDjGsQHF5zcR8UT7XdHqg2NvRoS++h+Sz9GA2sYCAI/iU
J/Y6DOO4IRdRy5xSudvncgdbQaBtyEou5JPS1aNjY2cuGNFkOsgo0C0ROzeU2I7a
w6FNaAjA2SPfvrdH7n3Vn9OTmUnfxHR7iNMUzSs8ScLSOwatFmuYAY562UB3QKja
1k1Pvj3QvpRfPYd1R51NeT2mSUH9ZnGc7ZJtV1h3qTUbHuCUMDmxa2n99f5VmbZE
ol5wBe+dOtCnUStjPFwb1avyw9vJkP0QODoOHovgHIxut014GdtOL9z86fjEJP+r
3GDv047FECHkI1xFghFNJffFLmVRYrYK+yk9a7ef74TJ8yQ8iSq48CSSe3H6APJO
4rYp4gHBL/pCiWBVvlgKFKKsxOM4NbBqNvcOC0cy1yqMn3fJkugIYsV4fj4I0sgc
NJ+BOxJnxLOD3PD8g06v1Rs5xo41HqcC7msiyMo+rSA8R+O7nBviEDGFyKhlp4Aq
wABarBVvq00rIMipWcBixRQxSPHHTWotF/UoCsfwA1Q1m8jy2TNAqS0Tv7A9Ukbe
aJLuD96D85h+CkVYspTmHO5zKECXB4jvHa/kRySAt9vZJIxu0PukuUU20bdofkKb
y6LG8u9AnpwnvDJCTeLCpVuBr8yJQv0c4RH1F5vXyJ56ulR0xRgNVf7IX+0JVNIS
4IjvRqXwanKDCkozoyJZqwJnzj0uRtHb2oA9ovFIY0GXFfg71gK00lSCjlBl24so
WNPjUSrfzF+RA7qhr8m1GYG8cwepry5jidrRplxu4BDRWfkUG1HZxgcYdKToyP79
6m49y7X9MrxPFgvldR+f7+iDm0b9uHjCvRGntY8rSOcsoUee6fniBsajauWo9rrg
v8l8ZKV+jpBuvS6cq3EvgF56sfiEHYMtr24v8u8p0mDHHzcGR8UISHou9/JOmchb
bd3wX1k1Gfle0BJklmadabokyQWTbwIlLoV0Y5uOcbnSu+HNG42cmYLCGfU5rMNe
ESwOpx7KsLm9ciXvaX3/Mbi/tMwNLCdT14i37ceA76WKAZgi3Xke1/kdOnQ0eRyA
01K3e3gaxO9daj81LCG6KP5htxLVUP8wD+Ewz+ZYLViO1X5YIzw6e2RYENm7apPS
SvHb0IhR3dgt6/pKI8FCsoCFw/D8G37VwESgYB3BUs86SUZ/GQjDsoaDdZB3fHrQ
qKxkQDY5dfJP+DKVgeuoWqKF/Fpw9U20C+iDmmVVbHCM9lRWVoPJwXHFZSrOqr+v
5Sc8ZiPt8pxgt5h+ZFGd0OSTApbYLXxIJmD9okmhj8c0sVIokx0jTqDEh2S2i6Ne
xQrXoQbgnSmRgd3Vwa/O8EqTDpv2xE8lxNOQCQa3vu03f0JAvQ1jE8GKUDuhykZc
Ec8/1lgBo3wwHCttFH85D3pGOg5YO5lBrS2I8yxh41CCxPGHZtSaQ5N6Znjyya3Y
DGkvwVQVqEtUvKypDkZnWVPlycQQloizautZq15SeP3YlkwEDyhC1WCkOd0pQV3K
TOuPMzekQAhTat2lrn5hcGiGJ0pDPCLALiKHhY16WqXECiNwUUh2de0D5kSMNXGi
ssJOXQ+BrRQsbpEfYaNcVPgUL7os3rrez0xsqQeGLB3nee0zBv57mX0OIezuM0mB
hwmF0Tsi/Hej2T4SR8u8a4aacDeQhA4BHUHSooIHD1H0HrH6+8tAC0B4jgWdN07K
R30A96m1yv+Ylt7GYiogg8pqn3/UU31Xu8UpRMMhZtrrVAQUeeRKDfhGA7u1EOTN
d2fa81sQInmU5kZDMNcbfIyEDp8lhE75UQLlKVOa34Y0BIKR5yA64vzZ5luWZ3u4
JqZqgltyJ5mN5GWrJMwCfnGHErYJz/TMO7SKHgEBm7dhDNUSXgqOQcHE8iXeOkzZ
5/QMX+Gzuau86ckHSKY9l28YtG0RAXLI5x/AnpJSV5ddMrLGCZroKh13GrYy1rIt
Z4z5lOi6C+ABe/frccymR31F9RjBnC2y/NgBjrzBgrt9bU5Zph0aULH9pJV/Dmc6
yCK+0Kq0ZMa6e510K4OwSjKRou5gjpsn/SnDOt7AV8S0mMsThvMDDgW4QhnizBMA
zvTuJybNffqfCWS7OkSnaHySzID+0gQeeyoGn5tPE2tcEb59r482FzkfmV4MpNkP
A6M39+DWT50IbRJ2yLIl178hSZDEja0QuvDYRXpzJX/xcRMl0mpqZ7fHIwsqmW44
auIw8BaO4ZaV0LE9PFvPj0E7r1FYNidT7Cy+V+Ln/ncfZd6xbGCRFYik0d/WaIgl
9fA4mCAP/YW/khLsf2/R0ku5HgJxcV31TwjpCFXeffWLO5nZCpsXLAigPlJrYtmh
A1k6nh2i3C+QU9mWNqgiZ8nRp2Vk/oDhoVqKiX1hVMe2PzcaPispxK9va728WtS2
h5jjTVT8JiNvEAoyoCstQ/OkCOOXKHF6FoyLHZSQNc2eBb3cU8OJq/COr7cKHBWg
JD7aULu5XfLvR1EWWxcuNXyPIUGOEWlUXx9QJWhTc+URuJzNpg8oQb23ZATlwYsm
r1P3kSLksJkX+gDOJpkJPGpylBkFPxXYtSAM/MpbFN+EIqyEPu4IWXcXPEcdWRsm
H9n+pFmT/2LXn5ARaAwKOr6Yd7jbMAWzjnGo1P0T5YOU1XDaC+KVzTymcBl0KX07
Uh+7FFf42+Prl2e9Qh6kiD/v0a8KD9CNGe7eWua7pt1fHgxzlDSbZ72eYn4pIZQg
Cvs1wP0c06kD5QmDIDUuUODdbvZBneXP6X6wfN8N06/NSt/Rl1a3hCjl23yDt6aD
itOV0RmMyspX+6ljoX6yjCr9rhruS8kk8LFkH/4C6NKr74P6NI9fqmgZR8Yl6Tv5
S6tVNX3PkIy1PJ8JXfC8Rg2QO71ymkrKkXiIR+wX3sAsk7GULdHVQcI8783STc1/
/eGiyEBvLFP6YhElGSC/mLUMpwThPj27bBJvU9C+PoUBwBtVI6RsN6yaE7MZQBt8
iu1Dy9FpQBIOhet3TbNSjytVyW4vRcs5ihramWwIQVNCvmyH45jog1zIgxot6k3x
P4wKkU2kUq6IC+L9zKEiybGBAfr2gkHEufwrjKre1dWm+aCWZZlgEoPUG+d2h7/v
juzXGGrHfpNs12HbGs1QH5PpAZPC+75No3HxnYg349Jlagz44+6wy5XOYOpRMHSN
fzc8noBIcPDl3wnrdaHv4ONyvym6IXdIZm9RGZCxlUnM0Ttuld77mgXI+GcrkNVQ
M4DdHaN3+39P+qzGB6XF4WmyAnECeDpAdupeOipy7tkR/uGNbnohP1G82LsSiLGx
cbwoSgg7ehWjfrixwUW72jsaCmo+7prA6odqqWxStery6HuOlqEUmu5HTULfZIf8
YsnBf9C5Y2U5IaXtMlskHFe+u4MslJr0MGLgwDlxMaA4bvk0c7LEBX1VOIJGOjPf
Nd9x9W1vNGaXmkgbBoH4HklAVBNbfjvR5Y8GACX8waJ10eBwNQPz7d+cSiGafGwr
kCNUIVlw4/5vl+/giR6EveI/AKwqSlbdGk8a5e6UH8rEiY/NyERRiowUPZQeJG9e
Nq7p1ukGqMHZMcL2vEMTrZ0RUZ8iqpTQH+eYvNzesLM1gfAZr9CM0L5yQML94yPB
COX900Q3U5Qqgwe0Ve5Tq3W2ONSD0pXnCqNCzfD8jMPNBR3HqTe+ekxZDggvW8OR
2JlQj6/E72lfAHh29XSdAtm74x+n+4SJMBLhq0pU8Qar6W9R9fTAamXioDqepqJZ
`protect END_PROTECTED
