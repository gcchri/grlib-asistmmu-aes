`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GoQDvjYlyBc3ttgwdpI8d4GOAE0PVto4sbDR9wAt34YT3jZ5IXT8LLp3WBDJLjgw
UH2txbmzVhS877R4dCDhPv362r/MIzI1pSZfu7l/4r+tLftbTdrTDsJLc/7YZfJC
ZbU/NZ0mWLTcybspbc2H/0STeMJ3NRNZvK2dp67I7w/KWwE5ZwXzswJHnTQzpWMx
w4AVezRNE2rRxlQe/ZPi1fC9Y++A2xDiyjq5V7T1RadMMSJ5YYpi8qPmnPmzgriB
vp92AvnHT2J4aS0MAQ4MW+Al+Pp7WKliklWdXpUMDFJ87iZWTTmww0DoabP7yyyq
i8tJ8coKSTJVmwY/SLwtZDa+kwHra07cp1qOQPv72y0N2PMSAgfkG1IIAv82/O84
L4KoQT3y8nxdACS5vuFy+6QX4j0fKdGBqIntjgNLqPPGc/ZXMxbiWjHDIpV3sw87
jhibllyN3EBpdfUUTGXhO5FS526CNQStED5PZVZGjO4CYwp/R6liX+wKHAlS4zQg
PJkmmpjlf8lGZAdH/1IIa+WC42Gy9JhmMlWIqZxv9aTI8is/7jxY49MqD1uVYBIO
XAQfn3aMFKsSLA0VDLLo0uFhuB4PNj5HssAbaH9K9gqDzzp0FIyK3jTsnkixx0CH
nHzA9USqfMXawlRCEKcIwEi3IJMJdKgKNENNdGGu37rliH/FAxmSNPid7JJBMBqo
GnQkmoyh8vcbqcqHDqCgN+F7Ksha5dQkC1h4rQx3lAsIsE8mvUoDqqjmj+OG7Q6d
ZFV3X6UEzZlNGTyA/CblP3Fie2IoJkH5jpTJFz1BfaV00V7Lo0Yby2XQAHk/WL6G
t27XJo7eNOLoPPFQ4kRkTTaMpl6htyfafDrkefy82/qxXnUwG+6JePBnKTy+L/ID
jI7i7r6InFp6DFQdfdDbqbXAeijcOE4Mft5o1aq7XkKBGsv2Vy7r7+d4DRSpp35+
ezYeh68tC8Y3MvefNhBzEBtpH62ZfgiEmuqKkPUB8fq0KRjOOdzbzMMMdbVLnH9T
NlSk3BQuZpg7g8yivBiT6ttXCxQbSwa3HCZK3Y+ngId5OK82R8epUTXJD8tIAzGH
Ve9xdSxmnXeKLelcewdCt0YmFCBzXfSBI+qLZkWsKkypNrWOUyRCvgmNmkdBw9EY
YOWK8sgHF6obuVw1gXFzKeojDVf250PS+CmOoCNkN5kVPE3VqNLRzp59cnxNBHGE
Kza9Iaz7iYzOzRVN4FLhnq4hwAhGNdNlWpnPoCM6NuWmpvyGnVAP342XxC9/UoQL
sVwSqP1SGO2FQz3MZ7IBD96Yuie6h1C4rb1wmzDPsPOoyYDaf5hEMK9WiQphAYUB
xYLKwFnMK/WEdYAZTAhK16x9cJLT1L865Hde1P8gsD/4lEIuHPvwaFwF9feMhTy/
NdX6/bwbf0UmJ33Qyy3V/eQz/Vl5Y7kH2RPDyDLLX+OIVUvmtydeN5iLgSSwf616
c+MtnXDYRuEgkKqA2hXeiTHAUB8oum+zHA9KxNuZu6rjKWUR9MUj8cxS6Wo2LNUf
dBVBS37C9fRztQEPuQGJLdLF5XRpL8T5dlGDY1blFHvOhpUYyn0KowOFk2HqxsaJ
ueUktjV5q3JEz4FZ6ngBKH0mB7T90plux/DGEOvHxOrDyrjjIDOdv6plAE0atAst
FF/jwb9H6VpztsOPXunp6F+k8tVfB8oHUJzjaRAa/AJrg032ZJRl0T/oUzlV+lAM
3SJw7ljdw+B4wBTljHOsk7/2W+/MGFWntb1i8pm7za54GR45jwPGRxn1UVx5VUw2
BnDoQq86xzb1i3TDPFEWKrxemhvc+ivceqJzWH3v23eNEsVx9/LjE6cx9pctOkwi
9ueSexJvroK5ADRk+09k11eB/SrSVPL3PGe8CJwdsu4oEWejB2qZNlpKwFeaUAj/
jOSWBo0b6DwprBvlnZpcZ916PBo0GOyzVHVwu4aZb30SfgTCYarkQFmY07vh0h5B
D1ZWjR2iOzx2LOp8WRWQWb19WX84++/lf/wrRGAtGWXAkH8qAiFs3fZUGHQRjUIv
WCp8Opap1E9qxZeRs8gGSdGWgYSelBmge0/bNKyXM5eAJinQICInrAiTBwGp5Jue
2N3ZCbmSk3ZJkIAzE+kVYXrFIUVGBVteLIR0XnCFpkqoM0ygRPW/glJS0UIlMeUo
770i6VJ+CUC7GGBat3dc0r/9Ss0Cr+MDrWWlaxLJDwXoijqVHDHs6xawd5hm7EXN
M+JClaFanVlYGLQnM+94rOqtmXi1xp4YGp3yStv3m1FqW8AsrzfAeiVu64GlasGa
qOY3ZAVf2Cm1AhvVZiqwP+cwDOu8CkqtdHSTkdDnd7Ht9GgjlSboikv3Pnu7j4gP
FKCZLsr8/fzJ2DbO8DYBQ5ys40E44xyzvQ7iwWHPxJYG5PJUIU9Gamy2VQtYHzz7
w4oqANuGUBJIKZkA83cL2j5aDKbhE0PhgYlyIxHePBit4QkX/crC4x/W8e+Xilta
7bET+s41sLzRgRLu4GpRFHUmKvogYmQNzIG6vj6X5UOcXbksVmK20ftgEfObzv6f
b7NTXyWuYEOkDoDo2aEGSuutlA4lV2KIXNKNokf19CvN2TuUTX6TiworphvreWjS
HimpGbTwm9bqVySdM8siZPgYaJsOeqq7QyFdL37AId2cqg0m9Ou/Dx0o7Dp5AVxq
D9EMX9vHIrVZspbYYs07H+mN5ertf/A6NNWx4q8FHrpqAzG2Tk/Rqqgkx7SUWTbV
C36FE/tp7mWlLBI1XGPGftPkzFMTsMqvfVzfE8d/bIUCYgbBeETL9clMJUCgBYwT
WOVxIYF/9ppLOOx7SMkco3k9/mXBlU0aPUeJPmycyL3pZK7iF/BEiJcMoiq+N5TB
y8SaQb8ltjKwzaxALWzbxMdeRZxLNVRjY6/WUaJ08/o4nEqehYHdgUDdML79av5/
a5TTRIrC5NvyydDeVaKpvr8RCgoeZBrrAeaDZ2S0WfvWnpwn9F87lfkn3ZhbUmsU
YD6AGtTWvVoglfPtAKUH08LU783O5pJVJiKNndkufAmcEKrP8bVMRRxhb3NeOIj9
fYkCEIccLBQ6W+cgBFoprhhOvKnVBogFtAhimBgCBvVOKmidjq73iEmdBTNjkpnR
/5XRZHJrJHVY2hurIzzCl5Okso7vg6+Xp7wll2alH7igEkS0uZ0uNLLqcSC2r1/R
E2vusJJJ4b/H91B1R8sQ0AgqSvzgWInL05eQwP6OxPmqGeawflek7IVBAAvWFVUi
/CV9OfL44jbprsop4lvz0LbKlgP3lmd1Ph+Fh3k9jS4DfptLUDR+udwnCdc1N4ze
8aKd6GJmdD9NPA2ISIShDiyAQBGEwQVLpJdbW7RKgMx+2NQDAbSsno44Y41RFCA+
X7YVSQMawRsV9Vm0AUU2rVIfx+xjvzWKTcrqN0SbgE/8SkekSNjLIJpdI9VcRmvW
VT573CKhFdbHEz4YoMUxwa0lSr9G008HcQKYKPCHZhPvNCwxO+IpNC/qc7EYndV4
7PooRm7XDCR+uLWIkblzoGEfmOmgS4h8EtEU0fGh/A3HPfxLB00vvZOaD9AAYTv1
lBRiZSO1QRDvaaWSw+mhHnJWF0qYR9PK/5ciVWl+qSoefYwmSbkowmxT+crtrWuc
lad63qQAw2GqEQlh34jF/Hu/FF2PQvg6lZLz7ub7Z1g8k0cQrlMP1kGEaMw9yvEP
K9ksm6mFmtQVMb8fgIcASTR+tvmO2kogbtdUmxAh0eifyFni2zCobOxoJC8v0fwW
W81ksNDpmCEBuWlOjUKpZRlhOqTG8rTO4yIHaDM8nI/MGXXpsW07brJgBy9h5EFE
NIMEMJy6ZD0Arn9l8j4q54mOTiWv+9erl/rooV2X5gymJlM1P0AftGwaTCfHPcT5
zImhn9cbn0UY9hTqTVX/PO1wHyNYi4hCwBsrC2h4ZIg5LEKaC9CKIgNrF2UjMiDR
ktXbfRZ36RkWrQpPisGhyHa1pwgTl51kNRGlxqj9RlOoqlzQ9H1da4ezsqk1huVu
xNZCeBBib4ZNq0CCl8HGpjR99eSyozlp7Rdbjfj8Vma7+yAX3aWLTDBLxgMcBf4x
6c6KQVJnw2PO3GY0MsWz/ZFW+wu0MIUSPBkZw0G7i0FkDxfDfvhSoNcl/AJustho
JDH4j/xtIdil8FKOh3kAqmBSHhLUoZng8g1nkqZgPaPgzDwc4u+N7Zm9u84+8n5U
dfV2G3Zd5GM62B3CunLRDxL4rkAak7hVE6Va/DIYNURmlLkF0GozYxy0sxtaUnce
ol/fY4ncIUlLEJhYUMQlArmlQkoZpgt2mCWZtNGp/zGl00opoAa9J112bmjKWF5S
Z5GopElHEofveEOtMq88zSkXerz7m289RbG6V2sFd3HqZQ+FurN0hAzhbqGLbeo6
xhKZWgzQRDgWn+nhHuEqRDoMlP4N/keuJ/B9e8nHcDj7vZ+GEXw9SEjuXYsj314g
+/pAbAme+ud7+5kUUyqUdVXN4g35bvO8d9gKMyoT4Keh/o8BcAqFG4VbKeem7Xk2
tD0lJp/bZ8L2KgJ8JOTtLLjWFRdN2f7RDnJCIP3hz+5b8t16mrUpny96ZquKunYM
sYJ5EqarHK0Wsglu1U/38o48RKAYLB6Q1vblZ74QAJXC/5PsQ7PWfMAjFLuZe4RM
YR1VgV1QWIfdFsG8JHEhS5lLrlHzwXY2Hxoxcu3ERU5T7JI2nwPBAvTQ1EVrpfGF
wi/SSuZY1fqXVtm4vTw+BnAuTdeEFObZZdN6yTufOxaE3iaDqGY/hob1e1pSo/wy
f/7CWECdbBTh56MBrM2nNgdh/MYrdwu3F7n+2KqqqJc3R7H/aTMTzlOZLCcwDmED
jxv+pOM/NLZsWNPXBObsGPy6ey5VXfyiNKh+qk/AqwypnMqmDR+6MAUMpWgnEs/Y
ySiqAMEFbBlEAOWr5U6fwg5qPPueDDCA6FFmb4jF0LhL6ooJNQi2KxxMvgL8V0to
Oomw7dB7n3J0gqtqN7Xc+EZyL7VLodMg6snlJIFkoX7oL/Dn+v5OD1mbevWmkUjQ
/VM/QZEam/ru6gOk+pFseLmPSUC9HyrOjw6hnITbAF8U0ka0VXBXv9ujvP4fzUP6
RyQ8isV8eOKSXX+S9Oxj/7O0dAhQukk75qKdtZ2fll/jgQmOD1GtgHRQ0Qyv6swg
2GdbRLecoo0DHoqYoXiM9Uk5IJCabH8aDhQSxP9+aVkkkMVX6c+qx0OCQQUjuSEa
PuwcCT6oa74bfD8YRWGreVBTZoHd0frc3HVyuXPKj3sse0Va2n621vqQJVL1i4WE
Bflc6datYJWGmJ6+rSpkx2MiQjC150Ps/o7gFUfn9wAGA22+bGCU0sijW8flK9+P
TbM5sQkJHZsiE5lZn+GdBOlashKiz5+tM5J4rOwczbbz0HA1yUGGIoPXI26CU9HR
Aa6/CEthcu+1Od+AnEsuGxJ9oYw1I2RXR/zi23DjFGm8RpsmqW+AgNgJx1Wc3fwJ
gQau0XWYs1QwO/oUEZW3gCa3248eiaLH5YJcO5Goexsd/lsRtu153G8j6kors+hF
pBPJqh+tf3iOB3WRdDY5KBQ5C4A9Ieemd5HQ6YNv2muV7Y+7DtRKK2WR9pmHto3U
7gwQObPLMG+b0h3Zcw+hZXvfcIEVApwMLDbzmvHW0TLty2bco9EoshSlIOkUNS8y
8o9aA23BdvEISjT7RQL4bLmMREVZoCl27Gn57F1YZ22WcW6mjBmx7xdkMCNR+UlH
ySzF6g4bxxic3eRJRasg3CjradDHovRR4A8Az8qNLKttcKx7lkt29p0Xt7SahpXU
iPWqlRh7UuaDiqSD22JGqwyDE/bYOVHGR0i2PzfFIvZ5r6w9GpYKa/H/C7cVU7AA
FoBpdThD/d6wEPtUWSRE5Vx6o1ACJc0/9hR9uEjNmjVHbD0gOgvLNP53i0s7DOPE
qpO2SClBGCzQcwDYcHDEM/Pd74EyFtXb38y+C8wMBZ8Bk8RNUYktd1ZV8iT2GSHr
fDx64Tz6sEKYA0/V8VfVE4hwIGoo9saoW4U6SvbSxRg4WoVgMzuic6D2G8vQV9eu
f4Oa01lWHNnHB3ZbBa7J6M61eMpkSPJvsh/qQwqKM4gS0r4oikpT41e//qZmbZy8
5GnfagDurKML/ljj5XMEH8Yi1TiwbQPXZtlSCFn2ars0fbSJ8yNVTyXgH/GUH/vB
kkKFQpG2/p4HU7043NGk6AFXCLpsbdyEONEE3dtT8JMV2uETavi+FTK21VuvQ5/3
A+IRe+eQfJWZLHb3pZPB1o9VfsLlKPTRt3O/wnnKMbLPX9RG1Rq9yHbjs+k5S2B3
cYk4pQzzS4p6y5Fx2FC9iRgY2Dh9STxLWoRABoepy04TK8DY4PIilPWs43IFt6qn
lwrDpnH2Wd4RFZkqjoLj6ntuFa+YnZQU4FF4oQWmDcxrl12cdqCoB1Pam1TaS7Go
CkNyKMlXd4ubs1OEfpMGPD0PMIMqZhyR/BHXtnV8IIE2YE4keAplIAn133rCH7y/
4pkeIhDJmAvOo2FQ0H9WkfbWdBC1iC/nx9fOV19Qa+PA6Aq25eLIbXcxRi2PAJyu
C0BFUVABrHVZ1YH6ZjvyqVKLaqXKCZycqYE9sPAcGBQbBKgRXqACu28lNSikmto7
vKTsAA7eLt68nPWH93mMSHeYNEACNgkdEqvjkm6L9LeTZw8iyD32aGX8Q+J93fA2
4NqM4/hjO9cLYaWUX60b/DjB0krlislGxeI6pJYzJs98Af523UjSQGOLUdE80nQX
LyiZxhNbFlVmIpa2W1pulnvu2hHsjjDFxAzVKu4S3vWrOsLlCQ72+fzIi+OQTUxC
2g3L4zFIXKOEXQHZZegeBcCRau3ArsVGposy2fA/UFBftK0KBusdF31j51g+F/El
WjcK2nCi21rUbHQSQzOT97MtgXFqDWyrAmglkM03Q4BIR42rJQR3+1GsRzVoPKzr
jURLUgsPBeuCUeYLtJZYS1J3xgdfhdv8zVmWMSd2Goo+LUa+Efor3iArJoJdaLTr
gsla+LJeHERZxb271tgn0JDUKIJ8wcPki8mXBJSTXx6PQcxCnaEHxFAvrhkWQGzr
WKYxrwtn3c4ctV9KFIHyxV3uDrRJsH92g6gAdZ5J8+Vy0PcREuyaW3Y4alAPtw1p
GEh4Gxq/klSgak3OYedZeGaaUjz6VlJmqIs+33ea+GwtzpM9330icAYYwYdNpfVy
I5zlyS+afo0+NfGwBcQaA4Pj17i30/BlXPo/M5WP5Edh99mnmi8C38ucAKedEm4R
bi5BekroCQjgYBrDFMICOT9HNRxx9M1Yq90YVpd4PARupq06CSyCCbmcEco75EjU
KbnazsWxL0DrUurwok8xdT6vZrMX9ha7V7fzGkxV2TCo5HpeiFjC2kp1BnGHp2oa
tWK1fnfiaLcFHqriO7hkzjnb5ZAR0yfM6E9qyA/pUICWpm1C8Dse80mOYuJneHl1
uBBRKlZMUKzOxd2kKENMSM9HZT4WOZ3DFv45vNb+5+s1F5TssbpzaJEi0B4XYwob
LHcU4wZtb/Feklue93pPkXNU6OXkIVtDZgEIc91MbmuUC2IL6YBMYweleMxMiCCK
QLukdZP/e/toCw1Gq7b7/q1rUlutuT/asI/9KNvktrJ/uuyeoEQVcK/PqzNFrPJs
yxAtOC2U6mE8YdCVzNjdETfmEYZdVzd6Khar3zI0HjerndUexFrknNUFM7i9Ka86
eenYoxfFEA1Xj3gJiD9B+b9Xd01rHhQXqPpU2KMsXt98geruDwzACJYYZJ+g/tN9
Bs60VHc6wf3mnVfoICD36cEty7tBfMI4qxUAIG8/21Sy1xE3eBtpOXsLtffaUdvk
CPo+WtMwjWC1nLaEy5njUlQ96G4BqdP8chzbvNnYnmJJv/uUvx7SRvIS/A71wMNb
fMPSfGTfcsILAGHOzvem2lnDBeM/f4+ZVhy6xHjtZwd2kRhPiXTyij1OwOhQqAYH
syXxZuucW+tARr60HwKYvhwWLqUoVJ5ffnZEdYZcewhildVUsAyHIqJlbxQdfymy
thjuE44ot037ZT4CnORZ3Tqf8Ah8aD3DIcey03PPXEIBGbVyOI4+I4ilhxodPFNJ
dY/P3w+bpOAo+c5AlJ2d1HPOff25wbkcXPaLSe/25Gy3P1gDTz9fYBbCM2/JZxp0
CamupsM1htu2iLTFW5KXpCWCokUWIhMbCB7KcKVhXXwqPGyUK/m9RuXEP+YqZ8H2
AtrJr/C9jyhQB9k82iETSslPQ5T7fOwpcvQRANKTAQAIL6iRldoDGpCPBf3TGPKJ
iPIJWe8QDMPw3DgnMn7wId1hhXExWL6u6GnjzCQSvWg2QkJ02bVRDFXKVn9g1qAm
xRgU2ckCiaYJTC3H7Uf/fApgDJD+GlLxBvW0mransILx6SJHfPQAuUxbwScIjkh7
kKW8ZvBIdNNhP8JvmJPLnjOnJcDdi+UpZZUeuaYBL6fhdNjJFRYgDwyXUEN0rLv0
NRlhWeLUeqVnOnKEdYre+lKNgDEhc/L1D0qpqSvarmYS2+NG1nXDMennAFA1FWig
s+FeCOxXrsXtpX2jjDgkrRZfM888HinSpOdxdQwrEczJRfg8r4aJb8SzhM+b0ShN
Z+w0Ki/nBkPNluDec0eP1Gu+NMctCtyQEMhzxPMesUr1FuaG5FUbJdLBnoVw8lsO
dlNuof+luKPZn4N77kjlv8Yeya8gby62QLMeX4TU93YKOSbuOGomM4RHGxcx0mpF
iU73HFatO2grrKxHU5ANh4a5+0OgaUb8DALoAer0lBdUEEf2hKlgXCwNGtnj5hBg
rASIbkMMEBg2UpxjOr7PQaLcs3jP5kwWhqKA2zlaSXbRnSaq0ZZNzFk09ySMl1zi
v19iUEy6cCWQgOnBhGoVYkd77neZT/59z0E+yit9EmjRJuWkYhNNSgnXDaOYM3DH
1fdg7M5JqFGdX26ECqpqnDPLG37kxHXXcMIhmLNDS69h3ykppu8WX2PAECDdKUw0
gGMZohv53vbgYaweosfKxUC52dTT6qvNrDiPE7WhNqRIIDQ+1m0rCfH3mvWK9O1i
wsSmExWAbvJMf/j6mDuVCOh/ckEwFyVfv4/POaGSIuohLTLfvqaA2NNMNAKIlB2c
7NHKC7FlBGoeFWVFoooi1e8LCYKHeBU5N+yaXEXRjQi+zpuXhGlz9tWXrm4i+cwj
2k4rXHqKPEKJYFlht0zjrRLJHUMnYRWfaOfRQoqK2BRYI4rDeuyubCsL36uZWywb
9rio25HoPcdbCpnu/TVTNZ9N0TrxosgR9QM2Uxn//qd8D5dqcUdOHQsL0ooqdAW8
vSzB5vRWEZjXUF3UN70khspzs8I1qDnvZrLBfcfhKYZYG+VWmxPF+UuHvyY/YdR8
JLK2WwBN3Y41hZOMnTcrc34uujxoOcTHBsvBlMpYYA/D3R8m1+zY2BAV75k1Kunh
88MHSEZrV8/I+zMvI6ATUPW5E1dTi5iTQMXfPUtdIqHykycYM9eMyyahKqLYiZTN
6DDsYrjdWw9/1tivIqa56tYL8qoYH2AL3u/uIES86GUAGJYQCRWzV15D3sLucKBy
Ypv3se9EzrSQTmCUwQ1TvW03RDKWsJ4aF1trqukxEbexd0hQo+LNtkkYk4CnCvWk
ZTsU36RmgTpfOpCx5FArYZ8wuEQfGAZP7Ly3NxH/3tAOkjj6ywL6Y2sFLOh/LxLp
aS27L2/cXw0uQvu4+cyoVScDb8BYDihzw20vy79iaXpC6awjb5UuzEBiz6H7yifX
ipfaJriMYmyfLiXQIle58xHjcMcLYpi6adwwrjzlZCePmLeg1Dq0t6ODfv1kLkCV
BqKK9tbEqDpm6OApdHSCG23lzf9luKnZACS67mPcOjDoIrYCFPodTfGpjQWw9jSG
BnEOwgvH17IyXlttsidV0g==
`protect END_PROTECTED
