`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qs/3x0nyyazMuLpSLRc4b+NJFI+33DNoxWflhq556iD0MnGARI+kwmhMemks4EKX
cP+BGLXmbt8MkgKprzAvcttrj7vipjKI7zU++SKWVSOseaZRaoehuwjGRq3hYJQz
vMWpJe8Wr7CrCmMN7plM/WFfiVgVpqN4NzCO6l+FRJNwLdu5SkyaOz58V/aTRNiy
fLG/83nRWbMRz84O76GwJ+ouzEOcDzNDt9eia+pXMwFDUk6pqX0xezDskCV73LIb
ruhNcJ5KCMVrHSi+BDifust20fVRI+ueOs+WbQoA0m+03MMKRuD50rTD/i7RD4tl
v0YazW8mMk/WJRe7/exQoWPyXylZ2PRdj9kQR6l4SF6rfhlZG2Ds94AkzakDp3xS
J6nXjdWF5+yHaw8dEVWEXbeN+qBPwqhLHFPTEoUTmWNdIxV55JCnRM0rrXZvwMYD
th+nwTs83H9uD6sHrhhNIRLkh/KMZQQZH6b6VF3JH7l2OcFwh6PZYEp9+uTjZ7Cd
FmmbHlghK+N2H+wN7x+S+fnmtX7+Qp8wOPuaDZaS9u/zUDxAONqSQjgOWz8614b1
DA+HgrIC0ducuX0ESjlA+TswpJAjVnnl8CDG2w7dGogqNENTScj9VvdFsDGCtHdg
berQ+nr3RZOSjsAKP8KYFg==
`protect END_PROTECTED
