`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fSUV4KrzK+iQ2yWup0E4QS67H4s6juvrDZ/HMGVfVQDmQTKOh6w68ImMjfT9k0VI
LcHFElHssTnVwnn+kPU4qx5FgQN/juiVzI7O14I5vHS4ixCJLoY+yRXxi6qHP9ZH
mCNq1uJhBEZmf16gJfgotU2NkIeBjbjsSTxyTJeZSEQX5MFgDj4YHaDyhzRQfhnZ
vJcNZhRdmD9gtLADkR0Nf04aGbJ6VzzMhbEm9rqh1BAKcaIDVKRYXC1NGeSzmQii
AsngrEM6RI2G3jEgPpLJfqJ/kqTHg/o5rrzrM+CLDFfNUoZ+2z7tXzs3oTa27cQg
bcXOOcYT4NBU7BhLFbyF0CuqyMX8LyVW5Oh0e6x5ATMjPCduf29I6d3xZwE4m+a7
AVGIVs9J0m+oGkBgq9UtqOMc+9AWoKuIuZcLXKHZuVIoRz98wetYbfuORAiL9Vzp
SGD0F4XfkYiR6Nmfu5d62L3vRUmHHvyIilS/3QmAj05fdQxHV6uMjTjT0Dl1sHz+
YdF02zAH6Sb2BKmm+WoA1K6OthZPJFhp0xLNhmklYD3rroUiazmTm7bNNdchqtVn
`protect END_PROTECTED
