`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kGNL0kgkhBHEyD3/ymWqTkAeiC2EFs8QrKiLNFFtr+FM4jx3L856EeDv2Su39lWn
yBz5AnERS17X3B8uinooGnoIqjFgXl5YQ0XJ2LGBWIekMF7MNIRemxGjkbUBZhbG
7/qdlYemUhKe73oDKrrg3DLtZvcNG+JflP1uLKvow1JTiLDN13jcYFVO5piJ0YVi
8NcSwHGNjP6hcAOiuiIC6sQsNlisPP/6z4Gk6VQ2qkPqlyw9M0lmn5KpV5AXgRJ7
ybzIXGKKRPxLNcSnA6N+HkasAEniXaJitN76euUn2xQWo4eFRXhTPUJA0YZbkIu4
766YN9sAaExmNA1xt8XLLEVfG+aVNMHZD2PvxT2OUpPp82QX4oPPHMiFP6bNuuVh
5B4K1fRcmIhOnj2XXaS1LYuzU1ihKcTE4EGUEk0xfdASGqjDPPhkFGoic7zQiBOO
qnnBejhsz9InZctgXTaKoTIejxkVIJgGdKhOKjQ4N4+aVr8hAieo4kbxcH+e3Wwt
5c91cDbtqltO/28PpcZbV7ueTH3aZa/+dJ3A+YzAVQ0HhcCvWt3W1PXFZIyaDsKW
ZVltwpn3MHe0MmMj98hKdUj6cpzaMe7f0XhzpcdYKxwk1rE9p7JR4z2xZaobHeQ3
PI4AHnsXIMOsBn05e+gbaHtOWgppVS6p1jQTlQbrvfGmNyFvzc33vakDiq5UIcY3
9Hz8NNpKF3ZI1SaDymhj5JC4DYx+FNWa6/xOlTsNS94KUwxCGdeCQ6XCXoDVbBQU
XxBdJM3h/J8lEY7I/OEudJVmx0Hgal6/zeZG73ywXf+BJt80JpLxfdhQOArXtlLE
xnDzHz/nVLQdksjGdnAwGml4uGX6DicojXv+x57Emvm5y+UBxDhmvBva+6k/B/a3
Ka46OuiOkRmXx09TbwqidAJfMt1bwLiiVWCc7ENBd3O/iaEUZFvZWIybcvEs3w+I
nUxXcrHNsiG92aP4n5WmYZM3JUoXwAXF2nNcoYmkyz9WopMW8MBN0A3Vbgrh7O12
qNnII8d4ewfjWLJgVURR1ljlpjm5AnOxUsyNjMoqxxELJAvzGQuCmTsXU1E1h9CG
SEh3qWch4h79Fk3GKrY7WU8UQzlydPfT2W2ykQJ9LtA/vMddD096K0xPRLRREYpu
xRnRl53aHbgs/+36utWcJQUpQjRsrNOgRDeXkGjkbuB2c/9uaZBbaTvjQVtzgFap
j7RdRDV2n0CJ/G2H2kqChnpT+cb6/hgaqpz8DEzk7y37tixsywXHLG4x9lOSJtdw
30Vja6n0wFnQ+4luOcLqIeLeYA4g2NY/eOlO5nTHBYYkWsMLAFSpERdE3uriDHbm
I6NfyBj4exPgZg6EZgiG/EtMeOJSSz/MPvFRR0k6o1fkIdJlOvc1siuvXUeSWrii
OWPGmL62TPCmrfjF0E430w==
`protect END_PROTECTED
