`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iaiz9eKnuRSND0ZQNIXdxIyf+WyVHJqQ4Tcjy4eNB+NfuDsfPEd5szfQS4oB41HS
i2eYz/IrOhVa3HOvzEhyL/brwnnNvQBE+NVzxsp+R/Sx5GlZ6MA+388dLzQxbHH7
2e5KWAhDg4AetoXoNrrU/5V4NlGa5FxIMHGrfxZpkhNo6lu+9ElEr8NTdJibPe4C
o32GYKr5IR1t/TUEFOGnlIWwzwhlSNXeZxlZotlS+y7ZdCSQSki8ek28JGEHPRJo
z1vEJg7FlbhOvXGN6pAwu59TXmdbm02I6OY6zB0SSPDj/urqkB9o7LRVsQsuZaNr
Y6oaHCM1rVw57N+mrnZdnoMNFYIgmUNQL6UQKAptLXJMtXZhDJ0tzT2tL6i94h12
ql0+13uBOGoW9t4Hx5zJ/Pq7Cvqwv2JqQvQY6VSNoyoplEcwliU8ea5XyAWA7Dsf
BKxGa2mZrCoGsv+T54J9eUyyz8/iM/mBOGCGMfv13Ow=
`protect END_PROTECTED
