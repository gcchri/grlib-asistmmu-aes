`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L6j45WDKtS9gdtqlqCezgGBHD6uyg+tv76v9te6P5V1vtrNcOePaHCsi1N94a3pf
Xi8mRcnak7jPSOkbL2Ui0hw4uJKW0YEA7usLN+56xiLNt4rXobggOLGJ6tF6ihF5
81xpRjorkLOv1EXhiWrkD03FXDXkMp4agSnOOp5LB32iIGlkGfNiLpxmoGGMfYiT
rE/ybqC6AwdezuwDTMy6AlVvL6m5TVSV11pt9ky3WQ5mJTdDNkndnR/lrSvfxl3i
6HtYvjjKrSIsohX/Qt7qcN+9JcvTQYKRHkE0bT38A6/NU9Xie2m0+EbMbePbWjOR
zGWZfIIKqzBnYfCAigKTxC+TdJccilwjcAXz6ya3c2v4TzNZF6+KRhDIpTYkLmA6
/N9vKdvmSB4BNF54K9Lav5PkF0xX8iZTZcTJxRwMW+8/5LIt/ycVLXqWse1Xe2R9
TVikuj7J1ZF3OYW5YV6x7R2OeGEAh//OLdd4hcg+KoP4O2FKosGOaNV6O1ibL7bw
KSiANkEg/KM9rY1bjua6MUi5LwyFmf2d/zmiFhXDx86ecsi+ttGlhUTb69L9FtMs
6TYcLSORh+nhG5tSgVtgDNw2n4ZZK1m8akLtxnm18u2Yjl+fFAH1Y3lIpmyOLjKh
QHxEJcv0chSKoehCfrYECeejyk4qVKefgbqK20jTCMxrFZHX+IufDHyURBYFgUMf
44E9XD/mSN3/ZPe6g1MblbOlZWpThpGLkUIzAZpmZFA=
`protect END_PROTECTED
