`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2MHvNtLowlWaGvGyjV5WVZTGulKgRhgA7I/xqlqBvJZjVTnEeIB8zJyUdFl8IbLN
rkhpCWZStm55m6mx7NJyUcE74vBj+W1PeGxY8W7h5CwJiIxr3Zo1MdqE3xLmKeFS
oEnGyNZrq9/B6I6FqsTZsJAmxGlyQcXFKXfvp/U4gTWFINyGg0zBkewIap7Q2Uab
yns3nZeYVRrAAF5heg7F2PT7ewxIjND+oijUOYX8fUHG+h7LyNkChCSXxQ1kdWWx
U6TbY3k+uzkREu2zFi97j9RDGk3LYsgYs3NcyIaD7VJY30DFSWV+44CBMz0JIGLp
Q2dThvmRSbwYLUiTy/jM9KGsVr+mjwXmCJ2QdIBwjSkA8r7UnTiwTQQfkWEoa5QQ
PcKCxbNnHYX0YEhP1ZMgoYW5ddGHYztNWSi/6YT435FV1R/PdQNprHFQ5uz59k9D
QT/hbGUNB2306RHvkYGYUq9rJpvsLUmxC7RmrtVs1U/ypYQAMK/Pp+3dRAoNQo2l
L3epZogxNbbEQ8P97oHA/PFrfG/JXw6sCgk0K53/nIRkMS+tK6YI7S3B9CpSxeKC
c5pUZuNa4zTOcEJI0toEYwWrKIjZmpV7ne0lKW1gtBsyNuOUVxrEgXSiBxwiPHtz
fqQN6sla7uPRXfSgiwEIh+eR68xjq0Zh25I0LlBH1Ez0Fp56iQhwO+2YK7g2K5+x
/gVcrLPidP4ndWRt/0pogyCnbwagxiTz4Ws/Nx6kvnOMeLIahIMbAC01IhX30YFZ
TncdWM/by9YAAqFu6wK5DQ==
`protect END_PROTECTED
