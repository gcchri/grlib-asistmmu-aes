`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JwLKEt/jMpQQjteltXhOFCUhGQzJAC89AX3fCaEz3rLcRhTqGmGMYvSVx515OMYI
XZVY5X9SoRmdek5fyBXyHUkiNGDcgvyQFEECpgkw4Q5ZgtU+i2BXQ583x6eaBO63
MCHPLaUkeNB2DcbPWcsdCX6/6jO86Ix5lFj2hmJ31yrnpthnDcjsbX3iLxEAAj9T
q+iHSAMOUEK1Z9XhkPB6ZhVY5v1zpSAFT6zaNgR8DYI5iBUOfRPP5ErsyQYpndmg
6H5BUmyeNEJ7hB767BdbcGBCW1tIcnyGhdHcekP3qZYyPwWMkN/FwR5HgBbpQp6a
DSjQikIfScSMHJn+Pw35T6OFQzb/u9bp2+9j1QthW1X/vmeIL3O/iqgYUy/Aqkk4
uC/G1psGQeTEo/AkY9kvMcuu2RhsnW/Gv745YXihowScGWZxYhK/A7iI4rvBKJsJ
xA1lwhyQqYIdZvCGSN/sqqIe6Z6icBBHOP+1IjZI3tNhjqz4pUywfxC7egQewlF5
dhUCbREZIrCPzFbT1355O9j3BuqM34XPdQWuFKfV0d5ybMno89WoQ81UyiTNttrJ
g4ki/B4y0dPn5xji1bXWQ38/9dnFt163uztR5KKwpM0UMHA9dfhB1nG943Wi+zm5
pumNuG8oI+zzLnlTvuYlZA==
`protect END_PROTECTED
