`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tKXaKdWG4qU9ScrOiGM+nVbPXsRY+KzkIOcpVNs9ErWnTojdKVMcEYStkP9/MLoQ
kYXqMjq7jja4GPGrxXjR8sXzHxuBYVYGtM7H50xkrDh+DzFsxpN1Gq0hWb2IZW80
Flx/2jwiCdtP7QH5tV7B10eiSLJXrcAStIHAch3ZZHYQbRLC+2w3tBDHtJWfRcqC
ZmDDi5bsFAZJMa/kotnfpyf8BfKw74Fz5jrU/bXwTaU4XecmjsaqGGCJxmbCFnFP
1Ra0KkKHXWiY07Y4qVIecaWInwUPUUSiFIzkSdtbE1kV8o2lYkid0f2GkPIg/Sk2
srui3AVqIkewUFRfkOytIwHkDgxTLLFH0Wv/IxXPf2BcykqqglruXxThdxWb+PTp
2tjId+rF5wpXFN0QwN4aRkPHxTVQ6XJwx0bvl4irUU/A9Qlz6aTRq7TaC0H5XxfI
Jitv07jmDBo9AY8ZnOnWUSJDWjyGZZFrU/JjsFvq2dynZO+te7vEdHoATM7x/tz5
gjw+2IeJ1CLIGpbhQaN4/pLLmJ0aj0birWehejc5LVJ81g6igu8MPcRzva278LBU
fq1AsID2oDdOeO//JSmMsASsRtErdBTLqV8MXdF0yni0mjR6TD0cQi9pSiEVkipu
YVLGepkkOqYxO3XJYK6eB+7UMXuDAylv8FFRTQ1U3vMNv325udi7JxSOc0AeSI+b
DImk2lbUBuYzmlltyn93ETk0/4KkE+7+foeNiKPWKFpFzMkYpAzeNAC9AfR8TMH9
59f2QvpFd0cicMkGCopFwISp+7mUm+uxhGewk131Qu3TaxIjQcsrbVbwx2qC9iCs
0R05TU/S/ueUcEjSYQuadVhb/k2bs16uMwNfrWgMWvPvqOcoDoXKdIvpUZQnajFN
FZ9mZoZHzofex42hCVGUsOxZrMrTRq1lWh8IpGkKLGNgKP9t+n/86x1W0mPUyXuo
zPJESWF3HvfU2sbBHAA1F6fSzP6hRWpTwJTKU9xjauIN4eMy3TpvGXEOdpKQBeoF
aXKrhGrXGQcbWVZMpWDackLs7c4DyZhL16bxk+afXsRqdZr+F9/v7vJQu7kiZXZm
TN9hEN82/IaUZ5phYmzkbgdZ5Cr0zlR7atWKYvYHJdhkXRfzhcDsYzcalvj88zEs
2jVpnU4qjd/NiiijTBE+eeC1pphNuo761E2I4jAbyVv9E9u+bMrPMtOMXEezEsao
L8MnPJlYzw0Y/kYCD5jb2egSl9VkoEcUM/1ioQbViSIT7s7MKj4Arxpr3mMX9E5c
cwEVBrT+xrSGVuIc/3598CQIx67Cde7ai28jeMbjDLAGChNcBXn0EGIeiX2E7ImL
GklxKyZ6u/5s3hpnqC4I+BQZ+U7RhSDOXsTo1gKOIa2R7OxX1oiuE3+7/1xU/w3L
9vig/0QomNdDR0jBOSRexA==
`protect END_PROTECTED
