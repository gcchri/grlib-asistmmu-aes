`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UZ9rzJdZ98zycIC94Zs5H+MFdneMsyjTBb9ou7j1bNzdnproP4Yqp36hcBETL0RZ
/Zc5xWcYfQLru8X4d1fw+M+qdANL0qF0Awf+nzJJNThi4ntxGy7RkrA2cvl1eILM
gL7tkZ3kYPpZrHN3w65uK0HzPA3EZmIDo26ISPLIEAZ3xtLoIyjyxOzbFWXz3ezn
J4fdRI30UZTok66HXnxjT1KcIvK/wemKVviLUT662fk4DCJNmsDET/0B7vzoV9qN
ZrL+860UhOVABrlk693Gn2DynOXT2xMcod1khH3mUhD9V61oAy/DvFJWhoetF9Sb
gKMW3T6EtuqOi9q0mxSndqdAfMMP/z4fqlQlXzgE/r5Gk0enfTZWFQmy+tyxUuQU
HuXJQRnFcEkBxLUWSTSzTSG3/2BdcauWg4dwEzPX0201lIzzB2RL+/uYhG0BX/gc
ALt8c7kwQQ9DkG5bKe/2wAcPbibqkvJXPvi2bb1pcGdh3/2+th9IX5q4HHLyarcF
zXwPiYHhKvykFYnXkYjrbZvS+SCGj3LSN9+eBBF0QwQvK1QAzsKarn40Go6FDVg9
uRP4hqX4qxSAOBgdZUYXShxTlTWjzI3sd604H0MlGno7nAxtqZVUtgjFFh49DXGx
z2JGQl4mcrbdUsc6kR9mOgW/dArXHKz82xa1eoAcSPecsRCC0ogSX6sy617aeZ66
`protect END_PROTECTED
