`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rt2rY3eL1KadrQHrR2Xv9OJ9C1vH7d9U9f2rw4muWI91TgHxHpXOEWlGU9+MDMdp
fkO6FnSAbF1lJbxM8TeaWQaZF1VcwGostw0k9umq+n84GN783I9lKkNe4Dn6aJt6
faSVasT+f3fjhJ/qeZzL7E0SKinpXv5aWLgJhq5lCv+HAV32b1bzgWS/5eF363EJ
eZG1Dfnj1Eu0/cqsujKcNAimsPq+0swPM7EGgrIuvQEtqPM+A9UONsvNmFsyWYNk
nNPYt0rYq2sNBGU5YNT36rr8b+6Iku5fJSLhwPaXtckBuEAIu9OMktPlIHHe9A6s
h9WZn3unCZev/W/oDp3t9lHBCzmQdRqoXEMeTrefNpPpcr8RDABtcKLG4+DJBBLU
ruqmvqWPakINQMV4/JCBcJtS26gI3fTcfShZcpnOflFxx5Z61Y1UpKFz3TATCBGW
TIXMKnOkQIJXwD9DuUB1F4zoTLGzKcUP8UnvlPtZn+hd4vRP6+fs/CGDyh7j+7mY
lCnetTnp1Y/NyGlywSaSPD7x/vbao1z88P7WJe7jtwfKGVUglyoxLazgO4NjH1Yf
FkgIuEW398nxJm6oePoNcLsxgMpPKBIl267Kl91/t2I=
`protect END_PROTECTED
