`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HD0YzttS053EiIhthf9RdeePSD7cDYlzOs5J0caFfYFL8KXSqSr36EH6AT3aDBNS
hNeh4STylIm5IELMk9gHnTTw7LBtuKA3FRI+UB9ih6FKHRCNCbx9vLpaP0jdRXGH
EYpa4eubfEfsnhsa84RmUEMVYQPzH0BMehbD+Jj42SroT+fErEgQSZBRR25zh9VE
E8IGNKUnaOGJEmj5LmO2K6yUCIGNjauypHTBqQvTsuIpJwsZck9AnjuRL5D8c4av
ViR1CyTD4LOtKjEvow+X1hEG1CnqNrKx3x/oM2BWN79NmOrVn0vRte2iX4g4knrS
wJ0tB+VC0pxfOu6W2F/xXVdj/wh5gqfLdN+CTbV3mUOtnwvZ8TTEJMCI07yK+8Ki
zQxqA2g1cy4V9Fw7RNyknhcmklFa8iYgjPSiReZ5yheDaRCIvbosx++cIPvzhEY3
hWZAxxtEU6vDz5717OcthVmqZYdAWW9BC2bf7hWGqTM2J4SeiWCa0D1VdYgNmdpj
L9fxNKIJhtKaby2eFziw6USsc+OiQ8cepOgfp3HvJfPRnbACTva+OJtJBPT5Ja7Y
RCLhZWXNzS1bvaS9EbnlfU9h/slZ5Frt9Fvd+emLrICUaIgq1P1PJWCmt6mCyA9/
PW3V6+4NTZZoAr2utbspLaCo0RnCaWptkT6LCLuR0f29TTb+CMY86V1IxF8/nQcq
l8+9xHgbQlh59/7xAmtYL8tiutIbPfCGKP5+VlwlPFqp4nnbXrEMYvFFl8ZwKM1T
`protect END_PROTECTED
