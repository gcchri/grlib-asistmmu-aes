`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fPpNST2LItTIjyx5aHeNpQEb/yvOrcjQR7SyessZmI5nnGTpNeVgn6cOTn9uqN9Q
58oCaEfWfa7RnncD04uHOIHHxXBu3gljX/dwYFCRMIGBuzwelkqIthLZm+NKd8Eb
KmsuC+DtNgzCNR9WSTmsO9+G2jVEIoTnhHiU+mCG64b6fH0a7nHyJieTnJZ3s9Tm
185DG7ylnhiFH/vT4OjoPWLtSybAqnLpaj3LMGBHHxWVzA0in5DtwwM6yw+psUyh
QBnIrGwmAzXRvZtdYzB3Lna4YV8dg9sP/ITGRLlhy5efWmyaYJ7wB+0SQ8i7FIqJ
4KrV2X1n+yj9dGvQM8FZJr3sGGfq/9htlRNqW+a8N1wLsoCed/RWsu6nMsD9W68d
`protect END_PROTECTED
