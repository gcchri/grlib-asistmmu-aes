`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NaQ6q/LKVSyk1RSf5cEcg4c9qOVaUiNkB3WXk/UabeJyMkJvXvucxhxaiZPSVIHr
WH1I36UUE42CCaJkbBRbWa1cWM9UfBTC0oPT4bl+4c+XB9zL53LvkZF0hxemnQr/
XSBJLQuZoH7+QzRL1iEWJl1BcHdasVC9Q5eTRFfBXQZafnHy8sh/h46aM2RvmVqN
bqKNmEwfF92pygKM5uxRx902JIUY4zBnZ0cGVcl681gbNlTLfDOXCWmPcvxY+rmZ
+M7JPnq78m2Hb/0763D+yOamfAJF4TkyyCsmaBfv6by4p676DsV3itQdRTAsQSJG
UAJUb9u83QrcZD3qxXQS5mu7agSI/3u/MsYHhcr4QvfaGF2PrHIhBU1xYnADMEJs
IYd08z/fRxCKTEJSutwO5Q46ucwjh64v6GUe9/0+1g8rbJJJLacfl7sliHo6/YBa
jfGCCnynTlVY2vKSAP2HECxIWonx0drMUifpTobfwCHbuvCBKWv7a32gQnQIj6DU
`protect END_PROTECTED
