`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VU2KEUBM4CPX41whvwKBBkmKRibX8KESYuIoLLBMmA4m0Qv7Z+gH5FKZPRpeZ2Uk
K38m8MTgFuhLsx65EYogDqylmIILMNMsArqfY9SQ5KaYeWYOo1bap7iepudyjBcu
UKldtiGDn1VHUxClu6hqkNWOsxWSZPfRqHTXte0Z1iJTKNm7kB+Ir9e4v2IxO7Ok
x54wQ2ILaNCN00YvZ32k7f82XIDUILYXIgaodYLN9v0i+nan4MJ52znZGpNyrbdQ
SmBIzEW1JF1jQVlCoLUToPc3VPbFtMEJgYbBsR4LdRU=
`protect END_PROTECTED
