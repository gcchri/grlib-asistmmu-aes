`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Mbn+bCouMJD7faCXVRSnBgSsc62y+eKqW408Bm8UhLGYMybLvDnFc1LNjFlVlu0
K3EVBZu2KlRmlIUuTyi8t3mki8y1YLLDJoVxRJLie+vzfcs4+/zYtuncg71xspNi
kaVWElb3HjHYTkdNRMp0Z8DZsWzoBABjNe9Og0pkCGPJaAtPBkScNW0+E/uXNHHk
uG+cVRw5Xv+m8yvAgrNgrW9/OLrVTQkA0ymT+eGnBtHzeVnY/B/kwfEAgGXxUJZD
AObC6rnCeay0lamAqolLI4Sd95Ct7xq1TxD2wdODZqQ=
`protect END_PROTECTED
