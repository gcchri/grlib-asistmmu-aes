`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xEQGZBNM22h/oQn0xD9h2+25al5Dk7X19EB0+E/nZRtCAQlHcUDlTL7q+aFJ9CND
2Qz6RLZaCsyf1rbZ9WCq4+jJR6ZuRyhzzCrDhujPGCxgaBG3XiL4uWori9W3rtQj
/jZ1LoGWKXxADMtkFBqCPizNYM97nas4px4Yr4BRQhsylnE5HCf6fehzllhvqMa7
WY5QMtZWdi94ZC4ZghO0H9BWWKfhaiA+GuqNIdF0OV/6FHUTXbKthoVwaFTQXF0X
2TEaoJgHjoK5ZP5jX1/rQruHa/s1iTu0uzGuJj6pkCAnHuPcUJh7EMPLT2xCRmd9
FVHUK9/elIvBJpX96kLjWE++BL0S1nPh0cBVX92nfYcwUEE0D/G4rJ9wS6v4apCd
75LM60b9IIIGtJjYm3E4CdWbcEYc8pD2cdDFsIcj4BLTBxL62o83530WCvgY3Txg
`protect END_PROTECTED
