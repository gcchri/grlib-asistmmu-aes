`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l64IRdBSc9tsS3E4vvDWgWUiCpKZu5OWY6K7mCIRyBmicyrjiVciAkFQ4XhcPVYZ
dKQQmJR1zNxoiem5hnnPlMJX8dfiaNLXMy4VW6zTc3sbynKXDJvIGzi/9ONelfbw
Xgu0vEZwj3Wv4NlKfsimXk4eGnqZykIm1tQykvzjEiw7RNao3q0VG3jzgKMsCtxB
OGQr9nh80evsa2sAVBZ8HT/2c20JBRqDYEvkmB3Gj4K+vlkQNgE9eDCAZZkpfFuu
6JINQzZ1sLvApUMiqoaEO6P4g80u3SlC5f239b9hpNKtI9Ln/D/qrH2JywK6hTwh
kkWtEolPLpimXGK1lDtCql4LsRm1leEKmV5BPnno3rNgBMafjclbLhMtosJy2hRA
U6jsZinuNbAMytN+blcEBMA78Diw++5Sm+NLw7yUkQtAdBChPsXe9YrC+A/DGHVz
eFpZimhADR5tnWwZqrrNKESJgDpRwfk7WWpfyYVU/EeQiiYgudIvXLCHqCvL3d85
AjLOkTrVMrl7wyjv22gpdT5QwOYSdyCAXkc+XKkOIe0xXbrHVyBZdt2IzzB7Jqsk
jgavsMz2wwmZ+Jzxa2HETQ==
`protect END_PROTECTED
