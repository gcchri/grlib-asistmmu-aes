`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iWS0fUXn8MdjpN9yc3K+2SG1lFXC6/6RNxMeWsVDiwR+VX/ZtRrERdWgDd9EQg21
7xG9Auxqf/N2Mb92VEs5aXd/+Qlc0X0oRuxAeZeDcau8EQg8AFLYbg+pP6THnVvo
3gYY2RUcgGGAO27Z9t6qopwswffb7ryKji80Kxr1wpMMV9YAnWVm33xhtN950KK0
Xe6TTlHypDFu+bGuWZtH4dbBEwlfu8Gvzs/MWcingOfMZ9ZQpDL3UEvyX+vvuuK6
W1rPyBqn8t4uik2r07SAtSLkWBBG7U3uhNMPsD+POhT+gTqxV5i5Q4aNBwdiYSc/
m/QUmnLYZhoDbcsfxgfVpIsrzI7yWj6iN2/BXfUDMFYT1H+eKEM6/sgmQ66/xlOT
GGYlH2sT/6B5sP/6OyIclG27wHZyvsig+HZL2W5RWzw=
`protect END_PROTECTED
