`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O0eF6VQraKXb52XXSt0ZV3/kGzcC6/b17QRLro51/mcJAkKwZiKi2RFT9UU41Dfw
wJo2Gaw/T87OA0NJ8lNA8t7DfSBHxLV6byWJGhdFPfI/vBoljzElTNho74I/ZL+j
uw3s58Vro/Ozenhwry6mZvgnlYLER2UrkYrZbFWAjGOSDwaY7pGch6ebqVncUQih
jZwSUT+bv+C6SlBkPs0NTa/gRPwTdGUV7VvIpX9WFqAAo+FKGxILDMRmyYiIErNN
eN6qoWJZSNlKNzJ+c6JoM0lAXhN/2yDPJmupr9CWYo84do5ssP+36bWsoafmb1Ub
h9/ROk4TdvYa/twNYBHdMLVNkC9WwiGGD45IOLMxC0uSOqwAv8/1WNYqsaUzcXKq
NGHOB2kg/Erpgx4RMPjeut1uSI+vXVdVVoc5kAo+0c2dsDDNeWDvIVw29+jkJzrL
1P6VeUDGJygxfBpTAB+J/JpLhnnjDckXoxGrnSCPCdSBus0GGq2PwvzFIAjtp59d
IHvWIu4frQ3f1UfAFXgbodu+kHprhHKxUwY5O8GSORoi634FH3ufv/Gz5JE6hYdj
3k6m5NtbRVbx/E6jCFcLDsrO5lt0UPeRNaY1hOiTWm9EYs8m2h5wVqIGCxrk7+eb
iNfxwRzlkuIxefr2SkGKvQ72fXhs+hWUQkK1L/GGHNGwxuW/ZtH1VaXHZiYRi9aF
j2eUs/aDXNqHu2A4KlN1jhQYWo6mO3bUJ2eIDzBH4osWCI6JLhEfb1L78ZbvCYVt
CBlE6Xfc85SMXjyDxpWT62GDenMCdd+qJxVADkxjP0k28YXYqlgHVGdFu3qNGEDr
zfBOsmkHAy5SvODx5t3klm8fM1JiAIw14sgqAJf62XodM28kJC+FMHMfPRjj1yGC
tN6vWBkQoMhT1lvCJH3vp0p9pgHIqLAG+t9Qyn9/Gz4T1JQSvfySuEmLf8lk/+Vc
m7wcPOdoT4ErWETIliQlV7Xyd5engakj/x9eaW4hbB4=
`protect END_PROTECTED
