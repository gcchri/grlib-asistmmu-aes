`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ni5JDqq+V+in8IFvLpuQPBGFekW+i6Tmw0Q++alGqKtVcgFx6E+zO95OyN+2kbiP
Lsn4qudUYR2cZBY2mcFDn7iHWLi8ZYSjWIpktPaJ6qjv9BkNYx3FgVvjQkf06GV/
oT8jhY+g4JTzOI79uQjPxp1bEWpYRTqaZN6CY3NVViVvlcsEwZIHtXv4mXd2pXxC
oPcDSfOWbTr+UuaOAdlO9LM6/+BgwAD0OnVhnrB7U0Vq4RxvIHJWqwD7zbELaRo9
bM02UEHOpDKUyLKJ8v9ia9O3/3q2J3WwkPdU42i0nEpSGByjn1Ls/jj0V3dQT0Gk
ShLpxyKZl/GliUxgH/rgRgRQPgF5UgiPxtTOvJj2zUolAAOHU/ve+nLwg+o3GqQT
gtwWJst83cHhWhu8Jp8JprjPgCJSrgiD7CH0ApEFK61z5O8CIVjuSsDeCArpGvz8
D/9Ss71ufldY8zpabToWdUhVtW7pzae2mwhyQzGZCvrPeNQ4RB66a+56Za6VgTXN
8bitR0vo1VlRrKPFoc3+4WfCtQJ9zrIvbJeGe71EsPAVFvRYVKVJ652G8eGRSXrH
gxRi6hgI7FKiC6CoTlB3JWmcFYpTmeKQL0kWZ6Tc60m+Ax1VtrrBIbIC/hS8MEoj
j8rBhwWoOQkUo26ma4ZjARJqXnGiF0qu2zVyou0H3NYnGS/lmANTxfAIYaDeCGHz
ll7FsduA97334VlKIatSKQ9AUmANN+Tpql0sSibgQuMJZupYu92/MJCw1D428H2d
mMkjJLhDf6kk+0hecF4zNsjUcbjBRj4Uo32ZOYkqCVgCfHR3w7O0fVosJenpCgHs
r/oDZkkLbIMS5yHrrnkJhiuwXEp3uuP39zuDzBjOsdiwLV3CAStD39IQoUK7Foem
GrwU6keL49r+r0jYlK0KCL8PeQe7gGrIJCPahJw7cYe1tkwDZT9ALJPouTMK6voi
FIFVD0IYI3ClGlzsxVCp2ivCOLSVU+B2AvPy2R1CWBrg/TghhbRMJHHJ+3eNbLYD
9OwDU0zbzNCR1+Sxv02y71gOwQryxc7UZZlMdVcs+RgktE2zxa7336YzqDoMr3Ed
yyfHouC8bxAS/oS6wAqmNkAyde7l5EUMiDtcXMX6bCdB5Q+hNJ4r3ZOxAk6FGCNg
Pl5upkC4koOHvis7zrgN/iHg/9j2JY/pVN48dP+P3de/8pq98QvxT7VooShV5Jd/
WF0s47mj1poDrOpxK1qf6WUNudAMicl3hWaBlZiHxSBQ/4LE0JGQTfhnEw/0Kcfm
BJNCbuRM2tViLkYlM+Zc/A0QGwLxg5VnWX3OH5vY7VfaSPoHpEUvDZ0L42BNhnjJ
RPkevuKS3GSV3C9yFl1zXEIm+AKIlC75nDXBgtJJ25twQDALl7kuy6DiWnqHRw6q
U1aueAeew/fdhs8caGjHAmaHEOWMcBjxebRwhZHflf4dGBDU4aBY+WMqjgzFphYU
SXDwxVG2A72m1QvgMbo2pF/MN65Kku7TXXsZ4IXYNPBbILS+WPpnBivwMRwZvm7F
RGaSWguDsQIUSpoYbAdTdz+evZKNOzzQUORo1skWdc1G+nHtHVZ0b0sduAj/TG6A
ecgf9QQ5HbCTpPQoSGi52HMfKPhfs150eXTYI8DF2WK1w2v/Pc80+JgMxU3Ex2Iq
XMZ13t4kXoDjXWQRgitlRdxwB82uYfL+jguZCe3QjppywdIeGl2DQQPOKOYbJ3WR
YwCzAMFHiTgtZUK1IwluoyUMdbQbDKpco5xylgivnnYQjt5JuaNxpVRUEM9ShZbF
0H0N4yvk9HoqL+KWI8o7MEv7AxdmaD0D2HYTXZS3XNvEoyXfncvom2PJ59DiyBVs
mc4VdkSwwHRhZ5uSKO70S0HwTXJQrZvktSETBDUAVtTjWPUZ3OdO704tXeEgXb++
pB5btAJ1tBRIFEpzcGsoXUz8f+qfw8eUpWYVAJaN40SuqBORj60SKF0haYSbMEJF
eSSpDr8pDIECHaigY32psrj5kkC2+KlmrMCa3nZNthKKji+RpD4QCBu3klynN/tI
34FT0rGIYi98K0nNByPt9cip1x4f2UilZnR0BwkDATew3WbqAk394w4XBfhnM5be
MDjuZIiAw92SzraVkdE3LJUCFmNIcdf1oREp3+OUL7dINJah82dXfWoGOm4va39V
7q1bsBkoIY9lnfDDy5WK5NLfpXwlEL5p1MkKsFwu7Zo5DBMC1ZwUq11Myd2CYU9D
v6QwPGgeu+k+5qJwtMO09QgrD6mDddhMrYYRrTbsSaKGWbwnxGh0cigkXIKOAmY1
YJZfyR4oBzqIe117SU0I8tRc23KoVvDE8Ty9kb9+G0ks/rJr7oDQKc1rzlkOLigO
h3pQxyzFfllt934gfLw/N7XharJfHSOJT8mc3MIp6+2KXRqVtyjBiH1rrqRBIqEB
fl5JcZ927m9OIhSffusWbFbtMcuAlXnaPW1qAOr7c4MHJw6phfqdvMLcohLjLmO2
HbgIcGt+WM5V+mhP0pRCJPytf3q20bFrXKbQoLB2TntXbmZZ1clc9YtIkurXiwDZ
TGyzr5wTdT8hLPkuJwPJhNWRb6pYuM0x+6RvWjmoIBzVsLGsjSz5xy8DAiYPQAhO
SPAo+Cf6v+PQdY3maDwtKHYaQs8CaL7BnhcgENeNmKZB/esNaz+ymn65QivNrSbO
Kl32wSJ+ZncfIypoSA3+L+SMK7r+pUB1/4PrNOx94FOh+oHntqcgJOa8XaxlWzPi
B2uUVCiCydGedOHVQqIX/HdveGAxYdfGZISnPM6Mwgn+jsPxtYfyW210+ZXv3B/Z
giVwYsWtBp5A1K84XxK/CZltzKeCXKlYQsLvfGAmSSdrgYEneoeOxk0QDWzGKkQz
BXC+2ZRFVhjlrsCB2+aeA1Zn9gAbjFo0uJr5YHgTVdD3E0VSWIitC6hdo5EkGi7/
BQlTMF88NUDEhLf8vOyxhw==
`protect END_PROTECTED
