`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uSLwA+PXiCSfjaGQm+rf6/qD2DDRN4k6sO+c4oqlTwX8tLQMj4bE2lSVxV3iC6pD
wlftm2tepqPDr5OJvkQqq7jloeOybSKT9q3K61O/m8c3n+D50CxCXBYi+oKS3uS5
/B2fRV7dPaHqijSeb+K8fry5tEsq3UzZpbkU+UxaruX+4svMIwuVd16xi3PRUhpE
WnUCdty+jj9BsXJMdLRoFlW9bbofio5Ua8B8bsqe/BG6rra9VwUwltY9cJKiFkoI
EhmeE7257liBFvnOb0Blag==
`protect END_PROTECTED
