`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M+VmV43A7MWhuyPvQ1JBLpQRtmaQS2RfMndorr8iEm7upHx2XyWbpAfSdVc3t3kf
Foby7wU4t7hOakeZQbxVlXAKoz/2Dyxgm7ZQ32JWYkLhvFa5QeFi/D4c89gdOSOq
Xj+EZ3GNCS0iYva86D2HRREMR3Q0e2vVmQMrWAASG/Aa20CxlMF4melYnJ4WlKod
jnlq62ew0crZ+gbBQwp/315bNDZhwkNbjRaOXzxJWWbkkJ3yxVRUfpjUBKoCVXMW
Vk17+N8aeICwTYfdRGWSUqZqGgv9ay9mdrrHv349RrQ4CZeR6k5c0Ue2Qy/yqV8+
Lm+eAdMk9XvSvpnK9Naqtu60L5akkByraqlNQxBYbEMwoGvM2j4o/59ox/6Q7BkG
QMHI/uNjsPmveujrX0ufguYb+MUMUPI8Tqy6tG0E9Ng9fUIpfz77B56huvo+v1r4
l4Ef20RQzG63OyEQtc2luHXpdClh4/zqVSA7C1bGEBnyEDSJg8EC6I4EYvRDB8IS
QVlx4vGuh3a/7RtbK2+mbAWt0KI3htHA+0fqG5AaJLCd6+hG9e6IYTuH0vjdOml7
xmsqcQEwfCwM1lnQhztC2fJ0ll4fmv+MGtpv7CVWSoRUCCBqK6vHILkJmaZayZuE
l1LyE8cBGva+HCX7+Cth04MgzSinn+g6serl2helJJIxBruCDjgErQj3n3rsjoKu
XbAcAewTv7lbc2nhKr1ZskH7a0bH+VIMD+QH72b+D9s6y6qg/fcNeCfRDFg+BGBB
M/++ViXpkLgwwlQmffShoVDf//kO9v+8tJCqjcAM78nbyuc4vw8oK+I0Cjp5yY+r
5zAHJQERzrakXksK/iSbMlXSnvCB3vAlPKcUIZTCMHt6iYMlQCkJyMNlHmQNQYAs
jbcE6xCfrybb4O4O/hntvcRgn1K125cTOf4TNknGS8D4qUJZw1Sl5eFs5z2vm3jg
2FPdSJ3mm87ZA/D9Dgx8Lakp2tg4Qowflxg2EZ3ZLqMEOqhFvfsuO4/K0D18ugx3
EozlnxEittawilpC4sjvxcgWMClVnc0PvW6MMaL/3e6rlBjitgU4HzPYL0KU6UnO
sQ7X6hJlWrg+GqhndfeDzvV9tm9qb8J+/Oqxwsmz2otzhihRAjFJICmKkIqh708H
pwlfQtj7paaRjpUuj6hQTH6YBOM3nix6BpL7XCP3yBRVSXMXZIvaiC92o4YEkQH9
UmVCGKGCbOnCMcC2gc3AdzCmT7LFjDuUY2g/w1cA63A+epxQ4rJFoc1mW6sUd3tw
/IBLOGArLHKR1w5ARhl25uIPyJ58XHXd10zPMvFrOHMh7yk0kp28+p2UU58nVNDM
ETr7ttdJ0UgdtKhS7HWbFJr1APYR2u8YY8tfEs6oP4qHiFXm9E6/UgXO7EhYrKOQ
6GDwv0mALEGAPlErK6KfSiaXtNl29EEjPbgnAMULektSYf3mJZL6yyZ5QFROJmNm
CG9/j5yGOPTmfqGRbZrbkzHfuyFeXc8ioWZAGgwQYISdmBIr15X8KNaZ6zOBl8mK
eAmn2jv/X6HFouGiksy9ATGafBPl7LbKIw5kTN0XMuOvHRfTjVCShm5KBeOwn4MY
Y8sY2tA2FUMmhqQ8TkF3LUVprWYsGhGupaOK8jwZ4MGEng7eZAk3rRBO/dC20Vsm
9UPu9s2FR0lMgetH2zsmbcpFVKEqKmmpnDuVaA4Ow3o2Ci+L287XMgWgcwTpjwGA
3ljcP9cuYza97P5Evkg9QNHj3K32ur+iBc3EAgH84ePf+KWnacqm6LIQrGnkcui8
lwnEvbq2kASlhH8np5khryIYC0+i8Ozb1X8sYxRwdOhvmhE+F9h6OrX1GUI0uD1z
p8+e5v7UAWOcExfp3E4AZobMvnlfKZKLV7vGC4Md8vVjAIGbolyicT/FtlY67ed2
JpfXunwUKqyFRRATx1YgSxXDKXPWc591darhMmM8hhqvMER+VBAUd/UOyaPsancr
xIvfEwYoB12LMh2lovWk/bHDiEhsI1W0XvTnsqD98PD6MWq/7BagVUdTtg+U1Z8h
E6xEx0T+KkuoH2mvtj0tCnEp8QalcTDU0qjQA9b8T1mnOFRBVP5kN4VQXJWV+uuz
XOZf7qOSIBL+9XTBVKiOfY7rG7vfmCK+w7b3qTX/XG0zwsrFmqAtuTHWEuYIxj5l
lo9oqkufC5ZiGhO/RM6KHtH0WjonCTGZ0HtdJ3KkHJbP0E5N0LN5rPMTkoXsTqfd
Yn9N+NJhJhUqqPIbRbt/zPIdya5O5P/R0juDGmsNluH561gT90Bh6cjXaxWqtNvT
noHpEUZROHadWWKX27IHGVx0ukLUOA5cmiVFKkwcL5vKG/2K68RSErTSqvBVDueH
SXoORqA7WHi/4qpOcZwY356qf7IKMDCEx03dL07kA1xta7qDEkycKXGYpWA7WhFi
I3HV9YQcPXbdS183xC7TjNE/jalyksSUhmLxaAx055xlq/SIfXwhJQEd5nZDHMZW
ejzfloWuuiMbpSoyXM8j7CaSbmrdCAsWeaC++/+2/j0xzfXT+eohmUhEvtA/5arT
QWWwdURzZ9VPVm72Gjg3xqZoqSpOmxg6V7Pf30Nv5iT6lZNOWHBwM84ErZBs+Czw
nqjDhyOyK64IqHlIixec1Rr6nrBTvzxaYzX9QW4uD1yIL5ezaHfoDeCHRcOPqAeP
RGPdwC8cHqZeW0Mi6PT87mWOi0O4H9KGQGhbUY8QpugLsa1xF/Pq3/MTmGnCmRW/
de03csaxYD3BR1evoyKCAuo5JegfV1jksky1fDT9Q7yzq8lrvzFes1mYPOSUGP35
7gi9ihvrwcvpCQdBYf1mhCr9kWBmW7WdC9PpJhWAYK3ZYzS3Xf0aJZR/z+ZOdfs9
mJAw6OY+kBPSaVyj1JlekjzltaOaYQkS22edcIBBt6wfXeDQiE78i7lnSw1gMHi1
hrFMraeTG89XgfC4GaUZ62KLc2hN0CSuIscdgiE8hJiPk+flaTMuJhdWTC2ANCP5
QrVSflED/Sd94FZ4Rx5nyQoSTLAEvXDzsqsah9CkFsIlYsYSV9P2y+ZMCiQmpVWR
a2EMjlHDlsYiIQ48CF/grVsPsjOYX0EipRoXiO6xSTAZ3JiMQzH/BHjp4OCowoJx
gs+m5x8ue/iShdpIDbXtrqKswxoPYSZgKUWi0daOMvKQbDkdNTbunboy2lL7CB3N
UBuP9hjCHq0gQBrce/abxNT5dl5F7P75ypGzThPy/vJ+KrxTwuqLzsDLdj6fvSNU
W3cHdrsoIZ4Tq97m/r53eSd5DALgHB9mp/eJoCivDw+u0GCFE5HDNd8gaMUbEyzD
LD8od1Huo2gNVfN7Ih9cPuS+KcESwpgdvd6rygOd9xNu01GNBTQfy/ErQPtlLqi2
NVUbv3VgOG+sma+qv3omSBg1QUcsj4kJYj2lIEdU2aAHmhHjCyzD9QdtrIFtWLEl
NTStdLRsIfFmMjw99GxB1WaQC7XvBPr3ISAZu76wXg5J0keO/Qm7MIXsvT+VhwZ6
/RdyZQQikzi3gMpwtpIwwvTJWOoCEfv9iNO2fe18T9lU6ZiplzWlqInywJkoyE18
Lic/WDSrMQ3Kfj5hgsBz6buXkiuH1ZEf2NBQWYz3j5SHvcPkrK+mxiWu7anbPxQH
+zm1/QZLxQHc3hE5VCqSiv3HcBhUB/cxn+TfTF0UQaGg5UXFKpYilEvndZIIYxmY
VOM5TfZpXqoKHfMgCMEuRujWayT3D/9fa1tWVEmpN6DRh4PVhb4J4jRaLFqmZ0i8
s1ENLhAEkfVtlPVMJfF8fN60bEKdtvwquWoHBhCcNUljMbdUTIFfDdHU0xDrE2RG
DrFhio74jwxEKhtZFJfhpyXgDh7AXI3mY6ej7FCKcQVjMBY9w2Nf1sKcIIe8iqGf
CpMPCiZI+ffnQmGKUgKPmKTvUlyxSZKEm84okGZeDjtbTB7Srn0kXZN52P8jfUdD
E3UXSk9EEWlgA6sJk2P+myhzGmbn4K75Lj9MtT+z5wnXHQe0kZgj1I8HA/ALIZXP
hQ0zVTMzq9SixWdbsuZrp2p5JGKUVAVTCZFDGyBJSHPrk3MiycsERIIT4Owx9UBU
ybBPsZGAfDsV1ylharCYV73OKbKpwmvopmFXfacAcsf+ZKg4dj85HhJOkLbmbwhu
Vi9i35Izpgwnju4XLTpp+6Fhbx//AimWWgIUDV89fgC1SLBxPjpQwyGzvZa+Lgne
sveQXNPH66I6jIW5d6U5xuoiSvciyE01BBuuTsebZZGs2ALZKxvPrPJYCVSXdYy7
oFqTgUYcobiwc48l1Ot62s4FHGx28Ye6A0lbmyuCUl/TqxSGlsvDZllFlRLPiquP
V59LE6Nq8ayomiR4fo9H4mzxRnXybQZbWKADAYCTwuVbBtI8KuwsM4lo/8yD83ZU
ZjWIeaGXMkyBt6ebB6GDCd8kF+iti+u0lZeSMKPPT2MM7hwrLl9tJb8GXa+Yz6/x
AZoCRJawvay/RYfUhkLbO3T6jQqLompDHex/rqL1DQDlrImt4EBRWbrn4NkQ3UKN
3bdMslcxdhI2G0JnWrzW8yeQTNQqW6naHXGI7hhtG9pWf26t1P3Mu79sEsDa2eDv
sV1MDS5ZGTBSl6zkZ3hJgGK5tBQBrchZdE93wXX+X4fckRaSrfCvWFo/aqPMtm2n
wyMmsBfWP43U8KzSAy4k/4TPgAoz7PPQ5yDRWCzaKbrdYCRV0lBPjZxQf/C+en8h
0o1Dv3i50iug8+HHChT8OA8LVyZi4d1PEiSJ/YUESO+1Ard6KAHKF4+uZFqXSVsF
wHjWsLYFGHy7JouREsVMNU1EF0nZNMFO/2MaUAhDQZAOCvdr8AIPTCpHVZwQKxzo
1cXDdXD2QrBVgpl8QcA5H9cZHQlK8lYWZYwwTYS/pHM7OSuIvc/YDhzo2kZZx0Gz
2Btpwsn6LdHlVhX+fl0bGgjzjSbgTIWpoKuCOxm0RFv0g4EQ5+uaYyv4bOxR+nl3
AgFnF5wvu17py+Dhx68ag/Pt4IbBb9wqMNR1gFv19BJA+Aue4Zw0fKlrGwRvlV8D
5QX6m9sdDwg6EyLF3NgIL5YYBwMam0dONqkQ6mdLqMvS6LDTqaRgUtlSO5jigouu
5ly511D5cZfxZBZFAMrK7977rgcMnKh1A15mXcSJmZbbEsgWT60VzYHh5vEkHvRY
l/4/b8UJPxneFC8EbV26vFhtWODtCniTHo0iyoMJ51nmFzjlPXsHy6ZA/RrF5rox
tSiQrXDe9U6Z+ust4Q+GTZp/S8HNuxNOXtbSMxhSHAitzHB9TcL1lqIV0OkxHtAf
qV4g4w91/kME/kch1j9M4T5Z1/j9KEen6KxLOsXs8lQ8shszQoJUCSzTS9SVhF/6
Lqvzd3Xyibr5A3qD2ZB8L+btCGnXDx+cMkisEOCIc16f/S//xBZVlLqkpDWPTYoQ
r4WyQ/2y/Eq2oIcjYzLsTy2id+IK8IzgbSUHetM/U7w2rQewlCDrsywrOz8OA5/C
2ROAe199CS0VFXJCczOOOvcM9V6HB72fskgsVpOC3cQEUW6fE7DKBmQq9vPnAd2W
gT1OL96pD0ZAI7YMvc99bAKYAbg/HNYJ/xEH95/NDK3k+NhpHKs01OHR0GGCtk0Z
DgT5F6GN6XRCcsI5tCuBVDENxxyMNo58aGLl6zf2SinuuJYTtkWe3S2Rf3wetTim
C2+oZZkqhrm1bR+grlC2TGOgK9IcpE2OQH1zPVzxeCDQJK3wj6OxpUMa1BZ2rqzk
+tJTZ83OFCwDCdX3COYZYHUAZRu7/x+KleXycwVY5WcYPg7Hgsah7dhk1xelNBtU
RXt7yjtmfr//JmMpHtt76tUgis3aeVEYJYh8nLRmwCXUGbMUkqwCaZbk+qieRQDA
OLvrJTQeuQfkotRvMCgMUoERmIpZX5AzbZzrfofRgFjO9oYtXRcrZqkcVU9OUPil
FGhuFnCOGGzE9kgrm2rYSkFt46785Rn3kF4xwOQNsob52zdzkcoRGTLHmEWnrzr9
098dQLgOSbIoFO7ySdzc/jPsGdL7BIJ4DhZk3NFL+Pdx810kd1JNf8EIe1R3VCeI
CxrUhl0BdyrgOgTZlCjcBZhguP9gs7LflXBFneUefDuBzvSkO3it7d27ojJZAEQy
C5noltXL+5g9yse17+WydWRKruE9O30NXMglDD62G3HUp31dqEKNSeQL/N+7Cuvt
cvF322b3vLB+eWgrHBQZySphPGTgZkLRu/MW2OLvfCacPF941sw5DivmVjf85MSB
bv/UCOd04/uZDgGmGKHIy+N3H60MEClQmOMM8cxbl7VePRvR1Iym7PZqg6PkY39d
nuWc2YXGoPtV2uwQTKLCPT8XibNp3WSzJEBfTD4STyygANlprvADtJy0Ubvq30KC
XPuNAxstiJ/NND0wx2FP6TB03ASr+Dni9S571Ito/87Ors5Z6qqP+n3l9HbxlbnF
MlgTvMO5taRZLbUlbMSfaY7zP5NrKGCnW3ctRWAL9Kn2HW2eo+PeERtcCC+tzGF7
Ics4zulTW9Z1qSmFg/EkQXbBGPZfJCAPu67D/JM0sNyhUGzbHrvNWMtVQhe4FzeP
FexKP+/Mi7GyRHDiKCGNirFNkNSRgwwDAwUD7DTGTMY1iYGi3FlyCqbygh9I/ltD
71JjPaLAf3VeEuCoYlmM+DGmSFiG5m05DZ4DIKQG7hhO0ndAVRAQI1/KaO9O91Wl
gm2mnQEFzvBzJZhR05tKQdXBYSJv6DQCEPxCFm4eMxE8wrerV/S+DR7JETSXZ8X0
0a3g5ZvtAMNTqF7ZAjIFHPviwnrJAzhadJuq8YbSI4Gv+ltl9vCPKzPEfehp0mZ0
UU9UWNsyGKR5vEsENW2r2lScHF4dPsNjdcIPsJCKGfIeEUaJGeKG1SPrBPLDSgFR
uqaaDmC7s70SvcpflW9YxxXyrmIGrs9ouj5KfGps2qUW952v4+nCYLUkkMVKWyVu
dK1u1OkRom0RBcOAMP93z68Zkl/93OXVbFp5ARh+5ijUe2LX5wRz89LVrlHJDBW2
OoMdg60Sp8pleXUy32LtHRjqHt/QlMZgJpXHcqH8FD4j8+sS5JlX7FKr2ClAhxn9
eoYe2yw3OTs1NPCVjrCpCBTP8/sZ2J1rk+2O0VSmMcfWuztlsAbT7FJCrUIXHIkO
cq5gv0F6NQRuTZ6ls8ekljAGQLb2l6rJbO8yB/EIxxWA9SQSlMi+zHrn8dw30165
txPjPysyXwElMszAc+rx+jNhmf1m/q1iJUgZbXSLybpQ84vD9GEhe+3xvtdT8tiZ
VFowFXdcV4MhMe0hUtAhkWFajOMCuaNQvGjkv+lrKFchXPKxD7zYCtZU3rIckn3i
OUmiS/Er9N0c+8wLod9CHoM1hgdHDhGtOKqXYv8v8A0VXaL2v5g9dauh2KDDZMwV
pGLlERIXOEmPB9ZOnvaT9t2TQH9mkMrPCjLDVr4O+8J2VCtAZp3aNBKVU8JA/k8i
+JPe+mxJ13wrhEGUxKA0QYzt9O9g7qYZMYsrBck1NYQd7fNnEMs35Gfb94AGBAX8
kN8129Fc4Zx7ZiCzb2wyU91ki5JNDRhAeL//aot1iwT+UNmhyU0Zi9hp2tu2lICd
SVMfwxZPel5dOg8Uzr6xZpw3pLq9NyDMbMOP553RBhgkqIgzf1wwzPQFxodcu2Ok
7wpYd8Ra721GhbgU/MqGVS202i9lOZ90LV4m+bWrjU1s9PVCDys8AmBW2p4iwFN8
HPBeaLEkQQGjxbKzT4/TYI46qyVtYSbhXiwL5avSsuivTpFF3aiUtbPjuh7QzpPq
cdBPm2PI9PfgbASxj2iBxfI9mFY+USE5oDAfyUevbhpU0LG6Ibk+8CgGJXuVxVp9
VcTjB02s4mvQJd7u3OOo9eUEOIEAyXxRKkH+vIHmXwZlZMkoB8RrkXS425JqaTvE
HQkfxthcLH1sS+Es5O40J8bDLElw3r++aEKwYJK7QqCWwY7JQVeE4/bHHd5Kyyy/
lKnJlPsfsX9FJmlY+AYURoRGFYJRopzMzXfRhMxlF8GgaTVVhzSSX0XW62xxbCUW
rk8MMVN7451ek+YTuwhMzEZi+lk4/b5kNxvR25gpLD2s+oED+5IAt6vOx4j7zd+p
8ahAMCn012qEzjIwu/2mHFv0LzUUoq7L79diScQpxp4jHHxTYsABew6yq1kuOAm8
nstk7KACaw+vg8LJrmRsbdd8ZfiujpQgyYeHcVjQpztFRlsQrkkjYBH1lte248Ta
9UsEmWVEJRQYOR60sWKPyuSJPNwvQbONXaqOf1jp3hajfoOY3QxX/pGOqxkGxEV+
7EJ3dXZhA7z4wtfphr1/hFRyqNDHck9JnsuScyuvaKHI5kHpQY4bi2cymXGwsmQy
UbgRWpVyokvYAkmIGKa2ZclvFO6GTa8jOFMuo+wBKRWti5A/86k8/QK3KJ9Clx+7
jVF2CXxX+3Gc0bCx03HWpkUUxrneV0rokHLEuebtlQS0f2+zsCo7sg06HpP9OWMW
d1X/jMeUyrubBEDxoSpUJN/L0d+EBY2kaZ8J7ACmjdWk6wZArG/WyPkhspBNe1cS
YPhb4FN9SA5HdX+xXvN9zXPrvL4tFphn/qDs76lKn63UrG6LZG8wWyZsLQ8rNUzv
rGscjrb+EFzOeeOGvyWqK4G8kzj3PngROZQBawaDzWW6VLNemp9jLAD4P+P3eUnF
6zuS69METeBUnZkNc7JNzqhnZuQlrcptk5CyGJNTMJdhJOHIdRf+S2UiDWc18Xbz
/VOJD+JkrLk3DCXazE+pDGDJ/NPl37Mc5B4z518btcoEBvGMUhkePW2a2j67ElUY
NQKCIHbiEjvyRO80l0hIL3kbMJ4Nt6TKYCzX6SUXVErIVmmFhyEM7YzuxbGAl9pY
B+IfqaTYncMAyRILepEAxXS9fykXky6ptmaqX7qnqrSE0vy3ORkp3Fm5uffqqfCo
3IMh2geiLYx6otu+ErvDftgN+Ako06sO8SgYoo0exTaFPhCx3XF5ibtzlLOSqED7
6bjcbDgoDfwnbXZkVdDRg45DHWaxaJt9K2+L2UcqXMr+/faiCB+wKaKh9qo9PYc9
6i3ZPKYwh8DttD7ED7J1yznSybe/4GklcN1FkV0Yj49QP1hG3UJMrxGU4w48TTDE
T+meggWobmuOajJhyPmSMx/DXACe8X8zrVnmzaEweobj4eAcd/EMEnz3GD5Jx+ho
wCXZNjbac1vPFNA4fHlpih28itls9eG9fbQzEQ7Oy6N6OlHuR1E/sol9qh94qV6J
iliaQ36SuQHfhiGgHw3ewxlmkzsCISaxh9DkwiH1RwIqKDUKA5DFzBr30os4XG0A
BewWmjVre1GFxuz34ITSGeVymsmq7oZlCjT/O+8Qszk0m88AHlQDVMmUaaiM2Fb9
BJFnF6zoMRpP4Bf1vXYke+IOFAu8QmLeumyjSTPtqUPPBDFZH5h9SyqqXKaeyfBl
dtXQO0FY23fs6WROshnHBP3S7iwAaScR1oyWSMx0GVc1vz2B0wlytcXAy3ISjxfz
MyXvz/deEb1oH20oqb/YZD7pPHA33ddouc6jJCLPNyoXE96SZLsbALkHGmGaAREf
/NWgDFTpu0/RHaA0xDysNXrX6hHrRBElYC0mKRxGS1uPCc52hdzMMwjWMrBtUAGX
zgoEl5JnL6UZOVv3gP7jVSs8ySgOr/P3YHQ2O/H2QPE2l61wBNiWFTVugOZmAuV0
smnK9ZnuTZYfYmmo9r14suPp7Ez+qUkNAGe98cHzcHOFwz/ZmfSPmhu6e3XUELT8
Z+kJUSGKAQEnZEqZzcY+hWr3F5WJrzm0ZZvKBzrlZ+MdU08wdWEx4icseLhjcccX
rHF8d5ikXaej0Mwt3lS+0dFnycnIVu6NGMulA0ugzU3IQfZFh0zDMMQn7I+X9IUy
reK3MEhQJZ/aUyqHOS7f8ryhnwffGBz5miQWB+rb8P0Fn+4EtpBgdYEEhwK/7yey
tlVmRijOV/MdU3oWJ50UrjqKGT9RXr4QnTwyFQQa6gF+cbc7rfwMegBNqTO1+Lb8
t24KTyy+2E5V+KIPOuE7d9ho8hxJ6Vs1ag+syJVS89suB7uFyOG5+8mcm3taaH/f
SYF/PurC1MguJHtcRAPVo282fdt+pbZX5bCntcVEAa6QhunoFzK2VM2y7d4EwVSn
dmOofF31QC3CVDqYiBB2pdDJzcV1ViNdIjcuyH09yTYI3eziYbyeOCxXKTtaHWHW
mRNtL3h1Eh2UeWMpUrxf0wz4ItjSQwCfez9DPF6CvjUMYgyuxup7CA8s1ganRGBa
0n9l9Ena5lghga7dyMbfOnEbNPyirlsCZ9Pww6DHRzpCeyiZC/tn3M0REvs00miC
5Y8O24dwKgaKZyjDLUlz09UOGSHXX5KgiUXyqxHNaCqUka2JmpBlT+wygMOtwUU2
4ewJtatWG//Jj9K/xZwELPEQgMvnBhGzXNYh+uZQbJD+sHjxk4h/Sh67krixdYH2
ozEO+haS2wl//Qe/h3u8V9eCxSq0Mnon2OnidcYU8OwTN7SnFBik5mhDhq2LzQhu
BHMDqJaBetnJyuefklAxuU4ltSNSuONDyCr1jlgQwWoP25T5OIEtnAoWGYzhcDvQ
aC7N9rssPJf4/4G/CEbZJVsgEycZEp1PQXz9lYEkr+nOM/j/Oq8gy+jWeU/HV+NC
3VKFrWf6IeixKdvaYv3ZUho3pOtFR3srk8jJdJO+jizW52/fP2yV6qlEVon3KX1N
lJwsq78D8auDMxmEWERrtgy3wpxepKMZ959VyvVpkl0JT8iJwp79K/DVcaXr7vv/
WfiFp99S6cJvt35ZL2SB8h3f95+Tfe4STFiiGZeWB911Hvor0yd20oaqVHahh2jZ
jwtqLM6LhRKz44a7gOx1Ef1upbsJdS8yL4zAa8rj2BKYZTiFPY67O1zOFMUJK7dR
Yzda3tT1Q7y/KDWaVi+yV5pMFxTBfvZSwFD61f/KI5BSr42I/UFj0OF0qPQsfNq3
bs0briR1FBUsTbr1Lp6PwUx7OBQiNwTEBGh+AZHP1h6lEZyKQyrjJPbSoO4v3myp
lUCGeX6JkZWmlKKMtRG4IeaKXvKDGXFDHedXwce9k5WRt0M4DwUmzosgSwG+V4fe
Wr0Kg8Juo51UWm71jN+QAMshFdsS/81wiBhOzXVSu6GUIS2by16CM42WfbFrVSRt
SKDsHhkEx/ncRcYzVW6oxb+0S+YPR5NvcIpOgAfWj2me3n/TGmCvX5S70DO9HRYk
43tC9OJHM0yxScGveJZLdll5aMSDNe1KeawIpkdAzd6DlTp6bcYbK6mZImHj9u5h
3sRS3xehgv72NNizNNx82Ydr7mfavdQBV5kFPOJUi7LuvKLYEU1usReRULsGQrEp
zHRRNAs3ofFqbXsaBFktDHNFR9sCA+kuWq0UcUiHS68S11Qg17MO5UVKU2+WZlwD
LLa4D1GwnFrRD+53AGkG/ZCuluTHusMB95HkNxfo/2sx+w4t8TvkexuNZgOv+1U6
6qzqDvB1ITEFk4+SZVC8lhEJBzVCjGhh+ULTbVNEGvI/y3r4TIh7au4X1V8vRPiq
pHcHVM+ZYi1lPczqpsFw3pLrzq5gtFy9WToGbfzyHy9Ou6yvvaCthVUTd6daCWIQ
tB/PBejdg5Mx7VBOUeCCwplOpekDIOBqHaCnIK/c8PRqPfBYiNkgxoKz6PQU4V9X
bPsA51enqX5pjAPIICynLOB7/oDYPAPv+0CM4MSmi/oGAhu1rbpBZG2rhC7FYGgg
g6bKp5IMFei6xMYPhr4HIvvGrOdxjndb8heYSQDIs5mnMBGxOfjDgd5vT8JZF915
gIi6+/tsLPJNpPM11tnFrOeQc+EWAjWdD52CMSYr0gAqWrJoFynli0dTScbwZC6Y
USEVsSzrlbQC4JuvNZSHbutXKyUr8u2eIWi3TVc8IBZyaYPdVWeaR1zOctNGO6pL
SWnamuWsKf+YTWBtcYwWfWmahnW0KdRlldUF+7L0PZKfN5zPlGHsT1bybdw59eQQ
o/BCgkGq/ife1beSEhy8ckllobm57geVzsGUhExgbe0n0KLmjbfCEE7MV3Y7pywM
CijtaKo7P+tVHYr7G7NUMCPSrsdl144cIi/nZucBShr+3l8uUCZBLl7OOFDIY3g0
bJc64A37yXnGp+i00ALK30O1mIjojAbBqZPB0OhdftW+yyyWBmc/bXLDXUtoxwV5
Su7jgG1VKJwXu73qfRjS5eqjk+SL4uEnUxGDfrdpdr7AFUNOpgDmzo1FePl2kuyF
f7xu6MhW/xisd1r4iS+QP+6Jog2BJvxg+08X/UnXQ4JTWFFtqWEB9rZlzD2XU3HO
uBRC3D6nNwO9WHrCbrE1WzX4wTJLGx8xhbSMDx1nD4NbVM678MLqOT+gpY8Z4dgm
gqlxIJnl1FPdPx8N0WIpOXfeM5gwYfSZCB5ch2T0AVynSlDR3HtGKIALr/lW7eN9
2hJYcGNcKOrFhfGd1BDmln3VQMrt266XCkAAqKwXZlQAF+jHzfXDdTsCfKhXe0ae
bWUYqnPfpcEYZTupwqmzT3Hj6MryLVYCiOijh9rUJkFuZ+M3VmEUVLaXf1wguHO9
scTpTPLox9asoQkg1vzkRVJKPdAm/mhLcAlO3ssrr0jTCJQmxG0Qk0GKQUJmzYIQ
qILoAYSCvNtGv8gDKPQBQWfWptTaaqnbKAacbKf0i7uZPoLSJZN2SDSta7Ly9eTS
v917lOzrt5dSOzCVTFj3YkNd/GIJJXZxeP207oPdZFgkL1elK1bVDPkp33wuPH31
8tX1QUwwF7OygT4aLnjlIzRb9juUeURyAN80mb5zAvI8SlswdkVS6FGZ/ne+WiDy
saefnTz3taH3YXQCAlYbPRFjvDMblzd69m+zDBfOa0bUOFYeRKsZmy34OmWQzf6e
pA88gJKxHzJ4lzTT+ylSaw7nZFouX5scCJ/ZAYt/jI2Zg2cC31tD25aiR73YpRIr
L10PEnwYwy9hxf2PDtSITGSNVSSRWJg8HoQt8jckDCmrtJ5+2m/K56Ymw4iNy0dY
E+JxvVtDfvCFz9tYyb42Tn6+rPlWklJHNOoF63WE7z0z3X+gKqKjlonw9adliR2Q
OCa1T4zFHBKnA6e5UaVQlAqgEtcNZwTmU4iBceBA8m21NF+/Fz79L5z5wzIWbWkc
zjJgG4DNz224cz2rh8f/mfJte+u+MY2ksxbRjZ62qMe40PY76zA/TN8j7h/pkESP
xMkU1PCwc8dPzcs0toKqJztcXM3nGvHYKFr9qyU0nu3uU/Ua7fcF5QXKg49i4Z+a
QdKvRBDrIbSQiI8w4fre8x0alXTkJJhnlMR60cq0LAGjG5u7TPzxTtR6vGdRcbFp
hKmWyAiqsR2q+Dv0KDz7g9CbLfR6SbPozJedDcIB7gKG0YUatEus8knMvo09+/1W
BiQkrGMF0Y6o0udxpznWxoHmYhXXuf2vwRXclN2zpVUsP6rwKlOenmM1TzgnmFuG
5jAa9ZOGjkgXYpdqdW/g2HGK6tMTb336c8YuOhhq3n3SfwFl5xyVxaCxV76Juwa8
aYOVKk3IEVdWerWQg2vkLxeP7M2yIMm+lZsjo21EL60GnpfVqcG9Sx2rq3e1HKgK
ip4pMkb1GC23rnUZh9EuTbI7CIUPS12dq6KncDkHHzSwmo/XZpUknxdLwqjWiw8d
h0kddpO5Mo+aAY/zPW9pfHwbsgGCXRKQ5kym+y9I0vtKU6eMj6yNMgdHOmOvKeOi
d/bejCfeD6ZYDElP0SY/HFDQLDuUXHHuqDqEV700VEE3agfdTSC5UDe5u2p4BRwL
hRliKnoOTVXomS/fFLDAR0DlkJupHod9LMz065UG679VoUeAe9bhcEfQRvblalJb
uc1TESREzWsL0AL2xnHPd7MBBAf5BaouubnVbHiShMGIj+H5Ds2DBkIOHTQ5O/zb
JwpdNw9QBK+3D96lMkF3uSWD5xy02gGHlcIY5Cc/2WzmLd8/0yNAwMij8SWcyMJ5
WIoe6Zgven4KGox+VwB0b+3AdnwCfWHkGWvqUcef+Wizy46yjBQDJTUUCYelTJ4x
qXFCiIiuqjKEJ2VOBt5iJvY+zG+qC7ZlF15K19BjZ+4ydsq5++BFIRXj1oB+NHwp
V57VNibBQqlnDIAQKiFcNvxxqqsSNpGKJpqYBxtgwia5Z4yrCAWOunnT+ZfKkUjs
R46vmJBojIU2aKcTRzeuQb4XwMuxvC562Mx25LNiEuMxxlnnLUGvhqrp+Tw8CFFw
zpmfAOWoBRE5pD/suqTnxW7CMHPJ/CZP+1UEGFc2X/rxwhDmIzXXHF9bD7abxBym
LNbhZKKW+iUPwKZCAmGV1ZGL8IE3Hg6kmHQkmAI9kBaSAqhDj6Dx5xHgx31jneO8
5P1nJCNSyA/PnQ/5yeOZkv+GZKYtpV/bvYIf1qgVPIk7003HErgbNyWnuPV5Jwc+
NOHmjusBWzXb7Xy71CGoapakRV3EQo3Sspky9XlhI9hHLiw1dbBTdoFly0t7V6oB
lqONb5ukE7R2WI3qKXKgPe7K7ekJaizx4nONb/O6yP2lIxZwVfKmJ4lBEr9w8Akq
nbuUigzaHb+LYTMCTPE5oyoJv1wUAuNpiOolt/otI642DaXwYV9lvQrl98JlEnaH
4KD6HzdAOivrUS1y8CF3PKdlBmNqg/H6zPIhT2LBjVllM/e3ulThqDLnyPEWuqxQ
sYjovkDtnSMqLj8NS0VwHYMsyRvfU6CRIkv6JJY9sX9p5dsp2vqwNifEOeUapLsX
HqED3ZzF4Tkh5ERO3Sbpz0iIYIN6EPywgD4RW/pD8GjGe4Q8OYbbQdyhw+56uSTB
3a8grjPUTgIRPX+6KwnqyH05eiNb3yDcU7nKcK2yQOt26iYCwheqhcq0N6IRmfw2
Brgbta2LIdnGGnMkyRTn3mri3a5RJRvtFSovvNJ6Nhsuohsv5cqefMUR1bPh0LQ3
NHjDTr8H4YaEZSOaDNFd9XtUeJm3hMzOuUHur1b3Ppmo2rVpAqFqBcmAAQP4TXlq
/UE1yYx9qFgjMmrO5/AVy7MB+m+KNmAHWffXqscSmFqAO31Bb2C85Pf8iqIgI3N8
sQLjQSwJMok4DVz4QgLXr7cR8QHw6ztDUV1X0AuP2HdKwQ3rdA+xdevKnO5dW98S
sGx0DroGKSX9PMgw4DQ1IWwhROFzzdbOlZnwJBm99gPbcF8cYo02p/U+6QT0+C5Z
tuGqYUpfOEjtKietOYoN/6afMRyiiezBxBpouV1JO6tuy0vKrUgXihkKaXW6rRjm
dj8t4dqqDs+mycH684cGfGmBVLfI2ih9FycFwtkq27D1L4W6U6eljkYId1xAiWuK
7wWySS0H26TOvjliZVoWqYznKDzfvZLdhxfixEK/lY6woEViqGGiVp0EhEIOOpHH
3Zb7OuE16mWFC1ew5l39iURMlFsA9OvefiIwIYr4yuFRWLDU5S89ysqGUcxo8rp6
KodUWzTneLfhBRhc2CLng7pR6a8FoYJh54XBkp8UD8Ox/3ortFU3uxxLgqZYBulg
2S4T6sNnWS4pbz/Brl2caHq9BrrTayIJEfx/m2J1fad8vfI95l11uag/kDqPKPP+
K1s1k8ZW9ndW/OErJ7adRtgiQYZAMChOnMgN4SqfuOl21n7eaQslIdzenRocNfUJ
uP7MSo2VrniM4aVh9IaTLFXJEci1ccMIyuFELCj9JNEPudMhiL+0jSISxK+bG9pW
F1pr/6+XZk3dGJMyj30IEgFzlzFARrPrCHTbhaFtqolwcM2etmEf//1ALG2970Jn
KQZ2tIODcxBnRY/1T2W8aiqshubJeFRTpgzybqnmQe++z7jbh6KI/yYwE8p8qh9N
dhJrHMXKZOZh5JVTYwyH5CozwNNo3No9vQjZqZK/n0U2AAN0cFw4RzfhfKnkIige
gT4Z8YdMO31OGSVubMJJovS19kBCatKbX2LHuQIKPbFgplo7xmUoh7wkHs05k/3s
4u/ZawzLhNu6+RQjvNaph9W2sITLPLbBCcWGLeEk7fOCn4Nlt8vAF8s3d5U60unH
6qIRboq4AP1NWFq3gn8IbPDr1Rxl6BfrHrgCSvLAgVp4bFEtZZvm4Vcf0xrttHsn
rv3xIXcj7otr1ofFm+3D/VeKb8rS8NKJqKpU4Z0xnyqNIPTEhW30vGQpodYCXTWP
EqbshBi2Cfivpmd/T/Ues5mQ9fFRVIQc9VESwA8xt4YTTb34FqExOw4hMv5rcugA
Sw5zT/E4UeCukkuakKwW3WRFeQKwEGhX1U6Zj+4dmkHrO3pDkvZsDjW5XlFXQhXw
N4w3j4/8JjTavOEu9pFiMWCerfF5GHOdxfpnl6FmTJSxvm0FBJhi6nI5CosC7HdS
Vr7FkIzgpihk1ihOR1nfxTrmRBQlAr5Yt6AtKcbOBMRUkJoJnIMzf5pdlrmB6laE
kp14PUqVytig+UXgkDzE53+VpaXqSdkW8w9Q/BxSMUDSY/DwY7Axz/PjP9xrc8R9
8MAqPtkup+qz0clG7YctMNZ/OWLZ9uEMX2+vHDK3uZAriBGHpuOWUExj6x7Od+8/
+EzGZGm5Hn6KCw9cLx80ePGLun37G54DUTFzDJa2n8Q5LTT7PvTfiT5krcdERVWr
Ofh5C5i1ocvudyDbkT60H8md2LBpThxMzzxUKz1+80vsQh2/syiTJjL1sRRFeJl8
2u4NOt0ytoZWzJ1clW1oi9NB3QpNQb86SCgLsl5mVXEKiMGkmPkuj6Ak8XDLEHZZ
a6XqeSytZFvKG95lOQbi0mZ6Di93vIXPjGMbaO4EePmZTekKTJ8QdWmtiA3LKyzz
kKLXKsSNhWBqbsKzxInffQCvMCLROIY1LkmhcZuBwap//sCLeWelbbvD1rn9TGmt
tZOhIeH8apESXPgl1wp5MlSicRQmvFiYzjs1HPwDMRW4ldRm1v7KN1JfnxMuQSbq
N1XnnGrlXp34BBpLV2QxVrXmzI5sqCco8lRr4TjtXEjogj88HluD46vPdKZ/MHO8
2wF+pMgvVGIsEvhRFdL9kTiLM8OTV1XNZl8VV9cQxH5sxG7GXO/wSLcOmg0szrM+
sSaF5UpN5+rMg5n7q4XhG8Oh2OAEMdh38IfNxEtKwlZjFu+82an11WhZe3aObG4H
uLapTm3o7hoRx+uCcF7zfCGyf/LJttDeX/YXXaC35cbXUE0Xu7GHb+tVego328WT
/fbdT09yiFv5nC6baoFkDqE+ixAfZWOYgVDMXIUGtQ9yVI9qqxLgAYMGMjWez6kA
E6JSVKy9FU8vaTxv+7tharp+B0G0dtUN4hhMJw6+SNnhWWCR2rn1Ujc20l1Wqruw
zPurCsHfYV818et/fTUvhcFPJ8Zs5J7sAL4J1PMMFqaZfYgb4+UGRDK+932Rx8pO
MtXzoi1hjzsa7HorY51io+JKt/EQvqJrEuvfpE/UIctM86ibOf9OhvF+hOYn7MFa
g20XpAVKwUTbSvgD2Jj/zstBA2fxr5Tb5z/MgII2TcvhlUwTbEqZuSLbQ80wVETU
ib10QHhHsQRrnKWS7i6O/+MsdcL5N5Ciwtsy/FWaPBlOECrOTi+mAyDSKXRfHoQz
sWal/Z0CIT8GOXzcEDdeRTr8sg4GeJ+YnXdT/62XSGkCTGOOmvgQ0A+6rDwf7Pfl
79isL+z14NZl6zT3uHvb7QpW9yuQfUgG+y0QLXn8pRpXu5vrPW9bpeEYvpS+j0/D
zqDg874riHfZbjXnq16dJxNPiDJ674VIInGdessYBbKZ1KnKMb2eXQFq2f1RNAEH
d17hh1WdFAih1E3xKiuiCZWKOyj3UuLLV8KXn/f2nn52TiSZPJm5UsxzolJiWECG
QFp2oPwXumKMyt7bHstIWFQPcWaBqcjtRCuHo8T2M0Gs0FxDhScBMlMV8Jj2Jt0q
4370Ef6LHgAY0F0EGYw1+Ubm9macsm/PMq71uTxRbTUYFkrD2UwuQt9gPzS0azUr
YGXtopdYOnb116YuW0z3sCowTsbBxe67U3/qhJh0+T9WveaHPUzKjxcQL5YiHsdw
7kzYFV+5O0skMoN8yApxGBRbhmva+U0A/9PEqc286t2R6RbMkVaKwZp5Q/T5xZO9
mflf68QjcsB+5+rGh4xSySl7zZ3UISxUlCu/hpP5j6ufm+6H/wlTDDxwT8IXqrrq
1zeZhkbEQ3fsXx1Esa/wI3LsA9fuMHYUKsFkk/6pJvOS3APmv2OlxBATTvG6LIsj
qScqSmuE6CDxs7BNibymjQU0MdewhdrdSTenZEDJACvXcx7fb2p8GnfQkXr+iQu1
OF+MkaiZHMfghkqNiyVnEqKmyNlCQI31sI2cJNiYIvC+LWZzKUhVwEks/4BWrIQE
BiPQXq83NqDtJ7qGJSIcFTt5SSKX9maEGJs5dWQ8hlQUBAQZ79mcNc1rxcmK+Hpi
u/TO0uwkIvNIrF3TjpOUEfIe76q5fyU1v5jyzsQCPWvJCur+tKH767Qcpj1VSECG
6nnv6ryNVGCEKgoNfLv3Sx2Xm9kTk6x91uO7bETwW17MGhUgx1gmesm0At6QqylV
S6cxlhaGFsR6Fz3PvJpxo8EcOpHqXdQZaRYoc+TO4VgJc+LVV/UJP4ovNdBbiKUj
3Na0dcmr0WtRevWbahSrmJVs8xoMpqqGtR7Uv1euNvBbCwB7OzDz6lQ13C9TVvjv
s1XpIF8HLQjqDSSaP76LP96PkeeOeQ58EmvTyAtHN6719isAkBZj1YLMwts7X8x6
IQWEBUhYU2oZpSZxLCitAsJOMCaIzE4+92zXQC2twZkI40254w5maVAQoAaaQ0kV
vVNHdwUQjIcpJuactIqX8IBpkNV1ndNFv1SfOAgU9kKcLgI6/fE730HQ3wcTdWsI
gIiMFhndaJIbdDuAzgHyCcyQuPrJCooeT/mS5/Jd1Hj5hsBr/5yIy0Jsi6X+ncvC
t8aty+pKLyMXOT2KFm+EB0puoCZKOLyZqJkBYiATjjyp9lI/HF4VnW6sA3uqEWGs
wv4CRdLbDFPQoObVhcycI7anZxmeNsZBa/ulllRpFho3+i1OSYZ2j6rCUfwPsMqc
MoX29eqkugHQST1XV3J6pFShsPhrL8KF5EZfSrmZe+AiL1c8UOjGQkyRrM5kHMNN
pH5gYMvW5KmKEAJrcOx8urfqhx3ZZ+rdWsixs9dYeOB0RtHc3j6WLlE4JK5ZkgX+
uRsAF8e70J7Z4878pZJ0F2pebhb81BrLnt4duGo+gG3A+rSMJLJ+LcuTlaHEJDHs
O8s0IVQTIdr7QemutETyd5gYV0l8u0NtSX8kiCh/Dbw5ZYrVX3i2vGPHul1MZibM
T3Lh+wScycbBW+4eVuG90rVPeckJYoq6dngQrWiA8m6xC1ysXk1rigKOTwjts04m
OafDXPXaN4j1HAjPQI/LYRCLDkhZfshwCbygabNV58b5YUu8mys5xnVNOxPQsD0Y
9BQAGI6n0vAeTgci+2UEQ7Uvl9MeJuc1QI3VL1zRVt33jERGECFud5YAR/QPZw+h
jh7A66KBaArRWMudL5CdBT2dCBJA6TxpWW8ze8+U+K+6h/FEgpXR5SShFBme6KIu
FIsUnWGBW+nIW9uvfNx6lIJCxSAVbi2zbllz2HpDOhxbP78o8EghLy5RyHjbSwRn
TUOXIPVPDjIcMwKVsWfb3F9BdfZSAbJxKhO8aw2InIG/Fu364Rkmok1Lnm7PYSUw
1mGYjwoeUMjc8EsZ3chHSEWlKi1SXsvkFBVRfhiMZyttmwFoJ1SaaXtCEa2dIxWb
hFuVfUxnNyL2vleTKLc3Yr8W9FYW7UScdxWfiIMPtkLeCoH9GScuStgFJlcbNy5S
Ztc8B7qOzlnCLPIDzbZk3AkNcNUXDOoevajrh3CB13q+PJ450yV99HHX77JCQxsd
7ykLu7Dz/daRqsIxplFH8DxX7gMPGMv9CfulJk3XI/+jszhsVPgPdOxAW+zwBtEt
s9SC/PVbcCNZkE1VAJi6j58JYPzxmlLgBHm1MnPAg/JJNTv/NMnbkT5/gOu3s2K+
p4gS+iGpwucf6oJrIVj84CubufSfIWdNaAPyo/G9+Gl1e1lzUyOIjvcIzlhKKLAQ
YpGw/gLSv6m2XHvEYRXyZeNQh65ift82/3Ko/LsFr7n4rGZ+LuDxTTMNNaNu/esF
wLwWs9EVOwAx/JbMoabr8Gadz6/L4gxeTasblmcNXpYBoqA6MTOWmtjMYiLYApI8
VCHGa3aimKUDIJbmWHeTvi+ZfjX7HmDDC2LneGUsucs+1O/Yy1/jw4cO6dbg2bnS
OlDBVq8oUZJhrWIMwEHImuGQa1bcuXrWiLQMrVvsW4zisMKzZ6oQdYGE4ClBseGW
WmkCETVDZ9wdvfRVEO6SC85GZ04lOqmOxvK1vu9+qYM+Xff/ntXS8j9CP29lTF/m
zFhuWf39uq6k3KPcrJeWxz7cv7OlD8IiwY/4Y6K9Y8pilb2CTERL3kdrPtCnnohw
xhuS4Mbh3ErACLBygVa66WnafH6rVgLitnVr00G/mr+pxinIIvfQmNeBTz6YXBS+
1qPUJeiaLZmM05aUg8CvujWmouzhdYQscUUB5MF4fD/QniL3lWiz6YpYsf9sZkzN
ZfEaxdZoZFhwWghpGF1XiCk1fBf7MmcJGZsPaTBYerprQ5x/9fjl2DGNdk0t30FK
qKZ32jW1pyCqTZSpmFEAl+FzD5zBCUODs4bpaIuM/VeRHN4D/62wmaE/QubKvTd+
QRYvHwK1UojxaD3p4Sf9yUEhIMI2mAWNcLIa1S7p42TFpCE680kGJ5VoM8J/36w2
M99NbhTQyyh/k6938H2ZVeI7wSeooE+l9WT391/gDyQfT0NswpMPJR3umHnfHSi/
svtbP5qkn/3/eqLU/blutRXmOyzY0zubW5GMO0cTEkLMsweHbthiMWBcPkTI8RTT
CyEtL0r6h1gBr0aYXtT8LpeBvjoz4ZPcRiWW8LxrePTqOoCg7sPtQMaCRjKSzipM
GCW+M8ocYbGBl52uOL2Etw3dDbsNvUIygVz6xK+ajkQwIr13IwasW0hlHN3QU2H4
t/AVRa2yQo2UfLAMr2wwjeKYtFjGcXJ04JHSC6I4nWYFIq44SGzw7cWFrepCW6Kk
Bwpv1l0unfHbYOptUzxAdOZj7jx0P0m5uvw0a/Z29bT32GVLASh/DCRNZsqoXu9k
nX5vO7JH4M2VyCjrUwNU+RJ2o49VuWBF/k2IxWUcF1VU6glHgufXqoSwxnNZOn48
TFezisdbvbJxmv5ZJGl1nJHgYmW5KqOEjFAds+kHLodQ8n41lnt3NA7+nVjkN+Ra
sTo1SfPDbAPiZaHpywG6YqQ6pSr2Z4pR02bVt+DzCw/MMR/ZZ1ijUToxyi0WxRMd
Vtx526TfB9/coNU35U5cghndvBfbx01eMLsPqD4cR9htxqhesqujJUtAj9hfNrfd
YclBYIxFbxikVmyRVMYoKyXqilj9Ej/pV96kVxRrmIQMtAybVnE9Y0bciihjfxpI
vsvHJX82kioaNlku/fOurTuvEyIi7DdCs9Z+lA+bGiH7LxbTuexy/22QJNqkd8e/
tsBPQAJhTl2bDIfuPAZAD2QqBJCaMkRc3E9va4Zx9XR0h3xKn+Tmc2NFEe13V6WJ
sHTQz4OMYcg46NwBj6CYfDR3k2ubAOPhq+eMl5cQ/qRRICXjXeMc799dk8UDP9ih
JZw83g3JtoCzuW7jjCE85Y/b4XZQJQYMRZ5Icdea7QJWejuCbBmLXJVVTcOF7wLV
5CHnZsaDSGEV6H6tcr1XPrcVXju7QmEuqjITANVWe1nUjyhyjZ8Uj5289jJw+jdN
EHlNLwxz8H8GEgBl+hZyReNbTYt81Sd0PUnO5dmwNfTE3V+tV+4Iauij1WExMNY/
Em5Qgb00RlOB1nVg++GuxJwjeUkvRuv12GuZyIdjkrLrnywYt0zHBTIJmKRls3fs
OfVn7Dz1+fWl3LZjgTPo1J5vEQmqGQ06yl3PRuHRov2EfeThfL+WiTisOJAYhXPV
JRs7xQaJsdFmUkBnUTo/DdRbiyHCUPgURnsBO1bvhiYp02NsjeBLphQ7aZuXshyi
eV1lAsSvezvzUAB+ERSMlfFUdhxLccP4mDPN3e8C412/hvOoG7jvfhgF4BGh4G0M
s7BivAE9NrTGdBPe3Sut3RxD9WhlPD3ToOeYBl1siK798NKwsqAAceWSrtE3oJ9R
ObWNj54zSt4bzjX5sFtUhxR7kSa+cJ+tyYrlvr6g4nnwhASMgG0UECbvIgzlmHuV
2BaWsV2cKDFYvA7EPKIVjAdnZcivMjw1SVbaN+p0wQdQH2tItO3nrV7WStzqpwSu
9IQp4YeAeHmF2TlBOS8gwVAXOUX1g2GuKTsD4Dncs1b1dTvsM0lhuNQY3CU/cK4n
8Q1m1Y/nVHV0vh5HhtESJ2jysgX8Om7q+fx6dSOL+AesSKKm+0JLaEQ6gvRZ8Xxh
T/knflcpcm1GlWHpbc/TL46NjzNMoOwAyZj0vIcyGly2M6X3f85Jx4u2v6u0kfzF
lA7awTuzDSw13SXTr2JryRQiTUEHnH4RsDGMMUlXbzf0XMCGjwxTgegooYZKY0l/
nN7NwWtMYRwU6CaNie0/0KKNsTwyZafqrhy2wcJHGvB4r15+pAJ/lG1O8esgbvdo
05wpNabggIZ50jFUnV68fKXCx0T0leJsqq8q0PP8pGZr9pH6TlgvhWPhp9J0I+GQ
OJWSI5ZZDLAbUU39KJvhVHSpdnHdc5mpUlv9JnHs/E5Iec5tliMM0TUShn6kcuJA
SmAiNfuaNyiluPYQnrELvKR1MUUBvbxkZTFc97Z4RxUeXf9Z5qkwJz2iQ7YOeHtc
cFFnnStj/ctGjFk6LbyQFeRlH8emuASyo28gSSXb20dq3tC4sJ6lstLp8PcVBuKE
RQSfLGJr7/95vARb6IEKRo4UIlLf1nj2LNrhsBHukPvYC6uxdu0wMZ1IYjlNIdUy
CYbh0dslZjcDWOlNnx1iPqsBdB0yzGo4EK46JiDo7G9b4Xz5qpEYDwhbhS4SVySX
pubPm49av607owX3nAuHQeQNZtelyNQsyxqLnnxgZMTsJu8F2DVl622ZrQ4SA1VY
Pv8BuqgBeqQHWszRXYuchk3gLO56Bm0fdq+A18+Z7RCG721Nu/8JcJ6bwZLb7R1F
+8DLM0FT3hM+aNxKK6dk+64NdITZWihfZSjrNcVVd4xmQnSCXk87O+lzl0N3btEb
i5neiC+Hn010I99EVMnU/XMndiOnbcnPF4Z3DetbapVSAh3u6GGgGNb/y9KLlZvL
T7FAOjKe5+fW8c//RvuV6iD8cL/CBNh5lUuiP9i7rjZHm8h9go5MtDA3pOkEOnTO
B/6BOeyTYhw+ISzdlzO8J2UqGV46qml96BI16N/+GSvV+1PjeUE4ymPV8Ris0/fS
uDHrY96ggK0Fqx7WC96XwaXuYIRw9yuTqkz2S2FWrITk8FLrS71nu5+Brj53l2rO
cXQcxQslBj9R0bWWa9Grn0J+lO4WMhn/mSq2OAWTsxi/HPlrWSod5Rl/SxbN1KWE
uXIjqFTpKWrY5U75GB0pPbmqVYgmLZtHPxPXOLA/S99mGCs15pCaDyYeK1EIC6f/
UvXOfYaqE/AmQXZCqtHD1mxUTrYcobcSkHtc3xzvCqMesWdkBXSFdajOlivdrLGL
uRjLJvTKa7uqLPkRFrM85VMwpZtYN9yfqvTqtBKtdpbAqHAjvkYSy5is2OYQUtoG
pAjMiooi7MISb3ppf1OOe+gEER+67Kitl7yF6C2va2PKYhu10a86XLQ9viYd8trH
B3gMLUw0p36ZpDrMOsL8xLQLi0pRl0V7L6Sx0BN5hWAR8iBbeoRPDa4HUDFLRGVM
0LOv+GG5cfXGaEUj3L4bJ5ePVsV+Ro/CE98qxOi4OASklQkfulW723FUXtsfW/5F
0gQCuj34a4ovnnqXZ5rl11IHMCwN4ArzeN7oUYH6jAll8SlzhvmDO58aMvtg4vx+
JdA9uL30nliHV778Ci+eLbQdWUTkyqLx0iMuhGFsdVlYA8Kth1/oWP7DGDomLobn
YWgQVyo4SflEU9rvJMCWSr7yffEzTXyFN7tIKmZ1rKljN/Qe7gB8hwpFPXZdkyUV
FR7EfXyko5kKKOud3om+7a7/U/FQH9QWAMpBWU+E65/p+Q88YAwdMVmw7x2hEFkU
M03HJx/0/YdzGHgjHQgzz+5K7erJBLs6EL5srpL3O2mvTX3BTkjy9VSFkM1Ovsc+
mKmAnHYUP6tOE1Ip5o6DmnjmrVypLtuDUeiEfBztie3TWYfZT0uwfyQHkw1ycs8Z
2uNIZPhHt18iL8+0AhpZf6UmdRBygOB7NTYkp93Om8keibkBzcSAv/C4nSvUl37v
EKwanfAF7T+RD/IhnMLgxK3jatV6kcSsm8+gnPCKWyAEuScq0vb7WJKAa1eqpiE0
i6V2gaF9VeZ1WfznI1Ke38fSRrybX0tm+5teLqFLUSYZVS3wfTIBVjQmPjHKEFAV
dUW5uMXuUUh9Tuz0iyLwv2sDRtrt4j7TCUL95pgCiLjUPX2fuSYvP6HXGPRTaVNo
PlCVv6bb7cKKv1IiTID5F6yhmHnDJXXcK+BWQ5snVT/db3y8SnsmhSZF9nIDNeMm
/+TVkJHXZ9LpTnM/7GR58/cDSMDZt9qbTVoVx/pj5jDVHD6wWweWdLU7vo4I/jyU
vG0Uz8symVn3fqbWbBDSs3zW2uVgxdHHC1ZsC9GQC1XgQkHZXKPMh38tXHMZSo4g
qvIsIve2B4tfg6iKUvQqUgYje4w9KDrJ78FI7hP8LwFhSHrgl3WC0nSz3Y5gcpHw
6ayblUtJKD4oyHsxdZseUxy9A6aFtbyX3SvoCsYOSJVO58WHq7riQPduuEz4TCqm
jbq3f7YkRcn4MpgLeXLcnNu5FBqfYn2LnIDMBvsSES7d4g2LyBnqrhkBkx5eQNur
BVHIrJs4jnrnBOPLrJv1P7MPJKkLu/apkaiPLJUO4qwJvECBDoT0c+Pkq0/YtzAI
8KTirOhQtMkv4THnFyfYMopWfMO6HeXqYq4hU+Bxv26d/R4bDWANcefrSGgnUuVQ
xQS15rRPlUC+ukkvIP0RMbeGV1LBFGls30SicMuvXB9OUX8UAQgsDMS4UBNDWCnM
Enm2/IkY433Fxxwxcy9zRMJMp4X05QToEpPQ/zeVIPm5eqZT/6Ru+bcyGQEzz9FK
jsuyMm5LQALCas0ZrTC5Bs2nNujFrEU4ZVfZI3l6vHLiQ2KKher0XRgfwSr4/rnQ
y6Vhy04R/szIvGIyeOws4XVZeiTQ05F9/kJs95b8mV4jnOh02LNafkgzrB2mRKld
ghsiE7FQQzLlPM4jR0N8UwHHUn5MxI2VzA2RyZ7nYtzCt2KpLpkE5fh+ot8MAtyl
oHb37scw2taa9+3E4z4Zu4zUMMac9aok194A5zUxAJPWZTOR8ahz3dGTNHan4eYk
9O+6ZOMgJY3i5Hqw9/B891tiU7L2m0kc5xyLV6lWDskEGt0PxAAA+uViORPcs8im
jgnEC+tXNwDlE0WZB3v0e5fSh4wEM8PcL5GIsGtWjbQiccTawht3uM10G5PVyLHm
N4V6uBcmvOUy50iGeQgClzQn6BxAHaWBgZkB3wRB4b3TMxeZMFw8x5cPRHVUHIwz
gpBYIFuwhB1uDGVWdrDXlmghbBQrSTbe9LM2bntgRh/EsAsXbxJ+BSZ2Ww/4YE9N
qpJtr9ABqkMpQny5kU8FgabL25Nf4Op5/QZeiZjTK8sNHj4lPyy/f75NCdIRNyAt
8ltblzzD8q161O0X/HD6JC0EELFNM+ZSQtmmPpyA3CP7YU2rbya5teNAJLot1A/S
0mWdhMl9OLydxvF1HIJkmJl/g7AKSR9uwTqQXH2/zhhEZkQ7u5aKcg/ReIqGd6RV
Mx5dkV04VFAfVi1zvBFyzdasztuka6AcSF3Z5CYY69tV85pwzK7Uw78XOu/kZN/q
CtyBFyWgc2fyB5Af0MFJVt6eZ4TxYcc8inRmNNMPizQZ/huwJmPk7fz1ogjLQugK
8qTNcaA8qtMA2jwoqzq/xbHJVw6WWLrc3NOR/xKTLuN7T3hnYcjF5KeXuJmmoEZP
polizbxDyUdp+VBCklkTW/DTJAkm8SoPytveoU4wbs/rELxpBeufndGrjIpOc96t
99GI9CsRqmWQG9U2pNcy/1eSnrmOagDQ4mVfgF8TyR0Ip0jqQu2RbPsTqQ3veCZA
4yMsvHXwNBiv4s1rKPLmH4NStVm08DFAvDzA4KJsOKthPEy4gGODvdvPm/2Aw0+2
DvRow1thSwScct1PPJAKCoK1VmsiedX3cRQouLqmGVnqxuoGcVhPHP7DNrqnCS/l
S16244rdKBXtbYOjzJqHZB/8oyhInGHC1utCeryClGJzTMWUbdI3jCYXmRaNYajp
e+kgwCKrupzGYKEzFdMhAZPBO9BrClkhoUbXnx+V1thSfY6P6qmtu6kymb8IEnpk
ss3UDqHEoSWPgoGuV+RaJVVz5gWm447/SmGg0QFAuIAMZfMcGDKI6f6Vrh5sVDrc
33oyNKoINbIfAH9KrW7O7we3cE/YAeKcIhBD3ecSRXQVbYu0t1iZzfpTBTyjTNW0
C2CBEBBm7Y++fhLE07IEEbODOR6kP98LLZAhOmraYEAadnkW8B9avhlzf1mrSneS
1RlbU/fUQ4YsOge3pvXysbIZ/PYpVbFWsBumbMbSvYNLKMjbHJLZT3lJXns7HO24
FtIWV2st8NC/zWzyRpJ+LoffDXsTHlaRBcjeGdXNXOMq8ZyErplW0kB4k8LMtZr3
K5mXZSoi93NBv8A3DXViqg4JBMN1Faet18zBgpulCUG9OeaAbfkmrif3crT36nhy
oPbPKCvipF1iaLioHRVv3xHbMofrVKDy7cyenGYIVbMO/ZO805Nly/zTohQEi9Ry
28QPAakKX8sDHi6/rQU9gQFNj4bb5CWusn0aAA8zWiPxJuS2DXZJLkLZ+zpjfesY
A4h3Es6CxfMttlE4T532mvjkqZJOo0J1NKzTASjdvNa08i0mTcuDd5Af/yFtDoti
g61+ZEW73mmt2/7gC9OsDA+CeyQPiI4K3RDd7cWqs9QODDhcXr14Lm/UMQ893JXY
hMMBmjl+K/b9+I0rdzEm4aVtE3q/zI1qbXKKc8bkKJR/6UIsLFg0JbNz6P42dD1+
9Lw58ajg35lQxN13RWRQ8a0Yji8OX8psr2TkLg03dZE+mFMxFOKZMALZFb2zJxzr
OAYZddB4Od38tkr0OCNWLDyex+K1sHSU1F4eFSLQr7vOsR55w/0mYDSRptju2VOj
xFO2RZSEiBs0lNPo2IKUZBwbW4yskLzmjj9kqW6PRINHDYtaMonMbz7dzQMsT5SA
KJflGdm1WZ8g/eZYNafvh/x2fMQ8j8FY7kBy8CmoKO7hrjcsUkU3ZXfCRb7dCygu
RE02RDKocF6b9HgQ0aOKAwmY4VMviq6BbFPVKJyezRJE2/7E5OUPn+KuG/iER63x
tdRmKsXFLGO5W7mfyMv1m3U1Rm3uTg/X0dbO0JFtvtYJ/uQ0p6kQXaw2Ru1f58m0
dlu/AhoBY8wLfGDDFWughcDhyJR2gHQzKyTtbhkGqUIM4Ov90akjISz42lxCaZb6
ShrB5EbMIX2a3E6g98HrjV+pGv6Wa3HoYv22eOU6anIsGBSN2O3WjPamKeLzdqLu
SkqriICzIbh2DyQ41CDXnoBa/2uO9A0/0dGBRN9tYZcGtJWohcF7qo2z1EihbKds
3MYfmyxynjuFioqt1RQCDgaK8bh9//lE1Gs/BSg2iYt0NMLc7mjZ8fnMJOjykigR
x0A5KfXb8cFFHKsbC/4o/XqDZZXzOuqYoQc+wMyifn4eUc9SXyOdd2SgudkNg6aw
Q8zGzFXUtqpfsMVpiW5arLOuTIqO2FGpVEKfV5CCyEM+874tuy4IRrIHFDw3DV22
OegkZLVZZn5qilt9vJtXuAgoLZzTGR5iqbq5iMe7EmC2SGFFnuX3XOnXukW3zb9t
u2lCP0GN2MsxbRUHZrzF+crvIeBUGQCTqrIip/gaqKplNAbPMOh1FnakBOoVrTCu
8cCpJqeDy6ZTXRNsKrRmDvzJBuAhjFVqhT+RyFp8c2kf57bm4BbrVExSYmMbAxmt
NB0gKKsWcoGq0zR2nzoEivNfC8ILOlN0JrwH1ToCmO8p63GmvwenlRVYqKpArz4I
5HYOtnrJ25jZV4U4ljec50hsgkw8zomOHxUuBUUncpSIsP8BCGq/ZZ44PPgMENOx
SlYIbsS5xzmpjuii7ssXUzJnFQr4NNDfMlABtWWSCpmoTwmct8S0/B7ZkmbliDSj
8+u3QjS1y8Q76JoJORQy6sV7SK55JjdJj25TVIVURF7ihCx3fVYb85o0jHdQ24qU
/Hzi/BVT6rN/dAFNgJ6ed+9CwwxNyS3r9Yk/u5fAGsZNFvZfSMYBZxE4BuoELn9i
dXGxXH/Ix1Jl7JqVNVe9CKD5G8P2Hd3KsJAWY78CvWUwkuJ1keVcpksiFe+aQbGQ
lodY9BikBDC7esu6dfjqqYEGUWeBu+YrTFO1BD1VaQ0N93vP3AWFmFPpPHocBxNZ
Q83Sp3/vFjV8BRRRzNcWamPIuVQzqY+kV2oeouIVJ4Uuy8dq2NHYePpHU57Zusau
5++ZtjSe6YW5viLctRfGQxcJzrOX+hg1H4LF2SYFeqjvbnhHNitP/zy+ivSRL3hA
YYCoLCjGOh9w+Osn4+/+EGDnbQW2LyXMZwaRbzAtkFzPMaOI3G0jtbPYjj9SiX1m
QKEFIm9SNkFBAsHQM27ZnnX69vkZ1D8Nr6M/zlAyrmZNZQrDB4OswRsojgKd3cVi
VqCSYMSOaZgfOnpFGORL10ozZxFaSB9SD4VkaYWWn6vkNCu9vqy+MMe9OfGLFCHY
Qpypyu+j+yPBJMK5bXEYLek9idB4ekMRGpplXxVrFwSxk+TJvY+ed+okaIBOzNc4
8yIaZKkMtIPe26sFCD9yV/kv6Ir2E8zaEjaPSulhL3ce3J2k7fB3Ffoy/v5LA9i3
x6GAFyLSrBKz2O9M3FbLzWmyAn9ViFbYOOEnVJIaqRjY7EvWjsn9s+C2FGn3i2H/
BWzMtWOMyour+lUB8lUWVJFWrEXjyk/cVudoOLjcUTV0yM6o2MXGL/jBey2TuC7M
MtN6FPoU9GuJn5n2oLnTOGhtgFR1TsCQVzgdB7f0eDElDnZdE6Pn8P8tIanLXAY1
c64FVsF93o12+jqgfmk1NcjQVKAO/dogVlNlmJtUcie0X9tbv/jSF6WtTt+/JGdB
pz6VWbC2o3tZImfiTpyOKyCHadQYfARQ5uYMIekoYd1S3MlVmStQc7RZgoOYIY3T
uLMi89H9meGo5aNXIsqNSid0S7ULt/G+j+1WMkklht5Jqgmbnz3BVnQ204lpkcGj
8DGDSK3zKsn99khdwtQEufUTea2Ojmxx1Ji13RQWv8MeCLuuZ4q+/hJJ6ZuNv9r5
GxycJgtD8BlRw1T8jLY3N3SvtuN1OJgH+LvktndTOSwiNfb7BsZEQqgrioDcnxi7
z24NLRXxNylseYZLi6MyYB5rnm8bCrVa28DizQZYpZv1QpgPxSV1CYP5zyo8sC2d
2ooal63Bq+q51YvVDBKvXTOGvcaeW+gMTtQ0g7/oOnnj5kzI0bP1XgZZAOdXzi/v
wA8DDk81XY5qwYkuO8INHKyJmjYC9lOKiqJuWejmZhttg8W7cneHmV67SS5d5hRd
+SSVT2mCCVq/HEmNrjRP/3ojfZu9YNJ/Jr29Q338nbAgh90dxbNXd6ke6YtQiwoz
J6apE0FiV76nDw0B5oEGX7d+tcg+E69tMbl+CJYRdnxt+iZ1JyxiJi+qruDRRUUw
w7CdvZh4zsphkWpEPAA6JOcTct9IYq3SLMMr1/YNdN75bu8H+2FpOmP3t8xxENo4
/xF+n63BL7gyHYUS/H+8S2cqclGOxMGNvCA8WEZe3E+gOhZNR8VLfS6B0pinu06b
pKLoOgrz6WLlQMEvzok4nkFvLxqknbvAn64eG/+SkpUYtdri0uJvocN+sKrlU/2p
GrRLkjiVfnOb026SgKB4cfem1kU6/4bg6l9Jnf0qD/AQMc3b8NkScSJI2HtPPYYE
5W6gqgjvUnyTEgZ0OfcEgXnKxLSN6wvkK2KYdmiXOpGraGVa9gVb3Lobm41Kntia
trZpMFDh8N2tyg5EuKciPbym2rnqIJAQWCZ8+ttCiKGdh7MnBgIPJ5L2y+VEQYyY
VfNrcmzIxcErhgx2O9KxmgrtzE9xHUuIR63KFZNvFwWEMMV2IgNmFAYcrSeTfrR/
2N/c2AzHRP5cceWodDTBRtd35te54gDg5ljUnhMpfAcdhQ6R317Nom9Nl4xSv7GQ
p+a7bSB/PW9tFWuMQcbcVKVuEHz3yk+LekBFGGLGZmmULiAQ9Ge50uPPVz9UOwKH
L0/4cZodnwiD6I6mVJj+xzfdWvnvZd1YTt07ZJ6ZdXdrBauYybrLjAdfzkAN7ggV
hJRoLQp2J/P6lXvCWccDIMN440Gej1M9hBa7RBMcduy7vFmyd1gg2/LJMOJsUEmb
Ik3uDWzaWoXWd8BueV1H1JklnDLbYcHl6INdgQYVXCrZjonGX0ebgg4CqHrXEWXn
VsuNspt+cl0uCK9xmPQZjSBlU538bOldDtFJdkD9k30dsCt1VZt2dmG53jjndd7u
2ghK9xy5ab9BQXt/KFXa/D+Mc854yRtCGRmbd0Cpn644FJ4Zfgl30kKxlgbW23+v
Vc8PHZKj1lBDaKpQtelMqz5V8GQeifbIf5sNJ+T9MhfLcXbSQasPhYlQwVMxTXJV
8HezX9TSV6fiW4VROy8yuySqIHjvUWdOjVBqldVo2LsYil4kD6q+s0nhAMRa8m4k
X7YIz8UYKjrspXkw7oX612QnmLcJGJlCa4FhHLbZoI8171ujHtek50TDpPb2r/8d
4egH9BGr9zygjPyS92ApBh06R2lSOJuXmUY2X4Hu8G0PDm1VvjfX/WtNvNJLEF19
exn49giivFTYiIsDLCNsmkteOBlS/lnFnkhHZPSfvb6wm4QSI2F50UN9F0mdm9yq
wS8ZVWrxAfeFWvcadRKE06aOHd1DkzPKASS1vQ2uvL0QrG8EMNo/JV371O53WC/E
qjlDP3IUQdmuxTZ64/GohVP5itlbZYnasZASWcLoKSqcVKdoJuglFQaJyaKedAmw
5q7znEm/Jo/OMVxtlSkkz95vAK0koKt2hZFpPq7K6ds/WmrdAmJZPdi79eRhLweO
y8JCI/SlgZPVruADqIfvs+CDbuxiE7hyRx10X+nGjh7yeXupOvi97CUudljuEdnZ
NYN2rA8Wvyjfop1Xn5I9XUcyRTcFJltQZKaAhOg4b/JP18oHTpOh2DqXYbyO8EK/
+eIRu2gMoadrqS+DZ8btqpPEWZxgkem0qUwCJfD8wHBHHyRTribmoxn+Hsz0sizI
eGGKlvVv7njZhTPspMJyZLJ3Fj7chtwt9A9aFh8A0YyzCHZltzAQ+2y8cl0OhjCZ
95nOurTxy+/CPu7+KsxfMi///yVG1KNuyhAxJpVoANyQU1vnE/nSxITOrXwtfMpq
zlSFw5WDKcpsObolFq4zpmlVPCjOubqTwVar3uG1THTzIWy44z0ZTHVhGqY69v1P
VBMa7Y36MEoXU5FnbvVaOhCvTya4UymfBJaxQY1v6rPsbZ1oO10V/fBo5+8FEW8q
2j5h/1m2+gfhGt1gvC5HuGxDNqEaSFHgWp7H7vvFp6CPhjrGfgOO5Tc3gyN0LuqA
sw28vC0EALLFNc3J7eMRAMim+PU5CalnBWagcxRIsm18uz9XKrxlD8iIuDX9HeRL
3u8vlrk3HfDYeD5ffEFv1RLZO4TB5FoU27vAhU+vg5h+RVCKkxbG0SQFO4DplYcp
LK5HFKkW/fGe7a7yb2EKEO8WWjGEySDbbt0ckz1iuYODfWBwLhL7fTYFCYiYgbtH
Yzenn40U3oFHaQZNWsq77/SooNfuYXXrV4QJ26ttP05sg0uekvZ7njw8yZlE1RPC
5ZEP7GgV1o+nGs75VYi/WbuLcnwqruDUgc3ZfMS64qeV3Dz15eJzKCqErPFxrhZO
bkyCe80jasVsg3L/wWnA1EOkzgXx6iQzgcebCAcRllDSnBOOY7r7d7KR1Tias1mF
2HWACOiT76RsFIVc3tPVkC83UrCvDmeeX5xj1HLzMyC/+Is7I8QSCjbwA81DXPyv
PU2E7RpcOHlFqNZAJ6hZP8HAlHiUsY6U2kH3wpogLHmjN7RlqO/zxdvAgGwN4RpG
8UMfIs+TDgJPSLSJlE0uV2J90bqfy3r7GzT5M67BSAy2toaD9ukUjftWiLujnd8c
WlvDNFCfu28EvZivgY981Yg7bzfqbT3TL5RQg2iOYbENuu62ToCzaXRKec0205sq
Zf1RVDUtD6RYW6bXJaOmBpPfjCxNhKwPvpHFqrR1Vcd/+ycIK7vM2rdBLbOqOFn9
e46m6TSBAaBRRut7bTrnTuaqK92nJLLqo4yqCFe9MG2F5LxW3efQVDvSium+ClDt
1IVGbff1xS6MXtD4Hc1mUKzw9K1ly6busFs35ml40I1pfOx8zqXN2+KRgHUQPxT7
vM7t2wm5magiaeE4PJOzduY6Fr2utQ7T4Zgpe9oNU1/YfB2AneMPrw64722uh0YF
rolf571ReBiEDb7YfeuHzJG/NmPqHNGDwSqzdlcC6ExzGSQJYkTpJ2C0OTQYbqTh
SUlynBJJqmmAPaMUEvcEQdOfpOVTrc9vR3iDY5aGAYW1A8nO06YEvD73xYNnL1to
LHcgmevvMuMl0ef0nOAxMcL3FBRhYOfcRB6L6r3eNkqb3Xjay0wgC1JbfC8m+F/2
pQRzKou3+VAV0xYfXU89hy+pCtJ5cdhYAA37LEXT7G9AmKYZL0Wb34xueN6hbwwd
9Qk7v3jYwU3PAeZv0OL2nqPD8TL01x08lTjmrCeOaDpm0GEIGgsgU9mY+IeZ32HU
FOPCPC44ytJzwxQMjynF+UFNeCQBEdTKFkvG8A+2KGeOESGunXBKXUH9O8qxNhey
sAQQjPglyvgvVu51nLljZYDZQohhtxu+rTsuWNeHIUij62i4HRaafx8gk+tjbdAP
TQvn/MeAZMaFQVI7p721hGd7w9mMVh9yEvIpl49yXOH5qpLYUrH8YfXzwZhIFtHm
971aeXXdbaAhcq4RGqqq/3w9hCeyPpFcDk542gJ1K6AZ2mhyk5Se3ZcVDvoEEFP8
xPmsg0lVbf5I3SzS1+/23VxLs8IxGYVPAUwTdj/BeTs+lgdR1ocMhDhoRddwfyPL
WpXZBZk+G/b6RX5YFecBMKqXXh/MIqU6s6vfMuWKdgVMCWXz/IJAyzzniSiEJtQT
ghCHtC2bkdrhK1ct4pQyhdlLX00MGZqo8D/qyRhXiA5xj3+f6oB9f47cZzG7tDeb
6/iLo02KDYiboNwpLdJ57SxY0fd5usJtCa8SDu38aAR4+8KsE7R8N5yUQM4t02Ib
oOw+y0Ne4gx2fphDtbF2MA3hikL4VR5wVomeOea43a3AT4oGQpZyt0RSIfs3KN+3
9t9+AYUgbmZnLKiZkvO8JOLuRZ/Xa5V/OlsJiPWi8eGY13BUdmztAZ7L5dKdZPfu
PC3kJElSWYHWCXU7i/Svn3GSjm0bU4Ha1Nf4TTcHTUnSbBiQc9hXruiq0u2u9oLp
OCu+8olejwdOeGKdGUmm1T++6dp7tumyjtgmx1I7q1WnqpUrMuJIZuAnfs1eSSTK
auEWKVfecZecAqIRk+73m7nwaiTEGUFHmBQJou1xApAXIXDi5a53qf2viCCFEFfh
n/pv8fljTyn1vFAwcb5lrGwKMG4jYagmPOFT0h3eJEe7k2y+AsKZ1cGuTLzHobHW
YeI+Zh+DDdJw5zj9zZZPqWuXTQOZUYKvI7FmX6fG2lVAYPsGY/dlBdjrx79uv7zQ
Ty4C6KQ3VbPAwp0UhbgRQp41/W6gSrbCOWl4asOKKisYGW/K5MCegvxOQNOognck
m9WZS3rtM/mBRs5AITHWkB/aKnnueRAWlMPbnLfZ5foR8p5RKXY1efp1yOzEMsJg
n3Tw5WELvm+POEt/yiepF0TFDwvQzQQN0OGoW9not1RZT4C9DIaIU0Hyo8owEvek
XDIeaqrfFTtlFOvvHo+dIBKlaQtcFlJMLLiJzLvNreya2dtruwqWXyFpXTnZPhdF
Kqe+vs31RU3IfqQ7AWGv/6yw8qg8AvpYVKiXvIG2lgGDbKex3FO/sFnlSq+2J6N+
+1VEdIp9AFczR8/kQ4wLEQoK8f+sPxZCJ9dts/tMLfj/O775BPmu9A6RG/88VdCK
UPxEO8If9kgiSQnL3MZWICK/lh/ETZnIcpqKMw2jnYfU2MuLaI0AFBRMzoIqdqpI
Nl5EQF0ipDwzN92vubePJEmzSdgrmXbMMuDHHfuXdNEVEDDcTWdk1ekC1rHahaxw
xSnuQi5H6dqMQI6BNmaS+u3ywhgBIFoorI4lpVVR/cKYdvum+9jlllrvBYHbDYvv
V5UUXyYhmfGBBKzmy8a+JIU49URdCJbuvXRnecRCaXvC6+gdIt5TDf/z+GXcSJ0g
/ZUiMJ3R9Mem8+CbZz3Tc9rQvgYEdtBuG/FaiIRJLsVyTpqsx8LWPXzgUgOq57OV
yPHOTUciQeVS49yF71kQd7nX6+C5+kJvRhtssTd1me/VLDkp433tQYxVQ2HOJm4z
fukiNoiExqtL405+Ff47tAeu/HYpWdsvlKUIBWLmNUkEWAbgXddsdPHsJuelu3YF
61juabwDzQceeKtXWEHA63BTvpg3dHC93boIj/0rSiZf7ZK/S+caLcBpRBTcmBJo
TAEJcTSk1lYg8lDqw4iquaFZQ8c86QfM0s/+JfLqx1sN//hh6/j7xtZvXTHPZ+ob
i0Z69pqwUP+2DAtwysJnh2YNYoYXaJknQq39qJL4+Y32K3VnVRD5iU+pq2jJhXi6
Bmpbv4t8ArQlYAXs5FHMbtUoAvR8bhM7wC/RASMTvA0p2e1y39KuK3Ah/SPUJy2c
qhZzDIH3zF4hpuCh/UEWJd/yDSR+U3VtT7Wl+o8xH91S/+Zql2lSJpXJHvAVRWRv
DaKojwgPLAItRIdwC497zI7hmU9g6WvhXK3ADzPpBPseW1h0+XW+oDbz8wn/HJ2q
sXdMEKcYfcQh/fmN5CCv6WU5GXIEZv6a5S4lIKgOM7YCB1U947Y04lUv7/y/H5Zc
4GQL2SXjo5HdXB9T7q6g1XLAHMxy4U8frmeOq34eQ/Bak+gJwBSB9z1bzmys3kF5
PRYdfZalSlIylysrJvom8QSUW5XGLDTmJvHSreGB7kQYom35qnOIW2wzJeAi+7HQ
/0JNqoXVJw8oEI6uHo6gI9dL5xIYVTuk+obQE1jbn7karUVw8RgtO1SVrXFERvk+
do+xC7b8JaEsL1QGXsPwN5mHkRFWSZAVZZcjArgmjKIBnaMPu5i9UzzVrOcoOiss
PMunAlSVXWeP87QCc9Okd+WI+xdPHx4cy+C/cgeUAk4dDz/1BVTtVZ8Sc9PhUcvU
BaVAfOM70079AvTAPrL2FabDA9nuPkD83CulPnsabfn9AbkQEzsWHC5UUCBpTLBC
MF10aolFQ25zlbJm84GGSQLF57xwC3l9i6UEZjOr56eit4Bj6qkFF1cccFyo/fvs
K4BWTBRY/+vMzGug8pWM8GlObn4gZBl0SqVkomZf8fLbN8r+ZuNtGrzAZPGxfMbI
xbpY54dIFLP8q9+RSGgEIgydoKFNFhrHY/Cc90Pk5CHkhmwzisRh3BpIxsRaA9ew
+sJX6iy9tX20BgOh+dn7K1K/Op8CNF1GWsypdZJDFW3X2/P8Y2vpAhNNiY9sKQp5
1nZq3u1Lr4yc05WHrckxeJU23PnLhrvdUmpsoeC0WHoA5b0MZFiLvLOe7KxGKogO
DP8yTXUZe7IigWAQYlPvfce//6COQJ23aICE3tv2qFBFMz6nj91PW7cspMyAB3go
XBnbOzmRLzAlWpvtWafE++ZbR4JDJyQZBGF7/+tbOBXemISN8oovMTCEvXPuCIyu
8FUlasY8RHYHXc5h9Gqe9kdZ0NH1Sjp3ChUesSsA3oXIqUngfcG4Sz1ba6IgFYqD
W+IjCvEJ5KRsGP0Bo37incuifj0sYi1Lm56WkmJDZk73k09J+0MRiPG0YBYThL50
w2M1CPAP+c4GaRgn51svr1HuztCFAoATntZcGgbO6ZgoOLw0IlFr21LRZEvABfrX
jrGJGpeyomOJdC3QRFZ1cpebJ0+4975SKC4R4/xERXLzFoBbcTNt9jByjE4GXXtc
dJH7DDYK4KFDZDu4T+C9uL3MOvsc3uLmb0dT/jKsTl0b3IjhjDeCjuh72bNVHJQ5
g1GUJsD6++HVGtAZMtmibvUSO2+NLuxTtX/J7WuH0JWWpJ2yQpKwIAKXwzfH1AlT
ZhHKHbEDjkC6BJ/N7O0loHge6qoP2+hMgFHt8Nvm11f5zj2Vg08V9AtXXLA5TNfB
RnyetSNIrDc0o9y1YvT0DWYcv99Cnr3yskRC20IuIUsWlMMIl6PWgwYeB0YdpFHE
p669i3iSWKiJNNTtuNRGEoK3nF2ooVQuDUe4Q/W+qaGvckIaZIO8fZiFVaOXOt1e
UwOaWPkfTNoNkavVLSLX861kUgmaayAPd2jSzu3yP3htceRPe7iLIZx+lJxxRAJ1
hcIZGCt17wg7YUPiqcI9JXKJHStLFBO8wDLvOsH5/hWf/URAg1MGYA6O62TcId4l
Q924632JI1rRG0QTSLiz0A/lW6Qx6G/4QvGCGvB49ovhCmsisR8lBr8JlOkDsQa3
0AK5ekijKXacdz5XeodsOQv5TJPRii3qElQWJyczzfvpa7TISUB30pMn1VlAtnm4
WQFA9liV8jTLrlLMZCwGSklrxv2XQuc1KkzN8hWWJYP+/jHeS1zL9IIlsAmExjZl
m/xYvQvXfDp3AOXSoMmnWt1eKM4vzydb7eYX7MdaWUyKuqpIAuEcCRbi/Id7vk48
fBAEuD2UjYcTNtwGmUVXwGWXH/rGonfb0TSYhojJnf0j8+aduXRc8O1dfLCS+XZ/
kROuOCk/9+kFTQbQ8H1zEgf8FoKba8J9n9v8GYzTE9qS7I5i4QPi7bgFEjOBu9SM
qsBTZAk57felaJAH2OlcCQzTjRuIo5n30nJ1Jlza2WpZXJbnIirv8PKf3AVYU7wZ
nDXPbStdiyyjIkFWonRnyV3OPT4IqSJFCb+dVFYKbKMBhqhYbEX1oredQPmLfahI
LBjf18ji6YM/0/Ue96VOK4x3frrDWA2p25Oh6X06S1c/IUrCpTC/D1fkQi3Z4bul
PZsUepba5vATHf+cNUWP4k4oGHTnKUNUPjsIpEZx0izqd3uL4A7wO3TyUfeo0Nd2
GVduYsB7PZuUW6vc+dEnMQvzGie/fxypbiCVxh3Ox5KMe1DQZ8h01pe/aDJ+kidJ
vqS+4/pKYaUtpwF2+5mOFxGc9L0YyX4TbwgPmtsmIvHDraBSztQLcxLsy+qjSSeH
4G9q2M3kQK/Ns5tMEttR1Vincho+RP9cnme3jGJxF3up5dkpUYHlc8ix95gvSUPN
LVf0ddUKYHrVBHChhgtAMVH20rq7Tn1cSuKSoZ3K0T5RIzfaHJA7yyjkdBQo3kHK
OYZUUywx1Myg38tt0gqy1ziiKiJhQH+DJKmzAJxoajMLVbfUHVcGCmDL7/ofsbtB
wk7JQBMIPhpV9e2aEn0hklWMddSl/esXih6HJ16Z6A4XkbDO2MKLnFiifCTYvd/L
HPgBNZq03PoSjyE6TEgtfHmIWlmqv1+I2u5bTCwfSJcFpS9uFQoOOtXX+ZH3nllH
CmvydbvHuwtAGb+L5oGmbZwYu/tCepxqerkw7dHrXFxRP0BNRfTlU9byAKNWm1n7
1TsMXvPj19Dcm7W4dbk19f33Dt98ia+IIK4OTgwSwF0j3Svk7k7Q7BPBzhXeU3Qd
aKpeCWUTtFhOaxU6tgaXbZFj9Ieujds3WraeCez064fmeoy6b2l/LjRYWZTUx/NQ
JIa+Kep8IPcRxjm5T6E21YVN99opsQvsIMELRB8E1dq/0XfT6liK8ATO+ro9+yju
r3FOi1akd4J+UPzbFU0BdxoPkQ+nieAjd0L/qtRkQ36vk2s7BMv14gZPFenTrVJE
/vMm2txFipULjoRhKfD1KQB3HD8Np/rha5QO35VIAqLzu9QBn4TQRa1cX4u1gwrE
WgHcfXlrEFa2DitA7oFjX5GZoTvqYt31xjCXL7WGaddYTsIt9gfSarJDzuupg5yE
57a+ISjTkMwzKz5iA0QfPhgJ2bIsKp3dZATWRB/pgi7L8gLaMGxnk4LLk+KG2IJR
wPtlYDJBCOaDYx2VfaXUd68RbvnkRBA0mbOGUIo3aXHH4UCULY20LZv3lsvswUCw
3RUdlSJMB7Zcv794IF8pAzXyyzo5qbaXaXTEwS0yrYCj3+ofGCi5e/4vIeKwKnm9
nXoyw3c+JjI2AARkEfbYX9j6/cfp4Hfv7ePrARpd50Gv0Zo9qirVo/6wXXyjXqmd
xUzVVVwU4jYn3/067997kBGRaFCu52MVgJtukKVpsCyWikq0hcNGlIak/4an3Pku
uLKROVI6EHJ5hYi+CIe3xDktMvA/I3Mw0QBG0r61eM53szlrO/CUuItoZig4kcS/
fRKu0XXasV57VB1fO53oeIKBdgbDqrY49XyuigAPY0mLkfCcDcE/HZDYtD+Fo8SG
FwBjDcD/RS254EnLM6aOND2A17ksal1b2wWXv0UnRGYO8Ah+mDOW9N6yRlg8GWSw
5HXbQfNsASMUG/gdg/tst6FEG0NxHKmeyMGiz/A+D0XBHXWevw2LKtJCEF2KZ4ZA
vdmxhg8JTr8n4NVkga3x0yE0N1+H2wpmELohMNZCDXN/zAp4TrLXUano7C8Nl8dS
C83OHPgbZKW5/ScwFEl23TUrGIJ5JF+BpgZg0OtJFpyJDtmGnKa5/ixdidnzmx0A
jiWK5iEz975lPC6ewBwg3vx1u7fgjYSqxV0wXkSfOASWoxy7wUfWpbgT+sieMhq8
Fv9g5QiDcbhOhzeYDlH+kzYyPeQvhrVekhuRArCry+zyl830U71fAuUIdVDwmEB1
3+8F+IaFNWbPMnkXsesOc/1mItXvws8wSXbw9sLxRzk5EvilygOPN4cftLNOYkZw
THacrGArBWYqruralCuvVMhLgbwswFcTdrI+kfTSOmzistMu0VCjtGm40y5WHUB4
aTDGM1TGKdNaLpESYQ4R2hqFVqL9l4uSgkvrkrH0FXMCF56JqiOEmEh/pIOxhz7d
kkFYIuMO7mKWTy/6mrnARt72M0qjwE/7+JH6BM4sP6fefElDkz1Q+YO9dIDmjUWg
K5ctDCrsQnM+dlig5l7/r6LVWPqoXhsGKCKzAHfrQ/ZoaG4bxvs27/V/25soDTKB
4PLpDfZS1xgqi4J1uOb87FiCgOwH6Efw6eVk131lyMHYL1l2SdnD+x5lnhymmGXc
Ke/T9wUhSUQb0e6mUKqP7hsmB8my0tls56Tr7aIkVTXmVSDaLrqsy2Tz3NvrEZVZ
8OkiPVFXLFysQMjZer1AFW8VkkR2Q4hjNZvWMJmn8jkUAnI9bpHgmV3LSs/NALjN
FJCvmulr1L1E+ABKzDZEgYJ3gfJr+0eRtHVECvC1Sn+l58VbpuaoDrvkb1lUGskl
PDffGCsd2EuUF3itKD7PQuKqvFjWrZVwrfByVgDdO1sTi70ZK4h6Gwgu8ovI9stB
XhzZmYhwE/6MRe5FwUDmH9zjXUQwPDHcI/Lweh7DrkCBmqs5TAncAIGyWshVlphd
jh/YhwGXTbjFIoFkI/084WmzdwuxRSVdYstXBPD4GusqI5kw0RucGyb/y3rtrqZE
B90PUeC3K+p6HFyWNBwB7SkzSSGDPiDoS63rHvDnCEpqu/Gb9WLJnrl6TuVOCWp3
q5pG8/EofD2nYUiechDfU5yJfVx4NFWivjZytckYwqyvqozB24FeK3H3LgXAhMYT
lZgLviuoUcbJC/KbOJDf4Y3oK+pzLYer6Fe3Zotb1eXBJMuglcvLlhb4h/b1vzmD
uVXU5v15ho0ocXTYfkY7oMqb669GRwHQGsPxAeCGYZ+xXP8ExO/0CmIyR/aozcFu
biyvyzh6sCiI8j5KZtW6n66EO3rTv70RMiGNnPAXH+nLDGefhmcKIcDPp0ZnlrEz
sG8fWdw87T31699SDk2GBNSGm5JGWa+Xgf0YmpXgEihPBlMzHelTssxjm9UrMfKK
nM8GenFth+aVs8uNS6hYOAXdibivS4Lom1ZeuH3+qMO2VUIDRAa52XhZQqtlmKhX
x+bkMzBT4L90LrJ+riTj9F1+9izN0BPulvO6QUs5U/qrJrVeDE7fCoOHksy0qxg7
9L6Tid+50oWN6lwgEbkCMhpdKNxi/PNJ38DbuAHtovmrJsbJFQHdN0j3gnxeeIXv
gto777YiS26iGwYX/yeZTkYeRu1TPJcLdKKYMAgxHGXbgh4Ety9pCMWpnTIb4zEs
TvhTrvARmoqrK+FJF0s2HHc0yhAEHf3eIM2rHswrqE+kjUWUN6VZtSOaLZ7+ZUME
/3YnKTDZtTIHHt2UYqKo8g50J5WI9nIbHQ93GQkRrT5NJ5eqgHj02I8QVhx5AY5e
a8kw5TrmEKX/Mhis4ym6oUbVqOi1+lvdt5MSggpJ84FKmx9kbhTKEOT7UTMGFNbw
e/qu31+YHkwIIA29YjLyg1eIoCIs13i3BjezC21J5J6o4AyWOYbGJra176Rp6xfX
3i2vyIh4DaXWxYAghc+L8CR0lOBgka2qUNX4UTRPqzVs57mjKceV5Ebjz80h66i6
3b8VZUFsaF9VaLKxwY0p8MnZlv2M3kauFv4LGv4rbqQxEbjvOKg4tPdlRjRdwqxA
Q0qweshWl04bEgo2Nm/7adsaW9exclwjx/TbJ7iessebPaH4wXsnDFmtCieySbgX
aGh52cgLnbblW+biLGz7FvcEw6+g/FEpj27ScGCDbuPBCLnI4k/qBoEst1ZfTiSN
HneNVyaHOJOo7l97L78jUpfVzbCGquOJ6+WvRqepi9OxxJMjrV5ejbE7v/a2UjPU
hC2OgUokjLdc6GAmugDD6BxECb8Rhi9jSATAwhBEnta4DPUhIQPeHrv1J+ODxLTE
pMv0q+WxwKbLD0j/v/vNnP8TAJ0q4PPFyURP++Z2YEC7LoPAtimKqvJkP/GFyuCU
wed3qxCJoil53nVRJKeIYv3WktxZ16uLQRm5CsD+c5+LJO5YHqVeWFTIEhyLaylK
HA7350q6XXvx4m3FLaSpvbJogjQicSJfVQ/gQg1CAxU/2uiyTGyic135EfGSIiA4
tnL8wLs8/kTwdyk89FAibh4Hb2nMjLvh3XTd6grWBcDkgtdM1JXS+04shiiS0UAS
O6aQeriSAN78BjJYOZ9k9qI6TtRqNNlu89s+2kpT6JTZwVV5OBpJwNKtrxMKgCsS
X/52jGS2lnPP3dArjvhy0DNPa1oDBc5848x3lk9gxczq9IxMondomc39/GaeRaaj
jD/TQBhs6jXNwpRIB3Abl2AnE17dsQoqIbAKUVSa9FXs2AUF8d66HVnC4fNC3t8i
PsUR3D+Olgsi1IQ19F9VLWbzh4fXonRwa/5bBFKLxSv0k/tcuhYQWMUlmFZ1FRzk
RdXIsJn3i0CNDUYmIfJY5ZoJyU3ZlVKtKaXxdyVlSHD9nQfHBX8y2oPEi6OEFNIq
NNaj/bxUoCna8KNl9qhzMdMD1U/XqTnPKl5pskxMIeQOYweSW4875cDHpA/xG94J
zEMuF+dTNPqvqHhs7vzKz3IhHjWdmMILcR9N415z0oMp6EAma9Jknh1WEyvEjS2B
GFVMBjVA9tpe77qa98lr4xrzDb9tsXkSslRqsS1mIU08jUFTbM467bHpuFaeEeeU
X6e3zfaWulx4lRT1X09rT1eKUmGmlcJseFOH8dK1zbvZvHepv/falTONmymOG/Nx
Mj/5fYmRiSNJ9LWOl3MDF0E1cShAjqCWJBg5UErhG2kyaOULVxT0gzZ4qk+8uU0Q
AUBRPkLeeaSYzLmYKX9CTCNR6NG2PAGKt168tJklQU2KwF0OZbNvGAwuTjhMvSy2
pbmQi2UBnXZBD7lf6BspgCuBZgS0RcHIFRH56ZFf93sH8VTQc0nAR5K/MEg3k6Cn
rPbELFE3IoskCJiBhPdIheEbBoEYwXi9mPOWhO/r6tZ5QaEH6RFLuGV+L08BKTf1
Npjz4SRiHDUgQ1NmmdujwZ7nG94T1+iIqAk/9hqK1u3RyJ7oHCGXkjdL5+0PmEi1
WFZzyhVEm44vu1tufNQV8wW3mZzsYGeU0XiFJI3ex24iSMR59NhuAaQ2JLKO52pj
GKLFyzwt7DbZ9KiYYWVxWJ877K47CBoft3oKw6Gg+mBeOLHUSkiKbKmZLa4xXDRb
9DgZNCPZin8vR/fj7Bntmi1+x9UF89WyHYqjErv/VlhMyrLmsS/3TomNfaqWIht6
ThQ3DaNzaLX4VhFTO0BW0FCRLDbUZ7hU3sm9l0VkeL623rMoRYuE8k7VB1Xs0u/O
WNAJK8tXCCW61D4iVmaFgSCbI+WQtR78vQhXz3aPMZkfo9Wm1m6J0O+kP/ilE2gY
lEqU2w+wIHiJl76YNfc5BTbAMRlSTdfcjot/SlJgempldYW0EIJnQEyHvwIuE8/n
XinLMcdNnZOdxIRHNAYp+M0t70P4jXCZnhEXSOCbrlUdMpKZnKpqEOjKR75UBb4q
C6rjRiwR1iCEReIITH0j8aDVJjxvuVJ8KYZ5LFvtggT9TSy2i6qWhQF0cpapat6T
h32//OFlI/sNTp7T/AtT2QmM64TSQpPB/rSol1shqGtJOtEs294XbU4+QV/1/OJ9
z9OarrOi0DgQesw1HtYt768oX8TkjEzJNfYVNx4s7vqDF38d9nNRynTRb2seG6+c
ppie2tPLevfL6qlJEUoONXZYVi+jZzN1ZD5ISgCDF0jo55ACo/mxih8gFMv8l+48
pUc0Sw9ZxmgIypmOQRv972vGwZzCC3/P/E2d3av7NHSF4Z2XtH3dkPg8Kardas2J
2zptiAru2+174f3HZyZ8LlUx3SEnoIjzQshzAIsJgowE8rMOefBdc+v519ue08zQ
IiR46/+LTICJTYIiBI6MbzQ+WU9n4F5alxZmAZSJS6FvXTweU8jCjSL7w568bmfM
HKuCXnpjZXzBGqoXwmW5IoIMQlL++emgC0L6iqq3xLBmMGD6lJoz2Vnq8zXS+nZY
SkiEUV+EG2tRjFsqnFz+WLbpOjCswSUhfIYh7iid2n63tpPG/ModJCpz8iVQem53
5kKDCnzeRe+Fpp9wqG7lRSt04eVf+wBLG2JhmsVGdkHT0YcwXAF7inxAurkwCPPB
AxTgLZbdsTB10j6q0sCYNnw+c3UCBFkTmEZ3EadqrbVmDALjABRZyOhV7OXBR7Vv
OsZion7y7r28zYbrQAedZrI9xUWl4iPm9sFsJluNWqgr4QLQYzAfGKeEaURp6uoj
GlreMirpVt9wOiRhH12svW8Hc88Nec62iHTI49VGTJ4wV72R3K/j6FFWPt4xY1nr
+0fEO63+P0wZbfunIc3SeYSx2SVUF7SIb1j0tjaGL6Hp3Pd0jchjxKAs+AQ8CRo0
T/VDUWpVFsZfHbB45uG1S+fnNyqHNa7KbeOYSbxdiOOYOl1lCreulWdjpm0ZpJMR
9oFQAktas4wJ2GP7IjLdtbJVw8w/Aeyx4ZNqu3waxQSe9SGE2FO0f76JqSHTtetO
hjR23X9ElKWDmB/4h7zILgOwbV/YjZQNZPdcA4gS8y2tE487WKtHc2KIsQTIP8LN
kgCUzOS3hK/lb265zBUevG/GCIQ3k7ewrFmcVrIi2jbEBLIR2Y7zgRPtra4X+H/R
N2vF5RdSxUAZ+52guQzZa/zn+GhV96HDUl3+90sl6CAZmdelg6+zPsAZ0Cp0zPqW
6SaXd15YMWT/WCCrgPhQu9wmdqz0VEeinoUJzcjN8yR3hJtl3mqS1XOkZNc5HIqm
v9i25tYv9LKcGzsi0y96phmiDfxm9a/XTLMVO24M2LbMXVV1eHHsTka9c1snvXmg
m5+l9xSJLaHUyQqpIIn1MMXJxRDnGCILQYncRrJqEwGwgsmhwABCpd0cDr3epM00
EiOR+qVqS3QPAxzMctGHP8I1WosIwC2wZvR4CGyWkWpsFdEgSYk4Uoi50rhlHKJb
uun4JZWll6DmUtGqoQerXJopisSvikxhbK7N/J1fFkIck/qneTF2QbgEPZMwAQUz
bjnyVG2+bq1wA1e43sFxfRLBsA9BPnZIyU7wHVQRdW68mwGLdSMmLQuhlG6OGwDu
DyoqHTUhPSJ7kamPBx5yJoY4hWbJEndTW9xCEwgwDPzlvKuG2s/VbqHl/0gt8u8b
6uMJ7j+v9zNnH4SrRVk+17EttpaGrE6l6Ed+srdYaMuyyqjwPkS96tgPXQ0AR6AH
7zAbyA0rQxZ4OtNnpElvMvacJnhIvnWo+R8vTshPbgI+Re9L7K7QNKAWljN4M37M
BASFFWprnSmGiseyg1Ahal8kvE/4BPoAjkU8JM0oLkKplg3smmGAtqpz7kDpt9rJ
FxB4G6THWlJ/qLliIeHqqdXPoj+Uh+RBIaMBBVuzSByGDfvyY2bzI9y8vMpMfSfy
2b1mpDqEknlI5Nc751aZrIUdCIK7FgKjcoskTbxxElSdx+rK3wWA9MTaUkANtn+e
AZNy01A+8ETUOfpnAzbHfCV8+raOu7m92+omf07YSEBxuAJ2bqtA2TA0OF1qS9Uu
tjGBiBMM5QhAETVjZv1ZR7daQl9EqyhUGQ2WsKDrbU4PY1tfYwgKPHYIiK63oNt8
w2qjpSp5M4D5QKQSwcnTOFLmaWRUqwOmFcZNWUnlLrvVikTkrloEQC+X0HgMhhSN
5nIgIgJAtzlrra9RVghaF3ljUH1XMDSG5cbusToalQwWksv8x5UlDrhw+OHjhSGh
u01rOceEM09j4Q2WQnXgeQArqLJpr5hVmTNEP0JmkyAiS83IaXGTvxz0lj8xTT9e
cefDbjJn4dZhWkbu10YYBmoDGebWQZUtJTmTJSPdyyJbv2Wz714Iru1UPR1zXWnp
xjhxSfIKe/vkK9LsQAqN/nshlbIO4ToQaJGP2Z0Vm4PsPjKYuHo4ZXfLdp/Fbucg
cq+gnW/R0KmhhUUS1KzMsASIDgDtBmV+nmlZYP6TW93J4NJKD6sXe0ElKU6jQtcQ
byWFc+syKUwrsZmeqxZhd8MIttL0rGfCUB7fALHhF8sR9xsa2V8IyDFjT83UQfkF
G86jvX+BX2bSEc7hAWNUe00RLQJRILLB7c2crPlkt/U1ovWEJfuSbkdQiTFVzHys
d1cC31HGOYHOwaXb9Heg6metioVEBEtn9L4ZPJ0yQ+ydO/27g9AOkapTMl9AnIGi
4N2QZFXrAjUC+LLXgBgSJcRc8VCJSooThHRhCz0/rn5hlzH+J9nO+rN2Of3OS/Zo
0UE+W24560vlEn3X0tALXPRKuqfZMOAe9/MFXztUg0fcf22+8lt1te8wsQ6yVxhj
8a1qB8W14YR7eK5xuzaRPYmcu0KujtWCiqbCap9t1fdf1RyP/Q+QLYYDKadhxA45
hjEO6So5FXkgdDsb6NxODH3G6g4FxivvsRgEDfi4Hc6zGGvdkyeSfz5Q9XnMp36q
j22FZr/OHkFZknZt3u5gRFR+JSjVeZsdotGarpvtB/FE0/+9IwZzsfvVhFjowRbX
ffEJA4ETzfYWRJ22nfIpkYxBZZKftdtcZYGJpDh9lPuYgh+rcl3zIV6u6ljlietu
MlF9ovgkOomcRbWg0NWd6Qf5pgLzqA9R9qETL6U01gvzTAfPuHnB56PXoU17qyUo
VJVWWUbur5VFmjtWZVCrDVRb0pzNTIVeLRQnIlP29n2sYcEdPduZEX5EXQPfoFWM
FwhXYVpGrgciLg9RIWOf7rTR54QGsIrvEetKHXOhChwy93mxwnRF6FNzg65J0diX
/1m+GAkA40jGWNg/J6gikXq/3uDz+31LccdEQucFzCtUwkOLCT+eKBNoinZqKpYD
NAZuCvenVGTL+GCB29pPmcJCakft8bhREleIwjDUnaFGMdC9UZ1QjReS4J0B5OTx
0YdIt7irq1Obda35C7R6DR+hSp1qzsWoE/yvmB1gstW48tbXEc2+XmUQ+BOhE6VF
2N3iLAkUC4XHPvDfdFrM/AA1q49+YYfXsXWtaI1aC49ncDvKABV1pqeOblrpdg/h
Bhqd0sv+AiCJPKT/pQ0KxyVFTHqbQGePjXbCGxlHcdfHCv1jj4JWRgwbAtSFxw3L
4jUdYAuZKXCIIf8eEO7T2p58X2z5nNRTbLYHAs9zxfX5LgAi0EbTw2sW3c/Ic6op
rJl5JzQMc9GmJ9RJGUiuFZqAOwQfOyNgZmje4GpBvN2N3WniJkPgfyqdP7B/0TCh
10nOlODCCeF9OO7KcLcWvmPvQM/xyTP1ByO8B653mA7EMahI7Yp8bH+ezs7Jc3iX
L/8ijcOaGsid2irSeMLDaX3Fcl3ZIJPpTnWz2sU6UKOllZ8Nh6NSJ4KcLFOSYDRS
g+6JDoUflZLZU0pX0/Gkn90bGvGszHgFDCvDCOmGjuIQ3K2zh8uiI/79iPJIAADO
GWJihzViCus0RedxQ4adIzPT9MCd/yNP+ytqf3vy3IUYzKGVQthIja0oMu3ZKupw
i3WBLt0aOVFsdjB/vWfJvG+p0qH8p3arXidxJrNKhVUmEAdTb54I+GyH0qDyWht6
e/KRnl/WZZKktKrw9KzjOQEmohT/PBb+Zld2R0GvDj8gn3MmXOIipYsfpeLbSg/y
VJY4AS1DSmTN54lQeNORT66q9fhByHnUd9D/g8/fZdadyTN1tarc3hKOVyCbnLO1
J6D7Twlgn2cruS4Tmx4CfZS0LUNmf6Yz+/CU5qj81xs4k0Y9M9km/hnSXJwEAzob
etLHYzRVPNFiUOuhLoHqGQew48Z5atxzvNFPBBgW2GdRTbj2OQ1IK7xbJRWv2TM6
POR/XiwIrgdNLG9FwBtHnr8qdlTAYSSAILMqscxtsi+nLW5S8PqasTuFzqYdB76q
1mXRsb8u3De5YVhzYtqWlm8NU1k06yE3MmfheDQjeuPwls1rTU05EM5ALgXrx/Tq
GZZUmfpJowYbTME8H+AY9rNWDyPB4s/mpVTN52X030SlxsRKLeKvRgeSF/avl2MA
DcFlPPSXBEI1N6IYpnakI2kWNR94QT5TEPFNTy5xAJvYl1TBUfaam8J6UXlh/9hT
UIjqGxkS1+TNsKfQwfNKqcSHiZv8JTlx24SpGN8GGxOVXt+algw6N9xxEJbLr41p
3oxvAwZqWd6LYktIBMagXI/oPlPr6N5uAcuvW5h5NswAVwcXqS2ESpP8L3PqaUJR
kYjwqd688BZWbIREj5a0djVeoKJDNFtyfwQ6sJLuZHd/RJl4E7GFU7kg3gR7Y1jf
9PdwhIXtFbHOpml6ydTDOoqtx1EQqJe1nLQWUxZw/iEvUYT1OSY+zzc6CvlTyC2t
eXX766FTh3/IHFShRLlHimYVK5mThAtsX6MoKlHFpFMjaTM6djJQ6gy0trDWsjIv
67DMc+8CyWG2/VJqp7lxZku7ONfhY84KZ978mtiQ5JwEnNg5vpahJ2+t1GZc/nnC
VbKQmSJp2Qyh48kRCoTi4uj7FgoJ/rHyXbBSS9pPCQ5LcT8KVkWqHxQG7P2i63wn
vSw2uqbCZELrPYPRIaz6ZvjyHH1FvK/lw7drUAmFmZ7VTAnVnHcfepaOqzL3Sfje
iFzfDUlwaqnRdc6AVQlgUXhAsrTl8wxKtSXYCfFiPYov7NZ8np/EOoVfQSr6/nw5
WNRa0UL05PCRUJ2EBtPxYTVZ2+7AUXhaZJ7yVaE51ka0WP07v64XlQ1D+Atw9hx/
Ath3hTe8iyMZv0EDoSqfBwh0oP+4/u0bPs4em2rpLjJvgv8GEH3I9naIbBr1/tNZ
T+8uy16DpWu6eRqP642zAW0z5slAHNsvJDPXdMhSlt8Pp9vScM42H6TYGPUMuFmC
62c9/R73NwoM14XR57XUpa6qIOjt/ji50clTBm0X8hlZraWQcf7zvx3Y58qVVWUC
ZcxXwBGV47E8FsxDXgVQ/gTfYH2TFoqQQbnvYUtl9JagwnAHeLbdPkooMK+CfEaI
7t1BEa1owIBaGzp+qEsk2/nBWm5GY2RHRrTtM/1rVRHSmCBAdbmp6xBo7SGrvBky
Feel6w6CL397Quud6dsZKiHJjshYiSJCOQ0mbVpSmD1p/cPMUdUhvo3KJmUm7rfe
/NTGZcazUNCQLsMDNyrTiaTR9iEcQzhG9nwPfVAfy+tOK5HmKSnqstk2zNRREZmr
db0NwUzZkMUve8WNakz5H4Dxz/O7CRuHHjiWhxEy7/v+/86z0LijYricvuABpJhe
ftuZL58pTobK5qnQEToZ02sHGPlj4o+t5O/mYhCYjSHcBLRPtrSW92zMvsDSAN5V
EIa7oWchF5/irPOslAdG9jibA6/ftYwpbmjxZ5gfPZIkAX+ONKA3s3YHxTnoVHM8
Ma1VFfNWqpxy0Qnezm/gcx/3XBS/0ZCECdMFklC+0hJA/AjByhsOji7H3Liqc8HJ
Fnk9movEXiZym/557+weQdM5u6o+8p7e5GFOo2SUbjvffEOsRiuy4UtbDoE1OfVH
2mLxmQq9rNwN75oGKoHyUr2wzOLXjOYPlWkK1wB6KJGaM8Yhvi3UD/CX3ztE5RVc
me4vz143zAPbyCCtv6lr/ghvGP28QggrIwIvLa94zpQGUJfKNi9w8SLqCtb9XwRk
sK35WxRorgKeUFYxer42wjHnChNHgRs+TP+Kb0W0i2bJ0RnkVO8UbS6gl//lO5EP
8+BqthBXz+gKhT0Sfrn83hLHqjL0gbYVmDjEQZMP32Cent6qJ8+TdDVsBhMBBdum
SLz6RpfLMszDIzBBUU0677nzCden94rWO244D7ZoQfRHmYLCLFGyGN17Em5GTEPH
Rvd0Vm4YvS/UYczQl8/99IHijlnpM3kANSLzMvPwk40L+nNNUt3wu72xv3ARomyR
aTC+IJyCkTg3WvbwwHPbWOoIMIs1HkvfnihXd6QgvVDpGzjGgfY1lpZX+b5QmfHI
JccSanbIo80lyFHL5v3GB0LOANIdNQqtJJ7FEnXR1glTooMm3YKGchDYqKD2gfVx
AFVxTh7mL6FqjeQHOShinxkit0iCQiaONzq+nANpHe2S6Rv3YywA7m/a2s4BXSTb
tBp/b6j1Kv95nSTZuDOGLSbtihC2DC+NZUrjFqtKMf081Ig1O3TaUyVDsx7bU2zg
yY/i65hVMzQWCCbQKQhxqks0uiDXxZgg0ELXsq/3CK+aIPSEMSwPa6HWJbtf/NBT
hijVVsSCTz0GNbrh6Tn0jD7mSlZjea6Ptma9tXs3mtYmL6piyooIPqcg31QZZ1JQ
tMDu5bzf9E3E53UKuCejlOYxPDKY+tj4ZnxjzMA+wHVS6G10Fd6qXhAQGn1lH/T4
8G9qjOwejQgKPLU0OzAFAnjVv7CfRlQ6Y7FNaMmQsFnrK8aS56CVYVVhGUe/qA0Z
XQhtnwoHiosszcN1/I2O5tIAHZKzIc6RpRRhTW/HNwA/rb616emGBBVEEc6EagQW
TTnbUZlBwo0Y4NEIioa9JkdHnIhUAJ72OkwnsIFRLNyN/gyJy7OsEEpMA2ew7iL2
9vGjJqra33Fi9eNRhWBk4DoryvWJhQF0A5ItfsFfdK7lq/MlOBExSyl9m/ihJQ1U
WoQamc8hzuGa4ilOSmN0wrRmIWz81zZE2UqQNn1P/FV7Rx65N11YL+ADIN/0Hv+J
8cxuyOkf9e08aBkIRq/kVDFza1aIYoZ3qHQUkrMtN1aghIlO4yjoKt9K8zEonrmF
Q1H0pWaBUHTNXxnX24pdRAQdvsd0IAA1zwLnDR/XrReBNwipl450AD3//ogiEmzB
zh6iyXFqGAzgFzTsaxo5/poX0Vboos7dh2b8wboTkZnQfqfmsZzuBgWD+okuPH4t
b0+ZmIjmHCJqOIvcrl8RptfmNEW6mycGt9B9n9rzKzMrQxiGje9cam3h6tYqCyIq
XPTNXV99MiVIJwsug30nQU2Mg1cugAkaBF6p3UySMLgQfUKezSIz4drM/Fy/draD
hQpORC37IhUHTOTh74jhd0x8OBoRo1zPgSc3q6qyN9t6ghhzVwPhaMrfVOWJ3YoQ
THNZpkAsZoXH78CEEzdLq7gcGqH497umpphpEitN6dFdzILQoSpDMyFG3l06p9pM
fYscGNZvyzqzsamXTHZnYulcLQx6vzK3uxLR6ajK6uGYmLIgdaU5OGMbJNXfoiYV
xeo0SG6k9TRqU4df7D0QnKyaVBKa2/FuW0sZXzPeGEdgf6HVqoUG6HqGtZKy2yUa
NOPA8J0Hn2yOcPeYB5p7BHmJEQTNMlGsr6FzjE6UoEFWtyq7JI3xW6CvqUjTx7vZ
DtpGXEwQ9ptBn1yYUgEW8NMu3pQsaATd9WpKXXu10c6BCueVQC+lF389o5/wXRy8
K837npYXdhUQg//b229lU8sqG8Z96JP2R4jLH6XaeVenmRldlRGcFsPmiTV69lsq
5m8fgSlxMdRNGxt1uisptbyGawI34/1VhV7lflobhxA5g4Ja9W/rj74L2a5XFec/
Rx9zhx6cc6AuqM5IjBHMkmPk0LM0UN1FoSBfszxqNjC1XneSmCMx5TNUcUronRxv
a9cTXcOmjAJNFwB7KkWfzUWj1g44Rd3ZZT1sCyd7ayHPlIFbOO39aClxPdz4/t9r
/NkHjShJfDi+eRdPrFdNuZAJOhgXzSP+ceoM6VUsREZSUuqdfHva5042hPH98Cqx
f/CiYpm0PG/vcIGveoR9uPWIFZ6d1VOc4u2+gijcZ5UBSTSemFpONyWFZrgbpJWX
yeja3wHu/0Orc8zdFFCFOnFrOeUgRzvR0KVeus0sSbvaAsqHuwck0zAFuqtpGL9S
zc4GDlkFSzEP4kZdM9sDfBh6JOI9wWJ5zsqY4sZfAohlRCBLbXRTTd8Vl/9Ppwe2
2mmWV8hriH3t2Pwwa9urzOTEGNBSQCGCabw8S+0SAlLjgpocLa5gEOtbAk4qwRw6
QD0AJwn+lDlZQvYgyAk+KkiwAX5niCrBSptWCPFPoUq8U2K8ctD/AnzBanYuXpmt
xMzm1m0LGIn0suOVKHoGTOSpW08n46nXJKD/cYPVYi6XIcDFQZXm9X3GntafwFNM
kaURoL6/aAgWDkttizZgBWhhwgcjZJzoMEfr1TnbcoifWM5hw4RbpgzYLIQTHbiD
AlX7vopwCGdxjz5l9rh90quVX7to8D3XPVJu0Twb6lGtfrzCViRatTk2DK0zUX/t
wKOc1DBJg+zgie20OqKgUUQenhKtKBpbKojvMbydgdQg4WBr5riUepoUyg+T+6sA
DzbtRVO7K/N5rK7oJkL+rQ==
`protect END_PROTECTED
