`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EvzsVGsX8FfFTA2ePBZGfrjyj+389U8z3KdPhDcnibKBKAdYtqCwJ/Op8PF3EjBi
EZ0hcBDwOvb2nWQnbpc31Hs9PTngioA93o2Ofu3B/uH7HKQyRMtIiVpGNDyR8rdt
l31YQw4Rm7W0/+ToMPbGwnMr1zFzcpntHwUSR+mgrujxE/8BxWDYW21B5Ey8zbO6
nA9VD1CWFW3J1LSsgDqygaiiy10SVWCKi0VkEZdTlllTBE3Op8M28J0Iv/2qZRg/
UA6HnrzqD90oDxzAG84F5y8xamHVQXpl2XqbJLoH+q2C71dEtzvg74F26VGXfBh3
y5PcvKm53Pgh90MbQoC9g1ABR4JJBe5wqWsQpIIvgDh18clK+ZTmd9yOlgyeQwtI
LbanAVbjykBgk6dKmo8YxqiwvVr5EWGGymYJj0K/H0OI9JzJxvl1fi6MwIa1/TPN
`protect END_PROTECTED
