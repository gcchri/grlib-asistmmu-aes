`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3maPXdzx5KDjd1JtyO5EKBOk2emZ3wZRizRuJTlSXTWO+wkA4LZZnuPqOB+clt3f
jPyMtiBe2UrzalhgJ73p9OVsyNcnLwS0zVJUELfgmzOd+KGuBbkH7MdM+uypCdlI
TZb7tRe2QvVs9FZcXkyVKFahvqnB66cCUMJRELDMyaM2H3HihSGSV0pVPAXpT9t6
VWtMzrdAm7AnW77ElaBZdSxoBkZ2YCzztOliscrpVgxgJRgThSkvkmovuF5X3VTC
9LVHKZ+IeGYhT/3/CGejFgIK+1nd7xxwk3YojHB5ob/zEBUJlFlUfvEx9LKGZHTl
agEAlJ+t3LFOGS/5kIXQQgUuO9NlbVsuTroUsjrdNZffS8yM3kpKFwKbqib89jwM
gT0Q1eua3gOGfHs0riYY8UcMKh3J7AxlDiJWDRH+qn5UtQoJWCYbinVNUlwflBEZ
qZnxceXw3P+b7nbB+kWFoKVsd02oDqBl4jb2ngizFikAC/Rg5nFnJYu+sKyHorsa
`protect END_PROTECTED
