`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n7ssuK/Vl6jV0eKSwooofcmd+ISo7jmWYXlIW4mJIJ5nK4QDUCzV9tfIkSgL5vVz
t8kspQ7uoHLwUqPLTDoELX7bwVtWzdj6XTHNbPnXrt8JtMpWJUO30vAnzBymCPql
U5tIqAwhxrUbnriRPoXGjrznXKTHyaQY8HAtXj7CO1x4ZEBrEdZzi96OXYZzumR7
MviavT7mcrQAzw0AAQAHPD6r2iraZyV6tbWDOjGZW/MaMr2o7lAS5prQwledjusr
kqoExvXeJyzCdFVTIbTCXJPbnQTotAXRO+wYIuZQFiBAi9KL9c5+Rkd+boOsaPm6
2NQl6Mw8bYrCdklvjtFMVAcmEZlJ2uz03bytne+H3lmjx7WTssolEbjnJr001CN0
2Awqv33qL3iOKaGazI6Dd7DeH/El78mujgYzpQlbbLuS6r+fnFRGyx4ww25RVdGh
3wJcyvakMAi4cta4R9ZSSw2fvyRQdzgHszaLFXHhxH+ctyGWtoHFU76ijRVEePvs
37dgms2esEMRZ7kg2tsdWKEk2xAGQnRD+RRan9B8GUeZrWup2tsnM1twU4PO1ai7
xzhyZFIQrLS3SnSBl70zCGRD+Qt4WrB4Tmh3J1zyJX0=
`protect END_PROTECTED
