`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zQkXTfI/OTPRYTy3tld1linfSoK1UfG3aaEPRdrh/lkYpKoCgMZIlkTJSnk4VyC2
vHnDxPBMwbCyxt3WJzir1+K+bH1uy4Wb7cPbTOr14OidCoIkNYmOpPcNjwximeRT
MsCcImaDxKSw3FpSCG7a7fSS/7vjpjszdSAdyxoRki46C+/r3KOAY22sZD1YtoJb
L1+Nnxra9+VpCxw78jYgydXxAV6hjwHEFJPuwkInpNy+RN7ZkVrvZHUjuja1YV5p
CElNIlUsYhbNO7Ka6pj/P8Y+bemNCxBSkD5FCBO0ofv+0wY+9W339NI+Kb3ePgkQ
aW0XV8uk4TcFj9T7mNIt6uNartdTnuCaEqS82upgEnJCnig8YWvNKz4XZiq6VQ4q
2Wy7bSK/HrDL4FFVp/PoM/E7XxOyGRDKOnEzdC2hjz2TigOy0toO7LZbHgeR8twf
W3rRmb9vRuCcoHwP8dqVhtMym+YsR4fskO+u0z1e/WJh9znYzaw3F9nJ70CcRST3
RdpkTn84y1PMidbhttVgdUkLmXJoSYuD/qxbropfujThuhTmTwE68bPy0MvnaQOd
4dnboQDBYEZxcaQYvAzHBcY+2lr1PdA17/tIV8Ibux5xcVzmX+Matmrp0zcCRL+A
y2ERGlsF4IgL7TmGdz9oKSSyExhwEmw3v9cXwiNlD7iBJ9nJGrcL6I30an2iQqlP
yptyz4TD8Thl6Pvn8IOPaM2ZjCzvZuNxcelKyje9c8gJ3Edg54Plmkmrzz3QTR3R
3R5kmF/aob6gqhD1lJv7PGjSIPcFSxqCJS1D2lW/RsxrAN41hWP0UAXOLAxxjBun
/YMvurTmrjuUklb9FtKkitBfUT3egVorcSqJTF+aQGZ3vOZAG5QSkx3XbKoatj8+
Kw6Ye20Sw+Lb3l0UOM4ZfQ8kBf1ugZ5Rez43kV3oE9+iWs5bKf+rfDSNYAkizw3n
SCekmF+AC9Ev6Pb4FYEdc3tBCvSLcO9iuCmKwl+/UssZj1zk07TjGZHc9iqpk/4q
CFwYeBDjDHo7fvNoxqhQsDT/ohFVQbAQVlw3demGccp/Dalum8lpfP0/JBnbQVGj
l15EUoitgYZLgRfMIkkf1tYMqP2fsKFZqgeLf3NepI2wvrvRBa9ezYbIhodnuJEo
`protect END_PROTECTED
