`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nVycdLepyKlIYs6PwoMF/+ncj7YbuoSGuln5gl5SejHEHuw5gGFdcztHdUArcB7U
bhl7p1k57eVidNfs0pbbRbqW5UBPg0Ok2cipTPHYSJ2aAB76PhVKWOo8bfpeql0r
UKLmNAL4PuislunP4b7E1OYO3o6tFzeocCurdmh+dOT/Kd++/Q4hSZedhdKPTlHA
UcKWwVzjhhOYzqmx6acMrx/uULkwKWtTFnfNtE/+SGcwZNCCMha8IJLD2YQpxdfq
2ZXxGv9almhCdu8xc4Ced6VQALUdjKG7Wct0XpTelk4=
`protect END_PROTECTED
