`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
meAk2v4AErjiFEn06iUDeIfMJauHzOxnnqHYM91QXLSf47WIam2RP7CMmJBgNvWe
XWTSX6csS695bjln9ve4ro5GMlf1lnO7V1n0iMTpg53Qb28ITdIDdnpR8UegO69Q
sH1/Q6z14xK0YZXswQTKrPZf6qTzU+CfbIBi7kzHHwoD8+VlwwEuoQoTgyU9WvlR
7Di/yQUyy/Z6U/5nL8DgVqku5SzxYLPf5hgoqLhiwdD0nKEjzQRPDfg8adQrCEGd
QlzoBUDec+LDiuYEQImxpvOQj6yirdsrbaPqq0+dDX6CBKEZ3QEzl6BQxrm0zhO2
cyunAcXm8vyw8cYekfIUHQ==
`protect END_PROTECTED
