`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ee/UR4neyuIUW4YFRfMgi/UixbAd5hJMqmsvfbXf2B2uSQIAUh2pJmGR39an44Ll
dymV7JgiCQDlFjVBEMYdAOklkdaOvQ6zzt4eqH6jFs60eyHvoksh3OfO3SHt20DD
FR4io3+srDu1ttRISmVAPjftZ3y7S/Hvb7obfra9LLrbxvcE2KE8N0Y+Xe3L4C95
y/12lVpdvms1ep9bGa4D4uViVi8y4Apfi1w+ppdxZc7RwXjixoIMEnUI4ERrwa60
ThJM0dFj3N/sAEFtCm8Fn9tqpkfSNRPiv1VdjAfJ82gljZPaJTbQHZvYQEMBZ8ZA
sAka41+ryNtWXyyqBK518isd5A3f0mWlXQsKB7N8inr5hBIIxrNrKlSWR3rrix0l
BWznGz+hF71JsiUQfAhs1qCfasyCpiiHMd6UTq8rNBjVKNQVLaCZrCj5ZFo26ssa
mEn2viZbXZxX3rjM7OztPNVp5d6seE75lWL3TFU6m+F3ntUPk8AyXW8Myp0XoiJa
6Zg0BYPTTQADd9DnK8tcxWUzkBNGTmrCxqecCsciyyrAC7YqMhwhD99n9M2DM7lF
SBYfJvkQjAiMhHZL6MaMmg==
`protect END_PROTECTED
