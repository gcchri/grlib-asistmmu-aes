`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sx1E69Za5Uk7FGgKKbtV0TGSB1ftmCIF3JrTektjCxP9BlqcoKIvbSwoYP+GBwPo
rWrGBcOmYml31npjRGUy1CPByUdvimaiUU8xra4Z6pADk2Vo38/gtrOCAVRAcCDT
1uv1hOz+W9cYoM3OCRwtOQ8TehODJkc1xyNFKlUn+9BItZf9hLRV6w1hZn432jqq
Ps1DYpmTvTPDfVjXl9S3q38dWpE9VXyLd5hlR7OtyDIjqptb9KmwPAW+Yk++r3ut
1GsXHkkbvn7sFJEivelnV0UDMds+L5gknWoOKWPu6kcCredEIq2Fg+Mdo507tAdo
Pt/ZeiRUr2Jp9jhFvrncJg==
`protect END_PROTECTED
