`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l9E6WBACF4hHpKHCJLyu11xbCCHGKGjRNAQp6yGDCG/2mqf7fEdxt4CXxC672jBA
SCbZy/fh1zdi3tGaky764e4MRI62apKCHbSr3BqBqI0yaXeyXwjtaZ0V0DnTnH4t
pd45wWukjbzlLvRMHpMsEgMIkY99grbteJ1QXf8yJmOEFOGY8Jfs9M7sRPdT1Mcw
nYoye8UUUcI4otyf78TLkrdvMPQgL6XbN3pcIF8Wc4QQ17l9jsr/LvJOaLSycUch
eaCA+hipAxfkA9PlKKjR2PcaQGkN5CyvaDEJK+lojHOz7kToH87vJ/emKfyJPQXP
Z4OfzN9Rf1Vt6Nxf+kTNIvTFJ0PRu9cscuW6NneIVLiVUPMPmcQzmqJNaQphhV2C
/fmR8QcSK/wag+yX14i2LMZ3bbSIYIk6wGQ3WDuTJ6PzPxr/Y4mJ+jVWuaABVgEg
8NGNUa2Ez9eOzXF6wi9jcFJOZ1Jl3d/GyhxXfgfxjnNMVhIUFQ3uA6HWeRCNV57w
uLIBM6EMYNOfMT6XDsvKbZtGmMFUvFDJ3gheczw3/lygq4gd0TPtzi4Jlxd5xbO8
D0mW9854JBnwdLWJU8a4mjiCLd7m5mWZwM0Trwlc7YILuYRsvQmr8U0dKiW1DQai
ue0MALTOgVixp1ENJ6PtNJK7VoAoBVlJBaQ1fHdrGY6SsOnOwt4Q0sg5dl+LOgH4
5DcQsrCapacIEH/qqDNggU965spTIPH3h+MkC9JtJbqvJkzKRLKMVPkXaLOFEnxG
ZrarPodsy0Kz93HGT8RHFFrL9cQFlVfkdD1dEjVySJnp9OTfag9L3rXQ9TJR8bKR
nfcWQLgrw+gDydKh4J3zgP5pQAO7LVCwHKqTWpNE++kQydwASJsP6YcbesK6khC3
TeAq5cGOJgWVHMag1lyDLI6u4l/DWu2tdVdaVtRP9EqjeYrjEgyINuJi6V9ae8SF
nle557SVYj8uMbojBHrVyEM+Thy5r3rFmPEcXGPytTyxY9923VvRRjlIjmgLLqHk
aK1F/THVeYMjtl/ynIEt2LHwoy3HviKG+YkUnaEREqRq77cccaYhzLiM0S6ZtQ2A
jF/WxuSx7js3w2JGITko9ClLRbRjq88Cp9iKEWU5wWyuhUSXnNoKgTcqoowq42CE
0gRZfzksA8Uesb11/t7/Gc2YTmjMV23pPkjXqc/Jpaw+7w2G3E55aksvhfajQQTa
oIYuwUKZuLKzHdRx0id4+Vt95mSzfF4gQLHY5JGMAlQaVLATr3Tc1TF4+EwubEEc
E5TJQi9BGNjgnXhe2M9890PfLvh32gGGi+CR1y40SEeGGsHj8m2/mfTo2UhbTkN2
E6WNMH4kUZFCxyueV+ygdvkrzbKkVNFjRfqd6O4eEQfchP8e7BDuzzrO92XV5Lae
U+0PS5KE2SQ/PJzEaEhU9Ay/O3Wni3pLshbg5hrvm226ac9RJ4yS6qcN01vx7Qhz
NXGdGhDTj0YfuHmgdB0fmPqVtwUTZo4JMEpBqPSAa1mabSLAx5E7HS9Gm1IcP5CB
+X9x1GMFByO+waeEzyIvdNP1UXxEys7s9S6ma9ZQm+ZrAutO4VMnmioli4wRdAqI
sizOjT12rMj6qFYKaIiaQlmNa2RJBs6Ppku8Hh8+3ks0ZIlBt+zJoQ4J+YYBnrYt
y5oJy7Gv2mxDx0XeiTMEasIGDMIb0otUxV3vSzLYzrIpPaLidbnY0WbStbcC85w0
7h/ZsAIyB4OeJ4YdXMg6NyJh+e0TIMcTAWJF3AxrmkcgmXp7TrekNi6b3bH6y8YN
iEudIjy5dNnQxtg+X3dMYLq33GRyndb2E2T5Lm8m1WQsFzfAUgDLobxF2FjoYyXp
aNx7CRACJUWrO11OYwPWP5zs7+4RaMguWXrwK/Z5uf2JvghmpdG/I+ZQgaxeLRuL
Wde8zKyQZBfBDIeoYU/i9bD1kY0WHCzOrB0K9RC+cyXBUzvhA4ciRNkGlf4NwTQL
QuBjehsRLW2E1J/z+b3qydcfeZV8joW/Fv8YqJ28hOB1D1MydGXIo75/xeR84eBm
y8plrNgMZJ4WIq2YbCvl4blEE5W0jWxqxJx+bvX2fA+SihvcvZU3qF4xJWt0mbTV
w1ca5MAeNocRFj0Dmao5TiiD4Tqnw9CnTYc88GX+ylcY5OBEns771QYPtPrnHPb/
jKVT7hGqizL5LS4XFGQGyCq9W3lWrcsg1k5DpRC5eJpa3I+lKh4Tw0HmK96dL7ux
nqSbtmmsKmsMn90g7/SGubpiBBchDRJtgqkpuL6x1zkYqy2DltGYk/IroNV/FDVY
BDO+NgdxdBQh2C4Xilov0bwINQ6O/NH7wooImqX/Qq25gSBUMO4Z8GmtzyhTRq2x
laVq+Flw1deDSu4uoqr4gZZq+xm6V12/4g29DcSjhtA+1YvHNZvIQ+6P1Ycc7fjZ
fjHSdkR7c4gIfJKjjGIM003EO+UJNmNBmqH8CJrgThAbAzOBn/CSnjhzDFeN0YGB
Ljq4l3a0Ui2q/iUkMqlCfwpQKYvamAxM2hc3klEFsdctINY5tdM0XM4zmfrcmlAT
qVWAFIXKrkEI6uKbOaF7lAUtIMbpe5I7GJV/ZvSiv3Bm1LLiITF4+7FLGCe1P+9R
JkfrLOPumtinM7XVITm5htlnRWLUoHp7YS2QDCBJxHIatdDtbjFQ5Nl//mAJMkPn
oPieR/FTjNqnP845zKABjvNFb0VLDGoH8ZS2wvg6Z/xxytpodu4YtpK85urg9N3s
FQ5y/kHaSJKq9iV9Puoo+k4wQ7XfMs8CN0kRs4tWH59ZjzoT0ClLjBp2jCDA64vF
VxY49B5OdcQzu43Ggjz1i3+A+xj14s0ZEoybv/K9CJ0LsDfsGAYDxJKbJW0hmM9X
RzvIsFjH642I78mtzjnohFaZbZDLj6wHX4/Efp/u2pR+Mzhzqc0OFApzgtrf7363
eBEh3n06JMhb0GsQtWQe6iPz9RzI6M6YUewJRJ2i3CAmvQfdo0BaMgvvyClHTxYS
MNlSm0hqZkWxVl3gLYJNmtje7vxb94dq7nRM+Z1AIqLIWDVPtxOr+7g+lxfy9RJV
teB1eQTJW1zfvsN98sPz/TxSREf0192RndpSIVF/ZywcvNeUUzsavPZwIsmgSfFQ
3KAUn/prmxzysFGLMD+SNpxBJLuhxE5ZPoZD/BbXiHFSulS2P7eHEqf0miyRewxl
kfhDwTU7PbbC3deDNFhmtixWev+kxjRYoRZ81+voBnahQ+vrzYMH5bVRleFXcrPt
zPf7C8NEogNPXN2qi9arhw5euhw92CQYx0LLkT84HK+J/8jS2G00wz3QKGc6nXXQ
s6wLpMJkwyMDNfMDLfnG2lTeM7esyzOAK5ts+xD6wfV9ip1Y/Rw1CeS5dPdkhMoZ
nEU9rXjSGZV/RRNBYX233fL7SGRRPYC6+78pG0/RKACnqIGTlOeTqncTO+sVinAq
99DShhu5uK2mY/JAGtq+0rNJ5WhCOEs8n8L6CeXZyPu6RWZOAgtuz0OJj/goczyP
LWyGvbnBIjmfUmCY7BbgCVv0E8e73OmNTi4nwTq+2/izKAa1wOQTuheLagK5YuB+
9IY1S/HPXtcbzeZQQcd6jnuccE5jvWkZjTDrEw1n06jdDiJCnnqpYJiojVFXpvcu
KVPr891lq1ZXgYUNLCKN+KgJ4N+BFynOkmGUKfHiOjkYlalKRsZrPh2zxzzXrX2Y
EdKcla8iqNIAvttqlkOM/BuNpvEmT9c0sbYdp/jOV2m7R3unneB5/QienE78w42P
WGo+ZV3nW2HCkKtx5Vyj157mDRQRhF54Kc78IuFrsQWC+cypGgE9aM5KN+51u4V9
wPy+vTDfFE12sijqxzMziOVmFr0VXFDze8m8pPuLLh0MYeUfZ1vKRq2twKx4oOfs
M7J8Iiu5H1ESUZA+6uyd/WSYE413P73YcfKT8boo1zmLKdcuMdw91ZEYb8+foCTJ
eCa2AH1dSo6LjG8WDoQSlzqQpNMDx9AUsFWNLCl7aUKvRLSsnnEOhPeQkuT+yp41
GvQiCWmcJkl8Zv1wN8mKJz6q9Nzj3Bta4rb0PT2CruhYQ8dCoqa3CYlM9yPLmH3C
vCV9lsdVCK52+3DVMwSP5/Sm8kjSnhgS9hXgjUceYOCl56DT6Be5cDK0UP4W8lc0
lUj4YQHoFJK23IznVhlL6gjufTI6QsfS+uUn6dPigSxVx6f0xjTlIkmdnpFpyQyJ
lawbGGUZRP/pSYGro2ayh/0oJH1hZUYs9tsa6yYv1Tngz7NEmpadHMsZqhOkkSWs
kWtSDInreBWtGnspWaIzwaI9FQES8ZHzkfJe/vKBokw/LZgyCSdsbjdjSUzhtAmw
kRlS1FCj1gbUB7NrmJziWQjWf5MejJRcmALqhuo1UY/Tn73k5eobDXdCoWtwPpPe
C83AivpR78EvppivVH5njqWMzMMjtYJr1llVhRSKYi/Mmnrd9LMmtHw4/lziPGXw
vXj48pte47X9mlhR4/MkN/5sD+TdDrsV2l/BFMro4RTTbV+jFnSp94Z0mqMlz+Sm
NaBafgL7pf4ph7MIHd6YRw1A8PgVpR4UzgOLyFR0xL4Uw47P9ASoLH1iS+35rael
BRCXHzzwaEkF7U7go9vAvjvbdbWKNqi/Di8IpU1e73vB7m7536kjzWfVVhs9EGtz
RlJO5o4X0+MSp3hOQfGn077gUic/vH3UVUM7onUnMkGEksCN6lUQnMcoArHjw6ks
D2kyZCU2vXMQWQvoGO8zIRpyWVMwnUInNL6Nn49CU/KgwlRx+gPLF6jJgt3IF0xV
pgbuH/5R4Dt7loXjT/Mxmi7/AGDI+gma7xHZL3dHe6sWj5xinxtrNZedWf4hXa0v
ejdBv18z4rnjQkRgRSRRZ9nonlIybiBonGkadCnqnaOZbcKoq3GKRqejYTAJv+zr
RRTJYs4kLRAGf5wz5JjRFGPqwen+nS7bu9aVVTkqdGL6EnlBOpeQ1O7/H6cfj2Wt
vExSUIbndR0/qFYbAvRCAiQgse7WqAYeEp5TzRgxO/4FIASzKtUZc9hqx7DRtCO/
UttrTKZRHBh7cBe3QK7pU9AK0GduDSUuor9D1+ElQrSE0UzLeMEMe+atf/osvW7x
I+c4WSAl2GAVRq01l/ICBE2o0sSEQUv6ed5uTDclLwHRDvNtKIpTpR+aCOlYITmk
i4LmTMRlwqIokWY/BdhZenQlvv6btP71j/iq97iYWx4HSCpwCRCxWeXVpnupMjkQ
LvNQ/P52eC1NipsQeiJMw9B08873lFmJoHRwlgHw6o5bXXTmy7j4fXUPfMSe3uHH
nlL1k+oPM+CnAYx5hWlHVr0NerkVWMwN1GM7vbwjsUvao5pgbrfKkgcFh+AZaprd
pkOP/oyQNLX4nT0jSut+HU6E4c7D1MHfXnZE5DVacOoVfYvGz3khuR4Sjzn3v15d
sH8XAZAkpebVxatOJsnCH6o0htdKrrkdl/CrzkQQ+YZ3IYNj+ODvStHu2fvnNZS5
Q/aHiRASLvpfbfKoro/SxYNOPFEbELyXPd7nJxqlT2kQXHHH2avlMOyPTGocbTdZ
HgTBfBSgfCYJxYrWYN4CBfvFGEe33ePgq/R8gVN95WK8G1eJ17as93v7pXOv+ofr
2SWithDoyA4N3y+KlcLVJE5Io06kf6Vgap0JkDcZxd8evU3++V12YZJhGZo4W4XG
M6GtiR8KjgBJj7K9EOxT/rU3zWpUQL/cMJanTn/mmFbrZSX9vuq6NMraBGcTw7WI
Egiv2hZQ0YwToCuQJcg9d8Cegw8yNirXNp2axKxQr3oQJjVivSZXf41KF3P4csWt
DbyTZGLQjLcxLhMroqFeQ1hqAGVcRASrRYLEQddtdfRetrpJsKNZYPu01nw7f8OD
TXAFlnqYrdVRoG02/4NKUzJDdWV+zUVT2UMs61wPkcstXETdTRMdVu3G8Elf+gmc
DkVFxhUxuEa/kH6nGshWsn/uopZGJmCV3Wyp5NasUGfQ8jJGoAbsn/wb1hYVGqdX
k3q0CYkPE8iG8RihwRyC4QFlgnNQNnSfUVODpog0B57gv2eyW3FL2DluNdH5oW3B
K7CtNvZ1O3jaNou5O0uzq9K3uucnrcL5WRJCmRa4Aqtn6w5HqpTlFrOTFR3Rkah2
Qz2l34O0FnEy78VSMFYLHuNeEYBSE+uDvJgcaFG/tYiBwE2HQZjsYaWXERHx8SJc
ic43M520obhpTtwddVxrc1FlAhdTMC+GvCUPGhM4x/ZasPyCBsDeRKv042cP4uvn
3j2zUTM1e32OcHgxjCp8T1iWVxEvhwyJDj69Kfwa/COkm9z2BS5gSgXkLTmS/l7j
A6Gaps2nAMNQU8sgQe+1ekqnjEnIFsUbSFMEGf8z729tAkC7otrel9g/XAuBP75s
JfgqjmCk6X/ibQnqWIjLHo53EcWkNs4CYBQyZb4G0ZyF3plVKx1KBzbHxFbPnCM4
Rycv1aqhfh7D44RGm6ZZKFyj/o5s5PA4Vl2HJIJIWPU=
`protect END_PROTECTED
