`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ljs4Fa5to0sH+m8DVvJzYOqCMa4bNu3T+4F3AMmsUbILvxjPrMYsgSjCdTfzI1MI
ZN2LL8Y5KA++3IBG6C/b9/l5L/jcbW615fOJmxc3L9NA67AYkDVcVQBr6i1EImkw
vLVdUnVsf+OvnEXgAjjizhe4psEtVyJUk1QXos8iatT63NJsn9sEco6HXp+hdYkd
3X1C/2EZA3SpZPqU/fhxwaV2KJ7hfL1HLUR2E7PiUFjK7c84QjkJMMEUle/zHFg4
7GqYoU7d8CVlmVNrsAsP3RBzkGcyJoCwJejcR22morJfWeq/ikpKL93rM1xzFL8w
zhI/PdsUCinvcf3jXCO9P7RPxqZ2fWJOtUoANCBTU9/LVEw8gATHmsLP7OLNRrPN
4LzNo/QtdlgASnobHeScX7LngfzDtAylzhLtNJxlFX6vQsLP9kDRl3UqVa1j/hE0
s7LklCnntzfA3RDwYydYyPY7t6jqfyjDV6QJvd458NJZzbl8FEVpHWzqskL0Rrkx
pT5bSom8XBc3wnjOVmC30i8NnXut7Bvenu/Lk8DvknV6lpFzhcIFDl1SItVDjg4h
JaPfCXJPGXrwfoP41BNGJWVkAz5ICOPagqPGvgbuhVgyiuzH1fjM8QsfOQLCi9Kw
6zBZWPatmmkWZiAnDpow3eNKzhQP1HlrAe4rBQzoTu8Taj1+tWtUSRHQhVZ4bof4
BUOTMLBId9as03n0FhdYhcEhvKkS3v76smS/vG0dotRkl1sBypcZwy5GZLRn+Q6j
UhtocCjRcTwNyCtWGLVhl3DfABiVmBH6J+TTOl/VawPIjrbEQuLjRTO3lco1S+gz
qg0CWFW7w0eG2x6c26zGEFD2282ObImhCE3sbc8HyvcauVyJXy8lByolMAxZL08a
i7IiZtcw/rsJ1/ZIQ2BdpnCSj/qgbSSKNIrRI369fjH2JxhTLtjbvaLS0reyFE9X
7zWksONsrSRKwUNa/SjirfL9ALH6XwVsvNnGTKDDHxIkUqzckj+DwORXQClqS+FC
44at5OcEDRBpWRfnABVdTYXSCgRxLY4i9f8vj0c/b6kwsXghX/3XComFGHG1jSaL
c6Wmi39G8AovV4Na6GvHhWN0ljRoWMVbU/qFcRbavs9ljCtIE9UwU1+1LI453EnF
liAHfoxc43EWormnxtoMus/JFmbldJie3nlkpiPhPhgdtig4GI263WATydG723rj
DA/YTOINsAyBth5GK1Dj2tvk3HSSmw6OAzOqzgbJjBLruUisopQy5OtiMcP3DRrN
nP5L7+H8GXT1ukFnJNCzSY8+oBUZ3xgo+mThY7Gx0Rga+Zi7zSMtqx+NLgT0MvwO
jy/gkthMWkPdG80vc8Dy5kf3NrNMvNg8egKQ4ehiqYHaHXvD1xGwfd0LluapySTj
TLY66d3OvEtln69lMBx/k3V0Jyv7cGmfkA/51ftycsAHiW0hEIw1WAa7RZnS7Rlt
PUb2SL4rRWbeuEYCbwDBWVnGYxdqaOxOzKu3Vdr9HgP3moakGU5EfjlANk1ApWUQ
gXi2WXgGZZWRnjw8s5cWmE43OzBxniXqwjOQWP9JI2AnDnufXyLy/CCbzZVxvKiz
1YD+/Ktps1Hw3zOQrsJ9TWXjWLFM4wQRBdGResTeWTZXkSuuAvVLgAlLawBZ1pga
szihP4rpnaFxfH1cdE1/Jcw4KokebcP6ZbOUY1554Xn7LGbS89IwnfUvenwZmoC3
6LL+xxT8h+YRdQukdF2JrDyAy0LPwBIl3QsY/Evzv9zK2vIIDoVkBq/FT2J2OrkL
df7khkF/Z34v50ecCzh5G8D5yjj5/1v1HDNVwWGrEfDo5kKzcbC83cQGETm7cp8i
ChbvP4FsAr9hcodln8C7lSfrd6gLfeBSCUrBbw21WSY0ozKsAdPcfHlQ8xCkYEUD
pQFn54xt96sr2rjlPg9/RkOmVPr5iEM1X7e24zFMYin+VVQZSvG+Dxn+ZtaQOMyC
TU8utK0I03POa/QK/oe/aN1+hyOOes1dwKDJQvdhj8Aj3cMs4SqGiaoJGmfzRapX
8aZnXsl34IJJxe+k3eScTjG5cXRqsSMihrqN9RVOU9aGZZjcOLxtsRUj8o/hhNFo
oW1OmjXSPVKojGjC8G/O3WuVOByf1MI2nnZ1UClYWS43Iv2JxY87d2TtAzL6dCKK
d7BqnOlltct98RV1Cgfrj3Y8eSvgfvtWM5RAiKzQUqsAXmss2CMZ6DhRNH1jSC+n
knzr3YAp6STP9bsXUmyRORYsZngmbK9HtUvt3EY2soDI4qppU8pHdQZIeRsWEsdR
rRawP4wXY2v6+kuE56BW3JzCmFRfxTuIu5x6hH61dioLH8dXQDj3G7tdksEVm0wm
N8MsuWPW9PsOLPe+XFZAjy4rrafcAlrIFvwSE2obsSILYA5yJXYerDsPMTp7gW7E
4nHDRlWtmUabwCeUhNntD2Eh2gz6kAPZu/ePH3XoBv3RPEtp4jv2/K6nCTTuxQS0
K1Tg+FAZ7WCohmBgM9oFk7FhIN0moHSW/hSyQIgZDK6rQFopvHlqQoaN6eBgnbSk
G1awXTsiYc1dCSNdgCQXnIAjDFsId0+DRKX6SWNLxnAgp63TBgcDnkx/hYwrUBh5
8TNabIeW9jFFRFMKHrh89DAgpykOaiT4v6Y66YLu/a9A0akxbJhEvoPXnt04uw6k
LkNoyfrGs4niDJEX3Y7dGFBr1fm27q05K5yXEjmKfyPr42Yx/0z/qsZ1QTFvrmqu
v7VacPcCnDYS75rr9IYzAQoaovfdFIhliNhzu3KRhLRwJIRCuVITs15yDUcXHs91
WoZh0pkiCCF/j3nxOeN1ntDt4kuE4fJmciginMNQ8Nt2BI+s4cqP4ZfTJFT/dDS1
vFBpJ+M3wKJkWIVWhkpbSXwKXDsJPPD6tf3vcQ7fOvzV7DcV6OhBaQCG8GxOIaaD
n2M3wfEgXRK2M2BvFYkRXo9/g4Kl25r2mam5bWcO3ABHmHzRgTzBb4I9MhYUouio
o1B2sjgMsdFT5WML1mdTZBiDBoGpl4BI8jkaCL4DAi8xi9eipg61N6QA3kD5Ov4f
0mhlLLzq8V/ehJQUtAUSd72sZwkZHhN+6yltzHjO23L8VkyoktJ+uqvnMnZ3RNYv
AnyJwtq6bNhr/QF80KuFXd9phuBHTMZ1ROMJjLvbT7ljG8Gpr2FUWmKx4rNKkypW
/iDb6H3FoQxFGhF5/9Gkw6JJsg+NjXTHYr0HK3sfqfSb90vFm5nDDXj4lqcAHN4U
v/pJCNM4e2dAtJid/WAsbHaADC0FaEBIbUOqgD5HtBB5UlaFZXs/7TtZa6P4ewYU
41p+wgA8TJFKvP1PUGEtcg8Ue4th4aSItlC19GQIpOfQfMngpIrQZO+rIk/ym0Bs
3Q4v6cUSbFiIlidG5e+Kw1qq+4OsWPWRnuKWc/hC91ZJlorwn2tm59Ip0NHuSc7b
ndxrnShH3kORGA389jCsb6iyzZfCyaLOY9yKKdVGkI3L83TWcDSFqj3aHTF+FGsq
zNbo3xBJOOW2rYEx2tJJCSLMNjGGgt7ikrI+Yzd31ELjFaL/HY9Qav0wr723JOpV
f4WSxySPN7VM4/Bm3sBSn9NR/aLDIWkwFmLHMRvQSYCTUDXfBwM/2vecNHsfCbx6
aRV5/TCjd+o74fDj+KgDA4b5USNQob/qFLFoNnX09lLsS1iOih+juBZWGPU2EmnN
qeEqm6Se44GQVDC92c3jB/vA7MJRrt6Ka8Z8CEV4htEnQWP8H9Y3pF++7nmCYrVY
6Z50sY9pHzJ6NZsSw29NUZFnNPeBnl6zoiP4QAmCNcpXv3HO0FnWDuI1fSRmK328
hywmkIGeuR9AcxWRa3xCYcpNOsBd8c1dnukZ37ocf0VAkHcmB1omImRYbs0T9obB
gKwNS9Vl1+6v+ik0tdmq7ce9aM0hiuyXntpSTdXaRmG5lFocj0VWGB+DTIyo+QVX
7/GyXVx/KlJu+Eeba5lBRiKo+gyfY+LU1P1Vw0L8CfhS2jOLhXPyZsq6tRI0X4AP
OmslDPIvHfiIHPu//lg4hOhNqYbPugoBkqP5ivimey8iC8IiBDA/Z7fKS/GoU/UI
RJpgt0Ez6fyU/ksn78ul85cwtOm+8nh+95Wv8MPqL6pFMzNT+t6Os2Ij57YYK4oH
YHiB04vbx//zZ53tM88BT4yFNjP1VklyA4X8YqSukLPirjeUgWexiUMztpRWxZNO
A947PXV4STCv7AgszfXMAsmu18gaAqLj69TLjy6sUZKo2d0n4B5MGAWW7/3u6V5W
9H977vKuBMLwQWcacVS/gQpDlVJGvsOn1X2LUPYI0lFnHkjHMPSu1GLoOeEkApku
XNcjb7tCJjV08nFBmW3UtNHbq6FhAjUXu5mpJMNrX6bJzfeAJIV/J/RqW2ZyebJq
ZAjq8Q8YYmmTDclRHB7fwSxf/q6Y+RtAb4ErF7TXRZlgc7I9EtkM2vPcjKUkiRlo
CspfudaWwG+k19Ddpsh7U86x6o+CWXscKS2W97BlO2nIR+mN6tXPt/31z+VishDS
rnas5vpnJ0mCiSEayzPWuXFuX9UdvaIBFCQmhAL9beT4z0/912eLmPrjuT2dyf7V
qTNEN4XM2YtCXP9d40fa5Yh42oO/rxnnwh8u1tJ3Gvnlkeip7eJwrD0ha499z994
+g9YHu3MZ2bFpRv1gtJvrAIvtoe5ava+HdICKiZsg0o7zjEGe6ZZYaPgiRTj9xWf
SqNAbXh3yydgrgGmIvH+NPGVWdPZ3VKHheeuK1XpvBjA8M0ih9ZMndCL1dKD9HeB
MFf/J9E9Hnz4CDjn49c6AkewGYPVZh2N8c6lVVSzVryZ6NmGWEpMPzuUjDHo3jDv
xsta2WPP4hRQ055UWHKfwk2cC6zVLz8Gbtep3Y/W1uV+jsV7rNxFWBLbI0/uS58f
ghs444fHprXZ1tkZ1sUySHoJ6EuifrPit9h5v9mT8H2cCTaKKGYsSW8amdIZQLF+
0afDuoH5i+XmFE3XmsQcR/uaCbHfi4FVN2vrm1pbIdaWUjgvmMhhq1tazOkQQhSV
fYwR9g80DGBYYc+hx4nhSr/OSCB8lERaLu3kmaxBD/fElIRCnH1tPNY3x/qzk5KM
72yLWapOhRGDWeZR1p/ti+9gEbvwtvyWrLYM1dF8Hxb+6eeT+rRnDaFrxwisFY6c
anpbLhOhLmA5lSIDIqxiH2kEnWd0nZBGBSqKzjh6LxsthfCoNLrJnqffeiuF9ng1
oRr3O1ZIIzBMypoZ4JFC9l7Re57ST6JRjm1zMhAubWQ6apRi4x/GhsSdch7K/X6/
7+V+3mILAD5Ti7OFWA5NJ/0ll9oRF/Ezi6TuGbKlLUKvYnHxIJzeULoGmZeGwPbO
izWfci1o+5adDCgjaK0EQl3bsRrwxyvB0jSe8zV2RfD3v47TaXTBP6RsxJTdqGCC
OKgwWO3DylQDDhNthtXLh73QHNbo0ciyxPVCmJPxKHu8jAZwSb/4r7NizlUdLGro
nsUvfquo++NmU3/zV+dke8ZvKKVSn2Pegi4jBI5n4HjLJqoyWQrz/fS+e2Y0A7W+
EpH2LF5ZF8SFvfhD1rEGv1aMkOHdGBXG38MHu4RisFnDda6cx6JQAxAdVHQfTEyk
DhmU41qjhQytiH1dstkkbDPSgV/l5CUE6ff2LiGF8AP/Pgqqkq+8o6dMr7tDDj5k
CP2l2CZ4bSsU/jUOYks1AAfICHJHkkE8t0Sz8k7fTeZpf6FWNtanBJSs+5MxbrTR
D1ZF6o9qIjDb74spXVR+aTD0DeYa3V6KKA72bQKcnrU12gr5oR0ggsVJWNYRclh7
G+wL4XCSpoj0Hs0gUc7uDeWGnFMokjIIrL2AKscSX3oMbkcVFHonkq1pV32A9o+x
V1vSfdAmqhAzM+Mkz7Y7uphQaRLIgrQvh2bnkvXg9nXolqnt3z46U4ytIl14JuNY
+tlmhV/MbXRUePi/b63pFwAyqjok4mNOEGM9qDAwDOcb4/MtAiyDZQO4VaTIAV8K
vzgL1R5mma4hQIUwRcHuKv/AS+skHmOcR2mt3UHOeIoSjX6BWAe5ik48Y27rO0Vm
35AXNHLrm4QVON/ccswksG0a1++GNQJjvhzRKhemiaQRtqj96lH2lNdoaJFXQpZH
f7ic2wBnyTvcI/uO6QHPAiTYWhe++KJ3c1KzQVz9vb5m640nr/tCw0akD3b5xGiN
w/D+wnN2H0gLNAHXJqbOzdXvKExBrAnzV0GmZ8NEyoscMPnk3kaMwV6T9GUHkE5i
YLdjkMHZmbcyznBqpng676qmPOL2A4qCsMssPJTNdIZ9iDdY5DDWn/uqtjN7s/Se
fDeFR9lW87tfGnTxxdfTqQwXCTmUcqexBYFiboW/nDi6GGdIHwki/ic5jFz85Eye
pltRJRzRxjZno34/BY9483b3opdtCR0Zb/8XTx+5Q9h1Zba7/b+pFFVvHbo7G3yW
lkLH/lADHe9gbfvRCmHSyplttDH0MFVAxodaHLF+S7R5OQj9BndnIagKsYNAX8Wi
EzBos1Cm+jQ+lvI7lK0D7PZB4U/0BHOhEM5Y3aMNmCx4R89QWGu6ZcsSdIv44nCr
0yL9XIjjmCydBLbgbzaJHHvPsCU2V9JJ52JDjgJT9dJURYJdwkzbL0hGbweJO2ys
7/RFv5GMAmh2zMd23NvFGquZktfp1dCDnaWLrLwY2ICNdfKgq+71GWgrx4XcIAxZ
m/caewjO9XS5d6g4ASa7+cXPFL0CYY64xmXs8ktlftzilE9Ew/CRAaDD+XeQfLTF
Y9q0d3s97QHhWwbIyeoAd3OccRVkXan8Wj561JiKVqi7ddXHhK2N1vp9jnMCjtKk
+19uopF8BHunSRt1NS0IhoHkUC0X9c4eBLJwf4f5yZDT4X7dkkqA1rNpJQFRkv6G
G6R+PXx/rVmvFh4n72rhgyShl4O9DGPdQmNPzXse766jpbpGXzxYIBSs0lwnfa4I
TfJu26QGPImDcqZC+djcTp0IbtOSN2KtjRJSbf7FrPTlvAEsoNn9XrNQL1bTqf8l
eK6vnjEdY//W5wvJCoKLBkTv/sLV/huwWmxGHfFXgO7q/fpmoxJK5a3ZPn8HgnYs
cW47UmmGtDS6A74YVeI4LAWRLDL1/Q+EBLqObe6I5+xCqW6yW9z6QfiHgNr4pP4M
Q2EUoXOb7kq/Fh/ZWNc12BTjpkHqvDoLzDLZMAnMKtauFcuKQ3qvyVR5KTPI5oow
j376tDBGq/O8XF/inP5flJNCgQeQGoSQieazqhRAKHjhSX4fLJywz9fj73hSdJWt
k6T56jIk0LNsh+Jdf3+PojmoIGXD3+HPk46WHO9bQ6T2+51D3ONht5XEk+BZW1AZ
EO+C/WtT7dNrSMesFwvieXU9WxorlyBW8wSo510oWXXStEwkNd5XAfeECwTbRJ/B
LG5mppgDaL0ASiD/l4eJbdbK0Ws+8PwfgSWxkhEukvi/YJQk6y6lnFDhJjCgsa6m
+uUBK+O1/7zDfLTGWubR8FzIRjxuMIAyCDsaxL59y1NYS79YbYxIzDMINuXEZ5yW
9HunuufAK20DfhJcApbo6w0Im6WHQf32TpmE+JzQL5er5ebs/7TY7+UQJIPI1PLN
TGOYKo/mqnsiNd1XWj7s2OFaE0wkkq/Wac+s5h6AU2euRDPXnjkIUnLieXQ5XWOY
V1toylN+JRLCvERXgIMQAmHqKb5LiUhzjCGM6cfd65sJP2Y9qrgwULCwLFrmSvzR
yhBqNbrTfqPKx5idlPq5OhjW+hDDpa5UsmGsTBfEEHPVowK/vOsHxwZvrv0zC+da
izMkEHzCUoPL3NUDstey3j3KezdoG9rXbQYIrx3hxrNT7H5USt/2hJrqHuxTXgJH
cCmIlIYupElUnABa/Zcou28hcUW5tRr96xh8+LSBBovNGxM+9TeTpXsUGJzWCOA2
dS61vk0KmvruACx23oBLhIsYP9xQcy2no317vv4Nf1jaDc7AAtfB/ldNWCLdD1e8
3SwvaHYbOka3ANQZgKEeiJAXhcK+ZHkX/yT82n2aKJzEWhnd5lolGGngNEwWP2E7
bPMSGKKz90AYp4QK5b76fISdkLCNzs6Aw1gUAZ6UJsPPyD20FWiTkI/xQVbv8IfP
rf9rrugXtGYJx2g6evXz1/fVdGGOQNETPXBNcr07EbeEtP+SJ6rSXVsRuE7iI/Wa
vlbZ1+01TcV+5Tx3YT1CJniAnv2W/PAjWYlfM45sdUj1ozdzcRrTz8DZDyYGWuHx
+UeekwEQbIvCpzdas/c/RB6NEOZzF9Pq406KKjMQmL/y8fyQnDobbS4qrPp23n/H
FFYa0DBFpBDH7TY28JBS+vvdhyWxA6qoD6Vg1vjwpKJEhISdAunbNRhuHgArJQN2
Aj/0e0MblsZa7O+4Szqj8OQWjL4WfbR8PkTn3OZ8CCyAj9x9hp0FyUrQkkKbO93k
xob4pHdRN9snm2WMhhKpIqxT3hed7vb4Ki0c/fd7hBJ4a3Z796i/RBfT3wvL6k+4
thBgLbX8Ph0p9olWTaVG9dcAdoXEcFLezU/A1s9JQbq5wKC8wBVLp7PnliHyWfhm
TvFfiRCY8UX7RgOeLOmxEBS+qldP1k+2BZHEzAvJIuG/cYfeu7jhEUVmTi70flMQ
4jZUlAMJ5YIjVJCVAGgL06xTpqp90OVxmz238cbjP7BF5pTqJgx2IKjHsEeIBObr
DQ5Ujlf0/yAiSopM8F5kExanRZ8YsDXN3EbRVJheoEGW6T83KS681VfcnBdQFwfV
VnkDYlKTMkxBcu9+k1Z1Fv47YyUP8svDle4/0QH8zx7KJgk8sqsLG4URSCxQ0aCp
oKyVytVt8ZONRORiIVL90Wqvxf6Oqn5zliQerOrNEZjSxpTHbcfr9eR0BMoH/WAS
jzpAjNPqjfffeK+IGW2BPVE+LTs3XNqaFP+k5RcfqV8ydiLEsEmc4CeojwzZkix6
9eRk1hihhT754G8EnX/cMIWc7fSxQ6q6Q6mjtsUM8MSFxq50kcLpEItKaYK7VJ+2
GOLgNDzamR8UerQchp92jUESZWWWKoBa7hlTb0BpVUIRax1awU7gJS82xY/Q41A9
2PAIwCKzy1FFkAayujqqCUlD+sA+60Ar2d6C+pun2IRdVb6EmKpRMSA8j+HBcodv
YaDiL5O5Y79jfBX+KXiqr0uFLIWlCd3AsQJN4lXjQwqVOBxRRYeLzh9u2338otXj
uGZkFGp+2hItwVHVbUx0JtJNhHrZFHfp/jLlZgE+LbcwMfG5jPa8dpf9xJOhv/U1
jErAG7txlhrJaNYS6O1EauRVvPGVH5jykMMWeYCWpOX4kdgkOJfE/ODOYb7cVqzR
DS5kPor34zwVQ+WaxWVq5urFN6VXOgSE4xNh7KYBiAO1YpCzLsF8VLHi5qGLNaw4
MQx31jun//I0O5w9oyQEGu3iUOYQrjxvwME/1VklsCAEmjXIYIUzfJXWyJtSNJ0Z
XsLSgQJBP0fl/LHNj0DpapeAUrTbjLMzzI4n9ixybckzV528zWtaEXug1aBPJrDA
8FLxL3FXH5fj1Zudy+uTPYd+el3TRdT8K5jIIJVSaWu4jQgoZ4PfbQopXUypZWWQ
gr1BmT7jGABDbeLKf+va94Tre52KPz0X46hsGtx+U9dC65ItmOjzcRHb/Z3J3deB
uo1AaHw2zzqALdJbJNrAIAmrftj0FIc+8z7KEbJ98KTPIf/J4mww1M3MiXHfi0Y0
N1JNS5/9fKGhDnAhomUqam7Uk9Gk7mkatch/OUzkRfl1OxOcmRgQTtxFumfYmKtH
2ZN1RGsshNipxo6pC57rs9KE4jv6lGVVb8gWm1p22xujd5KVd2OSLXt1XQYZ1a2h
H9oYYu2t0A99uzzPHjv2/s9b48PogAOUJX313S6GiJIxg+WlTl/h5EHHCTi0SGgH
a5SKbS4FTpdxBV7BUNn/3kWu9QNT94FaXMqx0THKBmHAasDA2pLQh9AyPakCmmw/
d8Yxw0uLA42EM78iKNYJAW4zQ13NAtCfobL1q3TKOAJ6/o2SpZYXgbTCaP7wU6IW
MU5uIwXRhDay337nypD48A3K7A97XNr3pPiTQZCUFIZcy7SQ0/gnTTm3/NaU8/3J
bFRmqFoa28RlLEqTVf8Es+H1Gb6rfi+mc+o7uDmGCpzT3Nq5yv/tfceziOXhbcju
X17jfYUWvlhkV0oaYTcQVvNmj5fofWAzrxn/Ee1DAWH7AByVyZaX21jxqzhhXxiv
KU8D/5epDVl56cs+UDv50mBC7UbSdmbKzFuTO2ySqkMoQSqmDoV0Okw1fgxZcIQJ
X+xOq2xBgxpmEp2qGbBEvdYcuBA7NWrmY/Xu7FocPnzQQxlgUV9T63WDwSHqkqr/
hAJSsbJXkOo2wxTXdC+GzeoJwDaSLrClSEzZqGfwDjMRnR6lqyQv0zP8dTtz34m6
wwLIPcfE5FdJ3H/ZkZYEPvwGbRzRu6PJ8e7eOg5QE5sPJcgC+YU0tb33SvGBXT1p
plf+e3mdWVmJkfurVkrIe+T4IqVbUaBYqxXViaB0gbrGzKbDkEYK+7J5IVZtyEZs
YKGfQPwVOdbn9oKPD8c8VePkt+mnFSrSNSwPerRnge1YRI8CCDsrByuwfdT6+I4K
YpMMXyhVfZ0s3Rx2Ab8h/rMFKwpD7PXBSX7sH8ey9Zk4VHRgXPWWVHNMMODx5zch
225m1GJuV2JCt3MVwLKPqnqahnVZu7oRq/dvxuuXcjfNjJ52lm6sbi7HKvIBq6ae
4oUhSHhkn2FHVQ/ScewtiHr4dp7foxQbGXa4hHliSwPdHcDkpB9W7XtzmG+oGw2a
HAd9Mu4A7/Gli9iHNkpa5bsyaKP8hhJKl5iFJBGdBF3EKiZSEK72aICuNtPknPJS
5SgdDs5ebXUAY083vSu0dXv9SejHZEg9oN7+wZiYQOz2Qu+ATxny/UltHKSuWlml
BTnrl9vrf103dfZfwcVI+Xq7+oChuA3OWmiNdPAa/iJA/EV6Oc9Zh5MNe6Uty76B
cHL0J3fkoNfXdUXcd+s6H/I8iiZ+atIHEwikc6tO9shsXSnjmHZZ6lfw3DFj5KFE
LWrVjjUS9T4V31NiHnzyAg2QzA/hEdCdeBSEbzDjF8LnMjqG/AYAcne8ZRDNfK0P
fJB2NNPBfGm41kacRDi91G29dyD2h1RZHZMnRJtasSSpiW9v+G8jei8plhfX8Tsg
fSiuRyuLIBjh1ECQ801MEOYG8J122f/KR/BmM13F+1awDrfN9TWg8x9JYJAc+8nz
DBadlQQsw7R4Tllejr0UNTZ9V/3BbfwgodDL2XLfRxyCo7i2zhZBE1z2xR0cq8qw
m8XYLoaL9vZg3lU/a1V+/rFyml4mi5GAss+OqCt01Nkv2Y2RdEYoZOB3876B49oY
X3cAGEkNlWsX+HC4AGACoX1c3cV31WDSvtnaqaW0kptpz8fzz+AOqn2vBRhBOIqj
llJTIkKTHY70dl9CBranIqeO2fGpdLQb4OSG+X1x/a9dXSfzhCE+cCxORIlbfNmL
VPOY1WUA6WX2L6UEyARyPsDbIfToEzLEMHCwSGNhtheQYXzTUn2wDxduM1FxjrU3
7l3Mnbf7LrpzYPIyda9i86hdCiW4rRFevtpzNhFy3vCPksO1Cl6EkCyd+Wf7pNB6
g6rdqUQB/3GQFecgYnQUTqgck5RGiOjokiY4dkFPAe4qJjHbgTEp8p+ohHQ03LMj
HSMPtJZPgNkuU69KuaLZ8lBXI+Ys3jEP6J1Q+Gv3YI7gkAHCE+MwomVzM+eSgOrI
UP/h/ABc5Miv+OUn6+3TNePhOqkEtYGIN9eVnh7t4ewpSvQ/nQBg2dgtZOmv0H19
+VOSiwvr5x6jJIBCS14P3ZzrUwHa9Mf/zcpv5POHQh5D9co6+3isKF4y8IqVN9M6
vZPLHRCufUoilix6vBOJVTNlgYsspjcWdywaWONifrh3yBGwxiX+8717gfjbVQhF
YdlH52xwilDaLKNeJkncslKXYWA+LlvYPiqMxOA6jZ6hcrPB2RHrSeMczcUpULyJ
rcwlvKxH2CI7x/aJGrLglZRoYRYe4CWQvhGBEG3akMr6fBjPmU3ougOurpNzpeXC
9rq+c9hxwuJXzMJ6MFAyS1xdGTmBApPbSXi/mVb0NimyUNsMfiYQpszATgjHwyqI
ll12u9VuIts4ncRDBlljIW0KD5PwFJtCJO0nHSddsW0jC1sWeXgzdVL6SIyXbz/t
kvznUrqFzFRxWU4sEU9ef0kL0xBW9vlHoanhu3SJq9A3Tm17iNt8aEZI/ZAh1DEj
HWtS4Kub2mgiUuqQCrGPM0/l0Rc1w4WfTjwMP4yBioNi4Q30dE26z7F6tjQByfbH
d4WjDTYSn8LErmq0apFDsAhM16NP4qqqAS6M/i11pdCrZQNO0qdC3Fpn12q3quG4
C9cvJ8Jlca0oRxxsR4FYWu/dX68iS0hnqTwThdka6l1J8UnhIgUMMVucZuGl1CUN
BNk+4wr+03GXWDWql8bQEeOcWmpQA7Lpq3pMSr5NyEs5m4Qx75yFnowo9RnAptkP
jRRhAN37VSTIAeHMEWp20cgf2m8+KXuO6Q9Ar/ABsDi8vKOUjc9j+bkGHlfSK5H5
zsgG6FZTAicMNyvAQCHo1XNEzf/UOa0NWjmkXzIii2Bxwnli+MULd+AkF0gZfGe7
574EmNVrNq3OB6WmRj4XlaNvDnFaOLgjzHIkVQCq1l0O9tMExAR7lLqEe2A6uvzQ
nLjlYchfZV8esfTFDqNvO/7aTJ8zje3UyQqumqAke3vSKZeYV4a3KG8LyyCgWBay
2mi+1SLUXc7QXe/kmSZ8QydwQRhEmzFihD2CEqB3CUeqUedXYBCYc1NJtK+U1Fk6
sXCP8uX6WEi5ORTOBdR7amZcErFGXdAd6wBUnQ7WgVcbGLhL4t6e06pdUs7kcaTm
vtQQr0YkoByI7KCO8vcbqeSuJ09/L40/omDh8wR8T6aOAP8gf7Mj9Z8E4U/PDIg5
jblEVaW8FejQ05TObAk16ak3dXcowNpwfbY2VuwTXGKNPq5M/dLqgjOYB2UuzIN7
6/qWhzcyxKvwf9WFZ6TKbA/kfxKiIEAo/WaTFjajDzXlxSPV/i2IVqSw5OWyh43a
G0RIbY9ScD3VRC/Gkb/m3a4LTny8W8YdXi373wI3kOMQ5KKNh4V0kiXj4T8ivXtt
5WWfsBotDo8rfuJIKDNx9lxE1u6rRHP1zbhlU+I/pgepDdhb/3r9/SDtKzrUir+9
RMi/Ce50ciF6SyyTsPu4G/1BgInjFhyRpSjIrIGp330WqTlzx9veEZc6BOPgRrEP
uEQHyWKoN5DVe63xrba9vGhxDCRB2voT8eZ/lII9+oNtxkAYywsRJ5W/lplqH6Dj
X5GranKdwUv6SdFwoVMO+AFR+3ggO787Sf1MUGyEc2lDGaidC54K55bMPmYEBwgD
ZlFrJWvLzxRSYCmOuVXZc6jyExOwx140KzwiLHsUTWkld6d3LZN3VKa7Qi0w2o93
Ve1H2UVbNu3G8Z1pKGru65qUyN7AK3RcLiX5qRry0ZD5dM58ibyFj6a2pZrJNIL+
FauZeE5PutgxhJdcS0KqVw54vp7aWUbzE1nWqk+9llEvO0xy5IgpH7+c00yUZt0b
EVDWamu5wxLiLQrACSuucmR/1dRyuEFuqLS/tijyKxxO5MYKaPYoaTlOpofT8VlS
2fbK5cBogHQQsAzxiDWopAvZMeFU87wL8B/oBPKGWfxauGE5mcL6/0owqYh9n+Jq
kGQ39RFW+iDZ4kNd0LadHujITZvwCUYxjUhWaQSwnIDHvWJ921JRFlWhS+v0N/8V
2ChToX5gM/HAyhzQJD79TekFZBsy1RENrFDiKLqAOy7AmPq8kUch+PnrsBGPJZKe
YFWKXlQq79KSWrowRaHbTqhMZ0VG8opi3RxeASZ4wAldOnGt7sDiYW6ppAxCZ9/r
wxcZ4hrlflr7QkDleuPiF7tZCeBMLJsFS2iw3Ai4c1WHfbAYPpzyPpYtSYZkpHdT
CPyBiW0Q8zBUJz0AeYdvXrYtSDhnW4A7J23xD0jP3p4xxbAcIdJKCrihDmtJ4HeJ
Bgs3ITRk/7kBkVfymV+gpAguTMwi6gbfrl7E3gGBAAOx9N/KG/BFLmIZNRK3hbSz
EZEBdgHceDB46BQfHAejxPvXadlg+x4pzlKFtiIaDL5hFjHihOr8SMPAhCIGtyG8
mDEJySUpqsABT5DXxhAKxLVaSaL+ZFtPoEaobrAoF4kTNRcPAYZeCYP2Q7nTNaHd
0PRCh6fprDOVjk6rgRkhNeMlKYzDa44VOWB462ul1bQrW6WDXvMn1NFEMlkNxPoT
N7/XUggm3OLXJWipl0bnIGNaYeycRE08er52smOikgRUZBIovvvpQixuFk5IQjhY
pdrBgd0S/NhMCTOhQ87owiIrXoO/ElMPRsTay2Q6+f28jRTlRVbFs2EQBf5qnNiN
kF8eHAMsOBLd8PZ64Epvspw+aOYZTZMTFQY6fVA8zGvl+cLklYTLPmgvP66/JcbE
l4U28vEuvKh3ILyia14TcZnRDSThpk+8wWjpURdu4lisM9XnzGUKYDusniT+5csT
iPHCBOWabV2m+VSZRbGua5ojvha7stlAe4CCOSZ8lOfsG6JY8OVrACkKa7bB3Mib
PdPnx2THI1hjPR3+8lyHMpCAcnehw5B+UUZOh0BUUQu5E8dllqMye4kGrLMxHdAz
Rf8K3qChuN8jHgIRJMd9AhpGpdvj0nK7+9futQ6Yce3jxrPlG4NOcEPuCd+Z6FKT
ccWSV2OfzPYnDpo7JgFRorRMkmAjKHm9/vd6RpkSTv8148ZsJP2hkIyWLxPfgDnk
sDr1LUU4wQEwRATV1R73y5yYRFemEd7WSNlgkaStKl0nHetxokRg7HcI8b3DKjRr
k7MZqZ3x9mZVXc9Ape2cYzda1WGv9wWpi5pKFiOF9f9LYP3NFLCWt+vD4Vna0PSq
9RAoWabk/wpJ6LCzLy06/Fy2CnG+0pkOo8EI5GiqTx+f1uOTpAOcAItxhvFUC/AM
IemrUBwnDG5XwYQk35ac10Xb74RvrlJH3dG8PpI/7ETNzHY/we3LV8VNWi7nHN9n
duy+0SPi0o2Tz7l22xD+lACRslkCVyFJIXpWapZPknb2uwCPsXbjqTsa26Fc3ejF
9fzERkTbQNTYaOOXxdoZ4VxcxatpnDLEh/UMKa4c8mnhD3yzXmP9as8G5XBp5dCe
E633YD5ZJXCWTk1C9VSNoh8RKLbC+A19dP/2wKwnuch8gvisC9YbPijZUKQpQv8c
gA5KTScfppm1z794KRgZZdM6lKRUy+46jqYSruMRPmNoU6p6cyXZUPp+qDzoS8aH
Q27cA0JabBBCtfwWog9M/Y7zV55TlcLUnhJO94zJn2YlphS9y0rYyY1YjG8mvzrb
hlJDvowhID2YVg7AxoUzJo2LSVF3FQsI9aOKhO/Nr2GhWGzY1ehJeZ6IbSJgqjic
83z0eZIpnfKO2ORjTUvCVQJnP9lRMpKIleaZzIRI1vKm9lc/eJaV9X4AZJvfjolg
K8NLVNK36ub/JnuyKFlluCXWNlLGKZFcqsnBIF4aBoqbfHIkF1yUHwiKpnD6Ugff
wsKSpM0Ph8TbKU9JAJ3wQFuAW1H82dQOTOa9umFR02nGasgrrV2yQfiz735vcOAD
0CAA3LllTrjQzovG6WKqcnEnTfPFJHsoL7S1sPQbS7cdPpn5YlwmgvRe9rHlAOMt
niz4QnESBgxkWvUu/BlECj2UgiNJZscVv5TkV/5kxgZN8b78zjZ9nwOJAxn1i8PH
XkDgqimyOczhPpI7XExnQ7+9z6w5ECtaaJeBGzeIhGBcvUcYn8B3hghAxnZ4kGbO
rML0jpZJ5+PI4/L71RHUcwFYi0+JH1sT+D5RjwGfS/PW1FKE9+gQ+wIAMzVGQNXe
YH1rBTLa0WjTZueg8wQ6ZhKDBM7zFjXXkrU46KPRyvf38Rqmp5Zo6aOc/21qgtWG
LX+cFXed6cA8y26l5wYJHY5vORF5vUVQawFt2u0jlC8wE7zJ+y46E0dEshu9s+yN
M3NKe0p9cyp3PrJF07jBAgPEBEyb2N6K+hwGH0RB1eEM9dNjbrcKfk0u8+I1eKe1
JfTwNusM8Ra+cAefb1aAjfvgrm5KfLiVYcae5C9FYift/5X2PvcWL8EVlWxd2soD
ZLJoOehgai19hkKIgn2tB5irq09JuXwjUugQ84Nf9esYoC+5RPvqGbJtcNCnZn1R
TgkXXSC+BFKEKCXqmRnoZAsK0bNNMTypYlHaxtkKqmIWywod1+gyo9cXDtd+uY6G
ViVIemYwK5XqHVZITuYFADWaCRQagfaSFXVbZOkSPGMkmUbnf80o15SVUhBf9MzY
YDhYWr7A3nM/wtbOMdVC41fMgeoaThFAa7u41JieMqvBM4K1JC99u2meyww92F7R
s3ZLTAHclcj7HezIJb6dic5Z8YYOI3V/mGagczHEHgUBVg+pKtl6EzXCple6FDup
3O7hsxO3dyEQPSuHWYmdjhh0PZI0+G0sTZ/HEekR2+jHnajioM1NQdavEr+bIg8v
LAJ+EM6ENvWxmkSM+OS7oe/mnvoudtram5PUY8Cac1IhOfpw3eX2OcDVSDr2/D4G
kJiIoBU7mZJh6i4ys0hFJsMHclRC+W5xsY92awfswAaYkQyfwVuIgdTvAsraqwmn
PZBPj5eJmkZS/Sdf1YMCGTZCG53DcdYA9PkM5442qIP1TCo+cFO1AZPmMzq7SBoY
p76Wpzz5nj/yCOKCKLTNiobTDKeq7Q5sec029fzuPvu0BDbjLJ1Sw1JxOw+oZfn0
fwyPy4dB/CVKt0GD371JuEVWRHsGIvbE7VyLehCyxiiLcv2r36FkhOvNqRJ0KHvD
8V9grmAOK+HZTcrrRw2yvqkXiTl9+iiWbU+P7qAYTGzXYT+HyJ42AapuOxO9X9+W
pB5UGnUK6c7gOC7ivwkh0aDv7+qMZjZIWAkMy/jqBBUpzDz7ax0JeCaeQk7rYzVB
nWdjsr+YnBZD5AclO043RwY5ErhmNShMOiNvsGfHtGjXnmXKI89ww7tHvuX8TELR
XD6R74nXJ6Z0ZP4Mq3CqSloetisYjzNVhGBfzDblUpptZFWF9Sca1iG58y8vV7b2
LKAhL5OrSjwsmM3mnD5/EOO/9ijCNyAlbil8ajel9ranD+GSnr3mncUU4sg5z7KP
I2WCUiNjlgusCFxR7LyBwU2A0ksK6GAd0MjWw935dJj/zfr75j/uOsOJhFhwmAPX
mqY41RUFLnhoEuiAyzOCDVmEWgKhpuIDR2orJykvvOqS2pgMEBqEejyRja5WtFEx
friXQRBCnRgRPWr2b4E3s7tG2NyPqAur6FzFPKfkcZt2lna77AtnnbKDGIxmYdqo
xZJ1s+5/UOV70UeSPLUGDwcZfnVJUbnGsTmpjA4oNpTE3pbJj+ZiBUfKnFA6OqMO
5xL9/Z87lOOkGvcoYZE1iL81+/TJb/1wfUH9aKCSNiyXSBBYn2BPJa0vJ4n+qcrh
eGOdCrOafnZgfurUv3XEqgYrpp8ZXfdq/gEnmvOLxFR7Irki+LIG1mgocv4VSVFf
6iFqp0qzZTAnykLZpbuld8KNOXc5/UYbYlB8PziWEr2M0h4mhp4ay83+hR0W3Bdg
PsZLsvo04CdTWmZClVvymaRaOAvGnDGyz18EzTsFuiEMzJAsQTl1Ag/FZeLJJKgG
NOx5YxYZrx1Jo766oCKZOYDT70KRdl/IHT5mhBTMZqJqOu99I+Y839dH/Nug6BAd
d9Ge+6z5/7ayaFycRwNzC1iCgwCpFO27XJa+QPyNlmHxQTxBoWgwR4kn4kLfgOoi
wB/IGqGELqUh91h5s/KwmZp7C+yFnXVlAYDq1CbXg3NLo5g0UH49RArO9X8nSB8m
a6mZrL6aIIjJnmV3WYLt0j+nfKoH54i8Bc1zpCEcEJYy5+Xc2u6wjKKL/PyUZuEa
dQhVvSoiexKdk9kN2Z6tjIpuKd1wSjZA7Sb7zQWN6NMGuG4ngwF9O/8oj0eMSX3C
t36UuvveAjO2ZdjvuvOv7qOn9tAVZ1oCH4CfmVwTpqBQCMvrizSBxitHhxrr2JVN
YBEs5CwGM1Q98v4O+n2ELPomQEhBajMYYmjGZQugrKUvve9CLoDmbGtHvWXWTL8f
4bZea4aPrMTW2EKy16c5vMZRm2mk62YBcInvchKARbZU8/JaPt0XSY9DFR6Ae5Om
S+9V9oJ13YX5Byi9NC6fybQ2K6zQnywqfDk6pAZBVdmTywRPhg9KRQpMCDWIyxJi
+DT2ni+v16zLqhtEzgi87Lhictxt1/O8pB0h3UmxHj8nBMb5vk/s8Oj4aaO1Ky86
R/Wi8noBfSBs/0plRGeS0e/tpt9cWLWkgT0AU1gpXwdB0GgrXlWpeZk/2zwOA56X
u9yD6XqXqJi461//c0mdidtkoCVqDpZbW/dJwR6Kjvx2Hup8t2eXuMMK0sxgqQq6
YYYlg287bAlp6Hf4UJIQDYxYzhhA1CNZvkVWrsk+sW16iGeZ86SvMZOJeuPKSHOb
Rpr6rUtE/EM/yWMfmwyU5WT5A6ngVlEjSMRZJb6m6Cl/eiuSoGVnnCJPy/Edpaxb
LKAJtDD0F655Ap5R7ELqilekPpqjGu+UfD0UECKqHzeQWQXg/c6sgK94sFIqyqQI
j4RwVPt5IFcDMhSvziLIrpJYuIbGISk0HCS/Kwvdy9/rCY0iVl1hKuUhE69hMqiT
wW6+ds4NeC3CZm5EFrbZa/U19LD821GeyKfIcYJuNdPnMituwwnH5SFWmGr1NUrK
LUembaGoUhKw7jjqh66jdB8EEurGYYlsvjrZM9zG/bFRBJ0jEtO0mRwe3QO3C4Rb
MmWr8fON7fkmQ+w5/yfSug6m5HXJ0zHX/xfhA8UK0p6EI2kmMIb/E4ZwPbar8Xpt
1fWM2g6/HbYeAmYDnpKo7WvRZESkQFesYGIaT3rAWi/G9xO9lM09Zyg+rccoxSgm
j4tDC5IjbkF7fp4kggg+PtBKGDd3Pt1V7oTVDxCW2yZX0Ln7Katzr2Wm24TXOVAl
td5vExjl8ksUyUKBCv+CKRcQQHnyPBf0eX7hPDXTUXCqeR4UwW5nyl6hNDwBoZJj
9Gj5k76bw+AQk2c7SJGad3V2UFW//rcmS3UwLhCuaGS6+1Mo/XLQoGV/Zrr7G428
k4Fq+WHmdrpc1qeXSAO1ol1j9fMEeo7LyMimT/flhJEiI3EhcMkOq85ToLZyFIQa
h1dClnPC0jwISh2YCDqupohvcweq+XdxR8Aj1xdcVIdtQWhUiI0QsLvzo8ceaJvW
FL02hL/FifgqJFMok90NCacwzNs47r1PE/v8j3s8SzFVAmUtyLCW8YIu3/0WDAde
YAFGX+C42gGd33tRrjUs1X+lPPObAGulwPQybqibuU3qtvb0PcZBd52FrkQtGcvj
D23DYG+vFlhatxADAP7+PdgylIdqleeNelgbagDZah94UiACf6A4sK45tREQw0DF
3fJ2IuAduDV9NLAY4juiLqbiDjoYh+tjMLcIUhXR2igohSXYQ3cOluq5GCi+EnGT
NumVRFS+9+eDVWVKqtneaUtnVen2bi4qAukTSs8FHyqGxa89l5ElbL2FqquOZ6ER
7VjDu7+0Fi5gdriw2iEFOK5IH14YDFD34uDbEvpFQMe6sFUs9vUu3Kj5q/H6hkMO
OdLukI5dgsbaquvphkVcFvqChcutjiXokErhFm060pQMmVCFgcKrb7r/H/gpFI1Z
TKQ92v/XlHYwye917hiBN0CoQIMycL6MN+kvnbahX1sUBKGEyVNPh5GRUXgpiM0j
zQhloVJrgGCqrFB+yTY2yZfHDEErtdU3Q0+lFu7oscQ1vPuEm2ARGelCjCNXuaEW
n0EJSuMYQH+hdfPOQh5pxmsGlVyjNlECfFLShk4HPjTmDL2+4CU0XjtbCilPW7dM
CJFvDF8nsMRUOvLQOCc6hjoVR2UI6t/NMWrTnGi5sEGR+o7VkHZs3AdkRUPNRZAy
bGSKGzxZ8Z776gq1rRHyNOH9cMKO8r5LTe7IGy8QTh8mVPmfJTXKQcJDAVBvYtdD
UYFMefdBOLCO//6+DKIOTg6hLVr143GSSYzR7OJCbwiNGlHscKE0RBSqSluYWHM6
pUYrt0tMunjiYamK2INvKEzO3Ap/bYurxGqskN6yP/EoU4L3AlIduAn9mdDiQ1RB
ZcfHOr0SZ68k0PL1VNCGvOYtwY6RoYxt9B35xbgiV2b1cETVqgKU2qE0P8jXsh0i
0i3Goy95UQ0poPycaTrGpuo8UqN9w07os4kaH0k4bPzd8nm1wzTl4pxRFkoyB+im
qZQZLSIh/4RKDBhQcbFVgFd9mZI6gb6I0LAiOVxikUgGWfZ+Qt6Bi3/ZJLds5bVL
biC4Pv0wA4e+RftTCeanwBKdDeAW+OxOlVqzCL6izQ9rOEjHj02wJwWsrrhwrKAV
dYbu0gbQLJtL8IbllPd80X2bdzQb5sOzfDMxr3JiLRN729WVOagA47+6uNVLN6Gx
uTAU4FDj4A/qop8cAWZ0EtiSzpz9f6N8HIwDc/3s/f8iBcml5hJKp0bLmqCfH8RK
dEzPrTqBYYc7dxcuUeO+7tYwn5C0pRXMwT58r6xgfIJbP088ZEWoDwCZCQ9Ku3Jd
AnPzMTwmN0JI5Uk0k4j89LpG5VKnl4X20BTSbwYuYQ2amuZPk8993zM/S5Ww3kS2
8WZ8CpYj1LHVBHXRKsmaPw0eCsuQ02CapLoC4xADd2S0ixo6g/cxcgTnLOQIyoew
oI4igOhb1j3koRsPa6Ls8ti6EOVXRWUaCnKreiAwDEfldwEDJD6FqCQ4ofDVvC1r
3C8g+V7EPC5w3Q80YsiZ9TZBYAvlRFOP1Crhg32+GGdDvOBjqVEUZNqy+eA18Cs8
mOZtPlEj7jOdb93BcpWkL+G2DLibyldDip7BwpYdi719dg+32aVkLX1+fhbnbHF1
rAWFOhYLzRIE24J+HYyUgKKrOG+n9O5x2OV5soGtzF0h1d2jewN34K9pM7oyPauL
7dj0RWNSAto3vwcNi9kStLLaO8QTxoJr2+QhPH9v4duJ3A7qzYltIv6xxmD/QSoR
KHXWopRY1+CgGYEfXdHtha6h2bjUgK9tdYyorXr6ENlW/277OSoY8ZZcTGMdXfbb
YlY/aqYmnoknaYBYknwsNMVjFoMJUmgXgucyPun5T64XCekh32rVkUq05k2fmF5t
ZjpH/JNZPBBXhfOo5T8Bd5671JNgtDmGHVZhADIXBRhIVcRjgpbT0lJbHC41Adsx
orY5zae7ILbcuGA5OiBS5DxmnEtTML0GZ8fONtjW0l5VMNPFMFSaQWqhqVJQD2S7
fj9zqdgVVi0wmmrL0KvjZBrYuDTjAprjSfw6Y5HuOgSQaDLxmCY7lPlMwIWKOb55
HooSps91opzHZx59D9QulA3WXp1RqJ12fxhvYDGvLmzM9UpIOk/b//e/JLyt+JoI
sxNPyv8q2SOoeLBEm9DYtY9Riw62WnH5/ijU1yKVXCwH0dResVMUG9tSjPsT13Dt
AVHT/COFU+fNn49uJlPD3FoU4lRrM+67gNDLLUoCNTTqZBSrKowq2QVFnN5Ecfvc
gm1tA4V2ozyh/An9NJxaRk7UrFQxtIkujLnfxeNfFvPJ0dFu9vD9reddz52uKXwi
hqANoP6LLtvKqWNUXRa+tCeQ7kcLB9oal7i1ixwex/PA5QKXzsF7tWRLnjTnIX+W
hxHq7KmzmhEjJEGCsLFqEXAYwg9upWH62whzwr7+QYd/K7CJEixoJHI90Z80DWDc
o2wrHwOBWp87tHRP6H2QxK0iNY49cf0El2bK3fG3/pBhmjSm4gTgZjMAkIfvJxkL
1/CcMLL3S0+1fpP2dduP58W2Db6e2ID3HE+Ox7gxkbe7EFCkscfoNTZhKw91zFuI
yoPWlEM/8Cc95ddy97YL6+wmStDnypZ1PRs/b3o6ZSP5QssaJnh2/H1Z8Z3W2kRV
DXII7P6pb0vmS35uOWJd3IK/5UEAhq18knWAjLFtaAqHqli/VzoyJr/hn7zIsTg9
xhtCtZM/xIda/KkE8djtZaN/SJbi2AXSyyUJ2+N+JvdzA9S9iO3+zF0SbmQOcoBi
hgN6U0TZsCCftJ1rRO10p0c6W8B8sMAtZQ3e3CCg9acM4vK+cYI1J+jbci3mK/FW
e/vhrAc7UZg0KMozUfA7W4kcj8qkN2EwrRVEsv4jIVz1Vb08QyP8qkW5WGVSAgGE
8QhoWzuG4ETAcBaVyLtcdbku3q0myByEpCzmNAk/1YRzq6iGEj38v+Pg4/vu1CJT
y8wqtsaXtFOKgSj34Qg7FDTaRw/Z6mCRxrPcSOzGd6wMyS3NLOxEGHiuQ3IOjVLo
Pk05BDmHzjJppzFUEhb5QunMCQ/HWglu3yNoHyM2v3boYjF5euF83EKEdyGIhRY/
gGQ8WNP8VsE6x+bFwQxG1rvOm9nj6lwAmTVrljQIoxR5Jv9uQt5abAupmKyssOJa
sWywUJTyMfSIjqXzgryGV+zVI5hJF8d/Ami2flxc7mxojyv8nj8hJOV+To9KP5WE
FhX4V0e8kJwugMSSfujrgkyzT/MoCNRmG99VGFTtgcF1WM9E13sq31b3z35dqosY
eL9VsaQaK+WTV8IVOAiazoLDcxL9xnvekgotHW+rEVx4nb1RwBknXPTRj85nLvkn
spJjNFO1IflLt5A+d+fYku1x76Wyu76Hd4h8ppfvBA8M2ioKcsfKRAMh9hkbLNrj
yZA1httQ4+Gs5lps/xRlQlF9d5nyH7KZ71/FcKlpZvUGhPoVnjToYklXv270Ag2B
Cb93bE+1HKoJ3Upze3rtjO98avwzYemE5oZ0ehkLmYcIMETAPC0nELNzl1+7KjtE
fkgxjWw3eFpvH+0EqX+PVQ3S++3g/GmgIdRM+iuy+FHSN3CZ+DXT2oGoCxqPFy4+
EOdm6CaNLaQGM8RxPnWIA1Llr5yiKv6AifvS7rgFOHRwNHJt5m72RiLnluLvIRp1
5Mhi0KYaktcIFJrlBTTlXfwuiHDmwEPqqs8VSANR8c9CPbJdkPFGDRV3nQmUllvB
4gTZczqin86AIHnN1vxVX1ElXizK36+FtEnxKj2kdR22GaJAzM3IxXUzKyB6x2OP
rab7Hp43N62HwK9yiyrVk/LMoOReVNII6BwUo1+V1S5wWNCYmYhyhSdm+5ICun+O
fDNGic4HPufQpDnUFzDM9cY4/5gWm42ekjOTxJz52enClbwgMZ2+qxPC1fO9KUha
/XiaohZ88fm330Hm7RPS6ZQtl0AwVOO3g3Bi7z5bQDUcbB6abbjs5XW8S/Q0PgQd
eGFylGnQ2n7k+o+MdWTFTl/DlVA2YJmClvuY7C6+seRDtTc83BhbWq9dxkYB9iHT
2NbnYMaxh7eMb96qcumTumqnpyuIn2gfjdjl369vLg9cqnzuJA/NIRffEHNkbwu/
ZOs+ku6+wvRG9c+AUoeAWTPETlF3zvkRkand3Sr07NmgjHjKaU6DadVBAwU1StWX
wG7io//ZFbQp56MEYxx/epdQhNti++BKL6kG0b/7IO0v5udIFpUOKwJfXhDFbcQo
Z83YaJJKuOgMuEZldxl4nHJnyFevpJCNzGDRQ9g0Bedwh5ClbJQzTPTSJ2NGsINO
cmBA+126zB6DS5iF748KQewUVWnqp0pwHjkzUoVWgU9pZHURD7nO8NR330alH663
m18sV/Mw8QF6kmmmJd0xK5RQrL7rPiEoPVdFqXWWcRtQKiSV6ldI3ELQORtCh30Y
ZbnwyygV1y3iBa6+kFSE92+Enq27izJKC/J3Q/oj7N5t08MYF38GTJ3woZ2jIt8U
GQJhGFcZJAWVxS4faevQllKK1TxV1/0AzdkOZ9Gl28J+O3vI3Fr5BYf4icfCCr23
CIf0HuEuFQYuBKcL6JcbSjWJypnNRZ5j72sZETtembSSZr52nWcgnnFXO8/d9AN1
juIsG/u41mhvRtHCR2t2kt3WE8ss+EQ5d8IGsAVD8qQRuDdeR0pTiPZj2zXiYTwZ
S2/ryO9XX9+ixURRxQbgS+ng9qS7MGd3mLby3+SMhkOgkT1hBM2eXXyqIEVf6ts4
k0X9Gqb+SwxlBY1jVKTmFFFM1uYwnEHJVc6wIHrwCzrRAzpYCmX1Ifm3+Uq/HtbH
MR9ZI+8TfAIMHF20jnOC2k3v3ezN0nfePlU3LTKezWEaybABxv4zKAEiJF+G8lDx
HkbkMvjaPrvAKGQqvGCcNHjzZzkxR9utVS4QUbH0pjwJnU+/KDzwigLvWk90YvvZ
GOeVhZb/4xs2IuoKcgCH+uUYWIK47vnucP0YT4T6SD1iQFFLaGAiew/8GiGn4yqE
IrSwCUCVfVrHLDEG1owBokGed/PDM4OYn2ivR9ZYucjnFoFLggwgigkDPXmzPPnx
b8nPOY+04csTpb+O2r4YEhaB+98o5MS1ySb40IbQBJosVlsGuadHo9pnT76fsg7v
0usUqPmZakKfSE3Da5l4QY9jXN5KLVA8fzbwhRwHm4mLXHaZti2LJYyzXZMLeJWX
87zk55Xzhz6TpPh2upn5rxJ8S0V/ZZf54+Sf015EaOZzvmLK87zUY5mwTU7b9N4E
Ju7B0yt63yz25Hr/ccq1FhkyShyJrHUSp2X1rBSMqe6bcFM5fS5ZeEMQS679njp+
KXw+3bUQgIyDcrWwkWPuhwRczdoBwn4RK7EsV3pstaVi/TSawG+AIGp0iOHPIJ+Z
FMiQSYfiSAu6yxXM+nlKemxFafU/HEx1J24p7nbZAFOhW1Vxt1L0CPeaQreApRlM
+0Sl4h/e5XCYa2OMIdpzM9Eo3i47EOOOmRQFpe5X8MLbFirTxvIklIIz9wnS+AiJ
uxhBem073UyxpnOEqVRIPB43T/4Wr9B2kk4ydanm1ruEMbtPdzO97o9vkYJ6M1g0
pqN3suVK2arniWyhROFqk1xUblk3Z2ZWldOtEmEsYQUhb5Y6QFXSTXIE36aK6C75
El/vp5p2rn65nvI7VDBUIfFHpW7aiLE9/0pW13DmF4ebIfvasKJ9OzqaSnoN1KEB
wSg8CJ/ou/IK5w+/FBSqsB8Z83P2c3Kg8DwG7xQzmdLZG07PjwtU3VwicHS2YCyZ
Eofw9Hm55nda1CY5qBokIl/oNmciWIVf6pARjON8G9SDlaHH+D6V1bNizncz2ZCj
uK0yH09tafrNxU7BmZJivXkyb1zQ8C7M+T/l1RkyP7sPPktkniuMMkwMPHf0REgK
jK03m1BRc4Bwi8Bh65UPQUUe1oYUR1rRZTaT2Pn48ELSPET7N8UtdQi9pgy5fduO
MGxp2CmVbtfssZ3D3/SXPZ1pHpuu9GNvfzV70VpBjxPooPRrqzVsFEH8DOWHxwMy
iMvns7J31Jgb+9Xshi951DDBnoKYX1OnZz7TwGmJv+Y24AeuSdzQOEgLKgyO+Xtj
dVrT0LJliHt2s+EOZiFkE99akGFAjqEkZZt7yIWth5ITJ6JOuUz/m6U3770Uu2L4
u1+pJUgu1o6Xmy2DWBkOqOc30iu6iv8rJvZ8YWjr03UZwI4rTXuL4xqCWahXppOM
rRop3WyCSw4cwUjhqUV46wxSsfHUwRrkKpkkOPSeTaYgMvv2KngQ2Pc0SlRGMl1M
trqim3fCpHaeXfO64nBIdiQYFrWpVM45J8SZE7SbhqQUZKmXUvX3JFj1igq+b7p8
OBLhOoo31ojpZ/i6nv6rRF8sT7o80NP+/S7tI2v6dpSg0EgWCqPs4OpL3PQ+SeVN
U12DvRzZwga+dfadeU1lwHNG81h+VoiXbvAQYoBC2TQQVmQiwBURR1a6/xHLdaon
CvaowuYcAIpQo7He8cZibHqnscpCiocqN3XMysBBFp4flLwiEb6hs9SzHrtgvHfX
SWYygKnLeINivg4B8S3/81yWzc33/IJurBm+/RsnwE3fSK4NpN7IoWlZbmEjzu6S
IwqkDh32fiS7gazOrCFZ0L318nQrMeNEZO8vaQhsoCQZtBLzNSWByoo6IB5KJL9A
AiabmwbVjsO6zvaao5Ambnjag2jOsgZJUp3P6hk/GrnE9IBsZQ3zRQro7eTcKzF0
RISZHgG/T5K6q7gsWVOIlmmnoqz+rEeqO8WjPu6TtzyQbQ2M8bDefY0lgESNchEt
0MHsMbI/q6IYxFBrxDrV/AFOZeAcrITKimGqo+5kmVZaZ/31niYz2Cv7oMI0a8dA
YdNBjVlmLsr2B/p0pZukTAtzEBzt1QyYmybUtKF5Y0jGBCkwHY/dDEu2jr/pjaVx
WPb5KScQs3Ktefqyb/QNQgs3qBHmPvc+c0c22DyOX3Rh6+2I9Y5twPGalwRjKPgD
`protect END_PROTECTED
