`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OmNEaYDAD51k+rLgpYRoX0jcUjK2Bi6QJJbSKXEWXcgmg7iOI/YqGe0/ogRosKS7
WxScSso7XXvPLxMXrIiL7rOsRCvIfNTJz+YX6fU8Pgeb8YuLAa87icvzFn+PmP2o
AzMgLps2Cy2esBBIHgiR920jwxedZ2lcUBvzywHECXm7/E9einG32mcJUmDSspoT
1AOJteun5bNohTeh+/iSTLWnFJ0ZMrgAMTTAdcXL39omztHqfQLiFIHk/kbKqIUa
iUJww3ZmZjnLYUoaMlstk0NpbbCcMY1YtoKAYkKS9Et9ppqGJtyndKtCfvRfgf2t
ca498rW5g9DmDHFhlNSdBFW2z9kzP1MAweBvn1I4t/0COWbIJ5EmrEMQE0Ykb4jy
MtoT6FtuVzw8d5vWFCyLvw==
`protect END_PROTECTED
