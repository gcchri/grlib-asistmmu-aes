`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o5ewLlhNsqpskmz4MNlm3X8htu58oOm7CsWMm7S0nFgap/VYgTkRpafCiOB9oBqp
foyMHl58cbpV7WWhCe+LfpaadbVfZE5kT3eQ1v8m152nYeVL1bwhMrNSMPm08Zl9
BoMqBN/IrUgT18LikYjzOVJX9VDpubZficQxM4VHOXHo/hBzS21atGF+x+Qxj4Vn
RBwQ/77bSDd8qUJmc5wpixUfXUOWja7rMgdzUj+EEZ3acXeDzAwanrIFLdzz2P8o
MVcMg44+vaPNNXhRmJhBIjmHOU9JrlXaiCrbJ0djcP8=
`protect END_PROTECTED
