`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xhar+8FL2TVZ5WerNT4Ma4Xt5tWrjXJ4CtHQeAjNYCzxe+Dm8mTyIcGhYtXFfzQ6
N1M4P/zSf9pjjjxoqETeEFLabU6QBBjv00wOwohcouWrWtDV1j38Us8bRuHdwH+N
otAxW+sn/Vny94WVilrCATZ8yzsesHSqM4YcGflF7OJhq/FhAZ364A1iHIjT8aSy
vGIXhjLpNSfqJ9l3iAWBdA0o1KW9GFCCwx52QpQEs24+Rcpq1Al/yRlcWCTXnuee
LLXQokRTMk6va/NbCEdZ4MHycIkoFNu63K9NY2gWgew=
`protect END_PROTECTED
