`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nmt0kAthk5kUV8NYC3dgyZFUhdr2wteY8KG/IZqt6ZpkPBZsrFz+jww46j4aV6kY
7mgF+qedQW4TQj7i9PDvkmvB1Jpq0rL58wo8kiVG5QFy/su6jInph4nBgMadqFvc
2QoqXsq2+eOngo1rFSpmhL/TTYLX4HU4aHazriVUOtH8RwY8N0KjJGzGSPAA0R88
U906wWzyVrO61Ujty2pOqwQj9Eiff1I8moNn66SKfkDwLtC/ng76glpuLnpdsnpV
oNQZqWwrI92t8vFzlCxBAbzleH+ilneC/F65o/bi10cnjOdUy1MdnOyK8dY6y+CX
Wy9zL4k3t0zAeFhCbUP2n3iOE7ZoEFzO3GG1CkEW83p0eJaRZ4SCKSqgCuD4N7nx
oNxBD4gE9ZUSwXulAUNRTYLQD3GlcIk4+TtBC238T+M3hTyFjRAnTJWgtXJqy4vQ
l7ZH+KHSaaCEYU1Z+2rVu7K68kdyYWOLC+mjwszSja/UhOqIkN1CGQTf4PmmQDp2
2P3IcZ7AlYT6hXZER8LKAwvGmbkw3LK4CRZLpnReCdktk8w3NsCRJmttpDDfg3cS
HFcekzfwfOQy8j/6MgnW1vIhZmozkaMdYLcgH2291nGyCGpt1hCm+Nf10OeP15cW
ZXR55jAhHmDzjBnZLkNBXkQif3qBwJR5GqNzrkrSxcNHgXLWnfs4T3NRXTnejBhK
IYGf960If8okVyZ1Afr318E/ysPJ03iqj1LzKqkD0upR0/rmL1moe8zvSx9fcRba
XwcAe07hyXZK6myY6OayoqnZkltPkb3+38/l7EdV9barrNyXnR3MSUcYWbF/lkcC
OhepYxkH1civWz6X/zAxVo89ZakeodY1AtkGmAAoU26siuLDYikkGDtK87Upu/Bb
7BMJWZetY+CVCfV6Aft3NFonYrwdrHwp5ubYWiQUHKngOV2xRvW13OIo9s4qs0N3
DiAKxm1pLgunWqJwrH+A2wjNZuH52DRwk4Pwlg3yEkGosY3G1//Cr+eFQDkSaJny
jRfhT8sDuUR3oAcBsRye9k10HsH1G7gJ9WTzcHmNrVxDkXp+iTbZGw64Ioj9kwF8
P2NlRG5CAuGyxPGpzIMkag==
`protect END_PROTECTED
