`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JDnY+XzP9FYe+FSqMFdpA7YR/EUl4ToN61xrU+WK2Rape8bea6bLmZdCo3i9l/gN
ovt6RLq5UL8UiWjFfK3/av+KxDqocay3HqmG2xBJlGmqXZvWBfqqyo0t/uKyUK9O
KKO9rQeHK2svtqQtwxYOa7V9yNwV0X9l5GsjOv0DrFNR6NOVkwOZjPWaRB2j4Yqn
07VBKRfvIg9JMD7kdj/V2i2QOAqFq12NzziI1BkcW6yT0rmLoojQhHNmG2kw3sXT
Zn+pDDLxL2XZXhDGCM02Bu+wLTJkBfINZ87QdxzGgeXbLl+w5vI+DJSn6G9vJ1Qr
qtbwiOfrnsMeQjA8J2t2zmAVDqedqVuxapWlQw3RtDO8TmodTnhqDPeknv6WDopu
ipeVzmagwVk2rq7x4g9rWqkpSIhz5RXll1T0MsplZlaLz05sXyp7RlqUeQNrzfrV
3BSfGv/+vtxqkoruug+0oeCPZpUJsrGiC8YMGQMM4QxqL3ervkBLuvhQ1N3Jblth
T/ankCwdOon63LKlDZBe7gJLAiBBq2kERgMkC99vmkgx9ty2+MYWIbwz7rru/hQC
9SBQ/Bi/X0Uzc4XNBSgOEiR6ZEqx/sk3PxRPu512a4ed909pYuyPqpxjMM0unFxv
qUIMUAUStPpihvdIWjYRl27b06okxsgI8I0sG9xRwSWUpfIh0qgJEOgSVsLNAXvl
L1STSgROCYnAixnz7WpLLMaTncr89gYW+NjUSTj/W1BtX+cg2NrWU5jvXGjms5Al
wCAF6kwKw4tGxBusl8wxiBz4aYnt7hRhFrUfO1ThCBoEutOlrHndCE6eh61ChKAX
ASYqUv/tn2TWFQ8NjRxTHuhbgk2wq/PTVkzPFLXojb4+QaEb/jCTHZEntGXeNGB3
vJoEyaehbuFi1ENPniYFzKZnUkuMvZY060C6EhI4/p6XoGIOGPMUD3whES29PKMu
bBMprzTo4M4EHH8qSAYPRlru+MnKVY5WBn2NZtH+dUlTb2BNUP98fx77euffUK5J
D0UD67CCFR1sTUWMUi9gsLyykC/2YSxItk7zJ/tuCL6NflWKgQrMIatNsQbhSaD1
wfrXdVtU0ls6lz/smbTeRY8wTG/MZJ+bfiz8Nq2byfvhNAdTWT5+TYcS+8wSv/ky
rRZFz10y12R0CyH2r8IDpJYKCpXAMkkx92rVuljMxcGQ1jImLbqBxaKBlYnY2Kql
070JTeYc+RJN3L+85gKKc8JKj8k9Tn2futesxdvTNWid8c/H6gRLPvlYkm20zZpq
GIb7WNqtQ4J89SMp49sZczLEK2wH5eaHMq6Gl2PIbY0Op9TpT10PRBMLne1cVfNr
SpAscuZHrzFSpE47I4OhmiJXQm4UE/USzWWw4Ux3Ms2XhhIpTPuHJgYey1XSo47v
F5cc5vr5UlL3T+tS0ytFmTFTuzkpZfJ1AQrXUduQljQOcJSUdpmVifGAHhrp6/iy
23/LE/TV83qQGK2n2bskscMlyhTeppkzEwSSKDn8PBWj6jhO8ZG6Il7DsaBS/B1b
K6ytj6VQEHnqTkrzQXk4N1DR2Ny5pI6jIEmDWzvIKrjgePXbribD776v+cLzAhrZ
UZvIh/DpOL8r1l8aTMWz5IhsIUN2XuUIYinl6NrlFl4bXhORZUbk6GOo4QxQuTsX
k8yj5CJxMFGKsDWBuEOc3Tj8f+MzixuAKU97SLIzTWoeCSdUoHUN+uccCziNcKRb
4iN3hU6F2P3IsNIhnL+E/MIccxqnK+sY/VndUudaMk9aEI3HNnX+tK5xGoavzncO
XD1zo6q+AVGlVYBZ9gEkdQlt8UOSZJtcWxVgpuS61SUyvEKtG6SjJXQeItOMVyur
p5VgRjIAohDbDawuCe5G6EEvfXewWCOFNzf0W08feQfZlL2W0b9QULEWq8KT8tGO
DSkF95h8rcfKZ/SPw4lr+IrEnFSa9sbWFkqA0tN4kDwgBrEFXq1Rhb4+eCWWDRK2
YS1ZOEe6uJYkK3RiONgypnTEMvxIxXuFKfa6U1iwhDm+Y2nLYMVovAg32OPyRwrR
aCS4VThDIBgLGi06eLaOW8NQS6LmAYaL+1F10h7Bk47YKa8jFtaiLk6t9uICyIDs
ASt7jaLReLG0V4SRK0iK/uxEs/HNunLc1fTOE6W4jGqKmR4z5o5IiEWdY7m8K6ha
yFJ/Pfl3xrYDI0CowaCNzz17iy8ImAdMZ+XJd8JdB2N7PL7w19lc8BltvHbkhuO6
KpMIhWvTbf+oW49wa7aoy3nsLwVXOmaMNezWoxBVRFkqC25ond7W4mQCoWBLIkTV
`protect END_PROTECTED
