`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Qz7NeS10THKCOF95VWTxZ4+aAtdj3CuGzZVkbUOi6SGdhBaVmLGAys6s99p3Osy
zyOd7PPiG5hIIlINg48SEkvl3RABu3BAnqLiZMWFIn0KZ20StczsvZ9GOjsOslay
vUV6oPVHF5yfxN6tEqSRm+lj+C9Cc99EKnNzukx+vg+RnR0EoVbBHwI0JQP/AYF4
cQQesdAxxkygJEjaYPBJffFIV/9Aw6trBzKMUKp6DdYF6Dqbvb9qt30mMWuXQqrp
r6aZNg7bd9pP6FST5w2HsNkw1yWuybv+8imYAt5BnshwYNaaHyqvmVa64wJGNa9w
hpzkftJKKCkZ7RroO/DwCYw55pNKJMzV1oPIeSzh1ul0WEBpdPy5aOPNZA0N0wDn
Av10wuR3dbPvdtWna8oJdAxbIJ9FGBd3lNa011gUKzRDljpfxnV9xoA3E818RaGN
HYv75TMH2LXRyDr0LqCNxDBiXF481jTYMnxMj76zeNHaV6HVX+tgVOimSfokB+ZA
xo0bnf5Dse0jfVN1XwL/k/3YYnwm8n7EDButdflGjZJoyvzNosaNfOfHmPh0qXHi
YD3CRvPsUeJ06tGmfieX97wOIxi29tlr4LDO4UbT4V3RQnZn5ibsFtpQtX1ygLsa
oid0UljrFdwWaLGfjVzWFi9VZ3k1p5DkwnNYX79VPzIEWhrwRi05TFY2bEzVfoTt
ex2AVYMHiLf+EAqRp/XN9mXZFLD9LrrF+kxQZlhUhkJEV1jWawslDmGRbjojmlUe
dHtQTf7zERQungmeYGh9EA==
`protect END_PROTECTED
