`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wxcYenM9AhvjQb1obsa5FhaEyf8JgBO6UwcpN3r76YbDurVdRHkmhwtlKVnhVi9b
HxFJT3U+Nnu1suFo5NR91DcixrGXDTmFJ7u5dycxPpiDwUWpMACh7ZOr4Us19cvh
ExzvYQeSljE4TUg3bYdU/e1JmGcMgISXOuRF4lvENMXT/y7IXfW8I6y3t45JnVbd
UTRBHCXcdQxQPoB1ffbiNC2pGwdCkuQ1hZSwG//EFiJiAvSTU6pLu1j0eRzPCCS4
LlWBngZQOWU1yU/qm7mf26rZnl7WmTpQIKv3Qd4mLO+2jIPA6MCo8Tg1YjtgfvL7
lJ0/r+I3QUpR2pHpIUXys6+vnbsbC7rQJ9Z2P7rT1LhtmLtBhq7TUgT5FGK7LcLc
SWUXSB1h4gJ0SkfJrC+tF0hg8aD93NRyPLz37CL2vRM4U1heOe3ETetqqIkUDXdo
sHQL0TTldkZ8z3RriY024Fx/FrwR4I+zcTcKqi5fil8oExTFPYUsy9iQeVVPKhqv
rRqTpgi7/A8N1SFHk2tkoAHcQz2J/U4hhm/3bnqUPYbQNvaMvSa42OcaGXFAZxlR
WiZOYgGY1aF5FAvAu/WJtRIhFPa7EAnVOyjCEqs68B25Xp6RTuaEs3HBlrbgkjDs
ZzeiihRaMkEMlOEuKvD3dof07UU4cngU/iKCPzu8YaSfHQELUp3uhzI2VL6HQgeS
vruKfR8msdvF83Ziq7s4XcK/47n50a7V6gfXCy5suZ1xJ0A/kl3c/6OefOd/j7Nf
DSRE8HVLKJRGss75282BA4i44u6lYh8gxdLlhxaFgpYuZY35tYMYUA2/rq6pqW5d
SewoMPpNMHDRwdlQVfxmJVdA6hucm+YEJDyL8II9sxRTW+ni9NnkQO14BjM1IA8u
ItUcPa5mvzMq52kcFk8AgfS7IP9ew3a0WQaOgCYnNdgQOobc9NPcJ1P3Ec1w5d5U
E1b48ZNe29gffZquTZ2mbIXWCFSFuUyM5l7rlEG3nju7XvNVSIwBd65ffiLkHbhu
zxOKhttGc0o0q5GUC2bF9RyQ0OTJhwPLCLQmuiZsA9AzDX23XSn+R20S/BcwQq/i
CsYAsEtpttMgiwApP8RYcsWKhoH9yjUO0cXbO2YjXnyy/bSB/etGsb/oHofKfIlQ
szHf/jz7jQ3nOLg/jmEys+wRyUJMQiR4ypLr2c+osuqOSIQoPOOLpmmVlJdaNrSn
mfMh7Twup1bTA0vW+q+taX36JEW+kWzfQgx6/QrlmmpWhgu/oUYbKmHOFPLxDi+p
4VmtevQU2nzSiUjWMd+uTfo9cKJpd9KPYTTmKzEm35AKelsL7cupBe3L5dDZI6VI
HlIoMoPCYw1qbjmWzGeSwVdaoTwPsHN4UKRN5rTvLoyrdcTCBJ81IPCJh2E5gXNd
a+M59XAacw5T/wFKmnIN1wcGQylMLrbl4CkmFX1qctlZJEWUf6f7rx+TyvLBhDFB
BsmdW1qJIPBfFLxzbxmBe1gMsphe0tO/K/g3uiWEDgzLtI4F91bcqFA0B7eKQjNA
gtRKOb43UwioVZz8IP1SGYxDT0m0v47s+pWY8XKU98yhgmthndDYN6uHl3E4WJEc
927vmudbcXRRmvxR5sug9t3teIq6F7XfWHAsiKrJ1D30YcIQik7B+i8KevyG+/Qx
mkSToYJyHvXVCDn4rz8o3K+QG87uuCw0E5aKZVOw+EsTB14WjJ5vKCIe/+JEMU0R
qYbIhY3YtFCiwFApNhWjoB4OJVLSQstZruyLlvEa+CKQuUfp81L5/FT71RoCwgQr
zBMI392GqyYbuEvKhsTK6igQibsVwGDF9Plo1Co+lhJrjp/VmbmXYrumcKYCjGxF
R3lMByrA5PDVfjG/GYczZZLurR1Rpsag6FsYZEc/uRT+RuW76q4g+bZZExNt+OLo
so7Ev+wUBH1OGtmOcmGdwsTMwtZ37vkLkaoz2PILpmvWiZEqO/yOyEmpIw/dfJQH
iddwVqadV4maIXH8HSueVOGwg+i908Zd0ESEAg8+xng+H1/74+dD8z6TJJTCYAOR
XRhlFttpTBx5Hjg0rqcXmVXMgU6GGat3jyn5hpTn2ysZPCh/vsRqGC4IS6boa+d6
EsaHZImp+lflfeqeYeZZSzK9gLR648I53+5EU6u0hHceYc2+3saShfrPU2pqyB9b
pD05+cW2XX770PELIi9pldWeenLCi7MtTSbDDWToktCOJ+8cyYm7lemWbfRe028R
Es5z3YR4rf0hKi6lFRoNDJlXXW5bY7u6StQHZsHn9AdKywaivcLo2yEDqNTu8iXS
kFD5vBu2zcc5Rdd0b72pHoJsnS9onp3KOvqXJPJXpFCTuFYRBKUxxuq6bL266PUX
ebQrII8xhWKyL4qWjGtvK7tXoF6qWTi4bXTdDXygw5Wwi2iDH9n6JTdHNM/VyYdk
hsprz1OAE9QP9HnIvXu516pWD4Chi1zYo1TEMmnGjCe/BSY2eKpL8ZWZ0LKrOiRj
At0lakevWdoRCPkUnkwvxsPs7mMSpSbtwsfnOiIKuZCH/GzWESTYkx1qqdzllm8z
kj/74a5Gkr96lkdDSQjmhPAiS3yOvlcfwQ5V+1fmmagYrtDbeq6CoHpy6JQHthV7
rShTdCAdfzHapmP9POM7qDVJg3A0qMAUFnDoASs0hvz8Hd3Lk+F5bFzVdvnr+pB6
CKLA2WQuX7SLcxNq+AMAC4EqUmtvDPAP5DBVvryfb29Q+UFliFvb6nn+Jee9bLeS
4r3utnm141fvF/1S2OZhGS7eDWCEf86UEvS+KGmFfYs=
`protect END_PROTECTED
