`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rUQtfKZ+H1Egae5xviryqhQL7qw6i2rCVBT6Wd7pgDqvR8xtODv8JRaXsoUvFUBY
wWsS1mXv03FQ7j3qbsLMlSy7bo7Mz34qGgsLSn99KhdlIwA16JhTomUvGFWc12NB
5rZIYe/nozJUHyhlfM7g60A4kj/Lj/iAPbq9C/kChbRouqJWXC7x1Y4ZmJTLEnQP
McmjmndrKN6L2HTd8RJu+Ui6qEykNQe3sVF+tHnOF1f+Xc7FQXTvcDEaW2bo083+
30HQMZC4F6YHLI/gRBGieQ==
`protect END_PROTECTED
