`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EjMDk26sicrIw4BC6psC5+bRzuVGPMgkNpVfYsdPb+0YZZTXRtXomXUgnAdJgdrH
oclHSi7PAjFJXdNfXxitLjm8/65xiQaLLqGHnz5hln4Q+mvW5MmYLckDg23tLOEs
UvddgvMEw4Z/GO9ytSKksbKE0R8oGaMcd3exKGDl2PGgzp8PMZHiFJwJf5h5B91u
XVmc0aoULcth6fiTkzRGa6e83MFdzLB61VahLYLyEIU6IhH+EZLHlxy2bisW7tD+
rrvrsuedngjDTeYqtTfwvbjLhqTc0EnBRO/C9lzKuA2LgrPozCJkdQ20mRxBwCc8
o6haMRtn6tljIr6E2yz2I6rpuYqFmHEFB+qwugbaaxZhA/9RzmFE9wXKOdd1M6nj
32CPMMAVusYbWAbeeBCoHhVNUKSAEulM9xj10aTo2g7AbeiRmVGlEtxjXjRWYQAg
ubcpfFRIVQMkwdC8u4dXgkRE3KDgCfqf6mL/MES5hxe/CWSzrXBeMyEz3T3ChmvW
r0sZl8+LvzECWfUWD+Ka8DqHEHzGWDoGC2FSIdBA1bitFXPSqL7sNpIE5jDYxKMQ
hIumEKsHC8PfOAq+HCWyCTBvf0AhLl/l/2qu2+sdapBoKaMvUQ0fYHMGiW/VQenv
3acFGIz2NKpScwbPqpE9fOfQvlFoAfCa595btPHXoFk7H44zx9k57XYie+EoZFd0
nz6fDhT+sp21AOdXQ2eZB7+cqKv5twZ7JYUi9rLBzJ8zi41VREcIjau2YUA5Fr15
UMmqvPMpoDHPAp2eJbvRf5sohvtQkfRq5f87UMqOHC3UP3IakRRvo+feW/q+4TvO
Z7q8+nIFU/nCqEpUx3Dr9jkmYXPJ9cqYA8rR1BUdNowrEC8AQfGNgLU7DhV9kEEZ
I12JWhxWfrOPBpEzBwQi55x9wz7YItiijs4EfXcZh8Q5b36+qx7VLoxmXDJxSSGl
`protect END_PROTECTED
