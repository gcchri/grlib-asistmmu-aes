`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V8/54ALFc5481NxrTFUdkfaSJtukheVHIO4RVfZ+Klh0llwr7QYgRT/Yg9ZzXPgq
NdU1OcnNElBI+XaHePXk/3HYfy2BKSQ02FIKgmj2FShL+N5gu81mSM2BjWnHPVLi
sF7z8dbSeqgE23ubg3E/edgpuD8VkK2PMt5cbGw1nn9IQRUi/XslO2Ut6u6NV6+5
tdI9CgoBFli4ehrADyJ0IB7Y1HSI9GDQrnTc4RfKs87y08KqYMwWMSygGy4ZOYy6
D5KAWupIcf0oOTovdIotoaWUln/KNxXlzGVlsFoKgpM=
`protect END_PROTECTED
