`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iJv/x9BRBtHIJWvR0gmtGlrmM6JYVhPJxZIkCOwCYq12I4+ig/D8sW65ogcSV6ZM
D7tdJ+MBfeGLfRxlccB4WhkXgvkdy71BSNyx1o8vTvuE844G2C+CdHWZIL3Z3C+j
W0/OnpRC0Mh53BCYk/YbLgeeZTIFkh+HKNtIcHXCGyQQTJalzN6aBegfQtvzmgIF
mn6XXymFpVlNPW1OSiAGVDz0H7t9wlxgOc3Umm6ZRqrKD1NUQQuG25DMKm4ssDwr
inFADYLZPDDU8p4VIUQrdDuyLBMzxbh50eTogpv6LrY5xzxflfyc1hMQgfMT412L
DRAHSW7u+W9f95OnFuT0mUZsl1TjNXDRpJH4jHeyliYKpaOZL/JFhtXGGpFHJ6Ai
7pAypgQI0nc46/UY0GM05A==
`protect END_PROTECTED
