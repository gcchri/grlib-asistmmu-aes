`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pb4bSIBpEuydr7zfewSoAj0pM0+Ts5Ma2eJDr+dSQcRS5uCIsxP7nBj3D14oynRo
0nWncvE41tjzYYsFjEiwlpYarJqmJOqI3fYQEOLHM+npsgbWGTYm4TbCmB8V/0zu
2tE5+0FQtXA8W7MVgfY1T9WlZKXBxkuAzfIShTv9FvJYXFTd6mggzkBWo5S+zjXc
ddc9fapd9sHPnJDpaLDiz5rQS+Vb3WtpJ71T4YaJy55nKmG0jTe9vuwrfmw714Y3
Wd5AucKxvcTkE5385qikL0/zTwhSMcncU/0654SIXS5WHSmHnztsGs6lYfZXeME+
Di5hki4tpq/f0DcouTMI1+G0wy+x9AfEZqiZwcLZQgLcb+gNwCEtlal4s3Ss2y/X
O7vt/Y7qgR4ILboky8icMoON2NpkdXMeihv+BobHHG4UpFcGvgJijqfDLmMrFSJg
t18edcUnvM5pYaF5vRi79554csHCnPNg2DvuyLkNDh/fasA9D6EfRqRfmYYBMevZ
ffXqWWj1G/uh6gnMAdz6Zt7NtDxMi+sIseZB7njCNEuQepyAyD7d1RGlgNml1JbR
p0QWE/zV+90U3UGQlc0xWNhcKuopRuLe8ibtbNUnKak=
`protect END_PROTECTED
