`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zeC4bJzwsDJQbanNrXkme24+DFeneNEXh5VHN0McNTCgNiYqWOMLpw+c5ZUFuxsj
E0iR5RKsUwIxhmCE/XrOsG0vAdZW5yulf8eNHnD2h3hFf2NFMrs/6NOrIawoZAhE
ICl7UZZcmcH5oo/w7waHgbubIMXDkkDJRlEPpur/NtEXYenBypFrKHYV9FKQ9SLK
9vTRF2b2QLMshYg3c+jxeRdVpm7AhRWIqRZDrKFUQag59s3bVH/IhaS86v8FORff
2vb5K/cDGzzAdC4g8zB3f5pPKr/x99KR/3tNqqBR7UB5qoDi2y2JOAlHZmgTSp53
RnkfLRAMhCicD07pi9z04Mnd6gFGVVQ2KlRaqEE8tvL7hgCEFOgyU9WflcrHqFEZ
HlYQqxigPaorkyOai5BuEq6fjMKzdBftFreTIrOk3w4=
`protect END_PROTECTED
