`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jiumWmhvP4abTXROxGpHS4IbJzRKyjCsrotm3aL4d5z3HnbLfJenKOQzxFUCD+5C
RxAGl15y3nyV2LoBc68KmwvQn18VcIwaHKmmVHBs1QKGraZW7tyb9EtU243I1jQX
K7enE8AEGC6+7F0ARABaGMvRj/wE/zmJce4nDuJu6fZ5aXlynOtcnz1Ucp3y7njJ
FSovp7M8cnSgKrY53Z/8RGhME+SYTwybX2vz8s9v6IRxqXvOVSfjz6MMMjMOx9Wd
/RGMlST7RSuUVZSGMOavqyLdWdAz8B5LVxmElxv+lyGSq0vaXlAVGRQDtg7793sN
Tdka+i7/62otLtlL2qOpAveJgCbLac9oVuJc6DtJzEj23GL64t0+WCTlyGnsrZS/
JgRG0YzBLtN5HlcpYke9MKR+etCEqJjQd87UwQXfUNKTfZojFlsDDb0+HhhAy5sN
0pCRr7HngS+BwbufWaJK8yV/0+MrvLQS/lMH9THyufAaAXUhPcq+aLHGQFRcgrP3
SoaIi6wFwQv1iB3Iafen+FjQVLqdoHIylSOBjBXZmTAHyl36frVwg22kUIPd/sgS
Kpm8Mwro/x1xQDDARUgPGeeUqL+khNYaaFio3uA/GA/fZgPs0wLywqB3O2RxPEMa
Lhds3wG3lCMHXKRVd036+cUe6dc7FqYoFycYV9p6z5/e8EaVq9aX8nVVGRb8TztT
T1CVVh676CRlwXCLslqjH3WMiAtjsvklTyYEDtTQlWqXyB0Vu357E13gZgnzfVEI
muR/6CV1cjC3F015OM7zTyxoUaCagxQTwU5FngHFLzR2mbMvtp5stDXDcDCt5tnW
ajnkZpeXixEBzPAOaXeReSEGIqxgj4wGmMJw0EIuITuJy2Iaaf+plM0EugQytZ24
HO9Jb2OYZD1WtzIc5uS8iiZAV9u1enFIUxaF40lGeYBxxsOOL7bqmBAOMGyZrzsd
WrU1Qt44vVX6Qd/vJCoHG6RPqqfa82qWnlR/xay+5aTE965AQa/P9lTnfXxBmHA+
JRh6Basz5h9PneyB5wzdyKRXkzhdFeTYmOFl4zU4N6P5enHiqzJXFgvGYRfYzujR
6BJCDTS+OnP2ChBih5UwuUDoryaQKUjD1K/2ppc6b2fwQELJyWYG1WSWXzGHdiA4
OgnFBXXuL0WurFKhszh0tI9RMhFGvOux1jSh4U/k69/WYuJJVIiaN26R+6y2E3hU
7q49sSJb41BK68Dj8CoryOS6GbFmaVTMZHCjChnhajobKMabyS1xU6o6q4+USI/x
C7lTvZVgb47XgLG2XvIiTl15exM3/Fbu3t/sZUZOfaMvq4dyPUqzRFl6D23gk9gu
Hi2Be74+hLJTix3KQOwuRWyVOXJ9cJjQkUZQIlF28ABurxTf1A6nel/C25EU7Y1I
eUmOT5u1Y0WFS4AQoxTCWbzfYMNnfA4oh3Vm02+jOpB09kDR53rrogB52zuzrAAY
5R5n6NNQV/XYWBL19/xn12XBQX1qcoDVUPB1HCJBdW89GpVPSjHKJzsm/QZ1dFC5
P4b3HhITh99rTm3YeLwXPg8L/K07THm+1O7Iz0bwu4RpIr4P1NAIDu6D47IGocay
5Ts8D0DEoB0rM6dZqt3UFlHqfvoEDvPJW2rI/0SFGIw78B6a8y6nmYD2ru7lci4s
zj22Sr1AfIybLonLA4vy3+n+TQ8WNNdZb55sDBosple1iwRcPjTYvUTjTO+x4cYM
+PCs02Yt9B6Ys7GhaAQlbod4uh0TKO/ahoxPuTvSPhVb89TYwMKGORPbFvs0Kwkx
DuvurOnNDqugcwFIoAD5uJgMVAb+mWbVNaMGi7xaCAkx6LU9AEOFo3QW0jlnb9oU
+b/Qkkb1hz0Wpy0rKLQ1Cl+BBA94cstNHa4lLmQ3qpqKPLxj0pyhdAgMLgCWyc8s
tnP5fnsntXwxQsSEm+eY1aHwUwPQtQNQ30725GY5DKpA/UR0Tv/b0i+zlhKE5Pbk
vdw97QCm4wE36cNBPiHUiQdkcQNVsv0XIaJxTEscG1VzjjExmuQyHab/bNZifJab
kasLNXZTJ5L2hGuG06P9w4l+U4Ik2I++i8kJII8T6TVJrYXpSmB/YyMJPOeUOQnt
8L3FvrokAFC5KiLnXRnwZyrXB15LQTA5DKSLIIOkU8cO4PH/TNpa8L6huPh1bB07
VG7sq0F3wcR/20hHRkvBh3pUcPjsaPsUxqkaTA0WjL73aOv3HWlA4uLettKr3ZDC
1wcr7CjpUuPGNv3DgrD78Ptts1OAikmrkVqNjKQ8Rxai9NS2eCtIrdq5knvOmNQU
YIKF4wjZlsR7cZE3xtnxu9WxK+QxPd4B8kTH2JlzOdesb/ekVF6L9bW3iuVmqHfW
mh3qeI8c3AlZamDbK0Jp/82b3UjgudIarITvZh5/gDaizYHotdCIrFGmPJewfF20
VrWb7IEPHipNxbZXLFgb9x0oBhbkJjdCwlgzX4C1ozvqLwAjRo8aJ4pDkI3CYEar
ZRAIjt/cNNMRL9aQ6ZtFpDk8KRQgopbmz0YDVxIPN1NEop398dATw+10Oeq4rRn4
4jLgH3Jc8WblLd8lVWzIZ5pUsyce5feKReAmGuocRgFOETCEruMj0yU/TtuINRDA
hEwOGA/walSJ19NRHXAElt5t8SGz3EoxyRx5GqfdxiFVA+AieJ28ncGsbkeSg9J0
Ic3FUKwqzgkegZs5Q9c3IcMLxczvRom6FfBmaLAYtzij5szRPxAsM6iWlNgPQCMh
adkwqTSNBMFvVbqgfYrynkYvBEh23BPsd8R05AbC+3mY0prGcCE/r7tlpwbxVnSd
Ogd4Wh1Fdm1qy+3hoAMFKaV81c3GeKdRfx2T8O+iCVBGD7ePSTbY6knnUWm6Fgtj
Wg3S5f4kEdA0Kn/1dL6pvTSwroNGT218NqM0frb7yukF4eMPdEtFQTYBkoKtnLJQ
SdnJFFgHqJzUm8xhqJKfzdNuQgMxp3B/IzCvvVlZ0Ec0+VfIX9PIyiAl23CWOV6b
pZ5j/zvcSDvcII8lQQ9CPY/OYl3D2aDpT17piNINDnQCqrJ5ImbGjHImgqsq98Kj
t9/O0WzGrhS1VGWBx9SB8RJ1NUjnxqNYqXsiFhLxOE/6k8KE8PdrXjIhd/vIzdwG
El7utm6JvDZMCztSQQXZXq/PjTpipZrZWQRl1dnrbqeIQ8srJtQDWgD+1XyjecB0
b+mEwUNjYmuDA4WgUpBZ5EIDCkF4IfmdSXrW80LMNfPexswF/Irm7gSwr/iMGRvi
NjJs/uqMMbfSvjrr5jJzboI4XAGz+d0/3PhK7kDcBBUNHbN7uKaqG1HVKRldLM0I
LNt8yea7xXR0tvY1TzjviKTG5jKx84mMQ6aaWkX+8W1KLznrzLXw+aCfaAhlrDxg
rlhDsYYmxSPt7sLGIkr1qRz9XuQnDvS+MZsokYJmrXLLq3lQsl4yx0aTy8ojb1Ln
/l6WZX7uDkCFmor+DKLooTY6+HZlSkoT8yCc0lrAQ/ZyoddAVdOFyTGwXSyw7C3S
kiSOtWo159Z0d85f0FANLPGunYiEzV5g/GU1iA0+mN6mHHGDQ4Jx99+B8x/CHwJh
c8TA+C4haLZ10cEXZ5DrFYppA3agGclxU283s9xpA5S/3TirOwrlUuEWPa+p+F+O
04XVPeCXgy3EfqprAy0WMJLGzPt/6oP630rHWGyDlOQUWypDX/px+z/NDnxSgTe2
63r9hANA06V3nilrAkv7JsOmgmdeFN4qUIeTRQQ7Huaooy6/S4kVDaQSe5s7vYN2
4i+ZJQy4uufjewmoovzE/WpLxe8kV5els5sGhcWb2/oD2PdG2v83qdEquxVuKxOm
0d/Xr3ky2/NChB7EoV5zmaNIYSUu6oOkoSKRdlAqydIxShf+Uc4zuMkT0l5WCOVW
Yqlojs9d48SN5cugkl5IWH39OGgtL7/OHfC8XbyeHDyMVsL+F8nhx6NYjbZqABiA
jI4K9pyNcc6nOEb3fWrXTfbMo/mCl0t9pGCylt6jIr5jNDdQsVd5v/MgW7ijatxZ
FRByY4OdehfGAeF9zKamWclrQ5Vsfftmlh02mcq+r+hg6dVhtTlOBmZHFpFPTMTz
O/9IkrI99M0Em+rOZL31GM8iPjJtOd4GwILZsO/YSI6AnspC6xC2mXi7dsY81Pjm
Z/bbX1fFhIq8TkGFbHxr6QDz6W96jb3vhULSxH681a2PNftgjWPMo/DNemv2wvFZ
xuwxb2AcqmOLy8jG7El1vsgqGas+uzUWwKyszYCI1Dk9DwX3dzLmfTjAySjcWJDc
gsdzSCrCciFHPbsXqi1OwJ6h0gn3HZwhzlvrOS5ErsNr1ofV6EVjB4CxNhDdRhG6
SibWt38KobKeLgZP7m+i5YNyAupl7+9y5fd2YrHXlbt02Um9WOGp3bLfHzYFyN1Q
ZueeFO1DI0HX4z6OA3qDzCflR53/314A2dWhQY6heKyT2a1wCdhUe43Lu0HQphfb
l5DIMM7AmRiAyxZBHIlkqHb2LJ+un3o2ErxENXT/qyfPNZV1qtqZJqOItqpZ370n
0pe+AXLuPw2HW4YzQIyWxW1UBymu2qSwUlaHUAYIeO2SBzUU0h6+IZbDq2OCC7XG
J5mIByZmtw/7NdF7+RBtsKE99DvxqJfPgArRydEyIIUIIBoyvtG+szga+sh3PRoU
YdyEq/+PxNE5Yj/0kg8lywJuBOXX76i+S0oihMi5e3avLjfhkarIskL+G7MQSbQS
WI4PPr4/mZomTNDgXmCDBw8kSpqbi0KV4dANecfgxF5CC7MFY2y4ypcYpTGapOr3
zEQ2xitR/CsgqKTFne4r6sTbbA8+pR5IK/L4C0NkYEMUtHjbqbjNYanm+PcREJhI
XDmQe4ZvXuHjgOWbZ6WvoXHJkHf3FbTaN8dSa2iLq2w5O9sqrWNtMrK98N+Fx+PH
HLuAM2FL2yDUXIjv9PbGAePwsm1+joaB+aAm2QE2oZBt3ODW3gb+Eu7HnHvzBR4H
UO+v0sDYzQoaPBCwQjKk+sp/Nj/DWn4GAi0KYweXq0xgDBU2SaiqccucXHP1F3bG
iYxa9nL1zwtOsNDTLq8Gad4tr9o6pvKA90p1Q4DzUT1/IUmD3dLnQ/rJOyxWoo5f
2jqwQpED6kEBK0ujdA4Di1Wo4/QzZXGb1eGQM/llqy2rRPJ/lFaweE558p1fiX6E
NF+Wl0xkKfXncTLJqOdOPcxK5IVYnskUjI/t54L+T34LW2YjvTfLwTLcQVpRVQRG
I81Eh5AzLUhFCKOvJNTI4J+3bvpPa+s4Z9NQgAlCJ9aWPMJoX2Cdx3VxXyAH/5sg
+CV8sSkgx9Bvx8VEM2Q8br89fp5+m/LIgqSAYDAzbGHERrAiAA18/3HblHXFyDuI
SSUcD/TaHaAfvqP921jVyKCz08MyYxygRaltDTOZJ2DvFVvBKu+v0dRtDlSGpCys
Ffn9NhbOERljbwXwB9lzvTcy2X9jcoBbgTI55d+yX8XcrcQkBwPRnK5DsykHYRC/
TTooxGGqTfa1P2/cNS9J/eoyyMBynwnqMgmg69Tc/CCT3HM9anhc/GOkIDvDBjZd
d51kl23gmMiLf3DDtm2LRw+YHRn8fA8tQDqR/E/Ppk+ZoHf4zjpr2bgOX/WW7wrD
4aWDxr0ZGlKmQSPJDB+LaY7qJSh1MwfRq/Hd4CPdcB3FIlT6dDmUtdpkbP8Y+z/y
W3lLKSZdwZKTr2Lm/VY11PWJbiLaB3VQb98QtmOeyjFiszWrPTRXyXzQovK15qDn
zJt98GTS+FORHPPFpg+n825DqKSKHZot96VXViwk5eqzmqpLcM9Oec+YyJBI6/0z
DTiwgIb+qAQrj/jj3BWlzNI1f2RIO4lA+9Qeb8befogutZFkhPsUkihx7qWzSqxh
2+l9nG+yLoeVZG7DwUF17ENgu++XekpLLWlgRTQMtUeFQY8aiHhoPy6HVrYmlxO0
ODLRccFddCIHfRaZ4ujJpL5j2VsYE/Qrn44PlL3Wso5C7X2kQsbKaBySr/K/EuI3
wFc5zf8dvlniF+2rdVcDbBbgmogaaD/DTtyuwo+4LPA6vzG7MCblBqEo1TSGX2PQ
kUJWEeiu4kXzMsyAmmdFb9WwSvrb+OfO0/nRYSdZe77QRgQfBSM3R8yKOD6bnNuR
EiiBEvXwdacjUgA7GmFXniMn7EfVZFwPJGuSuxAzxKJ+xPnYP1lhKaYWO6cfVxaS
McMdumgnHpY8KT0R5g0+S5jb+7iQG0GT1iNHKnd04pxGos4TUi65fGOlpF5N9W5z
irftCNunxov+RzlbZBWwt3J1GgHJgXPZp9VElFKsxbfKBDniGgUE6YeIFJcC94TM
O7XLM8KZJAPgkRY1O6QdrCP9M51nmjbTXvRM4AUx1wxuDgqPCW2255S0dzZ/7t+B
wkERJKKATFx5WRqTd1WWCum3kykxl5R1xMV3X1GoMt4PQGeXI+VObIJtrpLXtkiY
H8+QvLDkuJqHXQX/fLmn0CIb38HI2A2TmYdMSXy76+W3OkqWZTuBxBkZBA7xBimz
TlBoKTsJNTGWQsmjUK6pBvtCs3sZI5J7Ybclsxnk6bOlqoM/qxILUAH0eJEHhM/h
eCdC2qDJW/FD+/TPBbIcMXLwI1tyCHDDy9JItgs/GMNlcFTzly8KAXIxtTb2+QGg
7sx8LKPe7UPh5NItixm783D1886g/HfM3Gv3SMxc0zxYsgrdDnQdFQ1n5zc18ROl
j0wzcPfysZJCdkLw+uraZXRdpVRBFzMdPEP7fv+1M3jEAmNUEeT3pNRMmn3SRLAk
hoev2XK0eersjglBahxY9LhEWZjjeY34YCMyNHvAajoL2YXIaqjmhj3il1JWbB8Q
s93eBzt1NWdakOzTIw9SP1YJ9kJAh+aGGnqo2Oy0YwtA3wrmBCrbKkaMTpAGmzgx
gXWZU3tzZd1/TPSR50N+byj+CWKmzgaznMyYlW2Jhha5iOZg8B8wSQndRo2CG7+d
Y2a2sW2thm6SWb6XHOpkePZ7IN3JQbo5FxIwc7HqGceZvtN1ZobfTLcArdrLBrWo
+aiXPIiLx07lVw9d4Hx5/Z1T6QL3q+GjL1PlmZyFuYyYJ0QbdtOhfdDRbhPIORmv
R/kSNhFbMxsh2J0vi8kfmtnc5qxNjWq+7EY8kthMKpqPd/9kYEiMF6CM8vS0uI5W
EaPHgvmY2OD241t9Y9JCMeMuP3dvvwcAOdOvq0yyzOWCBcJa4s/EWBQYaj+lRYNe
QhAFaz/41Kyr7p0DCteiA4asv4P1hFHahBoq5ApC9DPdRhwacR20Y6p5Xinb136k
05BFRN2ormN9IriQ4YsuoKgexgKQJeUh8p29XUmsHkHuUdixoehHi/0yqau/2xIp
cPbUFcV67mavCRDMGuawF7M2hjcnaeAW+hyreP/cHhwqdPvy6NQwLtgwIw+kifAz
igVdomEbDH5C/Sw42XQDoI1bhcF7qh0BhlU/qx35zxew25CDAZylqbEfqTyf4ROp
D7Xz4cAMzsY/xCLbWgZfOITSzRfquQhzj4SAX4SL22wyvWya7+fvyDyukMqS5iwn
qKuuy5Gz0G5HkAlqZZXwlQ8v8CWBjLSUtFJtHViwEneHi7QiEXFvKx8k9j03uBvi
CuIoT+FIUaY+eRwU67uIzCi4gD8RPdovKQHwNg0opVYEhQ/BFRkDqsoGODi8jQCJ
UVmmqNAO93vfyCY7E48PDg3f1sihyj1gvd0GucEJkM5OFb6w7BTTUjzFDejXElbD
CScTsxl6d3KsbCEY+/WuVsd9BBYOsqD3BNzjQTSC3Vx8hf9LeHjXXpoKguv1ms9Y
n8yTxbUUWaWjGepWUhtMl2rqK4N7A51zQJ7XC/ENIEJl4rH4beeIIK7xCZbd23Eq
IinGGuwPn/kIIWiWapxkUICKNO8ayI6JPis6AzckzfMY34V5er3ldOdS0D2sizQc
TbI3pPGrY/ChGvOTZ7cEXS4ZNhkpjxdIUA5peopyjNPAQwLs+TDZJTJm/KcMO8lN
hv043Ax5MyEXB1uCZ5wDaGf5OxNEBBZd2HBbeTecVIgHGjIoIg6+MwLzywHRU2AR
JBoQ/r8NGgYYyNhPbBiNkt/fjUzF1Tw2MC1zu9NaIc4ZlwdKX3K0CUcM0KOlJPtC
ct+b3dSLruFeXXQ7juTernPjtvIsBSrNxYTQoXYlk/4WzWj+98c7obETcwAUaTJw
lGNf/o8vGtvb/sEBVpSkljjVNi0mlBlfNP8/G83FeQQvp0YZ6+3cj160Dl93IsJV
jCAb/3Sz3ThJW+cwHh+NHuyY1TYdRD+PjXqaOB0rQotfkDwMCl3Rgb9YgMu9KjJc
hyHsZw/Oluz9A6TcV+PtMGsqiTS32kKP9dNOrE1WBOnd/OhUPhGZ5uWaJWekFsxE
h3pZzV4MrCpxpzNpZu7AenG/ib0LHuLD7mNFthNX2WKYzyYMTgL/s4nbZgMcvLUB
fzShF2/ilcTgMS0tEtfnVJBHeKhKGSJRBdX0qA00v5LPOfo3S0eUmcSHJF/lt7re
P8w+mI0XsKS0A030VSvmchBQkRSwvvFzjgYrd5ah8pWvMCrSyGltUPrJLSuZYc9j
+7ypIrHzd7Zzc5yal+eyeItA+PGuu97Vk+vF4CxgVWvkA2jx7NpBpbgimqHr1eSr
0lZCstrBrX3W9G/4f/3/sMr9Aq4aPAOgnSjjUAIzKaRCBApPwqVeN7c/dLUzZ7Cw
1Xvb1Er8HS4C3GWhsQblUEiJAr3rjXpKrHGGvmb4JawmvqWNqleRm0zHMKBCofts
4JStnBmtN4ZTm9JkBfZxy/fRt18V4W3uWCtG7CjLibhoeXX5OmXE/niNjLOMuykC
HAhkU5eJ5ghETt7t4P6AgSV5E2+MVlnLEkllwVz7X8FqONe3PQIZm0aWkZvhlkDj
21dwW7cCNyWlmKwukaJkVf4KoEpJuVs0O1bCAK9vIhyo1PCMzlC5B5suyv3sciRy
xXD8jzoHadOi8M3NxtR1NEEFnjcGYtibjkciSWlf2wJltf+ved2bPSZnpTSjjYAj
qKncE7THoQ7c6CUiAYRO1sCsGU4GXIUqfcm00QnjWkxW+DE+5n5xe/gJoscW5d0l
uHis3YtUVCpfAAHEJKnUNjDjoAK6DnlfYNxFRGOphROYkedoHZfr4H/QkI/QMQhq
w4EDHNK0rwT3yZ0UYRAcvO+j0o/t+rFv7AWJIlYYEsbK3+tlw79CNwxbsJWJz9RY
0I5FtrXe/Wlyd1Rs26kv8J0JJ7qUX2/dTX0XxL32Q6s94HXz0WPlG+aE5GA8jU6W
uZY0gWaGIckIm9JnCJcsDYcuUChkaeUehsxjg4gQ+30HgPqe38F0vN3p+ttj2WRy
i+JjY/75WfEEVojuIQbD5N86q53ZU4ZROqe3tAV/Jox9gyL4LQv73nsHawA9ONuD
xOFIZcLyZsPiCKJfkDKsUaScri1RX80Ercmh/FsT253l/JgnawOnsJau961G2nTY
osrwHzX702zG0Cs7kLp+dJp7mLtjnEXiw/6bsRGimE+048NNKjUCQhLcGxWmq6rx
2qKGzow8ND3IhLZdUsSpdwXaL+12K4EMQ4fgGkd8EjutLtHNDe0WeU1dq7VJSCn7
YsuSsW3nEHU9+Bc+bqGqBeDwobk1KQ3VP5/jW3Ga7j8+tVHFlmHsM/IMJDQK63Cv
qB5Jm0p2wCrOo8h0oVVrPVPqN9DU70RZ5/R9EK6dYgyAn/BRPU0uy98jhqGJjJz+
sDWfyBzXI/ZX4Iwl6ozF0gTTLbnpb54DzGwXYg1IDRGCCEH+Ue9auWT9t04j60s5
erIW3qbTetrbNhKRRh7WQ6UfVUpOCGzTePuxutcrg85wCXC9R0oG2ZxIwVo4FIad
I9Ewrb/9mob2LFp+oJS+3MNVdkfUvYRQX05Q4IVCtcmqi3aUfflj+gSR18PeYPq0
CU/ZA8ejtUvmyNpqEIFGZEuIz/qG3voXXYxIEN8LVUg27YTS+Ig8W6kXwzO3tM4b
BcnVqOd/aroieLDN5p/6/Z22umbV80uJcuHPw8SwXQf6+OWqipM9aiRF9qgklxjQ
BxnHW3XVyhJimGXkK9qxgoQnlx5LgBgivgWTZdJNEoML/AdoJLMt+qLJsY1YC2r/
uuTL8w9ajbowD+RGaD5qPsZv4y6OwoC01H4JsTZhb5G+V0OoDT9iSvACCoODjoCX
7zlCu8seRI8cL4KSFShUc2KxvNZiY+bcXT3z6mhdXPUVv3qsnzSWGlq8tfLXZWen
JBj1+iOWgT2Eki9dE8lUXs94DQxZ7XWSd7GZWrwAqE9ATsWxbhptTLJse6+cHlDM
a0FvsvzgVQJLyWaceSLgj8be5dMmoUeKU2meAaJFvmBrPs98fH3TVWkFLrFMc92R
SB948I6lqenHpaMGSjwjjgfAUmCXQAYwiuUFammw7ggNGioI+BRkPCHNXO18xI8r
8f/ezXvlL23dCn7vHrHUDjoU99ZXVwuahXq+r9Sdak/3txCfT3ge4D4UwOXkVxn+
t1xKeTWU9HrVjdv8nVPykH4Yh/A/hyXOME8rE5rVdDP/dEQnHfxuCM0KPTdzdrgT
onJJzt/423xqCfuLYseXX+VYawqBfB8a7cXsv/cPDYbAWNNByvYK3Bkj3JvNzvhw
7u/rQpLbEdocFkcHhwksHzNdQypayukQYnF0Dd1SfMneK9+Lmep1jD0UFxU7Zyy1
B17KmaXaE8ZGscm0GmUhun9EuGBled9qiRLJaZ7kxx7uof3hBG3S+JnUrrQD1B62
724AHPrNl9KPWIjiAWcgje4eBrzBsm/62iKKVOY6V6nj3qEFk1B5GKBpvaqinPCp
K7kk+34jEHDRu7HjY2l3V8o1av2+TZWfgtJiITJEpcDOzj4CfsgRo9ucO+LAwQdd
uSxVrhmor0R7YX+DxtBfY+a6gBD6AhIsJ4P5bslFSrZ21E33UxKPluzYzjrkh+/E
gEfdRBG39g1n6tpx/Jh9HGMDd6iz0ZiZReqj6br2N6GjEkuPhyQDYmjxUKqrFgNO
KkPfqOJDK5Z3hDdXQ9P1n0NG/MtQqWBvLttNLjWuRYggOj64/ftT+1GVwA6GQl0Q
G42+VETOCXDJ2gYtH2KerN813RVFehPE6lvvnSHLzzUWtINnuS2cGylMId2Zrn0E
pN6Eyo42hSIGFKLl6wMbV3ZuDouVj2Xcyted/DEB/esZXx9Sr+4DFSX5r35Eu2nZ
9myJW6PDGgioFz52d8jDdgeWolwnpwQAjOPpDTwJiVPcHQR07QybAMwaT5XOJ90J
o0FDmyoua9PBYh/OTz3wRN3bfnMeC51GIXAl0sXc9onzoVk8KBbWGGluSq2LPKPN
9/nix3KAvdoj+yS+ViYAM0e1liNI+OqDTdQWzM1P62c3+Ct0rjWd6QJow3hpxo3y
dLq85EJknoPyf1Gu0rkzHyA58bGqtnEuPCjUUf/jqvhXAq6g8e1rQccdbuaN2vZj
trbshbAq/U8BoXoAdrjqpMO5DIAklGhBIrGHIdnyJWYTzrWtw1CBPykqUMJxZHbH
PSa1sRWFww9bB+yGVBBDtq3OwQGSh/3bgq0UVKHiDEhilJbddEwNUo4oWWmFOXCC
kehGo1YPXhTnDxR9t1KXz2WPx9Pzhv+la/25zGXwGzbW8D7pIdoqhkHryRYlT3gt
UOF8NhqK0kE6QV14Zmx0cYkgpgqPW/X7mIkxC+vNFR0EslRyqBgKK3RJk4kMQvYl
CDtHQWL+HPIBKHfUsNJOIatKxDVAfu7LrXqyXE2KvZYd873OMOQQlnGeXvrFuVE+
+AeCpHrzv2tzuAD2OEYtK/i8+DniI7LTHySrjQ65rUaV6c06jugtB5Mq/JBfeJ5x
td5zrGgH0066c8DZxLeHMdl/BneqoMb9/AevFQD+9OiQD5u2oLLElFaflJAsRHY8
/UVnRm9Q/uy45nc6rmzZ9DbRxyfa9/0geMHGTwmzvUta2DILToSzRGjmilrkUyOg
FBA7pS9oNbf1/qlk3yWNBINBYKSceF9/8QkhrzT0N1Bc/eEl+ZUJKvL2i4LJgaf8
XhnCK0yLLiCNtGADOy170HrSo0CBuSh2YPhCTSLoFvNhhEmdh9N67t8M3acrQdAO
039ydJt+h5kk2khbxPf3zGUoYJwIElitnuWN8nfgVJW3OERpN4FIA7atYEDWc9cn
631jmZctpdMi2vsiMbR3+HX96xLVRcrj7K85zx+ysY7IXoys2Yx9C+0VuiG+75in
hdBYBulAy+WayICDm0S46m990XNb7RvAiXaB+h9qe32Hs6hbRjLb1KzZppNDUFuR
eLJmv36mwYXI0jK3t8hgs5geeG/FQl/DKiFetW0RGf8bIBM6xnPfgSI3VhzMpw7R
1CSapcRvYo0bdVoGcuuiqIl2gsVih46o8wDlR5Rq3m69I+9GTSxJr+vsyZjPQDCd
stHFEHDHXXXJEcdW4douuHovgONCfCjGCmU1s8HAwZribWP/0iQ3wluNMzixT9sX
MAjOAuikO92I0ovs9SmYRl1LqUOc6vng4J3632D34GDKRv04/lgX3oJQ4rhJXZAS
Wtft7wfuujv3KBNexr5zu7ZCvzVXaNxb7DRUKhaeXPZLyWye+425cIbMEzUlR49o
kE2YJWBhW73uMbcAV1KPn9DxAkfRuO6bSlzC6l07ZJix0noeFIwqDawaHMeq/HLq
LSeZz1ZrVvw+npSo9sbaPp9qz+E+oPsk1mWwZwaabGpB7s/AJsioBYqQNFhnTYkC
mo8p6xE+Qh+t044Ogl06T5oKS7JcI9V0V+1vyfyNLoq7kwIG0AjhWlucyKyF3T4m
n240DXg62i8HqO4a9Oz1DGtng0GJh3heND/raonPnWY3eRlUY3+c4us7n749Ls7N
/UFxjheRE9NC6DmLFtSquMY9JL1TS+WW5GYL95h/Tc32xyEN8T8Q5lmVhA46SKVc
kIbHRG9QyZVpIikp5Dgxt60RrmEUIKUTpAFDISTX8WEEPzWm1jDeYNrEe/3l4C8l
tjf5UCm1Fcin0g3GzExEX8WtpvYhq+fRTPcdoLE23A9J/QEGP50frbsoWtpsENpD
POVsGf+5kNULJROA3ueVR1RJfyeiUsbNby8PKMrdlTmmxFQNN9nTUTnZmiRPCHbQ
noYTW2fb1JGfLtFau31MbSCKnkbUroRT3ZcxGHj6SnFz7RdsfvuP3E7svB9hSjvd
CAJFBBRiTUl+ykMCPyM5B6SgR7qB9BgM/aKPhjeL4oRNuwbEG60xK50bU/WrpncR
fZOnzZklcTsDWKCxOk59ILEEw7tGjwfKv6k1NjAWkKHrebD5qaTqa4qTlqlw5gcm
idKLoLzeXNywfZBV1+/XqHV/TLd6mcXRaSCdx6+9sLlLcZs1kqdUnR9r0YhrSIcG
RHIYPHuQwz0HmnFg0sq30MA5smADCbk9KVm6fSSwX0eb8iHcZIpx4g/YIVnlENRs
rYutVdAV9gdvCEuSTwWWzdEzT3Pa9mePJfylemolI+/I8uHo6tv8oaTgakaXmw/n
gHMTEJssxe8avOIYbWNZUKMxC5x1FKreiNeDVaDZe2qEvyKdFPe+Ipur4E0E9977
qTPFARxCbhHhAHC/kq8RhYsNxQa9safX4Ce36yHHO2Z12ya2iUDmGX7xkb3AfCiX
YOYM7lMpsFNBSbi8MiLTq6BhiYt5zVFD0c9SMRObGaE8Rs6X4k3LYINkwtows4i8
XKTYjxM6w0G4vhrXCv3WpcA/vl/l7BoRuSvxoRWPvfz/4RDdDGna8U965qL8aveK
JebJM+5abqgQl2JEyqS8akD/1wVcLUdNTT5IH7fqD+4h1/P5aavBrpbjCzMI3iRp
22FEdtl1LWXZ6mpyM8OJb2CchwAU/qP8rFYHhrgMx8/awpBSRrNxgMr2TgkQkSRI
eVbfo5rbW7T1kieSykXLQrpyS7PTcZMUL57Hr5p47czdH7klPXCWot501uMQ6wKf
nS3V6HTMa1h9uv7ELj4CEGaEtKNsCU1fzi+yjU4nV+vMOPG/ikNL2xiuvXD4+NBx
eef1/Qr5YKQ1DQCoDqFW2W9SHeAZwDmOHyL51r8IaqMqgpaJK82TdrsXjKdKA+U0
dbqhwDxHe4M8SjNSyJrup1HLyevNwBuLWxB6zVe5cRETjIAfEU8mIz5BXuoKc2FX
SSQAL3EcLMqOA8/qAUOn7QKWORgRyQ3763QmbnfZfpZZ+INEf57xKu5SFGW9feKG
`protect END_PROTECTED
