`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qOE7cIDOznsBFQhkn4DHEg4NT8KROXOTyvtpOJ+qa84maS0p5Qdco8J0Tq2KXef0
lkPWX7o+oVzWAjX19XpPZfC8E0MiuNs0HT9kt30o0uzgm2wNqi4RNjzCnC5W+/B3
bkHuHHWRkdlGHTzsPJmEIzw1Db1axp2E5+D/ZLRaR4oruQljZA2Mscy0clOt0KOC
lMSfoSIog/xs3gR2KitgvI94RH5PCVq9U4T8uomT58thbqoMpsurFeqKWHmEYd99
QPGiyG25Y4q5QAY7bBcb0Dmmtevjd/2UW74/Ss9M+2L8AnSni40x0r02t8xH02yW
G5Ie6ccgKm4qBobZopNp7CKbjYJtsJnHi44Cqg3Ndee/nnf0YRCslqxiiuPyPEz0
nCg8DxPUyrwHB1LRi51iRr3W7YHlqk965H1Y2h+TZ9NRAsBREofhJIJOj+jNSO7y
9PMQm32/hkWk4uHbnXnOK8zD6PlD/Exwv9WrAVkAhyOTpcC20MEcyLZsm+qBPaNT
A+TdljiItUH6R9Bs8aeiSz/tVLA62T8ejimA1jlFvoDX7lyXBjn+I+kct2aaXODE
vqWNNM/Goo4srOPk/VBzFy91/v/T5hoeBIPgKZymDxpID5mXXST8EGaVs6OQL1CX
UobHsCX7KvdxlUw/0UQMhE3L9lRD9Bqq/xogfNtB6Og2vvbUrVxmHDrESKQWM/zS
cmPJU3cwMckJsdyeJI9nvHt7cTLcBnS6947lPW30h4eK3eYCihE23iL00ap3HH3P
SVWbpPaZL/9W82tFoiH7ARO7nqGf65EHCN+pWFlZtCyprtLEpmnUhDw9wTQcWBk4
de0Rb2lrwYNj2YgM+dCPt0fh0ZRd8lmmisAFaOXuNy6O0+ANzA9A96jyT0Ft97ig
JMTJIQwckCWncbVTJ0sTSBSwayAMo1O6lg7SkTRgB350acw/DQd81sm0/2KA5wQN
huXPvxpEi14KTWUrryefTdeOqz8ag5ea7xT4DNkUX9FfUXpE35TLlluoidePpMXE
3gbj7FXqxT3kf1ypGEILGhmcpN1EvdpYMDVTRr9VK/yVeYhcPybCVRyOQl3dv6W1
VYvkq7834xj1E6UTx4bcMA+80HB4bBIuGpI1LjR3xIbDr1THXkH7bm6CQ/0vGFaB
AQoNA7UW0YfaxcvCB72Lol5cIlMReQSWu54bI1c3gxcNGdvx/+D9gxZMRSzTb8OI
ZiLwfRgcfdBea5wNiTQsNJMZQ45zNpwAczS0oTAXOw0eKmH42X8KqM3/nHq3XXi2
dSSy/d4P8edIo6UqHKmJ7WPehbS/WWaQPP22/GH6MFePjf3IKE9tM7Bh9/lmfRdN
Eec7CUiPw49NzSQsCGVsVM5mH9JOG17TmspYpUEEJAzhR/MDGV3gP/OOZdOIdeXK
KhA46Bx2Vqp4zFxhfZanNnZk/yOlAcxEEWxN+g3dGMJ4HN7DhRvwPo/GB/esgaVU
Bbnx8gfyT8Xti5u9Vbbzfe8botdD6r9h8Aalz6UBSSfErer58d3K9KPgHakllki1
`protect END_PROTECTED
