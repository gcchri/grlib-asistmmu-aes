`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QpvUIMcsC5yMy60kkNHI+hyAjBamhuBtYOwN4lSS9eAYkZ9C4AFjqI6/CLROVEyv
WMlB+Iq8CIoHQHlQIpXpDMOXYLWqsOil7xZGiO3cG7SErcVxKKwlE+QzLe74R4m8
aXp4n1E2HEIlnPMxlyr2CscvlUkkOSxO5+y5mtRulReThL5xoYKS30QuypjwMyZW
ct7osob3j2pfs+HE2QnBVtEA/GPNyxeC/b8tMUkg6UuKyjLCzpCTl/CIFDPKUzsJ
NMYr1lH6OlhBW7DVn9BCfMt5qisXMkq39KClvhYgsuTMxxlF8aC4PkhwEQN6d7zX
/Jpa3PJIDRoREi+TsK3xFy5NQ4ggtzLXS5ApnZ1UpA0CBu+iDdh36rgAu/njeo77
9pGdOhB+a+3Dc9ME6U8DvY5Zcg4KlLRuwi1GP73pxc9+8vXzLyi0VolwHEImVvXJ
ETxCL6yPrs1jlPUB7eK+GtECsehF3bT3Mgf8ScfYvxhhOxvmXIevTm0sZKLrCMzb
RzWFgSswt5vcLzKSvhKKSefZHtHLgn1VI4JV/8C59A3ecMRSklSP2YzBUdgVdJjp
oNOHVxcmXzHCF9k0QeRarZmMz6oBWB3ZjZwRyKGnr3mStPuYa1VilW7k36hNuZmO
nrJ8iZXchenOvtjRcEzmeyl2wcEfLLpMVMelI5NAeLovqvJ4UpSa3sceT6ekcB4F
w9RxE1onpcK1c+ff9PuZKT5/VUaWnKvBZYgeYBuNPVezjyzQ/o9OnMbc0DUMi8h7
2Mxj0YwImt3fM1yC/3OAqHUoR3XhwMMeH0Yvm25kOJC0xciKEyMqvF+67U5NfB8O
2Dfr1bFrX+FalgIby17Xe2mvLJ0KPVCAVIelUtPyU96BAdSWfP9+Pp/6TC3JIACl
qf+5qXwWBvnq3yOsefvU0VCpfrcW1+d9UnI/UNZptJKXMD4vkgWmM1uAwhkMcFUh
vW0hngDUi4le3azga7gmkfu+XumgGN2+sgO+wZ9/6to0jGr8gXebRcTBc9kXSDFm
JSmrSTJOTj0gc/oNdnT8CudWwyjEaa33lMq8X9Zf54ia+BDO6FChH5vsen9eRtQX
Lw+smJzJtvboGZDOyd3/lCcd7Q28MPEfRM5QLLTMXmrR0PGDep6E8inqH5Muhyu6
5hFEx+CNMe40GIKNegFnaffY9nDthlKDWcLDh+fMUJ7hq7d5ll7rax+7zyW64NSe
UJiF+Y1yy1QElTM0VYtXuIy+yNqnz15hlhK9glcO2iV/0FqtBk5P4G3p0MIWHrUb
`protect END_PROTECTED
