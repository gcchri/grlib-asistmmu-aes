`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wm9Y9JvjVcTkl2HPrPMN+kHZOH24ewEYZtTZ087KCMeBgtNm5IOJKG2lzv+UwgEq
/P3F+NiNagnssdd16cnr1CcywqYAvvDiNRC47xbcQROeuAWVLYuRGaO7edXE32sl
NRcvy043mJx/c7jJmzhsaORMpemFOww3Klk8JFLOddpVbW4v2FvdCG7AadZMuYyE
TjJ6f0bWNm9ZIHjvZYZFHU1Kp/lWJ7R7US90pMYO+l1QD/rSSnhatmaCmg00ZmqT
tTBLyB+RT8FLYCRp/UxPlQ+y8AuKqkYaZUm8W63rOfmE30wISq+n7Zs6LlVA2NGz
9XFezXvPVx53XeuXjfZJtE7aMCq3bxeL6I8JBmEZtZSkvsJUGIEhBQM3HMrn5asY
WdubVTk2eJtuLCaDxh3XBFCAysdKvBHZ+hnp+N7WnSnZmd1x8iIXkJgKrRXaf3Mn
LVRRGv5wiwhnInlAquM2TauvZXmozfjS+jgD/KLhAKCHEaKr1eBpZ0SybQdLzXBf
zL3emvFaibmNpuJJReX+1sdvnxrP0o0PxviWRPU+AJ/zVjBC/FZOqbBQvKlOUreS
3LL0MgrshLgzHhKGXyFZdYZUNxBRueEg3YFwSyy174qugOn2HR1yqjBT8UHBJaZF
AUxV5/TsbovDsiakgKxWrp3mHSIsRupsMCLd32/e1n6CXmgbwKJW8q8urQ7Sev9K
zibp+X3gba3Y6f4f2zk8jg==
`protect END_PROTECTED
