`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xovm8WW3PefT1+sUZfifUe02mJf87ekInk3t4qZDIy+pjGrC5S8j8jsH58DwMM/6
yleuWDESDQYK+nec1hHZsRF5nNWDltcyx64654nYoq5spO6HidJMX0Ah0hrsvJl2
1mUjy+cKu6YtYJHaUy6hNBAyWQ7UNsEwiSnVeuBzNUf1/ykgsw9hK4wx11rmO9jw
RKeCitwEnpV+cGtLYeV5N3TTqktTVeirk8SToF6QYM6zMqfJXSGhC8DApUn2HqjP
o3/nmlPSZISUBuaShnG/hjQA6gJlhF3dH2G1xZdbPsFxglybxqOP5QCTlt4eW6jV
zrKetz9K42fPXjSGYSkMHozLBXChdow6h6DFdpsNwjHAZrotlBInREehc6g2uW5o
7dxFwU2tNX7BNeDxQBFo6bf8XxJeGwPhtGznCt22DVe4Fyl71kns96Z1NmPo2VAK
8DEWRBcrF0nbve+H0K3LcqxUsLijpOKh2uGCoOY0yy25g1DWJSWpdgg1H3qrP03d
x6iDyg4KsLtMwGpKufBxZ9Wfz7lVt92oW4S28bBMoPISBRwHupqEg824MuxWbHvX
31pNZ+NcuJteSSwbsY3qdxhe6DUbsTN53d0Ue8WoW1I=
`protect END_PROTECTED
