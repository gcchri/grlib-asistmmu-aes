`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8eno708Mj2Cvcpo6geOrI9uot38zrushqNALmjTqVFQ4dRp2Gmvcta71XqQZMxdl
r8w4giTqt0YMQd7GixBNfk62MsN9plupPJ3+X+phJHv6oNy1V2JbCUBSz6oJ2VIk
EmrnqVIVANin3iSsLGdOiQF3MBuk/n7rkUiqLWBtmVApAJVG6Jj/L1kX1/jo0Sw7
gvC31vuIjEtTvxyJBNFOSP+YWBki/1RBnZcLLdG7bYHPbI2l7GRpheq5mIkRIk7U
eHIhEP5v3IQxHLottZLmqa4lJrnaIzVNjKhKLohX97VdHhTEIROsPyG9nK1i9xEu
EuKblmd11ngo5arrqqz/ByRUHzjj+Hc1dWW1qVFJTFdfEV2LgjRbIk/LKyFK3E6a
nWHeSTfakLGgJpCqHNYlY+QkaEtZHlqw2FGLysR2rTm9NEQom/38n4INFw4vLgrA
oSWwTKrcv9YA9EHSH8nsizCVZdZeRkJclMP4yTV4qN+yJBZSAPWF3aHTwp5FE1qO
9YawYLPE+XyjEF3x1ski0RVfNLyUqzX41CoNEiRswr2+rpkcVPzezPorr/Yg/uJr
nISLT2j/MsDO25NGUiWPfXND8PvR+TZghOPxQgqR5+FK0R4d5NTINFqpCImgf6rI
54+96YGZh084wEcKOpt/f4/WuU4BgnFJ3ChP77vrJ5Fkhk2GR8QyeI7C3JXcokbH
P1VCv9KQGMHckAL2nbFWgx3p6Sip15eHPnn/ALVMKy7JH4hCy5Stz6pGdZTPc7u5
cOKqyw0nZUz72eJsOvjvWf0WQp1RxRRcamvtbwpyRIuF62qJ0mE+zYTkb5YrA+DL
hs4Ufp8W/UGVJ2NSjx+gab1TgF6aM/wJi25g+d7NrjFZEdso9+73S/7hu823+eTF
yMu2mrbJBRJ5RlPnM0bpFYYdYvwAkr3/uvkqCvLvhm3X2mZ8hJfK6A4I1oPQXILY
Lt01sDxUKBQ6g7MI/uxZxPGHuq83HbLpC7SEbExuhpPSXE86bZdhFb69odbF7aVV
1J7MkVcy1s5yPOcdT2Asw95Sd7uLx5hWaffJrF9BZDQED4kSjWY2rAtU5AXBDLpe
ha9nqrLUaM4qJZWmy9HbvKXwqDwas0SAnSTo+4flSbEVNOjwHVC+aZzDKdltXxxQ
EO0uoZcWaRc/5BrdxeH04qqhQyvedUVZCc+JDevCG1AvoDvV16ezXWDKkzwIHY1b
iRv9ESsdJmMfYzJLdrJxk5lixhp1oJf2Q/u3tN0aRryHb4EVQyFmpjrYfHohdX2+
KzAU7Z4xQUuLgol85G8g/fQPeWqeH+9twGzHywPh4iecIVUKF4Ah1JElSUoPjv8P
vCizIckT38njVA7+sN3E++CNnsAuOh/2KgrqzYi1HUErS4dSh2X/GEeo/PDoMeIq
Ppe2cI0JvbJD3uhZkOmbwlD69T5IRUQuave0NrKB+VRF8ZmnKkzsVnJXtsD2gAhR
WNqPYwIjkzSoUVJFEHtQBH1qYGLiJ2ce9J0LyJQY5VO9jKnegcynKEuN3L3ZloVz
AI4JKqIJEr2sikcVFmaWFZahax0a/aSo/mB/jZvlcazUhcQ5dRV4Wxn4FuOOKvlA
uoahycLnf5BzYw3GJgkKUMg50fdy2X87/wyc1aR7Y8Ao0JYlE9og/1RN+ZB7Ry9f
lUnEyFSNWkPx3G+bU0m5sVDnbr+sEqaKYfO8qvbb+RVJMFTSAEHE69Wq6MGKswxC
RmdCwpd1lLv2QMosU9SO5HAwlMVYUH+nDLdSs2OM3hQd707JqbLItRxfm7LMsSAm
0hxkFV8QhRxh+/3CsnuDbCS4pQsGS4xGw1F3s/P0j8R+uLnbMwGZpSqjUneq4dZl
65pLUn39ob64eEC1T+QwFdTuZgL8slrJT+3Qzh51y1WBSe2JtVO+TGE99nrLWLEM
u9lUFMgdUi5Rb4xblwINYrlD+HEalI7p+Mbzd3CNKaeTlRS7Wlxn/xpCXi9ov3WD
T3OaRw9pTiS2RmaO9lJ7+8r/f23Ja/wLygguPgILUm6DT/aoN1mps4mwX45DISoz
SB2JgQrB+SwEMd3xIPvBtdWIo1ZhCfq3UgD5Ix2ZlzlMTmHTZxjXHb3hxw83m2Ye
LzeJzta+3aFaeikDS3gdyGDCQrSBOukgVqBPRGzuG5EyiYLXP8/qmgiN/E3rbCMg
v74Ya57j9EvmJ5tx/qE35k/OKZ500iJm0IOpfdtR1/CqW2r8jltVrq1SjAZvxEKh
KvgwKVzvUKGET37oucYFNVIgIh2e/Z0Vyhu6+SxRFH9EQUUA3XrSclXoRw8Frfqz
YdDPSoBUv9QkDE06JJ6mL+kf/HfzVB/XSb7T7Dh9mQpO0cXldrEnOaZhztfYjqgP
TQxNHK/RI6Kfd+PQnc9ou2lZkT0t3NWG8pDLGAqLQp8K1P8vKtYmvuKr+2Q50P3c
3aLipSf/Uitbb7mC7w3tlVlQ5AvjO2OaUM0uXEQ6UbVbcpqR7Ktkl02PUtLS4cRl
eQqAwOEr1OLd55uLd3RLi/tygQXlO0brPYpV7QRl8ChdKqRcQ/81GToOLk8JyrGf
x0N+RzPmSuGQFLmaKLqKD4GRrU2tXEjqyzLT+f30iVw4q5xkJjYj8IiWOTVbrn60
ppnCqsh7GCIP9FXNfeymeet4b5BDCdTEXnpIsjphJX+NDZ2asd1I2YuzreDu345j
fbGYybrPgu92//DZ4sJjng9fOt1EShEZaIRWalu9i0aaq6SHaRplRaL8aTvLE5Uc
WyzyDQ7bk16N08xET99d8+hayVPfouyppZvY0uNjm7TFbPboFMRgmxuH9v3qxKNz
R2LMAVl1jB4vKfIqyBw6Kg814MgmncKzu17caFcYyXpHLI6XU7GEszR5+5yM1lvS
AcZUfFg+Kq7Jr4cFhvXY9JmRtNR30WHWDEnC7wUH7dQRNj12aE5bsIoM5tRSj7MR
Ydd4/tWhfq17Aa+9VGvs2skuRVs/5giXYL8JSKq8191JBwDK6YioHEhYLoWRLFo5
E6TE0fOmqSTbwGt7Ux6snW2oMEt5HdEV4n881+npOllkpS8ghA/kHQe9HCKfxAtx
YxkuN4/ngis/bS9agUoe5D6BgeqHZ350aDRX6IHwTkMYw8m3VKE/0eCqTJBjUgsb
+wLM4vIDVJ6Hqh1vOZRNVS+bOdFslC8opTDQmmf/xpHdf86sL1iDGI+OlPfzy0uL
xshqGLWYhLMuuJI6/Dco0oxEigmOSGTZUQy2Feg6zi/T5aUlUs452+nx7DEogxK1
`protect END_PROTECTED
