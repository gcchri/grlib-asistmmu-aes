`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E75M/vj1VdnynHdtjjWZLPETTOQipRAYYjXnxAF9iNEtkW0YC3kHH0CHJUBayTcP
7H4qwqJH+lWLMKPXasty4qYgtTBcEn9T0MCjWz61vksenuIb8IfJvC91MJ5sDP0W
Jsce45M6cetHzxDgn0aS4UM6CzHWK6QZ8xydoMJvZhwN9V7sFbcWbgdnHsYdkjAB
FM6MyIM+AJnfwbQHO0Dj5hojp2w7H6hpXpzheEEcLQ/NGHj9gHq8DERFLRTHlwE9
GLHjDL4/bWo3w6W8SnVS5vFPKVKM89iboqVTXdbKNOPmPb4R6EsO7rG5jhT7/vIZ
ezid+yiTfznTltG/LK7neCh7MZzUMkoG3TcwYmwGNE0R/WqOGHuKPnG4u2awan3B
`protect END_PROTECTED
