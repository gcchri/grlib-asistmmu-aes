`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YNiUga1Nmr9wW+cxVViJjI+6Fl7u1ETYciNk7qiYQjjvj7yIoyKnMpJW4TG17aGB
6G7Vhdr+B/ilkH5xhkgaPGB5tiqDGuDM8dLEE5z5pIeTZyMPnFye7NttDPXas/cW
fb6u+hEeQRcf6TVTTipw12xeG4he7NCvytv/jyYa4Qu3fvIadvuaoZSR/m7bmzw4
xFLsTGTynnNRQ+nmc1PFOY7cM+rwbx9FYkoawziZnaQdFL7bnxR2VahG3u7pe55n
hSgKj4q4arCLfhXelbf9HR4Qh0zo8eSn2Yc1gyhalreeFpo7cl8rtHV+lI2i0VKO
9/8CQsoZ3GpzliI0MvdsQlzOAd9p1VH0LE/+rpiVqtA=
`protect END_PROTECTED
