`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/VmN1rsa4Y3G6y4O+Ooi61g1YGUSnGeZxzUKd2QI9nCNVkLdX+E0A11+1B7fF0+S
YPFyjVvbFIhSN3GNorgjic+Rr8AfrVHId/cFqdUyyTLla5UpTyDnh69P/w7ZtHmK
5Eg7LMVc3IouPIkBaY30AypjNTt8+PuxnwTqNPa1vjUbhBvcDDMl0oGkGTMk7qO6
82kB4/LCjg3ts46uXFdZ57Z4gjT6v9yRsP5N3wYYb9v+mrj/IHz/9Y8QdzYSWHCG
joArrsidGtKOgUvYSJ0Wgf+k9Ywq5JoYsaIXk9fzkjZ+yf6wy1fHqx476oxts/Ys
x9WmVHgymYO0d157jiWjEN0H7myWRHS4XBZSJ85hW3YQGHsPznvXtmav9CleTmEB
mEYMxzVz8iJgR+bh0ceHwixPp7Qk7z2VkhOJvHNzF/w3surOq128sE3Qw/OJMwXp
sKVuZvIYPmD1ys7xOuW6eFUE4SLR1VD314Ul1VkTTwBzKpipMC4Dke72ii+8l9wk
696namHTR9tLQ2oIW3FXqNYIDkuRB8jkXAo6O4hV2UILH74Y7aCqtSyOetzYhwO7
F+TDgQ3QPliQs5rFP61vsdzmMXdaE1JSDMJGvKZxbYpi4oTTaIkXgav9tiAI1Phd
6OpmwF+kyWHBAsTWYOBdCH45lpMTb5rbzUKGnRDiSJs82t1RQllPDiNwWOJO6MHY
7t8XMrsjDV2Z2B4QQtrmCiwGebl3h2SoqV5bD/cnDIPM6Z22rlOrOfLMlDsSsYtg
t+8r5RH9mxOybkYqpR79/w==
`protect END_PROTECTED
