`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yUIs5YGNLGR+MNoa/jNzEBqH/4pUkbxECe/i0OkHX3FmqHzliuwUfgWgMn1JGIu0
v6AqljyFKUhu5a9k8Vjrl8Ke9M+LxhsD23uusiWoBl0HHa3FUfzIke1mG2tmCToW
et/EqDeDMvqpVnKXbSjtK13/KhiIhxDZO+BFHBuGYcq4tVxxBTcYGGtILont7cJK
wn2h+vofXMBh22RNcn/n8nUEmHsrF3G58IU6GOd7Lzemk8k2oVgpshxgLxixkHfs
sQoLqkoa6AegMHsjMapbXsWEJXwjTkbzTWAOskrWrSYxte7U2B1OZUIjT2ymcSaA
BNJKujgdCa9ClP/fwFsVBfXY1qDeQiqx0rL9mCNkngqfsIfbkXV8Z3g18G5mTZqJ
6G+ET5ByvQvXzaDe/0tle0LVgw1nDLG7euxWIDlvp2f594tlyUTV2uVVo0+DwS4v
hYjQiC20VOSr4yRK9c+3LJaWndc5GQM4E8CJ6/igEonBcMWkMDfQCzC+/R0HiE0k
MkAQ5cjLKe0N9/TccFHxHrkUZoIF/JHeEDc+aqteQKN4x3HoIYdxOvFR6tG5Jd5Z
gSpP/mDgbd9T0oWThHhkR3xR8PXU27QUHcCeGHf9JZ1Sz5rxzWHMzoYc41YkQU1y
TbUSmQ5HLHyW88PvBG0QKB8h8VCG8fSrlAeMkrwly2KDjzviABkRVjCK1VsCRIeF
+N08Mm0hKNsG8qmPHUwDGOPyjM2qRKrkIXiEXXgoboU+ZaIySs9YUN/FAsP6coPI
ig/6V/sSmyKx0XCJBsoocg==
`protect END_PROTECTED
