`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qxUxZMrAPg/BGmg/ATnsZ0UmT6sX/tEr4P/LBagHWXJK5RMN1HMJ3FDp8dhK83Rb
6S6EVxqiOfQpzxw/kzEXO3SPsqDXU+dtFFtL8Aj6cTM1hE2jDY4usje/FYR+MCsE
IGgedPfuXFjXznIqZg5azoRQsLOGCKNPcMumEdhFLyt3fqEtP6xbGyascv7PTkHB
p+dxhAWtY1OsA50tLwQtERt+6DlqZUj0wGBBNZWadTLRIqQcthS/A6V5aMV5/M+w
xKfXrd6s4kdWI+4hsM2eXI++7dtXP8sEQeSk7NOHySptSeECy35VkK91Y1xJdhU8
u8BXWKyk5LMez7cvSqAWdSDiNTOy2rVGXxunZWKzSBLRtN0jE023eLW3dDu+DXQF
kbSo+z2I6TGzQiS+vpwUk70Do/Pz/knAu5Ws63VJHDSthIJET6evgCvPXwqI+ap0
p5UFo7jPQCUDQ3qGN0nz/OoufSJtwtUscgzcqHan9NwXlBFh63L2ZkpSkrGjh4cY
FA8ZxXkE+hd22B+KIzPJRGoJWaUXvDXA1sUlhasl0IQ=
`protect END_PROTECTED
