`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QDkCWycqn17tq8H9odD4qxliMuvzgszs+BD8lz2efXish7q5cE5q9cv652tpy0U9
H9dltN+KyWNtmTk44Q2n7r/Kr4WmDYEPNpd44psCLd7C4rJqE/6PZ7S+S0N5/i4f
23ClYH/0/i19Fn2Gt4CNscOPNr6nEuUyz3uEAZgvaC3L3fQwtVGTNGogbwdsyla5
lFe90Hy79uQLm+SLokOlnVzXC5ifiuxUUM3Ecm5f0nnwCSKZ36SJ/j43gwYtvdkY
aDkIsOEkRxtwhaKy5AbcLhxhcM08tHAhE0+spVFMZNzXjFxZOH9y0baWZaiRu1Tz
F01FLHa6wbIGYXRU6UZjGCWYNcW/GYffJZdUBEJ1k1NPX8HTS9+hIYHiu5cK5UjC
Fff+xzMA6QFX2Ob7BoegFDk8/aaeI1W2rmvbQGyGFQo=
`protect END_PROTECTED
