`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fg01Y4lyjewRgd9s+6jkmtvxzFlBIrZz2BssYC9yWAbVSSybMZ5aNZ7sKXquA4hR
FOryrs7Y1VASyt43yObOZ44Mpn90XDCKWWXuXfKpCp2xEAdq/QLWvHbTsbzTPeY8
e362Ubju7MrJaHOC3AncoSuwLDeMr4Q/x3aNhdUTrm8QOGyvfgfgsBGc+EFbR7/L
3r6zCrSVCUy1npdGvvY3sqwSNfs12ePlx4951v4nMf2Om3e3+/FmotpVPhnRaH15
ICC5gHVjX+O8y2T8Kb8XFHVIzCN5PBpIsWY2aGlFGaF21GsXF6tSuBteu1ItYTW+
fZahD0imqXsjyCGYrBq+5wHWG5PFKNo1GrR0Copn22RqxMlqpdPLbWIH4ncD1kg8
lk5jDx6uY32T13BpeXruiTOsCGjCgbnES93bj6A7ieAj61lIZyGtfBnzIFclqFj1
5Mc0mvX4FGqAVALjxA1wfQmuPTrMJcAeKPU40KqDX4u9/jiCt66dQ6oJHksu1Xtz
i4VLOfFpSvi7hH+DgkgljKfxJnsVcuZYKjF2SMXx45IcnEZZ+BxDBQ0zczDwi1Zc
wVpf37aYPxRaGz7PLNQ/ltxy/yUjTcTT9HZ7TwQRD8g=
`protect END_PROTECTED
