`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u0sbyO7fbbendhzm+LHzPOkXZIAJJtB5RGPi3O/2T/ZIQqsopacThl5I1AQnzWKx
bW2ZKS5y6EYtsTZ5SuuWl5r6PKClVmf0MC3B+ZFmiDj3N6/Sy/G8NUEaz7AiuxuT
yOLmESK9Zovz+cYqXJLHWUvnuGrIF80JWl3CFwluW04Vix2PITvbHT5lUatDQFQs
9ZBA1ySSW8gNQHZvlNmfh2GefzfCFYYBd2Aj+CGrdPQ5HVFj0xCu8+GJu831ADSQ
z7kNlhCa78c+iLqdbq4BHnAh8ZKaeaCodGr4j5KTeCP6CfNCRV1Ecadd4wwdgpTY
9TtyuE12kmPC2wUAh5VrFeb1/WZmYPwtSdtRbOcYNSq6EdIfLA7FN+P3xOTu4F7r
YyL6wvfF4X1dC2hKkjm/gw0bRucX9OeGedQRAeF6JV/p1Iqg4klF3a5uPldl2OYo
mYC0areDr0o+x7chuxck+7D9e34FmzSHs89z/AA5WKuaTp3yDFU10KCAIU5THDLr
H7rFNmi74FPwC7ruKS+VaFFYvHQE1ffIz1l5drzFwHHzfCU6+QSwF58SsoStg4U4
AcNShMAD2SpdoWwgwXhEEIGMYYtn0ZzvG8TXxKlnUWqc/6Gf2QTyXWt83Pr6U8qQ
k1UlQjdToPnVWj1Wrwk0TquFrM/9oEE1nnb657d1WFnbCQg4iuxsW2WPjfgdvpEN
N9CPU+qiK4FIIZWPeJci3RhiuHL7cZYACGteFB1S7rh5KtmhYl3vq7zZu0Rhngrq
`protect END_PROTECTED
