`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eVYB7zcd04Jr+ySWx5qImwGpMpb1yRy8/tcRSFhhIcV8RWRpq5gX1T8MRZAmsGaO
uLCI3L1LfxhqcrKOCKv4C2pT3yPl97PZd9VMW08e8BFGort5Yy5/hIw1V+rDqXoh
uxL85i4bTrQEDksS336bYxyRxM+bukQWz5dy8S+uG7ej87VBTnUry631IxQ2GLld
l1JVwPRTLXQo78GO7J202Iz8vDoxyDK53QfjcHPQn2wkUyfb+i7jDB0F0AZsJLN1
RG3wXS3L0QapIg0Nvu6dYgdOLErwVAW6hOpxrlijmgdhblRmNbvCz7Mg3R8YFsJY
`protect END_PROTECTED
