`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LV67cjxvVLFisk4pjCu2l22hg1eLI66cotq2oykqnwS53zXeSafrAda74YPeDTuE
s/1wIwSjPKhBe0c3pziMkeNDSb1EFe1YyTRutIMf9VpSXAjO6rqZumQ0LNGZM3Ku
hZV7qKQaa3xCjCwrZTv3qQ3X/hd4EP8dqcmHJ13VAA5wccGtzFRPlIcLXXXo3Xf/
hXIXZmA8iPJnPvAx4kQWOfequXdrtopSQWSM4/SkIv7JqkTl7bWm29N8/8+bdpG1
IDmPx7+LElMqEEdbtPASfYVy75pZqlrBUiG5/3cdV6XqwpNTJvYXnNmYeSF90gN+
`protect END_PROTECTED
