`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eaYyGOiewoJkpPwlmoNXZJ0AEMvZp60YCrXhEK/MSlANGINJs+BtuSdcnIoL64I8
BVbxCihyqc+Z6a2+L/LYS2E1Nz6dusQ7LqmWLkzQTvrNp3dJTk5x5aorDuyJq+Zp
2TOyt1Gyx+z9OZSAfksB8Ru+wBtiIhxSZSKqTnJTSbuNEfKQYFzbYmq9CrT6ufyU
8xCWhrv6VRTfksRhqlHm1TpxoWnJH5UD3cNdd3qo3tg3ueb+nBCJruTZ4nZSl5ob
TVP6q78eMYBEacG/OKbhcAIL5GT4BQEOUM9dzoI5CeYp3Wnf7cRNGLjUs0OYT1pY
Kw+a6EA9bfBI9w4/rKdv0/DXBceP9nLnFq8tXxCNxHsb8B5ZU1gWKnMDcYMLiY45
Fed7uyyTja6lx4SQkfsyfdfkl6KHQTvAXKedHzXs5oKUr+6xTXdD51Ni34cnMP2Z
lz5CKG42HIFnhDhOJHHMbH23IFlZZlrNIFl1wrGzEJdCIE3ZvdwpSDXiBsOfxWPB
iXyEjcjV33M6Ex19XevSxDH1Zz9fxp+sP8E5SV6t9DjMIh4QeeXKUJ35+h3raaZG
VKyg9jbmPtn4uBW7shKlh1otYfH41gR0lNfGmNvAPpS7bqHCp4sP0Fv0kt+nQ/92
u2DkoxG/8Ny6L0Q10lBiak52ff5oMKKFCz+q0Y4T1E3bFvyt+ZNXPfnUejy7mobv
opW06uhlLkktbZaw2OeQnw==
`protect END_PROTECTED
