`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LaAkNdK/FH7sWUx4SUueIXgA/Q5m2c3r0EhJmvs1mPsGe5abunzGIV2Ufj8kKtQ6
GvmHjtUEUjUb0fYAed9n2krDYAe5fj6qqFPsPcQGwfE70BgaOpWr1bUdiFIiYXkK
Pr3sZP/zgWZczwMeRpFe5ZAniYarRguS2SUGsxfZLrLBkM1AxwUWLUxRjYgzTmOd
9j0S+jLds4wykknXVJgTA9WSacMkFmkHnbVbZAuQV2uKggp9rg8x3cmeZhbMahR6
JfydtuS9mZUTq5LGRGz9fEIQnJI8WjE7BrFL/ijJIBk=
`protect END_PROTECTED
