`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o1pZQOvOPtB4pqCy9Q6LOV8FmSeDMijwr2m/Ram/GGzGq/g7LDumTKtKZzaBNDZd
25SCVp4UfYlzWysip74hcH8m5p8i/iJ7HU9K9POpM9K21LyOM+47A9mHnSi0biZh
QJXh+/JDX9E4am/Lm6xVdeiH9L39+XzFlGcaH4Zahj73wEeHccEmF5FoBr6fui+E
E5Pr/HGUefWyBq3V2CEhP4v6v2JiSFXDs24ZaJODHTf/YedTq8UtoesTJ+Vo19Fi
Wr3bFqWV23w4yvWCPWbKLakIKUa6ifmtfCCszOJza2nOsCDJeNI2yRUsE2UB3Sky
zlarf/YHcDVBNS3jG/hUZCgnAWc+TBavg11IqGaBGw88m+Ji+mtCS27un0RB8XMD
0l4VzLga1roBxqVL/CLNtpBhYi3z2Wv3c6/DDl9KSNxX8zC2xsyt6kqOgtjn2bEj
2rGXuTAhTZ9JcvDNmzzb+iyx46zI7XWxJklW+m8B8yl2w4psOkwHSmehEpKNib4N
AHKNUCGBEnsAVVf/lYp+PixC1gKMUt4Tvr0ifutGmTggZtga26FGFqGSt46Xqyv7
tCFMzlIGq7j9AJ8PIhjsJnQlMfeoqwghz2hIbYVjYbCgf0etkmiffwGJpWHP9HaI
ni2iwJGuHA5FjGEisS3QHmVuS0Kn6DTG/m0yxNCTZJjDgsIisjDutOe1Bw6eZxB/
qwbVd9S+hVg5m4ZyN1yaPB5YhjgnZlvQM8q+quaP+TYoXUm/IZ/eSYw3I6WEDhIt
ugCMrj1Dzt6/NomaDHe/IkS8N8XktBTQExC4vHZVExIjit5BGBpnjFHX3aiVzvqy
cFxQRZuwthdzgOYjL1in7fg34aFISDU5g4mIuHAGKfy5BxhE+8WSEFKsMwPBqHB7
4MJeZ7bnh1x+GLlk1Zr1Xlrl7naSyxPN63ob6b4ESYp/S1j8BoM152RPqjdS5gj7
9MrCpXgXN6fF3GGI0Er//V+U3IkCkkwbPUTkwoxEKyukja+vPwSnysBbAOVJhcim
Rz8wFDQdOLt168nUjb+X+o2R1+dLwA+7W8Petm2OEuZTkPloQnopD2scmPF5FAh6
jEe9jomL+uMxLvAPyLmYgxaoQYbI1Yits808FAU3/wNbFS3vw34B3vuZZVQuCMt7
hBpVywcKURDAKW2t8IwS1Mr/dTBmLQRmFTNStvFzhl2UpvK2O9W4e+56MFXnZm8v
Z5fQ3McqjLeEdYgwy6ToEpX2WXh9Dytpn6SvTKh86gd+cH+p7MHT1JrKLrykco5e
Y9CDnmVNHcp/mLuUJ7lrRT25VUcBuf9yQRDImxqVmEXohSRhDADe+n4qHVDkGG0t
7CKHamaL/JEnOw4sg4ehyEoksshb6xTbMnjsU2W4zJzWMbJlE5v3ks+mjRbvVePn
NaCqPH+bK8cYF3jg0UqX9Ok8FksbnmioxXq7IPqMTP++5BlHCemDXyBrNDp+bBnx
PeVG2qGTOZs+3VSGZbF9m37Iz26S8W1E0mu46lp9ARSzF5MYKcxfIsQPaOf3yLY3
EYy/1uXcyf7erzPe3HrOOKNI9VZoWWrrkuQKsy3k17cxwQRkHEMVos+p3asMpKbj
XWzkao/JLyajfSKQDslx4xLzHWGXQjP6JgSBWOldY8AaTculwWNAXt/hCQKHxSqS
FJfP49ck6n7mS7qjzCUmy6pRAqOiNfSClrxVoXDDRCycGza6z7YZLvPpGaFTMJM+
Rrcr3BQ+VYmLuzb/7dfJ1V1Bh8Igq/r2cNUd6VUlEn1QF/wigC5ady67T6xlN96I
ZzseXQERz0rMkUfdge+UUmgdM/ypxCLAC/vIOsLKeM0fXG8vPI7OPmCRHLVlV0pp
Q5Takoff5qB5cNo4wa5BXtPsW+9R/YnlKInEnNyobkrr0vfGnN7qIwNgEJ9ZjfxD
QVzsBuJgHOVE62+oJmoWT7G3RlNOwOvdlanDlUKTxvEX/aCpTJUCY5NHB0h0zV7g
g96jEvR4GzjPOeZZrifKhGx3bkv8z5o7T6FxPf+FrFW8nvq2VOyMLP8QBKLFQpda
Z6OLxSFkwUKHOp9W5Oj9XKu3UfgOQKM0/8sJ1YaO3mH1bwBhKMGdYgg5ANmp2UBl
dZ97AKhAVcilFZEvzWxfGVtlgHNKdkMxINCSKo8nedVmcF40BKyu9sndOWintibS
BKMvQsSF+Fl4fzh/bDaNr/TsvAThgA0zgZt5/TZlqQCFRVJl/tHvTtW8JhnIsBvu
f6IPiQEGGK9JcdjRS8zvEyzBge8r0NdfoDRsWvqJDRsfup340eC5RTe0/CMhGAvJ
5jc1k4b8Qh+GrtaCRUImrnD9EZySLsqe11Q18G+X7GYLn9Kns3ICQ5+eLsTGtiq5
O+v9FqYsj6JKT9W6lxLdaK0PEFy2ZsyZVS8vdL93nwdfPj4yGeI0fzlydTHr2eu3
GOqVxOpQbMnQxuJq//ljZECQFG4LmW6Pi8DI9yEBYDIBqJQGS/iR+kffQurbjSmW
eJlzGYk+c1bQ1f1oufRrqNZwZ4kMX8CwpJMiOx1yhDOwiDjfvqK7MKL8W52i7ToM
SymUPc7SOG6JPP9NBDDoKJiT0VlEu676HZ7JlA3QhfBuC+csM3gWPjeEZvajBEgU
iASgVG8TzvZnZ7jDePjznsLv/A259KUQLdJU53dZJZ8qCpoGXBrM7yWruZAXqXmk
+xWaUwisR44j3U0f67U9FN/HknYOZRC3oKBmI19UMBcaMDZFvc3HlmnelDABUbMP
xCcUhtCX2OVEMGvzp+z0zjudO6ige7xFs6WxAECY4B3h9T2PACQaPHxOkrLHnIk5
AXmBXCyR8Zg/41xgpOQe1Uo3JAv+5EvJRY/u+MfztOC+AaWaapZSp1Y1BCB3EM8K
OOgc+6YOH8HyE8TYWVBCgmVpM1Ol+VoqJcpX61AX3DV07p8Kmri1Po7EKZDtr6+0
Uy051+NCWWMfBU5f6DQRZQJId46XdlHRrrRpcx8SELN6WI7yE9tziDGiX4SXw1hl
updo01TswXRCoTKDCRWsYYpAQ84IVmL8lmHp4OPhe3PRO7QBIZ23rKbK4xgZlSd1
L4Tx/6F4Nj42u6wygIQIANeE9+kTx6QZ4kUvXnEwA/ZnyP6s6z0yzNAjRGMEqoPK
5bP2V3LBpOLhWo/kvrolKMB4SJ499+PAIHJUWIRFvnJcmqvarwrTX+y7JYxLogir
dCTlv847npBeyLp6Sw5r9eX9F+X8q+zT4yx0StUdVa0GRw1NAvkbHm/ZfmRFQJYO
tIL2Wpak9oyzt3i5GesNtziBk9arFGEKUeP/e4o1Vmx3yTuxj+3SqvRbZ4/8CTqo
FXQwoywsdsozqpCmpz2pGKLrMn7rhDrix8lKQ+GNkWuUqQgnIHLR37Qy8z2+57WY
Xu4H8nrvPdZKBJDQjeuNbujaIW73j7Q8He8CERE1NkCRYW5LcE9mF/kFJ8BDAt/7
GtLT9kUoNa+oUNgXhHFAQeq0kUwA6oJa/aw+Lp3KUxdjbeShu3ci1tY6wDfE8LR3
6T+ua1XL+qRkxFi+ZGbv4EV76+Kh/kfB55YGGRfQ5PdEvVUfr1ATnYPy6hydXdzX
ecpzPABwyHzlCvzjVSs1rRdNXZV+TqpFK4+zGgEbEKfRvzUSMCYxEcBkbByN/fJL
IkOvyMWkK48zf5mr0fcmZCtVQACvgm+eeJ03Y85CQ+9ufoth44xKxW4UAD+1eNvn
iOnyvyDjVFkvLWa6v+qGdJGNPtl9gxvPPXJxxez7pKwmbwGiPbISGddsr0x29BTq
dACm/yt7TISbThamGvHMZJioMp0mQf/jMUh58UIjx4N5ZJUOG84o53HMWBdSqo0v
8+Cb6owDuvysQ7ci4EuG11sN94aMXBhmW3VKp5TyHoRbn0KOA7K0fC6CNAJNJsaY
bU39H5RzrcWNX4tzG+8pzgT6l/JQ3i0pSDsQwHSS3MWjzzDfUjHwVcgZd3tUGVQk
9ifhP+aPUlM3htduWelKmo18JAQVzhxBY8216ZYvrAANdVPTDCn+orPmD24rN+bQ
s3ItGy6lRp2L14izEEQICCOlrGs08DqyzXEQ3Ss6zurXnRjzU5OixP+qAli5BtrK
MeuKkXbQX+kL5oOzcuOAdfaEGXnwAYuY4371x/IoW5NH+yrV4walR4J3lJQog9/Z
SIiLk7nMM0uUWYXgAhyaBi9A0N/J9gNFhxlLNogf9kxythYkF1rjL/6wYe6aj/Ay
E5Dm6mlTfS9DF2YUjELDgznXOoGDMFEakMJJjBWaEdAjzqK/NQBL8nwpQZJvxIqb
ffr1UfIQAIw1C4/SA4PqWpEHcAxeicY0tFnaGQ0y9qRQEh6lS6kH+b+aQ106y2qj
qNMxMA3Oo+wvL95BvTli18UJTJTQ8+wgCarBxGnR+FFeLy90x+OdDZo/nc1ysgug
dNW23lP3/eBDnKyO4r8dDGhj/SM4urChD0399428AqAtvzWvsLSHQRNyQMX2yMaY
Nn9WrAo656cBp7cdu9aH2cJ0mZmeAOZELaMScrR/55DaYjGNzuDE2SGJIRitovVa
II9rXGuG1xY2IdrL98NdBFtLO4K6ghuguCk7MZ8RYN0QyyrXiOuUh9GbGH4f4EfM
sSJPL65/xRoDKpV5rOuDzHOLQkPF9IMVyreGDSprGrWF1bQDFb2weWd5+2MfXnUj
QQ2XoLWC3UKAwCISc9edaXmu+yjsomp/GTXY+JF/a1JPjHWR2FW1fouzhqP5cXom
Z/23o5WFwLwxP1wd53/gN50Y9fTmb5TySDEPpjf9AYvaZ9Tkfb5RxDXDX6gyPdNm
PGspI9swllrxIH00C9xmkqaQofO/z/3pbzuiv7NbqoreNAxD1fmcsX0p8wlIoCGG
XAZ9E0TgsL/8ISideGzQyPB18w0GKaXJY76yOfVJF1tCDNyPSTIqbtNitFbVuJ0g
s7ZQWtQ0jBBLzqjbPQisYkKq4OOV+pTqK4n8spksPdkXChMPxC2ucBLBM1QFJHqI
wbW8Q5SYOpWaFFhs5clF9KZggod7r0gRoHDqEO12SCt5PrMvew/E2ZD3s2J7ymZq
v1cDtvOdM3BB3gdmZ4d2abf06mSXxg0BiZEDPZXkeq/4MMwg6OdOdWJRK3ajSO8p
aSe4rD4r431pq5xWSR3jf81kOoTvbp7fojrSnl9jApwhaW3U07najMZvRZS449qF
MDtZYXzXcvSJKKBJSNyNyDeifeCkJUT+hwCybqrKISm3BeuyOQVzQep4V8OXpglx
SKGQzxEZtSUlZoy4GWi1JmOxMM3HxxLaKQqihPM2ldH2bCvR7Nx53zbLSsIJ+ZhK
jHAsVUlVzXYezF+4u9RuVm3amM/fRQx3917EDVF1+cMrFXPlfloToPIYCjpO08zq
t/iirG75k/1TJzEo8tGFEX0UOgJPOWVkWJGOhvicafU=
`protect END_PROTECTED
