`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W6dlBlBuRyuCaKz1FXk1cRAIA+bQb9ZPrtaVxLIoqsYDojCuvlQ0m8/VZ0P7Th94
8K5rZ+ZRyc3OnqJCaqO1ItqWxzUBG0x9pCiRkEHjF6xq29fvc7PoELVMuyFawHJI
ROW9S+LFjgI1AmcC+Wz/TRA9ReUTGC6c8QXLAfz48guuFbvMvlbs3QTN9h+XDx5s
535mtxKyeJ2gTj5yAJyD47mfKBlbWGpKtSUuQtDzrkZwjsFRa4HjGBbMbeyvvXb8
RmkyE39Pagtxr+xHzoDNYQ==
`protect END_PROTECTED
