`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qNkrkKZ5I74wnkYnugE+GO285RfVxm2xSINuYlYk+3Xb7WmzL9tD0636SQTHZPqX
SQw4OtqXmpyVI+kVTJJjgc/31d0DArn9WG8Y+Nw6SYWBFyk9xP7/fk0LAuSeFttz
FcmH6ZwBoyLkgYchi9vfG6/4U39OPj9TmZHHLtfcD9QngKQs5fU1f+QYb4vLA9Yq
Dwv8guVpZUXl+B6hj0B7EQN6XWl4HSq9GCi5F6NkPMcbKHM+7ah8RpUjNkKA5R6k
64QNQnPVP0IHLXPScr9QndLYMlRujFAuGDS2Lv0QX7Vnq10UDqnGJHCKIZpAhwlo
6bmqt95RFdlcKg2hq8SgUKlJZp0YWO+Twrw+D2oYBY8h1OsKF/jm5MHF1o2aKdzh
u9q67RJfpbNHv0bqNBpv2afhwM3qOEHqoVCLrR+4fLJEf7ElU0r3N4WZnhImTt9d
RHYWbYF9cO0uJoW3RmjU8w==
`protect END_PROTECTED
