`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OMK9kwJe94fMgf8Ihmv0fZ+NcJ1uWuCwkY6hP0ZaWKrw6vtnlrwNv/naUEPWxp0S
C6TVhDaLGHLq5uqDD4x0SMy/0QC8vZ4c8FtJIt5K/jKhdgS6Yimzhykv54S6Wn/x
tlpFqB6TJUWvsF1Dj5HTDDepEN1W8AkPfbZT6kdt8EzgH9/t8C+g4EB76N5LZizx
bAn8dUNlpO15WII6Y/y1dqSJY29d+y/WlWhlMe8VeWuQjxgG9KZTZa6Ky1D15fWt
S3DTZZvXUteyrELLttmH4hFuzWJt4HUkRaB6tBHvlZDNRa9R6Q+pyLatxbAqJHWX
jYfrQDJMpaaDchKx+nMjXrgciR537i8X+tnDc6kqKcM5m3uVTdaGDF5pBrzedfJb
LvA0ImbrO18YK3qZQ9NX9LDUo6Hmi01ULtU52r13bcqKJQ5hScfmmgaJiTcSvwBp
o0wEvzrM5QJOB/ZwCybYc0m2JxWm1GDy3kLnaC8X/YBJPKQBpjz1rthfLwpgwzeA
P0uAc5eSy1enfxS+47/Mzc2E+iTOfplNMIsWnDlIXyVosAcObFVgbcKeYoNJIp96
DjpGEwr9QP9CRqZ7eJWCGlHfxZ75idaulB17nj4LQApiZpYnWH2bQmHy0UicNaIt
G82yWu8lsdAoWBnsbnLe2xAhj32n8NOcoifnol/2zhiGyky5ZX9kGbV0YH3P0jBx
`protect END_PROTECTED
