`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qDPut6/TxIx1tgvgsyAi6LAHw9lWsQNNG2lph2fpfUOikHHUsSmZN4PdKfKRmc/V
xjzTcKJbX+728RvLSEY4fxeksvgE0JgY0OAiPGdX27fFTQRoFT4grzLnldC5fFGD
rSMfwg819/LJfHp4aacRBD4neKl5bfJB/Nmu1Voe6Wi9QBy0T6caIdNDsXHNKb3G
7YL6+R4YWCg5R5GnKWbFTWPxxf39AZpEPcPR1Upnlaz+gzUQ+LXHkLidZvnSoRn1
`protect END_PROTECTED
