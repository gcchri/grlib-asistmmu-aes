`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7syGqNjqmb2ngA7JH0qarQbWQ5lRKNQtGflAgyHj7Vxx08NxxAf0LtSSNVgWAVto
vPmTYPS8h0uhH6cOrEnQdn2Zl+Avge6HK8tsWP/erSchwQhxRv8rSr1VoWiswTIO
d7UmT25iKFR9yZgn91iTJQiW69OCaNGYxQtG480bsGXlDBPOhcPZ9Y33Y9ZawgPj
PsLCpOwqsRQCgbw5Dm8duJbiGwVs8uzReM3WtpexHWW56mpxvi9pPgaCNa+Wx+9o
YuxWtNDwBMeCZpgo9D32sKtBAxGZvu57ocWfyNRryjnO5XwVAtYZQUGE0T77bF8v
vUVfuOa98tYPeHGnziiHw7MS3vjHQx+1xN2fWyuh4eBQuTDw7hcgFmH0os+oZjUE
`protect END_PROTECTED
