`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jRQQYh9iuFhr5PEAd3mm/rxV1piMd8erR7+HYCef8Spt4wrFsIxzpMiQXmw9CGra
/Y9VPadLIlkIMH1zOMkd+2zZYAOu88W14j6t+jCs4lGan0FUVb/PYehBGmGxf37I
+OUI+e5uYBhdOAI+HUiNhf3HzD50TMQJAOMmq67h+9c3pRPJErZNLqk0Y+97I9LA
27ysX5ay6blj3jU5tBVYqzRXkolRW4uJjj52Z6TrlQ6F3BPgVZxzHsBnaGQN/+9i
aDsBWXXG5sDWx7hxrECG7q1b8LBSYej34bmfICPjnCE3wXyrpHm7tWej/9Yy4N//
7SvLs0jcaNjUsjgJe29uTRHHbhQ/RKZWE6SlkedpP6sJkbJMzyjKQSmXd/DGR4gl
QCTKjehLp2s+Z8bKLJSaYg==
`protect END_PROTECTED
