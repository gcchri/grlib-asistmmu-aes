`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GeT3bGXjb8+ch/wSIngdGOiWaLTBqNOeZWxhBm9LktRuh5kIYyvIl0tCEWu7b9sD
4G8EzgnQPdXm3cZgBYlB/KyRewKAS8qK9GbOiERuI3eSiL2zTlyToVBFnFO5UobB
7mqJSoklNjjGGJYrqaWkWuhsoy+0pJ1W+CRwC8yc1epusg0Nos0zRTYbSn6XL5RJ
RWiyka45PoVW2lWj0BGJ2M2XCZpSY153CvnaG5LepWszWvap+1YTaYdmOGsyZMCy
NCrjw+G9TtUZseL32IFTumbJiGrKqLq1RoRS1hJqeRVAFCp8VNzfXuXn+FFi5NlM
da9+QaOiapx7I4cL2ti7JP7f87ygnV3uj/EvtUdIbzmmdBMNqapwHYv9NKP6wO96
HtoVIDO433xXxp9Cz9L14WvIMI1JEsihExODa6Oja0WxuL/O0yNGBeZjI1C813qd
MyW1e6sE7o/Z1gp2fmBQlTOrPtkdzXeowJLEt2SJulna8ATu8khVXkQa10BouE1y
GoQjglR2kzB7yP9YZued5qw0daqpNey6soJDWrn8cGG4uMnlFcEYmcQ5j3nwt+rN
X4/bHTrRjWQyO7bmUh/LwdGdy0vs+TWZH6TWmwzzR3Q0rHhsZjkvAwB+E5Xq4ycJ
YK69pmw3V1wY46pCFmceUR1zIdDgoC8cldbvGVytnVLdUSTeCKzhKSZvslAOrDew
5FeG61zPC1lt5v2Pl0+ZWOC/G+169QcR3YHBDk4KWkg3auosq7tChtnaVAXVmZ5b
o+Em+ZfsZbbD5Gpa+ZSsFi4s/Mcman9hzbz5WSdtxRyUYq4QOXsm8RvtqP5E9d2Y
nzuYRa7ZGxm/OYL2GV4h9k4WVCKEOgg//KZOKYFl4A1MOdVESqT10tTP9ip5nEN1
x/sjKQRYf7Aw+q87tFA6s0GNqm9v65+q5CkSsxpeB2+1fPjnI2uiT/dY46LpzHRC
Eer4wQmWMrnNhua81VXoM0xGi8ILHiM1MRqvBvSpzMbmH6ZjKR+8kmpx0H8GxX+X
I2nBBSah5wMXjHJLmPnv8tmbsKUEOUiwzcJaU+a9ff67mo0Xvz+RimNXsC1SgcUX
jimBMxOoubZtWjV8OXta+RuqjvRjMe+WB5LfnpyvjTF43FJBxCGDRhbefGuGs+bc
ChZB+Xz44FKmGwMwrFsC+AYVEDnA8/bjxU9wF61hFp7BIuofClENQeKpacxnGe2Y
opWMTPnrLlU7v3w3GP/VSeD6MIlygI96ZypK1gIXGXu/6UTqrj70QBwwmEry5Deg
vH2zIHa6QDDqwr16e+FO/guCrrbKgv3pMstf83rTzHCJBo0iM61S9l/qc9zXZwYa
Qt44dRn/ZP7r6CTv3bgvSi1pLUOlwlpKKWYjV2cWEZ5VOkUtVS+n3H8Eu3IJrlmW
Pa8hBT52YCfKx+oSxaROI+yiJGavpcnN08z8LUbUco6AhvcbCneq/RJY1SBs07YH
1AtbZJepJIj51KW+dwBhK+5tXvWSO8KiAPcX/zOUjlZGibBJd262qNVT/LXtGmLD
OfriywBSq+C1/FGjIryppwYyoUQ64KpaL13A3GSOGy3a4hEb/watKOy2zG5PZx8b
2/lvODe3FieImayvPYZOJv4mKzpwpmQ3RdcBfp2Wyx3a6jsakAL+0KOFbGn87cQH
fT8/1nhWNrkhMFg+AS7TqZgMKE/yFQ6gMfKv6hRag+ONT2FqZqKY+/Zszc18SlDy
nJDEcQcSZ4k3yk/Z9lTNeAlOXQJnleirwFNbVuoYa/owqvnebVrMMHea+36MT80j
lR0BWw2r2UuMgrd9nqM0ORf0Dqu0S34LAvp5eflT8yqZ8J6cgXWlTb6ujcw8Sxcg
ly2x9bitxj0FCUeHE5kNSVJmbApWD8HN2AxsqAUo9fGLTABuispxqIPHLnXLCbUR
Uffddca15upAtcGGYxEkDekGr4OZ687kv3x8/0CNytVmIbfzV7pw+rnktKxXSf2s
nUBaCKOiq7o47Vl7Eucsb3TRkFOjap05cpkVSxg52h5prpk4CVsDMCy8WrJrj10f
AqbQEDQnYOT5NCmyTmU7ioq3CkJR8OYoqiJ4z92ma8Mz9ogXQ5whrlTltL6Qi0VT
NOhWL0CiQny0MNXro+60sdslyEuFEMHD8beb6MHZnI6pArYucGFNW+u+2MX90/Bc
vPFgK6mONK7izpRscNZVn5HcH3g7HxucfDXD9uxedrLHfs4A41vGMhZdpI5+IB5Y
v118mMSq1i0fFMBFHYuOTXX1kmBxkXPirN75yea16hcw/IjNEcxX1nLixfiwS2PX
NXqWqFJwVmB11cx61zi38bkMFaeE7QnNalkNAczsbBNIx0nrU0Wq5TnLbwFmKfnF
pBPhrWyE43AP8zMBRJDUMegdyzH6xb7R5zO5YqEeYLOUzwZ5QBC9FYB2co6EG6TH
vGQ8rs3ID98QI9gtSAs77obfb0/+denqTvBXgs0tnbdN+JawJlkreJGax7PrlAwd
9U8m5ixcUY8zK/w9vRyejoYuR3visTdmG46PEbNLJRgs2QE7/FRK6dmHPA5g2Iv8
HxUBsaaVFhyv6uh3tFa5pTLNu4xHuydz7xRNX1eiSNENO3+wH2fa+bhYszdR5rhw
YNixJ/fTuhiosEEYuyyEWzsjVWyT3MBfaAmDNfCz0cSikTjiN3sb0/6BY5jioQXq
WSPmsQq5RYH9S7PfID3cxGQm5f8Asz3+i4GtT/0NP+bvvYTo/kVTl7Zybke3Mx7O
ap7gFA94VGUeEq5JzZoug/+cGmkX7HbwUPoRHZNQqUHFbwBli7q7t1BhgydL9j5e
SkTcrr2yGMxTqUiJKdF5rlmE9T60ER8znApQGx4YGK6DQhrw981bG6iLYgkhLtN2
neiJIIxXtd6+FpUfUN1TTkVSwwyfP0j/BLhB2ui5VySjMnGOB2P1Ijx4nJYBfX9V
AEJ6OWimVP3942CSJ9FrW32QIwUCJndk8MOgDtE9w4ATgpflLpz9lKcjM0HaauxQ
MPlYSflci9b2CDrpMm7+Dedno9mm+7eHNonav0DRUptMm6DyusRxuNJI+k1eKQIO
N3dQPMg1f3jujTrqZTQZpXgyt64ZrHd6Nx3MN9wSqHWwC6Sc/OWh4t4nWyVtvS7N
SkuZpK7oxBkTn2Zhc3xtk+e1E6UDkfBkCcp0mvFEOW5FwM3tCopaBOs7GAyyZLra
AuX8sD4zrcMT2l2IwYKJrbGMykKx8Dvw4usTYSGCu0eCu4+52h2rF+Z+8olDrG/B
ppiUtdmSVE+zp2GNclV0TyPBotWmxDKSpWomJd3ZQoZo7lcWdUQWDVyZv8W4+0zW
Wx8lBVDMMx2SRvF7KNQk+RjYGtRQEz1oXCpSPphDbgIDmy2+wB+sldfv6OUMWZ5Z
D+S0Z75uunDwiQvWnC6avowY6GhmEmu+mXOMQUQDuPFLJo7us0TJv0E3nGodOSDf
H7bO3UIoYE2NV2HZag28StHGm8wf00N9/nndiSWVv06o5SXYynduHfY3XQB8I2X7
1xLG7/i/hvHmHE6OXgZsA2aFctgEz/sJaQBBIS03R7eKZrYj3UFugPlQPTJeiVF9
5rOQNK1INqJPsI0BBF6xD5nXViQfh39PQNUhZLZOK0H+xsjv8DTL3m0vhLtyLPhZ
qLXcqzIM/0YCkCvdGZZiX5tK9F85DZERucT2NudIROAbf+5WpChsDut2xq0y8IhU
tDu3gf85a7XvfuXUpQyTxXQvUWCcDahsfg1EskUs1ghBvALjqbPOAzrFnD9rmOlJ
ZRX9eIRwxQtHza0TVP1Hab16XcyeIsFt00vVgY+C+PItLGbcYjMhmSPUxHJ/wDlX
UWmegKC3t/zmWMX5yqwVgQfl35TxDrjX3EMxd4DC7PXpxBToTLrMA5m2XENLrsnu
/IR/Yk7EGJM5javZE/oe0R6RvHk4FgdgFW0XRhxKpJZGHGe3+/pLyj2FZOGQmEYO
7XGs6D2VDyxHtMVcIULEat9Z8ZtOqG7HGUsfeOQe1tGvvUJ85D8q3vqsqf2eAy8n
bW/fjkuIB5Lfx4xzCEr8n3zcsqmZ24d5Px2HbmikRUcf9GzEJN/PWq08FWJsUIO8
iAiSIC6Y8Zo6EBVnFkDblL3nTLCyweu2fP+g6qQfc96HknlHVmvSBRt0kx3u3aG+
`protect END_PROTECTED
