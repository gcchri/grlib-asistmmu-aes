`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TI/zp1z+/43QWIbw2Ms8WLAbZZuQs19ivIlyYmAu20GLeBkyT4lC/Bgqk5UCNZKN
4lT20MEsRMpRLk81V88rpgGV8A3TcV102Owmrx5WhYTjYlvR5dbuGrnCsrMGNv5f
aVuwdlJk3+8XmulxUQC7mY18gnG5H4BByc4EGBYQESBVnJiQ55/lEeRteodCttzs
HfdwIdihQqTFHujR8hMkZWcJreo1KUFmOnTUqDF9lEJbM3f2gl+yFbVfuHUt2N1s
qyHqQe4DKoOpKplbIkEfZabjS9Mr2mjONfnMUAFEGzQPdNm9PyvFe1lslJ5wiKn7
Zw6cxtSjPJltxHqHROfbU3uFba54vhqr3jZDq75CQiBrzXx9ABk7rJQZsdxbRSKp
4bqMfNLrgltdZLFjwQoVC4kHo81JB3mAv42GzK0CoZQHoQ0vpYlZV8xVP8ChAG2c
AwV/PS39RQwPV/zspNCUp553+VhpgljJgzLdriW9kHYcz1kHmC6XihXfCuEQpVdZ
XOe3tQkb1h0ItR0OBGnnD8mkWTqnQEep+qw3at0Fdfk=
`protect END_PROTECTED
