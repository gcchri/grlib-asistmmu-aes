`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8BHCkg3nAj5Ml3jZNvDKapA+efPkLgDeTQayCvwX8HoHHu3Eors9d4kUfvYJDSm+
0fCK6Tgxxz1qOAEzVNYkUJd0SS0EaBX0i/fjWn3vEgLkffS9rcPh9IJsmasN7PMz
T/o8GyYssgLtsBa0cTx0IFxPKtoLIIR6N/m4/FrbwvjTLJQLSMXQ/5Qv5qEfSzA0
wTP+52JUSzMdXisY2W+ZdaFLA1QZdkwwYipotVBtsf0JQ6dRR+6+P/psxwcLfSvP
HUEr5ULQ5qoIIaiX3cKGkQ/yVhjSCFj5GZvOqc2PswM=
`protect END_PROTECTED
