`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1LcKSHrdh4z4XSNSIOf71MJR+3vUKe/cTv2Sqr51JqGuEDgbsae3aXKbLJQdyIMV
x9/X4vWK0Q9/Id1kLrHugmLWFbiUuzR43Ns0QEoF8ZwLhzyd05gauRHMw4/31jfm
Skbw1Hvf4IjlBxLOxbEwKzDbz/Vd2YpLBgwJaQuDlZGZ+LzJHIXxbax05iEeYWHo
sraiNoA8mdLAYcXeTduza9QOA1d+6G640HbZ2707WeHEw3tZO2GkSffCr+00NHZY
lyb299deT9IStPZ/jKDdNvgqDcU3wg2DTvyPGNCzVMHs38oCHp2P2bkiDAzTfG2P
YtkgPkvgERQ4BFdP4fIV6g==
`protect END_PROTECTED
