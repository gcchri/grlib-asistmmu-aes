`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BFxyT6j9sHDGKa8rTyhVyp7OCqtwnBUOQyxMhpZNeFN+AN17fZU6FuQp1YutEC5l
TAPqZ5GhIi7E5b0wzyHMRYpFkAN5z06w4j2Q0mUSQlJCpp5c1e2oGhP43HL00F69
YskkvgKgPmSCZjnSgH15MMiS+8fopOYnXjtooK02cnul5GelWsTMNvpWxRAip/Ay
dwgv/t3urj6iVLYjCdqAbTIR31LXmy9PISxh3sdrRXhnZxA0S82JteytICbeZMgg
XcviLGSAPjdWU6PugdGenTby73TttHA8l4dDYGvcwIgAEqIKIwWONFZNmpJDoD8y
Kdo54TpvFdrZmd5QIBb2YiHH+jwobPUzaulldTNeKApbkgctDNpos9wPeHGWvH9D
3LD0pfC8btlORYFcdyB2US1e97GzSBTN+UpxOk9yFLcMVawpYLN24szWga5kO64/
LSWv9g31OmedbFI8U+uSFOcRXfvPChEwmo0AcABEaSvkFkRzu7ZhmWZYaniFTX5K
RnUW26E2362qugdpVlEYudQUKOYkoPx9XotWlB/ClCVKnVw25I7UBa5sYgpr7J3b
da79hGHW6OtbvMCsLJ0rV4C/y1V5pNQt0rhTgOJswph6c0YkwI2HD6QCE3Tbnjym
4+a9zyqmAKlejrXX/qu9C6gyHcjWF6Hi6oquCZ3bsgOmSgi8hgCbJGYe/jt74cT6
QqdmeXLf6lyccpbbtOILUUJP4ENntrP3s03F2v/VtM4=
`protect END_PROTECTED
