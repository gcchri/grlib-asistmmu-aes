`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MKWTyp7Ht4ftYO3AWpA3CjHQ+nrjhrJo3RXSE3SgI2h1fC/H6f1Cz8jzThgyoNpD
2/WLYh3gUQ/45087y1Ywhx44EZC2U5AzUKBaTeoJtbsgsnHb3qlXQyeL7F8qoEgE
G+S3A4kQOJUVNGFDNz/JNWo5ExP9X3st/e+6un5f8YmmaGjxgDxdSHs2ib/8qPB2
VXemYYeaESLsWuEKwipvG0HJkzewF01yMQhvE3NgbkFsaNH5gvvfORXt3LPxBBbb
1iVOZsKjCYCn0bFo6nUybjOZ5DucRKoDwDxfI4Kmj+maJZMo0bcxbEvZSZBOFwZL
Uh8SR2EIr1zpcrDWGeAzxYO3cVNk4xDDYi3v45YWnUzsko16D15w0WjM0qznaMDH
cUp7Qa0HC/JZvsUh6QoUrBXmtF1aft3XigSLo86+S1fONExjiZixNgRjXQCy3ILZ
7Ne7bfxLQm9D5s+gejHJ3KMmM2jLK47d6Q66VwwBgE4=
`protect END_PROTECTED
