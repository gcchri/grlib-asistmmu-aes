`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5ClVxnCqH29LQwJGnF1NbLiSKjLaufVWeeSQVljmw/HBODsO3KH2gqUASuOFuU2w
x3v1lGWk8juwXo0MPyrOXlBwjY2pGmh+Rrwy8BlnmBtSDQCjuBXCQWxrB7+fZId9
CE+CpWvcCPNtldlr0o1CPcZ4fj3eA8De8Y0iBLyl+1bsp1escZ2XqhFdGU7CVigv
7YNxhM9FQYzgL7h8x6s7hO4OowaO9jFU/b2fLCJJvNN+tWjd7W4KZjn98TiEyKV9
6b7+frJYyXJO0rM7WZcEQnpfMT6fE7s4GlBH4fqr97ZHyjdQKYF9mjJvTx+G8j9F
h7DhnKaM9OaSRy20zPT6HuCkpK6XoWC3/ArJR8H+OiOmVw/Pe1Hrl3wsBGjw9oUM
YM2UOfYacFa2zSvTWo8yGwWWJAxa2IYRRVjcVPNbMSLELWvzqboZR7iCqGSxNYnE
P5QCycIHhox0PGCJw5sHymbHMT2zoiLPCjKSPjVOYjCqmMBD6aJQabISlHQ02Xgu
dCvdwA98NFiIyWPIrGKEJ2jY+iaVM2P0urnckLgs0LU6LOWxbb0K819JY7sNtt7A
ZZLmIoBL6h0FohGCgD/sKg==
`protect END_PROTECTED
