`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CsiArTaNjPykdcNwVohknHKTRex4UXjQKXlX9q2bIQjg2cv72+h41o/SBFBDHDCc
EwK9zGtzkm5i8e/ezjWRaPSUQVwqmWtxOqFSFl+3PD6x9JGBfxy+yQZXxaG/rrvj
vqdGFeZ9vQfBWOyQ5pWPm6wmFNyaVcMSJewOB2AyzL/wPyQdfIoghVeCdmMKo0fp
xFZB/B98FTx7P0BnE2LlGsBRl/mLRt0e1i8OWL//JlABwLz8JtPGJEmlr1k5Y12J
XupD/zCno15d2oLaBYrhpWX3LJ0Va4GbkvMbtwZKkIMvmvwXAW+BkAMyPrp6Te63
3Z6lHVNP3zB/2YQ2PUJpnob0tRPr0/04XhL7gHZQf5+w4iFGyXkFx+dyRC1+Okaj
stybCuMe1SOtq7T4hAcIqlo7IJPPP1GhKGpwEvzNOZAXZLK8tsmh/uzK9nUugesh
TQKLEO6MNUplJNva42rtShHhiR8cPFJ6+DcGxYzbCoxI6TrHuBoBvKkpZSNAXheG
USYqG0u1PURs0lqy9oWegMgCjftmB6wgEepvZy4F6JmUgpbqXJDK+0V76RpJv9hm
GZ43pcz2T5WNXJMBHzpPx+n/9VqOTC+s6jJgahDVbMRnsSNdon6/la/1A+qyTtq9
w39wU+EN4PTPO0CNme9twpIDA8/0NXn8BG94oCyOR2bWDd6usqp8WryxbM/JtFJ8
jt5jzRUI2XqI+TYvMndziA==
`protect END_PROTECTED
