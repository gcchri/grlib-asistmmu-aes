`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s4LrtHc+VpB6kUXOO82omkOVlfS9EiSImkQQ6ZmyrZ1Ry+R3dYIVPtbw5mjnYhxx
5sFLgtW4ADKFRYl/hyaMe7zX8zLM5vz+tbpUT1r5ATUVIdOtVnCOEzHyzv9BsfCC
/u4jMl3yu26LglAwp7tcN/fwfKRj7Pavph22ybqMNrhxGI/PrfMbdnzj0FdF/Wu1
V2XtDI+/xPXFDuUdbIHrZff70qlVbSdOxJ+KiViHCzOlfSvlfqvcmEHo2h0UE6rW
jvThi7VW3c2dwY3vXwf+ezemYVkEASEeub5zE+GcS3mvMghqgE+NGZK7fhcRJKHa
hvkhtwn8F3QA7ZBJHtOeAPUFg0xl/Nj0CSjcPiX90mWpPwvq1RarVnjFFNIqHHpZ
ySdrxvMK9T8HSehp/DXF+m83IukSuTiv35fQDxnomRz5RpbfyQuv1LYOx0v31IUY
K5aOW8pHyD3rn7b8wGQTtyGy+0YTPdMSYU8tZliM12XoyjksVnGk1fAdWC5m4GYK
dl50uinaNz27F97VLYqa3k7f+Fb0OUknocyvQ9hni81mkd6O+QQBz0K1IDj3as3a
eVt0xWbJekLicxn/BW16F5OkMUbz4PfKtZpwa2Y5TutYHDbigCQPMu7mMXzL+jTl
2R1vOmRii+xjqv1fYbpQXNtMF9FGTZMGe50AWR03u4s=
`protect END_PROTECTED
