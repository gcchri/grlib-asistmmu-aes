`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jUyshCU4SgEFwx5ZSo9GWh7o/ysBojHgq7olEhDnb51Icqu5hwy8M4OF+x5HqD4X
sBCG6r4LcfKGVqBLwcz62UUxZq4SrsILP1iiO+ckLtSiFn/1nnpLWwU8Tbxy4vSi
MtzkQi3mG3npQk8UiNTDC2tbluf1LjrI9a13MWBbJdM3sEeNgo/j6Rd6IzFAmiXT
iPtweFGWNzxk7s6cRSDt1vaF1mCxhrVCaRlpPFyI+0IVmHvrl+p5yBf923wRF1AU
wHqIKbBIorSUdN+jM/DdLWpb/KrdDVeWFH7hOGpJWq3sBh3mkeJkPmXqW1h1JX/+
WfTzxHLTSOmMcTgcJEktu7ksrmDnaDHjBTWDeL8xjjgJ8HZP0MnpndZIcbuz92jD
DFtih2ejPSz/BfXpqrBE04mcQQVpDlI57PfVrDtaiUSLc4gLiuUJkQUmgBPCweuW
VJE2hPqPeLRveMfK22hBzct30PwCE1l2zVQ3lfQ5wJnRM6aLdt/wxUse6vAqv0ex
f95ALpoQjWkzffl9habd+Bk+nBlvRy4x/of7098CMZKooT7m/lwHU2h2TcHpvbAt
Ng2F7peieeZkhq4ALzXlNIPpXDG2GI+aRa5UTj7tlH1l+MwyypFgsSVjw9rCsLQE
ru7Pi4fkDJbNDiVvLMU3gu5Gpev1K7PTinFgADtVPZLX4T9f1kAFeTBkqzIfrsSV
KwllX6PeiLeJoHR2UTQ5OZl1L84OcM/s8BAo2eMx4ilLDKMkFQowjZ6yh1tbnEHz
iGC49El0H++UFSrqTZg4Fg==
`protect END_PROTECTED
