`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hg3qpsQ6eDqVQX6bdzGCbJZGcFRR4owChc2NIE6FMXi8/4H6UspX6CK2dHxt8MSs
xve4MXZE+nYDITn+OJALY7Ek8lLQVgySEc4KxnsBnW95hAsKcdhp6YqnR7isw03P
mjkfNIiP8LIswo/V0X19GAc1JhBhJ8WUseVI3PEWsW3lUNWZa5XLboa09IYSuCAx
GVVqrEawg5uGFc7Nwo5TOm4B2jVLf11bsZfuUZUFolt05Q/iuvk5sIl1nCHy+/X+
nazD7C+lyiAb+t0Ohx7acgugQfee8kkIaiBPszYcOsJXlIPMJOz6S+DFuEWgveLj
85O2d9QzYKw+ni3eElgtJg==
`protect END_PROTECTED
