`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YlmkcKPZSF4Rfw0lRbDMHYHga7dameVHlWE6SOEPzWyhqR6iM39pPFqiac8gapcW
A0DMSPyQMPM/UN87u65icvaELMCgaDts44mqqQRjVkdASe5Aqi1SDz4I59TJdK8U
oAKIIE4dj6jqYxxvD2pnSj/fg1bzFd8VWMPDe+vPneVQfpkaTToW3UDyKRVmra2w
4ONDGUl+GSipTz/4mvtBSc0ni7D3zh/XodlLCDsoHf9rqwP0nxOvDkAN7eVcDNlC
sNx6KtMKOqmpbKnDXOh+yDeTdS4LJibnLKVZoDQ3cREMlR7t2qDgzuKOv4K0MXhj
vhiTaMXdy/CsP2P+FJ9wUaUsR3JjembcGsCMqOBVRjZ6Lq/xTqJb21Ufa8BVAwQV
NyX1etowJlqNyeqy5ATZmPwSkvSOhdMsmqIDcfdp4KJ6lW5mzbkFsGuHBSR3s5h8
B6VOVJ2c3+tjecItCLuPBNQ1yP5/CdeaI/GU6E+oGjsM1pwEccyOtsssjja/dSow
XELU0Bt9l4YAdM+r1bIiSfnezxGTRrnJs91I+LKIRT9u+b8FwlWMqPJBhmlszO99
07YL746AeJHblYwRr5dRbAg3TSqRtPSR/0OnPXIMoOoGk3qjwmOCITk151V6S40R
0XuozxSj1kO7BLu7n/6LM99Bi2SMSZ5hQc//I//GcIjn4zqYx7szDHJCxVHIUzBf
dAM3iD+TVR9EXQhs9nHjnddZ1N93s35ZSzOSB6tHzDRcvOXV1izrT5+Q4M8+R5Lt
BwJL+zcOS8gJO1BQkfVmwbgH6tVtFLgTWY7cjzJAOleoe3NzUFTkCBoaRai7ILSp
j8kkSpj7un4kn2I2mlkUt2X7Hl27oLxjfI57QOMWIHQOGqyZjKC/KpnTneqjgUFJ
/nxDkPt6nhnZ8Kvp1NB6yNfU8DSD+XwAAWj08BDQj/sXJk/4OjLQew2NvjAKD/70
P4cPFD47XNPbcXLdZMGQA0W1u27UlRQfCHXVo5rlFGKLvHdENN6CHIIrqQZV5PYo
rLTL6d8zh2bwJBI5EbmAULoIJNNVExo94a31MTFVagajWUJ2EuqTBz/bWtamDaq2
BVRAXI1h8985StWHzuhiu09q/DN9UqFfnDLd0ZtopIIj5ufgwlBG0Gm+NAdKO0y+
8es+8PFeZO363Map6CsCld01sA/6sbgrjYG3ss7MsF3uD21QfLqoQjhDRWrzGndm
CgysT25wbfEoU/V7YWTXyP+62jz+U8HrorPNVE5IdM6+66rqhTpj7DawGCZo8zqO
awSZdOVkJbrj6iUAveObNq4YYQzJOV/4T/QBWSqFtkzdu0IhJ8NIGKa+viTewHe1
/F3ZnIJwZ0Il2GlC3oMo3DITt+a7Ih0rTI7XyY6mci1ds0SsTmZu1Hv+RNrUy1Ev
nIspqu9wH2Ug/hq7UyO/0lSMZEGtbYj2tnV4b+3zOHHvbC49bNfr8RrlUP0pQXBs
`protect END_PROTECTED
