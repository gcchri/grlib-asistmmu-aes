`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IOTF8M3BQatqAh73Dp/cmuJPrfIPATAHnPBk4UIX2c3AQfu5EfZ+il7Aa7IhDD/c
th9h1zdrdbPiWocTBy+71jzI/W0HDLus302VzgNFyd1HBpG91VQ6uO8U7klgmJv1
QLfbNa0hJWBmV4xrdUQ9qtUpupDu9fbFyfjCh9V/07noY/cirhE4VLFSdWXS+ADW
gcaxQBDWwLuOXO8qyNJ+y32xOWLfDziX21bYPMDQ7TpRpAd+wscYkXcE8rT25eJE
OaKvocsLAyVo3ss2eTJdXhzxiW/us21IYk8DDMtQMkqMLGc1j4gbpCFfbpcL8k1o
eHHIctX2mKzkpNGF0TTlC6Eg8H+bvQzhJK4fjn9HRPk4Kmyr/z6rW0Psrwle407i
me+5REPCRIlc5ReLy/d7+5oJBC4fezyQHO7dIS/XjvmSDZvC9uw4vLAMt4JVtuA7
`protect END_PROTECTED
