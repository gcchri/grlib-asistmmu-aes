`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zV81G4Ufagj5lzPWh4xhJ6MIf3XJpfqdkd+5nzdQQwhxTuXs8+agnpfg24UwKFTj
TBld0yjc/O0fFtO8TevT+B04avca30PlPYegvg5E1/HCzTnoX6E19Wo39t+WolO8
Qq4vbJvroW4BBfwdQUos2ScqKjXb9iJ/nVUpFOcW+O3apR7iAc6I1B5UHyuNbdZ4
xwYf5vlLxL0uWB1kBk94k+Qieyp3MsqdTJt3YPHaCc4xKiUFoPNilc6wHTcKdVP7
+Fpu76SneOjDP3q1/YIZgBAFlOhSqi0SOwqyKvKxEUuh6Trxlg1kFWuvreWggWv6
O1rZRgZvLJm5FyWB6rL4mbmYgPWM2aXqNs7fumD4RW6Q93Z/pDvVkTcJYlezZQof
J+6kUu4HGeIGIMV4OMddjthkrdIFmyfvIc9IlyIRm8Djcr7mZS/nES4JJwMbr7/a
qiQh9rvRuyGbtXMWe0TlPSTDQyyIyeLXMqzkz7o/NkVB4afA9RUIBynk8F/pe2rE
Q61YL/RyZAlRZ01kNMjS5DkXus+Usf6vg+TCUCLDx1Ydm8yKw0lwlQb/Daqlg4+2
5Q9gd+DCc2phJJJQKrw+4jk3X+2XyQXz7UnwDM9dOa6h5XNF1AmKcP/FexBDMbFr
H0Jpf2V8gCtzLB753ZcUd+nIqvfki+YpLEGVFy9COFN8taxlGxsSyygs5P3pGqn1
LrLhP3AmfyXryJiw25t0/cHuMXpI915vF11Qw1wV1vDPrIEVmYUOashXSIIhvu4R
UijiyPhK/xlbD8bFHxWMKQ5ipWcUT2vgfOEqMqUxKvlJh/KhACDb4glSBCRq+3qy
dsLNKlE4FbYqLqRUpuhVyRLk3qGvVich0yGR4GnlI5MT2lFOupVnj1Awj4Kif2Fp
I2bnAtIviAjX/n4X326aqVaaoyWOfnXKV9FrVJcWf39e62OjLPFti8vhDtgY5cd8
6tydAbOCzP9zkCa/RrrPU9Ll8UGw+aryjSB7q5bOR4XdclzbTfjbiVUESIGCuw39
NksVjP6o/dT0kkIBIsIpYpmKICbqdpGPQuHCw7wmnigp23wwjWOQnaZFSX1mly7n
XiiT+zMpIF7ISO4uVusIEql+tJYJ0ekwMsgWXiJdVF6aMkSe07DMLXkS0SSfuuDn
QKJOtPV2cuPWhi4PXonPI5FmoJYiTuT3plOZ4LSmJkwZ8RlDBsnJ/5OA5Fy+GAxj
qZzHjUv0F63WluF0N+fNmascSuvqgMvbFtmuWzB60ZvJZCjLUk+Rbs7a0x8Ic2tL
Pw8Z2AhotgHPWuWetcNLPPHW4WbxNG7cXeZBigawZQBpuinry8qGeYUqsJq783or
DGjbZqOy1EUypZ1RQ3AUMOk/pzWn8gecCFKqKbTLs0ELUpyX0wEF9TtHvR54KB//
eDy9iF5b7aKcUfiQYx1pKktplHbPQAgSFiZxtwmlKMn2W5PLDFO5JItheOmKoiwW
An5kY19o5TdW1Nf6VFOCFwW7REhnUROY8yVwfGdtw2ym/OT8Zy3WA33zFusgJoA5
BEU0UpFy3+QdWk7SgcUkfLBzL9sge6DNix37vyhri+zkL33i7E68Qo6pvFrQzDAZ
W83fvDwEuL9gZ9JHGNJmeLesGTpAYnPNaxNWi+eX38czAjOrPwm0BHg+00jkQHpb
xiKe1odySaA3FUTtktFGSU7+eKrfZxeBTkteqwD+S6FpeHqS8C5guS76WMnlBkY+
bn/PyPbsS9nb7Eo20gpub/8c6SfzmZZ30+67gmwU47+dXSeh/bYyObvQwAIn7IuF
N3HKrR1PNLmLQiOKlMG5KTRSo8eDquRD5byHLZBSncrMoQvvj7VXPeIw4QWenYjB
D7otRfP45trfrKdehHEuiaY5J+HkNJV80PxvhfC/6/LHq1jVarjiqKlrBaLLS/IX
P1wFQx/Yz/d7qlTBiqU6wpODxcbpBPdnwhPVe+oLnFU1HB8vmCQP3OAA8WGF7BJ9
FVqyNvH1t31MukTRjodjbAMkEFLA05SaTcaFbXepuJXC1JZhfMKIC2CMV34KCFjk
t3u7p3VaxzKR78o8yb0PvTy1Vy4PADI0yCAvAkEqKNEa8I99dR+PHD2FutPKqm3T
Qxnw6BKAwSbl6pBTZYAI7UyaRLBwISeq2ZT9rd3zZLMtJCIQXcwIZ4BGAtAgFOuh
qLHWxtQTGmXuh3s5AF8UPqZrArE3Xf3p2wCGoJFNlr3KxMXxhTsuSBJ8Z+fPX6gp
a4Ke5BnEinHb0eHU01xNn26q2ymIJU5isVfUJadBofXDHBG2xiDplu9RBD2WjV1+
dKcu8qCsT/Av4+NXZN3AThrlg39YMRBMqVOc0uu4VhT2+5tT2XYE22Yswf6FoFgZ
iwAxCg+5YKvcioxYNjkisZk0MkZA3r1POiDTStkOf+vdVsKljaGCleTD9VZPgFyL
k45EObei/paFJ441VxZPN1SGkUCRb2w6S4pg7Hn1ZyIPOL+1EBOS2Bsqsw7r1S0z
89U7Z99WyhwOKNS1tTGyYTaB76N2izJbTx0UNF0vG8y3/YGq3Yf1uTnh5H91anca
htfOgmQXGL5TcFJORkAzikG9cWzkBwiQcm1nInnl4PHyrkvOkZ3ypq+bEsXgRVjQ
1Omm2E7H8nB0IKTtHbPxjx2kB2GSuAVyUUFZd0BAq/qOKlPI9ZtNQyrhQjkzXaZG
CflL5R7nG7DzEoEXmodHjn/g4dfPKPk0UNIXFcoDEzYhLcVGLKNJg8AuTiBdBNGH
SpdVfGsWeaUzpmaQR81aGAzwgEDg8teh2ffCWVmosvpIBB1TuLietTCgBx6IBpAL
122B+OpieVAt/RO+9UPSJ+dPtHe60BmexVEEq5KCdKR0Sri8SM6NsPozAlwNIv0I
qsZhSIF6Q1uHfF0/SNw9Kum26Y3s1zBAfjA0LsE1cQUAMcO3cGxY3Ag5rXLPHOaV
zwiEwg4pqK25BU6GTyOZNhPg4cHc7yQ/kAAxM9JWGmhcvyqoQbZ/HB41YonsF5mO
IQUG/CHzdlTPuPj/k6Djgd7StodyvN4LJ3Hmsj1xQWdxrqgrQ1ioDsKqxFHSucjb
8EcAdhGUz+15i1JCGinHKUS+DTz5hS+BchMgHjchaF7I4QTVzKAiqjM7u97Kpxo3
3/+3Kf9rY9YY0XW8sVdqOtCJfK3Do9xCVp+9VsX+IBr5KRTeTpMRXmKdS6ndns1z
mbx3yr+9bFmW1U1/wMsFfDVGu/6LcZ5Y7ac5Gcok9UgMTolAYuOjF9k4sRVHHZOR
8eIcgx/62LFJLxglNQ47XSeM8nKDazk+cgEPHXn48k3vHL39rivxgxlJln9I7FuS
P8IKsk+4EoCdxHOYY8zII6bzNpny9IkLrgXnKmNKg0vR8NtOQ52MV4EU62HEdJHr
KTldiaIcLXtDD51cFal4nskU4lsgLCbyR000SLr3FVMD1crKulmMm20rlQBsvrJ4
Mm3FCcX+KIXvsnSmK0zhlyD3/yBBfQZXL/9W6QBL4kbAgU5M3w3mnNmg32BXnQxE
e4o0e6UzWK3OPhRBMlGx/ry3idp6IwwHVEQmOCRzRCiXFssb5bM1m5nwAObSaRKi
qsgFe/VDiAhQY9sHHZJFtlPaKMv3tgmgvUZf2NG3k90OzudI+TqWniu3rvUI63Vo
KgnrNfdVoTQrjHXPlEUbgeHC7IMGVIDL6VdokzuLE6SHh9I4s/jZ8SdluD3vFo4w
tk/tNT+HXrOJVZjAtu3pM6mVjEv3m9KGSHFnOOY4X0YMAtAgwScj3Mwt60WtbDhS
ARvcN/44iaEYgxR6QlF876SZnOKrwRo8UzAba9IaoIERWlcasxSMPAID7zT7cHIy
UkoOnUlu2TF6FMEC/obK7RSCYH71lWY7pz6bNttpaHFsbLVDpJ0Xgdem0EY0LSni
UMHUooKU9XHUV74NB1aEKUypGuV7ggVnE3CfXGfmnGRgTjKn8p3ALv6QEb4BP02q
CsZQaFWmBCEe9Wq5qApl7cVBpnr2xi7mCfCZ2XK98o9STKQh0thSKaD2yTGmOEdW
u1aKJcxoLKJsw5HkmzPIzdEQ+hG57795bd3gZTe2Z5E/1rWfev4bsRCLOxOmMjTi
gSd72eik2myjpGskT5lG5rTPyllrIoC7sOivgTbAC+/WYg0dbIJCV0de+MwBjCQv
vyC++XdcP2nfiuRoflUTn/1cocy9ksXlmZv187XFtd9Rum2rDgTRIyAVe3tzWNrd
82PwMuSUDnY8e938Rn/1Yp/vswX8KLig5HPHJw1+HmDqRI6RtA60KRvrE/BlCTb7
/uzDW+c+kN5Ol/SI7RmeoZxkoBC7IDzxeVYp406RhZuYpqu8e8+MInusSScMSK57
klj9Z4NgL3oNEmufSh1N+5ms7KQZJ0JrF9Bpn3zOsf0vv+zchoXYnLcMNPa17qG6
0Hk3rB0pJhJDYr92MsFbzXUGrBuQWQCLx2TscJr4YSmrrv8/CnGc8kge1x6lYD6D
YTDUDA+tuSjUd6ZA7p7wC2LIHoNwCOu7eOo2lBu0+XBSjAzvarno6vhqvKf9zHnH
xAEvnM9FG6TXM1C9sn90Cv1ZSFkn+3gcs0fp7+cie6VB2lDP5zsLltW3xt5DOhPk
3mo9W1+PJ5ny4c7DzqoDaPtWq9GzwftIax2D/AWVBUn46wxWOYYgTzbE4XzMe3u9
5kH0Nh3nJE5ig6IUiXJU516slsw1cNlqosWQglQJkunemZDF/av0PflqzSp1Uu0A
T5GEpGTkbyvmPkSBpduffW0Wx8yvR7ilPyNDARaQ0bIyWJYcAj5AVUwrIRGKTvH2
ctdmTvgjfC/ye79Kbd/EtgAUjUs+iVqR+d4FMaTHQKBOkmCbgjL4JTurkCqEsXMH
vXeL8zhADiCx6YbdFv3dL25L89V9fhGE+XDm0uio02Uz0YJGvUX2dql61I2HPa67
/njO6zOJQZXfG5QB9fwnIVmBTChBDKbuleY4GQ56FJXxnCdZ7hx6YRpU+GjdMCEB
pRp1wzrw2yfl2lS0cJAFvo9ramSys6kPIMmy+yqGod0Y7DHNNznRudiH1G1KD8jE
+2ZbuDeEHDGibNqbW0+oImva0tXYOdT5C5p+hDYc8ue85l9TQ9CiDICW8n2S+OgW
UttG6MDR6iDqACnHUvaQpUg7sQpnXevRN1MGD4iXBkN9kSY1be+TqfCZBWkddbCC
2Dz6ElcZf8SKu+r6jy9NE67QB06/PthsRC4G2dbYrXYiY1uxjodq3bwXMf0cB+zT
piEEINz8fWT4jrszUefbUcAGNOb1EbT4CDy0HeHQmUdDLCwp+vyXW4+8bKtu+tCd
pucMl9lykVbi2YvvlwvhFgIR+XL24c2eqG9bjNJb2gYXHC2rCKTZVP+/mhvbOD7+
ktxI/eO41gQ5If8YJ/2ZZxCeBg34om+SO+X4LINFhkEQUI+6znoCjcIrSUI3GFh0
6GjMyX9TQjKNNrrStj3lVZs4o4ojzncnDUvZw1mhyBH7rL3ZDrqRyH1gEkYaCTbK
kjw1NDgppg4Tje1WEmQHe7pPrhPJkk7uuAlAQdiUoIoRPDVuQTkfOIeDOLxAkgYn
iAuqLIjk0cXK+DiKI7hfpoM3ubVGJ32PqsckHvKr8pyg+W8WkuSURcm49FFpBu92
dABjVmIo7cjlq55OL3SnGsdQv5cCkUNGfXEe6YFuf9g3pkBJU9rjNtv/Vo1P/aWc
aaE3x16cW5GP4rqpjR3eTsMVJfAYh3Sb4QFnelYWpXDvWoyzZbmKvJDja8zQZ7qV
nZX2KkoNNh9j+WsTyUxSkk06EL1CvFVSbXoA6Uqp1o9krU3dE+UGy8PRayJChr+V
9dO4D+ZLIWlXfHByB+KxHv6wqfSwigTjaGp1AlxQkOjfhrtD164pe5klIK1xsNzK
0ANbPMv/xMGVHlZFC8cgQFP00GZVg28C3f5Nbt/jT1ete+sUgCEwG/Z3FVcBI262
GXNuWTsJ692xlgx0tfFGXSQPOz6tYW5qFercNWpUQc+Vpocy0zVxsoUBQFdgHphH
PBd67w2P8wkm4RLeJPJHW6EAL33MSaJ3AnNLyawXQqnHlblFS4bUcKJ8ZJLQrHd3
tnJuzrDVpzd/hgmUVJC4RTpTOL0Dav5b/t2PVml/XK5gn1z/BLrIoqPxnmLoJw8Q
Oz2DIZw6R2aTD9Yv8cVXTsBBwU33NmJS5zZhjVkumkeafDlQj2SLuieGeEyRcJI5
OqbRr1lntWqJ8WfLaXOdgDzN2zVTqdHjchvq3z+j8cYjXQxXEEBDEjj1pV1VNsKs
SUEcYANWWlP34mpep4ldNEPsElLrF+VEPkuIQQ4R6NHRv/5ZUc0OBHF9gCJ3mbNU
Hb61RzP4J2yflGAxxV6TQc7D5QJO3/5SyaKD3pXoJ2/WpCN74MMIJQhZA2D0/574
sOwW0CeQcS+eNgXXBwXS2HkIbwbw67YNR/NHo1mgAvVwr+aQcbgOBVfwKaGWGieV
dxY0aG0Lgpl6kNUbHfZED08Yj0esQt8jmrCoqeE8F/ovinifv0VSoW0ISq9Ebtx/
z9QUeyWP7trNN4nYi6hj6YcQOsyg1pvDjj47IOykV2U1GkZ/F6EuBQXU9+ioqaZc
NKSvgKTjuacXRlvyq+cS2dtwgY2T+wE+6ReeHfgdvP746Kb9Wtns/gygmmq3W78l
0TVoGfpZrLmaDd5mvLj4eRMW3vHAG7dG9kiszsZX8BqfJDdyIJIYQIgpHGGJzfRC
CqRXO9ge35xv4fqkOHELngqoV0XjJob/ZUfnu4f8m/CtBXL9deSlq5Y5zeBRZV9L
etQm9dBNVI3YRQty+r6XMhL+OUPGIsPQNoFV+DaHGqs6dPXw6+JADsykAKjwFtaT
Wyx0K6U8ZxPzFOWwK0fdSiJTYsauY00wiaBiIqG5fmoOIRqxKXfPvTIq3BmBkwZQ
yEeN2mGhCashTKlhWT1Z0ZBWI7RGoaUhFhgYk9UTqln28DoAuzmz+YXkh38J+gtZ
qft+j4r0gGir5Qq/EAqKGPERvrDbNZaMtTj1KP1Z+3IFzeHpaTs+RET7oQQ7sL9Y
AjDOie9slT6BoxqpIYGeFU9psk0CNTjV5rkuIFT2lzV+INxfYhZF9nu1MsnJu8Dn
hvxlWMPgswp3hX12Ahml41XswLC9JJNH3tOLqGKXIlD/dm/8SQ6MQ/V+btYgm3v+
yjbZMTWpViyid9KEf0XFlAjvsO2jqEQ7PtqWso8x/T4ha/rbC+l1S6LZXo8D/XYT
I/X5/P1lFZ/PFZuKqdtrLe7cWZpkPKsShTEerixPTjAE5Qb/w8UvnD/OlSfckh2N
Gl32+pzgnbu67jFoJoQ7QhEeE7N+h0I02Bb6xdlk/Ssz35K81XdUwYDLqA6iEbFm
5PL7PMtMHKbPhaAldD7ii9TIdN2Se686wkf+EaMiIUVWI1cvjbktvPocsDhlnPRD
ShHb5KCv8POlZEKZaAHV6iIo3eGWypnuAVhA8r0du3KhQdkilGonn3bX1KPGcsPJ
E95OEdk119pve3N6T4OjxSCDg/8slTQyH4gK86/garCaQ2rB3kohY80cjY87bLDu
ePJsrFZYI7taFNmjHbdyS7HxGOU+Md6g8nqZIdOaS209BVXkgksVoxfvTV86kvkP
h84iRhyA0HqZgXil1ny7OqVSzP7+oCY6yJ2VmA0ZCKlD/SVHqP/sW5yfDV2ljLF3
yoM0X9cRVfv9Wk24ztdkobxDP8/xeUg3QQ0e7dGtn+bXU6mgucYbrppvPryH+xjG
x7yTeXUbpMd23dmSenGIppD7BrnuGfJxTJMzJ0eyM8OXSg/8Z/HMgu0UIXCLbYeX
HQS6wOkHIf4qJ3bf8CjvA6pFEDoZhpVaTVDsaMCbybNGQ3uAg6hhNAGPrfz/QpeB
0ufjNeYDSRWOqIltaDfzbdzD7Vjp45jX6uLgzaxPWLG+adMrItv5005UVROdOAa5
5VHd38aVI7p4f9dQ7BsR2uAA47NPlQASLCxRPS5YzzlWQJbot6jxXRQlv5fcQgZv
FQpG2hZkurvpAayUt0QX5rJFK43ankCmvjhDl1y7QlocFJaWSvxVJrMuHhd/XZoL
8Ht9kB6mMthcrTeD7HxHuDOQjkvYUc2jtHuUbsej5nVUlhNrQa9wk5V3rczTrfKP
JXIKwgZANWTKlLMSTQ7K7fVb4dJjQBNIkn+yEmTmZmKiXhoQolJaGcM0dvIBS6r2
XXrGX1zsoYgSNp/Lzw1uaQ/gQ8mfef6wMIJ+yTNxsGa6r1iVyW+OHsJJlF9bYyeB
Te63l07x8hEia84pPPAepJltySnRSQMRRh8zOJO3OtNft4pP8icu5NBH4iZcoloU
sI4aeteUjMIEAj2FRFh1D5mpEWvbAxJcTxbw7lMQnn5KNxRGVX2tlBm/4dr1Yqlh
crHunDUvjEyLn5UhCINTEmwwJdt+D34Rct+I403REs7ucMb6malJqySSfrJ0RLrP
kHkr7baT1XY88YVfOkDq09hMoLp+Y7yzZDTxSlnIsW2sfSW06BT9APnnzS5sLEyu
1Hk9ML/D8xz7+51nHdz0S48EZmZ6x6quZTtqE8QHyUfrB8IJl7OQLftwLjc+nyCb
rP4NhuuF5m1KGrbtAk+baJ7WhQReiG/bYzWgskyYxktpsmvoB+E4RYdL+NOpRGB1
eLP98A7XQORUoebwB1LqUHDgIuw6OaIGbQUaCeOxL7rLEugx9e5uLwA8cjEsyZ5r
+1qD2QmKHFi2x9bZMI/4j+QhS/FDeE3Y5HZcSz3kHRI9V7KrsLo2tmdIN++HYhB1
UAgx/JDXGDk1vhHFlk+leVnvEjDYgVW2ZN018qlI66Gdac2AdMLfXde1eBtyG5ZH
M1gisVBIxrVLtPWHE0e3ciIivSED1bKaCNLb/m6K1/yyJQ76tr9irw2JfIUN2KKL
m7bW/9eYFvp4sh2xlA/17QqE0eJly35+119kKo47h+bEvhITHLMwrjOusMseS4i3
Kftl1PvUO2opUZTIpE5md+pFs8TZQe68Y9x0myMzoPXe1m0+bHBK6zZPQSsCYx+3
f1piJfTBVgs1++mKCtwxNSoMGdTt1zIzKafeSkS4monsaPjOKSQy1w7cQWKZLtul
INz4wckSGznVN4jux4ryxkozThT/k99MbikL/qnZFzi5wtboaidwJlBIDtPdk/pj
h3g9PC4OXoR/lQPTaAslsykzs0y391+PmIvhNGbhN0VCnAEYWWI+uL3mxEOCsu4E
+H0OBoZK2ec20jFu9C3o1xujjU0ATohgID/+KvjEHanQRdzBoBa9iRUSq26FxwPU
zQd0SVsnUv/Snzjh1e0cUCwRyPrjKCtLlHnjS/QpCEjATDZLSdlfXVR9FgWgM7r/
zg82vN3+84iUb1lF+sko/N11KLzmkb3ACMOiF8iuacSBS0bGMvt8x+4wiCwkEmC9
3D5+lX9hxYWbD5LTssCqqhy/RwnzUZfVIsse3aLpTedpzukov4VpG1fWqO0RwD3A
TuWT+98z+wTNNu8r7DhDMI6S0BCMRrEn+hYI7yH6UlfkAvsYRbSq3edW7jlSPTkH
aO8MqFRaj0DB/eOQef6a/BF1JTBu5PKEPqCfzarjKfxpGHF4SXWyZ8o0oSJgW8Ea
cuzAkhSSw1dwIlWgzK3UYetitUg66VOa06LAgElpg9O3FUTav+gavYgyi/2b2V6C
LyfGC7Ls6NJpJuuChDT7dlUl5B93zjfpORVTihK1+wEnTFHcLCg3qEMXw9FE7p2r
22izEmY793PxrFc0GF6fiZXqBqGb+Xaq1F/55wpMu25AzVlR0qFT4piEh0D97B5B
C88qSP7YBg6fR8VobbPIxuKj/kjDxb8y3tCBo3qWjhp7+uh6r4SHFBBJuHSjfIsG
NJ4gFMlaKIY48j2FXJ2UCl2P6UprOBMTq06lTeNjJF6whJ8OEPMDZYvo+hNmpEzC
giP3cOwmyujBy3vhspcJUiELdsVT5aPWpx3ywbGajWIxbZwUNQw79/drHvy4ur65
sCzBUcE9ZLcUxcK0FiSq5y7q9tcaDcuCPKfTa8cJ9k/MCnmjAhUK62toKClfaGtI
XzsVsPr0CI8Yzj6MVwTlojMRqVDfqroxRDMUHnfrEJa3UZ+/K1rBl6rAXNP7oYVk
N79uK5Zp6dAxqeSjjap4aDjg5tp/4nayawYAREIxoPp6Xpy55NJCfTuuZv992efD
1yXqDThsy3Z43ixSWL9Z1Ha4cp7IOvY+7cwgRgesngspy9lza03tNexVma5oR3VL
1gJ+uPoMFM/L+hJeXoiclknxESjhBRiv9UMk05RbH2hhJB9slA/i0D0ID2zkEwcA
B3qjWaw4hGmGJ5AmNXhKv4aXehNeZvF+lTXhWi8SPie9DKXbLOlY8KBIyNYkhcVS
f+J9ESVytDtswRRee8AFQZo9EKYL7qyhLSVKjt6/XFQdnaDg6hRe1WEiEtjKNtZQ
kkCPwxi/itgLo3cgFDNH4IlxbC22ELr5CHw4Qvl/kfD7sPUyfbCHhFNaddsBxuoq
p12ghTGAN1m2y7/GRvqOY277NWZKzAwxnU3EaL0cr90K+nc7gxsVJma9OC+WwpWr
XMt1icfwgQOyYRHST151+4GgwRsQvhU6IWPFTB15rvSfrafQg9WpULSNeFlZ9i1o
Lar5yNxZZ/LEUcxuQ7z5zC9D6jkF0OLnhNGlJCIspW5Q3fRL5atRpvoxpZ7bOB2e
j0GepzVcDCJbhXctN2wY+J37PxMMu0CQDvJmg9l5ndYI8KBaoKolcVVQvL0kXT8V
1WTZK66JnLIt9O2cozS5FOD4KaiVvKXd0IcyczZCnp6jBRx2KPPRonHo59moplkt
Xs/tpayUuinxheDCqhSLSW5LM3UpGxJ3EiJHa3JVcHUV2wzWeUOBcj1us8BZeECs
kMABt8Gf8+6WkJ8Xee6/06FvmlImeqkk1SGsCzjrGTUijzqIedApx+jt8tLZNMK1
st/zClNnWArBvpvL0dh8EZyGHY6yzl0X2RXEF9Rcmu8LNcSin3ZQ0rGQmg2hY/zo
rMSrt3G5sI7QwGxjV8uQSTnFPvUx/bXjlbLauvdCEcBogIwb6M7CggQXXmEMbEy7
4rnt9qftPa8zxN4RGPfMPS4R1mNflWHDtCp09s1/1JAq3WwsvZ1i7S5HZg0vF4NF
Z1c3Xai1JW6uDIJixNO0PP+Kdbc+eMGM/k1j9KZhAeG7SYDMrYe+UJKldHOt1w75
FZQZGIOVojFPKJA2StDLT/mtz4uZIZYQIpQ3yBAwHSaPp+kx/aL3GQpOhnW01SNP
PhNi6hJ07oaVDBrF2qECi+KGu56Dnoi3jNeUaNLApOgA89RRTiiKtMGSGNYjEUL0
51K75aqCKs95Ys6er8rWa0Eq53EA80Bn9Z8sYb6PVCEjzuWHhotlnTE4HUxyi4RW
QcF5vR0rlRPzO2A0qdlr9zwgbLS/UVAsvATzhXOxb3mUuSuHznkafXDtgcrY6E/W
eCaQph4r1rqYdMTdaF28Bf3JlPGNayAcYdw2ZktG3vEoitMB85+oRqsQVoaJ9ld+
3Y/PqoVBF7sfOpRUTYCq4Sn6bLsSbMLWNg9G10YmVlFh9PScl64RBoVtBD7V2Ii2
JBGgaW1DIu7ZYC4AG39UQHm9vNAvE6I5hqUtowkFOTHRQoHDDIyGOZFpp58kqz/r
7UOqGhY+C86sPzs/Q8NvaKs/CQfih1H36joVHKBZ7VDQSa7nFsrAljVXKJaqyh2C
h+PogBGZvvX/AwSy8NUu6CyAM/pSJcOtU/u9UvpNTj+/upN4fbkp1WjwqzOrrK15
EQ8RMt6wiqgQOkL8AweQ1e2MmOwJSMq6OlRt/4qQScxjaR5fKU+wUwHAvpD+8uLf
YUqCEQcQzptXyPz1F/B8mdSfqAMRw54TMLQQR7fv/z22fD98eXvjCg8kWwElkZzB
MuJZYyxEeUeDtl1ue9ueJg0E1gRjjp0kMht1AM1EsYUJq1+sCY+NJc6erDa9eBxD
LLsW4CkdCCGXE9OLfcw+jBTPu3xs9lH+LqtlfvYHJAv6P4PXOxl+JZ8wBe8e5I2m
UpUlgUADYqrgsImrznckb7fP1njeJSwwb8wOjj5YMdOS73q6Wy+qoS0zNyIG++3g
Aipbd0KRVbsbklS9iQc2Wqk0JvlMFd7mtfNNqR19LA1bQHF4bLy9p/Yazt2OyRhx
vP3DTUifxlVoVpahSzyER9i35Cxupp+z8Y3qn6BJr9fsRVmC/Yj85k1wiM3WxQuH
v2RD3yaKYTLio5EeTCufu22l5amrMWn0K4LFjG7nUU2vuevDaJbv2s8zH7skz/7n
gyC8DbSMxou5MKpyhnshnYqd8MRi6U3BmACGHu20mmgGMpzXGLUGvG8kKqVv6hYk
BneNrV346QOWDKEJkO713ZETH+9lua3uKHJBD1sHLQ8QZusqHJEkhwUbBVaM8V9V
MDaulbjFJFAHBnQ9zzqMzHYOg4HCMIFKTML1aMKGm2mlMn0bysrrfgJhAA5HYLn2
ygQIQL4axK9uP0ted+FH0dBxYiQVW2mmaxraUGLdnJ5PLie7s+oa8qYDyQiGlW9W
K088/JMPIxG8ebL4YuB0xe+RxRxs/+zQV7RGQStVjKyCBqS/l7YLLCvutGT3JLfA
z5chkfhh9R1X6ZcFE9S2iLz7VWSJA9ELb1GfCC7cjK1sm2iza5A0rHCB5d9be5ck
6RkujdyQdHBXXfS/79Nd+ehscB6dEv6zKra8/Nm35ZlkmpOdHppGM1Iz9uzieYxK
CFx4Otp1OzRLLgmh9Tv/5jRoiPCe2dNhN/M4Sqehv8QHLlJNkm/2PNh5rcZbIJy5
PPZoa6Oxq0tuODrAh/pFMwdSRRTSe9nmOLHYe40qZ5NNcnI+ZvdR+TJS2COioXEH
8LgwAuqUH4yOfxnmvlPWMB24sM6Bf+2IzyLNyznQ0lZS4r52ufvoT0FBmmJ+3TbD
NC+MX75OnVS9dJkcMasj44aGMhvtaHNdqLXrE82HQjvsOr7dkWzTMtwgn9xWkWRj
kFMvCn5TM8jFz1zA9qphKceK1800+n5YfG1hNgCCbGtluSbhcWVnolERh+pcheb9
TS83bfedIAaTSXFQRiGH2x4sPZ/gUDUVrwNDGxDMnkqxGWPOWVKzHYKQviuAr6Rj
oA7x6lmh1GdwUzXAwG1CONKE2tWIkGOi7HYYQRIbQp2pcJM11M5c4X4EAqvX+kW4
wMGloiymcK9K8HPRPetTd1VBBbqMyiyKcbxbdTb+XgXQWDFBe7eeP5KCSYYQW+DW
I4pxV+KJ6hLwPgZcvKD+ojpCIaFYDtkR7nmXX7CITk2i4iSaoe0jYjaIYg3aSDSM
OyRiustasqAFVjQALnakxM0Qb2n1NPsyVB7tFTFFZzoL1wWUDV7l//XxlsnwiZza
Trn1PJRtz9tNiQXwmtJzUz1xEJQKAeJN7AaXiPXDMdPwYhS/pJ+tx+kyDDjmdFGr
Z2+TkVprIOhuIfsocPRPsI7+K1okhaSJEAxoZwzRZmMwHXYEMaBiFCswmEeiCUiU
2efOst+n/doa12XbrE7/ULbbKSu99j1y3UkvecoACF5RK1sesr2g+Q1h5o0EZ601
oi1JyWXxzQdqlmHaLWpaOcarwGUdkHqPPm/zflADrTdQKFCWyxUtC/qE/ao5Ipx5
bd40cD+xT+blP1Tu1GWpihTJfaCbb+xrjXcS9d3ysxK2jPJ5vJu9Mtzgo6Gu0yX7
L15kFANuFQ7W688Y49ImH8auOfO2IfhkYyKk65OASc9h75PIDaTCb70j2rUU/8VU
YoNhpg5NaynOwT1skljonVgH9dj9rJR9wV6Eu37zoUOPVweTFivlRvrUFpmuNiU/
ii22zqaoZUhqHnXS6pcee0eM1tQ+6fWjBixFJl55pH6nu0NdS2nlfYzNe51jiLQs
r64f1xotyYJcEwWqPsJzj4jyY5dpgd9eWRE17ovqRvJbSu1GsaQzVcq3C+AYDbcC
x5/vVHHGKxQNJKSlPE0S5EWf/Xg6IK9lzTxYNwfy/W8=
`protect END_PROTECTED
