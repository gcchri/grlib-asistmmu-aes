`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qtdcpsCP2NtTbGCs+n44O3VrbJMuM15h13JVoZwijT6rSKlSRLxESrKGpE0lvZ59
zSRk4PSdFM9w8H5i/uFe0V2N/2MrhmmDiK5otMdqMjB+91THFLmu8vmy0/6KYiTZ
IPTaFzePlF8RfRYA20YwFWg5/wgZNqjiZk1wgkatEu/TEgf5FMVaw61kdOblZ+PM
rUx3Gdu2xcDw9pX7R9IqDps8CtD4coTDQnP0Ech0bZmqdOG7Ju6DtV1HB+8y7c2b
jnuxxI7plNbtmFTagFCxzw==
`protect END_PROTECTED
