`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fs6vpzspsvhw8ChHaZt1gszjNOmW1kG0ksqIB/5VBk2OyF2LxCS3wcLbUH1mxzBS
arWB4PmZ+PZblC+fmGadmrlelqGkW7ndD67yG1k6kvz4iiXdM/n0qrVf/vHvHZJ3
JDregeBW9ZIA6ttkoVhrUbLdLK5SDKNR5Ucn4QW2zRt1UETSN+crMBcSFWl5Il4g
XNVlTAaBRLY4LohpepjWujd4JqqQq55cI/iez6DXiFGQVMRLeUw7wMsmB1qgPvWt
CblEqqRtK/XPcbmMz78b7olis3zarvFFTtNDNXZxrFP2H9ohFReo9hBb6m9kG6qC
ZmV4ZH7NsieE17TB/c3SygPx07D86KhVUHufOtznM6u/Z6CLfBagusxJUmpcbQu8
rhck887T4SMTO8cVuXuF84kjbeMJgmEqqsY++P9y+25lECUDddodgPNL7ZsKWpmq
6hdmS7MhmTQMWek41s9U2IRNcS0pVU44vbkFEvZDCKcHKRutvt4J8R8CmAMqeDvH
`protect END_PROTECTED
