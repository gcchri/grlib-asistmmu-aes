`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aWnkKL8XGaOqI+5MxNqgntvkNFBlaJsIgdnVQdKjB9W8QHKY/SsdXQs9O0iCPNeu
h/tqmWUinuWGwhnPuyLI2KMsIdz8BrmhFyp4UzEljRMSS/tSn56ARwOJvsd/zLiZ
BC3aM9VP1Dxh4ed6k1pacJ72kP+o/0tCFJUSdEvrDsJU0TZFINFyJzE1glBQkYaP
xZA3f+2NDXZkDLNx653FB4mk+h97h5AkWKKn6TAqkFqwLm5IgevINnYxKKJ4rzNJ
UcaOXVwIzdC2e+0Rm4gLZkjbTffKxTqrnCPzz+MVU0xLATLNXUMkkoCeYqlvdXzb
viYRR40Az83CeK82Vzcr/kmmqUdxkHj/t1MKmXX0JRWWLj9r25ULR6cOXVc9tG/A
YlBOwNG4WjLP8x1MskDffTT2IpqiaP3q6zs3onxjvEAmo+fDlPQStfwZshbBCO4G
x6fWh9FzkgxXjOmQilXZu4FxjbC7WsrpzBZwsak7EU5ISi5c96lIJuhISrEF542y
ZGD/1TjbkiZCkhnqzVDOO9D12bOx88YWaTMjaIGl5EEheBsyqn/dmowhVli+clt3
qgqwRQuiRXWgtcSwKidNyYqLPxRUTVPyZNjWpL/Uy9SuHlMHpaAIRKNxAE+6o62m
+xmbXiUmlZLtzU0ZA1GGHO1moGBmCyVjuhrcAzk3aIDsS7qnldTgXwHdT2EIaaum
GxATeV9PgmkEXlkiLBQdxpVrucO3bCJkoav2VEDiFiGNV7x5ul9lF2fRQnY8Py04
`protect END_PROTECTED
