`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jEQOfiXomCbB4L8zdVttDP8zaq31OSRLFu+o1z2QYp0RHLHa8NehwkPloY6GDkzC
K7SX3FJY4/eW/4aFwxeL5uSR/1+NT8whSTY0Bpw/K1VX/cbwmnCFDtIlHxiOrANr
QDJJ+pnolpXQtQHeC+1LpXD8+RrLJhfr0EI/No/Uigv/O2eXx4XAOqijT0FaADtH
lJvDI+VsaqXaVIBVYWxmw5jh5Xy3Idjb93bX4NhFQ+3ejB+1zMqfb+qnZI6hiJGW
nxE/2XNQ2xv9AiI2TbNa759AiQcl2QXlPtMxaZpncels50Shc8IeEEWNdlPv8VBN
6eN2/f3HCkk4lDVjyFBp0hjluIUzgGIsi/plG88TKLQFhY0rft2eufHX4MPuDT88
4c+KCLVRV4RNMhcuAUqNGfpj/5UkJRBc0N0jGMdXQAhimHJRBC+j/8Qvo2pq53wB
bcXNo251ZzMHquwlLgadiTh+5dnmJ7YihsugzCU9wUvBm0BqT71tl6T6IOqE31Hb
CERTaP5KVycAhvjSxtTglyAZseQshM5vzU8Ljbdf280fb4t70kCNR8mKEQ0qQliv
d6JYY9pNZ0lVREsOOryU/9mXyo1n+DCnP4HtRoG4UmbAzcqq1Siie6W785PGgC49
yLQSM0mGlUwPGcWERBfytpENn74CWdN49HVJYqPUCTBoTykV+WkgDvSWXBpGx6XV
DRzaTjPjasQyn+fSRV+zn90lAHf+aBnQaTNniNPNORLyj/CqCxCPGEwnJRzZXEy5
AsBpdbbv7Oo8tHxAXsfp8l+gFu3hoYZohL3si7R0tkzA/UZzF2AWplHRCOJiDkOH
yNuGGWDMVuLpf0rJyr+WM+Uu+nLha8pSscN4buAkTmKvGRlQWCA1O6uFdHhMa/q8
uxf3Gaa2jS3sAbb8GEEAigTFAmwYRvcZ+4g+tPOs7312f2oVJra0ixNtGf46/Lll
j1Fo7LgLqNS2SzAqjVYfrz8nMYrMYkf2YIgM3zQcLairAdMtzAdzaDcdZnExqUBJ
sCdd/Dj7TsNMkhCvETPuwkn9m5PA1JErLEE1gjDYGLtNi3Xrosm+OsabvaGIkaT8
r4ggCH5qJNZE0OWaFqzO4G66noO4yQjrq2em3l6QzKP7R5EIjEqAWc0TqRPrJTUM
rxrhMxNWvwiGsWUpVe3gm/ETWbbVTh3+m3HynIvXuGI=
`protect END_PROTECTED
