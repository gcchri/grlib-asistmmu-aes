`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FNSzEe/SW5BQLkTUnNL1mRO5DEQAc2gpzTgu0AChySr6dWf9WzRcbDMyZZItxKLo
f/Oo0mRXs+rnUb4DcnxVJbqxH2Hyg43KIangh9R1UIE+F0W3B/2Jui0ExVejsS+U
bHDJhFcPGdR1p4fI8CLdIsQ8R1N+Tjo5nlXXoxIfLXjADhwCPixPbwztk08ePU9l
fKsvMJ9s8qjlyx2pe+RWcfOiq3KhZj7UEMwZr/d96igLowDCR3hWHET4m6EdAy7d
6VYpFm7eFfsA7Y+i+PMgKuOHvjraUsGGq9kQjKClsu9FBh4TOcLRevEZ+D9Utf3O
Ztu0DepQ641PFb22GXeg3obsiPexaRo8Moir7RjElEADxH4qc5O2lij+5SJg3Wjr
E8zOd6dk1/WonwU/6llUMtAcyWk5kYTLQLYFkTMkxW83qIDSjMCJRCmb2OcNE0ZR
MdZO+TC51BvtWQw4nsmC8wH68CxqzDog7e0rIEKTjajb1yQXUNAH0PQWi7pUdweV
XnlhDFevz8zgprTLwBLfugARqfLP01ZKSb537blEn+yd2xPvQGAo2r/gDRz3nmIk
4dpOibaKYxSZCYKIvd7rYATLWQAJtypLpMI/CY+UTS5DNxdMaZjBkSeiLV0UMQt5
3+QC46KQw691sIhenh2nQIRvrao3ZvhlsK+NChnSTFyz8msPQYuPIr+YV6YXN1sb
gtWyS1KAB4AVL7UXv8Hij1v0HawylqqVbdNRHCzpCLU=
`protect END_PROTECTED
