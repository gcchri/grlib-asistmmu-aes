`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0RAGC+DGwNtmX78BZZbQHNSGld+ngoTs9G8yBtJO7VXEpNKZSGSfJvxDppQkxWPw
nq9Den05a0uz4tm9Hz+mauzyLxIl2Jws/h4kSDRIhxI9apaArDhaOF1uk/UC3EF2
qoAZCJsk1DtNPFxE7Ilka+EjJ+slqosFuB0+6dd/umx0YKiQ7KGm9bSz4qd7kHXx
DvTj4GRxKM9sXItMlmgHwjMtQq+WxDRNtmjBeIkduWBnzY5gSjMoHLaQIirL2tut
SW2KRiEEd0NaYKNwifMX3ZFOoW9trpa2bShiMcOwBc9CIc0dLCnGcwuqj58HpvZX
uleP9CW570DjLuB/UNGCwH47gX+qBoxJyC1Py1kP48mqp52nI542vHCi4RhrIuig
0JtWobjteqQhTmU7yDfDwLVXzqF0nN7RHm3DdZyZhy6xDMbF31REXofLnjT0Yqlt
P22TgDb6c+ki/siwqmE+3AloTRAYowM0aELl53/hbmMzuxftBrKQ79ZWTKUvvbYL
bAdHzMfDAiaV3EYYncS5qq5VQfm+QwJ1Fsy94wEPcr91M+iv7jD6F3GnMH9/Mlj4
3EhS5YwpgKTGkc+F3Z3AP+WmJRb9HagOc5/oENK5ULNPQ/4yL+shY76IkppIWPiS
2GtVohIcNLfpbxtQyg6AQf3xFXKmiG8upeUZi0WcPkoobFB7ESU1S8qdsWPXB4jr
Me5T+GNBCxgvhCcG++T9m8CVIwG9ah4G6+2AjUVBwTDkWVyxFuvbhJEdT3IYl1Q9
VjW+Uolr4K2sEvHnmuf8QkKk5jXHwOAuBJJPxkgefA6Ygmv87nZjRW6NVLpvkgMF
IpEg7njdLD5F+d2S7a0yyVKf6Nr9FeIPDi+aW4Xj66bNZ38KOZDZW0wurxdCAoPr
Gx33e/J+trse2t8uGaz7SnixZWwsbZxJBTyC88rdfrQsmEV1MGlilW6OwipHwen5
3nCt+Su4oAc3lE28fkj8U+GNiogtvQw2NVvYfFHPwjS5t5NudK97O4xxRa3R2YtA
OezS5xmibpri5nMNhItJT+IW5HPRrc+uMLz2CRNQGwKjct+oBbngF9WBDbPfvsee
gRJjSXgFx+8RhtLSS80QsXdVi8uudpDV9Xe+1YquuT2AesKTrR49SJ8wsu7YMask
Tis/gHv88k3D2A2G9FxbKq9oxiLS9sJhWspL8NwFARj2ykq2mzpAoqOLWcZu8uK+
jZgydMSmVWUa5Jb8R8PKHc2fyL4o7dD/8VeyBWCSH6nN9h986DQNkae8qgG+9NQh
l7TID+rWsc0G7zYz+hdhpfBC7YBPeyVShEhPardojoaEBiMcd4fFpagpAK/8Ll4O
IL45+QA0mzBR/4HDK/32fXwR8a4L6SW+fq+TobCMnAubizCytvoGgr9TKwGImSuo
ZoDWDK2SG+pkk3J5fllW/fczsa7wbtSE2yCazNaFbcNYhTdhUcBmzKYqVc4uwW8p
o7hOuHERbcaZehqqNMZZHTM5DkcnwQKFcxCI1SVLHoJkx8lCkoZqhqfPSjg1S4D7
l3Fsx6a28swfxxbImfusArQ/OcZ95YaTRcnFk4ePcXovJV0snWSMLm0uxaLlx5oc
50JPniIDxinJ5J0kB08WVy4EzLNZe0a6QmH8dvWzQ6z3YQSzXHXDOq0ROiA6FKep
iDG4JN3DqJATnKOArki1VnJGzKsBYf34H3hpGX+q8JrUHeAmF3g6BXGIJuWllgYL
L1Dv+mRElq2MjNjyhwLM0hs5Ugs0rCEiOyhWAJSzY9iX3mUEY63nS1rXOVIjMpFN
9hZgc6YHFCRo1WM/n7sO8c1OTw5IUf+uyJ/AqVfq/w1yIugqHQMDWb4FC4nmB1/A
sR7ZwmcfDCQqi12CVBGYY18xah4y1gzXFd4eS0yWfa4qUZBSK2fU3TvFxwnMtkCJ
jaUUqDJ9vaiqMj5S/O5cJa9xt7aEiSulISvNab5/cgcg982nSWQlbOJ1JhSbOLYM
oPIabx4C2zOtPlL1woX7/4liIANDGWJITsf/C8lgIWW5IPq6ASx8ugENK17xKJtk
DgaizrX7Km2//lZsU3Dhz8LtP7cbdIcbeqxb6Gf7bgoDry+w4EFnZ5cKgeb9R0KS
RA6u27lXaSXf7CWegCca67Eqqj/PfKgKr/14F4QqCrAEivMU6HH2EOubPW1sSVxb
`protect END_PROTECTED
