`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CEVZ62fHLMloKx+R4GuEUfjMYs+FEu9C1MrvADV5utBOW/BBVl/nhdjHoLNi/Q6X
R6z5OnLnq10larUY/qC4o8QJ3OGZ7LId2wAseqwmQSlmXRJgzo9VpIYg/5NS7pwK
QHb2a9/ixFxge8lerVHrvnr9fBpmYE1dH6W8cjamkr1yH80nxib63XvuBTE/qLAO
bvK6/E2zKMyC/fIcFcXwt5eJ55C4pDijYC7aV1cuzG//ZNXJp0iEYJNLJkFxZjOm
dKr6N8lyvPZnVMKycQ/aO2Wenb2w2PR88GWWGmR2RKBkilDJZUdeqgkQkGuZiZ7c
RPlqrgPoyhoYiSbiGu9J5w2UsnQvtiq/J39eo/TIvpp5QabmmhLr4gWtTbFgse/4
jH9lJnc3unq2QYABinjih+7PvK+zqJFstDw+zFdftG67v5H8QYJ/vShbx7+N/d+m
zgazjxuecsIK/18AobCYxh0dtDF186LPvKzOrfPxpRI=
`protect END_PROTECTED
