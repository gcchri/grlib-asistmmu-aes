`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fmGsMRA4WcF37/znBTarygHHrF3wSAfkoQuoOvLOUTE/0iHxXLimm7cvU+7E2gAK
BYyhdr6/CFIMwPHQWzd4BjU0FG2bkVcxC5nbcpwcOxkd5kcAnknpvHVQA4zPqv96
UvJ0zrbShcSVIvz+pYjh5k5MWf/7y9dovGF8q0id5XNBCeC/bOer5DhtO6FyHeQO
jfsG1fUXSCdYq9nKV4kWrR7gekgu5BzV/FDvtLZCHNBv2gWt10YS7uKeAWJAmGsg
mfv18sKDZ56zZSGiJO9Bt447ig1+kUis8UnfCIanDCRpf0wV6qFWmjiNnGjCUMkO
w61skgJRL0TmssQJ+j/n1zRnp8nu9ARwve/ogWK3L6gaLMvBxGfmhm+wbR42MG1h
RiTtfnsk8hc7bLpMOl2KH8817nzHzZKU26d92s0+fiNqRfhkZLGedumH4nfpqK5b
V/v6R+GD6mqnwddyNgNDCT4WZMsvm+By4kJvyacRO24IXuUun/62HNZ2CJaaun8h
`protect END_PROTECTED
