`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VSa+ATryrS5zNI5qZrWyDsIWwwVM9/iR2xenDZfNjAiy5jxofF/uA2f76srK4CO0
vbkWy0uWo8bzjf5m8V8ABlwNG5u9bZ4EfASIfNjoUHmCG7ktI6mdYw19ZQ9dSnjx
fjH35PW+kfveAUPRwi6oLldP8m4ypZMAw+tYFzafRmBVRwIJLIzki8axugjpNh8g
hpCLSLcsYwa7AtyNHuknppfdxKB6W2Ewn7kYHdOjyK/NVGPajmzk//Osh1pa4JK+
1i+LHqJglmCmMYH31hNUN8IP5kQumUteffqTjIrNLbZPmNKN+dpz8saDhrRXBArG
iUBlAn0s+X2RMH1ucBD7Zg==
`protect END_PROTECTED
