`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h9aRyCos2zD+/BKqOcgXaVfiwQ07kmN+u7USGHwkAafH12EQ/PX2t0hThWEW+cQ+
eYXJGBM+2Yk+8bOtwbkHs7xa2A13bQQMOeq44MEGtLC7Ap5kZeXHd1pBUzNDGTI0
3KnWH/HJAVpgt/51o4eotHdaQzV3XwWShVySjWWMRvmOO3Z7+srwntmxy631+GXc
uv0u165o4eGEFYbzwsW1ORvDSIPLpVqz+vRtVn94pkTnxtHOMDfTEj5CJRp9VA8V
xwcuVGve6YJBAmklU1/gPjasgoPppegsq1KciBlfJ93+3Bu85CWLGWI/wx+WXI0o
cYabdllJZBrYWvn6tYVI2yL1JiKuqDeU/nqetFRHhgfNSd/6eWaOFGU83fwn//3R
qicqCaWzvvaLvh4InZ8LPpadSS60RjvD45Hnkk2UnXwHVZnegXjfraNXmBNmLKa8
c2WO/jqaYj8ju3R19L0q/6mysKxnTBqm/dH7w4nSWyhtgx1Fj2QFQF1GOl3ymMaV
I6ueNfszUvwP+37I2lVXhWM288yskVDkDsWJ4pirMV8+R5nU6My3QphlG9rDJoMq
yHopzmSSyilCNbcYk8TnaVooImgR1bgnCORk1fD14N7Zq7Qz9Ch3GwYiAaQXlWFd
1b6GDazjtf6ZflOzOwt7M2888A71LOby3vW8t4oYAfTama2Syl5mvUfQRTzu7oLS
sUJAFXc4F9fO0ZkibjkGpi8K/6XvGL6SA73UiO+eggTAa0egIoPNlAjZlRX/HUT0
79CzENdmtTqdQbu/V/TfkivXsMvgGIvXH39DpLwRRPXxhRG8YuINn/S7hGlpWnFH
MCtijOo6LGR3eS7u4wiy4IT1/hsmOX4wsb/RFj5pOgs26DJhUmfeeOHrXI5U1voo
KeH4qaKT9H0F+woaTx8OShLQcWNSnlV1eLp5hX8mFxE3lkdLvxSpwndpOs0anFAO
MzjqcFZ+6NQ2CCl3CnXA3MAy/m6dIevSPR1ZvgVc5YIV4fwxyahSXcMB1DuPsJTv
Ocs0OU3VbpREzVY1PEUBfG1qMKPYeJYFZWddPaJPRnMk+ojb9UbvsLrLNQsdZYl2
6Oma72w8EDMRHhP0/I4Und2MJEnH4LNdEFDVqUHV4kS1T+ecQUyJC1KnTJzror4R
6wPqg4JxsKhSC1geE12Wbi7UFtJEIRCgYcuuUg0ln73g3qGY7JqaxRyLCNuOgEeb
mfhE+uEj24AMD365F0G5S/nv/IhbWvGW240b+LyYgydl3UEudmcTsjY+/2vfOvXw
omkQKMJKJjj7umv5VLrT9w==
`protect END_PROTECTED
