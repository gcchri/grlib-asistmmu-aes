`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yI8xffH5b3MvrZ60L0p+fdqy+Z94zeBq3YP0kGwXa1LITZm3ZJflin521EBAkSI9
RIZqRohSTUYPoQnbgsuJ2CygGpB8hheHqDCzSziuRfYzU4a5+4KodnWXOYL5JE77
uvORNoYF0cuPqbT2QOzevy51IiOWXATqlUl71Bj99AF9t31J0diDVdvDGjj7Lr+s
wTIbvtewbvirwR9PuaGRGmFbOxkFafjS48UNF4DtOU2DHB9PC077S8ymK2vY/Rqa
P0DqF9RdJlYJedPqOLwJ7q0QLZpe8KMxO4ItbpI8443F4r9d34bTCUeZ3tqCvvvd
O+lUje+MHB2tukxeoieKlzGf64wkxrYwpvgiT8dxxTrr+cyEFAVhsO1tjVaxfdQx
5+Kc/P5IBPqZ78elrqMzhMdrcBAbI7gLGN1uOhgRNP/18iNu6fOJnC+0PwMRJY3s
3Dn/7O4ivlai8KnmWR0Qy9s1Ad+ydOpsnXVBFDIUcspedPnMHXnDDngNAtruygM7
C0OnqPPW9iaEpl2rMt7Xg2GH1H5uhkyYTFS8deBirrSk/Zl98keYZaflcXNYmXSV
uFTa2OzkEDuwa72vBfD76PHu3sO3o6csVNel8fOYk4y8BE0MqUkwM/maeXzZrtCq
nIL4DUDdEjsFOdAJ9MKdVN6hUAEJeM8cydR/eTILbvTkNo89JHheXqR5vCapaui1
TaA40XJH0SN7biOD2KVW2SExYtG0uvJ0sgmFORpzdN+PFy0oKvygrws58sSAUktm
TqExQY9hv18UcfyBjx3hNp2nnk2QcyvEgAZm6T+sG/dy2yOKFSiJGPwfWfkjzcy/
0Po/2d/auvTsSBvW5QqCAw==
`protect END_PROTECTED
