`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s04Z+T5en6Ei5ORC8fLeINcf/m3rD94f7DW7DkG6YInDPv7odxY/z5hT9O6etP2L
A1gmf/7/mEHBE2XOV/psXXBec2tnNT8YSLhfZIRYTTEICjSP6CPaDMfhR/bE4NxU
1ShsX8kZ89vszc44+NdzLegdu0sX1Gu1nOeahn9QfSPU8KaiIvTRQfyI3G7USggf
K/B2UOOBl76T9pAkiGUQLgeFLx9Ot9Yl2ywJQ0x8/aMDCEbSxaxyqQUTP09wEyKG
Kxuj7Lq0S45gyg3eMN+ggYnf2GmuP4+qyqNYuVdiEqhpLA3cY4D5n4nHQtMz/QO4
RoSFCXVJqrzU/TvPUws94sZlD+8PYAd2Z5bmV1TdyZW54DdBxHuN0AYnEaYJsVzH
rJPRnOmwYIZTcCyY5++4iWndL3PiGZHchzlyjm9tAMm7LyII2S9Nu/0lBfwX7PAc
cZjshC3LNUOMLh8MC0bSZ6I6+ExGGxy/IquZ2tBXv+Wdp3LWU5kTqpjHvlxUAq7F
yu8sk1uoQRt/2zHzN3AIyFvPwnPAM6rVsIygmSQNdmmUy2TzEQs41lYHX1Xa3X7c
BQncMhAkK8lYIIs1O2S6GfIbMS/qnsKX+uVGpCO4RlBdR7a+pB9a9QcYnb3R2kbb
XusVznkvI0ZAJ6uW90moPUcCi646kA/izPQ7S2wszWHGZblX8xD+C4l5ckySZBOg
xkLk7eU97G4GSLt25/0w/1DNzcmL32EolllsmnCXSbKMMDtcobF11p1FRlqW01kt
KvnX6iXzxODuzW0069miScXGTeIJytO0WsM+NQUw01UYa8CtJfSvImhxhxdsCwm3
JWTHBdF6laj5pXQ0sxI3drISVpF/exNbZLGP4zadAUh9M3Yog4AKXRIA1PYfxqO6
iftFd0+UD81bQplVFS1myzAohIGZL8Egvnowzlkpfu57DBAYSBjVKCK6CX62vjmo
vJMNTSrMzTrF2vMZNpqRQ42IN2SIKj3DmfS26ICecU9DmpdSQejNXxfq26DiEHJe
RwzRFbqjB+yklk3J9I6irCjDVKWPvDJCfYj3ImoF6FlPICAUZxTk6f/xlx8MWwtn
`protect END_PROTECTED
