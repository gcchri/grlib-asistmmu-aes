`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rOHrJE4Zx6zd2ScjJwFYotYkFpKElDDEQbd8XjHFdnYeu/K6NuLK8o26lJBefVd1
WQPWyKGgyM54trRG22O6aCC4DxY82LTYyvU7jLkcBt3vZCOtkGaL5gdUDRRcZiKo
Yo/X5D5CRrg+rQte50CIgo+5i+DXPEkN+hEudZRHta6NndQrlFh6d1/aFPklxSt0
x0DSH0pUqNMn/IRz9AnfPatgySsKJP5KsVFuzkfVJHOz+TZyHYoMlzN1nXZhWKQU
j/p7UwPsuZ+eI+b2KuxVJg==
`protect END_PROTECTED
