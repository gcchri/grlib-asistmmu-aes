`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oOGcupVvEkf97cS8bNga6DgGXlNBtXonQZCMxtZ+sRqK+oQF5TaIEaAk3B5cewyF
LYUTlKTSKnu9Zjw0oPjzOOgmxxbU9xl0PwOyZSmCrSHv2AN758p1ttN0E8bTzour
f4L9OZ3l8fQD3haC/aFjlXvBpedv7hV55ZrBUkhIQTc6+0xThyhRnsLXL6PxEwDi
S38IjTvPllAhRw66x+X53VwggQHpBs7oGfWYwn+7f40rPFZAZiPfaIJ3h8EM3rQs
EP+vhl7SFCFJDOmiahFJgaSKOF63T7kRlvGtYGYrzKrXA5oBtTjXcyXKJlwAdnjG
6n+vcLbkpVI1NpF5QuXrvpD+yNvDbrp0jd2BQZwzv54dWl6kI3XelTlAkyD3rYY1
1UPlPJgq6Qaz5AkvmZzXOKhSbI39/7vjP69imdGlbTJ4oznZIdwNx/BqyibT7XN1
AlzDYPjCk6AvNmwoB+D6t1SJ/C5B4Yrz1VIgEtbPU5NoU+Pdlz3sl5mmW1ncCNdH
TCHM9latsO7SEsdy/jiBKg4msxxXJVwotK7S80AIz6Zx93BscFtYWJPvfE+5bzYX
749mTqFgaYzBjGP1VtMZdeFoON6o2qGf2gb8IYCgHh1JbYW5gSfp1dkysHJAowbk
CpSuU/5kFYL2ggKV1l+uvrriXnoeH28/AraaUmFwkrCEesYfGtueNXIGhBkFQGvW
htd+9AXSo4dKkno6mww8i9+EvQL8g+pAQISNolJJAhBU1QS3/VffqDFy5mVmwzX/
/edE7BrZEmi5aGT2SDEisgjy6reVhoN8Pv7ZNYyolba7oQl1PjmihfIrhzKc38t4
MHqWaKXe4+3AXci9pVNkIWNhcfpUmmMbfE8U7M+fQj6GgtrvqQMvNA3RBOttODAF
/cltM5ETCns+DwE/3zvsCX4jo1v0SN2h4QjqO68JY6CHvhcBOnG7WkUIf090ckq7
LwJD3b+/sJj5ZmDRegVHquMXDk7OnNNpe6c1i8rHw76J1Iw/llnktiPEC0o1VZ8F
zTAvRaMP3nde9UM08aJBWz6pRH9jF+yBixe1nmX4ZanGxavQ/UZwHmVeQuQWpUf6
G2oN9DDKbXglZiVtKvEuubE4cRqKFt0j5Fkjp9vWkgQq3ev3zzylM70u1lCkX5uv
TxSCfnSOV/UV5lGP1dlVa3KOSIV5WccBwpApWyaZdG0+XjEFpiTZ0Ivk6zd8q33L
CxlIUmWu2jOqhOtSUhC1ZAAPy9hJc2CcsGmQirTq85TmQANsr0WnNFhm5M4cx3oA
ByUwyJsorjT/a3H6dk/n5zUqqJovrR9HANzmragYt8WKzJJfK8jl0B9ZRU9ZccD8
MHeHuqEWJvulqBSN6N2Mf6LsjNEPURp0Xqo7deMR3JKTRlmq6JOQFGRw0MhsFANk
v3/ItunUX3UFxmUQrGrAUr7z6S0AwO6NsTIAyIRFQe0oVrN9fuagJPju4NeMgPLR
0PdUljY8MDIQNOzpZbVpZIo9g4Wk25aGAuimbhQCC7XdiOx3LmzJDAhBj6za9R1K
QUDt8PSsVfGcj/vgaYZMGWurioeAwsrFQvVpf/9W0d0/LqS+XY6EIO2OgSfqHKzm
SNzhfLyaHaMvUeZKi+faNjGNG/Q+eFnPnLbUXzNtlyunHuNIa2GOydj3DlkelEIi
qVV+4f4iTVrQNf/P+Xz1xO3t6tF5IIVtH3C6xd/O9zXbqXn79tu1kR5V3HnndGAs
FSmNzKaYHz8P3FdqfJvy9a4ci8/dJZQHrg7c3C3CVkE+B7kV54h3+CVRL5wLTY3u
D4w9UCvpfRHWek2eHjoH5AoGh2PbDfHSFF6pBb7F1RCh6fqVPBBjY+YdRo6vLc+K
MiyNSnwlnc8wGmK4uscbmUJEqZxo43+H3uJjbgVQ7FK/IOI7Br1sjAU5rmmzMMCJ
Ax60kChrZ3h7ccdT5+Q6TzBiYd7ttbKshPjJTcdTStlPS6rKHskJlI+2eULI9r89
onqwYBLgJ/ZjWXL4ManPqJPNkK6KGSWCMbukIS2E5eFTYsAWSgbDwvUIVRNnrWMC
fGlQlUwuQHC5P4NgdkoRM31qONm3yBefDaHUeP6u54ANj4lGmb4iWKUJa67ZLDZc
+6GcZcbWQqQPmasMyOByVzjQYVmKPWQ4kibfnhh/Nu504QE1yt+p/VCU0/toi4tA
wqm0JON8dKtdHiGXB92SkGrizwU+jwsqTAx7uGGZDQUDQ5gBjzsBJes/B1fYsX2g
F4PQxe9fAu977JnJ6IR8pttkbLyuDxqtbb0KMVR8qWX86xEqCdicr/Nze2ZJr/+Z
BYDdUgiJ48htEjHNfIZiADRUmiSNBeV7VpWpcuhmpnCJbvQz3GmGUY+1Kjy9sdns
63i9lAsgL4kkYsMKvxRa+zoH0H0DAHnXuUpkUp7PfiF054hfOR+uIAPfj5Oie+wJ
lDFU3yfIIEtFdT6g7iOTuYjP/1gsjPyXP2wiNX+ZY1T9nblAmYFd6/uSbSDggKDn
VdfehGtL+HuyMs+Hv15ZHfmi2ObpJodnilxwh1vorL2DD6AGxRf8ofS/kX1AFGI+
0fZ0UZJW43d20iQn0lzawOTMl5UIgQw358K2CM/kTC3hf8+xW+T0mj6zwlVL1p9I
V2kqk2vLaGvHEz6u2u24uR/oTkPSHtMK17k2KnR/ttr/AAy+tIuxQ13f4Q2OVPMe
+tXRwGz1DuCPqn59MsrZo68+klbrrA+tcDGtjznUmeJ8lPgofsHUQzY6LlQUm2xX
0tY6/Ni7+1jVamsNscNCHz9f03iUR4/13QE867ZSz/uOo8HxA4C6GmbEs8hmW2ol
4nGNCqBcV5Qbk2c/DFntLpmgh6VU1LE680cTGduc6/KUnoxDoRbtMu//3Ooyzk5+
KQ6ra0Cw3Ot0CM5R614sPMm8okBlsd1llYRzj3Rl8PXQLKVHTgrhmmyNRPTno6ur
ZZ47bN3fmPuz1zASwayx1aeyZvG2xVFR9FJ6sj6O8SqWzWLg3KDpu5UivFtM6Wyb
nu10gyerysz1ILW7yqTaiCuomD+lB/jAmsbtLBciMDTn6kYLEaEOq/Ho9FL1XYEX
48O4vjo5XJKphPNIpi47H2L2LBUVtSfvB1YmoYOTDzCAiWS95oVnUdc0927ukWSC
zSPiOHLLObUahinNWTIimT9vs/0xCw7YR148H/bjQipLFCxEXEeppnE0UEuPr2KK
Tu6tOBeDM8fMcc6iq4r0CO1QW3eTBY8Ty6FWsxhFFF9hE0Zg9Zy38ao2ppKDbRsr
querwtDq6UJdd4Wi4yPwFQYr8OZw5IodCH75rp/9XQLKzd4wAaEvXqM4XxtNQAVZ
/ig+tsWf8at4kUMTszrNuVdr9fi9QM/LIVsnLVaI4i0EIJIj/4ornCiN/Qk3/J0A
+DJICymLhD1yyDfLEUv4ZvH2i0ImvklTLez+7//C6VEshjReLvtYJOL/a3mhL4nm
CNp1v8iDySj8J2zgidAn5O4KjDGTSOBkn4GoDGLlFxzJplQDVdC+wkqxaOZzRkzU
3t2A1mOEwI/L2p9hnk3guUVEQXzojg+12mz6LS8Pp2/wLgjDyP3uLXdSxhmLJT2/
Pswhp3UolVmIZ3vSIWldsS0nU2eXN99LUkNDy516wAi14srvCSwfezOHtB3UmcE8
7NLH7Kprb3nWlEqYP5nl16TlK2e6zq20pDvqA7WpWCDddNuH+aEQiYhpTpw5P23t
Gx6EMD4LLVD5vSCtziejwbSzwRv+3QakRNisqfULHBELAO4TGefAw3VjwFOKLTpG
lpyXUD1k2rdPZU/ojhUXFEsyU7PY+JjgQXzZXvzQFG2yeAZXyaDJgskL/m1Z5+HS
/yEcKlAVerLGq1BkllzV4lBZLHxWED3P4mk6B+0yKCsskg17vwbcWlZRxRwCV3xf
0TEuXxuBQvif3HbiKLvtaRTpLwycE50Uiyn62iF3CWlgqW0AZ7A1yLe4dBHmohgr
4ZiFb4nLNaM14jnUv4jCHcY7nj4Fx4r79BsYEqLgM0srsSd7PkaTgbvlzouN2icC
/I3C2vFfRXxXmv48dcUYJTlnSCUuIAOyBhmdNy2IXOXNSoPqSvv2n+DzXkJ7sG+c
W8O0Lk6YJZsmcGQ+aLHiMH4Ai2kR2iOtHROe8Rl5MJ6QnVR2V3R1cfAwUgwACroy
tag6XeChEVLgkwnQx4Vk+swU4fa/ZH3MbZ/2nlXKtQJCT/W9Voyy9mmdS4brbCr3
ym39hClkW4AiDluKtVaowULD4QxWrzc+7iQE2T3LCIh2B3oFO95aTKU6uPr1KXKE
nAwqp2okWKrBQSFruikhrfyTBy6IWcaTeg6Ode0bWuFGE3Zk7L2DgSPgKEii47Vx
fbAuY/w12SDCkJTUTyUo5W3HGGRVcF0LBA2hkg+6/z4uPoGsH9TmqBocx9iGgrZz
oKo63rkfYKh6Q7DOl0NXNYM8/TrNicaWDV+dGy4us/h50tcx3VfDCDsq8IpG4A/S
JKbI4ZYjkN8oYI7lUetSUHFLKWH5dFNsl9ABE0edXAXMOZCVA/B83J44opUToD3C
McSvf1RI+3XkuiYhx8wt1kQcdPczIWyDWrfJCt8+ngenQQP2s76PTaMiWqaIF+Qu
g7ugAhOn5hSf9wc/jQuD6emYTgVQF4CArI8QR5c4vU8p1tJ5RDBrADNw9ec13s2n
U3dyizlJlP1Ts7Dve8EgGybJN1rnJxcvlBIDmIU5CisSBrkoP2ahxtSRlETpRTUX
sXvSSkRPmhySWuzw8BbPg4XfNqho2oJFELYTEe/L3ovVxNv01xL4RMrnOhAA6zTz
KKmJDpVg0epr9Y2dB2x9slaRrSyggZku/9PwV8oqoTEaYpcFMK+VEAwGH470HNpK
c8BZbTCfAIzNE5CRkGfFiVoDxU51XK2x0itqK4M3/lHYboULx8JAUsjwvxhkSuFj
1VRsgNirGjiUbgVR9ac1Tk3CwwA171a1GtJaKXa5aFe6b5kgxFX2YrNiJG+1ZJyC
La7ANpx1iYV6W/3CpNZ33M6GTrE6s0pecIr1eG0YhotYZdvEtBahIXYfcsnSRfdu
4dk12HphIJm2gj6ka6+aE4P8eRX8CMcxAzVd5kCsBEbCz+A2H5WJTIIoKZzLSHpp
wJWaUrgGUfa5Lyopb4fsOo5ANCwaW5R4K1qlm8YQ8EFuGKJLZHvqVfwHEfCN6Y9A
7mQdPZpXhyphSn1xDDbHAGTeE4ERMViLXcIP1MZK89uukz5uGW9slmxCYToXmaAI
IzUQNHR4ZPaliha1q+DH25+ZfxA0EHMr1d4SFAmVC3KgGdhZkKT54urbO/qfG0hM
RnWq3Gxefr/3k2R4iykL+KnUy1Zb8nM39h4TRl6mGXFFuk8CoiddApnUC4FBf/9+
XL5mvvl5D+7zfqMNZL4JRBUSVLen3FNtDzAxMWYLlYAFkq4pssovrWi5dCghPyu3
EwC10ezx5AylsvlOmc6yHOcw6TqAN+VAh5c/lZ5qEdt/DRPiKvKs3oDEqycaB0P7
Vf3JPcea3uR1dNg+2dkujTHIFQfFi0eLcDCQPCNB9yc9nhNczMTzx5YG3wUfAOfT
cgfbvd3I0bmtbLvSxaKKcNY4TroMI1AKJF35sLFJA1DDAUgQCuLZWtBl1VZCthm2
GUSaZHy3bPlkKxDdtc5Pp1FrN900B+9JvwZcvsZFgtnX4in8iQ0GMYUFs82pIaER
12C+x/K/FVVqJ/YTQCUaPXTwz+rpChHzaY0FGAwuiGz0XbYKBYcw485t2WLekfDo
bapqXHNRVqDD966A4+GB4gQfcMjaW+TukWnJPHw1bzO9apB3MufsKv6661DwIDpV
tHXh6oWTjD8BslltUuw+OsmExnQNL7lX5+SNsCkDv94yFEagbuBtjIjaFpkg0nKd
7m06MZtSni+9L284h/7rw+2xoIhrjZ3YFZgoB6+OkOhlT2ei5UPidhdfpBUe2QFU
3mpRBDTFKetkWfeuuC4PjxgY8FcrTkrsgTwhVOfkH3MJR9p01hyPcsLMryI/VMdJ
ccIaPh/khXmOC163W9+M2MuJl9WqBBBKbW2IOcszDB+aBXDuGppegLz2W7cajYb1
/NLwH8vrXarl5DkfDrcprwKNWyGDIGXeNjP+Q7Y5hoAYaDKvHeCpSLHFpks/MR0f
hxxLP+sRhu+5+kopJ+zkdp0aGnV5Pihrz1fQhogAN4C5TSBBBX6cbitj2s3D54cK
/NY9O1AGAPJ8XL9aJB1UwoeM95Wy0ZmMR+IaOxSnbxdqfikcQOrOx6ol/VNZAyTF
Hfy2Mg0LfpbKszZGP2QzRHsKbihsVJ1z+IbyI0aRBF55y1MnHX1FUwMyvoB1zGMR
qtUAA8odV4AQMZYIlQiweHNaAjCY2f3k0eqIS0WQBb6HMhjgRNSoXrW2z7g4aBn3
VrlQz/v82DIM50eve95WDiRUPxb66T92R+wNQngXxHOhdlKdj+tN4vPEuRkaLS4Y
/6K+00d1+cVLDSBslCt9Ig9Gcu3R6BO6Wx/gYvS0t0ICVFzB8C9ydtUmRn6+sWBQ
hC5eC76ggMz/UNiw8X/F9ii94NkcfMtzjp4RWIueRc0Y4YJ4OI7IiSiuQawOqVSC
5NAFguQKq3sil6itADkykfrKuanh0IZuDgUYNHhfIbRUNOB6NguPF0ofwBp7yKvT
zI0Z+7heTteJ9P+AQHM0/69tT7Mgy7FltPrWiX7cDBA+n7Xqlj4aN9cTlQISJWxz
0Vc+ledzbEhar/kWWVtup+N5Iu+9rrc0ov7PYP5n4QEfaQXHiD+OsmEgZEoto8eO
ne8iNiSyXXF/6Iq4XA1hXmt6ug/MR3NgqcTTAxAsLxKYUVslJ3ROVzzs7aAWYd33
vll8RCL1XPfhRwz/o2ZOLc2FDZ+/RX5u/A12WHPMFcvwokEAi42//OlqaV+rFoi7
9R94lw45RUI24N+FfTFbiHDarPqbkWy4ON7JcsqR0XjcvlgRDDVA3uvhF64jXAxM
dPf7r4d1HwtsOWOFsPWyNf8oifcT1oy1JM8Uan2FASVG8bZVxr/wq0VwSmLupEIm
P8mQoitoO1xKw7d1j8d+nkp2f+pVbFIwQOsC3GayNnwgYIhHOPDyrDK+P6b07ILx
MEva3GKnpLzEsLg0Dvr160sbnaQzbuwj2EVb19NHw7Y1IZ716pXx4joFQuDwDJ82
j/MVlYbn6QcOJEwyLYZC14ACyw0Y03MiIGfbkl22f77bXRL8dCF1+wzmXzTolSP6
goxXnBInb7g2ut5iQIhDBO3TSXMu8SXX9PXUnVzGwPOah0Z2b+uP19kylAFJnEjq
1vC/+RtdBB8u10zxH1lzi8EOJ+5Wbk/xNnmWoxbpuB1ZdizgmvMghVFrT9yr+YKq
7V38bYkFdHghhetGx6AkxI9TSc4KLB6TnyJ7vKPvpSiAckfQl+NlP014QP8FpW3K
yVkMwtX62ewDoc3rbc+xG0REGiZ/7fp6xEoZZjCgo+OdH1521G/rhRtJl854UZrt
6kPPLjWm2Anom1o527IfQdSq52msI6BZI2XOxWnc3HOpBJqgO8nzWUVRdiHTMoF3
BIxBZMZ+bvbLmTeUxqppeJudAttni8WWrlY3vbTLODn0JXzm6DHftuAwCr+KSyUS
ETta0GYDYGd7rFLu52AAoA9+Twpk3fPV+NL2+tnbXw0SJGeEvWaNC8S+JDuYwiB2
HyfZ9iAr1oqMPjv1VBM2h0ELZNyeSq+pz3gF8QmahbnMpV+nlwJxAVyxl6NaPEJw
LNwUz2pGHzXDGLSD8A9RWflR5CL56FikPD7jdSiko9k4kHSGGO44F30f6iGcksuX
KgU52PrHl4wWEiKsrucPdRRo89L83xgXzoH3IpHOodJTV1NO75rhEMa06cBwZePF
KP9HPOk1rx++0+tocxNlKAjL36EW/wfN9wmlBwoLod/HVPz1c/FVlzi55SOYgTjm
XgRaSCAN36fKAGt2+/HKz49EP2qBAJW+pPNkbsjba1//zArd7nUNEIdSIdu5UOPA
cIiXl+I736tooqi5FXBlxxK/XgNn4QpTPfD73WyssbGHNn/CiMhqWPtlmJuRrqX6
OgD28BqR9R80ZfNy+kfrNwO8zN6AdjjiI5ALvW5PT4a/082+mweVQMFOaGX9QOUF
DIM8hneS6pUv/USALuHMNCWkVdn4tPbzBYXkeDfE6Eb67n+SAVxhBkOoPciuB0kF
wJf+GkHM47AIajJrHf31faVVZsH4WUCES7Etv/659jpbwRyZhoUyBMAgCBs+L5bC
TsnWDdxUzdcwIgZ91DMm94g4X5fnmif3gxvuvsDe67gC9/sf4wQOYJI1K2PCnHjB
Sg3ZpaoYq/G6u1Kmu/8qGs+Hse8ybqmN8iWKVHZISRncCZ4Ly6sTC4WcAlWu0/YU
ebJvdFCyuc3zQQSvI3JXmmdKErnDx2ap4P4uVQFP8HlYFtEC7hwy5hEbxJ7dUzEs
Ct42mDkRSHuVLy8rkfM3Rk+oKghgRilo9i6jUpmhhWHLmAAsvoGqEhzTwXuGGedu
pbY0RoIQig0QlzqHHKyYdrLrqpOhRblm6ltElc9FjGCgD6Rr6sfeFIUzo292C8Rs
RLLgZ3luym6Ovu6R7EwunZMdPDp0sY4o4VKVRRGdOmp7eHtWIgIsgOpGF6OMdmia
RYCO4LgTQ3NmuF0if1MB/3D0aFM2XtVhLQuM+Aa23tt8U/YjeXmqfNNCi4VQ4wLe
P834OiWw0PtSdxeFFabAPBu3y71OSq+HQFfwkkn9NUI+Ig+EcsvFXmOdeztOKA8I
/R1JmB4dQzrNmY7jYN7mMbvdL1XI1R5yEDLn2K0ojJ71pqAS9MMJdsDtX7fdoHj9
Ej5CKp2iILW+tOz20+5gIwjn7gYqn8bmuBtXglgNM/Lel0k+i6gBk50YuahxP/32
vt4tgsTQ8hGcyIqiJblD5sMHzzxdQMZnUFmo5Gu+6+VmGXiI5jULVqqmjRQ1Un0L
Ivc4oXmIAw755ngkSHTMEVlS5rIdqXeLAIZnmOQuxn6sWyNGQk4LcCdNOnLGpF/r
bVZPegcGq82MIRnCNG6CwdDmT34Dksm0qepyYRh88OA9uf3uEFCcQbNv8J2kkl58
cnjFvL/lzwvXttBpf7H0LyzZNdpzABxEhKt6n6dnLelFYP6ziWEeTxu67Qyet8Lf
lNZfCx0iZznWKjR9kgbLBRe5lKiUT2pEA3jmyPlj9uCH9NWXSfg4NFJEa8ldKuwD
gSDCBtiVotnQp/Tgq3mwlJ1eAJTK2DmDiKk2jTJ8BkVPPmAeqNvp87jmSE9QARgn
NdW8B8mG+JOuQDGRYQheTQcvKgl0OrhaKCr8krVyV4yI0uS+On6qhysqdgNb4Ahx
DszWeHqoGPrnmcXcOLW/A6dkWJSBRHiqjNjrGE4YnKXm7qKQb6qHcpZf5GaArgxH
7Uv2S1afnpI++oDjADbOpQPfzYVwwRoyRA1IYalIDCR23Xc39SXI261jKsxSGyY5
+swWb+M8K1dnGw6ewwAWWBjxJz+vcAS6emQw9zsoqoa38R4lrmqb9pLA/YAfFRje
Pu20oxYfWHhlAz7GwAUzEh4unHkCfLr6Gz3fAxdlyU677ALNFrXrNCiolgCBIBGG
D5ooYqz+oxPe+XPowJK7b7q0qTSXwYxfuOp05y/zASTdjOm7bCWv5oCbrWyv51Iw
jPM+0dq+DsQqz/6dgKVDrjFOSuAgNGG3699XM/ZZkXAqI+CTMvulBkQhLWnVfBgw
CQ0nWDi99X/hYrpkcYvGPV+ofsLUujT9su/UEgxTVp0VbfX0eT+JsiWyVR2GoJqg
JZqOfhkT52q1UmH+F8Imq7guCXnamsomEPbnIfnCWJ/rcmMtyVunHmQi+2berpIu
x5Z9jSPDXORyVpOjyWSbDzUjJj1UxnI/567YaAtq0xJlXsEwXdcF/tI8PHbeer8m
O0hhUaFhWT+bW6bNIp/FcmFY8vaGiPJhkKCqo73EbyuFR/8vE1aIQ2BcANzIwq/C
Isg0lPZ/lv9uuWCHHdXGCsWt889i3t0Fv0pAFjHsLAOmCymkfK9txG9CkCfCWSCJ
0d7PT/W90uBHZ/YsJHGJKDUKQg2tD3s44jcdXhghNrABSo66T0C7/DQuPj709wJE
gVe9u88N9OOAiaZdQRHc3d1vIyB82UBNeT36y6s6NsPkDfRplLyQgU4EUsLX2jwo
H0PqzM4nIRga9D9z36zz8kbZpBNF42OFPUIgdvfm4ozgIgQFiEqCnY8lo1D1jxip
LtsHIRefJ370m3jRdAZBVhUoVW9Pcoo6Q/Jxuz70aqiQk2sd66UwJAsMZUtfTK0Q
+Z9F4fjdnPh6uxdjYQdizVjAAs+ESWMXXnE8/1oKtjTClE1z7evXy5NjFZNIz7fG
4g8NbDq1RN3V89v91IbyzHCiYC33jQMAxQjcm5hrMEuMesK8vqQypbcE9wmv7i+u
gDHqi5WxxB6WTqSR6gn2fLQZ6T+ZYS3H3vpRc1YM+QtH9r3C6SXQlLnskYlgoxvv
nuCIDF4rjQHHXEH+AEo/HLGQVCy4EPZ9uf+mVZVHTah3hyOv5yt67I1/H4YI+7r9
6d1cW2Zs4uEqJXFLuznwoBX4Vq1T6dKq0XssOEprOqdWVm5fdg2iRyIqX27K6xzw
fMs8uyyIvXznzX4JkT8oOoDBtN4RgQYm1n7yAUZBGYDyuVjSB4FCfT+U/Cxl5kYp
thRucmN3Cq122pBpnmPhsANneR2p7a/YaD072StMFYAw5yZow2gqvoeTniW/iiYS
6WAzEpj2RAPWNByiDCKanbQYrrzX0C7RLyySM89rcRwctUk+uWmOdvkgmbTaIffW
sz6C7Qo6QbwXJn/TaB57dBNS6b/AJrFqlyR24f5gAZH+OL/b6ovtzFGvv5GAqtLR
KJysMvYsQUVwudkmcC027XO0z2a+gpOojuzfYcgVfCZPDGRCDVISV3wMA+tSTh/I
WEFwLGTNjUXvG9BcMKU2sBdsPMqEE84wumLNTnPYvWeW9C+nryp/oJyYSisoSJKX
bcI2myIel1Q5TOxEcBHet+LEqfhsn61K0KIBnC1UnDNucQZwfntMYxuVGCgC6Tuv
4fdOf0QlYUXxZgKYpS/DaqBbLnoDLnskAtGzeB/iWD41zvcIr+k57xg20jguOBby
Ce58LCs1Xbq9chgzVCDk3zuDQm0X4PVsYiztm2U9F8/9bc8ZKIKbwA+i4DW5OzT0
0T0Ch4Qk1tsfuqf8ZlLklDRxKWZ+UYCka0sIRjJB+XGQ0bdt88xxaJ1tB9ZFSGde
85cGtTEKY/nnzkKae3/yFNwrlNnQoXlbOCHRPINTKWRmwncgU9vmVMgT8j1iv0Id
ZAHvjg7/5tr63P69yYPA31jHzM8z1U/W/poyEIECGLDbaN/bFsePwoZq8YL9Eqjs
EkLc+FWzacPweHgz8u+9fJfzATiwDK/OOQzC2Rnc0ZWNDR+NKXihPwyRiVNoYlH4
rzWZJUBFf8USqoxwUpQW/OIiTt1Q0YEo6F4o0Fa7uKNPCbVtKQpn2WQDhuPZh6Qn
SYIZpdAwTDLMSZILA2QHWbod/zvsjcfPCfDYRGBdOsw38eINwiObELHajFSmN20/
wLaveaDrYws+EQgKX9pArIYS3N2MP7cElz1np8oGlPc56IXiP+vr3mLg1aX+bLdz
zc7Rp47RUW7YUWv8VhX6dE+rYpsVjmey/x/0sIZvo5ttcsgDc32QiBTBSO0AfiIH
KeSddp3FJ/1k3Vo9aWzt3cnCZSNzvBxCfGrvpOKB5gZGZ8FFuMtjWDIYYlm8g9WP
2SAaBiWqBdUY53S9ikRoEZOXpVUs1WIV2fcZozPMoHDVI+HmaQvlSFl3oZBHHCnj
S+jnx5s97vr4AqXlumBjsqGtDcv0k3HluzOWb+A2zHpYuqoYrTFg9Fasna7lICLZ
/pBpf1FEX7a10ounIiCRWVHuE0ixQVYI9ZWEnWEYoLm/4R856RbbG/dYucfx84el
+W8PasHuqvGlDBENLH+oqC9v/weW28tsdaLKUv2MjvNwoh9/0VURanqttmtGYGV4
ddAWTfcB5S6yKAT+sO7CTbaHlyR6LL/lTPMwUHllwnEjp62SqnkSZNEA4DJpZPJl
PNfmnuCerZtuwwLh/Ge21iun3nw/n41/zbXoRjw18pTnR4gIsaObsiPwDWIXHPSf
S30IGr+DFUUuTpk35MCT7E5SUsdwbOvG7GHpBfdQEHoqWW00APCg2QcGQi86VEHa
K02Y9pPBW7dX5rbB8D0HkQY7n1upDR89K+USJ4hYXOBkHl9WXuvBebU2zX6iLHcD
EU2I1qUowBiHMQ/5FLz0wJCPdaG8gvFN+iFUeHOMlvEMWtT92Kv6UYS9jc6dF2Hd
huOG1dK0ajP8dO15adL3bEZ6IwrBuD18U+awqvGbVxkIv4O4AXs3o4I1P/cztH3J
ieNABRFmyxQ3tQAx8BdDrKoi7nQ08GJIMPAQJXGFpmCkwiuedwk4TzvexmmixnIE
+rztSZnR8vwdW5rqOVjIaF6CJATSH7w1Kqi3R8HujCW9Tzt5FFzVU/psOrVDHaV8
rzVH2oPW4Gt5G2FbQZWm9csYqZbvdf/ZtxAs+2bhRr0=
`protect END_PROTECTED
