`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PhSheYxKYloa1r3Kmia03P0/Vc2Y2nLyDoe5x7dVGVseLmEARCxLfFwqPJW6bbRw
bTXj4mVcUG8UbbGD+yYBh+xfP3o3xxwSP1PquUQgfpReKgRrW5Go7ZaoZQMKYtNk
0VslL18b/IbleDtG3VjDhQC4qSFoOgTAVUIfzQ5tiqLeQBOoB1lJxAJYJoCbQJFK
ktLFSuZe3R4xoswqlVRzYXIrkV1CU0/ILo/r/hG1hxRy2xpyO5jwe9dpzB5elU0r
z7miUMzsn8r1PNo6R+sDJxUdWslJKD5c9kRMqFdH/eVCXbwqKCo8pcgPUobYqkej
D84FyRkXsggxCSBHE82icmKy0yLqRQIKCuQo/ZlewwI8cRtCb18tsFG6mvXcSD45
PYa56ECf3Ud+BeoCXTekNFG3sgDz0Daj+a9PIvehjFNdpn4oHPomRV5MN4kJtLRi
2+7RVJ6kC2ekkaB+R9elK/uch7A8oEkcFxToZwIds2+jOCVKOLl6PUNw34J/rMPB
0lZeftJw7A3BoJooBIe9/oMaAR9VwrI5yRltk/8aNG9tGEk0cZlCuRO3CKV5+0KP
RtgUMPrUqObz979rojywapFV2L+NP1cBfnsyhYaDYhSzpcmo7+78XJ0JXDHSLtK0
ZXE3Q+WS/sb3/rf6kAL/chfaicyqyDL1cLWigMEFKVPrqWpZmVhPvGtYxCswwIfV
hRfJOz4JZSflrtSsj3LOD/cUyV9jgubjv1TSiMvmVXNsvCwBk1dXdzoxVobv56Q8
kUjdPWqEfaZafW4zfXngOAWRRoQEstId9TrXRmndSwolEA9q8K/Eb4owtJx5Scpl
1Njpal0RKfhPlrOywt1EK9xdsxqcYj2OwV2QUNSWGyyfh0xhSuPGKHplweNClCDr
OV6Ogx/2SeC1eFJf9ufqybCkc2zfWkyoTOqdtYIfoOXu9KluU81sq+lWEVKB2/ss
A0Uoxw+YcXAyPr87LUfnVQCv8xw3dnljmIXHQY4agn8CbEZIqwJa8v9J6LE1UyPJ
fjT4YOQwNgfldg93cuiXI2pgXnaNbXXTRC3yJJBicXrTf+OscdMA4DJ8ccfzpZdy
Mi7dIbd3vOoL/kQxb1lGQE4RnRBTaJj5edwRs/F4PTYwCgiyTf7gZ1S74i4YEC7J
nINuo0Tu9GSeG+WhZu/IZf8/8m5kol9Ik5Nxl6OldVvTpdIUQ1OzEh7EdGtNnziO
UZPNeQvcLSC0r2uBVz3fqf/WY2Mt2i9MVK6VSqpDo9Tb1WZur/Svmdd6pzhbNWqf
axOnguCmqdVHPugalMQ82pvp6DFUJIQIiNIjxyRqpKRbZqLPzRYR/zxdxA7BjBhx
6Ga53wqOGur3ujQdLkeig8QI7JMM045tUTY07/n03XQxxXM+VThLv4xPfWCpQ1ga
/Frn5wPoe7dsyXMZdg6/ZxauIPjVhwKdVJVVdzf30qkstfNRETNLvCkvZmXryvEt
xJkrA+Lja+eGBVID2L+hNg==
`protect END_PROTECTED
