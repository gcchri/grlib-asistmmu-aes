`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ADn89/j4FmpyMsyvFt4ESWFz3HsEWWgOsP7KgEROunEtZfSwO7y9hotq3e39fplv
ije0q4D4+Y1KFr3LVtgvLNbIIjTdp6q1DInKmFga7UK3xCUb4lAXaeu6kuTsoc/z
isLpbLrpkT3XexkFch0nkVX0TI6/vxlAI5DwSlAScRGTAofSbsITi+Mb+rqapW7o
Ce0MFsb1h0kwC5IMNJOR9PDWhMu1IRw+RgfcY5UQxTShYQvoosRLyTgHy6KoN1ju
BFvV5fLSMWMPrXeWBdrGDEArEyHE8gXMLeBb8SIh98X+3zTRtscsWZo5etAkKP66
0SmMYu/s9ZQChsJWR2doMegJNHonrEdygSQWjxOv/scsaRBl5FJP6kdQhB1lbBNY
gILMFKunGdTBAl15IXpySNJlfl5hRZ8ae7UgOqLvzKztKqzzz+pvKIDfcQpO4nMM
VTXeXqEm5JUBmPH7hbiM3tcKRsh1FADalmMU3vZYIvKd9CkNSlT1cdGo2f8ZQ9LX
2unBmbxWE3sfCy5FgGfld8m5ZqpZBr3O3T0m8LSNc6z9hcBlwDChlFfbsUhf9fJA
8z0PLJckxHECrRoibUQZ4hr8kPhBGxdtwM6rE4wxbSIo0Qf3qG3riLzBK7xZfeZJ
nftctWIa6fDqFGJURlQwPULxvlJjp93Auo/4N0JjslVuloUhlK3+cxFTS3r8Z+KW
3kksgu51Ku+zpEhwQd/WVavAv37AGGK5ngaqTbuaRRMSOc+TrldgotdksWX6HRDS
gF7zfTD6hzpzYGoZchO8ExhxssGbz3QfaZHCUPeCEcoFf79MMuQOEjDh7aB3HRe5
+chb7AIYnQlIwdTFPlsvGihDMVlJTJoyuZpR7uVhLha6tUcG+sawuN3p2o4kEFzt
Kd7Ry+csv1m10Ov454HCXzZmOqJxMFO3ieR/d5FeWrw0vcTos93G5HepIbPkWkNS
uU3ysBpOIsn+68lzWHjQe8mKDZgSNKNyRrv0b52reVUbLMTHyhgDIbyiUCLQeezE
rI5pnFn+Pz4NG7ou+9Hn/dbO+h4h91fZ/WXmzcvS7sQ4+ke3lqxTfkV1OqLnACnH
NRX35qK5SMXb/XAfdbmek2XYfai7zXSOyaYoQpdFwxms0cOqi1f+ZjBgDC99J/Ps
OXH0u/kXvsXLeYRZSoautGKoxNBQzzJyI3ayGXeTKp40yPQVyP8jrH4lxqwI80F+
OFv8GU2tyPdGZmkmyMrnbeXV4yv0xfczdn2LrpQdShBZE3wS2M+x92RlzzpbM/d0
MRXsFLmupnqeyMb1iiXWjF/XwWRUQTCtRX238MV4gQb1GS3LqIJfsTKm2f52jfxT
EBslN/JZ6Wb6Pr1AgCSUX9UITqlPUjsvIUJJdAFcoGxB/SapdVhArAExFYF4hCEA
IITnBsJF586PF1x5r1idtSuaKkNxOZVfEXG1SUqubXOGMrQIN/fu/55cp/jqzTsu
QfqQFri8DZBpkwkWy4Bp6AialPtWWTVJddtUs7r3GXfTV/lIqcEl/aeJZyBRwS3R
8USgtrP+QcFlFj/4jDPeVa6cK2ayj7MsmSryL7vLtPF8t4KAw3D+RSaHMw5rpZGf
Hw20nOS3S8IBlbgwQ/GZ4cSJZjkrpOOu4eJ9EkPRp6/j1O2IfuNNJZIesodcrQHL
4Tf7drB2TTr/zVnGOc/pYnirNWJehKvABj97iIiN8M9HFmnp8WGh1Xlfw4QT6QJL
Cy4W7HhUz+ePL/pPs/tYWQRX00xE59frb3y4IUrDeTUesJ28F7IAZ4YzeQCnbNs9
f2bJer1aSUJxcj7Gy3dE6P0mj8lbbEva6dx/yh8buFjjHK9HsUfgjHkLLapnsyhS
XdQ6ObEIAb3C/EFGg3Ohfy9YZAgtp6trP18WPgOhwBRANidjQt6rhabvUGf9tRF+
dVqdoGVdWyhUf4McXYsmvw==
`protect END_PROTECTED
