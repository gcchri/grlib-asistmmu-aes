`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J7RcVFaFZvXRcyNUjP6KXvYEg1KLfuA0s5lJTM11yzuXxT3svzhbaYvr9zfViaY+
wqn4mragLjH96tMF+cGgbfMRE16Uj5jEI4QemtDY1732gPocoU9Ty6UajvM0ZmM5
0kHKduOmj2z6dW8XnDRGNw5EvSen2ERp4Vt09rNnQNaZVX5XCDx1uBKJm/xR6BH2
gPLLDvJj/vVmT3vzr9kAhlXSTiAkM63HN2DZgX7tQ1gzTUWVX+uwHP+kGfwqIz05
StmsvxE+LCQBpvVYXBHGSgGSyO9JOEvL5neG2W45269/0vGNJxXX3HGu/3NpfwLU
hftjGhhLVni95XjfpHkb8w4TVwBqx3ZB2KpZfVVSUsjohmEYKVzAiVN7voLPWWuc
`protect END_PROTECTED
