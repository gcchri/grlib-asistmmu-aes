`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SYaI/HknkltJS3BPn7fc3UBvso31Av/D2PcAkHIFPKmry9dC2hUJ7X27joWisVk5
ElBbKYefhMoMdhbSZ3VK1fZorPWolZrK2PSPpihw6CsWHX4L79FUWRAQAGxFEixj
fmBYJu2cq0gvRZl5C2/WpTKk6EMnZLAPRKql20vyGz0UuCyW8Mm9I6XPN8EybrD7
tUl+9pX7wGfUKuATC8hR0mkCBjHaFMvhcEZTch13sjQjwN9Jbvnzoen/K7Sv6WKZ
Tww+Moe50eeYjnl68YXc/jT1bLkDJVGQzY4iq7xhRRbst9a1ul7Y19EK7gXzVaG9
MaZy4pXiupjF4hrlQSU3nAn5/lc5CEoyBh4kv3aR8AjG0U7xG96PHN2/7CYL2vZI
p+ojjibOS8s7VN+XGdzMqtNCtNc6RhYpyUvhUFljAzfgPSEbX7HN39NLlj+Cwncc
FZER1Ft/q1XcKmGEMuVyUkZ9Fp70IM2o4djlBem33awMETaNDfHFLsxRTlZyqQbN
ymxKbzwsr+JOGFTEOz/M1iNSJLkTLP+XH7P3414lt1BOn2pANCnGRARNF42iO+wX
NDjqDgLL4d/wDlNWD3+tXShu53GZnkGXaic0NXcuNwckeIXLYL+VABnekIcHJ8nd
Ki4dOQ9tTB0AWQStHo8u0mnxTNR5z00gLRqwsOl9rjCzkHJjCJo09Gjxx4fAI+0S
cz4Ph9CLsMM/1NNerzsw5EkA6nBRBzvhxRP0JhA53U8o3pdPJvviXMI5Q/IGq3US
cVOfkhjeZhNnlCCLse+kJFG9c1CICA7fYPG8OBl5s+M5djpUszjnHUnAzSG+llZ2
CzcGAvGUk6Bi1NED+LCGtk1DWLNReyc+b/0Q7P97vCiS4GxH59tl2eHr9acquUJS
kMWbxHVgfLfeApLk4DoZTkaAb08AjiTM+zWp1wPuMMp5GW3vlCQguyW5uS/m3c4Q
xrWkfOfR/NHxIiwLABjO9p0EFVwj9Bvl+nZIhJdvhnCnRRQXL0OUBMqwSfahyTo5
wJfshuiPJ9VgGYQzMJ5iIh9IbG1VabSdfkSzZhsZSlHJwJtuzE9AdBMvoS9VA7Ee
T9i4eMp8v/12aag4MoGJoA4M+uJ4rN/vTSsZ+mbeILp51XTGyCd1xqhO6NDLAoKv
n2TCIvvy8746Fx1GIIl3iljB23qtX1WOKMBkJbi5PDVFblhqsASx2tjLZwA+ASca
wFeFyR4IyYrlJvlGHJ97+LaRXgf7ZB0UcFku1VDyuTzWc1HWFbe9DP4lsqEdcs/R
DRfs3js0L1ZPXXoBXScV2ckelv942IXULcyaTlgxZEdRDCaPPwi0i4765Nlv3D6N
US7N5ejmuSkq9SmbUP5e/aCwXrC108R6x89SLqxG/kHmqFk+7+1BSyHAuHc+sRdK
W/AqNU9uus2jR1AjmIn/mpTBHtLtM7LL/EsBRlEvqANRQsB62gmz8xeM+OXSNFFn
wvmaThON7zNVC5HO/A2ZAisCVKFz3Hbx6LSbO4hX17aq9Q36WcGRe2nNg1QQxKy8
Cb5sVhNti3q1k4WnZzJxIgNnQq+xXU78cjJnJ26wv+jXsZFIiNRr03jvBBMI34dA
40ZJKQcnMw5wchm7tI4CeyE1jZ6YTAkqdf2BCcxKNKEc6nUmZ5cimDAIfPOUAL+7
Hv0VYnRjfbjen/Ft3jf2rsP+58mGWWfgI2biY2th7sDtruwBvo1y/6fnICZ0QkhL
YTkgJtqpJ4siUW6SY/hJW26J657cmNOKRndNWOAxKE2aJ0mRX0hKxMA6cfc+lh5J
ZD1G0Ixezl9tI0hmHovd2kF/R8vssyBpVTmocBX2uq6tzU8sZsm+rki+r4UOa6n9
c+zyEqd4N79JDTzZ1wZjdpCn2P+7ysaLFxUsKPtpM03Q9yLT1mxYJKOVT/k9vk1L
x1bkd/MjDb1VFYexymnhkJEigSYLOWAdVJkR3uROUz6qu+lseDe6fz5tmxr9Fdf9
haSTGLMPrUGw+7SGxwn21wCyDQZZo/Qyz3LKsBxO3SvfdmJkDpn4gOjzBwVrGkgg
Y9pOWDnN2MKYv2XM/C82R5t39FhWxX1I1urovFLybhBK1r15C95aQOnGWwx6n1Lr
9fVwfOHEAF927Edlxn/c/vQ32x9g78BYmyFqTgdJgMpRoEBYVmtGmVitt4sUormR
glYjqz4R+VLEFAyNAlbTwwCpsDi4YC6c5+qqDCjji8gPrcvrAH8QadXGrLzPWWZG
UuuXquYPhpX9jUpLCBYAoyD9oucHGfaAcnq5OMwmKbwd9mWeigFcNLdfESmkDv0y
/beTKiBl5bFNpWWPeRJMn+sQFRShkRX2BUGjUht4J9FQ76WVKJmvlBv3CQqMSXjJ
6CrpFM8c1N9kRD3GVpa2zYq0Q5evpAS/eYoeYs0UFofn8VU3wtGSUNdSsKfsVfC5
ayL+LMOUZzPgK0btKyHQ5sHVI6wJnIJxAO5ecjQjnBH5LacHP2aSJGQMnEYzOc3h
+rUNrLmixdoj0rqXiuaqRMUL7Fe3ipqZGRVA+1Q+F76LA2QxsbIgNOXTT5cfW01y
F03nEy75P0cHXNvusHImJp8ZOg7GrlNzus83ijyeqpY7eeCgvYnMCVr0e/l+SdVi
xPun2F67WhWRKFIXA1+9xw==
`protect END_PROTECTED
