`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+NDatOsQSj2mwLdDByotoR6pzR3YKD/GSlBGCHoysA60xIWsxxyGTCE1c22TegZU
MoJ4Kmhsm0WRLfDM0RyuTSNHQYOdQC340d7nvozCBY+4nZrkuAVe77fujpQ2jYRQ
Yzru7OmU2CEobuJLXhQVmfM/h8jA+9PbHkMTAj2aotUXtdqE3BKNssFeYDfNSr41
Hlhk2cxplWw0HbZR1B03gcyz6IXpeLq1PSTKyHjYlmcBMTjt+GUomnfgu/qUMTsv
L8xS5QIlYBGVlC4rQdD7NYAEXwTPT4qOgBk9G+izSVqUCnRa7vh5QylgXKY2U9o+
uxByoBu0la8kZeNFKDPhAN7KpFKQ5mP3CY5AgIXNy58PFasHjj8DsTUpRdFba71m
dD4HwVYcBZ6kyU0WXQV+QbxRv5xH46v4t+DjuSpCYcSqk4zwbmVl5gtaFqfXZUto
kYcJPoHjmiEYpU/ocvYtTaK4dfl4uU0h9igjW3+RVzHIRcuk/8+FFbLHTeSxtLoU
MqjP6tqnJnOqjS+mLwy6hb4PjT2LiCLvaWqW7JiyS20hUmw/WKczDoPFXtrr2AB9
MgHpYwmJHyTv5SVwiHJRmv16Stsi7hc+ke0yKiSQHU1AH7hI/7q9xxdZEA1A6MbC
auxS432ERQqleMVNbtipZzW6Qdn9oupFNILGKbPqKpcPAxeZtIn++eGzImQUHWNz
udh1yz4XcW/Ed9uKOeJfCVmClmxbZYh6PVyXXSu1AnejkF4x/KvJ7Xv+4ONRb+Vb
xirocn92NxHyYFEmAoZjw7inskcGjuKEDHYLKXdrvvapKoH/3Ztls4RCNXeZY36X
0MMnmTq2F2hCEV3rJusobVXdYN5ESzSn8fijeEe2erAlWqmDZoxyGgbHD9fiiI70
KH9rmekZxqyJJ6tunZRZ0g==
`protect END_PROTECTED
