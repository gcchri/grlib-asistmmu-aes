`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Iy/ge2au4z/t0leNGVDs22zPT96ULPOR+OuSt5YY5847xiyw+GclNEPmTaoDJ6d
ew6DllmefOBD+wa84eiOkH/onlne93sGP+XbbftAk/AMhQKWWOk/vryawh1/80iJ
7CTzKWnwt5DB4gzPKnhfp92nFF39h3rLfIMBW9uJlnf2qhSi7/w8cE8xFjyAQ7KJ
CPFs24Hqy4NfSnbw/YN0Q7IFOPO8eZyYZV6E1lL8ESXQ73tAe3cj8/gyyIiyTRwa
k4MAeG3kcEX35xIVB9x4DbaJPAMbfFVbQfhGhHglQOTKZXYsOPmPTKLbPq0KjDD7
gd+o3tLIa1rUlrnPGjwuNz4eXR1b6VwM4ydvwK9H/5pkAENOcmiBowR2LIMRmgfJ
hBl7m5hT7Q4zbW8SOEt+w1FRc6ZWLcCSIRA6Bvh5ydfMR6YggLfg4g2HEePnb4vE
0YURuj8ApADqKRNhrRfo5CPVGDrbDfJDLVceJWMbI8g4oddOqZfWObid+Bp/DfLa
j03hxUV4GZmzOiqUiMm1s7uB70z6VRP8wPa7AVvrk1ZCB0Km+oPhiOAKzjVUuqdR
aUaBJyGbI2fieDYOSoqhI0dk2Uku0VP98R8hkbwZmi3E054ZpObcw+peTZ/8FeK7
P/XoD1Wte3SAEfSslS7OYw==
`protect END_PROTECTED
