`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VG07KmPa+h82Jep1EkDzsp9zH/wh1DurShoJacGRDYXQQYr4VtLmFDd+B24RxdG3
9BSqjB5CHNCbZP6N3SDqoFsp/QymX1PtY53SZnGfimU0T6zwsyA1KHJXcTsW7V0h
0FoNm2D+BebZjuWmkEkjsDQ1U7dH0i6Mss/4+aZVsBSBqa4qneGzZI6WpsPFkepi
PPyxPzh6OOk9g/Y4vnn4UjoErzDMulyi4X7RFH5Ary1URjpZa4thm6ZTzQE4rwDt
qQiih9OPKH9uYuuolD5swmTuLsFkXn4Pjn0sH1BkWGRIQphjG8n+D12wR3MlpRtb
A1q8F2gbW5T4ZHLpj0khqQ+z3nAehNXBsayy2qE4cJGhm5TbeAMN+ZLu9qqO8cS1
gQxVu7asWveVFfc9lcf184bKYJ5bs+24wTPP+Ibc8Bgyq76XQq+M1Gn5I9mMUIDZ
0pBdZFBpmCxd78G4W9d5Qb34EBY+wzYLay0rZsciRQtPQrcDBpLQxVYkh/Y2O6Ob
/7GPft9KQo/+0m1J1drY4znxwFfsSbySDMF/Bb2DDgEbG0e5O36qdi5NmJ1mb/V1
clwAOK2mVmghbDuKuNVFjfBAlG35tElO60dFe2jfa0E=
`protect END_PROTECTED
