`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L9caypx3k/m1kKk/jBQVsfGQxTNDutawpciGNsrYF4gc9JrxIwHiGI+2K6edIo1p
WBTXP8nkF6k4l8DoyknGX+B/aVDRWr91dkH4xPD/MTgLO9xXlLbwW95aQ/Mo0+7L
UfhHO+07AxCoycLflkIYqp6uEFv9B5USz7YN03qw71lMtm19V64Gte8SvTeF/YB9
ab4PpMMPAw+ut25mIDx9fIDskWgin67nABfn7xvnqVY674Kil0o9FpyXF/U8ZSe+
KX9F98XrNy661wXw2PkXNQzcx51GMMDIPJlUpTPf9mk=
`protect END_PROTECTED
