`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PzWU6ST1MhUGa6IrWrO+2jlT5lS7petQLi5pblBAlT4jp/iRlYW7YQ5jFH8JC72W
z5zvjza4fLGBvKt9jUQc0MigPgnO4/2ao1WImcfAeiKWQJ3AH549MuFuI2rmWzEo
4mPcBU6QXl1ovaszL/9SvGPoiYX3VNgKW+6ouN6YWtFtCBUw8A9lEHMTkG1/PTRJ
toevPzu9nih61Af6fAvc+LX5gBZzNaY3emmiuudCxpB/ci7fQVs9Ka2JuY1x7muG
xaQOiauRTAVaROF3DmlK+5bNa4+/bK+MgoXgIjc8L1HT01foazlTuYddQ6NXWYCp
bSBhuYzOHbvyoI/Y1PtNXPzHxdwhDdr3yViAtMjsKX8GxGrXGAdckmZDs2Q/iAsv
QAdTx3S7xfMGnbpAxY7Vt26zTyXCHmO2QFgtn0dluzqZa4G4IkJZqrW6Ti7FUekp
EJFHhSbDTYSCCqaeDT2fbyryB9AompmriQ/h9IOjGjeC4ae2cULSy9Y6l9G6E+D2
TnzYfLzVKkZ/fD6mdiQqMhV6AlZQ1uKTuFip3h9yqiPyUMAkXDOuH5YWTXaf7nRB
Rif/wPdPCO7MWRv6LiuRCqW0eKNyKWeIHZN2YALYwqzsmHpAZF7Y4b423VOsW1G9
OvSCAzvdH76wR7WnWu8v0hABq14E+y4uxR9YVrqELHfMz9O4kC1iotgjRb6A1Fio
fwXkGWWldFkbW0/q4d55XK0XogAXTS/FyDTo/fyLbSf9jp3JkDhXfsm8Y5w8Oxkd
xNBtl2MYE8jO3uUp0YcYDiHC/yCb9fDVhdO0MSRLjQjThXRrmQDo538+KRKF9NmH
MreOfOMZyIBl4sSxmgMxZ1g4YlNtAgvK0MkbMXQKvjY=
`protect END_PROTECTED
