`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YAl2itQmnVjlP8oSWzYSy+vwrNtRqjDiMIK5VdUHA8c4pO28tnnyouKsVuc7ndd2
STZTsDtQxaWiYDrm5uuSgqsRL8x9FL71EqqeqR0mb/0IB6Guv4N8CwvnCwRwvJW2
5NEPg0Dyn9d2wLUHXUkT3CqyMOkeigsDoM/fFzPLncf/AiXg579HjH1crxXHSRjk
eU3cTaFCu4aPP28Okwsrw0tM6nj24nC8SdjZejaywUBn6TBN6fDBZHKoDRpy6ALQ
Ag2urgrnZV65Npi3AL9zM9GyZrjdY+sPXIOmF9N6/dA=
`protect END_PROTECTED
