`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HwKxKU9BGBFuL5Onw61uXnBp4FLuvIhCH7OGZVWKUOtR2hnCqKoVXsFhh2FIPrRE
gpO529HVIl6uIx1eC0ZF+g29/+Kbtq+RipJwxs8I4eNJZPDIrZLc8CkTAJqojYeE
wVrRg4SXbxxEZdEswlgT8dtGbUhP+zwYMNKwVMJ/HZ214s37eOQTZr0IZBc60TPS
dhtbojtlCl1p+kxBdRqL0a2+bwGVJpxCaDiCFwdVq7487hvcP9eXE8yKuufK2hP2
FAlIMsvyFbq6HX8oNwlgQjshL9oAkvFlGm9YWJrf7yM=
`protect END_PROTECTED
