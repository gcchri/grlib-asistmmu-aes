`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tTb5JnJIhY6DN/ryMxgCWGcJRqu7wQT7oyMwsxCK19vcJp65qdhQ7xPiwAenGOT3
NZpG+8E0X9EBfzrpIEwABVIw/E8inY06U5g6DU5s97RyvUOTSYS8wkjqnPmTXJaw
eDG3R7AQ3Vch6g+XMFv/f9MLQ/cnLcn6FrDIsatJithGAlcpaGQwE1jgSAXppdls
L/Bl4JerLpJN7T2Rb3O7FPYGDN2GGN6fso3yZO8OHkKEquL9Rs9BVM6Z5n2uj7+r
jY/1wz7XE+Qv49Zxk5RmsKSZNVpwW39yBy5RWhsChEnaN6acDTQsgptMDreR0q+3
nsneHhybwuuCrePayAPAvD50H+uXS+ohN9IKRyhDCbVWjGG9SHB7pB6llHC0aDwY
f0Ob+zk2P1ftaKLudJvleMK1EMp6jj8UmDnp4vx8yT/t8Dvt+axSYX52yi8rSwIk
9w9qfreuExnW0Swdz8pgUt/GDInNB7mhrBIwcXZ//tC0joYIYXxVBZCxD/2Gzytp
bsFEtIYm2rEwoB2xSzeAKknLLgy3bawaJmn2SvtQ8obiC9eyQhgtMqkwjTCXtVBg
ZSCT9Oke0k8lnfMxN8LNWSczJFbakd0YoGHMR9wVN4ji1NExcq8/Y98rIsyQwbw+
uT6bsZpxN2pEBvddIibqpQSeSPhycHaHW7KU7QWKxzqE2u16YDs2dTU/YOolBWln
3QHECIUn7uyYU4/sxIRzE9kDrUYaCdVRAXPMPmROO/Vgv1/taAhUIr+/J+SjEaRs
aq9A2hSH7iT/tRFrdzo0XBnkqj3mXovzxTC9mND4c05S1tXh8+LLvPs3DdPH2mlc
3b0cx6bLQDS/AfvDRZm3Vzrdmk9NtAIZjeaKJwvpFxqXs5UCz6HLkn6t/E38dALh
0JCBKo2BfkPqTzJ8YCVOYtY6Buu67rxhyB9V8i907MkipGvMs2wKqemX3h2yJ060
YhUmn8f92+BjyUVbVEkAhsRGH1XKq3cRzd4QDRPEUAZm0h6vv42W9X5K3EHvlb7+
MJwvI5TJAMdxRSOVX+jdZ1gJT9yGpadpV+tMLZs5v21iqmVgbfke+nalwy2KM6gh
if4iXyAyCoGrSKRQjMRr8ipF1H7WGxDv138DEt8AL2q1+QTrKR0UMwJOzvs7CBUW
osyT4inVFWYURRa73VT5wtljT7t/4pWJw4mRTK9lK9dlZe1osIhk3ovUtrcTms5y
ve6xZpzxtWBMMIIeylqkE/1LbpVtvZrW/4Js+WSGL6UFf6avD0Si4w/AQIVyKPP7
D/V2/qS9D0HOpSNTX8VJ8B0Y3jgD87q+lVhpPXN++vtxY0adzcg17mAEt0VnXdOj
Cv+2qLn/UTY3kvCS0JiFnZUkboBfUWpz0WpJUwF6g7og73mK2qFss3udLtJCtAcn
nXe27HbhwEYFBRlF0gJ5LmuTRYm8CUn5kWA7l0bImpWqHrtsBtnN5RzHGrka0YEE
rsi4fg4i/QwgoaPwe8nZZW1mQT69ZSQ5Zz6eG2PyMAnH2sMxS+TrkbFI2RlK2KDi
RpPccbU3TY6WUK85w4zESI4oPJeWbklilW3karOikBScdwk14ATtEC3v65s3z7ML
wBUA+m6cRyOZw3uH/pmdn2RIaANgBHjvp6o96E4XhpzKIbi0matFQEgExXa7T59t
UDytAYF62fvWYdrnEq/7oeL2uObk/3WHSKRwyHpd7f2r52kfRL2bu/P3wjIXhdyC
JpTQYgOQiw+UByjQPVvz1BPXX53sZDZ78jg/EtpVfqDnBWr2sLjjHHglOJVUBmCx
+wiSNGZ4GvsXUCPvcFG+tSod0TdUW4ezo1g44EUNKMejwMMDT3LdOFU5bsCQfFlp
f+Aucv86nkR5RJErihK0iNLlrvYJr3vvu3nr6hVpCJtRTkiwQMrxQ4XYCh2rxV/P
CYvKBIGIgyV7rsty/aL0HfHhj2qq6GRDxEZM1H3dXDrzciWdWC/sPXxSvwOczLOb
DLv4Bp0rOhjwtt65hdaDYg==
`protect END_PROTECTED
