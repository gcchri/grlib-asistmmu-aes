`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9cRQLwPk1wxVptArZzJDTS/yurK47aWWLWF8DCKG3wXXbt3DUMcYPLTZJZlcG9u7
YqX2KIGSnqmL11Yw+vpE1uo3fouXV3uwqggsY3HdxPro22bMXNXgpWhd792P8Ffk
zCWMFWR9ivOnk/fqc085NMCPUVGDs6hukNACQzT761g1j3CePaRT9Eum2RllWMNU
4l0lPRF7dkgcqQ4tWlaz5zuMAh2tcHopfKIz4wsEZ80W0df6PZ6yKAx2pqkn4vQG
eIJwNPAsX0fXMU2u+QTsVKVkxGCNBgUDzlqYp9fGizIirLdE8uG8J0AlRYV2mI67
uHg7MWFCo7uzIpHDSVs/YufGpV03AflqaQwV9lb9jNi6xPknKz5bley6lfRjbwyJ
`protect END_PROTECTED
