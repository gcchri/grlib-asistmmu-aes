`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6oFYX1TqI3yEoO0pVu4PRqmtD2nU8qDp0mjPUDxKWAlDtoHcb/dAimA0eYuqB54x
Yw/+uS872wSicPHC2CL0ZYR9SkpxydyJQwo4v5qzKzv4Sf6D+eBinVA9CAiJN9J1
1IQ+4aOvEh0qXHK+kz3oUsdzklATGF60CoNQTcpBIIywWGWvZrM88nCYMzJhiDpk
yy7zNyV+Fm8FJPkgDxSQhGP9x1qvIwjJE03a3S1sJPblSaHJlcic/FUu8GPLG6ad
MFnEw3J0cx9e6f/S7EJKq5aVoeZIucq/h/5aieZgvObXCLBpBXj05CXH3b7eMHlC
/j83eyogHxPj0POtjCqo3LIXjPObGr31VM/nWdKIUBonL6wQPpbmOrA7KvjydKXd
Hu+CpUCE7r4/wuyPdAfhDCdTeLL62ZDt88+I7Q4+AWI/jBnbLe5YWaEXmTOugv+F
hi3dGuTTJynio3zev5hAvw==
`protect END_PROTECTED
