`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GMCq/NSj/q447xXmMZUiTXJk+SSDx+icn0v7/v1yF7BA5UxiZoM6INMbWdBsy2JD
uxHdZXAyW0LeT2xpV88QEZrpdtsy4WnGQMyNtuVWQgvXgE1yzvrMZvNplAjD0mK0
4vQ2Rt3WI4vwrJdXhRn4TvIq8hOUheQ9ShsNaGb3NU02suXk3znClJQN+EBnlM5Z
lnYXMWGiQYNJ8zIivt20BCH6UCXx3IWsuO+IFFh7RWUsM921zsjvZw3Lc1GcLxtS
79bgDbMmQx81I8m4lKDTxAXEFKWHv4dJbRFgq1uiUcReAm1jgMBrJMZP3PAn4xQh
AoB/G+8d7anH2HnMN9SQSvJdJRX/jTaXp/yOjIiyf+xg9Sk+mYKdrvCnM+45VKTr
GfiE5f1bIxB4mVa1heLAkn+ElRKHGOO8MrueF34cUSg=
`protect END_PROTECTED
