`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z3iXF2TE3KnrmziFdlAByhyiqEfEBZr9Ck8D9cOfkdr7Y9Que3UbWYUl1owcYQVo
6csqRg6AcKQ0e2LRGXutsyNUWrxUAJj/Z7M+5AqhpODEYXEsvqQK+aC4ggLromrI
i7/HxgdVhjAPa3XJ5+AakjZJkPnU2u7mbuAGm8DsK9uQrnYRlJiUVMgls0ejJzA/
uvC6inBOjt2XQ0ifhOQAu6wY5fBPgeTX1mMWValb5L3weHVlIjMfLBmoUWVMeaM7
7JDEswr4ug5F7P9a85TeexGXlyaM6FNtLEzy3jXYeNbPv8fymju+MoK6zsUdLL19
HETRuheYFZ4IGU8o8in/yOHg8+kXt9UHDctfMWzuCKb6UsSYZJobcEnLS/LgYkGI
d8ZkNpZd1d6DtfB0Lk9BIUJdngX7HpImWzeaSHYEk5BawtnTJ/N0U7VcEBlWEZNv
`protect END_PROTECTED
