`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GP+h+onjpdAEa6N68BJNd0OdsZNXFabLGJH/Iza/LQYZh3TpgeVxkkZQk01IuXho
/SXDkZnY2TFurHXiqpH+C2Vt5unZ8OMI/q363mXP8gwkTaxU1fQs9rXXEzKra4uD
xdYnorHd2p/pE6gCti9J/h5/um0cgIrCwzdG2l1R4HFhCjBs4aFntQ0Ue9rfqp74
HZdcXLmknyF8U/Dpe1n7Bgifn3MbwAAwnGQaeDGYqdXVlvOujJq8k2RImJ5Ubdur
3DXrz7Wunziezl/zqq3fzq4edpxRbnus9GkO33O6aIECsTzIEWiC38YpVEByBzDV
buzlspEuTSDJDaOV7/BLof0IWJI1+KVhOESSGln9QJFqCMGS5R68w3kWLkBkQhs5
woBV1p+NPNs3h22GAw9XUWxF9ArSLZevHTEC1wqNATCyZjrRi5dErPYbrN6X/WjF
`protect END_PROTECTED
