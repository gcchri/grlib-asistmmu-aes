`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wC727G0uzo/QDdRvXO61JyEA0pNIkWoK73TZM9Hd0m6zrYgaW/3KDPle4/ZBhUow
zosdWZlkTDKeTk4wPWZ5rILs1ZCCXYmbUfU7rp1zyZFcxzlRqJWXnHvRoFNm/4IJ
AYEzlO5BMXI05FyAhQKhM1LmPj7osEY5mdIYHEFsIsMNjl7ufv3n0zmsS35JHgNe
JfM52b4hvUiM4v3uRuYAxfQt/e6syGAL4R4g/Cp+0+9/Tq+6umc7AJ5qcipEGUgr
WPh2smpVBnIWRZ2f4dnOn7KUzr4oV3W8gYH04Pq0oS2bVyDlr/35jDP1i1DhdNqs
p9RxjgOp/KTvm1gGkcJQTX0ZNeVYAHVA4nHeEahhw8HcMVqtwrKixQSmnEwZM5TI
ZuPOFeQ46F/3vavEtdYuVbxebXCEXF4IMusUlaeT2q0j/MWii+jDxA78qcFX2zkq
rkwjxJeoo+AHKwzaJhbi2cyEIuw0P7Le5ZnJ91dG3lc=
`protect END_PROTECTED
