`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sDwQ2mKTK6nStiWYE7snS5dr16USyn8esmXVxMR5B/1TkaeocqlGzYluq91OAgDt
g7cRd4yTu+ZdkyuGeBIaCrXKQQg2aQVjHFJTdxTyBgJ8r5/lqy3bEqMsGj8QNRLV
Ny46A4oT3xNGwlcz2BicFUwrS3mms0/nG/gQA+Uhq3cpi06TFmNNKr76INqg/W/w
aUnIaTRmVUTInve4BJ5RsycFKwnVRBeo1m5jBpmObOu9P2cLlZKT3r2mlLwTBrlm
y3jFDaHxHLxXUiHn3JRLGjd5Cvy2oJOXXdSqieBzKOk8aBAjB+aohtVQBkGnwdcw
Ka+YnybVQoKaC+Giilimo0m16WSvzSa9O+Xb+CVMywAhGX4IUn/dhwN2CsW6hydW
JBFLai1k0/6xkDdo0FCcArstHnxot7Bx1qZ0cEW/QHDYXl4FLRoFuYJ6N11aICue
OGOimFDBVWPK1T+Uy2Lhosf1E9m13w33S5mApwWFY8CCdWzcZB49jkEPNGkSKQEJ
yPZban5AhAG6xDRY0uH19eyUEAunl81GExsrStU6de8PaQCxM6sL2t47h93PMtk5
hxJPcoAHoHL2ZmR244zWhB6jpgGLgJoUGdd42KXw07p6g+OLHIfRQHsKAuxInbL5
Xavy61urZtYx1tqrJbGNGx8/6c+ZexzvJI3/qV6DvhDu+aPgmlNs1iqoYbCS77TJ
seU0fP1OkRGSAR/djhNPi9nrstS9tXM9ORJlWkaKnblBaNcOCXUdyF6wdA3VNrdP
fyU53mcWZhNXZWs6vp/NnDIthWJkPb8Xp0oO4vjENR4ar4p83M7+DBoDk7GmQkXz
`protect END_PROTECTED
