`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+LrqRDLkyAnpditXATpgDXnFz0wCq7grG0pAJilyzJk4SBY66kWgNHGT3yF5H+vf
GDfg3oKuBDwHPGD/Zd7LCoAvjHbv6Obocgq0GYDYTIBgT7IuO0AdjPC84TCaYJt9
pggADty/hFxWoAp0/uMxZTJETQP22hPjPaKDq2NXd22DBYruDLxC0fHk0y2RzpDH
i32vEZFQGapt6smD8/D8cYSt/L5sU0CpDhvrE5xkxKaXw7zCxwjqpYe29sT4Jfx0
+KQ6e1e3WySAlIJzdVx0iw==
`protect END_PROTECTED
