`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wnAXvWQTRkme98CK6z6ZqiDssF/IIYe8lbaQ6wazl/+xiIMn3Io1A78QfYmI3UCd
JcLuE5ZL2/cgQbIUX90MPc/aQh/7ONrIXE2UOAx5mWCbo9tGHZyPDqRnVSkVpmbq
O7djqgGVGuRDxY813u21U/kcF/Ro5Kx5YcHgVdPXX1S5HrsvvurhGFvJ8zvoEn0B
Ha31qi8l4CMITOW1QzJXnrnjQkyq1z0BrR+q55NDn2BdZoMMgMnKsDmQhRnqbmRd
jF51/kc7J/dedHKDZ5graoKCYxe2iTlp3JrvDFkv3XzANUN19yNcSXLsLgxpsZTI
EhqFSUEFUAwYGprvyfW6yEGkf5rILatVdzdQSaIq/rZgvX7KZh8NBDj5olTWOAiq
CAM/cbBh/9QIJaNKjqtL2eGLRVV3eXovsW+1xh3rBSvlv7qA4smMrbUoo/Nvsc+i
6ERp2WxWL/luKKfzVmE1lHCubYxjR8rpaeKmosIBh5yHGB9fiiIv2KapDojDcFHK
wOMEFkHefqId3ZlOctkjuaw+CchbQuG1Nphdp/E0MxE=
`protect END_PROTECTED
