`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/g5hDzyrTdupqgMUhY7h6qi5j93GWowc10Jk90bQ19j24ZVJJ4mbLnhQTNFN8AiQ
jVk6Kvfgh6zRfzGpDM421TpT5iHTlrQH/HwKhy8h9xSWMUKKalPS6VoYK4PFgbEY
uDOwt2bEFSKC78E9v7wbrpYyLAZrGZL0jFRLT71puH+YZdFJnf0DEg+RL0m0A99j
MFBtx3aVgZCKkFEXTYyYXyqBDy8RUsi73lVMhdBjnMJjWD2FoGUTMEAaDrxOoY7I
/8Cnot1Qr/i3pT5W9mWNiNGlRnXwjTwNef0tGyfd+3etUp64eME2ZUfM/BprO+Wt
ApQYGaFn/oEZ7mPqgxBrWg==
`protect END_PROTECTED
