`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LMeHXjCuHLbWL6uiZm8ywqXsLH83WGykG8t8dfXNzAJ84vOZdoZLUW4C3KOgGPjC
eDJX1j83/bSxugnAJDTr1/R+ziJ7hx+60zHAk2CK9P4Y0t+40gcc9U2bZCHfAeT1
OuSkeOCGl4Vn/DM6nBEWu6T/tAWuuldQv46aMvFaCUVAbGsvTYooMDe2CR+KmUpe
jKpPnauqQQxEVuEPi3A1Wgl828tEcYBxHCF3f8CUrdmXzWpmmEpFzLBmd0xCZ8zQ
eUByJLPfk/TD638SGMm9v7bx7kFp5PvEeK/sU8O7rsADyRtXfh33tYxLDByzOASX
av6P2MOl/BYf6SKEOKlSDWQOy2W02sHXYmAUznyhjULhzw+h2j+V/lYJ6L3iSFkd
YWitkeh/4+fGuEb1fuedH0ACkrKgw/7615GCE8EWtkLEUZgqPQ66SLNp1kCxnTcm
OWWm/ZZUTLZRxzfYL2xUIsigU92O3aDgpOCZuvDXRmwtnfQM7u1kezvEjVchtTuF
2QsdYK1gRPlRxHT5kh4gy9gjbRWg7J2nUztdiS65DkGiABQNGnDN95GpN4ykd0fT
rYUDwMS+i84k60PUVgEizjEAf9N18kTIqqc9/8UMbm1ytw72cCFa3jtvfu1CkRTK
emRsf7vo9wIh+oDcng3CC1K6cqg3hY5ERlZ0m38E7KMkfqQmk/fFhey3b1YAixfP
7C3ek7m7uWKmM2bK5zM45ZsIzSIQqFXCsWnwlO8raJse0JM47Rw4hAnfbN4pRKIW
fyxIYG2anGXBE0kRzhIKhBwgT41krXNVzvaOeVVCtPP1ge+2mtEvD+zMIdtlZkmj
CoiFknKC0m49mx2tOUGg+Crn69Ki5cfdTF5AeAVJKsbB7JzvpuA8poCubz7y0lIp
qNqTWa9+MWLZcyUoMxvBSW9CwIlbRSx515gdRu8mj9y9xbEfIeBtZWvOkaT1wiNj
qe8adw47TIQRptDFApFFncP4pkqUazHUk2HEQ/eogANStxplEkV3W0QbFdjw7P0r
X4mpNbtiL30IgDEynmL9nRtf65Rp3lCB56uTAKgecvoMBKu1XmBT1tTPco6ZhOBO
PJMstZTYUBCgwbfX16p9b2McO9+XlqW9F8HI+1X4kMYPQ9fsl7nxwS2ij+/cI4Md
Q4BeSS2oag3Hybocez78w2twCQ1nvb1/erqcdftnHALEDQXxGFW9hoaY4r7eqEXo
YHRXMoEGO1TbLMvBx+NshwT0BXevixa9AL/NdM4S8GLKcJ3Ck0kDsjx+aaeIwVKu
ninpaF0XFDDG0bvXzfC5qNaOK/SxqGEMsQiYR/fZYX5JwG+IWkHlIrwaD1p48UHI
zOfbNP3wSb1SGh5JpABd3ElKSvk/yVHeIyFNZCgMZ3hm9DedklJVR72DCaPP0GHe
ggbbvYUPMUrSzrP9Rp0vtcWZO6MdhJ3TwrWUd4Ihl0HF0/BjbbHIqWf7jeiMPOMZ
S02gJsc2FwqE1myr5Kte6hNtp6WsMU+PPciktFzXLjbCGz1av5+ADeaA7A/a6lX7
VsqhgcEKV+yVKV3BYS9q6ZKgMUXBS/VfOy/GDoZJRcBEhGIHDRT2/hHhJYyob5Z5
T1JlUFJXNZOwmfqpd5sg/FlhGxHD3Uz7C15ACkAE1Hbyp9zSSVKjUbTgDuS4TQK6
V97HYogQowoBq8G0Q9yOiHySaRAe3ASS7sjxLXsLvUJtA4qPlF8UoAEYMEAIu30L
TOkvLFxCK+fFy83tnZTLbMGLlqgh5ADHnaA0p/A9fs9+1PzZVvt71baIRGEiM0sh
/Ni8TWRGF4o9kNERPhATVKwqgpwqYQng3eeTT+zrjFhcFVOtdth4W7JV+zcgFttv
qjzxenIZ3tan+4RZUP2e+yEGKOIbSj0Z5q9HNbRMdMTLxJbLP0AtWwAuuYCjXseQ
aifM59I+IBz1rMy2fXZjWKy0q3IidmEnvyJP63cOK3mVYukuEvLtj6ji6DD8pUNq
ABYe6xK1Rm+jjgNCbouSXcL3ABNKw+3jmLtJfcRJLhM2oEEZFmUKOEsMM61ET9Ik
GtFmQ8vvQBz0eTeULbblFBIrMRdAjxuwPcglDen1V/CEaLAfk0TPY5SIRLnXN9d2
PyQLKccSGUnpDpujNl4x/eOpMXY64wldKYS3OjcFnkTzsgpvrqiFTIrbOLa4PaZg
xE10bq3cSaSX3C93VDjID1MrF/SmYx3pcuJ3lE2pijl9Eq/B/xrd4RwysRD1jUS1
Hfk7AMKvXax6AGLvQeHZ/ocs5zwxPGfDshafSY4RgGPppJipz/TfdJu+v4PhLL3w
AkNlwbbUF62xxsbjH7feKvzLpPDxDSekBM3xdIpSIZ0I83PMWP1bYT+qsdnA5H7J
6eJcf72iEmrhcGyDH0LY8jZobEUdeV+pXNu1WoxmOrY9xUCtgdzmhFiRtAZASJC6
6YxPwOgSa0cRnEvNeyXo3Ksa6m+hkIWA854nupyTE6rTmPE4A5VtsrNDOQXcioil
kf0wvzjVBpP0tbxjU0FInl/K9+gc37F5z5PBpMpankRG+0/w9TeONj2vmh5E7tlQ
gDVPe7QmnueD0occ4TnyP/48yXYi0HVlsUMZbySGxuljVk0+sXCpKHLj8PvVOb0g
m65lUz4NAXCRa0zsZb0PkM3qmpeEdfdPJs+m0J9bVeXIJQdMaRjF4yQj2qTZ63Ln
2Ez3hYOISgwknHgj2Hqyrj4tuw3ADSFvEyS27bgJQfvAby6ZbAdWI/g14wjQjJcC
tsw6z7TntZZiS4oYwIa94eIP804QJwMcRYgCkDoQnDHqj4kKdkx6HUHstTSQaTPd
7aFfMF+iUD+4W4UbDZ+k68zRqE22Y/Z0KgavhR3M2tlsRBGVzIWhou22TMgxjxht
c10cZC5nCwJhI9tEiZwg9pJYKlWZHw8KhBevvOH3J3wUwml3/TfkRR67xZmW1HnZ
BaIQvvdolv+6VMzBcGL2/Ib2+2B+Ku9oMi2ttscO+qYFYummczl0FWSV4S1gDMyd
zwPUBFnQA9af2hcMpjTS2++7SAkv7aaSe48ok/cmLEwBJfQLTtoglXWjivX8enE9
M/j9jzAxY/z1jJw0t5ky/MCofCj6RdsgYlBRBZJW6yyyIlkVseUKBYOZGLh9zlcC
HnWYQGZkOSOqbn7Xt4nmlIYL0vZ2XYY38QSCUBp79aaqTXr9hTzJzhE31pxvFGHv
uoeJ5Fp+kEFkQJN6LErFdsG+yQW/ESwcqr0vDKh3HwbefFcd5kwcv9i7dlt8IxUL
5zpAGjQgxL/DwbO8KBDhn1NwbgUOO0K3Q28pEMxPwKsd9M8X0j+jaIOzRNn8eioo
QdcVm6mukaCJVw+YBSYozXqR9AwuSCSs1dt168mdavFmq8O/D19xw9M8DFkmhfUk
arDXm6DYbPsmX/FUDzePi89qyc83gMjzv6thO3VV7Tlu80NgX0CT06gT1SCzE/bp
OJcAOYtGHq9WEiUqn2/FOyWJRt3gANkBPqloZNt0pnPZ2RebAKxuot3YE1/TF/Iz
br9shLgdIH0PbPP2JhOnra7eaxsrWynb3GKthh/dbbmaCvKgOMHLya1uMRvz4sjD
K0uC4cjnnf9KU6QCjyU94lko8BbcIqJW1Jceyp06S2+OdYpteqQ7Y4//5pbwWlDl
dNIYJ8Yp4kaoSVz1byy4q41lYE5dQZRNKK5P6IkLuAqO1mmPtEjagIzptc3lRNxK
74EsCKsMAWKTB2I8im2oWUHw2XrrJLxKkKfkN/F1co37ioL5vsugsgKYhyP5a1Jn
`protect END_PROTECTED
