`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
27pf4GHVt2A8MvrueQG070/7BvvdIlz05e4OkfI9Js0PP4w0HX9XxAK9Uqq8kmM5
b/Al25mlc2ZZyOwIkUN6vQOMaCOYq06DTyQBHwiN6c20as3uJWBH2CKnXhqzLwwF
BKUZv4r8LdL+hLl4JCfFFqmzbZyNYtR2g5Ai8CzcZ70lHcV1MVFBS4BIVooTmeSA
YQKKwEBVI6vZq9PYZaxMm8A84j/1OsUCUHwz4apilXHcn+kXxt3qimqqluouwfqH
Xm6z+S36YqZHMBJPasuM9knQVctSAyUcgmJ6jh71InNGLyZLj34rUFdBSJJd4dtU
cP3wNRoIepgwVtUw9fmhoetdgFjShvomzVyQ2nUjRfBSUfg7eh0k+UKuXXsbg5RT
7O5EYR1DifUAGXdUfkTDwYjAfpBbKHCGMlU9c6SvIDo=
`protect END_PROTECTED
