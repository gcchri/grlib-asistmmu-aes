`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ooGOai+wCwrXpT+KoJHIaNsTDJi4vQgq8kzxx0x6V8FnpwCQv3sIzfuGv5qYffFZ
fGbTK8ngMXrE8WCb5a3WsyPlgYX/vfXKObE1Jstf1iQQt5ctUf8BloKHh5WXV6Er
c+MGylC0G4SM0S9MBoQPH2d5349sb2LemT4hx4jZ8wtpGGc0HebmlTR1RelyvLPC
dU6OeLSb3mX5xj0AlkkF6wifhZtfa5GMuEV/Xo3EPSp1mOb80/c38JFBPKopBYfa
cwfAtRq+gLnrar9EKaCNtjguJwPqdmgu+K7gse8w0bMrnU8v06nzq+HqMkhwILGu
M63yaek8bGz1ZBdKQweJjSlUp1T3FeJBxzjgSiOx7uqYqWUdFnNgw09Kfig/Tgyz
buIQGP9vrYYAmKP90Duw2YsGh9lf41J+EN4pFlkgRD1KuIyFr0s+wYaefvTFxLMC
4jzopaVedKtaIdaqf6/CtHGnrNkTSW2jJXC61J6GTbNPba+q02CbHN17jOxz1/EU
g+s1KjZTOQ0CMy9B83we411JUaXe1D3Jf7IXdHQ+4J0WXzzPwtOJqN2LL77xioRE
Ym4iDr5jVaMqej1JUX31QA==
`protect END_PROTECTED
