`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AwOA/DdSoQ+zZoB87mtgn2S+ocjlsiPjU4oTz0CWYG5pVkZPFWToeM7zVXWR+wMi
K+o9JS+eNuJvFv9aduVCqQYnt0xpqj232jaT8Lzdz1A93Z/9e5zWCP/239q81pFe
eibss2rGhrTduIfXtIS8+G7W/wcMKXJ9NRMulSiAug0=
`protect END_PROTECTED
