`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
efuVu+52OwrrnzvW+GuNrucoDuEcFlH9EwHdPIlZgTPAGHbbQqP5IDqEZ0arUEvT
L4jf8bs8CfZOxFLCo/vRv3/1PZVjyug3QSaRI1nF1HSvaFrgvqwxC/++C496TsgU
053+1Xq82NLfBLeMWJLoZs24kzpN59t1SK0CdPH5D0ryl6Le7Ma4nTJdSve5lP6f
/Wa3ts1rKplXPYz8LX/INaWDxOXh/B6ChojthMjDMwy67JqBkCiMX01BghMfKyc8
liaZ8vZtIlDgai3C8BDXfzPT02i7n8detKzn0/ZchA18kteebW0JPoNp3ZAo+y36
E89mhL8qhvUi4t87tuWC3Y0VvjzQs+uMv/J7rAhOwF9kiKpabYvd2jVyo/2Uhkuz
9M9314jLM7q4aK9ROKi6u6WgAxPm1chsX5CfBevOj+nz4trRnB1uGlJcUimOSnb5
woJqlvWXVGHspZ+are0BdoazUb8Ik2k/9FEc1gr1Ip4=
`protect END_PROTECTED
