`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yOUZmgz7hNeaGHsvCdSDzKBoAQ8tX28ZHsrcQ8cFpEXqhUqfJQKwusG3S1iOLgXp
KVMPWe3JWq4PizekXiyQZf522hJPJ5q7FxeISve/CL2s5aWvjM4PXctpecl4ZSu8
5MVr+tmjcVoq2Iq18dN8xc9NfL8x8XqY0xY/w78gIuaWjQeA45oXjkmLI7KmmV0p
HrjzXQA+ZhBbYvZ5Yx7ECdiHKSVGj0tobYGkyL1lY1NzINyKeE5dgz6BORH8de6I
glmey+0M9ArFOppO9mHTuXm1Y9WYBbQnPOZbVxFB0ZH+cCUEl2PjLO7Oxx7cfWms
ovqnthl3FGXdgIFbUUKN9kiv/JF06Jq95Kfj7s6PI3Pu4P6NHBIVqRGIgLSDln9i
hI2fW1APiGEZZLUSLkuSpKS/aKnEJH464k9nW5PX21f1E8O3uKyVb2gckvYWihcg
`protect END_PROTECTED
