`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WPml3Gtt6NSs0bzWicZqVAJomQtubccU+sPoTPKM4L8kxL7Ehp8XvicnbLeYgqT4
v+zL4KRDgnFikZpA91jApn5E0UWQeV89m5YNQA1I64FiOM2mhvmXuPvNl1ERFKsj
/zd41MZ/uHec0f6+2qEd7k7SXzeCRvBItXoY/ezw/N97zni2T9CWiXkcSppd23M4
w15GQhgf4UN136WEPsgmIMSBXDSdUrLSH4glYP2ajzYK9T7tm6Jawm8XHJRu8fsz
zbdoZVAgkgnReH8TGCKRPQh09W+If/wuh1iBOrSaMQjNd570j1EFpTSY4dDVh5h4
ORVcKebmxk2bv8anU7BsADPbPvvGsYWxFiadBjv8y85htx1vcv5Onzn39CVCtsdQ
tTI7YU2QQtJGFuYOiu/S9Iaw3IxSEoQo3APbjwVi2aA7u7BglJWZVGhCEnpqcUBD
cnoWawRN/MwiGiecw2rFf5x1pJjtD27mwSyZrTPx2sH854aWT0vMPIyBxpBl/uNa
/5zHieNpSTbQT5ybNuMEDEezUZ4XH5N14ntxClapHUOtRS4PprPsNlfGlFiR3myg
/EXMFb82vVJ1OHGRJ9G1oQ==
`protect END_PROTECTED
