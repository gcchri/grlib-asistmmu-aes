`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hYb4hgn5hH4o8g1t8TUe3BkubsO4tTmvz+Zg7lyS+IC4qbbja4EhQuDUDekC61bZ
0EN0yyALLZTF9CFZNVMJkH5wuJ+esUmBrju2DdjVj4nVI/pTnGZd0JeP3zBIODgy
/kdQkXvuRuwD8i4YZsPiMczF7SP0pXCTM4xuD0L5c+W07uOaD/BjbkAXIUb4xa4X
HqKQTU8lck1GbfpQpTdZASkVFacs4N4SFSsjt/nm12jXWXuMJyjxVaR4tFeVZtAk
UR1BtK1IpY35Orne/1XkCV14YB8KY/bKs63Y/w2SmROjbMHMwrtgubRpOuaV/TyG
QOiaSKXzs/QGG0pEdX3z4yYXVKwaeXyHdWVKVcbhUX5Q4ODaUtjwlz/9WcJ16BqG
joMUBbXeTHghEm9knyR88HmhgSoJEJNuu2O470Q7dSo3RH3n7VhHEizZZky4DhNW
bMsGo7uIuK8U3w/VHrLzJnDWWJP8ZbG+NUd2KyBjB1ULrquiIsO8oLVB4MoDcg5W
A504JqhCLalJGQ2YzbH5fXSH43RFyfPYldZp1MCskiVi7j7qY1E3V/UdcqlSFCgY
N0EePSnk9WeZzYo3+uG8tQlO46aV0y3NGY4RY80ADUMWcRZX/EOjM6K2k6K2c8Pz
6glEDr0gygc12+UfSxLUDMQ9+j7QV/aFaUq+aCo/0hbyFfxufk6806dF+fTjQWa2
4hEWnRfMH6Ly3fcKv5emlnXJuVOaBSWEWWoZBkVXvppGzf4eaErQYPjGzGDV5F8n
dhGTAqeTACQegIFHk9Hz7/RKdVEaaCOJZT2nUApHnfdHWUnMhvjvk9OmYjmDcpDb
mhmS2AlDXTjx7RzuL8xgoog8lRxwYJON602cSF2gIsl9mSjKRLPlCwQHXhL9VJ7A
fML6Bbw7kSU5P11xXNefyjNcQDlrl9P5qnT30LUUoEUM/scNA/TTKpzYrYwkAKAb
bpnFC/nJ3ozDs/xbpsdfVKo0ItaPDD4R7cLgJS+6XLAcnEgzUMmc/C1k/5Y9h+jA
vLdGrs621/ZO2qLExfQsCuDsifr0g9V9eFPuTak4PEI=
`protect END_PROTECTED
