`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M6S1a1I3Kenrc5glmAELdCsMk43areYLn78VBvGcFYqCSrGfAseoCw1eWcj7uaQA
Lsk7bu6Xn9vJVoRuibi9hCAppGoNee+VLovG0IuRsztvwDtUcMIIBPY9H39N4ljl
o03k6+JAy07lbD017+TQ4GYYLg+RfgdaT2n5s3EwYqn2Gwy5dY891x/3OMw7CFxA
pCwDi0pyA+urKkAvAmFwOftpF+YnSyv5flE+w/5HhZwgsqL+HPhEMy4QJx9AiyCl
Uif8ZJBFOF1lGXkHRbEFO7ntwHD8UEiarY3RpJIwTijG6j3JGVeFWzuR32pC2yqF
U7EnY3GxR2lU/E0RlSFaxp+CV4J84W7D+fZvHUfpTNw9T7FnzzsqmVtCdpBOK27A
oqCvaaN6oTlCyta+BEcE6vF7VfWn9TQdDfuijiMyXP2EJqW73gv9JaWeymda6pOO
mUBuEqBzIPiKKkh4jMkaIUknjfmBVqj8ZgtwNpMlAabr88YdJelJT9ozlBVSgQiP
B5X1Dj3xvv/O7cX4XpKY9ES6gOklQnO8MYohdmADNXEcUAHh6ZrHfRkgInFPZeCk
qBKfxumoyPkogYGU3QDStWupapbLSMWdJVx8KwHuwUYr6Q775wzBh/wMyG5MWFev
7ejsZe4a5I2RgiBlLhyY4Zt9M1FFPKq1TpJGtJkWHG5A0J+7gqiqPgdUzkLGmBQs
4xNJBqHBlqCFhp5TW+I0EDWr/yp3olloCbxtnQgwl/3V6egt+VlQQ/mNkYzOWp+M
pvbGLHOs1/6jig6yu+MHXg==
`protect END_PROTECTED
