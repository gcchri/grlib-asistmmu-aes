`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BP1pCqaPnoVoOfkhf9TbBGbrMTv7g4ufYyYKMXDO8V4iK97CQNcYNt5fzF+r9SY0
BxaTrtCmjMmEA3YW3pftLUv6P4RSgRasAPGEqb8kT0daJSkKmZbAHq1765A7VEbi
NYZ6Jqcsvww49rjI8Bo9ifBEbhNhuhlUpLkIyy91DEu+wfG+0QUDVinIhUKakXKJ
VPCxJYJ79bnNtqwMk9Bs/QwidE3kpGAjiQ5m72yMkGCh0vZ4FicvULUVAmE/hTOc
UPdTP7Wo5R02Q2MNUH4Wm82yTnhw7NyvY9JjNBsTz4/pOoW8z4hFtFx4hV3Quf5U
N4nSJg4wUtqzt8fNlIWzMcPmYzumaO48h8DDx3HJbvJMTxilVO4iFrkkivx2694S
zBFysWENaQQv+nbRwUXUreT/AiD62huJqwJolaxXdO+1myisk8l65mz09TyHRcB3
FbyCCj8BM/nLj7LotTZe65FPP16ECN6Sstpn8kwTPpEWrJZGWPvfH/fxa/K1s8BH
wFC7Mqhrrwb/KmZpJGmfgkI0feQTnmTpBduK3ULOtSB+/9Ezpmp9BHacUJM7WNoc
rAv1q9mHtqcsG7thCnkPrcKUapTTpjJp+spOHrFgQwo=
`protect END_PROTECTED
