`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q3fkJ5KgS3TXgSCJDbd1UMPEqck2/oJTV7rCGhqwtiup7KoMFaHnyYK3HXwZXNBw
1lPHQU+Tel113YYSh/slr1sDMJp2MD1cnTr9hLu5FjgeNWVy0q29zwqmlfdAie/T
5IdL+ZB/I2wlks96O4fhKpRamDUEj0bz3iJxl3lLPeXpaR9anvRsuCdk369JZT5j
8fAbGY79pO4PlgUM3wagcWHw76cwYqV5ouwKVhV9HJlQ7HEVx/h2Vcv/IeY4xR3F
1PAfH1bDdS8tj87OT/OAUGlwHyuPodthxOk4Ou2K7Dqm9l60fQIiP3Bl7ZhrcTvL
vraCFD8A56XxeFxmsLG+n1Ymfr1TyJSsOoVLcxj+SNCw+CeStMf4h4Hm0XXwP0T3
l1FocAzI3JcK19nyuKuc2Q==
`protect END_PROTECTED
