`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dQe1TQ6Yab0HiHSA5m7exDmq76NTYMjVnOuCh4LzQnJbjv4Vj+swnMJo5VTUxF0Q
P9XXaWK6w2CkNQbcCPNBwTUzV1ZwCUH4NYlXQd+GAaZIjMciF6MZBLaAEWuDOGBx
dy3VHSqlJLVFuUg9ib0Gcrqxe63c1A0KYBz4wOcHfXz+mZo0rBflhq6B6/o6F6Gv
O2EXvl5brUdf9MlE+xUQbUlbTM02I5wEesugloG/NJDhSEOebkDbpDOL5W8wFTcx
KRvXwT9i2seFrBoDvWeq0T/ynaokO48xYTuBgLxc0YDZ3LT507Xi2eGGpiBOg7ir
0EFKN2L/iqd0MaEHMNQg0Q4O1oZZSzqh3SjM93uhJWYwn6lRLPminZveDUk2VjTo
XyzsgwVzD+fPzL6KspovghePvxzCy8IIboqTIAizEZLMVhy7YE7jXcjCCsxrwPG2
TFB4zGWy/587+CPSldRnjOfrhVpp9CdNBREedPMxEedGwPzAEao0qSnBe+MzfCuE
50qvcSe3m75PlRgXqqb7tQ==
`protect END_PROTECTED
