`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lwJSwLca0ulPWoKA3++AxgdX2yA/8P/NMDTikUx1GikyEf/ezEfsuTbOlb9in+DC
1a1mce6U3+aVDzPmxPeggeW+fP+kZwz35WMGZ6g3MMltcJElJxFDVuom9pewajNe
u58W2sigZcmjB0Woa64OD/3tie7sGsuFzSwfFJUt0rEdnxS2/RDaVfxGDnBs1giT
2dQz+t+jKpvZppV2+PJ0Bf/eOVk0CnOzCsLanazGUQD3iR4ZdGN2A4eaI4a9aV32
nMpfax6FGscVoeMLLEtQgpqEdQdt1k+tXwc1gglVbFgYzC1KKgXc6I0DBdbvuomE
RBlTT0UA+wqINGQuFoZ2moPelrlBhLeW/BiRPYF5HSZpxs7Pu76Zn/YVu5pJ0JTj
8iJUAH9Eefe/PQxA11D/vA48MipMSqWN0ssGu11r5XawIxv0W3pvwWmQ2qCroY/f
kGVZUzgd71VT4U4h3sdHuLfKcTVdSTkQxwv/uuyy2sh/1u8Br7GeGYe44HKToyAR
nBkzo375g+FrNmVdE6W1nj/rLpVUxL3cBj+tRK1MOF1UdAA9gN8uBcFdQmqSZXx8
ppTAUO9bufPYcxnjL71+Q5JuHaaWjRIJtT3iwr3mTDA=
`protect END_PROTECTED
