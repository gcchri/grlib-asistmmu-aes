`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nJxfIRvWVmQGbd0EAxCffIvC+LUws8qtvJ8xUW8/TNJtIPpAjhFWB5Qy2xHI18Z4
l/W0w0ghl9T1NDe4/Wqgm/xTBzwc+Wgj2liAlu5sEht5lMg2ocqlTOhM6UfXrCbS
VEbdR0xpR9j1bb8knFNCLy+hB/7PKZX1YAZOemvxzM9RvrIe5nd2x9Xbsp/GWhCv
GMVHOcHCAYxsFSsXWVkPAKuII5I6dEyo+5+7JypkJIXGuSuudVNxdoKJUHkVWChw
evNENjQjsy53VjmwhG+lNul94jAvAUGJR61538PVNEAadqgYvXOmsscijOvkxk6l
kSGiMNovOOQ1oRfYpMNXyc6e7+YPpfByqmsrdOuRgDzdVKppVevNXfQVYg45/2tG
1wXX3sE0OEbh3jTervOSPjzqs5tPR4jLG2o4Md9DezgipwBN8o2xAzJ8ieoVZhMf
6gJ0pMEjjWkLTmt7uUDKzP22So/qBm25L3F5696yw47ASb6SqYCVq8P6tMLfhUc0
VY5iI5hjWSOIGQMfy6Rn2xS3FlUI/a94lQPwNG9/7bgBgcdpiI4bgXm6GhgJGKef
2c9mE6f2c2CC+VkhUDZq5krhbSJBTqNiFSfPOkuitQ7KFi/7BsgHbF3U1xuSfjIg
pVHrEJOnVexRR0NhMvFTpnwcQ0snSdY5j8nO7g/GMmcL1FFqCGR2gwNe7Fgog8bo
UmbnD+SM39FAyeJkNWddeExw59DGBOmjcH7JR1OWDoK4QvO1Nep4XBwaF4T3d5od
vgTPiJLksmfBVVVyEePF6KsZIvK1doxuAHNBfespoEqY8kDTc/8EK4VQE9duLK2f
zzX9jUeFbdgLUT1u/NzUcqx9ZEJkK6/WSIuyeW4NQHXqoezzSUnYN0J7aScvyIVo
bjqYlqSQApYATzsCIMxLQFYc5V5D9hUzsoHjXLYbENIAg4QXCw64PL4CJh8uhMa2
PwF8TfEmdwpUqSqOSKgumk7fNbwyZ00dweZYXsNQ4cIC8T4DMUCl1clB81/DHDhR
iZMR4oGBDDKGSLIm3NnRPOY887gUJOsE9B4Vnajd3krmhg3TZXMRvdqNrZQBKHPA
DQh8lwVLlrSj2yTKMAftFsCNjsqZDOJamsgLdAFU4Z8f222bzqWSDpzYhSGF0Vdd
gUrj2Jn0Uwae85iBTz17IkrxgeidqxjaaCe7UZhXG7zkjPYkiRCmrmQVcIGMkkwU
0sGcoPjoOv3G3WVLx64UMqjoKIul+YiD/87Euxm87I0vFU37s04sqBfy1/Kk4gd3
YIBYI+7DAkdpeA/Hb77DIKRds/Vcbg0qDqxXfs0XsB+qt2uG8T8RFn+/1FQ0rb8r
/O0l9reXp4aafCUYeDkBuBMPIEqo0j4HItP5i3/flhgYvQ0eZhpm/SK9oqpBpSrM
goz9vd4gEq6nCx25Ijp1e28Un3mMCKeYF8aBU2ZUr1cx8xsHG5iTD9bgtvXiYF3G
n5fOMBffSDxDSb17NHwdW+OPAgyz5M/UZ9rmVSeTulzJZgv9SlyTwalm00V3AbFV
OHBP0kqJDy5A6StS/X2KQkafEGgsxzKVd6I54BiEzhzkZqUEmSUuWAzVd7MlegsV
7r3grOribsc1uLU3iv+0FI6B1eN566X4ET+BSpRlkNalSEj85TMbYl4GjDJoWg/M
5C/+uKmabY/t1x9mxHodfitrpQ8ywy5/XzNC4ivyl1tqRVuO8kNBO1bEE+/UXsd1
ZdlGtzagS4LrIRKQsHuNU+izSd7P55WHQIvwGpIH4VMKaj+Cj+BIQSXH8UX5284/
PQzHnuqXfxxvfp76wyNNx2JCeji3Lo5c2IsON0h+zXwjLMt1dIxH9pobnYr8xK6d
ndMdplIxF4VQCkTd9Q7bNuMateWmVNVjH1yylNuapOp8StWma2tEx+pqXD1ijSwn
eUobVes33X99gnVbhFumDm8STtPKm1Up9RPcdAezf7Mz+pollqv2vHhreUgqjr+9
NY1HBXrS1WtE9JGQ9Tja4Xi8ao9fDIIn6kKdRymO2X2XqcAH4oxiwdED7GsannIA
ZjtkCNlie/1DXN7q1aqgzgK865V+g6/Lz/Z3pMsfQzckyTvaKEyOsZ2UMYUusmbs
0XXcZaZLUCj9dhiV/ETx15DfmY200IVLgumtI0+BHPoj33zdM8qQ5Bt+f3bK8azr
gtOaxoOEvSr2NWdABW4X8Kovt1BEnYPF2X8R+DipjGJ6vm3mBUpCnZ0NjhLfS4LO
0Hyp/CAnTtQu9Qehr1nNSFAWS2CE94Ow37zdp5JTErOoggbIc3ewnRJ4OmD9J9kx
8BicsCvXn//4rLK2+iufDVXsrpuoU4Db7ZjJahvnNqqyjpZ4vX1CjEIgmzc4oArF
CREl/Kwg/hIWjcMsZRhLzs8KSpjYaPv0brqkGL0w9MzyzkCW5ehdMPMhZr/lFAPW
NalOTG0P/IAhnHIqEKQjFBjHOuYWCoHqqR3FfJ3pVLc9g1J+E4ezMtWvsl9ZGiGB
aAKTpY9cHwK+OifOhwyVtD72GMKLyAG7yqJEelCMBwpvo8z34bEHwDCjvcqQYplZ
lsIrDEttFYVlUQ3C3b6GTmvPsOG6ADjbNVSld3S6CzM5yKhxWvM+VL2sShqEFlWP
HxOqZ6nVSZ5lYdSqTW0uW4HbDKhrICnAcPAdAbKu64CiZQuWjA2H8eWPOzLFw3uA
+lDIK9+erMw8IOqnNcooHMP72wV198Yl08HWeM3cvKXeGU47J3gYBNZ7jJSTD038
bDHDE0NJLj6FfwEkBOp7M0V/EsJd2XOASGdCmG2wQoD886Q8uiMGv5r9Xwv7ZBhW
PDOfpIkjJs7EJCRrbAUtRdAVWBXC3dIFIuWxpJNsfkX2HeWficcWlP1fz1g+jmFs
gNRKS1Jqhsod+t7LYb5PE+D//NhJyPYZWe+tbS6jFwFaJVRy6Wd1EM5vL1p1XfLq
v503h7DQ/mvdIezepNzpDDm1F2Yd1f5yQTypLFkrPf8fviLUhMyPQUhgg8S1xU0Q
3/vIpVvz5r0ZV4PwEzvgJXvtxUlHXpNoufJ3MGcwadkngKEogLMX/I2HN6EVBYDC
uCq3zkegsZ8aw2XA5U1nvSsLViuPhzho6kXxqLPkazV2M7B5oUAkLN4bFSDvjzGo
KU4X2uB9WAHF85f3ykVBhuGMWfZTrUgX+dMX2qZelnemFBn5gyK4JHkJ662fRtpl
OYJ8In7CSyy6xLNaK4qotJdcoKqh8EuWkBEFxxYf4KVkSFcTNAp2Fj3LPCR40uVU
Ud7zi+v6WRDTa1YkNmoLaaa1jwQIEQFX8FaQEKsen/oAv2IeTimKPps5RqfVuWo2
vguZ0ng6NiLBOfTTmcWwGoF1H/A7eJrUAQSMgW5j7ib0DNo+1MVQvx2zLR5ISVFI
6K753kZC/cG61G+B9VTltIMD93IwOnHG/ae6Ocngs3TL3bENI5vM2ltBmyLEBskK
VDhJmZEnrnLJbQEp5hrCH/yEWlTKrguFJocnxjqJmIYVmUu6pLc8BwI7k+57KlOO
/jS41bPFjNcOPEsyybngRZ77D876wmFbqE5NW3J819JIk0xFbDEKwwSwEDHq3Gxi
d8rGMVOhPe0uwA76HvV6Ns5GGzt+E3TbGdUJ3rHjEH8TU/MbMy+m58DfkPj5VzjD
U3sEQc4L3BmBMFCyezxrtJnTkc6z2wCHVmqfmDprRPXgGYWkUxTXM6jiQqijQyh1
wNNPjJL+FR2vhYmf7bx7RmB9qWhvCULXQRBzdgH/NdhgyHo70HrC9xJtCpGHG4Tb
T61NANIxAQrCDGlV45EkfaNtPkxMQwLofXL2m0dOnQEIxEX532PrW54dhZ6ycdJV
A5WM8JVUMqlJpZNB8K9mJiXCFipvK7KKwccGul5VWCwNIy9No/pfkxi27VL5vEm1
B08zIxLID5DiWcBR5RPu404cpsReXgFgS5GIGHt+CtsvKpUolb7KLuPyuZUO60LC
YqydVideCEfVWO+LnnhvqGsjU0ImOQ2RGpdzx2ia0mnRgHfuV1S3RO140NKf+BVX
0EsNvW+O1sLHb+6FSqAjykegS7f1lfGPOkOj47ei6mbOwpnqfcvXC0oM4KDRsTA+
1I65vNWX65Sq3c+NrJv5GBLWc/y/z9kIY6xN7FStNyX1ibOC1KmCRJ1aYkJh95XS
LFu14cecADh5Gy4yp9nGjBzGqJGC61XQY95zzi9s3KYIkEGNEcdoX1iFTr/nUMC5
VtEjKQGCYzeqOsX1nUHTugbVWi5bIOqOjDjfT8QIM1kOeEgX/GigN1VLwEAOYg8D
uTXqpUYGCY4jB8OGpGHUc4E3e1uQlp5beDxgLyW69ftTVh1Y1NawJF4IvGHrm69B
dyNzoDfzy5mhQcL6gS2gEKmsjEE4m86CPUMgtUdl1SpV+FL3H/qRZdEhZJaxgfrL
M+FK3bvq0Sk0ZJNLDXvmChpw9PrvM7N3k2gVuIqIwABa7ETpKcrZ6mNbp1KRNXXG
bNSe9qizDdKg761i0a4WNSoSB7maE5o83NIar7mN4DrDIg2SF1XhtFVDaxPnMrnb
cSO44QIVP3ItqHVd4CeE+PzBNlsRFNsfDuA0iOod64z3GMoQRl/7TcpSZabwEEzo
2JeMTtbBB6D/spiFVK/Bm/5VUfIRE3/Aj3rWoLJOP/bLqfzsXt/y4dccqu00Nhyw
NkBX7oSjeoyRQNxT1SErWLG+Jo3JKkCbXr3nXeO2hVCEeeiZi2Yq/YhvHl4EFBtn
1LukSIw6qyS6imNKMCQs5wk2ew3yYn7ibj508huFfxR/ZydahcuAaNDGOmhywpKJ
4JpXCfK3M/joVZEXpvWS8ozIbjwyTiUMuGt0gfcaJit1B0mnsxBxchltL2sH0o1k
nJUATGVytyMGApZ0d8Okr4Oemusy9yEh56BQyY/gDppCzIJqKd/82/MsmJzpSDay
myzTZlSQooIsxOtfyWC40F815lKHPsZ6IU4whH9MPMAVB93sj9da/Rr08pBcmfN1
k+k9a5vb7fUFe0NXlR6SKBWvI4Wn9iET6q5/RC7D399M8ymHIp2P9e8GQoSywjjU
sEXxkOuGCM/ToutTYIY1LP/OwwFkvsqjrZN9XLsDMGLYTvr15t8J/SP5eMHBzEat
2FaUlBdCPPOzR4gXVeQaSoRDoPozTfNCWnyXBVNLZmz/1RuVABQtWAt9fvvl2lIG
O1X4CjOclLTgUNTswpHtbw7aCOuguX6kXDcpdhpI1T5vRhyJXniGstQuPfnkIXMF
beGOzYQ6by1vGstKE3niBYxkoDOW7WMqPR9/UX11/i5g2msE4O+RBhUrfrgdQKG4
kgB7dR9fkQswijh5JJx670zpb36edmTkVuSqonOSxg5ixf/vVPnjaJ/v8yjm3fvq
Tcb+8P3AaQKWtJUpiSEHBsVNK2NiwEo+m2Nwq+vDiFjj5FpXuC590f7KiHSfK6wi
gmKFrltsKm3eAxkAvIL5PUdEUUIF6hnrDSZan8h3e0Qs1r7uU3SUl3ySLncHZjWG
Ze4rgMQumRAZD4CmuIh2w6Mn7iFOkKgdJ4T6gjJQAQRHnXIRme1qdQ7wGIXPJKkY
ry7NnH4bbfJKSpuICwNkiC+P0bwmplZu8QZ+TuPplDzBy2Dy1mFLk68O2MvqYytj
kvzgDI9tCtJINir3Jv859Jla89mta5IMtb1TvV0LqGgh33W/VxxuJ9j+WuEvZzCO
rf+9bINf8Cp4XBAviGQmd26NtegQ94r8ct09qRmNBmE0xTgzR2OFGSFKgy9yuQNR
e72FNDLRx/m6UP6xMGYtHDDnR2RhX5PH6S6Pcs6mMDDGmZRMEIjs//SFg+Ud5TSK
FpHOshbAgKYD8qMTT7Z9/O2/gxu5/E79mPO0ZMWTILgKbE7BefVe+bHA4EMIkTj3
mfGxYHQFLlX/ZYPVfx9oELJgUnNj2TZtSvU5YhWS1RznIUAlOndN5LR1V1keljcP
WGGd+eGH0ZCpRBjROyOfncPrgmAJYPs+C4B3FtW5NfGQTmzRobm+iY6xjcpHMpl5
5gj7jLZhgUzNQQV7zyhV35xR3iGFsuihW1F29uD5GVF6mvSLtJHCKG1XbEgtVE8e
1walT2PL5wIhR3gA6Gnbqrt5uIViUdAgBeCS/jS79yUmwCno4qj1bgV0G6fPkR2C
3+/nhcineqc5fhW2d2bXqO6h6V9kj19h7aYhoYFdwmF4vXRwyt7zAHlnkyhBAR1U
uPZk6J3YJTzawe3n5cffb9rMOwIkAVPhMidLMQXVS7NfU5aBpoXspsEBc4IPpnnx
hw/0JHfNARz8b/1/Hwvj2Ws0fJXlhFjML0idTGcOz20QY/WATkBteo5p4noLK1jL
cpMZODR+5vyKgWfQHE1kkNuyn6+3g6FQKi4MveEU1VPv/6VI+RHj2rm9JFoLiiU8
WeONDQTbAj4BBvKs69LqO0nIvAvvJFGDG3Xrds9ZPdF92rLhx06Xm1QvjHvk+VT3
wFuGrVJkcvQZ7GRmjR1wa7x4wcQrHqzHsw+ox/mHm9ikA3cxcVTcsaTgLyVl/qTm
Kv78PqD27HziJPpQvhofl1VnBTEYuaztQu4z8OZqgZw1Yvo0yhtqQlhsrMH852YX
KU5L9HZWAB1VnVw83HKehRYCTQe5xNbbhhcbBwQRL/gvGuV3h2TZAx4ptzuko8Oz
bmzb6c+P7B+fiyVE+rqH7F4mXaya4e2EoW8lZJaVZ0JmU1BRXsjDBzC0OS9sPAKU
LcE4dGq7jVAMeq2bA+8LV72BWPOItyhpgONgCVAOoAsuLcYs5RBadpFWL+4BhQUc
01oDhsuWBUvkXy+1etSVI+gxUeJZS5lxbk21HEscJfYXRyGsnATaGo20vINoL9EN
sGtm+d5iGkCMLnxq6C7Z5WFRd/m8XOE2iLn802EovOt9xdHRG6qG9Nc2KxbrggZT
`protect END_PROTECTED
