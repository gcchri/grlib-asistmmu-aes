`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MIYCNZLDVDD2QAYkn6Reyx6VDKR0dGsTda2kKGMr7KIYFZYkRWpHlGVQWVmnwJBC
3RlIcl3nSuIsnPq/C8Ngj4GrWxK3Sav+RRcDGny8C0dEo4ESZZfbdE85YJauoxID
WLWNM9XSwaWkiNRZK0H3OMbnJ52I74SJLebvFG7ByMkFWnpKJdIltpLPYJfMEfxD
8TBMvjMyqzSYHp/Wc8LUrWmAVoTOjZ4sBRT8bVyFcAzHBHZFsDs/8sbbBFxLHUlc
rO8OJFVZvMP3QvvRgnJko1Vf9bBscu6e+ltDaoXPGjcWkheSu5YkHl1vPNHInQsu
la04yAFjBpDQtx4+a/S64zdQiZrO93LIuwbrVlC9akCtyNc67TClTw53vvewp0ez
QT6AGgKgv+a4Vxb1ip/uPKI+iqIu7olidervIOi78ixJmeM25UScgJ4ROcliBBjA
yTR+3cyiY+euONtlQ79ECFiuLuxP8Mle9ZaNUGLGdoxB/qeBh36sIObPt/rxNIGp
68MzEflHpzMe+KnWbfUBnCYQMFy6FKiZKSNyQlOSXgjiJRQs3TNAdk0GT2WTpYTc
qvhnk+CEbhBRnAXvNxX3V0FhoRb3HQhnmvTKYqQiit6MbTdRtG034pf3s0agIHvr
51ttc9o2Tw0+zYDEifrxI/Wf50NfZy5RUZLdg/ksiAdvCKyoQmXtz1Zf/komR78F
0Bdp6RXiazDAZTwFyIurLpzajA+OTZI+MYshbU6xwe2LmfgcpJoRzjGH4pa1EYN1
2vIz1hhER3SR1H2tOMccoJe99VI3zTfAJQc5Y7ZWEZ0YjG407Wq/u8VJl6vT6I1U
V8InzGG2d6W1Zkb4cFhRqD/8Z94aIi6HjA3t6Pa0mXXHNxa+xeqrzY3sEfwdDu0U
3hX4lIo+k5yshrtA4oCaUfb61HXoAVDLsKBnKa01sFHCKJPLJKhm3fWLSYNtPzJK
hyb+IUERBzuBTKcM7lREy3O3+EXrnbtWqUemMzxyPm4lyKCFo+zWUoK5i9/5VWPM
wrvQTYhM284OvNW5Babc8x/SleUnYi7U//UrF9dYXDU/nt1uheN9rq+ph5Kjm+Al
NW+l/914uKu92uKjllvz3IPo3NiEzM2b2c7CyBdYNzM=
`protect END_PROTECTED
