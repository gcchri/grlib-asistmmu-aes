`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8+PzRlKoFb44cOz2O9tBDYdLxms3P2n+2s2JnrIp94cDH4HtmDpknYcTbElsCV+L
poqe5w6g/BKs5QAnHVLp360fVLiAPLJVtHGjC51HxpXtvUX6T02WOYh3LTaPL2w5
/n7vvDIMGlZ+o4sAidAm2Dio24nQ/eRJqOhvkZDn+3sO1A8ycf2EcukO6K/srAqL
hdokIeESeBUxuW7TONvjzHWGGXpwNa6xSIRX3oym2A/ciEvFALELCzEneynAIl8o
eNU9Uc43nYBA+w+CORwATFfsDsce7g4CmjGJReCNQdhUlKXp+fqkHe2eo/3caTOJ
lxKKGfgou61s6xKzZpQvMlEHl3+2SlUwmby39dUYlIr8toze0PKA8+mC+YqoZyZH
CWfLQUI487XTpc1gA7VzHhhenGcHxAWEkvuNYlbgc06vnk6nYQymlpBtYdZc2yq3
2LUakdurOI6+D08WMrZI9IFcXjCM7UScsFFQ4QEX6tn3kKGAKqziS1tvEMTL94gP
GKrRv92qOvP4CVCXEeRXMEZHLl2arn78dx23J+V3hBahUTjtUDboKrYYJa+AuWwC
bxAGI8gVMZhWkh/vOA4upTwn6ToGG8SB9kl2moG8vPyJDhV/zRqXKsF/DGvR+/4S
dAMY0zybzXg2VoMkJUDLV/+Jn65n+YqCRE9Iwy/SDB2qxNM6B4Rej5RzATQdSaNr
8pSgq/+N3pdOeAN4PY350JotvfTQrsxEZ+XgkLgLFP5kX9SMaYtTwVEVTGB2XJlX
S62s4R9Vn4G2Q02Q8YcSDDcHXE4B7IFOhl4rknkW1+4Kwfnn2ftAEmEMXWOerGKi
lES3UunEYwY3vvtBwA2Jgb5Uh4UK80nOcoWQZtMDJ1MXOyndjzR/ZmWsKFMPbtTO
Luk0SMDmSVYUmxkIS+TD4Gl2b5ndFqo9hRdrNEBPWdiTmLRvfbG3y8i88G16Dg+O
VXcD7LDC1tiYChCEPk/ijVLJd4HE4Y8DCkTfRqQFp2nPprdZwYX9E2F+LpyuJdce
P4mCuBwA15EHPVDm49dc8QKFAa8XT/952u+n39l8PJSpFqbPF/6wV1ZjUyk9sA1X
lnRCDAPfgoCqV88A1TxYSJzEyJldlTkaSZYDHusuRWSSMJQ4h9FhUzXgAy4OEyic
toHauJ9AU4hkv1C0F/cZZCHH9xjdbmgEtxw3/qu5h8B/FXomikrlmJRFBn9MrFYl
9LGXiyNYZ4nl2tIx4tqQb62/WejsFWx1twTFJVp7Xk/nnaHDVDLEyQa2GQCQbSmZ
53Qa/yqhFznhoifxGxQuKUlX+LEr9UZU5U0Yaj6PdyhPVebdP/4rdqm6/nvXbPgc
Uc822OiOuKoNHEvQr3RtlKSraEg7qcKnFSQisMl+eHAQgEkPwHFLKqRO3yIhN5wa
IOUBLi/Op5sf6pGycyLJEL1VzEcFMvr5T51pANSCWLe7dP0ebvgL+KvKthK5iXVZ
mjSALSSZmWTEZCY7IlAkgduxRvNcU1tSavKbBqcWtOv/m7za+qxTL/cYC3QJ3/si
gI2W4laXMc48ec0fUiegDwx3QfXxMHLE1lCDLiv+ras9WOs84vq4vD9jK28ZlqLS
m7Xpuc8OZr81xIIiZvFQx4E8MTVYmFaC820UoGdVqPEpmgtDqhaApmNGmrpMFl54
3Q0FM93aWztQ8p6jdj+XzPVAcDLUfGWLuyCm9cC4UJQp8Nw9pzM4uUbgGLJ/nV4s
23P5wo1o7M0sZMw0sfRFjJxNu7qppYl0H2LwoSMAW6AhiCkkHWIDggiwW7IGda4D
Ej8pjrn6LdjF+SrFIdBi9ypXNE2ZujePbG6qs2ArP2P/wiote4VtaVmB39NQ9nhw
YVGTqkSxg42mnqDmM/GmAbEpIGIbNlnSOrNS11DVSYpP/tGz3BIPPC+hlAWA1C3S
7vjNX3vtBXg1DGH7jlUlZfdElQ5YGCybZDTKbYAcWbuUPwC3IXuTEQe3kZYQk8KM
J9bYhnE4IwHH8B/+F25M2b25XhApwY99mYkMv016dDUSsQDyHEDkg4iZFhtS6/4l
679fTVCW6SMw0fbgFvQn69aEEkAtNt/6+vGyRrdCWjfnLYAoYfvpAY/40A9caWH8
zGaGp8+tAAyCJWIc1nFQ2Db3c75XSHPIglbENYqrLcQfXA+FZA4bOT+Ie8Wa4O6O
U8OFoSoDkR0v2wSXdTDtHMfSOa8NHIlNvzhSF7DIkxFvzS/PTEj18NsJ5zMk7nAn
m7Mn/o7GVAIDnHP2NMVdF6y32Iai0nxFJmRV+7mOupbwr2hVJI9EWefQWq7jyoTp
u5164bre4K6EH0RPRQd1eIKmRtw/LFRoylo4McaoGsxqLWwSydlNMKC2QWkFW9Dw
yD8DIgO+tp7Xq9q16ozLa+NdYpfAmknB71R4HKEHNsq7PX86Be4fFqbPptfvSheq
UZehjCDxeKubfbYoiOE3g1pfeBS7mdmYsBDSj77Md0tzv5nqSSQFniXtQ3RmkiMW
PerVP7OV1oGOzuKTgODvD5DUTKieQLnMc358DLcKYGi1Jik2qldH5Wq/GNIrovuZ
elVwomVEzosoPbfEYdEq4F1hzvMvVXJqIuuIH9hvy7Bkfh+SHK1Zfo5XGA+fl2Ki
GLvx7tXVYX5eH2yiK3CrYyDN9iGsdxf7GFJuRx65zywx8mIu3s69ju8fleGikJu/
x23LL19uLzKf2lgZKuMPlHn9StO4tN+A16zoaWXZ3/7PbYQUljPTxGTthdQzXgKo
77DQkyWgNU6QLV/4RedTaIpjW/nWfABQ9kPN1DZIZol6kAvvE915OqqZUAq2dc6A
Sxs/Vaxn2i8ROsVxzR99Exn4L1ZTCN2wexTNtYx6JCqS4DwHycwUClBQPX+RC4uL
4V7tz+vtrsJQUa3329izFq7dEs2wwB9FMOdTUGPvPwzNceo+Mp/rARrWHP2SfsXV
OqQGgnL1GkToJ7eyZkNl0X5TbK9g2lRJuzbE6YJuEXoadlb80YChc9Vhqa3qJnJs
l4nVN/1Qy0k5XHxKdndBuup2f2vBj0dawRW07lPEHi/F5AEGWJimMDz1JFTkq2iO
hTD3BftyBV6TgmFA2qBCdr0Ftbc8nVas0nueKPAVliGB4KAqNuwdY/qxEaYj6Cp4
wW9YwRvGh+PgYOkwha8ypalKce3YcvPAyTJCXjzwK7rn/MNP3+J/tceYZUy5f9Vz
TgIwun1+mGf9/qPduJCWXCE5RmpVP9/oKmDWZSZqYZdQ3v5/IgvbOtihytlGj4N/
D2lcb1eJPEZZMvmNKDrc8G30fPSHMuOSUIAJ+MODr48D06GfCNiACV6MxIb7iS30
ancaQo77ERUpg/DEQvrupMbPMeCtlJZDcLWmN/V45IXlYY1aE4oDxKV/ObPUBuP9
59nTzn1Uqe6wQNu5niuNqm2N2n2JD3u/O8EHjqcjM39ROWNxQ/4BO/RsuBNHmEai
qmKUzWLhP+qVZ+ruOUyldZ80lmpnLEE7G+VsT9ADaIyes+9rZ762zvsFG4ku87SC
AjIj1pN4+/XcMDaOIHqvwQfYgGY7Mme7iQUhdj9VOaL5mByf6Tn5Yt+MAKyo4b6X
L+5V/coE2IR35aRm4qk8rdxmYzcjVDmWF/E/fbkC14VPVO3wkfo1BTBOpjktJUt6
gsVZPJFZ3b/AUxtNF4sxKg7Qz417LPSQdQXZ0ru8H5YcFB8K2YBrvOVQZB0CEdPj
b7jBOoSpJXtXlYDZBi8D07FJTqZNkjqRp80kjLHT+4SiCBO3pKAIxRQrjsV6ziFk
jxyLCw39sFyPlVaF+qX+Bwf/lb4WXxFk3k0MZjXPJrIHcsc0Extc8j3DPH8cZMBg
DSKarzOwUUQYTrMEJAoejoAl3p4TJhepl5yDQj42BfhoFAsd4c44rX7HIfauj7Qx
bFD7vDle4zGT4g9eg7nlEUBoZo6WkltTF0aBbcr5FEHiB52vAbz5PKWxCSXcQs2B
hyY2K5bgtgGZbxABkqs69KbMeuCYm/ojgdjT2q3f8fifAIjzEmjlcBI7ChDfq21q
pAAXPM4Jro+JtXvpmGk+n+5n3dy3ZIdpYswwvjngZAfHlnTI+GNBG8LBuB/6BFHx
hBzWCqc4dt3+EcKdefn4pmy42k4d0FH+0ai3o/uWuh3bG9lA9d5wJoN/yVBd5i2g
BeR68tIVmqECLFGIfqE9fdNUK677JynQj3a6lEmkeSCQ2nNJxQhm/dMBCj0xzdLY
TcUuZXtz8y0pC+Q5lyRUuzwdK34pfxPDSoD4t3DZlI+67AenWzo5djzKFf/uen8p
jqUKnYLBkVJYpxF1N6fUtKVQGq1wlqOS78vWOnjGbtf8XZ86y6k1EPNb/3yp7ilG
k7OfBXfwI6YIsTUBjHOO2yL34wEQItfab+Cks/no3VAKi5nLec3AG5/3PqD72TRm
aoK+j20MrqUT2S2TYCwsuytp3re61wjfCC6CokO8T2qH1GTRMfgBJ3D7OD7Ee/EV
/9qhCsCKfFmV9tc6lY8eGUtX3xN2bNfZFPI/AkECi2ddE+3TZYPiOu2Y5K/9cZWD
364AHEocYugeUxJt12Wv9H6UW2wDmcC9cAw/SrR9NJltEwpLjpTnyrkY+CPvJ4rn
M7wQ/IO+G8T0cPTmtR07oiSvdfy6K0CMhs598flbf5Eww+hdinLv3+dtHfMyOr9Z
PcGZXePkGNcDlf1ampr4nMyV/yMapYGwhMdaz3XGNhKkvmXNqm2k8Aj4FxcK7e6z
odFHOokuvjyRB09w0WFGDS5yfUb9QFscH4Y2Jng4jFfAARMpQPkW+HhOCBvMCKx1
OB3PjZaTfnBOTV+1QUStGXpn6D8UI7dNsCxB2yZ21X4UlJ8ZUukB7rFoLg1Qw7Fx
btX/lZFR5GAY461dyiuCy1n44w9bcccLYiShXnIcgk8Ug0UL5Q7t3PPg1rJfY961
8Z/QIeUi/ipX5rTFDoHPHcAo72DoBim3VVwKdEbwzxc3N6mlio0yYCfMeMdV4+rS
fSUu+ib7JIaSnwdHLIF4jWHFtkq1QnOqmCh2krdiM4vUwI/pWvn2MvuILetxOOPH
TIY2SaVj47qllmJLZ29meez7A0DeJpDe3Vw9p+6Jmn6215eG3wf2+k3pOdYzrBPj
a8CKTyUbWei6T0I3GG8gb4+iYy7oeu2ZLYELcrOAJM/KNH0SlgaOx5Hmg8qmOqP5
3dRAuXxdrJzKLc37IZpGhA04zs/htASi0+1Qh8eT1OLKPk3RiU4K1bfgwPWIzcmh
34E4HN0X75ItUaP8dMaFSlEta/vQZQyqQ/g/TUwRqsBgHexs/nd9iHq0Kw/C3lQO
lc5K6lyFeN7ALxI9lvnaNwT+P4Ig84zp2NAZWi/vefb9f1rnq/GmLtJW0jau2s8d
Uv7SKePEHMUtPQnOf1STWVrviHdjKPhsRSoPsprLvU9qjlhAhtfRR36W/8b4Gshf
4T2wJ47kJYtRx5vlZikEoFNViJQRuBve4ghznyVq3hdREObDENY8gMPhYb2IlydU
XEWJUhsacssXQYS0RmYCP44TH6OmPScufx6SkOuYXZqe/DDeH4FOcLR1T8hyJk6b
+uaCb0/12kwUN7CC+oFLBlyhsqCaU9K7phtNu7M1AMNufTBKvfiIgARZ+vV2iYQl
ovfWqVmiypBx/rdiknre8P4heIGNb2y8k0UhBEfmsgjF1g+qUfCLrCmydUkBKgcW
BFDX1rs1fKlmxD7guHvQfxzSNN3KvUFZO1FNVd3vVe9+B4tSxMSOs8CCtNwgbzbp
+rzW4p/oNgm1ZrAfHMC6/QGuUm8wsDRLSQl4xtkrnD2VBziY8rt2OmHaOLXMmHT9
BO2Y4itY18QTGM0rLJm5zR+geVubw8dGu0UzQxBjRwOVhgZUAC3BzUpY/3/5q5Gw
IE+zjMNx+23k0xbaXgnpl9jx+OeErpi4u51qMctzLh4XjoLbAMWOoqGeY9glqRI5
FiSfC48WM2Gw/oasG2LMf9c4Uag7CpZ+IK/fVSG4toQL7MqWbMC5NWnpOthq6gvx
SZ2MDRrIpkKEYUpvGtCwvqjtTNmslLGlfeVTc4CcWEbsJyfZBKN9ROclfdPhedtz
92tbrZsiFZDq5jBA1r1jXc9BWu2brrDNsOqEed8Smaox0Lw6W8MWjBR/SEi6Klbn
B8MaW6iDD25iE1xcwrswFQPWQr1ztKVsmye3AFcudN8cWkhgoy9a+BeC5wBAjsXA
i1QkxYPhXio6tMH2GLOkETIQfWrrMT1Dqw7alBqJG/XGXUSQEFyqBulcR1ZR88+p
mcifgxEBecq+WfTi4rsBNBQ3kcpQvLCLTyxEUY80SouI0Tc3JV6ZiuNmrj/+TLOJ
D78H3nn3cL2ICT68zOgjhXNdxj1V0tWfIlXU/Wdx851Dp3Wx5GNgmuv5rG5WZwKG
JhsWXwd7r5YABXAclnPIfqAkum4bvOb9tMhpaR2q8MIiALmJib96fg3C5wqyNemD
1C6DxslIUKw+ZWkJO7tHmetPuiOruPnLFaziQvWNf/xsbpNPOWla4z/CY62Yj70b
3gImur+hX0K72PEuaEsJ5g7jpZdbIr2tccrQHnlXzVZ0LvZMDAUtxTkwJ4uD96N7
x7kp4XuC1KfdFPfGI6TDmbvueElUwqHjWv8iTY0mhlocfdgve6FjgVOV3G5sGLHE
h+2YhFbA0Own8jiX1brxjvUBzKYYjqIaYafCsbTANCb4X95vL+CPW5rKONGac7zo
2Ljc3yckkgigO/klK2yI1gFJPUV2kBlataQmGRgYNFKTRYL4KA+qftn+SFmGeXSO
cR3Ohrw1KzP6esAczQEGPHsimivOsmWQIgFZTmdDtTRRwno1P8NBye81p5J8Grtu
OFJPasporlsQcXnDDpZIArV11lhF0+C1/Sj78I7JWooVA1kjIhzZ9+DQg9o32PKS
GOthyZ9V9u73y+SfEiCZTN8rhpK23GxLf/dC/OJOL3yDod8f5jGPoY3YFmwBUDvN
S9GGW+TIBKIIiEf9wy0Z6zETVapSmgr1Yf4BNkmECNsMv51/wfEWRFfS9NO8Ta1f
yrFK8SfvV9DxIz2HxUTXkiabGlqF/IVqekrTKUAvT7EWLbvdfjwGR1DyjvLWH2xt
sd/XBfnPPEoKXY9pZMDgJ94T8q7LA0tb9XfiziTe5iOlrpNbmEd6JaNUHbQAur/n
Z3ZhbZZoP2mCS/mKcgFX/7y6DvIK83v7bo+5noU5OGDwtTZlXG9KQSczQKa3LmKk
wIAv4kqMZcl5duY7Wq/GGWBff/RRjoJOHSlsYwl8GiLiHqktjd7YkIixVIJmdk9Y
kfxcmfytsuI8q4xMKK27gbIwAc7Je9XTfoDKoIxhQvf88u7kCTARVXJG+Zed8O9U
jeAH384E95E5/mfCFz1kiLKcX/JqmhSVCdvuyysTOsUy9PtciMk7o6e/YqQEvVHM
Y3DMgjOI1Soafl6VLRv39P9LRagSC/hf5c6EIt+vENIj77rDHrisiQWsedS/qqc7
MPjPhIkc0kQQrvrJKWGza7xmAYnBwwr4FFYjHARPx+4MMPvAhhTN7yw3X5Uw0ZKZ
LKzkf1W+D4/GFIrSg3MV6zyY5giznVRFaza1jGgu+GV60q67ffJVagWm+1zkey8L
agbftm6NfMZE8VZ4fx5tiohiQN+1KbNClXyNpTds4fZCWsXMMk6vX3DetsUssRXd
kYifZG/TRigSs01v6EbiaUa6vU0AD/v4nzuQQjWkPM/uw/eTQbenVOeWyb1kbzK9
Yf+FbCp+s7e1put381SK5JbeZQvQIWYP+PoFg9Fh2Pd1kdnOeqFUwzi8P06Hi9E3
pV09sMbJTACnHnGulhWUAXbVa+h14Ch5796gNau9hXSouR6NCNS/kjomZ2pCT/Mo
QUETmQkiniJd2Do4v06Dc0eU41qw/Qus5vSBB/NDU3Ts0rJDfjZO378W073C6mLV
BgAuY2VDOnIGGD8BHjHZ02uylIQYOHNS9VvLOvI30c5LEck3QL+OjquZZyZrrfV2
4DYgH4d+RBrdYyUpH4R0DVv1fxj29n326FtGubiyhKmLJAvMHcx0yMh9DqLBOyLN
FgsHYPhmd6qcpJ9vpcoBrV5OVeNkupuQsz47BM296KlRf9tGSF0L7dJhCV7PA13t
KYdSORDCGNwgqhKMegplRMtH4maZFYw9tfWirn1CNWxNVTmNDWU92tapbhMyi2aN
WAwzX8mWjiTxl+gQ+5D9IULMnA51VrzKZ/BDP1Ryc1db6o/MpdZ80XM/oN+QtmPF
k62Ws8c6kcLZjH5jw8801vmw8bWvlCcOYSBKBWNfyfkufAwmpDVRcgQ/O+AG0PNl
Tw03TdBnuCh3Q6PpGu2Pig69qOfeX6QySd58OZMq8HSdGm+sSeQFwvB1a1ihM2bs
M158gHv1RxQCzAvA5wiaE0IoJ3uRzMrOQ6M6B+kdxzSpMtDP7MvhZAN+iI5UplI9
sPdOo0KhpfVp48as/GpCsNkQ/GrbLZ879mS4b41QeFgPP27jDPC65yZYo6uBN2h0
CevNXOMvoDm1d4oi3/+YfeZf2+DtNQwTh+uvNKiNujX1+V+apZxqnvMymJzltoCX
SYD6O3m8pcDPti21EHUnol0rH4IWoNDi46uggYczwDt/rVKb+cuI8/6jRUHAHJlD
UVezCtPjr3fH12jZaZJBcQZ4ctkkycQAYp5YG9+ECxRDPL7UV1iiXSbzcOQ1Ci8M
STtaZQ4ElUcqSXK2WaYsf+vZehrW8rrbyxJfe7f4omJ50I8yOixcPkyuKQgICyHg
XNZA1C5lm8kKZ/HL0T7BXXi/GAZ73630YA2I9IuU4PG0myvRo6+uZXuCVWghZ2+k
z+eMeOiZOKljMfdjo8mrqKGXEzYqJh9slncUOZYBJgUpjqD9INsc6ga/+yNY73lE
4lgjNMRsX8/ogokNDUZYjKcChv5Adg9eOcZvzueoQzE3c8Gg+Kza4r1m3u8rFrpi
NdbAEbWb9mCgBtwWeu04fY3qHTvwe3sMcY6jeCIQxsBlqp7+oQ+Fwl2KA7UE8iey
YX7Zs6smcaYg3ja9M3j7lAmACXjTA+NjMlI5LWXN9IEdGohRE3sHhrPGOx5BzRGW
z5SgoO+JfIZ3SJs/CK+AxjQhmW72lSPRFRN4vts6X6100HqOxOuEVQSwjCjHVKHm
BOeIFIyGki+Ds9mVbJlil85IdzmNeYcgfnv+OkJ8biQbujjALtiErCZafZ9kG+1W
fM7wvnhFSh4B92VMNsGwPta9CmD0dCrDuXFZK89RDR353Fi6SsYQhDTrpNj6Z8M3
IlCrwSvHvCPzGrOk6OOjqY/KLJ4OLv9/2pQch4VptjTonC7Inru5roBuI0ibz+89
rA9csGQ5nlE4bRYX0J/Hj4nWiubjkGJncjANdvskkht7XzTAmmwz0o+Akk/o7jdT
KrEnz473aTinOJaNO9bpSIuhoSK0bzKXP7V5Bv6BV+gx+iDqwsdrJAnrSkx/98lz
tql5Lzyr1MaFz1Ig0jOiTGy+XqSYpnrTxw2yOoFxYtOaOciGTG1goo442Nd4Igdd
GIQVncEhgUzZz4PxSMyjX1Zg87ZKdiVBkHK8VAsIf/hAy6Vz0sZqYfrSN+Mx1bED
UXza8L4yPlF4SZSBR3oJZ6aajVDMtjNwV1TpJdBgJC22z0rwUAC05QMPn3nsNc/b
TzcGQYVQJ1OVPbCVn1opp5hGaxRwoE3BKYDOGB2X14eiQPfqsQ0YJC4n+uLuNKX9
/+P9nHx545bs7ebtLU1BWV9Yk+3sLSBo0NMFqZIx8EMOaaElBXIMSBhP9GgIB/yg
AStgcGnp2XKWIBSpf43352J7nELWIJkH9wS393MLFPrBOc+qp69WPMOqwfXHejTM
n5kjSPHwSskUD9wj+3ZkU26FITst5LZZGv6oMVJvjV3guuh6g6Y4jJWOq7hi91HF
x77OzrQc3NVrh+QyqcCoq2YCrIfU8OFSwDaQWRY0i1woCtoPvWLnElakkbPTHsp5
r6/ZQaF3oWoYIzg9HBYP6AwBJncRqZQ55lRcamk4ySHNBtGBa1ypl05vHfHmzQRD
ytKhd7rNT++Wpcnn+RkoeBCd5iVdGckja84rNVurM2ShwjxeQiP+/jOafN94O45S
rqPPmpYfRUQvoXm/tS+TrLHdLvWkwxkkWUoVV3CftL0yWD6leu00SCkdwG1tzl9g
YqzFh+ekrp5YOg/1o559/bplIvQYVtwaBnijTHJgYVJjHjUfvhxeqF1Yv7kFAlJV
fpqW19BKx9AbChCZP4Hhn/scqX+JjwaL9KZwgT9kELZbuXwBh1NsaWxJeg+dNQnI
FSY6/KTya4JJD9GzeE+ASYUFUh8VTVqflkVANZFiC6w4UVHLbEU9YMfIttebsUCz
HEqnomhgnrO8gpywNtYXf7jn/mFMNBGj83qDCTwOYfnAjl2MwhxBKPcDYTCi6UMM
LzEZmBDiFa7+7/amw419h9+Qre8R8pfmYKdyiJg1jD8INxZlhlzcKPPy9ltoFYSD
GpuQN5VnslB6fMWa0WqOhQEM0PH4UpjhWnhOA4fwO8Kg2Jspmmtp5DKJFRlxiaAh
zZJ6Reu9K0psCuKbsnffqGuKZv2xpLnBX3BC1Gy085pxJFoaqoXavlC7R2baeWUB
WA8sRkDgEU6crm2OxssXJmJw40XdsEWDUH+ggEbOAB/qWDHHpPixDHxFU+YmKI8n
XagsCRJrQhJJ52gegUdw6fLDq7aNmYj4hhPpEvkJarQf75ivyNQPwYuJPe8KC5zZ
bFNmkfWi5Czny0oi6Ml3acYQloqNNMnzxQELOcu80GiTJdHGejA5Xk/RIfvTFGKm
lxsnH23gca0jwgqNsFTmjH2fPKplQEKFU4AttTn5hcmp2FpQaynpPmPPaXPpe6Tq
wWPCew8yoaFWskDF1iq/uF4mkKjT8VF/TD7G1NJtA5rK7jygtZDdXMLSy3ONBssE
Y+mAjTzHJ7qHI0CjzdxtQ233fyCQZk3GPl8cxme8XlUHhzpxblzS/etpYwkMNmZf
bEGG5y0zdBk0IwiFSbbZKn+BL2TfPbBwiVXusQOzhtbbOVkG3W0vwRG2wh3Jlzjw
kF+s9S76wLMlQGeRBvxneLMN7Qaj3Du+dsSaDB/Bh/hyXeZbnHned9I3w5O1FQWS
xCS6WOmSYKk8g2G9Jms0wbwzJd9aAViDjKMBTvVxPOdLG0bq85QPuuciGb5s+EwR
f90YYkuNfIkGcxeQ6Vnv/f5yV8JEworr2Q0ZxPvE5H1SbfnkTNBHHDsQZFAia5fu
deNeNtJ8XNnFds2+sOzLYpVtqOhBMK0DWzY64xdK2iXtX7UGPoJsWlK1EJwL5ebT
apaYzTW+kO5pZkgf1r9hwIibt4zC7GkWkWgQr9J88inNJkTLa49uoRA9o320VRI9
rzj7KhaLhPPV1C/2XgMCwrW9Kc36OwbwOxY5eEsfvyB+Y9IzfwgRoUf9RW+sqmjL
9+hYachqZWA1YBI3GwYAPcpqaPejpcj5L0wmLHNJWtGGy2PhIOqIKjNw4ZN9/xlq
DfOALJrLx8DGaAQfZwavV2T032WxkNn75ShFjOJtS/FzAYQPa4zvobxgK0iKMGIf
sDfr44qjfLRDtS3Kkckl9s61Owfd88+sICMI+2l9fTCnrbBy2zeJ0sc7WzG3xAuu
pmSzjbNCW5460A18U/5JKHRYSvfMyZfx5WBrV462xuLKNZ0hZhXcijEGAVcx2eGA
A+IhDRKb4yqRY3kG3hshQljC4XMoXtaSZIwtdtcpVKhJdxIYZtOZqWWX7M82Fl+A
GgXqn5AaaWcaETyk6PqOtO8+VZJvdh0kHG0GKKExf2HH8Tqt5dFYgJ2QzGlL/ngb
DVqxtlaltQjdczUy+seHPwxYn/KHJdVIt+4wBTZ3XiDW7il7XbV7j9e3i/hgB1sB
CCyRuDPXtPMHcKJcv4d+XRciOu5/qc0zx14UzmYJyz600MkkiAntmvKMqqwtVd95
Njh4On1Z3MKRVbeUwWMrvLLK2zq1Nrw/8ncWmwKXEwd5DtSrT8mpAbPHgCxr55/h
ICTOmdEMfBcI7dEW1hX8IUGf9ASH+OXs7DP1OgHiSPu3pdOxjZDV0mveQ9ZVfZy5
PMxu+H9K0m3gi9mdEEyfalftQU8YD2MSy21Co3bAS807Mc6f7g/FURHLMLyHCUtk
QkGDFd7O000189BD/KeugBq+oOk5O0JikdQ1VgkGEllT7tAauSX6jBRh2MYuA0PI
BreNN+L3D+OJQGfoR59SXBpVmDmJ56HT82aQebLF+rDcjE087cXyhJCMjwoJD3gA
Qhz6hacfPxGYlJEO42TSlufb6osQx4MLn3s/uRPqfP4MQXgBhUXhoX/0665jtwRJ
sWfzoWOfa0q79waVT+x/DmcgHmKaWYa+FkMa5rI0LrFbY/bocAKFg0/lZbp0OdEX
hbqaBMhZqFiLerkhC2oFzLer323Ma/6Fmib7CpHXyLh/H1g3nTmDXFpn1ivL0NNc
pFZDaTqBQ4+eat46lDfQJARHDKCtXB0BR3UUdJbkhKMhCLRV33OCouJaAIVwQS2J
+A7BVlMa9ZZj0KEN1msxVbFlmy6y+EYbljhfE88QmoRLQGbS+9Q9eqcIuRngXZtz
senU2mZPnSF9zUtJgIC2vMqDSrNXRRAyoq7Y33TCywzs2SAg2mS4eIxxkqzENlsl
ylbZamwvCcgaPxcBxYuBVoozG4s1D1zBrOVuht2ERbtRf2yy1n+0hZPikbkU5/Ec
/DD24IjjTx8Bt9TOgJw/2QDovmd/wL5GY92KBV0OHxPFtEQtkHRirePgR7avrGxQ
KpKY3+faQG5s9yZDjMt6j1cwDHBHHSYMjri1q90nkHm1HHX+M+oVBrvwEcSPR/sj
4JTpQoiOM3eTcd8dmgXHf4oBsVnHENOcd7gZGAN+aOxXk6QWM1vgZCfBDqYTWA3F
v0UAEdx2otAjueOxv63EeXKG8fAdz4fX1UZpx6jpgnB6LVxSOr6tXQxVyZxpJFgG
onn1hTdDTTzoj8Qr4DQOaewqXsFgoS9GT6TPy2uVIqu3p9jC92fxkVeGRGGIIXBW
Ejos3bpvVeglFMz9d2GLSzNvhClO7LM5oaOGtMcpLk1UdiuOcLjJRYg4ZzOQsPuf
DukxX/yuBPADhKb1UV+l72bMkhe8vIvOUCGbb9SMjTdARWqyWMdWm4Z5Rt3+XauU
6Skj78wC5G7pkfaBR1fMT2rB1qtfFbb07I7ugL9heHUwy6LENwgqXNuq1kUYXIao
Iqv6v62eF+P45Y1JxCFIH7XS6bWMSh6aPl5UhAHRoYmPOfaEe5FXD65i+mvLji3z
l/09yUWlfqyThdZJGH1Oaq/VGsentMnVmvxuTh/lj4t2no1UHIRxZqMF5mE8qLet
myVjxB/3fFYnXihWzPaZnDcKCoEMTLEUpPQk1TjOtu6fYAtswMNw92fGys5zyHwL
t6p+zbsI9WK1kF5szQkthR78y4uDglmL9jBufo7Y88rgT5Bz+sOvsxOWBtXMSM6d
3KJ2R7k8NlPKMDcXQftunRUtam06LIxkSniTN8VruBBa+f//rosRpJG7bnniuqN/
xxeN6v8l+rXaVhuCaMyFb2nmQm5cRJN67fHe4/ejfMFJSNmEwWlnQzU6k0hOizlG
jo31S69tqAlJCjJ5P1kYyJfNHJEw5N8VLt7ymluQnicn7C6D0V+PwdXGD/dAU2R4
ItvvfjJ58XsiEqaISlvGv514zd67SQO6K4QpC/olzKaFDkNzPAcShfdTnOXBtpaC
gBpDdjHIe8FcTxkDWWEIkNq/fHboXGKybhYr81CighaV6KRE38N7zNtNvwV60Gua
ADXLCIfQEbpH+/uEpfHJsid3tYB9OH25QmOk/AV0+EKke1D6/48Fy6v+wgxqBo3l
frV62WwvchT0cU3Js/9/MQsI92Oe0ltpUqezqZs69FmqkxMSImhd7/odOvTlVTAP
Shx8yALhBgN3pm4Y0J1lk09nLjVaoLOyCLdZO3QEqNvTtP2i4q32AegeLqrG4K5Z
ETkSRhgbvqGTvX4IJokT7OPGxsVWlp4akV3swUJ6J/JWSFFcjbUuyMNXd763N4lz
lm/iiFhPuAuoC0aUs35IqDzWhMghpyreyjfFgwrDzdORl0mSpHh0KDgJdOgnkrMd
JhAmWZVmydEWUA+zQri2qLDsJraWMw1csXoxxgG85GgKfsb5TnkTjJjwbqlApSAJ
f9QpcB5/UeXbrEF0P77sedW4MRiM9Jdj0KU6flaohukdnFOJ4OBQY0Bz6kasYksI
vP4ad7YCOLuDOT+2pOyXu/fV1GLD+HMrDxXgMkl4sHhqmOknEruCDcGMU3tB2mOr
CQ7MSJdvK5p8VRDDJ4eED4XDYCEZl6irW1d2awUMM+QCjBIr17eltPbB9qwtwFGL
66yP1jDjW3yhawLbxiKnB3wJy9GmkMzlN/fTL6GIrpXRZWYjy+5D+mgRwO1yEUMI
e5JZBMXcxYRkCJfU6N81j3n6bGqCcO4O1B7HMAM+4UUO3apdmySgFt8yLEj547Pu
Ei96Ye6J4C4kgCi35al3OCJRU20VgJIxwxhAUDm6ey64bJr2XCuzJVv0bZIHgT3C
wFVX2ujOJBo1suYUz3BIMNnnqjo4V/RUJ7NStH9hcsf1VAKciaJxYuTqleWsNl6/
bQYL7bpytL8mIz31myGFbPiVGWE9HYk9VTkqBY0uhjVhagTl8CU099d3OyEBS9/x
1Tj5cblAXJH+elRaBElrYHRrmZwe+7Np1H45kKi2eNRDgetAOspQuN1eKCQLit0Z
X+dQvUZ66NnGmdlLQAnJK23N++KIPK2YJYeH4wodHOdcwL2xPb49RjWs1kE9aT5I
e8stmY1BHfAXl2YNn5A/odbzV/TnS9YjExQfex2vsH/6adPWtCHl2Y/5H17wonqZ
mNr0fAsdm+lPnxiV7KZeepF+ydGpAL1eWz34eXpP7OG4FGz6r9+KUzDQmJnN0t1w
ZLxIZmfnRuXSAPWdTulFanpT+Dbi0cvP46DHBD7wmlPJ4rDa9O0pBqrsbJIZu1C5
u/Pd9lk/XUbAwtMB4sYJw3hOCSEAsh5i0N90K76f5VeNsYq1EVp+BdJVExN1pL1K
pmQYJGCUVvKjc7HOMA600CY31tmJZLZbgbhnwXQRDHVgviLuQHIimqw4YAK/E/4n
x8ekIAOrfw0UMEPktoQwF2f4WBmR3XnYscH9c1/7YMP0zm9UhEjEJlC01J7t235M
F4Aesm6bFNA1m+OeT4RW/ATvizDAvO6uwgkwnqmz7rsiOE8oaIDavkQljewI++S8
ucmoITo98mE3bPMgQG9GB9xoY9ccIhcFgGHoba1B5ZWsa+9ZlhPN6nPKwE+ThM37
di/yTRVseM9ZmOQKhbZMMnlXkQUcH7VQnoTeZC5iKkC4wZ3l7dEkY7Zu2BRJSBcm
JIDEPUMAdoQOSeB5kXkHVNLV1hCELUPd68DxiB4lkE7tcVUu7maIfB3lII9AbT6r
P7M307uWqJnoNM577u3mhEK4OIZ/ezQ0PhAMbvdK2IEgdJ/OqO5DXCHY9/s9WUDM
VKd6+keZmCq7fIS1bgP8XU1+x7hFPY0D0vHoPUW7wu2v1P+yTpyVfyMtghJ6s1yV
KIs1NKigUK9a71bGWe1iaHwQQwpoItix4u7JNDV3ARF/cfsPvWopN0gszY74n9Dw
NZ6ZywHAms2Mk8MZ8u9FA4x7QvoVHfZ/a8iYBrN6Jdk8XWTQrV/0PJQRvnte5o4D
D+Lb6yvveMmLKovgM4i69kPTfuUxpcSF5x39P3jtDHhbEDpQQfoQ11POG/ndSqWY
DBk+7NxYtzaWJh3kSPXnCGS/PcJefAk/aDr1KPFl0uQSNT3cX0w2fWNThuD0Eeqg
5KzGK6Q9WAz0qDL/yL98wviuJ3rahz/X44KHLWEBtggExa1H7UZpiZGE359tnj4k
XRmsLxqxPxLUyrGuhO772LkIm2gnMG8sihX+WpBeCOAmqWkoPZIc8DcBlERcc/ws
jf42RlUXFRRrohRQqd1TtTq+Yby8JiQ30exio7oy6kuZ2YEqCGwUmQEDb75T4iTZ
ByAgxXEm7hiyQAnR8aPUoa2+biZHvMv6ANlDf2iXCfr/nKhJSQqnN5UdS4ah6/WK
N9PEfe5A/2dfkLVkVLr+8d1ld2uqFfoYX+xrNjrFAuWNbEFiyr4XchdL47KDOh+H
qmdy5q2WuzNTq7Zdx6xfovd3817Z20oXH07Yb5EpjDkNV/GpMCJLryeqYxBLc63h
8ofZjmK5IHMqjR3Cmq4rilH+ALtVkJXbFtCJFP7iXIbmyB2XaZ1IdthLt8MmThqt
wJ22MsQDD519tLyuEOt6qmss2I5sAKtjSP8/pnChLDkVl4wfi5Jkeb8uBAZAN9LZ
tuOWjMaofxQRhonlZqPwc9VA/SthBLnmZqPCp/Zws4kvFh2/57md+DK2BUpI3UOY
vJL7zLhuqXxzUs/bUbEVvLGk9pJWA+jk0wV5QNUcpBWbsorjyV+tmWcwuA96rcSc
h7deIbKp9nj+qJ37J8KcP2ZSj02x5eB+oyPPt6fUBBGQXwfqyQCunEIndZjfJP7f
Bak3OKoDQqAToHbho7iC5dUk+q+LEK3iVZvk8GtSMTQfe19TX9zY9RP+iTmnN4DA
ub773Z7aFyc1y+fnC/PRfkEcKMQ5KirfSrWQHm6ZynOhrsy37bIQan13nLjlEvwF
Ma+mLN0macNAMNOMOJv+/GF+1M2GPdz0iksKW53x/Fy3ALfIUx6PfWjdy5fizuwi
+nya2Mtpo5/7TT+WBnhaKy45s1jpLCyuf5swBP6kNYGuZNovJMx0IdjdrmwZtjAc
nCZrwT9mqZiXZlyxNXFlX9BPgQtMo2XHm3xn3VHCtbA1Y5or+T8cz/49Bk3hS+/p
a9/ZInhGHPee0xOSCafkPC5ALafuwaxY+TAVMEd3Dl5bGJeGms8U47gseBUnkY3h
be2z7AQ9KzBGrpZhZ46wtVFQy0NQcF3cFvj1Vo6iW453onHpa0CjksFVKeRWOuSn
DT2dd7zEWbQfLo0i/LfNxOvzTeGht91wDlRX1TtoOTFf6sCECyg7f1171rvJWwZZ
sw9b/Uf0oBwnA/R/p7v5rTXsilpJIbPnD8OssPryQr+BbvrTzjMyQ7+0SAB8/BR4
EZbxCkQffu0B+beA+n6wgpDZKBp7VMDZcZKdZTsoea0wKdHfSyC429MCsgHFGmpk
+JE3zQFhdnk7RhAYg5IqPvftbJbM5BJenc10ZST9hF6efzHcz+4duWemWkdPbMD/
7VpVK8iEWS/wnL0tkp/mYeVYV1qCjPJFlNvjGvp7K7lzhsvf4zl5ZDkToZlDJ9st
AAAr1hlvQ5Q83xbRmnG/Uyp0r4ezKXIyJMdyWnE02b+VqJc4QiYNFLnMVY8Be+wu
p1VMmc2W+P6X+feLDZdNzfQ3S4cpnNRLzRjcAjWgocE4bKKMjKl8sZfgw+/9u9Dz
4dQX/Nnqk40VmzUiposdF6lleQw2LL2VK/VUMOVK198xvlbYXqr2YTgujzvgHDMO
klKdmaAaPLklB1HoNHEES5Pipv+AwOMav+Qv+N7/lQz4xyofNdAFDmhVohTU4kH/
t6FDDzhdexkGxnv5y32NxFvUaxIIJqdNehH21Llf3TNeGQ9BjsxaALzxOigsLJT6
cZZSvuQZw4IRdq8H8Lorj+veNVYye1+gLN6s7yRGBzcCNdpokXrTtW/eUQiCWRnE
5R9VGJgWbWSpVULFsoQyIHknHEZTPmRO37lDRXqpUXqBNyw0WeQrakaSsYqrWqf0
1147AkZrtYFYxlQg0GwNzwFqn3V43GeYkmm9ENmFDPkn3qdgccDnpAifMkZPIQD3
wYLpUA4yNGy84ezgHVmL1nEcwv4awIjQM/zoJCFc0ZVJH9Zesj/cr5mu8u8MYgKY
o5f637dW2NUl2ip1+l9fQaoQycD2MLuoXQQH6F8eBOHejpOaC8ymivYgdWbO6Jrq
DjA4SjE4hSLsle0Tvn/pXp+MptBnezcKLr7hJ7fuE8OwIZS/6cXowLKDYrtMDBGQ
2ny2NjTxiK66D5g5dFgrCuE2ILAZy/vBy5koaW1d5bFioR1Jh5+UQQMIi5z3wSZp
vG1dNgJtK9XFeSSQ0ME/R8Gs4zNFMEK+j+vt1cY95f0TDcHOKKznEoAOZ6Rpg8fU
csKOLdb1TKaTcikK2jJqHQRWJcXyzTz6DSXZZtkAUiyrXIOYM6v0YZ0JeElJx6Ty
4H2ZwAVV30dsw1bekZ4Yyt5cQ3ruR/LQKf9ufk28RyTGToAEYgtvyMyYF8CSPdnp
iYVpoMG76/of3iJPlKlnShBQleCSjBGCEJyvQY1z0hHkZD/zTnW5IypzK41pIc24
SVZqdK8LWOi0Ie0ZoMA2QKmH2h1jUFOXa+qUbYyE+ycKRGrOUbBz4PbY4fSwBneE
BpBwxZFweTLs1eKVlK7rqQ3NlJlA/dTPAC+qpB3nBItZyPA95taaYNbhnOCCADiZ
fuZ9ariNA8S+F+UXB7sqRjqUeGwVxbg1CssZgPmbz3royAmgIL60cvsF2NhnAjOd
kFKR59ryfftDkS5c1fW3UZhWgtEZ3kXw9v1I29JdQlpF8/aCJieN0D5+0MGMBPsf
cGwpMPqOJtvsFt+khDLfpUfSnLWhuQFHapomZVNPwmLixT23pOXR7Ua1n5YWbGk1
NkuEqZbLhfHM4MWOCN+/Q5UnFYmGpCUn2ZLjvMU5A1pQ8q+AB7CuqRH7KFsa48F/
yTag6bbjhHD+MgYUw1nrmULKT5ZMka8GSlni41FzaxFzkg+5EQlkSdbLZsKchiIF
r3SUQe8zHsscyQICleftiY1Hc/k8xx6vXAa/t3mJhyCOhaQTruf10IXQoGra7Gcp
lPizOAeJwhkbIDLWwxiTW3F/CeDLJE8hSOIkS9ixBtBcKSx08dnwjTJ2BtPtIq8S
7DZJ5f756o8aAno6LbW/Pt4QOgf5agxg/Ue4qt3XQGnVrGCFcSz2dEs9lm3+ZD6l
AKmNb9OcMnum1ZqjYaxDaB1iLPc+sn7mJgBBnzEtgQwQFVDY6XK4IxuiI6E7imzG
c4wb9hq4krHOwYvQfiAEhmv3a62apNEL8r1KKSrKm2ikCt5sCpH2QpQkuOD5yA+3
rdwVCSeI0isZtbRCaiXi74Npfem/3niJlxhelXz1CrQjZ2X8OUNajyDJpV9pI6CT
WgYbnVK6OX1LoLivwLgP+ns+je/alMm2FkIjaYJNt6lkVMDgi+oZWcRv+LX/KaX3
hOFHAQ4Q0Pwg/Q7NoN8aGIK7Y+8puIN7/I7XmOs6D9zBq3L1qJ4Hg32FTmqufH1K
+30lbnp+iqE/ZiTsMnExLIa3D/M+ti0HWJTI5j0U1MYavbs95Jt1M6YEnJKNDUFy
3P5ZLb+jZuql9J3lz4Ci8CrbgbaxP7uXAPj7VofYMQfqT/3qE8WwHiICr5OnAU5w
KF3A7MGTknP+bN5fzQ6VPrtT7g61tc5arBEzjo0GnerptyGPcVCUqRvuf0pv9BTi
AXZtYVBpvaxzvMu5OBITQgu9sM8mv6FHDCLeiP20ufGvpV5gKn+kxhsLpFwnMe+p
jwr7L8ldwYDZDQu9qtTPsAwo2JoNHFb8VbddHD07bgbLb6CevlKRdkZB5mn7DX4e
SfRCTRpyYDso/bo6XQ/xv2DPyJI+WthEp1wjdHkqoqWG+JuGYhFXPfa/9t9gZq6f
okzW/JbylGJ4LJvHQB8wo/1cMvt5GwJ+gtaMror8bX1AGY+LsJFkHXNLRLhCiTwe
Y24TR5/t/sYZDT+ZePq6GIBUm3TbeqUdFsFj34NWzqalcMyz8clC8Ze9humDUdxx
ZqKmuXD4FYEBp+02J4PE+2Ql7qbFox+TGdciySZr+obFzq6NRN9kbNqRWiLW4o+G
9Y/qmWlbiSiwXeG+I9jrw6BK8lLo+5Ao4IDS3qe5cNi9nSAMW13SBSX57hM9dI7R
TtsXY6Mhy20VruoCsM7V9hnqf7Dmas68akrVXRyxh0KXGzzAhX8WFOHmXPSNZF/4
LVZAeCiuXhbYjlLP0D8x+EjNotwwzakOnkhexBjHN69+SyjTOZ/KU50KDWbx+ug7
6R3mske4hpl/NaWtoJKit42NzHksTa8a7cpdcNuijGArx/4QuWpA1y4oz5VQWpjw
Y1sEgffLNjHq28yMWr/tpbCcbDU8uHLp6yAY0MyTbLVCfcOGxo3MbXctXGJn6zKR
srWBOpDt2Z7A/zCvzU+pBWTNeYD4nPt3/YnCJ85AciWkCPn9ErpPu4xQ8kiTb1yc
O2O76RR96rlaIoop55XmBXLkjetP2nDP9T6gTsIeoat+L8/+4kUXoHFnDaehH/EG
h2GOaVWI2rPae3pdax+LHsdLChLwhIcP3LHHwlr/YQrSYC7r7EwxaWfoweRVDaJl
iDqXECKppzcPH5zPeHAsee1dm+UaZWW4Vc2tqU5Whb7B47QHdzJReDnhBhqBJNF2
zeSN8LbD5orxAT39KYkl0B+u9zYprWV74Zz9tWKcIC255wOh5kIFiUpaEWk6K83V
hU11/ZFGtZTCMaGWkEdn0C8mZQGetq/pEWutwO68By/V3nqBCtKmoWGgSL5A1u7/
SW+Bjff3mfxDszIDEeBTGtVulLUK+V4tDIuALrrD7ry1Un52xAIlcP7ZzM+luslw
khgYj/JZPVYxZqUejeWlchwwK+dheQ6IU3K2/I8/PaK45M9aFUiwPG0/GZCZH5Bx
tq2ISAh8CjnyJFO45y5PcLAet/5qPkSI2GOUdngtaJnh86gGst8KA/QAFaxpMfp/
kSQhvb6tnVDR3LBqxBxP+BWCEOl8eUohVkKgbrmkdUByWfdwzDy+FM8+dhmWNeKv
vJTs3Npq/V3ui5VVyX5CuyJvKCkmsAD8p53K4E02CTi1l5UMvTIJczGKh27t4J4n
eAdL2XSNRiWaqaFkUWKKJC3IIOHrhqwia6Y1w2i9cvrjQdh8YEV4fsym73v3XHPi
Rf63r+yUI8lQdhzzM22UlHCzsl+gikYUq3GyNR0M6SHO6kPR0O+23sCUkjtWGiYu
brAifGczI0yd4n/PnGgXHRJtJNxLj2/cRqiydcqUfgFd/IkN9OD5UZMT2d2VSRqt
YregvCM3WjXK1hecsNO6NWh1rR6j5Z3b9+WbbNRcftndtY3j9cJ5rGJ9IatlzO6X
K+hcSoH9zU2jkcoERPTnxZ9xTsGUmTsvaq1xUKlDekz0ksxd5Pw87H8Ccp2Dg0sx
1caJySF5wiLV5JQ7IEKrGC1xOtDDjS75kww/syQ8+MPW/mWrZd4LVaKCfDrc27NY
BaUA7MWtTd1JIPyfiPId5aIY3A7ocnzvGaqXJkYbTJZPWJJHs/tVGv/xmXnr+H9k
oHP6NG6UISQEf5P2ubxLgYxe/ifDhuwQUk4H24MyGPOqJ71GgziFHVsJVegax6/5
h0ECrP/ym5+yjWMsfEQ3t8ZC+/YNXCzakifQaZtr/iUagYbT/diLfojXW/KY3LyN
tCnyGFUbmEFC6S6Iu/PIu3/0qjqTIu4zCJMC+6w7X8jH0jk2ISoYloX+dLoSxbX5
uErtImnkE58KmgPrsTw2CvowxUZuJJdqyrN/JAocp4KB5iybiQ3R99G6Ud+1irRt
XOloFhGZ3Ed4zdBA9JWywaQ1h4QmpFgLIwov5kcitrCRvWwEBOP636CQKro2Od+t
2Hay6VnSZWQNAdtCMXqIs2BPOJJsItVugwjGzk7TI1l9VNG7Hy3AXXvBbiEhLWDH
N0dO7h0/QxKt4QP4AQeTDDtFC3nBw6M4skktTuvQwZ/H8YQ8H78UjEyUXPBPDUZ8
ZP74c5d+IFOtRkq/Nj/dlt7P5sBmgSvLzvxW1/in8MXVagw5Zb2CCLdKRsAeAs7D
/MWvCXxIFuvd+iCvbf4+iz6w0GjXevdny7SsKzDzeGPiH4T74AhfY29+p5j0T7WA
Qwa6RKNDFQxtsppxt4T1z3VnfgqpkbeAYNESTjK0GRyWOsLbGy7YzwWxQIKbjpXm
y7lXBYMcImmGHIP3lqeL2/Jm2P1LZtKFvKy8Ze8rsejA6WZeTmORGep8V6jEtp65
kaMQMUbHESa/fAIcWu3To0xPZxd94Yx4DXvRdGWZbCzLivCaJ+XKZseNUSVnYsBC
IrbPpFaj4ZTnI7h+1WOism1fUHBCmHyWgltWLFGwHXb811GASnAfmdWBB8v260q2
BMMbSQ2T9hEqBmrU1Ysv5Z2GwmVL8bNhxIiFo7yMye76cKMHe3/SlvTvkMNYSu4Y
odHO9u7tlhxx8xuz01w/uarjaNnaLCKftMC2pHPaTyjGWO6+t6xiZbb5flklk6LJ
aucr9x5oMWFSum9gZ2JTsQfItQphdSDqzFkgHoP0iIGTFc+cz1V6BAwJCEjv50Op
K3FV1OZldJC4xIBcayHWJVrXKcWNlRtIu7EN8fmlXEy2XNkl71TMxyEUyTtJSQ9e
sE2mFKFvhrggYJpY8OS7Rs3U/P13AtBHem56Xc+nirU6RxPPDt2K3mG0XbHNgdO2
TT+mh3AqnMICjGR1TRgD9ZgIk5WJK5scc/tZehc4nbNCtx7J37iuMbhxPDTOvYbl
HKIDtJeiIVUzopF9XTtMdRp5WeT3Rym3GvIMwpb2ENsfmQ0Pq9DFa9wOBK6dBlWC
IvN4cjd2mydXH3HOi6eqFKtQimwzUsbA+Ncuo05Jg66eKgjBNkfn09TfB+pHm7tF
B/WRLjO2Lvvfb5AiHDXTtGh8e6eX3eDBvjVOz/viPcFBh06A3uN9xMLQIxfZEmtE
n+5CK5GZ5qtQq+UDCu8KUfJfd2n2B3LIQ1FTq/fc/Y0UkHWFIqpor5b8M1apIcVU
40DJifLyPvQ04Q7qiGFcxDLKK/Ma/K8v698kc4pEFwTzs4eANddxEYPEOHCfBNHQ
vvwl/n0dWbM+dArfEpZvs/MkSczaOMZN0iLWpsll5zk3cS0AY5d52q3hiFxB2/V6
P9vnYmfOTENoAzSSVZ0B3onHr2ot2qH+Ji5FezQdGdYmDez/qjwmoKwuG5LTbB43
dpweYF6WbzLLzIuXSjOPVIZFcL9DeCGjQcJo5XZEWXmFobGLs+3re640p+5tTSp9
ie6e9Pi1Imuuq9MevtnnmrCqCv1AMXvLUkiRdlZZG8Tn0/o1n44t2lJavhtwTyNp
ZoAYDIrw2g/+GKWXhTureizSp+8gj1exXbamY8uIrqQEDMrlHP7wWIV6lN8syctB
u4AMwNMCmngq3GW6aAjf5mvhCTsx0aLJL7e6d0ZJx9nkkia84lOH4Fcy2UyPXN/B
eoxqws7kwSVKrFYWClwDCRBE914eOLZPoHagmvstX0lky0BShMLkOusV6Ny5au4H
6mQ5C9PssOg+pvkvAjgQWEbwB1zYQ/6V4NNh0oVcEw7k7dbBeWGEyjZDUB7Ou0aC
TKL27cTJAWXMTF3eoFhoVQr+fT3ZUv6I1BtwgTD5LZ325JpKPo3cIr03jNpzQDcx
LnyuTI+wBd/hHETNNQP+8VDRsehxguaS088Mwm+lw/g7vnNl5e6JdQAKjeSvv02z
nknyhK3MW7AgmY7ENU7bbNXGMCKeyFF0o9v61R0hsIFBWqkHmHhD5Hr2wDQjj8Fd
0v6Uhm0He9V2G6W+Hx0lz9ClwIjM1I/wctZMAgHpkMpuOIKC99s2UwDPlT54m8bD
W+EjZ6niCT2jz9V7eJ37JDMbRdJKyr53ONGnuDngFYmTPjn0YPEL8hWE0KRghxR3
GIC9b/2W3UT1UqHfFPE/6R62yr17jh55/bufiF8cXu0e9+96vAyAR8LW0Z9Zsji+
/YdwXLVSt1bjEInDmYBPSfvxNRdhtlis2lVK50m+08S7/mg2xrLAvngk7QqiW7cw
7BquSKGklmETbswnij6kv41GEGsIdZVUAfWkzwgygfPSsmHkqBha0SR84FukdPPG
YKu8fQhg7W/4WpeCTvhnnAgONf25nPuS1DBMt2K4dxQXA8ZCavCyj5TJBGGP0Pf0
4ton2cu9P8cftomdHJ09QmKnSroDjvNagBZoE9LKjFMX+Tza1YP/OqNuX329DGkd
2B2hlv/AMFic+y+8kL8rbFNH8PxiNKrEuC1OBFr2Myd07BCnlzdD180EpRK0bUpv
jaChGumuUBnqZtfhgLKrECLt1Za1FMpnPL7n5afZvn/cnlC35dCSsHfpjtcnJVj+
AfdkOe2LQq8Tm1kDsiZ2qEsoA1ia6TasW4gdr+nXIQPHjocSiPa0i1VMWxHJYNSd
e+AATWK2FjpssB2qFbcHIfjLSfz+AyLyjWVe7OcX2/9MN+c5gsGWzdSJKVl55RDx
DOPr321sIDBGgL5ExAPHgnv05P8A+u5SXeojA14JwYDsNlAwujRTkJk1yk+Gh7lx
UZMGC56BMODgPdZmoye4eAyw2gBV8LNtV7MR3Xme76UihLBQRO7U8RFC0J5ZPZ9q
FGj4PX62eO5eCgY+1Vb1pyx+ysRKaxEzoIFljaCPPHUsPRvctdBYvSSFPpGfK9Mw
7zb0FCUgWTy2jwfGCIe26P7EQwlnlDTinQBaZNGg0+tBhCDdVX1LT3Zx+ODD/O3d
m5NTZXQ/H9bpAZZTB4vMiy/8Pr+ethIu0V4T09ubyvns/IstOJ7SmzNPS1AwOFkk
1E+5MEddC6WbM56rDS+KUcG2wztNVfMoLtH7HRPiCWZg6wpKcbGhr3Ya0bUt6BBb
eXLhkkc/vEZKmh4XY9Yy1EcFsv03f1HNLFbPDIZkdDT8qKKxj0t+7s7YbHQF6MOv
lDtmYn9/Yr43VUtttHEfGxk52gEhuLlLxRgbKBqoHdYYHKVQjsWpwx0GWC7Nz2Tl
A4ox6/Jdf7IUGrSMtZS9sY2xWgjRSe2+KzMLEatnbcq19DWYdaCPhLlOdjwlOyIu
ReCN2gblmZrXTZBW1Y/JI8fdF6x0w1fpYH3vwTOmq13XxaNdoP+/eVrNjDLJBVM4
MR5jydLno24OdzAfY/wVUNzJ6RsQQBBT6RGUPkdTCAsHO5KkaVyBY04GaCIDV4Sz
5GPvTVvxWdIqIQpgGjzMsHQcHJuPBXBmYqCbgmuE5SC06jpIYfUkRo6MOLvY8wo4
GctmRfKKX3y9efOT4FK3LeQsFcgm7XcTausbkd33QX5h0MOgSEzDTQY4INkJCPvD
PRgdXHBqSGoyDfB9ORVhYa1tFBK+wG3PKa0HVEJTECv+L85De2dJWfKT1lBNvUXt
h2y1Ilxd6MI1JM8QUjU/ZDRHw/xYdYhJr+WXjEux/7+IDUlGZkt+MHnKilLonUXn
5Xd7op51kjE7O3h1aFJ5DLbSgppA4D1UsxT6z17z1URPkp+OxYq9Uvo7vepWxH1j
b1a3jV99ygZlA4BpmGIpPWbpxWs7swUqjJdVGD3ECiXd7Ly5iTtPpT4Qw3/Kloew
t36ffnhxlHN+q3gB5hk4oR16amjjx8kxb5M1QcqxnjGQ/80Kkrujo3HaeEEpd/fk
ilxk2Af6VjtXPUTVbLdhDevgJUBHs960aFFGI/3rNcKZwvGKtg16VlHBdNT4QnBT
moMVHVBFlNvslY9l8fmILUhxt4+4Ntvo8p9J1lcB6rfdK2n0bQjn3ilZm7X6WJqS
+sYltOQVRf87RVAl/B+m/w5jol1wBxmji8cGk07Y7PsXKB+ZntQ4lUz2YBdXDxX2
ssCIbiqVOFlSQU7Ma6wA7a+KmNayDzoZgsckDjl9NV06WKkHjubxKLh/UdrqcIRE
ccoV+5XyhUdNnS5QsL+KW3gF6yuQRhAoEgYJiipvQUvIukk6s6lGw7ZjHrN+4Pi4
e0LNRIXKtM8ZvZbyy0J2MT3x60+bsrDQ95Qv1rnm6+fqLrCrR1PO9pjRSDUsuoAj
fjRbYqjePYCurM9BV+7qOyEByB/s4jh+7/fr1rj/HbnPS/i6sNgkRuk1C0QXv426
FBWWuttoujGFKHlCKUfJzPNrx4Olee6DKD2AXTPDAOZMX4/5yzweVsYt72DmcwMA
RJ41UL07NysWcuH+RRU+nX5ypht7EXEZFHEg4d1e7FFiLJ2jPluvkGuiPhNIQzay
b6SyUAT/Qzpa+WcZN6h0D3PHANBkpr3K5INPOVDoXoU9AHSFGivaVmfGzfl+EnqK
sMv0Zkeli+7mZ05ianKDpZUzC1pvN0hrPtQs29PRUHVDAmJJ7J93lNjU/cpYvv98
uLi49ZnTVhpmXMc6iM/R8gl40eTs7SeMQQxOdCquPxVq5sjtU17HN7ca75eF2uaK
rlNWvIlDQa3W+iPTzSAkbebbMwNVW+DcLtuzIvHpzf4T3XGhv86nJmhw9kdYYa2P
lt1A0EMgg+H/eRMA+sk0tmjoPWvGP/4d77E1mFuqn6BW9MjVtJYZcfiyHShkOkDV
+zCIm0+648NTqNGmOydJHbLY2zeuw6HSIgunq5/rEc4wc8upTnvAvzxtlMi7S8/I
hjBYW676o4zRG6pyDJ2Lj9lXbynNRz1m31DQK7eojlfM8z3lXTRdXPBKJ5BnhKef
ThG4y+oxoyhv/yPR2Q0PJ6I4HSnV8oan4+LI5nPNK5oBAhmgbVMEjvKJY0eqGMUQ
8Ocju/+SXo3HP3fGh/kVr7Gq8NDfaXWvLEmN3opVahoWJnlkJQUNaVDu5nLEsmfG
VREwLhPnOEqVg7ymxLEtJyfej1SBDZBnxfWV03cV/fP58zodGZQn7d30+BgaHRv/
m2t2vNQuOt63ZK+qSsERTRxtcxna7zGCXYHuuyU/rWoG5H1w99Qn4YpM8sp48kIF
icZq0MB5MMBUrHl/rC2JcBDLugyyo5DTBCeZgnTqLgqB/lS1yNOlXPXaMI+GkWen
nXhFNhGJCac9IAM5J9vJBtRuUOim36qxEInOjohFDgFKxP8WHVeZivq0Nz3/27G6
FgXXTSt8kbhoDBXnK4Bz2P20SPY0G6jXyUe/BCHJ1C9wF8J0TGpriBB5pL5drT6j
fXTm+Tp9NGHVLs7ONnFcas6+XDHJc/57dLGygYkgYkO+GmhGXaWMMZKaa8ybLD2o
HW4I2Nq5MGsxNTInWDSoqskAhAHQt0YaLFOQp567/NY9cIWb1nV/891qPZ6CUDkV
9kWyZdzyEABEZDxrsYnnsYitcopbQ8FuQskVf+HFmPKphgZ7v/bkNmch6+R2oysu
GtTldsuaavsYpOf1p+F3ms9kWqi9LlySId6RO41gTb0rFK1lI+5batXSQ56mHZ80
0IpIRrmA0qadEWZhiKcf7ihvIJl5ZjFKA/uSH2pHUNfDYW27mqj92Ue2v/US9LKe
CBlOtk7A5VB5xi+AmD84SMlXt7USEzIqNLRT36MIm4qT6gp4sQes3SgacaGSeseB
094zOkUIeUetyBHC+f/bt23DdDYPq8aBmVYduvijQkopwvtb7FxmjgFDNgo7g5If
u6BlPxPZZ9EE1uApf+pieOe++JhAJNBxk1+YGzsGs2sUFgZFZcEl61TvLRK4ye7M
OFZoZb9SSLrYG8wVa2n86vITnvw4lqCJtDA2Klz0+V4IGJGXUh5k+Pp66jnGZM3z
spoyRjJtoXPRp+kMUURuBp3dLdEfoXi7DvZSYOrkn4oXODfU+3ONtuI3C6txQ2Y3
fAV0ovlF5qpFnghW7GkFfLK9pfo9eHtvbNMcmtLAqCNb0g+mUcrZQeUOc4rBt9/L
Bv0FMfWVA1d+qe5Yia5nDhJW5WEtMNs7rcOwiAzfzO0pvbMkXzlqpkRGorGlhk7k
NUxpyGzJ1mBeHev1YsGUhUNM/y5tQrkku3DuTqKGHmdcldDTpLNC9C4dP/7zLkTF
b4VqMMfaetckqgwTl8W0jBI6Y7fWPlonoc9BzJsbrh53SMxFGYb22ukkiLKnlceG
gH2RS892ajpS/zzUfK6R4krpAtaxK6iWrKjoxHTZJWpIJpGaxBEvmMvdqw7Q2+nO
U/pKuDkf2cB3qw5HL1XAL/xd/HMCy37kee+W9AeJf9FSdDWr41MFcJ8g8TCnC/yk
xH1MULMe7/1Bhjq4pEO5rf+3QG7L/NeqWf8F/gZeZXs3oL6ICf2FuOo1L8KtD15l
1gWj7RkkhlZdsJvdHEzdmQcQIrtFmroFY6U5H2QdjphQ1B/tHvKmvFhBCdNxgh3K
InaT+HYS4ldcDCIZBP6PZQmsX0/hN49nuly5cQN9jENOCFpo5WMIxE0j/KiZHnW0
YVMLVO7WEs0O49p8aCN4og7S+5XTVz3GE5YdZdnYd7gdOHQGo/QX2K5pRycO5xdI
B9AhF4Mh91OhlwJEcBqzblS4+Q0+3ShqQIhAUsLdnFjFKvuBO94RL583EQKuBF8D
Jv41hrV9a7gpxkuOZuYGjGNAxDuCXFLqRYvTyLSJn6+oyDs+XDdo3LEdzXthnPXM
UkVRX6ts0N3tbuj8lmA09yoxxa06qo+FmnZB7GYRuemV0/yQPaLGbm3cNtm8Yyr3
8BziOWnD2VWJjzv0KKLC55wN0vPwfxXLUMj7Ae5eT1l2lwhhnAcj00SSK3K5rIGK
Kp8oe0dQ4OAxfLF58n21lPKnleamC7Y4o7bS88qpNarSzJNMA0QnA6bv04vvNMdd
TxnpnhtfVGdM1PmCvLlRoqqUXytM2l96ZRz3JgZ/fEOmyM9C6vepcFizutuiFAZA
tuWcO21CDuoOHi70KTa2ZCvsRrD5wbwqkQq1V4JuJxkUx7inBk+kx1ySm+3+M8J/
/kLMuTJn8AKgTfAfJwklIRGZ9RTq8f3gusyFI+/Xxd4rN800lL8+JLzjqujhbvpw
Zl5mr+aSiV9F0lm7+D/7egJefInneeN4qiT6d+Mfp04kM5cvG/Q/B90YfP9Wt3vE
Q6OhJv0XBcTLjVZb2C4NyxVjGTyqhY19+Oo1vJIjm1G4MjwMQTjBaXYsNS0pNFxe
4FLfVywR7TQ0FqWCnPbuAr1oEkB/XoNj8ruNs8guTXOcCSy55qGaUHBvBo5KQnYg
osLlnHMbwFgSGM61D4nDHuTsGoOCs7+i/ZV3d1dHrpsFmNVDuWpWRACsS3IQ84AU
0WkX7cwOHRWwSfAJLKLggr2zE1RqKmQd9Lopne6tnbJ7fU6S1+jDhxdF2zQubNd8
9ZV41/NzXoxbEtLVU3KcgiPt9y/InS90FWhgD45iiccxKb9VIMZ10NqmhhUacI5j
d3I5iH4Ua9caBGZs5FrkHNHk2bvSyyKjX74VGjf72Z0rrPUjmw2wCA+Apc9OusvP
B0oStom7ewG0+7Sp6DhAvY97XgEgVSGTMCpSdbK8aRK2B9LBWUrgg5cawcuORN7V
+EFeQ58pdtJzYZC6L8x8Qj8ofV/is3qtkg03ESrXBzLCD8q195pokLZF0wy96TDo
lerjiZtQbDH8lHqb73/EBInmLemlT09qOo/YtVuqRITdosgKqbhcQtn0qrEuVwsP
CsDaRiU4l/Bz3z3IgSOaTUX2XeORzm6lF697AjwZ0/UuqvVkJM0VzbU687ltIH83
O+VmgpMKFOiG4O5YJOgjNySPKcltcbDaRphyeohAxfpdwlNiJlMDo8yd3H6ZpYs9
isiUsHHcJB7ASg/WOlaKfXT64CLEaxKDCBivQsCS85OKW0+o7ISQ5/JSbtdha/xO
JVKEUQ6gxPJRW1Nn/wR2zp7kvyKa3xCPSAgk/Pv24oLl8VswVX7uQtDHRNHrPrcS
EP9KeXyWHDXp7rPyDSsyw0kMXjrtZWVgIWMExIo3Jr+wQUnPp9K8xlf018ZZ5/9W
507tcskJ3jO4tNcMj9sf2SSIDvOGg2oR0zszUTKr0YeOl6CvtTA3MHeeaJH4Vv/h
hzphmU6NHCDzSkLJger/RWvjxLyY6nHW6DXjnQZxa6srscJTkSZE5ahE2Wawgr1+
Bjv+pL6vDSPiMhXtGfRtBG1CezI18DLmD8Y2xDbhXEZcH9FavIYLLeQgeIyvJgk6
Acn+7zBplXeox0/CbkU7f8PtRpOOVYVv0Vnlmm1esEofjmRG6+gxh8rE+JD4JGKz
BuAuKS+jRCnOW4paEREBSlBAVkJsre+PQmh3gorvhJSiTs7Q53Ok22pMjf6PtC5D
JkS77iXRjPvXBkZUxAOqeYZceqfrXHFxojdoPD3aY9wR7PNLcDKLDehyMLtNkeDu
vUH4PVYqN6xFLNfKXaJvpIvKLdRBAxk+5pKfuuax1V6/D9nK+blYrewexJ1Eq+oP
A6p540dNuPFqsoOKizpN+sUyhEDfaA7lUaxod2fjKeOa8t/0FmjBIignem+/Lu5q
6cLQxKQwnW3pU2pwKtlxaynNqDZuu+dVlVVkeMgrSr1Urbict+A1tQmQCtju6+Ve
o9SccfqHthiondVM/VP165L0bOoXLYHDt+ImD7HuLe1ORYOhq8EVcy721+PJayqX
uGrDuQDaFovKflCgPbBUybcIT/Il+jPi5MmTC2AsLFTPvQBuXnIU7NSdNc+qLcO2
5an7QKdApnqrDUr57tPWVnEdJYaCP7cm8n4Iv2dvc9DuAyF2cQE5Wubkkbi1cnKQ
N5mXeZIX4H3NADgScTN8IDXdugc1Fe0QZrEVAuTIKQUCcTBKxcrH2BFBTVS8UZYx
iiBOJ6J1uxi8fnVwCjvkZX7yhkUVtxkANQKJVoUrtK1VOFbKjjZeU2L0QVXjxOvH
BODw8lt95UHxhsTDUaWf0gVJ9Z0IIVhV0ZzKvw2iy/3SyIbXe/8j7Oq3FyJAwYiv
m5YHlUv2rwlZf41GDS48dSnhadgKIpXZdxKIuaeH1hLsqVUeTsLiBldG1gGg9eir
UxmLn8iURtbdza5TLW/V2BIvI2wunPj3ieYalKgJDeJv21jJySs2+oYuBVdGF/Fv
G49VFDSIVmM6l8arJRt/tEm06kjuC3gFI+TZQIMmbxBgIj+2xIjWWUSv/fGO/DFr
sf/JuyLcW05qTz0Y3IUCT3MXeig8N/x4PsdxoyrfPvHIyXzULMzGs68xluE+50S1
Hf0HRbMCC4t4jMqRm4YujRRVSOU/q2pmFfNbHWOTEJ2f3G9QNcH6Rp00brDfNoi0
aXIMznRqk32sCSRxBLwWlIpP7fFuwTzO5WuBieBcjSyNmdo2IK7mxySTOI1yvXwH
nQL/HjM58CITeVsG48413/aAbYFOD/huUa7yRvUbJB/vxAHt/RtZvcqjy8ARkJCI
hAbsjn97GsTPG5wK1RqCxeKGzcLaQ9RjzJaCGUz33/sqqAhYbDR+juK+c+UcrhL4
ooK6DCIv8WxT0BguR4KFJVtgoajiJr29FLR/VNnRGs0ya84gRj9B0fBOqS+46MT5
n8mGMf1fjrwuu17lrC/MKeGoe/GExhLLTVo2D5BjV8jIKlzJGeqGSvJ0f4aAk5uP
2lJCByfq0AAUT/U9yrSYlhahEDyGSqS6qeS/79tfArwbmcYWUqfua2Rab+tAw8GN
lZFzCTNPoO9Ns7ci1v6f3osel5+/NFDNqiFrnGjlhqp6BxVMMov3EmMXAlKi+m/I
YduiybEvDOchnIjUMKzLqwuZ2WlCd1Fth/4CZtY7yYIsaGSSRzfou641O7jMtgEE
pAvbwcK0DufpZtUT0846RWe5PDQ1cXJaNgUsq3RsnvEP0g+8uQm41eJuZHWhs9jQ
2rvnP4ODsdOB/H7HBVzN1PRypb+PTjjJIZ6dEJCH0sYtHKJ/ja6wV3nOIkcw6Tjz
+NIna96+v46Ta3Y6EoA/fM/bBvdkz2FTHEzfCD/0YJjzMhfujg7Eq1nwoZz3XVDd
28uX7NuK0RKQzeenk2O/pev/LLcMNDjEy92UftfjW6q7jeXYWQLifIprTp9OoI8g
RysA4Yth1tKmhdUWJcVWnoPM8NAmXiVEx/WAEOk72pbxI8XQovIHUL8Iy6Ru/1aM
5xlnpsKlqqAiF5E8D/D9lWZUUf2whAINxb1jzeKbLaDGwKeiW1RutAFzSjRsqK8k
I1jb686Intc8BrlJs1svHam+oHcbSi4vdU6Dc23wjY9kFU7eKSyuadeAaUKPRJrg
LNI9xfo1ZT+boqVz9syUf++VkaBu5Hk4Tk8c1parNfKtQnAxJRpGrmWg4QonBl+l
ZCu9QoIKjS++5mNJ0e/dnZHrOYDjd4Iury4VLQTVmIqiJGQrT8Y3vWoj9wq5uego
lK369B42YzfrEsUB9ijUJlvPbkTpSX+KQ7OFAuhgWNn9JLcHHl7VF9Uw8x+32SqP
kUbe2BIcqMAmT1kb1nD1rHQ1Hnn2ElAcPHGUcRV2vAvFWDI3I7rxHafklaQh8LD4
9PGeFgQxBbAF+q9Opkq99oUetequ7SmfP7PYC3M98YpshTSEdGxIY/WEqqgVCOr+
w9qGkcqzktU3mj8870FxczoA2LyytzDwtuvc8QTRTGjxz5d0N8xxc39Nqukf2lkS
jlXHoYSkWJLb26nwgvXxC4U9p8TmRepzU+KxacAejRymasehb/YuPZIy9L+ce7Pz
Ldb4ASxAguArlB9y4/D94mH7Tj/TeQVNa3Rb1C01//zBCbcSdbWgChV1tG/8eN7Q
lsu7zjzF9P+4cymeq5CvHRyRchOHAsjvKyKj007p0YbiKmRQr4/+h2vlRuYNks8C
naSAwmTui2Mygh+j9HVCMdxn6qB16gILkTnw6B2Cg6s5I+NKva31SU9e3kAnYcVt
zqw9BFtKErEji5bvlwNu4S5TUdyu+33gyIPSl+CHoYX9pJNkGJA54bvw10Hdtl1K
Nm4QZ93YxhIqRpYneSBku8r6GCdNRybaPgEItjDjrl8X8oXB2PlotkeUsZXifk1g
D97Dw2Ka/hn/c1L6Wcw/o+EztZTMgYYTM+xefHYl8SdbP293CKGwdDLzRQqotuoz
NqtIONMFmdsimfXfiGoVZOpPZijnxvmFvMfvmg/RYbpIHQ87yD1dF4XHXwv0H7Mc
hycIKp0jgQd86aR42xyk9DTnAqWCWT1MaJ15R5s/gdjeuBlIWOe5OrL0vwDBjwoC
/qWV5bu0nJs+du6xB4hb5wPixlZ0j6Dc0/1zQBLPSBEq5fCNzy2vDqLPPtZH4y4M
uqW3ZyQ8l2aEoFB1AQCfH0GcgHAB3z/QCsMOX38aMR8GR8q2C7WJCJM/QeAR9vs/
h/tdOayZyoP6Q64YWG7nzwrL0fZuytjfuAt6Lni03WgrS+XQrx+L1cnFxgjZO5Pf
r1R3B5xj+66KkpN2aJf/AwNcTgRaaJtRcf+yO3hhgzPXefbFV5hvrrnqQ201c/Ys
+H0u2fw7e6bmLanFKne73pZoiCDDIZId5XCHTzS791dWe8s2KKGyMPQeYCeu1w6Y
e8lTWwTilGQ3g/o+PG9igW5kxWAa8qpBh5piiomuvrINgjBxZcZVybZ5XmmTktBR
GnYSXz0IaTdga1xIgX/U8SKb2xQSGeeR6GI1qu0QnGf7KHDggHhh1eanUKv1DS4P
QHSKkplfFDgb4T8f77Kqt/FHVbEOrKQN4o0HasPWdzYYO4OX4DLAmNTmDBOk3yvK
cehxQt26zIHpoM8+hIS7tw19ZwmSydO1zkewiGsIvLmUFqDXBQ9K/lx79s5GY6Tn
CPIqpaV5ESEZamp4Sx0d2znvAOpmIfUZsvyzKh6HPyuOfj+CmKbB0fotHdmNpc4X
2DpeX6tVqni8vzlYTO8pNfpPl6A/1EIqOpTfX2OVt3o8boZAKOXaRollCIrHvPE7
Yp90s4g16z5Eim+UBqXHGI1XzCQWEyCNV7qYFmcSPRdpXbiaOGyaR1B9Wuc3dNSy
3gOzs8m53BIlaNaJ+rDGjBDFsiTO4FFJfc9ZCdGxk6RghGDI33IO+HhjxdsdMIzX
1aBRHYi0pJPTQQD+WA9xp3imt3WAbTrc+sCfvmWUXxactL3k5jF8zB4qf6jKkyqw
MR1gx+EXsO8Su/I3aky/TXX0ymziw5W9AZjFr1XEAjhhWgAq0+NOI2s4yn7eBeT5
PQEROOHA9gv1mlMKYFwRz/LYj6/t05H7Ed2S7etuMV+OBdu/V24bCRCrNhaqJEYU
vXBIAMMgJ3t4I/+ROx1MGxm7WddY0baKbARg4jAguypdil2VJFFL5mc6NSbR06mx
gS3T11rVwL4HMKPNFrTglVRE38GxO/nhtQ1vyCvfYwWGMnrGr9xkfZxh5KB6Af+x
kprd5OhfZ+RmGMMdkiQRw6g4hUn6tzLW9jJKVKVHoTuoCW0lNIroZWxVA7Iye6bP
rF5Y8nXsP2os6y770w5ne6KwwC40qGVLFWR2hvbR9GCpmJNhJ3NbZAJi/O+k+90L
jhWVV/0NLI1fV7ZTQJpv4mpGveoEzIEkK3qGtdcLLV4KUAUTc7eRGEwJcUSDzA5o
DVZlz/KxbOFlMZg0esW99AiUcXPcUNe5r/azXo7bss+fQAIZHyviM2tQ1ymklRKi
w/q1e7SfYjBjglIAmhtY2DKaOBK7C+ELabAoXYgnL9kxyu2TsMgUY9Z/96JTboaS
ZQWALS0W0pg65BGfHZjSRMMgayyFjt9P32B8LMgrqTVnPdSm2oc9IKT0TaOlU7lR
xdwi7XXNsrLs8ntgvoeYPmsgqRPswmc8+iWSTwmp8O6LHXTtY5JPU08dBViMWkwK
Sz7j0HAMoXGiDgSlR6YJ/AAZnaft2aEncS1rLxWuxZ4iftXYM5JWy6+E2+qYa2hQ
4ns+MOQHm9/FrmmkaLQC1D8FVjjTWKvjkvdGXnaiv3QFB/SRWUaoCgCWSKHbOe3T
94OMfdl1vGall8HWX9Amb7j7JwpUsB3S/auDAzVGK13+pZ2eUcuYZEGH+7QKd1Jj
+eJyh1OYVrQUSxUbfavO9vbnyIxLqvYhEjTtVi+c+gJ78wXKXSSsa/09Vd0FNZjL
Tf88BRSjm/badX0X9oBUTJTcfR9zhqTssTb+jaZ03mPDjr9R9xvR7IM/tq8c6l0l
X3UAYO3aFeGmt5+eCSTY3aPQXUBqf76kZftPVUt47g3Unl3ruow8w604lQpnJARY
FQHLcoaw/S+8hnCz0nFjzyfONwxJeuUDhMD2e7Ym7NGseG/dZNTmsS7ZxBiOPyGR
fBGHSu34uN7DnXSHp0X+9ePV7mNJssp7w3jkxAVYiBHzEMqBK6f2nA2vSrF0g4FW
jnrXWkn+K2A25g29DUTs5mrxU1ZRdbPStAWnR3pQ9NpZFiwm7l0ZFCEL0HeDX+tj
VgPxnyeYNeY09EG51nYf0xYTukQj+WLx0Q+hd8bwbt3XJOm3sMTnrcQufkvGeSJJ
/vgN2i+nunKT2Nk0R2D+r89E6eql4DDsfw8p2Dj0Ztyrxbji2CecOSH4O2ci+JoK
cleT2xq6X42BgPAuXyX1+wxclinPRTFTGigKfIsLy2z1iFSibcFNVAJMyOZODqfE
hbdB632OEYuulpjptlEWdc6fMDXujjqU0QEWXHXl8FfxbhBwKPi/F7OV5jMkuXOK
2Yob30t86Z2WD9S2RGT9oCQ0qxg5r4zXLTLMWTVgZMFZsYUWcc7i2yqp8LE5n974
9V8C6RELRC795gjxZ+xeQ9EQpVHMKby83VaDgIiwJgjwB3FXjjv4SoiQ0WcDbGTT
fmOpzkvEmcDOv7j7JYTtkGxbadBBfH8rxZ7ypnO/8f4KcpmkGQY0mj9dBZjMTJ+g
EN02hUvq0RP3QwsqDvY5II2DIVL94cQbCiVju0Y81kCf1LR46BMtcim9CcuH+I1O
yHRQRlB/f12pufX0fNz0FR5HkTU7q74eC0+2OCj7ocbWIGWx5EqzXgT7HJsApuYi
QoURAlO38jsTw23eZRao9BOfpqckEAysKlN/q5RptMhqgm2oq/SIXLe9aPiwDR9s
IRN4JNLbKsMzXlaAnmvt/QXYQsr51sXRpmbcA6XeQLwoeMBUo5BLMDYpqF9zmKGv
FyTBxqUne4QVFDrRdLqlIbn+K7szwoHkW+PVPcAJ59abXRjiV9awVgPItqxnl9pC
659BQUpuzsf4TDfWV8L9cFiNgV9qa3ZlkAAbbbFKSsgo4B8cCma3KL+FVinvMfrm
LXSe/hkVoVMHomjsB/+NWguVyHMqwHwY3YPqoY5zm2jqEhVk9B7ZKa2I8r+Iqs63
5D5CceaTdERQCs9cN0vNvHkfgQp1EsoKsMeqkAXlRIf/kfMxss+EvnPbvDUDbUwP
vaQ8JX2+o84hjucSTkSWYmlKO4ZsYok0/srsOqYkzWklNxAlgmUBh7NQJqIUkAe/
tH/lc+mq/ANuVmcGmDOOBfSzcfqj2Svm3VSkWjQgV+RNM8zIFzwO9PWLzELVci/Q
+sBpWXedvFpbp4xX0Y/zUWyuuvnc2zaiJP0yrCwKrNXtlVqHsCugvXwFRruuh8FL
wHJM41mwgzJVVrd/2fA2U0cBxsLILMvk9D4+SrOojlxunyXPYn2h2lA1eabXXjvP
xGmAYKL3KuQbVEoWOWNKNOIp9zN7Hdar0DlD6vtq5VfLEOVPPb50rFzoWE8KGDhI
8drti8+lX25txDU4sWWGLZZuDVfXb17+dZk08P9690oDQ1bezXNDbFL+o+yHJ8zE
aCr8ZMqgxrOE0AYoUQOqP+tT5r7l/DwxF164IgiSzl+okZSfLoOHtJHkxMNFuekT
1GGZZ7LigL301ulDWUgAxTpyyIWyN42Ay1u9r0LrhDD3vZRcBEuDdGHl/Fp7bJYF
cOzJPJqQ6Mq74d4H2USyw79t1Z2aQ96te9xE1LPdBwzEqI7UMhM1zM45A1T3lcmm
zzea6lICL1NOS56SAztiz3ct+TXBOZ48bdSND/CbhioG3RF7t8BG8lzAJFiAzxWU
zJPij4vXaVj7nc2Syt/uGz9ZzDuKpzsyTclWGER/UdTjjlS6BWc+kc2zQEMwBGc7
/YglMhGwrK96xcQsTZUTIjoDjLcfpzF2zy0obdC3OUeY8fhGU0Ak34QBUxWnqOc1
weqA8CZG9/BEFSW1u1/ywHvZYzmB5d/M0zkPM2Hb4cVAAZ5sgzTHb3p/lxZb+U0z
AscciI3LOteWuwi/Jdqk7IgXLbQz+fUEiVgCImiRt/+fbvt5ZcLxUetd7dDij/sK
ib8mhO8TeWLA6GtMg39CWH8CSyy89zbOCQeVTlvDk5rVT/HNwuR17sWKzpbCsPMa
lFERM4UELP83t8pR0wJWx9KSkk0Fv+LAXC2y8aEVLtxMiuXgvTLK0LatEa7D8xKF
WPcaD2r6H1pispvpFn0K6Atc5h+GBoJNpSApBvGWXuBZQ+5cyh58aCz5mbKwTogC
8ur4eGwmms8ngi3LVo0kbojNyOpJS6Ni+QJsoxH/gJrr9AycZyi2/7VuL0Qn9XzE
oBQiZtIyeMGHULXCUAdgf4If/+cQry5WansqYGdioYWycobhy9F+byQH33uWABDU
rCqrwe7O1cGEAA4X8T1a8AyV5ZkKkK9SZ4Dj6EMtBL5nseSMZxzdTaWlUVcRkoac
7Pq5wZa3GJzSFeq/2niXsitT1eooNGsO7W6mfF82MVlyFhbHDzIWywafDmHavqBa
BiqZLVUdkqL6ea0de3aUHkfBdBQu0Yvl8m+XJI+d1APnHF/MMvpjHnLKPkTUe4iW
Bu87h07JAkdlFPVWU7pKmSky+xbztIL9Xyqmv5+/oWXEF1y/eQy0dx5pGCHdfplN
JSePpOL6DLBNgi7E7uz29v6bqblx5TqEYFUY6jg3qFCjU9Qnzb3dPN+K2bzlchYi
v1M9w62iRbtePhqOMlLobNOc+ZZWYpEfwqD0P2+ajJGlvqFguexw4JgEqRtGWtx5
S4F3fwWNvXyS22bWhBpIy6HQLPVFZ6zvSAFNrBnFT4RnIkiWyu7UKvSlIrCsbag0
ZKig4GzM3fxdjM+2lwTmBasJtniHtCdBP/aiXZ5pM+whQunlQFZsXkS5+kIxGg60
EC0CM7n4p/UVQq/goeJrdYzuLpkeqUb+15ClepTLEJabrjUVlQU+98wtHxtN3XqT
OAEl2lPvO3AgDe0jAxRbgwADXF4mQsk/OrkySSMoAgvP1iIJ/nswdVbEImgWuYCq
mqjN6LXo5CZ9rLSE6o53Lii/KBYwXS1VYQi6T/2FMW4XzAZR0kKGi+gzuSoE+i8f
PTzrWDOWbhNV9whzo7Ij+MYTCuzKZKbEDctYSxTT1arG5DLVOnh7s1CIY7B4YicP
/41jgrvnBIMpNhMWyYIQG0BDfX74c1oZzpPISBOXXbo/+ITFYck6aCT06+/1QiXP
hDPfe3S6utGOWsxpdbvPX2e3EcWZ2J+ZunZ+bKPXJ9x+L4HyhbD1y5Znbo/OIpb0
GW0ht+DrENrClQBZKWX0ZNdxHv/cyAa/NKZIrQyG8Q6Ia8793TW3YAaAmxKU5dK6
ERliav/UpeH/h7QsqhdgePvjnlHhsnMBsouvDvtwrXZZ9xKcRzPQCd6cSLx6GVXY
MVnrjbJVnl8iG/dHc+rfo4RLUHZOqfqaRtDjrDmGdCIkF/olFahfktZcFKpy1k+2
msLn88MFE9S652uXFV/1ApGotR9lrxUELrsF03vdvtWSSVv32vacyi4iMCXJyeci
px0tieTmzHYJAm6hR/h/n6qSBsM3nUmWWZUXXjnvKuSwVwGkTSQtdFjzmktAFzk/
9ukjoJcRzhZO8nIVZGZPT8QXL3+9a93affFvTCcBR0EB5v+xEMPAldMC758N9I+6
Sk8Tdyd6M3JbvJ078eCV2wngs9O1nt5qrOdrgDYHUYVssoJorpL2d29I3aRrUK2y
fBQ1RwuQpQi8GKXEryZwqzEr6Ggk45uj00946CJhctgX3o7hUsNkXjh04AlpF3J5
3HB7uyCYH/QTIdriS6lHoNV0zOBv3geBvSrZlF4Pg33Kl27D9zCH0BVZNqnhsECz
wfl23v5ZYd0L2YcomaACtNScpTKw+q+sU9mrDPvCboWZFdVBPYLZHudvjcgm6izE
DNboL6tbCMs01Ol0TyXzFJMPMNuWM+TOPlLThk0iFULxz84yx6uD91raP/0zGAqU
kcEpYnCYMnUCOs15heky+N/EmDpYVuqF3PQ9RVkxgSFzaZE60T17f6ANZ9k3dCcT
SALf33VyREjdvNRvGoUNvAlr8E+2DKa4KA496tMgk6nAJANooQynKfesXjbD0sbz
8a3aIQYG+Cl5wqZzLNVU1ehJLRFjfioyguMhfIQ+AWn9uleaEm11R2W1TrLyd6eo
M9wSYKX2qYLx6JVRTBgF74SLAibtTHlMfQ4ZXF/HG5lr4ER+V6CKiCdD/z7j1Wds
mxEj0y9mF8S9GaGkY4icJba4j81HSVAJOKSdqHqk3nfpKhZtWVYR85Z55Dm64jPl
Y9CQHRG2VC0O0Q3mokxEqpxl+y11PGcShS2ZeZak3EIutQPW1Eg+XQURZOwONGz8
KIWipLqrOrC7GiBp3J2ZRfiIYjGqVS0575X/Zwuh82bTuH27UgQFOaaBKW+qEte4
gxwo1K5/J4DkCTmXDRpHNpJt54H8rR1yRqnCQPDp73Bs7zYaJLot9ywjSg0IXcyX
jHMOkxtUD0l8O+Qu3cSO3ZP8kAhEf3OV0HE69HovntoUTGdptCvFXWR+x8PSjyjI
PF5o3vZIb1pTqN2wbjWRQ0EsOOvahCaEk4/zZbMKqpWxDTfTgyrY/JaWFpUOSLzg
g9Z45/Hx5Z6of3yYok/WeiT18/sQozh8t4OQQHjaFFBU3AFBFR7HY3ZQhmKx9JUT
V9Bgq2qsyfGwj6xXN2VJZrPI0mUmTocXKSkT55lWwQN9EhuGcHq/dWth3GOpvqSu
y9pxy0R8SP00M/aHfTss87G9sP6DdokjXJPVh2It2z/JLZBwoR7+LYIRZdDve9ol
SNZ6NaJOsyAcRy7EfBdgkb+DyxAA6fMJNLlrzu9kAx45xZ9Juz1Rj8jdAN56YimO
XY5TUJm7q6dyJ7W8hqktzAv8UXq9ROhQl4sBYrDN7ttr3L6OJd2dCY74YrkMqCHL
ekMVyYS+QBC7VqjktaM/j9Zrl2KSfNpSVTiIScKjhhVNtbkIAp4fSx1BTS9zDIl+
3Fa2Xb3MaHRxoWdlmcwfV8a0NcAYeuV5bXuUTn+Jvaott2A5lYOoJM5NiLWFoTQj
DduDH5g5rYIlTQvJlUXBXVqXqDwbzzYryFbLqiCKChuOKtlZtrCFd9RI5qTfNjck
K9fwkHYC5eImlWj9bUdw9DiVea8rh/5jTnbJOVy9upGIxEcbKfJlpL8qzHgFZHKp
mAbWHq9DCS8YnHnZI0RnOa8u408sLI4XJGgt3YPIeS06Ux7N2IHtQw/1aua1LF2s
fVkUjfGWUwZuVB7chqzFM+kh0WasmgmOmfWTSkbEwG63668mK0JrH/ZsmKtPfsjo
8/46AVzU50XD2hQv6Ri075efNp00S8HWcMB1nQVCwX1/xYoIW+8o//BYpQZ5pfaF
XDu1J6IhwAAuPOKtMb9jd6HFF1xuiEeChbc+4IT9WMzBY0c17SLqZdEqmRWyX7AD
jXGel3wUhVhjVJxKI6uiVOSDQheDmEmWAxcYH4T/zXtoFsTsWdiaIszi2hLVVarr
EsB76S1kbBrMeEhGpHCwkSwx2YDtE0/HscKFDEgGQwgp+KOGoKVZagYC0ts4Ds2G
hBUcat579rhMD91VEpyEzzGgAKCMzFKhpffh8pnGtFFAXf9EFPjby07+/UQ1J2aD
cQnRqzh4FuK/fov0LskrSK1fCQCeuUuzm9r5nw2luoy17KOz6vXkVSlMA1owpduI
b9jcnFOJtaI7WEWVLiU7eSEu3789cICV0R2C7tIM/0bvnTFV/bwjgCEnp5iN3Wlh
ZwirOxlTQ7/Xbcqizugx3ep52dYaPaz/hooBo1EC5UOsyE+3h39+ynEMRPYGVd5a
r8RR3GpNFR6M6gGnpvDGUDrrL5jD9tc37Ylipvw//5zuufNPyedKEJa59EEKU6MX
SlWjFne1CjqdzY/kzC3twTKMqQ2za5sRM42fn3MCbn8sOYJoYBG+ds7pminQWcCe
RlzGAIET6afwH1ciE1+XJQeySPU7W/nZG0OejxrXKEjZCsZInM15sZI+aoqy8/hq
K5gRD3W8UXPPWQezCaHvkqlUSJ0gDKo7bQ8eVacTccoRLUf36u/BVgB1f4FOLsVY
NTYhbRzAaRf8Hg4Oi1AeiddOEx3J6O2s0eamIADWXZpEqS6qUp/IMGxclINKuwKD
YWCj3a+8lovMWO+ghundTUbXbpvkihIT2auAbz0ftQGYAtPWJgKMaH7ww4k9EuU6
hkKzSPTrUomk3unAzpG5rP1bKfCrkUP8iYQvCuwzp2zQyJwWDuex6RHSUT+1vCou
b764ixJ02E9TtNtad0m3IAqbws94eaenrhPFNp+8pruVnrBBqURqGFC0miZaXnCp
brLukxoY0G66ihmRvdhnxqy9vNnlquuUJVKvD9sVws8ZhJgEXnlkGeL4vySmtXH9
r3yDVsruwucBCM8QSemSNF9EFaBF98DUG1lqUVCaBw3eh5K2qkVwhX7CMFZ1qlp5
61tk3npJoG3Xy3CzUaWtQzrkbObv6S4Dz5RLgDMBh6FO/1JdikslEtoX3OrzuQNe
3Z7krpW+b5kNW4GcXIaDRv5rNTu/1eZJMYhWf0rZyJGkNa/WmCSN+74PU6Ln0ijg
xxq1bzdS5l+qBABAB2bnXWkdHkZ9IBbm1RZpLE1kK/3S8/BXM3+RQySz9s22RMmp
bklKVrT9H37rVSKmRB+koSUS+RD1otvVIBuwzXl1vII/lE5iXwgARA1pUGij6ajX
0A8rlyB58JCISPvs6rFVWyiN1wZn2UNIR1fHCEO0ex4xBv+U3ZGAQHlNWisLKv3y
sDa7OAmlrjs5KDOJ72myehwgDcQDXcBF/LYhYKKegw3KVq8MWx7UuHU5iqZ8V+3C
Z4aCyPjzFP7ET7kS4cBFUXS4Gl4AD90q+GDuafZwW/CFgrFr/faayAcAgBDBl+4t
TUVykMnUABY1iEHcMdmCKxXbPjkjUQnYHdRU0M5N54q4RPWXZ4hAyJmWs4ms7aK3
f1PajGpk/0RkoN6AX2Ff3goxT4hkC+wZ+XhxLZfGOGOb7K/0FCTy8cht3v0QMSxe
lz3iMamTYbYApgHIscBNbK10BsnaRYDeMOSkpNHSQHvjZ17BEEJWwaU7A3izR/fo
N0oSzsFXu+XRV1YvejUrheyT3osuVEvgY+ymQHbn7M/5rAJR6ty6m6qv4UYBmtnx
d6dy4TrAifWPCvJ7OAs9+PrSV1GeKRDG0LStYTU+4YEdnlyRJm+99Pi2ami9/HZ5
aSqIvh/6lojhjN0pzrY8NBswD1nTvSC4xpDe0dGy6RJP1ZH8OM6uIKpdXkE2tM/c
vywyW1qL52pUVtmaPLkmSVylgy273ut05h2zo1ILskKuJ7OwPkRIPVDjickQtXMz
1GW74cT28adI82Hsw4Q0GMaFYqayrgqns7/VyzVBqHZ/RQebAgKtrJEbBmnjy7j0
rhS/Zoy1f6Y1L445RMjB7wvKdirYXAnFO6Pm9UInNW0EpCa/FexUCUzFEZ1yafQZ
PLBWVN/G4fvDoUJcjZfUeqhFdTpo6p/JZdNKgmd4hjOUAOT/g6PWV7NAcMh2CfPy
R4Ta/g5XFlmlp3tz663KukCMdY/ueXydqiw0P8O/XV6zPc4Z5zzG/i9VTBSj/W/i
RoVyQygAfOsu8DOm0P6AS3UwOY1fJYTc/ArhgrekOTuh9a7EpWXpLGeNHF79sr2P
at89o9mcn+mt7HhTSYB9flNX2Rsulp5sP9cXGVJorysuvG/r40/8Xi03p4/JZd1H
Pls9HPDLqq//0RBEP+BE5JmMzvlInXq9YLZh/Sr/uNTNRJc5bDSQDLg4uiP7GN0I
uMJJ3kYKeY1Iy30IYRhYO7sbQQrz6tEpHobQ1/EGlz1t34YjHPZdT3MB6OHImi9U
7pQICwSCxugWZ34Z947o4WdiuRQFhIGt6zJjpynvya2E+0IPQelLMIpDNg0MTHGf
lDl4R49rostlMW4gEYhFRkG2zSlpKRu4QVekN8wUIVcLj1Cnnd9M6+wyAGaVZRDw
/P4ITetU8AakMoz9UIhgoRHbFJ6pPPqRaQuDcJOjYPc1K0p7oQ+xQQfHn/iIEHr6
zbjIkIvrqLyCSjKeS3zXjrYJgxf8Svzgl/xmP2TUEED8YqF+TfreCGDQn/TWVynd
vGTHdjxIF1x5C7UvREUqxxxxG1fNCUhvle7itWlUmQHZ46lOrg1JXSRpdnXI2sq/
6oZHcBb8dPvmG+FGCYqtNjuxvPaoKg+uYfj/oKeFTF/cDhwMfhSt7qXiAv58cYso
fLwhAnXTejofCu0vuj0v7nRkgGTS2gfAXn7PlCYOcCKidRhcTft2qe7ndTtVQ5iU
l+zD7d7avg7B0MvTOBzaW5GhOL9+Ri87/f0/kKyIcolp4piXXYI2OIh0NjgXzsLd
r6rmDOnv7koBXombLP6mLfad91hMl223YRUHMhUz74EVLkvsYrMfAogzI5NKwucq
31TtFHo/EqvZ77gyFRiXqSDjDgN7wyXjmJtA9Xck+4zZEcsD50PeIb0x4a/lTsOw
+3uCbUrWt0tBlCm7YlT8dj7Uy937ZkcZ09Xyqsvw7wigbJGHzp5GZcAM9k8GYN6o
hiybgG+QmwtQp4JOXfuAiaIYSs6jcyB8Vl/qnycLohnylsCxlQH/wGgFCpQK84Co
cC/CdoyVjq4inQMRX6laz2pSEVa3FWTJ+BuaohHAFNJZ//01qg51T2ilQGhqSVFR
7zBREnHtjQ4JFqBV7qSwzOn1LMOCCc/+ztwUBpJKKdS4t0QAIIcLuNAuyxCBUREc
IfsVkv1gLKN3Y0NOHsR6MmDqZgQMpE/MA6Ra0F+zXKmH+eVg1qb/g6nXG+HlT9Zx
ovGZM42becRcAEXfBf8JvsdvgUhOQ6nZ50pEItHhcJ7yQK/mj05Hn+gHF4uG83jj
J3/BBxHxCBK1JxzyV2m0MLPLB/RuqHRco2ScBq+5eArj0Y6wJrYL5tDII7jbGLsW
vKZmRBgIbDuf3JbWorcCR7eUIvlQVl8d/wFXun3xx2ZjyFRp93GoxN2f1529mAM8
pRa109ohZmdWZfj6t9j8EqxMvfl8ao4OAhF0KK0SPOt8t5U9ie7I9l6MpN9mhmn+
9CJ/IVvw4vpM6yjFr8x4p2byp9+OOimeA0BgunzALfqiI2K4TFPXdMhPVvGvzEbL
4HmIu2OGsciKEXrdNMD4T2hZ1rjjTIrbznzNeRNzIJNR+xzhjiYE9g0G+AdZa68x
29UrTPH1AAfjGzZRgVc3fGwHojIWNHS1JRtw6BO1Zf5Fsgk/bLP1HlYoC1nK88r3
9qXTfCwcAjhS8BjhqQJ6GHLFcdf/S9xPTBrWfYpiwTzVFyWLo6S/r/Ufw/kqK8uo
RVV5VaUdYq9N8pgWtkudloGP7Z6bVXqwqJ2MlVa3aQzpwv4Hh8a5BAFJ0gBw5lag
aZrJIanCOs+hkmzoPaXhe8dAL+Rf9ZtzXCGUvvXAlhDjqUTFdI/iVoi63sW6tMES
yiMilw4VPR1c1lDR4dpSJYiBK1cEwhxxJ2MW3zACxibu92kr5UGEXn4Tj2bCKVgo
a3C0GdmaEwGW41JAU06SS2f0z54SNNT0h5hG/3KYFpi0yp3hYQ5dh3VVOEn9sqUD
5wx/LN/ZUJ5AzNwcNhdktqyovqmqmkAGImHRW5o49VY9PC2ir5wmW6RyxnOeGmeL
4P1gXlpD+xhvjc1uesZyIOTjyI2D0MUuy6CqE/AJJykK3oBYYg6xOxyfs/TK1a6W
y6pgJt02m4Bw2CuFz2u8sQ4xdfvJC8qflJLhP9OFzi4H1aDKEnSzqoK/UTHdny0E
KA2OJD6yh5iFLCbqH/TcScfkKD+WjKoOWD3YRL8m81qKZ2oe1TSAb3bIm1bOBIf5
9LsEmnK8F7u9rL4pPJShndqvHQCRevT8IBlPuKmywtoyyQwWq9YTD8Oc0u+hnAqE
U8qlQYpQ7ffhKjAp7mJIP89CN5JjD/Ov0Lp3rvWm4Aew9z8zPpUzwDFcc+vQfzD8
OjYIuGBugKxfej8adYw9npn8x/SApw7Dbxv5FcPjPY9T8lFH/HWij53iK51efLEM
wZYMd7xaev3m3ZM7UdhHCh8BlRG+Algg2SN3lBfYE8rS2sBBDohzzfCjREtIdMUg
eJ7l5G+AbaHB3d1/Nno6SnKwi6c9ML/RYYjjoAcoJC85/Bk8AKYqvqFHFTM/u5PS
NUccJysnFrBYW3/Vg5WsAqR31faPCC4kzMKB6Xg9HJwRIU1Y+btOcXBiZ3QShESj
iOJO/3Z6l+Edd7Vp11bIKj6r7lwEXdZuck1GUbPmfxTxhmIghRK7FOpmYoVptRNZ
e2/r69OZAd3GE8oAiJ/lFkqWdDa75U04hdjnIVf1PwAc+XS70FysK0b9aspDaxWE
Ishmwy+2AcOdhvvRUTuh0VtQ2Q8ZWjzw5HoSXf/07rLBSL0qmlRz6Tz+o/NS6Nv7
mZghAZsKDwN33EST1d23H+czHbyp59gwYBcHIilOpyTJIW2DG9Zx8hgJh95OUG3f
5bPJrQMUK7+15/Y/1oKVKobTvwVNrtR/nvz+3JU7Tg3ZfHbzopqW3URYKAIYhiUF
nwm0Nl55zbHcm1LqU0J0Fk8kEkJVIICf7BYkyKQlnxFLaj0Z7TSnpWPumq9BqsCJ
yX+xrNw5+X6vCy4ykCWi+mE403Vg3j+GQS1V8WfrLPWLlcsWoeu075Vr/p9uwTM8
8BX2vVQNZcmeMy7SWuGwcujzy1Qj6r4Ejqwh0+z4qq/3ojJ/WNyI633tiMRuwKYk
KsBUtyte0Lg4Z2DyHpjUhAA0/8skSPUFv7C9WLo4aS/v/bHB1Iew6LzHncQfqHF4
SrzgamlDYVvK5t8by8y9Ci6t3/IIAIcDHuW4un2e7aeI/uVYqY8f2rShLfxyGe/Q
8jL8zhGDeAf0RSW1xXWrL1Hsn5VI8Ou+ggzrwAzd04MBBMKJ6aLIHxcYwcTCKVJB
vqDaSP7XbkpUxieKzV06jhVTt7TEdBaEisPcBBJh6QndHX5A3mT5YwduPMjHztkg
2+yCmz1bMuxcoGwrcNyme9f7+m8wVKelO2qLG22mSw/2ntHYDvB1WSuk745Dcr82
chuyEEsRsIdu+PsYZ/4yDlk1b302DqVjIvxm9fiDiPH944HVcRP8sQeNYlhTaDwO
ZTb/TBUaHHkwBfYJJtLPH5EmR0wJ6iZX4sW8QD0h8pDEgeMrHwEmPsgjPHt4EpV9
TWrDaw+W4DvlDlfP08dEfnQlgJEb0p3pz5NwvfAwuicX/Ri8JUEKMu/EGAEJkVqD
g46ktHY0Ut8ofI5ktspmFz0PllEGe+hFgF2CCmdNR4s/BT38iUsro1v5Bzt3oGs+
Z+MNzRVXerNqF2wPXvKn5STpiCK9RDwNjqKCz7u2lS8cfSPS59ydzjZb4E1y1j/z
fjpzDZ0qDvl86OkvG0ulIVNj/UIZb3ptFHWAuG/FADAr5T2uiXbOTqp/KK69Bb6N
/XRP0wchTMyLm+i0vzYE0a+dC778udnUaPpQMWYG/2Osi9sk6oyQuz4W0qRC3xte
NLr2ey/FSWkdZAVk4dsvmn6tcEZ7Ps4Nu1/Zrhrb0XQ3Pq66ETG0rrxly/Nd1xY4
LZQoXS/IVlMU49HOO+2nrag083MV4J6RvzqHLx3MH2SdzJ9z+djUOcINxhF2nzqt
9HcILTIEG8PrHaIkVOI/jz0ZM8hGWFjR5LcZ6Liny2qPU4cINdiwHLvxz46WT6PJ
dzVqLPiOJyg28Gd3DwB67aorgwbZwlS5fHE2s80kteZdUVG1X44JhV1oZQZJvLnj
comkGciGIzFfzcsa0+fYjuXSp5ok0rrfPH5xh4DmRq8CCXTRywtw/kYEfTvaFn9+
CUm0zSuiHp/In1GqBKeKLhLsQoihY/0YC4kqep5YYOL7C/Pg5DuMpXjBsqlnkODY
KPs5zz23MH5y9CnHYMOAc4pOPue6+WA6aB85OcB5jTa/4inXz3FZcw/wS/bWj9Gt
ejsNHgi/4UcY0ZSsj7Z+VX81/WBItVQ0If/1OnENm5iIuawfhdh4ZFdae2Hkyr7t
00a5B2ij4GRlcotjWrWHxNuG0y8B99KUj5uWg4lSja20PWmrT3ElDfzrPjmd9Z1A
2ydQ3eO59NB5nBNUbStn82GPLRXMJwhmzaswYnRxft+yy3IvX3JJchqIWgj5XZaN
lo2jnq7Fab8+Vs2z2Cij6YDhwOEOSOQP6qpj7MFIe8j1TCeum/ani9NEnZzWyXnO
E/csU4P6mTQvZD6wb7hvRFHsOWenhxdQjRfRkEmtjAcX1c+TBhmvWJSGuHnrx0QW
lBnVtWAiNPlsKrInEyJZaIQUwXFU2YgwtBuQFoPaOlPz+I0rhdab3rImgwJQDdOI
zDDq3YxId6P1V8XP///Of0R6m6leo8+McX/jKzzsVqBY7uIfzlWihqbzFgGqX9w7
LzLZ5FSAtEMXnsOPOJdEIMJJOliUJOaCz04ErRYcl3ov50cfR8RYuJWEfWIdEZcb
Nwd51SJbKbKVe2xiAajcHdjsslvH4pgYuyvM5zwb9NnocJywlYpOkPnNFEbu9l3L
Ys8IfHS5JmlgrWDw07Tms78IdEvUq8vib5/ywBiHz67OTpNQ5NOkxGc16YYvbWO9
TpX5AD2hzcbjeWCQ129XvzW1JcCIGu9QWs8/5bRCtFreqAkK69f9AqzUIcyHaCWp
ELFPM8eYFWJKxhsrDSVCqhEvxG0OSfwcDeNJMAYC3T016OrP4SYTTWlxz4rU3Vst
n5nt7uuh3YLHrCAIV5Y7GB9EHM3kP/pj9Z/e6r5vnvYNQT/c7UpMmvO6LNsg6sSl
6GrGlm9PhEpIYjM1WYPogkkFO2A9ET8VK1UjPfa6zu3c84hcvknHD1CbMu3pwuv8
s2YvGgG1/D/L6iwPk3NQ2gJ0B1059DR5Tr1S4im317bL1cQ4QwESc/uT6s9WXZHO
tny9AA5pXLD/gJwFeVBEQZ5ZB3IJtd+GbOqW/900XwHA94HLf4xmyOI9Nm5oZHoE
FnqqabKYnjXA5+yrrCMCmed6WXZmUhSjhuNm7lNxa9pO94ysrSI/U1GR+p90y7YT
66+cyFeUHINRkZZswDpiM8Ivu9h8ZW4dbeLwR14DQ+d+b2gVI+mt1Bs5/bfy8PCL
AOAFXU0sOec8BWj2hVs+0b1fDzNf1QL7A9AqgagPPzFVSBS3D9IAaRZ4o7pN+SXz
pNxh8L4R0C0LeNWz0CwJOhabmGnx/DPrKm8eKKQcHWIYtIYa8z/pAFWnlvA+UNmD
6lLHFimUm7KL1GROa8euue4b84G7S3Vqjj07WBjfztg1mXbivjfzy0G7ohnWcLCC
IgtaT6g+6Fgi1yw8eeoUuFmDpHThOKyo4gyn6DQHhYR4lEanYCULWDHVFbZGc147
gqhDuq5KKHuvNuLagdbuLpozaDEbB1ounjyAYNDohl/sh0lpjcPQV4/M24/nVXUD
MZE/A+nXVAAIhW6nubkHqVn4tufiMk6ti9SJmzwh7eRqcR53VhzYNjJT7BZcWPpE
Bhj5Kn1J3XZfE1XImYmfwpUOrc86gihB/RTKutwsmQVdz3HMxO1HBOd3vP5o+OeH
jsdjr/B25UEKlWqAlTRaJTVoetC57mD/NHEui0fP/qMoLi3NRR4OK/jwKwKLiwzT
VObrc/byDbtJXYSralAQVv3rqqgCat8A6NPhZxx0NaLzcJVLNZysJ8a2avif81k8
d6b4GvN1XrTdixm4fuUwUwoa76qRNVRKGVLDU2Nx9dXPgm2HQeXecU/De8HMxFRu
gAZQV8lzF+H0juV18KkJButUHtr5cuj3kpXOL6T3/jhZga1fFGMd0JFca6DUIEsC
YMXDvgKn8ZTHG2/8BOkN7TeghyCktDX/wpEctI7nmb35ha8pNROwFdm2cUpqnruf
xxjVf5AQ8v4ZT8eugFYxw5Z93rI3Jg708KchRREbDv9uKs4nn2AzoTDCnoL00mNl
gJVBAzRR/9KeuCrS4QkplW35NbovoNNm/TJzWHE/mhL4T77OZDsYu9rQ5+mrnCTD
lz5BGT/EN2f5YVDFI3NsAmbj5ZrTXBIg3hg85GH0/rLpvG0SzWugdkFrUFkGvhtB
4B+RA666QymN4Onqym4S5JSqHTzjChgBPeedTxnXKpSGyEdmQOdCWGsrs6Ly1JmB
H6dVbTl0r9CUN247z0jRMvFYi1SAv89scdoobHr8TDThx811z8MKVDXl0BC5wm/P
FxSNhiUK4zygPwzo9RI/qSa0LUT4Y7gyQ+d642d8grD/Oo5QhncxTizXSrvyi7Cp
KpeKyYAQVEO7QgL2Xvy4Vq93SfptdFxSxjUxHjyCNWoj5Wb2NniZwRZo8ox8G9sw
SuHUKK/Eiq9z8RFO6idQydqD/+U8E0f5rW78I7S9rD3BjmRglKEBYlMKSVXWnnGw
Jw+Dqs0CIxlvQQ4jtfwheKIHgeVNNc145exnTK3PcxnksRhnsxfwF2zB1ib7oRd0
EKI6s4SNhRGNP3S7oiTDVEI1zdf2VF/tfrmdboC5+3lIJ/6+pifOROO+P+TKNi25
lsK929XXUTySxgQonurpaWdABV3z/Ttg0duxDiyc4B11PpssptX7nHmc1TEc4MYH
cHFiT4QPnEBFlPnD+4vRJfsUXMEdgw/j2akm8xpU6+4vL0vkPwLHQNzFkKqkU/iF
OqS0P69stvPhrtynx2Z8DC3z+YMK/1tFB2VUT+zlCISOyKynnbAW5uNWQN5iM0g8
BdbWnlxfTJqTzNgjKBRcKNnIHfzta1aSMJg39PhPMuaGwzwzqo8a0wTvBqeLwDo7
KgVmdKZJ/r1OZqA2/5XzZrhFccAfQuMZLg7vhwVt8oFJz2ZlNqnf6O7zMlxlcA/2
nk9Xuv8LXuJmu2cItRJXwt68Wl/i5cGY+yR/oMlvzHLdInxAAAFlpuLeffu1ZLGa
LnuRZlckqffbwlOavG8haabhVaDBiQOfXCWhqmlxXjeHTJJ6zPMAEVLKOjhSlMvr
h3rHgKdhWV4asMfNW1j/2xclOIT4tkZNi2grAV+vdsErtMN1t0B8o2GHjZxSbwMN
t23K/jDziuDLJD9tcVs7eKK2hJSZr/ksM+fu6LaB74/SM7+6Nks9SbPJ6hpFbOzn
CSUBGEQP+MIzVKYLVeSoTRq4Z7saLN/0ZPtQxlxa+DSLywqBWiwhV6o/yCAMHH70
so+ekPEbSlX8lvQmdUIc267ET2WHRmQC6x9JAy8kUymGNA5v3wgBgMqXpN4ro9Uh
wKJrueOdS25Nw0dWzL5SGKfvu8vdPgVHZJ6WZZHjSgjdgy0JpizqMFsz6slwTz7I
UiWkd3SEBXCluTMp3261g81kamwbnPC0tnlRn5V2pI7Gzg2qjxLGR2dysCZ0+5sv
YXiUw7Gxl6OeqQxuqBMSBecBsIkDeP2tvbtok77CqIgbRgDcFbssD247RVDk/zom
sqmjvWxlhnPBeQwazvGzNJNepUh4yyoy0pE2I1UfHWeVR4+jlQ899HASLxA0NeiZ
kVwDRl1+i1XTFe8r1J2zsXzVAV/kRRhMmviempqYU7HR5Fr6m8tvhh4re9kVUMjA
uo2wviLzjBZaEtJM5nnzeBaOlGSnSySbTVCR3wJ50F0GvWCEzRu2tsgigzBe5oFW
JD/NAcAxkSIcW/Cnto0BwNbSxxbYlbrn14yRTBnMuUij2pw53RHZwyHgI3YcbGP1
mrqqokBIiePq7DjlZBDWIoa8xMu7c4tJbAwcqQz22KBIPHfLw2t4rju5cz1sEn2l
hOVryUv3Z7fIRgnSKIF2J68h2aoRBVJZrJDmoNv4SgtHa4N85lHB+RayBiqmBXj1
NH5H9bUVcvYpzUiWoTGYFW6nyfdhJbYCkDGsbzNGaQuQfLs9tDindm+2MoEnvcDZ
/4mdvI2nGtc5uauzsiEY8AiCamp1PWzu8e7F3g0aJsi1XU1kUALf9w24NQKsubyE
zkyhO3JfwT1K0hFMzSlNSKq69+NB1L6sQ2gJPayqL3HGe7DLoEhf9EJFuiD+TqyK
sFKCTi0AP4d6IMgcn7YoYPOnhj9w233f31TflitXAc2Yr7oZU2W8uPrsY+N8dba+
ubH1P6S4U0vDtM7B7FFdjHh/tqaeW0rOO7nU4V9GxAK4fXnAD1DaNDMQyy46NgOc
ZAHhqYygPfJmF0aA1simeUyVvank0Hugkli1Z3wxpSz6W8mgBqeObVbWKY6gpaHT
/AhxvKxHdehyVxMaki54H0ndr5nIHiQrR1RL42tbioNC3wIjwPF6OlTT1oE+V5RW
uUvE286jXLhJBh14KYFAJxPqPBYNvgzfO7+xFya//zBnurl03e/CDKpvz8Elq1G+
Q7qr5O2btt3j49eLTDIAfSdraFQ1bjPr6qH4ZY7ja6MSfwKQzEDFtKyyCsTL5Guk
7pRiqH885irbKRZgVN2H77pl7mVmZEKZ3TAjQY6YRXJiT59Zx1DpOh9BYn4GEbER
pVC1JDgybCH6S+TuuYz7RaQ+aFvNhj08fQXp+s3sGoctiDsM+1/o02FSnvlL4HYb
HIZBXdZIjD8oO/QsOzkawK6avZEWPdLrHxf4JCX3VSWTXVWNXPFkIQaIMprfhQpy
6kDHifUpaMPJgDf5vN9B1p1nv0X9AF0dJE7elCRA5ai4L1hu3wK/RnOu6uvPYUfZ
IVE5pOymuxB60S2WI1wPL2LvCXutdkQWp3/wotHBo6uECMAaojUVtU2N1u5SETKH
O7vid5bV+tKxYd4FSG7GG0tHW7l2KOnBWe9ugznqXItLjVWbmCpfo9EU0UIk8IH6
0d/P8fLG5RSHy7QTI6F2mMRbUTkurAC+CCiwpNkrKbNjcEophMLkaKn9pJGse4HH
VDXko5Hkq2tPRpyp7HVGIDSG2x6QUc8oAQdW+TBqoW3M8bbDP1Yr9OMWejxgoq2R
i2bCx6e3KfD2BDqab6/vFWYiaseWclRkAV1+lPQl4O1Uv0URZHPQDH2LRyprnt0X
bcetMt+wsfYIR74v+8wjD2rns3DrziWRZPBJdtfW73p0WJE7RnHLyfqJs5CRdWHv
KbAjBnXLVZyCPhu4Z+0BGF4eH2Sjd8hma6k/p9wR4Cy3Cbtcymd+lpuyGycU+uJA
iQm9+0xePzWp6DG/Wz0yArEMOnWfqTIBm7dseQ0j6hQCVY4wnPQ5Bz7uKHVMr4iA
H1Q8VjhmyWLqg3IafM4eWl79ZEXtk9kNzw2f3W3zZmIcJHiwYxgzqrnfsknEUj8v
EdCXzZLrwvFUxjEGowVoZIdopdikmjDImBZOYpvwi4qZObDO1eD4eXY01uz+y8ge
a1GeH77TAH5BO5QSHqW1y6lXMfVK1qzXlKs0ixTBlTEG/95URUNaktPwR1n8ZzmQ
t2jj4QBaeRbiH6UBeDKJ+BxnoDTbgXM9WHXFNP72b8bVa6N5n+fK0sl/8A/UgXnz
lRvo4zUGAnYu10MpJ3zhWRa/a5qALAmQzUVjZ+60mQi1/3F/Z17ur0pMCUhOemVu
inP4QHkQQ2ntrXBx7Zi9M6U7bvu1tUjtPyIufWjQSAT5Sy3dePdZPsl1AMFFCtFr
Q09tFr40e+GydlaVrI9phrmzejvh5uF0MHtLi8qkUarruMwOSpYUu9lZ3TPLWe+A
FwVwukDHQ1hgbyQMOVKKk+TcpHKxS9a916B1gYvCNVv9JURDm22DEzOmPWE6X9Wo
6LlhRU7yQ7dYH+XlKk0aHitPB/zB0ndRrylUj5Vko7OReEOy4mPqLWgE847rTDmq
Zwz4d6Po24WI/mlwNbVqNfaRulCvuIgizpTK2uaaZTmHgiReaJHdo9XpF8EU1svC
/DxxD7RKU4G1WHSXMvoI9+rpgIN/ZJNyQ548ilYmMcFK50jiFXJ+zPfuQXmaw9NM
GzNjxA+UElrVBNZlGrRju4wjdIDkPgGM/TaP2OQCjgtEs/paiWDNrqWtr1SmSQwu
9bmqaDSkttMI6nwuJWZXrvb4x/C14OEIJw2qXm8yajihnrCR7rBFuC2D64s6cevO
BWEVxjTZm1FE98ptX9y/chkttfqT4fGAfUTyKMVgb9edp23A/pHPI4EwvN5ve8y+
h/ZrhCA5aOaW3aF+G+Snaxb4l9m4WCbQd9NlH7tHmD8YoBoUgBdu16Y31C7TzXvD
Ni2opwNwSJ/FgR8WfTWtH2FxX2hVFP9eAW41uS1mxZQN3rPO61B70tWaeGL3zrza
ETTMzzKx2tzDVNQDT7u6CjXvuCl9QCyHvwII5NtXGqse6F0/Ti3haNBi59ruRRZ3
NqifzHd0pDGHngqQYwoQY944X5aYZt+GjOzT7t5yAoiBUxn5bWxK4+4vGm1VF1ab
ISgQ2+dH2NlNSaBTsrXR390dQp97P+VxewCfgGVWE0iFJfU0K0OVcf7nZ2zNmj/F
Q9w2/bklt8t8Ol1zCBdmT1NH/jfoTnHzNvKmR4n7yPojseu0lfVq9F4eElnOW/qO
Jp59SiBvzrqIA/3A+ERHVgIGXVfhONrMsg846UKV1Xji03SiSorXMn8HwtMvqWqw
dvCmcYNT5rFNuDdhnoYuJ1+KZHT/ZgB67JzPyR98n0BHW/PhmXw2aCuQrorskdAq
MBmypVoF1+Ex4KJGKEeS8fnmshLdZx74Ja1Vmq0QsBsNEetRCWLXP5I0GlUij8zq
d52ulWWf0etPOwrQqjda2V7/vVWPzEKQFYPlBZUI7YE8eJlAL01DUKUI4itTXxc+
fWcg+QGGwrMyzaScxOoHo+bIicMusfn3Ai9TZFMFUoIit/8ReJgOjIM1UY4puWF7
IfsxeAMtO4rqYaziVBIpBrqjEyRwZdQQdxRg5AgmN3p/B8tM/5aGDER7q2/PUnhr
BDrt59umQQ/poHrsRSWFvoCNaY+ZBml9u0ynuDPOHl8V4V/5PQYMVK3yLTMzAylU
EB5oCTLgMi6lx8q4knqdf4rjhDYrJ2txV6v303tvacZfxyGtxBTRMPovWVJUowAT
UHuTmTaUxoI1Ihl25lrspZ3Jrig9u1xp8bqL4vYRQUuQsH7BfmRZtNu+bv4kC5KE
sXezZ7fv2C67ASRLj0fbwzSzKFDGz+c+P/uZLsfrsQYy4rORdXU1bGA7GjzSabiZ
cWlCqGA5VFbIUeeMU3+9N0rT8pkas0ytcAw6AawIOhR6DYSnJZqPTijnPTQVfQ1b
FUXC2O+JLsqvWXEwsI/PXNVxlAu6lVzYRMMvWl/EXchU7m8wtsxheHg5JX/+xvuK
Zr3jXZ3hcPuy1mVp4Xf3QlKaWDIbxDNMjO3Lrs9XPVxe7UQWAZusNv9cd10l2WVw
86XXNDtbb0vSdHz5XiDXoQW1KFntj3FKQOR1BRHYNcQskSh1/TfE37iDuRZak88z
4sP5h82EbnXWNruZznjjZdRU3C+hCJP40Z/tAQ/NCDiXXZJvTiPFNYLLM1YoNQci
OYZH+tfKpU08BzzPB+6eqkIinsyuN4B1hjXqRf45Zs8r69uNztGQPwP+qOg+T7SB
`protect END_PROTECTED
