`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N5SGi07ABkdXX6VgfLav2bU3/VH38bUp/e79BIu8Pa/5xuIohACzAv/Cvm2oBx/Z
xjc5jUmhRicffpmPlgXp5y3sKMq27OhsD0Dvc7efo6IcV85C30NyWt8jrp9y/9TP
zxBcVPV5VlQGL9Y63LrFgMBjC486Uplm/DZUF8KcdueW17Udid3SE6lT5ssNUAGw
NCFd5LRw4/XbOIMTO7j3V8olIkkb5rft4gVsTO5Mt6W+u0+UCx02izrHeSFTLByr
xnS/7Z87q8PypdgFmI0srhVv059yOgUamgAZtZ4Nc4SRzw8Gneqt6c9KiEAUYKAX
jngDqoGEIGFvtU5qzuHBhM+fNvsxiMEYt/qAAriy2gNNAPNB2aXJD97OlnVBhoAm
+6u8fN/gXATVVbbSqMnl0uDRqPz36oxKYVIw8nD5jbTRtQUKwgmRIivt7rMRVjT2
Puhq/Q8I1Aiw7ZdLJUxotj7XWi+Chql7KJ+DpavOTkE+xP1Mc6960ZOaTEfSmR0s
M2ds6qBVSvx+PAtdHN2dAkks+ohUOedzKLMF7wxAdhTyxDKExdPhf3vAkYvznFrH
Kv/cdngjasVgbwCRQyDxYv45jXzxq7jFbOQ+TrM4/FEjsufjTDrraMC/qbqksQDW
7Frp/iTzdPI3nCTy0qj6zW6BM0XT2KbHyFHgyMKEnk58VwHioPtfbyl54Ks6jjJl
iZWGvqnVE47x8zG9A3SyaDuawigtplgzI/bWeL+xT7Sp2eJ4YeKbHLh4t56CMooE
o31tirTQMoWFDvEHvvOup1QA2V1Zw4pJL9k0RJCmP5oLLqgDrM+v55wKqcIJLjnj
3RFW0SxQXWw5eh4xCIl1JfVZcXwXMHhfM1WHn3iWkC6WyvAWJu1e5VPfRxbwZLMP
s4K7xruLs1gj81b9zd1aIDOQ149NmcPZKwFLquPdKnIziuGulDzDfa6ScT906glI
2eazRwXvFcNb84mgjRR9/E/wz/ZCsQA0Zt4Z8Jt6RCH0x0npDUz9cqkfIk5A7tt6
E8ziiUtnOA7o9adnaFwZnsPKkoMF3YUeoyJew2hfS16yzdrF9FoXQjaTkBGzx+DF
dc01VcxuzzMI190Lj2SoaDf28BYUVgNvxiQeiLYt9JPFpTM7UtaV2pgbmUs2S3+F
StQQVM1I2vdgkqBa//hC34SfrlUkJtThimO4Gj6BwWdK5mpqn/n5NZKr7QtV9lxf
XkmMMitJSKZiodYLtsmkhYYs82pLXl/XltAgAk3UNJqELl0EFhwxrwGGo45IYd/y
mXSPPH7Uys0LUyoU7yjZdb/VQMNnWNMJDZ7OwnK/2UP/U/QU6cL0un5vLzPu52mM
a7UKA4PkCanzHHlsQDSHYZgmi9R5n9YvhlSAYZhExVN+ypmGpzqb/9RYeGu7SpAl
ulJWIehSU4bzC5418PIFX9HGyAUI7ubutiw3AgZ3LQaOsVgqs43bzUmEzqEUuAVd
iKu2bOL2OdbwweSEanpxc+mYhkSY0xw7eiVLIXxe7Hrc8du6nh1QJCYjHVq6pcCm
IS8lqbhcjRSoxByOSU2W5Ol0hG1mn8MfvVQCURvdeXC1nVICp9amzvYFrr/nYZ9n
lp2pHRUMYcwkwi7rP1J+BFuL9nWmRSsHnTq1CQL6dHvjsesj2YLOuQMFf8YCPn8y
ocwfgOfRHA2ACENsb9Djg8Ce+5PkTBI5SOFPmOmkDpvkS7x7xGKjpZEaBpa84IgE
paW5thm9k3BRf3l2IdYHKqncTPMLMKQ2jgPYfA1w3UhP+W0Wxt2l8x1NOvDNxOp2
hHQEMk2ARPZaeKhUu54veaRVK2PEsqTSp26Q3++Z52tmzDTs4t0cFlQ6W+3ac3hw
ROUmsXl89LhIHfncs4sBI0bbKq1wfCVXqO5J4Z1J2NVDTpFaG9kNBsvD6FhA3Ns6
10UhjwzPImCRFbBBfRWVgn51Q4pt1mnA24LDjClVMOg48j3VHLe7TDatc2I1mXUZ
6eX8Np78M6Ti+gxXDXIw0AblAJhaN/FOCAmy91QEpgEZh/3ZbHXy6VMfDKLv3JvE
7PPjvONXJ91m3QyDzG4097zwo4Em1W3+Ml+KcES8DSxzx1FurmR3Gd5z3Te7W5MU
b080j+Egnw1xpTH8wAeRj0t3/Ej0q98SVe9DEwq3pLUXTffxbc4tyQvvQVxBg7ao
JjMSud3L0AJH9Pd+r68ONDiFt6nVGjvYhWlIhe46nZsafqCVORQ6OLGe1+CZ93HN
6xk2R3woRIr8PljjumW46WQaJO0//QzAUbl7hzqo3Z2S6Bge5qx9TZzbMQgUvzGE
qYdyFmxy59lyTGzkBcEWZtCyUKhRWHys0eYxaMvhCKN8ybWNDLO+/mU6r38w+Fuz
YiidP4iKtLUaGw/YuxBFyaFWzx3JfJAGkcHT71KQp7FIDpvyMHO/xvF13+djfaNm
Gi2F/Hw5EQVc87K7PWDhXCmtvH0wUYGLCMxf2wAz0p9ROzyhWwPatcCCgGfuE90z
QiW1rnnZWQepXtS1ET+MvvyipDxeBS1i0BifNEDPegzWdku3pWQF0R/xfoXRlHAY
cDaI1WqNOvV58+6mUutW9FpC/Id7sjPwVctW8xI7YGiFESb4j6tZ8U+VI92f9tDt
sDO0drTkPyamkdBW32bVexAQDxCDjy1/fzyzUFQPG6nemlD+r8yCh6ufQ019sOZH
Q/GKoR2dD7vTxgBtyYL5dYBu4aQsUwptiGYdCXJIFef5cML0lwljpIztOQjmiBjC
lsrO9J0OcAmt+awRNPY8pv9nw1GOiBh2P6KUCr6sTCalI1ENX5ATForY6J+mK8bN
uR2KCwPzRn237mU5+t8JkowqrV3OnxcE5j3vw7/As+Ga6GCtB8A0ZQZhvJqZ/hTa
tEDik/Fj6BBTDsoegGAm61kMuVC+i5SYdtiA0X/Sa6Fg4tsyvHMCF2THmaBefjTg
FYzMAjYwHs8ANusmn28FPg3FxDsHgfZPCMWGTrBBY6HqwBsacySVQVwwRfraby64
y3YrEdULbtUW5+IMTtdemvucxXM25CTqgwVrFgyMZcuw5lqTsVvjU03azJIi3aAd
HoMKuofZtcz5ZCQ/KsU6nQBNun//S7gApZmO9k7xJZGrgLemN7EOmc5s1jc3DOFW
TVcCdVexbnhtuTld/Wzz4IGoFPOWPhLOcN5xu7qpLgRnaIFeD66Kp46l8LrJ/2sU
ywZAoh32SPFhTcaacmGXvcUIr6IBnDj/YT4Y8Y9iaDwU14/P1nIp1kONYHqS0hPd
eaq9MoaU8+suyHNu2ecrEbPMEC5zEPHOU++SIZJ8nI+qxiHKuOS29HNyTDK4Od9Y
dYAZSmp83KMUItQ85tj791kvTiCufPS0ZgLGQ6q1D5TD4iV0uxKZyVjYfbqdxVtv
toQy40i1hV1EJ2Rnbqt7M8xx3FC/PxcHw+lMbVBUEglRZywwPVLAInuLAD+ZlA8e
/eahAD2EPoGENDQ5v1f9KhNzx+JMYZAyZ+JSO+E6ls8MRrLKrSkk8DbaEO4aPfBN
qxVoc66aHO0nG6QnqXhH4t4KGNmo0Hg2zM93MWUarGBxYbzxeMUqQm5dh+qpUDV6
sgP4YhG6t+clruISfeLPY9IO9Y+Sk3ODUr01YJH+Iir5jBOPtwcSfAF6V1oPX48q
fU6hhZTjNxB4GVOlRhQ6Vk8zgWvhgCpvSat94XQyu6Z5+NEuwkQ4ue6RYbpqoAyy
kR0M4qpH6C4nvODn+m70j8KXidv6pJ5zr+zLieguk00p/wq8fsHlDXI+qAYbS1iN
gHMZz/fsKXlBSjm0WZ8xTgu70qeCr/lFojLLwTL7hWtVENs6O/t8U2sqhjml4ZQF
YuPXkYGD4bLpDwAciLC9m+KZIT8O4HD9Soo70CMwfNQFE9YRxbw7PHNWPcoY/t2d
EaTEYgo1JUFvxTNrvX718uP1ra9sDwKvXdxR3A2TyYaAQJr1se6VmdvOHQ5bhZRk
pm6yuUXr+AFJM5bJKvHkKRex/N/chzseHMBvRVnLi54Btf/c9RGGVirtK99AOZKC
l+010ByL4DArKxf8v+cpgwjJUaNXHOXC9WCQdts5YsQ5xBzBPnH8pZD79QL9N04j
4NmFiBIuuvsKnKxV3ODDgfIQz4QtYV+ttbTn1saetqPGL1rnAzOl8pUSsTAR+7Ks
e2tudIN5b7FhKXAFTHs75duRdZq1rrAPkH8BAZLP+g/4WH6eRitzfSIeWWa288CF
IhFZ9qV9G1BTY4C3/Cbg8PAmbVoh7zlAtRRqZFUuvU4If5P2ep2akwcihYzj46dn
iqD+3W0egf+2sJAH48F2+KWcH+dzThdJjzFVr9867SB2hud34bqzkvlshPlJeLnx
iPWrVzUpbVLk84Vv8SAWnVwkLrxu+kijUPVK9ztJVcSQmTVjc1+s4E3mDy7EMn83
n0SSchbFFFGKt7tXlKEwvygH9bD66MsmWwdbhNPsF5EfGSQQJbSedduDmiOtVSix
/JiWUoeTpAD1snVbfvkjLXNXbRJ89ITh9/ObAij6DRzRq7GkZhfbOY4m1ce6xy/X
LfgcdHJQBbQ8cpmf4GjyV/PXJObO7wgJb7Cq0OXUVEeCAQeLZcuE9CHc9/cQqnQK
N9YSvEk/lHsKHWUi8JqMDjUc4ycRtNSmru6SmfXZDFPGdKZ9C9B3c3L9KiQ5kDml
zvlvdWIQlwZZWl8ZuOG+QHtzQe8ax0ZMyUwwip/89jP1HPj5k8U4mdOK1Zv/A0YW
kTUrXgP0IpaeQO/b3SDAaLPPwC6/kcAVbMiXXgnNLGTf3SxAXZWIP62Dn1tx6Xkz
MkC6Oyp3/xKGCQqJsjqKTRLUNbF/eq9ePzQqlutuYUSehPNptry66hbo1EiX78hy
AMHWujjyUt4pZvVP7CMZt1ozxwK29JXkV3wIPdXLGig0csclxXcP2NEmSAf3X2AP
yU1rrfClmd1RvE+LvC2LDKNN3R4zrC9vAyv4Qy4HqtZPkMeWea0SaJKO4gDZqzuH
LDaLE7wPiAcaFam1S5lB7SVziQOfzxpk7KvJNLMnF1ybisfCHS0vORGBl7ulZThP
W5HpGtbdTVrGG/qQNleZUGXFP3Y2H5Bn2ZizTjGkXU8PkTfjn0OkJMikTBAvz2ZL
EPiavJInqUFoTBfLqKmTGdA8k6NU9Q6Z9JrlnrrETN/VYTtc8BUGjNzbDeN/tk6/
CpBb6h2mz1YwCVsQmCMGqWJjwRLPLXjKebxszU6adMlNkLf2wr37mZh45GSefCap
/LxYwFtwFr+ubD0EgAXyfT9MOTHoNg29eDJq8qoSS6miKiFnG0idwDU+/uiaAx4M
QpsqwCIss+i74pIzeCykgP3pcN1SqvlNl7B7IvxshkL2Ax3NdTr3U9kira7Zu7wM
lqB5/5Li/iA5Q2S4mz5qDPd146uVQaWJYMGH1aRN+6CbYZ8a38V44856xl0mBj23
jUtIK11Ao3lzzJDLJbyZLHvoE5NWLYAgba+cRdWMEuB6A3zPrShWX3HIw0D8LZyx
DDJJZG1PGp2UC9pK6e6qsf+BrN21WP9U22nzHOJLTTzfEtHRkVggteuKfNjtuGnM
fvGaHRU/EcmfAODcLy7f+kCxPk6QrkcBTgSe8UpaoQQP6jWgEdOmvei4jz42+Ave
8Qvv5QT/47F3B6CpXbWXfgSAIYu7wVYLQcxv/GmrIZJy/GcIo/xH5kv2fXmr6a+6
nbH6W5gVv1oMVAY942F3kKd0Tb9f8XmHGV/qJq9kKFOg037EB7WL/PzTD4iD/DBp
t4S701D57BSrKce3KmexF4zqqiW8MdGoWDhjXnHaxnpfPSeHghRU04ZqKnPFDULz
jMDdzeI+P/Lln1hwEhGn9+uax3DhsALBmjDL6yWt8wop1d0qF2x0a0Rg/JtGAu2o
PNDJREW7wuWbcCb6EBBhkkh+B0KIzx9GLMku68tHQZ4P8J1Z6lA+613s/mv4FluV
eKiQentqK8HvjAmJo1NNPr8n6WVeLua/PkKizjwO/J3xTVOyMQmdihKkyKpSBLn+
/LsZ2+5WjCjqGS+BmusB9WY2edjrRKog61ycjzEFEQZq2k/EDJ50cgzDvW46LhKR
pd04yzdoadCPLgQEYe0QZnMZiWBEc56gGaiPVS0fy2skVs2cf21TqFuX8U1BQ2J7
EYSP3kcvBLPS2l+ELYRuoP7vNTrOxb28vfMqdql8AyHqOXa1BOxclnexU7Le4vzu
9CzpwscYUUuhYfhYDMQ9eqA8fGrXrWqXQyS5ct4wIHHR9p0F0LNO858dJIh3W7cN
ggxUYAuaPDTmp6z9gsaM5dMRU7lnMY2UJZFHqyVhlk35YX8NPvEn2kq+8yGvF1DB
SOyQseSjQ6RYA7oIc7lJkpvG5Iiqp4xXqw5LvzVe1kBPOHLm6HguK1zbd4j3qeGa
iMcDv8xQdzKcSckFuU/ergNP5D7ATwtxhY8tsCeDETI3k4czTnRmIIxFvLwz+V2T
JJOYzJnYDYG2b2YsPnW53rc6O54VYk9VpH+UuTQhPnoIMXn+e7FD8EoIylCYzahY
1nG4Hcq0Z3N6geBAXkJ+RLOtKkeE4qJs99Iu+TvkNfAd1SQpkAb9lAsIlr94uV0+
qzqjSQAW+GeFeu9fdvrMAYezDSoWpVpl6skNj18+479CKEuqD2cqKsEDF/Y8aB5O
yrUYLL3pCCmSGHL1UN+ij74vOp6lF8HYWg9zboWZLPpieEEmJBVRuXafPWlu3/16
0ZBEhBbQu+eUOQwzzPIDJh+ffX4t+q8Sx+iX8dpv+cLUYBGpFIeSuKW6GLroM92Z
ROMMEMAnpLUpUTQY5zVYlRFUD6fsKdbOfIEU3zP+siX+xy/GMSssuJGZphyU/dIc
GHQKWmjpvvtEpiw5dPpmM16vr8qpNl4+54R5/2BuC2Mjl5Wu2bMLn3mYgQKujR+j
mRPamR+Xeu3owvmGlbZhG/k0uxm80Kivn6Qm9H/P6CBfIZs68EO29bE6YgTjmdyJ
TnoA7rAL/EPXprQ7hpJ5SRs9jH1S8XPbnq3rAHIIeZkPLMXzzIfZl14cij+YXJi7
Gk9guI/vpxdnkdEOv+KuuV1SIbhNIZ5y9h9DgCkQ1e2yCv4LX8edaCx9snsldUPY
jVlqatM42Kg8vOKX3p/OxSRc0AETcwJzSOP2iP9NCyoCVAgnJzWnv+Alekc9Kju2
k71+cx2B85kzcbZC7Do9ug3azRDyRauOLpBGKqy15GBwFDxerYIV53jEkIVMLtWj
APr0UvRwpxmbtEHiZqBz2ZlNDryY/DwbfzFPYd8fBy/aOXVyhfLQGGMxicCvxHXW
dxxuXFXFmYAGXBb9Gmgd230K3LOHW3oVDeHxq1n7mxThYOn58y3YpJ7vdbPDSPNy
TTqc686SOx3c4SXRpoXGUUKJxAKaqO1eXS6/BceMJ4ZlAOo5RvSRcYiihle2gfNx
HlJN6Lwfl0G5GScLfi2eC0dbGQIpCpyWKsEw2ming3vKsXaczzT8lGdz+t8PS8BL
FVnk1hXb478SDauVuy7N2HiRPCleSkhOM0DDXH0mbEI9OP/Jz6zWGS0j/DueMURZ
7oxv3DK2tonxZQMa6q6S/pvKOYw14m+OZj4NtV3NwwVQHr3FLcXQwpAkA6ohlirU
RHg6OjGWCv2OkFjglnBzPysaLGHizS09n0me5dPyG+exZRloGEEo/H3WT+97TAmV
TAkgZSGh8fAd/xMhajosUqP/HsO+e36lURTGSfEmyniaA6AnUJFiZc46jmZFpxt8
bYHwcTrS4C75+vWPOs1jyCJnsJej8f7t3Dz0OS+c5S8n3CNBONeiRNngD8+De9Ta
+cQC6OXe91RzICkUxnxlvKgGShaOwL0fUsQAYWy3M+oExO2Zus0SPvV1coMW9FYk
xXx/62tNkG5woMKp7pc2h1DhZI0XVZbJHLG4QJ/6VBE6yICUpu7galVcya1NOb0/
i2n1TIzg7YSfwQBi5zSs0vtyYUKGj3QNlUBfphh7GLKEruervD5+Sbl2rKYQMDGE
edcBGeoF3VRVXKSdaE+DLNY1MXrUz8IMV6uUnAXsM7dOHgPZUTU0ouJ1gwlFxBAK
XPObV8twJAziWTqGBBqnevKcI5WZfDNeGd27ndl893CUJDiNjeSBhhovp+l+FX1Y
ZbO/I+PfJz9Ax080sjE5QdP1S9KoUk8OkrOQS8FgBBMIDUjeSG2CfcrdyUBJMsUU
3DOAoglcBl9h0ms0fjwZIHbW/+BdCeZ7VPudYIqlnD4p6vq66bsF7PS2H9drgGNw
ToPGf0h8LQQksI7YWmlgnvN1Bvr82krPBFKeDP0wmaGOvDdAD9G0p7l07OPZOUPV
sBm7WoCWUOYZnAZuRBey/EKjtgxb7C9JolGtLjCydshj/HW5OPYAUH6uBikU2OQf
UjGvL0hvRJQtL+ZFmalHawzfYJIfPKsHZnaIoI+lh2fzav7gVgfzBnhmVPhUAW+T
L+83c/7rGUKCiktN2djcTlmF9w2D6KIHJYXxvUnSxYBlZuxAbhcSqPsmsAvVzPEg
Co8NzwOX91QyTQ3eY5IXV27O3hRIMuxtuuYk5JGPKb8ZCJGXMbKrpK554KebHLfh
ohhbAJdddYnkTcL+pUL2BzYuz6hEcja/sKWCdxzogcUe72AYjiFbz1YjjWUwqVND
i7x3arfCgHJU0S4CnTioM/aG77Vgyz3AsrauE20N31N+tzBNXigHmCuEchOtgOS8
uJRigKsmtQHLZsS2zHnN8YwIQxGcEs020hFQwQrr2f92vMEpBEEb7Rj4cKh+iAbW
5bANgTTcL2zta9PZZTMbn8OFJ4XtCuFXnPxYN8IQwLp4zBeHlDZoKMxQrL+IQYFR
cNbN2oXrS4ZYOa/62c0zGt3ezRZ27aOEUMqOixI6Swz2519LpJoxoMlz6qSGKsL6
iQ3/aHlvH+5YoaK92EP6s23yG5dcYAodtf7v+ZT0gnEoxbscStfASY2gpqeOdyAq
oWIsQ88N6X+Qb2Cd/F7+YKmJG7uFRsw0xoMGKTcUUe250elepRt2nlIgIXrgQ3uK
QS9MOxR1gAH+8zN4ZzztUiU2c9YK6nBruBC2Iu2BUs+QtDqzMrD2U1ZzPuFTW5AL
zQffS5qa0yABuJRVWi7eW9JwpdO+EZ8787exr6mmfnNB4NKQQWGOohmDutzZx/NK
G6PXBdBU/FMsIaitKWvr4TdkGdJT0dwSmW404ovcTGBPgotcDraBvMCUX1S1Xt2q
nL11tjjlOs3ryM2ztswIe7t63Y1hyTBy3Ssjvw79oWuirk80Y0gd3rqVDOXH2vHe
InNIO2kfcbn2RQPs4HFQ+qPU/y4iQYeGLTAerdeldPV9eXZpnrloDB1AZTBTCFqS
X0v1sq4wQ7eL48AuWODD2XyTQuVQSL6FdWEcupyS8em4WRyBSpzDd757nqK/hGdJ
mBnipyZgvYKeZ4EHxdgM4WxY8ZuOsyabTRUu8Svzci4qJyohfIrCHp+d6+9nwSaa
7HipprnQVAK1Jcg6TIBn9xX2JWsUlRKETXvJexO1J3UGBacLvKBX3TCOVKGVzcsW
dqmK7EBWkUM1E1YNIr6SMOUGe7H87HTWtEo9ddee0wu9gx87KovzgvkN8AOMzSis
fmyJXeDo18lpQ+kYoWfgDlLxso5n+cdkiNsqQiwXeU+2piy8+OIX0GruGSMHdUs/
cIgo8yXvbB9dXCjr3fCNIIjWoAg3knff1oFMLpeLlgmegmhj4vbytRCbDbmflmF1
DmujFOmyLWCrJRt9E3VIoEVh6momEiYg1OpYjHldonTBeTDycDP7SVOkqKKF25TY
cH9VqO1ci+g1f2Bzo6fYWTJBzEAVPzTSfkO+BA2UCHwavrtJeeUaAQn4daEVTlbV
2J74hxtHqrkbdAmbG4vfEvJ7uA948ZSzlqQWNP6IZIidDp/0rUuk9Q2O2Ed5Qjy/
vxSG7C+efrCdTGjQLbjfuLPcnKjwrF56P/dWxGQSRTq9G9EAwDRb5DS+pIBztd73
XYiKsjTvit8DtnxTmWXNQ75RfGphsd5nDARaqd5EElauIyB9INs0yEx7QPY38cSw
ZuV/BVnTw0LXZV6rbYa0d12m0gLl2jJ1JXcjEP9dy3Wi8RnTE6N4uNiqV0GgG0lv
k2Vfgib7SkNy1GkwATqd6z+thikct52yXQg5xzqyDcZstuXdOStsW8wnYdQYnMUZ
qGZKhWHopTQR5BAo1yF2x8gquyXXBUyVM/oY0ifF+cGNE//KqZLl4DzKussB7pw9
5fJ62R6HMxYaB5unqMvkUIS9aTlST443XHfsnd519/lm6W2GhUUqspV6clQ7mZgl
oxoRaOGlZTuPSwof2/ACakpcw4/K61CwGP4r7hMkczgyS1J7cvb5MEbWZpEWrYet
M9liG+CddtOst0a2aRmH0p5CoMxkXuGpVA2SJG8Ux+dreus5f+be68Ga3zKJyEPk
wtlrPh0Scwk303u9qTlSnnj4lbIIPUY1fcRI/O9a0MFxNQwqkeoRaWFNtozIAGTe
DR5vlyhju+fif29iHEvm1J86qTaAFSma1LcgNkfrEtcHiRBhV94zkep0D3JFiDZG
RDfv4I8KnAhGbwCAEUXyd7NgktYW/Kc7R2NGJNaSMgDi6AzlEsNGESXXlr1DQMox
hOROpcMhQBvhEG02G2HbfzNfIA4/SpN4f7lCtolcN7Uh+XKzIVc2GMZphD2/mCw6
wIrKkuw8Y1s5PlD2LT7MsQ2p5O3g4IqfjIg8AmkjjonX7OTwjPdEudjaBcJYBzV4
T8BMoa+lga+qdTuXhYAf9H9nLa44/sl2YWYBr2x8O1Ps3rbzmbNFnOxqqOjcxHNU
/zAc0VDodg8OzQCINjhpTdeOd2x7FIbM/Lx0Sm1XQOJrb1YuYTO4PmmJQnFIlK3m
1HU9qBhn09i+XFrbdFsVHxV47MVlEDT7xgLH5DmXK4bpCi0xZuqcFf60vTs3OWwY
Bxt/ZdMFdijjQ1Zat/8IifjayYLMZB9cGM4FNtttms5PBwLUbFTlxJeJhOc4tRjc
kMK6KXTigQ/UjqBLSURQ5vn89bq95oojvSBYf0UnckdAcJ0wKWLvnm+pHp+ttP/B
BcB9HT4u3hGzuT2EJNeWQNj8ge0/17bA8t6pNLi9tb+kZUfABHbB8spV8Xg0ay/c
TTKlbjp1Qs/rio22UvHWN/+A4Oak58QGj3dt6KCgmW+i03a7DkUrL44Yu/MJwAjq
DHZJsnjorZvoHeglMT/Pz2oxv9QxiKYpfnMsyIlEC9E+smYV1qTFq5sGHb3N08YL
qoVRV7kLHN2lj+lN3gPweoxLBWnEHmrW7Lbt3DIfoFssZp7ubN1YjFcOfqm9CEaB
Ojm3cqaLa8V4dEHrk3WojxIY7YOBt59ReKasDBfjH44HvvOO0HdAZ6AtHcbwDSJK
t/kXlZqgduxYPVCh53Zjus9e22aBNFcHKk7GOdD8U+Bi5J0igoXED2/X2GacbSTg
/QdIHPPXQfzkgZs9HmOOcXr3wIp7IoTfp+6ZKO59BM8NU7YjEWdQMnIw3eB0t6pd
v18WKelCh6W2ZuICz7gkkxYgyUONhpPliG64FLZzgp4znqJ+Pj0klJltJTNk746w
zVwU5/t1r/NqaooLJII+YaK2qkLPORDwb1UgF9uVJBiw+mUZPLpSPS/CVPdnBoqY
0cswqcH8j+vZQ2mfwEO+A2NwGrjn/cL9ID5brEU9M49W7wMHzSz+j0PzA5yjn9pf
mZIHAmZNe9d3h4vpJe8j5XVFtJS4/mEWu9/HWigrChTkuoHbtv8wxLqnfAhfTxba
8y61pYSAog3Yd5zIPyyExiNYVsRL2MPC54LF+26C240fhmyNEnLEoD3O9k+issrx
o4hmGRJEvmXrsmhJA8XqxMurun/t2aSxQ+FmaenWEYlqyi972/qlQAM1As15r5Cp
Toij/KHOWf1jfA7f+/4t4yZvWgTt8Vdcb4fnY7YLzZY=
`protect END_PROTECTED
