`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JB2YBenj0wU6DP53n8TIp2Pth8GnT5MWsDE6IE268bZlKAjs4MVT4p2JyVOev7Nl
cmnMPLxvYJv6frSc6amubCBrhcBTaOZS+qaB3tPU+YI5o5WEguQwj9GguoWGFAw4
klyI177hs+86osIOb4C4WIvsPfPOqOsJ4ksgKk1uL8NJFDhE5h16ThDT59ULrj6r
W2/hLpi+3y07cfPlarmmY3195h4bCQ8GjmXkn6nDcT0JiHXGM3Ex6w9VqMl/gwro
RbsCiAGJqDdojXjOHQxb8DeRzSRxvc1KQQ4PA1WrduEd5vHNIp3KDOvbGS5McsVi
aJnEy6fuF9dGMZqFVgCRxUIjVIZLKqCmdasaDVykkG7FhUODppBPSWfn6ngTAz0w
3keXNI/GTLSsHOrq9aMSkjueJZDB8nCGiOVqcI+zD94=
`protect END_PROTECTED
