`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b0z2WgKoRtPJPVatKARc8zmWv9NLiD0eCXkmprYf2NlwHvl44ZzhigQzXyJZihRb
GgDeAd+V00/IcGoPtkLeTld6A4GeC0dILF3384XFQFA1MowXZvDfCzCZYimd78iZ
j6uVaRuGRaQKZIr7l6CXkqhXjFA04JaqSPI4MV20HuwKQ5Ud2vMYeGmxQhEgQt3D
n+tu3G6MwIVg/GNseMFj/+K/QNP/KKmggoBr3rx/QV1d0F9IaAaEfeWYjgNHmE/q
ka635nlQ2yfPhI+3McxgtV9b+lq24iC7k5Chd8xAC+GMD583VHOKUBMmx9RKS03A
42wqorH0PKnUnXaXNP+f8w==
`protect END_PROTECTED
