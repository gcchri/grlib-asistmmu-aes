`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kFP63fjn5aciLbxsIwoQF3+4x/5AGxEQ7g2oFXrYm/euSBfrZGHJPulOkUIwOrb2
Tx9FUy2qfXofm8NN2Jt1CQWRgqCH1ygrcWrlznGoOKDF47q1cXEFJL+s8SY1tWoq
Hzlg3bo4LU4xUzI7kKkblY1zwr/lYj/N95zF2Su238AhjZFcyYRveRn2MQeE76i8
EDRx8YoghGw5mNR45oawRiFG+HVBQhlCld7/ebdUSMzMyyE1bXDj47yYZQJL0K/b
EI6WCbO9Dmjkl10vWeB7Lw==
`protect END_PROTECTED
