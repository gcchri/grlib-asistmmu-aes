`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i4Pln5ZNIVaH56bisJ35l7W4PSL8Dgmo51uAAcR8lSVtqs+dKI0aOlUpiLe/m9pH
PHWWAAEhb7X+x8NZNIeHtqA+d3ASZdnCTpGQpjgavnNQMDSyewh95YKFeCIBYehF
b8k2ZUfVFxQuMa6zFjcGcbC3h6NNq8Jq6tEmPALz1tPRWqC9DdCw5bMx5IDHhh37
xu0/WosmYrOQ+TNThwXnMzfVfUZuA1mDSYI/wEYAe9nVTQkmZyKdJrnPns+mCWcs
4dabcIfYtJ0PG5htTHwLErZcn+3rWrJLMOnLU7yCMvHxN4veLiAY/b3ABKSb2/DP
UQyRuacXKdUS9cszaQDpasDjb81pyXJfGxRcmf9xuQ/Vb3j/c7WALeQL9Y9skWYY
JziwOccIJeLc57CLllQrvSg3vnq3OpuZBcuE8Y210Xz3ZRcJI5BA1iFOJNaW6JBg
cjoM9E+1jPdYPNRUT7kC0soeW85lA0+nTMSMiWk48M2y0dk8usAQoAblV7ku797O
LaHzF+FPYMyeQBQD60d90fY1Wiq1tXE4Eau0UOit4uQCg6/KkNZAMaceAnf7dJt1
wrLvbsf/UFMCj0PPPRuwO4ImYmFO2f2VBQXz3jCIL52YAjdMEFiCEnkXvCK/BHnE
8kMaF8xwLqGaqI8Ia1oK3m+CKuFTFLRgVwkNlUi+I2GB6IKauJrKiX0A1lX2sY/O
zbWySlrYc9LDBLMcPhk8A1FRbPBGm8yhLIWPdBG36GedlIGcgp1pbWs907Vau4jD
N3mSgsBwb2MPckKtEAmowWVStV6iC+gfDllCQax7a7srgz/m/H1sYrSJHZydwblG
6UNzvj8z4M2OWtETpaFLgj9tWI7mUuiGHLW3ce4kiv7x6n3kRNUKOeXqhpKnlsAD
nUn3uGwRK2jmuwEpPIpGBp9pC9HOhq5xguwrrdw8DmAT1nouNIU69cIJQZWK8xkc
Swp/ZYCnSTcm5MS54YjRGte+KYeT5/ExWj7Isy9mWbN5XeseAcmLQ3tPzzzYUKEt
N0fteL/RA7sLbNmTjMa62jd08p3YOoA1dOpLO8KoNHnPtU/1B5qC4EozOQTfhwkG
ecEQ03cr8TyxF3Tjl1QN2WVfVi3PZVnAuVAPj31jC1CxcBmshMAZsS3wgYDiQBFh
Mjdg5y1Rrzb6aKS2tzUboYDfNIEu60zp/jL0k5OXx9JXVuLVVgV7KiQFI2ZBYSMF
x14LgwiJSZcCIXOsnMFeTtWYNB287kSqaRcGSF/dSkRoi1/2Quna5E84hvDl5HdK
IXILOLgx32Z64IpgKF7B+sMJBN+1TE3E/s28XFaYGUWcS2cKR2ZqlriLnHTQ0Uok
SEqlvznCos5ss7Ljtw64vEaLmw852+jv2ytjNWBlRle+K47LL3ttlo6AuWY9bzUc
ySrhP2TVAYrYNmlwr7AUolUDd7t10eo5/LXaRGLoqIasssDBPIMa39092Pi4SKTj
ax+R35HaAZ36KWuN+dDjA4KKZXAcEPL2qZKGWyF5blIiSHu84l8HIV46vlMcfgU1
aZSH5D4w6rygO2o4IUmRXc9elFPj9vB8XdCxHceW/3UZ5MkaFFhW7721J/pQ2qn7
PA2Z1oEUB+e96m2esvsPLeUY4Qj/KL8dvjdFTg6wOSRIkJjzMght1CAmyeLFG5nn
bLwqCMX2bBs6Tw5ATg4royC1Dy0qbzEnRqXjyiGmdRNEHXryF7CesBsVncP11OAZ
0dJtQyTe1cfkA8qJmlF0FQtpMI9fWcNiWROV2gnpvq8H2VssmJSrCeIpc//jfUdy
6wSiCAqy/vTptDWgg/fXJHdPfs+CZRTUXVEkTRPFXf8zNKHT1lAFIqeU/5bs9s4r
`protect END_PROTECTED
