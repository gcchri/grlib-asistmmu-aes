`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0hITf3RMWWHXP/z+ldVoGoPVLRA8BFBJ47HwB4GZOfPFmSPcb0Ina1rdaXA64eJw
77Xf5GTFiGsgetPbAo1q88dX7Pk8gvmcmgmzyJGOc6udYsPm9XPv7sTvK8CCjXHa
mwiRLB55d56tE3CrX4BsGiqNBj4yMhlq3xa0FdRUb+TEcIGNC/WZsldI1jQz5642
5Dl2hNc8QAlRSGTjgFmAFijZk50UCdKSckhu2FY3DkZasmezoAJOzO/uH1XF+TT1
IbYu+Kh4L3vObKtWdtMr3HNbFJwSeyM8ip60NIO2FxCBri134fAscHItu5LtxXMj
getRHIzYjN7mOLovoOuSnzjW7uQ6Lgj0ZpwHjoC+y6cXFRMqRYGYT2XdB2gTtyqt
sWhdqHPKeLHbtAOzq+mcdA==
`protect END_PROTECTED
