`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FQuQ8QWpXeOPA8o49zQRRbSXh6fLcarUCQXLq3uE2ZCcNjUeHHy7mP0FoBRhiQrH
chFr8B24pVpM5SMsaid137wxrGKHMffeoXE9YqxcAMUCaN10H2WEqo83CrAvfDlU
dNQZhauw5KuxGmH71Mb0PftAiOdoIqyULQXWcj31jnw1fD8S1zOI1+iidY9MNVkj
juhOQKtR+TO1Hn/BDQd1dkBIx/Z6FNDdYi433zHjL3LEk9HE9Y+YvAG5WaQKbEdD
qu487T3Q3wFVGKejL6uLA/uJpQU6zxYjr9Ke3BV/mqBV1zf4xocuG7EdfQQybeRZ
i5+E+mQQti7cFuSMSeO5H+4UVytA6QpYm0RTrCHuBM72+Y6d7VVyuBcZj6j6K7H1
woCPNGESKBoJiTUsQoGsr93BTR1ZS3Ni83o71R40V3s0/pxTlDvgTrzY7K4s0OJE
Pn00io9PTiKTGjofb8x8yHvdKrvaQjNmb+envoJUbA7O1tE2VctIFYeBjXFH+eyb
obLRZHzswXUZB7SHhmVqf1eDzMwj8scrZEZ/0uNXTKS1chWxWLgcaCAQmMEJfo2m
j2uSvfCyeEdxAndmT+49XvkzaAP+LhQIYIGkxgwVI3lRaFgIq4vcxr19WTsgTN4e
2cuF8Q3Xz2ow0XS3q+zmGdMTBmEpq5C0M/vPeKtzh0SVaq4/Ljp1UFrCOPG1K/78
FB+zShGwB/fZFefInwQKzOGeizgOdeAuPvVcvNL1kIHktuLNO76B5J0DApKo9KMk
eth6ZtXzjrRd3rekurcAxfkRRgPOyMdxnfuaKt16+atLFgKYMZ4rsupaEnNwW5eW
x5G+gAilKHVSMCVuRqJwG+jdLilmHIUWfyeK7O/+lHaF1C2Db9NhV5wFVvD3UB2p
7oFwv0UQ/f1zPOhLxe7ZlAjt6/9q8vFynY+Q49Xw4lLgnrS5Gxfcx+wAOS2bq/x1
QWf+eu/rtqa/8SYCvd/V7L2TVrb0YiYNNEh2KoY1TRIj1XhD89MqOhF/lxyFmtcs
ms4/AKDdAxT5MLYWRALnGEbFMAOQJrLBYQzcYoPl244SKOFnpmtLXA3MnU4PuoYj
9Y7UKyglE8UOCjq5+Ihdobx/ZnoKQdQQ4YFRlizTnFRinsGQyP7Lv7fumOVVFrJ8
UjpVS8c30uFc3i2b2ez4jqzcCSCrFnOayzN5OlE46Lmurvb0uqXGmoJRnKe+MaSV
QFR3BuqViCEeqJ07a+uuevOgN6+pB1rsNXftBGuEEscSCO2z+KOK50H77L+j09fS
/p2TOPJ0Xwxu9gMOcD2lcM10A4s4PuxJwDVN2Dhrly2h6+BEVZsYRmjp4iczLbiJ
2ooMF2vRza2Bu+X5tC+jiZJSPium+wawp6HZJ/sP7EqeuTlqG0EOo6u4cs5+7taG
+uY7n9bguUH//knOSrO/dNbPHUoW0aco7MMcI3uOOUs6D28mKfTux5+KJjh6f8Zt
aEJUi4w5qcHdYhFCQ2mCnm6lmDF9iWFZx1DUVwnynZAohzJQ2g1SlpIWTB5Oi3uU
MA5l+/QFk2qksHsZsYtLiWtsIMa958FWPtoBoLI36nrz8wmBpJFygaAXO7kkGsru
7mr/fuqb85F9O+IKbEfqrCsJmvZKe01HDFe2RJd9UiiWUI1+4tKJbSvCMSzOuRSY
wVviD/7sf0Z522jpurbA6zM6HgUaew7PyUPB50RbgU+zyov9jKJ2bM/0cQu94bdL
uWLVv6/ZiWp47ZzwF6PEZdVpbz9TNR0o0UTt4MfjPbVwi7MIppBpkK7YAPu7nGrX
vzFMf6hbFuXv8+Qaxr0oqRS/alRBmm5Tl1tG/42ANrwYtp3JYZ7xGpuHmaueo5fk
S1yBVRmpGvvIW7gIn3ZFf9yv/rsrlCLZl5HvzUytzcvr98796YPeiTYvBvXUS3m3
Kkt64yGFEcnAeAzEXH80HrazB9CXR5DTxN/xLS5iRafN9Fh4eq8jwWlLed1DOxwl
AqNDzN239tFfIIglRwRkfm/0bB48d/N5bnBJXyx0qbc3elQVLkyKCi5ZpuBJlhBm
cO1SYGpyeDYZx7wHYXezrxEUZItMnm5wGIBY2TtUIOGEOYuXxXgdJ41xhQs7u3xU
c2wpzc3VTZXhNhhyptHldvX+C7QTzwvFAIBa+M0nAAEuCy7urqHifYUgC8FWuCuQ
sRmJQcXrrZal8XMTO8drCS7RlmTUaKpXMWi3PS0/seox8hZJ9pkQ5qMQH8KRT7vR
1hEV8ivUWmoUlHBUUilzMqS3mw5QjEOCZ+R//SOHER4zcPbnXcZ31yhsH2jtpQLZ
Cp9ak7igacjmdwJnZzd6noo/Bx65hyaWaDEQLFrE8SXKzPHvANnrV9gca3JCo3jf
iW3ZgNM7WewzbJiCXJJvgLxBSzjmZc+Gcwh4NdvLVLWqzZVT44l3XrSv1g7WoJKb
88koVF6Z2kpkNe4X8uw563wqMUo4TZJkAHB1kizKbHLNf+nqAkqJkzTEUOoC57VN
CgfPiaAkoKZd2mC0FfaH4Tskke+gdL/pvddnyA9cfnnc9ijF7rvtprroAbBn5P4d
rIt23aAzRM6mkOMcTVBMaQxNIKMdi9HRqJEvbUTu49DcKxx+9Fd4X/nzGS/CGvDi
6iPx4Il6PM14cO9sTGYykuw7GWj6dDzaL/C3KSIMkH0ru5JE2qehqdDN0kU8S7J1
Vt7zsJr4N+qsfGHWjoNky8J5wzXo5vqv1vMlTmfglZQZt6H6xV6vipwe5DKL5sC2
JzT1Cdv1q3DEH0eaWKsxLdH3mm7vV1cxBcP6BZjaGcjx8GrD+lhhzMGWwr80/XeQ
r2vgcgiS8S4RP+QbURZOvO2tpNSjID1ZA2NhFQm9fBDHPCe16pCyYXSLaPWJpG/e
ZjlpbVRIxeZNvQIj5MVRJa3tc0xxsy2HPR0aPIukqew6ZRbfM5UB1xSzYTgf8vFj
0YcDO5trIOqvaV1uSS7HWv5+MmlTvrNAVE9HzcBdoIjtAmIfqlY3GUcQLOuMpRXN
mLOTY5ZQJuIM/AXNZYE0VCuWBEOF827O1aF6BwmElKa/N6bdmkFmWXRCHDt0DmX2
2Z5g2hTuf4acXOp5qaOn9hFC8xP2s49fnbWg+axA316wtcJX0GX/LqPYdExV3Vac
kqIs/Xul4qy+oDfmvb1NZb4D+BiiTVZ4CPSqJRmlVHvsYRWCEKEtRzAtIkJ9oq+r
Yr7wj4Eb3MGs8O52GTtW3z7QWIQZFPPlfqqq/J8FClgzCtktPhCGWwoQp0kbz2zb
ch06+/b06/ENu4XX3tXAdPxuOwKxNV+lvoRWbcy3CBKmm1TRqCyothq0fMZZQIlM
kx/h5gdXo9ViDr9mQQ2MSPD/9OihFrZwaIPMnpV8vsYr3MWs0D3i3eXfkVK2t44z
TrLwj9yGcLV5HnxSodtDPFzmtSAHeM08i8pg5YMvbFy+hUOjSIGmBRwkhgaf+XKZ
AMO8jnXzzW4yhDoBLTznAwwuuu0sK1Nk35l2/09MnJmQ5uns/McPj6OGKpZKN+rw
o5RXUDgX0u1czK23kZiFMMaPVGsoi6J7/s2rq6lba55UfStf0TFsJ/8gWymE9Iw+
wbfICpbfsZ21lkdzkqPgIeJ17bRps/dSa2UFnmsoFbU7w4cZSlkDgWP75luiZ9Py
/Gyn7ryYRleGoSdZKU32oKvhOB4G00ki9tXyHlcICYwtFuNDH4tKlcYQoLQhtLXw
LL3AnagzuTd3nvw6Hgw8kd4X5QYiA2zuLEW/QGNXPvKlVlB2nXjSNdDgL1YmNFiV
7I8RT3bdYB0knS7j93I9tlZRHHOKiQw9XUwRw6qDR4Xrg+YF0DsKRgvpv9GtcVu2
NF3WHs+Y99s6mCKDxjZ/07s1wFH8LJXCkggRwRJEGruM33ZMF/kn7IQR3IQgcCRc
mySS7IdmNNYqMCsIhC70wJuTzfxpmVdL1EPAr74JjrQMHZywYQdXJsn3rwObhcYU
8ZelkB1R68wlVxEpWyiwkjdBuu/kaa3lQdwWBhOnR/MIIrUXM5/9FglJVJD1b+pz
YhmbkkF6iYvP7D8t8yQaPjYHeb2DFC/Vm+pg1CLlwQ4U1pT+Qgh2xlG1uOta6eGb
9x6sJ0Hh/r7GgGE9yPZJqzM35riK3vNJl/MdYCYzHxeN/8IZMbB4L64KVq1zjuKL
lzcb6KoezhgdiIHUKB2XE8zITgiBxvhQ6ZX7rQUM6U7CuiDvnrhSjvjQDolpr0QW
PBu/yjZIIU5VXrZGoYnScwLOhJiadDzCP7E3Xo14w5PWxB8M+GKhgD3aKMtDBjAR
zTPo/u0BaBZ2AGtLjKQsWRAMEYfwWAzrqreP/0CD2uxNwYAIR/bTrpnxIbDQYVsd
aOuVfmn6lbqSzwvQdtHSp7vYMrjwXz/r5qSv3dREbPRV5tWrB7p68uRmHPc9LqXI
3RrFOVBOVeYtAeSiPGr7jdeHJY4hJjUOS455DhqxoRBw2y40wnwPrg/66JRNG8m1
JxuW0Sd8tCKKW5T+KXnajlPW+gyvyBBgolamt21+Jv1hX39sJZ2cvPWEsCscLWSZ
rQ0EKmlUhpuAOYwWEm62z9+ug/a3oLDPxnHJpD/YMfDdJLG7+hNawEsCRPexjKTr
kI44O1AyXHGAmg+wKzx40niAI1pGsHYkM/0Ig95mgyoeIbsVCYhcJpHlhwyQzhWO
ka5fZTQWcMfiq24iR3G2yAh5oPXxZpZFOxlHmAZXnyzwQlz1SKHgMdBXXjhP/LIi
OYac2dTzMGLF2g07JcQPHv+Y3O91+EFbVW6yB/sWUdnMINMeTyVsZbuhyhd/6VGJ
Zccz4/P6oXNMCo1czYThnUVCaIqzhqOTvLCNwtidUKPikS1Fm4HcXVjPZ/Qu4qEy
PDySPb6uGpYYI/ZNWX9QvneXOvzP5G+/UytaYiKUfwhY6mn5l3YiPN/2cm9uAP5K
VRF2BR6p5wH/ljQTi/nT7iLlRCqEvM1tjsON1GjWtscL6bDiENWIf6eEY6FmlJNw
ZwYAnUfY079K4yxWinEekiJ94MA7hrIPwAeFRPN1N6UvWOq5AHUoEskKYRQJLTIl
md/RuIf1xT2nWWUN03f+9E3zbIgbQWNN6XBCzBnWJ/wPaRWkybqC/IvYm9ydUNbR
0s17Bk9JrzcDLXVjASbk4QRg1cXL+vMe/ZcEUcQRyJVJxZFHAnfVykQCg23HIQCo
QV7qbsK4cmy8xFnFox/H3Q0jJsn26armTJyPsZuUWxEVaf3yDZdHsenmmwcUMI8L
cAWogj3JIyHf/ZXbyIwsAh66jDahk2XGqdooQQpIE4cMgwwaUG9un0QeGBVurATV
Nm006cvygOhFuZv6XbFGio8QLITGS8h6ZXQ5pczRcEP0qCjGZPkBISrMedVhrt8O
qh/B04efu/EPJL32C4WKvbGZowaiIMCjCYEOLnBdPJIWS0NKROgoKPzexGAHDo+2
voVYbKbYENaF290osgEn7SShrZtLBluDoqf7NgP4kWqaXMzXI+/pYXwRRkCXROcT
Au2Z/Q29FriPFqgz3X6O0IlBV4RiysuSC1bAv0ztwPjUBcYeMkLwAOz08GxImM/h
ROCYu/QKl5BqsjlZLeTNnSUHIpAQzVNukRqZ7p3e/0VUC0RhEISqLUV8i+T/WXXN
/dHt373z8MJw9pyzMSorMtIL76r2xh8uCoFlA9rt/n25shNviQK5X5Vu9sJEU8pM
J3nKzVBUSp8T39uFcPu6y0wZnWGf62SRexJQPpzrtIzSwhB0MART6fPPBQjbTbgk
qeGv9kk4lGYmrE55Mw8jXUjJmvwdhbeia3PghEt6/oYnooeXMliGV6c+iy8a+nWV
+xujyifgl/35GQhtBlSFZ9FoLybejzJCXrRKz4qhWdLINaYvQAIpdVBeZynkJI7C
Lsgcwyo6HI4cOr08ar1RChy8PYUSGmLebjp9ewdnyiwwZUmFm2Wy03T2dMDoCNy8
hNxi+WfVb4BcOSGXqmifxRdBHUG9O3m1Y4D1um0lu4D4Si3rnCuFHPtZF1qPB309
aSc0xJZDli1CQn/dKdCv9v9p7BOSpvPiLdjALtJQJZZkrVUbgZ96CciiuEnmuMMc
YhltS78Puz0lgpj6af8TzUTcNhTSdxa6rNTDlg8ebbb7IT+PPQ0yrhDTpBUXx8Am
G1bGNMpgQbyodv7XPGFRNzUFP46/triwpeK+km7RZ/z/9w++LCFzkD/hSmWIneSL
alHAKQ47pf81QCg/CXqddVE2VIR1xLc+GH12jGTfVztYjdlGtnWnLkyVZVP3a4Bd
tviw0UfXrXT+QuimiWeRcazwIfWN+yfzCtGRi1MTmXsNLRQofvwt8Ubj8s2flyNj
r56a6jDgfSHanpIrBk8n0vQYuU2zsMhd5GltD+gpTl02R1cXPyzbimKT+q8mHkix
TE0nHJ5t5JhXV4KGBDStm4fiR32WE21lj4OIAGqTI7n77AKXtWbwAGGSL+70y6fo
6FBilbl3/Eos89KMcBK3LtuJYdRwFpx1gjKi/MTLknH5qC0kzFhXTlODJHfexZPs
pXf6UWYnu5Q+6UXpYs3HjdPIsguJo1NRI4P4OfQjHrEpnxAaKj1oH1acru5qpfo0
lOdZNxMrWehKK1VK+gTjkJy5enJmkMnD4Oyp9218N2b0KQuPJFbg0MAEJ+5zLJuc
ddINYXlxhra9a5eiTNasC0R7PZpJmomnN+LS5XBlcxLZqOjqO0r9WIfAoQ7M1stx
hz88hk0GOQH4WnftUXG1/AOK2XoOUpDqZLtSGSkLlG9ny613OM/1VMMpirEFz4iK
l8GNlKeqHMpSieN3vAr1tUF3M6nbT7Z1PFL9hsj0BILhqHWNYcOZRCyeFC5IOQh4
ei3NN73G55k0C+UCOKFKazS7pUHbCB+hjUsOxRxyVPJeWK1zQgO4iGk4CStfs/BI
zWgobRwWG/FaWAaov6BXCzZEoyo8lyaBo+EFOX1lma+2RE0/sCcT/TLF98rJsxjc
B9k9I/5eJAzc2l6uYj8RCjdBctNEbvIGdCxgzxbKeVBDvehUAzOcZCx924feXWqU
ZkKGLQqveC6x8nTmMoIsQb8y/6uteukV6BGieI+iWxd3APvwxPtadUVGg0PEl9V2
2lEa00kgJzQaEk8E9wE1BK+dUYC56AxBFGksWvaZbVI1tM+EDpo/sLnjZe5IZX0s
OB+CWTfPJfdR9LuJKUJJeESgX7DpJHknvOsCmu2gjrzi3BL4O7l8HCym+acWhooI
J1yGbpUL1hhbVeWD8Q/ISZk1hWmaTKFV2cnHZJxpqygFc/h/ZQAPiQrs3f6UdfcK
7C9SnX41ZdK1HHYg20kBmsaDTVAqFDlUKSw3r6oIfjl4Z+bbZTZ2YzEadW4vkHP6
YU/YFQzFr5aP9caEa3yuehSu7jcylihwPcT6yZIjGmFo/tapkE4RiT5MW0jVGwFM
QqZ3kl9sywbq7apd+lFdJ260ZCxkXWoLIcqwNpRN5RhEJezWxxblGZrEdT2mftUz
T6eOkjiwrX/APOWz+mKC6HfVng3wPXwZhhkYOqzxY+BVOj2Xq6lTIWQ9OW0pBufP
GrfBmdC/EL9r21boPUAXfwTLahreolrh5PqAfYuiGAmnAb02Bm3hhJ9O7TwZFO2G
0qQvqp03nV/BCJAhFndhraR1o3U01ai9HypLLKvhfRx5CthDUyZdT6wuv+i/X/Eh
FLT/+pPxk8UgbiuZAcUA+hiQR9gEnFtgSwyzO3KFuFUngXjGxjtuSCHOTP3EosFN
O6UMZdG+BaBboHNjETqBclZLwkjpxUlEhM+dT4pMGhNjmRHEmLGL169mhALpvnNj
JsFJ7Td9qVYQvDhLD9X9nOgI6vtf4DvaGWrT7yPr5Z3M3Qu/d31F+5fUe0VptaTZ
PhDtwWjBQtG3Q6kSyb2IDFDRsMnYNpkYk3ehrfwjSMigEgL2RFgacPLsXsljLTB4
07F3DP5EVDPfp7bCdhXRlNyGItH95zXszXOnJGmdCQ7anVMK4eXIyIam0OXIggBy
xzdmVMEPHv18KIvuQHoDwEXy81fyTU+XmVfby6OlHRZEhSoC/tHnT5xP+NfYj3AX
roxnPKQFCdocIwiFaO8fHMEMqcNwEqZcIjQcF9Al0ZF1KYfAqms0mspiprzCXPJ0
XLuL5SjWBwJU1Gh4LMjeIYem5yDLooKxHCjhDlyVXA+T4knusZJw76wKxFi/3p1l
x70S9M+7TxxS9MOxxePpazHUeB2ViYIlQAle2sgc0G3FHyz/QzCCBa9nXpRQ/0yG
r1FKlH1qJD8POTlqOK0pZBEf2huFcG0V4wTadkaUg2Yh2+4znxAdYHHqzEkU+rLG
m4bUa5a6Yxcw3hb2iYpybssA0VgSX+LvduhV8bsrEsM1UHGYQ6vpVpE6FNtzIlOf
HUJphfAhZlS9J0ZmNGJF5MBsQpMkBRKqS/xludbng/UnPVdHYMU1O/3lX3Hmw6WM
xrxM07LEv3NLThgd66ONMGTttV9HZQ8oaDK6bLWPypLTrP84ZvwErg9QJSJgOc8u
btHOdx78rwHLGHjaQtRWp/mOLq6Nw7aIxIz7JAmB2S5mSBKhQfNuaxAA3+5MAR2C
WvOxxjZHe2MrJidcpmXOmDAtqqyBB2uxlxkbhVhUZoPHfVOQ6ds1cEyaS+qHyzor
4KGzVNO5uNdga++9FsVGw+RsHxRbZMcFMBbkZV78jmTs8zevPfBQAoGq07+16jh5
3d/XK9X9ZSCTT37fnKWQ2tXY2CyyMPIafJAh5+3D+oKuL65MVoCb/XPeFexvbxvA
lfctqzNgb0l5tUOVqIPDRe1SdGSO8IZsCadha+KtsICvYg2MfitbIez/1zUY79kJ
W0G7pChBrlRHQNzcdGA7rrYQkVki4idk1nFlRY0TpL4alccV9EGWlPV6GBLUYsio
G3lDGRparawB88KJZzsoADXs9fjD8+ZVMEBDSiH92rcLLP1ZXT0yV8m0k1lYsfV2
oB4oigVmxptoVRDHQ3ND3WGojK3bkFD2R/MAAk0C7n8pSsaYOqT6CtsyJPahVyrv
FmPVDxwTtTHv3lqSV3N9Wl9Ubnl0WY3D5B1+dX1orCpf+MuhhfsMOz0CGYjCISq6
V65Hukbvw40N7ROn8zo3grwPSi6qS4tXfV6PNSy2TB/G/jGGlfPwBMw91W/8QqS3
IrkzOFQvvX7JfDT5TlYxaI6NZvVRhqaO1L38MQrJSILQNpGEYx7QKJzqDbxODd+S
C60Smz8Mfe2dalezpvx0aQOmBDN0KYtSC4L924bfKL3gi/Yph7gxA8xWW1trLW/M
QnlSZ6Q+V9oATlZlAY1H8qCR7XB9gP4YtsaLOlgs78GCKXs6UzQWnZXOPQjfbIFH
MS1ds/LrHAwylbk4yvnPqANOZoO+q1K/TkbYPswwxqTf3PmscW6BYS0seLsNNtyV
YcAr2qDTBcEEW/2TwlNUHudS36LyLZ/TT6/CQKeaNHyGGnHdewiHX01yVVZIXnci
3XEHLAvgK15mn97GeBGVKYBxpBDbFh3HgfrhgykOl5TseKJn4p2F9kxfzccM3TGD
5uXPhuqkYIxhgYH/Yfbl6F0Ur497Lk1ABcyIzTSuEQwYNpodH4UjrRTYASqtdO89
COlk8mgDB+QSTlVfFQ809006mFlciDZeWUkv9F64o2GIlkKzGIf5zesEXExMNco7
UNdvEQFRgSHhvZOmtbRwNoS/yW5EEhuTolzPGp3zryEpMvSMzWBsTwfyfDnRbVjB
505/RrDnl/Hq2KT9mJI9VXoA0UR2FaRTRgzz3KaUCdVNmCnug20sfTMW6Z370sT+
TURle9SVQls2nAZuSEphiQZ/933XtVeXAKZ/l+tp4Y0fJktx6YMWlVC9NWgbKxpa
Cbt8ukJFOUpIjCJuvY+Ud4hq16exikdcNt3o38/uffEfUZFw5krvoHN0v5AWkD9K
i3vJYQZX1vTdcfCc8dmTXeGVEdiIPpbUG78FIvsm+XKw1LJ1qctUbspx+tiqlBmd
IwCEj1vI5dLRKKgOlwxDbYPI9pRLvWaqkDU4tp6wQVCnwK2zFIydUYuTNme4QmU8
80AhNKQKMeXj9wgoN5ZjjZDYIy6Qir0xje4hCOtlggRYAfLKrl6/CvO4/TO7vipO
F9qBPeC8/R8sZrTQ5vLu6oqhqOcIU3UxQuq8VY0UbllMYvtgbbHqSdW1zIAT0bQ6
iQPle4x6IrPB3Qh6s3zCt7F5AGQi86OsBabLyoj+OrJKazRIecLZ/eHw3nm8qXK8
rFqa/onWknzkuidHLxmUrpxsQGzFcvDwk5JesL4RYuApIWziSiuxZeb4xGanijIq
wJMnWoKoDkVdvhNdcRjnIlrjiuTrXLSEPZnEPEKmK5faHGd9xhI1dOVeHcJASmFY
1q6+Ps/DpUW0X5cvQKprP/xYBtRZNeTY3PntzR6itAle1v3/37RFFRsIjEuRBU2+
0GDWAiNfIGb96gUHWO7MuYYvuAfv6xFcbffy0/pgcmSWPmK/NdE1oAaMIQsvswVV
2P0KK8Egziq7Hf6siwCqUehQoQLIK5DKDu9awU8TV/Wh2VUyoBu3V289RuM3wo93
r2eHcfRF9+byDfv5Ku6APWqO4FLPZU0jRRC5BAWpCow=
`protect END_PROTECTED
