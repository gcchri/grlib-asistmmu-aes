`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ehWur/8s7R7ex2zKWaBM60cYibCIWzcBr9EgGFBparaqGmjY9eaVXw5tc9Wf7Vf
R4m+ILb1TLjphuK2a3tFxOC125/SajmvNK4drMXRgrQS14S277XESoqCPc+3mw7o
olN3i4PUg/Fn/HXsrTA1/RAmLQAJT6KiCDHRaWq4tKr5hAjM7bQgOmjpUUuT3fLX
6vXbEh84O8DfZwLjjSkCrLccZBWLLgYh9Q6Gcn88zz9+8LP4Uqbw6DElpt1eQAzg
CzVu0bRJ7qxOAAfUmF5EsFET5BG+pm8veQ9ef/0OVljFIqiUOQht5Jz5vs+U8Fwt
vGCKGKFolsxsf5en7MWaQZ28GaYvFYHcKNuXTAB2SQWrzjFJLiJD4kUaKrPAE2Am
jCTyaPd2E/YMxOD6hbIhpb1FZ9IiN8SUdQt2/CD7kTauZdKtMmuDaBI4Lyh7svHo
KA1Kh4NAOpQISFzrZa6uc8oXRLmubei2dDiwozKA9E/Pj5Kyv7dq98nQrlkzyZvB
7UZWLPxaKJlng2ZXfZL9uLWF00eXuZAFVhOBMbYatsYQPavZG/YWF4j4gsgnLHVJ
AyLcIhVKR9IP1rNFiqdmRkoVVGjp0OIbQp4zKkrpKvzuCLt5IrtPBqml+f5XndPa
Ty+l8F+KWJmTlX7u9ajValJXPbgyYK5uBHHm0BtvWkWCqCMJbNuagDlCSeFU6KnY
xaVU99X31NJwW0lEGcKkZZ60/8pJcKNTnnulPLVvYJUneU75hF90f/Re5ZH2YYB5
4imLcGoS4tcyw57S1Y0XpX+pMowmrRyx0Rl1y5uBwY71siDtvmAbYaYkmAF1MVIk
RNHVsM8p1S0fkMFBWt1RL9nasQhYPwpPn4ucO2MsJHtcqWsFdcEZjt2UVeg4MYCW
ljF//921PNj3ECkSWPiEA4X2YeihDFTf4H7WovXfE6AbEikgwXgaqKH8zCjLO8rQ
QC9Da2a+TdmQtQwtQ45hIRN+ruKeB75dMY/ia7egMx/QaP2psSLeytEh6IQh9OeH
Xwx6mdtGX/MUmvgOedFxSqS5oi37Z8VLD26UC67vaYMMdvPTbpUbGIYHYx+hkE8S
Sck0xDzO4sME1pkFhGTDlMAt1y3WwxlROkbOA9jzpLk2Or5bhQ9lOOF+AKGrtqey
NS9Ky7XlyZkzV7b2l3t5cFM1L56dYfZCgklEGywGF7nnTCi0taAmsvgFQDOHLcVS
0fga0vNZn2NHrQGcE2plyAmlkoHTvdpzveQXULH2q6BnNmBWDuIXpTcXK0VkyKnJ
9fVZGb7BgevQGvvSdicEGy/TuYWUUz9bBe2nCXCOpHNsAAjzZQO4ioPcLv/nvHje
007TjxwwfBUGV20afkU20rpAkKlZ89G5Wlrh7YnBAadc8KWCCB830LJBFZ8lW8ia
1+973R00b2d/1Wj8Djv4I/kz/A7OdmfSzPoUDI3sg/OyWF/n8DsOd7LwYYJ/ZDbc
SNOn7zUJ5tn6kzb5QYH5jqFO1VBIAs1RMaEbk+h1qfRomphtd/SOLEmedEeP1shM
i7YQWDTeasDU1sIttu2C6WIfEgknFR53rT3U7LI9kkleNFZXMjyOwH/9M6RjFmYf
YN0vCT7Dsu195+UuDKebABMe1eZrIafXLvrkzwTvWJ4oC89S3ZdcmoluYeG/6tcD
4aoZapvqkbYGY7khoP8vAQKFwBcZNcuMaBZBqH8oyMZB+WetrR3uDep8Pe3hO0nU
SJ5Vvk8mmqzpchI/yirIFIgCblTrueDgUy1/tOpF6SX8OXS290qWTbHXupCDAAhP
0Fwoa/zpt0TSg+FVCH9HLEjVivmlqfwXx1q2KBrTZB8963Nr8DX2Db4LE4PY7SnD
dkk0YkWqgdvgT4tvC7LCMtd+bqM8XOPxyM7tz52yxeQJiEKe4AiCo15OzHWwGtA5
Vy5NjhXwwTiQlYkQRWj5iKA/3bzdzJqN0ZX2i3/nLDSN/toih44u48SB0VkYoALv
Nf9nFtyGjZg2TkB2CnDAn6adhZl5kagtabJsmn7ksxFWU0WZbGPSXUusqd9bEEK5
`protect END_PROTECTED
