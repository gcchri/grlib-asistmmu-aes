`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dGQA5Lrd44DaAJdgnwQEnFqBoOTJDepmGvcbtvkUM6aj8h5y0BFOIdTXfm8hUU6R
OE9WWEfEotBHAgdpDzrzitY1kPqq8W8eOf1BefFSOmh+owPrqT6hg2hBP0fSwfIt
oF63pQHC2ar06AV8B8/9HlpSNApKCsWzrrm/Jrnd+DFVfLvAby6PMOqf5BV4W5C+
pRT5XE1JZB+/tVc99Vo4mJK6jn7E+q+SBwHA/GuA2dVRnFPHckmUKSFW5j4KHqYq
jvE4JV5l2Tlh0KAQuYztlvIsW+Tt9zgDcEm6eln3yECXZyhprXeZj3H35dNwIHNY
cbCx54Ia4bD80jSq/oFvKtTsefgqq3eYvFPgu792WpScI99J1d1LFXyfgDq0Ea89
8rHtTiu+tIZi3k9P6QWFujGS/g3KExz+mo6poPGSn/DbZ67vokaUhFhyDqTLqdKu
TLLS9EGp/Brj3Q0t6r5oIvKI/Ey2LkAQMZ0ULdFDR+iXdPF/W6Bw0sG71aFWi60W
FRn7Y39zsyU9ngGlfmrLv3xP6S9NvwF0gB6Lzy5jMCg=
`protect END_PROTECTED
