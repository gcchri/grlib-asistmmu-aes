`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ve5TJSbJdJrY3PaEv40ng5vBO3jntAxVFVDhHWSlTVB5PFFQlvJkZ7z9AyPdTv2g
XjrWYYsTeVDngJ/ctiJ2hM11HCjHkDzKEB9FaLWSOInf/grWwE8BKNgwOzLeTDQf
Jo9y6/h42NbtiK27qHMaCbIJo0Ox5gF+JBCc5mGXCspqfqUXvOPZ7R00qYk7LMBs
9LWAklOC0oEhh/CeQ2mL1jjeJNRsFHGrkDjs42dOrSzQxn4/063elhhhDdW5AXrg
Cq5IsxFreALaJsxSVMOqYmjI/hANjoIiIZOJbmrfQkWrL4+SPH/oirjAN8nw7Tv3
/JKfmHkWHzYheo0kBDTnUkSDmhwJQ5zbCV21r3hHSvZxtattvUcY+a0PSDjN8yX+
7awHSYem//p/qayx1Ah0PtEA3dRMAdcp9GT0408SaAYy1H/GSpEBybxfyVbVyaTV
gibuytPZV/oTco5krpehTBx4wHS2bomaqODCbIia67zZ+4DCldanrMsYC8WUNABL
QGjsSeUopj9YLWK2Bvp/bO+uMGdzaBI9Bwh//wypP361kDOTEHomBWjW52Yl6g6i
sF49KslRoyqq8GhaEqY3Ak9M8TR+NvkG1mFAkhW2WJ2r6/L0cRE9rJWS2BUSUZ4y
bt/XS94It2mSzc+/rPtLOmsa/a+ROgJKNBU4ljJVGsZ7FcKhXtcpt1d/cWWjGIUT
pQnEHwqe8aY3ZM6Q6Y1upS7/c2JX7IDAWss/WiPaVcLFzoxwvENwyuEeSk9gPbuD
smptqgmowbPxiyM0NrSfQyJmF+WY4tRhbTj8YBmCLLx5+ZZjaznWuQZbBkjEWxLl
ZXsq5Mj7fKzN81J7baj2kneFzg4lXFaWqFEQY7wfUIo=
`protect END_PROTECTED
