`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QovJtpvdiVWpcF/w5b1bOZRDRBsOkZ6AxNM5c3wPcd2eDhdvJLgrtj3YFoJ1xA7T
7Xufyr7NPWOmkeQqHnmaS581Qt2IJo6hQO98exkyqXyRGJIdVRETfr660uilOg5X
yLxPcZIiZiKf3j6VGWk6VP/5puzMMDD/261U3wJ7/Epy94jcDtid0FB+FQUcHR/Q
1nQd0oBXYevSECitRTqF2y+UWp+lJnmZysnJ4AzM9C2ZvtV5p+twez9pql3Lt4kt
NnVLp8OBQIyDua1+Y7lgZXZ+ruM2Yf0oQfq9ccuN1RgQ8Aipiv96gPfiF52NolOs
vHuNlePu0INN35T3ldEaMJKhhc0yQcFH2rdr5D2LytQJq4Jk66dQekSfGNFi4ZN+
hknQ4vbMDGP8fCbV9p13Iu+4OiRvGWtXFYJ3kaJjArJnJEMDBkwClHt4zAxQukyS
eM5pGQ8jGy0CICZUndpzCJ3z9YTu3ZN12dCLpkoysJ+D7Zf715nJYW9fhZeljIU/
MB/Jc1DRVOJaZDiqy5+5r7Yhzc9fKYlWPlCXjbb5l53FpiM339DZZAurxSsRzq2v
BceM09yw1gYghQ7noUACjsSkA3YFVdmOrb/1vMsjZz/LGRAZ3DX/bQhXmHsGkBTA
g+Q0BNyaeMByMfRsvz2Oo3WAfJywm/GMV4JyyV+fQLD6EFMs8KGzQ0G3aldF5i1z
fXeQ5L7m6FP87ctcNScvQXjoIH3u1320xGsbBOmftNZ3tDaf+eivs87XjK/hmTNQ
VnskKJpHLV0GqE6fvbPn51BxkLPdVP5iANdtQG0ZkHyqPT/u5KTYGVLe4QSRbfT5
Av4+iL9/xfRaVlxK+sYglGGhO4H82SqmAFI9pYSLl0htIy7KE2BzsKSJJvtXs2a8
vJAFz+XcpSGwNg9nu6HKu6Msq6E6meuH7nzzXskrQsFnGimMa1bHDNXHJ1PaIfSt
IIPZf4372Z/QBHNu/KBzZKkE2Y3Urf9syDnL5miXnKTtcSsfDsNgvoVp21pPpzra
6e5mi+FW4o13d63iQkDbFKEDk4vUHFTV45HQugvwUBD2moUf/n1f0GX+TVu2ujQ9
Eb/2HH6TacXCSLo8G3+zp8LKMaTnRxrD5bR0bIKvlH8178MPJ+wQmzxfCJt5/mIC
S4+UNHUhG1ObGjPk7O2sUN66nz8slNF4U7CmCKtMQCm6Vghy4KQGVUTaoAb2moEw
xnyObDDR/OHzF0BUXCnyXW4ykA1pKY1hMO6V4gg0X4U1dagim2K23QTJs2zRkjb0
Z0Tx1i+yZKFWBRqN1as0sPamSxVBHExfZTpPLDs0LnmJYtz0eDlgV8E249XGOnpW
HTzuY8Pd67FKSwLTc6pJvZG8ijgDo1jULac5TyaWhHsi9xqG0nl60p8KPST7VExD
A3eBt77xsYBTWG7b9cy76ndGLXY3E6PjQWrp5aU91cvutLF+AFdfvbuB9tvUOCLs
fcEtMlscqXGOZIrj4TXZzuoRFWnP+n5Y480oWLhyevPQuXLyejXvFp6ViBICOLkI
YSzYTEyWlbxesq61Ly7h4OlkJYmrX3GO2GU+McJKRKHjLrkbBqOBi8djqZelmvo6
iPtBn3ZZesw9z/DEYsU8dafm1TZZujCxOjDIMA7ouBmegKzYRIOLxshOGmSjvRcz
fO+dgM+9WltOAkSCGuPXhyLFVZY4hcYotbmvyXCwzl7RCGr8XhX/8OeXXMoxpJnc
JsPtthuCpFQfvuX2KUhWOSW0m2arTLTZwQSG2VHyeoOmQwBE1s4lLn/tiln3rCgt
Of6C7DSCI96wChDdTgXlkiv6OCSFzfX8YY3XknfxL254uiFobPIYiz39xg7FFfCp
sf+b9LbwXLGyFD6aI1p8tMlu1AQWIwlmJjHNqxXrbkUn9eMgzZrnmxoYsVeGKouG
mkIw5loQ69m6K/JjULQA90Kba8owLish8VyD61PxILNtAvXHrd9p0lK8O7sHI9LD
vUtRtNfWe+XqfHjcFAayl1egGQnLhOM3pyCkvYmON+Dw3/eahadWxWanT9SCcAV7
LuuK06I+w80a9rN7nj4HqcVkoV+cfEnhw+fHizeqlfuo9dMK/K1p3O51WWtGjsGo
35pbIsSQLgMOWTC9z3AK7rpzsL0yXplQJthtCVxVrxuK2fR2JuWak64Uu2BrDLiy
99u9UmS2qf9FOHPtxnyFqs/qH8/2e4mqqVXuziPH93oYPCMYEoLxmagGpJ29Sx64
EdC8BuBbEFqB1IwvCytcMngFjKIQwVWiZZ2Q7QtZLXj3sTW7rW5f9PXp42wC84cJ
12lLrSIsGvj4uMekEEiP0iwFrRSQjjdK1areNdELbW9iHwlVH09Nu/EemieDwC07
csw0W96gavAyCZiWme3nDfplDLotPoW1p56YUrSeWLzab2tEWsbPJBln7ezl770U
cYBa6ZxGGHXzu3QqMDy8qeCZ+k75gNDx+bAe7wwehRpCBTlc0BPSUzihpP7YbvlR
g0f0r3U043Voo2+E5Dai5Fl+qm5zZBNsov73aWo1gW+1SvUf1x2oWx4x/jg56+xQ
MUjXaIiDqZRUoLfrlRXy1580/rJQ3Rfhi1qZo4fwKTsd7C9TojEVXesptDUOxoF+
xufLjogPyUYHbK9j7G77YbnqgRneY4+s0CF9uTAJp8+AzU3/A+FyEbkx5u2qN7Vu
hjc4IBlOqGFButDheOzSzMWgG8rhg+ZcXD16XnO9Ycl5CIXqyupZ/d7m5GGPKoxH
j0koa5/zjMTetuM7eFZWWG4nlgU48FL2e3XVQh5Cnle7kBZd8nVXT+czb3n5vvw3
NIYzO5ZfFeqZIcEJz1G6pp+Bwp8+0VWART2uDS2E3qCJRofj6JDn52JoJsupUDaS
ftP7CzBVYnPuPk4c67PuebD9oD5+N75dqOlAtbBGPN7Y4XtgsIG6PFm7nBeiDaGe
LYSw25yqo6Vptq3JQO8GWmc+2AHS+BTn8NBE5PzcWSP4EfQsinmh8Z2KWsVkjwoS
9VnxflZP1V+Q9k9E2CNLK9fG7OQ/FVVNnrnerxmmDhGBCyKx9Wm9fc/QXf+IN4ny
eugXeqS9TD3HCyrkD9+fITMVI8oBZ0XZKvr3+gNkrerUjuHUvDzQknquzGY579UP
0Mbr0niYYzAsTeMfVrRsKLhLEzYzX2L0H2m336JvjRNe6+MLqWizXuXVrWVaXHyE
/ZMT6nDDw7SKMOvCdSZz0HJKvZsNyik2uK9uMDZyn/8eYSuEeWq+hqeW/yQ917yX
70xMqgqIPyPnPUnqUZbjTHU08HisA/wyIsaA5yIUWhpeSw2eng/W5VFMshjxmHUb
xpIO/y5aC4r/1BtguqOAYd7V+EWw2CVdi8mtANMCEerDJnmhFqR0dTaun/WO1LBk
b4XVEU/1NY9mkL0DCD/X6AiMZjEg/UnhiWy6Cb3BPhy9Y+eHzrlY0KDRf+PadWip
PRAtnoR/5S3vTJQDviv4bQCNujXBC1fKxEnhms/COTR0aPZzHHOzY0fV0wvzGc56
v/lLUPST/v4bNX2THo4iBu67+3GdocVyyQspBPP2ROnMopqtyFHlsODJ0TTqSdTN
GWou/6dekK9oPXhMPdnmLIBkpU9Md3fqr9BBIapXcnKO/u3UkM46zmSl9tUGZijR
6HhALdhyZEB5Q9y+c7Br6RhATVwKXZJ29j1i+wI4aQBDoUzHnCJZvkuFF2GQRQyh
yRvtf9mz3VK14CHSbXGpPZ7QvcPt7tY8Re+wA7Qufs6MhljmOnFObXZO2W8pTiU9
vDov5w4ZDCDO9Y9YbCZWwY6gJbCVNCsazmsAw5kMtrQDjcpVyi9CM47NrEC+8RcI
iFXTGe72Nh0+/wKtdtbMtmaW8/HdBnx9rtzm68AWophEaPhmmM0qsckdM0wrydKA
7Br8lJLUFmrPkj9hX9R68EOGKp3onyEpQG9tTOb83waEbzknu46qAISf7W8N/m8p
R08JqnhFj1qpyTnCM3Lyvdd58qCS5FfSgpClM9Ej0HFiNWZnssJv7+mM9Nqdkkvc
eaS+wTd1CG4NPcnHHpTbEjVr3RUhOuJTgnrcdEKFYapIhdIaKNQQHVo7hdZr8Q96
aqLVBLAnBubGZeJtiCGBcv9eHEiVrKWzCx92sZaRIbWpcuuXPawVdWRAfUN9Ksh+
YKMpL4m2PMtx8mDrIzEUXj0hQLDR59veg/1XVrEbq33I5qPPUx5olm7IOS8I6cgL
yaCnF/72iC8jB+/U/ckTEGITpNm3V7cx3mROpqSF5Ar1eOOpCs0N+sD2VpLqle8V
MbTIH8p/QSh6dSVbet5tyI6Fg0+uMN79yc/FDOz48HvKfc5hNR7d0RjhnDniYaN5
8GN+V6JTToHaMrK+DuahQyCRvtPlVL8BkhIgf1h0ph0XJfL2lVjwVWJAsr5O/jOj
h4DCtsyiCYhghoS4Us0cAGk+S/2T7D3va2io8+0lugX2FxR0KNAPwuzSAS+pCcpv
9B1v2iAs82DwMxBZqmjZLYTfNoobk8WU9/w/WXAQ6je6FJnVh2BVcJWZixysjkEb
jcqIS6lXuLYOVHQccO3fTNqfw4TZWOwmdVjnCXxdA+Y6i9buq7QddE1YrfP0MW33
L5eg4jBONKTOinTMmSY+IG9r3hhdiHD3olM5gTlTiZRfF7Use5kdKUUnGbBuXD4E
mRotc8Cjx1Hi9znKuPdW3hPC9fgLjpWFe4vhl7AX/sIspwIkKiwV0CQMHIJv63Ni
G5n/oZ4YkSzPhv6yK0LRHX4Rmbdb45gzGQAadUkbMinRnO/W0x9cSdQAZqzmsbOX
xv1p8XTAJ5zu9JFPvIEM0o7AQYbsMLEY9b0lB+Z0mZbtZHDfdgDxCr8WcrMynN9l
WS0VlKbpiFc35ngNOJBW2o3ZrdUKDOwFDdwkX0/0DWa6jJrr3nW9u//UaiI5NdM4
4SsYXUXIieqn1HzT0JXP28djhRQZPMK4Vuj2lOFC2/uwTNolS9Jyvv+XBNlMFqgl
0EQUiZjBmKPfoViYn8wzZVGveV/m2SftSq3h7Ws+4CZtBc9UinqGpo1dvv+lEwCu
UWBUzZjcKW6rq5GF0XKSmkje6bMDASGrNi5wnOIrZVGcw6l36U6nJeIN0hWRUc8l
VK8tVctOnojRMSc+ALz7MaC7hJ48PC1JC7UTfnuNrELcMX+M9MkeSQty651Q0X1F
0EZI6ORef1RS+AsuEO7WA3LJ5UQYeNyMJy6w+2STpL55bqhFgwVMkLFSTSnXwY0U
lAxspg2yEFwqpflyX9cBeUs8i9oA4MJ80zqOq6xxIndy3jDWY5Ero8UeEsIYd5jK
+Z34KLHc1DbbgL4V/m3QrH/UMixtrjlNluPNUjY6a5mMfTSe2Dhhny4UOdMjTYTC
SGMqUbDkPlqyAW48Th+RR/7O5pFADFP3DUWSOykbPYTgOTul1MIUNGh7/74OLa5j
BTwWV+pEFvAxRTOwVvd7KyfuXxQzuQLgNBUjiJVrhy7C6f6u91MG4ZurB/vojA6q
cCF95uFeL59+w1vUkoftnaQVn+OJ9Z2h9Sx+syObK9sBHWURMA/sqma9pivE71vD
b15vvGazKQSAGmphrLJfaNxYxaDyOm+ejjsr2/85RkJ1qbGqdnfWlD++V8hfD0xb
hHLVRCVtMOBQaoZncZdPR4AeuFmzRoBS4e+e9KyO9ohqU4THRxHhq0nXJosKJJEM
0rkLNo+87lu4XVWRq86ZG3sMYWzirfWXI0szEP9emJsNSNmKDttF0KHWncpghBpk
FICCWtgaFKfz1BYbiD217R79aMSvQ2EgWfh9p06J9Pitnj/r4hlEmCAfEapkpgHD
6m3ctHWhqEiHsnYdBQ2SaaZhzRvM/zM9YT+7GsUW3u6eWmqy/m281783WOPrXR4S
O4lKUryp0C5kyl+90ZPRvbgrmCtz/BvY/H06+v5Zj5UMijtklFMf+2UtTspZg4cZ
0mjmog15H6h31jj5A7ChR9BCHpCRXBIBomNgjAS7oHC8CCpFCDEOUcZioBm3DF+8
VgfrnAvNBfpRxnG19mbyUTjzJYe55unF5K3Jsa92M4YFmRDKS0eOUQ1V3KfP8zu0
4K/T8ccrwmADIA8FBEUcdEu4vChfwfRMmTCUl7Xb1ppxVNr3Nl9TEI80YvNqzgSl
X/I0pE550U+xpPAEip7gTVvj0kD8jTvH409X4yTHwlHAjvXIJOyMmf7oxoNqNjuo
SERX4kihBeaRl5DbLarOjW8FH2/f5NBZP5KVHNXk+6KMAvD1YatTl67VifYkg9jy
aRug2nb6M8Txp4oO7dQXjAkdrg0HHIIrf/raERDtgYRgKhGWuTlhrxe3pm+lOiV4
poxlyZ0d3CujuwFgCklfLeKTtF8HIkuebV6EQbIEraflWFP3x0825MQIFIlpRSlf
qS/XDKUTzz8DExtJ6u0I3BgvWoC0roC2m0IjfzeYWz5DasMdiB4m/XiKVYL+T3NY
28HJoHQDrbT3uPBi+TJbevug/eGR/Sip2tARrJ/qA7PuprC4Uavau8lya1DMIoKm
CHXMdKo3fnAR2YZZ+9ib/z0ab2PnnU61C5r/TMwt6ezRMpQFhhAtKeuMYUTHnBvn
ZZyIdiqC6j3L+7XF7SCxClwuaD7NLUl/UvTJ1xSdMm43GXZbPcyV9LGVm5AbwN2d
b4MqS3W75EkCfopfpGtFVf2edyNm0zoOxL0Iv59gL4kyQw5wwiuElo/ojh5ZRpNF
QLiQl3A19Ann1JiclqsfjpvonKNEQ0b7pwXEJ1zVZAS6pPa5WC9PlqrEBlZTm2PL
qS0KkHQGme4vIv+fB8Dze/PYg+HlXDa/+r4/CJKUEcX1/4posRcoWDWHl7LJUi52
bZBz75QKXnGTK/Vo1MjDNx9yZZhsjefNil/PZ6BYIDnXjOX17RLL5qGtdvLobWGg
2B8S61vIGXOww+PM3UNhl4ciGvNfekSBjRn903DR8t3PINPFm7ctBf5uJEdEEcWq
N4oZqiYhL5ycnDA/3p6uUlRT0gUUFRj9ujejdNvnUlaLVu4NM6m2DkzSn/LyrABs
de7KIXtpq/SoC4tNyGl9oB47MR/fz7gglU9+OSdPDR74QX7h2YXZGG2Nned0A6eX
4lfbkRICahsFo5UgOYtzovQls8SEmzsoKmQyFtIWfNbD9N0LM+jzF7YQfqPcJrNK
+nSec0DP38HQVqKrWPSJu0wmGrqGDf6QCpn0JnmrY00RipwCGRu+8ys/CEOfohZ3
VoC3PKieapAodSHyRs1dDLsD+P+96fy9yrc4xv4UJIlRJ2syMJPQkODROPCczugd
EV8gUU6ZX3772+Qp1Rg4+yEMMUyJ4cL29dxYPcvlbijdgvVcCVUciGraJkAK7BwW
aTKzReShvlBSY02+WoisK3s87OuXRVLH29SHU35jSVaBYYdwyLljPDqHuodMGFgp
afWCfYBpWVAMGGd5YzsKPgVhObdQu6Q/zorDRyTWqSZVbrvTxrUHkdb9tKOF1EvP
KzEld1oatjUUIyXyJtNmRT0wHwfGC82XN0zeklyXjc0YxY7/CquO7/NpEIiYVf0s
a35MlTxa/6YkPg8f026rK5lec0GdIFDaMmG539aOfhFdky84TmeHHE2G+Uewq82e
+oEUtqYoA/uQpIZlbWL1APxWCqHvDWRnILc4/8ZUuRCgJy2T1DVPR1um7GENb7Em
7YykCRnEi7C1T2SNcBH4yY57bpPVIV8v9eqChURQbf6MZ3E7MYya/6D1xBt8I3zg
uH9/JoII6TtSebALQbdJBRglFE/igWORpowUSdslto+jmptyHvFg20+VpCPysVuY
N9k3H5IvBgCOlGkdYxbrqi/KkBHEkG7Agr5j9ynDssVvXCfICapbtqrNL55AadwN
cIWzn8VgvBJ1JblN89qGSJ4d4YlBeFeDONoGi8Ump1YyGiGa4k1cTYPVUhWRk4ue
tZekSLPgBixWcb4Dsn/OHxFxuJ2t+vsbSXI0v5yPImR7bi1Y1yYY0N3CUDItlZmX
xIGZx52+ajcraXPH3AoFLH6jT4ZvRSrGihcdlcL8meIyv3ZY2qTAoCQ2DFkj0Evq
VabX6rWpM3AsOiGbdGc357YYTUoBoC+Dueq/sWNRxjBA9NR93G8WhbZtxH6Zi3nu
B5u0TTfOWA+MoHkXIQ0OM6d69aXCIU/cKmOAKq3AXdvpr0+q5xbcCM1tbUGWA775
h7/ytIE7gcwswaUa8Lq1yCT9iDgPKV25VduMS79odhA4qsU9WjQUzSBDAxs3Eoc7
8nbUas/RpE8NosRGnyk9c36V785GSQoAUG13mmvxVC1Gt8wIxwQKXULndz+vkXPr
8ECOdG72ZpcQsLW802Jzr7vR09F1VNgB3LF9RHZShpQIu5VxabK0Qybz/QVh7ik5
MaDbl4IrK8z5pnHfQE4nTVLo2rqnoPDcJGkaRyRxHDlFSCmBE4mwUSp+4b1FPa73
oxXwqZcDU/4OmpsHjULTagLcHvwb860KPt0gDQO3K803f1QozDqLCyVnjwW50a2x
HUBf2K/mNWuTYR6o+B8Ee5J9Y38x6q2ghLPFsDPOY3jDv1T4NzJJZGVZ7pMqb5FD
D0cYtC2HAfuGvYPbygleCpFrFmkzLrZxPu63WZD5zbzsYScYReMfR1uOxtuQsdZz
kxEllfRwhGRG4votkBguzbhNeBnDFFsy8yrKsNBjIkHRK7wfQ4hIrjskVJELQdUc
mSd7YncE7uQ2vCmfNVvNPyjUfBWc2WRKQ65OFoDKbZq1xxLviZ+XRG1yZIpCMw0K
BtGCQrJLnSsvYhGXzEjAtsQhsYXkiixpSyHG2zxnaadhjGZwGTlNDSZbdyXBU+UF
wXOTxn0WEceJpXr3/gk3WEK0WaeAmx3E+remlzCf/c5vVQJh9m4No7aSerJIk0oD
YD0S70xg4+ddbI2dKnkk7zsAaSAoazYW4dtaSYNaU+1lWfPi/Dktc6h2ivAmaHv2
P59KBogVl2KpGMkcWA99pLc9Wh+uU4xQIOfrtbm6AHu8w+hXVP50CAKfrAHtg+Ja
TTvltX6rtjrTuwarn/OiRchb/DNsaHs55Y3PPOi8adc2/k4cmZTLzpj0WDNcVCUl
cpUPKRPjEjGRkCO1q7q/VTt6obeQgVbvw8gvvmVDXPJm//RfUfYfgSJW8cVNIJGq
Sm054HVMw+JQVC+Huv8g5eZiWwUvYWS9HVaBtz+/snzn2c2vLid9tHTh3IZ335jO
mVERrhF+IcUblp1EtJJqwBHdrEqcFibjoug7kpKvLvE6MPEe6q9PZnIH+NL44yhp
jxdDJE/uisLUMAxb9lmzRPDR0QSnaQFRBiSduwx9sNnZ90myJIopz2+GEA4bwTdK
rfzSTS2Kv7+VmtU6yakodFIw/5FaUt/fRS7j9CXH8DHBnr5Yr0rE0lj/MULoDawj
3qpqKhIgxV/q+mPTs1mbO+Q8BUKTU5Z18ZUf1MCx+hN/1AzKv4ZMmuXI9cIprvTS
xFVJEYPX9bo5KfXA7mX0/RRVsRuxvgXoba6YiLi0zS0qMWp/2cpLiNHF9Jr2cLlm
qw1mOZB9Zv5j009AYEM0/0yk8y+BB6qn/mGptg2ciIf5U2ZHALuMldc3Qi7A1HTY
tvL/wm4EibV2qUvAU4L/qbVoKUsXJyiSUH/XoeRi+UnjCfOXaCu7WWgY94aq1R+0
y2fbXqviWX/UGCaNyz+6y7Ht75k9YUig2VEejeJ7cDs/B1QmFDKQNfMr6pKOQToT
4sP8be2bNcBfyS/MrbEBM9J55jvap704qcpp+oFrP1OYw0qxnfKEVogvMKMlw0oJ
5obvaPFWCq6C355wURcMYo7L6HMUKL2v1cJgDUH9+hlGTgBjI6ueOfeurjDahwKT
Sg5ybq0i43QK5vG42yh03vMVhyElyIs6bNCmgkL1JcEeHP9kpYfeUvteGA6bDkaO
fQZ5vHH5Au4bQS5Ry9UhIKKKellfldTiMhlNzVcSw4f/LX6fwOdbqes5GW+JpIsn
SDKfi35njLVzWDIeltkTUuhien6kiNdqP4GWh7OSv6gyYMTed1GHdXe08MEW6sue
CYkpPSz7N7KpGMYYYwy9BzgwypE4k3wxVP/wyEngQjcvxWsJdjTdKf5TIWvU6/M0
8mJV8+UBjh+MDrgb3Ow4EaMbmZvymRz3YQSd56v06566epEBVLrx6CCfnuNEX7Ae
Lh7Fx9wLAbQ8Aylbm/j9YUPb3uwe4nDA5xYbeYV8RDZ+zVcsVgcWuzsa9bH80Spk
VdDGSV+7d+y1IIRpIHWpOi+tciolNphbY+u36d1aUmQDYf07r8w1yfQucLPmBD27
RWz5Nq80/yG4Jk80HzCDZrkpS96PFPbP71IBmrkIl2W3V92Rf3dLP7HbwIuZjjpD
3q6WMK1JUKzi/vvFilDZOZbTIeF6gcx9KJ+EgHX8P5GcvRNAGwfY4Tlle6gCfvPq
7K/h2bcnCVO+wLE90euNeCZMls/dRO36TO+0KCoIfQwE1xaRuC4GcK06ja65Qy4R
PIgPb1aZFJ2+oJksm/UM8GmPxklPxVMKQq/Ps1sb4rkw1/WrnQa+nr+WBgUaa8rX
tie7Ge35JQYw8NXYaU4ljPIfUl6OigJ924jjTJ3z1QDO8SO/I1bvjQtBj/o3ysbs
2DjBuTxDctsi8X9p6gujf/V4PMGUKOden3HS7L5+/r5nb7WI+AEVZU+tshsVgXcm
NeQbAPE1C7YrfW/xdGtkHCyM0AimyXkrfghuf8y0f3pBc+jUCv+aYpgMZcaLdC2T
ZFX/tSejfGAaToLPHGaaq2C7f3WZLDyRAD60Yd+3g17AkIesKxZojhguTcLX1OqG
Fim/Rx5uFvkAeZqDO7/9G/uOldT5aqijzkgemFeUP7DXe6THLMz3Oi8FXE4C2bGw
qhlR4FijUwwVLAv2iDupL2L3I24rQoRdo3pILBntWmjO+WTpiWNt5O4EvMmuySEN
9PrFQO/XUNlDLTI3TyZTAohzmDIPNkSU9fMDNXNJzEVRvqFKkC1oBtWHYY5m0Ajt
bVO3ec0ShX0428YOLti9cn0eOsNz75hDHsv2xfHFY34XlwqVdu6rxNu91IAY7NEw
L1b3wP21uZhRVq/0QrqZzmRyl8wZ49IKQVFLrbOdWdzgWd5sZ8RYSfhL2zWyJkor
rHunAjgDnwtUz4eej+YqhD/jEYISI/Gh/VVj1Uji9pE7KkXYwGRVF/15RreJJeWu
1zRg1Unq7Kq0QG4GdCPALyPTugj+T2iGeSVrOZo01/OHS/ZhoJjBp6+r4PjuZCcZ
gxz8poXNT+Qs9CyW5A5oLoS+gel3msGUKxjHmCUKQOLMWXsSc8ABuoD1mQQYIaWy
/Y19BohjJ1oNmLDt3ciSEdhtp9naAndbDywH24oI03442C1Bu3RL7+8uNWVeQQtl
smTo64nMAbl50k8Rx0HALVDP+pP7YpXBhDdkdujzV0E0FUhtA6FqGj8gXfGeCn87
26v7JkUrdHYgonIgiNDaaD3Ovk3e4ou1FSrRvJAs5UyzJJYC1/yW+5ZOMEIGbGFa
y/NqHbryV3Rco1gA/SH5pUPQPVzvKJLsAvVjJoWAYM3bIu+EJjFJ2ZPic5sQzMRL
0ASCMk4vJ1dNEcsOnH7fl8B2Hyen10lJSqfjz1Z0x0xmQZ+Q0X8a2uKtwjMpx9+H
5ADO++K2SCYw0bhOFLv8ETfU55rMbhSEHqsIbRnAP1b58009LZd+jh7XVPeOuFYB
U6d1rjaP67LdMtv7gVsfGkhUy7GMfkuacMwC5HASDSFZLRX0SrTprn++GrYR4PIH
XgpFoGTykEO5FUmcFnh72OR0RoUqQgAzmcuw6JGlfOu4cLs3nxKo+flyYkofN3bh
i8Zl1JHQxth9OH9tMC+U63eEQ829KIXVpS6yKyGiwvAtDVCwvsrvjNLSHX1OOfwU
TECamRBfLfejERVoYwenRZvYsAkxfEmcUhZH8INxGpEk95F+eiUruZ+Dlk5hr8ub
91fzhzE9YlHQ38yk7fbQuL1YRDxM/IpH9tE57Gu47LaW+moNsuCYF+NxcJQ0Qk3K
XFG+kEJ1TtqeD0xz+d9caqZPe3syqZW+Cx5n09RxAim2QBjZwRdAtBBpF7sPZpu8
Ct2B1Y6zXA0+MnAb46wQT/NCtdbIPcFaaIDKmjwq46kYkLS8c58nblZK+P7QNeRy
A2n6nYETVn9SpPEGKKE3oULxk9ZO8x7nfE6EJUUQTm+sno8rjM5zf/kK3Bebv64d
gaGrHASthOWyjUt4EIGMWSjyNHCvUQ1SA6+1yQXTeXxSQvhPjNmMPaagyCigjDBG
Icq63ioU6f2pznF1Yj89b2LZm0AFTv8bV5qApzv/wGgzeP3vZ/MdqQcajteeidIU
ahrRP4FPf6GW/oMNKfzmG/X2MkMB/jj0McwG3ypIkpvchkLcgJdfDHJdojabLbfQ
8YBwizLloNoSJvx80I/ReQyl9jDWCfe/rp2/lmhBkwCO0K3pRB4Cn8fpkOAbPGIB
WPZpiznJo0LMRzi9lbHPMFMiQN4yT3LEJt3jspNvQR4X437/u/4YFydLZCCf278A
+x0+zs6lqZbN8MghsbjViENma6DH+LKzQdDccnLVwgp9SJ2euen+pKb0gr3m6085
DhM+DJ73DzFVZuePzj2/Eqpj10622zXk9V77xpEw5xLx2eAT7WjbXLLjwqUktVBa
04QVQ3c6vBdVTKpUEjSg4xAPz4/1lHVyeMB21RN6pSRvNL81dUCucTJaPMUezo4v
mR4WIfzWI9Y+g/71BFomrFwmVU0qHnCh1dykVkNEf8N14nlE7r9AlhyltqlvJVdV
+mJXcVwYelxjZaZ3zSmLCIWIWX871qSZ1oQW8WodfLgKadt5vPiLe1VXZ3E3RAsL
znrTyUL+eiy0QwDsqaL+SPRFXmZsVI7gpuSZkuPcS6TFcGBxK5+xVWPpsLfY6LCk
MSlmkhqDIEjwInztbBBW1/ahlohx1N3EFxrXk/PvxEPJqkZxrYE+lad9tsikqbmu
mpCZR+nxd2DkbceUQikuI4pTNaiTuFQvErPlqp15+Q9dgJ/D+CQFJlT+lvy8f9Pt
mJQNK2EnEkq7QQCU2lw6icLiYo6Eead66ze4XD2uN5NyUZ4lAhrEPZ8Q41hcoQQQ
yhMNc5jamIkeiWrCCRpxsV6UrWwdmWvpmrU+Yf67OEVe9OuNL6Thrs5gBVuSoQ9/
AEwLgX7LlZKUhxzoHPFrO7Hvh3PFzpb9Qswg+2/zUOrnZLpOR5kaphlGhHvWhJyL
YV6e9Uy9OirIAfUylfqMAf5jFl2yVTdKO8baE/POQlBb+Q4yMSUAgVRLIDhiDqM5
SwPSSC7Pj/dGj8fiTRl3cPpDqbtAjabeF9oUY1ZorCQlXaO3ejT3zaVV1sgTO1TT
1bWFQuq7fcQxvfrQBS/X7XZjxdAqK9oR4GxQ+d/oQjGzzcajQi1+wL/6edUi7K1M
77m9RmL/fA2yYhR4E+13s6xs8u903SbkYYHeaIlFSjpTTh+ZAz1bDM1btlXGQ8Tz
rgI6OQFoG/fsBB4ad6WRnGzMAXhwBcy+GnkcOedIcbdXMJMbhtvoZt8Oc27cG3xc
LtheK9TCqaK7oESkYWjEa5tIzGARUmpmdkp3LpewG2hu2TgGD+5TCYYkQ86dhREk
bBsA5192oYxxO8W9MJ0F5g2WdGPb/N/4fkMy2xGkcl388gFcCdDV6HRwCYVMONMn
5CwnZewc+zyOasnp0fkJiqtK1fnVqnh49ubxvIU5S9Q4ljND4gfnBsSyKQIMi1SY
1jSVd0Gw48qY2/sDBNlgHGYUjHgr98QMafah+O+NsryvXqlVVdG0i4a6CHih4Hfg
Zu6VkGgMrHliVbEiVPHOO6FS6DYpoHUaxdguXTLcM17XwuGlkQ6elu08m3O2xjkJ
rh3PQA/qnAp/UPWnSDVAm6yhfPTXCqD0eSWSqWKE8Em+q+k4Crw1Iau6GVgnVtSv
IAUoj9wiyB7rW8eaDIuK3lSiCQ39/YjK3BNvbYRTXCQ1a0Ir9KOMXy3CuwKrovwz
IM0WrOc+mNHANZzQ5SGG+464eJdRNe27UHLmLAu8jwhgqJv10yjj56ypvIGfACaz
a3tF6DVCk34o3ISOX7Idbggq0ImwfJCAiE7fOnbXxT1cFRi6B+iYo3d3vDcJVknX
oVElv6TLJPVHHMSxJ31cdAuzG2pMgfQbCgeB9xMyNybjmx2fkkTJNhUESe9gjpq9
kLhOx70c0S0ebTyBUJcSYa1li+urI03OJF1rTSNG/e4yHYlWUIQxR1q5hA9KFaqX
0X3MrX8tA6b+xY4rn6SiXtNv+/LQHTAoZP9o2C3ZKHCHfhW+7uVLjoCi357zKj+Q
2oEZapxogEZH9v0zdThdCuCS7DgjZwRto1sJNddDq9w2PYfK0CjW4Vv3YrOVlkiI
wqD0BxyMKEGQmMTrvjKDMC6zxp3L7+H8Rji0vwwyR/AxcSprnBjrpLyzMvn5rUeP
+zBcr4BR0PiIzB0+kab3qd80PAgEcj+moj1fnqXI5TxX6WZA3Ft36KfnkpnSzPFg
5gCApqVZk0oNneguv0tWXuu0eajH1KdKNbCBnh3IdMxgsAqrXNIM0R+pyWZQFJFh
SOOh/CxJgMr5yCqJVFlOlk4PxiTuRHHIlhth6qCZSvZEB/8fTuV4nt9pLlW2WW2f
6wL+Fy57IeMgWqc33vccMWbOxnpyoI66eWw6uYBOz4MPF8R36OxufLU69HxnY+Jy
P2t04Jafl4t+rOZX5nyv34zk8Lhbmy0RNZEymBHpbW1z99FV2MOmOKWuXpQHdi/Y
vpU1NKuBb0n1zf+kGOk6Dw9JWg4TX1yTUrsDXDB2rX9KAETbsoHuyLmaKqnNkvZB
MWtGhSXc+46kh0YtlMCgWyuL5ofd2OcHAY34UP032/85vwN6IylYYvrPIF1ZPPjZ
VCjSemEAYRU7nsdPxdG9urvwJzG/y3QIaHELNULP3PfBFC7j4WOdyOeRXWnjzGag
1dxw+dzBXuilrTxexgxHM1QfRESmrXcQaL6I9UOtowOVm9jBGBuAsDvK2H3FgMci
boIXhz8AUYemqhaiZ4sas1ODPp3B8he+I1fl2Ls3krtjIVlvX7lCMDZmJfsnbRyu
K93UxP1xtwuSr+5VCeMsCjG8MzvWv+RtsWenG6WFGTWHqTjTUZDDKCI6nGGuS5ks
x++47k89mZ58VQDtABKj5AmWnmQfIRn0l31haDTs66xncjm/VoqN6/3T+ydj06le
7SlllH/OlG7vIM1Dbymu/3IjyKPOMYZSDyU9Y7zNJdeglHN5nTtryzTXWsok68LM
v29GYzM4yRbfEk5e1/h4TGG2jBsCErmCJz52JTa7I4wsMjQ5rqx1tcmfI43bj8tE
hZj1vDD98Gbga1YAg5vcObRgmBzJZCm+B97LBwGANZY+Y8EfXQtWt8Fv/6yti8DF
uf6j3KHxkcbbjBSgJXJ4ZlKWdMHIFAKGWIAH5WVbnkp8CSSklnIBFC7UdaGPDRAy
nadU530YuK6CL5l89O0hoC4xh9LyaxKsvVrZblUfgIvnjFdKixu3p+bn8Jmv5NIP
fkQB/CBouww2eNDZTCE/wM6NaF9kvhhv9NVaGVbo+iFICc23sMhBUcgz32aAmc2M
zzGRCOfZmOrjA8Z2mGOLxfqDbUPMXTkU9N0mpmWxP0blh3niOhI9Yw8HFiCv0KfV
hOBndHZLtzu6gzDI2Fg6KHDjWrV2bzAhTujjuolHR055ddkMvPnR/pH6NaA+aTIm
ccmU1AMJIX9x9no7YDRIApVV8+IWZbJlW0+o5mWf5wOchnTkp7ZUqxaxoJcgUrIh
ShFL6YA8hIvNQqjOR0Oc3CZ13EouFkw1iCjdU4wOy2HQJtlDuG1UtJy02MsTye+B
TBsCUpzUkmJ9t6Km9A9Xy1FOPssITFow6jW69YAU4+4+I5/mV05+xXRT9AJ6TLu3
AEtPYzmPj1Tbj5KyJlQqylI0gpmlD2m1mk4IiYO41+xuA6AEKodNoVnM0losbkZF
l7EnHuNOZ8BX9fQaVi/L7vvQZjRSB1ZanpdXlIYgbFG0BlmKtiysza4X+lumHAKY
8N/bDdUIPM3cDzgrem2OXCz3zKWYTroDa9eroK9C2m5Q2BAC0Ssl3lt2bxFXhQ76
KbAIZHTYI7LBa0s64ykzTYH6QH47m+NQ9EfRkp6XqQQr07r6a2/RCE7Uiz9TFc+b
lAFkGs17HqISJ9BAZ+Yd5L0WWlVp2QW0xIJ1jhqHJsDA6Cjy03MoTPLbLCeo+DDw
kb9UNyFxJbLJisOQknRNUQh21TRNfZgH0ktHVZbPhkeFSwKiBdF4PTjlw7gmgNFJ
slb+D9MyZxcF6mwslD9RGIBTbBHnCbjkOaAlsVR9gQTCf5SpEX+rSvnVVvjS2Fp3
fKlmfSNDCWQZjgQq2xGKv8T6HmXynmozR/IK4jisBkTOEIimdKHR9FfDQB6tiXPZ
i+ufUCXCCKRVR3MX4fOEFRpBTLuqcDWy7aQ7E4rzAIv9qXjGk0jAUIB+AVQMN7jw
AXl7uyxtulrK2C3x6GLWI+PTYVDF8I2oIGl6pcStXBHS/nhEFuhjxdDnnuTsvKyj
EdXW7NkAUAOQaWgTx+z6Szr0S11EiMPSfszdZjYw7NiB2MKlZ0jvigBos6ygGngc
IUmTKat6S+zCqRzMrngBV+YhRqObspxBdnJFu3PhQ28G3gH1qUjklyvLdDC6c0SI
nyc2aTPf5ihC/Wgcparuc/flpqmzYrDWvrzrWGLWWG3K/z8R4AcOt4QZ5xWKmsiT
QpgfrijQ8637Ljx/nZhnIQrd4NLI3/10KMazHsmcHj7pWCbBwzJ0y7yCx6HvCmzv
e9WqEK2wJdeM2OQsoiJbSEg8Sv9GdgSofZe9gZvjWgvcb7QnytXtvzGDSNGZ+KA/
4Dgy5mOCyXOIJCr8HjDmym9PbL+J02ZrJxEd9RFtrIa0GZbNIaK9Yc3aD34NpXcv
tKQqArlZIvJGAAx+EGC4PqJ1c20JmkzZA3GV9woJcWgYnko7uBDDDrqZbUXL7T+4
tUJ+VzW7yFSs4xdY7ae/vkzJJ3kPijkS8fZyODY1d98wYQ6gTs6tIS7G9bGTrYN8
CQIyn2xnft/JG1cDif/I3DDOtniXPFGxxESy5Ox4z0E8P2dVyPi1d4nw8xODBEOB
eip2FXmNjKK2yx2BD9zZw7zTDoOXFa1j7NpliZnqiiOQfIvA1rHNcxwsKE2dUlOz
riG1XFQHHDqZRs8ILy7icrZ7LVZmH1J1698wva4kXSz7tGLeC1WOyw8pT1tO1qzg
hDZp2HJrUmsMJ/QIBb+0DbD1jFOVz4NMNKKMeJsDLrTHmfN8/PZAoakKUycyJ8CX
3bkWzK8B8JcXSIMXfyvzjArDuQvEwpHZXkh05J4/1FkkU9qSnva/14UMlBrKiej2
N6ED/Tc7pylbh8jeNIAbK6zaiSeRcsNXlh9q6EI4wrHakuyOkVniqiar103FGRQ2
+KX7BALc38NNH1FbN8wUhaGwHQN/mN1nCPIV/mSvIUSs14LJBoyP9aV9HhoRIU66
u6dW5//81qKU5tTsbdewRRyocrK2PErdWEn/ZVKGFe1qT5vKJzUsmOirS8vmayva
gkEb1AfADsDo1GgzT428vTxYKaIVl22A5VnlFbYT6ZNSvF/IKrRIEVyQuxajUB/E
PtXaBW7+MLhpMNVgXrrV9MkMRsDEilEfvErby0HlUW8y/HWCUPutQAzSqmnSW3Bf
mYOoMzllYa+nJZMDIeTq5HMlNjaMcivVztZw9ZAfACSd2alTXcUN2bJj40RxYw+N
HIyHAnuoLDjXTF/cP/KMYbpkYcSqoj/kPhW3y3G41zFAr1wwD6YGj4piiVdT00AZ
HsGMYLfOkVB/PsINnEBjT2z3ImVYnPEcrBa1/0VZxUUsE4J9Wpxcn4jJwUzyWnYT
7nuqIOrc5b5O81VPZLgiMWcKGi2cjuzHxke6RMoVQNL+VKPoGdC8a9XkIoB33+PY
ZqqVSIgpKifTyxfkjS4rhaWu7U1nhZKIXHBj8om5dFN3g0K9PkTxO3p/MdMz5QQT
Y+zCy4hGUjBDdasyzSwBXS5uSx6zm0jQh1ur+vpk6XG+eQEwWL3pL3zRKZraKE69
nRp/x18kNKrtq82jdllXxePUNhvTQn8PM1/5S9yuosJTO1BPR2W4jB1znFC/oYUl
7T6ujKP5OgG8p9LRiL9HS6wdDYmexAICSB5wcipGLc2qP6HM+iNSuScwAXZ/0zFI
g3xUXlkViEq2txuWBCzMiIo3asNsOD9y/b4+/xeCYoEAUuoGfQWsFviOecOpzs13
jS017ZCVPUvPOoFhsfrKO7gIBpJIrML5UZpcMORA1McziTsuHP5E/mYFbuejxEu7
EH9feX5CBIlLwkdf4Tu8S/+mUNvRUwk0Ff6XKxYw6Rt8aOBsS91xVenPnfs3jvsD
2cYxCYIwn0hiVticmyYBp66Yjj0L/GT67sjvhbHYOgo0B0Iplo0aEqV/O+tR94ui
oOhm9psktbgyaxVOrFIYyLVQ9fu6a46cbL3U7Tfa3wd3pcXfkhbMh2j7P6lnHygy
rq2MmtfTgqT+S6+Naoxu3SXzpHcNVbfGGanZwqnpmZrBbSoFaFpL9+kAy3oP4P12
YNJbQ2wzRuJiHHnLkj2hTQyGpmyQ7KYQHYNTwsPpNw8YbfCJkus+z9r9ZSTvi3E6
/ThjXpa0aq8+rTYTBPFk1CmI5JVYZIdT/kMNSj8DsTMS3f+aPaQ3YlY7xxjFzeYG
3PUka5jje41zzhLnB3s55JDzofgSAbRzPf5cwd2I+5uPvp7V0CSM8VYHaabX814n
XJ9/l1cD7nZkD1KgzxIVEzK2b2lbYOgnfM2hQ9dj7XiPDXxOYnYe/BFtMrX0bgV8
YwOtqdycfVjY//MehFhwsgwRn1q1v5AURPcB8cCZTw8AKRtS3dNnGbciS4QBicWK
NKi7VINRYPugeogYdEPbUYeGBcuBgj1W9mzZvIxpz4bxR74/kK7s/bjFIscFdR7S
ONqd+bIFrdTDjOSLfgTQvUpc8N2YqtGPRS3WGCud9QyoNykzI4JAlzBCJO859zZ8
pWLrMeogsx2zO1RmtxHBN7kwJOSn45oddh6Sou0KTh7i+na9PfEjH3CnWEFhHvJA
yyDzBDx7UHhX/BQaKV8CciJE8NN/AGfXzDWb9kcx6CqTiM0Ogt+bC96wHrmSWEpE
AW8S/AAnawpBW1xgDxqU6El4kYDsg2WkntiTNdUsjINVEGmd7NerTos0cXzY1BZS
0f0vBDM0nzjSv2oJ9sD2XZli5N4DHOkXoSCGfQb2ica3Zp8nCEKkQYJSi0ByS0PL
wA5rCPmFDoboB6tbQl9Eu5n4iv48/+iYX1sYMXrj9PokeDPo7VfU0gtkw/R5gIYM
y4JgwCscZutI1GorbWnBh2lMMzlWEo1pZ1fTrBZwWQN/0y7gmpbvqQdI0qJ20cfp
iZXbamXhguS8r0uLkcTNhOArXSaFQtV0I+MRu1Av6ebCJTjcDWhZqtCUe+5+FNoA
JQkV03Na4xQO9dhlZoQF3aUZA1zAmrpjiILMYIg4kQIvWE50aOWGIQkS70aXRX4E
KNKTP56jmYTusqZhVH9cYJ9FNRRlaFVGd3jwZCLycFUF/c3A4xkylqawia3RxTVn
k/W65QBxlJmKIhu4JURJsWq50oBK1oQ9Cjp2ZcSmVR/ADgkXetO5LIfphPmPdcQu
f9C2VqpxUxJY/qvUm0/xeNXle0eHvEUWGOuahU3OwTrvy0nrui4TZcnbveid6oaD
xvvbgDIoBuqIcqC/Iew9y7ODBcxfOsoqs13Pm1jA/XAQOcVASzXM98ypZlo9wQoF
dehLgrBnSR1UgmY36N8kqFfn+rBJ6q03YLonp1sqaNNViHi8Z7TI+0QSLywlX40q
uJvcCLeiQ+hb2LAS+HIL2IPWWf6oSeNszcGLpiL1OQDyOwH9tMwBf387oN/qehKw
QFiuVt4ONYE9hofQT7MOMKq7D3n6BriAwQnJLoOO/L6200aTNIYPFd46eqkuQqNg
ftBD1Db4NFQrTaUmhLi443FUZ6qh99CPO+FiR6kJB0C7yLiN6yIEMmPNMAzrtPBf
8lJZAcLug7W8SxYWeYDDn6bKaKGme16Zhglv78ehyhNk7E9R/ElAGbPCsgPjsefi
Ogz4TofLVqztU76fGs9Pt5aRSS95Ddfsq8uuF0TPRUS+cIc2Vr9Hnec/7duKhSLS
MV7sI9WCV3+1JFjeR4/mxPUhHsO1aS2GwR7rs5ZC/v3L/Vztz3doXY4n2Y6vLuY3
hxsutBNxEVNWHSNoA2uNkHBto4HCdVRP00N2HtDQAdHcVkKI9ppAjDDtqHAZ69An
p0dE/DS5QVqn01PTcQ2QKfjOm9wGRdHUptjujlC68NIBoxLapCJQXBZ8FWQ+66KB
GP0xunNdp5i60O7/AM8jDKVj1hL6reL0NrpQPXwurE2D/qzeDTiKOrkzCiEvxvFc
dWSIL3yfXSerRip9T6iBUgD7qcaF+kwRMTB3ogiIujDkujLCLmTNGFA0Vj3S0Myp
TlOj9aFoHs0AdFmHdEqZCQZgE3a+Kbe0p0sRNgh2KdUAIqWzQVVijLGUxlanrkf2
3F1hzMBGCLimt3uC/aKC9S4/m1hktE4j0imhLhRZz3bbWlV97cXzXM3060mQpecI
w7BIQooedsKX1L1LOJIJRXWelIIJmEBCDq2pxFrx1m4B2kpxE2CD4ku1h7RsvL20
lE564ZCXeiO5nYunTHx6EVNvnDNgpINcewDLcoMJdmzGhqYE/2+mg1wbn8rEVmbU
9mZEDIMSXAawCTJI0s3IFWBsf81S4GwNimDQb8Jboc8uX+EQxtu3IgK2+e4I0tHi
c0ZehHsk2wx61dvt5opceivhcoDt0DaVfNYK+kfM2RcuPxr8/1pZKxC+6nItkIku
L+Q65bkye++Ss6Be8Vi7dUaqT5BZXOkTOoC5QrYkWXf55ksdFRrW64xD5/Vxdt5M
zrs3ER+DH8bC/6e8qJflR3oNN4Ha1gKkptUND3dCl4+swojEQJyR192jN4TG4rEC
ftk8IZ55GUGfMQrpV1Bx9M8o/xYHcIft9944W9J2KZzB+IwD7PMmaoyHc6Cz+PoC
4R+hc0ojYabS4yJ/s5amv403z2xRF12W2Aw0VkIXTLbPikRJi1IlaA+R5NwoL/0I
sLU9f3x2NkRFA2CeP5VGwk+6qriYA1qP4uXKHHp448fiRbPaw4i0l1BGnidlOO7J
eWi4Q5qtEM+fKV5Yt8ePCj0JXjaWeZIj/HLajOhNtHy0uGTTBKaYS/HjTrrwqsZk
P1UYf/q7jsum7D5RAP5/uIjcfeNVZ6/TYTP1X1vZdlY4JThpgp56guPX6k2mPasQ
brsB3QZKs/NJURu3+PlsEqKw65MIxROrKHqmi74km3n/WGC0ROjjo1x6AifvnS8L
VsIS/4i56APa9kNXyCTD0HDaU9bRX9bg5xMffnE0QGBGOkPpEXvFw7uSp/bK632s
wdxdrjk9mn7u5ddjKSLjRZKZLRmDH833gX0U66ZpVwWicJbwH9dKG4BJOyIIl3R6
KJXUSXW27+GWN0X5Z43/IoKHd6YVDbOLj+LSfYlQ4szyh7Z2EyGb4mlLiTc54g9F
kPNPZmzIZG/90bbumSv3kq56qHn4LR98ruuCI6EFtocc27K4xlosfrUSlMIkGQbO
Uk5/uSt0hHEQhHIHLkwa5ouTjga9GMPjGwEoChuAn3sxaoHqWPIZi9vdehTpIpYa
OAr61CzrswvBkPohxKLc8kpw1ORcl9bl+dWfnJK0GuZdY2owbgT/w9M3xMxtSaOn
L1nhwiswXBNXAOhMd8dn/GefLLjqH5LLT+/yhslV8WQ9e/QCeVIFoD/kOGoclsgE
TXhBvC9rlA7PaQBgi8RnQL/ZsWzUm0SFfTjG/21sDqCn+tyUgn5eqDQ0uAVDI1Ib
g9C2PZW+wc6RV2Wy6X0zV5hmGdDdXpoMg0wxx+obmuR2A92q+PeOz/aAUsWAAAu9
cei8/9QVv41p7YPNVsuQevtXPtgpUE3QbRui6Bo/PCJFkD6i7THP2cA1ma4JmNW/
2vbfATBo+hdzPXdaT6GkSe3rAoACD89+8GaSBl8rnbhYbD6yUIkVHxaLOpQ2EH00
QLjvEOGDJrCARV/obV2agyk0/d97vk61z7tL97dz07tJQdNCHL9WOS5cwU1xMFBy
x/Ny8iqCMOVIZBB7yQXD6zGfRQb7f6iB2sUWnYdWlqQsYCfQfGOvSRxmLZEOMh2b
dpSpdARUlTL3Nfmr3lC8eZmZcXHgzifh3qyoujyrFwfDGmp4Cp82lcRCAlTrthDa
Z8iL1rc3vnVNfHyXrA6J2ERhLUs+mP8MT8Fk8VZxGzOudskVoGIaqeOY6nRxrn1q
9SBD/Mw5wXefXJJUZD24HMQL6B5LG27tiZc/YmO8XTE8Lhhcodx8XJOhq8fM7aZ1
Qtk62GWfcGbTMglpxHyuUdcCvqcyYU3uiCoeh14bKOh8U9cQiXWNpv1iUqC8PEgL
CxgrmjHt6Fia9361k5kyxeb4MnK47VG+uhE4DC4elXk0Tjc/Ldz9yT74LmKT7Xpe
1zxmzX/d3scREs4Vjgh6fHmDu5ytXDLQDtHMWqUR9vXXj5pVXLJoPer2iYiqI6y6
JeiotTmGPhWofJPRu51Ew26S1bPeWG/lrPK5NKvrQiYxdUttJsT9exICQnIDPFx0
0fYFyRiV35I8Awodd1NEU5BUzPjvqOeUu5jSY/QOqk6ySIqHnhsgr3ywNngfHr2N
XaNR+j4dTgMmrd+4CzQBUnFavUpgAuT2TGlkYD00LfcgjJDtR7EQywwKw/PihJnU
vaBim2cljgudk71xp4CJaQ9xFuA4bED/n1RVkP+NgGQ+dJaJHLaMOi+C0fOeq3iB
JeFQ8j4kTiAUfBMJj+xHx5baxM0cHP4ZNT39aJALKHMzwSNoyXoo8CsD2/KlksUQ
oBNwibqT9rk0QsZ0fBmxx1r39opP+ampqcH+wPD0Hm65rVNO+CaxxYRvO+T9kDhP
A7zzHxi3KjmUKKv3HzWlTGr5EdiKhD2LGsZubkcQUh/kBq8bDRlABvP+PSbbXwgS
Hu+8F9r7vxA5FzfmWEY5U6g4np1rM/7paMGpobCghgACNC+XG1KY7KqZeT4G112M
y18Mn7/laodMLCwkVdvFX9NOKqLtMHBF898OyWDExFBgTLmtDnQszR7jRdUb5PIE
fRdNlhulLyBt0ePXWheU+utau2QtjrHS1rpGVnbtCGgHj6Y2qCQzoy1JI/kV+dCr
c5+Ta3ukouWFDivuiybIFUS/fr2hyPkIy2NJz0jSjtGOeduGLehruymWcCzNitNz
zR6aXZD6oBCA7lYczcZQ9vfwXW0i3qfN/55n9KF4rqed08vgv43qfKatoNH7VKAH
p02Grnt/MPJzrQotqFBGT8wuRTYxvkjfJaNlvnmBCoSm/pEbrdtmuWk9v8gYvifH
MaU4TyI84XEkMERzNxINFFhptYY/lV42XhDjhJZCE6ClZtRHJahynHONDJqE1xJ+
nJANu7nVMtT0Hyq9giDLeLUAiS/7ZlYk2aLeA9P6hRvQgUrDA6ufpi1W7EOn3x8E
kk2TjlSvegABgGG8elmxeBQLjj/KbbfiMREpw3NePk8yorMPC5CelsrKyqmnPcB+
7wyIcUhm/CRQPZ5axsK6QjGp7nPuRMt0sAKZvITYx23YtVJQlRdM88zxwETXiVb0
qZXcKCn4V0nFocKKuy/sjzbhwJOIQYfwqY5RFdtrJOuNGajjqz/09nKwOfniGX2t
k4r7GSaTYvp9wSlVb5BCJWzvDsnjtDDsTW4UIYJLa7OZq86txmZDgbgtKu1OV6cE
RkK+ilxxhC1coCix++RqHqS9BmcBJCbuJk+3hvMeECDEF2iFyIQnejEwWriwPnUU
BxcEslq+ObnthIVvtgfERDsn5+ZHDOwI775pwCFiF2InI/AI/7XVWSNeUOF2GjiZ
mROoR2FrFha8mazj2h2tvSh57T3wmvvNhd2idl2a2CSGwycnIlBIj9MZT91z9e9i
0dcv250xUHux6utEhK/SdWN18Q82k350BbK8gvHaP4WABaJaBE11giou7Ew6eKDZ
bzPgt1quQtqF68PlnDMu+NdofOkFj5C0DkhtdYw/MKQGrbuG8SP1xwrVTMLjgAzN
Sh6z38KYt06QO6YDEkiu2pMg2UaeCUfEFzIJlSWYRjDmWtcNdFk+vqVcZz0Xzyzr
ekLHFLrUAvGrc5SkWx50gkEX/XVprSJgNf2U574JW7jxYZ7IZF2fJP8uXtIVlGoc
ToH9C6aSt1bTD3h0pDRvwNI765KfB7WKxAqCrpjUnIqlmHvr3Rlh66OFRh/MfBep
uRgMx8+UWf8fHUVIA3LPamZxkdu6KmfyWxaKdYVktMTn5GObWHpux4Gv3hspXIvO
4RqOwULlmll1rVW5h3Y0K860pGX5Y44WdhfoJ8UA1KKLr/B7l2mAyV6NuUMBcNFB
vVKmVDEnt3x7b3F8fHzCi4g+cAQfcz/GXXHJxUYiKHrNUs2w38dO0h/KePeu7v4L
djPbs0u+f4CjoZTxMV9yBf348r13lmf5B73ObrZg/E7yCn8AgMBzpjyJlXbep9TH
6X+S5E5ZrcbANvHHuPNZGG0b0FannSyqPThHN2QMw5d45npTCjveAIfx0zo1eWEz
ypKpw+A6ws039d+L37iMZCFph4oYFyYEjOMULK6nxDMEnw4oPQNmy9l5sVAJi77N
H0RLKz+65IfR/xhpGMcgYaIDiEa/FaM6lybUhC3uD0WItY1b30tURM7RqBDVmxAv
r1cphXUTWE+14z0r37Zm/Xn98TD5jo15hVMNsSsnIQihurBOd5wCYSt7ubxJtXdU
isEbugSY2W5VLQyfAn5yZaeFxZIjhhGdEV46R3QOKRR6UgsCLyiAh9GM/y/Tx+CM
qjP2PYqQ70TMgeZaOuOIUDxk/5mikzcS0SvgAB9dPZ5mHSRiSxihrgwmmZvGmtJy
sxT1/aXavjlTCPBmHi9y9ZAuYTzQfh7VAUAF+BGKpHuETde9QVgFLRCyMCs1Whgu
4c3I7RkpFCPMYz4BbgV7jbwavTqpjiREY3jXiuHBC+UL8aGKfrHEIjACUQUgWXCC
lJHt4msUMaBCJlcgY1VLOWkA1bUt0z27Weeq/NYaQMhYRpPMPKjm5XxWTGxFGLLA
uIk9CcdZMCJZM4HPMGwkYgk1u3OYe9QOLZZwSDVpawJUnWWVAUow1UMIj8MJfSIm
9GRrYub9RA5najayYPc5dZ7sQDU2ocLqI9dPkLmiqbRWdk56/yYinAbSmfIFsAcd
iLNQsT58TIQoODn3oTIF4fx5kwue5pfpXsRyJUbAOO4zNDUj2C6xE2b7M+YvOzUC
xkuErScAaVzzy7zI7n8pPqkHKLUDHyBB9C/jRwejodWQM32RPOZsCmCGTaAhis7e
g/1gO8gINjMzI/RmlSxQE3IFfrerDE9MnLQhau9xtcIDkX1puqzL5HF9rIDBW0l6
kF6hhCyTzVBBvPD/NHYG6N3aH1WBz9VUpdo2cqLJEdfS+QC+BcIF4xfzmy3Ezm06
xnDSJQaS6ke0ctR4EM8Sru0ng4GSp1c205ZPUojN7N4OCqdaUxE33nspuur3dcG+
5RPyjBfqc1amn1tmtN+o8c/sAmZe0H0nvwzDNWxiv1ZNSivE1t2HDktUyfOSvV7F
E06qzXMuhskVGjGZa+esv6xEirEVE0LGcJzsm0wzQwfjj3XyJQvgYMbYT+z7Cpzp
G/PVUirF+7o2eBtcmBku9/XRynjHABQUpUqka4j+KEjdvBV9yuSGZ8BrzG7JdZ6S
AnkPiFKOofWn8GEkwA+zjRSJb6Fi3y3RTQDiCklUQudHfLMcooJ1YezSxi+d9HtB
IFZfc55f9Q+Gs91qpn7l2p7kKq6qtYQd9RO0RM0zxVv1HGe7W+1xtl4Ypd5iMPXm
J1W9iQu/McdUO/KSS2uRQy4pIiDlI6pEgO5ItZCB3d7ahNu9PvlIbFlZeh6e6ZS/
/2h5oPp1sT84BLUZQ7QhFgmTEGAqlBwEcPzobdhoT1WX/ncr8EFlmqKei9aegrPA
ilm+MKqdZLcXf9nDiNJbpJ0H2QIz4oG3GtyoCDGcOs4crWcPXMO/wTL+bUkf1swn
V0fnntn6J/e5hOUNuk9tv92wrYu0fvbc0yuTOzFBqqKuqPc0hdv+hUJELj+NtTDZ
aXQYOYi58hABduv2eF/r2kUiNpUdy0iJAO6o66GYhNwF6t7YtMS7wgYF0YmpFoRs
Hwna9Jgb/sJL9unrnI8DTUpmo5himIxVAxcs0yisHm3jkwVeJuKZk6xOZgnagnRb
051Gq+Ew56eVSe8APbpKMOPjG5Rh81ga4i8jGtuzc0h71f802lCBgnnqgGpJVBDf
Zy73fdbNeVs/vGdw37bCjoRsnaksviWT1COWayein/0Efm9mUHKYzIJ07hiyN6ow
WU9ba9ZuL/SXFsLVC1aP2iKK/T4rkv7ELeQvjcpJNwu7Bp3Wg6EkH8uLS+VN3no3
Iu0hA+p0JQGISA5ejIIti038p9d1Vo6eUD5cVS99k4LamdrODN+BPGn7rbCV2gt0
yqXE3T7J/cO9IDAIagJYZbvp3Lm6EZq6whh0VTOzrwsgmoHPQyc2+naFux+7099c
29g9FeqWs3rT05JzQPQAzh41E3cQ3A6kvwtpxtJQ5cQON37ydBHibAr8X92cQwEv
RKQkt1BQkOvzH0irJSkxJaxtwkhAMZD06540jUvSfNinZm2Ccs4y2P4ATN87FTfD
m0o3PBCVyWgcE3V30FvqsbQwyJTDP5bNdhTRDIojM8IsZA7QpEy/lHKgI0R1PrNC
8oTBAQ9DNlSMzTSqMLT5YvtzwrSvARPj1lTlNKsquD+GScukDCeWQrhWDR4+qljY
fyka0PZM47tyexT5HmqRP2TiPJ8mtkgCUtlHuVZQBF3iDAt2spakj9aWbIYmdwG/
r9059dS5pQzMb6fO0QMBZzuB6Zyi54G5esy2R3GexD/GxinB/UkebDDVyAgCcw36
YWSrdDc5/jyCn0UnNNtKkDkBEPpHplSxZlvwXFHcKAPWc0g8imP0/dzpDi+9btNo
WB39arC8wJYzoFZo8YZPqFKObh3K6Xpk8B/bHAtmnYn/aASkYAlE2gIAOfSTZOkh
mbVGvALxNpI7UF0nlygtyaKMly25CVDJBuy3nkgeVZQZB3oOHORqkX9YG/py3PPn
s00YWS5EDL4ySf8bca4KT5PQhW1lf7mLgRTcGQqgQpCx9Sa8fzBKg/ruq8rkOHm1
CmxqpL0K4m7S5eSs/LHUM72+xble9OLDtPZnJKBZ5QtduJ0pylRoIctsHK63R8x2
mqEL+eVM1rz9t5PtohXCMd9+8e2oWZ0Q2lWZV8+hLdUlP867f6TqiTI0VxEIyZoc
kD9r4/Oq6lLQjYj18U3HcVDigaSnBG37bYvxALrHwVs6y74n5LxnTFzcFJg5L2Xy
hlA5rSbS6WwUg/R8Cm/SoIYDAMfEuuJxy8R+ChsVIl6IpjuWpmpfnXbPS2m/njaF
3StYVQb3SDVlUbTDiIdhZNDZngAFCvn9nPl6cOSt4jS/lDhWvvgtOuFNnzGF3xRS
13FRqrdvypf5j7KmYLYwVxmqqw6uA+tVIELzIfBYOz7DMb76afCm0Rvwbz9wU5iQ
rzxcBKrf6aAGSsOXuoumxb3NpboxU6UBI2zh4g4BTNXyN04rupW28m2UptzMVzYe
SWcT0ZuD22s+yU7udd/cYXiOb7Z+QW6yd6uNBJHyuZwz+HUFqUQZPrlJy/HIHb+L
N3kB1ytshfuJnysrQUhFIhZXK0+t6boVbWse+RX8M5InceLrQ0QDOc5CzdwR9MG3
GvvXsVDFmjRNDEsNg/JMPie3s/CLjrJxpT18GU2450rUP1PMuedye2PoGnIGuhpn
azCivV6YMqqCs8c4B7Ufg1Ioi4GZGBma/KV6BrmtLHboc6d+pKBGNUBTF7A87zIv
mOgW5Daw2otaodHSCjwKalitOEp3O99xSte+pXEJuxfMyLlN1l/VrMFadP3riFBj
51q9PkBGiNQ7eviGnsxbNZ55kMHBJjrAul637AX/PiEZIBNxrIolpLlvyByotSha
zY+xiWIjG4AUuk7ZGPhsZ+bogqtDHa6sMl2BrUJXAKA/DaJKBzdOyimOa5gLf01C
LddszTuP3z7FQCwJF/l/1u9wsQIBr+xOwf+xiV6b+HHciDFTGDbdth3UUO7CiBzj
znQsFEsyxco+nzgWiJ8nbc8M36A5jb7doAWRTeRS1PzQnlt6m0V7HnOI3y8vECzH
dH7hGV3cN0YjswzVBFTTJO00eyemyDQNr/dnc79FXF3Nig0Tov3F4Qi9yq2xGHfw
yU+ibB4DdlMUPoA+isAKmqfAkz82gw6POMa29yviL/shXgghf16mUFA3w0ZtEj5Z
eOfAfOY8yPMvk21l5vrLaqnFHJT5daUO4AQP2bF+dAxhnZWc5/Xw4FTBb/x+n2bz
3o+KSOeSPuGqEIAfPL+2Hmjjttunci8IZ45HGpbqNK24s++z+ZMQ+8p3dQ0SKF2T
tKxGr34nqfF2ZPJ2pRZo/l5nJBc47zeSdlK1I33Gl0KU+yCvL30MdqUDW8McugN2
NeboHKRs6OgkqfjtZHhEaNV8az6gLXT8FNPTSTzIeyYHj2JsNB9wRlw+MNZQ5miX
OGoJRKRf8mp8P1pTgnlC8JKXa7H5PreH+qCzhvBtyfsMe+7vwzaFv6VSXbh/0YLA
iuTstDhvnbMe8qoz6xuWIZwTRufOW72CNNnNY8XW18uKel4k+YBf9wEZfwxh601v
e+FkN+G8h3hdNQ+URjM+DIfN11u+8AiZaQht/4+k6lCD1vrATNshccaD3pNhBMjZ
FiLRV3tZJmi966dko78N9xL3TVB8jY80J8KHTO+lw4aMCWLSKTdxNY7L2/UKG9si
uiMbdzrwgh4NQIpGCmvtwxxDoVsFSupqKX4dNiraRxKdafCozRjauqCbQmpbbhoL
no2vSy+pA4ZvDCelEjCZ+sT82M/R0O4qHR/6ZKsUymYyfAY2GTx2HKNGNy3Fm6ab
YI2LZ7oTNUP+RCKyVglH5Tc+acUYTF45mg7L2sbz3zdGj1CkRWB3bI4lTVICImZL
OaCNcEK7lEE5T4K7V5zqEpV+XxboxTmcsyq21EM+l5W8dkp225FiRZxV4zJYIhpf
QBTjXz4GZ3XO5+ear9KsJb3u+/yIyLI4S5DOhPROSOevlOPWzleGp9PvvMmLgE/3
RkgRghIOV6BXiRELgoNV6sFCnNM9HzFn9gfU/hmf2MNTMpWTdVSg+AuzjlTKjwrd
HoVbM7SiTasLoyZuxbuUJTdXnTLU0/ahRJOccbnblDCzNhC60fim5Z9dWYQGVa1p
YDhTII1MBWpMJSXGi6UwKgBI+yDPPP54Zh3bMf8sh733LG/Zz6F9E3V64kAjhKRH
5VdGagvXRdxviOwbCfCU6kK8Zng/puGAIbhGVCWI79uGb7h5hMHdPgMnaP8CYafC
+CqVgmPLfLP7yc7ykle3ZGHZdP6qi3FzYKQGtqJuY/lkUSQP38Vkx7+ZTQk3Go5I
f4vAYmUkPAuY1U+Zg5EzWhwivXhNgf1uo59VGifm8pD1IukkdS8n/VAZk7as+Xql
LL5lk6uJDeS6ZKHBqyd04ICqMOEwKlBFUovs9n+I00+ggmAiUHnu19Ky5Lq9lcvY
IHHqw88n1rCxV4cIr/AY/cFgZcT9Xkopm/zpJKwNNrhrtno/rPtC7NUE5bXGogs7
ZFztVJS5PoLWo76yQDEg4N084DipWivG8lZyAhWiyMoNJtKOdrDP0iLESnQjz3Qf
jiE1ZAn5BuiX6XNRquoNpDOaEt3Fmlh9LTZO444DfA9elPpWtId6Ff2uaijuT22E
PgELTdB18HupSKalrlvYtfp/p5vqIUfgCNtANth84o3p5L6zvOtOeAeVYD+5N1cx
SwM6bdES41Qjxo3PNHwrweCOKM6JFTMr4vPggaR4eLUlHQ9QY71Ve2WCWKCl0g0c
PRUf1YQtWwpRnSmUJTAdR6xNAHBTyuQe0qX44ZtdTQhrEuj0ZqNLjMNjUIGAhSH3
wTPtdbBKp+Vv4JuE2Rpnga2zfHyTPJrPOhJBKCF/MeYN5/mEQok43qgDjOG8hQUT
5vAk56jtoP6x8/71aORZtP364gd8vPhmYGOJTFKAPlpIelIPfjfSlWU0xbrQYg0C
lh4349OuOPR6ZBBseG0G2vDCssFaWS5aTgauGYRVedMl0Uvfd/2vxh7VnjXsHfs3
0jT+RC1buyspN0P45tL4NjcQP7W7P2+QOCVCyaNcDFHUOgJ0lDtodHdRuuNb/ZFK
d5NlQY7acdo3ekAq2Te/1KhSxtkBr7aX7inH1IdwUiRI/1Ucd4e4OkvYdhbJIjnY
wLdzCkgw5YIyIVw4TWPDJONB8YyCWUkPajSYXMHyvENwc0uf4V2qBLFqlwuh9bIo
G2ncJ5N8E3fVs3j27IUhUbOfGElgMXUsASOYBfCBn1gaRgA6aqufdlgAQYGePXOj
0kdsRs8+f3lDBo/krxZwRi4ZwSJheo2yYjIg5qOB9dMpKGSExoCbjZoG4gZZxt67
nIWrk4c39zFuuj92Eo/DkcK8rfxsEpfCewBOvEdcJNpTadhU7v406hFftA1IeoR1
1HZtebAUe4fCKu9lbJKGPgdAiIrDpT2JU5NzgILrQl1iTxpvlA1cE6mSzIYsb4ZQ
eC2GbunTeAXINfxuegRb4c8c5pjgVE3HR+n11wuPmLaKEbvQLImRVVftcrfxyf1E
lVW0ma35pMjDrucSkEDndA/Us2+xqW0SQ2WSVsQ+kwGEMbkppuXk5jDHNpNafK9g
+VFB+FP45cpiVJZpIVgq+z+9xBAIcW6ASW6BKbA8HzHV+7GI/qn8A33fNKkMKT5l
1S2AtLO23WWqdAfZTKZfPnn62c2f0rVTJM12aNur8Fas+9iSFYdIyTcSUPdMlM4i
uzNtFS8UUoFFn3/pnQHjCflAeKB6VyumjQklfwQVNQF9o91kdyW8ymDYnFUwIj46
7TGvnYdnq8QMbtylv8vBVWBcZ9w8BgE4/PTKFI0VGZuWtrJpWsxJI6Q1NT/mLXH0
0Gwrl4SJAg8vtKLL/ues+vyBMT9GcGr78KhuL6w1oP2DCTWmz8l0Ho/wALJXoQu3
BhmX2zwbOOPlf4hY1Vr351Hc9KCwajPyXo35937GkZu8BrR2plmWnF1tPHuVqVsV
Of0xhPMSQtbZM7BnovejcEl4cfrxmx7UxtLOWs62qxwHlADrl1pTDPvu9a4POfal
W6EjrQRCpUZSCQ+ASyINotOrUHayEcTPIY2w0rizqVm/dDnrN6iv1Id1qEeY9gz2
bRLWfqVI6xklhlKcRmJuEVKlj/jeyzj75lo9QTghyiFht7VnlbIy23+aRjYideal
7BMHm2l4DapYMs+Su6PUg2vHwPFulKIQ4NWO1TMeKJUChCGBlOWW79eojWLnmxHW
WXD6OKZ1sNRrRanWDeTLERLZchxZtQV8ZYWeqoTt48lhnWXxb+tMGQ69seisvLQl
DCSQqRYGDdiZ+okxIK78DGDkPFScz43LbYdKTHeTiPJrqbhhoLodFpq1XdPr1ZfC
8z+RzzgEniyUYLZBDo/PHfQSDXoBqL9HcdDlBZMYm6sqQOGmUEoGdyLjD84DkJs1
vRvNzTmROSaSjQH3qVN3Pb+X2OacWNIu4f+GK9gmAyPCgn17HlrfCnMR1DuwjDlr
8m/cq8n5Rulex3oukrLIv9pp2L+p188AIUu4dJAZnWkQeFvmF3yLcp3we4/R5VoX
9/Bub/g7s1t+wu3PvVY1kl3ER7nIJJghYJVTml6+vdvOTfc0AaTuwXPCsrWx7Kx7
B1iHaXQl3dj0JQ5ntgDAGS3DJS7vOeuPa9FElPFVzkbaYR9AJIR0AGJFocgFkF2J
gvvtmgfG2dnAsLmJIik/P6nftM1H9fH3dIhaJYQ9PCLzi6Hb2GOhSPIr9b91DcOP
7GaGth67RnmQHNlOzHSSMuohiogpvJ+if7DuRjrXhqovaSm9Rpd1QvNnmyxEghF+
jHmx8QfhXKIC/1oqyCrDxACUYb+2mfAHeGbwe5hxnGKamt1oPRD9CdxYxQ2XuFng
JmUNPhEK7iZUWrS5rO8H18r6DUKp2YKkfoJ1ezhZJwDPRy7Jvt9xqnafX5p3PgiP
T1pc08ct/TWcyXv503XeDeO3iL2KdDtVVGFXkT39HA9lPou4ADUpA96H8kWpez9w
P3oMMvWBemBE/WytE/lBsBWm/870RGxZm0bCAeCXZOO0/otUPCw4h4HRkQpRlWSq
YjVy/lvQJ/5JAENpaVE90CeYgUPO64GvxCXr757MdLXaMn7J5cF0JqTkHFJgR59P
w4nFtMnid5XJyhJ41N4adwht74jJE+qcpF2JtFN/WlIZMezfabdkEuL0Rnpjjl45
pkD5gSlUrx560iGZI8wYloXEnpF8KyqELjqvogb8xRrsk8l+ntQbpJoZhD8AO3gy
b2w3mew3Q+/DOzXtyC7nPe5MTpQcEIwGVIFV8+CYJRfHZ/iDeqjGAQj2Z5cj9VKl
FwhQ9yNAFtH2kD7tKBm/+enZxjUN/avwv93Z5dLD4dnvlc5mLG+UB7TVUtWVhUju
3w5AfJOd9CT5a8EBXkmkpNNLHooYfAIyFlp4dC09r4AnQWOuL4ltbJljy4EaLCOI
QyNdDjxMXode2wcL3hrI2alIIUu9vuhfxgCX0DBM6FUbL/VVA4Wd2RlN1y5+5ShF
xmyhUztHcN3+5kGfkwAtanXNtboiM8zCnfynrpal6vrpwjOlLHTf+MuXvLqE3NY8
aV01XgbfF1I/PSCRU9+BtuP8Bz8FZbLjF7XvMcqo+TuYwAKCmmJpMHod5LJ+PVSQ
0jjrqYCxT5NVkqTl0N8WyxEHA1Y6t8pW4wCmvz3TBnb+cSzjJbFfeBL4+GN704+t
GYGwRkrz3pWcHizK7qIaOt3MkTz7NgxDkJ6oDXhFh61xvbPwFSEt3GPHBfjbDPDi
VqV/qVW3kWQD/xcBAR+nsKPqqEyYI9WORsmEEkSEtQYcaGTmKZiyocpPxkyWs6ez
PfJHfF8kP2/hl3XgUAnbr58yvyMz7QpIF9pdNqGplJ1xivfzuZOtLlilxzABNoX0
c4uglTsxjVWnz7xlaGx6+ijsFQD4KfDw0JRbTjw1JIIS5Q6LBz8NJ9swpYdluLDU
/f9e57Vxx21E/9OvRjqBTBcZ7JFAtpaFhvst2L7EOWRme05DSbCcXQMpLV+Kfxor
ohUviFwwjhvVvDiXdjMu4tptAPmzpTFOJDF4AyCVrqtP6OyIZbjxn10yzCwLd73i
nvLW6lFGWoSSlmdWNv1GLBG+dXY9IeYTqk8wU+ujVreXeG+chRzlhTK/mpmSXiHn
l0IuNAwMswy2MdJqht/f1pEz1WMOy3NIBsUcKfbpMWtJjkriMrfsAk2izLVjLYyO
fYh9Wo17Z4RDxG0N4MghdjERqRv4sOON09zGE3I7YXM0X8Sa2cQt9SC4MqUmBH07
H4xv2J69Pz6p1Lh5o1Nj6itItt3Z0lLXbyIradn5VxXPUBxBsY2h2Wk7niSa6kyM
mt7oIbyXMFMogKacyQpHflktR/GDWrkxSdZ4Y2GsGhzVtuJ2A/zE8s7U9rsLs+KF
CUvnQWHEO99fqIva8MuFLQpVgqRJbXesiP7CoQRPUKZfjhxsJyJ2yp/29mrt3Nv9
vu8zBkNf4HyfNrGFu2zoAB0b5epGLpWd2lQuAocO/8LssS1WZZQ/MGp8oWPiz/4A
eIIv3XeTJl01X6/VA4Fv2k71AoqHg3OyYUcvTivVovIMuoVP2JvK0+QEF+auGnOc
GLV8J53+mF85n58D2EL9A74jNvS47h6uOvPVKoj9n5nR9dM9AdFdAd/XhVH14Frt
cFqwL9I7ARHjXCphpkpu6exzagnNJe1aXfqGfmD3jSMj0y2M4p481bvKRX49iwm9
MmaH3LAWjJlXisHn+elL9vMm18pHmwyMnjuNmYbaMTR5p5zAmm5+Y4LTZPmtFCZb
t/8lxuyKplBDTMCawGyGckYgKGahYm6Z5sqqVgLfrAcAFYcsDlQ3uHQzk5D8Fo9K
Zmmh1drvsliLmxN5icJQ4TzKkDcW9VRxO9p/YY9h+AqGFizJkGzromXe+VgGYQc5
AtOQpt25XRg1Kph63PqmStOXFbm+hgxtSMhyItcYYmf+VpkMHR4nw2T2DWrA0T8n
CyBi4x86LVoCtoIRMGGIY06xODTXsUZfghNF6V0VJUvHd/7RKIxZvl3/F7eVVqAU
mEbdnIPb61O8uUDDRSCKZk9Jt4zmzoXXVhm1TFGFnKnBjAg0B/3d+b9hzI0s6PQe
JjgLr8ybtwNQbpA+AQe4KGrKmQKCiEn+NFsWngfOhrVqKKGmTAAHd3ecqkrK7fSG
XRoPlqb9yaNk5F2xOomWcluPmZ8J0bhtyccFC4CYISIusoxuMMBC3DbELA7SmfQj
D/BNN01bTOvLvFmn85buscedUHyB+Iv4mJ6LZzBpOSMhcv+VYARBoBBBM36Efghv
6oHxz6+45FZYf5bwflZ4gAu6S6PBa0RG2CxvGsjMtt/3qNF2skPtn4y6KNbt4Deo
euuzKteGVbpbG/+4DvgvoVx9EMfA59teS2mOgK07/4Nst1+Q7X4FCB+cusHoBrji
mcFAo34E2DQ6pJuT2G2wNdXc2t7yH+IYAiA+OemKUak0CzRioBWXQFgJWBNrboV8
tmYxjBJJNVK9DFhqZmwUNjP/8LMzTbaF2TxLZ2kSE6gwAl33zfqk5utcmixqZ6sp
ld9QIW/da/ipP4fgIGVh+VFR33O0wYT7P7OdAVblV/PX3NYppyrE5/Stcw+9BD1h
SUUlNXQZMwwvy3YHAvZ+zqjlxFsVU1sI1q9WToNmZzMjYaLMlTNO8d54DYW1dHX+
pHkIrG0MUru5zwa36uTM/qx21U71aNQqgB9CD+XsyhBI+7/gAVzttCPA74Ojxkyw
wZHnoRwe0WrP5K0eMlvwLU8PPsFcaQMSGPl+1jjncvnqznBtN7b17fQZgg1iewhW
xTT4Y7Z/HiSpsDuvTqMhYZSwCI+NZLqa2qqb3waA5+sWB3FA/x0Lnqng7Pua8/+Z
tgaWcTc7TeE+ggdMKvv9y5Ax/OH6twszNRHovZkL7L2UviLb+f/SnGL7+zKqj1vr
0r536+55NJSd1B8g0kMPTzDgyyng1NTUlYT1sY7ksM+LS5Y88JOZ9BsIi4ljrFWb
GgkaiGkUY88KFjBGZ1Ji1/HliajtCWkpVVMfHnfR47pTab5ElhUeGSlWjOa4aKKz
/JfKWlYmwJVVbS5UZc/bEiuFxmyt/Gn1AUQyapP9aTwXeY5IWI4zMgEkoAxKcrwR
TYPu9PSmjgl97lBugIYhd5TqumxfkgA27VCum57qjYDlaYDvEsLgU8mpSDIIQwqe
H7QkFFvC2iLW73EXWPYjwUJMakoI3tJ/XuY639CJjdyMMOnuKeZnAFxjcMgddUcZ
kIY1BGMURaNNZhTCnHGRtrjSDMhOEXl2JfewxNFrM1h6PLEwdWNl5aacaZgw8Ews
jlhbHDfuh1nSg//J5jraJpGsqlw4T3NKJC9NcF63eY6zBgiPhZBM1O8DmcLIaV0y
ZSB+ZZQPGSHQHtyE5VcDhQevqe4KvDeNzaY7XTlCJDHt0nq3VSDNAcq++2gASkce
jodROeCWI5SQdcu6X9eoSKOqdUXJsKSWRNkGWkjmP0z7aV+Wm8lA1Cd+rRmUH5Ci
VYAgOqDcbLNr/WZZHMYxHTZ4HPgBfd7Xp8D51vK+NgpLcYk8AYfr9WkHk32ZoYI+
rO6Gr1Rc64Lr9IHxaFIw4bMtzj8US40WrVSIKwjuIRGLfILsBsfPDmUIbf1K23k/
ZyJWeKwcaSJiNaP/4jYGK+xxeLgIuxUmD+M3hG5wBCx9gQnSmg5lnuC61gdHYUww
+wsqLGUGhlc1Gajk+5pkkzsqRZqIPOgTZm/JwUNtzIdAIYNORuP9hy0ZfKCAVPaZ
elUTErlrWoo/kPDqHZaO8tMhy8jmZVw5nqV4QQRYANTaguSxRlufvFR3KNCNY6Me
/VGSeEGaMRnZ0un3ssWci2sJ6+d3qtwBe0ueFqGhO2BFQH5bIhHsbIfkdW6b2cKx
taCyvuhNVaiEqIAxVB2/L0Rc/Y51ACQ2ZWpE01jm0WZ2B1Gah9cMAYloagR12Qlf
s9InHDt40P/WSp2m3fb1fWO0sh2aiGv6PMC9e89fKuKS01hXFNAwuWwb1D3RYUab
RYZip2t2heLrKhJeCD6+Jk314i6nd0c1iAxJcqSVY0F+WplpTNk/U3ExM84fzPY/
nqr4aZMkwzEry3o8g14hmSBepbjYIOEx83MpERRaFmwkoHNrcm4hihazjMz7uVX9
xZYjjjc0HaVHH/wzqceM2eVdGzCo37kJCDPSrNLlzNLLzP30/FslMz+pWYMoDBrZ
kKE/s61lAzTcpQOqpw3YDFWJNwRX8q48rv2wJIiHC38dPLgWrm8L2eX9OZb/+t8b
uAd9CSubFxqiFO6xc3bsY1ohgk0gr6wozz7NbeyLW+mGbroB/TMJrSehQXo2B+qf
9FI7wJnRKwvHzEDlVxfnbChMuy9bmsuEmdbawV2rlFEAPR9AK7fFXZDmY9Rd+0E4
9ztiW7QTeTiwG4tHDzExMia/CR+VdilF948J0Pd4c5yf3/P5uO8jlsBiFq4NR7LA
i/tzIYGPEvYj98f6GmrBhbK6LG62j+OF8OPQ3uAkfEk4JyLAH6kvasl9Zf6JnG6E
gqNhiktAGb00XKDqR1N5yxW3itd9sLR4zJB1nJtDpBHQ3qC14Yl5E7fWfYinYR/R
yD1gqijMhhnqz9t2TAYApngY1auGV2j8a77E5cOiQujNxAF7SzkeVBhR5I0VCuv9
Pffw2mZPtRbI0JLBFgPdmBcDQ1Zl8HGhO8PpihXHnq9Azg/fTc2bGi9in2lp8ohP
nSW98w8lobPi1IJZZmt7yhpD+ASTDT4ZhvgXoXSmKi1w1mm54nm0BFwRWcezB+kl
IaWfXi3Nd+YVci4pHJLHCTGgRWE3iA6BZCns7db+yx+5G4tDwwAtgW2ZMoB/gVDh
RMAg2BwUhD1S0aFCZiwz7pkmdsQIig2M5jDyRHXBoXgY85mHm70qesWe+WvVHC4T
DQDRY0BG8U2Ui/458K4Aw/R/+1XXi76yuZaVsHOi7j6K2akbA9ZvONMpvJtWkbr6
IYpYvySMET/KDlHPUcUDfgXbpW2q8hi8muTT1R4ehWH8Lv+Mm3g2DYEQgMb8m1zg
7aICx72dD1SeWWRtcIy/x8PQFhM6PmUdqsgq5mvy5zmr52zkg9PuzCjc6bbBa7F6
MMRHL9KRjQtx5zBeehei/KuoLob0x1UOAwnaulNyE4Z9xFaecSMO5oOREeGPxL+V
ElsmFI9gNrNmSlOGOWxPDyAf6nwMEJ0zAT1vW9qArVAfhuhOBgdfmmZIoC7so6D2
vsWz49kSvJN1XDYPSafoJnWkSC/fkHQNeUxc2lKqGk9P2WcI+8HWQdlel16YI+o8
usYAjFhf5t+uhWtVum7KY0KWKJildbtqzupgIGi8g+swF3zgJNhT7j0zCRwrWhB9
1Nhk2LM2oy5XR3fB6b0JfkjPUZEmJVqUxSBzgTgBNeAd8g67DCX4d91bICQSd+SR
TakzR8w/f1i5Gxq8D/U+BqYSJrWkt9g9jfVZSN8tfr1CvZLLKeDCX/Ms1n3HOR8E
YVlDuRgHpP+dlpSGUJtee59h+dJxXBCVVNIqvVPUzy0olAR7PpIZMRdojuQCiNLA
jcVdJsifAZd2VK7RugBgJGikJKgiy1k4toPmu69f9aHHXTqVm43SOs5zU964TLZN
E3p3GuNhnuX4A20EVWMvF7utiPPeqJi1DVmWg6w9YlX70/7oS4CLygwoQkavb8fJ
K4DQmJwgU1PGOFzLuqjyOsJI24UCW+xLEh3u1Kq3uH13QG9zYgxXoGs9r7x6KFH7
H4r8QrLzpV0EO5KIjQBPjp4b8AFdSP2UvIZMDBpQVT01a/Ud8OdjDDfz7ADQkHil
uRkJxNlAKlwCAoYR+K2IIMNbCCUyntNC5xCBMMflMmguSubDKgvcuMLliAYYKAcP
bUt6HWgenAJ14Wib5s5B04Spro5N/rmmJnsaBrmAzpqZXYTYmhO8UCM8m9fO8gUk
D9or6GDacBuRFtj+c39nYPeB2MGF6uJGPlpXTn7kQtVF2x7ftal9J3EEs/Jtyeh3
U8Z8FQcnfQhk6bNNFW2mXsGLMU+r8Gh1cAme7AfELLrle9Eir2c7NEegkFPRFkQx
XqCaS1+lAIcrvCK73ogyYapeO8f01Bwy+aQCehIjo9vI93pH6Gno/fo8+ZRzDUaN
S6IGoNUJJXDnsrZlETtK3EFVdraZWL4z6g5LWdTNNeKRKP50k23m2cz6973VClbh
50VgYp57o/LcJLNsuK+M33sE5nz9IbolT3bOTF5Xtf3MyE3FuGADiEmh9b1sFjG9
A2M7F1GzCFs4M/VQqY8s5Gt4YtNVWzMwItx5wauzTMzYaVHpk3XlYl+GcQL+7y3G
M7CmRKowH+kNp+46Yp/stXgMBzwWLvxsR/VIVkdOLoMxEH4XaO+Dqc/wqTFaKp9l
Bx68hywqPSvtbT2EXH/8kdnPPESe+aI1HZoYhtPjiNtu7u/zMQQj5JBBn/+rVwYC
iZ0Uipe0IItBXdqx0maD5jxoDdKM22RPaqpqw6kmzYHTm7BbMVZRL5/lHwqsoNc9
MyIA1Jk81GGpUzcgUhjE7V81JgGVZuCGsXsPkzulxcShpt0qjVYcFhPQeclXNzpv
+NqmDz4hme+wBk+b+yNoxfLBv5R2Az54y3xh0s58JJt5fdko7mmBHrxD6WnbiDfE
EB147AGPJK9I5ujo29jWDYHRif9O/43j8Qx96gfEba5F98HqR4amESNHl/+0o8bf
mdzvc+juzGen+YBNrSGO1kHZVBWktwOUrbZnDJAZ+GUv+YP5hSwxGQ4glDddoI58
449qSnD19fwBDZL4j8E0ruO1E6g2candzSFdcWNba7NVWkNPQb9zZ0ASrwo2LI4W
wXtFSWuRS00QIlkTrJmE6B1VeJi8BFlzdTj4XG6MDimW/QM5Nlf2j1EIjvH2qjeJ
IXSysmD0K1lx0SMWO7n80qZMJ6uBapta3Ayr2BP8q8IdZuF2gOiKJxnXjpjd0aTs
lW5aRarAHZLjKyU9PYJFq+j7xFn6oSnO7XS5LWcvZ5bwAys5k3KZ58tpFf53WzHJ
RbartBImi4z3c5YhSRGFCuAFFe7Fcds2E2U14zpFbDLkqtjZe8tfYOtTS4QnVhA1
/fMqR+bfCh9MhqCDS1Zf31q5kDags/n3Xrtll9MyRNPmttUggxos+n8gsIxFxoiL
+XntZZ+srFUk7Ozcrnse3+2JCNmjnWAeeazSU0VMwteLumoSOtrVcVK0/B5ec+NL
IqeP8y/fnVEY9o2hmEqQo/EazuDJqk4nEVZyK+kikamqbyUGDMwPwyTdvU1BsqZc
9ef9iE+ojLVvxcZyD9wyegepoimrecY88F1WXq2wQbkGszHfB4EzbeLMiBGwku5I
cT6q6HtMdKc0GAKceZtFMDdqK8qRTUhAN7cp7vR8/3mJuir62aNu5u1Z6uDdOlO0
kna63g3ALf2sSUN98Y7vNXPC7t9V903otpUQCwqlDBLmonK1vgY6jxs597caYNlG
mXnzqn7vKAfj5AiGiCw/beAb34sBIHilIWCRG+e++YFHiLXmm6mzQocUQAzqpQMY
TNeDFKBYAeSf9Vj3tLoBzIJ3l/K3XXt4PbqAtcLJ1ZxCsUb9g8Iw3N7jfkmtWv3V
/hw2jZje8xN5WJvsq2VX4itPVY4rasUNwdfnDYCAle+VVez5Innw7V8okihExROk
uXDXxd+xL69iINqkA/mCRPz/nTZa0vLfgSP4riSxk968xJmK/jHx/B634gpmmrxq
VU3X4MISOrNWQ7hZVXFWJK2crbc5BjKVse6HgeM0snL10sqA2hK/cxRUPQfz1fz+
zZ63K9eRtUQ35yJM25MhP92Riyg/zhUp2V59QJauGX6abDHB9c7NywUxpbhH+a/j
p5SCmF3eLycsarFyJJCu7wOiDVCc7CBsUUR3aCPkn50D6KrCKrZehAwQoeK/s9HF
pcmEZm8nITobjDjav9qgvbJDZwZiS3bSS2rgDfvq2D9nAL4c6QvYMW2p1Saulkhm
8+a3utjVxua2S5Mj/bDgBIzLyVO5s/K8z5uLf41X6ewxZFNQ60COYbPjlh2vdhSf
Zh+rRaIWQokKKeu5XpdAy9zQQqsSEbq/BGhXavSpLQ1cYQfhrE4JHT9WrcFbx0eD
xSrAuexNSjWCXdApkjGSDWUusl/OZd8a03YXujvz1E47XBzerb6wUVj/bGaQHY9H
Dr+GlrsctFqBPb0x6a2rZvxmTS1yfRhf+sApCyBk2AtzFDIcO/SF7t9QaHiYdgnJ
qC4YoKSEwtW1x+eChmuVZT4ymIL0DHYoMASQh35f/6bwuh5g30PV6L5i8AQ+9z/c
t9omDvkbeYE1kphnwgXI6NNd5RE4ulsXA2uca71NBA59IeIJaao6+Be0yF/OWaKg
p512MeVSlajzuL+xLPF7b5Ev+CzIGFHckLQgLZTxRixECXKvpE+oyQap/6UpcSEN
74ErgEPH1YmBK+GGO/MKRZ58ha4q3RK0CEbhEc3kuF2OATIyi6Yp5OmO9/WYDX1g
XKOptcBC94mxxORdsNQpulP8c+8sIUErs1GvYvPvkzt36ZhQGaewJXNjEP2aM5v5
natEU5aoYXqbz6ZGu4xvtDTQcVCyxyjD2IolTthlwBSBBUIIE1eh+VkG9b5Dv1Ui
9BPsIH0rQgnnqEvpk4Ul0vxlgCI0rQriCxhLjj+GqJ8w70jvO1JFmGlB5lgWZPi6
XpP3EglOZd24c84winCHivqbGu2mvKKIGVvzDKNg5rV10+jiy8mM8VJdHraZmty8
5TNy+q1o89i6NMZ3JUbiUtSG0FoUqMr/wZjrqHb8c6yJcM18CIdDFNW8OD+dJoIt
k8fCGANyeTWb9HwTZ8y5xYnMJfsMExDlfKB0eJhN+QLJunJ5SAq+Abhr6RF1tkQI
r5dGqA8FBdC5JV7CXsbxtow4PYhtagAruG5zHMpzci4l5b7c7nOzXnFTyqoP/rEf
id+QDh9+DE/5IkykD88eIn9brvquLzKI++bUH2erWt1//WhI1X86Vo3ooGDMa0Me
DbSZ3iidQr/2wwOUY0v3PYqHjxOVm0FPO2mfmE9YokcBo0cJvQdxmlhyADBHDFX/
D18b52jrgfPOXtTnkhRQ7ZfFEhC/4+sF8nuGqthJMLYTbpU8vKttAc7LpgXZtTFF
foqGM0qSvCgRHNz6AzM6O29S7qHtRmUokKa9Q4fzjd3c0bcWR90kXgkFAkYlAu8n
ioFZFBzfOfS7F3OPBoOtJs/crfzmfUUscGYnmqvSmPc20pumOysk915/8QSLyFqP
te8nfNyJWtXWTZTH21smNC4IUxbXva/r1anXMO69CmEWFo+D72HEsfgfg4fjt2w4
EAF/QloVSTIGE9XHWSg+D6VCulFjRvlALK6ohoNyLfT0+lm2qMHYhyzDJrPeovF3
l1RdySXV0UEPpFdS1JltEjRCDr14UVX183hZpqNWN3MiP2yMmZoA2GOyhN/1TTuX
xSj8+XL0oHVGr8PVpqgcYo2oLs4167q9RCuF8E2aLM1moFVzNG9+3A7KWtl2XRTn
7w3NozX8ZLCeWDarcQABPQM52Z1tH7MlX/t+SMFwByI7uKHTKTt/ngqJz2ib9oGw
CfyDXWalrIeP6L+smO+x7UYOAFQkqZVt5uqbdvrVqbqQPQFduuPChXOYcyNgyRbr
Ey7uOvkYAkTeAjA/llldtTqXmhOMV4PrMqNrIXRkxdTrOUsHDqZe/6NlIWW09PYC
eSGL1YVZ/tQG7kWxvM1v07Om4wWGqJqlm1SgC3aU1A791nLDY5cBs9XLZcwf4B9R
wxOUPqidw9EEZkBJSLVeLr/xFt8lDOt0414C0ZjbHiWRDNnU17r5sPgIZ2nJKqdJ
+X02q0lAakKx83dkZAPPKaZopfNnLrcCcTz2ijmuJBadC+ijTR4F0jzE9F1wDKfq
0s/q6S5FB2xqlKw+b+Z+CwgVw9n4dx3IRVR0Bl9wG4T1Ee3cG/HecHzxlCczE9pz
nGixWFqwPZ6crdv2AbTx2ck7+3FpW5zJ/KgDFiWr1p8fVN493vZS7dv8Z4o3sXNI
i7za36vrJAuTwpIXiguHot2Hzw3h7QTqKLPmUjrLNBGv/sgCFZ5Jx3RpwVg50hcd
DxTrrKHheE/SD8ONnbyi4hyJAK1V+TIV8K4L2RtU/b8Iatw81ERWGYtJyN4DAavC
B/m9HUnO/JYOC1vXK+EIvScZ2Hr22o8yyA1y8g/x/3TZVJgll+MYo4J4RUZd7pqH
Djtd4fZGse9nxBwgJ38WlviXvm9EgR+ng5ZQ5zVVDaVZ96Gaz6AMxZMgrSpQA8tz
cxqbiurlpueEPtFkqqF+PGr8dTC9Rgfb3FIX5AMPQlB4nupI1CNHLZ1WYUefD1Jn
jTNMjorY3H4Pps5a0cpCMTiybnBt9JdhNbxWdM0rmbAaV9rRaT8CYkxvsXz+9fpy
wZRuAV3ZodMT4h/gcEhxnq/z/Vw6HTejFJ3gM3CdAIO/KjA0y+qYjCeyNJuzC+Fj
28IB2S2jzWUlUQd0eT8RLXq7nnPQHzfVkJbdCwcMq9D6lAxf5NjgLy7lkgkvd0jE
w36vvfnwKOPlYRRQbMGGYixY3hKhRgZaQwEIe8jLc/Z1cPrm9UByuZTX/M11V4lT
NZOJolhHWYu3JNnyYu4Yj6rn4NBsc6Si12ujQpGKI8sksHIrPtbL0NsCCwfyeMKG
KYTkJ9n0awT9AY5/smwgT24RuZY7ISLutTh6859huInhUx2AH+2d6nOHHgJFEC+g
d3Wt0oV0r0dKOV0XoYqghdD7If2vkbI0pWLNCVNvHvS+R3b6HiPlz2UzV/bukzzv
9RI6LltVylag3652TV0QXIXT4/EbVZT5/xXtiHu/18pctCruPygZxa2nvwi7jgMN
qtvEChiDlc61W7G7gIJAbGqzFF/Joy2nG5CihYfTu9oWt2/sEdo5XWCZHCwMqvmR
o//GUHnVJwOJCa28YlhQnH1Jd1zzqugTetCFvM1jEjWuQ5SM7hnhmQwTk3dxGzBw
dy1Hcrf/hmDyTtVcRWDtWO8ZZT4NaVU5e7VfU5BGJSjWVfLWVKH9xa4aAR6PTtsg
iNRlQD//4HYFvdkthPi4zsVSRTQzQj98ib+V1pl4+vyh/r4277xOlQ0Lu8oujb9/
MLKbT7Qsdp7gSw+gm/4RhsCSe3EW2KSi/1cMU8tUiJHKO4yM6GgzY0ZAm7HFh2NX
vgUlUzo+S5sks8Dawjmpd+kLxnInnxf8T7Ff1gDxMlX7FFBmMKZ5Bc9eo73zJHhg
hnSdc9VNfnpzQxzdoNty4ENayxYZUbOuqIhV+hGiKEJS4nXOdxVakjnH8iI7+Sxr
Tc5rxm5dJFGv6QAs3Hpo9qYq/HpGAHOJ7N3ZKIcLlGIgFD2dK9B7wmnZ7kEG6l/8
eTK7uyuTDKeoqkFekcU6HjskfmhxaDPyo0o0WANZbp+RweebJ4pMHBdD0QoaiC2X
3vt8SLPaRs+BEd++QDIsQQ+ewZB5UdlhtHODyzjxioyMV534wcd1OUwQXKaCH5Ys
cUopVxPZBoK+XZyhEI+7U47Jvg+UGeasyKML8dNMtz3Kf8YGs1or1wikh+/2DfVu
H3+VU9IiGcwVwqB79eT13IDezObHZrVOeCYMH1hlW3JiXciQWFjlzBziX4dVArLA
3RrUdAxqFZ7aBIj1YF9C2Eqa6UWboybi40/Kp4Ci/Ic+Qt+uV3t2/tiyBiPAPEj7
e5jTDyNNJjfhQ1pCXsRrn0R0X9/MvL0KTMMMg5+Rca+MgEP84pRWDocvFPidnzFK
MyYPooyFKJz6ZXiwv5BwZF38qblggAWjeTgZBRVptYBb1A4BO/7sf5zx2P9UnnGG
ck7SeT9Y4QyJfSFr8kCIo5pqMlvexKj8fPtIi1XhTELOhcAvdD+hjIsm8YHZz6FJ
oH9U3l5gyS0r5CB8/C6kPpqPWXWyBYoLi+3x3O5wkwX4PtQ8N7xH4ftveK6GWxVs
VdnYFR61i7UKBO5VIF+5NYXEx9nuRV+HtZI3JZzGG4IdWhdi30B6Kib11CzLn6Wg
+rTitNmAYfXSDzezPzLYULLZZIsT8ptfSF/g7ZQ1LmMVpHcWBWEFO8kw5r2sca7m
J31RmF3dBGstyikG+0IHDkEWQC0rCnVSYgKAJE/xUwQO9ykBvewEcyQ/idUh6FVY
BkCwtYCaeuWXvnssPPpUQzqfeDPmqs5Q7ZY9xC5iu9vWzblycJx9mrhaDF/A6R0H
S+sCwfcu7f4ddrSHU2RC2fPCFFwC2grAk+m+ZHQh/0dtU/lTS7gpxtB228PWZJTC
XoNUISpfhCv1PgerYSHv2yMwBMqQ+j0XNgfkeGYCoyNE24OUgSVNmPL5SqW/H3mP
la1YqylKdW6R26Nj3rNDGqj8cSLJids7k797tEkR4uLBYuWqYFF2hM+4fZEkzlxw
5y3STaK5Thrb1H4EbwTz+VSuFFmeEnGo725DAQEBQKu7oJx8T/fQtXmCMAGBAAFg
3eqH4K88ulPaaj7d8DUlh/9TA4eRNggkgs2w4dBPLwZhG3UKx0N+d4is5WLbwbQD
iyINAElhjr0Jo55ausWODM5ZmaP13cC9d2gUSouNk48IQ7Xra/tn5Jn+CNojUcij
8e7caW8DHSW2eoBSRyjQBjnhIZOY+jqTLHPP8Gh/S+OhUDjBIiAL5QBjXqz4j4lM
IRzRajQjhraBB7lv2PA9b3E9w5TAoErd3skK/WN2Id/3efri7Zx66VnB1dizZpaz
o0cRpHZ5LvpYuNzFf4vbqV8erjn1f1bUupV0LMkEJ3BhbKGXSWz6f3O8I/9HU2Sw
+GBz3edAqn8wcoWJaeIfjeuT33fhsUYoH/lwCd79Ldpkwo51lqpmf/aVEqGGLp7+
HhBiJQ/mLsZDg4HwoRO2Ihsd89T1oFDLn1mW173kCfsAh1Ab72N/mWBi440IiUEE
AA8FjWW3LJf0lkVcpoq0DMRkABxIwuwVLCRwXUo5PPDkHjKm1V2YRL8M7mw6V24a
fHtCEuXQIUS6B05OR4HgoYmKp5iqWmFj+uhGlWMM9aQg9EpPEBFiLU3vu7vps1bV
7ZaOiTkjEqat8Ygx+MP0WCgF+npUJuCdp/J53Y6WTjvDFBRAPJBfI+JiYzDpB1LY
AeIoUzouFRrDd+yp4YObJlM3o6VN1prDn9Hc6mfHKakIHNPwBEYtI7nMipZ1MD9g
4oFLUQNlaXZuouAHZhXZJ4CTFSrWBhdy+g4U6uWwQ+WLOWCM5wRlth8P0lIPiMXz
vDdYQQnMY1r0/RgZ6Z0gkothOmU/oFvW3dKTOVP2zZs01lnlzhIFYuBHysTB8NGn
mLvB2E8aSN+yccsNLETN22IeGC5hIEdZCKpb8hdYZDiARHxfa9moGKWRMBCr97KF
lvMgFdPms2JckcuzmkBModze5pfYcw3LpYplJKd2u9+0M+go/G6Onh+Kq9kGLaqS
jVngVzLAJpTMhKw8k+Gy7g3+jtOKHwYe1w7gsdb1dyA1+eIP8ZmkJSgPsrvsW6+R
QYbJOrSpl0k7pTvWp/1H02vr+y2kgBidEzaoyMx8t3HTg8cRBDrKxERKGyvcwPtU
iRrb/+chIJ2b8S1c12BPUYEGFJXatdg9GxqdTyDLyK/J7v74OdHEm2vMBw2OhGkA
gAKrz6yS4OpNhQAMQJEjzrfetfGoMBOMuddqOe6ebSYt7noComuI7dUSLvyhSpKk
58kIemvPppRB5GsdlpT5QM/H8d0rYNY6ePU+jXvdlmIHbtWrihIx5aBDjxWoZE7F
GzUXLTyLcO3+/GgdWpG50Zi0FHcnd83JgpiBv03EcJKaMUjrsVCEV4CG6NLSvfo7
ELmipB0t6d3IE8xiUSLJqLWQmCopAuhZJe5tQA3uTDfUOAftp5DgP9uZmgylUxKw
F8doHdLb+PNK3LQhGxnXGinjMX6wWl1WiMJO8+ylCTOs+gYJr++nxkgPV7Oh4Q7x
kq3BfLM6eJRP6OUM5eOwhkdCqXneQpJF7OClG6+TlP5/NOaYS94VPC+BEDisjTC7
atq+hYQfDwCOVApNHcyZe4HfZpjSm1+vSXDAn0WwZPmx8YZwHOEO0Ml9gtOYkO2+
x+5uI/cxGVVdX9ZdZNpxlQjIJNvX7gcxM/eIFU0hU1YQMWiIxNPD0xVhGY7S3xGC
OVoY5CiE/Je/pwhxvDKzn4SH38VGkbf/IxcB+/2L/V6myUvvOdVbQRzi7gfN7lF1
gAwxRcrpgFVhOPqbe8VFeh5TQour586RidlIURYPe1iiDSncZlLu+XyIyK+eZxVu
wU1n9FB2Bu5ysp3zUcm6Zt66IU1XuTGqSXwLnsIiEdsZKuwAa6ssJQMuvl7ScYcV
3efXz2Dg2UKS7W+8BI4DUT2s6l8sleusETuucsjBPoap+gUMwzeWMtXXhEm3+oX/
Yv/fHPPDU5o3zojDq+OVicxnSCpnmHdZQzIW0Xl4FBhdaosivkBkurl5p4+CXrqK
+fGrbzxXqdhH+TX610VT9Gb/qBQbN2rU43yWm2pvbvFCuWjlyFx6w4oO3vW8dqPS
D8XMPjwkO9xrQRp2oAMk3gWs3az2fnk1MMy9t3a0+zChairJATEWTeI+k1Unx/DL
DtKIS+A7SZF4RHQClB8W6Gg+Rrpaa2ZedcVk8IC/6/EdGikJPj4nlKmxUo0wd+cm
Lmo9oL1ShjaA+pyApc4H11hKM9YvjQocABIzYdaQHgTkpy1J5K9DlZ82+SZceipP
TXWEvccqWn4+JF4/H+FLgRPkESNddm+wtTcUZ81RfmM1ttR7tzZ5EC2zWAKnJRhY
4BWYN3+Rw0WjvgfeXsyHR0/Cxd++XhaLWmZQ2rWW0TUPQf13YeFhlCj5sUGC0cG/
6tgqXiwEkGOnIvI2hc5hTtwue+Mnbr3f9Qjxgks78uGWh4vY9ZC2r0XCCm1DuFo1
2MAAHSZr4ax/THXsFTckRDUm+mQUypwSxzRpjipmWPLAC654DsOJbf63FxoS7EnS
3tg/0FzM2eiDIidZRjCzcv8Yevh/EVp4n6M244BgeorA2t9J8EuouzSbHzdi/q1z
q4g2NQutZzY3qnD/LMd0RWGFnotGARp4qdqVtpLztJCXBVrp+psnxRVBUGgDWTvd
Mg1ieCKTEhd7gdXC7uLPYzfC0TuROgM6cUqpTDvqsJP96QIJtgnALBe56Bh/JSIO
MOdHjnQ8wAoX3UqYxCCA0esA+f5d8dGK5rPqZvGbf4X16I03Rm5TVrpiY5aWUdtz
f7UTifx6+gHlU+3wxOfZF1yjlYbNPddpU8B2SCW2FrNN1T1BEGNlLyvJqsFnEv97
iW61zZhOsvO8C9QBQj7e+hEIPCcTqsagvB99dDkX/IPKILyoSLuB/VraK/WLx9SE
ZqWGdL4Wc51fzpws2dcRqBgrec75B4rT+JMdINGTdMde4dYsNmiWaZBwdhhDrbcu
mZADxT4uQGwK7f4Cf8bRqHg4O3B/sRfSaThV9aiTPIO3ZSkrTkxUD2h6D9qYz8j7
Innu7TiQGOCqFKfkEJ+YY/0WbeX3ASwTgUZ05JUclF73O3T0qlhumUHht/qdhToG
SMecRmYtGp36gGep6ja69TG5Qh0xl74cVCkCwJURUQv2dN2a8z2V1BAkNmevVhJc
QlzhnC+Pjk1BEa8ajlbeUaEhe0JpsjyajOas7I+l4dT1H/59Z34nEkOU5AVd/7Jn
u8Ds+J7t5H8JEiIcZEporVVK4h/CWkCQghduEk18vBjeSaK1bZAoeCnWdvdyb7/E
lw9t64yga/sD7tIRd4hrwoP653gWYcDydZs29bmd445a+ouMzWUsc1LbH7prEYCo
AUce7/KJhvGZtaCPQc+b1oy+p3CoA7/Hsl4eC4PcyJwV1aQLDyXJYh11232dYBxw
Y+qo7MFIqNrB3S+pEff74gK9LnK+xYWO8cGsz5tcT7ckMvGMttpsZM54Q/5esuGx
w9Ql8P166K5YJxpF2eLjRL43rG+HiyYmGMXsmYLxeQ+fcHivQqJr/WOGDCF8NUsS
LxjHaWO25/MerqjiWXnIsbJPOKPNYbg4TcUT5npRXh96SoPNLZZQ2jd2Ca+BYk0M
mkprrHqv3zDeXoQug1UK0QJcYz5mDHposyMShu2xtuotm6pPl0Uk/jiYspY0at7f
e7raIBWvm7U+H0fd/oDyy0+5YVUImb3a7dw1kIyG2GWFJ7AmSP3Fd5ELGqFeWzYN
e2hqvLctgIRsNtNltFlNTRPH6bnagNvhcauplpfOtQMGNsATyLARUyceV5UC2UxH
F4x5188cKLFk2mfQKXInyrz9z7KBp2qfnXOCzYztIzuhuVzNkHJuVIW9L/rIVHWd
gyuLxlSwGdqAJwci8FD+CAst8loTCBsYwJGTWGDtlPFWLNVmU8bOWNLGs9oR7g07
0mcZv01swfj1TlD/Xyqhpth+QH5IhSH86q1X8neYJE3Oho6bUGW8d7tGlYyhbvCT
YaohBGymrD8yAvoGd7MpQ9Cpc1mtNtXFk6ENBvdumB5AZYr7/t2kT0HbtBn+SRm0
pXmzlg6MR6iBmD3JcM2eJBbs7x1m54v2qaadcq1WdU+QVBfCMrwny0favgajaDNj
0zZ8skwh5NKtOhwAZVYSnApmkk20iObQPSje58O2W0MiQCvTQaeMqLmQgshXnlR/
d+4iFcJZWwLwSSVSyx6Gyu8yZPk064Vdb344wSdeQTqOH9Z9awl50feEqRzYwNPF
wRgPFG+T4l9tLdjK6hLV+4KXHDXEvMEnSfbiE84crFNZE6IK84FAPC7iRiLJV3uP
5hRpnjEeRny9tR57CndAUUbJPG5G8REf9Bxfr2TQBkz0YfFISVcLlSir6Op6KfZJ
6S20qejJdQDGwhtJMMQQzo1iwF8EyTVa2XYe95A4gzETa6xrN3m6v3UTuXwkgHLT
5VwIFzqypTudBkIGF3/mfVIizFryGXwAJWuXccJke/loCagtg8rBTBZOt8rfoqSB
dtNq+SZZm9O4El2vsxFuDxAXxY0SVUcXqDZsxBgFD7fzhSFXbycppZ72eUaEeEP0
7fMv3YuJiX9tVQTsWPE/N69Nthf89PfEREOEC/TZRtudtXzE99gqDypPqu1suc4y
+GJ8kozgPOS1ScRcaGGOpc9m++2CvsGeqAJLJD1mHSZFK+jZwiRLpbQnbQO7fyhP
aCLGVKzSvknm5bxu4JzKlbE4Gu2upZ31aImb2U08BjG+en6NZBV4tw0Fk7jSeY23
s/bFkXPCRl2VSUk4ZyWQ/3haXL13TiourxCvSgxGcfVtRq0mJUaCMT/Gw9T9INJL
qE0bO2b5Pw/3LrFJhV59Pk+WtqIth3BCGOPrLpggNQeXT6cmG9rivASe0259/00S
c6N7+baa4wfcl9uotliW4XSEAaODlR/YUdYpY4ecuZAO91tJYicPp7fYjIpDIkJr
olPbGbdoFWct415o5Ml/z9a1ZTJi5q15P0IWt8YanoV0aRaQ6lKYhn9uQIMOPrdV
CBgFOZ43wjJRLqN3wWFYWvgsFJ17SmiUURtAzV4mG6/9sO3kj3eHD9UzSCCldfE9
3PIfuUJeoQOU5m0Ao2fn5shwCcr7SxZQKdRvjjWnGYJJdCLJjk+zqEuZNLw48TcC
ynR/sz8DocNKp9Hh3fibm+i0nVbnK0ZC7/8T/y8ewrk7VibzcpeziUbwa8bhPEqo
J+0neqqUrJwDeoXDK+O97s7ThOPJEr7szzt7D++jir3ForSL0pupoIgdMs0afIw9
EDIZ2Ht2iH5t3aZ1WfPnQ91PzZ1mkLWmoEL+buKEfkb4Qu6rzvWfpLPXaBEIGz2w
MG/3s9h+JzY8QhcBCdo4r6Z6alxnSgPMjRhpnkgWyn/kGAugEOQScapbFDH35S3C
52MWeTE1By+ie3+oTMXyitj23mHYBe0Ua/52roD1zT01CrcOPil8xahmZIBzjF4o
S5Oh3+zWoIPTbNxDkP6+kJm8q8Tc94Lq80q97IPjIoDy5SIbLrrQ1cF4veQofV9Y
J1y03tVgS6R37rdP0mpX0WpbdxngfuX9rdqhUtBfk8thmbzKrQL2Ilv57bPSQHVD
/zwo7ZE7YI6SKGhr1dgSJZ3eeWKLAyHD3qpeQxwRAyRGHsB153B0a6IWY9GFQag6
d7FR/zUclWTTln4LfQepqSNOrN+5XdWe75KVc+x/7S+7e9ZTK0v7sQBYTgrV8um5
soYvdQ0Txtf1ZNCf/s6y7mGRElFTClnneyRnfPxxeRP4UFN3qxG1pSN9BE1cXHHO
JXAB8UojJP4Xbev7VJc7FpusnijoGuFSuZ8pzKWwAuFhbZXRZKB6ZNvJQ2CuFofG
6HDzskBApb9T/aa0GqhqtamGr0ulsJsuAuUPBpUCxPz1i3qZrdYPBAKtCVwxUPTo
rXpkdBESWYY95wPLsumaDiS8F/OSr4PIQ0CZNGomPLt3R2IMcttvRhaI7kLtE9Mr
T+E5HdkIO0UetqEYSOWlvBYuk69oti/bqv8jEKpdeFiJAEMaJP6jKz48PgbV/h6q
WrHawu7zULF7RhFP1Tqh9419sHv0EpFZ9njTE2yfxyyuDLdqnnWraq/zfR6zSydf
wO7I3IV0hau0Wxv1y2hOg6yreg+xrByiVmjWDMZaz2CENi7H+taDJsUQa7kL+a+m
1cFdQrtwj22famxrltEJzE/6sNn9o3BbTfhwsULKphAmETZu/F1ONJf6u6T/7LEN
2zaQwVpmMY/8Uf39D5EIxxBhEtZtRLye53AOiXAis5AW2fRuXFntluc8Oa1CM1mK
DJygP/PAJCiBC587TxmZXwXLFFDKn3g8fGKcBXHlUY98qKWfgQGRp6vEKu7NkMYy
+LQATWJf3b+r5ZQ0SIOU3XUivlT7eF8V3BwrUgxiDQvQblLuwFAjSqZXUvtjacw2
2WyLfwRdePLeiAxPxVjuxyAL1efPYjSrKBrVGCrJtWh6qkljGq99VynluwFd0RN0
FEFS5ML/9TftXixp65MQsbyd8hMwKGiYU4g61P5FYL4Do6i5YpL4AIM16coK7CZK
vr2pWY0f91IvFZeEtbuPmatMQuqPFKk57H3uSXeodXhRqcze6IANzu4TlbgAgPtN
TR7cq6badneCBKVISu15aUkmMMs/h35XZQ5aT9tfVEXQi2KUR/YWq4K6svvg/ekP
XwrdogTEieztaqOAGBjFTCfkeyi34cWU6c51asi+POpbzBFxQ5JkLExdfqXtRizF
hBKA5gtwH+a5PvUxD+vVxeap3Iacs5WtYeQWEE90F60gqqr0GCET7FF8JXiuNXnF
k/m2CjlYn9l/aMRolHUUl4iZ76z+WAmM8DUNMODTSkmVJtAMX7RcDiR+jLt2OV8E
mR2aEua+IbddN5+rEQc8CsT5P8UKM8kSMTuI+hpgb4hbVvxGpznRisXXQ2m/hX5z
x7U1nVQ1pL0jG/0dNhIpAFBu2G6snx4RFSpm9g/8ZzsEDtT2MTx3qjJUW1BTS2S6
bVQcHHmCHyvqA+AdSebmgJd75q3c3kJ5JcBI+l7OFYRloeu3EvdkgYTe3X/7FUdI
I5jnCpxLxd4jLc63rRQPgEzWuaU01K9rphTJ3OgsG6X52y0CFedPQWgyV5TtYVxO
uef0/CUkORC8/NWVtP4CgMT1qReAIsutIbA5VNXSMKbCbHle5LKNlqfJurURSr6S
ZKPGy+BqNXQDDRos4dqK9kiZIn5cZGjVUFaQv7M+eA4WWkjw4QNmfFD8p6fs22gr
YijBxRVzyhWmtM1ptVn8+1vfoTiRxz8VHQoTvOUTeSKXL2SC2KdVr2pxQCkUo+/p
eNzRIfOqMFV5v+vvlUo+sPnMTG/MZF5KrckdJVEuARQfHHlIJNvH/n8nfsMWGbpZ
OC7ZdVqlRqhApjCPcn2Ap3gMq7EYztL77hUTV45dNBVivDIiUucOIBQbiSXwOHcX
pFRUvJZr1ZhoEuGjxhUJo/MCzZWq/3vkx1WNRN4kkvy0rwIbhlpiZUni/VyI+mWq
J1Nezn0T2nGbhtRkpQX4ImALtj1EH7WbBSyvJo8fROB2EosC00LQLoEZIHVYEDvb
4H0yCIExpflCfqr1RxBncAxl+TrA9PstNQuYJZosguNcWVd8rr7EAi+8cayBkKFm
IlEivLuIyxY+tlIBPpJE4SI835MSXLURtBxA6mXRdxAM+/SdvkKeRITguiIFVX/L
z9QMCVBe8sciYJeGjM0ejuDrspw5ZO1mCwtsEeeBx5kl51ulQ13aGo7NKMpGVd59
MgtCuTN9CicHN4rZjW9dK2+99dSpCfxu9LODrXzPtDfJ2KAF1Emh6uO6FwsoIO4I
0qB0zYkQfLunvRo1l9tSKxKECNUaoXgltSorerG6EXqx/fUi8WVJh7Xxub/gQYKM
kjGY2xlxwf64hw67E88XIE/KJjPskq3YUprvPvF6V+0x8MhMtufv6Sdth9sZrMuS
Y8BT4RiS0s2QhNoFWqfFuFoV5JsUa5CMIinpdPANKnm+v0GGNVsnKROE0EOWCawk
UVCIGcts5V04Be05+nSa/QJ/m+kG9B5A2F5bUadihu5j560vO9Kmi/RoQjHZqBn5
GKZ+Rb6R0P/9OgGil9dHlPkqSvccxwk19W7W6pyFLpijJ6HlYoBXpHzwen5dyj7/
MMxSpI382f3dkXFnvXcjLq8NbAxxbwCxZRjM2dFSmUMMdI6GFJRQbXuqalrwQsjL
ZhV613EwP8nW0h+onEybL8Oo17BtcloKtu2KaM4Y23BPnJi+FjjJN/LyKVXP3TAq
OzJTJxfPzDM89JAeHj6RaU027K4oTEZDB7miE02cME57HT7SJlv5EJWJ1nLqeECv
fY8mZfJwivJyjr57QVOXRdrI8YidUPQmck7EFMMhL9t7bKK4ienktrp5i79id5Wo
4Ej3HzkEP5KZikXMhno8YTxRq0+RCGVbmy0mlLZ6ryZyfRBmXC/z/fedDYlbO0aw
vRAnbSafw6rj0iraPuEnFkXQHYAnGh1GrZDgox1khsccFvtKdxxiP6U5Y2HkujL0
Nfpdk1xJRl1Dq45wvBNL6M2pKF8EMkmSM9noU3aAzrw6w5X0xR/aQsAvuiz1y6R3
Q/5EJIjIaf3NYYbBb8JMDDqWqHW9xQvMwWv5WXgB3Zo42AbN44w4XgcWKAx6KPnQ
la6tGpYtz6iXraWxsO80JaLG/n5JgB9K93IJJru7iJowg//RR1tFw/tzcj03u4+/
vTI7kNNx5+Zb2T+qBlVHBpVco0Hn6+Aqj8nHyocDHeGaHT3nG+b+3I7otgz8RHOQ
2HhQAJXzaMrp1ysFsT7yFx3FAZHP0LVze4PJ9FBzE7Qgk1+NBtRVapegFPjJrQ0n
eY+Ryvpk5GlQB634JvMw/cwisp1CLmn/gglFyMP0mEr/BECfwF4bIL7UxSXQ+NdA
HPjj/HBIpR6BaLzrUT2F65IQQAqosBnXlzrfVsbzWPvCp+vTwXeXwqppy+mi8Nes
UwbKqGKtOUBetBcnUfAI859g1rz+PDLvIJi974lAkMDh4H5/YFuOPlEIxAbhH1pc
raMH3H+bCTAUu4uuMXUlPE/2hdNjIPoxHFDxlxq8LpyzLMDLAQlKjQlBcgXV1O6S
3uuXqtPSRQD7MsMRA+2z8fvw6UakW/sVj2Z6qQlkREKfRx6Fc4jMQbi5IRzQ0LBC
7MuEjG6z2uSyFkPGi+E+DckoVxicE9Pt5oDVhoDjVrNoXWabCZzgh8QhglUFZnNm
L9972rgFyV1nB2BtzN93HzPVJChWDNwAH5mhOIQoQ4vuQBap7B6Isd8/3T4CO526
BtSGV3x702YHivmGjSFxqpTNwk40S4XhIZ8Dh9h7XKWxXRWYhX4BotmTglMhc6bW
XKTVXJStUSomT1VCinEygrYU4WbNi8xBKV3Q+nT9L+jPH/Eu8TL8IgstDPXOWkqj
y/xRe3oRZaMAlvAdiRPYn2nTpvafzT9E4SJwC9YIgK7slskcQP1l0Y7D6Cg3MyOV
zO8eUDnS+N9/Vvf80z8XllbML8DlRiJeDSwapQrB8dt+v+lnBlvOvM1Q7aaRAop0
xkhtlsBJt6G0r7cbkm05mv9xLFSLc9fBO3WMQL341PWx+XzD+rr5G2D6aTfqRAX2
RL/n0yHhOeRyVQLAzhiGs89zkN1iKahX4g830GzOeO3Ix5oXrFU6fwEv0HIh2EQA
RjPBL0utj50OFKlKoFD/2SMRKhjYvWX2CEUXmlcVwnnyk6H3jLxdMMYCe/8XG/85
nAXgAC33n+cueSxw4gnrVZonPYLSt01//IbBihNsXOb6KLTcqs3dESG9ZECOGxrM
HWxLsONuCUTPpIGc13RH4fuqiVokynYpEtXIOYcMnaEI9xyOi/W/EhVPtY/jwJzm
srcLHpMIySdAY7ZxGiIb6okLGtkx4/qd5hDMACi7zyu9womSxuzIoT7eXbCkOAsh
knlK4OY9Pk58ShIojM9OsTciDeuujgofec1Fmg74hnty5wAmFvdSXczZL9ljJWTt
QAWwnZdTwpiTId3lpZE7F1+5Mah5Ak68NX0Sv+vOrsaYZ2KuEEWs3X5iAE6YXBAv
lRLkRjohEHNv3eWJfUDHifY00MFFaS95DdVqIpvX/W5TOo8za//SF4oYQS4iVK+R
53mkPPD1wjWS+ArzOvoKjpX0sL3ExTWH/PHSzySkyjxJONkmf10frG09pqbBDWPR
tdzCyuCtql1rcSF9OzhxDGvkKW8dGAxpF8qWX9knHi+5dOS/n+nuq4rNKvurvNQq
zypsnRA1nvQ6htNYlbH1kQrWfWDVoVZSSZMr96A0rFLruN07GhQFluC47taet8qo
khA5frQo+hyjgAvfAk3+3ioxmFwadTtfq7J3XVAMSSXLsxfAXrvY6V8fyaP4VTtZ
/jL3Ao8k8dX0m84U8t9WgX0xXlP0i9DPnR5TyylyWi52bDGdzkn+8eWd+qq8OrEd
MKlJ/5Vu3x1gLtex9tAYm+9KRh/7c8VD4bjuqEkYtMsjQk/VGyZNmtO+r5+ixmvo
hjbVygPIGqCnzk4jSVeaYQ0sOau8VV15m/BOqmSE583NOrZ8VAwS5G9zz8nBUgYY
kVgR8We9EROEhB/9sACBpbAmSe6uivCy3Tb7BeePCqaY6kMyDISzYpfLpVzLk/QT
vtkNpxk+I6VmTMvsxOqa7jw6EDI++gVAxB6YwPb6nZHIhvdtEuPAqysbBvafXJV3
KAIP5nx6kxvdJhfESQTDO4hQVZkcv3GDPiBpS6GuVPxE9ymznC2iX9ZBPze/Crub
a7C6o7Rz43PF7soJqvLhem4f+BlFnnioHHnwLMbD0D77Bg9LIpRobfhdZ1kyP5Qv
tu7KQL21tUy6hfkj5R72HB525bwU1S1iIbrlNgGXtJSccVkZPoQTTCH6E+hLT8CL
WBIXuQz86qjFIpJuCJLdOEyHYktRalOUulR/t8XD1rRKVubUSXJMSnBG4m7vX9VP
TCjzt1SJxHqqpQpEFa4NsDucShgmyYX7vQ2gvY9J8iYRV0g7oPRiwRn4zXWkPIZz
/gXo4Mr7KZu1KaSvN+irPgcD1XOhqlDz+RuGqO+4om7F0Yprjez6ZHUHK3p53syI
0bINf3845CVxXUqP3Y87EOmjNn3NrsRqew9VKCFuW8+t8LCt5yjMBloRLelmAuRt
vDKB115ushJEZRTFcB8VVn+8NJ3l+VSveCNaXaPJ98kTFL0QSoOay9IAAEUf1xBL
r7jNSkOgUKX+DaWbdt+/jnC69BAHJ/Yuwu8DpWBv1eKPlebRAb8HkRdcYBasHlXP
XXZAGWoPAJ4F7ZwNy35UBivZ8DLue8on1M7B1/H+Bnyk2mhmimFLOdhM7ZlZFxPK
e99MLuI7R1nzhzJndYusIVi1e+SjxJpJWQ2WcYiJFmqeEW1mlYcYLWDgEVN+Q4HZ
IdXQMak7t7EC+somvwZVeXqfI8W12PabccbQWLwTrOTHMFEfhxyTu4b2QccfiPDy
IIwVQeRbOASXIuODZXJGr7I8znvfYy6HKLnlCaOh1yqOyT7CSG8agXchUwesn7og
toVPCNcgkpu9GTXr2dSSUUxC+490wv1wHT6rLpUlu8jLYCsi4BwZbAuiA+Fqua4o
rwR3M3pg4eQxgCpscpQP7hFSduQS4TYJPMsmznfhXR6TcVynG+47d8vnuJm6yBXx
MOgUAtAZMswf+nYDy/7vYLo936qXOv6RPQNg5M/j5NbW8nCZtIVm2iT0lkXKlAHA
Tg6uT+VsXEcOu+3S00QOKeWM8jpaHmB/5zPYbhlzxeF8mPneD46jVCKXz6LrvCK4
e9hv0QFTssa6lCCrttFYhIgP1XXI7AYu2CRu8OjRS+Nqqmc0T3vtqDqXnI09k2e5
iF/V6p2RhWIoR/mw5Tc9PI+H5BgJb9nMhV9CPpL+gLFibh2kbx+EJqAklei1o+gS
8tpfwFU9Z4wrpszd/II8GZVh/NDRadpcTMmT0S9+9RsJYoflKn5muC0elGEzUWZx
u5UfHjby1DlxuJgkV/MHSTxJ51mQ16TR3kiNkkAEpYuIKxQHKxIHQdjN4XOntJVW
2p8TI0D9kGrgUHosJOc7AaqTnyrKyAcjWsTgHzk9mA+xQYZMfysiMMoKc4CoSUPK
h7Oybun38tp9E0aWx8F3x3eKsw5wLaha0EnMzXguXZzIj+0ZppOvdJUKvtRbRC7j
uEcmwJNuR/7dIxBEL9cAWFF5JDTs+9hAKIKQEcj/ktG6YqZk9j81mnWrzkGIrazB
vMNJIN5LgKYOJrxvaWdZbQgLUBWZKiy6LSVBDQRtYxOn9/4Iez3uQQTv+7i0/dSP
xjj53QoxvA/C6FFDL6cq4oenLMWx/Z4EhArGyjAxdJchwFdZWJxhEyrJIx83od5V
xnw04uXbqhnzrSWy6xtbTVzV9Vvyt4d5xSn+H6ux/oh/cN9NH0scQIetRZgz2a8r
q8zO4Uu1swYGU9FbLX/yfasIQ1eUg6/GYvgvzkGCgGtNZLlh3rAm6PoPMCLNS+B5
YWMJDjXKxJMYWtjIGEJHbA==
`protect END_PROTECTED
