`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L6EOg5yXxsL2bh7qZ3snuHcA/nk9LrvZtlJ1IlLXH9PRsLZfVj4NuMxIwewtYrWr
H4MzadUtJEozkc8gE4Z3L2+XN0kzQDu/0QGv+UfASW+3CHASfmuvalM7dLdc+5f7
OTZ6YGbwWeujeOyBBRsMWTr2KHcR64VMYcWMT2knaN/vhMaUFf4686oEtt/JKPA0
SRcHdjXX0UIxp5tCwVr9lb14eaD1GTaDYJM2J1gl9LCURLIOYzdmCIGcRvaezGfB
WZrt/MabfPVHMRw7p8Pg+PcYW2bnEAOZ9kI4XDBIIUn7ExWQjMOi//3kZJsTwhZi
ulE2YK96162e9CfEnQmA6r3jr3in0yD/VlQOWdq6l77NgdoCwR5CN1bKx6BjTCHQ
pX3A+JEkhm7VgLdTRNvXkfn29b2ua9kXTG2r9al5bFyXfqUaoFwctdhBwMb5EtL0
VBUEo6zVDW7G+F8JBKW3ptEzPPbRKJ8i63N0nx/BywhpuIzl7e3rxjw1ifEVmaGG
BtYjDwkqJ/BY15UJF3bAwkn2XhCZtgiStv56e1qECoyXlRE9kDehQh6TjvJsj6xD
FVAV7O5kw5E7+FBYZxyXnOv2+7PrgP9AqNf8bA+n/B+F0oZYvRNT3IALRlORmDmX
dT9Bv35fMPbUONT7uOqaxIZekX2uA3EuPHRimqUvQBXE+tnu2kJe16oT4mTUurtA
H9FdUuQi46oTBqyopPIZEyGhKRS7DvSQtPwYZ8P4fY5Ek2UPjcyUwWpliLGYQSdN
ppuos1fDbbGpfQ7kz/OexjKCt8xeYL4jUZ9uIoOYKoIkDyKXrEpe+lRM9ac/XEW6
29teO/lqS0NIC99e0RsX3x/jPtO2QwKOoKeF6u3BEbGBonciXgSoEb+TESEkUyBG
`protect END_PROTECTED
