`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fr88G+NyBX8ll1R4yHXt8yoZdXUxR/jBeJTV0vHPMNodUcflcnM+a6QiYPJ477Ph
seGsrCFq0q3J40xl11RUxciIxCpwmWdnOLVLx1D9755SLqQzdvR/rlmmP32+m7Lp
Nt6ra2wy6wG/kSCiS88vkFxDkqM/f7flbnDGKK0rpZnLoQ4Oi0w0o1eVZ1wsyKEw
ilSs112HZAsgpnxmTVz92fU62Cq3pZCfwsM0e1G30BgzvPwH4tHzs9AL13VPovao
HkmFa6RlKLDXcv2Zy2JZ7UcHEoZdZbUJtBge1ehdtuOFGju4/e3nN1dUxuSNxlQ2
/wbu5LWmazw0GtGshQ0r6AI5CMMkWLDtYwXS/PxEdtos0TMpnjAqg+uhYyfHaTCL
hysdgVUz0dbIraZqPZ0x76Qvo+4E9IrXQ9kpL5jg5DyrkxbIeAovz87hKboSaJKb
ReKqF16XENBybWWwT1JWsXNYTtdgexRR1mYYBNv+qyPnedbJd6ThDbu0+5LfEvJf
uU25hwfFR/cDuez9yCptRqqF08xXseCzUu8UCugTR2lywJKzd7bOdSRK3ypQTR6A
PgWuiBW3DMHT0m0kVNJlXi3vctJTpeLXJ8kRzzvkaMV/jicv4cSVnp8NyaeoJa6U
UbipCynJwLFuNPR++B4p0+guRQICEwqwEES1XIUEg0wehOuZEuot/G6JbeiiBi5u
TwfA9fIuPLxqrFPYF1ByL8/uURgMPwX0qABjw5yUwegJRt7xAwU1+NMU1L07NVcR
wQjP5usmMIBXSawoZGCler1i8XCKPmW2xU+X8PG8UI2dgu8mBSuorWJaNrCgtk7k
Q2s4Cyx087ApMk8hVDfAQSsCmbe9uL5NI13pgVDcOYBA3blX0DdxwJBgPOs4h6Ig
w/nZUjb0bWbF81ZP9dRJkHKddrj9Wv5RHRXgnIoYIgikkUGhT0eHpZ0tB3lDOQZc
U8TCE9o7zUzceKJqvdXCnXCCGiKJ65xyg66UrSyxKCeAcBP+IKO40nVcoRIERgJZ
MZSPk9nb6qJMP9nBkqm2PRZY255ykBy+ey/iCk86MGQpHbdzSP5sOmExkPJOwdD2
efXO24Ulk14ocP/XCG0x1iaihV4o9DnWl102zfJ9ta2lcDPsHkQwCZa+mSUn5k8M
I45487nc6y7Qokc6Q5coVkM5AIMiwjtOG4vHbnnxJsNgMQqEG3GC8aAUsYQARXuE
Zdq8v9tp4Yu+gRBCHCXq374BVzeSatgfDVXHiuAxBwYTWI+Zy+OWYbc675c4qSUP
R7mNx4jKF1c/dKtw4r8xHI7nF2t9Ev/2gn52YtUiN342noB6FLZatDEacpq5TT1B
gAt7d/F+O7PdtDZroD7TkM8ULCLBqeF8L2k3mY1J/PK3QUCFCHP3sKO0IfXsr7LV
6EE0IW6G7ke95WDXAKZhO4VHRkkfL/2BYHUxHTQKNOoavDgu27Mrv98dH8tBJQVs
Y3ZnVsuGv/uUwrRGRchv4M2uiH48/5YjS+DsHyz3vHgkHQH44nzcRJnD8P19qaUD
egrjaPa+6VgHsVxIZDBNd1H86lXjOoXIRGqjJ7VXyWGZH1chR01ShSs+c3akoFS7
xtjqXXIeXC4dJ6WU0TkHk4+AGNZwM/Bnd7fmiqKmtoifVj8Ka8GPDxeAqPp8186U
tKchUygrXTBwei61nrasELsECA8m2smq3Lv0wNNcKBdptLbpRdNJESkpgWy5wTUR
C+l8B1TKLVHKVXUJjzCx/t+WDAClWAubywie4wMqZ8s=
`protect END_PROTECTED
