`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W1kGwQ0wcaBQezQx9kx8Sn09HVsv8/bisN1VGkBD31OYyAXIP3wIINSc860vd1ou
jjysYLJGoiGICDgmzE5dMLIJRkMHjozpbc4RRF1CytfkBViYSO1T8mC3G+QhMGSS
CXHa7yV5ZEnRrnwUPgA7g7+lgypvsHodqb55a3vf7lhRujyEoT/bAIJLnZcQknZF
20hKCf/YgnK6i3N98lReWiuZNkp9EwtMtXrIBPNNQtaQH9TwSxw/Nv2wVSYu7KdH
BVHXAzNn0Mnm6TxB3Ic6kSDzQ2L1qeRyIg3RINUpFKb6NPq1EOdGkNtTzpTLV/3Z
ZOPosF4hJoyvvpEKckKbkrp+Bw7KxqKHMaUYyGrulxLfBrFMPbzOPv6oIcyuZkz8
KVGawncBiDofc1WmLGqtwGPNQ1X5KbtS+NuHGYD4OAk1h6RF8uI8YYU//en4hFgK
qVZ3dHIFAVFDQrGbBd6EnjW2HwnJsGigav1RaSYG0jHvN1k85Mf5Jx3krn56OM46
d6nOClmQAalvxcjZ2xsEwBgh5DSfjgW7bMarwkJ7msOX/qSIN9IEIN06GXdS2gV8
`protect END_PROTECTED
