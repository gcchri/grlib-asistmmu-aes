`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T3JsEcoHQO3XFNkJHwzBEJkidO3RQ+k7Clm0Xb2RDyDqHt0XmpDLF8UAZPlYkNSE
+m4fazkc6HM1vA156Ut6jmnX9hCLUK7fK1uApLBB4sKOhniYRHoxGF9s2iJYM7KI
zhH9V5/L+TllzJ5aONFFe+tLYyL8v3YC86iw6qGA96sjmwRZQuUOn1UdvMhuJgOc
LL+RuXRB4MJjsz5e5wi7rMUIctenyEmC+WCWLGFPRyQkvRhHvSJ1cwY1qKb6MELA
N/ewlxGlAa9EmAU5ITiMnSC67vH6f7GsDFG8kkL1V7RlCWSLPellXKaU+PwAM1Ep
8R5VO50wiQAVKhDB0WZXcHL1wEAwzLEF6GqFIwa+iDyVy/Rs9zNdoPvpcnofCF3M
8gUVggNm5WA8cf6nQJo242Th7ZFZ85u/Qdwo0hDzEIIoJkaGJMtOv//uVKtZHR11
nqwZ/fxuAfG0UBF0RxqtPMto7UTPX07hsAeo9dkuq/k=
`protect END_PROTECTED
