`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SaM3EJN1lCEvpYLMlFarSswUJwPUBUJIUsT81dt4C42VaWx878KqXOjqFngp7prq
hscAv+Y6Z0RQs+jIzysRA4XRgruuChUmiF1ghAx6zgb3/8NI+QL3OTlcbaWgQ+0U
XjbsVJnOYFPzq/gy+EZipcMxJM0bz+/3kcV1sX1+0riHzKkczM0OgDUGru9bvz3o
s3xQmNCZdavPaP+ipqZMv2IoGlFZEssw5CMRyNRFQQL8b1o1b8whA6mwv9ah3SnU
Uqrg2Zpfem/nUhTYQz/2ZA==
`protect END_PROTECTED
