`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ncdMgeAH/z90hkazCpJTcWrc+GbrVGgRbcvDjDG0iFAKEnmtYu/9FYVxo+2VrhI1
necl1CdbF3nm0kgvRgDYZ//s5TMHOI5MduxSWd7Fz3ZT3qe65vb51nUJFi3aUeT8
QICIT8sq6d0S2Vg13W97yU6mZruXQBBKeyQAkm2bV2Q1b0Z7SQ3/Yg+A9uEVQLOP
85i9QtQ1f5JTHqIwUKhIbpkctfnxLNJ/STI40vUXYVLlsbh9HXeSf6m7Gf9d6Pg8
DlQmd1hKgr6DcG7b0wm5TUFIkZ71Mko7iuQ19kTk3FkV4R7a7dkiGHsa5eWbJ39t
ahLVf5UPfEHCt4OlUfqwlswyxiTFTIBAgobcZYo+jmLZmDBuKiwxXY3zRZs3ftKc
h53/2p2Wtle+oMuADTJA5tWHkccIqXxpHRfrwRcFNPDa5PZKT7FbMpwOmDS77HyJ
vPILLoMxnDCuuEAtLmksRK44oJ1WGKgFF5ox43Tml9uo1kGIDXGp7Bmy0nHg7aFK
FUKwFRByAJV/iiJGoItRbCwvgntz94cBlquU+fluUsOAgfL5z3R+NtXwHuSsvb5D
DNMDM0GC9N5Csv8yBSao0yQDXRc0jd6rD1hfIKG7dFbYPPFnpsawmnw7wt5uSc79
1gRZJ0M4QIAtur2piFVEl5peFM5wSUyP6ZV1jQ3iA6F7aVjZ77LhNwhtYWtH2+PA
SV7kZXcAQJMf8P1dDLBUcVkUvFoC2dE58SWaSCxbRZknDGOxk/Xks3TBEQSb9to2
ocmdfS/2yAnulmUtkVYmEIANbdHLt3p0R5Aj/NOR2bMnjDnceH/Q4l5f3yB859Ne
Q0DUEUEuDf19zGFaIrp6s6PO+fHgpV3gr3IRsFIk8q8iorMUtXkaJRpxlIBul1Ln
UocREKSRiuxGaCSfLhl3tSYDTEN8+5LotbRUsuZh8oMmipM9L7lAKCzwHzGem8Ly
es5GmtM9Qof8FBeWa8rY5IloagFLccmIzgkaI4WIAhm/+QmRoQD/ktA1TyQORnXK
TvCzFl06UiLytFxLF1lcWuTX4F+YKycMdm+QSS3ccn65PE0LUBw4owvfmL26v1KC
JdDdad9jMwVT9nUI6nLUOvaf9VcmFkR8vVR+hm3D47u+ovgTCOpqXKfn4TOgKWvJ
JA3OY2neHtaFBpsQa7M/PjCTZPIll0PDdtOEsVnGe+hut3clqFDR0GUIQVS7fKW7
CY2DmZfcmxBzo8+wy1pXE3bl4YGzTdzN+NwWpklxxbluJScP0c5sfyN1iyfZPCag
ID5dnmBnq6/i9hclKQpYOkSxWNh3+QafflurWiMB7137nlqX+0pmoR+gScL7H5Co
jsn63eD8TWAqZarWUNlRvmF0KDmJBs5wB4cDvXCNPKfWtsWdo0jPdHUfE7JvXuxu
SwtvmtH1Cs3qKE+O21gbFUX5Wpis9mIYF14//WpdHLxzMiALIXe866wnk0TCGC0D
eTdhzMFSsBodFJ8qrRxelc5K22VkXLUjCRLuObaXsjpE9BcVKH8U8vmVcKzQeOjL
ujbuhtyMSM76+AgNjuB/7+QLd3YW8ToJRx+Q6EuKH7zWPfevQfmuvBkvZeKn/a8v
IPBDb6j1ZVeHtOxNoFAoZ3GCPWTOz29RSAJBOiZLw70DL3/f3kZ2ju7X6JMyiS+K
1+Nekp6tLid7qR1BAm/3ZVBt51tQKCFIAmJvTlnXljsNbYJUUZfd+N0T99gTi8JV
Ju+37/vPDryYhmYAjGgKCiCJfim+rtkjhUONgsafDkQf73DyuvZyvQ6u1IP0KPMh
h8IrupIWlpPVrpaBlcGGH9MdCzCyyL/f1EvUWVykT03jFE1djheCpmvCE6L+vnYZ
0T4zLtuhw9lFd0TXMyUwypNxojkPnsPG8JTwRT4hSUgfoE9Ue/iZLfSd740gGD9p
1aQ15ydqPkieJSi+NbUnWmHMZxust8Pk5oqICaPTC85vRgRl/1E/qKCdszLelYnm
emzD8wtw0AL/0knaYkdwd88YMmu+08cy6LdnKlMzg2IP3c85ZtPSPYDN5PfhQANg
xHMpXGMFGWYxQRuwintTsVwLacy8R6EYB0DTwXOzUaWwi5cVluJoJwxaCnjVGkDT
XkIuNpfSAcsLNtT/HZtYJW5GQagUpqECpqe+rQ+GnpfaAB9bcVsUIFWp2kHmC/xA
Qf+MKNO+I5cpwaPhedxwuDyKPJHaspsPOwK6gYJ7buGNnDSpCCKC5lWvqEFNBPJS
y2iS5umyUQoq78kE8FBHKzg+/KKTCJ1db/HdX7pc7bekpqi7NN8N8kWWLgyZdCrh
SICk/OeZdKefzF15N1fxx197JQEo82abXXymTBcgJrQ/8Dm+TkFkl81VHsoRR7Sn
vpWQZuSnXA8QogMVnn4Lrnb67Wza3vwON9g28iUNQXkGVp3jnsSQ9mUJfiOIQaZe
wuLdwHHnzdwd/BR9kRYptUETI7p4ZhsCsfkvWVS7dwTQu4jpIsvJ8l7gyu3/BbCg
Ya0tCa79ekLP0SFK23ce/AiwwAk9ttPJTWYNYe7HRndQMXP3utvX9IhxQOVPevxj
+94Yd2AGiD/g7kfbjsuGYNubiN6R3dzrSqBb/4BEWhEhUgMR+1ob0VlwxyJ0p7S8
XmHx5dzXJeWIKuVe5KfAOvaPDKZ5U8QyRNTi073pLs8dEybpk/lS1nFCyiFOorYH
dMDVc3GEX01LaNCO8bnD5x1UgwGRrO0m5ac46o/gdFISfHuv8pkapYoYxW+EgG5V
OgG5blnJ/dKgyA6dkZRu3XNDdv+5ecaL7n5THO39PYzUuucIUSZ13xjKPiqKXsFd
CJ5dISKZqg8N+N0n7VFN1LvgaQ0pPO5XD6CVXPylNlXIoSD6xp51AfpH0E9+wt49
QoUG2b9CK5+xSF19ajnjCK2lEO5Me1mw2mjRSo9EykhHTgbycWY5DG6lITKrMvm7
JlIBxHEY05lY1pS6hZDkQPk80mfXYrahzVCRcN4x4t3g3RsfF0qdCS5q2+WSPPzT
ybmUIyKCEGLjgFf7LwY7h6CTOQaITJ8t7mbb9Bac02qRIJPNWDEUQylrYh6Micnv
1JI57i3r4fZXLmS625QHvE2zem0U2vNqcme70GHd7kyJsZEHN++QNc1K9UFwdXwx
50SFIojwYNPUO6DEG7RmOfaHCl3yJo6i4LasYB8GsHbtBSlpuPJzod3rrll/lCJh
9o2VuxJALVQ56AZ1CHWpCh0oatROtZXjDAhRjE+SkX7DgWJDCy5HTFhVx5a6asa7
48pTLsfYrd0iNZpE/6DCA6kX9pi0zpDtgpVsgu4xP8UMaS12kkkmZDNQTy8zXLRz
TPkItjtE1/OZDsTBdZbLKb5pb64AR5N0ZmK8O6z62fqsgt0UJ19dAzCi4VSGCOYi
D2+C/Sxff8CIRRppuzLwW8P5UMiQjXtAcT2s17QRTmoJkab1wa7RF27F7LTI/Zre
fWQvK3AFrgDYRxq7t4y47wK7hIsC2LMN4wEIFbHmCk2ToqOJ4y5C2Mwlh3ya8W0p
gcPdMterWxRvwSvBJOCABD44GmUCAh3GIhD0h1pI2qmDxMa/JHGDarpNWjLoi1OO
WqTkyN14qc+3kW/jjXWvSG/Ckw0luo5uqcxuGX5ZN8KhsJdFtdSMABZ9Rob3WqIm
/VH2RbynbjKdwQOnRl+XW1+SsdvqtsaAm4nyMo6SrvjPwix5dMwirh0ozESu1t/G
4GDRCN3+yi3gQ935AgupeD+wAKskMZOcxMbUugFohZJKfCJLqodPMtN70YLYGkIO
ResdaAtDm0VPEVNDHPxAFJ02uukmxz+Em7oigMdN+YE3bbbgLAwbZ3hmfpkglqxJ
CFtxA2OeHtwc4Ry5Hgva5y7hvFmnmNcU75aMPQfdnZLztDgMkUy9VOuAi7oSTz+i
MEL7QiHHmwmRmQZaqiGD6e/xriC9XghU3pg2JBoE1iO/t0kvwWM31evKUasVmO8w
JVLdJbkzBxiCaVlLBq24ayhS4IgjATksGdZK2NrUO+9zFeZX93yt6ykDmpQhtQqK
gfCrC7nFDy3i0CN9xUG5wy3MeM1Gg59LfJoQMbZl5/blTeFG6mN+NItrXt3rJ6S8
guv0sL/0UPh4oGg37PNCHR5BSmZ9wHgZC81TRcN2KhdNXPySP08VXJ05prz4p+XR
CZyacjIF1AotcWnb/V+iOgbgy+cBKEJuaNqVWxn6owdmo5mIxOXKACeXh4oodNPk
AAgXAeDHkqapUS+nrvEb8IccABLxTZivWalPDLzArokWLJqZ8LMuvXCWVA1E5MqE
b2LaDKv3NB8WhU8aMqNw6SuiFgmRTuFO4ZAuQW1n1oWqTn1wcebctm/7sufCIJmA
6JmfQvvh5aW6S5vqlDUGuKI12TAAiPic/9GULavKzuI07973wsI9jp0c2MObzPQe
0dT4d/jfgXSH7uzgSVpHjiBoxhq8nuUK9LflhcrS7YIacele4PGdK4oi6uwUCRqF
/IzYLcT9Zt2xtndp65r87CVIOIG1HCOLkfwDJRjKFxmjN5YjesbgHWkYcZACwj/f
20fVjcdvxA6/u+HyttFakK2CpTAfTx40rBZyh6lcMx3b03rQScBlK8QWLn+J5COx
WcCgK8pyY78n6IFEiDydej2WxNxZI1viUqwq3rZqxR9i1sd9TQgoHYU/Cy0MEZuY
Bsyeyrcnh4qMzhBN5Rwj/ZtDV/UeZV78z76LW7w5+51NIOgig6Kn4hJ1EiPujR1W
x5f0i91f4oLGyGjN8QW0RTfxlUa2IGQKRal3obQPmat+UsnOvbdAQPsQewqr/9FO
LdEdOKagVlv0mb5YyYhTc6RUNY+22vwdBt4CbnrMpWetk04JIy1++rGoysQg63lG
ZiH6JX80IXh/WSHqs02ui6rPCI3pOt6izP7TZrgfW6JogT8+OOekPI3TTfLDJB6j
YNUjBoybTPWZxU97cxO47xPHFqEk3Ribbug0rqy+6VyNoiNKTY0xUiUZc84CHVeX
UJxAZYM1r9vgOk7q7LcgPs4YHNyqDbo6qYFKCVVAuy5g8rg1RHHe6BF/J7t8Vei3
GsNWAGDe9kPLiCFgShAgRdIA+8EQbFtEn9ytY+X3mJxFmCZP6XPLkefo/E8UnrP8
GSD0jHwjAfjmaE7dc15HbjQnFY8W2Ac7TO+C4u7c64QcrofDusd5T32djuCGN5DX
YhCIGhrb2ifALYd8WPjOAtkRi9SYH5fE9ogpwb7FiDuSh/P2ADZX5pyvN4z9mJ8a
1TPgZDVHWL9FGkqDr8EJ5De5XaukCpPIyu+gTeptxip24NfdhmISh4rmeD6rAco7
SqN3N9nyI6uOHUYxA2+BFfT2mE2iD4ZdkQclANbGuBaxrXbYdR5200uf//YW+G2B
RhOtVXnMKBcTLTZkgf2tl0TWpifmsEjMRN5aLjOKxX1oeJoQ8qnE46DOhF/rWrDg
doeKT5smctSsQss/yT76WHjYv90NAhRRVuKuwshT/bdbWePWoaxlRKFElCPw3B3W
jtL7vfryTbojyDrnFNPgqpSliRu1fay/57IUn98JXd2kovGy9gyUHG9OmVQdonM+
XpQF9272Qa2Y33z2Eo8gLoiDOQtrmkoP6mcqHhi2/RP++HVqZoO8czwaR9Wz9YoQ
aMQL0SG5LNaPbgX5hctB0sjkamsWamWYPJv+snaxJiQ5m/mBAY/QMVf/FYF7q01u
eYuolENmtMGAigdyI3PN9u/WRI96S8Gnh1614TqlqKmnVixolsL6XjDqiHSMw5OD
DV3o+N0GXKForJRfWD1KTpWMjaEEIqGC/XI68aMXiPfG65MP2c3L+eax85wHJjD7
kVTHCgHXpcZW1nXQps74i/ANlbF9CNSgNDWy10E2GxrBr5TU3MvC2Si5sIuXJjNc
h6AziDLbI8gIJAfu6Am/0zWW3r416fS4/oPge3VzRpFwOFR+uGBm+WbLdb6fSqX7
5jdSGVAQYiIE0q1HVN/IcH3lNt272ontJxyeD5F4P7ZCKxZHl6Em8ASdvW/ktYLK
UaODKWDfaVGSLvdzuO8ugLVg2VzFabLFtyZ3socauacRlZFh0qokWqwbcPeIa60W
NKscgYXmnT32a/X3ekbw1wy0kN9JSfMTyMK7C/2ZCyR1pjcUDI6Qp+h5X42VS9Ke
rdF+BViOLFta0Rkh19nJiEKBjq3H6CQaRwnRFLKAbzU9nTToZANn5ImGPXoi27d4
1D03jjL63H7hJKuKAW182fSBLeTq68oJLaK+FRvmSXT0ScLhgJz+B7o1duhw2nBH
sq4mWTr4Mhf8UavgVZGwHT47ng/swq9v+a2t9TPU7j5QeRRJXY8B4eUIQm37DsK5
yKaPjRF6QMp/rXthy49CRcFvC+rMQIDyCMs6sFfmBZ5dIJwkyf5/aGHQ65C4WHzh
J2ZCOKomIP+MrqonBSievQQI2y5ygbn7CqsWhrptkgJXyVY/eVuLbLMibgnH47Db
9oricI7piG1WxyPnX62gM/84dll5P+TKYhys+x6a5maesNNvYRxd/ChrCj3lJROg
CvqtxCn5MbAUgvQdVLjiImhgbwikgOFxgTsN4QERAvY3cWV7JP/VJ6QDJYpjNZzv
eBGJNQQemGxl0xmsh/1vBVv+JYcFe4QbgvD/fh/CCjzorglnI9gEYQrTE4tUDIZB
CN/f2Ow/g0Hccv856dct8GxpvEz2q0GC/UNgmO3ifQc1ihbJIwSyITu07iELm/Ya
f81MXp0efpbRctMLFfSDgzKvQW5ukyN/NXRMivnEb3Dh4SSbNqsC79D6PamAoG85
Jx89Lf+VGahkcSki+uG8yftzgC8HF11nU83miV7q/MmRffF9TNksa0h+7ZBMEhKk
PTcPG9R5YP1aX5N3YZf8LDspiY5/T9jfE7bR03bF1X0zLE0WlAh6YL4kLpRtW6Oe
brapoiM+wyALnTaBwtDHff0XseVbXGmwnqXb7s25Lc+eUsSWZscNpbC6otAXT1+t
Kl0bJvhTt7O4VY+uFDplZMgqvQRbJ7kFep7gvlHOj5zC0CNSdp7XX+h6t8UxQrN9
fZN3WGR4Qkh15/L4M1JhrxGQc3rfUQRurVMuL6Ea1nmhguer1FNoCc1pw8PvM9YB
ocLK4R96SO6o7F3c/XYAfyc2o/miymfknxIGK0wCGL5sIIDvgtooybigJ5clL3xy
uz6Sd3j4gfLHPeZ41NvukMn1tHU39qqE1UoNfu5ICiV9B8x9UZ/UAOREV3gYhDKJ
HvahLiwCpxCrpPpzqcg6ODwMKjCM7rBmUvI7ApA4ZW/QUpubP+OdFqDMhd8C3l9q
PRY+XKIcvDBt7CfPkrbqvEbxYFYiiQ/YDuDLbGIGetqQ56OzJvhiXi7dmlCPN9S5
qIhgAWu8aC6UXydwhWYfc0yXQsbtpHj7hbPiajbvQmwLWYJ6P/AvWPcSz9inSQHf
Kxx1W8ttrT+srDTRtHIEgKJp+b8n/J1pScOq7PfvqJiKmIRxc7NGaldc01H6uYX3
Ojl/iIOjdHIjPXpdleoIsipSKvactOGJooNpAo5N/r6Y+zIfjlNKL3TLmnewEBCz
u6k9NZAnesWnTVC9L8qSH+y1kSZ8GcR+QWtUjUHa8eIE/kzsrnj9ZHCoewosFkSi
3e3tnBo+pyhch0b5kfBsNh15OCmdFm6eJ4FDbrAGOkxD/ri3JdOWlnMRfalF0xP4
bUu4tQMFcls6rspYQNIBxgL45gSf/Gr/OOh386yX7zYK1EqzLE+wA4avDrv8fmMN
bCkPYovM0Ky493S1vcqdtPiMwLPrYN8wv72zr+7C3BoQiM9I34f6jswbFj4xufNX
ye1kt/fyjQE7Ttwsy6r0f5upfFYxOANKgHpbVWCBAhzp03sPjtK08tzxnZ8WUGAL
uFsC6fyTH+DZQYskDbsghhX+Fgkzj4FS1DCfsMsEiTjyZbhTSWv2L/Rb65IuGILG
+VXinkp7ewv585Nka66jzY2sqjrCsjymOJWT88u711vnxa7vbEGCus9UgmvAEvLe
/FEJ/mNJ/NsJojM3zZ2ZhldtU9JEHmp0qCx1PNBOG3sKExzeEa4J1A0RAefnswU1
vSi3WSvV7aNh9Bioq/1G+9RlMSdqXnRMCYGuUY9jFr7wFloiquDbUveXXNZVbDwK
UfEKE4HwGsmXZISC4rkXd6UlH8c5pXWcnzWnsmO1oQ485g847FRzK6ecJBLxcKAB
C09obK+Le5wlRkK2ZWcycWjQzWN0I9WFpuh1Nghq5gxe98V6T+Y0X246WT3SFJIT
Kh63GeDssbmQBbL7BEGV1qo8O+9DWbH2vKhwU13k+RPAozN6qzaLtcOmQvc/csYk
Hc8ueKH1nWILmX1nf5fcdj9YsUToBFPYX6WWwnYHZg4DWARoUbIDPUdmgrbf4JZ/
S55yQBPUwKj9MSrkPoYQ6IElGNReCXJVYH33Vv1PsSSjn6i0DdPjGBdeSiuy1som
wGns9wsD8NFSEXIiOyeGqyg1+nPsxM0oyB9VN2qVK/6PijdoHmAo2tVbTBfn/LjS
d/AMV8KxfYXIYDYBxSV4s8Ls+l5C5UbJjAe8X0IBhSLqisWv/YUWqcsR77Q6kDod
iYG4RZcisV6r2EGYQh4SflOiJUDPvMkCmi3SAHxnLpvarLAT3XNQIWqeziKo2HDs
v4ZX+qTzEpu8kG3woC3ouwdjow92ZW7rvMns8TJ0i8Q9VPmS1VrHqnBhBtSllgUR
aGNHQ1bysp+ZQxO0Z7M/WRjk0zir3iZd/h6KAf4N+WmIM1XEg0rf1lhpv4y3UWFC
ABZSlagm+Q/NoxjCy6PPGHE+tsUSCiq+dI+smszOVWBZy6rJJK3VXgPNKLJY+OK6
TyoHUsBnBpKdCdb9cclaoZVVqK3JuFlFTdQtFOssEZE/rSkjG2eEzNOe5DTdMRg0
7BoB85/T1Z1BkCsjaDnceBwGIik5epvloHELhfDMMt3uuTyMHrA0ji33aVLXEDqV
Y74rYq/AimwRKYX+xvVJABb6yV12eez4K/fYlzFHe6DxeBGYNwaPWIw0akrcx7LP
B3QzFne9DoGQAASiKeA67ACs6Nt37NxCaDiGhoGyaQYIY4EQ6ZZPx1YHXo5PyHuQ
VaolqMBJ74h2VNMN4IWgKIjnW2ipUFaDQgr++hQJQQoDS7lPt8i68s23vjBagqB8
MfqE4OC3fih83AiM25vNAWrvLGGK1mWN0r/8guedABYL7m/K1EYNlnYJ0+Mgj24R
CL5gj5yTl8qBDUelKxIOtVUsh9XpZN4HR2iLRilcNCGjcgqZFd9GQL21+DTofKVD
r+AhlTAGe++GAk89EQXfTA==
`protect END_PROTECTED
