`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sAR+/DYrblnEI/WbEno83uUkx8wzxGCi2cL5yvbI4DaK1q9IhQe3BU2IhwB8UGkr
hyoK5M6BQgNbImTQZiKZwFgGsM/iHVgWPH7F3ijBnngg3E1OgVIqEOuUK3OvBIMT
0c+ZUrDYlIlRKQbtwnYCDdwNtSTEf3+r+Zgf0BtWhKBV3597Xtdb2zX5IRXim7S4
DjUe3Xq3uYuMhUd9iVPe581k+BBG+3BfsnetnlNxjmP+tK8KCgg9BtvoPXoSHN5d
d8cu8TN/+MoQLjsIxCzhare0zwXzvGDGd47vhYa2kxPS4YYeK/XwbFjh6mVEtqN/
IrsYiMlEVSkskRrHhZNTkSur3WRp0tpbIaBpMGkKbenNVd/Av4cra4oS2hoANK4z
1qef+h0iYbE6a+kE5AQc40+aNs0Bw82sG1JsxHS8uvHQEiz0XaCMyZgMcguW1i4f
PhZCRs8XRl+Nq9XvsIOAQSYwDmnz9ffqNRRMwLpL0Avqr+nk64Jl96F5EXIV45Jt
2iCsYnkhW8S4ANJO9NPvBD8+09OFwfH32GXXK/LppApq/F6rKWGMKy67bKiGtr5i
xUbYHd1GQksvaNq4EM/K4GlqZe6siGXV72H6ThUubIhGsTUWj3+n/EqowHVjUGxI
4VmNZc96WNCuUwo55ytjS45jpf48VdpNazA16y9+rzUVIocfAuwBQ2Uhl0EtGX3/
2DxMkch2rgShPVa4BcifWg==
`protect END_PROTECTED
