`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c9PuJLRF4UYHG547b0tHtTscfepKJyu0qtCAtNZi3qQ8Jvbhh8LuJvBkPxWYN7Bj
i2I+HVh7LQzBdoc7MyzeVkiiJ0IqlgnF1nY2Y7TUMrV0oZ/ydCQaBj2v3BKsNgB6
TTOEniZpUt7+bBf8Ekapp7BlnkIh/DMfqT5xlRVkCAPJmfK1gAfcP2u1EsrMYPo6
lCzRcjhAqNsiqhAN556I4obsIHAHxYMmAFxozWKUXJj4iYALQLzdqfDh+tIgETSr
eXX09FRiB68Hn33ftrsE0t3BPruempyCoMtu1uRRP6lQv6WqUIOJdxzlrz3+PxVy
gPt+FE8Mrnx6n1ZHm9EFgaW3/RGkJUIgfHOj5z3bIPE+5YlDM1X3HqVT0IM5t3JT
aDJ+AsKPvtiS63rPM87evWm5JrRIZCswPaC5KXmUnI8IWgo1pE3Ohs8jxdIZWhi2
+4VJG5gwy4RNWuqVNrYSphJkFzX+PG2TwFywTNdqJPA=
`protect END_PROTECTED
