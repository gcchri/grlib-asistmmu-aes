`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fX9QUv2qGthbKfJIJ0Bg3u8OzUHIE1u5oGZeRkT5n3m8Enm3nu4JJydRevnDvWex
hW6v9jlMMavbC2yW1JQm117u2AGA6au2yfu4DK4Ra6etv6Yn3EdsikgR1vwqDJrp
PFh5YMp8+YDt6LlwOT66CVug9X7OzgWWmUS/ZykwvcUX6xzCGdjd7EtrOdCXYU5Y
vMApLb7X2db4LnZ8lWTyF1DBp/td20+ctHlMUtMYvWihC3qQDoS2W4v6NsfDRjsA
B1n62N3iNdOfnLiIW68mbmCPWRkksdN3A9STpaMYbiP0xHTNjX5mrpC2GfJfjQn5
woIanNxY9p07X4iVyOMNq/bsIdwwRNMjCR9FT4rXmCcn6MMMZwhEWpMgWaPOAaYf
BAkrpFEWaP5eWYs7bYkFR42YA8VefnPBJLcKTpMYpOI=
`protect END_PROTECTED
