`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PuE8LtN467zVrz1CDeNYvPK8UmLxbkMb1zhcHeg0sH4ncnCLoqVyF9HNVyIodq6M
oZ6NE+aVbNrbL35m5NvpFT+5kQUUnlYa3ET9orLRxzkDB1SyIjE1dYtTb4mBA53n
LGdH21/uYCPg8vkrrh65bnvKXtlyDhT+FOouMPOdt0OxaeBUAqFBRHrgHh2TBrve
4lhdLfY/rrgQsUMwgELwUXzJPQGuWtcPEkywjD7hkQfsuH5qpLPH86TNPnRee1L9
3XPY6GL5F45k2xKgz2Q7nSg2kf72XCGviOR8ZdhcwiJeo9d1lOmU1TbKY7PT1J24
aTIEojAt/67sRI0TFQcKZBk2w5cxwFQ1ZBl+WAyS5u9+t+N2xwok8OyxgbXQn5SF
+BXzbdTVhVkx0h6Qv53lbqfWT4f+hEbzdFePxd9jNhYqqzi/+UQ+PdKUI2CjFgmN
p+cXtTYzElJeubrjU2wGoQYpfTX/You9P6rhS66q1zR4fEOU+FRYnw1GUt1aBAX2
`protect END_PROTECTED
