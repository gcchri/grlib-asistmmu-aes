`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4NjGpI+sZ0Iimqd27iuoGLPNTMePmn3aF0AI75/sul4hXg3C4+90DmurANTzOwKU
zHK21dyEJGCnseJJXchwo0h8P77tlW5ICh5O2ueKVqdSejrq86TSfr0taMRsWWIh
gvxafXh55vgEm+fwZOZKmYrSY5PKZDSKY+mx/CF5GrDzi+xn+poSJgbWL7gXPSAS
RQgCAON93VEmD2wgAtkBsdcpcfmrsPaaZ2ww78iKEa+Dx//u1jTugscwBCGpz52u
FP+uB+Fw1WIWUycBWIkifMdf9Rg9f+/cnziM1r6DxELZ48JSV/DtKHAXiyVISwXk
vTBAXuthyclTWommLoWQWbtlo/oUxb23YHOKJO2uNoqgmRZuJpLNDWQIL2AFHqIf
wHtVerCYeGbgeatXY681wjrao2ASADNEIyLc8YuPUqHfemum5krwNghLjH4O46Q8
DlTirDgMZO4oSz1whrKbRhREXrndLvqvKKSY8WOWV3mg1/x/wzY8kW8s1epx47iW
FONuN6lAKXIUKKKZod3ZUrth2fv/YusF5ZOAXzhJ4fQKSdRN77mmsc0eF6YO67dL
U2x+rI/lXtgEVts/K0aMCCSPwrwdjYGkYxgKohduqwNT9ZvUkteNkZruKY/0X3M9
/MnacmB2pL7PRcmOIl19kDm3AS/Fcokstmfv4+S07x9oXBvQgxsPNxVU6w48kaO3
P6eRhMT9crJ7FSucJPVX+aBktlSWSib2zV9o1hi0y8Zp1jHyBnPyjQvg9XD/KWtq
I0ixtznwIzK/+hNczsz2QuqKA89ElNR4HneLOuxqUE4nnnJwXPhK94b7/Tsk4EOc
geZN8HrfStOZsex4eUGf8Q==
`protect END_PROTECTED
