`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2qT3EMSyyYKzcBV7ZKzn4qqckbt5SDiNrincqTszdeyuwNIB+0attyK6Rq4Rpz/E
/1WW7Yz+acwXMQz6OQ6qcvHexnvzi8A8QSHmGGOZaWgndJGNHBAq3os98tCqhqL5
7Kyd4bIQzB59oJdcuq0EXr0KalCydlbrzh01zWNKCm7t7oII6MS2pXp1OGnvLliN
KgTq2ZDg/ahUR94KiupP3cHplOwOE8f9DnhnXKK/p7d5xgr6DEcpU4ITuQpw4Uy5
B85+2QPF750L4qrcx4heg+vo310kanZ+S8KXvn9vGMFS3UzwsSdW7EWdwgmTHPrS
D5G+uGm6D0JWw3L8aIn902Hluew+J7K/uiQ4ZkhcxzS80U1rTGAS8MTMhcFcxeFP
wvCcdB0Zg8QXCrKAhef6qKixp6ivQitbc4Z8pWg4PrI0yGKQI4QSYMcTRZtO3N1g
uKcDflATOrAZ7hWQ6pAzQxdYAdk4JeCT+gfdlxk/4OuP42ZmpZCz3Re1MHN/J9Qb
N7pqiJ1Y5XK8vetqkr0rK79VQ9WmKatJjAItO+J6nJQo3Y8vtiBLw7p3mG2K/Osz
QJnjwpM/3W5Ptqiko23UR5xivM60vjmyRxumZYd/9SORPHHPp5RYOIB3yCCi0AMM
A5GSiSLuarM/1BPWmen7+1IaGNupQYDyXpcNCzWPi9k=
`protect END_PROTECTED
