`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BSk/S6Bfo+E/CCyBuYAWGZVQcibeyuwP5Mvyn56OBLShI32vz6LmbBMruGTqLiIL
pkbV/rmqtX5K6Kgdsl8fb4MPXym78tUtxh3FMAYQ6VhPYys7Zu2cm4ZEJDp7wWID
eyBOFhaJOB2aREi4AO2AhV+K0z4z9XJSJ2XqamEFPWT+Z9iDh58zYheejRxFc/hr
nYApjYUZU0fjEHgsrjyMUANFoQ2bKWJInQAVrmhgIsCE76PwzJQYxqyqZ3k8fWPc
vjuQb6ayT1psHM355yvJJESVJBTH4dlvdMXYQfVbU7G/4e7UXUh3ynkJ9kqhTePX
R+KGTN3W2/mVF7R5pCG/hjdbzrJSNxjBB6kXJ44Ok0bjBwAFLF0lQJlHspAs4W20
ZPWBcxBm7WHmESwoyASb6Pdgg06HRKevtI9xOCgrzLvyAyG9xfyaJRM8EQHtT1bo
HY/UNO1dpZA1kPzRCtVnhcKkFvkqL2Qgaty6188fqJ2Eze5voM2WSrgIMN/J4tBb
0zjd8nU40jZvSSayUoPj/vNp+xeOKzuKePU4UAK+WuMp9sPw0PczNzlxByF7amhT
Ah6QH7wsYlPFg2YgvlWzOQWaG/gJVUbUmYqfDYRkw6ACMbd6PCHagCly8Jy8c5cS
ZWWxEENSDiaOQT6PZL7dLVS3rDqrhz3IFSWTguxUyHx0c4Zqk5n0w5+CJwdibihu
5mlzTpdw9F1MheR+mWHWe0eBt5ibOrL7oOkXlnW/0pFCmyOPxO2YAbcoBznln1GX
VVdaOXGp1rEUCRERvxTVwNA+n45e7xPXF0jT85YH9rRiFiy4SiN6BoghbZ1AOgHf
ZHE2nFPt3K2W1DCQbUjy3QHm/HJ0S5lTEOh2Pcju25h5pQZZyeEBrC79CuwFiOq9
BXzbjzc6dh/41ie2lLAufYDN3EELzIyqodowtkNPfmw5ioZ+Z5ASTfdEMc5JVTGT
JMPGErOdkhmCHuX2UpOqUu2wn7HWxAXh3F8kCrXuTgiIWThIq11MOC0HcaakmO2X
RVPS554z4iEy0LpPc3egYU6toKL++p74cB3GX+HUUd8cXPcwmr2hJVvYEL1GxB1a
gRVOiLHNFzK2zYd+McNfbMa9Eji+Fw9Lk1Jt3jbTBS9XlIk3gPAkezF0RUigtVhl
y3L76CkyWVWgLmeTrarMpa9lr0jDvitBL1rvd2BipRs=
`protect END_PROTECTED
