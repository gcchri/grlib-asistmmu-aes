`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jh1+twYCW3O+PFNAfZ1+9ZUNOHkmQxWoitm5A+DNzJxGQjBzOjwRMfaaIVknVNfA
Tpxr0XvyetICbagMPrYQDQdj0zSig++U377wbcQYhXJF9Q0hrr5YiBap/8vOEbp6
VLAwm79A/IOEn2X6X5g7hvxdd3hniXGBqNnEIrEsQVB1TUR4dSz7DY0f2gcGFWE6
4YSnbvBibXs+bfAnS9a/cLs9GZhcujjGipSBWes8VHWGP8p1YX9bsB1VWVaaRANd
TC7RygSlWw8cnx780DLgCkG5YJHcf6imPScrum/bIg4DSrc7NcmucqBdU1CqnR8H
juV5SqaZ3is2aFNTMbdJGVA329LAT+1auTSDBMKOAwiLDPgFmgtNbZKCmkTwP4x8
ygZHsDUUFXO6Wf6Vo2dFfeMSRGJRmL8ceCssBVRW5o05vQOAfSA5db1905W4BVWS
bkZ8rn0otry6At0QYm1V0kuu8oi7+/uM68y8X4gzMdc0OFRoksTg26YDoEJc3YEd
EU80GL5wrRC9Hv+o4ToL0WsaP3AUUBonDFgdGqyUPZ+HZUuSw6VWxd6g4geiLiyI
ZLsQpUONtK14rkyJG39uILSqPFaraf5UHaZPy5MzmoJ18XlmkOteotueOtpUTzGq
`protect END_PROTECTED
