`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y1ZEvgO3DwDSa9hirZE8MBz6ApRRUtI2de8Y8fE8qy8RxY3AHDz6uUxiKfU1Mcss
MxIcCIVlxfWNd/pWPuh3/4UdMQkuaa8cHkEbQMUuU71NPal22X/W4Vax/UpgytX/
wd8sSrnMyKeC1gY7K3rrWhz1LcNS9/ZXmxxirSa0wOR39rE8RyHQIlJ3ebGMqhAL
2QPObwfl5U7ZIAUJkGXFHeAyVOYgUcKdkIlQ6VL0UTrnggUoY2lga0u9I0tkPtXs
IdQl6d+5+p6CW0V3+bkRguJThWN4oh3NpU4e4MngW3qavB2W1Qh2k4yV2a15qpDr
`protect END_PROTECTED
