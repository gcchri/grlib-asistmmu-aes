`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3JxQLXAkQ+tqVAPc/O1W+dI0LlsTYGGKm/Y/6j/tF6NSyuCqUHz8cNPFqVnzIOfK
EbyhUF9BSTpoRFQ8IDeEUon8ULB7BECuQqb5Cjv5gxgls5QeuJJVuTyFJIucKPwf
2ZvaiG2KzR3BrKc0RFyhLZYCnEXLnOvLlal0/+DiYiNts31i4B/P+Cr69/86BeSv
wDVsEtaAxGewLQUfOk25aUdamFYAu1deTVitf1aJkCUIc6VX7JwcZV1jTRNfGJMl
+89WP4HShPZlQ03UgosiA7/ByLGaK6IeT09vsdr8XTGw99Bz2tIxGwxwA5jQ6cJ4
tmcFTJ5ONqct6/pJmVbew3iK6WYrL1Ef6WAmaMXCVzNORZNutKM7CarUjZ8/Hp+2
97dCbSm1U9W/Z2OAmw3xwE2zHIily8erzQCOmSMZAhp3cr3OgVQ3VZ0uq6Ff5Cm7
UNqIE8h8pS0/EiEQpjgmRzWMezTaNsOeIn6gnm7iz3fy7IZ7Q8Xz6rbfcUnQjylc
lwDMNEfJ2mA9GjKkY8ohDDbUtvfNqyZoyeUuCC7JECouTzUDbBjRGiwqLWqiatwH
+35LKDPEEzVFUYsvTxlPEbFKaWMcsTNgxEC5uGRebH680BWTwfCso2SJVL2VCMd7
o87tG1WuPtk70j6qrnBkqboGR5p+Jg1YU5f8tMgVCMk481/WN0prCiExM0dWT/zo
/P2mOe1CyghiKhKiXfEMt5yYDtR4Z5xD4L2/QSx8QjzK6JUGsKOTlR31Qiwx5nlH
gY76bzcdqP3r78CMAaXowga71tcfIJ4t8o/ZGMtFXVeylMdWEiEyeYcfdPlhXbZg
nZLsoI8RDOY/F4Dn3ykTBeVXnw9s2D9Rv6zQ33Scxuzah0oiyxMiN9Vi28w8/mcm
c6v7WcRFrwv009AED7zcLB0zbRCYaK6ak7WUbWcP6qrcRJwavSNQQ6mnR4uJ1QI5
KImLm+8IzgoamHTG5fRs/vPO0s9fmKaflMRqopym0CLSu1V8fvnu+LaqkrXkQmJF
BSm11XxBOlQD5yPCSo+4C8nlcyMiIejsL4162z6qG5CfjoBlKzfdSDN5VpFjBZzC
xRhHKQSY6/gTtkkc3oF9T/GNeSBQG26PwDLxgGfKebqn+zGASE1UuHKkp8Ffi9p3
8plRsfN7BjK4yZVkWooAoCvyM2EXjqFxOHiSrDEDnSQqhd++VhPm1zoJ5RrRFCMD
0Rg8YQpm7h7A7/YbTlzN6PH1xtxTV0zd8ORlt4tWw/APNLHEpGDL3CDPSYKiHcVH
YZO7QuM680qJ7A8iDYJ+ADw/ovTHnEhLA7CkOOtURCGx25qU3+gaj7vQ5bPFtFWc
vwQfu6ZBzsYoMmvaeNgKIruveOvGbfsSRUq8Hw+GahtrnRDxBHMB4Cs+bhpepfCe
1cEujZsoBcsSEW7exHGcWdQC+x5/7xScL667aa0UFBqnEKJCSQPomUe9HwVfe9nt
g0AZOC+tYU8jORrA/hIZ+6RhA9OrVPmaWDBLlbpwWb1oSsbn2LxAWk06jmy3MLyB
VjlNoVrE5Oe9BHrtfWtPEyZDE98hlWvW2fTECvhzdDJD3X0zl/K8A+5zEIDwB0i8
zxqz9n6xA4pkRVPICY430pmM73MRQeKEAydCJHJXceIcO/OJ+wwL2z6LFvynGP62
bGwufs9QID47lCPVjoSCWxsqMG8wj3GNQGFVIBtx9FYWNgtsG2HbSLmKYMq7WXIo
HtWu4VUSdCuq1awRsVfI+sMB/mkfjzNGbYFt9bnAS/Tgb5+CHN/X3VosXe2DcENG
afGLs9GJUULd9WQmB0PpnJkklVFsr9/9TLTlDFimrAWNcYKfQLahOCnj+gYXoaqo
Fc+0m/p+EhgZOxfwUQN1FRbIHKiLgO1sfsQYlOS0iKEUH9Byy6vXw83+s66eJIix
KpnE5w+vtdH0pN8PqXUjpQ==
`protect END_PROTECTED
