`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2/hI1o/Ana6bOvt/maLX87KyWpL8yMUg86ddF7uD3kBwtNxNTgAKX8k9UklDPJoT
eGqsoSFGMr0IiqjrEYVjQi8fTKsnvKe2i1/FzFGYT2aUgVqSLYiEuHFY88q/CBGb
cfjEtRaRVgAQqhftINIyIDuvLxvdZ0kPwQ211feRfxvL3oBF27XAUcQpf29k1uxC
chLg8UaACARMzJZ3u0bDhzQOcoUlEVmsRimqBTNRMsuats+xOrINTL5dul3x9rav
V8WAwi8Y4KRY1nwrc+U2+GZvIE9aMeh44HmeB/hM1mLEjwWC2KRSVncMDdv7FAOh
5Hjm5Wywk3tSrNtQZbfbGjmbWIOFAb9gfVGztvTYAAslm9mzN85lK4174O7TAbfb
nMnVcN8VJUT3iERGr+7ygz8CBEpuozF3ioXHnKwm12f8WzhD/wzv3lxJ+Q++IpX2
DgXModrepdz24KopQ7yx73sAAWrXFpV473MhuFTO0HqvfB+GcBh3TVr6mNUxoSf+
21dkwYlDn7vkHWYCyiXADiDvuZhpRRaL0/LIa477p6UvaspyfibVgkmtP4yGd1e5
jwy/Lwal4/ULtC9UHb7KTppp8lOZu5NtuI9GIz5Q/cvMjIHh6NzqDxISB1JgNcY3
DuNNmhCIlAbizA+e5V6VZBm3M0X/85OEN8HSuflpVjjn+4J21MMLQvAFW6S/S1y8
Uofo9Ub45mdeS+GB5FxtMbl0yG3gn++wg5nyQ8y8qLt6S3T7e9sQHE/Ehf3pEy+F
lyE/ZInC7sxSm7PGz4Oh9A9aueBWkSRcoJYeKmlp1tfzbDDRobcVTGBH2VcH8YLb
kD4/B3w3vhoZRXqP9ijNikE95OxqLN6ChGbUaIx1+0nmCth5fISsHWgkozjRUlmI
oomUbu2u+phrUXn+Rz3L4mvOKThanFIGvTL96uxb/L6kerUX+ijI7TF85Bkbt87u
WCHJ1PQPgpECtyJqvF+/cssff5iC/xXjGlJ2MywQqSW+xuiHg41xR7NeIgtoAQ99
AISWvLle5cFnYR/yR6lnUE0zlDVp0aTxd30rQOW2O8dBPNkfuVFViTRDLc1vetak
eC3eTsh0nBN7u5XJibVVTxxiOxXci9/8feXE2jJCWhXSXU8DDF7zg/NaBYPmksAR
XFiTYNvMB9W2xptBT3+RwnMltfiRPeH1BJerynoHuaiHQ1uQBY7n25YvVGEsZVIc
FvjicpGqCi3SjwfydjL0MnXo2xWwku/NRKZvBbv4qMWBmpNIHrZfGernJaCFgFXi
nIzxiqcwy2rIrSJq+PS/oTj/X4BDSm8i9DwW2BKg5gt2kD3KUNV6D1JnQAGUu7c3
4wYhdqYUzCtoGWGvE6tXQO4FW8PohQo3MfDQ+7BtxQRbhoxjoHIusZOa/LPIThlw
YFZTQXEeRCXj1Vz9XbmEmTvGj5Yl1gjmnGp3C/rX2D60O0Wv7WfZIrnsFNVYQaE1
ZJlYucYhAjjNb92FW73KBmh3HOhj9NwL3mcfAOZzhl2jfo+DrJyCVD4U1EXNVQyh
kVV/nOVCVS75AsYRYCju24pmmCH+AgrEiCpjoHpgxt+5R/8UQRnhAwZynmzAgBzl
7dnoCkh1WfZZu66tzOyizDUBv10ETMFVvPogc4y3kG2GoTM2wzpzJ+xiefx/FF6U
fevw6eZyA6V+Iu//YJTFd6qXJfuSEI8BkmB9cNwOFvQ=
`protect END_PROTECTED
