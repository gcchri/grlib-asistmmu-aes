`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JXR8eE7hemrhcnz/Nfqk6e6lXTcYpi+moye0unYMtomcuEIfmGcIBqmfTK37xcAZ
S3kOhtQgVCEIdqndU5IrQPhx1FS8yrMKjCfV6gP6QgFt+3gsbOaPC6cf0+epapjl
Iu6ZT7h31giRYU3wiXTuG5yljQ4Itr5CTMz1LN012XiJNMjIpYaRvR7SgkgBZi66
Wl71y4JVriwKev2wpyIJcfuvWLKTtlLMX2LOx4hgBI8VycVaa86KM1T1zlkOZt8h
YPlZ7S2dt6zT2/Z+sORlRePxhrWo4SG4MN+kDr9c3Qycu0NBdTnZ1uBkrp3ta3CG
iwuHVdlB0krMay4m1qe3bXPyGvbTmToUrr/+j31yON3yn44iPI6e3vRsyF0WZk1Q
+VMIOnLxyqMMsjsU+d8ILA==
`protect END_PROTECTED
