`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HdI7tXTqAuxU5NC48n8uQEVRnFfxVL2UMHRfwqbWmT11xYHHf3rjQWn8ZrxgnKys
p2mcofz1Ztt0wzSXggLVIf0FoTspoMTpUPqtP5HqRLMEUtsPL/JlMztszIkOZ4MU
pAluiSm4ySLPyboFq8vZJhRyW7864cX20A+z5UHsE3VVUqTlzSGPesLN07UCA4/h
cXo+VmO2D2uuF8+VWYofLyJT+VG4Rl5/9rvTr52fuPjZHDC/OmNl5qvp4F6AlkCU
quMolXzoQRYeW59ZulKcBb/Mo6hU6boKBd/9wFLriq7h7wCofILhXZNV+TAVKfbK
jC3xFx+QndOA7nSlea9Lmyw4x9k0y2so/jtWkhwKQUz5eXYgNks9B6/MxeMAdnud
`protect END_PROTECTED
