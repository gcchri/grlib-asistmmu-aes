`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l/tvFBc6Xz3NtNVvmmW3IMiO6B/a2DUmyIyqdmPu3HjqE+LSoN2CxqPGDd+CvNRs
yh/DsG2jQi1Emi5SYL6TD1uDN45hYRJ6dZo2aUXu1tUMSE2Ay7hrG5LJBxGiPyX+
+KtiAvDTMCXqxQvdt4Lbf2gTlO34m9byGEag97xqGRo0xhYNrEs0lwHmq5LZpnBs
+lYq8NH+iWVBqrgDwRhrO26GM0erMlcI+i/yGXu+kZZBRc0QgJFcRXSchvQliN8k
F/syEUnoEb52WrC6bYQHb78dhErs4Yi7TmFJ0w3V2KApuLcdpxfssL3HpaIw0fAP
ODrUYEtg/oSrHZbykXtYUFHeV5TkD2bdQr7zuSYaLlIY3/YwYUwggK9IVL8q10KN
JMx+Xd2gnmelvlzp0E6/ftpD16Uk2U4VvzJYLYn9VlboT5r9UbSE2LWlIAJbjv7S
`protect END_PROTECTED
