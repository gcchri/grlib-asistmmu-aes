`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LjPxmpagoREHH4UQ20z9QY7tlxzNNuIPa6WIfLluNsV/YVgvoL09b67lzr4uFy58
kzPtvKUQDeunlnopHrfGNUKQmBVAg1FjiNTKyC1/Y/jPrqdIPfzMbynxADmAh6nH
U0UIVTi+1fAXtaRoMajn46Nv/nd7zj2JkTTe0uLDZ6sBzF/yiypQybZavK5+8Ugj
txs2WxXN/wvqb1PjQwnUPERvZVaWdBotwYK6S1CYhExW7sU45MuSqmdVr5unPjOp
FC1Uq1VJwVWNtxcnpOEZBmbJWjNevA0dONbpGuaMgYYL5hE7lvXA/UPU4Ge6Nfdb
Jdf2109KmMvLawUm1W3+qVwkaZLaBXAswxAgF9sNt6Dk7cz7gUHh7N30OrQBNigE
69VoLiw7aCStRKOhcEEImV+ZrOPmOgn81MC/8Yb/VDxrjnyOLjJE2W/mpZHYNVYh
nPKuhGPx0NKMmMTfnVM4UzSyjLFK+b3srJb7VF3f3JU=
`protect END_PROTECTED
