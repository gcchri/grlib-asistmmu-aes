`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fwnaoN+pE6lPBZbj45A+IZfvuyJfpo8mCBpecGBLfHW3vVYmXdmxqIh52UYN8Rba
gpu7rEGe4cQAvyj5asQ9139a8rkloNsmx6sNzFPJT1g6ZibbEIhnP+3bY/tU0sff
ibFrWe1EO4NDxi/g3M05YLRTNh/P0JS1iUH67yvdHPago2cNldFVXQPtmHOKOYo5
Nt01tSg4EQ/H+PctpKHRYkkTrQyJ9B5Crau6uxVySAJFR1zKr7rLvS/JAzUUg6oI
daEgKGGBRzFzEuMEcuHbMpetjF9UUJhIxZNLth9dBpu6F5sU3g2FKfqb4zY6KQPp
A225/XKs/t0FL0tSMJGkAcE8sEKJrYyt5CMC8MWrcZDEjYbfy4vVQWKIZo+uVN03
MlAa6XWDZHLQ/2jI/R+zZjYE5X+CHOmiiz/iec2XJtuU6xpwaSuqkssvJTY3FIs2
Jv/oS2aZGnahiYBgTgY+e+M1E5Gyt9WNVuGucmCPqnR/yYL5BonY+/zgXhI3c4kd
ovUc9Alz01aknRnasYOM0+tDkyQEloVoDx+lSXw6XcBv06Mk5uzbYndEqdR8GcL/
g8VqD1tkdfX65YOCQTLjg7vWzne/+AsU/PQWy2KcCgHOWVH24mpFx94E9HpIjXn1
mJ7E9fucBXiaG4/nSedmpO+zoAeLzKwo5EQrkUvNAV7L4OBi8vM24pR877ucrXjJ
3yE48qKTXgQMYcbX5Q9xtpqXU5juYaqtFclbDc3YMVjvKYgrkv8CizWorMby8+Ib
YtBotO9J+7OtR7TaAefpLxTn8Dt4vVNuSe5NfQa8R5ejyZAcUoPNqQI4WO+O39WH
8LM0DImKzefUAMRlg7N+4JMMcqiZnP8Gbzbsj7T+qN6w6lBX7br92iF3WbBknU6E
E9emPCKDgeimot+QOANl2ipwSPK3E9LkuZyjRaFO8mICe+oV5uS+XjIAah55ez1j
8BmEE35mD4wqWoV5T00TWhETe09oJTOMA4Ulxpe/VqneTJpv2EofPq98Gxy/VM/+
LzhiVJHpH/k87XWgiFUpZ84Mh8ujdNBHi5qH7BUMIt79znxOqrb6YwWZiNhijCfO
0H+jldgWSmsdRbXoPpMoDfuZLwVE0aPAOMLCTohfpBUs5IruxHTDQfXSyVnlviF3
i59ubf5kGV2PUcGZPAPIJLPCu7TLv4gglgZGCjlbfwc1Mrzfm9gowwSHhMr3J+Dv
HAEibs9LDxHp0l2lN7rMRzzXySKD0Hxn895PqMvcI+iC0HHgMuHxnLmsWXqYgAaT
yY/awagOJ9bN+wIKr09lE84UuF7Xb2mo3jE6BivJntTTJE9MpyY3C8BsrLfKwklr
OFSu1+MoQ+/eB7n0EN38ZL075vBCQS9u8LMgYxkRviZP2r+t0GgqEl2w4DE5oUir
ZsOrIiT59qnYH9YBdYOcse5ifYazDM5VoPwvIcZDSMFy9HfgXRHHLaZsesTvUt77
OVgNQxuvsOO4OLjl/DP4niPr/JER/AqJHFuwqbWWDBztHEJqkHwg1VcGncOt+aDf
XlB1UxQkbirinYp5NZvNI5kf1N2wWS7YawTHT3juYVjSn/3uzfaDyxFycEhN84nz
x/bsL5yJklDITOLEJvsyLNmjgmhGwU8hyyNkraaZ3qFfmceb3eKp1xQQuzhQKuMw
8gpmwtBiGfWDABbDn4brOCgyrBCCraPqj15DvH0hzyhfCHEtFUUSrAZyuIhWCh5/
spjRMMFKRzMjWAYn93p+7dQ25I6eUSrad4FbKKwgYOdY+6NU1oFdx+l7Ve91xOHA
YPkl518YIwWx3l8zr79BNIZMixjO8W646rcWdMgv064nEJtUdP1r+LBpuSEz1e1F
MAQWhsCuLQM2x6yk9WOBmzBzt3EuAJqIwZfvQwVUA0nDms0+6cELbrfMTIRjSbvO
Cp2Ntq3QAZJo6IUd1PQAqKPqh6oU4KPgJgJGrqvqyNNEKGssTW2YV0ambjyvNCQu
kSlOAbKSeN62iUMHKdrmMre3vwWEMCGGs8PSWd1fjHQKldEJn6yrZaWKi/ZKa1e+
naxqk22z1uJqNiiHM1GtHcS4ET1ueDsrPTO90u5oNoi5+oAy9rpAPQHHV7aOaFYK
ULX4d1fqoeKlU7Z43IF2QhnVqbuDbd2fh+DhYmhSuV1+/zMOQgNagsgh/DJET2KD
+S3PBidKpSZ6lXR0ZJ3/EDGr0mzSqEmURt+Yw+2i2qW6X+ou+KnIcB/MJWHJMP3+
4EqzYV5wOYLpyKeBZcrdfrmvx4kOuFP+8HKQzExXbt+bBJqWW3xFlMKySfAMlJlL
8+2LFL31BN8PY9oYh+wVBrnxygVaIS4RzcuQJ210QxkkFxTEhKJTMy9BxlLbtbRK
+DCXVvPTurH6wxx5z7+/6DSGObP/pu9SMTy+R0YciSn6Q1GPw4DjRME3p68xTDve
SYSZliZhoBsZabDPCIhXYVwlkKOgb9qTf9K8cyQRW46GaF7us9rGTvI7ctWga6rW
VNVvrBOzSDXl53IckmYwHWwx1Fb2fZPIyd4FTNQ3NxlH4P3ZJCQ67cO8X6LMQfM4
sQSUQSEQZyT+Sh5ItEPggbRsHrfROrzww8AJZueuyqUbtqAwTmjptgmPq3jghFpY
1d8aOJ8y1IvIT1JCmhbF+LKMn+7bJvMMmn9n5p5fKyrn524pJ+CW2oc8sABo/hih
Qmq3syswo1ucrJZ6FsNGHPskMC9lSeIZoXfF5/fy2y8j2urtyMRjGEy485gPfD/g
TW6rsPANhfzYLG1HykIEOjGII7/fDs3mNvDh5tyJED7cKDlYLHz6JQSGeFtmqEg1
s7kagTNHl0M3BVBtfemrnZPRoXAfYnG5gPJk/An2jpBxF4/mm8F0+AaOmR2L/P2F
OzGuHV3EC3UXmuAwp2ltAgyBwYe4isGj33dVJc77bdRIjf++Y4gG6LcckoZ+BPr7
0U6TZUlGrZOcCeXtJwCj9DPuxD6zOciaiKrmnwAdarW3Um5+hDyK39uBKrBc+d+b
64X/ObMO9Ja4+9uvpsWxl3DtYD1dtuYYFR+cj6xAX5jv0siJSZDYH8bKi16+dg0O
DWvFJ7CwxGZYqV0ANylYyUQYYEygJM1R+71nw4G049LquMz7t8mZOgdSN7aQT+4S
JfGKenFRilDtMg1cSRatk3ophC5LLMOuGTzn8qhS7ffyFQbHwsgpQq2RXlJ/kWUj
ms4ck1YxkCCSv9OV9m3o5P1fNoF832XOF250erXRaxrQt2MDP58LsT1wsKLD4o+f
mMNyOuES+pcMS7nbURyolhd/RiTOUA2LCT07Db7ehhV0hidXWt4wqgjKH+xk5Ux8
5G1PF2bqqQBcK1VPfhTWdA==
`protect END_PROTECTED
