`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9eP9Z7ZHNcYiOBqVMKezRV6NmwiLXNYPACJS/IZlEOFM3fj6Fl5HskocwFqgTj/Z
P6lPBrni+iVFG6GSwQbmU2I7/LcZEwEOSr2YdtWUXZZUglUv3uZ2Rs0bm2gMUShW
4KUMkI6g6GXYLoBezPYOKjZWGBf3dy8my+BswJg8xkqo2IG55k6QV/YKVko22gdC
UcDuyLUELXMFDKYsC4lYl+5gfduc25pJDrGClOi4MPTh7702fJ/Phbu89YAxqmU7
014le68SdrgtFmTmFSkn8dJ7Fo++53lg4Bflu4zkfM4t59RrOp3YTfRWLZrzDBJK
CKGoKB5TvlDtPldH3eiQWRJ3erPGK2jwEnfqYnmgPYW91X1gkEMu794jVxwbHh3y
4CWxSiAx6hTG+NJSkjzFpqS2aA0uFdMXyFkcBXbAemfhJD7QLsy250lxu05yR8AC
h1iVV6FvK73YP5xFRn5J1tXJKFrH6/imHMVmLHppRQGuNNBZnu5JsKOrD2wmFRJD
o+Qz7xKqSeIWpFeojbCGz3A0sGxrqI6mVjpQj2kq9zdZWZdDz1prhw4OV88zIQMG
hvrdUIM6Msy6PMZ+78rklVQbI91+4P94pDDb21b3+TBwRv6deFYwIBRszxdgI09z
IdMdY0gprPVXQYwyWsEsmQ==
`protect END_PROTECTED
