`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dmTDdY7QYHYztMXbVUV1hpV7KDWQbYmbl6qlKr8FlAs9J6k5Sadu4cI8ddP8nXEu
OUJ35TGWR0cc2AhEExRKNUx1XdJKJYDu88BFT6DH9R1giyv7Dku7fSX85lEyiaCR
1ejyWOs31SNSyKCqRerOBc1TRsQhkRKh8DVEpOj+E0U9gxwYuZFKSWalNfTkGf01
iQ2XvJ71iOF3WK18BzNxL4sbMGxCXFYyxz6JtLrN3Gxa/kF5cW2EHmY3b/Ft1vie
HV4522muheVmYSaHavp8apFNrUVqVSyO8f2OsVi7/bxY753JcHwwee1pWzxNi4FK
yVvXH9WvrR9HnkwFScm4gfG4+ZtSVnN8iAC5Q/UajGHNlF4N8lA/gEtV9ZtJ7Ms9
dXG2Th4JCWIqd6XxMFwiuUBWjdJvf3p1hn7w9dUrNvtWdJJtqRJLzgFjpQDYJEGI
9kMeJBUMQvV4mnrryvOf3zDY7ATi8aOaMWGXHYpAQiUMC2Np2pj1uKQ7bWl5xknZ
8L4Qv9ldPeJKwmu5ORmGKIgtRGXdtbz+PpJfbcVCbbVjM/pnCSf8dyJ0HmST3tbF
+4GCCAIzigGXAF8ptea6Mg==
`protect END_PROTECTED
