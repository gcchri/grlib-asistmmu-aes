`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dXz/vld5PYKw0bB+iYH4ma5n2AK3rrtJhGk7aadVs0Sw8CGWq7eVUCN19rMoQEH5
T98wyXGvZtDv2MhyV5ZLuLwflTzixN0DEKSRSVGJ1QElA/oeXKFcPIG2kBcjFR4r
QsNIK4imS4xfxoDV4x8EkI3o7iSoxttkFZz4VAxl1HYUjIQ2onK5ljvCIwuMLEf8
y55aHabbZipf4gB5K3dfTGnHAK2R+hMmgx+TCZWKZ0+TDIq2ju5eTUjNX4/vkukr
g2PjsrdvhIyPrHrFj+Rb87zUU2uNYbScu5zTlrw8DAxxAhIOMZG5aQy+BsLqT9/Z
WbSZJd5uNfDs9qAATsxyqsqalrCR/WsKUem1zBdLGjRXlTaXn3mGgyKsuOus5FIB
CiAtTfMgva6cseYkhGdjuqWH+LW7aFDxMdFRaI/hm1CZ8wUzggyZpLhtf9WL28wu
gvzRdff5g41z1JzyaiDyJDxIFOnmpDVyieAl/euEwRCDOhWg9pAFZc+Nc8fKTV3S
pOqn4DS/YaDGOjc8VTQ5mOWe0ROEMOKOC4VDASCxdumQRVNSNeNYPn0BOf/wBP58
uKiiKotYC4rcKpCyi7CiWA==
`protect END_PROTECTED
