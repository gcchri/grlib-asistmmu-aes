`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9vB7n5d78eEwlPBVWOGsnrhst31snsT8UuoJG3kzOUCYTS+zEdj/X6/G+1LD9mLf
GSCWSRjF9rkN3pF/db5pHe1hGZUsCfr9Bmm/u3K0cPfaDrOWNYpEBLY1uBIPsAm3
sQ4XJiYx3xOOddOqjSSb48G4XdSOQ4EGDGGc+tGUnYXzPrZwOM2jWiUIpzgwZLxs
u0g6nGaR+DiePPvisaVoaxBYsP/4XgGkKfRGnBYdNv/zstwb+h7uH4V2XJwoGE+4
W2da/JED/VMHMLFNyXMcNOeZUhy8RN37FVhMcIKbvMQ+9STa+qqHEpjutXaO1pEx
tCYY/rmHBINEuVXkEiOPDWyYNojU18EQ2DV7ptoOgJWjzKUEQssSr+MHp51M4Pi6
hyS9UDLEQTOAAISvAM1rUcOq7o31JL4vD1UYqfKJZYWZkUTzl1AGj5OIiz1UyRKw
dyuYTXk6RQBR6+ATYi4jFzcC8+C4zBmS3720+5AuS1i18x7vWlT3RT2yrVdkmcuJ
DpGgrRJz7SO7CNTVeA7Y8GtReFYriqD8yaV+1hz/qWr/gzG9gEzz6MR0TvUI0gaD
lwdkWHdO9Vx4bElHooU6n21E56ehsGizlnfGPzEexZUXCyyxaR62JwyG9niBBqfI
cUoDJ7L5oMnXfsTokHgzBmwG2vhEp20mMWyQVwcsyyWMo3IWr64XixnsmvoI92VS
+GgELvajksQyxLuaxsHPEZ5NWyusyfw066wK/zOjl5e8X3Momi4guP6WFXLvsE5D
sStSfoUdVa7k+zWryCbCWXrSLxIzcX6jSLhANRljOq9v9/Rs3q7LAyyafja/uX+R
IQAHcexFwlc3dCCPR1ybhhC9aDj021TWXY60elw2JujM5M/b6szzI9VQqdxbQd2Y
IMBvv7Xp8jbjIKi1s286AFIs3NkW9jUoJCKrGKecl/oynVMriY//1UDuCKjqRRY2
J124bpdwJJC3BPjnfMk+GzcUKd/qzH5++AL1Bilzz8TccMGIkD0rk5LGLlpSjsk/
XV0JVtOKcoLwMTP4jIcNvNBtfcyZNjuxOaqfSA6jvrKG5vdsxHW/m/B/cuN6ieGX
uOyOAIz7MmWM/9c2hwJMS2lykCkOYFf86va6+lpSqfemrMj7eXoyQzZVcXlUwFWw
ZHvTKuhVGCWvohd3J6HwErtLT9zgkcLmuvo2UOtzHBR9J2gDxlq8ts+VnSPFKSw0
UocxygNyK8VgKKktKqqWr3ckBbTUKA6vow3nBibLNpuoNP1DSfPJnWX6qpMWKiFe
iaqTP/ux4Nl1rNn+Mnkh3Hw67HJyQOHLXpxepHsuLtqZ6mIAJqeE/ciGrMaTpAjN
MB007f6Zv5AnBrP+nqzCT2zBd01IbBpFWezoQY+0Nj4rKegHQOOl/BFk5LYiYD15
v1nKHQ95ifz5hpmGmDmmZTvE1PMVXaRK0H2lZZfxRGgW5Ltmnm0dST8W0OxvIsxP
20yIEp7deqwj7/sqMmIZfTv1z2lQxUIH3rrrb4SFe+Mc+6CtgbQCSZF+hGYJYY7S
MPk/V6iC6NiEdESKzCNUPojQW9AfveeMpgLGmCs41K5uNyRtYON8eOWCAYYD8ECL
4jJnJk2SGKqIjt+rEdrueURYjrWzvq/m7cYBv7JU7BYA++Kvzo1NtD3BdYxFyyXv
RALx6D37lbSfiqWWrvTaxglA0oTpUWmE7OOGue50PvssM+4a78bVDDF4WRVUut29
ZZSBYC3UMFI9sZbqhQxtxwWPhpYKZdQU0xkqPJKeTXAFNMW7q/tu48h1lR6nhVUB
bqBXEptIZw3gpx79IlMcRaNYB3mXmN0HJbyblBV6KIWorEBn9Sx+DhCWc4R/PsQ+
GlUlSvUIyI7vUJpCHKzkXyuep4960sxm9FVFjl+yULdVbDthm85VT+3kgsUxPr0p
RuBuDHlJpWYTbSdDbtSTgQagibvABx3dfa4/HOxxgOayU/+rYBdrL6MvZtu1fVB9
p7G7+ZxkF7EfgvFizDNMf/wzw0om9Rh/gSM7HRVlyVNiCyjGEStrilfZV4DDPVTm
1//9omlMSNTKz5N00XxovSemDdahSCupGt4/EAGUNPRiiwE0DDCoI0UO43J11jMK
97UfW1vCrapNVgp5KZVXRtx+/MCtJgcpznUldqira8K0JnnxmRvsOyP3SQktCLEy
WYfifkcti4uBmNVy3GG7XtLJ8j4IsJqOBcxR9KB1GRny/moCjU32xDZ2RwhR9z1u
LgHEUwg9fmMQNSL1cFnHGe3rGCvk1ZD9jWnil848Bm8S9L6pwUVgT5j+FLOTJuLy
suC7O23OKZV8x8BPlWZ1Wpcss337dXZ74w6WxR3wvqILsJg0k6jM88B/RD+AV7L9
4ze7OS2El/2i29zx/ET2/nXR0UHl197CWRk64CSDmPV+dWwrI54+niZG5feXc/aM
lXn052tcmd/NxGpwjR1HHkYf8Q5HqqnGQt1ilBU/Qc+gSKwNZ0RaC4ee5vr5tbyw
zaEmhZHoK7e4VJeWtxPCFjiR3pZ/C1sXPeMp4UijDnL/+B63Iq+Ai+vBuN8gEKUU
4Xh3JzyfYfO0AiPukUCNlT4oN+JAA8zxr3gn0Twpeik=
`protect END_PROTECTED
