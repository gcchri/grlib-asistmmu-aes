`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
brlPCVc/wGYgt7oxFGKFLVBVoKPhN7FlkwJUmtTBmzpP+Hp1tCfRzZjyHjcwJI2+
+qyAD2/FqB/fs/gDJNpRjODQunZeE8DMUnoFukEG7RXb25ubFV1LoLCfMR2QNamt
40DG2AbmJgVOjDrJJRgmqnLQXVOzRtujQyD6RVfLvhwVh6RAfxB/UobIKoJvyZC4
o+ULQ6usCpTtEwi+Hd6eah+ulkMF6yFgUZGfcpAKYXwUvARcYljTr/18L2QzW5Sm
Oj66zrj+bjIzdQPp0Z/Ix6iReF1H8yJCEj5NYamPR10aYZMoTKYfXsVB2W+beXGR
zCHKVaa+LBl5uvvtxp+piLIps92PUt8hYM33wZ1iuVDzOE0vaQ6puAcYmNtGVJwh
kechBpIUH0yE0KqQa+ZXu1cq0SacwCk5Egcouy7RbXtFTuazX5YMV+Bcv1wZ4Bm9
e+C9EIQAwHGLNJyHJv+Av5Qs+Z41qlGc61wnjQQxcVLO4OvqoGyqnVg7MH9hEOsO
nVcZ4jEsiZc2gFi5CCxhSdxPjaML1wnfgBmZ0WTonudGNnqKdb+sQTc+RHLQ0F/I
9I+62zRFE4+osPMymYhMHMaPIx7mdyGf2PA8syG3HFIJnwqjGKUtYIMn8Qp6nDsj
JqMAueVpFL3eqxlNR7tUzV4ON1WTTJY13xxZVJe3jPva+g6nGSSPQbtGgEj0vUx2
uZQXfJVUb/9Yfd7ta87hJ9suN3yqpMT0zEwKpsXMS0lR3tFsK/MZVgNQP85067oK
dzThszGUVpjOhaJWTkGXpdk7z7Catreb+GPlYH5BaaQUOAvwNwj03aSQWV7XOWZT
Ft712us/MSf+XsBo/mVKbzZ0bJRYKdJIr6kNx0KlPndinXHoDe5hw8KT2T1waUk7
9Mlp8FFRiVbvApgcyOZJa/xPTZKcR1eRtdoSjcG7BL4X4JI28oliitK5vQdR7Wy1
`protect END_PROTECTED
