`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3X4Ct1TRnBnuQ53p4XSg8AwkMlJZ2zMQG1IfZWE9BElajQYcZ/15Zde8GEGey30B
ktbr/A2hC+iELQ1380QGKZuv2PZJcBYwo1oqoKWuRQIZ26bwRLSGqlsD34ovoj7p
e01GfqdpGfCpTqnInc/1o+51xEmUflSi6G3gLq+NERg/SbZXPQbMHE5HbkiEL3ez
x6/XalogbcWw0uWNr4tSpkQo490nLrZdpcbRGR5trrjea+AV4OynNuv9DnVuFA9p
ZcJa+lLpNvkWYliV6fcvQH5y5RnAldQsMR+Qu6N7+iqDEdgRA15xN8DXzdzSAu0C
LzS1YcHiXz7rjQUlT3CN5+JB1fjfEaADOnuf+r+sfvfELgOezmKPxC3T/oNXrXgQ
FmmUfbNluY4HiIJIi0K3P2MgUhNMr+dFchU5nDDYHwKw8AwxQQ4drPoBxhVz7mFi
LvSvsUKY6SNFBX0IIpjmBmXYneGFoWxsj5XJyMo/I19Jr/dh3Zu1BaU2u/Q4cPP+
MvbgKe3mw3OsZ5+gFgSrvafwR34uTEdbMY8ZRcUumQZ8MPU6Gn5vROhHUrh57xt0
Xij77ylDAMhBVdEIOe7aHQ8mlv1BOkGl9LtYzLGh2eB7Mj3QdTmtB3iLanifQUqw
GBE7DFMwZYYhzb9z51xAmdJDQgllF/uFqJoVt1dfR1M=
`protect END_PROTECTED
