`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TaR7HWAgcFDKA1hF1SpWxwBJwTu3fSjCXDBQIKgHVLgRP0fJ70ujtKBd27S/lQjg
DEixjf9ReSMLN/ZQPnlDUEjf2xoJhgs3fi0gcsCxQcLv8MUgzmN1csGm0IcJ1ySZ
f+AaUOh67h3JyWwCAz5Hq8zvkPUuYRhM/o0sYYB/P+WGKG7PDX70YRK1Ybxppef1
bGo+0aZZ0Zvd8uUNQd334sMgV18t6Vq7Sq/llsTMaHGcWlBtHBwezqg+6IOqv8Fg
Y5iPi6mVjUr+jeLJQNJNWKNRU8qX0GcewbKPfP46kJi/6gF1jEs/Kmq/0TSPkHmM
xJ3miM6GAWYVUG9QBfMAO9oJxaSa9/6TYYlDWFJxfHMf3/qqzGI3+zwUhBS2VDPI
DoxhYxk56rn7uAyL+hVXd1bSDwC8c/ABcU/gu6zIGEkBllUmzMLQobBV1Ius0ije
agpEOUZXINjzikpGpj5KdECWRe6aGo+XXAtR73FazJ14cBu4mCVK+4wdYU/xBKf8
OSKNVcy2fwuPyvtjj/eQFf3gG2EmRuGx35w9DGwd3h6qfNtD9B0EVJUC7Rq/9Gmr
t5PU1AcaWVF4xQ87sqPlAM953lKX6wX8uKzNkctDvdd+chUCmUMGGboJLvJVULKF
fZgE3asjtFr7wyt/1iFn42RjQesofEoS4Vw6MnnqyH2XKBGH+BVJG7iyUpjBMkgH
DjQpeqm22qIr8Tk23sdAHGQCyfyMZJiitdWMNuXVzn//HavThw5duzy8BBtrRp19
4tCFNSw+VDfDPXSDzTGjpkzrOI4kUq4uwuWGlhOdSMySefGxgySp0XxJzSEOVMHi
VHqe2y/wy41gllGyjkV3wyCzHPEbY1EosCjIzTx9RCNf2yrXxAwVJ8PaaRyJmtLJ
zuTGqTLBnlECq9hCaz5RKuzq1+eXSFLJwVsnQSP7ABLeM1RhWgaDSvQ1MNQwI3wO
fLuG3w6o83op7nTSIGukEk1/DByN7GOjWINmuvfl4M8CU7Xo82lUYvpTJlPgvz7u
qSX68+vGmgAxgcHFgScqAz8vhmMw60ADGHVzCa/RSQePPeoLjwdzMNtFJBXfi3Ep
ERRZQyPpKRWDNjpdjWCH4fpVdI/p1IXQbGbK9xUpOY1OtdjLltbS2GF1CTobjIs5
+SnYskodDY50pDuR8BVa68mUNP14nJg192O56aYYdDjKhQbFJBY2eSTdNAzgJivq
GX9kaAYuO3rzr2huN3RE3P7LBRY6mvUxKxjSFVf9Ztnzbk6m3rMgnwvdBsit2HcS
qNGahNP2bBQh9la7iXCdCMylZVg12T2+7FmBMqua+AiyQz4rWSldf/M6+mituRx2
hRWnUua6cHAac83JsYhpA5g89rGxj1FjYT+iRFFWiu/o8XpNzei6vbA7tVYN1AFx
TSQnDnMc/U4Zk3MvF179WqNBetVpUh7gHyYkCaytPnQFHNsNowdHut7k0ArgHXPq
O2kJsUcILlu0wx9zs0P5n6zpz6C9qEQwk34gtbXsfbpxgxIolD8kZVvMZ/kvsu5P
7ObUqTjx5V4hBmwnzvw0DcVeRtEtwCTKtVtv7jNW42rtDBIZiBm+ZzOgU/Z4E4Az
7EKsMpq2sgB7jgDBz7wk69iIWGMluYu7SnTRHdOaK+jARHPpLRQQHYDvXe6FkbAg
ew6xuOYxR7KEZIcNNfqJJ27GFp+OyOlkjB5fFWlmXd8weEnHMOyBQave5T6UAioT
WaW0q+bLTvUo8KpUW1wkljgxIq6Ti/CU2Kf7NXYePTKoBNAna2hY6RqMYgkvd6Yw
RP/PSff09+U1+wdAn97l2g==
`protect END_PROTECTED
