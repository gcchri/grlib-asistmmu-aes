`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sQd4StNs+FkINcbkV/NNL/XDgr994V8pDgYuR1ZNvJlzBv5qOYJnpIerHyoGzPhM
fX/u7j8h2J4kAXOYdYxn1EXxhLwzQZt8Ov/yCcSy0NIqmz0+hrColah+qYn5esvu
lFqO4lWo1MNsKvAmAZpd2YA9uFasF46iIWRSUo9KapJ53bhPcxEEZZWcf0zO6Srd
i/OTm8nm9HTSDk1gRFe6aEhXrGEmiVm6/iLmnmDxdBLp5O7ciolC/PSnXcB832vn
dBjzedVrZUsj6kuQSXVkdAThXVKhLi9FAIiVjPdJU7M/LHDJtzJI6Y6aNwVoqNZv
ogaoJ2kznHe7MxH7IDG/hM7LyjuELPDLkKWsf0ie8G0u8B2ydyzoirqdHvGZvImH
F5+15G4JUJ9PWjcbCqb+KzxA3+S8n2QzYEGB6RwW3oVCyaOAcahFuIGdEl5wFqPC
iQSHsvDGxm8duIZ6HkQS5lTTriOvmyNAWXZHpC390RRIDYb1VX1mxLs5rG/snphi
fXhkQJkCeLQ2w7MKAmJZaGvIhO49YeaUkOP6EXKS/1KWniKqjO+6AJYjl+yHrTl+
bq11pqf6bWlayCyJ+PsBY63DVGcEubVQzuYQxJzWbH8b7D8aNRno5k77NyB1Hb+6
EbGd7zLWPIfuxqxbsQa2EzWXFu9BUx1cvdMuq6OEuGL027H88htJmr1hREriTcL3
5OeyG6IibNamcX2tBqPgqGF2TVFQQMUIHBUuJXkO4vXLwvNheXKhpcJtWYyiz/0X
Z/xNjw377yYfPPJfITWOZYdpzC7y83RX7AE+fvWN1Jp749BkYkZzXKBAuEDkb9sa
ROgjkEWciGBrhWqvo/J8mB1fowctMidoFW2YRBLTCNL3bBV9A59V0BS8wmPDLzuq
NkAAr7zTrd1TyW3eS9M2LKJ3FrOuuJsERIcJg/G2bu2TA68PkhsLNpYLWa1OO2Jr
DZmFN/urJPWCwxt9qNXXbj5inuQOKNYKH2PxLLeHOki839V1aMwjuQyQQPxYavlo
ChXFWhIxVROc+9c7Xj80hoI8jGIYcaK6pTtjXQbgi7eOQIaBkzH7J1Igt0/N3c+B
MG7/F5xEd/WE8uN+4RqiLtoMYRXB0R1nxLUMGPBSebNlS9PFBX4TVB3E3JEf7n1e
Q2rcRpeJGwJngcV2tLI3z9ahMFExuSZ3amZ58n9muod05CVfPW1TCb+C4+h1dvK+
inFQx/30nHmVjFDp+CUe56nS+HJ5b2MoV4LKPjhU2syO6UQ3SAg7C1nP/SWwkW91
bIydJJZeh8dIxi8TpPyYI1SA5tycX1ZabeOjX85X2mI5dKoc31SVXB1iQHi2Q5AK
zC9s9kRh7QYs7fEC+bQzaP8hzKpYtJrc2xcEzQKZwPDAE7tttEpDSE/yJZSnw6sA
HJjTKYK2+FyidgutYIN9ST5qAPSx94JbdJAsXyOo01jhVeoWP9lzVKC6BmosJszW
sJZt3O09mYfQl+KG40tUPxkoMN7TlifBdfzdXzNKSjFMqPFKTzKPQpCFuZq1kfrf
AifdzkbgnA3vtxMiuMF5lDdA/Nb5yDtGbd6a748HQ8dvxF8jsyyEkWd+gzn2G9QQ
GjyO6NGsHpcZsu+0FMwOJECiaSViJPMQ2c6rPDe1CbzaSq79sWwWMRYuL0LWsvwC
jAQCCjpEeoPCsDxLo4R82rVWeJ/lJkUSCGdsg12FQ3ErhFdHi6XAzX+hQVD8GA6Q
f5IznR8TpyySe46P+tASAHue1Ua+K9sA3LdCaa4rMHev0p1k43/BrkFwbJsopy2V
xpV05RsOU9nqiPtWIfvAEHHIeS5aO5mKEyzeUEcsN8yd/2BdVrR80K9rPwgXeFTT
Sd3ZaQXSO/R+CqWx33NWhjgVaOW2/lvBsvvsh9xT/YtoCdUkWwbQ9xgj0JZh9fd5
fFmqNFRZtzD2mTphis+HKJOKIBR9Nr58LBPXrpRWZI5QjCkP/pRv0zB/57Px1bMk
MUQ/t1pMgEhKTpI2HbR4RM6bsrGK5e82Gij0Tinfokl8fbYJIh60k9ZWS64+c9H9
qeh0YVZHKaeKe5Leyqh9nLmRaFbVN7XefBvCFIIsQeDuFtHJy9F/Ui21SKC2EkIR
8sobP3tAOlL6ClUsilztyvg8aoIpIwlX98Zm86ynjraNPWnyH4JmLM69393mBNHI
ADML/oD/5AxV0Lt7MnbJd/5t6WKxkWp3K1d3eyI7E3TVDSDnNCLnwhczxF5XCU0c
NuyB+veyw2kV1HVBp2zl+BPvPTPuw4soAslONz+DTiLfpBD0NPSj96m5pwy1C5qM
4FQVTvrDjLA/cWfUicyp1q1yx5O2f/uu30AazlgJFqCUq5i0TTsEvGMwBPsQ/j9e
AuwDt46G6OYPJrJkKV5aFcaEAVTyw25tjH/NP5PkqIKZWjw2gf8YpmMfCh8vVKbO
9oXT+gI5N4QbHMVW2sMu5hveIucnE7pb8c0mzUkYsKF0IgZc89SgkuLN3ya77Av2
gfqf2qNVOI5n411gxlWPzRyrv4CrAl1YTjdPg28eepwnF2to0Ctiao/pzUWN1I+J
c2WxcfD2/eObUOyPUmRgIB848n5ctAckmTk48FIdkLOR7mREih2qZozYQQkvkk9V
iaFS5HxPtownCVAzWcTYg856w4R9Iy15Y9mmBMfzIFZ+upV2V1HOhwVzWDSyw/cB
0tzQJUse0/9kBdcJYJzjjuHhKppBz3jiebsLtv3TQJoixEIojkIlJHuXa+Ftmknr
oklecDUmznMz836ov/g615f2qfFs06Bk3uB3DNJ/VajIYW5BsWUkKWJzi17iAs68
dJEk7pQdW/mz4TbVRJdHnwvvE1tQvhjwiA88uNenknca0B9PkESWIhiZzQYY88J9
Xkp5Lmb4EC7A4xXrBSnWfEuhVXYIpoy1WuWhR5g1gktcA4zuFEuc7Wp2cihgjjMU
2b+oJQt9rG0aQvbGigYUGaDpFwhRtu1tmWtnFdm3QZMOhUwz3haemG499se804xA
lezSuS5zfntqwKua7ju6FJN8i1mpPpfbq3kH8FNGWzox6xTsi/70X3m541SrUTf8
eWlASmPgy2jUOBJGcT87F9xgV6GaV85J0I7a/eZS6Qt/c8xjJzyuR+ZLENfLIfP3
aVl/Pq8Zq+1prg1ZlJ4LvJ+La8mIR6xu15OMZuMa11J/NcOsSTQNthCXrCHbZaSs
1w6wehL6DCSbr17+FphCv+MLD47pcwBw6SXCmb3T4w46MtWJMAhxYAeed8lx8OgB
Ex/Y1Yn/fNNanjGWoapwBfwCiephSlXY9V26ZBezOKMDBz0iIl0VchHfSHWFFTdz
OlF5Ha4Z63dF8Q1PEsA0YgB6S4jSRiNHFiPfCUOUJLmE2gGB4MhNASMswiJ6ADx5
CiyGBBlXvO822S5ioOWF7xitTWHLolSQOx+7FAZ0JfVXFqUcPjJN5SBSjvkQJ6VS
vCyN2kfFOuIxCKFVMGz7gtu6TkTt69s15UObPX8sT2dCnQtkcQmGVmn/Twq6AatQ
nX0BvAIlioZRZjzQ/daKlJmwZZ7ysxlK3GQJaNP57mIx7ymTunnLcZr7WHlHZSl/
ZjfQ/aSQHPWvc7gbTLOllzoeVt3Cb1zRmVj+OuD4jSZrzKwBey3YPgKYt8M1V01J
LxdJ1VZnsV6xewyYDrxP8vjUQYzZgUcFjfe/CMHmLyPIbR8UMYhj4Eq46dJz/Z4F
X5e9z5hzESAS4vxeKQ/CQ8yYR4cUSJ8xBokIO8aSE3Sye/Ur+q64UHusT/ZAdKmF
koqLCMZ/UmE+SPMwHemA4hxqYHYH9MP/+XVxc+KxQGiUaArkpZ64AfQlrLTS3fmt
hVrhMHa6re6CjhoiGzs4ESDVMEOZbMLV3KQFTnbL1kYUN3V1cJHdt53PAqgGOOh+
ndrat3c4hDftbU1eyJslhVLHJTKLQzKbIjry/Ua3COj7Rcpqexim4EDa36hpzAXl
z0BpD3Qd58egpOanyjBD1TEB6198IHtAboLz/VYTq1ZXyoUjauFPL00j9VUAcpN+
Oxz5LK0DB83ayUmMFnNrGXalsS1SOfKz812ZLbapDfhrZ/bS2v/GoClRyuoo3fLe
M91r7tFFi24vyy2uYDyIKTbTyKU5WrUo+j30VxzmZo4tXNDiAc6MVjCqex6vO7CQ
uvcrUIWEk9rLyQ0v5Ddffcqo0ST5NYraSXAzypcJ1wxeZ8VShaOGEZC3rIoUSxFU
w28O/EkJdJLxF6cF4VOCRH6rjPyqr01Ko3tJx8vDmR2yBXS9z90KA4Xy7UX3SS5f
tf88k8eOiHt/iax4mEsVEfxwye2xO40m9DxzhaSJy5+ttJITe5JVVri1CpzuObO+
3LR9DlpBmkVSbk20QUMhWycXH189lcmg8r0mZ7IiVlUvLemKDpLuDbgRjW+d/hUf
+sKrgmZ9DsDnh8FcVQxkFRWwa27WNbvygt7UgF/I8lUlO7LMsojLHrW2l9Vkmqxx
PMmccZkIcgr4qQWWbwSocDdERLR6gOoEFupGoz8nnD8iOdFnNQLXHJH1Rq6TVzxo
h7zNW1pz1//H3wTXBn1u+9mFL8SBJWK+08pb4WfhqMoUw3b0v8S+iwf+vnKDq0m/
2SD11oH14pP8WXdKT+aXpCzzI2k7vWzcQZuPdP9fEv+OZNe7mmg8dYZOX7t3ZORc
zbLPxBIVopTJZC2UTyKWICZaW9ntoKJSt6mcPbPI9v9Ug2TTH/lydg1ASyYqd9xi
E2xBi4XI9NJ6oUq/yabAovAy100Yh9jFbCX9YBmd2vaHEqwy8wtLLuvLsjKy3Y7F
yrCQDFaIGH73E8PDCQU0UkGHtYOaeWhTVKZn+FaSLUDzBO9bM+qd8V+oaIH6sNyl
2HPTk/8JMfGFohBLbohUa2tFPPBqPdHv3m7FwVKbvEgPSeIyhGf2EQ+laGoIxWzC
AXxQhv6OIbwvq+VsfYU/AjTM5KuvA8+1v9Hy8z2opkdZod20y68GfnTLkzo/eVEG
bvoDGtbyeuJh/wd3KQDkgEFP77o/obgI3552uimEWDH6R799zBdUzXiwMq9apqO5
gXvOuK1vvSUlBOJYBOqdFgfLWJjx9qHQt+s/R1jCTdZgbxj/HO9g8Pf5wVd0fZkJ
IxtMTRXxm8Uw5rmCpukK0eNQ7l+cbadOgFhgHQMn9SrHJeXl7pZ7BWRUttT/+KoS
cAMfvN90WFzD7eMtMcjNdkwYN1n1/EqaXInd7pP62CrI4gzOnzVIrkgZ/y/Zm/ys
dOTIdDEmgSVwhn7OOXh+DeTqU0hrTNTMPJlzHvIKigbUZcJgz/UVJwdgyK2XE414
CtbvUr0L0eko6HNbU7/qFjRvzoCV3h0gkhVo9OXN4UjLSYR793r5cl1gac377dCZ
jLj+xG+sp89IfJgH16bcyXXDgNeWZDvPc0T0TLO192ikismBzvweD4sDqZFQZSmO
hBlWwMyhTdNv04yyokpr8f70hQvb42El4u1KcnQRREdfxQIZEes20ik1SQCAxYhj
zRrC/c7UCsV/WYMA+m1fwLxRWYFnQ/4QyrRxm+0oQvvZDTA+VwqXBgd+5oGcOmH5
iu0bKpG18PG9zRtk/6xqT7QFTgGd7dZstYXZbrHyIzikh63UYG1Kk3mCN02tgkrq
J+hjgmnqUE/yVbSsLsWQ8Qs2wG91ZwY0wpWjjiZL9236TstWYkG1OBs1po/LUd6A
iNtJIyoogErlQd+SC5Y0JgIAer7YhWAukpP7zsLrgcHWKElLYpWsKINjm35wSHbq
BobQaMtz7d30UkvMjRvyiTfljRjNG3WC/r/pG3Z5mcuMH7yytvpO2w24XMmK+1a+
kxBGydGpmeNMjIMRZgSeXcGSOHnuxXp9U0jyGDL39CP1nsxjEOiRDXR5lIfRz12U
YV8XEqcYUoASnGxNi1La33z2r/A0k/Jn3jD6XefumKNqyJgPTjZajFxPcDnrd1D4
4zVe5YgoV8x2cOo632Qc0jzjt1OlW9PCGXPMfHBFhVqR6MpCSx+KdtSOIMRlJsFQ
bV7GCcrJajj9TVn7B2MBHqw5YXp873P4TvkIfAqEi7XkDrYgndXD6AT9+wDLcVct
6d5u2vmYcW2oCGlJNG/cxK418ZbY56ilFV1bWz40f0NHt+ODo4Ifa3n9xtwsVue/
/WhFzoNgO525XEK6KPzqk7ksf2H+3KKTcZnq6IIgwtrS96KuKkZaXQt/4hX9o7jM
oZ/h8SdM1Q87q/h+WIj2xCQHKzs8lFD5J238Tkfaafd6p+MezZww0wOuVxup6EnV
5OnI7Px+gjSwIfTrc6k7mmhTacHJRD3mvslQZ18RyFRaGXmLIPK9twkMryycPgwL
LPdWZagdlkxR32RjIatJTwOcSCk9jsQQfmfs+lwSiB/m8TvGBOS6khjjTjX5s5uM
PdODuqjAQYAM0JRvV2BlsHHZYl5SHWB41/I5iIWl+auSj1zlzD2A2CGNr37S59Hi
2eSPkgZ/8zJQMws/z4fUF2rSfH+9rbTEbT9ylJW9NlgIrvhh7jiAs8KaREqNgfLY
IMlOnPymUu1J2iFgVJzMnv+dgMUnLvKw/R6Tcb/8AMkE8XQyHTsYypymKrnJWl5E
nB8S1p4K3ow8gCOp1+wnO5d74XwfxEa3xPIcb1ngbPoFW1crNaY2aKVGxD/UlRZW
vhlj0P/0Wn8HOfLSMdkVhoDZB3UFgy3Fx7G4+msY4Phl3bGtYIm+g+tDcvqicOvt
N+DvJBGVBKBDu70SQSm2pR+CmFQhWql8yZIDlvlGf23NEVFvwnGZClMNT2PAHoTG
YP9Dfdk1cpzGqPdT1pnRj+0EoVJ22iKYhxq8UGWOBNaOyrcuSyb497K7xJwcOk3Q
jjbDeILqLVKewZVn0IoQmHWKIzvWiU4koKgqiFkC5T0WcAyTF38BisYIF6RDiKjf
hwXBgSNPl0pxnCIwx5sqrPXsuEHjl6s5kGVhO9gKMosNfOcYCXVMdBUNhqqrO2b7
ldBOt5GLLZvwkhQW24pFQtpTzy693UVSZ28q+S/WvDg2d8KuNz75hiRv12kSAluZ
s99wc5Wx71tijc9n0SmRCoMTXdhCqpuZ6Tm2y3i78udpfkOKW6lVVvEngPe0IDcl
Ft5KrSzo4sCNOTzAgmrosbe87RxDlxI854mH77/j/Kx6o2p+nGn1Phqq1qdy9NGM
a9iG7+d0sxPH6t4TjPdXMJ5EiZTHTG1hl8eMyUsjmDy2jgTrsfSO9FO1KiJh5qnT
wF+fbdpQ4gZbu4Ejf+3/mGZdFslpilvE/sWEid/pxK3Ugb0dnXN4q5GwdXXxML0A
k5O/b/UxBEFXOQE4z4BcdD+TAHrVmQN9OMyDzqoiIiG7UkoeNRAiBsGa7e3UEcJK
dmSGWBgIUbBra0CVjCUfEk/oH1icZXTz2Z4LDlqOYsHW6b/NMK1BRghRqohGYPRu
Yj9QJacjmOk5goXK1/TcEdKGOvgYhWmvX8iRi8XfHTLCG9VCv1o5bQeSwa736XuF
ESnyl97xXZXPyGhlbUCV41hmeif/cL3HuQJrPMjQXpliAxmBGhquIm4Atw/oRfV6
8wY8eIogeWyC/I1XxM4plhTmOh4M6dx0jaP3H/GqZl9St7R21C0OyQ3s6zbq8LNo
LsdUSOkGFP/aGYgXj4B0nr2Tg28yTO6Bf+PEGuqqii78GGJfd51alc1isAZ4zBO1
jASiWwKGTtQlugZ8Z5efkuR83ow97Nk2nT7DeMKe4KqptfEeJr7ckLX4v9ZHsSQv
fhHy+9yoLp8b3mfYBsEpLvqrK3kt1el2I6AqY/N+ql1ZTmgcGnWtQPkRW9SMjOFo
5SuGtQmiZ5ty8FTk+a+0HLeoKM+bplA/TR2J5IwA5Amn7c5eOdKj7ZxN4cIPkeTJ
IZ5cW0KNH5vtTd2wDRYriaQxfPW4VfBCEGBnrB8QoTVlLfyJv//qwVH2z0iQPGkO
rLyZ6Zo44l6X++ARcO0JEDgbGDS8JirRb5y5f5rqrg3Qih64czDAvzPReM8+PB2P
0gmmZqsrLJII7WG+kD59SMCQ5Bj656wH/SzeCNcIrtJAp4W0/ck8W+euTO6mDZ5Y
Z4e81CBTs5tt7pbFjMORa9IqYQlqPjHPmEzlLrR0BM/nUB7msaN8UbhGbJQyPaG/
r6IKV1iLN24mEWalWZCEbmC3FmfE8dysbAE51rhz4/Iw/m3nNEutKOef03N+P30e
KuZZ2D+Y12z8/QtrG4kcrMDPJhNsgpNZTJlU7PrR8Y/gL4cnk6g0+Yv3uevxR5ex
TdCLNStKhKevqDf0BjqAgBdgSK313z74U6XOuc08SVx3p0RYEXjILJghY2Pm4eWX
589nuNPIU1xhqWdyYm77GQgUP4AWjqYoCcSz58ZlPSp3TXAArn0gwYxmbHL8rcpy
dWC1VjRvmeBitHCcJNT6LC4o7bJeTh4nROGBoqOeLrkr5dGw4utLDkwtKSu81rKm
+ivDJvf/jPu56qO1ygNWj7fyjoRkaoUHCTpOOPSsQo7gKTtIQzVV8ya2pE3MVZQq
+uasObqlZoCvuytzbXCHGoClEAc/52BGIUlPz7uBc53OaBg0gF2yHTuA/EjZMTrv
krxCsAMw5W4uUSrxWVNIaSfbNKDFxPUtB/3ahRGYRF2KlVNxyzmg/y6XY3pPtGVk
+gC/gSAiKQK+uf5CdrMDZG+dzysoQawjZ4zVioWM9JVM0OB6nJegAWkIIDdo4+HW
qGm1cmZ554i2FkzxaDmeS3ztzN1irEoRZW5AulIz6pKKGpJpsKn8WCX30eWVuYaB
LRtuB4CAQ6jRDcxX850yLetu9NJQUtuVZ4HPOKcsMHeiHO2uGGwxHgoYqOuKhjFp
MXDWQaHrvARezF4maOC6aUMj7XdiRPVuS8fW5o0nfE8d33J6pt4wG+fxety61R6v
UeT8mw8M50FacgPLkebGVI/6h+UPG94J/ALrmVc/xAKZJoNFybWT0FuZlvl6qSwY
MdR5w6y32ROW7v6/kg8bm4JxrkVyAZOqgNE1mAAYhid638QAA4k0I9YPr5eOFyZK
DFWdh6W2jZDLfLQ581VPk2OW9gg3WGXEDuViSEpgv6f2GFWLoEUvW9Dj/h9AJcsf
wrppZVHrOjBk4X5eGqnDfQBJGAMPj65qBL20XSLQx1iHIeWIGkoxgqiRwc3f0XEp
2Ps2/G9NpeiYInDmCoqINwFouuzYaNZLWwOR/P2ez4gK10zb6Vlw4e71G3jHRHwo
wBl3ZkeCzteS0/YHx61OB1YjKT2kWNnHaoos0ys9BWIDeQqasRJVuwmVBxEQuFAW
9xRyFRBnWTD2ejMTEuRYyRFEgkdKo8O1i4EzySlpCPoiZE+DjWyIdKiipRi1jA4a
TYsnT9jEcZHafDOpEBQau8MFYDQ12lmr1N+pPqOFgQDPhl490wOc+KjIEwaf4EGG
SubHKgMY8frIu9TCKGpZoKW0FarxHhpcy0ENM1OigC8YTsFjyBUU8KxkEQmm7bNM
rSsu3+Ji6qg9JavkkU9HPs+bT9v3P0whcxkEGjDcj9Vrli57ie51Quv/Jk23V6j4
9rmLByUix1q6d33uKknnObHBa2caxbmh/z4usz0cIAoDCvbbfyQ3Oe475nROwAb3
Ej+YiJFEPsY+LF9rxlDv6gUQb88Kh6C4zjyo31VncRNiDskvitr5TZH0FQ3E5WBp
Unr46r3VXUJxjHjFR8uJqECv0ASzVrn0ZwddX+u0rHPduLCTsFo76JHx2ppMguda
163CHQ/JxpxmCkXcS794N8D5BDE7aRJfDbGxMkImyUJqcbZh7nU4lm8d2N0J5zHq
sGFGONJ5jViewRwjRgdoSr4Ig8jCpS97vNGuF9PS6hUpwgdP6AMfdWwA921ZuyYF
RjBHSOtatztHK4eiuny/3lv8hgNTAhKQys6lchO2gCff3/DNClubRYEAqxJoUUkX
yYyivj6smyt+vW8zI2EDcKl6A+Dx60L7tOQTP1wLOHTwnBVcP3UQmhctRncpATyX
qvrXi4teqcIheBvzREbGP+b/QuX79ncwWf6KjYN6R0uOP7cFBBgUZhkipoHJonTT
7w7Jgj+z8uuSVYYzYSzVpnP3AyQ5QLckqy2ftdGkVrN3QqT8GlmrdN+uQ0LXaTOt
I88xf3sQDtLozC6soSm+WuylodSJdoQ22EmW7g3/IRXNJ1NoOAd9qwFxOh+fDgya
UDu4KL8zIuAN9bkseXpE05k7BP5Z/R4XojLNQDBKpH3D+rG5YfJWDfyg1d6oDY6O
YGGgBwfxbeXx0UladKgLOPL14adtoggMZGiU2sT1Kv5FeIp2eXQnaL64F3bSAneN
pgEQFpaQtElmKt9sHCgwWfB79CFEg6HQzs1hPVmckiqxPlKJBASM5E4fe2oNmsf0
Gjft2xSyTYieLOlhDgbiKM2GfawkeJUNaSOuXs1NwdvpM3Qm+aPJLusACv20tTFt
MOIIQ52xoEVAo0m7N8BbmOFFl58unyvC9XNXKfl+gx9jSiyIbPGt2XMmG4IPrQcl
KdSBOAl2zDyWzuj+b1ykRyHhZIVhsTQpAr+Vf12n1D/giKrhRy6BT3hDev9rdTOL
o3F4EiPa6RK4D+pLxjVrMlGj6R35Ze1jsWfFswxhYQfB6iXB4qsJrh0sFwVTainq
u2P1zkSxTqJ2Sa+CA6QSO3r8nFnZNhrt4AGIvb9O7pEce6YH3LWPFw0REmb0GWf6
AnxhzI4PQL7UCeKsdkuD3Qd3pDBCUvTwUtysd+ZIGuzYUZjpEwPTgPD74q1xdnQo
0q39MergSn8O5QWrq2mn5qgTY5CHY5SjLEONA8xKIYtSC+52UpHlr7zhIsPDeHZO
jgvefN/7z+VX4+hDr2yBIkX8PfTSs4SMInoTm4ureggArh5orrxepI7wmr9rcrgr
mUM00pDQsHa52LIpOj33lB5hxITU0b0Izal/vR88VnTUrbm5dQS/3Ni0FfI5TVlu
u5V4YWNcOOZ+FsO9c8TIu7GuVznZ0G6gU8loR7Kf3hz+sA7FYPBuVKKfCbsFbrPF
jZNqfOHSOVuaeCdis1dMboRvO7BwyyqJpS8OeIlrj3nXXz5af1fVEnJMH7yrOfaE
bxrFcQxyYl1JfhkWP9X4+czxigkm51nYfUywxMiDDjZ4VjFKVD6nBp5ncMRbs9Wn
yWF6Oc4w/g1YQ3IGfjtOVcZTMNM578ZvnFtC7GnHK7bPJCqimBHcHQGQakG30Rn/
TdtpVTmi/Ibcb84/tbJlW4nH1Ob6qRPq3DaUoDgluyq5XUbtT+HCdHN7bFxpLe+Z
UfFGAJobl/FCK5JrdSK6VeBFzZ8VP7AKdY9wMXgUdsVPoCeoAiUKBWXEuzUbFbDZ
b16HHLJAz/Th0hWyJoNjkF+C5hY7J9Wh3a0AoRC5OY5x9fCaJr2U62T/F+Vp61Re
YNkk0xHzJZDf7n/0bPre63Xp+WbMW/tBYInPg9auH26ueZPBjzkbDHeq65ZzqiCR
C9OWDalvZjydYnZm50ZCEvXJLwdug8A4RBULVp9MieONaEJVZNMou/CXaskfWM4u
1FcXkIraQYrnnbAgfGzEmkeQ9PmGiq9NPrIt/a6dKQB8NIJ3SSxegx5+6SKNtBKc
qcdcIe/X1qNPIVTXeYjhXJ2BiJgenpub0MQ5JhALaqaO+gmWY8Yvzp7Bh/QbQmBC
pOJMtDB1cr7Yh2/ahNfXtxYQAabZvMMB1OQRzbWdmZXFpMc/Y1Aa1dcetRUjIgR7
wNDTWU+l6xh9w6mNpxDsNNATGIhq83ePVcFY8bDpIuwwpKtL6GxtTpFWiKHRKr53
AYJFh1Co1pPubBl/WIZR3VwEJKRl8j5bN/4+Qtm4K7XIkof/H+vFfIZP9Ueqv7yT
btaRBYaWToDn2RrT70Xh018fs+LYkH10B5G8lQ0gxXA8srWlCWIKQsyZxT497VIn
N4TGx9s9Ls5w6u6ZOWthJS9JmPvlvPsmYeQpyO6a++5MrFWkb6plqtS1xzRtcrhE
cEWNRK3M0GZ+F03pwyZtlOb8V30/SSFPC5NmwBVxUnYRavtJ9mRjlFE1ZHXnesCX
2FiXquQok82wEEmV8zn3FqZob5vWH9Ym4PlbOJXZH7+YKgHb6gn1Ir31174TPO8T
3i6Ft2JGO86aMPzyezO+hvy4noQQdwbfJF5sNZKNYLKBdMHnwv2Rxj443/zSmwJk
2mn2YRvaU4Lr5BVca7k552Mr0FL0Ubw93yegDHOswXQFSjRlbq3Ohp2G7qTCPeic
TC5a0TSjwxFIBPFAh3hTEc7KBOkR6jYPeLTq4Vv1pF/+/K2NHoOy+umkMsbqqex4
l8em06F67ThoUZT5ZDDXdEMg6Tn9V4hbtoEx7d+ACP35UY4GX7kRS8jBgtRh2zWb
UOt+yUzQQxpawKVAufjCK3nFEpg03rEvrUXoyWGL0wlQ84Q6nJIPaQR/TqZt6a7a
wqlOahgsxPzQS2ZFxrUWKZ23jPW8E1WPg6t3wffZXKZXLrm5T5xiJ0FE1AEes72A
ECNhmg0hatP3Jt1tg7yA81xOFKFO03DMu4okp2jNYU7/FjXulUJDIi/V7lyvdo9S
gULu2ZQziWU5oDU7gg9tUsY7DMpCRmFM0fGPbTOoSEOBudgezSj8hmUGGjUsvTcu
CE5X6RT2jW4LhuQFUPXNi85Bl9d513MuqIeIAGSravVyLR41WYImzZ8H+3ljpX3/
ABIjhYfs+vabBkbTkOmasfKQ3qDgzJ3aPoWbw13sKO895l5b/XC2K8kYHzgM8gEr
vBExG3fLSuNc0EY3R3MBjUpaHw/90ZFT+ojvFitg1I+ZjFgV4EqFw45Er8KemZ94
ovjkUPnFx6NimeuPb8UBP//SvwjB9idjxwfKidA9i36gIXFqvzjLc7Y4sSRGyrBm
jBdDZFJ1KnNTcRCe7ztydjRnRbwwI7evkuszRQoHMijEHcWu/hvTZj2TwW4LNci8
4uiksFUq9f7W8GbgG0tYQImqHDAwoCgGUtuCDJm7BG9Qo4iokLJvjtoigiDbzel7
1Ca6bYlqPDDUKLB22t0ALZTABIqsBidTbwnySk2V8hduNt/iccwRgaToJVKhWrlt
4ReLZTMQIC8y2beNO72Yvb+6V0MOROMmPfVT9fHbtI6D8bO/J+GM7+Gs/4h5iel2
ipJna+xJKFzBei9S3BAy66C18SVYl8OqTDKSdHveaUT75iDkwEPP6pw0BdF6vREU
RpUYqj0BF8m8XDiuZz7ZcRCWUZAvcrGBIEh/NsgBxQCBbpuxdiIMD4PH5IBk8yYj
QaG7VvAvIGPi9PBbfZK9efR7gdxFCojs6b6d1gwwEAYNlPorgAWDwD0KV4T/myNO
VvMWQDBLYP/1lXblUzJ+OdP1QYHwneY3QA/fBqeS0U6IcVpUComCfdTlWAJZraD4
O9l1fQ8EtZqjmK68Z498CZudzgv1x/pAyzCsJ6pC6c/TXOlBNFjs3hiadQEbpOuA
cKCFfjdETL3GE6H3o/tjJq9G71vekc/P5ZcxmOnjbKrmaxoPp84vvmM6EdBIX4WJ
Km8sJpi/QWncr8NVyHrdutWs96j+sJB2L6y//l4M5cm5w6cnjJ50cGC3tQ1rrlAB
tOxLvVS4X6nY5liXiZjWe4nXwt4ymNixg+MwudP3yDEw3IMewmtL+o5+ipXwTJdo
ohpU+ArwjWxErKtVY8MALq9QlbtqG7TG5QrF/3EIvYRTnwUwxztjDn2QcERTvvfl
0OhTr5hOxI+vfoqcDCDMu3SbmvLWqNoNsR2FhyY6DqLL6onmkNMCVbaJM9V+/xTE
rII7GyGcdsatC6ZlGjnlug+KdGWkruSXwpubJFTDaY4CiI9Bla+GGPHvIMEHB+4x
At6PoXuDTYIcUZ+/419BgkD62m2bWUqMEipPGA9ZSs6bAoP88wTCugQizIytQcUz
2IfSb/Dpv4lpLC0awkdIbcrfr2kd1i7dljQmOCQl4N7NFjWNCK8595zc8MBRR9Iy
TVfMuOP5MJCcZ1jr6Fq0clnCLPNZHkArpr2K2kbIXT99AxavUjcuK+eLjPauCv4K
eKpdoNTApSnIA+4JpY3YChbgE3A4tdjD2lFbAilNajO0mwf4AsQwxmtrEREyuJN6
dhPgvXjYN9fUH85nD5y7PplcNBgd+2YB4V2qJN5b+spi1k1GC2sXhW6smCb+rhw5
VRGIbN5//A4BWIU+mg3sz8mYY00pcrzGtGQU2H4W6KU70XeHjwn7uGa0ZaROnb/9
h1fjjqfSp7u2/p/3hhERrRJLSlE/SqB/3xQwcvQSwzB7ZeLa/AhL+iDGwu+88WAO
szvMVwQi1g5M2QCm5SaaTBTnEOgTya4id5Wk+EUukqafdhKgfvkTKejiy7P/tQnt
JPMQx710rE8A6QFflGv76ZWwfiRxwcBTKzkITZ1E4QyQOd035hcOvgwp9dcDNk/A
5sq84YCq2xg8uqHkAo/VDrrow9MfxAqUOxBOvswQVAiVCyTmHmqKijxVGQQSaHK2
1SegzA+t+yMXD+lcpcB1B9/5wPqeOXi4FqSp0pXTbTevmYHRHDdcElaWVXlpyejD
Waz20khzAaIHIvfDd3SHpvekJKrtj//br0shN5lnAgzEvSCUTQA+VGzb/l7t4ntG
cSK8gbrboO7La4McGPMAObdm1AFgJx3a6ypUxDrK9Ua4ZMEOnEqpAM6NJkBU3jho
eyYEnlPrFjuaYzSuX+ygLfXVdXpLOP+ufmkk621oGUdOLcucQJu2Fnm6KOpR+wfh
EUUGuhMxSFW3O8ZZBfWq6YednOmedvoEYWIBHBPcgEoz2k0R33COWBiWiXXvXqVG
gx81s6hgc/mGWHQkpgBQfmvdSWVNyHXuh5xZiPqgNRuqk1/B4U11L7jSbFmdmZdv
JEXSDV0OyFVqugc1ukDvnKc8kB0zr0n0ZU9ekGTsGwOE/BscM2tQ8DjT2OiuhE8x
+4QpW/rIozifYv+ejNiVArfSq7tO/YV2jV5EpuUT7i2YcJcBM9DVSPcX03+7JNTT
20kIT6TPK/h6syhMj4NucDj4IEeltKnOuZoNB/myn7yGa/TRUd4FkaD5QTcbGN06
lIqjAMt4IZ4LI/mv1mXdpIDiokPBz1fT3d0UWiSVt8Fxu8CiwKrhpPukIx5K0w6P
9fO5Mgi+9Mj1G9PPgy4NZ4vlOm+6CXXCNeW06/U2aNUpzezub4XjRPgVMCKlfSXZ
u7ygN1mMFerfsaFXV4/6aY61NlxOiL0j4+WXl4Q0mV0lQjEveNp6+h6WpKVC47T1
ZpAL9YQhZA5Gl4ZlOkAKIJRJlGMM/p5bUGg4PFRV+YARemnMI4LA9NEw7i7d5Pgv
dYYJ2YM8uw0Nhgj5OAh3UjoOFUzF3jHA4uuaWYpjFY64gPYL2QKgIl8JuKi5aBlU
+ow4oh4MaDHzssuAJiRZnjct+PuE8//9Ypsxil4WESr+OqY/L8tN5GgvK1naa+Uo
+pgKvceF+7aNHyIwtfJU0HYnQsLXgvW7msDkDPblhXKQtvHpQxNJCKhFGvcIQlzR
no5xcc3VLbjHQRJBvgGhQlaBt/629JIZn34ieESX0//YETiLXuOuesdY/EdLKCOB
2yKQinTsH31uWnesMgHsSP/IsXr/FFY93jW5oXcV6DuANHRa/etLZ2cpwTV7wbJA
Hlhw4Jt779F+KWXBczfGrDLr7GijHV3vdb5yYIaOOWmpS9OCNtvx7oZCYQ/ENS2B
B1XxZm0FR7a+aIKb7FZQYu8fFHQqAQfZ/2iLGG7kMZ9cWfvfeT2cvthFxgBghqZZ
Cvc3KSPv6F1R5aDwkuQ7Un5n4s8TjEh86sTmQIR4wdJlvPEY0PCkgyO3n6dkf9YX
kAYffjJ26uoukCc6iqtk6WA260EaKsj4l1LYvRQXHwjx27X5XxCeDOxynNpWYuHO
JuowCM+Z4vsZW0FsgsMDzfZorrLfniL058RfxmxLYZ+XrA0LcY12lcLghH1K8cQ1
Bs7uBYJDfz44RoVQzTqroGIv/1H/ir84NKxiUCz8HLGP1uvu0Y1cnGKFLG3u/9XO
zoZVp4hdPwQLarM0PVgRH5S0fqzHg4vrCukhO+z4wBQfktPxnxMYB34boX7YLoqd
TcSLmzuDdfXNh1S6TPfNHzk8rMUrMLOPOG5UnCnHEO6wFtbBnIEsYGroVoEFf6nv
mZzR3RkbRL7RBuOD9vh8+ZGGUp29mFX2PDCBXHWhTIqStsmq+q0++C32HShRYG2n
Y0sZXz8jLsaZjKH/KwIdMLbkpAZ7iKFTCPSd3+0FPy+pMUjvpSwdGSS3n3vVIYMC
rZNEV+sNpxAz8GxFwgoUBWms1x11D9oq9p2jDF19Y7IkYUQMvskoEcSdKjk0fxLO
Lf0WPjwC88n/w+MNG5ySkfZjy46LCZqbaTaPnbSJWJ4llaJ+mqZbbLFVdir1DnYi
Yl1WNJkS4xPh9VTcyAwQRSe95uHB0QO7tBDyymYwl4Zo3j9zk8pFRg4C/fsyWlLN
TvACp4agq03bBGA7ZUjpb03rZeogebad6JYYhD2x5V999sD273rpuLDg5lxpkTmP
QqA2Ecr7Fn4IVP0fWP+zqzB4sVAojsw4CIKPNYXOOvG/pRstr9vt7IqLQvdhvz8B
cE/jlpT1z3Tl1oEGmec1kLptn/EJUfv1rnKP4MHPajurk4SIERblOvWWFZg7wDGq
AdPdYeDfft/RSAbwXr6mZ/mIVm18n0FJiBV25hYB0V7azBwHcA6jzab6JFOP2cuM
O55kE9gpOcRVsNdzqMB5s5l/0Gs9x6TJLzHTgMtisYfKn6rz59S63e0dupMH6a2I
aKQUKHbdpAMxg7ZD9Xdz0KrE9BRcqBVhNuhriKlRn+AchsIRleAUlV8Rft3Qsw4l
po4/W1cJmkTL8yVZEhMlFPf64NSfgAFe/sT4Ymp77xx0N6+GFdTOFDv9QdCrsAUA
cZ7y+ywpUEJt6p28DdVWB/gfhdIM9sM24Yz2dS2Tg+o28aYuFMrsAG6hkoUcWZvA
AF/mdpStpB3YOZlFugoAQfgL9gGCce44Cy+PQ8Y9GmdqrYzxDcc8Wo6IRn9rcXQi
IopINaknPKt1y5AhjSsjeiEV1I2ClUzweObzwQNZwlA3NuM1JzzVHYz7XazpOyt7
JrS0akniqQ70mWEMc4omManT0yGbEmiXWGkP4yCLxBAtrIWRoU0TgMRrBlM4PQLY
kNl1s+u+M4X4VVXjXHxyWOh1gBfwvl0yDyIjBlR7Z870n2ZxyxtJpN8YMtFrtJNf
nbnIGjW41tcc19RpclpO0ADSzEp7CAVBbarmpVmzpVokyvUVHjLkCo4jdcklHNR2
eExyNG+uSApJjomlAx0RABa07qU1P8K6ez8bhOClARk2lXmJGLHGXOf0/3Kp7rOv
Cq33W9FKt+dyhTUo25ju8HuMMro3b9eGAALyLhyzOImlB8Hdmz89xW89vnOsshpf
FjGtBBq3CF9+4Qr0qjZz/nKTOOPOT22Tjlbq5nBNcxMFB12wxUZoHOPWf3idkVip
hcuxB1KKJouBsk0JE3enObanhN2TUV2xlGlAoN6jafoGMnzVATOqwGSpgJE9Z/tf
iSKXL2VyR/jeTjgJ96QwEtLqYK1GKRm93sQmB6SUUKNd+ZdxxF55602+lYFDRikS
y0+c8RITSkUd/4NG4VMCucPFTD2vODQPzQY5WxO/My0OKHIj+v99otqIS4tRwN17
BhQw/d/3ep2C4Cj+PzDqjn/Kowyk+TgAc6okUXZD130+r6ZzX2EoMwu4Y5wmYbV+
rydYrZJ5uoYudINLHxPUwKgUd50OupqlMPBE6rZjtyk/C5efaRelXXSNoIdttE8G
WG8XxnnWbVzv8LGHJXfZGX3qBW3JxeDSJJVU3UlJLihrlmcI3MzKXz0MjbEBbL0G
/JGzeAg8o5xu5KbU5oYbqPAt/AdxOZFeYv104DUO9e8EuS/gFLqppotDVxkZD8RB
9QfS8Til7vTLmIN6yvq9QxXy5QOc6NHuqN9BAZrzbBrHk89eDYirPPRQ0tgMDb5h
f0vjKVQ2GMjN8YsHLafaO9IL3PlwAU1+ohKV8SXNIXXzhc2VEdkG/nVUIReRCCN/
3YturcyzSzR0QTwj+zOfdpMqqrL1aixs1DMrxcNheUa+2X6BXfgLESJlm2OY6PtP
dE/JRYWU0D1JmMSjxJSJqBWVbOhfaCKzXLHyZvyrl267VCvCMfUFU5WjnElmn+21
Pagbb0AGG8Bs7iAXsETMfaIT0IkZOlN1SPVGXMqVlkj/fjHqxuekNqhc/J8RRfPP
M6e4hFqlNppghVT3K7wWe4WXvUj13d6gqH3INuzpUUblJi8+OHnqfRVAOINafbBE
yAHTN3kCrBNMNWH7kk5m8t80uTfcBkTpPY8GQHGw7ePQUya4edg9hWtcQW6IkVt+
OHwjA9N4wSaYMJBNzkeNhddx+m06xr6JbneyJfUK9HV4QFIJ36LF97uHVSadO66c
QCZDuQiqPDwSIv63tdnzESV/ofYlZxbZblG5W+Fm7NQ0+IMByB6byHyiLx3G6/ps
fAs4+r9cWZ8bJrPeDqptnl1WBex2KMBDQgPzXUWSUIxvGUirPEIeybOxqblKH1PL
nGYGGMGvsifCUHAsOyH6iRiVpjKC9cTGpfsXo6XSy/oLmLFid/ZCncp/oAM8WmEi
XXUA4j4ykhxGJM8duIcKZuP71xyo9hXLW0R2y8ab47p5v4pFMPdSntYK52yuTrwG
8s7CEqIAKcPXZewsZW8l2Gznlroxf3vvKGghhRowl30e6cQNlzJknLa6rM27/vaL
bm9cMRU+0Wn619MNLsVkDIdNLlTUxHNjFOV86/X/m5hr4i6KFJYObYR94xEScJNP
Yc0ihRTWFbEPgGp2v0JKAJwdH+hh7j7QrySJApL+2NNdiAyaGuga/aftXXAEuPIr
3BW5/rKMf10Af5uW+QUHXQmEiSpoxSOM3cXZYRbP9egHJcJtdqx36cZ140v0/WZD
mtt4BHwYFRpZoRBYA2BmvKwZ26WVk43qHYfmvURFiCgPbNo3tSKmor8TWPO+5+0A
XOQJVS6L/8IGmtdMsDIFXrzGGEbnXcPQFnB7thIMVkoA0DgWecCSKc51vQTWSDEz
yLjEC27xIFX/Bz/+6EmLduHdLyicEMXrLmOMTIS7Fpd9eL9x5vjz87Kyt3p2ko6T
JIZeIlUdGs1HtODkWHTTUOcNVY1mWMF5pclXlUwPosVo1/qCb+jQ/s2lCynwelEr
DHaJ8FLeGdaGtDbdKwi4iqTGhwp663+L+sQLcOaVUry5ROCXWjA4rTWK1YtiTFdD
1cd8MhoRZVUP9UqjB/UUGEag1Ril+gxTjcPjaLkm4AZTm52X/BlmPE6VGhICF5Up
NotU9QMa0+MeRMM+uoRxXDyTIrO1vvN3+siRDJygDMNJVLsHyu0hMPoqVwWoZ44T
Zrf9e3zGCXCfG/8pJ2dL0tL6Mz1+YI0Ej3ktrf3qWlJhyFG4bn7YrBYj0Cw3dbjd
DCsN6vKtF2+rr2eQkUaf1IAhpyvCmU3igxB9zOH1+qFrY+GUQN2r3uKSmpaOuRJg
MQj/A30L9Fr0LuO/a0NLXVk0L/cxEZoSO53It3gKW+BqOw/E4CYiZJy/twy2nLD5
uOfgufHtFR9sf3DpBfp2fQVHFrVRF76Ei5HqxfqbT3jmQYHgc2MfXryoW5Fdsf/c
+DeHj51FjRrLOgystVLXVJD8tTZvcYYjP7HifSkaE0XX0504rS+mFuvZtL2KTpNv
+He2KuGjWjNlpZxmuz9XQslZrOGGbcSCCx0PAhuWpcbD5satx61m6kkaD+t90YpX
RMfkPqpwrDi1R34RXHGbxyw8XMZVvpTcUq7V/u+1637s9M5KnwLSCHmyn341ch1O
xWR6OLuQ3reOxp8vBRqek5PXgmPJh/tB+OyeB1uMrxKjWb2mDXMtIgJ1h8pCc39Z
pl5eEBcWge2vQ0Og+VHcI7FCFVrXSCPz3WCJ1dFK/35ukddsNkGQgCt4+uNNIQFx
pZRtcWWVrDFDrJDf2Pz4Wu6v+2xFTYj7OfJGnfmrC8VCZH8AYIGsyU7XwAToVKCY
8gaAM3vv8xH033UsvwP0peFxVwEwFe62+JEPB7cJUcZ4cZDk9pBkjxI5vqM8gzYA
nTfTUKmXMs0dzgeruZAESGkO1Q9LhvPxOKI3A6VM53tpvrfVe5qy6r0K+EVIuWxE
xLVp1LhW1HmZzx9Nfz2VxNmB7dZt8Jpgrelu7wl8G5/41YyiyB3rXXU2H7NJ1DIv
qwjTJ9F5yCZDPsoJ4d7mFLVyaCHpcEG4NTu+Y15YfyXgRg6rd8sCu5vSvSa48tJT
FpDJ94SDqfbeXwsPKz0o7YUAFeuauOmiUIJLENDOksVX7vY7hK6U8mbRPhiC5Y3u
5qcaPe5sXFdNJE8xioETMIzR+RKI22FyW3AxwOtkr4JEiPSirOvUl3NjoFsIQlqn
z40V8q9NmsEF60MumlxMLfnJJRy1qrqBFNYmzpsbCBdNOnTibfyWr46qEzRptdwG
G5ICNTPJ8eQe8t22pU9IznGOoYjSDkWZXxf73wW+CSFpGTq6B1bGvDs/mCWd4xws
ShAK/TlxjIDlXgbwwBwScjwWLl9HJ5+7o1rQ8v+u8x8XLTrDJzF8OYq6QQs6MvAW
AQTKCNNcl+3tlPdGTzJipXpkcC2Ya5MwyJXLkZzgw1dVMKhCk71MWwVaDoQp12yH
OoEtgnoYC60xjYXqWd7QXHix9aGKEdNwIkurFX9MorPY07eJsjZEGu07pmtM50PV
y/pj9XmPhv1DXCzq9dolwLAdTq2QjQfb0zE4qQnoegPDolR/2Af3JKPvnI5MunLu
Hk29tXLWGepEebPixmO8jOWwoagZqNWUEWpJQtyedRK/mUG2hJryIfE6TSRu+1in
zNcsCJX9dVHp/APPI4tRvewCU5XxsgInWZPj2OtQ6mBbpFkOrQpcwPI8d/PNNaXJ
ylO9NJWiCA2tqI/TAIaRpMGVyw3H9tK3hVZsHGt//PxxcTNN8Pa8LXV99be9I8Ty
zfiFiBiDzpRm09T86syoaW+JAq5EVLwWZ9wsaBD1Jt1HuoE5fv/kClQmTmrwPJpz
Or5yTgZBLMXnJmEcSBcsq1uA+2y/y/gIlfFjgmj9kFaXGw4D/D3vNurPPr9dZmnR
ZEzIZZPy+00elaQSc9qa3dj22VACzCD343W2ThfXXaOlOf9WDkW6kwKpl+wwYyuu
0QVzJWUPWzoXQX9W0RLKychJdweQZd770RXmj2qPO/VaBy9DM9SXpy89S9oZi38b
HvMJlm/sMWJOMBb2o6QMf2hJZ6Vme8e3pza+1irr3nDXK0fRRh2y3XfMQ/VpQBF/
v8LZDloi0d4KDO2qyClnl4a/Bhe/5Jk7tH/PWG9hD7t8H5+tLx3XNK2xOjok9dj4
2wzHZATiujlE1eaLq4hXSDdCWd6OsHOQb2mXdAZ2wUA+12XY1KUGE+I9K0AA4AIE
yvOy6kPxf/kEy/3wiIWUjfz5EnZVRIClEly1U1HPxGlSOBHUPrnJdUTfzbnEhZa8
gJ6kaAnAEHtmMeftkV/pQ+5QYAMJutuyc27nMynnlF2+K/GBXaUxF21+CBORKDJu
Rmexn09ltmyEGl54K+FZsG1eXrUkU89MfbE+4SfM9mGAClrGXrHH6bc3a5SO2bT+
dbcDiFowa3hfIsfT+Ej4lMEDlYoXtQp6bB0Kxixqa8dRlgPMKD1tq9N86yh3kbgg
RutFsoOt+3C1/vsZUFcAPPoMN7rlVQ2EmhXpWVQL8eWFdbPAceQCQzTLJh4f3Ybv
jrmQ7JTjrUecR6RDQNFIb1MsH5xnWt0+i1pDPS0JNGLuKCg5N58nAgr+pog+34JS
soA7PpbvJcb1ui7T7/58+ggAVhCWDvQ9Wk3ZXBfAKXwgwl7+qehrc8q8wvv3uujH
X1PCG2keYtiBCbdxWkL8nqWVX8dP9pG+kYwZuoDPvNaUWgCgaYs8JU67kU0opexe
npUMEneVYZgEGQE/exiodL+4PEdN3cJjm9fDGehKKdl04h0AmkHC+rYmi/1SimVZ
qtbvcAzBBZC45796TH1GFCRJQ/6cLXpkmpjH4zyZer7xQACjoKd5eirTb5pdEqfc
Fv0p7NJMXTx5UgumVsOAwmrs6DtNS5VBuhKqIsawHVaDocAKR/sVwAqkC2K09H+M
HST9tY5X1Sz66bvPp9ucFkQ8sEfO3OBkt/quoF8JbFfGvjhLjjEr9fb6ePDhyrZK
EMjhqfTUIKB0GBSjm28XS67bMJcWYAdaf32n5O/P4blCnyr0OIkZ5qrYUBFA7sWS
yqalBdCO6ff+jlELBTG1jzdNMxYZT1H7ujcKDdboGL4RPCbtJHb17B1iLoWgR0wn
itoJW3k8oJxEY3DTrD3cMywLhnuW+yVHHQEhrErKgNXu3xnnGCKvQXhJfPfoCcc5
FkdLWtDJA9HxzY6OKAoc0HQLhd91ilDKJxizCiddTJEJ3FhQf+TjG6UxEU5TXY0G
rND111F36BRu/uaOALjka03rwyaucTgWv43DH37UUiKobqujVyXxipUACmRn0hEb
x7zAyZTa5iPxBXk32avaKYnM/ynus3ptQIBvBIyAlVkAbqpUwC9C5vcoF2RyST6v
QrPL+arxS3Ygl7mqlYc9g3ZZEChwRpJASOs6E8NzsRjvQiko8C+LrabWuZkA64HX
bFh1koIoexg9AOaSU2bSrl5QnzyQqNXpmAkkrhu7bmhrEEe34AYn+yuHsHr3KXuH
CpgqeFPB1Cs7HWiQexL3Z5v4VcIkCIAfiBB5XMTovH6u+c7gDfhMpnQn+BStpshr
8R/LfCmOWYf4W2X/muwYTXw7/vXc0qV1SKRLU3a2JfpVmvZ+I55x0War4/5gBERu
aZ6NFRLVUqCI+QPxkOgeqqtaYx2W09Uf5oPPumWFgo5AdB5lNWjzLUxQKGV227a4
0uKrXhc5EJ1kg9gPw7oORzJ64w/rk6T/K3rO+3l+W5F0QAkv80gt4Lv/FrvQVjy3
ItSibvlAiKg/aBNk4LZw8+K5fh9HY1ksRz4eTBJKBF9uh9cbBaSWoOfyi1SLJy+X
CqooqlTftS3Z+Ur5/tAAz0JKRZafmoYLbPqUxNdOCqWLUe4lZcK36y5dnsOu1+XO
5hLoJmvNC6E9xrmcRT0qMq1bTtyePbGhKqIgcWi4W4/yX17DFfZT6Xi6gE8ZlzZB
Nm+6/PrN6aZY90ohtJNsiyK3oc4GdPbCzoWuqJ2Mphg36yaAFDu2wO8UvQoUrXQK
zzsXhHggGO/3peDd8HmPeyqe4h9fzMkZ2R0VODXrDJ0gSj3PSkQ3KL+FR5mIexpP
FeNU2uINKjcJ2lMjzwO7ZWXMJzrxGSUSLQQsntj3bP4g/GVDwpJeQS/QF6ZykD7f
bCpO8mNLC39Gn0THBwE1pkQoGmX77WQV7T6UiQGSULUuBgWzColKJptJzYOAEj+a
pcLeF3f0aPqRh+vuMh2bJXzekKQSnDqlqDJZbk8NujvDxIDP0EeP7Tvbu1epkA4L
vf6bHioc1QyJCWi7UinVgkDDvrMV3CJWwQyXl96EdE4QbH9LiPk3QKk1IvSgr8g5
7KY3NSJ5VOGQMznrFJECHvoY0a/NTo9wF63Zu3GNQze6HvHaHs89TIOrW1msK/yU
NsCyBgP7IPcOrNKCiQuce5qlxMBYA/L9GT2ZzBcaHmnh62goReASDO/XU5t2xKJL
OMJEwBXPW8lZI0kMBSZ+N+MiioIxmWrVgCVLgscnvkzsthiaPpbP/eA/BNtW4M0h
PRr6KLVRg5YqeIu+ikDZBdWAV5YRWrOmo4ZTymqfhgYWpTDElOC8zftymVoUYkJy
9YLCm7gQro8K4hrMCWtN6z2wFfUzE3hdyfsOV1KQw8ivQwo6KcW0wr4SdOALM/jD
Nn51Jhtjqz+j+TlnD+J6NZggTVEWYiFhW7/rrlbpbIe/HI7dpCKqsM54290zNIga
4lWCRIkNZW+a6GjVlUpJtZd4c/2Mz9f0nATHUGd+Nh6lexLai1L/R2gV+vLINU0x
CKC7ZVNvhiEuchaRIj95qkDGzdcIUF+JH3idXqUybfppUTyjb563NFcv55ycfJu+
BYPvPPMxe31SkYJM1N11Ub5Fu/8c8fPD4HE3vli0WuJ8l6DOg5/3li17CKT3IDhw
hjF+k3ZmABAtnhM1boh6KSSsnukDFW3ip+vHF0sXbjm5hOsEDUZeoEERjGdWmVxF
HE3MLsLrb8WfMcdJ69Nuuebv4C53qpHVz5xWvQmvG2kDJooK+2Xg1ds38WFcSAaE
4LrJcv+sgiEEf1a5MJsl13Y7OZYeTheI3K8mPb0Mx7lAFbd0TgqM8tqulXqgaX0+
EXoPbB07sLdpC5QXsupFNYnDZuBW6GN9f4qCU5FFSRfT9cyfyXSn6xsk4cZWbu92
ZHewv1/ijRjzAoV1WlSEYR0LJfTSWY1xwn9EKBzXqETTHqPRZN54XwCz/p/T8SKT
Jv5IuzYadm18qyGmSN6bkrhJsyfaC/RkNefx5tvbEvuPSmUZKC95IkVmYTgRKUdo
RPLzy2jlxCMmZ9DxaEcK1UGFcsfSztrRMhANMmhIEP5mU8EbYblnFpKLbU2xvoD2
5K0Qj1HeeGmPXvxudLNhoQx2W+qhJVpgNLw0+x7iuzqAbDKSTaxRm94DwTDckoSU
ejWtiHJHR99HxPNrfahK2gwT3DDY2lRQcSVx7yGmH6c8dkHdAgxXdAX2PYpZH+sf
J69sbM0rghCjJCujNu8A2NbpZy//uJLYMi2K9xaByQXJEvGshvF3p5/fr8+Xrf0D
bJxsN7cqKEuv8zE0gmf9lrFDfQRdoGdX5f7j6WfP1f2qBSMqB/Q95g+g29864gPK
0o2BRn5YFZvdhwf1s1SKg0wry/77BEU5DfQjyfHTwPDj62mqyvGX35auVsW+4i//
JhUOp43iXp/C5aalwVK71bBHAPIEYKd77wSP+Btm1V3RC3i7btfdleZiZuEdR40v
2uKh99IRk70PcZFBhdujCNZJ+S2FzF8pgN/T1ix8enJLlMHK0S+tvtWyuNyh67GM
PKU69gx1WXIoFuLQag4yBAapSmOossVynMTQOsOBNOVAYmwekIaAYQKexy5URNc1
9uy0VsfSbA6ImH0CB2F+dkIIV64iQluYwYceYZer+Capv7LjOEpCM/BqHKl+BxiB
PCVNmgvqYjfkZ/ZIjcVueFg/ro48g5OIVPSYmkrmStJ6lg7UlraEhqHmAiOuWA9C
d6wlcXQbD1OCFiKN84ry9U/KTADbnbAmztIc0rlnk5xnON55ua8MYdGDBi+ZtpAt
VKYtBlOPQna9Qbn4HdNOIx62bkRwFX3xtq9L357ZvxpEJ9ud/blHdijOeh/9I/1n
GoX18F9CiTyVxQ55n4vLU7GH5BGuyRKUpYMrii0xG8wBhRUu8WsXYfkJzaNQJsXD
pG3uZN7O5fZ91xN1LQbo/gsT5zCCGhDs/S6dogSutvhGQc/joAI3QPX07fi5aZu1
eWXN2H+CeeVK/IZJxLUGaRGEvhhWm05S2N1PwbbVW4etvIOcLPZrtzEq0/f8hKJc
VFBwcpe9aY5ABqL64x9yPJD6OliEBXi8NUZoi3ZX9/ueDJRRbljTMPVV3CPhvuT+
XNKNdxXuFv9/CRJ30Y3P1WKwtq9k/PDew6AnoSxA1k+oLsRGRQHLrx9eLAi1U9ST
PCM/Na4Atkf7n7kjFo3BmvkZiHyxX2j+aBsbKxZKBQs3mD3XU7OHrMF7bMuljVnX
9hjA2OS9/AydnfoX01QJpB08cx+SsjKEEjzMX3OPy8BquUBC0F/DJ4EZ4D9lEO2p
lgFv2S9Mp0WVXiVuLjbG3hu1NdtPeHwpCds5A74gIyAqWZdEkJIBipV6g0KD8Kkk
x0CtprspdR+6J9ycUtjwQMJHDo85rhIIb449P92+nUUj2VXH/F1TTVjJe+7ebpZ0
xjRc2VZnEBQElu34YtGLTnZAwuzVUc+lZP8zyOmEbUoB1KUFNzUNZDq+S70iIUgl
7moedBO+QOepMGOTGsQWtKkNREjjUrim7D9od9SnhIQw76Xl+Z3InzgZOL8Oc5cm
8Xs1AgAwyMkvz9aZNjSxl9wFoGomXVBSi+7F6q1SmjDW+SgxrhVtfy6BZbxAPTfw
W7SpsxSKSgxZtecwkBJBEyWzu/A6RCmTwKeHa9tCVfTgDqh54LKI/T5Tv4oX52DO
zBwTHPfozvhwzAVg9Ntj+DkL7vk5t7Qjk6klcjIxGomYEmXmPAIfsOetc1fQ2MyF
u+b5h/IiXNp4ZvU+zzVOkvTXYoPa4fWLbRTYcmE+jdYd0EQyAwbHX5HkiyVM+wTH
XrBuvcaFpI14GlsnQQyuUx+rx4DjXKTYfmvhN/8Asodhp7C5jNVKeqOBt/Shs+r8
1QEVwAg5aIARgpjnfriw5nMxiMXrGxmkMA1oVVU8QZ7ne6j+zMyTFIWX1J/aOL8Q
S7tyIrCxMJTl9EMZVpLkyGq6OC29YX0Q8iIo14s6M1IPnhyGnh/BkaHY4HZh/npQ
c6se+zHdd6jg5PHQEggVKn0JsPQbQvT+Elxk/EPW86dgoEXtlLtxXW2ovCI1GByR
m4k2OE16LbVgisfg8DGhnDkP5RGivXfnGuLsiP5uTeZPgQvs4YF+4CMEtJPW8FNw
tY0SlL3/JaonW2LEHCZKcegFbvSpZC998QbArjHi5tY9SA9s22GKGrazUxyCk6TS
4z3nlVHdR0a9Ilw2hkGyNXPdlUHnLs9EgCq+XG8u8kJ03O1mpu1LlmEocFStWs29
8UfSjrqnFuTnG7V2ViMofgD74ghsKQbaUbV6SD8I6dZFr+e73s6HgWs6tktB9Owb
DS7rYNN/Dmv+twmyJfkAuwWkk4hQRRjqXtYHjA+mQv1UAwV++iPHIv4vm7Ic2Fh7
QAEHAMW373tyZRvjGhQKZfGpOrAVodQ3BY/Xg+1LJ+Oga+Gi+XaW95h2tkYWuse6
FhSAm/Pz1vOkI6YyzP/aR4UlrKGnVscJeKTFDAB00XG16z+Mb3QwU6T4Msdm2bm1
m8g/6GWbZuxbCuaqvqQZpieqFaL3s+cY5VtgSP1AUrTXdFfWiDCC3PyXH9PTvwyb
zRaQoYLcAkENigvJ4+3ts7YudC7DRWYIfxblP+SoByynZoFS3QpqFNfTe67ZW/Tk
4J5pUOlqrxv/WFw22E9O2tNN+6H3cOAg+xfVjZGHi/s5HjgbZwUqHvNmsLSsNxLj
wxbv3e6ZzIvQxKI8mWCi4ZT73srwUIvlWZATWeBC2BdYiw6A67QxD7yTc+iDLsC2
PM3bK44EhVRHr9Ust9sjFrGFJhAzq8xPG5AfnZVs/MFWwBQ3yH85xelLFR9bUPYI
Gdr3ihp3J7piswlQXJqAc4QeRMO3H8CKTl6bkxSMo736bOUGQGXwngn0pZSzu1zg
KiQ64Ot7qDve76uwyHPjZJxA4jxzEyRH39lEQgFSqwB6SbARylzTbYI1odkrJbkA
SRKWjs+5FqPuMICkokTx9dDh+q0pEo+CJMdwkz4zNhTsNV6ZKmUo+Vy6Mr4jtATs
O3X1GE/MYPyVH7WgPiO1EmpXkAYNpFHNX3DKT8YFsUXDHRiDpFgS3YlctKHs1A9b
rAjBIuBuypwW7CGMYiBWER6c/u6c8geMFnP7Yd/E6s1TF+8qUu9H5YvejCYUsvuD
e8vMpqGbNrdugDSWgvliXfHzVNxJO6OVE97/xVjEjTq2vstDF3ebFsf14jRy9uOJ
dmeIWLmPTedOGoOqohDzvMuz/LYWzNc8a5OO7wrhcdU09/XGEyKz0GBAZDuP6J9U
zC0A7sHDVKj82qxrtZL0koD7NfRAszCt7v2582D7tpMCXwIYqrc0eebvl2TeF7Hs
PP/5dg2JkGFKuFbTrPo7Te57GSVm6u6mQ9TnVU/+i3EX+ff8EuVEPxxbVRpiNUkO
PHYcrstFnNzrp6maS3mKvyBmtayTcJovdIThc0w1TXi2y1uJol3bSKKXbtRG4LY5
alEdU110BjHksVl7Vj+1KkDr+jx92BhzTpNQak4/pW1FbZDqz7Mvpc2l2HcaWE+N
Sp47MTMXCwGMwfbC9w+OwrawMxk0ZzsUCztCH6Cp7VhpFc1Y3D+ANJJex+kXACi5
tHv8lO21SfI/BcC+9Ug4I/Od0H9NEoWF6idh5bGJ+wEvcLgt1d+D5xSKoR09QYJq
h8GfkZpR9SVgAV4wSIzPLpd2hFBnPaTwi/TLpbMzwRMQnS3FSCQNKdgQLEY8A7lu
6gY6G8ugNheUZ/ZG4fdk7CacrdcAgZkL5tBQvvOpcs115EuXFiYrBUJ3/Av75xcT
gTtKDCnCB7MLlB1Ocjpjs9qb1hbGFyRpupuKzdwe8j0uqQdwDBHSf04B3/FkPf4S
Mii3JVMJMiDXpcju/bjh1bWHDEyjV/y9tAl3wn7I0sz6QJFW4GGE/pEKve25pcRv
3DrJNGZrWmvjmRTgHkjpbuKPAP0ZAJKJ3NUrSKLH/fdSk7Ad5UIEJK/K0lqLk7g7
o/BldiFvrNCQei6GO0PzM64mrWlCfE4fsFi4ZlXchcWOjlsMouM7OSLYdOHwtOtP
+ojH7G5JiAgiZ5rew5ajM3sj5Xxu4sQkK9M+a1D47aoni9Oha0+OVjcRoPv0mgTC
U5VhGm8EtQUOgDjw9jvwaIHEgLbNtKzvHBR4tPQnYA9hGJt8Eqo6/knu6cWJyRSp
CDp9knxpcSkVmX0HoREGQQSI/MBZ9vRrestqJx7Fq+f0Wq9XYIRBGX6T9rpC0NQz
9vJVtVk40030m36hbMvP+YWDwpaMGwyA9SN5rjR0EX2iohDrY607vf2qa+qauB9f
URPBxtpFae746CrKO6oEj18saskqVIubFdPs40p2VfpWpG1KgPkp6xhKboxypXIe
IBX72c0T9wtHAkxnw8boktCzqewxr/ALl2NLB1r/Vv3ei9BgzE3vtc2Ipq8QQQ+x
437ORmwwYOxKWC0Nb6F01uAZS+3DC4Bf5kO1/kf+pxnveWFD/ekkCM0hqQUqHIFY
JBiUtMjomcfeEtyG9DLH81ekOYAxBIzH2k5WZQZtv+YwzxlVJGMA6X/owVab5/8F
WyuSNoDEapvDo53FpY1JBGxsICqF7Dda7RVz0d9ehHasimvt2XN0eRY3/neMvjVm
JNuDE4j2i7W2gQB10iYrNNQhgTzkJ6NhNSseO4wceucuVO/dz6n7+59dV3Ed6fDg
T79kXgmmoTfiSxt4bCqAMuYR6B5JWZGaEACB2Yc1V+4Xwk9PrQVqa2O/fLVwC/Nu
jwMbGG2/8r21ja0ouD+IFK8AmsujB5sasiliV3VsgigXOdPqQua/oSho3gAQmdDq
+gZBqwxbyuigICXPZgetEhZTeU8m8LXfGuEwZbPrEqeyPCdr0aF+P5rZr1tbygO8
L/OYHmo9sZ5aX+IwFqC4wN4UsFxTb8hH/0h4i2AwKRhK3zrAgMtzH1flXTSKJh8E
phuusxbJqf1b/DKVtHhjU79RJ/wyO+JguFoGJtMbgXzY2Nzs+85+uu+H8EI3+w/X
KyRcbchktpwy4euN0s4lyaMCD63xJ9EDDWQdzr0Z1QT0mUI8gMImdsHkoot2unwT
mhA+wDkx5vQRwDR+EA1GZZOCMBLyJp2C0Soe4+8TzMTF+Dm2BAyBZfxtGEWJ4rEf
MQ2MpwyN4Qa9XECN86ejgzbHjeFxlQPOD1rHGxbzEv/Ca8nuFwz6LF2CQMp9n0LD
/nvhlJhjZ2j4KpjP2kZAdeoanM/9h0oAczg1NCqdXwz1AaanGCqW/5JMlN2S05rH
MR7gytEWJ+gUnzs7418Ck8BDT5NlHK6WqxPR4v0uijIQdHHVBVfeE5iARuODHfb0
qQKMsfDXFkHCrYj81lNKTMAjY5+J9BOW1hYxnaMC5is0Ds4CnDgmTHvU/fNz2/6U
Q4HDJKIEy18Nd2J9L0XlL9I/v410ImRG53SIfVq8LMTR6XKDSc1tOqLWGdgC898R
d1TLdp/4RRQYBhQsuTEupEIyV3JFjzgtld4CigjrRyrCqtr8XZHckehQNlZS4PQS
66Jekwb8Ph4hnLtlueroR2ipP/qCd5vn/fAiD1Gn7dc8YsxMh8a+yxK3TpSiPUsV
OTMmlfvSglNPEgzMh6hd61Wugwk+RBK/GrRpy/0gxQa0QvTOxSaupUV4YtjXp96+
+H3t1qVaSYliiAl37EG6vFWS7t89+ORz5CH4uuEXcdhulnu4Ng7NdF2mKcNbtx0b
EinK2FqLzkqp4XlJgaldZE5E7bJI89RBa+1eUglWdHSpd28TXiMkXrlULIa6676A
DZucxJLKTQcqEtKmh5DK0BLA9FFzCrbjoeliqr96xTWn/IVkCf5iS5jbmf4nikyH
OndRGmCb4y+TTfGPsfD2uuH68w8K8UZBikmPrJSsj9i+73r+OivOEQ1/hA9m6UVO
qQIPfjRjlaNo89FU2oEit2JjehGY1OZrRANimZWjWgceTeop1baMZ1AxpUu8umZp
4ucmPKDhUE2YzrOAWhYfU27CbCaW3/G/py2KLQK8U5Ai43pW1xzvOXC5z5qvPoxI
v2pXBY/yJIjX1gRYN7ghy+/hbdLMWqFJNHux8Nd2h71tL/KE0DeeDT1QGfjxeYQx
Nz+e/qqLJhM63N0qTSEwcOMEJUIuORh1lMw1rZp53stmOuSmDWfiMXxEjKZ/qpYv
TwV/h41+Scl91u64hHYwzTKz2ZxV+x9fMgz6yyGKwnhV9nApsh8hdANUSufZkl2+
W+TA8DDPVrNULaH1s/2+kW4iGV4Pgwib1Z7jmb1cAox2x/py+tYjgUwJ6jjWX5Yt
DvZklqGwBcV25AFKMP2o7Ca1YKjQxQNn9lNDOY56j3pE3aqirw2oHik81YNXj4Rp
RnpFiftq+ePmILQQbbgcnEVty81Kc8B+8qA21s/Fu7iFFurJWsNQ9ThIcx7Pk5LX
haNQxSUAViz0aTphrtCQofMgAt2NFbTl+qJRd+cq75Hk2kyfK7wYoOhzThZnCAq/
StRR0V2PnPka2c/2OgP+9rzTsrwjWEocQP58i1sTB/VCd1KuaQyWc75pKZW0XXO2
zfsNXC4VeFBVlGpfvXsUQPkcB8l43+fJS2gPcylN2ORhywBBw3EGzCvfxQWRODiH
JKWsj6QVTLYCRoBkWpcY0P6MGBtm5B2ZKrsD4Yv1u8/TEwW7izxuC7Z7hj+i8UQd
MseNZIKd52p68+s43KqDGKMZIwrbnkN1FetezXdVaWZkZ5Q+W1KUjqQiwtoXlBES
7coQ66EQiEyCuWq4MLbmhYMbYszNsXNXp/X8MhyopoO6jp/cvVMbX+o7Yqm0gKaC
9oXqwyHfUi6pJgoInSuE8+0afMeZyiiMliDkmkSmu1MfNhHi3RdJSzaDDG38LMCW
v25295LwDCrCNuB2Gb2/9IVeQ7PnFsx3xJjRcnXlSCwWsZ4QofoBoZIJF0RoOjV+
5wX6lB0DLZd7aWZNgBYcBKdl8BD8lpdakKzcj2rBKabK/4Yo4YZ9NBqUSQVFTyWT
LIG6yqyaidC3m18cfwPks9SiNLIgeJbYHOXbU3rg9FJU8NfWf+9CsbdVPrUz/nCh
BG1nJaBLfRzCtpzQ+cFP/ATZzVbxngzcCe8ee0Jmoej8mUAHZN6f++09o/VuewZ2
zaB0Yn3qLEZ7337EWtDQn0uZHnhbzHryEXMUtwuALqUE0mEm1dG3FWn4fVH8GhjI
m6WPkWeUe+dmgSxgPE3nnnLXkH7l8KxZ2Au2pJYZtB3akk9WXd2EWjUIaVNqSYQB
101SV8wG+sNcH/uw9S1zvXJeE/yqvz2vUR5++S11PZlLRyhDGZj54OY1gssvtLrI
2RF98WCGUv+DqbQgw5qWyr+XtCywT8D2kR5i7iUiRpLS0AcayLPG1GmvOPPRuwQZ
WntsutYsK/1WCIZ861JN7kr1KvIdZ+4/UGdCD+vY5V86z4B9LN0OS3wTp8CKKfyw
UK9ahEgQuTO4hPAI+GgFU0jX4MF1PLxztDAj6JJ0yzawIHLRHY8dWm56PUyvbfLP
1OTmVMTKqSWrgWawTrKciZldDnDiV86/enn4ayJTX1XcNxJRbocrpm/CPfgab2TK
w17QfgKczo2JkEKNMggdEriPR3PoSzdKjnF6qgE36iEYI47mAqVLl7dorbmrnlck
q95mQePSPUVJeA3uSiMTCv7pI8baNY3wXSAHquZxX/rUrEqfWX/KrJpJ9fEuQ8Ux
NuSynF9FR9CfTXmaL7fVgid/+a/ZcIg/fE8klvaFPDnJfpmoGSPf8jvKR5BINcJw
q7OLxhN/AeaWVZtP3y4gH+bPYxU4qEb9PaU8TCnmcVA4voTTL5rOD5WVi1J99q9Y
BZX5JVFYcjZuPMafUFRbt+L8J7rTMAR85iqCfXmn5B6ZiZPXHMYxDtgSHoBkgk2n
CbHONUecCMWrjhRYr6lf7TQgvsO6XvuUonhivz7a84EJBbTpxz4d8bPQ0xjPno6l
T+Gfkrjr2SKfJ6LUCNeh6FS86zjyrh/9jA/aA6cGCKOZe7ypZhHWgoIAC9LIN4JX
Y/0K4ugH/p5BxhgpCg0R5ws6oTSrF3UnfzD2ahz937azHOgaOlitnEHLc4dl5tMZ
P8pXqWXlYE+6S931qw2gW2hraCE73TrDAOT6KkOfqwTJdTjD9umNhH/dBF7r4zMr
RCQotEtra55+VeNQu+bNUsZ/Jm2GT+jctoz6iScVmvVshrsRngCUyC3GDOlNFH6X
P2a2Te0ArZqEsUYek7l1QRpzfX2nymmvIwe3I5ibH9EDPksXv2Bvy9vRuNaE+UL3
LW/eadgtYuzPAQlTDoOqLWWuGzoVG2BG7kfcGN2gsdmX2BcuvwdsJcAu4hrlGK4b
rWy2RQbjljBo0nlVlHWrlqaxblNMdQMfRypO1QKK5MwEEMF3LBiyVifBMby+apEj
a77ZKwEWtG5It28H5EWGkpX678euHAxJqKELImac4F7CoLwD3qeYBsQejMnPRD0c
LTHQoBupRUAfJQZ8+E3j64tOm6imCTD/+arvKbqIQAr50YU11LlD4tMi8R3QpuVn
yH4qCQVSn2KFgw8pNAkqdoFqEcEDIgyznQLrl8vWR9pSLtjLmd4bm+gbCwJVTzxU
eTYfsFA92q2lOJoEdxmjT/X4DohL9VmR0XlTTS+7TEip5G7Nj9pk9TkaioQm5YFA
jxHRXvnnt38s+RlddFYIBQS58wVdIhtaRFHKFxsofRuq+UySbdXYmjFlTFCTPMWm
ygqCC69Wr27x//SsppThQq1lRdlZgae07rO6pyll732JkvlNHAU6IoQsVC8E7WhE
pboh4C6uRgB8VQg3n5G1zLQMBYK4kU7bRXNEv6q0Vz70Em82C9cO8xEzA09RAT5q
ABIZYdHJd+4QkxW0O9hEXQg8yNS4W7hfPs3CrvRsbf5InuReoK7Z40ZRyVFGKD7s
WnxygrByNLEa80mE94gs53PXuGxdH+waOkQg3PpOEwFNsLeWtIue1Uk1gY034s8t
1F7WCOMT1Idnff2DINaXlQKPqo8UpFHJ+UOVQZV6tvFuzwsJzE6+UH7QXZeDkoRQ
zWVzS1XhndK0wth5VKzJGBL+UrBtpJXqtI2ZIjCbDdFhAAD1yso864HCrkoMna2o
aqK+iwHvy1PbWibM9S+TrxyurJPLPYsPPs+7Ra7BfuI5+19q7cdH12oFKn10Jydi
YxsLbX01bHhsmWDxDygItdeD0e5XiKR9vy+u8HIlJ/AHEYaU0SPsyCmAQwe5Zlli
RxFmwMiTXYb3HnTXkegeOxGZaVT/uwCuRhYcl1qZdtkDbK3sa9sW0O1afiEe9c3W
sg2uuOuXcHM3rcTcmeJNKvWSi8VqwMDb8IG57TbefVq+buxNMCzeGBBEvNLtrHFs
N2m2ebIB3DEd3PX4psUZTGcteX7Z1rGi0X7/KU1SWim1SihKqF47Lfw5GuzI3wJr
bfuqI/2lothVmJZcALFsuSQU+laYrOnA8vtM3fodYEX6pKMYBI2nXdepvV/7wHqP
dpWGMnx2tSOouuDK9loNp0ECah0H6EmLF9Qf71MLtFc7LdGJOh9M33pWWGpWYL+j
E7RtgVfkeb+TCUPgyiWNNA5/OjBSAFMSsMKgmqeb2ZiMhJuONEHAhC1HqeQK8HEb
MYdf/GjCy/g4RLeTTO/KnrlkTHIKtY3aymvo5ejtaD5OpPWFo9i1hyIr+5YSIFxe
zHqQTpEz+/OVq2nlH8xRTyErun1OvTe5GTXrOkPShNkF3uyBPpX6GPIQPxxB+G+d
siYfyTEFNipcN5wh7l7Bqn3vqWlrj50vEDsMkFs30LvQ6bxHS2I+4oeygi4Sx9XN
G+4aTLz3y7hjQh2Hqb9nO+zJk+pLBl5WexO1FCC+ed3r6qecrVrZiXI20NCNiIZs
1JlxqioYle91XKGR1KeEVe5AvtE1urH/oIxYNfAmmSEr5ujvPlrzUlMt4HOnqbdK
8IgpURAv7k7Sgwsuws2GzI4nxdxygjNG4aNN6IF2JQPRPtrhDcog+V0iLtIlE0wf
8DIHREhE5xG48a+XJRBhicG0upB9uAHszvCSJGqYcJp1N9A3HruemcznHR0MP+6F
8w3xbjGfK5M2MfPbvUk4k6P+Fjo+6at8yExPDYZxjt656Yq9bIS83hVN0Y6oDHIG
8O1soKad2xYEkImm94TS4+iICr4LS9rxJTwg3phxJ57ZrNMbzjBYdMHlDQF1C+op
79c54pjntz2M4ZHzOpn7eXR7Xf8VOWTO78vMVLUAN6NZuL0CRiNtIjZ2TeB8Cgd+
GeyGquygHV7uuN1/ywAZZhxU4tUdZg3nVfr/2l5aCV0bf30ijsFyceOn3HTIDs6e
gvvV7SQNBTqKZuA5vfZKWpuJQEjP+GPbJrCWATqmMQQptDzqvL+yUQgqffz6uoJQ
Y3Tu35//kFPyYwB2cG/3MiMfHJyOp7k1vY36r9W+A++nc7H4VGUCdKDzbT/TlQGu
KF59PjJxp0haD+ZnTP9pxcXvQL1gwXQ2jMHmq1AFfBJPjwZYbaGkL014XBX5cWU8
yHVxrZVBdKmDGswyeJnm8xa9PhrPe/tx2eg75CmWfTszf8b3t8SVNbmHQJgS1vWj
wbvCfKLuOhVfyTbO5FBDWV23bBtdsLwZZkA36JCQSHH6YA/63ceesyz1fM0rZEBI
GvRzyb+8GL5Z8S3N0ng3krlz1viUBd0TjwMZ6nxG0K6rhiktkO6bNzoqCCGB5M8y
O2VSwuUSemE/YRf4Q0l6WMfoXRO62GcUeMCVhqxK+u5p1nvnMJdGgnb73dFnUM/Z
60/wyzWWaziOjMVKirOTDJAtzndBWX8MeHo9MvvWUez71Eiqi3N6cKYQUU+iq04e
CCDrKOZOHCbhpr497FVX6xPFzvK43Y4Q/ml8UiSdbVf3u9Ob42M7XJ+gCeeFx3W8
5olB2F5T4PqYa0uaieiJCTNGyQuwVQNb3uL+zqrH9UI1wsGQDFxc1Alx/61AqaKc
SQfFNCSNQXfLeGGA4QHWHcKTtVpdLbgYxaFza4geMU6302OCHuHso2RXY7LN64pV
1YUfueOebUutbarnQT7RC1niG1tJ3Z+p+Sdze3JKFAEVN4weNakSu02kzUhGE5b9
xuOmg4amykBLDCV5EY8zYELx4Xc5BXwZlfg672UNvGVaS8omw/yW2g28j11amsLo
5cuusdnwqRSvjupHGhw279Ijc8Hxe5YxeX3BtNiSoFjM9YtbJp/JhAT1RydkDyDq
RMIXBMHXXEVEdPWY+Hl13wZvqNtEoC/1VGKdy+vdqvE/kZeD3mzcjdNlzsI4PEAc
fTHHjSzxqCnzvZ4no8gIdgtelmuTnfUTZJihOeDCbiqomfBa10Dqe0QX3b+caIDF
RDfCkQ6Tlfu/lj3rT2geSWC46RUXk/RijVTlKS91heJ9t82Z5yR8fcvOXjA+Rrkd
oqwd1Y2G6KzDoYL9J3+T6pTbg8zdRsZdGUgdpdbAoLsy/Gm+mHLzC2UbpmJ57ucJ
aNUgRGWxEAkiazadrW1HWq09lw84Q8N+lOOr7ET+gpHPO8gj8rroEEoI+P1MBZHG
P4UuaSfKemxl6X226iDXhTgT1fJ/5+AUBf42Edvze5AxKRNf21L/Rg5Q83LferrF
YWoJXe9HxHF6dgnHuLfe7q2RTDQNXt3lI8aBLYPh7ZRvJM4bHdp8LwOAUy2GShGJ
JGwOLXZ+8R5Crgigh/5nHt+LtaGQchjMLGGhDtlNqQKiSrtcC7rkvUiFJPl+VVVv
nV6MGFsNgewEECNcE3FGA/xjmkB5rb8BdYuOm9yfwWZ5Qix2MkMgdaQzEMaPnfvh
YzhIrkSkfH53oWS4WsIvK1AH1z8OMQc5BI5a+RAASQN5TVkPXbI8X0OMwDKfm7AE
6JWaOj9x2i6B2AcBK8jgFP5IZgaqPqTEWPDyWOU8JYJf6tbmSXJxwLbqln9Tr/Pt
MuzzpAc4Z3xHk8/3f/Qcs/rEVuuazNQ2xSylaxY+TCF+ITRlmu8XSLd1LNDLUyWF
mN0l7dSCLjOCJmvPrW8VQjW0rGMtvLXFZcyhLcSoPKaq0tZ38ZjU4tGTr1HiXisM
xkcoUd4j9Go6L02dqMHTSqzAXVZOHpPMr+XU7tzMkOXpK2fm4K65cyyrp1FAEHnA
umevlP69eNvIgvzmoWdxd2MSuhX2enIVC6mmGBCiGfseLjR6fD0RzGW972l52at2
EKCGRszYp9dEMcRzCCLapE0cgBkunTxf9gk8Er8xmN0zyAe6v972Niqlpgfq13cs
pr88ks/ZReCQRDsdVsI1Po0oShOddQEG6LGQTuXX+CVtI4fUxi1nxPuc+CgDswYJ
/ImwCqILxcTPPGWLnENxaVtVvnilFchUdtnOmH2asMLCMxA7C6zYqa6vvwZdFIC7
RXeSn8ZmhGQ2oeJ5CSbECunMblJLyLfiYvlWbxq6UxDEle0ukmsHPxUYNUYR04eL
zYT9pa0F9nJg+vB9isWWI0Z5A2w0MZX0zHLLZ2ijNi5Wll7NgctYWUVIXgPYMBfA
eVdmY1/0SyZs5ldv0/Q3s3D4EolHpjCfYDXWZf3yXBGFBEKyI5OmFsLgxDwFAZeN
EoDz59RP4QCgxfP4VfefMJ/SbpR+PS61A/V1RjYnAtf9+CPlWac7hA0nt+sfcOZu
tUvMilpIBS7t8FBoTAajkTTopBnQ2uLVwIqkJYTFNyy42hvivOpYzrnOYSSpaIrY
nTvwWB8WZg34haPpPqXeZD29C0V1f5mSQZxQIQ50580Tas8ljLmSx4nytIY1nkrW
dStHQH4Axx5NlesKTycbSj8IXV83BCgZ6zs8Yp40LCn6l/7mdlcec/n1hJJLHqtx
l1E37UuEADWTKUPRhkfMUNpsccDVoUcNDImXCBlgrpcrER4H/FEPZIHwnNYZW0oX
T4jxEITZOz6kuWqI43BJa1y/Hzg8G7UFu6IU2rp9eM2R2jcI8DpvpESSs+88J56E
RJp4HelhmM6XvnfcImzDP9HaXrZp4DGcIrDJD4Emk1Sp5BF2GoThZuUX0uSUzS0O
vaMc6ss4PjVusStdpN4aFCP/7LMxNKjESVDFKwaHrfHAm3qimRJrf72zJsUgijck
AOpFXK0PvjUP51Wt/AWyfOo78Sio0+arlpqUFXbRtKDK4YEAQ3MsoSmSCDl9oyil
iIg9G0frsCwantDYXy/nfyKrZzTSZadaGyEJreg+SmvgZLEuyTuKDhYoZ4yZ4/7B
oOGtGRyURL6T9OBpJ4FVz56NG7u0V34W+M4DTtt9oUPo0Hx5W3ryPGkuyg+IlCbT
xKA2Jm89EebUwSEuAro/JNOIoOTrEYUXsJFs6LwFN7A2+mGCqC8I4IUPyQZ67bmW
Tl7zHGfdGlCa3uCRjNO1TDE6yXcAU3AFKrENRxMq3HR0fjgbxoHePFFpWx3oUkA7
eJYEHMnOc54Gszj83jn7zY7q+tdVB+G9E0qsVI0hJinKLwqv+OxiolmbhxYtu1Hx
dFYOkT4YpiEdhYHmpxs8w7MNewu7tgc9FY/4ZIr1+5SpTl3x1rvyO7rcbsbhR7e8
+jfwj/E0OtcbNYn1NisXoD+OydrUDkiC7HUsl38OceveaVeXKFlJM3Oldb3CWyyZ
upGUft9DjWwGL4is390ZdugWciRE1G6VcWDAkSodNaOZdaR8l/CgNCV51tJLo1b/
1vWxdZD2ureKXB9RfA4oSHFMOTRMNmqgZa2Oh2m0PiHVTug6AFgJ9JgDhdQZUr6w
YbArsXhCZea8eovY8P5glgkE/NRDHFnxZge+cg3g9PHcUy9q6I5bU7grbbHgyBW9
ZHVmaPZzrAr2th5DxixfoAgMOc7vm+iGqrlAtS4oOb3qYhdsViGME6PgWkkKfRp9
EbOIRoQBPY13uPqekQI/e+eJboHSV2Gbpavke8nAGBXJIm6ThYwgn1xKw2NWOZLz
Vjbliwc7iJDMohAjovw0hXw4JMD/UDwe3CTMD3CO6tjRlS5XKgX8dkuP/9KVzYPI
W5U3aowxON6sAV86Shuq6fi1hK90rPcywdVZqvZy8jbedpco8TntJIlH2nrJdMqN
ypS2EgMvwbuBNHhx/ydyJfkH+IU+RN00N+fJ5uraDj1zv6p/My/T6I4qZCMwgHSp
A3Shi8tHMgCM77Wn4/k8hlDUARNjG44bBPnIHzsBKvmM+6J0LzItxZrpyuGdeVRp
7cJjh9XjJyIAp8ozNXcIBdDfFolh24cquMR3P3cgf6qBe2jEehcswRGsdNYtoyQT
D5HuUFA3udweFbgCGUnyYyWYarGOAXcZWG0EErqHXJNT01vB8c94o07+9ObF9Q5h
f7xNuJBsSjYS4ntR5MU+BSnxy6Yw5ju2gZ/zbgKZh5mCcQrS/KTabTG6S2+HRIlG
a6hMLYjLhkasP3iyYAOHpWSQFJ1EHH0Y9VPZI8eGfu8z02Nu6/5jXJEF1+ogPdw8
/mhmskG3TWCVjJLwtKl9G86VmBJneLcVH9js1RWHRdAUacG1YSiAhnS/mSNP7hgk
bNgqZu50biEXj4V9QrixBaEJHuhB1BJCwPO8ZxlByWhxqQ1UlzWDEijYLqcui09o
cDQIAdo/SQzzRQhuod3nO15QJjtUQw3+70uOxBu8+6u38kZwfHrBaoB35gIschId
d1XbqLuG/sT5XEGYfxe/3pnUwj2yj9tSQWPIihGBE8mtH2VQqaseMS7zcKbxZXL8
7sJKs+I+O5vYzo0mB5KZyg77U1NZIU6jv4HWFazamDSoBZXD1v56buqYOhLZ47wI
0z7BqQFUnHtkJ5jFuV5W0nHi249/6l8HT2y9K78VR7fdVZDiH5IHFAZwyKKwnw7B
c39raWOatUyq6BBCd+yycaO3Gv/UJLXr6PoUOQhDi3sv+aubkluVhZgn7NrNgtpB
ai90S3NZdosAAHsHIWqoMGCMnR0YNHbiZm5LisIUhbi3zv1ZA45JCnzmubCp98n9
ZNHmeEn8tS7i+ucFeYzZkmaVPQjheoI2gptZPKeVELVGn/NCOmUSospAERM5L/1X
sGe8gcmGRiWUESABLMtPNREZIo5gaIqwL5WRUJXmFR7o0Bs2a0LJa1sd1Jc65T3t
ZyMmY0evq2TBJh0IaaBLHVkhUzWLd+ICKLua11FBCflIG5aEbsYcrLo9vFgm6hIi
xf4M9HCLYx40QjhiqkNXC1l0rpCD8DNIfZMH9Mn4eNFgkOZ2D/9PM8e1DZCmwaoA
TbDbkj8vFPrDfd3ylKAl/oeVa7vzIdJqsskxSdejJumbvpcqQQZH5nTrzhlH/0Kr
mqVhoey7OmH9S6jXxGAMrH6uTJ17Kh2gmXE+G63yid6wLnbp+F3J0+t15hnG7Gvk
K2J7Gpr+NwJ9T/KX8oehP3/6sqt/x2N5hGMR23kty2hzDMfdAlSzbvWnvtFCwb6l
Sj3mDHtBJiE14GbTEInoBZxJ0Es+bb8/Ea4etE84bqjPcnDT052vkAqjN9M4RZaq
QTOpWpDO5/mmMC/tHsIFAg43NWD5v7BV4fulfk1PrhN/GlWHZwip248qrP4/ArGO
9qtXLqS50FHmBMwsHUNfWfFZ4O9xZXcBMfb3uOE8BMECGWZd29BT1pikR05cRLdq
AkREHl+woSXOafJwD4yzo/komlpQ7pfcRnW3Glu0yZqlF45+TbfwxB4aw0Cf67au
oQ2LUNRWjo2LmxcomtVMBCEFHYCNoSEyS76QjN5UIJaoSCrBa+3kCFu6i+hlbXqb
yLA8SORFf9QTSoaPUM6XmBmOqiKcNpThk50gH8ff5bPxZXgLNx4cKfG/Uo2myzEZ
R6l6Pt442ZhS7jf/ZFJnBovKAEFT8mW5LBFP8AmS8RmmeEO02wumybFz2bJPQ4ij
09UrGmVCkVTyL4QwiXlIOfCNZyfMqzkrJfoFmLElws0mfBFm6xAztl3CXoAKh0LA
D3w7RGMmwDPtxnpbQ/CsaCUAETzclP7yJUVueP69TgAfMVffwVBfVq7djrxuuGU9
Y5yeYVrxOyeLo+fD8bQZGLJsV2KNDfubScDr1yvFh1BnZOuLptEk1JfjFpTkW0RE
yb3EYArqZw0mIQpRrWIidDlgqYFVNCQQuhZTn8gE6JzG6srynglju8dOF59NnSHu
ZN6emX/+n6giYdbKaahCnm8ML1UPYelmJPxGRk/2DARjz6XwZMEOvwT7c6dPbak2
abE9ILwD8B8Kxs/shiQoVeyIpgM9+wJz3ONdDGbjUI6FvUKJJSGm/g3efcqEzD9S
91A8C+r3/pDtlcoRmWOBAtHRdM5dYgmhRRO8NwUeCZ/vjR7PjNqnxax/NmNOw8nB
2kWoxtH0KBhu94DP229WGaK/UFWzTb7J+CbJnRxWaC7Nyimta2jnWndZ/ra+MhvX
ve2BvPmvEq5Pns3VaBgZ4KVomX1sVgHMMUXLhhU/vxGl5FYmjZshT+f91FHY/La4
1Qngv8+BDWaioT8dqgAoyDlKSxMYMp8Hr8mahpu1SV7wO1eEid1cwpv20ROmzN+i
2eoZu9D8xQMBWjtjTDYUdb/iVPGb2k24DhXwG9w882KnGhJDAP4XG2glRv/0sbD6
DvAVOhoRSRKq/nZnD+FildfoAmaXkyvTI6LHThnuF7b9/7ZZ3/CsUUBaSl5GvcDT
3eUVP+VmPV1Wl0qMNa8vciYu+FaCAQpUXGKpafIfkbn1/ED9XZywW3Ap9MzEX5Pn
MtOrUHlkRmESROJq0RtbEq51kezgLRE+4LfJO/ZKIjof1h1lnIaGjT0V0V3WA/5v
DvVYyYI6J+eHEaDp+x1b4SNJStGf4XY/wmv/j3afgMF1o5ofu9GfSUSH9VkBuaeT
1WhYEF8Bb4BdknfHbWwobRRhcZCvILIJYT7rc+FZW/C5dJ2WBXOV2s9GNR4K+11f
rIvHdZnwIqt4pQ2PcXX+paxDWwlwXj1/ir4Wayhkk7rY9sKBgKpZmldN0nwiD2af
d1XwSCUQVgtt6g4KxGpj4BFUNNwOI0i0AhsE5F5cLNZiZVJ7q8sH2547RA6AlEnJ
lcI67ehM2QuMIzn2JlIvqh8nZOvEECJQrY1VQcuL7iKBh9jQfBsGV0OPQTfjbznc
wzPsNGzS61sJEOcJs41Kdj+iSHiGBHKFd/4qCPg+fc6koDS90j0q9u6rO64rionF
plFjmBaa4KDf2qHt/nc6kTBf8+rdz6J6h9BK3AkHsHgEywuXGfGgBNP4ELbf+Vkf
CToSPm8UoNLUm1mDBhK4rnaKew0OW51LyH3tlfvbGcgOWBqNftORSOaLo80ZOVAC
oKiStVqVwn4DaKelx0phfatp7FwX6x4iVQGpTXInIpIKLl+Zu12e3toE3KCE5UGe
COnj10eHYaWwmfA192ulbmQGwDU4eghXClOiNBiEjc8OQnuDT+d2y24K5vEQBQFS
BmZZ90tySucvoT86CUYJXx+WGyDhmp33EQ0roQd8cQ2Ig1jUVHApS2CDFGSnuNHE
05aIuIJgob4o9A+5h7I2NPR0f5oiNbNNHMd9HviC0N0zr3glzuT73AGiYaUcVVMa
Xx7LnJmhOv7ajY5hTiWv7XE41HWLDBlsEAbeqc1H6Pd6DWLU8qEYHJi6CFT+7Emh
YHuEIsTYeLmkHwTOM09oAwti8dYUnqFaptM7vAq8LtHySppjZOsbGKD+0Me6b25m
BFqi9nN3FZTTr/iG4G7pJQ/RlCPlvUzAhNo/tNWArMK0Tb91QPU6G6A5t1COiGry
UOvjdJwwMdZcYbS3yU9gdH7YOSCXInH5yGc/VeJk8QoLfbj8si1nP0ZGj8MPOpXV
zXjSlQvFsYY3W1pznL5ChBQtUXf8avqWsYfnWPNeWwi91TO+71EBa6DLT1yL/WwU
ivM2goq4aNU6/JUVzEdH9ACpCw3hweFyDVjz3jPodfnElm2uZoKqCRbUtF++Tfxf
BWcY8IpNoruTP9166ETyUw7VTcAGCZry+3aG6ir/OjF66UWB8WBHkM/Olc93Tgqd
ykTVK1XtTQA2DPfT9LdEUU1yR5u/qrDBrwQc97Ir62vPQb+uvZNKQSh3ilVtQAVb
jDvJFlftnTgh/tuKIrZNsRXme1GdvzMLszl8qDYTN16mBlv7gBE2hCeEcaKZM7b9
UFNRu2ZOA8dwYNf4aUDrMA0FFSwkyx21EVwwBHgCuyYtTAM6ll1HQzyXc3z7c0/c
K3cv1mzcdW+gjQPfGyh47zE8f80AGtpgbc7/437bwjp3VeNyJ+B8+26MSdQl36ed
03OD48Vj9/U0gFRvrZfVeowUVzLPeIbGObtrdlVpqfT2A3QLQoIlTcHtP+AlKzSV
gc+Gp5HsNV1P5P86SM7nCN8rRtOqjhBGhVfijyDKnzc2ovmgH8DhN4oYCF87XF0T
WASAeMO3HuuepxBMiS/W4Mm90GvZEXsUSrNEQbUxr3AouVSuFz3XXFN9khwC/SIt
n9w9KDwR7jHzdgWiDWMmKq0gkNlyFGSl7ubS7PKnNqJxs+OP4JgliibhHKRsZpou
KfKiSI13ff5Ygyv9RyEKZSyPtVHiTAvzzCBzOAyGNWCmMuifBdZ6qt55UdMfgVrm
EKtwtxjPlha9xIlvqvWdtSPpZDm+vGOsDH0gjyYHd5xPfK3N3JcEf0dhXaR/1R1k
P74G/8I5fuccFjBzPVuyHx4mLyTDgXrYmVUePWmG2SY5PkTSB0nPQ3mE/FCn+Hi1
Qzp9BlO+8MsBiOMlQIbMvwnlIK4LEl468pmhAphnHg961/jg0fXVVCu65CZZRB8S
P1VvU/avc1vYioaXFIFlf4V+qPUpg2y8VqItwPQsnh2t3CA9tiEpwkBCxTGUhcVu
cA3EWFCu567aPRyeiWznTuVSHoB4c4aynaBTKAqrrCtrtDmvhsASfm+vCY17B0nU
TEi4xxUKF7Yri5/aLdv/txS23YWIK87neIRTgLl48ETOYlxOh/0k09571/a/oLRU
FXBrQsDdUXF06yLwlWxvRX+zG7l4B0bd37PudpNIGXSDC0wx7qmisvez6syQeb6T
Bj5J7Zf+/VFq6m9dgapB2hh27KFT+OQwAislQmURqY28XadwEY48u8CCsoL41EtV
PUol9Oo5xci+QW3zGZUs7ZSJV9KsQPtw+qEhdYzqEH/yfShqVXVhSVM28ODUj2Nf
oPN16k4VFIpwm8ir2Pbm7kBs9kSVxkSj05AH4tXGPnULYdl4frgBfYXNo1IRxhRo
ukn7ssWWt+RXMUSjjUrkMm58eEVozTb3n/xWcCPu7aB9Rp761c4FzjsMJ5oiFGeI
V6qD1XRhvMBAW0dNPZD+8Rbr3vDhvrIU3WxtvXlybNYfLtPdysvQ2ccsvPnusI4n
MsyfO3zly3/VA6pgS5JHYCEqFs21kcpYCVgTfVeRDudbkZzzap4MklwW1hpU7fY1
uyMv8Y/RndcOOQG9F8AbRKU5w/LsThhD7/PR8pMaMEMBX2LOTLIWZ0B4eeMLUnQL
i02ztAeSHlZYeCa6S2XVPETjDKDUndR8Jq1amusjo9GQdgJMgBeSYW9YO2CTJB+r
vTaRCFOrb1fWYBipTRxqZerKAgWrAiU9sNXqXM/9RHmw4xZ8TjS2AeYOgPciXG4q
mcp+uJ81Gx7itqbi4J/+LcPeScFpN8QhLDOqettq2J0nuEl0YrszSmTRm1hQ7V8O
AwGUokF26wBgO+UcNFFPBN+cWfhGIPsUY/hJWz1f+fosn7Iur8wT8MNTb5PdtL1p
ff0/2cQlJRnRbmvH/S02J0cw4UjwP/MHYoFHWXYPpwje5Eg4+ZI0kFcZRt4L9xKC
FMZm+VGbMF1Qu3MVoBaGlOu1lzX1rZTAuvEPg6YXGDDEt2Y8TjERxKKaZtBHozth
kUZe3VPTwJGpz48fVWV2l5HYiKCUm6FF6PJbVny11RLoZ59wbImqYAyDdf7iN4RD
nXPRWWLTAkl2Pku9amJg6YIovF8V2FdlWt18B6tabLFpq+lwteg7HbHuf+QxAZuA
JvsdwupZEcACuoL7znELZZ1yp8ZtkL/8WbKMroLhUL1rpadp38xUylQPlHvn20K8
ZoRRLsDc/gpMc0oAqcSuFWXMJNftMFk7Y1GW5gc+N9pVr6pf4aEfpcudynhsB24k
gYSwfhlta5i9KjxSil9M+VbpNhZJxfloRdwc4CumZOMPmiHTKbdgw7qlomKN9e93
2QBcC0NLx74KW5y3XruG8vHC1B7wh2Wk6WMQ7nHnKP4AF/L+wjmvaI89xT+Fyq/G
jJ8QTb/9cnEiplT0GW/k0ZiCpRihhxnwP30bKOdTXYeQWiasvFppHIa7Sg3BBMmy
2LaV+QhHbgdpinsUNIvbf/5Pi6ZIWSGu0mZ+BvLYvgSHeEymdJT36AtBjJNCLL1G
uIlzwVW6m/pSaSUvC/Ggvfv6Ls0bz2OlAzyvEOyNf4mZiWwXPIDe4uHcNQe+EMAN
5mjsojtgdYqU+/eHlKrunxA/4FfCeUfsgcrt3z/105xvxYVIfM8WVYFgt9GzKbAs
G//rWLWwd4Kni7qp1ukLPHFdVIScCltQZwFpvVjb/uz/qmqDS0hkLxqd4mODEjDH
lHcNac9rLcsLTJ4OI+uOp/6wgO6MebwjsHPywCUHUSsOh4MHrdXhO7F6t4ymgSOy
E1vIaTJexTBmESbNWxqs0VE6U2cyqJLtSXfjw43BND6tce2uemC7maRnshdisu2g
9Oj/WpHywNHAMMuav7BLLE39iLDEhHldv2q+4TFW1OHBjVEZCd6dIydCKl3Z2NhR
ujfzZpNTgjTic28hJCz1ahJhljiffU8KKowFKYAxdJy6qBbZ2q+LNh4wYoK91wuu
3Iywg5O0LsB6SBgSBaA/chppNhS7ATvP33pJsYsUJ6RxI4h7T6gITGyhzJwoBoHQ
jXq2hyiwNXjDwAHf8MU6cEgQiE63jFDBNycbpH9Vh0+vIOifiHv9NG5dS2Bcj1p/
OL2aHijo+PDGxNHA/UW2bNM7hdeLInuymzB2Q15/tifLFhuCtfp0dRI6OKNHdfmF
+EJ9Tb2A/Lev6CZlVUtO2ep5dueuFdkJ5OlfPj+BhiT/BLQ/V8ad9jgyZds53e/z
eeF6s9NXUxMMiCmBd9SayNGsGrwmNFqiyZeP2RGQE7qUiZBHR53PDJ/MtWfkWOTV
0PKHwtr6XYD+cgrZ4Wo38WUFXg8XUifT+iYpESSONtvv7yXKXLw3qFndkewYGCA0
cW/gNsbyHDjxOS1eW1m97wlsQmz8H0hrVQjj/FaT/+39dCALWy2j/ijv/W8820fB
0FZHby3lclXb+rv9Rb2sNWKlAYbumv2ACKs9JVHN+Y3w1f5gE13zek6/vd0v6j55
63VJTXIG0/KjwfBm2l42IeYgWG3MWpQgaYuTwDS6mdl1JGVLwVz8jIJjxj+GlpQi
0oXINVcZkwbkCox8w9u0isPwu66oMNA3KmbF7j3WTwJNpcSiTLx5Qg+7Mvh1W+NO
JPXbpNR4tHkAvD5rTtKko5iCfhnr4yIwDClhcEaIe2+LAC3/j/lSg83JIDat8RF7
tBj1fkBq6h1JFzgVD3Kr1bzHjwBvt+kCpT0vLQKpNHFKFVuHxfvEJRRM9WiCvYkR
+Y4qlU7yXuX7novscEgMJqPVzdt1aGa/ZRIGfN0rQjRc/ZUxfvrM9pFJIBJIwwH6
AAiYUiTI75rHDGQb3e5CdtUL+iMJgW1Lq4Avos6j5vP6G4OJkliYvUQJD+Q2GxBC
nd4X9VTcz2VxCxH3oKL9jxy0HcmhFAO6ieCHhaLQ4JEtDuqboXAyRFTgVNUYDeOB
LcoTi8OO0DMX7W5g09oiBJPAhJ77cKAopSXwhz6Fq4mn+LnZCBosHGECTVhM3/f3
TdIC9Bv/p+rqUlY2iSDohS2NjqRS3skm0RkH1U62fpb0ZHfXcav9B10RkbYLNOL6
20HqqTYYlQbEt7/04uoWk3HTzGVEv9tck+/bwVjF3wNGITK4QE5RlyMJY+UgDHxe
wwKowd27xnuGrlXehiaEW11S4f34V18wclnS/J6Q0YRzWAORx/uB8MALLbqK8yuW
S0Spc4zWKDMTliczUgQoeFkKlqqBvBHwwJQsK6bi9V/+okfYL/KznC2vOg2ypu/e
gTtEo2pQWIpvwg1O89Lyu6UUhQcAnjISEc4T8IDuyiOuC3yN3LoEV48MqsaO5R4q
3yuZJNWd1tfcAzTDJhBHRGUWDNpB1OHg8BBvuUGJGPp2neXx/4mzQHmSg+lhqIln
PuQVYZKAn73/o7vBCSnY+9h3dHPsxqpL4XY9sXbIDaQRzj2eT96UUyTZUh55pk5H
MuSUKwluSW8XxXG7jX4tUBRHnnnqnMvh1zgYc4kAfJS8v/WbhtuFikX0hz9MOUyC
Y8ONWPN+xSGLWIIMsH+r9KMfQ86YWhKGAojD5oEhCeHB63o+VSPHRPDAIziBOZmv
n6NVNi4R6+UeNGjT+xB6JDcVdwc0lXYMU5IRuitkAscS5xC/eEqQSP4MYCW5rIt0
2We1dXk/1pK3gGr/7EU3P6jA2q39nGFLQpcSTzAKXiHfJZJ9Eqj1uC7ls3PKP+ja
JjaZPOwgzx0D528T0BSHidxOiRsv61KsTiIN646VTpiojWhHEIUH6nCNgN/2Zqvk
9SqYpptHjxjKbdbzHTswmQAFB+NsfzHgfFEFuHolmta6lRKOvKhc+sMmEaX7Tji8
ClGYSyZcTMLJgvZH5Z08vHXM584LPxtHvDz8ybAXKronTVM5ghout/6ToppFPaRz
j40laONNUYx+0YUKHuDKx5khnmTYvyU4zFS+puIm8Ov5OjwEhdV2CKLXyU3u7dHJ
tFN/jZZKnrudPXMsjaNCnlobz5i+BbJZs7oWj/giZPlegYea8bDbFECGQw4JwfEr
kr3CUyJKsncX4+hea15IJOZ+Nz7XQMWGWDFQpLVvOItdVh6c52d/osK7a1eBEZQy
2BzEq0fx94e47PBIaGX0JT5bC2kW7I/usBf16po6yQ0EsOZfU3DJha76a/bbTWnv
u1jhzDTA1A7ov4JYF6Cue0BW4BZjp9G8ma3cqYRgkNsUE5d1AJZSXSRI5LajWcW2
yQb39f8TecWBbf71JOAL4GI7skJ8fgHiKf9gbnDgeAdpqnE6JP970CkTmA2HDjyl
122W/jEXaOOJRvJ7Abj4JWDdYMmRbyn0MR3JYbjpKNJLN3UqGstT3fcwtB8ZMyO+
0JqQxNHWNWZ1viTWCE1jFR1ZpE5kcnFPqPmHYexJQXnTcMh84LlwjkA9qvXS+8ym
Wtuua4BLE9TUDKOH1STk/PF6eBX+D4+9pe+sTGGqRA+rsrE98YUSTayWCGBTdSDw
umE8BRUgB9kCWBnQOlBL/Pn8ZqSnxLeVGq1t/44ezidrDpPeqcmTi3gCVEjYYjbN
m1Ewig98KXZLdW3lAaeWqPKeVddYE3GYAP2KSYRnfBFYehVWv1W8sBGD1uWgrs/a
RSarLNMmgm6zZh4BMxrdvm06iuRRdsfruwDH8yPbeIZCP3FjQDVmEtv+DV5Pqa3E
Mce5fmXHrKxY7mxoZYBPGOKEGQlrOp7GUcMc85eJf62HwTpWHKSRDq/pLbkfnLI7
FTqWIxVIpA8/5xWYRBGK/Jq9CRKNxU0Ck17ClHuBCdFgn1ID7Pge13HxFTrdQqYX
NtOR52hZBkJPtrE6EE/TyJQe6pCNjuBIKw2T+vWTShlpa7rauLrU64KMvkaDoFHe
Nlr1FxBl4FnxR7QQz6jpEGMYUdjj7t2MvNH8Bu9BoPf/ZPJTeNVGfLc5ZKBHPhoO
8SdLs9ZPzv+Bw1R/d0xPNOrQGYIN3ev7p2GwUmelzWtgT0qDMHmab+/JH8VMuPu2
MSkkMSUq28PVIbW0GxzyYdchqe0Xlu4abpv6Kr2SsqOO2GXTGhDK/YS7Fkfr4DMZ
KCgdVF8xNz/JOwYcfhz/3vfFuUXWxuvt8binuovqXKk1R6D/cRz9OB9mur8x53Tv
1a+xTbJILIOe1gfl3gvrJna40MS5TBv/XK+TyRJgIsKUFDlzGdox+sxDlq3JHZ+l
Aw69xNs6llbFS/Ttsv1Tz9SCfWi/IEo9gNPjDzn49jvM9tP9zlwNndRIUwjMbzBZ
8EgfpUIBbc7VgRY7ntGDXxw/bnarUjYHZ6n11M2MCV5xt9V89K0gq9Kl8TRG7boA
zb17FnY39gSzrKSVIBf5SbRfr1Bk1DZR8HQ2Yovzg8vMca/HYLZy9u4UgCE7nWPU
BYjGxTCW3zLmylBjWyn1v1m79dMDhh+ldU6ENotKsqC/34Sc0Hu2/IyUtk3V+hel
5q7DMFPWYBX7KWOljL+ScZCPQ/yeUvx6BpNYXwJhd/nvjUfhi0EaXvYZHrfpFA4y
qvGdcIFOmAyp3w95r2ruvl+zIm7TxoC+6HqZgNDOliYRZJr3yMr+vBYq5Am938k3
GvtKCFsrIiZ8FliTMZpO0rew5Mo2v+O7URDocXDcckvinwt8us3+Yx+dxhaqiVMt
AX8pSHt7k17YkAfDD9eWj+yI/xB42QGAPLKYvTCqc9D/MQWW+wtGkGHdvthJGlyz
9dWN37J5j+KDSYFHPhVWcFtN7Ajx4iqE/g+z2HQQ2xI5r3WLF+8z39b4OGb1roFl
Hw6yWWU/JrOJyCfvb2piQIqNtYlbQQ2rAbh7Lc9z2tvfmcZEze5UuUsgG7YUha0Y
dQ5SJ9r/72/jnh+qPthIq7/Hcm82o4zLnjzH4KkCLS5BiM0m2F0Uw8zL9OhVaSke
n0/zag8bmRw5eTEF/7OyHYxt4weZ7VLBfMRlV5Ik38PAF1LdgZ5at7JCWE4Q/P2H
3QXP0i2ExHS9EHTbn/shRS9sODVT0Syy6vQfd0R0PuTU3JwY8rp466XNXOXIr6I1
PDz9kQkRF1Eslrp1v+fHTxic1EszojTdiI21BfVLRGfXg6kYwL22DPlXayhGK4Ds
GcQw8IHnzavmvMjWrqFVMznw3Y9DfGPf0C1zGb/6OmUwZ2EUiICqQq/8+x1sWHfD
hg4Q255QQmfaX9MIJNGsNNwzQGNp7ZdKUcVmcbXJi44K2FjnC3AcpPM3fwMm3jja
/aoYsojqSBJmkXONgiupKLjFipy6GlNf5rapcHaYYCl6g+y6qUmgYyLUMtvEGl6u
HDTd6sv98D6RH55N9cPzLJiZSDMEDSf4x/THmTJa2Ril3wM2qXJbR+iVOyqo3OF4
Iq2sqDyQZa1vUMAx4+xVrS0T/9R+H+Jd/Ouq4BXkfii2x503P82U4BAa5OHIBZit
SSdrwFXAkVI9L8iToNPsjv05URMx8D67pZgAu7jOlVEREVLQQJjDp/BcjqmKroDs
a2JLC5KYxo0RmrPqnDmX/M0mKX61wfjLq+Uvll3j+sbOcQMKfxddj54fGMXQ+odO
MIqPpnWkDotyECDfffNJaT+P7TnPguc5inYFlVu8dI+y2ikts01Ffq7Bj9Ah+WA0
K4fFx+m+9EsLWfzdjiCdacGQDKOHZhIbCVDuFzSW/gE8a8xyQnPizFKD+09H/Jsm
Ho+TNOQQzWl7mcLLD5JFDH/7FOYyocw9mBt2qpV+IQtgLqT3yTrD1ov85KIqgViN
OYFKBYrXtyTvI3O62wrLWHFXUuTMu+RnNs5/y+wqRiUtoW44d87FvHoAjdcg3mHf
fExWniwnwGPVV+iuo/lniS4lMFVJbA8fFtWvX96jXVTuRdAb2JUxLmOkHEWzMtZg
4hNkQkNmOQNVAlsQt21sKNzL2vKv64dF5jR3WzUZoh5C3eG3N1Cyq0EfZCMbJFJI
/dLklLHyplafzTFSiG/f0EObq+Xsw945rO+aLiFFGvSYRoU7SGBTT80pVULuVBsS
IWHvJpwLTH+RGiquapZMQ5gixjKTlm279DBYOKiMWoyXzfE1s9ghqH7hDt333IWi
04Zqn1bjvU0Rm+n6Dq+Q/UmxmcYdx5LEEDI4+2ISKVqS3pOM+adItK+NMyGXgjIL
hmneiZ8HHTVEBO7a/KjnxV4lrr9wYfXmbx8BrIpayrfOeS+T2ZgIkxA7vWgKEkST
gTAELg+bSKAonYhPI5wC6r9Gtckrd3dUW/2KOPB+uXQ4gyAT7uHW0IFvKM0hM26A
RlJoQXrwq093UeV8OV7coeYfdtjowhwZ726WQIlGmAk7On5iDZk7KiLB8Xdnbnfr
qztmAwz1SKMl+ZKAX3rlEE9ayQR05bNieNqiruunUnRPYSrs1VCisI6bUV6Ug/CQ
nVdK+pNkhWDCKHfMN20AJnzdWNiDFIRfwKfcZyO9PCm2Arp1JqlUTdbTOhqHfX9s
EQbD3zPpk4k3+/zuMVbM/UPdBGgB8AEubyzsQ12BWaeGFdIFDj5sgHSTeQ4OHQje
ZgG/R9X7ivcjpSA4cQBIsi1r5rgt1hZFSnYLprqOM+MU+OvVDAKt0zcfIKuYgwLU
XWYLL1iYSwplo1HPOdKtfE/0+YjgQwPsEG6w8inhyHnYahFX/J2FOslTnZg/iYKG
xDxxgUMekkWuVrobS7fAWC+KsddTS7yuMTY4ybuodIrhVbuNoOt8BVB87ofoV4DP
aTMIlrl9aozKiCu07fd/I6Ib5MAt8UJYM1jKtBRcqVeY6Ei9t/yiLjPUyamkCtl2
qtpKnKJ/BKj31WYTZpty24j0mQwGf1O3OWFD6XVGgzfjcHfMnwqD/2H9ahti5dA4
IN7dzNvTTmBqYCJ6/n+Gfpn/mEPMuoRuywaNVgFL5UhuvbUSdDiag/bbZVJU1m+z
ofE6Yvf0fhQU0/pWhwsY640ExIAK0dDPqtcLQ/eDBv7Qa+dD3AW8BFTy3UL6jF2z
i3fMtJ/O/nl6SsuZ58qFEavYW2ROQOiihvwTtoJ2LZiuLlhGTJ0DHmZ+wLkVV0Wk
VjiTLLiEqHwtxauR6IKydVIWFtmr00MGvsH3bYZWV4oL6sPM93ERnPdipzVEniOy
MGPbgWRkG0pd3Yi4LrsSVO1PHFZR+K7a6WuY0AjPIPHVRady2xFX3SE4wX73yDkS
y374Syn24Q0O3OG63EI0VXQ2xPpfuWhmRm9B+dVsgEDBagTAtUbA9d9A31ZwJ6ej
qMFu/TsEQhqI1PPdZSfzCKQXrJTPD80cn8ya1OVbkvmn0VlihaJuSjwqEYhqijuQ
2/xiGX1pubLVQEKSsFroVhSI/tYi/MjYGuOICMccRAALIQipFkowtv/huVdxhSNt
xo9dRqd+Dzvb/TARnLafxOgm/uTMv+sNzj+K9J7GQIcplMwLn8S6BQNgyofb+D8n
J9I5wRjNgEzgn6Sgg2ozOlmub2jZ1Z+4D8CCtqGzfl9Pqd6GrVTcjEh5Svx5jjs8
JbKMOzfxu0081iOGVlLdVL2/RfTBnmYgPtD86ytfEBdZCRh/AiammqjDoWDWOhQ5
B+617w7eH9BKRlI5Xj4WPMMQeMeX3ulvnUMkYbFwB3fKAFyWjZktnVku/GBjGCBk
j1Pf9sYfWP/K3b+UOvNPo6oe9w6bC+i9OH88X4x7yULRHqpx/iXlY4OxaaH9PPtm
m5q8v+oNOK2pwFXbg4trsnv09Gk9nxoMbVDRFOIbmMUb6wxlaBo9KYc6nNoTqOVB
r4d8djh1jjjwfHHr2yVE5BCoog9JisSa2HPwns3vjlOy7Q0BDBw9Pkd9ZQEa4nnH
efWrSKXF45bG2Yc2M+GBuQWrypM69c95dcOnqV0oLsEwgC5C8cXl900K1doGqNde
6ES1y8SXfHH9sFb+rA/cgnyVFKyVIJmM5zxGvRO6aF9Qz4gdRJzPLB2ME63CnsHU
ixUyJny9n0HoxhD4BWws14riWocVoiRO/7pAcAcXFYgAwsl5TpOFI7XdgUKmSt8R
ZlAskHRdVRCiOgP9WieH0ZPaGJrXAf/1H/MsqHNXilFWy/Ky+xartXYpG7+f1VfS
ln5lmLgTL3ArdfNEq7DPi0lAK8tROQ4db0XLU69UoRXPpxaRhMFrM/ZICQsu6//E
LLImHX6QttrPsB1rVAzZEYcSclY85m8lZdF7rAtroOsIFi3a6baLP7keJhTW+SxO
DOMvATw2tRh9Xd+4BlkDMQpSKThnbnGnNkVITYv00sAOOySCKH9mxgrenwHG+Esi
kl+LuarLlTXU59D/a4U8BvAMKAAdlyOoa9MvzUgTR9a9RFT4f5RZ4tRNNmD0ey3d
6vkmtiG6YFBFZ9wS+RIfhpj78Wa2zg2cejyWchGi+4hLI8TDhyH2c8hNJ6z8h235
vnEtflc3SsGTa+XMYO5wx0pD5IDVhKs/P7QVnjkdZCmrIwNlj8WFy2836qfUpt+v
z70uzS2qjK3rKbADLVCAn3iqSojAKY73Vo20rJRgS4lZzPSwbkKo3FoG/dVwHZsx
8ymhXZEYBpqIZsg4+zb0++tWfnXsR2/9vboRibRY5iitkuopDr27P0ewEhtDqvgF
v2wh25ftORuAG7EfWNS8Zpp3ouGYktTsKUGkPpI0PRCyfPIHc7nU5Zm8yKiTMDF/
W9ZaV90TOEIFs0WWuWO/pdrDzb6p+A83E8PA/AMMtkcabfm4RbRPe2/w1iAXnRpZ
rCfODhJGcvZ161JO9gvYSzjeAzcng5Wk+wHE8l2TXhwISNmqrqWD8Yb0VtreRHLu
iDj3qV8WeaDxHia8fORwSPTmAplPmgZGOD7RCIQWGGh9cs3efU/OW376TJJU5f7n
Jvt/ivvj7tpaQKNvKLy8wrT+peg/knziCHT9o0J178nL3chndT1pDq4pZXpDAgxG
OtEOKEF7P2CCtaMI/0kGn5gbFQdmayRYgh26tIEYotlySHGi7PBn0WTOIuWYJTZl
IjyhXWq7fJttHkAxLxqkiJLbV1rccIiC6AADiVazFalo5XM5mEcm3QzWKmjqBTLe
JM/wFOFlfQtkt8gyvyxGAOmU8R0faYrGxGFAaqC1KeghFhszbXn7cvDWYIU05+C5
OefgSQJ8RvUPP6V+wulfuSWMBVPeIhANMoFgd/EKJBt7UFKhZjPeqb+qKvtBkpyE
Fq1HdU8rM0CrMwirYwg7RunbDts0QtWvNjLFuAVchKWBDJMK1nQSoHBmO174cQt7
0fgiDSjwH+TrS6n8nqQez0ThsCpOGCZcmNzV9i2Z5VLfFVM64DUiEoa/t8U+Amr/
Ci7ql17J7qtGD8ruemfICfkHyJ9G+GnBZhPpZyV2Eh6c/q3IvtG9lzwXaNouG8H+
fBaRRIYKjiHx1DUvrrOncw1pMDeJfWOwd0IU7+GDiMOjOOIWyzHRXEwIi1Vhu9TN
PRLOIDEmY3iw2SFVWXBSjETQPCKNNyBtKFhGsczlUXMppQkU4KEq4svJxOPu0Aky
OBNchYtJSUQSaUSP7WzaoLOP4KwuNufR3cYBtdork3k4gB3RXZjFdaHKtl6sJ7F9
1OoxSxI1LlC/LEa8eQNmehlG6gHoAKNyI9AEMI7D/IOzvKSA28ZBo1Mri0npdFKj
HCdyX314i4/yJTABZLXBOakr69hCZP+5Wu3wAncNa4SA2gBwItzPmuDZI2j9w3en
GVekHKgHth0O4Gx9taebPngtQLXF15VMqhogkE6xoLz/FtxunlPV2285jSYvx7Pd
rnNtOQTZaq3I2LNTnDvS8ezZOsnSIpcjT7eNIDZzPzhK/iA3QLMq9qXOvKBgR2UM
X25zpGrApvE0fi0uEex/2pgUaCZHbttN8JXcEsYopxdTAb1kH7b4+ENCP1BmC2L/
tHjoJIYrDWOoRr5oNVRc829DOX3Jq+dGs5iazrHmNSTf7QZKJcy8f/jAOxByzOj5
hI2CP9nLFeWD02/gTviyUJQw/BPwL8/9tJIlNKr2De3iOcH2/mWuGUdyqAxpTtBz
BQffAEh0WxBKI1Drl3lKVp+iuIBHsV4FyVHMZpy6pA4TsbymHIB6NnFbgrUXj9xL
PI+VMLjfySyVGLGa7UU8mOroeYuRlAjPE1yvKjDkIfQkKAswBo1upj3wmOpuHbGa
trvJcwRkaErzlI/W8434Q891i7Iu1Vp7150QGZP/OXxPUfqFYPWhwpt4Z8kY8KCf
f9vvdXw3TTXNcdFVmQJ+y5cou7BovK2JK8SHgniSykyR1BlUGOeUcOKHBEjd9WgE
HhsXEt5aknO5bTwJ305Q8B8S9KQ8/OHydChzx4naUmay9084NphZTUBYgt9pxiZ9
UFabagflKHTAGqndK5jXLxOE/xVrOjoaq5+lm+LtM4u9tNWsAQWtPmtxzDkiWnic
QRRsxYnuQjJUyYvH0pO8A3T+qn7RHLjk7I/3GKiuQB7Guh23kFEEo2nllVRs04JJ
zpP/4/7ypibglBOjEJc8PwCqyTSgZKcA2LtkBgZSZPYZ8I2zOYA11Cm8HnMN9FlW
L7EgWHE/EprdR0vJsd5hC3u4LPCy/YOKFjBDP7z5i8cEdc+YZGncirHsy9r1Lt6y
aWabXFlT2/RJGrzwFLvhpQZoso9U07x/QxXkTmOcPOKZThbYDlYPH5HHODIvn3I7
B0WDCrtM/TpfI/gE+iR4SKxeynaOu0K3rZTnEvFyR7hFpMMx6Qu71Erpf3ZjwZBK
D8k5PDp8lDjHhvAiL95bavK7mosjYWSO8ZDpKuoSemYL/8/yi1iUqEYKIfFIAUpB
cmvcq+sXCMEF9a4z8QZB+P0fQXf5rDDvWf+bfKEdiNcMV3C1nsB4XcXTjV+o2GzH
ovNsthKJ6JBN2QqouNBQ2Rzt1r6eJY64OjIUhrac9GDkR9Gw8HjUnTlUKfqXqBU2
iTX5R6JHvWPjYRrejyygXPZOOHOXafDdeugPDjUXbWrWGpcP9f9Q14/97VEHrN1N
oBeKyJlr7bMxT8l5wkD4zrwNz/qcUAkqjI37fyAz2+s7hLpRDSi/JaF5jE+z2THK
F8u9tVrp6yzAUnhEIi55yq7PlnCjf4Y+2NMEV9X87ziJG9R8aLUnX7dv5IDNpmOY
sifsyB7MutzKuwp5P39CEmHq9MzvSyu0IrogwMPDvcByPKDRZepeSQ5JHWX2sUyX
1NmwEWd8mJ49GVXXqTBun3IamaoKN2TpXZvBGdsZx5ED/qwYsH2nRRfchBwmP2gC
t7I3cHWT+Fn2moeZclzBqOzhJc50pzECESV06wJoHeUPXRBuiSm7VOXuzOM533DI
fNQ5UVAJJNoUai9cpBLv5WWGxoZMvlojwGaDoD/r4Iqu3DSdZAh7TAhkjeKolujc
XtdbbAtkFbiluDpj5H1mxZvjOss3ndPRZ2hCGU13zGhSt0DFO5shvAobdy05ExdB
FveSy/dTZM9EwZN9EB8UlwrXA225pWRyLtSN8egUDcekvrQCEG/eD1WqeeuXjTLd
0vMmZ3u2ZIQaAsqhkk3fXbnft+9wlfW81QFuoopLtX4sV2uWNu2Dmo8phxq75bqa
+SoHuhqf4/c2Q9s/M9iU6upFF9uGb70+KmXp4tEB/PCdpC/RfacFQYTHhqWDnOgK
Eaji+IGGCXm+DIxRC03gHOP+LJc7hNLkywoRPGdinIuxONfYqw6cYvLh6yVIdTNp
2VtK++m+bAveXRdRAu0WPE9xAJuxEtASdzviQfbtFtzpTBCCfZoCxewTjImu2Elz
fEqVpjR0PJ6x/AM8IR51eAqaOKlU+565HsPeze7HroI6yZjO3jAJ8nx9WbEkrs1Y
iC9eNnhDNJ9JN/EObaaQ0ZQxil0raWGol0mc+dBDWu/IBO21ZgYdJEKxCurJxspx
ofDIUzH62IhzVyl8wL3gEM3fHyUXV/n9+QUZahR6WwO76ybHb68iJsTdmMqhdJfZ
uHZLqWph7QHzEWUejiePIyEupHKtF77rn4pFTMCKEXuxdrel5N5Cbual/WoYDYWu
THRoJ9aqgHoZZuhAvEmAHdhg6McX42GTWNsa4HGlCkxwzPtOMlAs+X0RiUSaEZVl
o6vw3Sk2EEo+Dg9HP/LlxC4r0BrTwnnE12jBnwF7iBE8iUMy/yrqcMvLgzsh92rM
B590Wn3YMEx4tI7vUQ2vv9+jnusLKJQC7qfzKmPsStKSzvmGuiIzN5mbi4UYEWy9
lyn0EsEZ+RzmahCcho20yn7qqh/nemPDxrD5NYxk6pO4QXs12RxL3wyVCaj5/do7
ePo05wNfw7Gk++MewMPql/BZuZcoYovNb4fQ/2BcaWp3bAdp/sFLCzZCrACbUmIk
XPh6vApNJRQW5lBXHDr2RAvi/BphYuIidJKFdQ96jWq8XXfdMHK6XN10BsrkTFBe
GrkoBw0fPGFgL2GdvzZ0vhVu40FtY7QhjAiHlQpoZ4KD+3+rXpVVpb2eRYG2FkTM
42YfpA6VmTJPDQ3eCQIaz6d11kvsYtBXyDWIPMvGg9w7GFbKusjfIV3Qcyi+YiX3
t4okpb1AiDfNd2yQ9nlOAGnhTlDtdwAsRcXwp4tXnoF8T8I82uDa0dluOZeTJrH1
HqDSacPOq8q/UsAr+xL9E+LKwFNSc3S5A4Dm4gT2RRgCP5xxW4eCqNXxke1YiYrE
NdTbkn52VnT8C0edkQUu0+YedUAI72RfFCGhScTwW8ZWueNDeldczfEJ/dGWJbbm
xGs+JiLhQPLmw0a/+q0UeMFAEcXSb+hP4mFWKLnDIdQOVVPv5cyfnrtY/tSCiFAA
p1q+bc2KWBsiS/E+QMYQa55Suh5XJRvp4N5dlLEf1zlTij660OC5Eo3WaIFaYgPQ
GA6bAuEZzSW7pIYNz5SBxbSdFX1q0ySHqtBHIiN+qRfeFc3604LPSCWWfDDAqgAb
rKgNe6JsAn3pMly66k5sPu5cN+XmqetLXTy8o8EAxpyL0OZchFhv+8pqJLPK9gKb
HgxHVRLAHx2SvfoxZoUr5heSUUzRx7x6lOpRA+ac8WEQMT9KPgZfvYGFpvR+FhE7
3qKx2MZD2EdCD3otfm6+8JmHE2wby6zP6BGDXmqzO4+K6QwSRZX6ww2uiUVVofOa
DSkZmMeYSZqhiFGW3I9fR9sUMxK7KovymcUfsKz8OXtTeiQt1etNxOIb1b0t07ID
PP4/CFTaDxjGqaiKnfUQOz7e+At3KCVpyF8JmUPnhQn4030TFctc36zhvH/2y9rY
7W1cv2qrSUWrkopnDlLdA1rC5dDkjSSeIJzePEqfeLJ49j8HhmZzwuTES4wshoVc
ZBAw7SYw+C+eNGlTEZgI8S72S3w8AXC6Js8abrC285zzqPbzg/Uf9CbX/Ni5RRlZ
h13AbXzRboAqjjK6bCDY1m5UGH7bc6DCuO3Y6IengkTKHNbgJF7dV8JItYrFYjge
KxBEPpe9xGaQjc2qfJdeeFvaTT5Px0EZbFB+xmkuysWcK//DkN57Lhvgdk1eX2IJ
0kx0OAyghBHMjM5eKId6Q62sM5b8YFcLp8QB0UbxP6nIxK541MxQmukxP/UHs+7z
IQ6FBuhykegNcm1tr438nUx+aokHPIcj1qI0rbiDTxP7iN6eUqa0YozT1RaVXTg0
7kaUeXT+TTVp5kF2FqV40BCz3PLMBjsSMhu6KtKaejAirPaL7HMmGxe2JN1oBhda
VnHpqvqOof4wFMMbK3pIuP8L9G6ZuKwqYwQA5H05mAtp5ofiK9N8yrH9ZFZkDiol
GLp/aeMTvmmLIUXMVBrdlTWlhrzzBZvrMmoE8M+BJat9GZoErB2tNMypA+GT6F/b
syyW2o5t95yKftumc09xiFqwizjzQJ2A6jjy5c8NJ8GLoT9LI9tsA6/8wpjBrqc6
lhF/PYQeM3zdGCqTVhpww3TKxNB7fBwSHeBKTQaJiWQvPiF1ff+M4Cno4wLUO80Y
T5bhoirHMmFbv40iIuhuwIXIGO5YBbaWVlRNFJ5fcgGNF6ei95nBian91IVXgP+B
f9XYOFvkLUsvD6I38EHhzn4BxJZu3pw3rS/jtej/kLcvz6l95MNwom4wdw/pHG+y
Rt3HVhNjDCl0ENaBLHbtNYDgJwFF0dWrv0K1AXV7pALrfm/uyzVMyGrC3hqwJ6qr
4zs50Ao59qJ9LXHInUIRWSL0PV5dhBfXzYhGri9RBzXgmDAh32blg/xq0oFjBADH
W0uNeULrkljg9HIXBeWpkvsicBjo/nvMdelqGTmUT/Iv2n86y1tPsFkQo5I4G0ID
iR+/UpMwS+oqfPJJf64OLSPxiLlgiiiEm3UZWbaBzeNmyBwhFuXPgZWkrGa68gcD
glviDvnAmZpPMU+bwi91SYQsR+//NBxWBXO0T0G1bKAOOPlxOat0VN5WnVEJdU21
h5GX6clQ9sKWvV5nVCQPmfiXqNymtlUDReo+gknHsAjgNtaSOYfGifC93xnso5T9
FvE28xsJYPCvjbUjhLJyOTA9XzC0Q8pPa9IQEZbN6arh/MGTG3Oui1O7Crc0CONI
n8bTp8u+DQ93zmLnJfYCDa2cNXa9NYJ+PDXqSKBnLs/9h62mVQmw624trm8uk4BK
tcfD0dqUHgunrrJ3Hh/5KxZL35eLY21sK/bJXWUJDDozjG8YULkWQYFVlL8gShKE
ojh39DBa46QODqYOZaj+txQE0BAA13+S4l8uL+n006OCJ/zNEWL/GTQxCZSGFPa0
2W/Sfm0Fglrff0+4UToDOpkJ0PyBgag7uEMXjtVRqt9dGMcykjTEnUvh17aclGtd
4bMhIJlIqgXZLHkhG0Q6mObv2IQDave/JEK+tTVLfWHFRzwqO+ubDbhVBi3b8y2s
2OrxOZm/WaGr31fVK7SbI8ncpp7D3Gujuj+xeGX/Jx4kFlP4SWWdTeOSKVWevgur
FKb4xKGyYSu8TZz19o4QAqz18L97qpM8CVCGwYq9QnV6/97b3nG6epgP0Cg5M+Zt
wTetgO6YIcrrPHc9uQD2yRdHCmXo1igWzWTH5uNZE6C9sF4Yi1NwBTQHCfm7TmU3
3ETHN+1VzSMhZr7xUEnfagXXOztggEjiMqzT7iEPrfmoOZH+GeUe3WGGrK8jxr8Z
K3Edo3LzC1TOlGOZEWtCSpffZFaxAqh6I3EHLJEKnZJlI561khxk+3PU9kJUYv9o
FLz+lIRBmW82vVfJ9+V+UaAfheDEzquId/ouMH4+FKyfYK/ZKrIqn3PS8ThrwSBJ
4OSRJQAW0G+FckRR5uS+79hrljYZizt5lSFyskHEiOUSOZo73c8NIsP5M2pufIGq
vk790C0/OkkZz0zMd8VSUYbjkPTXrVsQ9sGVr+7yjUJi0DF1GiurpHCuMzo1IXxW
A2l7ZhsyTIzs7ppCQqYiCwu+siGN2pdawandUyrs3+JXd5z7kcji7Y5YOm72lJmW
RIAyVcstoS8lrKrQ+SC+kU0JVNpED7KmmZR9+a5V+hie4r61A99ArtwRl/qMxX5i
0TLxnjhtmenBqr9iWkuXzgB4POCihqOmtYmr6PMURkwkLsqMN6Xk2SipctOcDt1c
vBILrTQgL63/c19hUwQIMyh3CwKXTHFtnTUxOO9fU25mlviGnwOmZpGQGMS0GZ7x
XLidy5iLDHnezh9jxWh7gIDZ+JKaE7DGshxL1A259mn28osO1SkoIwATdogMYsVe
+1iyxJjsAiW+28mGrFi/+PdNzkFkj0QyvYrLDCc7L39SIbkOCJtjdVRSw5078ElV
qaP+eLd8uYSpsMJd83D2XeMOWdbeMbyJ9EWvEwjN6U7pMn8v1tX2gyhdEkgLjD/4
hUsEIHFBadiF27VDZCRocc3kDCM46zh4cjqOwZ3yGOB5AJ5CMacjaCMr0MZ1HfeE
hQoB2CW0PR7Gy4oCU1UJYJq3u/NzMgMw5l8ON3InO09ZOBznafkygCi741pkKwyl
pPT7rEY0XPhBOtZ5K3tYkyGtR3iXGxeeetqkxjOOW016EnSBEcmt/pVVLG8jar2y
/BUQSfjEJE7gmdNUunPMpt64AwVbFbgsZzkXYXE/fGNdh61NMJ2pOS/KvG6RvQOR
NT7q7oRCSOVTdpzvd1MdFBbEQEuptA1Qgce5XJgbrzhg5wsmUNg7/opAVrKsiJGj
/a5/Ht+9fSqygfHfsCBhkNGy2jbOe5pcdma6VLxCFu48h1pY2cDDxU5Q6LQOza3M
vVTn3gnyXA5Zgd+IrmI1vjnceMDCYI9Pp2QdNuJsdLnP2zgco3IWsvKdI2y5VjUu
I7YWSUzuFJl7rNyZKVXXbiyb7Ej56WZedYeX4GnL3HfqjB9diRAw2zH6UlyJ+AEj
kIZlTwtSiCdohhIN0UTNnVX1ZYQFIhmrNn8QR8Gzje7Ttx4ydltLW0tjq54swxkp
6B8lVGmdhJ7J4u1mFLnaQq4BEOPwAIXSLi1srSQsWn45kSEKGwkPmZybzIvJG1oo
fyerDxuO18ucFevZwmMkgWtkmTCUl+gADmdsSfamaxAaQixM+w1j1hT61Ko0xAeX
Mq4mXFDEBjr3QV2c/6qP6ILlHVVTlCzgF014+xrqoce9MmrdW72oYQlKwA/5ngd6
uM63tP9E2bdMcrFVb/1iPoKR8Z6hqme6Tck3uNCA4+TDzE7qsASwoIGITfj9akRi
mrwDqWTQWE93tIkgpiwDlDpXXfz/BAcE72BZnsOem515PvsOzYPAP5xtRrlZ0/Lc
d5rsOys5xrJJ12lqXYAYMhWPuktljehpf3c4lp1oL7W9C6ckQNkXB6H6raCZ4h0C
xN6J8Q/dh8/HdNIWeNFGTOljmZ67ST7fyLe+uwjouz80NaguPlmhniGZxDLgdz0v
5VcaNcKXq4M4tNmtA7/Htt3jfNyue6pl5+2e5U6xmhPNhJA9+GAOIimdUlIFGEm2
pgVwylizMdo/rs+/6pZqjLmkoyLxgw1Qxg30v/U4YhQKGMsomk0Z84NUh+oUg0ff
JpMinEuIDxu14jRb/qZy5gjHLlSPtVVUQACW3vFRSrMtXPGX+NKo2YXKjWCFgrc0
jEa82mVBE/l7/wgTXuN8QiHLcx7MtMjoWc+YJUQpOpLN7b/o/Eorixh8apsAgfB4
UiFc3oR0Yy+gbV5vY+gTqOdlY8t3JVa9SLg40yvi2nmnk6Q07lvsFdbGAXHbYekh
XWLsWbi4WsqQxhxivkX/7nGu7Dkhj4eNyCxsPhQ2exw7Jamo23kGYlA8A1UqtzwW
rJEZxnQa4UBN8BOIZRWb9dJmTPb1ohwNLg/dhR4dBTEHrFepZR/i3ajTxNJADZCq
rWmvx8T9W4JB477dyHN6gm45Znhdg0OnLaQe83l7nkufdASRWxVg6VvwQ4OdvCiN
ASJazDMPwGWr1KdZFgZRREJ+mcjvIxD75Eov9my5iPYwGPmurYpogUNoEpF6DR+h
nMRVvysixSf9Z57Pv929Q3IvH/VurQsTinABxPmAkFHhOh2MlRsJ7gnjBybHUQHa
/TsgecnQ8Gbk+ATe5gm9R1a/g9WJPmbI6hEvRJ7Xf6PHPaXhWXdtVsvQ6TzxyU58
bvuEAuz5xCpKh0VJLD3Rhe9aT5QTmsO536T5+r9XGRyig1PwVr9N6xMJXES8Yjrt
rtmrchWae+DO6iKdqDkxiiAtTfIMlyE48ZA9ewxiF/e3gU/ohOttyHuJEqH7Mx1r
FZfSmh2E7rebRyLGoSgonWzvx8WCKxUOCnKp3k0EWayQMDpBeYLdwHP1PE5RDh6p
55gVmnyl+SXR7wHqTXMA1p0rXlXDFlxM7uvWe8RZTyaNyU9f5fTrHbiCuWdCGfH2
rT9v3SdWQHdLu7qj5a9nlzq4bHPl+cUWatSaV/slC1BucSze/w2cIhElb7bbcpDF
GrlvdrNCT9v0MuhbFPrPLDWlVi2Q6l6rLE3z5RDYApiCoFuOb1BcRq52GCP/79oF
J+zTfonRa5kp91xljjyuX/7392Mu8AVskiDPKghDr+0d+fNwIV1Sa73bNOlSAm4n
rM1NCMNWDCDE8dRJdx208+fRcRjvvRCT9Bh/j6t2SLAro5Mi29HTI7hsRl9kELQy
lU3WAuulciVk+gb45PZUsTydv1/AvQG2G6Pxo3lsMUaT/NxMCWizltvF9QLLd2E8
EueQ+MLMPFKGt0JBeY5u/P9rzgiW+aOQ6RvTVigD3S8k1e95tIZMbUaMzPTijprv
ukqAVtinWJM8OZV/S9w5BP5SWOOdZH/4LHR1sxXsiTxcLh2WsIbJvVaie/iCK/5s
4YoOPy2yEYSI7VJbI7HV+kpwJhZKcgd/bgNUpvxi2C/YdTz0ouZmTAn43uT2eyTV
y0ozL7l/Jv/7TeL5pMdGsiNlDyzd/P+5mLDDsscR0bHIJTx4rQJHy/snTbnxNVBx
T3sCG/Zx1UZjItbl0+7r86eXhMq1ye+W7EmsxHMJ63XvQOu8RE1WWYHMDR9o5D5A
7E6S3GLz6JJhDbU4L7iEuwQz/aV2rzk8jGTW3DcBvRfokw86IUcQoFtKHebxpIiu
DeF4fHc7WGsuQ3KXN1Ob1xvwf6C0y/r0ygdnQeOmXJ/mQrnC/wbe5Vpc8dNigJ+d
p/I06vvOo7tN7kEMwDGsWfsWROvfYtWGpp8t0NIQw8ycT07gATe+y1fwg3XbGKmG
rvnTaoBNOxyzbOqp8ZohiKLGTgE8oYAhULFM7vM0GUlYXvVubF2oYejwGiwcqLDz
N73fs7eFQCu42zBBuM3ChCxkpiW1KITEEGXuYC2nBPpqTIzG7wvNDfPf0kqnci2u
aOuCM7XMdbCWj6N8kvxV+KPSqnYNYZBoavOWiBrXPHkfS0ZZ8UqXWefh6M67Iz3H
u6MQw35wj7E8+YvwR8KAn/mjKIxvdyQpX1nlGXchPc/K+IeLGpxeErYpvr7zmmWW
BoaGTmWxdMW8UwZTDn6M7bj8+tbSEzv8XfJoIHJSm9geXtm2fjMb/64JHLYBVrDX
9MpC3rmCvt21+U16/ZmaEJdfj5WL3scUD2rhpD/n/mpoyGasceUJi53lp+DZ/RUk
VV1awyCUj9YPG0zBfOdBooXvdfwizBKsOi0z2ZHSlI05Tn3IKMfqy8b1EFcJ1MMI
s4OxKK7gZ1p9jRKx0yfpfqWWFAbduSLzP7epznZIKInZuxlbUwZM29/rrknwZ7tw
wxEpJpBtSijPk4P7lz7rO3gEBxt1hZLerHoNDmifMAo8RM1CUhjujB4P5tkvn2ER
WDRQVtyB2Ow5tuyK4+53wBMy5NupQ/cbyxRPvhk/CH5vewiC4+eFkB8Ae0h5mlbx
qJQjjqc1vmXHkLt0Jf5587Q71e8rL4m2C52FhfrJV65Y0+YMW1slGYk3izp1Q1Ou
Gwgva3UovSnV++DbjxE67lwFW0ds1vVM78UC4Jt9Pfeh5zm7JtckFWDVER/m2tyN
cKdMMhQTb1ItC+Po9XKRRSBwNIR7II6WhbvjwFTpSZp5gFCnJDIM/BJjCFn71wjX
7AdJ97xBfHzJQjRmJM/0SAYEqVyVmH1tw751SpGkk6kOk3GDVRE4sCe3s1+kaqHB
rtcwM+l8fJfKrtXACNx9oEL2qGxEWrmjRJReP0EqLNgvLHw8B5sCBFpfxjoPwtl2
7s5YJcgPBinJUuYUgawooddteVa5e/By9B6fk5jZgRPzH5R7/ItPaMbQd3TJodZ4
YPBpIYtVt0CNJlUywwc5Y8MLspZkv/c8k/If4o6fszIlukQBuNyaIxDh6aPAMY1Z
+bT+Nu83VKUxuHCeFbRI6FX0T62FkRbSGGTnZ5FzPaL/2n8UiZV9502LVzRWJ/8f
gEhASzbcBbHOVHIf9HfthBtnLqfonQbgpAX/9wHnFh0wUpshG1AcoeJ0lcUzGbEU
5SrDk3iMyGimg2Nc0X9T/C4CrouvVaBbCeuf/BFhOyl6nBTH1w5a83lh7CFNn6ys
VnTM8vLUtGL/bsnZMTJfvMbE8TSoJOtuH8DUrKcR2sf+ppEkiptp57Wa8Mmlzvfs
Ky6XYo9mI0d/zMKu9z0AnnogZfpzCHwtPeYrEB9sJOaefsMe8G/7OtR9laRWTqd1
mBugYKRkKrZZk3GKuZ0AiFI3NHJfJRhk+WHRYIjj3mquLuq0EyA2LwdASloY3qJF
gTXaBmKHoshr+cgH9cpHrzxoO9bdEsT6Oa0gRBkcRQHMVKSpcItefEFVbpsYyALY
s0rNFeaed+m3uBS4WMFKeumnyj9jNC4hET3iWVgz/zcOlON7SCPCxxgK+xgkXUt7
gZENXEDp+liXvBarLUA0ELaJwlEy3vVUEZOGGPzHcS9gZEjCnepYxkMiSd+57L6d
4dxmCac4mjedgZB9snv6kQrMQbw9Io53+qtUVXLlNh6xLubi3fKHy0YPoDXair9b
YlBXmD6ZqkKhb6O2xt8DgG79rz8oG8HUk16ihrUkEpvEtf9QHvKOq/2MlnJvRArA
pIi5UJqSj3TKxw701/9MCfov9rw+u4RmGGCUGhG+PGIikAwrjGtH5bhGxUb1PJyI
pMSEqn70nNHTLIrX5AnzajBU8ygBrJFD8xKFVR84HebnbNAEM+riKG+yBYfsTfZn
xvDDTaEeRuPMaeBBPU80NlDSDyNeQkBNYb87pp7458anhdLLZFAxu/aIU20ZGjdi
Qg27iXd7mZA7+xGkAWhOMOHkvjukhYHbensVbx6vOX4XCMmeiW/qozi3J+79oFnF
mk8cBvwy9LEfjux7EErSk3UI5T2GmlnT6ljHdzp2xIdi6lTCK6Ui4F2CGdAXan+0
fcSWnT8MLsjj+3sELycMkhSI7Drod1Q6JAboVgeyndmvVKFMhuwB+X/yaOrQGl6U
aiReqXhXwe6TBOeWeZC6CyVqkrx4p084JrJsiaZuy6WmWA2WWisbr2vaG3b/sN3y
Qvf7i3dlXHev5FO4r2sXGH4690WfVgWnykVcWT8WBDTSluuta1edFpp+nIyZpDih
0CM7i+2SYzc6F+4zdHhYP+cUtRR3rmw4k0Op9och4W+8cf+ftK21gx24WH1gWwdU
5weD+NFYSTqVYgfDEOM9a1T4kZBdr/Grpse39jgdR6CvDtnZVcAJvqFRUG/1ABhs
TrFHAfGY4anIWjPKLqM/tWbdZhhzOpx/kczLPipuq/ZYWS6aiZwpoO97WMoRqRj3
MIgx+izuQWuQTCfFg18riAv/ABGExiDU7WtAvL8Aau9YJRZcZGd7NHB//jxSq4rp
A8Ge60oxCdO0sayMOpOOmP+l3C9P059u1PSGtIbIt010824AkrXeGcBskkWe8DaR
vmjLNtZ8FPv1BhOQckQrZcIlwNoeiC87fDBJKBtiM47Bk2eMufajeT5hoP8stkE/
hMMI/n9UGZi2gWmmmB5AQqqpiBhIM+wPaq4BPLM7XNIGSLntHZJcN7U/39nP0At1
C4TsTFq3FJ9/p1eniPyy9jnJmCn3mU/IAD4fKObhEsWOROG5vOh1Ego3KtYFv5nP
+SQcsJyfPb2OC+nP5oGIZcX6AHzb/ka8ThN0tYSrG8stKyDDbRR2zaMeZPIUTt+p
GUjzgosELVLwaWJMoYyhnevCuJuzeU3MHuovT3MlyeobBFdCQHDrqDyrkjurm6pe
1JoG609lU7ZHUxfPNxsmHY7dzwSycx5Z+iPvTAHAuPw5qWBNO2foZDFNLn5nC0c3
Tkm8aPjfkVhlG1WPQGzttfqnRfBxYhrGs+7cCcIFhOMeHIGHA8ePjDTZL4FZooxK
PT8XtR4D3Kj78tYAhr7cjurqZCUpRVZEmtF9jU60UE5nmiZCX3y9q14gEmd3k5SK
NQc1+6zjz3H6cNCiP5iZqrt2LdxUNbiZ+194JzFUjDi2i0yzO3ewtS5BzSQlQnYl
hXkdsC+K3BMqS1AaEK2s/vCpG9QQEX6Iu7g6qUwtEL71+rCdInAU2zrP91TyXj3p
+cd0gpui/AJbDdcoYpqz75pRxVIl5RltktNRtlxexEB7mwl5UfWve7YH59fqTPPL
Zm5OTixb994RIgotFkO0Wl2tYKSyI2u/oA9CoCfWFOoyXhOCd2ZjZHWvasARONcE
xaDw898okyzw6scXe54AqVS1OuizPLgX1gWZbxI1IRLe51TVGOPYJDgqjwtWiriM
XBQotfMsYII4dy/f4VZIayEckI6hs6Uc824TuCR5l/rQQYl/bXp4tKDWUTK0WGzq
oX6SVSeCq6UHr0G0hJq56/m2zV/Qnu4eWUwgmDQqfgyS1Kq4m5MUdfJz2fL7IxYE
e5eTnIqfcIJbl+dPGpjIInxOYfUUBVbH/GCmNGHdEfzv4FeuUUnZFuo01GeA6cWg
zV7P3mnf0dckpg8xe1FVjzI0gqbAW8pesCoAP+w6+sSWhOo+UILpTX7YL3C13w90
Tof/uz6qwjuYEOkatmPPSOIcqQSrSsC+3yoD/c0ocLzlogdEYkkyt4/CtLI+hy9b
cgmArvPcZDCTSXTIHH9No1sE9P+aCAsOWYGhr81LUDgysyR8lzCpJGEBcdAP5HI5
rn7lQF0Lcz5muB1G6wP+bgFHHT9M3Hh36khNBfabwlE21OOIVYr222BQ/C9sGg7m
8ZCg1fysQggbTi3h2PTbT3KA3FkcBPdWFbeOWHazK2j6XHiuaTOSSTlMeuO00gG5
Bk2CV+jhoiIwnj2RKWsCj+wnxCmpJu5k2eYfQUbJO2eIhnIDHzyEVGlLQPTslSfz
QBuJi5V9bP0GxMZNVnP73enSvvavNczQj4nx6vwaVXLCS+eddpCRMnUXz7jj5oeZ
VC6ehIuAIeYBoM3sfbVkKZot0RmFZSZBoc3kldHknMlMT7BbQiGL+uzuPTu8+aM2
zmN/5qelwvufktlKm1dKWLG737aA9vLHhy5J0VSv06BbXW6pwBMfjQOq01G4wOdx
Mpu/4f7RSlgwEz4exaxcPL7x/8gDGmPb31ZDSM31tTeOA2uN8QJS+qZtOokHtcQ3
hYN7wIfrm5uyMyM619oO3f8wmY0ikJwivadigz0O4IDW2t/wEiF5c2laT/RJ/6j7
8aSeY3v7s3kWVaKamJ6wn3PfcsGsBW/E1KbHFv6RV/Ndmu39o3L/KflOu7cJF8Qv
836KwACQ2A/m8f+CyPfYir5+VlzpZSEGxFCZTIWyA7QX1eB3ISZS5rcKGFMIOEuu
ih9jkvXN/Kb/6jciW01WuB91Cu5n8cW10diJ1ylnw0S/tEXe4tcfQ8eY360SkgMY
4/WtG7JNXjs9je7SaItsayXpXiM+4c3szw7Pnf2c5Zw0NLUkAoSP3QdcsslOZMtq
WMbxmHg3tdTQc0NG19lPdKh65yimf6BLKtOVkdO+V27NzSSqxCZ8ujeEKpM7o9TU
6POYzW10OdoR7k3Aj/kBnnBHw2K0QwHryCU07fFtKuI8ntF6ElN9WR1N3LiIuDEP
L0YnV8pC8PWtG85sO0YPmVhWNxTsMNBeKnGUuncIRSpIO6ayAJyG9KUWm6j8p9JK
9rgYdGTnPPYsjSFJaWthboqA9lc7J3J5R8VrA5N4+rKhZSpDlr51ACsEqRGLBjq6
jmq5gF/kBvdeSOUXiUjJVVAPWIJ981HFGHhxNqanEAKSNJAtcaWmuqJj0PcUnHmZ
431tdzEDkOdnsJ3hz8vDxDqhmJVMbKnF3p9S92HZ3O22KFBjOkI99/RPt1BCnvGt
E2Fm5PxCyq97zcCnzXuxOQ8cMsUhoG2w/LVJhWfVovCB4B2MpQPDjV0Gx87RmPzP
DGr0x/xDNyiVs6xRxN2wUCysrGMVsw+14ckI7HTKV4366YSKn8ZyNS1P8LGjHCk3
EPbCeNeHygNUyztT7XKZoYlWX1St8K4gpQ6C3u250t/wGwgtRNXvAd6tV+pdfb3f
Y8Lt3s8lD9cmmxD94d+Emfv78Ls4xsy9oGfbDA2+HpXcbzkaT4iuE8BE8R8fnyfo
ZuXnSQCFs6PnQT85VVtY2SCuF8sWd4OmrcyZDv9vVMuUtgFR5iojvNAB6X3Sa+nj
dOEE6wKTC1EJSsf731ac57zEa16llPRMvasYaXzqCjcb2TdehkLUQXj/s6uDqhg7
AqHyz3yKAgyryNSj241Jo/udzNl+Mw+/KC5ii7Yvkpw6EMx8fgTjWe5XyJNIYWKR
7oC7cJXZqS4thvB5sXzHntVdXK/ECRDWzEpVhl0A8MhVBuWSNEbfCmVUwuAL6Wgd
tIRHb2H2eIz86IqxmwgKZ/6Ej5gEAASoVbTThANkIXiNLp8m08MdK6VFJao37yvz
fBTpUNPjIjMBun/3YB3A0JojIgEQDJKYG4f79rDS/fZ/V1BYRIpYXp+0+YzSeCfL
yTaDMsP1KjJuGefulAz+ITEam1GyRt2DTH84vFgNB1LnQxwiQRq614GJAMPrEin5
J3xBPxe3qr/NVI7kvboLBTDwBmpjZggnSN90La2U77k1ToqTU+0AwyrRNtRsFdmQ
GA0A2nuVec0uZIUd6RoZOIihMAT9Eglr1WLVpEfyEO8+BddV0e1wscIeMwdGR9Jy
xeVNssSoboaK/6cjDihcQKBtAuo5UQR9AhMH1owDGZWRcMSDbNYbdv26qPp2ypM5
D/ie6ZZHEagMvPCXD0U9Qvxq+bs3zcyy7Qs0o+xQabzG1KrcOsMOwY+MsGEsJQUi
Svnsx4/TaNnfoatnI79j3Z01R6nG3P1FhIzLS4SB3GX8oPmyiElgyUeuhwv3MXv5
+q2HliZbA7ue9Pa2VwOQbJMk+lEtfV1ATLZtLdNNRdJ8sIm3x3JW2eeu5QC9lImj
ZRmfUHyR+HWKcUB1FSJuNDEUbWJ8h2BD10nCDIR/NvpTFXTCGY8r1dNZKOPZ60C1
kW9NgwLqIuzNxXTiqRc+17Exrb9CA1HY+AlD1TMri3HhZ6zPL16HLpfHI/JImebj
yqLFKLBvY8XBO4oAUOI8dDC8gFj6Z5K5hNW/q3iFLeLuzifie30c/nH/NmbYC8lF
Cj8OsqVEYibMcKL6OkxS0VcjZBuxh/4uPXn+q/tj8ROP8/4dMJd/m9UiucNrVhLo
6Bz0ENOZFs59qeHdPMg+WlqjeXHLcA1J4zohieKY/TslbsgwS2M6kmKWOq142Nh9
Cif879VCjebK8H6Z+oJ/RnnZ15ZCAL7N/JlLWvOlKPLK9WnwmR6yf6rJxpSYR5up
cMbmV245QEI3bTf3Wb6NdQrHFnfEHnmYbU/o8eLqOyv4SPUaWRigoQH6o0AqXnBU
XIq9+QxS41FFy/vngivIc3nlAtCeg/2DW/A/hp7FMsLR0W3N/NPE5X7Z+zMKbZYI
+JTwZw7KQnrdPbxC0HM+477KvnSMeAPxQZgKj/d3xW+xhHWF38g5MLj62sUy/ary
HsGk/l5AEV9/X6/45n/3l6g6FyKm/O2m8i3WRELs+5OcjIQjiSMHKdCfM/N2wqid
2CKsJmTQCu/9F8GHl/ZRYdDDgMqUeVXKRgvr/ZZnZhf41L4LmRpkY5j2Un/nMEEp
SYIQhYNYL3UR7odpmC6ZZyG5Tt+3MdJAGT6r1Y5s6m/pZrSeVuATaGs3LBttVu9D
RpOxV4W+LsdSlk5Pj/cz8hhsaQi0+IDN/9K7XS56itkrJc/wkmXVGLuihcYY/vD1
2ml8x9vlQ2imNdRRcw8BPvUVMznVoNpP5xUYf3ViZpYAGque0reh03uCVoKj6sKP
bBz7dQNIf2fx0u2GN/fo8GjsP3Gresuc07KauMvdA+pGw8teYbSQsJJRRGAKRaO4
U9zwPshw1mlVR3bo7p57lIwPfRwVFj3nGjK81MVfgjvGL9Hbet8m7XXwfAbY7mLE
NdcUxGlHBQqBVFctEujiWnbwuH0Fid+O6lMvg+n1ePCVRcYRqtRJcLy8xcV4bLWL
qC1u8exn1ouhyQNd41jtCBEO1OOpxvL8msE7vQ+HhBQ4utc4psngt6v/puhRGH8g
Vn3F6WMXIDCov6My/MClIrfZ1XrzmjYGkyGCxcSsFXTM6L+zzKQyltxebLDRS28i
BUbDsH1/wgARKd27UQQDWSz7z2hWeIedx6SiNvGu9y6dXcrvyVFZiPeBYOQAbnqY
TEawZU0csS8Z1a+F4MicvJsFXN3isKR7Z98nE1yxAMQnmIN9RSSij4llKDxrn5iI
khDFuBBhdm9IpP2T2m5waS01x3YL8kbiM5dz+B7GHkQsS+j/MmJqqh4xIjttmWB+
oItSKD5fiu52dZE/Rhx9P/LzbW9vjgv2qnSpZGXjLOZhrPxHwAIrSa5Ee/as6jkn
26PQmiILXvxNAdAHO9N75A+o/nDMdY3hCAKz/CeKCCcAeUzmlsydrabQ7P9meZzf
LCvoLNdOJB5zjurt26BVlO/ZJK3ZVRPUU5Gzjs8H8FML51/sfpb/jzWOvS2XVCP/
NgFRUvxy2U9eLO9u0plUanOfQamLR9DgwZB+BxkE4LaWJyCZOwwEmS3Pj2L+LdTa
OjCgkda9XdHeRH1+25E1sxSab18WmV23MChbPr2JcoJ/WiESZyQp2r6Yn3I8Bgk3
603asxsrfS1CGCLTimaJS4d7VlEnAMH/7HdPk5pdxQSqGm7xDTPouux8zyqRN9T1
xDeDCmk9Zby+j8OgQb0RelJ7BM8Aqp2PPX1bIxg5pL4PeCogQ1eWpaVygF5hDFxy
CgJNtQxfAPgK+7/N2mfwM3QeZB1Eskhrjv7Os8Ur3/hjuSlUN9nVYuLTb0gsMyu/
c6THbJneeLXGvxHkbH0RkR3xJlRb5bv7n6oUA8AqNf1N7GWC4T3EgMT7rvmo0ZTg
+XhMFnWm07gSjUCASlwo+6KHAnu3pPKKydcd8bOuNdqNjqWsdx/9UzdrEb2R6m25
7c5dlbe/GBZFY/i5Dp1thtDI1Frj61DfJx3lsqeoiLei8+KVl9vCyTOuvSefKkYf
4EX2gG2DDqTM42MjX+cAfIOC7sfKtwIHsFImhjIegHJcRpy9Us6lqFFEEy0NPx79
//x9tG/1unbFPOhdetJgvAZt0dYSxQF1e/qAISQDU73xaozlnU0Ly6QxeA1Rk8J4
imI1lJPv3iqt1XwyejZrwNBiUObZ5ckE+FIBpEDdELrxDcGvgCTLY7waB/dQhC1T
tl3PgQbSB1irAihy9jR78bUQamTAzUXLLMQKfgT8oYhIA5UuoB4su+XtvJDLUE0n
ubh3qb3dKl9VwMv51LHJMpBeAgHx0ZCikIIdb4C51J/PLGF6SywrHCKC1sLNvuA1
STN2ZMZH96DJ/2b4aNh0ZHK6DJxF8+4KnSusP5Xcll3iOD98IbqE+b5H0SfzYlxA
x/n8aXw8Q8u11Fgzgh58nXKASlWO18C8k+CC0mpOtghZHg0NAE1619eb5FFElWK5
aq9ZQodzsuO4b/hA2z0wmKPKQzox/RCmdmX0BO1y3sXq6QUbh2wh8iAarj1mA+12
xRgAIvyj5qXuXPnAg2Hu0L0LEZnm7NXdXhhKvvstHeWyIH4rXePkUZBnMfH5I2Pi
RAzmhlh1FTr65wxdyYcUX59h2xMnYgfQkgqWsUdBZhE9cvw0Awcv33+ZH+IaXuWw
u0m2+tedu9pN0ag5PijaXURVjeZzCIhI72VQaIIVYRP04ABTVacnKQ1uNGO/PRCZ
g4s0vf+P29zVuQNoK0seVCnjS5ww5Q5DtWvLMMCq/NgvBXBjRhMwugp7oV7z1L+g
5eKX5Y9VY18/laoLiEdoEyDZy0V4MmQwDyc7W+90QlhnhVrYc48Ni/clh1zEaOSR
xxUvkDemUDV37ZPthuY1Gp+oT4I6YfeTNvtQ+/KUTgeNaxdJ56xXixbgNGqzK0qU
bUO/uJp+NHlrfj4IfW1VuOjVcdq8mwlo6Naz4jDAAnhq3oEhDkYz1PFowVXj/1NJ
D2hVlfyHbBt32p0P78q+hYASwaZw+lr5y7K9UITtexiM/APbSbC2WxoK6x4XWVMP
K0uDiia9DnPtvKeZKyZYjhxljQiEPoIfaeyABItgHHS3ex5FVmuXOn36IM8CNnr5
HK1MwG6DAyAM1qTmOzYRbTZSVuq+kGgmdgN2zW1hP0Ms/fRg0eUcHFDxIuwfut6B
0eJrn0yRWRtuJIyTEjz+On2nLLe1FCOM83iQKzLlhFnSdC+hMUy4pgx68f3hwtar
0PEBBi2eJZ3IARI79Ji2+WrkX99zyC+OM1wqAj2KDv9IosjRDX9w2YABwcCHevFs
Uz8oSo+BNt+7GGJ9qzH/yA3XtGEgVWKk05SDsT317vBiNqULJI4/uw5ADoITbEth
ZenWa5OPZWumxeUvvgZrkDJQoOs/bLjRNpAxm5j6RKoij7CcW7vV/FYA6Yc3aFIW
yh131YCQOsXa92KsO9n2sH5pKLyV9BeoiS14yKI4o8i9tDwArE8W1wZ8FhFtN0T8
N78E+BoBMp6mPTGNlNSXe1Ao+fb5GwbgYO2OkRRi0VKSVAT0p9nwIJrYIPl3PSY+
Hz8uFDKauZDpr+X/6ADz+pVLvtW2Vxo/wXO1CxLp6+8JbkfswVFRTD12aVZJ6u99
l2fp00lCKgdxSy8cpMFPlFgjKDooJ04pu8PNTOwBllAHRuq0s3ws3/WmKTc6va5y
N0TiH2Ekmlu9YQvCUexRSSZ6eoMIC56cLZnyAoWqOzeGphOPo+t3lgG+nTuNLKxE
DMiBIx+fqHGom8AocDNjVLY2cwzB4YLajtvfFJnosMcnGtz71X4Bp1nh1Bv1El0c
Z/aqY08SKCjsLt7R6Noc0N3MXMszfknFw+ebDCYnTBeum3/35oAJ7dcekfe6lrci
wCvlQd5Xwf6Cd+QIfAmxDq7MFE1To9+oyvejEgrmljdq0/Fm3RB3mPP1qVW7O6C9
L7y6yDEeCZp88QKs31/prMrdvq3dzkYK/e9MbcqIhfMctlWsoQ5Uk5DmYKFCxtwB
RiSjJ6alzOlvGsudnTQbCvVKOwGV8NUFr1fWKqN7xifsUeKBHwH15f+7L96SnQ7p
RI0B83QZ3YCtDgAcNjljA3Z7QHkQXAlLNw5aKYL/GiYRJxB0HIVtKjIbj5WmqdSN
c7mc2bXpoyv5aG9JmnIc2UWM4QtYrc6LV6zTjurTeXNG3vD5u7DFqMAh/B7pTlbK
Zq/yZ/UM78/H5BbnonZ6IFLYbR27qUP09tyGwJgOWJ5Hju1nFnzi3fnaYiP+ey78
dRsNgsiMnBROnlB9FNunXL7VqbNV2CjE7ilp75cIRfgNb5m0Die0/C0TQ9QLeXQW
XQl9icxASEbdtYPL07W6972QZ4DVTAsOs+q4T0g0O9eCsBiOgf5HUGznr9UGWFeX
z9tdBrstS3EoQQQ8zrY1k3+qXkH6vdw67DI/WZKgp3qCCKc7pGWLM/C9NjNEpaNV
jSnugHGSkdZv13usItwN64slgxYSYOAxkFK8odtfscqRi2is2jONh1xx/eIxbmx6
vADj4VqwJgeXekQCL5Tw60YQogSDmYHm2KHX4VVKcd4EqcWVXHhieu4N+nRntndj
2yuNS9vHGYGY8coTmBFzA+h4Tw/QCKamRVnpQiq1cgDt204myKQxNO2LBcuS6+S5
kP7MnaTkWvR+Y8tn3DfX8UVTHxaXVCqtnM6faxYay+VhlLqLYhoTZ6fofQLeuEXX
WSzIo0L/cFPsSp5uKiMvCOz8PdtTvW8LUI7kxNarYipALrGEDENR5i1D/2VgRqhU
W2yDCx2Ks3fvSr660MU03VdNVgZFo/NrtBRGzq4SXLabFEgzZikj64iKjfvOV/C+
Sshqml+vjKMDm4XbXcUDkyhTbKuPKH9/ySSczN2zh3efcwIwCwWcZOZEMYMmz67C
Q0mb7aB4uizEPoy2npFZFHbCiaheIs8+0sd/I2XkfuQWC/rDTv2pEu4C4ghNiV+D
mBJp/6KWpb0WelivLWDw/ZX02FZYFkidGnzn3jH3I/kireWq8//t/qETWb5HRavV
ISTuTZYj5nrdXqAaJGbxRtpVLwgDvt8amZeDIQxZ4pL5pOcjJTSUVQqAsW0UWoKG
IYpZ6w491/H7NVZ7CqLGL8b1eg37vL30t5PSeprxngFra3n5fq/TYsp4E7LkLT7N
FFr2wYuKk5ndZav40X1ZMjmBSU7gXz+nd77fwN6BrjPPDA2FvRbheE7m/vCv/39X
aSRXuAxfTJH88dzeRx/X4FPRopqF/343jeF4PH2NtkttMCfv5WqhrfQsWaKfpM9V
GwvYG29JsNxjIu3FF2nMqW89ODxqimJqNyzPsdGDyAxi2C9Icu5qSV0JCJGPdW9e
/nORODAsuVX4WiXk+VI7mYbGfA9OzU+Hyeue1N8z3WbtR4kGYhpjKixQRZ3wX2ID
JuFniSBxydcdE7Md1MHjmsWbjYCj+4GW03tuWvlur5rusFkN8edkCAs465mUMDC2
NcG63uVk304QHfqZiYSPafjtHUAUndeeX4NSEKpbPbPhFf1P9/TkRxGVtMyXlQGv
o4+g16eWxBfoSlf+s1AJAVUYxcEmYu1wUdRUytLUtzT0A8nbWOlDnPyqFPwPYpba
uAuJqamMP0mg4KsevxWoB0ShQKs7LbG2bw1JwRueAhM0Q8LbKhawWtoHFveqc8yt
7NU3YNAAN94Ub/Xqq1vB/zHfMFl1tsl7AVWhHRBq7GSqxQlSKJHqxiPEewetadVW
gLvCun42nXaGxAd7f0FlZKx9gYzx3mbY70ryjSnLlZzjpo4QpE95aoC7iClKzNiy
H9MQXOTGGX8+zML9sURCm5ft6apVf9BKr5Bz6NW0tkyMLm0ELQsUOyVV1N88RqwF
f6nL8sYHzfDSJcdaCCZ+79d/pQ+I5SLQftKwq+DfF7x7Hu1j8ohcsqbsRAqdQjSk
thwHHRRM5KP/FhS8bqFkEWxrXOWx/cdbvV47KGEpsQkeZ00WLB1AdHBw01H2BMmQ
SVbIy/hPIDuj1xiawSMd2hnmZf/I3TgF5xbou+W3uwCEYxN4PMhbHy/F5CYJUnm5
DyEPX11P422dBRG25rhvK6+gwRPWp3ZRCPr9IV58bVI2PqTuM36fc0bxp1LfWw0q
6cJ1PuXQAEi0q+BGkoCXSsejz1pM3L57OqT+L5PCvsEzhLGRag7DQKoN/HUOJUHo
MGUSKr7EkKzKFFk++BEDIX7PovXrEJ+z7yxcUdkMm0Zwf+8Mq8/0DsIPEQ7M+noZ
6tfaqlQ4Q1FJA0vA8FVXUt+Kvt7s2+H78U+Yrm2L1+Tnjx2WUq8IeGRwF/NwcuM1
b4A7LPEFj/t4YFaXphlR6r8PXy8QtAvfZI9moohmYi/V2ghdqrB6qA8un4y1EOvB
i1EXaKvsi/jtaoXZsee3mPomajAXg6lx63wmp9Mj06XKu/FFkpuUjklEI5idN5vH
J7iiOHiPO+U3VeLv/l621bRFiosu3aeZSCfVMxWGiLQCoJMf5XSPxrIJu8FMeKKP
7yN+Rih8lj4k7uM7/AT4mBXhbKk/x5sqb5S7TJXYbVwA4Lp7RvWc9icn5N5kYH7d
XGTzg8V+tEAixRFvGG4xsle3bGpzLCGV97QPaNafUbWluShMFgSisQTR6ZkI3Sc2
jbp0aofmMHxRkGEBckGT/33+n9GAjGIeGNtJLpA9rnvw5m5yLdGGyamYx+/0XqFy
GLVXaCmXZwTP3CkzA4OKhQunQhMcPuOn9CTl7B57cMbUv59gRJ+yLihlBiHOJIaS
/oZudptHIHU/cvWQbuJ/Q8a5jCVXzqDN8Ku7eyOG6EO2W1zUJsk2A+dKsGV8L4I8
lj/sMuUcdkC0HKs35Fs8Ylt9PwC8k0/VZEHizFOb80HlDs9hjgLyRWxg0D0ue6ia
d9ee7M96qyPT8CVI2ek2MeHwacMnSZtDXfMsqjYWTo+I+LfZqPApfNHitTa2l5UR
tmCqHorhygyLRIRKAHMLB70SCkXiz50V7WRetWvNq5K79fdwG7/ImSjArlQG8k7y
rIoC0Odb1ecNjC6saiGX5QZG3V7pA4Hqv7B9DNRyEF0IxGXt0H6ssB7PZgAuwipB
6B108cvbbGwe+sswK3AJUnFBZaCSDhuTpzNgluZY5yG1GswDyoM/gg9dfIaBPq15
aB7Ieh9nCf5UozLQWmFA2FuiVuCt2NtxNLJcAMBJe49PEn1FWlE1DuU8VCjBGjSi
2V9EY9P1nuRai5+iirY7sBZqENXlJvrSSUtIxy4WaZsmbUpdBtyFF+t4qwtVZyvB
qgseQFE2ONZG2O1eBrFHlLWzg99D4xfkOge0heVddHz1EuElUAH93GQKtvoZXDvm
4UvWpUQrPSketvJzheJ23g9pcxjUttUXI+sxXKkLuSEe4xtrClRsYuURXHpBWZ+v
ZT4L/b2gg7IYYloiz8JBZDW1Erh+hX4YX3t/myr0EAGJW2jx0BpiV2tSbq4zRN5p
Zyvk/vddfTAolmgz0UYvoyc9LcaJ6mEJmqSuozfI5kjlBP++B0FLA2+FLU5uE04Z
qRkPxprvR7rpTigUnBYq2vwFb4bVvHAeyCO7oxhdOJS9XmfjhszwIGHJtcaoeeTO
EeKtegCNHpQVgw9pNMQU34vG2rVJCrI/8hwJq82rXFhASOgMotTIObp23mdTLm9E
4OCN//6H/fVjIU1wuo8LEgJrTj31bMYDDWvtLA3noby1zdQkjE/5PHAe0ZD0JR9y
uhQfZbvsaSl9jERLDR0cNT4kVAaPXETyqKhsZPudGFzUpZwkkuIikFS2XXYUtAuG
1C1c0OlbvdKOI5lTvIW6wTeBMtNCk6S2Q5JdL35Klo4SKi2LKVFK2WbARRtqy+Cf
npopLPS75bOB/1fyg5+2smRxWgWv5lmINT6IKZS9JahKH3+ONHBcAxN+aBdOlw3C
DozFwMQ9lSRdZcoLpL4ZjeeRl45jNY8zq+7BDx+BtbiOMBDjZr594jSZHhBpn3d3
ls9SWXNexFVIe2qL60KHJF7BAeMMY0mhCW3ZyaBSGb8USTQiDHHyPuotULgavnU0
cAiOTJtcd9HbI58pG1i+aHpvX/tX8gzCMtwIUPR+aKl1cAwg8ncUlTN3KLxJ9DoQ
P/9+k5WIF6WfDLw5AZwqFUa4TSMrIJcH3cwTadUlyzn/oRvP15uB5lT7m8Coxmhw
UW2Bwr92tmf+frpPzj6jUgFkhHF8Lt1MJC/EomXf8QcWZlgzDjUd0yRi7WCfWNTg
9VkaAMi+l+UaFBFI2p7DW5/DG8PY5Ibq3mk/AkYKbD08Dq4kUF82a1v3VDFMYxnd
mOK7UuXXVTPWJBgS/tb12AKTXOFJQ6p5kVClfV2QFptk7Gi2IOfB5X5lXGDaQmXJ
dT0cK1GsOSWVCp9oYFwWBRguseJcK+rwxv9NmSBbqQCrV69t7hZluAl6ef34dpx7
bESMm7Jljv3PBe43mmy5O0gul5CpjfRivVfWoVx4TC3FyerKt3nZdFBgkCp+MWq5
jHl0BR85VeWOE9sTX72dd5YJFAGVWRTzhCv33yMl4qLHoJVl94QcEnz+8V2d3XC8
ZoRC5nLowhAxGiTDE3tzud3UH6HfDRcqFoHIknLdKJV5HX0oUN0A5RWHYUg7jUd0
3axO8120ec+B5sPn6hMlcdWmhBootzLOfr+0Y4LCSExZIp+zz4VRg8u/AmQ5mUN4
ABqO8zJwpBdxJ4DYT4dqlyO57wrL/AsaYERERbt0ltUAJGjq5Yh6zyFh3A/teneA
khTB6upiXFayGTGi7Dr9UoArUNWSem3Zh8VSZVbAyV54E8gqpsbls8hM4O82Rdlt
VLpn0/s2kPOqx1OZquhcHiIOPg+xw9kccbWOgFHSG7AUd9NY51HqeMJBV6KBfEcX
jckxe7BlOjCwyR7+RuuFv7LeMb3+Epv85weieUXivFHCk6KJJbOZ4UPcc/gM2wAq
JjNayiphhV2dJA3jkaQIk2GbzKJ33s7rNuMDzsqeLXaPuhqR3YzZU6Ptr7CKlS1B
WgkjnhTwUl2/z5pEaR0zYinJ/O6aiuMeV//cXbs8NbU+Daepi2WD7kP2gcCWWqKD
qZhp+/1X+shz3g/BhmsC1HWCBps33x+EYSWoVzvKq15i71GaiHeQwOCF1jrSo2p6
zSO28po9y9yUl+b0wGIfpMnSz9L4FZ8JpbF3pHHNAah6ljhOA882qfQu5OxEAFNX
/MhLF+ntUmBowPqeOuksKZ3CsSB0+bUh9PkvgvwyFsdqfW+s7/OvYlopvTvViMvt
2otcw+/lgG5V34WUTmV6zIURkanVK5Y/+xLc33CN2t9qfQEum+yNt68nkYCtflaT
xX8CsqMatU3sQL9FN2r7oG4E4BtkjI1AunGoZMi6kPcRZ9HiCp2/3OOyFrWYzvOv
swfqSSLWjRDLrR+ZiMQYbN/3DcM/4UDUcI8BfZOlbHK//7GfGuTtfDff/xfF8X3E
EXNYmldYpzoEL/lkTJP3x61M+Qb2JStaQ3sj/syaHwxmxGVXfT2YHQ6CRN2cZBSO
TwYbQ6gAVNQTMvXOzO4VjpbMjh3zhG+1ufJHcgbyPPKbF3VpFRosMfTVUOQl64jA
8DY2io9g1tiuV1ihZEp3Z1OgU9Uc1LEV92eoOgYsGjZXmFtn9w7pf5SNTBrl7ctU
BR4aFhIalQT0uQj+NpKhAbQYYr/vjKt7FnTgAtOLY16ljoCVVv1+n+L9Q/gtoIYx
MIoft0Rkm4hh5lp23HcFO1ucNIg0WZnHUqThJfN6gw/fxMvVoF8aW12zC83Jlb3Y
TH02x68QJV8snA1Yx+ofhGG0qNaAYqxank7rVcD7ELxVLRvyhXCG5zJJKlsZDzdE
mGt/Ky0/UQgPId5MDmcB/8c+3p5VJc3bRnZLbsM/Mz7lNc0PUsUjQgaYWABn/vGs
dDWlztm8Tit2gcM353WElkYi+PbRgJdUkPuL6Ul8xNDZm8OUVLHntkSueRx18dNe
lMaCkHuWooHkG1qJEsBMve/pSOJtaXo0IMS5znAqU4bGFSPIr5O3XC2g2LF9cQJx
ffRxXsyxdYrIB0H2uMpt/GRSvTMvf4Xy0yEphId+WNbKn/LgCHSbx0AEbbjO/Ng6
Y1ijEERLg3CAcuAseYOIUDrJo8+uKBP3grNwS1tu34JfDkl9iRqnx8pl5DbHVugF
EbvY4TiVxx0kTOxl8SKvcsUhhrWFb+td6EpTXPTs1WeesIot3wd4QOEjaS9CDNLp
czalsV8cJlMHdbX4Wj1OWTC7N32tlUhErEY3t2KYSD//LREfaqroJz2fEC3q+EY8
pWGc8kOS6T0WZTShybKPgjZbScrPYe8i8oRbAtOdEG9LqXgMNpLWxdNxfDth5SLB
awUFU8gZ9kxw7ZdKGzeUcHORDLqgk/FimnKO0HEU4ISpCebiwcLTvR0fJ4IOkzYF
oxazscIwlpvl8l7KEU3X3fm7jgl2rXWw6JlFv68jL+3tgawbPJV06lw7oDsrPPCw
zr6AY9DKNzzuVFxaIFfNv+Whr0Xz1R4YLSC+aL/xsyc9s0OsIC38sx977WC9rydX
4eLwVhpCvXT2+huV4DCdUejD+OD8BaHELdqEc82yvLfLOPc6Yf/+xVrQEx43mCWa
Bg+EciKCZPsiDuc9ent6Ji4SFau8W26WxW2Ven+ujzsKzjK1/6kATS+L5JudxLFX
5YEt46b9usxuToQfsogLzIR4L81AXLdI2KIXSAdGGA2CLEJmNBVqy3tsYPH07zMz
GEIBnqV7uk5PryPpEXVXcvAjkgHLUEqgIv+0tnXcKQnLxA3XJuXdFCrLiIIR4U2V
tj/dcSZY6lnqZxxWEJJkhp/UgTTL0MdwIfGTbCfZ14aM8srUjXL8kemUUT2FSgs3
cwgpD2VPuD3TsJaoOjzl0SfXrlzb3gkWZqPlPmH3i65gjo+0a1YMYryYDu8QtrCG
EEut9hDrRdEDHi8Lsw/IzJthm3uVICu4XrJANqcBjHh/1TR0yt9TxtrKvQemnk3/
SGraJMZ6sRS7T+C15vJ+9DwDt3NfjR7rmnu0ZUVsySqPd2Y2JSzwUy+ka3tSdqn9
ggv1itvom+C0oHpmIjzufGYgZDzgq4T1Gxs8MnZEuvtNbWpIgXyekIqyg4gbIQHB
Si5hlPYasJeEMKOzwTNUvIKIyNTSIMqsG6COqOZUxS/vYkCeVDowSNPg8iuM9XKp
qWReIpkQToxPt2jt/jE21ScJOit4Qzmiij4wYsmBVLG4bQkJLouGxthXfbBj3FcU
lJTp7qYUSYiDXrNSlNvdWEGHCFsBxHWNcRJTZhl7U4OCiu4p73u9ktd/4VYEf+Nt
pxcgUi5OHuoiTUL5+qSUJE7c0VDrHuxSsMhqgcBR1jbdHS79TfS/rNrLXW68SABL
OAI7AT7cW2nhBqX1Qq9LcFwN9xJ/punV7T7Ya3pwjehGLhum8RgeUvcdhItSVyug
7VAOQ+zzLbgTj5bB995xthVwIkMy4Sy7h7ktlFVH6pYU6JM5KItEPX7Kx0s7GRMZ
OsU1dbJ2VcvPWZAc2S4YPqxdXuIxPP6u7V79gcRaXr84EPy/4ggU9xX42aN3HqiA
kEaMPulZWLFTibTU1eaS37Q7n6Mtesswhxi6IhbhjlQEwnA9gjKnuL7SaBPzN3w5
+iOHQxiPgdAr0IDvQt/Jif8xwVXcrJlatC9rLWXvTtPUnWiluz3Pf2dYcHeENMJL
n2YS+RRCXkzcCcDImqBxcaRrdjwk8MdR3R16ddgLhSAU/KWWRTrVPh2Aq6R82Y10
5xU11/SWo7VqWa1jnap2EI0yJWoHMLU0rNf2GgvU+IKFZdFuuUoyLDkO7n9GB7oh
xuKGUjYYYEhUOpjcCKMIanUV+Tk8ZotmO7XF/mX2RU70QMN7Ttl6Sb59u8gom1ul
/XU3Qlh7dko+vDWE+xQnjyE01Icn9O2ZPIAeKr6egPh2JZBbv81L+VayUjedXT1N
SK0fCkEXkvpNzGehY8qHny8KZ97FyQq/baxJ61KTL8qasiQfM9wQpdrkMhl8N8ab
3nDUUP1kT3zdKM7xL9+BEOT4S8L0UTTYTPdjfTriOXRvbg75TYV7c7j0we3XSJwa
rO+K7N6rtsVAHlJIPf6XMnrrGTDQJ2V65cQ2dPZ84yH/DGXvAXYWpueq0JckA3pW
TRRNgw3TCgLrrpCDtZls3+hbaxCUzxN67qZ4M7RON9y+k5j/2WGIvvbEM9wvyUkD
Y6tL9e6cWBdtMfzrHeNkcSZsjfxfkehCukiAEIF1p7JE10FQGf4qZ3TpY59csVA7
3mMs5zp6IUwZ+Z7O67BuNcR4I0NSoLLY+pK2u8oGmVduVmwuxz6ej4LESQe71HO3
2DLROt0+/cOoBr2jHgYpg0dnDkaPcqrEeVtFdC3E+gQTDZS0gmm8wCtbeyWF9f4o
FT+zLWM0Drx9/qToyKxTJJWEpWH4c5PKiX5RYT2UsVBWUMcQAXfV3/jYalfNG3Er
faOyMKdXp1dTUg9WY87CdbEx93rFhvHxdNc/nzDGJb/gZK6/lZjjr/+1dcAr7Mvl
sWyE7GMfmHEr2fbm2wyjQaqIJXMMsHmCcJYtO20gI0yV+d0esSJjYpcA2FVdfLlN
GFt6knJ4s/EGXcsm1Sml1VIObMslGj5G2rV2BtvPqKS9lyKWCO6HnGR0bgVDgwDh
WpzkKyx2Gg51/AcBLxQTzcb7uboosQoXSpVDxj/RrkJJTdQCSXh/IvngK+j/k9OR
DbdL4OI/9skyTqJDZN+qh1Vl68uCAigYM+bViB2RFUVYraz8MJ9wvwRJiehf3TtM
mMAWGuYDTmDgnUJiWtC3UyE2N7sw9T7X78T27Sbzi25ASL7Jbg0iJwuiEHWUknGy
877RxFLgbZQSMUN/r8GRbr/oFCjrextkVML7WDywuS9zjco6Go8chkVEdLtfO5zL
0SgnUlu40er7WjSV9WMOSFgzz+mY692hhgR16LmkZsCcltIKlvpByXah5hMZSsh3
gN2C73H68+Y/9tyxZf57JnGh5QWB+bpv6mn5/oB9FYpW5QorzsbbJR52MC8+gUTb
hPirLCvu8YZeRMdFH6uMatZQuFvKYNYSSoXLKWi/h+eKO3gorVD/UI8xVzf6yW3K
AZN7O6IvQiIxWtMSRuStgJjOR55hHBXHV5KnN/bUcWV75KvH+tM+f5Z7VcnOwdlk
G5xpWuYa5ry29EpHIx9KGg1Tka4YyjjXwd84zNz0D782M+luR/Nw0wuzf0QFUbFd
Ac3rWQpTNb0q8hyGtujO6EYewtImYNbnqiCRJLcG2D+EwuLL1fK3V7Ao8K9fGvGK
lR0K9ygljbniMQH0KGpdkeYD95KWVzMo+WBQqUt9FuOSB58IteB8bN4qnGwYQAuo
9x8jqkoxw1XpjWizoZ78vMaaFeB4kFjth+n5qZ2DDKJWJc/goGrbJfxKiTH7xp9T
t2ZGww0p9KUIU01iLWo2RjplnogzCbq8OkWgYRzOLvoG8kwMeT3iJU62sLvoaajr
ozwvWjFVVPDqbn70CcbrsexQOA5xhc1SfVak/AYB3BLH5tFdHNx74zE8zUbrEUVu
G/Iq6CceYAlKAx2NkwH+c6F+Fvnar8/Rng/BekR/AjXN8PEjBQ6IZp87Mmq1U3wW
r5+XD0mNxG3KBnOSHvcgcNzRHMo0GNZJWurytKJqvWvsjKgq9flDlfZvt/k4BBjx
CvPSSAhpuwf+ca/gGPLufkdj1L+oT7Bg6GgzeMVe7vAUo0N4YDwQkUv0dwxR5w3i
OLCWP//XpJRkWk1vGQLl61+nCwONdROeJ+PsaMjLj9nwvwqJn59O47GZcFf1kC4W
5smJAamw8xWD9K4GXmjFgpzUOqFRlrGMUoWtJC2aniPkDNLYJAd488YAywE/QmCA
wdvVYtnWnPiaEvDC/HJNsoiLQF0CDgxW8K8gDFgTHWaKWOvcx6d2miGcCRtvcSmw
9b1A0+3uVAypK5OTiMwXMJchKd8rZYmZqkvR0fVZAQ0XcweA/+5OnX4LQ+A7z1ek
u9widGvVjMalYXW6Ri0SqDvK82PZz/2qy/RoS2lXJJPAd19eWyumCNVBlTwJYnjz
GpdAx3oJdfWxbzJ2ODcU5335iuIarylQT4ZfsdqKHN9y2/ZXvPlybsu+IFabNctT
HljidnUCpyeae6b395qBmQ8y6K1Ex5Gdpk8E4joiNq5Hak1dsTiyrFUv3okH2+J3
Rw5mMc50HCLTwpLFhvL0jUIxWd57SBl7CTQGA7ExBaPP2ljfIMmKj+nAy7xTK2Bp
rVYDGOMfrPahaHqXuqEYBhnCnwArHZRWw5mSCDgVKpX2Wd4rSm3aNRfueMxISUG/
nyrsUQk7qH6klHFBhjjOQXbFTS+21GySQc57ZTem7Y0XcZiGknQKJA/zgOGZK19C
hsd2kj2h9S9Vu60IYdbFEeWgCBhZ6RPMdX2RcOpyVuD8hzX2hEpCGA7yj+7peQ5c
RWr4r31wFNvGRtlXgBWin2txTJG8qgSYyuuUh2AUWcPfqEPoSnX6kWSrA/su7VjF
Ajs8liLodDbVuPZBh1L9cKuZOicFXpAy2eUliGe5l3qdpFQ+dNGOjWyZ+a5Cy02G
qTH46NqWSuohCYENCMunFBar05naXVb3wUBUXVKpKtCYigxCsInYEV06rnhr8JW+
pYm9xZ5eUKewUuyqlomPr8sh36q/gPcvDj9KA8rDdYImb33s1dWa0Dv2ED0B5LF9
Ng/0otZD8Ut1ZFVFheuMRSBUms8E0J2Q4JXP07k4Kk/rCPvjxWumTz/RunWDsj5P
Q8e7VsHTY+iZ1AjNyIHJqvae3s+J3NqevmwcYUtNdtQ8SuDQyJ48TtisuHr072GW
r7ESHcUuDLl4l5rgpEuPYaow0uHnJb5CL5f5yDmMKXuXIEJ7YguD7uKLxdip27sq
A3xxF8PIbVw7trunNDAQGccV/WKtK1WC1T74sDhryqOAth7hyKz8I4YKLRIugtcU
XuyKWxA7oZxT0ltBiHMXeDDHzvaoGMS/pTqhi2DNV3+SzKwqvX1+eXyBe5E87fi0
0ImZPqcxb+XAjwZidLXr0oMDDKejou0YEGaWQ+II+rOpk0+XpW4cx3dTpvbDZZRX
rmoymXe7OkowB1vomjPbPmBGhgHtgUzRUL8mx9HoCFUYFIUGWamZTP8X22BE/qJW
ENClnBS2A00jY6n+4M5Joe/zAjzm4tss6w4if7VxV3MaGIp42SVkw56p8od28ha/
aKyrtDKsf33hhVcjCYAyQSRUEfgZ1jWD7P4MQa1SoM1lo63rjKedSKkqDSFgBiIy
cMcRIn/LUS8CJjbKT5uO5LjAtbLHDPwxGGwf2gEatV4LKhKDxheBpYEVAs0G8fzh
gFCAEmu+7ZCVmY7lz9uzZvJ7ONsCSJGXSnFDXThr3QSbQRNfnDRcJLwYtTQ4WCTc
/OKicBxRYIFQwCi8F7Q32A3KiTYhBJah/TQIuD8evGsxKQH2SPjts469lfI/FYk8
L69B4B1ecJMuXaLdtgmltkN3NKBNHBRgmIPyVQSCLJH2c7PaBc7l3X86WO2OIh9j
E4xZIQFDpf7X1UNdbSf2qvu0zRfCqL+sWz+C6UIY/xIR5a869eQGokH3szFJxO+o
ok1JytRYbBOazH5g7ZrAAdHQamIkT7k2A9ons0juUE2Pb+zbD0v8k7tX7mTJB/7h
JPNBf1MWeTtFum1L4HT9ZGtWvgD6b2XYHS0/v5XfyOPVEPGR34vb9uPfOVsNC4BP
imAG4HcyxGjko3dL0zzNo2EF1y2HDXlca5aOAgBGIp0JlDPa6oSsF4RF4ZXaYFHw
Nm9inEtiGNHL8Tj0imquXE6/tKIrAllQJRHfrUfCAhaPJrrh1i2YaDy8eC1HdEq4
5kZsvW9/rQTtXlePSeDl1g7u5k5QT4e1ZCeMZ2lYUFLm9WbcuJYGGssHWzDiEjlI
RHw7Qr6u9j1A9fkL9ozAEAgouygCbMzRF/T3vgOySES/xgOTVUXH+wwC3Wp72vTX
2hX2OCFddh0DKOyHyAf5Ht70sOGJyNeYBmREfvoeypyf3GtRgMcI2+77n6ETIb8A
QGYrvW9//xwd6jLTO57mBg/wntGdnRPMqMrsbdVypMN4xZ+J0W/oTBS5CgKSgqOu
XMBJJyZjGvxdhRvbw9hFDD2qU6lhD3M+RKWF1pQWRY/M7PgqKwxYtGbDwWyFkVcX
GF38mE2vD2rkwsK4pNkMx57+ooTjYPYOogNMFc/A/jd6KrNRqZPGqYvuh602BsV4
rwzWuViyLEX9uuZrebUSuX5nRSXYA5LgfbmK7f+m1xKsZrZi8BwDb2WsluW6xSVR
Z9SMH+U6LqHMH0Ac6BbRMBvUZDfbQAdZRyY1B3YJ5c8HfsyXc/Ml1JCbOaSc4mle
OGQjJ1CykueMVET3DT9u4kKS7LybBLzi8OJ5EStGEHkac45fgN0xBzU0xiIjJ6rQ
8kVHh/cB8gq707t+21JiGQN3dKko37BoTWAiN1LnwH2298L6r6kXLTZujcfa9pA6
1eQvntyIZdjpf9anPIFISstD41hmXZguR9dbD1bZNjq8NnLI4CN6dSBTqHF9d2sI
beu7/t22KNK6F6TkXKvLeeG9S2i//xpfVGLw/q9F1jA8fXePGamYksZmcz4WzIM3
to8NFKasO0UfPDFyLjeA6b2Apmqc/fAG5sqpx2g9L5BSjGxVwprcvZFlJ01clhWI
fJQUYroSejJ3Ie7ZAHH9l4IJ8kLshMKCMIrrrcFBoGUmyprdaNQLo4gdNxU1wDns
rRa8xi74RJ/8yJ9ifw8I1gXu+OWQ51l/EoRVFT6pSdu8pinBuqlAGWafZ2v2UY9i
6/ol0G6PJ68G44nOxzELwvqi83p8T77kpPBHqX7hdKQWDIbKtMNgEdD2TKUr2Ama
CbaZrq3z5ReBFcdcxIWyH769HJJjrB7k7O06WljtMGni8RR1MdQ5/NtSxiy/w3Av
MT3xpldjFQqd0sT0Dq33y1ToqfylHOFWbPLoZkDyYlALnL/k5NtbTt/J1Ssm+2L3
Axx+I5wrqATwU+NEW6P9cfr7USY3hkTL+gklgOdFpw3lrJeDJbQY3pin4Pp3DSlz
rSuHPNNkM2DBvv92YvxqnPoFqhlImBE90uC2OP7ykQxNt90F22zURlzBKJPuND6B
OzqgrGIBLoCI1JNY1Y8ym7vAOeOvQtpXF7ZJLyqFTjXC8JO2Yjy2nMxRu88tFxES
NZv1069oFSO6OHvkfQAkkUaGLj+828V5oZ5QvsWbvnVUbBiTZok629JMEHsrMpHL
26YtLSTsQ2Na3w8iEUA+x9+NjBJTEKWbEoEw9+Q8tpe/hAI+7ZReaA43qP5umObT
oyPrcw42A9uqDUxg/xeegoabbvkNagrkFKOQxmEk+1Ye4US6Z/JH2DeRtA6mlbMt
Mb0woQ1rx+EXMaYbELEE8QCOIoLQdczYQ+oYr+fz4zj3Rk8PosULeaVNd1MNr1x8
3kUT7xGnNMw4T4R6NeJIcrCK+WMZtd543H2z46FhA1fc7n+b4SWqKIxAsriTe7Z7
X/s2A37dhlWBfUR0WrEs7HiJiiD3MAQGieGECZiHXrrOV6e0aOtH/CGlXNHwOIJc
0suyy0tSSCjyQSHdtsu+NTLf7wpn0/rgmxWTT/wlicIHhdJd7b/4oNucAkCDrgt5
cGFlgpL6VZMHaO41i2vB+iBxtr12WERIc4KyKWTDy+f6DK8ylzLbWyQ0CVdDQnSo
fpgBRKb4Vzn47eHS4ThuY0+h7GmtMZpXH9bk4+ZbxC6pXTG1dScoPaRKXa10ngIT
71sGFPRzDYSczMBydl5KRSFeY3s+VfHiVBdJs+M9raoHmjFVDfU2SlflA22B5RDT
eLN33fYIU86sEvT6qxx9cPhQ+EgDuMmkLelKE0Tse70KXL6N5Pv9EzTqzKoeumPx
AHGO5sRNafC+n9SbEjv8V0Q5+nA68rUqbEMcLFpXLkBuEG/8dJKBLpASMFcNmX6+
7wC2SM/HArDyvfLtii02uBOt98+dM0zZHN0sf5kTNgcSkfMM5JX7fH69MLfUwiFy
2OpwUsR6pkoSbiSC7zs0TXmHdaLJijLGhIjbbi4WCkt9pMEjooyC/GIa9KTkYTIW
6cBU186by1/zMw3bHY3eqlAYLyg4BPDVaQ4KDS+YmAeyAeS4XkTISlXkhAtuUECF
E2mBUUNHyEP3NQY/IMtLzasxbUhA8xuZD4/I3/nQHI2G3vafF5UpIbaSDr7UWlgz
2pdkeILut/nnvlNhSSj9PBMVJ5WjPLWwe2ROS+TryNc42b0ZyhrCUDdmo4jZQDr9
I72o5IHj2wWatLDhpKrCnaMsUzjpqjdc4VxQ11r2UUbN1Xi3g0zBD1dV7bMcjF3I
6iDZd2zG2kAfBdYlQZe9cvJvvO8w5PTXhfNSiE6Tj3j1e+Ekinyzrkf58FyUyIGB
wLD56EcKf6T8wblRBoTOzKxWNAEZOmdayvlxBlHW36aCUtQ8ONaksibN/xj3G2uF
Xh+vbrcNT/dtvomLhaeR8iH/kB+6gEbi6bNV9QW2dhJb54dIfO+jmWF0wdwCHLV3
7tczAExTaUeBfBbaxaIoqOPCybpWPzM0kyJ3faQYVGuKlCf9VnArutgkoqipqqDw
dBNw25wwvKQOJww3D8QXwMliyHgfs5T+7h8t0YRGrEoFHCOgJ0x7DnUuNRn9uZs2
l5g4hhfDCJYoGm//rAM+0s1/reeKu5JZtWJFcP7gj4d+61Tf5m4ArSEs0uuxDv7j
V3s2c/nnafffTc6c6AJgtMFJgO19B64caPWrLf1YCi0YQ64KZ7GnxpwzQwumc8Ui
/dPgHejkrX70fI39605PvVGqug/oAswc4ESg/fAKCkT5UlhFQ+afv2PiuJlrvqk7
lPivtxEpPhErwp2NgVmC6aZWjmQ5b/XkZzX+RpiluYLZ1Lppk1s794ByF2o7TJi4
CCJwYzFEfcTTVDKl1IkT4YLgJZzmjJGp5HAgQYn2+9mtxFBSHWbP5bmxg+Kc5CRu
O3t8YicNMJ2WHfqZM6liL/KPFEybPR38k6xdbNb6CVrqF7Jkchg6plQptDKX75zt
vdKq97z+kG1y9TRECHrUYbthRGbhhY0sY8Dv0thJp18Nez6V37rBBohZjyf03Aav
q+10hfTZiVdshk2F0SMSR7oDI2+ST1WB1TBQ5IsmmAHIyUyLI7ebUI38GgVPT37/
Ooo4OlEO3HqkwvOmvtViz49Um975u3eh9bAVm1fu3YiWp3loAeIvx34x2xM2MwT5
mN8udBpsxaICDO/8Qol+lGzriBOkeS2/iubi+tvOMXZCSSg2l6XfWZCqnGPH58PF
tLcTU5lcF4Hye8BCN91f+v+UE77V3havGn0lchvdecpnTpe8TL0Dvj5f6jxIK0PT
p25RPA+IIAd2qlcQZ+WBaLY6yX1Q+0YwYRTXqHc2Qqn4D0gjeoxtqATjl/tFliIt
syj0MvFbWbLWvzD0cRD+ex00r+vkwwGcDTDprP8gGODgUmvdtWFS7DlWZOfVbsQT
ZPhvBX8x+2eYlPaqi9s17hOU8zPVOUxrD6lvMIeFV7EnwvEEpL2U4NpJDBbVh7N9
jY/ie/qGhT/as2OhpjcDmbYRbhj+EjsdzNfbCGpBuZeJ3+cWlXq6bE2ZfYOhoUdK
fcoyf2T2q41iFquJdpq6fRBbmWs+yyGXPQZlXT3VjOI5rnuQyekYl9oBKxpxUSzQ
RtCWPWkWGZpSzUn3vDEl9vBaRAHCTiCUf8ah+G760srOcpv8hyKrhRUmD1yfZYAq
myJQlF6qKxamVsAJ6T17nfNlpwRk7JrNJnT54pWG3+n2o2CSE2kIg895cc6H3q8E
Q4nGwM2ICurbbDdFedyhohtsxGLCP+BBUkLEosX4BxuE4+mQPKIrVkB2NcwER6Mw
/AvGuJ4Bc6AZ5Ym7RdFTVhcf0jCtsE121CDwlmgu6wDZPIPJXLOIuWyvkudZ976l
BZITzaf0s0u5xwPKhPIEcerS+onp0MAqTusL4gClnBlr5E0AYw134hH13moR3DgM
SUCnnLw+PkKLTqP0P8PAFt+Az1N96yTc3A4/5yDC9hUKI+WIO7sET61AxIZLPwVt
2lCcsmpqHFU1CSW2qnmA6rM1E+VSIQuLmUIFSRizL3l05w3QRjZcRJjFKQ4VTGfU
zrGd4Df5ooFTkyKItqhmc0hm0v+T/C4roZeX9pAEM1EtkBXwxr48HOo4Q4X/GJnD
3KoYteFJtWzPA4BaYKeTRHTvtONfPo7yNya/pQakSAYeKci4pg6EeP8eF4pgubNb
5lIfO79JISfvlkkcR6WKCz61cyaZhAQV0K6R6ZtrUFtpnyvLbRHulPySlUTnkjR8
I5OgRmZnwyyPKvtHDqy/fGJgugXfjeqLV1A9v+UOapC3V13EbgUBe/ssKKen6aDp
3AfDwvPGz8BiodhziXfaygr81zv7kKKk9FlCKR/hn9w8qdeGl52ptd/GGIi3bezO
WVHzA6HHkb2vHCAnmwSW5yHbvVfWgVVr5IQukpeP1VZQUwlw+ULFq9BO3g3sFSIS
4NFVO+hFxZCKdhX2mv/K4GcSenBIH88PnGy8eguGhDre+CxW7BNpSdNYjMUqNjNi
B5Ukz9YTA3zK6s3XYYREdJeHkCW/ZvVFNc8crnq6s2JFncX6qYrF/Zj4wRIuoezF
YfLFMhfZh+eVsRbuPU7tj3Fo7I8qU9AdILNPMuxDiUecZKXuUsR/1LWOuaQ43ySB
Rv2UUx31Uih/+9fFAMQU0rL+LFD5AUQPKO59yco5neJKjXm/sJdvJyIFFInX2hFR
Ragu31oK/ecb0By9noqMQpM+zbskd3Dpv8DajsySJtsDEcUj/OrVRUfBNGA7k8Zg
TAFbtgzbScblb205SVoY+spN7M64JX1rTnzBiYKZqwuTWomcuRbi8Oqjr1kPIVx7
bF2FrSa17n+k79irAaS9ZmAqsWyVNiJ30nulZc1xBwgPmA0TYT7xPBcn3J7z6JqQ
pIaUiUHt2cZHOaADScwQd4+WP5C/gwDi+yK9/cVxhtHVwpx6sf0RQ0g5BXM8ySdg
5+L+OHLi52ThD9CzQuJw4h1rgNSmMErs8r3bwgjlIqb+vqAD+Rylmx1qe30iSWL0
GX6zuA6MlbARC6SHP911dVFoBb3vPvHaCIyTzfUc+emMdagbp94CY36iCDNIjwLk
uX/ATr/qa5PgvIAUOPPHk6Ur9Ns6TS0/C4OvWKxScub2/O1nzt24VQSOsmDLCd32
a2golCCAND3U+cID327KhwS9/0Aiv7jqZkqiAWxryMAhfiXp5wjYtwbKZk04hgBu
YVok0BXH7yVMc/WiXnlFRv0KNhis/jMEtHkFPFBf+oVJnI+hUI0ymCcRPGFeOJXD
8gSSF5/w1vQJ4oykS/9rd1A9ZGy3fLh+1yN5vYq3Oysx0eIbX1gjb3rg9JDiwIAO
LdWV/AzkmtzZ8TWfCdE/S1C5ZCHbbe2idUoS+bAo46tcvxpsqV+mzTA3zLEvw3CK
w8LfdpjWX4QFeILFx8cOCcDy0AqBdRhVn8m1em8Y17Z7Vcau2bQ4Zpt1r5E1jbzY
37VATUvqfws3FOoXUgFDV4ZoAEClUCj+h2IIfUDfwF0gBCtId5qpnyzWrys1ciq0
hKFSeff1Esv6XNRYN0tTZXU01sSjtSLOgPgc/6SZR+DJ1jz0GUF0rRn2vBAPZa2/
Qoc8XReLid4oY5Sfrf9xv5UlhJcwT7q35XkXswl/A90DZLOaylQ71t+M489dGjrA
BfGoawHa0Ig/uVXOIVHSizE9HdT0ARqyz7hgjM7l4M1irA+jktDwhaFdTdBE7HH6
00rdGEpEv/Y02NfZy+kS9WSi9QUmg8q0bq3khTCaClnm8yqPJWWubM97XLQVMzQH
9PM+zu5YQD9DxQd0t7vww3Is6u3xMzbpmdkvF6y50pjpFnF7zc1bs+IJffTEUjth
mwY8RWxSNdJI1t+ySCqCaOSgPk9UeVhwoq5/FX2fVHdOOXpihf7MtkmqCJ2ozlcv
fkZv1yh+O9k9bgzbk3WrATVyL52ZO8LJhkffJb3zLa24HkNA8+c8Ge3poezC+QLX
lDRDxoskMtmI5Qw/L1rtavbubv/QscodLYn+Tn/0ZSF4tl/qdAFuerOcXMQRnKp4
eql7PVnwcliulbFwspwMC+XDwhfhx+BJlKZDvzY1rqOkIQgaPVoau1SAZST5y2yu
UoL1Hmjx0CBQqwrpMRGW9TB9ReZhXwDnxPGCOKq438FDwPfeaZWvxX8oPcqXBVNV
TxsRQ8+kxhDNtDFV9SNCwz8s5kGBhPng6iFNC55MJvh1p3+mFkNeh6kiJeiqpTFi
cUbhZBxag6JR1GDvpF4Hq3YFivWkC5Sz5n+jBmwyhX4gxcAnywqxv1blIQ36mUYZ
12RFthElQN7KtH3nQ71dyppN1UOp1CKLfeMSHqwhlAfXqKVZw2d8LUSGwDS10yE2
T/3YL2f6HDIxvowDxEb0E5muVS4ZxnuwBb3hxOQA2JNxiQwxv9cdp/pCwcfqYRZy
POex/scF09urgyaqJEw/b/Yr+vqSpOu0W1T7aQQ7yR0y+yewZrOgI7g5njP86sDI
Webhni1jODE0+pqUQYGdkvd0A0fbO6rDx8m20AWxy8kqSSMCyPj9iVp7tbsafUwS
Q9yiXgSYHSQZSdBATCj/BkSgV5ixUijyYkV+nQFvrjs0yCCeAKm6CQkkkxg6WBri
lfdp/JfPrCQ5HHRJMSlWyRjYsf26xeoNILmVVFHUY1esnNnWg3guXeLcEuYYwaZr
NBGTHQmiUIXb5CvE2BJ+xLv0Vy3yyLWlcFIHQnh7zDDR/ZJMsMT87X/Y8cLY7xTv
I7mlv1DtPJM3JRK6cCRLQXzmlEhoxdu3Ucxr6EH94tLQ+bioG42hue3cg+RjJ5gG
ryZbf765w5DEzXRGP7frYmpSf/3riO57jFq5fbpVO0/qFwJNuef6ulZOLsWKc/Kl
b0ranPWPcwGoVbfHnjh0nIYvJRQWI/IWcKpBEf7Rsz9sQR//KiN/LH4j5AOEjei4
Refm4tlNL7RAyA/GuxHiChk5Xx794ePp6CY51NtavbX2nAT7cdzSoaHz7Y71tevJ
GwLpFdS7z/dy0pKkx3FPczgpNQlWC0+5LTOiBUAAW4igCM085kQ1jPaNTbG1/0IW
IoFiE4v6sAmzJgrnr8CqL8IswVXQkOSOyWex5wjzJ6R5AKe6uq7AY01zzYGNyITT
atlKtPGIj6W1R5sxXKauw+3ALzEcxTYJZJs6AsxfDDXXZdZvQa0ZxSH6Yuti8DEk
Ar1sc/df4Xin4/S4VIuThpC7wn37/WFgiK5q3dDinUXMfHNUx6G/5M9GJ8znBYtL
Iz91q7hXM1hvzwnnwePOPbygabKFUamCgUyi9ZKmnjFcWxh1/UbJHf3v3+lvZX7a
j6gKvqAemw3qKJ/PgZXeQ8/HwuX5CGC7KsKJmUKQtJDcKwC/z088DXFbsrQmYm/I
Ifn9Kfqzf3gqX1NS1Y3iMZGyZ/25yC7i3IiVR3khHShdyfeapqhdxUmVtBYpQmq7
m9rl9BgHjL5VDt1XD4ECisxpbGsTY70b8czLfgh2JIedH69hMiZsWUelwX+lZZko
HyIicM9lqgc/9+J/zpFBtPcd+rcMKao4kTmUmGcjLNPZ9oi0ALB/8nN07e9UbtZt
DHI+KigUmykYo8oBHMBsnXB1NRZKyOFVzHS9hXxFyrMJKhOdiyzQpTYGmRYeslBM
8loSlC80c1SVRsKjZ7PU1PpZ2SvLAd1f8aU9dVppRd8ukNwRR9WB7HqO2WQ9pPW7
ckQvBTNKV9mtKegQotrzy/TJ3NJ3FXZWGB6hiQvO5zOU36Ie3qLDpnrB3CRt2nvE
zToeRpLACY1Ru9g6LU3h9rhtGB8Tp0oOfwSXNkA+NB0XVAFkAZ+2/tYMeHM+b0yl
pG0JGRwsFli5F0Bjezka9WzNyiVugCFytUPvlQwlRzVshqZWVvn5rij+zVM/A4Uh
+OOLrl6MyvaswHFkY33RH5d3YmX2R6ca7dZZhrdfEZvG14VgxNDSknKa9keP50Zj
bvXxDkbYx565vOpZR6vJ2yEctDGiJQf8rWelWrEiAKyY+YVCC+OSCtX7z3+v9HQp
6DUCyCKzwJcDRy+mdD9T8EK7i4nC/aRu4ZfY/ppkoD8gfmkshTX0ZvzYDKtuzpuy
nwVVU9qWmZowrPFR3iuesmtTY8Y16dsz9wfsQ8+BwVFUhuhKLEG7SQsQ40Kj3LaQ
3avRoxu6/IYxBzQSZTSRibsXHPLPU0NpqkHDM8MzHl5+aETs9zRKS8/M50puSGm6
4BxrwJOTK6RJswC8gkuYH5aZNTjnAnBqb/sUxdAkbqFGJk2bg8pOayJ6JybVrMyI
OcudGLxvHlwgyYrXA/cjo4sYIZBJa6FciQT3TaQM8Q3IHfX7gziVUfmxTuCh3kjs
MDxXuQhUeEIncuLEa2iJKV42FTY6iykgItU3Nvqz9ePZBr3kJlNm/PF4HlTEH29D
KaABhIFwwHVJOjfhrGL+uqXL72Ss39qyHeb9FrA/RUR9s3bJ/Y3uJkN0X/403whV
WOMqkTcjzE4knlmOgWpJJ19hN4cUKC499NkNb1EI7LlUQoHRvH7tjnkxCiVp9cJ+
H+m01ZKsmKorQ357TWrNQ7b/7ZgaUrvhp1JikFkCl1RtOtOcsX03frPrIWLdQn6W
J2ZrCEu2SdSYmxcDYUR30zA+ilnLB2bnXPEfxo6Zh5LykHBlZcxHD6xHEHujXTbd
uZSRerb7cX3jeHUwVfebknO1Fn2q7/fUALMJMPAVUwlxsyV6gDi6Eoxx9vtESve5
GRHeb+sx1W00vOlhje8rjhR9ZC9945UscgbYvWtMLhyBOKkFFBNCgwqDODVwp+3V
bN2+1R4b5c2OyK7uMpTym/8/pPmEq1FbVqn1JTO0M/sjDLqjJ9vhfsaGXXBStnJS
e7TrIyoHzg+ELLwBgAXA8krn8DrTmu/5JbQf0ryyxJxF1r9aopZUeHDG+7MjycMd
IYAv31dlLg5nplvSMOycNhOMgFJ3GVaIf05DH4zA53AGqY/GBZDyIImKsWOYQt2g
d6BrJM8d4eGOheg54auPth3N9VZl4PXDyIkLu214CPGUQsP/399VWzGG50B86SFD
LgsRJT575Ff8P9ABkcjrxZX3BuyQhcTrkSEs8Es1sD/YBm2bUiPLG8OC1fBg/Hg+
vOH1xlR9aYGFSjQ+cPaHbqg54EVUEF9Jn6n9tYJbc2Mo6+A+bPsxcOJxaBGpWPMg
/K6l7sYAg+flGCmWL0X+hAnlT8VSQEyaTy4HwPw0pTbONrH1KuCg3+e7W2jUAhHo
z3UQnUrtmU0f1osTPAonju2TkhrXe18KILmhLvaXDHfYnA7YsS8+SAv6gxY0pfva
2sdQjFIQcjrp11wogHxt9+/S1WUsekDKFUlbXq93hlyVJXZmfIi3gKEe24vx33cX
JqO5muTl+lSbQvdnAUHUg4dVEdto2QE7KYLv7ngnTH9KdauZ0sgz9lP67+1C6sTy
W/6Ew7+cAeAQ86lKnipARzqlA8gO27Od1tp9nrFZabRonmjiriNNQQ46/9eiMbEW
qYsp27aMcWZ5jv/7ToQUmWIfu1Z+erU3i3U4nQ/ICksd7u5eFxKaj2h8xUJNT403
ZDM+/1kZkdKAr9kMfX54OCxwcfr9K6w7gIlcidm/fOQzpjyT7lXfwpLNZQJjN8ch
vDtzoGFQSyp2PrCTkS+pASSGa55SP2bZ8rhHKD0gEmApSOdLl3cd7sFCbQZSD8ii
LKL/J+7A5IrwzG6bZ+wIusoSJ5Eqmu24TicoyK6sIZlzSdt1bhmQNlJ36r5gIIdQ
BchRSIWvWRyWx8EqM0sMd8Y/7krMpiXQhjAkNZqPwe+ZFNf3gsCaYRBXXdbSE/xc
5qq2ueaQAqa/SXYf9L2FuuFuHYV300qGqtZLVGTvtfH2lLBpAll762Kfypks5RAV
DCtaDnByoIuwY4LfslnT5wkv6TVqAGNyAYUmnb3COZHDYDauiwzxne8bTy/l669R
Bb6HkfOMhoQ+VugFTXztldARu3EnQy/CLn+R6wGB3/HrAl4aEonA2LDSl1CpGWZp
o3xA9Ex4e/bcVaU8BZthYqyPYqkO414jVGTRE2uBDiEBPghe2iVCZRK7Rc1rMrRm
DiMCnFTqokdeNJNup9dooQdQuUFvbr6HpTjqi8j+PkpAcbVq5/Yqqed+KgbpDqC5
l5KWqXxAqBJShej3wvlivoimK1b5pEY9XPXbUgqIV2BbpSxKdCOOxVPzloL6rtRP
lxCVNKlrnAD0MkA9TN8p6uGWvqveYH/ZnyHmSY34OeNUjAi/IczJTrxgVRQC8cbq
gMDrPmuSQi4NJstMYQ/4XK8nDoxPyzj3tj8zyGu/sisyW+HDNDjNb6jjqO2NGWwe
/QOGw7ouDG+gV6xjEp16XFClALQfFEznfrWdBRKPEGFmc65MS4wh3RdNoO2tPRbZ
nyX8+gTMTOR2+Ka/guU7AS5u7/jsUdkvYZJmlzQeatEzJtC6BnNU+nO4N+ysKnFn
Vj8v/zX9Tn1qWY6uUb4m5OgAwTmFLkGZPPviykWDirh928FppERx2reJEAzrK5El
q3gKp5BbkgFkaIpC7Ighec1GUFouzznRY6lid4IjhCYDHdHJBM2GsQb5/3cvGLaZ
63a+psbjXl/qias95aVGQ/puB4J6J/XG9un9/ojFlfx/0cQhWfXmirh+uqAd5lqv
lutYgMWH8MOkHhAxKpQBy6NVYJEJenDDE2bB19Xfdwor9h1w/xFwkGaS0t9evaIv
9u4N4ASohU68AoEJ5qyyMQbK4ZhByeLL3/yGSObWz7eIC7+XaXKKQE25SLKimhG3
O8Vk4X84dPhCBUkPGKPw1bvtN4Hpbjn9lzbhsooJuIUcq9+wkTMk70fzDu/N5xQb
ehOaKH4atissih2+B/aVRi+dpIfcpUO+WdeCWYrq7yJSZARXQmX2XWmmozQR1CDG
uZvzg+GqVSODOctK/tJDqk25zB9gx/iE2W7NacAhOIZkdIe+LpQvbYNQkqyRcjpp
QSJCtTVa75681zKE+v8y8fMJg1v/CbhIVCwyrJ3IwjLNyg1bdBo6nEkET/WvjW33
KBPwb8Q4ihsHUTbUD3iTzZJ/IpqyFMMQnWycuj114IXq3eEIV9Gf0wCJx+CVrIIW
yDOCBondVZCWfETpTlcTBzbw07Ff3e9hS7ZgzFYN34vsKcvhYbCZV44VvpQv5v+Q
X6vxEEMFhVW/mvAy6meKRmC9stJHwLBo24WChhfHNeAcahJZHKngrpINRaaZmJ3P
5ufEvZkxR3yk89aw8nveCk45ngCvke3qb3XHd5czX4PUXjmQzZ5mOoPShkjBGqxD
gsCsaCkL84jzHQnL6AFQAPsa2NkiBe3qfhfMV5QUw2M+EwF/qulI4sIMmdqa5rkg
w4lzcanHY8Vpk9U/RR2owCfo457rh2+H2qAM4MWZKcuD+NsYVgQ0dXko5h6uSsMD
F+yFRAcpUOeDRT/7uCoQeB5/Gr1j1fku/0iWl6SwjuHFJKH0X3Yziet9XlhooHGU
iedFEb6MFAmQp8+CxE7qxidsTxDc9CzMFetnsPPg50j+mi1RowAAYBRH1PD9RuXj
RIlpPaTgjSPaSI+BNGTSrmp6ZZPf//Kug1CjdQrSBIhwlYyMq2h+1E0SCq4u92MV
LaKvlDw24GJOwHkUY+77DXMJK8Ov7Y0rRmkQyFyYCOTxRGi8OENWavVsTzgiuTjd
KH9w4NK+OM5oO3vi/14BFdyx1tqv5ey2KNx7tuTzOcDW6mWU8yxW3du2eOUj6P6f
0fUZGrABrSGYVTMoOdbWdMYLitzBaSkbgYklmnqDbMkKkkijPxpH8A1AcvX9vQrm
FA5t5xKj9Na5Hb/4kPZWC9hq9xXGvRJu6FGRK2WJIpjkIarQ0oLkVjcGMiul3zgC
PtHfZjhRkUD4euGMQPbIF71CUrs/cL3LvSCjlSD0G3cuuoBJGcZrTLjwYZ4az39F
myaq2dB+KbgDVnhT4UA56RN+iAwUa2O3a51zK2JyjvFSZPK/KvRCnpNn7lZ1CDy5
vlSpERRpax6sN2WOQ7aVv2C/gudNd/mnhGGuf61DiKyb2r8hDR77It8WY0vbsKuI
3piZIzwWMv9IrIp8nl4C+8Y+7CA5UHPfrLZunk3f/10mHeAPQsk7j4b0AXJrrIzM
OWl4EjX4dDlj/BV0pu6QL24GI/NjbUxi00A8e8Pxy6lUVhng0zfgLyBSYDso4iRH
/4hMMhdIzNs9LG66RkTWCnxtnzleNu+Z6Q1idcOmTlmfOZiTh3hdl1ONo9W6uI5e
ml9BOQi8CetmbnnJpDDrFkfQ1nZbMZ8lwO/Pd3Qv0Eib0xyTwtNzoVMCOlulSmFG
h9SK+ubCpYy1K3DumwWO6f+uExHLI6WfiJrT4fd7M8ymLNjPR+CpqZPx+R3R+ba5
saT4gYcWELXk7jNy96CGMDFsgd29L6lc3oW0WnRdO1W5b/wwEQY3Th9Zdgj4mm0p
RwQaybfKDp6jfCaoz+vlwqZ7RqKns2SBdzR34j1tIsFTdEGBTHhR6DBWXqLw4z+O
Fq0bJ/wBiK+VO3tiv6IhD3E2t0VEv9R7DcLLitBYq0mi96bOYtjHufVRJJ5nPzcr
IXsc7WkShNHCMxhqOf3G8iqq7TX2V6oma6+Pc7+1xyN0hz+Whj42QxkdUaz/rAwx
c7fncJ8bYJblNsMaUYGjfxvWCApqMLlDgHQ3RjUEZ0z67mERqnme3qPLMjGbf5EQ
Uzq30l80DtJiVaWUzXRqB7OKSNKgJfHm6BiL8c79bo5VisHqoIWxR1VxpL0lcIAD
UvNZzUkXfgZfsP3Zv8SwCCq0MTL2OpiM4TgAXJL0Tzr4nhz+bmA1obprD2HF5cRF
gEueQDzTsZHtxvrz+yAT0xgYPNKlKR1AYHGMgH3ABKYuHJ/NiwkZcO39XrALec2x
z0O1bI8q7Z6IfsJCv9mwpF+Hs4Z6MIDaStW+pEoNyF/n4mkGiH8qnYEY6VjqPEFX
hJbxzGMjxRaWKPqRiE26oQQqD6NIUhp58BBx9cHgaQ5J2eAjyLVrpOQ8Vi1+OBjF
Im2bnf7NQ6rhFgyAzPH5JVkwXK2KOnKPiiU9cTzhh6qVji/aY8QQAv+Zl6RAGjzi
fDy8dhuBOfcUXCjz2HSvDSxR+11MQyxBE0OlX8o4jz29+5pNg7VckdTTuqMait3E
YXzFfDySg/4aMH1cEseoBVZkTqToSP2qmG92CUTZCq6XJajKgnZtfsNX5ZThzeIV
V1NQoGD9OA+ySJ2Nn+yKs3D6yXPhp7xhV7IQLv+CZqSMqJZxVi84cV5oujczkQpl
Ic1/tYndZlxMI0tN3CzhEgjAPRzdm1fNaIahTldbOTiBCiVRUbpX1fvgvFAU1Ebp
JR9vl9fj53TD/27mbrxHfHm5+cEiw+3lpAiy9jzPedoHdSJ7dotrPDUVS2JiAANT
DH+gQS9KswjweHCJvDbOb1YkNfqAFRWcY6Uu6ZYJ6ccfThDP1syT5MgmgAFAOHF1
Xb6GwesU+UUOXRUITGNJ5qaLb+F7oFzNtyz0TdMU1C2o1luWn/M8YnRKiBLJIj9O
5dt4qXEJZnSSwrLb3HJ+9SulC/WLcDyTB7Gn1KLmpDehrluoQ/HhPtWVt88lLGqj
c68shbfRmcT+G0twSn8euI1HhomO/cRI9Dy3B1qmL/rdeiNjdja5M/NgN2UyIxup
ZZW5GR7fSRnL96adqall/iqBL5uqgZW++qLwF15APhg3MHUxbh8EcvL2jOysb3ga
5ZUB4iwIhsRcqwTjrW1IidEHNp4siwqVz0aNr7Nd7bLaj/Q22eTY6cJEuGJCPo4R
57028KWx3YBtg3Co/c7hHIi798vb+CbuBSsyNe7L23Omhcz1loQu0pe63eXia/4V
ql+e1j2Pwf1Fmx1dU8lAP6IaK/UnjGj2/C+L56wcIIZiBZUInVhtcMmtC2yQDghF
6yN9C7xf6Xzb8m+WZKQpAHGhBUlU2o0fKuqIwclWp0LJ+1oTrxYwnJvsUwOUGaNz
TZSwXKGUUGjXSg5ClWZhsSAZBPKg7QqVUVk+rfoqqte5bgf03ElR0PLuBho9e0Af
zv9C1d1XW8kKPXb9Yf9CtqtQCwO6tk7XiEfERPp4TB7JdhRwESgTzopp24A2qlzN
hfeKNQBTgdpVkVIIDZsjUVBSgdlGdZv9rmp6q4uvDvdsQfM7TMST8YJ5A8lDNHqT
lZ8xgxuwYlJr+jhEsTCkNAQZ2KP6RRfnvp3FyOm62GaMEeqgOnXlCLEUvHWSOgck
3nkAgf6iYgQWkl8h4U39Y8MVgf6oqzgjralosgPTvpKxfOslVEyEBKlCSzoMewhb
o1UuWgu581erYy0e5/gfbcdJsHnXHcOpszpppIgqDMg8Mkq93/fK2u4Xi2QsKuaE
p2agUea0BEywEtuX1ZaAz6pyiGy0ssD0PFzF1tllTsFghGJkkxPZLj9LRiY7S7/1
95UIo8OvtEDdvfFfWpdjRcpTRhyZZ8M1mblP5R9yQ2yvWItwy1EhqP8cWDwMQYY2
/JiZDqw/3gKatct5dzqT9tqBKAEG4b7dJxML045vpg1iW/kGIDds4WyQ4DJH92/y
Jx4BCbyRananCe0WybFN3EE/WSP052BxaHnxa3ZmHJXwEsLyIR9fthj1onwvt294
hy6UYvYxhAVK7Sne2Vx6dtftnD7Q6yh/c71REEvPP/nJhOVR6uW8VStWTTRhmBAh
7ocSTCavPd/VHyqLaU2PI099Ij8D3ni/iqHm5HjbYBaKguDbcP1ObBUrXxI29q2b
bBCekZYcwGg2Xf/ee0D7jnwRIbW899z1ff+V43REoEYE1Guw14XKaDsGSYtlMbOs
CjgFgokFQ4RPvjq95BrTLKEH/mzTtfuIqkb3eCxtjTUQZmTXxYKJVlYTHCT2b05m
p4PJiBiqNcEQljb0y3LRcITP0OhBOR7VcfTdX9dofwXCmig8MI2Ev30tY/r+zHHF
kTIAyDuduZ5AGzmTc7KxTibhfVGxLcosLzSaf3Ma9qGdm5S9gLb0Mqk3jQmb4duN
YI39NzsgsfqmjW6qvdrtoBWJnDNOqLnmrxfT3YSMHBjJAvfIj0Lce//XdqxW1ECI
DUlkbhLQZgwFTNsiWuI52bIYLyOmOf/rxzrqo7fAQaeKTRZuEbVzJQ4gMh/yqVxT
RaRkkEmdQsJKWuHwOUpmJ2Hq8PRftc5PuaISaWTsSfQgZ2hZdU2rjK2vxahAsf3M
xXbVOix1ANWhcMe0CtSvVMFpYq+w4p8+NVkxhyD5E5RDldEcmlOaF8ceOb9pY/Re
OI/RrnqoPmq0D4c6hou2W58+9ymzcK92mH2FhTquVYjfXrclYtr83sfc4A2JKTkG
zjv7peMf11XeQt6kx5p2RuokpjlsdfuJf8b9o+Maf82escrzaCWFBo2+M2yzleKs
E9KgldNjJ2SBk6Ld9F2i5RjSu513CAldhvuBzf8JmvLkac8YRTNS9SmYbxwL03QX
HXRXLttGne+45NHTvslr2ZrBv0Qm4Mc+9pToYjOK2gobOLPMJXWigMP2fxe2k6XB
EgaslBvLabthhths+4rWa1mhc4giIcR6mKKlX9JrP5EsCuNoVeMSupyY9opncQYI
nCyuyOAowBCIZ9BLXze8pxJDGHSlRBVtEwnWCtu3xuIps/dNzfkMwtmG5DQFI2/i
qd4nxORMQIizM72IN380w7g3UMoCoxGuAZ9velB9LsKIkpwyJdV+auYqsUXyxMQU
IfbWgYDO1vim0nsLql+pPotVRNfRTYWNLlTbYkdVfuZ4HZWpxcOrSaibdX5AT/jp
s4BKhnIb0uvP0ljedLF1q45CFFZNNBozerN59qJdN/4s0zA0Jo3NurMVOGfagn2a
ZAb2X5+icpUaeoa9WRHqKgtNb16Jm49rd+J6uj5sSjV1Y9zxM2euufehf2mh3icB
v91pE5p+BLglOU1oUx3iigTuToILHDk4sjJufpw8tYfNkb6fT8rZjXTbICEMhVOn
ta/KW5HclLhl+4qrZI6ccYiUeV+MoT5Hv2ldpBOE7k5lDYq8Tx4LwITXOjNROccP
wAprJMWflQjgJ2r1wt1Y/bamoimBssTBQ8kgbLkpad2ayUYZXxwrOizEcKCQk72D
WoHyU965VhP+YDT8AdEq2VPNKPPhp3IgKBTfwhw1xgzrCAhSc+VYYPxvbQZyDdAG
p2EPzqvX8Jqf8RChSLFqBJrL5HJUs9MoCE6av/Y79qEmaoiLZJgpmBxexmc3ZSQd
4clVyu6qOt8/9kpfiG1kCPouK0sK9g4k4CQtiHuZdSgqmq+lzx28AoZQ79OEH4cI
VOzOWyx0dWRGmsof6+6CJGTubpfL6/TIdLJFsiF9Uzkob45T3P23vter61Tog2+N
FLjNDdh7DRKluWHVF6ZFLxntCjwDVilnAQGpvlb/X9eD4wx1E/jFUOyIKVFU/PXk
T5hNbzSkq3MF+9UyI9e5ZOxkI9u8IkDGhtylDicq6Rh9kTOf8dazmknwvITveOjb
b7keRt5RkGp8r866LG5qhDvqWgjWq+yONvl1xBbq/ggGpplOWW8VUD811ogVxfG/
DpvwR+wtRp54Urp6rzCK220iIc6iMw2afysgJvI7IBSnocIan9tFO+3G/l7N7jhf
tH3M1d0X01DSxvXbMUeuf3ru4SlwnqkqMeT2RKnTvYEsvMxNVLvFu3RI04ayQZa6
3R+4pbwxOJFuOtEOVpFqq+IF5rfgwz7fHHR7ERmJp/S0EH6rH6bQw+bS0e3nFiRf
WXyazAZeaW50teD2OmzntFQ3Us+0/3ITfySGTFs+pdID+ezO11Y0LMfD0AwMHGJj
UKIcqSRjk5/1eeqZf8QvS2+n9fkp59sL7sDwpCNCbW1Gf0MfSwYcrR2nWZSZONNK
ystBbO2hM/wNhDsQ76+4EVEJEUNVLmXY1PXruerGcYWYenu6RKdMe4Jt37HrgHUu
TVC4k9gudKetAyyvoMcz/FSsy0tzmwy+rXkLZgNQsbaiAfW62C/LZxjmZmsfodO0
CR7Lh5VW9PGwC3p2ICJtIZ9jBs3XaUnsUO9XcFIZv91OJfXzIpCraRiIq6RkxxzM
NkMFpR2tOgzhjJF1+PKMBA9tZGkv98uA7Ncws20p4wbXG09DLy9Z/48AR3DeL/cC
GHglo0DLCO5nyxH+WPncDFCPoqM1ne2SyuZDzfrQDjbegQZz0GIUf/KDZg2r9L+a
5bFtGbyVyJ5jBGYdqESTQ+eJ0MI5IVqRR/gYkf76eoWCtzjetjcMrh8sQnLaET5C
yhYy89y/jwimREBTRtqyXyw+HWRGRSAb7dd92QfZu5Un67KPdLglmxQCgwA9Nj1C
qHMeJy/bgesX0JyM4UeQQBBlEO+BLDkn8ff3+vn5PlqTcGZmIxeHTd2r3H2GXHqT
ZIjCY74g55ctDdYFZufJVoZY5jxFoytFYlOab+E7CHMvXnEDIK208ocVzIwDzCGM
9eyZx6yPrxpoJttr6gAOWB1JDqWwytlH2UfQ8oCVBR/cKLZAFm55qblhwyLNPHoh
s2lsSBr/ZRtudVbv15Uyil+z22/7reYiLxrQnYDaLuNE2W0IvTE5PdQMb7XrjwBd
PtpHrXjIR35A3SHkmiESwbAqsiJSmJQBKhq8ayVZORvT8Ry3OQ07w2jV/DMxCHTF
E2+Lr6gyIkERh9SRq1bI2yb2kF96zb4yJj6jzAN2D9xD90wrxFAX/lFJ8T3+TUqs
OEFe9G3RLTr2CBpuM27vLWNaqZad77yPbZ4lwDr+qOm63j7n+LyoKz+vNftDEmlX
NkOgqf4E6H9/a4iD41Mx3nBSqzV4OkyEkIx2uaWF5RTH3J+oaqfzE0DDliESIduD
FjwTIm846Ahts+ypVi+qq7H7EOqoGaZJYiNeFLBsJHquMtdZ14+o1nyR9LFSrn1h
bMcSNSI8aDI+mGRqHO23aVfFcWNQtry6uKITankWPrJG74wrqAE39p+bXoClxV85
SdGQaMAq5ypgSpn7gX5pdno4CT96dKvOhlsVtjnXGVG1CKhDYr91IgqivKWI4iIL
dwIgKO5tJD8EJL42Nk/S/nkMxSZ9cUJ46CeS+zz6GFQX1WG3+3UiP0TOwcwFZTEb
Qii9s51Uce3cUsHxG0XxhDhsaYLfcbE4npWpefy35vRQJHsHfYklSImwDbOzS/fZ
cdBpaELPF1Xg2fGSytb+7D15MVCpcfi0B+6C0UpnkwD39Smrfbha4pTgia71NOgC
itAsLxpvRfvAkd6xozpDhidSWEu0jKUs5kUAehxnwJuSoOk3T1jOuFLLJiWNq95O
vCd/Rhzjco2qMfNyzys6C1D41AxtUYjPU5uDbMGdLYCGwZuUl9xVRqxQqU/FoCqH
6beBwjmgCZPgh4+oLUiY327f5o3O5BQhn8k9lTHAVXqYi/rgfw7ep2K17TeM3rjU
ErP5PJkm0m0kkwAY1ieCa7xuRDB4njjzC+5DBO8V2yQvDcK0KA2nEjHL+Of4Sfrd
skQAhjXGMohW1wsSRu2G6A/PFel9+y97qXmeLMHK3WMDn3sq5pST+cDRxEI/LncN
A0pa6I3z80zlQFk5nIHdDH2Nu7+GsDn/qolUDz5UmJlsw6fZx93svm3YcE64ovyC
Mii9IFrrJYjjP+yrHtuun1dpXZSIUMB3iA3Fk4l7WhNRF1XiYqX643c9wEgKIMwy
7IexBs7SIYBkAqYUX2OovOjZ4lI5D+71ptgZKR8RkUpAbaeRate1w7bqQt9yMad5
NoPOf2OgT4pmpqNCxv4O6NnAOpfjStYLYbQw0rDshL23rR1YWJoemzXb2MJ8soFp
jQMvpzTyqgPOkYvahO22YDCJVLyNNiGGbNuhh/kCOwxknNAGiCqoLXekyQ3u+MY2
dGeQzpnp2NmGc60sU47xJJ06InTMWYAnA+fik5Iahvrf8/fnA4ENmoO5HhsH+N5Y
QBZiZ1TYyRoL19ZYgFNcokCp2eC4Rbi7MfvJCHLr9uVSGPI6FJQ2aeELYgEUzUzK
FWmbTJR5kfa/XAJkydgTeLeMaJ5u8HEkzq6ZIOSctCNfvvEzyEICkCILArHWw/uy
h5uN4Gs/71aYmk2ZtbKkQUAGhk4BOJAu1wg7lgswUoDxuqzI7o+aYxcBHsB2cweO
suoP5kXDZgaQiZkqcyTzteaPKDUWoqQNE7o81fFs2NEqGVdhSKMTYvz8yhMALouJ
/Zp4aAZIP0Q8uoOkC2FkowunnGBh9HGoI+42YCQqTIdId/aeSQE28w781rAThtrG
biOZ5skCou6+YlgFu98HFsMIrK0itEAMyyE8u288ecdWwYrGV+RX2Bzb3ZzxtV3E
7ib+QJ/dD3FsVbbxZrTTeN/gpiCMCwInOqrk2YlXsmVCcAxuW1iIp7DpZM7lxMn7
9njBTiWbI5soATO/WD5I2eFzN/BpG/AZMfqvZMpvE4eKdhU40tp77SjJTuuqPGiK
IAwPQUuRC5uQgKXx8yWa7updc8Ndv4fEA7DnaI3QKNr/CwHGJRGIBxIMZNoNQxr7
c+MUpVH6M9N6XdjBfsweL81mREhX2EN2Ldytx0ZrdLsvr+cjMezW7v+zrgsqT2Zs
DsyuADKPp09ipdWjwV/uzowah8+2bgP9u6dodWDthdRz1PddyJ+Na1C8pXobS2re
xhadfhggrCt3vc78EVJATfWbgpYhkpMSOFKIGbrSIbE3qG6ZCwL/1FCuO2ystuvP
IKrajpnpB3ZV/GNhrymsRuoRsupK8gNTNBvF+QMD7VqXCzTqCUFCtvCwMMMH4TNZ
v3nL3kb3xhtau4J1/fxD3zCXXkIWFv1k3j4XDQuhCYJLT3QSqzFpBlOfKznleV8T
kk4zI8lsa171l55ym8Bx8GnLghcxXVczjrDZ5z1ldhN4XJn5bK/lvF+2OT1ES/Lw
+QHHx+tCwKQhl8ZKuzDkCBLDHkNAIO8RaMC/YLHo8kF4J8OkZqpm0wiiiBrSmklE
49d9IGe0TrLX4Z0+esaUt6cYzgO5vFrJZX+Qqbik2N3cPyP/63ZED2Ye2XdK/QAF
0pSg2dxhtwh3rC1qip4gNYlUPW1i05X2LA6OEhzPFQFwkXRc9P3pcpEzy4yVd1B/
RzguednKj8Mo1D0GDloJ85LF7LTWq37jVhTPBjsyf+YVxZTOwYdsYCj/RaonHyKq
RI+aeMKjDp5eC7Sr7YB2oSI6YyeGh+UznmPfgghKcUMf4ekJw8JuR3zgBRHDFQqP
ZRFyDO8EU+JvCNx3EoDyfg26YpyPMKarJNnDpGZmOVgTEtQ1pDI7f0LxomugtTuL
VTor9YeKlQGCCbc6nNaicjuoqvYQN9IKKoArBQmn0iS96lcU30pUqlT9zODIpC8F
o8egIPZATd1SeYZaE0lc3PmkQ32I2x0I9M1AUbPMGy16hPXQe+ESRba/ZmzpBMHT
G5izG1XGFD8mOTz9etDwB74x0bT9halNKDDIMLf5yh9RYDHrp9dEXgb0omxClAOA
eFOC0yyOwy/o7YXL9F8Eq/4OHvDy2vrR5Qsu0z3q18IYbQoArd6S0PRLWFeBv+TY
bf/ve8UQdPGm9u4jANwoZBL7yJ4Mo2KbPFCLZwvXdGibueWO75E0Fy9lo1n0dyWd
c6/p9MWQtvvm3nBRcvYs971WoKT408W2OGC/7Al0doFi9Af0S5+oFg4XwHIr1HZt
7sFyFahaqlPb5NUDd5Aen/QuPnxz+HliYGHl0tylpDKeCQsao+d567j2hkMMbl9B
z/2CEK4KtD9DLmljMxudiXS7zWejZK6PXSR4fztYPs3i1pZ6ozGnVyAbIYWCknXn
ANvqYxA8nsBetP2n+1hlCe3qoq3UdYbKvJ7kZjvfqmRidThfpUOual2UmIBPfVF8
lYdWego1Hh2cSpRAryFPv/Fxh6CBV9tKDTkc15t1aSwb6uAJwTaBtFqwZmd8qBz1
2AZ4iaR7F17eEXJKiLFTVaDstMwhmuWtJ4iUoE1mhqVTT28FzGSa+NWAckdnK6Z0
haWnGcLxYL9SfVM7M1Y125KWqPWcDMN+p1deGUfosXSx21C7JhDufX3ShujptcdA
wRa+kBPuvjtFNVEfGzVBb9hOlunTA+W0t0otZLwqR7+SsKeYU4ETZj1BYbViqG1R
oOgy6ECMxzIJTe430sO27OArVBZIc/h+pzct/WJDqLopP7EVg5QJW76U6yADe8YI
V6XESJbvvZOMtUCFatelWzJhfnk0IG1ELTZoJ9twHyFEpC5+3LKP3KohpUDWDT5A
sT/8YCyiHbcDJ/6kM+/+Do3hqYrVcAIxua9oeNgJ/Ydmt6ZnuLx5XplueYEiB1eQ
RGD2v/mplMidubJdS7lrDFypk2htqs4i2eqyrVZnxu4gaW9ZvElzGb6OPUcSTQZp
MQliQHeCG55W7t+4KuHVY2OUbyz+lEXV7ZoJZMckfS1ZMtxBE8nlSyT+H7vnY87q
AHw/bdzfxuhMooLOQCQoB2oCKIZTPiX9j/KcAMqOz60Cw3Tkvv49/aoRXAbPHH5E
5lvZ/jNejrZQf+feNb21kmbl87tgc1RFczWZefeeLUf8Tbqr98ULUYDy7dG1zrC2
3w+54V/5I6NRoQJ7Jga7dAhRxyjEj84ubxTLVu4xPrLOUYvFeuM7iv5mJhIVBOfa
3tnuDbEEfn6V4xciT9y/V0EEpU9jprH9mUo17eEE1ahdknQ/e01YVrhPalN8PDwF
JtTuxFtb1kOsPq9Wz6iDGMYaEKXLqT3SjTaGudvsVOH+OW9e+3V/XW7OwTJW+eU9
v6L5Frw3xWFgOgr1lDeCBOd7h47Gte//L+mOF8kJ4J2RHmBaqasn2Vr11Gfloj1i
xY/NTopR8BDDvlsbIiW8QBnQtObRc9UZVydR2XkwsP2tJAsJxGRA+7x0t6WywQWA
38wRR6o3cQlcVvNLynUQmPBHZjllP6VKNeEg58MnF6mnSJDREKRuUz/y1cwh5eJO
NOk2j4vpPWSEqxbdmIINoZvbOvg8N/79aZLzMx0RSbBT++4o5NLSWMj7Ms0XLE4J
Z4PEQ1yaxtV2KLRih7rvj+THQ6e47eir+dQBLEP/z/3TnWaRLlwHz4rkr1fb7HLM
yxRD2mPRLzvlccIqryHyrWe3puU6YnOpFZgUAwZxavkJKceu3iC5JgZFj8FI06m+
BATLgpHQlXDL/0ipf1eNIRXbWVXMoBmGD3XD3QvAnkAWqsuXl5GVfn3gJDIGFCsL
2NrypIV4w5kVCVhjXtZKiO6jLComUVQi8CeJWEqqp8qkyS2JtZT8Sg7xIWbsAkEX
dtCN3267JOFojxhzS4ZJgPl00zH84bI7jdquYZtzRusEneYm9ioEw8f0CcbFQWM8
lY1LNJNughxyM6s68hpw7oTZLBc/eH+3fgR4KH3P7EIyVjKCrv/n7LmpRIebmg2W
qc51U+gMFikIKzZoqDkyEDerafYrDRLCLk+8uOorlYVP2eOShOQ2d73TPRYBPkzf
PSlOcg699bp6IRe91HZ/J0dxKaeAzsF+797UlRPGaWl/Y7hOHCMqqnt2+QflxAdK
jJ5hEK+cCBWVBoVR9NEZ8A3ZpAGZN3qHyHTAmYyBs56TnGgTOYnrEhRNW+F9kFTe
SWefEfV37qJoog2zOJMP8C2981EtqwlPtyN30yt57QjymbWg21JXgjICXQfMQ1PC
CVql0G+/5rJWgsMmKWfrh5tc6EuE8RoEPgyIQZGK+H9k9Gq0lVOiEtZcYDziEg8+
EIhUbzWCa66pT7OzrekzpHclmGI+alsQUwszAEzgRbPTD9kMuhdw5GfOW/ZuMnHh
vi/59xjT4LDpPausMjqYDaU2JychIm/r6P4IlWBHB5KaBbMoxoxuyhQcKjm8ZxpL
AFSKgMHAqWz4xMw9m9u6CukxZ9xxwzXHOVlw5lArxL7Km8tCi/xzlwsz8s+qcQtW
rgUN9D3p0cUXaUOg0YMQdxTMAU237oz5GmcLM38g4jl3c8L9Z6wHEf4wKD18ZNHG
/CZs/Vwp14j0KgKsgJU+q1VHH7HaR3hPsR0FDORkV3xltmIl9f+OzxrLhM34ja4G
vII1uxSp/BzeV5X4RfYy8IeSIbkCOGqfDyTf4ylOB4GLnt/kYvHxDYfQizOTF0fh
1qnYqmeXvFSsxtiRzdq1exvB41wKPgd+LemQTsB85wyvCDZHVlUtz4W3pH0/cyuS
dGcoRGJUJEtvzmjm6lR39P3mnKkp+o/c54lDbVaA+3Coc8iotexDE1FDXdurIpye
bM09icNeQg0EFbEUjRaw5gCOpaHJJLJ6lZlaBbhN/VZGudpUIralRG1/0ZTFyPpI
qEFHBJJPmhqKRe93Rvd2LLYSpuebP5bq8Kq8F3ggyEfP43bEj00HysPFyN9d1O+H
kzU4Qkynz65lQWwAC6cDMNLdxH3SW7JEF4e1iM5ITYhHDpddouI3q42YguylgURy
d9IhOviPjEpWQAVh5u68o3GObs1na8hlEPf3Q7qXxt8BakX17zruTGt+Dw5dQtmG
CWFf32AxAMwXc9+pnBVHQR6v733dbI9kpcZd6+F7p/Zlf1m6bWFo557/U/SuBUx7
LVyjVbtTk+V9x/kgHyxNqRCDInkIBK6rHq55epZsSoBII1Fb/OkPoaIIxTyrBYnA
xElkgSvHGyT1TqpccRXfdskXAdKka0lKWqOM+29H8EOV0lB+l2RF5bULXSuh9vl4
DqEQqjHCZ0XNmj0TLwNscQHUiupZXk6hbVkVEDVfEBLSrP+hjEyN2oO5YYWGaYIB
rU8+chWpvUrvYgue+k09dgxXFNJTpuAC26xclk0I1MizMra25EP89bxJXAKPfnqT
pFDU2xpKQt37z+7GloDzZAHgpp1+73f3wx2H71IqwBXq0G9bBYV+PISfj/C40oZh
Epam6SEmCfdno4sXb61ivqEZxRPL5pLAxZ+Vjbm5YEkAztugPi2GfXbvazpq/BDY
8Hbri8m7LM0fJtGphc3h1+snW6zLQABorlYcQQSn3MGN/QPUGNQPiCdvp46qqgVl
Wnwlz5OW8hzOMK5dunQzt38y/bDYrsASWJj/1ZMdOf4u3EqnVzHyuxDxvlNtxuim
ToOzIcviZ4KgEF8lOxXlNQiTEXQmbMCYZi0zv/MX+mo1cI8nvXyGfzPm80JEHPGF
nLDCqDPXowbBYjJyVYdERyLT1HK8jGS5on1gADc4SfkCBWN6b2K9obVRaf2R+n9f
5uwQT4DoJVDzsahaTQcMKIC3YTxKPwUueVMv6Xfhob9RBVluq4psXKsAsf8jXpzZ
FTGcnXGjVvXBtozu0YHiASXW2iTyUxbv/+wPQmunixekUorVQxN19fROZRtFIdCM
Lqjq2WJ0xTUset30y3n5n2+9v5AyHre1bXC7LBzA5anc+bETj8gsRXw+SB1v670j
HU3h1I7KZSYCDxAcLJ5hBgxDet2SZuua2Zd8I/cjR8bjxfwP8NsxQ3rVzNSE2Gl6
jPdAJEXR1zYFHM10ICZocO6bfSLu5kzC9d9r8qFj9OlHGgKD2iUfQktV65/f9sjr
Plt6JfAj+qsd1AK0YiljpArmE3Qx4VhRAwDn+axgB8u9otxZxgqtQhvPLCWgw8M7
g07KxdCMODgMVOsPDepraneItAtgoV7Otwt46kjYJT23/ZigCCWffxvL0uf8GR3e
LNWT/LI5F8z2FoU1vlsKFbXbfEC3pCgg51+agj8QBeIJL/H/4GwNQmy0iQPDcnRI
Ml1jL6hPXKudpLq+eLLaCYG7WmMY3wjTeISFIbU/gMFDVcZAFohloZ/HF50uvdQl
Y144id+IhAqed2AigoW1L8BQKyuPh22uXxxG/MNQSNtRpg/OD/wFX9ov0xDNeB+9
Ho36t0a/OUzhBa+/1oCUCpCPq72g2bIW/4acxLzJqZwE2UJiNc/tR0ICtGQIeujr
IZ8jNkb1GyUxpN05ianSiFTccMJEIaKJ8VJzv9hT3vGFyHreMQBnS5ARR7dlVW/K
dgBRXLhTNTCVOBOqUDouh1S4PO1uLmOlYk/5jaquknHPFFKTZ6RClvJ4tAoaERt0
dbkTrAtn6kmQAIvl9T1jxR8QZmhoGSSdIYGccv1NDludgNgITsyacZdFNeHfnSGP
d8ea5Dw2tcdRXoJ2bVcUDhi/WL9MN3C0YrNqzwT579MQqchquv7m1PiZ7JmMaiOO
kpcyBeTb4sPVNNOOSiYP6TTQn3RWzwvYw50gZolGYz8BKDJNUwip0b9ffrRB+fSu
YOpiHx4D7gEtLN5HIPC0n5UV6/ym9IEa9mQgNhrrgAkjoPQgoyYgBgxDvSnpyWDJ
E7hz67IdiaP7m4bIci8d47HFjNIrtHGLh1Lo0k6BQono8a6QM1Bg2CtDX6yHREs5
s7fVjGT4bBcCuc3j0Qb3h5L1P9xifXWgYH9xhFOAU6lZK2FkzPVfhE7rK06Fupnp
F2N+PlNGpcg2xBpIKjRIwaPvVP/R9YjCOJhCznM1hHgIApoYr6zx1FKKu8cFT38/
45MJCkBaKe/wP7GbtX657OuxJQr6ho7EuMm8tkCLqlgM/05UK6W1SEcsKlQ65fEN
jfZl2fNJ8ggEGLB9mjYNBwP6b7cpIumDorLtZ9uT6MbyMCsfZ7xArsfD3Oke06qv
Kc0bcq37rusxrtRGFbXYyJJNpPcfJzJ4H1ZvylL8aSWHpMdPMoUAkTfmJcmbnc2F
skjPcnQc2iRTT0zJlS5P5Nt5GWxOTpWCx12mMa2LXr1tcs6tMIhCRH2UFO/CG69U
JqZsEWDUdofIrZMKK1tbRy9kYAAezHMnNdnrS2o++pWokDBEpNrnAIpzTmddpECU
eMEzBISBDpIC34dPd2S2lkvoAdMNQIlssimTcxPrHmRg1+o8FGj82+TMtiXrIoNu
PwQ8dwZRI5LOX/g6nQBhi45pN4zE+T+mLwLR5kvdOCPDrfpT5jBMQts/TtQNfkRs
hnhT7ha9aR4og4tHtWcqfFxmltZe/6kU9RERDE1lScYkg1jQclhkSGNkpPd8nrqB
h9g1ljR0Z+p6qIaNTuz4aVXI0Ef7//6kl1wh3T4kK9I2ysbGeWllxTJHsbfa0+qX
QEr92eJmZEgwmrXgVB3pDTPSbMvwPGBE9rtlsQrPosHCOLw9P9ZQ1hBMRI5arHsm
TmaVYw3KYb1DIJuS0GaPlQciYlVR5rQs7G2/PbADgffn5CphkB5W/QClhX5TnuSc
KQ9RmSF4NotSgFSY3Z1QPJ3CVkBxvbjfSbBqfhAFZU8WX+awByN8cHYaqas904wi
xiXJ6eINcP9Gj/LvcVfJItPcYRXGcAhbI2ApTPFUeE4KMRZ6Q9+nWDKSWxBV89c/
CGlGrID6oeAdfQMI9X7/TfGoAeNAZMmM7eKxSvSCwPEmUstnAE4Tw3CzGB1tO84D
kCz4i8tAgjol6nh4ZMQ37CFtmfyMzkxSP577xgeiSFSoemuRDERbeV+a6vbWf3nz
NRpO6CQr8/r610cPz/IQG0KxLi5se/gv0jyKJxXXlRteEHBkpsSz9lptI8yg8med
5DStEqnYnn2pYsG59msiv1pgEe8rXvK8OlX4mmWUHHWr+H7r4PBckNudO3P709nG
ZyUxsOjPMURUNxxGkYMXwpv/K/pE4x/zd6VcY3Wp8enhNiA8GZJJVVThvghIR9wv
IGAQalQANP2vQoNRlQcOw9UKlTyzEsEdTr2rO9IGjYpxe+qQbd9/ocbkERr5ssyk
aMZxhntQY/GWj5qrFmM4HdYDS3TLPy7Wpxu1ZdS/CdInzjzAnLSc0Hoy9oeTdkpe
NexhF1b9w8mAS9SVihq5WoVBKgHqmartMDxIL8itc6dTdNo8iAwid7/eS3YMpig+
lNbWEo7g2hEkpAD98M847SG3+MeAuOoaXKL70L6hH9R+m+CfwHIonDf0E44RKY4f
ji7t9ntjTKInUewGlcktyG6OwHPiYhzMckRzeDbB2NTawcDxUW8WD1w1TkO85j1w
wjBxQaM56cKGqnVup8dyr2C6TyIYxi+zEd6tBtTYhNpGhp3pwjxESKARXspEpTk+
MaUQsescbctZnE9hiW0VmZ1BANPVfh3maeUPy7dFKIyC0gWlyjXpVccI40PtGJIn
MVHpx+HfvxWopX9+8V6l8QWfW8XD1Yunmf5jOVjX3hPbTOL6JMJLYNKtYBlplSkL
/UmCG6DUYRm0um66HOBzOihTxG+SsTdDS+z5hOV8G7q2aC1tFgDQma/DwmL5tMxW
o5mINEciY8FwT8LeA36Bh8ATaWRo6ZFLqH3lNKl2IjuLp6/p9bIgXMYSn4BBqb5y
Fo364kQUKikgNU6Frk01pt2c3ZFbMeEWEmnLgR5oePi6eoCoDXZnferNir5F553e
RN+M74YUpYifoz4RYznj7vQROqGcqcYS8YZf2ZZlHUEimvLoK0HmRsJ4Cn1oRFr4
+MY6lYnFJ1fg19QHOGlN171TgJ5gOst++GaWS7LS517sq+tladeHmXY6z+//lW3l
8FsN6kAgfPvdQHuxc2fTU2BHmr6WXhaVD5aqPwN7QxMPtcCiaPyubz+YJ/tZs6tl
FbfMAIY4A/b8HKrf6ANnVBe8HQ64lN+Hw+ZK33UP4g0LwVTbkwMq/lLH/ADy5ylQ
SRZB6eLejH3Pp6qlr0QXV6bcqMK2cfP5cP47UCUB9dVffZPCKOXkyQ8o/y4gUlmZ
l4ym/mHlWaXZDqOkJLikeTZ+97hHN5KgWxZcqEaaVl1GJAa0oPXsISoB3TahKVFv
J+TeD1KFHTghmih/PblflLdtZSjptTS2JyTmPBv9rX3ZnDRTahYnbqpJLVi8NgfM
PWY72ahc2JwJmg3HUeFMipOiMiWiNmBFAEVc384O3+KE0CQ2yPuYFvhjKK8scopp
pUVAe1e3f4Lb1dCUSu6E9i3qdExR1qAFTeu9szd+UOz0BK1H1phcljkiMjr6rEdA
KLhuFhWtKafCa2ahlQcNblITOoNtsr0o8cwDld+gWVeLFXEWV9ghRjYCefiuNioQ
8+Wb/+4JaE3of+cPZUy2VPSQNUerHlvwT+hQ9xDubVZwaXdMKsFxd9KB7LUiXG77
M5PpWXtY50b1YI7nNXQoh+x1H6Eec5DKtKeJqQKzLQ0zAc/to3++4mJ6lxqobigW
oMy7BdpcqypKIDNd/VtTjFuK7kLBAwQjVshaD0OUe9OsijOrGqjxt23t+JwfOeGw
wnXJ/gH+0Iw0z/6UTjUKJdzCLPkQ2mo4HaHhBfPICD7jYzXqCSzPz0Oo2ue7r1Xj
we9rrB9CURWsMxYhSsx+30R2CVXAOpn6/1UKEnW1vEkGI1iXqQlfF8jQZH8o6F3J
m84ZZ82YtxpW/4VEY2gfU1wJL4/B7iTsCaB+TuFGjhLmX3QhICAraYGvFg1C5fcT
BwL93+WRrTe7Q5oiwjvq+yz67Tg2Cn/hdJ2RaQdBFrgYt4Ft7Au+h2wq75zeS4xF
9cP+HmetRANtOEOLr/KJpgTX4pE9uULIYMxQBy+S7Dq41amg7WGd4emNNxhiN31f
QIoh3waSr0TnOpqC5kFxQhEmltMw1EI9rSJ+mcpbUPy8x140sI+rQHxgkOw8WEa6
f5vrN4DTzWw+JszMWXxDzYsQrsF9zR63LEXES0bc21XOiWG1Tyr8qvjS1Q6jEa22
K4nzABJ7eBXrP+N8EfIazs6lds71/bK+57q/oqlvmpDZAU9/pXc05+AfN8XzcVnG
HKBSl0JvZKOINNeqIccSZcB46x+UA/BJf4JXc8zjcqLVczvN3v/3Fm8QMXFqqA3k
PpTWNLoVoycI1g09hjqflRAjhH2ymd2/yea8olbhyH/o9RemRat4JZ6nTXfPgBxo
ypc/hqSwmZq/jtIcF0RZJvW0G7GV8sTKZllQu8TiBISS/NenLe+bfyEVZTqoC+Qg
ejhK4n3JWe4BlHMrV5Wqh8VQGyzC8rwHxvNF1bp86VhQrg9xV63PO3rpADw6kgM3
bnv8QrOGGwEforlqw/NfL1xFGayEUy/Z4u6tJXBICzEmSAaEN/1qtkO5FQcGgeMp
uqEwc38VT/OnAY/SJ1Ap6CTAmfpv6fClnkS+IdDytOK4icb6uUg9//q0qXrF4TNj
CMuOMk99Q1OOS8rinBEVemooqggJQPGzSU+DZHEMD6kxu2aoaPYYCDYNj0tgkLQY
EQPotIuQnENBC6TatfNKZ+40S+UV/Sq+aVOhWJI8XldwBVuRgxJRoXDRkdog+IBW
tb/I7AZ7jTHhyvkHQrrRgmV0BMb8VrvhtRneRcwzhd2Udc1mrxSzpshx6eKCpfjd
pzGw/1fgt92g5do8vI5wW+BjGNl2GKuiPrQpvRXpRLDr7AZFGFOEL5tZaWwFIAsx
cbT7kUy8Rj9p6nZkjIS24VAQEZ5yRP5e3sQHZng65/z+pLCxlM2rIRXQOl2wPrvg
nZ42tMwXjvkeCur5sdv0wIjl8mGIT5LZCZBJuyR4BN+Y2lu8t4frasptUBDznbID
/9aTXvJxaHhDE8LRqdQMFEeZVvFZnwkRuVggY/yPkq82wBbmErWpIPKJBpG84PFU
IM9un6HX4I8UKhTIiceYQHBU8XPHG30RnIqdTT6BtMRLrnyipugUFxNhuoOWoYqj
22VDUJCEzd+4RqFczeH4w7jF6liV1bY123pK4JJR92FoKCXkmGYFUHCpXZuikK6F
rUE724lBJDfxlxniyaw9Wp37wPnAkhLJiLMP8EYvgHd7qbi6kqaddI7uMy35H6G2
JvG+uVXcdaYw3q64B+i1wpJErJWjl/I4SC4ol8EpAEsYzdK4ZFesOOKMTG66ZOo7
HnUvyse9JO7vDQFA+P+RaNQ/WXUafeZr0lG4F2vkSid1DxGL85tetX1gAIqYaWmR
bM9RqagJwPp54kda/trb7cJmGjSrTiy5KEoYOMtkgo5jtxUq+ge29zbTgAuXujOU
y7/gNwLbQfu21FFvEyj+XEVC3+H/luU9s7b1lw7mt4a/QCAUBRCkN5SKhHTXUK7v
4ex5Jpq2mH6d5cTvywfuVigqbqgdYgBjrlE5IMaR3UiIlHZ1wwNq8WX1oR41OXT2
x4bugyIZqlTvKdtWpLHccXYQI7QqSCnfWeI/FJ8a7XYXGV9NEp75sZOtcJ7f4MQk
kWY7X5tn6GKlZBT6CXZGIG9dVx+3tfUrT08c9lEaFMqfb8F7U8SyQTAH4wUFvewu
7hYujh2/Gi1D6F2TjqhNyTNxfzQHP8d/onm2LSHal6WFQr+PPU+Wec8D1DCtVSY8
thuDtbt3w8BhQjRGcShlY6CytDbvftY9JOAgkQHTUDkfJamsPKd/ILL7P//UlnIa
WXiaN9fHDUswy0/YlaStFqicJKMhvTVBA0rSmfHV79MeYRx7RXxpvlgbnkfRjtsL
8XPfAtqiJtJDfgC+kZAGt4wVAjJjq4wViAJheTapQcbMHMVXf0NDtQ4XE4fCQ1S8
u6AfEHrLuiylmmNb/XvwywqapIg80K0XUfrGCdxburo5LUvAquXVh/ppZc1JUNqa
iqoS2ofLsFiHf2FrQUgv3LVD8V5P+mrIpy20T4y6DD7K8F3Jh/HtuMA47jm2/Buy
qqShr+XTQV4FmDTmAmah5BczUBuUtLjhEyvfYcfcn2Mmn2LBoQTBcm8YT+ofeqFl
W3Xj8QOLLhyn35/X28zK2bhWEERrGDBjKVlUA8ClbyaM0WsJF95gkxlqjaXF/kiW
Ad1YkkJCv7k5FqSDrEoeu+CRmCUabeYJSfwpZBOD5/DjvrGpQubeKMgeoOLbWjeQ
FrjvJw9rMishCYW3Ov5dsZDK05IqpUWbA6Kf0zrVtZTkRT2fs/7k+S0Xzn7t/Hq3
jtYk2gmWF0yEhRUToi9G0UkPxea0i7sn+xxsb/9c2/95oRq2NNR/UXv6zCsreKfA
JIC4rxY/0pql0/dgCSCCY/+G7eSF9p6Bp+qlwyrbOMVY0NL757XSta1S0LbHfRLf
yhAq8L+WLlm1xtwZAJMu7pT8HiilWyY7fVO8AQTi/ue26Em5TrOgUYPqRiI/Hc0W
LLGKgAm6APyrPF0OgyE+PIFTQUWDBvo1n37KM2XwsyH22nKNpqmCt93T67PRTGn/
k6TrS7o110T2PNF+FJGtMyfMAC4vf6ZWSlprGfh5slSy9g1scpYDEuwlya4gjBHa
27QozTDjBUjPLxUAxPnkNYFUfVREbYvrIXRfVUobqn+Z7wo7D7O0xOHCROPYJtkU
hnBL5drxGuM4TBM8INHVISkr/E3GJIwwFqPh6nYYi+Z1R0ltCdXjU8y276iF02rj
EBrky7L4YTwuORRK9cWzeDA0ftmw9PZ9BgpcOGazMQmeYJhO2g8xWWKmRpPr6foG
TXWyKNg1Bf6TrQ7/CKKSty8Fhg9mcMdu0QTFEELPHuR3w8CWeL2ECDH0H6fBgvQk
tYAPQmsPSMBUShhKaplgp6d8phWDtmpb6w8MjteGumFQ+WSmht6Jr1R5KA+Pzuhj
EiScLEnBtNcWnlAHdy+uvo7LEfxVOhGz5SNKgi7+IN5+8jgz1fcXPmyLYApgT5QY
Y0mwpYUUCpHkLCu+CiiVqHe7LeaBji05UJwxu9g2xSY77X2tCv2D8J9wBy+jSEHg
KGZyHy4hnnTl3Hr/7L7LB0GIuZtPMNWJVpjx/uBU3X7tBc11nn0ycsLLy0cFjoAV
GCK+iK/i0IAe7vBWGcnOqW5QwHsUA9IlXsfLGfInBrBLuJm7ToGTf8js6yMyKRyp
DOQVpOdpW+btM4wUZjrSRrEL7sI7uStXdeTHnmykxjto0KMBvxfkzSe9l0Sc3aad
iP+/BxYheDzju2mgE+HB6zfqNIR+K1Nlu2sg5vlOKoz0vf3ujAHXtXapAeM7FFzl
pZGMf2HLQmjYW60JNsVkqNhA2fRHM/QnflDVExyv6U3k1MQPwHMaF1lAP9lBzaiI
43b6MiMmlxXKVu6RISYb8yjiN8MnejRSmauRIz8/sAX0tY1jq54LrfeqpsaxpKxL
s7+PLIzqIQsE9L07HWli6T2qNWLgg+HvI7YvA+HMySn1G2DuVM24pgc40JIYsWgv
x6+PVjbxHqi1QAP7rqBgg6buHUSTAz2Eo8qXCxG8M5s94ESRWNJn/DhjP9y+yzHP
MPJopBE1vpWSwk6j1bG+cUDTLf6DylFZJxqWkp+1qb4bG5ded7nj3xuoQeSTQoEa
pQ/TpD253NwN1vKIKbDsFwcdLwv5eVkapGlEYRSkdBmjXr69OjYv+lIj+3Er9RTm
jXc7p8qYN/v4uVpBwGcXfHq+H4Wws6pffhAc9arx8yX5tiG9Ma7VvaVPV06SIhJe
8rDRt3XnAoCfQMU95XD/N/zLcEMw0esPo4DdNrVbFUpzwyGWrbCYh/EeL4UAQqcR
fSUxuL2dQ5/qMwiWLCqD0OydfjQiaz5/hky6KRq/mpvjY3+XzMVPM4Y8HG8z2UNh
F/Wt+4V/1uZql6e+l/OlTrxaza/rjJuCeUiJtWAYgzGuaz6v3I4vSZDhoD+Q79u+
NQ0hGieiJ4wbuYiXsI0SXX6ZuxYazHEvSsnvdUFwzBHP1phmpOpRKGYnmInMKjTo
43kkLg3lUmxlaw81JnwaJ71WZKkhwhsbcID8PAl1iArZWFqD23xoFk8JElqtMopA
VxT7EkY2KTt+vUq0lVxpCL6lu60gsnbAYv1pGtYYEK8XYMhiMJ41nFv386P+DC5h
n+bOaE3RiXzktOK4UA17J4Ws7Aem9cT+WH37/UgzO+bmYQdxuxgmPJqOc33b0VcP
iHnNrZwNLp+6ZylGsLsJXLG9xJoycgW3jaAbV27z3plCCtF8C8kw2bxBRmREy5j8
J/uSyAHthyB0ilHBLuRImXMRMUM4kmCVUn9CIrHKb7wg8oWvHCM8kaH58vdNsThx
So0O8xQStoCikt3vjkSF2B3vq+Ud451wOyBJMBrln4Sj7qoIhFn96zGkxFe1sr4C
GnkiB2hdz2NWHllFi0KtZlhGSnCfplEaILCic13UivzOq24eYTUbgkyEUmCKoXjU
uT8Jwr3YqiDyr3/bGDIjhPWzZtG8TinQiCY3Me9YrDiSFxoBNo3lxcBKdvVgQN3t
F+bNLP2pMBT8eIUZTwLNZmW4TexP/Ll4Ns/3Nhrjh0NKCF9lFf8V00b4W7qL7kDy
INI2jZym71+AGtNFWJcIC2NfaZb3jjryTqp91coFojBgLFXNy5P+ovByI9h4GDLu
bv1q6D+BR6Ms24zDe1mdovpPiBv0rXV2MMXkQRbNCJWQ3abNrkYrjVwqedAixEre
CjznpDsNzNlube0wQwQJ0Uf9uUrArVUM9DLXNJiz7WA16GXnLw3XSPNqKt3UNwEr
GBVtfQ4sLE42jXV9hcDggB6OapxLbP8fBKAbA0a5atera7js+paLYNF/EaxETH7v
o3DSXaPoqhpJc42ncnGYe5CRM6IQcDpJ6II6fDiy6tbJcgBDVj8VjQBl1R5NEpZe
oLNeCy5J1IYP3ScUV0qmTog8uEzjDDbbtr7RqbkRcFb1wHYP/PmGbCbGudDQA2Fw
xrtjhA3Gy7vNsvYEuSQouYq3YWHfYf/fTFvjOm3X4RIrFSwadcPjJupMFD9WUgUd
v9WlDxMgKf/Z4YDUKe4iuqpvqMqrK1XRtnjCQu2mHbz7zGmN0qgWiUekmW+tfD4N
LgwazuBEh9uLbl7sWOlUa1UQOndWCJUm8u9XHtwvZzMlWba9paA4GaTUtRuO91Fm
FETnisKVPnYnZeu9uUiqQojYzhkOqD90MVCV1bmVCd45klecyqPkEAnPoya5eJdq
YnKTYh0kbJqm251BZFAKsKC6eMFzSj5nxFUsYpI8aQ5Tel4kU1pb4OimodbXdGeS
tQJPc0PtBV4N6YwE/EivYq/Ho1TRcJzrTfxXWJapdVKtpB7VblHyQ8372szaUz59
lWu8Y+5kHl9/nATrudqPXBwv69/YsARBr6XE1pcmlHSbMnPFtQXzZWW0zw4sosj6
TY3knLBWkitpCliSb1buJB/jRTckNwZDro82osqLcFLXQsQtOe/LTmSlrM34fjyU
ni+Ez9T+xv0j+lNANLo4uu0uY345oVvQsmn/lmaiV3uSmjJjKzUkMtIJ3k7Kaygc
xoc3eXLjV0TwdoYCSx3tYtphMw6mkjs5whzEdPPpQyu8U/HXytaQvmi51MVvzKIk
NGhG73yj4OAj0D+obfm419p5AoN1RQyEO5+tYOzZmUziz8tgZZUJujPGyvqPExjR
CMRflLRveZtOqX+9eMt6D4zJbgcGOh3BBrclUPk1lb4xmI2ecURziuJjg/vp36Ay
RC7nH/m5g05sOzh4hu7VDK5xv48yiwiJnpQaIQxARIldfWaHIUWFmHSKJeRz8AV6
t5r2ndKd1jWRMB0PQm/sC/FZ8bTgQSn7r3CZSfzQkiI8LUbvW+llblKij2N+6Jro
eNs3oTCm1ePufF/OBdEKuAwiu+w6Rr15ysuFP5fJuvBltvuBmXus6L9EjDM29cAC
5KWCkQtQIcjtOf99T3sZa43+WTxopgqN+uKdmb79lH8f3EMUcSPZEajeOm8XrX1M
8BPw4T+jP9XEmVrL+ztravphFkKl0DC9Jd7qWQbayreWmuud8xZdYVvz65cLKg91
0M5zrk0S8uU7gf2/jJEXjUCZ2Ii8f8xOVjtx0xIWZB8e0yL1PiY3LeZG88Nt4B4J
p9NVfN8/qiKMJIkmLG2kW4Wvnb37oG/fUUF74wV0fkXYgIhykCO1lH3gEyMLdVqU
9z0Bh4MR3vB0I6hCWwt+sAj25ORna7KexYMfEH+y8e7YZT+DkuIATp/72I/UmAcY
e6NZqgwv8g3PtDDal7CX4Kch1GIR9Q0olUHq3/ikI94Fe4oznn1p1SIpIPYcOCE6
hCN8Ep3iLhBv0T9oWO4WvIGpxafnAhQlc/dX87O2PHwB/QvhoXtqsFDgIYrScmS4
6reh1N19IhQj5fkmNNFU4/BddcF05L6FeXZbiGsvPdsvAkIJvcxD9qXMTye4PFFx
G8E7EQiRUOTECao8qJhy8cX997IoOPJcwH96tvENeR5XvnATp89ri/7ynKvfMkLI
Yj/UpV3qVDqYIBuDv1Y+efD8TNB7LByFKIUMPESdWheTxrtg/gQOx43CU4sIM9tx
FQQogcxAmTqK3rLPDhCf6ZQho1dXgfNEBlXn89KFsBN7+IwpMXB6S4oY0eLdhqDA
cnOuPYlov3q9K2cacUQs1xmt0PyCuvoMMfWVhiT9Xe4+Dtmlq/114cTl0inrgjSl
r+GMKf9W5djZg4w/JhayIaIsuD2oY9x1420GZizij3ChaoRa7OH05J4Z4FupLBQF
xCYZYHSXoqa62flvI8dcw8YC52of/2OzUTz2oGvjUHa5vjKfwH7xPcpw/BvuzEOl
l50FAjmEC9LL4X0BwPbMed0lP2HXP6ezqrVKg/ML6S5S6dxsFE2WMiMa/7JcpGfF
VWhG+GSgDi/GmeDZKM4JKDOiJ+m5py4hjuO9sveYoxwMYDUvaE6iAryLQJZvCA0C
sZ+riNtxRPFT3efJbpPs7BvFOmT6bhk5uNkBEUV7A9QP4vG3YfTsXDsXF4Cl31eZ
0FfzM9NBQHpeCfp264xHfRx1xQEOXCLu3Y4QccRWpFUajpEUlWtJ72ISSPr77+aO
cm6+NTxtr8nlmOXfYsyMWbOKzafALC27ybaAzFCP64iLOVI76I0NKRkjXrXSAyeE
FsSRvZP3oletT2zmiEQbKxWsatQEQvjecWaxMcj5pibI7iULgs5x6lV0Hdby+rZO
EhCxK7PnLBG62K8aqEUAMYvWfmoY2peoLtM53VEgZdNgC5MCbnR5pqkD3eezTcrv
VGzyuAMmKTmfa3Dc8KRkoF9O63sA33t9dmibuvcU2rTe1AN1rSkdWuwyiXY4Seku
Bt7m5CRhCU5F/KgLIM2LYdrQFxmkHZ7nnS5o9GT+ZUfwu7VywrE5NWUr6Lms+zjR
Wl/QhIphUE2/LrRI7rfK7QPNDMXfVYEt523lgi6M4FYo3nyPnGD0aqgWKoGNzK68
mEq+w3ati+Er90+9Wcp3oQQbbwXKKUNmWJ3s6Lr7Mv96CSEX37LG415rxx/+MzLN
4KML1cwWYmb58MsKBK4YutfuSAiq88/lxIPaOSh30AJ6MjvnOk7/N0J9DjRxOTSx
e9utsK1SYu8Vwsl4FEa8IY1AXbZ4+jxeAtElokUW423ncLAiGgtPWrwxnxn4qD0T
qLNjUwQas930Gd7KIP0y100VgwKgCqg/2RPuRc40U35UGP+8HnJR2S/zHjITRpHt
4I24MjCfvuM0E5GGQTZ4z6vcUPn+8jf1ORUM+pQ98Cvc6dyfxBJUZaDJaP2ruv8W
HgFVJ0H/vLbVBj57V30GoZYne8G3xuWo7NVk0L5xLNTFSXr5xPCJ62IInUlzTnRI
rY2DS9AxiIRnQagqWQN0H9xhZPswWEvTcwEoOiJOE2cz0kN8oFhdGKiKe7oHROKP
WE6/8UVQE3qZWuJRP0zsBm7CO4aGr9wR4i53EhLEKoj1tiX565bgLKlVGY3a2pRi
RsmYRvOY/T/FdN4t4z36fDUEivb61rwn2bOFnizPY2ww1npTTHFQycWIlV4d+VcZ
y8JLdJJ6uePGMtYXD32USwWneyswk9jzG9nS66W/VHzMS4fimW9XMKRFMdfmZjVQ
ZQVI0f7hLrBOtHxAi2t53cYcdCPm3JLvgCRC4gtgEQ2G9l55sGuK4PuY6sTQJKIP
j8122USGPa5CrVSsk0WyWHbhDuvNgonBAPz5hWcKTQIEsp3lBxexdZJTCCcfEB5d
sSnPoJ2tSRhoNToVKngZDbDtQZW8wW6qWT1OxWSWa9JUTKKg2p0pGUugVlYL8eCY
wieDjK9XbK3uZ8FXisa6fzV/yxvtr0w0K6+C0zLjGlOPS/htMa8l/6DnvHRQkshs
rE9ugJ7kaeYALxYtqxyMNsbsCefNHi3RhKgUVqxEuIYGFqBJN2Fh9kXHJYpX/TgQ
sNDhOEvoxuuhKTyXl09yEzM3Ba7K/mbXlzyxtvoBioGVtzoLwsLZVDEkTHOw1Jnu
lzWQnRqIbM7TSa21lhYvEd5gv3vLDiHAb1YVihNCesVTT+e1svEK1Oa36NiDVfP+
dvGcuAnsm3WOSCQ5wHzUdWmugBOGj1H57PyRctcqxKUmxnj88ZmvMBNryTr3JZYS
2sAETlcR5mI89t6jvr0aro/LUPoFyylnfJATeuil/RS5dmktyqqgVwez7cSlGqvv
SiWkaDHeE2qlxLl6v16LF+1gRuM7YMhNtIeUUnMIJIM3gxXEnkCIbzCPd682sKCQ
vMSG0V701MgXvgk56R7/qyj3zx/Tj5IJJQlF36YU4odVrHMqCtNz4/mYpR+QE4yp
otE7Mu0GS9JsI3KNNjmbGnMPuAzq1grMyRsS2mb6QNtrCa3Toy0oSDzB1sAEYhFs
v5KbPbtwozVj627eJdrdpcxULPtLVxLKlwckvlD9n5rvcUTzSt9jQai1ZhfCJwGp
8JbgHrdrRJVZ2wF0fW2H4gp+E4wq+b8hKUkYMBy2GZkZzq2kcgbcYBFplIS1W7zc
SH8w7lMfI0qkQaTxoKBi3MapufWCzAIOjPaPxiCiby2TkVwbUB68v8ymWLVFjfli
`protect END_PROTECTED
