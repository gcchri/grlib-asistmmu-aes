`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ItP7DHLvyCAMVzAxMnSNxsP4CDeHe3Her+AvJ5A29fDZE067i0KGgahw/qr29DyR
o6pnZvj6fc8YtdTIe9f62ZN48m5bJivC5G/icUQVcRlnwF00V2O68Ha/wDOsmaiX
Z2EXDNPP2b97Ivwfb5hqw+reNa/dPGyZkztkRxgVU+SXz7b+bXZumO9eAgAo0vA/
4+wegTAxMKacHkn3qMLM51JDz3WeVEDmcL5FUbpy165l8CBQryAKu5BzxgCzOvCo
jAK22WMxh9VtABUmbwQantu7Fuis8nC9Jn0zXLlyRm/+txGPaMBbooYrNkki09vg
GT6jsaGgIQiFfRg2ucOd6Ry1/V5m4hCFDQjcB31MF90O02J0pY5MCEX8WXDLhx1Y
OgkaQHn1ArrZM8JNIj7zMg==
`protect END_PROTECTED
