`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sNRjjSSmNn17AqU7mejg7otR3qNifhndo3ULOp0DKz7+qxhLp0cG4Rgaw6mOaka7
cijwOoa7Q7sivGOn8PO55WtQXaEe81xB30lfDw1V5KTlJMu8Nm4A0uiuZ7rLpDZB
lgSyEFrSnqfhAOYDBFWyU6pPrWzRAxWoBTFrE1woL130LwG09u4FOFjmmCXtYAsP
UeNbmirYCNBSt3lTcnzwguMI2bDRRGSBXAcvJ536e+6+XQbtyMwk1SruaiGJprF4
O+0YWQ+hs2HGTwjoUhV+GQ1edsSJXmikhKY+kR07o2Vno2QFyE/De8H+mzvnYWud
/gkYZP/ksoSRmEllUbd7kXHAMvBpKWw+YgNiudAfJnYWEPVYzJu5cqW2pddnOLC8
tBGPPv4/CU20ZrJzoqcCRV5A5yKyqUBaBw0SiRP5KUSRqHO85NFRhWqCR7epMmKB
UbWf4q1QdY0n4TZKR5z9MwfJ8YykcRZOIgjK/Q3JIlelNeRIsxsfrorvyE0xHalV
m7DJq2IYprwAds/FjJFZmn7MhEifjaUVr8APhrHZY8vV6geYu9Fr9pbrjUf1elgi
uqhT9s1ZpAJMwQl1/zFz5YC/fsIVRJsZ/GjHBeK0lEHiM6hR/KXQ5XHHIi7e1vab
ojlTyEXgtmFG1uY1qV90MQ4f8rEVPOoqnbUKKtR/p0t6joofTBU7EcXJVo2sdRrS
DDwBtE58MQLEvr0L3zw4SapVdvg6+e7hFnMiDT8o5P2a2JktQj29il0T+gYZ+6Na
Ibp9EBpj5z9/nh2TCY23To4PS9nZ8CNexdP5zjF9kc/a2hYMlTW5uba+/I7iR1/e
Mkl61Z2INGE4R0vjZlHEBa0qH6FWpu0/Nqu3yqgJpNguMPpYLkK4FY1R0NvB6DKj
GloKao9S/Zbbks75zQLwFna28oo2Bu0pgFZDSm9iAs85RqQ4nHL+4w6wSist/5OJ
bHOqO/1GEHuW2ORJ10TXqg9A8QBPSVyvjJOdrpfEZ9renxOpqXC3vz4D34yUsxIh
Uuvab9fSp+IyFliQIMf3HfJk4krIFhfUmZWArK5fovCZhLN6E9GoQwC00QJtyO+8
bucjBkJvSDh0ydISEhKwfWAcFhq0Y7BExCrxPIR2hJ1pyu3L2UWjKYDGbPKwL2a3
WwcIjPqe0n+RGXZeS7z+yZpbqem3gpVsLAGiV+ZpwVmFyCdsbByxSX8a/jEPKgBx
ftZFa93xIhqNxqsdQaVUMw5WoG5cji3ORsaxSe+4ekWovLGsfJznL2pBfT+kLhkS
MSiPiAY07lHFi6Z6qM8uYwWk4O4nXR6TYQnaS8cqQlbnOiBt5zgDHFN8C0Aj2l3s
fVxF6MgsjPYrfnjUmOsv3v34CoVNIVfYTfUPpWqFipKYCrSAQgqDHK6tXCqfZlyD
r4UfxtdYTDtohzZdp8/Wa2437Fe5jVbeOl6I+4Sg3uXHAdWMZUYYpzko/Hruaj81
me7rPXPL2b9jCLYpvTOdLe4+DBYZZoUm9AnVbQwhyEApNXlVzcypoNhigORq0wmH
tPyv1DdlHcSu39iNBXosFW2HeezjTHezfgEcbBGw/jyqLOib3uRvY8afn0aTIl4p
3WZN0LLttOz2BxbxOTbku6y5T3S1zisDSEoPuJxmSMUP2SgbqQDcWxagnS62ioES
7GrABWl+k0nII7UBtjYgfayRTkBj6QO6nnMhXPb5nYgYnKj0CdHY4YqIQ7y4kedm
63CuzC98IreetToAl0FxgPElCztmHiBRLb3uGuxtaR8=
`protect END_PROTECTED
