`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n8uJPvHOiDsrTGYSiCr3INmyU6NVbnP5ovCOm/tFjl1NL242f1XoSf5T4+bK3dKm
L9ChBctGFd29Qt0CO7YOqUN1lKcE5MkhNp+M+Geij8PwuwMvyBgSue7YcDWfIjoZ
a2UxI6ZYzQ1mwPEpcRX8MUYdftEa+BVrEKWIY1c/TbUHUWuZC3bhGy4PlUpJvsSl
Vu3c4m3HHFsa8r/30RDhP1ra+xD/BuaiVwQCEy/6jsfKAVpfuq8kx2ruzTFYo3iz
nQkD8bNghWz4tJutV8jqGC9JC7yCLa92cYCljppeHf4BpKwqlbeYj49dBJ4IiTXL
AWiNCZbn4CAk+BPChgRgxWOaXYDqyPjc1rDrbytiUZwjqlzKVNsWA5EUOwdLvR2H
8GyNP9vEnpF/pLWRs8TmqA==
`protect END_PROTECTED
