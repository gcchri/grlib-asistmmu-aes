`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IgSTnWqGXxmcISmtT9RCVIT+RlP1KSyQmwjj2AfhwSAYkyLDRHJX1XqaI/ZkuzUz
ccIlxags9vkpPgbCMiEboct9fa4a0Sdiah3+4qX3FRNOMLit64rEd7Bfnr1HqoH6
k43v6TCv8HAHgOdNU/C/X2pgN0tVfSi9Sw9DZ9w7DFSK5gaKz9TC9ZPpzL+OCi4r
rGU9OXpEGYj7+lTiUzLcQ01uoR/5jqHfuRFzKHIqQzhUAcS4lV66mNwGkbqy8tQg
udUC4GFmHnPRsi7nMrWynZXIQZfi75Moewpu0/Vxl5/vn12husVISucMXkUVqF0Z
E8FuJNWgvuIBZdt/jIwP0VUtE6rGJXyujXDUfspmbXQzZGxSAAKoMWhRrQToHV4f
hquMVzIrfmWxVgLFL+RFsXWK/hKGGm8eacu/JzvIX0l5q4uqoRG3AkV1MXhbrMBK
tTn62IO1b3E2Ito4PvP7IpmSrZ6AtVuCaB6w2MpZgHlPdCiH8kMu4mhD1oVTH2W2
YRSSGoruEpO4Ug/VMQl2fJeAkqMFKru6NPkVUMNXdrRqjDI+5RENAFE+D/AH2hk/
GKrmVSqVjfc/coEwOe+LWPCofdYGMfasdDfBCzRprs7K/m2B4mxNV6liLKCtITm0
gihke733P+sOi8a3oTGUOg+ZGNMhjZyqkcVd+IPqgqYhDmpsOYhtGuXRSpNjXCmR
i8TCIFYcNjpXu03xErCF5FS8Nil380ZRrDH8Q/+PUHbMPHmcPBocZmfL/eEJ96+2
2VD9c3mlOQw+yU2Yqfd/vOWfDbhhrfgZ8/yXQIGLdKr5W3zz5tnTyLqpGmPajJ9Y
avg+vpH5T6zd3gMqbvwcIPWsvKyDQpx6eUdC2clQh90MTAx/gpEcKC8L9EDPxDKS
cJRX8AH4+nzcwO5P0oeN4KA7wn14IR8CYLaGA4ac65bGwGy7j7jGAf5bIBuJEEom
n1/6ehi0dT7A6vjkK26VPJdnSpNvqwoJRW220TCOGtQ=
`protect END_PROTECTED
