`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GqMlEQKrvc5kLQH4tVI4pHBndtyOD8k2dD9IhrI5JP8SxyWdv4sblLGBv9jMCyU5
U5RaDLGrfc0741y3LKaCBfKtzaJA6l4U9SfqXtBO4F6g/B2xNY3YcqS09b/IUuTP
ujlRd2ReVK7JL8p3n7BN/MPwfvCQubeWvbFhSRAbFRv1tMtf97jQVDz9P1kGu1V1
9Ci8tXx/8fbRyAkHfpNC8ADcz76dqI47sbtwErxUoj9XJCsYrQnj+4I4q8oBhMBg
ooNc3CMJCCHyiQAAqUGzhMXNwvOK/heWOCwtn+Q+xzT77y6JUguYHibKva63pyXF
3PS/4ha696vjg+zHF+lR2g==
`protect END_PROTECTED
