`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k7Do2SayVPx5NQ46WTik/viFp6QG2x2f+o3ovRHE0tUJaOw7simxoSM3NcdsNTEC
GYV/Z3hzUsBQ9Kn4G7b4QfYMDk5bO4tbOg769wHAschP0vIweFdJ5wiGdcUXPZVD
5I0gtDnEBoOuADCDuKZIOq5bCmyfXVG9YG5h4/w0CAD+VdmCDxdBSXUtGzrrnN7x
xjK8K4B8exomWL1TfTQKgud6do0KmhUIlRd5/vhf0SIFUo4X8R6AYRkU3qZdYnvS
UcfO8jAOebBPwnRsPcI+5xysjbW2ZhMA2K3jbrXluTYcQW+Y+nwT8MOQDu2LppDs
3y+8XnPLiZ2LO+K/H2v1PEbj3sUSucLAlKuKWyBrmXowQqCofdXyvm9yLfK/7jCb
/hTZlxYAzHch4K9Ih8RMgOZXp/XU05IRi0HXSRXwq63HEhx2EYddDi6Eo+Tt3Jqj
Tu8ExfutOXAykDW8Obof89QmlTlD7vrshenk41IrUU+XlYgRnWdL8e6pc/QKzInP
GysE0yzrC9eXl7HnxBYwuwVbfQ+9gLvHGsVC+86yCNNdT8xmBy4ZB0JDeaDPsYzA
3OP1PZOyfAntUPzCMPne3aHK8E+32Qe04vPTD4RxL3A4PML4nfoV2WdIoU7f9Zcr
8LHiZ8267fT9nLBCOukpAYNOWtZ6Y0L2XsLFvUs7sjlxYFUOCyONB9LOJMMMGQCZ
u7XgaWsaySUl2tDXQY8yYz6kDvnj1u+P5csOx5SOrhIIll0U72b9bYHrTGzcle8i
ACVVXsu8dwzbbDLbw+eu8CGEr5btodORixZoe2Ux8It5DwINoqbG0gjA8csremnQ
rS6ztbyI83zMM3flXWkTsMalb/8nrZHkHQDDhJfFftI8HcqJ+QStoy+QbKgtxOxk
TB4Hch6nF1lNPEi2N2g7in65mYI0Y//FI0I1Bs2/iWFcC6Q5YQvrpCjRWUQPKEcv
0gqjxObYbAIgO66bMjhcoHiUFNbMR3Sk8V/v4USAgU2MmHrE7e2I0o40R6e5mDqi
zdMTlyn38d9e3Fc/ZNAlP4ut2ChU/OBLqf0o138oCd+Jof7hmGFHAq8q1OQBRgvJ
SeDzSvtWHmxxpgR0aGBkrKjjN8/9eNmFKISFO3gWu2Bk9yMVIYjrAqKXIxgBbDV9
Xb41zbR54lbmFLe/iSsoMHBM3w5a2xhPAfUuXYoIQvLPS7M05+HFmHmc+lb/cCgd
GWDQiaDCazJjuVGnO4BifLSiQJCJdO130Zn79J9JFLqoEuEuauXh3lqwJrIrCdqn
TShYGHSF6xhycfJhgJgBkn3ZWjbz8LIx+PRkF85CK7jaGij30rexJM9WCS5spg24
wYWTBpk9g/JH9ciqYe3zzocQpcV7rB8TnDpesb87L2oXNeJ+fN9Nn9P5ujlwJef0
qAuvqN6wQa0usA87QYJXvHoQ/bWgoQRTLh/7TBAj4GE=
`protect END_PROTECTED
