`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dkbS6tZWaR3a//aloaLePTR3n4vKAkCaPgpMyewKCdLeD1VxAIonXG34cZ0Cjgip
ttHHAb8c3K9HDY7Qy8S7C3YNHh7H3+HnOSskqP44kw8s+QZ8hU7zLi3dV0pQYgfA
8WMgpTt92BauOxmAMDt81iNMu6MIA6SqF9SLAp+qnlxmUUYvKxv29TNhQILzFS83
MelDfY64Y2Tdh1tkrDRN5yF132ieQuF9+YarJnkal5sUOoBsMmxDvE8ULNumxH5H
7g14dP0Iskdzq9XEezIHbofIDZfJaQZN3OLBZS/GpBy+ekBH7eIMGy90g/AA1dE7
dmkRCXxKNG6xp6/cI/PWwDcKEqtOXLFfR2Su079gQ+f3hdB1XpWHd2vPk7Kfj1xr
LtspGYNlMsd0hGC1O7DLc7Nk+S2HacOIGgv654etA6Wjpcv04jhLOenxK1G870x1
`protect END_PROTECTED
