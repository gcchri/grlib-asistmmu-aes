`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GXbRIY2myFpDA9uTvv4UkL3Mdjpoex7MjNB7ACcw89rTmvg28wfHwJ0tXYqzV+97
IOJTlTCjw7Cm+BuKa1bWrvPLM+oGfnWM1n222tLgNJMBSklMDKS2Yeeb7S03S7Bu
synmZmy9hswIhXIo/clYFTvV+tq51BPh2W88NuJWLItb0IYXppYLEErCIBMGUGsb
OT3VqnZTJT+4oKpPGIIv5Wjsn+zrrRfXuzZP26SASRwmh0oAIA235B9oTc71BsPt
tkFIKVxkd8DNoEn8brApxEABXHc+OvWtmGUUfvLwpluEKVfcuT8xXDMuFm0X0vy/
8q7qiGtBMayhU694BKJNj39c3bX3jBt736XJ6Re5UD7L/Vb0ERFptzCKE/q8IzkC
eeijJzNx6pFI012IiVYFwSpNhryqqOaTzgK45jRwuKp7mkRlSFALDyUzL4m9diBv
KCXZYnI7sRczs9ecMnJEk8VlDAVyvq/urMxGC80mQvU=
`protect END_PROTECTED
