`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qbeTOJOJMOheUV1u4KlUwtXEro8C64dqYS6zxjpksLjhhraj4btYPZQuhTsimCLe
ftAlnQNj/vxayh654IWxUxxZLzXFN3jqPGJDoMku0xJy8OS2HrKUETJqTS/nrqWt
69pEMCX5jKhy5UzVRHFyK8rg4sbmdU1xdv2hZ5XBexmvnPGNH3vxR9UFWFDbm6K0
uPN330jcVN4vEzLscgXCngeET6IS8MKh3F9D1RIP1Kv7uqi1ypt8UromKK9A3iUw
tLj8i+liqTwX2M5hGDCa4Qy2V3TNWoqiRs5+krrY303/uu+On+paHgFgiiF3QCDm
LCVBywQGepMTGmOWD2X4P8j9pmSk1BdBtoX99LkKSXE=
`protect END_PROTECTED
