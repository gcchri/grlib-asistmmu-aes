`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7m91CAaywt+CQczWxvYGUku8GmtG5RHv5G57n3FhA5jilxuqzsj8W7BNmfUIaR3z
f85aYttV5tPl+QmABr9lQRR9QJj+Q/ByKeWNPP4t60uybbBzf5RRZVCbTNuSMtKT
JEumzQjXpFS3cOgfpCA2gYUVpyIxvbqvMOXV5A/JXJNQO15fownNBvDhnbQf1Jlc
AKRVNRzQegOkte1AOvjcJ8dT9PXIycmRofWc3BtCj/YJ0qSXw/lHD/wu7Viro39r
1DI7ftOUM+wV4YpZI/yX8r9iuE6GNepgJ9aJeLY2WiX+7QZyoFoIou3daOE2FaiE
8P9wQgzIW/ZQUFpuGcp2rGYWEDuJXxoQ7/SIvUze5oGThsPQZAvGkc1s5LYnjQ46
o2gLH0ddRc1wevEdYBpf2Md/uopGRS3O5ATj0X4ZOuYF49QMJsYzY9Bk2GUcfKKd
+prjv10XL10K8p8/+vW2uQely+f5sBUfTt0RZHal0P2vh29iOy/563ZbWdZUkJi+
AiepZxmHBNiU9PP+1HmuDJfVxC/O9Ro+4zdq86z563BB3lHYT8CDTVE9Aopx+89F
P1Au/z9AqgC68Wqf/7aDbczS4EMx3Gn5meD3NIPj9gLr4Z/f5NdUVy0dkg0fy8ID
nnzxptlTSyYiEDamsA8XKL0tQqjNpQribtpF77jsgfJy7vn3rZFekEzkZFXpL8d5
hlWoND0mXRfqWjjLVjdRRAanRG73wRLX0elGlEJ56dq9a+ZVrO8X9JfcjvfhDU+c
Mm9yd2kNHCTUT/az3hq8UjjAGHI7xK4l9LwQzFlVrCJhGum6fELovaSjOIGtMutw
6ZMQBAwLKs8wVd3UpKEsJRo+dxqBjBKKEkRPpPe65NmDgpqpNTlJech68ry3VOTG
Gm99XyO3p0QDlXBjYBm3GTYcGUHcQo7wXWEjUyFVJb2i3T+3vPVDnrwMyFdRsmWD
`protect END_PROTECTED
