`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ly6iIhN9WE/ksv506IggHd+tiQgWx7XWY/CWGwp1DxHN4dnWPooX7VgatQKlGdA5
lqgBeuJaJN89hnco34wvBxaEz6bGHfe8FVEsy64nC3aPkp9l3Ay70t9xlv4ikZiC
M+y8ogvoqHVqR7Ekb7HIltYmgJ9VlmXE8o5PDsXFiIWt86dPuTyvvsQPZ8nTXuIB
IGFYxK/nVdm6KAwDOCL0c1+O5Hzi23wuWAPy+C1cp+ryN7G+kEx9MHaMWKFEw3gD
Frdn70IOyUcHY9CfSTjKOets6a08k0WTtLg9DgSny3Z1wsnnpTSEx2ZKANSBvjlg
aLmhWwDuyY/qa7kz78y72b7m+U+7bdf0/qMRvgzyzfNx5S+LHLdUxHmDq2fHOnus
0lHrTw7xFkSfrupdlbW7OnPjKMGGnwAU1pdAMd5cJc1U6VmkeWr57s0/MBSm2hoK
H+Jgsh8VFIXLUERzxPeeQkvWZMjCd/XBQqtQaE72oScjzMgIt4ngBt0Y72RK2d/+
`protect END_PROTECTED
