`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
38RUOq842vRnitbTEQiCamhNfUDm2OT3dVUBNY6xl552fNUALsHJ2mLeHG+sO3wT
57DXAWZgn9qXoilM6od0T2cxcV6ZoyKIAgVZneu+eaeDk5myovbmGR+PQMCZER8k
9mdWJYVX1cOFuxrNJv3b31Lbl/3jS+66kV6jJxcHOk8ENBqfTmzq1LkxLjjUlpaE
qk63+5/uGqVEmtgGJQvnRBsvRsy4p9KSSTRx9tZUtJb33YDgiCpHMBr2EdvbT1bI
XW8yO+b+k1AMdeABWBABzwnva9AkHENaei+sBAUQh+9bow4wDLuWsoX9sxmJoYcy
X9ssdYRSVVkm43B0kmX69OYjWhKApIH92nGQInc2DhkvsPikc3NRylEV5pgO52po
TeCpzm5wqDousmcPs/IzqJIA6n0c0YlhBGbKXiN5GR+skRJGqVzeCstZ+6qPLDR2
JX2CiwUdFsCm9Y/UoIo3TO4N3vyvwrQ4tgKB+3demdgdc0NKuUVcTSiCDvadXNgN
WbkljE//6fAUFoSAeOkAFMbl0dewYYDOSEE1TwuhJUtTwbA2QNYZ6n2ButsJoKRR
0HLEGRm/dC6ExHHR/zok7EtYtUQIKfRolb2gKBtgQQCGx+qmOtZiZfwA1o7NX70k
tVbAzuV2JMGBAKtISbNEnBRJwJRZkukk/tdYUbib2HafzQ3vFE8hEUEXAjqMe2ZF
Fy/3Q10tu3+eYTEkekcZMI6ptZ5dLtp0TLkrQmQq7lQ=
`protect END_PROTECTED
