`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WaLT9i4dkRF52U9C1AKCTmyBytuMCc+k6xMcRRWyttatNJlokKB4LnReR+HPG/Qs
D1k1PAFcfS6NukkzJn/VHFXjMP4hjF5GNj5iAya0prHXymY2NMMGv2yocCyi9a0n
A0d+WbrXcjZi88xWwF7s+dMPoA8Cn4lshD94R3ZvcID+aoSrEYhkKYwBoCn0OUE/
7saVfn2dSca3WoL5KHSOkAaozaX2WbvhnwB5g1lapxPpC20CSGVRZ/Tr72J2Minv
LsqFm/KWt86/l+UxXx2ycngPHAl+zvaohdrPMHCDUERBNiRX28QKH6SRHo00T6yK
2/zgjkjF4ZG3IwLihJaOp6ozotL0p+QTLM0Y2Xy6+/9ZObkH2VIihQLFxxIr04vu
Lvjo0136U4VD9AeLhN4A/Ip8spgDStoBu16SK3q1tCjaUGeEtc4cMn6p6jnDPt+i
h+mqlnI47b5vFrfqp59X2F+GO9vjXpGqa9LQ7qoW6ISplQ+5YNaDD2nTKG0waHDi
IyKsq5oTaD8jtFd0rTzfRSUjkpGCd5U3yTg+tYROD3wgp9r9vh052HCokjOtmLox
mjWXXC7JTLSq94xfA7sX3eBNxcUx1oMVtOI+UeBPMvGmKNUeM9dVhzBPaffe3Wt8
wIu/NdMp8wop4dEfESZ0IvDCDAL6CKwzfOi8uWphXp1iiOh7qFxOGKiOqwevOxm1
lkMaBfTelIRySSeFA6vTPg==
`protect END_PROTECTED
