`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0JFxzCLhmwuk5z9K+pwPFDyqK1acRwQ6fD25SU/mN0GlUobOdzp4hL5HM8MfI3Om
0eRmusxT/1tDN/2Iz0sMlofbliA4hvGrO2RBkUHajOo9qwqQgKrQMvyrkdX4hBax
rvP0LouBj/0g2dGa3hY93V2JqA0BdC8u4pNNN7hSerWBMF+15k2hAOEf/8pK1P6l
xflJPc09m27cMyG2G02ltiln2E7DIGe3obcfi1e1dIdJ4yUV5MGtuTmMohLPjLxi
KldHzDMjNgVjcPITTe27tKTIYYdWa+y7l5AV/EASgJCCl+xI1vNykWYQQO8THND7
GgnhMo6rX3mr1p0/bc1Hxp3EqjG1AdM9jGW9soCm0koyBTWpAjQC/0mqhq2lCfVA
o4waEUPurv7FbS0MW0H4vrTFEE9diZ5HZiH0ujM2HFAXRHIz+6nHFZ2AKyh0A8pb
m0JzatLwxYBJ/hTrUmY70P3Wqtrhq9yN7+DYDaGP++eklI2PsStQ+aHC/DSkrZ6p
ry0gLaIzDbIG2fr+2wwWtoTkE0PDvqu81HR9hmk+YBQ0py0VqAc2e+A9IU+o6KZJ
d1QybKNTWFCKX8gA3WC45OazzES/UTZz3RHNr4PtsuNpX9J4eMJEQNPV8oZg/FQ/
MAEpLaN/aBKFMfl+lj55eb2QPlL6+QERYvnJb/IfdNv20wt3o2bLet7JYO7pSGWv
3mVeVk9zKJq9JnZ6c4F0daYlGOM0ipvJ2gm/8dnSp1T1LImYoUctDjOqhWZ0lXZ4
zujwwbrHAP2Z/kVvcyla++gQ/qqQEWr8ranraWOl5yy29yLeIFXyRY+J9QfEGpwn
LGyg84oAsgD6+YS7xdQooP709tGXXdMmUuayxKunj9l9++dXJe1hDcnke9u7+L1I
9muLWilqieQI6IzjPDHOcYQ4DOZMJJyD2TlaJAKwRzFSaRjEWt08QhZwC+/bNg7J
CwUtrryPqqvmjhz/hCwTsu/UO6utgp2981UWZI8iU/mQi60YjH2Ho1YU3lUguUw+
2Oy2Ns0ucDa/tW2SRLfspS20YMOf87Am4mp2q3DDOfIptkwfJSq1TYn2jCagjyQD
nGrT/2PiNXR9dUuT62LiABcv8K/DbuMfRgTba8L+0xBsV1x5osxkMq2XaLpsLkVi
MMRluoT2jVnpnqXBdvNpZBOHoYIU5ZYHilrnsLmw/BMt7LdWzFB3UCvKuHh+5rl3
wYnQaEOKmBC0/UZknuDCt4In7Q2QCN6smJkoN+lXOxIcVyGQs3j8CURfCotTCzHk
/YyEEqeCuI3nxDq3ASB8UBx8uF36ycI3KZNaJVRGgdHKHitADHubFwcMduDvn0Vv
O0ljv1XYePPTz4CaO6REP6AKjekXQ90U2bhjTgxeR2Gnmi3dek7zNXpe5Grbl19w
JrpU5A6mcDjY5ZwmyLCgxOppIRaLV0aRo98JIn6+xt7wtZIDAsRP13ovYUWyeekR
xRODbaV14dOGuthZ8MLo5/YsD51R4rAqIbEVP1LpgPk09/pIuHR/QVUdsI45KTZL
N+YWl5cKnkNEUA5RKD+8vCICZQPZQ4n1ulPfFx+u6VjbHwbGNRnVMDiaJCzjvjoU
NmIE//eStlGIEP3Xum1hys7Nh8tedDBVUL360/u8uKnnOcOY4013TQ1T0SLeS7YX
8S5Sp2pby4sW3m/E46ZuDrxCvZnfM27H9NMH35o4sspEOi9lRqzUWbrJ1X4rLGka
NCZsX1ffT9TurNKaFTgMRwHks+2oQ/o3H6BYy3drS7dcPmLXQDN/2KSL0PTv0xMl
SmKt+qDVwmUiB0a8UEZDbF7pvqxVknIi+5LK7oKj576PsoG3PP+daPRShoJAZwGE
UmHAmEqm6ickcjcPHJwDvm5PlGG7FELouNhzgu8odVhQg9cqOUTiAirvh0vfVVpa
WfUFWzujIBZMe8HDII4XJ1Q9SMsg5rErrHRIiktJb/aHGbUlDzUsoHLK0wqrB5Ia
BO604OnpM1niUo1YZxcQQB+WTsFAG7vXWrCexPFZ9h9RluoEEn2ly8Nj4j6SvGxE
z9Dd0arPGqzG1tE66pewYMFl07cLkKumdKG7BKlTayv/jGeVLDdb9mi4isDxBMY9
7Cv8TqcyqVck7ylhdnjG8lkgQlIHpTt+cUgzKc9G+yr6EJWvIfYbZ5B1Xi8MvCDI
dstjJxLT3NHCs0X1o2JVT8gLSE+707EVXj7OpfMMlYBbQoyYxnAiIEzffq8Bcbf7
QqDC2d6RZXSjc94YHnP9I3HSK1Q+U+W5EiUn16utQFXQX0dksMaWKfDFaYCN861x
PMAtdpRzrso6UdkcQNjsTcjtGuUNRql8o+45+eAy3UTqIe6GzCAjCerfwZZSsmaA
il9Rpfm3/eJFL9kGDIeG/aG4Xd823cBv+SIyVm0WABTt+41zt8B0rm46PBr08BiZ
vFpS303wrWK0/bxyoQDNSNbXaUHwb0JPUbYygXylrXm4UlVtojpWg+RE6kLonyaD
1lwCL9p0LidHYmIA5Kc9pnm0ELQAbxX+74oeJmVdupa+S8IC6+4p/ALKLNN2xS/S
rqng+bIW5m07WqCFcHg2Er/zqZDuybdbIZlsUh2myyZtANteqr1hDAb/j0P9553J
tFAsSpwx8k/8SThQ949cn0QiMyuOkJHCl5aeejMMEid/mOtIu104ZxgZnSO7kcAY
vQpYX+qRxcN7i+Qy3lSWPweCKDnbgTVF54Uj0EP4G9iAzeVJYAFMeqfQXUzG7VeM
5/6njOwp2jGBHUK8ina8gHAgkK3ddosJOjhZV2i6ge4oDV1jiS3+p65BPKBBeG11
rENa7iCdX0QKzcn8UHn5z8GBFJG+KQaVjtZ9z6DLoglIJW/rLwPSPNXbQjeawPTA
4gLwg9CeQ+Rpt98K/2DJHya38aCOv4/icME8xZqkkU+mwAlVkngdsswZ1/WiZUXY
HR/lRVd7QCfuxJMJenNpPD70bYaNgKjkS7aIM0WDGm6q8RoWBJY+Jvrim7KghvsK
DeNLM+yNP648QguicHJ1d0z/cT5E0HTFNj4qx69FHDc58b/nxl9ZshurhoIT+cfe
6t4suk/WbyxI24whHlnXwpXLfhlIFP6wa97jZ6dkXzgVieMAngKVywQWjUa+UUSu
yrXIbY47je/sy8m4PTTUJCP+y1Zm2CA4Zde9I2bQT3qhmxh0iOUDuTAjZAukQeYw
/GsyLCSeY1Q7pYVay1Hia8l5eXlC43l6yScac9UYO0hSZD1BBIWyE5zAdpc3Ajd1
ZkTRq6OlqE/8UcCW39v2xg6jekh5IasDkkMUgXLtXb7dpa4fPVCWUS75g3lBDsaQ
APihsQ9qGRJNtBip642c2AS01E3BsC+P4r6w7PWyrxgL67bnZatev/WA2l3pj5CN
z3XzW+aNhhZJLZvMokIWyxiALpSUUISItoLMRxwK1G2b6NlXnQPLH7TsRVC0NA+h
YESA+Tkrpk5oF6SxnKbuh2DbmomAAXzIz1iwcYAi7aIQzkkOYSaPHmnB7H3R+S/Y
550iSZd46Q2s7KIfap4qKNNF34erknbQBcJJ/0VrBcLyBJK3V/iaQr9bI2G9vlIK
Ba4fpxjMr9ATRdtpo5kDq2OAGxv7b1GIPAPfcH4kkU7HGBqCjrkTM2xCfVMpsFnh
nNVBEvwA6qqnuHkhjzy9moD0uEZ4lQhydOkoUMzTkJH9ziE/KUz+l1SMbl3JD6/b
hGyauS4Fd2kubGMlBv02b3NTe2/3tiuDGMq6uK+MoU/V3UUh6fjHuRQPa2iTbaZx
fJK3vj4JY96vzGp5OaF3EsLZKCmxbzEsw/tdrrisPNJEe4rSPjcmSqfw+uSHhTxQ
uUfe+LQoIrTq8A1LzW4qyzGRvO3yZYvSDzs7Xz1imK7lnTXFguD/g7MS6WkSDdBM
5LoITeYJDRyFX7efgtqfcDKSR4zvAEHC9WiXDO7fpFjXDB+yJ9yp1+jddVnc1asv
/PTOhBGUFk5RF7l6HMHGyQa7f1z9Cly2ckiAI8LtwYKuSZCNu/+xx8hjKbMnaWcg
LQC9XQf1tLnutb5k9ooIsx2Ae6CGIwQNpCtO3e+asPcMQUnViIuajY9wT1BylWsN
nU8fxgY/1IHQXTsAKQpHE1liUV2rmxExXVbPpn72Vbl0/RD/A0PlFft1YOdg3JJE
hHsttokXxc8Syy0ioFlN4vX3y80Xn+hTVx9rxboKeSifhS/tpNWUOmMzU6zrV1A5
D2ybr6FicTl4PPKWNYxfZpMnbFF7BcJ1lL/1mCkbpCK8s90oTRYnw3Fxde3YuXe0
iQyBdx43/wf/g7BRRvzjTcQ8HPfzGgMj+8DToXPuy6aYBxgS0NAY81w6X8vSlzRA
gp7GAUqsQbQmNz3azlr6D4J+7uz/LvptCvP51rMw09n55BBkLxCU9U2PtGkaYR2R
cS/mh6l2ciLHB+d/OLkbKZjD2QH26mAZAamOTtOqAgTePuwPAooZPFx9GxkxAUhp
32PXXkpZU6goYQ//vIS0ARahOd+AF49X1I7SANxubv/6Upj+c+jw8Ji7Nbx8lvK6
YWZsAnzaWKYlIH/0DVC0MB0xxEuA3uqBlaN/3lSeCqTHw0I3jtF/pxrsla1yBPOR
cipAG54RR04t6ioWzbvfGQ1ren+noIwngRzvwQ0c1gm+h2LFjv/W+SWvtzicZZvt
Ocw0/nwxwWP9ZeWczt+GzfOW1cNhLlkMGyV494YdNzEv5JROXXdz3bIEJdzcmb6V
Rk1haMMbveDZBqW62YwoBlpzOxLCrtrxEIrTC3cx1fJ+8ebmRk4lZlKaeaPTBbCo
snJ2d3K6eIs6HoJBDyOEqiMU4jboARl3+9gkoz1elfJ0vuGawlVHnGeNLjMoejNZ
bkRFiyT9NSklGGKQxj/6zuVuy9SyS86NuWZJ1yt7lwVzYPNa9gjcSGQdjEifXX6X
utiD4cnhCr0NEHpIOMunJ6M6JEf+7kXwadvrccb8XJfXR9muIsywtxJzir38DdiT
YFxteEw74YDNtItsSRukIm+wQo0aS9msyBTTjLNo7smHxyZLdU4YwFzyfc8sBIsj
j8oSK9SQNjA7HekPvtPhanh1Iu1SyRRiydVSEo0H7BJlvxmR8yAExmtWGVh/4tfI
/FdJhR8HrCw3MlglGXBa91p9oOEVxWqTKbP8+3P/uWTfSYeL3McU4RHoEri27v8n
IDlNx3BSt5Vg7nMi08fI9H52rhYQnXxDrjrwIG1r8M8sz0E1EJMUKUhBd7pcVAAa
7FvCpvIiXcxBU3dq/9ACZmk59GSuYhgpRY647+AETqmRNGQ1Vnzu3+H22i063mp3
rNKZmNwg9lHHA//WVbKpRT8vr2EHWh93w/IP6bLl2TiFiosfkwmp4jEzUYjaK7/h
t6HJopEwFYcCo1B8xT8GTd89d5L7eUZ8CrQIKID7xmy6tYTxVHPj5Q5xC7jv32kq
7MtMvxVciPC6ULtudDH/8h4+Su0wXS8ljR+iy4hsEuBvMbJGEazRk7jrdBuHcZt6
uEZeTcWrC1ABTBZHZHHoE4+0hEEa5Mkzsnc/yoMV7Q6b6kelF63RhtZyJjloIMQ4
M9X92lV8eFJ41JetOK3+SQiwUkh4iMlDGB4SMs/E9rCSWWYCYcoy5LqaLaMNweXd
J7DbXbyhyj2BPfMY2uUMiDqtV3KoRzoJA0cIsDW92JbvxASdJ5SCQrNm+nAbCbf5
oDKR+wxUxbfWMVZD7/YmJ/iuvv6TMOSGuJiSgRvmUzHodAlXJK5NaSb/MBAilCl9
59WA2CTdJ6Ymw20pTDFh1BvVPjkfRdOXb3Ln5WN3iIYo5t8yBBOKXmAcg4vNl97n
UgiALQnhpAhO0RIJCZIVCPRy7u51DT096TONmtrJXLOmg1kZ2cPGTG410lCDY+W6
IZDKusXVwPcB9YMXUuh33ECRpR49Sfdnis+aAkLOSktc+7XJXxv1rLqt7BM6Xl6E
AfXIJJy7oAQs3wtO80MAAp3zkRVS36QOajgLash1snVi0nnAKJSkJroNWxsc2xT7
jnkgRUD5VuYCN+9CB7F7WpA55NP/QMx7YV4O4ytf51UahsJELFjEd7uwkui/shU8
UzuZY4WPB2ZEoraORMH/qJHcScZXWND6t2VJy5c2b6pcBfolNLga+6iUp4Gd1KYw
ZIxum0POE0k2RaLkE4eLptNsu+sCwbhEVJQpmw1WHHYKOsmyg5ttZjZsoASkf39S
7RZotzexpAWDimMZY1Wf/NCZa5+D9VmZa68+PHYXjtpdT8vBgl07sYWTI9Q/2oqz
SkDZ9mvBms/tWYYUMr8qnMSR2Ctt1VdWNuZdKp3G2222wQI97VMqbOVA3aBVzNoG
B/vkPhvBLrt2Gun8ZObSUxFYqhZZG5s0un9q/SF3L+cCcptL3PEs+qMnuas4txDf
dQdlNOhebzn0Rp8+9RukQ+ocoPfIaSn/E3mLSLg6pj4thEE7Z20/UrSssFODkFt5
4v0hoDMWTfpri6ECIpnbKwbrdYVuUm6qmnH4mC5kQy3Sy0miW3+bCtTNoZGMyKeU
aqf+mGKy93Czu4Ut9DJiP9lnWEoG+5sAZWBfHL63ecdD/dLTjdbO1T4nB2GNKctT
eS1dVA9FDdzDGb9dTsJuzzNJZkE556witgdLG9x7hn+hzpklLBxiKrGeX32uZAra
r8aV3vkbM/XBZ8sO/3lkolgsmO7G8U3xPlKl+nuBytxwMrcTDboY0SDRCsGMHwHm
JXhW8mtNW36hxn8VKVbedZ6Qlzfq3042QSWstADkdFOaLieK+sDlo9uxkOX/Jgog
QZhy6wNUkmIZ6f0LrsuaS5onlVtCuAS2Ah01Baaj23c=
`protect END_PROTECTED
