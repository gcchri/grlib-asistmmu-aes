`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pdWDirHwDowT5UGHswoJz4CyiYwpFhiqVh6MA9VAy+CIit2XgPNzxKuW/m0H6XOr
xtaTkLOWlb4/4l/R/8zKagj9X1hVx7PNB0CRX7Gl37wCgiYxKxk/5HI3qYFqPDKV
GIp7fbxWS6oJbc3QoqXGGQRCYjhMnDpq1K4WzrBxV6p7ej/SvMeeFIf0iGXMGnvR
yZzRZAbp8VIekzcZ659Nk0DuyLujjwRKr5MuIK1hdpfbfHYQBVmtZaLyOWHQY3eC
8S1xCA8nA2lgQcn+2ztpfKqHyl+Ltbc82d1PeRrz2hcxiUL5uSar82QgpV5xGt5X
ktVkqPPunJZe+t+VTamt29BMQ7ZUTXMl5ci24hnSm/EKYiGlAjC+QXiHheVQBGYy
WjGIsXvqTt0LDDdsPTf8ABTgrVA//hoCxWW0ER+tK0wbsEJMV/SZvE6a83CySiDk
L4TR77Fgpf8CzYia64lLDap7kxxh7uRfOYxeNhIekNgV2VHt8pEfRIY+tnTHgU3N
aF8QkIKC5O++NKSMWe4TSnFBCaMSZHimixasTdJb0JsDooStRIewTy10VcqUF3Lx
K2V8wQBzcimjI4NzpeOrCoyRp0vK/C/MZYIbIicUrZ5/71gdYaFMtiw+f4ZgOvov
AnmNEPYAgkd1R/d+H+QW+DYv+DI6yi06GtO8l5LR+NOkJJBCF0lVC7uGE4KJR4d2
8lGZwyJWKzWZvnvNoYIDB7DUvBORPo9JtFolY1DUocHR3qizayAEv/lRRbYRboeV
6bIjGNdQ35RQkJ6ohO0C67yniqZUpg9f+UGXN3PjLHFS07OONxZSup/0rIVgTz9U
`protect END_PROTECTED
