`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tN2KT/yXnNAd9xTwqYJf8Nfl42wfD18mYp5nBHQM18iB5lI+wslLU3OlYA0mWKQy
ekbM3FNLuLifLZyT8LJR/Fh33IP/ovC9kZzNjxq8q4y/AzsKaiB1uBQIDxh36Fdm
ggXOSylnQDCL6JHlHhUmj8usPo1uJsXue4xP9DBTMmy46GPvWnc3xTyA7bv+wnA8
TSVBfq2/mYEc2KOMjAIbOgsOgbExo/yHMSpsXNp7feOy8FEaUYaosE2PC8R4FV0/
QaZENLq3uyUZq8LZAQ1ZABvXByS97rP6gyW31zknTY/xXjmnJ1kkvk81Y63i3RzV
Vxgnq/b0M+iggyEJNdQunOu9EP7i14q51mqi0v2DBwwhWSdzmsNkcEOJD0s0FeRW
knfqk3wJq6Eq9iJ4ZSnbL3kZ83KXJm9K4RIgExkIEfFodNmc7zKPF+iBzD/I7Eva
UZVS9cH0MTp3NG9n5+KMf7nEXnk08muW+N8BOb//hdu6YdzCjLAe9xlUu+KJ3vGY
V8OKjFwMXrGoVBLJbZ4NCbbm7HI8OKRnYWmYYmgqnosYR2JG5YCDo6V/mewF/T8x
pLPKeQ/CeBZvHI0X2DNrgA9xxD1X7IH0If2onKL6zWHJ8ESB4FIXAZk+1WQt/Zr2
MGTAIHGUkxWd9it+61NdBRHXuSPjaRRNTfvzhGv4gww=
`protect END_PROTECTED
