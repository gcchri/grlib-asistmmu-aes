`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VF1gfI3aLmCM2JFmtUXcaBHM1lxz53d+/u4o7vuhY7WGokkrsgZwZH25IhFWVQZ0
mrlA959T5Wq1v/Qhe8yJso3oxwM8WTtmW5ECiBeHj2HTa/sOFocks9hg5h8m8shN
oRlV8zKw89x0jt6FcFf1qjoNA5Cb2O7s+ZWjW6m87JNdgB4jra1aqWa0dha5Vyn7
XpNaThRgNVFLKRdSIyAcX9Zf4yfQaqSBSgMpm4/dOr95TkF1DscVgDOpXb1SkrCv
eXqS0tjRtwl/BpYErsnn9MaZlF2JcB4OZm1eS1b9MFw8+ixTvxJVIy/1zFxdQn+G
/65mVHUqzMpWjtsoeRtZXmLckFFPFFGt7riUS1iCfbn9KFg9qYvgdIyPOJkc9oTk
DYOUyqXc0hzaZboNCWLUYSk+0FZtrrf0QMEWE+g6uNA=
`protect END_PROTECTED
