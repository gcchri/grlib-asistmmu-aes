`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XF1OS0Z58NV9Aj7Uu5qCQyr2Z96EYEgpVWO7yInFtuU2p38T8soVkG8H3Vf5ek2d
c5Ceydz+douJ6YplksXNh+VplUdnDn5zRImtYt1LtCltHc+XdxxkE31R3B5HSql1
gI7AjFS2LeLAkiFss4sUkFvHzlcaPBftNKwej+x67AWzUbXdLrTMFrTx7aJec+Nj
AKMew08fvHozeGGvB2Y/H1vzjZxqASvY/dvVVhq9Jd8oXxkNDnzuyLLJL39i/i+a
tZn/gRqB90xiQ1XvonqrpKIElu9Y6sBluwGnWF9CyrY=
`protect END_PROTECTED
