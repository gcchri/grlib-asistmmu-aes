`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iBDs+dAwL2fcr6wp7u4ypH+x8KB1IlXoeHdUlSZbRjvPRKyq48MC3Sq0u6skntia
PFe1FEcMoUP+OcWKga07NVunP9822Qi38VAEsvivg3gnkLrZEtvk1krqmxz5qIfd
UZKy3uyI6OwnSKEePtyegKxSO6lYzKtYTUdfmMpi0rP8m7YvK8G1/azonhxG/EMa
/ypdU2KRmDok8xkFlZjp1/BZui5hcbkOtj1HsauE2/2/1TO0HWuTSQiWOfnKIgG4
kqF6OIUJwUbF/Y6IugR7qlV2HN25KzZ7+jMi9fmVvqL+U19YdfvbKP1q+9IFmrqx
QUPYSK59/44gXov3RdvnQBjOV59WldfW0dHd9u/bAJMBkP1NVP9Fvj3NoJ7SgSyl
pWoUG9hqZtpQZG96qMGTCGOjmimN415F/K2LIleRD4gyXWd8UDGFF2Svm5/mXft3
zB3JtsG3wCR6znmQ5hYcQzffMwZIz5qWNoGDfB7gyU+hY97zNBp5PjcbLm52c1R9
dlarJplMX9WjvFScyTp5trLxh8myyEHQRllcQEFkmE7jHBGkIIinbODWwk5F+Sk+
QyPbZBXzGYpZXHn8fSRSQy/X3d5qHKbUM4I0h9i/4TIzZ0ppYx+1y4pkwusqDhJJ
3loY5VNQuOR7CMiIR9MV8qp/Bk5PYjCM6ktxouf9zh3LVPMPmAYb8X60R0plRfwR
JstsbFjRhkO0k92+yDcPEIdFluzEIpSXIL7WbbeW6ITXDWlPhW6g5/tI3hH7FqDF
+B/iU1uekojCcX1zPpvl1YEec0vGKtp3akM1pYh15CYtIJZoJ5CTl5I9mLtkzpRr
cYTrMxsvPGILtgnQyiGO2WWLJihlJqhwkHO0xHx9QvEKWWX4udXDxSx6BBt44duh
R2YgdrSqDv6cyh/BrQlaBDR2CRhc7qqCLUQbhpZYj4RFAxr3o729FfQB4UMyC52e
UNBEIv9vWqxv/PABJFEBMCPHtO1YUuYrkYWHniaxSnxK/GmyJsZXyUQQ8qg095MV
TpXEWOmPdVdiHLrnZiykOCMnRaklUON+ppwNd2tW8RxssMAQiTU6ksf+L6OjAkNR
lcRRdQafOzo3B/hxXBEXIzmbRWCvJBWk9Ej+2ZOFQfK6868n4ixQe0IxZf8Vv3GJ
tg69ndhSvieKNzFlpNbj2vwznh5N4rN9sHqaOIEHKqXxJ98Y9V9nfW5734DNac0T
AKZnA2p00LFoEbXE0TLdg3GReGpA8fImDUgWyIrurY9e8huhBRYFIbY6zSFIy25K
CqZLn9KdYwVxP5FXaoFzeZmT+48e9enbaB3JdmWbrDcCkZe7jWwABxwmnJNuEsea
E4mS+y359OC55OHTv4hb/Qq9YOrGBkpG6fv1DVC+/cGjhllfZLHNA4zs4wmHfqYp
Amvo/tc9sJy+RzRwRuURoz4Ub2gQl51+dlexm1wfIqKq6DiBXte6cfKkhRpwj7pb
bst/OGZmVl/LueGetaq/d/LNyJlAtkc6sVO7KyaiblwkZge1BJ2I81ytyTTZ7Kad
LB7YKAv+vsx2qgvUHXVRJKplAg1koCjCaXaFh/jvJ+FllY72UsQjmU5BjLhDtzIQ
tcnPs6f1fYndEwD0efAekthUPv1CNDf0H6oon27XWrJiUz9wHMybnMzohrcQgRW+
38SOTNm5SBKHmrLTXaS7K5oSkPoALSrNPwG0LkdzgCQb7+dXXEgGTCk8fyZvtFGS
OTK8hicJIYPhkMA5h/4tNcBlVM305wCO82lc6Rt4mcNbvBsK7gIdx6H0qyiJpZ1w
OQV/u1/0Eh0dVos0XDHyMWsjNnKIbqS38aLVllVCROJleaeR1NyOBMXJry4mD1A7
fXN08VeG1zXRFd/WU2NTXhkeSdRWHvMnii99k0U18FsMG9xICoeYoNNkLfT41bdE
fWPXoVT5tKIjaSCykbLMxztqBR27wXB7MhFHNcyRSqEWZHo1sGYUGbMfSe+nTWoc
LWs0X+fXq7ndzojSz4OU9A/GR1Ac7sskuSZZB+HDMlFn5hg/ETtV8rkYeu//S6FL
dELuw59TjltlM3Rrak77n2ibxDZebd56CfzxucXpTeVA0rgjfFokSjO7Jx7FLvDZ
BxwHfpALEq5xzoKKwwsBZQU5TQ+8o6U9psARxwMiFv2aLguBgk2VGdT+dsJ1b6RH
j3yuUbRu713jxx8406uEpONB/PAARNdoX0lqw/ecu2YOMQYtAltFON/fS4oR1qZV
oKnT2joYJrtmYJZShtmDoy1A5R3Bo9qWlUNPtMIsjpePPFxbec7bzutqOShEeWnu
/aSP43PmCFJeAF9ibWcUoca6Wn5y3zPglOwkHsVwPNgpsY7TfGqIzwi10SVyHLCv
TtMxmiT7DVU7FzLI9yWyOYcci4ZTOKuqT9m6cFRtRCR2i8PUoIPs4Qp942Y1hyui
mgPj/tk8/1BCgWCWvGPQRk18iYaChYJYObzuSF+SX8tjw06Wx4q3STPK6YVg96ak
1S8fG1bbiVOar7O9zYcJNJ+DtoU6QSNtHvafErQN9u4=
`protect END_PROTECTED
