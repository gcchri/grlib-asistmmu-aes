`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pXXhUGy4qCh1S0xcKxnBmJv4poatoyQov7181HcEGx3OMf3wPqjKPmSzlnpZK1PK
/9kgU+JcUo9Y7IcXwDXPJXa8PxZXqqRGPuuud3A9ji1kBmRr1qBXwcfaQT8TTtTj
+/ELGNxY6L4DBJvW4ECdhICvIaW9AvmIP/8V+KVSoKgW6dNNrSRgmvBCFKQsZ9V9
hm4rJJMlBh+8SxutEWqNcUbk1xt8HKpe+J+egeZF/shF09b8vuI80CS9OQRh/1Hv
cEq8kHjC6es7Hw02s1DoV90vrFgRPcC6YbIeY34D63pEjaxy1oOu7zw8gHBfOi8p
`protect END_PROTECTED
