`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lQJyXO9l94wj5/KkJ3GNdiPCxHxPttChQpFoFsLk4N27qR8kxAcP6IUJvRM+AchF
aS4K8zy41MfImDQDydcxSHSfgDsI/nP6OyOFr+38rPCW4PGVCSNbb88VICpxu2vQ
w24B8wmO3MHN08FiN1iWHd1bzZIe8jTAfX+Rb2vjc9OzireG3z9IDIV7YGaQ9VB3
+U70u6BdWKUDvCVQ0FpcUPtUTEyBkIDs8FK33HaUDxDz4u4gMYDANpxQqUePgDQM
aESIncjOY/M5RPfFLNxBjkkl/mMqdHgdM2DEDARnMAyHhnQlSVhnGa9rOK6shk5h
qu3B9dQga3UvF7UuP0nlVHdaOLQ1KY6IYhn7LrOR+sL6gZpMrtPwcRYv/OEwuIT6
9pOesV+08oErKlRofemI5cmig6QiVv0/CCs+WpQf/WgoBqLAhFlz7jGXV1mos6bu
T750XOKc11wp+XZtp3odctJSpgNAYa/1J0tTtNdMlYwy9tOXQJeClt8v+VraPZEj
ccwAhkB/ZS9KhZuZuD0Q+vD7hcAbnf26mapUHiM29SyZ+ebLiulfhsfz9YSXnLf5
6fVUpy2+5CdpfNhAFCqtqg/dY747bOCyiV9kau75VJyi8+t2e+dHlSVctvZnLaW1
Oe7rlVUtWkYEWfldnBz8tmDJpv8Tv0m4MXXyEWrGSm8IVnW3yj2Jm8wn0mCnIbo6
rsOah/PNPHuXbTfBUjwkCS0iM+APbULJfHMjgjX67R4HCGwpvfKdkQF88QD6vRyW
A6k5iED7vk6ouWEMZYB83ztqr6hMxXS5fwv62NouFYDVxdpx9gzB8Hj1669V2NzF
jBqIJ8y7NjEw9gkQQWh/aqbueGh8vAPtSGvHiLMVjm2mQ5ipvFKdZmWcJ9/JLPkR
4ee0+O0FO2wqRs8Evzs4Obwc++Siky6Iqv+H343y1YcH8du/6d5Benh4xauvigNg
YsT2MFPo4EpF5+QUyDeFRqApWJjchE3jJRCQ1h+mSWNdyH2aC6k3FrQpnazNbSnP
HBNhhlhiXbdwfiq0dx44caEznAat8cfXVbgABDHwxKkm2XTgDrGNYc8ap2VBUbLi
L8qXZgE+sFfABx2dGu8XS2lBvlExh022dlduNB3pbhm3b2521b4myFShk094o7Y5
IDNJDOFpBDz96uiVHYpWD0UHVlS2ej041RhDmsiOx1vL+sdypq0rFOYkBbbN/RhA
veJ2UazHRtkJB3yW/R3GMTmPr/tz8bFjPcToFmj6twQrJIWhuUuaJYhei8QObtww
lgH9vJER24dQyhFVNbNFbP2uGbo6XT0tViQKkLcs7Y6UzjJIsoXirplhsEuxP/m6
+0ufZZ/Co5/uzpi8ZpyUC5nRUxKv0TrY0HnLgzT+aeYXlVzJSF0CaneIcbXWu0lx
SSFqPQwY3A+JKy852Jd9VPHuYS4mgU9it/XN7RzYRrArU8FeHr3dgMGtB1znrSIL
Cip0ElED5vMGH+PuXtVa/WRBU0Y0P2coKoc00iTmSzSL79vrj4iSE1k1x4fF323G
mz5IWi4tKYcJ1zaTVQlKbjG1OvLni1A2M+W/iIokPbPlg3HcG1RiSMSZZrArUG7o
nuZ+vMbfVzsDJfLF2DbPqi5e//mn8qkyPCncgzG/Kh1FE02HRHI+ILxH+MuSJm3x
BNheFeyROlR+/C4fhUg1tfaWXMAI2HgpMckzgnG5OB8odznFecTkrGP6Gav1I6Z/
eXfK3TbCW0M9OQnsdvWZnCJyq+8ZBtjbu/y52uXo9NSsA1XB6ZsLrPnLro9aDD9y
66UardLIudpcWbeHO6Q3up973xFbmevLU9sBfqEHz+B9fzJwfLYKGDH4hqlJKqJH
PX1i5m1PqOM+Yer72sbX/0hbxE+go7z47G8wrGyTMhrRieJs5r1mn26VmMqGJsB6
`protect END_PROTECTED
