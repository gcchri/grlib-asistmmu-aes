`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1rfgLwYq6R6e1LP74kI75X6X4Wv0wBqQqEf1yBTWvPe1DzZYLUaTq/WRxQCL4CHu
/OCEJdp8Yhyc6ltiLAXof9uNa3uoSp2l8Eal+0nsM9Q8z/vUyYm3Aa9pytqnUBRK
sghts34tB2QnUocRylQsGRNBQsAY4dX7+XmVztYtOjwYrKWp2vfgfAQKUtS6DXrJ
Jf06AtridnloOR9GoGhYBPA2KNyLVdyUVnZQ0kooKzY2HMzT+qGkSG6yhEalzsfv
k2/S2kZ0K5SKqd90KYzAkKvnIwH2pmZeVe5GfaHIFlNZ2AKSMKXhZt2Ifxjqi3hX
NoIqWx7taGlFsx2baTEWLTS7lgmhyFOt5SXyCQOqozzfjjxFd2scg57zmizLYJOA
fyxZKtWkDyfxhFknlS6bc7OQ069/raSRTobBPhuB5s/et3jrMe/jNz2WybeEku+S
IRLarGwhT653QgC4KG+FdJvsaNrplwKpvkiHhcJ68T4FcyZvdpA9afaawz4xLGYk
pHBv95GMHfNj4c91Vrhxc9SLC2y+WWAHg2pyaOK8PXZQK9ugJdu0hthMTSfovSaz
cgpBd8/5Qjz7JAXUeDQch6hjs86SFO6fW8c45qkb9nRamiIQdrtBD4gwWVP24nfe
1w3WaivvULULyAVNzl34tAXq1qxaO9qvB4K3BVT+OXpKz/eqvaUlnW6Gb+uhEcGW
W+oKcRqJqFXGGDT5/GPuz7AgLMZKCG5dPnzcGtgLjgU4WuvIw83yZ9BoLiGqBJng
Z9Van5HoaGqac3TiZjxZQQ==
`protect END_PROTECTED
