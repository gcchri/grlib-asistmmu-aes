`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PdfWVNYEBNlB9KP9OxifOATCqZHA18YglzsmATushRmgislPpMNaY8Jk6XwwZg0l
3Azze1qOz/Xg2MUO/qg7g2pzXVHGtSZMgH+IpeN6xbsxJz9J/Ny8+DoPUZp1wN98
jVSVtzMW+0RttTfLK3MdG1tYGXSsB6mXz+/XFRivyglgisiqtQ+Gq1nIMy/GYYs4
OsMpu0YprRL42181Dx0U9gGA6xTC9hGr9QgbxhcWztjDZkf/op8dTnhkLr3UfHcR
Txcq5nknF1PEZMBJKtS70vcdfzZCYaePM+CFgwjPJCsZ7CccAKTpIYkz74Epf3ty
oe3ZWBzM4NHh+vBFml6p+z08D0z/A9K6abxCov25gPb6fWwJhFRY18A5aqUoW5So
XNY4TuM1DDJTISBKzSV2XqCCNNVfpP2+liqR/9OuKXutSaBhBdd57HBP91xj/y6O
avzZZcRWFWDZvLNldTEkKk5x2czGJ2bR08eVem8OlfaHrVswpu7NXQcfbxgxtK9z
kZ3eUKyLhMgAPtJ6/a5U6pR7Jw/0/Q6kWpfbs+3gMOCwFvWRyd22THP8/rbNboVC
bMXVFZQ7RLIpqD+tR4E7940pPbIiatQHEjgYSBuyNH7MsyPdf9MQMIxND7cGUh3F
YuoWolzHC+hTyQ8VGScTL8WQq9zt47xUywkEKgKOsAzOzEN3d/MsYGbH+JVOml/g
AeqtAF0hCSGbj3SDX46bAekzRfzWrpP+SHWe2dQ1frcxQmSJXlVBh4yzEi2Dqfgf
+A6ePppl7suPrbcymGHTuIyJzlDA5Ji2lhw965RySZvf6DYr0dRBdUlLyta6L4mP
R9IcbwtYyw4gKdugimEu657eoTXdp2TXNPPG1s+6tQI/IJC4n5HKPfUKwDMm45uu
FLfNC+9Wa92/Xc5xk/VUCvgZ/89EfCMl9GeOyruXLOKrze5psCxmOJxkxvynOPxl
QtDlTu4Ps8SPYANiTXOGSv8aTl4D+991T29Zpwkv3bBjMKb+m/pq7J4wsJSU7cF5
ewqTQcG+xyq2Sa918LQrb8rSwP8zCZ8hqAZsJHTjbySqYHIQkK00D58OvxNDM+GF
h17gr+2INBsHbp3hGUMK0CUn9j0KtLTHtbi/pmoI69sV7BdgvGqbIlH8kE24+jOE
`protect END_PROTECTED
