`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pGklak560TNbus0CR6Z3JCVNF46Hv3MqrHhmIIK4fFQTzKfbiYxbDGf/eeeWbKTl
VbGuXbYTUpIPzjmVNn9zY/OBedLX9nOj5a8nDOxuZo8vQjyAytelIViBc3yh8HWH
c2wnlWcpcwHtiieI8JnF2HgvGh1GiZ1ZK+QiSgrWQbSmBRRmBb9NksyTdy+XR0Y8
ieTUq4gXgtjh3UChjA5Ord+qQ+mSFpJSrFXkBomkiVlS8m338mf5V9C/U2EZ+skA
Cy5tE9pr9jZPJrpjqMvExQAIYut3ekYRo4+h0v/0JM1z3pvLM5HvbPCyV/qNEuHj
ZuE7asC8cglI/O9GhnpOHmmR7GGrWyhoTXvL9Wr55itKtNRyJ8HiIftNQZCyaHLs
yUbJta64FAYjKPGz2XcS9jvWciil4jS38SV7/31/INV3+e80Z8R5+pKXfF0Ww1Mp
tAbJerhX0EwUESXYru8KfD7q2vSb9k3+W0yhXWgn3xFLobsmiiFP//UFMOgj/Oif
otf9u6fnUCF8J2C9cka2rE2vokYf5N+9k4ZsMow1f542pgOynIRzwxrX4D5NzvuB
b6kUENjJ5z3fvnZi5EH0aHKVd600/z5ju/uHuduEEu7Wz8suw6MB8wKHTOm/Mnv5
QjuRu6kIzDlRVQjBbTAqh/kAiI1X1Ot2CyFeNwwG/Yr9qYBQOg3/VEWoBkU6qM/m
R7AhbGQGGf+SuI9P3qkWSS2CHhx9sPA4cBvpntF6UaDxQXNeLtSsyELB4GWXRWDU
L/if0y4i8pxXnZhA5WwBdq5R/e637SgS3CTjks5BbNQyuVU9uQknvFPr1SqlV4ED
yL3cv7uAmIvm1GEQmY34q4fWiapqswAy6bmFyE5hs7+eZVghadAnNn7y6SFuGbgb
I5KTrGc2obFma//4ZeJRnozaTlh3S0FRCsRHdC61DGybG179bae2uXrjjdjNpxM9
7aGI6POqODpyp7A96WzqWgNIsN3dg1OstiETUFPR5VUL1FIRIfSsat/oVPTomF5f
E98N4lUlJbJtWz9THWNJqYU87IrM3urqwXkrWDls+bbVA7np2+PlQpBEpAAWKJhU
/fvEV2g/wEl2dK+HymNDyLpLBc9fLGUS1lrAU7NLyC++K6ISWHKC6V0SwKBezSwy
knskcJ32yV/9aMkpzME+a0opTm1kqPBp3oFRFMOF8Yeaxd3+lyp0Lt72QmBL4LCo
u9btPpV1IJF6qreQPEKIXcnFCUsIOyDQcXZ6q/eaQVPDTPKtgDyHYTX9wf+u8SA2
n/LXcdx27Eougxb7MHZowGu4Uaw/1THMRPEYI13Ykf2hwhIcVpOqTXE3sH3om8q+
L9aEPhim05PzxdyR8FXYwUHxZFrsXYPtVqg2Z+QPYx5dC03gXC1IZafX2pIEkcWl
hAbKqjN2UjmKW5UJgw1A1lpcymew9Le668+WCryT+PLNMqqcGHVaKXpxMPeed3JH
KJL5P24Kqv3Mx9kBM+R4qHuzTARi1V4Q2YBrXRyvDfqkxMXu5gZ3JUU3I8T7DouB
ohhMZH5LsuzqBxrhI6+6i8U4flixl3rvG5qGxesR6+YcNeXli6wuOYA3eaiavVDZ
2FjhuljJ97AzZqiHDR76dhP1mZRUsspYzHm6Tu3gsMkH28oIQlsQBAZbQAGbCeeU
kDBELpHRK6rrgsSqTOCs8mWD2Qrt6GY+swljW8DFwS3zQtjQEznI0r6qQSPCFO07
OUQ5+6jigMdoiQJloCw/BRQA0GV5DhW1AWaDC9awpHHZFOjFDA7AENQyZS2KCzFr
BygME4mtRYa7MhGBw1k/SSbZbcU77SKc+8unyxyk6f/OC/NdqfS5EAh/AsvrQfM4
U+gGUjbdg5ZtcaRXx7kSB0RsohlnGA3CBzJjQYY20CQ3O3kS+AL04MYb9YJclffO
36woQnwkdhPAj484pgzJUy3Nzg4zwBsl2bErD3NpeBgG/S04rASvJkA8A7iG4Gue
HuicA4CWlFsoHXsxdIbwbBSFdYDR39+CT4cMtEA8PGWlI3Yk+CbkX7ZHEPlQUzys
zvqDmsaKaJ3cE4xPdRuOov8s4wYy3OghNDBth0XmeIvleT6LYtnDmkKzx2o0YifU
DlJV/ijA+uOQvqgsHXd4lLHbWy8SWEmdsBpM6gV+RioaerRbQnjNtSkzbW9ipOQo
EwCKf7gMUWZt84p8NhSvgUAjRFBbrrZgOH/+HuP21ezOpPJ5DeGVHhk3xphB3ABY
QfOufsbjDJhS+bjbIokpnuViaZUVhWXAe4wWzoPk4ieuMGsLMZIpjHd6LQyrdSYM
vpdyRai5duLGUywRboPYDDXclsQ+atH8O4d8LH/MhCl9oV97I3ibY7KElXNFs5MA
ObB4FY0BFlQ1GprcrZEnqtPkoL3dhuz4P4QNljX00mXYC3cCuHPIAi6VoAgSQQzH
kKuUZRfxDS2Jx1xhxFAbOvJ5Oqv1E/+9di4af3iTfZpqhp4yeqqjbGC+cPI46htw
jXLCgUWJcNXJ94ZZk21FZDeUF5cFy0+5qu72GyCEM0v0VWAv3Cpj/tJrcJoBI4+x
vSUp5t8w37dH26ZuTQxsdKKspKWuoQI+fvikp++0DWupKDZkdkS6nOH5JydnAp8D
7OW/DwJnfgKZfZOdHSfUT707L5ItbWG0eY/QDpUrKMrM9KwNQr2Wrs5J9o8E7s+h
IAi704oBWFen2gKDbm7xI5FhYieSOBNG/39XJkOtOWvZL1+Ndg8VjNQmkKbkdgq0
XBNaEVnhzWrxPf4mIjk+RJSYicEK96xWygaiY53N/YrThapsLxqzVrGGNzoWXkeN
nl5Mck8fFhQzYR0oj/5oPL7w4ZRz6NnYFH/wTFRrb+HUKgFh59yjHsotIe3fAV2F
7nt0SgOzFr6UPqjfN7o5IvXM/7xPZmOr0f3o42D9Z0v0S2tgBZQU5jf8c/WC16IW
Rbt6/Ny4wn8wFfhtbnyWIE5qN4Qv4UX5HpoCJ0xPOjY=
`protect END_PROTECTED
