`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K6+5kbe+gmOoUnt33zzMZVWNyHZU2IvORJAoU5tuMAQ0nfGCjvWtYa3o/2iYE0U8
PeQ9NFnxnzx9MAw7ceAo/ICXlQtUwtF8qvgkIbjOhxiyHkgZBJQoOaNwmIEmr6l6
JpPjQfFRRIx23fpszDm0PjTpvIidDIKjuzMDuj31BNU5SCrXetTUbjTpcwZS6yxE
TfZuOhK8Rl8vFbbAhLA9GptQcAmW2Epf5TZPvs4zIqhKNK8YauwpBDm85b+h65cW
3TA/ttpq15uOrc/vYuD2dHNqX1NvM500bA4KAgT3ltv260tXQike2AZZUq67cCgY
l8/xlW4Cv51jSa3XXZCb9x9MD9Pq/E2Ky3oPgMmFlQnL2G6eA9KDZ7KkdYsQ0XK7
mroiVShAGZ/YEVYZYqaz7D1Wk+gdt+GtBJiUSZ7OotvXBeFOFW97H29X0Cp44RpY
2Iz9YnrFIB85GRbZ7HUaOhycND/CmWazPDU9TGglgiWeiYkmuWV7ALq2IRsY8aKa
VQPYrOQza94eL6an8Fv4/zanmvK4kj7TtRRI8V7z8s3fKeTCcmqNGKv1XV4x3YiE
VutMvzVZ97+LBMAYRD67JpvOGSAYiN5cgGRmgtyegUlaYpvmtUtFKpH87gtRD/iG
KhhVQsFlfkmIKcbvczyBO4ZMYIyGGLp6KG8VlMO6LHGRgD96F/Ix6F4Gg7x+iWP8
xDFema7IhtYnijSxACReHbPXaqhzeIqrw6/O5q+N+WS1tpiocKAKeb2I5wH3tZQw
LiSPeSdvbnFyUYXiGyK1RJ/kqIqgvEzICbjYzjVaUC+Szxgsl7UU8wzCqGfg4TtE
I52nEohV3EsI5PXjo7Pw/5Up5t7Q7gYc7t5joZ7R1HqQf5COisllYLmDiZNhG7Cz
31RcoHS0FZJwajFEXeNHQXA57VCC1wIksH+tJKvfweGSTXcML7nhTj1WyX8HakLa
4MmatkR4kV3rn1oq4AQBWChCNoivyUbryfxw6FNC2tyj/+YuXeytGspFRGucC2D3
Us63+M+Gkc/aqMQ1Ia7kINDFKFM3BFx3EQE2BxsE+b/q4ZP3VA+uNfpVp4jcQfIA
k2H0yXkDPScWikIWYpeFkNY4FYH9WmeNxUpLOG5HDKW/vdhIiJh20EVLP3qmQawh
1X1bqO/4MSUN/9Fe5qLMo0K3u4aQceRQfFJkGYC/Jv7Pn1DdQZRrWnhDOyYHuF48
bKQRQKvJ7rLdf3R+FVUyiOc1F5FAynFa0KqurmuK9GB79QxEDtIr0y1MlT2T4hO4
gV8vqiVhq5Q1m2WxHK3f2PV/7r2t82PHiuuRBlIMY93pXpAo+G0xJqpSubWlqoab
wr6uf+sddns4iuVIukokKmRGx6AF/+k/TCz/OGs83/we9QeeK0+7XCWHoPt+PcmC
P0BhCHbQqLx77Hbesvir6f7ERTrBlamHHrZ0AqbrYFfzEOkA3j6+zl6M6dCNE3sY
wsnHfM1TA2sdPFRdaIb7bH/2QHnpDr+EXbrvPbfPmzLxr3Ovc6KkLnHV+ksUpMu8
1myA7CWEkUQFhRW7H+Iu6egjCivaBwG9Ys6YTMFvm9o2rieCZHsxy94/Sbz98UTv
ZcXsjTK1FFYvfT/pLxVi7/DFQjKOQPgcvvyOGwqOC7iuJqZ3drhfwYN0wr8JzPEJ
FmyP6mFomJVUCfoU5HpoU7J7xNuBtyotGxGdTFjDvBVi+DpRsRlO/TbdZtvVA5xe
IXpe6B+gmHwaXLXbLgRMXMvHzUzFExE1a/GDbnT0R351mwrsh9d4kVltFRaU0k9R
wC71gu+kkHQOborrTxJAUFiy0v1Vt13Ol56R/5j1JLJOnYOa/L81uZXuwq5lYa2k
gSfcxWfDUVLNdqELzAdXb0IrCArbAqmB3e9k/2Osbh+6MhIAYCJqW2a+VxSmCkdn
ZGqBsxhkqrPBhLWqMzKY6bHpIpll1WqaVsZmNI4DJantQCIKFCJJ5aEibUdOXMxG
NAFd9Ipfg27S9Rf9zmKc3aG4T6kczqF/vIc4wyZ2xLdRERWyVr4tkHThXIo5n7E9
8nfWrjjhPD3JYqS9xmCwJG/+V4QF/dvPF+ifj/U5xmWj37EL4IHQ7MTRm4bmCeww
clWkq3aNniOo7ceSXLZ9lmungSbP5G+N2z0Gye3LnT10/vmbvEpFRBVdbU7BmDFz
2ugR4Ixr8bC1r8haSeSh2zPIOu2fMlFAR49LSDkPmzAEsHpa8o8Yj3D6g7qM7K0m
c7NouYw34cckVqRCURA6/sVhPD0kO+kUpvmYw6kgW5UU3DPd6LH4QB1tiRwaAWkM
pG1/T0Vze+yGE1YYaPQmEznf2PSoKhwAZOq9krci+KDmBakLvaU2giYa4avj55YS
AGZ21jBUHOPm0jwxp6mT22wwV7oB4qMzkEl6GbGFfKLqMUbPVMsygc8VDf2P05tq
EBg3j/IdzYUSFL+0lwFgAQVW+uTnKTp2FikKvJ9G0siNCaxA2ZlJ6fguV+9XevkD
L15PzMMWjLVyeaNGefvwVH7ENe8U7DO5ucWXeJ3TqY+F5JRKPRPGx2MhxBGm1/z5
68cp4grJ6UYsWXXkdMz7LzMVkamuhS2p9MvWG8ZwdcoYw2Wtu4NL2QudtaTmWvNZ
ZTZ1CiVBEjmJ/5BdMPg9ts99uhMlSXNsT6d5lifsuuONBrUyPIS7GcWvAGRJ4vuK
LMzqHKgjpr+w8SF7vtzu17kkMaataJyTrPK0THrysinWVNOgZl1/JFol/l8Nn4SF
0KxBREVrHvWlXx6odAXaD7y0Q79bo3XEFST6XOTBMm/zYz5Aw1xGOlPfzbLuX4lu
9UHpfoqx2baXmOYXtD2SE1FLF1FTynzBM4h8D5NW/LcVJwdv9RdEzwfmkvIZHWUE
m/zfQNY4nCUvUwQwT/tNeoDPd2GqZCaH+wxHsQmeJW6ZnjRbjegl16K137eRwgc+
Is0JFxhYqLbls55kkPriqHNGjYoapK71uDSZ+vRUjPMDsVOYnR8AjaqkNDlIUCv7
baC5qxo0iOZIoMXCqOBzSht7p70Ah3JN4S8DZXp4Ah3Y8NuOQbeyflOQeg8tQOEy
1XV/oJiBqs7o5hLbNUyFRVR/pfuhvQ4DXiqymo2IjUWXDex6fpW/2a/J4OaaJGiK
exs/2JwyQeI7TIPqSolY0GF2buYBG/M8LbpRtm42uK+XW0HYo0lYd+dxuQcfd+CV
MGD1+cThq1BtUVZovja2K0nhPR9871U+VRvLWkTHkyqgc/t5fz+0/kmZr88gjnzb
LZlRvvJPPN+uVxlw0fdlilrkh1BzdRF65MKZScswD75s2qQcgcFrISGgbRgKFS8+
W/bYSHKLN4t01LCcRU+mIBh+5i+ijDGO2I5+xaPBhGZm6zbQuBXncuJZn31sso4G
O/dPlhIi2mXNsDn4UQIVdMRcE9EpwzhKX7/2JsYGkjjaa41vOjvB/k5AhVw5u0yg
f0hhYwP1fFbc+DY7hS2enExkSKyywG3Y34CtxviOrBVW0bAXXy5HDiUTqf7pzPS5
7ZWtPlcela95fCcUJB+HcPxuArrNYKD87Tf5EPS9dROnBsIaGnKxhGOjemRsZhQu
Axd5fgSCC0uittfkWiSjifqZUHrzCbSDSCWw/AOjgdA54sChe0SvwrGjkQoDypvJ
yBmU5k+fYLpxaCeDH9m64vswn7cBNOTFbNOlv4Uwnq9A9jA1t0v8FGl5jL2oXqBk
T/2b3WeBH+CeSUzVUf3YOseBlBXtQmMyJoY9M9BUzONetHSOgpRK2QvjC2fbkTbB
AaQHi/WLHHdOynHjPewfaDlvOwQxq6EKfzPx8Mo0k5aa1Erccl9B+ICl3R7k/vvY
1JUy9Hq/QX5swUw/LxVRuk/D1pqm20NC/ruI5/OTDXvQIAwtkFlz1GYUT1TV+jiB
QAFPwG4EQsdCcUvM/ezVqlpnq5UHwCktcb1zd+esRPtk3F22Mf3p8yXKLtwEQp7u
/Pc6ueNtBKSosEIBt9BzFmBnFW10/WkzC+UxGWlsvupMY1kaW5P2NxILxGlWSzeJ
EESk6KfLvpSTNm4/G5p1jCbYcmHJeF3eVEmn1sB6394Y2YCniJ7L6pX+J9CHjicd
OZ15IcnNXiKd9NscKwVtYKyw5NtimyNKqVsP377pPdvhHln8BhHE55KS3aSifNjk
b5XzRfevYFrfWS0SMiFq+F9D7ZEKtXU8ljCt9dyWI6w4ka3vu2HfRXEEq6OHdtMA
saFNtToJqATiQjZzNUowlySsb6Uz/TcA4ZW6sKpMlTz8cBSxUTQRmZc/l1HKxdrs
2L0JbAJJHgVQze54qEVZ6DSslKv4EVNAM3WFsUmrUULRUEbwq74aX37u3UAbBqvI
n5hJPYh1eIFEwUQjnOLtzeGSC/n5ZQ8mAL0LpfN0yUjn6OLzJivzAvJH/LR6FVNZ
UpfFrXxHqSu/pjeKSD2GjvBmxxleUBqN9y5jrwRynASNXZUgsihzIVW1Zr6iYPyg
Rdm5aiefeyqnKW6EKCrdvz84sXiGDw5q80+cSQT0/awytg/TgqgI0oeWz4AxH0WD
HRdhkQ+1rr6h6607hWqDzagNBOd36zu+vPIidpv4G/plcnXQAo5CYclSD382FEsz
C7sL9cXnZ94BJT0xNXLnk4GdT7KZjfjgKQ3giSw7Bs1zlg5Dbj6+Y/fq1fb0u1d0
V6DNCcz/uucH2XbMk1FeOq72I9D9MfQIsKlU0QHp92DdstH9z1vijJlh+fN8rGdc
5KOM9ZdBTXZsc+mvqpSRCMpCICG0YCW2HeqwZv9tcITA77DqcfUmwmyotmPRtb3L
ERLaISSZMaL4P+aUsAkjOOA4TeSVdquZQYjOBlMky4heKR0hF7w5kbra6Q7zKAB7
DlqnaazQRWbWF91IzFyE+/3shkiWLuR4qI/kgd3MD9avLiSIQllnEm4+VNtX2AzA
wdIsTi9Z1n7uU+0zqmsmVpJ4E5i4BCu1OwZ0AWKVr+S4yXD57q3lJr0AYhXkvA+5
4gTomtdH0PvhfNyAjX15e3di2uR0DFdL/D9BqCxsB0fyZ8ZticADyjYDCsWJDwDK
Sj4EMfy0m9i4UcN4dbpv70XKHYKI13nWt/tC7l9/JY2tBnAK2vstwZkf+rYojWOJ
LnOk14+dgZcpLtPdtERf9z3rpGyVZ8FMiG1IoP21pgz2Uy+DEhUz0S3TUXjJPlms
Yuay1o+hsgAROvpOKxKh3U3Wb/UMaRrLoJTo014Ky3YcJjjKRVlAnDk7m4Zg3Gaw
w7ZNcKDLYXrqCIYv4gLL80lEPoMazqbVrL8EWEPxzvPJXCwNpf5TaIQkApkDeb/b
ACL6ZFxvhQrRUd8pNGtTpqUW+AKxAzGNgWM8xmHH7ttziVSjMQsSs9RWnJCjkDfO
t5liPnvPxKEy0H22r3VHyasshp0d0+0jyLV5l7iw+4uSCzMG0Uc/DQ4ZEsuTRRz+
PeFpifPnjBC2/G4fYmlPMZRRpnvBu9/UzPd95w33kFprkUJhe6wVx1rs7KqKh7pX
O+5CHF3dwzi13RyGctdwqw==
`protect END_PROTECTED
