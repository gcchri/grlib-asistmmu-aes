`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zaBavTKVBwHVLg8vGkenpxzdf251Dy5YThuLdaW90fOX3HqQpFaVkA4degWvMno5
fXt6lZX08BPf4GkZs0szFSXS27aO3uREVz71MK2Zr0tNt4gHAVWBArHqhpZgt7uG
NmviJmJG2hDV9cC28eD4wpWgi823zcCv/8IVwk1tEqq5r6F06SfH/4VXDSRGZxSZ
Lf6n/O/rtYqB0MgS4Mh6Rjzw9JH9lUP/a0b1o+6B9s5nolsuEsAT7N3XLwt9HojV
UwyC7fvy98IbWrX7YC5EJmcFtapYp02qEDfa9TO+XgofNG6u+aTHc4nIO/eH0KU1
LnxK63zQiBdbATjuBNuTON7NeB3taOfUzQusyhLMYsf4otZ8y3JJoxSkWhLl6OjF
0KRJ6W6+KAaTpRAttQuvgTzlh7gHI9MudRXp9IU9Q2UMP8Acaiv4n5gU6CmtQsCi
MwPY9Vk340xVXLO34c31qg7G+e3c2Cuo3i2d4M/z5o8+SVzjsQFG0+WWLvmii36c
J8RbMcf2crnNOuXn1US44K5DtcWeCUix7bRu4e7LFUTsh3sS1CDW7DbxcnJxzTGL
l3vf7lIETDdXlgE39Fa3QcwSMh94RKcCUherVRBhEe8+r8d43sTPr9reAHbemFYa
H9F/eASGVETHWsgAPwQFBbDVZVG5/nNCEGt++M4faatvCs01QCOPDJaP1qd0HgEG
tVe8GmNqck3NwS3wn3lYhCIZTrL+EPKyruM0htwUm5J8StG3DUMOICkzS1CnGq9C
EUgLws33IPC8e1U3nsMdbUa6MOoy+NdKMmZn/rEvVPMIZnhHybB7i0Cg3yLTI7LG
1IZvOX6V3MuIsibeu+oKMJfeTgJzUN3n0fBMaBmBJ46wW9V+LxSdskrbsiVoi7l9
3OcrWliS+cNuTGc4JM5KZCNLqYjPVwIOiZA8sUD3YM4h1r6jmPB5kCa8V/vq7uI5
`protect END_PROTECTED
