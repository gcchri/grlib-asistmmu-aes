`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JQsxaISc8lxovjwBkmqY5cVKVyHEjSrlQABGxW3kvGTu/cuzeKMS7u8e5yUs6AW/
5jQz4lDyMTjkaslhoqv1T+NNi0i0bZavGm02dQj1Z1JfkgpCx+JYh3UoRUv14DdJ
uLh3PnPDo7pyJZ4Xqzka7oVszEj87P+9auYP3kZ2ij37v8i0sIK8WQp1esthEDND
vMgHbzwkdxQusF/isxeeD9w9Y4Suv2gWvYlgKa+rV+y7UQwfe2VUFj0IykhLG7/i
`protect END_PROTECTED
