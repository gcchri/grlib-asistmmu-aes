`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
urbCUaIfH9oxnuhRXrZedqw6Lbjjnd4VB/rJfpwBOE3amiZ3Ny42tL8nQT2M8P2N
ET7TBw74h4vQyGSdZAqhTBPlrG8Qr6n/NSsaxFTPcMSHKP4XblT8MEznGXJ01dwE
lpmTtsK3gP50zKvISSC8ESjy15OwVWpctqCxWkD/OTRVOuLCK1yzt4m+qavb2/8F
bfthQTrAMeGbDlxGyuBBidOckPFWOYvmwvydqyWCwI63uml5w+arML/PCNas3F1N
NHP87e1v2wBv8KZ+q7UuM0VzKSlHHLhATDdyc6fqaIYs/h/u0/Jem3q3ai21QV/B
MTmONJWqKTQ8iff1bK56T2Qf8iXZ4pq+2NdEQxj+F2v1GMNC19pkFvrd+k7Wrlrw
TeFiISqC9prk/TlILBGErwYdETIC554g2cVIjoknmWvRFI+KU4sWPrwXTe+R23lo
v6FxC/HVkNnWa2tfhPlOGT4aFCTgxUKEpdKNuhqpGz89FhCVw6AjZ5oyBlF5IEKz
yXLTX5lhjQLKR0wkhisVT4CkiZIWOJmsrYDtG0i0TtuJYlg33NBkXyWIWrHJxKa4
deoaxPp2tNu4z0wmtjRPjXonXVRP2kA/v3cU8tPpjvHP89rU0bNGhTzICjmEpjRz
zvgynvGrhrChHM1yCw48tKF59tgjr8x9RE0QT7wfdXsdTmPYCnUL18uWtLI6SodX
U7VO/UCaPA9oEajoeaMmJ16D1PqODP0YkNwXfIjkUoU4don7eAYUI09gTkFvhada
F4UW3zmopWcdH8xp++gCAl9tHVC80ExGOKdzpU72xAtAzNPcIEowCp/xEKM9Hpp0
o9TXObZk5ESK6x4mK5KEhGx2JEdm9kvYYRvvIakCP+k=
`protect END_PROTECTED
