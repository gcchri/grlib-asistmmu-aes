`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o/QMfuIYd52XOx9HCiWqwbWRm3p5z3YLXjNfpYibmlFNJIPX4LrxMQM4XHGpI3k/
6SioOrCaX0zzS4XsKYp3i6hdvZJxkOTU1p37tggTpfwYy8HLJq+mPwevQS3uDKP0
kCx8UYgHwef8AHgOr5mSg9phCOlPPDwDE3rQeXJ0Kq/H2eAduwIgHk470efClR7o
ZQgshUgJRUHLFjUnyaroidhl8lYOQl55u1YThRq+KORzw5wOiMKiWZJKBU5ZeU41
OmgSyQ1EiESsrDr/I4EW3XxbXivO9+SdNzlZ4C+W0PaCKF0rsd2x5R5f+JDewmOz
aYeduidiCg/2tdKwoE9gJ4b97go7/TdAr6aEdHABF1va9mIJcU+HoMTXCiiA48/1
xSxaucujNKL1z35WODBE7VeDVbLlMjAfRuZN8BYUeFEzCIPONFs3xDZsM4aDI9de
`protect END_PROTECTED
