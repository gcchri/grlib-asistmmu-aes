`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fqrjX1azds3s/r/j5UFKgp1xdKrVfnyxBxz0K0dpXbLURvs7evoCUgCc3UlP1jEF
9HnMLsWkn4lrA7LCoxA+jwOTcVQ8SyhV9YjJ9HsA7B24OJw+nl4Jvnk2OrG+pRWO
MZJEMRjuWbq7y0uG7a/v65TE9ig4oxvXkbg9LwLwW3PvJ7sbLGA3Sj+aEKAeZ7t5
FGzBRpfe1UZyAkQL77GnSOJKUOf7hU7Xd+SruGfDiXC2FLgevoq83iD4EEhkdKxJ
BYm3T+ItqRj990jpOw9cWwcmpIZSPcQ2zPGKu2ncKi0l7HXvZ9741oBU9i8oDb1r
FQnL4a3MFcatO69xuAS1xcHxJxEKkcwHN/IsmwGUkIKvGzey24IznisdB0GYF8eA
tSQl+ayEEIBoE3muOpWPOPCAbOo/vpcwQq55lp/a3lorvi2KiYpN7j9PTKiFNvgQ
7mm8nql9sPwedgvo5epWnvRjClHkhgwoE++5h/A1MIA=
`protect END_PROTECTED
