`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DyCGaE7m5/X1CwPkfmIKoskuE+KMNxuocQpC/EQveIl1S2ixx5ylanIJxvS5qCfE
NeGiKaOf+6a4UfgRER6xhUHhNLyQFR1XR+PoXZBLUT8PIy9obnNpbLNWxFrRfCw8
c5rK37VkJ0Qk2R7uW1qpi5XcQOIIOrpFfIwtqFwOjko8wzcw80WJ4VRi7ObDnryi
3S94aO6c3abbiMCAeaur1Nw47DCTUhO5DMBl8EFwDg4JyAi5empcSluLIGO0wR0F
wOSbCUj+4sgquxblENClxy/UJPfCWZd5jIHrnQlj6Xm+8HNtt8zsR34RR4BG4LIr
geojPrCIsrs0Oz5DuoLPCZUz8XR+y676Enz9PlPX84QyuntD+imgAz4SkGWN6nqp
oOBb0yH14nsxyh1eC4Ul5ikatMi3MbYB2Xxa10mc4rEgrmnizSdIwcdhW4zy/DWK
uTO3kg85qyhZt82pf2+eZOvunZflvdHy19RZNJBnwCxAYf7bRIR+WWx5Y3M7cAtP
`protect END_PROTECTED
