`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sM+PV8kSw8JdsfNHpNhrjH4OC+rbTvr0X7H5bQ72CD7I2qQoKpyaTjywlojejoKa
vNxP1IP17qYjLy7gxisSy6uRKFzdaQqr87a4ZKSBGlUiHiAUtOygRUeXxcuLWWC5
9wj4TP52iE8kE5QAFv+1WQKqTnSvAHWbEj3yHEZahm6dJljkymFP3JYna31Yv8vG
VF3xwZ/ar9ssBOicqTrKdlKHcjchbexmRvRsITkFRLOZK4rWTwVKDsYcmi3u5L03
vjLczrNuyBRyO1ApzDvvaDHRiYfVYIz6aJ/9Pjo21qqWiNZ9IGLxMRcmcNN4WtK3
OSVXfDWxeUg7TUFghGLJaCY5TndT6SkDkKmzrSNPXLj7OkAzVI48WC02Fu5Punoy
8fYhfB2ZEhWKEUxIVSvX0sv1FfHAlr01yXGAB8kKhSp6YdvInPESL4KzNq17a/Vg
J9D9BUmBkKoXEsVCC+yL7TgG8+DGwPMxcs+CAf4CCL7fRqLBVlUrU0uyXgjrpjeo
3ZgLagmIZ1oj4BP74sAUGHq22wqHFtxoRxSytvtfixOn2Danx9ChQ4HeOEztZVwB
fKc/Nl8OVp1vE3xiOjGX4k8SwrdD1ujJC67ZAssVqpGzVY6ChLehe3z1vc8nD5dy
LL02seaCVgwrMs/SOjcnW3FSNkDTePrGtfUExhgajDWMhI1lsPM9fsM2r9abxcrz
2z7rF5Us5Oe5vhgySQZXv8YWkLZ2tMhZYR0BZEKWf2G4+KYtvjlT7TAGvWcjiV0f
t8iKCCfV0aCvoALCcHyxAxbbi1JwVlb6X0iHYREm1ZFHiONQ1bgZ/KsaBCPrJdix
+xwZ6iMjAtG+xntet6MzWVpXXV+uH60840pGSlobZQ2m1gaKYsA8/PYzG4p52UMB
NhoPBt4VI3rh1v2gOqfirpCdgw6ZfiDL4SoIuulVAODP4vkWuNAToDu2vExZVaG0
kQYqWzjGVE0dDFHYA1Tx1gUsDpU7/9qpxQvfGJuhALWIQJTCd43rtZR9K0LI7Kqa
DltnExRP/C3USHhfW3pvNbM/8zrJUmZyPCLwtpKHkTKRjXoZA/00OuJ5+eVJaXOT
HoDAYi5EImP/GOtryYsgUrZDls+VmjRWvNb3mRXZPGFp5m7weweakoq8YyIEDQyp
o8bOJPw33uKrD9JC56gwf3onGx6KBnKFxOAo9lHr/12j+kGo6F4ks0LmCrTBAh+S
lrdOTCmdXAxRjMYcpXZUgjq3CF97WniI6CnHP7kTqvOLBZUOLb5vK50vDe9gExsv
PzWtj4QpdpOlreJGtbeAIcqVcV8OTSLvKngdx5qbVbWwQ1I9qKh6xUwaKIlGi4hZ
L+L6hpENq585uuj3WriGX3snYpwpl6tWMWrlOD5O5eiOUgTV6zHeCey7MPm6YdPk
3ZY4R6ZXVlrcotjE5ctGvQ3DUaPrC7q5DDmnX/gxAQcS904Q8uxYpZuKdTJmQT1F
/Syrf/9rM8m2+cqTtZlJVtmHIFTq/t6hgx9EU89NhIowPTemsQ6UFFpbKsI9Dh7k
QD/8r0jFaC4kH8tF+WFPLFHEQXgsI6pfS5XHMPkY9+pSNZ+Q11GxN8lPBqIBBGuX
LFoxYsbmga8dZVLOlLYnnWjNPm2FvuUYCspmJY4ydqwzPfRxmopQWpOyzqTqXyA9
6tXwu3BAuUwGIJob6+sd4nLNmnbxxrRuO2z7kUgCcIa24s0U7HWn3FlflyPD3lBn
2Q9vPZj2Sslo4qWymaVdGoWAgXukN8eenaOBzXcwq8zH9ROWegjR+H0Yg5zeOJ3F
sJYPDo2pUb2layBpNhY8fZx5T6dJf37vsPisyQ5zEdEQ8VnqXVdHk9LoKORv8Rq5
dxnhsFqLUPRnZueqLANsA1ILHO/46HtKDQFP/M1biZhaEMqkq+4wQ+Ah77oB00mt
iz7zv8t7Cou7Xk9z8KKs4UmaId3+IAHGC7qz+OpmZq671IRqXl3HABqS0CUoMmwa
D6x+3+CZjy8KnbXFsJzkpxQ/YvEACzmwmy/IVKXwFYoD3u0da8RSoKGnfylszTcZ
+2ul3OHbi8luTSUP2kES339ujsqP4Bd2GYpia+tVDb7wsG9hCFxLDR5WjHt+PSm9
Fe+eOWHW8kjkXTNvJzVwxsXS50Y1leNmY6ntnkj+cXVVuE7l0CdpA/qh6O2Hi4We
zDm5jl8OPZM0e2RcjoYCAwvYFgr/VvywH7TrN56lranjMruQI48jBmx99zjUqU9d
O/4bOHzRESwHY5XjWlRsp8W3UmzTES15sF3SZ8OuYBOQ8IBCGzwnTM4huuzpoeTL
jMJ9FoxXujS/pMzH8CYKIMGbMk/zH6DX6GiyyWaJyyQ1WhC8nQg4CKvhKk9v7F8/
umB6yICtjW+7twGzzq/d2CeHFPKW5CQurk+gmmxNEX8Uzm/JAZGBK7Wn1y98RNR0
6E3aw3qnPogTZSxjTTiiUV17YbhS1kIGAMq78xk9Ihd1xWktk8TtVtyjX30OqseB
fa9ufhtnYVOTqBSuah6Ebv2PL8kD1ZHgGkZ9Tj059Q93dfYcVll4DgiOL8x+pY61
Ojo8EHVRkhRawuvZk5KHZlcm4uwfHD1T57sPj9lfP+xSfD2zUWqv3AuIc8lT7shF
7D1bEzvWvHrGSn6ioE2Ud/+NU8thB5K6It9TbBZsRkqMPdem94ZE61VzwPWopWPu
E3zJNUIfU1Z3bC0R0w/L3eXDRXSlEH5eh9wDa1p9FXQHTJBqPbI6GwvUqcdF/Jdz
RNt3UmK4SaRWJplX9c1uxRCkdbwkcEA84ebE12PDVx6CTLLwUI9VSW+wAQbYB+V2
0kayc+nQW4khJKHMIIVNd9B/Vtx+2VZkHrCLAQqaK7kLyZUf+ViK0Z+F4iamESA/
10+po9h8z40wurzRLk/lub1YuCjerdzzZNEhOJb8ZQITmQr8n96Tt+1iGdd/1HhD
AhpEPinNEr5f/TkwuoK42zzafv2IX3kcQEUfq+awdwF8vNOfMV3bj96aGvsRsRI3
TKiT/KyWqAhc1s7TFehkvViuDZPnQ7xkeLgr8HYABgah8jX0D0qXLu/pXKX4JT96
l80OLWmjbwGFhKKfGCkVyYXBBoAvhE0L1+5gz0uO18N0+pxcZ3+EfWDDHUaSXQe+
wljWD4w0+OOSjnaOxwcW6ZyvTxlg5QaRhhPoSOebYxwwmdZQFJ8t/gf7Nd5ACZYD
oLmbxiWZrFdpVTSzdHyEymj+2c1XZAxiUOrWpRhMqYm9gly+WADugxHTrmYK3A2z
FMHML5Zr0rYygPSUKy9mW6SzltCfW6kDrmczP2kxrKveM64yuqg9xjIVL2QrQKvd
lJC6pPynvq4eLqbB3lmfiKWx/K3+rPEgYxgnAWiyUH93v03pYvPRDROS5tSJNE3O
96QHf2HwpxZx5hy2Q3w3XrApW6IhT2ydna900uwqneM09XkVOhiqsjGbdg6dk5gn
reoemVfbX2KtRIlKWmul1nyLQEFZRbEwPaZ5MJzoZXZ9zj1KshRgRPjB9OD6XKlq
1/zNYOq2mS09suqlepcpKGcaIrLDfbO7IpGM0e8LIRuEUdtNzn1AGgf42PGLogeT
iL3gXbBy5k7vSiSKNRZtOGtgvW/Q9B+J9L1OQIBw/E+bwo/0U3RBr+O31IHm0bpg
FRNhHIBbk7qW7AvhtLO+Lzv49SyunZxWu0uDPKtPvTLouWEeQfwnZ0hHOuumQfJC
wp25MCIskcXttTmZiaINCyF9et0/evgkvt0oxP4sneT0WkxFZvTBNdvXVL4d5133
q7CYPvplzAKuBDxvKWIynk/LS+VyKXED7cPJIetd9hyJG8RENSdNoq/P8QAPEfnD
W66IcVNCkaQMA3Q9FT2rG3wPxcgxeLCbpt/u/UnOGwvVEBiEn1nrwG4OGZhO0FR3
H1k4fbBBgPvM15SAOggiaG2485tP5pMPzMhgYoNGEJXfqynMSlggmipGDN/YYwj8
oLq3u6HoevF1gMSK5A1mUAkdwufPKwW/V6Pj7jsulDXT/0eZzfgzunH9todq1T0o
M4r4GvHhsjTRppRp3jG+uWJRpS91Kozp6AeeoJtkQYwyHSf8O/CL5PXO3Q3KRdmt
R5RZ6JqsE7QP/QrkHEHDWMFGHCdtlJv9EUItY74is4oikCVYLRaasyvAPFgCvomJ
HVqiKBTGe6zJxVOhRUN743CAk1nNEU537oQUX+tTp926PKLhbdrldCQyrc1obWyr
+s3ixl/Odt81vzHSJEyx1hpdMRc0oNe+Aqq2hUClYmiV1rnkirFIT4p46SxEsila
uYiWJlIXOu/Nnbj23TJdK1Cp1u9aLc+xHqt1GP7gLP2cRK86TXxfJx6mXplDZf+k
EPrfrZq/4xdB+YAMglxsEb7blDpRSxjlGkvI3OtbMrbc78Abs/TnihvR4a7FpU6H
sJh65sSYIhHLJyufYDKrxKxBTow7q+mbLYVXvbDPFJccX6umBJlZhKHotrxZkab3
7Ui9/eHbhYSxeWgSJQDI5mRpxDhVu//gwRYpUCcCyPlewt9uy2GW7v9+uEeMJnoU
ocUOUP414V51xAM3LQJQAf6+ukGbPqG1yViJrY7tvdVvZ3dVlvQPCp6x1/ry/1R/
hzbc43wWjMSSV2kW8hnL8KPJD7+feKEik/JxnE8n/xF8yWsi4mjDrN5agSpG3lgr
E19dZg/ydMMgQrJdo2Ll9yazAl1RguBJHwKlhQpB4cy+PlYLtLGoHKghMl9dx0sY
DXShIWuk91ekWYrp220LT/k8lUmAY4EUNP0zhB3mFPeKu5j6pfRVWmstYJAgBK1z
W/YRZQnJe38cM0hkPTRguAfSMEpgNCKRrR8Vbju4hQCrjAV58R7UI9BYNPOKEBUX
I+1bPEzuu439qQBUMK4Nldw5+Ji867Wlj+S42Y/2Urmio98qbBbcDMTsanxhyqaM
Vc2naVHrB62+ldHY5MuUs7ST6P94n1tn3ecFt0TqOrMHeU+EEVeDVEbmM7+jnVLv
AbjOl2mpw1Y9woTmt3crQlMcp1fAECd6DiuNA6lBHanBDB77v7Lw13FmIv4uNnsb
iMOu11FFhMBzjwI5mk9GaKk6Zw71eH+kdZPbC7hAGlC70QxskS/2gA3Ha7QQHJKm
nE29PQKoXx53/EJrZU8Lrhz/e+LFwzfD/2N5gcd7XU83P7TYxcpE2xETYR0oPzDL
8+2FQbbjLMJltib4rkkPKommFXrKJeBUrIj7WCPyM3hjOACwyQ+ryzbnl/GzPCY7
RGUKRCxfI1BBq49F8d+aQx1Y5Crc77zsw7XrMfRKRbpOFPSQa5bUrFJpaldxV3Ra
JizTx26BCd+lQzrl98sj2cYemLoQlJq7nasVnm2itNZaf1Tq+oYOdZC1PM20IEpq
N1Ce0mBqJlgz6Fc3sHq+Syc8tuokvt2NuYwr9Igt8BUtySwyO0dthnUCa+3hmT9s
6W7bCbMC6G4VfD9djmT06/vje9LXpVXuhhhgz7In2u1N3azX/3f9ICqX90F4z+MI
8/hTyD1hdywNU9c+76QGl9Q4uj5LB/rIXPklW+ibmBcxHso3NJ6cdkxeG87TUFI4
kR4B0uueEK/kzFucGObKBfcxUnpGHnmC/BkkZv+HKG0nI+ah/MDFxAHNSAezv6PS
YICLTlILSNOknLj8WP2Ie3ItdbmF6OUL2TZ3VPUM8we4MLlRUZdrY3idIY3gePXo
c9EaCzs9U168kTwss5TuiplAc7zT6HcYeXO+zPsoHePEA4F7vi46taouJLf8BNPw
1cpe4ryy66+kUb4VbMKlrZNJ8KiFXRaeSr1OP57wRQ2JSM1PcSwt4ZukxvO3hhjC
DQXpQnucl3qoo1Wj2TFPSf+mBavV2KvcCjXo3fM2dOk6M4Z2x3scX5P2EPBc9rzO
O9MPiMQvxMizo48Zf9xGNOg14tO1nFkVuzgLlWlxpsgVt0efjMzX6Ft+RF9eflmu
kGGkJH9kiZqsNSR4qdb8dHpYmcS9/SCThnRkT8ZLtbplotIotD7LRcH9iDUPutgM
7cs6aHamycdjm3HWTzFnacZzl3X6Wc6Q625Bfe/agowjbQBXj2kk/ZwlMrBzNUQt
bfVQVm4VRNmaxDp25rxsAKm4pHLDs7+9MMiL6b0a1iiw1NiQNBeFrIpwz1f+kiUX
lv8EQjCoefoe4XL+6HRSnsR8v3KDcmmhQP2Iilyj36UtoeU2w5SRl2JNmrMUOD33
E5JWr8U5CeH0C/MqoCLEEJU9JpO4vyzaJr7T96rswkowx2M30qXcOtZOIjvKMT/d
y4BdGUMx9kOgrRrHkuvK2B+1W7Hhkz7+9SkDgKCorFcKXpP60/7l6akKytbNZw3r
TDHIq8na7hBOO+NvEvXiUH2S6jjV7e81FBeYEJA9GCsFfzK+7rDQOb83FJvUX7ZF
n+1i0VlYn4asFKe3dY10dNycR1FUfpM9ZCgQ6SVYZDH6M5P7biaQNfqkFUb40kTz
C4QRTC0Rduiq9mK/q7L0MYo0TPvgaBnopsMwAcDunAlR9jePkrhpdjE3o1xRDHep
vDDJxr3oCLOwESfe3a+k6HAIZQYmSRVi5p09uT40hP/IDYHYOftQ7KqVZ6w3qzZ2
kO67hEZEBa0LQgaPLlLI9M+t4T00Rqh3JU5O4ZBOnSx5s7EQR0SPSl9rOjdzSV/b
famxq2fubPaRJ1yJOS3wAs6zZDy7zCl1biyDzwnFY0HnXKbRzQv1415nXzHjAUp6
8Wo7lPLhmKN3J4r4QV6elw0qcuTDBwZ/ZIDL1HBMPgGcmo2J6UyL7VzJPJUPwQEI
Wt97NLzAcvnwLGKDDmmB1QIR1xkQmWpLdk/LAyPbP63+y/1BWRLoeCRY7rGMbgVC
eSWCLJcOclZVGs3nRStvCZHHJ1fc2flzPjLdrPPMy8+HeWCmSGuFVmTuRjHUvp/m
AbVA7WKUbqnc6wIsI5aUL/UeSDsqd31ScA4kM0WvHMP7rANdosOCwHem0wuYaRx8
Lp4m3dVWiAprw8kpmIp88ex/bpacg+7mi3E6JyukgtmwTPQVITSTMhqS6zKiBhvX
YIel9Gk+/U0g4WhFZCOQ7JRopj+axABJZCLqthzmtQubuMP/G783j37KkfyHMeiz
v9UY6FrDsLJFlgj0e9cccD74a7Z+AdoiV5JicQ4Z9+Z/DsNDXVRofu/q2B+kX0a/
oGYpnmOZ2NOeXRu7cjBUOsnGqcmA2c9slN0hC/k24rQdUjKTXxmWeSdiJi1sQBph
8dwLQuTbwsGJFiZLTFUAX1iDXJYoHuWK+tuvpxGSqNG/B4cxzHQajQy9fSFGM5OW
u6F85x2IQztq9VPGo/g42WgprBUgxsLPidt/4lbRa9J15i+qvJo7JWxQH0kbdtIg
OWRsr2qwWwn0ebx/AOjtQ5Ditmak8admrufwMszOJiBHSkLvhh56VH4eZiIr444m
kAPA8TgqwmqA8xzWxJsy8vQJj8pEH9FIUj1SiA9/LqjRFpclbHP+nrMlBCaqJBKR
s0OS4Tn7bEmdE1/IDUboqBCkgA9iOjLqrjL2yPEtbsxipmYeik1lfXSbTzZAscCy
f8Ik7BOoMCM0fhDpLHo5711nROi93Pje0mdkUclkYJNvr/7ovExFk/NKLywLI0XY
QAG6yE/x4BMKl9uI9SrrkCVrX9p8uQuTb0/LQdLyMU5lToFKskB5hCFfi52pHlUo
aJBdvZEAh1WnvLRyycU19hpYCjzfYj3om/Va0rXHZdlY8+QmUYmS7vI+9KCjB69h
Q3EWJOmlPLua84Qk0MKpo0KqP1S0t+deu/FOGmTnkyzjaFRl1wLQkHsASNVPFi4r
ZeeOuBkvOsarN8bOBhUEIRopMhM59gY+kNonOF8dO6puVxZChbAOdNqipeiOK1Wh
FHsB5QmJzcj0kwI78q1a+JS8q6zkNntb0TjzjgJgSo9lD0KmM8WeJmJM7QY2h5sf
YZCD7FTEZGuY8lkcQ3oTTDZkWGjQaeTaee6tZQ4WMXXhPSgxn7075ezm6rHXDbW2
HVMFEHhdG8irfk/MGe6T5cDJE3OnSaXfbsoZpgKVKG2DzeVm5bZfHGFBQ6My/Yff
F9KkQtBVE0qeJtlgxKdxpOBu723rlw+0zomMlacRPVeEqdPJesYlnKl1NHCV2rWa
wa716mF4K8EoYJ8WXBPsVGBtIocKPcTGOfzKMdaRM+p1DrdxR/vAb1EBM5ymd3sB
eO5hNP5uVc3eijohYpHEYKGoWKphqfUkY3nE3sj3ZLfduwx4bCWZo9EWJRVRJ/px
GcvCC8B2eEaGfaf2Oc0le5jZthPxR7D1Ht99+8EamIVP/1wR0AfqrleyLlB35D8U
cTAcfi0kNO9SXl835FPca//ef/8uhGeyWgYQ4+TA3l4rESZH3CDErGMyZA2h7pct
gMnZM6D3KXjhRn2ZYdI3kciClayoZK88dkJYpwMSz3WUkyRVfhQgwmlstpoUgZ9B
TNMg09GTWBQB7JjgbsPF1SDR+kzxmOcy/1FcramD6RGgpKpT6AqJuhFg8p9kW3Ut
2DDvIhPXjvM1U7gQ4TxHN9H/Isex9PZ67PtllfirMWvhu1tsop3RgicGt4Gg3sAO
39vLaCnBZAkmN+oNHo+9KUcJfySfFg0xoM8cSYEX3UT0+0r5mhKGG0nrJzOWX1xu
nQ54P7nSxGohfyjvuAzom3aO4qxd8pH1UIULQKxgjvenqgtk8TdsXhkOZz88Yoc/
22YuV2KUKexyP4UKllChW2LTPtfz+zUA5jvtLbqVBVOSIbM8vcIlwrBQ0dhybl+s
FfUAqLL2f6+IqMqZRoe7hWNWzwidBqIcukDA/imTkL6aVuBOUgWxfHd8VGXcVKuL
SNBUb+En0Y0WzarL/89t3sUa/nf66lxH0Bk+Ru2DTBE8searee4Sq6E9Dkkp4KE6
rn9GAhbnVqO65EHh07jRXxqVYmSwjG3vFRyafhFRFgpP4P47b7TqRCv+hamZxW5N
D5Js8P4nw325qLGAkvUo0EsWHL6W1yhnS6RhX6WzukwPdTaA7f6H9FLeDHAyU8FQ
J9eUOg9PxZZj5k9X1XEEeg1bv6YY0QGph3n0F5VdQCQmFc3UCZcJI/psEQOki0k9
qq9cANkhd5vSGH+qz0rAwTPTtzhiamwnaaUg1LK7cvPjnv1oasJKygnPjw7jDa1N
wqdxalikMjzfIsA8IMi+0AgHLXewQtcy6ClFnRieGqfmGTS36YxbaQ5bs20yDeYE
p1solRiMZE8lfq29hZIkXGqpjGSZcdUDSBYjKmQZf9HnNgVO26ay39SJE0jed8nz
C1bhSOMzkf/LwQgzWMkXG1ZSy62OX/cV+JZ1PWL+iRZavX+GZqIExBXGNhZBiOl7
+660LI+Jiivk1MfcuWYzAcBXJVdhLJ9g2Vy85BqQoksfykJVcNOm7Bgnwj/Tys4o
SsefHv7LviI9C0PbzWGnVfxt9PMvxrvd4jXQmokWSNT9qz9PgKl4jMz+WIdTvRb/
i9UVI4TnjGXzyScdQ06tuRHqByGPV85oIVSa3e2ZLEOLVT5hgxlZKfG4mk7VntfK
DlQxJNLvdClZ8yIHf93X4nLVZKwrSWKk7/r+hc5CH+Y2BRqamY3u4Adoc4/RM22M
nLI0VQjDTjAB8YRKpBsmg8EGsaDWcXsslO3pBR8sA3qb3xpOfWzzfrXA9M3IJ6Hx
7UGKEcOGbrrnI/Mx8s8MufvUQMiebzozg+IdBWz9vNJlr0OVTE/GCY0KR1+UiR/h
B2if+DP5KgmGdF6o3ts+4XuAL66p3Gz317Jon1EuBjm45JsF7jK/WFPt1jDp0G3V
q3C0nTzPylzRdgcTg9oWRUquT/UGKpH6dqAbwxCrNRrzXiWE/fOZi7snZ8ClFc4X
SltXPEHmE+66X2OtmxiT0ojCtYW8/Nj2yVpH/1D/5paXMK5ltyy755Xk2A4vuPLN
wiI57TGCNFL1usVDaWf7Nb6ZfcGqnslX54fBK6JsrsKpzxDN8UzOnfDEIhGr94eP
boIPnFgn+v+k1bfIBUAHGETIF++F0ugELN7C76gx0eGxVvy1wyy18EOkzUkphWyx
KmZqn2KlboEBoN0WVJJPpl/3vE7qReQphTMr44yhGnt1iZeo3LuPYKoHuFPEdQ43
BF6hztD3jYTkLaBkTKwef86+qsBSNdBAha1YoOvcQ0msK+1czYxLx8+KDtQd5rwZ
l9gvqSwzAnkrzScm8g1praCiHiV6PmlcPBkJ9jPa59I3mSi7WkZGQhxFZOq7It3h
xLiQYnZV7OWh0bEsUS3CX96drL3Hf2uHsd/uEMtMZ3EDdK7Rgp26DCmgXFuLpdVv
vxr5/lgPI3XeZinK/WRmOgRlppsjaWFtwG9JuQltLLl+AjJ8tT9d0bRgV597pft/
P6P4+vma9dNMZCBNuiZawHey/go0Jn3Wh4Nrdlc37VKelxfHSr0VfD2iemq3jlsG
7HkY4LTpmhIDH3iHNAJLZSvrLfQqAqmdZSBTB3jINvr0LhRwfAx9PBw4w2F50vqF
gH1LdrstHku1Cw+2VpQ7ViJBo2Md0ex8rlOD0AYGEZ8Tt/KOs4aC3ds2t/oY9I4O
W3Fk8rjgVoLKIlz1+kNZ1GAO/TiCuTgIu0ASmz0NwVcxQZ7CYgzYqLcrhoGHYNfX
PILIrbxorlY5yUHa33ld6AKxzR312Y4/TgzDnAvrhTGfYJywhJkqauAb6KfTCgsV
maCupYF2KjZ9A2nGXrNU7Lxx5KdkF/C5mxoBDEGwgOpno2pH9+M1PHEMlZCCvAAL
HwdPNYqqJKgjM332FFyuVYQ20YWE6aoZ0Puy0UjhxvK6KUhqP4cEuVQiHqv4HxSn
afcXiXCPUEnc9USMo5+qu6ZF2PTpjJAexbcxju3J0kQJ+tPh4H/5jJhU7VDjgAFM
G5zjk8t75FVTHUUtvLKv3Y0m5C1uMItgbqz3eG/CjqaSyhMNGedUcdU19M/dFv52
7O/H2hAcFuajj8cSNI+LPn30EcVIpv4+91/wDH1PEe/zc7uSul3lKv1LVAmBEB/t
9kgnwe/DmDpnsWdE/vUhTEUiJMM3GziH6v5mpPpZ62x1ML4lhvmIeaNHK0xFSpIU
ZiJJfWPcaxbtFn9jy/6SKofimFBTZqAo7cONe2p+XMniu9Bik4YhT5AHMNRL4UEe
hkFwL7SjNB9UNYr8jIZ49O0GR+nfC96ghpy8qZ37jdC14P+obqf1st65TiXTiNTG
yhzj9Qh0KS8pJykbkYjthc0ScKQ9CnsRjxefSUTpygrSqhZHb2NTXeg1Q5MpGdA+
JMZ3xVuBswT4nw+MK7yHuAP7ULIFO7Tw4k07VSP311VwX1sxpSCuWskhigVA+VHR
WsanygXsu2lljua4gQycswBQ/RjSj7BC7ko5O/Q6MLtQaU3ed+MoMFdjkq0i3oEj
cZcfD99LjBmyhuCPd93D52cO4VVrl2YZhiIS0D6XaZf695Bm+cJI8Xl996Kq8PgG
hTYRmFupPZwpdXOModsnsfZtrUhYFxODQPFpPuid7NGSuj0Q2AhtqZhJ9wZ8ap5h
1WH2EtHO4tlfuW6FdPYWQeesWwBH8M5HLUZWKaRiHHqflYOfuL8jZzLgJo3jdpn0
R78HrhgoHF/wk/Jf4cbXyyxaWnXDADrbb/LLOZRHyjbr0ZoaM7sF1d6iJM/2gNof
ldAuTIx3qawPMNhhZa7+c4w56Ow2agK8f2YeUuXJ8n0BKEsjnkrW23N57Hg0vInQ
g5Wo6gNpQwJJg5b7KJPmujE4f7OjNx2N0m56GP8ZRSBtsHev5Wg3SxbNAChptSTO
mVi492T5BVkGBazX2G62xI1769M012WuQqMmCEhRIjmm026t5YCRV7dhNZuzCn4F
l5g1gWiBvjoYDYrrf4aPsVjQXsKI+TSLOsNU20F1d0muxV7lIBuaUNtJ24WGnal0
o90dqaQo0vpebDUEUM0uokIkGT/ZnEZAp+jmapQyegheZ7TxuNK9nI4sBd9jNynu
dIzf0LLo/bvDTbT3WXUSSXdCSBuc/m3fULXpO225UnrYQQk1KVUrk7NNbmGWuWqH
ab982vlVU1zk8Qrxy0lbCVMQTozV6O2jPYk5uojAy0sIYGbuvFlsgPHXBIRPcsEg
AhvwcJuWt/WaT55ie0+z6Yi9A+3iI2oweppcSn8lk24urVm7cPnne0igk3RmX9Dg
xv6Qw4Tb8dLcUnenhlVVFB0fxQm1mCq/Hm8sIw0QuQqVekU7wvzmhr2pIVlYoNx+
OyMiIClPcJEwAMm/Hk/Y6YlY+83gqLjn+soBTLn3V5B5Sh69shpxC5hhEpWvyxEp
Kmhtdojm+WfcwEfUcrm5Fum3yrDfjxYFUy6qphuq39WYuxHmRvTeLrB0AlOOb5SF
LOyCLegU0ITWRgcXWhpeCllqwK9TpdA2MaHNzTF0LaUVuOxzejxpuyxzXgTTXiH6
s/ZIBJJHkogXnShS+IGbCVCYNWMDUAA9X6LI63ZSE/oMIO/JHXCXtUV3jUJ9VcIT
tMYguavHMIEiNyL0JjVRftXgd92exWtL/y39iSnHIsmwWchYv85DLY9If77IdPHb
BmHOEfzCG/q42J1u00y03kuZGptR5dMZ/6WCb1ssc8VIfEdKPeFubq5jNAaTQ/30
hZ05aI1mXB0x10LV/jHZNfAe+OiJlBdOZ7mUQqk54+u9iLK9e6Cvb0cMJN+VvsBR
1d66DzmwsnGyntAYVZ4go1vXWD7UW1VtcnRu4W63aKbDG1pcqXa7kO0pMbMRCdHY
wP7OZQcGjn10o+fnb6Aw8y/+1Aui5q36k2ql6RiJFLgqBa+7G2XKek24HsUI5u9V
NFVQlptu8bU226kLiBtSRUOOVQlxw1gJ3kvlT2DVbZsQui8T60GZSiFbZtVCo8UQ
76EaGpFrM3fH5vjsYBi1s8GJZBOSVGckDm3Rhgj/X+SedLP7SgErxiec9PKbkd2B
8XumQ6TNZwFoJC3S3CyZfuCi+RIEPEPwyuu6v+/RnBAJBQempmg2DNrvKHd1nANd
RETGFcTl9yz+r37LwVjrXQSipZYzTfgqY1iZpvypeJsx+zoqEuxZA+DnRVzDryn6
hF/Nre1kOXLf4cAXTp0DJEkCIfnggadv1W55AeYoM38cM6m890mTSiBfk6Euvul8
uK83inCgrMDeJFSbUW+x2PQLyYOBTeHNkJl/NwiBFBceilOr45loVhxm/kNuCW1O
H5aBiu70zuJV3Q/yRQeG511UPVAx9+Xe0Wl1UuXDIut2FGaZbx2zQdAjEOBvIyS8
KNOmafSnuk2p+UFxiQMMoXFlUlXl4hayHOIltOwZbyqrFP1emzkrgz4ZqQblXEbC
LU+Nf5L925NnErO8734GUj7XrUol6vxXge47/Hqz6lTGPv3VLW1XaUS9QDuzbpVl
sMuGJFzK1qNKDL6WiL2VZuZKyT/vH4k0WSr3NhFUrmVuykRYv6fULDdWW2YQK89D
yEu4J58EfIQUX0OHnTp9P4W3qGrib5B7ef5YhHPQSqus/UtRLE8l8ymYxFCE0fLb
VhtjEiR0UrVt+pLh8g3zqy3uvxVcR7l4eneQrT+ogdUzl91GxxVCju5TZ3TrhxM6
4Lr2xdbMk3aLWV1t9Nz1A8Cm/77jYeXG5pstf+kVbZIMqrBK7Gzohp2OiOTUIhoz
acykVA5uFZ+SAB2uPJ6c4Wxou4g8LZ3q6lr3itcQexrr6v9zPyQ9jSJvFLgQ9/MY
Ya8fPjY/1YZyBBS4rLMqmpGUTumJw/atkdyB/DOHKIwNHxSKWQsSAgk2YiWRMb+N
XwCMmBnsPk3f1JxiB9PjutMAkTzA6LA/jenoBwLfqCYzL+TGR/m/Pc/dCcLesr2c
qDAWfZ0HpIsTnq0gecvFiS7LwNGG4YvdVCaXuey6mBb4wVw1rDsuzHxjW7lPbUBM
UQBh6PtFyXXAOqqDYM8c5zpg1lDdBYHAMqqIzL6weG6dNGEk7NKhfycUXEUqxjuN
lBSpnLAmxEday4QdMaIouJ7tJt7ZPjDmLNZIyiYhGsjFwBFVdGk1v+pdJ+o60rXA
BQ1WHqjldXw+TBBYyZTyTBmPmKNqXLMKr5dABQhwBbnZIoHWwTecEOe73sMhRgBd
8eWXulF6mnMrtADLuRWYHnrdAsWjQwSK3jcfV6XBWZbvBVDf5YcY7LDfvi3uIw4R
GSlGwLSj0dSPxfD8gElQuK/kJOwO3VX1k0K+vgC76vYGNDu7kEpBjBr6cNuv/DUU
Qn2upsqDU0xQNDBuTSj2zfJom8gNYgxY9CyMY0PWUDU7rQ2a3hz5qNwlw2PsAPSn
8uMo8u+jOSdvT1QHrG76n4SCr2uEgh0fdrQOCG6tXdaYmcKHqYcjsajChgzXMo4A
/wPXd5ca9pgA7zryUkjoBPNcmG7HYnyt/psxIhivE2/dI6Ky3lNHAJhLxFIaSTa4
6Rlwfxw91WiW/a7VBPHDXX+8ol1aN8zds0keTotsMwbqZ1Z2Qoc3BHzMODp2Ttn+
uv1hkuM0f/m+BPtBin9XkEbQCZDCIGH3G2kx+hAdSXPzCvSfwiofRfUxP7AWFdag
4vQj97cqA3wIs6KPG+odnxAT2tRUDB+j6fzrIAxdfsgAGczCb3wE+kj+LzLm+Ktq
D5CJ4H/aP4Lkjjoy/Qu8VEWDuBA/rc/Vy3e0bXiYkY5iZxpwqsBv+8d9gHyjzBUs
AjnWa6DCNkcRhUDtPH7N9oN9jv3yqfvgJI64fzw3Q8A+/2cLIux3zUchuCde/VJb
Szvga9IaPhWqx0IMLJhGgGNvaQjUtjPTWMp7yOSULY1hqRpAC1U5/i4mgReAk8Ja
L4PRnWeArQh8G59VMa7G22ol7Cd6ayQAIjY/DIHN18yBMy38QeJXxGwbTLjjUsgf
CK0Hdlys/LK1ea/Us7LmZLRJ3CGVixlSOIlv1O8LwoeBKavA2FBEkwxXalQuwb6x
qFWYi6cZ+uXw7f7lGMwl4qN0kCpPciQJVXQ9NU1e4XYntGWNi2sJ36L8EHsusCGI
O6/GdyJFphhr9tX/terPNMvMdU9LCal+aePsv2neyTUjW6OjHomcgdaRlmHYJATw
Q2ylM0D8dwWuj4jt6XkiEVQoUX/XPhkuY6GHDIPy8FKQIzGzDcK1VqkU7WtRN+qG
2ijIt8HQX8vsFV9wj0EnzXXckKmt5BqfKRzLRWMts1I3lqxRDLXpD75DZwHujl/6
R00HOo6ptKA0gO8GFS0FIMcF5MuYsCAqxpAHd2x67w3SbhR+x3Kjj+d7yy1/wLlv
yByvkfWQXNWZRcAL0QRhkKupXg9iHOownGivUSvD1Pon0UFckarAmW4Q+uoH6Xx3
K7aGd6/gARe71M5PWqVVMMJahl+QOFP8RU3dxNflDyIzAqzes+MFzi4xePTB/3o8
lOTXCJ/f6R2na3//UW1wirO+OqJgEATkKUYphSNurqgrjal9CK6ton9nlwSXGz4R
u4yqHkRbqGVB/Kj09l7yzouClcO6NpTvqcfSqIAOu7cbNCs98sd0xsQXGoMoptSz
sTqgac/cdtJJYQOUBiIoP58/cr6fthZ+E+bUc4M5oG/du6NCKEbYal37X3arTgcJ
che+rMI9C9mJPZRP7SqS6psAYgcI9x9tv5uun4TFwMe72PlTagi+4HV4ylKc31LT
xob7zfaG/0do7KJhg+V1IA3ZHoykbNONiMbTk9RTa9Oup804YQPYY2wAbGtIe2Co
VaXPvDHGypAKMbI8TyWg3zePtoCyZIhjSAp+Q6uVqc8mm+uTCLd8xnGS/4z7zkBy
/3DsXi6/+iiB1lSuZWOEnJ0kbQ92iJdh+ut7U91ApNxf9D+u84QLMOBGThwjW2iv
0b4Tys7W8L8GPEsr+8EZMqa6JDNgvPGWiBFsxZUaD+00tsNPnLY3aDJdSOyP3XK2
lHjdgkacXy6WDgoLb9iCAFD/6NkBSY4pRMZAG6SKIM6SY7dHNnAFUa7jbqL3kRxH
mhOeJHCPkDjEPlM+v7PGwE9GVowm7qBJrlEkGRFFs6vISDlP6GCNvPU4sDFhxkS+
oMqKHCtAEAak11z2vU+yqxV5wi0sMNMsXSLyDhlPGVCferAF0uBTxfeEa0AaVSfL
CSnZuaILkzbqwx605ZtQUrF72h4fRRen5fWOR3a01Xlt1eqL3bYeouFDJ51TQpzm
+3USaqPaVe2fgjMtOKKEHJfhCQ9D/2qApGhBsQyC7wOrhN3ccJECTdcvV/7lj8rx
WQiuITcoo0SmX5lcz5GlEMkFAUcQdD5FuOema5H5gwnKvuKyvTnoEynbHnNDXFf4
sQq5vkqidfxJv20MsNAxEuiUJ98ASutuxqkekgeqClYmgg4qQ0BZ6s5ZKYVOavwC
/VTWrLfESJDjIJzt0byfrvKfyyrbrLy4THy0V/2sZeLQqGb6W8P35y4yFvFIoAYX
EYGaEmMkubPO5B7fNS5pvrB+3jHlVpQtuunEVtU60gD7j8lTdj69mckrjYJl7zFK
+I1pJdd7rzxrPLd6i1gQgHs2RCndiSi24qMiQKlQGUQ6hYt9CnVM+7WwqXPX/jTx
DiyhEiAIRXTwDfvKCJSb16tWSB3e1ZWt5pybLAI5wxsKXv1F6sjvL9eIDFpgjEJl
3LawkDET3QCX+oISjHZ+BLQqQHyJH9LxabX69LAYppiHLzFZdD+k0y10Q2PSmUJn
468lHCAtceS6ykMU4rqIls00m0F8RUuiBhi40qqfCALtYeR8hzfzeGZplRhEZfTN
XDruNFVkgY3uwgyOKAxg6e+RgUSPwD157UL0nr4/6x/rljS/U93meLq7oCit+uJU
pAGgBsqU0N6mC3AsZHS7QENlguKTiOVOfvvFFMTrBvN9DRssSEcUgjZIr+KLaBta
gxXclJUgaHFuEaWRLWDVaH1zWyyu+VBtliuO9Q8KC/XfWAQhs21AcUAAJrJAIiIL
wtogYPz9421dQ6xjKqQ9XyDXLZbDUghEnHvn05EBClW2Jr+w/dlQNMovZyhXlvGO
BAeZwK0K12mAgZvmMGiAp0hNcUNexkWid7KZrcc5y+sWQGzQWV/cfGvOZgwvNAC9
1K8blo9KbhHy/0R/arcY5Ns5Qkycf4nUfWBODxHJAug3l3ssR8/Y1cnVaoxR+Lno
jwWWJF5RIzyrIfrSWMcMCOaEdQ5yt4OZv4vynmtGqPk+Qk2FfSrtJFQ6JxcIbaVc
LHgTRWEdiAQ26lxGo3KJ9X8UlhBp65ZawSufa+Tpnj+9tmi/k0gy6wD/nkqjLHkI
WC/Er1SBcSZryp5pm0r9vKcMsEb0HltmeQq6rG/12CkaHYO1qkUp/8IsFdPoxXaq
4sk9LhxZYLYSE4rPTMAf9AUxN3ahyyVrpMBSaxDQtqBYsY+TdKpuGgmjCTwEyYSv
I2UhN8bVp9+WF97xO+HiVleam7kvyOZXM5Xw7mr/i4E8kPoILVbuhaHExAS6D8Zm
H8d044ja4BfqoTDwuG6/QOrlzjvL/JF/6z0em3YlWVYlU+HJg7zIO/kK+n2MRu1k
Hx+T7Z0K53AO63lcBUn8kn6Q9Rbr0NI3LPzwMUnZzOlfuKSzaKsTl8a/FN30morQ
5TPDjGGQbWcKMeeWdEkhmOSpwPijkXy2Jl3Ud4oX5ecliIFct5bB7y96WKFEn/bw
Qv3M2jnvTpCPft1wzMrzg6b4uOTA4eLTwb4MQ/xaKKpjdaqynzJa4gWVtF4OQ15u
oN+brXZoYLxxDfK9B9s+mitUW51rjUTqQ6sKgrd07tRFVpRL74Nny0NSf3amhz8Z
gYX7w/pwV7qEUztHgqrFey17kOq5yMOsT7INA11RJMjMky6KBLXJnuGbmJD3j0zw
DcFj2B00dMtxLk+oRPb9a4TUvKIv5Lqq8l4CqkadHFqdP5jQACwqMveQQCCUYy9S
arkzaNEcAHViX3ja1lMFSql3gy1x/5evp5EfxV230PeAXCXFedRASfhFPdmsG+Vm
2ilJh0w1i1+aejKU6khxtATJUG7du0YAEO6reQjvBzjaTCwCzWoHrSgjk0v0djrp
lv2isBugqjSYqM2uB0NCloUv6AXtIWIp+T1vJLFK72dFDZFvf2K7mR6HHR9qJGKn
HnQ+6kdRanxO06ISH0CcYs9qb7Jap3cgvEncXeqPkZ+A2MxaC90cd1dpj/jBQfUB
+1lNDtgW/xBqMHneWwzK5xwLNuSAdckr7uaepwZZuShxY9GKvjPPQu4N0yWydxII
CDWb7kFVsxrTx5BPC9ydiYeNhVQBkAt0TmUuIBFuYHCBoVeKbBd0nWz0VIt9kYgY
BziwkGMuXBmrrq997bbzpqel5Y2nBLPnfj3q5hKzMuRY3C9KNGeneoLEqYcd3wm6
DwKtyYh9YJxG4B6LNQsVM3m5v8u+dbl5OXeYsW6QIGi2Oxn+CEiM74yHNIpiKbCg
0XfsFIA4+6khN1aJRGbuhwCGhJ5ifm5GXemqo3bxu9zjwpJDYXm4AmnwTzNBFo3+
m4mROl7HKHx3QGa+wlyBDDtVi3yRayo3ju8tSuOcdAcfWS40tAOy0hFHYPd0azFo
+JSfcylbgWjaqndUZTQNV3kZHkMqoImzxArZIIxTr9pbCGmZVIKlhWeYVo+lw6Zo
op07AnJXP4bGhCKasP59lBzrJwMulmVaESOjFoP05h7oVTvvTeyDDeac/0UZx0aJ
GrPL03Y5jyOIfGHif9uT1Yq10RUGKMfQS1dXbN+NRw0UkuY/NCNq9etTcpDfJ2fL
katxBpMhDtbcZogbJwiuJg3GoPVmfgMlswTfSIRB01vgCrisFh2a/kFoFQhiRhH6
gkUcE96iBWY5JQJcPwX0uRVDD6MqaEsiNJw1iHp1nYwLgyugQqSva279NxyyH2At
ZhRIsPyAjT82i7vRGqHgqwPISv7q5MK7xypG9zwi89J3dmt/a150BenPaAidOsXU
mtJ5GJT2iQL4q+3qqn5vHO8i7bRui+I11UxHx9QbHoBrMejAIRffBORjuzOOKU6i
PuWku99/YHiR0UneGAOmlzNrbtlqKeMVmUFSlnZB9jHvcELul6tamHfewPPfOh/U
o0kOfiVRuomCJYW2kZhu4miSHYlG2Hq72tgmI6giWebSgPNsHvZ72FUAzkzXXDj/
qvPWOS+3I54YIKaS7utMeJ2ruST21LnRreSpS1LaBURHUOifJWqh7aM+6i3FY83j
SdBqVVwMYaT+nShQv5aBvJ4+jOHleVyhECMNZtb80K5nnS1ejYh767dtFDOJaL5G
Xed4kC8wYFXdDcUxOK7ytbEH/klrt08jIzgDLXnqGr8w3g6jHMIuTIu6e+IJ5FJ0
P4ug1ypZBkEVegYRH4RWBiC0DmCIRe24rnQ9oFppYBNonQeHwx4URPf/hET0AJTM
AbZ4v7vNgWg5lIauEtyksxX5KC4sDR2iAIxgmdCt6eW3DYOi6rZ5I9vPHY3d0Mqc
BKEZ6d8prWjLImrdvA1CtMTfQZg2oskeBHjy0lADGQtdw30rNGszeLWeayW7sEpA
8GqTESw+zQjLfITFreg0VPyppkTFor5HuYkbnDSTLfRWcKOOYeFqSff/g5DBbO/4
d24/D0QjAwNVDBSN2kUbP/h3sWIRDHUI7zOMV/pqIDgrdtRjU9wvD+wikRHUwgjY
rqxnzIloouCLWQCc34Fr+ujeR0LCskWuBZnMUjYdBB/6ifhFtNRfq5G6ZSCflA3k
vntrglsJMEaVtk8LiDhwq7VB9aYCKeV0manL0z4iuMz54qpu0KFzmrroARr2283s
2IKFZJ9olqCeiAw9lPs4UE1dquydZHfad6of1Oz16bzNzg2XC6XQQiWtZ91fUBzp
BCi3WwEWGcFih1Yaf4kDgeWvSnejAnZTd1ur+IbnJOz5cVpfM4v7CAklrTQ67Ne3
v8i7u9Z00FNa/8GaGiS4t8yt5rpLpgFZATRuk4PVAY9PY8rLNkrg6QnxXS3i1zFy
BK6rUdEBNKQaH/8Th72D8a3Qza2lEqnma5P/UDkdA+bnDEb7FWXRRZlZj9oEm4F1
yYPNEmJg3TPXNuoS48+MysewlkcbelRYo4w90lwBWsGNCE6jKdaMWIsqJ0sUcLkV
/4bMTMb7PkMBAsVTir8ZAemjpXYohPnQ+cc+ud4Ww1RtLqk1K0tjsIV8SuSDk3Dl
6NhHvH6XEcD+7+eiPrKezHhZLGu80gvr3m1O8AK/BmTeRmjQ7Wiu9Hy6AkdFAKbv
77sJXTC2uWx2NScVwINE47jhKccrxDFg3jE7MArd6PaIEBeOpJins9MJ4avKLeGJ
1RAGfKHUqxR9YD8MeGNulsWRdBT44KoFYYgeKBS96nlLDSo5Wtyfu6LNFymwahIC
R6M/wF3fOkoymUfbzTn1qN3qUMra4Fjf9ax8lFPLmBOV2w3PSu96GVxJOrZy/TTu
Yt7mXl/22hT8yopyzjHLLxJdY/l7dmaJPdwxHgrHNe6xQ10Lh7f76d4pRbxgz0RS
+1QfBwoGZtcGE43R51P+hA8U3DAbyJ65R2qnOIUQP3XdNL0bFR++TR9+zcEGCf9K
OhYy2ebQd8ag+KK80ck57AiBSGEY6+EnASaD7h08vjm6Sw7zdgRdDjlhr9Oo6Lz7
vSyNxULu2QRsNn7KpVfhRej6t+1U4iwJ3RoFA9pbjtpE5kTDoxoOsLdKM+nqJ9rm
QrXGHk+uIM3o8SHDnt5LT/U9NoZzn6QN2+XwwwmwGi/NAOMggSUGW2zL0QAJeNDi
fptiFa3Pm35td+olof2Zb8etxBHnlXXBArheNQt6At98ubMXPEZf9d27ZBUvzprY
oel64Pt8tlyAFYD+17zM4VKdzOtSd1TrBnVF2W7glAVUcIEyWxXPTUnFsUH3d07q
p/xApoFbmhNMNOxXKNgFqDBTXpftK16JEbaNXqJKF6RL0NaXPdhypqSmHRjY8amJ
J1+dzVUlITPQlt533F3cLCDXUyVbOSALimx+Fy0IriOo795WKmN/oUuZA8jeUi0V
cqGtsm8YNjcMSioX3QJiyf8GMw1+g6/Iyn8hFZQOKeTshbWPFiOI39V7+OaSmgmt
QzPPyeMoDRM6BPpl8Fv/B4leUwbQxqhhjkEze9/0CaLdjxmKRCA3ACw6qPGsbrh7
SIb6zqifeARauv93p+XyzpqwucfZB/9rKZefnbP6+QhT+IulPB5BbN2+yqDs564j
APgnt68frFDJ8cg53V47MRltVD0YPHYh7le+MLDICyAoa0KWySXIt5KwBrxtm52z
88Kb848ihMnXhrbnMg9yhNUhVL+WBvH5zAnHtYJcHC2W43N0Nv3jnfpZwgXV37rK
39kkHpB+KyuhsAYLEcmX7lFZh6GOqaRz7b9AOrdoeCWuOoEk6fdlmk+qiuOOwOmP
XyQ1I770w/UQTHAyfTFDfQ7yZqGCZDOWR6telVbomTRsaT//99iMyjFhHmIUU7sD
X3tWTC86B52mEii25OlVAQDftMVLpzrzr8D0gy+wTCNX27GANhU7oojCjLAaCob3
NItK4xCk39v4GW6kAzHwdasEjeR6H+u0wifXXV2qR6mTOysq7ZFFlraYe0ehw3fc
hR6BraCpjdwaOh+VONK6VQbX+s6r11HBcpMT5OZv/qVvLucER6IQjs4Y0RMrGHRS
6O0qUGK8WYzmxkSXO+gZH/u4SSLckJ//fEvGdbJVpW5jS8QVbqTuchuoV6mY6Ort
NHVyY3Ez7VDaTgjkxtZdGldB3aRZ7bhWuuqV2dCL60fBfelrSEaZP3Hh2RFfc71k
DxUHfg0qraLSFvm2Lu+9OJouBRn3/vYxd27OphpBMiMjgYS1/tc53p3yBZBmC8Qx
Wkl6KFKrd8CbRm9xO7xTDtzJgPt3g8d7QWcoULtp/a5Kp6ggWndg+u4TxVS0z65L
jiJg+T8sBjdiMGNE7r607g8gRZHHcPgA2JoCmPuUkDYCW5PdP7Kwtm1KRuEDDG72
A/2gRrhKSU7OaqWbIE4SZNBEyd2raxWwdkWQ020it4uYzGwb9eVo1E+I9JbuAalm
o+gP3ke0jVpmGr8MDk0wmFrTW8juatid5seD7rL44FG49vbPMJ2NY53gH+rw9sCZ
j6IftCzeEEMOmwr1UYg9ZWh1iUq2tez8oZ9FMs/68phvZr7x5+LaoKCOMV6eoziG
Vz9Kd3vgT3HjpFWbPaAvLjCI9RvUZTuR07nj6cvhG6lGSDG8g0o37Np/NfPg2T1x
VozGRtr5ezeAWvdfWUZwSSfdaaivRXK7rOUs2/4L59vDsSaH2aBPluGMcsiYyQKU
bJlzzhb/lR8UCLxzPcqOqK2DhidXvoXfFSIJAgX9lZ6RYykq/kPBV4/lVr+0feOt
yeVI1Mjr6YYYw/vzGvLmq01f+vUCVnv07KyxIwraTLzXnHbJmbwASWM7doZ5Uy6h
8XVOjF/YxiwPRM2a9cQsiM48kOU4iznVmmcXExLUbLjG8JxDY35aaFzmUH4Q2+pg
5U+G9jnTqU98DTcOOeV1WHFunq7L9BFJx6HaE7KRCx6op0pCkbPDFZHzFhDxEW+z
juUfwjA2Wt18Sgt3Hcg/mmW5S/JPJUdt4k6C4v4k83qVwP4UWJ0Nr9Wfb0i/ZtPL
kkAxWRRFev/DeqDRFB3AEs4dDrT8IHbnyKib4usPRH35M+/6ehE23spaZzYxR3A8
rmNvPK5BpmVrkXt4nPwRuiPs2AQDnTIXlXYnpfeEnzQ43KehhJ8y60xatJmL+Xy5
QfIDTj7WXGbMpj3PTxLzPI8y62AIAJFYNoz8Webh7t0+TZKVPFxCVLZVQ/sg54uy
4MQV4sJL6lHM2Pw4kgmtLYGwQtYdFpQentOjfqoPzQpRpPh8eAqov6NqnSuD6vwk
+iJifDd1EHU+py0Gmi+0usJSGvfEG3Z6bBCtezwxwjD5iCSu0g6Map/IyGKenMCQ
pNoQgEfo5KOQK09TWsprAzoAZytkM85lfdNKj6HsHuAyU6u8vx0WWSlwE+o5MHB2
rzZyHTi3enByX5mP72GZJx65HPmHvU43MIqUIAawnPxQX7Uih5z8AsardJqYX8S7
ot5j6h+dNumkktehslVE/T76SCMb5sGkzcfQ47EITTvz9O7GBBmVO46EH9PPty0E
9Aa//If3hY7NGWSEVr0wTaWPjkmeeQnlQG56gwrlk95oQYhKuarGYClTfytRJy78
PBCWLH/cI3s7mSd01qGucprpcK+34+f4Qdo4ua9iixOTHcuyVqiFMDmHUe+EIZdH
CzfnGRCVgKLSMSkp4Zwb2reOTGGXLPS+R1mYPkx3F46E8HLWPP0+AI7UscHHGMUR
ZdtpF8xAQWHZPbSs/MWJtr3bX9nbI6Xj0NvNlvIudONsQ5/ky9NMOXsb3+JwC3w9
McWtYD/diIgbUP5p85fTXp3LL9ehEWuOUT2NFuIDQoeNWo0oKDIvxo41p7JiDWOQ
WHkQYMjbTXTKFpRPil5ey+7iXAqOqWhUoph/wiD23ko3HL26+7b+rptEhnXF1VtP
1yK/P0sRrG+IIZn9HmnS3y8cmsYGMDidmkl1dswLXQdg26uh5w+PnW2k7wpNTLLZ
2MPm6FCGB/MhQnjZLViEMqHjyoZ+6Xm9P/pNy6++LD1pO1AzAxcdZDIqhnrNO8c+
NN/lP1vthVMPO8CjKxSbUKb0OTAyiMbjmnzRaO7GyYYLLW3tRSw/wZyBSm2IsH4y
pYIOC3E5ZDc7DcKrQhFx/cvAo0MO1tmmeHYTcQ4XcQv4/6TGKO5b93BcJ9vlcgau
zvBGOiRNhrFnYqp8iRuNQ3yShzj3G2azpiDTl9EI0GYQAeV94za3XiDFw/gsxq+W
WBQTkTQ6RYTN7pluc73ghHeNMgkx6RU8KwFt5ec0jG/K3llLOvaee8PcJwEZubUI
uzGDJgk+Ow3GEtE7yK1TyTlsARvUF5eb8tAgULLL732T+Hyui4XBbNsuLVo++69g
am3QOdRZUgpjaLuporywf6/0O8/rBBmmmKLv7Bq27hYDgI5oejgtt/D97JiH8eM5
OTH5YqV+0DjV73NpspyaWR+H2G7nsORnvT5ey3MXmuCGi8WezAeKEfrqTLN3si62
85jfNB9FVJIFhWDDeHY1HHF8jjqimmrH7DUFNn8KgvTcFsnAoanHaGYDQCxWYg/M
V6OQjG8XEynj+3n01bALyaTL+orblxz+WP8logQ67n60wCX3up4ri0rrUlFfMaWq
Z2vypPyqWy9tWWnzB/RPAYIpcOUMKPvdyNezzXEiu8ik1ebLP8cPpfXw5J/tot5u
JefKxjznSVqSYdiArC5D3auY+MRBoydVrIiLV/x+e1G78MspnwKD7rAyI6aGGovR
n4/pjmpGkBgpds6gCtNJHd0lTV1Qwaro7zuLTwtXxuyDU3I8N2XDfuvX3urMS6HU
zZ1S3g1aiGromS60SodbNp9TJsyYP4YDjlBL7cRXG6Hpa4rE4snzLYSuGR6eGylb
wQE6yMF8jj5Wlus9OaP10jC5CzBFFFaHVbaGIbvPcU2oV+n+r0ROHUGZcW0OpU9o
MtR5zCBZuuF4i0TrignJ7i79lo8V1UMlz3g3G0L47L1sDLpQDrCMEuoiGzEdJevD
KDi2ViCjDc/9Gnm3rwHjMqG42ZEWk1vmDe/qxaSFmIQFoAgLt/IrgX61x8105e4N
LBk5t1d84XWn51DgDXROfjhxjRxfXhK9qmQ/CzlWUHuG1Y6j4F3QWN6U1mij7M9q
eYPosLJCeSmuqemOJ8sHwUsJ/y5p8begJtv+mWM45Qnlimzwxn7F1oFqK2u99vpz
nlBLQtbjRFmScCW2i8Nk0Q47PvCaJ8JaeTdgH+j+ZAKA6j31VYjcsOy0v9kbUTtk
f4Vn4GIZXxqZUgjo/42qLgS3504/NqvTpMf349qfasmtK9VO953IcZGxWDk6h9Hg
yzV/yO+OsdFNuyi7gwWkj21Tx/5QwvWDrfhmGso4kANBPbEogZ3+BwXmzkk00tuY
Yk8+xsjL3n7SpuMINg5V8e58mqNp9DnofNTYU2pLs/V5ksUPrH/imqSx87zxw44Z
Iii6wEojjznXc+XcD7dJ6ucCEeKHgYtbQk2SvTz59x9MH/e3KflTcEKjIVbFnkE5
BO6kKwyjVwUDkjX0Y0u50TwOL3q+4KfVO8gxQRhNOhC4vHz91UmsLWniDKwYL/C4
rs0m5G643lKl3158uKoXsBVURSCPFgmRI0l2sH0360hd83Q0MyrdkKksVVGI2h15
dO+9W3pT/pk4JMW1YKxl1Echy9Mco2vcgn9F3NQvj03HiQ3jK98cdqIPtyUGqJtG
hbCNOg4PWOtDh/4sp7yOAx9Y77eUQPI6bylvESgcly6lFRIDgenZcLKRtjQceVif
N19SjwLvbKv2jGmJs7h8BcjfgqCN/6dU0NzAP/azkoxzdrWvYIuu9cpaUHKL+fTd
XvNCJU/CvWxryITmHwu2E3wI7Lratk5NCx8CjAQ/N0y9vIkSmDfy0gFdd8O9HuW2
KpKn13oN2M1wsJ90wZDQal2Ohvle3FTXvzBiQ4yF9TaLT0dA58xYIGsBjjppMir+
SJf2fL561mvkJN7i6fK3BP4HvXOd1hEbzWknghMdGQYq1xQJE/WrlqBr1jUWtyDD
KmB1Zx43TcW1iEp4FYHN8hSRQ/lnke7TKYLY6k5J1Uanfwn4WT1UZfalXocukxEx
++64qztC7RXWUBX0HadHJpwB0AYW7DhSkMg4J5BYXxkVS99pLqa/P6oJmsDG42Ck
4ArMmMLgYM6kAaH6yBQ2w+wJ3/IWwWD4vRVTnYjG2HYaNEb+n7VvOqk5uPujen2q
8BI4TmbnwyUpWIlpc6Wq/iKpXpTJyB1Dg2Fdrz5mIq0ddW3I1mPf7GOGIbagPc2p
2QFznyiT+MBiTgZmL3sDyEmnroWUb6IDEi35QLKjJgeheOBQDgWGX9jlk3ASCXWi
BB3DLp5t4Ev/K2GmW6h2FAC1SoSC58CGYLzjKaa0NjLfi7/Xnau/tvedvhE8ICyS
R3UA6sHtaD1rxMyWF8GWvvEFpEoTQ4qPx8FsVNFNabCnBh/TRnKwKjbzxhvp2Kkx
m6/BY5MFalbSImRNDfsAVs5AUseYZNaaon1qBjtCjiuJkQ72DtZpgBAX7IjMijKT
KQWLWt8/Gs+rCU68FRIKDv26jbuSgrW5W5OLVlI3VdxrglWkB2RfHeN1JI+wRkNu
+wLJpISaAYNJ0as2GmaW4nlmyXyIh6fSP/MX8p+YP88E3Xi7aGsK9ouUebd6srhh
UCHUwFttJ2hEW1w5nCZ/lN+aJ5sJ7ijT/UTzR5CDSpr3FkCxlMpFH9/UXWhQ6VXx
e0CO0VNyH4Z/+Q8YAxdRDxx2D8dNWkl7DaIPuSYLRN4XREqbOHxEGAJXG9h55E2j
M7nU1Yjy+9RB1DkIREnR0dewm7Uw+WmEASwcNrXFApvjyafLdNOmi/tnGnRLKTVC
SMXGgujasC3pt/42W612tLkvU7vh+DnISNB+QSTR9IAigPlphoFfbkt6WoQdYMV3
/eKLSOc05VfwCj3ESbpZ4HyNwLkjd2FxoZqVSS6jKA2iq2JEwlCaQXkOf5l10DG0
clw4Sj/uzkuoGnQOTXQgtbkObK9ubeBPYLh2/OwQ9hF/tsVuVkkNn0iHwXfEyY15
N04DthHxeb1BayBZjgzaZ/9M6kG229RIIMQ+3KJZ9edFXF2NYIViWIw/2BbOCWd9
oQaWwZiwzjxSUmQ5cuOvZThujVuJO75aPjAKuhe8IN0Omvtn2k9y3XBFVtqcqaa5
zi6v9u+Q/1xgXPgR0EpDNVLPspQ391roHLBvOgoUff6xZ5YMofAxflj2+g8SZ2m8
fbfUwU3VT7hTWgLeU4TiouSPNO9K7LzMmP/Bk1m388K/yDY6OTvQA+lyGRzURmc4
4gH7R7BtbhujRqvf514+KFcyMoWP5YvIyShldXSQ9DDE/TPOw2ytPk8AeRrO7wWs
ocOaa/e2w7kP7zXpCW45awB6OClnplOOwMrnSlGqtdNrHbg/ysaz2C2qA+tlc/aR
7OnF8hFYX0DSC9DtZfhnxxa14rb1bICa2+ojh66BTUmFzUsikZgp8e5u7w6/Ny+Z
A2hJAyv6kq/H7PMAfZnrzos5QSwMiKqCmoSO01zmP9wWkOQEBztTTqA3Esr7gybi
QqOfZtmyEag6+HNbvLABlss+dycgNpdu0eiDCgylF1fa0uoqouthiJjXNwNvSYYu
wLJUDlaTUis8xpSJzVV31iiXgIl4mRJrXseBMTVOprz+EziC+a6mF5YG/S9pSkSB
VBsokdo+T528ZYWTDmOgCKDUWJLlGF+CflH0JponG1HN4AhzZRc1xpd+KyjbpUVF
S+xo2DFbQ1NjZXXxmqxD4UAmwBaV6zmWwjcXhULwqjr3oOfbDNx/9s6LLSB3seaj
Eamte8MMDWYjQ9ZgXmU05u0zMR9FWHN6nP9zwm94vQhjdwZ0lCGf2myOamht1BL7
ppkQvxw9bvyF38Lg08jEdFuxyhAGok3Sspabh5Sex28W+i0AWoDxg/FTGObun4QY
oI2GZep3MhUEvXRFI8FOegvrtBAJOBtYEWE0qlMpYFBuCsBqEx0yyfDirXXp6sza
ybkyRnFxoFkpp7L/xu9kYPoELmkQKYo5fF+9cKGa7mVmC5GhFSURVHcrLiITxiFh
btN93CS4HWRIs2bN9QLLGVO1I6VpOCvrv33BZwmFxRZD/gWaKj0XtZttRb1RmPFA
GH9mQRTRPRBYEY92fI4lcu9jKdKLA/UHpYFnaYg4jJcmbdlbpEu3h1UC/zoLTWJ/
jXSPWAmQPkYls7jmut9MeIQPvSijAKCnHpqmj7w11dFs9wzbmxRmAIfodi65ckOH
b8w6ZVCCwmIyc8X+T9tZbDR6gjd81ZgZUVm/U5pFplHR22Ym7duQw4ADOqr+MseY
w2KZ4M23yi3EIc+PYVIIL+eQ2t+Qs1MwR63tGJYBDp99RjT+tqgy+XTIl/putii2
jvIUqhD7z1BP4h6p6cmB0GLMg4SYfzXTzdRqcIfqrDFoWtNsDV3/tOOmkmjBWLfo
Ej6+I/vQYJwUa1ZcWkkdL7GOdXj4ds476anOT+FEgANAwjmc9xTnpP6Yj6fRN3o1
xjQwN+wFTZd7QxEySF2K92BbGJWQGlVGEehNt2MMFKKESFAE+Rzd+gmIPbJcOd9M
WdzKbITDV5iD+36176gJX91W5w6KS9Cc9uim7BLNtN6CLNMwc2of5MJTLHTArsAU
YhzVsrCdzrwwdRV1VldJFF0lmMW4Q3KKG2aM+n2MiATV816oS7AtPYPDNwWkyoB+
K4IHvfz8JgkCynSutmRZPp5fAhavJ2M0nluoS9vBSpYhbqmpQGf3OI/kCsRN1zfi
ymM6MEw10zyrvkoQtTh2+HxK4fQBv3tFFwGRzXmHR9Gbjhchjvckt71sYjgMquQX
0/iQy4WlCv9l9E2XtPDcBPLmGUTxOpZlE7/OVc6RpwzXIaHFN+m4iIB4wbAVL63h
INgKdp00gkVZFHHy2Gq+vcJbzg0ZbQjohqTJtyyAV9GGp/1st48Sl0PKfvRaN1Dd
ov2NKlkGZLM4SLm612iev7jT8+S9F0sj+C5Tu/98kfDnaMmIXOOhVMuqSp2iUmlC
4pZUVNjZ0XfX+6M4szbVe2mQ9fwG/7JzBcz32jDSL/HQrfy/sf3SfMffmNj+LWRt
IPgWxrI/NRNXt/yxAL0NSWOyCLuAsKnhi1ZdTBmEURDrQQ14jYQhzTVaRW0hbSvP
PJHoZiFDJ9XD1wMkLSCnS0lcrhbQelyD16tClBQB/b8uhVO3NXRXByPbCGJhJ5aZ
4AamseTFvfIfwrGGrkA/uCE6XDkoMcW/QL+px065qoMJhNf/AAPJamGUWS4DAyh6
lPK2eF0O/9gLs6/k6U1xWsulSDu+YlT15WOvyRDdlra+X4n8xqsc4c3gwegXgSwL
CgA3enkG3oNVAGDqgHL4yKHhWaESzpw93m/K4WcAGiNxi3b+EXcyIrXrmw78sfQ8
HgkpcSfTHjtJHvXA5nKIXmRnkz5IHVtL1VUg9q1V7JpRIbuQc+JYFr+39GEwRmPo
yzDeDIB/Uz/eLsCKXzGQJhS0Koe+6bI4Ue+52h4Pd1lGnELJRQCwn6fTFJx02ZK/
NqE2/sJQPeGUI2IiiEqKAxacC5qTPm1hi+rxVIXuN/INaHYf7Dth7QHAIXMBMJj1
udX8DyKcN15kju3aUbdaTqP8fi/seeWdYx3K95Y3pwDOI+ougpfrH/h28kv3MiNC
HXqB+/4ZMP4HhZLi88fB7KJ9bHTfmr7HJ4qbz7dkF08RiSt8cV6mn+xVtRDDSI2+
U2NUR9qIOZLZRDgR1OPxPjvdx0Hby+Q5qy5aDMbTe1VGfWwnE53Q7KBT859bNHN5
u2YHlLEh6NBx2rYGYCpR4qGJYiNWYWdGH81rPMjbROVumVKyWtLTwg5H0ttPsbj1
vie4YwkI099UoHGJ9jm4CIpodi40SH+U6SGmbz/3szr4kA44Tj9+DZXZZv/9PI2R
0/p5j/Hb+wQEJpWczkDG0eTJ36GLkTbF89CVTikG1OOmjxwY2+GrjSVjZqwf0mwR
J3ZBpDshw51hvyr6VqwJUpycuw6ghLWvmOQeThPX28YbyhOlBXZXdSGCQLUrXj8n
O85WUFDsrYnLGzLeyikPcd15S8DA3ai7lhyV/X0yhJBsNN/PoWplgyW3nefdoxGy
7gTS2TGb6+h8t0BtGJiqB0o6zcVOAcDuUIejsoFasIam3Guu7R9XeKp9Gu7IxQ/g
kT606rzXFXjOkqwQRwQFnHqEG69cWvcV/OcOmK5FOGeorWYmeR5DSVt2y+eTvOrE
MZJK9Z3VGbpbhcNwX2HORcZ27Z/OxR080A2ujd3isZwsSLQ73EQTAwRBCwc6lDdL
+HrGy31obr90GcrXAteLufwD1G2Mp+scKrtKgxWUX75bdmUT+B5IkswIssr0yFgh
baIp0H8APCrahnZ5bZ+QL6G6tI+4fvf+fyindhLaSJ1o9mmFPHqbnI8ywCTU3R6K
MbI/3KAXKmwW/gWrk9KyURN+jlJO9Kn3dVjNFBHXibRiEDtdVSrXTrazjmHC6Xuo
nD1AEzDP+/lXT8f3PYOzRMvycvSxUrn6av1y+c5BnNtWFhdHlDSavwo3B/5lf15V
7jSgu7UpIYK7l3x9pkc1fRFSxVFS/9RPWe6Ua1Sknij1IacsSg1LgeP6MCoNT1zV
WcUu1OyCPqdsLhrdaU+8aeAI+iM+YttLdfw0f3gQ9aCW1Ajae7ib5AnLDga2nE0/
IkwRMgFyGRYsRVnEggRLuUaPqpQ7W4bIohjqlL1mleDPuZzS8WF1tLmoCH7vBxTe
8R8XYyeiijBnKvoEbotsApCWL159ESefzOSpf2Gff47lCVcxcVdHN0vVVxXk9p3z
r2S27UrsmOBsxBwQoNwxpAq7dyvgS2yL2/fTGy9GjcWRkbelxoNFVfgYbHq4fOvk
jMqLQGaQiu7Ii0U24IsTCuGf58EQuNbT/stqCxHCZCyCRQ0Rq5WQZStlnk50mvQ6
+wdBfwpQ7W+sm7erKg9TBxligOxnrhMzRF7qsCa2UdsGAKhG04EkwEuiWzh17CBA
mmRBUCnxm/AN3EcbythoC6/sUq8hwmCHcMPWJA+ZQf+kEywGE0ha6/NY3FD0/Pv0
NFbu1O+fm7rT7QjOJ0gAdqXnpbFbJywMVNxbykr/hBG2y00QJrgrIp4s97b5mP+z
Ks4jJ9/DwCWKj/Y7QbbiWyqMc7asYyzhviaqLRwHPKOfOBJfsKLAPGuB/sakSzEn
fvN5E/DXNHuSw4w8PUPDmOH3QQm6A6aUzTRcP/Rxa4hnokKrnyJguGlnONu7+sfQ
iNwkv/QCVb71sIVGMnSvTr2g0y35LlGDipEzi5jO7cXvUBYnlNikfcvEC+vfd/lV
ubWIPWutGMBA909OR9gwqsO7IiWkC7E9LpinavZ2egiviMOskhIJwM3kdMA9JOKX
OhFXdLM2twh/jJ851j2CpWITAvXbANZqRJxkzZlldCnKs0OtO/3kh7CYuXUwBHZp
Dqq48kc5bGYVGURWbVBrinaOSbrQQuIFUFr70Nc/lVA0B2NBGZvaVpv+uBFr4nZF
GkNbgHsLP9TAguoDuucxSdh8PYTrJRXlpXn6br75+59c82Qv2gWpNOC3jrSR5VMU
r+vOlfBNVD061cGWvENHlpPXuBkR6vKDMMOzDjTtYqmprvXDM6I21tQvR5Ru8yyd
bsNb5Q3CytKFDA1161knXpb3gWndEkwVBMEIWA1pUxT9yuGNmj9k/6Sjq9IkZh3T
FtAfFV0mwq3lfxBPwMH8p5aYfno1sbgq5jpymvaIhcYntgDu3oPF3R7VUrExRIMX
f7XNvqEIEPr8A1x2RUxzh29dfiv+ISHGbVrgzWyOzNYzZemnHSSOof4eiExCNtrr
PPGycOXEo0t4iIXSH9wm76Gtrdx8Ft2jyuy5KCq0urkXrzb5Y1z2MKq4Xacc7Ho/
/QkHGFNpJwt5nteB19byww8CohsuysMYhi8UG67gw1QiXM4K/+8oOV1ZMGsat0wX
2Anerd+fmRYBS76RRTxArhE9JoEuJQV2lMuXVhLcMrwX2SWpZzCGyAqn1Dcjpqum
VOTzzSfZv2FcMy9I/87EH9JWVUmLFRIvK9HjZP3wgwNFqBS/kDnmj6q3i6798XbB
j6yUitg0mDkbM3QJ+6jj/HxuV7jrplg+m3x6sfyFFNLsXsoWf+s+Fi4o4rCim2re
4iooEQi9Dm6EKjKiwhw2IaKPeeez6gawUTmzZoQAb4lzJtfpWh7ASDHvXTsWFtl7
RWAq3ruDb92GKB/L4LOj/ewOj+N4d6yoYL7VyZqT84gGZMfxC5NqiOFjeyLBueaF
x1C/3dVKjAzNzRr16ZX1Tg816BZ5F1ueFjLPR+zC2d51NLaDLcKEzxunNXVZlIKz
gAvEhBjY1ylg+f8u3MEAhw5qeNT2hqJy0eow3YtH2JXY14VyQZC56LQEGyM4XzXc
+Q4IDpFjr0FdiwOaXZ1IjOr9ROA36aU0Smo1qobTxzATryq7KK/O69K2MRi/U8nb
Y9YHoIU8R4CYQqWFv/+O5hH+Ked1W7AUZAxFrNfkSwCoIWdckHDiXlkkUnfz/5uI
T6Wdfa5/XjROMIACbH1VtcM9otSQL8lZ+s7jXmbeLeamj8KfKVk1209Ib2YlK/QK
72EBDnadaumBs970JIflu1SJPoTVpYTMFUwsMqaYvv1eMADmRcfbBR+jPPwzsRm7
GRRQiY2zuBIsnoOiV1mISVx3y2Ats0yVrCLxB+CLukRnaadnKISvphbDGaiVHvWu
j9xVjrgyuMqLcyQNnB//Y0L0oikKhSwJJ2xGwt2G5e6ve5oYsE6aDi47hYCBDzKU
ESCaiymbAc8eNplb8zG1iKyhywVwg82rwVTQqjywrfEJSAcMZeSGq+vXAYhn+aFU
gRG5W/nkShrb8F55bd8fs2zmHFfzJrO/JzIbon3wa2J0cyNARphrh0VyxA2yx+nM
pF9ZB36lRCLUXsU9n0DWhkcT5/XNhTynqDmGaBNjHkeWBcdhsPSNsJGmk5u94SNp
2KoE6vyWFcNkZ2fDyo7N8cHkhOhg/N6f57oE/9Z+ePVbjeLW03HXj7OfVJRutJcl
wXLxBY2ujCd5BSmEM2HtUJ629sdvnvc4xuUt1laEhNP0518L24N3qrXwJ3AS4UH7
KwvxSE4gnzyHsO8KsY3wbhuJiR/3A1UDxC3UG/z3lPb1oummQpXnHPrXU7dfoU0o
JLf6SLBlqIEPfP0supRBrYhAQ2P5NJtbi4W+rhwN7+rBiROAlF+0LlsUIyfxt51t
F6nDbE5JrYK1tdYudHqZoP7PMx4+pzJ7VXHahj3OAhizxEVIMOthEjIquoa4KUH+
6Do3JyF6IBt0Q5QHHoDDX1XoXST0j6hK9aM+eSrCm5braBN/JexwJUmUXhV2BrvN
eI/6TnLr4pqluWI+KzjyIi+jikiz3BZU04rv3sQvo2/mxLNFNTBQfcYryMIOaLer
FNlhNn1kq6tdVhEiHKvwaQKdJTnnk85Yz0CZkk06ndu5YvEbi4HpnLzasR6IMXZv
NdhAH7Evwf4nuSOiY+wBXGBQAFlV4vLJyGyH4yaql3xjf8vz3OvQW8Woy3ZH8xUr
nMQ55YxOICekLGX0+ZvSHCJsMCjvlLNaiPApZ3oLQm48knyabv5OCjkuMWxhAFeY
JrqdOpTniC0owNy7GHpqPuKb9jPjo6umM0oxaTVtFdVoDrw22RnO60UsdGVrB2ZY
JLdRRz+UXr/8rieWKCU1Ng+SeUNKaNMwQL+grtez7jCz2+NEhq4gTSS+8rdLFBeW
9fEAyqloNPqx7HK2JE92ggBlPpOAaNTaAziGM7LK58Bj2/eFm4OZg711e46ET/l6
J2n9MFwDTumVECw8z8iu28hYZHX3jy66HFiUggF2NbuXYau+GEsdAozvCYbVjDaM
qlVsaGu71pI9C0zYDerqKnMKxcASfBNPli9V9aQ2Yc4vZDwd5HW1QgOiMBg+jVLB
GZWC7JDTfSsnHJQUBEl79DzyW5rCttXWhdqvHqZZrzVhejqey5IyDjQzOVUDAlQF
Zg/1rFUfTrka0shQJT76ej9LhczccUbNIioERc9hxt/y+vkuPRyhz/9dIuidtRZB
fblAi8D9a7h+FvY5okdWaUJq43ZpHTHK7q5YK9EQqk9PyZdL7ApyxI8CUmkouSLb
S7KTKWX0K0uaw4edynrLGg8sdoIXoEjfVk0WhdVRrGoReQnJmH8hfv9Lhf3F5G9q
196ek76m+d9A6tV0VAzuLJJWJIMVh2mIa5aH7Bn3sAf/mn1XTE2huseK9yEp2SSM
wuSBTpL8zvsNHnWDMrYKWJuZdcdoU6cWcZw3gCd9z2ubvHv3/gQwXPc7QgLTRTTP
ynHqjdRuKekwRbNmnYe+tLGlG8jW5wc4WOKX7+AEVxzZ+GZ8UjkX5VKSWZUj1w0q
mQpo+Cp1ESGpi7ezGDIyxds68y448VMpO2qhGbl1aClrE7glBUihzg/vUetkpyG7
Hr9TRHV6G39Pg/s2p3R7D2TvPCaZtkLd6mYZBLJlhT7J6IElcIshrQuSMyLypDjZ
0UHBE9FyqYgkLhBnWBk4k19iNRgGnC0RnJjt+jqhV9YbeJ/NlVktaTYEP4M4Nvwj
PFS2N9OYDPsbV/+3wCWXyUmmaYMfdIP2vv9DPSlwjBq+503SH+pnxs5kC5+Gbvyg
rilDLzAuT/ofTXCtgKW42uT7SmdBgFjYYWwnJvjlNjUpzAwMQNyGrosnQZ+BBPHS
ToVAv6u9s8x3Pj1qW+AwYss5ULZDNVr/DzExOXStDQDZB6AviM2zfBLP73imIwQh
Ubm9x9RvfIKBaBvTOwJh2J6ct4hiK9XN7T8t896NqwB1ku1GeTRLADWIUJXEmDmk
MSe5y4CKF0TxNWLMnSEqP0ff2EIwjoDc1VKSx/VZ+wpPiwZQWejan5Q5zbMqIipt
qrnnx95ldQqixDJWWtLK0ZHsW0BxERSHEJEhZw6uguN8b0BTvc/cJVa7D2Ula1GM
h/K1Hre+xL40gaipPmCbTnKyqBtIEQaR2OBMP3Va44GrdrvNaZU8cf7v0rTP9a43
FnG8B7RGg+39Fpmfq4IwYc5t8hzxHcIivm3c5cMM8GMQ3KQiwx6WFEAUpdRevSxc
oUR4vqvcWlf+gVfFTx6KlBhXvGMuN7f7WLVZy6l8RSnTLPk0AlUbP18Y/k2dfTyG
G1rBBeL5mFcDVXG4xmNkue9d5Rm6CE/HA3rxEWBSyncwl06dHbGeRWymLxZTktI6
DEM+ONofESVc6t2pezqjtxeGvP4tJRr7JkVhn1gWjbgWeyaR0Sz7GdWNetgevHv3
WNFDAODzmPTpEtCqXFTcll4FruuAd34EZx6yqQw7BQ6i1KCByVIf15QcyXVIHdcJ
ydZDj2F+AIulrnrMLc0BswheCrxeXB0apa+lcaXVBVyU8pQz+yfSDu2zc+n0tQQ7
j6lwqqrupkRt87TN91AOv1AYj5abC8+b619AoCLphNTHrXar51sS3ZqbOboPugqi
K7KMtsTi4Aif4OZcmilxcXEle04Wn6BVwNFIHKSuEq2vvjUkbN5C52sRFdS3P7mT
Eq0WaklFspPqrESwMCkWMekfClVkYT1HewSBcn52T//6JBP/KT6TjBaQv3vbQS2z
/QvrMgkOZV2P6tTNuCSFhNyHWu58dZQCBvexLFnhPIoNnX6fNIG17o1dsCMEgGfA
l+3af/C8Nfh27a/BNsmP1Pr30nHynjBGFwn4UxNyDPvdbugLuUJI0/S+P/3YeVih
2qhiWXIB2DRXf7YUk1jZ0GQNkNogvfL8vM8Pg/BJpxHspoc2YQO5Hy8I9EpUNGSA
gYD+aO12y9Yxu3KU8GMOZLkR/0tWu0+PCUKaSQo9aSCtwY9ZNlfxg9ukp6fs+nwY
cdAp3cE/XXN8G2ZBrylfGv38WPJu+5W/67GvNoPGYnSaiMxnQ+KWpDamH2rfMOlT
3laYzjUEU4itenCnbFflQOuv6J4ZTnvXVoh6GI+SpBOL4jn/BIqnOivyMupWSDQy
C8BDNFHKt4iTqjbM8wJlLVUYR9tw7wEnRf82evSNfLmwJG5dDNYUmPf2JRx5/FiZ
F3My2N0B1O+E0ZfWnjBhMskzuWJj2s/awIzmqiesjjbXE1m2aNyuTcfRj4IIiNTh
WQYBz24xWcPAwgQHWpGnynksyw75yGuKhfa81gIG7DIcyYTX/n4N5zpMnx7FmwP3
n0ZtjUUqM78xKc1YPKoVtt/EiXJpcXvZM7zNM9Kcx6gPaB//0g64f+q8ONineMgG
0UP5ZlvOOAoviX0e5leCoO7d+wzE/jGzlHAFgFvEh6EkRbjhLSFgl82pp49tlBSk
Z94K4oeb3/OGFKT8+JYOg3Yigb5vAY1Lt5bLziIL3dU6oFZG8MzyImCrrudsHMhw
32g6NLeSSneOKxreOakMg9/r4NZqc6uODupxnDi2XSwFvDc1BdXqrxsB3SgdylyA
ayqvQIFYjiutPBklER1YWsa9YHVIC+Zxk2fkr085Oj9hZO3WmIV+bA7W18IQZL+2
7RKNk2AbLMn9ljHafmLovLQGrQy9OlM8N+yDqpWbYmnkEPni7fvLLHl1oQ18tFJx
4Ql9XgJjJKnkixas5Gr+CYIVKWHOg/9QerOazhtOMumFIplvqN9Lc2e8u9zDK4Qr
Nt1KwRNZ9+tznkLs2CTHrprSVo4OotjG+ZjGXH9fWdzuBHSbl3rUz5MUso6nuULp
fTy1eqrU+Ios9TsaxEH7emTUOp1R5TjhD0P9wubDARviXR4yNtTUdTzOmp/krCmD
5t7s4WvxkS9pF56eIS/x6/WMtVA0hpGd0DHowMsJBsJKabt2ahUFeMChBpcORuFt
iK5MEpP6Qwm7ng0oHeFUDSb/18nlejC6OMCHKJpHVamY5/93guDBKxfGLPO/JXqv
RKInX+EAflxo9YLq/uCo/nFmZMsKHyIKHG+jEEfl5PvtsKJRCLHq4NQIN2TNlmZL
LArcGtHQ2vhEvaphr7JMYMw/djx9gDZ6MdvT0NoGcFkbNibuXTMTl3ld0WkHLcE3
3O273unpJmz6xtesK8NFzufAkzuGfhPvRiHVuLrcZ82lsgkI7wyGvT240P+58+4X
dDXF9QaApMl3rUhB+vGzv68vkpOuV1/WJ0F0aedmdTQGmeF8nLEJUpPvWeh6bRxW
tjHKxjHdtPk9TLrQr96ko3eRSRxrwGnDaFKX4e+xAAtwU2Sw5ItnC69MTMeRdyS/
eLUb850sMF65PRlwPwTCPCkJL9QqX6OIXhM/S9aNeJ0AidmJSKFjzOi9bpVJQTt9
NfDQp91vJ5y7oiHt6l6ObNVhntUzlnOKhdBJDLz+JScpdFlVvt3JPPOpH3lWKWBl
3WKe/3gCB208H0Ti969neEjeCVeKNfwOm0MDW2nxPmEcve1RHwRKEe31JliqkBsR
8C3dOq5QOjoV5ZXgg6JmLlnWYrFsTOku7z/RqanLvxIhK7VE0w6FBydbLLBhl37a
IHCER0WHCdCXzpUxt++zdhP0NqfQ1YrslVkqMYwFAXe0c1h/0Qu4DpBrz/V3yP27
ANEJn1+AUc/Q510tGqdmPNP7h4squVa/yokgx14RuD/zcTYYLyKGyAVjRg1JVW1N
C0RKlp1xq1AMYs6hhOBSkzWiFH8Y64Ft9Vh4BPUKeEz6u2fLbaNCeFCGwyyvTmFN
kRdV30kCQCooWKUMpJtRDC143O6PPxzQP8WILlku2ZqbHCCS5OgMP5/OUL5qbD4z
FQ8eckmnxDwC93MLKI88YZUCHFlf1fI8xzbDoK+vrB6CkuGkA48GHB9lTfWjrT+4
af5Ndyqa4Ht2Zs1TshoCzb+ZJcXpO7d7VdDhgP1OcP/XL88AT5MI+W6Cdvoq4m72
jSF0YMPjeYoJ8R+BlqBZ6L0NgotM8Avg9bJ5UZTQNUTVd1eluwFfY5FmfIU+vvoz
dMQj/LbrSnjaYzrzz8mfxnc4F+V7dVfF3nr/hKxZOR3aACBOVa1Q7maCFqluWnw5
PzoCSlFgMm31PSk+WsKtIbJ1Ta7E+MURswM1WY49vxkeEhjS9AhBYNH7NlOyHkSr
JUrYiox+qAAdznlJPa79SxaRhaEg57UtJ5Dp6xBF+GHoOBji2mEmfMWt+sdx12wP
9rQxMi7xyo/0HQdlStb6vKmOYN92og4MKudAfaWsPesa0t/ih3L7FGZNkJyrbD92
O5anzz+dKFNFy0wsK7La3p2y5ddGtnOQCT6Ie9rirvUBhStMdjMJI8OQNTSJatS0
nXQ5+QUy8nFUBCrWMqcLlSAMGBypRCewuAKWxnWIuG+0smlSDdavTc2LFAO+x9dH
UDvOGsPx1kk18t03ZcoPpwk3JecBRrOVOtKLUZnOn3m6XIiLezuwwL7GQt7qlH/w
m29QKA1c+ITlZO1Be9UepKtPC7O09327sC48zt72lnDmAFbyPSqxraTDKIwgfVc2
KoA4jkrNWA35Qqcq0BmwnRxclnD97dhtVT3pjAfUXq2PILjypCLOrGikc1+apnb8
gnJ2ONAi0Dz3+iV7elSrkIdlV68wlHrD9GINeBzDeOSA8ilT3turOEK2Pvax87pO
JbMJtNkr3/crf5IK9mcfGFJelKIphGYz7Y402wBi5+wTnCrMrAqnRwANbTpiKbb4
zT+vsgqejhqlSjH11faHRhsx8ahoXt9qgBZWA7nZ1uP5GQPf/2OTtRCAfwnU+U/L
4C83ui/gAlJq3dfMiiK4pvGl5m05vUbkuJmmw7ghLp9iucte88H9Jf2qFyqwQWwW
NIv0ALwzEL/GMFJpKJTGLLVkpB+YDmT1mxNDwELtkBnQxh3u0U3jRTFQFOsTVOeQ
f4PeKltgRzDCQswZSG70M/+KIH849SkQ/Vr2Qk8owgf7YGMhOlPfmfFBwh6HmTRZ
ejeJpqFQbwPNbq3An7+5tAsDNIz/IGWBFESnppkUEdL5BjHrXYc7xUWVi+wNwtNx
bZy9D8jSPtMIH7xFLbR7zqjSfGdGKLYCAjY374v7MpKdJU7pxvJayBx3QANo6XI1
W2MgBy/DZeKeeT80n1D/fFmankKqebUwalRXuf+5OPz9vHib4Hzof7LxRCuCNueo
stYrNypqaGBy3QpYmqvjllQF19LOuG6VVmlekgbigEWplZN1diu2AnA3ZzVl6jeD
R7mvub7+9svJLdC2/uoMEYZkW9Lp7GVlFEBMvsohezyrFBowX4DSppaFK8JVfQxC
JegMEee/Llh3MXJRou09TX3VeEyNxYKKoZWNxG87FbD6Sum/MA6yJ+WvWSJLjNRQ
+9FvAam+h3Fcdr+qeCBwFZsl5O8gWZJLdTHw35QUZOZj/2bstip6yqAd+opBL8Jg
Fct/N7bRcvKTdQyH4/SekDsc73LekuVVKdrePm4mcaRahhsNhJ+5jRH8V7fwVSU3
/w/dd6qZSJ2Kpjv0j1fgOCEwim4a0qxa8fmcNr0Nb2RLg93hBro2DJW2AB1tymcH
5AVrmJ2fsP7wd9dTpzUJQxZ+IdruEWxXYmHJl6kK2aSeXrRxmh5hx4z0FYSHYjJ4
shqYBSiMstwB7auB2IUbykQEkb6G7Jp3P9R/OTiGs6N7sOQeAhRYnykaV8a5e9ml
LyGzZ/rbwY3s4eF/MwyvqUVK/BhnSDvscw7mV/9+Lj8gKpHmAxIbiuwcf76f1QOO
vub5HN2SCo1RkCeSakjnaFM+5Uf3FW2RQ+7ovMCainwwR0jaB31JO95Uie4M/1Ki
Poi7V/ZjbYpjIwSDqQyJBfCyF1T/mE8V2C0p8ox3w5K9AQgBmT7BdJm6totscGff
lsbGUbLJ9ANRopqhAsvfm/EN3YVUKW+6M6WKOLkhnHZxVDkYEJ4/u1YMfOBr4+G0
efjKGLfXBZYmFCxsiotE//RvMv4DFAIIa5fGsq8+pZHCDmYU9sLmgopzhUqvaYH/
JQ0LDZlIpyF8JKFtrB8aDeNFJp0DBc9vUFxjiV8+GZ87EVL1NNPUge3oKFPqezVi
M6rzZQM4peBtFgQ1mXkPU6S/SBwAqIRD8nu5KHOsW9Z+yuXq7hqQJymrzMnZ4dyL
3QL9SJMcZcrPfNFwI7w2QiKCNVC6zWElcO5AOOjlJ1SQuA0KR3au+hLoU6CKWxyr
qIh7JlmoGlptcHwKgYCphSwFl2lnzExQyzPSkM6r/27Da7Vnn2SvRm+ph0lMDctO
SDsTHyh+CmrpazPHYj6IXghmtXymc2oSVOSFUqcRv2UoEEJi7AbGg8wKTEZqx/I9
j4JXGfuUEVMMs/y4dHuTvHoaEbLB5KaSAtSwBOvLGeIliZwrAZzgQE9PM3EU7RCZ
IiIiL4g/ems5+ePVIw4Za7XiFa669fWTA6+YzlULn/Z4M9MpgsWDmiKSa9lFmDh/
RfE8mP7jqd/WSEWZlGxFs7C1cGbl2NDiwlZaKtn5Af9zXN8jW9dZIBWTHmOD4vQU
wePjf+BDiqzv3DIzD7yc4nojQvZAmRTDwOrhw84V00h19wsYQ/7LSXcLDiPi201B
hLS015XloAOoqx4Z17lx8JVGSW6WBmHy8wLVkMcDHA//MdSAmawgv5muvbAjonjM
X1d8mUoiVEF7PJYEvDcqCglLwYE9XdGZtF4GNUWYJj176XA58bSYJmY84sn92Ruh
aS2Z5C25brFjd6GBr/6Toc9KKoqWoWnplqTdgTHhpifVSyk3mRl/Dw7dt5Lm17oQ
9mBTkD1fSVuFH5uY/IK/Wo2ZCA2+hS94nIAagK9KAJw30sIMhxXI1r0sdREFl+1V
klLd5XeuIcYDL0RiGfASDgLYL4aItG1p5M3cF3sBtHYcGHodP792uGDjAFHsn+fN
LSBA26IoKMVWWKa7WF9IcjtWpIGcTPC4PizvLCEx8L0XFb25aQjdK84VmDnY2SSE
v77TSlTahsk+F08zjCB4BHOTnJe4ip7MR0o3UK4MHNL3DGL+21AgMlbD5SO5CxKE
ovGZ+CZMQBEoX90X5rihGHlu4FUMQPgFDw1Tw3vMX1ObqCIb/PRfRNVCy8Rnu9Mu
dyz6+c1Ux4O6I7IzZ1qtl6szMk61k3CyUd6QMgLLaS5bS0y1YQtRISszjqgmTZ5M
wL1QludBU0qizBEmmZz5D6T6FTnbcq+RiLessHMK3bIoLyt0wLMTj641wviRK0A8
3T4Ziaou18ryXojQldiY+0KKAa3KtSV/5DD9buQ1NtgKkxc0NFKwKs0B1SidH6XU
wXxjkh/qu4X/vvCAnd5uBCA0Nfhp9mU1rmljc3rPKssiqq2guctRriKiFRuqSDP8
SITon3/oIn6Bz/MOifQbrZYugzhoiZPNMzL3z3jll0CxeAWOHeM1QKMOhvjNnH4w
CXlaiKleTnswZalduby4ipojuH00L/qaH6OagWPjmLHJ7ZFgq0cLRVJVHDmEtu4E
DAVHANNUnFJYnOwhecUb6bRnJLUFF8tq02zty9VhdYRMh4d3MCCdniyDSuVU0m1E
BG9qKmF4KifzxBArAkqfuvXLCt6W/T6er4xgiUJIom1e7k7g5sWYi9pp+M/DrWq2
Pu3kyZ3YM5Iztfy27laJQ5CqEsvpGZs7awd+3rqGw28fQq2kQ11GlgvIi/AQJhCE
evobJR00o74YqOGR6LzlQ1rDDh2CzeIrTlkJi3tXhfMzlmp6BHRfuCsJyOoyAP0E
1ykwG5Dn1BeKsZ+ZBG+tcIm8/a7C3q+VSbIRe4b6mkqUs59A1AXSMvpOKMhkzCyO
p6/TW6MQ1t/5lG8nOReU8je/d3x4GjvOLT4tac4+biqBcdtOl9EwXnzRuZEzA81R
j3A1pC+WaTDkLeIn6f2efjgiNIhFxUHmoQFTcT9Kx9RvA1KTT+rcMBn8Lpkok+eU
rzc1IRgRB3VU6ufScMhqXc5LIU9rYFtEX20cVZK8NjWnSKRz9RCpk0rEE3qk788L
liWkbyjw7DDHD2nIblfvJHIN8/KSmNqhgzaaStwA0IznVrg5PlX/JyLE/GLgEn0b
xu0ar1mjUMw6aWKAG2OZumSnMK6jyNK+OGWDCr0NFjs/BUr1p5xWcXFicZrwSTt7
o5ysLoNkgPWApx6U4qY0j+VYwwZYSv81/o+LHu4i28JOd73qnNQETXZNv4KfUSvh
dB2hDOlT8gsxnoIUlsS8WezFF7dhC35b/h2FdBPG7+aIueZygBZxx+ynvGE2Xhsv
1LjoU2kPgR2AKbxw2XgQ4xxRsLOUdvrHZQx2N/1MqyTLSfNoJBnTNQT/TfI+HWNr
nbialN7ThnF+BhhEspDznYw5nfnOHIffcZVkaONx+EZmrRFmwYHg1XZnMZXEW5Xu
KLP0vFzDNGNlWcyCBm2FTW37qUCSl9cvkLVLHA1Bu1DLKQWc2rCRBna1G8PHpYi1
KJlaB97JhETE6nEjgxynnV7zI8b5048jk3GoNGwCxnjMHjmOTOPpgw5T78wFRcR8
G90hY6nAeV3KXqGgSo/ynEoOgpzaDL9uhDUvFkFpijgwfvn01hKFge0xlrBs0qj1
ckwfyEt/7agFfHUkc61VaE4608nuWCzpapFxAS7bTevLFkqteveBaHeOK76GzC1T
pkbHZLs0a6Lby0OIl7HtSKCJx3ne5HSKW+qFOHcuN/wEOT90RW2kydqiX/NjxRSH
AObXeVgH1ZxdJOW+kE9ahTtneZ0EcSR3wS95yM+1cObQQg8Y270hzZYQypEOMDS8
g2e3HLDg0YMe/jOGVUKTk4K5QIgkPvRAFG8qo8olg83Lm5eTgUNVlYODWm8GtO+1
3VposEjnuEzRnSgwimDkXps52LeGMoHD/U5Z2jexJI6NEYobJUQp+BzcQP89ZODf
jf8TiTEZaNAjlO4VqR7JgR9R9TORwHPYx2Wu1vMgc3rz6x8Q304PSlLCfAW7qwo8
aKdaVyWg/cZR/aFIFWJDHi6Q+CNQVhFgpV5Z8fPcFVIvTxmgTfRh754D5iqYv/AU
Fhsuc+N2vm2tPd+t9JJ2kNi9msBLo+nFK+p7moWal2tYTJAiaMy/KSKizOAeI4bw
WEHoWhh4Z61NsS6K5ZfZBdyyhX8UCj+1Bb4RiGxs2kXMgvu7vhbUe1jvF9TbjG3v
dlJ77qmB64RK+K61jVd1AIc+DsH2gtnE2hUu8irjeH1zuZ2IKzpi3w4lhxIjCZqp
+v7f16twgW56w0UD82SqlBlUUP7pMUpsqjztyntfkW2nMzPJa2seyJzDZqUwxQHY
e+dAMqnYPTWvX52eWEiKXoGKWgAILAI3o1jNlJt8jBY00PNeZxpTd2ef9rbUR5HF
L2gvqpwaWkolEHpVcsriqSmFBmeEkn0J9AF1N8BuwLy6faRgXYaN062UxAXQP+Oz
O90O6B3+JuGljx5wZdoWuWrHg3UHZ7bQOAvSBb1YtK0PmK0a+iKkF1+2bDDJZhMq
kT0Al4tO008e2bwryDX5+NGjYTzHRMwVr51E+ETwDZSRSEM1RKK3ejzx6s5ecwEK
uJ2HTl8euJBlH7woL3PHh46yzsC2DBE5n3VXP9tvxAapRAqR+4FAlBiX+r8GE4qE
X9QbzfDBvGpZCh1Cyv2hdxewSzlDYjhAs5lreLnbM2/jpsWOzUhB1HnWMmdtNC0v
Jn6pexT6OnKpnzxk2LsCqv/REyxvA1QNPyhx66A1917SdWxPLzBi4osJ2iJ41PPb
Br79l+9lNqP/8cB7/em82V9ehwzn6s8cSJm+1ZOeC4uM8fZdzkZQzXMIZ0dr0K99
GMO+2IKN64846EHOzlKMv/xXKOH4Hb1W15YWgI5LO+e5+6WYrrEqaPsn+90T7fYd
tKBZ8QH1qKvapVKe8iEvJLpLzro2m1aJuxGcbgsxdzEBRBQUrCOFeWJnDwvLTANB
pfFS1d62LJAHrLBfIYKveBw2M3etZp3PJH29QnLUNujD1g2sZsxp4JwUH0m32YSN
bAWZcaMqWDmjbBeOee/n+mEkP9UDsHb7J8MpNshnUl9YWadIMQZ73INb1V6MfHCP
ZaI3WH7u/co9aC3hfGe/VnG5FH7CHZe0HGo6SG8hyByeKVP7aAubysns0qTlJwM2
tq61G6QcoYVCPiXIPMo6XItecEmDnBEmrc5EM8NBk6k0gGlaEwyPBULP0MKXODJh
OM+B9ba1dNTCDNQiIR6T75WRPFym9AziJ7/D9Mzbybu/Jd6P7fuCL+wnMRUsnVFR
TYka8evNLMDk1i3pBh6mWbLmBoDYM7fCqDZTEZWZM1bpXdTBG1367cqwz7aGg1S5
BzFRE0mXvIUTnW2OlJclmzH6ID6lNX9/KfEKDPOVksyQWSBnyt92EdQR65sHfEhk
1jaOWRvjqTuRo3CN4U0D4Jg2lnc305MFigylCnDH7TpFVzgQGP3/cKZ1RbUVZAHd
3yamvRLpqqAXKIKXSe6jTo9Pu7k/nUo+3fX5syawaN/hYxD0W0H3dBfuM+wLO8kr
6KfQ5EciQWaSgFrhf7lLsExQ/JeoQhyQTYcFvTdTrqery/zbsJEJp9v0gtYUOolS
vwMxKEAW9pZEAr5u279TDQ09rz9L9mU/aE2Ix+mfO32JZ0cz0INjCW+sM8Ztgh0l
4qfuU343O/gGYf2YZvnLOo9qxGydNynsKu4DGjzZuN0HXliMLgtc7GJZuTgdPDv6
iGLYSGCL7kH+uRrn01OEOtJ41zxM5K7v3ar/KPK1a9J/G5FJwerq28B/082BZWSS
hJzKNNXutecqipBhZx2Uyl28jpc2NNihBMEfdd1Ii+d+NPVUaj+0qheFzT+84a2z
r8ncKOoPwQfP8eBm54HpCrBBmqYe3f9SFELT5O0ZpTa3LdFIpfgPR4G3KP/5JJai
n661y3bLxkKRSsrDU42vj7IHWtP2ZN4YdMLJdYtsPTzqLQ14iwi9ZCjuhArzwbvi
icjeq0RWrKAMYx8l1bQeOQ7hyLMj54FSQdgq2w3BWI0PYNlQbs+3zAClt7NBbmDL
D+rPVv0A4Fo3FXu5qeYs7up9XAodtjnFdTCcvcKgDVIobs4CWma4WfLOfUV0IGBl
yhDMbV5RZlnpsF10xZddKDY0DVJe4jr6Ni7mxYGxneqgOlhaNdUxzcn6hBmI54v8
E/B+A36ljRuTXOOp3TOAfE4BgoLGX5+Wbx8VLSItmFBuh6zRIyfow+XlY2IV1Xvx
W7ObfRtXXxD4HZ2ARTWPcju7g1Q/zqFaJgBoqYiIBN7olscOH86pKk/SHdC+c/+g
0rGO3sML4LsaLNy/3XEFALuHFM3I7KeYGmV0ZvTxBryDoB+x7tKgSXCuA+IXqdam
LZ+W0Ra5Y6sEV0lTQWJ05SMJ8ugZqVFjD8A4owAnls+Nj6rW/PcAC6et04a2Hu2G
FD2F5mxlj3MGXyfuVjzxZZEQVublUc+fI4ftnszNSoCIb1+DX4pjDHeAKwS2ZE8s
28557uqE5vC9SX/Fq6pqL4oxR8RwAKh0knI/sJKpk62qVmWsPaq90GdYyFc/SArp
dV+pnsRemw7BgGVi+p8kwVEVsO6S4z3RtHGyEmU264tRQStP+gT2Pw2vqaNPF6qH
7bF5GqWaLLH0jis7SAOwBgkWCJcYUJrCeGa2eyPggD+wij3vypXyERMoxZVnmUJV
AzDPPyS4XLe1h+XOfov5TlUg7AlH3OhrTxblOHbKA52TL90GkZbV8Do4vUN83yAz
H5xymsAQF8iW0vbrekUgOEOdS1xCYW4ILeP/Oon2KASQPk+Ckr7g/tyh/Wl3kvZH
680jVNzCUQhuaJEJdDzjZymltSnZOfA6aRYXCE++zyAdJCIcUtVdXtTYJmXM5bID
vCd7Mbr4atjDU3Ciovzwtk1vLWJvAyWk0wm8tyPFys7Cl4uGGukC/YYm05NPhbPJ
HUn63096gPUnXGcTPiGaxc2ZJuVSoZDDFkkgxXVJsZ3AdnhStyzIYe88iD7cU7kx
dgsCnpgKoBeyfoiULml+y8x0+lVgHienEDwc/Q3GpLUJW70M0GnW5h7yrIdJ8F3f
W9GqvpuutxBM359nQb8NAesdnkckQmPh9H2zlJTFQLhMfBKX0Ivdl1bgmmPYAVNR
HsyRkcv+tYh2hr4DwV95zv+93Vj7Y9aoxe4hdUwPqL2fUpG+0O5fw6dSGju6erYt
0cpyF4m+sfyo6vpGOvIl7dpFVPxSwGjOYgJkAxML73inXhzQgbfU5uJEu7POLJV1
yPa6tw04mHAqXdN+MBuDrmECKHksA6F22j2FcPbdl2YVhcNUcCHemPPVkwLfazxC
7Rq5qBuBNIP+GRiYHCTCoV1iUo6vogrTBgWOq2XDbCWLpUsGx5IhKr28nrTAEJ59
Dj81TZu678F3PyRQcz9VAPpp2AdqIpE0g6+oOOVAC+3Xcp+meSrNkKlB+q6cJ350
JfJ3DmhAQPl84HwPiGoxjfyASXf0dqDlWjiExqk+OPlS+lYWCoG3DKqQadfgXwUr
+qCSv2XYwM+3DDqrAyQlCE1L1ciOW85+966FHD6kJA6R1Vc7wcktcXGVTlGzX6MX
Bv1QYOLYK9aEgVi0SGIRedqp3wEVHaF4SO3gSH3tm63lXirhCxAZogCDP65n7C+D
Qp0gc8lA3OuqfQSON1xvYv8e/ahLmgeNvUvNjcQjRH+Cz+uGRUkAWq/CTUVPmuMw
77KGAvchLczLKEMYm5iDaqPoSxx6YuufijYeC5RuNY/R2x8W7my2fzFv5JSlj3+V
62ssGaQpGDXDMZA9LRyMho0HyCntEhUSP6qlFM5OPy7k/7OFCv6x4XPPG9pCTcy4
LzPzQ4g8v4+OwaFOQbjvFrcioX2I+kI7y3rnFnS5eKXxeJKVMAWqC2rJtk5cjznE
d+co7YDDuaCToFsuJS6f5Gsvjy0vNPiYXS09MspRfGobObqPG3s2vsrZrFd3vuPZ
v0gS3X8smUy7hbZ41l5XO24fKVMkmgzPKbyOCIqpUkAaEIcg5aC03pMsQiqz3sys
rhZl3AuEI8wdr5WQ12KEOz+sYKDcID25SLJCK85GLobz3spcw3MYGhnK5gVcXiSZ
HU2RKQ/GKILN5OJ04hmd5gtNuVUNZ0X6bTtss7Cl9R97l8JrGJlN7pn5ISzZhH8H
KukgdbRaa9XY6qP4MtgieNRgIYh/H8K75fosbZLpT3wiv0R4zRWGjaCJa5tr5YRO
Pi2I0ViztLC3Dwoks2dM2MOPz43Hyay93QYK3SAEPmBZ8VMdB6ELGZv46rtUjgol
a33ZoUpGxOEu8NLU2JyrmeZ3IoJf3RM19uihI/7wngelxtYGow9v2ZlJtx1SVitL
t+pPPlqorp/dc9rLbyFpuw+Aiaqi7VzBL9cGSheIb1ZiCRc2VBUmbClwncjZGdZP
UTkCq3k60TKwbhfRxOTJJhHDlqaHhp/26WWxwI/eMpSewg0+tp3tloYkiEDf9lKE
0Oskw9NEgDgGqGF8utjrix277CfMHHWM3sE4GzID1YkfY0874Lk0ZnWlgE1ZY57D
AJyUIx1RIWUCCS2n59HcZc1OE31oVaDzxCQ2HNQOGgy8GANXG4W7vFseahAB3wjp
PNs0v0e0v55eLz95KbD7cZTsnzvRPr/aR6gQM+lS0AKm6gbaOEsnO8Nmxu8GeGmp
cmDkmNDzeKUYHqfAW8q+1ysBsAjEHOR04NVCamr4I7r0hiM3IpQfuohXrg+XNYUn
Qfqnac/zGDa9ezYHLoV0DZ+g8mfVxb5L2gSKKQbGx/jiq/YNNHmbOLxT2L0F03Yj
+M29WAprP1W//BJISBzqMBePhE+oz7EHjeUq2MNlS/nkSFylFrqCc+SuAIr+bGNH
HChiS26y6vJp5RWAPW6yosBGS2WcQErGjjHuCPKGasTNJ6tzgLIqGDocN7BFA3BG
STWCFlMqmzQpeLY4/gEYCtGFd6zANRNW6dWczYvFUf5BAsorlSdYfE48W1lJz8F+
XNlWNQww3YUtDiEtBksXJEUJLpaTzp1g49MV9/jwaSjonKHXHl9D0xwiPSeFlSxL
0/5V7vRZoaVXUkEDCnuTYTa+Psgo6dCLsiFPvoPHI3XSOdaRh14SURbWiBW6YP1d
dQiBEtMYO6ZZr3eAeeoaw/IyxiVzceF/OU0D8T9gCx0FIKLDTVirJHAfCtuImcxc
N+Kv/IwHwvQ6qFSWHomPHJPbkQ67nCd7gGTlYHUfeeTNL2Jgu7JQC46NmF3TkZy2
MViAqHfXBjfKmPXtwQuhHHDFCTcChJnSapUgZ4dO8U5JWr3t2QRzG/XD7PUYrUTP
9wb326dzb2+dvjAYy/X78dhaWIandYwYUuxu3deLgMB70acRpFJgi2oVoMdvPsyU
3o9tOsqfeArM/1OuwOb01CJY4TFR5fcIXSslG4xCHIceQzTsZLdd7Bvhf1pkjw8j
X1COVzyHHvZofaJGk0dh41grvkdjS8eidl1Bmv5H+FdKsMh0e+ZqxWvPBC++XVa8
HNDy6lZjgs+CfLprtdsb1BQnQKB5JtMqaGPsDrgqkobarJ6I+JQ9iFZcscdx0m/6
qhQN4sg4Cst+zf4T9CE+RBWPOJxmsjBPtukYGJF0WYWBWspWmQTP4PxL+Nc3aqXr
8sEONjo7KYzUThUE9hcRjp3qrrQvHN5IQX3mJGV1au4nrQgsPJMDrcWa6d6oSTgO
iGld3qbOgZtwDGZih3l7wSlmBvXH1+eerzZKuUel6vC34xv6hvup1FcFwNZ4cIS/
cGZgLe76QcmuCaHYkLLpkAR+CLEPSdoJ4Z2LKJyV1T+OhRq4SlTtI/SggWpMwCqo
mhd2yinixO+uP/luFwlTidfmuXvyhzHUhmIdvAkvvt8jybyTLC8/62eonduZLiaR
wIgph86c8J8olCdfdcWDHkkgOn9s5uTyqVllIpXvnR9Dhen53yWk1vMb/eTIVGdy
Tt1VZCMVCoXKqYmopuEmNgOehv1bOzoRQ3xoGY+U74CJ63ElUJ5gbRU2eFpjTN9v
R5U87iwj1/wfsepmWxM3TB7HyVI+Rfp6/o5Z/SNh6OLmbqmiZWjJycwQ3vpGogNO
CfMNPO5JTS9GiV1SVCZu2dV534azPcNxvCoy+3myTnDs35yGfqLNMGXIjc9DZoY/
d8BF3v/AMRmWece6epLCVeQn2knEw4Pf0RnPUMNHmxu1ovxpyqLmNevZqYAX65kL
HHxTk9ffvw4lo37Gs6PESOn8kqAbHl4T491bUjYYja/UE9tBOxR/5qyFwTKbYlQi
Qsxz4XwAWAyBRwhQkEmX+lIpoPdY6Cyd8o/Pq51uGfsBrKt74skBCOnrPkRbGlKG
L/N9BqJvYYqOF+EUnkzda+3dW1vHZfXXQgicPt2Sy+MPfuHEAc10XFBcde0aUaKw
YeCOejjx594pqOG//VqSFNgPlVKtsODi1Ne56txhknE+5Kym9diOe/JOL8ztlRcJ
b5QqXvuQOWftWKGIsx5vbK+LLNb9RziSjSQUlswMGJ1IPviu56vwS9i39Y5VkGZt
VKet67vSKo6Gecdo5WhRaVuwjQKjTK2M2OPF+U74KswgNi/yY/0lTS53LyIyhOXW
IcVihxjyDdZasKo31S9CqXL33xfivws+lIpEJgPyWt59jQ5rw9rQwYPhT8xFGiOE
SODGdRkj65a+r0uU1+vb7gOWNvlSz0lMRXCZn1VK4eWiKsvx9DkHT848JRmIVPjg
IxptmEliEzO4MWJRSPD8tChnjF98mZ6j6SwabnRgVySFao+idM/bEIEypyuHPUpV
`protect END_PROTECTED
