`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hvgICNnjDWuuIpuXzHxfNECUPEwGVxyuZCEZrGY0lIyO4CXGFjYRJZSiUkzVIZbX
KVkOYx9d+7c2F2SEyMFAHv/XDnfH7eGAjK3NF89GgVcyB2MHbR7o5cF4A0UqoQwr
Aeu+398taHdEPOPVamX82DuTvJZIPWxSsHfM1tnxSfCZtkm2wbJb+t92BXB5jAvP
pLjICVJCJLZ+zPY3BXg6l+QmN8vxCVfyXs93Mz3ZTRuxJNR05PdcSgqK9UMCcPaH
Ns0VTLDbO3kjuf621CUPh+4Tacvvcldop/mU7DxPKjvDratW9qk1UsjIPYuIZ4Us
yA+AtMvSxNvlUwBzhgCP1OjtDEy1Ujhpim4h1xPbFqpiRo4yCYpX4GGvZZ7QPpEV
l0lunR9lCiR+VPqz4sMlt8t3HrVX0j1G7Ioe7O8B/lVMZ7rYC3H6DlysZ/hli0sI
avHliBB7myKlxl/4wY4xSZFy7uHEoMIe5I6pxCJSK9omSLSXq69RmXyKitCQNxXu
2UsBuwAsJSmI4Pi4ZdDAsyqjS/6MaR9ARwuYQIH28H5z08YAbvJkfTHlkSA5cjZX
/gcf8hYXYfgyS79erw9zaYj3j+eALy64appU5CcFVToTOT+/clEjLU1agpiDWOhg
e2Q4xkcdck5XIRj1K0POSlGDfC7xvFXdXxh/14c7gWkv3Ki+bdSMyENup0oDIf5i
sBCdkOYOhMAWb84zCvDAjeQhMzci3AC9ySzUB8NIucs3Y5w+aPtwOnLRGHCErGLW
PA5Bd7NtkAZtQed5PRmtTYnmweZdlo2VD68OukkZkqZqbsoYquK2n4yfFFcBj4ky
79PXyMcR1an4YfxrzkSKaTuIBKWgl+BbxiZaUtEfzivxVUtNiQNYm/bUN0XMCnVa
9eTp9Gca0yd0CupCVdbPPtKVW1D06V+bpmXhafmZylXBGW0SyyLZNhuaioAbONS6
eJAU8rSptbt/UUNhDB/DiWNf2/3WbZTzrxRcPRL/0lu2GCGiSVHYtE5ye7vF2s8e
K0XzhM/SXxk37qpMvalLN+dhHR06PA0PGu95FVGF/sKlkTlkWR+eqei6iGk5qdWD
0r8c6N4MqqD/ZlqtPKbqutoKAv31VKvPokH6wUuHFRUwMtiklhrdB8ATVLJZs8FS
jLBK78f1lsyyGoou7J1lj118HAmoYM2s6mQqM14CPO9VhCEubRiHeWJ5W7UbRR84
H6mahndYJlKhBZkyYr8AfJaIneEUGQ6DZwcD47gPjrjA39XFtVD5l311D3NYaf1M
Z/6OXGzXB5QYGyLyJqKmk7GSv8ujmqCr5LkZKgl2H0f3sxmmibSSXYLZNPiAMCN4
C3m9jV2VTCjmTS0SFX3LfO9MbeeUflQur+4O3JT3PQHObJUkYTfNhCqMq8/36hzQ
sg6iwaOulj3KyAVdj5fHiIvoYbeEAyl7N8cwyPedEW0ow9SuA8himylNNGf2fx88
es+g020B9lsVrl4iY2KpCuUn4kSOnYWgSNajDYd6OgWcXMyBFFkJztw7Kn1JntKj
QMDmgBJBjTwC2IseTEtaOPNK1NWtES78vWx0T7KVYArY5ANlEeHqIdlWeQdE+lQR
V7iSDR5HPar6PiS9UtvRQynMHB9V9O375sRlKEiJWe1pNX5PZkvjx8NdwDB2djWV
DfTqkPznNRUD7vRl04a6OJb659lOl8cwYk/Xldwxr1TRtKkIRfkpFFWTQoupFuOn
hJJ/fbcNoNekNbf5YOLet1UC32GPk2e0Bybep/TbSkseu40Vw9oXUB4Xu0r37sGG
+ZjaU1yBnkzjDMjJ84s+f+ghRjp2m2Pjvx60yhf/rt1MPxn98hP1W/hRHWPTH4gI
/sYiW25PnAQyhPnl+KRBghI6y9aCJ5VWAez8GvSApOL8jp0ebqXK3m/7Jfu6tceA
+PpWjKNCBqich91+OV49vdYtlY3zTj2CpUkih+uWNzvNxYykldzmMmKWoX/wRh4T
NTn1FwtvZI+ffBDwVHW3ppVkFqGU6kRoxRemcGkmBXYBc2Lgw2vfC+QzXV5PXwu5
jHCVF5VQGCLt3WWSDaOHDmMcoI5exRbfyUGDrZTzRVdYzshJ4oUOdZwFNHXSJbME
Q2T8thHOCIRT35BQFLhl6coBFvHPyz1IwM/0nN+y0KEETrdkAE9vxpgViaJO62B7
7ypAEvgK3oXtjGaWVVc0Cs6nfJXB5qrATrgFi+JRd0vmGaU7VTVIhe4UjxdGBWIp
Ub0L4dB/D8H57b+LeaFy2oiIvjTS3ifc9AM6+DyzalnODeI1mqYQegCP4pAMzffT
`protect END_PROTECTED
