`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G3m+G5oSyx/Vj08ty2rSD4s3rNzOSFLoItErEA0n4/LYy4r0u+NWVxkDhDZX0rSN
20NvRPAqeas2arxYB4J4WN1pR4um8uqiXOwkYbI7FrSzjID686YVeUNv9Za3p6NP
MaKbT5gEXsoUxYHv+UuOnsNxOrjsY9s5r2+ypy2mcs5zg+wjBdmIxlcLvKcz6RMq
PtimLDHhj2nrM9B3kjLMHok5l3SrDcBJRnpBI/DMfueAzvQV4ww0ahMkdjjtDn6f
SJB4vvMsWTFDnKLWxt+V9w==
`protect END_PROTECTED
