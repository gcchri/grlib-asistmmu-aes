`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k8qSo3eSdAP1pFnrLJ/Y3T+zX+M890YXwp8ZDXanHEmKcnAxVTtkW3g1KC1sQ66S
jbLKAQJAcCtTU13aAuVyTOPJMW56/6gUeT30iSrXiXoGKVC35PP+SdTzzNqJiPJQ
+b767Tcupt9it1ZUs5RXcIGc8cN4mbx7u3F3WJFdibsNDtuV4OWB/+S5IpprwHj9
fXVdEeM5ja6kz6F1P2aHBIEYCAscXQqcRRkzRqljE+OclBrq501SS3KNDaAhAr3C
8XHcwb6b+rXSpsvCSSBJgStw4JzSd18dwLu0cRbplo8L+Ac1Uwbo+oN1EitZP8fZ
9gMyqP1XShgS3O5++z2rJ46yvmfLLsQV5b516o0P1y9/EGYwRDNGLmduSgaXeGCA
rFepQFMO39ClnQZULFppLoPbDk0VlSoOF+fG6O6yxo3tc6693pyOuemlV57L/beu
b3+LiR3Y/aSlG5MAZhO+sMZFaYAvpIzWePeli87doN8qtVif+P++kcYkD3SaqK82
KAVu/HDb1dWo2upuY4tAOFyNrQu0m+XTubUB/G/4YjsqyiAJo/Ksck2uhV1woGwh
8bs+JdIjg/nz/GrYfgLjlaHNNf5YcJQlCfOJJ6ZMbSRjSYUSrwOZztHUgieS5ce0
QEUXsl9e9x3z8RweOXM6MBvSwpM8c3yPAjq2PE5Mvb1cZeDNH2dtPpy2ZvpmpQts
XHUPOYkx80CluY/zXrPnfml1STBOpGMqQRuQzpf03NJKZR8cVaB+HGCWXhvNR5P3
SM0fOJSRNsbpcSir/eGdualVKlQnHciTmMOrfm5kLN8h/vBppWFnboqn/HsjjZfb
7Y6RygIg5KklPTbODaHpjiqvBrsOb54lFnqEukTngZevPExl0xU98vj4J9Z+gihS
4Mlnt689L0nkB0BBPl6Cvan+Ng/aiCoBWJBda0L29UCfDno7Zax8ipImzw+nyTYv
0Gkv4bJZscg0TslbC+/c3Ycq7MYtG/I/EYWVsPnAO1Nmo4ma+lxwd1+BJFEoIyn9
CYEMBnXSZ5Xyo3+7qftFAisU8yGz8b+872CCaVXXUuhAxQ7VNqIU6QDN9mivNn4z
jp84PP8MusTSV41yzyZ9dUilq0dog8TV+Mm6rtPth9dmDH6iNsTx7oQ2N9bJKdb8
SwMKtFGJqoqstrD/coQ+icamKIi7tZ2n7ktqVkn6EkY8gqex6kZQLLx+ATVebITw
hXLN2w8NRDXw+GK6mCjugg1SNZkagkUw6ywWwf1k4LJBewFQBngwCaybZvFLt1Hy
gfSR7MgFziP2EsLK1DM4HT9SMNhc1SvhcCWp9k/1a2OXF1EkYM4ik9Tbo7oDiBxs
h8lZaKCWjXANPACI/U43CmL1rdTFN3p0FCGkpAQCoC4uZMTY+MSTtuYQiRtY5r6F
jmq3glhDW8TitiXMVEUbEgsWclFVE9cjqFVTH6nIxMqq8H8fvfJRCAyGxiTlbTfO
cjDayVSP2Rn4wg4l24Z5hHrP8Glp1zaLU2Zdn3CmQCuCea5PhXG1DNj8PF4ooKiz
XltoIoEJ8YPYJ3oY/JF8p4LhxNg9JXlSpoV+nTx+gEsAbDpAo5WXc4MX71AHScWp
VgdQjJioVX4pQBcPI9vWTXaLhE2EaEMHVe7dReYbirBC+lPTn6TojvLSsjxRItf1
OAsVBTnrunoH4jrwc1sTUJiE9a/h1BYqlCp1Yl7zn4txXGDWLoJZOyPrklz+HJqf
dPZKvstPusYm+K3DUbJ3gPrbF7R5HKiAvgqWK07OcHntZOXKCOUxCRH5yPl8kYqF
aFXVs6HO2yACTFHWnW/v9GnXT0/Bt1+6/9wThv+w/nxTzDTKy820QdJZrrDP219P
oH9BY0Vj9RRtwFw6vfudXKlVNOgb3O2zgc0WdPj1UwiXllvNLz2Ml98Y2IEHfow0
HKTm3GRat8hWIfRVYbf1KNCOp4VIEPcLpkkwISMcR5HX9Gx8UNueQCh8Pu1xT6kj
Ho/qF0dQnSUt2cj42Z6bu8jjKIcXTTefd8KKeUXJOxtEwlClw/F6P7Jk4mXNlKMZ
3VUg7MCL2OdiehGZjTY5lxXaPXf4hgxXpyLKEz3bnJ61CYBuB3hiTjhRIIcLq7U/
v9l0FypXMmUQpX5WheSLMORxOgzIrI3kGMe3Xv+ibgGvlCvpP9tA6TpTRlZEHGFG
JGxtqKlnSuwkIdACKCDLDC59cyTLwhzcb41csRnhp4vfwz9o0N6bUbh3IBpn6FI5
vUYFEcos80Dl5bo+K1fXxkugg4wSTfYTlNa6FUjUZzfUM4CIhLtw0golNVqYAXec
/DoJAgYERfeaItsSrg9SkXdQNUfvKBDdPkGYy2wEQAfwuRK6kuIdYWgTR7Xy1cWS
N9zRPRTj8nDadOgbFCr1QWFSWSbhpaWQ61YSKHJFWQQY9ZUTEo6uOIJjHcy5Ix+F
tPFr3NztU3e77i4Ahc9knOjF7wBN/W7UY8/SzNidb+vN5vMQrmoujxajHNqJP/jw
AYyUwzwb+T8je/lexE6Yytyl0TKaQA1VSwsAlplg5r4vHp9cQNYOfvdyGQCtqk1D
qyuvJ6fMpX+5Xqs2M65V5ACpzXMs7YMU0JdgjwIpexrSYoCNv0xc2zhCH4ki0Uvm
OaEvhqCljRXHtyafAD4JQpfHht5eRT9sjInDjYG9tS7RX9h3a/U7G4y90YsKiIC/
Lqlffo6PtQo7evqfZwVaCFm5kaNoxfpsnDAL9XXYvC30R0DB6RHWCMJM0ohZWaQv
dhtLhIgehFR6xSlR5vPU/NX2lQsd/ICpAGDEjaEW1mhbYr0guoob0ymBGw4Me3Cr
pr5B1o/A4lBW2tmXULx/tVNQmDuramue/0dyclHXpJzaBldFUcq6CjMgarmFc6Wm
PAfzGMuV/mgH+O9NU3V3JEwsFI5CEbHBP0U+uHZozMxeq20ILw0+LcmouIt6m1OV
GlGHYGcU6nGnr9FwvyavmWeKBfnYpJie2k3Dpo8n3+cOYs76yI+hmwLp8G6lwtzf
1eE0Favbwf1oEh6oAlF07VyEZ6SM6gzasKqM+86y9u8Otj16S3KdgdMaaCc9OpZZ
CqukqooSVQFzxAn9M+g/jfOLRjD47Zk/lefFbYQcm1+Jdc06H3HGelqgrIK+WOmb
OWcrldkpXJdPQAXzRWcBzANlX0NAGxPXEOIAb7OBJ9RtV4eiCC9XG93PPh/WXFLB
Sc6p7yRN5f8mvuRizmldXat1Mibdb65p0bid6UDgSdb+89gyfoJeTrrM7KIqH+j4
cgDad1hhT0znX+oAyTnTAuCVKgaiVWLxDjF8Vrx/wxS9UAUMVIbZrm6aqQNOBPwF
W5/qECOnC9GgKDl9kHZRoJdPW+gl6a/bRufGuK5483HwCiGZjSC2n9RcUMtkirh/
j/IMdL3j0WV0XjLcqoC5rCqkWzDphxjn9P2NqjmIW9nPlH7AbYLH9eZNm1puBuUm
t2lG/QhKJMh9diD25thfH5m5OnGo3K4lpn0gdPNOHaS3op4IwAzwW8dbCbKQoY9O
MHvl8JfY1XrQgXF/JLRdKMQ4CuI+TeX+cVjlRfpySBA9YQw+ZP9WtpKBcaqQMsPz
nfX+hGheBhAFyCrIgpl5m6Izr+88eIENt6+ZbVR2AW6O90i3Ri1+6w6/NptZjdyV
zfD1wZChISQMgZrU5eA0MiQzaqusWaCOOM6zLQhE0gb/I/KQXUs9tEQ0MI+YQXe+
xBM9FC3ob3YX2e/ntnolHPc5JGByuBeIzrOrNvsfHGb1D7mJh0qZyvu9VViPpCql
EURDusZ0A3tjDDJDuLrHFHlQtIjd1H8U+2GsnY48xi3h8HeqsH3sIH/XkeyoKx+w
lC11SQBwip5bu81aMClCNGIVWBSrcR7AAhfEbYgmS4wbhJ7Qu1IIXMkQzOT/jAUz
arkL94chc8mLspRzj3PuM+xDun1nayKXBKjJqwDlpAE4HP4M3/Zv5c8WY8Bczfh5
oZN79khILOVX8FkR8nqSR5KWXnlxl8cJAwbVq7FsoL42p211tNQlQBmQ6PwnSTZ3
JKeMkkqWSC5Hpt/LOvjfG6iCwZKuQ6lXE5DvFPlNO9LN0R3f50dCyssGLtAF6HGe
3mOo+jdP2+dcEgq9KVBnVW719jknT9i4Bu1fya/8HgUbodMzrcbDG/lvyS4qkMBX
tbFVev7XgP/CsgekfdmNzLUTuNuk8j02wcPZsLDNbvG4wsRPHKOs9qtYlfuea0Di
zPx4MvG6OmBfSRdPkJooD8WahdqzRsQtPnMKHczlS/aG3WrLeTg82HKE+4yCq80n
TEUP68NuL7bGnmbBj97trN4u/8Ug1oMMf6VgOLkq+uINrrfjmPFdIBHglXrTzq9j
/4DOhOpC1UGgw/+MCWwKEeorkx3XywsUoZt0yjvPN7tPa0LVuDnvwFGysO9U9kba
pGAp0IjGBa+uFxb4O6nZX/drsYyUv0LF6cU3MnNb9ffNcXsEULsUzRHdItvTYaQn
IkhPHdGtsR0fTQCkINFta7gr0LZtdEVrIYh++pOFAqdd91h9oXZVDEWYhoImBihB
y0iVK+pl/toi8CQON+CSF6RNq6qTdOOoSJWKBzYBFitpt/nmSCop+N2T03a9yJqO
l8+Hyf06jA7yA44nl22tUBafueDEKT/USNEkmaOp/v/wROnFtwIaKl6mNP3fhLQG
bbTEqhZ/AhUDUL5KbiwMQnnrOz5HrmGBHYQnFyqzN+G3eJmdrqX0n0i0d3Sc1A0j
dmYdvDZXG65h1qUKVL6mLAc+NWdsOuTZS8XLOiYC/jC4UhZQwy0GAgwLttVBSWI7
g9xopn573yNZrNfkXsMUH4e5xQIv06pqWhZSjAGWmKWyq2ma/RicD37t+T/cwNJJ
I6iqBP4fXyOQuWsIzocZhZlhBrdZt43e0+5WlZCtYPTFuqhBQPYrR61YGsufErBM
E88Dqmkyj0i9TO66C3wsz7jD0AchFr2j0Wgxt3QqEEkgPp5zZ2pBczWHsLKSrlTk
mOq/Gd0rugafwMtE21Wz0tAuIaeSufbHVMaHgRzZJp0cFLrXmwizSqO3/IdQtHSl
XBYRiEnFJ7MZe6/5vh0l6rxMRvgVid8+h5hil4yDlvzXf49lYfa3iaImRChHPAXz
KtFu12oTgMbKepFfIL8NV7tQNZHUB6Y43K+L0F59yGooxBExt6IyWKIzQh1OiMWr
kvB1BU50pNIzm6I2XO2EaPnIjwokYtI7oEF+ML1fTbpdVQ3FjtOD+7j9Iv4ETf9B
uWqLJWuUTHP+xuxwtywO+XYsltiqkYLjgaFPThIyfK5duU+i0stuVE0yljRybXTZ
xM11e5rZZI5LoF21cNn6eOK1h45x+RVqLSZkdfvR3uJk2l0Rxm85dCQgoJpUUB/W
t8yHVCHYF7G13fA7c0SU11V33g24NdlvqIfvfvunMDUE7YQMnsDi0JXa3P0w/tzA
6QXPmcHFzgEGsvy7scWWwB8gmU7B1bv8orIWdJjCuvZnp2VBmyxmIsD9ohBr77hD
k1LnpBI4Fog0T05chy8EJzqc3Soo514hbpNImWt7TG/mC7NjDYcx5pnfkUhNGVN9
e8hzPcW5O970cmaVF7UUpn0S2k3KSZXm5SzJqCts66C1H2pE6pFRLbb5s0c3JBiZ
apzxh5VMUq3Iumcyt1XKihYVlEbpFRSgQRn5p4vbyaOcLnxslb49U0aPjID/3YhJ
CL4/pIyCX4PweKWH5e8nsOO69tilVT/RUt1krNB7hFma8Qj0pTW5tigrcMkLvLiU
+X8KwruW5XopJTUsrfelk8uEKiPQzLnrjDIuUCYDsSNYX7ut/wA2qdiz/V6Rd2aH
cKhRhWnYdCiUhYNc7n5adLZLsfZmHXDgYZkidEyehWi8Acv2/2wrFliVZFTRUv/1
SKNrN8Y5NhjatBodcx6z7dIdM/XwnsmmEWjC2WEhvM/GSVXHXN4Ihn68daaQ84qD
AAPmKhvOM2ouT86W6+uX9Kpnj+9DjHJs3T1Aqd/i54DTb46sy/1S5YmPor5NfbUo
ZxtYRLK7Eq9ckCsaj82/Fk+XDgQYGRXyht5gnXCCbp3y2CZW6AONqtn2S22ZX2PC
LVXzUX6HFOHiX2072fI3SI/pjuk1+K6RHM6R+GwnAfJobabhH7Y2C3ByP1cY98Zl
lY8SCaHmM9UEpLgHnCaXOthKBGpA8ykod+bEnC3IRqqT1AievRJrUvw+0yeeTFLP
3ptsBzmAsY0yKDSMfMTjWdFshnSf60f/irAEkVadjd13D43k8EwguExpyOxIgp6a
M9/vjgWl7OU9r60pYGKgpxh/rMVzvKF4n4s9Uhx+K/bNQqsYOz96GaVblyMplFeU
SO1TxVU3XShiC4PpJr/UCtYZb5YrOTGSJBZIfOkLlLFwET9WZZ89JJJmNbzfAT0f
YlaG/+mOwvWLgDBgxZdWuAMT8SWvFqyIe4v7v1LfnxM01GXXfN9YyiOHBPRYk9H7
R9HEByF0EX1HSFScYWSgUD49EC/cfiDkiDwqOhpDuN0IUFEP4jz5A9iUwpTPNtJ2
830LniVxNTEB6f8B3BKNsxyHGYev+BgPmRhYIkhRlMMUEnGlg27RjNtoTl9NWqM1
YXKK5R/YtLQbOI4bakAnx8njv8XxTxP0GbgG9ycQoxOrWI3EkHtfxaLWTsjHFt/j
sQ35qhc+17QJii/KtppDQkAew8bdk3+aKJIf/PPavR7eX+dhuxYXpHqm0Em1b4nD
VKm+CPPt2OgVF6nwi9gQojPIRDfyUD2pBmtRrIfwylJOzvq27Sw3y0xR0PajvGpk
5gen2H00xdvuZ3u592KNVvl1o7omf1vL8Ly2HKHIpkWq8e2xPPUIiN+m4TMpzuuD
E7WWXQT5Dmqbl8aoFSxZ3WR9yoUtoixaOGgMxAjXpD1NBGcfjs7uXkQS2LPmfIKa
aVdN8C1hL2J+rByJfnKq4/Q6L8+1VV7RIGF1kyGSOxCe9Q3/jHqibm90HWAK+1Pr
6Hj20ukz6r17tFpP2z56gzu+VtHz34AGtteVZGP95bmJbgeFS7MYnF4HmXEQsT/J
scs5AhdhpOnFc+15mysmOg2dYWIE+HHR6sdV7BtDfM4JSh/Oc+5B21vQYu593Yq7
QE07gSI1K3/7F4DzNCldOYK58VBzZBhVWXT1ZWHuvtOJmv1nhKrVa0cGDxZw6qeX
tCe88I/F79w4cIN8BMx6zao4+cb8G3NEhexdRJ+sB+RFA6aMHhuYGJBqqV9yIhXD
UkT4SqSaL6QhPgE6Etki5NE0Ei+AmIYvpFrt/ESUp/3hFhVLNEQ4KFMlF1Y6fxzv
c13WYQb+bAf8bRWQKMkfERA9n07HQHmBEay5LGTTuPE=
`protect END_PROTECTED
