`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JZXIjU/bRVqSDaeB+1wWKBDFs8LpmqpuQHG1AfsW5M7/vU2WqlyTMoQV+otwY0kk
9YKsxKJPUjPQEd3b9055WQhoM4dmGUhM8ddzRoH2zXcwLVfLwLNtt/xeb9qWITnG
ObwsjEvQjssF0NKYKfhiuDyq9dmjNEnZwIWUXg0VhbbnhlsOmdILcB1ePzYhY7BJ
Cqy22DKTT3/JoOcOEa2sL0CfovPuHrmtsq0eknVeaZvMcTAhyZHT5XBuqSOqZfaz
gMPguWa4bR4kf0kxwSVpLU/LSlVWt0RuUEygaD628mx66w5f174fIgDFEMdDDZAK
icSnV+DEaMSpRoWM+pBpNfRd8VzWgIPxkYOz4gbtk2Iq/qYjeKemupriGU7+B74H
6yWW4jPrg9KeEEjHe3FYm+SdmFLParDa4ZflywvnKlhHM/Al/IcGdHUKnIBO7sEh
LaRIv9hmvaDkeQVbut4EDJMaZaLqtATWFsoUyVt/hcab1BD7yZ6VifzHt5OddbEg
R6NNqZSr+W0fxZ1dyfYLKpvy0b+f/rEJ7znOIH5hvoVwyyYVo4dCBXdZthjLrGtM
89AyfGdMzOq/T4DzwCnyvxgWsinUwdooafVkQzTKmczm3nto0x9yZfX5Y8CBTCB0
8wtkVnlvpdRa0oWr4THA7WemseuOM4etUGzDnb0ANodggzNcmwgtpocnsZ+e8Ucs
ntu0aR0CsrqagQL3ZIGHVR4KCaZdBS69xY8APv3F8fw12LG4JmStCs+IE9wzOd9s
fTyvaLJrWr4rooXblEm6X4zDrKPWysLUzRveeeXiUylDVwyVF5Y94dF+WRS/H3I8
B/ouPAaX/RbEmjOYDwbQuFy0SFU07mWhLxSd3I1mOI649d34xIng7ZxSOTkNk5JW
ETWy/+YFp51kZA0UmTdCEV9oRyVs//mLNHkB6Z7BKRbOXCvvWThCBO4zUwfDmimn
W1gGOBNJS5/J5dzm4o/Ho45jc3/4cjWEdUQzPNaDPFB69N66EAtM1QMtieb9Va7k
u4KouznIGXpiaUuvJf7cnbpyxxEfE8GonZfV8BHgFFWfWUFpgNrXWW8CvrmPd5dy
rEDTGobm9m6fgTVGZ9ebEVIK/YOyitbhdKhlYQ5K84U8PScZsC7p+M5zut6ln75+
Wb4XP7+Ew44eanCga3rSfk1Y9IizPBqRKj+TgPlxsq5TUS7xQ06xFBFhDARdUzgJ
ZjBKAc+dhTVOR2BhPjRfWKEyxabi4vvGH4+k45PYAhAZetYhDfufLjRf/QGpetJ5
rPgYbdRx/WADvUDHgm+h3pI4s6apNFXyAERV42GzKgbifDAyQsbKh5dFOSpAkgQP
hbyGRrYaYIFX6AbD+ivBsZWG8Ts68mW9REPPVdqy9PXuSLQwLUbBa7G3XcbwUDFB
fUit31lGqVEV3a8Y4+wXmOOUpVVXhTocUznm6PXJ9hrL6nXHLRwpzQKQh/l9dFKb
+B/JZUxLNi0UCQ6sVaBV6JoUDkhVEpHqG0JoZ/RUag9WHK7fytGK0OHC4AjV1XXf
BBzgpEw6YEpTebgvtWOnN0RTb3lsggnAhtlHWWqZxR53lf0cOMZu72zCasl4snGH
3sLuYZEmptb3N63I7tiEWzlScqGf8wg6pVcrQs6UyzacW8JKsfO01QpgTn0ykHrg
OunlutXqVB4N/Q5nVHOfIi7jXf9ZCVAng3vNw2EFlHyo20RxKIHfsmWTGAN2vYiS
bGx0eyHyov2iUP4vKdkE2oF8qaJDx4Tr9CgGeKW7bXPIBysAgg9jrPnlOIknchLo
SPFP5/eawZbdeW4FFnxW/UsBTDnVo+xV/oJgxaT64G/mCYaK1KuKoueduhAce5sz
oueIG0W3KCyWDOmtM/sSLk6o98qiuRmrlpXU/a0mSEyyDESACXx/caLY6BEOAJnw
t3LbzGIQ+o5GdxcoKsaKQw6u3R7KfuQ6FU4sidCQBsmCIYMVzr+SWhk9p7y2udkB
dk5D3GcJxUBQ1jZbw079AAJsIEHdjLF9MBTGtIYfHEUYxXvBika++WFsJ/69icQg
rRUXVd8OgJzYO6R86lC1jHI1vWN1yCSuiglHy0AN4BxzsEJc8GaswNtZmIoh1lga
y1jwk1GszZrp8N+TDBRKaS00bmMhOtDsxItzGs/fovsysoMEBfR/qEvuyrHCtWRU
rgXjg5QxwKKwK6wPdjMpf5DxBDEIPZOSXyzyyKc0Sidnh+iBG4AiwPt1ncUomY4v
ad9tnmYEAeguP+azU+j4RKa+5JqB+0Z0Ug8m4SmOt3oywES5fcGTUrXPgG7GXOeV
Z9BDAzYID5wdXTcuEoSl00BHCpFRCTX0mhFeB8nnlzucx7w0oXQ8x00jnumlRjqd
gBb7MbvdAuCL8mqph/UH1pISRLYYiDKsy/cx0AI9KBrgcHxn5Axjr97BrMA6aH9a
j9NZ5Bo4MMM5y8bm8FfQFEehtJPFVoBAC81dC/6yWtsV3WaPBY91cndWo3oGiZmp
r7NO1PrjVDadNUhAn5NT1JY8y07TcWSR2aeK9Emt44eVLlo0WCF2XViWoiONMPDO
9BSsVXaTbz+xsJftLcydxNLpJkZUuqTBbpS2Cts/QM9FlHpXVPHSg2N0epPGXBZ5
QW2AAd6bL9w7w1y9HnSmmMSEn7pKuPXLRynM+gUnxQiLfg4Sbhl/88isjTU5xRbT
HHpb0BNuOoTatih/EaG4bKoqAo4CkNG84WILNBkY5dXm7GWZ/5Q5BFsQqQjewc5y
Igp7acAQD7diwpti9trg/9PFeJgPJ9ufP+Bnk+h01kPhC5Y/qdGroFi+HbrTYxM6
tMlDFawNs1+IaCKkyVOGFDQdCspQ9I9tQCxfU1uyeHNu75StigUppGnWk3k9ckVp
eByCCg2qNf9Fc2cLs5CgHEarSEcPpi77FBlGa7AwYO6KgBShI7U9xSl+mUW6+3FR
xWuXkcpE9p6sqyH0CrrFJhiKlQyMSLbmj+T0FPx/p3JE65eN4zg8rEp8fJm2kBZA
g+AnE++YdehXZvVj7KKID0jPSccEO7JlZiN+77G0yc77gUviCfLihpyq7HkBx/D1
hY/M5Ff7kDt/Lnd1BTO6qYUCll1sxYF6gX8/OyezXhoDyPSJREPzRFmqJWL5ijGf
Nt5sseqys1VVKr0LavScgGSPMfQpR0UFoKBvuMpx/p5Ef89ZC4uSaVvMTvL5exvN
K2ofzcdqhd8x8ioxJT6bpz6MqD9QPs1bCDf0p2haicObd1qgTonRu5NfpUmfaM0H
WAyxDNbaOBYLubgOV9Q5Vg==
`protect END_PROTECTED
