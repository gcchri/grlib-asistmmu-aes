`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RXMtlHrsRWdmp7wud/3gQiIN2iUCaXkgBBWhz9JOpkSuJn9HbvDwiynCsCczR3KY
cfI839JHdYOv4zo/kCneFiH9Tgfm6nRU18NGYl1F/I9txvEHal0eirLic/HAejD+
CtdSIkTsmg8tuAuLgnd9QkGsEMKE4YoKEaP6N2l4uyMvKJ38fyyBrY/Z5cAR4GpM
uaMyklkIb/+GwpLaChb1LIipgQwZ6Nr/l4Gr/WKq/i3nxvGTId6AlZEvEge9/kTV
LR/VmbKTMsarJweO5ejQPg==
`protect END_PROTECTED
