`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wjnv8T2E4XR6i9M0PxHTRhKm35nDwu1A1crnM/iad6DKyizvd9jfLbH8/MgNObD4
wCOxORvhHCzZGJQ6MJir0WLRqjESZAH2E5AC8uslZPnycLGXdi5vI465PWh+l7Gn
YxlprxJVaeik8KpcKRPMlhog9wRt1NwJN4gBe1CILm4gyhN11rjuKbjIEJLGpJza
N0jlS1Ulh4eXLT6WCBVkKdtL5AxcfPldstfuIVkhBtpBHKFzyVHpHzqXbAYyl3N6
yUfZInWuTwzugvdUOe+GMLPju59uWdyusVsv8628UqfMgJ9R8e3KWUrU8xNBpAZB
kTq1viC15KVkyAMMxs2CPhO+CViqoJQiUhlXmAEQyTT/D2PnWQnlmXLPyurdy9FQ
YWI3EerNFwIZ5IjCTyRWnIElzvZwQ6nwcDcyBGquDMO07WKPMTjrSmVlJ+6tr2gW
B5TY0QImCSduHa9yKOtqT6wz6H7mV/6c4bFt7lRy5sdm5WytsStp8hUwuRn55EJy
GydXfORvvi9Czz+m9C4AsmJh4WskcWushFteoKRA66lOFD+K2z/alKN1qyTo2osS
MvdvJULxId9Y9DyF6AAtcLmS+9dr40Z6K3qYycxPCW7xpmUDZBi/VyyBUNPyc66k
eTFfRF5p6w4sXS3SAzJyyZUoc1G2L+y9A2ZRxi8RqBLxZOOqa/ozm5rPc7DScFot
S7AdDb4Ug3B7rSwry5SdI7xhrW53wNDi//mgEplK3HrauHG7v2zowVnsTkSHccqw
4vm1BKW0OgVjJmOG6CrYoFzWsqX2KSmvHuQIcpyHmYytsUR6hvBwNGvVsIXW3c4v
5dAJdyVpmTM1AI/zSYmGOfMLJ8HBPrCEKlCn/rJdQj++zsLQAKFnI9r3p4QIPLNS
v0/p0e/ePiHlU0e6drUdLE5PFH8TDzZU209r5trBOhIMdyybro3Nzu9cgz3kwy6T
`protect END_PROTECTED
