`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W/mRVpPSK8hKJJekowngANiMhEehWfjFlBVh9Rk2EAGyRQ3ZLcxr+vI/2/fVddfB
ZW1Rt4KLf9aJjHCpspi+WkMfxZYt1k8PZ9oOYO0/p0CxUskKs+bLck/VIaBQU1Zv
i/QPDGyXNHtp06qjGr105Gcg4b4AjSLNmg12y26zhg4=
`protect END_PROTECTED
