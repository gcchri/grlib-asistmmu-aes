`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ml+Hl7n4Lmur8f/KHDANvLkEFwaGy/4xCZD7/iHkjB4lJRjlnL6XEu3ZZ6eMvo8r
NXdCWeITjxv7mSmR3btedmJxXc+2CM/DxO70rg8WL3Ds3/8UzS1KmulQfIUu3LlR
hMmZ3A7NnrqiReNy8c626jNY7ZNT95uiK80yD0PsAbYS1JRLABqndQqsS7U1WbNI
dZMyHqf7QQN+ObGWcZC2hVQBLF9oRv1L+wRwzCrtoB8pTVierWWlElGHVW1BbKus
KDCpIl2bYeOTMohhUK+bJQnokzDMT/yjNEoBkqM4/JAuDDlxnjxb0YNJWmWwu7zT
cI9oSaTKeGZ2IPnf+TOWLrYwDh7YDS8u038HYCSaFB68kE3xCUAsRUoZ1gTbCK9q
O6mMfadh3VfOiip25PRTy2mj6gXL43kWYUh0G71u/Lp9Cq3thXzCRtzeJ8DNq+6x
WeXxoeSiD7QdcgxiP5wqKmjRusbzVH/nLkbBPG4pi2koPrn9ygGzhmPCm1BPMSIr
u5Xp7c98A/3G+kDdoA3sBFFfWusmcg7GWWj9dA9z3kHiGex9edMPyBNpJrq5+cNO
jfVPjF4yOBnet8QrNsTpzR84qTjy7TViynrjS415gPQhwfrAHTm9rpZaAmugJq7D
7kb44npsKEo4kSleB+7PZVn1otN5VnNUM5ReFtHBFGfZMIrYVNbMlDZhehiEJWXS
986Clh9oj3wUfz5dDnKWmLeJh3lhzPppcj5DXPxwTgTUXUOtfCbm1NYGCa7LE5g5
TtPyVpHQmLqbxK3Lb/2WehD7UdsdhcDT2KNRgGsK6VlE2Ir7/yLtGgc3WIUZ5CdW
pRMlB8cs9HFnye2/v9z0f/v0ScR+OL5WraxnCOKLEqS1iOrTF/Uz0fZ2RVktqhM8
klL9sQH/er1fFVcPGOw0+iaqacCaAPV7MqXMJdp1S6EhX3d5KQ3VypBsI4vg/sPS
p/ivRwEXAfvf65LsS4drGHNdtl7W1t81cnmAty7i08Tj9agN5zExehYhImrN/Rv6
7JeBzK0AvgXC83sFdk0Bl12PPYRF28VOvjwcPWUphYwWVxWeOLxKVvalPdiFJxDa
8LpJsJN9ygJtCrJYfF1tDHNQzFK3sznMQvJnTJ4K8EQq2nOD89k5B37qdKk0PF34
xg9io2EAS8QIc+w/JsBbTn7pGtOYB4FjMua8la+ts3GW6n9VKznnGTYRQu2OUis6
bd+c4gbfRvqFDcvijXW4c+ud2nqAypAWpyhu7QukBSAHgerIkGsO4iyblfmAVzzA
Ql24GCuEI72XdDX/GdWrWeirxX7kI1j9f0UqF9HC3lLxZfnoL3kC0zjH3p3Iode0
KMm63c5tBKzRxTQv+ES4wux/zsOtboQfDsr3qG5Jj8U6O2SmUpn/wruRdeE1+KbC
pXbz3epZ07YKoc9Q54ABCmSr/HCMEKvbjhqGetdupBEv+nGum+l97X1o6ZEWLyMZ
FmriHzb12FeqPafcO6VK0dgVi8OaCp8C71EOS1zggbDAfGi5R8BgE7H0EBD+zJmP
4zxIGiQFlOqRXUkKsbsEvy+Dk/tSH+9HxgsV6lhFn003IefP9bxoFeQqNuDLSxK6
VvAL+oiXAQuIkmUNkutmmhgVpkUbRmXfFEkynK3KE83755cRbV+vKF9hQI9VVR9S
v0nvIYTyStosxgx6TcU79gcRr+wjQeg14g06zmX08F1GfL9yOTC+5CKeaBiQsARJ
`protect END_PROTECTED
