`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3FP6zcAi/IHxXa2Paq5IJBeq/30naPYA5QdVFzXufkgQ9qZU2ypfbH+HAJvke8Pe
lqemtbqnmDKcoZx9gGSq5Hi4G+ywINN3izENuQx1d6wIRy/y0YoTrnJNkQYeDadv
7OJbB8MMuPrXZMTcZ6p5LWC8Sw9WaNu5YGa+b+ARBjbzHSxLpIw+n1h5T4Fr/rk9
sO4OLf62/tPkrCMQVHSa3qGTZmYsdu3T3t5Ukjh8eHTTab9qrpMXHQQYUWccO9+2
Q70O1Nx5gEldhz2wJltR7+xpvXtyCRYUgSyNd/5gGCXxXOZXt+Xn2KcJbkcOOb4N
TH0GQ3MhSas/2NdGzUivC6AuQRxULWVVbtxfQcIXMLsZQ1eIvd20hQKB+cibcMbg
ATVNyUwMxzh/D691Hbp1xjDp6CQz3SEK8kOwMliIGIGHXwB5LpAhJMKmFMvUZJip
oC0hSLRqsd2e1NjdfPdWRDaIYsEjHCgZMQvAhPuOfVLNRRkDbDuBXxvLknIC6TzU
xC3yhGCMW2Tc9tXVR31JPZBvEWdaK/Cz1JkY1Imjg5V484ALLtDxepqIz8Z3piny
a+ZTCFczITeKfHugwYYtBpA+86ntK2i0jt1b8l8CuXZULPfz7HRpygU9In8tnNrE
4M1oX2VE9q23iDV+T82XBXkQv7hlahtgftC40URzviRC0IfnuRvU1gdItFBaUuAA
SfsVdssJNsAxI1wt0JpvyNxeYbV3iZAb6NlX9ZKEUoJSsS0Q1+ZEm1F6FhFrOymL
mMTe6nbrvVh+xmX+ZV6cqGabXkAanJtO6vHw78ZYlZ+aOn13BsI3FzFTRNPCYWNS
ueppXrgOc3Sl4TIAQT7MMHM/uJ9RwgyDC9u63nNHdGu4k8bCA2BxuwyK7aBq8lNG
bqpYek3e2DndVXandm0YwdAXdWrSkQr/GIUo2nMMNyzeOvyJrwT7oEnwN9BWNIhT
7/yicL+eRvnBkTN2Euzk5nJU8+NILCQzygQ8ts97/HVxMgqABIS3Q7kN4iPyo6MF
vdjBM9BahlzRUrorhxfZF7I8pNZ0vdmqAOnoYQoqVHnrBipk5kMrWSljMqAyCjOa
JfqnrzdBY4GJtftO5oLZAHMtTAnbmhDh5BcpMOR3/X+DjOnOTbLjbMaY2rSWJvTN
dSS6SCmLZtjiAo3v4yyQWV9TqsVQQ1msIFdWaL2nFRPPukSujKeEDADxI6Ekf3Bn
nQcOTbtVsgyCAn3Ji4HeSwhCbjhaFhkj8eABsbEkXkqUpjKAeN5+wbwAaGLrTdA8
oJgp0+BbZ2RccJItFXybwrj/dCA/yGV7saZ1QFNCh0XSeM4IZwvzURW/DXTTYM78
7WsN/dO2DqEXNHH0l/w8x8ZLv1iRz2rFd+TFg5vaVxtyWGXk32JFBZX59yOne7EK
MrWKI8mDB5gtP4yYE74tkTNj6edOkFIB46Faz1ZO8y0vX+Zey/iCTd9kzUAYZrFC
vJ24Nb81oPXmuMH9ymVBi3RcuvxTV+QdnX/NSMP6eh/ELS6RGU0q5tmMnTJBbd9L
7ej0efdMmap11XfdO1MpVe3e2gM+YRNE8E2MQ9tF7xDvltkZnMOtEb15JPwv4Knh
OyNtweXjOhplayw3tFBMj9UUoWC3hx83JtOmNw47tnkW+gJmqQsBcGl3NGGHWUzu
QDY/m3TlA6Mmfp2j+h2axBW3MS6y4HkdHC89JbGAwKB72NgN3EYC1MNUJc+ch7k9
OSHeVIhhQQWj+SxJSLVJRss/p8qrnQvieCc3cC3UHFyvrQbTx8wKNUJ8aVvYCXKI
xouQeEfzAqLcIhiCMjI86NqtSauvk04ZDZj5nPqmCQ12suwG7/B26aX6uzq0LZHU
DOpRnyYs9kcTYpO3lvEHDewFXEK+Y6DOG36T5AxCwSe9icRNp6B8VSIoFIJrRfTp
Z3ROy8WGw2EAumPIgXGsIirN27E5HpQK1lJzWJS9gXonji93CVfN1YW/iW8SsyPS
Z0P4sX+8tK+e94SbRo1n1QZ+7dN9ioJl2Xc0asMQw/kRKXZ+TlYHzIzlEobbmM6s
z4h0emlvaWutgoUNMbPIEyi/RwHgsR2J0WeyUkS0mLM5YoxdS8w9mXpPRa9Dyzho
i8I7vu8IXRWy2SqQu4W8O61DKemYnU1xPVU2XbDmlNACDrE2U0JJ0uds2Eba0aor
Bx28YDbNhV3GrmGCu4mSh//xDMLKXdgTAxfq3Vrs4fu6w4bjc1Tclrv/94ve9ryD
bL7WwX4nq6JbXaOTHP0hlmcAffgX3E34PH5bTYtd9GY7Nw1kca7NSs6pqhRDWRdh
v4AOuCcmXDmUtcc8lUrIjmf02hPtcfQPDpiP0Dfk8c6cWZGGs/t0MFfCDBBocpZ2
RmrbqzSBRctjzb6j2vpm/poYE6ERbNAd5GhAItKbEWBiPy8QEo39lkf29sg3GLEw
3MFMFEK2gZY1vrkvOER1xGxO+PFsdiPZeKO0SIlytZL1yZndkplLMPexrNzi+iax
dZ+9uezlo3liAtFuOlBEd+prg5dTLyOYORDG8rPWTpF6KgBCt3uSEfxidXTHbvse
AbIQ/MGmVv8lcWKDzSeE/f6Ou9ee4Q3f8nUUSP1AmVpvSwrPl9G2jFkw61OQREgw
mHzkihYkT+eibQbjUxE9y3AePyzzulY0Hon1B1BzYiX9vMiSOPQ5Zj0LsnUj7MF6
8KvkdWTunGjDWfJZWowIIgqE+iZ+AM7YCsTkoTGXnvHU/NH0tBCdrkFt7fM2orEF
nSsWxICCZsFsXVChNPABH2ONzainHXY1vOz7a/sly5jm8fhujGPosOxW7i4u4Fj4
vN2ju17T4aAfQlo6xsPyqWS4qn93+hRP4E3qhc1Si4D6Nx4qQVItpDsV/PjXf/YN
Fr5cMSciU5YmmBnrZKd+sY7+pgqQ6V1HmMFRuFqnKlrYtczQGSTyXHWAf6pBQhoj
2hTiPjm953/8Pw3XE7EbekPR7QrSFMFruR6oLRtdA7exapGNxuDxyEGZZXadqqTs
jSjQ1h3YBBsJ+yy+VJocxqPA3cbt/7yf9ng/gHMeDa7q1Ivq+ZZhe2lYndN6OxTk
hs2GB7m+Z5NBtWmuCW9GFam4K9nRsgYtW/IpGM7TkGfwEjA6TyEDrxHLmWoqJTnG
Yi+10dIhiV3OzrJeGCkRDUEhwJS5cnHx2lxEc8b0GfqYqVMi/vTGUVWj9v+PF4JU
C938zqUfweiBFNxqO71KByTIzUE966svLFeM4URwoA0dKp4fLSqkqLfsZ2hVt54f
SuA6DntcJVKzuQMQ+MTFM7677UCt2vE52lBocYFiJai2nEZdRPrcs7bONL2pcjqD
jkfG6nqpE44ftOfYDQV0YIeIkYdKjlgDH4lLtd7bESsFcTICxiPLHiSTZ8XIM7mO
b+qkwSULInZw/0Do+ufjzddAq8PqGBirYxu7e3bnAJCsqwFkz0D4Ozbf7s2hQFuw
zEM7WtEjAcE5kXDdCEhIea23VFhohzoue3oG/YAtcl4ELaBNYypYUmpKEHxbYg2E
xseTQJk4kP8YCoxv4ywqCfJ05VR/lXprY1xZ/3FVYs3Wbn7hhjtTUMCDGLRFZTBm
HevDqeDV2dLV/SNto1d2YwPKnFL7g+f7rm1Cca3dXYSdHgh9uvguJMQAKdTnm0o8
d/x78zoEYiLIDlwbH6+Vv9ak0UuzZtDz2l5Z4TMFsnynrf9Ea7DHPBeFIclKQdZZ
Jv9ZCYRcGuMeSY3vPqpQdO7kT59bWDPWh+P0d2gHFQ9PCAkxQ7BSeQ/GDO2Kwkr4
Ul8SplsNQ4xSqf+x6STmLfzHs3DRaeHRyN66WPt9L4zlFFxeHIUpHvH6EzqL4s7C
KhZqkGvv+7Tb0JxQc1amYnDyrCrzkSewfl7WOa/C5b/Qh2GEkGysqiUPrDjc7EGT
W7iMmDm1Umbhx6EvFg4rQaEWZTzHVHXh5sKwxDmYcO46Op9Z583YAeBmbZVagnOy
mSg1mKu88HTMMd/ivQyLDhy/AEkw6OfXsBvVBxTOltLmBVJ8k173VmJRpEiSfckZ
aKkpWJx4CXxB+tyPFmNfMH9kRsTQjNAmhbhgQQgyCwR3sYNLLdMKvs2ePZcwAt7w
PO7lLJDwE3jUAHKdslVYvd+r3Zo+dUKatDsjdC4LUlOq79w3EU5ZBKuLOQCaSjA0
DRAGtxmiW+M42lTT7uvGp/gF43TmasK5jZZ0c75jpSLvFLGmJ7kSTBpkx2ZQx9Pz
sfVT+WqXf3Ki41DjlpIWm0dcXWAdP5tepIF/BTVBaID7bu8l0iSsgQtbUgRoliOl
1iRWVVz6BDTCRAIH3TYt/yUTis5B9UREmHPDToVjmsg5ibzTsgKooakYWXe3pLrS
G+KJpFRIoWlpTewHBQe/8ApQY2u7GoiaxFeWfvubFU/WUSRXXoeHYcOtkjkE3LsT
ofl1rJe4jgvqBJqd4vPo//AOjutugJrh5Ixyx6u+2V7yvKK9QPsK9vk3+yGXWFl2
7OGT2mHAUmYXmHkVOA3ED/T7aGsN1uSrp8hg4Na+GajiRLNozZtfTPDyhXjyMteS
1tGEKD/1eMKzG3cdLqjWD3pMS3j/jznrb6qmxvcUDzAsP+8WqkvLoK+Ap3JFiJCY
jrZxL7ZK+Zmol8/UqZKGETGb9AkLyglFLUoZjHLYOH+vlo8fzYRqcYrRsdyNg9+y
WQth6kWEamoc/UOZkAoyxkswoTo7HVCfild2zKXEURWV+hBjAJps1NL72QrMctvT
oEFKkKNHMSlQNbfpb0iYs9AaT/s/LyK+iSqImvHIl/0JquVP+hWmFl0usC4etJTS
xX6oSQrITfuCDxAvy7OGW/iGggHkfsJYdCCnb+jWvg8K7l09rogxLZg4IIAdsihW
B3s4Yvay2OUcF7hAKZMdB6WPxlc2kGYNH7SA4nxoSngzT4KhGqT3gAoTMWq1oGi+
RTzlTWZbD1lTo1hQilbfoXy8MMMa6yZvPgFhMtPeLlJFQnZaMwtzLqnK7miLIqtG
Zc/3G8WTMmvDlA4V5pHQIaFX2hOe488eprsf6sOXRtoaZa5UyG15g4SRSo8tmdG4
+Fw98tCS3YUxe05Z83xgFF3fBsmi6P/g4zCO33lWcjJJ8FsAW+q/DqG0oGrLTzi8
+65rDEmOcKE4zvqRbdAiwPIb7kngAp99XmaYxLBCAlxtMzKG2GdGQQxP9arJ+Uv5
BFtqH1aAdfF4vSjFkpqiWGgbacUk1Oaf/h/QuHEZ8FehtHP4/eEnrS1Acnjw6ix8
cVJQzsuxVzH5eWgyN/kv+pCQfuodleBabcOQ87yposcwj74FJwW2gVBalB6MRoR5
gYeRf3GyOZ2f5H979ie+Z4wRjYb/ScUtI91o7GCXKsHwJz+j9w8UQDCtysPPjrx7
hqV4U31M0MrkzT7nSSxyd0Q9d4a+HGN412VfcOrvSEN/zNQJdQiXP96hM1/yFjST
ilWaLhSVrVzgITyLe1ZOkCx7+Pc+i0J2M3mcG9Vddkkb4euarNGGwN7TFzplADwR
kRqtZaULYF2GMPCz1ASCa7Z7ElRYmKltjEX1zofRjthVuR8ffEmEG8wnqozYiciP
2hLIIX/bqLbZNqI/sXy0nkAdgRLKbcj/V50aYV2m4+9ZuAG+AYb6wHzegk/NkJVu
NTfRrn4KXwKIK2qrFZ12LiQvImMqR9Cskrkw3XwASUqlYnyIe7G5ELaWrct2Tcsl
0GrhXGVA5bo6aghqvUOcdUFAc393xL0AZBmxE1PPCn+QermZc6pR7ZWE6WTF3D8a
1Zj8wZsa2UfllNBUMrK3Dye4MzcDhwsX/2gyL/B8Yn1+yrQbrqZts8H5jgTmnB+M
JZA6CCUcMYUr6ACLwuDwysgjEWipduvGiI8enAVT2s97YoYB+1NtPWFftDXqHOsl
MCOiwxmGbQah5nS8k39rDHkpfupAvtAa+S1v35/11NDWObnLa3/J4HKPRfuFFGJx
HxxKkxvkdEyASw7nvMD0FjfaHLtMaXcmmak/OICYbWOJNNGAxTD7Ineifp6EcNUy
KFJSNilixdoV0Woy2JiXYauox8pChRc8NTdXU8qUf8ujmCwaE7Jw3SY6GnTMlODR
e1z6in5bq4wuT0r3AS2+DdON6MwU+81/uOM2+D7CYAqtVLNIRVCyHi/OxHezdtTV
W4aVYwRhpqNNHbiFlW8QDt/Q7eeomkVgHqgMHGqahDO/oHniWHxFlgA/cPDz+Fmv
xDhw1e6XRnUlhnOXytdAzypoeY8RVw+e7lBbxfbvzfYmMB8ZWdyO4/7XHBbKgOkI
IuYVIW0LIvnuwM1+OjbIHxuY2m9d1zDD10tSL8wYO9W5U+k298DYGgIrw0xkGn1m
XASBi/qMNNfODPW3sqNT7/xv6yVUUVBMjwX720wPGcCV53so2zTZmY18C6t/ax7H
H4Vmtastn8Cefi9gs756HrlvbWBeD38VkF+OX5nwo6swmtlZU4cRKJ5Y2L4RoF8q
rXXsgDQosPBgT1L0Wz5x3WcnPIijw02rB76FPFEvu7/XYmQktCRwmGSbJHl3jo63
OZJdOnQMTzeyk1dLvVPWwwbaRd0Jvi1h6mxCtaLR+VPDe5VQBAEKnqfGS+Ayy/hb
mNGdUzdm6jRe3sJmtj2adiCVBn5maJmRUWpxSRmNA7rftzTrqNgl7B55kRaP8dDM
IHZbqyV98hJgqNTGKD4E4g9aS0r4l0BAyiYt2TXL4FRQnmdCm7uh3W3tSI1nWz+N
KClr4CTOffFatS/LgBnklqW5WXvD0DskuUvY+RB1+WMjfyKHs7kLgP3Ifx0WJDNp
fr+yXIwa65HoaiugYVbPrWdBfAOekNa6K74hBYcq5Iy8eeTJGDtXvcL0Na1JL1MR
z3XGSM5RkLiMRhMRHckZapjJ8muJTWtnFi8JOAIskmtdEKmC3wyo37Y116+PEllv
oPHTdBXTwJWGUnUwiqDFBgpWWNBkjPxVG4fYyuwEn57MRX9Ct9tg5cg16woa4NiM
H038DFEPgvtQLj90PpIr2DUNuVA3pEzFZzbBNIjBLNyBUP2EpwtSLqDsg+2M7swi
L+Q6QhKQfIZP90MdrhuHUmac3Wsh+swMuTX3/C8fQIQLraJqIn7V3dKTeJhASyuA
LEWye/Q+vofYbZqxnGw6LKkcyxGhTdxsIAYbdmMXU8cBhIJh2el5rD/eEd7eky5V
4uqWGjfaLJJsaifb1vYGFXFu9HgQrKnhVo8z38Gn21L11QT2fcYADHFRqeKGN+Xc
sh6MSCAMMMSiLXhYdg5Gg2Epmj4YPQUkq/e9EiiRcnWK6tSs8HRgBevltdvY0NQ0
XUPAuc35TSWIW8+rsXwzixEJnN5znW7sdPe7zxr/luidkDQbUc9WRtzFe2J0d0vp
b+TkpqpVErzPx8rnPcdO6eJ0bXcrTp+0liI0Ff4yhVYtgrEdzmY3aQwa4kiByOad
CRhMqdFtd4cQPSUWdEN4fvJM5xhaoW6RkReGVl7E0kP87fJWKWAPVaKqJK8os0VQ
eZu5G666Mq0Fq3+956NR0Xk9lBXad3NirHQTKgtiYw8gD6CamsMtKYALL+LTroVU
k9B/6X5NXzlvOWTuoXu+UwdvjHuzWgMKf1hmzvn8A9u5yySQKRdZOzJaoa7Ro6KD
QEqcsS/P9OzDy6iPxNkyul9537g1h51xBKacXxiTmPDum09rAcrlui+9mGfslRFd
/bZGdSBJPEq8T8CIHPJ4/eJkjdpTVNpwSps7FdL7taRH1/Yu5Evd+DdynGPhGAzP
cXKYCJVNfwfG0a658qzviuMjaGxZLafhKhxIcoytmgjH2d9bvPpixbTx5kIFBYTh
XdHbsM43ycMaJep5853OrpISk3QjfcHzoBSjI0kpWhTx4R8CUiDpk78WRXysyqRG
aFX04T4TR/1g/bJehh6e9/M+gxqynITqT8HUR/JJ04I8+cmO6YmgFpiXydkJdsfm
1hcal81vzI1I1OQKeo2g3XHXv1tlGdBOPE/v0IKiwgxrMyGpuEk5nKp93S8/fUng
ONG/ljJz81PZ4R9yJ0MPyA1RrubwjLmuLcZ25ha88g63tlSSfWwsKOnr4oFlVsSj
CD3uQkEgPWE3JZVDZalZ2Wbc9vaBEZ4uWk0CIMPiUrgEdMqYIsh+qVtorTA1poAe
ggtEBO0sUW1YMBY7WbF5psaQ/SxsLoyLGkm91fLT+12l6VY8ojNaVQwvVVxOSESD
99ApkcX+vy+NteEoJ62DU8IHnBfnMrIsdE+K/yFalUab1NTyB55QgjmhUAdsd2Qb
MZMFLvyPyuvF0lDUlRJ/HrjtFhY149kmI+/rku7boSqtwODZh52s4+KUWThXz3wx
wYjMhCKkqSkZv3U8JhKuHZyGl4zjmDpQFpThm1fpRUC/o5JJAOMLLUxzJnCVdo9c
nCmdDJFmAUvAHwFI1O1kNfKLisZJuTfhkU67LWOb1meHknQK5zkQN3mxX34x1n9E
JRnE6vD2jvsUjUZ458zJVBs1i4xmtqwvhsrSsOgQADi2s9rKt6qdrlcsPZlyMibh
reqyGhYvyotN2c4rVgRBsueSWh7zIfGBvRWDXUAwGp8goR9yivWxDY5Wsc8+f8/h
SOYJVynhOoQ00guZqRmSoKDDOUMNJw6mKZiwKozYklF9HZncvz34UdLFA42CYQ9o
3ISCYxwUrvncEMo6M2IRSelLJBIxaVuTcRCBLkzSBrFvnhvfygUhSFSrq61BMv/q
2kKxAHCCysajxXOUtScwhIlAhKjieeQlJNjcZgEc7oLwlYEx58Aj5sQssNtokXyo
w2/f870Y+QV/8DFwY6CsmCxtZI55YDSWyS5dDxBDFaZeqh4DJ8g5/oTXPZNQcl98
FzxVCrBvFn/upIl+WA63/kliG7v/nFz0v826BtcxZQ2CO0H421lD8qole4stTue7
Fps6S0kDA5LAL1PFpdYpEtYWsa6syksBbLLjWtiPLB9SRoe3+VL0WdVCRmTGvVho
6b7j8qRj4W+31J63z267AzuAlewtcarGmE/MHA7fxBMXMD05Dp8NW4/YkFHOOD3o
fnVDU+Pu57jcXaNjwPeDYyWxevfJ54cZI5A0s/V3aDb9GsvpvGmi44K0bahD3jXF
4xG+b8v6fCW0J2gDMARhlG78nxEkJDeEX1ZF0SFfql7vTe0XdZK7L8vq2OkNLxGO
k6zm6jelakKtXyxD3IlRlal2egxmPau2U5CzBF1v2oh+OzhNisRhOi+0ltc6b8ZF
c3rH+rBvuYL4TciJuS5PHo8QuKdJrcn+EAWFgncEMhsmQaanAoiuPT/tIPY73MYj
d+qQTNeKwDS5++nMdpzryeuX+dPSCM867XcHlHof5CWNoNOUbaPmiaHN8QkywmsY
UowK2mFqGS89tWaQm22QK2Hk8FexkSgM+hT/OAbHnelcIQhrKVYvCI3aTx1YUQc3
6b8xI3oW/0X+8S277PBusMRLWUFCb6MfDm8LouzTGvX0IkTLqddUT3cIsupyR9lS
xadN8k/H+HHJo6UXYYyqFD4dPhIMgdVLWhu/VzGWB75z+ytzZLNPuZJ6o0Aj9diP
8aRRn5zbZ6TIfEoYIisw5EX4Ibun1G6LQ9i8p5fCGgFi8jlpJoCMF8ONL2vmGLo0
63ckEDOAN+9AQbRa8NwrPbZhTZwpoF5KdxIW1AvTjpocT4nfFqgED2Y7jPFXn+vM
jCZnRbuF6LHJH3QVue97Z/beMt8iWKOqJONOEyGHYHfZSNgxDtn3+XfQysli4S32
06oTKHN6J3FLLS2r/w6+WJDTgkGIiqRyYeSrX6UISvsXZ/0zESdgCMoK8FtHByEN
9UCfNbVlx2z4xkQiT+3nhNRoDGvQGJbRNroTQBJyWvf4InP0wMRAsrmSn148kUm8
9BxAGm9GAYCUMt8DVixnjIii2zfxYlOhHtrmsHnsFxktvVzRXgfXIEy7lmugQoi/
h2PetTkKMdrUXykwDHDZ9U46gVHQ0DwFKUYPckRK2ji0AT7FAsHdMqnMvzm5nabv
Ao8gIO3ddzrrGxv45zd8HnqxJ+WN/xoOPmgRUFtZ5bttFZoq1QvYwJHS5U0lKxHg
3O8PeIfTDeei3ivXSuJKDDTW4tv8rQn5zDLvkH//mQTXi/pyyYdyjzgohfhGEVK0
WSrppv3nddLSOOLHCw32IF0Fqkk2EUylWkFiE207LkPjclRocdnQDZE97W3PM/nW
R25Fmnxx1WDjp0LqXK++yg0Z+zGg5PzRqJCMJTDDfe3OUDlvWFhHBcY2OX+Su4Y2
KBEePktgEbVPGSxwCqF7oWXDSq/qrJ4sYpOQvnX6lf5SYTtr9tS5V8dYzOH/Cvjh
XAJwsAUpJFs+c9+KXmF9A5T5zGq5DO1zw4rV4mSzDfTXFv97PFM90dpA9AcmyjPj
KEl/3cfi3batkrvCty2gSfxm+K98HwpZ4Ce1fSPEzqKzVj2yKVLyq2TEKXEB1FSq
68WD8n1blcpLqfbHnb+F4uweO+q1CjTMk68A00yB0Clt4AREzWnOKSU+6hjrgo+a
ECU9qoCUMUEVHZUPswHYCWHzl93TFjmK0UsCeNAbG0+atMIn06cz7PaLERBLXlud
n/Xv9geUR1PWFjhc2NSqXRf02JSwWxc6vFqcCNH+x/PcfUOczvIGlBpqJpofvaHe
/aJkbNtCecc79rH8hqf1KdnBqPV4V5MBYI9h5PEdGnJdEiLBbziicyAzKZ3lMw1A
Jn6ZCW6aoGaPP07xyd9gkt/phvnDQoxN2Fu7t7loTXAq3yKXC+OfezvI+IflWlGx
as6tsmt/4mt+0yYpAzIZGfXeqWXbHlMj1AShePd/ri2GsdG9xblS0TSKIT70YQg1
NmXrw/k3A+PYL8VTPSF2GA35YEXbMnjdz3jPqE+/PJAq1IJ2fuxYqU/8TOqv6CIu
D3Uc4Cw/QzWAjglXEBgD2yo7JVVDUGDe8ezVrV8FJPYTsGKHD+0d4vDVjWqJtFz+
DBVYffCFLiYsMZrWLBOaWxFRWE7si17ruDoxo8Q5uM1n56BH+1LIO0pYdnCMyREo
n0yean4LRklC+m3aAVUTCLR4WSdcqLxxV6z3tdCCVWLnrc22KSGbsodQvzbpxez9
g77Np94Vv88ZeaytPALPadSJtlXZXdHgAb+eqQt1M+1WhSjPLXgy9V3sQY6sZcNp
2nwQIeA3HqL/SEzC+eVFHwGaHCcdqt6tpntNHhFmBou3YKcvTDMPtQDEuT013wOC
4e3j6Pa/gS4KSPVASK796RALWmPS5oatKI86DRkO6+pibVpjlJsUYffjdnop80or
VzCiwp1Q8M7DVi+zb3hoHdNhrvb3NGjZ5GiC1HKLhxZCe9NAaiCQxIDVaDNAiL1e
rEJRlkUeLN2bjVgA+s0B3tijlB52TBIs6Pgl7AsIHacETbX9GVGe3cxJsO0zV6Ts
Y9IxY60VfWG9ijW/lbZ29RsZgdoQ/jrhn6D3LpasN4d4vxJjTx52vz8SqMe8KUtU
17uzp/NCbqqzabzgOV09uOxRJXlozuPXuWjsSW0cBgBzUpV73D/JWxpM5AwE/K79
uBbYZWGnyUBeRuSEGP7UFbkqFnpQ6duORNSStW0e9ci1XFrUqb4EGxKTkKNwMQK7
JfaOCZFRuHRfE/G3gr8J8umu7zA8QL3+cvmuSuK/GGtJp2Sb3LVWE47FOlrw4kYO
rK19qWeaUVUBB6zuz3j7nKdG7SI03sXmZtmqtXypLJyo5P8ejVenfWK6XaGv+1QF
n/Kozh4zmZxHyyWZsSnBpuAofaUxnxUhnOLW9fUVFnpgE+9Iz3LveF+WAFCirNG8
Zp/Qh7hLxoN/K22qonYSf32kbbbC0nbQEu7VrKEHmwwiqv+HVkWZklvBEXNvhNB2
PurA2uNcvb9QW7nmQn4Uu+WCdH1uYo9ZRHgrrB8YV6ms3wJTIRpNPKDe67Z0D75x
fGLawBbJzY8YCyUEEZTOpbWfItyoaukt4UekwgyxdVT6rUISVLcku/d1UKvS86QG
F/h1X4gi8PeyGrCuHSRhEYv5LV5YrV7xl28lpBagjY1cx59oDJoRx7RdTpDPLsJ0
FJkdAkK8ZfXKMcAjc8/d8NvEY23USZ69HAJzpYxNEvP/LCGCfefPcjpIg+p4Y7Ai
GOMqvnah2HDuWJh9bj84m417CfrOK1wgK30TYTZUsJ4=
`protect END_PROTECTED
