`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9SDueF3jMpt1xOWOPO3qNhzp0GzDfyZQ1Ul6uf9gsE+NGQ4pooHX2ykURqXWkzuL
OS4FnDC2d/OYQ33u2lGaNFq4RAx2hxM/r9mKJ6Ek/ktVQObA7J6HWRfsLPcbdqIO
ML+0PKanHM0cUp6jE6PWSlwgpQIOKOrMe3/13QO35hM5gtOzXx1WnF2RSU4YuifO
RRZ6UZwuunB9C5grMQQfCvrf759uCwQrMEv8RaiA6n0X46WVEs98Ok0ZgQ8xGTt6
MIJiH12bXbVcGeSKIKLbgjgxJM4skMtciC8ZFb4Mj3dWwmQaBbDDNUBC8o71L+Np
ilVpEO1Ht6d4eMr1L10wcSKjCmv8lwSD1yeQLF6Q7CHBkbHpdGDCcoYcofGtooDI
KMJUBIuUjrgYU5ThCBDmUQ==
`protect END_PROTECTED
