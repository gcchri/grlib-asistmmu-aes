`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
poQi/pY9SZtzeCMMbp5t3WB1vmaH/PcGEp7hzmZAwmUvejne8/bdMGrMpZw29PSr
In2eAbywGwr+57XUEb2vOVpC8WbCcoVR+5OYpKi4a627XWqwuTyT9wuQyFpR3I3c
hDAdipXu/8qp9BVM9MjyvTjbVo2HLfg8zn/Kvwe51TMs3PI3LdasVt18V5ooTtE/
e9dKYe3zjW8M/T8LBZb5sRggrRAh3hpP6NI0fnz1eC7U9iKTfhuEJ9gtfaCaM3Y9
itABR+FMm8mXMZRMc/mi0SxMWFSvPYT7QhYhLZCIg1CB89Ase7grRRsQBSM5Ii24
2u5SMSiEhCkbU7lriKfrSYgh4VsFyi0Rh3aZpj5WVnnyleKtLti+7AX+M2aySYRP
GIst790LOVlXi7DtO8OfwF1/UAvWbzyyCQHW5NsqXI9uwF3ASQVTW9sOMQ0Gaiav
nCkAmHstR7NI/FsczAjsw5wWK+nbBlVnCfpT+lqJjEVi5w+N4pjRtwqfs9IruDGz
9W8qp4dBIk9AARJL9GkLPUtvkcc/guPf8Vw34//0RU3BlFdiJygdHBWBk4w40D6W
nebgin5lSbT8NRJEoCuABZ1vp5ZkqzGKVuzES3VFEfyUFuxi4vBrikWzAi9TZgUd
zAo/UJ0xVybhqAnWHtnPilPzpFk5U0+5EKW5UNrOPNIM+X0UU72nGwVKUG2RQFOA
+5Z5PH9LOOvPKHAccxW4TaGs7XJohOuICywjgyYzuBPu0aL42ev3K1bs+jWfjkqg
frpatu71cS4CVga/fbyNTHfn6gW4A48EovwReLZ+QvA=
`protect END_PROTECTED
