`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1FNzp/Hl4Nk38JlB09eBAmk1Mtx+DYWCVcnVLPGcDX1b1J+h8e7Y+G5UoXkQnQhi
bzIUHrYoRcm3pyHX2aOxu+xbyAEnAYExIeo+nW83iEN+AebdnnR/jg7ot2tG8TQZ
5kXQs2fqTygzcD4DEM4QXPseFiTWWV/gJFJSOyrNxmn0UKyRZEDmJh1oVwfj4xgp
CxmLJdTeGikPxGN7hG5biwMz1U28pkihz/hwUQvedGuyFM+Lv28QNvRZWHYGK2Tj
OtKU2lA5saG0cHGIDW2VOECzAWt/b9O/xIQhjCYlXg9u+EDF4Kmr6QPKjf4UJ91L
vl6ZH390OWaIFw81TwBqG32O+bTeZ57ImBjd4rC3YFVAxRMjbf1ixKrNbM3L5eja
fN/3LsfYVkkhsGNHkUeoDkb1AVy5vlg1eUGszAItLmj55tl9lCYP2ueInCWPMVbO
zXFXVmc8+FVlJY/mOG+xpg==
`protect END_PROTECTED
