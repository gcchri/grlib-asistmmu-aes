`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wlwvRCsaAxBj0LEeSXrT4Mo7LQCHYYekv1lXlFsTA/5x7jAaiH6hhJb8wwi4r4xg
VpWuDjK1YbwgIHLLOvmeOqw6H/Avdku5mgPXlZZ4xfzjAjWrw2FH0U9lbmqi0GzO
VzAIX1JpBQUAyB4LEEONgkyHrBaK9xMxnol7wmzVOzvwD9w4ig9gLYhU0FtkUQMb
4h3kezhCnwyIy9g9BiPrhV93JrWE5iOGMNfkQqZ14EfMxBe0Xk1NexUQWRZEYT8O
qnye14ezMMA+zW+wLxbE972TMow9DygqlP9tDsV338caKVcThGJLxGkalYkfwLax
rQDQf3X+oOQ8JJv4qvNyZw342PZbwBu20MlMnC+Cwd7BcteQy5H0g9zcyi/IdlIp
5Qa63hhGbuL458V2yIAENSYeZMRCHxkK48ykTgOWgVCePsDH9JJGs5fDR0OVrHl1
Br8WWLUORam9A6wO4d+ms4m0g5eI4ROGimKm5b16vZaQUeSriizT24HjkQQanQ1g
9QId/yNOJD7JH/C00K7fCV+rhCn4cjc6nvsvMaQa9TO+4qTi2eeVThY0bQuPQiBk
ikR9sJ8GDYyeTdKXqoFIatRQRzjtuA2uyfcZGlK8cLLjOx4NFwEHQVBCLkXDbfb7
D5X7qXjCbsrAER5wr4w+NlmJ9zzilVoLs7oEhgvx7uikTErb9QNBKciUJi+73u7C
wGc4mWlmBwSHp/u3BoDpHw==
`protect END_PROTECTED
