`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V3OZuZyNlBOR+jpBb3RntBPPpBEQYfsTpbUm4fuWneIxPkM2g0lxLZDrETC0SWfX
GeaSjpNVTubKFeM+BcfXYGt/ljOk9GFc45gszU4ibbPCzEPTCYJlY8rVU9Z6muk2
TCwipAraiKc8hzORIvbuXGiXcKQUtDtswqFk7xBtl0mNqdrD0urYFmA5HOuuWr33
U1XC1IG/1UBF9L4MD6qmJ8JtjFO3TQDl6V1yHVENpBzNsap5mHMZYKFW/Ki/WKwT
kSbHrjGy258iX2furb5T+FaXWCck1VMlByn+jDuSCQjF/aRGnAUnb9xWYg4E+BwH
ct4O7cnpZHRt1b+PiZdBN8P8MhRNfUPvBNaF1T1Wr9ZDN7MFPLyGVz4tzaqi35dU
0RKbOPGtuWDO9aF5XEgH2APXMI86GftT6zjocj/MbVyuvTU+E5ArrVOyky53SFCb
tBwKquGuYa+IPDg7Cs2BuA==
`protect END_PROTECTED
