`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rSxTlj1GC9nq6rt/gqPjeloCX2BWSd0UxoGNTRcu5AEYE6itDp9iAfEMTdtNJztn
SJrFUVMjsisYSDC3ogC3eAa12wOPQ6G/5jKl3xBPAjMCphzjEcdZbX9wGOSnsuHi
DzvQ1IK7G9qdU2J+qBhA5FUK5xiCBpmANTVF9UdqmslZPAb/a/NBY5wlXMYHJZn2
Sz1SczlzpK7ImYFF5GJUAoHSF7tpD3uPF1752HFcLiiXReES0mAjQpoLkQkl0SI7
H9OhdoBvZVpMoQUWYzz9v/6iAQlvodS2D0IHV1xT6elkgwEX283vroMlL9+kIYiN
UFYszHCSnpDHr064j2JPgnodDeAKT39nhDahbInXvqYkzx7RKtNjiKAF4CAn5gyU
VI/XTZsSNccta/lbunzNi6Kgs1iGjUoxy/0NiSXV7/N0Nd+n86ra19Ev9AhytNSa
3Th3cq22svkHNX/RITiMKqmvmyG7tjsPKDmoB3PtlprJA5EjgTQYlWIeaevxDq4E
iUoEZZE6P7H3LPLbop5lbwkHNp0x2QwgwDdl54DJyA271KD/I3hyCVkNhHComofH
DAjztzApYcBNq+vs1Gcl59I46U0ywv0RQQSE+Rg1wPf5Rb99t0bxa9sHTN5B0XJB
3FTf/nOxcxmDf9N6JqiThw4DvJ8u7jo2TqmGRB0MiGCNRWBXeWmu1UDNghbKea8a
wyZvPh5b7L2PcTBDJJXiwt3kTYtebI1IWu3Ge3CuMlFwUtxy7hAlLjdyVxApIvDL
8hNRID9Vxy61Q/tbLJ8ttpBYXtEvcQlG5/H8ZwonkPKaL2Ou0mnakXdo8/a2oLJh
rZUi9fXuDKzbriiYL9Z7cWjjAGFNopy2yaA/gmgVG5NosCi7Pby6Zi4d1KukyXF9
yItWxdtz2OikBkeJQC4jRTKm1+t2tEHoufzN+jAJb7FUCS62pI26plx/Nad0Vao/
+Pkn0BGpaQe4qGYSURuJoWkAsA+wjDtobM1FuTKX8OKCPJvqzeXW8T2nNi5kEunV
Oqw+JEoXIL1h2IwHcQKQpLdH4pCS/9WKUxpedPlvBn9OjoSXk9vt7Za9Ev1WsAnu
KwUOR86wUrTw76NCnqQYspr4zOGLJPFxek4cq2YoAWnYXqoPSeeab11I1IV9J9sU
OMyV6MQvjyIKRpXYBb9LRCyzWJ48J+BkfvvWnonzJABrLVvMU5qP6+EaxldE2QsZ
tHv1OlDBLOfMhL8jZQdwNPiqlqhn7ZoFpkXWzUQCp9nqLnmCRbLywkLK/JFUjL4D
yX8QuzZAIKZZZVgdZUkfBDtG6iFinMSy2ehsAZemvyj+smuSmfXNyQ1KL9Nfh0s1
nyx47lhV2oqpI949DeqOhZGPl4jVpbrI34SuoGZagnPlQYZ36wzmEuNXucWr9e6Y
oxsDeKAHfwLlRTQ5m7t1PsUzBGamWPfEU0Wzn6P3wuItt5uzdnGR4bhLni2fYMns
+NuLMB8i9TVAF7xhxGTZSUu6PQnkd5CURTDLh1yq71rsf9RHCQiYdrEZDD3YwEky
Gx1ZUMUvdsoTb/BnhePRNMEM6ZqtJJExqyZhhZNbveBFS9CkEumvIGQaTAH3YZQt
nDd1xc3ibHnLJGsfhRJVkg1p+Ypaq1hqTY1MMB+PStYshslYIcL6IUE7HzPBScyU
TQYdIRCaRFOwD7K1tvwUCkc69pmNKfVRN5jQfoDtwYwXWvXYmH42CP/oFFNOcH0p
C9E8EHvbzbsQlVWdaWRHwIlLmuu9QREQxmgUaVTTmPvNtH8Js3cPiniWDzZZ3vPs
QpCpHQ63ZC4dLSuH1I0ipddINI8NFA0oyAk+Mh576iD2D/9M1kn+p9vP4ZSr5nf+
PFujep/6Ou455cQXcZPUHzDNAQFaMysXlsGb7bIW1oN12A4twM37OobFIZjAIM/7
hnHh5mPumpZgn0CPItwG6YM2mr6UKvDS4z1LxVj587aBVTYwNf+iwVf949Af5mdp
JyCX/S3J9/7F2+p0lj+oRokC6rpWQq3iQDxB0pWqnz/1ezRrZ35ySUBcc3U2JpA/
lobdDkpWPll13zYTlIT52+nKCXMuCdDRkI/JhzlHNNYHF/WS+/BYJ5UgIXmj0vQI
imYOF3TAQRSpLG9yqhjlMOQRD/zXbzavp20snaFQPvy3VyOHzhYNTmd/xf421Cxn
sC+AQvI68bnFWdGYCxpFvJ2RLmTWCWKPy9Lthn7UMg93yBrB7ZMkrYkDXHIl+SG9
0ywd0p2kYL4QfN6WffAeylSvj4QYjxUbpB9R1dn4ChJJsNudrAXjqx9IOz0BC/q+
s5u1Ps+ji4X9FToKP3d1IFLLMI57dVNQinEheAJ/g9EbpS2OiO7/FD4BSyqzKZXU
4PO7973hnCOjtiXbTz4lSwAwcR+77OKp1LXmj9gb4ialict7I2R57p7Y51sZkm9z
dUJv4iHouvYaMmfprtUG4uhIi5lpt1xldePNEmUlXoHQu1a8geOqPqrB8mgetA58
7TRRTwFVhiG6nTuEasghWO3cX5jPE7uyzjJ0dXlKE0k0B+huzYOEQcHYe/f921ql
e/TvN5etL7+I5DX8U0rVDfqaxqf6uBD8rF5yDf4pA11pd764wnFRfsA/3yrARjNK
XMVCiZuo6H6Cjuh+a1Cx4nUQv1LOfmEg5cv90hTWNI7H3wtCrH1uT+s4cfbzJkYr
zwuWf4z1V7CGVnCNHrX/NfJZi9je8bwZLKCHl5JUQ4yfez0OTvhh6lVG6S+3Hgxp
pzD/GEcSyfvY8Sj7qFuY8w4Y14ZyYrA2VSoTQ+m0iwkL/aWvbWqOMyMp51ZPf5x+
pgCW94sE3/CA5L8L1YlWMxzFKW4CS1rFaWLGGxpsKETbZFrWKkfwadiA6p6pccAj
dsE9dtDW+67AfUmMhPly8ksO/8dWyRIzA/naNB3bkIH0hAyLDn9jEPLou/e8AEe4
z7JiHvJJa4LCsCrIAHrpmQLhMBdCZwKa6Ysvj9DaWhFmgdxaXq1svBf0wWeu0pvb
kMdrXhKABH2RLcPcpYqF2dZ8io3wn7o8QPx4fcFfDvd6tThmZJBa1jt/tmSVdjs3
vpsT0AR1PdMFfr22dWTnmEGFCTH6CUFc+Yl7d3ZkLBUEkEe3AqeOJ83zivFAM30K
0XIE4qFQngOQHlFb/wCE0YSv7+GQMTPrsorSPyUl2HQGKqoisyf3s/Q7uZCNj6pM
s1OUqc+l3SS87Vz01uKfuZwNRS+oUHEZXJreT1Mk3dMEfCviFKPCsXwJNQrhWL9N
iQJOX/rxdBiNtUM9xKh0Xun5T517ZmqSuJ2Pfb4twQUjnuMy6dTCmWMnZMAqCC7k
arALR3AwzK1ExFQkqEaMTkhv3LwzKxHLJ26CxCNVdCg9Gf8ImZ6B6mMu+74jj4ZQ
3N0o1b4Q6zo3nWL5L2aWeuDFlnjHcIBzQeERRG8qy0cMOZvz7lzVeQzWURZj9xOG
a/T45BvQPqmR1a7J+sckJz8BFpo9DOCQaYsphU8eMQJIq6xpuDZfJNxN2hwoiL0X
Hsb3wmpZ8ydFAX0cuMKT4K13K0H2UHK1buYAzpD5AFxUMQzl4C/TRw7fxmztPLsm
mjpYUenWmryHrVEGttO/PbHJf4f48ZnaGvKk2tnKvgEkRw1PbgcR0S0lklh+hSk/
vrfSXdSWHeWX5Eat9bmgvxOTYqbZuuH5/Rks8D/Sn9ALaOeZcguL6TV64IYsqXMt
6sg6gAXCac3mgbcSRJBjzdMogoDb51LFA/Asw9CnhD40+eo0QvrN7ZIP0M+1/Ruf
pd744rtvCubTQm4G9hvm6pljq2YZPnTZkPNJYNN3S+JDQRVBiwT88MWyWWVQ/J+/
1XzkcBrvHTkD10z8slnPBGVHp4LDFC1asaLnPcQmgNA4hUlQpsu4diP9v8U1jRx4
+Hz7Nie7vmVIj0/XztIAdP+bOqefWR6t/o7b8CTHAcJJbfn5k7tbURf/9in8dgv2
3Ldk9CXb+3qZiZYxHh8pKu381lx3yjj2tsdBhjOXe6wZo1HmFyGJBTWyXEJhJl7I
w0HwFd4xPoNvUcxDpwriIm63GrCvMG/2lvR8eZdWe6I6xkk/enAa4UhFx6eco23D
zCF/CmDdHu68kf14SnCp9hZvOEcJk0LoTdLQizqm/4G2fFSUNqqMcq73OhkfofMY
kPyWP4Qq6h0DQCm+AmcdvxVBPVEeKchje0A7gWEMlItuB8K4Bq4TCo3vE0A6AIT4
zVlusYapaFhDBTHYUt6t/cP31IXZFDSkswMgo5bImSzpwr0z01pPBkUhMVYkU9ml
4BLQf+7mNtu4/9K8c7I+m6NprZU5Of5gvuRHqxyZ6E7IAI2gJboiv1bcrVtswAjR
1T7hYba7d0PIWLhQUYro7kgjbfmkDA1eT8PV1y6jKeHGN5dCjnASNUS6ej9K0FBg
mYsD53jwITEeoFJ6bt8GoAJhnMXSip97vKcKiJlpXs9NAs+RTWoqvtd5mp4YE6Bt
+m+nr98rGwO+tvLROw9X4nVkDgnjjLWNrnD+siFCXU+GTdongiwxqNnzzUoi8mDJ
gQa+nbgw2CqUDU51Qi6V6Om3Wrn3DDvXzO4X9K7o9DzbICI+SfaBzghSY74rHDNh
MmeTIKiGTh1CUrpoXzJY5NgkD0/5SWmyobCaMvElS/snDg1Qng1oOqS8VfkzqrLu
zsstotvcFciOs9SghmRHin43DowGiJ/Wqkz1z1Sf/ZqqDZUqZBVCpkuZFdQyQ2iQ
y3yjSabL1QD6177WsQ1mU6zhfYLWrRrZTgfOY8gyDlftOLESkKelghx9PD5vLFVV
S+OAmLSzfubAb9X/e7fQaw==
`protect END_PROTECTED
