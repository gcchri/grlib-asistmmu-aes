`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KZgvToomplnmvKgS0wmezocdvY9RVbMV1EilFevKhBRxRzKL9H2MFBWa2D3vtovO
N7es9UdkJY9c6SzinunnTpoAirCOGaQ6dE+WpoGGxNj+CUCq8z82v555o+cal1Bi
nwsUg/MY/S+MZeLKCK2F8oIekxo3RWofa83bH0CTYBykQSm7LWKjoOI8zcNOGjwt
ArsLoYOxt3aJNjUljGSiFicSrYxZwRNIKUEU+JCs+EWONm1BHiABEidgKxNEmX8D
+KcSZnwpL8FJifcmBz3GQxdR5vTXFFLtLFK9jS+Ni0pDQgtxwAw6BzpLRLMiuwU9
SPKo1dhDIWSs4syAGv4MQld9YuWBdUQ15ahF2GbuZGJANWNA07eT21W2KkkXuLD0
5j85E5bhGmH9KH7qhTslO8Vd/9EzLWtLNEA/1kRDNGH9bHn9W00F4bCS+1n3MXJn
tGQiIIIbuHOP0jpEquVFH5wUd9MBvMvWonFAvFYanjEznnHWhceCKzFSQxHzR69Y
c4hSIS2iPxICx8jUlqqIdOW7YySo1sT1MVmBxz3/oGV4DebbZ13Gj3LNdzdB+vB+
`protect END_PROTECTED
