`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r6T5rbR1jkwwhFH83j19PFv3Qk5GV3HJDn0t30jZPFqUKgz9IhhvUosb59fNZb0L
AveByne2gnIGjFGgwsJF0COGZvrN1PqsZbMFYKKz7aANF+k8PtJQK8aFVtSqZCNS
X+3qIOgcPksKgWKHAX1jtPdiw++jXr8yp+u68VVoGHWJ7p66vtztLCRT0W6/tRSa
dZPw/OMp2Hof2xKbxsjucQD+FAnRtjfgbnANBGL4IYivbERhl7/BQy9zALJBeUKF
HOSaEJVrDsLEpDd+jQBQ1wqX/7JG7aXYjbQkgnEtuCnsFx3Mmko9K0D3d1hVW2WK
fErD1tef3mABDmGMEXuXbtxUPjFq88qjW0L8Su6zny7GPWdZ5SZ6X0siG4Pn7VaZ
Sc2MtJaLqvNrPyiI5R5y2R2H6GNraRFFgswj/T1DvzRUbBz7orLYwgv2YutuUpLM
l/uf4xSwj7QdG6EH2kIOVXkwxVwSUrQvndD1qzm2smKTpqbhmT4/YfR5nrcuNDM5
vYNjCpLYUXjQH4MUwSzgo+Jt5eASa40dvNjSFCk7xmMi6r/rWNkDhb8hM/e+Rpl6
Do6yc+DFGuvltZvzkIzZDPFDITwBnAwVUfVxk635+jPtBRjtuNEP6/cANRLx7naj
VFazNfVmJz5tfo66YNIk9n9hr5o38z5NfHbWroaqOYtmyKEdgujkIVVNBFGBKcom
AqBnCNtBfCjjzvSLzp5DWHhspmQk86ZyHRxvNoDgD8LbGJ0TsAzkLaKFdyGBTKRb
COMyxuGL9aF+fT2JuUqCMyg4ZMf6LFCP8glxynwXXEjllTIb4ney0oZhRft59d2+
moMRy94DA9SVaDsBjOJN5GUYXvkFaghaPE1MiFgN1REV5TakAOHHXJ+GgNvNQvm1
hdJ7RMZaC/un1CAW815MucpevL9meBirz7WB87eesp54vsKP+jLWdWFLxxnCLrFR
gO4X9+qDfrmSN5/Sc4M3lOXq/iHyqo2KlsF2rRJzbaov6Jw0Q6apYJUCezEl62vT
KTG0UuYWscJQAGGrRWFskLqytJCbFN+eAlgsV3bsYxcetRwcN7ICS1m9jD3NuNGl
ofOt0t9UbAaJfOSJJg0w2sYfRl8fNZQ1ZeqVveCittzyMuukku/cx1vBCgpqi8YJ
oDEbzWi2hhCR9+/jl+lnmEl8VuLkZ4dxLB37tsQ+IEHmfx+CgljQx6BCOpe5NHdo
lKSQzIwu+rXhm5sejNy8f4/YpczEibPijCRGsur2twIkyFX0mWHdDZcujJ21ci6+
`protect END_PROTECTED
