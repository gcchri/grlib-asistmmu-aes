`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gdiz5UezY+bed1Z7eOLUsevyC2Y/2yKQavh8rpUHkWP8531wMPehPE0PF1udv7cY
Q2s3WpjyBQhvXKf7EmPz0eiJ/OqPAvFoFVAkrtbdt/v+f1eA7MEBn2hO+JdX8mQ8
Mk7YvgukjVD7ezXaVqKw/vLXhfi+7VBf818Am0+q+Xt33J9nroAMJvFIyd80E2Mm
4X+mwGXeNb3TvtIp/bI7rGUY9icSFMNXiCL1ZaxxWvniVe5URaEoD5lWT0bK4UKa
UCBsMmI/CwErCfUMi1adWiOHFPvess41UrU8wfD35tKy9io3DRCTUblxVIrFuF4W
OtW06Gow417IyniS/MxkI+hThAd0bPd2RhwHQbVrIiNKqTJdl8NXdJNchirulvjb
tuNHxZF7ZJx/KYtzByEyanqmCQcGr1uJUWydd8SnnwKMLuPO/x10772HkQVykIpe
LqpydqBaoRTbkgQbnLr1gNoq3iilTPzLblz5WOxyhw3UKaCIkQ0DoEptn2/i++Dd
OaiWT3xOSQeKZUDH8znNgZUnM8SUdsFgjhZ+dBDac7ImhDE7iU7LCXny8HV2dsXA
pP+KrnWKxhAc9vEdV3u2OqbULTLY6G9L58Vt5zdy/mtF4p6cBo9jITT1GINnS+ak
`protect END_PROTECTED
