`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XNEGGWV9eJvDx2ZW9s9d5uk9/PlrQJXhn1ti8/N6wHLhRcYI/oZexo6O6drpGTcp
mZ1bFsN3gnRMjLWECUEFrK3HBEyTLcGc5JqzNO9UQTNmTcjxJrWWvsZL90PIhMQN
QRlZOXPNMCpLc+gEooFg2h5qN1cUJw1PKVLf2B6x4yreMeQJmZ54wHYZkee9evnt
73l0+ILjC5YucLoN96oo/Vs21lT0XMeYXUW4QGb5nKLlgyRu82ahg732r9SbeBm5
WJrPdvRl3rl26oXF0DndQzwHCaUebfLmaTtUSCuFXPI+rq8K8VvsHBtdmvAcqxlC
nKoBLjF0n+9TaNH2i4GHcftOMbRTk/R9Z9wdCG0dj9aoyih6NB8tOgtrfScj3c/v
35+iFaWwtR4+txlRrH86LgHOEyhiy4cUA941ut3K078Kiu1CKjDZsgoEMm6UGIyk
`protect END_PROTECTED
