`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZKRDoobPrFmIs4ztzdpanVBZLFCWG22V+73E0ncui1cBoAE3eMk7wYQ0Wxfx80AC
mXrL8QCQZwYNwmcDxdinBxsQGWMIuzRjZKRaCEHuyo59l+skyvExpLOe3O1KHvxy
i4HyOKMzg0YletaESW1JNvUE1UOGG0W0ECemc1SMZnoWLhZr0jQ2rEu6irodTDlw
cORIyhxvw0/DcC5SNGKT4k+mVDs+jviDrx0ntKx4Caowfl/aKOrc7nEeSKcz75za
RZjLJ81u0FGFHQB/vxj75WGZ0+ourrFCL2inMYM6dkDQG1j5WbtZbw4jcIuM0t6x
1vlKsgPASVpWNwYiFBLUH/lbDtlibdr3GuuaUyMxk/7qBza8Mq6rqqDdcSQ1H6F6
4QnbgByH999aPkhDiM6B11vD2E10j4PZ/n3iwCy/Ct5qLMCP07q8YJWEfI4+ZbZg
RC1PaKhj/qLbHSu2gXATisoBjD1h3nlZU74faqEIIj6GfBYnln/4eV9gA0+Bpcv6
Jo/tu956FVUmbpUSU21sgqCg8lVWBmrMBMQ1qF8yPNXqUD0duCgLOET4c6Dbn1Rr
6Xk52Z6bpzBs6LESm2FBJ9zMX+LgDqSNs4PpQbbwi/zYjfyr2TqPBtryfbRCNb7p
HDtHuCek2ldJ0l+GZGR+sxpyc0F1ouChS9g2P+gvjyxJiEjtSq6KV7lY4y72vrC1
Z10f0JozEzYhVQn+Xh5/KrLUboq4rdxdVlEnE5+3y0nGnXFdu56kXpWJD9dB0b7F
fI8PuSdVO7nlKh+iXpAfNYDKT3h4EP6tivledOvgMFTkraPzZGlQC3I4clWccI75
6CiWswNavtL7zVtgrpWpXGgbF9FRW4LJuLhsmDn3q10OO/LdYe/HDnKS75ALSLB4
/uCU+ArdyeLE0cy2NFa6IswX5POFnk880zBr3CevxWVc7X4gWRYnRY3zHULgjP6A
GfE/kkHCvb1BINC7HpcOhMgTua7wvds2940XndFRihus00yS0qPi8y5loEM+/Bvk
4kL+Wb18GuCo9LAA8Ws7YIRm1TZpj3vEv3Pek+IQRnfBk4cgAZNsZtpOZbmckHpm
oZfDSBgWy3nHmSGWNtWsMwqgza8BHBelM6UMv+PdpYJNJLkidEdsAJFfNNmdGdUJ
nktJGBw03gMnPTdz/A7l0lGoL9wMIjxt86ZPn/7Cr+bGSn5aHkmCaMnV8xxuNsnj
F2eq7hCYJl6K8ntKkeXx9eEcL71+FqhACtNIGq8bUzKOhd8EpLmzBftwy1DwSfuG
GBP9jdljpNC7vLLQmWUjLQ4EPPDyeUp3OjSEs7cX6m4NpwEyKPPUsI6sAay3YhXe
86jwd+EfnIvRPhqvZTeYadOJecLvBd69xXiAbOKa86Au2fmFKKZDAXyG7fdMDVgt
gd9FX3s80EPqtXLhJJYVPb+tCY5B28bfdjhwUu90myOrzyFfp73MsJpjariGcHis
4gQZHHZZ68/7PA7kcz3BVWukd3j9WWzoujb+kBvex7NcMniyKzZ5JAs3AO8Dxjes
ZLm6pXQYwDYhGgIXLJWSVBETl3/FrZhH6SggMgLre3/uE7EaAjFRod5HUfb0Atk4
b0TL3cP7HkDxiLAJoFxBj0s61F6YCAczBWUZikTQlVjIP2ceHTfiJJ688YCURXV3
ZdJpnRz62BJGx/JcUuA/0YQudu0EEofZS9uF0pQl6i1icSYbYnHsJhR0ERI/dhDf
J+0tNUGT0pNIZG6hy44RttP8RliTJj4yo6qwDTN9VIKtFDGmTKs7Tbl+T5he5M7C
BaYgZT2JWpn9nAFV6JOcusdxc29qHnbXo/rFn6TrgXZNHNbczdhj77iAojWlc45O
pzk+ZoJvfuW8HbphPa1PttOgn8JCyBYKteBWP0+ovS6SA3kMuiky6KnQO2stmBM5
2Oh6Z7V8FW9Vre7sZ8pkUQr979KotPoPohK8ADXO0hyezfNu8E4NQdULckneKs+a
jcm4fTw3mxxdRB8TsyhBuFkz/Dd4iNC3VzprcA+KVlj8kEylzGRQRI8EOnEy/UiL
dfNhSigTsRd4KWEfLivo2oYRsvc1WCb/F3OK5bLCUb8sQ5cnuUbeQWyBWNEl1HCK
VsJNqsEtBeBFsGybQfHx4FJcbKcw1uzV6pIEnXHhXIIi94vp8hI/nlzubBG4KHSn
fVYV5kNWalGsk8CSfC7Y8CQm4R4e2Bn7xUtR6vR7aCz6ZJpdz+E4wIou5vW0nmzo
WigHYCpMv8qxgBMtvuykbgwhLCIV5dpR1wACvgVNUHzjDsmfL2aQnB+cjgkXj2Ui
L/8OcJg8pBQpjVUvwO5u1oHwOepyuY08DWq+XMFhQuAgTwEJozCbvuiPrOWw5WHG
9ULsrn4wQvrZmWWYlGTn6uP0nLKsqlnxNuAg6YvfvUl3s1HrolmDW1PrD5rS9Kfc
VsRhs70ITzv0bH2cAgbRMsEYzHuI6Owo3/oboVCG0wEhAIfCdgcO5Mhgkz3GOvlP
kj1LkWT8Og86yiQec00r0BLofsSllmEhHlLZ3bCSnT/KqpCcv4pAVcSffQG0Krgn
2xq7Eia9bbxVtXvsfTcrruL5hZYwlo3O9PBQlN6DtnXoZZqgiVcoXKaOt2EBnxHG
Z35681fD/1SBfA0ts8xvzAseBfnu06k3e9DodAf02rBHrdpjugPvBP8/anUhLsZH
5Ei9cSr0d4d49wRDQczS2Pl080UvM44JnI7OIDRpesq2QaNwtS6dyJ1sKVx0/1z9
/MY/DE6+zHcz6zemWH9Xv04O+/tLgarTeyUvQ3DA3eREG3pJ7wmp8eT8hWwkLQnr
NpDoeqclwqHN1o+Zysx2Iq9d93G2LbccehyTOZbEnUW+uVlNMM5Ya7wdLrju/hMN
pd0f2V5DGF8EvnWivsEtwa2B3m6LxQBC5ljA1VfNUobpRrcROi7GpSpvsyefTVUn
e3/xm1MbP9Ix6KirTpgoW6AngjlHtGW2UC12JA78Y8JFOnHgzgzLhfO2fwjOZPfy
OmNU4D1QJQj1T8JoQBd5EzTIi5g4+Jhjf9/dgsgNVr68e3PKlyP+IkLa/e1j/4Cw
BMf2192nHcIZgTLzXSYgyKphiId5g1Qs8owLStqlevPdIcLGflaVu2cVaoecUqKx
SO6Q05zHzCTiIOeg9cLA7O9MMbpJ4BejjBXuPhJ3Bd/kkWuxNb/z8lGQFucOptez
rOLhESvWdbb2ngfyTt/cYNS+KMd8w4jwfKRhJCMGyvo/KNriiaBEZc2o4a3/s6yb
+zMOp9rHNS74IMwl27bjSeJFPAb759ej+trDoLMXnyJq6nIfZ8xmMWube57YWtnI
8EuSW4SfjVUjChxYTkOybvmnpqqy7wtQiJPqthegxqz34EpOUJqm4qAmJcTRnZdB
gyn95PAjGmmSGpJ5gubQc0YlDt3ol+C4qcjNi18L/m68JY82UeZVamDFI3PHGMR3
WlMfdJGr48wKAVbbRUp4aW/x5JcHrAqwKW6PVRuqa6GfAMRUR+NEKCQ76U1BiMSW
+RG5miknVF3Pp/dGcDbL+NROHqgayQ9HwO5TAOKLHJcGQkaBBSIoETJpr3rN/1iw
BAXzHeu02E3gehlx54XOog==
`protect END_PROTECTED
