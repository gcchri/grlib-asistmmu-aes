`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fG270yOXksA1yeNwyMyW82sC6oPOq8G3dilooBSB/vQdVbLHEhwK6kJ/dyYHuv5m
sforZdpSffY2O12ki+UOgL0U7jIDrAJ1L23G1RvaNyE36+qMP73jNiPR74QRL5bV
ZgsYt52Rd/n0Ol0TRJw9ElJPFfhL8FSVOXKT+CsKAaBO41GaVCdbOds6edY2+ahA
yHidKC4D79DkkvD4Jiweks7iYwK27JAy1H3LxG0XeZFaEHrZbKRl0HFmMsIcV/5r
ALRZkZ1b3lON0f0G9z0SPYvLnLDjTUh6lhjQPUOtrtglfqRYu/HxPXoR31YBzfgN
xEXQT/3sAC4iFyyj/Z1/faeVcj1r8aqJZZGLp4N17OqbbsTkheqGAqgLgQkNldfg
+3/y1uInh+s1l1VkRVUWZtEMP27Qfkgp/yOoEzRviCjN4dYQRxknnlWo25tgYDGR
zn7VdoK+eLFd161P3Rfnos8ztmRQ1gdw/htaEvh9/QKeyiU8D5M1fh+KTG/mB6zl
OyL+1RBp0B0jv5b5eSzCRyNq1PywMUjJRvO4Kjh6UAO0HL0tpg6G/Mai3lRHnngQ
6P0ITjCg/1CjtkIjtdIce1bct7CRW+dUquz7A9iGnuqv5v32nUYirIcyugSMRC5q
qoGHNlzxqEUm2C8891Wt8qCWt0dIO0W/eBiUfv2Hmdp8ycpKOFBdmQXNlTMA+ili
uhRMAPa3OSPkP+iCwlnAB91lSXzwNPkmzUMJ8yJpfeRZUhQOyvk6vgI5943EichR
pRXxe5CKBng6t/di6Ev1fiEJNTeSFlnqER8BJcfO+24lGzHUT+DmFzOR14TJ0y+a
oQtp5A9kPACkPTXpSJ+4whxxTzYqRBRrAQCRq4/XvGv3LfR2spOnxAyeWzbcKekJ
WvjqRUU0oISphq3cyAjgzElx1lII4ilGQOrIvQz327yKEMsEX9drUk3CbE8Akwq8
jw18joqZvaHxTywx5wg5u4wwI3DtZvNp9XExM4qfg8R/4ya02cOQtyrv7pHcVP5F
Tbe8Cej/j3K9ZMLANR7shj/lOIRU1HugPkeWMjXleaLU8UJ2+ToegUGLkbVwxEvr
xCaekxsSrk/31h2t1TGfMPJeoIlmzK0HKaWtJhiX213yM1jMl5GDIq/Hmkbq+8z4
x9nSb8QfZiP0eWo18zI5wjN+GmrKNvGonsfFfaQnqYZ8FmoFM1IwALo5OWBar2Qy
z8q5AHnD67CaNlthYYJkOHefdAJ9tJavuwU9zxfBV0r7NZPM6Frv4V3Hm98WtrsC
fiPxA7dUt4nYPn+mR96ZsllEsHjorNVHxDXUG6kD4rtu4H03BYcEHvHyMTovngE1
YCA7fHUcKezseRRNUU+2pvjEyeQh+mRydrxep1Zh7pPL+RM6q07MOuLSV64TZbIT
FjvhqUoYKeQH4qt/0WzRug7Yaq0Wql1wYz1b3M0BmfTdz3xlX1mvyFAgbbrIZviZ
oKqbPWgWmwJVe5OnPPdpjK/epiap1dgzrmZz+oeDLKqXAKfSSyzABiKZkMeR8/KV
+6qEhChtYG0Wi2VMG5j6PNskKmKtig446dKlACqvnT2reS3LZS5v5RdNVC026hS9
a4xIGpLxjiVnys+8HuE4Je2YNNIoJXIwIPXZLUxthx5Hu7gXO3rNQKFcX41oj/oc
ppobnP9DL0UvVdy/IKA5Fajj0BYBc0JBwoGZU6R+Cjp7zJGHgIjs9cXNaTSA09h7
CCGhVNix0LGGPfv9PEFgcyFIAOfxeduLCkX5y/epAmeNfRU1bTn1K/Pzs4iOV1dr
qjQmY6X+aWxezzqE61uag59II33MeyrRsb9Zi2aXvbbGH7kaRegLC7tB0p2NfXxO
YfoLdRHMvVKnGnjX2tFW8jaPzVVFTnCbtFztj4D++i5xcl7m1TFMl8AKLLF2HdGx
LiRv9iNmsG1ZjOkHCYfxew==
`protect END_PROTECTED
