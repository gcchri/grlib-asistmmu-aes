`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
daKj/1KLtDj2gKY02IGhybQ1+FvsPdnM7/9VIzasnEyCH/6xhbvFjSYaWf4X3JzH
Rcx31MhgLsU4VAgnaQnS5RAchWIkL4uVvL/c15g1SFdgpwwkyi3OdtfB7xV3gyt2
QKDxYjGdyLYSqbU9qZ8IPbnBRqkLhKym9xoEwcQPVoy+6D9X/ZqN5+BOGBDPmeoV
RBS7yxtFFss5sbWtS6qJBKsj99vOhKECk+EUN8n7FSIWnYD08rEbSQW3Pd5WzABV
QEoOmw0Pq3CSnZgvrh2tFWoxZOLb5RiFR7QmVlG7r/9e8ptv3pzrxES6mpu36dvS
2mxffSzsSbM5mCjkvZWgHWolahGeVK0h3zzM6lEebxujRD44JOh3emhG4WwbKsfi
y06NTV5gC7DjE/9yBRnQ25VNFE1igl5HGgLrCH++pBwhG2ca3yepYHbFvAbscwbz
XtP0EVYWfXIpbXfZxe5ECyLCi0/hXwaWjbH8jFlvbTCa6a1Y0hodwmZTQdA7owOQ
`protect END_PROTECTED
