`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kIB53HHFjd3D0n08iAGwKEgf7AgTzdBg55sf0DI8p2aZtqkWh6xUiz/zOq5WISDS
+AUvi7kbxq4N5lZZs5eBJmS5fSRhwHhXq/xQRG2u1vzUVGQn9BdWFp27lHDDmQcD
ywgfDIX1qUpqntDi2NX9WffPXsGglrK0/0ltPAUNSwN4NInRbS/JjRVX/XpX2/wu
w11mvaCqk+NuKwsRK65/M5uixQCn5+wz3MitSxrJ/k/1XeWK3H7VLR4V0Ojt237m
ZA0EJevFxx/m+2QO6M+mUWSCiK38Qhzp2eDkD87sa5LwG5KZUdyDtEGwhoDrfJ0Z
ykyFzvjc3ey3o9LqyCqNR4P9kPso0WY7STz5KyyIve17Eul4FdriyZonMk4nKl6R
iLnR9POCXWdPwxkriC+0FAxzBV9kzLqG2PP0gv13v1H6nTZyH91DZTfoXFJYnWte
`protect END_PROTECTED
