`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jiZGXZQRq+bCgvYkfU8Dv89PcxR0rO3dw03iVSknmX6yqpPQGNdxMgLU0b1ieWBH
svNrSSY197uIJU3MgbNYgP8FGzwFJ6N1oXOBbH0V3rh8DdJri+3WwDw4/nzulpNM
HU1smJsk9XG1FiuYu/Sjd8+GGqmesoXeFUCiijVqYRu05ZSbbrutuJq3JVytO9+5
ipTwUAN0co/FWjw7RAS5BthaWLRJ8ItT47cPdVJTS7xKcsHEO26ZHZpEFNTRKm/n
334Gj9cYiET7Ye3zcb1wxfCmolVC8dnXtUssqSj8F+CpZm1pE+wNImuuOhltEeJH
zb8SoyFbed/Ix7pgqoISdC2RUtetcW4nC7pVqcW8pWFB+wU+wYSThX2gSM8xKSvn
O8KnkQ0OlmpBojUXOXO3OvtBJdfiJyhC5/x2OUHIlJpeRro8XLJMF1OG0CPY4qdT
`protect END_PROTECTED
