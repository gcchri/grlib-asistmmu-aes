`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dCIm7PzehAUW9niLyxBuHKzaqsWwPIOwiNL+58pFjAlehMauz1l1G2K7VtwRciWO
rjd1XIAF+uD4o27f0ygiEx71qbrUOdf/ntxIIkajpScXLY8kn77j7t90iunvrWr/
78IseJ6cyQQjaKNdX0nQdNH64xnAvOJorAtf1VW5oj9yGv/8b/2QYx6VdVErwkMf
uS/m8XfHHqR4M/g8GQ6iOGZtZPzd0CAyMc9Oct3ZpWZtvqTe0KS3qdWtMf5KzZUi
`protect END_PROTECTED
