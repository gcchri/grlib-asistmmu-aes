`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LpkqwkcooPYD1QLCb8t6AzlIFQyKeeJSHmSrYAOFkXBc2DNtXk5lTMz2PnTFzhU6
8gNtukvQ05qZKXsU9zywj5WoWJHPQpyfdUJ+mr4bHkI73ENZwaDrkarMFNkTD8RX
gs8uT9vZCnK1RoGYj5RO4PD+5fZDRLZzov5WktwZ2hlNeIpZYZGalFRQvysvBjDi
9mL0UADKjMp9UFtvG4UI9oom7EofMeW0oxaqwIHppOiCz+TcObsZm8E3EC+XYfoJ
l+HTHDP1sj+aUsycSlu+tjJ+rrOqgE1jK6u/G9mS5j96jSVUfsmEjX0EH8C05lZr
0g4yCe97Y4v2CO9s+UUz3wsevXfOKuzJa2vZ5jxdMcdujpgFOVDILggMgBHZVHYr
WGD3+G+B9NcSBgqy2MZfDYcm26ilTL3lFtEwFGzkBY+NEY+Hz3QDXUQsCfby8D6h
lMiG8kZ07f3yt/H0fyfB+ZD3RaFHSAojnPzIAwQw6DeEOLMA0dW+oR7Qkxf/KG5x
pbFz7N445uSpdQw/HH9j9L+qTTPkmxo0HjzwbWYCgPopVdpubJc55pB5mMw2R6XC
y6j1xa4adpTv5x5V+zzOeVV+IhV+t+YmYD6gnOKn6OD13+YDMtnaCE3mixHKX3t+
8J7IUo0c1p8t7FXGqHZhbo/WkG6SJ+Jxm5lJRe6FcFQXuh4P82U9Qfs62PFRht7J
K/VCN3fefxHeWcNivGYLilYpDjsxZVRDXSe1eqhfxK0fFldTRXV54pjxG6/vX1bv
r4BX2JrtJz8f7/YtJzXCSxW/lJ65CpgY7pgZPw2R/w8xirTK/7rJg9nGo6bMwzgF
jDdjblBqb76T8FfQDnmlYKRiKiBkHI3XArP6+7LelDoOiwBFyGeYUE5kAYqnMDcp
fN7m4uk+tD7zCBtYKOOlw5H0i/gEl/B1R4yDYLChABedaOIOqijSjzteQ2f1cBB+
c4TY+Ihc0u4S8GMX8IN5R0EyQw5LI/QZfbECVw2xgITUMwNNfBC/+sShh31dFkeA
P4VmIKwF57ORYYIG0VByQPa0Kl9TJOL6ErZ5pJLMCdS0PkUjl7zcoCj78YOgo4+q
+nE5bSAgTBGofV72vAYskg6GNvcS5SED45wP8h7KB0fTdlH2fZ6+CYSYzRBhUuzQ
HJdiWbGRWka36pxxjBldtTXegyW+/BwfCrVctifEZx3WfGJqYSXQswMkJz5aSQtJ
egDplW6gkkmZAtB70KwtNG427dFgCI1tPJ2kopIJ0jqhR+SlPQeHhgPJnFPxsbD6
J5Fp6ZqNsWPlWREdVquXpZSG0Ud9QV47C6QXuvOTwMFvLebB6wIW51JlRW0YrIMv
Xk4yYPpHJa1Qv/cqrEfc9w7FOkXC9O12frZgtFbER/LlV9OmFbc6X3QEtE3kGFBM
Z3GTuOoSICn2uuAVo0VZR56hGd3gCUEkmjQIxKWEZA0T1QD6BnSEjTu36iiegkoM
spo0IGhWHkkKKtSNTaWJf/atM1IxH976OKJ5f+rLpyS9W2lsB4F/GCJYM1mXyBf/
Jm7qyBclcb9n0mz2p/Eo3P4oPqjQgmwknwfTFmupCYwyIiUjff8GwiP5mJU4A74A
9HugNUskTO62ssHjKqLrCTwH7EbrkxiEC37Hm5u7biy5bL534BzhBjuH7nTQQ/UN
GegPK+ZvfGsM+GXR7M3WfXTqCTaBFJFQ6/JxVdi/4R9DkVM2rPrxoeQXPKgxJfdJ
lqCNq8XzEwGgKzmNqeEkV30F2LAEWMj0sE+ngeHq95G2cF5YzFLxp6pkmnNSkjnt
/6EPWWe1GT0A35Cz/w+zhDIudThO2RCCga8Nw0qMGrrSZIvvcfQ9FQ1FYAEexvgk
x6H3er5PaChL/w4efmwDuOmKtHhwb9pwxXf16VHpMSwQLwz/dp1ltXKnDmNd0nnE
BnltmX7mo/UxRqDiOwDBRxwJy3cB80bRiQriPh4/bEzOmQSY8lZX7N9Kr4CTTUmx
XDNDFGa8m5p4bA6lylhaIpmjTDDJn8eLwgn7PHS3LiQ7VrwdZvJYyI81NL6Kaigo
18QCRMOtEM1ssJsmiNkfcGxE/M6Yh9A+kcQGWHEzgK4=
`protect END_PROTECTED
