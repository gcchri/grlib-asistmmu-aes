`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qbw9S/ktP894S+4TxwVV6HAftvHnpJzrXonQWrcKG1T4cQA7ymAZsUfXRR/iG/Gj
adi535mWHJUETK+7x5frMWy1FFgHFT3lM7k09l8kcArBrRgjA3c7li5SQQcolTuH
X8iPiapKfw7eAhd+qfLUbfhDy9CQy25PxttMniG6t88ChkNvK0CeIFUq/Lxavdlo
CFwd32vW4oc/kpcHLXXYaNeBgEHs01mCm60Dee+J2ybG24T4qwsXxBieLBob/AwL
mzkT+De0iStZJ5T45xh11YWpLPDMRbGiME3GI2OJV6rwLJAxLvo87AcUQe0lKcVO
RGDxAjSCp8iXcd1yqWtcG4IwqD6MuroqnixbApUd6A7ZUN+y83Fk+jf1iJMBv5YJ
waWK75oPwbNcCZ7f4olH1+kR8UF87TRDh1v5HvgQww62nGLySzH0KI9gU5MEygVZ
`protect END_PROTECTED
