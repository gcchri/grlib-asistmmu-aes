`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5qv5nBmG9wMbUkfDt08zqMVEBSFm91nuZdDuf+F1bFRvGyzgB3KygqZOu4rXygQi
DS/w0xAh8EEWUWLDg/TsCQ9CjPCZH0HbKB+uwnQyaTmSsI9uFM1WvmMh9e63yRz3
zxa/EC7Ism5m6O51qcAnDQWQ35VJrkYGa2MWQVduXoiBwxGwQbH9FOar75FRIMeq
NJnk/xjCPzyFPxhUfI1+IGJ/dHd3zYrX0hSV9ZPlJRhUOuR55jayKxwsuhKooKXi
iUEWMppm2XZ3xMR1gWtB5xk7kjEfCSIsZpJtT6H7zzyd+iG0yINqw5xuijckUMqg
DHePaEDcYAl6mVhBf02T4OgM8cpxTBZ19ZWs2Em5SOqo8IEolvbr52gMOkHV8nxS
6CDOpPnbG+hTfLPv5pzlG87fd0HMOux4taLe7PwDVWpSn5uPMEif6IgDWp7Hp0wH
`protect END_PROTECTED
