`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vx7WUDOcmYWfAanpyjVowtVZhVwrZfokzrhGNCLY4NXWCTy2O6STPG2JPDRb6/BD
LsQ48oOpqncH2U2mhXf8xdgCT/Qge6QdFpSBHV4ylF8RLSThSG7YXDfmaOoCKKK5
5pW99FmGhSq5FXSoFdgw4vC/uM2YI7Oulm4B7dLfbH/jJKD8NbLamwT83oqDXmxU
XqshVudykMh5j1mdC/08IcUN0yE4WK9PQ9Mf6x3GuBNrMw9pJ9R8MR2ZPL0k4ftj
ZirqpssDJnccmdaV0vFcHkof0fXG495ydUShyy5a+Sn/Ko/rG4TGWACDmEFnd9vK
lvH5n3s/tw2kopP7RDjOLA==
`protect END_PROTECTED
