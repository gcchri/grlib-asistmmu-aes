`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IcAdLRca4F/xDeYFMIFGAyvPs03GtwapUZY+xZG1YoXaWTzoN8hDO3iN+XBah59l
nCwBNceJ5BpBCJNiw9KY2OWXY2yWjLofaEltqLTR1en9GJ/SE5deyUbo0eeuNjLP
bdNl9g+NGTV26yv8zuklhDRWHTzo8vkd7lOfl4RBOzR3bIwvZwLU23ni0gMDnAbv
aXqgidVYHr0NsIZ7eXq3+nSKPgzJeDq5BU23OmYAs+T5k/xJhV51/gQqJV0wWwxp
50Qhgu9NOqsrqcG0JmuyV/pRUbT5aAdF4Mf6kegOGrkxRoX3CZ1qTg8OWNypXeTX
YXxfI0GRHpJD4wXoF9+ScKd6b+0e6yRwO8HsH0Ykhf4qzfM4iy3rHL9hhOi9+EBZ
ixJCPwd0oVV+75PKuXsvsqWfcVBXvPU4aRPr09gkhWCKOkfIOP2FCMaX/cUwySpd
tMp1zC9Jv2waylsDzhddnTbrQ0rnfeybabQ+IkJwZ2cOmlriAc1thps1bss/4bIn
f8a+Ph51pu5J3nyLP7YhUayfgjovxBNxAHY+xBOUYYgmw/zXjFazIbHHgi+jJn1F
tCoF6XFvf4Ip8e+Ls5GWZ1kj5gk3gUY0aSQVp4pQwKtMq+3ZJZKYqvQOcvaberVc
vA17Fn3fZ/9JMfu3kYHtxmkcu2QPqQsZiTEOvG9P7Z1Cil0vzarcGBbxjM6HpQXQ
HRgK4keXyDCH2xKSEvXsPTmGl7BK5wM8ctjkgzUNFRD6CAn4HFWMOgwRW7vz395C
ckvM/cHsI+IgLhbxMiU3hIZktXIGNDH+McFDaIqSixmGglS9oJPIvBoaXlz5qKfx
5wJx+i6F94jUyOofdg7VvjuH89sSfVxzSbIyhbm2IgvZ6jp9Y849CgOoQRQPpqCv
Bex7XFnqrKf9eCXLX4pM+w==
`protect END_PROTECTED
