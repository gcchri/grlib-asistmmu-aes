`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7E4j4Ai4QBPaU26t5tVlVvF12IqIag8bTHMVuaRkjy5DW+ivvrzTNt3bvyATRPXy
ah3hEMrED+68qWCXQJl+ZFXeY6igliASQ5W4i+WCc7d/A3fD5/KLwcqaXLytTQOq
Zd66zw3Vzk9R0IeKTcuca2X/gWEBoBXkkg0TttuvsAiv7VYbCRX0Jh8XRnJxAuGN
VkbseywlWnigJ88vIWISzVVGwK8YAxAY1OBhwWKUKvZ+bV+n15ALY4gK3WwJa6Mm
WLzevZ91ZTNNhNBRKcfWTyjq+tY3Pz1qRgd7HpNO85C4uJ7NR+vY/W7NE8aWT2La
`protect END_PROTECTED
