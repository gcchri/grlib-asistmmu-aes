`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JnEk+SUc0Q42gDidlSETjicOwGoiRp3R3xQmZhbYP7LSy+dwY+0psGE/pbf3dcp4
Z/BU/GSc7eb7GToKZH0dJIwmH5YdgGpK5X6ENLwdgWglLS83YiGfwZ/B4L2BbTGg
5kDZjm0V6LCPPZYGVxUA4WCvO/oSP2woLPklDIsgOYprQVaPtmcoGx62tRi1EwEf
RfWnQtPuh3Y+GgycZxsdHcOE1c5Jjgzoe9xgblyMMN8gwUw/+F+dT0c93iONvYzX
vgl3xH4zzui2GDl12eXT8YPHDQtgPI9/neZCaUl9C/CwOiwPhZf8F1GGIyg7OWko
Rwg0PUAwwe5HWk4Cu3B6cQ==
`protect END_PROTECTED
