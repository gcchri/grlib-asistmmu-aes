`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Vh2eEBFrS/iTwgZbu6vlo29QLxtLFPfMqHq5m461JYQdAwBxouIzHc9S6cbcN5L
fXHSk5wLrx61QeVrC0Say6ph4cM8D47TxO0589GZyufGXQJS032qgv8DAuczDsAc
nsOULFDut3SabW/1RDrwdHvmPYhAN/xbgrRzW+PreGpL0F3s96gwCnHT2oyLpI/g
8CqIyTHolYypqCD7SDBI/RytHkV8NAl4YsQi9/cdfTCgQAElZDgNlD5qD14J6D9b
kQ5rhmGNdE//M2/4kmI7Naq6bihBQiynZ0e6zhkbQFN9v//BB8w4uq9rNvJr5dpb
kXgcCMhT8zuAMMapplwEtdP8zTz0q3sxJ2IXU318T89y2T34F3xAeMvd6UknmsGV
FSxNPeZZgkygXL5nFTRjHpUdBdmXd8A+7+bGLiOgJ9N4mJbkli6E1CWJwEtKXeO2
BnZqVkLgCuYpHds4I+mqKGwQcijdp3BbkxW8q2bz4Hx7KuZB6HM5INbR5ZwE1mvq
eEE7nsDcDVMpxk4Mf9KkvTP5PDp65oJP2Qk6BFAb+759uWWNp1mEGKpk3W7WAFM3
jhZBH6eMQ8CiJ2khD3hxhYLi/lHmD82RpPCYHKqOhYA7Xpgwh9ZFN/hVDK+891oz
dGRqjBZkjIkaiPUW9KiIGZFwVZXBAuEZK62qkjl2Ws72LA86QSDSpQhbaZ46u/1M
86SgV2La9h1i9roNrz1rnTXpUDLNzPgsw0ErCRub1bKBYzRiT5PDIynUyFHxh4N/
JFacxJJ2r32AgeiBrt5q9Z0SRkI9UvWhF7XQCo5nYR6fZ7KC21wIN4XPMST5EMRw
rgOBisimsSIbXaIhKAxJQV2i35sMNNDED4N7fMMNqm8Zfqd8rlpF5GYXi42rQwkW
//daYZtsovWEY6yEU1JWUvMty6qPmzKIAdKWMkMuMgBhDzZ+gItESdXFq97DEH0Y
RsiuyQWndsEqRJjl/JlOaE5Emr8bxdDQMk/41AvZvM3DBiaPIvmBgXjV4RQPOuna
6mOaVNt5iDfr3xFbu+5BbD1aoVLqkVFUPv1xyeTJw7uDQoxqzWCc/o5lE8z8ck2e
MnytqOesGMw+Ic28JXep1xUpFgPhhZiS0Aa0hgFewGdHGHnqKKtegfjT4v5ID+3l
aGKaUnU6B7CD5gou8wON9GMG/MH6yPyN9Sm70L4UTK01rGQniqTaw+yLIEFSkNwp
3l3mMIBHp2twzoHyJzVzuxO3ruNorB7OwoAHTAF0NJOk29v5xz6CRtcRlD6BuaK9
H2wchvzik0N/0obSmP9FafdxaK5JhJIqEgwKclOTrAcoKLdvrekh/xiD0F+MW1CY
dEYrFx+Dvs4uO3jqGl8bDpsNLXnmghRDBSR1XPnInU2wd8im1E1pOOmoSHtdgPbE
P9fMeD0/9MmCeUWhS0YCpvsqC4djWa9zsldYt+27yYA=
`protect END_PROTECTED
