`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tAbhD5hALec/BAP7LnpA3pNUXEeiw+zBK+PBtVGzqGqnlzU82KPeEWM81iewRj0U
56ENn8PK0H0foOdCRo6TvuHo0FfCARo/hNLV90b+fF/RbvZTis3ZjyYvdBgJCt6U
0zLli3c9tTFupBw5bWaSkuTCGjfqE1cRlLs27uWh3DiWcUJXT+R7g/O/LoZITLF2
kxTCfbbBpp/yoZSkBYUKJ/TJLVH61S8qACFZRo4I0dRkuZPYfgTs2gY2VGFBJOJC
yliOYXJ4leaSSxjDE+3Uc9ZGsFMWjjXitTBf+Z7FbD0=
`protect END_PROTECTED
