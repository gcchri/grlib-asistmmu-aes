`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iNNXEL02Gk1mR48dmcg0CNzwmN0F/2yOsdcXTPQIA3eL5HELTDhoV4WFStLydh88
o1Jj3CLdwJqzYJebK/03LooLs8TjBNllpFFrECLTsIW0e6CaOqfmQRR4eq1GE0TC
fdxhbnTDnbYXA+5KogSEww0SOwIcKvnXnGVhRyv3OYJbQIwq2/pFSslggLLT1/qW
KwRZojNce0nQwbuKb8lcD/pjUzotAhlKvdauB7DlQKnI4/FrX0AkhVy7zHmD1n/i
ufU9VBynebguXkGAE7PIuu7rdsJMGnrNlk/uDa7dEAI9ar3bJ41d3ara9sJDN4ip
FIXcmrIvTaIbspxoaNYTZH4hs8ryISDgtmTg61m9IHbnr2f9LldzT4d/l4w4Z/SN
p5xruXMqQY9BGUO/MMXu9KejppCd7KHq9U8rS/cQop/ANVSerx++OTpF7mRD0dpp
s8VlD4QRifkUYtYfEPLnDaqwqPyZlfsiYvIgf/zD6EBX4Tl3yNSrBbLyWGP8bt95
9EltvC4npT/r5tZEf01mD3UJ2j/wqJe/f+QORMZgSzkelb28WDGPw8qJAPMkU9vx
UpEjCKyj9FCqUWp3kDV7iz9zvIVMwx438j81+1CuxhvpUafrxzdJcfmNDmMdVP3k
PrnUO+rkUctk7eCE/m+mLWf1trFGDQHcGX/X3svKqd4kmwtWuZ2GBIui39RQk9bh
6Wp+zPjCt3/y/3QKV9rQzE6WsNvJS22owsATomPPMfd+xpeqxLpc4r6+/4oDgT0t
vUB89+aGZ56vpKpgpw/RpFAuzkYrk2WynEERK5ZwS5NfFAyFJP/5KQ7zuARhKei6
Ig7mjrIuHqrOnUeBjBa3yG0xTFWK+ThXEp7ipIl5V47v/zzlWelCvkfXkw3XE3ce
Evxq/NnSJy7obXJEph19KOAR7QsUPX3K8kIlIOegNWrNgFSb67xrcvCmFelKiCEj
iAJy+YeyywQbYjZJ6NAxE+sqJhtEJegdxQUx/QkfDOtuPY/ZDtEpdDNUnBdxn0QR
0dkXKRC5t2BvgXon1s9vLSdzweTkcbE6xZs9uPcj9zgVCj+oVML1/EWZTJpfCFbi
rh3jo5XY84zAl1C3pN8M+qsio5vmz6EuTNPlJTsgoj+526BLY7gSpwYolCf7qhTE
kJEH1yAXMxbO2q5oNC0nQuP+iAD164nghz3w2aTAYrYNl00h5wBHYtHOjP3xk5+e
5Z57FP+NJGhKHd/r5q1eROaRpwkOC/oKZDGDP+xNJVtB+BGhwuyj/JjwwsAEVCHz
n1OGq2gOgq7j4tBzMWbJoU80wFDKvw1wTHil7dhLrhNZk+vMz3vldNuqT8FcSno5
3fc/RYgoGBkR/StP0HuXGhcblYyR9P0vuaCy89f1XJ0hbzFdFFrlUg1JY2OS1yW5
JS6mLY0SgutWrohF7zXP0ccWCBwfYT6WaM42gLoKjRNUAE4x+UU0qcxLa7hENgbD
JPMlIQHWBYojMf7oiRDgca7BKYTptkhDpCip2FKNsySQAb/NZDGA/MPvcWYs6/SZ
GS7TN+9sk2d3lgtVE7FJDVoA/D7BiodZ7Bo2Vp43vOSdbRT/YaUhXn/3A7H7FoET
fYNTBWMhKBP2HwVm7z6vyIhl5HcBa8WjHQGlT6NovX1LInYqBnyJtUu9UbT0Ty4j
7EbtEzGPt4sxYmpaJIT3GMtdQVlU9qgqlYzvl9kjoJ3KoGHpJ3OEnDKYLJEHPafC
IbThF+I41rOFdzvreboy2gbAycUCtwGg1K3h3QZDpq5nZ9EViilQLs52rx2nVwr6
7Bh1LHTnJv5EKzJDLHNYmC1YrG/Z+CgbFqqPoMw2v2kR6IF9R2IkkEMKkZ84BkNC
paCuq/qxL+8mT2XtgI2h+0ouNjmyttaBZmaUL6FbrURvC66QwvUMit/2ddEERoD0
uEpDu+rzcEPLbnnG+A+p66d6Pxc98jwGTcfsKY+WJGHt2huhP3AnYf0LkEzo7qSK
0Veyp3dqN2OzgxaAPdtSBw==
`protect END_PROTECTED
