`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iDIcQ7lQbNp0N+m77rVcMLm5/UbaMf1Oj3gNqcHnYAeFFTcvKw8DPVlUvOQDb41D
8CeL2OzLjfVaUayPqRT1nmb2jP2eN4IH6znQNtriOn6CrgWQ7RrkXtei01m7IIQq
vezEiB1EdimBPCwNlmZZw7bWDYtMwX9oDR+QegW0kDaZDv0r9da2YczeTw7sNrNf
Dt4OfqKYhPbuGPyMNQsX6PpuRt6SmeRLNE8Iiqm95V5GGzq6y9p5ncRZTLGeto8U
v3LYZ5c3BH83VpHho7cUXb60ydOFwGiMRvPglHx3Fe3hqYN+Z3+3B3TNnF1xKuST
moW6WAjZY6h8ezNAZ8pra9nqXaukk9CRfj+oWYSS2OGIZCqaE+WXrDCg/9rzIHkq
fxlopTwireWhx5oi/wdjT8edaLUGMnqKpO2uGuUkpBwmypTE/L0qwNEyYG75+6Jo
FPZ3h4uuSzzj7hRnHuic3x4HhBKZLaZktpUGCeHX70h10QRjX1VCDTE9KsMVl+T5
QdjOGMSDxjiHZ5szBEveio3iENbxeDOMqwIwKwyP3npmOATbykPR1y3YUnTcayzP
oEMbzhTclpTekXAY0Lpbpg==
`protect END_PROTECTED
