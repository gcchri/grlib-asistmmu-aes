`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eAUZ5gJPZ4VzrWtOauGUmRlD1tZUL7UwJMEu+GE5UYS08Qfru2tbdnDGKooFlETf
9JEMTyz2Zn1WWACBH+AjHUHF+x0se+7zbB4wv0k/8zYoVzzMB27Ha+Oqb/pPhmJD
A35TmAEfKExb1rBcOLw02fcCJqEkDmq+W5nFuxr1VdR762djYPenS6Q+2O4XF6Ur
B+onvL/nADQERVDx0UttTdwQlsCt54TPTGLwqd8+X9h551UsobhG42416Xcs0nTq
UnXBgJYFv0E1NlqhOBVOuN8tPpi6trvaf4K4iYZ6yKxpYhxml3J/X8kQAC1BhL2x
Gwjuz9Byb4PW+URZNpyRaQ==
`protect END_PROTECTED
