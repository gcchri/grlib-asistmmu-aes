`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wPOjGNxAr2IIM5N8dJZu0ODP0LHB6l5tED87HKX5LimQwEtny3hBmQHjkO4uBtpF
RvJvOhuAh4G/Kn5+jMwQKcD3RF7EwLkC4AZ+2q7asLQyuqtcMSgWBiKp9Ob2QZgU
GRd3//QBsql4RweGi+Q3w7z08pDEcdvarkfUO/eKjp4fYlT+wb9iq0TWmfE2wHff
+1W9NXPdekUrl2nNOkkfHR1uc5B7y5xlXrXOcBTlI4yVZUjB4KEVidgd1m9oFCqV
XirPxrp3zLF5A7cBA2ofv4qoAqDNC9WBZpUKKMqH0UR7NuU/o2rf5vbzX+4NXmXe
vOlyN590NH6Xy63AiEuozdTDmbi17ZbFI5aToUOify4mvjaNP2b2jgPPtuuec8K5
x4y207OeWXQUXbEPQwksb1NBAcvAza+e2o5GLXu2sns5wbfcIN4jCU/ci+bjGNzb
ZnwHoBNvbiJpyiRkuIz4eYwFU4rI6/o/rk9NXKAQcZ8yHOaSQV0WnzA/ARLLV36A
ECfwRSu6ZMerqWHUBLg6WvUCq6Xsc+Gh9QZsOXKDxWwT8uxgS8CyDQ3V3sA+8zid
ubgWeyM1Fk11On5CkXdTVDMVOlMTaLZBF66Ecf6NpNyzn1C8JQp1ZShZwNBN1UkE
nlU8d11ZvdpNhMLoSBX1KFV6sY6iNhQT+6FHVa8FZkuX+s8LQFpRzIGf8lxlCGw8
AGBK8WwcPng/aErrqU3JlK1WLHrXnl051F7lDBDGtSAAl5q7yWYKQeJkt5CsrPcC
P3wlPosurYW7PwmXesUHJJ/zoGKKCcflejpAoBqFVfhINcc9U/3S7AcmPqATd7Pk
ykAwRvEaQNvpJTEgieCiB+JKhIGFfz1o2K4Jjgqj2y5mympEDbwx1/PgYBwvp7hi
E39BD1olVyOqhXxQal4RuViiCAiXQaT+qkJFXDwjjrvKnihsj3mjuQtHvRp/nD9W
`protect END_PROTECTED
