`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lfk/ecArvZhABFZ/IssrkQYhFa7rM50c3iY7MUxccdUPPXGG8+pAwB25RSLBX037
e4zk/y2uG5u9AwYtXdm9HBQORlJ9fhpgFBug3gqkGMZrSL4oQeSxK0RshKDmy231
llzKuYfy2IkjAo10kfDfmnqy4sAtVwcaQ+eJ7TbjVHIB32hmvSXB42zLlagb2oo6
BAclNCJzvyYOFafeIB4P7w/1usnOEsSNSWCez+p00uk8suvZZxLD69Eh2c95MF0G
PwwhIH+DgXgNZyd1lONpMLxsO1Dr1F96z/kM11Fpv/B4ehsHPyX8Ym6QnXwCShGg
CarCKT/vN33t5fHfiYvJZw==
`protect END_PROTECTED
