`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/LMWnPjyqtBOGZhT1NuboWMETb2z0HExJly4yimMPoaerfOA9KJAgJ4NmFghrlq8
McoLebc7vyRCFb2b2AXPLdxo17UkR+kIyT3wNCo3+3AREn+WJMGAzcLEnbuTGeub
Cbk+F3GmSxath3QKuszzE9hfUGwzrOpyjTHYaMZvt89ZJzATGm+xoZbgseJ56ys/
cqkkmb4YVtjAxuAdUXIn9GXBwCB1GafajMYsEpQgqzDTOWeRGhK0AaarnqS4ow/c
IcyUZ+S0IT3vlfB4DtHbK2afUNx6ZInlnimz2oEzdNXjR9XohWG+AypTnBvhv+CQ
t6we0MVEa1ZjX7zraQN8Ca8mK4Tz4Xh5+6PUzaI6YIKrw7KSG83ftbNLmE/Z7p0o
4OTudoIx2f9F02KNYBVTL9igZwzI5BN0w7yHX2/qo/48SbFkAftEAAkBVNupnhJF
ghq9NUVOQuNSsBpclksgBDWx8OPH303GVlt5Vr5R+j1oH9GxGssOm6e69Q0RkhMD
`protect END_PROTECTED
