`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x3I3w4ockOZ2u52LzM2IPk2jMKYTcmCNvmn5iyg5ugt6lG2xcLs60Uq7TU66B3qz
ISQMZR5uU5hBuTGwvZ76TjcZveBs6znDIG3q65jBaM058WDb3YMzsweIYTvoBcxL
FvVrMP9GVM+HL9XZoiE2xCOhmXUszeOzp0lH+f8S6o1b7fkcOiF20noMjdBgCqtE
MwYS1pN5EQnLzUCGcQ8wGC1jy29axU4E/szhCWlIKaxXmHMsfWdRlBkXCxBQ21JD
wt64k3OYkAZ7qUlFId5KJyEWIzb10Kg+y5klXAYWMTfQh1C4QEsoozFUwhYz6ENt
xPKOR4YjMcJnW4B8Zwa5OWo/IgMs3O9t793BMpHrY0sMdGpv4fKoSWZALKkfJtsD
xXPnqVsG/MSnnVcmVCpHmg==
`protect END_PROTECTED
