`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IUvI37QhaAtcKyTZTTUxunaCjjm+f1BZ6Of/7qHFOv/wQM3VMasDfXnBUMe6Lxra
5kjvOG/vayo+R9P45RBoFtuZ0cl5d1SJHEKrQ5NkMxsx4d8athV7uqC60q5TXh44
D++52YbZlg14RT66f+Ww/cF5zSvT51wKdfW2LyMgJ6zEG0nPdlFmJVhtiX+u0SAL
kMzOxpjxaVepLdnTn6OVtVGny0xMoOlpAM2ty+ut1612aTzYjgmqnisZNLWMrpaW
mu1U868w2V/9XR7TbDroN71Awcjh1/MsVL3jayponTGuSJP7gNfYEC8lS/BlAsMF
7e9YTW0zNWbkCZL7IoBHg6GAzj8l09xU55m/9dWFv1Uy6s5qyDI1auiYYY8p+/JE
YquDACAxiQJBGPG1QM44OEV3yrpKY70XHgPiv4RbZj929q8hMaYQ15FatBD1aV9K
`protect END_PROTECTED
