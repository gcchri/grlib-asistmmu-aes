`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YJ1qXDHRyyd/hFDiglcKWO26UAB8eJ/kNOMBkeT39xH4s8NqY/+49+5Q0uI7dREN
2mAHDc2R4tHn1MHUUnumVaW5UfMFv2BMTS39wAQqbxGYFHSmLzNYR+VlktqdppKU
S6Cip3B2sGqq0HxCf3pkCgfzP4oMJF9nA299OFY8LgPTZIR0u0ZYccBOLc4SNDBS
JINuHslF8Y3wapJjP3mXFhsus7WDLw8J8XOQASG7jzQM5FvGvStSXyXisdPqjtuY
o3YEeTerFyAo1inbh8L5kY2BMsGU1wK9o3lIVzIAcwh8JZ5laEuUDLdgWD4qrGSq
wUimwKzUfHr/grzcTEyiLw==
`protect END_PROTECTED
