`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JdGbbXoJCodk3RqqiQbfNXCPjclSW4S8vhhI4DUZMeejROhoPYPp9gkvBRuuLABt
GCL8hxDitblguXyE2+TSVdskok2BRZ3E0kLom/v9skBixSqBMTfBawzw002Yixnh
g1qgBQvHHBxdrPncwDMTa3y8oVgvKcLNefn4jsNAuuwDC2dGE5KZGlkEoLG8ZhzC
uqzLPDLEvUn+x2Yp+98tJmeJcvA6NAXNy6P4gytn9UVppmgN6yvluJ/tzkOrvO13
uk6TreH0AEttRpGaIFvX5zrJKrGvzZPt+XEUCNB3PM+k26i5RstVJwtei/SvdLQx
A/CwsWkFWGKYzU9oBoS9cA==
`protect END_PROTECTED
