`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FQ4seH4EYzbWWzbreLC8VJWgzia9vVvsS221xQY4hoTiIxZTE7QwBKnVSUWBE1/f
6YsXiRJ1JpM5rvFVzY0FCZ/8bRvJo5qq/I6Hu61SfifQL+HpRYB7Ic5tTigfFKGe
O2IVAYwmHsBhTum4ye01gtCt+/p1VC/BWBLiBUjxWBczO0Q112w4buvU+5fEOfpt
9rRZkyAbeUfUwk24P8sYkaLJqoWVk9enJ630xHGHpQDqhbYWLCBdtK+hhf+f2f88
Z0dSeSNm7gYcbKMbvSdBCYGp31NWJ8q0ahaVj5LG8Lc=
`protect END_PROTECTED
