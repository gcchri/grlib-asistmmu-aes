`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KoBdqShJNKkv313t5UboW0SNk4rUYM7Spw2fsZHjGR6LisyufFO2Y+SW/iRAsLZc
+mS+c2dK0/4e1cL1dJVlWsRSLMvLBpT3bXmAy8wjmBeC7/Fx35gG8OshW6akDcBt
+pTJBIlJqbCWJiLWgIER0FYcp6k76kPNdON01ADgMnA6Bd/hqPOb3Z5UORYHG7BH
IQeDPJNI0oE+yt2FD70YCmAzI7yBCznW8oVSmQK0q3Rlnyz2Fj3owHnv799GNqNn
L9iAWKkRW944+9ZKQvuoPUWB1Iy/LXL8w5dqQA3ISAB2g+1BCPRVuOG+DebRtoAj
4lPsQScxC8g7W+cTR/Dlx2lKS3qJTpl1fGB4kaKH8G78la6rx7V8wGbnA4WdU8JD
PiCnaxnVqxFUXHm8/xGcW+tTebMFxwlWy9G8hj2DxgKFW1OCFUGvODzRt/7eCxBg
5kcyQdWZevkXRR2Jcs3asf+o5iXtvMq37ptmdAeAc9EmLWv9mlLwHwQXIEEOSAMo
KcbusEuGwlycfKIT3UIGjFn7VMliZ1vBEsIemrKAhO3jIRAYB5gNoRHx8FU40lD5
AuPaptACsofE4gGtFFA9Y2QuYGQfJBrpibRgiVU56mC5CuTYl62sINT7k4lAS+Vu
ZXccoLG/hHgQmh9YRxGjfA==
`protect END_PROTECTED
