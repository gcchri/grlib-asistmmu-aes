`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W2LPQ2P91mSdQOqbUwxqvuKpQelXK+rd2U4itBEEzx/SnbXN903Faj0xHvsLChGS
tv3mA+OeZD3jDKNo1x8voo5cwBcBaYaMXVG2+ReOLTrQ8PnYcM/H9M5v47+znMVD
W+5fCROpLb3f/OZAnHdLJy58ot5rO7rv27AiIoUIobl6chGQGqseHUtEw3kNrFL9
mFsQQd3ToSvuaRQ56ygID2tOQfvFpruFSoJioorcAaCQFkl+DxBVtjraJunm2raw
pzVIm1Wvi4c7WhSbbJuqou6uivPjuVcFIjetMPGnASG0av9KXXpjRPO6LQI/x7XV
gx/D5Wi5szXNu8pk7UmkoGGJmdEFYZvS4adfgF/HiZO/D5WxzCuwn6MiNTkM+mQp
a6O6ehHCRmbMt0L2cIOslfvfeCAGMzcgishWuvGu5lHgIMu2aNbV7eVztt9YFBtc
YCbETnTo1GybKKzU31YqQtEEdLCyYb6CrUwyKzZOoKfjlpYn105KsXYYk9Ps/PAH
UwVY+YcA3zpsrJl0uMPCWxQ0WCHBnpjmpf00EpBA/CydPw5VBZF5RqoiZD0q+X4M
`protect END_PROTECTED
