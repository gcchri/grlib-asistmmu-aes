`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rgqgten/6zZWO+SL5scL4jwL7U9yxVvBIOWDGsOz5pdKi3gNRD82OMBrIdv1MBQf
+1ZfFXxmXLuq5SkdNP2EsiTGQsHu6Scz3iQNN18z1lJKOtVNXxywtMjwXkyUiFyO
iVl5D2VUM5wpqL1Md+/FJceo0RdANRB0xlnjO/WJSKYJWylEwzM8WBj4KCEjaV4m
RMvz3QdPO39i6koUdr3uTM2sgGPJAqt06HFT70ebEIlrWhjPnPmAtLjbkJqbs62w
gue8RrtlR/Q4wmPBtvjEDOUeEk3gIVbazPCNzi+OyKSpcSMQ3gGRBmMJ6u+OjDNO
`protect END_PROTECTED
