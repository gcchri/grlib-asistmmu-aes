`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+iOCFrbq7oazjvJUKTOqTlEKYdVrCE+IevMZ+a3eQSY/UAi/XJ/QlCH/GqgTOYU3
aju2eh6yGNCj6U/86LcaZK2eOUV8IU/gOIzTLB4nwV1uIiRjfUiuUu0dTLydf+qs
ARjMPa18XRUdlag8otJWyZEUdb3aLYCJ34B0DWKfP+wgbbja9TCU/Sd77gpTA9Dz
A8MT+UoIA101+5hN1KOTQGkXEFDjEf8mfMIWwbr2RZO04GFunMhamoRQXRtmV/1p
sPajnI/KJaGKj3dbcCwR28CW5+9SJYRgp5m4+sobnJUGfJR72fMbMLoCkPC+R1WL
n7YRA1Yri4dCW5QrUng5OPuT4+elejsU1JaTOMHzsPJWaSvFjpDTyd3bObl89V4T
xq7e+qz4svjWKOmaLY0EP39TsHBT34yAz1QVmWLDMv9pWoLbC/Ceq4jo0QVF+pZ0
`protect END_PROTECTED
