`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
youuZnhIvspu3cK0FumsTBbamCkLvib2uUeWTfY5o/M/7V7efIltQJL/xYIkmAQ/
wu86pZEEJPvWC9Qe/LZoyWkhcURkEBnb0JfXRhTFr3MQhxbX0JVD8uSP34LQAX7t
UKG5Fp9BUrOxq3PkoGqjrkQuRdcoJri/omv1dczxScGr10naLdmqyPknf2X/7L7k
Cl/VI03VamW3lnDJxteNzJ2kcrUgCFSgr3x5NGppq4mzRdiUc5YrF0CFosRRZbtU
M8CUlQLzwlpHxJPplxGZNzjvZgMdETVtTTmF8c8w2YjRNEmXq5jPm7U15LaCbtI/
dE1rAo7/kZuA9e/+LWhqit7Lq3kWSTWAdxsLlaLRcRMsoWXLxSJJw4ovRdJKgteh
TRCF++d6MhhPlp0yJpOkIQy5dIszOGkIZLwVRz9ofr2WLKfhNlQYa16XsZo+sqOD
gMiinARRSUt7vkF/U4SeZiCl/yUYBwd8e1i94NU42Jekp47y/BaFLM1xUMjNQrs0
QJfRQ/AXW8Jq0hRjj8O5xNInAW0AjgCHAe679XjCXLBtdoiiaGvGsXB0gMKsXU6G
`protect END_PROTECTED
