`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7l2DAMuj4e63E39soa9veS9dIOfvnGikywAtfO9jbONNostyh7zStxIwwAodSP8x
TjxIt6L6L6DUen22MYUcNyFViZTdgft4XlkBgJh5aVrhKm/gIDY2CfUInkrf4KNZ
RemxJ3TikL+vFzy7F+wMOrURiJKb+fUh8yt7o9i6z6z6H34T8rSzzPqizVQPNKkz
prIo0c7wvM/Xuj2xaXPBqjGdZXxawmpJVPu3GqNPenH3DIp3/HzHu+4bffEvKg0R
mZTqBOYd6xSC9Qw7Ro0z3dCqwIXGuOvnY+XvMO3qQjszCu3ONg9KLjvDjbwA9gmt
Usv5CcLo9vL3QLe9wujrZbiBpCV8MZNchPKcACNpJWcqIzeGWTEi2Mo4WXmQyIId
EsfdJdsBOTHWMeBAf7rw3DeHM1Noe8gbmFpKM2wis21gS8BUEC56p0WV4j0+XxlU
0Lxym89oeDSz7B9ZxCMelGtuwlCXOYb1+jsz2WYhpqJzI2t1KIEdq2UEIY9Ee5aM
`protect END_PROTECTED
