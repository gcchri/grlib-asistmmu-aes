`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aHyp29NM4DLfuZoh16koWy9Bi7/OVPYQpZsstUzhrgOKAXLWsVKUTaYBH9uFBy/U
w3Ft5AcKQ/PNEEU5hGo/b3RROV70oEbMbGFIaQFqvL/MpDzza4db2hzMDiSm0lIU
s1XgTtBy4sTFZ5ocHQqVT5VYCWl2NXzucslZSIwhGncwNltkzx84mAmk6giiIT9s
YCp6M1oZv/QJmLo86YdIZzuohNxvfXonNApm+bTExMBt35BWXQV9HWGxHeqvgmFf
w+7nFj9DNrNPt9Zdd1tBgwNwIRDK6ZKxOkA0l1socuY=
`protect END_PROTECTED
