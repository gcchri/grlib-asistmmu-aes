`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CQRx1yfEXgxjU2auwI9VYgeIWemPDo5JyfEgsOvyeBS935WU0RrqVxg3B5UKUsqX
Sgb5nFgZiDfBQMmiSbUYIbrGAykB6MuQPqc0WfUcFFO828agQotSdRaj3AmTqGE0
SYYS0oHCh1DOTPFW8rWYrQ9tL33UWQMhbo0w5DYhxEYhlw34LHjO7R9H+g7wESqU
cEJMTMx0AjN1pjSuDmdhMzQmr0NX4TxK9jYBB3hi4ypmXnOYzetqLxWkJNyjsIAw
MZCIM5RMW6ZYbGfv+BvGCofb/13bW1j59HcfmqtI65vb6CXvMbJTn4oeTwiXOeiw
J1FKshdJAfGTyPvQamBEUQ==
`protect END_PROTECTED
