`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AHUud1RTPRGIvPvF0oEQDqQCS9327GUF8hl6+4liqPfM+4Po5EJ+r8p4PcyAkzR/
OMIK3QkLSpswXO/yVjF/tos/vrgnx06AA6UbOKI4+BrCr0pBtzTOiLNH6sfJRylM
XyfSQL9pTT6t3eOJPLRHl5+aFJ8swUvJsz7QNQ8PQ0hd98WZCWoaBLs7viv0CFA2
5ERlvIy0b7hgeJAYMLUy4wpaTy20PQqAQL5gnA3QJSqBWYzLfxPDJcfV+M/R65hf
oS+YPT/exjPBff7nV+kS6ArSs8gWkXC+d26XMXOevNAmnW68VDZTxeM5Pzwre2zx
hiA5DEZjWzxrDI2IMHd/sSJkgt0mGBM4DtTeLujJdajBYBNHhYmTzkBn16oCpgrP
JSTj/qs2EBHfxNMU0+G5FyqEkfyVcBXDk/ln/bNoCSsIO8+m+25bX5PRtm9lRt3j
ZV3OyGySM6TMfpEi/LWb0xb+7Ir33DLQ60fBG2RhGU3Cb63vVOLS3PSQaJAEiCtw
qz4n5JWu7YEpVW9QyHg0JvlIkS6rR6E/bUafqV5MazaWIB+EE7I1TMWPX0eZmLJF
SeeVxpzzPErRl3n0jjk8Ga7L2FxSurLLxOQbZrD2J20kbuygubyu2dzDsmT9qZTA
Ei0mOwqsJpNeEW1xNWz8toC2sY5T5dHlndZWCy7aQcimAW+xqtzxX0hTt2ntK4IR
u87NFIAcPIwFQk0yXD/JlMMPmN2IfLxR1lNH/PnpusRDGQgmsBFggWldIU5+9yLZ
gC5f4B70YMsjjYT4MzRtuRmaElyCVQJi4Z4aNYpoPpD1cAcxFIrCbYFUb6+s1DlX
RnNOd6N5Id9M0NjAZYvR6egGSjtO6Bu+3ZA+9AhRu2niiyLB2J9pEyTUC36BQa4o
+mzyQ/fjevixGI4aipD1LMWd+5R2kUTKVbKphd3J8YU5Hg79BPnnQZuOjD+Xb0Sm
9tQl3gbHhIgrn3NyfdocyQ6u/jxl28RxD8Gne66YQFx2ywu2xLZP+0/uEdc4BbYg
89t6/odcAw7IWnC4JYoITG5nHMgjT5sLkQ511bo5mi8=
`protect END_PROTECTED
