`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vtSEMYT+cag8/4i2ebkXjfV0ahKvXJgGKviFZ9GExid7YahqyuAqUeQKyGm9N3/5
NlhbTtSx81ry7F9L6ay3OQezMYFDQfi4AvEyF3WriFXhMy5nfa+w2p8fWhJfpg3x
qGqVDGkNkKYPLWOjf5pO4RnKpnOMIDoxtmffoTNqGQbBFHQJvB7391TtBp3AmQj3
H8ZV9KbV8/uxJrwrDbkDdIowITx1OFO1XC7WkqDn4nwiCnXDl2SDfxYq+QqECpqY
bVa7u1fMBv+9me4vHkZzSh8dI5cf3SLhAhJwDPn7Wb8gUXAfFZMl1N35EQQYK0kY
PUiF284wlHIQRUGdQmVZXThAdReQaySwqA8Osdlzn2zyH0x03MRuYEOq2tnH0HEo
nQdA6dGM6c5pZLSkbkWvDZ01cAPycSoAOu44IyFoF4r67Cn2qKpAKeIvgetiviwn
f0CznpWaX84co1mG7KG4Gf5meFjE4OOBfSMISyePe3GrVhWTUEHWiP4pxBuQy7kB
Wxw55NDDp03tCpJW7sKBoypKfWKY/Ev+HHSim53PcSwo7PrjO+VJp58zec9WQXF+
ceo1sq2qaISTK5llZizpumo7bETcIXzl4VSiz6APPfM+2KEnzGyHVtP7HeRgAVkr
DiVoed/CXKKpT2XkZzdmbskk/dwfmXYkJzfGEX3TA8DyqVo5E4BglRU8ru+XzWhf
FNFHNbANN2TbQDe3A2jashCDBFqau7YM4biROPbEmnWWBvnACoaJNNa8ghFGpxlg
izA5MdsLfrU7R0gtQ1SyV7OscF994gUvjPzPZshAzm1gECCL3hX/hs8y2UJAwX4H
nL+5vP8vNt/ddjgpwkVzX3uMQ5f+7ZqqUY5D8R2zil+nCLVjYvJXY+SNyDK9gx+P
y3GfYGYxg1aqzToNX+F9ZEO0gCQn+BlpCh1UVtEOkGNvg2+YqPPlRaNdtz71DFas
9CRoc0APvpiCYcaDDaKFwwF33LiMPgzMSqBP5+YiUNtQXZtDCqrxyJ2B17N9tXhx
YXQBlD84h24FX6XQ/i/nedg2IEUCt7pItitRH5hc/SmEbt1PPvGUwHtrECgAW/D8
uL3odzmotkPo6IF3G5QsH8Y6UTWPeHsqma9jHk3eTME=
`protect END_PROTECTED
