`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5H4TYBOmJS3rchQddnoqU+MNcwsD8qouSs4KRKuY1eFl9f3OLXqy+FaD/qNCzJvT
Vr7YxVnwI47IqAeu4PeEsbZukrGcMr4+tFN9efxw6V7QrvWz59uO5juMJF8Xvpo/
WHvrGrGlG3PFSV0XO02321gjThYNYT0rpq6/s/RRoS7umD/2xzR1fAV7aOS/t9Yf
iEz6JhC4kHT8fDzUm99juWlGVeIc/eE/e7tvNf5KgDV9poq3Xqzgy3j1fVLJsShY
+Hu09v0yPBXSz8DJqIdhNlvTjAm03xw2JS+IwCRtyQr0a1hA+p6wKrUFEVXTsQso
`protect END_PROTECTED
