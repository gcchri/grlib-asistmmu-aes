`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vWpB3DocSFFu3uR/3KWgToNa3elGjHnoHN730wsF+gh+FIoOnhGx7sbfg7sV4HgJ
skpuQ4k7JBW52AcuZQ3WEXPg7wRAtl2GbFr5pNiAZ1vixlg/1prNb4cASk0GMppw
B7UQq/tx0KvU1tFAuAiLQLi8Ya7Y+YUi9UvO2Od3pYG5ruJbr2DrSFKS6FVu40ba
jvPDAf7YXy3aDEZmQRViFtWmpfRE2BA81T4jdw/OWdBx5eCvQWguCoiWfCEk7FY4
OVxn3jVSMvDjNzpx05aM5JScahEn8fgibUexD9ehZg85sEDK4bvhGceoqm7rKYm2
TC1w1RoEgeu7R8qSlIoD/4VvNrbLnY0WZAU3THR8g7forYeYBCWqlesU+aqxNtSv
R2weNfq4XOg3Wm608NOca+j1KeuMBYnRcM5r53sY9HpD32/jCEnzbgo1o3LctqkZ
wbByawWeS2ehfUOhX8G7D+mxrp70AkqKwOrl97XMx+BsgaRZpSIB5QC2hk4CWy/B
6OTY1FAgRqDaj625yPn0VEd2QSlO5qRtFlXOeOttcROfA++BsyAPwfmVaVKctVHp
BhPn9uH9NJSGq1uOVwSv7UykU/hx3LPRmVcA0VYZ1JtF6B0rMk0upuTnnwUqjGi4
xTW9JyvyUsMIBkqCEvV/b4IfsaTtKbqKcVmhS6tDUs0=
`protect END_PROTECTED
