`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S3n2QU9117C1sy7fbZbvYIlbp2jFMOwX/DPqlHBZWAMjUxORi4CX7k1gEoAfYX/b
nLOzR5jAASIDiuijkJB1HppfuifRi4PwCh8LaF6OtJoElKLAFaE41Op4bfBe9nDS
YL5+/7MB11m76yUhYNXFCPeW5vUQ7mOeEpJe24vbrkRy6iMcmyUJFtHdw7b0xGwj
/UOc6AP/k0eXYZR/gFscavshQXgb0z0vgTdgWvO9wmS37sA8SnCytMKefdSPzPQL
X8BGcnpQSWDI8L8G7W+ubcpc8i45eCZmOik8kWSSn+73sCZx39aI6qbY7OeY93MP
ndZUeoLQX5mwxrWziJYWvqW1WvijuhmeDQ/0/EM0T1Rh0k75e88C21nfq6UBw8cA
t8PcR2DK7pwPV4yLPWY6+zz/XnxqWOskGcKTyjylTcgqdKXGglrQNIAAwmGwa0F0
`protect END_PROTECTED
