`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+kZ4yjvKhnThWTzhklxvNNcc8y3MKqiANBofYMqgLb8Vw4J5fQpbWGfjRErXE1N+
+nyCo3ne04gWsBtUR1WuiyGW9P0DjeOMaZ9tsa2C41pO5hmF8/kJs5m78k7MXG/u
LUedf12akSxNh/F14OHO1Te736RO2ZRMit7qeoFeIp3FO0IxQOyo8QXlaTsWoCtY
ZsbIAvRi5qRgU0MXKWVPSvurqaF1FlwjPquztuWmGv3PTAndST3YX2M80BcBmnJW
eG0jZWvmC19OVy6R+3H3IN6w3engnqphYS+l15QbUP0fXeOBnU+zwkJzlj1dOpQr
u7bvrnzTX19amTUci1JQ8A5Omt1WrueZeA9xVuMYmyYqF/4+/265aCRFYkJtE7Xx
IKaR0Wc3mJFv+RDsLQ68zV0cmB1S8bvWC5Cd79KqkJM/nvIj0DFRx+TX1xo2Qxtc
9Hu+N3onEFpDND5iuAEACQGewXdhT0MxB9sXIehO3ml67lW0zWc6VSKM7B3NIO5Q
OcKokY8SgJEjFAIAEhQ1zDF6ezCKduXI6BDeiq4DpcWNOE0OMz9cN6X0JGi7wi6W
vvxu1hzeF4FJSLltc+C8Lf0lGCpLRXEcUZnt1FTPPCLTCk4BsV2gSsmsUd90CMRq
zr5FGcFq59MZzST1/kJ79/wlm6sbLHF1Yf2kaw6YI+0fzLWoCmqKKLvuiQ/BkWxW
pfXLBFq3N45spMCKGxQJeduiAGfg5ph/Jh/YFbFnRsPATa2XJaFSQjJx8diUQLud
v+zWOJO/mj/dRtrq87qniZrFDiVlBlKhHfaG4KMEfP12xfiBIFPpvZ8IuVWkx6jU
C6YQH5cXqx3uh8vdCHSPfHcfuLTfkqYaR7D/kQw70Y8NDpYe/DquLmWB9WGnEo4Q
VORArTtaVlYSlPSi0P1oOyEnwXb0it3YRvLati+GC8lfvEU3Y5zBuxASQDAMES6K
MGsW/lORstbaSof5UuseSpVVvXxd7NdEd566IupOWKd6iJgBW4FwipgH3TokVtFg
`protect END_PROTECTED
