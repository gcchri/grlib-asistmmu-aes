`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PBCfta/JR6gZR4057AkA/HFum4BuvGmdJIx5X0hbzTrCLQXI7Q6DD3TDWItPlNd5
ehJSY/c9zu0XbBk/Iq8XGY2IdWHFQ86KSZ+rvrjoGjb+fjEihe1IivnWLsUALi/W
f+f0xnHLOGkk833O/zDQg+NUAWpVOrO7naNAATBC1May1hxwAkEaVSv3AFNhMlIq
NTJoVTx3gCp1gL8WXaOdbCYhx60yGGdDoCZoYXBG88CreFb+BScCtFR/KG2TWjtn
o+uM3W3jqBxouY94RmjHtgHhDfSpgwOl8zdBysaccGO4+0tJ2SzEVvfwzEc/UqZS
`protect END_PROTECTED
