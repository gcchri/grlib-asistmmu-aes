`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KBowUkM1pQQd1GKdeS6FtoZFQrmw9aimoF4+5vb0TqwiW4iLTMKhn+W8/a52d3YG
Oj2svofOlQ/JSc1ueDZh2jm/oQjENYupiy2Ag4qsJJIbKEsTlumUxReOOCjxs0og
NsWBx/vMNSEa90/zLpLa1enxLonPqQ5k1erIMDyEJBiQK7stHqVHgyirYRnVxirX
A2JoWQDH14YGRR8fWFV0Ek/Vn0vlC3JdpeRLAqte8vQQZwRrJt0So1SsGGpamQp+
Etk3Q02uNEDPFFESCBhyizkP/FtoKyrWKBG0Gt1Ge8WSUJd34n+DrztPVK1BEGrc
nOuemvQ+pvzEE+oIFs0VQtbycO5YJjtC/54hXN9WGI2yC3gTv1Y0h6NjrjZPPrdB
qO35oxkfjLJ7LB0tHFBUrKqj1obpa7HJH7HicKP85UxmqB/GqOWHWfUBFx21QB5k
QxKiYBWciy7zViucxLpIL8fIHW0ICe5MTphAIt6E2hvyzdg2gToe892cuel6HhHq
fP51xK6J8CVcwfwi3iuPWgwjFQd1rUgfFsjmJQlWSyEpGiNYXA4n8VeyvJ20ZlTC
qz3LafMrA+aYDVpPXCIvMbmm6qZthJize17/VV01k1w=
`protect END_PROTECTED
