`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tDvEvDnmVJz5+HyR1YZ/LlvB2Ao3OQI5nIjNfRwuyXGv6dmVGXW0GNzd/IAQcJk1
QEyOngYceMbK5ep8zBZWLS1G+BA+e7jFuaWUrJ8Dgt8+8EMrpOAz69oqxe1gwiIO
3Hk5O1sxDgAQIhwX1FtGenhogxGOFfzBxpm4UHIrWlYTAUqmMSNEd7L1wLniuD5G
1RaYeBlU4AfH4tMrUba/p0jE/PVAzPr8rTd2Bepxw3Cu9jaFsfDiXn9fWyZ6F6Ym
E1rF9ublYvL7k+6MNxMQmvrZOk5/CEaaJvE+KR7L6KHCiI65E+ybb7DRTrg/76Hc
sJ7a6CmbKQhVrq0e2RDL6HnAWb3IBJxM477ljbX5B0HSMCEReMZpw0MqLgnyCv9e
xh62v81IRZNqL9EH6yW26AOS+YGWvwFhkjA6/g8x9t3xfqBxCTTVipcYApSNKBp3
KKa/NU91pAAiOgvOM0RJO0KThXcDs+sJ+NitlBfNqbGwCTKq02vFLkufl/iqZV99
4TFIlKCZ0G41HfwFKnHpUGW7HYv1AO5fhZtACkR6OHQWanT6PA+YD0PUtjK3Fryv
T6aMdTkaPXzRN9IS/cn8Mdute2/on7hMfmpQjVWpM3hQaFDVKFYrB9VFJdlM+ioA
hDTTWOTSY1x4jbQaCYkXIzVlE9zF4+oixIuLO/20CyN2djmcfeR1qx5DeIR3u5E0
Td+jrxFd5chyi6AuShYwMKishJfAWPtQ0WVcs1TYCoQ3IrkVouICCB76r+2AWpvN
gQ+yFgWXMVPSp9XB4oKdB139WoKMKrl6vW7SC751Q7/zzriINWQo8L+Huhu9WHcu
0iIprJ47G1c4v+T7r79IbDErRmA0X6EuKU93rWSLoiU+fYdRSqYG4CWkPC+kN8rz
UO9K+nCgUdwVRfbHlcTpgo4ewi3awynt23DOfeNkbrwWuWbq5ykR+/2Q5a8KEtvM
Idk2cKmmjHhlfx2U8VaLQJxEQlmMzKpZLXIQaeqECBadZTHwuEf/pZ43A9rFHb/9
9jaDCINyMBcavKEY25gn0D9EXdQ5aOeG+8qssg4NQgSy2yLPZctFbMIGl0oaignb
h6boQZxkXYiwV8BAepPZkZS2mXMcVhyqoyc2gb1G7iG5LFEi5+1mI+SSp9GwQJae
iqyDqhEcEpgo/ox429aOr/O0zqURZjrLQT2L3jCW/Vqu6Z5V/MRXxUu08v8m16xl
bBon2iH5e9Tx28nSmmyFRj15iTgSwktLN9U9OebBAHzryZtWZ9WjNfn+8JZCu+wn
TN9XVRki1RC2z4DRAtQVBFAsc1zJYesZ5dtEZ0+m5r0sP+C7vg0+EESIg29HaFox
lSPlpqKdtaC1HSmoqOa7rzvZO9bT9fCHCD3Zxehg8ndbHM5tFKR2cCXwnlO3fbmk
7Krg6/654skmij+xaEJM0OENgkVqegkeTWtxlY5NHhBKG39w3h1ivSzYLO1gxfzT
SsS5YXe5GPSqrFl/4Rj89JOYNT/N3YyEB4mgBCUtua7xCAE4UepX/GyjYPklFIK4
Mc166ilvehCVvlWhEwwnvitNZKHIr2PL+R6t7nPHt41zMWB6oALU3GvjfUJQfo7m
ZvZk3VdZS5xOkU4QOqrwVQG9D4f5X3YQfw1fsiNkMHg3Kf6j45RDFmJRmRIyOSeX
ow+BGjiQUe3/0N+DkcHEOYXked7/WE8PTMCQU4/NHxqGx/QSg1OZODcAcp/tTtkX
D0QaCn6V8HVf+LEeVapxfPJvYiT++kHpQX2MUruXDKFQxenqNWT++Mw3aXEf/Cru
zpGiW3qwE89+LkBftFOR2YxlDWkWWchIJP9PFXYA1xAsNPlM+7XV4Tag2XuiLBEl
L5ltHx5iadzR2U1DKe82TA==
`protect END_PROTECTED
