`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
khQUi/wuDZFVdId/lEWL8PTEKabutG4g8uGJsUWPtozwvAuNMzjLzi9+oUK2pujl
k4dNuwdnGEWtAT7QFNXRSpq5U++e3MsN+CjqjhiBoVcC5jt+zirBvR3WIdy4EogJ
xHGwG+qaimtT24Ac+b5of8T/VYEWlJ0OfhU3Lf4OGmbglvGodoF9He2FS7o9kZpK
xnBpA8e7b00/jIGkFz1wIoO78jdu/jhc0WCiz3ZuOZI/+SfXfX9d38hHWTDH5cBB
gio5yHQZZodggnBWjHlEVUnsB+Apk9lSMDQnLu1rOA8E+/fSZXqrupN6j+x8HKTk
QnUQZjqBs1GQHu6okBh6TjNHunIAHiUFY7AvKK/zd/Dx1OFhPE0QWU2TXDQyLV0X
59OdxQNExkEiIH0Z0WS4ZqlqGsW1cYuy08N2gKrvlGRk7W6ez3s2UW8FsLorqffe
j5fLjKJ98N+IOdB9jSfSSwi39/CIlhFyM2WC+TXeNmntVG1GBvFhzaUm+GdEg9eD
mFhFe0yARMJgm5YZWtlxjCZ+pVVKsQf1I4zq03hDiKF7r+hxjDG6axsXGAbuoTZm
CGQ1URJWQmgNAPe51mz35tl7Mer3XNdCuPk1eJx1eK4035hhu8h3vjJYdYYdKEuT
Z0i4SYMELJwKAL9pEjqTlkn/5Q/TWI9w7gHI2um/sQBAT1yJtm5pWNYNvd4WWN15
QOYMwKoL0Y85k+Kh6y//woym3HeYt27WhPb1JjAa4To5fkEcqr4A3Yh7IymupbE5
fvbe+0s7tp4i494Jx5W3TlLmeQvUXD6IfCpP4v8Bo57iDywMRHMZjoKZc4Pz+P4z
7xQHsrtb/Y3l/mOLgqxbtrOtDeaykBJsUhjFWQSJH4ZSdpcbLyf47vzqVSxDaEzy
Mona/AKAn4QbaDR6R+/QbockB3mnotNjq2f/4FekXK1684bFM4Yo5jRDSoe3XI8k
xLoU/ehyL2ez+qf84Wrne9EQ+TAcLIUrGe1I+F0emUmovlhjtznlUq/MqTULlK42
ZC5XV/9DUtBOYpHxyxgo8ruEncruZS3LXgD8n8hwNrSmeqOgi0C4hbUdEQEL0EYi
CfGsiF4TdMfuXUSuegZAN10uFjo7lZ2ugbty2e7xKofc9MV5XHEsu3BzZcTQ/nB5
XdPul6EGegxaWC6sIlEnS7TTn+/mBm4bOKQuMjNaySRK4GDNZe4T1Ai4BiqLIKkO
o9Wo/Hrv2csDPDE3YlPzeWkfp7hhgQaMbi21El6pjD7eaCJn2larIePkBuONDAEA
t4VsOZueBeF1LTkEv/DuPqsn9An6JCEwaNFFM6nskqNlzYH56QIqj4VJ77M/8pxr
PXt1EzuDi17Uqz6+4lF3F4OWBb+zcCy0vMw9MC2OyAcL5otHTleCaI//ZhkyNifP
clDEysnL9kqpjgNHvWA957hkLm8WwTHsNK5MkuECAQ3PgIQROp02IA3yQJ3wWrVF
NtcGJSjdq9STY5/AU7HlhMFf9iE0SqVFK+++LNE5/4reAgO8FSqrIULEt+cHmyZP
IgiD23rotTIb/hFrSFajW7HCFEkxwYpJx2rrMj2j4k3RYHwjyt3H/Wc5Y6tdvRm/
VthxYSjYDYUwzo/+BPStwbpKXXUKFXJNY5KOeNTUIg+GQMgseueU4AjTkQW67tj4
77N9JabaszXhhaBsjLKX4heYetvvL8Ocnuws6Ps7l8E7lpdEFOgP84gl81C2gORO
SU1kIyCnBbO56mlmKyOutlYnEQc+RztJYH62nQOX7sMO9cuEdFIU6MIAA+av8kh6
I+VvvoSTR7pbT+OmKw8xfdj+bwSy1FXBJWASBiHP0v1eUiyAvNPGzrZ/ekEWe8kj
UNfUfH1P6DXCXX6y3b9R4X70rhoExFcBRGUzhu3BPIX5o8LT9lm5d7S5nptKZsEv
nh7c0Gv5jjS2EkDoVhkF/Qmk1pqICvmnT3mG/CFCpl8FJZ1Lvkaa53eytlHKp/u/
sY1pHfv/gjIVteka3wvXOQqbQLQVg70dy+9GFqy5b6tg0bLvJiV3AIWUcQb+wVMJ
sN3Jk5RO7V4Oez3lwc+QFE1t6Au3fmXWgL4rcmhiR8GTHu9nTMVnTrHTQUhwpCuk
RqTst6kQyZBLW94hUGNCnbMQStt64WFK6Rnt2F1d0mn2nj+/tQT5YEuj6IqwwNub
+arcNYtqMf0vDVLlkhx96z45/ldsBYWnmikxkEFnhOcoQdvdKyJ5s2vbfaL4hgmX
/tGnsbNORNq+/OwKDWsmyUbXuYKWMm9UHLrBeby1CfzWD03n3EA4IJo4LlBCvPUz
nmTTROSIpCZNojjvjjUXRnf2QVoQuR7AEHa+eox22LYT2skkTm27eP9r2fdLLf/l
Ya4k05RjPuo4ZQkoiPxFASb2kIwB0TN0vVYR4JOXODST14nokJEP9pq667IPnwas
EbH8dMLyKRNhSKL70qB6FbAbPA4Y2QnQ1M75gjeojY+wdhEA/ynCJsvjD5NhBs7D
5HjXQ3z8Xudn1md5qO2SEqjYWvyIP5CiUl+EAkizLvF+7RRVJl9NORmlcOvhR6nL
U9HCtnEc1bafvahmJ4pIxraEtc1IQxpjXegBZB9401QEuILcIEu5y705elduByFs
nz92CM9v0JBmpgSONo3QRg2x+LZFfGK6i+fkaZ3iNdLEXflS3GJiBj45o00gtwx6
jF35kUhykyDKNmiIA1zmAGviJOCwN4/7zrslROkHn8HvBxbYiyvWKLFGqDYjYX97
A8QJMr+aqUNquAlkMdTteU0SiLSgRimQf6+8jyL5ROdbJhRPbGfiVkq+JQX4OyaU
O+IyqZ28N+iR1yysiXf/yRFh5YM6RBS/kS/YMZyz2Fc0nP83f+Ys2K5CgDrCo64b
CmNuH8MSUEduteJUx/wu+izt/qEpBgQMKdZEB1+zYN5afn5gOr9U97r3stXHln1Z
+r+C/r6HYmVoJMl5NbmCjAujNgA7ZqdKuB9SC0Vcc5nUFkQq0F989D5BON/3uWba
n8cQMQIzTL2spNi+WiyWuGqa5f5YN46o6k3+2462Dqng1B/pYGRDi6s0Fh/vqmIR
rk+uLZCmR9EwwoPZam78HY+HVESI27lfU177MOoVZVi2Ex+FjkWFnAuvlNEVKvSi
ekGnDEkXA01JOSkbcTUwg7t3f74YG8LA+rgUeH+i4B7RpY31jIQUime1nGsilVcR
0bE/dR5V0HRnQjhIcLLrLH4lWpO97sfHiQgG9fwm3Uz6yxdCraTNLaRZ+8v769a/
6DfjE47v1DY7RMsvOtGKqFiU1FodlssUSH/vkqSZ/PHel891DAe0RNxHcfWOoX59
rLtrSWr8AM7p8F1aQbYx+2CFkLqyoL4N/a00JO2loGRFMho8mWNDbOTXaIwy6ci7
sUAyuA65MV3thxuWkK07Clt07M6WThLgk6fWzHDq69ua3otw1fHWVrlXxiPQ6Q/g
Or60AoSMY99ewjnZVfRWuZjh4bMpDCuXQuGx4FQLe8WNQYPeNl3ks3tc4i44A+IS
iuo25bu6zn2BaKZZjn7/hK015p4ZaYVNgBA0SeQaoFususeRF46QMlmvt2DpCON/
qQ60gxyVZ5HG5bOxWBgNpotuSl7gHrJfMR2a0/cte+JBwzFI3IUknUeo22lucthG
cprjY7fIbX0Sg4AZ6MLIdqpb1W5wM31AHQBvGRdhDACsq7k/L1ivb6pPbvcPLLRS
6QqXBYRhDbx9JTdbZgfIKotDfvwbnaCEhllgG5TLhkfcksAcE3OEwrwlptTb3Md4
sYl00cJSA3jI7Z47k2t1hU3TmnRMiGksvPG/0kr5E4+3gYXaRNLQDPVG5zQ7OD9v
k/Cg35OnKhSjVSUUxEGvtB9ncbM65tGKYjlzXUUEJYVL3FXJriWv26LDR0FdPu7j
Q/59xnPPxq6lVq6ol06apCOEbIEyThiG6uITjCEuj0djx39M8s+D7h7905gH1mNw
dxPgK5gZ6fVjRQfsFDRs+t5hN2LPots29ieWd8IA0LcY9ZpsZGHduckhwBsYG4+d
7NGc+MLR5tDkyGWu5PehhyLSkSEJvaAiJnphB+RRT8IWznbsB2BqnLMVoaJauejw
6VxQXr0+IwKg62CdQXLZGPX8hMHlc0sl1LgwUlrQCgktT5IzH4SKxkxp5bf5MRJY
kQ+IyVyDSpWdaYgHciJb6LRtwWp8ORuZqmfu+sEA6Vsdkdv7pax7V/FFCTt2wTb3
TgREY2OOzjghSz/rL5sCmuPhqLI+ru8SJQ3Js7vi0rAoUjT/Kq7dEpKkl8QYSp4p
IcbvSgYODUTg/C7SwzwVnKDIEdFbgIfTFwmB2Ak75uWdgnM/w5H9z0fiF28LmDG/
EYbNZRoG3i+2ShvfyxXjHFP03iXcsIeJuu5PHmU9+kOvF3pCp0Vu0RIaLb/h0Ng9
igRYA1TYqjJJj2WoCSqMWiwfoTB2pw7srD1P/y1GoDlQQrHW1e2AqFTSlI6FYdKz
nhdX2giCFiCJGcBUiRsRvCEGvCHLwQZVDzQ57BE4ujcPJpWrAey5cOrlr/Gfl9rg
dITkEB5KGTyEyh+PlolX2Sqprj+BPfTSE/JvfqD4U5amH0cw3DFNEyk9WbflbdeF
J6RTXRHFystYQFteH8gqehhJPqNGa+iq56ow2MUN+Si91dPF+AQ1jPqekLAQN0Ty
OkJwU610p43qEUK/qhrdJlzY2tOzXmJVXEYzXUnG6l/pk1lY7pBittfVwV5xFi/L
O97dRh8N/R3usKNizsyOn8+8nD1DjeCtVfVg4aaXPPqKqlpsHEpKJqeYL96UVOFk
aUVtSf9jI6eUEYTSoHxLoCo+xzPCZkorYKV/Uka8cKZfYLNltiqc1S1Tqd5DhW9d
r0cyo7vMEranWVBryw84WyuumuObkcurLeQlqSrfJnc4aG/J4dDlSzqKz5WuTkc7
Ft2pNz1W56AmCRvSYpvOPTsD164GRAD5fdBY44cp9cdaEa+iqkCS7OMDlKm2i3X0
b1/XyG0BmUiFWfSJNlAV5v1klGDndk4cscuvePqrB6WHsm0Rzc/9DBHmU6OmxfxK
hH245uqBkpyt2YPEtGldofauigP3IKl3SS27a5p238ePKSY92scGiP84kgV+Y04w
Wdu6wWl2JW0/qHl3FM1/9WiNES4uwj+cHZzQZcGXPQzLE4EMCIifzbAu4AxxHcoK
+OvH6obpW1wgaH2iVpVF3psLYwkq1lSEAuiz4bL6GgWNlQWMOkO3qNOWw1OZm1dP
j86dM9r2wEkU7IY1h/VLGhN8fJMudsYklvenINyl12s9Qc+OV3B+IDfnC4ksvkiD
hT8ZFw+d9qQ0kqYYt3Svj+3QvWqFr1IOzqe4G2dwhNurHrCDSyS4SfBtnOX+2WJL
X1aiIEf2zkjoeU8NmWIh7ErnvTEs4fQ85CmkgbwcLHG0ctx0LnYGWDE0BGjbUInd
Fy3HdBXyXG1egjiWhcU2agGOifV4IbLB9bMBrcF+sLTx0O/82dIfV0Iy9cQYoW8c
+9wvTYY96SZL+bpVYpa7xfIGog8RgjXpYBg6QAEddEITdt6DbtzL/Exsr4flCwCt
lZqJTMBd7REv51shdTiecO2dFzZIrJ4I1CTj4K0VZ9BNNN13/3z8zokBNfaMOj5c
/7iCAnq5pc241EvGH+SEDoz9clOmkrErSD3BGpkd9fU4OOik/QU1f4Zx2NhkHigi
yB1wtD1GUWX/UTcry3Wd0kdfwNU99v/mN5b47gciL7HQwrYaBl8yEiSh/QAEgsY7
I9k4j2GngJGkJ4PckrSfBruistGVj/ZBxvzLPphSTVsCEZbJyR4ZacjzHCxdOMSF
3S5a3msNlR0dkSpuwK7bR8Qf2CN2/PxVfJnvGZlYwEJlnTv7FIpvAQA7eUBmBb0I
jseXGYEOsOR1KbCUPcU6Ui+xcU+7URZQWWYY3DnagSuiMNBYw4XikBvfObPuHyhK
D+kZN1Adrt/nL3KoyiK1b68620/34iyfBjandw78mA+ADV+kF98tHG73mlrKs2W9
SxLS+dMPci589SDZu74EQnKTyC4SCKmNUqaooVRavof190QBuYUk98+G8s7LrwpH
pHtHbHk136RLgPdn4zrvSDX6qlmQ1rMarbcsyYz3ULfI7KKqQoOr3BLQbtJa5nlu
dtsluuHzUEq15a5FkoAaQ1E6YpxdzQXLcuunkIF3qVsfBmieJNDoORzeslyRXqC9
k2UdiOFH4+Sz0LgZzNuGAsTvNX6LxjY3OOkMg/8vQlEL73z1ZhUV0HZEomuO0QR7
BufQaOnMeOxqIc3HGxosRb3SA8WSgk02rho7HhFSgrq7cOpJ0YMAhO8rY7g4+LvI
1pmOgotiK0iCb0ZVi7J3ZhjJWxkhH6Pe/YDRja9YwHKHFVGZ/gJWWL2c1wnv+PhW
afNuCWEl81G29ZBW/JyUALxBfP4jLneNiezf0Au19mMo4Z4SMC4aIY3lOvX2o4Ej
D1QgvmeAT3Fywx7mylVxqrMwUS0mxUs6W2VlhwyNXu2SVF0CQN8No+7v71+Ga9a2
DhJkDAlUO+4alfycPgXdVuDjvgeE9Nyz1iOdeedlkXl0w3SAnqTJbYgumCILhR4x
ITtffW49dxOs+HofkUOU9q2i+UBOET1aHdLxqJzEE5ot7XrSC1i/ViVxleq5t207
SF9wuuwyNuBat/R2W1X8ve/YwscJuZ88FrJCYp7Ut4Sz+kHmkZX/Tw72f0lyRsKQ
LU7oslJK3RtVTFI4hZrXbvV3XwPgC/wI7+LLI0Gb/ZHGdTUVxTIrUwxznPXKQaMM
ZxXG6d9Naoun381DFk4CVj6J1s19Rm2pc12p5DjvIqlDUtc1X8BhIBzCwAhFqmEd
ZcjWVZa5mjXRunVm6S2jddiWbg3haeavsIirdXeoefNURi7sHpJATcneGV3w6Zi4
2Oqgmh/1GpaRwig7LwlvNMewe0RaVtKIMPnoNbvZBrspjWDLNC4EvOJuCwsvsOD0
ukw64TKnfqHuraT5ECjlH0Tcrckw7GxfozVg/g/qplRwqq2V6OOMoJZyePBfm3ok
adMNXcPYH8mX0I6TKmop9336absO0W7MOj8Bb2dAPhusWLFyhmGhVHTmHAU62qlz
QF0MbV9lHCeZ4jegNWUp9dMuSqnnbfZ1OFW7yLOQAPrvm2mQJojv02Z0l3NTSyqa
FjdpbUptYJSfziH+/m+s90IOwLE+melnkJA2Bz6cIsvM/hbpSV231ZSUXzTytNxV
fTT66m9q9o5gTqeKjV/gdqXee8Yz222ZXHzwS58lrsMnbKVOhco1a0t86rtMdm0C
tAcRK2bIc6s65RrmCE2tdx9z+/AP1U4ieZES/W1JqMOUqwlRzd2hRIimem4dk4JU
OkhFIWyOR3s/I2t3FC0z/nfjY20hYDzdfaCvgOVsAdRRW5mq2tomou7Xl/AbyDhk
+59apSbGIT9YssdD1yDtnbBeOOJ+i8S0nSV1FpVKKtmHy4r64NPkKXgM9WGo04Mj
dqIRn8UxQV6t87HIi6UkDUHfWhIOCspi57J58uPqJlmyKcfICuhOCq7+ey/eMJpB
7kyz7C8QbGFTaxwAtfzwIcWsPEkcqLXvTld7aC1mUcqGHCnR5bCaZJoCD1q+bJW2
8g09H8m/4VL/JnORbZlC2uouEzrBohu/gNtWNJWCNbwJ0+3+PiC/NhWTJbvlrYKF
yNBSpk60usSrxX7mDah4PS2iwbxy+Jn+WH3Urf0A/njAC+eAHLYRNqqBWh+lcXzb
b3kTr5zLvN2g0qDUvI8y4dzumDTMT/P/ZqU3GsEk59QK5rFYXM/cV90I25pmlKH/
XAwW+peGuKv6iuxLbFWr01VazEj9eowsr1bKbagagw1b8wDA4HfL7bP0aV5nzV4A
D9bMqI8Bph4TX0JPaZ78tyLEOb/37WrENEMlfr3hgMrOYOy/jVRd9tOosHbmE+a+
j5vDcFeaOpMlLE7b/P+ambz6eUiTn6mno5+fpZAY/XINxednBc7F0sUY+YNrnob7
xT2qaIDUljDjQY/gBBaVGmUGmyuEctYvV3QKktJ3XusOnZ8kBqACNB/QvEv4Ozvk
qw0LK3xEClzbupc8xnA4DBIKk8/jBoNK+d9ziYPg8v7yQG5AUas5DkZcFq24NEnT
sXkTiIt5M+ogCjzcnO+J2uabF4OMrKQeXuZ3Kju2kVzc+QIMskZT4EM2M/X3zQUa
eIOozR+5jtDLOcDPgNDul8+rl7i8eZIiXUjrG4/TsvkX0Aw/mMJqHxcn2OU4H1lp
N+tuaDeLiYFuDamlGk9WWBPPP2nD7vQvUeMnj5IxZiYTvxQzmq6MNxaYldT/30R7
5IxHrzWh3SIKueEeLUVtN4ZMZPL/YqqFOaf7iZrhiJdY5vmareA7zHZafTFmOnnv
kzDhhswwcUBGgL8OQZgU7JIVa8pPZpnvYEkruWL+ocrm/xgdWjZ6b/QMmJv2cItO
X56KBHKc+Uv1P5fi9sq79/K+mUTifgh2aQeUDQ20aeC5QhDMZz62hjThMOF9oe+N
2fc21NHXeIJpGZbcOxhCQL58yem95l8DzMhb0hCovjM2p7OPlbcfotGEB51439g3
pzIvkn/PUKdGK14Fkf9pkIN60XwnGrhfOB3yPFZEF6g2tmqzuKGncswWqFQTmsnR
Ynk5v68PG02L+iFEatwC2taSzR2vA66X3irG/9wu2k3mihD4SiK9SQ2cCFQj7JVc
w4SBZPlNuBi//HzARpdhrfH8DzulgjxDJ0ZccfQqPZQs9KyOhmVMchljqiCQl6mL
zd63hBJHFkG1UwH1B4EbGNBOURjJaQnvQoiTg8vsSCF5WEyRPXkhJ3VzQ/rtaHn+
Cgu0HdImQeh3DXZbH3Uf1sYKcyhJaO2+HGxz0ozJZSq97i+KNCSWidRbbERCZFup
1OrRhHMB/5naMGPdKb8xZC7+ZpdbmJEddGAiWjl2MQ08r/Q4JOrOFPLKHIIRSsKc
lzjslcnrra4HG/rBZi+CF3TEgvcCOZcooC2qsKn5kM6sZUVTotA6C6/WHBkiFq63
Yqhh7aHhW88s1t+emXpyyxDpZP/Y7f3k0VHlwEftdyTbzYIlXEVhrwaCI7u9XcGC
6ZJB6tGWcFnALBhzhuj/qxu3lHqP7O82mnZGLzJl6WouftGt73uIp7PsIT1lAIhS
yuQSYFGwJnkzpj2sFgyyhDh264lBxviN+J8Nt5VyqomIPRoplXFEwsL1aLKRFG/V
Ywx894BFPmu1Svh7Z6v2obW6CK1xLoCW/f7VcJLgdwnIr4H7HQR/LPnyiPOOHHQq
TSClCOA3qow7Zv1zQf8L4zwSf1yJObRFTQI3DhecUYinuY26KbJ3V6tOTDgRV2c3
b00skrfa1ByvZeGqYQbYjHtoGBHspKZFcDV35LiegiWU0CQ+Emzu4vSQ59obnYRR
GyNr9Rj00Cc0aFYaEGWF2WdJ/wZ6uq+wdJO66gQxQTg+Rtbb7uwRbNsWEp9DoAh4
xSdYGqANl6N99DSzx/ys9vL1WbcVmphwo1F1JxPwxjlD5lPZ13jnPcGVRtfQCUk7
Vq8+VfcoPrDjfpV6IDxeNocQLaoky2zKccgk5/9EFhEY52K16uCG8gBtm4nXlKbC
gNNgclOtIi6tQgnMQR/iC2w83LFf+X7Q/lU4FoKf+GgipUnATQ1rWyGyiusioLtn
i5Lb2cj9MAp64cGfOa9PktbWqpXxoa6Kj/oG4YzUJPnmTpVvAHQmU04T8OC83xYC
+IdxcTPNJdOFjZsX7NSBGqeUZjQVSWleOvr/Yjvi4LUJojZDVkxSxM8KVX4iU3Re
4PDsjFXeZWZrKD93IkKJ4IzBORJPOFYsN/D4mkCWPKkAOp0E9+qTkfjkhXJQwIvi
yvzn9SD1yhCi2uhjJW1/f9Y7LgUrjvp8q+QaErFmdJ8qUAWoXWx/oYqZmxXMqucF
CwKuKbYxireXhUJOzQfysQBFEkE3OzMbZRnC3ER4pyxJ+exaFX2fOuRzBOG0p1C8
0GWxXyhmvf3+40zoSRwnCfh/gtbjrffxPDYH/QP+AQhmwQVGnaw5aafv6H1D6Zz0
mXQUmBNjaYnw2zh8RfLWlOTfExGxQQMRHUADC0ClPN3pvSTvMkQ2/eFdtW7Um3/I
d2K26CMqz2oOS8SI7VYrJYZbR7YQ3RqIXr+/3D3hqjJEuHAoJcWJk/MelOBs7mj3
9qZSoZvJQNIVfPWDS1NTzAFQfdkaFg9AlRZ/M/92T7dSawBoDuQKFnw6xxNSKBRz
lJfZABkFKyXyuxvxYo1y7F6r6/YhRdYJce/2RQc9RLoICGfvC35MD+a54W7QYyYM
KcimPZTb4xJbRjt5O4dEYxZJyCxHnp9D0oOamVKTwDyMMQ2hWgEh3UQyv5R4c7Ke
MIZeq+aRhbTXms2vJ92nuQhl75MQQXpeDgOfaIqp0nfKzQ3KhZC35LNPkiY380ht
9FXkefHCmZDR36tR/tYl+CpYqA56+CwU/XwaQ/0CzQ9feVlLtMr3QSMjSqy29Uh6
gS/V5qV7BBtOrG5o/KQ40A1Ie7q9fY9d5VhxEgdz7F69WORu9KMoAzd5n/t9ARMJ
oSeqEYYVQ5QF3tdGZEnDdIz8gcYqmoHWY6gTD0+rMQwsAYg0imk8v3OEVJM8Px5w
YkizxZyKeaNyOUZlKQoCEuDZdWM0a4Xnfg1jwLqBtxIB70uJhcjPPPiqF6lfDebF
HxCHX4/wogrYfZSowkGLI9KNJjMHNuMKuGeDtrL6/uAlVctPOqK2cNSa2dj+kmKp
m5N+Wupou/0hZsHITGJWvQdgxbiudIDdhe/ZqjJTCKxmPddkos6ihj/E+jr2OPoL
x0R3xm+Ab20nC1aUbL2rXE/uNxygCzvXbWwVHa1vIcO9XsIDULWITMMMGpcKDbze
vVN2z5PY2AvfaMcT7YZ1u2u/RX7dDJUD4tnYbnqDWc6AOYRGFpjeWOR3pxyuJWz/
WoB8QGdj2XB4DjiosV0WDL7kA38+c69Fw1fuLW8C+8+sBJ0gHb0+KM/xy3jdb5+r
zLMNi7b1VTBA04otEO1WxKtxpeiBo385kunjHbsKWXatjU1bLflThPoOOWo4ARB2
xvj75+pTpYJRBTcXssNG+es9h1E1/YpQINxzDHRP9RZdSoT5dpZSRKD2ILOi0LoC
DOiQE71gR/00p3MaHEIFJ9qgZfNVttFlQPFkMG1Yl6uTmgSM27x1bHCxLJz0mSc0
9xHoiKPB4uE9TQDzcbPoM6d7h/dznspoerY3dHl2ORr2+7V0Sz2IQO0+ug0uhY+C
3OIX/FZaIJCsRT8FtK7pvbYbeXn5BSnFlDcgW8dz/Q0VLpStZ2vStnHq5VfKeQtF
hxpgviv0SnTEkuPGDXGGX0xb6wZ9QJhLkQAO/JXUTVOR79/KLBKHCuGQan+dJHl0
pBs0F+n/iNBZHUcRIeaUo9j2iaB9p2CTdB0uboEBwsMYGyXTVEbNUoKLVm3+s7U6
CS22g7UE+z68aMAOohw0Mp8pIcQR0g4oSeprwJAmmTQndXFeHJCYmP+S1Uty3x4/
XyX2uhsViFQ9w5gLLBUOjiycbFyejgK3UymRoD2ye0qzSVG5tTejp4Rv3296jQxf
mQphoxdiqujqlG41gSNejYbu6vIfVCtBmmBojr1y3jb1NidDzYGYScfVZgFUWVXc
FvkRyxdKCyViTFpqKwPTdezjMek33kxgmASP1FG5mk4I1dWQ35Y5tLZshvYnGzlY
7Ec41aq5K3W+sk4xSKRlVb6Ac037dU4mnEl4eN3xg+tIykHehXn85CzoiHJIkQ1z
y0BsZtfJYlKswdfmd1RKLNuin/I4AvtBlVEbRXnZUVj9BP3SejoYmVIy9Qs0Dc4b
pBW9j3gWXv+a0IpgSj3IHlUR9piPykOoD70oFQb59kqdSeaOXHUA601l9Yu+rfUM
D4ybVrFqgTImF4sZATaUXufXjTl3p3jxcFUXZywpwds+26TcLj+XNkN9kfgWu6J/
EHptMDsevFuG1G94pMYkZ+/TtvAJuhqecxMUBPYia2rI2r2ZELC7PAF/xCszzleQ
pgK6dDGLxtK4FIKC53IC4jZXWIiV6UIPXef7q5pPahLAOGhSTIfwSadvKtXVBHSM
H38pzknw36QgTEhEWBdC2lKCoaP3xXjReYXQ6g1QkWhoKIuyDHImyCQS6xq0RYJC
ywONHLHX/QNEk5ng1nFEkDyAMCDU9F7bUGpokkGs0slb1nss8ue1zOOgwZqOsONh
uWFLTD132ttxdtSKUz8Xah6VnfX44bxrrXDou7RRxUToAZQW5AzbNU/4/QyYHb6n
CwxqJdxNLrnapNJn7/gBGaDF2QHtkWoLP5wdqjgpW3hZtBD/VgNY+m69MqnyePP9
Je2XaimOv03Zk+B83N3Q/qV7FA9XLG2G8/mzYk5nfrN4JKOydPjUxh/6bbQsRBqv
YxwvqLbfOKTfkh7qZgmg27evnXDr2372KrNosfmNgknFa5tLjZfBgFHZiCaaJmbg
rbLhQozLxfvvYqmy1NK9n0TR9GNFQZ47Js3zl/6mfWAOI1ZWInpHt6bXzNiYw/vv
6nJ6SgE2tE7kMpx2AjCs+r1JHxHskaBKLY9vjuo7WSOu1/Y2vyMEv4tcXnzAIYU7
G95XJ656IVS9cpFKftsyesa7KhE1K4MkBWD31f4firQRkiIbr0H0BO6s8MH4g79H
TDNajxVAXzojcs3f6HYsFN5EKDec9bId22aPLYTprzEpyr9aLmAPFEsg2iGdp9B9
ad2QzZM8OxaBHWfLIHA4jUotI/tqjv6c7vK8BxNcrpoNkisvNZhrX66t7S+TTuaD
q0E7iqpFpeJwdv5JSe7ohsTSpf3oA6vqaafUXfnc2kpmFgcFRyHD8U0sYjqTsZZA
PvETLEqvV2SUSbiq2UlrHUfub5fOGhGRjlu86QqnQz8h61Q3iAXFyY8MZXTxapII
o52KXhCCla5o8PMNZ8elTs/wPxTXulZpu5qnYmQzjxsyAnPmlYsxjYWadJ9OK3yU
YZ+ekns0QYbqgpqYKxIBWNL2R72py++/Fi0H2I7ofAJ8eolimEXkqrSdJZrI5v6W
p0YRnZWRxUYahbNLu1IB0PN3P0MVzVph1YCO1gCw81VfVpdQ4tpaiMT9I6EQuUo3
iyeK9MlVXw56ZW9KIm7DkJQ6B18Vbz4MtE6xpb6Sl8mInM4gn5yg7OwfBW6lk5iN
OUqaK58u8rz8qotCabfesT26IfNvqqLVSaJDkhJEyE1lovE3btwEIetSiAM6Upit
0ULJduolGxMS8OW0UG5h4ovukS4K+97DMMtvFnmyl6Yy4X4fEOBTShoacop8Lp0F
gbM2AF/IToQa5CXAfFSsEjOd6bLypMvMz1DHoxyJyE4/uK3xF4n6v/EWinWOSsHg
2a+/kIcukk/qvJdXhMBhMD4lyZ/tEfGrFyGvNp4BczaVZ27ZRaLcc1vJONUpaAxb
9KLhRQmm9Q/7hXaFoMbaHMHIUxBs6q4SvZaAYWEUbolYMxcxLaD2uEzNw5W11P+N
1sTBaWM2TdBmAclVa9ay796Ft2FuTI/k4pv5vExP2hRsXvQ189xbof0gPKkMQBjq
LUnMtOM704Vj6wH0MWUoVXWAsWbUqql3HFpXjBcQ3E18ZsfbUWHMlB8MYZ0rmk4v
BFuNRLxnLN9CufyJJYaRu3DY/gP28O78gy3N44Kh2QtiTKbZD47WegNJ1gK2jdYj
7nzcCOu4oTKIE0606xeoCpW88mVi23S3ys2NM8+6mKPxKMxyC1NSEkkBfjx7jJWW
VVNmwcUMKvkcNCgneMlivcIH8hBTskSnAKoDjBdhrsa61G9Pxu/plw3Cm82JqUSc
ehNsAk0kVkpAi4B8lnnRktTcjFrAp5jhpHWv5L3d8pj3J4N0HkKZqwi57XDYN5xw
WqvSyTDefY3uTNSiAcMUzaCbtnW3XFNir4Earuo2J/WOsXt8LmI8yExJy5ON4qUl
KOQhQ1GSppnP9cXKPNdJ0v91Hy6yf31ET/MI91MxSXJL8kTGVDQbnLEUu47XmZr1
pkvo/7CT7dpdXF/TjwIgvKRpgqWc7wzXcUj1cVyPiiW6ybFBkEhOR8sgG2IGZqVM
/rBNAFHkvB4jAJ97PQUJ5nj/6o1rFIIbVAgiCGRLexrlI1uKey4fIF63sFb3MtQD
SY2vFuvYou9YEhca9AjuH9EBXSaTh+qA33+pIGH4GEBxEL+9edH74BZ3QKQza7Kd
1fwFgMo0DogFf7kPRqmIxjydk/BTtUzu+e/u6Z2y6LI5DTL2fhNKOwhQR0IChhZ3
oDV4lNkgfZskVeoSZs/UvSNOoRIdywSVDyqRLvFID2ePFgbRjEWAsra7QQYSTUeM
K9BPqEfjD8RrbDvfFk66TuuhrdjNuDGi0BYa/iNMv2kmlpRHo18F3f7r5MIhclyI
GSScKvNu0EUGY0ZVTyX2gvOfafzradE1ee4kC4AOVDVwa1E9os42pWqFTCiSxMUq
B672aOMpPBVFZ1InY/hEo8zKyQbwWjLdbeFQ9jWEbI1hpYOGYmexwqbzop6qKeeB
yjkCMt4F1XZ5Sv2ycfdXgcaTuHjH/g8mQjgFEj5TXzBAPVRYS9wnCFKDgrVsXwyC
e+5cdSnUEoL5ByNpgPPX38QtjiBQJ1O9/9JToN4iiB5AvHhB+cN+F+LRmczVQ323
wQIYuLL7hokhXpRt7nhqtaNgI5/2GMVr79py0A7dQiA804q2Eimwxr5pDEkMwEWF
bkKE0xyxnfelQiBKsLuyIRImsopHEtMeKQykfzS7rh4MjcQ5WrgSzmvCdE7TRd21
0i5Elu+mPU2allDtPEpVYJ9BXnfllx7farrvXS/gAe0qSq+ld1N3HihZN0RdGARf
ggORDqzBJyvsqEdcuKYJy/F8y2+h3exR1wkK2yjBL7BFluwgcCeY+qc/1KOSmkIG
4gkxh6/lGUcLxFY+ZD17lOjXnwvzwDdmAzxNYwtdHi71TLIOjyYwha93usgR7E3a
YCu766D+KdlDW+zewdLCyFmKHtrrg5zsG8LtSjTZKu3lk5SEfduttmy91qRKuzR2
iRC//X8wuxpqRjpCE6xWeKRburI/LBRPXerRCV7W749nQn/cOjn6Cqvd8Az158SJ
V9mp5R/dS9zhWWdzo5raMGXtFhgdsNpMmLj5KIXpipfQb1E7iv5J3HK3XwdVOSYf
vKOq/Gxfxj0i+tPqYvmqXVY/fRk4qUUvlyZWwkrz3qhzKWSQfItPUjo8B2Er7qbA
AbspeQ29STciM0c2jIr8Y+Zr7EbLwvRt8SrH9bneBuKzDtpdmCqcOVL8vey6lm9L
CunGLkop/AbgiYKKh02qoqdEWIhnZ87cGNPQzqfndDN2PMW1db9EGoGxo6MxpT8S
zv/TVgxPdx8blZcsB86M+HpFx/n8x1ztYG8LdyiVX5TLdB+XqJD7RFN/qXmalUnY
mIKKNm2Zaz5bh0gkGd4yxnBvVlzD58WF9aZej0MFH1kMz78IIAEbxP+HKLQH/MJV
ZRUK0tUSWQs1W9hIoUkZ9/TcjZtLxSTGR7G0SfXtgSBl8mTgRZCRM2V9u98w1Jq2
K1fkzdNl3jaEOYvT5hEu/sqXSlEx3Kn+LUKynBM6GrjOyn73qF9qF2AcZ1VdZlHR
Gd25JpVq+ZTSzOzIT8DB+Lq6XftnQvX6H3Bm+JdKVdBzPmdTMJpzh2Pz0/6tq5Ev
tqwI+5iUHB95LLWXrk7wFGf3eWQobqbKbh1vzq57uYsub1Y/4m7mPqcOpY51q11c
db4pV/g1AQ0nPDK3P2J8j0nSb8QGzROe/1jFi++IBy+qEqnPAKBkbpdtKJ8ne5B4
9CSMKSxdeW21Idw9AXNSLVkvLQK6eNj9ehA8ejjDaMhCnlbEE6DmOzvcEXs2u263
OU0GUT/PAZovLIGDln70CK2G1gT9YvigPlY76GSkp9NqbsptVWdqpzwxxRZ42iby
ABCB4yleu1/KsO7iJPOzzan6gZptIdB66nuc1Vzj5fHGY2WCaoovDGBa4RlPjTBu
RZXW+GbBXeB+XIFjZnB6Gy7jQDNvbMcixvPOiZe2cXwecAqaJi8picYm6BX/+O1A
CnyDNPC3FBLsqDKySI0oECwc/ydeovOuJNW0iqcV6lNGJPqKIf26iYoK+E8Yvb5+
UQKFEkSuOkTpuDiT3konI6zxJtnGrcBDFBcsM20/OW1+NJISg3XUXWZO4hezMqx6
mXVPVLowXTL0v6TaZyds6gVryNYH7kZjiwKi02Z5KzR+XZ/1YcpayoJ8bGUSap10
Tb8SDPN831VK9AWC4qedO/dNuby5ngML105o+o0Ax4Eh1aAfGmxv6cpXtANeK9Le
VXegixBR6dk2dxa7LgWbyTQfhe9G8/jZMUNte+NDVBlzR1YWrEjseHziyj2nNg8k
kaNKGr9a5IxgyP9WeJlpTclc/jnvpBNELkDJsSLfwV5X/eeVkX29r4HqwS02qKVr
LiDh9is56B43euKiDUhzxXb8hJutFBJ7GW1xVa5YXUmQJNtzd1ZKVXQ+4peLd4o0
e3aiCf1lwQRIL/u3H/fZmnx/QvyaFQj9I2oeidMcJkEqWpvnsbuhFc2o2ZR8o7uF
N7UOOv74mektAaWMC09lUQwTKW05vsSMMmNm2ahLwANyhJUFhhAffBycgF2F39YP
05q6hNPPOMOb0Pd2xIV7DGsMLC2v/I1oWtqEihPzzi/bgAkUTZJ1/tYb9HR2Un9N
PY7Ng4/2P2B1n9c+0nyap6A+Ws6jFxrwT/3m0JouDXgRFbc/TzPIXGamNmsZKYNG
GyUzMujSYveVV43fICmAYhmW8aXi9NUD4wuQqOoO/XWcU+f0e154gd3LJcHak5Nc
aytZz8rKd7/YZumLq+NSVoquB+zn+EoFuZWlZtcn99lCPYcA+V9CkrYCLhewJ1Wu
tz84LDjDzLoPqcuPzaCtFfwskr+5cjPiiyjpUfUHC7xAYzyFFGvlkFb5UEXgihew
0e/469s6928h7HsRnFBtnxy/gl3oZCzjLxTyR+o7P8i1xNhyN4YCOns7jAmE1Sdv
BZ/O0PDT0/LRMz8S9WcBJMHjGBMZjR61Ja4Gcw8pkyGEky1b+8iJ+4ycMDLEo48T
Ef62QahEul16aD8B3IqAVJC+ziRKKv+F0G84aUF7bnmgVGSmkAGCCbriRIXxfENK
7zM/9r1N2lIjbw9HjzxKmaOmVcboW2EXBIWKwqm9Y6Zr1SHWRZSKpjAmgjdGNg9O
bfR6aS+UDmvMndJY0zfN7YKDtYFjy5+Q+gz6H0p1PYPRlVvEb/eg1rbXo/gJXoz+
+d85QDM7FsU52liROyeIBXeo8s0Ckr4P1wSf8saYcfN8hBvf3rvaCCW3++wSqvx5
dfhG62kW7FxmJk5d9GHfg5CwlePZDhmQXNH1c1+7RcBvBTs0rkM0qQIRvtE3pqN3
CFfMf14Q2UWGAJMcQcDCe4CU5PO4t6+Kpga9JBKEoMEcsCLVZTTy7if5mVxv+ZLw
1qIZ9ETACOvYbEoglB8dlWhLVECXwIHyVWbWz1dOGmRmwOB9SSiLRR14Tvh4gDY6
12HX+4aeA7652iAI8Mhg781r0A7pLoJq7zRL7yE70ageQ90OQ65gkoDLmeogcX8X
HcGnfSRRDeNZasoye7KBWr/NVJqfZymdcVcaO7ltRAHAk1Wldz6ywMYYifsWw+FN
+bdhVrmo2i1D2NtWyEZ4n1fcGrPH81Q/vtedrqS5ybDi0cLlBGp2si5NK35pvNTG
Vhz2GrmcZ0YsRgEJrSyr8JGEQDPgvMQy9/olUnRfN6RJyDJBOFbzJQIJUaeKaiyY
9wd9tWrZ9NnNPTqJm8Z2xvqmNCbsAs2K2BvH0AlTaZCeya7EqROlLQoaf5K3676v
lUcwLuqd5C7w6wymgN9ZP7T2u+XA+quU4VOKz0HSaVteFGaFw3zjQeUomAlFB71o
56FYNuZq2b5BRQx+3GSayAsqm3Cfm1Q2B+NyXb/nzALcU1hF5kb/3t+KGrRBCaZv
+b2yn7M8sGyfIfZ/JAWdsKGFSBFU5AHwX4QBoeLauxRbCRZLx2UKsHdGDJa8ddMU
Al5954SJua64pWRkDViWiNopinJEFD/8qNQZx/xnYHsTubiGt6laltFgapuy6z3O
+/iPGT6bLHROQZkI0PpGCPxHSbKXILBgHPLqZLx9S3PovINbsfKFTUbmzaDSjtAs
zwmUqZb9LMDnkOcQMVWmmDBgRw+k04miSHzAFO67xnGvSqcnj7TZJcqjTh1eKAmn
QHlcVdfr9QBvD3137a6RxdwpPdE9874kIzxyBkUhCHmivSqKPsUin5bHU91ZnMBd
ZiI7l3kFrmoNjA0QmV2D3ALtWQnWr9k1po+ewA+8CFfoiVNb9dFdEL57Ovbiy8KW
ISQGiqHF6Gcq7qd1v0EGmtdFQop+WXWgVchPqWol29FL+QRVE1/M7spGW4DgQJgv
Snqo5Mks3ytuQZFSMHb8coPjFGQd+vIFYVpnWFDGi3FFBubpePqUy3XYggJ1U9ZY
L5Ax3UDs3a6oqtzQ8nMJgfBqslFq+pxgENd5o3Y2AROQGXVpX2sOjNTpSCy4t+tG
e38Q/LUqGN+TMTXtQmhW70cE2G2LhKF8a/oD3KrLlcQxCHjT19o+d/zjPr+GPXoi
qbbgHBmAxZHK7qfQKBtf1PckgIp9a8wXnDRZXqdutz2KYBOtt14RwsiC+kVBfyb+
a9Ql9Qrx0FJ/qfNXsBySq5WGIYLb8FnZ/bFaL2CT+lalN9XzykLIcfNWE75zz89A
TWocxoKxt+zyRRrC+/DSbNua6L/to/et8HC4v5SPRMTUNrnWiflR9p7LCdAp9x3r
BJdx1Nv8xGyF4la0NJANOYjSnZjne5RAC5W5NTt2U4LAa9i6qiDjsOmhPbx8BXLZ
K2+KisjdBuFvnWlKBgh6sSUSOx9Ov7tg/9ZWvMGzxqbBe6j1xNn6MNXPM+Wko9yQ
eqCtagcnHZEN+bP20q2b1dpvM/m1rGgn/alqlqVTvltZBcJ3xoj6gt93hpq67uFP
f7HeM5iGL0BtqYAnxfC8hcSD2TI1vtNTjDP9bmb5c04imdpkhEizze9ODOdyh1rv
aEwyVnZnhWVHFoZVm3GIVnDEd6Fi91NTVb8ZhvhzcfHZwOL6zAdNYRyEhOcxzB+7
urJlfaW8RwLmubKKti+KMvJxomA4oetNzTe7B7nBAt/n7Pr7CaKuenzTvBm6NLdJ
LQ9Pq76HrLS1aoOfwWxpFU85p8DhvCd80Fk9y6xdyY1mg2G0r3UFeJPb+Mjzmm+q
wuEC4j2rnpVPoA7GgA3LszVpxw91U3kFyPjJU5HrtvYQKiyRC68NfX/ZNITwQSih
KOqh/gmtsyqcaI5CaGHfPDKaYuIBAIF07+i7r/1HP9IqsflNBiG/fsEOtqJgJUwe
V2IBDnCTN3S8DgrtRmTfzG/0ndnGRCAUv7y4ApKG4SoyvFRQAlIiA/3urToxA1zW
7m3CzMTvGCicn7FPN5FUHBStoms06gRT4Ef7WmyNtOTP7e3PlBBf5hji0fJ1GWOl
skO5/QaqjlEhrzkwCcEYztMHoU33nYCLdeUDCMRM3sP9r+eka1EtoOKNG28FPKpH
JzIv9nnuyGs7Cbn0RR7JWLSbwzuGo7K62Ad6dB1w+jeBkGGB8F3RYznQV/p6Ful9
m3hleaf39NX7gQ/SvxvtclGX6X6EzGdFtNzAoiq3WTHpTOojXRxR/BqXTtB3byzx
W1gpI/0x4C1IRlobQOAcXL/W3FZldWKq4OTUQyrpTEz9J+KjO+ENYwvpIGlaEipK
maJ5G22zJ4+8rW3f+RUns5EaVpXATThenxgprYMBjd6bnjE892jvb1wAkdGw8Uc/
Go03H68Ju0RkCnWJOXAjy5NkthXqitUEujI6F/0wNLZKSmBkcUpdTi19j9nMahMP
APwjWl8on0s4cPkXRctd8LzgXVNvZxnqJ1cihyKwjJH7SD12eHixG7XvDxogqFUP
eC0JN5EFvsBpXG5U1CI3GhUPUnhMDX0Qse8E2/pbnp80XdMsnA7BT4pD6pzKm09T
y7owBFuLli54yPk16ImVNRMyDlDnbGzuJ3zfYj/jm/VDyBC2undMRUD5yLIm9yDs
oJSJNrwaNTvJD+YzfXcU/uIRK1+ScQ90ngXal4ZikZGfBV22XG5gfzrZJFpbeJLx
H1gpnOlclqKOtKwbi+V2Ia8jZT0esexp05XzOMgkhhAz2rOgAO35xZsVfBIwHtoD
tNEIUhi8zdI2niobUZhztM5CTVueiDniZ3iXqppidjJHefEEs4/dseW7TO59XJ0m
zZZMHkg2gtyAz4Ne/IkcblT3RJRGc50cbe/7OXh49encS37mlGkxJnrpJkyRxJwk
oBFbFklcsVfv9BxHhFtXKWoDqZWdMkOrc88PjBJE5KVFxliJeMXhCloUQ8czfRrL
428qjpUhN+aUvTOSVi/ytUC6xwzHAFLt+Sncglua2ievavehWUqOZBJGRaVJMYdb
fNTxTvpfbD/5Hlv77XoXw6/PxzKujD5BRRO95rZekorjHBaI5QRrENYJQgPxcptW
PzWnFw+QTDeQIvmsuEjiPfRXmu0BZ7w2X5XL3obL4n4kKF7tEpRGlTftT+PT+lk/
U7CrGQKwsB2qVRQ/uxdsOh1Z/+ARM5uag9IImLHca0paXksHE4FU6GcPP58isBX/
VYhj9QdciNuA42CeChYLnz8FsokQj04vfzPs18ezcvqgQCC3VmHErAUq+ue5bMu0
FphM9U6gv0R8AJpP7jCWNcelNAsR0KQYsA+rMcp9J7WQIT3LNWo7Fj2Cem6d90WS
7GJhSTMd90Zl/3GrnbJx2zj2w34BWZPZEkt8zdQxwjjH+VK8Qjq4oaA1OfvVNpSp
OzD4kNVZMt5udSOqyF+tBktJ4CVhlfnLlB9GNSZtGHqXoYHdmsj+14JXyhViQTl2
zETxUODLXNvapVg8n3as6P68E3mzBwnZiCRgBTCmorFGKtgEp8echC7NMs34tXos
PVdLFZsAOodk85eEJvmC5nK+KuM/4WpkEPS3reFTBupnYfX7cn/5KzLIPh4KrQsE
xTstI9rr3sRY6NqrGdm6LJet32l90Eo7PgbvLUGRj3CNlUhJJCibv01KIjTYpV5L
9EqIz1TLSdrIjOdYAiuqwU5VQs0kyvQCjIp3TlN0AlNDg4L+8yKXz1NdPLikrmKJ
N3Eo+Je4BXaRSyldVami90YywrW8b016jfvhp/FdIl1flc0nQ6a5fzYyb5cm1wVr
oRmjV82D/MOsBzHigvZMVSjLgXmYTrjfHj4S2LdpzBE86tcEtcRA0ao+OaZZCceB
iQZENzlC3F8Z3ngoyGhUkkPVOnhTkiwszSKtVBAx3QAeLGI1zQC+pCPKtsALP9dk
oMR9iSiVm7Rccnyq3ifAX77giQ9TW9xSU6xaXuoTWc3gcvIACM2ugyrfgToASCVC
0sQz3O6gf1XTQH6kV9MEGtMu+huGVYxMKyuNadXSBukefUEvgaqnEoVL9BXb6XSG
4yM6DmIgoQeAt9+XdUkOEW+zzfSeLK2Is/kVUnO0ERnkUHV9ZK/2sjs8OhggktDV
4/rgfV8pUq7nUCPNgWF+4Ioffqe4kipw6h12QPCio0LfdHKbAsaptcKYvCksKbAz
pwh0Sn/FWjhTkGRSa2RBQaD9o5JzuBRhR+NtaUAxyt0JQaOKYXk/EOvfFIzrvgT2
4BZQs4aSL9X8AqVMIKXJiB6OCeJCFxs0Q1f2hbvjvZWf8h3C9oYJkqo/CEcl6TE2
H2Bpsv2s1rLpOJnZXQTYFkeIFe9++nm66LULpUxYtSUC9X8w1hp/mAWqkRveRXrw
IisvNPrs7nSu8540QspmRNLanMlD2m/0f9Ur9pW/xbPUF+W3bWzK9AELoaXDmkoU
vIQrwqikXORYtwDAToChpriWidsu3estKzksH4HLhZ3eisx2/6FjQlbtqM4asG/T
+Co8kJxl/TK3RcZMmZQc10/nmIZo6q1PbhHIthNpohzlsZG41zQPqM6dFjXKIQqy
jgOYCH9c6oAkuNIPb4qllG9WWlqOtyZN7IS++3a0m0941IrFRt72Bvd5hSjpMFdi
kT7Wd0WNgjyocq9y4tWJKWaMBRfp5xLEyFsbE6qGj4SB3r+S9FSrGltfmO8teiOG
icGIiwFIvl95a6gl9nccswLsexVTP7ZS3X3zs0xikuW1fWQXJDgZrfwSWiUF51yM
Vj2nyXKe2yxlKVETe5ReEjA4NG4VFBof7q/A6nDtB8Ny2RNgLXg/syYwmowRGzYM
Ec9wr7iM6B49SlzYFdDym5mzI7xz9IfbsUuiOI0bGMJokU3nMlskxJtNj0a/WQhg
OB39yjui/JpLzfAhwcXapywTZ4IVXvWhQuYcKWHBdg190n1oR7y8xKadv/2BBt77
uuGjQEe7iKNcXnydPPJtbBapLFyDwMKuELCxChQCS+SZRRDhguuoB8z2RUmMg3om
ZUYTxPN+DbJtANaBb7CE1PVrh9cx6Lydss5ZhuYuMh1H0MlzSP6NF+a/4vUqyLaE
AdBg318s0SBay6uCINJvCB7L7AOdpgn/kNoDBK7BaH47Xt+b5HMIg3F2NSZFR1WQ
AE8/55Z/Hf36vKsAmxDc+5Ju7/zqKBoXcdYLismt2yo31Imo3HRUsLzp63EhOwLl
P0Bi0+T8gSs0k24dwHUq6AxYqkqdrhOw75UmukjyQ/xm66BVNYgLTBiT6II34Z0T
bAD+XNK5TmcoKZct3MphIq47le43YGUnD1CWLwp0xZnP0B+OItdX5MvcG2NmoEXC
YREi7k0vHRHbqqtQu3thVSAq2TKdAGm+nfBif4nMiw5WTsscH6b+OaHVELI0levl
T5CU5Zx5Grh0wBhmu3n+OGc4pvX8l/+TqQVenLyZ5op5BcGG80RsgzlPbRveick8
+FyV6Ia3NcwY9lmS0QxXWRiJzkdlh3wW3NCTYpw3gLe/Zo0Jsz5pBIBby6XxqqsJ
exjI1n0+0iQpqt0QydAg+DxRalbyZ5OP5TvdMPcqTt5/aSeShdsW6yLGoVAGusuh
dNoZ752GO1OH1fNDh901kW14GqsksWAL5KGWHWwtMhKwEnhke6gbfNDX76JcC8fk
XCSUi5wbkXimVWKmDCUfwqdnsd1u5/kfN2azKuBWksoBQY4dH7yW6x/IFmtqoXyW
LfLmbwQA6Lepq9chI18dU5amseKeqhbEex3Fex+yC8CoD+o/9cDUALmDMw8Ui2X5
P5oRlwGCJ24zriN4oGFW1co+1pD4hfpZ72Qf7XvxIgV5nMOCrTmZHm8B9vFaT7xi
qyHvWC2127VSvxymO+LtOEQQXRhKnk3y9SJ4sWCOzmlNrcyXv09khahAAekDqYD8
YVgJsQ7t5K1T3FrafKxvAmTH66tLi6Ld9+idl9LEKHrAO7oZRdA4vcZ+1nUx0SO4
m+qKVkO5HsnTL8pqdXFZtfWGlMptvfq+6BNYZ2rZws8byyNWWdYRIDBHLMNJWN4+
jlwBojlVRv0Hvc3KbQF+o/wpawPh5zP+jUpH7NfYZ4Z1fqf2vB3L/bN/ih/BGVw8
GWLw5m0Ak1NmbSIkaptKUn/rgAy5/cbkWRWOz3BEEuowtZMYND2PZKTgKWs0018v
XNYYXRX3bEqKjFqJfLO5xnr8h4gImTiqRzFP6rYXZEzwdvT9vjBDdWwmdQwqbrHe
JPGaTndBx9q++smreLU8m9EBrm5krd3LyxYi3oNmCpvNU5x4O70T2XYV9yqP6IYu
ZeoW1jAk4InO8q6LIPjfs5GAf4HiAJUWruaTo9zDb4Iy+xZuIkM7RkJgT7Zp+C7U
oSW2sQ9eLtvbsjhCnuAj3FB/wETXyr/SaakPvJDY35o571ZxvbEKPqLu5ejnl1D9
9N4xzUmYsxG1WhZ3sDVQbhLQTMi/WO79lFhM2joCXp89yic5uVAmGMsnX7hf9Hoa
iZYJjUvioy3O7d27r95ZdA2eIMIzJSGEb3BunUQrDEudFoNadv2kBhW2Huaq84Fz
wIvapuxVrCEvptvf7QguhmAZifzvmDzxvxXxYW6smoaU2FtzaTZ6f+FFJ0banbz8
Doy5QAPckVBHuq+uiokY0JmX7WZofiwVTIVfO1Sgtkk2oxTldlppQdRg0neUbaRP
JU8mjyHsCcufjAVthurJCPBTuguv+sSoNgozC8hNzsY75bA/GJl8QA0fEbT4r+Cb
zMyCPUi1IS44mu1aTWzp3uSxVY7ae8ykOK6OXWTDgjmpWdeYaA8kctvBkak2XevL
ecU678UiXrhWs0dEVAF9NnKvWI7wUdSzugMYmk1QDOEqYz9/k2GT2s3hiUs8N6h7
Q9vxZ2klXO1ChoSwFNrsP20p8zNhoDfBn23fu/rvMKMqCRBYBsUNN28XfqoTKjKo
UMAuuQzgR/2j57mazy28vhj7A5oq2QAYLxJ38gtUA7BcOfMRHvduCKH3wp6fqi1Z
vGDH7zH3b914/JD0TNsyb4xGvuvbCOFbXzYT5eVJ57s06p165bHaBNyZMup7Fv44
d5O77+A0KQq+/rroQLhJ/5HvKX73WyzpLrqnI570WvyTcMp+B0+n07Dx2WAyk0Lw
OzHxCdRmfz8arHfQuZPZevCgtDtMRA/N/LTObgge/ulk6yNu6B/nUnReVDz8Z8Gn
95C2Z9F+srcHsJVakgbFzLK3q/SeLN8ZW+zyvCA1aLTwMK+TWoUTfTQm9OBLBqmj
TJXkL7bHMUEisW/FZzxZSyVLpOk2ndPu5T/c0pF2SceT9vlceD0dQVq0zTgMfUjD
8k81gZT9PqkJZ8xgIZIMXcAypIwjTVztAJDI26Vz4PYO4l5oAAKzNtaVz96Cd79F
LA+UbscMQtSISksNUGrE0VuEw14p0G3724I+uUKZdRQmRLfVbzrA0cJVT7vOQVdB
IdPco4i4ryWkF2ViRHbrZfRpD8469jc+huxfK2oaU+FkpZkvBa+mSjAghoudlK8S
4FBt8LxQCPGczhBYzL1hM1CjoRoQCcDk7AAa4NvWn82qARGnnCVOUJWlb4K8raea
b7YRGsd9aqrAyBQkVkKOr2WDxfJ8O9rUdGbo90vRMqFA2zHtKSM1pdUWwHvpRP8n
EdKNkrD5NRUKrLW7Rba2WkE+ajnsvL+3oLw2CgFiEUofSbai75qB2BXtKeI91JN1
bb85jYsml4CzbLahdjFwKJoR37w0uge8Mg9upj65v/ag3+DeSIL1RONw+rpNKfXl
5noBa9vyr5/IwAiSAmyHFKaEI7Z6BPeR/u10zn6MAzVYUhwwsJjBptNBnCIfPJHg
Wz3wBGJMJbxvYJBYMjdh9r8O/AI/oyplb8naVZmTxqax5HST8vxz8yyOACBTVDr7
ADA50SpN8ZNjd2eI4CkLyUfItqxvef576MFyUdheYQz9nhVvj9a2R4y5ETCksulY
thiRKlSGehSVvsWgmG8OOUxxJRmaOJW/26QnTxNaVIqJ+OlwLvwHUNau6++ZwYxU
dw0NR67L+5DDrbl5hlUuW45JEekNUv8nvblm9EumDH483Fxot95Rv+Gb9Gk8V+q9
a7+AkCFSSoufAETto2DuY8ham14eeoccSm+HWcnyh3Td2RYHKt13MtfAmoAX3mvS
qgbr8E/GpV8VB9z4qSxcUV2JcAAveO5nOB2/1zmQmOfoRNhtm5XbKvzg9z/pMKT/
6YejLkfiKB4z6TjOeDKjY53z7rDfAISwJMvVjNsRaa8I6DXk3OBJSN7gdrnFx6gA
zsbXjLVdiX94lj7/7TagSBjFyhiNrbBFqBe7WqrTIKVFqjbOs9a8hVUuj10ZclP2
CLrEpdCgOjnUppK8SKFYkiz9ab8+Vph6L9JKMQtvRbqqRHT2jH2aFuk2BrUl1Wmh
bhSTO0rjsWpnb79k36JAwmEaBiH35iGiVR5TTagAJsRanWcMSW6GXkACJ0fYf/Gj
CYyC3XbMNhYxgKgEvQKmyeqYPkkksaNCxIdOaBJtWmuUMHl1vuPCS92ZZs9Vyfm6
yEPsGsA4OzYSI6/+VNt+KKytlL3oSZoIzLdDa+hbWX5M7lFBHslCdVqWbOMqE+wE
jSQloaluN5zzfdGqRJiykAQbBZ3ZsMO5XAQRkKwz+HM6R6/I+mzStrGJ85bITKRa
lQZYBoFU+X+ATnslRfsQmkclCEFo6oWWGNXINkT6vUbNTpjQKgsXI1Sry+wwFzz7
2+DqGBp+LcnvfB1ArloVC+K4E/hUUDvssUWPbiepNsSTRJQSMniacM666v3MX13l
ULKrHUABnC0kWACu6geDj3uZvYnjdNABsJXWfvNb0o8S4rXh9l/rZLAh1208x6Qf
CKvIeOt+eoH5i8b2oag/Pf+0a0NGkh4mA/WZzRnbtc7P3bQlMPxOLYK6iiKR+XHP
u7mLkIEyM93nSY5D/t99y7bT/2DE85fkr2n4ax4OV8KgdTyIyCWItRiEZLselyOu
pO/uf0mEBqyWdH5RfCwLO/2HeovCYczJC/OVmnkTdZIPv3H3mYpbvWd/HSNzQshE
pT7pbPtjeSgLZreJ0qTXtlDzNT9u3YBKW6koOSl7knW3qVG9BGblVgaRNGuNlgIy
VKCiiZbE/GluY7AemKW8gBSJrVJPc6Rs5LIl8vsXHbn9rDeFRY8EhyIFYwy68I3J
3dJx25iWeqNr9Z9Vy8ai0JZ/RBlr5R+iHbhAeHPcY9rVp5NSRnYnCtHB/GP6JclC
lv5GHcJqNOq+C+5SiDDN88y698HRTrGOBtBmJ2/lauKIlfOrUMNz3dECElr5Jb/Z
KjCdbGo6kwYWOf0TGa2GD7uz9fkBOO+Ldn+2gog5Ele9qZUiI0Npl4PDWWrgQjKj
Cwxv8utxl5uGKP3BrN75Zjl0fh7uWlVKousjyviMqER3jZ0hyPYdtKA2/gL7E1Lv
4Q4UQka3lnsindgC/ypW6XK4ox/H2wvbIcBvMh7+YJ1b+JPf2rjgFuirsTZsdZ39
x5u3n97IRHNu7KJA72vUc28XWDZLM2hOnkD1LhUk5UxzMlQh/5unwfWdHCebpCHR
xmOWeYrKXydTk2BXvzDI/7XDlDnZoEibxklDTOiYO56c1BzaIjvn9uj8t3P4w6ov
ZTAsK9wSzjH8IWoHR3nq3kVXkO1X5M4r0cZOUCYsNRB2By6x8GXv2L0ZDAvULDlt
jqUPc82dtdymmiWSmm1khkV6fgxlgl5uDeWItNBAKS6TXSOIqLupquwwxVkzQWoh
OCJg60CsLhjg3bIzL2tI9ghB6IqBBLQGhVHy8AKbeJsQxHlQNy7mj5gwzmIRfrZN
d6bEZbMfoG6wsIGsyVe9CLvuwYzLFo8NF5HR9vgBAZgwn3haGzR9asPIJAUgkA3K
lFTVYA0RRXQxZvCt9WBoaWClE7KceaKjWZETNyTEKyxmNSAiS7n5kJYwVxSiAYVU
fxoHDlXobI8Ng3Wve+mWujzw6adJPLLSjYha8wdSTkYfgoeXuzecCRbff6fLyxZD
d/UzxQ0NXIP5YgT6pn7kwz8IBQv4GDuB8kVAVP5EnmMCDA5iuEqO8FMs7qUQiFZv
kgh5x6/unwvCGWZiOWwVrgGqsDAXJIyaB/YUmn1PjBix93wCpLbWnRYPI4D3ckYH
IhnTeEqFtbFCGlU1TfcMY225dZ63Hmr+WhIPpAJik7y/m5jHnLwCJ7ko6AXBWdze
qmiloxW+Fw971u0LGhzNLDhOYf+4iFJTFyVXd27S9kLpZ7DbKNdMzti5uSGhCg8Q
H/8pcN4k5DFpyQ5uDpy4mPT3sQz6c5pSoW9KGtkKPY9/8BhtuBPrfg/um2BQqUAl
tTB69t634/zgdnByiY2CHAOT87Cr+/hILW70v840/o42mm33znVIt1jV8YmasYMs
kF7fDebUb5BEPh4ABi6BUJpnlLKJdiS6DiBdYFBJ8CY0Baq86S+JzOjPODPmUaEV
H02qlgVgGO1gZiTEleHe+VdmyVbsd3q2seZmf9hFXX0vCGpZ3ZhZ4GZ+60In0P/7
1Z+/lzObd8ixZYPCvdNFwiMHAgbkOJLbEnRoJaeLJlM1LBKHODSQxD5dnX8xniXV
Eumc1QJGxWyVp7f/qrZ3txiCLbGvlbeudLDDLGpa85K3q67tZGgfkJ6vi50J4kwN
rd4sOUUcdt0dhhNQ6UWf7Pk3ubpGj90eSJEHdn+2XXBLWTWhsPaHxS7tX5WEPTrg
66lrU7GyfU7XtzUqgqDKTY0a71MSj1z1qVk68Po+jG9Z5LlI+RPlR/iXF3xa6j5V
SrpxEMlAr6tlsGjbQVRhaG+XBqmU7vwi75L650pAyLU/dF6oR6idRQ9Le+BRXM/W
fNB2ihFV3W56K0mHhPZBJUyK6gr4oHkrGfgxqWPXQ7tmMP9foYQ9iFFrNlx/zbmh
4eNWS7oiavWbK9ui60SHp9hvcspVyJwpNx/wewbIFo8pfofMLox0PI7Qf4HXdj/t
C+0xcy5DlodmH8/XMayqC7SNnTkrcnSk2K/US7Nj38GF3sfxY1b/5DXUc8uvMn9r
VVO/A5OJ+N3s4IdzZKsu9zp40zS9mUuH9FnCdH3h1c1R0fSaJnM46yC3mkOsP0Lo
IE39E753EsHgzk5DUhF6lw69Bgp/FdDks0QjKIxuH6X1zZdmKVjn2NmPJIqoIXHM
iA88kr3f/omU3faJnJPdQX6bK4ht2ngNV4SWstlOpfhtRkwCzu/XXXZt44S8Y+MB
JLR+RnSGuP944bY85INVVP9rtUxEms+6vnloPaRTQkEOEVDTz2vjUVKx8cN+D/G4
ckXgltjup+400TwoMR0ksm7gAxycYzg20EV3NoWSQA2CKq/rXLDuNFsqbb+NE7pL
ra9FAGXkUrwEw1z6HqTUuoxrKIqClvJjixXS/zlHWRgNop0kk72/ODJCsKjBc8Sz
OS1oxj2yk/qMgrUlVP8dq+mSusB+rR/zo/0s5RvjpsPmvAHsUhHp1I9NkzFng855
LhmpGoprJkBCX329C9hRGm3hz/l4DPIWJ/S4Zi8tfyQPaU/qUvTv92064yZMUU7P
Rm0WpNWxNza5FbgJ7mU0PeGmN9WDgQruplXyuex1sRc9VnjtVXH4u135YkFSJkNL
ePLhRNP4cKadY1GXdkQcNE7FPc6PdAJIZ/h2f6ICT+P6LEcijszqZE9sloDkJKcc
FHHsGsHZUcBjpWHqT0eLMuKwt++uAeAkyo1bbu0GEmMYEzZyKWUjDges2ObVfJco
SbcsRBtiXYgG/vD4Vhz5FLUX815afpe9f7R+ZO6xBzL7LyX4SgF6YyWhqbqUtxLo
zUhCg8Me7/aYyi6bRNzAWdjvB3oK0HJfL9CuT/YTeVgGkryLgEx+H7g7BHuitH77
6iS5N0RXrxpwXVM/f3rU9z4vxZmmGE3kXQ760T7ImlySVTTBy4WXao/VDEUTOytg
p+KnMgt+Q4XSgjSb8tcgodQJ2muu703wIJUaUpOU+4Cuk2CQhQc3J738rWxaATmk
m0XYQwhVQ6vR33PHyr6X4znMe1aCi6jMJ2+YztPT6Ah3aJDOx+jI1zXHHZaYQc0U
KdtDugaJi2UAtj87Tk0n1ajBoW/tJ7Q15rq2fT1xRY2R95ZRWUdXB8qqrK0NWGND
s3RcioWTWroRRc6UpF+C3iQhYyxwLvEc0PLqoqmcpwx2k1vp/t6uFvXvLe29sPYZ
PjI8ANA4WPdrF5a5tflGWsmGLL23Qypm92XHboj1vpcXi0cW+hbojwoTj9f0QMl5
JyVjqW84J7QKsilMwz08IQbtu0/U/6LRPfIcZTcFU3JccJNnBbaXeSIlmcOdguVn
cOAVxMWqwlo978DR0IlmL0E5T6iIjHbwhU44/I+APwoxJV/nME26SCXlpC/7/Nio
ZE4wZJyKzq1g+OJy+o+v8k3QYF2CflkeBX4ERV1es0pocxGpJFWJjv/Z9pLPVbp1
RySRRnUyoUfejL83K7iR0PFUkYvlIHyO9iTLjl5ptvH9X91Ie2WuTis6GbdzSu7u
a7yc5tdJqmzZDJdgpZv8ljQol6/i/McyLKnZy+JbUazzHTVeDjl4CZz8cSzZn84c
sRBP4cJ4VE4oxJfXfMcmgGXfCT3ekn36EEp0cb8muBBCM90StTx792A0R0EHEKh7
IuSLlf8FrDbFrYKejESWqOVoBD685Yt0QNoQ1j5PmKMS/S7Me5QhONgss5S+Auqv
DDp5IlO+IJfe45jHJr/rdRhIeNK9EB9wXETs4h8iK3SrxxjP7+4qoB2dI1dlub0v
UzX1rjgAFQKi/kXmy+rd/7CQXieTBidAL50opJUbWiRFEAJ/kerZkL4B5LxebSla
Z+HqCUFrniS4+ATvbTmqBLaOIj08rIMDtjaHfYPX02YYCaaxZ/TzkzIWl+5a9nlz
8GXi9V6nkNFz7TgN+2YXosgvRE5ADj3/UEryl0aftxsv35IrVNXNcG2KN8EQW0/r
LX901YobsZEMA7C5J6pAQAqkBtrOKjnwUq248PsnX5B0Q5AL8qXkl2zfh1ePD5pE
BtxKfg0sjILqyE1GoU24zbW90BCB5qDZQQjuwNmBR/vvH2OolvbFBTVL/wvgjL0K
zmomWQhFMp1kmS2lrZ1PbY9LGXS8zWv+rSD64Qz9MjUEN0y/o9j84/HtMkUE+HU2
WcPSuZcegpWrUjlF3tU0cU7TK3LsiOVM9kOcp5cNrqpNoIOx/3tmnf7hr0iph51I
tbvsMXS1TqCLOpLaJ2XeVMcVAZy2woUlPtM/nP/F4kTv6eVZqLZUWzMmDC2X/QI2
emUlDgru5NItJxHVSiNEgpPahEG1zxjHl/QsI12VSBb1oAR4DKth1A3HKFaKCQhc
bltBm4mzNcBOtQ2V3z4w1blBqPpY7rIlkRpQyGE9XFfkOp/UkmMW2RpQLlN8vFSi
+JU/T8L1pVHxBe2k1jSbsNFjGNvzLLzIkHlkHpQVbY1lJaSCJm9S4zaGRYGHSwMS
IrKP+QOosAXKFBCrBKxqmQI6PNOvnKsgRAZp6Rd+8HZSrsDY9udqFaV9L6eiYMwF
iiMu30QwcE7Z9FMnGd76KUQ3kWVCeE//BqW859iZ9572aQBGP1kmWUX0dydvRNBJ
0iQdGx91rL9Gm1DWb0MObU8rYBroqVnV0lGVLlgurAx3B9eal7M4PBorPyUHN4ni
KpvRa7dgyOTVeXI2+kCZAQrRHc17wS5tGonf8fofkdX87c8NcPbkL3uQkyLYaff8
uQgGnh7/Sc1MDXriQphHKkUb8KHFWGjp658vX4JK828jq8zvS4z6h9tEPMXswJO8
YCpZmdMMEsbGXAwgyujgoBu2YQaAQeBlkhgrDoH1FKv8yAuJ7yMB51w+LbszVVvS
RacRH5Mof5W3eladJ5ctTI7CbdbPvcin2IlU1wLrQwrBJIUum1HWBavcMy2HrcJv
Pjg5Fq8cFspFHtcJobDMoGuXMWfo/+M/51kNEreKbktwRU3dtHpringr4dIQ3HWI
dT3Ul5h6yqUmN0OvFP4+9/X63jRVwUXnL3bwBjHN/RHMxH853B1HsSP0VCPTZPe5
6cDqhBILjyC+R5kp3iGQlOxABBhmLRoFCwGctjAgs8qCRuwYmElXRt+RqnLTMEiI
A3PlNEdicSmsefhx6lBNtySDSfgVwhoWu9TB9f9JrhUMMJiGjVMSD0OV3vuWEPQK
/ct9usjle2ydVqMi0juL9xswWGJ5wwKzt4K38Zo4aIWvNKELVAWZPFwyk7ANM7Oc
X2TR+L3GZV7BxTkjd6htOrgfAWIY7G8LcXkeUEUZEaf4qx4kxrKU1d/25wTUgs7d
08S0ylNrgvf9EiB++0sUZX5RLPurGBUqV/sXkud2Q3xfxMuIRVLEkgbsZwh3Wm02
9TeZp/vW/efKeEb2gzUu9j1Y4XVwSRi5j0LOdG0ZnXTYGp48iJDOvGUdMB8wX/Sq
D/p3CodcmlvnCsTwJ2kmVXCmTdGr6wgHiGMa3rbJulueX+WQMpcDWSWmIvs77zuV
D7JWiAwrE9OSrd5t6V1JW6rlWtcxLM6TSCwzUJLJFwwD1Uz+HCPcaNGFkQT3tZCh
X7AjadWk2xx2LQxEMPHzAJ4Ii3Y/zDSIFY3TOy1MIqb0lYeSdpmtC2pnKdq+UDwq
v0F1W4wPbe3YcVEJ009xD9+08tFLQHVRscpvxCDhAmdRjMlAaZfCspw1cwwg9B7R
Ns+QPCHUiPZEA660Q1cnYF+PZwyn/ZNYcuEvVlJmaHv0cr+7Ub/zi5xhXdIXC0LJ
zvE7zwlnKnJ3Oo+jk8kE+tf5QTwdmip1hHbwa6lL3p+XLcHWS2mRlDYSdEiU9G+E
X04CZRZfL0bN9vXy/JPu/ga29FdCwHztri0wEvp5kD7kuIDs0MnNHYY7xP+rUnUE
CrxLZUB5QiS+JuS5F8s3eC6Xobzg1xj9ttNZkKfXfh/3wjBR2E2cKDCze73Sg7LE
/2FUFiNHfz7FFomNjtUifV73jCh0J+zIE9sJK50ZnaR21xrcj+vtUUJ7Qponn3nC
hNAuPT1ktEwT91CH/SpRwXsCtedT87dFTblPV3sbCYzzfa+VNqUbKjcmYvF4XNvJ
diALG+UvO8df6224JphtLq5oot5rYvMGfo5l4m1g5LyamXOJE/wWZbkaNgvan9kq
MOTAIws0hKfQkXVsfNPMIXm4q1nJeNnruhWtSLOhUtFxuuHBN6ckAh3Uvxc/llGD
YJ57zpzIXmQ1gp8OxporfXJ2z6uayKvvo8bXRa4ZeIfdBKPZxBDpBAvmAc7pNMk4
1rFlV5ZHhj6Z5Xca9iVx1Hck1RWYXsKS7bOndpL+Ir0cb2ipSoJqtpuukVFcQMuH
QS2sgECf9/dmGxm/gxTIusR5sMeJDzwXYNdpaJtr22ryqIRop+/AlhOi6RO4/dxk
tj0IPaWHwVgCSTDF9N5p+hxzMzfxPlGbChQCZtkOH0TXRvZXw/BpgMB7XlKzsPjl
XYYPEyKrisqqps+u+pT1ZirYcAFdqn/IYjWZ6sTIv2cW/XZxoGcj9Rx/OuUMpzv7
UkPeP1ow612XUvUVTS67JDjmk37luTHWPL6YBOXqbmOuE51bchEoTH3MjnQEgyu4
giJYUYIfIuXmMixZLmScnyEdiupGrjQi9UrWhAuauZUKjGrBkEiSNO053Jicp4Jd
U/6QLI2x5AkzgaZCcGm2SM2Dv9VQH0ShQkq3hmrds5BHNOS+nuIgKbnP2bMNgtgw
SUsczD1xf5YFd8ARY9gzJ+EVJSErSpqP8iEivYWgSJ8lzCJvxrZbgXpKeKhcfz5X
jpbxvH19jG4usR5nBJn+i0XCMYvlYvfuVG0nBn2B14Vm+EiBIqPSqzZ3oKyZJQVl
TTkU3ab2djf+rBwl1m5vMBdrtgD+8fUP3TMQ/iTTO8X59Barusnh4hCY+mvaQMD2
g4zsCeiinMjhLgUnwKo1Ry0XpS0QxvlHV5+bAt/k277I0924vcYezsADQJ04mhkq
tF6z6Sgy8zTPnG7zYzhJLGfM7TP3MhKDHot1XhWs86JIMLM5ApWYDKoMmDV2oonK
38EtuAalyXAzJUu6AMATIry/q17u6hGJZoQXZtE6HdlWpUJ/NCzlDhMECwyVD3ZB
cgjWhQ0PT+WuBTucVOR8nGIoQMS8z+c7nrCc82vof16DaRxH+2yG+4/MIhpyy3k6
BiS9W4yb7XT9r/AsB3bAE0zShFDGW99Jg5Y0UFHjHEx/ezdireVmTtGw2p3X/tEy
LWVgxSHaWf/DVS7EBowkIzXky9BJWs8inTHcGt6MRUMvLmJNSQKzE9JCDS926GTD
Z5ADTBrLnReFbs01BngS+WSp5jYznqtxNE+KrtImEK3HrhBHwSP3Unsfo+Acd7yn
24eXN+atKykGe8oXccZIK0/o9bTSERIpWSJaGyEN4l5Y83hcklsbG30s1zCgJQiZ
6YmPssCGeFOU/Xp+iR8lzTprWYsSOza9VBeTo4e3EU92ya+9lZHp45dKKiXplELO
9eB1D233hAs9YcyRS0ppWPHeHyDCRr9qvQSfsSWnb1fZ8TsI/7kjGjFnf57K6AZU
rNnWy0XtzlfKzEdAuVh5/5/qKBpFlsfV0NK62y618J0cst+LLUfIFPVGEVoodH44
DwGcmED0SVOGkadXBXqordudKRxbzar8JcfdJ8IP1tMaiICDwkZN7MOjAo2tP6Ep
aPL23nApK0hMsr2AO7Rty8BCR88mbQxlhK0/2YrQiMgvYS7yY+NqN/Wa7pABWO1I
OCIcBREeU/s59nxPBXoeswNCr65+RouOer5d5EAFod84jCz6smvUHGZELcK2Bzwj
TiHmcbZW02v/hAVFzynmfmu3gU1Lmjj3r2lSntpAdp6lVJ216SnPxJO7eFAqxa0L
gPpdn4bhxu1okX6AfFgLnHMl5tjW+UBrwbXeMzHTi6kq6Ey+7LjujEjFsBvPwb5l
QCBBRdPdkWWGKoxQtal1Tp/5KDLwqgF9jGiPMRYX2oyVLHM1zmFeQBk3Gz2NxXqY
PXZOAUWIZirO1PHMJlxxhFYa4zjuQmd1EDMvycs1z/vC/KztrqmID/8yEbyJapRR
suBTpWUGPqDnhP+GCTCr0GU0UZkgsxCSVtEHGxfsy+LUgUOkm40W4sehLr0O1d38
1/HixA1V2e7GD93gKQ8lYRfmh6pP97zl5u5z7WLHVwuykeo/nMar2hxOJS7SFAYl
BliV2rvtgwPszx9qg9Scak/8QW+w8RCao/IZ6RD1ubBNbUefxmz+VGvhn32djQ/j
mZPtF6DtVkYRVvBnIVbfC2F8iVkUqnYgrAMy8Olk9EgtKK785Wk3JQgLWYomrx54
CjFGnQz2EM3RdMNH08K5asy9nn52t2BgczT6TMOiQajmErOrOlP3+LW4ieHnzmDv
kOOzxHO0ovj9dQCS3/X7ZT+U+MVI4BkXo9Mh5C8kJupwjVw7e+OquliZXc/YhmT1
9zfvKE7ejJbClmCGDm2oiffg0zyzD2GSDqdPuIgfZeDfgRA0CNsOJpi1O0rP7LYT
JIMYgarrqCIdt3FanK8rTkHWoz8/jjVWc+kbyZqlUQbE3hjgoelbtgNcniIWPLoA
8dG95HQfvGL4M7ZbKJw3g5Hlomh+SjtvVcB7effO+twqTv5filE3Zjd6PZNvm2UX
tB6i3JClnHqHBZvIR51piZm0ycR7BsnWklXpsZWn3u8KCASWbU4RY2eT31SGHjxY
lBGkWE6BQMn1re4gugBTYIL1xXJHy3VxqsP3ks9y/7fI63eGirHb/2l+fbFyFIZC
MtmDuouvGMhXqC3JHy6XLNF/ljoGLwSJEOWVW+Bh8snSJmjjq3SeQKgrBvA++Fv4
eEshVWyETJw+/d3FWyyVkAX7ISBGeRJEN6zdzYNRqEjSkxe1PiN9MOsrEdxbjtdG
eaGgZE9Dsi8Xb58uVlWeSlyO6v1OFRVQW6GPy6Q8SSoH9jnOT3FDqkia4tQO/t4Z
OkuewDyxOla6u33Huhb9p7X137xAk/urDhLlm0SODxdWOvLH8TG8acsj+WBwpmRM
00LFlu2EySvpxyjQR+V1g4ujd1TVMB8YVI+W1+TZ5kNYQNzckLErUcVnNKTxcgK1
G246gIjuEBhTOLr3/GSB6J0al92cZzh5ao3Wx07KhxCfGUpw72SxfYbS7VuHRPhR
3omHwWmiTrW5UXcyL3YoNeIQlr7z8836nimVifOeZB5yOHJr4yp9crkJoKC4rdV8
TH4JU9fYjQ0j4/hEuCFNClG2PML1kn8ASYR5NYzq+37OcZbHCgztxB/R5KlqXiBp
GlftfANt34EtCroISpmBkTctYqrfBE+nvNfm/rV9lBmT5HY9Sj2usGlq6Qc6FIDW
IdMLx3AJPthC5L+e+BDCn+4U5ykz4fYMi4SGzdFif4QM+hCuM1fzJFix2AxuON2y
n9YFQ/u0082q6eNIt6kT5LaD5n/G1VseciC9JVJCO36s8hi3eVlWJYiEYwbkPimP
T7tKusFL5C2rDHKUNiXury8gfmtKerc4s7k6mASBIb1c2hjhnsZhH6MzAwQ6Qkw1
oirKaWyppVxbi91bz4Z8uKQrpXLKeRXRLeU+Jrf12RmCoXNTAZB4FBla994Evz2L
tevBRUSKUVEr9Bo53Xw8cJ92z4A1sI1VKiYWkyP47RrpShPs14KEIrnG4loDglqR
Y1NTiv7elclJFTcDVkBZBv4m6Pq2OEr23ePDEnWCEu70FjIupkFoHPoId2qfvFjL
sBzOeFz5xniz+mqcpjJlWzIQ8aN8KuE2N/XresgpMqHnkjQxPBkknRYngmiMtXbC
+KBWNmi3M6c3OjGHnHuXuZClu70Jg9uXRSy4zLGnlGWDiorXRs/lhiYuUz3RP9MR
0MIcAnyuIWiH8Kp07xgseYwNqV7C5Is9zhyaP8pYWVcarh01PASn9UA/kOSnQCXA
XR17pEXTaqt6zuBj5G4hcTDNFpEBlLrwGjN3C/XxoO1HDVKYtH+FJD4dvlHPcTiJ
UEfoCAq7EUv9c7TFg0MQm+oG3JjftKNUt/AIcqlRnIDFNyc8AgK3FiDlYVr54DL1
spJ2yEyZMhWQhj8kyPUjgGBdzhrqNRQM3bWRRwekGZbWPmWTGSXO7oEWZPBAwazn
NGd+VwR648FB5Xb9jau/nw6Pl6WcAJ1UpFHi9W3BvSX28KN3MK4pzw/vXYgwmNfH
cHxF3qNyUxN6Mx29KQuT8mLG5ZYXjqIw4AeS0RxfIhWY0W7ejolsB5JYfYKh9SmM
K0FPFuehfWm8Ia8Aam4jJMwxLINerFxLyb6Tx8NzjMxr0zevqqUUAUsGdRlrsNUl
BL+Z37siTG0VvbdpaQXg1ye7hwd1CLEYJiFIDktjZsNj1yBIIOej3KSxGCh83wE/
BhuWFBa/eYaIPe8svWqxOAkrDkRqCKaKv6+1+TDbHyR13+Dlaa8HTIxBxYliMjsP
8D8IH5LE7Hht2eY1zHZPQDqlmWDgDpkv/9WQrqJGDcWpwqiKL8WfEGTkVvQ5Vhrm
g01tWzeU3L7BwLLFXPbrv8HztW+XHy/OtzkiphloBnvrmSL31ZF1ztGUeCRB7egt
zsgS6bIVDAxelZ6eU7TXyoqSBy8T/7lrwQE/2kE2V+ih47TNvylXy02oS75Z4NPq
CZloxh+64cMk1v5TjhKr7kKKDJd0r2uDPqCjQPNbly3kXsPGYlQxAy4LbzpKGiUO
4TDbbtqZZ+YQZdVKMPzartUFAQouFUU71V5/5wjM+/c6KYLf6J+yaEqmm1fcKjBj
2f83rEJoO85g9qj7lrecx75GWJSW2+WTRmZTgdMZbgT8WU9SfUdQ/f+hsgN6wGGK
R4Y4L2gHfu35c6BGIppQFfbdan4F+EKpYf37AiiHQI2a1BLND4Zw3FglvWnopnjG
yghQdt9C6U/F27dpw9byvqIwCVnhAoO/nr8V73Uo4u9gkeaiJ4HwEsXphuk7OWRT
gzPbEsZLT9kQ8i78vZop3SmzgeAW2GG+UjELkpK+14NfosWoCGZal4M6tBDxTWmS
Ix0GKt+RP6G/T9l3FwRwuN4xKJhPS6zwtnlK67E5ztgjopIgNu5sPBR0sLipfW5J
zBlBIg5SPi82klQEeJSt7jaLPqnizllkT3wC0whzyHapSR6zJvjV3+3PIDxiiaTu
SbV3wiXd8bYLDjIeiD41g9CtcxjzBLnDogFvsaoDgk5Oh9wnSPjCjy9W4rdZ0yur
os1Tl2eMUGTEmdfgfGmQxFSQX9yruSQoInhTEiGQUTbblLWQ0kX2fS0fDrPa20Eh
k55/erJipXhrFL9AfmNbEmfYw+g3YJemmZIU6hc7zLN8YtDdlRzq1lyeEVWBuXnr
PbQPjh/Zt6+2Trb0l2KhmwK5leC4cx0GAJ//i+7ux1lK5m90S6US37o+Yy0Hldtt
D/VKqHpyiWJh2fhenaPJcZL/EZaG6MKNultjpE/0N3jaGhv3+BmZnffMF9st00KQ
ibRvT27cz8kdnJxUPsUocfAA3rY423NBipNV+5cH8eHpjltD7hgsJfzw0vpqaC9l
xua/ElNns48NHy9M91Ws0Q5Jl6SYavtFYchAwiEyWntWILYdFbjkLHffa1doMgv6
UZRxbeNWG3VmBenenIOLhDfVx9sYAwEOaqADHQgbpNp9F56VhrgY6cdH9MPggvO7
cRR82iAuFWYnCPL3zbewbNtTWFQThrGIyVcp9pL1qsmEw6WUEfePgyALx8aqWP3S
0LGPL902QhYFC4ziK7JA136rJMWX3KmMSQiVgf4o7OIO5kjvQr0PdOdE58AKOmqi
GDkkZwkNMuCvM/aVpfs0CoRwYjIxS+5EdBNfvy2KVA+xb6S8Je51LK3J5HbkYNoK
qii26ddQkxLhudJAeY7lkoHivyJJ6XaBHZ0thmIw2g83dGEo2bwKaDe4BV6F+yj5
qerS7/a4KdK6EJHFomvOUj1zIBR8KJAYEHyUxzqyga9VoPrx4LIqeRaFtKaeFIT9
mRX9xkSfQHnMw1hf3t+63HVAYnBVhoP9oDNXvRssxNrEvAwBdOV50N79fY8RY5Zj
8s0DI3A2DN70TFQqXiBpzWwMQveQAy4jm0IH95/qsXD43trvS8UitYIHAcjsk6qg
q/kTgqk7KOq+Y4qLM1u2jNeWHxD6/UGnImQk22zHUtcNLM+PawyfXUONS8TFg/3K
uD1lRPsXMcYK2LfScy9VFB7NDe6XuBjgiMZjCQewLyZKQxH2b3JoBf/pvcjqXFip
uXLYTxm1KcciTIi6PSGhQlcDsctS0CEidC51/tb54xaoLa+GonzhBgwod/2vN1UF
BN1lJdynlzDq+SJ8EOUF5MK+8r0/r985a8OrKndJNW799hW/11DLJZNYAzILh06d
O5P48FKLbN0kwkjhbB9IHDeXuSU8Vdz2E2X4J6Q+KWGqnMlXgMWpzVTQ5qIYrr8E
HjK7B0eJ2YJOGtkXo5AXI/V9Ok5zvqhmZy3yjY1P8oDxFxfGAoQ7aojtLCm7KlOI
jk7/pP8gpmWHy9gDO0TyYyLx0qQn3le76qR1zKY2Lpon5pxDCr3r8tOtwPKtPpqs
ZSOD2//Wfm352e0j6chJXBgzT4667u5cBBtArlSNlrDnlsp5TJCLXouhDoGAavCz
vIbFMYdzGdiQSlBUrguX+SFel6C+FhoQMikl9oUVlRHeGsDKMJxJS3Juy3BqCrGg
+nbRU3oZtvS+gUfZOcya91owLxRw0Ip94UP0yktphyshK+vj7v2LO67yuvG6ClcV
eNNdnE/zbg1dXulnFowbOGgOuEhn/f6NtAcBKmZ7U3xKwCVSaIWfPBIs2O2S8HGv
12TXYkVgG+9jrqhrA6TqTQH3NC/0LUft4L+Twy9WFWGkGZ8TTV0H9Bk+x4Mj8uji
yOnCY3Mm8BlUERCwXpZDxuZxo3bVzOaDohwsqf3+KqB+QDf50qdnb7RQsUQnJ5WQ
XJhXbdfWLmEG3woYbV9wXMh8SMGwUDZ/GzvtzgG2/mJCw8jIaoRO/6ZEMYzXzkxH
hBUmp9kccpRm95S6ZjZ9aMgnQn7XTH8BqYm0Bi8Y21NDZTBcfFDjbKPwfLyZquiP
6cwBniRc2Kal4IFN0AGBy1sf0PyZsTnPM7EYuxMvw+PY4yepuVJ+67CGP2QS9Yh6
aA1AqkT5NRMGJ0DQA+2jG4oiGMs0Kp1kmasp9RCZArFWKjm4on/yTK275jEugNwv
EU8cfVV8lS1P+PtU+zvSemPmiNlT+wu+W+klu2rYqIIoKrKnHDNpCN/2Y5Z4glCY
Z9VgFBfBhLYSD+msXKakDT39MDhst6CuVJzoiKuaAo03VCRvZY8Q0DyraEz8MHjv
qL8d/akdVrL0mRvOMZfGgOE5XoYpZ6tLYvW9P8DV+DelrgmJILGMW9wNYQV7CHHK
M6gMB4tS0m5xyVkeiyNC1SjPhAWJq1lw46/GTeK6+qy/ndvfWxXsFiitwRVevOjP
8c2H15seYwzIuam1yXT26Yt1JCccn3DxjbHEemjlBBjaFiUuZrw2RnoNv6lF82Hj
lNAixCawVsyfUl8oiQK9lNcpsaUsTw9z2mCyyoRkkPUEcyNbPN19ZvOoeoRIkvfS
3ddpNC3NERbJkf0iBTcef1AYxwp8vHADqiYwgqY3gbLgXHDrkXQ2NNEZLlsdp0lQ
u+bt2XEmuLiq8qHDmvGReYbjIB7CQO4BPkDZrPLFp6g8NSS8BB9c0VjB9e4G5+bU
e5HRXOxRqWqR7B1/5d4avwseiiTkA87lSYRCl1pqc9C+Si0yi4d18/Yhga8XXVY9
BwFQ0irihAJthwXDHV/mcEk5tuNONiQsSfW1rlzCBY7UR+Go9Qu83EhWzPUT/MIp
iPfBW5jhcRHchQatkBps1REUTHnT9838OY74zq0vtTlq6XUmEmVkaiaKQ89RBRZa
Nd6jq6z38O/KAjhPI17A08u9l1X+2rZw4XPMhjjcFiu15oic2nmbd/IEx3V5NB3X
lfvDHK4G+rBRnjNHCeQSFKTokAVGeXYs1YyByKoeTv2N1k6C3a1tqQdYTIB3vHd4
MxkKqnaMbZS57TlY6nktQm1Kg0/c7qr/zzhFuLfw1/2NEOM0MqYGxKWvbb3Gxa6d
e1uApTKmvc9M3+YWan7jZzBGLgs0jA739CBx2c13wHq43slwGt8E8AtmpP+6JSrd
sm4gHSO3Do963zUHktdoTQsNV43bPQvyGDFZM/jwBrhcQiHfTqyx1OnPYVi2+/Ub
zhe2bXPks7otICLwgEXnwZRNna73FleCkrb2W26kloLV1qA5wbeOIZbQiYK3igpR
dF5xbRS5GQgO3hGfX5d15iBUpfPu2qTsKoXg2GmyUechCgV7XStBbK0Dk5udQqjQ
C0uijP00iHM0NKuQMTpTCo5eqNWNBR7s1lpFnpTSP8CDn/++76Z5ngQL22mGmaRb
PDlIoarZE0K0/htt8SvJksv6fJuq3TKBYjsD2m16lUn7yyrAgA60haaj1zmaTT8U
NO6b8ZwIym+ZJRsdfnu8LjOuu5FmBBb9HFoPjjpaj4oKt9oyJADa1C5lzJiULbCR
TnwvjihS9CJIOWqWfUd7P4JDVP2RY/8BoFOBso+ZIS/i1a62atZ41RzvRTWbWe7E
hI5FyhfRBsxOlhGpSZtaLw7wRsI6DnQlZ7YccimxbUUzemyyxeFYZYlviooj7yyq
PQ7BOGTm9mzNZET23ARE3UDEkB2gjHgxe9HXESse1wVH7DMgMzBbF4a0THLSY0mM
cLKDuc6W376UWr+E8VsOnlzbFW6mlTpMVybBM8aBglL1F0ypzpudFx1SjNtNIjWn
et7lMgjbpYDMiN4lPM02R5DSLhK+0F46l48d3rP5JMfdvxci8L6icFfGd+GaL+xS
k7oqe56iTLWGXzXiXEvfCcx5HogvXAN0Bi4OSUVAVgfuk9I3WII2Zu5r7wk9gYhy
IA7IzpmyFL1swNN2vQF1YoI+gKZHwX0JVOkfmUpe+9P/1wM+sUDkbX5HQODdpZvT
ljigFUez9W8LwhVdrAFXQoMgcImyxTfAw9/7p+gBIa2w4fEkNtAHgpWm4YaCq136
dELDIe8LSdzJQd2CK3ODa4iZpPqGenO3jiG60cxRuP31fO7sMNaUIPJjTCok/P9a
n9vKjooKfdfkqVBPU1U/SMILAVmE5TRBZZirLNccDg/JMFms5gTXjDO9AoYAV+S3
xESaGfPsEimk0dn8Ko1FdL6xqjBkvaX/uaW6UPKtFSG36aZVpCXq4yVibvrpjMJ0
0u55pkBNqActzQoc+FDXHJfQbFolWyQohK9I8jfGrKXyIEzBhV3v/ic9uBfyC/T2
iK4bG5nIRT6XbgopvDlbrybcubpWk4ZNYxi8+OBuLOOhivHM7/lyQ6f8F797sXhV
L8DHUS/H5VvpVIhJKhNTk4rbVsf5INTss3us6skDFmD6x9WlsMh+AWzOA+BsyPXs
JmHCuWJ/6uvWgLnlYHa67UmnNUXIv6tNtJxltP1g1fyKYDkdOzOpGWu9SDwkpmPO
LmcPxxeMegpOxqgIUgL0m2RPEO61o1vYgMRQVOkWbGs7Q6C4+/NFPZChz/1jEBYK
lmUjrlbJBcFGVQVtPi3mnYwIULV6dx/Qvlo98D4YdKT8ArCmN/pppUgs/zXvdZZW
LASXDpyS/m32YyrmI+3aFjwHx++JRJpTVCV5oJ3kMuqgjdrxPcQMzqx9wV5kgo3C
GCpvHtQMcJTsN6WnJXTLHcPJysP7H6YC0AGRcGtFut64ysvsHkwdtA9hZsTZ4UFU
JviWh1m19nsBgeUqRtnimHsID/1it3FGiubjyVhPSi60xs3MiaGRitI+eiTZpvNU
tKO3GIjT5K6vUiVb42z6CJMQeFlGncWmzXpvmQdXK6TkhaV1j3//vSOggGIVUJc2
ZyBpCphGG7gccXIS15pNybyodUy8YnC4dVkeR8eLtsssBM+Vz/p7yNb/jJSBUYJM
Z12Buv0sFzTZSmB1ANVq4IQbk11Ny7PhgeTe9p7NnTY6YlozCw4BZGmqWC9u2xUH
5r57DSOhSv3qG+vS2DFOxzq2TYdaQRiifwF2IYxYOe8wQog3UH8HlY7HOqcvwxQ2
SY5ifKQwQBFM589xRJhUphsubvMYrlFizEe9zXTpzk76IMfWSGgBv/cdm+qROanV
0x/g9MCFiq2t7ziG1di98PX4lBnPlDhXVWKkfTJ47QM4cobZGp1XvtqBf2zxshej
iXVzAZ9xoc7tupBwSTdGh94f4fvT0aut9ILMKlvTbmwjLfwc4txRjoKqiddorVQ9
ToxLVoVgWRi/Mp5SuQm9We3cMu6qsJbbWaz8nxPT+k2WHNsZJFFMRl/u20XtUiD6
qYWcXOr8GqokRMfVm9IT5jS/rDLbMMXjYDMvTEAMBErbzlhZu6HuACuq31UfGFMi
3OeydZqk9UKCPKGqLKfcCTRcTtdM5Xpmv01ixFDLECp8UUlBk5f/leldHozW2xQR
bwsPSyppr4vvRJDe7fKooeh4y2aelYV/GXDEqjVVNABz0dqi38TC8xhdmnnX9Lgg
00MRlPtF4bytRc73hflg8NpkCZzcKjtdllYb3A5RzU+L18uKRe+r8ig2wlyULn0u
W2PHpHHzSh99DXZM052v7ezp92NdiFR/W9LbYxhAuqkz8JqohRzGEjQEQCAc8Akw
g0hVO7Wa7cnJD246sOoit26hhqW5Qm2BTb/eX77MKEFLy4ANlGJtKb8GcKBMDj3y
/h3fbH5YT68KRFSAytocsM6PlajmXPW/38jcTdXfBuhBDbRtM9PZ9OJhFrGBBye9
q9LvbsZ9t+XMFRtUGMOdxQN1gQ/KBVJEdQ8nQPlB7WOiCksbA8SI8nevAF7g7cs+
9AIamXa8ocCFO4skLRp+U/c0QbGB5QhlZ51JI9KqKgGhhQFmgIogLy1ogV+85Sx3
9Jw3wG92EWqnG2NhJN5HxZwe08mO93YCdcUI+AJpC35OWE10SZ7ZOz7816Lq4k82
sXSHzw+9Ji+W5dZwEvykSv/a+suO9ECrhm5wzo2kYylss1294xjxCodYsEZiyCiD
k8KCCCde9hUQluy7lE5whkNDx837fRFZWhGtbnkt2nOnCGC6saS80srQRYdz7xTR
QsyHypdNzv5hMfnOs/qN62x+ly/Irndxy4qoJyiHrQOzM61kR+CGCqWMNyDyDA1r
m+CRSNRsb07EqEpLIxTLaX1WEjQvzejTPSDDqP+pjMzbFj7ox3Acpdb8ae57q35+
HARWhQ0vsVp9oxjoznCPhB1AojeAmIy+yHKCoy7saFwxoRmq6EbfXMc5kQDzBWKc
KmP6TI+JehwK6X60GL3OwLGI+IyZ6cGZ5hucxt+9d/GTREGzpfnmOIjBjLRENsyD
/TCrETbJMiCRrZ8R+S/VPLS9p3q518Ylw56yaUW9+4YbhtsOHNHzMO3R1nbWctW7
oNWyVYHojUpyqgbgNaxs8stalLUWjyjVf1eHqMorGKazBngzIvFBzVc1OhRrERb3
zRkXprtU62rwegHOwo897og0LrE8PCk7xyjd9alD2R55E37XrfkZoagfITJReeSM
IaYALRX5cxISd8X2GA2u9hteOmvgEC35mF0T5PVn1faO0BJHUlL6twiscshzcUgE
Tj4mjAq3+oJBOpg/d9kkHBXT7ttdRUBpbT8hgjlyVj09C2HN927S61LEXgNSEicJ
u10hQibPplOCYgZd2Hur5aokNLeHXEu/D7bYq79r67i4dmYSfgU0Mju5I64r17GS
TlNlBBGb5qDt9dFuuLyt7NEYHJpgNT9OA9Do7WH8/8FCpmxHtM6ynsFgs28D4v/H
vmJ5pDa+w+Tfp2EgGXmjF1CiGRNAKgQ/IPe3Sj2/XW23P1yCI03xWWI9l3v/uHit
S6NNqx6cBzdoiJrgDSmE7Kekd1uL46gdpcTw6WtL5jtiLkDfMpA6wHSw/eELWd9s
b14jH5WlZcsLmeCdaQGG7xwLj29w1I4AQrWl4chVs3NjCRgYUIRZJoSPZvx/VHOS
cji7G+zsooRsoO+qkF0QngVPV2aNJ7FnfC9B4jtOMeEGlMmZdbTz5jG5h2Bn/km0
TAG1oOjwrHyfYY8re3TtkWHd7BVJuSYjW/iTFYVr8jTQnJiHb3zfV9eD99JLy4sM
NXWMepKg4M1bb0wFHVeyWWwMURgYmfeF4TN6EAmcI7P+pu/0sxvVFWd2rZEt/8xB
iTntPkOa089kFArmaXkY0Pm08Y1Q24723NyPBCdHqk+XPVg9liVAgIxvVMr1/iiy
UNxXGu6DBwyND4yhSApKSrtMMnKAH4OO+CM8HpL1CPXi/j+aDKtjjQBCdMhZPCtW
Ki/6VSNc0LC16HSLDCSPbVVjU1DvGdlXS6S2tzK/k0xB1APCz6nlFJJFOAhMo3gc
JWlAifKpsIdZAmcxXVWKNLP3NivvPOWVZdK2yUqd2FBV7UgpGKsV9njtt17YPASZ
faLyzSBRKeuqblrUhw52GHKc+zJHV4j918MLBOu7A3s/HFHqeXI/XwtZ6GD87BjE
Zp+KXTa7GzFVn+chvUVChaOVVzFz//gcR0Z0rhLr00A0aUW34PuaEXbJEt+2tEXL
TXpIUE6h5C94WvAz2aKb7gxVGgkZ2oyrILuxtTdcBTjv31q90XRdaGJIAP4nOstS
0ih++b4JwBpWQWlYlvxfJzSmrV7+BA1YbVqf4w2lMQACGt95Sa6hVttGpKY3QVtG
wQZOJqK0ox1aM0vllyH5ze57eGJDNL1x5YSqjHQUd9W2ZqI9dHf9JhO97KEyAvj1
OhPyGELxds5rtVqP+3TqB3QOzxj9yvRz/GInmKyEto5UTaDgWfC3foIQNqFWzrs+
U8fFCRLN1D4OPCjd+5C6LbVt4YqDcZScoaWPqdVHTWoTZGYcghx+EY0VZQaH9+le
Sd9jkQe7pJ7ga9Hoq3GsbFdXY3EN1gtiooWS+4ZzE1+8ycdTKnIWQM7jfM5Sqr3X
G5TFU/4MUl9Il1zRxsqKuPnrF64JGCNgzMMUOXfqgE8RfcHRhP69eJE53C31QNXY
0XUWDnIPl88h9WU3JF+lvlEbKmcIwHZWJgqA67JMmfVdacyY5mWPIHMovB+0+d76
k4NXNJfbkCp9BYzGfivRgKlbzKZBlbrjd0Svig6nDzgXyWJpnT0FtUY1ckjTSsXl
S/PE1KttnCWqeEoe104vP3S8YyBktfW1ZjAUUlEiBdK64ULKkIo7/tBy0h+kmiPZ
2GEcDOjE/QCAjd5sPjFvlY61q3nwQLwvjeNy50gGQvFYHQU0shLRwCK/6pHSNLM0
HAuQgfIs1bgxnApbV3YqlqOuSp6plVMFLkPSdP9gn20DcGIIDrzzalunOpRSjv4i
cfTh/9F74VJlnpE9/TBfXZyRKDW8ttZtCqZCBLjVCr544EJHZQ4NPe0GB09/aGej
MFrWycZyLeQT8YQxqAnlixOmh1YrMMfZH1hTxLksAZflGXuc+3MiMtw1kd2v8R83
6TZLymf9Z9RQTckfB2pJ+MHpEgaMtPr/uLy+Rih1gGJmmiOjqTkWJOSeslxatyuA
mFf0AA5sfvlA0lZPVTNwSrJJMz7Cm2bE27l21nawkylWfMLZhniYDayQLk9I3wWS
ZEHXuuzAEahZl26RPXDjn0dDSzGqeCaqaixyVpAVWqujSo3aRKYppF1IRFJesnaR
zAomK/3WgzDJBJzzFEjDskm4mPoEq8EdFwlYhWfNPWE/w99pfzR7HXqzTFSvMevE
XIDjNugMkRy05dN/YskR8SfbjCdpzXM3MVBl6swd3Q9/oIpNZylvCubnyxZ+CfCw
bI+jOtXawOLAWKSgh2SrDJ6JoPPfzBoaDKCgq9EEMjU19hn/IGW6K0usnt41jZCY
tYMiBClGc9bbcO/9UY/gv2fYWm2heUs1DbzH4BsfnInnMYgGbpaKhpfaeXGoXx5V
yPN2XXXDtIVqbpOAbqcjA4OBsWsTIUcI7c56JA7QVbuYmUZazJ5kfEciUy5I76tr
bYdlZ39rDLSO61t1Zly+pj7zEcrljBQsO++ne0x9ONvFuw2UugxUDqc9CIrzxx3L
8AXl5vMfdVDRVzLNNIKTjLA0Apxoz0LvgktiqBm1f5B/ZR3cEipXxabh5bSPIn/k
R0UYIBHK5A8mo289HTPXs3y0m4v4wcTaTpbYDhkxYKEYuhykB1u/xaeTMUREQFnl
GEaU8paP0hwQld3dEIcFo14zKBc4l1ZuJAviBddyr7EGk2HGtDv5lX03hLIn8OWH
tj03d4Ym7Acr/sjfI7slcKpxBRGXFEghTiYtTqNi2+C8qDvG0Yrwyl8iB/LrDT8I
T28CTOyF0tDw2SUolB2+M3y3Zr7S+wEBXcZKRRSmt5yofyzBGwb3M2f2isG6/smn
u1BElgVNULTX/znXLysMuzdQAV5rz5RQCNnXCQsgNQXw1UHHU023P6N2gR7ov4NE
dfag3Z8q+uTRWZLhyWX2BHp9N5F5uIwlC86zz//8aXQhup/ijVFogWUZc+V5ohnN
j1TbWLQaWngFC6lCDUthTnmWPYNGlTv5o6dpoATod+b+dne0ZUkgqJvqAdaJ2U93
jKNe5csiCnNfkniv8bI/CgDp8rgPHHcJtykFSFf+ky4De1tKtSoDKhmGh03k9mgx
6Tw/qS/hKS+C/kjw2s+C6fgNFly5X59Um+kOPe57uT08sfIXvhij+hTDIqmhNblf
PPG9HvCIs8g9dIoCxw7isyQjR2ABtJp1Mb5NTZFzi3dOP8pOIKkZUWymTB2/JaPQ
yj8BrF28+ZkHGNP/74dH0+HImdZqyNQrIIfWmIXTb6zL9DXeg6/LjO4LXk++5B+A
fduuDrsbnNGOFS0Prhk37KINBqJcfIYbS64q35wiuPBY2O0YyEPm9BQjrffSoWO2
rQKFiLSipc17rp6Hvfb/56iS0k/mg/m5Wf1vOhlG8oUBbQktWwXIswqTcRl0mEVv
MoDQvgG+spgIPi0Z26pJv8HtEE8wLueaeck6EaH0UBNk0LCaP1OuPSkYd8EpJkT+
8127E/YmHepmRNutKUgRVR6DxYOpONbUFuKDqeFnbD5Sti5Ic13NGy15W7ea/BUR
ZN0ECi4mjlUsGkT4ab4aGTZGzZTZWW5JjCZ/X8KB918E8hlbwcUup/p5laHdPc7h
nn9j+ANvBIubXKrMRqrqABIMkBQRFDR0hCZGDY2EEI6d7HVaod/0BGipLIAps+W0
s888atfC+mzND/KtIg30jJ1uJHOOU29RKCaNsd8I3ClIp5P7kbhhmsWnaZtZhUdP
sIu0YRcEKalx+2RnZYMuD2Ng3jexkeLCbNpBllluol8CsbMuPNiL15zEYARfrt4B
xugWKIo7MXM1KNgNNjvOq4Wek8muLf6kQvx2RLDXvjxc2vHH7k1CLQMF3ZOpYzM/
BsV2ZNz+/XdqZEpSMwPaIJ4vFWFmNdvfstv7qwX3bxSObX/YZ4W6xMIMegjobvlq
EtEbwFZPd1HxltTch4GGtyYUrw1Rc/fjN7mBaVZsgoc8HoG2dlZMy2HbqsXrPBBU
Mc5JxxtmOsvsl65weoAq2J1AhDCYw/ZrnyiFAbth1EZExtEAsdPtAVZuGG4RGQ7b
5zTDYBnMBndj883M+44ZafIZAAQAOKT9I4xdAjRse0RnfQUXDxg+X6GJTvBXoptI
YXfs0grBHI1dLzppTXEVYPGMJ3vv9DORxWy/EKvYSIGvbq4/W17ju55YoLmep9Zp
76bWv2cWOHg++y3C5AK+oi6SLQgkIRftkB2h0Zkv9ci8/BVbMDu8y/BKSuGRCbNB
bsqqgkwfzMcTk0JxJ1Vvd2J//3w3t6ugpNTPEbtzcs8SH32SYXFCmwSoVffdsqo5
iI6dq5Iok+hB0uixv4qJLZWJn8yHH5ciXzZnEmN49yH2wS6xbEPxB3Et2bA4qNJm
Ya5f8MbRvArbzZP0nWjBhlEqlCXkBkwEkY+TVyNFcTcjPrvsNNX+J2glKQ+gK229
c1+RitF5bZzOLu/kyKnoxjYQjsoOSfaWFqOV93W9SQFbbpuzWqIAIOb11D3DQnHl
HUDhS6f8lQymIfY470+3RHj6TUfzvLWuWj8j1/xCS+ebJIy6PLlPKcgbNcPL2HdD
kBuoTixV1HeSF3tTpRXJKyk6oQyffU0SQv7D0WDdRSyc8KtkBHC7mtPwpnCQFLqQ
L9f2nQXPceRHnkAMX8NprSthSMVyOR2a8pK6vNzRUbJWOTAt1Lfglr210ss1lGlo
q2v6f+E0O+tHXNPnX6fz2vBkHElRedpSJaqWM0oCxsxj7Hkqvai8FL1dIk1Wafio
9SrRFkvqbStgvD1Shg4HjWouX6Tuda838gfgJ6JNT9kITI9EK4HlUk0A/q44q+OK
JDEg7rHE+f9dXg6ZvDz2P4sx3gn1m3tVn07idmCRFXx6xqo+H9FvNv/BQIhZIIKP
SnN4tZ8j2RQyYGyEF049I6pVkgio8FfigVMFnZ+JHNAXZJrUNxLnL7/rp/4/S1Os
Kg7EdWOpct7N1juXtLvrs9vYyU3CxzCP/208kid632iKEeWWz8l0aeew4aNY1Xdq
aelL1LsjJwy2yRAiX6MU/3ZusS/NmcvpLH64FPAU2hIeWpiBKp8CXqqlLPc5bj6n
O/KjQpvSu/kbHOdXQYOxnMialPpMswS/CL2E1N6f7E4ph+/DWNfzu6pFYk6fTOh2
89/FCW8ZBmbge6m3Bl52IGyCsqyU796/D9tLEb1FnZZZV7Zr6P8wzF42cpVU5/fn
TXkelw9jek27iYGtl3k2SOz65MOKkFNqicaQm8DZluqPEPSUK3CFKe3gJ0itcXEp
V3UGDBlnmP/pxW8HrqgsFZZ5Dqpq8nRp8haymWoM75NZ9cxnhrN6iwNEb0WBhroy
Yliu4T9kb8864B/j8wLuYEB0d1jAZH1+uK5R0LUU81k/UQq+ChoTmI7TzGHctgDJ
dmZSFjKhCrGObAehA7JDXogb7GZeZ2gg4jlJOja/VCzRH1oOjR7ex7uhWd1fGHqW
/oAAGaX+DUNg/x7B09w3NyKTqBD+rAJyVzZta7bc0hQoUrbVB1xNqtr74soZ9Uew
QnMZIQNvJC0GiuIxQ4sDPMhokizpkhdyEZdLAed7PqQ6HQFy5m46WLgjj7soUg+/
Dv5soi+qAaZA8C/TLsCmpfSKOgQzd+OIQ0cb063A7MP9zS0AXcGx1ecWfnrp7ToI
jbeEuTKi9oAhutJw+HPWQmk2P54jJg8DgOUyBHtsyf6/jGRVKNmu1eeeWAEUE/6Z
XVt+KILhl9mipXwydO/8efvX04ocuKBfMVyZK5OVVLP/AC+HsFBmKtBDwdU9KZXe
Xiv08eVXycuyMrk14aiUwiMK76WXW5fdIxxFVHQIlSCILixZA3+GOmp+QEIylpdu
BQ4YUrpgwa6ZkldLiwNGNA98pmRGpAPrkeJK9h4pugYud1zfjE7YKu6BohUSImzA
joWzaCnjM0kD9nC8WCg9KtxVQo7Fs3iyrTegG1qISANLuuxlh7CXNDgSma+RmDNP
UswlRY853FLNf5e+SPjGRxkZOkHm6jOkpXM1DDfA6UldMTPrFprowEWlCcqNWNyo
9QoEOWqrHAniwjgZaTuI9W3XpCHd9tbcVMs6OI1S7yTmTF13bPb6lxuADV4fPZM7
Du9CVlXr3fTjKT1NJioC3ZfVwtt188zFV7NpZ2v+LY+FYRRnfyd8+ckDxT1NNCJI
XD+lw+KobxXyPxRbD/4FECWaNixHn9LRbrSSq01XDh8g8qJy7tm5XcvguDLHQlvR
gGpC48q3ggqYJ83doXbaL8VEt3EcM6YoyNBiT/u1nxxuwqkDq7bV346gS6cIKmnV
IxlWHKc0mxGi7p1qIZhoQDctWnkna9nHZStp4t+CkKUJnzwUuXGFFdp+rd1H/5m7
PB14elXO7RGk1AaSkNA2xGkfL09Ta0mB1cG8anlsSQzO2I6Huxa3HZUnAsVZ21Mp
dcApFtN8FA3iBmfsjZK78DHxw8XmKx8jlTtWDpBs9937SSVMv+hIM0omJua3bu7F
If8JOXvp76ENnoTig5HsRB/08A/JorRl3BfagPlWih09p9GYLnqdfGrzaL7wfK07
nlPv1X84klNOURaTByfRDZrYHlKy3fE3v5DWhadk4Pf45opF6/dhbzcHKqfkLr8P
wP7JluFBFRWC4VOY05CL61UxmTBXMTvq9Q1l8YSU93x6aPaqaiNpknEs2FIHbdAV
21VlYfKKhknN8mNH6WQwSCzZF2sRLMMPe0nDTSwyZO1y71G8ZWe1qmrz7kS63u37
wh6TVb4SnthNmww7GHfpyh2+76YFfQpRr55g0I5QNMlkZHVBz1+QPVgoJtqGjw/J
TdfaHq8Gtt63eemYRYHl1l9NfcqhK33zUL/UAkL3yEWGecgKjcxTrDK6j+Ah5bBx
Xbk8mL9t3MI6K9hwPO6RjzHhHC2mgvJePkXmn353YAY+7tpGIIK2E911KHgxZ56m
xhXgDUozDrXmcWo8w7N3gxP0Q1HVAps6gdETGr8xFC3p490KK8u+qLDRTLqcfIud
8j7qxKZU6EyGFl4ODa2z8ymORC4Vz2xPvsiWliCXl9G1ZCEDjgO0KySXn8esaoG2
0kOVV1vZJj+yjygGsRbijPl4I1Wc+ypus4Mud397xPBK1YIRzi+go15f8S1553ov
LEpSGqaldJQrwvVHRF/njeXu3adErO1xnypivQ7ozn/vTar1ISSkHHaCyex37GfS
DNtJGwz4BzegcIAkhIoaXeSJaCky9+ei/7lZgbAgJVi6q7h3VAOGMHrSPkwVVXeW
8NWDU2l+2J/3nfnPp21HUjAgluxqi6JxfqX1n34b/jBYgcbgFmAotjkC39bzzFWf
YCmIm03VRhKwdZ5RTbp6Z/+vAwxgvVWq0jULLHKFitNJ7xlUlGFNME+jytFH460R
yfv5eXD3HnsSNSmg1Hl81OgzxdufyZV93tFdT+nBVgQ3nGoYv0Z131WQVhchquVI
MS4SdBlAeCdaFwy6JcIsRIhnwqwjFf6r9K4RqhRkZhnG46nV32M2OlaH5adoSPwH
EFcrT4HIbbQ9haIXMzn70ZaLPsliN1b+/UpgMVVcQQxlG1usvilOkZRc2xUsAv/F
DPszj7XQM4cpwMDbTChB+f0UhSfBSiDipBdwu4p/vFbT3Nmz1YTMRmqA3wq0y2k1
SA8Zrtech5CvN2EeBxxeIoJ4KTAgu4bQg/dKDYWvVjO4TdaPxs3Muj8FI3aaAhDY
gvxwT2iuFtjbVFCeEsaTqmZAd+KCJUlsuLbCFxiDCR7LH4egO2DVIl9YW/UiEuP4
btraM4VjCMnOuuQdnVl/1KT9SVe5wymKvRsWNq/2nTm3lKxvT6jcgww8V57CBeQj
HBOh5cFFvstgPBcRiFwRzen/nuFGA4AXUodhbPgm1ZQq4cmDH1os+rpzBRmS/Gmt
DgdEtFzoML6HRqndUvB4hhlF2eop5iLR11KCN1QzLKU6x+X+3MfkhryWi7ngxlnp
solaiy7/SlthsoFb+N0jq4aU9cZ7spvJnNr4ZSDGVMIWyaZZYf7sPtUxBTMh59Zf
h4mIBiLMGQN8y+M/mArTX466B4QgMaDCRkIxx6YfYrFD+SJd/PBh6mrjo/NN/Cvj
xS6BvDCDIzOkGG3HE7SsyAGNQ7YMLuO9xIfGS6wvglHsQYcftYpVtVlgoGXNC+pq
JRxj/qaK2h5kB8uZtrWd5ZgXZXmS4+hsioy4BpsEcgzwNOAzH+AtkOQHYYvgLy5I
+x4W2oNl6V28oog7tt9Z/rvtVqa3WfBfc1sSdBLBWb2wS0RfNuM/YnpGsmMHUWyI
onY9RHsT4OmHdWDt87w1LmREvrWqjmiz49U4IAd5VXo57IOIq0VqiBKa00VWmMkb
Zxudqn/LcygLU41mua7xEGCxXb04cTQE94mJ+fzWavsmQdi+bEceGXFDscjh7ClI
2tCCeF38/9NkhkpSs1Y8js5qfbPzDpE9kvh+KU2k4T+9ev9jH3fFNx4ryK37LfOu
l5S+jQKyuH3QSpIJYfg7CZLkcVz/mrEls+1i9Jprb5DalxD8lGCso4nMy7zqI7Cr
5c9xlWpXUsNpSh36C+OlKAyM2OiLMejx6xEYEUxlUO8EHhHE/YCep7EEhwEHDhS/
CERbTzTPalDdg20h0vDoVfA/8cOFf23sHzUp4YFJRrUCS7MhZlzzryDx5EeKLSWn
HmUI9MzBu640IX3wTOBNPdrBESanOAx/JDinQJZrfrvtMyp8D7Bbxk0UbBjGgd5g
5JneH5bsE0HBLTBBgtXFi0mFZn+4heHOrfplPDcfDz5Mh1QZbqi2GLKboLN2ll7z
wrGB3AVkfei2BnZ6sdMQwjEJULYIR4LQ/KxWJHN1Mg7vlUz7Vg0G1t3jymYYBRVB
0NAA8B7yWbWUmL8Jum+KV6tR59qGE9QIW6JpaBPfvHxL8H8p2xr4KZSSLAIJaNnt
Gavm4iallKN0LGWJkOTFJOVUC4Teg/nSifyCiI31dM5pXK+UjBHDvq+kvM5N9oG5
4VDobXZ1HHkQwgBb2LRgCjnZqTCRNuRytDXjtznA122IZl8ZCEfCokaYhwqmEAqZ
Z4y26OrJlGY5AAK15Mnn7JB/ldH4iItIfAnxglwlkCFTb3LaZ0O+Suet2LlJ73+3
VC9E84dv7mtz7wxpP//T2hiB4kPTBQWb4oY+fRkbg+T023j9wat8sZq7PbQERd0z
mDfvH6eeU5tkzVRgXg3t23x/7C6kVfh9bHFuiPbXZlLEMDOTAyqDtrbSs5BI5SvF
Df5BEQGvfHYett54qtcVlZpFBKtXPDPNXLx1486qgT1TxeVeK9vhBEFSjmM+7NFD
85r48pqEDIS3xgSjEJx3hT8RjxTEmb2b1thm+LahwgdTqv8c3R7G+aPxkT5yWB4T
ew4vjokrX5PvTUr9IAZqte1bU3oAApVxWnkcCMzT6stW/DkMS97Yh5JBaajvGc6t
H8hOp0BfBD3SvnF7qLjxsHq4KSb5KX9rhAuhSpc+5QxV8q3EbQUtwKyfCmryfjr/
8YW8lUPDS4cbzdbUmsM1tSw/SeIdL3uVcibl1c0AY49m5o16MIORsCzdcTWYSO/v
iXzCkgcb5DaqY5J2Ot720u5zMR2MsUZD71EkzoOejH8bTs57p/svCuuKwxaYjrSO
SVZBNwhqv750oJNd0yIJI6iCQEXoaxhYkI1d+avUDgrbBpuzH8vQ32jJm2xX89is
VVtJbRPhqrFHOC2tFVMRuZFxvkIUHMUji2RIA5rfrtWergayiQf4EZ3mGNFZ/Ynr
NDp/Z8PQxUIvub/0rzrGWlkcuAaJf0N3g1cUICSFJJQZp8EshjqbLz67Oek3E8Sc
m4rlZomy6uQIDr/Rk0U8UZCFNF1HrgJqkOJ2Ws1n4KNouHmV7gy3K3qM4ZabTkXa
uHKIQPWeL9kSxT6pVI7CNJMdQQv/54P6Utn0E6bLWRWpiTQeIM6VZoP+FCzHhKOA
rVToUSwEpGB5Dy6lzVikeO6g7lDL0uq59ZVTsK/RK88NKuiSCwUQ6hBABBHKxzhr
jWepvw8gFIuyFKqN5VOAWLdciMWJMBjgdf2VCT2QgHODNaL9MgQI443Qujf52Qxo
kN8BlWNVuW/Im32piJWGJ1KF5RHVvKFzEdfw5a1pib9i2YZX9qXE085Bd9DpEsgu
+9FQ8inhvEmdC7nuAablJlgCG0IDojg0tTbwVa0JozdzwqxXzSOJ6fhy6Qxxx/ZP
/P8E7hPUW1+buAxvHkvLKDGDc2LiBw5nBZgwWy61mLxIqouz59FMhkwhBzjo9t0J
4FOX9yJ+rPxOiARTTtvgN9PjtbXQTkjtUVRvIkAN51Uu4e8XZwIFDOGlVn3NqZQO
C1QsBz66nsJ4n/YChJvUVhFYeZtzvipIpx1GMXN15zkDX5d4XR5erSGMadMLOFnV
f9aEstb9Bh1wOav2ZGXr/szINbZ+TGEXtitPiIMuUdDSRQ+LwV8oHCHoFhMNgzPP
jXuAxE6ZrwB3xWSakP3gPY9G4QaIqH8YYwm1IVLwBHoB9qZZ1cgyHgkrIxeaeW56
5ZgOvb7KiEyLMlj0lBkfA+bWzg88RPNwo6cD8Nc4Nf8AM69Y9YcazNKXhT8yw3tx
mk/B/azFli78JliHZqTsCh9cO2Ak+ddBKSfg6cBq6mQE6OU6IGLC9nmk8ABFWQSH
5XaHMm2N6UX2N8/EKpLAzyjTGcPdcyP/OmchXm2Kejb6KpvmeGrXNknQaAdMKsfq
XHJZIy1qclH8508Zs8oEWJI+0o2jV9HOX7gbBD2ZiAIjR9lYQ2PpWa0URZVZ39Va
TcpGtGbk8k0HcnNDujfF6sAkF+wP2UwlQPuaCwJguGMjgh78hLjXcJnCbgYUIVq+
TKM/eCbu+9IIq/LJ6qrB2P+WjpAILtgj8SwXTmWTN75Fqbnu/IRZ3xssQpbB5ktQ
atr46RlsezGpMGtmduufnfrAtvAonV0ey9nsGImupE9CqhS9sgK9ZTBezU7L2B8v
ZIzu6FazWFcea23izERODztf5Lhrvinz+fzbmtTqlUu4sXHQXWT8rz3g/vMg3ruL
Xw25ARbyfx4JF/CwpwDbs0BYTNkXZbHI3eLt+RdlVHy3OdbxRKAKRORIWVxKhBdd
8mrQ2rCKdsxIKmBWtnfoLihkGK+XNeb7e2ISxrkbXjdL/Uw3twZm50NauuuF6rPP
UsBkWQQOm+bkxCaIX6COhW/x6CU8ZnFE4krG63uXeVUxvCGftKx1N7HtEivbfepX
Un5tC1JAtpYX8N+4E1jvpI8KJGLfPGsNT+gsDi2PBYSjE2Khtulu6M436tW1gi1q
4UQcdHadYgoMS4/bzQY34oyTxFyYHLKKspb4Ae8Zm7Z0h/cThELp4F0jPZMv9IKr
Jq59ObqrKcRTFuLyfAYPveU43n+SWN7wKL+R7ycOI2VjhOu6hb+NJY83kmSPCvDR
km581zkWTI9f3ILexogmdPEVDp3fICN0YKEc0YfwfFNaxYgVCj6JtRcBnpMOAS1c
ir2sOjU8cpTBbspb6m86LgIGvyJPNImBFngvZrNXasNLB9MkCe0ybo86YdfPVxou
Yla/3dbAJbL9ygrYj9imr9SpuE/ReooizF7F7nbNmLr3wFDH370h3ITE3Dkj9wHb
Aj38yEilgOUZZXlKTPFE3A9eURVf16r6PGckTkpLYjVSaPLmfKaABcX1gOYUPur7
XiWLzPNnPoxxwqbg6obezjIAj7grNi/UUKzDNHKOo71BVDvJCMpcou+3OoYOG45T
Av2qACVugpR30KgvkpMzdk0U91YFKbeyzu5eOEpPiVMcoO8iKkLrLA983LYnclJm
eWG/iPsg+HpbVYC3Ssrk4yx2Pvbxt7rf+Rl6yMFrBbzyeLhY3qJJd1XDk2cZtmCj
TZxm9tA1RnCJWyo5BfjkWkfO+4bkfVS/Wilyt5y0Dynusx+l0CBusIr79i2o3lmV
exBJfaJtP0DNsyndKX9y3oOcuQc6pTEj4CZTMSAfnVdqKk7y6wxRYiCJB68OPZOO
2Yb+MAAYK39ffDAyKZ5qq85F0I8IsFktphlZ0SIqh0F6aEaT5fZEjT8Zyj+MYLWR
KVtHRlofAnSkvMORrtFygdcRcpqvs/kuWKcSt1TgYDKzMgxijGH6W4RkKhIxbBOq
wMTPzH2aCaPpVTQuAppmlDrZtjPkU1WjML1m5L+Q7LJbTMyADuaylTWLJv1ByZWB
iCD0TSbaTe+TlTMwfr0VukPxAlgE+rQFl6xKUWdDJeAGeSgpE0hUS2DS3kVmE+vk
e1f4h2xB6af5hns/ZxIYbT747aziP1QZStJbwoDjzZ+6+mNmazpSieXNytK4zEwU
e+bLIgvnygOIAVp4Uhyn75d5wyxa7xFYcSjVhxv1EhwS+vnqzM1Ec0xpP/+LI1kE
WpvrwVGHp+urbI0pfwp4C1n+5SOtDR6DRMOMmwkloSC85fWpBm3H5F8vsTzQDXTN
6UIHpQFJFS+O3R68oksATcNzecFJw0kVBACnhYyk9+a1bO9cl1Rllfv1sdirrQSm
voGlYGucelRHQ8eMgJC6RR4w+xPJ2n/jrEnoXS5d8Tq6wtURb2s0ebRSgJ92DgG1
TAmZb8/DhIVk7OX5RC+w6B4BG5VNCaFuwyczsLwFz+AaPxwWhEhq6BfCoi6FGU2B
d409zTYwXCotHNr0Ewvs6mA7WMZ0pae2UZ1EW9+V0NMrR46zkUzKqQhmqSbLMRnE
tb+/mzfAUyZxznmvtsqKMnObNkbAei3Flf+bi7qA2nfLiDPxqdxQCk5UqCtcPM5b
PM6NjeI8DTAuSFY8WdY1mYlVWhkKYLikffLjFJw+S1l5gt70ij+UzbhaAgiJVGbP
+8APR8RBR+Ze1N1K6V9voFi88zfu59bIDodOmljBOsUrBiQPiGYCC8Mkm9GCvCwS
GL2ayU7x1xpjkg5TKtPCUqWLUMWSK+jXBkCqjd0iIx7yxSFGoQaS7KABJJ0ZJR/L
jp131ATwTJZRmGXGVE647fs35vSLODqQ4lgnNHsgqXIah6NnQpMKi0HwMINFD/zg
PrzhNYfCaCWUizP5kekZv38SHjD079dN+qNH8Enl6SEkuUTGfgYrJrclH2LzXzm8
dZkNngYnQ7tSlQMvmk7smLhDfBXz0PWuFfEYOzNkEzS0RlCie9Gi9LENCB1DMwca
QjL8xb0RQYE+MeLwU+YPVGqqy/z+Uxa8wFBasoQ33WEq7SsrHqcLITiarOy8P5VU
jx7cyzsOLV06DoGdMAq3xz3Odnu53HgjNb3WDMui1FbRi+kVO4hmIfgh9SIgIRLC
kFj95EsyWxyIXUOz3/kPxsya4nKkqz6wGuHopSQpXILEhOv1g8OQJrnJestFGu7k
VovuwiRKcoaBNaXJy/VtfgJll2W3//g+9twhOUYPpyc6RBkDZ8Vly7LCeBhLlA86
ek7jh5b9zbyVLCsR9k6V+rVkOSB2kvXMeb8ozvCtuWTsy5SSAWJpsLRjA5mdIzCF
ohTTbDSHfqdRuSijqgsSOfm3dlP40fjbFxSmb/r7PIVNBWZhM9b1RATUM6fyKcmQ
TvqifKEsLBijn3seHz2TKiq8gzdcd34KtKaqm42BJMcdyHby4kujR1HfYK5nNQR5
fC4keOlhTsFzqbvAqNl7eLp1g/5PFkZMnd3jbaY/x8wrjSa/vkSwzYTD21LtqEwJ
8q3WQ/CUdVU0aUvzO2D4oxBhwN7yf3v4VHwuOW7ddc+1TTVJnYTVJw5avHIM29wq
xWGV0Mgn0DGNPG0zRw+EXjnv5TRVd5Kawfy9zghPF8y+cC2kc9tMfvh89krzdJhS
pqxTfw9ragQI6WKqzIIPxD31xnPBY1h/WstmY4T15ZE55r6yiBIZb6yLPg5aRnDN
YMFXYDBi+52ga/KvVMOMFpEAzyjlzoic2CCDqYjX7bLhJSUuIwbzLjDSwBODBfTR
iVkhoxa0EqyTDf850xacK7qx8KekG7bCohBO03dQ7F2XGPytnVoZ9Cq1ZDFGfXXD
3ffuG2LjQBAmVUaWA9j0X8C6x4nqNC7ebca05LrCcKEUkQmkTu1+rWyA/AmNnq62
XRBF/o9XcVaqko/UbFoSoxQyB06hbev5LJIgfZZz1d/sAcz6EQqovXkdhk8PfugH
U7K6krW6b+VEOykUyn+8hY23uRmaiinVqJyBpZPc3uBRYP1xRBdFLt2pqwHCZoeF
+HOLcqGNqhHSD12m51Qge0ZVk6TtRIizzYFBnhbgVFKtrU97tCXMeR24gaIjkxEH
H+gdFbdshFvQs6TzvqkqFj7+IA++JKqrCNBfaPfKiuHZ9qV3MeIeSmwksCuOqrIO
pHTz8XYsNH0bCZ/kprBaYQt2qga2DswPKFNWBg7cwHQtzDShNBMTczUMB2VyPg3p
dmqf7PDFwb8FqqZDQn9vCYCXHWi+ZWIIO4pGnr0XJe6QBMBtBLl0BKInEozvUm8C
uWWckIZz5pDhcFWJrG7LQnStGBoRaEQ6fww9KC/b24zlyIkRn+SdTihu2NTGrAFq
c6E8nXJ5VEy3yhovEaDsEYMVXfLUqT9X0qSlmIOfo7gI/wbl8ai4KncXsF/nY62O
oFtNleGEf/n+/ZxEnuggmsup0Uc4yBHt6f27QcjKQyPCB/9QMKmL5lCowR8IVJFD
/pG6Xqr5KFmrcQMD7+6JVNhS76mBdZBGccZOLNRdh2iurgnc/h1Vf7MmEaTmiPao
JNBmO1hU0M8OFdZLN66LNy3CU6VLg8BPXDb6u/n6YRJSJFDPtlvkd3DgZw/406gw
+/jkwmEsbqJIkUGc4gcRp7C2iXYGQTNWQt50bmGn8Iv/6GXDvyh8GxgtnRLRXDpI
yCwr1sMMLqAh2d8MDVmL5BzzUm9aJ/hwpMRR8WfPk/AJ8k3c/s5SO9QOoE3vkZg+
lfuePp/7wbLVGVxIWJ4mdDtn9Xf3hxgUA9BwP2D3wSJ+NFKjfzWCz9VqYakWYQ77
+WbVJEdxmbWZC5sADQlcqjYoynXkvCg3TZcv0b8O7Ng1FRN5l25XIu6ioqfQu5BB
mctgTKuuuJy7kXHhZB+7sl/EHVDKucR0cP3HGPStMlwbWGqJDokfcHlhrn4ZI2qK
OxK/jiOhOkqShQUd5+0EV+MHV7abjgWyo7bS1HYKR8J92OMmAZgfYQUao9LZNn2O
frFb3fqeuB4EXEoSYgNMulmce9Q6p/9i+m9/1COTSKfuFHFDLfRCa7+M6sPf8+BB
n9zwnG5jn8EmbkOz1Z7YzUOnaDzRst2oj5bIy0AS8R0zR5D95TtFYrGxbuRGAP0M
NDrsreWBvx+mIw4WYr23xo3qOgewsHorBGuXwsT2lyYP2HrNyDe2Hks3ABN74nl8
ZbfkXP2bN2DUQK7r7ZO1qNKa6WkpqGBYq3LNiQ8m5RPDWFNGSSx/WRgKvKlTS5nJ
KCFnOaamSDSo8cju0NSf6PoIcLYYx0OcsF9jNPExz85VB4AFRxjhj+Reu7QEiuqI
xYBqhIq+3nFE03ZHHwY+dx+1pKBfWvhIVc20wwnNuELHFSb4XAWnDvs/p7kE6OOJ
1xlzUMy4TNozbeKTk9ARa87JfelkK01q9ndjghKz/tm2pS7o+1KIyQ91r7yNKWtf
9Ru4Rq72nrjSWgNnJwU5vU+Mwj3v48hbRI9oS/DLlygRxMOaTF8OPn4FO4qSUCtc
qTjAVA37Re/hYM05kcdpaUxUkT0OSDTdGs6GqbAC25l4Wha738NFkrveQrTD4Ql3
vCudGGcCPGzGJJUWM/IktIDofexdC0JgZebmSkZzYXJkNf5i8kvH0HtzsvnI4lPQ
c1drMaKIz9VF6EY7VHvQK2bvJamwpDt2vdjWhpCFl26qhoxp4bBEqYydKD9ijL6P
OKBUwdZ4UCe8qfc8tT+LtYzIPHlzCgMj3CAvwBh2H/bgEbP3uWtSWmW28jaeXt5F
9+UcS5P00tCWuUvi2ikvLkPZTTqSuhcX/HjT2regI1DyhVVsmY9tWN9Kmdhzl+h9
hBlQvz/+g8fofdoThK/T6bPCIthunmc+Bf6mXn1Nv8rROUHXXq+hJIeReFnSmvXU
snP1wb97v2kON76w6yssy7/M1+bhFyHjf5U0lrTNesjrdRkuMzjl9wglmvmDRSXD
AWSRCCxXAXhX9+hSGHEjjc1Fmm2Wzuc5SnMSYxN5Sjti3uZiYeGhfOp/BlgmysmK
CkwY3Nn8VVIyUcQMlqyg7/kVVw3rTgMviguIUq7To0HBDDnqLveS/7+KxUqOpUF/
mCiThrVUdzZPpDxccHUv0SKWazAdINEeRR/mIYvAE2XT2obxfker1VC9V6zM5xnT
Z3VnvNIU9r7Wt98SQt7bRpzYeVwFTPgtG318lqWkaVCeqw3gveKkBSnX7M3piDLG
z0PfVwMpzWl4lWwAOKBpNkVGmDnEw2xGh9kfrSoZSpZSL9uKJ2dRJTlzmuNnZ0FY
ebGChFw4auH8wpiLLxCyQf3kAS9Z/IvBBjMzBmtikGgJl+o7DWb7jV6bQONTzxMR
DmxWoYKh0ZLuZN2L3N0bhDbUP/xKzmTQ+H4KGcT+Vi21B4O0kVZ3SjCPcv+e0xVp
MT6Vs9Hzze0qx584A1Q3NJqnDDXTZhpDNbRsd7qgtDw8kkHW8gY0DhLIb1GFEwqn
weGLhQwBnRuGA1lCJ6orvynsTy/VpHj6MothPjOQ+8AHBCwZa11Mj6SEPm649d9h
MwFmkf2K919STPkTzHD3HIr//JG7/B0N317YdT+CSeWMktMgNWSGwhX5ViK1Cj7l
edYG8P2MhlDd1UibIvidvQLnT7XBe75KNRNTQmBFy8kNwL3JeIGNZ68cXobPet0q
xjN5ruUUd4Aj4wwIy9rwlBngwlkYUZhylan031mNLOtofe9wqNGZnoX7wuvLiBDr
zMBsf8raJFhMpf6rw0JTDfSi57qdgLx7l2YdOYo9IxQGNObRmbbKy4afxTa49FtD
mFQbZZsFBTahK+CwKOZmO3NAhofnHJiQrLA615WjZ87tddKge4lFlfQH2PoYm4Z4
Lf77b1GBUUE6dhpdkkXoyAX/c0UJHNh5577rxQzBScAkQpt5dn1+UcuAQbzJSyrm
LZ56Zjx8oEEVfmeUF5sF9Vs6wisu5Lgmm+lXLNZ0aZW3mHwkl/Nm+9YgWTInXv59
bazd4NTF47L920ZrgVmLLf6d329AmsSYc4Eo4fPtLM1akGij5XSksm2W1cm3hqo1
B0xkppj2lSp4TYg0L0SPaSan0gKuKj7linFq+UFq77/bQw9PuAFRcDEeuda4HYBN
v7hJEvynILeqQUZUPcgaQjd1n7HXpgd412CMkTJH6WIzoFRY69V7tpF4YG/+yXR9
P7sUJ4/PnP7scXwVh0hEhUXAb9e/eiepr8OUWQQ9L7Xi+DuEwd2pMlLSaZFkdvHK
x5BNTaxOFt75JO5zhyLsqFbDKA71N0IrnYcvt0MRmLW5algrqiMmRsjTvIYgSAln
rgSXIPBii2qjpDCG3smq2ji8W/x7/j0KeA+6IyRvJ+RsMSZNTE55v45gfpKjc8s/
rt1q+O5dxTua/q8DXSqj5ZQZVeMwKFbNZdsmzTLT1MU26TkTzt6HdB5adtJ3Znxb
XvRth2f1V8n6fINO+Q1faqUZ/sGJkhVMBs/zE5Og/FV5NvAJ2c85+PNeHo+b0b4k
cGx+xLLukaTJN9uwfe0UOVKMdZvRNo+P1RT/6zOUyQa+9Il0oZpzp759Sfr22Fu8
m/EPEi21aHiFNePbwgxyeIurIjiSSgB0sMc2y9rcLm7q5bBvuRvk85hiwcml4Qhz
PsxoyDUjJ0nuH0wUP7Kqwl90XmLRCmLTCIk5YFocpM2uUusBXXZrVwIylW1VRzyO
w3uhgfNTDOUjadGEz15t3FBlgvaViuNs+IEhwsO4fA8NQ1K4oFoZRz7yBzVhzl79
wzkj+7x2Zl7xqCK+ig8kB0fj8AON+iuHXdWHqzEXxBlTKoS162vwrwI0qralkXxZ
AAgUBsE2P3gefK9DbONDYeyg/+T4jr/AnUtlkaTIoHyfII8OmgFkvD6tfgLnf4YO
Lfo7h/TnalngCwq5WEs0O23uMLeJO9YrUKSo3iXVGASrC++b9DdA0ZEd+pCr79hq
vcrjxbvOWQeyjG2a63jPPmTtI28YKbfODozdtCBWm5lYTHmdnC5dO3kZ/9jOMpi1
TkNAgq61ADZn6aOCK6NQj9b9h7B874DravUiW2BrxBFU8Y3LumHauIngwIMSEjXc
4OsHoU9Q58E/FiiY1oRCDetMXGeyeohy6YmOMjgWfP3P9kbEZ5oqBNMUoGJewzaH
eo8Q8ePFZV9FZR314e4c1JF/Ca7dDVek/rP+0puFQi4GT51N8VlhAZttjwRRPu3q
9Ci8oNd6qjfn8tYNIKRMQsTjYeUMqp8LX4HTV8V+xUSMZ9ikr9ZucPUXzRul2oJu
lIdYZPlrAdNwV0mIpIKihEcL6VNZXPrgrNrPLa6re5rwGwNgdCw4DxxuZ5vLSo4C
/6h9HOX26lmsOAza3g9NBs5qMml02kYUqOkOb8dnB/HeUE0ZcotwErxnZoSnj7bU
Xg8e20F2MPq3s20fzoxl4U1OqCI18o/1oCWdYCxZN/H07PPNpg5js4jWhBbkbmoz
+UhZ2TsuqArdGLYuy+9XYDSyc0MvrCluajGEowbD49+kFNv/TtGyL/IHpCwhnu8p
6caStCnnlXcIEDFzvdDO3ToktcqSn6cObDJMpDjmlfaogj8eBMSCSAdV67a9Hg8I
xNUCHwLZEtYnl0XjpGhLWLSX/Ryxm/XTg3Ws4ElJoHx8osrwYdJjdcwUbefL+hQN
sxjXXMXjthfR4lI+c4cAVLJz6tkfo0HszUwdL3QiWKfYKSoylSh1D7wFjVS816Sj
Xdkx97Zi0xE9fs1wia6Z5zYBcABFhoueW6qLHD2kvoUu/Zh2up1h777ZlxtED/Fm
D5y+79yvR4mvmX0U0E93+to6OCcOWaibCbm1VdaAQo4pVBZJXM2+4BgC/eWmOoIV
j5BE3dWLTCwZXPKGeHzZjoqqNzKTQZu2dwEoa/AjW7110kzplM1B/HMj5PZCHFjO
U0iFdvzvaGQ3bHi09Jy5QEO1kdTec66hHzoH0r0uHyJQgsi2T6l6tkJ6h2UoLsIa
GxdxhtYVU6uwjW8ohTNvJRzf8AEa5347xYilXzQ8CQhDJunjjMfm4Jtv0JIC01cB
ysvjuqaWna6BR/p7pPZXMqSpBO0y0KMSGJXHkuVfD4NgDr4LyLdBNuG6cmVX52kr
y9c+Zk8EHUdMYq9bDgFdWvcUuNsx7pjRMATcYpwWv+Dhz2LFi9dGdrinlptEsF03
u73BcsRPwuSyc96BJpun1lE4gQvaVtdj55JbzUjuU5Ll8bs1O4qTnYDxSTbcwM1I
jZF/4RMPL7D7wZbulEKxQXDgM9aOX9tvBjuHrC3tXtOsYR0C6NelvCM5PoPDoHtf
f/2gTGrwE/W22h1uqnoNfmPnQQI6e+9ov8mKZpFPVUk0QTHziXRBP2gxByNvMYmv
kSLdJBRa4DYPaF8wFW1AlCmi7wTuOIb/aggye5DvYVnywozc5/7xcY2ZoNr8UKNx
KjzzhcvZKKTJkW9PY9wZjplM8NpqNsgdtRefF1ZN2Kf+fqQwvxCpNKRuab34fGl/
I85HyprpicZQ/4NIqcIPngcqz/ssEgE5GwZHbGh3INV6eSKWtTkWhtIwtsA/FA0T
Nc1jj1xPCZZPfMte8J4jX4MXe8TVftjfVhRFI8NU0wDw5JEcRZNq58eqkYlsjLJm
WyP/1dDbsOHK1azX1oRszVj9GVcnphrFFXXopAjcX1jeVO9GtpisXIWKOy3rDWiT
N31CxR+jNTRkXCFned3FhtC463ud4pGZT58yoovTRmyAOcOukUq4qAcPGpoB7wZS
pQJgYENmY+0lxNtlXypjyB95Vr02ceW+4J1VvY9p4UI+jPWGQ7R7Ib6cflNzBOpE
MFkd5VwgZ6goVTAhJ/1sfAY4myUFewNRGBS3J7DAUfn46xtqRJ2bQyd3f8zyZGjM
FGPnup7aBvechbb00+uEXOPONrSgQKbX+eu7fkWd5ikHq+O/J4U0BjkqNDcH5UT3
nyGyu0JSwwVINgAyhypXPooszdZBtq258N+WwIZWn7EDQE5AVvBuuq/dwM0t46go
C7pKKvR72rhyVx6TnwvJiiSJjwqN8f6wSaebTyK7A3H6s6amDXgj+Vd//08ocQOB
7hlFTG2bcNYwMNxCkUlnsvAA0FoQDeLYyA0k4VzdB3QvDADX2Q3xm3a1JPaJvnWq
OTiMobk6zxtyDCjZHKZSKJMKPtew8RrHl6U11jsHJE0JMQF3lMJ/YTmGuCxUsHpn
8/1pGMcbXUvinPOyOdLR0KHBIyjwxzQIBgz1SEqGcJWNcZ38eOG30TXb+YZpA7kp
6PXZox1+BaVD39qHsmNp16DQk7vNkOYLiRHkW+prd9TDpPkKO468DPGEXdK9Dtjy
x1+5aVZDxU3jScs0bVqsJL24C9zfF8fBRBMoj9v5utdmLTkvpnUABn6rdy1fwLtR
sd/EnXk0wzdPvnNAXH1LKZlf0vlrsvW20TIAhOtBxaQEExqwm8+STzGRD/IBR3xU
N1kZvn2q4C5aBMHopG3iG8EB+V8xtpwPM2renx8SsD0WsuyRP07P7AOHXj86EBBh
QhZIayY1XXROdCXnCilN55SP1TlVM0xGhhlawq387NzPjQzAbaiQouspE2wjqYjP
s9jnZEKxlfk9YM2xRA+0sGCQkBExhDafL8RzMXD3N1NFw1yKKlOPJOyZlLxG1ocD
sdIYlLXBRVcLRWTgIosCK5fVmZ4nuY9uLyhjsfawlsR3xlENH8fYJ2bMiN2koefm
cOGt72G6lmLDdIgKawAGCOg4jNFAwuXYajhhTZPVlIl55sjcGHygRAAxJWs84xnD
Fo3OUUjQ5FvW2u/XfadZEMwdXIoDWyP3YLd+EtRDleYJvDg+mjNXGh1+xLV1PBkt
xbW5mPnKAmK/MPjgrsg9AQKFM/LzTP54xR6vRMHNzEDHIIM4yKTFNlCZcRRZvz3Z
iSIcx7Szvv53aFjKkP89TXNttoymP6FV9ZrRVoDU397nug6mETx1Uj87m6leTbWN
l8OnDzls9ur8WTe2HVinEbCfOa3wtUxZyrv24MsvoL/1cTn3f230fMcnCFWGhk9z
5Q5vkmdxI39cy9vq8nhnLsUFVU+I1Ls3r6mhychKuxkbFGiHjhVZPW5ncuvQh5C7
d/I76hSIRXKw4lMwzGNdQJO0hkO4AYCfnVi+t8FPGl1z1RemR5PdTB1z01rxJIiK
R6fQhc3IceW23NEtEmlsLvT1lNNIjPswN+Z+QYpr/EVN+l5RGYesKZ2rsdkQ8tcN
bWGIOYI8v0uzzBpf+TIDq5BZroKYkQrlDAgsr4YW6dxgQXBWCSiD0n7ftnkFgtFr
Rz76ySzc8ZX0ahucG3Nt5WWKb1NRC9y0bnquAcVMJPa3tQqTfBzBnZLk/gd6qil0
PK1vXXswYcdH9NIi0nR3vQyg/CvOBS1fMKPgAOd6MLGmIZ22+KysfdxO1n/bNdAG
5ooOmGZ2NVfx05XRb6GrawiPUhlR/hX1/rqfzL2sHGPaoWKpE4KpOUDWhcEM70UD
fVnsmoi1SEXMEucZ+Qnq/uZt9wqKJ+X66nQUCrDnXVyMfkxhak67DURGoJYRv0TW
2zk75T1anhI0aYS7SGnc1ZFuKRk2dS30kkgtN9lrXvNheEZKSPuOiy84ZFoBc35l
ckWQeu3Px0r15krDv1LB4qpy3nxrC2u+jPE/1QkeZ0Py7FkP0IfdsFpZZyioGC70
imKL+L0OtSvkz5PIr1Vt9T5rkSUSL5ycMCYw5ULPaQV091guM+LGD38z9b2fGQzC
itEb6pRC9flnEW16gKEeO2pipKfKTG3gWtipPQn8uHJLVLQc0MuunhWnP6Of4NUo
LDV3mRdeVPpGnZvtMXOhaW3ycknU6dE/4xGyaYOm8qWheGVrxM3iw6ECrgWtdOxL
FkWSiwkzmCasgK8ydgaiWE3NpwpFhmSYfAFZStYtt8zx6jkRdzzlc8C1rzxIQJuk
QeIILbgA/5C5oIrVaMEd5mCW9o3VePfODgsxDnko4u+V8PmU6az/teQw0/1gW7EK
sGeOg4fKC+zc+5B3HJaNy5a1zBhCpgi/mkcfYgX+cM2A3Z3OrTKy3Xt+Bbbxbs3+
EYpc3faJfxnRnaAM0OlzVBBJXiqIHjcp9OkSyTAhCr19ygPTSxSX2xwKXKZ9Ibg5
FKDdnH4FZnUqxVRiI36ei8TQ4vHotluyq+skRlqyGyIUnXxAiVNjpY04ccFk3Z39
vtJzXuxRwljI6dkWk7pdAzYCstGFB4vPGXzvzQ6gb4M5vD+qshptsFG3PKUrJ5KA
hfxg9lW/62zosKOMhe2eZYeXRPEZvDRLaEKF5z7qrIRyq8xd6Dmqddkoka6YoGIW
6PqBxCrVvRlKFp8WkPC3GqIvTxUWqFHkSm+IH+tucHhnBfMhtcxBJXr980OCbCRg
VsnpBLos0W6RPvAlajJsYLYhV/lpnJNtnLPdyiSL6xxDACGdKfkvBXg02vdgQcd6
74X+UrVS3/5MLUtgb+Yj3vVE2fN3hDLccmJyUI5mQhKaaHz/h3zVL4U89KsHImyx
hGEmyVxeO2zSwfy+i6OC+TJIPSc7fc3DRbBKNh5IZIknVZilS5zJAMISOL1dnGOA
u4KstETfaPpoCPpwdhYsJFnk9NSaFtPfL4AAbPlNBnZBQLIi5AQ6arVjb0ywD355
03y2EVzIsV8rTABrAgtN8JPfbsvCOcr13aEDWOSuffaKCRfoZDNR9YeZ7KEKX7Vs
UxRs6CMf2AnzX1h6DJbgzmRre+FTu71umQv13f7cvfkq6hNwfnSn11nHHwXpEEkN
86pkXrPgu3HgtfYdyTKgdGlahr7L5mieS4TeCMWwBcxm/xL3JSiNA8c+XgEGi6p6
NobzZbh4u1iECtfCoLmRyZeSqlyShI2Vc0mvBe5QOscyiYx2Vb8javpurxQE10Pb
AiXVvATfdqEN/muxJ9INLiKq6YG2RXaJnBqwmB881ScDuCH5bmVIVB5ETaeByczz
CihrHk3+yetaj1iBWxMKU1bcm2gOUT4MxRaDEvq/BGQM7wdYygWe6/KKScJQg8ds
7RF1C7t+6NlzSIpSJa7fJ4/aCYVfutxevoynCmroym4lQa61xsWrMVXMwkbkxtwS
YrHwa3DZXbTRqY3F+0DbI0OF3eXw/56NtEqqV1dOyTSJRcWNF/MYxqOk2DNw50IF
7+M8i2B4qbY9/GqBlU95ldXZtBPRjVmEmuNTWKYoa9WQvunWhcHCdAw+IUaoJp8n
6BeK55OrMdyaDQ6R8Byzh63ApzfAppjkQ1AyH195oLAWp5PZuxR1VD3y2ke7zN1g
AJG0MVGIu42skTVcDgYOyI7gac13Ojiyk9eUGyOPpm20a3HOpm7TyUVPkyi1WvZx
r/mOi7F43LYg9WNp0k8u7lFEVVzL8jGGyQSjMkJ64p2sjnahA3uqenQ45oKAjGfO
TvZTJGCYl0/1zbn/WB3s6JpKtmTkxBxuSxnkwFZlLu27Tq3fmROo1W81bZhsxbOM
WJD6fKn/yYxyJNIZ8ru/LKPfcgGfMvVJ9EVRgT3uh2jC19n3OfMV3lkHnsMq7pTo
hroTOU4ibd09Yg9xm+OuWG4O2QXmdrTF+DI8gM1UmoeSKRYWUaHOjURagtMu3SK7
jQGlPE1tR8XOUzXml8gGN4rgR7A6N2KEeZ3C5wwDkr52o244+Mx//XqqWd+4PPo4
QF0f3197FLgby18wkTHTOMIvRRGd3aCFYuoIvBZQewrz9/1111DyO59Nh49wVGaM
cvubqUJUj+nlrRZp6ro5Y57Eob9qZPyK3kG1ma3nvjViuwQZpdb0qR0pDOlHbYeG
ju7Z/6g2I3o/f7/d8M6TVZS332jfnR+QyjYY+R6XRnVrbjliyjUHxnrwdPNLCwvN
gIbDvOLrPSPN2pH2CmMKNjjeO1rNVqslhpoQQQupxYHZLxmdvYmsi9mzDK/FaxEi
KykJMvuQdVo+Irn3EkE6OagnsFDYGyrmd1MGlZCDaUxLiphKkGVXI8CV2XDpIxVG
zEAPJqbTIRDDIMJ7LdwaxaSyynfwlG3kubZ+EDurk0UGUGz6zjE/s8ZpPCEBLWwf
yPBmDzRVRM09cjHdTrtSaO+aSTwu2baJLYtFL1LnlBMvs/fHrUtN+pTb5/lWbM1a
Ld4loviaSQxYKTAiOqgCgSh1kzreAh+dp9Ti46b+eN+aUvpYAVfW/F6UQjqpcuEt
IZQlT4JKbL0o8r1wHzTde+dPJ03dvNDmC41/R9Knpp9JT70FoM2gvDa5Vwxi14+C
23PUYqmfvW4H8kDFixYsy2XB9858esnlvBtqlY5/ron44HRIt2PcH6N88gb5hmd4
FxH+73rt64VGsCq4zUhrOg5xC32v2M2i5DBmgPGGXm71Kr+dUxiDM2Q7Qo/CrgIH
lASWQa9cm0scU7C0ecFMLLLUz3pYGHJfs66YHYM9JTn3gwdi/k652VlWh2bEPbE4
Lzv1IN7u+BEICGeJa9KMQRMmRxsPdUPCKkE+yfd+ZmcqSTAQJQcTD4ObcHNqJRrU
yeEOCFlS/BqZXBjCZ75eyrBQsENNCTP5BjBxwIvn0OdKAZg0OoK1PmK1ByOikyaQ
mTfdq9/0TwZFbQ6geNhozqglovSI9mAiUIlhqWGWHzZ3dfcJ4c6t0KLzDp7dzr7u
b9VTg7WkI870gqB+ViV9gV3C4DpuyeQJlFiB3626HbrjzpfzOea/49ZScDs4vyIg
PkFevILN7j4bbAVT0JCeLSawiqNtwcXqBSXudbS6hJCOuLVu/HA4fqOPFK+hOAdD
bFHAJjkVWZ1ihPZVm+2Z1d3ZGRpXGYfKB8hKnYt3AajDr6LBUU5GGUYFY6a+wWeg
LIZ7K900JZ+8gyPxMrRdbuPGutCRL7wMxM9sXnDE7GP5ogWH9k/6zuYyr/RvxjUS
+rx41XjxHb+5IV3uzpo33EXCnaTqpGKT7oBnofnHMYKebPbaH4bRlmdTkjaNUCwc
f49rw3aCQmB/M+V5POWpbOiMgHccLoxaBzviZIprmjg0D7Cw1zR/Pu05fN5y+mjB
02kJ1fD1WtnozSZ+c1VM83J0pBUArB+28xK0lT1OF/VXvEPjuc3DYNmUcLX4xhRt
8woDwtL7WefkEle09TANZUZyo+/EFxynm/XKVDiqIehwiWSsBAH3y0Zo27ViwsIx
4lWMJpC7z6tsfnqD/c7hXKtO8UBlXHDwEOgY8ScE1u/5UMYqVkV3SPT0ILp6XO36
CkOLTTB3tR+v/x71eZk1Mov3qzVGiZ3EI2Ra/CEQUMkLlqVHct0bPkvW9tCcctDW
aGpZoXjvZKT96o+mHcyTnxHLDtY+jYtTVtKsLn0/HhYZ7iQhrag9QXwdVqfbBsOj
jaKINIPtBJE2AbdsVocm/GgeCYYvZEnccBj/X0OPGwvHqeGJUV+7nh5oaw7winrq
lIur5TO3J2XqDZ+W4GlZMAKDye4CsvKpqjgU77Bntq1CyjnEsUJtWzfJfxILTBkR
bzoqxBk1WUTUMfL2Ucx6mhzYIOKsW/ZNW/QoefzKV41M8hKwk1yhD6JIY7MKQt7S
+RxzTapYdHpEhpNr2hoHMkB2phWJDcIiThv8zRmUKboLC9k12EH66IPjTVQuAw+/
wTpGHkJ5ylewOpsMxypYsivG8uMQXayQgQXvEm6+BzRfniUQlVHI+Zw+sqsSjhxw
/rXflZbDfitlJ772SNRlIWDJJPSVVZAQRSlDirP/ccxJBaliehfqaYS0qQ2LgxQ7
2e+PagbkT1UQyE3H/7iABbKe6nPywOmOmjOiOkgxXEZt9gizUVFVSyazLqwhUMsO
34LTW8Uj9S9QhpTwz3K4q8BZ9ZFozLGZc2vjp7sWtOC9eS1kCB2++K8ZUKlft1L+
XuEoJxA/eEBW9cR3t3pTQ7n2OhsfKfJaomo23YrDoqV3BvjamMYHfVhxTg6c1cSC
PNe0F977yEzXF2pL7u55dMsVl994155VvUrkySXLFWxIx4OVUpodZ0CAKDmm0Rdw
7TD2hHjJUAqcSLu5/V80zOsYpjXqnkkd6y/WFoHZQf7cPjx6QGEkln9Lw0Nl1LAv
P6Ggt/3h2otynaTNZepvxcUOmBHuPXJoxxYa7S+lZkx0C06i1+iuHa7VqocaV5HO
MsEiglL2b+AORdI11M1df9y1lPPP511/XINEk2yevtZcaWI1ryMNbcWrqMlXAALv
LbluRtcVrTz64nLfIN9TP9dSMH40eww7YEUwwcyjc1hWu9fU4MYX1B3anbFdA64x
gaKHSlnB/Cpc7xcWpIRS4d2tvAQIJXXePGcm+RHcg7g1ghhHKXrg/CmKaq430xlH
CqxFyzgh1RSio01oo6VlVv8tgWrdqpN4aL5b2qIAp7QpLaqFg9gsb/OMFdob9B5S
f60Rr+2iKahFdcEhiyQQ0M8+i6HuHf3aYVPo9ZxL9LxcteDg2jX0XRLbInVXzrtE
267r69qYXil2Ozdg+ABVojiSVx2wRF+Ah1tJTzo/AIaKcQ9vXj4BG9jWPEUl6ot9
7aYkvZ/ld59GWTS6CHSw1QNUndjkzIqI0K01354oVTxDPdEW3p4EOCkS0R+m4z8N
EzffPjOFdYHSRP/En0b9X9tiNrRayv3swQQPDfFm34zEfh4UK9Sc889ZrKSu/W3c
SHZCumV+vIE963gajaKXNrIz6HrHvFnWCrURAaD8DKIfzjN4r5kdLijEyoeLA1cg
ct7w1e+2aQO/jUlBW+M4CYmPFJeMDDKmYgbhHPmCv09RgDgBfZbUXhB3GUQNQTA+
MMfWA/hUIp/47SHJLFgbmithQblvDMUJVkkcI5omIu5iHlwgcKmmuEKQiAShgUUg
Nd3Z4u7DBPib0/ZkMY0fzWSqmYF24zElL0rUy163c5Pxa1c/sA7qnmj4GD4YtX5s
w1zCxU/77bCwpBT6jjQwlnpA49srfmdzbMbkKV/dP/qwen9FzNbnDDssOWq1i8vH
TTZ3Wm60Bqstv00jF5jrMBMoN6K1Up5qECMQB0k5baRX1Uu53wsE+DzHXx3umkP2
p+B9loc9kCy+rij9bjwYKwTIGyYPqm4lTXzvaijRfSVDk+tgYFyAFlNrvdjEJoGX
NRixVPeO+rRnQcn6intgQfjONDpCkOnylkZSksF8Bd1Xbh5lu+gJf5tcPzJ4E9PM
Q7GGLrVaw6XjXTspzAqMGcujc3GXOi6QoXB+ZTz4op5qRJm/XBTbQTrgEAHMn+ym
gWniTIGwqnV2THFK4/e1Z9rwj0HKbrk7snrIIXdskLB3H9DRe42w0VdkNHw6s3WC
UJ6NaajysujJzuptvdQG3T/20S2VtXNO1nd4J3KLmitDFt1Bltf16nGToPR5YqPF
C/wKzwM2tDqv0Nqt8s6nNSd1/RmnzTGl09F37eiNSgYJCOPEuc1+zVYeYSXgCI1G
C8QxPqcffHMdL3haWGbu1VHzS9uVNYQSL548RjFm3+bZeJ/FDkXJpSwGWDFLNjEP
Fa3SyQCIjrOZz55wPO/HyxFsJhi4PdKv1os6OGRsgqqhhDx88aGvj+DmtJxwjzFV
Bw6DXfhALbg+48xWBR1F6JBy210Zmdu37ScNUiOLMJ1kI7QMsSVub0VEaaj60H2B
QvIThi/ShZFwwc4p2R7prL1+r25OnSmBWEIhr4STM/aDCLYN/fd2WL0ph07gmxaJ
Tv7WnDp3jr4uHHyWfpCbozn8+Pt3UUMxW5cBUaNOJWrohOBPPcfUa/HtvLDXy6gp
ohM2c7QmgYubdzcBz5hQxtb9T2/3t7pyN3po5IPnu2dH8YD8/h6Yu1sHZg123352
vTSARMo9RYVSlYMrzOTH+FwoKCyQ4+HP/+38YYJsdpLkj2rcl0POtCsSQj6ypTYS
NCbj5ZnRvZq6TmkarDBWiuC6q1WiZ/rscMvhSr06//hZ1BhOJZGTwz6pPJ+5VjJR
gdHtiL0MA6BGEr5tb5vwPVl3ZdKhMiPNlmpMiobmeLCB8g3Pd4ExY5jY6Tb60DjY
mqf1ujdUMkKXo547orGoc2aRHxdxFKPup5OauWuk5GbSMOwAWX/I4jkpAWeOFI/G
dlM75k18CpGxXY8YxpgEpQ3dTSd1RnGRrz4ZnoXCDBwLm92oxoNVUIBsXMV+qkvH
KluJsoM2oZ/N+aKsOSWKslxcCZOifJU1Nw5regeM5/YDa2c3TKBhYh97LctvscOw
On2NihgCeOUtIeU8u95ogKK6DGCqi0O2K7w9Azs/Zc/NIDNNfb/fCPRhpzSTMLT4
uXKOSfbxZ7Uz/kSYHjaD/dyP0j4b/Q4KG3z3BF6iEDi7bVCYYrN63PnCAe9nXgXF
blx6CBCUCpvySbTEWzkVhkX6bqe/UF5eaC8ucpQWxxFI6Iufff14eLi9rG9rm1nZ
c81YQDrkFuGko+9dsf+R/j4Fj4trOHfFWtBH+OrnTWYRa1tDZkKbIo96UfogKy1h
o/N5VpfNTac7FyR8NfELneBGvA32tWVXl17tAmb7zf6pJ6GyvxDEv2gcIky3VxAg
nya0zzhtCure8vhjFNgsdxSrHHH+jssVugHva2aT+8bXlTTr4YkqrpUJRRxZViB/
8sXYjVrUQfBjIAcZpOUFrp9ZIpG6V2EmBrumjI2ZkcH8c6FD5zf1OYay/Rn/Gvj1
7IDThFj+T1K6f2OPWrI96rYqQ9TYqr4yavYY4Vg7Rnj+SnPJwwCqhLfVSVJGcgoM
NSNkZxVKtblubMIwtUbvJIzGPgzOcez512XtuFKtBMy5fEdltQNYzD9+2Ab1EMHD
H5G19ANB8vhNGWy1RT+ZGSEn1cxFh5pvaWXq4w+JB2T7wDoe0WQjQ9EfmmMaA7y9
0Tgwfk7q7vOQyyoxsQQnhGNFXB7ATIHS0sNHWgwK65JTK9GQU8rK3+PZmi3g+JQ0
M41td1gT1zqMxIg7hHRcWdfUZ+A8aujOPK7QCu/qQWBi2wv93Sjt8ge4bmW/miBa
3KA68eiExqWI4CVjDL9E7w1Xc+g6TXA8aoQAOxBVxOQp3OucfHAFprEfCkrCvfgf
5f5MLaT6/QF10MDVvr6pShZDZll92ZRCosHqBE5CRn8sC4S6S9kdQ5HhhDsgWEBy
oMTYmlKOqvNRzdNZ8mhuoCzrNiCV6flZUyn3GK1lOZmdGtrmIJdd3a9iLzKWg0Rv
NeMlTBkFF2s8vNS9flMGWUNKhnxz0pZDhjvfjtTpPMwTr50HtvrvQURisLfWriW0
edCs3W4A+MvGAV8OsJqBIp8q/MyWh4l206i8MHCoGVBUJHotlwOxE4bfSB31BXl3
xPeD8Y2Z/KVgCHQDAhWXmzJnXz27u4r6aGXmdnfKuhopbW7T5UN9aYLbqhJEtHrU
YTFDDa3yW0KVZq1gZmAQ/1KduQsXNkbipXh8d2WZOFzG63KljERK60BdS0NQtCCi
JY1psTfIMHO6bpiCybAFNdeXPxNT+9/tuHfBHqMrmXiKXM5WS4FHnYWlmiLVf16d
bGBlQegf5+FChuTcu65IF+ax5udd0DpCSg4vQqe8n5bQzs79zNYk1Os8YPGT1/mk
jpLWkfd4sCZ3OJD67MTpjSNQC81qh10wQyqeB6g1faNKZYv4mHaVK3Na4NX7bdME
rDBMxTNsXOf8msgmkR0eysxBuATES6KdUI7pINxcaFvwdSpfZoofwmHSL2vAtTI0
x8hUhFdp3MgrpUDhZyx0DgY2e6livmUi+rOWXjxAfKdnlFTnpkoII198tSbNYR3k
Brkk4RRtkPfwnFiP9qxfJEK41sCMrIqbY8Qg4QtuUFHLXhXX5c42HtLGY/fu4HfS
V7c8q/oLurmUxyItto53MBSzX+fIi3hPVh3nwuYB4c+xmf02wKrsLEbvNMVkAYRx
TlWKzY7ELtws9djJ0pMQ3KfNN/DelNLtlMuepsvpKcQ6UhDAZ1hb+NwdKUucKXbf
fTCrXvoMZLbqsYZ+hBvNpfNldfjB9NdOjOP+oOYxjM1OUwMQYx/qPXyexIdimhmy
oj1Pz0+c6c9lxLrXMDbhCxYLm/tkDjMjOqHYGFKApWO04l+NaDu5RhS9rMYKjL8+
bQTxAg9txwYjdYLHRvUfFcLZJ0RewcyKGoafFHZymKDDIfgi0VC1ABB7QEn85XpF
SxgkQt5l/aLor84QYAdfxhIZVy99B6qF32mZMfOBgyTEwUVgec/oK5r9Mqnk4w8f
W5Wb1O+CE0oQ/88eotnm0rW4eXYk0u80OWgLrk55atrOQhUys5tFxL8yy6XoDqkF
rRchw6dTkhKLAZuKQX86XVQM7LYp2crZ9lttoHZ7WI1yAnBzRJQGrD6Z7KHPh1hv
YDwOi2lUgDUAr0wmzMtOUB2I+wh3X5HdLe2viPZvEbwMZ1pWnU+uGqbh1O2HkRD3
ffIazFBDpqgJ5U+y1PjzuSMfjCum4ZFBT4Qh09Cqb9MCQvZ/bcsDm80zy2BHmVFa
VZ1fo/H+aY4M/j/gaUFHWjRqXrrWjZdfJDRa0G9GqP6wenVFpJvvaQtL+IRL2R69
eN2ZyAFFxvC1ySQvmlhCCdItgiayDuVNFKn8sQLhUfuN9PQ8wlBfFV91BMzX3TZE
5dAJdVO5/F673/LQV6iRJ2vssUYbvBguyPhPmef51kD2UscldFNnlXWTilKqqkuk
V6kyaZw3VAG1z8u1MfHg3jvV6E8ttPo4we2rwdAejpM5SW7TeTC3Mm/OzXU+mjrq
JCoZhWANp9YQ9NHokULA3WF2EGtFV11FSahq0wsn80VGfVwo6inHWNv60ZL7A8Sa
e16Y7AcEhoZZrrSS0N0tBCLpmFAKMH3/Gx4OPuSgmJJQdMZajTnAkgWTEAKwhOCW
9rxES4M9I7zxqr0/EBEYwEf7dCZHcbNxsWzVm05IyAyj2rgY9aFOvpTvw4hvo9RX
7EjvJ2Q6EvASa4NPzsSffdsXN09LXrawnBEARoDbOGpfHtQyzgBMVbMdUHYhe6SZ
Gzp5M7OpsC9RjdKHWdjuvneSHiwve5kzfIoAYjeF/40U6ZRWkmvK5aSC837+DXtW
Ze0G3nHlSdomQPWAYdoutUYmWbmm37mqoi4e+ps65GRjvp0cn9+dwmUa6/R93Yd0
68EYP+11/gaEq0XsAyK08SSQ2m/Do/xuUA6BMeBiY4hHtKggDzkJvy30p1DRGrvf
kVKY4PutCUCdna2ijxGgu9MHl+27UNxsZkYCz6k/k8o97JfLYYAkw2WE/zgjdGSw
cE/EG0Cv2ChmpBBRSDqK28bpXqPc22iCVH4TUW79A1yDwa0OSPUnJ6kLIjt6gArm
t85c1xmHXkDlfgYdJ1mCCv1yYwa3XiUM6ggqM4GfGfAwhH//S+yoXEHWMeZi9ExB
FDLMowTmRrW7YyI1kvizT8J7og5R0A7gdykkWaI2d75/VPJOllTu0J0svXBDSeb1
nIgFedwoz8b8mCpyDu4WNKfOKCwqOknJDGqeKTvw6FMS4uKBp5hEcFK5fUKXgLak
fwjwsV8i4hpJQ/Ueqdu8yqd+JTgWHO2EPPW5t17n2pZEb2ZaxxjG9h8WrfU42dSE
PrU3XMb0qkneaPG0uLJoGSuegT5pUgDfINc2QY5YHG+xtMoK6ZiuLb14+FSsGjOB
g4cyE0pHo9PcyMBT/gvQD1tuQP95GwpK3kP9ZMhnU43cYH9XFhndfUGKzaPg5ZTS
Ta5Goo9NXVmnxeygKzJm2LS/3WF5QzQRjAPDVVjr68sNtIehGP+G5iCw0KCrNYJ2
vm4KwbsL5g9oqVdFD0+MueeGFtkw45QT6s9dhqVMGNxi4TZsqdMJeSXw0Ac2r4P+
i0aH1YX/TWCPS0vDpstpa6MMp2fT9LvlMwG+4Qu8Sng1wKRjT6kpS/lqxxW7Efmn
K01AOxSjCIjcNxrhlkGn3xNGoR8U1yZ+EOyspUtC8qZjCt1DlMbTYbzCpQqsVKxk
Yvn17fEtIyXEg4yH+Y+fMIgZ1ix95mUtrj5HCz5P8hgHubrieFNx+hFwpxO3azzB
UN1eOap804pRD9FA7cqOvcHcs+dAilflgzAO4bk5J3vfUBWsVfYGwxTNtQjOqVWp
JIQwm9ATPqj7eM5cdbYrNWRMPsvyi/jvQ48DFTKTPk4wPG+wYWBpKe4FYlbBzbHN
m2kD0dXH+L0qXLVAsLUeMCzapNPQINE/8bZWnybLxg4R9UvhxqoZt9kqvB8pudtu
Jd0XM/feU86Fa3ObQTD8tCQKAII38+xFiN5jkqbz8wwvj/FGZ1aWKxT5FmPb462Z
g/EtExTmkCKq4MkPZFO9fBWgsMYsBqzW/1OoSGYaRRAi9SpMwQpI7I0DkEAMvmTT
1iEyFEJUS9n7zdSCynBEPPGyfhAxAqKbXAvLE6HST5/GsQW/pwhVl0Jus7w4vc6a
8c2Stl8avwYS0XlsXUQKEh3R0m5Un5XN9BAzRlMkqBDSQKKgeAnFiuLJDx8qgF/9
5XzW1cfKcihPQfM4BDW6mR73G2Bf0AZ0dv/H/2CL6nZWuabgeqmFyvuyleU8Cf/h
Tp4IVtgH0dzGl1ZHnOKieTdnjRG8zBdT8BD7DXeBgy7v+YXkRahj9Bn7Vrt+pw+2
eRfV9kIUYb2KmkWu94HTCXmE1vthFBvZ4OBFLfmjHDboemC+Fos5ubdIEKJala32
UGBLad2+67TkcAEJ0imH3gUn/NVSF67MI8vn0/p2BWXNh8WB+SiK363v7PXxsNcE
jtZiC/SnGziXY2j3JGPrt/31bQdxMXfCXBabmv+jATRLmAWoUC/RpLG2HUJ/D6RZ
t7AUxmmgOp9bP9p9AwrQqMTlw36pE5kjob/2D219hPC1D9r/TSCWmkSDv2fuEk/O
SCBcNqbQ8PPmXoEc5lgpQ8jPkwiRCZTzBt3vB/nf/XOsR/kR/+DDuReGhSqy+fkz
NwejZNSeo824Jrc8WRgAVhyki0ZUMbWpNrEsVfzcR9EyU98z/DfH9IMvo8ZF5v57
StuKOhAfR9to7Lbfq5u8SDxSRk6hvcBbZJFK42fiadUgKbzu5x8UTwn0OS0ESWS2
FW8FLOnuHHakjlXSqwvS8zRb711pQpysKExGhTZ+mzWM3LpU55z/0y/+mNl33WaP
afPoNL8B25ZXCQdPjTRnrgKxDeiBLBqnPMUeKb+VuUszSggDBrO5sjAGFrL3tGvx
6ytrjIFNPpdtgh9Qa2WzebgV7g7dfrSO6WgqPhBZ3WuQ67NIsUJbvdPgL4AvDvqx
Bk6tHVYluKiq1ZZfQPJKjWohcXeyAcFlXYJ8kX/S632EeTi/g1gDY5pr8190dtfb
peULy/r40xd1rZ1PZg/cEjx7sbrbdBR0H1ajbFCSopTh1pQpbj3c8MDEn9mISamY
O665tTnvsMZpDCJuxq8ZoospOElOZFd8pjRfYf7U/1O6Lj+ZcAQV0ctbJnzJyPrp
bW0fJby95ycY6DJSN2fyrQ80qY2sJ8wHfOOOQzOBEu+BZOWKwIVc0dwQY+xVbQ0u
E8NVksP0/Drfk6le5TtXsC5F4h1eKeZzHBPV7v0PdoixVBRAAzOmu16jqYALVNou
1uwpWW5otMGBAUuuw8ABhT4Rku0WT6h+9BS/ND/8ZdyNKqinU6uTWZnAkn1K7Dwm
4j4SA8Ze8oRbu1jGrTAttf6evvJraXXVteqOkptOUT84Xf/l279AvhMrEPvE+vEc
Gd63W6jOSHezBcpqVbfLO/LdOdGhNDnZSr4geJGNbEvIbwgNvx6y/7OKFkVoyLO6
oyUxaHzBnFmISEQCycu/Q5nlnN6DLZO9egXEEzfzUJNopStVTwxd1TcJFhExQGd6
XRxqh7BiRY80Cn4Xr9voI2QTsG2HcIFwxEp+7O9XgjC5tTYcxrC1ARYY4WJj9WfW
Gj3c11Cpz/0x93kbzuU3UdlBxIQWsT50a8O57BuyDLR0Wwb856YYuTVL7Sx28Zxa
/YY/AbHS5L5pNlVjbShDL5bUK1idDvTxI/c6OEe1jeIXadLTQapl0UL9bM57FT2w
dcR/6aZTQRiT5qANhGBimRG+1mvDT04W+yUFrLYo007/TCIE8GSc9uiWUf5VJIP9
PrP5YRMUhFgYFmzlmLDQZp4E/+1HvpXso133pMCZ7bD5mUgP3LhCDwjzaooAXFAU
ii3rArz1vjJ24TuANVtAB6ZckOlj2uj2NSl7iSCHdaxLaWjxrbZsl3MU571DRHIC
4q2yqlXdwwUpcNpmkHRFTJrSh/eNoG8BZq47siIovY+6L0/4Wecwz19D8P6bMukG
OC/RXOmlFE8KXI8czX/yLLO37xtcd1CqMck7G9psPPX3jVkflS1L0zu5v5Gy/Kr7
SyB3AcGlcR6rfHXTghsm2TAZ3yscA295A43apHO+l+49oZxZONEwdEFCGzxdHkWg
uUFqMLqnmFPwxBLNkQHtebMDX4sWRK0Wc+3URy68jjpEpN+UIPjDIRmwPcGDtXpA
EQkDrXaKYr/lTpGlLtHeMPcnNKbOWlMqNOAaFkmT/6Ww6otOPoJB2T5gWWnKch7g
JexoOFbC8/Fvz5lOVRJWuXQx+zh9OvUuvdiIce9ewX6Tq9CZoPdKW38CoY3RGg6L
GVDVF1dqfow8ETg5Ml+uqeAh5KV1E6s9DGYU7zOcuhZy6yzkREpdsRLuAyQQPOXy
xZIUIA1mbgwf3Br8MGEoe07GqygnX6ReOUAOEoxtOW6PlpY5k6BQNgNx0JmZYMYO
Zd+Wfzf8DJvBOm3X95iu6IeYVN+XV0H150zNBusgTJ7uly26oJvyQy4YHfLoSl0z
Ya5hR/PS2WxKpr8FmaLtYvC5mt9KwPn1Q9qOa7XHpWugf/hBulLjhXl0ZI/fdnkp
GW+fvFEsjvREVL7zovLyLvdTW1+VUxQGGY8+eF6N+JN5S/2LUejjBGQPNtZbpkjW
wG1sFqMKO7YIgKqUyY+xMp6bW9DJlfdopce+v3dmJGKQlSklBmsvK3J0s1NPE0bk
ww0nHFkF9hLegenLYrD+Rq+IdyADOV828kznEZUQ6jlcJwPIJvxjDWRr1P4pcgwK
1JQpOpiqTp0xU9gzbGohZW56Gkx22IMTeyggW+AK7tEtuQ5rJ5p6ZFlHdUFXEtad
fcOzkwkWtuWtS+oY1YpQGtIWM6V+IrMj1nJsq5G3CLYYP8LqK4f/zTruEzhhiFio
QBHrTtk2wzEdta+bmSiha6ithoMgCq4JBWjTVEDDCXebAJL8u1CaEIUziP+Ojz8q
C/ZrXn/RK4MTXqhSitwdyx3oHuKpqWD9Bwv2E7jSh8RP+PEkAOaH2d02RjfB7uaN
JTpQ8PNr8ldp81mnaW7N77Cpz56iOnOdEww58k4AoqCc88o7xr3afLpjIdkbXMoS
SZi3+2Ve17Cv5GJPJ/0ttC0MVrlG2TfKugJYuatrhhB98b6JbM1Nt/01o9YoIMyR
Uah7s+laJdjZKVPr6qCZRxm3J0wFjdPIlUvSt0/yf/PzrUDqHgyv9TRhE6tbIudK
6VsB6Z0gt4qufikFR+8DfoHzm5ZFvquk8qYNP26ZMuE2wOuteaqY4ZlntCMgbYUQ
4u4dpxz57xnc/IikHNTPKkn513n51SheLF8pHCd9xvjT9S5qGXglz0T1RhJCzjbA
vZVm8yXLtME1elJTHAuVeSTT8A9FodM51pNYsjiw5jUpkTwFUEriEvJBBD8eLv4+
6abMJEa7cJjgPO6Z9bN5N8ZDFczBD4OrRAclZh3YagZdlLj9iBJY2xUw71IgqT36
1jUEYec8iF4Ws0B0pMcdIxu1oCywUedMtpEyzHYyPKCMOR8Ue/ZvnZMS+GRXzL/t
palH4kHdOyj6WgFn7/cNv4md4X53z3wnuX/rsOrN14kgt6GK0MDPb6688+88jiK1
oIAzQIyeYjyE57PHSgOJ7c3mY1qGru+hwFdZ8LHYYfzBvQSfDQPRkjLTiZHvFxMZ
5DthqTBa+RB8M/qH8FkzWGBa1jj/cCXcBD8jSuhjsosb0X33VMIV5oYhHdML34V1
DKFhM5CPuSq9zPDIVQS9Oag9uYr6JeXTl0DTJdLcM5pgxejHzQkp6E2pdddv9bUE
vdvFAyRtS4Cp2SEA34z1SkIQf28sjCYAt4UAmrrE/TxVhYZMOIyk1TeOyQZEHFf/
O//9ElWSbvezeSy3mLegRlPqL7I8TH3HKf3PjJHfO5cdKa6VXl42ZIVlzr9F3MjP
eGYgyhVcGPsHX/pBPy6m7QvRHPifbAxW0WjwrhG8AulWu2OvJ+O+mCiZ7oObtHmn
JF+s4H42XEvj5Wllk1KGzr89zDunabiz6MHpvSMEypZM1VmXGG7ni9n+A33iBSwu
0yn+ZwTHyZqvBmgS/S3uBMk3FB4eY7xXHiVMHr4pU7VVbJMKqU9HZWpmAoRc03IN
w8P4usLyFfy9ADM2WlU33khO8d+uIBNDjIVdFVxCQ809Un51cQg77fNSoiAqU9Nz
lt9x5vOoZFK5h5g//k2g+vxisREYfmd7YJDwzVYkSztH2JvQ3iEr+ndg1y211QFB
T98tXWF4x+MMKZUgVm0w0WEoxSXFRFRvhtLDtms9HYWKcjOutuGw2GM5ZXuHwXYI
I0V2DTDOOrtVDLsbF2dpbufkhy5ludHxj+hstOrh62kgcfN1+gLFfllKv3NbqBkH
O8Dh8NNYPwqkDGmj+NYJWUBwYNQVmrUCyPuzuf2t4Zha75UPaB/InC1Gj/UpolSX
4yENPML1WxCmCKbQpRtEIflfIf8b/1vCwP9bAzVrC+Z7YcI14bF06nL6ky/+ATtP
PISwKea0c7E7DRHFIUYbk4bekzQhBXFyFaXhleZIh/kA0TubRT896HrcF6JBV01U
88Y56Md1HZucXBwohydxkuanOXWkM9s1/3HteWpvZm6eXtCicYLzF2jG8OCKzAFZ
hWprDbEV8twwlrSUyujzagQ+gc8qVurbe36C112qZdcoCyXoGfnFJgvgyrqJJbps
kldWBe76LGQaJjLWhdzGd75KxEj+pi9DyZCvBscvh38SIVOEtWDNleTManWTafYy
NHpw6La7WNvnHQ/wBoWKMA5g92s5nH+MZPG4n4LPrZWDUpkpYN4zwi5PtP9uRsOm
sP3Loa9QbvRcZ2AnhLaZwdbV2mY3c9CCHzxFPy+u98QFKCahOCa5UlYPM+EsmhRQ
lUfiiVdijAph/RyKgTfCBYP+KTbuP6OJaswTHAnruIp3N4/2+rb7ojsIdR7t+VQ9
79OmkGywFd/nXySZ2Brcow0ilnnLWRqJeGZ2HnD/EkBTiV2BXFHexRq5JU4Eeu32
/RjVxFUuiBbsohk2c0VGrw6brmJErfyc+8/zrJ1iOeSzMNwrQ0/TVn1uSuhwFpvo
AwRgohp5j6ulteG2e+JoAZ84kjuDISHj1otuug91TIld+8awVTZiv0ZOgsmYE/5d
Pl/GJ89SztXW86rj/GV4IknLQu2fRGcElV9R+kshIJgzVs5ejcbNGpVgp5aBbYQc
1lyXcYrkbli/tNeNJmNLFg5fWjHxgtOP7YkBKoAG+1Jsx7YgOkgW42je/OXHOgvf
hRPz6MgrCLqzo+QPLb0aYqOml92X0s+cNFSCf1j5A0GvIlVHOzV5Z0MLvZImg5n2
jGBKX40qh04nXqFaEvr6q7K6+X4R04ty35m2xO2Vv8tFKqXBLCApu2zlFZkDnjMh
ZIvHkgMMsFpmWeCmIJP6FIp2bg8oAc61piuNOLQvBze71dvuGXmevXx2WeddLGt9
lN5aquw9+ujt2zyTkwou+g0VNBHiWiCU8s2uibnjxZtYb+mOMa1Q16fLA4lspVrU
4rtwghNWeyWyPRXaoBDPQZj/Prxuw3or018IiuQh/cj02aA1B2V0H95vB2z2KDT9
z54FNBIJ8+1hyGpSLSEY02jf1QRIrbUvirLZmn+QW5/CGj3eCRz1XFw+zkq0wkKS
ajNIidfMQ/vWQuayO91LQ9sUJEpKz6gXkNQvVVQcjTRodlxSCGlhWYrQq9teV8Yn
X23FRUofmjFrWLFBHPfRsHH4oS14jd9KDCBpVoN7YzHKMYti0fSayNXaaRKwt/d1
E0UJT9qsLAENmhH/q00Jwb0cCNj2E2/Fbf33434pIS/VSODW9vWLPTdymn99uP/G
qU+E9cuV04FDaCgIyrnah1utyN4Ad9ftLFym48Bdh6o5ishL2acZ5rYU/uQ8Zskh
8M0EKTxwYZtYmyBjh0XC1ZpjOje177O31gocfYyGvBVqny4m0c91XufUZIuui2Rn
Qs6G0u/EgY+HuJZdTFhUMLJh2wdX0uOh8FFhW2k/CD2+itUtJtkCo8qSRBNUakGP
tyi4zltp8MoCj+tRxo5R2KQWXWsY/npgj0qTaipumS1MviwRRE3lTsD/DOvnegaf
6HAcalSxd8LSmY92gbaDyR3KJX4U6LGqnStivhJaRJnzpyRad9yAyD2K8FjoZK1j
KgNOZpdqy0V9xODAZd55nC0uV/UjfoXmR292zHpAwIURUXTJo4N+nY0OMBtvy8WL
aXmR6kWMubUbmoze0aiYslvj8GiGP5zoTcSov3dN4poRKl/9s4i5B5e+bhlN/Rx7
mC2XzVnISsr2d1HnK2F8RhhSeNXlTpj7I7HXhPPl/4RkCs5MTZ6JhlLteIJeK2AW
rvs1e6MBgQRv0W6P8gcxIH8BkAl4FVhJhV1JI6TGvXHQ+uaekvi+nsYSrXjWpZJc
U8CiNxq+cs8FLkF/c6mkfOizD1m5+jaTW/uTaIm6RkJbutT00hJIHtkiHMMXnfno
VOg2K7zttt1hAtsPU+3VfBhM47CeAuAYmBeluZr2oIhL1tPampc+tsv9XlCu9ZRZ
+b4ozT8Pocx/sXGTEBjqQZZT1EnXhnhGyDUJSM1ASElyycycaWwQiK7gLres+ozR
5GmXX2rEaaKguuFlu5oYzcNoCIUpA3h3Q3wgLRonVyKwIlGvHIxwUX6JdzUrb/Qv
nKpTTQi1yaqol1nAqQQgXYfVcT1GbXeMsFtXqajbsREqu7904t2RCK039rn8lv8t
LGSdV3aeGia8E2sbLfVBPfZVGi1sS1jhsZPoQGLeG+A8cNZoDB26nMI4+tKLdhbK
M1VDE0EamfU5e3vpFmm1EQfYsHJMvAzgez5vgatHpoPHM0hXCeVk0hOcM8MYu4ir
CKnOrGOEtI/JHq/yGKliQjkZdtlkYkeUqOHIniMv3X0SX0VPPNxNDttayULIFuE3
veBkXFpzqiRyLBymXyPnU+5ohaFgMQLjg8skEuegbMhq4FfP5s5fgdBKW2Ouuo+5
XQFQK6jHdgjtSbe6Bh00iqD5h9jezvhy9zVuHRmnqn6cyXADRDj9J/oA88ERVdT+
E4qnEWsJlyu2lfT//C/n3CvC8LeEyQzSkQNGkoiMaP9VZCgovTKdGMj//LQQRK/k
Cke8RsQL01553d7N1pRbmZK1G34C+GmYLklHRgGA+Tzs+ciekHnFoMm0g+cRGSjC
dgv47Er52w2TAUretZErnZ5ypIH8HmcViANJsvStAX1ChY8rCW8t4p0c4vlNgC6D
zmxgwHNhTjvS0G1udstD6H1H1VmfYYd370fXBI1BaA49YPq9qrk9V6jThZl3f6rd
+g0SbQ9GDYbgFAQbqWSjv35X+Ciz6I/GdiQDkoaRXLs+NwFmGx7kuTK25wUJQ8ol
1tzbaLXdo/YB8Fzpyp8HBMM0N97NckWemudhpHBlpZWSgEunl2IyH2MpyFw5k/dk
t7WaB4YrjRgfRk3h1abdzU9K+w4V6e10cXDwPEA112Lhlz5imcX1yKJguRzavkbs
2+E6XxxTJ9JmwIJO+Urg+ccVjs3la5icaJ6FEVAqm7MJ6jYVuAIp15im5YEE9fNt
aFuaLh2wKEOBs6zsQl3tZ895GGhcvW3fVebowQWOawNa4+KQx30YipCZGZTworCS
qO22Dsyh/KSGB86XKNASg1LdiONHN8z6dqeFn8XOFfs1eZ/CivNyp9DnjxIV2Cnx
A2XXmoprKlg/gOyh3AWO5UIJHPEow2qXNC5Oa6VfQQJd2tec0l2DlMP6TfOlxJKc
2J2GwEdVcTtWbtEQ5kYCiiy47/oY6wKOVxXdiwmfKzJHMnCjcQeQ26BilRP/rML/
PuGmb67koSO8CHjovTYjZ22Tm3CIoK7T2gRyDXrDLvvdbrdIntlesw4vNZNbadPk
63aNREcjq3Bp6TyHAw7zrenARp9h1fzMdz8PVs1kFl5KnYJhv2zfx2FAzG46c3gG
ahzVP9lFni8A6rxQfxBEiGtGNWdHO3eE5owfiHxPY1iSN0ORKQU3LZuneVm9rPyC
a5a/P9q+v4OKqOYy0KaiAUqOQ6u/xCQFgrb5ZzrS8sDJrgPIho7GkGoSuzpm0z+Q
+D510uEtQ8BgQFtTodEfujZqB4nYTyymLX7h8+sSQsAfIQe3FXp4WM5kmNCirNum
YZEFFAzqR9W8nBYCbGOCU3KHbZZ7R4S2yvdxrmo1r3+3e0eqHnHeaAqWENI2fs7B
z9qu605SonCIvKBL/6FjOc9roCY4WM7L/+uIjBwy/kcMJpUzjXPf7m1S0tiSfdss
8yawAtF9Ou0mISUGvd2Eism54W8tEg0ZVWFKviT6T8DAAZYCocYkQ/e6IojSrFxQ
b5oHuehz7db41k/BsAQfyU3hkU6Av+PqvovhCJz+E1zRiGCUNPfZ4qQ6OzdnFq9D
N3NZeaC9iol8xkPnL4m0nkZ67awg3wdg7RUh0iaO8NU=
`protect END_PROTECTED
