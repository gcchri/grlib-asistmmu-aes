`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+tWpPgGaDt1oGgWAmRO7Rby/If7vpWRUd+627SDOezV3n9BDpk8/fiuLMWcmyMy/
Un0/Yv/txGzVevY1Au9oISZkV1a1RGSKB6lpesqlW7MPCVuChUDQak19VsQyFpxR
p7OXjQJcN+L7+dXpYkUITO6fh+q55zKg2uwKQMmASboEd46IxJR3thParSlCPnM4
IRGAomboBhThnNI+pak8ZNy+IbzndhLJoWtA3Z8LpRrXsQhz81R/UzcmT5KJLnHW
p5ikMnwk2JiirleTMYx8zfSF7igaKR736t6OeXqk7HBCkLFFGs1wEZrUr71FxrUI
95IAK0DCswyrHomFqVA6jQTSGkX4AptrtZPH8oL5+5GM6E8h7+TKyOLeFr4BTbb5
KUg6INKpGqEE9KUiHFvFUXnR0fZHebhyDkZeDoShW5ZT8Fa5tU9RG3lim/sabNfm
dXPL/tjgztjukvv43FFDUJb2fLVX/u7B5xl3lQE7Lk793AtK21DGocxN2rxdn3Kr
00EUW2L30WNahsQrKDfvtCJW8TkZ3f4Jj1yXiIrjWs7IRsECozp6XltCQeGaB8v6
89MsZoiW5F6MUERZDxRBOA==
`protect END_PROTECTED
