`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B8gMThEk0VJd0LWKiKBnO+FRxVuz4DGyHCy1yxSfbBt+zpeqmmgFEvQQjT0KOkwd
xBSK7E8qfxvrJCR/R9PUwXj0gnOYWY3TygOfPCpkvRCga3GhNh2CB6JgiKp4JTwA
MXLh0QVA9MexDLrDQv/SlkjJEsEzLPPC/1Cw7r+96R2fZfvtsQN/hXSwitsB1KZ9
t/Hp9yigBCL26uELhW2L9PGDRACuHbitKDOTHrL7l16tqVL5saJfp9TkNpWX6ImC
XaYciCaei83pfXuFh3Fre7I8yHyKcFKmJXVnv2JQo3uMH0FOqXA1ipGOy91ozoma
+NcDisVTAE5QMXt0/jwK36oKP4ksXpyFiPOL4SUvASMI6VQ02G5NmMQvzM23D4r1
9rekdMzeMR1xe2xrEJ5DgqZLU52huwuNQFjRa/4zs7QafOZ0u0qcYhSwuLYFlOkC
DwQArr6NhFGCsgESAfFSimNOVrmSpivLKBOKUjq515/dDbRATkL4QNveYemWri9h
FnIPMHTyyC2r8stAPZcOhQ==
`protect END_PROTECTED
