`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6MzdFoUBM/Ig68XJgoXI1fEJVx3u+t8CYR8UFTNCc/h5oDQKs0bARkYGCeVazqB5
5LlEvonaTxISQV/mBJ8p2U5O7r+Jz8vu2zGgwVPw76iXETyN+jo+QhAvqAhBeT8C
ZotwI/mSyI+wTe+TV7ya2HDa5IIWG/PCqLFFSx6Hz0ewSiNVwOU2xN3SLckYaXDL
b3MQpVgGlQ0MyuHBJRC0oraeoecsxqU3hUsnGcIxEhcBhDMYabd1QOjpmCyUPLSL
9KqeL6YYn+L710FCR/ImMUvs23jrbMVzfJrGBzK3pYxFcec3NUGO3tzysgRVFVtu
4iMxVtu4leQn8Nu1imPhY1WmTRwWiambbtbOKItvacJK38zBAEDIX3SHP36zwdDM
G0Qy8Ns9sh8+FxUPbCic9dQVGGgN1xd2DBJ8c9EpJnlO+XN48elYzmykHu/1R1JZ
EyLBkA9/Jn1MDJEifEtNpGhqAwc+gDGS8PVixLAqFirvCiVYAPJidWxe56S48Jhi
MsH+xVUGxbSxtPKWT89OGX/Pvy3TEpJoe17StGGpSiSJti0L8hEtJAPaj+Q72i1B
O6ad9qAl3N+NHTkq4QZbXUMr8YEXtRNIPBw848zJIv+T7c74tl4aeFnDpifo/CBU
xi7mJx65pRoFPssj2Iwl43MJnICuHRqwR3sp0wC+d9FA5z/VIVy+lW3y8TlPqRLv
efIM1gohHWScL0JjWUOaZg==
`protect END_PROTECTED
