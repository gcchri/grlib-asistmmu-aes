`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LoxlLAQC3mVXA+I3h4rkdJJZ+hViswzDmPn870J4l8Azg0xMahg4a3RYMRXIK1Kh
swapRtAKZxkILyRLXxx33d36pw/2v9mVdY3vhcLsj63bg0g7G3uyEx7aeHgWE5/w
/9vY+zja+RfDNM6+SplZfUj4Y1/k8FZIpeYjnpy9kTOnw9/OCnDwQqyWaYp5/28I
LrEKzxDZWPnQ2tIAIouxxpncHgZ+2sTTWpVdw5aSJIb1rPGcx1XPMc8mYl1TbC/J
tmVOGzY5Qoi1CsJSkWtHQx4PeD4UD5U5Erib3dNeBIiRZ6LnyCsEDJYA6nu1LPik
YePZJ4sG4k90N35fwnYeoVmCBnBmzHEfVg+/GDBAFDpkmBxEGnHQb4X9eCOVNHZa
k8pM/0uTR7LqYa7HhvEX7HInsK5T6WdkR4UoUUvGF5ebZBJ+XtEJxuRHbOEekT1C
HFlA0XAOvpikV76g6RQMbphdW9FnvZ9I9ZXdW3htdKRd3cBIjLvBOqpZR7anVRXJ
9crShaEIk0GkzXf/S7tZDsVvVjik5pQyJpqDekUVPCuQ1JBPqVaSljb2do+xOAR/
skzyWqBr+NndO2EAiPHR1x++deo7bpysiLS69s99sNFfDvVIVjYjts8/B8pkEKzm
MC9XRcjT4IwRy55zcrXxluCRhyhDf25p8gh6odK3svIqQvMKMH1Ep65HBeK6LHoW
DvTNja/GQH7GpW5/YxSlChbUwMfiAvH2UyrP3oIKMehNfW8MFJP0Vby6t7RbWBPg
DPPBc43oIB/Pvk8PsOUve2NUsPFRYey98m+sXbWYR4zQq9KrlxuRimk7ozj9Xugo
+df4/Xn6A9tGpfV8hm/HqNw2jUkQCA9fzRhTDvDu61YRJC7wFfzoSG0NWlh7E1fv
UEMLim1y2Jxra8N5thg5UaeGz+FiSnSiaftPDk/DNFcc+nU2sEopeVXLo6lC96qd
Eg3QK9lxcrc+SDjLh2EBoq0FFXTNd19MhoREt5urKmoucZZyJcAid+BUoQTqfEGs
abKMyd/WjsVdluvaliRzY+HwIjrdRE/AVk+xJuvgPWkWYaygat81CbQUsitF0fpt
BOgNd6Rwy9fyq4dKrx55X4JWFQIUIwNvx0/MZtx3NuDqn2BfMl9vx9aITP+jjLmZ
biG7TWaMjszOXO20XA7AWiF0UrdAgt0VGKpPOpoeAZ/egP6qedjmmPevhF/gRNxA
lNNHInvx4JOwXHer6bTH7tX94M9cFN8BO3bwF0YVTzy7drihTnYJRMc0+jeDXeg8
pK+Z7rIhZ4z71xXDiaX2Yg6C4Mp3uCRJenf/vNvFRvqAbt7T2MQXWi8QzBkvl3y5
o9ifeYnbkxiPx/0ptPungNksMDnl1IrSTpZgkxFscwlcNkBiJSlloEc/HUtyduV8
eQ0x2p9Ml70nTbnSR9TAFGHHpnhFMW3SDaIV0UHYQbnEUsYyRH5dB7nwQPJXTxD3
MZfNYdn9vXoEskvTBQzodlCvw35U/Gvp+XiWPLwE3/tTZJLMD74F4YM1hMOjP52g
qRULCeMmTYcd3G0jQyb5oBzwWBxo/1wn2usLQjm19eVsf7OTz6EiLx3JRGeKpuDy
pGOBH2y5qPY9eGfGFhSnw2X8Z3czuulSEtdYEtn81DzqyXDYohmPfv0QFz6qxZGL
iORJ0IPQrk1VG+3lE0+VDw6qS95UUj3rerEEZcD8KCWZIILvekV4YJiaNdOvH1i1
8gkLZRY2kXpMTf4KNXH2WF+e0WwXK0duTMcsZal4Bma2VG4tT83yWcH1VFfp67RT
TsXKyXPaC16OPDnyQ8y+2a40RQlYrVsHwnjZ2hxu5EcWXuXsNG/sc8iyjOl07Ve6
7wvrISNv7fabxX2RPQXabUS76TsIxbi2kyGULBAMQvCbbgY5xbBjq/LLBpl3y+KH
23kfAmgBLSlfW5xgxN9APlncAZWPjkQwNTc4Jh5sc+nogRM48AgAuQsPhkrWfGFc
DrcnT50RwQU3QcHWvN8erbHL49ok8b7HkFJIiuDtkchy9xuvWIsXw3mRor7s7XSz
+H63e1kYnyupXqviey8EG7rWn4q5W+f1AufqH+PcvWZcPI/y0fPJkVcEOPV0dQKn
z6jb2zeAE3/tC5luc6ZJLPhqrKwyYWzcSVHCED/5/hXfnvrxoZ+pahYySA+3RN0B
NhDhZ3nTBPNBGF9WadKBb5vIuxr1hApsQAWk7bkwpoPYjLViLr45aTY2eVHtABBe
V2mFCeNl8D+JRqou/g/RwQa3ISEc7pV3ot88bb9pddsEpZ7eNy4e30l3uCD7K9z+
l1/yltNlwKx34nHkV2Uo8iR7VdONgftnmjYtkWNiccj/Xrh4DfLHlUckd/9U86A5
MwkSY9nt4EJBZYx0UgiJfvFGmotVLbJmnRY7qaSN66uF8dgAullBW1hY6WXmbrX6
Ag6/w8wQqzkCjOTHYNrvx3MjVVeWOM+lvMhyAsNp3hTCEvxXAp5hZuwj63SIdhVd
r+Wxqv4LISjyAA7/BG71j6VMekXEbtdib0nC2KfTIxoXY/vL6RIFEg04lx7D5Wdo
oc0q+cKFCHP8+nercVT4sTDLHqxa14+Jv4S4yb3QvBdGN9VjpTXPj2C9FOArhA+2
KQJTY3z6deB+2fZ/d6Wq0H9dWLbMUoi+K8rbqLZI4nxRcttX6uEQnUBqAudXrTHK
t32yDvDCFmIwEwi/MhqI0WWcVPesP7STjIQ/b306HZ02YbUqXQsjC6ql11gfd3SD
cXSQ3IHMIb2HUTol03I+3ulP1yy3h6S9hROfZv6FMQYNsOaRAst9wzmab6wsb0RE
5xekIJzi914xwIX3NbYrK2QwUig4NpuHR4o+AJBSyMqPmTzxZQvIK94iAItEN4ge
zIjqqDwDL4o+lNIoIXEZjfSTl1PK9fB7rAcupMAv84PKVHkZ/Or6ChT76mZ2m8Sf
EWpZIZvkfeujqM+zQp94AK1mMD4fo3UE+uYStaMUK7w=
`protect END_PROTECTED
