`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PUTogd1xiYFv2QwT4DWW2y3iJN++A2+0y3S5n5bDKvo5rW1MMjy1VP+C8RdANYLu
vkSTyHntRQpftNU9qwegxgoqrtr4zN+Ho2F5MmJB9S0b2NX4e6g7m+6yFfXlp1H8
uMqVqOsbwre3qbID1wZKC4mcaO8uG/brxEQsQIMxSDqNv4DHM9iczE4xRVyvB7Zi
kcDYyBq2lQWEzdGgQhV9D8oAydKWfgAEYMSVMX3eN0htGbcFNgkRkedAZ+Uy9HgY
Xz2WisMwv8IhjYgar+dHmzc8tMOQlZp+WcS59RYrJvyupr7YVry4Yzk0zMni0Ruo
+TT3/I+qqS6nov7diQs15WyxfD0UEmpsCYz4erBz9Cpr6hHA79/ZkdadWYTe6pTq
1RPZ1ZTLhzV2zhzEHGKz1A==
`protect END_PROTECTED
