`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HyTWF5OG9QFfMmY+CBj4/RW9h01OS/uFUsll2oRBWDyeQdaVNiZEKHMk6NmeEAGa
kkxRPI3qMXKiE6GjMXRY7YlkfarIDR6x1f7gp55lOLEeE5ocIkc6x8MJFa4m49u4
ppMHRUysW9J6rJtYaxhD+i/knPChGxLDLdCdqFGuPmrR6Y6h4ZL0BZ/aGmV6HQjJ
zrHE8tqLWp9Nqn23qyP/LdWc/f/La1wbcR1EkR/PaM+Ag9Ojq9qqGLuNMuQI78YP
iITHnOtMqDXV8q3koNkrog==
`protect END_PROTECTED
