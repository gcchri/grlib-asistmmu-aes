`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ot1ONd5xLO7VRBQ/ETUy+a9D4QGtTjVjTB3AORB4APBrJZhlNARSHTiHvbjfNFi1
7tq04GvClMrHFqPYGBVFygeuttjj7jPvY29Zd+lkcV4ViVasuFmXaSo3hhXC40wf
t3EkrHK2XxjYP/mnQOvVP30h1LLnmFksA1R6MybiNGyQFodjEc0LtO2l+EB7nIn+
FftZFUuA3uZZDAr1iQ033F7jXBdzBM7nCig0fgXqN0b1NeMSwFJY4bLcS3RtoDKI
L+mSV6uls4i0AsLB1sQDxT0fbgh3+yAhc1mz12OmbQy9Q8Ncs78gTcMGnz4szSOj
/A6amy4tXCazLzMihTWbXF0lw241OJ1qcETSW+a8IWeTWv2v/dHte71Llcm2Yuz9
CP63leETBPnqdTHSpxBsPms9cwTDQkO4hsEYl0DVNvP5GUGuXP7U8U3WddoBRYz4
Fa4Zx6kV7t/TL/x68D2yXzFfQzbVAUBgjkKgUpCRd4EYhg3Yr6Zm/uChAFfZ/Ijj
35rgb462L6EsXG8PLzF2UsXGz3myRcaOex7qm0Nl1uE=
`protect END_PROTECTED
