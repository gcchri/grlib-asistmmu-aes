`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jnY8JY1KuVuZsA6+NYuLGx5mr7ufsgTzDzMRh3WES1M5HZ+wuVGjBhSvY17s7igh
8YkqqH9Qe3qjDi0q+Cj6Yr44PPLs7V7u+wvtjytn9DDE4dwfOMs1IohRT4EOGp3X
WOJ9ePLDAjih05yxMRoO6QLb9v46c3uosUkUKN/YV2BiPVxywRvcoWizYMTq478T
60//72KcDJe84I3E0tHxxQZoe3Ls4KLFGQ+I0106cFK+meTolDcDqXQBzOt7qc2X
ugEkYBBCCSgRHqcNKFbKNS3pNfv+UPO70TEdTE/Rn9FFUgKPTTl6MrlM7XDCh/8D
qBs4JSpSlGHyE3cDshJwPQkP0jitzEKEB1M4ySAx4MZhZyRlBXCLc6CZDPAE4/0g
UJbBJvVMGOSOr8ofBQh6d+7yHXdka+Rmb5xO/WcjKGQ=
`protect END_PROTECTED
