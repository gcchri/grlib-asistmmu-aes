`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IEfh4E+RhIIywI8WMxeDfkIkvFQ90TugEI4SoMrujJWBlvY3rdsFwTy4bwE0HJs5
qyhpBPoeomnw8eAntKw3oKQA8qumkQEl/eTqG7F2ukObGWWRLRzGMufiKXd5AL22
JevefvT267XEzmqnqicqzLQhlbMjKJ/kWYqC4jE13wYjniOYRMbv1vmSjRiw9A9W
HvpMRwN/zRH0y/3dx8ZX/j8n0yCDiZKeZMWIgIobfSyfa6nB0AkMXtPzHaWVV+it
JTE6ALQSxh+SkfOFuQ/AyWZBobXe89rRvPIrA6RVDIoCI6mIDHC7wY9J41TXx1vh
HQRJR6liKfYLRH/7NYVN6fq3x0gwW6zgEJOabUkCxnc8O+yC4mn47Sl7NKHlA7TS
qPJfb4RFUXltY5kdoar4Xvmc/7XK/8gLzrLA+x4lYZXOcBcFUdA4vL5ZJemadni7
PbKr1GBo9bkyfoOwuxLy0EslbJEYBNu8MiLOnOqz1XCcVuXTmACYOsx6qNPhqlqA
KpifNJ5Ut5U/m/P58EVe4nHzJJRPem1VcGaA7uW90bGRlurHiyhF6cN8rA8jfIfX
qeFyB0ipJq4bfF+PlyuNTw==
`protect END_PROTECTED
