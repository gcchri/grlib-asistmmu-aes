`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9N6QANaRF7jVzuAfDF8gUi/kH2t1+JlYBrTGOXJnZGULT9q3uoOVjyU8XIAUoifO
iQAHLsNMw2La0Ga2PJxE1YW2vk4x1r5ojjESHb+2yI1xjTX3d0Uh03gDSQxYMRuR
3qsii88COcYOIB8nguyI0pdBQsPgYB7+5UlQCdg0fqXBkzwcaz7qivQJJVbe/XSP
sQOsJnxFPaDj86SafP4j7+IQelgMzdfoH/M+J1tyEfS3t6gA6AQRjcArcVR1bTYm
52q99uQT8vVv2bIZsicbrYCrDCj64jfnvBLpEIzlMAKB7IO/VWfm3a0vUgBlBYa/
EehoPV5/aEc6e+xf1er3ZCXoK652isUK9CfDZfUgDvC8CH0lZqeWfyG8amKR1TAF
RigNd3T0yTDRlqdj2px6BzSpyOaUkK9mjVki0LHOfMdY99/Y0dsnqvqv+pPliS1k
fo/hwmH4QY9QP7nu1RNROa0bx46Veyyj8AX/ixXH1Xx8yYdQ/f6oDOcXoD3MUogu
kP/9OQqhL5kstu13RH/0uXpUTL2GsSS/yjO2vVvyYv+z2+XF6+e8gv1beU1ld8gl
wKdf5do+qvSk2jqCBOq0NNu4UwZKNtpUdN9rEa2v+Cd2rAo1QT1FHl0VlsKUgol8
qN+CbwROYnArgu7O19lOJCJkp8x7aOw2XP8yy84guPY=
`protect END_PROTECTED
