`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uZTxZbfzI0LpXXh0Z4nzmGq7S/sKw3Or+7O0ALlnKTJgnrVciAppwkDikUvZVrym
I1+IcyS1EfULD6zuuSPBsoXCnDJ8SsjDmwnayYDI60Lmw11uonbzIpMYF+tnwzfa
XrgmIiaVait2v5ylA8xTsfZLo+DqDxgaHczt6zQhy5vjQnsTo+gZGMgXNrsglZ3n
9G0uG3ejKPJ+77C3pwm8yO5c5wY57Nbb6AGLRXkOZ2V9Eo1aavhA4Xss14IuNaEw
4a+oJ5I+eJI0QWywegNok5029eHxjouWxSHUY2xN/Yqmap4LjfWb72rfySsNsR44
zEScLLvLbvwsncqlvCVcIq0NdgKlJE7BhgjcV++UHFtOag/tcK6vbWBarcCHujMC
+fxSOGaK25xoHrl1PfWdNsmXfh8lNEjFPDBPbg1UOzN5vPgmrBbXpUf9mhT0KAxf
e5gABC+08wo1OSf8zufaQpWXR2veVZHIj8Ctn0bAVm6dd26hKtlwvqIS8B9SzYVk
XIrLZHxeodknJoyscAEYa93faFIxO++5kvcCURjivygYkXmF+JaJPlb4M5DH+PxN
bszHu5vyP8vpkVVv7OrDx8ag7Ut5bD/A3ci0qcZwELM=
`protect END_PROTECTED
