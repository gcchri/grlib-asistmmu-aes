`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fYvsSdocYwF2KVpbK6ju9mKFoRBw939ZYbA5i4OIv7SFQyfNbSeUriXUWDU1wmPq
q4JrnaTd1BF4i26bnJ4eHrq8/OI10aMn1OeGH+lHDS/kYrIb3EkFDRqPUvhhOuwt
NeZdh/pXkbeI6FAMxUYlksjIZGV2nz/9advOyjKQaW0bdJkztMqiJD0bFT/5+KF3
riHoUnbljjkBGb/1v/BXOJFIKW/iveIguXlv/OIW9RrkorxxOnoQFBCOh+nuz4yL
ZBHrNvAA8vpa/rlg1gTYzoXmInZ00zfrKFWsimHrPfgQ0WAX1PIGZpzZSzbWgXoC
vLpDBH+4AJO0Lbvh7lliP9Q9nWOcAOVSULZcYyfB7C0RV1W9fsKN24Lv9w5ASRfK
AUBsM+1vTYmSdFP8heDHrKgcoON7oxdYPRpvPdPX87CqNYcrrAg1IPGn39G8b2S6
RbyvC17JMfQ926NDLe9XInlo7godFMTYFNy0YKxlx1KGF+xfAE/+5nKniXi7Pk4R
1fj7WUKf/ZXCf87inD2BSuqhy1cLWAAvzqMEhIw4e/sR9fnXabXl+QSXbRmF+93H
yJEGf16A/0XFs9MbatMr7OmmVlgclfIwC6aSS8wB78gBaBHjU83CiUkiIXTzBWbb
bM9t73u1ol1ATmGS9Jvq4XL+Dio+uiebZFzvUMkThCMz2ghftSvZC0d+BKsv42JU
z1CKc2uKMKqOTpxLHjlPnd08StIqHp1isx4YQRdjkwoEGrDUxDcY0WCA5DeBl6+m
F+PnBQygst5lFe5aEb+V0cHRsQ/EMEeq+e1TesZ7n73oYuyIltYZYtz8rPL5GMIl
SE9Fbi0ljly0lneK7l9Noz8WeEfyzmE6FWMbnBEdcW7fSUyKA8FnY+Bn1OXA3u9Q
hcaey7WQ2QSpZhjcLbKfnfC6FNCVhmW0t/oxdMjKG8SVv1B/MykA15JyXevSebqO
xzQ2EFlQt/nlQdj3HJrBCv9SybGxE+Uk1svM5j17hT5v66PsmG1IFzSsNHL1yF/v
4+efPtA17OfJX73NBcsdfqsP5lDteCy9NpWJ8uZ8SZbV2f38sAKsEIG9kABzaBiF
AbJTUDptC/x/9JUeOw0h3nvfo6PojfHMbv4Svge6I5tt7vdfAERbLaEM/W7KFah7
LhtLK3kR8sqKhrPU6Fcw9vk7WfRRbGutBDoOUpBPKl6fj2MXGQ2gLTZNB54EaEpx
Gr/7ERPmksmeAA/+dV7nM6Rc3yXjcg5P51aiuBFQ/qw6PoRP/P7/bO5i5viwxcuW
IdF4a7aEUGF2+6B9wBvfDZKlLr5tvVqEl5uHehxSjKWDXF7YMB2yFVWZ8DENQ51E
EzgyHj5bewSflGh/l2+xe7NOphKjNuO1DO3UpDt0BG1WQdLlVmrAfyXE79TDwPRZ
wU4a/S9GpAOABEQNDtPGZv0Hm7NIdFFofOd4T4ScleVaKiby+RB8cwF7mtGPaWxW
L5kaDZkzU2eOql8DNdaMtvdhYBajsDwR9b5dwxsfTMUqKmIgUUjfWScZXYa649ma
l8oWgGZQzfHhKd5DTcBbaH+DIm7lWCIDDY+o0KwLTzmyS6KL7HHaXU2koLt30C4S
7ErJv33BTtP44Xv+8spW786JQsK/xglwOWjijbrK8Is2QHYNkXXSGfIlLyTXx9to
odaqfxLxI5bhETFHMsGO/4bEcuJNu3TrjymxDy4ylnIAKrMN4O/9/5YkYA57Bjz5
AaLXw5VQe0k8ngYhh8476tz9KlnzjGsRQVvfXMvDSoLDUlmNgyQOkrUdENdYhg6p
UgFK9q+uIXhCG1gYgqi031CHvRQiA2e99uOqtInUZ6Koi03U7s+A/gecWvQV/Z/L
7v8/f+MyXYplt6r/SVxIfheriX6ciH6j5nQFM2gOUd6U+vak1K7doe8CIm6RKRM4
`protect END_PROTECTED
