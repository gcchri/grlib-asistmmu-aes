`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oZ+k3TW6lYave3jLFFFnf/yX1K+UQaruN3Wj2UwNfvjC+rGJNSHhEYdsCkoYZ9PT
b7mSiKCxQyz3h2WsbekwzYtGZWPjHesQzJTM6O5e4syIIdNjN6XtzcT7GL03J7Au
cCCBq61V8KBCAGfhn8OA9Nt7LnSJgJWcAZ5qQDaQfJoqzXVPCk7s0LXauW92DSVh
HDsOXinzaOxqSSMB7fD4Sh+pF7KjJrf/Etm/qEGycObKSiM8BSQTccKTIu9Q4AYH
Uef9jxhgV/aC1BfjQr1jEG8rw9uO1g8geEaR1ehw126vizxxZcKmPdjRptG2C+eQ
9mIFfB9wiw7K5xbErZXNZW/5efqp1tKOb4vLcwzXuya1eiUoSCrkmFGEWf2FwKa5
+wz37infjX/kv7DfD93XS6AoGTIWJe7EbfTgLvquAcCNJmnxRXu2FjEWRfqHwqJc
UlR4rans/caHPaIvXw6x995GCqVzYbZxL1vpMpLr5UM7PCchBmYDGSycQ64rkMrz
c67s9CpkvIuCfT86/jCN5i0yU6esdEsjqL9eSPLQm8TnVOPIbUKmqOQioO9imMuy
Oq+MdSWrwhKb2mBSchEWQgxxCXc3PRCT31ktf8R10e9ScYp8ocWFa5gKllWAyeGX
jn/T4vVo/Lbx7xxMJK03Q6cGMvIiy8cqKWClkEH2miJreKyGukfEBdtvWiiYUctG
QEPXKF+vVp+goZGYyVSTKne90QsqsZGa6ZjzewPyZCNpXaXDEo9ERCqOMVSTwSfp
+attTS39ITv6CE0wpTSRvOFudEHUgTyeY6A7P4MPuroeGl1IsjvbptFmFMUCLpd7
AP6RPwI5s6dPo3Wdvqn9ulJarpHinBk2o3Jbqddy5XgRLo10fie6duLgL21uQTXK
QS+Sr8yZNrJJ6wdlTfw+ZXJHpWaA9YuVBUIUpCLuwao7fVFPp7KHBUjelHaRKTep
azsXmK8bJdBWYxYA0lDyTdj9uuKJM/0sgcxEbsvCYRo0TIt9otkqiyJ2cHG3Ln3i
TEUtdWptAwoxiAd7aZDgOwGg2Kp7k7gSlOOp1wseO6tuVkgM4itvc7PNwSKTUyRE
cArA1txS8f+qCuQfU7x4e9zqa18ibPJ/fxqSD/Df9lA6xP4bcownQhqqHZbxh0Vf
ZFgU/x+dH7zf8yg2xEspDC65OpU15/fIMO61flPdhmeLGvVlPBr1MjZh3Kg8vSrC
XF3NLtfHVTOtitg599RT70wxJIxl0RSvr3EyHLxoIcuj3tADcu4ZE60NSlJx5O67
BE+AOX6l7Ibl5t4nQGc3zr0CdIGd4O4HPETfKJwjHGPHNJee7fFbaVPNkf9+aNRm
wZAEpmADpYoxhEd5gmb/PnOY+8LhiYvF6oy4mboPnXn5MNJdxV3EPoW9ivY+gpwt
ML6Ejk5U6t4xtOu+3tlcZpMEF94LUrGzUTG2JNHOLhelIeTXVrNxPGszwr9PjLk5
XI2BMTDHa4F8cefvnfJOvoYnSSmJrImPk32FMm0MyGncs7eTAEaKGB5pWjDKI/xe
slcT8zxB+Pbc6QE9/yZC9uen+2uFfY7bbVprirSofTZRBf6wywSkvYSJ1q/vxzDa
3xenKOyK/6SSdnveYmnLnDZhshCyof5oULfHyNJEYid+ESMKufPrv8+PmUP1dNYC
QkjpYLLf8LpDbh6xVt22/jm7LUwc/hdTZyKIKPqYvnM+9YmKPL4l+ToPCqw6VmDb
rveqwF3sScPNNXu5h8jnWzKnFJijliasettp+Tq2v1hpvQhWwz/aBPhg9773HaFp
+XlzZMVyzzDWILBSl+Hnco2B1O7S56rtoog8ghWSt7oBvCXV7obWGvN1JmJfmF7h
A04eGEruFKRyFScIZzzHQal/JIXrK5m3OhThm15S7WaRbN+RrNTICgewjlDhrY7I
chfLjL8B2dXwDjHa922DNMQ79pQWWWnNp/3ZISQ+um7zSgNYnXC0bLUxp3yEIxSp
GSOzAdYIrFB2kJzM2HlbVdOK3uF/zqjMUJDUdaz6eeReTPtVWLwgIiL68g0UTgxD
e0JeODmxhtjMd009OrZ3TJeRc9GDq1nUPhH8hmYI7BpjQi3K0TE58U0hWMlSEVy5
xir2Sib9TD4KDGWh/z87JJdXYXs01g7PlJKR0+fyszYrGgdYWW+WwV761BShLFLB
zTiQ08JCRnuJU6TBfJNVKyXVYhA4IpYiOkM66jVcIUJo8aZ+vl3UJRGaSPgeExx0
akIlozRnd7OoWpRV3bMKUGt+952zINEZKa6YEUsOfSZPOSUxqJJZnTSCybqQpgfG
jeXbSGXOGCzNLU9JgfXUzIfpDf7NuCFGikCps86mKmpglr2FWKiCEhyBa655a2zJ
IbBnIaIhed9ZwI78TfT+quFs+ugPUn/jgxPvJj7cnejKxcFQJl5XB+4o/SG9Q78K
NQbDObZPYy7f/I5xac/yeHDhR9XY/s3twrtq4YQnX0GidrVpC6dN1EbvUzZvT5p7
94uJrzs7Sx2SdUYPZbeQos87ijLDzak7TXFgDuuACPsKIXkg/UXjf7hNvHzbUxZo
NUmgrk5Y6zLQp2TrjSSAPP7vpY+rZz7iMFOX1FCWKB7K/s0ueUclcF8epGShY2jY
QToAUMP/8A0LorX5Pc9h5IzWETT+z/d5wZHzgiPuBKILAzN+Uf/owmCYpERbFFya
KGmJY+lGpHGMBEGA2VyFLPIyGrAS7FetSCUzyhfSmbsuiq+qDOVmplqwKoTYBKVy
QZ9CyW+XQNOouXsO95gquAzOInMx8Kq+k6yOCXdX9szhMKfnx9k7dweNBy3SxKHX
IN1SB6xFJnxslMyWZ1i+U/uBOdXtlbLz65j6TlxAvFZ0MYuNHHXdZIRi4JEZNiwP
Iv2GG1PFOHn4zBrDBFeBk3siWwlgy9W8ycFFWb/2beo6V6q1T7+z7yqALIOsOKtN
hqA8+vtDMvkPOHEfY+RUYCwmaX9O3m+POdW3WgiBJwL38wQzUghswwQA9+f+TTEA
MkhoKBwpDVAd5RE6sjKeOkMCX9L8QIpspAP9KDgAvoYjcW+1C8AzZovgshWf1doP
OIjLMTY0vOswt/pC77lTx+5LGbqT2aV+2I6WfSGRewEbdC5hdLdUCerU/6TuFJpx
uLiht7OibrWmRTQBdqva0k0pLZzkaiiFWHnm+NjA0ylvxHhpl/Tt/oBXoYrkJ5GC
q/NztpFlwxGhiHP9OQ5+mLj1GkL2ilvttrmMgrTbER7AgGa5bCVyq1vfybd7Qdoi
Q7Vf5ODY6B+NPwnP08LcnzIxZ6ECdVhrZ7/V7bAyO1pgFmpbnCLuzEEir6Jx62vN
qoenoboAs0pgvcjmSAHDhMcs3FklVrGgePs1ApU+dTnPco35JGm0ODo7cAMVfLCA
NECDcptR2OmHAypE/2dwk9ySTMswoVNkCyMH67AsE4xyLYflRW49vFcwFXPvJXkw
t5iwC+iUVrbgiVNWk3kjSwsdQMVuwjpxERvL6k6PP3z/mLLAu1Fb0/8Fg405HMye
Bna3rHjeq+fqUI1yGArEQgsxHTXAqs7XTgnPkPHyBFogid3H8ZO7TasCQ5h6jCKh
I6hwGldGf0aQqiDLm71FyVKg1YiwCbUQIqN1SsF5dsQ0TjEuGedlWxlWks6tDseF
Hj6mnD75DVdF964BNnou51U6fEUzy87fzEbNcvOhtqQFE+Bgrd/HoUu/tTQknlRK
GzzjLliAsas2ADcY7X57h7+pXnUhm6nlmRg9y6BKJWYrIrTjMTY5DaDu2NPY6wLf
79vwuppqGcGCjL0piCitI5dO007hNzrD+q+s03+7kZAkrGOE9CeTl1c7T6ZJZuI5
mixB+b9udqn4rK20NPW0ta8oCnH5F8QXtlgjorRXt026bZfGLFqU1IeBgyQNm4Hz
VKFOz2QvZJn/ACIRfJq9nwSq6wmg9l3pTZbWik+7ZSXM9Q4qOJ6pti3AhFTPdAha
fA2NEq9bODjCMLcLWaBvgEYmbJrgaTCNkkDMxR5WurZhJ5o6BI0yvMsk7BT4YpaN
Fk4HI1IkMD+COFRQMx7Ue3K/bG4CvY7RTIllFUeai7CCvsa6AGapQ/ZSGvtiYzcK
3fOGU3pvq74r42wVI6IMIeGI6uW9zrsBU1aXUi1JRNCrfTEWjqRuiLJqRyUtHYWC
ZmorJ3i7jZJgQDnCjkPSrivdd1siyxK1f/9EkfertZ8mFjXR3bafKodTPU3rjQ0h
FksPs7yKbs2tpcZnmCDFQATuQWTfiueBTli5i8El9EzJqB1JtySHIBF0zd4y5KY8
yh4kYGPLNW1sVF+iB1F4xosT523xsj5Qu8A0pNKJ4VfrTH2vUbwpBUEg0p7I8F9n
UEldqBnrz+WefQD1l1E9KvSvL9sZ0DWJFw2vNGkAHgLfl83y7aFxNpCaG+GkKBP1
ZWAemwFiejm4gdEexcLqTYuyOqmvJGLCF0XlyV4AT22iOq/RI7lZdDxx+MJGGue2
KvLJC68Z1eZH7yVP/rfA9DW3uiC0TExHJRUAVhMjZxykUh0dByhnhRvo0//DXyUb
JW+wIc9RHVi/5RDzovLJKx+J5xwEezm775Iv2iYDb3uoBJiaf9/rQFNOexPnUZdY
8mEmmRY5bZ81qQkhphSwjj4NBnodqrKMTCZp6f7fRuPBG7f7nXL4zNM1vPMryScJ
QjpFk+BfBQUrTgqLobBxkxBEBWdOndsaQ7AtvmsUcsZQFM9kA3HxX/QxkcbptDdQ
01kez6zsB745trd5wWsVFIPQ9BzpYBif9guFh1FdQtDzce4ykD2TOqoTfQBgUozO
NzqYJLbCWsL0mz8mDJjfIAlurfo5zc/kMW7n5Mwfh9WfUkwIWazuQyqoPiZS/3kJ
FPQZMO+U3Reb96q/LJ/dVuBUE10ThA3HoIpbgV1/IiNK5vQwzEjxpC6+hLaQLznv
QXJyuBYdKtnTdVwUW3gyNsFQ9UexyIvyB8x4Rg7DFzmwd1tzkxiWJq4Lqq5wkMC9
WpesuPnJRxS/6SZrFTYrVan23oq6i7XN6yhRLhcdORF+iXtUKv/eMxcw9m6FZsuU
NNOVQ/x5YcI6tmF+YfjihZiwm0WLpQYFOeqhGOR7lOps5feRnrNCzBHSx7D5LQN3
7rxcIhWf3/wS0wh2HcwPfXqIDmz5rQ9UBoNNkUQJyxX4/t0tlggU8F3ZPrcCYUDz
voeMHdH0iCuS/G3Yrf+ExwOKiROo7Dx1A8tlNVid6hM6XiZ8zB0liZDdIQHqIcJa
WH1TwZWZXb+E3NHtOEIVPSAiatm5PPQVSG37ZAhDNe1rSQwLi9iyYZCObJptRS32
dQ0bCyjmC+OPs+oXgzVWePsueXxrjSVYJlmIVMhzYV2M8jBHEwaqDQ1e92LTCe98
MCEVVt7SSqWDudHVEzJEv+EEv+uMX7wy0tnvqbf3iqPJGRp8wyn9aicGFCe1E8c2
KgMEYNJXj60D79m47hpHTsmlnwERL7RcP6MUcfdqsvWrtTz4TWgLnztzjn6ULis7
zKZAqXQC5/9Yp8rhgX1h479Ae47WOipfNr/GmzQgfZj2tDF5xMCliYpY9H6ijD07
hDfamBluAARlsKwG3BardVYej1JKO1o1iQ2WtOYwKdh5wek8vuQ35PgRh7rd28ln
plvLsET45UDxnnvfLJeNZc1Sg7kjsnMmxeeJkc/n3lwtpeoeyHTRxKnk+i3KZAJY
q/8SobG3ReqFm3nsipW5XMvMWn74Llie5ULbP1VRsUAYYC4QHEla51bfkFY3XC1R
j8FTrhc37kB5/CUgCfhA5KfOC0s9qUwESlEAW18oSXQO2e0DAp03Wcsa9IhIxrhX
B8StMO1AqByPz0hrKwtsUlwDwmuQvVhLQ5d14xr7O5X2wSpbSEMZBpZ5awr2wkYb
UgzTXxP2D9HQrS6as8Lbt3rQxyOHNxJh+L8HoRqxJNbVzQykXlJw1PUi6A43BObI
3Lbojh85AKKVA3TfSGvx4qWDIaQKaS68JR05ng9FlwA65+LP7mIsLLn9hQAStbY5
oxnQzXj81q/3vnVZ+FjMji/ZwD7qaPFbi/GpD3jzP0pOQYdad0esdCdBwngrbvM4
+feEGhP2EoLmepAHFWHP/+T5qnP67rrVawa62gI1DoXsozySstRWS1PSX1fyhki1
Md1uRmi+slSKfxl5N9JJoFsPr1slo9BsSQQeGTBimwqXU/GBMSN60fH3kuakwdfV
J1kjxYGu9ZI0hCs8V4bF4GgZw65EJGKM3qnGT/5h48BzvuES8f2MNOgU72lj9X16
NMW9GcpAVmqt09K7XS2P63rTOo0DA9Mk0IAfxdZeRT+M6MR27qEgc0jCEk2nNAM4
x4DsKSYGnau3lshNVNdCjHRWw73BvMxE6WN9Dl0IvgywG2L049jaNk4yh0yreUxV
8V/pvDVSj1WvOPLPYEoaUiUP8HMYOOgp9kkIAUVbU5+ZE5L4V1fGeyRBsf5X/FIP
StcWH8GI/89cZMNLAOXL7a4MFW7kQ84hyfpEE3jFr83iO8k1ua751nTfKvI7kHH+
W+JdD2c7XtOkAGiT4yUjL7HUyRvKzjIRSBVrmOI7tsUzyDos00qeeUFiExcEc4Fi
iKXa7d4cipHnctCRBexduHCGLCWPDKvCwBqjgVrOS/kccsMypoXlkys/D23ngvMo
G1h6aLfMomDXuJcuuBpm4Cf4L5CTDdV2ReTdsbqNHplW8mI0LLFm/aYeFBcj4dOn
uGVDwETWorqQdpbWjm0j9Cw7EVDCeNO7hLfq6EpEnIA4u4chXxMJEbRc4ldMOoz0
Nbv8UjIPrYFq8u0lumcpbyGmazyJ0dgiEBzLMVnkD4ESw/SmHU2M/29ghP2T0n08
aYjEW/lLgg4RvvY/oYGGTfRi/xaGcU7OVjEygmW5nfaY3S3uZU4UTE5gDxUFulxr
4xpHTmMv0eoajgrqsL2iSURMRXK7AHTsaleuhIuzkZROKdEshOLXREn75zRg975i
iMKbidjCppWJGeR0WYhlTrlVxLrY/B0Pesh21i15dDG/deXe17cr5T4OIU+5oIiV
udTDobhXwr2RIwNtNS2jZSqKa+ytr66pnv93Efye/EaCq+bHM0oxlWorWy/PtSZe
d734fu1iEQrnbMHKNmcmoDJAaLRAAG8ujpaGpEbMJ/pDgh0zfhdPnw5+6+QFDT6L
G82kya6cKEPdr/FbEB+ZBxJWG4WDG9ydC6cOx0vRAE/sGJSCY7q/gfzXCmxApp4P
9RuEM/V3sWlqH/vRwmN755/AoJVB6Fp8R3pzZ9X48AWDVnf+EmM584cXQYKo1E/S
c0hq1mHu6Tc7lTgUzAdvBZcmdACIb7qCoBND/QuXUKTh8y3A6sIoPiIidRAct9+/
yoXJaKd3P8xnvdJ1b5B7YPnjN12UrzxCjpLcxR6Jh1k/qxFPx/RR+o2rKibaQcPS
dGHKmNqc0kkaQEQf0XYaf10VbOwu6/5Ica1vGa1sq8ck8AVskx362KERH+D6+MgF
isX3DQdEbeMMrJPCP3/R5XYkV/yagdcflVtN4WyyQ1VArgx+aGeGNFX+KaZds2h5
9R+p74QHCCEl4ZpC4iiH+BfCpwqiIUfaIthiSLkaz5Bd5KZNQWnL8ugSgeFJI0/3
kuWqX0A57vt0Y37dvWqMoRJDYs/8Le9BKmZSEGiIl9nsmzoMoqYw+Tk5/f13j354
/0SVKrJLDFD10cukTvFRxArbNfDf3kDwyAAFz2NXkp/ArTHa3PBneyry6dDyYzRL
vMJxKc4IB+Xlb07CktGWIqM5B+Y0G48/j7BvcW95wdQFoInwQgOXqp8/Eupqj0A2
Y9Kj0EIYQb8hRP3TTsoic7YeR28KzBNSRP3yPgwv2HQb5Xgxyy1jYyQb/ZZOSLYa
EVOEoJhNEFohjmDiHTVuNcHi/jYiyeiqgSgh/aRjrb2nWFrTy1+YS8QAtjCkVxnd
YGNjL7RBGER30wtCRN6drcR19uvqFAJJ3d77TkXk98GPd673aoo5dVslvJ8wv3Ld
LV9Jq8ssBlh5urkJNiTAafy1QqxZMhGAwDYxvavdutkEPHvm5AChzwGKyqQWROXJ
tafZFCmwLP6t8TXqdhvQ1zGGT/kGOlLJgNtv5ssciNoiBfUEB1qzVLvUezKNiGEZ
4pIZde3V1nR/quAnibs3HrUDaHuPgpeJhWD1lD2ekVm0rssb6s5RQwhXnyIJiAWu
spSfAxtt/eIrhT87d30BoqQe6u+8+69+80lTKTRQjfQk6lpjxBAZTy99jVxz4wxI
WRzTXLtkDJwmR6l130tvVYyNs0j8k4BcxXL67Std1ygFiTih6nwamxjwA+5xaT8u
iwr5ksiPBb46Iqa7ORqm+KJxxvgblKo2RAfRInkL3e4uuNnmpLERphZUgyukJqqe
JFsJw4fq1XNuRM3RqeR8do8au2yf6GVFUZge+ZUbtJ5sB/zwL7SrsNwpFXhz3SPr
k9IprCtDTDQpiJ/Gh+niX3U1YGCNnOrJpqRDvdHgtoVfRDNZvz0LADINMPSCXd+N
pT3kRQx7afvbN0FB1qWzpKnpAL/WTXjWot/ejNnKRYUgUCyc2tlSeVADQD8aPq+s
2NdYTPc3mmJ09+X8wl1u3pGV3zAPxyPpN3UMMmJbvxgWPcM6aO1wAezuyIMPpwN3
68iy1CD+K1vxJyDvDayf0BsdZUIy2+5wU1Zxz+a5IpLO5ctTBxHAGGXGGCWppwbt
MIU0q8mtYjb8QmGztvpnR2qwPKNpVsm1zH39odj8Ue4rmpQv7ZPXVaV9P3YGUE40
6y0Js7LLH8JchXFjAZIilvykqVGzVkaqCwLxZgxcXVUIHOLO4+xB3889rJSA8PuJ
Op46YTgl5xeYAak7fHEH0x/SCUxDR/z2UPrRzihnwJYcVj4NwKiUqR4ZnbhEZkUO
1nGnbEwqrKeDsWdb9rXo3j/SnadDAGAlUWtMD+38x6d3bm4WP/XOGjEyegXeZTKo
wnpPpeEcpYZkjtVZUhSRMAetRJ8bBr/QH3QkzWer3RrI/0m/K+TArvPXufEbn3qc
fkTSlgVLNSr5P9cBhS45FM7lJs4C+38aKX14d2Nkn1YtfJ835R1dVPIoJpQFDLJf
Rh8/oj6sXLy4lI/thTmn4Y/h6ZhtMGe4lxKPxOC51iU0wrH4uywwFQk8krHK3CJ7
WHgZpu3K/DNvd1vkcRS4dlf96oPowabRjobElwpwTnaEDC9zIkar3uCxRkGE7BX0
eljI7jrfFTov6k6RKG1S+il9XsS/+MTcjuQIJA2LjFk9mhGBd0YFJcSwYP8rcR4a
rDij1mFu5CBbB1obstE6/111chiXRhhHI7UQyCE5IzR1jiVXhbIRDJzM3N0bkQ4h
AHNBL3qMJlFWNmDYcwwEpR26zFDKdxchTRNFIpM9g54CZu3obZmUKSdtIuV+QepD
gEfxMonVRhYLyH1PFqO+JDN4BzGA9O8JDi5EijeQtB/ZbYGGvYuDC3FlrH0WEeuW
H3kvnUa9TuA4Fxv1XBg5LgqtuXmN+LxruTUYIf0244QGVRS0mgs9Y4695A8ucqfC
/EeXjCgowxKQ8XdQa4JmCvUDZX8++vVb6kGMb/7hWCDNlcZ4l/i82B91BYNV5rgX
0Wo440KK/5tZH5U5+NgRKxAJMRDJvQo1JSzZQHX+nfoyuCwIE16pgUJ+3HdCz8aZ
Rogf8mpewegRGRmHLVLgNn5JKOdjZrPcyXuZziueVJqRs7pXrOoTTQl5pgY3pKaQ
X0DzQr3bNbxa1sgaZvMnTdKuoOcRjS00VeY7MQDD2ADGIfXuUYpzXDmKI9eK+H4k
eF2py+yKgq6ENePK2IXbNXg7DDVxz2+lOEEhxUNccdC7zZV6GgzoFutJjLF25/1b
1HsQ06VXLIIFmwxdeqDskw1CxUskISlVZEk+3zYFaIJM5iUrk+Iuma/tlftTxVKP
pIbjPrS+0vIi6OkiuRFWjgqRmlwlAkriRPn395NLPVuLtsuunpvSnhONoMqarBYY
TKDNBXIBa49pZ0tce4oSwV/rBp3ocq3YINDlLl2SEYVA4baQMsSwuxRS6g17CMP2
k0+SyfoAZQUAVl0TKM6wqEhjEl3qR6CmEkmMyQCR6Br8flx/K5u1oGx/Qrl+JJMJ
3MYn+a3dvfH+/rgt7DRZGhcDkRRALH6X+J79VmaLa+BEDJaoUfGgBM9ETM5qkoUB
BrwiJ6Hi0G31t+kgU/CgkR3c87sXu+eTedEn/JGZWuIc5aMuieXNeYli+VVzJCIi
oRWpeoDtQKQQQWns3hrqFRCK8wlDdLLXt96rlhIktcgqezLS+YLZIm1d52BQ/h6x
TifPgxS8M8ZM0dizg13reNtLG6+MJrVV4NcLTY+xy4DTO1bd3KVyAorhwbm6PHnR
ZsA3lhiHjA0HdoWefY5AC+EMNGmITmv/Uu3ROuUeg4I2+DWASLQopvQVvrwfuOQS
cNXyKjV0iuwJWwwjsvMfHAOr8ammnmLcAAc5jL2cuHnmoqk6HUuH+MLUp4H0I/8j
Z/MA4/wUPulONtc2okNft84CQmd/+3F4pSHtILjdOys/YFwt4Pqm+ZLFGwfDLFmH
E8MeoQbepnJH4UqZAs5K0b/SVG3Lddo8opeH8urreDK9XR0pC5dCP2779XWUV8fS
LlF8pTBV19ZyjtUPxXIZNlGX97v9Bl9zhK/JXyfqXaEn2TblJ2LvVu6YUuaI3Av6
MhYJ8HX5D9gO5D9JUazA53bFnAM0ck2Afwe8ONTWniUjzRsZTEUWqtXPCVPMUxyK
uSRSo5uNkDDcXk3nU5xISZSU46ln7s9P/pH+UgZoff4/YA+/HHUjPcfsh56vLTrP
8D728xE5T4EnsqPafNc1VlN8hf8cycJKOcgsC824WOFIebipm8gfuqBJ4pxCZEdv
9qZlUjTMTuC576v/FD4cAg7Wl7QPnshFPNpFs38Ql0bjUeyu0EzP+qcAiALW8OOw
Xa5LnnAwJBgzoLF3EEb6hBCX3JSxs7O/CGRg/9FmCkcCdradaSfiqk8jm+6GbVhM
5laxQaAsdIP6RQxsc1Cbeu+Idwo4uQXCARLVgTmQ+wUhAi5BoH8qH+jIxO28JNs2
PHHT9lCk1MKzGrtAWrsfZVZumoyWemrWyeVodBKjYkBDZGwHWXLBsO+2lB2VcJOu
qbR1NxueRTHpCrUHt4RF5hQBDSEfQ4vOmLufeUgem2pcv/oQJ6PCfjbDWd/fHe/q
3tqwCqrdkNO1UMb0XrmJ/v3Q9VTf2a+MwfR1BUyk6Kt1lVH8cDUpMFQUQvFbuJoQ
q/7H8sgsL5UPnJ4Srb1irbkrvA/c8MHgFOQ5RAvUco1dm9TRgLCPnscuoYq0nIro
WTXYpIATJVEzx1VEzoy4Q+vd5w5wK0O8GjaBZEYxaYCyNh7K98ibqRER+LkjARH7
+8TrOsab7x8Izfpg+TC5zug75t9stjvP2lRLJszmh23LErot5TjMoip7zrsaAknr
+juGjIVGPYLi4sRRQ17u+Ap6GbidO8TBtg6eJl7yjJfc74Bj42ZCaT9uTQRUHwBP
2S8Zd1eDb7TCfNrIvD7PHgRn64yC90JSsoyOozDvculxslIGmCqk8ffVLy9jw9Uj
iANW88BGyD6Uncgzq5LLoTLEMze7R5+jLNIJYlhXS4j/lz9rRH4Gk4ZYiJtz+ook
5vWaIFB1MJppmsLfLG2tV7t3P8JQ9UtMJyBEozvUvVpB/zOPtD5zwHAJpq3Zax+S
X+TsIaBPeJfi+hy/yI/eEFabfBA44rDJxE60cH/2m4DuPXHdKGAOtNTNO9Yr3yQD
YmlWkOG2l/n0lcaxPm0Qfut7H9I7KVnuCw79aq/g8mXcyv8Zp4AGNX7ZGZu05slD
06omlrH3aqaetkQm7t5sDhEqXmCzkuc8cxJMzErkri3og3bSsT76FQQaPpKmsJWF
VeTrqb1BquqrWrovjZXYWJdxpyeMjowuCPxXrmVMbMBcJz2N6cP9U6hIRcD7rhTa
04j9Hin4vlBhgHAbJBMZUCJ2F+DCE4AVy0UpOTA5bfhBuWoX/s1Xngh9z3Ofqg65
6TAcsPwZqgweb9BqOIpL9toFvA5mXtZGne5aP5uGyHmFvInfwZlmKF+h9m5M6HYn
bttnrPh2XxH88EoCJzvp089eb7Kb6fR65Y0YzmugPggUnGgPruzwQ091t4CD8zuv
EVQw09jwDmifqNuXyGPgCAcMApMVuOTA+UqpH4BgfHXHaItAqg4YH7srmkReNcYo
d9lEbleJNYXZ+D92rFDyH7+vxS7v6H05/bEouLgxAL0tt0YwVXciwqSghBFuAxIH
QJLWd5/jFpzSIjc7kVe+GFBrx0UnOg6eYFhOpRgrUEgA9IE8oHncaaTEWHxMnBAB
3xW37tqeg7wZLAexaP7FGQSiqmNUgAwVSgmOskWCmTqfDPBQ9fENkB/VG+QdmA4q
3WSNcAOoM5BwExL9v6MU6ocZc0KWBaemMJfXFqpnO6clDzjf7kC3uBuOZPm0MQwJ
mgXtqTv9peV0I55bYxk2jZzEospx3Ypws6341ec+4eQBkI2JS1kjBHbtMrAhC7Bi
RmcWMYNKG2HyzFxbgxiTQJgvNsNg6Lagx9EkWJCB8GH8RrhpU0+daqsdaAadKbX5
1DeilbzkagSzkaiMi+JZIgZ3QO2eHEs0epA/QHlU0oiJtYSNn5jJoAY/GtGqXSyP
NnnrkuxJrOMgTVscziduwMRdvSHhMXJzqZHZFtCKc74FltWs+hT53kW9cFol+b/x
SXqb+tWuhMDav6Z/yWY8BmDfyXzUqIB4WZfIf7/OLmGz0HmbSBQuAvjNAOXp2PTr
enEkg2VwjRTvbbXFBwiY+f61JlexMy7SPj+y632kM8SDNnDK5AO4jSVjpdTRjwD2
8QmxB5kowUkUn8fxRgBuafcadcyMRI6Dnm67yFcsY8X5dyeaQpcg+T3RFOiKQ18+
YE+goz+zedwXNF814T6UbVTQxLsGPaSv7cTcBhiLnjyFN5U6O0tPPgFEqCuI5MZr
iWZtuGd7ZN8sDbt3hOPO/+1nGQFv06WQ4uBKmN6Fq2cDXwxR/FRJKEjPD7Odkfy0
HXfcOlBRb7CiGolBa827kqLOcMwaxjxb2hH8FiM10t5PCCdlWKdEOUb/Q7sxqF+f
mm5egWBpzH+AIkBc93NGKSEQM/dPVTzJs0yZNfkX6UMyKY9sx2tCejhcMBzYS+dV
esa2IoTQ0uhHVKZSJBglNid81wXjdYJtaDTPvnkWwSmY+jGWE2aVzotIaMMGPduE
UlIgbhL2pBwYvcUGxr0rf3yMGk/6zxES1dLJWMV9UNX+pbLYuFI5wTApOOsAopZR
0A7cveayRuekOzJsdvb7tN1XgHPHuMinE3Rc/vZwLQqqLa859Cp6V0IvpIHajkn2
bMr+nYE/rD5dMhDV4XtSVWfVI9RCdprS9s+x3XYIsMIUkJLz8EDk9FX9I+bWxLl6
X1I3swcGI8pQItpba83u3KRDWkHehG+ZVmhkYsNGRgQB/UAw9wCFsraGv0hfzaa1
xIaQxECfmMDJXlwjseBymhC7+jyOFCSgFQefgw5vp9esSbDek15SxCQazEijECvA
rFq9jee1DMuP3u5KcWTPDZ8gZvWZ2KUdkRR7Sxb+DK03APiwBE9kUOR8/JMyvf6/
jcv3lMcatzVa/FkH4ubVaSrEUnpWjimcqGiXFPixbYOSEeKyswOqcsXbbqQwaQGp
j7i+IaVaPq9sU/xh2jkFxDQ3WsoNqphz6OMBNYnEH4JLRoxCtXH4yGrLkkNkL5dq
LHRBLeFHB4uwB2u/eXrXYwOAIl6gtJY1CRFqHrUqlEf+NcyV0KmyUcAV6iajRycK
Gj4JxCHZZqbNtXr6bmw8D4pLj9wTi/6nHN8D8RyT/0rddPYnmr1rIpszy1+Rv9Ra
m00l1kiB3iCP+omSYBSTtfwdEB3ob6TIFH8K10LE/osP1FYv9qzgYtlIz+TTGI9u
IASO//bNsIV2AfwI/eYg1i+IeYaAdolJ74zlD72l/FADA+kIF+QPUzzgKcMZzUsg
aGcx4DEQRHmYHocAEcMOfdcymZioQbu5azOhcAkZcXdRqyeEfXaPsnc182Slm6kN
g08nM2jyDx18fNdwwmTAzEy1/jVpNqpff8drfynA9TmBUI8a6XgyzcCMkEDaYRf3
lAPgIqIjQ7Uw5CdD/E7z0di5moGX8XYbmMPGlFmofifRA+Okm7tcLvIhn0MMb6cq
8ZC83yZnkUupoAs4kBpMC0rcddQAaePSmgabnMZHKaAwIK4FCQKbB/+cTfcmitBt
gUa7chKnX4und4Idtgj+Wp+yBW2L3arqs0daxPK2XuABk+07d6vEc5ffFyzmI2B9
gUi3VHFoZphQHtkYY/oLgzcm6Je0wOLebWXsunUSjjSF5IbxuJFvEi6tFg66yPiY
udlBMhKCxsxboQOz9PJVl8zSjxr466Nf3p7yvslUpBMlGLxpN0L51QIyJ5FzAKls
ggLoIM8zLT1DnDb/7jxBsacXYhaNdwjEtCcLaRwD4leu6dFhdvuEyE3yVhXH7NAq
m6L71M3revrH30tMuszFWSPNGZHvD3A8tfGI7bIoxbbnDhc0bBD7XePhcu4Nq87p
hdMduB5IuFUSYwdBEKwhwA==
`protect END_PROTECTED
