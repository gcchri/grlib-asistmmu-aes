`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uy8uTwo71liZNqzBDQriWyyjJD79SJqR2NfRk1+WHJLka1rn7wR7wskqwfavdWJp
rV1VOQwpWKLI2OUSAa2TFEFw0eIDzS/JAGsYjXWzaauKYuRNqcNZnssOP32WAri+
kSHV+gHShQ/fd04F/2t8omQ8o96yY5WwrTK3POCmaUa35zQc2k7IGE/1rry0uU0k
3zxdd8FE1bYZStsJCj3sKmKOgsK3t1QLR6OLdwt8elq9W6GYurDkMuAS3kBpe3LP
bJBEv3vjWK4uxCBiai2jy6WVWswz1t8lkzBM8Ih7eh9KVibLYkQo+FfcYqBiT2UW
FNOh7rwLIl3T3PhK+Zek92gyp9iDn+WSbxG2zmJHGEXPMUNM7gSl7wiYaiOKcaW6
Xmi6IphoM2H48UN08W6JHJZReLMyMjV5o6CN4+F9iphoVNvF/FyQE0UeZ5/sIMfJ
BVroI3Aw7cgRKxsdcd4Udb4NPR1Qit7VkjZcPES8iy5ioHakInxINvR5IdxZwmnl
mIGRlNxTtfirps4FVTPdvlD/Lko4tQZqhZ1IdpppMSI8oYH0Cdvlx6Z5OqXWsRjN
AraiYOwuxHY7//mU7Wttn7XD+0tgd0xjwYgtdolyZvQqq4ZR+g0qsxI0g7zWagzN
/n7Cf2nbuZMOuV8SHl3efC2otjW658yly/An9p0+agfjIsFVXaJCXUCly7xDRC5I
UQiVVrVwJTgmG964t90lU8jxFPbiBx0mxKlF7YQhapOowvl+e/rR69VImouKqnFU
U+64uKladSZK7SVAzCu7NmGE+OFRf6Z+QljEhtOD8FS9QOny9J76y4dP9w4Fr3BS
OPCuqX5NmfzXBx4XzGCbGRzC/vgxhCgy82dZEg4HMRwzuKLnU3sEVhOiCl45RBsv
Xgra3/l4B5/zkjPRLWTWTbNRYvo5deTrLCkQR3FxmqHlkMntgZdUE05BObqT8awY
VYIYkbFsSBdUQrhQLqq3vGkt+UlTXm0ecroktesJE1vGRdrj3Qn/1FoIDY1CUCp2
JUhSb51djIMxDwQZYVM1CAcVNk0Vj6rv0qYjFjaRuA22YY1M+wJZzBeu+lRnk86u
qAsNVhwHeSZ1jnFFc81TMgOilnLJNx6sVVhvvHmVVscnyGC32wrVmVPTsaiV5soy
`protect END_PROTECTED
