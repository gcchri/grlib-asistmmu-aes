`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JkNYJJ7+uFhtyyfTvbvQCUSldlov623QJx3EcegFV/IA0XUvgxuzQtzSrQR/4nmn
rLV7aWQHmDK+Y++PUQXOLznOVc/u9ulCWOo/hERONwnils9gJAjX7rrqbA0F6+31
hRJGniIEug/qGvs1L/LzRSujoe78Li6/JCSAlSfOjD8+n4zDNzB9D4cMUmdnFemw
VRulG70BulLNjpVkMK/wsZ+mcmcJYhn1TDf2kzkX/GFMlrEWLnK9ZJyAB8lsJS5r
5K7Wl69YcoeWO033+AtpoP20j2ctHgrdfHY3zc40/1c=
`protect END_PROTECTED
