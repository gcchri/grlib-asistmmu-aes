`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GCW4Ker63l1eG8CnbrciC6fNH/1A5Zriq5dc/gLQF8QBRZl+Ger6oDxpLH1YvuVe
QhkurVjlbP/OXbpMUSdB7khdhngIMVV0rtlEREc+XZ2yH1tBIhNR0mAueOm+BUGp
Wjt9qGfUjLRrFA0MzzMJ6gZuggIIZAwUlF0uwxq86t4eyeHXA8noQ2aDgis9Z9le
ywdyDuqTG+ZMaNC69hzZ5Kk2K5yLB83yIt2yR21YgxzJJYMsd69qU2HhXPpe0IRn
nwyKZD2ThIjtvG9PepWbwYi5QCRzj3xCJyJLAKqed8HlDIRv1lGm8Ai+sOWeCRkc
Rg8tgjLTglcwEN22N1E1eGFkAdnekXVAUJK9nmdxJfXL4Y3jGGo5oQj2UqJ4ShpZ
8JnnPxk5tqpY7FbDbsQEHOpy0xNgMFckddrgSdI2Oy4=
`protect END_PROTECTED
