`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WWru+KyjlRD+DjXfvATI4lLN29OG8f8YDrACifnkCdp8htaL0tKZAWbrE65pOTEN
n2aSdHqYCO4pcbmlOD36dcJf9DkPyTx6+6lxQzWlL98ZUdo++Rk+LD1TL+k8ptzq
KT+ZCyktMg3aI433LOG/+b7O8Z/uq4uG6YEroHqZOuNorKxbtb3TaIzEYpC8ZUVC
zYhcs9RHQPPBsLH1y4v1hJGZSlH3R64Z5NMmUNkVhPqbBIw9IxGl70QRl/tj9VlP
fSONRSz7TByJNZ7KvXncZWh79/yKuzkdNO0FvbGX9t61Kk96BMvPEO7ti6FEzhQg
00AYXmvaZ3O4qjV7CpD0YkZvI2nI8vl3IkcmBrzMS/VpVwoTGlkMgsvfbVWiKc9X
v4CM6trOxzc9MKIFEXETeik9BUOFtr6j7uno2amTkprHiKJk0VneBleRsSAcXF+U
UlPrlTbWeJuuaKIv+ypgl1KFAvjN7NXw5axOWAlUHnccs8Rzd7xyYcROO9E8EkE5
nMykP9B4glgcFWNAisKCqSBbQmmFNz6v4RHU5HPXTaRgyeWsfvP+125rBoolWgeS
D0+xa2zdbyjt4HB/vHQZDiLLrtv4NVX351fl5WWnKdevrtfwY7WxRKxNGHcWGESi
BBRHTA3Lc9L2GCpI6Lw57WwyEFsCNCPF7jbbDg1PdRaeR3U7pcYkiYgjbFhyXFPX
y0TxzvicfxA8IJv085zu4z/5SZlS5lh2nDFv6tV0943lt/NtgAijR65Rc9RdgA9A
/lumradhn+w4oPNOK2tKrqk1RxSvhGnmVlLhxdqPNcvPMCwhrBrnFEmeYJX3ehnf
fytoP1cTBLSjFqwO9rpMWhxp6SGvsnOCopZsVBYSEaR5tfK9ggoA0adWfvRhtbOf
r7t6U8iC2+1RjLTrGaziaXgAKrl85skjnQR3HxZ8427ylBTlw9xE0A5cJZOIaXvG
5Menle7pZXcfzJlm3GAlPQLauo3pivKQaQeMZCFpQrblqlR8fG+9ukW5aJdDIoO4
4sPwE8T/zjqZQXaZWgunzYezQijZHD6bH2J11z1XUfQU5svmOp9TM3BbN2x+C7hL
oXCPe/TfbAYedlqww2P5vKNRAU67kuszwAhVwqPY/yOt0F9zC9jxK44Lfbw4yYUe
Ukk7rfNtQPdp8neHK2ozYDMRBKyUcYO4b67iuFDtoUER2sEQNuNRNskE0pB+yazD
tI4rG4Mv/XY1X0TajJHPGIBEmOKj0ZuC8MxqbCYA+xUvstuDxHBi5ImKwtTmW4p0
`protect END_PROTECTED
