`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d158gu3NjGcPEq9LFKlpQu7kqH+8CpKIrZtisIj/jNdR00zSUSbPofQwuedOSwAD
UWM/x8Y0M4zQS14EGKsnVH7MYQohqvCpzzUMLjSltVsQ2IeqFAIrau4nP2prTFbL
04bDUc+bsUtaDFOHKQk9du+4NDs2CUVsO/faM0FqLaBJX869CwXWd6si9Zk82xd4
aEiQfK0s7FTC/k9GkRqNPI61w+qC5rpopOouspTRgVh7WtL4PCeJRyJisoOByyZW
riI4QJ/OX7/Z3QvRMQ/K3fQFaBBCRI+v/skXqS6TwnaEBUa6Su1Iqb5I67MrHgej
T2bK5dnLloQC0ZVnOP6z9w75pMTKirRG9OMleLTMuDYJP/UJ3MuqFgSUvuCW3aWv
+8lcOQ+odwKJBVHYaj47To3CoYLesi8VMscrW7S10dRwJFRXsDVC2v/DsqjX/+q9
3zhDb73ApSoo2OGfxqSlTYhpCnSBnahsj7hpG+eNVCE=
`protect END_PROTECTED
