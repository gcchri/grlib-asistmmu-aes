`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PNBjneyBvZTWeFJq6xbbqFqxLkHEYqk81+gBHn8RAyqCHz/CXByMbG0vL9jTmX3A
CKJyzLLBUsBu4D4lJS4+4yiUwIXBWFwWEsfFUiOrq6JwyD6KUhwkMKzPvDjZyWF1
HGFMWic8Ynps91ONEFlD1ZPZQFdGQprq8g7MfKGEvW5/vZE36c33RCJaB/mJT1U3
UZ+5Ae1BaM2ox8/hqpFyZhnekzcJ/09I/0k0DVmdNdDbmkjVRuwNVMBgwjsAHZAP
IlrLfashsTWVUXz9y3fd+w==
`protect END_PROTECTED
