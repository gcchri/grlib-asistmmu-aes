`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UW2Ucx9qsyy0ToUD22HxDpc7wiWH1/oeqMFaYKarPi0HspQzDYOswdcaH/FUEPzW
e8ur5//rVIc52cmWwc4QZMJ/M0Qv8gDqMMKpAZWouYoJ4kGSgklotnwm32mDBQCS
vThuUcUYOw7ASN1S/JLm/IeEIXxHzlU7FnK8/ijc3OcaCNGV1yuvvOpn8Aj+taAq
RUEpfsRdBSWzmcAzY/ReKnzW5w0u6XPWBtQ1sqwTZmn0e2l9ABOcFEBYrngRaGNU
s213qMt225vzTKfcuIqV6JFuiZI0pu9qIo0H1N+XIfGsRG2xKH87P9WWJeCo54Pq
TOFOLWsk4pc5htrDszmiiruYVzIPeK09JJKgVZ63RvJ1Sw5PpDn3T42UWcOrUWy1
9Zz+9XMGNXmVh/CIeo+mGadDHd6dDulCmlJXwIKpVLk=
`protect END_PROTECTED
