`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XMFpyVGKdEJFoVz96ILTWrbyL1QDPn6lF26rpiNqZzor7wwtK2Hsj8cwpBBecl4X
JKoNjGm0+EcYVEA0aCLRvb7yHfBkK0N7MDHWo9kRjWMokYm3M/vCP+2RRo+svGYz
aSbVv5CxE9U8vOJIW3B64bTn8QrPqarnYTqQ0ExBrsLq0c4hJBUW1nMq7WouGFr7
N9m3BA54mVK+I8bR5eUcAhzcinXX9xBMCzWiCBu0FC01MkGq0U9SMCEyWR/mJtgX
7nqmeHUrmfv5onAxcPjPVIeqbtbHOU3rzdZrhXJyj0VBoYNSw/LRvIp7QOww4JYL
qb6VkZDhoD1xsyUPY8jqIw==
`protect END_PROTECTED
