`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8jkIo5D98L34rxEjcckjKBzZHk/bKaHUYMbvVsDsK+i+sYbornKd99vqF773z6OI
Iw09+5M2smXfHF283jDmiaIdcPn86mtg9cUL+wC1LMSrWAbVzGVKVOvphjwWvrCY
mKNzTtNNgwXdgPChw64Qg8aWYxEx/+PnSsvGjV/TjqmUkANS4iJB2brVsMbT1Z4b
F7qQg77s6zTxbd5Pv16Gx6murlHSmHmPZuGysF9FJ4C2qdgjYLQpPTHZ+J3qEXtv
0FvflPyMINXjKWRAncad8nJQjOR0jfnGZJD6ZCIKwOAjz4FE43AkFnFm+to9G8j7
mYgSsdTtKnYfl3TOYbozbVETDTJXPiWwvDX7rF79seHvu1ruecb1XB0G4NWwMATT
KN9w9ijS70qw10TaO4ll8rVIjj/R3W5NC6vPMAvUkjXdUuLs1I878vOQi9ZyLEHx
`protect END_PROTECTED
