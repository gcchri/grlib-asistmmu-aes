`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BvZTWpxTxNVFSyndXEMgTxKDNxIsLkcCvgZxJX5LJeIhiD/fe9pFPXVHxAfJtESJ
kyNdJSMal7JYHlGVTP3yDYPSw0ye8GgF/gZlPSlbG3DdjcPrqv7EdCKFEM4UrVVo
HerxyviRgb6OGxSfm+RtC8O/XZ4i5Uly3aTDjlRzI3fqRC13Fa3diRdXTuT/AYaX
Ra7WDI9PxqtVW6AgnCBGEfh4yOUqS3/hI/uYPieQKVYk+pJ/rFKJtWXEkQaNvyL8
jpMIVvb/yjovUG4k9ku+lVoTg0yN7UydB/t5qNCcVx+t8vlJkmngE14jB9K4JBPt
cjHEm1NJhLFCODMKseVbKjXB1+3zunvY/WRtlZAAapk9EtWOZQwev65aOPydXUtv
vKMAN3OskL9EFPczzxaLaEraIH+gsktn04YZnn0ehqm3wJMPOy4WzZXMx4BGuVeu
ce+wbpBnVESby/L7r+5Gg8J8+di4hbhkkJ7o4ZU7xddWx7j6G9AkXXzbg/vrrinF
yBlEn9yAR/ahaM0hro2+robSajlxT7Dvxtd4UXy2jZtmJxcthy629F48lepWXDaU
cHlFT4FRMCOA/9XZnABKRhviuSAg1dYlWLVZexCvvx15YmNdGNonzy10QtHt8WSu
KCnW55SPTUp7p9zxViqFtogWVdUb35c6qJQeZ7fYTpAzfAeHV9JN7Dkph70Ky9Jn
czdCtCupFXtdKWf6tfk5XUD+U6adFnO9feenaYGJaSKp7wty+8g/z6F+nUMQqsbt
`protect END_PROTECTED
