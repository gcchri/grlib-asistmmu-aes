`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R54rL+98clUInjuCYySgeaSxiJI/XXKwUW4jMDnWcifbVyQp/24AVxKUw+1vpeoj
q89R81ffyYuJ4ZdjbBMf8QLnBaC34mtPz4tFQYjuo7IbnpF5bSRWmxYTU1ODHfqU
2sG9cevOI+HiD9CQkAi/+5wBdzWSyyLIjil1c1yXEIqleij3C/17V2Z2r5w7VtG/
IcmoBIikVjrgBjeHQkAX2W1uI9JtcfGD9TsZX2I6fd5DHAwkdwbDUJYRnc0HPwDf
vxH0lQeSnKpJLt2hu6ECzr1XzJ8WQ8hs3+IoMUcyBnVB+B8W8F6ECiNDQc3W1lrK
rrUdIxhAQBe9Y4EFRqI7faU3oziqtqbVD1gi3Bqhm3YZia5cdajcnaNPA7KT5rgg
XLXcK3iE8UU7QFE+rOPccgZQWRGcye6XJlI+kIgFxqc=
`protect END_PROTECTED
