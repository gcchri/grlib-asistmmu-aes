`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xzr4CnfRQ0rT56pi81TlkoOb7cMrgJRk0OoPoPp2NkDmn9QflJG3tb5QgYRw7cRi
hAdo4Y7YgbILM87Rf3QglUVKc0FvATWsMi8e2kygYPRHh75sKh0zxENZ3YRuKW2I
4OoEg3PPHpVL8G+a3KHfqKcG5n+1LP5fdmjWu2AuA8zzFHjAU9k+UbAtuFhzr1/T
4DC78PDZQArONEYPKSNuKJBfPVfL4/XkJd6DUy6N3+bN9c6kZF8QvA9Uyh/5l1WB
uPiRJlgQDV6O0qpqTvjBIxMnkZlSur2XKE9y/Zxt/wVfL+mEdbImX3fgOM0uT6ax
V28taQ3KdouhAGpDS6TO3cF6VSiKuKd5dQIrPn2AKOHGUogUCvBYd15fOe9yKlQ+
XPoX+1tnsLfFaM5Tc4LCufAwItDll74NzOBXZPzqDar4CUNaRL96rgx9lxiPXxaT
2of/Bbe23FUvNrbMFgM/1ZZB/8CH/hByaAIi8GfnzGeJOYPf/Zdnz6D4H4fEAYbe
pfEjXqGBmxs0p7YeNyfLDRt6EDN/4AYfZ6IepTgcfvBD5o2PT+VmkNXTrOv753ib
OFuROpW5z39oN4Itg478nA4OwXM4A9njvYZ1HIPAt7yTS3Uk2NU2ZKlr3lZ5bgkP
HPfVpHXKzkW9bmM7I0lH/Gov7Wm6RltTpDR6CpUB8Dg2Tn65Nd6SgTfIuxH+yL2j
QoxsuCywUCcsYkRglIPQ8pA0axnnFwC0vD/khBZR0u1SKxepQNPb9Kb66H39ftpN
q6e1BZnlt2EGc+Si8JjOTWwT+/pGDCBjvRtuGDSLKhKG6MchIi+vV+/TF92SA497
1YVG5cuLuNLbbe39dGjiznw08vLjD8VPO1PwB+vG9deu97esovNz6adQjceT+aiB
qGxUiSXD9NUB32moFrLb5ifePJ8Z5XSyhz/dmkgoCoTEYS05AtdMelBm9zCD5Py+
0wuVE5X4lDgwucGyWm4AJrjrJGbg6EwTfQ+DjqQMWIS8DJT6/Q5GlqUBvNVe8GXq
IdVve36SDgNKNp+TvN/NDV/7P+ct99HAGzJ0N+LnOZqbsEZDza3GWZ0hPtelQqeA
RSoq58ecFc1C3NeRWO636ygSdnks6t3bPc8mSVWN3ASqJlBRwSJbNQmqBGD1mI95
DlNOn3kCPL6nsrM8SePNVQaSs+CPaPOsggFCnyAuFvrBs/gnGfZJkjtPS4Q78TSX
4Pmmea0An8SWtRe03iYiZNMarhxG99rnTJjgK9c0Q3q6Qud77pdOyhxpJhjI6WgV
zAQWIiRxG2QZ/3vRCX1iVJQFc0Im8EDGQmNgkCmjrTz54EizNNc+jCMpuZUNHMPW
sbAqXTdqKcOG0B3SGVpVCxFbpWXujnOBWo4+UEkVhRQsk32bPi+63caxtsBUHykK
EhbgD8mVd8yKX7msHzz/g+U3qX3azN40HqpDDVfFKPOZijrkFtud4QFav7DLC8cP
nEPpl9y8UUfDfuAcsQhGDQqQ8v1+o5FXv8L0S79OMB1VUnxuJDTqseR2oKt85AZJ
nxlMlqHrkGNBlJzjg+FXyrPLv3gbHxV3ne/KZH6Itc0RKhSgBAdR1HwHc/xcPIvl
WiTFUEoMFcalrVorAvLMGFDyR8eZzfLGNzNhLOqe7B1/QHj5IJr1NjV1yhdGWr2+
yS4FqV8q+taU/iLq9PA+GUc3D01T4dUrv0Mp04FWw6ZGvSDmem7SDhePPS1ook4u
17NjpT77LrsESmhGixeBo00KCBvI652cabc+V7iiB/YlDBPcWW/hClTChPww+cNC
PzzNyJ9YA+MFxtzv5zUrPimOROKYMgN/dxlLF+yJREK6c9T0iKFkmJoP6vmeZPnx
ztYByiOGIfm1cSjwxtQfuoqyBeH2asa/EXObcWXi56Edb9x3l7vVXHa55lSjG1GJ
y6Y9TszIITLfeALaicP88rZgP12SjpNhQbrOYNpJTWKpoSCrNYCzaGP6/68YhEyS
pdzXVL4K0+b9WR+nrrwgcz7b4DotceBlAqLpgY5k7aHdtZ0x2ktfpRgRnaiV6wVX
70ozAqjWITeeNbBG0yW9LaEZ/8RZ0y3hr/wSVYW2li6ViHgRm+9HLmyW+/3W6Jfu
vO7E9wVAmcuYnFI1jZWWvcwsZrbJe8UwPX6LQEarYDWFwRb6BOnD8D36fVppUHgj
a16wka4s+z2VDt1n6lvf085YGy4VkeOAj4n0WJVe2UIowfyBANhFlc6+FFMMislD
99Ezz6rmV9tn9JCD2xt96KnwhK9cbPadhsvgmvq3TdguNdzdKSLJXiDmMhVUAnI6
gtvrh8/6HNwqbdu1kx6LtW21bbvygX8kl+9uDVzfdKCzus6G1I8w4FSRssS2XqoB
/nfy1JrMpCnV3jtFzT6LFvWRbm5PXFd1n7xcKbEIp1GXDwC/vf69YTHeftkXFip8
1+a9cKF3e388FOpaDcdbJv2oJVmUS1AJ2vcc51OhhwLRfOByUFcmjelhSFoE9GTe
IDOWssM0w3UDWXuCgRVIzJWwSz8V1/ovxu2aGK7W4kng+liAFjX1BnTxNC+0bv+7
dD35JS1+HDhdzDXxRHhpmGyvP9OYkCqWeQ0DYxvZDRybOpvzjn1F9ClvucqILEAV
USyxreZHAM5AF5RCM0pp2tlGoqHOvEpB4MDO9dnOUBfx6Vj5LRhopwCJk2Lx0rqk
sQXYhyIOlf4RwIWBMRI7q60nkyjsGCrl3dhyQ4c7yG6M0AcX/ab9yuIVdcy9kORe
0BnAz+sGOxeoROPIAwkSYLM2BQCTty8+KYUnRUza4SIzKgPQBjTaQIz5uIZi7Y+W
AHBwzKhEIGD1NTmjkw7abcdMdoHKrvrDwpAsEhkcuPS1RTB6bo2+zHf1msbzLg0A
cz3UCR60GieRwVM2xqZR72do+wrQ0QQp545VkFqxmrnRcjjQlt0orfmN3lPwiATS
dkQ2/dGE00PX4ukAgSZGzCTUEc0xtTponsnT1qpZ7P3NUMqLuRsSnI7OMI0fWeoF
cwm1wdoolEbBMQO6qGCye6EpIk05Jj0drAiIgXBne2IjA4vTOmkl1dhhVsTaLy8z
pkqGiR6nE2RWy8xFAbSfghnZftTFi8jtaR3tLFzc45SFaMC/lyn3w6OM23DxC/Yc
9dUk9Cmwc6U6giSib1wsyrbatoCZHsDCiHQKxhpH8YSAgNdICjPtdjzgKomsAppx
YEKh1oAJwLsnZY+WIn5lC13+Js1P361yL6TE426t6ekNuxTKyoh2N4SOFVTfz/38
Arkh+Lyy6Oq9HHEBTeB42t3hHVd+h9Nd11NSBWczgKV5ThBbg2nzGEawa6VNja/V
t6f3kD7hoajVOUDJ1bDl9Ld3oapJk3+nxsCm6nSurYJfVjf1Yyps8RykpNQYaLgS
t5gpEDwmZNnPpDpLeqHJxonXw+ZVxj6fjq7B6w2DqlqnByPVPgI5kD2ot0TXd1aN
i3y2D609JxwLtktFRti+oovp5Wz2pDqH1+kk5fwKpm06kF/O6AU9ePwBMzCkAMNi
OqDDkT6HPNlX+D7fT71lQcRNErRcpuUc5mLxNjxdhV3FuZvrmhJ94QErJ2jr/Vrq
g21x6L2XEfS9Uw4qgWMBd7Ni6ERfKjPPeHat1q+6Hc8G12+WbbnbVSgNN7IB9mfb
1ADj7uWTcwJqINlxSoHDVGWyZ0m8X7tlMDr2weoAGeStsOhoVGgtHrTGH3dDpRk8
3yKAcS5hg0pCLEqfeSDk0rhpjfdktPyYkV/KGKhB7+XWkEWaf/K/U988goLer+Pn
b7xNfN+cv6tHozWPQ233l8dhiVjU5Cx+OpC4twAFph1O6CiuPShQj3PKzuMdQIiG
4UrXmg6wwKklbVnc5yCqsWrBUX5kHHvD/PARu5vCtlOUt2Mkn0EkgLiSezv/ANtQ
eeeqGPgLbdVevw+kHmpr9U3Q1kt+Tgc+AWuObXdW5yctmLKUzf+F0iyrvBfhh2//
p6mXOm1dP36rwLR5J0m4lmuMAsxoDTN8BvtguiAXDCwlCF6wvqqyeUBNFkCl1NOZ
D2LsLHt+xpUMa18gqDZmVfeAq5nnPvo1wuAI0hOmk+n3h1HWOwfSJ71uES00fDts
nUyLytmFIuecatVxHbvjpjcFi5GwqqonRKZpg9/nBi2Y/UNcFO9SCD8ag18CcNFp
USSnV2Dw/14AelrMwALlbTwgXQDG8G+mhQqjG3J/KvRcXlE7Uy6EnDy4HxPnB+RA
Ja5wibdOF0PVNbxy80TeNc5HhZAQ1V6LmJX20cvBQlim/jRBL4EaNlltpdyPDtNK
EWdapcJWV4BZkMUiImD2Dtsr6trDLqrSPUG+1pyJKdhpBFwKTjVr2cVyMytLwqD3
cKNVHGwQpgIa1owrH9wLJvmkZldNLIW649sQeViM2rnj0rkzda0qxT4H2t3N26+h
gsz/9Op3XlVEanG4fb9x/+T+b4NGFkjbkT2avmoG+Mr7YrHPbxU78BuQbRPEW2mY
3LFQreHPqRgX+c3CQUG2qbBvnzcktX0gteS4XlMy9yNJKD97fq3YlsDuWLy1Wkrl
8jMcGi0PcjMcmKdanowi5ngdATfwVfFNVisp3Bpu39VyvxOYhmkRNYDEnc7G5Prq
gc17ZP5o8PUq045Kp5DhWTyNRpIusoeJfJt3hV5CZ92nnpzqfLPxUT47DFxKgJjO
1O83mKg1ITb3UKmi01woufS9cHfFlJzlNUWP4tKRGZ5H0IIxpRptNRZ62u3ekXza
d5pJBgtM3fvS3SZJFSez9u7D1fJq3sHiubdtApagfI53clQ8dKhIoF11Wlaw5l1M
nKb1FwSHNmJxAisXFjLAdIQPYfM6SkUyzLtwcETkvtLAsqnovwVmfL8ndypjmOJf
9roNIWGiKpoaddob8mEocXeSOcLtocfGeGCH1a4Nx9iJRJg42Thd/TvND2jrxL66
IDwHHenERKxfL1bbXz7f1+aA65aR1laZ1Nc3i2mNofAV8M30syaewI3BNusDafNk
R9YMt/BwQsbSs1S+esMCYy6euoJIZ+JJEirIH5YsoGzSsq+fLbddN46bfnmL/CNL
+UZZdJp8uok0uZQh21GI0wkg8JJiUM2N/0Zx8yULmg5K5Cb0z+GwdAOPNPFxqXQV
jDAB72BxpjwdN1wkF31+DL9CPgjEjpLdSa5JxvKWe/OWj1aDiKqOdun19zYMwAOT
3wLYmDJ2JKgWgN60glqSZl5HqeKd06NMH2xKZrSNk3bkiMBxLAoBQnXEOzXMZd42
GGEhCnHDFihSUh8vlnZYTrE9pfYy9l7vlEXccH1+DqgJ6STvHi9+t7mGeLOjN2R2
OrzLPrC5UhLR9UVKbdu03NEWmaexSGBfqu7wYetQ0RCMXS0eZSAwlZOslJ4PcOfy
eBqC5L/Whbk9RgGgfeyZyI+qSEaeLhJFkDS42cm7WHKfhq3cwJXoGAOUc/yCpocK
InLf2Ty8IwEHYuSmyrKCBpV53Bv164UR1cLXtArnEeAVSJCTOCEDMGOWB9qVPclA
JYtBbewPyzevG8AZz8WIXaxEf+mL+UHhQiYRSXlIyWOUfoO4ISV6lqjf2U0FD7TL
Yn+vDxGaeU7tHGdh72XQrHEU960ENAmp9t8yUhev55tIk6ra3vWC2lSv+XFwWIqW
CzTuJGs2GUpAxR2+PFdt03YDBF+Hj2lX6SmWE77mSBO1WlBndcRc2IfhFms73UVR
WJ0DoCTlm7x3PjHAwWcxBe/28tn+x0cK+bK2K/SA6zsY4a5pYiHBAJPtgLWxRQQJ
MHeYLiOkuYRY1dIHmlxuQ8kTlDnvTX4IoHSNQIDepvRfwA9lIR1dY9hlelwjuDFk
/RtZfJImhQfA4jUBpM2gg8PfQ3WP202y9WyfmoiJlQvUZCdoXdJMDAFdvlyBZiJ0
4Jn4Xft6ShudOiu3I129Ykkv8wZ0krba+7j0a+qFav7BzbHWFwxreec4bwblzlwW
yf/sgFhwuwoXs5YHTR/IvDvITws0nDQ4w5dGbT5duf7URUbHhU9Dvlsb5ecJe315
D0pgSzXRiqvqHfOS2tA06fUsF+h2fTgfJRnzO4p8k/UMtOYYbIvZYI+eUW5LaCvt
g32eRNuOFfluIZbO7STOX/W9wfROSEVK86UalOXkjvHVyLHmAJ8orfkJ9ZUDU11G
UW1p9LoscLYuX91MzaVnuEtTF5bz5kT5dYHVv8MZxbxqmGhy9VClprkqmwWmGmpe
AJNNIhQMagPQewsUp9neYEPV2/2M8G6uNJ8H60aBKDemzlHhejpk12czNXEhDcGG
fpMkTeamnY0yq1Lz4a/WLSfLfjpOfZaY6kP6JrwTHEVflkX5+Q+tDGjF2X6tswxd
31mm6YuEwuQ6OY67P7tWXVrWhaKBYLfLDDp42cpsSS7MAKzBUVSXgTAV9v8dhMbM
er4wQfwWf8KteNmySa1+muBtf3mt+ZY6OrUuxqlAEhwC2j1DpZQdBZ8iyGoqnYHw
VR1KXFq0c+MAdJsQRR2X6abyXtFa8Tjdmh5+70IEYOGbMz2J8qkb1aDboRu4cmIA
ju0CClDBZzFctIIitsvGrYdQ/LbbA0Bkq9iATsuGogh6K0/5WSUw7X+71yV0O9g8
gaqdgarPpGRofdVYEWiDvMvMyfS+38LaEMzT3UVO1iqFj/AiehlAGLWOHdZX3Dma
MnUJYOvzzfRcT7jM8Qnc+RgMPZWE932g9T0chLEI7ALpHdyyo/YndXccjU7GNvHa
Wewsdf9oWqploLWkkZUcYHU2KOhOcVRg3PJdFafPwecU7mRsobodif/jNrbRuOT8
8jODOc+gDPegLT7U/AK/7G9CwNCbVso1sMUaxiEND2rn9v2ZtABY5Y3iKcSb12oI
NetymN4sDph+sXpHIhEXfGVpOZE37yUF4sb5hE9UjyjxAIoEo1JduVRm3x8JnfJy
OilJe3ETY68v9hPAUNxP0qXnSDO5ahv/Dx4AK4YD352KuMKwIR6lFrsGOfadAufQ
IkiZpuLRXmwJi/Wqicch3q/Fhz/Bt1mwPil9IwHjrUMsAtkETrNjO9dRr7n7jFqK
`protect END_PROTECTED
