`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mtspd1InKrK9aa5Dyqnmi3UtQzDU+Xvq5/UzgIsFHUrdl8y/RtiVemHhOsyf7bK7
ZEfQP9znNXelqHp8WQEkUqtaFZnwkChtlM6/WO4J6bsZ5PEbXhIJh7nTuvH1INJ5
iv7eT0a71WxHqfdACAuKzbvS9OY0fPcAYvAMJX5R67zRTqssPiwHbTpNcMEP/KW+
hH0aRboYg3wbOpHE3yW5wdxQ+7ktuVdBsdh8IVeS7YsxHYd0VM7qObtmyBIv1V1V
INVnVk86SjfFI/eAuQCrCPLzwWmvziEwg9czoSaDchBE2IA37LzZtdZrNlg9kzRD
z3vZ/y07qiqO4eDT4pergNsOTZm14D3+6nu8L69w3Oud5PDqnzu7LuhlSrIE4TY3
JQhBKNxyJh9WaA2wopCnJglX0W1kueviBhjSbR+qKvZWZteSbVKr/DXHnCUVVqvG
Gs1UJstxrYcCiT44FiHd96S/JcYXR4458OBNtP//JNzLG2G+9Z3xteCGGeG8sDtH
OGfqcmzG5Ek3yK5JW0/EUiAFPtdLLkRsUrfLaSaZwofN19NVrwqaZARe6qEHaBzM
10fdPlEEvyBDLSD58pJ3VxrodwW2EEGIyvo/EbTI7F+3u5bJF+MuQ9HxwFejILRy
1B5v8cqnjTBBc7me4BzS+XuFnQJ8K7C0+E4xmFfwI0a9+SnJZCIccShR3sq/r0dr
gjm7WnU4+7ZBH+OQJmywQRMhJx2cB5W6OGJPZYeH5UJBIzbDE6PtqbJK93XW550i
TCjkVXy7QMXCxolhzWqWqy5o4tENPs2c7403nf/A7f8YMoWlhbYEGVbD7r9Ey8+w
q8Z/NgrDia2TAacxgTsG/A==
`protect END_PROTECTED
