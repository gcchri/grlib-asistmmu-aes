`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z9EpMMuRyseWiFRM73EnFl4A9/Ifb24Cpk2NqKoilzPavXJ/dS+NwaLF0Inqr+jd
2d0NTxTZymXnWvPQswrteYMnCbj0lif9G94x4np4T4taI0J3PWXf+U+WM9YK48Et
8wViMb80YCxAFZV40CIx5Iz1ZmUFvxAeHXPCvKCu9d3qR+vAWe00//sHt95FFIJQ
aq9HJvtRqFgPE/hz/+Auzle+cWRFJqRKs2uXh09JZTaijkSWC4Zamz5tD1vVD1TH
1MW+maW3FV47fGt8XBOXMjmTkzCrJ4VDt2L4AIetaVxc/aCvupdJtMKMai/hZhFU
Gh5jRgfUMFVHGy40WT5s17pvUyDEppHdHC2Apu1zCwnza1KNHvKlPyvpEdKgEGod
TDjaIF/cwllfC9mnYPlT05Z7lWNKzn75Sz4FzM+WyfGwU1uqUvKko6khdVB0vTlB
O7iQHOFYVbcOu1B2DofQbOQhlTgh+QrTPuOz9u8LwjdJq6woUMZacx/d5Vot8pLd
THn1uiWaT0mcIsffz5aISeF8rRXmngvG6ZnbnNRunPS+NDqnPm/hv3Ly1Rt85sCF
KI4JW3lDTtLjA2uOrxSiAk17U7HoFXWdBva4WWFKa8eFggdg15hzt82fvJRSvhKc
TVHH0cnJV2ySLc0x6bnuy2oClhvfBcvmUmBxFFOXEgzfDIAXr6VD4mEi9Wb4sMWT
YfPL7bCAIudkUyoPtTq9hXBdVt//fpWK52E3DjyOakwHBeX37A/rBLULz9W8t7ZI
I1CIuXmPCj6nuqQ6ciurtzMNCsLv1RjKB+d/KkfDY1D+N0HDDbbqkY6urZJYzH2r
NhrKVIRzt5PfQckpNJXs8NfB8vKn5NXed6ce5mfLFl14+xdBWZhs3U3C7sItWRXU
40wfN3YitX/SDU7HgDfNUs3utb0FPHxChW1Yfa8U4zBtLPoWGGR02XqG3Axy+hSR
eVdvU06Roc7MqHRRsq+4VQ+PLNafF6b3SBeviVPfm4bu3CR5j5Q58ccHk7kOhBFP
40qOa8gif1yWikZiibYgwCMHsQdOm0FAF2W5wx6TbJNw912Z/cg0emKt1APyNLe0
EuehsXL+mUWRphzamrnTevIGhXAwRYsToXias3DIY/MiwtWRoNuk96J2YNEc4CI7
9t/vm2YMfQ/K6t/dKqE+Dh7wABJhFvcj35jP2tRKecS1DhhU3pcKcMCr7LTvQdr0
p5amCox5xS6pZixoJaOriTk1Zlv7Z9K/0IOdCncMsa++CYEX0bGawBAqingA4kQB
CMAYTYjSQFjIuvtE/3+8IP/Rwy7daeWZm21Vdj0nQtBSUO4kIzlXPgvsDtpFzcjG
BWLrtnYL33FFgD0BqCCNT9wwG2u1iXY5DNXIRY2taRHQHwMxVBKcIWWYRssir9e0
rOlshYK1vsvRWPzxqQqdKekZ2w2rAUjIJaG8jVtUzviRs1W8Pd4j1ivosI3vjMFk
ymz9RJXwzCohG8kOBtuVJHMN6XOXJZ+50mbHMC1ITg+ynFUkbyY7k8/8jPhjRgJq
USOgNImswqLHJ5oDkQPPzw==
`protect END_PROTECTED
