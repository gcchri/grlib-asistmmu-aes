`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dg8yFVys7HEo7sDr5dNvIPohug+ctn0yn1Z2G/B6FskJFUvCEJPprByxiZgbtT2d
agFD9XlEJkVtsuYYAnQn9r1u77qFP8Y+zwV5B5sJbOtFAmRAQau0n/1QpmRmD+jx
R9UliX01HLs/+MCXLbfCPFnyy7Bsjwa+EfmkImvPRFUwNTDo6ipQgcmMnG7IXEfO
cUv/ijyY7jsli7bAHB2Uvauwc2lG+2+qdPhYkI9UwHlJaUp/DodSEEKUk0d8t4m+
tgsf94EUHymjC+VS/vnu5V1Iyy2EIV3S+nMRjbSEqU5untIfZ4sNVBDELdXi/LJ/
uzVjbanVzkYIRuj5bkyk4ZGzSSOen8h0q3hGyjgMEk1zjBsvF7eh284l5g/zt3zh
4cjDlMd3RDhVKEYNdNPzkIeIspndBg+zxtlN+ks3mL7KXRB9sgWiIOQZJnQNMmJw
mkcRc7jo/QZgBVKsPbRv4nrMrKNebMbTZgBlXm3rekcwbJd+XDvE7MaVX8UQa/Ra
`protect END_PROTECTED
