`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SKdrhO6K7e12fcsliiUh3s16hlih32Y2XK8SewLkak0yfoGS+xjPpJc+j8jLr+gw
UOvn007qH1TSU44xFlsUyVEQxpVxzqEFCD9pl1Yxe6l53tRz5WPqbJrecfFMa5gP
klfw/LwaHEQxJnuzuqjeQ3oQjrQTN/oK37p2FD/6Zle1VLuZnkYJy21oDiFkQCsT
4f63sFgYmzEF0k+o1foaAEgFTmrJSt45AmbgG1SKl8vJGNcodrFrAs1YUzCk3pOO
UDkRHNA9H5Fmhb4QNHVzFryFQsKZKNzyShYfr+3p7c5KlLLxeiRiQk5fA1A8iFuM
pTQV5S2oHcUJvX/HSvlRznxemc3blV5taxCGYMbj+t6WKGMuTu/iubkghBy83vZF
Z1es7bzO/JMl2Cd+zn0OTw==
`protect END_PROTECTED
