`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f6HVtK4RCE1DkXQVzwPBWL+zA+BD9/vghkYjhVisl7rwax8nPB0oDFP5y/U92nsL
Z1OsN29CMZUuLKJx14FD/Ie/JtaRhpR5vzy/AOy8bluC519I3s9j4mJSDjpZ2b2l
/qsEHW6sSm2UGveAxly3ZwMHBPGOUv2c+ZG3WpBTkXiZ8jSFbxVB834cSSimp3no
DwvYvOGXdEqsKOfjBDe6oO5eWTJLvzFGb2liP0qYdyX/RtSBuXV2T8Bwu1JmwrF4
Gf69MBW2cxr6k9tjE/IKdg==
`protect END_PROTECTED
