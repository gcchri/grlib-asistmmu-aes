`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Id5I7FN1Um9kgrSQ32SBMBhj8rvo4yHBj+bjZGCWWTNhERn6ttPqYhU+g5BvlfN
15eiVU9QLD0V3PfGdCBbrafPuSBUV47kYhgGk5zpSwDtJrejjAM8TcoMBNrj+Ceo
wtm1zMAboxAa6OApor87oGCXQVbQVOzxGV/Qe9dn8mqjVFFfjf7EDX1dI+PHFnew
5CagSOvfR8n6zgstwF7FxzJ/GUfIN0M6FWV90jRHLw/padGWN/ZnNBRm9REtR/zi
YUjPJSI06RaA1f+Kq+jxkix4T7aE1Hqlnu4op6PmSrrvOSH3hkbGeYbHZwsfhmEq
OYpi6aiL81YBqdqjOqRhk5zwEY5hPwRHbkmzbBvRGHhSpgx6TzAc4GlLAL9wI+XS
fxplGbZmUe0u2tJc27g+9MRmm0QvbmLqzVWpEJQH/yxIGOs9n94EC8UOaJnOQdmz
aazownabuKbaIR8oIEYi14opCe1B+3zaBcwFJLd3vOJsYyyvOVGrRfUOovdsHGiq
UVnNeJ3CvLc0JavwLv9KKVjIIyI/SNJltEmpU62zImLeypHqqSBBKCMaT51ovmmS
IN+a9LdcuknSLvQlUAoEB1fP17TEwE4iR/7HAmn+qfKcKqsIvjHPlJKNaFGTvZFz
iwMgY8QSqbtnKMqguVIACDjJeQ6AOc/Q39CYVkMnbxJlVmmV8//joCgBlipe31sY
cWIQkIX500z7JCec8eeve0nv33xYQeIbnbEuMimG0129VM3eh9+e0nSaJLyxzlvO
fc6bTS6XEpcgwTLhQGmyjrkpGXVqkGcoEQ/42FtoDBKrBIJGEmjTrzfXDO4lq51A
5WaO8D/IY6d85/E7YqgqmBeS46GUDRqM/PmgOuPABOU76uq8hKDYPVLZvN/DrOAz
jSfNaDM8vbEyi3UEKTd2FDsqy2Mk84n4igQwW0MkvNA2S0ttPaDVXlvWRiCJTjmo
wBqDD5PGSYhkgmhFLQ0gzQePjQspFr+UrsiQmrzIhb9TdxTreMfnnVNTAUfQlH+l
kxa//aag4oxoybxt0LLadKaK6OwscjV+ULxQtquOT4U4XWCLWH9pAHEZbrNCd2Gb
VfHS5XUViWbe5P27JfCicA5MnzRnvlvsAwQQrgelHj5Qe0xoBoOaZMd9KC2p+AH4
5jbsP+06IMktuLigNSuOw3wzzavvHVsaG3AEjt3BNmJtceixjT25PaxNnKb1QyhM
e3nnzdFyJCOmatzGfYrrvOnCiH8wvVS46FPH7vH0aOVVzT+STgXh6dsPMul4B6v4
V3wrJJl8cBRULVNTDTGW6lQEsVjBUHzq6eiVQziJ66zrKENPTN9S6GkCuE9FKYms
eOxEaqsISmJQ7QLRUQBzW6dpsLmss/kbGkP4vnAAfNKOG77x7Bm86d6EPI2kuISl
VirHXMzdBVxHGvRWjags+PFIVSEOAVNNoK14LtfMz/CvS3p24Tzp1MyvtQ3u/G7+
ScR+pe6eU4BeTDIQXRa4iwK+3Fhqy0lGbRG+iANyTXCX5VUGzket8tPGzPkso7Jh
4x1zaz1wmTGMao6HOaocgjpSR7DumqAXK7vQO83sjFdT1hObPsv8wKHDDAiBkGJq
VPL9wCFGCIo9Tpmn4h4nOyvVTDOkDTd+XvN28Nzdh+0D+6pH8ur4EvoUeA3LsiAD
ll3W8LA+ci8NRTEVp+tlybw/Xd/QrfqKqI1NHSNuzdnmKk8f/ZBqAmJL72mxRZiP
EyWrjY0aWHSu3mF6LycBdScm6qOjvGih3KG77tmKWtuwP4D/3dgpEzu2v30+8dcK
LG54zORLYMHDEASTGEIhxCEIcPuy2248N1AEh9g1bLHB6jcgAAM37XOqzJXB2VqK
X2H7Gnuc2sNPeAwG3sZrV0g2EhZDaoIMESiWz51ob4dAfr91hcGQ1QrtzeJMpW45
OPIhVmX5uFqwHHcZP9zSdX3gqSYnp6YtkCAeCwk/cWNAjnTq3hIvB5NW1NTiWn4k
OpzrO1J4Rihi0ZyWD23XikvKBVoBy1kT0mkIRJ2vwj1X0fdAE9B8exENXZ5sbF+N
ZOcTt4E7+wTntNWXQNDn/tc1g/OSltWaMbmQ3g9xafQyL/M+IV/XlJSOoMNKfHCQ
1hNFqMdeXDU7FNIetSYhDCtUjBB015Ym9WCi5zrYiyMLnI6cUB9u87rotOhldAyk
sHcJdJZshQjaKtlHxo2YXFC4PTGy9DK6pjuCyVSijNO8COc1UsvumuaBuBy56zCl
kCvJfbOrsbEiuzWR/4waNCAvCD272dSw4roffW8aFxYkkDF6x2MYsJQPe19WVUu4
aoA2yb1Y4mHHyHJpn1/Oex1QD3Yz1Ucp2I9q31Carc8YAbG6QnflVh/WHNVsj/id
LXI6Jh+00ptG+JCyHyS2GdD9uFGtxPzGG+mpe5NO40pUroj9vkPgUW61DzQRD8B0
cWwhDgBSAg0pjFOkjU5CAmnQWUbY+QZQ8qELyCGZdSOE6ovM06DZj+8Jjkfxm0vE
yrEMDNBpaVU/sAJOriTMxREsaPkyrcC/J6QovX/LO3geNatkiG7r/dFWBZwmQeCx
B2cBOO16h+V5HvkIIKB0HTx7sVjc5rYjL6cHkQdbiJYpaZEzAY6aitMFDR5Djhmj
caOx75xK4DZplNHVYLqGpEUF8GiDI0xAoZF+38IvEPiF1/QhAD4zfTkFUmtVqjGx
9ykE1IYW7WuaXJJ7tOmoyhzhebhZqYAXeLC3hnIaNCC3KxHF+jtGueYK9bQ1ubyv
FDoNy8D0ZGAksAWslG7vLFXJE74oTUr1TINXl91SXHJ+ADcPG1TQ+OSmVVmx9Xco
AAbKgfYOp1FI5H7cCnXE3Cn1w0pIODuYPMe5T9FsdP0mZCn0tepIRr0CeMt/rzZb
vVcnlEO3L3j+PnpY6unBMiymS70AOypPMVr2ByNYwZP0tQaEUMTgKBmAgriZZvSr
lSHH+O9Eh75JsqyYzda9FaY7OfD7RVj1/YOodrGdREZUgesKbqRnKCj8OBWq1ys/
X5yfAbyvoA5/JMQ+QIwAjqxuBS1OxA9g9oG+fMVo3YmxpryXVq8fL09l5Ox74dm2
clphIlT7a87kd1D2vdP4iLiqyJJvbEzTzN3bw8uqYSjzQI0dkSXyUSiNyWGoHwzT
RXRn5ygXgDmdTQtMOJ2IKn575e8k6sR4nCBGUDLoT4BlrsBaLivylP7RXIkGO7Ti
TA6tfQULSOrsVz7Hjz8y+/9V9xFgHSUlt3J/8C7tJLYVWM5rb3wHbByY2BkdGhCQ
Sril8f/m/YChDUUjZS7Wne9FwTlHm2UUahl6hpkbSIhwBWeF0psHudMbDeDVVHYc
XRNinjEt3UmyG+DnqXWB8YbOTPb0yKYMP1wlaCQWbm+WrdJA8h6dm42QhoXxyn5U
dF3Vtevq/HL3Pl7LfOaDeFD4FUJv1/AqcyQ72+hqPBj47+OIoWwvIpLYi8227Q1p
/0or1TXCnBPMXhIuN8Dj8z2U8BGaC9PYrsrRiF6TolA7jpsDP12oi+8JyorUoA/a
3cik0oge3NorvHnnOWoEvYB3icV7ID5aSgqXEgQddsKrnh1YxsWuYTeYyvjnksMH
oU6pPLN57YHh9onJ3cwD8MMCFfrV6Zy1CK1Ib8whWA0HTydwyVg2ejoCJj82wPZQ
pz4Emlwzf4ZuwlkSdW4knCzzLWOP0HaAcK8Stl3/IrB5EE2wEokQMouQLJR2mSiX
o3QtUAXybcSNU4ugam/8vePLzQsjt5r+EkWLCbBsBkKC/KGp0akz8/27l4xSe+EG
qBMKAul7eNmCFbTj0HS2DrR1azHWhLJNPKktdMNoWbleHi4/naHCBM1G81Gh8wew
k8Oz7tsmmizw1jXBZyYnyeHSl4MxvgiNPQgIOfhiNoLhzEqOPXr3+G7juCQ0BlaN
7aoQLqcdXKXilU8CQ2s9Erh8BhoslJRHwlj/qw3J/JvdRHnLvLOlq7LQSRM1vlqi
bGr/tWHimvCfiRrppKpm9zItYFggI/LzY2yt3wqRSNv62Jjm5pvehIvHZfZ8Q2I9
T58/uK+hwV+Fk1TEJEohgWD5nAaG/HeLd47yCBD/T6tB/Q90u/NgqkJG4tQ02FAN
GFXBGUq2SAp+KxnAWGhGzpcJOXe+nOzG9m/t/XUonaSAhxGeIj+6F7JAMNS+Jd0C
OLHKDnAZs227uDc1xt0FV6RTiZy59AtWiOqOyDGwi4OPt+6Svjnq4cjXzc9YCY/J
Wcs9dSZVDEhjCzZ9A1+hOFY/B7bjlUIMwrGOZDCLI6fND4v6IMMAFPxPNkKL4XCb
7HS3QE2MQq/6cKfRvd/fnQ==
`protect END_PROTECTED
