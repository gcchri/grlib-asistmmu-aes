`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
By9KfhTsTYROsUmgfkFzFoan9mYFJzNwOFcfPMIBmKRVp5cF2FohyGqHuAAJVzdF
B+5UdQj4LX0udo58oZjKVMj1h3/rkJ46hI88Wah5tWfqyvk8iw3eff0fw5Ae/JI+
ncA6PxHcI9oYgT1o5PZeQsKweIpKTjVYfmLJAxba1hudo4RebYqusqk4CsBQvCZ/
WrZKkbGzSlAEs71mLSsBAHmc6bWZJlDQ1iHUAthoG+mVA9u1UGukMP2LGREP7JjX
asHCH+hp2z8t1MBoyjSwQvZdpmHguzO5Mn1+hIvxdTJYSxSZiSh1KgkU6RyKZsjf
RdMSDHBHRYYx+5CKGC1qrFQWs4dIpzJ3RC34t1S99Zs5e3+u1E0R8ce2w+uB7vhN
c3TEAAc4YDQ35eMuKrLEffJApJiQdAvs5Wm+OqrcPVI5ulRo1mp7KqOUid8xks3J
QuqVAqpOcwTsNha0N4yTZyhteOrKCnPucFuTwA4Kpj2rLyOlNB6i78FjooLy937d
dJjZtOiikPTisrGMiH+XSx2806rHHlCiBvuLbxCWV5JBjQikbLHz9HerMh9vW8ie
Rfs2PPr3GYLPnH/P5OwIULcDvF/pbV2HVKZpkggkWAhGst6JxzyiIVvXj7rIHvex
ho76JOr6R1obtvW3o6PXBB6+PsioLiMYUXKO7qI0j0kmM66RTp0Tw9f2U5Ot2hA0
//BjhxpbCDw3hpgSZ0npwZdfIiA9LT69TZzRWjNEynXnfwwvKusIRJ0D2gyhkZvo
YQBrVXAfzu3RODffAhaavsxxrO2d5YQBCt7s6zOWb/6OItaMqbsWsb4jH6vQJ88B
iw6fxomTZV840eYqhVhQ6iHFOKAxq+im01tUL1N1Pu9lYJEYkXnM8dYDp9yA5Qd+
bP9Y7tRobZnUhWyUjhfWEIaxWgRf8IYXU1vinzNqz8+0wxNRq21QvhoA/K/mEF4L
dlPyXLG2Ch68s7RhwdmrC97BWPx7Ws/aTaVSs/5+kDepju/MSFJWg+x3KVebGRHg
2RODutQLptkocMZ69p2pDHOJASbcXyyCRUlXlWAsgvmYwrBxItRSUofciZIM7VnC
Q4gPDdRajWmOlrfIDMxR0kC/G1PUKrQ4sse1+VLwdZOjzJk4NQ/HuPUR8mf3yBRU
E0s1E2BQ5AF8+9AYmlOqk4EYFdFG2/y6WXFab4KBfFS4FbI/YOqP7djnjm7opUx+
Sh4HnYSHZWjAWt97X9YaCEU6KKWs/Fwf+y+A0S/cGqhPidkme+Hn4NA5cgg7H/oG
BwfSrMEr1dnRsMa/fJLQTzedLKi11Jgyo0nLVR+JuO6Vwmto5hYGNMzrmcYG+aJ0
ymfA4zEdIMyR0YCs4iY2heMn23psHsux9bQdzA1WBqWMt+pS5qypug++Mw4z240r
9SCI8ImHkqn5jn68rkl/I37UmYNBmnIUMvh2Ug/vHNYBuZNE2a3GWamnBeYlK2Vo
SaoO+Sod1VzZ1ydyf7vpGaoVeLEm4rxTqUNu+/WTeB8r4XrMyp4W0zHyaP9AOt5S
TPc2MgbPukBh8haFmKhlKZxVMQC68sXxhaDvpYUt/jrCBOyERsCKuiCxEVE7AJYx
rVvPsjTf9Qk+NYqa3ot9qgTkgT+woxPF14yVowFb69psFGkKKDY2zUUfl8Ylof0X
tD+RQB2M//EYmE/CiEZlrhpSIISr+6Fr3GnKD7CobLa66bCC/EijQFbqamhIDyo+
qmHgwQN+OaEXBxNiQx1LvaALOBylKItFISpKe1GUpQl3dQXYFKpNcd3KyioUxN4S
6c69Kru7rTWO6fFP27kNRWeHyF3sRBNzayzgVCeRPpYFrsQarsi/Ag8esuJIcsqt
GC14MQSl22hmKD73zlgRFvA8wr1jtsuvtZ72mK8n5S1E0IgpYNxHDKTZ+49BK45H
iRrcZjHaG+EL/TJ3be8b6bBVNio7hz8zpKJOQ3FWrFJRvON1hxegoWWByttB7fyv
QvgWl59biLgY1KNa5rI1CjLxbUqSV13aVOrz+1dmQoMeTtBhglw/12b0pZZnCcCC
86L/8aG4bV3G/KWrXTi1hs8WqrG/9Ot1p2cxUg0cZ8hxcZlb/Di+b1a1h1UcxxTr
uoFaZNVOz7p7lY/E+DD/v1VbAeyvWUYrmgty06TsCjiBQ6gO64Dz+at6FcTymPb4
FqGp13Flsoz0pgwM/0ogVVMgRaudmIbXRPqNtChVRn3XFUihkMpNVWmdv8fqrskW
nYAA+L+3U7FhTUv9z6lSI8xlZjxcFJDeCVtiI3Fu7fxYSOn0eo4HjOtCxQaOXnQN
0tUq4cInt9eRhM1PDcqy8iyRnkxiG6wTVpRlK3pQlH/fYywCypAcvzmrrLxx7YmI
+NRnru6yHluHSgFrBs0X20Ayrp9KnwAwAzAzWHj8G7VXcpuattmZgJ7yNNxmxC1d
iQAdubWYVdDAqMRB9b4FSOVcIfmZsdMS36DxcZ3nOxSgwqYEpsHOu9JNyaILoDTV
skRJhyXoUBspjliSWK2EKQ7FwAMTY3RJmAkyh/FRUhlVF2MSS6WIPxSHyvQNEeSl
384vVeC2kCzphDnyd/a7iBH6kF7y80NRcg3ZsrDxh6iLqSlPjooSDukYOf9XOViV
Bz/46uP6/UUUyprxCR/18ow15irrKZDZbGuKWorC/jXJtErOJsBQhveDPc924me1
aJyJYbIU7BdUfM5VlKKnU914GsI8zzkoIdceFwOZWWfOrkFSskYJRsyGcN0BNVi5
uTzoivRI6UFTiZlMU0LhlXn002NURNOSv3xAscKT8dSSIwGiR561k+tgbAobZl46
fwf0ydDsGIc5zw/nto0Pxm3OY2hOf9WmrzVddugdL871+9k1C+8kozDpume+fSDq
EhRHyc9f0ZgXkPCu7xyqGcs9y5pVcI3dsOzDYaqjFpPdZUiH5YA8Q9rfuPqe98tp
qarXfaiWc8MugJY0LZH07w9UPcJ1i44P8kmvfoHQLR3GfmSM5ClAt14zLrppmvHI
vVOi53EOE/2WSn6mtmXGKItu2QRJFhoAucI6tJflh5hqLhYC7XYOPkcj1bFlrjLw
jKoCY23UowsVri25kALf3xHPg0d31sZa2gBZofdYz6zynI5eR3uMA1WcWsHb2FnP
IAE10t6gy6032DuLhUJ1ehGWlm4aBbBb7Jr57RnmrvGcCs7fwmyM4s8cV9hHsZVX
wHzpZCvo3Z/cBfd0DsTFjDUNQWgajqaHnOuL59aVqAvOhkbbVYhXhnIWF6gqNHmE
iS4yX04JBq03RNwShvazKgPBMrXGXaMS8ehp1TBuAHmgc6L3Z0NiCAaUHM6hxoNt
xyyeLuiXGmLSjrMKdWb2qVhQxqG58zEMyrf72uMwcARV7ruJk3ne2XmAu9QYjqYA
FppKo/FqBhHOe8xjddESZmgcHMCZ3ajXbUrWrQuyoHP4lY7LcCyMf8/YWBOZdoIq
sl80i3/sIi8pRWvilhHHFdIERK6UZt8IlYRLuXp35IdaMOFVrFCYAg8dlH+sZvAW
PjGECB7gA+wZKwhNpDy0rF19tEJPyC1XJuYVeeMCM8aZ0m8ccnQcBDz1MvUG4jqu
qw/Y90C8hLIb7OvAZGcd7wg/j75EMEPhJbipNsK75n6XOYJ6lRba7SxEo4A7ki29
2sUtUlepf4fgyAJiX6RNsYGBh1XZoVFKeK9c3qGeGoqchx3fw5EVNyXwHkM+0fgp
sVsWR+/Sbz+eRqSdCW+jJg7Y/nS8xbML61WN18XOW14nHP31Mfjn1QD/GAu9zaXT
/Da3VXYaKWCVI3nzjzSWUYpchA8eFpevs/p0N3z1bg73P6K3VhoQvf1fiQXSUh0y
/D/OV1S/RE9qeSDyViLUX0VAWAWAyjqzA4bvJ2scLSDDCULJw5+gbb3+i8cwQflN
i3c4UEVtJ7RbSiGpUx8uCYldoQY5k6NXHf9XfJrXzWVPrT2/CeY36UeWUPZAnD8L
QNg1oAN89+oPTq13FCOjAX5Qa5/PZkklCGMnQwK5IwYiI12NT1L8N8eEaFy9tJ5v
NpjRcfLqfOkytd7ne7ZfGjJXoZnU5XGVVuQp+gXxfqdteUhgdeXSEGv2etQQWTXI
CTXiNdIenpL7UEnujC/Sssg9lrdT3iymrkkttJUO3TEMljd7YwzXCYfV0/w3Gi/c
H9ooTocxCuLzfwkL4wqTkKLB3eCzlTAKxg9bHy1eahjCYiKdzf5HtmBn/Pig2YsT
kcAzLHX7k14ihqF2NkZmF69HGxrUV7eZ5Ij5Uq/3Nlz3vobMiwggmv5+KUyvcVvU
AIfmnmTTBXIxWogkcobMjWf14S8HD7y+W4aNOszQuCFAgRAAu6YkZ7LlW5NX3yGF
1ehLbWU5W/SkOG5HNoEEnGXuuSMoRvdzHxKXmZ50owETfuoV1bX1l2jrMYYkyWUK
iUeXBdfw2ZSFPNY+mu9oAxC7NyYE3S1B84AuJs+1wx+dmO+SX3jNlk6qy2THbMAZ
DBKsEt1E1DdL9bl/mqFaz+Zdl1pFiqxLiwG4bna+8aBDzlb6YnLp36e6GrNXW6o3
`protect END_PROTECTED
