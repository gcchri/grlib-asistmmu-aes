`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zsZDKFmgEkHGdlzwZWrCEQ/AQKL0y9C5N4CLpMPosF9wuWh8O+LaY1zrp9sQAmI1
CXtPy+yPT2oY7GK6cZH1Xk31+2u9Tf7q4glt/yniMThXfBNLm+z0RzMkeaIZ74eL
IkSiLqMGJEsrwRzoqY0OJ+Em+yaMW/ppuWfdP8kwwWbcqLmvxJz+EecNeaSc04l+
lL1o4FAPQQvoSWnqpalXFhRjmoy/8T63iuyvjsMJzsGJuZtWuYyNW/cWQ5124iEP
HLcuIAZW2eL8a1Luu+0zYnb9LZQfODy3jiu0jjMFAnAK+pny394r2yDlDSki7nss
tci3KztQzzwKXLtVqJ6VjQYNRkUL5cyMJkpHsPyaZmEJrb8n+8B2SFDB6KZRbdQC
N0KpDfWpI6jKTqaKSaCcbYA8WTqIWYm81poHdPVrEOzW5YYw+GZuvUuo3/1ePNKJ
J0II3SwsaOzK69EiCPZaYg2Pu7OU/4jMflS0kSlimzVisrmybeFWZ3SCgED6HRU9
Ysc3kY2Qe92Ep5sQxBUkdHP/B1aYc98N6RrZhk075WdtB9XJH3QAoKL9jQMA8i23
moLlwHJpinpzxCIW5hTFhfIbVUqMVWjn3PVEdzo+yG2ff3KNAYwquOJ/sAhXQNAf
VJ6sMfZyWw6+CbZgkfVXI5WlUjmpBY6FN0Cw0WB8IAiuOxkJ+cVLS2bjLs5dBEZb
kDIvy9t2jbsJXE6pzs0ZGSGxoc3T3xQg0+MEt7+29P6R+iV5RNYj0uqPzSDAdt6K
EpVQN5BliUyEIldFBpXvEM+L9Ezxy7xqWL1s6y1ehu7TOUvnbGhC6OETGGVkXZeq
0d3vCwzqYFHpOZnsl+v07t16x3naq1QdlobOrmFqnI1q9cyCXqL/sVKYRl6TnMRw
gwL6/4ZQeRlWOzwJ4jILALWjNKdhqZGlPtg4FzzKkqD5O8eYk6Tu2ioHNAzbr0ru
90BXFKVaU3jKtuUJVkgff6q4kYqXdlk3r/vIRubRke3FJJigEJ4gQxsVbX7HOVri
NnNI5oissEglINY2YjwZoWDHPLlEuXnk0dBY1GndTl+Tx/+K4J95cMiKvc15XGui
IJIoFKyGodDCY8exBXOQeg==
`protect END_PROTECTED
