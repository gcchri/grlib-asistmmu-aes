`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kL11dJVrZrVHwRnZEbu4Va3VYQqQU/jcWi/+K88LVMZ95/VF68GOTScz41+XcADY
wd2fLzZimLl6izHLYK7jZGUiGURgeod60BHlIuTIAeMFomYarU9wsLCVJr7uCI/m
QalQRXp8V5ahn+CVykbSVzrI+JVs25M10CD8oYLsR9U5dR4bT63P0aYrQwFJs7hE
rULl5dxUDxgIZIj5VWxgnIdSWFzm9slXvycFslrVPksDNmMbpUDdUqHhdn737P89
o7aUHq0l0Ti5wdnBG1q0gGTlEVZoA60u0wKozvXmA3PVFumlQQUVzEw5tfkuFM/j
Hr6iEBP+p6ts6O9ZdDckiQ==
`protect END_PROTECTED
