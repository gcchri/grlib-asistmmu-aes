`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OJb9MkjYlzQk986O0YCYe9lA91BX8nWdVshc5/pgNJutyxyyZHvxgxqppIQM4+ug
6kcy+q3i+0ZtiwHEI0oUxQhmHP/clAH7w/M8kPa0qaMnQ/oy0UanXXoBsGnHf587
LlZayJ8KUpC5I/tD7Ds90K+O1A+/vHoHXRCJwZ1pAJVMdk/ne/MpD+JTHLPJMa/a
buFTzNYtzTlCyn0sa3Q85XlDy59mVujAH63pQnKKttjJim568RTOcFpsDRYsgY0M
R8TP0tYQgWARNEtQcABW40GOZ+9XixdKLIzOSBAeb2o=
`protect END_PROTECTED
