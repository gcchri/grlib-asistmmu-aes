`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BGhFN7upPi9zbvzhWP7v3hgfehAUfmeZ8wO6A85TmSkhwJbao8gTAxusS7osqgkX
v/HwBdNWLWkPLDHnID+5uQ6T+HLd1MJxsWUQD/ajUWyCB8h6sy/cQW3x9NjCgySu
IpI5My7qZbvhSlPHGvzIq29ZFu0MFpJ95sXu3du03h5zixRqwXoXeHPFm1nse0BA
UfM28Zm2ILu3MYcU0bNSgC2z438mlAGBIjn3WDQdu2jVDu/GD73GUgzJ89TgXRsC
rObhMCdiGsr0RTDh/f6dHpMCC9FPs+iaSDbRhKT8LbThyyTzbHYA0S7emaGS0lcg
4NqmsujmbbrjkU9C/kWCJv2hphbZV+Qvc/6JZJybJWoZ07YOPAo18zarcU66hiq8
RkMAKb+q/clcwHjvIURsG1X3AO1VYMYgWAK2zXeKZDoiL1uvJHqOX4OycfjBUIDu
3ssRULnmwvN2W/oNsztz39kB3BMkM6mn5+v2oe5CmoGIYyj4R9tlH0v4krIuihGn
r83jOTqWUXjOmJTC5UeUxwOQxxMYHTiX9yq+SNx3hR3iLlwZku03dcF8pUmcN/hA
1kYrZT9PMdEa86YtnPpvmDRQoCMA5WVAqoIX8dlk/fu+EshinJfU2o5WOAyJj1Qy
BMhJG724XR2mEaKY4w8CxR7jtdLv1Qx+6hcOJedil6pHf+aHMjewESOaKaPdluX1
wAxB341pESXvyhBBhuFpXvKb27aE6a209eDjuOiRd1H8McS4wpX6xz483/TRV+D5
Tt9/Xiq8p4VP9lY+HWtbzexZUnUOHa8T06MgarLvpSZ7JaD2sosABBh3mPJMHNbO
ZliH4P+7Xsj8Ax8l3LLcyAT9+o2LeaxbU5mYL/pHkn5y/GEkMS5UnYrunZV/nqQd
Pis2C83BC33aQZRfXBT8+xwXVI4RjjgkFjWkybz7MmvaTWyenMSbR0UVJ/Uw+DE0
raYV3KWWMP0603fvkN2M8SanVX6qztL8L6Ye58I6RbS1FFfgWnKNpT0zMxSfCrBi
pcDQaP5Hj7ztUrJwvwEr0ZQpK358aiD3tLhxZsB2+8mcc7QUfYUlNxp6Zpd7gs4C
FZ30k7Td6cTsGmpKk7g9wBoYGCX3v7yjg3tNHCJ1dH+3IVUPvfN9kTQMJRGKVi3y
AFaGGtB/IU7LStWyUxrN2Mc6ETXTAneDa5xp5ywSBp55awLdm5ET5tlmB92GQywq
i4PxXbvq/Xbr61Y68B/Az71SIGNmpAANFjvg513WpJ4UNsvO2vNqiuAfznSOMOAm
Bt9yNsMl4Q3jkBlSZa9E1XNWnkOuK0dGgKB335FfbtmYUFr0LRCQALPOpyw1wL++
3cnFC7TPEOMZppoQF67WOyZ9J5WXvQ5UHU8qBs5HWabvRvijILp4l5p98c6a1+xz
2yGjUudt0oshhE820Cc+g1QpU/+7PH0CZf0Vlq6LJUhbqGqNp/MIF22BzdTDFlaF
6ecIm04lAPc7n97K3R0+lWPdsZjoCfvwv4bfiH+/wW5PQVcWJDOa+bAc+RZt35FG
MeFQ0kc+2OysLT70v2n6v5SrUUKcISbaNgBVBo0Se+swAy47bm8mKV5nKLkfVek4
hfyhKG0j5ugfoMmpl8b3AXRYExufa8jpIF0oX/GnYkSDrORoe7mZcfAC32TGzvgL
SDjXTG7Ss/inHww2ct9fRARd80AjWiA++Lmp1XZBkpE801Ur3pGbkBpinlI0Juwc
w2vqGM5ylFL1gp8a1G7P2bTZGi2r3/EngsshxeS59In1aG/lj5e8SUCpJFQtLN3+
7ttmZetf54eHXQX8Qhxcyg8UHYYM1RFNeteloQX+W1YeKSHRnERAqssmOaKlayhH
P+VS8sXz32cukuxaFLBnDhAPdYoG5Zjv6fehL3b9YyGLGt2sYcNn0EU+DfRejQTC
+pwWF8M5LqXHzgaeiHqTxMCVSXz7StW6jdkpwkfot2oAoP596CqPsq2//g7oErnz
42Ogh0rxVxxPgOSCO6NTkNb4+HqvGaWJBwLzvZ9bShL6H/sixQqqZBxRVUJIQJqE
3q92kB4/ZmZyCPok3utnDUiHcZ2iCwca5DEBmoqIqBSFPexUaTzzVMLFNtGbGyFZ
JGbZZn7UrHYHpoGrqMlP0xUSq8EcBDGvZ0cQWX5Qi6t6MpO8/ezikYx420IF1Mrk
hFsoC/PNfAFbLMYXH/dEWAuGXIOXdMmJLvOAGdCojzSKGLa+jzcPqRTizBD2oYBX
gtqQqnq0uqNQAUCFN9xt62pIrktugRMGF0AiDrtCuVOVkf3ZuMJvGU50+/4lZnUv
TzLxvpvT021XA8wZjChGU+5sC9RszMdTr19zlsLLIjX69mcaZ4XV6PBFaaW1Qfl0
QrG6w5ZWhfO6bchKjfgisRUvCIasc85tyyD2dc1u+H35mrE6rwtxz3f7nbzNX8TF
BUH7ZHQ/GdVtJAgNt23Muo3XtH/HG3d3c1AvjKJUMg4O/8YZbwrOhpIWdpoVtY0h
pRBSBm5YjlQmQI9zcyyDK2Xdm+H/jBD74zwM7Y6eWf+j8e32v2oI8pfKoHYJMYqU
wK/n29jYgCuXdRsW9GKep1n0lvCxTRl6mYoCUEW2Qw0DbUVCxtvpEAx5aOkirxgl
/Mvb6XHebDUrNuNTSMdCzC/OlzSbvTpd9s8lfatO2RG3c4CWIUtaylFyulgHaKGf
bKHvcKZMxu8P38cWe2YR8P390mw2wMywVdzqB+twxdKPT5pagen8DvnzUXTVXqIT
Ygv813PRvKeEaE7x+KFIMHI5B/+z8WKiwATLW2uul+mlZhclMGjPBv78IFJbQ0YF
/oRwkoOAA9JGyVOuZZndsRb2EBfe6gBVdLPBXx8yJ2Lj9FgeYvcdH+mM0VZ1e/r7
NZ6cDEstul6O3xMz9GP8cG1O0vgvy6/MLqGqqKERJayYkEsgF+Jcwz9nmLvpX6M9
03/a3ZpVNPbZSfsX8KC0yNiWxmHpLbGqnBdx2D6zKh82XsoJZ0DDEN3DQRKo7s9U
2ZK9TuH7qAcV/AU0xpzLXtS016U1+7BmPug8stwj41pAYNiNA8nXh46+WWlgOUZz
WZnB8HFDaRssOaz8wN2LtpY7N1GhQpbX5ypKpmzCJmtizmRk07MeVT9JopQ3aqBc
2UeT2199CVje4/WbtdM6bfZxei5IZ6kLICssAq4eaDHr+jJzP5tPI+FM//fCNXlF
2Yscxc0PUA3rkXP0esS+2fyO+A2qiKCmgvznLr7agF4RqfYkCXOEB4RFwmmFXdvR
/AG24zXf5iVukY64kop1+ZOskmBptR4SSWuUcAVh4m2ZT8REeLjVr29sm3LXLFp1
oywtfR3JHQvPRgpem3sYPUbHAc+RgBh6atS3rfsOLSLCc5lbKFWO0MnKmpf8bkEo
dAOGrYKBmjxVJ3kSAMiLQ0XnVCyPuzoHJyWQ3o3GTNBFefXg5z31TtM3rUH9xvVz
uG70v/IWQ997g4f2i9joBLXkZCR+MDP7qu5KO6YXRRjTmNbjPhkLVrbE+Acjev8j
U22VaSj54cJjbNoa7uOLG0m6avcF+H312N0jfNO1muSf5kx3tCfSwoYsXp/zojx2
VH5/zLMB1gGmdaTo7yNlyW6btMzWYTiCrXABvGd4RpjxekiCV6t3jlotM6Jwsdg5
dmKQldvyvasKj0LiTgxvpRSyOmDHP+/43n0wyYjlt59Ryowei41wREBIn9RXkGUH
hPPCKFFvO+jAOGDMy6lnXgBOjIScsXOSUV76rCcYkJRsBkOKW84uyqSHn0I/UERM
OkVc+WesdkE+AZ5WLTeLLa0/Be9GeoBhtVHK+GY9jSI+82xeLrPhtxWFnHZwRzgI
a4KMFhQ5EXxRSQrJICMvSA==
`protect END_PROTECTED
