`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
apiAkm/u94Bu1ZvWt5mgd7ujHovwxV9fAInRxM1L85wH6zfty68Y5TT8MMUwKADl
2durWGi2JUNAC+VRT9iyqboEqO5bWAvGy2kD+ia54XtGrdc02DUAhJbBhzzhBahN
I1uhbd5y2/ARtFVJsFpsJ9L62fUKPnKZSIO+altFf9OKOcQQ4sBlyqcK3L92H5RA
wIHQYJRJEyerxtyP0KgXdIruOhRqI7wixhVqudyiIJJZmmyX6b3V2dEFtpIrJq04
65gumji9PwUOizbaqMbDkSXNsBgjPQHGa97RXh4BVsw7nECsj+G7MkRnyzTHxy5S
am7kEG00jdA9DnEL1xMfelV7LpnILFLs6yud1WxSI+yQcyNydHOZWg0V0yOoqhpa
2yQiy/Dt/HR37S81U128nVDY7jc09UKRfTuOGXfs9I3RsQehTxQ13USd6NL3VFXS
DgxBNA3+U9S3/OIHGUq62FV0pWQq5ubeCNGxNKWrbTKi+uAlS52A0YbMTLEXkGAn
dJm0B1sVG3orNkdsHvh9kogktBdsY5Buu9OSJgNTMfpMTNzaVTPjwjwj951CgFCm
99foQno00qpiRa2BgaSxKW4ieWzOc97GtUN5XwrhV0TMDmO0jAijLyNWC2VrrS+U
BORVX6umUelQnrMIaalkY4E0FWdZ2XK2dJl8EZ5/lCdBcU9icd3dRTO61wipCxjN
ORJB4Ks9rMQbfoUVlA2YBhWBLzP9VqkNJF4Mnj5FrKrfBpKh48i1DbPsC201xB8q
8mnlzA/lhkhtE5Vz1Ryw55HH+lZjohshSk9tKU5ljavCMCAjagzAGR2q8AghojnQ
alCdZFodA/BBLkcwkCpgCttUNZ09zhcqtShs29wvf+nt/rHZemK/bfRtYhf6npmA
`protect END_PROTECTED
