`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ob3ZSFHH9GjjeamtQ2PvVODoqygihiXo4MCYOnmRmRRnPbdozVs4txhaB3YMH2IQ
lRMf+XWYFA232mqAATM3JpECTwTagd867Vy4SmdhZHXpjVQZFXb7AdxpoRpyw39/
jth5XoeZ3NbcgBtcD/fbWGauVBeItsISbQ+L8k5DuT6uaYW4DBNc2vDh50bmOZIq
6lei0khJh88Gu9Q6NcFfbeRU8CJFSdG8q0djg1t3VwtPK0+aTZvtB+IT2rzIy7Cs
3mDNJJRdPYFmfpjyFA/8byBSzXJmqKZnh+v0bIlQZA1KgUqaIF7k1ybWPTlszn/N
F+/nFOcY2W+31gfJfBWXKLaQm3SjvLklxLojK0DQ7ACUI9KrwJGeR1cAq+6HrkDL
PtuFhIbWAfUWGGbZw1ml9A3IYYNpAFAH5WjFY5nrsIUjjvfugJ8WoYRIEJlNwvjf
zUYnSPS1CufRi3cQILgwi8WbvasXzZh3RLMDi6tYIYum8qfTlSudo7t6YF6RXxtO
BVZLNibVk5p5FqrYpcXEQDsuvdMt6faePSObdG+J2TVXWj4Fn5C7cJLyBQRqzmwa
qgf176Bem/zLbpyU0lIy09MQng2c8VkYJQLRbOrFTptvIeULa0kzLBrlhpe/IdK2
ukq4hkvuwSbPjt27KcCX0R/tKTCIbHeJ4UJ6YH+6bYZ+T4xajsuIdqGXYMlE2mXJ
vtYPOXDBX+PcHC/DmRM+jJDtYyTkgmagkweoULFseXpSN0pr2hN1Y2CPuxqvbSCo
/DmgvW+SnMJIRqZjAM01NbQjjUvaegiQyk6UZQPXEAKET7UfcUvwTYjvHc51SOY8
+iflsYkj1zpu01Gv848YNjvAOvvM93YJWqd+BlSbWC+hzDeUYa8G/m9aPRM+3NV+
tZ2HnjZtaiyhN7A3OW2tVXutx/rFjeAjwz2o0x7MbWWt8DAOTZ92FP2oVmHHBvsn
7Hu/8dkPSGN/FpGljTnRYYjV227MslurPzS0pIPWK95lXUYuLPxMo9zoQr7SnnRl
/AZFxgPgpHK6tVu9nMx4DhcSfWDAT2UD5TFYjEyw5DU+kO8CD/PlxHcDFQWkC/37
HfrxD6VBSAyQR1eYI8gkU7bDfr2CPrTePbp4cwNMNbxBf54t4j2HvTkxEqVC0KrP
p45kowEBH4+7VzXFj3d3Tb6shOztCDOmlI/pHBCJzRcK7eScq+jlHNzGss7QV27u
Sd2PfvahDj93hwhDpWJMIIsFiIzNMZVkDq5ruYaFBk+pN9VDDTGHXSkKRwdExxtT
d7w2jnwxkXyj7xi+m7zQcjkMRHd7OKfqVPc3Nv3X1bSCbgPeS3cPWXXd1Ks5WWoQ
5SeTmB2t/YhnZnI6FrK0nHDhw6hDnE4nuJQrKxO2z+8Ce/zx7AYBgjkRmQdgrDjU
KsrDu0KqueGJKLjmWPD8ore2Vc46nmb4h7MK4eitCj2+blcZGcg8I9uy3RTQDB8Q
MTuipvGCYSNgFwEN/M9tPzjnfYxvk2DXl0Ctg6aVuIz+2jFnC1TlE6M8e+HoY7Vm
yGISamASHHksSqEbphKuLX0nW7pOX79edDMSWBD8KB9mUONECQmjMNH1jTNXovbG
BHi3lzG/WLRjOnD5IMZMIUNtnLd/wXGNCpM1adrCK5ikskGVe3mXLOiNA4UETF6v
veNBAXlc301ADAuuzPh0Cy7tD/gPIZmfLMSAko5bjqxwFoGkYkbfudC/sfaIvQvI
69PK/E7F/yAW0RszRi4I9DvY1Vi4jLmvYtg5nmmxN7klBUtHujQTuE7gsgxepYnq
6KCiqYrwf5UgpdIbnxUVRdPIxCwZSoBAbbkrCl8Pl4RihyBqM0AZCfIDIGAzbjni
nz/Nfmcqr4d1feZrvbUEx9M68au6C1yOn2EavvOaTv7fwEZWiTFIktR+gso0Iv0g
ndBv2A3TqisAqV5fk7R9sG1n9Rexh54GR6Q2tkMFPqwjiUy5yViJfluQCjVeK77Q
99ZaqVeibPTTv+BIsTYqFsmhR63/KJJM2iV/9f8FLteGeGTMRMOPZc6HhwosR40q
VRDb2vH/8hPExWQ9EA4oV2kjm9oRJc+vDJoPu+WOcTndfamv6hAzKe8FtO22I4s8
mSQ7VQJ1/oq1yvFsh5itmZF0Spknnzu9g/NcrRQ9d9U=
`protect END_PROTECTED
