`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UUlUfr5EiFF52t+V4axgdTISlg4e6rDaN7hHmMYJYHzhVjaKojJWD7HpTamOC9Bc
pzEW4LTorpnakkVVzro9R/bGlKf/jUb4SMotCHd6eDabQdTvpqdYBtgOt8Xm0vOW
PgPoxC/ZrjgxUngyPisBxXQSSNGM+BAwelOQhYczJHJ7JYxHk4fMZwUhjDkS6dAj
6sY11/T/1HWxWqoJ7f47N4lHnhhoI4jr4g0bH2FMtXQqazC3k71Eix1CpuAuvtrU
xilhFg5ik1lpvRv6F/5iSYlaVDQxIoBayUzqCqsYyjnbeoCXER1icoUlElEIzgdg
z+61zPtwLf5ed2wOR9wBh63kkjhT9K3aM3eCXcpBbFEg2nE88SPwKqMExMhRN8ZY
4OQ5lESPhi29E7YmhTKAKg==
`protect END_PROTECTED
