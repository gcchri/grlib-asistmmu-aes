`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8L8FOyPc1FEWmu5jJ/VkyGPts/SbA+blbzugMVMfroaU/C9L9oZzX9NYd3TUB3Es
/NGFZXXahKIP91MvEgirHgVwonvGn3KGX4et4qmO9z2ab6iLUHiEm5B+vzU8g/Xa
bHptHJKgjk0dQOFJozYexht9ZU5YcSieHX2xMs6ZS0hxnbfx4g/5P7FOBSVdsvOx
9qWF8Ji6wx9q3II/ku9jGo+wNyqmDNEctEvwmRpQ34YidfBHIl644XIIMSfJ0rVD
stmO+qGmRqRl9TJmT4T6gDQV6TxJMoj1SZfAhPccsbK2/Hh3GDYN8v79BA8bxJgx
7+5oyMKbmEM+THvDaFaI29ULBvBYU6WZKZROhSdIr0tFew/r14JsPQBx6exAgBM8
EE8hhAon111xEL7iB4Aaxg==
`protect END_PROTECTED
