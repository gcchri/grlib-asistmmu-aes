`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yy10F5PIsF4YX3MWVpS8/pnDFVlWoP9E/mSxXekM88mC5UbH+chTmMlBM7y17WVu
u3vo0qJLPGSntf45nxycmxm8a3uPQKucBBEhpOS/xo32YCAFU8j/IPDtMCncq0Mj
qO7QdUBtT9kOSn+0Lxzoo80aFGjPljBpl3pH8VwwRTcFA93jaktx5y6Hnz96MNNh
jCVsppjEjM8IkXd8+sOJvBXxq89tQHxn3SAXEql5bOSh3at8w4UyUtjJ6b1RO4RV
NU1tnI5rwMvKR1Mkm60Z8NT9J24op4A1RZ59YQKpaSTzKk/QHY2A5mTYAIx7300s
/0rja1XT8pFiiBnMjNxw1r0ba5n/7H3hh36fRgm6Or9+PcDtc2QN+8yUnfyVDExw
AY6pYG5HCIEoLF6BFyw4PvmsOah+H0myK1MaxqsoimBeZ10fvuud0E3g4ArAoLMg
tYBJArFFf9/49X8l5VY7thIVvtaLTq1uscbFC30z7btyFhGYWUlLNzV1283jCKAM
mM9qg7ICTDpTHM+dKQ8wLfYEv2TgXNNg2IQUUVG5Wvz2uAZIQHE3qQRzHQRAsLAN
IoyKHS1anqJHko9VqVxMJdxLlNMCUj0WdJDccahr6poIuTeAB7/CG1eN6KJnGbYX
q3sxEH139yohXbNm2tSzpS9GTB8LSXXSTB9JXoX2S1PAg0FR4UaGmAELfb8YvmVv
m59ltvVy94ypuCj7H0yBsHWFIJxtRh+U+vMyUbXiCwu+5WTLv7z8i/QyEVQPR33o
wCkOgYJ0EgXp2y0Uq4Qz4uSJHx36ZFi+fh6qxEkhn/UDTezMEyx1BvWeVzrEuEl/
OYTlXUDoCbekJwqI4VzDXDbcYnwkt8/i4AWdDQQbpjqIEDBLkG1zX4Bxw/o83X+h
zvwf12HPDyoYB7o54TDgEt8KV1ZCbmCGEOca+SDog3CEZlV5YKotbkEBhTslTr3B
3dB9GUrsQkWjqSnykgz/MYzlH+m3eb73okzN61GRYwmL4alsZ6Pw86/LcWGYxVk/
R81iE8cPADWJzIn61s2m7yjsXnmXOUCqJExrJ6NnhZpBLvFqlwgRaw0Z1rxi8lhD
28NF0QRcwV+eysgd1Cg0htoiaBsMnxpk1PtuJSF6Q0H+VpJOllN0cHeu7GiuWaTc
6WMxvlvytrBRpOojv/Yf3GuaV/J47zLRHd45ZH1GSMx1bYExmC3DgmETJN3wBjIs
O0X7TMYEok1BmwVDKbGPJL0wiWIPAQwEUAJDbBRRSYooEC1VSBwWQ1tNzy2OQlaq
bwWzgxQ0QIgfuVNaQEkJ4ChzlepGsFzAMmlaUZiVwRsazLteizqRHAQ5pe4fFkq5
41oJnFenv+FpiSGt8mQmONxtBzm9DRji1Tn9s4zXeBlLiC9CRamZKT/0YI2XCOmM
Z6rO5BKzuPoQyEDvM/vNz3tBwkoh5Nhf65JpKzPhZQ0avFb1w62NVlP5si7Rn/lV
30KEry0TnkqRlNPWrSJ4Oy2PJkOMfzKJnCwS1RHVznWh23SulodeApDSXJiXCV3K
54/IebHRheOOlXmG+a7zTHw0B/HDnE4Sx4D9xEpMFjUMvGp8gxOSBlk3EzinBIRr
+L12i/T0L9VEsHa5N+Lf+nTndjMpOvP/HcOJuHGZvTfZpMRhy0Mm4PWJvec6n7vY
SX/DBDwT8Xtc6j8/0hiWRb2rMN5BBgkzefvVXxCKltvotXiJ1Q12DT4j8UtlHW7w
Natixj6Tn8L66HXZ5+6ZdZ3oyzbYwkgHfbB5S8q7C+kZy3MmyJ9YaR1dCx6d2vau
rI2Cm58I97/Noitp3SHAFQ5WkvzzEhJbnteGL8A8hDpbhzJIQg1stO3tsxlEIZxC
vFg6y91M7HeOGogfdS6kl1ql/bGM4zay4F4IUXqTLi8Y+6FgBTFfD/Y1G+9LT/z7
cEkTaloopqTVhAvIoEShM3jWxbJJqKn2L2vrQgqigKMFkJhWsZ2/G1nK0DYkruwP
lRztX52P3R10ml19pIkIYrHAA2E/8RvnvNhmGdW+iHPel41jl153pOq71cKofMsp
fRqXGiYQdDRFd1LojSYBU3YSpRjctNAG6ppBFfWIlaGSR2jxwHvLHvXflede4FZ2
TAUnXLEmWa4zcKhVJ/0r3Ucnmg3Izs6tt9reuUSnp9mYyhgRUOlVUTQpzo3Kny/S
jLSBUGfMt9Hm+Nj12oGrEfi4ApvPtz3HNKMUlWbaTHfEfUGcZXsLfn50+H6Flceb
IsccZR4lFTIm+qylgOaPvbFDwqQI9bpf+Nl9D9cdBSvINyPs2f9fYu/LxBQihH06
xGA6iMmHwUxG2p74lByRhcCXfEgnQvVpsXygHbxQPEkA7qfstpw3imTjPjaydsXn
F+T3t4+PawIn2LzVRKf+BDip84WaX/p62HOktvqRYVqkj+LAVvj0nGUjuQPlsU3Z
/r1xFkgn47L6/CKnaK8T7Wvx8sMvlxj49Gv7rea5hMen5AUAF1JxEni9mYQ4tgDD
FG49yQ3SM4D1a0too9Ufwy5esxa3AK7nVCUGP0m4XqSiilSx3FgEmdrvyFhSgCYJ
huqAT0+5m0GNefUvj2Bc6NBEoQo3Msongfhbe4rNBwAuEvoidS+6NI0H3DCV+Llx
8IO1SB72tIdFA2HYRXMkj13BB1qb7ghLdu+npnypoTbW/obIoC1h0bKVE/R+mJS5
oCJ5xCUQn1h50vTF3hyT+RO8S620cg6dYsNXguUFjlEB4Gtu+E3s6nGJhbLpCDd5
qeA+ovX8QEEf5jn/7InqFLYQ3afZOtVR0SSRBpN5e+Aw2NA6z0MdasNF0nR96K8l
2nNCqGD3OTdFBqikC4SbMA/IqKXBXarC9NTtTtRDuA9sQFeR8jq1P1B28rLwEvdL
6kZW5ycpioiN8UumsVzYl40aOsW+JrVL3z6uuQNqaemzgw5O5IDKOlVkb+Z7pI5w
Q4HQ9kUZqP9q33swfIMpkPGog7r4SiksSVOfeYgOgN+o7Fhi1FBki3214sQMAiAy
spJxTZqS56Z0ya7R4HR9sKbRPESFEr1nzsAvEGlsLVo6OUfRWL/HgNruHaPdig9a
ENwPExHqooHQCayfDeJpu0zBd4hs+jr6z7SD+c+YTi6JjSFkAfQNaKg9P7n7mzzL
MpJpZOnQEuV/V0TI5TKbyRk/Gxvi94GkGd0w4eBG2/LBHZyJgORxcFHyzQVSrYJi
flfFYnR/5+002/WesqA0mjM3lJt+hh3J/iY6JfEO+92nlgyRYEUZTO6IDRpNs+yT
k7GljqwomdMzitqC4EyI8jTcMqP9ICVzKX49uzpi+DXnNonPOFqOQZw1rWcJFzUx
GdaOzle4YFYfp1juO9Wzx4if87nkBg/DfUJuiEs/cUflHMxYI+f/vNowyifa9kFB
96BY+EwsueuIuT1IsW9+/qE3XghOjurZO5QuxGR8en2vp0W8YVKg/YgQi5887qjD
Ai+lVkSCn6aOh+QhKkmuB3YjI9nGOyunqndViNIz0byzbLP9iA/5BVvpJbGzSTf5
Du5K3QefNj3GyT3DirqUGqXc6cfAaWb+yHtN/KepAiFfGdveg1rMgc1nQTXPUtu7
5hVE2y0o8xk+1gZ6acx676UBo0ouf97JVoi2IRxMymIrCQHAvpVj6C/CmfW2msFj
VdMQdCMniiubVtR02QVaOHv3o6JkFZZC/XODNJxewA74h7TvCkFr/3IVY2xY+Qvb
0tUFLdU3GOTaVj4d1g44bfeJaTR8RDEzNl2NIC3f3ukJsHS5w861hSaZbnM4fkyq
KsLnU60wHlQeJkCkXUrAsh6/0guYmd2waIgHJvOt0WVg92tsC9bZUnrZ7C+lkqNS
1N9UMMgUk6oMV7pP3uwVtaicGlYxImQChw4FsjqQc7Vuv4H/nPEnwxe9qLCl8z6I
JDoZ15pE3bs/N1+mrupfKkia/nDrbH8/thqDqJcnUxse7ypd1tQr8MuhlEk9yGad
oekvR+KgHnGQismrYs697vPggGtmqJEFmCCikh3fWMJbiIlJ6svxN17vH7LVkBzg
V2oVEiQtTp8np+uXckUpsR8ENNNuj5Oz4mi9S6A9kZ+S14dAxAZ41h2JAIapIGOy
x21Kaj2RWzAO2aXrCe8stPwVA5rqgV8RliDNsv/sLfV0t/Aeht/ifl8ilRlSTdTp
Iewmx8TrwfGFlt2gDfJklpH4vb7aLTwM4KVJDp8OYTQVKhZEBviAMHUUCC59mjMt
xPxtBu5UgluK2HzbJqxNo0axksm1Icw5OHzMqaCaEo5Bs7Q5iE1ac00tBO20Gncf
sVGFpitfaKjX6f+EmORD1PTGjWZkOU7LnYLJZbLJ55XEBUMkwYXaSQSeC9Jc/THL
9tkCxq5kN85gDGFoaO+k3e+L5LCuEXT4KTKFB3jEZUfOPnOj6m1aF0oWDbsno67Y
lRFpLUl2Y7sFo7t/CUpZjoy3hRcQf9xDrNzMfX6o9/dezWPcP8DmxEkoOWgZkAzf
GSE6+fe2j2LP95mFU2ML/QIzcUTpoRk4mh5JoQcwp7JFDeBseKT6QcK94vRzq/yB
cZShj2Vb6ux+DUse56M/weqv1MePCLEQYFnTKX9zA/QQfJQFJ/JzEhnpLNNbI64+
Xy+/UBaeiNmzYFVe6rHyIlMRGMbHE4qN906aVj2vdpCeoj4m7Sz/uLTyNhI0IEUC
zxrG1z2exOBCWk4BeDUPfBjuj+aNE5S75F5P+GX3ZtOJRjspSkRK0CdlnYxft4eA
cC8RrY+JybgQcUFTny/W90y633TdFVueKBWuDTa69RXIxy5+EuMobWX3+gaEQtUr
iamT7xjQxju91EouzAxXUv9EPQploJbIrEb+07zoCPdJ9bpbjQgAd1Vr7KpDoE3W
bdKFKoD07uXEM/LuLTgjeBQ8amsTQEu9h+vWaC242bfDoHwUCH3WZshp+qR93gRc
2T1Aesbyf70Ll5/4eHkBsbRCPR6HMJ1EoI1vxq4Vn4Fot1r2yDzdcJTbOJt+noU1
SkebV0BFttwup/b5G2tZH5FKa2/kMkyHAhYY1PsQA6nO1EDyUni9Yr1KyK8Uf/3E
a11s+aHqZhNL0XwmKOPMa8dCs0mJ0XadKU069Bp/7npNWonQiEmw4C880r2mk9Lb
XiKK8vWvX0tahMrzV6RyR/LaL9WbRWp+dlEtw+H6IwC8q0b+Qq0Ch+xu2ir7+8PN
+XCy55R07BqCjUjpLId/F8kiVFBvsu3VBUpWXSu+ZYBd/axb3Pf4B+Mh/wEhnypM
RQ8RDA/p/43eyaB2qb5o1l6uvR45a5Esn3Al9ZomeCT4ntbJ2Q1pn0K7PpskObTK
RFTDNpijEIAvSs+OA/jfVpY5IJ95H8hrDJIWFNacI5g9VfL4FdI8of9SIEDUzvvC
qVdPS0wwkc/k1kNay8TDJWY65YAzcDWqhajKhbsNX+F7l7KRQAg9F4Kbe5HJ+lXS
NpRazX9QkmJW0YmtuE3GQe+L6m8jQdeniVOdoc1HZO8BUV7zk6Teyh/yjEzZRN71
ekxahJburLHnpxdiS/y9CL756UZqfo2HBmlOfYHXhSIugOe6DxdfCihVThTQUZF7
3qpujfSKbT7AWetJKP9eEwgCEZPxWFebB4uIU0IqgHmrBUyOx1HRpSjSaAWb1DoR
bq6UbyB+Dx6mdswCqO/qA/ivO3NdpVNLwkVcsHNRARPhUDmfGu+0/DxorJrRhiS7
7FE77Zmf0O3V8anu3ebNnQLnINxT834s/MAPPyYYy5jAC3JfEYOONrZUMTGcysMH
hHCAntb9OMscs4QXpXLUmwbRqzJUX2jKK0kMXBMgAB3ByvHv+tA8UqP0j4sOAh0K
vkeNw60dvjM8ygXnnQ6uaBlMaoorhNjq8yY+0VangOF603obmycwpJIkAYwW3Gs0
f9rWtMO6aOy3MY2gD1VnhGEU5QfHfD5YbvR/vM1+HLj+xx+C2EHejkp8dN+qaaMF
qh0i78udEcx4uYgp7dGXjmYv8CqwCb+Za0GpunwTvogenNxvaBiZ+cr5G02lWWJA
YeNNtPQ9RAX3sxifxXT/Mf8SUCeC96+IpZpjfTScC0WbrKv6oNMtIdYr0gKxJz97
fX9TI7wmAFSu0RDc48twtJ3ocFtiUq7cjjdGKPr7Lq+WJ3vXmWkkByr7j+IHG7SH
7ePqfIfCm4KDKPbZjDCu0Mf5OT5+7CwzmH5OgFqmPxFIRMRIthKmAPrZnxRwAJ54
Tkpe1zAVa/yG7WC01g4mAEQig5pL+CFk58dG6K+2m+1W+IioB53KjNbARnumQtPC
TLd5hhDajxob9sXV5TjKO/MadzJxPbr68WR5VXDdLscSzPccx3hgSTWePCMKzCrp
s0C5DMfkLRTyoAGGgFZvl8igwa4KlF5BHmNTZG/IM3+qHs+42hT1N9EgGTTpYY5d
dm0z66NioFxZuf19goZGoEQ+1StX+5djITOVXWV1lF146WmQk9BSZbnCSmQrGos3
I17u4DyKmG6NvHPxbPCuw4gT76+aS8tFVCh1oiK0xUinlSVvWvnD6j1K3+mv0gWU
2w9vtvEg3QjnTpEy6EjP/+BecHr6erhYQWCRv4JdrsK1614UgRhEJoSAuXgvEBot
IBIv+Jz3fsBO8BcNbgVcYntRugo2DyiKt9f7QknqdS66fkBHYCX1fVtIt6pPTwMd
C5wIwr0pbE9EEUX00Q1gZv2NtOX9cQVd8Gg4z2LDDQ07e7Hd5H4imSzfHARo2niw
+VND0+03aLLss3WXUMU13ouDvJhZ6V7hKE8Yj+0xpbI6Dcgz7G5GPGCuCf/TxJUS
ciAb4KHHH9Ye5PlkQD4ux628HypYcbX2OzM9G6/Jdpu/GaoJ7p7p5P6+i7JFD3lQ
zp0Ik+wmHlcMGgsH1XGhtzh501Ff31IRX6Gbudh3iv2PFIyyam6jh7wtk9nQf5lD
pUwuHAAQjNuKw5+8fn7+D79IQDuXWpXwXc78+vcMFsJfczfsC8QrV6QSQdgVf/b1
S7YDvzoTR/6WYPjx8VR+WDYZRGNSUifyg0KW4ne3amZhNY0wgPeSvjMg8UTKuL0L
0LNaJCtHiW1f5xu78ZhNGFoSiUhWZ8dwuhU9YL4T+5KZ/wmSNKGPW5D7wItT282K
KcgGn4u3cr0HDjmHE0U/zMXQSd1dxueWId53gCniLkoZ7VOD+pCU1YST7PsM63BA
mtLE3sZgHDsdbcPv/Bgeeb3wy4iJIdlK2RNbnZbjzpqLnT86j+0yZ9CjkfaR1HIc
SMDVJbQLmgDXTkQKQBuOTNyoAH6t7FyBB+VGtJml8YjbJmMrE8oOE2I9Gsf5CWVU
MoZpM3qOvdGWjxKdFrkZJ1Qky0mGgTA06UNdFC0UiG9+D03OTi62nLVKiIpJ2Xkr
EoQwH5+ryIruGj/4QFSwE4ZIsdTi2gNyQYPycN3jPvhV1EwnswB2KRbDNr6yIk7s
2Ax+j/Zh5Xlh+yc8zBIBh1LeFr2n/kELreyvR1kuyO1Az2uVr1i4zFUjkKckEBI+
7OOLEQtNcUZDJxE7xmNN99EMygEqgdPDhy7o8Lh1RlvYJ2/L1RjlEF/ym6bzptFA
X0CnMekOc++XcLrHEurypmVvAGHabJHCbK/EVoVe4UOZn4fv0m7Gxb/QEgrSl/nk
OG6jVbIPgAlRymN4hKijPqVoY8T3Z0gnFs9h2P4mn4Pzig5tytNMZRKmYFd9T5pM
YDEHXmG/RGw2IfK18R2MPqe5q0voWYAJI0PjpPu+SamVH4+62dH8tR3y16woKm/Q
GUWPcQU8FzYlWcHuBWpYqIIZQaEZB1D/4r1TyVPw1qycZvCyOfKhdITv6/nr5PyT
U636f/ax2xnkSyfxV5SR4Ge1o3919nFxBp2Lbj3zvqxoViKuw+ytZMf/xsdY8ZmQ
8jUNTDj1tp2Eg49/huitHF+Ld49t/8LSYwWg+4FCMA0GuuC4lNjNlbX8B1AfBMp8
HLZxJM6Pv2/qA45IDcD78rH6fme78sAKgqRoofv7y+iuJUFZLirBE8BkB71PXYgw
hjI+lPMIvXUX1cHbY6HrFPMq6qDua7a1n50ECVp8wWrjUJ05+3PQsUeUjzQ8lLXk
0mHBywIbgwdH1uAgEx1dvG16z+nmEZRc59JyZP7oDTQFJYYTQwibOHRcYdvEh4ES
wQO6xpaS4O9n6UcG2gmvan1G8dZKkh/4Q4NnIrDuGblGdLAD/FHziKee/Bxmf6ms
bI2yt1PqvgJM3r4kXp062gRld3lLyXfWR46LT460q/rPUu1aKXBl/Y1q0PlEkVNe
dm1JOrAkwdpYRV9KIyxc0R2Bdd7auuCipLsp3Qyfz0//0pGTFBPWRPNvj53+RW3A
cIWD4Vkhd38KMeEWbP9LIWwZ1cX7HwPl5qUz0gGL+98m5nOBMoGUBAlse/PSkEgu
k2RLDS/p0MBg+0wvBXh1GbHqzZJ4FGusBP7PYy3ckAlsKLfBAA9sNcoVPqJivuMl
i6+z8+bZQ7+zIW22YLnWaP8R0KwpIBPSV2EL6b39KoTL6FhUPPWQnS+s//ZeukxN
qTSXp6TJtwP0Dvv90bPfPBQFbHTZ0MxRmuqoMyTSxMCqN1T8l8BPGe0Y/UseBMn/
XN2DXPPB7KUGPgCLPymnad8gkEMVWbaxds9tB/Iv1ZZTo8UzKFBz9njmK2IlmVl3
5amzj6MDhKFFZ+Gom5BAIXL8WYtnSzkM6H/yfJiCJPkEmZcavhtgV36zNp0YWMIV
CLFxqhpewdB0x7suBgASmNDDtadNabu6VhjCq7ZmlZBH9BcwsUhvPHv3esMHrwEN
MDkHxfQ3zfjpSED6F+RL5thUt6rz6Sxzl+3qzidq7UVNMYzKl/nHIjxgE0Y7U7Jp
24HlmD9JP9lUy/zbC1U6bjWI1sJO0boOFBqGxm7N9DOYwe2OcguOrmlZNWWKVlZv
AUjvGoE41omNnO91Kvi6fPD7tSCin//OlvylljxjpriTwNj3H2mtwFSoFurj6nNf
b88babkFnva5qdLAPjRttkvKMLcD0MDiA+LwUpJ0Z6jmDT5TKwoOX88X1qiIeZLZ
T+QzO9tvIrnTksbaxZXkTLOmJgOZasjKpAqKYBoGBQlNlSxKStou8cLcuInj4QlB
ggRs3JoIes9mVprznChAiLJHRocOwnc344a4+6XfGu62EAV2bg4cOoXrMNdr8YEK
LPzjASA+m+UY5+LrtvU+kztUrIin2XkX5HU1CUUVgcILMuLyx5UYAywZRd5XxJzC
EDXe5ByAOppuIcEFRtZFfFIVdFh/ENdbEdkiT7XBLZ5Zb8c7IVjZl5lAhR11LgC9
7DaRHSJZa1VWjF+dpN+9KPytiSvSoKh16xt1gUmaID36hnrGO17ieqChh/7Tv50T
irnCTwXeB9a6raWhxfaUDcB6wKPOHR/DqaOD90luF6dCSpfU8PZiwDsgG8Ke+fVj
MoTDuIjSsCS4+kN16sXK3809L7jhw78BS8i0ZmlQjwPwMjgnshBputZkRFXYEso2
6HS3+t+Ru7rqPbVjnfF3lcHZefMqgKoo+RYYh5iR1B0NzbE/o84bNL5Mih9XLnoy
/pi6vYx+ElBeWapzUDkn+QsrucvbBuuU7bdtC51vMH82PziKF3XaJCcs888r5z5u
WTcXiYIOjjemH2aL4jTlpgHBwp6PGTza5dXvWdulAYLZ1BbeYcNRmB8uZxlG3KJk
GFYDbf+4v3MA3wYleETrINeK+2Di49VkmPdpR01/1JH4B+r257M6fOMip3OZvzz8
n7wX2LvCgehFwEWcqWDHM5wquwWxCnIaRBS5NKyS07tawRs0rUfzV5UG7ep/MEsV
+FBmJaxJQgfIRotANvDR43q5X8X11jVHtzHCKv7WBHNg9tEJFM2rwrST6HsroXse
llt+zTLc24Mmdd+kPBWTlL1ZaLsHO8M4cjVsQGpAgacCMS0ETPV+r8g7u0qCp9xu
kFaSX8n1G83M2ANFu1sEqOnS5NXZdNtHaCvYIuWEkokV/IFDOF8saeErqTOAS6ka
KuCwUR0DzGxslAoevmzk8qJ2HzgXPjbDUWbs4qDGTCwotyL+xxekqDj37UyC3kXY
eqcqwO5h8s3ufAa4MSCpsyeLlNg+0mWhuCvsog06FZW32kvMMo6BeoYO4Mrezral
EmtewgMb3MAtksDXjYy8gSTl7i7dxnwiVZdHBalCF0IIGulTw3OwcDL/cJn3F3ZR
CqBGUPw0tfXE9XEoiidtw61MpDyRXh0VzGlxYUMTzo2C0LCt+HBE/b/bHppJf20g
gdrRjlxwkGYyaigX1keCeo8UixNCd0KqOvT4mL7AKs93GqiGJi+0WvjJgiECnYkG
RIZUwMvP/x7YHJ/9848K1kk+yT55+foywQI/zSZUBTrN0Enc0+EWymyFpj4IhlFT
o4ii4d/KZqv3EsJCy0XVHbrDoLON3d62LBmHPNcjrKI4s7ZXGt6WOmjOyrCmFsh8
Z+eO4LwIsXL1EbR02P4ieG6WpmAyuCFkEO8sRJmnDjEbgpUe2ZUyK5E7kqVCxb18
mSukxNca/M6N4R9zPggVBFLNIQ6n+oiBA+dwvcEEWF6JA+a3ta0+WfG/2d6chxJi
cnHqD08GqSJMODOjqjbA+DhYzGCIB+9thiAWfmV4fyk/qqhiCUPLvNwBNqK4HDm0
SF3F5M/xiPodvNHgsM4RN4ug5+ylDwnUyT7KsNQIgiAcCPW1tmopQqZF9By4rj/y
TKaHTCHgOikUxB0gz537t/qf8lcTeRRQ2nc1f4Uu6QXCnftdbbecHDmSyuBYfR44
CE7M1dJd07UG72RIzwCuX/Dtk+0XLrGlZXXF3Rbu8KZkrLthTPwNm5nBvd6/jdG/
XXQ4UWjpefiJ3yd9d+i0Trv6SV/NMfHU9/wAIf8BtKCPgcnxZODImcbKjazgwa2z
R+r7YuGokLG4Ia83YwociG4OxkFd7WfbKLqyRWofXqnOlByhTgE+Kfsl+51/yLga
QiTntXfKyWlTsnXzYb6rQXHHZXl2Y1qpWmkU35I2sGr3GuAmHqii8umLEX9B3tBX
8izzclQam2JUdlXdG4pfJb2CR+AKAxVlsXn6+oK5NgO20YQ0xvw6DvGF5oaQBOSu
2eHAz7dPV/RCltrM1g5pwV0Q6MdkGI9ho0jg22pP+Rc+jfb6NiGsSUeumxEv0y2E
Nq5cdhWwNEW98gPEWTsyg8I9ZW0Xsyc35q0z1t6j9DZT3s1lTFjorTtR/HdpFiuk
T03Wk2frUIRxrw7mS6Gtnp2uHafrU388afWIpC9DuovLkpmXBQuujzOiTyj0JuTk
kajHvF3BtEuJhc8joX2RYJl6mq4C0dBKsMDe5Z5beAHT1zv945d3KEKZEj7FRIZ4
laMvHp7akUXTJpjYu6kuwSlL+OBaadmi2/nbgdjp4UlERPN1Go92gyxpEhBct6vQ
EJToMLP8slBhXyUKX5jDcSb3pcKKJRi0MgP1X9MFP+wZntQwWtnTSIl1AQcsIh4O
sjMkkG+oBfOKkK8sPz0OxpbKDblNdk8MdjFgb0pGnjEsa9mQLTDTX7Aa+ZidnRIu
ekVbHtsez6p34upvg9sAkHStDjSsHi64roWvANBNKNYsDtUmxI5RITN47wx0yvim
2eom0lPp5z8kOl7tfkS9jc70atrJf2wyVlMUGcaQCcA/VfUTW9PSEvzjwFFw6GFF
a9Y5iQBmvkFhYfviYqSoRNTGr5MFHOfhuURp/rf1r5wcTHn1GecP4VaNAxSbIFgC
sduMbJvUZVw1iDyH6y/oG/6BGW8xZ4rf/TPTaasxMcBsR1jXQGmWqqrYtHjHFhly
IDt/MyT9vg9L/4k5DDQnNO4Dj+vy7yfrYFIT6530p9PesLdbTxp2PHFGsgVMIXs1
Wicga072TFu8AU1DK5FsqkFqvSJMMqtWRcLS4w+j9iXplHDHR9Qn/qBDlNEWUD+I
h8QjI3AA+fLynxcsU1psgDwg588ZRPi8PPxmLtaHQTNAL7MgA1V7vAfcFLlnzURN
o/MTdcm7aF+R0YrvwFmS8Fnil2bHo76iX+3rSOSLJs+VnDa99xKXeH5E9OUOt9y2
a1ZrqonFiSI4j66D4/HoEKEnDUQPBySMwgX7PaC+QqRSdd+E6x5udFVkAi75peL2
RkPT1TL/WQEjqMyok7rA3DJuNY4cRFtf0etw2TZyF4/Kv7HURgXXJ3A85J3zueIK
zO2HlVCb1z/h8NTdVB8aVd4KgYFi25XVJfsXNhQ/sW6dZUE1FbDdrd+kpNxM0a+3
8Vdwqzsabe8QBgjKij1oEn+eqLpj+FpJb/wmgMGlkUT+e58ywL0VcCtTK2woOJWo
q8GQT0QbY4sK5koHeIPfkF+YYvaPnxda5iwFC6psL1z9yoIwlOc9ASLx+TlXp9cy
0+xQTEpwMrtMYuWhpqXxHP3ueysNif1x81e1Be47m8v+TWoOpUSDbYSvrhAa2mJL
YDtCgL1z1zKxUYQGz89JiHaezawgxB/VAG5xH5C2oGCnV4Lw8c6iFnzKVP2Fohue
pOuMO9nywvxHDQdWkBISL3CGJzzY32amon1tqsRYyZoFUH88saWOsByP9Xz8hn/k
p3t3aNxh6Pg7YGcQABxi2CN4ojanyonzsJh0uyktJX1mDobnrhdt9OI/2UAYAfY3
iRHf8TrjQmIOPqVatJWsaf4twMxXv/6HbzxusXCudFeIsK27oErtQoRR3cAysKUQ
LfttpzPzYdfup/xbNCJaCIw71l0nrqM5HymnpQIcDQ1ClVAWbfB8kBTJpbEK7eF7
DSvrJ49BXzBs8vmgPOclbn9eNyV6n0y9cVaAGOzCjLhiO/hl6YC6hsz1TLVlcDI8
vwgMzyn94IqaHv+LvieyV3/GI+HK9kbP/o7ktCj8vG9x9zs54hbMgju2ckhUeQtu
Wku0ApB33j5zXu7afCZGZ7lvgX6cwmSaQ6Yc/Mc9JljE4wK8bUicK0pokzwrAAoc
xUegYd0h8w+1xp+RiYJd95rWzYngRuvTIeUesCoxzyp8wrfMPodb2UvgLBKXTPak
51C/etU/a51N/PzvNjOhSXE2ytVAraWrPTgP04zRXH+Thr3q8SQQazXJC23FBBtb
66GDCuRxF9x0cVWO4MlV80s/5ohYL/Z3kr1gWE/7QSrBfM3QkqtEVvDZxoS5a4rP
s/i8u7qEmvMo0Dup+hQXMqZJTER/55X3o/0AF4MehRuEsWkKo0UyQzlXPMdSDzf2
+mB/f6/VG/c66JqjbwJwRAbUEfWh3/NyH53O8SCiN+PftnvwvQMAPa+iL0J2NgQ5
cq6irFxuelShTQd2yFIEkBj8SbYWy06xC58DzkEfdblCdK11r2972j1OO1kyGZac
rIa/Qzq+VIlprDemr+0tvWIVkReqAkg+LefR/OHtCa6QxIar0sCF1IQSFMafojaQ
OPbbh4SVWywL8RlMPdcO6OnHeCzTBNiz9ZYYwob2bRihLc2qb8xq74tKqSzqc81A
jrLQEsJgEHdtP1uX3zlW/zcOdX8RM1tsGk0sJz03rvPiab50X39c1njMKd7b18dV
XvXQvFwf29Ruunt1yMD1ywK1N4apI/1krLW7SC7yZoVXFUePv8tbUE/SsIb3CbBS
cMa35ubx3x+rkj8DFjVw1KR7WxHsahT4Ke0ZjFCLB7lc4t0R818tab1/kNzoO/A8
dpcV0YAIT5YfVtt7Ya579oNqz4qLbG1CkrpVXI6eRfklHFAjR+PKn0iqWwL2+6Mw
riTHSjJfFu/p9mCfUI37/w2o/ytP2oDjQW58KD1L87yTAD4u5z+Jh5AymqNCNX6w
qpo8tSYuErISLOSyQsk9i3fAbJyknG17Rq/qD7BgarhJ+o9MQvIHbl6DPk3lSe6w
U4CBfu9Z9xTP5OIFZnDOTITtIwotVV16qVkBRtP/2MJCHqBDHIf8rPV2iZcMFIkA
PhZ0gxNi/3IL8s1wc66JuHDz0vWOsTI6a8lnHYDRVgNF6VFc4I9tG6TGAnIVNPZG
H9/y7Kef65FbU37sypJjvmUJkTX+hGOVdngmGiMlFD+GeA+Hl1BTrHkCQ0gC6Wkz
mYpa71fyF49ZCiEpo4qVWBk1cJJssPnp7DNfD4LhmV7pv0ZcDUll+g6bTeIGrNjZ
6OKhnV4UqPgcCLE5LIdIfhsnyz41bFz088nSB8QD1fJNTSXOHKjHUYbx1dNGMRHb
JjtFJ8Uzu8xwSz2mPygeLYptFrwxVroCEP5UmkgXPsIBZLk/ueJ4/AVvgyCwxdnN
+JjSmRFPvPhN6Y15GMMIfHyAJsNMzL2p0hhKrv0NPXV8LapqGiR/S3NNPo7IYM7T
EKmKdqDYzKIyeCAbNv7RNqq6PprcgkrkGXftPVtiEkxhg0pHf4112h6BT38/v+Hd
Lg2HdKoeBmhiznBaprB6+ey8wjuUvR2eGwQK61nn55f4tmf5lekr2jHrNTzCfo0s
UDO+qvd2wLnZO652LWyezlrl1l6WlCfcqr+RegYvSq2PU9cDNGSCQDXt7kwpX8Jh
UeArqrKZhfXfvl4HlTKIJzRShXGNqivNVRS0uqKVPK8h9p/HimBWy3ncEKu4RPSy
nlcUsFq9/RWTy3bijcy05ugF3H+/qBO4vw+WQYpIqgkuY7CPTzr327sM1XxBA6kl
H9Jd/feMc6rEophCmm1xkrBpqQy7Gjmg8Y2t0M0hVMwwQ4uUYaZidXjtVSIrqYuL
9F1PDQkWAt9wt8fH9Uomo+NHoRPqxOSAqynwwd8ZRRD+1LQ9RYbnW/dosP2z82zI
pc1YsXKxlZBEXWy4bX4DqMM2IiGkz9Pxzs0KnEDBNldO9s0BlxwFQovj3xlDmjm9
AcjWe2uHz8CGtzs1Rs/Zq+EZIIfNljnkbBbGbXvYAUfbPEPaRMqf9xKEXjLjuCFP
kvbFYb0IvDNq5M6Fshju8LmGv1b96vOBUlMJSYmGDs9KQw/jFAS2eubawuH/tWq7
24gQK3ssZ7aWp4xokcc3tFuM+tss+X8l+zIrVbMOGDYXv5t6pz28DRbLyISesj4Y
Ri26uYDXSAagPp3EfyewbJW84l3etseiOVkNwfZ83DnCnmxsvLaLAPRN0kpyDteI
qzFYBA2R4mk1G40PhFiHfiUjGPKUiHBKBXj14kIyfB4HpDZ3d9f5COOeqw+yx3X/
g9ALPZ2oCtlahw0FRJoddHkFyQLXD3qejozpSkrXYqnmtQoJhu/YYHwTjjPzscvO
ADUWqN+jO+nx2puabX/k9Aqe4GFF3C3+d85RO+/gP3H4k7vCFUhI7yenQTuvxrRh
F+67kZG90fdyuHnbeB6vfHCP8anFbr0flDOnT3mySMAvUgiB3ZGV8FUWEkW32heF
kDo2rPawxe5wxEIE3XJc2IVj43lIGhy5WencP+lMUe7tf1jm0etw+VUMFe4Za6f7
bsQgXhJ4Yl9UJP5MXIvVXYcQoa8+zuUuDjzjCsWHSmsKjOEFm2wNHJLvaY/W//EN
mKBC89UO8pH4dSgYCv7ZxFtW6+yIQU0M+U5tIp9U1mmYaGxZNFl+Ole2hZkAPgqQ
U0iqrlVW8LpmR3AURgSDm75iZtiWxqMK3Jo1xqjWm6F3ggu15jomocr7FCY9aI+s
0Hp/AfR8SWa3ex2SBRdJR/swubacSoqzllirNcgjrtbS34EM6q83uC+Y9myCIV4j
pKy5l75Ksgoxz3gXFWnQizPI2EHKVNnEU7vdEgDq0YN4OYl++wmw0t0Q+hiiI9vX
O4Gs4rwfmCUIt5q/JJm1yDpFCjQJD3V9muLP8tFHPDv2AZaJ5GEWaTE6nFxsR/vZ
gqoUY2nPS3mOmE51G33oeNreyJhTRU96g11/dNzYiGwxI/SZ/L2R/Q4HrO6Z+POD
JsiYc1iLsewMNCh55O+vVWifB53RroTSng8a/jQyvSyar9dnisbZbAktd7CejPG1
EDWUKBrxmagMoTnlMjlumw8NGCtDqugI8KaaftyPchjqWGyO0a8mqnQU5whtKR2+
vGXHVfzB6isG+tb40GjdzX2+pngQYKaQXozl0wP+lmW/IAiduHM2JQiXHCBk53AN
3JvEHLSsxxBYld7iML+k6zFlsSGUj1IfCuZMmLA4cFfOZjRKZQ9fw+W2JKJ49lkX
DCXMeF2YxhZvtURi8/Js0yn1Bk1fR/a48XDrtlZKRPHfmesCZaqHGkhuSaLMP4mT
NLUNpAMNLkO1kVpeAaAnxm9iei67Mfkb26ropcy8HDsvHN0G5yEAeJ3WfG1MzoUK
rlaJ+NiazR9XyFuetYU7d75uVqBgh51OUvwYghZlb9AlBkP1jQYQRP0TDlbgSqQ8
P/PoclHr0ohpsJDCVDzGnUqsLo/di7I6RCt1g1pLKFMFjSgOvIIlnI7WvFwjZcvV
+4XIJnMNk3a01P20t8e4L5Lm+sS3f9ZVNqlGduDtAZRDaexOiy85VIQUd8kbnpv7
mAxqX0s9kBHD7dA/D9qiAjt9+eoI1KPhJrL2GCxoqnQzYd13wiFLWoSdLdp+Rr8P
1TQXjsPCey1Y2NuQcMvmolpWtY988Etxq6Q140pZJLUh36tHC+JYcrzqHMTJN4cW
z5z9LhTHnqDpfcB64nMgbyGUOBcnRilJJERCKKVUlOraUb2DbHI1ZN4C7TJjzeEH
leLDhrQbkzf+SEuJrcu2P8j+gSMTKzT0W/ptYiZnFARwC61p4ndUqZjupjN4hnb7
0rVfrzLm05wGrvl5RLxD8q9BJs/agxg4UiEBsHXJ0FiLPCkuca/cTKqKY6tXsc9H
VQESIcdoa0J/IciFkwfGr0EjIx0tjkex2SEQP8502uGz8HDS0WaMfdSAfliIs7mv
PkIOt2IU5azdrJU1z/Kcvmm28otRT/H6j2SydxLK+uft51IzXplcZaz+Ll471/1D
t1TTwF5Jj3B9OkxcsE5npBHHvd4an341CnwzBhzzdwpN89lDBs6cYA/7vmmN4TZo
Ou8R6vH5zKjUZLbnYV6dr1KJHMRPKSQ8qnz86yMhFUG97DP5hnSEo97ZPxXj49qY
xkj83LBeJXD+QwWgKK9pArwQqYwAs0W0PDOe5VBkpVQJdXNkOVa5gpEzAXI++P7L
SOabTknrmKbOnwAvTvRpiYlCKBIybcKkY0liPdqsJPD1z0vCgX2wWuiRFR1CAKEs
/YmBGfOdaKtUw/W8eWesYCp/sO/tWz+c0YfvW4CT2F4l1Z8bzGorIwHeubs9bQAh
wLcYzWkDKg6ELFnRUu97/mpEE939gp5wgK5Z/zDNuYnI+nhZNgtDZL6ombgcGiq3
MIhFrFd75Gj7meAM2zZ1omqBZqRAiD/BiWMxnVaXEPh7TISSNWEmwsa4U5e2X5dR
B4OVdPemj6enoH5k8xRcigdbbiZWhnHTiBtjwJrBg9ZXtzLmLPVbfgF/4TlgpNV1
zj6jS1fI5mKsRv0P5nwOCpDZycW3fTDcl/A1EsBsImwbo4tf7QWYAL+ylHxvSYuY
eESZQl7MjoUhy/9bXdk+XTL+wzjezFhp4p1HyxXJFbKvXZtDriulWxWJ0KQQpnJE
iTa6e6RobddVeqlxzzglMtZ2feqrnbJO9nzs4q+ZVly6mP4W4YQcmE0DOC6MS3+P
5/TnxrxT4KZXyVqDXxgP1Bwwg9bE7Q5RkuB7JEMtcScSwWaRGOi3nIOyiYrAW9Y5
4tfr9e1uHF5iyWJn0pQ60VqIT+yzHaNH7IeUs33pnEEARKUJq6mpfpLvs/Q2sMrh
GmBDaDlj/F2XtYK4HW/DLZISqlg42JVHkdIO1CoN60S+m9WnlTyvSLp9sNjz1cwg
Qbwjz5bj8esA1Th7kWOrb7rAUadzStXsOhIKoXgJYXBjMoGUV84Cmi1u3uVneNbP
cex50MDOaNXJF1ZtL97BPkaCiAtH/xIZzYct9s9xPdje43GM9DKL/JhdbNbJnA6s
p7gwJku0QJbJ2A4/7ywwdzXbLY0NwPCNSNZ3CODH/4fRneTKGWKUIbXCxX7BzgYd
2VCQYGsX/VoSTkxZI7Q7uW1YvQehYwtTndDUMHkOUtJKxxHh8MFxBukcATrt+53w
Hhrh1CeKY4jXTSJP5ZmF6u5diXZ2eHsz9KLQJ4MR26OYPe1wfBB0HtixdUHEnXAy
pLk+3UfEznlafJGKEiDcyjsL3BycdIcxnmh70kZL+QBNtamYqdwcmhe5Fo5fAd5K
7dFi+GlkHzxA6Moy926xgo10BElqwn9ck54RJd8rvWH0aso0R8k3HHwMPlo/UNJL
Knd6Nr6gUsU/lCWjtNhfoyF0pgvzcjAjm0epJEWS/j3RRMDZwRLDcUb40m7YmUQg
s+nYK6tYu8pmlDq2k3YBgzB6fhUTd4tK0RWAJEFNbVrS3WRcjuq4Nb9yc8TcIwr5
6z4uOK3WMUJkgfXHkCQw6sLcI+DSKX3Wyw8U98TkeyKhJGkKNtsiE20AgN/XLmN8
/PCbUm4kKdAMOpmiPvGcD2NnbHAc2BXG70fSiUC49H0iF2t8i3tuVc48ibJbfQxw
q3jiIndvjOpAUspx0LPxcD6phRKFgp5nfE+DHENxLMv/ODyFe/3YLdekiI1EwFeN
85QFNODBw2gHCVuo052Cgq9TzPHY8MvEMoJSiF7N6rpOFr69JxxPDjFciX6FZxE/
D8CipNUmMxs0mQfzXdVtTki39AlsSW/dSIKFsIpKvX1rDT0RTjoj3McZKLMTXVRZ
h0svdMCFqO3XncOoNENH3+eEEZ/iK55iGgCp4suCNWSnbPthpOaXDM2zF+Mh18G8
RmvvvNcu7PUcD1RA3ffPWi6FLuTRjMp0vdpx2ouEkVvbZ7judZ0mgwmxJNoKsuzT
+ousuHgMul57lIKX4SVPHQK+F5Bn0uXUN4XrHMgef4Q0NKrZH/HLfoXx8fpHJgVN
SWL2UvVpR3QYVM6eMa+jBtRfgyPT2KcS4EcKkjpXgHWbS2p7hvnvEDlFt86YsvOg
Yw4KzA6Sj2r7Q5VP96l4I2GFL5TNMWsmvh4IVPtQw4XzusHAtBc1ysJ4Plr8icsk
hI1EXGWFw0hnDX2U+uHkhObxIUZ0GjKrp3sOjke0dYcwXLXrSjbaHQEo1lv1Ani3
Lkm61htuoWt5JIEBglvyjyrK0/6NxgIEUBMogvuB21X1YX6rHhqKSqvLpQrx3OEQ
gUUFf5AQgN756NOdnTnOuk+dlA3aQj/sXHxDL93J+RKKvzjPEogK4t+bpckj7vXh
g28pywbHI4YOeCcP05BWGCdmGl0Ijr5yu0/DU133c35WiDKkQDagknrHa6+x2Cw/
XUl38dBJRoSntY5whHFg+eqLxeHTbyX3+IL6jC20bso1Ikiv6Vy0hKtsgQB21Eit
ZyEmhyV0naV/0QxzZyE2Z5GRVbCDWhak/bXGhUKsWLa7ncvu+2q4gUInEFPql9V1
4FdrhA4IxnqSjqCJUDi1B7QbToJ/IYUdewAXLgGyAqIzgHhf2bnnBSQCc1RNwISN
iE5wR7dickWbBZEdlhDLh9mCXoXRMRrQua4qruWKbRS1q+o0aoSWUR7ZP1uXUbfY
dHB6dcADxsCrvK+VvnfFxVckeXz/Iv1HbZLfqPu6SL/yd++WDCLMCf5nQGO70BT7
dB+79jABln8KMJVQBXa4C4eJTCVLmZ8LGYl943NLBq8rpTHbW4mPvOcmMffdaMDz
kmDiWuCgtld24pfZARQZHyW7Vja4obhesR0/izCiOKJLalFCK0un9TD9Onw7yoXG
H9Rp5Tq1uemmWynV9sgjTeMtf//NilnQMMRlx0VZgBORS0IcPePNPyhqA0oNPk/l
/KfX8GI6+xHeXSG2YbNuNBlGLdBuLF8im7wzzHN21JrBhT17ahzFurXP0WzrygnF
TgoITySalv3CSjUVT19H7/V99XS9ZVN7qfhsKQ3bqvS2g3ao6PGgy7ET1yBy13Ha
hp37IST2SVYTerzyPoALoGTaC1Y/c5kctth8/PBUkV/s0WC1P2+uA2CQ+criZFgN
fGzkIRHdE1wS53nlO0bGQ43AEUf17KkhIXDpH4ngWlgeiDxVd0x//vSBlSv7/rMm
S7k6yGB0qvxvamBR5IU8twHM0jEZT+HaZG6SJBl3gpJ+Rig6l2SJ0HUWY+hbJkD/
717eL/iXH12FYoes4uU9MXTsT2qziptfEX+ltJ7isVAx1T3ZTVJd8UCT+0J9/oFi
K3o2TquUwSEBzC6SX8kfXULeY9TkE34ioeCdoFPvS05OqA4UZ55d2cYoLFegNeL1
dhQ7skvUChN3WNb0AaOTt3W+bUt0MxpxuEodeGX+mZc4ZRRzMj29Wzc83Cj+bfkp
eNK5hCJvC3EjjrG/bTK8SRVZ0sBsz4mpyDiyRUtbrghLnEetYrC6j0umASOhLxcA
r47/rH4wbyQnEfoCwlqw17aRBcH1DtRWXLERX+IBs2Zf91bsvCVYWdmBDbVZ7F+y
PJBwKV9QiAhD7Y4Bl4D/H+HxEFd+SsBWgNCzhFaG326Kc6lERDgslfG2Ts1doZ0/
j28w8nNRNnBOV9vRvX55BsUVfkAEBUY0BLTIK/bnAYvrrJE21OZr/wIdyeEzOfyk
8qPEybPkmYbdr0UxsPrH3qnV6Ji7XarCxuEa7DhjxznGZ8RZ4/mxeE/xqeMlNzRW
4OpQ90ycAr+fpPMOOgkEDIMqi6gNd8IMHiHHNxTIGnKIhFfiUxGKNh1zu5fMtJ+U
VBrgEiCAKT5XZCCNUnyQv0gmon8rH5Yz+1AP9QN/+CRqstvPfN8W7j04Tcnp8vkb
Ny64/kKiknE7WvTcF7zvYTu3BI4eWMcWzPjWJcErYg+FLSF7YI4dP14uv1RyUnuZ
PGFRAb7jzkOGDfFBCztX0ebC7gOmYgd/skZTUGcTF8NIs7taKWmPuLdVu96W4vo7
gXAW/+oyWxxBYYkcEV6ffh5ZBbF+WRM7HN7tRS9FcJdETr7Gq4LVGtlUQpljtpxk
paX8h+3qSWftX4AC/+DqpPFoZMimwv91sYgVEH+lSzOoEcYeg58tZyI1n8EPAAqK
3dNkl/14D1XNKRYPCvSDbFvjz2eCWQ64lCWZ6c+VChEm7nA7pvmbU+0zeSOIg5L2
W+TV8q2PKfKdEWaiTpOYfyBVPtwF2B4SVZLWQcRu0Uau2/MLONJPMs0ICf+tgm+t
ATASZrNL04x0JSIZQxhNHa9XVWzu1wba2Kt/VlbLHJkeZVu1gH/3KMDZKHHOO7XY
CVx2hJHyCrZB4MsV5jf4nA5t6ahc2eQb8pBlCn1qhy1XuLMtRAW+vhDI2rtJoLNH
FlZFWHYJwb9Autvcc6Zh9UEcEd92ieZrOPJcBgedPu2BaWPBv5VXeYrH8kKvJxVZ
L8Jy0OKlGN6EcNq+82iRcZISButrEAufGJDdqFQQw0K56TDxo13wxFGJohmobq4B
K/shrxnvnZ7HD+nWKj5nh24Zi7Wt4UIgLUvsLEyJ/Ki8118Zbd+47Tue7dB8QpkB
x1e+yhitM/hkRzhJhX9tDHSEqPintLxE1a5E8FVvGqnP+pFhmlJ8MFDuvfTOAJNv
xNig0pETDlJDCC71OkoMLSKpK4EOPttNgdIAaumZ/WLZlIgManhw9Rhe6K/1dDHz
JI27nmZDJNnXAMIpO4020tiO9AfQlqcwB9EYiAJUXWoptABMJd113RDwpaNI5wN1
hPR3URYdlRaY0YbzP4ivAxoLMYzsybZYltVC+f7BOXtjVSTDVRvJpo//ACjtaI2g
ve8vSevkwsHaUYXAWdf2Q0FOR7S3C96suO7fekF9+k0xBl28CI2wypPimxo2ohls
R0gT1X1r5wqfqSHDZQtLNx3958OgD9inSFW3GVOCy2DI8RmTxywV3/97vaD1whqD
LGqsLyG7hsjWWxhkxrlkKgFlLMBEbbof2llIG3JMo4U3AYpzQfo2vQmzOysRgEl8
OXtstK75GsMBEVVwynXnkljAZX0w/BA1ACGXXWPF9w3YWL0mtBTSaeAw9HHjoEou
Pv2qtq1lmBtNS9IcCRQUMk2OhQ82HKttIsqV5BNEVvdbLb1q8F5qC7RDuH/NqKat
3m7Dvf2t+KyIE7CndJurUXd5PMGaVXa7eWFK4NqNlFkEhBXT+q4rLH7cU2JCdm2d
xh/ukaw5kM0uSOjTbwcBrkf1sAf4Nwg4alULhRSPOmGw5dgIPHvBAH52Y/zlb+3M
g2nNbCz/QdKueNUiZTpeCw7ZFDoWbnvVX07A5UG8HipUVZfAz+puy9oBCGcUWySN
XaFdHyyOQXRKLbYjV8QPCKe9finmhPeAzKM47YszM2V4ZmaegIFHAGxXVBCEJYQ3
r+ZtBaSmL7ve3jwon3Ut1g+L39gibQM6t1kBNr/BVkVNJofhEM5bbJpNyt/kpQFP
0HGAHQW5N/20sdtHdJsQfB0Fn1hEL25acCN3tDKHOpBrYC16oebUpAIRKWqSoXYb
G5wiI7nOYhkWtFPK9yccUtEdn0eFypasI7cGQLjzCjrsUp7nDJWcivtX3hyPRY91
agHDSL4AcIvJ7nOtToCBJDqIoR/uIeY+ePc049++ZLaUJEIJNTCw+X8E3zjBv/MY
CNgizmJxJak0QbsWzUkzweaJUjTXojwfwRTW6Tsfzwcvs0in6d/3XH2BqCWoNiDZ
8qkwdYg3Xpp/VQnTXUO2eM7/ehmaik6bI6yOB6/l2JmdK5SSFUgBi1NShvoM9PF7
EH2BM+ko0UuyqkuqZDIBVrZlDo52MWPIVUEwfsj7C4C+pZK++0l57xx5RPmc/RHC
XCj6cMgj6HoL4HCRunwxHjfy6pj2E4gGor+Y6HwoP2f6cTj6cY7OU10lsRt86ad/
qwPZl6nw1vdB8WURDT8MY3S8DtAhURJxXMdw20r84iyV8redTT/VjUBbd8XMMHsO
Mt1Sv7qpUI+Rc55CeFIfWubkW87hnAH1fJOdV7wWiZbhCSKKgCoh6feL3BPn7RkV
D1aF81KOeqIKAGtHxk7myG4bbqIuPHZ58VI8qZkkKWrkxoM6LbO8nzetMTV+VZEE
KeMMBy5D4z4zdPRpfnIuQoPVOTNm2nOXJ+uQvHX4PlsivqC7UdkfwWOugFZ/WF4j
bw5b18J+1xFdLfgZLvXE0xBoYQUEzcXSUNJcEeH5UDm9is2OIIy1CwqEoM4YcLVd
S6qAFUhlNziACTwmhrmp+MuYNw2axFobKbzCBojFoW8oc2swCWieKlHuYOhVRrZR
KGjjoguisiqQv/l7fEYOejRI2P5zY65Uo+jMYJovPVxntIEV+Simf5aV5z+9pH8k
AXl7+6B7iIODvY+9llXCVDcqRr0t8cBJ7LFR4OabEwxfbhe3bQi/ldFXWzKvRHo9
2/3jM1UcjXuKBv6Fp2C9fCpUXtJWTENVoab7XT32/kXIb8dg1jeZh9MlD6+KjDoI
/gbXiReZfgr4WvHWTL7H+WRHjqkZgV62JJXgxIxxXq97hDXlzEs2yqOMwccceuNU
Q3h5cKxYtL5/FHf4IwQGOLnrdGHzOLLjsJSPsbhw8fd5BgVN3vsQQg4NZNboy10J
ULqc4GdCETkAbFH1AG3yMqg0w5c7Nkdoba8Pk1fdPGme6jEe6Vo4mIYQ0QNAh5uD
8JRxX0BrcBPD//uyfhbsRv2EjnufQ8qOJTFIYeAEXmevT4GReZL1Nozas7M8B7Mw
42NH0iInp48TcGcyBneiWnzqD+01GV03HWeLVu/GaFlA0UVEIgAw6pIOVW5uB9/N
B83kGjEoIcC84wrhL+8gIV/V+l0QnbYRDIVOWHg6BB9jFfPgG9fDw0yLBUgHH88h
yXKyjPySypKI3UXcxHJJ0bWAmsO72ldYr6Xd9zztoBv0U4LLZ++7GKza8QhSYsk4
BeX4OzLjsB2/wySTLqLr4JjMxYlrKZhUw5ZvkRdjBrccHHFD96AxOE915ZECzvbR
fp0FqC/i36lHNFzy972XXdou17a4yv02XAU9tLpE8T1wN6g8oyA9wWQhE1+gvVtP
CgTzbTEZ2hzBTthlx4bAw+XZrv4/BR7blNk5juvNtXyZt68Zvq/BV7NINPTcQnPM
sTv0rJ3zU001HlNCxp27ZxvfHrqyg2cqCBZgY9uaAZqkyRCCdopMcj4pRt/hNo3+
5A+bt73jKO6JdOtalK7dS7OUATPR8veE2yTfl1kdYikzgwhpuvfMhT82O4xOrs4z
TSbVwjW4sHyHbJKKvKeICMVety6Oq4EV74elCk7iCLAj8BiTDNiCH/5vJVTWN0lf
g3GIRdN3tSiXgbjrtobJQURL1SL+ZcrfmLVs4/8wMtMddD8JRLP6KHZVKQTqg5Po
CyQ7XttGYWiHIxolOE5khsFxAMd4RUZ3lNjoCRfhiheo3BuOM+4WJG41P4v7L7s1
F1JsK4YT9GSAAVTgJKcgQcKLKH22XRqFKQqeIZtD7kfQGXo18o7Mfd2FrjFMmqwe
diN2uW3GMflPr0pLqU8eDKBM1bWmSDN6y/zP8DhT0nFCtj1vuvGyszEF3d0T8nJT
Fe4GfpFfMNgZNsigfAvJcX1Kq2G4AAbnK9afKW7wJ2BamQNdTpznQIYf8G6ucNtZ
3X9cDYj8J5ibyMhmx27v3oTQmHbFjOCwqV0KlhMVfHMiGajDkQMVZm8SxihIheP7
0NREgNmiPEM8cIGrO4x/eDyij5C+wrSTCGAN8F1EqoAeMKcjweywM8ON20iPu/wn
bVmJn1iq/ecJY72hPy+c4j6r9KwEnS2IJRAwO1dSPWwlaMIgWmixUbu7YNBH6LT4
oYvegLA7kSvrcwe1c/RGD6rGC0rPMhz/aMvPY9ah91g01NA9+iNhPob+9fAUSJEo
hbQ1Rb5pB2kcnMc5vErLkgH8v6xO92CiB/znvhzI7QnRHDJy1u/zvVDUlQnPiT7V
p+8QpnbTcstAhprHLPukcvCOeMuWHzIK1dppxh9DcGzei43x2+C0tmWNpHo7KCIo
BFGNxLMeJetEDaTE0pwNn/lF7IADRR1m8klG3TJsM9OZWC8LDfKEELWFaVCLnWyl
mj+7WL6S2IL79ZGUKkY1vleH0y0rpA+Mnf94gehd2AL8PS9svSPZVlQI/TTTadbW
5EcjzqjluwvShDmlwTYomSfje0soTw6Lnkqf5C/+7hsePWfB0XusqNYHTmnp2fRy
uk+G78+R1Wg6JA+6p68jCj35hP36h9kxuRM05wIhvL18eMBHdXX6CFs5y8vDbFYp
WCqbWX4yV8RceXEO6OkF8KLr2lipS773hf6HihQUTQp/9lACx20DuUaZJDMN5XXw
7js15WxEYVxCv1d8ddEwQOTn3d+kkowmMSPBB9T5OQhxOZjGCMEqwKihEEGEhyb8
Lo6/hZtjsniItSL05Cne0sNnAEN6dTeK9gpFNQjt6EUjr87WLDBxeMNEJZo5PfTB
XhV+WujJWeV0lrYMAjdl4yMjhmVQ9pCCGwDFJMynKu1TqfRgFJmqOaeeY1bXU8VC
KQYAOsFDr0a8F/XGYL67Wnhzq2YiFWuQCkhpCBkxupNJ0fRttgd2MEijCRncr12x
mdmdSIfmKdDUykQIBd5g3BumQr8Sg/hG7PJuqdGVE3ISF3XJ+yhNBKU4a7U8WVFd
6OBAgG4K/o6QjvQCWdPC+mpoWfCZArAtKo49r/8fH9qZIp1/QgrF3mzf10boOoQF
c0nE3ppue8M1zNlx3DWfRaDLHhhnFS1xF3vuN7Yv0vYXHbH2/bmWMwwn1dHLxhz7
hQDMxile04/lfp24AC8jT+dI8oZmhANKuFJkvM2MGd4RBjo4VVXSvYCAkMc0vCjV
0Bmv6z8vaRfIrKz+DUlr/Iwz2yGqSK2giMrFHKMNoGXjyDWr4coXj08bXacvEZof
DMCHiL5JoAIVXO1q/whuTXZSKwmR+ZzLed7/ylF/1mmJyfUH39V63LUq37EoNaaw
F5J/ePMoCVDV0hErFgY9gWV9kLJgl3xUec+I5Fp2vbdUq70b0AN3GuWjciNR9U1d
AX6uR7ubZHYqgsSL5qJo73KUgFM3KHR3rgL6SfhkEWNakDNa/ZB9E9xF38IfIGe5
rLd86Tn5qU3JClt/QNC8N4YoEDJWkhRd8oroML3/7vB72U1xKnHYVnDJ5ViEcFbt
r/qKmlsz3LIiLBFN7Z3oueHGfXhCnRjL/cVdJ09evQiet33Ew9WvVhp8kdsPX1UN
k5ChUITg08Uma4GY3IAUtAoAxJxltvbvQhIGmcOo/7TTZG9qess8hfnDNMLPKSni
WkLwZ/kIZRUJuqEdcT4eloDSAup8mVKE8GXKbuMONxshef7vOlZAet0RMBYIEuLs
n5x1feDLnaMNXmZv6ZGhep/o0C7aeYubqWhNivaqRz96rRkteNpVSKt5qP0hy0MN
G4NWJKKCrDOxIMLgSD69mstuJz2Qe1429RfiKuF/z9BIITs5e+MmwCbQX2CsaHQY
RLdpyr7Q+QiuRTwSM2s/IS1Ee1yaRVTvW55WBSTGE8A5Gf+BKpOx6P1qVerEAUz8
6jspc9Rmdp5k2VP5uXvtdd/c17XHeEFV1UHk1bZdmsEvKz88cd8H78928qJ7LhNH
3LH+LFvr37hyXsiXx3ncsyZmvLooY0PCLcr27WwdAgzhm6lzUXjS+T5W1fOVt1Y3
YvhBGF1AzsB5UJGgQ1IatIokNpgybY9dC+yT8sb/i4aszU+3k/zvMeNJ3SEPmjM7
92XxZlCObsoiaJVvR5oIJgXkG6+KD43Vq2eArfaym2GLDOJCJ2O8bd3sYP5NwN0t
mK+qhZadK1eF4OOZKZuEcIf8CAtpXobffUTlQMZG8NXCVCv++orm+GIcWIXjGpHf
6nY/T+Kws5MXktXDchS1gcri0PDAZaFiR57CveNvsOetjMF5Ila02grZu7eWdCGq
Coj29EYL5Ar/11gOQNXgqoTO4N6cy7jI8DcEA0hvq4ivsaTYMm1+mGS9ylkw+7mm
8gWwU7cUhzvk4meSGmSYmqIDDoLaviCRlvBMtHuGtD6OoaqgvBfSJAWZ96XELYb6
/bEYn1iOriLv9AdJNuRYb9ov9WtAiK5efyS6o0o+AyEL2U+PC918tTBj0chFdDUY
OeYWUphYqu7lqHad3/LtmNlyIMvpLyb9KAz4+OYoKRX9oVwni+X2Tea8atmFlVPW
jPXC5DqQZcpvvasmlO/RqdxYWKjWvghdZT6RbIxXR33xOw6gTh1W4cliSiOY24Zh
uV4W3L6soYxbP7Rvfr7BV8e83Iyt1s3pVWmv62T1sgGgiHV4rIzLjretSUqQzYTg
9LbrnDIuNC+1KfsSDsFVi38XbOiNmS3zaMolxjvVT4sPzMj6g26zeNf4dX5ZeYsU
Uc9H2Jv4jWp0UpbLRG2OrS7rUXxXSal5NkA2pbQW3v2vwBLFX8Caw8axIlOagHXO
PMaaLhnhBZWjF3UZOSlXn8konMdAaUKoTWgx7pMdELm5Ymr9G5DI0ua+1EBrt+qj
CPcCNDjCnkZhDSJJeVQ5EaY3zo079PdxxYfDlbBGZJ/FG+70xalYUA6nLOUrW/6Y
gKKc4k5/aIX66pqrYnEijCdviWd5mz6jPu2o4BHjX1lqkSl3rbqq8KtyfmArYpkM
kMJM6/4xKQzN1Us0PVObkVsqA+QcFf8mbUGRLBtuZFDMrjRNBuwvN4nDuqcRsy0+
PeyFAj0yhH3pue9TBKryXp3nGljlTg7SSpHTY5lLbO5fYHDyh6wjJKvdBFtI//UV
QfJ0bSogtqDEgdZT11viG+98ywiEnVZ0ErrcI9rkuwyGU4p/sTOVKQ/Om2J1eNIc
HE2iNcE0Xr11OuN3Ki9wZJdiPLNyBzPw4HuCbtf6+IVdDhajfaQsLcdkOebeYvSG
zDi98OvenGzB0XNzSbsuqZQOR0rhYdPnIva3eBUrtf2oK2XwwxkHy5kwc6NlimxS
IpW754Q8ZgcdKT2kJ7D2gJSenQwesJSgcbo1o3YMFA29YuYUyGTmWOPH5ug0qhzs
8w4JRgcMr4ZxmPyIpcJB008GZ1+zH5g2g6WBJALWs2LJJrfnZOtXchMV3t3cHETM
A9KvrjjRbGibhDiwxiV5xujf9qbPW4LHrnmP6CTEvc+r4Zbr62rCbxM7r5iRRFrj
xVgRu/Hlm7EqkS+g/4OUB4L2awXSRvS3buEI8veUWUSerK9DxUEKpS3w27Jk/W3C
b5e118rVzwnxNiTN5NP6h/FLt2hEJLmWV/whuotG+PErUnV1AGkjpo9OljLgvsEV
fbrGNO/MdMer4b1D6CFqxdxvQ5/dNRSQmb7RVMnJWGqUAvz4kly1aM6cKGyXzPuO
8oNmJNu8dVnyavEdr4CKhCbwgz0yvRXFS/ZfOtWsLhLTqtPKQpI6GDbujO1Krj5a
9ZqBxAle+uy09dh00+WEX2WbhcFYbrupVGUGm8AxigIf3JQxqUc4Sx/HGBevztu+
aBfaEfJN8JlFpZlenaUGhn1/ydFPOs1RunhcvKVk0/EjTc0Lo6ia6tATrSaDOVa8
faT5W0qjlofmRgaAo1C63hIH+7ZA9SRiqoahhfLgFNvqB2Ta8LMViVeuqy7iUsHj
XDFeaeF9f7DP6McqdPMg8UmVmrFg9jtmallnsi0YDz++QxlQfBfXFJP2qLtF7K0C
AKgYURnTsB0ukQUipzFxWYDxhX/xPNdG3Uc25YTrou4/X1q0z+q/41+MsO2KEZM8
E720YESrQ5v5pFrqPOWfi5QfUxiVBY/OgiJ841eXs0DyTZ+rh+ORvcId2U2MD+Hu
NYIaf/JXw1SW1xJP92VjZLI7oQeZLvqCpEa6M1bGYwVR0ox89Y+XHufGzRc7WAEg
gGdYd9lTqQ8LKsENrDfqQpnJlavm3QfAc7VR5ltmQd2Rp6xTQxUcmVnjnFzGCb28
vJY7Cvt6izFpXBBM0mz1ecBq3DwDEtC4H5SvBoEXlBh2Z8nvkhThope6vCoaJH9/
8RITRKKCnH91fERCMZkmSgRoetyRoayhpLdWJCV4eQmZvW/iNg6ePH7GVABDGD7b
u0qjQf3y/iND0M9wEddcW0B0jHJWOH7PXs8XIha9Dkvo7ByMIKthkYKTTvlUyH0w
u3woXP9tNskjRiAorGxiHaCU13lDmQ4ELB/JoS7W+fSGfqpPtVfKgs1gujpKQSXP
ssclRiTyCr6VZeM4nV2I7Ik0LV61HEmqKWRORf2eMQgyebL9A5nNx9NlG4wJX21I
9SQCCkIAK8F/WxKa2KXljD+fgfroupw4y4zRwKVYpg0nUMvb0lUrGiFq2DucZccL
ah1LM2P9i/wIRWLyYE0gy2uQSlGyXcM2iAIvQA8OSavoa/mSYF8pT22pnnwmNulR
3LrH6sRGTGHi0vTn40Bv3vgbVPEQ1xJW9OlE+JU+J/h7KjbHy0FdoMoyG2yAU4YP
+9iCotc89IP3/tqVg+UZtCUlyV+zYnIvUOGFTNMJnve1T7t7l7+ChSBj5mDyxwN1
sX1m2N8mUau4doikMfn2Rp/C5Pnx8bwK+IN5ZpoLhOUjTGRH7zRlOCfFT/LhAITj
lQXKn4rsoFwuJZYR5A32efBNzAa5q+x7FBGO1EkxNJJgEwKYyLO/5gG3pOdFnRa7
j0e/hGqDJcIQwiOa0PugrtZif0lvjL1LfuWUNA9FPasrM2YX7o18miiNTqs6hT87
JDj5wMFpDxL21X8u9M9ud8vj31PaBeaSk6oCn9hKdl+nLAr8CCi9pMcRf0IwgU4Z
8GTCQMuqcRleO+urhatr0SNNj1NoauR8piSEF9rv0dWd29SprJ1rDfrxvXNONrxY
irW4WH8EPiF8kMuZ6jrLBirt0RL3Dx63EGwwKmigXnEfFxOxk3a7XWJMeHnmQDlb
TPJPNdHXoDQjsu2qWqcbxaFFQV9mtT+1eQket606ttsVVPN+qcmLkzn7gesfgPyP
v2C+PSkVJ8L6pDNAj5UTjGt2kLplwjZwMmeyKccPCzKiFtXFayxJ8GS4ag2bi2G1
RyXssvaLCbey2KVxYE4R8QJsMxFjhtsCw8m7ED9rRELuP3oM1Z3q/LY9YoZZBGLf
T350vODeBx9D1L6Hf6FFqjtla9r5dqVAfZvtQmmfF0M3eOejdqsJpTZ9xPvwRWP/
LbJY1LqaS+tsBGG0SfGktFJJSSO8+0NMgGtUslfiMklIwF4+4A9Ail/2t1uUI7XV
YJRSFfNcQHt5M1oGgu6Loz8o21flo2s2OksRSB25YOaNYXejhPs5mYFrcL63Zfuv
PN/NfULUbi949+zRAVPmlw+cJSbSN+T2q57sB3kyz8xZciQdVZnebUvwfDmMqDFY
xvXPrhGPfT6QxpYgIcd5s9wNSM/JuFfVnNBZLUsNrBJ8yScehtFKaVadj5QMedV+
BKRUyaCoAqhBAOKUwttKCx0Drbw232gYwBIsOQpoP2ZgPj7VktJywHN2IeTWGSs1
0XvmhEZ586p2PHyynv8/r1dJ0XIp99kWXGvuYdN5DQdhnEzA1PsKECwgOKK/Vzm0
ToNLsdVvYsBziSygouLw/qoewptfDavEY5EXHnnY/Lcm/lusVo7xX+KWp3JHnp8q
gke+/attbv+ijB4IHoLqOuRnwKgOeYIlNVWkAFZDli9jku4pJOaelfFjc7nwENQW
QU4/x2QZHuBRNWByU7nsDlABqw89/ef9Sl75j3dYCdA7SCzxQKP7cyG5AMFtqX4s
WEX1nDVTdLjiEjZL2UhLA8yhZXo6D7pTS98K28ziCLioMpOcgL++Z09jBSmbp5v+
C/pTwgSUoFZJMx6WQ0gON9NmKuBmaqNqGwjMkTFnY0kL1qdhsemK8i0KnLWv/PSI
0kJTo8FmRL3NroaXgPGLBOX+yVB14gksS7krb9KMnrjyJJZwbvmMo15FCEidiS7a
zofTKl8XMfKSgK0vdRfNuDtdVpp5NESW2Kbbkk7+tjKS6vHmoBrKcL48UlO/7K+g
IdBoFkw9UNA64DadGH8m5OYGVugzYKT3V+TP8d+esMrdut9VSYaOES+N6U4TqXqZ
I7XwaWZuNnwEOqx5LT7I0uJdXq8QXCdGRWbDlTQf+ChUQeL+Hv1OT7YgjkjvwK4j
vWLXG3IbPUw0sDFmo1OyCCOzANIqL5WAflPXAqS+BVhIUYtIbRBZidrndzbjmvsm
17ovMpKOkDD2FI7MJRNGleIaU7L8xpo5/CSvazfs5+i6pxotxbIrhl9d3+SRqcdM
37Gfn5NtfAFs50NBUF5+Otwn21m/cCJ+irl0NAtNJftXQpxzBJZuVya454CX6x5g
mMKAX3Qq3vXPIk5/zlSLNh/fQ0o5pRHrGbP9qdSq9/k0I6iu3apxhfHkbOMsNhbm
53fKK309uC5qlg/RoXvGV0CxZ1LhosKTpSHJwNTSUl7Vo1+LEnK/xJoLGhvJPuFe
rtPT1TSeK4Xu0IeYUEDU4fnIBT4mJw96S7ATlFNJNLXZrTxLjtp7qLC9eN1Wk7Ei
7dLq0QvWk+hQFKbdGJcz0ecaEAcVbsSrqIIcy2tGD3V3jRWnufcffHtKbHCiBa+i
P54v0gRA7Xtddg6qwST0J7qIe2Cnd3dfKj6TSfJTqb1ksE43An+YaYeBPY4OedGS
v+jlXchqOlTAYhmoc2dDjKJoRAyRCbUDARHkgNYugPhW3W6/wJOphCqeuQPYG6Mj
XVbKm/RLrDEpUVF4m5Z3NH9FtB9ZQR9ypeT2HqZqAQJS8Z9n49IsV0oo0goAtZjI
qpW9GLB596qjo2bjUDaslXrUxX5dIXBtO2zW8Oyv3iRIeUqcgZpI1nNUqle3KR6P
UGxCBcoEsjnxJEtJLquA6voAbovju3TwGnr9hAdmXEiJfZ0kSxWHiHWg3c+jb2fY
tLys7GEw0Mnxjs0dFA4r/Xg2gNGY2ugsmkYRoVz5a7W45nRLElxT6b/wo9W93G9n
3cLy55KPEmH94h5JG007TYp70YwsH2t7yiKGd6Tcnl68kCbmUSYS2E+BTWJsDVwr
dJaaiN0BUh+Xfyla8Mv66JV6ZEjOxgSQ7R8AWAQZrMlQBFJxs845FTmle+wRWhLL
j8Rc2uNevZQ4fgTlTjXQC58VUThxs4jypSltTl6uRjIZyw1GInFGWVEgNQDzhAIU
xI9ElNHOAKSSefxI9aav4/e5Eu/XodBjdgqKVUmIb0oae8sxJdjz24X3oOxaOLz6
romO8J1jflMNIne5uKnuYJkc5odwcNNOFWh36qhahm94bQR65acXu195IR0OrDKf
43rzfnKUtYDWvLdgEl2yHNSJgwf8jqxt0PXD7VaNgQxHTZCzD471HLSnN4bkET5V
7CaYrLPQ81hk/dBKnufjHPk+o49ti2ZIvd1p7LGwbUyU1FmRWAfDQwvHIoPpmqeu
iBtKVpO3LkjYVzgrCn/KAHqa6gFTc8XYzmZovv1RQZYTkPI1mdGbfKVV+2Ahfyxf
LRtUbw/OLjH2oYamW4+IjvtpUKFyssQO+eAykWXr3DxH/7zjoxK/5+mOkxT36viw
ePXeCwQ90OFoz+tm9NGQ/F438o8fsSdvFqkExagcD20VPAQuqvTtLWjF22SqdE4I
ue3HnH/zvN88LAMz8HSMlj6cFgNahBTu8OxP1S2+BIhPtvhHsF6HHQPjKsZGajsg
J5fRy6eByRRM00qEeAvtIMBiW2yz/VREbMUvQX9J17hC1G3y7F+1vWo4OjTMOM0z
x7CgTgBHels+hZxYhRmvsAvLEL/kNgfT/B9OfJcr5MKCufmpvOWGf8OSTmtX0gUN
RAV3q4yP6g7F/1VssGbSb3tQC2pM7xV1jfFn9S6mtmzTpVG3Q/1L8oekwK8ZhY16
9Vfu0AoU8+EoMQ6XdkDal6X6qC+HFs55IKXXNsHUp2MhlNb2WBsfSzWkWHzUBqQD
llzXZPt4WJkNHKHfWsup9ty62wQt0j5tZSX72wR/TC8zixjtNuIT9qNEYSWpVKQF
Ja5j2kAkILAXMCAqrmXsQHp0siGRbjc9X+uLg9wv3o/itEAjEY9SExjI0FyB66TK
pdSkvipzWemVuymhl6xOURnEQsX2A7vwLcQY2Xkf6Bvr+H9VwogsmZDM2QUq5RYR
QkMRTg1gCY92EKtTzvC0JCCqd8iyJWWqW27BBx2FISc1fcW5CYQ4/L8+vRjakIpj
L1A1sf2ojfPK7EMvl4etq57a2jzbi60o5Yk+N4P8jMzFUVUw4mjmISPS7fmgmohZ
kGsjVtN4CQU86cFR2VBonA1sVhq9169W90bE+L2v5BOC9pRYHNj+QOpe1jqenzUA
d9mcJZLeyyQxFtHRSJWioTTG8miShb231INTVtIbYmk+2YbUJ+QildkwEY/PrKBY
y/aqspy5Sh0BvFPR14QYHjDop4G9rRy8/AIkJEWbUgDNLyNjVdfd3KaXf+PKnEAE
mDTh5CqGghioXHTYmeSGyD68cBgOVmaWLk5mAA9NR/AVWmgu7JVsF6VdxwZjWOuw
oCCleHCwe5B4ActjV/UXoHl4QEj55vWa5zeB6x/i02x8H1fs6mdL0xMvuihYVqq3
Z9kpsLz+rls7Wja7tHGqWzvH9b5kWko6EFRXQbD2IX1o242nwcwLmNKKlMg9qcQ0
xDuJcfYjDrBCx0odr4GpdPSA2LmZ0yt1ZWjsJ+xJ0x0aJ3dOa7R50dc1Syrc+NdR
ukhEzcxCPDW8Ntig3+8ZlIXKZIo+XWoT7cRFKi9U613AMht2ct6kDKHoNwjtlVTc
ATKHR6kvnRVhssr//In9pIlbT3kF64/An69XU2LdI6NqzZu/sj81dIracmAtNYQY
h05KudwV0zGHozxmYz83xTPn+ihzDr2MQp2y/hI+phFuewfRGFvZ9lJ/qTmPA72y
0chGvTYH/pGZVomzxpho6nHHw68qNWNp///ImlAmT+XMeb+vYQb4YXCZb3tQ2pND
49lIZW0J0M8EumXlD3Emljs0LdUx6tXtehtk6HQ5S9NBcXQmUm/39XpRCUw34iMf
RU0yYKPZ6e8b/DA1/n3PS9cJkEXIvQd3+iPwCCL7HnR/wPKzr/d+To3np38DVF4l
e1f038VBLZRd+YQEhzTqd3IuHJyzep3Ntibg7wdSrD8Qgzr+rlgqV0pQrR3xKOgl
UB+PIHkTZTfNjfO5ly+HTOpS6tstsW/6fsYg22i2YgZvJL0P/zE6JnEu9ePvfwcu
7jyENm2ikhgzbceFyvn1zSD8i4Jb8u0ObPA30JVaXaVAtxyZEHY+c0mc5qbzOao9
fQzJUWArxFs50MFectbku1Zcv/Qk2N4OtCRMnO0n6m2KHMBMrnwnS8Pswn5NA65H
sx/hyxTPLVO5zAthpisM7ncBmtt726nLVzWKULEPfDMXiRSbcwtiK+2Ff028gLfV
D32JTHIksDyFc0Nu811tfIe2YjxtMjY7QJMcBieMIsPo+LNtRl8Mn59JOUHJL20E
Q1R+BojlSjRPXwFXl9DXY5wtPDucivNFcWg6eRflejG4BedUgk6f3yMH2kjptCTj
UCs3jvQmdN8kIWAC5aPfVt1DlFUlWyetCTmNUB9miCiahms8X2zw9qvsLjezIuzW
bY2Iv7w6Av03muy95UUJDhbHh+zgqb0W/J8Rluwn1eUxNKRPs78gc/xU2JQD0fIt
d5jXEFKtM4K+jX5uQBFauHYS0uAO5NYuYrFIzQxM/rfV9XVcrPdi5b2hVuSCDV5C
mmZMPj0czBlnPRuksh3Q74U4/I3plOAt5clR63q+0zbkw/i/SUtrYm2JV8L37uWw
c4f1JK39WCEMrc0O/cZjmzgB1iW1mJVmJFo66ALYjrlNikiqvZD1MJteKtGLVVxc
AwZZx3p06PYZ2LwgLrFInvwv46cemxSNDSKVFKltakFTAvj0tdZdyoZf94b2p5P0
sqen2P54VTsw6hogRwDEABftl/+5QJyXWRJSzcz14n4xQ7lhF0Z40iPEfOCl22+D
noV6pOBwSABh2AITW9YXVOy5xtbKuQdW6c3ShPZax6P27RiQ6R9joYZ5zvR4H1uz
H4Oq4x/qOHMG8EAT6OdNEaVQuuO657xJHpr6GmzRTDySPbchpvc71QipWnSAwBGf
AJoo6vnKrxxlWSu3SrweNj1cXDyovq9RU38okmaErQ1+LCVdxB++O3lCeSFOeef5
yu8zNHzomuJH7gBpsUSejRZjx6pJsAsS76coUbGUUhiOZUViJ0Q0i1FdqTMmn0kW
Zr65R0Ee5TlTffBW7uhG/ZdeS6tfpGNdXd4JnceZITSDoZEixkAczmoGPM1jjOkC
IBD/77IhVvTCImckVKbh3QiP5wVnvkAPML1oHpzDCSb9mq7BXXXUTXSSlbtp2l5C
N/VBLbaJka7oFHL3nna+90DJNitobSKXMer62l+dAGHJDYeYhbzThi2vJXX0/1Q/
k4psM2uV5R4b9OlrjN/i/2oDGzSXNzsU20ASAJi65vhfEIBhvX3Al2qj5lq62VLI
9JHgpVTc9OmbuP/ajIaOAcpjWTuiApqM92V8gDHvPiJl7H56bXM/lwWyqjn87BP1
cxvtQTvsm9Ahz8NT8N25Gxuf+mArE1khxIhr09qJn4u1JUb44yQJ0/C9t5U+Umiu
9gq+d/PU68HpoXjOScTMnlUDkVqJR37D1AoyPUYWejmDuJEZN1QveidAl5nuyTSE
0A81DIQWPpla/KTUS2BHxJuZcVkmrVgYHsVVMfShhDbqSPc1OYM+sKORnmEIqmXb
x1ojtfzX2T1phcPB7Ven7087mHFsF54fhVstLrrMFDXcroEr9T/g5R17Sa0vVM69
mJdSwVJOBPE5qSP4M1JXc5ErbrvAwoEv9dRfruz6YbozOJRXWuEDzvTkwu54foIp
yrUwkg1wASOJNmTTl3Jg+O3IKt9gVLGXifMeY1M2dQXYxTplQNRKoVI7YFU+Nbek
usTPeAlrvsAOAqk1BdkW4iTgdZmEZ68Upoc53kkeX9dLhMr83S9339QG0PZDsLDx
BBMZ/UBbOmzL4T5oElg/Sl21UL3LZOzo0k8vCJVDTrFsFOtGBlC+FzxGwDDwSLdy
nPCwyCGDKehNf5OtDIXMYXR47I87BogNLCkElGbVEo8ngYXixobutRlgzdGxrCoj
DTm2PAt7cGlNL2FxZWFjcyHJdC37fVni/SYG7Ydzk/zj4ZVI8xey3WfsO9FKWUeE
dg+MFdSG5hdd7gn3lLbOgb07RXQRcOOa1rHblk1aQXVTmfUZgvCIJfDLMd25+jOZ
cm51ZCFYhNpOcXKw8VbDy0UPapppbcibZAYdHgq1De0JvJQ6AzFOK4mLBm7W6mpS
zJ7AizJsBIm419Z+W8DNytzHRB6cEk7285K5HbW3ApD6JTThqrsVDCnfKxrvAQ+0
h2NQkN2puNE/TMaEN/YToRZje7hZ2OtlQe7edFlwizxhFGjG6inANM8FcUGRF5iG
DsznOPuJLuEE52X9m8d4n5lOFoz4iGY7NU+oN3I10vGxQ4wqShnDjo3JeGbmlkSX
kJcnJ6O1tVvJIj0rS+9YQr8zd/b4UKThR27X57mAmdDyaM6995L8IR1wTiQVn+dA
PFLtL8bpRJP9KKckmPha8bjU9vFGrO0K3dNs6cT50WQ/wyrUx4ACh7xDghiMHi0A
K7KPL04anfyRQrfhoo6czoZDMIafusRY5YGipDWWUPoFHgrUaOwv/oO7SoJ6MBWX
kVG0z/SNXJVDEh3DTXe/m+UYo0S4h8GrSmBmXgiYmRqkXA5v5oR1i5AOOullVkjm
iYnT3kE0j+kA8+zsth5UYZp5eOjMMvKHn67aFx8WKtM41JKHpVErZTzuyxCj2dJn
3av/5DRfR/u/R53wgveby6gyinpJQ4Co6VDVVG2QrYGDYkstVD2VE5FGT7m9avLs
YYkadWJugZgyJiOY3GWGBikANciUvyAogVGrKK961lhduIKdwuDczmAkxPuDaYcZ
obTqwSVlKm6+7mGMasBKmSy5cE5wdalNSMdbYv7jrwGhQCTlKEs4g6n8WuQNNBxp
mVvmpPLDBWkJ4lD7vFl98YMInZz0EilvOQI68In4ZzGm+n+sCGqaXNgNkakgCCXz
zDa2gI/XyzzlRJMkyy/Cc3jX92Hv9h2smVFxVZMaOLOfIKYJd8udx3A3ybA1LD00
4aL5aksE4GAv39qfE4jwG7yJXuY5JD2/0svJaJEM8Y2IJk6yIaTWEbQ47kcq9NFO
+4kQMyeANTT4h7sq5SnBCxdw0NYF9wkiNTND8ifakHjPlilmaWnU58CxvDlxnq7E
1LmLjT1ApKT8ItR9SKHlKoB9uHavmXiOEA7ZflOmI5BXj7Z/kea3876bxSx8/K7y
lGolmw9xbD3z7rM9vr7kGEeJlbr6rA/GvgojfAu+yx0GixE06ZIHSR9Bcflfv+TV
qAhnGbkBC8ATamNtwYicZol9zMORAMVlGOg+H00T2pH8FtM90Ck0g9nFE671sf4q
kHzTe2XUbZQl/GXKUN9bdpYUPahbF/mesvcSCfBikgrcbSsnAgVQ25jG5J2sCXUZ
+VnGeOW9wTg0EJAEKksdp/k5nhRD760CM2jYBYC91FFJSqN1S+vDIlHDcIdZ4DaL
KWftqHyaXGa2eJnbiiKKRwB8kXvPWN6QeU3t+3GB/IqwpqFl/bblgEhAOe1xF+RT
UyZr8gYRiWy/YYMOselCydQtZ3E0i1OTybzTt0NKif3SbvuCf4RJSwQBM86dYb6o
FooVJ5nI6MKeFJGjKD6o4xPodm42C1LvfoZ5G6wSSiwoBj1L6FVK++6le3msNiOk
TtMyWm6wE34Rq/KWqb/pCiCaWBeRvDpqcaO0MW+GBeSfB1z+L852uGyKXvK9Z7vH
JLtgzD57luazIQzndJ+uN2Xc877ia8v3ByCkCJclnBx6QQyeinuhxGbz2x4Gx7GB
VED5akbg4uX2fvewOabKTTaqrBDAuJPNbrG2VjDxkr4v/iUWCbrYYMiIFQ5JnTkX
KacVcCnTOlKDctamcnWHzIL6PottLAx7YtcrKSvlTS8nbMYSelsAovR02FoVWbKc
g1FODFrHkaK7L/oiCwLem0ABPFskgQ7jjTUe9I4QZZUBo20Ist882IuDioDGK3NV
KVNHCGMM9WCF9CwEXjenJMrBtPubPbJvP2RPvCaMZev6C3tYrLjd23xB5aDVf2/O
Re2p/WsgAlCP49Mm4VGY2BST+aGdD7T/xveBYJTvcAzpmPuQ9pwv0DY1oH2ceiOj
ok5DxiWGVaCWBjMi/aRNA90rmYKZ0BNcXKrJvv21jjAk1NjeroSPSqEQ0g1c09tB
25v5y/JSnXtCAvVPnGIrnpgk1aEamhMrvKfAexD3WWdpNnBDRhCCr/UVPEOgtgb/
9CIqPIjBuu0LseQoEx+DXi+BtYb3MfjSUlnSPezyZhOjr9tAJlbq8YHWmmJDS19P
KIdOqgmJGlSR9LEuH2DpLy2EvMhTp0qnJntkcIRNtAbnSu6ZzeB6esmIGBufv6v4
3mhDKQSl55+FBQrbpWEJkOMim3rHvWlaGEuRDrqwmNsf3EIqXWXKeIty0sBcuMsq
JQPHOnvTkNIrifznfesBpKDHCw0zLJqSATl74jP7S7Eo4FHBO/fPQs9SbYaNi8EX
sGatIO525/jl89WIuSwAGI9hmcx3I+786SR5CCQy/DQy/sNs0rt9ir0akFBYjFjh
QdJpt1/UBu1D/JWgtBcg3gWxipZqI83yjEWEfhuVWB51oLKFGR3AC0wtoM3tTQMO
69cpHSttfqo3hlnESnPKEtHBfWF1oy6qlBnFGMjg/mzdaIDcmGVeVrMJiXU1lKtF
7FLIugLHwPwUprIZFOEcHyHzDh9ubTb1cxYw5zreBgDqzsP11veE+GMIntijN4FW
JZUSdz2hW5K1uCOK0baw35Y9hpfEID/nxHyakHSaBXtWxVEZmi4gNe1N2RYlxsGP
ue07fdJcNAcFG82KkOA8Ip2BfCgzSXqCDqPM6lGal9hJELquJsuqMPIbwnt/Q44j
fC81/xw1Uy1n0zNQHw0Go7wmhCN3daY1KSB2dVlHKEmcKw2TI3dnkfuVLCnzbJAc
3Uv02B1qB/nHkEZYYxKxUUgO1VYUXDHRox2zcUk+Pl+OWW9iMvY6NKdDs24YbAOE
272cJukcEUvIb8rlHpVmo8JMblIZZ9JoAj5YsnfMjc/m5UTdq6aN6D1+3ET91MAi
mlEKteotV4nwOyH8agBaMLHr20kFUhPNkakXN1qcjeRPkQJFSEjR+OsNCANqn1Ih
c0QcpfnjGPYClyk7l7CDnexejzQ3m61f7Hu/Yf2WAw1XRr6DyZndY1XuyxuDDH+O
TzvAgfvvWIJTt10Zl5O5sVL8nZyeNsLIb7Tx1x6Pg+XxuHM5HXW3knmLBnnIQKXw
DvwduyjO2tvvdOv1YqdSg4rnV6wXK7MImU0Il+LfFXIXzzWu7YTfSOcK1y7Okcdd
hVK8BwTxZH5xow45ZE87MFocsmn3bTAHRbcPE47ojTEtjBklvIeuZUixmgBCWCAP
vSIT0MLVrP8udzUfjYmxrCeDbitH5GQyixICEofOgGcFULqM6b09aECQ7Xc7UBuQ
8xDAkZth6FcNRbC7YnQXAI7cpuVNXPmTyKvGBSnZrhlXl5pyS1k+2ORevYeDNqlj
ruK10tJH4awwSdEmXurBy2s5mrTWzb4uTNI09cYBnsMTc20Tmzkxqg9MgZ74dgQ0
s4EXKwvBGslOfPsnhV2dmYLYUoNSJXYnrD1IkiR9MBMQPPmy0XbXA7Sir8adV90v
Vm/kPMxWNfKXgZAFTrQBSVfzbs5XDHsT5Z2cEjZ4JbAJ6C86MUaWlkjBPtjLr+Xa
bZLuxg3tcquonVU7A0H0hQq9cQL7NoZL+Mnp9SLIYO2GDbAEzOqfX7g9KCBWYLMZ
BWirt0EOWIyUM5UeOkFKCcyrvVX2sLW4aCA1KZ1tOcDv4Mu4K487PhY8CNuTz3RK
5yk+78PKsoRIzAvjv7vkv9NPTtUDMo2icC9hA/ggpvd6y1VxZ23qs3rUgVBaMl2+
ytuypIBBzvt0wDiS8j5X8noQ7ya41qy1rUUx7s72BlA4slzvPbYdlOF6w061WM43
g2THLGouteQ8Uk2jJH/l6OiGvMcbiuwS9C7ddcKHy48cCrWABla1Vf60KsGffSDV
SByTsID67BUU2PuMzIMKufT6YLQtCW1Rg52zjXBxvozSUkK3EhZMszqQWhuxJVfS
vOyVNI2q6gYoqzWXoyaaVRvpEm0TwOIfTp3eNmQs2lanr4LHhfa9M7NnNmqbEHX/
SSia0asEcIOk4baUub8Ddy3NCJ2TB10OcNGpkg3yQ3hQl9x48ebUvuxPM6wdKnve
GeeSLC+kdMWt40eCy8cukx/CW9vfQMDCOi0bbX9H8yXhR7wEVN2zXk4RxF7YVoxD
oymzbbadYHnh0e7xJYQ4vGjmmKpLp/yJKCc4jQ0bqiuVfGhVIldMU+9smqHGn491
vQn0cGpWRKJmJ3dO8F1WYSSQsElgfC7pMdVPS8vuA74nWHzgXWEu9jbxXGR8iUgQ
SzBOJR6LVLGEW4Zu89WywQ33hjgHX7A/kMfi7gCbsVOgfLQzW4J5YkPPwQUWxkxx
uQeGn8S/Ml02p9k42vCNpOiCFadtQczSowGpMGZkfYa94M+5Qdb1pXe+jynv5Db3
Khxwrub3KpooQi6NUct5Ap2EJmfOqM6XTCypI/mPZNzI12f4O+WTe5lfArvqYC1Q
ZpOVi5HE17BI67YiW98Jrt7En8qtwEYm5lCtcUf3ZARgvx0EzR3zPhrniWzDq1Hd
2FI08y8XvRNG5lK1FDeLhykZK65qbLecp73aV0S5rjZzFehIkuNScMRvGq4aLyPC
TWhQfFVHX3R7hgHVY6emr/YzenvyHdBlla7e3dI0vQtN0T1dIrZl9ZRGFDhHjnzR
HyEmQKyKVZsBxT9AJiHtEuwDtcOZZks77mfYz7oi0C85M+85WrO+2hFrr06j/xV1
iaCESZmozVKgHtTxliu6S+KZXY3sGe3uppbaOel5dblHF4kViCs6ag8y436+Y7Dt
4y7ziUdHgI0UKVce833UjXu+GFEk2j7YHeL1f7hWyldtXKwiup/Q3iKNg1qn8R3k
3tRZFItLPR35ae6xhsydnizbHMhdAFrZwtu/d9Ou88H/6FbHyRA/mGaoO0H0yOga
qA+pUfEO6k88pXiQWlSRkWAcjmYv9Dk7VtfgZEJkeOZnG1R7NOD89KlZQTL9e8HN
Du9jIYe2YyBmxfXoZ9gFsJlBmR1Lo/oYGQ0FgNaoM1NOytnZOhKsT1AzVkzVGPMh
Nxc/cd43qv7YuGROOetyHHqSrye2qNaLrjZLUXml84HZCogwsQj4I11lWQMe/rR1
HbrQGdly5Df1ta5f9/WHpf7Xt8rPLzHvvdblibSAYzdWYnpEpbGEt5Xxbqfvw6nY
fK2TxRskO/sno+H4RRm6D+lLk3awRXzN3PZWegYd9VPYN4OBl7EzSv1I9INXsiiz
2k6DlUDNDKUFc3TDyS+sXHBz2UqZJQ0CsVIq6uPGXY/sT8Iqm2sFcjjpIfmj88AX
FXPlIap0TptKouHAglPOmmyo0nu02YQAYjtM5Qz4hCtkIX+6Gdfo9xJeQo3TzDk7
vzEWKWqp8rkcHvYNgIOXIw5jfd31vZ7OCqvcBqp6YFUkFWQX16vHFXLtnBSR1Jf3
ARYGElWh0GDNcnHxW1ub2p4kntWhNS/45uX25Gx4EjL2Cj7DX6TW2ne2kcOdQDSt
abM+jA/7jtTA0S4EiJGEDOIb233IwfdGpC4/ttLe+ZDOwU/ObF7T+Mrvto8SVo7X
EFPTPz0LBvNMvA0kF1n/C1N64ZKMpN4zJWU7Cnu/rvrofxv6Ylsc7DMPnipn7Cv6
6W30p/+Nz4KTqCw5lgdqkrz1oOc3c8Kv4DzicFj6K6hdv9eX+ry+5ebd9eyvs3+T
tqVcEfDdUKifjBCvOMmRDpBMc2bezu6mDSTV13OmOx2ikeX6sWMVOHkTUuQpFULd
nTARiNc69IbRg+1f4gxK9pUmESb7fvXPehHZ+f2DHePHP0aOJMu89dHX7UtnoY9g
a3Kv9HZa8uzlm13CeqmygLiKXjiBtxrBqobY+jhnKUqIOCNaMMiCTsKQStSNrxaC
VDI6lmFXjucVO0KFlTg0heSG9HD1g8hVFMEDrpxgzJtuvkjsTOKnPLnwrQn9ip27
0798kc1fhQZt8GwbAPREdrfuGY9mwANFTz7tH//pl3xUK9C/01dSsG2HpIYAc+dd
Y86weUI87M8Lx35VG5w+Q2QTuzX/GBifWN2xx8tYfBdV6H1+9StZXeZKWunhRneB
+AW7n/cu1s7grdDFQGjaPKt42sjM0SojyV1D0JNp+7QxkBzQ0W6C9z3Wvxih3Tya
ol6tFfSwfazDF/iMqf28t3LBCEgdQyN/l1dTbEoCNaa5VFScydSYNwnhcnBCy/Sz
1lHEhfTg9WXCWkOnK3iE97PHhcwmUjf7uDOMPwzbJKt+U+pB/I44f8QAnPW3pdA2
uxbPT1EQhPDwiJbCx0GCOxBQXUOpAX90b0pP3ahYYgnx1AiEkcM4VYNqEUx40GEi
94/rDrR30qz+jSNDrNL41z3He3e4yueZQ/1GhiE1SvJUT0ODpS6oC+71N7S39XJF
DuO6pUGY0e1CMLd6Bco9LOnnZJ2qdnfygwB+h2RVG3JFqj2sUYlVtzMiYSJ8Mj4x
ash9CxCzpp69/cnZFpdUy4k/QL7/Z/sU+I8deQsItI81Cg+tcP7s/ze2+v3l6Hcm
hwl3Rgs09eR7RWhrTWRFgimmCD0Lh8v+CxoS6MkQTtgEbpvMsYvReiSbY4t98V76
UuWGRjwCq7ihmkJNCPRtFT704usr0aeTN5bqGCKcelB4T+3ut5g4qbmBa40+pIi9
ToBREc96qCDRzp8DXn7XqQievPehSfIBf/jJgdUJ0TE89d9oXc1oJyDbIXmiXiGe
o/J7Sni1SRr1AReIibUlpNyzAbPIIdN02iiUyxcGwXaBcDoHe9uOBfevyT0cii0w
37v/Y7XFY7Vfbcsq5t95wEvPl6EB9Bl+w5TkOo1bGiZssIGx/b+orcF9jprs4rNC
6eeoK9M/kvWy9rU8yXB9kVpicxEYjxL5zCjv/8JLXLtXRSYLLcEmbmXxczqY1SBF
qa5FnwScVP8kdM8BtODFAP5ULiIzux7GwABr+ClTIQ6jUxRlPVFxBKjub4W2MdCe
NbEGushRN5IaWkymUpPsmpkpmfvEkTicK3XqiDCOVOVztJp4pPotOE9P9YmDridr
RX16J9yM+C6nxS8gjugwYTTqyYKYrs3E+etliEFOdiBFJSAtzrVbZeSwwumYSciE
PuOlc0MQHA4vjnlBmlRGF8EvgCec3ljOWO03m5HUIFgkcjzqjZN0Y//nVn6zmrmF
49hsyCCKLs3TOkl/b5R4LQibvdZEdgdns+Fa+iwqbmo/TvMkxWzOtDsoJJin+hl7
YnIoqL0aTXqamU+YVWjYZHX55Y9ortB59tXU3e5uTK4AlC3XaVPC+qLDfvzfJH5m
zMeJkgqakw+5IR96fnZbabtP8abJ+GKDDC1KxUjdjdaGp82jCwXaN95F92umLRN+
oE9lX61nm6BBTorWi1vqshG6xquL+vVB3phdamRxISA9O189xkFN97DaU2htn1ut
vTDbmVybaWX4iIlO7CxBR13AN6Xqpvmu4uoQ5JqQ6tZIRyupR8NB6Fqp4J6WKSDf
m6+QmhchrtO24+Z/0mTBXoB0RgxwXGoX5S1B7LjPCPcC3YMhgmKkwIwMAvgLEXiK
GIxy7wBee6KBNyPBM3pm+OyiECylSBw4GQUdIWlqzLmxQTZD9L4TLkJCc1AzZdzN
jSerUHiww/wMv4DF+npI1xSHp1QP98zXryx+gGrCscyU5IRSeVI4gJp5lS6lvKFG
LmqaHpW/LK4ZevmNgM3O6Wq/PyMtUeRnVl42+H/9Nf82qMRzWwMz+RF1nSkdccQ1
fzv+zrFCgYRjTIZv0kiC5rHm42E/UGa1IiPKikmWsFYe/i7ONAaJJFWbFd/fZcAH
jl3s/hOnE1Z6hWqTUi39agZ+wrVfnYEGguxHg25zND8f4GXwgp+HKLL+D0fXmGaX
VbxLuxIs1Bgfqgw2+ZaVbpZCZQh5t81XVxTGGY6sAnmHHuzCrFnE/8nPgc7gQGTA
GNZYolSFJxYjCmYYC4yZNksXz5gCEPf/R8PIp4hGix/mZUFz/iBv6clMLUeSU1KT
mH8+qrLcmmrzzNO+4bvSY3B5dEZgLGIBlFyRgKzxhmtX5FZR5ceeN1qcBSFs60K6
m6HScAtt3PhMzhXsg5NQPJs7J1vSS9215dmORuxr7rTQjvroHqr2HPntNHwhlTt+
zn4lt0UlS4RevUup9mmt7M3z6lg+6h+dBixTNFi3zOa62Fg9OrKkvvaS1kskdsv/
GMrXWC0h50UTQDF5yWgrErYX4AfZgYF51z4N5tDXfXoMipusJqnBe+AvyxfsSXAK
s6cenTSyFbt0oREJkNLqaI0R3ikeqmT9L23J/iMWc+MdawzCNnn6gjOCv0VgiYln
T2CT9A0Fblt0ozAOIxP0WwazOUh6YVJt8TaOy4InugHQmC0XPjBERHS5NOjd7mY6
bKCpHuiBIf0APEXiywLfPVFncLAN1uvCgopO/fv0KhowHsfh2JouBM8sqkjpzrD+
GyhVom80AgsZOcQ7rWjpO3V0zYu5aH+TlQKKwtJNmhW/JZAebx5eSUw/fQtM301I
5enUZupuFtId2GSvusFIFwxSrbqtrFhI2n3S5HSHO+11IiDJL7jLXsN5fNmWASd6
5+cCzF+aHa3CtySDiP+PHKGdF4PVCk2LPrsUXvW7PW5c4xOVTYx59FK7pz4rj0yA
fIzS37Y92lVPRKzP9N3MMVwzPcLSBFXlGX2/0D0bzu8inyMgwoAcRt0Fi+zW8wUE
1/c5l+jT6GF9MU25bUAtgIKTrBkPGrCmL+gDwkDaupdsWHzDtDU7Ou6IdOtZboIj
ID16ZKBhYtTWzjE8atYOaszOtYVQunylDJMB1IoN7K58L6k43VYgsuZj3lqjMypO
IJBu7q7kTIm5SyymRFcXdrvWqA5D1+MSYUjkbGwM48Yy6bVpeQTCjcL6mMYImMSd
pUtYSIT0Z7RSX72dGHUyqDl95eq33VE6J7sCZpkyPFaw6dQ9mTA95IXnVxEZH7kz
3DO8mFSHJCxDHQGswps5Dkg9QqH6fJExcKKaoM8dDdk2kmCDdG1kJ8f6EqcLXRJQ
DiHgLjBB/UVq+Klou3MATg0azD/BSyWCaZSNqM0hzciqzpPlRd1Hbc8yhbo5ScL0
FauFOuXYGg24XhavU+elDl4c8HNVTnRfli4GrIMqJeNGAaQSTGSveHe4e+s6Pg/I
AhQE3ssJ6HbUlD39fygGTSfozGXVzIMOYO03ngvnoaD1AIx+PUfD4mcjNv7o5mqq
olcg5W1/YMNFOXeYMaMf0tVwHod4Pf3hjl/5XsaQeND7DsVutXX++NsFCbhXt+kt
4+/Dl0BsOCNJxUEUi/h5Ry718jQ8Nck8eibTh9KDs6I7i3IQD6oQHyCPnnzBxPXn
6YhziKlKSzuWxGRnd5MXb9ZylfDUiLQHZpoCxDavZNY7/HpeQgrM7SpD8FNEjaQG
OAkCyLhoAGcTrMWugidX0EpKRC/Q68UIElfjvwH37wHEJm703WmmGm012daKbRzk
deM1l84ukIBZHziV4/3wiQRxVWzbfCwKAxZNYROR+hGgM7U9GfLz1n+lH5wWA+rJ
6JKX6lnHzHtN0uWMywEo4hKFekcIIwBvrCW+12CTrW1zp/3me9mcbGBrhB5EvdfH
FBcx4GqByneZDTd7BWH/UZkKqJDq+blJ5SJAg0eO0ApV4G9dmzuv2gVUi4DJdcqq
DKKf7uC9qjafyg6upNI9elQIFr3MnGS6IISiRXqCU41fHyUiDmqrAZyzPRzUim5C
IUfNjWnJN1CjyQXIDv4nRh7/JgtnyF4JPTOWF4SoIahZynXlUkPszeYPksgm/TyT
G+fmS8ADKxlckw4dvspMKctSQS34cHHrSY90NnKp6pINzfxmNxG/FJ90Z0FZVDLR
GPn1RTwP+/WCqLJrNUIM/f7csOeS+yy83w6aXb1PH22WwYyKmblOZ6kkfuWaN9t6
oaLuihIdnzsKLUZG0wQi0CFqgQ36pNa/ZphZ7E2/vHyToF7u2pNJi1L7NTxHd6UW
ErP1lMnPkwBFgWk4O6UsSc4mwZEOzDVvCnZ3ZdoeSc/32zzuXv/FEY5PM4LHeDo4
UJN+UN+e5EJx5K7DQSv5ScWSI69ERTkUXOFRIQ29gE5+UYS06lDrKX8VmigwxYIg
gK6epYcVzzy1pOIiZFaJRd8rQ96kv649wlqCKz2wkYxj7Q+tV1lST5SZGVoDRnMh
PH/PaKIwLqPXx4FAk/NL40m9p1CwAdovsWZuvfAaj8eglEbCI452IHvPUwkbq5rb
R+PENXUKAGXXHS1QnlPCWYednWISB32Um/pj6CnLkt0yOsautKGpj+4xfMQrzJeK
rqpKjoheWS6zNfnFnL/ALcK6ZGDsa28kCdByeItmx29c0rnY9m5nw7I6JiP3t7/L
ZkCvLBVxs5jgSTpSXU99Y6LS/pK97tL10mFa1lLyuvOLHVA+R9Adbv8jVaLKTiYr
k2BeFlbf98R190bLntSnsIefmGJLCYAFT6trTTFZA2vkenEYMigkMKZZ5+XMiA7C
nDndhOzv51ie5Qhg2ooUyIkPlSsOL41URUKChgly5W5Ifuadhq2ukHE7vctWxwg3
pOr2ieaHSDVeKLmKTTGAkLLagIMBtx2rHcc5Pcc0lRhcAqPSmX/P0CbUug2UR8bz
k5Y8jPaY03F2wI34I2Vlwj3vZxLj5fJ73nyeKHJpJSlrasrdyLQ3fQ8jG3HjRsYv
Du6cPTkZ/0nFvmQZvyqJKWCWe4QXoP8fQgKTOUsYdGgc7OVLRPeEoZL61CJZeViZ
9iVJu3dbhg2IRUb1vlAb0Y9EFGfTukWfh0ixhjcTEevrby5zGFFoDkSI1BtWbQEu
Ve64N2LLEljFCNniT7IAzuMW8xFkC3caP0Bqcdo2MKkhZ9w7EkJj4mm52bFtdma9
8mrYcIrFg2RI3HfCLZ4JkiWlPaBXCbhd74vWjQ+BSGRpl6hZJD4CFueJQrxN4/qh
85DH40jCTzBSp2a/Gw6OX6x5NMORk/F+JPQO/LLuHT+yCfBGTd8GlL10s/D3zTFr
HQNVZ476aCTKvXfcAZJCltWZ98NR7cCateqpfEge1JOomFx+dxjbVG04ZReE2aeM
WJGJ83yAHQdhQhgnebn5+Sh0QogGHTfudmfb9Cmc9QRFytBIRhJIA+4F9nlRhBcM
lAVoEP9StWFgw9rTlS8IBWAeWeSXqCrzLRhFBYmJFROzrpaYknBVza85seHWrVqj
L/mwT8RRKhyrVooyMxNAPTuyHSl9sOs3WAExQqimxNo7OPqIOnAapGxVyM+MuLWY
pvVwIqmJ/3Via8p4qVGAixw6aMhcEaSuqPpyAtAEie5V93jZscbBZ/M/fNY5Sy1d
OzVo13Xr4K/BtJ061DghzJ8gM/VaxVQCRsLZBhvgxEo1YVJydV/PSQVFJROJAM/8
DAgFccIENifMT1HMmxy5SX8n/VJzEdZLPE5DA2qSXPXlJ1J7PBydeHuJYpYgdNjV
qbkmMqVfFdSkCWt+BS8zehEOT33f+hCapCaNGKF/ldKy7yj0Iepko8xz+czaiR1Y
VjHA0YzAN8wt055MN7L35Wfi3PZKBrAX/hy2dr3hgYddhErWWZpLGr7ntMNFDGUI
qBzWSX1slmzL4CmsmGhjttIlI5DO2/052hIR+7kHeYU+SK4hXTybWJBpdHhKNWTu
z6pfMsFfUYPY/IZNYFLqGZaEfwhZYIArcl/jNK8xO2fRZz9uBEU2zicnnE5pYYTn
4xdjYgbmo9No6iy+aN3c8FRVKC8T/wWLC/vrOYRrz3tGMPssruOEaG2aUIHzhpyT
LUvDy7del3E35SR0eT2P2tQpQCNogMOQ/2G0vb/24zZBvO4JkxPbreLQdWz9D1XK
HVRRT1ep3L8Za42AL1EDuXcXHkRtOsudb0Lg/DB7PkWbM0R3CtJ+FEMKCM5eLIRa
5cYTieLUCO5Ym5ZgXeqqkf9pAAuv+uyQY99l5QRH7fwAs/NyvSMY+cn7Eq2L09MU
N7Jao35EvJlqeVXjwnQcDSTMb+h09MG8ER1sf03uvWk66uge0iGF6EjaqwWcc89Q
ts8mLyhroAwLwtpWXbydJK3vpvocOaL95wo84bMos3N6QYaSLShyL/IwCIRv691d
JpK4j2fFKCHipXRz0Tk5kUFys+illdq7gT606QGtbcetp6yenD3i/YwRxS0oGlUi
cSryNB5K67LHV8aWi+hkJF44882wpHsRdfa9rVMwQex8uYl6GJEkonBkn6zy2b3U
sjKN+Fbe+gkXPApAI1FvmCyzUw6VY+I3W19kkWMsQAhfd4UmuxLLQrPwOEbrHDqo
4Rxjn81mhqHfWUiT6HGOanrokWxXxxX9d1/+3vDea46JkIlwJd7+SkuVyP+pk1aB
Tv53+l6hdGT/UMM4INSpTDPMq8o2yYTd9ht6HAEp8F9LTMv02J9DGTNKeG4WXOj4
zgkBdMPB4mzZPuHiaBhVGz4VKWMiaAhbrHRikl9NGUh2vmPq6qVv8WVbSS/0wv4Y
MynSa04q22gITHuRNNmMG+ckrFJUtf076GGpsFgb+Zrt2teS/lak1QzvUbHNQema
G2NtiE6PS+h+C+11tNozMOAbkHW6uDI4G+p7fUurqFB58HC9O23AnAkrc+QjLCbG
flwwUYyEMefWGNLPg4eF6zh2UTXcRie5IF/sHpgtjbv+eOcwqJiR95+gMRDsxC1w
f2PTKXNi2FXP8P5Uef6ceNs1zsOlec6VEk8zssWj9n5r7/sZXbl7Ku6z+ogIJelU
VVn1lVBqtHWBEqMjqzvx9qTmZfrW3SKvK4RqWz1g2+fa6N/sY2QkwT8Xnam5/hUE
1oIkNEuTRYKpwRp9paea8jkwOCZmAGQTOvf1GSB5peohafZU7KPvdD3wkpdiSxXr
IE300ownDaFzKeTgLc5ZXJPCXe1ESpawZgOfen5qo/3aXYOqltehXigSStsvtqER
lCczOmCQp4MYqXahUxcE8FHAOzaZPQiJEyPQkPch40f8NjdmKdlD7yjdTBwNYPa5
Pe4dDx2Xuo/qKOUHW3DXxCd1j9R4tyd3pHO+t1drck1Ximvt9KKflgwcCCBSUMjY
IoeR0leoETnt2OhR+y/6QiKRE1Zz3HvtzLwF3vcd8SCLE7kPcD90hwwGG939jAhs
FKovCoQmZ9k2QdW+MJnPstt+8sv6CLnIuE+PnsMOgJJ4I4zReCvhmMpvz0em02Wo
uEnW95Lws8A3k6xJdkeUbTdudSjDJcbUUYtcH2RzRjnL15nuI6ilneQlF3wbCwYD
76sP8kyQS3IPACIrV0eeKbKYM3BjKfppW+lo+PBoQcpL7CGvg1XAPpIcT6dD7Gnj
vYiYFTgAAbIG13atIJ9rcwQF3fJtoLnxcZDVO/LfdanIfqkriSLkDO/Pc7TsWyKn
EtRwp9t1kqB89virLG3sBLB6/s11PxNSXNNHwruwOi8O3rdpXpUwJCUqD5cpaiQQ
zTjT4M+wLmgqmTJqi1DR+TBHkM+u1YZfTlP7gbTWCeAUZ0lyNOqljXVeB3Px3z6y
HJdlcNTqa5Qjhz7UXYA3HkKpwzK8Gdo/rbWaQum8I9arZJ/w2WWHkXzEUYAnlEcO
iGQBujhhPuGGpWpxaJQTXTq0tar3pqp/7h3eApEhjZnuvoOfGlPpxZKjkS6hol2I
ySU/I3kX+QwnCVjPfTeowBgM+bIEmU9ap1SXjVWuecJ43pizlzwUNj4eqEGQod2x
JI2QiaA9cvo7RHbTCpF2ofWGo2/A4s7MkGJZsCvg3fpBlqGidSUdmuQVj0JJiyn2
SnawVov6eofnihP+dG4+SPqzIPc6FS4Cht6cPtyhcMWEB1jovAX+cA8bMFMee3/4
HyAHCmsZ1UbFsHjEVPtpe+uAPTG2mpBX3ag5Gun6815VH74nS2H99RQnUjxnk9pB
wLyqXbKV8sm7nAsujezC3HxjfKmr2CiBKR1WCkh7HZLFORswWcoTsPt/XQTQSShW
Ye6VWc3HT0BMQ+xppQU0rEUraHGZXqgRKVgfIz64t/1CMgR3PiDKQiUybYeKkn/c
iThziEM9PJbAw2CwlqX/Gnm0AqfFhiLDtbUKSOyzQt1I/qfUrb4/omR0HSDbnEwI
0pzoXD7IyDW0d5iXNJx9SzkVFLYEdjmfkwLFkMBIruXbKDNkZFLEweooE7ZFZGyW
Pf2G/0rj3OzzY5+B9cfvB18xYleZ6vm5uuivjXG+FfiTz82eceLD+ZoLDJ3j1R3h
cPwdg1AJmoWrFgwaCL/AC1HPe2whHpyAZjJoVwEVlwyaEpPVR4pZkZgUe45mN7Lm
lvt0gdrY3Pn3BKAwcqpIG3yqIPeEALXH755KYFkyJTqi7zlf153gS1JJsjSLVnMt
nREQwnBwceFK9VVSJiFrV0rsm2v6kaD6SungIb52NsgbZhAJ60TunTlUW0PM7Ijc
xIKsSvAF+fBj5kHOfsQuI0iLY6YiOj1CEM8rUIyEiX5Kfi8O0KYYkJbVPOEHtvin
MA69oiACPJElvwCuM/5kntTdKH8YIm7upaBTQTwsVSuFtJXpYN/Byb88n++cOR4K
sPRkITNOFBqc83HttV09B4bQtBThwJ751tRsoVNgF5Kq2cWAuv7N+cGMGilSnXW6
X0nfneinEeOIoCQDwfqSDFH3m/beQZ7/yzKnP1JnAsk55S9nieHaaQ7DubVBcdRS
FM62/YT9UE7IIMqUycltqWfFiJTtlt/FpjquhBAu/TsYikH+x0kLTcNdMyV8YuPO
Qnif/uShYv5EgV4o+w+6LVjYlegBhzqKCYqNMDmgKMIoO1oxsTj3EUAV7fKSs57y
qI52MSz3OXFDmqFa+bkNqr2VQwIo1akFxVTHT18PSpHBI7t+R5MXyuUUEgvAbZyS
bHvI75x0yphLRZjAG/H/b/1xULaVYyTs7iLAwU+r0XI8u1UkuRpqlisMB3wbaEgI
xr1jB0g/iuQpqMKHrAmX9VbHLIUpOk6Veo5wRQLLWCqiUrI9sWmhVkSvb2xcSXqv
3fQ31i1jdP6MrbuDWcQi+aRnVA7X7nVdF12sZHm0f0TNuj7/6LdwBX4TeCGO0uMf
gUgF7iYvALKgEBpCq455/RUjZnURCZQIV8Me84MizSGO9vXdOZcxI4Lkp+tepT2g
jzyHRej9I3HF3Eb80XI6bxk/WPMkukBCTwv5tV8AwxLv1fDV/isyieBKdQ1L31vG
8jMxd0eQ1BhnXJWWVbeQNjc8hGrw8TWE9joRLSSPmxFZrRI8i6qbH0ORzA34WJqP
jrKYW6HO8Iboxolz76beQuJvtLV8wGcFw/uO2UfddL+7fsrCxyCDbQN0t2EWPtWj
C84hq0PDW67kku1lFO085RUQJgwYO8Mx5V4PLNdpwMrNqACSPs+XvkyY9bLQbCF/
PZQLgX/hr0ptYX2940XOk5NTGzqFEMFygAQqW+A9ceEPj5kLcJ3Ho70xUTd3NfHi
IoUKCtnU4VXVQtjUqnEhxZE4TSd+TOQc7eVvwdmj7f6Z8kAWa8ApRr2v+MPGq10g
ytgea1VN2TGllWsMihK4zfluw2xnmwtqGJpZYzQcOKS6SDE51t3pOEydlIVy61cC
c6lZxq1CqDcOg4n8JmQkXlP0shjRvwIEGirk3ofKcTQf8VL5YHpWYSO8w6BfpsMb
bFT/Xcebs0ofno+trOME0sIV9jQakNyPV8wnNqb1fr1v1CGb+Nbuhcmhn9fg9WlZ
LGU2EMBdeVUfyoWzr+G0rIzJHj6HWXyny2fHD1rQXYYlDY2GzoZcUqmSGFRzL3ZK
7IThz2cJ6Layi/69+qCaTxcnMNfDS5G45Egf6aXUXVHyQsVb70F9U6B8V6MST1zA
F4Z/qnsYs5qrvlVKzdbNkxoxrurp6fz/QMm4cM1HXVbk3NVV5p6ClAKrP7XggnvY
EvG6hz0kMlN7qdbMfu34JD1OWd/Z+qH/2k5BELcHW0C78Mq31r6+UjAVPdGkTL3j
oK6RX3I7zLh/htWom/FnK1/2cu9xQGTI15l+NcFpCXEmbj7mqyDfmn9Ou2MUcI+E
7iH1tFJAcZJC2dYWlCXeeFfa9reF4dfXUqd9dWp2Oc0+VmECJ9bpFWAyM9I/oWUz
YRE5YqRxkG+2wSowJGUpAsBiUM0+x31kE/qVI+ufueMYugn53HQlwB6245/aRk1x
8Aoy3CJrSJHxU25+kFtwOtM3mep2M/TxFw2KnaDseeXP6YpiQobJDIzHUp48iq8k
yoZ91mGUMBC7/ifFtdy/wCV2pNaVCjekalyUoFVJokfb5Kq9SGMlaRF1f7A5OOLy
Aye8FwehTtXvLJ6WID3zkAb2q68oOJ4HBZ12IwiGB3SH7k3vB085me5lR+I5id93
NMtG5HsbBKgMLg17GBZSXLx2ubqMIjuwtVPas2tG1fMuDUExNPP5ATNKYaFBDBx5
LayD6ajjPVUBi1S6FK/3NE0rMFbch+j9ufJ52cKtlQjTulQBzer88KpbYuWoKKbt
8KeYQdIP6pQMQxR1vECOLimo38eUM/asj0cmzfEbyJ8tRHDS4m8u2j1gE+MOurly
5Wzbwniu/zzgtUqnA+OfFQhXUxZqaSzzNpbHO1NiV3cwrqVD+G5IMGfd1FF08zo+
z3cAOjfUGwuNuba33fgZfRAxLGjJTm3ujCZFQEVEoqjHcSO0zKAxx2z8rlmrqay4
W8ZTTfYPSCo8ZZjCHYXbuetpgu+m3doDOXi003POudSgQB+NFRz6rEbdLQxCAN/o
TGyhgp1UiY/rkUDkveBoXGLefG/OqYA4WpHhHYUPCce6Jcvka3uIWv2pqFloXrL/
87AtjPYP3b82Q+aVX8iJIhfzS9f9ShqcM2fVcXy1S2XVDlwxu6oK3o/xlZDVPaFK
xVZQ8oNnH5YU2IddCr+L8c+vhqNieHHx32nJxy1S3uj6VrC2VFTeUghEHt27Fp0I
kTFQUjR5YYPOra6ChiG+PDpUWMGNKafe0F1Aakph0Kp0Quov79uY6/hYAhRaWE20
u9uo/2KnCL5J7v3eteUX2QnWAFdBI0AuRfzfriQAdYnHrQeCkF+TZ3tlIHPE7bSg
hRNbtfJTDswazRrmk3/4e6SVca0bxNuXdB7jizuxsEavZ4r/6N2i495cqDvhcPkr
t0izYp4HyJfg53Jnno7pE11GANjBq7xlB0pTSrf8oq/d8NdmpejwHnseogpJzipe
Z4sfBRVJvhK/hZh47/GKVkbq+DUxDDQzdzPk7oEGjgmATi57Q7VwmKZE1SK48Bbb
iqoG/RKmJvsO1bCu6peFJd6o9HJBh8J1lv3K89A783rIHSylNZ7F6a8862G7MMSB
gxrkWEfqLJB5dAtUR1OxyazSCDA9oWsFfIL4bhTaYxEyZ/2t104iPYEZrU7QjbM4
B9ljU3SxqnMQv1rwS2cBB5RXXdtlF6wp88mGChgZtHoNH3DvcFZ/ikLPqK/TPaMO
QrJ9FeMQsg7pCFcIP4Axw7m6VwXeCRDmV28YA15nbrXSTS/uWWlVPBmE61spvMoU
qNaNRz/1LMFpDq1/YUfys01NaHV2B/NWF21krsFC7syherzeca833gGRNKR88zP7
rbjqMAyftAFz4w8DZl52KTy68/hetXpblDB4LN1B6Yt8ltWeizfdqSybnuTu810V
rog7vfxUN0YpgrQLSmW4ZxsGeP30RNFI3AKtfrHloXsvAKx7px5tFcGWPSkCo1i5
NOKz+UaO3jI2k/2gpd/7omwvVHP1sygRseTdYHUgW0HUmxpo8OX60GVulH5PKXfY
ClT223j3cY11wjOn8aFNTU4rP0f9LlWorERRfFO0lH0KAwRtocUHiMqPImEv2gN4
ArZV0VbXfxzOI9AAnKLyBGs3YB5WP7An+kn4DeipN2Y/USWjYWNXMEM5/Y5Xc8r+
2piveQQqMoAhW35mCjoXByyXoNf5EApTRCrF0hU9PeQ/oKfjGE00D2AwyHCgoy5o
hZ7FdHvgAmBDpmcXLcDoVcEy4aznNCbYomoowSVBvIYl4VFFq92nLzwAH3zsUr+O
qJBFgcmhuzInOrTwNLchZvliKEKSkqHca4DUllL4g+JORTYkg9IcYj35xesxgNLP
vhEEMC7V96M8iApaVW25CKRXOv5vAUncviej4gp5SFeagwjfxWzMME6wKbPZ5jgs
EBuOWah4b+1Hppfr8R3bsME1ZRhgOSL0EKyrqcwNOwHCSiZCgHe+ZleiUj0QMNKF
3wmShGE2kEQoVPiscRMUqH3czwcHzWfygNsU9RGjE6CsBLFTfZJGaIxLVn2IVaOA
tdVbvdtZWBhASTy7xjV6cNFgQjugYp5Uf4ufYfjsLfIvfsqcexuRQ+vaw5/KkuRV
5rMvNA+kDcdFrKK+0gAVqdMfXtHTqOF3MikwReTESyVVFXXKsrWr5fRsM9aPSTNR
R2EjADwVWS1qtHC6PKEow2JwG521ECCyWAZFPiomnhc75b/d7MYHPGJ/oUWQkWZp
YKf62xBr1gla73t/E6znt6N1TJZQgFYk83zeNSnsHZiWmMBxGH3Ka07p2sSnghIX
b9h9dSV9ihRe6vbcsOdyl5x7OIfFDZliMQb0Hs2B0J1y08qowAnT4FTtynUC7KHc
TzxDgYa7V+OudFTLsHXOOrQvmgE+4sBp16eQTD2H4XpONvuNWFx+fNNCJAzhE3ux
jTN+wiiOLu/T/SzJJ9az+mbUjrgNeleB3MKvs6sC3tB2sjzM2CHEiBMgRn86fPnx
sbjPABQPZgCnMzB6Dk+Od/3TaOPxnDm5iUhGl+z3mk6zui+SLoib3upvljzAlQjv
ZbhhUV/miKAzVfmT39q8EVIfB2dRemOnFxbCV6GBiGxr8Z0dUtpOc75YWGKd6bvy
20zHwfMua81R3oNVl3Mxkwv6DusUa/kx9XEnsMQSfsMN0rHpiOg38SaA8ZVyCIFT
cHZWdeozgpmnNVvYT/fE4HAH63VG964P37LRpMKvvvkIg9l+jQy1hMd81GCwBO/S
Lad/JzmPlmZ9AWRak3t7g5mtkMqabXp8TKf6bBmOCTAGHnMsPKDN40Ai268X3QOo
SHgAurqHfbk5Oh5gH8QOGRWq0I9jlzn+M/VLtVnnC+lZbD02J/vRZL9E8LCpn7xM
8d3znvGdBZlHX+luhxa7dNY0fx58mIlq1apIPgA0nlG1YRkDxFdB2Yvy6WN2nNom
7Js/WVxzfOGZE8MZ47hcu4vYtXcXupjo4OGV9MzXY6OpiGWVYXTicgBqoOd4g5g5
HycfVJ8Zqvn3eLjTaJtDIxwiH22J9xotVdDz01iRs6XFD4oMilCUXSf1shuF+HGi
PlfwaDg0yGmq8pob4F4O9P2VNFUpvbtbZcCn/QQVGNZJn2clZFLSmDVR74hx6WZa
THRxD1Huva0IYpdS0RvngDaBUdHVNdI6zfTz8cxlJIl5tIebkDo6d6C+LxbOQx/U
XkcAEwE0zuRvFjjWcWL1G+LNtUFYbthLT+mOzMlqU83Ahp8hSd3g/9ENo6F6bqzd
XxQUCHwtDVHUhz53D60EOV84Vyag64XCGWH21gbAO4B7NzlwZVgYTTKkGatIAcAC
cABGtS5KYfdJn8qkSYBKBQmUL9SRFX8MCp/tT99O2HEt14d8BqiZsZN8A5+aL2kh
XvbNGek1+MQYuT/ZC9nT6P1R4g2yH+BqvMGUHOYmXjjSPQmTnlYYhxuspDy3ISgA
XBhMXGISMj7lFT5K1g9Q7HV1cz57w+bZGm+KIgbQDtSipNsBHwT7siW9Fx8bjPqK
aRLyvuYlw/BOip5pkIi/dfNm6tuSuL7ax6DvWYkmpUYCr/PaPVsgp6IDPT+CUkuJ
XMz0+23+KATUuU2NnTIWFhslbBzp9CsNyowoG3TYWyc2j1310i0BtceHgohnmXIh
JCJhQhXPBtx/WjSQGtfjvtjNFhqQd6Q4xuaFMq87p5Sis/WnfabvVN1QpDO+7uPf
DXogw/7e1ROvUw+mG2o1TyAc0Lrd//A+9AzSggA9df8qqf3A83Oftukhm2qU2gNn
KUcFTFrbCzItD26uJ2YHLIlbYz6e2K8fFIHN94eOeaImjFUnFEZtUOz82MbwCxZs
qqrJJOChGiMkDnr2gNtDOm3kfGlDEm5ylSzD1tIiEkCyEzjEhf3Y6/wzS+RzzwPK
iRzVcTU48zhp1QTB2jOvcoOCal5jgACT7FfrversPlglBInQv4Q1fhaHnl97cTY8
ajX2z0ABPYF6Je/qVB1qEr0YUQ3isPFF5CrRdNYQVB59iYY1Wf6r07ZUIruMZHzg
RrWyhxoPFwShjojTNglFtOJ/gfKZYGAvsA5a4d2482AEs+oOGkGTs+12PFd4/Aqj
IKoxNAwNaPL6lVYxrejp01K9Bxf4XeyPS3bfWNiyEnkJyigKqi5Fcd6YY3eFRc2H
hZxDp0OCzOYfmri5WaKWE3ytWYFGYVSVhnisutQwNfcHnHHxUCM7dDG0HVgZoj9o
DqEdpfnLC6QrAxIAWr0XW4VHpFla4msoZk2lWqI45vhgEYHI2CTxSWurR3Mdhjsh
YZ4AE/VB8+lCTcRp6eZwuFl2RiVEgWXXRlYHAbUCCTG/OtxdROPNiS0nhBtJ6QiT
SBI5t+gYhyhWNQntnCIlQw/2tj8ot2xDeC3z0Nm3sawOT4VwxLdf50ss24jU8u0P
hj2JQyxtgVAGxFUyVqOYmLpcKjmp3eBNTXrVscYx025BnlDaZJjbom9Gn8yg54fR
14nAFPxbuann3unNMpiz0F85oJ4NhaoDbROVTidopCWfaGwzRj4zLA3WHTHuibTF
rv42v/5cTti2DbInOg30NlgkH0x/veHiUFF06qaDMOmv75ZbuvwW34cn4mZhTyyK
Ya+lHKFOuwF7TkzuxDNYF8YP4iDfTrH/42jSv24WE1OxgNIY+a6Xk9jmYRbUViFC
Ase82rJQFhD6zLUrkhYtXRhBYr3ji5K5yCkq83EztR8356ttDUJiRGZf6jp6AJs+
vRXwl+27/+8SH9BXnfd8BL+HchTSCFU5JWSkHcCokXOqx8mrYgf2tbC2vmP5aQUC
z0uo8rSF5q6AyWghHTbIi5FpI3kik12FOU9Bbjzc7+aqC2Qe8lbK1muXSZl2mQjz
nRtKoQ/85JS9mJWjOtgkHMNTr8fMbFlI6sl2zbB2oOc2X3INmoHFWzBvuhBPGHmP
rGIykdaqCMNXWBEZBzbP/NYYNyG9GRjkT7hIbibPfzvXk9j+GqoDUapxFH7zJsvH
eg/WnRLHwXO143gaaMyBn6L+LDvSP38OzxsWBVFlZQn4FRZaxvBdtHx4QR4nfv2w
lUHvmW3gSohYtJ6ufhXnNASosGQBP6VLzgFwwvbgwnb5Sn8fDT4IZHOmZerQ3qs2
i1/szIKyxGFY+PP7ScvdeKlEj4XdiToF0t7W9VdOUxJanACIdu9qWQVdlrmmJvrV
IMjBS6yOeUJ7sriqL9bZR4yKSrIt9AGjwyHRs7WZfAHTJXp+ZoB1rlIWFP5tTpSC
HcogbBptWFGIfFi8NumNTh96/wAl2/78lOM1vgeyl5jLfn3YoUNN4Cc1QkuiArek
BwP0qSMpwFdpd8Z1upKxlLbRRM8shSmyxCFH+6u3wy2QblH3BMysGOkd50bVgtny
YFuVRWU+IjwfnuaVajF5iOBZbjhcgZsmdZTfica6+aIua4VJBAftqWeRJA/uUvTH
6TEReMeB0YA00fIWmglfLSB9kBqP2tWsjQZ6v5hxXq2I8ZMwVb0+xOZJrRXwcEN5
SB3RKSwnsbzaI858sp70F/zt7YDy2iso0jjDDqnEcEVonS3IQV8+EPecqhVJ9AWS
2GzmPCRlCwi2d6EsFZjG0k+KMvvqcJISjOo3+rbph1iNoV0XVizpsqUm+wdM/Eu8
dnq5ofrBYlcOV6W5dOKo5BXKy4BKKE92OZTBuckZS/qge6skwPy8GZVZ4A+BGUiB
ec7AaU1qojmvB0tP8XBwOqSEFe8OUMYbJ4fN0exNptqAI0Y86HCWxkpUeaXO1RZL
3Co+aPMRsYxgpkpjvOEA70Z3ZxzOw6uuzpSVygIoEyO+aYR7DIMNN4aiD6M1tERx
DyYsJEYhcqsOm8ahSaj/fWeNFHzTl8zSSzkizFm2ZNZBSK4//w3xX2AUauqwWqjb
krN4k+dcAO9ICwV98TLovk7sgW5o6ruh+jQZe001m3k6WZTvQJiKbn3kz7iQmh75
qlZCd0hUKSU4H+rNAyD1442XKsjcBRa7MRayC5ZPbEfe15c/8pd+vMUidMu8iV/R
cckIkwjwkeXkACTalOGptyYWbxJ9D3kyysKRNfhlulaIjuSfbjan7OSwLyt2+ksg
Q0ufzTT8W4p2OJcWGKY1addC/JqCGB9etTM9VrWaz+HIQ2rzEsOeTURvBTcR9Sgu
e2nymVTgpycKJDywhpAp73x/LkcsMQOOasm2Fy7WIgMGOoRpXcaSTf0FMDKzOz63
w41+jXWHh9lKcgShHZy9I2T+2nKdbA2xZin1Ysmn5zJPf2hPCixdiKUO4aKFJLOG
Fnhp8EMGupepzTc2iWtGZ0bCip5i+B4IQTDWckpu0IffVPCW58UD3FnxiHES5IBX
HGx0qwTRJ+7EL+6b5u8KQwa6dxMH0sJt+RMmCB9RFk41XtjV/tGIiyM+kMRz+YxA
ElEd6Qr5xzzUAelaSW6/rCgyNFzvgGWjGSOGc2n8VcyOqNENryoE9vdhisxNFBOV
3GQnGj0nWDQ6l+6BgYilws2LQUmWYzG7X5WKmpQv5tOZPR8BMBTfA/Od3wzr6doW
TnN0ZYqAiQFT3lihoZOQG5BRqb7/krQNkv2ngNh5vzUq+ioo5VtUaZMQdSIdkcnr
hpwCFZtxob4b8i3z7ufEAbG4mYZS3syjVeP8wR3y1e9Juqxg3WqRvXpG48+IYapX
qXRa0kEy3NbpmidTUOmeGQBZP04KohrVJtpwkeZrS+lDHhraEpOUCp6nhVV+bOTC
gD/0nfK/NiQSfhGxHcPxmITCCwg91qrTi/Xq/BzxtJJFmUXSI3mrChPSSDWzAsXf
9m6bMsIfxz44e7heYKY4xSSMsr8I6F3wWJBAR5yGTFz6yloQ9Qp5u5wgrpQX/KJR
jyAYfg8ppVARsyMuw2nsKj7go6ZKgZipFr5itOPwgFNvUI+7wWxIBNl5Kwn1b4kc
3ix3bXC/phZzNkAPJQgUhf2eIioQJgzrMA51MC47gNKcrBDFAOS3H5+UFqHja6IH
N4H7oXIl6TEEL0HaiGu2PLe2aunhKX7WDyeygDDX7uaPnwdWP0hMAPn5X49/kCJW
hmSs21yfQfhYRIN3ZV/LCC9FPEz9O8DhDdkD+NHAh4luwecI1PWaFaJspMV2GxsK
D4oTuH766m58OxGW7WQI2wsARv3Gsv8MsqHk3bcSLrcvF8HFYB6DoFHxA2cV6Vki
qNHIGR4itdDiB6VWQP8hXzR0X0DlENVlpbw6P83pGHNXnMZTc1Ze80f5U/UzKTam
dnLb/k+4+2vAw+Q9HHhEBS7gIdbgQp4aWSYn0A63HPvaAsva4ji+b5FY7sR/2/nn
sBcNOc3eiSJHxWlxkOXDM47OPJ6IHIHZAGMuMidtxz+axC+zRc4lDRH3gBIt9B+Z
huulabVcKDkGaq/D5UVcDwSXKDBMF4o32vq4VIn8z1r9n59hLJV+awp0M1jExDea
vOJYoirsqFWoDF6cUKiohynt4w+7DSrtL+mddgLl67YKfRDjGKb4m8NgjkT7rcjE
LmnTMGfu14vaSi5m+N34eur2V7+ESEd9mQGtDWxblDGvroAIChv/hmEe02ZHlyf2
YWgELXGTBUg8dN7uirwkHD7Zjmml+huGeDm3/9h0wiyg6qURrPDcif+/tTC/WVIl
3KjRUN/2waseJg9tGKARZcevDNNNTBDxqYtPs4DH1TGhspmed1DWO7l+VTCQ/nbW
gzmgaeui6G90O33cv8qRYRwWoTI2GPSTPTdctHrZ8l/aJDShTAlYNGThFGY+TVGk
y/l8B9IhTVbgPYihy+/gPAYgWrasaRbjiw9nueccHvi4/5sRMzn9tQ+JRZ8+TKRh
igyewx31u+YsctwfbErty00ZsIA9uebXx79JER14rjNXyD5+3ozHLw1A/w+tbopL
Y6rL9apejWpEcq3rGis3OG5vDw92ztqDD2ZIx47McPiRqrawJNTfj16Y+h4EUxNK
XWGkjHrHFpBCKD6XCllS0ZMgYw8eGtcxxwlrk190KhimpFoAngCVhOf6X4s1lbxR
a+9txb8gHDz6ji3znMmoey5SwR6GjpL72AMiP/tcdflRGmBWZo6MAMqBeqAbnNhp
qRbehMsiZ0b/wLwP35JNO/KegufJ2yPEr3TTZmCrPKcyaRCaYt73PRtGbVrzlBVT
h5Im8LCf/GoLuckeTp7KuVNct515i3PvW3zHaBpU/UzGHjxg84G2igNbw4ZqW+Em
JnkK5qZw3XJjrFVazP+FMwoYiP3TTMENzw1fgH0vqTJjuP6JQ/G0qZ3wpN4Qlu9B
KcPSRYRzR+TVHYsZKhiBf2jZpDKZ1Zum/jsOIFhyUhanWcD4ECCVUZ2eGkPNSjv6
PDjvIPQpvwnyuEDVRdffmelgBUaNDq1Qo+PGZMJoC62KEV86t3MUtfaOR3I55UwI
jMi2pRUwFb3SswkRD/2gSY+4G8wOGvZec8AvtnzUME6T1fCPbTtEj7Ptxdagq/wY
w/xO/CYVVEtQSkkb2dMO6wEzBdoEzXsxHBeSO0UmnPlnGXazKuLC5l8FHMMnoUZx
vRvjNvUUUbo04XX6WlBizioUYWiZxWm9S2GULjAao0R5MeujwJDYWrTHqZMGLdft
JZYq+kwkJ/O4yBoGeapzQuhDggWxC/DMZITFUay2MbFUpgr2UGcedRDAo05FiOsp
Jz1yjiNPWP/zuCkqdMboZxTDhHEJTg77mWE2UUrJz7LeZAAHsUkcogsvAZKLjYFW
sxz3owacyGa6HfVt9X+XC/gZaDnLvyeakNGB73uCxcGAYH2qzcuHldabTFU7ZQ2D
OKZD1IJTbslQQ8bubjodl2EcHFMpe2PlTkkYPK1MzySUpnDuqaHFmi8Tjb87occ4
9ffWf5V1ZxN5ZFuPxzV4G1nWBXnPsfghIR/zK8cuMRAtAf02xPvWAuVCfYTvWxJy
OBkQw9yLZB8IG0oBniBpnvGEFSeltnHasHmhwh7C7Pa+JWHcJrVHE6KwD0DAnQ9/
76MT1p/o9vNyzfondLFc5eBgdYYxnwbCa4vBBveYBNNFfMvCIoozSvxvp+H/0rmH
G4WEjm3UnarZuBTB4IRHvrG4gAg60tWKWMQPNSipPHGG3hTmgcw5P9uX9Xnz3uoq
1MFtdGcSE2gNw6quume/zEKp7D0h5wWjqsfKX0e0Me+v8to8BIK4Z2I97A1CqWhv
wAprWXMGHKaTW4J+4E26oJ9JFNU9V0RPqEYKfCeTedgb1WbnPfcDlw3RvWxKXyEe
2/PnuuchoGdynEasAZII13qkGJ+DObA2McaQs6caGbHT7Sk3Waor7HejPGg9ZCga
0G3tA+Pkj2eYb0TKy6HG7kDpBvxe2zJF+OmQslSt9dPD7ijk0UE1ANr6/Hk0yBmI
famcP+yUklqJYZtU6z9Ab86PRnBqYJ834bWY048NU3y4aBjeqCEoP19oJvDaKG9I
EmQlxf7uCqyzitXqEdY0MoAYTjwRwk36M7OZk6ypzhbk95NWtj1b0P3975dqbhcq
opw1F1Jv8352BeA1V2mNGNtbPx43/b3Lmh2H4g1LoVjTn3+O6GUwNAiUUnbBwx65
W2VJHHv++qhqqNeeYuQuhpkofXZeYq97XbtbQbTqGiyJ0RSzHwW5y7dcvgXVfl4d
88VkSbTAjdcROVHPNPlE2aY2wD/whopffhwlPmRiUFtLTdCXI3fswXjUyaM7ob+G
NqeduOXoptGEfnaX1fouwMBH+AuFzbGTqTevN4KR7Cah4zhLgRlvla6mqweXzYxq
5/PTEkeYsSfBZErmH9plqQLX32vnCqu5ZinxuiJHZr9tWpUI+UjPLsAh/C9NgCMc
QUhKJHQuhlg2ajfyzuR/VUdq0A172oNoA2uRTA6jBP+wnJ775hv/XNTxyPY55Oal
3rRAsvK47JePm3MXLHsbauvmsCWES1tUW9/dJ6j22srTcaFMqH0xWkW302Kk5C1p
di2BDIsIXk8zprkiQGkPLbUiFgxlUk1RqefWmzV73QZ/sWpOePI6c5TCXIsSjohu
9zqUrc9a+NEcYD11r4C3DfOvPhyqWFDKRJNFRqU6utFWXPVH8af3WGqPtOxOU7k1
JjYIv06BL/20s7D7HRl3akUdHCkiVNfXEDZrr6P8+wpnudc3Dz/AAkhJQ7jn6lR+
0xM29NmvtN18lDpyxw1Xza548HvLt40lrW3o4TBqWAKzmQTFphtFTHytkgXrBd4a
DkH0EsdWrTzjNdL270ljUk8YwgqeF4zOyUSzcAFZCeNmdnzmzs8oolv73FFsj/QO
C1RJy7RxKVSApAn608J2NO9jn016wGJ2pbNJe4v0MsgDIfXwB1oljAD/RY44F5PC
Ow8pD2UrBvZJUSIZzQF/QLjAm4H1LWx2zm5ma8RfFTAEdLFq1FnorPV74nu2QDEE
/mWeNTE0lxWB6DEoGl5Fj2lI8EhtsNXXoFlzY+FnhdjG2RJA6N3KuSx74xEim6D7
Fn2V5gUTwZmGs/J1922WR7GT8LWU1ujr5i4PNlzAbw/n9k+MaqmZ+pTTiusUQ0lK
FUdKaO7O6iyAvBrKzuShBmKX9dA5ECeq5SYjBrxDMbYHmoIUEio57YxbSO8J18Cg
sB8sZi94WqJ3I9xMPwpD6oPR/MRqYYdQ3kjVflPiCsNl0c3jkE+jbBrgsr/j6d1z
Tp9l66ZvGy4YFfAJ+fgC0j1YNPbM/aKip4h6VU/o3p7+7GKDyCG6IWnNZMcQPQu8
JBSkx0HOK+cTYzr2r9rLNZdLkxLXe+H0rzymthV/+uoSw8ZmXqf9bEkteEX4F6m3
T6+QrKTtsgJs004XCojlEkAEv1iN34c5enxJGEPeOBOQroMM96YGA7YfbMgtk/gp
mYosf2VAY7Nw4iKDlNFmRCeYs1lvaoF+T93d5Nr/Y4lWKKTXu+34FLEA9EKTAYYg
tFOYgNUf9wGgkJFlsnAbETs8my4ti436h0QQJJF94bpfi6mYzahHZogd7FzEky+c
9zJI6EOz2/79BTyah59HNVlA6kVjPhAUE0xMkLg9NQXnGgK6K6jAJcWqAgtSXgZ0
R3nLxR3EYgG/6TFfYww0RaqUNnYRN5PiJjOhuBGgibX//wA4yPoingDi10ba4bIR
EAht7AroKqLuUbcP+9zOuFqyGH2HW3K0shTQHdrjgVRiRcAZSOe+fg7ac3VnLPk6
KCsu/421VEAUTs7PBSl7ogD5XcUkgES9Lkv7CoGz+e1GB+DsCJvjepZ4m8wSxBbw
zolWdwQKrnSKsbWqdeVyDCdzecn18b9SzjRzPh1G33xIMKvlIVgIe1VVTZa4SSPV
wJBlYGPCMkWdQSOXh/ib6jsEMOauhQL78C/qvwg1tgm3M9Dw079VFpd29iIk8mx9
su7ROVKBILdBxfxWpohmtKQrGwj5TBP+gofdRoTyLrkLtF25ctjCWiXb7B8Z559A
NLClyOoxqPrh3P2n0ltvs6KMeAiG2MOXxkEghog7Hr2bVxK2d+bUxiyFbYJmw/2I
3he52RO5pUssUWNLn0w+RONbekTsBVpEvZxEu8hOR9Fc0TnziTDLKCpRnqqwH5pA
Grwn8Ut4drZmkJZDmmZSD3d5uFTgQYkY6vL5PKco7jSMb/lue9yAOI52w27oCHoc
WmtywmE4wf9Ex+dGeQU88FKIikqBwv0JUJ393QURAuaaIpVr6rKRMhDuVdfFjfS8
SFRYuhpnsYyuS0uOh8+ZbAKCWMBPdte4RxmHlKrStqegS+8coDnH+Ssh8Cq4/k1d
+ryjwdZozgQPGJii4R+pWrMHn6yuc+lD24xWixJowGfg2vkBfspxEXlBlXshykhW
xmR85uw0pcdwpOu9jCE2R3Jj0mtaJFsqo2Hrq6zJ93FeUivmI+pIOPgL6dVUHcLN
OMCJLKq1r9sSVDEL8RoardFt3Nr+i//brV05sXTzVSiNINyJrFoy0u4AMgC4nE1m
NRPfvXA3fwGfx7j3M7rBv6bKmvuy1biO/hLKf7JNbYVeuj41THjuegnH30T2IcjG
A0FUrgXGJOgxqziUvOifiUTn5+pMFe4IQiMbROf+sIrcqoADM+bEi922X3dZlYIC
SfIKQKS1cuD8drrZLykMi4oKkryCFAOElBtW8Bk3KRvWcbbKS1zq9AaKF2BeRf2a
Ra283hx3hYpwal38FNk1SZicVWw/5PabEQZqypUwbXT6/KVY8LSnE7DdAhaYFLhD
m8+vv+wD5tzRvPVi/a2Nkfmj6LLHQEqWUW+bWKxKRhWSLLAoyGxlScOIMGhzOJ4n
OVd/q8KUgjM4OAVSq7VgR2BjvjZLmhxSW6YSp+PistXWmEVKwOYqO4PMOQdIL4hg
ubcCDLUowVcRNzraw35eASLkVNIwIFYMHyVaTCxhA/btVEgaE6BNmR9B1Qvrw/Cb
DVs+L5+MVqTQlBJYUcq3xPAMcUqdo/D6kY77uTIVV17lAwH6WW4aHgToDFGkTpeb
d2cwntz6PGlRhvPyy1jobAVr+sRndWlpWg6MuZgMusSgKfLI24ZdZbt0ehqXdDp+
wsZcVpDzEKkjZRf0mQcySHRGttylKQtOgIUs0ExuPEDARJ7VfcuE54MklpzwLs2X
z3WTv+GrR2aRec/Rbz2xDWtX8oXmRSqqblg/PTgDIE0qvQp7yeESalh7Ju4xo/en
11Er/tewprdiNTrq3RLKkuFuVZEiY99fXWeXe50iqfOeMCp6fTTdfuG+c/K0hmH0
jdmEt7Y38c7U9TTOj21ElFOQ6blMxX7Yo6ZbzBQVWxD+90v7KUHuU7x4HPh50F+8
VZaAtD+KZH58rjt+3lETEDD/kOK+P3PZklzuxCdSJ+3/ImxwC6F/X65Ehl0z8Q32
qVrV1qAvbqHeo/9s6Q4EYX2t6qG74tNzw7dtgiYU5IWQI/i4/yzgshu9SagjLmor
KBRtfConfyIfPUNj8aNf8YuhghCab9UwVcwRC9o+EvfagiE2unHmJdrUn5sEYDTz
OHWvaluFEVl+jdmWwdRXBrTD6/wPF0fppCv8Afp855igNhNDAyai9OboMjaeHIG3
9/2ZvFedRk3HvdyGsXGrz7yATCWqbODgX8xsjZvh2Jg/LCp+2VxJih/FO+7Yndxn
YssFa2oirYr2HQkGfRL7oqO2wMU39EsC2FQBWNgU2XSy3nqP3PXI40o5SI+/+AIQ
R52g1Jm889OeGyF7X9fd0EnCZoTYT3fnidAV1FTXBVhSC45Ds1mywAw2/Trz6px9
exui/jIDzm5/6Amb9g+SV/O53/He57RtAdfSdJZQBhWpe2nEuoYJXIU4bjVKX78q
0Ckj8/HfBEFri33QSJ9UqlaBD/brRWVeVYqSPjCDHeI/Ozej7oOKa0aLpwmRjKRR
E5YqoMZXCw1pYYNeoXkFyuUBb0evjskxzBD16/+EVPLEuGeMa+YBlQsGq6FNyH4M
Wuib1tvtJfpVxC8GhlYHuxSbsXu9gkJ27JR/6VGQYy6ikGFwGbwyQiNbIhHnFoDe
9zQvXkS3xhbVzeC2nmMhVdoYE00nJmrVBBkk4QuSHnJeGjWue27DIyIPORED5XiJ
6MUs+HAv6sW1TZonyXbIrUqnRfO64uOV94cQdwnzD3zQezj5CyEcMsE7asF6SQ9x
3h0yHgajVkDLW8PtBo6wYIwl013Z6GRaCif2Qu7IWZwspILV4z/yGmusAQwrgr5u
yEskrqcFKM3NSCtoxGFqYO2c8dRH9D9Bgi7bAENBGPm2KjBF6MFaL1r2rcXnwjSh
NMBEUUMn3syUVzf9ByRy3TE+dmzvIte13gPi0UEt9GMxlORISdf0C1TUlq6vZ3q4
Xwf9FjqF57nLeTjJ/OdvFwWNYkLPqndeQV+yqBDNNGwREkyql6Po9JCEArmmfjOs
ddJZGieGFChdeR/e5hj4ddtmL4SJxehhZKhfPlZw5nKvFMQ+PUW6d0e9mxGmuCtf
Z5EI9s1VLbNJBLZvaTRNfCegh4RxDzOBakXkf2WJvaveNFka9NC4/WWW7YUe8z4d
Xd94z5hknOhZrd2LJyB/F1EV3GxuYxk50URQxfAulV+Cy5xYFEuUNUA2JuWE34PT
peF+PM9ZfIaWEzArI9rs4VY/+03pd5PW9eEOpsFN3e+ViyXdcdvP0xfsEnzC+ZnA
WX7OtWZord3njP1MyiYFBrxJ4IzMfUbiMjClCEt7dXswg9DCT48h6ZS/AD+4MqVH
aNJEOvWyq2yMOXvo3QHPoyePIysBqt/2fXYit+qRA85c31UOE2Zur7JjPjwnOyEh
+LndU0V0Zn6xGkmXevttvtJ+U0ywyxp45/ek+rJqyXcerd0QGLoLzx40B7YlSsWm
s5a7E/I4a20rYK1ciX7xKuG73iKlKgiKixMy0d7V3O4XZ2mbCvCrEwMFOwoTA32i
XOhetD0jo31kM9mNldH+HBTKOFadiEAE0sW60UXrTKgVxkTNAs0JpqyybHh17Tqt
NKLXkGXgLoKDtx+c+jgqRZmmpb6qC7UQI2DtUUC0vDvjC2Fn8/+1FgLRfDhv5aPB
NyJrMvqnxiF/muifGePTn/bLjTkESk06jtkPAb+R9mUqXzDyXRBcJKvzwr3mh8nR
Tsn1gUTRRN2sHTonLYokCI7Vc0oaxIJ1HNbA/aUX29WbCSEdtwcZtzY43n9I/tpX
wST0CzVXpeJTqPx+RTSpLBeDRX+SIYdgHY40Wy13fKx+IVziK4fC597HJSQUWFjb
MxM6he9YQTgsJdAkPrazA36q3mnBaAC+PmqaOuhUD2Ly9HOFZ3F8lDw2h14Y1lF8
L4eVB770SjBCvL5UMtJhrOlUhgDLwWIuA3vXJQl+CINiWho0h7v8+dEAjkeBreTu
GJ1mbdsDC10TtwMh9rugb9cwglkllA+DwRvpi5tyFWD+I/mKng12FpFyHVPYh+WP
koAd0XZJ9j2uQjss/dArpyzEYgObE2ttQxepdaLQJU7OCZG4IwJ9IUZ7xldGPGNZ
WtdZ94EPfbzCtdj/ONTInjS/Dpl8tpjqsCnmeh9Fb4W+2QqaS6UhO47lfXzjUYj7
Q6gn1Ugpo3Q/OJVNat8Qhbsm9IauPsG9QCX/RH8yxywc9UmZ+EgzDkEhLqS4HHNQ
az24aPwcoIJPjHP4fiy5lcHd7rhmFASv9ZLxI3Ue0FZfTrWAh+0f0T5D+02rLZM5
ka9o2b6fi1UW31ANIBW+oo6hPyI7ll88FUQtFQqBupWTvUYH+FlEvSWgE0kqPrnH
OE189jT1qSkgb1ise6/jHqxVwXZ0rdIH0vDmxOgK2c2mAbhNsBfM1o9pn0RQH0Us
T5hqm8YZ+yjhxejAyLzYJ3ncpF6RG1L0OL7bNxd/9QuRQKqnKFukKSPBb9iE5Mzy
ugOsphM8jCWqlpPFYS95Q+SjFqV/8WEx7kZWX1/g4r9xvDu7/mO9zzjOX5cQ6HwS
Cf88pqmDL2gVLsFUNFarW6R081fxW+dcGbLyluowpVnRp4IqtOn5THrNI31sz1kg
Lh6iXBHphQsiVamYo6FFdl+9aYuLLl7hrYGmPhNkFpG1u9XHLvhdLGT/Lxr/RWZW
uf2ZSF6vPZaJBy3T/hG6OZyA9b/WrRdj1FpdlveZm5A5wh5Dg6Ipf2I8b5JkutWs
hT/zpAvsZ2QDfHP6f4+vfXGpRLFHjK/Bg4CxGltBqWC++oV50zyfc6a7fW1mB0JQ
r9dGbX+qwfmP/BgUUE2O9/V13n37oy6vEEuerbclB6oaf8SNxj5zu4deUvNR0nWf
RfOp8vtZrYXPIkv6p3YtReFZDbTKzt2t+mFALwLHOA5yGA924ylHuRbwZUUArctf
1Bslj40vrkoUu7/OpF+XG2Yxrt7BGnWQn8+qGVluPvv0DfYE7q8AfWseGqMzv0nm
qYtkszO8uiZ6GykqplV6lzWs6sn2K1vuMu1TXP9+wjVnGJJT4+7ZIcf24u47HTV7
WQ99oQ+hSA3p45fzfbC6kOe5mxMd8GWilLh4A7T2Su9LcYSpH6VfTkK1PJu2dAai
ylQ9h480a2Apw+gfKSKzICcCOoDqe0GA64lKWuC2EgSvo9D6tXegEx6X6ZuIJekT
KI1F80PAAjYOLFeM/fxrVOCsT6/7O06fuAxc6ZataI75KQyS7cNTtxhp/PWc8LAw
ug8phQHGRmV/HIZvn3NzlISKN1MK3b8m3LVklOxAWG8Q9A+0m+cD/cnMyKpPJouX
ZK/1bXx+ntdWb9WkJ1BbOFOZyo8h6caQHU0a47YOAJcZEz6z/Br1X4WlhIKCjZew
zjTZmLA//bXwCyfIYqVvMF517Uf/nMVeYL0eE0vpFl1KCB3kHISYnjK3h+/ccrZ/
4L0BB3c7YlDq2Pj7W60cEeGZ4zveTNuuo+q7XE8oc0u+SvbCb/HGp6OfFRmNs8U1
lmwz9U/m8deg7R+ZlEcaVGtmDYlpFu6TAFpAQuosMPzriEMdDvJTTUcUPGDfl6vY
j5KYn0CW5KGYFZmUaMWCNlHOmD0ygRKYAOMcN6EHrCs1iXJBQGuKkTsawSNy6pyM
gLmcdqdiDp2CxeQ0BlV/2CMen01nYYKMQ3U2PjoLmE0LZZGNSXvV/FTtQF+j/EsZ
brQ/tcCqiBZqL18LLSNl9D/HhL2v5/aNbx6AcMRApUoUQ7yE4ZKrHHlmkylokVC+
+wf9JjyZsW7dZc79cdQ2SYL+7S6ZLXIkK4sxO+0EJmqdD5pNBHJQLgp6EnUVGZSa
DjeSTsisBtUMJaExUPsUqoxOBjulOjxnO2aGB+JiVfJMy6VWYQpNG/gf+khk7VOQ
iN084bzmZXh78q+0M9dznpblmtYTMEGX5JaFhi5ZgzZ7Y9AHz4oC15iUgW1xXPRS
2XhWeMsSOjXeahyFpGAnsYwOHFNnBWRXDzf7RMlxJndHSMcMiJxTa+JqZkkOkSzf
XU6mGyrI/C6OtMYH3C1zwLpX0SvJPF4E/pqGdtJ/K7YAepfVNp1QW6IXW/3E/Srr
Q+5AJWQV+eEqwlCublO+C2bhRenl78sFn7O3f37M0nkP/6yqDv2VMKCDW7j0jN8P
tndnF5mvBoc5dIspwb7RThZEjtbSQZh0TAjJ2SFF2qa4tSYbX+4YZWjPtvUOENTa
QNpAOZqhYiNlrzKhTP3hlNtlZF1zNM7E/+uYrYrO00ObbANT/lyqJ8t3JDnVgdAy
qd6KYqTwMHZRYperC8Ry6m94CdrgLL0haN7y4m43omB8POm9nf6PYNr9VNtXhJVT
ynm04CIOmxqS4vuSaAQr+cnkzVHJIhLQI3Gk5AyGuY2du3wddldg973kTcCuDAbj
LDNG3kw00vZ4GbFeT+fjVqhBc4zvR7nWpNZfU0CFztGRpr+ScmZ3hP60N+cJpzj9
btkJY2GP+tCD7Ai3Xwrs+HqL2lqL2/0kZfZ4ukVsX49FC+xH9tZVnnf5RiqHPUgO
WwEbZTu4L/tZnKCeHRDRq8urH4HFaLU6B3L4UDCC3P0bUxkM3NQuJjwMOwQmBTQu
lLoDsiEaZlFi60vmu55Yq3NMMbbkS3koYNMI0UTAM7CaHpRts6bxdwvEP682FoK4
FuDYK59rNFKSm6/+md1fNgkgK88OBCtUlb8syiQWKFqyuTUpQoQdHmL3Pi5fu3t4
4l8BSPlZxxtyZ0XzIA/Jpi/ChWYjKlygrc/XmO7du7y4EmpBn2hJk5ygW8uwjuUJ
5/cy9dV1a3YhGraZwITHt5XPhSoIR6e1pJaovylrlV45iee91wcP2H85xRw7nuCR
jsQuVgQZEX4D4rEIYEePihBdhdhm/iKcg0yjL+mueYY8C2oXDAFiJ4Gh1YoLxCVX
VRvElpfjo3uiwrHpjsjxqiK3zpaOnHXv6I1NSFG1uZrlonUYZVNIqxJsU+7O6DG+
Vh4QCMDswDsHokRZktdpAzfKaxFdg6qBszdT4pGuIpVcumwQe0adGKcfx2RiPFpE
5EF1YDYaqYktRQZIXHpDER5D/DP/SZnA7XVgPPNtAq42qPY7itQsJeD+VxgVFAfP
9pGEj6EknYV/zuxymqQvobhAqILHgdoNqhAeal+F4zZs5khITe6R79CUqCXcCCbm
F/Y86dnGgyxWuMWKr13T1UtykZxSvVwqVz6PeDZiBTv7rLUQHRIhz+suRPSaRRfh
xerKLdRft769vBRFPFyP/czUE2m5JxxLXYFNzkNjELNHneRPcplvPyBCFSgFszvL
lYXOd4dddVMXhoqhERgR9FdJYesFL2qjk1q6XN1EPTe5fu167AH4gznhwWAcvo4O
c7H3sLNX7YpEZAx7XXNWCu5NgygOboTJb6Ew2arTDzUbje30OiT/QH1y7e95jTTU
DFlyGiZnWpZE40pHJWMfXlTvuf0x+IT7nVhd7zjJEkFTM6VC669V4Mw6V29lS0ec
dxQFdl6CzJN2GZi62UGnXqcxLETB3fEnB707OBCRSio43GpfptlT1fTo4PJCVALa
dUvwQ6WxotVQsneEbrG4TLHmhse+rNSZ7QzvdCJidgjmUIm4ppLApcYmQkIjHLb0
O6oWSML+D6RCm/VLTle0cxZv2rigsXxiBp+FLiZWwr5i5xVPkafJNFpFbUSeyEmu
QHWeELTxyfNy/egxS0ZiFbhQ5mmf39k1iV5z+qV3kD5ZHI0U+nH2WpfCEfVfu+1m
ETAJc+jSfEK5W/5pMOBUQWtY1kn4ejIBKP4fJbvrSuIG/7UfzDeuf+0D1vlaCk5o
3to0DtRMyLjEUjKPYZOi9QuERRxJfh6bFuZQjhu/Te0RjdjL4/p53ilEV0nCQPlo
K/UZ2JNRc4IFcpyGySNB4mNccVjWmU6LLaxXAePw0kcmMrqTP4NdKDcbrER6FnRG
/fJ+8DM2YJj7j2uSv/Qv+TFn2XX2EsXKHVk1IA4qtCC+n5VL0QtuzHjKp6bBTfXq
5teLH+wDNv5zSlu4rKN2/TCw55Dw3DWFrtzvROSgnQw1P0/OtNGSBiqlq11U7P2z
cQsJ+1ArONR7F7dTtPGkCyy9MaskZeMrhmn59G/gz6FtwKI+SMI8Y9NcAxGA/vhn
VQu1B4XXQUmvBF3gtt3NmAwyCW9mL1UXrvPRJ1Udv7pEXN/aOuuOnppt/QPp0W89
Nuc8iGzCZhQ/armW7kNqIIpdoeqxcDAQwTOzgJ752pzY+lBJWWX+kV5W4pNsUsdS
lrHCwjwOKesTlLO/YY958yhRytF9nBz9vHhk5zXuR3/TXJNqo1lm9vMQYnBCiI46
vNJp/OM4dWYa2rjzNTFUvLrcCepupS6ZTzLzWZKDZZhkUD73mcR6CwvgyleztdoK
IzhxuDtEWcbLAxlPjr1jXX0F4lLc1005dj9igX4ZNUC37PWL2qP5s/jfNuUClNRG
V+dOQ+90l5uWu5CshuFXfiLTdO9SVlMkz8RI2Enky8hU42e6RphqRuJgLOqrWiTJ
j22nuxSTY14gqIKFD4orJtq3cepdlVK6tIGASBspmAV2gUQDghXHCVYSQYUMSclV
1wZcwc+CbPVmNC1pOdQ1eDYcgyJrR9tMFr+VrixpY1zwhGM3tg58bDNHkYKXg9+k
KmMCedopfquma1S/v2ekWYbwlCy3zwyQlIp0rkEsURFl8DaCiblPi6ulztB5FhlY
TN60Xp0qu/PmKuSDhQ3MfpvBi3ZVRX6RNED6fLC7sz5OYqT7A3djmigGnUG9HVod
mKKdK1E4uJGWLj7BLqoUEoft/Z6mkwIeRcGX0EBEToSRUW+6JZjNwNqFhZIkMsnW
/zVu/umtirXc+EQKVRPHQbtnt3VX1gVwKwz4kHwIoIJp7exJcCzyYOD4ftbrn1R0
BeHf+23TMlA5TtSkni73uL4rgYtl7S49kon2yYD44iBv2k9nFaSszTPsIoaQ1NN4
i2KmQO+5kBJSryb/JfCibTZ7GlGof7CU6xsmvTbVMxBGFWurRMKTQ+5Yk7Rdj/a/
rqoc7RESGmzQKk/U4zdMDulSeTkMNWCj+MNvgfNeMb6Ymdr7Gpu+Iy/Q1fgCqjrZ
pF0wt0aqeK2a7xkLfJ7EWQq1071I5Yazrw1afbRtacuXYCEBP9pe5x1hRfkkUnQN
WmkGeQ6vZukQpDE4b8lwDniM198MafNmPWgTuC5ZmGN1+GaOxIBR2rlrP7I3c62h
qsaz/wpOPZGzPY8aFOjJSMQd/YVqgU7Zg98u3r8qZkv7NFaS2nSi2Qs/imTCAxcv
6Bcwtwn/OXEyFzl4TEeX+znnSAY79aiACkzjqKnMOMIudjSLZGeA24V4tjLdowzH
0YH7WeE5lqapUjMhOXeu+PZXB5fEddxtIVgMdqp/bSy/Nm4XI1osMfq9uEJ/DBsc
84Ed82tBSfCajlE+h8C8kA/46+2uT/v96nkfMYhHNVGfoQBeecnXx6J3E9bjhKyd
Y+il6MD1e3MRZvMexjcfcyDhVBv4KxusP7+0pyROY6YvXT7jq5M6U4vOE3+em+H8
G9kfoKMT/AhXPqDsa/yD2D2VjuQ+kgBli4xnCc+aSHs+8QfYYZgnvpqxTk1FTK4/
GHRyj0LVCv25YG5fCOIEc9jxPobZoNm5WkZBFU5qrunmXBFQ9b9iKpzGq9fPe73I
IMIM7qhyK3nkJwj0J4rkong1uq8k8U50BZQCRi2KY6ix7Xe7bToiZO41Lc3m8xdD
aZQ0NQNBMdIDkMq2gnz4gU2NtG7XlrmXNWASKYq07xtaku65uEW9/2d92LaAOMvR
aPzilK7anxEh6YSYOabZ94KHCRK+Gf444RS1C5P1sQiyraFpRlhsGelW71Te1Cxh
h/lp+rWrK0nI+lswM6nyVt8THKHGpkF4wCgOKqXgsCQffnofhZ9Y0J7whZn9UQ8v
HWeRVTl5DsI+N8ZUQRPTpREclI9NnZ9qoUx3yMH0N726osAxw8OmBTSCtU59Rfnd
nY/dXvDAGfEx681edsqkChxatdJb7I5nRPMorT2jhhC4Cwm1fWYUo8UQlt/cBJEr
Evu+z7TXiPN7dz9JNBqWSymR8/guhNWU8HZGvoMHG9gxFPow24PJ094crkIXIfOc
1CBn9Ufcr9RQNufv7uuEff7vOw87Xf2Z1XrDEfL3QCwrTLy+QJA6zG2iNapH8h55
GHPc+f27eXlaXoC7YoNd0iw5seDhoPMpfhr7N6oJ625P8RmKbDtEUsgGLohYG0Bl
EXqrQnlkVLe/35HxRE778eXBgyf0tFcij2GJ1qbd7lwDoPsJ7Mq1+To5Gh4ouVHE
8CCz4T8PYpwjaFVwEdpEbqAgJh8Oeea+/eKg4Mh0Xj3DBhDfMSivTN2K1jBpmNK1
wpXL61SNUO59yoI9OOLtZGRADINnCX8OwurWU+OzcAXMw9fvRgD2tfzBNcdxSJH7
dts26rNX13q4J8RX9Abd/38ey0c+ct4WbnXxqWWQztb9pOZZ4xUmamsqtEUh6FOg
KI58I+/NqCeWIz3uGROnpf6oTJjd6davbHFAu5+RROZVYcQvykkC39nz0o7y6/A+
gjYGNQ7ZQMdCkD4TWud1EsjLyn3Y1eig7jOpmyRsSYRYfYwE+XWOBbBd2LfIkX4V
e/lBYDQ2sIZ7mGl70FX60EeqSRYOKHud5riuqfswVFqMbVaUWXS/jrhCGxtGu2ie
iG6G0Iu+uk8Jc1FJaZSAtOyiFu8BHZPBJg0lnuzo8EhR0JikAaf+CFgGo2uHDZfl
jVk6o4ugtQstu+mSebOV+TeUA3BKKca1BSoSKM7Fqzwbmid864wIgxhnWvwxWCnq
7Voc3TTH9E/2G21jpBXtuhgXK2jEfvFdSReUuzZJvwA/oPb8rrHa2vYPDyeviLc/
eu45jSrcw9/o61t16QKFEuWK05MfyEGJ+S8P6qGJ7K4d/K3ENG2d0ToHWzrBGtzD
VOYzR5N9V6i47NiwnFeO2Auzcv0xpvIRgSRvxBoukcLDFj/jcAVM5T9udL3Nu08T
QZw4y+IS4e8ikC+o0Q0k9NgtKZ6xiIHq6ldcw8fpSfCHWA5/zS9BkaBCji+1SM8k
0A8iKhLI5wAqRHgStvd2wRM9oOifLg3hOAmZLOs5n/K+TSBx+byw+T7nmqVCaSJP
0ct2m1J4KfQXYE6SoLRVGqXks4lQcFwKwxF7wqI77PQDjCVKNeNMK53TPXN9o8sW
ZV8qyUafQ/Fd3ttHsIVlYyRTMex/6JBTRItcV5kMxtW3OJ5ibkV+kFBAZWUmld0c
X7Mbq2U4HFCZmr3uG9a6eJMh6OuYRxsVD2F+mDvLFuo4mYoTUpYs8gMiQIte0MzK
g/d8wXyY2h+wdEEr/9dkbq7d8sWpwj0Qi+s+SF8j5pcUWtO7FPi0XzjESK5v0irX
LDDhnaknaAJROHVyJWMWLx7OwiQ9kA7itrGnLue00mE/ox3GyQlEDgHDQW+LEPrI
c2AbCbS+uy6n5aUyrSHpmuICmuBRJy0dhDid6j6c0FioN//ECcmN933BWUebJRLj
Ol+HIyqKjBzgcv4weLtRfX4t+nU2DOxbwFKDFO8jDeRjzbDXVt4fs+AZUJGi6VNn
CA5EGPgfzB0f56pRFhMQ7vSVDS7W4j/UaKKt9XzDUEtydKxWzGoZTLkOOb+8uzay
10ydJDpgg/oeVT0Yt/oHFWt6TpSeHQY0fGQqI3KQrQo9NeT/fByNERzAycUFFltd
9IORllR/sj3qsgdGAQXcenDln6VHh1U3UUdaEC+zMrWsVh1Ah4iwiEd5dZ3LeZBv
RURrCWt705BGZweoJZFRgINnZOv0LoPuHQfOxpv+k3l7W9MBM+JyqPWkvxCtiVsu
03CjLHur2q7WhDGhPJUh9lM5y7g/OQfNeW6ZX+9L5ZJpHTbSbr5dBnH5Ssjk2ep8
gvhj6oT2C+BTBz/RtcgTt6pdTxH110Vgw2/dmKmcvI/rHYxrM5arf4E/rpf1gOdG
ogZtVHN2SDUB58qG/ogFBf0Bat2TSsYGWc3EEVBOQuWpHTFoJxDm0qozzaN3BjYT
l3TYGrxfBEjXebDSm0NvJId0GPrBgjPJA82UFco822aQ3zhnS6+EkXWYdwItm8Lu
zWNwglPya0uED4NOPen8hf0GYtterr1zdKLmMIo5xLHZIamQCBwwympnSu9ggeXy
4UkGB9SM/tPHXrTRVoHcsGxBydNfEQgwdOQ0AgnXgi8jYJHNXRRG7uH4M9kkBvos
1AynNdtoO6HYHw11Anoui5EErZGJXWyeGUsd/JbYIqPmfqbcO0BdqIsdyfpVcNIv
zKRnyDHnyxer07c+BUBiRj57+jJHoBNNdJkgMkHIwTWv3k++fqWOLM0xKT8RgNgd
wk0TnfcHJXSrLr7RilgzlUeyixxRmcJvokQQnHly2Hr4z3AgKJSGKLFXG1JGDVJ8
bsbkr1Jf74sqEShgOFGKF8zAW0p8GG63gkwspP+XO0NVfajJ15xo609GkWrRcb7N
niUApNESqazscNj7kZ2B3F+h7bZ2RVynrxzl1vN/NbkhRuQOMgh4x1wBU2JlRMBo
rRBI7mU2jsFWZvcVhyWq/pwXoYudQWOkGgxvWCjUL8+bPRv5iHjuQcDElBM8MITF
kFVRdH/DHpj3mJxz2tkICZ4KH5TnDMnCGDan+sy6rhPlwVWm/Nw6ZMVA9PNhiA0Z
j7fChKTFpJGF7+fhOG4PXNboEWvEr+/G7aU58Gnnlk+LwRmF6jr9CELXdrI1To2K
Cwi4CU+ZM0gu1HJ/GF5jEbiKQ0k0svUeT9e/CPf7njCjWJMWJBqL0y5wW0esbIrr
m1zjdYrJXaHjByT+ZC9xJXW2hdeX8mFaUNHb+67RpKGSkhQTmsKstqrstQxcIRin
4KRt3Ar5zQHOHMEmFXGNCnsG3VT4GGqLj3KyIrXVzCOe7/ESX3KYB1LYAt7w/0l5
nDpexm90T6XATdYBQh0XQRRIktBZB1EHWct24M6BF9biGxNEnIZx9YQR5fl/Vk1/
UMaGxdoqMTbQNnO67bC+Y4uQODuW0v/QO0a6xI00I3IdIZh7Dwn65ASZbHX7r74D
QDDL2P74ZM7GtAlDzKDyCk2i7UTk/bOhhCL5iCJYfnRVak8bbbxGxOE2XOgYuSxU
YT4m2Y9VkMD8oQet5z/2o2vy+DofSeATmCbyLYmu4pgsbOaboPxF1iz7UpmW3/mK
p0VepwrVpZs701bpCx55729kWB2I0rJZf1vQILA/yQj8qj6PGAIWsGv+1m3IRnov
cXHgbz4nvTkmq6G7q+Y4NBr+TH6DYLVqk0Gk6IrUlQxblXhhNauLn+k7g/Jty6c8
1A/z3Cx69/TCjtptAvyEGirf9J/w/1P7tlWyVyJhZY0g+nMXEaDJnC61XM7YHs0D
G86WonoF53eGJG53SiPfAoIcv9KqPRBDh9rMQv6lCj7fUHfnAuAxQ1/O0b/HblAy
Jp4sM8j4DmsxQNWNpk8McihpCKjf/oLZdPLmCWWa/uWy3QGn1KsM8NT09u/HDjF3
Q0zeBoNtT74jU07FXciLIjv96p6GGSsYex0zQ/hGptk/+UP1Inllnq33LyUtO+E7
tkpQTj+uCFIf39Tn6kpF8THfd8rg/pC4imLBdwBo9aL/eiInT/skZHp2iTqVG0lM
oGtEzgctFWv1EHWUAgl2BN5EnesM7DKmcu6/n1BslbeK4Y2nkcrN2RBKBrbZxysp
A86bGW8ZWyGVRXFzHYPOaYj9sav/Vivf7gXH+LxFsqmR0fXZYMZ6zvZznGzb3hx+
4+y5SRtbX3uexKc42zvGARQC/E8f50ge3c0yJdrF3bPp5QQbwz6ym9tOIJKDxD0i
4Hg2AYU+RtlGfBHGptoZxX3mEGugqMKG1nm0s/I0E5eqqb0PE4K0YXQI/iVr2tyY
DqVt+j8D34B/+757wGcAyZdJU0lPOM10VvNIwaYFoTFW49rj16OxJmWtCPW9RxvJ
OCdejGyuksGKLU62/tixG31EWqZkcHNPU/GMJzag1+dqQi6Rvob4CX8TgnG4KqCU
8pUE4QZwbr+8dX0tk2bul1zI0qcl0yTQksrDcdZRGl7VkeQZwEhP4bFWrQ6bQZyA
qnqckVcYeaSCqDvTFjCGtdwuaEaLBrA+Uvs2dYouxLKfZP/QoFm++ob29EBXk50M
d6qB8nIfzHn9dKI6wNzFb4yp0Bn9qudobDOuIF8MPQNOWZQ/KPwQoTzntrvxmPDW
gXilNxjOlOZ9BEveww3999SqBpZ597aJqhuZ7n/uBGG7YsvWgVQpj33nrhMLV7gY
+ak7A2vvvTGaChd09OjO/g1uybGk59AGJtJnGp+SfuFdLNs/xkIma/4w+TfF9+zo
BrnYMQIxGKIbY7zlbk8l6ByrwWxEv9Q23YO/vW/bUyHqQ7ARHZcU5uu9AgIbvPi/
/O8dBoIlgCyQKiO2HhrUU108cP2FY6gNbPH6mveGdom9Q5SRZ776mSiRC/KunEix
zmKywCzQZQQTBavud4aIWTIU0y32Wbb9ujtxWrynFvCVdd1190OYB20ntjXP58kc
R9tEsoQoBop0qD2ITdTPSVbQVYF1FYHbzr0wY6cace16u2/a6X5CtaOyPFERYusA
N4dRMEnfLW2ns8KZA2Wpzdwpfm7A32ko9+fXGL5Uk7M/zM6Pc2Jv/fc+9os2vtwi
7ZKVtNdhJ51hLBjV1LOi7QSoWbNCfupFg9YS1SVhnrXjoNFHR8dAuQ41dmMBkMWl
bs+/jSMXAO+IgfrMVqVAlhu/CFgE9iJG/JiCavCOh5DWi8zHDQXpmKKgzmBUt2bo
qjxuG+1KFBoHZ/wkdYPFLmiTJc1lv6Qm2y0mEORJB5S+iv99X2N8jzbfRKug6owG
52J9CArYpeABThBumwToonVhjFJxa7z2M/c8vJ1GUjb2dp4r10qhZOWkUDvZNXqd
q6uLhGl2T4KmtEUc3u+FdD2m/EYNykNv15Jx3Yv+L3aS07lgeYHzg6issoE4y/NA
Zu55RQdsn8LM/+PULxZTJ3FNP8cP918CH20hnojc0RF7oQibc9EV0BYx/AJPnRNP
hDvX33kjrin4LYsmCcWLgPetGMJdq90PyBrfEqefqENU3oodl1YMAf5SDWyMwQzE
opwUgdPYGZx0MbAEh9pd+4Bx6KfWedwGAzu+jE1WT2CJMF2wW6waGXMBfIo55X2z
O9+0Vr5m9SOZ9x/fazLURLUF5dhianNUqcSK4sJ9fA+rxm21NnOIuv1xDM8rNPJV
sFPIqkPgnR3bk8LWJ2Vwv8NRgf9fFkqCyRqRC6Nb6lEXdkykMjIXfCINExj2Cdmc
rGwJygHZhrNm3AfFn2zA9ppDU54sOljJWLvuBLGOHe999ouh78tnvgeY6Fkv/xFg
L8x0hRC2QEbkqA1KAHbz8L7WC+PN1luOerhbygqIW0Fuak2bKg938a3eZQ8ltzmw
o8OkI2E7HY5wgLjzLXon3ADomZlrlo1W4rW/4qPVCkbGouAc8r9DMEj9b3d8kMjQ
cPUiK0in+BhjlE3qAXInrKjtm2W+9ZRyKbccsgULwXpeN3G5QW5FshxswhK/Xq5i
og02UrVlgvE1crvHDbHmjO+kryzGBe2x/l9SsmsMg3daU85s6SGmZ0ehszCgeHJd
6rKe1+lx0DM/nv3LVi4J5POkUPetiDgSSCf5wesWQg2mNMXBk/pWzfL0ntcuxCan
vNLVFQY/qDoLQPO73sz7SmLcFhIv42sn94mHnhqB6Uptp5lhN5lnP6ND2ycEl53l
a41OdD4X+opfi7oQRu2b6tRu0uHqvitU58wJGqOJYf95hExxD2VfhR++E9Tr18v/
xxw7xQi5Yy2M2d+sEScM4lE3zk6WZ/s39vxXPBoWpgy61ohHM9/8rTE74KFP18T/
P83aoZKFO1Vlo8/0yS8w3QZu0aX+MOuqwjN/R+Sx/mwd7Qhh1Uvj9df6mFBiU2zS
47VS9icl+gb01sQUFd5nIDRZiFFtrbuafnFNCTj1H4AShdqPLDh3ky8UMevboOuV
0ywNgj3AcaQu8yBOLVzX8vf2VUBT3yQJbEyS1rJv75WvPv6RUzqyO37XzZO1iQwg
9NtNGgu4OMg/m+aFdwjrgV2lMKxhhDOg0v4PVMg6yLzHzgLiQoaX1WNe28/qY0k5
jRgc7FmeipeDpshRCVCJYi3kyEDoHTKw2MPVGyZQJWbWVOz+OWoWRaXKOAkQoGCP
yecOAA90cHBI9hGOBcF0VIqhpFljv+DchU/2W90M0mJ+ba8+q16U4mhU8wRQe7LS
nLa8mEPnkoNrY6nhyvO3kihSTOJWbEX7vk4Ous3CUU/MtlN2WdFQwnU8cNR1Yz6a
vj4SAKYir55FasnNVsNQX8UaSbnxwag6hQYjdzdXQCNPmrt3AMey7eZte/cYi/6B
Goxp/I0nL1RdeWBM8BBSecEP58OwA6PRkzc9EJsFs7ABFy/4J5PqMZRJHYDhWboO
emlGB1hlaVrGJBWrHZIxpTq5lw8y3Lf+LCKeZxI+3DuL1lvxTQu1yd8h8m7Xd1rP
65K0DbflqXTty8swsRZSvrzkneqntXPGRC2+WEVoRepEqN9rl1anpSFSh2YXZV2t
fjTY/hB0M7EKKZjcimW8q0L+2DtLV1zjJG21vauJJlIFhj1iCJoRUWfi/IH4Utrc
IRCNCepI8q4/oRuHw6ni8srRh4ggW40tmAPfF/fXMGpOMhoaf6C4SXPhi5mW30/9
SqJUkA0pCQxYDF1+sUgmVvtuciVD2saszL7ir96vEAmK97Trt9gc50ud1d7JHRyy
rgOR6ROJCueSOhp8RrqyOA1IZqIkKGoSnbRotmNPDC4rNkGX+fL5uDbZYO6ig82T
fzZhgbipPBzh5RzDY76v/WohjhyA1W3iwgcu2paSeWDTlGWUFGwpNkLsqyLN5F/d
BYbNBd/s233zIYhPDBaQRc7fZTqwDD02Ezx29kDbkZC5Flf6H3+gzT6bIpuUTeC4
gXlQmV/U5e8z26mMxBxQ5NoS7t49kHhrw8Dy17WGiI2MfSI0KzqjuFcH1BkyCIK6
a3KBGksIC0sogE0Dgs07Cnhwhg6Q2vohxu/rNu+v8fclP8DXwv8LWd+1m6uFVUWk
BsFG3mx4bIZPbReULGPQimkWuOOFFilJeeGEdwzYut6lpSQh8/KCIJIGp48tzA2V
fV4GDCwN1WbqKZPvYX/y8lOlyGNhE5IaIVYZsBdlEHaaBYsVum2suREiojsE8jqc
kcGETOdj9+em8MG8ajLPYpm95/5Bf0SiCKZV/Wog4TyJvw0RM2yaPOA9IjFZMtNU
y59usBtlG7Dvdl/vaHELvcIK9mpLOK8FJk478rwlkvL8x+CPYxuACZSx0gKvm3mD
pSAWhSMIDTdMfDcJqZnw/G2V8L/T8I4FVjXDYVIM1/ZByh3jn6AIaK4iJcCCz4IJ
TcFA06c8SZwJQvSSrey3Gb6qD9wZnXyCrmvd4GcoKA0yYE1x2wyhDBLQFQh6hj2X
SxNnKiVbJqipL8iQSRArWcs7EPOvCC+gp+vFNPN2++AajwlEy3UyGTNnHZU7NOQZ
K/D7PjZVkNS1v7OvLToeRz1aagcUtbqssfZAr4V9WC9qVw2+3k6r3dVtuc8WICME
umu9rgukKRKZINfcgqqKG+38qO8kpSRrqUPdb4a9DKSRZc1zwAJQT0j9yacTS5/k
0DkNG+WquMDibyr4jO4RVEF7gy2YBagmtjRIL1FXcmPj3YMhy2OStNXEK/7Ck/fi
lXjBgyEuJ595u6pCArlj3t352ROyBawe6yK56ubf8MHmSIIebYHhCj7ETrPl+0YW
ZdvCFCa2mJ1Onpjxk4AOCG0j9Ab2PQEOhnfhaGJ8/ytymWgZeaYWjBuj89s7g6At
s+Q1HlHFbj/ay7xqWu0WTsB50HrzKhcspo9H9WAf7Qp9Xx4gW9vmUUJB9Sm2Pk3q
VpQUt48cMSlVumk3SecRw2mEkDDkyMy6JamsJU1Wed7pSUP9m0G1LIHKo9J77z6O
URjNA8hWF8Xz7sJP56896r21+8NFHfaJpJhPEYYAsOPzk5Ut/RUK8f1OMPd/rr0e
uCWv10XltQzDFs2NI7081LscZ5jcdGHLPLgRqCw8+D7psYKU5U7FkFiAk5HSIz4E
ssvX34vYQaPBw74+O1Eg/De99cABxGCRojBKcEt5HaEum2qwSMdLDZwGRNBcYd+y
g5jgzczQQHUIYBSYo6jzRv/RcrDkbVEv3PIJza88Nq47lpCBh0EYeuesyECUY3Dk
wvtxcpy3lKmcVSIBmKz3JRyTt1afNusOtp0PMccyGyY5H80rbS3isO5IGIMjz1Vs
l5C725z5zCaMV7+uSXJz8MWyzezMf7n96X6ZA84rsZq20+55ltTZgqjs4sPKjLM1
ZL2bxZwJyJdke81COulAwe7Q8LdOOCjH+JCTJ19PhgpHE0tGV9TV7bi5ZvrGiDHZ
OPewBxbbSo4Z4MTzKUU0Jk6pIitMxmmZWJmYGyKDtPyFH6W733+ksxx48yLfeAUd
8ubKNPL1sHInLIzrPGJ4FCiDUld05TiQ/RBaGFULhjeha739UQ+D7FJni0lCdOWE
pIlAyRendBpCbimMu8VXEbNRFDXGKU1EMLOHpAu5gOcz+dDc65tKgvY9Uhs9u3H4
mS2WxJNqPLfnUD1GvLcheOoUpNfCF0weGUQpnYJScNp4Txw5Car2ne0XC99ccnn4
giW7h86OukztBnVNXo11ci5mZz0hXx1WXBJPClx0xft//PON9/Jz06c6RJMdHwKt
YgeCklrZGfw8oetuFOhP4Oayz/aHWbgceOKrp1+/xyxuVL8LE8MHGuIXyUWyx5ZW
prxfk8BOO68fUaZw7WvspdUXnahuq+QublKDxF3NTMKDCccI4QtUWLF2yWJ0dbh+
nFOJz1PnG0GjjY246zN1iBkZB0Al/Xwzs5REbAE7Q3hO6cxKD6TpH4kTxw9prM4k
i8Qlr4zNOPR5cyhMgTnLodlEU0SuaCilMrVY1Usg/Eu3oUcFQ3Lx9n7CDZXEMDgS
1Pl7z9wMNiBsujgg6S3sTAiUhJqovq3NuaJNmWjb6k2GVWFuyk1e3JgbPgS60LcR
D7j5Dxa6x3RCbqAzvv7ZxRoWTD1o5FBP74a56Q+Us5wENBWlEa9hTW/4yARZGbwm
RRg8vgwWr6ZHRIrwAnRlBIJxJGfwocSlmMdYQepo6cekisOCYaS2bWCBL4fCkFmd
Eln55SDonKqmZm4g3rL/rj6doh6lgQs6l+scVXBzd7QMkkW6ic5bp7MN4JGBL5CG
t6qdc1An6sN8GviuKlxCF59bJXR5rpCs9MJEdRgDQIXzIuJUPJzqnqduYuED3ZXE
Gn1bezYVEbgzyW138xxfN9Fqwt2H49Swc1l4eqhfeE/DhQtYTO7cu8jLrTol+wsx
z82BtNyhxXHqTAg9P8CUSz8DlpHzQl1GgR1Cn1pm+zDZPI4pDz9CzNZDMJeCHxw7
C9aLxnO1AyFX78V1vsg8IZ0eiOz/Fe5BAS/bdXVfjAZyOF40B+4rs86AgxqltfTU
UDjody5BggV8jF/MDuKP31kd5XvgtEoBxGBktjx2oZx80qcfu5uMuSTldsSB6FTH
C4UbFZ0Wdp7bWdi+6MYnVfQPLi1+v3pGVfM+DJLx4D+ap5EcquNpJIkVJe4wR1Vw
H40gGdRHLRvdDYl7xEUb920iT1t8RnGKworbMsuWpU1V+vlplNuXRJ5JnVLZTl1L
poQXrsl5iY6JDIQ2zzisc2wSv/Wh1uX2ArTn2KtEBSJhp0EenSmUNnz/f5iKPEtc
d5w/oxnkeZnDO7ck68UrdgmjejK+z584lLJr4BF6IGT08J3kpftTqGKK80SCOus3
ZQuIogFAB6hV3jXuzYcMsEWJcvE7+1zsAh0m6oEPa7j/gVGjAFYXk2UdsIFe+ywC
u/dxp/+PgKYlWOgBNinLs/FHnGCpGNwZI5z/rqL3vIQLfS3QyA8jDJfbYYSpEhyn
OhA1NV1H2cH5X7QhKINLBDUGyQACVTv4JDwpEhVrccR9PqsrBGxiykHrin6jEU0v
W0GUSi2D8SfV4k5E9gqZKG64VauWfdqfX3OFhgbiL3QE/O+t+qD17RgFMSru6IV8
wc+jx4xlsPpvsz5evNDPnX0JQlxZcw9aCRRgRR55i6Pwjdpt00E3WBWO7/0DYGV9
QiuUBqkle5LDj7GIH2Wb0zrWy9JNltx/nPFxB3YQCVdHD/Xf3ysnKB6cYisWggqw
9rYa+pQnXsXgxc/nxJzU53E7Bvp5+iWKqoZ6xldoZCxc2f8Ff+jsHiM9sq/XGAB7
KlRhwCyeODdDpyiGfj03H+lYOdLSqCrUy128HRmU8Ru3kAblS/KCCtz+FFl8yuIb
WelJDIArV9BpVc3uS/4r0TRqH8/gDAlG34ogD2azsTMp03VruPvmbjSHrDn2ys47
6jRYFVho/PnbDtzErgUiDXz7xis0N16UH3YfoD0kKTND3+Qm+9LC1XCf8i7E06Q1
5azI9UtLOR7E6XxA1LSBNsJnYwWJfIyB+752UydRO7YgNXCaYFgxTvOQJxTLo5YY
0vtyS9/fd2B28+uiD3RuFctCi21SvxK4V0Fj6qwjB5jpYMWcMLGJYFH+HyaztpBN
QKlKU2ys5Kw6zwhaZAPJongoOOLNJL1MP118dRgSv+ZQ+5d8KPHS4A/gvV4HZr3H
vRsMhg84cSCsgLZAaXTSrDsqsR2jF/iGIv7icXe5rpMmMEIaHE81H+4b7Wd1jer8
f6Kgt+nH53x0Q7+tCZM/MwpbNQ9xqH4SVgrkzzHgKet/MB+GjBxIjm9NjFYk64jq
v+HpWHeXYs+rAOH6SZr7vwsppVlpVeqCtQ5+kbTM+U/Itrbo67bZufpXsUtfK1Yt
89FmjkOt2aGdGaAXA+hhhMShZ1sgUes7ob1zkCcxoeBuUt9qqsk+cnuEV98D+AKQ
srDrs5bbHqEm5ODtOJrBhJI3i3gSDrEyHIi/9St1/XcSMOkVwryMmLZkm5BeOmxj
2/n7jyXs8ZEBulX7B+auwTQs0pOlSZ19Rz5gma8rF/tTtpWZd71I5+BsjsJGrwXZ
rqtZP13lus7+IoAJwaVhGx2ZHmpktk6hrGQMh9+JYkOGrrWvU7H/HWRu1vehP4ee
EKJtIi94vroKNArAGJqLr7UFrYVkZgBE/aulAvvm7ueXLaNhUPgQVhbypV0flSB0
xDSbj/hXUw3b92LARXdD2h+vli+1uSUi7uwkSIEhTtKuRb25IohYm19O5uv/S5jD
IWxQY0F5Ig/h8q4s17evJybBiD+epxt9cV2FOKi8+uGm7UNAdE7i6TSj6uY3yfnM
sz0V9FJKh1ziJ+33ZvgyE3sJd9dOh88iPP9+ZFpP1+YpEETky1DnV9vxE6JI5V3G
gq0ahrWmxnp5TwKdxsXkfQUZf4/FNl0XOXvKpw0Cf26ztnc4iwtz7fvah+nq+GbE
5ctwTzoIzUVe1LPFDTi3Lp4ulni+BTZfIa8cBvyOqfc3wc81+BC5AWbF9FgmPIQC
zBcWN89LZgg5Bj1SbjiK0jP0lSTxfKyGGOTBaTlRmEdyqMz3IrctR/qgXMeF1QLM
eX1iGXYZXkB/pdK82brSmA8AfbvaTbdP/+TANBS85krrtQsyeg1lgiJXliD3yhFK
IsSmro3thxK/4yAM+oSWRe5POr/JvX9XwYpY8cCCXRHLh3+M6j7Jhm5F4fkMnKnh
w+U2KCczqGmdpr2FapHcI89qwl7Q8hnkqjXEpWgMENyswVrfvaucBsMt2RM5TJGA
Dxg24xx2LNhtpWo+oTz87WEoBfvlG0mJZS/1+1Ed8/QKP+64+c2DotQK1WKyRP6W
SwHuc9CzHSSUAceequPLvTD6KMyRAyfUiF9YpIun+7y74cIatBsBG5DqoWxfsX4Q
xA2+SG+YMa9xn2YPhXnwlf9SL8OxinPHlh76ybkn2rE/fvF0OH+M4IcqAqkHZde0
vHre1OAQm4c1MC57PcvYc7GxzEf6O/8UJqLCH5mypS73SRwv/ExQJFQBj5RVf76x
cvmkdYwuToB1lForYRHC9uIdQCFdMw8iEU2WZGvs+HUgBVTRoXhZMHqqFbdmSUX7
egnr2Pj11ET/kCSFQULeTSp2Vn1nhIu054HTWML5dTUI5mxIQkIqUOgtsBmrA/Eq
pKcvVrl8cNvz7nh4QVMPEgrfynfjybALlR+MsofquxleHlJOHq2S40+j9TKi1FeR
vgPEuqfphQTrXJC1deksozezh5+vne45DTN3tmKmfTAxTGw3at18yeSL4UA8Uvbc
BAMfPVs27HBj+p0m37Y8J8A+H0qsfOQt++ewAjLHj7tA/XNXPbrQ0oRxOJpf7aZV
gbHdwAzEbimBi+QocEKMPuBrfVblQci7MMXhnDx8StHpKfMPknC7lTTs7EnkoFEG
A/JoELL2DFVuLBMPykS/TrhHUVwIz0XsZzNDsDAV0+yhaEXQNoVLtR6TjXxUV5h+
8NVg1RXPZ4hItrh8fzcmayqHFoD+32NLgrspjngHD3ejhK33/qLzVZ3qOTlI1zVw
l1HdJaKBteqUXyIdZfvOgHLg//QAlsXj+jL3VFgt7XnfaGWgDMQjPwBfBAq3pKpC
QB/r2R5yVg33sZejPYDf+uoe8qjFgRBGGiD7SFxR9TgeZGpPMIqXCYgLJtzHkVaI
NgOOmhjf3UTDazIb7ShdBW+io9EWHTBhQeIxvUr2jVes82UHrAV0shpp9eeIHavv
AVnePv9mkcLbC3aKPcuadCMdze2a3xangPALJ+IUZiqZWhwyma69+EhwrNmyWa8u
yJcyP3t8nL3uZW+CdfetcNbHK7/nFlEoMZmyNY5ocjm3iukPosHUGipQg29rYueW
Q0NnZOb6v/0vI7LrmhC3sheWILWXpp4N53ugvjT+TRQDIrCoooJ+MzybFBnr2UfY
tAobRTkrsafxWe+mwDq55AXwOq8TZGCtwOYxeBWCon4+S0vNQhGMOEaP3K1hswfR
PkryZan8Pp5UMUI9i9BvPeY2hSHmcAAwRJ7XieJLiqtDFARUobzMJesCD/aFVmfp
lhlnwjkpVwvnnT+6iT/QVN9FZRhOt+HmlvN/WzDIiwOhd6LOxKn1xSU+Uc92nMpq
fbrxc+yRXwzQ4KSL/Z6Tc8d2RQO8em/YhxsmHnz4ZZfcgYF7uAcP2TKQuu/O93oB
mn6VQXpnP94WS0zdRxNdywmc00v68QJ8z66U0V2wy/jhObVQJ1ahx5gY6UkUQx7S
JVRZkpcPLZmPDeBqYLf3cKW8fRNxRowBL7vXD4D+WljAYF/udJUsUa/RcT1tqg6U
FdQWJlwLVTvKiCV6zpRf+aLf9DCIq+JeJ4a7iGpuakVg+MI1bpgxCedDegrshsG3
NOc8EIfWmO0c0WTYP0oOv10CYwjJX8LZQFlwzYavb+aPeb2xGWk6BHrAEWQz6rPP
6N1f/ktEW3TWRYQhBlo6FMzCMOEJTtqLw/dhAVBTvYP0Bc1q6Lw4TCxhCs2lVJ0x
YepyMe6OGm8lm2sDGopYsRnuW5EnozbJng/B9ganAVADS7rPZp/aNOqEnWkgyOAz
Ow2LC46H1AZYhOCyWT127x1nFuGFwhO+TZS9C28TDUcnxChgyR8zfDB4+liuPFHE
j8eq9UMuHNMI18oGgK9MgP6qvoHyfrDiJ9Kf84DP+GEFp+xflNqPi7k90MAoTqq9
XOmWaGPLKat344KphFeILoUyjJrluG25EbnBIwJ349GzUIyzPXOGuXYvdKFzt5M9
m8aV5oqKhAAtAcQfDkUfIr2OSIASxeb5ibmp9NDggaD05xFN0FPVIW8gUP0/VEGc
55Kej6Cr3g56J/MVnNWqoya9rkRzWaZCkzC3AD86/ogPd1yhRW39n+nHe053f1Zf
J0XRS2Eb4PkRM9jt/jqjVrppCXrYGD1Z7iTqwOrh6AgMC5GgrdC0m+DftHnUhdSt
CJEDHk2YQN/xpFKBW6hjXxElmbEo9apMTk3+gcWSkfXQKPk0vv7b54t9ATHZDdAS
F3DjoHgPx7FgcyUjmZttvoT9lCFnzFJaQeNbpOXHoWKnwPUJtIlizGpZScLC06eA
TNoZddJR9X2wTHNEuI65sFcqvmvMTdrVHNJ5xA5m90BtX1RvByYo9LmeOKTJkVqo
QOCyFan4pChVXrhCGHglx2KTSVApHhaD1x57mStcuKdunHD5pon+HfzWxFxNAsRO
stm+WGeX92k3cAAuf4OLn2uySHPZPS0Q43eP56DPq+5VTwgjsTd/SzZ/2gT4DJ2N
8ghHfP8S7dm3xarii11eZlzADeKMGhq22/2XdTHMsQ3RnJFSdgTsyBSBTvZ8qhx6
9jf5As48qblmwpa+o+4S9GfDQVvGOFS3gNf7nTYbKHmqtmyPBZaTMF/zZ5vUJlDq
GBjJrfk7IJJlzGijLnR69W0Cu0IU8RymwatxUteUj99Kf4A2XiJK734oamDHumYo
/2wpk/CpP31ZHK1EsZnDEemiEN4YS3F/8J6PVR1mb5m/8aTKdpWRO9MO64CCnqCg
6if+I8+nVs46HG0OSdABh9aAOxX6wj7yN5xUuJqw8BgsIotbAAIPXf2Bix5ealn6
SE7hgMKHKKdQkYiBTzJUw3wZ+9G4sPqJvj51B2r2MT08IKLucBrfFS1c9VDc078s
Xt+1XKybj5xgZZsmr9dcVV4EpZZT/Xsya7VPT58OXzMe7vzBvEx3NxGQRhjCeZpB
Pm9/MOqCVaA1GH+Nn0Xb76fUvS/p+988/vV5nwDkAjq17yUrx8L5eGvOjGVrdtPA
dAn0E4lj0qZ8NgYV9moIco3TjRRivCUSRNFom1PUIY8FwvDE6Kbyatn9zaw5xrAD
Eg2kPfJ0ztTwZFXL16nlneWIG0HR0+wHtcowzTLvGi5RPcYjkPZ5OXv5DUQF03yc
6K9FP51ZoQ9wbvXpw9IqJvvrF573ufBI+yCvJRjXQQViRsE7/1OlWY0ZZ6pyZBV1
jhz7+qYHSuVHvH3uM4K+RY/KuFyO8w1xQND9Srz3PQ3B4FWK8/ttMjikOqRhGMMK
1buV/uXf8SsB+O4ynekFyKodlAFzrTgZqO8MJenxBlfv9LjXICFB8T/LIvaAucMs
VJdvZbrXfHjtlwg6q3KrsWwkdcqwHniNS65dFmMPhAK4DN3UWvMMuslaZLlWKEVI
3z0ExykkpUIra8114SANG0QX0rk++7S4hdi5J6rJVuCasYGBdDwgOcbgUTAOVuxF
iN4TlCRvgiTU03gSqufMrZSebmmgx86bWO5vOsCXnrQDaGyMq37PrB22dvwB2yHQ
/Yuzbjag4YUy9LoaSVVrrd4ELAOL3SNn9yso8kxRk9vfyGDOna6oOGxTtQxi2/u1
LPQtaHzfQrG1ajCP/vL76wE9hmrsn/oKD51StheYeRlEHm8GBShOIUXK94+OlPdD
hjSmpH6jYtXphaN3/cDtRtTEFs5SN1RnqOZX9b38zoChrOcDwnatlt2rraxOYpUk
L1yXI0GIlXvw4PgDzrQZBMX9oZ2SmClpjhPv4fLBWBLcrgN19Vq0ruLfj+sdlUkW
I5dGdgF3qwEPxBmFb2M3ePk84nxysvOCgm1Z/JwD13RNbKdbakPAwq6iHxpZIUZM
1fNGOocywgIg2rpX5Hp5IzZZZrfO0VL1Ik6ShxpUdImnzvNS2yljIEsqy2yniuWc
mZtb59OZGOQOdaB2C7qwIKUfPLrHKQiSi8Atgrl3wOZbu+PrO2hq67MxQEr173DY
WvkL/zeb1vMmaVamnyRajEQiWejA/DfMhV370YfrIPd6SJb+rngIGz1TzO04aRfa
Ytolssea/nxZ71cWUEWUd6b76On4NAlr+JoxGYQblPj83O2cdYN64xd4BDycibmR
SwIV+CMpt2yJpmoCrhECAo9j7TRpvkeZz1W+yqgxcOYyBd7UOsB2zusz9BVW3wa1
bBVTrONBwPso+KIpKR2cRLm9HskimOq6WvPHlDfNssQIrMygfzRWQ9CpD32xBwTn
uY+IoB9eMMd0VEVY3jmwNxLy5zJLRnQAcB2tX3G79Hb6PF78eOe/NghE9B/jM8jd
AbVs2f643roQM/FDyB15Eh6QGX2FY1kSRnVRNFMuogROUPf2XU6mYZ8vJC1d9LO4
g6JZ7KY5qJrQWDioqA73mH//DbfzMRq/WXLayzECrqmYzccamSOLNpu/DlqnMTcd
tAr24lP/06uPh/o7AptLW+EIOpebw42VnmTdnMYclmAePSZ0kGyDaVdlKjiGVrfx
ShJThEuT0O5jSFbi7igUyL6fze/wTG8RngQ6I4/dnAWGCjvoQzy3yZzbt+hhCQKF
N81krXu1kaS+DaG24jB/+yp08UgxL2oOgSNx5Scbzvog+2Snqrfv5wlUAGwurr6a
g6Ul1R4sYd62hI6g6lwdyTA/1QpViJJOXUe7XvGQWcmyEpjv1AZlZzYXS3yh0fat
oCNCHXbAbbM85RRby82HPoFbGGLA673x24W5AVkvJeHGonPIgjxA+Hyt2OG308Il
9RBQ89TnKhwEm5sJHhBH8vHeq7/bmmid+iL8fk7cbGvlDhunUx70yrHkXekXYObK
fOGCEnSgKbZHm7JMddaCbQA1ngXnDP9pvuvS4v9RjyH0xGoCLk2PmSXhpadiNiEz
DokIVZ2uiFF1YOCdDCnqwaqf4bU/J7QGIPiFNwrOh1Zm04shoaPqbYZZaBJxmls3
f9FMgizOaMkdilfWt0CyRwhXPHOi9MmojGjcq0j6TGfOzgh4klRH4ip5djrMxDBl
6Nf/LES+WAw6GQciVVnjWlvzvL3ysfsSZaOHzU1z9/mZlwhXUgdS3oVpspvKPlMk
bvgD8sgWTHGEokRmQHM/CRHn4+J/OpoGL6xXQHG1+4D7UJM1kxHzeaNVGZkNR4j9
2AG+hgrRNOa8jMSrs6+3cQN01YoXJOFiry79vvwbOus862j7PQ38i2XrguwcSyqh
7xde1QrciUkrKlDB1Y0l/nDMEip4+z73nwwPnW25bT/yW4ro1JQ/3FFt1B8gUWJY
goOqjOf8+cJfq+bl86ic76+VLzrTCpkO0KPVWbR9YEpnB6EESGApBdinJ7pqvaLM
9Y3C4T2L95qYE+v4lMSAyOV8nguNMg5h8yg1GVjtQC7FhaIiq1Svswkz2SUojZ/P
v2kB8SGmOE/RjnebdiMbeXwISzHnZHHv6QWLt7w91zVZOl3y8oKbLwY4jbYX9oO3
0jRPscS8llaYrMB6SiIK3kdWTNgFGb2SCdzZMLOolyZqGGftUvvr16QV5MCXPlcL
4zsOsm5XHFE3stSLaazqydy28ViSidrGiu798Qh37IUk1pzgyB5xXUDt+xZn+MJa
SIxLiJ9eUQydW3vtWcDL8um9noed7Lyl/TPH2K+qqchLLpBp8Sv2hWlaMvhdH08o
fLRZoN0vTYqNk1GDEo5dHUyr+zKS0bocbY8dmhC3j0/LlUcGA0A7WKvl4SJ9IHqg
7kIa51WPdirT39YVVClOLOeuv7Lv82kiP3UAvxvCihowcGGzXR6BGwg6mIP58Y3t
UwvNYp8LL8Nhdo8MNO7xb1V8TRbqMiqIArlK4DY83vgXBIlvrP4WWo4u4k+YaUPk
hGi6GKIj0xNgrzJNbJ86An3/JxK2q406KzZoSQ8xUpOGfWiEgjsZ5qFWDZ22G/CZ
0DaJbsbZWMHo2WK4H3Njfr1Qjguim/FwCy9aBiDsGF25f6fqbpvqy1kW1NTM6mAK
MeoEKdWTkjLQGD5BXGbHZBrsuJOckNiPJNlfBtdmJV/Z5oEPg1PQKKCG2ICxGdEr
KwSGHQO9G0IDwvzS1RkFzOZMHnRhRPBb+DYD2UOB7okXJWdzYQw/TesXsZ8/ljw3
23BruuPgqJWJZBbzFecaqB/NL8jOyED9g1uy+hKv4fdHMRs5NEPjfUXNPmKRVqQd
elUFhjD2pK9KO1R6u/+GtgKWLVN83CYOhHltCnZ4hyjpSVR6+KJeVT3qyiQ0vsNe
rq+cDtWsoR9VlvLRyA1DbuyvHRmQFLXL0Kn6KGZ+LTc7E0wha2WVtBVln87w5BEN
sjViz5i7cxD8r3teo7EKy8+etIsn4BnViwpHngGwP7M2uw8cZnGf4x+kZZPJctSh
OrHk9GkzKyoIWmN9S6Mo5l8KQ193ic38qRIZ/vp0nc4qFuIpqFzADA/BjhjVQC9M
TOhABkviP/m/MxNZ6AqR3O7koYFhD2sADUdzU6eza4RHOMjxs8lkkRmCw3j7pnpS
/X//U3kAaVBsKGtpSvCDuOwk8B3fF91kTmcJX5BbP8hklKb5VbwYIJNNZ8Y2MOdf
aP3UVie8+yypyV7T8n2TwoohxX6j+mKa06dWpMOVLCGJJgWSYF74DVnmkfKtfbdh
db2cua6NLMnS28AFxsoZbXBN3pG4sQJGRGojct653sgm66NVBJeUGW3H2jlJOElJ
+C/7u0jhvVWn42DOGGAunKmbs2y/EhT0tKmjpeweWiy+p2nYnFNXoXbAqdPhnREN
5pWRPp/PWE5IpSIkuGfdIazpZWkmeEe2AImrKEtgT377gTLCKAFqH+tWT6vCX3Kl
p7UFSlmKIXgB/HStlsgWnTNoUlcAFUPtDOYfzX66BTWhll8d/I6DFTx0c5l75CG4
DlDwkpiH+lIKADxCQX/oN4g/pxZFKQLgqORNfKn81J14LfY369jDvFpQqbscozVB
a/zdcrIkMzHWrugP24WkvflfMOvxPMsepu+vziYmkrsev7XiG/33yu9DVjNTOiDy
lxNnXuP9UjNUrbV3+YUcQoxlsmRhswNhrjnMonxkRlqWoWcV3EMi9MEFHTSnB+FU
hvx9uZX0LnM56FYUM6xku6Obj63gGXOaeLDZkm/aO6NquTVb023yN1Iza+AVrIox
CiY3GTDxAdM8aH48dot/3a5jFnj+kspvm6Q5IPm+UfxmPr2GM1JwmDy4SWow86Lt
Q4pnSRsb24idIMUhtjlcb62XOg/Bv0PnWwmGxPKLAZ1y+YdLdU5J6wb9sv8IE+O5
XottCiJ1+oC75zPtormA/jVT/3cBGOKzP8dLzIxldweg4i9/UMg9CY6KOLGSNrc1
6c0tui9eInOpVqFxh9xBn3P+AjTCiSz+0tbuvhZTL0FJJRWYbHY5EY87+A6+BplJ
wXOtUHowsWcst4DeCqQ0dtCYGHxl6ZOya0BzBNaSjXoZ1ex0t+5t7046ueGnrDqv
UU0dCGJZY5O/RbaD113RHM1IjkeqX7H4d2Q42piW33DmYIU3FU7bCwLBE5XqiWU1
uCo9BzvOyQe502S9Y80xQQrXODZDUfqZRzmi71zE9SP4T4cMh8r5nRJnGPlDBo85
hKKFORNrEKxvxvWm3sPYjXjkOEyw5eQDJ/yq7Ivlgm41EXN8FclZlBRley3NrBRa
na/hPXbMPhT/gZu1OGyaXUtv7SAs/IhZIOAqJpTAm6dNPH6oupzlKI1K3y9AsqOV
M4HufxxBnCV21fA0Vrg4xIs5o47lRZJRiAtA7cpt0w+TBKCuVDF0f7X4LgJIY7vL
1LwtHvVzeEUuz+YmIFrTFPKeE/yzPv+J8LURe0X0E7836gv67fe+Qprm2pRhM78e
bca54P9HVKofz6Gjg5o6lPJqso4SS8ZPn8BlEHnvr6vLyVxE/0V9wHZoXZYceo+Q
y4sKHltgkV7MooQYDfKtDeTSwTyloJOEWTR/5mkF9LWwgVAEskDxdpSg4QyPyUOC
yTe8siUtg/sDv4B4lAIlH3FfSgAyxJGBx64d4Wa7Nnzj/OFJbwOUsCHKnU8tB0pO
niIXUpAB+wVFGYgRMLTkIjKfsGTyfJBVJORQ5rUtbtTHc7guBlADNNOydIOgJJVM
b1RYeb4KFlDqNP6Sx79ykpK5hzqIOtFl43x0E7jC6VvRzGXs0HY9ZDx0jd+xG/hw
ixkT1EhSx/3pf4VwvQPk67QEEg4hxJPvllDuxX7xPJ/pxHrratPiZnvX8Fttmcfr
OoAw8aJXLwGfMA4ygAxGpnZhNa6OodgPBp0/3Yz7u/8n3/w/J8EIkxTFVGgAhj4E
Vxb31g5G5Do3drTxFT9q1r7ULsXqAAd1caXW0c3xnRhOY5KQh/kNGCyWRPejyFtK
Y1ttZgJ2OoUG7gBIRoum5rPzQM8twVREHH5Q9oSdd+8DgYRSg+XxLhMfR8WGEzjA
1tA7CoKQtj3Ofu3B8/zojeOQX1G7rrGjzJnX7YYtfPxxE7sR3LzpLJFFg0wxEgFe
LLGMNAP3xkzwsREPly/5S24mgXx2HUWr9Ej1q6stqDY9yNnM1YvM6yOK9IK9ZBEm
PnrxAbXSyqNgAT68S0JNRnwT6l/xun/wr+glBbmPcHejvWEWyIJlOwNIDRWvqB7v
K+JBmME4MDh5XOMFoYRQ+7w9A1N5WKxvyWEXo1pkfYuyVpmX+vvUey390nu6CqXc
l101fauqUpDdNZ5WYvsmTT0t94FW+msSSS8fzWmLGqoYXbJZ/Rx+WIXFvKG8wHgV
luFmgApLiMFEzSOjPRkI9hlb/wEmXz1NMSGfSV5JNr95rDQ72U/x1VD/Al5Mtpnd
fQ+bzCbCkQOF0O5iVUA0CSP01e5FEI65AX5fZEnXS6Mp/0ubO4XO8jG+1q4izDqq
t0Q0CYrjt3wglp5rqtULMAvuWWEc/i78u4EvhZCAwT02iUXB74CzgUKqKQYCg2rE
83ZO7Ed1q4eWd8WwEL5sWLrmT+ZcKkdpmU8kips3AEj8MWX2KudxF/+NQOlO84ya
maUaOWZXIHooIM146DHxeg82gLYvxfHN7zu4HW2yq6bPn/VEY5l4teVjTrONkMqC
5mIWXRabblMgUXkQyoE4MhYse+R+/W6SojVlVHDz27I9WWOqActMpyv0oUFnfiXj
gQJfPVtZm86C49pQzyRVrpTc+tCSxGr6CogQVP0WNn4/bMe3QvxnWmHbRtIZngMA
nLyun3SFxw+C8NYYMu3erem/f41S3VGE/enTCl7QN2O4kawsd2XGf9NAE67+oUB+
w7WbHtkXdGdfdwEqzcQE1+cfSMS+Rze8ipKKCOKeq6KoFUdnr3ByggFir1iSQgnS
aTyLp6zORl5wnweML+4ybYOhgq9CRNsM/Sb5/A+CFvg1C1xlYQ1BOSdNBIMVcgGi
q+4ZC+Y0S4HQGjLOcOwMSSpuYD8l9WI7XigTnvGWeuCisEGv1LVGP4F+7TCYzESC
zSZ0n4nJfz//SBCd/gav3eqmeez84ktXHIfNf2HxDWmVhXM9HyTbsJPuo8s9Qtsw
hml3ux/PQk6V9sUzW8f4y64Let/q/+oDdsap1j/RxkL55QNp5HX8NsUj87xjgV4G
jNvPhqTCWoY4vGBDLhTiOSLoXrVgulx5qfFkHc6YHFLbig8QFpUlDXysTOvE79ag
tFUO1uzitriGivQ4x7UQdrFbt0Il981yWRkQu9OIMVXdyl2VKV2Y2b7eB/3GYHkc
C/vLIHDVmp70/Dc0wYuuhkOFxHdsg5vngQgBVM99FMAw5lzLtIbt2j7yLpsicP/1
XZMRhh+2mwGscu1DA7hw2bTHaMf2VEgqcSUeHLON4kjHXlkZxAMIIum3Mwuqi5H1
c9lCjiAqk5jEHFH0BGmzBpYs1nvnEGzD0w47fTgnWDCLb+p1kVvVYZ6z0H7FBo/f
+hvVZ1lb69a/not2ePpGh4KvARD9UsWSav6pLEj13fiDv9/C6xCony+2Zr5BoJEf
aGEaNW+F9NallmjEwiLuusrNBYYyYWuOtNgCu+lVW/BelJ+EaizUpEeqGb2ZAUUA
eMxKvMhK4dHwh6I+lP7sUHfmIZGBuXmK+QCKiLu+pVYTArlZIAznpf1Yn/ZuuFJI
/wp3sYK6HImK8CtQZCrkHObSWtu/ZrKo4sAjL2FrHReEyDLYE+kfcUXundG6JCKq
gNnlzkcDKvjVcLEOK5OA8p0fPkJuVint4E/aSGR6WPxPr8Mvg48oX5A6H5Vqr0GQ
v2S3/gIrJKyni0jI0ayx2xVqX92qW9GbVUyom/ppIOjtFX6OU2nGuZUGg1OcDBQ1
ZcWoD8J8JtONPrwzfDsmAkFgaTaa09VM/1OdI39LZGU+WwqduSPfB6j4oBDkh8sI
pCVbhxkw09mNsqb4oGIvdTfyDi9w7F5cgjZse/fLxfqXrQyj4MGp0GGGck/9D1uL
i7S/SPlNUs4Y2PPKe7mS/gaV0CEEonuuTi5qCSZBJWO0IcqwAbjB5KadVIyh1xb6
zQc3v8EpjvhWa70LasOrRtl9PvXkRB/myLvMweK/y8/ckjrOG0gwWledZL47AbUH
GKNKul6uxVcNfxwcZFAKt8aTDiKL1zFb38cuHyavrdR756owxabAv0mVfoRjGQwM
dKWJztpQezgcw6AW1W217O+4AS2KbtjwcgbZmlxMM5C2t6ZzLDW3hz6Y7b4puJM+
307zbFSC7Xx1f1iSeoij9PSOon2octhgvQMT6/fNjeKdZ+WFU4ozDWZTPG5b2MiB
KFGCp5Q3XfS3GOqGO/ti17HipRHcpeCjMh1brnhmIe75g5L0jU4dCtGJBg7/5+RG
2cALAJexow3DPAMDIQ5O7hDIOWST1iDoHOffWmNPu1VMo3N76Muc1Rt7lt+/0eX4
2eOPsw6WK7paqTofG3H9irysojhq1OuXsrBv/C+j+jXZU+jkG3mpsAwUXVr+N18T
3QyvhAVM3s4xGFZ4GXsQh3+1RT8MIzsdbb92tYQJb2q3f6m1+T9I6loYw7djeGlt
V0Xzph0K+9uYTPwSvWe5ZoLSKU9IF23SNRuhzUBQYn3Kmd10BY0+SiUraXQemFK6
4YS0cCVE3QLBwP5IZr6VAVY6Pu/hK0RGNUROpjIgMt0+mY0uzwUjuCXZpwubUWRN
d7arzxeScZ63++uzKp/Ota7NF7N8sbsXfgVFjzqjjORHf5FeKp1GCrt/4uGXgh7G
CHFj8p6KwOn/zhFvlJan3D55xjozIQc/PZyS5pUiP4chgPDF7ehNCs4IfnLOKi5r
GjtDYenWhZKWxlsZs3fTiLTBLV3199IpnxkXEwBirnSxnvsVPSl0x9VXi04F7UN5
VP/LvQdUYedb8976am9I0kouEJNH8laFL02I9tBu+L7G4LMoL1uO8EJKXkNYolF4
zyPv7NdRt6txmF+VgMhCbVeA89W2aL/4ILyQepMhuEX0suMdOAqMgR600RP+wy4w
2QHtaX7+wyoZV/qdBSdS1jddYC1lCA5f+9UFi8Hg1+s/4bjpKjoWui7Hn33HtQqX
mrTIV8vqZ3WZGrGDTn4eQiskNnKy4NYEfK1iJy1RmKwC21sdQOSHT0+Qj5WTX4eW
xYA8tFUkzMWlT7SX6wTyFOu0PMZemXPfTWLYDaXBJYZUVz1LVaKUmO8Dflq5kzUM
FYcHE2l/B8E6FTuXPwaetkEb/U6PD6qCL6XL0VP3eAnNVKb4lqJROqWbsSS46+uU
qIXxQY5vKZb5z+lyDVnLD5rCTvoiBsdnPHqbry+HsnDPe+zxWtsFcGmD4+j97CSu
/WKzs9rBfPAqJf4S76HDDnoHLCfHT611Xc0jKM584nCvW7HTV/Xtdt9DOrBsVTQf
3Otm2vokBkB31SBiu6WmpX/PcM6dSysAW08S3QLfl7nFpbI/cG7BKSE3dCgm0wmM
6U6qR0wM50tS7Q9x2kXiLoB0/bVLXOuZNPbRfbOrFtos1bmeQwM9HcN+qCQCZ1hD
TjsKC/oCJEF3Bt3t+Poc09TvpRy7/XwFZgpj8YDRRy0dA2EcyosUJaHCfaaQkpIO
M6THDRzpVSN4z8l3ORlI9zxIaZd6L5Cy45EIPUc1MPzkuUC2msU/Rsnib8bUN8dS
GmD4RDpq9yDucWePjb25bFPITUGOXgmfdw2puNv3v3KVuylBS4NXGrgINFmA1oYU
vaSoitM2kHLArstj5CQzV16ggJD+Cb5cP6jHwWROw5W9QiBx2ZOzUpRxFjGteB2p
ybLzWpN9qtYMO4/Qw/Ws8Y3M+FrG0gEzFUMJo9FPQ+lqKGR60w5ln4qtI4lbBDhL
vKNa2rVNS9ZFg6F++irILjMgZfQtq18Bab/KUlGAef2zOXFJeEQ9YX0PFOn9N6hO
/snZTL9H8OCL4zyH4/6433P+LvuRguCjMT6EN+MQjHl3jKTlJegNOHIT0QeZVPg0
FLGvwgMs+QwlGMBaMmUDVSLOFW7XSFhrS5DsjKR9sibjvtDcMFVROO/tvB47/CY+
DnKCv6CGrkqJr1GAOqDUI0Bi72NrTw4KKW2V+Wlc6bkjBn94jX8/IPJF4+aUDjFo
z+Q0+S5PRdme8jtxMvXUOlg6Xw0E5PFu5K8X0tt5C7eZxorfQSLTqVdtYcggr+JJ
qlPwfHTb3X4LhtkSeiC+cZLBE9UIcz0FVGWjugsnS4/rU8PQH2NaUanfY+G1Iurt
1M0s4COcZRyO8HPz0Q1OYvMzbUbQ19/DBI/JoeT/vGXK5VcFF04uM/JQjwWoO+Jw
4hpKVJCsVw+/St3uueLIvMN/nKKwMy7weZDWGEI0fuea1Ju1GKRlI/Zy/8udHPou
qK5mi9lsF8FEIjY8jBfiYONYHSom2Y7AEPjnrQC00SJNAv86L6/YnJsmvztfa4/9
cH9l7qbiF0qMuMj02oqvnskGIHO+Z+5u1WF9jL5EFtR5DhXIz2U6mQ+Sx1LSnSit
uKrzPAkfKiUKnSFc8O/5Uoz96OFwBBQB0QIRAkYscr2SJx3ZqwB43KPSssYQFUkE
PArlFupTH6aMN4O1q1YOQW5UACBw+5QYHBplgz3Qz1ou55ipRL9XgzpRe6b2BFmE
HYVnjCFBkh5yTQh27+R4d046auMP4LypoYGsEVs1bPlmrS2aL3dJzoH8VHqKXov5
lJlkNSgZ/hpIZ9081qvRKqOVbpJdewvdW7MVEAwXhVdayAR1WUgNtLylKhUmuKFi
7YKlvKr13LGbBBaiMgayMagd/+6klLcWc9G5nCyOai6KnUtJsQ3PcU7xCp1PaefC
EMEM579zFtsXy9ZWL1cXLJhGgbgZuLpRMmVk6oufqssTCPhxGYOrfRGOjqjHpEyC
I/0z6X27b2wlvxB62KXY+NC9EIOMN2O7FRs6gAhKaAdRyYmdHyD2y+X8CykVFjOw
RPwLgonJ5EC2v0sHV6hZhZmAPt08dETch7AjArGaUnAb1SJ/zEFCXhuHcl2ix+0d
AYrn8KmwvOLch0Edqb7KW/nWzlv1drBIp9PeqHKQjzGPZSKNoBBtm/bVM3/h141l
jReQG76Hiyg2BzDyOOGRgJGrX6zhceXEUJs5ltmyfR1R+QRvuB7FeffN2eLLQgiG
VNT4PN5it8s7GYjSlZ4StmLj6Dleh60YXRKckuNY2idIrTxGXJF9INesbBmqL4gG
SnUvBNh3323af7gvZNbumAcyiBLpB43kQwe+p7cDrEyaGvuuR6VA3sIp1mz97S+a
bP7lhgSNSazDBw1TaNjxx62cnzj3ilV0xBB84ilRmQnQQUyGeqImwBJoALXOc6vv
2fQHtmA4pWgIbTpBhDa2/q5XAMMa5dgghAbKRORXGeKkTBKY8TSHkuDkzK4h9d2R
OXDc0xUQxymnUvbNgWweujJLZY0rYO2OWVHytryZHq2Yjl6sBCy4UGmgDzRs5J4Q
o/lDDLL6rlCaiwFVEgfPmhGnCVUjLBuo7/zzMvkIoYVa/RyDshzkGsZNypunZPbC
cT1K1tqH5Ft40IKGZpaYxA86/v3hqeXSpMUZ/wTqkM4rHMoZKdta0hWIJA6/KTSX
lLq5b2Tz0Gmfi1MwEk1jLOgE5mUXdNmr+cv4uwSVa4e5jaRe+nB48maMZYuczEkV
7ZvFXs6UcxghPH9/WSnzIuHi64opyFMnlfWd/z07QUe432xdnY4iowrBpsoxD62h
PYaU4RLdf/oZF9uBsDXDQWwCHnDBhlpQn1l6A1f9MOCbZDhzsuvCzZI25XTYfP/q
clUL0K58yeLB9eMmr7zRaKnzoWbzsStTomuh4ZFs/2hDxQB+rOgUmzdJJN6K6uM4
tD869fMhsFbodbQcrkg7/o71XWz2XW1rHovQXc+W4mt1ydcNT1q8T8YyR49SAtdS
B/6fyXjkz9BVBPKCrmfzIKJqXt18egpQJK1XgiVsVAsWnZxA9QLre3yUyRCTbrUg
kcZLY0KCFexPFoD5CU56MbBacBnewGKDLz8Y9KTeCgH7JHBKVtWdyTeeb5KIcejA
I2e+3bmRSXlsD8BEDIhpR3VfoKTejphTGDyA3gDYUK/nVKCSpJrxTG7z6l+gELpp
PVajm18AhUkgCmm337TRqxpvNgVjuuaFHaNV5QSbsrHkIXI05Pd/akFBUCZwv6gL
LNIFNCaaksMJ3ZR9CdEOampWYwg+L7TDDaI6AsHJms25LXme15ky/DAp6pkGqxBx
iSxJ8tkRwqZo07V/KIWNu24WwMs2ageQZ+5fNWgLN6DlOJ4iujSu4Oza6+ap3Hkt
7KfirwRNt2CB9nR/pWYtLBxixlQuR7gbp65K1quaKZIlflqZi0FiAV1P1bcFTJtg
ty8QXokaVPJcGZRtLl3iy5JSch2ofj3AT1vgNicTLadBXzDq7wRemewRRwkW8NFg
YSUvudkWU+jy+WlXDsGtEBW224dlro+ZMCHOvTcnNoRwxWz8xb1oQzwubNYD+Ktx
igK8TCnDMW5RnLoxyRjwhpktZdsY9vXEp6wqQMK2vN7Kvd+cyhWDBXqXKjVFvFph
ADJJpRYZmDpxm4Gwxw267s0Im0v76F9keli5Aj+2ekkbUEM0FdzTF8aNroA/xoft
yI3ICr55OhThxb0PFgz52S3lswnOcD9q0BMD/rULXFkL93+SdOGaPl0ss6YPnJXr
m22ti5vXm3MdrhJ22luCwLvd7vq5wG7duLltRRQa7rwqSVde8dcAc4u0JbJ5Nv65
93GK4jjD+CaAcqQZlpPeQmGtQFYJS1RKXxNakSxHrTA4FoUsTGCrPWj5QrVrTb/4
UCJKt9MX0z18pxbPX3Vx5Tk4HA31E05QgdP7kitr88F2Mr825LyepDDG797Cr5LP
WQ7Vr7s+3zs6oYHYqMZFhCbx+XYRwB0jz+K81sGZY1bge8ZbU5JmPdCB3B7j9hcD
Eg/e21f612RPaty10l9rv8oMDWVaz4eFypzKV3ceYpCnfwQRrH1n7hAUxHGhKK/2
yczXP5/5N07Zmz8Ak5NMzVdd3CflmVaK1fcLTR4M2TharNqUKIJziH/37a75SmbW
nC2e+ymfIIEhAlNpsnYeltVUK/SfaBljRlMoa+EngR0Cj4JselNkKTkvI0o3VOVO
jGubpQNFXHiiN/V0f3y31Z/IUYdhrP10X0/w+xajUEmXkxEnBC4tOvEolx2xsUzM
66aadN33mploAYUGs7Ha4/CpWxrsgoG4i31P4mBB2YFT0qWWOBlVfL0oEOvRya39
jajfcFPYj4jnh36xyRpSaiCPsW1VxQE4dL3sp3jKZ/Vq9efLpHBRXmdpsMMX/TmA
YxCNhCm9kGMn8nAKEuB7yKiGeVpeExNdhXXamxT61wnlaM3qF0Mu8+bKb55bOdgv
Oq34Dcnc4GU14X+7TI0upwqlPc3dPQwVrDcjpjWDdv0T4p9OFIFoWxKjdQXIRpUv
UYNUyK42kLI1ly3Q//7Nf9Y/5mqTA2QlEeG2CtZrDtzd8kjda/yEOIvuQmum0Yun
PMN3WydvN/9J5aP9GQAucOc4KZdzK4/GADt8yLXjQOIm0mr7P5/QrObY58P5rBys
yyNGk2POkyDrwOttdS0baJ/onwgEZXe3w3cp+cb6Z5JdSBXmUlIQYGxLw60TLOm5
FTexMIfnZCBsDg8RzSZkwsG+u3+uNDWRauEuWfZB98ErvwujNi5D7Xcjox5RnFwj
t8bKKkwPuG63V3NQNXFrDPWGKfCtDENggOXrVAzW02gcV5Qv0X6z7p1A1m+ORuZq
ZMZS2mfbmLTfiRM3u4tBeaqoc6b+3UY4n52ebuUL/vr4ju4dMvnl7O0GD6V2P1lq
/Vw9g3jLRkltolh1dsJqoE69GoFdOiu7nOiYia8GDefefbl3fh3f/1um0nmXPYnx
9sCsY1oW7mCsQzuG3DxsPbACxrjS4BEkzTKCSPrAonP2DLKuH8ZdYfjLdIzrxEbu
4PF4J70BLt00heegmPgqmvQw7NwNbiQnIZJ6eEtcgZAqnthMwPtodoTslUmsLExK
aykAKljaq388vVmxJ9GoJNy6SjG0S4s75egFP8u7F75icbZCx+bMiD5Jc0Rw9M+R
cq7/X0oD3sXZ56e5MQk0M06VJ3CUA7vBehBxy3Fig2UGdgePc3LM/zZHhp5LlyJH
AK2/kY/E0NVErdrDVVMkm6i82waF8t2FCS/tfYkIe/UagQzcjREKMp9P8R9wqj2E
yg5S0Ek6LAkuuYGOmVdFCN+MOiK81PEmGZEYUZCXb9AfJTgNUBdPmIexa8c7ptFh
VxOcQqInHt0DkqxDx3vWzKx/opFtb5+EdB9ITH3XHbBjrZxsn68e9l4jHDniaEqL
pNJBip4QWMtgKtocgBwddG54eWjIeYDtS5GhR0C/WBFOvaghCvGBbiwTIiRWLDoI
2enwz+HS4e8DYqeurvaaWygGHXyYPg6FPerQJrsS6OoK66vab4qcxlxBBzAEQy0m
DUeQkfIgy0WjHp04cpUoqd1UR8UURrDx2qi6Y3NKyW2SQ1LTv1x7pUPmhx8zA7bg
8Z3y9ki+BMbty4aUL//iUe3DmhDVtU60pQNjB1QkhDxYuD0lD6Yt/2yrvpJmEyWS
caN1VF3OvkUmbKMmvgUSzNz8VG/8NSXsnxQKeUNDeVkZn1ZTjuFW2OxgnhJJHvI4
reKVAcE05649b5BNZgqvOANtiZ3x/k0OwwNIr4ZEyvpuN1EXp48HwIZ4nX929m7W
7hYBebZ8tGaXylXVbGdwC/swyLyIaaCOuDAnDYheB1bJyJlAdc/ILlnYBRgXZOK9
404YsUvBM9mphMem3dzQdFvyqdWCBpLVXghTQONNh40ukzTLVI0u/8IrzjijmCqA
STYraOeRVSH6SoAvltVun3D+Vw+RzAYL8vIAhhVX/lZe5W3l8IUMSZzGjBJiR2vY
3ntQ3DjS07SmfZ/TxTnr0JvypXS3JWKsqMwc5zBGseUxmriSQ62bhe9EBOm+2qR2
YrRMhGHfg+yVqGUjCvuiwjoDui9U62YOgtNXTy6U+TvfMknOYYvZ9j/m3Ral4hmG
QfvUG8i7AgiVowupu2rKboey0y0peX8PZfFPDpaA5H4YgUr/AdAnU0TDn2GFSHsD
3VM2Hjh8AOb/19NN7UzbpKI5NDyXvLJLfAvVTcUe6T6dvLgk1LWrRPV0Nekza8y6
I0p4iFN9ksnxHXH0WPmbz4zJOkonFgWcTTqfnM/02dzBsshyFg9pf41BAA1ZOVkk
m/q3vee6uC/14/BwMF+AV+r84wKdnm72Igf6QuFr+Q6lc5EUy5eu8RJTR3zP/G3I
BjCsfavf7Iczb6eheX94EqHyVx/3+XUE5+qHQioAzuWt8uoCRtElgsw/f+ISCKa0
O6i3BL3HblGYhObmVq7fQILUBIJyKnmOG5M6EUSp6zWJ57M+UiHqZCyppYxtM7b9
LYcFUpd7uGDHzXTQbAynl/SyJ18rqC2LrKQ9YhruUF+ZSF0olijH0Sg0DUaYDLs+
NVBBKagZwFauD1Uzwkz5s0IBZRK2E9sPzVwx5UxpbKuZwvrxTZKRa8SdkqTh/abK
zNHr3KTNtx19LcnAFdgAo3zkjwu6BrsdZgE4NtPPwfuRAkoMGonhaRILSmJ5fmnt
flTzxPpSZQZVW6LBX879izNeo7D/Upa2cLHTsDqr1b1ojl86qFUv7c+VNCTV21RU
1ItBrBVLpoKzwZpkb30hM+Hv+duI0/GYlS/MDGkws2j8XHVoLmWqradcrY4Fvk9s
rNSS6tm1fgzcnTqib3I1k8ryrx8EwRz3Q2N+Fa/Eq2lQmx7jOlJYd4dq1uuhWnac
3HNJvvkQTMDdA0RklQOIlFvzPmxvxF4InPGRHI33kEs0Y1qoU7sg5wmhDLk8DbPw
CsNOnymqNsaAUe1uXUiePgFS+bVqjJKA0cFGXg4z5X6UWTfUZif9e5NvpG9JgnVT
BSPLBoluGPAB24INCKd1q0MTSirM/sk1Ro1BCzaEP/nu6tdLEf30YUBw+doR56mU
CkMO0KVc/6k5Mxj9KFkRaICyMUS986nk/L3S5hJRkJJWb8OveLN0MK2qptazK4GR
zeZUj+yLTEAiUrbZOc/XrxcrS2/ZdVsWEsPJPASTygKEVUgJjGIsnDDQ29BUMiiN
WrL/q+AfH0j7lPbHkt4e6TYmN96wcQWThAq6LVMCGL8HEmdrmqaX8oyphJqlVAWt
ZTiS5HgoNJm0kfEidkZSagEgtHijtblO/tuzsa0Qbg/wZYT187Qx2ffATT1+dg8C
2Ye6bzEwFyxyRQduu3VSrEYF9yAoaf2vmD6xE9NWYQbfu6IgoZQTWIqcocc7nVoI
cxruD95gD3qYsceD/Q6NIx8nWf4FkUHjAAAuwFuC/CMnImhj/CdYVD9OyK5Wu2CI
Vp428gcx/k4o4wspI9R4R3Gc5At+9R39LA8HJy49oC3lx/j3OKsv9nNAljGBlI6+
/juo9kh5LYJAAOVyIQg1R6f/zvjEZnFXvobtIEcLdLB6Wu+wFpF/PZa/QoVLdQBO
OfbIoRzDd3WqZBY3SfRlidU0fMVlhOY5WPDw1Aelqrezmv5CKRPJB+lHrLiGc4f8
XWQE80p5jIv531b5YG7YfnwF+TraNN2YTN8Fmefol59eYurF2ZeQxlv830lVgbzj
FR2DOy+umdqDqvrK32aVpDsfQ6E58gi3RZFuUtv2HstLOxOpThkbXIXpqZF9NOi1
zKWCYQHLjL3I38YMEnB32RU82Pxfmol/UQctYZ2UWPaN5H+9qsTm4/fU28OKI6QA
1yTQ7jwO4j20dGUzs/VG675xOxmzIS+KD7cLDdD+QNaXVNgCK8gt2/RCdrTeBpWk
ulcV34crvQo7HyzysQWbjgVEHDo8ZNVGKPzwEUAHDyJX+Y/Kls/l2xO4SVTPc57U
qzHFDtbMJAX1vK2L6upPYQ2wp/598dcmzQ2wbTtCrSwXxy1k+Cw4z1ZDKBzNhZqE
OFY+RSMEJ0nM7MGHW+1fgpqBv3li6aa4LTitEh4sfvbHAP7YntDUYTNj/k7jrME8
yADFNi6NXNxxu4hTKCIZoleCSeDrBqqEmqXCtF+hPOSLtB5u2SncKTXF2KOH5Nyb
aXqj5qInSQLVcRa7J77SOp3Ca36RLUifs+9Kt17l6nIj5XGUnRnQxGmQJcBL5Q1u
nIY6xyfrx7pmuOyLdALOEQvmof7csJ1vJOKASPBhxogt3kPC0x4W8UFU4UQXGTXj
QLV0Ir6jkRe9HU5ZEAwtmbBUZhkWvX8zooZwXa09jxpd7RRuYwJIO3ZJ1bLWTd9l
zjZRftPP6SopC4E8d/q9HxRWyrWtbHJuNOOpNMK1ZrpyvciYeTZ0SCjOH+eny3ve
5V+b0AuB6XSqTMFm6rEYPh1rfKDfrt61VoM9Zbz8uIP3UOeieUw8JnpGVn7G7bUz
26U216TrAXuVS5cx8I0Q6HGoaWC9mvwSCjayDpt+OYdDfcOADaPi/WV3SRACu9Ff
fQNp7lA5HPaigirn6ZJEvHzHAL5fyt5SoVoVWYZaf8Y9iofGV/Wiu5QOR5Ll5tA5
G+a5UiPLF6IKMsOUtWswopTKHyaBEkI1S4QtPxb+nBvhbBmYpvmRp3/CjyxzwSY8
QeH1t10sBT6xl4YaGtv5beJHpbuj2hloFJzwSho8X2WSdDxKO7AWO64M6nu3mG/A
HABkfd8U/9PmGrLll6cwRfO8tOcu3+apmrvadqgpSsmwb91ii6bBkowzd17+un/k
J8jOoSyxK0qg8GAIgi7t8nXeAxESzFItSO5EhMjwuyDuTdqnLkgvB4nNv9rhvq2w
WqeL4GY4cXn4nxp2i91Hf30B9xXKl9dcI2EXhxN+HqTzckWwIsrDDlU6Wa37TiFI
Xi5FXzNsx3BW9y55MEtqc4UgR+lhiBVbSNI5ZN3TjxxG3rCEG5dPUApDSIS08Jx+
XPxWAnpoQrpT/Bra9n0a+ckr0J3Cf2ee+DYqZZuTF5h99TGghMzfbBs8KIDPrkQl
SYXzNCOdicQkGM6WQIwgzQRNXBcJaLdL+Bc93Qvb3D28t+PRf8dvzhHoBFdcxdtU
FwzPebS6D/ed0hE7XGvi341pRql40P2henGZjO51P3pnUPkhYMOWP0veHNdMdtxN
XpU6C3Hsg+P11Y9lpEgfVGTWLOLqkQoEaP5zfO9G7Jj4KGS3CvSwoi9E1S+oiTKL
mos9xBDSvGNqDdLehpBufYmTs5v0A9NEjvShHd10EM+Sq3kvyC3UJfvVn11AragZ
sKjetcYsMZjaJXV2nLl7Jdq4tlJgLqBpN+ssw9L++XsekyoCOpvDrCpuKkcqnkxy
SK13q1ZUlbDzxzXEdJuJ63Cb97q5WLbcJnxbVL6NRugk14ne6076Rkw/dy/UQTpt
/pjkWmDhopUeTKXxXiYwTVahD7zXJq6O7Yp6gUV3+msUtRy5oK1SE6FTfIcMxHQ/
xJbKMSmL1dXmqVgxHsGyTOKNtMSDLw98xLt6aJsIcIRFA2PLKF65H16eJW7TkKDm
gtcuj0uNjcZGCZ5znt1NKgifixYWmq5hqptPIJR7UIqEU3RmHQ7o/MWOqof2ELs3
B6ahx7OKhzKwflIp6Zoq9g/N8daq3RnHCmwWIf4JgPSmMVNR3IraaIll4YgOY8sr
J1gBQCkQPm/Q2K6Xkg7LZepiROfUzvVc8RpSlMFCtR/vHIkTkA4nM63FPW2y4GAo
rbSDExHpe1kira3oZsizlMe49GRuCG3cRiuaStKQFocuzFxNAfu1hi06orV0p0ND
PEHsyJ9TrS3jWE2dDTlySZRd3XpGNLxgHRQ78NWE2yfxiDBA3gHqTmkFHMDh1bjH
8NLqVV4R4Gkek91iE6+p2oqN7stsWDz9CKlbr+AskcW5F451LaMMd9EP6Qq56rYZ
PC5Zu1x2Ad5Q3A/TSjoXQwfJmaMmlqNrJ0rELuQfaARSfzYgtPaa2ATawrrEwFZg
0t0qvWzKGMPBztqSijINK1euT9+1V5gTcXR75wqhFpcQiLYa7RhmjnbPjPs5zz/I
Yoqo7VowTUUNpzP7UGgLpj4e3smKl2b4rlDCtg2bFo9GjSKB6iiWfX+y0bInipcm
hf9sb7fvABJ2aBVZ4dXtl+XVd11XhIWlZkga6NgsTlqLs5XNdSxEC5cpHP3c+vJn
J/G/W4Prilaoqi+nHky0IcnT8DHugW0Wln3v9p5bx6v26CiW8dnnBh5alQZq/8bl
wza2ZrvoRovqPySnsQJJ8SGhLYNOXyKTYxs0NP3L1nbkoLWKO7Av6moXialMhlRf
PNpC/1qlbimV/7oDrfcSIEqbt6GC2wMdxhRlV2hNNletwVl+VD9OaQZMQOhxzUkO
m5YxbtRdZXmQ7n6insYdIIiRQ3Zt2rO1aUmA/ujT7XxfUSr8xnr3y71GfD0Sx+01
8472SUBLPHXYK/5p1748USoVZgrU1Vq6QP0pHt9aZgkt+EwL2ESwenvVaJrVCP4p
F2sKjpfsK8ut8qSUA6ekxnqhbeEEJA7og4fzieJPGlAXRreMd2pOSoR7b/ibQbCZ
ZAIk7ADgZlezF7TlDlHL1hlQQi3dt2cAvJeiFKtDUyPC6Z7tQLg7TxBxKPukyZdD
xAZaFLymPmv+yVVP8mMJTDw0PhYlK3iX8rlsTYW7gBSE8sr+x6y5pSPNHUdGZzLz
nGb4Ym85C2TCijYbvwmHDYjsddhvUMlKpe87D7/50ucJEJWGKw+7FGDHrRU6bb5X
utuwNjA/BuRaK6CMKdtB7deXR+8tXWkfFgmniopsdy6Kx1yVKdDqsfBN8+wcjvKl
Rk/DetRtrmB623/s0R6Yu7NUgmQzsQNybLDZANFBMUxZnysKyzqASuqh8FVpmQyd
A7NJFSStxlzwAyeRAwUoPSzmOAtWaGQDNyPcoKNIaeMBuzs/PvagPxbyZFrH4A4y
Lp1jln5M5dhF1//7nTKd3cPXJTgTrO97KMgDpk0OSCZ7943b8YIZti+ZNjABwg5X
NHVF8KMis0q+MONTPcxdlY5Eu08Ol8/SGSVoF0bu+dd3rt90qkfnk1C46bYMelRX
WICTb0zIKZqIh1t3FnmuAVeu0yi25jZInjVOj/0Ku4EP40KBo8V5sy7bAlNsb5Wu
HxU+6tayeLH56v0bOlA9sejv6x+erUPEFG/RyPBsWXo/rzkf0MAKbgsW/UTIJ2Ju
g9icBb6yAK+pFPLkk+W4rGvU+n6CAKW/BT9dEKrCqkFZ5+TlIqRnC23LwX1C+FF/
Bc2kLytOCsoNy1cheqcFioeLCwmeVTntX4ocIJHDkoKKctrXd/4TK6L7gY4bbjBo
hMDXKSGNp4sM0DByTl0Tuhw4O6nvCLER0RYUogteG92NTJSzG87DI38HoVvAw0/W
L54p3DG/jju12V8ZGTObJjOlsHA9U7CN4Tl8xjlRxUOKvPQdpDTRaesFJUacEBIJ
d6heFVVHthvVGrBkH5nLgOWD2Wrms4Prb4cZWzt7iETe3/b+5oVz3zj0Nldub9Xv
o52YjByvW32putdutR6hTYscwenN7wwrfmuA32gOh9zlVQYx4fB1w8HDXHIBjnsN
CiJZrh4ZhyaHmQzD51UgV3yfa9ePlTUWkHDb/2+N8FiWfzhdmdHQp1uM58stTJqH
mJCJTewjEU/2n915CvM3rlYlERdVnT/qGDiTP/HoMFDdDwHVjA0BW36g5erFmsiG
LcITtvK/T2jifPg5NDjrxXts2jLy2gzR3ocV3vMicRlevkpBmYOh17LQbyoDTTZB
3LIiiiIBTWW1oekPTxdoDZkFIpJMRajhc9Mtp5FvAgV7tjMLNdYiuviPkYnGpNhT
jq/JwoY4zsytSMI2mrnDEIAsTfIgNxn3neYvIJ06TLLeQ8os5Lubvf/5+AJBHxqX
+SbhMotTF0/9z9v+Jdedg9EBVwOxj5e8KQMQ3BipPnU9bqTWXXn+tBN8FwpUn1Bg
giICG3k9MyWJdsPYgrNo9qYwrRKOieVA1Nt3vzKBtcukU0dqBeBm8rPSaLt9/l9i
eDeadraOgoZM47beqHz9PoK0h+SnTzK0QhMd1rSYyUwxIX/UdPkoP2/6eS47GmI/
ydUmbRVaf24MbNE0kvNXSkhgxPAI1nEjkBxUBrZiLntnWKTD4xBLx4SiDspQRoqg
qGBtp8iX17Xq602VFqDsKCVSY7HA1xJraycFxf2GGUHjpc51lQ8iyf/nUvT+5iVw
RQTHfE2avG2mPjMgmzMv7FWcTu3pMW2ycvv8t9eHCtwhnqmeNzO7ly8/7RXW64qM
QihIQr4JaolzIVei2qeqjGnfe8Z5eygdNP3xccSldeotSQdg8mDgaHA7gjwasiMO
FDjOSnMIOHz+wiCPgAC29VJ+qOOolT5US32b/2K/LqYKKq3Mz7DB8bhxHpLP9l1y
SLGB9FINVsfW5iuk2Tjq4yxQrgkf0wSD6810qZOi7Zrk6C2rAKzWxFGDmNPeodvN
KwgJvKI4pvHxb/LH8HD0tq7VwVKcpsaqHMEHmlK0acA3epCZB88ZJnwnPE0+c0/h
4N2dOhg5czS3acKPR5ivPapWd5pAYpt2xupm3JRJXF8gRKVZM0WfrJTvPh5Af5Bh
COBQJDbN9r7kU0rRDhrk8ubscViP8ZdwpMIphhnxVvncyB2vjK4+wB6EOxnOb5FS
cf2y/D2aqZFllOwdzgLjU7jRZOElIYf3c52ZJiYas3RHEFVh+cu+7cStliKVCWYO
ZHgVA7zcSok+FmddFSyUlEOjIrnR7/Yxk90JGzkfe9gW/ugpBg5Dge4VJ7MwZp7b
5rezn6uwd3Vo9FVQIEYnk1w6FrHGnYSMpv2T7l76IGAzvE0tYw/5Y7wEEDvVQXYp
09uOJgENcZECbDq+b/3kFJko85W0kfst5l1rMY+8BZ2RbEkUVwgM7ZsjTFJza+TS
NaGvYJ0HbdsQRnIpA/LFQNWx9gaknh2ocSgNz3C1BRP+QidaTwr6Xb5PErLupiys
279bm0k1BQe7CyNRaJcLJSWAx63Z3Or8sIv71rGuQgz1MZCEzBYQlPPK2a7oq88G
2LaW0Jp1ZEu46+DGgdv+8gliMaQNtSIHIB+qj2EnepOAsz51CRerDAVQ+YlOXiWd
pTxG5AI3Z/c291yU5Krj6PY0rhSFHXi8XKrbXhEHxv4mokkJQ1NGKG+m9KbrNXMk
pZ6hNeBjlsTzHOXBmELdjIfef+r4z39zP6uXpP6Xbb5zOwnB8Z7JZiFWYlh35ViX
fx9ZCYtYq9HsG7RWmM1yxBwh4symUJHiGKTA/r3pXv6+3axSBOqcwN0hylO5/snk
qsraUHHTbIDXIydCoIeSB1DAwcS0ey0f9TI2oEJz7WotuO9E6pQ8tj3XUrDTueog
euVsLD7BMneONW8saLj/qnLjRDIh1AhOTW35oFwmPq4++XbEyRW5qmB23F4bqh2D
8kYaOAdZNFh56EdKXCShNbue71zf+S/cCXPNqwvQOMtkAukmhg1/zE/K5SSpDazl
Kf3pMbUK8w44l/u+oSMeUt88qMIYCY5IZrTceg94/3KXxxxgi2rdk6+JUIknRA2t
xQJ9mM/IfP7aXqfL2smzZFTh3VdiZy9GGwfoxHucOAtSIkgmVMOQvqyDrDy+pCHZ
+PYx40ogZjC03jRKKxP/z7h5YDTmEZQciverxfr2x9ZOkC/f/GrTU3nw+fVOrBrV
9/w8o3PjCB/mDCVVODD+inDiJRAUkmEV5yQd/P8bMIsm2p2H5KXeqWzZ2GbeQjr9
AKhM18gIJ6+jh2ZRcqL3MPMG+yABCgb6D3mcVCiCtNAVOhGaWBxewSHqt+Py4Mp8
46QJXPBqtvREDzKboJy+aP3ot+28ZghuaF+Q/XXVPB/fhQHGOlEcvORu6G3q5nKi
Kk/687199jUsP2Fw4j48GMstL9w6aYs4nZnlnGIVTdauv56wZZ8S6q5dhz200c77
6auI3CtBtakefrmLA7P5vw+Bc3EZDmMhbPXYyfikIAUHfmMv6KOM7IvwEMuS790e
alGx1ck3eRW/lB3GdDUCdJAYikKmkOxf7St/u67JdNM97JxmmW1txz8COzEtWOsL
K97uzVy59VMCsEKJfSAQSsUqwCZE9uaZCjHMEZeaWGiaLTJWzrnz5cAA8E+eAXvC
7xTR8haBOhmiAtBMhxrI2rcG65l+TFogEc4YxhpCI0eL0r+YyTsQGMCPJ1ct/jQT
qX6rT2rTZqFV2PiiX9EEUVqp+Ukrt1MYFL2ufGAHpeNdHUs7nIBsZTu8AQhIVc8f
6xwVx+/g5Hf9uBr3pulxHIHHGSPIr+WtjriU3XLWqTvgs38vLcM/HH6qWe1Y0IZp
mcaD5/BpT5dO7nJRZtlsUIKjEGAxCN+yMuM6afLbl5okEnWJtgBQMzEHml19OhEo
u0ufzWvnj5qy64gufvM8XU6N5OaBC6U/htI2mRfGczsT1q+KdIQLyHmayIXqQs5U
3Bs9muy5EWoZr7gwtmK0JBqn2ShsFk3FOgCJr8dOkQMNNWF9RCua76EvRfurAjv2
jxFM+3hB5YL4vC+Oils4fp4CP0HKua6tkYd+kngSpQZxTuUbpeawWZtYaj0GoNI8
dJYSLtq7JFf4Nqu+qkrJCeZMFg0ahs2eWSETC+1Zk+jdy2hIrHE2k8Welz9+myPH
uTXADa5gCmuzJB2vdE15HErusXXLlHswusi19AE7drXm1u5e+lzDZAnwmYVpvDxI
EOhy4ukIa72xWRVNflE/G5qeu/aimJSvNT/ryuO8PaCi+yyKcjCworia2dXTzpDu
S4mnAjceW1kfUYt1d7uEuKP9WkMF83pDUXIyma/64e6021je6efakMf1yLwFjVLT
XqMaj22joncrzs4Gj4WISsCAnHB2K+HKWa72h9LodjUnawbXfbHxoq1aZPJIGJwc
GswY9Vh2JvoCmIceCdL/Xu9qFQx59auzF10wbq+NoIMQZPbEyaESJwc8lqRtve0A
8WfYt+L7M4k7OFXR5PrrX8NOlL2q1xv5OScxi0mQAcFsk5dlbdy4fWbKuvBK9iq/
5VFm6AXndp98iWwtD9wqOCaH/uYpAdlYZE0pu4XF7zTarDSy/38VdaRlg0QUJYfQ
Z7NJr8WsDRq25TwrQoDLFxWnx3EHT4EtGqYzPsPa1tfd+NaXQ1CWOveMpde2PkKQ
rXMOM+xCLhX25yn5OKOi9kEn7Pf2kcLPw7iHSKP1I8JH7kybGqthG+p0qhy7KVDl
0mnAv79kJVViGVdM+MeNeWFuqI0Bi6Mygrsfgpic7lT4eq1B9+bhIo/UYkH8wHmU
xtZoEY9MVbRZOUgDyFw3mHl6V+Q5Ri8YAjaATj/F6dY4D91niRKmiyVfqVwO7qGR
gmIBjY62z1g06TT3NAKwoxs0yibz7Bmj4blO74Gd/u6BKn3aeT7ckK9VulCruGxD
iTGvNJpGRxsVusXjfN5Ill3OBLETIe9iB3/rgVfe5wCKCfNb7FSPsz2mzyfcIs7J
KKGb8kXiSdnsQfe1iYPBrFFZMvuPDKYm7TRHY0dYq5KmkMWyIQVeU3Rh5FP0UDjc
MWOrJlLk5QzobW/f5m/I9BU61OD5vFftGAUlKQU7r0Ta/yO3Zz9MztKJ/lHksgDx
5gibXBcp98kpFiXwXA58D8wLoq10dnkeCQAJrWaQmoHz9dSCu5s4lzyl3J7RlyOT
lD8CBLxtSaGH6FDPcZTDIXiqMqlpVfX25xG1SPXyS+jzdLPdlh10MHVccH2UMG3/
Ni6L3NrzLN7BrMBzHVi5lI8Y3TsotIY6UipcHC/D08IX3tSmJGgzDhtEoh25mh9t
w3+bTDTrT+SKkG4Sfg5EvI9v7wmajjoR1SN55nXmBARIS6NeHBR+pBheJ2VUfZQ6
JMVini5VlSMPDNPqtqbKNOJ0hX9ZzjFgl8aSMf8uGiRHI5Jgeq8XzjXiFI65ZNKg
CI/fw54rO3ki9KD/8rw3EGlBfsh9gxXxoD8W6K9eYoY+8BoBHMQHpF9b2uxwsPOM
ttpWMZ1020Xuf1y5VDTUmpRdOaYwhWryLS2EfPdNyGne53aHemx5CwDLY2ePA8So
N0Bict4mus6lvb5mRNLmEcMg1x5+FrTRn2zWc/bnfjYfPp8EYqOueFgYtqgVPiwQ
ubpHx3n+I3Y6EcbWOF3uRKcPmNyCvQuv8K04i/8wFv4ohxaz6VlmumQteXzLDx0s
31oTZZoi9PhodytbUyJBVqFFE3xu/JVh+MWZqApioR1rnARGJoD2QUk7B8Lk51MV
mBS3ALP1KDoatwpXs4HAcYV1asIxei0zoG4XtpT8nzDAgB92+RokmslZ0PJ6ntW7
xCjX/cIylPazLkeYhklFemc/NwirLWq8xkC4pW8Rp+au8V+Bk/6LZyMDGO4U6tGr
rF33s6wOoHtTosn+NnxlqT9EAjvTgzQ02saGM96wHEBeg94eKIdS4A9tcClswVl0
W4z7UWpK9mXD3VDzo3xQLTvHTeZM379XA1nR1yqBieRcxFngWS54lx5Fgmpib7m0
Cbhxd1VqXtcu/zZ/KFch8oWfSwCD6yxTf39lGfB+7TbPvdKSYXnncW6IFah517pk
bu1rDLrRmf3On9e9ReA1Fkl+hXcmyZ0Zq3B/W3ChJoNu94Co8IuymW9HPlSL79tD
zdSlA15GQ7JyLP+2alnIUWplgulhCxBHXVMX9OqTQYlewg5uguMCfwb2hEAIKjfn
f6qII3mxQO0FxC9d5CoLcbAbS9PU4JlshdH9Uhj3XZiPAiGkuAviFJHV7zK5kZGE
wUBIXhgxBOfgl+FKm3SwiYwbmZkC9Y/hNJD3LCn20w0pQ1IiP2B0qetltYJFWnUA
G9NG6tDpKA3Za9h2VS/eBycE4FQOZQzOW6VVfZR4Ut1meQ1zaLq1SNiUhw4XhWyn
sbxyXftk1I4+989CQX9IVEzIE8rTn2o4t+DiVWUDalBeSk9FFaJJ9f0dJVoYoN7R
5xsd3IZ9U/kGbaF95LN73ZmasU5mkkDV7VMmQWlkuQxIYJemVHe7WpiJ14XoO6/2
I7HeWcBKuEbfXAZ6CiErhgxTtiPTSt4P3MSVT8jRWRFeh+rmz7UAo9088u4VN6Nb
mXccwLncaiWb8/FtyfN3cdiIdd710en6QH89SOB98VKzfAQ2ur0Ndnv/C+NIOe/L
tUx7HKWk/lm62O1FRed+Wy2Ax64UZvojNrD8VbtZrzdfV6ozGKSV5y2m9/nVE9ma
vi44lJ4ZTmt2/nf34Xpp4g4j4lSPREY6eY25XmRgteNhLtvRSXa9g+gOstJFgyGo
M60T2mr1WC8+vcbWnF+SCaV58kRnRaM+Nc/Qp9YImDaufaRHx6BTc3DmA8FXsk/b
MbBC6RVXwfYJ1IISg21xdC3VjY+6CRrQxt/E0G31x7VHxh/7p7plAUaCzFCDtmXW
61w8ZBJBsNhwUSp+SBBfI7zIp2aVj4KwPvp1NMipMIlApqQv8hsAP+naR4NTYIeW
Dui2WmQClFijyNtWoxgueERYSQMfIjLzHEGqV4bzG4XQ0gbULM+jGygPSTck2cSi
HJVeVdSI6Ea0+OpxFLHfubqPhaup+Z+32XEgvkolbpmFTWyFNaRXdIpn07MnoHTC
VdJRinLVaznFtGcTLez3sYmL904sKDVyAr0UyHbatYqVHfRNDquhDIVUvJl090B+
nmqd3WDbG22oqkkHx7wncw66D2iT6xtwTkgYpjtiZ2NQZNCxnncfZqnb5aUyA1L9
eVLJ3XZOFFkIPytMGo/i4JnndEZ+00c0DiPLGWm2/oKk6qC7ALBL9ujBosQYT3C+
9GLo50Ixvhn/HAVgihX/kT4kxmjOhxFozsShb3ZRO1BG7k1/gUjONKdHU7fXZjf5
+yBEdVQf12wblafXiZL3X5QIvwYhsdICl0L/95VedUvqQNxGtx79LEfRpbnLJojq
hutKzjLO6SwqPQxm8O1FfXh7USg6oO8rPkeKGvyYglyXcOFjXCuFCpVlZDshrQ3I
9/w0R9iOKHbWJcZeQmN811UTTujPxEgVDIz9C8AfD3kOJ1OppCKoREMQheGUfKM7
D1egJe2F1Sl5b4Zvce/fGUUXBYocyeuzSxcNGoj9/oMoFEWDSWarbP+70zEk+cMZ
IX5iZ2kgPi4UyO2f3jKC0k/OtnP6KvREYsDyLALEMypCwX5BmscS+992TfnJfz8j
ElL08mXqT5e1AF6b8BD/LX+7lFLS1UWWSOnzseWjF7J0ZO64oOSOVsyquj67lPTS
7ZCfu1r5rgsyrXub/+li66d20eJeZnoIE0OL/GjlstXI82V0LfoIElDhbir1/U/P
QVbhFIIrRLVstWytKuqT/7jlYTUSixWw55TMFR26cZd1puPaQkwosMMnQBRUHsQc
pRHAL+ldgTNMfrAQ5bEYzfFXb6ofOa93bn1iZHjUnPKUdUhNa+LI5JaZOYXw4pLE
bXpodeBRqHamdeMuxl4do9ZZJ01lIAthT/BU45Wm5h2oWbqxfvYcP/3wFSfv3oQR
msCd6ki9VGFKyNmoAEfeoQXVL6m5QEH/jheMtKKlkO2OAw8ylafPW7QKOb4fHJZV
NOm96Qz4oaOzjyNPyVFprf5xMRZjIG4v3r3Af25nzbys0VytDJljV5FitDQO0c3O
/aq0TgfZ/gYRgYD2cwNKo+OGxamnC0dU6ZAVSo5+tJxg/0W69zWISOHtAFb5KVWb
Sb/E+n1RHSHQnzpHiNxnD0mvaE4i8/zaOncY3dIq7KKgR6k2bt4ojl5EY0qZ2raw
kkO6/3aEj2agvljPf4mKIiKc4OzyqAa2KtNcp8XscRUglGVFtDP5HfS7jpAABTsi
fToLvZhrEzXvOZRLJthz9vK9hq+A9SQl8HXs6za5LM6xjWtfE6/24Z0zsCTVnWSE
kqTnB3iLZUj0M1gXs7CT8MQE/Hyak8f5jQH+d23U49gf2Isf9MW0AjDo2VuRrljM
W6LulqWAmQJFY8olyZG3SOWE+SAzI4i12/XoklROC37hd/Q6gGjkZHwJRI8Mz8Oz
N56EUbHD8Z6XKZQ86ACYqQrZL+KHUjUruFjvRcvTd3vR6dxb6bUa5Zu+rrWAJJY9
0PrgUxhG3l9B+KH5NBkPWXeAi9FWRDO/xwFfZHwbjd0N570CQ2kK+88g0CJW1vep
mFLmt1veFs8i4SHw09PYTJ6uZ+KFxC6hXwasP4fe2KNpF1N2dSqCMOnOXofDbDIR
kJE/sILkO7Qif1Tl0H92tglvJqhlC7FDdSKlIYX0UX7JBjJFrPWJRcCiIVwmGUZN
UnSxPcLmA0RDwV07yZBRmYGiAdttyo9vfRC1AU9yGWbLXBrvNm+JHS2bWKpZEuLU
lqkQQJc4vF4Xa/pQnh4+6FsC5Je4I7R9tP+Z8nH36x0oFdrIJOK2naOqG0RjjNoZ
uZosw3TYasYuisjkAA6lr5WYS7IpaBEUqQtXBQOM9TfFGOOHAJDBG9FIzWtWVOW/
4o1F27mKSYMgUGnPdOqbA+FmdOt9jaRJLCAwFX+FPzFHbd6vxSEA21USFvdwUvSf
31IKId0j/LKFUT1lBic5qZg9OTlvmmBW5xR/8pR2kXyVAAMsyQyZAN6Szpa3wkpS
CY6zpN8d02GUJ/d7m+PuWYZeKzLTyD2NTFI9zx3QLYmgQwWFnJzAgrDtvXxEER+k
AcKk9ZbbivYy+ZY+Ljs0vrTLrXaGXfVYJNRuIoB75Ux9mAjOD+OlUwfV665XxjDC
/J/1ya/yJiFLrsaCicVckKidbm+RTpy8OgjSYi5ZQyc/8doZ8cRxKlTwnMJd3SA1
PbOAKOEjExR5XMbeJSnjH9o8yBCeD+ykSC0I4um9jf0HUaDDs3QpS8Z6LkM2GpDF
fj1qfCVgvsGIqt02QbqoZVhGwpFzGoM0tHsfqScDpldXPqvfm8EWdX62E4sCHrIX
m6QG466Zmy6wZvNvUQkHHL+SVmTl67l07Tf6BmS5yS9neEh7jnR5pFhov71TuK1q
DHLriLuDI0GVm6izQ45F2/0XjgIWxFlMgtAHJ6kbd2h49N5mk0UZtARs3ZvTz3+2
J8ElRnmsuurMWbS9YqKvX40/SlOb9ZhOBYYI5UvOwpLD9tQnTHoA/MxzJ1yR+DXl
K1A0SiPNXT/TERQ9MHR6Ty8aJSE/Md8oM0YuieiIQvBHBX1ir2wpHieZAo93VxOM
WsOChUa8glS9sUZ0NJjAj97xmf2ZhxcW7j0Q+2zVN7qES4fIbGkm2y0FCca7vzRO
qeDRSrvZ4UfxJ+ZLq8Oa912hfH7h4vy5f5LemKEFNEJage/3CfiuEakRVi1uIvw3
+1gK8A4M3ci20SOD7UGJfXPBNRSsuLr5L3HW7OsQG4uTjqlJqYOvb2RI2S6JJPJ0
9XBMSPxfrJrlgxepSu5WKYOXP4zXNKpsjX/54408yOMYtiXXJ/GNgO74DtHzv67y
Ar1GY7UCvUrXmYCyeaRdQpe8u5+JhaUdFcjHMjc2l5grXyFSF2VQY2YS6GMG9Fyd
2bfnnXLbncv/Wb03MAxkHQddbOnstCTIg1pkevzHzaYEaYRVKTAIV4E2WyEkZOaP
pByKQCVzvv8i4PFB8wBs6tHPbGkDvtcrbyr8zOr5KCW9eSbdMUTSsH8UiicSAsLe
geqRb8qvhArWePjYs1EkGGvkc8eDLeqIs3m1kdyK+BaP/KA/bQm3RaymGTrkeg5E
iCG7FKU+Vhc5i/qy0iBOts8QhaOdZr+7dWor2vHT/lfdvpbxkjzQDD/n9nshkYNF
pvf/RdE72Xea0DtqXv6FsEN2h8p3spo2pFvtljkiEcNUVFBGYKPKitwaiZbh63UA
NqiB7bWeanIVNeGJS5C8bjPY2F2Aw4ENN1g4b8o5u83jlStg/Q5IhdLVVuy3g+xW
5O1RHahVmfqb5YP2AqCBttZJvcbQThuheBRg9eDjngPPz09j3CqHy3LTyl4/sGPf
9cB5Cl9PbvlFWdrIjp+i14BAcggGgB5kf5YKcQCbvNIPdX32SZ2F5e5dvudeqtEc
163qgyA/crHiKfrvL+49nhOTssReXPNqnXWSLciFJQ5pB9SgPYrJK241y5AhKZpa
FCYrwtZ4BG6mS/0pCAE29ry7/hA0zUSiGFBhYXlaHLLNXK73eLPFI4BiPW0cuN2B
aA4oRbEfEk1Cw6RvsOSWAyX+EOaUJo8t/UMwuraBDPLJSXqK4Ajp1MuVg4ZDdWfs
ZH5ibPfLt6eboaX+HxgsrxdWu+jvNoeCAmETndZnMsR8SgpW8mUKTBpGDmw7FwC+
5byIwpVkNR71AL8LtAHPC64jK/2JDtd6SgRn4is4oS6jidJr2o67vyynkbDSf/Y3
LleOZbmnczIB1KjyU3lqnB/sa63N0gEjRxUTFPKJ6ddGPIG8OLHzpuy85YFOIZBk
0D51IkbZS30AganjgtTOP0Dyobbs0yrkERfQRUlL0DzJOXuFlyX5922Rb/0oQT4X
tKei6nwK+LQmKxjvEyso/RkWCjQKTfFcZOts6QZ5hls7jviTuK7g6apE5fzmJTYt
+cw8fikOONNd3+GkUvPEcN+mCL+LACwfKu7elWcQukfdo7T3jNEFtTKTSaSRNriD
a7cMhzPa5zfJCi/MrLMixurDVe3nTO67kOSdJnTJIdkV9ddxKpd2y5M6qykGDXXC
hfbBTvqFoRIV2x2uArTXjAANmW0FX+iMOTcfFflmN/1IeHPYNd/ci5nC1uUqiX3O
9qGr3UOkHgQFBVhTwzAI4jPPLBu3/q0K81nzryFjPs5CiiujJEXH79yvKT0liWcH
H3WhCbqLNv9/ho6Oh/gdKiiPLUGbeL95P9Dk8YJn4lmujSedpCLZtUmdZzq7fCC8
DA0eneeshy4y5nhtkbywhry0mrJxHTTaTx3hIO/L7DzoTw3H3BfwAdVoX+FIBT19
H9RQgLjmCKy6kXeBeT8agcuN7vKzLmXwYNHx5RS0EiszbKPaFzCvG9gcOnO7kh1K
RopIFKU1v/mqkrm7PMH3fxSHpEUy03nYM2YtdEleuEoarvOT+qh0x6+r/sVE8qwU
mBKXdDOB9U3FeY+fG/rcyn91QME3JiCoSK58kmJbsTOsokVk4nMi6WHpptX76S/t
LdbLAWHBrNcTNa1p8MwcaLnDjVog0DSuAYT1XAcMcBhQbAmf4PmkLg1zqgeE33/P
1VjzSslWV0LdOD7I9yG71RB2bO4l0L8tia36p7PAt8hPRy/20NxLUnpZMmRKluSI
qzx6ZigDhujjzY5UvlK31+NwsfPIry+RjlMPOC13z7tfhy84tIqIPMi0XlJPWgyj
FKtVEE56FzHYrEvaznllWlpaFDWhcFIAvjimQ934J9d8GLFnAZwZHTiOSaX8rtyM
4O0tJmbfg2MTUr5woNbth7UspHxXCH0qGlaxsEG9q7xsDoT5gWiB9sCqUbC1GkbH
7dyzku4EoTiJqUmb3TKCVRFvWEiJTQVaYU70UJoysgyMguAnX5tl3qIZ50Bt2MBV
rHh8q7S5pcCbCCp0w2oUrfm3/ISxD6Hs6eY3N2fpK3DxmTaUw5H5NBlXrZdR0z7W
5fm29fr++tA/rX3+O1Jp+S3BoI2bImuIxi/X9SgAlze0n/cYuO/fkAnmjOnuaRlu
X33fEA7EUVNboYCWaAMQxXEyyZmhiCBmBNaSQe0hgfbYW4p8hiDOEv3ufovTjJwQ
8jOUmmmVs3tpMTPuHY7EXsOUbROm2OnUiEbRRjE8lOhQaZ8CcwrawRHxZHs/S3Be
5B1BZbDioN49Xq8GYb3XPBAESXDCftPUMBLzNCDLvS2s1dFz0ojGdf3qQyaefzLP
GvZsdktwvUrzGA1AUBdclkkkYHbTMkG94zwjJAlNKfMsF/xll7dYXYAsphimPZfI
H7g4IaB+BB4bXEMwYhTEzWtBdMnrX/JdcHf8xpzfD8CqGPZXKBUy+kczHdLpzZC+
TAi1JNUPaCf65h8MIWIY5iGTuoPtaibOkaXR5F/icqxINWNGSMpPaNO2YKJ1FbtV
7EH/rl2oSnhy6R538DjIFUK+/4zH64vtRme5UqSi4tRLmAGbNBiD7vImdKyDz/Xs
yQBIlTUmWERyArLdJ3pDepjWmkyJufLMmugIECdpVxNY2Idwcct+spUBQBDl7gaW
vB5+Zm1Yy/KXx3XMXR38i6Q6ytbkjRKkiV+1/b8skaV8wtX2LdEg9OPIukbjpw++
zkV0k04xcxi/n7Fn/Jim1nGhlZ0IcYdJvNKLgES7MtJoOWMh2wnvFDzGvCG2iDhp
1t481AGzgZtVJkrTrqpY6AqllJssn69pei0nIlC8SNAV6AxA1Y/z/MyDEfGDJfIG
BncJT2w83WdxM3NqwbkLkfXdYAnt2NwJI0x3RZUDCPG/5v+qVebK691UnH75Ls64
TiPSBbmOkLo8EXrufsbRmRtrqhoyFIZITve/XptulVO1FIe9Huxdew+RrFJiGqPk
Nyk1e2lHDHgpKdg5qmPURUceXwY3o+ckWzHiyC9eg+Y8ZRivcrwupVHVd6AOfoUp
EavdaxNAF49uGbXHziqa6hqbKyGTcEXNB4RuPHrZeuHpYrBTAEvKAmIm3gQ1c6Yk
toXb2Dg5teRxID6EUVhRIOaRiU84LsDAupdpf+/PCGnVhS+x3SYFfd4Rb59W7AUO
ckwu6oVw9NPIRJY1RQIVRsSRp15b1NslkK7E+hXfixCEOgnrbnlGqWrqB4oAUMBy
QWRfBKHpC0x2E/M/7p4cIe45xDcBuuLzOe63jEA6Bz6LdM6eUkIBEn9T+mKtbIXv
ce72F9Hq3u4hpEUuzshUDimpHse42mj6Taghj9tlCLtHLMfOYy2fxnAhDJaXvYWj
hcoWLi9VfjtDqbul8ERfkvAfMRDHM09USFoEKxgTcZEM7J8l+2sUV//TObCcroCE
R9Hr47T560IZ7btDr5i/Kd9T/KAye5qpmr5mJputXiQpdMMkfQZ/JUBiNW05W6e5
i7lv2Oy82+FMCYZDE7OQFrcmOGyyVE7pQDqzPthZyoI8W3Dtr132vayIjcW6uQJe
fKsH2pUQxJ35Wf4ScP2umWb0mKLGcxFMyLygHYNR9nPCuO0HvNpyuHr9Xt5By1xl
KsqzfHTETDN8D9c84eujG8lmNoCiF3KsjfSv0ATh4VgPSjAiLXNIF9qUBSKtO2Zn
nwRdDpbKfJMx2xw3mJbYEMk0oRdAhK81NE/S6ohQIWkL9GkVcjGrxxEYjVUWRHAf
DnDokFVrWLR+wQRIiNjA/tu8L5FXQMq2R8zeNaIMA5meubB/Hmoh1BhXdlFuliBI
xn/aPGq48ED/JFjL3redicovJDWdocTTQOZWJMTexAll7c108mllukaInqsogQxl
eNHCwZ1jwXkj6JxGprkptU51NQo4qDjg2lO3oCjIW2wpt31JKp4P58+g87Db+RnD
3PevibPLzwnpU+8tTvyCv0PNrl8T8YQgJDOM4T8qNQz5StLICOIqDCU+FT8BdlT8
X2qnSGglF9LT1qdTzDztE0BlQDt6Ks87pFyaecIYl9JszrJHQbmZ5OjeKip4bl98
SbBfX5y1lDkYdvsH0VLuveESq3g1eCD3Hkxf+P7bieJNB22dgsywRoZxpaBAdkGR
5xFRRTNd/ai565OmTISF6+M12AfUBI7KKWiLZsuuKDgB34xBf56uMZDgJXxKz98W
Y6zY8gaG3yx4F0LwlEeZvnd19L6qSo7qKZP4zJatt1l+baD60nTuNqeITpunBwZt
vLo+7dVe02nEgrgPqq5Mi1eRlxN3Exv0Y/Kw+KtVGn4RG6DvFCzyYKs3TnukkNj6
p3yXR6uTWh7h1skIqjekoKfk+AsrSklktklWx9guXlxp3y+cbN2oivn9kbprpdEr
Nftd4qC69D7KAVS7lbwQ2RTXiAqUISL6z78qyOsWTp35y+0vClUio6L0jfdLV8pY
hlTNKAjgo51usEfqPyl/iA0xvQwdoya2+a3TgY7j6MMGZ0kciHaVYniE0Boq1LWM
1AnPEx8qmcu6tV++c4M6BgjUhbiWooe93Sz0O3KQOfOX+sfcR7ASZioYZYdAojdV
B1oed6eVP2z1zU5uXwh4bv4XGxhrwu//ryn+F+rLx7HnTs1BjSYMpijAUwFTqO4q
heoVDVwgUkb+LU+FNTHOqiovjbgLPCtQ1EBWv+lMH2vcMUjMkvTNT07ojd9cGkPS
etKNtPPyzyuiJZYKFBe6kuxhp21Vg+UoAQciBZ7KvuI3ot9BGnjE71RmG+J6UFO0
xj5/2fv0OYIXAm+3zdFxpY4HbGOrbS5bfMmiuBR+w9rzgMyzWPzKcHnNJL/42xYd
bdMWoD3HMBLvnNFUrq+SEsrED/26Z3Nn4gSGqjfsmum9f4c1vYI3XpJk3u0Yhupd
7Quj4jjHM4zAsrN05Oz/LA175un7P1suyzpkzOsyzaa2fr5PX6/aRpb10KhOm0aL
6SQjb/8EbpxYq2artyur/v36HRDpAHixVRFl6ZyAK/SP/m2jwaw2uCOTDhn+uZ8J
w37FbJGzcDwmBphXSawXWZkzsd0/CyjRwof6mABxpvkM+yxZakeGmUFImr0SV3CY
CcvUCREsPfdrXVhwS7ydQjb1Dwv2gsvhXr+b5f0oG/Fnz5Bsp+wXrCIHhjKWtTlx
sQzCngF7EWJt05tbAtywNFbqH1Bnw43gHCNLE3OMJlLGkzGoTWzG4yb2TlV1XZLJ
uKMeJXIqQLRsyw67LJDGCD3pV53yuXWE1kevTVHzMUy7+AfMLeh6X82paguEvSp+
4Z7lchV+VC3ux+2EuoPfdv214lOjqJyj9SeOB7rAlfPphxelN+ukCUd7M13EKnYW
jpQdzj0as4GNtfJT/Ksdu8235RzZiYXnNmeoxC4tBjsVhu8UfcO+jlR+dbWg+GRi
pd85lEeV7+91o8RwfIFJbyk1IYXbHzB3s2P6tuhP7ldH+D9X3e5cjvDE4lxq5nJ8
NhLQz1fvthiAeZwLJEE9d6R9/BzUmVuWGVaM+H5C2aT+gvIkGmAYvTawRSHVvQTr
3Qm0O6m02lhbKaW54QX0GxHNBcTUAfVFz+cqr305JvUYwHBkQayF6zUITWEJ8+Pf
rcBJLb+m+E9nPsaP6vQewe4cseKJls7oBetddL3A2J6f0aPPKCOe/quD+nsvWoB9
1za0YU+SfnQvfUBSQVsDDz8SNxwNqJ+6laDGTZfaW7sqLVMHjXv5sPK7al3p5c8w
w6VTxkJNR/yQbfVU2MIGdP/n/dM5dDyUkWI8yY7pFXGLeeFd8gfH1o7ZlHgl9Z8m
oCGyPOJEfxSEHmWAeewtPNkx/qDk+nAGvvgySAmJd9uNNHkBC4dYftBXWT6/W91e
ti4UfQICnsZ+xwTS7CjonTHC5pwhf0JwxK0n4RXq3X/UeJK44gw21Uzc+EVL5Cw8
D6xPENfUSAqfSXWEiAjKp9B5JZKZq2F8BGqn/8y0s6NKzTjS+IaFKGTXcFjQ4v8Z
b33D1Z/gkMXaxYWjBt8tJtSYHv6zuydjFCtXSVVKrR/cqohjB9ZEsC4C3to/2VOx
E3eIRfEqQ2aZJNzuZP74JZJORd14CYqZXTAM0Pf9rlQUo3dAILoZ0Toa3Cbhhrfa
VIgl5rce0c0L/5cA250MSGjH1w4nBZnpkmhM4H6GoLu3DuCHYSrSA22Bu7jo4yqf
WN3CI6bTiS+dF2/A6jQgRMLevllxKVKQNqIBrfijcMMY4dUE10ZhEZYXoxsftpiy
XJuolX2cPJKD9nO3YfPLfuXHAEVcEzUL2Zr2iIvLpeE0dnNSwKG8X7nF/IRI6Bby
amHY5oJx5ZfUkD+7eZTTGqcynfCSAWFSHZjiWTEQXHAHqzEYDpNB3XzY8M6ii0y7
feP5VRUxY8/H9FHHE20f+lhkkAx51WrrpdvpfaaHLgGdGDDjL0LUJWYJkViKPq2m
TwBuw45rVPw1PCQOEyeJax6nUUK/G8uQxQsjk34YolZNrGCUK5w5UJKwJnqRefWR
ExuGgd4gkQxJQZAkl8NpHXAOlsDOJNi/gsqeN8PiO0GRq8KsZchC05UyFRP5GFBw
M8pSZ6+3/sB/EhwLTieTjflBLtLBragg5hHXASnBZsxordLbe/pz8Kex5QFdBIZX
yKpWj/hrY0C6BNd4jd1PHWAQztJvKRThrjkYjn2UKaEOL1xXxhEzDQWmB/qEhcl0
aTsCI/cDpYDuG3+8BTRe38wTVl7nWaB6c5ZORLnBxPy6deQWypsnszVzdzjDDYAR
dbW6ppS04EI2J9TRq6T3VyPM5bjGQ2LVNb/fw9s3ePu+Xs2PuFcSD84q5GdFhkom
lKAQVXwTbHnhr2qI96EmjGLluOnby+GBzTH7kPbqTIoOqQzLn3Om0YVLIW4BOxOK
Ac4P9bE5+VX7hqld67MSJa4AgSl3VsqCkt83hr4CYLXBnNR4CabBumYpeXeqAwoy
9JHRot/gPoYVqvHwCBV5cK/XXfGUUW8fsOUnb5uBwaRgV+zIZOR1wz3vrdOfnCAy
qJScGu3l5D3E+hBQwdvJQ2aHsEi8yrWU3hAZ/S2RdTYHLcqoTm2IETz7SXLEWxdw
jsQDvxZrcMAw7jLlhpqpibTigwgJS1JwERta5ZstWSDWBC7NJrfjAEwFRYbeArvD
s58E6YaNrkLfKfq284dNhTqFkyt/cbwEn5T+5MN9hyP2R+m0yr5OOk88+QQoN1dY
YEhw7wqHFsP4OiAwdQx19MmDwFx+S1I1wpVhs8UuwZrmFeQfuVpT2132z8y6jySI
fW6AxjjuENIyo0XWp/yMtk/DHJNvLEjDugh4TNdt56X5Ei/HHB1rYXPfLMPHosRF
/2l4jTDyW/JKAYvThT7hVm57IbSHPORs8kjt1TFLTlGQtllIvTMaQM00uGhg5Qvo
p/QFyXmiMo2RkNCkunyZEv6mou4zVLCn6T2WyYuEkTvRtPNjhaCP6cSzg8x3/CcO
e0Kj+VciYj5xOXyoTlyuW0vbl4zV5aTWva0+nE4afH8E25kLaL7ZxC5YSiW7NzCg
WUJ/JT0H6w39zhSXU5obVxJ42eCA1YK81OyMGrlP4VfTfQ/jZqRLhl5RvCy/zXm5
gZhWnfsnZfMwQT/7eQlL4r6T2hcVgczR3qrzNmcQP0yFpJEH8w9A1c7MFmxGACrY
Orj3n09+0MTjhZBza30kwJzsGntoTRAZrvbP6Wc+yYvK6YOVZfi0uQVO5RjJw1yp
evEcBfzqWreRSTW3zpMH4MnL2Gl4mbhz0DCVRSJ0ntp2aCG+3SlflzU4q3KWSUTk
M3o2IlnBsS/pz6CfbDA8feqlW7+LBO1V151cQ4AYoGzAYGdaLBLCqrsRnd3fuiBI
qWq0QkWO3jau7PWTQCgLX+ie30hKKy8kJGf9E6JsbHXIs2wLrfHsADE1OJ7cHcez
NkE5DozsGtyMU4SSGPxhfavbnJfR1rTKGwNQKoTywyKY+Yalc8kCKTQ4FA8dKemu
BsZC+hvOpHcxcxmG6NLpm17zO9V2Cmsn/4EbBEvUeixhq0PkxKopGky6NJQDLMYz
SNebmCpyKpNGkkYytCdA6+TAvZDg3Tic7RS2F3aRxXKf/TlGnB3ab+iQN/lHMF6M
3SLdQKcjQ+7gEnNSaKOQHmP99ZfSSTBTsA7tvXTiXR3DwHPg8uVFROk7+PKq3mHt
FoQAuBhUHOG4nwS0EGkP4JqcfUI6ow65jWPgTRMOS9SOp5KLgPhQexxeqCC6Qjdu
q88mcVX16JrJhvNpEfc3et2LI346xom5jja2e4LnNNXfTh1JmqYL747exGJQor75
TeinIxjDoMHs+EcgFYdE5JEJYaJtKNl3/jhoc4CP1DFu7q+pUbDBxYTwMxFte0Ye
SqLIGThToKMvjCIOKpFTmcZtkW/PfLYUG+QP4Bc4OD52tek7y7l143hgSO1YgVcW
Scy3lfWeYWAxArFXK9RGeioEq1DiLm1ZikeC0E0Lg3SOnPedqqBB9D+ED+a9mElE
tM6FPfgwJh3bzOZNY2YZDyUmXxG0BLVMKMNAr5p7oMne1/bg5zKKbQDvGoslSMBu
kolKDy4Iyhwe11RibOCl2Bch5ZJH5aXMDz6RqLXE/Zq8x83x0958+uVTD9vOzKeY
iNPNUMgPEiI2exB/9SIBOe+A046x4/Je/jahlaDf2n4bHcdLI/zN8LL6TPWc4NeM
bcAKqvlbqQWrMP/xMM+jz7ct15+jq7TCyn1M/HTceh42dH2eLfOjUvCjYUCIU36S
I0bhg5qZ+V3vCwHR7xRm9dhvzeehYNXiHaWl38vePAU8+HzetECnf7DYGSslzi5j
JYjrSIj8JO2JA0Y1vWfUJL/OHuFYVCqtlBT50JwvZriFhysKR7KQMJSTfr4GVXAo
7/HhaaTbilylPGfhsryqdZCDpxE//d+F+szvLzQx0BLNlD6qR0OsfBm89FhPnZcF
ydPoDTUeJQfWxSw4Cdba4QlNMAo3gj/rxHP9LX1RwMA+fv4988NQ7IXowY9TGMhP
trJnN/a7RgC/1kpod2/Strl7a/7dtDfa+HO2/kTDgpWwRIvIRkruJOUsI15Jdvb/
JYxkm3fPx6+YcsUudhYXUQsYwpaiIRYQBqlHm/9SYaMv8XSWXnpFlrrCLQEjgTD2
/VRNeV4vqMYE++EL1E6l+zvgpD1ZwqucJXKQXvCygJ9NtB5L2Lq8ub9GnolUxdIa
Ao1pXHA8vAit8Uivyo8RqCnh2gJzG6K2Rql7uGFuesCgF33adwkTtxR0yjq5JHjw
8gtY0+rCL2pNtG5FxgbkPbT8cYSOkSogBxnjazDlvJrPoGZYd1HpLrsLRjEp0Kk+
MNv0vPmoHJ/Wl1w/SD7EXpaWLoAIYJ0KY1DPyV3eIzKlD8/fNe4thmlfPEcUbEd5
yTMf9CpPBUFaoMASQ0gen8XuR6xL2A4yRnANNBkTvDt7Bcpf8dPuYfpIFinbYoMU
APBOGYljCCBtVNQkETuWrdeG3VMz7ZogRFll8u5AebKbVxk+MVAy9VPxuOb5FjrZ
uXQ2x1fO/XPdHbs2ex17pQYJ5hC7x8FFDQeKRh5fvOwI4hzF4WKyxF0AujK5X9OW
KmWQou9lpdqg109Ydl6Kf8/3XVwUWVqV0jqDQCcCQU/H8DXGBFXu2Ka5fEhLqiV8
o2/jOODOH1wIJ5WlvPxfK56QFL05HTrwUo5oLyPg4/MNwSRJvJhiXGSiY0RsEyy9
e8XKSrNUry1zQcH3KZvCddZq/Vpu3C1GkmNj+zytxpEcT1z1yiWqAHn5sv9xqWVn
QnZHbNEMCleuMrNuGaMrUa6Yc9mJRQqpEd+8B5nEGWS3pu4lSHmAc+5h8H1QdrpA
TbcQ0PjZTIU9n9+V7s/5ILgTXNpHrNIVjDZbtF3cy+GYevS5iQeoM06x6v26SvEU
+o0Ajc3r1X/kdA+XBfPFkR2IHFJt+bKdZYwZbNqt8x8zXySEoM2oVkLgzW4Qy/AK
+jKOLJVpqPHA0NgdNh3p4Ng+rAcY4682p29TRJAhFGvWeVZNC43nO4FARbYUEVDq
o7OFV7GnlhblabFCVVLRYznKivrKwq2pkZRPLZoLGODZch9S/JR6KAu1NJfN644d
nBDq6vAEbVAzXbsplCLKLLPnyNhWB5yoOaxUTJ9qk+8JzY46W+RbKAieu+tA8vba
84BjW9ig7rF5cYOE3qv0EPEZRPcEWFVOQ3AReeOSQkCvDmr1sdFtlJ17QAaY2+Zs
25AfwrrAyNrH6ouM4ScLH7dNWDbTQkzwOWBkQ28LUuPoEKM0BO9CHcyso1gSsp7g
xibW/ZQH9nWPryomTp8rvH9oVVeecRUgznX40wRH1j+bgxaZVGe+x6Ae/l7YtEqb
aFLiLxEMFrD6K2VTNXk5gJrzE2wKL3H5WI1uMxB51FxbsZVJejWhCpCmKDZmKvrR
PJNvhjHlS4Ik9BKBpE4WeI+J3mtUSesy7XBPgDON4jBYgtyBZNeEA18CEY20Rjaa
0ETznRGvqvbqpO422z7iixijnakOXkla0od92q7IFTXdECGbXhVsAjX61T0l4b8J
c6N+PxC95fCr7P+WaTqmvzVFfV3e4gNcdm9wod5osNiO1sM4+1AH/5qFiySUysig
UMS71D1L+zp/PujD1Kf/TxVkActAN+jdqoGbH+f+FyEyWpiN2dnG6n0+zupX356r
JsVrnvhdGvb1DYNlQhpGjU8BTWw/6nF+2SPA5K6PvWKN8isfN6J5iAqxSSV6lA7A
+6icKSzV6vYM8sVq+34JIVsnR007AhFdsX/gW2xJmHsJZxYXb2s9u0uV5OBk0xY3
uHPTGNMKojNV0vP4XQy4LDVJnDis6R2XpMpUOmapQqA1znh/PmT2wIqT59cqs9kQ
cAR4qSH4Z4ivGM4P8d7lZJNb6k2TTNmkRe7STLNTWGCplRvoDZIRNQxxOR8JXWlC
gKg4hnj6A8U5OcHOfnv+nLTR3ZF/RWmfN4ejtxN3U3UtDI1OQ17lDT2LWuyo3YmI
7xGD2QCR3yG2z6ax+hu49ec9B4UVKcqp9hIy+7BuoopRLP9yGkQDaSEv0XtbWmve
He4z2g/YQkcRLqW+FfPvjwIgo5ORqgOIgd35oQXwz6qoX5FCfnvSgsshMPPoXPM7
z2fsW5StiDcxwJlx6WN3xLD+sAaryBtfRjgng8u4oOMOuDLOBwyttY2nX6+BEn3H
Vsu/uWBMgeNG9FotzS2bcTzTvlVN2Wu6haxuWiNHD52iZtd7pdxlBjIfq3ehqJ74
oe1IX18jVqF5mu+6Fw5tpMAWoLCojjbatod4QhH0UWmviWNGTan38umcTIwEH3An
V4YnZlQdIceqcey02mWSzyQt62GL5D+HQ6XkcTpSo17DVcmn4P8AaCMfQlSAcEml
9NDUWSsNCBQhhIb3TinEPSqnJpa+du8sLH30KjYu0Q+cYpRrX/HYUi1+aBU8+WWQ
myU7K2ShEjve50QosKS0ikPtgsfhvTbNuVQ6QsB4gKPtOQiOh26QIB+r2FDVnUR8
+0Qd6SABlDE1QD/7APItjy9eM3m5ZcDTAd9vPfVP28v/OhyuOP9NmzkMMPh26O83
g1qCmlhrjVBwQawbi+nWyppq+vlDbKp3g96xVB92vhcvOvqevSLV/T3U/ATkJtIC
DibnAw8c8qQGJMu7+gcxl/scrbDbtY+wytOnpDpfDq7SCby8L2UZbbomGcRm8K4D
H3FzBFScI9tlGo4hPfvASONT2j2IkTwCky7r3Ky6N6mQBwmqiM0UZCJO01zMvjKE
rSdtIV5ZhIamB2e0O/JHB1kPEL5pZqH+rdGyyn6cMfv73hdrvuOVFCoJRl4H6GDz
Gq92LgEcYi36ZSAu+mYtKIWi8gPqNalOwozmczt74WFP86WF/fgHt01WirLNhBZ5
U4VFJ2ba8VOnwbRbe1+8Oj83tkgCzgzEuCnyTlH6lMV9Ltapm6wSQg6Bp4ffMQY8
frH7fps/WK5xbgi5B/vOZTTjLDrevqZZIHgFG2dMSvGCovb+2qPYGf50nmTmyZZ9
i91XNCvN3OQ5VtxhzozNIdvDJYx+FBwRjh5PdVVQeYojY/lLK62wdcdVRw8x8b06
0MhQiHpYCc0BntJykP0fBxVsfpHQ9L3yxcjjtP9V/HRbUc+Gu0T44biHbaLvFnpE
6bma3AUET+61GJHahdFc28HG+pjaYyvlGxuSdv8RMpIsz6ykOOuPUCbwgfxRQkYD
p35gWtC4lJgxXdnG+jOen/e/JbHH/1RtDt6/tbCTKpMHRjc4fW8rMolTT80L9eDy
K1GKXF/yU6Wyj/N32gFWqiiVXvbWInKzUP1GkzgKyKtaK/14k+v2TP6iYbtp/GEG
QQPEhs/iLTNt7rLvkwqKA2EKJTD6NbFLNVfrSbMfSBxYRi1/60ZQJB8+g9k0FFDg
P6o5EOlRWPaOEjGf1UQPthig/joX5pkCFfwRN6Il/nt88S2XMwmimKd3Oan+t4tm
oYYUl26jo8THMfcPbwv09HkbJRtFF7UEwBZE/4/Om8eZA0xmhhsXOMQ5WHykyQD9
iQygettNgKEdpV7zbyZiTJqx1E/HdZjEMkVfqMNnBNNXXAMoYfvDEsPOaFAznrW6
EBO+q+Ld9k6uyYhWV9rQtUslwRG2Egx8Z+4TW6P0n2rd6VAmzUYusB/yhWqcm3pi
FM34PQmWPQMMKx9QUInuXLNVXFCdNAojGlf0CztApUrZoCiTvAIW4be+Y2s+CCv/
ig38T4hetFAiY5U7fgZa69RwLVQqiGom05zCyJEBZiaQ4swD2VyvbSRbgvJIxqYZ
PGmaYc6O3cYV3HpNhqpxGltpYL54/U6KrO+2ygfQ5gSWXplAjIM706Xv4tILSZea
fPb/GMtiDcT3QEoNGIddpjhdJ8DdKcRCUCADxMTmzq0JaUoGPRnGvInp50/Ec7lm
xkfevrOTnJio8/1cxS06jV5jwNKr2eM3W4h9+5V3TN5yM4F9Pt2Rew3DvKkGMzgz
YmluLyiwknASp0lLVJwxV0bJqQRK7O+/FKB6XxshoqMpEiQcnqtskx4XGQtWNwc9
b4+UkNBK3nYQEWaiM7IMYIQmaE9VLYO+8cPrE4rarSCpe4AWyqQruRz4ynmKyMEc
evLDEk2kxMFsyiq+luPNuu5o93+/O2aByxlHlau4ltof6RLc1sXs6M/W0OP7FcuN
8uRqDVTRGTUYmBZH338YSHFjLvKOcJ5hg4zT5PtbMwczabFsZq1z139W6N+rTi1Q
BVjT2FIrwImvYBSOYFZsfM3vwL6VLqHkpBOgu/XKIx3bM1CsDI5vr828eindSfTv
zOHZbRtQICbg2kN+R60Jki0VdR5ivGNs8rCR36w+DuyypdXjLHxUAwKYCiM+gRyQ
4WFA+Ci414Guop2kzmh1Iu9u23y6wgU3i798vK+nzH5phajYelvrjcSmrxHrMopp
iYPtNN29zNQETFwwRW+FNaKJz97iwVRygNISLx01viwoDGIgJ+UQvgZ5iVLQfkUK
JtJA8WfO5nvmP4x7p9ZprXd6WksZ7nrKsyH1gLCpwLVc/rATc7Y2RbELm/n6io2x
ofc2kqBS127Lq+HGci4+N0Y9UhHPfW+iCrPoiqotmDe8yEXqlXdkq35i6lrcW/i5
Sfxm8JSG7s9fGiAvP3nWaJHA+n/G0olaSJ7cm7RM098pj9Pfix/cQOrk6DWxxb6c
trs5KhkdDnefMMsrJLBJnmrlKmjhaFRGnAiIUwLItp5EeS5RXpjnhGYmef6/CmCO
3Lkm2mSuAdrnnB/cyEeQyqLP9RejumGuTvdTsqgmHt40ZkUtLnLzOzUPw2rbbBiJ
eOkITsRlBZujlonbIhmlwBzTaj7Wf4ggmJf0a1CdjsOCp0lprJG5xT4peYCbP5op
28lWN/JcXh1NjSFa2VHKhHzYjCAG00OeofW1iVcpIVQKd0/UUTlKN4shYVB3DaGD
s2aQN244+aFB820+z9BrWTyFViFRuMu1bPvuz5iCLrJqqjpKv65fvZVKqJjEv7e0
RCH2j+S+ZT8kNxOV0J9ot3tfplac7aXDchYsF9ud37s3vPV4QniYnkhkL23klTZm
KK+ZUM78DqI62R1wBZsm/q+vuIshvkkeoV2CrfngnUlhvAXCx1X4HNBJkOV08mlS
2O3aKDb6CxhBixgKaDjy46SXC3+7ExV+tR8uQqqs+N+6WPFSoCp6/jZMPd/0tJo6
K3BwedkDlYkhuWhblth9l9u7pbhBLhk62+kmg+gX2UZgJb2TViPVKQTpyfw+wL9V
pwdKwA/x967ZJSaW2yDeI4OcjuqGxxnaVgEDbAndRUlBf0UkCaGU0CqAlPwyGEFV
lvdKG71fyq6jI82xTVH8Yg1WRvhTgaiZ8mq0DK2YlK9rwnnI885imHsMmzEPpZlf
DHIZv10bVYunaeRqSJrhCbM+bvVu/cvZgFhbRkl7SYIKetKQatTQCMtoQgrt0P1a
kNLGm+OHXzf1Oh8UbNNfgc6FIsYth/CG0++Nx2HmXNlaDUf0C8QUTgF6k8JJRA46
rdeIJsNjdHtVaL5WOwyf364DER2nLHQUMznamKwwnfNyV9lL2yjRIC8M5LnQ4GYw
hGa9/ac7sSS6X3Kl5wYT1XhyEa1dS7r2+Xzy7abS5vhoVeePlVHB9vyzL5BibUXE
DjS3zUHuZsaB0s+O4/3S+jcAz2HEwPb+r8KHRsb9DrMUs7eAVyoAAr06en2nJdxe
UHnVnT/4ri4bK65N95mOIAt9gOgxr16pqMOhNvyjnKprJtiN7OdPBe7lOk9CQYFw
eGmGWOWoqFIvRqNVDKcA6gwCP9t/l4Zepfx71Ty67b78oqoWbSEOx2OvVgGSWbCw
7/G/8lUWCDYms5QzkiRJN7fGw8QfivTRYvZsifBYbJ+HXwbm3SSIaBJ5Gx15YRUs
FQMCVqEoyKTzhrROE4POc9vGuS3j7tYI6HzR7tMhmhI3goM1OeEE2j1a+XSOa0Tu
fMxvrWzn5vyYkb4uFE7V/qhbZWoKxYLLMQJWvmBLNrDpbsPx8Dh0kbbRIVaR6uBE
rpVqkLAcRltO5Toi4IxyBup/P05j5+zkLFf+2vOwo18v81ZPBsqdHRTkcN1bUDAp
Ugpcwww2CiYkZ4Rl+n0ktGDkKz1mxXg7IF54HgbQzs5nZro+DbEDl54e3R7r/gJG
HvaSm+3MnWK6NnhhrXnKi79vcEJcjbSpDJc8uzH5Q93Ar+1VkJN6T/Q+XMP1QSAh
4nbZupnLf7Mw86k94iczgkweabuSu9F6kKQm/p6k+KaD8Hav+hfTL4e4V5qed2Zp
/duO23QA8MnZ2tfkUKoGrp5IyNaTR1B9x+/icihWfqVvO82V9elEZHZpFuEaAOgX
2yVPvggMw09vZwCWQgY2v2FS9//X57GgfTSQHqq8o4ELjAJQBrWD554RcoRDNPMV
jjFSg0bArmoMZDdks/wtyJFVo5kFft4wEU7/gBuVHmEirizNT6ZzMOWEzAf5uGpT
GtcgdVdcDKkisyNsrXUYcMSTvfhtb3BSJOzQrSJz+cTSFma1T+ey2DgEdgOb5JQf
js7MFkOBRKBSLAbkC/TA6urFTC+c6IpNjDyFD3Ldrw7ZGM8tEKr/pMQWnzUT5Rrc
Kz9mHC9A57+g7oupig/PCnDQrN/9GtwSloNTiflQtD9LNtX8OcB31kgzpHWJuU+q
PGgbFJI88zSbml8Q4FIqFjM9kv5An0pC0XTQ/Em/SQMGtQ4NEKHIBAYvath7UAf1
8EG3Y+Dg8iaYbPUfkQQJkEPANNOSQgruBjMDfYV0E755MO+dIY/s7pN0COaczAhp
dnDrf2uTPxAooRfufVM7Ex/f4mD97ukfbcdLYz0J4/HeLZkR3T+psjl6MOW+SMpk
YLlhr5zJX1uzmwqdiACemrpN6vavbRgzhoWrfoAFggQXyZlz+H4KsG6K2XHKKzQ7
I9XEXQXZBrGZvBB7AsglOSxLjc0r7ldTojQttfq2nscnEwKQAx8PClZuUvKS5ORN
TtZ1ysfmFpL7zR5pOUFBUBnJ7d27//UxeWRdbbFnJk89T6R3JUrX1FkMvtxAIEyi
uN+uCmRYDIGk3eDYNuK7fcagdCfhZcDoX+uHh6qDJejA1zOvgd9qU7QmCWabwhE2
Jd4EIQgUF0ucK8lsNhfs7e+vUQWhCx/A2KigvwtR/NXz8bAZ8BehSDlTLzMeZFef
pWihcBdj2Lg47yg8yiL58CoYa5LHz6iRPRqXpwPKkCT0cTno8c9+MN4qLLUPw96b
IviGSC2mxxL8hH9VbYlbZQoMmu80XFavjo5AzjpNiRuSnT66V92mrmJI9BA2FpKy
7mitfbnqJXaNsYrOuNkVg3S1rXhj7djVRBDLWovQxj8TyyBsTs49gpMhOT9IIsl3
ZFkm3VaGU8tuqdKzUSTUTL4Z4T5O8KMBcWK0nIN8c/9aLvOxLEApMLCjFQE28Dcb
LbODknn5IaHpOMJzxpmhv6Z75AUFCAqm396tHCbaetiVML8O4Hj1Xr+HVxfNtUV2
ij3xGC+RVdzR0LuQ3kt2Z5j2nGNK8TPSDo8bjVwdkmSlRKz5URfZ3CwC88pJgQAa
p/tSdbtoFWdjpFygJ+Zs1Yoq/K8UPcgP2jsPYPyd7tkfBNjBVIRN1d234HjPZBO8
thaw7+/YZCDOFtLnINl3j0HF9KKT5C2Z66/cTRkT0atZjpqWQx9OcXqTxtHBeHIT
iYtukJfJ43EbfKp0LQkFy8PdsCBPN99DU1ZdZKIFWZXBQ7aysPPVNtmebS4kqRy4
UfO3Zz4qde5gS+zKNgJyCgWbhXszuEFnKFexJaI0wR3BkTLVP9Q74Gdtqx4gCoKQ
CwScjSunkW8GjaFqQJx3RJXl4smFSgnN3zrKX0+ztlItYg8QsDmrfYTWTt1/dBX/
QdLIMGrKUE8m5h4FAdDmglu26DvubfVWA++EsM6vFVoFGPf3IvwMrgbQEOSI+4jj
EycW1QG9Sv9cBNCu9Y6uZfEPU3iRxEnknexImYIaFd5BZ87QUw4pdXOmEAyH2Y3c
2pusIfIxDTsCLOtPhm7rbuhxcLicPJVk0xNarrhCA1IT/B2WgjuY0tnxKO/IPKh6
NeND0RJv0LcTidDpy5FpjpfZby4v04xeqXsxqZSPrOQojx3bRjmopg8H1yIL3Ogf
z93sWU9yvL8JTjoYrMZLjC40/KU4vctlk1AGUzUQiKcjUzrpBtMMDF1HfP9PiJQb
DEXvcwMRpLeZeQo3FSieCYIvRbvkhpKA7BpUJtsjgoj4Bzfzwlv7JSbKRVC3QGME
CehKN58Bn+4vQ7mJ4YwPjyhh0BTkv9qtYnYBiFeWuTJUEnqkUzIACcOM6gWJ9VEM
Ch0i5klliHrX3RfNn7+A5hbybs07LGLtTJYMcnP/AT0s3XzTZhDHKczxBkW6w7yR
Vq6KHbw5h+fC8uBujMUf0eb4wFbB8QuGUcRl3txAiKNdpPSdmr872FnQhY+TIB1f
FTcspVGCg728mysCL7ww4P5mDW3v8dsP9bXS+kUoqrMO+RVwMPeMnr8fvg9hpUX2
2soJtMGSUrJJXoEY4VgqNST9rt1CWiNb6r3ovCmNNeRVshuKeA8x///mQjVmpLgp
7SrDOHFnDsPvm/Patu1xljQ9DhMPXbd/givulFoKRECkn08tibHuuzRmHrtQ/jUW
3EzZ8/BPIHJqfYbeABoum+JlxY6iPWf698pt/YOhCMfAlH5ycR14c7JzgB7fEfRP
JYQ8/6r40GK4H8SC2OlbS2RAJut2+H86OaSZsVWoI03WwS4pS5P64DQXqJ6E0P6S
kIiajQBUs4vonwvkCdC4c/FKKhAHXxjxkP7PfgjzzxrAtaS3Q9cQA/AawzxB9A+B
GE/fNFPTm4yYfz2PLjPfdf/aI2HGq6OPXXBnrX37LevCcnEGhxYFlp7UWoCJdCd+
o2sCNywShlLPaLOpU/Vp1QeVLwTeV72Ke/WO4Lnsv+Hf+m7eU6i78UZ4ekbIGAM2
fo45/w+UaDlyO2wWD3DG7wK4V5PtqV+HQQMJUb9DXpAD7zzUH6gTjDZ/psAVlYlC
JZWbBfL2RrQ4r7MVjwZpFMzONnoKFRqyU1ipAJ2G+SJTQyg52vWc2j6zyhuPm2aS
z+k8zkxJEfBnQlRd3fwN7oexy1tfogL/oWU+/QWrGOlk0/p2QMipPU8dvxBjJYxA
lmec9oFG0QpaWrIH++mzDwpPjzV55c8oKASDR2Jor4ZP7u0mHiCrr0Danxzw7rXb
glN5wYUzkx4VlLy4bj1mB7U7gdiTkNYOu4LlyWLtd0QuS+1I/0HpybHFNIa6VsD2
+dmYCHdmG0wCZpiQBczJ1jZmwtF9v9QgG/GyredK2DFWK8+VoDisNgb7xm+lbS10
zbEu6z2wht4ngGfQr2OIuyouGD8Z7rUcHzlnHE0Zy0RJ63oAJGjwga2SLPjFpKw5
Cc/H5b69ZHQflA7HL7ihOao+spiJZMJVc3CpMBDxZ1xdTn89apjc6doFq/azdQ/s
ALFDVX0Oi07yAdlsyKk46ndwimtejZopeWL3TbmTvjLTrCTF7I1REXwkOnGykfeJ
J+7NCHUYmRSwEfQDtsE+4dETW9uRQOaNmLxuZ5QrvS69EUMSvqJAAnqQXlrIJVXD
fWLmmtQJBIqEn0xWOpXnC0rh5AQ4XgelPbEIRtjm/xZl9rwggzn7G2vJ1G60I6l1
eD+B+ZNnO6iyEAP8w22V4QZyKwT0qPUOrKRKd3tocyJwhquR1VjPCT5YV/HirqHs
PVV2bjuq1q8qynZQLNKO6fbDA8BGUIhJ3ZDkVZlSsHqCLAdc+cqNQSwl6JPld9vr
Kt7pd30D2jtOeUiL7kQQ0ew6vADQ6ME5xp8QEph7FUpn6OTFhMrKbSWH5+MnL6/d
LLJ+yI9XzTtEW6POKoP1AyUsy5WeU+X+I88KGbIGXt+fzKcjpgHBlDmMQV3jD0wW
zyxXPa7iC4bqM6VAC50pLeVMfnj1YGiTa74ywv36TSwD3sZyyJnLYxkiDO8S5HFU
K+WaiggRpaYsHeXUXF+97OwcPM9b6QVydGVcPWS2LEyenck0zzybtoZHj3Z6ed6g
LgpBkxPgWnVwnmqMt52iq5vcUIxEvjCMToc9Nk+NXKwVWWH5mrvOqafXFG6klpD1
hBUQyMJ9MJHI0PxDRtc8xFrYhqjcXuv+1PquQy7c0w0McMSrashULIX9TKOCYk8M
Bppz9v8/Xavt+d34EibRfKM4Ptp04RNsRGNU4ANbdyIhWFAPC8U3jyKkL72Lgt5Y
pjQlI34VvlbTupFxiFcvDfWJvHXfEi+7KMHih/na/KUyBWgIyVagLmKZM1QovJ91
sFvwK0qhc/SVLXd5JCkYE5O8b9Sak7xdB9x2u0KQkt7CBea2LZqreHfr6WXaibyD
vIdutYSwPbtDlEZil0oYGSYiawc21Kixv4+Q0Ns9Dhi92Zy/kbFXY5ubmwDJBn5j
cZxy1lxsOPl7Cil422+/aDIhqcf55UMhrEV6ueJZpEvUoSDQc/rh+gt9qTfR7dt0
56OLWX3am9o8LytFSlCIrTTGhj+cNYBkrnt2pnB8Kr5mmJVtMXk/il49tUzMgxv+
09Y0esdRCaObxSZItEaGPBXNFZ/4bUL0tar2rQm37DvYVkLTwyWZyLe8Idut4tqP
+HUdPOBDWg+C4N6ygNPUDgBYKa7tnrhJWei1RNv2TyUVLGsIO8BPACxhRcc/Cjj4
H1mcu672D1cHKk1OlVg55PsJQtQmlaqQa9hx3qL1Bphhq2YAcBjKcDX9hR6oFUGa
qFk3w0cWoLPkGYUIVjRI9GEoUYtzz+2c7YrnCczvmT6ROfRcaTrbnGMrnRyfR/BB
Y2LiUWlwmFv6QYahpCw8USe3vEMIpLZhFsyH6LeRL5lbdeTFjs88YD8zyPI1Np5l
OXqBmk7HlLinqSvrCy9dbuRGYn04rt/J9NmEn/S8OKGNJUHNaMNLb0U7DAoiBYNj
Im6l7iTR3X4OqZa6VY0uOhNJkHACPm9tJNmhYFsl5K5RVCgZRUeOgXFt4KXOj8MT
t8/eu2WePtIvOPKwjP1Pf9XK0Uy4QQZtYyOpLf2WT+V5SAXwXxfV+CBQIK0EAppx
oYqGAsEhIRUpghV2MDYFB5wfAA4YzZ0aADyysf+HKi4wncKa+cPrEVHcXgnTDZZv
CXyWAcYEjJLhqBSYC9hWJn3OuyMdl7K2YnZHBUtvBDYM78Jkdt+/wxvr9bpt7pqB
lMnBL3xobCsdB9ifhV36YFTCapgO3cRKjlmrJ5db/hhKmhMlVHk1GRGuuy7PpeRX
bsmsEqrbJqCu4xgJouh7uSJhT4M2lcAZkkk1Ym5iAh1qTi4+mGu4l+Hwuruz9k4+
xLFA0ke5weZZjoIIHdHrMQFO/iP133Nxv99QkfgNaCL5Kt7e/iWv3/hwFOuKdPf+
h1dqvoAffsZp9r4fc1gsafJjrOcpvPs7pRdNIg2D6AsmyeK7SAh4erq7ZfImrygM
F2Cin3WrU9ZjEelpDnZpn+N+Vrxman7D8o9nsmUyVabH90gooaLYal2Dn7s3An9i
nZGemFwwP9Dn2L69HsvnjQl2NO/vlF78vToP7TzYbCvmf/v3DxisouTOIdcdiNxU
6JqCF57skydo+pvziQR9lSU4VEkB6dVLjeAKzyjgwsANBeJ8M42o0LkRdRy0uHye
q5mGNAbUkKxZSqOWq+Xjyps729hibcRFUQgGaMKPDau1jzgWxl7AIt6d8CYEPAw6
FOOhQ4XkHGcT3T1AxMxBa9N44b5cQ1E90fIBmbqSZEft9I2Qlotu11DyrDr+Rm4q
ou+HUorFAK9rXXs6c7xVhfuPez3pJa68VzfB3KD5ZzgtFgG5Hg9O5x52DTOgJx3e
3yoTwGpSGiBB08I8ZwOHVZs6CUTprkeb0Y1ok8Nc0ch7UON76SvBM3Q3ZTGVzsZ+
gO0WBwE75k9flGCujMTesZ8Lra+X/HbXvAhgE9aAM0OJYVFxUycKuOgm8AVwxJ5y
BlSIJHroiDOajqNq9DILkhJNucaRSMSj2+3/5nLuRIQ0dqJengAGMGhG8xfWaYDO
twRCWyqEyf2bYa2yPTY2odA8PLpaMW04JST69Zn91n4TtdhL8lRZhQ2IjRBHE5gC
vZ94GMrrsYTmORBIs71e1NVSN+k0ycP+F/ylrAA1N22WWNPFwe7ZpeBOY9Npz/Bt
N2n/WwplA+KnNjymtD1Z4S6spNT//7JGhgUx8hcTUHjTg06LioUSvnNlC5sVOcQa
DspBgHRakAZDLwEF3UAl521Wow+9ipLCKIvMvjcmDlBXNMKbLPgvnuWjAKd456ub
dG+QXw6ZHJibmGC/b+mMxNxn3Tp/DwyhRUubqavfAGcUu/SGn6rrxkUDpcZI1PzX
4QMB7rCXIvBlTlvBHyTbLe2NAM3/obHi6mAi4NinChvmXembQh37xm7TNdy6pJp5
YXIZtpkTIcANbBqT5MDHIZ0QeCsJrdiAOwtbiil62y8wqYsS/HMUOwfu9v117IM4
yH1Vyz4fDcj3Y0VFisxkA1lLrB80zhsjrXy5eiEWSQg7oJ3hUFR5F3WL5GFLvfBV
160kKCethdEwqDddxhehrdIgEt6qVSTiaqB9inaOYO3UOwd85lD9TTQs2J6LgFun
bV2I8h0fYUtYEm1PBJfywvdE170Y2XbZg9OWoMTZRVS7OY2U95vV3OQAWWbjErG9
eIKM9p6hY+mUBJPz1LSLGhTTFGMGFZZaDF21tK/MiCLps5yEgSejZMjfbIDp2Xlc
3hDoL7HscG0oQhUksXZvhg+ZR1iAIH4qu+m1R/Zua8TSV5bc61grjMe4hPJBKnau
VPp1YwIL/R8YTNguM+MZinvkAPNJMY0HdviyOHL6QSf6CZGO1SjzLE8tdI6OipUm
61ULug+YBXPNwJZHGCgUpSBK49do+7eGp0aQHaFOw0GmOG04XONIgGY8hboQ/Rsd
lnXGNfzi49/ALrMnGmgtDftabMN+Pw1ckSCqaeR2B4J/kuYEQ9nSKeVjZtjZv/3K
l80/dhXjLVUrNWktbKc9dIx4qdPBMwlqvEV19PpI5iKIXNN8SPDZEMsn6nzQKXvU
fpAdQSy8L/EDCkXCDKHT9TLR13R9nPi93MgxNWLXuSsgMV4TvdKx1K+h8NQaKCo7
MMeB7jKk9sa3C0mLMGIDCQlbs+RY1ZDnWH3BdgC9b/dv6nXUPMUispThuCqSyC7D
c8EhGcYt8Z4UYjLmOKyoFWyNTlYDXi1sziOm3RXMLe/QCH0UAeQWw4ATUODmWKlj
Vq6l2EXe5cgpRe9BdAl+xVH/je2/iObRVOCDXwdOKkHSz1WKzwEQqvSAJ3sP3KtW
2Avwvn5Ysh7fkU6LRMQ1CVl1OKxM9Xp84CYqKbDKG3A/Jayyck8JhwB6FaoCC3fU
mFQ7S55ZjCZ3/SDq5H2rYJjMWOT0YfI3OFPYCPeNmGhvJB6N2QC/MlfQM9RJtpPU
7E5HNyL8CA0zp9/LgsKaNUlfrXBfHT3MIuPFt3ojIAmQaqI9ueJ0MpDrmkSyOIsr
1C8OYU/yvbPMCiHe6EnGT4437jTBri1yzOj4yQEyaA8menFTVAoMSHmmkYha+DYe
itcWTXgopGdq6Jsj62/kYA0wwdeeQ2ndkkmgyZrgu+FQ6ZA0ZcC+NolweN+orK+p
vXYiPOzzw8vtKhnfe5vTh6EFSKAeNC80ddCxQseEjBVRR2BBajvOeXCWMeD0TM7J
XnpsePYgi/6MPYdmcUdNHNYfeSMvzfR8+9WvH6RDWEgooqGXCmEELnZd9I9a0TqV
R3lYbwdsFBKv892Cyi0lvGfW8zHVza5EvBnXAuC2xV5akbcQZgvgybhiUYZBY3TL
zDvlv45gJAKvMBchXjRcGZOeQTU6LsNQ0tKdtnedxsr1pEYhn1/twJkVUlKvMMDg
8HTx/H7E37eAi+43wMca99kyOeBiH/GIA7N4MlZgvXpzD2tSwDTnqeXD2i8ONAa4
38wzA2UP2PD1c8ukiQ64yNQ31rNon1Tj+MSb7gNPkl2GomulGIfdZZdV4rfVUgTP
a3hm0x9IH/KOBhAgREmdks7sFHvH3hvB1MnvVail++1++MU5GUGwyyc8oVM5uc+r
dXqPbg7kI06LzWWCv/q0R7xv7bhrybtI9MSiYUgyHYExjFxaW0uBv2RStTSCIFdX
r/tfGX849RCznP+t2GMTcc3trovGD+iCg0+bA8SYuFY1ef8T/eFnIjAN08m/wZtZ
2ThKAuxpqIy+nH0I9Suj2ibA2EEUE/PyKxjIObj4XwZhDNYjpjqYS6QTOzuhkH+V
pj25NYu/iMLy4EepVYmpovja70pHr6aLiOn4zKM2IG4xaj18ZJ66aSE4h8Pjoekj
qRMAvFPg2VpPqpZA3Wc1OUmH0J38yqCXKNV48/DFZfXFflfraafBP2KJVC2vwcPB
qYuYgmNzdym2TNM/mXwejOkidVHKFSpwnm76xcjBbW4n56Ixu8uA5ggInn8JvQZv
DXMQjnsjJ0GyWiB9QRa/ovBdYugosHAysZowLmMEJH+VHqvw2avZeuCifDUpD6jS
IB59JaS0AY3gI0bcMhYmerdn3uQIVb7P7g89nuYKrMJWb0K/1dRB8e/t6h+CrYCX
PUeUOo7LtSfLeN/8hqhUwHnpWZPWqqAsIRhdsWO5DaSaVqL6VsPRWsYDiyMYYPzL
uJO5D0kh6Q6HV8YvSl9glCHO3Ial+Kp8+DlBOTBtqlqxKIMbUP98F9OdM5iThSvD
uV/n6k5uW9YxKJcSYyTKWMUFlIgOEIWnjeY2ahiPWTBhIopBya0okNSeWWRgVCS5
QhwYjj+T72oHesdh4xpHvbT8Vs9CwmcIaBSl8B0jhB+niLxS3VixhAB9hQH0mWsp
KuVQvQVGFBZd7irET+ume1QDSnLVwjoHSLxOHokrlUnDq137D0Yq7fDNsmO8JATB
TSpHB1idb3WIppswAF8DX1q37QuSB2TbBu6oOFXMe7PxVIqXdkWWwDRe4pD9Odn0
dedAcAj1xdouDE33drwl1RqCgER5mZzW2lbE4LoaYVjbPmxsP5vvR0nnJZBSd4dB
S0AepvrAqlds1lJpYjBi+6JSHsXuTCjgF5/HrMV6HBJST1TOkgIU2tLjuafMNRpn
tB4stXWDElP4N+B19XfVbJjfb+VOBPPYbj8H+yVVCimDlm02t4D1OwNKYVosPYfW
kB3f6QbrFHjH7IhAgTKNXJ8AeL0T3MR7J6JhHrN42XRm+3tsuc326iAQWgAa9est
mVcFrRZNBWq+f0TJB32uVlDTejY561yZJUxKmoiw2/IV9kdgPvhbHroh2ybJScDj
mGKK95bEU85dL4XhLeRlR3DFCW81V+RJE7rLWa+S0nYHL5IONVlcTfDF2myQcVXX
qQ5XVtdJ85JQvZ7vD4rCcQoZEii1fUJ54+y/Qes0j/mTVt0UIcSNn02MZx1mTlCG
uo1dBaUH9MD6BpvlG6/PyvkDcZRPE7L/byjDfhP08BVBPXpva+CEP/oZfjfxWiZ5
sfgbwmPM/6272Bo553/kwIgN7vC5aV8lSw5f340FIII+N2LajtR8RDnGpcr+EAg7
Wd+1Gezl8OMwG54SnO/e+bwpASQQiEYFA8wOKvBV6GIXKAWT3mhssjS5uC405YeJ
IB9Bkr3ldWPvIz1ZuLj1fOqTVKJpIfUfWrjHeaVg2CnmDDTlfAPBzGNJVdTCmJu1
vXqXX2ZrJoVeEG7XhpWurJCo6p+j0SawGD8mb+DYJsV3HeHZPgXxrMoyD6RehXeO
/f2nVP/gesLJriulNd10uPSWIL9qsw7mNGRG54aQk6qLTOPDqwPR9HTC7FcUs8YB
vyjqbKJRC7zp/KC5SskQZjieUPDQ4nYxo4ubOedYZdo+QYjcKrcQKv6tnc5sYScQ
ls1f1mPLXfLF/b868/FL5Txzh/OJIBA7dhz5Cz8N03iTbci0S3sYHfTgWCrq2Ey1
pmQVTRcTTgOepmrVL6ONIGbgSv38ENJN9MIh0ipCSit8SJh5p3U6/3gLGgs/oylS
Ss/nuJOEUVD/BGUJMoju3u6ZMRx2v9kLWQmPutyVEOoT4B1sAhD3aEFF7O1ObpRh
WGM47bCM36RGQ6gPrNckt4ClAnYhfDqgjkNsq59VR10JJ6QPW3NZY8fz4mqxYTLL
gx+ELfVc9MHKnctNHlVaEncvjasPN4pK2jvxchCONdMmbWZuRs3O8XWmcXzmN05A
FMtckKlTO2oEbXyDN3ebpce3adh5IQ5/JeUSQoNZL5lEgmx0hqH3dbx0NmWLs0hd
gAOoFW0WRFyIgQPW2t5MRMVJKqHeYx/vCHuQXZ6qiX100bAwpAwwL5uK/XtEvn4n
0p+6Deuw1IQmUBSxHEu0b5lf+25FXkExuFv7ZSPeA5jTzIDAlIbI94dk+ZDHkbzY
FCStrlttxk/twf6Q0V8i8c4qFRlAvUm5PNsm9YRvYoXC2TcDI3e/Uo7n4OC63f66
MCTDeOJMF6PY3OE22G264Q1xDmueYisE0+oZUiQ3OrSYC5N2CFPGLWU59f/FCoAk
kKlLSN9JcOlHcozIbg25mlLhmD0JNrU+CmO8O+BM2CS9vf0/uuBeAnzWIYuiODKF
rvgLGu1KnYIXS9rqbRGMDOYvd9bjoMm1XMaHIMOqpNusndVH5tW+aIIFODHrxFAQ
PY67KD+odahqyNo5cqfj8qKYZduAKkK10c0FAdrY9KSm7J49aEJ3yfkIjsmYLV6k
7wivklKIlSvCBt9LoCiJ/OxkCusNSU9k+DQULNfiZN1pY178BTPyv+r0QVI/i/Nt
Fv3FV7+YzyRuKApq5HCIyfFe6zFBPBvf3qCd1IezN5y4PWME48jE0rgtyCE80A5v
mNOHJoKtLkZObOViu8d24TwUbQxK379t69EedhZmNou9QDwEzelPqfHRkm6fkT6Y
l9MZfbGRsbo3O1zGHctDP0xsVgoGcya6WJfvA47ZzpCPO2W76p6tPlRAzTyNJdJz
SnTk6GUbXRU10fIs+Os3xdM/7jauu4eGz6AeaqUfAOI/ZmmV3IuPCwSnPDzW9YGm
QJL8YTHyGXLoPMSSaeYEtdECTLrrUy25JCkCWvAV2iVV6DMayuoLTuGk7NtAsrFH
y37Qv8U8GxqJWW+6palMp7MjbjWqAJ7f4WYuWxvnJhUcDKRmfE7l+YXsNcU9+XlX
w8ALY3h55dvHfUL4ARqL/TaSOrkWhIhOeNBxKl1tuJbtQyY1om6IMD3aT73bXGVa
ygtMWDMVWTlLXBxZjwNVpG+k5BOyqSL8ASOdrHLCllEeCADPtiNM3qAf2AklUy8c
UeTcjtNW9C+VBPAeRqMAIJg1HRUtVJYQRrCdYoeF2hdXJbmG1i/quBoRDPe3Si8q
JjXgVqNJbQjT/nj02pcvAuorEjmFloF/JuYNeSlYwQ2FD8CZY4EZqhlKi3imWLkW
1Pl9J2dA7qhbRQaz/dr1B88ZGKjs/9KfICbfncvdlpeyLlEHNVhk1UkTY9tGTD27
9YMVfbj663I3vqL2vAE0FVx/M36UgdXq3NHGQZ9Ir+SqgrLndLbE1U9opnvq6buT
p2p5nwZ3FenxGAXzz8czwjvW2lqVtMoRzhkmBAh+Xyl4szivJD7J3h8Wm9sJOtlj
TIajFtvUEuKMaSjwfPCcT1Ww5ymsd3VdlexuztrDjCrvCCpw/5MgJZLFQznGsKgC
mRmtMf7thbNmal32YYJcDjzt6ClGHQimpr0f3GpZufLUINPOlgndjetXjBTtAS08
pzoew67ZOpDudXXLQRo0/bEleQbTvU0fiBn6hTOLXlEcNQIVkI8jvHwB08yvVgcX
7Fz/opgOykAnPhyMLJqeYUcNr6Dg4/+ZhE0MAy9kxZxAIDYKhLlnXAJNghUPgZfK
x3WX6eWfyTfq3KCCQEd3DpZ+qPVDzADb27z3LXdXDBdiPeHCXyMenxwmg1zoybJi
q1xMpPbimlM/u/bkuM47IybPgqe+lAYnhodz6LgSG2mihUB+Kc1f1N5XPmZoZ6pF
jHeOxsFo0HyfpaReVo4pCyXsEPQnWKSP4c0IK1uxmhBva8FKJQOQ5+CkfRBq8euM
jYYXrf/t+uQ5hD8xkYi/bynXVcUt3DQbuhJbYM7NzrEnen8ywyrtvMZ3/yeF9GSV
GxeOho1gUP+FCXZBm6NTeiEHIPIQrszQEnw6NWqU6gRBVJ98/OLN+DrvZ11pMvlA
FOZ811EWgStm4KcbgdxZCz/BNUTdeNXGGWNWCg3GpbynXtxKdst4kUtyP4cZdeUD
1s8Fe3rsZ0V6tlbU+8CpMqakgrhrDOTL4zdB5rrP3exx4R9SYv05mjHyiknSja8m
jTc+AtT/69wnqmec1mJy6gzKS7vsmVDWA6So/3qk9o1t2IsVpDijLX7FbuNDJkjR
C4jNO72HqgaVFVie2eKhCqzdyqMpEhRijBOHn5KdWYT6uT19z5cRvc+fWiOP56PK
8/UAHkFcVf+mgiCQD2KD/y1pN2uGa+/mbu9+wvk+H179hEx4e2LuL8C61xcTflDP
//UesZctE34y13JwA0nU02AjY9jCiW11q2dwYJgfnjIIDH6rsJ6vXCFGE1syJQud
/1RG6Q/Gos9zXf0az+0fokkmCh42qYBJL0HXAd0XLwqext3sGxSyg4n3Y3pV2BF7
vJtiy/54IUNfcZKsbxBqldPkEggOQ3PPSCvpqzZJGPVLnWVQimhly9IaRFpazQb1
mKTf2APJrfKlV65gW9vCyY9eAELNk5pLTbXmgNDFFGXG00nrV5fLyQT8UcI4fBJi
aad4X9tLjcv8VT0umu26CmgEuTEzzqGp6Z2fE8Djq88sATNe88Gs1lUxUjMTzV2r
2YZeUQmkPhmv7HQ1h/P15xRaIN7sk4pjf4rPa/VhVZEkWg7k6sUO5Bv9m3hQK/qe
NIVvvKB9fepyKimh3VIoOZ8hDqlPG0RI2Pzs8i3Wdrt/LX+s6FqMQ9ZQm9GtJLdQ
c+XsZxYj5nRlDqKLTgEAd5op+kkHEZ7/lHrbzS52WTYhFEy0VIbm7EXybrxvorqo
5bYzmpTwmlZ1W0TpgfoWnnz3pOiGF49E25Bd4kNNBpV53mHd6MPgdTLe19MUfDjZ
iHyvpdxw41TQzU+WjB/tagtDqd8KkNNz7AF2mz5j0CC91KZgFb/7V0T0nJQ4Txxq
/vGjA5A2G4OLkBTt0qUCbR8y3vile/4I9c1WCFKMZZw6lRG9n9i5OObqGz8rVy2A
pfECYxEQRGwjqW+ThFtpaWwdHOKThkZ/SaEMQDNp1rx+XoDmuvt8aYqbMa44BXAj
YWBfUZwrjSE46nXe4Tmp8jq6n005hpE5r7xU762jPx6Xt5OBFii6lbO7yry+LNWW
sVwj44wW0tboaFiFRNX488H6jwa9DB6bZELgtG+U7wMV7vogacNnytg8Jf9fRqgW
3k/Ifv1uQyzcjgtLhciSfRryv18VsS71oJwMWH8hw4SdZ3fdFJvbbFUp/ANQZnOk
glUUSOHJFqOgndbDsXhwvmJtovRl17qzP+rCHCgTGf1kMZIDsnmynOLqovSO/1r1
wKzDYGNE7GaD/+2Bs2zLz/Vf6lTRqLjs1rfkw4/7a3iX5IY/eeUhNLZPRRbyv94S
+patGvjGUixZXlCzt+mrc9jX5sbjugNdsSZaABXwe62v3HWRvKG+lbtd613ux3XY
oa22v2cfaiKMZLqWGFBgaxpOFM3GzvrFTJCEzn37aCHho7oEeavFucTsqi7QuKZJ
lksk/CoFkLpwVkrEQb/qfm4LbVMfeU6cl1z26Eh+I93a9jkYT4Oyr/cbhhwfc7Ym
jq9fx+jGUgX4u31FmTRN/y9S+AHoHhGXl/QhcbtGAdMaAVTadCk6Q1WhEv9BkYQO
tftU+452NYz91kvWbGYBOM6p308ok1L6YOTYg89f5iUMfhUVqzBkDQxAYqhOATNd
B3r3RQNX9LiRFoaAPswH6/3PhyKUhQ7ZIA7xaX0uGQ1ie5K3Yg9gY/d5ylCeI042
LVySVpf0+e6Ig+zXIbRsvGjTlva8fH0af1fIJMGQGxayLga1TJRP5AQ2tXwaBCBS
/Lo3B3yY3RR8S0w+YE2Y6VaMDFHJP54IYzKyX4+Hgn8Grb5puDqL/EsO3w01vJM7
oFl0gBLEUSJwc5SiLRwfKccPwF91tvf5y90iXARt2jYzx+YQN11eFJGTalmF0HJX
Tt0HBQIDwfct9y9FwlJ/kHXD/h7AXXAO9xiDPLOjjsbmiNms785Lz7FpyIxrS5eW
qc7cQOLW8fI3/OKbZIentzMhyIZS/NZ249cTMBg8KyKPDVQL2ixnutg2+u4LrhWI
HBHbFKqkiiqfZSxb/J1rVuMe0mMDBQj4E3EDcLFm+tiG9Dua548y+B3ILVsxyNMH
aNyDUiy43l4f0lor5CcQK8D938KQVXV9tJDZCKtU+C4qq+utJUADxsHh23dGf1Hr
98bdM7axfLEY+2IO3v//amVdAMY1eHQwxeKUnCmlVNsuSxBUflV7WLKYrdslSrha
asvKVpHVPgIXMSSJZ9fh40MahjhYxwBsKoNptjBp76RW7nq914OKL4ff7/up6bOi
uS0TAkq56q35NlYCV443k7K3CFqsNMDZetHhiT5mUhoThK9YwpWDHWyVLxQCuM61
5ayG+H4k7bzhTElPOFAtd1AvIYt1OoTEm0oOCJY6feDteYOfHqASlSnJnFSkdsbZ
JRj1iymW9/kO/M3d46DJrc/6mqIlUt+QUlproybo1KHtqyQjLuI6BdPvjsmkeUwP
uzUZW9oRqcHlEamCI7RDzfDbz6i+5VkUiX2lgSTFVwCabEa968FsoSoSAL5Rza23
JPzIhR+EUU18cgR+Mxz4XwXMY/TOnEcSRwgO26S8Br6lkhNjbXStq+suZp8wCfgr
NBU3jCvqHf5RfYPhxYZCW8952AVeEawBBssdscqkNCCjAJbvZQxzk7/s+QAkLOrm
gMggOCr+rn8LzWryl5cU0hkbt+E2bKeFOYWGVxVN+VbwZq640F8C7+OzCRSP+7QF
axNYcpp4gfHcxI8lk61fhwCywkYTHkdJjdvbnOSpR5s+1ryMfFyfJuR+o76vSxqH
S4kqD720WuPL9PEFT9XbY5gjADc3YFM+Aq7z7XYa1/7Uvedq21qqyb1hl02FOKjZ
/5hQgTG0gIieH8QxHk3CaFhgTzO9j02JufZnpp/ijCiNmENPQn4HtLHZNXXIvkVf
O3xqURV8eW04VlxF8RpkiSKnyw+m0sWJz/9s4iotINoaDwm3N9iHcESArhNTkLSm
GQ4oAxFHcRU5ZGzKp8W9aJTptn0IcnW1Z2NsB5122Ee031QnMap/FHgyIXAK+3Il
atuno0VYXPtpgNR9Cqi7IFyYlrzlhfkXv0QNWX9JORJ72OnDKgqaktqpUJMuYo80
WZpejjgWgOD9GHnPLy3SCW0/ddBzfq9zV0mBumChHCuIkduFVMjvtPM5mmPwSfss
20Ix6j3+c3qohRK1jEs9ffhTz0M0Bdj21h9prfOLQ9p/0+lQi/NnOY/E24s2l+Rl
wmil4w8bv1EFHJgH5E3S17v8My/wVm41vJ1tyHYH7yV4nj98NcNai3Mi3zY1Uyiy
6ARIsmB/PkFogje1Ja8eMIpBLoN+1HBvL0oArrnou6g1SXbve4YScH5ZsZ1QjqeE
b1TXXWpw9rv+j3S4Cma+k6rer07U8DlrPAREsTUCg4Eq+0vBCCStsTALt3QjMMTg
c/cTWGlbnpTvhjPwqNF3BKxtC866gfwWNphlqtnTyzrL5ZDqdV4hqZsCVUqwmwax
u7/5VSlKV43lUJKSdx0Fl4Yfzanl3GNrOIc6H3Yij/LUpRZ6ZzI/I3VWD8z5vD3t
AOeWJAdWkCKr+q+DThCNR6nOTSpyBfvavnFjRxMDJLS/q6gQm5odP41HUW1JMXDg
nMGxNlaegPvgH6vI3eXwRMM5ple/2GnW+B3jy7u3XcSThyJU4mLmc7CNrNQUgwIV
tnQtDZnX8FBmhJWVBq/gASoRItZXYcD+IVJsjPNhEngn6E1QkXxx9A5hKr8rNLuV
lCkhCvrRs66fQxL8T46xYScHMSpRgq+BWIhWIAeJq+qDWrGVlMJYOi7mpBhOShD8
KrSpfeETJ2VmT9M47+AVyyhYIiR/VtMk7ocGgwgLETbYG+XWIJ2IZndQ1vwsd/mq
ZLKs9VeW8m4FeLBnEYVq4gCQFs+dqKCVQrR8F6UJjWdVSXYgs5flbR2y7TlP6cpb
8QOmEsVzZmXCdZleDU5SI5Qf7ad5zv6bFbXGls58HZhkrxPFk1H78gG/Ovdte9xc
ZCrSsYHWLx5ZBLmsRI4MP79oqLVDFTE+dWACllhqx6ruBm1qqTXqatw7rDx4zO/G
S8JLpzaDEw+N2HNr/+ms5P7kND2L+pKg3LAb3SBVGvxPs5q6jbzZZnlJV/+NZo+N
GRmY8+QcTuhl9Fe+H6xGhGUYjzpqbvQFiLA9aPEezyOadVooxAZYo3QiWr9R0Bcq
Z6BAwfUeWkxc18hqWFrPz7QMUvMeWBLmoJ/d3e8QMbZrzd52Xh+V9wvjqDCnW94g
UL+rLI/d/WtgXKn7P5mUAf06QsxOlAXEcNICLCAiedlfvLlNDLlpFSWx3SbbPcKj
UNDmVw/kh38580Fgi+L7zV4TxxncOQNwZB+jqnFTXuLrrCQyZGrieNv9Ij3ZRxKE
ONvlSEa8OB3FI5rALIMVP4e+YpuWGw8eFKb5r8SD5yFe697xA1TM4VCn1ZfKf1sT
U+zplpp/KK3ETIxkQvdXtIZ/G8cAP5zfrolOvHUrDJAR8ukaH09pXG49tkzhePkb
u3K4gdPQ3gHtsQz6JDv2myI0t/b4tUYeeBGehyAQsB9cvfp5jHEzPadJ8PWYXRIb
UZT/ZE55LQlPI1/3wY/2mlensJjwJzeTYcfeyq6DA+xRzCxpQcaz/KtE8b2zQDwy
HxM+CwVIHwoSrR7ftwjfu+aeqOTx6gzVE84cvY07ACBDdAs2CJF3cXnjsmVpNBbW
dAHNdqktT4YFSZqW+dFhoiWoPJAQyT54sxdBXmoUyOdZ12tZ6JMX1UqFuH9KLnu4
RZpid1XMa9eHdKuXOPpgG7ODCYP8wvkA5idn/xQA3FsSeOA7KyVZoaRUEnf/jSYr
dCKBMME8nbt27XPUdUSTPk3y1zJJL2+fblsIIIGiPkrvdvnHQPHseRFuBz1YaSFE
GDQqITNv9bxK1sjGBUlrKyIzXLkqNrY4kbdMc2ww2356mBy5gqe6PHEWNpmrI54y
8WIhJ2wnsdLKTgZ9EbPBeXsn0gF2jBAjCk/zt6OQdYvKzQJ0XG6eOoNvXkBhglVB
r+QISW7DYrLyQOHXBjurZ1lCrUQY3eroAqRxeiOnlUWtRPl3AzJxboKX4hCdlGDR
FdO8BDZFfQzUagH2egDr1tEKHdzOPblgVwYGthY+ktK/4zDPffcMscOXzO2wRT52
YHbpqxMZVFa/h157NemVdQpHdZ6EHz8e9MrLP1xFD7lB7gJaoEC8/ffaWjk34ROl
cXSGUEe29UDlrIO7XgGLvgnfTDtAnRYm8AoR7JpavGd4RpaDoRwxoEJnEiQtps/s
7Hd1mxin7G7qanmupk69o/eJNGrXVj9g8zaBO0ttyfdrEOc0HuE2gbERn5aWDsht
mMLftlWtHo8N3hs3vRTpfk2Q9npgZUscn27rJrLCO9pfCqNrXuJ9JBog8XvmZqEQ
BBu5GPt49TQ89QqybiJYMhYt+8fgm4xdUjzd39QC1r7Bvz04UFwimnMWpIUdFDRU
DprXXPfjFL5cUR6zwr5UoeTK31xYeSrkfRhK5heyYjDCTbJ6CoGlm51A5qxWspCu
+gpU+BlGeE1IIDrhNiTNiBkFXJYZoZe9Amc2FsL7bMuxfQuWPbjaJv4AP9cx6XUc
IIOkKCaWcBRGJTOARLdmFb98I/R93kRsObf9DdpXAijxpHyo4Iu/Y/21IfEr6iXB
DEFMyxBiRPmQRKWLUxI84bgizB/iOj3MFrvJh6Q29f0QotQJ7wi0aKUfpGh0O8A7
WK+gjlO+0aiwy00Q9DrIb5n3vda2WzOCMepUf9hLB8QUxuOgixOVejJsejnARc18
v+ZgZ4/iGtqoOwsrwsuFy/Y8+dQuXAboYlqIYMWQb90atlfcNq45mtUD1wGSRxpc
CD3/ySjOjXme1OnRLauwiUtm4FejfsJSvIHe0AYX1Sox8ww4vYWqhulFGlEPtfvC
/0sEzutOZ30o2buiO/G3tRFw46F1z6xvcOGgX6tQMlNezSN9el00LzUzAqBm9/WG
/6TUEM3hMsNwTcqGISb+NTZs9juFV91lrBkX/Pkl9X+3PyAj0KBwIQE5+9LSdNIt
mLcJYzKrjCDgmWwUzfkq4hHpzCkW1yiuFnV2svmxIp0EUIvhUrlySAFgM3p4N3zg
rkqHcSyAzE8Jc74cdiFupke2frxStMSPMel+N52ZhlRdOKwJAsjHxPH9E4wXl0ZD
/M5ELK/YWjpFJ6manpgo88aMXZ+STcUFu42IDgSWR9SM90kUZ0IztKi6KcJ10vSM
M0GunirPY4jaTtrB4GUmg7WTu6dg403E31ACpXbHRomKQn8JeU94rUm6fkDH90CG
17tWSO4d4LhokoFwa72PZaWbNY7ZgIKzRl8sjeOxR01XiSg/MzqVNq5E74FBsbcO
P1kLecNfWjqCevqunV32GXUKN7QRFpWyCJTmh4GEe+i5+d1XeNgTQ+0TOc1ABkVd
FkqB3Z86Qc+NiGUIE6tyti3R3H9xT+voKTA8yPAgDEkJI41RvhAShzud3q0Hc9f+
Kkk9MCqqwltdiQ2bTH8ovn/osThS1v+2pUriVLkWulgtvebih8MJzdUwYXObQqvk
2NjeFwt4r4BqiJWBTZKjUtWn2o5e4AcP8124u6apKSl1062AmcSne2C3somlTMrP
NcwvKK0yg1aoy67SVYCUqRvMS0DE+6e79plh+c5BoDrqkq8+gR07v+0q1mr3yLK9
t8gIfHQD6yg8CE2POhid9ianAJ6XbnIbdsP7YiXANoYnpCiMP/4efGICaidbVsyr
vYVOMbonL+Enofm5mqSIuBkr6C4NQSniLe+866dgbyB6rNcUpJIwp+cIUtD2H4Kr
4j49k2x3+T2oCwSd7jGCyQAqlkSFGPcrTvr7S7WKeom6IuHwzyuZ2VdWyI6yniEN
uzwIvBzidHv4zc2anPIfEsQN4PWZu3tI2jdhsMJTkk49jti+nOglN2Sg6hbSwWyc
tuT80Km2r6cW8yPZzZfGVhQ+tirHZz9TLPNnqe4n0nVLWbf6ne/aCmcll0cOUeeW
dwwyGWFl7s7XMl8DMyI/Dx7oAPQhyMU/flQLtEhU0LQhNF91LDH52uKAI2mlYOT3
9nJLi5UBqwoK6d11qd+E/Xqo7aSACC4uwmaoKXBOXHwa12YRm/MVRLHhqgHaaoRl
nDM82kUARRMLPCaeDuEF0HuWuRBGsBnhdhLOx3jl4sWWrjkQlWem/j2Fl3igYnXu
zo+Qizy/1cpb8INpMFR3CF4Ola8itC2aOlat6gK55WnQkk3MSnFeEEQZojv/UvPy
2285nb71mGP7gn0ECq6GSaynOYoAgUMOWJEWRgQ6mn6+b2p5jpAAOi4VTH4bPfxd
sMYF97H41KdYcAn0w4pyMPBthSpZ4lBnaApdBIVec1yKzZcA7MkdbODODAnW2aNu
HCmQziud6MmmtDgMaQnF3xGX8xve5Do0uz1wcI11cvGocvq/eJvXS6Bc0KplJ/h4
EEVkALGSveERW180PiHTYKZ8238BkZrxlWPHhd/x9xN6UmcrJunZILug+qq/UUWh
q/f3tq8hhFMmGFnXrt15mAKr8QRn0aTznrl30vZFQwUXcrsRzvFkL5Dybsk/Jfzy
peTDozcbdwaLletktHMpn4JtjgycGrVIU8dg7wfgJ5VAL35YsnialfAJSQZ5cFKE
nslbBqd7WSIgk/e4r+YDkuyVyQmmiH6+d8gy1uUPCsuAjEFG2eyV9ePf3wlnX9lu
ijAIVZA/UYhWrC+ksH6ICXdgA5oMMBqHXwOZ68Y0rWbTPGozMIBfH8PvMxYHz4Ux
TbavNnFlGbUpIm3bXIXAWqghVhkl0kvET1zk6C5GjK1Evrvqe6kEZtUvBaZtAW+n
y/q2lR71t1lQpp0ijkPuyfqgCNLDxcyEjA6a5VVnonbvx10HT9iMDCpg4Kojoxa1
XBZqnE6OwrzDL/ozvheB8Bs45CBRXyiHy9l05zkvyLxAHtNSiBaURey4Xy9NVIPQ
JmZ0iPjR40fUxEBEiKsZ2/7XPqQScR2a8lIVFBFdD44IH0waATpLxNTAGNXZsmrQ
9urgP199kSV79Je7BoS/RKHFGtEqVHFy6X3Llaix0aZGe3Oum0RuqNbs3pLSzBrz
ObymLeX7eUBDYm5RZ4H3D4bWdU/azoh+7/ZLgWyBiAEo+1458OvdwWqSzILsq0Le
afJk1HrjO2ffmDCc6yhQ5r6uP9aWn13Xzw/ESNdnA17OuLHZDXwZCMzrUd+5UT/x
qcuOnNKrlEV6iMO7ym0+I40sb5CugD6dSKgdqMoH9INW4MmoVOC4iGZ+c24RA4/b
03qJP0wMusuHUQH9txwnYhfdEN3AWu+oDAgMg0srO4b/4wu1GPE+cXdoh963KOvL
cOK2yXf08Wyrs5JPjT8KjhogIZdKRnJyH9os2DQJgMbXYkzJVvfvd5S4xwabfrmF
q7mEDZmfs2KiAUOYVL406nMHoSZByOl1XDPzkHMf7/VQwQ/GjWqtrz9ITcqch9R2
hMRSGPeKR+GthdpcX+VJEPEnXYYCyTIIetASDCDdr0GpSW8zlV16Xa1FmnByeOQm
xDijXskwiISebGywpfMDHKMMkQ+CX+mQNfEUdVxQ51AdMvRmaJdeqUXDWLxMWlm/
XOmaEI5juqRbBlLgNX3bfHV+VQEK8FfuZv0zN7lNhNox0a27aPOEjwTHSzY7tOwe
+aUEgYSUPqflLQ88Hq+23QDmu8uW/TfzdAXZ+Quyy2aHKTsMbUQKDgW0TCmTtC/R
rax968uOlXVWcD9WgbE2r2jb4OMYH0qXp0mE1rNbXoySuvF5N3VVo3Rkz2rac4Ok
bAZanJjk8JboV9kzvuBmrQUZW2DsmI7xTDI3+OB34y6rfXbtZvuS2QX0eB3dVU9l
Sn5NhmHcvVXmKFBcBPKql+vXAU6QhqKjzah0e6uwiv77CwXmYpY8bY1d4rp08l8O
Rmqj5GvnPVEbFxlnUj4ZKtqfAVyVTsVKV6gF5D6OZgtIVtgJDAWwtorCsmtyR0/q
Qr7YDTtlofyKvw+suwbUfroXkCGFKiIBEmbbXl9u2NSo8eYaDpadya6n/9o+Pu5e
oNuoogwmP1cH2s9s9hY/GaRh5UNPsqFY8+B8/cfg+OXGFPHW2tBExfRwyqWvexSv
9ACJpRDrQriqp06h5Gk12Cg9u3vpwT7M28jqEfXN8smh2gmh4H3H7sxQ6cAlVqoq
5J0DLqVmpwhL7R850O1n54pKaN7rlO1NH4H8xEOj2pSXnvaU5cIGGyV2zhAQ/ACy
POqfJljCLNTA8JEiEiELVx0AbT+JCHVUYvilREub9cdkVcy5kcL2GFRchl1XgLCt
83bmMsLanwwnAplzBmqxzcNMyV3S+Q+9Y5BeYsg/xsWLeBVESNTNuaHUH6L5oAIM
4DEqHCL+Ss8Mp7uJDFY7Tak4g6RhU/WN6e8g8uZY7QxsURhE6vs/+cCdLTD+9JBm
A0g2I/xNqM5Y187cmZWHFUd0XGaUwvWH69z5UL5xAtTyZJAfjL6aOKdT6GX6XZyi
nCgrwfFQl0XV/e2rOCbvEDJYdHtdQ0JXNAdkiEemGb2K+fnnvbj73U2xk7DcrEjp
nz5UvRIE3njSLwrz66yY2284ZZjDRU9PCgC4iAJy6Nh4afZMAP7JB/+CNDPQaZiZ
s/+eepK63CEVVhy6ZI3acVKclHJjho5RUFRrpF9h/DyCqAxWTjglQmZl/RnJtO0E
enjCNwzz6P83H/NaY3Mg4FOfX5lY4zvqeBfLY3N7O32HmhLBDACX8UiYO4u5fZ/v
9CEJhY5jXJSQtpchXPw5ry/CUwYcUh8Xe1gGC/uN/sh+3sgq4N5vgsKrQZ8Teg4E
gJBYo2ycW5SWx/cajKo/LV8L/E+up2g/7ZBbLq8lXqgJ42WOSNCHVQkLQ5s7Qtt6
mQhEwNdWD1bL3J7OOZ1OkCSMSMHfJ8Sgdu+VygtOK4qLuV8pmn8WnHPSplm3vbNn
0lRUKXbLwgcBcFZZT1bTyl2gwMFUuaKleRgNa2LpxbsEvKWHaiDeCj8q7lwlROu5
VE0oOW6rWB1d0BrfZGealGjsSVnDAH14RVrAJZW/glHY4+OYyiSv0M0EgJBIqNVP
gu+ITlH7QzxLFbANPHO7nZ/+L7SRVPco+aoPMNPWAsPd2D3p4yiO3uxDRNa+tIyC
+OWhr614xrSZEhgqjrysLk6XrP06XWwL9lUCrfMnbI/3r3lyIgUvWxQFC+2i8CD8
hbnbSLnkTd9wfzXSvYtqt9TZOgbD8GbV/Rlw3rvGjsIKooUhtt3woE+B20XNl5RP
K4lC21+Nf1LbjrWsez8t3bpCN9znBFRmj+9a563CbYkUfHRTXh/SWGgdmTnLv2gm
n/sPx9f1G6UY7vN8QnLJvqDseFWH3Dcl7YHIySb3fJ0EyntcOplq7KzPgG27cFCt
RFn9OgHc3ttSNBS7LYEEAcGsNtPYuBXOviqqVjXN8ugeqlQIhrQrGB0j2jnQvI1Q
PMToy842LwU5TZTQbztHXkzrQU9zDg5d9UNuWIWCdgNu2odOD3BvbbE1A9tYVwtu
pEKODjWa5z70+EcCAgT6L4UfKXTXd5ReBrhzzyYJ234Ze9cUB2unO5mDA/OgU8U8
Xlcx0VbVYWDbVJPN1chTQ1I5JkhFwmJkBbO/pYUsf+Vm12Ylbz1v2nS73H1Ylhc9
LhxnajRm2WUJz0/h6duIJxE2Ny2Cus6tE/pq0IFnFlnCFCci2Q1StH7M1kht4OOA
yYWbJu2BX3DA/D/pChDS9t9I6vsZphBVs4yfvL/4HoavhLotgEbIeu9nuGKBSWcd
RMfRVP6RgAPqqNDI3nyToNekUiPzYNbshiUk6L6DE5hHa6zPEu9sbhWRIwzPQq8d
gVmF8o2Ly4YhqV/GD1CDTwZarb+8XrMi/xGMbIzHrSYdC6rS1RDfYAquM7SZHChF
0keMfBtK3TmUA6E70bEJQkFixK3EFc3V9eIpml5RX+HzYP806yKRpNnbLnIt5bw7
Sqp3zzDUSLCERClqQ5yb6UNAnzX9gy+qRWfNQo/e60GvPky6MWxWhY6rRE4YZcXY
o7aEicvpkqQOjpOfZMgSAwScupmYZyRv82ZZf6MY54mEMva2I12hU29aREVAvEfE
68Dzi1mvHA0bDUaX2UWcnHgYrIRqZ+jwyo6XvhFFtY0Z95dH2ElSb0rgSUs/Wi90
0xarFNRjM7TGSQXu0U4vldYJfmwS9vB/DJd3l2FCWeWbnlrP2RkEb+swF9QDa5AO
j8F5v4zCXD157BurjA67ysS3/SJ5vzpW3XLWCZkj3rTd1UmqiL4csWMkYPhPVEBT
e8gdlxRzAvro032P5dO94z2JQVFzS8o8nWKE3+Tt8AEvvU5VLRR/fh/4XEBtxhnW
ICNNoo8syp7CifEdGNN0kSvC88eX+WTqn2QlUVnQcEIaftWqX+1HdDvCOg+AEKvy
xVFJp1WlL159dxoP/aTkneJqtl9bRDPE0IsePfYk9SysQ2vYzT4qqxlXhKObue4o
vl0m4BSNV/Zb1aHoKKokE3Kd6k9iPYztItTGrSr3oi+S3LiynowlVRUYoijekGVx
Canyal8c3ySaNQZLgYyrG5yhs4YRT41tu1EhpshMlEQHkTyMQedjilvsCRJ86xJg
+XVtRUmbZsoJkCtG5QFtld97mjkfiej/FfVD8mpvwFmT7xJEqmOBh/zbjboI1jUz
SagZet9BwKABnmveE6hp5/ZCS11SvVphpsMwrHnTsRWwS4EZKGhAxcA5fKlUi/8s
FEL3AH2A7yeXAQoWhckz4CbrLoGvIVpQgkVwmVhP6KWSe8cHZGAvvpNlSJhIybQw
MVXXB54ToVxOJ3408ZfeA8GGymS5Q5j7mzBLfD3oQpfH2qmOXqZx2sTeCBysWNEh
Rd8jgxfJ00oFE7oZ99ZN+6DS8oA2XITDs6SNwK7zxDSWsNK52Xq1ItbhnCUj8GcC
iaNXr2JDqktKS4zim8fjccypBzi/mG84pnjGY636gL2DEbYFRrdZfKQb4jbsnSeT
+Q3JBfEoCvJPH7FFGZWA4lk+E9rCw51ttrYvQ5FTS2OuAurFWC9fYhJKqqz1l/2Z
BPkSfsqgeQZ4Y1J97PYo0N5ke/s5IZILmw63XAryEUhMJz43xcERBdI0JBYXaCh2
WzqOfhGkqj+P8UtOFsSX4SdgrEmj8aNFZzUh9yTmHUskTDRE/k+6lNt5xhgTRAo9
R59pys2jcmb2XWpHSl1nou77S1vjmV2/ldAKc1on56eWW2/Vb1//AZpIBl3cICSj
0haJT9BqvZVQqHUbEoZorRo/yXbv0BeApA7MGl3Ko+2xDB3kisonWIAJ2nglKyXq
zRDEVFfVFhPmK7SmNEIqsvlXELacRdq83fdlvYfQbsiHNcOANyhqikiDFerapHXh
u7h1MmLXlheWi2ycighB3RGC1i8tZZq4Q9jWrMzdLe7AFIKnHiO2JEa80MRUV+gr
A2VSbDx1qujNXkurgy4WWx3HarfPmdxsNoszqbXIviSZ+mJ52dtj4fvgrBWbgYsR
REEFHX9sWE7BKXOii7OTqbWTVlgp+9kxGWFQ9JB5QjRaKyacCdMyWPxRxwR54uXw
90VT2WsLp9CVSApsLGLRi4/tm3XdLISyfqsEDKUfHr+bMcbwLF333XuXYgmFN5Yf
1TcEbHLKvvvkvDGgV6wq58xCk/oGy/wGUF5QhhVdPtjO0HiaDq6z7TvMzV4hak2p
Np04vxzImwBgZCF1b9+YJSH6v63HYSzAyXdsrtzReLP7gEekpQQA5DKaCUlHGGwF
YDiOjw6RCv3lFlDMpTwkzBSHCAaigvWHT/k7v+hGQbCIHtAPDAPD4q7cJe59fatS
vyTZR9EYxjRmjhWzhbhe5I/JbojwQTY2gdACAcqAFqxYr9oTfuT2Gp1tEH380WpE
ANWim/ZsyAzEbQO4l7jtUn8yS2cVtk/t2k4O7U37+8OtRSwy1yuAskIeT/z7KxCg
//sSLwpSlAP4hbLcrIbTarkzvEDxVxH0zUZsXU1oUHIGHpX6t00zuWqEwVxRJ+hF
MALbLn+81KBeSuiFEGq5Rncy18EzpQmZrj7gTo4gxMZ69yFm23EOF/LLBFiJJgst
LhU+n83kHU+PUGXlsZ1rFe9U9Cqc67n54jTj6iM9KnctiNmKeKLHe4ctOxCaIjGF
A+WjMetZ7On4C6faZFQc2rEWansz9lB3kniJosMcGZFQkK6lV5W5CcZY3oGOEi0U
itC7hG13qYyPm62l9nMGCVvVrSSbeYm6ennoLeZSaJ9h+pSCIuFIsqQy/nsddYhV
SX1D6JfCUpCXbd0OiGEmMXU7HwglN0hCovqwtfmLMvQqjmIUzc0OmeJld+NEGP71
VRgcdM7f1oMhq+0ev2oYpy3CbNqj1SoEofgMLYrId7p7IksWxR7HCS4q7NniAW1+
J+lnb6/W7WUSZNEy2cmZYb/nuuC6/Mr5uPVOH4uEV0AZ50bBFK8VQel5Ar25uFKq
GCCHYm29vdjBQHVpQWid0vFzs7S8BuXg4/7R0LHfR46p3BzfrldW7/lW7oB+o7OT
kJkg7pE4I43S2YgQywcHPBgcQvnVRGcUEmoJGSEwwAfu1SdybuQPs7qtJc9U13Ie
9a2ifmr8IFWpuWMcIGwLfitinyGq3SZISpwLc6M8PRDObboYMw4iBgiJOANEr3HZ
66TI0Q9q8qIrf6CSFjKLi6x+E6fCveK44WtzVEJrSxNbpKLif+l2tDhuUbQXpaSi
kmTmyIbuz8/gYPX7ILM4QCxsShkTeWg/AswNjTSkRbQkqKGTDUtwL26RcisSQ1g/
E5dqr+j4eGsfIqNLvqSxQtcCehiPfazb9jUw+PbvSPjy1HzTexXF43wayIh31ueT
n9x8Cq2WzfJyh3GT9iBEZ/KDC2ii0f9eikl2JbbDFQZFi71wWq9/O8SZqLBwUQ5S
tWA1Rdn8Q4Pwb6+5afYE7cD3t3FykX/h1wQ2CeP82oOrAo7PQ0g60hLcLEqiqZ2P
MJ+7MqQ3C3dezPIMWKU385ow/pBykEz+BQCFLWtIHWLZqo84sb82jUhJBDDoDP75
X7k6sixeKrdsY0tQSKHR1YRNvYGPxygoelKDTGahNkjO9lYTFMWyHx6YIGxvVMwX
vw8fvMOSTO+oY0JBSz03szBjOWbfsLMGr5iKHV/JjVgAAX8KE2Imdt5yrBHnsfl3
BPCcz8Lqyx4pJuEVYaU2htt4sjZ64/fSQ0Vl/6QcxuOhcmwNIl3aQmEmRM9QQDMg
q2xy/PFWo5yN2sruR1ye3b/DAwAvPQd+PsiS21qPEt9fly25Bt88KLOzT7DFuuCT
4v5Z9a0keRAmK6Z2v+mU53YJ3TgKR1EuSYdJhBYqKKlwJo1PKuFsdzNrK1kTImYj
zXW2dOVT0U8p0PY2IGcbeBcNIPpo+jhM+3XKJfgDFZAV2d1wmPrkbfV1YWFl+hke
3ioz6Ep8AHPwtIcqDAeYEPIpEYHoTK+FaL+IVyyaoPpVyDiP5A491tQUWqqM35gz
0aWffntSCIZL77H2mQiB4JZnbkGTXaV9o82uiob3v7z/hjG62QM32MQVND5eKNp4
Quy9nmaaiaonVYMEEEbqx7430wJaLJbQxLhcJHlj5xlx3Nk//QV7ShhmX5+b92ac
BLPhNGLVCRIIiE8xmkkSoCN1Gr7CPpFSVQ6TaufQpAg4trxqY9wYEe7oklvZeuS7
9r4KjKHPvELi56rHwUgY9PWZE0sNp2hwOXQMczyolViHS1kKscEG8TpQ36ypGjYG
x+GvRs2J7ablL+JqbX17nmmqNt10taoCfvlnA+rSkwVcBV1wZ2ck4IQt0+P86Wns
LRT8C60X64rlKwv8pLPO4nQ3s68Lo/tcgp36ClHSActhsEmA/BaSlzfG3lU6TGup
kFmRWUxw+ZiQjmh+uIT/qMWQrarqibCwUTmBZvZnNF2ZE7Ey1rZu/AEXFhAnb8z8
Wka1j/zj5bo+SD9Jgj3/1fkR63ACZfgamMy9cc/i5Mbm4djEHl6qX0qepvILVtgM
EWafJax5mCjzGUAfYa+0xo1L0Q4lpqppBHHjblURmB2EHLL+vc/2YgzmQ3ri1+tj
D7v6wozPoDvqQE586OzEWQsZ3TiOFioPUmJh6Bkn8jYmeez8s+4CFmN9EqoCrSBA
tzfnia56gTvIaAh4qY23RA5URm3a2hpb7P48PaGRuSO8U/CpY3iRhcH2Ei8rHuOW
p2T4zy0OMArj38qwb5+qAOBjv3Z704SwllVHmrMUfsRGVmuh8w9pnA9WIKTvGUgs
w0b6w5NVdlNnW8y20D+meHSgB2yrXrTeUVFUL/DQC0gdY10Q7ez1lSssasya74B6
7RVI5ArgsTn5W71++jnAFRyv+H11CinCovkZUGYu7xUEIEdRd/YRlwOgzBjlA397
lvNl/rqxaiNiR67mrAsM4e7WCCMT4u6R98QfnkdqaP0DLlT9WgiY2ehRwtsL5y/B
/xv0U+WkpsmpX7gJcbeCbDlubHBwDUOzu0/ABKeYv3x9aeWp2li382JZjMsUNz3H
umzlaz59V9lcPNzIfbZjP9N3caVr/fh0iDTr7NhWH+QRrYEc9//F+9rpoz6wsG8Z
X5QU/zViUTTVO6UgpAbZ+NMDYyrB6yxqQIZtdhkva8SK4E0tXxpw5sm29K/5Bvk5
lSa2SezfTdSV6eO43L10xFokjUSs1zG3eqlPTnQBSeJaVd6wPLPN4XngP+rUSEx/
g/LXG6MI+iHG4kbSB62VXbGkS30D2IwUodolJjCDtfgJjT9jOIltRTcRLPSQ6Zb9
8NG66hJAyT4DhIuBztBmuMWWWrJgOw7EomvAmp/3019sgBAbBPiSPIKDJGKyoq0A
E94iRvouKjeB47DayUM+qdZi5jSt3cxG6ALzYQFFWD9agHEabcb6tlKtmhnBYv7d
TXt32lNGlm7iWH0bMvFjbRrTTsJhKmfSbd/dhcGf7ztL/ef+x+QTatS4YFId9n4W
nWMbyX2hBmgEoF30gLRdQM4F/nFrYH8qSV33IDzEDlwSM3vsDOeiNAzneBwMEvvu
s2fz3DIh7ATPdhsRMpDPVQlo3836XkKQyc2xH8Esnuq0c2zys06b1kopGSN58BWM
W/i0j0CVMx54n3c3tILEHSRNdDJAHzR9lYkvvcTPDKB8QtbON3+ILLjSs8o/QdwB
n4tLCDD5dfSb+qBo5U4owVnfr03Igopm6aBRBVNygaCQ3AKakEh/lbM+wpK1kWEh
dkahdEwBo56ZYrg9C73jMC61oNH2os5J2dgrw5i6Ui5kc1MReGpef/QF6J529rqE
q32hWfrX0llymAavbPke400c8uug2sAWGAnjqDXXIMfdWMTfjiFA+/mVAgyrnKxL
yDLy0v2DVoe8G67LtdzXpRW/lAPsdoypyStNwYqPyyccWWCr0z57Doxj4JzqDI3d
CbTL73VhwiEtHPBo72WNSak27lJEMjJhid/sgZpuLTPz/Chdn2oN9uD3czcZvAVq
s/8s6UBm4NW7wnxvEkk3jWkAUe9ZkNmNCwapF26BKTHLKR2J+WImv1yIKdgAWbCv
EJzEEj5ZKOsSeEd+fhOn4DQo4XkLO7C6cQdZ7802GsrY6T8okJpG2nIfUcTMMQcZ
YIQbBmMyeb53/mx2O7eHrwPkhJhCaKvrBU3q8LYNgEFbooNF5G9kRcWKozqlfRdh
tMpjgZ5gvkKL7MnxYINf+V/5gxhoBlV+hRqvBAB86ovWs0rX9GYOyopZ1C1jasrb
hohCYmjuzZgSk1XiAVipCDMgxSc3xce4gPDrVAV67ZmQ5d6hRTnKvXoO3JuaqojC
/hYANHxgORBcKwhyeKjQcpSbsJOlgv5sYTqak9st3LTlq95aLAc2xysLK11ReIaV
W5rzxeLxY6JYrIW/mG4q7z8ImU07c2Gsit58dryQNoEvUDfnv2w3NMKcaeCHeWC2
T/C4S2o9yXZTOLj5U6o7OgYK556ih2Rx187jGLkpBIvAKZxkl4//lQkd1aOy7bPf
XoIQD3BGmt5hY6w4CnSji7nez0PlVRZQFx5ecYnTcXGYjHYSrP13J+VshN3E5kkc
+Qg0aPka78t1jtPR2l113xrBCCaZIDSoe+YaR5bBlM0hvCKc6D+Ib59Fdf9kkQV1
EHX37Ofz8FfiUx74iKJ+u29j0AzMUIrlMriwIGR8ZrRP7VHeXS9mbYDjYVIsCD8q
I1TgfAjkPveCJjcZ3pMak3lThZbPrf90XQ8UJZh+cjKizdZZtS9qBS2vJGqwEC8r
WZF3oKXRWjsg7ryXVamu3N3GVvup96/4L1i+ZZq00hu5u2JT01945YRTy/jczWo4
RwpQBNgz6/9Ur5x1wA56EkldfJfAkzze1iakF5y74w6sMmEbrLhzyzV2FP/UgLXz
NIjTXBLA5/2/RtxRGpVDuOSzNngwsrysDTSup22CmSfa2zxUw7G1JFBp9CRyMG/7
SXTWSvN0L9ag1wHm2mzV53efZ9BACuUKhn9+Inuv4GQFEWkK8tSBltDgigkfP1lp
s57R3BWxng0fhGRXdM7dS9qHonw4NWuG7ycrQ0kNlK1y2YoEIb1h/YmVFl2rWczv
U7Kws8QT82qMkk3HUX+A9qEyvYAWhaq4Bf1LGlIfw+OtLh5vo4GkY8pE2mflfquM
qWUcUdMU52Yvu1o27vKTM+ovIdqAnl61rI2IYU7WwFoqEYhwKHbcaSMBe8Ln3HtJ
opvaYXx6C70BUY05UVEImCFGuOHSW6BkVlDWTUuVgzWxAHCQdLIXZACbxfRfKanV
8Xpb7/iJfyy6ag7diXdL92JtcCpQpFBJ5eVeaHKLLl6RLxnKHyqdxtvumnIm8J7p
tmw3GDynGYbHqowxd96UpaCrpS0YFkTllZmAioiKSZlnqeJE5xfxLT+YDzglQbuY
j/yWt3Vq44/Z9GCgoidwa9uJBjLl3/00tSLRlD6sVPze41zAnMr/Q3y+OuoW8O9P
BO3TSEbFR7BNnfH5iiZ0zZ4vLkSJjK37xBc5IWN0FM3YUWeV22jT6emM6by9H9F1
lXFIy75SIkRUjbbbrbotfm9OGNV1jPixOfroV4gc0WO/psEwgCkmfYclJq7cpzWA
m58SSenz7wm8oU7lp5FGAhK8VtiWf6Lz1gN9qvJTJY1EQLev1H65dOpGrKdIMFnh
Ao6LRjAIomWwEWBzzXuMZnk+X5K5MofLVMvYXUpWqiGq6JwvA5LLvxmmXSeIzYv+
Yj0kF8hKtj6gsNLckd2aIxay/zqhSEsELzfkr+MPwQpXVHw4mDmMy038RQL4xwvO
4BMTLBjxu+5PY/aiE/33vbAGnkGMmy8Cqw4rAItlhDQY1gtRY9ufjgOySilNU9RU
00bIQSbCxnhQGWpB54pK+4SCSvJ6xNVAiDs8418UPiT/0aPF4NI1D3tSLxg1SBFL
GYk6g5geAmgO/t886BH0QeGo/Mlcq91xtcZ9RCII5dy6zOw0u4Ouk3nrip+ba0VW
3TtR8NLrBxdMWymgdVdFqnRh20e5xR3Gh0Xi4uFoz7I4DxVuvFSIdvpg7K1O+qmo
dboJbUa5oCHAOBK8kaJf+O7P/qcomJgU1fOsyxFZEYPkwnQ/ZPwwNViLgcar5fnD
U/zoNKTgSdCR4kgAv999Qj5IKoQ6LwKJH47anVAeJEy1Y5EmeNzh1KWIJk/BLKJH
JSwzqKTv3tCnYXTHGOf6wDm9NLNw+EOpium0I5IBcpLD3dsaZRulRa1edTtJLXci
Btpm4swRj2ArcQDJQNOVr/EJiDM2qzxtxFep+XjdlOJo701GXvgXt1W/p23WQ2+x
rMrDFHC0mygBtuaLJOap9PGmr8aUd526x4lStJXRklnioswgXt0aBartOyz905Fq
0b4qoHxHNHzQbVSMRMbwM3FGr9rHdifHP/+cNNhX1UKHQrc3PDw7Lv+juJNxVTBF
h1ekgdYT5CY8soG8/+jiyPH9YzEAsYNf5qfWx86y0T+oRHt/Z9jrq66r6kqrp0Vp
Pyt8R9MXKJ780DkiWPor1aVVLDvZoKdBavnMw0NMgnkmYF1r/KoS3Wb6DRJnFFua
aJH8S7IlGCbIbvoTLyln1vQ8id6YX69rqhSl4DWtO1+8dAu+56k0h9tTFrxvTRbt
IZvp1M5UQfY/J8ow6fC+jPNtWGlfQLaSqZrQ9CiasZe9uux9hqusHiip86xBhQS1
dQnVDnWprGPTe5pfuFaQdC/jDQsUGt4t59h9Vdau7Jq4jrs6wLnHbNLUqt7KH9Mj
rz8zsCOF1Tj83539O2bL06xLdh//aH7lnDuWx2bW61JXQKuZhLpbEd2ydwBcM/g2
De+z66bmAO1hoBsivWPKjoy5cnFwce8k1LeoR/VC/0VzXhMBb6ck9e0B0KAZKkRI
m2Ktr7D6PWSmNLNzab+SZnrYOZdn6vv/E/KcqBCyFUs3J5w0rJxejzmHy1oTzKT8
/rAa6IaF+TiMFerVi5nJtd0kS9OQYwOvvxtHY/1PdUb8PkP6mrLLgHCz9bGSe52G
JCeI0W4SsrvuAOF9KSBm/R5bz4rOhCHUZ1pn+lWi5It8ljlWt6WPL4DxZIl8NSUB
bVJcecWU4YM2BCJu7sHpbauearvCWHG8DmrJ5yq1sykdc2JesF/cOUAqNFc+aiN4
5tdXYNQVtgtdhKb0sSZwDE4e4GlMwCoenC5U+A2ImN2jbm3S6q9Jafyhw2eUXceW
+VP42wKMIEMoQDdD/XpYEA+ZXSNrcoM2wojvgzO2PebBxbweQKLju+Gx4BX+Ii8O
Lp4EzSR3NCCqOOwQmA432ck9nGBDlLraHIE9d92bcqnYdy7bulEoIEun0kJ5zeHH
SnYHbfXTBb2ZE/bD1rpdVe+pmhvXzS3Ah8gmedeV14erFCR0UzsDnIfgUDGAeozZ
OHHqHaSStH1mhwpQBTBHq/od5oz9SDPXopbHJJshAWR9sQrlRsvlk4jdSorLLGw2
+LjmRf9h93sR1NHnJaNcsTyUwip3wjTbuzRA5jWmbr6LTYWZQ0vv3wK7rSkyFByX
6JozucpdeNwpN1Jm2qFYPlAz/DGj777SgevRfNtpqb4XxJKp51R6xpHD2p78JODQ
hMWb9NDnL9jBwjY28C7yVXUdeE/u8yeAWNMz0GBVZa5bOt9a7atyeSv6NzRvKzJY
7vAkQ66QcZPsDN0x3ZUBCSa3olU1a3fW3QmGJ3iXjflo1GnvUXghEIR5VuXJvy08
0fvBdJgWAF/GzWSYCFcbhDCfp+Ed011LcUIHPTIs1IBoxD+5EhNW1QhxkufuIyE6
HXctMGIQq0WutFrnC9fdEVACgzfj99AkLNLSLAulx9XAQSnBNEtSpyPM3pfcTM03
cZBaDLHL6E4eDWf5y+fqJ97xkJieNoK11mVpoQb/pqxasIqIYD3pIDIGCzKiRmnH
D2iJLv/QGvjVv8uIOHuupbb+zqAm6SbTf6rIePihMCGBChpo8SNoshg46n2Kl3Ss
9NRG6+Iuvj2ks2Vzm+x6bOjBRguuiNk54BicOKEiyiGzDAhETvl1/5ojSk8rKjDu
DCjYKVjQQy06Pekv6uePApwRixPmcDqcwsyfiPQmAS4CZGOY5U8Og081D0S/QUS1
0X3ArqDcYVzKB3oF28cPAUGhDhvWrJq7QTkYolC/9RJYt1f0q9ka40OyZtSC5VuD
hha5GbMNt2NiukbCeKWarPrEqiRkCCZCQA0nlPKOa0ezRxqYlnXsMGi9T7Ej2+7f
zSFYrViIcn+2cUGAbU4/qlSWtTCVIllAa58TnCtFdvIIU9nVBQ4+iWk4FpRJeuO4
kjaQc6cLFg0H/LIN9+0D0VCHGSQXAaRidguLH8kqdxpwG3GENf18NgY06oKxoNQ3
gnwr+UbMqFgQV41Cl0974zHSE8rIHRM4TeqODIxfxYTZ0q4PBRcNkSO7GOq4QOJu
EriUrrlYpSughzwcR+sMdFH9eTaQmHbL5lFM1HYx7PA4DuyxGxfV08gBjsqMMcTO
ZXFk9t6C2zx0oUW1rOo5Xll+ZXZM1R1GYKyt3dbL+BOMKAjaMzGSUbx0DwaJllwi
Kq1YUQlWGP51yfxICyrnVNCSO31F1wStauTflXoDpoL/1rOhLJW4k29G4I20LPSO
FNFBqN62vLKV8RBb7C2qCnHowBS9/tnSquBOIbnHTa3gvIhhsHtn9DXk1IDpEhEQ
A8APOamXR+1WfU9KTzAKrbF8v1LZOF3aOySECv+X8oUedZd3C3l/Pr/JxGW4ajP2
V2LlJ2A2tyxR2k2WRr5j9iuh0HkXmacOY4AcUXjYHNK526N7SPTMTIefj4yTUkr9
yHVYt+vvA+B92hE7IyDX/s3GAjPPZPTU4aTSFFC/P6o5PhA2VflIsqc+ORtRJreQ
g0KoyoDQTz2jGpEiRc3V+9188R9q8bxBNoT5eyUmq1dc1TxpDpiNSZgLXhzF7/qc
qobUel0edArCb964bUMuGaakgZucILYYmt7WCjTw3Xer6KlkjD41nUo65bCGdYEL
staq9KvDWU90ORJ7UxHNnOWHDP9W8mXdKF+DZKYe4ucTcEJzP+NzTCzzdQWGNpKl
5nuZJ0jFHQ7O9kuR3lPtg3ggIhauR4y3KypnzCVHblVWZl1rsI5xjh9z1x+A/lAk
2WjhwQvfFF3L5k0geDaY597cQDi43Tqu5mJ4gY15eRceVPOetvFmQdHUJgyX3zW5
+sDYcIXU98/xK8/xyDLSFOJfrSHCGPSAga15D+L68YeJCnFxEmMWIAt2g4r3gCR4
KezMrODVQKenquphFHxGkqkazo75yg6ypoSKvnfQ1LumtJOyMcT3WMHFHpAJvZH7
s3CIqmNqSKMRq2ZHI+GuyeY/pd3DYpn2Yalh1qby9cm8UZfOAsk/fQruW1/ip53m
/+l93oB2kb3OonUXEAgf99C/a4r/WpWkX9ZBIqbyKTKI1GPLuwhAVttp+IuB/BHl
EDNFBtRPnWKpcDsGUWuD/pMEHKLscpCoXEtZrrE+YJKFs8MNiGmj29BHWUT1ncCs
qV5ppImhs70C3VkM0S2jPaZLdK+FwgXttJSiDbDit1zv3kqmlaX6zFuKekCcFU6A
Qb68847OijLhvNkyItQJYonF8851gsOrL7rV4aZpm51ph5r8sEokvXxK2rT1n1WC
qZ3ECW0aSAEa17htmmbjBLgBlvi6cA4gbDGTbkhmYwEHJxdkc0tzo0fDTkW8EW93
eNzIeqqqAp14Aqp1w/jHSZ8TYpiloGHXP2zSv7R5P9s0KC8m2Hj1Y1HaAIkwccYX
zuj98qvYqRy9dhmqGtCK3Te/LyuB6XpZOjO5K/eNJZkRioauO42JTG1q/gNW/xCy
TQcD6nbvdUL/DeITsDF/R3bQnJIXsPCe7F3HFYteEiId3YlmZ/yKZKnOp75A2Obp
WilgGkOnwIG+V92g17krBat/tFXM2zF4eA5L7xEHtx0RRCSWwnopTObufB+Qlekx
2DjHO2NlkKiF21lhAgFFn85a/YQgbymkFBTN7c/j2xMGAXTFX+thSC2EoW5pWyGT
yHYVX57YJo4IbWFQFUoVfHDZgOviaOc9ECiaoa4uJKNkmIfIP7bY+8Yx40XMVfz/
Ijbp33QqrX4Fle423jJUBiNkkNI0xIiELEn5calpFfETA8BuX8NidqOqWnVyauWE
MlzAe5osnusWD8dt/s0Bm8qvwbmRN6ihV3ehYBWqoD5XucUeFfL2v9d6ootEH18+
lhtEaGBBzflv5VfF8VLkLHkm1K5YZFoKcNVXxK0oYIXwjEbt0vYqzhlRnj4szTnG
p2fjmu9jM/B+r3shK5Oe1nplhm1UDsZHfuIn5E1jFKBIjqvnQnk9aqi7QUygt6ZY
DRNjS2SjYSi+tTgieTFKGFG/aAiG8kkSygnSTmIwFDVXFQ6BFuVBMemPIaS2SfXT
VgW/sE65d/fokBhxV+omQlqi5ik9e0zIXk0ctwSvyLMTqQX/LG1eFbd2wY/PZTWF
Lw7aVQFAbXkspzwMk6wM3wcaRdstdXtdWkFBeEgjL3XuTTLaWtYILRHzk/3lNEs4
vvdxBR9ISGUytJBA3DJV/gXyB0lRvI0+nH/DiMicCcMI8Z1bjw9fRbaV34IkmiSa
OoFYsEJ3z0ojlgfWuPUFTJ9g4z6jvKMglRbxm/pQdIaOh/JkJ4HAS+uIzqul5VVE
zy+htJ9mB2OYCra1DDzfW/+BlEYPRVQ2ubSzO8b23hY8y7q+Iq+VDPMfouKW6EDC
z9kdtQgkNhs15CbZ/JlrPNOOTSzpU9+0cxxHrs7KAcaCHeAjn9oH5FG5k7xjyhCY
M7l6KeJ0V4uyzHyCKlaCmHwm6OyoohvgS3Fab8u4+0WCh3aQfI7AgLgDvm5+3SjC
yq+MFAeYeotCC7HsOBu+ZrDWDWJxUMwAb6mnb4rIo+Uk2B1xC1uM18ezhnk4Nhue
3ZtBOzlQvd19R2PJUoxSrRwYZlB7lWuY8sPlRijqSMrOXypo7CaIycOv7CtyPF1G
o2gJYt4Fmzwvw+iPzEVVm7JCPADsHqusto0zWVQSV7saJuUMcdPYUPQbMcajogbJ
VqoNQGqYHPvMoepM4Yih6i+Da3WmUeVhpnXB+2NM4nK4zF+tTIJ1GEI+pZQpe6ba
tOKlUMSzK115jf2OGi7qfg0kemVz5EFIKxX7P1j8QrY7LUMamOXPobm/RYMm8aQF
0boClcDnamD1N/CdoIRBgPgsD90y0DQQtgVDcVKwmIt7+d1NQ5Cwj6wAv+6xrB0L
Whv6mP7SCgAneOcu8gp+UtE0rqXD0iHORQ2kPVXKMvfwiICtBckYiFOeCaZ3BBVM
PwxGXS+bsF1WIyviX2D3ajVOvbP2M1ZWAIGBnSxHHFlh6+hYZbC4nvKYU0/2lsi7
I9XvnJNCMLzkI2ev8hHcgxP0hb07asrecG52Hrs8cJXZf6s//U9Lppb/M3+6mTjL
rXT8wqxGmciVbOHYjc/mfrNdmS/3dmrkDqoI6KmrEktb+IxutvoscCdQ8bC2kv0B
OxYOvIUXNABC1BYaIAWy3EMurjsSJASZ7F5JvXuZQhmIjsYQMR9kRGmcAyA3Hv+P
+b/aghkcX16uahPsJIow/7qPZEl7J/4+1shk9gcOCOunFUNxe0QEa65V81UTdflA
OIdFqa+dsAmTltl70pnUnO4BVgmkcgB21pMrfCwhZBgbtHP41+1KoEGhIt+4+Mpi
6M3IGElde2HPBJzWWL7qrXFymJQsG0kszq2CV6LDhnFoi0yuxaKjg9FTKDuVoe4k
ZiNeMKSHXz/X7i6JKXaqq1+ebZJ6z2+ts60fHm4q/rQvYN8Z0vFCWIcC+ALP3kPO
YqAX6BngATimFduhEWisd4YxEZ7wAar5PHrCyh6RztA7UQbI1zK86d9e0DFcOX+m
JLBIV0YaTaKoLw4tpW1hpP+zvDYWTkoonTfEQrD0jWckg3xDdUjUWoLD/vwlPW8+
tdabLQx7f6TAI0IYMT5cIcUL0cwwEtDfGTwcSUb69nTtWPpz+psUYmk6AMlC0Dj7
oNMF2rXnUbww+MpnVk8wL/z4+vBSNMvK0b3VnogZBU4DoJ2lWwd/YSM8nnHwT5oq
1GD9Jv8OL9TiEGWpkR41PaeaadTyJs5AYb2FYvHmPegAfYWU1MhwSSeA+9TRFfKf
w/FAl9IKy0lGMXbg2p25bUW1LqCeYS8FdUWsBRM21jsMoUkysNIBODItQxSPPM5R
LN3EgmYwUqwteOWmByHacWuf+KAQ4UPTgHUkHSGYZe8L76rt8ILdLRhZnwa8184y
JzQzffq+lz3KZtGPZyx9z6086SbrC/mJxMucKQbGDyb6nh7C834ANBVEdVlL6HCi
I4KL5149qIPv17hn/oIHKaxBdY6ZqZM/bhdLv3RDD5otTVx+ZmN7TpU3RJJqOLW8
Wtq42o07XBrYl3tK916O5G6JXndWbiWFnmcmZ98VLa52MClHaDCXKxbXBylbfEYA
8lb3q4YCqcvlTLkbXB0YiiWxa1pPMxq1GYXBnp4xQBmy7YQBKVHprPQX/0AYVYNs
r5VaSMijQ4qSl7+jxrSWlKh05IjX+gPryAiIe663aYvIjRAhchvv8queHdROso8r
v9T8RkyuRgrQIbFGie1eNLRld6ogWgBeCE2Ixv+tu38c5qWBmmO4TgaDkOYvWTGd
q+FbZt0wX/jQzOV0TdB73qODRVKsmB/dJz5uVyv55Gjjar7Qv+eJnANpxLNpy02u
O4t64PaWl6SN/qVyWqdAHdkhCkz5cffcs11UVLkBT1QcS9rror+A9sqNTlR5uUbC
wEJywxnd0tbAhnaz8H5vSqBrUeeHopn0dzxwGOQCOM31PEGjOEAeCSNXdHXup8jG
8GzCYEaxYLjnAgZrV9WMbSU9OPeBo2zTSCr6cjcoNg1j5EW2X6abDiRBxgPkBwsy
eP0ND4fQGJv5pEMgWrA2iR4gqyaRSORDquau3khw6/QeFwTt8duduk5Qv5LfMebq
yoWKKr60yYWwxkv+5kBsHF6PL5tho4IYKCARRI8rxGilAHOnPLG6o5h3U1Q7ixBY
uIgc6SX+ISw1hT0ueLjKrarcHyDgFDs5hc0xrX0PBmR/FJu5f4IogoLn/Vh3xXhm
0CJGMGMIOozukVqrhgsAGqvm/pVypdPmS1K3rcn8S+XXO/NMT5Lwvxc5xvGzNZho
joH2w2d1uz0XcY93Nfg1Vc4XJCvznLu6iuEzeSCbiV6ZIRNNO0yNq1IpHp0del0V
voKthWXNWHJM8t6fZ1TWpc32+6lUwxgiB0PgVCH/ADMch+efaZWHRsyb8vYQ0EBi
70gvSPpzhb9sA2Fd3R5Rj9VE6AgQBU/evVFOJFEFXM6II7WAUdQorx/pH/FBPA3Y
CrxKxud1zN6v1JX3O6XiwkmT/OQW+uv7V9tGqXvmAW4Ldo7VpfsdKnKy3bwYDnSE
7cb1jThoaFe5llsXCUOsuRd2g5x9Jnf4JS2b+ArQ9xOSLIJ0Y1BKoBvxq7CzKE3B
HONJKVwgMQ1wrbmnUdhJAFPwVjM7LF+n8SKIFI0fquRJ8B+T5L0GpEl+WpBI4z13
pGDfUwSY7E9NoXGOYgRDf4/A66FUI58uW9mjRv6Yy3leDkA37GESyzpt7Yw/Wa0g
vH1+G6cCM0DTWhDCqzySWQEqsdg4sgmOcMZVYMg1iTtNOVBLgovUAcH4CKbXWQHf
mEa9jG1T1m2JUfJXtmvcFcxQbwY3liEIxI5X5Sl5HcbCYf3bvb9eEXyWyAwvkI5t
Rpsj70SBY0C+2oJPSrdkmHx5F0Kc6IhN9Pysq4Gx69giFupMRLjuoSlYJuralD1B
dQeO6mlxG45T4+RKi+/uaXrwklBgO0zUCXhI93h2khN1RShcli0L6I4CHWRsZ963
JMFHn/Qw0vLdz8lik5y5G5eJnuxGxyd30Q5mpcFfAGOPJq9mLgGSeUz5F55gqbEy
DFjWeWg6kcKhL2ua0MbU2mEXyhHFe1p7sK3Q95CBFVPEV2lT4Z1iqJfqf6MxST/Y
Y1paaS/dZXKzv0ospE/bVhNhHMQVeMnChXEvNIxQB+b4ABjSmr62vWi58CLzkQlD
g8aViUwAf14sjEbQHCoBsQHiVUkGTZHxrGtZWNsXD9eeMuYKve7k50XQVTkIIS5d
JtKksgi/BUpOWRIQ1K4MyzYCYxygyOqW3oBqYFmkbgd6edtR92olq7xgtCT2tnmA
VApiN+Bs0Jc/tvX7AtpDXZCRFnlRadg5YsLQUTu1uPDWjtQxFtAlPl881e79++8X
WG6kjYoMktRgoBOSERvlxI7/tCMaRVf05pc39T/vybdEqafJw8DtXA12x9UgFv3s
tgeNaxkhInL0OHsc2kc8/ZcmIlFNauLCgCfamYpMEq213hPB8+08R/M/KUPBJV8M
kHBz/3Be13o43Qyiz5hFPUxTtZykMB093OnhxLC3QlxkiC7CE/+0pO2wLAp4w11l
e3v4P7qZG/PMdzYaPxkCOogOeJSz4gmX3S9Q1+0lANxvDuqxkkkijywaZh/gv9Ye
wU2sy+J7eRhWsp4rVuvH6MVoIbk114MQT1LA/zNJA22BEu/CjBvQ2LTuW02qZdvW
mwZJNCociqGy5msrlhN9DZ3gAXW+blfP5FdDHVxnaSpfGMnN6MwQqT7BzkkX1mOx
lt6GpGMPTxFpsqilEoV6Tdv9e/fcBW3YDjYzwK9CWMzP9QMGcF0zuOVjm95MbaMP
fwuJKtyaWkejhXKaIH3b/pbJz2ymvW1qTLen7uk6EXGxq6xaH84Myf0EM0kod8tN
UPqI7kCP9TugG2K36/e8E+8OAVNx8CNDPFtJYU86sIH1BFfFnqHhDwQmmT9PIcLx
TKk14kalPc2nmuGBfmCfkWeF3iylRwakenbkEqk3e8B17xdC0prznqAmv44O7ZGC
XhuHXfMuh8oKTnhKzhZ5s+zaRIU9sj2q7qLOvPOf/RjHU35NyJRUPaCWZ4NG46eT
v0gcIhKmYybWgIqMeUJWwl1Ulz+AQJyhKuhlpubfifSbFeY+LgkEPMk5DqFa8PLG
GfHOuSLGCYTjWfyEm9QJkNryGPJWdRN/SyxbryZ2smH3Ts2CYkXoxP+OM8a/KQkR
lzaUBk/G3w670oiouspUfJammBoMdJWdpQoFEPzCri1AMOqlKbflbZriSC1kpIaB
hwyLbksc9oBzcK85Bs1DQXIaE4lxO5uTLZ8bUCtRFF0ttPU8eQ+C2pVyeORatQYC
VKXEWpEqATCm6Ak9N4O2QH5LLB8YsEvuu95835br7oH+oBHCZ0cUjBNwtQuSw5wj
AWy5AjDbW8eQ68cRe4CT5wsRjIauZp8YVBPoQr6WC7zuJ1kfVT9j82qdpHyt7fYW
gIJiRKkuE8yjSrAOYMwC5FT3yqGZ5MUihSeAuqNUoDFRukFN3uHkwoWZaL8cirOh
57q8yk/43Wz0jUkuUOqEZkO46zMQZJ/Zp9pwcQeBAc0kIJdXQtB6Nokl17l38lRo
sxotygP1CANmBEa/Jvi4O862/7EBGSo/Cp6oQplv0HBo6R4N7zuABKZ+Q8IJ0/nI
o3MX1513pd9AVRIcMeVO0MCIJ1hFQ90gc8I+K9pjzO0/RZz+iVqKrNj+Byy9rBHd
OfUgxcWuzYfFhd+rHU8pFm+r1PYipl25+pfXbAQ19ceLczl7kbC4k/kblKS0xw9H
2ha82lcRlapO2iaWQnMpNNrAizLPbjkqnD9762TMSBsz7sq9umBdIZohw15kEc9a
USTw2B+60WUGxq8WxWQ8vDdJG/es2LWpABogz0+pGkzpg45595wDKDmxNwbFQL09
gSvVcL8LJd0jgKKPBEe+xVmUnehq/cBWMhTd6ts1TebwKFnqdYJQyNpQ9YQ0Kqd3
GkrZVS2yOj9HLSCospHyiBP/Ugi7w1Gz81UQ5ApZ1VzDtY1nqZP3fbigpYYXCxv/
PUO5YyqDtNo+ojTALQyutffL23jPd84gEZW4FoVPvzvZdTcrEFgUTblf3Z2B/h1K
qBXg3Qz2lcoP0E5jdQFQwYrb6iIW7Djj7sKvp0GKmfoVOEPazMKLLdmhtezPMXBF
slPX7S4TOzEd9lSi3WcXTrv47kk42ZbIDw7UGGFG2rgmozEbn6PlJ7q+Y5JWDuQw
qBinfSAj8Q1QJ7b1qfC+Nw2KWU4ZefHet94IoSual7Dtr9IGHhEv8dyeutzTPHlP
SWFWskuriAzzyJR7a2tJRGw3wodrUvakBtKFLSd/dlwDSSmsjZXgoaoPgfZAbSDB
5pNxpICQePjU5spl/3DLzb+fJVv8vO0FV6QxnQ6vmhiErWdfNmwhvsSjz+PpgG55
UdyqFHq9dXG2xf6NAHd6Fs1uzroiq6gyb7DHUwQWOu9aJ6yAd/zc+nHDcL0vEJZZ
lM8PnbZ3M24lfBjnii4bimStf5+td6oRMR85vJ1SCaUSAuWFKkly9CfPfY4aVB4t
Vi6qjw3GadMVtLTfKx0J99jFUbp80ayudemHcdr1D9WQUydvggFaTMnpHr2Q2CVH
JoSmWzNjk3A79YYtA+1Q7keoYtrQa2RDamBcuaj5FDfPXGAO/diygVeZK6oqdvMC
H0wU/rLdVYn6rmZAl/st6Wu64yco+Hs2euP7S1LikARxynHls+qhgFod4lw0anDj
MnNridqJVKkZb1/zAHLUAu3jr4xsS0Hp3F16HcoXgus0QEk3DxkHflcYojeqbYf8
b7V5CgUBhxWnhSV8SLkC87OiwTv0diexAo1G/YhSYrKluV03kvVVL94LrL6vGMb6
RQA0lmDVzVRm//sM4GuW48pgaAtbkNN9YhAH+OVLy10NEdrOrNgQJFcLm7rVfDZS
sY60jU2IsDSncaUTS5i2MilnuYz+UNLGkYSXMU3hLa3c1iMvpP0horBUUWbO1iIv
AZZoc9w+l/mLIXdYD/HZ5zXjp44cFpbOSBEIXK3jdisW3FvS3RkOqz/qa6SafAue
rFYlfp4F60oOqFTl4Pt0ODBP5eA21mpta5KqDSEq/x2rtcct+2Pkp/8f0O8eaDer
uK1yHbWZBShMtz0VoeAyYFtqkwirEPiaZsLOyMQWtvhhZHdxP1QSZmx9Ov2FtxMz
xWuRhDLNdWJRfcAyOFy7NzuAI/p2veFS3E0QGcxM0kUaEbUaq4jQ1LLhkPNSWXYm
6DOEzHGKC0NYDTPEtjtBCJkz+Hsyt7og84bymq6wzXD0nUqlrKvv41RiAQLtZZpR
pttEZ2hulsu0+WQ//nlGtk95GYCuUNJ2wNCLtMYFD3Bqn7vT+q4GSfjwHaTcv+YH
dXpfc6o2xLE4m1cZUPBIDwcAoI4KYWfQ03OQ9fW9GyA9KmERFAN6TqWHd0rhW8Zb
3OXOK8QD0O1LR6nHcBIcDaBVLxbb413PrSosa801OWsvfWpQU++F4GVdqlozkmBk
hwQd78lXqguBGZbRo5DQ8iVf4Hhcfy7UzLW8shQSE0XR+1Ira0eGTMJvpnA6+A4m
8oXe1k6mMbZa1ARNi0PIXHkEW2nD2/bmr5oIWua4D74H7W5PgAt/zvxDTQc54qza
/3LcyQYv9UQooE+nFdF5jIN+uRnPo9/tdSAzmf6XOgI4THwAD6nZS1RBcYcTq4Ay
HrOv/HX3hOnAfd0ILCvVdFU8QAHd91aMlyf+QR+l2O1uEw8ARXD8cRT39pe7vc9z
KHHnYlPc79xwQ5DCGdpnhyxV9siaOr5ojho3SIKeqYAciA7+4xP/84fsU0EjyPWA
DH87FqEP4SrylwDq3fTzrkdI9qR8gx2WCBKEGp7zO7sLk7P+AlqA5xgA3l6oADIi
09woU65c1pzVVblVYnZ7wdXEWU1IP+IQDhBQA4GM03WsgJmGgLOJN1/DIiGv46KO
WxE5OGhHpXf5UuiDnPjt8GpHq3EhIwtDMGsmb3lxUP30vCGZhOM7QhrDmoUz+NMv
2KvHbhE2fNeFoK4EzfdiYrE01LuAMxuYHQCOII4/I/zeLc4KzakcuM4tUUjIgHY7
9KVRc02KVWJKk0geofm+ELnVeaEaUxCSRiqOw+uSo8fyeKK0HsiyYujPvGhxzToK
jIlcRyvw3CN0XsX8Z4/Y4O2jhQJYDnnNcLyfFopoTACZDZjNPqQCOyyUNbTwomLl
AmV4UCIW4juKkS1h8DRnpuX4Uraq+kX3EUNtsHmATNb6lRCQNd5UQAApKart8WYG
fvBXvh7SdkPpVWqvwZEmKsKrmJ6mYfrC3LaTxiSwjeiyHoJJuyAiJgEqZc+21SHo
Iodo7UpH2y6EfdqZyRu+ZqQzmAcRdwo5I5JRB/IZwYyN1/eYzIbzzPuPnm/8XzPy
jSDLgK3MMp+MW+uC/RDay0LIjo0GZ33PiZQjodKDi4vJYkyAzHungfhAgvVso/cE
7aHBPUnMkgw5RZYFqYhjDc7DClosy1z0REcf2je84sr776aUWsFQqiJorPlz6V3X
vaKtKlk4uF/Yd8nPFPA8UiIsDtLovzAOduiPC20TA1cfIkF1HC7wcs9+Hfzoz5gf
d3lUZPcfPKycKNbTPy1KwiBXW1YZbvpE7cJKIUW5g6eXgGnKVhBzT7JPtQu6bS/v
HlUIcqZrdQnEMHbEGx7wJ3+BlhwFWqPn7nDpgwNteL9B8qD9xYWg60JSlLc+fhym
iBrIgdghtocX6SFy6KEc/XoOcXiwWzta4zCMhhQ6AMrBkhSeaZ06xKSDythwCrOt
u9bsW1iPJrI3Pd6spZ1SFwyXpcLyw21aW+NM9sQiHhf2WBtULy88UgL9ob7BvrPb
hAjJzFnqNB6/8g/LXTYU3EAOgSjMpj7y7o7DC0b2AhPqCCkfRctrv8GN9QjJAUR9
IBF6chLUhJjTSafXuC+2SNS010PWtHTxx3Y81fE/D3LrLTl4kz3qzUMrjWyABW6J
NlVNijuNTN4chjSLuEaQSda/enj3ew7LTZ0Q8NyIVzGmB3bGXBNmD1bcJWA/vqNz
QdgJR9vx9Znt06Df5871tRo5Jm73PFwMdhf6AYTKkVSNqzXY7S0rBJvNFEdqUD6l
SdozlWzbyR12yejhPr3SeF9bOt5+LMqT3PX+4AH8sAy9jD0qsQIGJMsxKANcvBdO
bs0q6nyxtX5qWxkF8v5oXgBzwL83IZHgi8r5//ShPlXKdtflG7nOxJPQeyu0oVIT
V35DERV6MfPlj4KAXVMd4hf3z6gLadLHBOdD2tZkfOjfE9P2HcMmsdEWsP0weIzk
BA/tVZmetDsCnzB86QpEMauEEFwfiF1ZK51soWhSxAlyY8Cy8O2jFM+fcS/ZEpV+
OPxK6TipmWT7NiA5FQWO+GdIxJt8ilQ/YC59exTAwG6E3PEMXzildwuuic/DtW+5
D/IvgD7ecQErRGVw2RybmWw0ZeKSyJi/ffglWvXUvHsSFyQglfWeqsAptErG5krR
r4j5z2YU2T8+JACigIFyV5ZEltCzP9io+/cqC3s1PkqE5x2y5Vvm4CBJvU9SmQuv
JNw20G8dxxc7NZwGJv+pXu6HnLl+Px8YZEpbLEgDCt0SGQT9nvkDzQjLBVEDLSxJ
VYfqwy4534Q+YEYOX5/EKScWoEMAtOV7FWrSbljoa8sq4WnTqzz0EzmNMQKhTMWG
Glg7JcVfVmaal4Re+8b5epRdF4EuHoxr/61//o2ixFmBKXsxI7DMBMOx4N6WX/w6
f2U6V4Y/QD0s2vOewvA7+chjNr3sHlTBicZZlUyeYND5ncd0fNihV/nPgVmWZRkb
VaaOeBW5iuYmmkeJgmoV5UB6mZhPfQYXQZQHMScGjGb9s3XrNboN6l9UATe+C5PJ
zxfAAn1MGGPKmgvKXPfvoqKNk5JGB3b8LznDmxX5tp4C/ZrG6d3ShB6JVLOq1FEA
hXmKARZ0pSJl8EzUQXIpo1t6uoEU/ixR9kvHP5NepYjjGvhmUViAyq1cDX9s8pHY
yNPRnb9aj0CxlweFJUQF+szr5+3MhCPdp0JPac2/mMbWnIEYhvAOfkLU2nBdHBdB
jDVkt5AKlDFtCn9lYb4iZqrHO2zOHXVQtFYuVnyIvX3PvykQxL6HLRn7G0g4tynr
NvNgvb7koUCAyAff+52bayiz/Bnt/IPxZVoHbaQoqiBN6AF81yvC9vO2RIwNLEKg
HevftyMVsC8Tiz8RNEvJwBP2YxnIwT4Nm/kz1CNkA6d6EDIa0C7R2oXN3s24uRSi
YAksrTPIXQo5pws04bDi18RtWClmArT2xHD7R7SNqCEHuA5E1UKBHOyVs0Nckqpb
c8SVhnK2EwJAbEj5xs2wNxdWLvw+ApZOzOSbDUR0bpD+A1VqJcO8i5Lu8VpAn7Hf
XTANJ1ozQpC8Zz5yY7G65S/usxCw7ePdqTWfgngJZz83PcbDbVzUUzogCHj2myti
7B32OTex/zTjDbZO2ltApJ/uMz4ZRCOa1BRKyum9j4H8i07fwlitcGo8fCT7OsPA
9axfDHezI4ICWIdiHo0k07GyDSsNjuieinSv0T/vW+nXPleVZGF8CAnb+BkB282Z
BifYp5qvm/H2GRS9oayuvBI59h94xu9W5SGMLBEtHJwEL6pmuyrTke3Mx+Ej8l6N
ip/sV5rleEouuBWMM76ofjZY8qXOBPf/N3prWEKqVPgoeaLQS+Q+xqrNYrLqO0MO
BJl8AyUppnKEtK9QsDwEP8pulXAzq4MrgAlkxQEPVhaCDyEnf3etSgWpgTKfT6ix
lBf7621YycKmz/U2C0TdskVoXrD+tukEU7tSRJ/6nJwmUyyY4TpkouAZfq3EU9Ai
O8lBivdJLFnmGjJrA4BnW8hB2ngFBntMpOCD+c1vgkkNnwYfq7BQstSixTAKoCPK
UqiUb3XI+EAwR1H2tSn8AQyDDCm0AiRQzJsSugnjvLDxiP3FIe8ALZdZHOFh1duJ
TUQwRwjgxa0eGs4ynzvtavI9w5z2R3vmY9HQ6f+9OeCU7ziFxiOcJeZej6ZSn1ku
s6fTtfUGgXe7vLnz6otQxUYV0/W80cXhlgi54Jy57z39awLvWbwQE5nitxw1cnLt
VE04ivPFIvbTaadLpnegbb3SOr3yfuw/BvyaL8vZ7RPnlUBjgc2WVdWvKLtYhIyS
n7wUThsqC2xvgKDpJUKD0wiULgx7ZpzQD9fBs/h8KSf5KDQtty9QZKqh2nCJoQoB
ehcf6Lc1JSRebrLAM/4O/DRUnDRluqV5TgqgzgrGm6rANgEvnC1/EZ3q49BeFdl1
oLb4ottr53N2L8jOBRjDTwzxfJxhodN8nnUwlSZEsZPs/METAjKK7sawzvFsEKin
3Qo+UDBA8fYm3/d7Uw9zf68Nvw7iyX3xj7B+jOWQYl6YUt6/5un5vg8oH7AWSTJk
1U54ND47Pz68BcmPpotP2cfdAjE7U9dyRc0+Q09RY4YCU4S7k9TBUEVdgQKW8Gut
ggNYjSiXyUW0PD4jOdFSL6gvDkxrekac7xmtJgiu8cLuyFa606A0zDLarbvldEOC
mGCxVywPaou53eCD0XSsRfKp4wupMUEf9T1IIbjsw8hM+9QycjhXIwM4i5zQY32x
laGpoV9pPUyh/2cpnItyqEOFzW06CgqYZn9FxoR+/PqpsTMhcd86mbggD0wdGvqk
KkePzPEk4bpjZLgN8lH5CCNMT5NES96YGz+7hAYsgzaonEb0HU74GOLucSu7G6pK
FUTm73bXutQOGOCuvzX3czAH8tKl3+idBrNYP9e6ebzmne+NhVsSCcrP7sIa5tu3
Y0vb537Xx0Ajxj6StLJeYnc2qCEA0SCrmHYAd6gi+Lwj0KcoNSGaGE/ZfuwCbPSZ
wyFEiZf77FeNC32/Nh7xg9FOgPj1Kxkv/tiRJcCRV7kApg6tA3qfZVt/h9ZMrIqV
94mqkoCaFVWdCwWySV+wszFzj/pMIwVqakRuSc7KD2OFnQ6tiQcP0zZJWyw4Ezlt
R2Udmpnqka9imKwoafwUUWbVYXtZi1l/kmHdF1/2gDabR54zDgP0yCZfT1wYusHB
lkWozBKxxUnys8WMApTKZUkyIrZcXvbxUE4x4yL09sr62z081mgg+rob1M8fFN6N
ZpHPNDQHC4guRXdQgENVjPyQ+YNmaeqG9mQpVMec5T146GUsFJyt/gKcvTPzZ6qf
9xRWp1ay5rVxVHxLEjbR7I8nO2VOH/AhP6aP2jEbLfKt29c8t+JvCkZYB6TifLDY
x5h1Q4jfGVA8mJEMoTun8vh5GQPcMD9mKNInO/kl9iQUvXgpEpJCYclGpcrm5cca
vxaAyB0VdmbaOi+mwUNgPTnhv60Nwypq2c0GHO7p2vTofos5WVC9jN+mKAUXvktA
svD5YRX9H/wBHEGO8KnzBvXhCCG/TKcukWLKrus8cj3QyOite+4TDBZ7eJaVNq5W
EAPLmhHz0PSoSLPJT5PgVxCNC4JwkHTB6dLo3vGLqyy7bb0DjzGgQrnFG19jnxwD
TugQe7kQ/WF4Pdm8k800TujvL63AvDLCrQdYFHsg5yLZcRX4t6MmQl0DUJVTtToT
Kd07C3JiuL2c77r+EgHzZBAk96vVssvaAolUEYX2xJk2To8jDGqwhPWqVJxqjJke
P3xg5wDbtdwCa6rn6P5cFm4TOh1CesK1mKYFXvBiedV+CIOYwYBm201xTTeTeT9c
gpeJ0RiQl3EGbNISrWgfVPrrj66Sl3C2XIBCS4J1Y+fD2BlQsIqFlTXpKgcJeIIz
RVXKq8JTLNZ0MtJaJOj4rK1Y0t6AuAZ4NNoncRANpFemE8AUPU6FXLTe76j8MPm3
Dw9vDfaHnlVCXfXoEBb9Frw5FhBymFjSniKlzTXW7cCHua6D9MRd23o5fznRy7Hw
vrahWP4IFmj/Dl1fJId2q+ySxbeSfEcQnP+cfYIK8qUzLdi8F0cqQ6GIwIbwA4M2
OkjUcMK17917T+3vBgASnvX86+GIsIC/x1L62FY+517/1RRoUJApsReC1i+Ye/an
UNYEQFtq8oHucU5uctpbV5g4Rgpky1lMaEaBdo31cClXQ5qens3OVzj6fy4HRvHf
UzN4LeTQYAMXMszUrxSPc7B9eb0GMKeyys+1uKnMCgXTW8kqUdX4hijDI21eVhZ/
0mZcdkoaevG4Ko7ex3WwjuyNWjbjxCoegy4NI0CaxPc9v2i4/9ZzauWL5aSC41OX
bCUOJreMo8q363J4DZzK6HIRRRl2uDFQJbhTBxB0LQ+Rn3enC3sBs1X35YEfZUU9
Q5IDmnGODOknCiNv4jKr5kh3HmjQjMytyy8rx61+W16ulJCT7bQyXTLeIYg2xuWm
9/+EQZVXCcKYpBbcGh67qde1oMTwPwbwQvT4+idwe+yJQ7skdxj1QrK/pa/EK5zp
XRrpLH3rgjlVsFnlYlBG2wUI3jKKSN9eOElBRDoJkUF7ES8ssTg630x5NKsMu/Hp
i3ctq6ovEAbNLAjZOtAr4x32dwnFDaaqFqLnHEE46cYyQ0OaAqga4u+0ep5Lgvk5
Dn3W17VFD3D5GzlU9upnxt23x97VQNfWdJfpUhguOnXxugY8twbCslU5k9HXqQsJ
o5kenGZEs0w0NfM5bJv0Rn734rPih9b+ftGXr0tFtamTdNuMkhzf9n4XjWB2l+7K
4D8mQcmZ2clOvkugQsE7ic9k2jUO7XhAC1oRcQfKy9UNwcnEEcIUrRgkBsuDoChB
yfCbo1sc6A7cLUvLqZ2kjT4lK5qAXKcuEuqYfjVkrJH0dECuQpa6i1iBg560bKTt
/0AehEAS/uUDg5qUBwFv96hmj2lkbwCidCFNRpCs/tlchDUBHAlKw54pduOTklie
aptqT1j3W/hiQLUWCLQJsaFIaHrGeK9GTeZ10aIwO1NC1cMnesyrxHfBD8MhsKne
aIvq/yVljDB47EyA9c+fQtiv2UDbxMRGq76oBIqQC5jPwuvBBAfD1RcQsqpIZzyJ
5n7oR5flqBdm/og8wu+WQMkfr1t5xoyEj4L3/9IqOY8XPEwCKkUNn3lTU7yATkka
ie7WQTj0l3XhaTxik8NwuJ/UfPxI6nXcYgIuiKh6okwCmnHSvUAnIdek04txPF+Y
Ake00EveXmA3ulR8LsGoD1/pzS0Ve9kXjyQYrZDdWtz2PRqoKcFma/2HShkEr7tz
FzIZIRyHfHX+xLTnvW972TFL5minvoa66BHkppiz+Au1fq2JsPKh6R+NkdSFoCKi
U3wrJteUEn3Appi8SMO67Ldr4Ju4PUBZ4oHzDLZt+82dUzY5hb4RI0J4Am460YI4
JiWiCJxGujzseHAYnl/pMTyAkAC6TWrshhQm3yiizTggicLt8g4uVK6ZwB6eh8vK
7j/NPZp+0IfR6YfoUgGOTbheoMTPxtsKyF6368+/RqIJrymherzrfUNim0J2v7d5
sMP5n5l/YOnzSDJ8nWvw5uiLPjAIQKSPmRpiqSgaQvp3/k5yRZjtz/LPorKMMhLU
GwJNQt26T5SE5WYF7fZqAPZz+gID3Ez0LHXjLEOdWukKtYIiMPMepQZNVmdy27Qb
vI5Cy6B/4hNUvJ7ICJKEADYKT7GOoj9pfsPGTL7ttvOdA0u2fP4siU+ykz2Q67k+
8R7/YjS5yXpI6KIadnuGRHbkoAXgmROioyRxoRMFH1odjCUiDCzzfMF6wMA1e2r+
mxsoWhDt9rS+UGuimUbSqalQW/PrpJQYIoHfwypKAMPA1XuPm4XruoA7SMQyApPx
tmKPn21i5YI0I43+q84AScXMYdhIlivr7jDeiYe7Z+6lIdEeh9b1T+qg2fHeFCcq
gvrGlPrNGwOTFXnfBai3UsMLi7w2HUuru/5J2dqVmOk0vVTSfz+9mqKyx/QLqGIB
JwH5jc7i3pV0sNWTAKXL7xIzgwA650CaZwzBBZgb4LBh1mjZ8mF+b0TNzqZGClZU
HZFg/fYpZlR6wE1dX6nKzhlRGdj72VarP8tcwuofd4+/gB3zJ4H66EReQuaJpz5n
ASPZepxsyGJ7aXLrH/nCEMvaV9t8b6oYLR0IXBsAItxCt+MLUDJnfLSV845Wk2Hw
3w/xHpfdVOvCY+HpGnnXaBltBsfXHhgfVvGAK22Iq8iEcPy6IbxWrIeS7LrHjsrU
OSelTuoVYpj+LVGAJnz06Hl/5Z8KhomSZMc1FD+9tXZz0kYRKL/Q0uCPYH1GbgHi
PVcvWmQ1RTK84G86j9OhD0R3y4qTEhJIFQrhtBfMOn3ksCrbHvswxFM3TAZSUFmi
ETXqdgangqKPB6Es2B4mv4RJXLe+35PCkIKiclxZb+ehytzpa2ij4AEy5+fgmoGA
57mFRJrM1Wd40/y5ZNiNA1qig9ojBPNl8wKDail+lOUzE0cqHozt390IQ6gBXF1M
MR4UolXSThLz8kXsiYypM1SE96HXE0RlxLdk/1N82H62MgvMg38LNojfhEBucnjS
xyX3Be5Bd6dBafJhyjQ/MynmkSY2x+Xl+NWD9g+269k7ml0iQD09qd0eeG9zIaN+
rsosVC96RIWg22Uwbax4lgI/GkTSpv6hqSjp+OzsqYHVi099J7860h8vSDXADvXn
6n5M5P+q3rVAUIZTEkSyuDYgIRMMZY9JTvJgusEb8s0JtC2vQeW0WQVBDy5n2Zty
iDifrA4kfOJOkQtIhQ3yplpIDDBLMQIXeKR/G7b6KisM2Cf/iPnBWAeOwC3xnUSr
p3/UjMqf/zU8mTOS4AC4CMDxwYcvF+driIh97xP4gykq4384rRSpXsKNUwO4oeoa
on+X5PVx+bTvqqxfc4dSjj9UuWA4TeC0tSyLA5vHncAvY6eZiB70dbeFxLeaGbMK
YXb8D3+GCN6EA7lf07M3l+pENfMDdDoHykx4doz/JW/NJ9qqRgbuNjKBEZ6kWNfI
bGmeWCHD10YhyCqCXe1G/LpIJh+sV1fhqLLKlmbfwVQv+h4drzs5MI3/wLYwVkGp
YZ6ZLEjWt6AvCXE6CCEjOisZUy3gJxecV9GYlTUBZ8UIK0LFyD+8Zu+jnRp05Qt4
D9q+jJUNsfaWlBIIcPWlXTblDobs5m4vmIdYSG7YAcyFjiTyGQEvWSGE3HT/eAzh
Tk2wAmhNqqIjahKRznwRPFekNAfDpgJW32P5X72VpK3i9PWWQzl6chNuEx4Kaenj
cB5H7pt3WKbjjbAAgfmyq34LmiXl6l0s7auVEcJbTqgqEm4I6tBcEKJo6ubHFr7F
c+vqBpDxB5SK+C63s4dB74CvXyWqtBJi0GFSMlwriJL/aLwnpRySs0WoEVvI+S/1
BzbexYlj14yhpH1zNdKc9yFwJcL3N0pAIYOo6pLsSZC80erpETMxb3fY6r0N1lT3
VsZKvJ+T6cm9YoJAk8rvjyo+8cIanZ0xZLw8YBECHTRyZG7vWeXB7ruKgTO3Ey0q
SaKEJPsoIa5nu9SRnavj3hUhJERfJBxQkp3sW9RY1Pm8QEMsO/x9PUKJKa0huXNn
23+Ma4y/h/xeycuBd6/4SGrs0kqRmL22/jAnTr81PThoUDPxWryG+Qc2UiRMYmcc
2oLZyJfcOBMVXFDqq6SfzRkhYL+fRxelrSWCSj+CLc40SpvTzPGIoF93g9/A7Itf
hnikDpQ9gG5TWfdW86BrRB8xe3/aBzq2UswR3lyxLBPRROmlyHHmvTFyiI6qQfCt
rsVZEIPc3hZlPOoDJxctMzOXHtW8XlBTjzpZ7gOYN1NHxL9Aq+5R+SCPzciudFKp
Tl7pDYa0iMleC523Fo0xt+lecFRRjT7+/Zbocw7+6HYpcaEW+X37nKPugTC9h4gv
mgK0k4+TJtGGae68edc8SHCXARlDtv7uX8LJ1+uZR0ZpbtTPdy7oDrpJvNhksrSF
UcRkaSaajkIi6cuzH8hvXXOzoGShDQkM8wyYQDPVTTzgxGmKiAci+YMw8M/ai1iP
2S2OAIFga2nzodI/lzYpnckpf+AeBhHanLuQgSpVSwBJH8BIO2LnXYnuByUtwPHs
npgIkgCjvpuRJh7u/o/nj3PC422eZhnpmw0cRaFRdPC7fNT/FPirjUiXEM9NQU3E
SKeRP+QDKP2TKbTl4GvMOvMbvUyFQe85nS9miQjC1FsvSYI6ekV90JQct3vuHPt7
Msl05TmYXxrTyJxLxbO/43/ORd8upnJOGFA9ZII2Sd6aQJXB5cZkAu6W0AdBScqT
rz7inqv2+xGAPDSo9ANnvayuFQvby2KLpQTCw1kx9UE0g8UihgzSWyJtLTg9y0DB
Y+HHyeRMvQl38mnR11vUSYH+jssaakRMkvGxoT6U2VI2PzKgy7Ae3GziNdOuUjuY
a+G8RoRr5eBlbnDegf8/ernnsrpBVs6E5JSiRd9DaG8wPb/vw2vOF3Ow3+YeICRe
tKrU9rHztk0jTe7mEWL/P0VscC4NIEPZHjmLWQ/BTVebMWnNn+XDfcO6c1KcaexM
7NHMvpSVpBIxOlEcq3uZoMS7LtxV3yr5TDQEyCS8vAsZ/FcV0iakaqFY8CqLQAOg
5qqG0VuDY+pDsW13oFQtGgf0n9kA9irEjXIZZIzbB4iHuKr7n3a1mz3zqJbtXVYx
pw6a1YCxVrOE5GU19FO/EXqjIHq1CUNTSOMLNhCbmXdtzZ4TbSwf1Qb9a2Dwlhr7
9ahb5D6QdO2ulacM6Gjcj5EIBakCWjotg1CmyONzjLiizQ6hxaFYSWkjPzpIUYds
I/JRTJp66AHi3L8cgr8HipswnPQ3M6yaNgQzICkWcv2NCdXC11UnCa63UnDDr08p
/nNCgL29hV99f6FAJqAVkCUYHALEQevS1jltShQwxXvW1RRbpmzZOhYJ6WS/ayHd
cYgPeIcZ1d4ztnwNX3HPSApBOUY+BgeJgbRI+Kxh0tE3blI2asLTFRWdNGRb7wC4
eMnUGTVFXzg0kd8QYxYyiLkcPm+cXj+E9R7Lf1LpmmA+sy1T4//F2m09cGh0p1O/
yCPbyoRwznlIH/XPGPjqEG3n4+LbhDXLNqlni5Edc1WBnNeEABWMmh7WiYlJHwmH
/+kJcv9Zg0UhvJtqNmSqm5frxE5KRYqHtGF+l8MPgHHl+5BPkpoOYmV2VA8cRXwQ
eODb7GniA0Lb4bJRBSEK/El3aIWq7QS+0II+Cjshki6/cnJA/sFZbE43dGj+IQG7
rngm1mpS2/rIFwiZGFrjR7x4Ub9oOIOLOr8tQbGm7Kux/ek6fK9dYuvsgi5dnI13
XbhdnwKc2k1scsC54jT2tpfmWOGYeYlFiO09COVL7u0747DIzKZIxUdCskOQUdmJ
J5137pcqV24q7815yXOXpNxNhQtawJK9KtDvmvgU2Xbvf4pcY/0jBKAuFjvagwYi
KG8DDr0fgz9VeGUo2YqeqGonHDClQzWI/7eA1JSn1VfYDbLhcvvAdF8392w8/HUI
OyN3c7gg7eXnTYErE+zpQn8zxlQeCoipf+2H72vQRn9pdazSmd8yvfzJ+xkKecaB
n6k/iFfQLxaRkWwUXspp3oi1xrx75s/84FikH8rFsj2m7xMwcUUtTzq6VGqplK8d
uFfbqLtJVHkBHK0iOy2dIaobY7iu1W9cxJwOxzn4dbUY/cbjk4E6MOhlq28iYB4d
kG0uYyABB2UL8Wdv5vgIFPYNZ3VKQxAbPeZXxJ43pG8zPsdGGRg5JwbX+wCbPfsY
y3Es9D8KvdhEQDZIESwjIn9fI5sinfb8v+Rveq6EGw4FDhr197pTngeb3eZijjJh
3knYrc7goJeC99j73LilDf1zmO4qoGGlacosg4+YLjbzSA2hBxPkrSgEH03zPcH7
dx2KkIW5bzV+vFvI7a/5G4Bmnh/9yO2/hCtEu6sWVkMgn8GJVWjMAi2IuLHEyjXZ
I7lAVnXl/5YG7Z9DVoAi/M8AN58PMjxh4fO0qvRuw2elvuRBEJB14ZLhIybNAlUx
0llHlrnjajMetLEkQcNL0784nitNgP4/7UpMD0vllu1dIuL+rytYGovvUAwEN2FF
Stq4RWaVUeNVEJ9HgMqRyrEIE3SRQU4RGIAVXi/Ops7ncz8I3axVNCUN8q/QyuQ+
4RMLULN13XOupU9aGtWrpmc0ahQfsKyOBqUoQol+hxhRuffS6JWCi6X5YB4rPD6W
+HU8Gh9GTWVpj1nOvkOyUR/L8F1HVGhMdCR3946y5iVHG+0Ty3skwZ5bs6RBXvqs
my5Kiu6j0k2zBkV4BQ2T7Qh73v2ouNhiUwmIrKOIMYJU/bYKaJNLjzdw7maoXXcQ
Vztu2+K4QPf5D2ugQo3oUNbPVmxxu9ooKSIWWAZxnKBOnvRhGxFm44TGa6E2Oun0
gn4FUIMznVn12A3Q/UMbwgIPiUYMASs94LCcTE6Q0IxmRQyYAoJQFCRzKHEvGP45
18ruPCF3iWMQiqJVhwYzBcbJAzD1GVwoNPVqwqZdoov2f7fHUr7rnfR4qAQ/67Or
SkEE1p0ocPQ5p+3Xtygl8zoQz3bMS6BgPnLe6KkiBkGnQXzTvJ39Mctq5hPVdBei
27ScRatcxv4QpLK1ndYSAL624VtMZIgU7QtA7xv627K6dapG28zCq2Xg1YYf39eM
ukjkgQ19hUMLqYJkrd1KHhhdCkn0dIeodZQQEN4WNSEJtY8PxeviHOLxy1vDTcx2
ZJfWzGApXKaqM+n29crmoEqD7LT+j3c0XOgMe4vqE8xQwK8SkzT9IbzaSqwIgc1X
1BQEG0YILxqqZVjlvV7EC9OECykCWTtsXEFYV+FVZLHPD5yrxaqoqkaH8b43nhOt
3vdgfQvLgbYFUb72y3oXzU2TBXP8s/+956YOo8GvxmqmFlwsfIXnwS0lVKF1BGYD
ADa/lxdQqk05RmN2jjNlGdUjDgPHQ9jH2ZZYER/mkQ75iE6RrXNUJ8fEMyocDl0U
5abzCOKmG4dTDCjbg7VmZ94yyd6LIMyLPkPoqeElv7mwek8nEAP3w4xEs91ukiOi
x1/m4/x2scK87Nd9+Sf+YADsnZR9nfmDFAz/uVaWaSo3foJFQuQEj0gDXW/OUOGr
5DFlDrgwV5+CR2pvJBWrV/JzzsdvDQO9tY7sVrbZILWqwGN4RUWVN26dEXKQ2lOy
PZByE5gco/HVY2tfIpsuuNjJ3M27j233jOnLBTmZsGT+pBI+d1KU6juazusKfGh9
97vtuqtLSJG6yEmiV+AoFpGe3CW0hbl8Iu3mZG5ic2hYcXMX/EtXdlc5IFqF31Cu
YzuuDvf6JJwVy3M1ndW1kvERj14UBk8J91vejjJHMFzrNfJSC4q8ImjtCNirQP4F
3v3NSmmhNM1qRBRkzADfOvmiYOBOPw2kdwPKZYxr12YwGIkAo1ajVStv1dnLgdTO
95RGuGmUWYa/+IEiBx7/FS9uZjliplHqRkjMbKBb663O1ioX9HGSUz1jaAOiDvt8
NA8WAi5zA3jCTnBwhy8g52iJrPRnDqvhhg/lk5UEsfbGQgfjI6mitQW4hJkf4qh0
VvolWT5yckO80wXB/Am68eTkCRUINBA9XL0NeT/mV2pwpvw61vip8TKapq8N9rlG
SOG2uG1Pbx/L8jPAI4CIuWe+OAXDFWJiXWtKE8KZZ7It8h1LHKKqr2twrOzKCKTk
DyOq92qxGNXPddvO8Q2xF3w3zHUhM51zAVWytgVMmM6A1tbgZCkz6fEv0NYM/mim
pdwzYFCY2imvpwQmZhZs6wj28InmOuDRsbMLtfVs8Yp7MgeFeAgIOL63fyweEb7a
tnqPZbrb74O5NQleSJozAUX8uZwNJv4pchA71122FbYk09vq9EXl/tUsZ2zeFjp2
Q9lxpwnL9W6+nml9nu0nceYiRtUCeJ6EFEFJ5hs9T9DZsh2MyCgOtDDALKN0jMLk
RH9jci6YWR+kIALrQLGOz1KuOiAEf9OPnOaQ3IkEaJ7iM8JWDbah+Wx3dXmuhGIl
jbDXXb18yhAgUTTvQXgBe+z6I2KSXYkkMsBP5rxUojb2Ogwv2fEKpk+QYUUDV39J
GwhEnX6AN4Ez71a1vJPCpb/aHIpInkEzfg2N0IOVRPA5CdfgPZz/5vFOU2Ldp/Fn
v0dhsD6orrKVoqn1xoa9b+AL5d8hfO31PuQGXuCUiofXswoWFDiDClV+BjaQbgE+
8S/AGTSz7NJgqk5djnLrwHo7Hu8k4ZGZL2oThsycI7tIAa4zqTYsepmgVqJaWWkJ
3SjHpfj6DnYafnWNdKbhG5p0HY6uyOm/VazpoTlzE+ONjhz0PFh4Ew09pkgbgDMb
M5oIn/6zuE7hbNodyR9lSGeFzY7iRq5dw2IHuVAIra6zUTlfKqTlcaq5eqWKM075
qq6FhQ0jpxMNp3D5RNVIxIE+v8e8ohphsCE5gu6bdH0hs9MixPm1ZhZ8CiILG9Pt
ehKT8l2SlbJ3hH7Wkh2bzxMCZnpOe1KQLMERX25Bwevb/caKratseqh9y75v2feK
bdH/FIFHf3eLzPX6AOISmRMIDqo57vxP1eS4Kl7kG4hpVQ6y2VrkXvyw901OIWIK
CYP4hf6exyDV3jC+gviyHjJF7K1U7dVn7bBkMBtypfc+K4UyR7NAhdQJTkGUNrxl
LkPuqFQKWs047Cbn98xWFE/TXuoyhHIM6P+mZ2JJrbACn2sThGV4i14FuH5FiFr+
z1s5oLQuVG2Vb9+/lNUlppbX4Ph0kQRIAzHTMjLnf8xQgtr7MSkpwqy6cenBbX3l
PMREKw3cpJucnDTXNQotxVsa3N1MXR0x+us0qYwEIK9sXgnFdQxKvuoAvMpcdOw6
diVEu+eFRlnMv2DX+yLssvlAfvqO7vvTZZNRF5RxXrUw0Vq/aC7bUDC93sSmi/T8
ZPksmK2LFbd/7v/9LCb9Ifg2yD40bM+3zvwk7NU6H1ts9pJeOuTvn9tYQvYKyWMy
Abt4PbCDiNKy6GG86WTmzYqnu+rY38kY99Z7vkZmHNvB0t3L7GhMnHs1aZpBCDL3
Qv7BEHSjqWmcRYaVYhDgPYeJtf0mrXDgyriuKNRLG9Op0mm/uwR7z9wcGRHFzgZj
rYk+AL+lbAc21LCkFXmi7qF5Ns/djKCOS4Pnwn5uV+WZOu2+L4txYtrwBhmnZMPD
lQXTB6HSuu1dGzmvHzfHIBgGOw62kH7jlGsBRx125BgsSnObxAyoI1oBjQkCMFoM
NLOj0knIDHKh6k6d5E9q9fhZ5CDcaBSKvC1uLLvbyky80T09jFDg4M5iE3MO0LvD
Zy2uSdt688XZhpspxRH4d7yL/+TzPOmTYYeevWkizw1mHlWy33aPvXaYigzuzJVC
MFixCDOBXOtSMJiFrc/4w6QwNxrtgIesbJRsqyrADjX52t5f3eggkjgosmVkzUPn
VtbYFkj1jghhChxjYhh2O0HJFX23t/kJVnDlPI1rMBWi+qxJPCo+dYMIquRui041
fek6wwjBQF88H8MIPbNrZkcbBvXTOv5zwBkSzw4KdKBR7R9ajYFe4on6Md68m9po
6MEfwnALO8pLrCf3AZHEwuxplPPkQk9ZKDfRvxH8njuGflfaTJMKdq8n+kvUFRaF
5iHRks8sBrvaBbK3PDZwidflWSCpYbsEuGOw+MXR/WLUkcDxOJ4PluWueB8oBZj2
im9egMZfkOXvmgFFVoCnKcNflqBTS7jOkdw308PPBjhsanSEngF4yShgOuqhZgq8
ZOHvgadWOLrvQo7Fem6DzGPgLLZ0e8eRmICrvU47KvSgVSpkz4+92eQ6LXI5V+CU
Np+QcS/cKNsVn+85zqbUK/xUXkqei5CG/wCKmjCxcrZOkueqilodXhzGPt2/j9RY
EcbD4nVjTQFpolEyauQMvJZSNMRhwJz/TnOBqHLxts6Wu7ji7si01uqfFpGR/fgx
GcgqMLDYu5h2Z8SRW8cFb2nd4ZiYHh5TjRFb+kdhQMbJhUZBcOd7s2LvefmNAJXh
MLKWMSRrzJcRlEmwq3Yd3IXUB4QoHcj+Wuo8xqqsgbMSB6zq6DFRmt7urQLFZxiV
vOK3o8/VETxjsEi0SFLhNjHJyHj/VQNjE9ZDBBMr+3nHKgVYmJwX7jRpyz4n8oDz
+TGDfIJN28m0Vsu3AugJ+icLzQEtMAs5Z5uN5UTb4pT0V2qi80IefjPbk9IrDlZ4
QwzMggqCmKTz3fK5efqFVDNE6HXsU1u3/vNKuoZvZDsgo3fuo8ufREafiIVhRKXc
LitTYiYABqTz0CIvYaOa9YrrARK2e7r+CX1Mzy0JUXvthThydG5fNn7V/JcG2+6n
2GzdVNHumNQSwtZ/7ZV2B91pXGpebIdz2n55WIfhM77XPCwalzQvwhOBb/i8+Ig1
crVph98s7amliT+4vyVxBpz5YpU6w6M9AzWr7AN9LMoxBaW6szrFstMk5f4+Jv6C
Jt/QIWPaFKDFBEM838sRjlMxDpkoPMkFzFXzbzSzqQedUjC397GXh1nEI/iZIULL
LPXcpMeOxkp59JHZsEgZdoHqdRwL6Nx6QkPLSpzo+1Jx+MEwozGvtFkSREdFX/57
dNN2eVi10vcma6lNZ5beJMdFlkEkm3WaadEshMCxECmGWKHzQcF8vcxXyenzLPmY
b5Bb8Y9OscOB49j5eUu/4o23++mUXqQUOIlsO6EPEYIswDL0aqYMJqQ0WPbU4NId
ICojDypsfupmTDkUBYL9cwWeGpBO1PHFZ1kI+aQ56a8hQt6TbDYDuL94Q7VT2HDB
aZJnVyfeV9zZxEVlQt7Jzbq/bL0UgB6xfP2PabPRaQzsBeB+VG4Z1vvpqyMtrRrZ
NdJmFSqQjeKyT/svNUvaXjOrlwkYYF9oFFuTCwbMgtny3IrzjU5jwaxjHdoQhAV7
kmMLTO5IcdvaEzGiUrvPn3BJmCveIOEcFBbscBNF9cB+TtzJE9FbOb3QDg9IesoU
Rc9Mtfbewm1N9PMwiubTU/147tzRBKf1h1KHdDr2mU7x/lDh2lY56AhXfMSrBGus
bRq+fbgWK3un6JtNkV3RaMtwsdre4ZiwGznOdoIiNmIbegeFvEOReeaZM4LQ6Ewc
HzrvztpYTiQdxBQQWYsK1P38WvOqkUFMW6svd/ZcOJBxG3gqsbQB6VGYZl/B74x+
8TxDcEBliywCQhw7zwVc7Cetl/CvE93lxekICUk/9q+xJmRmIBYvL8zxx0hI7S71
wlC9JRHYzhvyK/gdfud8UgqtTHCWWOh5F+sAkW+r+P2fzN0sr9degTbyji0Uyqe3
OJ0w2ODLz+kbdNCm94UfTEJ/PeExucvQT34YSmyE6W4tt+MbvbTu8L1qnV9AEYhe
FjBMePXZqM+5aa8xTYXcyc62QTlqloBQ12Mz13gDj3W54GIgd+IKN9p3B/62Z5DC
af82TgPkUv7O2qzOl/CjNir+wcRmxWS5dxlIXkELAYuE/Pf37cri8GcZ/XlrunEu
0r1Uf9/6tSkwlVqgtU6I+XlI1M524cjLnVrlgccUvJVtuqRGmERoutBC0c1LMlhm
yl4+9XL5P0do9zzz1L7dBvMZqpK4I8Dx6RG1uhokVIomimMjep06fKyb6dhjN0Y2
DZAbmqGm871bAynUyPvl1mccD3iVENcdNdP0t8mYHAj8gFl/uOb7BCUheaM4FbYq
43So2Zm7UdXCj7lDzfEin2P2MTuyn87YXKbfOBLgDkHy/tHf7GCJERtOHArXswcV
Pr7BzFHW4QZyOTGaa2LVLwZ2NMzxcyP2/9jtbf/hdTX1r5TDXApLdFV/ZvlACosk
JbuPORpaJOUZ78Ws/7pk+4Ud4dEer+wCkc+i4QAgYu9qP4DlVFPyd2sTdTQGoLtL
h4Be+EMPjis6TsoqZ1j2sUrjzkqrdn/UK9GCPKWU5qAPeIxvBx9WWcpSKC6nSR62
p6ifcLxQnuuCoqVXBNk1qDSwFQ0AKH6+wOasqlPIewijbW+3ILkJeUdqAqHhJBTG
tUtzLAWIZBOabKRz7b+HDvI9KL8lf1Yu1DX+DqrFVyZXI/Je8LGQ+OhN6AfR5IOh
CVXK9FuwozZs2m+9TJcB72YIHwXKd8YKg1gjJPu3pGD2FncivxWiI3p9X57rJzDp
wFpphcGFQ8Yg9JctZILphrxrUGE4n5l4pc+5UIMhQXU7N+zMR6Q+Xgzai+FXBaKY
5ZZtkvmtCMKtco16V24CKRulL9F3iU7Hip/+mVX8CZFuceR8CuZ2OyIP68rjuBfm
p0cOKvOhpTq6m+8CdyUwTRxJixQginEdSyi6TqM62mUewoob0HwllGSCKVeajUez
4miT/meKPTNjX1jvNnFNu4+pN/HneJsZYKgHCpxt4ZoIWz155VWjVCXX5Se4pGXY
I+sxtn7w+Ypn75tzAVi+1BUcH7y0YFbMkG0dAvko9dYxGJrcH60x2IYHRsRKmpGx
yQIvc6Zc0md/TMEEPm7rMo3fDX+ovijxeg5k0h+BO8mZDBt5ZQm8w8Lg0Q34/UIP
tomTFSjicWQOEPimzT0fnqM1cFqrt9AgiV/Sizyvj+JDKcnnX8HQnHmf3Vc5psfs
LHd9/yxFI6Opqb6vc/V8FCWJKMR1snZJMHqZ5TczhZ0+AjpRPUrztBKnfUB9HlV0
ztIwb4snIzgETjoxmwE/UY6rzCLhS3kRpMKr+Qehu3elBAqiPrpFBrvTab8W1jjX
sNG2Iunv37VdjCBkPmvydk9Tc8LpYuQKKp5KBzON+BvJz9l3kypef9o23bZEKWRZ
4Ewt7Vlh/ovJUdYKB0x8Dzgs1bCYMkOQSlqne4QdNWQq678o23arCxc7s9Gu/l1P
y2KRrC5Gvj0Y8J++tY87DIqjLC5XdDrTtRWx/5L1/AxFbQ15ptlffWmaxIaNkFZu
v7fdssqy7Dx6dnuiUgWEJHKFedNpCq625BexBwoH32qEUfI/HwDPyMbQl7m1XEL5
fOIZAOsJUAttrLkUENv8N50Z8ZReEfgbi7kv6Q7t+XvkkDbanJXo0XgCR0VmnTz/
K2X0pGoZtliZQxVc+STp6kCq8dlGgXYmcx07eyicDFLEkIqjLN5m+VeygblTEXtw
hS5E5CLSH8ggB/0p4N39GR9aHh7SDYOzJPGSIels+MIUjeSYPHSmHnmPya53U+d7
69BLmy3RkwCOj1RdtXaSW1xS7aTI4TdB9XRI1ode/lqpgb5bYsw9dYIs4zRgMtyi
A0hAQKlGZ36LD20WvoEe85ltC6DAzMQ/a1DUlyZTf0DGwi1DRW2jLU3i+FFqoVSp
zgvKDDraUNLLwBS1a44u7alJSAjdKImLkQubnguf9HV5+USMPT0MbhKVayjP+goS
Q10TKUBDbBuNiaoQpGBxYAj7kGZDl2G9/vMDRrWVs596fMmA++F8833BDdPXJ+Kz
qeSu8q7O4ForKcjI+j8nAS7mpd72IqtiWl/urKoQImw+8+CZc7AFe0Bw1cn2J7lU
NtUL2VxaJEdLOhkRO1lAbWPyacxQTsOM0CsCc1z8wdPC+t4dlrqnB+kiAZlV/jdh
+gZxsOFyZ6TeaDOIXCbJ8yBzv8uwxZFR/ngYtRVfzfvC2Dhj4pksWKsBbJzZ+Dp7
6KVNnbEkTsdUsnCOEpqm5jMC7X2reUbj9RgR/QH0lnKk/wfu4SCPPKydW+TRkE3J
NxfHyz2+oZD7zqGPvgE0l8VgG5g4dESVZ9Tqn1oPrVwzlwioLZEZY/h/3YnXcUxV
Db7ydbi90kUT/juQVspnBwpXxfzrx68d5Io2STmtjxYSrvnKcVrogdzJrL7qmo8K
VQGBwH2ujT3lPehutKR20w/4hFK13hyF5xQCo1iZvLw6S3IBe980nR7aUbe1WYki
uOVQC1Vy6bsWWMJcoCRPznK2LLj0DeQk6oAc38/YU32Kw3OjOHdNmpL18aaR8i8J
XD+7PVKdCGCnO69z2lGtoDhftOlI6mTOLq92nfMAE47XPpDA2G0n/ZIZ/BKVtyQB
mwXjJz6t6XIHEcr76vutQvfg3uRUsUY957tXV+7pjXHpv/4SgJFnjo873/lS4By9
xAQOE90dNORcYpcfOvR3JU3mO1linynPcu1TmBz7WMEnqX0KngQXAGvBHIBlRC80
PyuYv8Ww84Pl/uaYP5v0Mm6vBbpTI8d6JNkwyuO/pJh3edSZTI+GSt43Y5lpKTR3
PFr8L0RPADqPHYpW2WCyaUdOLMIcZGFAPsYxP8cyeRUnOcGY17Cc3b/fTdpGV5u/
8ZiAHgGp0RpsDbt2vISpFUCuPDP3IIgvFe1b/kggOka+qiPKPMIMd2iVU+6oH/kO
MEfH+zAX/0KqG2/zKicQmsPvlrYa/5WIvOkCuwfEEL7KTguX9C6CRXBX+9iUnb/Q
wCrIMiI35KBWVIXjC3+eyWx0xyIAunzDcbbrci0JBmMh69UsSifatO9JUX59vFnp
CD9bHrmiqmti4n5Bmd8/X1rvFVObjUYkfSxUTOXuBrOBl9VGvoKIvYgM/Jzcq0Bx
ejVUCVy3hUgGpIWVD8vNpv7NOlZde3953MWq2BcBpU2d9ZzIrWp34C3MTVR/0QzF
FPD6/1d51xqwKR3v7ijuH02JG7nvwhDyVocA0Hx6dQHS1vSMU50EcB0HsUiASu/X
zdPkxHfnArNjtkvv5+8TSGtEg93bO5Mn5VfcvBad6jcPXh4mMQugI/7dPLFA6DSX
LkdDZqaeV7s2mCIPY0VBFJ5tyU/ZsElzXVrXDmXOxMxAwiNntphjnoSX8giPNB5V
aiM+Y2SmZ30f//+d+rGaT3YCl7d5mKgI5c+9DPFCn2IvHWgbBXkIEShX6cMLimo6
GhFNkQpQdCZ9LVQSMwyCbEmPo8yKkmuzfuDG33kOjljr0e9w3EjYtMKqEMp4MHj1
AF+7Fjm+mikfLfx7izy/iSf1JY9Zm3Axgi+RJxRzprdI5YNX57ASUCsZPLSnn/00
X/1JDIuKz77nMvpHxXn6iO19JKGH7/7Qrt463z+YnoJVJAvcyJq0MGbKrCWlnfo2
OifEBOjBE5X/9ZxAQ6djdLC0XDwzcU1vSy62dXoE6j+z8IP0qvyy265xCfiTkwEd
oHDU6WWlG9RP4QFRjh1rtPACpvQEhNvDY0IV/CQj13zxE9mjZ0g+DQrVfb6AL0r9
RIs9JviPBDow7hanyea23S54cWMf1c3GTCpvZh+LtTkRLC2AQ3x30g17gIuMsLMN
KJmMipdta8Kpuxy+Ldq03ztzBtFd3umABEisqrUXrWbjEkUJ8KpX3poCBnJZM9pl
2xZidPxolhq1ou1Q/FjH33LBn8yLlpM3oDCe2D+TWz+uGKVdKt/9Izh5YAda2Bcw
iwiseelA66bQ7i0cqlTYvoOqCV2JDDSWV1+APtrAZbBtTIyw84fV7gIqvWC/xHv0
ozU+Y0/XcAS2J/3+GRvKC86sUBjayAmKvkeEjkJk/maDGo6vQkXMufrDugWN+YVh
7WOYHJAP/oLszM0uww68z4rHHR1RNIQdxxqnMxGOxHYvOWkichA5vzPyqIWSDRC5
orUhrMoSa7+FzzOFA/ELltFKeYWNzp3WxancgrD4La5lGOmA9FYdZOYQ8TZp3/Dl
YY5jS5CfcHgN3/aRzJqfS9TnRU1QaERRk72qNaN4+P4LLwlH5uptzmMweVAfxoH9
meSONu1iQoi3e4cmvSVPsQ25LPVx6ux4/g3mRfhhtbg20+LS0ONN7T7auiKDW6sf
F4I0TyjUECXjkEsF6lb7nGUgJbl8GtUq6wprizyaWB8KEpgxM/7FFEAfQU86tQkA
hm5kHaO5oA9oKTZbVHX7xc82Tf7kmow0xetm6LmoRMIl20TEZ5brSIU6DilpK/Sv
ayPrujraGKmgBNRecNoXCLyTdSPzTwmEA80E1ZbZZ8uJCIa2icBgWma5/strtEAZ
kn8Nm0pd9PAtgoNlW9eyTKlwr/26lx49HJJr981skVYrH9U8eMC8e2Hf/7z39n9q
+AU+NhVd988q5aX6XEm+aGn+3lWsqcboKcUzY2TsGggNlZY1NdIWUTg1p0pCCBBA
i4wn72t3tOwf8YMyOLZgp5tNy7utay0dRAMWeFeg4VpcBrAlGmmd6TyK0TSAaC/6
RCkthrZ2gkQW2EllK5SWdfvq/9Exqrm5jtFH4NlXiHxBsEIN3qfe+4yHmx8BPWUe
BeDnUZN/J8NmOj8BU1JIXrcpHctkv0rG2IA0lYq0Hk3stm9HJEu6k0S5J55AtC0+
Gj5f7iWMGk/HtVKxset+JJhd9inUnUK1sQttuQnqKNovqVxkbXsp+DZQsJ2cuoyW
GMgl+rS2gJtCUJmSVfbkZD8UsCYynQdhorkAVJm49dwHvOFos1ZMkSmNunfwZ8Ri
OcmYRCOX9wN/9WZ4zHkKR3nRP3/Pbs+Q5M+8OJoVLpb2IXtvepsJvlYQ81dYpDPE
EYEOuoBsKLXxRHt2rw8To3JpqFmgaI28XdDYwipvjaysKjYwauYYoE7ZGFfKq4Iy
O+Rcub3PmnZFnPAGFqGhiFEUGTpgrs4+JQrJut1XYVNwjRJw3aTv6t4p1FZh8jsb
BnlYNKpbQzco1VDjH2sCVarEsh1arx9k0CuAyOreOnnHewJCDqpCP3sW0GyI5ncC
Gr4yl0SQTZZ6PMud5aTuHPfvJwf43BXns/0z7fe8n/bHoxKzKHfGRTgDwgYGE25i
azh9Jq6gjJnMAidEZrdpPbn0IzBmvpubmGMJuWkD9byalu9XBjYz3fV66rB+LPL3
BG+38Vnu1SF6giDH2ZOUo2qQL68ffpEe0VtYBlVWBVD+hQic7JGUcPE9GxjvaKya
BcVgnHL5nFn7FUAy6/ObkoEVDzLoxWd6/T6nyEdHuxhAdPIczGVunKrTONcvSjq6
gTET2Vtb4rBxdQVMuQWttHES8kCcfNsA8ZUvgl8DfLLkaC7lBkOxHdMPNOgQqC4Y
Hh0iVuNE/hPuMaQI0avc73pPg6pyjCCa4Vk+EoBjMljyhvNPy9fUW7Jj2w0/ptXq
ZKzrdFNxuDVniDc8ZJ4M82SQW1LiFqtUYFpgH2BK0dBkKE2PjKu37WR3PDehzBh4
YAesbub90g5UeX87UKWhiGzn6Q32GRJXXINxIWEWSJRN3XOEPXaWmI1XgaZwnTm+
ALpwDiY1ope1YpDdiA7KNVBli+eHU5HhpQ2Vk9MCOfCCjAZ4HH5EBk0BB20EXWQY
PNGulBQECcKrcB8Zw1oUqcYS1vKhOTineusajtpXQkA24uNo6/WhZzeEVXPVB/NF
OsP9rojdVfMAg+4Ls41v05N3azMiZppt62QOBNwE4W7zYQvApJHL9OhZWjfhKDfH
X7TJf+sgX3JvURgdLUVS3X6E66cx40THRXeZB5y/bxkCkIvWQ0lCpeXiY68etcdB
FFN9WntDuoj7KOmOH9vLwEfW/YYl+Z75PKHUqym3pSopw4DSBsVWlXuYwcleXhJr
qI4y94KVu9b50iCzUW8tuyXfatpV0mLlegF0BDYpOnlVCKP7NZXrmza9x8lXMzBi
vD2CAGRPGFyBT/B80ICK0Zbc44xJ484ssNLKiIrZmvKeXIwQEPZowpFbvk3XKsyo
u6FXh2EBYK6h3w9+Xgr3GRj+i5o5abaSuO7bp0bCmx541XARZR1Ptm0J+gwjvlZC
XnXfFGW3Pf5nWwXscsKfTYIhMcm4j8mrmEms62R/Jv5SiTC4Wz1ibXkop5vkSgtS
pOuW6Fnq3G4QaWegaFLWnhilDtQr9+MbUnsfmA4nB5bDMTGt8SNqoHlx05wGRF1d
obR7X10E9JP9SnIgyXNG7bmNVbrMops2nrN6kAyH9AV/8EWFWSZcMMYEYFUNBvZj
rUEiD6t7Zw8q99023XJM83h9Lxh/ZCPeTqpUGDsnnkhBrQVeIHcPsyKkNY2gA5Jq
RF0hMS18zAvn6b4b1vecGmyp4XEBf+UXRu9VwL8NXXEGFjgbvBJVjlo6Mlamu5m7
DXmjKOltAGKiruurE8Aen1PxZL7oi9JESDqCqJyhveJyoH3DsD/tv66R3rjsA5TX
zlDiRsba0oUh7t1T0xVpOhC8TVmEFG3JHzdZmRmJ+GnLyamkzKdz+iV5B2OjbtXl
8gwFBFjzWrlwJNmXRDZpU6Vv5rR5qRSkxuqqU0IjibzxSAzxRC287/sZNtvGkLVB
jomnuo+Fx7BDG4Jf6APHaP1U4uBDtLkDO7VboBDPIk+gsp8hDLT78J6w4Nsaegt/
eVTOLaNdQYixp2c48FisarTTAeVpMviYx9es2MLGTSJIRwXjZ4uq7hVaSIhWXxJd
VLJ8TZFPubc5jCRZWeJNVzDIrWGCZ1sg6I9TvOYYDSU=
`protect END_PROTECTED
