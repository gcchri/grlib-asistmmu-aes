`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ozal+bVGNLrc8GwQE0auZ3d2UySMW6AqKO0VMpdZO8Y0jtvynul3dADGIboYAdTf
dlpf0eShBK9Xw8WRN+Q9PbyRAEBCoYvvbJ2TYMhgNXrMJeR4k4sX5xpkzPjth4rz
xYiCWUFzPRjXQCTb2sa6lVZSl2zNvGgWDfUX6g63AvuyUIJF0GdtBJ/AqkkAdOkw
iHJd6zTJCmfdrxjdkBMZeSPEULvHW+qD0qRcw9/1pnsXhH5JOhwfutdVlBgkCuJs
91mEgODqY5s/pvJGrfMCOzz1snprmycnO9uRwciXWjVx7K3uTbZuVH57z5uoN/yd
3V66vK+/GOYqef7rvE3tmdsTVe5Zs+gde/Gg8bjz8fVr5dyy5EF0EmjdzsWAHTL9
JFH6Koppo24dR0oouHumrIpg5uhyXr7NIlOvma4QXScM1cxP9Z01vqqOwvqiFffu
qOPN3nIYJ5glF60aZEdXLIGcHR7W8VEdMWIqd6b2B4s=
`protect END_PROTECTED
