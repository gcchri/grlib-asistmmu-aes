`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
um5MkbOXI4VtPzwUOQu3pMQWGnaQW25hM+B74WEXkoVCQWjndzHjzreO4U8AJpct
so1Fj1rLuDEh7LAyyjJQDXps4I8Mi3Y0l+ljHp0ZWEMvFtCPVTdNZwqvzuxIJQLp
mJ9PY0NJwy5uKpSTow7EpFIIBw/LxWXoU5HdJvSskepOXGTDAcPdt8qqIP9rhF4E
KDOKVxr1wwlmxKCEaaVBeOE2vMgkPemerxRGcaa81PxFVIhUQuinGGSp3F0YsUXr
BEtcH+wYJ7oz8zjlKeQ3yQpWe/fHZ+npfDRlJS0dvTDUjmuEuuzZWHG5NCpdnyfU
GvD3x5UPsJ11ORc3BSPbvlua2wNmCLDu1AmgoNkAWCVOjEsPLTLPSAJEOTNB1Jgg
w8zgy2FirRUXILgNcRz/k96/rGNQhhLooKC/wYzvWmLrmSSiJ935broJ7IDhJvov
EkNnYyyTfOWoQFbtjOJlgFF1txyE0APriECUJH32PO4crxihkWxjvZJHm/h0r+Eh
4LqE49ianqf7wzM3TtIC+84T3xZKsC3cbrqFEz4J/Fv8zfK76QknzU0/hWcF+jt9
oUd8HfQV+9HWUSHVudoz4U79Ge33odYPUCz7masYeNzDQtwCjXoaKj3vYESJVaqb
kxmpXcQwvY3jzYH3OR5gFiWfCs6WlpZQAdTr/+Fu4hyOsKtXBMgy7l4kPFdzYJ6l
n+1uJ0hridle6HdYTPQhb0R9ghHFr/zFR5fUJfrklls=
`protect END_PROTECTED
