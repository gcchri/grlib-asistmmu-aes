`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xt/vJ0TYB/RaGRJE8RTd35NFg45JCaBGCmwxeoSYXf3gD1r7lONFCB1zXRzIdPIq
U8TPPi9ekDfmEiEHsa5ii9OphSjTAn9qssfLiPzexRgMjRfshQ6RA8eYEG2zMwFu
PVqMNN/pooU90ZYUmDizpu5p1csZ0UoX0M5F+pIUgCTlxtoQ1Kla90FGKN1+CmK1
T3SjQHo8ZC/GSKid7yvUBLMLb6SvCUgcXgqQnvHvP7xw2SwAmJvZsVoPFoimR/I0
YmypoSj94798T8AvvakdR1Hcfhgck4TNxAb1Qn5baHtFFBMRyg9exxoNojgv6Mku
RqMmogj3XqXJlMRXL158x/embfzTC476BPRZoTBn/BYI34F/codGol1VTsaT1MtA
FcIGRAhnYy5CA4vxep4+XAHEgAo3Qi1OTa8vcal9u2nw6hf/H/xvk20Dg2Pndu9s
ucHIyUeVfLECDgdEG9K4hQ==
`protect END_PROTECTED
