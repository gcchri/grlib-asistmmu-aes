`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0lqRSWyJa/ptcDtfS45ctcE2ZDoKsGzlBGW8WUk5RtgzqFpMe8n9fqu6sbV1wQUL
5c+O2oVINFnRzzeznBAl/muikWa3QwX3MX04ffbDP3lsttrUcx+9MrdVy5igRiE6
r9vPOWNBhf+6xmPnGlQCpPx4an5oDzi9Cdpa8qL0NX5y+dH5PlGLRKvrQ4pcWr0m
gTjE2Lj5I19agrax8ak1ii/tWHhkFib9HMgL2P1MdsYc8W+PA9UuUFr7JK7wqOWN
ZkqgSPQsaZdLA5Rd+r3oXQ108LNpMToc6Qww6JQhSCc5OUqAPb7s+ta2OZTgFm8u
nVVcWxliH2KxiQyr/oYkopOpVX7eZPaSw+QiHaGv3/XwWegwFfnycr+tGFqMvV7V
sfhnY+1WVzOBESciP0RDW0m89yvATw3nILEM5z99oVuJbAjZkEJrgeHUZXUl72YD
`protect END_PROTECTED
