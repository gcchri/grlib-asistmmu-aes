`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YGOyyEBBa9LSlOCaZbBB+yjwdswN6fzAucPpGG4K0JdQJUvWNpvhNo97hEyU7/+D
yZR6s9HZtbVhU0wC92ueYC+rkQ+e8sysrfuRwW6dzSxp9YaIJYlSM9q7yCU6wJhp
WfaGNw6H8l1WloPxUSaB00qPfE5mXBCpHkf3yz0IY4gVJkzh1SzotnTbUjYyfYXG
M4GmX2mu9a/Yd7ItUm5o3BMRkrv2toXqPPWja6UmGm8Gw/PdT1DKyw4Ku1+CmLnP
eC5oJ2K/yAUwIsbB6OK4wvzol8cNKcp8fX0XQmsTPm7uA/u6o4tlDrWTIOxbDien
X3auLAvFLVSuaGagPd7y7yYjXW/h4HBMOv5x/AhmFMxC8OktjSQ4rs4JeMYe9Rkl
onAZITC0w2NmaB72uizcs7shfP80McZgwr0w2A0QbeoDQ4//9aZVkOqDfqbSuwS/
K4IYKo/PpBfKLnTIHdERykRRkSpGfVit4r9UV9836CdicE/6EtEG9Q0x/7nvTy4G
UaR/6tjtVZMlOHExQLGf47/mbRooNVz5EXAzXY5zn63KHYlUje2EE6wL3J+kZE1X
M7SQTgK8f1BYdeW5QbHip1vXYQaYzhXAkYgislychc/iXjdLFx3HPavC61QQsnFb
Hm+1fw1sH0zS3WHiefbCmw7SUffztJR1aICErp2YJ1OsigVdu2Z2WoJw91FIz1vE
sG9nMzyRtPUbUFo5+ddhDXV9FdZPSoZnbzkWDb9WlE3FoO0XLhG6syIABsalcxEb
Ws9J7VhhEGT83Y0L9DRkTItrhgHYCnGKOcb7s6+fgSU/khjCD/x2bFkppvQovACX
yvQSkV1KSx170Y49DTvAjbakoUy5CxUIULvj7Ss0lR8=
`protect END_PROTECTED
