`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1f+XmzDhuXGnv5W778hUaa8OwS7yjqAsNt9M6ojAUGxZ+tqikmWVHenXVIVjz76t
KsmoE3Pc7Tqolt5LmhRBEM5N2Ffgh5sPeKtbZw/yKRAo8GbmimjvuNpVaQh5e5MC
K/Ltv5tjVqBme3o7o9q/+9zOEY5mdi3uG2AncJB7jGxW97rsKqqU+W1HG3ElFBw5
nWzl4oWzXII8KqdZkBR1zE95lITjA+M7OnGXDWE4qKRiqGVeb1eCTPaes5gTI5l7
cLt4ipPLvd0WEwD1arDJ8yemqBJ+TD3mJQmeTlaSjit/4n/lFZhGkhTIrMYRp4Mt
xIYAdYPzEkxwxqpbbNdg6CQX1CZfOliiTAOZA86djpMT4MMyWmPb2KbKXTxTKC7M
7v02X+AhQU/oIAEvYtrMZ4khhHVCXm2bAkLpB8xUM+rO89PFUuzJn28JOcEOZBu/
+E8cC220XDgSYJVDkVK5tw==
`protect END_PROTECTED
