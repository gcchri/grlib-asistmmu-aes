`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3rlZebl7XUar0dxMQsMLvfJjGVsOmyDnyhzODpfIkt12ZeJKB+5G3b8rcoo3YqcY
NTE7QpYZMwLxVJQFW4qBa88OETV+aL/YfhEHPOXZRcyv/l4sSdyME7LxAKeTg1Z+
Oh0s4Tf8eZuqBQN03mrv8WELArugv+FBowfbYymOoQX4QtrOPbZlynEAElq4HYOT
V0z32ZeSH1+SiECZqg3ESkz4RXi0aNvg1rHSFt7hkiG2jVkOLbj5lXEoGPPA8cra
jbeA/SeHljtWpZNbRXePiRcQ7OXj96I9bvfdLd1voKVrH3tPYb8EVcAdbcUO0SH2
28rc/mSp1PUSSENvlz2oIuYkzhhYvZ+GT246HwLEy6++dEqR4IXApfPutgr10uHS
sithLv7dALGEObV0MTHiWxvUAhaQ0Za3WuXw8i6RYu8HaRtKc6XiPY7syXF6zaiu
`protect END_PROTECTED
