`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ISTNjMiQ2jvAv8VQeFq4zjZb5ec3lE3VbHT/weC/QBVsilDFUr6SvwIPWfKY8joK
wXq60s07I2Gli//PDNOI/GoRQBLr+TcpbGuoZEw0yNNW6eg3DoebRUdVWqcOvKFe
LqgmMs0homWpDDxS1z1hvKJ65D0wooKs5pOlxkRa7AcEwgU5YsR8FmWSpHNp8yTE
SaSvruI0Mq0X/z58Ij1x0yWc1FnlsPNX3/Jwm2fqdCPmmjoWA4BRVgygPFbLVHLy
zaOWwwbfnAJKWcd9kLbqbF6qSOoqa09aADTSvYPO2u6VckX3l8wtzRJFQyywiweq
IK9m/jLiflSy5VXHve8i25d2QEmgyZnj8heFC3Kt30S52Cv7W9MsRswjO7DWLAOn
FQHWWkNSk0gM0yzglLkSJFnzvyZ/4vrMA453dJv6Sgc+PgYolABh5SHQ+Zlf88ge
WIgoMTdIXx+qP2jqEdtEi5RkflG6F+pPufiyvHaYfTe8nNVP/ThHIYXs6fBSgycf
`protect END_PROTECTED
