`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8JebTxJRVnbnwJ+rSMnsyUH3tdRtUpNCFlqOYXNTPqeijvM15zjW2t9jk/JWXUDd
cni8PiwsEcHziiRFxnLQbT/a37VOfYXNHQOMXZ4WTPOVTjEAwzbD+XDLUEbacoxj
VzvH4X3GGP9y3geOcctUlGl8G4qSHP2+rFnkvGOkxpUIPHglPpB/m81ungvSwOYL
hjr1eR0N+dhHmVnpOTk3s/ljSX/1OfkSvu000j9w3luQprwE5HHCtjzU10PvIxng
b3X2MGmPs4rIB2bxkXY+cpW+LUqvfo6OXON9x6Npp3eAk2FXJ1K0M7UtbCb+56zd
qv/73Um6sJut3gkWRlZqLQ==
`protect END_PROTECTED
