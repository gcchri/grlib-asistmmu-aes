`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ncdNDd1eS1UcIJiCDoJUtCRnIsR5121yiQgHuMXHygf64XPtM8BCATgsIcWLZafv
ft+83DVJbjuzO8iCc5YNG9TIWyIW45Ree3oWxGPxZ/B3+H/Lj7cdXLYxcHzO+f2T
kMsk5g79k32Co94i8UFCQCOy1EffDzsss8cm0bS1tDTOfsXLE3JGRwa3Ej+W+w/D
hypjV3z3FuG2gNq0S6xAcEt0M03oSjq1peJsaOHi9sf5gF7SVHeZB0hiCL6mawQn
wz8O5oKq6GecxX9gp94KQoYfs593c+B8ToBE/4vWt+5cC0yxI5vffn3gCvH5+dJS
D9WSCEowLA3XVDCv9PvXm29uTHvWheZXPmfLHMlUmaJt2yALT91aSWq54K7WJ9rv
X57JpbA90rDovfYOjbGdBE0fJYYhHGYeRiMH+1HKxi1zUQju3IM3WjT73Ei5DXdD
sH5DlHFHnrQKh2dX8XLjqQgh5OhNM15Jyge5crXtS23u0LI2yKunNdnpGlZBmE1J
HE+MS+AdHUED9c88JItAS++ZI6inDnFg0eR/ch0JyIYQnI9CwQ5h3b9UJi8XiP2/
7URYqMjfg2Ag5XAb75QqnH84I+OcWjrkvG90CQ9EGIU/WS/gBVjTEguUM9BjMgkE
tbF18Y8ymcsDWn6hrZZMH62pG+GmdnmrwlYzT7Xe4olqSrl9+4LfMZAATY0TYG5f
F51dtg6XUG8DVP5u5CnkrB50TZR+PJ1/dW75RsM7aun8jGq4/X1gIQDPGU0wIAZq
ZYSIEg8dWpE68dPMVoqZpX8KQofNGR0+E2fG+sDFwsvYsjmlzW5stNxiLWvEnDeY
TOItXw+mNqQuQiG27HPzGxcJOIUOyWKWCxRliuw1lruUCEUCY9QEk8QV5najIL4/
ld3mwlfaMaSBVkYyULZbTMPj4udCdMcZaJt22il9+6O3Zvhq/q4NJXVrmagHfyXW
qMqySkAtrLxCCu4T4NNVvK5LkqR2tuXjuf8qs6y4NGONhF8iuo8qtrjmoKQZQtiz
F+54BiSve2qITTRJG4Jzg0DlG7vSvbv2O4W/qPo+XAz85/S5uynPQC3D/1Y/OsqA
1XgYz727ad2uaSqZSQ4OUGX7dLEAge3wlsi6OqyhYfjIsMtiBJ8Q23F7dPLJiem0
EGmBzsq4Ba1t5zGA79VHxFR02q9n+VQbpihhP1NbPYGZlJkFyQrfwYH+uM1HGPBL
un3FWAS0vfU6D8iN60TOEbzm9wFaR8fCqx5i47Atqt0Y0Ianv1OamfVWUIsd7aL7
TOTYkXey7SrQ29HDG8k9LMLxDGwDuOooC2yn3VPhid5Isdiv0/B8iOVyfsqTAWUF
vcT8FcGaO2EyCqMOUiWoupXeByf4AfLzvQS6dqaJUbR8vDURNb345gJbXRwlFKEk
`protect END_PROTECTED
