`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HAEEA1GPr3jezjrh5CLXZQGWeLZvLEaTvxO5ExeWJnWjhPrM0XmRNfeU4myhHiF4
BeHtJCYD46Af3D/o9tvtqUzHXNm2SP+lnChx/03qrZptYV54AeS4iV6Yfe26Wgo5
AE5podcaMap9dYP2rfKUjWAjSVUhJhE4/leZ6L7S8NU+K87jLCQwiiKIfFpVymwJ
OAEsJUPTguOfSIx365jIlTOAWugyvCYBndlFLWYZgHtPyZ6t9xqgNlUSqyLS8BQ3
kKkwOYMeHoEp4hcvUUADeXSuZ2axQ9yxOkQihbwy8svRbqZBPizijYfxYT0N5xk3
lc+f+k+UpbL9/b+0uvqYJAOuOXX6zG3QaQccEuxIqGAO1iFApbN/FE9WrcdjDUyo
3vdvtRzdWv7N++6Z2los6GMiabsK26yzXUVtbkDEwvVlbAFFdTk2jY6IP6kwr5sD
VLZdzU4+jeebnjwisHD4Oknojc0ZPt/21ZUpIJHP4vMxqV1rdDSXKMi2TVO27AdO
dadPuuTx2ACupYBiGFvA7lVfMQKqO+f/rc2tfc6O4aT2GDKgK/drAedr2NIluWWH
yVvD9AP50te+/V1u6i/KDIb74NUsR3PkIXfKQNOxnSnsmzr0R0pegrCiXC3/P2WE
GKnaUAY2CnN5+JwkHEqepK0B3EU4EFo+/+KUrNwFxaLHWhdOKV+2wE84dAlyZdbG
xGlyKkK4IvBYSDKYf5susjy+3AAUOsy+L0HXb0SN+vnancccH3N+NmSwGvmgZdV9
hk0SbTaO1/FKacjw0upMG3Nyq9Wp6blhDiL5VhzKF4Ecqa7ga7gcnVfUCwHga3B3
8k40PEKC9Z44j1IM1/KP8IwkjFz3MYiB6Txlz6061WMw6VCOiMUopV+86Rz11/+g
CgaaRURBEQwE8H0LVs+RLH91uTluEXx2wKwlPk3SL/k+4Rdvn8GWt1WDfGX2Ss+L
/wXeh4mWAONoe8FrT98tL8Mhw1o7PjTpYpnQ8AlESmI=
`protect END_PROTECTED
