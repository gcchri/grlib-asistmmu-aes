`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1nKFxYdz7Uy4QMsof1dJmToPvwEqEgvKkrtmzE8QYcEEjwnFJnlrTIorYSt3yUkK
/PKU/ICiZ6FHjaXOEdc+C5BQLd+3u5XfIUmZBtUuXR++9KO27+E5gl76d2Zo+mJ0
/nu2TmLpyAneeVOSTGXxOfske4B85pKs1MvgJc0ZEDw8nzLVCLUZinMpg1+k9vwn
qtUjJ8UAAIR5ncQdD8SSx6SQUR5FZB0w1YDRPp3geQKATwDd3yGjWjbkAQz/G0dT
UnF/CKk+uBbTc3r4LME4xb0XADoAkqLvfp3ZSr0UoWMu5tyyLa5MngHncuouOjJ+
FYFy+m0uFnKAVi2XSXdEuw==
`protect END_PROTECTED
