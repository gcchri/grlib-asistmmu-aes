`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hlcG97X+wt9/wuZ0yWA6fxwZnpFxk26tqiGUmiyVMQ1CTZvZTX6BnheMMtqaKQnv
wX0w75brVmqqNVDtPk5BATRcDnP5EOPz0f2BWKE8rXtSPKBPx9wxBYzHuR2YtMZm
1q5SSGyaOdI2+jpM4VSfAxJwmchv+SkVrk90m7rtqYHnZufNGtwQhLxoZUwBxTr8
B8snoO6ImmuurwLmEXOVfpJ+D+m/uc7oLjsHJhpi+9T+vmEOzNLmYcDPVjWBMQdj
ZFMHURuyLNfcblz37OjZqrxbA5//dgApzzS/VkxOZ+0IAQBo0f0ua1MyUi/DrcYl
6/ptfxroqr9+wNbuY1e1a8yt+miBvgEnQflE8IlxCTDdykfclXxRCpYL6iHh60Tx
tAcDnOARa19xbitCnIFuBvVNQawqZlx4851Qo4zGiGsK84I7I4cPsRPibtdVwupi
Yx41Bj/Cfxzg5b90nP+rU0XTFS7ANBURnk0mXngXw4rhnxymzGbqrq+dCFLU0jhu
X6TXryWUuRhjaKqvvF/mfNjbCksOPema0m8twXMimYQsNN0mHFeNQhi5bO/57SGi
ahYGO1N2pfPD4RfswmEF5jShct1VlC6AXSs3odKTXSfei3BG025TaZxH9XWcEm8J
arNyzaI5V/OXrFTIN1FP4SA46RkUxWGn3HtCRiMcOPk3b7pIBJ8GCbR7iPOXoVso
vttS0Gdks38JGhxEcVA8y8FcYPMQQD/s9goj2tDvYw3CbxGtI4ANUP/SixIQ7P0/
PvHZeu5HfhRbdvZFh4V6fr4yHnx4ZXD3b0izk3XigoM4KBVkFly/WyRfw3Sq2Kb8
G+2xFTSoFMc+XLt25+btIarUjNF549U5fV4lRejWP/pTSt8KWm8q6sMQfwiCqLpT
5G4jjt1FrNTA8564LeEilLPlxt5KdEcLE+xED4zqLQA0ac5rlDZxvVqMp8TBXvrR
K8MhAXY+59lmB/69HXrVJIzvH0Gl2mqIVHSbJZQKthnLb1PZmT75WmmC9Uv0XdQX
S0gFoPnvJYugJR4A+XjjghqOvvpYSic5yY5aNEeRwGulYMg5zWeQwvg2tzrezEPy
QHjJ7XHLx2cTZkAs+K7aBzOllo54BLlkRINHb5qqYY5628BE19f0FUWKCbnCAIYb
ZasJ8RZPqFRfAIvMAc3hsYA1Ob+UIxy7iQ0DALlR7ws3MQXeCWAf7wb6N9qhBMQN
rZiyFXfShl9Ot0+yGNZBqT9hDvqmwwCmLaLv5oIyXRljSadn2r/Zg8MQ+WyuCLaf
kUzk43TOhXovhhqJY1TBj0GZXUC1j5Omev7LFHx9mBj4p0gbOavwe3mRWySvTZqm
tQ4T7hqbMd2rLp1g5lh75w62GNhemES3EZzK1DrRLDj4ws4jTeEdd8Wg+eMYkTRR
uDS66JXINjjgRQY62Rp1w9vVd0iFLJZC74OPSfFrIjXh5ysy7jfnAjnQKFDvFZ5Z
9q/DQsKnic/jN99B8SXLCToW9IZHDrtXh29n8kyi1l01s1r/a7RB7tWU9CfUOvE6
Wkc/VcxzJOYaZFEcw5n6lOn6340xCgBauntgOtYONpvMq9QZzF/uIDp38qsYExQq
/UUNO5SmK/JGhBXlDnP2mukR9Zkv6hTSlb+MUdOasCmcO2x8K905ThxEha5TEvE9
/NUri21TUdz7EdRq4RwHgzolspNP5W/vdGbcvOWCmPCAQ3SLMLhAy5zs3z7LgjYm
L8rOxvkS3aP8QiVPysZBryOw+cQIO3xw1DWb8Og8nK4JUIm02e37UE2SC8K8yo39
ejoFK+xnJVMkSeNJqWb/j1eHBlt16LZPEiZg0VOFz3fn6jUcpVuFQrucl3SKB8+o
8q2e0VUNLfUqmQDwvd+hIMWCQ4MrlsKyeZzfQInQzOoxMx8VEhFoRNt9sb7C6X9S
/ZmoPbjMeGFi9d3HYpZ2gqgjRjvKz/lXs+mHWgRLZ6QaSZ9c7tUa3ipgcNm2/bYH
8vKC9bp1kqEJoSsMGRkGmyjZzozjzq6WWQbGsquKA+yjqTS8uL59OH0X2q/azO5e
QRONzLugOB8j/W1/M+DvuYxEAvQat8Z9wyUP22EpAEe2BBRlsm46hhP5PuO0266O
BNNSbcLC1AYyx8RJmHe4+f0Pizl5qpu+Aix0gh7L2P6LiBQZx2KVwzED2RhKPDd3
eHveoFnDO1oB3hxy3iDJ8ojUxF/G6OO9GO/5cQ14Hrvo1dX37IM5LlM3GFrlcpG0
ghQttbPV68/eEC1ELouCKGFGL6MRUtIYLgQOPhXhG4/DQj0FVepbvlWu70qNFBUD
HzUv6kdtQSFjNBFGDhnJz5lR1yeyGZpBIvzp2+1iAjgnont1Vzcp9ubXKuJeEwnj
C1skNu8JXbf31NzzcoCTNelztp3TPwXEnWag4SBm2/ayubjthXdscxPs007XCAQ8
xs3eSObCw8YYLOrQy9uetA==
`protect END_PROTECTED
