`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x+RIubJt5gQJDbG9SuwOynlB+ApIIo8/EjlgrcJR8wgATIO/IbAuiF9rgEZynGwg
HcVYikQAdkwZytYb1C6lpaEyIeKb+Zlsn6Q0YWTJtge1iOzHmLoehKp+Ba6/ZY0D
pTwKHiUu56o5HiqZAH+5JZm+uDzTpejwI0Y0f5JWd1VsnkI5aYVCxK2PRYGDPdiZ
5baY9jehGVizXHgt4JuShcGoRuDgLKnaLPPsa7NRz0gzjqopjD6V9D2rpJ1aNRCH
2+pC3UafvjU8NWkhostcgKnWRfEDfgUgx2/yfHaASpCVFDc0VoDvqJxc3qggcFNb
bvIUmJhbMpbXj8m+7FTnjW8JBRh7l3NRMmx0RoDfnFywmiQPDJM/MPsuYMLKqXbN
8HJ4+v6RFgvt1AReqD7rR94xI9ALPWwyBtVendJtP+Q=
`protect END_PROTECTED
