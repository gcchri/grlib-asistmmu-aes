`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HqojAu9NMkcjhV+6C/a62niOfXcBFeLPbhlOqstOx3Y//7EEBhDXB/T27UUZ7GnU
kqJ928iTuvfgike69v6VWXQpKrs7a/cTGVOtZX/ezYQhLgkun12kE7yC83BXn/IE
boovuNdUgZjdWHw3Ed3M3seXZaj+SbKWJqfWmCNCbBtCEyoMtw0kp8y8Ot1WFewU
FNpOE2UiDW9qXxuUNR1IX9SHU+qJw2DC1qBMVRRzhkEir05hv+e6H6TkN6W/kmh4
UgKwX+Hj8wEk1WhOCQ25i6cqR5T9RRmdulXiaA5JTBRBPUF21bf2JqE/2G4U96Ae
t655OeCdOfREjrLrjb8sLgnf25o9hMa3ggSo2WURpc9xeWz1VQowBbyWvLUuxZXZ
UVvOmTPbRVIoA3wJ/en2eKAZNy0f0HL8IAwgOe8L/swbkKUUSFHUm/OrmHtAdEEX
W88iEx7qunJSB2NLw978GN+HMg93DsOJW1nR5apn75vRYrjvOM0Oi6dZgbYQEN49
W4VxY0tnWQiRx3ZvMCGi547nD0hFRxlOio0DELxvJYELAy53FOeXxOzMFIQwlMbk
E52tEyz6vznPdQUGuk0Gr1iOKDIqUd8s6muQXtCD4O2ekXp2onfqCILk7SOb2u8t
qVpbrQbxjQb1VAx2XE2RfBDz2deqezmt4BwSps92NyptZhJrrTWT9UVZXLmVCsUI
5ZN2MrPyhFGZo/87W/UbR4VQVuBJSSJRwB5Hn1c61FPNQ287OCg+6eg7uVbs9ypA
ZzZVDyEICHKq06FZEp+lL3lKckgmviIP9cdq7kQW+ou2W3gLDaLuBZmHS3GfrIXu
VYv9LrU/8njXHOFjuB0Q0ugy+qKF8fX/sQ2qZFESV33ti/Y53VR4vMxzlLiKGA4G
wCwYC6/Y8dhARisvJmqYQ+G60kHD6XmpgVp1QX15a1G5l56E9gDrRVxbeR4VNPQ6
kmXlFF6cD6mr0r83r9bQEQtzsA1d7Yp6JZ5EVjdrvq7A2vAxoRCaF1tPimd35+/P
sBHsM94dh+2THZboVuMCLlwY9aAcV+trpgUjF2Zj0ZeXFb9HcfV/XOhKLUMtgMnI
Qt37/jdpVZZyi3T460OeZ4GaGPJTksaclrDCoj4Vjo4+/15GIUrtS+9pmHTtnf19
ojdNrhlVulzEZJEbF1O8AfN+yCC4GRNv0Zgv9XblwKvMO86lVvmOjkc4FUzE8Lf+
E1CIPhKzZ55qn8n7T21KZOK7zqdbk9OOu2fCY98h7MeLx13YIuDEFItdRqVZ+7T+
HnBdjHIDV/hen/Qv24Z5KCxk6FwdvNeZTy//9M7l7hcButUvqwES/FsxdImQQSkF
huyXDqkvl+zQba+lp83e4wOdhBsY6epHqLJ6fneBg8c9tzzu4gqUQhP8CXxrNyKH
99FB8JG8b3/eXL/JdRh90nAaGSwZJF4LO7KJEOjHsZVm5d5YHO03qwP5Ju+2DgzF
OkyvKBCspjl1YmPZYEhS8yhBWOvSgMKkTgMv9UQIZLGlG8NhNXW1RdhaRx85LNGI
0yQaOAEQyiZg1sZsi7Lbsu+iIc0bNg+Iau5hHXKwNpymxREta8K5wUlOH7LWOt6K
JgIFQUH+5w6KoLsHiwOy0RYOlyxRFYhqb9eqARgn/FmouZD0gslpg3VPsh1EQpAg
qq0llJjyc2sSnZLIlZail5LBDRTCTOVdEWLrJhGOE8WFVR3LgpTaM84cvEK8Tkcc
+kJLekr285SBI1HaguwT/h04FPv1kID4guIq+KMmbpbK0/5z4CaJht/gMVsyEPgJ
MEW+PJuc7oh1XPXEVlZUu45opQSzCkJIRna8VN43akn0JiWrXB+gMOhnunm6VYxY
6QKdEuGzBhLhzeeUeGyyjvQBdUTCiuWRNEvlP0kSAKr31aFn5sSf2Dve5q1S7Hfl
sS/QQPQG3PkB5lFO9mxTATTGctVB5ACmf4KYUBSFdp87nu21qkNMpiyOWYps+xGr
VsKDbg599PRkiT7Q2higBJjmlr/dhEF3pEt17Lp7gPdPKC0olFbrg7jvLmR8Sz4I
C0ZoJsejQ7m7VgNskuyhMiKX+0lqbIiDgKc4R3WQ3e3LW5Ns4bLMSkQv3IEkQ2Ky
bIpMP8l49+u/NqdogYtyIWbYdsn8Tm4FV0qrbB3uA7IcvUzqD5E/AwxFvxiBhw77
PvuFyPbkwIT2MhLsm9m0w3Kb2Ete5/AofXwx94n+2JBBH3E4rUQ97kIVjwkEMklX
oPjI1NAkyiX7g9kRzfiP90mYl9gJgLtqmjIAiNSASQpS8xGP0jdLaaSij5ApBtSk
1prJqe2UbUv0JLm2JnLI3bdp/CUggxZjRAyIRhEYK2S8xpcUVfDJpK3OxnA4io0i
zM31BDXg3AdgnSLyzSHOfnN8jBBVsfedu9wv6ZkNK7QE6yAKV2zP7Sk2zqnxM/ef
f43vxkK+0SOVCtT9qLUM2xpqABhWZQ7qgvIK9qVoQoEAK5qJzaNmgVliMSU2Vgnh
pwYOITQGwtDgs0i6LluBmTwxwg8CCjUbMYzT5nRIHM9nSqRxL4PVoywrRgbDpuWr
0VkOEuQabiB6Z0ltFo58Gl/p4pXkDjtY6GCFXtvhydA=
`protect END_PROTECTED
