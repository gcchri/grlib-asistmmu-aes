`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qXw+obDwARKU8k8kef5cHixNeWaUIIuSKPG196QqwcxfWBHulZVcAO5KiCre5K4V
zVD8WJNJnOp+hPikB/5EUBs6lN4Zr+/c90G11ZNBQ2WaIYHfyqSggmw+VodXoBIq
TxLtKRJNjdBBe0L4TkzkjLRRJEQ+Epv62yYAOvyIc1S0XWLlSAIw3YNdyorjVTX6
VZ7Azdu/pBw4zv95KJpfLdehQK5wXuyx8LoDBE5sneGjxUrmKzO1tHVMNY4aki6d
U8xDTWVzexKYbVRk+259mbGFrH9YL/ALZOBqbzEKn8/Ic5lRBhJf37+8YdF/0jvk
tADopQbwM2OFPTnuX+VRsNK5Z4Z18acD8EhPORWb5erFrzZSeNY0mp/nSqvX2a/3
pH9n7tRH9PAvhD5kom7FnA==
`protect END_PROTECTED
