`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+SoyDyBGyjdfy/9xc07xkdYFUdheM1ksccwvr/wzMyHlU+nYjTnEPNmKaER2V3MO
w3yTyYJN0jRClG9ArQu/LyjuSNqjVsU2bB/vyyWApCA417ssHnrqKd0pjccMPybd
nV1zMxIGV3gf9FnvVDPzZkiD6RYDzFAh1tKTFJAsWNNaMHVbGFerUjOyqp1JV8hs
6Y5wUmIvViUgI91F99h/VwKQ/Hff8fcy+8P0Xa9dbJh4d8NNJw+DZDp/Y0m3+fVS
Rb9rrnnIHXDyyZTOdAU4kQ==
`protect END_PROTECTED
