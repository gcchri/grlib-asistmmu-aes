`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DQo4VsqMQlaT9Yq+aQXDfIkpXoVo7855DD8lvmYnCyd1p1h6Xfkv6vWjQKWbKQVt
30pESn6LZzwOB1UI8zI4C6jsx2jwznBncBd9yQSW/hq9Bq2u0XwNU5GjbhYT7EO4
UCxNQSMfrmKTpUgZkAu6xNTGHVGzlO5l1dWwtwLWOmZQ8Unum4MIZzg98zPvESO6
AMp5sVsPkHuio5Xf8bLHOk0skKMeoqPPKjynCxb/lo8NCyjngm/fEJqGPcLqE9bD
Kb/hkaLgjc80hT/o04hFWQjoY3KINGbFgB/Wb3ILUKEOVnSL2TwcDfPHAGF55ZJG
Mugk6qAhevCCIbs0lEc9IjdcBN1qR+uYiTqJ3ypdWWRrrQebZL1Gd9glQJ7DkIrb
IEnr/nYV3nSqWOKZp7EBdG08URCxQw12fDsaAsrMUO0A7qiWhFLI609o7SCLzGi6
HmYS0x38NoMHFZrOBCPb4S8ia6WtA88p5N2zVIOKbrRosLHhmweuoxKzFmr7ElDU
YydSGmikWgss3qd6VhGqMr3+bKnMYYIUxYpKNNXLj4ReZmVOOwdnPqRBn47r2HF7
oprOkYAFq7H7m3zfV9rU0ksO1fO83+zGdOKqiV5lGDu5h/WMqFCzP+9uX+AE/SUK
mhUEJYUKpYW2h1IREME9PrDtTlqd1LywVk97OTdL47EhsfBAJ08dhyLNwwuaM8q4
ILQIB0W5LEg1iAwbsPKpK873jyOnXVujUNSHnLDNg2khpSXqIsrULBBMl3+DG7Zf
iRoKwMtPJOUSOhKcyEh+zAGYPsgK7KxGQruGlyqWFQyUSe7u/yhItfZnAtW/myeI
Qs/fz0/aYfqDfy9BmOgmReh1Pdm/cHzkvHulRo307RS6ZeYXXXUqqogWv88acpp4
5NI3kWBsHWj29/b7G4vUehv2VdeaF7qpVtg11VPGFHiGQLAkDLoPtVekGukCTfba
MeVdP5Op/YFExbtiwWmUvDU1ZUGt/WYvUJ376q0Om8hI51O33kPct+61N9edtm7E
pQJCO2trMZkdP7JRd8FY/2jNS9KO8ivr/cTlsO7MsN5m8SmxhiczzirTO/OBWckk
Ef8TcMhNaAnhuyoziyv+pwjVi9S08PTNxuQZcGNlT6PvfTnQeqWLsgC6yfwMYsPk
NEZeXaHS0iEjitEEzLiDTfPouzo/HgB7QsemaSY9YIV6bDuPjX7QgRhnAuQv8eom
8CUF1YBz+UBD4ZowdCcCtpUsIS/KHOL3AAzV4ceJfuJoGmFt6BUcX5iG+RQu4kYK
JATfYaB0DmZqQl3VFx+Ffw+bOysS6JBWNmCc9eT3jGfHe2OW4rPJ7icT/wQajkn6
zX8YHSfU73K7+AYYytJP6w==
`protect END_PROTECTED
