`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7bihB5oH0MSjOktyV5y8phZoBbzbRrGpwAdiAyR6mmGPLGKXuOOcRQnxuw3ZPPOT
dJPsvtMv7ZEv1jUwW5UapjHYcnf/7fE88AT/9lFIzEAp4H0AtNvNbl/AChSDgrIq
ewvINlljTTKBQ+fDWpj6IbVZ943K/ZlkqaN2NFAs+rnLJlPRfgHwlL/EHHJbFrxY
At2/y03o5NWzgGj2C7yhWD/ESwQMWf0dL7gtgIEnTX0b2Fn9NzViYxozPUAvEqcT
dyFf41ZLBg4NOQ2ri76SE0Z+nwKFHhp1Sm4yBRNkrWd8r1K8YoD+cPkubhTWUOeS
8TiiIqkWJdqoCtlQGUwpE94egyIn9f9/rTI8Qu1HmVzs7nUkG1hVI8CGKl0e1bar
c4IzhwbT/e8mAlHY2atM3O6LeFb5IoCK/oq0h6RQhvtZwxwk822VxziYqPOShJgx
`protect END_PROTECTED
