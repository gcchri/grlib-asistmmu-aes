`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Am2egp4pIC2re0WIWdTGoA/QSpB70jM2uAMaHI6BkbAtK6UMTEHJYcbUTD1dyKj
Romu2s56GhSvhTQJDuPbwcYgedjtPuMHEETcKyB04spPmFfdvU+/1gwIocIlOnfP
V7AHU7hwR/PU2BvhO9rrdKeDFYxzdm4jobOGxry+xxLCy/l0eUSM0ldSnYPlPnlr
fzKS1rELkmVTFr+IBCsL3dbPnHc9UMHXtlgJ/SNsHoeV38QLs1opYshUgSNFBPSx
`protect END_PROTECTED
