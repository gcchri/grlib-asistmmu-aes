`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7zPryfoPqyIgTA21/8lkB/qWDE2QRH8vx6gJS09x0oWR/d13JKcJ8tVWAhzKMqrf
mt3YWK6LM996FxwRZD0mintqKxdjTxEbwpVqlSB48oC8lVh1vu8USxN2ngaiFyeh
sKFb0bj7/6548J0UN8ofT4ubEX9ySdZDbLVrl9HVpKKmfOc1XQGoq8oluTNHc/YX
AQdG4aicwVl5/cvDIM89wQeJBixuav9P4pNsPKo3KIIOIcGUCSbllKniRJYz9X5D
5RuevsAGja9PEm+eoTfYQcv45jCsmbd2c20VkR/EIVA7+KFlvMqE9HwgMsys9sEC
z9t8RUr5NkVBLiSiUumN1RyHvU5K58OlsKEL52Mo4TaRgFCWEKBZBfDkdwSyPQ7e
3e0Ky6qozNgnNUfArALjIbY96CtQsVfoCQH+UaxW01UCufMIFOZIhJ2gOkbYketV
84kV4WuAmdlRBQV6EHDAvQKFoyMTgnCKFv6AEw5BN/7Cqscvttbpg3hv2Px65nyl
gOR6MPCRr2kEBTjXQXuvgHKPps5yVQT56bSZQAeR6hRj6KYRn5C9pNO1P7K/y5KA
ccVulyoE/AMZh6LQKzilRzWC05FNVJzOol9ozBygHCDhxSLsPwHiUQHe0yowIUGN
jiZcrEyl7hML8zl4vBaFLRbPw9rPmTxUKYe5G7gJQTjWskfilL9fLdIHjWkmHwaf
rb4fnvA55Plbbp/6o2I1Im9s6z3wpUpf4pF4kxQMhLgSLxQtWKfxEg2kN8DC/A6P
I1B2L71L8vAQrttGp/sGmRWoL8tK2GoG9g+5spHLPhQL4/LPBxYMF/VHgCw4targ
23PgtLo2dvWl3xYB+HcXeONUA0nL1eKHNjBMs++JcwaV8QzyjEQ6N8spdIpdZ/oS
J9lRpYb7+XFR9pv9TqruTXBMydB3GdWNNhMcxbkGgoeGrfUjeBpKMdrtgPZZflQO
GpZx6Jl8eWwMEX+QEN2hIdIt4eaqqWY7CdiDpqP2S0z/DQ/A2SrBRbuHHnW553mU
W0aRXcQ/6BmITOzmGcI/dtMAXbueddzGDS/xQXFGM5qUqb8b0TQep1tKiLHaslQb
LYckpFgPvqXQpCWBEUVcv/lqElMbY/vHwSC2QKHJelnfitai6DmWeYIcYY1w6o9X
`protect END_PROTECTED
