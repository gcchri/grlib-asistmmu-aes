`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cXqdyiwqVUegsgohbjvD8M8GhXfo0fS9r14owx1EzkbNo4XvC6+iPfojPBUpnpqH
dv79sAVKhMuXyjT5kzjTK+cbrvgi+l0JT2PAf3j+WPk3/4+gOrhzUAM9Vc7OKc86
AeVbJqTAmXq6rkFUkUtEKVxL+ewGjsylddx7HyofyLiS7t9tto7TQfKrbjWk2pA+
tlG5X6mXYK0B7P7MysIVastAECy/Zg5RA3+ePXPylYEWHpzd/ngPimJDD2AKSY9U
rxzRRSTThVlo92klHuXyrmB75gVprlGA6NtyTgn4CDY4CaLOOsQAdnuO2htYioiX
ZMXBPltWmvoHCuAJTdKLRA==
`protect END_PROTECTED
