`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uvAVZWW60eEZ5bxbxurTwqemQm2lTvEKc9PCsJ7Vq9kWq/wsef5aBSFm9Im/O1PZ
6lNxZuXxVhyRnv2d3NDqxpric2TtqGvt0Q/7NXRVvQkD9X5HoN13JaS1v2eqCpJf
H87M4TNY0gkERwXZrM9JpuWgLKaSW+8N9/AEZr8thXcSB2ruFbA3SuO4cPrpupCq
7HNPGk3eyCQE/dbE+XNwICD9HcZlXELhNtWA2tIVoPny3ZxhVbZAnvE9GGTcxZ3W
AhuqqVG55/e7aIi/Pc5FCyrX418z/bfUJGrUEdCO4HLlcJHyfugFbc9L/cwGSqEN
SEYk/AbwUdVuwFNBsFdtejBpg2oCcnt1iYlQnoxcQ1j+jF6w//qb0rGYHrbak/xv
kTiGx9Yo/rvjP5QZaBSlGw==
`protect END_PROTECTED
