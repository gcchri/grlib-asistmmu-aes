`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l8QxB4cd6JTC/dVJKQa9Hau+ql05rys9mbowwr0r8vnAGbS1hQ7KMQe1z4vB8oh9
2H9bSMjRUsJoGCPBO7hlvel22/tRGh02PSenBPP9QhNV86uYE49Kk0myAnt+Sdrq
YO/yDbvjAqiDryNnDRe6Pt+uIV02rdbJoCIC1A/itYjwUX9pAlrhNdg0PRlcJuXG
Sj7TrFfFcl24p8Inq+7lo07UQ7u0x5lIHkVkcuKKW5x5Crb99QvlMoVBrp5fEe2N
S6qhKoiPG3K48RdbDzwBl6yr9LomDCuJ462fsNzXd5IQZdPfAbwiTX7/opIdiSQa
OV4EGp1I55UUronXqY5x4NQOqWfMP2EEZ1AgtK9lk4FzJyxyZHoegPjQCEBEFqTa
F2mUJzHNXluRFo+PPu0rOAbUWAu85k7EaKEnyUe5D/F8QsQXSbwCZ/Q9okJwAoGl
LCso7NFrk5FHvBoQxQZijgQzYa9TiaI1KnttNLZat3qg/Qb3WjCLKYwYKeK9HVtI
`protect END_PROTECTED
