`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I5KWjfYJqD8ntl0Cf4gRbpmqVsatavBsiZPaDB592DCA8BH7vkcAql+axZPWaJ5M
JeHAbgguny5dfiKgVrd5b804aVcUPpHV6Hoo0iet/XSboTIK8VkvBbPtXlPDaC0y
/dLDbFZKu1aqgEE2IzG94pF6yH1Tu5Pc0ypx/VE5V1jRmVRU6O/1l47BzGTU1nOQ
c+uqbF3F4chSsW7gkZUCSixqvNBZ144GbC7hiimMpM3YsHiO4G7zwvE8J/g4ZqIH
cMIZclVnUA7PnnBn8b4nTM4E5KM5hPVvrzRN/w9c+8vUy4mc8FbEBmFTo/TFGPcp
`protect END_PROTECTED
