`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YxKPmUd9dlBI5unF85W838SHy8vahIWUxYOtI/jVFXPV8DnQYnxtsVVQ1jLRzALX
5PWOo9N8oB4KjOq5nXOkypyeQgkm1MPSPjQ1xwx6upqFzbnCmrHqOyDGn8kopNdc
d2onR/wdUeL71VUqRBimkumoCfGC/ZdZDrDBpZqnUkBQwDl8xDHboxyEj78d27K0
FLpJazzrQ7lDJJ/rY6PpH9lTAf82ADlu6BlLo7V9NAp+GwliLQGr00Lj9jno0GCt
msvnGXmRbbhOkNbmKIuKhXECM0I9lf0sncKBYv4jUxXjrriuJIY2kEBFyJsx3qwA
KBPtIxcI3bPVyyhTp6PHwO5BqQhYuUa8u6vYWE3FAdnX7OFa81/sJg7trE2gzRH+
rjF46xRs7miQDKL347njD7k1DsQ7l+I5t2lu00gWdDE=
`protect END_PROTECTED
