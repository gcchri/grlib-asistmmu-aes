`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
32sqbfJ6ktKsOHzfLuDF8JAlmi+gvOQiq9Sjw4S5u0Mzt5ae1U5Ohu8KtqDNB1QJ
G2YeUUfzOFgHixjGkd9skVXtwltumUZc9y+meZ3dEECvyQiaRR4QJa1c7Gox3Uvc
Ni2gnA5A4jtejfF0EbObnQNzhXe4fxYS4MDWi3fb5W93nGp24Eo5M88ZTt0TQYRW
8++8y5ct+YEqwZYCmOrD5vaIhO9tDcx+WFvIPFAIx8DmEF2Y0pre/67v848Y/YhJ
05W43BCx6VnA37uXu9MrT5sGNtLNKSwokq8tbP2yRn1aOHngrxIW4XGG+ECh8nBS
LjzfhkaCtMAUTuVgIPQH0vebSiBh/TqGMFDZHdzINHO41D79aJL3kLH8YTeAjroy
`protect END_PROTECTED
