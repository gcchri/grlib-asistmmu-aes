`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X/Vsbvjafajm93MNORmtAgHQiUZPSBaplsAzdzKdbUqfqmKAcleF1nweUzuRYDNP
aqePsuYko6UwXOmXNulNwdQKq04t6sEdXh2MJpEGVR2sGSwBlKfXbBQb/EXB3Vl6
QD2k7tjwzEZqP3eHxPHfjXFjJndK8PlQRu6hBSaPZMX3H2ukQPIwx+w7OIF2GG2t
gf+jyC81OBOEUowPa6KTyFPcVowC7RdbX5Hi5vaHS80MGQH+DIPFmZimKQfdJ+az
j7ehGSawsqOn9G3QJLhCYE8o8V8k7XcLZjjlD5GS341CTRaNbm08FkyX7qRZyAnc
SYPYvWYjxyUS7GAGaSqwpjjgpBt3gBKLIAAkPQI9YdS+nns1YInTZfBYJOrDqTLs
nDkodJF5Eanu2fmaAxTKaIPb2wad+GymxV/LdP7a6+f5RR1V7vZQ3t/lhiI5A+HQ
q6IamCowIbHLdeWBg4i5g0X5sNyxwlH9RmecsJ9x/Oo0W8uW195ToewFgLOCZnJs
Su+GVZIazACr7tFKVI8LWLthlatkunVGObyWbMHaLabdImEb1hRKoHyBV3gpropz
+VwHfA76ey/DiHr0LmUBmiFqQPxIosJv02LkepS8mP0=
`protect END_PROTECTED
