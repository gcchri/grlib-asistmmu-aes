`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
reoP+kq62fcKcKtCx1vavOsvAvZodiTHB7H4hNPZ0xS7Nnl4UCsfKHdiL60abFF9
DWTe37G5IiAsna71gtpiEd8oAoP2qY+TQ4nmfMI3oa9ZippFYk3jvxOrpTWQLSJF
c/nNnUJlF2CUzM3nK59nCuUhHPFg84vWP7sjfvhRhUngdqLvNyANVOyXkQC4q/mY
jWKGDuXqHOdkf6VeH3Pb0e00sMC35N1LnZoU0vfJ7a90Bb1206EzljAI8Qijbj3h
eaFQaQ+Uz7nevWj5Gp2apECLZ+CJ4iWivfY4w3Eh+iKjVXrnteOvrI7trbteQx7Q
5qGmkN4worpol55MZX4NKEtT+V1ORTVBbr79ttHodMBwnkEq3Pm/Jyghja/NpO+V
odnKD9KWsQlQMnRIuMEWRxyiNe/qXi0uxxu5Azt+Nr6H8T6ef0MOhK8To9XWR4HZ
55aAl0jX6zBu6M5EMjKCFjeTb8jA696LI4r11zcvfKnOTUbZYPuhjX2LHaRxKXhw
eQw0IDdE+J+vLv+5KLiJmdIH6x3QpkEuxjJVBBgSbnhEEz4qcV0ONzxEX4VHgSoK
f9Q3RTmpS+is3ibn+DDyHw==
`protect END_PROTECTED
