`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HxVdZxcS1190tEBKPWa5eqRPL58CFOgLDtRltOWwJjQE4I7EM/UgDIGHTFbQ8atk
u9jTrU/kNWAUPwc6081rN5qtI4HCB/hOfmPurpt0ST4czMPX3F+Pv32m69IVoD1g
vvKuYbGdT/ISNos3sG8QitJ2atQbR78k99dBF3aDH7zrq84wMdp4vuUWjXF3gRrN
Rzd8/UNGK46EhduD5zZj80v7vJN75e03N7/k69GCvyHEczuts6ozIIEYsdI/7Noh
3Ch5dkZ/Bceykddxj7UQj8B3fyMs0orzfmc+eEA1xYPuBoJrIrvLgEX9H4YdFCbC
/+MQyC3vxAnSSMaw10fKAQ==
`protect END_PROTECTED
