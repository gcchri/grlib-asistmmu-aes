`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V/CckmiCdMac/GHNHsb/wL9XTw7VOAVfL4QMfdG+a17GoFuY9Uz5vulkq4XgIhAx
Su3QAwFqlcPTY7vtw1tTxEll/Jt7pco9IGH+e2FppWWgVL1kSAz3W7WZUzeZ0NGF
OInl2ne1BJAuG88G9zrPi0pBuLpkCokggZDpdZhCipacypFT7C/dhB7EToqu+iRE
ASzIFeu0S6TSgBOBwjqd1xM/IeVT9OZGwKY/20tqkCAMiuQ4xb1UoV3dB6uS8TxR
sBjPIjptF96Str6ilI779NvKRtuV4YK6etJgt7+qRZaev+wkcWjpj/4Jc2K8be0Q
R35EMEpg/q4lLJZEvSHOZ28Kd/OffDf7Y52CF6SY+V8g88ckN4uxg8WGbEaBH8We
rAxwpYhg5MQlZoD//WWx3wVjHv+VmQVYWiUvZz3/7lR6oyT1+uh+i1xD7xpzdob1
y0jIocxpp8y26BXl0TfqzmDZPLCg/CxJIVmct322PrE=
`protect END_PROTECTED
