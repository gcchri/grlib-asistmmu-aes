`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5XduY0w4NLoEpMn1RPpBhdgtSmQzKkSSKBr22GRaslASKlpcOAJv1J7HBQr7v98B
J4ELrvwlVc33Lbk/U35SmjLFwsRDGNtTg+/hjrXvHqysaTtg9UEA33EylAuTTDq/
dY2GLcV/Xp9yUcfDxZHBc5NbhdCG7D/NQ5DDWMt3a/sJBUC95q9+pIkRRQdMNqI4
FumBvENaNYzI30lNFLKn5iyy5/mklw+CeqU4NWzuAM59guZNByvY3Y6Rnesheygs
TvQ9uUeVkvyZNtLs8K8hmqmzZybqyZ5NeGofb4o1KSiwcRE5n4MzGkysg/5N4t23
BBiBtAa/MAN2KXfJppzmrrZnIGWU1PswDZB7mrj/82dP4szXZNaVvD4vjpKqIELK
Fgbv9mzSCLH3qY0r0rxSt7qKgLuXVr+y+UitvJezG1oWGMI0JgNudAv5KDx9KPqE
wohFT7aBkvKK5QCdfyToE+u7CVCBBkdm5NwXZjAIne4n+uUyPb0jC5fY2EC/Fw3Y
`protect END_PROTECTED
