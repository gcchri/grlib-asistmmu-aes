`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fsogWHQ5QTADWCk3s0/Bcue+2h0GtlLFv3+OC6vQEU7ZzQ0Fjig/liQaUpIjLdAf
LIQi8+k0Pkfh6uezVuT6WK+XlTiyxCJXPwx1oVSKau0ocMmqcshWzG9thKKqYM2S
PzPEmAYoziyoab8vnzLjstdDZFLl4Ay3gl6PYWMra969z3cilQQQkpL88gCQip+N
I7KyX7O07eYNCuGycZOvZUswKcVpj3CeISkOLHjrXz1CofaSh9MK6c+MACnmtI4C
qlnh27EBONiNM4/zOgp9WvjctJLUdc97d9vDUH783UDkfkWR7JBdYvHZbfigEHoi
+2q3GfNN5hDEyidRLDGUWw==
`protect END_PROTECTED
