`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vDNPjR1b+/mvgMufviVygZoVf+ZypX2zfMWd4/FZfPCdSWpNlw0F+5IXucRBBqym
uj+B00JY4GDreD6WBMw4kbXPD3DX6LeqRvvPh8XdbV3y5IzsqI9e3oReuN6P9+ag
ASWUSRtNA8mvKSlxxSN8zARlw3wEwJDXveEQEp0rIOpUaL8MNR34G186M/6k+Bk6
BcVXYvrAmh8n5uy7Ub2Sgf2tbjWRCGT2ROoMpz/bLHWpsco6kC2NwspniHcQj/Qe
eS+9SW9GwizaRX5I9EumNzZkW5nVmeEGyIgjtR7poNZCnJVvXhXQzZhOUbsgDhOP
upLc2CzuB3v+cDzP58dOX1F3RuPzF3ic7C6EZ4xq+xj+F6cCuKXfSVl6HnTYF2Cn
1Ub82GFh06x4rJzBSkRkjgUbFlR0APW83lgN4T4meeM=
`protect END_PROTECTED
