`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2GEbZxHUBdIQy2wuu/DQ1ck/Ts38PNf8o6VyuHn3u8XFpqQmzvNTm8BOR+rGyz82
6luvvaiBJhg5fr5kBpc0KVqxY7UkIbD0s3X1Vpl9AJauMUpt5ci1q2pebw8GSlY4
ndnJNjww8tygzUWM1P5IMk8QupzOxgZ5EuN4m31xgOeyj3i5rxTgH1whlvMJqABw
FhaoI5GRfKiSE5Cs49BU17ct8Hk7P/O+rAJSCdEKJRAqAhdY4x2x8NF0XSmhSvbh
FxBPFS7nmL2ExIbyLeWsv8k/Xt5AgRkybc36lqs455TeYHWA9iRWbOVEVOwySj2a
6hroj5Q8tNmiSabJnUKn8A==
`protect END_PROTECTED
