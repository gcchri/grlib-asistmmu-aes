`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wImnZKMQ+gbr5tDl8GKNlB6zhYOug1aZlpCYymiCG6HshOaXurxEL60O3ZN2ktlw
W4VrC9H5f2WXVEUMxAKExaTIv7yQMDkaSkROaecmDKAHTZshodC1Eg6Wjlru2Hne
9NmEBwia2hdh2stqSoTBGEc0E3kQbre2vY+fXHkDEcWzjt2mWmcSiz5UO3Z8rucW
KBPMr/1J0HEQVZPw3h+ajNqeHTi3GYApPremRbh6gMTSL/utERQ77GL3VRMIp3Fn
MBzplaXiWB5KPSghVptFozdBQGGkqndYc/is/REgOkES0g57jUcd4axbsfewyaKx
IOzzsWIO7d18gQMiWYzZjIZTNVUKX4FB4d+yOF9vdzN3NpYILccLKqUBlJ02o1+C
UZxjWHd13gpvI9qlJFBELwmtUbPZEZX8SHO6jRwRnZheR0fPcVKYQfLXEp9Q780z
KW0m2Z4eUrMn80YZZ+wdV4n8xkNxJ2BLzu6sWhK1qnW70QNINL5gX1R41lxz6gcS
Wf/1A2U6je/Y+04MSJTi49M/W5oyUYx2J/NNJ6WNQa9rUCuSXUOSpIhKlw2Pu90H
B8+PbX8PH0s4EJODA7NjyVCbUz7nnl+qAZaxh6dnXyNVsYDiHUe6YV7Fav6066PV
z87y1rJigMibIKzIW+xx5/q8yWnG+uRhIdiL+ng/rksk4W0onaYykAfIAKQ64iyB
AdTIpiFvEind/hSthkVa0PnfiQVV3E85QEgOYIX0qsZqo9rraqL6z41Y5FVGLTlC
`protect END_PROTECTED
