`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BYmYKQcL/NRoURcZcBEvZToTK2wWkN5q1ZjzhZA5vzlkb5ltOK9yyTGY3ty6ThFA
T2nTg6VNxwINYLuAVmJ8QRfX9ahjzydHEZHLVgC0Caf1NkaTIDCeNHFBt7IggKqB
YXkNZw1KKYt14Ex+Izhai4vx2rW4R3ngWne3URnGwyOjhlqkVpybicV7+LekRl/a
x3MPtaSRUQxFpLrg+J7BQ3oXn/8GaVxyJLPkmUP0FNKIArYLA9p4XfJz0DT/i3KS
mBG25oEGKdNBLfsCMEjpYMCKqSI96ySIvZ969konc31QsTEdfb+guMNUuJdUNDwV
wdQZV8YxZmoa1Xh2yeryri3Bc06A2OOuGdAobnnJfjDQBetO5k/hcqGE3NLvdsn6
rMhj5hVKQfOVvh3C6tnYCzBhJ5dj4z5L+zOxYZCvudHR5CisjjmASF7bv4Yqzvp3
5GC1ZF4nXfMbXQDyNDZIoxjPPGGuF2CG779wApJ8GAHgtxM+KGXa75W2VOX+0+EY
gSf1aKxhmQrshwO4tjGwidGjj27DuIEmMM3APhd25M8Oj8V9f4CvUAeIa5d+LL/A
ghyKEf4mr1vDEuKDgesXcE+A0Sjm3akzCrx3scFfW0W4xVmbMWj62KbDKIku3iE2
zeLjpqXcWkesIEUhMCAZqTE4buP8HpvybPUiWYyf6wIleV79Kl8CfFiA3RXqS0vY
mXII/9QilJ7yRbCa90pcYKVzMzGBEB8azK43+dgiFLPY7CJg8nAn/DFch00KxDqB
OJGtB1anoaEKW48eH8sLzAuJEawfW6nYNWWwObq2QDD+A++cs0VlUg7zQxII7OZj
UaiJPTt72Auv1fkCKTfMuP+y0IZ/VLU2zpExZmFNLVIJiXgj3cOEDzIkBiwtgoZs
kMWoA3wgm15m+npj0SyElExmHHw+Efv0+y7AZRq3IOAOT1cN3nBaoia25Tf0iCvE
Tj6es+W9Ne1qQt3uhsUNML6wDch5eJVlxEW/nbgkNdD+CLRJcOXZiVCafqoQ1ZwS
IwnPYzdQnW+V7zoy0wBfd2F3m917h2Z51a2fr94llPLg4crkQOga7QB7BOyia5zw
hJgCjtKMLMxxGb/n+kya8vjsCindBjL78rAhq6jm9Kg7gWFN6SNdcPqpFYyx5KsC
1wvCgJqZWiI+Ox4nlIqJpZylPWQ18L2N6+3R/ZvLp7skFUR+OQypMPiMja9xJMRB
nt8owzF3fC0lQjMxy/feFn5pFoKnleucXFt1J99AhatDtxgFBxpPvBHXZZCFOMUa
v4/fqQciI7CREfqENyOGmmwDU0IhXDX0TS7/p4HLQNaRIuBkqMSUOYQaN9KedjiK
y0jmDWg4l1Bup9poaYwnhK3pbHC73kgZZ2YDbayDyip98iOvvQLrVL6N17GQz2qZ
Iy8dyus85NFrmITplJlpXMllQfDYR7qslpSxc6DSQKMhha5FsVXgp8kkrcq+m9ZW
5V9LRj0RvLVh0v98B6XlaVtLfa//57i5/S5JHj0qgmvsdwx08ZGBYvLBtYutRWJb
pXufqyFnVvAH6E6Kl7I3Wh3Cg1JrhwUontkU6CXYHNQ6GrNGqGGk8HBIXPBuC7mt
AqmlDmxK3vF7F3zUnSRjn9/ly+IrD/X/SDBqAUv84A1Sq0jzVE/5qmnFZuy6m+QZ
vyoHTxzAVsN8XdMAioqjR9XLEi0a/u9IxZscnlyZbhT8RC7qdKdRP+Qkqd5XCosj
cKVqT5iIjyvPXwSGucXibfY5VHC1Y67RzlZg/iZdnGnPfl0fKOLtKMmbZzNvnNfM
G+ibJ53k1w0/E0XZbbvXuFHmMKAkOCFWHzYRRmSQXMnaqVbCr8awguBrW6ETRaFO
D1auncebhOu/B3GmHguG7jtPrQWDU7SV7rM0uKTVy+tVck2Q8D8+mN/E24kUxE3w
ER9TcxZR2i+kaAnFrNbm3HcYUoagG7yFGLBcEc3cK67zElXhu/GoHdFn2QG7pTgl
fLCbYGjCrr94WUB40w4OANsiPFEGKogKrVSMPGcVjsjGaev0dLNPmOwGexOavTAQ
dFSRm7I4JncehFRhyGeDf/BikZsffaFmEj7zEeWqcYfswKx3C3pOEBIH4Kifg1rO
hk9p1x6U0xoubniZ613Sd2sigSfqxLMqQeAaQVwNe3USQeQ8lmzNvgY2opuPgstA
LZ/WRnCVkL8pGWcTEgD/tQwBEMgp7BatEiQ1lCFYdVMyQpDuDSF5OR8S8lQf3F64
h94dcsATw+YFn+xLvlBiYcMe8StlL8rR3He5YK2yvgcgM5qnmbU7aPhn+yd2I400
PymLfpbSv9ByglJTZ4sL4pOsZZ9qR82KSE4rFfNQKXw0glsbVl7b75Y8zVINw9ze
EKyK5n3AKwODWM8HtxnBYF5o5dqgXOnwa147RJ7iOTyHDLAURo3n/hNfFrB6zr/C
MY2tT8Lx68Img6S1iX0Gl2fAoJ6ebNvQD3U/67E3HqT4x6OHPz9pS24L0Yyf78iF
Pz+6dgwpsMb7CpTgMKNK5j/dG+UxVAJokYziyfws7SxBt0lEq51lwgnVCCVkSC9y
w9TwdiWsWZ3rs+PKjmmKaQU9Tp0frQ9fCctNOMgX2XvNoLjBH3nJ19lNRI4As3/G
eradYtScrTYgimgRPiRHfb1llAQLVI+rBs4IrsNCoxf4aVYbf5yA0TnstvdeFRcJ
FSmZ/8TAynYM8Y/kj/D+jRH6xeDBMjT3by6X5cVImOf2j54KbTT2TnWg1Mh1RlVX
6Fm9yUKQwD2Bmgz9CoUZQMn4Ud3PCjgGo7Fp9v1pEUoEniJ9mDdZi5xhp3+vJVsr
2ImdYfoRsi+U4Iencw6MLflVUZKxG+MrIM+7oW3LYdq0o2UWmVqxMYhNuhBElgJW
8xrXFKBQmFhhxWJu18DHS6Ix7V/HzO1HLcFGG0YRkfxRmadVoaF0P8TPzQD+YfBA
6FK+Y151uCwpRP0E2jLYFhEJY3yT85N+yg+MDKZ8/Os1WfZgPZ1qxlZR9ws77FQx
Dwlj3kCtEF/On8ADLK/e1wLAttTctEmG6S0ZS78aqPp6xDbdD50mEfcLXzWTUquM
iJGDK5/acfcpnYABZjwEqx4cdYdthV5YL7tL0MWM/y9p7HYbChYD9A83W70Ncc0c
71VKy+gBYySQ/e2WvhhFeXLPzL35tYp+vt8NU0rjc7Hyt0Yh9pAbMOrzPujUV+jX
QVLRa4KMNlLZkuGciQsihduEkqC7YL81pV8jzOrkj3EOgmJBhlgej63qzL8U8J40
cDm5dv9FAJhA4eX3tn6PNXmJ728z9Y9D3IYoWRoLnjqjw9P1jeVzY/VpXHiRIOV6
G9zIZVyj3zuHwkr3K9MmYoi/8VtnwM9TjHMOScaZ+Kb55qxTmO1GfpabcUC/l8/Q
mSK8NJW3A4iRZQBZlY/y8V9o1h0L0CNfJdazi2bwseihVse4CuMqZmA4qpnEZQ1+
yzL25ffy7X6nAeKWvPLFPz4Oi/gX4SfNN87aD3OpOkuITI2p0+7Tpc2J4aXYUV1A
uBrfbunFpP4n6foi4v1GJiMLLx0+3usP5UcdPg5l+G1tI4ZtpVzD/TlDnx8jcncz
cFM3PNtCObQ1sB2ec91pA2W6lqNcqwH4h8I4cnHc66smTs2bL6wth9s6Vkb9PEgg
KA7J9Fw0kJS5PrivU75qri0LokT+pjJqlZpGZeDHDttA/enJQ57++lTVlwFownTy
zvbI1AjzLa+tDerp1H0y8MQkH/QldZ7bRx6wd/679IqfQxLfdzay7kf95a5JIKQy
Dhrzb3aIwF4i60TANeKBpOkUfleSViGD3sUX0z9nMtRBRn9ck9hWpudIIs/mk3/q
NkNhc+W3LI3tAb6LtJ3r5PiZobgpBrtD0/FBVgMCKlx2X+4ZAE9VSUi8A2HHdd0x
1M3x79lJdtx+EqIUAUWUm3l0mpB9MXTlIRuM/nUb5PegCA6oUAsolGQG9gTCQfcT
XimHdbsTjVnwwSU5P0taYBBn+sMEvaLO0UtGPTXXe7YFkhLpRoEBXk8YoAB+M9Ky
0Atgse9FjQIk7/nJmFYercnQp7uJzo9VuFPlDC5gqfN6OmISCaBrMZWA4FvNHEnK
Nd7cn+xkLgx3SNo7/xExiR0XZsfQw00Nn7eQkRGrJZ/kswEL0vdKad0Q6TjZRMD1
Vh2bTkFsxQ0YueXUvLTEzKgQWH15mwgsF76SxM3IP7i4zcAoIqB0CcblA/ckwu+r
8Z8r+NArsHDjrz/aHy+PH7FfTidO6e57Pf076W9Ky0uNEn6eKYcrrfZn7Tyt/AkR
uw2+fCyLVYqmAaRD/OFX0BCTkQwSlCXIq1v3oHejZlxLt8qgr7nXRnteNkC3b6Sy
nwDd5iLGklDd63HXMIOfE0qs26t1qrruF68kp++lS7bo1sV6Y2+MmVM5v64gQLKC
i8YlzAnUmDvEA3YsIVH+qPvSoLGJYxB6Li3D0hG6yb9gw3doKYzNZPcFY8KEIBVC
lS8i0F9kUjd2MtmM37J3FqqkYiXmQmSHnXRA2+YJMnrFSWPqne0nKzAAO5nb7Sjh
yqg/Pety5Jr3eBH5JqeNwR1vHktIwzYI2WYQf8bV3eO7GzbidaxeI5PFf/OxVjCJ
bPVElUTg0MzRxak4H5BOg9sPwKPHYBSZ90lek6Y/MLv5e9yxfml9w2hDxq3I+jgu
VvUEe+HLRi9Trl1q3dVg1bFEApRs1tcsbnw8ehDy6gUMyp2JAyq5JVjP69fmXV7Z
1RTfRwwlOojSoJRRAlHAKzzybyW92SPVRkEUInBEtTTz6f3DWu8UYkUV520eyfDQ
47jFb9UZH484KOeR5ZiS0Y8zyb55gn9WtD5UVDf3sCJwh0M72dLu2P4Nxys/MQ+9
parC/kQFdJZGCso1ky2SSB9KKKiSy273+WWF4DOuLfR58i5iTNOQ4RT0IUAQxQGH
94kfGR+MGLqecHtoM3SU7EYsFP3qr9yZTsiQY/xtM+XNOz0OpXnjT0mui5qYDX4Q
6JHeFTgR9j0NeTPxbSHfwUWeGYxKh12qMCVhKTfxgTVOfG14v4JSSc2DXPEx4zVm
mU0zY5QvIanfTkM4cin5SKlXjF6a1L1hJxGM6QZxoDQRpkCv9sB3uz9ctqlSHdUq
2UYm2+NBn1lwGZN532+LlA==
`protect END_PROTECTED
