`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CUpiOEj8ri9biU0s/u/Iwln3rsDySRX4yWWSGibftKQBoc/94hxLhI8yTQ+uGLh2
6g9Ks6hjuT9faqIEWtbkoMYkp4yJTg5NmXlvGqhRSP3GlvEdNZtvMteAe2jXuElU
b+Z3H95mgKL5ZoR7/Yua4pjIGpwIG+atPLCy31CYucJWBzRxWiSTGoxy7VSc5k2J
HHhXSq4hwjnJg8n7k++xEw6csOAPddWeO0ko6qKL47Hu5LxuU1bylYNeU0q6DOZd
3HCsVl4TZV1dTNbOm5RmL5w3nrZs3ZKnWmZZTEq3LL0=
`protect END_PROTECTED
