`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MXKhkOrp3LtUbH8Im5oGKw7ioX9gKhSusOMJsldgk5Cgv6GXAdyrzXzFg2GDYUMG
og/MrzGTxJKwwR/09e7ddRbb4mZ57uA4cYA6T2uo2tiHQVO2j6tf1iKLh5qtDAKG
4OYTtNCk3FtAYgvAUeWIlvjo/hfSM8vy7pqZuBtiuFvwdGfBkau5FEMY5tIhi7n7
OrRjZWA1wERgZOGzRwUfGNIrCfif7kMZgJ+KW71OXCyTsCM9luZh3jzHqXoeYxYT
VUnaSf7xG0dHt6C/26dO5EHXlXgTd5ZsNoOmfgrGiTI=
`protect END_PROTECTED
