`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Sg/3y4jyPPLJuJn5iknLv1e2FvV7XK6tbwl+l/0WPz65w0PO9JPagDh2dDQmOcC
Z/h7wz7xlfYO10qA1jka9VV7q+hc+svVsdYckNZwLOCN0FJZnS0aEQVy7RLkAeWM
9Fw5ZZvXIfnGOU97P5noRjwi8CrgD5q15v14BWztrVc9yFcX/DkUc/SwFGzhzoCI
rOS8YvAXSIN0ml2bstUvdPQWs6xtPDGARXh/r4odh2tAcrYOFzwnq0zqYYR8XHPo
x5kV/+DbJPkD82FEPEwJuHEmwn3mdemyAZFk6ETPd4k=
`protect END_PROTECTED
