`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xRFJqwmJom6C8b2u4UYWm2q/Q+cA5NGXpgbpdwRESTLjN4ENMBRw9OWiSe06YS4w
wlxm2H2b4BM+GIg35iuoeSDuBlMitqlvJ/F6bZMrh6o6fmfodS1sNNJoTRX2W0au
GMLKy1Wre9fVpGPzjyi4w24pWRr5f5bZfrtARsgcDQsOPtoBJpn1nMJAtAo5JxfD
18w0k4Sw2A2Pb5NgxTliwrRykIN363pxH5T1wvNPHWA+TfOtY0DTltFznptmS/Tw
B4KOli+t10HJSXnj8CVLhzDwLMZO3Nq4M45yd4Ygk5gjzX1AscCgyLsjDwk3/lcx
rwQPsDwzNw1YuDjAVZkJisu2vrw5V6JHqLZOAc1GuWKuMwrSsAetk9KHXDLDYv05
Qrn9hkO06NjETqu6Wn5yQEPcU02104/OrCimI20RDHEvcgaXzD3nMFP4hj1F4o9Z
RdwstDmkDA94RVWNFoX280V6Y4yULueK/+ysdy7T1/+3qZIryh4BhRfW06fNgfOT
iZ8HKMH42wlnurQfp/flqfraTUijhEFttwheFA0XQPVBoesGBdZq63fy5zii2Jfw
K1ZSSWGCguyKJ0Oxqa67i1SNd4yICeNrw10qevHryH9Rhlzo+rZNKgR+bCigmn9+
uQswxYWPTD9/q1BGIPotS7KY1hEisNg8nRUaQC9+YTa6aojP8SP05vXl4nyuJrdU
gdWU8od2okFXj48kXG1E/e7nr3FaAvARUkj6ilKrz83J7DZNIlJ0fqvl+Xu4yYfq
gkHuUUwKmxEt9uKSXTYAjTqZZ70P8kNPKmSRJ/83dr2xRL5M2GqLpNHgp3mPYCfz
raKvMjyhsr9DlIisplesmOZnzMsjCV9j2qRMdbF0IJdJ5n59AtH4t3+szMVxrOtp
a92W+mEZ0m03viJJxlZL1MVUtMA091MGQXL63lyENZlyN6YMXsBfmU83bWoG1Sj7
Qhrp4gl0zs1A0sNOXVaLbe/4qA10fynBWZN3GOCHP/TS9kgL/S6L+NyA168060HS
M3SARGQn4BmRYmHA9jNgB4InbNWoLj8Mnzj91mDuBQEO+iUhCutoY0pg/2WB9gLE
asSyVB+Cl1U7OYDJiop0YKjVFSabQDA+I8kY61LDvtpXbMyG07qsusFcsKCJw2O1
`protect END_PROTECTED
