`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zmyDtRGgx79u/cr/vVmutMHz7WsfwHsVTY3FHb4ACdVIBd0o4s65gkZmR8uUKxjE
x1SV+MrxmaMkEEJmJhcacaliNqy/atMELylQ51BX8I7UydX7kjHItIDkiSFXAqm3
hSg6G3gs69QlFfXrTfaMxCFQNpjiNFZIOrLcZXQ+ukR3CzYGHP7b3fGojp55rRG1
5gyRyoX4FAFHwKsOgM9t9rBG+dBH1U/uO2SmVF/7fjSNMMCXCGKMwchPzl7Dq29v
D3/iONLfnNYgClOUUvOCqiFO0rrzjYTJcW4jPrqTDmljbUBvAMKnhaJZhK/BLFlW
ZOhYjizBK+R5Va9sY+NO7tbo0Hyh0sBTRg4eUWYrRt/8yUei9crZ0QDE8yajF7Ss
rT565chrY26+5kBbyPzpI1hwD4rsDKflb1zSyXzJntFjidkv0mqeF/xXDTTbOgo7
nCPGKj2QXWAlBMWf+VDzvKQVuaK2rLRVBJaNtyS5tTiPIFvs1oH91vx/lh27c3rg
saZSHTMwMMylYEbB4Fzpx4P41km7A4IyaEcjKg0OAUH3/KFmxgVf9C9hLuR+M4YF
l2oGQxT4Qrii+uRFtaIEv8CjKNy8IjGDxTKKjTwnF0UWYLfZihyTn1lyOjE4EeSa
KVp2OoBRXbsvvKZb/KmDNiJ4NEd2hEa7NunRKIXstOdemWaoMmI32RxKHB8tJnIr
ndnRFrUN4NzhqXXIcNDv4bLNb8G5zuQHs15nPf3MBb46Itu/y0TppC1nS0ncK0Y0
x/L1m0POJj7ay3U3oZAKCGXAnAiEecItu/NKT7zIOYkl5SD6WuwHaoWGhmHiE2fw
NKYRLOz85N1Sh5zxoKmtmWlA+Yawhb0EemWOxUwyLlp3reQaMWOXFf+lnARxkOa3
ujBd7qnGMoCc52llSOq3bNMhBJ/dIlCIma6lKmcgqtX5wj1Er7ci42funzSnL8kB
2s7bjzdA4mTM6qND0yCHjxF+dNK41Y82ixfPwjsmpYPxUg7RZ1ZmeOHHd60duUsj
K5l2wdUys0fzsfMi0e+7K5Hf7y4lN/77swMp5QrY144LD2QiOJxqiHC7dLNVoR4V
REesWmWLm59HmgQI1OJe5brXlku7JuQJrkIbfuugpE5aOfINePCvXi6zYw8Tst5E
zuxebM9/QRpnANU3U/bot/4uXkhIAO1xx0m0csDiU83eaTT9zAOxLzWOx2+HZiH7
ev0aR4SnizPYSH3dZ+j//SYd8cdYKIBOCpHXCFIRSgj1pQ4EY+KMC5Lob38NR3Wa
r0mqDHJhBGM7cprrsiB3Jk/w3pfnmKaH7T/Wc4xHRls2T+TOVC7PlbXOkWc7Mn5c
YTTjmkofKI8P9j83FfgAXBEdfwf1f5DNVKanG3GYs9mw2acpLsL1H+NbN8VQ/zmv
DdMw86s9xBov4e0+03/d8nFml1332qtGHIrpt6M55rc7akOBy7DAToQppIE8QR3V
DESy6416XUkWmM9Dk337kC3rz1tbDDXCKbN4MKZxdskVDueLGNYrQl3wDTy26c3I
yGehpC/K1S2O7BTnL8K4MBEAdG4lcPIzGLHyzgzn8r1uhH6uL8CvHRtL2v9FvXeD
D4Vz0KBhoGCyjgVVjPAU/UDLH5TCmFpz6WPNTfrtxsbgBdjgRnGpPeeiAxGQrUDw
kb5S46BGnkMZHBEOpP/YZoINB4vZbErQJCXu9l9TMJ2kfSR2SD218v7G3LTg2YzF
eSgIXelUx1s+QEqZnLoiWK/WzYyjszgsLwy068UNLvEEOVmHtztA19yge7kN6/oz
5v9LQNsZDoIvC+9cs72mCgHw8k1LuwnzvnFukyU5ZsUl7OEXI1WUc6h4cXHurK0m
rmMP1y8hXLu/ePRQ5bbV1zvViPDSXgORto3u1iFe2rRaRKOaAJsPoL3fjHi8VWMs
xJsp5jyyNZEZWaYvy+aWqlRjJntaG3jhW/ga9dKCod1tBF9A0UZLD4q3nWzLMZxE
/LHfBf6nz4U1GUuVpgdGXzmdqQGedQTi550nDGo3z3SwDUAwUvaFGSfx3mOFG8wR
qGp16/NZYK0PjWy6fdnN2Uvq6UyqBI5nH+YEdkcyyHGORhLnV1W9NNXlVcbhZBD8
r1No38OmIPgGb4CdXQfj/s11W2Uwlgh/WjRHIW4sSNDEDWsPA8Ba4BFPioN4R0R0
J9Y5vYAOmZq0zuBL6bGvEJ9Tv2RDSp79G/fIIMBqgycDt8B45E+czuLEo4WVQCem
2X3eoCH4Z3ZFI7zsDv7YyEFUUUM0yd9nAYdp8NOvLochSbPhu2tSAAVz7ZkSwTJd
Gucplah8xskA5SjskWzmrBnHXZn8ohbiabz/+zOlmofdxuGwdYcT3kgTzcqiKHbA
c0F6h88NrXH9/qv5iYMLK1a9tKFzWNH8o6hJje+4FtQmAI/+GGLLp84Xh0YsGSs8
FvJv0Gl9pdpVfm9comj2fuDgafGAQ3NwFO7BuwmbQUsjbH+lVirKeOW3esn0w3mH
84p3U+WhNhkTh8snB4rBxPii6EhIMaBuQZIvYVQCdc4QX0g1MgBg/K82orPNeDM6
S3qbqZ852NoWhh7/3HvwH6lEwBcc1k8qE5h90YM0pvR9++0qQpYdTZEBsAr448Wb
mUOncXSkf1UuZDWLcMDxzztj8dJC4WBl8jWP1pXj+5Lvwj98DrhnAACnc9LwVHaO
R+qSO+D10w/3cueWxtYDtcAcSgLwqc4EN7yNgTvCRaRQQ9lq/5lGNuaNLgE0qK8g
NxfQBP11UHB3WnV3A81fqUZBYI1/gG0sxYYZrVQKm4VQp5m+lWP6NCs6jKpbV3OQ
C0mBQBVa7x4B2j+onvdZ2dJWQQaNVjbpWWpPI3ftGQE5qznJZsxIqwTq/CRRQYCm
mI39l1brkrF6E8IfXlfid0c6harhfey0dI0TcKZAUWURP7U83kypBbweU560WOpS
D3CXYNU3hkRfdn/Jab4DLWthRoN4Vs1LwOOK5004c/PuqnTe0PmEIl12T7KhCFsW
ykpfSJbGb4uekCZTMdS2kWtVlf+yzPRHlhhwlgFjP/iroWmp3tWD+6I7gI5VKbZI
+LU+Vfw6lkmNsZp1GrSWqkXE1CI4L713j9SDqcOCUSGhVYLwgz68nXw9QZeoK1LS
C+VKHrFAUmgJLiBPDVoNOp+MXuuHimnP5VnfR3Fpxxb5Kox6zIswJU0vTRsd3UK4
k9+dGKuHob+jxcfT6ZbJ+xpwTw1edxuoSjdsyulCjYkuTrOIens+XzfLk8WUSI/w
UzXoQ1YFQybzPv8/lNFJ7z6tob3z69FqjvJjow0yuhyssfW4AvfY88ONF6nWw6Ge
86WwpLmVgT6kDh6krY3hQ0jRPTxC39zIiW2JsvX9d9Z9TAPhMmzdurnEo4k855s1
pcdj0sOifhkxgcWtxmFkz2PegZfaxnWX8FzxAkp0y3Ib089wFIiIkiNSi3wGdtvT
O1WE9r3+/PBCXUUgmiQz6LvXQnWlh9QsbMeABCweye2BGVXdXv9okIrcbynccW2k
voM7PSAN9spx2hIBkzgMH0vkrprayO9CrA3GqZflUd0fwKVZ2FspbJhLy987Fn63
/Gd6gB6+lfLTnkywMgRon9yvCS9RUSF8bw8BmynGnc5+TngI9FRuMrWJaSqKfhC4
vmj50fbSgJEyMRa5O6RrxkiMWxfS9LivxTt2ru+j44GbNXn0Qq9qwfJ6yxeGR/Du
kFArcqhHoOuft8ZeeI9fyLMg2Y8N1i1o31iZJgsjzqer5UDWDOCDxShPAubsz83o
GiYUvs5VfD4kCswwszf28oLkeR5nGsfPZuO+1EMkPtcKryF2Iu31QFPaGgV6iZnH
UMdpX9bXulyn8deNP6YCQKXiaeingH3wd1PJZoYEP8S34CcqO3NQAS7WteYTsm25
ZlDbMaR4el77CBVtFxpIw3EWLkjoTzETXOCe6ChMiy80NM2mNg3tKRAPWOFcoJfK
nBHO3Az38GodVf5rx1lqHyCavhGjPo0nQovMvMOl7J0UMuxTiNyKewMDKoSByhbx
FiXEBQ0OznX+FWqxtyk7dsNnBusp43n0Og3YZTxGTIA+7k52/TyZpN/kX3P5q3J6
FL7mqpOel2pt2SR9R/U/FSJ9C2I2vuu/C3c41WqHczC2I8Wco8+ZgD654c9o/ac2
7im1kK0kFcnPgQJjntwZ6GipQc2crd9ZNOsggbnhsTf5uV6+DfXg0Hk7R/a0v2Qm
nGdhizHb4WwQTm/wP4kGgRorO3Vxd9P8R3sstRYdC/5xFwNcZm7OJjIstEYxMm49
d2uOgJiKglhAPGqwAiHsiIpmRPq+KM/IxkdyI2JFOgZrpOEfd3uE/Uo/wMTMJbhk
HG4RtiwHbRZ6uTf7AnW89qVO9KADjDzsOTMRvy5UwZRKc0Z0sCfzppupvqgg6mg7
CPAIZ+DXdSZRz9XPyMcQ5wg8d02DcF6rGEE0FdYsfWK2z4RB3iJcvJBDSKjO8BI6
qTXZglJqe6Ts9yVjqp7qZCcQEpdNCv48+jsMvlPx0vGsfnI8TDtqwVn3c8QJM4YQ
ObyQa1xk5JP+MMeLNvSlOx/u9UWoTV6GO/CT5yNH4+EGFKCCZt+iqzN2YbWzmmN1
eJCHXKT0XAlZQ6CCflFLujTLPHR5lGwWj0HsAWymLiSrUuf9prl2D9ecjHV2y+v+
zFSit/MSW5sNOsGBNzAtBqom8opZyTUtd1Ly3fXOJG+vpJ+S4GnmLc2EQtOXEmh/
LcYZGQ4ElKcHsEGFFePl84HCZLAI1s0rSgT/tf4rGb/OiuHCp/Gl/VZAvedrrC7H
LDDJkMO9jutall6ntFACOdyqd9jU5meqUKtSlIg9PwL4e8AIulbbmLi1KCvBN7j8
h5+2TQX448HeHcJjU/x7jVlPghR+VKM6uPMjPy0EozVswbPRHAn62uAVW+OR+V3d
wJ9fzGNkgmBqwS1OKSvUQy2os8NwNPL/sRpyB9PFKly1uQvl2yu68lN3ECn5qRWo
gh9h8KVyz/lcaC+0D4nJpubuyI4dqm0b/sPJfuxk3GKdIS5Fsvz33Bt5YPzqK8T9
0DlyA0U3HJKqaMHi6O7RKH4CbRI6MvGid3FLGXHy5jaj65WJcju2Ka9m5hvBFSJJ
fHapLG3KAYCT943gvWnRwyzaozJMFe8c1cTyH+mO+DbjVRVLheEUsw5rBdk0pUxS
/SptbsUuhN5LKAUKxfyzKZtbBEVhoa0AvMPedihMGbKXr4ZZX/TqSgvi5c66pW12
B9uk+1JSBtwF0u+otWCoJI98gDPfwQviMN5v45VAKsCj1jiItOAXJFwewKKj466q
iz7VMjdegVDstOxtJyiK6W+Itng2QgQDWnSFwz3mzFTE4VqdrNzNvW6T6YOeoEIm
pmKQSaxSqH+nbJ0f4ywKxJInmXfHdFZoYrDQQlw7zBKMMgyWmDQ8ps79KdUGvJia
`protect END_PROTECTED
