`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UOnS0eSay0rtFDEBAU84VSP+c/AUfr5IrPNihEM2MT3Vr+hY5uGQwbwxopJmRYd7
8gDFJdM4PNcRqs1OzLLJxCfEU1UUUcXWsNyAop+nIwBdxPHq22ElKORGPXqpD4J0
lIA7zW59n1dOjC5vV6u9qD8rOreq8i54O6mxAr8towKrWPqT32vxZxwj+y6HDOoy
rgYfi7lt8gIKaNzak+Isy6aen9K7Slympc6MOJnp3CQL3QvH2i8HIcASvGBRKSeN
7LYTT3x5pw2MFEVg4QeBegffysM8MORyAoKqCWK3u6DOCAaH8HRSpdu8HyPnnu54
+VMmLKtjNIytY1VEXQuysxv7INMDtUepLLwjxELxT6UWe+JU4dTwVjx6v8NQgctX
zUlltU+anHDwYJhEVvDhivDuie7mbL4m3ezbVjgGIbNMhOlwZD9Z1UnelfdirAFw
`protect END_PROTECTED
