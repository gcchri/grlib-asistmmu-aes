`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JQ4mjm6Y/d8bhNnhnSe2FGRc1WIkVUTyT2Z0+x1rTBQkFEWsABK1sFvCDyxmz3g9
VWBVf9EMyNmb892wd4QTRECypYckhgTNoAWWw0QEe0PORjYoTy49Z6tBblYC2VYF
AKNvcrA0+ekstgVPZJlinHKICQLuzW/X68LUzr6ZQB4K6qxLPIm2A1PO8d4Jy4Wb
JKtpocBMjM6n00Opst2kMCqUtb0ZFsD0WG8Y28bsSwzpM6+5pu1QbjRXkpihC7SO
LeRb2oGk6SWB9RlDmLItApoGLAuyqJ7EZvh/a6nzwnbcLwrU67nNkagNMm9xSlbv
S21Gb3ykDqYp4bXwOJv/GgOyGaFLv7Bavn1MnPwx6v88KFKgY5bhHpEuSGtVwmGz
Y1h8hicpUK2r4pfWJirsE5hgk0VZxX0pjZFjPj7yrWeo81JEn9pTsgRCogxYpdty
JehJ9WFyIkqLkR7ti1MgA58lKtMRqBmvov7900lygEiH479Jwz4G91WEuCy7PehJ
EPfUdyR941gkikRXZLrqqw1I+EbvxxWe2d29zD10a5ZfkfnI7sI2nfiF7zYRk55E
dvJBdOssdrrRwLB5I61eWWPSbCGsKb5TfBCQxB93DZwsz+MNChM4d0LT47d5HFxU
Ve02Ew+NdsuffHxu4a5qIso7n71k6k13LKXGSbHVtqdO4sehbX7JnjSrdbuKJznu
RRGgDa1/xC0fj70lJ1oHSAaBA2eglzsSqP3Fxjc1/mlbA79TKfyN8GvCZGmXA45Y
5lbaZmbiliYvIoSQhskLlErNFqebLJcX7U8qV5ZOTo2KPzAa9qASjCl5Fmr1HcFV
zRtuL+weEvHPsJGQi3cRzIqOYrg+J9LdqQz8RJK0iHXx8yyzSzOIKOnmaw9a39Pg
nyl6fH0Unm+/A2P4qFkDBEoTc8uZ3WefVZPP9b4z0nAR7oHUb1ss9jFuQT2Eo+a/
m1SZ8OXPccDv5sYVS3u2bn6f3FcSbvYGe68m/VkjBAueMxQfPumSYUBG9+TgO4St
oBZW6eaehf9R0cVJy44LLRL9iXXU0syZYVx3JXFWBCDCrSZQq2mFVAt5K/VG+1l2
Hrq3IlCbqaJQr09zs1ZbgRxqw8jHvBTOssiLsYb9jizGpPS3RMX5823DilScm4rn
ez4BpeJqbBT7ix29N8mS13KUyxVpoMTS7O5L9cEk9MhiasDdPkC95Ev+nlaHtOiw
d1WL1V2rD9ZLinWZ39lXo7S1AWVVflvVrAqEUZOHng5LQo+sdOLmFXroJlZ9YYdB
QCxB40rhmBVybzrhTBWIjLEOrZJYzK/vzhW20/yVxukslb6Ixv9wGCMoUTPC1a9L
BgMtI/mK1ek5JziaQU8yzF2SQh3fMhfOpVQ7Nb5S/bp60BMQYit02fYXWxl5ZL8v
434oGdyHnljAI2oE2E92uHms7AW7SXPd3tzdEz1jBFvIpu01hX1bD7NHe4j6103k
UJwH8E/DQD3tUgcYZVOpgq3EejX/owWfh1wtnMGHm2sjVgaFXxGzeVWUvo/ulFuN
mJVEZhGA8Q/tUi3VQXJY49OqlCghDcLvko4z0OnLOvzOLd3EsQmjYA+pkODYVxva
hOFsfpM6ETEYj5NcssMhFHjMIxvPpocrAMZFeefrXKVLNYuvojZhrVCaKxVn7mcn
82pO9CXTKTE6ltNQsofuMMiJWeHSzZ+m4VCMXIxOU9K2DqaY/Zg4QPWO5D/j+y9G
s9DlRLGkFNXtmWAZ++EaqrmfZUupn9GcFMnQytSm1WN0fhDeZ9+fqggO8tt/OtMK
xr+d8c0vlrBmRMXG0uqKbP9V4vaSAmqk7Rsv6x7+zS+WsdzFhA2BYo63ylze/HH0
OyFWQNX6oI5oDUA4308pcTpquaXvAOqQC5KjUX+yz6Hotv3zGdruSld7t3qox0ZB
tsQxb4x1waPQxI8Gn9bNaAbB1KJq0GGy6yZYpqrdeFnH3fxg+cmSe5IMgipZcHxl
VmhAzH6Sy/LUWlo0mZWQDsoxX4pdy95IM8SZ57VPOPTpxBKpVQvYxnaogqICJvMX
ISGm4jGSJKT1McLPkNmW3ma3pNQDIfqf8Yn7ydu5OTjl6ngwyeIsn62dKlti54dj
d+f81Wh6Z/ZmNjdjrAPpS8/vJmtFUOFPwBw4hZgmK/7QKZ7VIL9maQcKhFkemeJv
qi6019WT1YiY/Ud3Zc2FohR7BvnlEnks9OU1zMKcmm5LyjQptQruK2vAWRyWWjAD
OL3HEWyrQJUkMyrJGFSbzSaSH5Erf+GrMBOuNTw3+Ph44LZyXg7ASTWc8lh3Uko1
L7AzkMhvK07weEbmnKMmd1cCfe5V/AmfjrVzbBParxAghYZC5hxi1KG0Leo+jcLH
Iac3zLJxwDSV3d4CvromoAo3aHh3T7MT5/6nGFnlYxh8P+voN+0TeRAt3n+nBqvA
VlruU2ycdsnPK9iKhVjpl7MKobhcNsvtwzGRRfZAMrdAy41eWu0lUOF42UmQChVF
n5DGKpjokQHV5ofrTXOe4rMp3T7bRs1Hj8KdPmAYT8YgTKh+mrwErsq6Kw9/Xcja
IPFCkXqP25ERrygG4FvFhjTu+C92lDxph9XW4tq8slHERlb9JCsHAPVbjnxR6hD/
gT2E3Sj6QxL/KNaqT6Za1P5WL6U6NunlZj/mjoILYFAU+i21uneQ5Qs4Wxmp49ae
F3kH1flHoNXitm4Lp3jlSV3341LcVto7DRKYvvSz4vJbpxx6F39ZHExbLZbidDhI
DrVThUJOjcUSiUlxH3ehkUCiME88jI0+3qRnYEGILeiFiWQidOIRcp3Cugx09U3T
QO+gUQeUy8wTuif2V414aL5kF3JlwdxKLuNUolZ1Ss6uFvsTptrD2iLRW0F+mZxh
ecuhossn5edSPi9l9HY7C6Nps5qMuqy8ZPXF7Azp1ysCX3elBuCqmKNTvWkLWV0H
n4tt8DjMVcjq5h8sAgEpeakUDhrtGVvjyfptICORPZM4Bcq+OcbfToBqteMLFW7Q
N5/4jD44dNSJ1jftYt5424kIH0Or8HTbzpyhPOWXRJ7mFtpBFtFx/1SME4Mx+8jU
8m7GngUHynfVMIoGg3ErBxmx3UcdzWtL9TLqR8r0IwYJgKFGYFsMr9m0Rq3kyO79
u5Q1VZLhmdMD1YINutVxoWaKgkir9HvU7MsCjruk/pF2LB4WEx5M7HKAhrOyoAHN
w67wYP7bkyR1qfpn/Tv+4n0MWgMyYueKhmmuXFgmWlrIHGHt0Xs8XTZ4XHkbC/AP
O0UAcLvSGU/hJY5Ar6vmW4n5Kb6tDCNhVZyTZV9yJxGxMx+aELTTNf1j3Oi4VA+T
DZHZodWxsVBD0uxKpA7DFvdVSIsMtx+WIgdC5NvEjEsAEQXXaNv6DAZDO+Dn8eNW
iZWmCNwllIeOGol0FPPW6tzkBcGd2FNTBOAW+IzqOy8r91JnOKvLnLZJKPK/IcRT
AGFHYElU8ozXHFPidJP6/zl1kczUT9sxxo4ev2i2Os/AJ6WX8n2SoJboayv43fDl
4kZs0c758u9alPZCaJlrNOphZsGsz/49MMO+9rH1pZw4tmXc5FHypPFUPOOjRuEx
deUho0mQSn0OT1gB1BTuXB7ewB8wvVift7VqVoylryjvNwDDKQXroKZddKHAlmDw
ZZ/NH2aEwbdYTWpH8O7kh5+PyP9Hg7DHRkmD+ZG8hiJ58kaMHvBLQijiDk5B0T+F
yJ8uYKx080yp9U6pqdJFOz8oTyMur3khxxoyd+w/wm7LPcOXuWzLZq0DqfiUmpPw
FsEbytKx36UB2Y1C+VUMGxA2oSyF5fSCR0ASWh4XqGvJL/h5sawVRlDI1Lt7V7za
YUl3JoTc7ox7Bc0M6x2t8my6D2+gw5kkFKtHrhd5bHEMirA6nS20N6zaUMsEOzcN
uLCBwRNtySCzhNjRawpymiFwD3dXH8FfL5nlyxr0yvYd2dCshvvLPI1bEoLT8oek
+ddTqpja5moI9rvroFgkY/s4uKilzzRF/63dQLj6YniWokm8qE8u3kMhl13yuy7A
UTMOGWP499savppTu7sp/aN6uss8M8Ni7PiDQeld5ccEu+X36e6soQICoM7GGgjr
rcDhV0WZgEUkqQuu9Xe5cpcDSnLNeH+ixWrIgXhSsw87NGTL/6Uq6OWiJC1uNowy
Ldb/sX6i4m+a8r8iYm4AjpWaZHolDydkm7H4PsEoPXRZfcYv01WuavcJL5sZhFqA
dvUuyT+IKJgPvAXpyzgUJlCFC3AkJG+GwnE8higdOSNJyiIfsESA6SHuQxf28jWO
2yuWFKkbYSMmdz+m4emreKovoX3UkMeTbD6TAuUgHycenvynaVaXJN4vknJMZqgA
OJdo9xlvQlfI771POQRx8t7pycik8bZwVftzqinvPVUouKm7+Z0htPoCW0YvvUg2
F/1PU94CdpkENWnv+BmgC8kr/cCOyNPChYXhJejYX8Cvn4WrBPdQb0gccCx13j4H
Zmnrqg4bmGY6BIXf0qO4nmXb+2fG8dimRnpYJYh5bNIxwOL0Ne6JqjfLPUHW0ZaK
9h7HE/1EdkW6yjKzDU3D3ooKY0vKCAUGJVS1Zy+otgzo7JkfeVWksBkpEDsBkCea
eUdhjKbVtVIV8MfMUMfuLnPjexngtS80LIeXhUVoaMTgsHXmT9S2Z+4RMo4bqKn8
WU6t3iGfpPk3q7RnTsQaIeYQQo7Sem90fyHn+LuQEUbVvHh1vJde1ftigJN53YZB
J1tUc6bHqzlPqhQNmlECSy/BtxrouSGSUymtq16Vc6hrWdDSyx8ul5yYoJn8oJvi
ZFavaKtmXx1G0/6lO59bb3GeEjn01s6zBvJN/yXG0CMT/rvDXywIv4bFvyWA70YX
IF4Ik4Y/W3X12/DcoywPAmkv7IveG/2b/AuMQtjJ0Qjq6A/aKVYEg6K64tsuZVyu
L1ISwBpgMYNefJAcY6DxouuvNVOrUe9EuTMX15q4+zlmgSBzHgs+orYSdmjB9Q89
HC35os5zoLC3iyO0nIfE08XkanqazK+sL4sxb/NoA+3fGH0m8i2nfKgUMQz+zX+O
Y5A6iTV5mrcfXnBnePxsqmiLYBMScTinRDcNjWQynVDgRBBjvT3LDcK3h9uwLTt7
qOgVtKN16oR4myjML7FUiBv8EQOhtBO5e5ruxNNDg+/W5ulscWT6UPMKhvNZ6s5L
IjMsBK7QUAIQyCTH9COtPmMwsguUMeuQNGJgS0KKVW54ukmKNZq7sJIS+PnCPjwU
75i0SiKgEBnJauPk46V8Cq5AmIqjUYqetNfFzphcysYDc6KjAdXvcIwRyUpvHJ+K
OYbyD7f6qWjKIrXiIzAI0n8BM1eLMxSWiyr3KLPceQDqrUvj0lan3XBVbdUBpMFt
fgKxkomysVNx2930cLAwBcSphWQXtXBQWd9/C9LbV82bCV+O+SX0vVrRNhtlcXdK
dS1VhtY7erQKsIZticuzqwY5nFVnyXQGDo1POAO5OxfYaU+3xCnzg1goC1+Os0E8
uHOe5O8woVEdjy1jzf2PFMhKhDksRMlxZL9C4pZmUBDxmk9EYjObAHkUL9HaQ9IY
dudhiMf8BbkX8vzQP7zuUAMPkwk0guA4zTQcFUAzKHMGkYym6RODhKzi1DRC170m
hTZuZU9ieayYq9IQyOkHCmfiHOB3m0i8JlgT+urx4m5Xr9o9466/SSxIGY0HRBiu
1rimjDZbCclKnD92v/whuIcldWktt4di0k0cvN/pD0LG/sSSBN/XDuUv6j3d6+/G
6VHDuqQUQRLambJbUT4PoqlApA2hfcwAgJpNdTmh6CmULQn9SX2KUIpMly+ZYC8o
Mt69dC1sMKUyKL+ntPccqLN6mEnGVoccet299L/3mF4HMIbuw2DlidtqbPpG7nKU
F+PGU/RMOiX2QYt/mclde62zpMEMQrdqbLAQcqKYg9JDywhNWYW4qQ+pE4yl0+Hn
GsjSc4JBzdNSIhH2ba6cNYmQyjp2xTd97RwAe9xDQyqqXMtUHPACQtL3XyDu/fqk
wulzntNoMOUDllO7g1Wj7py+/hJ+7kUNerK7zlarrHQ/AyJvP50NultBDuVXBM2C
tfbJX5602vnG7sHTcKFhNu5chxbJKfGjENEhyPGRB3EfEqL8idVJ9bPoC4rX1EL/
3X7X+h60qLpt/EfaO5uu0bil8LE5/4/RYX231M9w+6RF73UITCHfIIWTiTWXXXmx
58iqPe7+Et6G17LWbfaO2DwR1wid8A+kGEnR/xJPBEC3C8Z+kNU1xbECxi2WKyHL
7Dp8xLKEEvK8VseGm5fid3SV3UqJFPCxfr4uWre4t193D6yOAHB4bnjx8WdhI7IA
1ioHIBkeu7xIcIhFsTj19mGA7dvXE/aX/upiDj1Zg3FHtmwP2cRshKuyoaSkllrC
caNJVhjpLouzv9z1OrMQ6Qgnu3lkdiZERjT65U8HbIvrQuDdgW3RBcQj2XAsV/+X
5e8xIk9Ie66Nii7zV+aYg00fghPYfgY2tID0uKqQHiRiciHYKtdXJ13MVW13SefC
EHXcIwjRtz5F6asq+gABeOo0Ky6iVaGRfrNae6IvtMCAnMFmDNUhvm7F2x7LfaO7
8nqXSZvi2GU45Sbsfxe8n+sYqmWA3E6iE9BPYd1YvoCH81HM7r3yzKBoSlZxXC6r
ar3H4slYI/z2WVVhAnkpU9wVxZgsL2Ye4qwNn9HzWi3qW861ITeyapYT4+lnunYO
jArwlXduXb2C5N+AFRHXPko6s1Dy+qO+MCKkEbzIt2b6oBU+Q8tTbnqVhTxIRF/w
MVlIe5vol3H6IZ2X+YxIu+vuaUjtCleLRYw99ArMxT89ZFdqms8ivjj1M1wxXBlX
zOr9c6cdk+Cx2afq4QX2jTXAN9z39zdefp4pGovDSMyXGtgJI95+vdjxWMcjRQ6X
CqkAl2nAo3npzGV2n88k+GefEi46MOen7ZFcZZrz3V7N+zFZ0bVXsyd8LDrSSnOP
UAzGVa0U4oYzKLBZxNxHiK6+EC7xSoyIrhYB/9BJod8enpGilU4Y67CEdakl8kk1
RdthrU0IHy+0HNIWkQHs6KZz9F5cDuSdehHdo51cL0otPqt5G7k/tlUrpig/+B5X
uM2jYRUBH3sHNFRgh9a5aOT1KkyxL4h3RI493wM4pxFmcsnl1tNiJwvAqcl05KD4
3WuLviL7RlMBqgqw7ERb1pUwM+IbvJ8ONOK2spuTMhDYBQm7bhZb2TPiHrdvLPc6
eWnTllw4WG6znWjHve9qLISEGPbxtItNeEkVjOHLooiTZHHCY1+ylmgA873j3PCS
CXMjoLGBx2+vmu4PIfk/NXVvkzgslLx1Djg4x17xALikc0hPc6TGHK1RC3rP0uKG
8duUIC2R265IJ9509A0PnW6idX73Lyuw/YhbDYh7/KijwaknLl7E8+Zm3Tu8+sBA
w54fXKvCQptltpfBnh5vackQDtH2bxTnIOM3YZMS+2QfCEvj9ZhI/3CQqUaPi+pj
Hs/w3VJ923O5vl5wsLG8ULIVMzeX5DHBNTEad1EUxfZB9yqfO9uwtVx2Svsgx5c0
2uyoW3hFwhpF0ud6RC91aiOaBCWiivcJF5JN56eOCwLJ5GL/zT/8MeOrb7QQ00Uu
d+M4pDt4AGnJ8IcHdDu/cJZTtoXhTppVlNaIW7wNfISVMLBOdYjcPpslOW1p1+td
ezX/ue8X6fpevXoU3u8B3Zkv7L5KqwS2zb1QrhmayksfkKE8hMWEYXKMv6b20AOc
l1ZoveJ33D5CZYyq/oaiFNddJsM6D7sJdCMcyHSUqyP/MpCGmQ1Gt43hCeZUdjBP
tmWj53iMjhgXUHAyTZkONCDWQ4XRsHZZxaWJrV2KlU/blDL+rUaweMmh93B/QUeO
izal4vbEJtKnIE6/ppKlQIcnOk04pNUqwPkzvYT0fxjqVgryYsWRuLK3RtYaVTU8
lP9cM7pRCKs6fSVILjc5miKZhbzoTiCmrjyYVa8Q0sxx99isZSyZ46Cpi9sBOV+0
S1C4GyTp7ejx909HfxAVa2ox4r6WVNrV3hEtNju0Frm/4gms97nKIKnmkvDKeNUl
u8nF1EPxvSZCjrAyGUMRwMMSUrqBv1x8TIo66pcTvc3ipt8DhkgPLZDx4mKsOBdD
B/f4IxbFYG8neskS71aNLvB+MS9S8wlqTMLqKq5hmN8UeqE9Cptxvac4k99u2ADn
B/FrNZElP6qWhICujDwpGjsAG+YZR5gRul1bjhyiFus7Q+HSVoe6lLkUJ0gXUZU9
+2DdgyMnqj6n/BbUuAOE5xBgDaoL/iSQaHeSuIj56zS1yY/vU3zHL9cFuHgiHlAa
rjDr592ijkXsKqHGFS3F2qRvMOaMW/r/1v4HLyd6mArp5WgW+uLlUI2uknWt3oAZ
0jpv10Zv36QgjmmxYKhPqKN5dDwRRNJNGt2czZNqZxp+FhAp1y4kxqS0e3MHeV0w
yMxwgVHwvU81s+W8x7DemEdHyV42fS0Z7mCLh95H827scqxWrZ/+zoHnD0s+Fyg/
S2D4b8cHUXhR5YjdOCfHWtaCJ73OclVEWYvu6hjTeheH2ZZj0VgBx5xgYEl/69Fy
nneifUmp1ARAPAMr4RtoHXAjWSBIyW5oePfuMPOr1hhoreoV3F4a/fi25uZRw/HI
NeJiJdaMzB7o9t2ITDdfpAxbgIhJU/Vq88o1m/VzFhe2gwOK9PcFwVVl34zb0Zu0
8ABfKjOr5O5ZkWpRYk3VxzagY/GM7pbfY5SsXbr/is3zaWycswcFSqkTJY1djwoA
Yg31ZHzoNV7bZ4IZsx8EUwQhXNzGC8OwVtBbLsGyF8ZYL/rfPtWLxocFEVrrOGwJ
mojuYGyXtGB18XPwFomUOcPRLhy4+EtG/yeL3UW5OZPyF7Ub8ioi4w2gdVll7Y/0
WE5qC7S73yDBIfaMjySsQUjtn8Jfr1M2xehoh6NFunz38GyvI2HrW5t/DzbUQ+zV
iUJI0Wv/dLL26X3jX0OJQMlyP0mDrKxgJdgk2hGmPbMMYtjk2GMbyOYOcePhQRax
QEYQlWZJqmrqAV1yuyDKJasQMvTiA30h1E3Z5Aa7XK4SBtxC+kZ8Cew7u4Q9AvQl
agn0N7H4q7gkJ1fz/8PzWqiB7wdrNBF4/ADwi9F/VYD66DWY9nxzOmMm7T969rf4
F+PfHIx8V5Uay5qtfij3maKyfQLh3OAY0SUMLlwT91kriCdrusu/QRU3F5pYwhfB
I7PR8AODnmTrOako0Ttq8Uj/tGuClUXcKh3MqU8t7t+W8N3w/+qMxNgoF12nhRg+
PvVDo+mNj3RgfuNeAdYF8pDTjtcSr2YXwgg8JBSx7vlPU2hP2RDUmvm2c1xz+63Y
ueCsYbp7enjEFBKkd5EQ0jJu2vd7LhArrrHgFi2yMC7KmfEWDE/z7EHkK64gTYhL
U7wIrNyVU7bG8USInW4w43gdoFiLGMcMFRLPc6Fgf/F6ktz9mPufb+bFrFTsYGk5
UOr4lemBwhQfipfDNP7hyTv9s7fJ92RlQScx++U2Uvj+E4GdY89CTQGLibUFF4WA
1CSvm9a3sc1k30VIS+EHvzrd791cLgDRo8MMmZhrCIeMAoRlR5HfPOqwWntehibZ
Kj+DEeRG3zebsndGdDMFtX98XhFWo3Ghd6OTtixF6N4QryzHOVzT94MAwPq7Vf+9
8bTnvrrONLBel5GGzz9JqRlzTbN2d/q8Zcv6Ikb7vWcmR+s5dJKhECuars+4aDRF
8b3TzvSSxj2XvtJirdxyyf6gSW25FYTQQdnzNKoJsco9YAsFPHBmWbSLh5sop4qF
f+X+2NJV6xV7IK+IzYfJpxNGHU4etIfrXgTQI7PViP+YKF98MEHzK9lRGq+LWzXN
zs+DsbciENH3xoZFkMytzpASea3uiREsKxkfFXz1+yKrP2ZHqwoKzCEk53MFd0Ng
N/J7Z6msTAI0C4+qFonnC0XgocTJnSpA4VFMVAk3GhFwJVyNOgjOHLsxzeMNUWq4
OBl/dEb+yR11Cri37NHQcxokFhvkLY6k5oziqsaBHUApp6ol5dAqRH6PXfZwuYC5
J6QA2BuCsCF5bveHOYxhrrpFVLcKkpyNxm9ds0xNbxmotd+WPehpR4OZslwy3hyx
MbO1Yt5tRzE/CJe8jdjUPtFr3TmuRHRqSn7+dmKTGvHkTfHsgX/f3rN4RkFU/N7k
b9lekjCM9ZMFqygZb+hLdDmFnQ/9JbGXSiCA6wHg+wGmKd5dXGC2Y5OmUqqzCqFg
Wjka+l/bjwFgUxKfWRSemgQx+Rihlf6k65MHy2Q6NzG7c5oZ8VngKXKjJs85yDQ4
fXZ15IkSFvic9t7EhTF/mKnpwFPMcHt8eJ7KOGkoXHISey57WoEtLzrt/vYXkhIU
RsGFqZX39Yu8DzxZd06CUVxi8kXh3vm38EVXXBHqtA0RooEEjJgYar/Luh6CCTS3
w5Rgnjbfk8I/t/cvKrNT5lfhZSg0g3VD1vYcWmrWMdn5yE61v5vyYtWWVschHYHf
9BKvyffm/kckT1k/ALDKGhTjI71e/dBg8Z2iwemAz4+QNSzGVu2JK01XiRsLFBSe
HsCm4Low4FcO2jjLtKIeAw5+KnxaxB8j+hFf7GmxepavYjAWJj34zTsnRUddL1A+
vfrwttyfYC0PaiTJ7lyjfXLFnvGlBSL0laohxRsADmn0X+a2rv4h32/4fuX233BH
Gd3jBW6Yme0b15P/A+dApN+uHD4w9YQuVHZ9J7M29tHxQAwQP+l4Fk551FF0Z+um
lZa7gAzh73aFnSDyaxqyOCP8Kgc5fdcnJ6VxC6iw0ZoFyUL7hEBbhBF6IdEwP4tN
Ey565141FQW41Wi/eMWvUtmfWUDX7IHq9TdD4PHX/oHt46Fb7qg+h3b/gVVYLP1W
E99IeLlp+fuxDzXOWcPYkzjNzZk+dl065XIU8PAIM4+nXjeqEUrg1HhgJUFHZs8b
hJilAYXgMww/4It08vUs5Rn1enSY10qcY/y3WCJIKJ2l/cLLtYi4CnM4AzBr32Ap
DFC3pXy/Lx44C7LKiUPKpsuwlaFBEbJGWlQs8w3wJk59GFL345IAaNw880TrK3Yd
mlV3EvAgliEqV3iJvtrCXunnQJqz1r9U+CUfzKiMjoYtdaoTZN2OJrfHx+xOQtBr
Je8lE7bjpVn4NnRm4Z0tPcsJIpVQTzfez3+7FdX2483D0ez0C+4kE0CKBKJy5wVt
7Qae57sLjiOvQpxUrZZMy8Of1nWy6p3u4YBKFwfX0aKTrTi1GPXW0i1OJncRdp0E
NDbJz2KvdKj+uXmwzt8CT0tRHDFQ2Tp1SKPn6MdmmOKbxhcx8myh99k7NPHpTkEf
RUp1tEEBv/3IUYlX8kpNi/XAovvYT2b35RPzCO0oQGg5a7eN8fNqeVjPKg86k2aF
ugvjUjC3lNdNX7JiXH9SaMEgUy+d3YWjSsSn/gKuJ+9EtLUTFBa9Hwj1i0w5vgld
KprAqO2xvYOrfybMek5a38RCbhbGTX7GvZAVJfNgv0frkgAVSxdJ5IXxHA7D63aB
NfD2e1bJC0OOqXE8gKDA4+OvdZIYa3uyWSpWaPFAf5fg09lX/7cKFOSS4lD+Kp2m
qfDKxrt2TFe/JO5dk1siZS/DQER3yunustnq5QC5yvPktRNKv8yCB0/EcnjOROq4
0Mklkg5qOvctKWJ8GI9tHLBokOX6X8+QzFA/r4/UIc6oAreMQVTOOlZCCN0LScjh
B8J3I2GxpCK0NnsxzacSnSEFaXxG9uj/FqBTcolI9rW1L51Z0gi61VapJDUlEP60
5zbPoq79G6Zwz4kaE9EZLKlepC4BVoGulsiuopCNaB6OegoUt6DjDYKrzE3WZcxL
YZ7109oAUU3GHpZhdh6XseR5ivrBpF3L934mZrxTSzOjRPt9dqULXwvaEjP+W9AE
qZ069Bh/p7ywueLkd7xeYGOERv+ojDlNajoAp1qZ5ZzrQ4UxNhI35e3ROogENAKC
4qcYw/FDeEYu0Fl/7AqeUWjdkAPP3bOu4tKCY64c1j/tmdqELSKMOPhOmasmhJ4y
OjQ/41Q4/CoUFtC3tyRkMCSgrM7vIDNDcCjwKnr+eokVBsm9WDrfF8jgaS0aZOqF
PAzMfahjCpH1io+wt6aYLpL2lSeoiom8rZdMlb8l9OH3MXxNdhjbTUEI+JhzA98h
98I5JtGoFmllt1ZYAvaw5iqfCXA1Ay7FewuBEAEdF4lpRiIV+8QZCDPQgKwyo0hO
Xk3hEWRYqNAqVUMw4vGKJ8516r7yVTJKO9RxVSX1lhjlXygG/qwYBgTVFTI358Aa
OSdbiO/6gkwfEZIOCxrT4BjExv63Pcj2HS7kizE5J0aFPkIp6IWf+k6tz/IdxANl
x01V6QsaQ2NWfeFEyuU7382QhVzpPcfkePskQ3nhQiT30oIWEPsSTtKjy+/WLIX3
zER7SdatcocQMkneyJG7CWkBiBTn/qcmVutA3WmWHsU7oTs3FUE+Ee9UteohD5+e
kT54+VNtRm/cBSrXT9vRsg1/a4BV1Q4orrBDH1UZa2s7N+gS5lAN4mr5kHmBvEek
TwdaNNuUU5+PJAD7topSc5dbO0WwqmxucY9s0AftkjhcXIbo0ufhC8/qqKgY3t21
hbnDSwf1K/mlG5TsMKSmfvVSuqox+m2zqJqdFI05XMyML2OBtr3nc1ONNvHBZwrQ
lXHIjDbXQ/R8TD7ea08QqZqmdj5LHKIOEwDr6LDRZJLc5uLKhi3+1oUmW45Rsfmi
JTI1lhIEtGuW1uSprkNgGf39SBSj2uDrYykwxgjDjCmaLq6NsUqcClDetLZxtinM
VDITq1NFwvTNkHEueLM952XAS6+Kr0m6pg9ZcSxfHEjgve6BNCNP4d/+e/uIxCeu
53WjghbPg3xGvzWX8FM677dYLx53uU73LWPRiq9gu+JGloo5gDV8WTw+446DeLtQ
frYiMJTC1NUWVgnt9XN8ReE5uvC7Suj/yzuEtpIhh24BJzVzA/Xzoxz/cgrlo0lM
CjbXvGKMdu18D6rPBUdkuzGLX4ABcsNsSwE68+xMzpzH7brPMXs20gKHCcHzMZUE
9hPQDc8MIOQ5LxGn7HBFQDTPX8z1D5GKPy23FL4MyCnOcsRpBVpglsnq5Rx6Oq7k
plwyfvXTlymlx5eSnIzauIXSmPtWUD5ajPHv6CpVDubr4farOMqITHa6LY/l1ada
teYphC911wrBfzGHR7poBtus6DK/CJOkm/ZgTUn6leGoMgPhUOjV4eGoFXqBAk3Y
WTt8CagQ3xe8PPTr8yU3/xNPegi4SByfAsrkPA4XFRnIvAysncBkD235X5JXQzVI
LQZL/e4L2HyoFaBX3td4N12vud98v2nS3bgcj8WA1w23eyGPu9/btAJ5BdWeYKOc
WYP2JvaVC90eADclrg9iYxLyLAj9/J7Bs1oxTK69gotnywz1LoJ6L3E1PD3QslMs
7hQ+NEchHznSsA6eQq49dE3lXHpnFjrKDp/2utiTdevJm15uq10rFDn5EW5WW83e
Sww3QLEo8ocae8Pb83rHAc0DyzI2J1++O9Qtbe/KSJUPm9IEbqeGOdCa/35/MbVT
WkOPPcYnrfVHG7MKF+6tTXEivzzyxaUVTi+7v9Cglcl3ED6YcAh59RdMf5ELpqxa
aetheQLIz8HUEo247xnBTiFPRug2vnFVgKYWdnAHAAEcEOaiBGGZyVPOJZpH29eQ
FfLSC7zyHzYX0tLyYWrE/0nkiHGUGrMW/aqUC6Cn3pC9lp5VkOVqmUFs3tWd5M8m
sRo9BftNElSFZ48rQsFvDvOlyvWfJr7HbkdpNSpfxvfVOabYKtK+GEimtDdPcvLw
KtpfbCuNhw6Tz6pkafxaflrBt9BdPZ2/V88k4BQqVBaZtwLBB+PmXJJJ0Rcqivn4
aNLakObbEvKYki2HouFuWchST5mAD5l8kfrfPRVLvXO7Y3+H5QCvmVjjCL15fwWd
KVg/UXfhDZDvmRPi7H5zjd6yyhKEEMCO8xl4tftKmG0DDO9oSA1cNijj3880MqOW
Wfu5VOXTM1pijxGCfIXxuE3ewOYIk1ybwMk7MbFc6yoiu0HBttSgPKpdlVEQW40J
5mZ2zDuC/jNY11unifU8Ehb0phx0FOZ9EXrCAEe3zTZr2mNESfs21Qwr4bKuEugk
ODIFmnD6kNIj0Glbp9FPhTWtU7Csu83kEixTBRkc8fc2Q4z+N/1ZTSvqcma+SGNX
nsXxBar9mEV0+BMwdexWf1A8qwT6cXoGo5k2ju8AGEZthV20NAIo4Y80VYY5QtQW
3GHTpqRlzRFlCuS2JboGuMd6G2HOW6YYtoTcoR/cAdcizyDT9jgi6CFifqaoohAt
7rC9OG6XftgwV5g1l0kB28KR9MzwZbP3jGpgy6Pfju+qu8eT0iMAVga5NqDa/N11
jVqxMaHRi4rVdUvHlQL968zZ3JXqy6ohoj/Xj8y44K0YalXNdPxJT09ig1Sh9tf/
aYvjwG7txpUJa15l0DfhBQxTrjFI8J2OCO+17i3nkMtLEevtSBCBzF8rUGsJ4g64
p7S4dJIV4Uj8hT3BNod2yRXOniKOTNySb6qWQ1/5imoZ8TZnX5oK7m+IdLD8GeaF
4OVnd/X6wSCPLOaZ9NPHaVqkkihFpT5W5YdchG1LuKyW10HmUojcfnW5sgIVZC9A
v4q0574IgbH7vnBikWOpIYuczSvC4+AGBi5n/iuB7fq3NrLEWFpowPpEhgExW7JW
xYT/3LqovUGkkVohMLtPNVM9pFktT4oBSzC/7iVGhwAcbFM+lvvTjsNc1C/IygC1
MBsDqR0lkIcH8F0Z9Y6jfbnrWyDoBkcu71gdGlStyzTFo+gG8WwT4j2SSN4K4zjf
1goIpge2w7wTsNTBTcGYllgWAgv8lEdQiH1czYy3Nph2KfBhImh1nc0oU6Mz96Z1
VthZwqsRNZguXmlDMkSpCiF32RXbXcDoP+lvYEch78/Bn22HRr6hAF6+3C5pXijp
QHfyQaw/72wTW2MOAjMM7r55un5ElQwLxQQMlcy6RwSGtWLXKCNT/vU89nheBFqY
v0f8kyhQjQ1ORL+Yv9bKnSw6lI42su+e4ZnUtwEpZi/MRdLtKmEEaWghDwbsR9Ji
xEnskiM8OZfWe5KzKfP+Rl/Y1zsSYh3TTfJFuMy7RpF2XCmTViK/6jYHsdcuCbWb
OP/N1Is+Ys2Tlgrq7Vet8UhyAeB1aAVFAgPoa4RrARH/xX5ATHlfb/Q8oM0uPhbN
l/ihS+98VGD4lJfhqT/dAO39D1cv6Ny/1aZAYaXg1mjFW+UpXIztVz9763C/ySrj
Hweg2Kods7y4h7LftybL/GPFO50B+Dmb4VNt9NzK0Nm2NW+i2qmtInZGRPzZzK2b
TS4ndrALOxptWFLjo7uqUnyHvpmNEMC2dy2MsHOeJ879JjdUKCc+N4v3venwdAah
9VToeSZ6RRMOt4k4T79FwNy2HhLbWcKayYnbXfkPfH5ixbwU5ESsPfIcsJE1czlB
26HHKWV8tlEK+HzcBEZ9lie1Qr4+AS6z2zQWH3PNheC2CTzWxmRaW5QNZjV902FJ
pCd5xiikGEB9P5ggAEBPV68LurB0PxSV+yKW1NB0DTt0wlM9xUS9wcLkII87Z0ed
DnnWkD6x/lWTM2iGEFDQWtih2UHNTjunx41yBgN+xXUKFkobW81AMOfIFPqHT9mB
L2TGQO76LGPaWT6tdN8+PhsJzor3Gp+ANHOrQ/mjxFWyRwTzLIL97Ja8I8HCxeFq
lnSjpXnc0T1p11F1KE2sQo10YX72ff5AjLVUzDJFsAgwjfxYiGUZqMpzJRKX98ki
4XrcuUzHK9n+ak0bz+SLbG+tXbthiIe12fMp6IbldAzCtJk4mIs3VnYDzbNwefKI
VkIxR/4H4CtyCBbTB5qdHkzRpA4JGt6xdOPQyjiS92CBqlj1mMN7rUlXNJk5eyvM
VvbUzwhVORzd4jamdPB2zlHPCwLvNbFAgHpJks9n46KNtPzVbYCCraGPW0Ullodt
Hu+hkybh1h+i30rFmFChRpJu9r2XKSVW9Icdk9NeMpF3vLybPPou/Y0JcL6cYhtu
0roBhLGhUdTzTrU1L/w9nQYB1KY7e8Ki7PZUuQR0wwsDJqC4pCLzpNh0SyZNlLx/
webbYn+funsWOm0HVNz7MumX2GqTeuYm5l5nL+FmVVCJxPB29Z28A2lRwBCpHitL
/+iZmZ3LfPpHoAnikvbg+IquWId/rFjN0bCmVnCGPtlPsgqcyz+eMizOwx5PcMT4
XEiEkgfazyCDUjfIYZHRytD3EnMMU3e7hQ9690olc9JRdC4NEh/JJktMoXj9MRdk
UgfD+0HciKNyTQYD1OGMrHQRC1rUNBUmPll5Ygf7hItjlCjxZkGgxXIMogsQI7aP
2KzNJrCbE9zyhvqUFUHophyOhMGcdxyhsra45lxl7CxwpRg+eKRfO4T/pzByyJSU
ihHAONB6n/gjZ5toFsG+4GfujtZpow+IGl3akIOKUv1AVcXf2LmDXtJWxPRTHzzE
/m/Bjp4+GZ1tg4H+MdfbK/VyutP2tLsOmLjVpfTYXdDXsb2efTqD87jGa/WVxa04
0Njj5SspepYBdmCKu2ear3YZNYRYrS/JbIt9puci1iOkTxEyiQVzYCPhTwl9cjND
FYBsF5Yn8mxMUesRejRbclQjwPgmMAXCNsJAM0oF0MyR3dzFvHSmmjbw8vz6H1wI
Svuuqroq0PdK6LpDkwZFb1Pla/tzw+Qkk1kmLEh9MFt+8zRtJm0jGBXCinrXrPT0
BRi/G5ULlWwh8eKXgw0LcppzWP/QJ8obifjZkker98u2+OFO6NtXursmficfuMjm
Hiqwe+/O5YAmGHnYo6X220/MUU2dgqUSRL7TTHqu718NAH7S+zoHi6Q3eYBSaPoL
Vml9m1jH3CkeT/+pFvm0ZQRD0eP2aqn/VFdpDNBhzdnZEbh7GDoGOMq1PQ274FAk
NjOWq1I187ZbrB4j5+DrJDlN2O6+x29t1ozXUmgxa6q3odDBjZ29POlGcUnfriUu
CR817d3DMnCYZKZ6zJjhnjw89C5XdKW6/uAJ8oP0ZQTuBadKQ+wQZBYrZx/8xip9
QOgJWQQzxA48wnUb4Is/dKwVM+Bz/9Zs11xg9eGEDHVpoFdpBBEEtax5bwnXDNtP
i7kqbC6vikOlT9T0Xz+nBJFg8sTQ/LWgLkmdo+E0AGVMt8Lx1oxbiJCWOyzGsYV3
AoJrpRJeTIgGfo4icFkR8+7HxqyRIeGb4sUT24SoKbdXFTEQoDvibpaQDPKSztik
T0bxmlXkV8M7Nh/JDH5fufxq4covGCvH03BPVjcCnvIw9j0am/l1+moVqtCykH6m
i3JoWDUiXI33QwIyD5SDldKEeZ5bmIGJEdnoSDiH69kAI2nSfUi06gveyYkN9ORF
m+0GAeX5fCusYrOE4aik9jsjqKvF3YJYUayQ/mOU67hDVHC9v6LVwSHhwFBULzJn
2WP+ggl2hF1Co6wMSO3M2ZpktjJHhEa/SOyYIVbtzMZeOOt6koEmMvopuWk/4Pge
nZAv+uWfXfTPUkRh0AObzE/YHXdsIkhuPgTFBwyUj0sdd0/27r1OoEikMI7TnoZ+
bxVRqfZo6GyazJCiwjThG0v6C0TwPNPSL1iN1Sau/ejZUmp0w5ykBUw4bB9uZOXn
ZE1drii64Hfle9gWh8Sgh6+uuAcy1fMKFvW/HiAtnEGM3fExZ9CwrlZ/dEFGcUYF
SIl9RlSaAqNP1TUDQpeFCSRV6iU8rhopl7uam4rEQQ5/wk0fptkNTIdeV8k35V6E
L/7N83UPx4FiTHPF8bspLn4+CfOtdAmErY8V5RXqlyAQ4YCZ/CqVPYItOtoE5aJz
THPjBWYmhu+x8mwWWhc3J3qAYEuHjnIx5r5S/cfgNxxvEVrV372XgLPJXYJQ2+3A
cY5flmHIyxM3+g7+xabr8h+r4dJxuupWZ/P5iTTbbY/B8IAx3i3c8WuNxfnliMpQ
ATjZeFrU+dxMPSMpVZip09oszJ0nJXjH1PidxrDeeU4eURu3X5NqGZh8iqbvazGa
4OSUsGQSo+yTIHgiGxQW9ZXdkBQB13ZXXOiUl0nATiPLIorZKDrZG9RVlefBzP0A
fejjL+qjSqSMX23JKPhGl6UwOwWfs0s4TKIyIBuA6tyDjdVNE9bNrGEFKJ0Eccfs
5LLMaJyUYWmBry0yDkhSBRdKUmDlTFnS7DSdnTsFKA6TwYXkm9Tce4M8t4QA1+WI
RvQ3V4n0pplZW908KbUi1LuQsvYX4V7C269i8r8PkhuQHY8dQhUpRWqEWq1JLFzc
b50FuRKkOzV32JQ584ftLorXF1MMPbzMXe4e0FgJ0aWX+PMP1IZxyEfdYHJsxjc2
MWzp6Uy60UZabYLI1EmmTaaOwsUnZLCFnWkg+x2Li4bXRrboXOTHeaUBunuCzQN1
+hEe4T7a6BSwtErl7gZniruEMfpcT4ABHQAdWBf33KsJ2hXNPRvwnOQFHZL8L4qU
Wdl1I5/7DezwncLQs1QS5j6zlA3K7QkJyworAzfOvLvTvIGv5Em+BR7R75CqUxRW
4gPSVZLo0KF3v2/Su8g2Pj0vmdCsqcM59gV0/AfUIDQ1WhG8urHJXO0dDU8ahwww
mBGKq6qJ7eJRkNf17Xkjo7Kg1O8G8DcSO6tr7DVrS5IRea2zDl8U9FAVbwMRhWQg
QWrXNs4XHk0RZShw2pkx9WvFtwnEo0vRJN34YBbzilymgkBW5YsYR7ZOIR+3IskE
nCi9NdDAC0R8/KzDbal+D2eN16YbiruH/Mr5TSnUEmfXNmAfeCkgOSSm/C/IvgFU
EtD4qBpS8EYyaMPntIbqaPCVNn2Ad+SuWJ0Bn8GDOPfnbz1i2/0nlHFnZYYeXf9U
2nVw26Mfxr0jwJjam2x4FWeu3QQegUUGxnt6vNIQJ+ZEjzvR2Q9+DbPKzYOFlkEQ
WbMHdpaph92ut00LojB4bUKtABRrYZm699cvIuSIyS+gfGhO40qiCYgAPvMSl9TC
GeDU37eb9gV8a/1yJMO/v0ESy1Ftw9YZ4fxfbqzbTBOrZDMBpmfzjSwsYjSHW0jT
j2K+vQVZp+iWRC1MPF6ddWNPoxZ9Yl/zz72giu3eDj9iv7tmyE7aorEiq8AgWABW
vfhfujU9qekGPG9sxUvqlS7kmemW37SGQWJhTj9x4bUYi7jLB8A2/tOLGDiUTOKO
8P1QFTV3Pe3kg2ylUANA/Bi5TvpNtA3HaP0DPENimWBO5cliQzRvm8kbbmkO9D3z
7zdQ9wf+djcqBM2b5u+HCV8HAQndwWFkBOzoYHlNfZDdX1TcnO5GPiJIUjWvvB7i
fKhqxc18TC3IjEDUzDeWze1VhsPs1UhwOvkNFwK40kOj/81TUlAeGxVLm2bSsKcv
0aN73utwR8dqOocn8rQqZZnUPxoiWlgGJKceTeC6IcR4nTy1IbdZsELSYAxhH89h
RTy+z5/RavVnF8kkC3m5/7WqMC5/bWEW3mxISF7nkohxZ/xR1YMDBInFyn0DVM+b
4KG0LtNLiDCWL4Pe/1nAjA7imAyNm0ypZhBo3ipoUQv3Ts8OYKPoy/obtV6lkhz0
dD4cEewhxQ9id0qmVu9Zu+Pc7+Os5LNXMA/nwfbEUdwuKCZEWWt3hbjfXxJFlvNt
KoAx9x6JqyiUlFEUXP16Z40FghXQjgHBNAWrI8FPc3ff0Wtdky8wH45Lz20/RuKJ
3Si1ejyEOtqDFtF54SCJbnrgQ1Kvfc7qu0seSnXr16BlaKJjHHcAlAKuBOWuEFat
U1cCk5zYlASnvx5Vr9r2n2t39Pe0YhLk3oXXhn7tnRcLdak5s7Wyg8YV/LpWOAyz
ETHVEX9kRt3HM2kOm14N8badGOAkG6f0nPfnY0OJZPUVosAY54aIVjY0++/Z8Whj
evXU53lktj54vM+FqBo/GXzwTgg3r51yrpMhZII9b7PVzY6/6mrPYJkoP50onDka
JwcGCpMDMX1FloNqvIlhQnlU6kpuRVChtnnPvKWQuR+AVt2LGEU6CBIlaOwmhsZv
YGrXmAHctecp/Pr2t7DCpDfRcf82tUb0DiOIRF8yD8CIQnsdUbBMYS2dtlvJk6b/
O+M19/HxA4iuTYUiR1rzZ2NORXuxO7ynzNaLhy+Qensme2d7RXxswNllEyMH1F/h
HaSHUXM/0EDkscsQRd9UvhPfjPZRyPtEyJrY8byL8/gBHAZ0U2+qlBe6brow/BCp
f3nvnJxsOwQujcMyEAWCQ1ZzGO0o7RtR7N+LZXjwORP/itbbDsf9JQYvvlYb3yDq
6viTXhom20se+KDEDhb/cdFJGi8xWuzL7BbXjpzf7EeqXY7pXXalmEpfMVEmhcsq
XghwX+0V2xEAW9exAnDjmoAeHT3+1BIyC0ri/K2N5SCS3ud/dSkKX13PjohS5K8X
ZgsjmO6XS1y7mPiv3UdvXmpLgSgR/CWsRlGVYZ2zVeRMyUZhw42PIhTeBogU6IKY
Jb50Vg2i1Fn3j1QGK7htioHDxjTVQ0FcSiIy8zvnZLoA8/PQlpxTBXSmFcvx8LRb
8hvU+om8xgCcvQXcHFonHfaJrf1SSCDV8J5cluI/Vh86i21PkQkigDJwU/WuI1da
T8X4mHHaHNLfZEElSkYWtuoL/En6d3UEjtlbSFvmNOKIYhhUnCh5ISuj5FbSKKPe
uYnBmFqe8FXyqWId6nM4RIMqhl916dSTo5ceTbyApPwi4LNGkleHCFsinQ08LMSi
dY7ney5uaob0mQBD7Pr6G0BJvgQpaNCmNBIziRakkRcfsBuKNaFAt96b6TpBk4/z
gePR4gyDPvEUulfhEGd3z4sR9qWqBION8AI1R8f1nmLruvKpVnvU/XDBZmMsgjSz
nEPv+Dh3VnT/kK7LhmwTlVe/UKSzLuYTwx+bNgXO4AGiUmFnEe/sH+HuyTjfU5z5
s8QkJVAFQ5J867EOLgBz1raD1TZiOaF4ZmKDAt48r5K9txq4TNRTtHbxlh8qJ4xX
0zMuC9P8PeWN47eIFAEN7jh/IHFi6jEUSJYNP0jPldTvtZQ/GD4oRin57O9v5Gu7
d75s15ASAAoY7nouEIb50/VbNym3vgYtvEYCOWt/ZYBTjUo0vqZxpXKChPJHvPWP
1DVVPGsU/q6IYiVoIz4eGHfudhK4YZwuRirvOBW3eQI9lE74SRUZcIIi1goGOYx6
Q+8ekfjvjqnO78XA3uVMBYsN4ff0huyTgSEqVgN/hGTU52EG+OphYOLff51H+QoC
NV2RhHPHhLwkCw9fE4yY9319qhnp2YqjVsdtV8OEYUNg4EVO/6ShiitCyzqgtNUa
D8jrKdriMooLOk+okO+AiH/vL3FcU0gK8PyJR5PmIGv4mD0y5rPuHGAeRlKn+Jei
CeznueCtgtmIwhn8UwrgmS1ssNUxeVdab+GwB4IvIRCqvTaCm/4IdZ592p8zXAMN
gqKuq8HJayNO58n8xzWZzEXpwM/BJAmeBtoAEQLNOXNjWhL8e7ALxuGiRR2HKCY1
4LkCtdJ59xkVFv7yZTY71ZFs8Z+0csapyjB2j7JcBLE2lVYxuaZEmWlcMFPt28SR
e4H9hOIOCO6zFH38fEDLyJx+ugyaaTGEPYboQ8URRToxgIe//lIv/3isvODQuzHf
w26JJm6xE4t5eCDlKDMRrkZ1aCbZ0cW8jVdC7bKrhZohjUJdEHZX68erwtxkl1vk
3eHzRN+x8Z6o1Z5JSCEXecDt3S4m+0MXgkDy1ju5WVJLf4OqdhIldIsUbFH8yBx4
GhtZ3TtYfXf7ngeB4Iz6srb/XzjmeHumyN7sF16B3+qACgPNwh0hYiDy4mANZRm7
/UPGCXJ1gGtjmNk5V15HlUwnNsfB0GKXmqwwNPn4lsoCQi+v5ZTiRVrSmeVLQzpt
HMJ1BfxaVi7j10NGXwYIhVnNSA9gC8rQOKFKBA36WwPN7BotlYvilYRzBt5KlO2B
y4KckMxmoNiMTlcgtrpOt7wsZSGz4Q/JDS5SOw4XL3XRD1MXdZMqqd0yJ3TInw/i
CyWZAWmGh6laOm+dBIJHH1aQ4GNisCThYpTMnlUrgeVJROZqJS1eMhFVTpmh8K4w
3vCtTQ/wSfjhBSh7wWnQoEKkf0SvuhlJSkxnkKa3gmElKzp9AvZpTm2lbzMeMBsT
NgDTa5/6xAvj2oNz8bF+Z1wURhrH535I7lc/Rx3VkUbAv//67A1+heu64alE9rxJ
enoEUwU7OINPhwuNExJ0/dSuTUOTaRjyplJaz+6eNCnA5aayiwBxJTEaaOzIP/KP
rrlZPfVpMVoJ3qw2gw8AtrHM0hqWow2MlRLTsEjL2/ks1C8t3QFwktDrwi7cF83J
X9BylkANX99U0oCFO8WO+X/1/T/Sl9ZBajUX+0gaGdq2oJRdZMOgsCS6erFiNKQk
/7XaRcE56dJgTKiIDa/0WV4DX0rbuGxvMHXhIsnQBuAk3CoLb2yQx9ufFXCpA5rt
DyHNY2QyrEJURojWh7PegdHVB9NY+ae0pxt69poCtS2tFdbO08efZSxBzFGPJCp7
RLGHeSOuk4IO/AhOKQnbuh7a0Ea0moQ4dDuo5iTkCNhY+SWeF4Rvt0FDJcigPcvP
KHeXaYOdUUrjUbmDO6Z4Ji8dGhybKI5NeLxk9g7RDhmaLY67siH4wUlmCejoanct
LInM8XJqyybMN3omECpjRvgwz2+Jjp8kT/Gb+buUIygWlSVAn+32xUImrFc2Hwae
h2YjiZFpPDeEVHwtrVddetfH4YV5SjwD1QYRk8scFI5ePkvwcm+G6mfw60lwclYD
Y7ry2in2TdO1BQf4EIp2jxxvWqyTqiX76K+KNMJM62PqQt7BXdfQvkiDGGuOPBUP
Eg6lx4UecflXWcYgt6L7DWGxvTyu2b2uPgxD+cEQVcX20vkKS9DWpWnel68UnS/p
StqzTB00b7JQJ72mpD94dM4qZyGSyeZxbZ4hST95xPM1OSVkFEfdQDG10wBqfnHZ
xJ/bYJt3YIf3ulJHTN5bxfPZsFD14uisSCqT/p7Zxou2q6WfOq2/5CiPYeq8E1Eu
FP3A19chLC3yOOzo/cns+ehHpkEnTXw2pzbZ7HwKjaMf+xV202CuM9ag9XSFdkzR
UT5n+6+WqdFVgoudEv1Mk0b0ytWq2OMjWcG2hdkxE7e8EI/KkLfsbEnrv9Q25g6G
BK4/Kw0jT1I7+7DAbPld7zp7ULlbWsa/JrogeifnflX9qzvrSU3K4Uh7BLgUx7J+
bXHKXv568352KXfyKNsQmB9y1/xmm8lcW2rLOOUqdcaos1m1L05AQOLScNk4fBjp
IqM6qArpzli8cs2/lkSL3uYifmgJlD6OMZrVXm/324pa+WCH1R9+8H+EvPlrifdy
rMqwnmQTmC2qBOZpfXkxkAfkmLw2Xl71PhWgnjnYwEj/GkY3u5DEWEwDl9oPJl5U
Ah5DBootGvWPuB97Q8qRs0JILrx+7+q74s4Gyf2QSzVPD0+EvINtKszUBA7NH+4n
j9kUbQcDpHQHtbIFmKqyvZ3jDc9W6fkNHnSnh8tzJ55TLK0rLTFmO6yH1kZVwD8k
QlCEW+GA6Y7tzw7oRDv8we4Z+zQsN08QQNvAlP/1b4DtRNwUsNqyGHZrqMp1iyLu
QIKmPSFzDOt/BoSdXqeEWem1Kns1L+fVH7BUc/Xc3AiICRdoFmGZCIJn+H9iMgEX
uD3lXyPwVyrK/eW4bvdwTILN9FdjYFIC+UgjzXe0O5h2anrhH6ghjjiBiInIcWP9
LPGrquSgAR0ORpavGzRHw30dYTKw/WECgDC3KAAqmCRqSnEKg+52q4IgOwSaKv7l
FWk3vtjnexCVoErUDOMc2nlaPB+3YHG9CXaCSRdgI+i22iPwv/cssyWH99Z9HQOE
op/zVz0MPuiOnM2FXBpGuPW2NnkTOCJ+z7uc70TU+Q7ppFJPiPzL7lYPBMqVmHkE
gUZ1Ntk/HffeYvZkBJP/ywtRcvy0uC7gLEVVw/hbIjcLhPQDxltKfe+kZOM6QQmE
ekPg+JTXKEDGmCrLOnH2F94AGXVmVxnKwTmBSY7NGARNV/9F/99P/xqGYafFS2S+
y5z2HdqYvVVMaWtxaDHHDJVvqJSp2tvcqKflfnmo8Gk9XgfNw9Y3dP47Qf/KQ9gf
12zMKwSyqX1wDsqSm/7iGfWpyrjf8FTgiS8KU21QnqMUpwuDzna0vYI6epaoGuqt
uc0BIzmW4ZaDPIMKJ5d/Z+o4+4fBlTKF1On6h3HcOkGtI0Vj8jSLeOF66LbkXf1e
gGzrSHw44uyqgiDFyQZtZLkoeirBqTc7MjLIeQYtI7DVysw/6J4miv1EYgfLK922
LHEO6ruvJQqffG/miTjv02DbMKNxk+ZPbs8qOLiEoui0yG2VUTK9spLLlRS6xSFb
BXdU0Tf84olfmxu9jpB5bpR3FiPP7jUcGPcamv6nLLk2srxZS/SbfydVi5ziVej8
qLKLPGid7ORPHDIExlDO7GNiU6o5yM3Aq+4NC4sxMNml5V70sw0q+IP7c1h1qStS
7W/sCgO6PjHg60deJQd8upqCfacRnQkulnZocz41ToKxyYTpebsKnWC63RbPedfT
5sL7ZzRJv3pet6ShFXuE2A9TKBEpglsBvOGDhZgW4ZmoxN/DhPQ8c5KlBFDlUiBq
zGkNrERHto7U4FYdT4UmYMY3gitHBBRP2FSrGEWAYJU906Ak0gDk43kWXNo/spgK
LDQ07BLDSPTPAow4T+nSHGtTYcULJEWp5lAiFxKZlDGvtvDI4nxsg2NnkeZemXYV
GMjbYXn4nw6fbWkNingYkAQGo6+/xZFvoaMaQ/Due4qo0So0GlpsFkEnlkZYw3xm
JFq7aDTPQ6znVUU0xEnx2qHODGauasYNy1ZAfIIUFRwfJOwi4WaLNV2fmf/YbrC5
RdhI06Z92zRjAvtOY6bNoCw4m6xo+eWL6fS2Msi79mnXshNYUQPaPZVolSHOuKa0
fHwUSwZnz+wMKQsgZTOaCiyD1SBLk1RX9O76RxO2qWOEE/KkFMFuikXq7m1q1JGk
P2E7B48ptgDbxGGyQz9lXSBlM13olHFrHb8NcQ5rqlmGcxsBrtYAnvi0vmZkaeDs
RkGZy1xU/zMBcizpwB5XfXx3RYloT3/GljZNlARYV/6pbQft9XOQrIDIrpghK5L5
+E2ahJYZu9OuFfZTEcYCuYOdB+CAlg/To/dA/O6De+gNsenmoSzQ8wOZCpq6dbeV
jEq2fK6L7KOB8RGMDv8o3M9A8fjlzo/Y2HBbxuf8yFWz4hT75Pzjf4gXJhMvMPvo
BZlQCJXyoYGb2M58IFVL/82Et68XgE7Ro93yyNZBtyNjf7Fyd+5va+WD52RdOHFK
7XMmnFRUSHP+mq6FulGQLnKWO/gUgUd9/RlrtysURpGb7fzGLFdzNyinxQc51dZJ
Cat9ozlAme+bSXfnR6ArwevoKAut2Y5FDcFiOWkW17Bu+I/+0HGOkgSHX2GmEjKb
M7fj8nZTKEreAyetWR9ynhwOCtVvhKSfOPdrfVUGLc0/aPRkjZ2nhgapbBhPN81u
jT1L04xgORlmc/cjj+eAMMok3ZtOmFSSB+z503C4nLYJqMJ7XO8P/9du0fLASnNs
yV91TdfH0iEKUZTNBhJ1zuznyMtBJtCNKcuGRqnfe0EPYA2dXMPwRhe3sz0Ge+Rp
fzQS8pvBPeCakTeEQRfbJx/J3bjAUXnIzaF5ZOf9tORMZvAwKEYc4Ow2uI3ObJon
+vXB+HGoguIob0+ZBWV+lfAgqinNacDTaFjA55Ix5DK9XK6TUgSO641f7cRlyV5W
coNZkH1zUzzWOAYOSaaX1WxGDZFgTK372ZF9qvFiaAz2ZOcbtDi3uwGvbesEDRNr
PXvfxlbYNNNZn8DI7ff+TbucmX8GJTK3OWqVoYOhie60B/PsEFUgm9pr0uvOf4Nz
ZVmpa4Vk9ds7GEUyTukW1pS5yeVB0nV3Dku8+hisw6Oye2n3xsUMkZF3V2439U9C
Q0QGQ/GvE9MEln7aDCu1s0L63wsVTWH8CiaZqCdqXEf6nDE2vhdAbZ5jvcSR+9tY
zTUShRTQobdRCxJFbLsQs+I28Pti27o4//JU4SaRAKr0/i1Bz6IRm/zqqIGRY804
LThJfkCDNFiON7M/3GrCrtppVIgcKuymV9Lte6GeWdge0ENG9rQAlFSSuWVPI7D1
FLIXiv/BYCLogq7S5BGG7VOoEf6nnxgqoxIPFaAbRoel2BzJuFcnLSw5TZknAL2d
J37hdc+X3CQGaYCy/3dTIZ/20BCyKy2bAiXGl7RleYI7As7ia5usrVgoVAdNk0Hr
RyDYv6S/evkVKR0MwRpDosqgTUACDnDcWI7VXNm27SfZ/W2MJBsqS8gv5TyBZxSI
71FZlGbi7/yLfsdrltHan9g51qjxBvjCK1QZOgrz8tBTeVd+H9Ukss2eD7r/X07c
E06UivSC0gxAL/foHWRb4DkVWG9AnfZB4malqyA6yFsD7lyfuKaG6Zw0KN3qbv88
hUWlw2Gwiosd9c/fx12GxbJimApQEhSgvqi8R1bs+2hXe8UQtLOWP86e9mrn7QKq
oYsLwjfDPx5MSn1dmcANuh7tOXT0HvywKRP84zQKlDPgUhZEjNG5xScgyorEnXKJ
I4do6mwt5jUraHbsfBRoPxZaSG51iM3l5pBPjUVTKDIN8XTpwr8utOywX/YyUTNh
2zBt7nO9KwMFb3gm3BbyqY05da9Y/qZ9rKL4J9DO6h1LaRNj1rlA+iFZG0baSrAy
FHMGZOtg4SnUnLNrOOMt4aNdcKjqH3Gm3tuipptaUjBRqsaiS3gduxks6FnoLc7H
rl7U9WFdoebZBjyDCfD4AsUunpVDCxmuM1udoVdQTA2Cdt6hgYQhE2D3p812u/Wr
xHPI9l11D5exaEU8QnNB0pYGGHsQDIAcWf3p3CbQ+3g/lqnBT84Mr+Ez0t4+4IA9
6V6JxRkeLbWvNv5fYssYyiD1bCMbGGqhzZT9oHWCz2F22Grt+x6ZIK4l29yBMDqw
noe/0TlCbV9iQVX2pkPh4ZxTz0StNaJMBYAFWGdJIU1fIr4t10LAs8V5grmmGZxk
8vR+XYgV1JFGXYYXB4CsinbbMvI67UxqndRnt0ia/3xe0xfm9cGnH2fVa5nczOMw
8pHmXupDQIHDIu+Fl6BVO4zxXmZA1n0OAO97FWG2ocKkYiO/DMMDIbHbfiFePmr2
JkDELvXCIMfCcOwjprJGBv8Y3g5rf0FEWvSGU+mVOCkwHVunRNehzlpiSEQeBzXg
NMzqSTIawHR+zSRdT3QxtcbBqr450E4z1sG6/70cKxDLdBvblC7uhkkOdEHu0ri3
OsGJzje+65yTVh3yA5+mpU+9wnjETvoAvPO9hhGoLAoR/ApSAlwsxmILxkyUsAGJ
n8u0d6jy4D8ky4qm2UK/SggBKf+j7syVFlDmuIyRPG/iYMn/y0uaepn/Ehvw4G/I
/Os1F8lOG/ajbJLixCBSgn4bdqMce5O2vFHxSfLcsVVl5hUBpGbHc0xL9t7SXdi7
1+TT6PdNluquD6pU/jrymqTCShi7MmLAyi2OasoxFY0X3I+Nq6FJhqi8MZdtz9f4
4GTbPNp5FtOneJ1CHvXVQCn+G72Yt0gHCkm42yWutq0uxG9fGCWSb27d80dfA8cf
iDRG/ThEP8oNPemIjh5kuk3N+MB5jsxV8dh1f3xym79cbUO/QDJINkmvMR0cO2d/
WIcXIbcbFwWldVB6bqiX0QZZjWzZiRGy52I0Y5ePaeFhNwjJfQnNJCb+w0EiU3t2
sME9CQdDoirmHU9LcgBhIbsSgdyGVRxj3vAlNXVZRzRNLpJ6GhiI8NCzm2U4ImXR
1nH2I+30kK524zi11C0aXfGDr5Im12mLHbZ6vW7Zd5f8o7ynU8iRuxYcCMMCxljt
jgb2P0x4lFTSRp1bS3p3Mzl6eg4BNlbWNAmSAERDe2X99TyoHwPmC5wLeRqq2CTn
vVM9GoxLG6ykrhmYg6J2MZGQIhpSC16AL9C1aDJkRskRCF/wlOOJJ0deQTxmhcln
aPmtd3vE9kpaVDwK9OntczvHDU386T3qw5/zbP/qT7oO9Ts9mwPgPQTZb9HTsNWF
sTdP8CUzN86v7lw1+pvM3C/xqRQ5AnnKdoyi2H3++03FwGaWq2r8AJ8SLgPl2ar1
ronloM55K16cOeVdFBP4kONsbYFk1QQ/Wkhh7UnxDPfdHVwacToWtshukij84uSi
nw6GOXkdAtf0Fk82EDdic42K0L6K509+3HQRhVnmsu7pS2WRKDMCbXTeyRdfXjP/
BCFj/W6NV8QDXrc14qKVITalK56inDZc99QcksLvwC5IzdfpVycAiV0hh1p8Jd0T
rpp9mZ/DqLmL11gdujx+rh3SKCLi2yRjlyyhDSbRAxOWVHZPQQZSuPF/LnpH2TUP
gDFaFcvC2gn1GIkK0hMZmfq/Z9oaIZvj+KcdtVkCojyzHrxt/2xM48RNrQT4z/cu
hNicJwPg5+qF0ipjuo1hKZ3kd4P+9/8DGxL4fcn7iYRIhkl6HbZtqdD67PV+Sy0v
FcojCJb5uamd6Vb+/nVnondTw+lDw+scEIRjeANwOLsdxpai6uhVlgLvLCRrhEEP
lmNhIJNentMYy/pzhTJR//XeQcrQ4gpv0qtJA/uelq6wT2o3F8f7V9XOURwuMsCN
AWSL0zTpQE16ECJUFT+7Bs7e4M5/pRaKbMWL7ow6PGAZ0arZyXwZwxi9cpzxElr4
H6do4NdZkv123n8TJ6hYvY2RhYx61p8gwUm2huaVCDgAfYF/KE/cSVbjrt2HzGr2
M6AeDhFfdlwu4jhl/syn3w+q1NzcnyiSiyIBNe/aTh/WgyWYyRyYYLJGrLs6Gnex
SPNotnc98b6gbSX0pW7nDWUJF8pi3Jr9g51Ktnsfzr3jMOsCuqy9Gb5X44vZZXZu
8rJHRBY9g/NHLsAghlmHOQCh3R/UAiDhetq55K1HdWI24IG7hKX6G/AntjS98rV4
4mae6QNAlX6czq4XG0FFia2pMGJGmm63/4RH+fEYd9AgFvSK4mHKnmTOe0QksXu7
1sM11eYARu6FNZWkV2frlOQnNI5SBxEQ2ANIEgepyJGYZj3baISmM1QjAQsoKjhz
XnZ6Yun8Z0JuOIlDJQFxyvVAQM31iHQKznI32CkcyMhxz2iouIqql1uMXWnlKPDH
tKgAabAxiQnjNBmmpOoGHisCWZqJAklTO33GWAv5UMIFpSrFgU74cMNdxcfQYHqF
0BxLUwsPyCt3ex9L2BmgZmu4Rx/bzqqaF1aurhWZEyBLXCN2owpomkjpI58wT5XP
5RQxBV3eJZZ9vdjEWIYScHb9mzn7/h4darfPFUHsrefs0TzwvLsySekvN6ldiGzh
ogVF3mU1PFy5d58AI0SY8v0Klnp/wRSUvlVB2XWjf7BA+owG5tJfUK8fqNYem1wa
CCQ5hgo88hRIjr8MIUW6AMqmUZq9h80OAkzR4faVFjZa+lF5obBAMn9AsfH/4VoA
0yZWlZd5+sAtx0TU8Hx7zigzevvbDjaXXMpPMxtRXPujUf/yrprNqX0z7Buxka88
6ojJoORvaVbkO6JWFt7LSIIvmVbaAYCl5m9NBrYfAoFK7/PcDcuPSF2CEFyTHh3g
33FF3Rt/pMCkf7bEarIKk9sKyQ08QZkTY9/rC7ApDM1G7KRgbehQ/Y1bk8ta+N1H
TZBuULG9qrcmQ1Oyu1lMn6ixVVTNM6Yb/I2QeHbM38RaU5dbL2VMI3cso6vUNXwt
5u26lbU+GR65cTrXQ6apDrcRyvK08cHLFrJWHA3FRXWgpVjo8xLTytK9XykoD9jN
Bd2uqB843pvNoEFb+eJZ7crle8xFpY471dsK4C6DWWJpOO92wC3zJ4LgX3UGfI3X
9eiJw3J7DExK4r03foImut7b7FiMEsfFXToIP2Gz20hQt0+1fIUXvuS66QLH2nkm
62TT15h2/zTMM6Gd57aoaTZYOikkfmrNyz4LwWiLZvDohU0Ec3GvXk6l0guM2xgp
B45NPcg3No4ypC6YMLLFqsLTHGli4kXnzbTHK1uM06EjXj/8FOrviS6bMgXaed3u
tH/xmw7PE/p+ajxB9Xt/dhixq2KtiEQHXVQ8bz+WmsNkWmBE5IucXyJ1kLzFvn6S
CE3qxEcT12SAcfZPQExx8zoqRhjX4lVG/vTX9VK7pK9lVENxupkYopBGSzrZKQ88
PS/Lh8hXBobC6CzaHY0dxSbLzwaD0NxP5SEEdu3NA+8s4r9QdeHePgaUDnZajAu3
S9hvhd5DolVUpNSvB28dalm43ZYdD4OYyeDumenKexd4HRYlYMn9PICew/7eaHFD
58CroMPRpRVEO1AOzEop+Br/+CW/+3R3/16OYw6wUyE4Nf7nygXkd531Jjig2RAs
24aF0HIHjqZL7Md8O/8vnkzNgsg51DmfFIW8unsQrCwxjigb9V3kwsFkqiQPtLPs
JZ17c27dJaViEFxIp9AhGiebEXY6AY0OLvfsiIjkuIgm9t3PGnosBZbbaWtA8nw4
bNSWUMKAxI8yvTmEGJ2Z/xV2MSM0OMXB4l1CTJ9YNLGsPwb56FBFTg/L4ZEKjqVL
C4n+JaJ/XoURCNmQ/Bv5OaeEFWRVYPUxdO+m7809zokMQJ/VQN0mZx0FyekKQDem
Da9WDCIfBoxNAm7VbwGl15Dr7mgsOn9A7EdBSQdRNVULs0K83qwhia2DE8kR+uDC
PBBdj+Fqhrciy348piPyMijBGd7w4fx/82fsdxba12NJOzS3fEK69tlIH0pZYbfX
0dypi02yeZH9zZkhm3jVwQQBAYVDtIQLaFps2EP/U4p13UU+itwuSRiTVWCcm2uI
ykPvFR8OIVZQWh5zFMeeACKOwFqhUPvVadJ6za+0/ksFX8osQyJ2OHfG/S9GgF/1
bPJF2GS5EFUfDBmx+Yji+1j9vFIBIJF/lo1rYWwSWLAyCd5DeRYvf+OuhV1xO+b2
CXvJ3LH6ytarxua9R8FZiomeK6OLC1x4IhlCYoF9BnfebUdtPVPuCVDGure69Cu+
FHbE3Mzzw/GHJsjg7oT7AVyTGqI1prLQeVFWEobmoAvIoTfOqDmZtUDYiTfZoaFY
HMT6g4rxr8C/NVAacaZZ/Id8Krh3trKAHeyp5WUupAmUnpd/BFGd1A8QQZq8m6G8
RLs6J2Y19ZF7y/oq1VjXVzPbvV0AgGUNiPlVib450F0ot3m5m+KWT3cnw5pmKXOW
xABT+y8Uzv3c9GZsXZA0zoa9jpRMrPYEhyPuX4965qfgYaPJE4vz+YUHFcZnqDQn
CL2aU0h2O1c+AiDXR4fca6APx8qmvBW4kFh88BW1HBtJ+mNrO3avC6ncEReCFaav
jsHMb2Z4JzRCqAJEhQf70rnSffQP+wpxh7QBJedSv9C/hX6XUibCzYh9P7ADe6Vc
naeftz5Skc0+jIsBSL+Yc+JvUDsaZUEUhtm45HBmgdGUs/2zuqlmmV92SyOyWTnI
qLH5HDIuTlXwdK7cpMLBCwsejIn33qqhkoMExpF8CTdh4w5PgIkHr10hognJyXgE
oZli2KyEtuUZsCo0By37d63CGgWUXt5IOQgfWW8+RWXTsj4NdH6tLsnpCIhscNCg
O2UQ9etPQ8hmhLUZCIhwyeryg4S0lktM5lZJtBsvNXMwoNOB1e0sgDDDWPHO0Xzu
CwWax2yvRXK3ZYuXFC9qqTWtQkyajj3qYowwnREo5g9b7pX8Iq13JeNz1M1O01X7
atMYYOOjVXCyoH/VLYv6zYFIR7Lv12c/zAHOQxONO7v8tyD5ctgx9197P87Ct3WR
+V8c9nd5k12+4jOy8YEzBHwx1I0+lnhht9M4Zbk+aG6chMnClo9PuyaK4GtpzrQB
e/hwiJvUasMBEqTOMtcDj2s6QepaTcflB0r2eNs+3xzaGzq5f2LMWPuBrgTv2Egs
iycTH5NrV5jhriyMg6V2vXWgtuW3XlHfp02gI2T9upTiDcWG7Upfa0MNuZEogpF2
UPhR0WC0Dv5NE37TmfI8PAt4wMsSNA0Ww41X9YJVohE19E400gML+LV1WX8ZEafj
L5JvNZbZvSNDwIOYleDFqSzOkZzFXhanLkF6Y+zy3A7nRk+49lhVYMw2Mlkjp0LD
M62cHQZf2hhJe2HdQ7Z8MW8kWgTRhyfJAIwK5DDsvLQKQGbTfjEuLy7KczQvHS08
bGaUtu2aopd8Z9iLVHgq/cNm6WjrCmwp4TPvHnXRpBaxncr6DLNLQ38djQjaBLjq
M15YPvMvUpPPXvrASe2iYLb8zdNOkhs/X22BTLHwv5ChE7AVWn4UNX5c8ZVsw47S
7ofPsF6MFWRaAd/QXaCxVff4wrISgqi6zlbEzFb/vsbVIns6s4NTrROKSoDRmBrm
tMjXj7iUzp8a2/UMmsXIcs09HHH2+y0OZVgE+PAod+4MUL2fz5cOT4JSVfBn2HlU
Lf7rv17q2LfNvVD1Wm+0DABJMeBisfRBj44xgrUqKKFFz8ywPAnZYzZB7OKX2+7K
HrSQp1+E4Ms+31SwP8250pImyvBXl04F2DLsW2KMdT9mXJvN69o8h9pPLTh04JAf
N+7Ekdo9O94jYxJF9keNs4OkzQGOZC7Wzn5GUVhfJy53W+7fAzmIauwV+cUaFkMC
qEKk9/ns7wgWOKGrHfQsbD0UlrP4UsvbYvcdKv+kfUuRT2MddFiDnNwDCe+wrCaY
+hyT/85wM4CpB3P/GnynunzGJaC9BPoGpwVgyig4yYmB0H/K5AOCJg0avetKxt6C
Ry30zN/xTLNOKFxkHkxh9Gpzl1rU6z14NqyR6DTk2jD3lNSjTd3GXh1M9Gi1fGM0
zM08JYEusmkQdy+4ao8F/JKvLtWdeR0E82WJ957Ys5vStL2GdcEv+hWjOKBoq2be
h1k0BNGKmaCkIp9Zy95835nxRhl7SdNlfOfgIXyfTKhag1lRTYlGk8r8vKzopNGt
bpaBqKFAVcwh2jgsX+osjgCMS51sTQogEhQGTmXTa+NZStL7rfWwwsTp1E/i+YLI
3At3AzMgFu/CMUbI19wyberwWCf09ZoNtBGEY9OhfT0O4iEpFEzZNQB4lZki42Do
D9TUyRVjNDedACcYhgd+1O69tbAiB16biReFvN7bpha3uRL2CtotkrokKUwsoX33
NJ8dE0VS/uhc1ZshQQIjhgV0m9Se9NXaTIs8JhQMqPIRKkP45H67HjWAbTRENKCz
f1+HN9NPZ7CqmDRRWQhHHTIQTjXiFZ92vPBQs+SCkKMY4eq2qAXVJzQJEPQR0Wct
oJtCvI70uX6/ztctuXpoiwFoZb4eEOBPzYmN+y+paVUd+roOroG0Q3qCg9UnYkKe
0iIlxE56WQs8jrtclTcuBbo2MU2acRXN5sfk9xYabsqsoT/5/jeKISEh34FuSXM5
AGoPBct4W1/sdtNnLVoGEwzk0H6wSkuw8HWUVAqp+oqUjmbw/30fvw8Fb1ymgr25
zb8MFQaoWyw9WspNusfRDPzXzQS69Ej/xzZpsvTz1o0bcnbMmKv8hS0E9rQLKrqV
0PzadahSLU/Rdwj9BZEs5/m9rUdw04slNQB1qAKlEzukopT66UoUfIlLKaNPGPuN
c42mugPxpBHozrTmovFZzKy4+uS9kg7le8gW3J9PhoeZis8KzBEgPwHBDA6spk48
weqJxKeVI5QNBRuh8+YIjd7vQHYw+NHcfMMalbt1uzDxNCOdERsQIGXVj0kc0V4F
2eDRceuUvf7/JnFPbDJPCNjd1+DA30PCeWgp3Xfauc/RXtT/s0DyIv1KA6O16Vgd
+ZzT4e9GwHK+mQNJG/dgQFE0aWeF/vd9APAbvh0G9eSytEfLyESHOwbKZN8s9625
RiAs/HRRwbyZY8fhFZYtabdaW8SYH/PMqaj3PQMrFvvF3cyarbGCrY8Hx8n42sPh
b5t0wjR6aM9RV1+Zf0Kj+1/IYXeZNBoccO9A3ue/nDkztTzdUKk/Rm9yul0zB9gN
O5Y6GD3reP08WA7pCQG8ZrR5ixC6AftRsCBU1KCrn5whn1NHr7wbYTcox45XWsF5
hADQKlJ3SGOX/mysvubpVr8tnQMUyOrzH/wcipp+iKQRyhCWiRulT83XV58PhNg8
fOJsBCETLz+By0jgJQX8XbDANOKMYv1VzntCo2jmxD1pOTGyEEKp4zpVdzMA/aFd
vl6KYspH70dgAcHSWT9y6DsjnnOYINa+9thFh6hkOfLpE5Y056JIsV2ZwkJUC9hB
C+WjZUicfsEWX5F2D2mzAf6+jsgG8QyjmtUqOpV6JOzre5KzA9HtepB4Gp0wAHn5
VZcGYo6lPZYuS1TZx2zGEp2US6p1mPl36hSdA+G5tKBPHT3Jwgsc3C7AMF5rn2bV
IkObM0hzOd0dyiwmOC1eC+vXt1bGHFx4ImkmjWhSQdHzzJBpIksL8nbR1NJsMS91
hoe/4MeLidlVgSziZlBVrFg4iLZwSPZK8HhLI21tl6XrpxrlBIUE6fHAVFRKy545
fiP1bJTXxmCssNhBN1NEi//E3sTgjYYnfAZF8Nt52tjxHndTjaE8+22+HawZgj31
ohU9+Azhc44Ltp65GcKZvtEKwueyO89+m103u20v5h2tOW2o+gF1QO85c+rQhejP
SXA9Bi1wJQ0KzbdvN3PZBEKd0RWGGU+zFTDyn5v32UBo1zuE18cqRB/UWwK0quf/
2EZdEgKISH04ngGDpvNeX0fGWpnMBdiw4Kb9MZVqvfwnizi2gCmlVmgbME00/4po
bbes8qdorwXuMgj6fvn5geOgmu6A0X1gW4OLEfxvd3Xs2aMtef9F+oWNx0BH01rH
AEbB5aYzgY05cuSILUgExnBWFIjnWVPw7VTPpKx8+1yvDdYvuivQY/3M38VToGJN
hTY1nURF666dS7Xh5KE0I5gj44ouyr1JjbvYLyyrHOCB//GyuWVfAA2erqfqbyqh
u4eImnEezBL9zj1OFjzicSfMJHFFPTvTB+aZgg9O05V67rM7FIxPLB9hA53SHB6K
7A206ayJ1dSksI97lE+PF5FjyPhYXicOyMwX+7aDcdFTCMlDd61CGcoTUe56L73o
icmnoDuv6Yvk49nUCxYEVINtoqDJnrURVRdWk2GYmjdNPGeR8peyIE9XaCmIZmaL
6wvHPbo73eXt8j+tVtZEhYucqzrCpk4R7H08YJIOaN3WSGac6/rzl9b8H1QxHywa
+9OxFOeZG0tgHULTfgGBHsn4QxjkBlp3xXFJ+joTT4DLvOmUO5pNK8CI5z5q087V
4hTpzQmJ4sc240y3llgVv+yyokbyVVC3sR6uib8Jkhr8Pv2VRRt0VOd6BXES7LMw
Ty6IO8+MDBgUWBwlxHy+7EUaJR6PJSy7WtNVtvS/DztECsJK3Tl12n21aSpvOiwP
py60d8zmK2jEZzWJ4Cy0oApYQluj0gPHuqsn2K4m3TuR+b1PPZ7do2r8EtTOciKo
ILBEeAHrS+JpKrTWZEq5vBA/TFmFmAZjsBmoiOBHf+em0SLAGGAdWANAAPou49hU
YKdKOvnOPWVgtUyW89Wbt3c/rRYfGFpeq3I7HfyhWQ2IsQ7lMCoNChBI00SgNimL
/B+JuGZVlHnErEnHjAk1Thc6qLBrTXH2WUmZoqxOnCNeilv6c8l215EVsWMWVO2b
bKHj/5ZpQTZ2RBgE6ef5rWHn786dv0B+05ROCKVZG+DEuom8/gAzrQWS8d4jgxg0
mq259ITDq2mNQC4NNh7kfgVgQ0uuFinLdo+fpCe/tNOHmErYEHQzaW+yu0Bs8T8B
L4zAg+27alF9/jsXkr7JG0X2MsYRyPILyMljJO9RhQNRbU2MEXj6D2bfbli/5Mhd
E+fteVfgIJIkwbjGiRmFv1pw1y5/SPO0bUi71h7VsA5AsP2wDe4d3pJc3GCNnlot
3oFPFfDMf7i/LimVt7ezGelgtNVRy9Qs1bikXMx+BeX4sFUceILcOqiHseha6v0M
kkpFw0ynIPeI3kDz7+r5IftQiLZF5Vvou0zPb8ybRzjXmNwI02Is8eiHhXfzCjQI
2UOJCd0d7Qd8NBQQrzp8pqjOfH6/npXsAVi+mlhaTK3UrlLOZx6+vrgIeKFWoGv0
OmzS4c9SjrgiCs++G2idBRP3kfxj9mR1bAtiJc8TxRGEYUzrG+B3Y7prb0jBVHHT
nUcjn0mjhxoNiW9t0rDzkdKsBvNDBUi08neyvHR6uY8sXQjl8kHFMdB/38FMAdHs
mdqIvqajWDoMPFR8z34+CnE+/aVGswwbdGX61NpOq06WE6INGE/uqBz10zWsty93
5nWshX9j6Qg1ZkjB8cfplK65UV5pejIPg2U7x2KzT40xl+aDZ/tr2awOVPXxGST3
SCa/XaR8KCCi78G1WUTsWspzTvMo2qUncV2d9gfIoHQ7NK6+2GvuIWD3ph4Wfz1/
AtPBb9x/bEamszXb2Qj9E2+VcDA4i6iftJdfPpgwmiap/wX3V/nhwg6Bu6N1mHZ6
NN15JxoIQV92yZd/36jOJ1XXAitK9XgB2/gDbXcgBNIxWTnhbys+eBNonqKoeUAn
uqFKrREmitMdZye/w+ZPSCMX3tUKQunJooqYWY2RtMdxqVOIkpbPNwyE9f6cLEuU
7WCvWFPgLvefj3jRHqv3K+PEvBJuLO9e1p0fbllAs+rxRs3aA03Wy7CtvRuYkrFn
AxIY19R2vyL9EyCYit9lJaHiZv3fTo/P8ZxCth86aDfhIJh9Wl0Qz9b/deyfMUlj
00YELjinNcmevLMHFxtTXDFJBpm1E2wUO9JHOKNLi517T6gkkO6RQkJKvhuzEnqL
J9Ak1Xsa0P1lmPzUV12NALVbfbMLi7LKCnLBmAOd+qnCIUHuKbH3BGLQzRCXWrM4
8/9LFQYfbAwDBxOFPgg5Nu56qoh974XtbUX31B5zCrNuHS18sgH3zhyzufzUegZP
quj/QYfCal9XTVnnJjz2qxa8jH923LqAHhxdjJzt2Dkn0UKf4GGjFT2GiqfLaWTK
mtezLaQA3g+NwQU0doSj4tP6g71EwnMVkEoLq8Dzf1yYVqSxmjZrdNsk3L6ArzPT
2e5tZ/E+IznZNNrnITmg+SRLlzIs4NcI9AvWFPdCp7PHg/NLOUFR+zjwg5+A4Dyi
BpKEaYhl6XF/aBsdCeOtCHwn3G8bF4E29srVZIVm03Ucc6oES8HydTjxyOGjUUlA
+u5Vynziwy+O/Hm8QcekYAf8MD6sipdIuAXeoTU00TKkxPvUbeSWocFT4dFwi8PV
86uQtwHyZxgVYf87OcDdLZ3oNgPxc75pdqhSWoj0cL/V7/gO4o0hLwIH1Qt9XcrS
xxGqyo8fZhIO2cx+CqsNw+jXcOArgjQDsR3hxFwwv2d/dx2+RPYrIUKpFcdI7Z+T
AmOFNUD5cHi/bOkL9D94RGvxP5IKcJ7G4fm7iFNwVjc6LD0qvgYm3WMaMkENMWy1
UpgkB5hqzess/APDnjntHm7mig+V7zGDkHbZIxHQJZuLvkIcH/4dyApLagKXylc2
kBwFMln3cDzmN6SGrnxIN5Qx7AVSx0Yzy43NB6VZCwmezosp2uVRwjjtSTXzqzmo
QeH+UG1fZnMEfjJFwbhki5d3FzMex2AThUUREZ+GlVSRM/8ydXQHExTuPQazqecF
Z+FIbmbjAe6adKVqIyfrw487wMHhQCzv57bxzhxy8rBYseZ8poiu0m+R/xjlWv6I
NO6yEAgGuxSoYz5HsuMaRpaSOGXO/1cC12y/g2VWHndshrIP6jejpuQC5wR7R1ui
9jCQlawYDU61+cZOWBrur8Nabto2x/0z0KfNpCT8X5tFQZ6w03bYChKUpMAF2Bdx
nseLJ71p14EmdtZPXymeG3Mlby6qdJYxe616/2nLUoDwVJOhmodjoHbS4hAbiGR2
WBS2ULAzI/alNWBWKru8v7L/35EkX2cat9laVO5LB0p6uD03T/tE61N3+rckloaN
2/FlySr/rm6vhWOI+fTmEwdINUTMq9Jn2YYSr4UuF0j+9lrNJ4iNU/zpl0wPh7UN
28sq2OHqM29Yi7J8cEhXsWRoAVR5PwaxtTFrUpkLo8eugYqQXZYELsZcehx4v9hB
i6C40DnKX08OaNTy6POMgF9RjIPRen6vdjnLsPgI61gCv12Y7R0x6hVUOwTeMOL8
cRkV0RReya5Gxp2NM3Q7ofQ7RfPogymLWb2VRjJc5kb14VUuLyBxgW8+dO22s8/H
jEDQ1WfZAIsTl0jDukzmXcCBiyxfuCBHRjUdQn3QjXqnDwLrNFIbZ878fZcJAHqU
u4g5gGuizt23m5NQew7irMdsagPLgE1EnizcvzysiPUYYuW07c7YfFf/v/j0gea0
WwLfbyRxkSYDGXGkaidyQp4nGzHudJjA3J7Dcuo0KTjGgINHdqfRQifougEFLJYR
N8+tRS5EEYcytoiUj4Qfd/9fIJUIRxZexQMMBTz0p4h/3HDD+yoJ3TpbOxyiG3NV
nr5oQLdCLxN7H3W7hRaFCK6BKxYXfn0z/owuKyrwAxQdo2eZp0diLR6XqUGdfmJ4
Q3eiStf2APz5390XN6sG2lNVYDxqs5VNlmuyYFDbsB7zibecJNW6Tg/saT9aA/TD
XOj2d3QVDGPCi21YO4ColB1mIXObZ5mBeGfC4oMDuchAyMI7IoriHlmeA8eg2hp7
BtGoPDosr0/Zo7DRdPTj97TfdVHtNjXmklVGBgJUmbE61lcKMdVBEOYo1J3TSI+P
PzzB+O5bHJSNWdtdGWgIVdertMI9iVireeHo3jPRdpTCL04oSA1YwSZXMZ+B/BQ3
1TzU3h/8nMoPQBNzxmD/AcGaSPARn0UU6YH89PKREUbIT3BFvU2xlFwK/LrZ2Xtj
vAJZLd16Tk1ZVqyxX9qXIEstbBtYAhOyhD0qWcJKh9vp+ty/eeUHf+QRLUMRcazZ
GH+dhcWdrE6PRmoWFAuc9GOdqmLyr6P8k1CIBmeSN7PA3X8Ho/DcDGkxGAReuy86
1GnSdZ1AmTJYapYz2UxdcBCX+ZV65a0CU6muZEqImvogxs6fplRlxCrqTKD6LkFg
OMmAmRZ9Uc9S/PMU3VEd1PFjpSyT9UCx3HUYeWWIuiRZ4T3bFo/vpbQQPWKoSbIP
w7vZSOcWx3xRNlk4I6ZAnKaTdwTvWN1Mxr73koi22V0ZFt+7z1RRGZphganaeCuM
9vvamJkJ6JjQWVTZtvan5EKZ0YyIXMmXkzs+07GoiC23zHlkVPL4sl2+GICN7lHF
44R+PIFfdWH5cI5Mk71I0kcfg+hRveTr6R0HWFzY47JCNZh1f9ZQrQ3hnivV7cvY
FIJcI8vlTnKf0jUiKVn1DsQkb6CBNL+4/g9uc0hZ79AlVFiUPasZdzrH1rkPCfvb
6XfR42Ol9nOM50cF+bp2XfGs9PIdOxDv1PmplolBz07jP4YLq5vtPOo2Vgg9RjGP
kd+PsRquGAG+nsW4GF/kQwfbtcKONOowqZB30Btx7jjvm+OI+ZbWmXcnvUTuK4Hq
P6JCdlpDki9gcmiDNqBlt08zT6rNmci3S9mD4bqwbVrBANlaeogShWz+EHr3EiEi
oUBqAxm6jf29tt4h6uIQopR6bFgqRGyBPUNm4isLG1BpZRJbHhD7yrXKttLMxIC9
tvSZG09pMIJt5y2vfiNGyzB1Z1NdYhZLzAnx5pvai9avrJ1xKr6z4ZsPYp+Sb146
U4PA5TKG9fI1aSpR+Ti9eOLhhsaaxWHuEUr5K5iSSUUej3B5TbMB9nZDIWtPjQTS
XmlOwmuZJLEVnNibtZRfoXludI0AzaUMeeJbdriS8R3bHskI8Wk/6WdSpnV/ZAuT
CLHQNucKcK5xAlQqRqsNTrgUOh7z6rXHqR5xrUnqf/5MODmHNVWWGPciUQCPIwi/
0pgGxCLBhH+epAiwrejw1tu3xvJorlfIyceXNXXoGGewcceBxEUMjtdjNme1i7bO
uzlWg/fKgBTy4LH9gdCVtNSVv3uDuHWHJB5+QWRrSUEUQmV4YskSXDNjhM0LQMVA
NqpVNh9pBHlO/p+wELtpUwJE8KZ3ONplZbVEpw0i0EF+iKaQubyNbZjCxCTVp76u
Jc9HuG36XGrMIV3PDoQeQXTjeHC8gFDPCT4rpnENZQIuAUG5q+DFOa2a/6Dovl7q
N9ip+D41dLITEMO9G/lNpF11RXeP0rdO/9g0bTHBxoDai0Oj+CqRSsdXHdnNLlPm
vbFDgqyE9eB3Aknm5PDZdmJfQOhrtfwrLNF+hP4DBNXQJBpe5CsTjETpVT+WD9Et
PHVx+P+2/hid0zlbO24NwXd7U+ohQ/W7k9anO8dtrhO6uqSxajQMIwfcSe9nsRrL
Wm1+s2viO2wfs0AVhmJ2GyMhyJW5qJoksSv55RcMCduk8hse7coCT0tKubtrBx/l
v67WNrKNQopv4s6pcuuH78iO9tPlgzVzlZ0E8q6+0v4rsaSIptXvjVc+Q4Cy/Qo4
XWEpkQv0FLp+hKk7bzIAImmSQ4bL+AVie9RH5ir1q8t5e3krjqf5NN7+Z7U90LkN
DIPNeZWfwoqYnhxTbMkm+P9onJj8mHVnZ9I0huOVxV5SqQ2wf+/f853x9NkcM02a
qO1sdXVvJ4J0ZoOVb4yg1qglXibEmwDxKAvFGA0+LqceMix5lGvi82dW6bfXOsqf
9ucTwmL/up/wQ8VRvSlnE27XVFlR1/1alYzwgnG1lbs/VP0qNcDS8IDo91Bdmu4q
0FqJUQLxSZo/Wi67hshxe/UdyrnIo4dNTk/LhrWJStAgOYvIfzQKgAnzQXYwmPlJ
rORjHVYVk+GidRjLWuyPZpLKRtINfZ7lXWMgngJi1in5a6nPiBaekjeKH1DE1IOO
Xkm9MNjKak/f3fnxvpynAThoZnOzP4g3AxWR6DK2sTv2xmNitlib7bI1OX3kLb+c
0UrgN+h6dWtZKRDIidBthF5ykZL2iDl4BdpOmn38YVTLe+w7xqAlGs2cF7/oQ+mx
5BSUS3RvbHPUSJ5r/u1E+3KhsUvkxbJ4TG/cGJKubJaGG05sdEO8bgvmGyXr9Drj
KDHL4oL1noj6mo1ewzIZvKDNwRNRFW7JjhtcGwocb20rSvVNijm+W4un02XU22ey
qIF9jAycDKgZ21vcaJzEICtz1qKxbT1QiVL+3ejDdlLxfZJUwFElcSwki5JV3lq0
6wDAVqus6N9AHkzRD1jqfvlTg21TMqT+Rzufq38IqX4DER4IZbM5NLwsa5/uOrbC
/hDdCR4T5X4ukcqeoKsni2IC2vQ5/9TECwcFZCqbVdAhgxsOvDGaPKS+LEwwUl6X
LYh7QA2/J6quQS+ammI8vt/9IgIWIGrl6GgVM+bEBOY95Jtaoqstv7KQ7pyUd/Qu
rK6ACzR4ZdSi95Y8sBsqA72OKv+/LWmc9K5BogE4po8gfu9uQ8zkXmyp6yJxelIZ
Ndr8CeNTdPLHpGTaYKIuYeaavaz0sYp4ObTZK0+hyFUsQsEARtXyf20HJP9RUx7U
jbhxqks9ODx5BxXFHRoXYH/J2zHTlb89DZIba0BKS+4tZ985XRiaWhQQNu51/fLZ
4362Dy0lEW1pAfzm5LRZfILrYtlf8usIbTZ2FDaI5QGqqOym0mEtsuSaYwvA2nNh
ix0PToFXGlvryD7sp6Gpfdw1inaJc8zq6LumaZFhQyWZt1IDODKB92iaaPOkS3rL
H8mV8R9cAmBCFmX07ltZnfK4qmyl/Hh1zRb1QfMDw7mMzT3MZIaskfXnnRU1Bt7I
zW9IErlz1zIsH0vbPK6CbV3yVvZ+m1laeJ6bw548aIjy8rOQbly19KDhLFQdopEc
0t1b2691gzEiH7Pl/Yl9wAB2k6Rzrb3Cw8D/QeAgjZ/NqhqrgcuVl+WnEtWFHyyJ
aKl5oGeJ4m0LldV7MYHYsKyucu80OmIw4hmkvjm0bdwQC+7ilmPOjixIv88St0cZ
skYDzUPyFkhzvamj2P9QoLSydG0kgbp95Cc+oo7UVFTvR3RshpKruLD61yohiObK
qcLqzCiZGTbFq4aj5jmACIMbNQW/PMvUrfbnertqSpUxuu/WIjMzCaSSTCwTNgSo
lC2x1XtFvDWX1wVm0wmkJ/0MMl2xuqZ3nSM2GhF9qInivRyR3ulGv1oH/1kqeOzb
2w9Z/SmIGvKEW7LtMEGDwEdJ7EIDnqlDX/gVVpMX5x5BNrX4BWFtZTsCEt7aNJRv
4nY9LIMlPY+DMQiOZg9OEQ/9qiBYBqd/igjRbB+ZVBNSPElo3bkSTAsrWZxzPG22
cUODHAUNrtRUf7SMbige6KClLWwQKN6xt+ao6fYGaoLb9007nQBPK11FDf87iTFe
wIsxuDV6Hs72cGJXJBafwvZo9fsXqiqMQm0ArY8fCtofFFupXNWDq7VxMv5rB/34
2e+iMYLCmSwa8vG+2F8wJKyMZqXavmhAJnrzFzIwvJHlYOZ4TLT9KS/IVJkhgSzu
8JXsGzfIJy9CBeHCMuhrkHndWYQ4tboyexyZxT60vAHm6GS0tL/UjZfqgr7787u/
GzhofLoqtwkd6jCCPzVBMD5gaAUMKYj1M8UIQdXC7+6Sh/CHwiIYzL/Rkxr1P4Qy
onhOHFd7eTi5z27nj3xHwmYuxdZ7Br+nwGHLnYPfqk+5BWYEJeEWHaIcZwaX1ZP2
kjF8kc5OxHzYf+dAb1GYuyeMVJX7zAeb0wIJg+oWEOmlTreMVfPALVK6oX6wdCHd
SGdZoAQGKY8OjpbVAZc9sC4L28g2QORnbY3Zs5O83x0Wo96CU4WVGEzTz1aoSN1o
+9OQmuTJ2Mi6V6jM/gv44yzuoHIpQOVvUyHMraRULTYFhKM3tR04SfPxUGuyy1m+
4UBDeyBc8I5PWAPQzNAwrFyulUkDsDBPcG/yyUriF5c7cfv6ILRxpRr50EnIShjq
dHaV0GCrDzWmOZHb/f6ccG/n45rkOM16Yopdnl0EcJtuc26BjI+lGZZ3rL0xpU97
8fUUPRpbyXW5/rmqzy/NdL27c1UajJAOYDWsz8RUIOP+kESa9sKpsLwipzcawedA
k+46697xBh2rp2Fzln3BKmI2RN1NaPUc+pF0R8QMqA7wVsHrwiMz9CETirOq0+5A
/qAgE1AaXlxAtp8qEFi597oqgSXA5C7lLUjGzOh71xsqWhPh21ZiQEQ+TswD1/Of
crTjiJl0dfbi6m3bRnWkVtbk9ZB8cKE92JNMFPXJLPkubujrSiRvIqCZinT1xcqS
FEZJo9IuNBmVQHeWqSQ1t8pOC5jv73L29umtLxt30KiGMBxekb1pGBvEsrreeae9
LlUF7wuCh3Ex/k0cQCl/+V1pHgthhq+ItzJODE8V+Xx4P3e422Sn8NFysuM3u06R
dsm4lW4DtV4C7qcGCLy8Dx+PFI4/2XgZL5IVSni30ZIUb5jqlyXz16KMqOxOsyfw
hQiVEg03A2QkfK7VQnBj8wpf6uNe/1od4ZGNbukRpZIeL6rmOPI86NB9UMnOJCA0
WLYgpC72uMWjhpx3dcdzYeeC4ocWk53gYFQSzen0sNIh8qbWzdc9htwzwnHAWtX2
oTJ1wxFq/4ryoy9EAMbn5knoGfId0x8M9oykDofArTrgQBS/HWcVJjpFoejpVPfg
O6kbmW88yIXTvq+0D/rsV9YZA4pb6fR+KcdtdaINaI5zas3uKpv/Ua1waMUI5Yoh
YJdA0JzQ2oqkMC07xXmzyDm2j4c2N0Z0KoiuXevHxfzP6vE3NmKWqJXOdkK49R37
f4MpeaXOT4M8325zMHJeSBqHNTUpXMIjxNQrnoqKY/S7WaxuSOtNeqqgXb9dLmpw
iuUqIFzTqGdkh3gLh9G/Iiqj+tTKUWHfbVRchpDAOutcmJujYxVHXtZthseSHEZy
E2PkZrqAzwDpdL0/HTCsvcOU9h7hHDPtLH+tt4KMGWEHyo3pHTfES5Qd1VEq1Hf3
WAx/pdIqcpJgBK41/rhKFnS9qXvYurHVWxngBBMd4p2UZ+r20FuiSjYSBiqn8Txo
k/R07U1Ez3JXLdP77K597fKRTX+Xc3atOrZ9/Mg4EpJqeyZIHAAO0t97Yn31bi8f
XHlptJi95ze0o9OHU8q23o/C3xrfSrpX3Lk5KA/jWvg9mL+xIcBzGNC3w35XTHDR
nJ7079Zlgb4+OUGFWEA6uXSkljOWNzqoOB5sA3BY3M4ZnZhGDtnSC2Ynwnu3RZZA
E+1Wzis1/PXQorLYwKOkflmQijjwWHeCcgC2VWIyGpEQcjkC9MBqXwNyZy2M9GSg
nNboZiPa1jsvamVmc/weJ5mcEEdKXt+bUNgilUa3JQfnoveXIFSk2kZAYP17UbjG
U8qvaQe2Nk2ybfcegFq2UqT276rnnL3FFwXxiAH2f9aOWGa5bi2WYcErKy0FYUsI
HA4uCfZqHatYAxyzGd9SzVjWAoIwU1XLg3nIQya6LApIGJ7c/EsZegPy3WdaeN2v
yUD4Zo0ZcLZB2Fsp7QEMwI7iOlmboKTstsuW6b32dbEgrzdXtDE8A4RVX73cLdYg
ZJakQfgPx75uFWdHFBG2YaCcIiG8TDL38CfdRw0gl3t+M+043blSeECcR1+SGik6
Tg9PUXY37tg167Zdx7EkMqZF00Bw8y7jVtCOrb6/U4AH9hxo/Pqb6rS9M2tZMdxJ
hvcoOGwcoT32P7N5cCfZspOBUcNmI6E165K4puHVLAaeYhWm7QlKca+aSdnpyY7V
EImCi/bueOaWJOXaG90EX4lLiE3DMlS1L+/Un0PyFbh+FM1p6UEzsAeXavj+ZkZy
bxorArSjOd5FgXMnm+OquO8J4Sit+jDDSTD2MspJcFjQurZ2f8EoRvxlJzhDmRzT
k8yqdRL/EajM2y5WF90Vgi4Yxv9o998OrC95S5ZYqfLQdC587oIs+L2LkF/mDkcw
2XeBEGUDo79V/rZxP42LDSrbRti3TU5etNs//aRu7Z/IN8wx3ZomqKqyRl1VpJX5
hkoqxJjPzBns0KpgHh2uyPUeQS3pPCD7mmOS552rsfM2fGFL83I6lXCXUpbtoOkS
erSakYxTMgw2U4YJwhcxnNmU67cYNA6owi/FJsNRtg+aXpec6O9B27MnuJycQAIi
QrCjcnFCQ53UavC+Hq6SFZ2R5V342Csuhy0xYAVlyXg5OMMfU4+j5mwV4A7Uns8a
MWyBi0q4cv4uC+vld9QJAIX08WNgqSVjpOAj2LZfJUFt81FLK1McqJN3Eu5vsgbD
OIYElgLjg6Y5HiANEKTutx9vs6NjuGkUnC4WCDOueqvo2/UC/NF+9VnEz4RTOPhO
QoNkTU9DhK2vY83HDMOxPUZxyfkRMRuJJVzbxOwp3bGVWnqgbqOojAG68pIQgVYe
KVlE2UbTw8Vodxb/AsYXlWXh67nCt7Pa+C8yBtVWkng/kV20EzdqgmM3b3OnZrAN
qd2CzLCNmOV1DgVLQOsvUZ7HVpIYhFOVJuK50ggLhpQ26yfn6cCa02EMYM+1Mp/9
K3WbTugU9UAFGYbxDs4F4DLRH6BoD3De7yXEv6aU/r6T5mxqBzuAl4tQGlXcdl6Y
YIDRcJAoBA7BRQDcioKzQiwjTC9qkJ3mQiv2dLDXAb2RJG0MzC9gqH35F+F3xdV0
e5Ps18d5KqNdcKYcmJ4GO4zsZpZ5nmuplrtoMmLalm0Qwbz/jZBtcHMlp3pMX9Kt
nJUVpgWUxzTODKrIGG/6eO0W+XlCY4AbFcPI+H1jH/H+p6boeR5AjSfS53uSYg2b
hmHsl7nCZcJBD91zRDI9ifEdhKC+oig3C0qYpkqFullxELa6oHp0wpjpKkD4gU66
u779784VByXk1KjeHUJushKSEGMeY3LD6JuQmd4iHF4ME10pE+ivagdWe0xFO5CF
xGfeY3KGZNNAdTtKOjKT0wB4aPbKubvNo3TMh/HAimP/kb079qVEOed5DWKZ0INA
IUbBgB/tDsIOIU99r/mhbQFBzb5TLe+dWD3w4h02Xg3ByxDJ/xzpCjgxHZnGZzAp
lzVZ84i8tbU+kvq0E+Xld822EqGuNOjdVPyKmcnKn7LwdqNPidAVCl1/ASeize66
rrx083P0miLWbHLx7cu3IFUGs0t8nqeftIqXICh62wp8AdNMx88jURwRqqqQRVhG
k+6A5POrUcjlhc/aGEYSk54jo3e0L9OYr054V42c1SwikTgKLwxiG1JsMVfqFEMP
OlJtaJegf+kBbgWC0wV5n+PJmuivtspH9aMoGK3aM7Efj5dElHRU75wE/CDxNEJn
HwA02kPYFfTv1mrsk/36CUMT2+H5+10hDNAaxoTJT5KGonjkJaHvPo7gRhenkprA
6lCsw5Pn6F6WH0Hsek+E6s1IitheXoRWwVmgjUsDCXtqGyWIn6cDqgM9pkI5mNai
1Df5C4vZAJzTC+DXzLRrky9zjD5r9Z4kkMqC4WVdrJrQdtCoojvPvagR5zP1aCiv
BbNLqcyLN1pUBaJIyDbrRv0+8o3vZJqr36byK/8vp6vQUHXYq7piVztBK3yk9w+Z
M52LFnglvKx1dd3lu8Repzwak1AaNOYqwie+SZJ+tMIjgyuJZRrzjE+vwDMv5MeY
nkgGe6CUNp+hvGHg2U606yehJfc0ZbT8FoxK99JXNpb2BbvbE5Oz45qQG8LbuIyy
GFy2k7lh8pcZ6JI1/2bGFIh6wAlOjn85glfpQIz8eyXSB5cVJ8c6mu8Y+18U6OKe
9rPjwjtqCF9T9OJlNyNahMNs22GzBmnuRQ6giR7mVEIc67O2SsD6AxGeCDX1s3/S
ZURuxmmDZg6ISc/ibT3Vnfa4420B2I8ekySU1vb8Y7+cJJXfHKFnzRN5Jjhf5McL
6L3PoEUklpsxvfXkXUmNVI1Uj4Q/Q+QleWgi05sIB82iy98McFAPjFEYspGiepfX
M1IFZiV11juFQsBJO8gIt8KkmY29bqEe3fOhgsBX4WrYa5EqWDsTdfBHyHfGw+rz
D6ELgagSKnMHATMUoWx154yadxK/erSW2occ+G8sgctaBL2XcGmhG3Jnqba31JIe
atITq03ncpwBbBX3Gchhtrw3P3rAk8EB59QzaFLoXlZmZ0xkerK2VmZSf0c1fz8F
/6+NopCRp7LJIyweAzO6HGFZ22D7K19v73SqRuW3ud+vLiO2Vcb0XYndAVvmZodj
Dn08rRLUfYOG7VTa/tGHrxt30XQ2oD/TMglaOp7xSctkHbas9AkWO+gTz1hjDTst
NDH6DvQBAVJMy3K/uH8PUWJAs3TkqE8O5uMN1cFaArx9v62ffjlyBo8dKl0L/fiS
IkYYVz0GflBO1i7pLLed9Qx4ggVGUEZMQyLIVX010AZSYWf/qLE1HgQQuvBw1eMH
QaeFXpCYffw16YtQ5DscaUmy1dW9foTWJAopBXuATkfAZSdbFOKZavJttfL5NXdd
OrzssLKTZYEoxylzUizJqjawwzTY4+oEI3C750EEnI5tB1Ht3+eZ7zwq2Y2ZpwgX
3w6M3ZyneIW/qQoYSYaDDTb8hlmRReArD+2iwzC0Faz6yzJk66GABioELwi3ROCo
Hi1KKNJFwWvx6Z8uiUoaQgfHV8XTKSEVhqfdOXAf+4rdT1Q/0MvvW/kRqcqNk68s
A49qR8ZCnIoa/DttCfk7H6mLllIL5NIFqcEZbcoqzHk775SJjA4qxGnlj5v6TN+S
LRxyrwfUM4Zh8gy1fBdFJlhauoWIihGBGrrA1r6UeS+zy8Zn2MceB5WY3oGObHTO
gPKsdQroVFwbVPzEvTbC/dL8yPoIp7LSs1xMwwx8/IFuUDQWxCATCEzwlIo0wYZ7
G4ptzqJXLImKTkzUi2kKu/l33NKTstL0HXf8wLXyaeerV1oAW7zlUUi/CdZrtylF
CI1CsOQXi8UXq0LMw4rgwkzAxahlSZk9JCzrFhXyqWmo2yAtvaMKdqCrp4fhtq0X
H+/nenpUykw1WrRLk10H8WmweU0Dgv2RXis+rIHy3Aw7AgDqw28enmYcUrZrrqJh
1x9Pkrx6Cj7VAx8+Xyatsg90Sa/K72RXj7zPWIunpUVeniM3yMj4I6Vf+LtCYtxr
/Ba5IgtWOEQE9SbH2XOrIRKc9PYV5jGCugjdMgLGQHfivifdUPPxggQwtjFDwxMa
At4gx0XxFm2WI9OsmKaR1b7Uhf2zu9ECNvfqE5LPHMmJHKsDAstea9XbQwyMETxl
rvDBS9MKt2YAuXPaNneQXHA3YyX3rGVpQyHdFsp8kURC9cswUjzIkgW8cbPyN+SD
m+Rfi2xqh0LgWmXi2JTax8ILXzeyzTGGIt7vaoub2bhKy8hwACQWTa8bWCp1bA2C
ESxo/LRYeQuLFcLmxV/li+i78G2beO+y/NwB/R1ceHuFfCZAsTQ8yAbpH4uXat6B
e3o9E5pB9LAV1/0RiKAImyUY4bYQVJ5crIWw0f6HdA4f6basiBu2J+UvNm3iiErv
6yuyJcJp8EZH28wuTEKXSk5qWjjdlw+ZYiPdrtP4oYBX3pmQn8u9rNlR+/1dVkFt
CqhuQhhAbINMdQApsiynVZvF117UgM/P5I7cFdBvg5FHTpCKx8YTQEV6ShSSFzoG
IFSOfkOtszZY6JkkH1drwAmYh6H6GOT17C37BgOcLo9x9J/CJNl5S15ERFwxxvaO
rC6zhJpK6SJEcZRDpN5EK4Otlamph1xlyRxNVKPrXYhj2iCE+b3GKzk/d9FCFSrE
RT9EJou5zvlq4NX+bc3S6qwk3kV3nl1T+2DZfUhjS+//dGDbW3DIqdHkAmlPWwhf
gznc9A0kgCo1xow+ZAFJHXcd0ErMCYiDxJ1ud93SSHIkWcqPnA41i+wjB6rGhihp
WV/6g//F0/P9Uq3M//Af4RNb68qoEc/kZIoUWLhDDYjwNmuUnw14vTNYQi9cUcup
tpdU+lr/8tRoa0yTsamRraw2lwt4JMven1Pw+Vi3/5APp+b507Mdtps/g5yClemM
Rx9jOnv5klWx3AvyE+1txDbBrrT8pzQfOCeUA3NxxvyR9+dA8R+KZwgCKA14uEUF
LK0Czo3XUnyNkvb1FDLEyrwVCO/yVBnZxVGXwlD1Qe2ZI55FYj13ahekTaoufKGz
PQCfS5vNoa9QmtaD7qclvPjhIte+j3s3zQn0RnNAVryJ9dMzJPjURI21Rasqqk9d
RVYY5bLTgLIiAXC/hNte5+4ZGGnsIcXs6fbdTHquMkjz21lmQCnUEjIzTYEAGtbs
ADiGH3IIcGsQSjmiu1ttPxW/EH9bHVYbiL3kuvDhf2a7SPeuIWVghkVyrhelR9xl
Qt86koicf21qyUKT/dAGzgq6W6yTNQX2QXPbx6jeJS5F6YDLwzKalFhih8FgIP1G
rizJAsZJrHte1SDb+JGW/3uGTmLcTiIM0gbJfR90hXEh/QNDMLmFbzAP7xTPjMNy
el+xn4wukg0O3/Mc8pKHxmoXJtLDzZVxlcLZgghQcl5XgzQP3c+nhB+HJ3ns3pZu
+8S4NJHiag8cxYFuClrHe8/MIAOJE8uLIxrQEpwH1eJ0/XhNI9hN7ZHbIUmTe5fV
pDHyTOXuCiVcmnAk1zD032rjZdbTDnHeJKbW35lzIlL1KSr1ei3wITS9npASp+aD
406KknhhqVN6zDZL8mkf64O/up92we4AGidezTfC7XvrdeTBJtYJkygR19Lik8yp
XHRgt4riquI4QcBBGAhhSpHwGZTFhxWkky3cGPQvJh0Bq+wjhDcmtm89sgYaZ1bB
oWXLNGWO5z747Dx7/NKr2f0p1u8zqsxyJLUBAFgXKPwFiYYEtruVWfQgajpMFlml
a9D1kvRbVWmz6Gpo9dmfjOd7iiQldFwrnIpw401bjuVNkG+XR6DmSS1wyVOORk21
NDkQ8FwcI3/7+dsMbk/vgBDEnRvv7LW7kIg/y8cqwahnRBXhnU4D2jldbYw6NJ8j
vaYwG+Jm6pbLE8OfZllGU+637wYafsqCtewB7llWIvf0WV1lwTjiPM4SOdwX5bcr
Jg8ZtZ3dbQjHK+PcuNwAXoYLrMZ/yp9SN8xuzvxILdHwId5+HIeZ6aDfy6Qf6MPx
5NgCHkuvWMDmWZNO5F2T5MTQLvMME0Zk9AQYDRf2BPpqdzf90fwW4Gjm06dqFj/B
cieplDANbpYXsY/D7WUkIySFV+Q83n8H6CD/PbI64OsNm31pBX3IqQH4XA04N/mO
Zya+DuocOjwLQOpwvo5cil4cTRv/eTu+QhsmTQGVxzlEObY7cMPDrXGMWz5YaXxx
v1X++FMEbdzEtzJgN1axA0TsGfazCE/W//37yqHEcwsrw1Fy5b1DA3ufl5B1dAhk
eotp/wOSUgqbuPoxGVvfujveYHg07qRi42SdcNZ0vL/XGeJl1EJN+GVlK5lCpd0P
2KfoqLk6EGMj3i5affs6It7WE7HJKs76dPkGD6khiTyPUIq/X0RaLntjtRbdBymF
isZhM/GrDbXZ5nSWw2mbgXkh0IjaONttdK1hSRAPNEQ9UQyFLxmUOW1JbO7BOlyO
ECFpkuJWD7+Sq//IbGQauBAj6e/wu3a8c4Vg06kVo5nDJcMZ0LF9J1G3QU2D7REo
cLju1SDMl7/YSlea7ZGgCHhGKe6jICb3ZtwxZfFOCvIrQMO9C0PQDhtK5VEgyPnI
uvrRQ0fYv54/3U3oHd1KF16DagoB0xBV1trchnbjDVzKXyV1c491qhkclgHF2aEn
fIi0qabOk6NIybt+/R28YAZlt1ztAgbmYez1Ugb2R9kfkwuGbdyOrhE/Q0V1pfmz
y/9brHU+d433U94qNwr+cb/kbU6lA1bEkaOyYyi5mYpCmJPPkblw3qV75VTuSQZj
BGPuIEm8GTUrkNm9CrQoEtLFI/LdX4PuPOpCougZUOowHAlDsH3H8SCkyYmaN+Zk
XHmZQT2lLY/BxhVdmLuvL4vtFbEoidimX3y4l3WcyEffs0tSI9GIPk0CsdN0neuK
HkkcDLxo93hBz8h1QjLHcqj2U/k8/cNAMGe9j+2dTdl2BwhL1XTfExoddtAtft9t
hSYjJviWx466Bp7BJnC2n+xp+04EreZY239aOtQmbesZfaTc5IXELJLGK7DfXOD7
rNXM9D0Zypg0a0ho7uwP2w0uRCaTR03KIJdFu0dfnVsn6FJy2relYo2nGwLKTUHU
tzE1Ew4mN92eOrbZq4Zk7Us46mGJWXd6PjN1q16aV/PeAQgZxy/DYxH8P0QLu1Lv
ar2O+IBhKdkwTHWL5DHhNuPwpw1F0RIstMPw12Z1shY+f9BpIsIjOQL9C/inq4gV
bvYWSblPxdiwGvs/47LlnK8Ggk/OrHocuY6lPjS7QV7u637rNktGpUXIDY3XYoWo
Dm4qwOWzoIIqFITB2Xdtd7Uswlg4uTkOYH0JEyahe9316WY7a/91gxkni9vctbt7
m9miyYQx8F9kwAhJdz39e//AQFSoweT8jwNPeZghrlV0UlwK3VQERNXfqvRfJzeJ
M1zVbeb+NEodiufHrD6PG31ot/6pRhVjTG6d/FcwWyHxOCOHU/UQTNkg07iSeSAr
Uq5K6ahAkpsi+xHwNMLVmpNr2P8A4IeqTHJZ2o8T/etF73mwwBFd+H8Tulf4uMIX
mGKTTQrw6YdZEC1IPGtSB2PJDJ3awC11vAjSDepZSTYKcEuG9B4Tsg+P8/Em9lAB
gap/XvwulNDFQhSLIlZ3QsE52FibXUaw6LPXLVgmQwXyAhlsqaDVR19mP5jlBIvE
JYNkIfxAGk8eg2FXlnox2VuofgVTzsfvrLqD9WMsWTB4FNCWyEZeFxN3/FRKl6UM
tE5paati9HerrkjGgQANn4m7ufRSPgXq+cKWCAbnblCLGRairk4eSOOQbxLYeRrJ
4miLO3ZRqOIdca6uQ+EWywX28ssyKOCItR+Fq3aswnIpGj32nCZ9QmljQV0hMti+
Iu3AYKJ0WUNFp35y2WksIaq7u5cKbmzQzAlB+y29kzXfnLnqWVY2dZUMqEqZZigH
U4pK3Da1ytILZ4ueDkcPwVpkeZIyNvxPbUMmYIHH0hRJTFHjqRoWvHuci9LtPeC2
e8r6vByG/8zitt0UenIcHkhsYV6Ynh4LQAboJG9+cpRb7OQiHBXuERz26YbmfdzH
37OuDpjaS+wtShJPZfUHzWXaxmk4YNWV78lHkjhOpYKLWI8A5jB8/fWArk+nM4FP
Sum7dWPt7c/iyHAkZAC8J+ioQb960nh+ugItspL1aAZizo5sQvSwDmxO1PcIB5yb
tX9VcoyGBF60afwLl+6/T0dc4CChiGMDqDMU2E2TW6qjA6Gqgx35EeHTWTKC26Rv
FGis24WLM/pgipK281V8h8/1PdJjE3XWILeD4iSiEbWD/7A3qE7MTLDV3bGh5RRm
FBmU5v3qfu4ZEvC5RVJeIv5+x5oS+wCbqEtcyZi38BmAfeXozjbqr0aRESo/1/8t
ySB+YgDLCTSZrlptgWdTboKHA5ov+FZ7NgiJtryc8WAylZ7quFRAE5Gl1m2kQxLd
1a4cgRfB0D24FGzlgYK55YxCMZBP884NbR8d8+ut3OSJoVExS+8BRTeUwRx5eHVK
ow7bZRO/en4kycvpYj1kF/Izbn5Pq+sMT2RM/eI3wTuBZZHuvChp7cUmnCNO/DB3
QQoPv4j+vYwx3JGvAlKYjNcEialk82HvWt5nLQ67bgBMxd72HX8p7L99oIQcg/tW
wuwZ6nRQbEIGzuyzsWrOh/5UeQivkYxr+HmiPXSdCf55sa4WEqO/zdap6c9uy0CW
jmZ2+IquIwuwm6P00gr9qFW6an6ev7Hw93W7R+xhqyD4tcC1dXgNIoGHccT6IjCz
ah+tJu+n7uh0GKQZbsz3NxK8RnjZagaKdvNy09MoOcPgxe1Seu2UUdc8j1wShsMf
iSgqIvhowx7lVI+V9CeNNnKdnwfldrokfsKFcRdtyXNnqKfeSygGMrCxhsxmSzLI
FAQBt73qZ5h8alODoO8R9p6u/3DsIjhy5c8o5DS75WAS2UarzFIBkgLAz8L650pu
tbEfwGahB0TLVo2v5/MBi9SLFa6j5izK9HRK5Rvyio6poXQn8Aq6jCYH/E8Sc2it
8b+vSOmeQwPu0YtRY+jWJBGoNSudcFdmvKnBp9ARiaOxsGM9/NgjjJA80YKNj+1u
1sLU+urIFPRogBrlG4UO4dnImXDHdq3MaLx/hjo5EGY+lO9IvkAUOwm8KKWmKKyk
BCxrPk+vd0VjRTZW+aynFliZ8eMKfpRg8UL35R/p4n8WkJQnW3S12w8hgPpFzey5
RQS7PyblGaKlw3UaZkXpQY7eKU42Ynw9va2AuPpD5o24TmQHG74prX43OcSCqQnj
xE7Ja1Q/AEYN/q5D7J/D6aQ6rJlgmC4n4APVOUEatag8Sz9nLYZkeVMHxfaQjRFE
XUtSTLAHGlS6OJcgq3nhYEcHKZFW4wkp/g6xw32SdYaXj8s0gtXkNUZNqIT3OrZb
RBKC8aD+3aIAnWFaTR6XguVZwq3WUulcwx87BVP1VcVTHbfglwmEXUIMOhvKmw08
u/mSnNhpcKhTNZVjSG7LiB+E3T4iVeAbQPixOoZhMumedako6CepasCkVZ9cQuL2
9JITbieSyKpbzfq3yLx+ynEXBWUoDTO6DuoYQNrv6WuEH1z8yQLo/uvTUV9jGTPn
v8R3ergBxoEcEVAQx1IIeeELh9BKK6lyJy/L4v5mQ90iEoZFMm+kQcXRF8gG6yui
oAGUDDjk1ErBPDveIbdsROPUL7XT2cjo1WW+Q6baE2kyWxPwwgMdf7m6+VCaCKgi
4hKJHrOLxitvRR6KBfc5X7zGgSC955YwXxbqS9uBme88JH3o9BqLrYEBdG8N3Vg/
sUqHTj5wUDb9pwWnai0i4nbe2tkR41znZ6gnjhTZzVZBskqfRZCQieCPNBK2n6jB
D3blGzZYokl1OlDpQXWF6rRWN6vlVQS2bmOGDZ+UcKvy0i0AsgO8rxdAUudEjZsO
2bqmr5IVGpkjPr2y6OpdREZtYFmuv8hq5Wp+TUvB57Elkh2f3JmR126miV4iU2RD
ckpkSe5WWLsIEBMjm3x15Sv+tF32oJAoVn/t231CCoaAbrFI2ZuyzBfh0M+9ugfa
sP2QBKhNOzubBQpj9ensKg8Dn4tkTQHkPDCOIFjf8gRyLl9jj37LLiR/a0wLIusx
DYkot8KX5+DI6PeJqempvSOwR4a7ef4uVfqfOgJehz6CGrNwS53N53dKCq8t2eAl
OtNdl9MvUteCtufHJ3ZCJGNosaudpm8F9vzy0OBxslGnXma/Z3wpIOHgxRsSjdMJ
DB+sb1bggo5xdGx9jyQe3Rdn/MaDYc4M2fwM/Ahe+fs3z+G23VhyZmfGnJDmuThK
x4G0J4nQxkHmSN2VF85dHcxvXeueBKKlXC9YsMDXVYv5pZeFizMReD7fBJhmI/If
Nf15cilxytMjxgkwU3dDi16JFhIHqc9qO3S1GmvqtSKEKjAiXcYxuYgc38Sxz0ND
RfInFNq2FZszoudd2z0iGpLKBIJAcNI9EuSY5eQBPTEJDnBfH2l/85wuDHjS6k3y
9XzzRWSyTBzi5kG5ADfGG+fqjyK8jAeq2dkj7/Y1BYjMkccISKhXZmg/4r04riMu
KVOlgtOPPCx/HFyAkHRmaUbKxdG8iNdgoE3ISfKdy8MEXunsC7W+uR/oEqHezKN6
BZYBCtC8dxRKrDz5vD9pHuc4qVjwOsTsQaveQWFK8jgPSVKzZfWwarwm1433nUQq
1sWlBt4TdMOzpo9+czN3EON9HmeBPKqVj3Hu4OuvN9fHdso/gGhdNW64+ROUHPfN
E5mr6MuhN/r9Bh5HIOFzLyVzk1vrIxe74RwvHuLvOW7mHtT5qexuJnl8+zvVxnM7
VnMBX+ximRN3B7i5lNxOyboUGDNZRuPmmaz+JN3UTbcZ8DUlC0Xd0G6Ass5Gcggk
AXvp/DWW3wOpQthusS01rzawRZpW4meLueE5ijNqvihSFPTJQFVRYjkr4OXR2tQf
jEZltcx8g0gbTwn/x6HGltTXYwMnIWe1oezWlKe47O4UfZ36VVrLglwnbnb/mvJ5
ZBqHNLzkR2hLi3eR75DYFcDE9PP7dGA7YHc42FLsGUqHRgHJyxHdnTE0ZFuT/5Fz
Te59MJIRG0nl2pTI3DPpJeOv//OImiLjmCpCdwqasW/K7I6mDd1LdjclFBvf80Gi
aTLMt4aHhZ6CsjucANnvYygPFGn70awvlBaN0gaOJzCePfvLaRqIjEX9kctvEaHZ
A3BY2mvs0dSAA4kO1mI9k8qzo20yFUo1W/u0ktgE64gmCisO4QABC2AhPPnCQVXB
pas1L7p+/+BvcQ/yJitpG/dZyCP/0Wu7/8xqwZ1UX5cm7pFEHei1KypHIV5krwc7
4vSOTCkZs1rzW1cffJgZQgvnFnCaRV8u/DAJgBIM6v7fVpiqOPntM0KEfnWK4GWp
HWTMvC6iRdkAXhKYZfIr17N0/Vkj5wJ8X4maDw2sGh3dWXtw81JvWBpY44NWrG39
4C4uF+eUKelAKeCu3kIJk9IE4+TbeSqd2DkxkRD6WNRPXmdmr0CZWgBT+Kecw+k3
O1BqdjJ0aNIAnarcjhL5z3iX5aIuO7nI3hA0RQWwMYKWw+qJUhb93jnQa1ZYupJb
7NRhxS+RitLeETrnb0ZsLL0h4Hrc7kXt+QlAiKHv3cU9du1doyZ8b8rCvViB/P5n
lOLAtiANmX0BlTkWxi8tWjxZA9qc9j358ihTAfI4uhOjjCZylx6SXtx8TrIH/ZXM
zjDduu5x4n1bBNd2H38voDW1BRipX95GRh0tCBYAFPpK0QY4S6y7WT6lzTol2q8y
ZulFQateEdd4NkzV+BNqO5fkHXRyvbwE4a9riIg/t/BZT/Y2nH2TVKoPKLwA3go8
qWQrViYpnpoHpdmknySrRfGImCDzD1qD8S2+8fIbVrFA4Lfcss7DireMaLdpSJ6d
6lU+pu4L0UW7juIj4loYp30In8ZuJzapjoJZU2qUDBkYjf2fcugDWUlVhZSQYYXT
GvCooAzrSrFSQC4Fikcc2uCQ7IH2aOhQSJIGzS3fs2FF36fEqEX2oQkedXbllImB
zxFjc8NnRPp187Y7EMtQeTW1/lVawBF89aa5fK/Gdr6/y69Air2E9uUcbk6abjW/
4sCbOxKsfVGbibKd7WNEHn4KT1Mb4Vo9G4Y6Rrj23O4AvwowOwkGQ0MlVehYbgqR
nCCzt2fzmSfkvM4d9cm4jZoQw71WqrH/zKFpAq/UtF6pn3ULPTONbC6A+K4Hy30m
IMkx/tJm8b7A4DFfMZKWAvreqelBUtdKkEj8VqYWRb4p0Kx8fq/S2+45JSLLq59v
xy9OVn6Ne4fuusJVcPpi9INR01U+N+cklquGFLPPAwg7ZtGfvtt20P+A5tTcPw4l
Yi3wJnvJyWfGLEcytkD99PJai8kOFuXDF9uhn7mO9QP6IMIpOKWWzMnvY53PvaPd
mLIuTnDtag7Xp1aI7lzf3aO4GriRQB6Yg/ftf9P83/Zdys6HNITOPTzx5dC0eKbp
/thmalbE+lPgOeLCgbG9jby9B+oY9Ss8jG7gCbcTbAh7N7eNAIz5tPu3T5QwG9oA
5PMPf+n4MsYt3x1p+x8AJfGRxCnPYiDQqj804HgkHtI/Fs+4p2fo421b+7JPpMX+
+YESzaPzuyl3kair9tqTbVf8+JlTySK8cXhKU//fU86Yzk7/N35evQ4u7d5EsaVT
G7IWNvS9LJxgkMiNBATViIreXZqU3nIP9rJA7E5e9v9efMfkAZxvgDeM3K61ja0H
ExlM+br01d6ancUISd8Fu2zYYGA+RSV6KXL9llPwB8VGXObbkML/OQEzxLg6QNQ0
Phl4MeUCZdBFvgLZI5I/oaYPGsx4lUm8Mac+ZDOjOTh6Y98Zv75ecCq6HOif9rtk
7ELMR9BIlGTWF1SoxaL2ahaRTdoc7JyGG3ridJCTDfAdXrBfezObJjoPBBIf7qnW
3/Z1NwMl0c+k9cb6cKOMNqTp4ZLXcQbK+XgLyG5I/7EY/btkjY6PeWXZo7ArGtY/
hgbncfLGlmsQQyWGuHaeLkaXhFLReSnQDilBa7+XIs/ehTEVMEa6LgbdNbSj6EgD
7cSbMVvFwodE1L3NKA/84Xi1VmPAk/uAp+tsOKXImZIBg1cJS+Fp55OmKqi8lI2C
JQ+CUX5HAZrXUC31z1kdtZQi5UoU8tH7iTt8akMrGBzcQiNLQTKVKsIj5wNS8g6q
9ctonJeiH+ESiRGDXY9khyp5R2vvRvJTNCZdyB2AqRHiQgx2qyFTaE/LlNliLWK1
QDua2esmCfuQ8M5q640ADVcy5jbkP0t2m8pdtIGrPi7t2eBMl5oYi0dIxtjZlga6
iM0x5yQS9M1yBbewJKxRN9SrUXrMUWCXW05Nk7biO6VNwdjveYJKQwoQrEvNyiPX
3vaKrP0sTlSg0x5NiCV0VztniYtgRk8ZVpR0N8UaJ1y0A4gc9tPccLSeSoTwrp5S
18L/bYcd6t7MeUo2NR8FzkqTog/4ImdsLrSdwl+AmdniVu2R+ljQm+FtkuNb23wd
pYl6KvAX/4duFcbQDkXkNo6/KU3+V0aPiSxnAFVEehBwxzR0oVNv8i5R9O9b6rqF
/Wt9O6l9lz+UwiCDlmHXCsFnaEwvk6shfKTdMypimyoqG1XTVYpvA0gMH/MmUy0+
zuwJV4bZktHfvlEtprigGb9Ltz1re7XP3G+RH4q5YXosO1Jv83/3bqOJVvpTT3UV
OCEPj9ueXGaQJWspnWtfzHDbYFrn9D/NNsrLw2JOFOcGrAXevsPAjicbfWmAHZki
uwQep7LGBCduQgRMHhbkhbye3gLyfexJpKHvtt0OutFhSBtZfoqyvtx+LmIzXTHI
24vQjzrLcPzgD8LtXdUSB8p0FN+BXc55XJuv7vcLqj6ERjI3/+SXylTlEibls5C+
nIYqlqo6eGV+F7xKptH1ukOK4X3trQZsobXRfeT7cqLjkQjFm5EOItaf9dErxNn/
JbgYTgrOHh67wWtHxRvPA+tYDKiy8DelPhiZl1+6xSwvDRHyqSAglQed8mfjlYGi
z7QqSehtnWeMmpKnTKI4QcaTQJtEj4QXcezM+384fGYBCNX4bHoTAYuI7q2SrcSD
AmEMoAc7dR1Jc07Mo1nfGrA2/Du4UTbJWzslqkPjWo/E59IsIVhE2uxnJkBVE1hM
xJQwowJ608SRgfzTZLNGm7oJlZRPCDX8IcJbqV4bDz/XAvcWoiqJm8aCUPnzQwX6
swszrcYtDBq+TrFh8oZIKSS1UlEEDywUCvi85nI57mxL+007FM5DG3jo00+oB5Nh
jqUR1ZUrEdbmdm7PULFCaXpB8B+BNEDQR6NJlmSbdKgGBjp7nV2J+LnfXkS4NvrD
mwn6TfEQbJpv3/2NSj+cGp2Q9d3R0aj42Oeb4Lc7M5C2H025kIWhjk8oRl8GFwJP
XywRgJthfaqkg7rPZ+4JHWHbFujQ9ZjH5oNHoJmTLqPb1dfRFWPpNGDvoZluiUQ4
UumpK2xD6E8M/KVA8b7QdXIxpCms5ceLHc35GVm9JNyN2EFyvUvQ9LRts6W3+d4N
UHicHnlbu8wt2uvoAlDQlomVEL7UlCCtnsanOgi4/6fBirSaTRVDdfkLdeE0dKJI
HMpmMUdd9ab09piwa5QibJjwWYDcvzJ0XBeKD0uc/tJNRnHIdKMslT6fqOUvTaQY
neQWPEv6OmTRDW6gcuWQn5yfNAGrMQRAmEube6W//f3yjUOwmuVcS0XuPPA1GlVu
6GwJfBZ/Ulwr6hKwFZ69DzMu0hpGM74V67gA+k0uAH3SKFNtv1Dr0ucSYXjbKBWX
txWm/3De2PHqC32lIL7kT/jF1bM7Brn52MeLbUcq/AAsk0QEBdItiQti/a35d2KY
dtKk6nGtR81vR5+qlo592no49YVbOGAZI4VJU85WRorz0xbWmVoUsKzb6SosC0Fm
+mBqL+AqdWVnT1ug2sbGtdmBCg3bOW4TM70mYfRfp6s2cEK5XN+tZcsQwrJTFfc8
Lje3Si17u57cGrAPvOG8kABs9qbltSllOu2BGq7if2l809lwprB3MYEdBijrHV3A
bGm0HLCi8lxZfnABvRuRTPD5aAdNnEljXdhJMFbI9YrFSSgooRxdOuRBAOZOJXBS
JDPWiPkkh4dLuH3ymM9ehIHEx4OYYnCXZBoDH6wsBv4fX8n5HaKcpXeJdsz2fnSX
Ia1NCkA+altoo9r6AGvo2gueD9KO8sDxqmvfxgHuUICcx7wY+KVUW1c8fpA6r4l3
PyXj2cQf9s74D0zIpN0MFKwqT2SgPhtFVRjxKcoDsckLz87gwA2dziJ8Z1lJZbtG
+O3NigAMCrFwVJ6wpgYU9p+6b4kTFuh2nsscIqw0jMPTPuYjKE8KPyPm9IUuhwYV
w2v4zIW3cOf8Zd/j+fS+3R3Lca7XStZXlJRryt2z8NeJwIPKvfdOs/5FHPYM16pF
qist6eBHG+sifWLXMSlV3Cd5cmMe5KdDcfMxT5G14Ay07T5lgskRQ6139uoVJo8Y
OCQeFOEDo0aVJ0/SvQMal5fnUTtx/8/qqOl2XgCJf54AeXw5cGdAPadkju0/Y8hz
FA1tqPlRdvorIHwtGYeZlCCQO7KwYlNlt2/30BqSLR6tCGTafInGnPD2KZcu0i3y
JmbNHeKgFw1utzt/IuSYK3FC/KnWieq5SWkaB1fymRq9IhjvxauNLtz9XYtjB2B5
+cWwfrbFVAkiZlvI4L8fNg8FYLrLwvOcW9Jfesbh+ds8TmorFzGGHX5LFSlUlWWa
T3dQAkXfGzdnUzhip8Uwd4SUN5goATpVwZYc6UmrUX/UhyrbKBUzC4L4tyrcHH/c
TttcBGlnS6WlbXgCq4+if1AH8rVn7dhLvL22NJZuH7Jzq+4RJ8KGRvwqKSzc5t+S
3Hk2jWVGfB16TK8E8gzKXSQntfzAYhOWwuJCMxh0XsTXGqJJSnfpaQiWQ5IrEZRd
iTaW7nL8xuLVuXuWq3jE3BZodpWUtPfBB6ftr6FNysqDoW6tFxv3XzmR8Je7y7MJ
2I6QJASMtk4CiYwqUZeCqd3//GJXGv7rMg9IDgk/mmvtTNPmxYj/xd53qSHmIBKx
j2+vJ4S5qW9OrO3eN4MVr2h/nP0uWkERx98D+G9YtxQNHFTkRzqRRLBq+oj8PN96
2f0lUrmvJWqHfSf0YPvgSjp8RnF6/DWLgFqFkFtrq2o7YwfRHifaHc2KWnNnlH4l
Uel5WZJrXHrY/gOrcJsLlFlssMSflhRxd205sX3iKfSw0USVgMgn27V+ZwPRfDZG
3zh71rDaHSTvc3b+RzPtnRLM1l9i6qyKnD2Z/8EOx+YopfhbjHwXX5he8vdohZ+5
/ePDhGpiTp3sQlPKTJPt6y7pHD4QhTitQskA2pte5RVzTBrO6bvRLisLfMNzWmwj
uuL2whVIDxdbI+liJYc94oNU9MUZaywYzJnyZOLrxnEUY+W4b0U0V2mvJUQ8Cop6
xJoL3sHe0dsumOHiw3PZ0CCV4gwmSyufcZ8ep6Rys4PAIG0htLDtuUpBvoKqyO5E
xM1MPpwG01KDjD4Wmqr7wyMnvWBzZx7pIjiKFM9Qq/oipqfJrlwBlA42df3PM1Wa
VjoB6AH4hs+gzZMMtEAFxclHaHKPU3+RXtXlNN6di0QVCw/zR1hRZN8z+DhHXuLb
OV6Dh5TYhj+eQzeSjqUtG5hZ9p9CC64vSD0VbfDbV0x/evjfIVkKSG35fSdxpmD7
bdhcVfVfOkjLm35nxGBnP2R3lVRsXbmFKWMzIirkNY7xDy4rxlp7ZcUaPllr23uK
us37WuYKTtJxyZJRavXeU/W/P3WYXipT4cSmoVsbWPiyopiXsXuEvLcZmsDuQ5XX
mJ4DADWgXw5RDseBxMDUavi10tS0c5KVFG007Ix4v9A4P3QmbKSsL6S8/fzFuYJw
DkA5cpSjiawxykgmkV2ua3xfi0KDoQuSDhYQc6Py1fw24vHhLHcbllDsLlkaTJxu
ZjuHZT60AIrm3aDfM7N9OK3DQyoibQBLf3pig2E1VApOa66ycengA+q1zDGSmMwu
kXcP8sAwt5r3xlnwM1SUO5TkdK5IhV1LM5V/LU13OFclXaDYa0VIZ7zn83PpA/ga
344hWf/pcg5zq8bwxy+no833ywUGkb9L/k/tH4XIHdu46dj8flTSa0zL8PCxl+EE
HBHbvo3Bbv53HxMkLzqLRTSrhNVTwvJPMcHF57jQbjc/8KYRA9b7gRYu/G5LJB74
B91t2mXkuO8KJHjAqOMI/e/z4w6vAp2xFuHn0tUj4i+2888PmwbFRPsmuusqTIIY
bSTv+xmKGpm+G0o2edRFCf9KOG0l0LP1AJwqAPGlADIa9v+OmlFck3EncRavFQB8
Oq597bYaqEYWrOeDWOgx1YCHLkicoR3uwAvrlvca1Ardz0uRGfmNWiwXZ0FftGHB
AEJjQFCgu4EieYfc/pl6kUZKlPt/FHFcYUUHM9ItRXMegy4DJt5SqnleT7D1iLNw
9t0yJclaxP7idqTbZZtZMw6IjVNnRun0Cej2yA6VEgrLHUNYu6CyAadVp4IBdRLR
U41f6jHZ355xph33Jj2ixsnSfz4/DM2WSapLRLACKlhahQei5J4TWTyY3RvKWxr1
s+kLp5HZ+4aCMEaT18dg9BemeOwlG0bqTvndEtKKc52j6rxSXULTAfXAUOA/giGa
ks4SupnSETdlT3KBAK6ogitrwlSNs3lEmIIKfJ9A40x+k5wg9A6tqxFDjLAb2bnC
nkyzyxwXLEZbrNQXjYZ4ORLeazr9r5rQOQ+URHDUSU0v0XxT/iSUR/fxH0xLm/kq
1SQp2qS7hupR2tFX7BlOrbGqrUULjptzHM7eGIffGcqHGMlMtxE0xPENFIbRsCy2
K9oJgr1jICzEnMhdLKS3EsFiPVuM9QjaFiv104UtEt+2zx8LqEhuPKIyI2/EUkpN
8qwREbAVGmq7m44vGYW3ndQnFQV0niZxzDF2WUtfE3nM9OloA6enwyA2ouEntUxy
oppkcoqcF8x0aws1csO+Qwv0Y4GIUHVg0QXLP9ecCHjDBzecXvWJWg0Y2Dhpfjpk
T9NuWUclTus4sOYBvAWlXjrY/gQi8looXNsqNmF0ArQKr7J4dqcPmk4MT1jYLk0w
xvA1AGxLpggccjNGWzeXMVH5tcA7qi4+tq5wPbJMkAVtsWbdIIPCpdV6sDr5GuLX
zKnbqg1a+9ZrTMUYA6ykPxJ1g/jU+iEh/L3YYixitkof5uRSxbzEbmSqLzzkKgc7
9wFOnvTNfDlvW0dCDNe2dNCH3IbKojGL3QIzUIe+o6n/fwF15T+71FzJFmFYfteR
DL76hI3uFDoS8FZJLu/ky5Bc8anHrx5UQjvEGNGvQOF1BIFlY04ZGQGeZCDQqyxo
9tDUHgH/0sChkeZzkRJdzPOssVJsh03kyx1jVK0GabKEmM2D1p2FPzWWozoqCZ9s
DjB+as/VAdjWNoIrEoGKIjijk1v9+JRDjGnriIRpsRd3u45MQ9lTIaclr4vvc8Gn
aoGDnAaNnzXy5xi+Y5c/fVo1l+8E4kdEXwenH+EIWN37OiLM1SaltMSm0iWgEln4
XtYZ1d0jm2bIHtN02j7JzPfiindNeIoPLAZlhSv0ku3A5zgHDuKazWL1pN+UiV6S
ZIOjNiFdwOjO7BqJd3fPtTFzJ8QBWLFgY+2YINjnxbC3abu8klvMoLWApQ+yQghI
YtWl7LTbJQOicD0rlx0smkQSPoRphecyA7TsWQ0C1HbSxnSoGlbZDzR78p53t9Ap
dBlVd4I8cqmkIofaN2tvR3puUPYJvzqsEAIkmHtV0wrsMRI0axn0tinVWUg4cTfq
Z29R9Z3Iz5nApsfzL31gqckk2GD/3JgMhXHzxjTUz3/zMOlBP6LmHcQFdgFxbZbn
IgPgp57kUKZMlPzXKR3eStyX4nPFs4oWtraW1DanJk46leKA9EHw2LADSx1MrRmc
1a9o4cv+O/NrJD80hzjpGYa/rE2oYkjwZ1xxyVOdZqolvR5FeOF/MaymTbcpVcvd
Fjo4CMpfmmukX63wg7CQ0OS6b/l4/PvOOqid//+1XTRuGcTosGwdK19KG1Z5GHwB
VBAPd6HgUFFqAi1oGThi5ZUEkXUem6TdzoxSvQ/t1GhIsNwOg6GUl9mShfKWzMLu
uq/4Gq43h1RosPQwaCZoJXVZRj3qE3zRQcpEGPaPl2CYj32pGF6L08cVDcDl8Nfn
swub/NLu2T5I3FlaLButMOdvbzKYSqC/cPpdP6ef3Cu2pg2tCE23vXwa/MYrS7cx
mjeCOdZ17MTU1XqABXNPqZTeq58qvrUU+bWqg8+P9zBieKIiervbwrxKvEaMw8Qu
mE3lcI3OKlBQDahQAsUI/nl7WxqxhvS7ZmBHzdZGwjdcLCGFWOle4yxPHdPDzEbD
DlZa+n5EYCer2Ab1v5v72lC6xWgHRdoGnereQQs0Eomgvbpa31W7RX4z2+jZ5c4R
Fc1g+y9D0ZaVJpqB2TcxniUYM1lEv+m9k35DiIn73w4nNJ+TR3jy9t6D+/lzfPU8
bdby6Td6HHmADw2imiS7Rl5UgVV5GetBOQ0YYHXSRAdKjYc521+mtoETbPIcxewz
Z1IxoGWtkCkp4x97aecvFwSsSpKuEEc0KQr99qoJOHmFFDKk3MFfutn/a0G7oRxS
XzoN74jNE8FUybBCw6oPWqWIhogEmfMen/VFEGO1ypxU5wey07B0AEz/0fIfCPAN
+wWnmcmfzh8RZG3WWki2FjcGttOhZaE4sdqDuk4NhCyJbytBaBbGnmv7aZjksYYi
Yz4y+z8Vr7P/00VVJwCJbotrUQFxeV4Ks840eJ0p7ikHwuGstcnb477ZigNTKZFF
HxtU5Q8bnQZ/opzcKxqTYV0RF1MGqu/GC46llphPXhWPGkj/aNZqU+Wfo1EDqtKF
J2k09AJWIHQ4aDHG/SGxxMbLENd1f433LxnqsXEMb81d3jhUiwgqOcc/3nnhYDaE
c8hUVPaDR1kkoikurcPrtlVU2IxKgprrx0SHZjkP/eJrf62aRmC6sTbBivI0fzJT
g8GeT3m00sgGpre0SIeeQVqWhIMZxj2jag9LkQjg+m94cE6NlGr9ksBDU/Z1UVN8
CM/HgiEcIwyUTu5Fpq4Xl/bo5F2WUNMyQSaAvG8uwo62tUODEhubr3v+KEBY4USP
akey5bghA7jpmGbSXrT0wZDoa5uZjiFpRQ6uaowVtvj56brixCsMKNLmlIGcDh0y
UI0eVWrEu9HtipFzKZKoX2uuWWZ2z4ee6Lw73kw8iB85ktUt2ivrv+ij6ekq9bts
v7TiRQYvGJFI07fJhrfy5sUVVKWejXmqcIX8BC1vKvYPqtnISkFbI2CFCqPR3VkU
rdlBCREvbGFe284mLub0UWgCmL80i2J+mS83hM6POVqHYBVEk/JDigitbVCMbflj
RUa36t9opbz47V3HeLpoL6r9Pg81wtrq2pVMpsWIaGT12HT7W3YprKs3tclhMaZd
ljbTYx/2uHeCrPEUqk95ChT7QuVpWhBKUnSDg/jx0v4GyIagn6ZQXba4MUEnMh8x
DUyTvZPc30aZKwdclfsvKRrEfOCTO0t9rBw7B56j2EsN2CLG7HX7EkapSbbZu3cW
ovRYsMYJewWA5Q+FUcpXzkLxijTHzDTYZ6wPJ4vohOf/lOwAMlYJ9ah6PLGvLMa3
ldh2QVuWv0ngKZVl2+yV5eDibHqXBxcAGforLIoM2fngSkr9RAlzlszOIPKbnb3X
OfH1TvbZT0OJWU6rb4YCFbYx9+eiQqGvzYAnpx0OIaVJGtcv0xW4/waWk+zEvRJp
RFc0ZMRzugEK+jjk8RvEeLz5TcYAZM7N8AGxj/DKx9u4esrYmuQN5LAcNXYlQzEf
ojoRMC64yTlgHrAEdmZ0KwZoD99BMdMVPD3rXMtF8savlLC147aTv7PbOpi5fsuH
1420kBhz4uYY4r9a27xlLZBrUL/GkTGGTYHi0sws1iktcpVNySWiERyA/VTkw5ry
osNbP30c2LTgx1AHrY0Z65jH57GyPwsFNe2v/9Rv5/CjlG13nvrzbvNZUNP5gVTh
uuPaIkFrDSN3yuwlMhpxfeO+3graEqWSQBgOct1w+S6+m5ppgt75xAnhI4RJ+bla
dG8L6fsmhctNyb0TOxa6JoTB5SWEpAcLS8yMMn44o10Ojq/dTHW+Mq++8Xelb4NL
0Enrc3RUtc7+L41joTDAYVLa8pe1g6+q6zHoDmlfTEfrAZvk/iB0QSgHmJiHzfTp
W6UD9jS5Fpbljx2zWgodEwLGeIP3K+S6T0AztJCd1Hyh/t31qz6NdexhLIc+j2th
Yed6FF/fFXOshEVlcRBqVZjCLi8f04HlomicNCebbEV2jXhDEKVfRlHeA/OWpU1f
iDiBkWrhJ5fmx/KVGxvclhDr8enBIN7CNcGTmiA+SwazV5LrK54Vl3zACohflf/O
wOzSgyYw9SR22cFUDkxqJKWLZaZeJzplqSgNJzrSga5qXvA2mkjrz++MkWIK263F
m8QJS/lhKJgKHFeBmAVDEQBlzlyfc3xqYPSssQWabnPkeczhcpgCk5EPXLAImger
uWnAEpKd24Q6NLZQLh22CLw1cEympp8D2KPXcwN8vonKOzZKca/vVthzE0R6Jwy7
+jvDRi0YG9rH+IG7rUjwXYTtCTYSho4j/jevzYQ4B4UpWFCLJ7VlSinDYaoekndE
hkTToQaPeqP7e7gukyqq76zfVdekxbHW4cT3aa8+BlCey21/3Gs6tetneDvwv46C
eznmj2NA4cEwyJ4EWaTAXvcPEE4kuTA0OhzZZ58M9Oj648yVvvqyWblx9+nS0zOf
EPag25uzJCNLxW8k9OaGPDAJRpIrfr18616TZJkvyHN47GifdngF6Mmb+uf6GP/K
CQrwLZHpG/x5cVnhNnCi/6ZoM+pu2uA0YL+akCj54M+Q3v421MTe7lyKNalQ+73n
x7Bp3MGVscoD4zRhGF2vlSk4XVCQqViuOdndwVu6aZ9tnLTYcaTG3np8yWMCqbR6
ALW+gHd/7s+YVV5pE5ZeOL7sMiGhd+cMargwBCqWyX+0NFU0lfly5SzgA/yluD/1
GotEzcSgeZx23713tGFCSW/XAgJDgXrAGz2YdwEAI2rsX08xC7/kfbHkSs2e1iD4
F4JboanW2LbnjTQjyH1vblPXKs0tqubg80/Gwtvm7dekzqr8EN/tnBiSFCQ7ZYCl
lOvHsFuLvE4H80vOMt90Y7BH1BRTnoDmse5fi0kJLnS82l/+n1K9cQawYo31l+L6
FNSsdRvIDTP+kwryRnTuqNN1z96fK2rrmcpdw2QtRquf2lFAldmZpVTj0HxuujT2
OpiYaI+v4OyUJjB0ImFTEC7+rYjpahxVoBPL15iSUn9rOMzxbqGjLuzKnmS4s388
RsR540r4yDtEPAW1AvYQTzzUw1+qW0PxsngCnVbDSupNwQu54N2iZsnT2ypPRCYL
ATlEjCfrXji46B2+2X+mM9rTyU5LgNm3EyElo641jBWMKOsefgYGnZGn3vFQlp3s
d+wXU4eSnQ4nuJ8ShrsGfBQ877jYRtys93YqqTnX+nHvhmLXnyi9NCN4GHx8b4BC
qyaRmmRwjn2buaQt9PMJgbnhGFclxxXP058/MUJ3zOTbNqN4rSG6kD2UH7QASV7y
Lbj39pbjjQwFlwC17u6+NHLiZvXiwkC/Oqe+jk0C4Dqo0oq6eSGFKvK9LyWsySj3
A00y8M+3x2ctipQwSJD5M50D0OlJBsTfNbMtTUnVQQRtsC2no57fCHeB7AeoGY9L
jtbffzNSD1h9q3w0poqTyyVahRuTziQtOykduASvVHMt8LNE8YM50d+2UkpTgh8X
QGrhCO2/50RKmzWkPkyJ/Utx2Kjlm6T2TpwVSMknuQl471Ann1LXI53IOPVCCN0y
KSd9wCySGSedmkoJMFNsbTDBWMXZfm6V0aWp5uJpsmaEKiAo8q1F/Ikw7grFqll5
rM8npQ5CgqeV9oQXm7EHBDZmUjhk5qno+QMv+92xiQQlQZSDG9t92ju47KmxCseq
a1evoD/L9pcrDA2UFOp2k/iWTIEQTR2nuPKQA3v3Y7iuz3sP+JJFcFPoYAioKjs+
lVCzTfcqgRIiCm4keKxu49g2g/5r12WcoShrcEMZjY04W1Rrdt34lWYq+VQjUYtl
M1OAgD5dpHdp1fzIsMdSBsYZj1K1EDWXmkPFSiLuBqfwANQ91TH2GCYdu6tDR5Y0
o8WevNa6ZEOV7VRFTKhJNQvzWyB4hKo4Jb7tQllUtKBYesN/hqkSYj7yrdcidlUK
YrNS324nIzjhjXMUype9JZXtpKWDBfWUNi7uQXzFKcelOmjTOgybN09Fu7RSNfF2
j0xWatcb6ldpsLxj8O7tBMuTzpo4eili1gY/ybMQ3NOgU5lmxvVG887HElpTakdP
nxaWUH6TIUpzV51wH1Sr7n0v8G+hxE8YSC3m/NTPg/+pno9iqCZ/7ZyTqpyFKAr3
aG3/cPn4irNTQE3PUK7lMymsxfDzR+3xha7GGqW2GGwvP2yhHxoIeiWfhcCedhrL
/p/ShRP4oYeljmk4v0yqzmuW0WXDsKRK3rTgaz/FLxPTZjFtNjF4YHFiT9lDeIfl
NQ7CkY869UEeOkaRBe6kn5Uh71Dfa4U7qHV3r+LuE49uOPkUYZ5AO7s9Lz3TXNTa
Y7ljmoAsnsTQXka21O+gSdpf0tIqVda1DjeW5I1u0etF7/8tNNm/8j4A+2DF+NxA
4PmbrODhK8gAU5ImijAxT3NZZojYmn36hV9rZaakIOuzzoQ0K18x9vw7mtvZmvzF
MSpfjh5POIXqq8sCUIuFlOeU6/HzmJUPUP4GK+VAA8UGey2AeD33eUhuJjZlYT+w
ntAacLehOre53uYWLy4Kgx+JWgDPy37f7ZAbatPtotLd+t64kYILxA2Cek1wo318
A/8chl3md/j1iaIz+XO/cELH+IVhYqe90Kn6dlq8lQ6RsMfOSA6cgO0DPUSaXWxg
6RRj0ZobWPvNuK2G+tvJzib67Z4ExC1l/3EwQcUQVDkbkgGl8B0lKVABZrNwYRCo
a78+BDTA1J0bhA2NmicnwMxjO/+KEUhVkSmmxn2DkfVwFkKF2r38v4THoNGjkREH
w7EwfoSoCUOopg7glt1oFD389BkkTi8FL9gVnDsK+RmHb26hDl8xRRL3lDn5GKq5
Eh0NawPRbQ6whbuHtwM4lb39foMWqtFOkhY20gJKRsBvlBWc2a34BIDOhzskqtGs
2yz9Cm8c7RJFHlm4jMIJSN+++p59uFlCf7OeuCEnnZ9e+gm6T+xsg15X8JivyTWO
RUC1tPNglH2SWLMVn0gOkGLLG5PKEwXz0cgj75H1IZMAY2fCvoRzj4rtH3e8ABrg
Wbfm7T63V4+8Dfb8dP5yEb+kW8/TZsrXenJdO0QK7RMo02oKRTS7Kw74YEdM8GFX
cL2ftCzcjjU2dktsxkAqGcH0HTqy3aatqUoASjmQ0dwIGLVPA+8Y8MW3gqBkAdYp
fZJnlx2t643v3pTw+3xsSmEbi1Hv46fOz3HZohU4QkTfUwebOU9ZH4rLWCNblXRI
FOV8gYboO6OCmLeJ2p/Z1Z/tG4Rd2jeUhpycjoNCE3bvBi0q/uCgwb+CbVeygYeX
vpgS7rOL3E68MKsCvZhOdQUv7/V+h5+A4oBfynZBbhLut86Qs4WeXpoUG6C31tLi
MjjDCqPpU6gah+x+ss7axWS+akkBs3nJ0O4fqgaAonSlVCofefWsqOen6yjZif1I
NgShMDBppIOzZvz6U+Lxk8kxYq9dC2fUY0VHG5Fq28GF2FMJmQq+eooeWBVU3LQr
ETKxHqGUbVEr/w+R/FOg8nAvoI84k2zJtYJqz9Jmj1RidXFotBcPD22yZ+PCE8eX
y9MWKd6Tng0XPptiVS+zvk4xXXeGEu4mnrdejH9etqf2QszmaSnI4j1iSAoJ1m8l
mw/DnCs2+tmd827CsgGUIr/uIs5oLR2Z7IEBkJ3QXXamMNQOdoDknW0V5WOf6s+D
+Oyz7EkXRQmPEhAGTTkXQTb0OFLki+tN0c4nDEp49EeaOCI9UOPHBXMLGB/2mv+9
zwWVaz6H8EydYtmoQXr+AgBCLrk8p3CP8bkvQfU+ZlvVh6RVScgHMqEYGVWO74UI
86PHIXjgNMR+k+W2qKzRrCRTS3Tn408vefjq3VB652Xc2nKx14cqRD9flSMD8OU7
j9P1kRzDlg7d6o9ORYJ/XBltK8Zm1jScV6UG4dJ16ogY/xz23EMnQdkYLdFSdkoo
G851/4TdAoYemnf3loe2Zfnlra1N4VbvnD2MsZFnyDsLLFUDK+dLTUSpwesG1z70
6G3ColuT7JSPCmK0pJ2BgKdqb7TjB04cIcToj/Be2/lIXkv0ksXnUsoca8hAFkhd
/t/WxxKM3dZhkUmsl2+wlpU9wWcmqEpR1408rOKHVVjFTnLAcfU3jbtBP4+7V0MT
G031QzHPZ9jBak6B5Qagnp1otcFBCuqOaRvSNZpNnACIJ4SMC3xV4XrAtLikWDZw
1jjJcgd+j25ZDFpuGQPVw/oYVfK2egYZjf8g0Plxx1jHQnAWbjUBkWgyXFV1MT3W
O2UqnS8sdBVz2F1uIow1v7ulFDB2y8wQeRB/aqTIuzKfP8jkgWpKs7a+n848NyBV
idwhYry+fb1YmCh3wVFH9Zo++5glnDE5YmsqY1SFY4DSJPZGPKiNBl8hXW7p/KJH
oxg8k/2aW3lYA/Hq1uNNKx+DpSt8lsgWtCSZgrfr2sly7ti5ASj/7Qq8IlUjuPKm
J7PgAAXSW10ya0iQbsI0h9IY0vtZhVxJTOh7udBP+qGPw8Z5g2HYo4mD3fMvp2rI
vknRXKXxGYnigZpGJ8EJ3oVujJTMINdALkECgcsG3xrEoFR7JU8/+tScuokWf0SY
SA0ux3xtN2Wb2WvAi3IvX6e6gdkx54zsw0BE9/3Iq+aWBWWzEtGMPpTJXeM4L1Fl
ejlQvfRfVxqs7kDYuXcC8xAEqZaWW0LXHPF7NL/lsg859KNq0t6Y3SKO6Tx/OgN7
eH9fpIcBEna2JzvzZNnhCVtXIQq+VOd21RWD4LdjZrJAdXbgICXmEL8JzwcROsV1
uZTAJQi/p1AzlFe+mRfXyo196gf7VhWg5hU/BEmcFFO8Xw1rI3qEL21bUjRhoAFn
2NcqWDVWoglMidnUeG7BrcFW/2VpUCTCW19rnDHQSsdaLeBVxV4I9Ch5n8V6+kC9
hcf9p7D97Ykc4bQjnDJ9wsPWv/BxDAwQoflJGfKooYwwKezm9E5+5o1V2pOoLSrs
ocRi2mFduxr2hXCxcuVBn06m1n2UCbx0IttV8HeC9+DkyuY1ryQur5FnehRpIuLO
0BEfa4HTIGF2VR3VaLVNfeZYsD67Ps+jUT3eRk73856qpAUay8dWMKD8MkIdt+4H
ojEgLiDnzKE4NIrJlUlR6Uo1N9MvtOU2bV0GQnRvD21EpOq7u1Z3CRxRjTZdU07+
zcS/wqHIef7P/tPTBan6a39P3XSjEv0UlaycE/79KetA7dp9tK1hU4qMgk3pQDoF
a+smX0lkwVMCwMN2BfkXLn3vDiOHcTvktvbN/qd41WeqC11EnKm+TzMCN59ScELA
owQfHl+u4f6x6nH1c28/BhpaIwTw8EnJ3623yn+N36C1lS+1tCYXkV/T+QHNt/Lz
EzVaCF6F4SF2lzVsMGmk/YuzWIlcrQY+C/wKM7p4mPWD7T1rgpevramdDxybZLcp
2H4XTjpnOe/053oYJnvRxKXjWRnpH8Y5PK1EWNBlnnBHHRKaR/bj8sz7WDr3zJIq
1Zb19oHUSn9ClSXQyVt4RsT7sNJjKqRH48h+cv3qzxqAVDsupRcbm3wJ1/iSkZtn
UuLyGBxusMMpm+aWCm3PcWRypa2CcfDzoCnvMUuNmnaQBopb59HJlkP1qEK5HRO/
Taei2coo6HntbN2fxXM5AcW0gywr3GdzkxuqlHbiLE8ZlbFdoAbjFoWovgmCgbdA
YkY5L4ek+AtT8lBdDfCJLA8vsPgT1OX4M65IYvtWy8VHgKIhFS7p92fQOyX2sp3d
9UKVtVhIU1x7LMSrCxnpg7XnonhviTZcSQgY+3CIB3O+XP0hYDr9vU1h9wN53pOK
civWmBJVLiSh/Yune/2RxjjdPKtn6iQxPv+u9idwfcrsyU30KQgPKE5ODx8Iphxs
IEo6kEhhQR4HtIA8CnnWmCUR93IBuz8yVWo1Ix/+ZyPHiyTnhWUdGnAb+6PU1Ba4
Li1l8YGslNc3TqIE/qE7ta7oAIMxzbnxR5VKzSKFxF+8Ks/OJjKwb3SuvTbQd1EP
c/rG5QDcp1Id8SH2mZGPY1Z45lgLju7ku36QPnjCINugGiuDkwHRXtQJgjYksb3B
vf4wmp82tkf4zAJrI/NT24YAXTN1Far3chMPgNvSzg/NQ6g+plA0v8RKtUUaIpky
ESG8d9wj7bIbhSwvx6ZJb1UAg29Y7B9LfRZRhVQFnP0s8hs9jQQ79Vdv5VX46N3N
yHehN3gxe/I9SJSEFnru3R6pOxhZU0WDU4CuEzkgFfQukzxeuXfaeAwq71h9X2rW
1Slxypc+Ump/8HuYBm6Sp+CKNiRjTpd9sQIXtzP9dKXThShLv+hpz5E6qimOVbqB
AFwsdpQgwNGat/qFlr+q7HhS60nqK0JkzAyONqRvzuletL+oqwlVGmq7mjjqJzJy
DroYNbksuAUEyGUOu/6Gn0pO1S3IW4/6q+FT+t2TvilYO2KiiqlMWHk4DD5+D/BX
YNTzIitj6AUHb/Je7zZAMqeqUzNngCT7oGkezkPHs5P4a0TpuxL1aKrtdhVSDyyu
s/wDhmFfSa7SyM7ReOZyEc2R/znVvHKN9Eh6dXdr8NlkW5Ht4S0UtoReEIQu5Yvb
q3hN4BoRWX5pcruC+HimdJKZ1UX066fnqpuI4ZvMZELBC1wd+Ee0YxcDlU6VXaTd
MBe5OAzPf4dedRMjLq3jJNGu4GsiCPdxXojVdx9QLTZgWVd0Ad7ny5JHAv8zibxx
YWvfj5Ys6yZ/q5tpdjokGyOwERCmlkg0axFXdntmElsN4oNJf+WHYudusDkrQvhF
+/yOM8piPu/ICoayiLp6QjL9V1CwP75yFBdNVfeo72lek+3ob5lQMstOjjoI4k2m
f6/OOPOzKSieWkdomJlKP3SpXwY6SmbhMupwxKuoDZr26oe4f/B99LalaCNlUxJQ
Xir+S/jFOezX0G+zmvtgemk3EnNXasu8U0twgX68SLs4cDS3aSBIJY6uzuACNfru
RJlWruY3hb2MiNunyYx/enp5c0rxbaoxmDAq97FACX2pnDN/9EgRRkh9qgkfWYpk
bk1r81+52HAS73AigdyEZWEtkYG2ZEb8Gy6dALvTosR2yvT3GInDEKfLG1QB0s/m
0d39PneNzfXlgG+dAZdCNMrA7FXYJYjuEAowRb74HvEs/foL/0FdR6Jtpmg5ZXP0
4RgtI8Mk7IMJ0pySfJVPRiZD62MQlEwdmm2FnRxGOSnhWDqLrYj0jP5hMz6y2SVw
T3yT4wFJo2JJjoDM7DCJzvUEZGZdVzKtTi21yh9rYmAInTq66t5/xVmpf/WPsCI8
9Whr5Oc52JPIT0iqSrCzVmOC6q4Z5j9yTPY67mmlx2figrm/IgAsSRs3QS7PdqCs
hzxOp59BQObTTfUUvTTYZiGN5K4TTI5B9L/ZZuCf7xWR0S6x9cQg178pqxnyHndr
UKgPqxh9gBeSNa8fuRQ2TrjTM+0j4rh9zBj7KIiJ+MN8ElGXdS7vLY4uUi2riqoZ
bZ5MWeWwzKzqybJUEl0ws+oXnCVJIO4eUCvX4X2vugRYGB12h3lMrPI6wKZKr1rf
56jz1F5mc0O350QeWhWBUE3RtXIeGMTYpoE5SH1pez9TfIjl36tq+EgaNg4RbWbe
dKE7zgdmH99J94VoelKjVXbOz0Yy6aAzwSCnXDHCHqaOjXn0LC5umwVFtUynaiTX
VAWhUbHsmOQFW8+65BWQYpmqJ78DJDTgVa0oR4XdCpQYv2FJpJFPNOUxJpKrTlvy
8Uqwb1mAZAATxLHnNRgDerN65dF52OLx630dJAMnDbEhAERLHapEsFrlxU+Kcn/e
p0iucnJbGqE5L23gCPmWjK01xCrg8M4BYga9Nrinz598m+r/okCvF+p5l6YiwrqN
cvK/4B6GY/dhV2MQPqu9Qj7SR8Sv2rZx1cFCTxf+dXX2n1Inmk60zXsuyXP3N4Dm
yblanzIHs5Z5xOAEMBv/1xTp+6gGmxtHRcj21iFWZCycEhbn9waPQd+Beq7nPUVY
KI8hp1DpoLxlr6nN8d2GCGKchV7HgRSqEYllPGpVfHF4w0uRBJve200l6Ueh78L9
MwB8BxCaHlCjUKUvp1hATDzqNqAxgVP8qUeMCT3HzYJLPIR8QENYfac2lFMAWiN1
9mOdQlHNKQYw1jDVz1+RjP/xDRgRa0R+Qeg1szOT8GdebE/DQhSUYsxjtE2t2g1z
670vACtv6sGGZgOk5OwMjY4DeU8evv3d4XT5lQeYchYMCN96u/bpIXmW6eXE4De5
UOednq6y6ql6a3uHXIqqyVbNbQ4wUdQg6a3Bcp6G7EHH3oZes92Hfk3kLN/WuyPu
9rKtpbOP51WfkVakym/bD0rhzVzN+dP5YYUoeYa4BnOBkR0Qh+h9VXOuBs0JM6Dc
cT0OGQm/2a/mf5GCULCwVqHo42oojQ6GljtDxtQpNsz5sUE7Rstz0+dnixD0fvvk
zap020SazJrcCteWF79VTBJcr4UKqoOexF/ciskKJ4DIdBAhMgOLmzM1ZrDnwUb+
gOCPzS6xle/vvoTSGok21TAF6Ll55jhowuknHad4kgBGxRwDWCaRyDSm1/zzaMvv
yJBhjYAaB6ZSMDDcXj9Drv6+5p5S+kdiZ8MJAL4XHQCa4sqM0fhPT9QDRZEPJ75J
WkRwrxiV2KTIUOXJMj2IbcWutQFuKRt1YsrdTspKIZ5FSWMR0awZfaEy9pbPYY+G
KpyeeLke0HRDdr5nOHqzxJ3Cp/FxxL5sTde6neZ3O1iNAncwgt62LBc6GoJmDLgg
u1MDTsXvsi36LCBI6dSRnl+lizLX5VgeRSP/vX5Ps/a5kSOyHIfBAIbBcQmexmZx
eX5gYxFKfrrnxNKa87vBTfZN1Erz5ExSJQ+v5ajUpT4rWd/3ZRpQla6RM6T+VRoU
yUQLiABcfoyFXoI7r4wlLQ6vKZzWTqpujejod9MYcQtpgIPv+7+F3OCo8ZkfR6Gy
KSTy7GjH1SKZ7S14pR6pOfQVFYYVhuV0BvWoa3E5U8nVIwLMsPsb7po5hYIcqGQc
gtqEXa+e/2dS7q2wa41TyTxNSvnrU9KPxFoFyltbZmwMJo7WuYYjWv16oXHEUh+A
46GoX4bxVbsA8XYbTp8XU5sA/XvrEPbBp0AIZbsy0lUdGItDpPJglTatr2uEfB0L
oTdXRYGeAY1ey1wOC9YsBJpKSrsuQYOsaXPARbei9jQyb3AxKKy7lTOrPiowEV1G
qgjaGw+4PSKb3uq07hcfAmcf5gEYn2eu8cXG3KlBzLn0c4aDVk7YwNOEPD+2RBjM
iWJzuuxL/a4ZtNqiZpe+A0ob8sQ7UwRAsXHS5lsfRw1z4hrSQdC/SW2f2bukFRVY
60FycA1ZWFzuW3XB78jsLK0z0YyMcUBsiytQTmNlX9YRPgIMIm2vhOhTiqwgasBi
QDXmsSlixoOvG6EYRyV8brSlxTWUxWbMs9Bo+sSe+hFBKZh+Im9kBN7Qo3uK5zxH
M+i02HbSjmfn6thHDzMVrTAFJHjuyVfSudX1Ut91J+NJr3a/zCu5LiPN3mIHDduK
kthxx7GroUshDYXEU+fDKLAFXGq3ua6Zjtt6O+L+mxSzRF+fU2dxpSm5ho7TdzNp
574jWWUDS/rrTrJ7vAxvaIsaYuKCtXeW+fRk0OuyQc3zt6WxwNFt0tJJQrtw5kEv
uDWNsmwV2UznFyRogwJXRWOFUpM4XkPfWtM4/c+wlLKVEf+UjPcZwTOWOrHJRTVg
ALS0HAYV7X9Lt/TihT5vB7K4SfIX/SIPbF0BGUMIS8cxxEOJUmGRAYW2Qg058ehL
NPvmyz8P4UjXK+VvNsLluGQtGN9d1C0QklveJi2W5D3AgoyFLe8ydiR2eCVAljQU
MKC5v8yaSis1cVtWMvQpI8ownZHzeaESm98QZji5wiX1UMAbh2g1n2w2etDVaBQg
rm7Hl0S69XBqW8J4DiE8PuFNCIxOCoOE2NeMWTvCYFsSn9nKBSEaW8BV4WoAUC7C
Sr9DdDMj0gK0XM8X25iDIO+V7TQlVy03lrFQqPLlqazMqkWpTZIygdIPtMsjp2D3
dKVeies8urzLAbR7a/ia/7K1U0XM5mxQnixb3f6VQhWcCwd2zpdzasHhHl9IAgGF
RVrO67dguPEIRVbbHaaUTDXs68qbYnGKS1Eh3MqdZeuIU6GHekI9M+9DCeSzstno
q9vlS9XrIEW1KVNfIweAZA9dFrdGNu1u2DALMtFW6PrqlRlFQ9pC/O++4nAkbkXh
yztNTx4qQ2DieV5iFHnN0aib5dWFKBnQwdCzCZ/pIGV97DG4OQynao+vhQGJPBIW
L+6y5RuPzyudcj9GTtCewmZwlj/T/xI7hw/Bd/mlw0NMEumRh9PmT5kmX15pCzer
mXqXK5cDQwj2PVUGa6plfHgagSybinqSC2Eq1TAhDPn8jE06p/J1sdygnlHAC+1B
8yWAa0/EnKZ6LrZjxsnZH5zN1hVal+DoDy+MPXAuHb1n1+OY02A9cuyc0EbY0cbr
Dj9wDZwjww0xu7zGVb6UWw4bdN6BUi5p7Ndspso8i9FH2uzg4QIVGdslioKKl0cB
E2f9obo7ucMU1UiqostoHCeu12N3jsV7cIspolmGVzW2hQVin2WGdv/yuIw0qoJ2
QDqHqAM2RYNdGcPfbEvxrB5UzeIcbZ+u/dJ/UKE9S+qefm+graF5nxOM1XDDrn6S
PkafKq5t9ruxYxhq/qA/lKTS2nrHZuM6sW0Cs7BMpUcaUJ6H0tn3gtZ1BVFOiYxU
w6Ja03sfzEanD6cp+vtj8naCGWgxARU3t075NiNYr7Zo6OoFn0G9TACfiO97s1Km
IxbJBIUHF5J0Be+/e81GdCNNh+TKOw7wjXA8QSiTnU53cZDr2afFk0s/BvA4RAKe
c0/WA1wjs1u/TzhF0gFxM69oc+YP01RansAPlylzeGVqxQDZSx54G90kH2mxX5FX
/51V2pMYRf8TFeUaMWSpK+tZaQ4gHh381Zqs1cSqhIEDuvlrKaJ6ozY3tyEj0Pfw
svo+DkXGThoQqZ7L5S4zPjEGAfjIcP5PpL0qdy1IDw/id1EtLBk9j3ByC/ushQ2Z
Po5q5AZknNq9mNL6DMMX45ejPQ1QJGcbYzqRH3IKc/ZEUX5mnxh5RP1UAQtofFBn
6VBC6JJm45XFkhpGxwfwamOXnOGjv25avDNLJ6gCgwdetvcpvDLdAaZ3BsZ3Fw3N
x+uMraeW+jfa1WeiAEPf8oq0dh17LL0F7tPw7Y11uqiNtVvkEL7fJjDc+7DTRMw1
lROV4jgcOo91oOIb47EF+o55rdApNhoH2LDrQ4+DxnPe4KBhJlpdInsYTKAgjeBo
lNxkb/GgB2Gq8LBj13zQTfQrRLsHdIF5MVmhe9M8esXeMdOCITjhYyprBhK/hDIW
w9MhjEdo6+hDtkbWNcZvM6pIg8Jug5FL70fIyBHkpYWvD9snWEpLwOysD4iScEt3
4P0TRIGeiYpRWSz4zfWfMUXhIQe3awh4IVTdZ6F7GJIRjvGk/7RqCnokRY+50LqJ
v+icT+MkzBQbKPoC98Q3QqtPXUldueoIvS+NbX2RhJJxgR6DiOxNMGyrM7EOp5/Z
8xQtg3fh3fudRF5GpanW6gNoLgFhaOoB8okSEYvZd5ulxiX8sUrnVlc9WsASby1i
quUL/syagkZnX/sAiOmqRQ6cVTbN4l1drUi6s2QcNY4MTkxi0Wx2x4GElvOyt5eM
1jnTDyhssTNDGPD1oYHSwQ4jpcYaaIOzsuHemVHALaoHlhGXRQG3pZBGboBMUSjA
/5irBUNlSvtMG4MAFYCCfATlDmbhSmyIP5v/Qx1xx/V2nw5U+2e+We2xZSt4fGit
epyolqiYG++/rsGvoCn0LTZ+5Kw2REdZGKrGjZ33monlsm6tMP/Y3fuX4vJ0V48i
ww53U0Ib4jW96WAX+O14kSyf0NL/ZZ25X4QwwclQsCcNadQC/GNXrCqtEJg7Wcoo
2RxC0p/RvV+D/RNCO2v6vzGn8oxixBs+FxP8LYmMV4z+j7Rq4lv13bB9eGzMT0S2
um+UB6HdyMLPYdo/qtL7EzGdDCZCc5c5riuNaRoYP9fKEGqOqKLaVPBYEZ1kN8Uq
0fv4WvVqAAS5mJmVijrYjIWS5PzT+VX/ARWy+pPbCVxfubKpc1PLJGWPaQv+jvIj
InlMSe+3ViucwyN8QZzUgOBGlYBZKx5jmVerLQnzhDBDsRRGh2osL3YahrJ3YsRB
eqDfaUH4tXogSgW/v7sbe16VfQpt0KzGEfpBnv9wC5FHOKbBu7hEoNbI8bA++oAZ
XCwXEI2ljxEBAyra7pjU8fqQQOD+ALZYJqWAxknuEZrX3yvWp2s0WKYft3xjWoDm
Ahh2Q18N2YLzsSQzuoYNbbFLllHUMWuToNG2LsVBhcYfJX8s1Ksjo/HmtHcMiCz0
gNZxHq/UIsL/mTATZdYCLcmjcX8jMb87+jY61B8DJaCLk3nq8KbJPaJraQyhtsvZ
yfROraJudtDDzKCYml+r2vFoenFGaCLC0xcDChWm0+wrMfq8XdR46WxhC5jOxsGC
IMAbSxcb8Llmg9BWKAP0aZUjHHNPLIP6uKr3b+xbAZ9wagp40+FaY8uBD6cfXRC6
VQdgqYXRRwKHYjCLYVqO2gnM9wrRVFeKdADchSkdo0Tm/NsfAKtCNoWm76i4lT5t
2sOxAletWpvxJ0gHvFaUGf2WGjK4p/nz8gKU/jhr2OWzl+sqRYTkBSMxz59DywAy
BXiQ7/rDGaBGQHDNsvTQ7UKlRlWTM2OHC1TrptS4/609/Se/RzGikJSMSkaaElzI
dRtRUsGYHbiaBP1cCC8AY/SikAWLtgn/DwVpIvjUIrSL4pCN8QP5eXxhIfVb1NQe
XAhr9+kSFuvW72Z1sZqN7YUYOoG5/ebVKnGoPwygzzR9PmpKYh6aABaEC+EAN5vo
pMMUy3y9JIiV1edrojDsT8ubrBY7xgVNVTdQDdxQeS+hkjBYjh69ONL5NFFFh4n6
HMEHU/jEHwn7H5GoxsrhwHrli/5rYU3UziLo/YuZv8FJbsjnuItlLTVNK0/T8l41
kHnCKHXQMG+cagyMFGVnCml0elYiyP1UgKvzgFAl24gt+QH1PAHXDWpgZeWQ9/xQ
jgxjONZl11SjsmsIfnOi0D83KVFsWcCxFMhCSR/ksCxOGuZZOPgHPHaQe5Ls6Uro
tBadDwsgTD+sJbGFeiJVViOPM4V4txtD938qimXIa6lmLYZL43COnHn0QReW96tL
fJHUiI8tkgUMI1aqzmAk/kL6Ydbi5A+LxBxUl3+TZ7aJ5zaKr0CMPGFdbcoGTJkm
Ne+LqdQyO9HMngwJqH0OsqdWhi1vJ8hJdKI2nQ0Cq8t4TozonZ71/feyW114rzys
K4cIR7OmSmsfqxT6JYA9yO2v0FB5iluzdnpgSkWECtBo4vIA4AGo5SfT26UGoCA0
bz5+KWwAIq5fp348ZxSWVkvOoHaToS7XNJw/ijNVSsPnmUmCDDfSpoMMZv860GBQ
Z43GEB+dydlfUAhP/ZYx0acZcut9S/jITXS2xy6Klr4Wh2r6UoT1EhA7KyorIt6H
QPoPpYXvtkoP+5U/l4p19zgNa9Hz2RD1cvcxvMGPCqaW42v1bUVGX9aM2qrJO2ii
zWsbraJQWbb6l6QcqZt71Lf+BzQqaRhBgcMy0oALwhdot/zPt2My4Sw+zJNY4MF/
UjzB4kF28aoFo2DfeX8RNcvum3DS+rJNyVsR5SxxwTOmi87bqOXJp5vs0pcaLtHs
sPGGcFKG94v9GpSW8pHNd+yjiG4zr9YGv8tVnnC8R/9buQ/UySVgAzKoO3XIS7Vm
2zzH63s8iG6TOWP4T3M4Q3u/WShHjLeIWGA1uXCWkFX2tzCveD1c9uc6g61Ey8l/
zhoy/ktd+QeqtZtReM+ZI3r0S55SrW/ra90NicUdJXqAe9oJmbhqwBQapDfu9GeC
BaZbq/M5A8IzxJ9BpKDy0yiH+FEv2k6xVFVu5ywG8ZR2uIq2T7sds3ak+qeWysWb
QSq+LFLjBQvSakZl0Bt/si3KHjZxXj/c/KkMmTqQR1nxBrT28e7MdXla0CsegMyf
1MQ1uZqfZc3CA2R6ykTpiDJhr/+Rp5RccbLosn8Orb6HxB/knsXumXXHlKbEXR3k
iKYROSZ5mPWoOPN9qDLcFi73feYJhswT9tx9kdwewaMxp/NfrFmDjpt3WRVekCqo
gMrvJBhucZ/0+JBfvv2mtb7nXbZ/ReRbrrzoopMyomlKb4qEYkkQwtdXRHVXc21Q
QG+8E6rLrUNV6gKT1VPkAgjELVdoZgOgdPdbIUSZ4hImrZ8TPlsfBHPcwVX6NBWp
LwQ6e3IYiGfqDjfDNYRxhdL4o021dxWk+Yq/3LMjgL6z7PKPGQ+UImW7y9F6rBdb
dXrh1Agkir8XsJFXiPJGTFXb2VJ6Pc5dJclTAG9a6JuaZS+fSfMQ4UACVMa/VJi6
DjwG8hWiyRzIxtugrVjsxiWVdtxR7fmvXSYahPl6+Ktl2JwIGFcOPPxYRbwYB3bX
JSejY2iUEfAd4BHg2fj64IdI0zFyi7L2l3EwS6ge8tx8CnfHBZEISkQOPiownlTS
DntxTVKtsxj6p0mV2SdHJhTFfHSffoV5KCDg9ZxMLSqKSg06fY20eC85uaEY18oM
iNI1/45s4s2HtRQ0clCgniAi9ndpl4D7Q/TludMsGstjyuMa36e865XU9ss53jxg
B37DH3nB14er/5zzMjZsp+v/fR2HDk19MkM6f3+RNEYR0WIAhhsIkek4BVKpf+8t
AeHOGkSMBaDsWWNO+ssF8YfI1LfCCequ1VifaWp7gkJPTLUE/RPE/B0wgGFYjIjC
Y6rptTQFl04ozAZ0L/XaohP47bY3F6jGGaZpK2xS8y93sJMNqyX81r81E+cipuim
JrLzppwcNCag4q2L6QvNx5ZA+2aKcj68qw/LBKaefwtUQSiU0+14dOpnBFbw1FW2
7dnRdFjWuLzjaaObi4K5i1It/9Wuu78bQdfYnSBZLFBhRgDDYTmo9yQlKi3diJ+h
Qn/NJYhKnTQFX2JvIcmf6Ls1DjwnM9+zfKQ53dwV4SV4r4tZXf+d3T0DalkanMav
Rs2/q7HiytL3NiOrv/UXwtpOxznSsS8kJEoqEDEj1OtoBRdVUyW7UJXiQ7KO8WR0
wxGBvFyxecYOMXQjbpJJoe5LltfzhhRYybvELIOWzUb294eL/QFt6VA0VfkrcN4z
1uSCXZuetdOV0IPMg2apbGzGAtHzPW9LgpQrz5l8iqvI424a7wSPS1As/wdxc3mf
Y1NueTZXm9dKtcZzLznNxcxyvr6jqTHZW+yQi5cTDrC4SzuK33inrNWilioTHIX9
jXhq6HQJCEtIVe1qc5nY0kW1XPOmmqag0UGVnur1x4kSy/XkKiAeganAhQy8hy+D
3anFK5J0Ei9L2FDTy+HFwkJJ4KIFZ54PdgaeYk1XzEBTtZiwr9oszeTxOd5yti3l
t+SocCjjlxt3s2th7HO9aaDaexCgYkejgWD1KftxVJraciTitrZd5VhVpUz9wayn
nAMespyZ4GwuXrgIMpVKAhe+cjxm5UA67YXF/oVQwPjipO0swLrDMYvcVJjd3Kcm
M3vuXLAy6JFk5grCcfTV6YAJGNYDJyUSLu4WGk8RIt7oAAZDf9Ea3THjz8GAm6O7
46dB2byxv2QShLjs+Qyr3ohlsOeicQgQFe4/Z0w79o3j1g8LTBp5mLQED8IPm4U6
TAIWoE1lWN74Bx+eZi+88xqZVI2h3NaOMVGyGBr+tG3Ug7gbHz1Ml9xfm3Sp08a+
8oEEYn0RWs72/HcndN/uYRzFLv+hdbtXi3cfHXPwbUaG+WEcCBuOhR3JU/pBza5q
jq2Gn7hreTYDYxAPZdr1teUD00EiEcplEbgrxzuaOgkty/JoNVYY8t6fxm9FxuFZ
xwgpnKRR4av5/7Na4DaJiwxurrpj9DvR2BNigj8dkcQxWr2+sPRfgFwoluoEgd/z
k5mYaZyYsR1DdRSlcXvBe3j8zEA27VQpuzj19mEfNrqhD/q61OsSa4gsLt9689Qy
IgVNRtyP5boI0mz+vod4cPLcDibGS15A0tkSOxJ6dVS1ZTmNuiTS1OnZ0Qr/GxsW
1eRku1viR/VXt/CogMhOBn1qYUiNVyZccMtMHPmldUYestnGO27EcxlhP4z9pIn3
w7vKjgsNQknvusP2VeQbGHMjj5gZ/eAXb3XWpq638gsSs394R1sqOHIXpqshmih3
9MGJ6Hvin8pR7ZwVuQD3QIAXcHWpXQgyA+IjcSiWEmIECABA+Rd5ilrP6OwJ4PT8
Y5H2qAIXx7fuZzOpNSMgm7OI+HaLmQe9yxY9kbk6VfdAw02hRqT5nDYcBJ42eSoy
guUtPf4FoISl0VN/nMFbjkahQO5g9cMaR5sowhZOeqbM1TnZbDagDzkarsHR1qI8
M8Yrjhq+oV7o7rO6KHE8kXjksSTZw1GiXNuLOuh6v8v6pymU8XEm5aI1ifJQc9Cr
r2lDfw2w4w0+OIZFvq783ZCaonQ1NH+TCiyf4lzFc+oVaCT6kkF9muy84052zz5b
HHJoSI+/2+oe5k1YuAVOuPqUcaNp8JyGb/7msjnb0+JVYl2I29vROS10zRJINZoG
eyJ6g1V4eTPLP6Sd53Ve7ssnlJC/FI2SG+MEs3zB73kFEa7zAExNb/TqiX5VAJ3J
gfF64csGZy3fyRKqwk3dqUgr9iiLwzeG7vZga3gdNrrc7iMCcmZtUljlO94XMflk
U9os7W2DYWkwEu6dSnMbFcoJFvquMstRLwZaPTVYgAQcrKmUq0UsHt6ZrCg0FV/n
/0/7CPi4mTeLRTno8bueclG5hSflkeMVhw2JDJBBD8DFkKaKz8ZNx87+o7MWwmDd
lNI0VBDan5QRrO2wkueuscb0+EOn+J7/qSL1KV0LW2T/Nyz+OSm/tXSVMlN05DuQ
rdtvg1IHogx82Ceg9pVGegI8um6NgTpFA0DCxk6V6UsxYOxaHyFa5uH2vEFI3uX/
PjrTLzq68eOz1x2t7+mdqKAWTVco2puuhm9v1x8+n7Qe4eYxW4GCKXFytnSB2lGo
OSGvja+6wlNGcOsfy/QJauZSzzNYlmXvcn7jd6pWo89RjZ3z/TE8VylZxAqrQoLV
qQgyqdFY/VUQyKnZCucyqnY/swzKFl8ObFeYMmnMJ/ByOh6L9LHYU3odxeWS5Qub
+aVnved6uVfpV+WkoWHWgCU/k6YYOmY9Cv+QG93xQm8/bx1rZeEBU5/I8AkJ6bFl
ec5ozXN9Mi6p6+tvgQ7ASMgykaP6FCYzRhNAUdwF0QFr+WthMsithymIS+nanylC
iKngquPwRV5snsPCnBeS8RHs9rE/G8KEO4d5CrRF5UYnfOizIJW6CFbveLTWOsEs
keCpRzwqCDfSaAvq+b9TbEC75xOoVMcDi/opqGpmCdJNb4hwer6/yJbSOpIuyNep
dZVYGo69iFZsLbOvEgipGqEo9dzY6r9DZu5KcTzJFtHl6P/to2tpXVX9mRh46jy4
lXxeVya46Q7XozjzOMB0UGgPNkd3tLLzrOWLCRCdiiNDI/FkoiI5ve2PrLodHtzh
XfndN1CA3OSzgyYuUXrWsqws2QwPeL7V/NQuo3lTSosRMJgupz4Z/52QtVFr+OQT
7w+E15vXCvjJXyO9au/IGgFVvx/KOsW4ZQrYzLYApyV/x+qkd+zTicQwE7/dGT+j
cD9o7G2QnFu/aUcGWQRS5CpNE+NGyl4s6TgoHieUkKpVqm28v/ZY5zAIWmqcibOv
FqxN7ExeZJavWoz0wcDilYmLvBCL9c2aBVnTiWXFu6XGXIHMkax1akwVOEmCaFLP
KOJkq9uwhESy2+rNbHoNpL2shwg4fTZcPsctqzJ90wCi9aUCkG9yo111wApxeT8S
KvD7/UIUV4LzW488mQG99vcpd7OeYcCiKzqWJcBJKBoDik3LsLFl3lUym7HC0q61
sal7TIduGuCM+SdhEI7jx+A3W19fnwlRB9h8u0QgVQ8aBmLCuuMNZW2+FhAETmK3
rEmFA7mVyiSCaFNmuE2vIWys7+TaJVTxO+sYQw4fAzI0Vc8S5KGS/7kzVfnrtFjX
LD1WzxHh8bWe++3x5GAGwcd9OdiIVNJdrbyxUHXIHKaDUqqbj0ew9Nykpw0CBTIY
BPtUF3Vc4B71maY8uYsBu7QwTHMk1QAVSw6QtDPHAibUrbcw+7SitmVnNSNWnSDJ
sOHX8uIlvGARQbf0b9sA1bCLfGE3yUfnfnuBqq9J4c0j4LMQGC74aQ3ULfy0RzCL
qlCcYdWAx4TZk+IIch7BL1PJJb7+f1fJic42Js6P9IrQXbQoCymDBan0hG4cDEtL
MPEdBfujXlw/js2tFIm3s5anERTXWTNbrIZZ9Jmyjv5eoa+UNyPOhwPDxA37wPH7
QoHr4RO9Y1uXK2zeq7lIeF2WlJSyglkGtIQW4q9K9kV73Ze2ndcYf0DCmXtys+zO
5XOwq+fA+SozRJJrjhV5sRjeu9dcsHw9ckzJInyg+LNfx0Gx6Ex94w0cETvy8INa
iOypdkbxt0VvHcX69BlD++YqNslR+aOX9yyNablMk7CtfG50PQ0V4HHuQbH1yOwX
t4484HoDaOGcw4RvKnxT3Aoi08E6tXKNrJ5h5C0T8cOZ41KQJPAC6QRnxnc2ZKcO
H3wOMR+eGOtXeUY+6VQglKOijBdNhmIgIg2ouEQ8zFda5h1fSLU8a3/iLBKQRHCQ
eBbRj2JERBKF+JUN6hIVwCa4f8lgenQBf+k4EnTAB7JyvuiPfq2LouIUbJSKQbQr
6E61zAn41KLxfy/wn6UdWg7u8Qjx2z1sgXpEdx6dr6MeP+DS5cfxFUwMwMM2d/5L
+sfHfzCkx6jXGZQs//G7txW+gSAyqwGne87u8Hh5ozRz4sDCRVEb+qa6zgwMU97f
6aC9fcErJo5JVHN6LpzX8XjxtER/GiqTGc9XSfeGNA+7680BxxN6H8UesTinzaVw
Iruz7hNLzVoUpRtgtf9YCtAjXtNARb3Y2+R0WqF4Lhw6gjANNhNeJS6+V9Dx575J
e6C8SbkI2fbiDbBSudUPpfW8bopnxmIEUslVbwAGkuezirZXV7a7Gao6VcuDT1+p
+yg+PrAOKSmWdh7fj+STqH2zIEZagkcHVMzvnHLWl2zbYh2ENpow7QMMVrpUuvFZ
ZtpoeOa1Ac/wRB6YPXQKnui4X6CADxaB3sJMJ/J4vLRAcEzuHyulQ9g00gRzVTc1
QY1uXtSa66wfi5o4uhVtxJeWOO5ZaC5c0LpYcKROTQfCs+NIWk8JqMrjTInOmhGA
Q4SNCTZfA1wEOC7qpQIF5fgr8gId1D3WSRlQykhZKSAgRRLnFuqt0SU5YrnkyCY5
3spKx0DYiCxW4d78cvhF4aQD3duFcMpqTDqAbL1RaFWsR0jbOWyVEKPrasvVTLhO
rr3Ge0NsQqqzDwIEZVfGlNayEmyw2MbEVoeTq0oIT8xATKnmMQRCCHmmU2ZgX+ZO
eGl3mhvEbzAHxr7Piyuww52HWMcEjTCHEkjI4/Qhy2Ze6l9B/iVMFat6RLbPO/a/
Lg9jhDcAk8RriFRrc6Z8KodRnrZDI+qnOD/e1ZD4mPOCKrx+sDoX1FSz4ZCqti/c
wmFtVQs+Pp4EOQGyz4QKCkfTMOOXlF22GVKfEP5bbZtpEDX+A+0kSmWP+mBcUTf1
WMg2bXRuzBMo3ggRtsMsSp1FcZtnkELmb3Zz3LnUbPXpvyHO8WFlD+nFZ8YUUKk3
ltVEeiAD0aOZd/Yhhzh5NeZ8w/alXBVlz/+L4urZVzjxTE6fpvtCSbrVKk+tGUYJ
ccucxYqFX9a7wCZ+YuwLsXF3G4S5NVL4oaHWGD6CkcleoJsgGvQLlOLf5LCeFNsF
MC59gFhMu5isL7j7dQsfbxDXxjzuyJEu6qEKxYc5OyAniCWZoNY4lfirtnopv1b7
nIzPjclHwrm7FMflWnya2fIOzqlRm7MlszOpSS0Xea/nZYw7yDX3o6quxoRBaqFt
dzj7UpCAZwuXPkWacWJgC65fsG2ypD1x0GQgNmpmz6etLPwm7CHSD7adyKG36W2b
ysf8CYgyHc1zGCjnIc8HAjaOyu5onCDPOeS6wLIkL/KAc9wCmDl3UWNILcuTIs9A
a0nPgMJP7wQPh/SG8XktRXMaps9abAlX1b2apR54L+t6h8bPiiojMBMQ+7EEgmZP
+6MDm2njYjs+bKqdqiPsTpPATuWNGKnHhCHMhcH1qRsoyctSqpIBijI+WyuW7ptx
bN5ZsanZljfLcY2AdRVXoph/pncmADmK84MERO9BtKqrD+Jg11NU4xgDsZeZrMCF
pDfBmsJEXpquJ25RrXPCHkr30KA1DkcsvLoZ3wQXDUUIBqjZM90fkQVNUaIFmFsV
vzIriveOMwXp3sckYccMkYNlTO4Us7Lf5ShxJOAAPeP8zJdp35AZou/a42OlMml6
6hnzVCLeCcXHWPancJaHfBI8Jqnkf3KuXc5vAxb61s6UkGXUSFGr1c4/K+aleF3s
9mG0rUrSnyTEM5ULlPLG4HSwlSjsxzxSefy0dQLKRG0rE7rYLtpykDVaVlivClng
`protect END_PROTECTED
