`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZztjX7AwtJx2Q+/JL88cP0vCgy2rm/3/68NLK9u1cuXLgXpzh1Wc2PitkZrUREYi
wYdUS+uxohf4BkLyXwTdiepClvYfydEMCHNKyoY8Sz01jlu7cs0PCreXAJ3jXi8g
Z/59+4n92lPWXEYsvQM+MqMQBOOcJZGzHa56o39RBZYU265kuBfY1aOOo8fvisjI
lWUJrXX++q9yftQ7LEp1PAFpDh9YOAziX/BXG+9lrByDQd9FIu+SQ1z3XdOuh2x2
qOCvjXUo8RqOkabHa+HSlFKlxSOoLrAm9IF/M7fVUy0UTxS86ltwGSlEfqy6wkFq
LLXNrpxzVx1arrqgpYzhJ8mgqMAfrnY+gSFZIhEVNfuq7g7yj7vV54dHdPx5PgcM
RK0WzghBXun4c5R0690V2B1MqegwaqZgilfCDuTqGceII6/lI9t2i8D9qlWzD0oZ
`protect END_PROTECTED
