`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x901+BycriEkE7/t8QxCLB6TetMr6oAwFd5slK5EX0GqxgZUTmqDNbKwp+rfpC1R
XCRqKBL3qVt19sP89xdMWfMsCmuEeoBg4uwXOLjtaC/Paag8wQnc9UFceFeh4KeA
ihPEg4rgpxFS0BX03pYnSsumXqZoLi6dIhfwiXVkuk4ugYJfWXqbI76fpbz3L6fR
ZrQE+ELkynvhu9DO61ccnLIYbyPRI4N4JKUXQY/zUMs88roKZ1WJDrgIU41nBhpi
7tsVrsZX6voS6nNFX3nxqpJPkFro6Ktno3zXVeGNS6eiOh2YNQrIP1BjU6kOUIBq
rPCmmjITDrJnP2UEGjkhPVOmn96eKL0E3OrFl+V7c3DI2huUXz8nHeN909/tm+Mg
Q5vt7RK/Str9kxwEya1SIpNnimN7Zw2/EnQKbERiZhpEoJdS6u7jWM+IWj77qO4y
GUq/2nKh2qnv4zK31pUPT5aJeQ5dY+x7d/FelRX33nesVTrKbM4NHX3COWWBk/6G
tIZkXjiC3tFH3w9IevJuK2iBv1VVXz4OBeV86mjsUqkNiFa5cvfraEyWQgkbF/6q
xheQh60bXgIhPapOpAXErNQ60E++LINgxVV+MF+KtaRlH6fgRYkVssDwpr6Q7gQ9
36Es/bqnY8tyeyLHy5v4OpPcZSbQ2vLXMtZIJatDMOk=
`protect END_PROTECTED
