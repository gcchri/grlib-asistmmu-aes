`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ghjOe+sji8i+BMUOtQ7hgEq2WMmPQLQpP5UfEki/O9wlwAFaW2fOrYahgol4klr8
hbpgZVQbSb0kyLZ/CGbR9bVASwnzRou2jsVNMeqCEe8ZumqpLIpp4d29FbT/c8im
ZWOJTXISDHfW09ZmMgzkaAFFo3429LVRHTtNpZnUPtQ5dBkScnszdKpIqeivt1b3
x83802uecd5pDlZMQV5/3XAtddHpuhmUiSEGh1BkBw1w9zlEjV5ju2ZYcCWIw3A/
xnlvdYt9RlgyuBWqHOsfm+54PWY8bDkrmLIjgd50/2zm6qMar1CLjXDdMShNMMG+
yYJaaZS9NFiyv0tplc3SfE31liD3NEVnUh21991sB2F0eCzSxm1iQ/PYjhp0FdGm
fQFKDmMynm0maUYe2wLdJyBo0EGkwsvAXaRuSGd3QwTvhjwpLQVd2MtEuyRb1TQD
jYqx04Vo8fD2uZHN6gkd9Ri+hL+XmGJkiU4n2UJrfxP4tOXsEmelaJ7aMYHLeF/B
SjOXb/8u79tkV4jhjwSnaNHG9cBwJo2EWZnO9eFClNfTAsciK4M5trQ9gLcajk+H
iMHnNVI/6R4xlWx/Mj9uf1z5zh+gAFAhoV7+uW97Y96w217kwYdGY02bvhJbLvWk
ElkY5OdJdmTiEzhzojn4mOXlXfCwJwiPRgcz557fTdZ0EZAsc1O/kdOgzOoAjE61
W8zJ+Ms1GVKzlOjW3sMYP52KtlC6MU5bpnUls82rDI0IUdv0SSwZvzGZMpbZm7yw
ErPMRwUmXEWuDE5zkGg+46PEONlxlbP7pHersF+oZNQ6G3nZ30ReHan8F5ujrh8F
zGTdLcEGdx0jXJeboRsjddN1hEzEvqZ26IveHwbFCKfFfWUBwOtxSWpUeQt/RQ3K
57azSY6cuJsru5X+7XUt+UeFvPpHG550KBzf/x8cvz+2rGg1FOp3pjNaq9Ivn+S3
iV0XTtL8lm4rPuLQKSW2RlNR2/pUzn7ByTLs6m7rLGp/bykz6Syuk2rPI2wykJ/H
`protect END_PROTECTED
