`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
88gbg0AMmj2wFRAa1CEQQyWXb1cAthsJcYriWTIHd61ow7h88Z59GnU35EJYpp+i
v+Jg1CahDPAXmn0MmIlevX2o5DHj43TiVDVXNHQ0iTpZGhtxVVLV3Qz3m0qrkjkd
ce8ufRPdtYn1hMEXuJKHY8ErWC+SOPCQ9hhfRndgeW5lOSKWLkgwrpah1D5hl1Kg
Belj2hekvdipfjijZtLGAnzbL909/NJQHGg6TO28SWLuFYPn3IS1Xfc9/Dq1ROyj
ya47ECmY9o0d7jylb4RcX83hY08a/v7U6iYjrMB3dibiWRECHHx3Hom6pOBOzMD3
w2vkE/dgF1SCkvzIaBBSemNwJ2BRv4u0Zidt2z7KDgTujy1Lqmje3Z+E+zOqHKED
zQ8Sfrxz9zrtfqByUYbxgL9bgt+icxruXx9cjJ0HcbTPfkPqMll0OTL6TmawkBDj
G0M1RrI+6BEHo+D+gxHXVgc5Jq5rBp0UaIVb3eSWygU=
`protect END_PROTECTED
