`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/6rDAhX1cZUhJjzOuzsk/cN6LxGFUelW6yspsYcaVwhF2zXn9PfzFKpVvCBeJykp
Z8Hkm2rA/DIzu2quurFkYtRowSvpL4dGt5kev2AfDL23bt2TKJZ/VSRx7ybpqViZ
6Vb2720CAUycpki0+aoBCm9ZQ7Wm5qwNNPRBItVReloDlXs1ZcFU9v7NNYtFygOh
c2ibI+IUW/CEti8jpJUSW7j9huY8oF3ZfK3OPSwlLWXjdZCMlAWbXam8MKQ6HlrB
JvtSCqXl1jytSZFQ+r0/tw4H345ZMd+vhWplAQHMzY4rvUDoaXx86/C4fl1vDRuR
sflKrZaVvCNw+PzaqCIgBCvBORhZA7KvPNopby+B7kCq0XXwN6LmM21P15VWKii/
PyLFcdiBbK5taO+p06ZiTRqlY7gFjB3ef4Z7mQksAqwx+TFIoHZwy4LcCF8+Z2RA
fATqwG7TRXhUrwnDR/gNWQBQhshM46QFpbiwywfufhpZ3suHxEF6jmM5s+TYh1Zs
CdHDlp4eOQEbqxzr6q4q2Rs+onhdyegD18iCqxdQvf0Afic2TCHO58qazU5Zm4WV
0iWqzPIUSoQzXfso9dbZ9g==
`protect END_PROTECTED
