`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vc0Y3DrAes11JlJlSC+bQAyIF0FI0iQy4h5MgR3HFJrFqA4eRwgyr3KtMB0M9xIJ
RIceg05TE3ZP3O4RZ3eQTySo2RQB1RgQU8dWxv9/f1YFJcPNkp2j/Pnraled0wN9
oapwdT3mnZpsair9G5NhDGIf0VY7RBlSKmWDCo55MxtmlNJSRXxZjoy4ugV4tLOv
cOy69k102cPXBOuKTJrw6TP6J1tg8Ph8ODgDWjeqxaD4kGT01KhNiRe4h6OV+Ns1
4ZELCw0wHOa4SgCzu2n5CIIbGGPqzOOyUDn9/E5Hx7KfSYbpaQ17EKIMJ8TjXHhY
aXfTiHIytu/m9iARZZcLD8oy95lj3B/vEAVR8mP6xOFf8qEwWTRjdGkbKPme3WYv
Gfl9maq4I5dTzHD6hgRLURuszarzXa2aWqYoGk1WYnw=
`protect END_PROTECTED
