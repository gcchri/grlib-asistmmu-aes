`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qrpCv/kLFhA5wOJQ4cutGJHWK6YEhJZKA/+8dTXIeQXG27M/daB+LgIsUqSK72KD
GHFXSy0u1AHcbuO5EkAJOnxFQgmTryLGROR+u4pkgp/r7t7eL7DUMYLAYWQksOCh
u441HDA0e2EKKKlnMou2khuj64idAfcYndohv37yRxHtW9vx6sBM67DkdOAY7qQH
2KNQ4ZejjJJaHfF7as4YM0gMKv+qK4Byb11Va601FGCe3rIUBMOi6eAXd8Ar0qZs
aaA/yBqyjSo5SRH8TnBj0gxJSRIqbaDg7GereN63taZK8dXRK+JP8DZbkOrB0TNM
zd1wK2ypoQbK+5hIsl15aCbdOWeBLOD7M8r8l/wMhzMlz5WQvQD/IH4lczmGYmBJ
56xq1cmccwNiLMAQ2LXNuA==
`protect END_PROTECTED
