`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X9kSX2/BTg7U7fK9VUEaolXvtHAUqHKpFpvVh/AlNik5RDWHncGuX2C71QrIS5lJ
PDRwH50WHr2TOXd0w5xffLMJnCupI4Evv7gI4VFSHM1adHCUPaoZWe6ZwPAEdRVq
DXdRPlzlf9Ib/mmKYgzt1IOgVr0a/LPxB7+/zAkUJ1guq33AdWM8Um429aRnmpjr
3Be1HdFgsjE6w3yO4XnXJ+j0gYz0W6pamuTmwHGExwLtobKGdVzwSw9pc7AuClQM
DsTPYar9mJfpAHJWpgIEd6PuPmCGZLDMxYCjMOrnKOzBxhl5XVrE9sV4EvfHh/WO
Nm+VASsn20VuLC7K3YrB1jJgMoF1IYsWz2P/+kfLej3RKy4Vd3lc7RlVi1LpfL6l
XreDF8jYUHapUnePo+F1+hoZIGLftgtw9z2wUdMrNVDTgKBCQSyePsGd/8+EML9I
`protect END_PROTECTED
