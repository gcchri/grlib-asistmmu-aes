`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ElC1BrAfg/z4L6oMtfcjrcwCOtLdrfB2yxEMqCppyFrGfxGE/lFXEhvASK66sVmi
qpI/EvHri/up9N8PAbZLCKpmpV6VuCBoIz0+Cju7pcqwH05CiFOG1+a1WohYfxmk
0SFJMj+fni+hNHTv7Jp5wZd7cKOK8ai4MFBfR8F6vTPuqeYbeY6NH9jpOrajS7Ta
CTYKCmkbL8W8xcbMo3O+uWmCuw6noxkVfOefm8rus79fSh7ZUHo7Z0uHalKpnipZ
Uoh5hf+3yY2Vl1BnB17Bi9oyHT8a2B4kPt5of1yulu19yskU+rq3oBmVZt3KOxdV
zBsxZ0fZkDPfKg06UUTqxhw1qVmDw3CQEIO2F951NIS5FXmzzqY8/U13ookD5Ghl
BQ0JEsIHR6bx/ghRT9i8Q5GoNKDSri9fp4006a9RFoIGf9YGS+8LV+BBeh9fmYhc
d4LDvBSc9tGqs/cKz8EwOUy51L9S8O2mIzfF+ipWMvB5W4QNjUj6UjkE+H0WSQiz
fraPL2hGfgUBzou/o7bTysVmWKi4qyK7zS1HtaWFWg4=
`protect END_PROTECTED
