`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FkLNDKdMAMXAC3Y1n/TFaG4AfvFiaVBMZyftzVOQq3cAZxmPEpE1ffwZhBW/R3nD
0dlq03desFyBD/vZnVmXbsJWFPJjc8XXtM1v1YvY05fZ/sOUoTpD55o43R7Vi3kg
vhjT8DiN5POkFcQRAsdqxkXbcveaC7CYses4Tr9SOeJqvf3QXlwJ1k1q8BIekJNa
1k/cAM7lKxbHRxf7hZ3Qx9A2sBlx1L4il0VT3Qwv7zb0V/5Yzh+30onh4Xwnh6jY
v+AnTdOsfmL0Dam3DsDKfMUijVuFE1j0V9tQ2BDX0jLHNujAXi4CV251J9KlahNW
qYA+kmXtMeouOYhiliLB7S2TjviTcSEZEZKAgRgFiAd7agluOGa/utdY/XZF3DWW
O3q8KdnarYoG8mlfMtn4fP8dDbK34aRFnrP3FKNlj2LbSwNTL3cmurBKHZ0Auyw2
SRycShSVw8wrdZWV/wFdqCdmN1e4TzPi7L4Ypsrt4OfQACDq4DVmjJZwGZg/0m3E
XBA94qrFZAL3FWc3moXHQ0IxPgtoewNZmbSahMWY6B9fFIn3l/tUjF32DAjfoagG
6qz6bWyIWH1HbvPeBrum1BeebZ3kHwfuHXdGeoJ5qRhurfq6+5FMa3WX6x2xmFaR
cFYiPpMUWwpAA8njJG2+BvNht89PMeJdvn7rzDBqskOT4G+zG7JgARCWRivQfTmK
6MW/MpyCpZeViCFu5WdxR2F/7q8tuOUzs+4Ni/q/6kENUYFrz6pjWrH2fncdhc2b
uhvguti/e1u81TfyIBNT99s8kmZbPm01iyCdqyLQit3KcR3uT7QPhEelOd45Ybsa
E1kWMqYs1kWSIFA/R6GjA0VFGQm5s5J9M1fmRCj08ZzTIC1eeTtgyqhyuP9GnAt/
70VpDEit7o1DDdujtHh18EpHkbn6y92tgJdk+HxfV1PIxaLszta6zjLbHRw8bS6v
5hhK+gKaILCCwxnpys/Pwy0jT+1p/3YC9RdLfp/8vcaT0EfvUKkDRacqzJBtPWPQ
e/dFf02XDhGmFQ2r17g2M+2RNaDMIYrcnH+a9o/uOM9a8zTgzhK9VgnPbiGV6h8T
qcty68/y75leL2e7L6AdSIwt120nsLqwsLCTEfaWQ4rir7fACSv46HdlnPBtDjkq
95gV/EZzjPl28q9qwr8DZ/XM/VTXAT3RXg3CH9QbRVdZIARmGgv6uYl+e596+7PN
+rW15L0JPurphA+sa3RUH3Uhnz8bYjDiz4QiTbYNfJmNsCHpfqyjbIkC4xNkjm2/
lVEgwZprMxZE1ME1sz3vUJ1tFdfCGvn2zqpYD8DKa4OMI0cw+4XS75fuXDlx2BtC
syXTH/5FFNqWodusm9l8HsQFjm5ye66B9D7wC4zZBx0GL9y2IsYNuDuJt8LXH4qO
G7x8HZrAndPflr6cN0KWDLcwlSdLLDjYfnw/4mn5B4vnE6G0kZN/Abc0RfoTXBP/
/qqAyODhb+5ERdNEBbQ418XdzumTSitdLiPxMCBMxmEQ4vOW9JSr9RW1zxrtxJBd
KBIIxtuMuysoq00LxpJsUlj74magoxHGg47LklKGeumVtcm42xteIiUOl4Yh2Kq7
7ZriLlU+PTQN/kv6eGFxrxx7WTbHwoVS/jdOgHKpfL7yuhPfyPlINsgwvB+MZIe+
L9xO6P9DbDqIlF7LZTk7xLzJs/4BabdTS3XkKLF4BMiRrGz33NYaoGFrg6S1KbtM
lghnOwxaA7w8jE+5QyuueXoTpsfNjIj9cZfvdWVyfI2O9AOpZztHuf+Tc3PIQ6G1
98KQzc/ef//wYQjJJRRK5ic+go9HL70tXxEUV2zCYA9fWKSAsSn1KVYlHQPAptVv
icEBXypsq9pPllzacukvaI2JmtxfIZTlSYxuzAmvPxIpdJTnX9uk0XDoxPAZwFOb
nNgh2HQrhoyCgZ227spU8tWixwuwVzc/4G+d0FMkYgL2c1ukAC2m3qu1LtGI4q6s
1A1wPccwf1h6W5NkRFTtQzH0PhmcUQ8+htMoYKTJBRyq/wH2muprYiQxoJZ9gLpG
foi+pgoiU91xTSLftAEo7kND/BgIle01u7BOkfarZ+sPOJy137SBcJmv3Z8WifZu
zwTkaLQqTOrl5d9C04ZEl5peN3/jNIFiYLoUqeEoQ28p97DSGboTbyVggjQcwRW9
P8gP0w7PegAXy6Sz0UaI3SOAgahTesL6FHi+TB2E1moiL+iXAoY5iH301GmIy1n/
Wjd/kgMRUKXD9uM4jZM4L/cNjNlZ2ScCDuJa5PEA/iu0i2PoW1qV8BZa8RtaRs9U
xYo7wIIY07eMqjJQ8WcVwjXw8CVZIqlyJyuX6D9Tek0hstzaaosdxw8irwAtIQ9/
0L3CFSCwWjVoyogETgKQyDlRcXpPO5DzjLeXmWpS5pDLVOy1TezsmbKfSVPMJdbk
I8mr8BViR8ThiDZeSiBq72RoXm6/n1mpuiE+zZdArr88+EaR2Z/a5z7G8vRJDu3V
lFE70B4c+H6PGub3oO9WMKZyycB76z/ujfSy74zxzmS5D5hijaSjLTbMqQaSytOY
mxdrGRuJ5xkDs4PgBZ9DIXPUstyetSeS1VeikvLw0DIXhO4m+Mv4Y4tHX9tDsDeT
spZVhgawyTaZWf2vv607qOI30FcBUHuAUDu1iPeiHZCuEBrsq56k6oh4QN4ulWJn
jJZ/VfBPWUGRsJKXkV7/5bZ/x4xOCfFFt1u0xwmfjHu6Iszk9pE+88Dm/w835dS7
xd9/E/rI0qp+lfxQtLk06049TccUqvZvjL130c5lQqfbfHDOBPc9LLnhjgAsXaDw
Rtei18tNnaY+S5X9gaurRUV+cSqPuwDDfaroD/fG5wlSP9T1aS8+jc8VLYbwHiGh
MD9vrs2VMLfpj9zeQlrzNBYxTohU1pvHLmXfLZ6BBP9Tsda7IQr9I9WDRWNopa4t
VRCunEeCYGgCa/sHRTEW4gzqb80CCYSTrN5ETM7sBaxDA+rLNh4Hi3btO38dcOTs
GtDqbqsnesjDVIshQpT+SKrr7aWZQexzdrM0zzbtewjJ+86HumkJQL9d74YKbI9r
C1m7YDipkmkWomOsEE7aQv896d8KUkt0Brov5lNwPwzGq3KOIjWB7vkL7+iKouW0
Rv99SVZLGVgq6vcGw6WD6L8BnM8kBUV/rFaulc82pPeMZ0x+OaGxqjHtY05uwhGb
L1pA93hDqjuLX4SXzquSoDMCd/PvmXCHLWZ3XeO3qkRpyeaK8czzIfbIesHugTrr
h+BBFvy0oEVLxnAUzu7YArlQvSppHlfyu462yAcYuHHnzSnOS9GF45ART5cG8WWs
aqYrZCFzJrpgy1MrsXgcqybgCIm9dNqe7u+5jhk+JJS4/Y74df3sjNUG1ElzK/1W
QYKS6ioRe85H82roQy/4ptp5BzeQiDB7tzaTx982/tMPwPy8kLwyxI3lvowm03Wu
U22Q7wiKcDPBr5Td3FJ0TOR5+F0WEM+jklMrYOZUapGxM7FsRz5MKDv3GPMIWFPS
HLUY4NjHm9B4XPBExSh1jekrY1KKY/t+NUfqfv3stx9S4p4cp66pZ1U2OErrhaBz
vUCnBqEO0XaWsk+TUUXaGDM2bq6c1lJJv9XT7w97vmdQle/gkaHBbvg1P9BbaEY3
9DFKVeaEcptc7A0RooBMXV2PKWatS5prd4GRW8rXxDygeTkHgJ57YcpvZUIg1Ozp
S096HnwQJslxE9iEOhuNf1LyDr6++NEbXWs5eE4anlPBD7Yvq4seBgMzjFe4woeS
QB/L4KBTWYaucsb7oQkt+svvehS+fTzeIZqn+jcd8PIuZ+BPqjCcTumn/i8gGBJo
14Hw9YhHtK4lsCDSeT2cgDuieCqhVwfqn84Ev1hP6moGsQNNz6XaiY7Bn4IakAZe
VcdkVnASYBcBGdNfl6Hje2O6qjqiBct7lTHQCWMnZ4c1UPICTpXhDVVgjy5WAaWD
ILY41sQ6bPRqBSruV1AwfHT1vC4NyQxJM23kPpt9KEYHBYWQAc+EFgAjSoPRLTka
3Fndv+W3hLutlxSTq89UKU/3l4+lOQsd7lk7kyKfwZYePGw4CSfQpFtUnb9pjr80
FUVnlcXVSh67AzKBTppBBnAP2ygfl7DC+c5bjB1486o7HiyDyvUAnp6Rn2MSnVIx
ZQy7l047V71R4bEOfGSjpbJKeeZ66snRPNWaRnTz5DaPPhuG2nQvmj8cnADsQiH+
MU48gvt5BxgcyEch4G2FfQtMCLlWKYYX0Sf4tv9YMo2W3OIsCG/AIFWvG46u6qeo
kB1zwzEkPGygCaBrDr+y4tqiI+pJsrJwOfw9ly67IspY3qYS1fMC2puinVAwngLY
RFdqhbmxEi57LmPf3C9576BNxzcj+tQ1H/nSGeyzjhYUYJK5mMiAbzUCL3FdPFVi
Doqra1EcFES+z75wrNhHKxz45xStODCzZRIy+AC2X4heE2iMkxHp3VKVrk1DdtEi
AITbKyMXuPDL4S55ZHiL4A==
`protect END_PROTECTED
