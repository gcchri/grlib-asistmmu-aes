`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fVHUig5asqkF2WCJK0WcTB2NDG9cEQqRqLfXlxQAZ1B1/DEb35u/uw0JNOOpRcRH
zwMr/WZL6CQQgbeQh/KS4uI/ZeYIj2e3EU9nOhnOBeOA1r9sBOA0axN8dsPzMxNy
Sj1Gwt58+Kj77+GzKlv5Nzv5iQsPBVuueIcsUImdM3/rr/TJMXpTFqUpGIs/m2pT
VbE0xk1Wa7rdV3mteHkIywjm/y5LgcU2wifyh877Y6EUycNgff8/DA6dK3ebu5Pf
LcoiVTLEYairbhQI/d5xNhTR+VHv775UF9JzfGB8Inr9fDmJ5U1YAjHSoRt6bh8E
dSXIcZRWJbufjB3jzR774qkfsr6Y1O8K7n8dPRadE6vCCYoEQ3KaxxFlrt4YwNdv
MvXoFQbEC3FFcsXKfQq+yNIErkwPtnL22xiULxEtSkCkYJCtS8iB5TMlyEC9+p7C
8G0awuuNjj1cEDt4b8iqn4jzDVL/LXR068pUCrjc3EjRBhv2/U7q7ZGAqXzYBEOT
`protect END_PROTECTED
