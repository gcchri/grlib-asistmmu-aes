`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eg22NRATEv5dIg1lTyiEFTU28ZZi37JQhJMXfrSIhghQ4mUnRlgEUkJL23WAIMav
z/3Sbk6hIVpg9lUdvZMhCeypWum8CokoRszlFWarwduykSFPrzxpTFB03mQKhF8m
molGibA7cRYKZIBiwAcqg+5KPclc0Ni4kAXdm2x4V5WP4+0YmyBS9yWClUVNu5p1
7bkRqMinofQjN/bAuhcEsmm5/xnRbk37XlIhKTJ1eEDYsYimC14Hltfu6Fe/Ij53
nto/sYJyrQpzJeSMIoHTV//CGFT/Dm8pvLlye78WH5B+i2ZtlkghZ3A5QDcWtE3m
AVm13+7081Ela6UtJGfaNA==
`protect END_PROTECTED
