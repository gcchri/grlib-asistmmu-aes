`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zw3d8y0+ilDFqJ3SpGQvT6wVWcOgJamEE+NIJbEGOPfUGyW7KX1J0uy0ywYavCN3
xWP8AoX65Cql1bSSg5aHpk1axw4nLlMuDlVUGj75qWjr5CjMx523i438/CZ39rAO
zDrX4atXkIHIUFPqS39eVZZI2Bvn8Pwt6R/io/v8OCTLjMUFcS+UeawGH99WYoqo
+HNHwzX/8jahoXtBYjn2alt07f+g0RUdp9q1iXhUa463vm53zY3OdH/A1Tb4I3TC
hie8cvQrBxVT4DtcXoQQIi9NzvNrj84FjEOPZ8SDb8FUY3nIijYEjvgDDR506LJa
ax5+lNa8CFE2anb93sfCZV3s+IVjnH6VmurRhAI50hDaZu7tjBYMeVF67ZazVQOM
+CbuVSz3cnmTWvjib1iQpEjF9cucavJNLXVszaBRWgwY9tMfBW3hP2DYh36/iYTG
7rFY88kC9KFSDjP4b9IRfiiHR6S2UKf9F2r9o/TcMHOA8UhcpaWjebj2PJcKwESx
1sVSfWjSJLg0D04kqnXzbk/4cUhBtTGHdJN4JZHPDLJQ3Lgu0SG0T+WltyJCaFjb
Q/JnTU7L1NzrQTQ7bB4zYKCzCMP6iljYYq+TDPJE/PtPUAmTUnr/VSFagm76AFkH
h8jyjrghYB8wI0ECsI7dZMkY7IfzDCTRCRzPkRRz50J4RlJmLH1JA4fn7DKsQ+sl
BJQVU0tS8TDdiXEGb8hd5Lyph2s+fsNTz58iwiNhGQViMMZr/rP2Rw64zeIDFT9r
CeuRDglz99mxW1E40Jk54hgHWXw2bqTHamvwN2J1QubDKbFMcBm80cyf/7Zy5utw
AkOVhC3IfDy2+/p1/rNUkD/hZ0U8DXD2OmKvofJfOjgGIjJqvQDBRtVsvWDTnlHb
qZ//rPa6K5afbEjx8FHS1SQnJuaQkkdrTOE2a2XwFhqyaKG8GtLC5ppxVBhxneQU
MjAavmm5cBfopWtOPlGTC8ba9N59dy7LngESNAY65hypwA9eMmZih0OwKuKuTkHk
T6S5pJXEMPcuAUvwOUhis7EkF+KPIpyHRt+XW0ncpNSvdecwY0x/734O0E6PAfio
RMbnkqD7UbvRkGXqEW5g8jXAKZtQm+RKV0JGFsm1lahhOldcoMacd7ZSAXa86PKQ
GI7O4jbz4fESjiOEkcv04nUnxMOPVkP3aOFhDMmWP19M8axw293GSG3bikhyn0g6
0Hwg96HWjKYYL0LBxIHIkfITLU6+c22FOEUVAaGKx8J+qcbf74OgSaiJNZqvdNs8
Zu3j08mcK/9Et32VoZ23tqY9tKJyNioYttosJfd0M/g2hqU6vWV8vdkI6C2ZrUfe
/J8Jsr32yQpNGczUJqr7tRIg6TB2kHr3PNuUEWmUxMHrWE8FM5rVEMzl1IhcXOMW
0ru+uwGE+qES7eBXkdLqERBxkTXktZ1K0xdU1sPX9nezBGOz7aVVs1kPL372K58z
zgY6gv+734OzpJtx5Xj0Wb14wVCTrMyZfYEadMwFsFIl8EOPqripPUZD7q1eOFl2
c4zK6i0ta/qejFRDSqlf/T2SAq27u+TNSc+pOt3jiiZCCVVnl7edBMte0c/xkYjs
s904E7hwzcfhU2FiotZHpX6bIQLSV2AhYCWwaFYIQE26MUzhz6kOQaNATcwYrW5H
pDL2kde+Ul6wM2UF9fmDR/cUvdPG5UwS1a0ZCMf2KP2XEyVzC3EAqhqSy9Qk85MA
DVP2QUxYG+bABv9X9Jd5aXfeRR7pdAh8XLBn/aAsmb5/SRVeBHxBmxOxZr/hqY3n
l4SC2fbmRrsJ+YueII9nDqLsnvnuXvMLecjJAv7dMedpxEKbmUSH2VbKt24rD7Uz
W+aMLlXO/97byT2r/H780s0zxeowXK+QqnbOi32pQcRcIMC7u/6Jw9NccRVuCWsv
SOnBAplUii7HUluP3VF0FxXLDqm3BWFAwlcCUanAc3Lf+RAyGwRYibzPwFDSOtLR
T7ky9eGxhJtn+TqlybmldTSjS+mrRVEH6hlkF0tRGtg6w7boEeAvMb2a7IDR6tc4
MteE6ugsT2omxWy9A/uDME55qj18yRZN7wNG+DQ6n05ebjkrdn8KATafRiF0IaDJ
f7vm5iuSE/crSr5HwAYLu1MaJ1EcD6ZfsdJ06S3DsrOlwijXvJHz/SrDL3ezm7wY
QmjC85FPh2t86svBsmOYuA0WQtm1wjuyajt7ywQDKynnJWo7DQDDqGxhcjC/UcXw
K1mqcKUU0Sk7xOt6SZSJiw==
`protect END_PROTECTED
