`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qHrCdxsWlgmWJLYFzrxHk/+GNsHfd1B5dsedMKaoJrrGiKtAB86eEc2pnvaaZS2z
JGf+zV61KOOl/WuuW3ElGBQy3VvKEVzVzZFi+kzsrrTqVc7WvhTpuEJE7fyvf4ab
EqVC6uBNCw525znT77E/UHSVpEtytKsW96cQMLbfwaiFH3mYlKxxyKCigZmDid+o
Dq/bVKi/XCJBRlPS82BQu685R23apkxvPCCwLsjie7oU7KZLgiuK25/N77USUdmQ
5jW0Y5rfdWaLmSu1ulR0seIyEFb+yLjldNENEnRSB6MD/Qsy9n4BjZDO+tCn7ntQ
Xu2YIzfxDLAkOYo6oW3ve7EKnxewGfQQHHgDmLH7jzn2OAcAq0HILCm+Y+smxCVV
/oOEoKhHOl3UBb1J2djpEvuEoWcYJ0C2m5v80wZyqQk=
`protect END_PROTECTED
