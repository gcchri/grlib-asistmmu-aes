`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tBEGBA5o9wBhjXQAbnLjysOcQAaDxthTE1xR4qp0GBOxsJ1vs/nVXGZ8rsHUxZOZ
jEgjxFnsEI5ykNmzQhLfdDs0lWLiX0YhoRzzTP2e+xWQkSFNLTS40BEgYjgplnb7
cSxy61mv4QUTX9O/Kqk9em132R0eLI2qzjTQNsxHWOidjgzZbQtkz+QfV+Kqq8gn
nxn+N4tr6VCkABY35fqXxk/4prRTdIm1Q1kU3N05lc+tjKA1gg18zUcSBpx+4Dck
UMMH0tGwoRsc8ij2jxcLVHPx/UvsnE/MBgDman+/4HvycybSxLLZKh3oEslNNC+G
ef1D427xF0fwAvK1GoHON8qmG6TX+aCIQoI2b7aBYEQHZsYOEMGHtZRxP3cOVDdt
MxjeADELpTG4Cq1iNXsFm2tXKKTS+s+IlBRTcctQrzhnAB2RINCJx7VZawqshD0E
ooGjvz6Ufo1NofFYf2O1NeLZyfNLvHwyVa0ULSOfJmRUuLnJzIqfiv60JlR6kdo2
79i1e5N8ajXuhxcDTpy19fIe/r3ho41JR55cC9JCCyNwKGWwG/F1qTe62rwf26J+
PSdgiVwZTYBJ6dWDCNeUv6WQpiepc3NM+cBN9RGvb+ZB8kAlXyMT4In2L+apeJ/s
1K28OKV/AHLCZn0ioJdGfT6u6oB7EQLbjSLVTz8fJKzx0I8/pHYhUwZ7CfXw52g1
mjhCKdiNXCllp9tAnwIHfD5jCukqWLyot4Wv6m9LmExTM5zeWLhwDqL98xEuXvZ+
1dHHpzWECYQTkefth8r3ybhFoTKvykV9rNpujMraKfosPXEy2UM81G+gaQYnnpK2
Eedo0s7yAH8sXrUrpm6mf0qN0qmlDH9KM32++9wsoZTnZVWYryS9CDshTHwqXgoO
+GLQfdSeZHHlU87vwt5Oq3sjOdOi1CynpVMkT15/lN+uuDivFDLe69UR+lnX9/Yj
`protect END_PROTECTED
