`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CcTseKb50MQVDuzXu9ZqOAnUCcB2VNmHEoxRbG1IyZp9VCLu12Ype0j/9E0Pbdt+
/DT/8CDuEzs4sH4i+jIRgFrBpVAi8xGMmdJDJV4Vks7eT6xz+yX+DcaOqXULyQEr
W2EO8rh4MBqZY16xNsl45GFSRPMRLgvrldBiPqGtKc+Zbu56SlOYxoDZOA/WheaP
4vIbI7tAZzbYU5O0LoNmd+WXGNTjbzOWuuRqbSjM6RAdRSk9E0EiAcbVHnYp4+gM
d79tpORjG3Mb8Jascw4sVUW/zvBrVL6GFLJYg0rWFJbzRtihz6VQYh+LMH7gQM1U
ugt41yYIxD4mX9LGJt7aZND8tPWZ1ZTrsrDtsEZBzZKCqZ+5rOzWUTFccNjqS3Uf
sRMu2sPUjmL0P8N8vHzRpdF0Iyzg0U+o96LK3BPIJHQpKpI64DU7YaZXN2s+ei91
RvdwoMp5WhGCtXtTIgAjsrboFerTCdJFyVJjiAGEwG+bQMa7LWows5avFwOwVP48
`protect END_PROTECTED
