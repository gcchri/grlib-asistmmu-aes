`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sxjjdBffIPkso6nWkZ0n8WUUg0irDEYKO4YN1T8RmlWbwchn2p65i/TAA/ypJ7xt
BixYRKWooIK0ckOqwc/TRi9AMHAvIuWFa/R7z7I3De865ym+qqioNYwP7kWGlG9g
w9oOs9svEjMjiURYQJbzDYa6O1/DeA5ZsvAR9xfMSywG+RXpz5Aww67/vIcssyhW
M5CWuE0seC951R+qcOy8tDvZKyrU93XucDjW7muq8cSIcf/PDIkOqdXdFJclPgjr
7T4q0OI+SSZPzBHScUExbd2xx8S6auA4ZTH9ZNLeml6MGmum9dxFv617C/XCfejH
Z5gtzhYz8u/Z1zCEQ/VRMuYi7zz6QC6kIsxn7myQ1NzC1zO3ANlW1pz8K9EyVIg4
bM5VeaVsHfWpRQek7h4zoVpkTSo+Rhd1L7h66ZCOwlk3SPmEafGk3tfF0EUecDqx
Ef1+Kw8wKu1pr6y1Qf/aORVtr5OCvB1qxwjkgEzGhqpvBy22khJIZfseBB+7vOCx
d+MShycEP4VwfBo5AT0Y9tKYD937uPRHfCCgt335b9Pimg05N0e81cq76Ad1lwVU
azu/VFk4bNXfbANLglrCtg==
`protect END_PROTECTED
