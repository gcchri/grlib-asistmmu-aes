`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lclf60vPmxqX+vgh9TVsn3P+3m+CWycwQ24YCWtVLRgiNhPyPpzSJQWwPf3tru7Y
q5EFwB1oKbaJ2IGqeuX34tE74kKgK6iq4nxt1rjHfuQCpCh4unwuo149/ykocJf/
KIj2FZIYA1bsVFUt6+zMzNHYRu9rSLXIlaYRsmHemEhBrRLv53GXNPAThQX6DvJh
Ez0KJ7R0ALMsBxPCf4fwz8WHtdWQYj/dOVTAoCkgvXhqkE5NXxXJLa+ShUgmiAp2
smWOdiuXn2yYerQDW0YmpW5N2c6u9XBsvylE+tpy0ZQcBpx22VHSoW/W3bJoW58f
fZy1CTGYRyhOZ2txPA1jajA9+pMfndzlDALUTan7fKHLoVLzOdjaCRrQ4xvQswNa
s1PuLC1lYWs1dkKmxfTx/nhycSBJ3h6PgFuWHjXo7SiIrxO/mvORXdkVb6J3mEEh
3Mt/s3879bE45DhyN3ASBl9TYzN+Pxc275QASDKvyiv4aQQKXYxXb3om1QUajBkG
GxBHJDU9VMR9IatkZaEjZbyC13cTgmsomseE5Is4UWbN8wcQtwCADz50P6OWMU+4
kSSeYPZfElcTLDPfO1htxzAYgtLUpDJdlCte8GuylagTSBW/f8FCffCnPC/2uNj1
NtgZSNup6OUhlksxE34gUXaKrTPAF2GZ20MgGG2POdQGQBZ0ukDO6byNrU3VEX2+
pj76Ul6a+B7O66az4aL5LmkRuzielAEwL/pz17zRsLF9ImqjZ2gXoPtkp+qRxtOu
Nvw2Nss/hh0/Ve4PS5OirEWZXoQNzQ1mDW4MqhoV8oDmKonsqy7Hw8zxyoT1CE2a
v1q9UGIBAVFzW3PyyV3OpDQJJk7PS4umX2CYjNMD8euo1lRyDJxpCGRoDkTPbZ6S
6BMqQqbAWhAQCpacRzFGEQ==
`protect END_PROTECTED
