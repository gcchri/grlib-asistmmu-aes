`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ap1FN1r/L1pH29KUTW0AkKmrbBEWcGFmF/U2lSHpyPHL3SaWVDtWAZvygoMpII6H
uqBktFFJs02jQ3d5+mDjgWELJqWrncg2sOrJD5T5Kl1C83fRK40MsGDT75PRd7MH
RsVyCm9DgpQ3xJqvDtMsjd2PYlkNlQt4yCRLex3fQ2vDx+pi0JYkuMRZNwbGmY/2
5hEi4ziC1+0V/s8Ls2MgBDtC7Ad2IKFYO/GQGyZhEBXpLuNeBTLjgx+14hQquk3e
LfYdIK7W7/i677+dQdwaM814Hzyg+D8MvL0w+9LUEJRH/aj+YUuberoa3MlbBgI1
2xNWfdsTxbm8nd9eubCJzZv8u5yYs9GG2pF1XvaPmllj6srwOLEqaGvn5Sp+pD6O
Z6eimR6/hoqAeaUQq/HyenP2R/1Z09dm15GyRtOqPuyEHRYQY0rizfsNOjpJsOcv
`protect END_PROTECTED
