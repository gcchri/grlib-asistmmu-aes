`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SlDQaox3IzCBFAiJ9rah0emNXRkjbSCrbrZ2YQb3J2kNMHIV7MOGt2Q1/lkX9F1g
sh25DoNXEDyD5GAXkZyAIB1Fmd8oQV6NRcmDXIS8gSdn+LzQAS9PLwNjHvdBxAl8
GTX3RO+9HP0PuSEM3fgYs8+VDCPPxr1I36mNox1jlA1PM2W8HPDyy/3zN/8ZMQbl
MPHVTOLDE5lLWG3XPK6m+71ESL+aMRrCUumsQDpv2F7n2xYsgzekOyZEe15ikKg/
JQURBlOLIuQEO1+BceWmT+RwENWdSEEZLZr0mgiJiUU2q8HghjpPLBjpz7wdf7jL
2KPpMMa5IkpMbOovHvdfDyvatwRjFaiCEwEEv6ary2vQP2mhaL8+h8oks2apUHEu
0TmgVeoC56LnwBP1ajmDpGIQJHCYNPGUrACeSH6K+KqRNErXJzAUoosVX4G6ADlp
YznR+GpnZrqjiUtrtCT016foJHrv8ot88q64b+Q5tMFsEgjzneu9CFSUl8m4Nn+V
`protect END_PROTECTED
