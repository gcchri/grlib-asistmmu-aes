`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/7YrSQbu6jpjHJk6B+T2UfZmEv6JFIWzfQ6QWaBAYmCzxHJhD+TF3m3qwCD3XBLw
uEDVngy1tCuPrvx8Nt4HamRO/gZN7mBiwsMlLPLC+Kgz/p7X7f20DaVE93EMK7+G
F2Jjf4I+S3X7iIVpEWLJd4xS6bAaj0Iz8D4ejB1lu4cCBXdc+p/9K9+EKF+LLgo5
kG4iS4cnimgmPY1q1R9618dqYqhnOWJyxxbeByfVsxEjiPL2ZlSQvmKuvXyKHjj4
b9Afk2zpqvjPCiVmQOadxxotkJl5SZ2mEGl6Qf6dLiBwnqeUOlwDzrghKp7JuTts
bfck6yhKzsPdQWW2SJeb8q23a/eG/qrvWmdxlMoahy7JUhFATwO0C0ZWgdjBIgTX
+5FuRR/k3Jtb7LKmF4e9Rhn4HDsgpxV2dWL2KPPbHZBeog+/u8OMJDUJZ1Wr4Ixl
AC4HrK8G/JtvzhXJT+Wgq4D5U/eviaQCiDODqd+59NMyAmdC4oczocWQGdEvdv0T
dfvkUm6DbxvaKghhtBgcgc9YV/W1ImQCeWERxO7NL68L8whpSfzm7dIQtQj4qHXy
jl2RcFo+X/ABuVcYQE/tPvZ9kghlnG837fYVLoAkJ3uRmLwi+Qd4G7XZCIrE95Li
JVl+Eier//ESOCdcIXovrzEbcEBrEnutyLtZnI9IKArX/kRbxq7Km6HOwesDO4d4
ezRS9tK8QoKgaL5In5Lk9+ws4WlBmAWLSFBvV1iDDZcZYyvMkfkPdpMfMxwvNG7t
LF+GcMifAR5rboYfUj60cM2AcA4fuGtiLYnW7qqE5AFOYUnXQwiN85fQ99CpL9tn
4WROMQ8tJsmO11BO74kD5EntzqIR+j4S/vGQk79/yyxgISWf5RrLxwJxFuenxQKC
sJQTnyYF8GynI4GadMIqZ6+TZ2YmRAWg85/dfG7VYB6+DrEzHdGD3cz26Lfj3JUZ
nVQ1l8WjgxXxXl/i8/Rq+iNyrYyj6IOSc1aM/tTwP3s+1QYDOyW9RnrN4aV+MD/9
BhtUpRM0eMjw5M+Rjf/b9Ub4mkicvg3tICqMS5YUBNDJPHSvI/qTSmtrneayj4mv
P3pfo2rNGp1XpiPQL0bRijlRg9bdaGlLMuoPAL/JENEN/wYYJHVXZ6hsYWcchgsU
tx3gxDUc2zOlni/u6SVUVLtRjvkQhfTKjEBHXTl0BbLyGt14PHs9Ml4TFbhZW/f2
wW917djb49AznvBv6lBwmKjONXz8Tx/wXQT3ltd0gKiw0GptaAXkoLpmFEtLnCxn
U3XQbFFcKtCR1AjRL+loWCvYrpCLLSpuhG+EatpXSQeJk43fsO7mlMx+NmkYCuej
OB9AqWJL+RVu/Cz9IS7m7G5Fa2LumpEdKBXGL+sfwbQPH11X8llxth/DjJ+lvaXE
HQ/WMxC9sNkjCS7vR0JWloUMcoJOuJLY+V6UPYSom0Wij509qIPpoHG+3Ze2nYEq
X4VVJoZn+q4J7rqIAtAAJT+t9d1uzLdmPgjjDsLVvlLs0Bl8JI5/ua29ZvF9PZS5
10w/01L1Yj/02go589ctDXsy8qvfruJiovDetYZXlb1AByak2NkwEVcENhhd5HaT
ABJteCJcG92X5lbjIx9WHXJft9brfhApXAVWX9xIcu9EvPM3fCqPpn87vI7xsDu9
QcnrLMTZNUOveF2ecgU/TyKGdos7rZros/Tul4uPOvmaRak4l+QfLkfi6qu4Qf24
NNWez4GA8bXG7Dxc2bjk0BDateUXh4OyWgqrC9/qMbI2WG5BGCNCqAuvsAkMo6kE
zKfzGTl5X1sGMd6kSYq1726Nv8ODqQpZ8NdHMLFTgH1MnXLvJO0jnZFGkATyobYz
agjr09EeFZN2x3qubG3o5sskpAnXiTAtthx0Htsngp4tuBArRZ1YeSZSDNNxIJm9
EsEXL94HZJX9byQPEdHmmhNbe+GMbUb062bg7O85WWv2wStuYBZZvizNReU2j7My
yrhzuGUuWG6FstlI2mIVKgWTe5w7iFPkxsdJNTVFDD8hAJPmb9QkKsHlgq/TJcLb
Bj5QwcMrxKrXb0KND34YQw8Y9d6MLqu9SktuHT9hmc3pFRggXL8b/IZ3aBRfdpDN
QCdgk2cnkxS18FJvrGY3Pg+DRD0uqIm1Fzsi0ZIPygip95kDHWfve1sL5ORdc76C
FYiw6yyXa/j1PFrwB36UZ90+ujuayiy/nDGuxyoeIZR9MdaFpuhBmawbONVKolPy
ZlIKqbNml5TcXRx0gbGn2b7qp5NnHrKbYWqqbPGkyF6wyuitpC8t+TRIOBbCTTom
cv7g6j5ojPwtityUoBlfXbKnbkC7aAy+D/qMuIG+kPPkRnEP5aXqo4RVR6GlQP1E
20simVTIESH5hDEi77+HfnE2o/LuRhMxFx6+gmsTjn6lc+Us163u9Ir7Ea4ZsgMb
IZHJXX0ziPzsxj0YJrFshfuvn/ayU0wmpg5iO7fHzIPK/l/hCjWsmXhiLU5/+JRG
zvO2s9ezOqC4KN/Cr8xfMaGMIf7BEgRSEZqBa8u8+rOuF/Z8bW1Jizr0IeANN/pO
1RLcVeJXdih7s2m5ThuoWmwdnKxZxo2sT5tWf1eAZrOIwCDWcD2EGUBWh9JM5W4M
nVRE2+EysxpVsaZ7UctcAET015bpSJ1XdwlTgtcM3rV/oCUKccfLz9LUM5VQiesB
RZ1Wis5lT9+UPJHIZ5Wydpi+J4QqanP4BR2sJssRpsGeRJW77BlLr+kB4U4SXAgZ
rvhALOu4vJnnKLbxkeYXrvpF1uWEXK6PCmXjtauVgkamidgCj4Vg/Dmt+qLcDWnP
F/8bu5oTSmK2Jgy78MbaMgriKriSMzMi1js7aDy6le6ikmThKS4FNcY/j4fVVg3J
bAXtdQpCaqDiOfncpqCvipg8JWoB/aNa0F7mejUPwy6ZmXjxOobNfOoeff8/3gSv
cXf1j99J5GZtC3sklh6SgwVNg4I78FgWkusvqWC99Oca58qTCK5EMSLpMwJp1jQi
YH6VajPtgYui6VgqkozbX/3eg9jE21To/qrcUx8UnIDMRZIFgwxsjnCdOoQpq6bc
7w8IfH7DylpGx1c3WFz2b49TA8DAd/L87V151VtU2u2AKrh1VvDr0Cz05V+jfmp9
foBhRZWya5pTLDohSt9w8JWuEOLqdkYCs8nYbWvJEqqxJy3CBW+eFy72SbkIY2Yf
OX4tLxQPHLsTtSJZUkXifss506J73PP/mWSCI9yZ+EVnu5DGNH6vyag1wp+QqWCj
nUHRZVUb45LMsRjSmfMUi+OPzQeBTdSp5faCilYb/8KuvW9acIzam+Fdeun5EYc5
Y6nxmMGR2c+vDNlmUTtG9wdv6MBRlpO3kkq7PTo6sno+eyUoHiwivgSo7iYbJJJ9
F0c0PRXKzanEPfjbj4L+oU3SBLoCJpPCKTy5CDCfL2GWjFzJjD0u3Xci9btddLPr
HykHc6SfahlKUczRTSBHGkPAvJvI5BqrcgSQcAJYz4cnE1tbYh4VUftJPXAt6A0/
FhWzS972EPEZNVE8B+0qWFBNKcgMffP8WuXWmwquc/uhD+sPlu8RIxcZe6T3WgOc
cjAEm6QBCCtv9kpnkzsoV4ofAmBPSDH81Wi8O1jNeaiV24/YdPWw6n1i0Jp0jttY
7lUxMVEoKXNAqlX1DuVXqxESAgP0GiIdvS1afOcDj1LIW/eXpWPdGof1+bG78gOm
Fkma2K3Dm90geZspk8EAR5rd16wYbkAqJXjHKr1AiY5C48gxjpe7TA1LRwKNxoXl
xjuispKOxnumEzdnthXRLRue0xnnlqj/slKo2O3QibeEuX97DbDtJYUTl2zTvCwk
Jg53zdne9ZmtsXJVSyDELCg8yLWCYbnKCces4pE+i+9YMBPMBGmXpRN3MXPh2kYa
/4Vt/xh6cK8F0U0d1JLhqf1NFgj7q6A7bj5iQAF0sLQosIehwlyXNSyCW5u629e0
T6c47qlY1yZaN65EJZOPYVP5YEi5YY2Xy+OsMbf4QJlzTJi0f5vE6N4PADNQY9G2
SA8/lsW0TQsQBqZzaVgCytBn+1ihUFqnyBdAXt6Jn4v5oKW3c6l4ggE3w8Od56z2
VNBvOAFD+su/EFHCdAZcP6eX/zz0AIjH/fFQoNPymL7TwXctj2fby7XT2VFEbEUp
sagcrtL6WQ+sd5btLqVDCeFEHN3Q7+JcQBd8CHjsSlKQWMWENbMmMwUe0AZSNV8k
IU/NRqeMjPWa9T+LWHrEvahXyqXWtO2JBnwmgfD0PJaJPw0Y+Bbz0W3yisxGOzcd
`protect END_PROTECTED
