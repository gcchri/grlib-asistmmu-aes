`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CgP4gXdIwtxQhdvIsiPJZ7yXFeBA1Ua2Yw8WMpCzj+U2j6YTnXj4z/9v3XTz/Uvb
OeXDQnA+au0VFZRxs4HehpMeUZlvf3P9cK+EZxwxu0D2CbBtnMloNoexnwrq+bkd
5/9Dd5WPz3ysXI8tTIKiIBRatVfAOBo/OY/L46cMbDisjau8Y31WMQuSaLbzF6gK
0CVSj0Ptg/KmgusjEXYF2/q7qDmSpS5h5exXeJS4HQNj72ot3kiuoX0eS5xlrQ0i
`protect END_PROTECTED
