`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lawv6AWAI2BabHjQR06FchvFzyaoZWYno30/9ahAhorwTvD2RSw1rCEBPIp0sQvl
Rcn85hi+VpNuvQxWB/q1mi6LDg8PslWnN4RyGcXDnXzJRuzvDo/mlZlsUKllPslf
9vcc+RH1Bbz9JZ4GBppYdQMaCTQoaf8iaAWYiwysLKijcDj9zcPU/e3c2D5CUAP3
SnxmFIkF0/9PiI4IGm45kD69/0kqVX39T8E+BQRWtDYKuAH7IALZGooCno7v9/y9
eq0NZUOprfLSdDxtmhJCMdtmiKti7LnHbZ8Z0waglIgBsOgiUBbDzILm/iB8DFMf
ulwSHXhqc6/Z9o1v4xUcxQElStB1vbbgZzsoX1Mt3hzVcFeJIxXmTlF/BEUd35On
3YobK/EH/Uph4jbrCjB0wpaK2iydneTspj+zNjJ5kwTIRwnAWV9nAlJYBdW2E6IH
ITssk4c9v2a2cirkUhE/BI4dCD5P0H6Mll85tQk7M5nP03HStC4EExv7PNL247Pq
QMpCZhFS6dFXWi6VGOVs/ugUmJnhhx80IDlZrdiM7KLihRoiCoYd4aakGZEVie+q
CbAqvZMtnjGPCDB0AHAHI2+1DoW7dxJt7GJHRuDQrywX8OD7ttWu0tuSKIf6VlmX
hL9A+dA47ck3Nil5vXyBgLmybN7inqUF0UDTMAqVaZKUp0Td+x9IiKEZz732ORph
rboOpvmlxzHO5IgUroXGkz3uq+rdgcMEZXQWPiAbtAb5JphZMKcpJ4Bv+ERnPWP8
Mc/5k60PAbVdESmY4t3EBMqrf7LerU07UzQe3s4fJhzhSuJtqupzrMos9r85wRQz
vi6tGqrGnpJ1xp8AeRzKzBatiulbMrSZUkBku82ylvxMWXCXx6TjiJKfGjGcj1RF
AmMiw95lhrZ1vTurAdrbQQRAMEGkUqjrDNaimjdvAjBY5kyiGbNCKzTew+bAg+dv
N/176I53cGDMpAt0TG5eM6AngRpH01rAtmJehHfmUoSQipR5GrFAPBRHjuqsX/zb
6uX6Lpmk14wSUd9FVvSLNJ9D0WcOHgHxum3qZJQp+Bfr3ntxjNqtgtabxnTOhpbD
SxjamyrgHwSoYXOWr6SjdWlPV0esHDpUiBbEs3/bWQLURCDBBC5zdpWL3cGZlOGn
2vManvgDoDsgc1aCFdu/t9arL1j7//1/mVJ7+3NBSIpoqseTsU/qY1gPU+KG3OiB
zFmOIupWeDk0C9z10qXx3YZ4EXoCI9uP5WHwvWcJINUZH6kYtymS7BNDXLHYmjpu
5KZdZ03asYJujoTgOUX3FX9QoyDZh9PxRQszv79xKC1YUo+3gOZPVd90sDTeU8Y3
+iuLdv0gUz9SEmsZGU19HYb1j2eEFvDDdcmhZwbC3omBOZ6lMo4iiHUQcBVbnPnt
1uXFDa04EEzVA4+sXPXlgDl4EuI3mp4G1SA5HShWflXksenhuZAZxyn/16j9e+RJ
57JNhrF2qpPI941on9yFoguqb9JJJGVOEPNBInMwQWKI9xsPBCcL3gHC1Xc5sc8K
bJGgroa6a5s3DrsLMGHnUwsQLoHHmN+nhcZnYSfaLuGdHJA87FYMQ3czGGLSH8tX
4yDXs4iE8FCBp4MdQSvXEqOV0dY88mebdLcW2x1Q1La+IH38fYEgVB7vlUzo4+LB
wzqm1armA21pGosHJV5lkgEpTaZUsJ9bBxxCEeISvUfBTVJ8cPYuBj9AWMuPZk2Z
rEoZF2PsZ9WX2259Ua4OUCYKKEkfdI2WvRj5gO5wMIxOFRNxf7MQfF/+dg620YkW
i0NWzIdiR/NXg6DtonYm07Uf91C9aWaHvbZmA3M06RA9S9DL1+gkmVlKiv10sjDx
rY4CfWcL9csaU7kbSzP7l1IO37TXQ2GH2vmJfVqbeuvL3ZJJT8gVAP7ujK1ZnxHu
3Ik8AUTK8KQBCdf1VAUUiYrLA1U1oXL/8xjMXKqV7efTUZt0HSFr9Q1Lj2uR74wv
wYAEoPxOGj3kkwaWvfCyEBVzyV5G66oKmb9TYV3A2lYr7aqDaIrFk/8erGL3pJSo
3l0lexiigoIz+mwvoe7iJVtE7ydwHoGIVrYvT43Pfl+A3s0NXWAiEJ/UvH9CF+yG
shQc5R1DVtMnJREKnwArgLyyiThZdFHOvF+U7iyfZaB+XySH8us0qxWOirm0L4cy
BunUYSPkM5y1ewFtR8e4Z8jIMYBfI0g1gJvr30s5Qu85mURKd/qoeSOOrBJGA2Iw
zeBsWedGielmbLpMFBNfqg/2TQ77yOoQ/m5pYV1OUaOL7i/QgMAdvz+m9VFiZzq0
8fO3K1XLKvxh3DniynxE4z/koWzPaabNWvZGJUR62NhD5u0OQDDJnZnVLYzbeRNU
+h4/+S+Bgi036KiEkVRe39nw1qwP3D5ZDx/ZaVQnjSeNcVGMgffqTNxpcZTcz62A
EN/h43wG6aec0rNiGRKsDM6WVfikCsT1DtWvT9HbS7ecK3/k+eJcr2pQDz1PV4XF
9irxuOLE1uuthv9XxsKTFLsuAdn2+Hlxr4J/FejWzgX4WQ37g3Ti3xchUJ/cDNUz
GTB6MDjYSOaO6+EckGyLI0q0iFYH/kaNMdkrjLxiHwGDZLqGjPyVVNK6HRhkCB9+
tUwjoM5q7ywTJ/Ij5y+rEm2CXGttDIfvE2iMfHCY0r6Uus+jIgtto3++OpECHSug
irGxlfZje9UwPB0RftMvUCQGLq+BG6g0UMQFtTAlfBY+xiiPzE8yOIA8WrENbtce
JTeJAhy2Qyfi6npUfQ3hDr/Pt0xE476TpEUUjnzI0aVRTGA+nVOWzUX+BzPBlfiu
H/RqQ4NGF3GlKG0AV78bnHB3WsVQlsQ8UrMWd253Kg6Ws5pA7cetSRsqauDT7oBa
O3bvlidpWmxKW6STfD8Tm3Ziv3EWEDwWu+G/7dHiIhC8frg81mlGxGXdhox0EFPQ
4zWYd3Mins90q5ngUJhRapRGx1ieaeNFwwAUn+5weMWgVGzlFddg214IublJGjNV
moSbeY0IsHPXMN5N/Msg4TptJkT2+OoAFNXr6x28bHJEk+tnW001bx7kxupHEMqh
IRaWqURantJ7TMPxQ/XKUg/M3vVS2goqj8umn8IwiZulIixFKpM9fJlvJmrtB/qR
gO0GOmQrHaYezqgJ/kdpMHz1CY7hm+1QX01PQoe+dGlEEzJcEVHiXq8f75lwitlg
SwBEfBJovzkEU3kL3hdTnRBdYV7u9vUCsu/8J15UfEECnjZvHZCXjC9JwMXvyhaU
VxHc9ZyTrcjufnRg5N8V//eED3WoCqBs1uta0+cR49I6iw6bfVkhkEe/dSzmOlLf
R/dOsQiDnc12SGaEiwkjKj5aqKXjA0jXocWoBL8ePZgEEixXS6r1rxRTbfgCp6ai
naGwQr85S8nAF8LJhepaxMPepWa9zf8pgV6sBDUDZhi4sjgWpZsU8P4IHyPcJWAT
+4zusrngH7ITN50+JBKGYUJOpetX4U4U9HuTqNyy5Arn0sJfj4SIYDMN1Vg1Womd
j5M2MKxPkKcuhxnjMAD41HFTgqHZ0p6DunLM6PKJinIxBsrcD5GIAsowXgnB/wMg
Wohpe+5G3PhfisaxEV9zK5ri5UhhSx7+jqUxNadWGOqO1NbRx/33e5e5UFCzk9ZV
Sh7f2CBXE5d7bTvGHJz5WMbuVW/nf7g6ZrLHrKkpv3YWnekT9EEXo24roCbR+S/2
0PH8RHLZwxf7JXyb/dAA7xW1F7tVjta2gSTRnituO1pAL5RICKeS89IyqPEPhphp
ooDWN45xj3+u3vIrjdgGTqUs79MN6q5Nk3RLy27fof65UBYOGOQmiGEDsFrWVGhk
a7UdM031AQMqTyFnJbCGXFlR9X/aRfV2cSpUZBVH4KS8tIyLLZq19oViSlrDCjPu
OboUt8wVQLa9Vh//gbyh1Lvro0e1oUbd6ZGb5/TKERAC9LN1/uB9puzE7qRM9UAS
4lEAQrGNHXcvNYCzBg7KQWXPZGA0e7mI+uErXNLcZT7Louznmkatn77INkNqzvn1
zXAeP2uJTNfa0jgi2ElMTbCtmGsMpaNV+zSanO9ojI8ey9/vsS4LKuVJc43oST/Y
W41TBeYJKuAP4h43Y76Pq3hN35cRW/poRqkErm9QYhMBBjPH7WqxDEduukm4hDmv
mtXX8lCXmfHbrOiN+ercqSN1IEd/gFiSCm8d5S9eC/kEb+o+0jbJwHUc5/1XofXd
i1RZIKWNiJx+iDWHNzW3AjcM3Jmu2v5FKRUcknnGmiK1OR3Mr6no3whxs6fBNcWb
pEWYBvAegGSY8ad/wklwbtKmMSz5vTEC7u3ifuZEntv8HkpVP6Z/ni8T2/hC7cMW
7RpMZSy6SNcGqf+E+SRX3Vf45MsRWFqQleNj7x2qWypmL2TXp0z3gSip+2OWV9L3
uhUmgVgS278+G7euHSz/vTh3Q+84t8tDf+U5KE7lKYWK8Y8jIKbYRN9fJ+4CnKWS
/SDqBmssh9qeLTxwsWTaC7I2cVPv2GNGh4Ro0w2UWh8YvaIk6LNTzIz87jTIjbov
aF0YxC8fnRWcKhhB2UIkEHtvYT5UiwUKcB/7IMOblajNdMbQ56X7V953kMpogXbE
t/+5klHwb6U6XU9+UNiDmfzg3RaCCCGme5NJm+Ahh8ccUwunAIVidamZS0UwCeqe
Zz4tBpqqrsNuL1GkfkimFnwyZKfHHS78vuByDcy7oYXPBGtmADl57cMNUX6bTg4D
ZOCOThzClFUnrb7WzhOitEiy9LZyNDRxsg0cvXudh/jNmbvg5nTK6rQUnHU+wQbE
XiFnPoMcidDx285tseeIVIqrUru8Ctv3StcUaqoilS1vf4EmukYShccydY9e3hkE
kUsp8svK8iHQkUegFQEKDVOcbZWY5O2rmXq3bnsv9Z27P+WPEvdSLZNlzBX+XykP
fBbiEWhBO45dAS+CsvuNvSqiq1m3WKQ7dewdzR/k5wwX56xakDU3uP1n6KCQC/9Q
pI3iAcmR4tqnLfeVZaiJNz9CZ1RT23jqgAsOp0gXufUoCrlOAJ3pDF691bpxl2Ur
YFVeGrhp+MvSWQvcCVnEVSVzYjqRMAq7zqVokE5q30TIgCpLR/ysxB9hN92is9f+
FWRxMv31vsFAfGdN7kG62c19SdtEGVs8Vm91bLiFWohdEC8i6bNJ07GEDOkMlWqz
AIqRInSIHe11SQTlzDuMviKKxg7a+CEPhNTnPXNZbqbYR810MYGwe+YUKTTuCU3O
DB/DFaAcuoac6tBZxKZ74qDeXYrsMnYURpFHDQFqvcGlPLjBz5OHGsAGd7t2twaZ
dqfsMbvDoHzx2GhdDb29AFHkqk/aIXRnwcb7ca02EGUkPji3QzzgBmoqWQxcI+ie
LJbmEhUlaGrce/YuUxZ4046+yYai5uruH8lCTMCQnyGd4sdLRo/N+FWd+6hDYRaA
wEuHJoWZTeR/DCT/WFA1YaVJOlH0lQgxit4IF9ppRbAgCBjn5Ybqy+RcTiph6qhY
bXi0/+5Jl7HFVR9jP+eFKBLe2C/J7JgdhC02CSK+6TgoXzmL2Ai7hb86/Q0gKvix
PhZuXbqbOCdwqdAU9D04fIwnyqlD7F0QP7IjSZ0BZvPOtdRb320JZbB5m48mCnqq
aGiQqXJmRAHMfG//sMBUVmaR3I+GPXnieHfIajyr5KYzNHBIh2oMA538sb6ZuGgs
ZUA3T4TfN8EOp1vMHHVecLGJpqyOPIoFW252ue1IcTFoAyl/6jrkWXe9aLdx0RuX
Zw2tILgbwmu7XRb2chvsdXktudLhYmCCU/LtwKPb8Ftw4wCyDRijgy5ch4CnPRWt
ldQDMG6Ag9ymav15+H6BmAF+lrQaHUxvqCy/EiQz12WYh7HbclpT0k4ZqFEeEEP7
gtmXptfwKIDjwq2V7v7rPw9J+OiSJmty348sD7QO+cgrw9fzyjOREPy6tUVa3rWb
ucbez9ezc4CNEDsak7vL7EMjFxXefr1cYCHGzoNrSidbVqxneQFfcoKuye+eplmp
ZiKUI54RX8yx2WcmB9Zd2QlYnA8iAtQ4S1FXCoHhJhzrqAxaCBNjx7XV0zuesUmP
75yHX650FWcczFCah1FXq2nrfTgItC4Fw4ss7Vhb5BHkCG59xbo01ror2MZmv6zd
0V+Le0lXCXlSqwjlG9B6jsohr0ysRaimS9p3il35LqaZzWCsrQ59RxUPeX9Un9Xd
OmNEhCqqgZx7eyAsIpxXyPl8u/jxUg8ZE5qmewqTyQyXfjsIAkN6uUnwJGzSFKVG
UhDZvnFpOpBnU4jDwFFvuOWCKPSoheZ4vQ6wtruRwkwTJDdmtCJWw38YLdhbt/Bb
g34AGDBV4S/FOzZfS4Bdf3/8hujT0PmoUUWCupxMW4z/DR0hFwup5inhTxhdh4hr
QYoIr1sEB/79OFe32AJvBE4QoIkCktHxBIXBTydFVs7ZAxkvudMWxYj7lATWDcII
/wCHd1tj5JqjSGtxnUVkSIj3eVLGzdVC66lydUuUNtkd5lw+QwbqkKhvU+rF2S92
putBjwLnq4jHjVzAJc8TSIDrQaeTKDIaI0T1vmyi8jQzY0B7AFyCmVn2zI9ArlBD
KGcbRhh69kWb2Qcnx0ecLVm2NUqg4mOnpnWl80B51GFbg1YoR+spg2tH3GIqT+op
At5L0rgRoPMj6oB9HQtXqWLV3BSN+8S94z8+By0WGwtp/nl3+E9egnV0QLuQPOZq
AVIRsZ0WG+mcAHQgPEg3u8eOsNxehLL5VfaeQ7+bc56taouJN6siSTy0cCuwIbXS
Hf1blmhHC5UHoV2vsPyNapvF4Oq0zaP+hsBb+e4MQgL3jIJ7ldojVZaqsVJRyLOF
DCmC+e700C4Kbg5N8hkOpe03wLNsoKm7rwnguUVuvOHZpCmD/0lt0e4SCDJCvOnb
`protect END_PROTECTED
