`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YeuDDDAyd3KmqWZhLS10yf1hrIwplF+o6PNzMG2BPj0kfpQOFlOZCHU7s/JeUZDO
ujLqVTLYqyJohnNjii2Fash4tIkV7sjXrcKi/V5G3eqM9X+DJ0WDJVJhuM+hQafj
xuU3KZKz2SwzEmJ3Aouy6HywmkG9eZKTh03ogwOTgSCfrZCwIqwNyR9HRE66vdXT
VKdbD4sqdIHy5SecYJDBnpBK4r1dKk/p83aoWQwrpM7gWKOH7DEAekuqf4m+mRfN
GUdp/HuRlGXFUFG1eOKCDg5KRJ+r5VM6WhcPzkpmbU0=
`protect END_PROTECTED
