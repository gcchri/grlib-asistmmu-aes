`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J7YsaEDIv1dsF5+6IlgHWZUg6HFSgbVDyO54k38UOcxBT+cfPRVx4DntoRDvxxhu
ge/2c/EhcS1v4vuXaY2nmdZ3Yqta8V9OPcrWGmx3C03s/sitfyp04SUgpnJJjDuV
K4RYxp5kWQkCSGZX+15KtYxSBiXI5cBgU+PA4MAXTmWnVsjxAiWnDoShhz/zhHT7
lnWhGC8JVds5dQc5q1OnDwscEbBEONd26MavWbCxvtHiv3Wmz9vcPi1pGxWg2hGW
vV5ToXAInonp0nLwBxr9YMh2Lh+juIhUAXp3ePYBlSc=
`protect END_PROTECTED
