`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CsJngSw3f96jU0E58EVNdd0yWitOiZat4CKuccV3uDF95aOdWglDFQ1zlROI+mmX
uBet++yvCDsqG9NLVEHVgtgU41nOR369/HL/2p3Coy1twUiNipn0M9AzTUgqnK4y
nsinMzmqlJ3lzALMpqqFvNpiNwhHCAG5k1yL+MPg+MMgcTvqxgQFLPNMeODisrpy
9snFO//oUGZk/l4U5qwCfMigxWU6pWl128HAwanLZDRyPk5cwDQMniI5tl7P9okT
n4p7+7DYxoP+g53PaQBC6Punc0Xb6KbFmUjX/8f3Ih4qNFSiA2Bz5sKNuvrEPVwB
RaWfJclxPCkPw1TEV/yjoy9zTocUvtnKTmqhWAh1kT5QZnwet92HFAS8wgb6I05D
VBguWbuTI9nAJNU9bvKyq0NUt4NWen36UlxkmJ18gIE2uP3cjBm6JUCe+obll/Va
fOqiePVl0vLe+suDgSiiH0k2ALyOvp5clwhLoPqM9GbEx5c8vus8v/G0qn5a9mle
LxfUiEEd7D8ExmvCW2QlpyfMrcMkZVjx4C+9gj4XfNojgOtifyoT5wfA0CXEuwJR
PgvH70Mf+YmcPdoZ7Msor/yApeQxx7q2sL8IYW8MBzrXbTGboZZwVLxMWm+4DHKN
y8fEnGAe7wd69m7i2knayW3lbqKCWi9Ucfj4Afzg1d8pAd7A4bMHZdc6m9wMXfRg
DiGpC13sxbRlGM+NWw51I3KHQMQYykusdfNdhmwJ6cduxoeCQhN8SgebxP0lykyV
KmgLyuOSHksq0iLSyrRwxjgPTX8+9aFwKfGR/5KWx2J4sgVrgywX3eH4nSnjii4v
5FZWxuO27Gpb5JKmgchaV9R2D4bgALW7iUdJvNKlzG47cvAfvytvjb5FG7KdB4Dh
LZBpBEVktsGcrLtCHqVRvNvaYynaMeram/OaJFmCJGq73g9IHIb61sNQ7l6ORyKZ
0Iw7bxrAu9IGVwTOvj6vSTmXFiI9D5IoJZ7l4z+F5EAxFkAbPsso6PrKtT1Lgffd
ZhCzgXPVU5hYe9bAimEvnroDA7CiB60FgcuUq/ImMdM/unoZO3WTjiK2Mi3J+D/j
lkxYTGXx3PkJwA/PNdll5nEm1FNG+fasgqJzoY+7iN0r79xZQ85ofFIz706SpLQ1
8UJiJMCU0a2e+mPVfEnKGlsqkPGUMG3KP6btlr9O8B68QOHETduxLn/0LThlwXeN
yqTJCnCvy048fY5QRqYid3kQbe0L7YIG6nH/m1ogzyCMOJcInVc2bbMDbPg5fOgE
zHbrijpFJvMqUK1GqWcavBw+M158Ud2QQE0MVLbZh/VBlnJTzZh4ycKGpT26YjKk
BxBvcjJCxNlV/dMG0vDrulJihEPLj+sFiXrVuw9tZpe6OUrqNS9YAIzLoghV3r5S
h+DgDEPzHLUf0Q7hTttKrVGMmiX563HV2uYtDP4ZmfqXOTQdUsVV0sz5olO3GNlK
pIAv0vsszh6zoSKXbGScmUj87xqOGPhEdyWbjxwRHG9/CW85OgQBv6sJv4mhxBIx
OUyPrkOkUOw4/r3Tqbv50SVAheloHrP6Ootb/h8bdS9XaXFNGtLPAjb65feMXeO8
aV1H8LvKhw/dPzgbptHTXDeeIERX1P1R3OvKumofQKMGGh/l1r65cSb5ksve5VNw
mSqqu6ClJufHdF7ij3mRBsLfdWq8bYkCdkkx2oUBvZ4XhnYZmM326CqPV2t8seUM
RK6HEr/dx19ou5CFYYwbFCqBunmGZry6UAJscMa418ta0/67nWIDVXKTePpHu9xs
ENLfO0j//4uqmEvyq0xIrxjRd2XUJEHAiU4PMd+HAnSbOYm9sRZh9axdKqIE/I9X
pn0XRrVlcBIR8s3TjCM8tQm8YTy9IzRK2bvrDPmsOUK27g3MgO9yknc50gy6XmcI
A/cJplCQgMEi1rm8R9CVKTFuHip4ckjOPy9gZcl5uijWB1UIF1+lvf6Ed9GvaFSG
0Xg76FAufhy/kz5NuVJYRLR8X/5+obSlJRhCzEIsdZ3B/VpmGbvtVAe3Pazm40Cm
9sFKnWZOhnd/pHyAzyNv3uhvzDGKNi9q8cMRP4m8eVCWIfCX7NdG8fpih8qmdb9I
bDhLvCAKgSrR8CIeGj5cFVJgwqgXW6vRfM/P6ysCy8aLDWIHRtAy15cCg8FEvbnF
o6lccgrKADk6sZB6N1VpgptHDTd0uSt64/7uxCYUrrdkxkmO398CJz5iVqCrKteu
b/RNr6vmv6iS1e916i2pRG2B/5xJVWS9q67WZ0bP/5HViasYeFIxy/r/caPpcLyz
kkb18+FVSN+ieRKfxtDm5IvV9VVPmox8w7SrN2RKoFP9/TbIoJxLahffl303TWZy
UDfNwQ5xsiAgR+mn/Z+bu4EqXQNc8CCNcfJLbKruUYqkVvo9Pi/dgGVY8sL9IVEI
T7NDbsHDNDM4/ZKMHezUC6IKrESrnk657uNCloR8wOhsd5I4Sx19Ouqo+Db7WK+R
BkQ4Op0eDEvInrVeVTFAeKHsIDFOW/J6vb/noady/CPNrftUYAGOOetaGoLbduy3
pdTAjU161jr1xtuP3vIMOci0CCsIi5DiNmrPqcnBnez7cYhgVbISI6k8PL6lFAy9
OntVK3TFxRV1x/Vdr5zDY/QVHzFSftavYDPNXpOiD2cmPTp2VyEHKciekRqnJKB3
1+w3j5WHtXF7iQsFaj6Q5B23MQuXDchTJdIcGQ1YaaEnhqEiyMt2OVtWiI7I6tvA
VPEU3xgiEAGNY7GUvekAnOjxHB3zLDJVNjyMfGQe3rHAsz8EwM40yzKWWn4hJK0Q
qFs5wE0s9y3IpxX+rFUSaRFrMWQGlEM3grPxynrQSGqLpZGcsSIJpLWI0yf3FivO
Qe410boKuhx28F3kIasJ1gCjTTT+c+Brj4rwiicA0vIoNpYj6Ydz1OBqU9bCBWXy
/9f2QWKO92a+WkryATkMa1NWIcRhNG7gG9LYzMngcbr3XVOqTJJ2LmvYaFvStnMH
M3UjJCB26owWEHKRZQbw2qZf07KHAg603lVQ5xk0MahcV8bPDDAWTqglTES178pA
Cy3+Z9yCzclE9KuMHxGOP6g0tCFYcrwytKYnDmz4GqulBiDo2cnpnx4kJK3fmhKT
lO7K96QT4eg1k73vppw0ZcLDckQVyWETi6TYIOzkgHsjQkI4z4F3ZYcVg+CWFoYP
Mkqyi6HBQAq5r3MpA0VwKTZW3zXEUsuZnfT+Mpjj94E1OAt5Qx9iBpxR2nHh4Qiv
NR1YM567fGvRV42kx+2uA327Xk+yYRlaWaojoIg6yPSMXU2mPFnGv/cj32LHv2rd
micwGGvNG8YVLDOkEYJCOjlvQkLpwDYTUi8sOHBtZiA0lv1eKdQ93W8Ma8dJUpKY
h7rUE5gqkijvuI0w20hBX+17GoVFJMRXpSaOw5DZFkr9oh+wWX721hlHolxWooXe
li+KRQwKXxNque++uaHeAhhut8XcbsRdQ+dxOKHf1IDehLKWNTffM4vRw3zWneRT
zD6PivolLk6Mq5UhCsjnLKSanosBy3dZTbgxtYiQ8rzf+jAidZEKLXNNoGPspqT+
wED6xo66bSQ5UnqFyaqB4kByJFbrQD6YvLxSZaYS9HYBCskSDh5DwjdYj7GwTLMj
6ZVzNb7XA/deznSRkv9TzZLw7OXY1cClBLiOTZPwT6w0hI0QGaRONey8JJGXga9y
VJn0ABqYfcEBKO1TwcB0ts07zEkr5ycjs9AmQFu2zsrXV9gVIwBeIaPRTISpP8yE
kwKv/H7tsuLXCnu8e1pIagrvpH1SiMXOvnhLnQqdc2NMtnTZaOjDMKuwYtQ2TsXu
Yuum9TBs/aHfd0g285CaGX9JVQj8JW1TQ2gARjTfIzStnc1H2GgpqGIQwEqYZ7L8
GYdmTjaTcDdw6K5Ckq9lnXCfM19+9ZJZE7k52xrF9OAlTwDFcjj8fYif6Gn/Ea0b
UIhWEAvHFlha9YieDwMvjw1y9SaORzGr/zVS3eLtUOyaNG4AOKUveqJ7QCBu3jrt
H5d3YXDSIkrl5LdLSmfqHTZwgJxB20T1IwIauPC6eHiWxruh2e2ma6uxe4wifntO
Xnd0RxGFf6dXJrNu9sA49jzBvo5CrAdjtKzTcAt17vwOTXjv6TbI6oaqsYi1htY2
NCfH3S1mIFu2HqmD/A8e62E4DmFh2NDGohmJnWLmHJbF+q5lvXtOYhzyAbVDTYJE
ZwfWaT9faJLMdMPB/tu/Q+eKiG2Y8SxAfkT9idamOqXTjQ1FonCB+WvO1UwDNVYb
syJc3tJk6t1vqi6rzOl7baSxfEh3rC94stQDJ7uZ3XHq2R54ar00+pq41uoMRoTR
Ugq9L/bU1UBE88h3EenQa6zj9VqfND84B4xe2JQBJYEkWcchcZqaMsMQ2UJEJoJM
EhPm0XwCIeIJCqtN8M7hoIMluQZwwPW0xwSKVhAvzJUVkZsHnadVuqPPKCJLEPtQ
dcL+Hh1dnCXiLJPmSibyLuUUY9pzh4C+AzyNXO3OcImz3230vXBpuEctJTzDlspN
mbcYEo97OH2NpXkU7XAJ7msTMWrRTMqwg5UbQWXZ4qsKuunqbMMzyWe7PqEvZq8W
ahrh7HQpHVCDlIoxNVRom8wxl5Ob+i0pWXGOoXdtT7ytGfBxtLpUvJ1jDqwpKH2G
RuzqUMtdk2EeWJl6V8cPtq1NeBu/FpS1T8VWvQXTWxS8yAcrY54soega/b3bmBvo
69TyXh+Y5lfMKkYGMYTBLGRS8BAIfPHuM0RkJLR2rm3ySPh95Vkkgxdl5SnhrJBz
9meqawe4NQUDCrKmoA3rm5zdjN8Fqu0CE26Mxv0JUIErv+1oAlkBOTRtN8QfOrWg
aefiHm6EHCGlsThcLGa9IW6HAjcLlOw2/O8EnSLBT0D9YetbzW8CYIDjApfsDcs/
qKxNrnfsTW3GtQ+KMCWkqOWoT2wk4o3ewD7QwuRaRvuMnxwx5zywHUgu6q9eA4bj
zKLKMpKf4GjHuLVm5OweefMPkaG8apVhqzZs2njCRTgLmwR9O1pwzh62FmbvoHdP
V6u7O6AblqyrDJw6qEHOBQt1ztDBhHRBmv1bBaf+Yah3nL7yA3OCV96lzIlsCvrx
ajkQhQVcX9GyyD3nSye1tqdwm5/fsl96Vxkurtt7VoW0oki6ZWwBGar731beTP/k
IF8jen8awNLZP6Ts2qeL+Lyew9ZAT9GlcsaAPtT9NoPmQj8AnTqE512TYqGWwS6p
yokVMl89D3M+mph09BL6es57CzwCyJIgOp9JRSlTjQPr0PxO7j6DCJ8QwYw92EA5
aE9eh7ul24xvASp4VF26g9e7Kg5NJ3QSF5KhnWlR6F7j/I3rDTWKJPkofgnzQAE6
abyyEX/6wZrnwNnIMcj02ForJuQm/Qvby7acFq8eBlihQKovvX++HYdrAeqoZA/f
7xa0Ivmp13HW7drTMg/jRP6mTBe1QIEV6YQd2x4HzQMbZkURCim5e/jODSacxe89
SbAmLw2oUmhYTQ2YediL7eAtttJP6puD+o7zHdaqW67L17QdtZK21jP7r+8VEQXM
h/oVMeIgiOEWmKWHzWj+FWJzPtL0qEUugjqRxONhhg4ZIfJulwl3EZJDD8rLnwE9
YODodJL/s7a32atDvOITs+Sj96cwpsw+qNRW/Vi88uK1NmO6/6VDOaan9+Pst18z
IC7dCo2ANpjeAXxDBeghoan8zVt9GSsqswSnzjgj+JLZ30d6tajsH3g8lubLgWMu
CVZEg/6LXnEUjWx71AtuVRzRtt4qjHb9lte2Zf1EesqCr/Of2XGED+KLXnFx5XIE
NuxpVw0JR2WQqW7UKVVYD5DlhSgRFXEq62a7XWc5azfo2NrsaYsrmPKFscrzt+5G
oHsjU3qoFIMCyq9aMr3SxXJk1Wc4/OMDaz8mUQ58rXSe/6FXWpZEVbhM2/yNsMvB
9QBY4Mo/rXM1STtWcajo947HK5hCJms7UbhF0vHPYn4U8MRqAvpNMqqHvRPBUmrq
bgWkTZlx5mG1CpSKKvR9v3eg4AEH7Mp91fbFKP6qlhmLY9BhKiXi5vXQP8tgPqM3
Ae4aBePtticSApdbx28dvzPC2cn29e8Mk9K1A1ZoJn9mUAhPkGBxqtA2MCOQvf/w
PVXsuarPbiNHU6SdWNGhdl9T5re18MBssIHkNMDsNXpiVbHGEYNaxO9ST1brE+KJ
Fcsu4cGJBig9L7eTd5NwIRGJ3PNqHNctlZ4vTkHu3vPVEvF+YOK1quptJ4lCukkb
xmMWyEXe5Mtz4nPVLzeyHN/91A1H2ckB2LvRkP3FG3/D8ClQcIYT/AOIZL2n4GxL
UzyaPsJGy8C192EBulmhXy217VpMElN6Q7x+NBgOR7VEMwGglUpJ8oZFxxMfcySD
02D+Bc8sZiCvSlsKkweoEVwbWE27hnODSJFUFbSOkFblkzDc9iUpdeKIu8vNj1Os
HpstLXqLLNxzRqsQHW2GVGgWu1xZo2o67T7Cy1jkAizyVi5HwuhVaS3wyxi9RS99
mn2uyofneB8oOlFLqy6BpcOpJIKpq3OwYcztejoiq/EirJwbsiBke/NwulYOR/8C
pdaoFlyMZmG3uOlI/HQOdnlA9Y8oKwOHkFwSfGyjPCLwp2vHCth8rrilNilNHjMp
h1Siu71LazwZXpt1ahgiIFo1MJyhxdilpBPibCdJ2wLe/LKtsyMYoBPBBKFFEaIM
upAPOkvLG7uUhjWbgmk6eKp8OSdduA+TKCHzTwodNEEvOb9gO0Dh9PHmqLxA86YB
gMrPhygTCywAsQYLJtGMDeNMk1HDbqcO4TdTwLwlUSmJfAq8MbE/akuc8yaekfmi
mCJ48jloLM12I8MoZbFvMCPfTmvbw/w+eDKm5QLxxl2eCv5SsS/ZZ6hmOPkY3tAX
iHEkhAi/TbWbCO53Gd+oPtjqsO2pc1F1EravZ0RHjmmu1HI3llAh4h+Xa//fjSw/
CAUEvpI8WXLyIvNjK2OqhRjIgVF1MN5XueZk4ZFgpOkAqudfIdVDzfOuFyjYvhfr
w+Mv1Zxvsw5faMKP/WJ4j28HgPtc/yM1+FQCqgQdIMJ9czdPMlWTnuVQTPBy/mB4
D2jggFVsV6rmTH2i9uz0rDk23kfC5hyEB7loX32UjqWGiYycGvoCZdL5HNMTxWPA
cWqKTEX7wY8OeHsiDS52V/LXwklsYlqlpAZiQUQIFWvH7VfD1UZfyzsvchhDAgYK
vwFCU/0UgKVgNXJqGIJ5R00Y3smEvY+XvcgsNWxIq1Oe00Npf+l5YUII9/KkLZHI
CJTrlj1nZkb9DpHtfVP+3R4fA5Eg4asQZRD3bv7rSJDI1MeAJrUbtdTphlPrpEZD
BwHJc6WrgD/ZDp/K9F6El2kfisFpKzOcXUUX8xAEFzEtU+/xj2uBt6zAz8wnw2Qv
luFgRgCEbUgOMW6i9H5sKIJrfs5MfFQzxt1teoXeWz/G742at5mkQ1tcXncF4ak8
428x6wdMXGNkwG670EeFJzsrxVCf5oUy9esS7nEgInc7uy+CFcyjOcW/iVNIBvvT
G2pzGoEy49fvw2o/zzvRjj0FeTtNRmMwXdaLTWVEI91ZT8Vt6eSD11V8rMd1Cruc
7dEzWm7bJQ0Zs+zzd6MoHf+kiIE5MtNpkV7XQwHLAfchr3FMlaHr9hSYC8Tlq20s
wE5nydnlCY4XA9JuOMV5a6p0PBSMBC/fPLkhD9QsxijDRbXZKwL1dWzHFlLaNHl/
fivHhHsOPG7uMnAS3TsA5pX8pWd3pmuBAXdL7m+FwihC86GJj5YlrFNoIhdwwNCk
dFftZpDsr+0bs+PcpPr/vy8gkKOcCJq6WUJyKqfE62Rx8mJbskl38c0OeC64nt56
hmqagjpEnhfuCrCyztwutupYuf3GH5dj4IVwGwLXDCEFzgMcKCtBxUTtoT46Eri9
EGjOKfg1l6uP0xsZb0aFgsx0f3fGLluIxPIhGiHXwY7J45DvkrnVWuLzNOCICB+F
d9caRsiK2iaYpG/6rvC9eYp6Fgh26NyGjJ2rdVah56fLOw0AYl6Z+gURywa0dzZ4
vWOVApAS/C1sfggwdjnZFBMHqRuDGt2XlIXbLk/rpXhhZymrDi0qufteevRn8M3y
4TBSHgs/O+BvpMJpaqIHU9F/dHaGZz0S3ne8Y+ir7eLTjiQGewJFF3Gs9zFBlQvC
G1cQ935g/J9NHKS3rQ+AHaPKu4Y2YhXkVhT5pA/BR/hBGAXnV1VZZE8eZwYzLFGe
V4AHalS/AvyX0LBB5/1IIA2nr5p3n27bGpjdSciDuUXnBc2haaDXxhTc0cRNy9xg
/QH9Vq2DmahFlC06Illp8QSXEwGB278MEzHczD95x1wVeye63yiuU4SWSbW0ZcK2
whED/Z6hnyscQ/aDDmF7+TGNiaXjNRhO5n8NVpqOOesoliMDR+Pvv7WBI80tsvsA
BTw7x2FyWW1UNU8UiEOU6KgDzH/rX/dpbwwhdOI+D62mkza3U7WvW4cowDCD4Tid
f7/vf1L56Po0mQX66FVUB8bC8EGs+9heFLH4Nw5uwtOlJI7nEnCLpwxznCuE5ojB
YgzjZjO4XY4nplH1hvG5Pds/3kkKJHFiqW6sqj3ZS3JXZOQjQLJ0Gxwh5zEw+1Y3
9XKEy7omBHyWoogh2tQQE9ACDik+i9fEm4tNRCP2WDGnd5c9AabhQyC8LQhfPvwB
b4iGfQG0BCiZ/mUSvnKBxPz487jIcffbmIqWNZMFC3nTUSNvp5UMkXyXCcpvQ4aG
gX65XZGf1Ol3gMDnfWcIHfZYYK8fuD/HZeP6nBgQybpUWf0feuWWNPV1y0+nX0sg
g0RWD5bddCmsSNY6XNOky6Y+xVRgZVB+5yhJXDxZ3LUwlAkcfh8jEzks0paGaNV2
RL5cdL7qVxPqRUf4DazTMmXTsCtaZCfa2d/Ezx57cXoJcQc0/LM3uTDYDkTywMS4
VhEzq4aM9SA5GQYOgYP+g7/l3V6Arnb7qKIQqmusAadSFVwQ96sllDS8cfaAf53S
rE/pSND32ygFGuSCwRUGR5GP0VrC2zn7R0KXVtM2MvnWkjQRjzgcHeyBXnSEJh7X
8Ai4cZLERqz8tWW96D6Q0a+C6wGnBQ28VUnBCmavfqMcspVCmrlyPrAW1xwWrJ8T
DD6vPACP051AQwqBnL0ABPI1+oI82CsoJgbz5y5wP2q1npWI7Y/Ebbe2HF2s7qxl
rk90g2gk+MnpVLWZb5dKGor2BRWXtI6rqAFF1wo5aEHEaANoe60wYJY8wnFpGi99
M17m8Wj17oXlgw1T4gGvzEUZOtSdjUFti+ULF5KvVblKFFkH/CqDOk3JIjM/R18C
gmQnIfvomGwonV/kdFdbPKAroQ1Pp1fM02CBT6q4oQWxQYkD3GWbMXext/ltEbDZ
ApWswWWps7u1LcpUt2opl/+dObtMgmJ6QMnAPdDiey7wVLaeq+FthvfbbfSRlLM3
d7rYdrpILVukV9U190yR0OzU6Zyi6hrsR80z3ME2M6XKBgyeeHCj5GWLSIsAXAfB
5LK172LC6TjcHXvssapZJTIKcgavV1ND5Hm3swpy/oXVc9VzSo+Cfzma9ILJ/E/t
oux7JhI8+u1YMx4h/4I2NNBRHZfJA/HmR9CurOHNGzscQPT6jX8L//aPTCvRR3ZS
49eJUR6nbHXJnlLvHF1dqHGGuYQxWCpHMD1L/Zfqnnr3nOYTpkPPH7G4Hm7lIyea
trFpZbD8MQ8eeCs2Ho1bDn2mbpRurZWKe1xGGqQ6CKST8t/ugVSNggi4Y3QcrlCE
3QodjuG18lNvjAbT7niJJTxaU8NupEnJpIWx2NKbbGxu7AlqJrGxxD/1huqs1R5w
lBYTWwJrR0DmzMCs0EIVQf2wlCdngbBi2CtVV/j7CZEsD1BpaLJ2YRBMgpmyv1ZX
fLafPZa8gG78i7WLD8qSr4Fx4c0oHhwn+PQOn0pOIknRRsF/dC9Gepfcrv2/rM1B
BuAkWolf90wPUUWP5xxfi4XQ9KOZheAuyil1YHghNKG04ziAaPDTbe1u3OCEp/Xh
rrq/FN7wc2VYQ2X/7DR07L3HK7rva/llFgt84e5KRW0N2HPCdgBvD5ulNQ+fHd16
ThPSYSLXJ8ETV7HJHgyN6PhpjhmfEMn6w2WV2f7t8rW71e1DlCTdbGj11zSe76Pp
opWICRrkRZQq72d9py9sEhYN6/YKTxLsCOwlde+3+0eXdD1kViMdiDU6X5A3PRfo
QIkBsoB1QwR1Pczed8rvoQ==
`protect END_PROTECTED
