`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ajmIdj+wQ/w8sCiwiXA5UBYdUZyFIbkBdeLD0pHi6kbyFugFel6LwlHcOQ90vAVY
k09Hi2nqFZqhsUhGSYBloSzDGp8LQlsO4i1RMvSfgKt8b4yYHO52ujn+rkqt8N/y
eT4chlLWqaf32tNTzNUhtFewX1i+Hx1LcSSpr/Z5sg0xU+4zlj2QVnTtcQZxZFM8
1PU2zXWlOMKzLqgLnowUvvTEPYnYLKXKYGwAOqNj+k87uxMfrJW54vG4YdiAfFXL
ULP1X0LfJvXfL5/S49TqHm6mV5/SpeOUBClSM9FllX+mvKWhBnDs4OHZQm8Rx3UK
JPlE7/NqaQG0ormi76mz/JTKacm7DTfxkxAnYpULe6XjUuhpofSLQLG5AFEiOUqZ
`protect END_PROTECTED
