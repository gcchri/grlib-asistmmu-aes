`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+czozf/YDLkfvTxp44o3jAeaF2JnPHTeS9EVul6KHXrgog9dGOC0qcDb1vYi0Upt
cEvawidahXnhGPKGFN622YJ5FXBq+6vPKvQfhgLsritMRzm2i+D5jf38LTx3RaVU
OqYJQHt2P0hPa+OVCnpP+PBuVvARW2UJ71/5PWHYBLwn4CCUEthgMt8baQOj+HLa
BZ31HtLevXn8/+Ub/AizCr8CxZotFnyFKmfpIgkTxwU0LjFoCuY6pHOJquFLBG8Z
ZqFDnjn62AXfo8lYbTyyLB7JMKg0Yy742Z4gfDE3TaJozuB1twCnR9PPxQDH6DXx
OmzVTeqj6ZYHZU9UQXLIoA==
`protect END_PROTECTED
