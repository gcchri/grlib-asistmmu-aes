`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YFWBd4oymOIp/jy/nkb+SosE0iJ14jWz7nXl3qYMLNo3hSRiT7eELyot5f3QY62F
mpAbvFAnM4Nhty2GReSmxN8KAPcTP+VqpC8FZqcu+rmB4FUq4gS2LxyLdKNH+y4U
862nQDJtnvrkqBPIPPzCPGssZWFQ+OgCv+GejjDbZ6DVeZ9KKjlOs7H1Rw35qWpO
J+yd3RMvtXStsAsffGVDoZTS7OE8m+oILY3w5g7EFbcJ+UVTZ+4pvHyL4lAEe3+3
U+MKvwqO70CNeGaY7pfYNZd9isNikgKzFhtQ1IIF0KcO6HbR6NMnzcravzqYCxhW
n+qdoHJZdzrUfjUbwHclfWmXHrc5ZXu66irw8wLZN4azfX86Bm8XEJyi3v+U/YM4
5rqpQUUgtfw/YJZaQv5PKycfOH4nNtWBopqw7J+Kel4=
`protect END_PROTECTED
