`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
utnRWOUg8dM437G7UaeP4iFEiMgrj7V9YaXNf6Dn/SwwOUreImwnRarh7uGPl3uS
0PMue8Ze0YtdvJ88Jg3Tf83wrmwxMWhialjoe2jkDxxojrTLELbgnQ+DfhR0460H
G3AWGCEAQoBbcR5Q01auLUkPfya+h0TE77CvaGFR6CxngbWC11Kt7x+wn5AzWSGN
rMK71sanPB/5wYijxf5ChDsFYVUA3iw2pE8EIeNhYtY9SAgum7Ryzgxiu51r8FD6
37Viu7ufwzHnbdq8AocX+PteKGLHfxGMiVEIYAHgf/d5Z0JOFbZVqHSyt1l8TSWw
oNLeD9yX1wfXzoD//c8TY3D6tr2CK+c5dw91Hy1Ij4Igga3/diAsQAhxa7cGdW++
maolQcXGwSs7ZbVva7BoQyPD6jNO4g1aJe4VTDOxMwQl9ExCliaJBQs8uH+gEdB+
GlJVNVI9NQnhdfpzLnvE+hQovHFpK8+JFXfv8Y6X2mQGrnTONkf991HdAqR3u6zS
NLEB1ly9uB925k2gWOLFrMNx4hW3nrqdNajEgu8LYVDqLlACPPm3Iiwrm3uBEcE2
owSFqCcQyUgO2XUwYxPydZmOgaYw1rDXUe9nC6eiQ7mcVaBjc4OmO25hJioOOa1G
m6DwFYiQUN71k7Z8zhc/May+2GeGxm/JjleB005qk1BhGDZwza/GWNlM5IJLSMny
7uP0xE3ttwDY5smL8zWVIPu3O1cERZzrrC/3f8FaQZTjKulaMMHnouLxUPsOd4Zb
`protect END_PROTECTED
