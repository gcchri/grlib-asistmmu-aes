`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F9Ce6HJ/x3LIX7kegQEP6Tzys0VR7jpnJTLBkpli3eNwiC7btk5kTxCCWoF5Pu2n
/KnwNyczBJP0KqIFaodIb/biEeuMrk6T6f4aJN0clZ5cfAxmVj4IGeTkhJRpzWWp
nwM5EK93pxrk2bWSdWeCNPBksdQe8tzTHh5ntEASLzXM1ua2byDDJ5ONeY0UEvki
rPoyO9cABmG4ndSOkAUC0wkFfTGSO0+Di8xIoyRj2w/R9dgRDQcgxCsJF8jDwTwo
faMgtcgz2uRHOAL5fmBwycJZapkH1Z8fgg0Ow36fjgJwTY+DO0lIfcec5xmVpjhB
EJRX3LgpCl6Bg311x2fVhHE8pgQglMgMxbn7UXbwIFLrPpNQvPXePTcRqQLk24vX
bD/hWAnHXYh42QgKAu5bYPfyKBiK0PaFgo94kK45miXXt+6pMjQjDbp/webx3gYP
Bz17KQrR+n4cfWI7liBEs0Ne9pGUNFJk8xSdpAmiT3jAJoSlzBC/qESehwFjLS3Z
n2i6Q4yCQmrf4wBK4KAL6YuHFF8nxCMZJCo4d9TqaWtTTILS8BYZ/D6SgzgsTg3z
ZMfQY9DAixoK+rNhi4/iH51cyh8fhZzwRgwXM/zBv1Bk8ZQDdw/eolMKtnn/s4Ff
RMcOQSpC3Jxce3Q3nHpE0MzBiWynwBW+/ZjjJK6q/qym6YsnP4CIIP5saB8PTlOx
+RcDaRKYBQPSjwIwYdx2RbRf2axo4D570+h51LH7AdwjSx0OB+KzbLHQgHSn+i4P
+gLPrknsZSNoZH5hmKOZrZNl77QI8oZqGxQT84mTP02Ss8rlWRtWt+9QH9z01hey
iTjIronOgQ1kNtZKopyHoXU1w+LL5DGqHc0R1obig3AtfzfcjXpKYAZSXO1rht8U
vY5qYKDZu9/QsgKK7WDebPTKOXJ5POu7vy4UoARO1gEjvtg93sg1zeACtU+oOnUS
gOvMX+JY0bjUPnLRVj2ToU2eFB/a5HXuADfrmySEQA0/NDeP43h22/ueQlWIoYg6
ZMFECRSE0NIQ/zXJFU6R/gNWyyb+qJFZ/vxsPg+ju8D5q0YPWiOnUJlO6q5VhQ4J
tX7+CLRDq2PhShWtblUTwYUXpjqsRL8WQGkrawN35AsRE62hFcjshgL1MtdusOv+
KpEpgqrkyavniWmLUkbM3WWSSR/VhpmB+J+NWGDWHM2bxsXL6+0lBrwoPtO8b+PZ
9+igWhcruaOCX0xmvSdtkQK70c2j4gIphN6WK1dmcLUVoAGcUilfwnVRWKAhqsYy
Ahmy+pYXHFz2fBK6LbKeR6LDiQdnT2NqdXZYZvWR7i55baNfWA0ZTrOkoJe3AfKC
R9/XEMYv3mhIBCGdW2+hK6XzhpDn5/8cYeSQpWUysQBvTpmJpQOrNP/seYxpaWvj
2o7ouK9EvlXJ3I5+WqbsrC4oAHbp6KTVrQ035BhmEv73Nwb1QMCkT5MRNFPjm9H0
9RLNtggDGx4TVgXtljk2QxbMI84Y1ZueKtOdzl0ZY+rtHeAmArLwPOF9WW6E7xrY
h18aEa+yYARCMKAvyz3dMCbayd2SIg6vMJBDHsf3/lX+yTwUcCdkZ9Ea2hHsPpFZ
AnUAXsJgYX46Cr3svS8pAhVLd7CN3A6YyYH3pYJBuDkwiw8odPY5TULBkLSH0+kK
u87Gu5FHJ+X0Zdj2kVw9qAY/Oa9iXAyFalVynzqCfTvAAyxShQOAEM0w7NK1vT1D
B+WkRF9ilb08vraZ8ayB0ELDrzeU5qeL9vjWDUpWPE23h4lfxrgPECUXyCDdl8DZ
QFoQ9dw+k/7Yns+c3V8Z1g==
`protect END_PROTECTED
