`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x6JDs789Sux/ki8L00QYL3xr4wOwA+p4AR66LBtUvh1E/vb4R2pjnQg8xgI+pG1Y
F+99o8gHqwCNgIUEbrtxqgIDrt1b9EyuQry9dTglvhnnCqxelUSsoTbtiEdy5xk+
bpMTeVpEtpWYHBdxqhieh0yIAdSTkNS8VO3XP4zOOpjQMNx7kBVRcjNDfUBVUvM0
1X8YtO2BG1F4Zwyd5EW3y+54sfFeB11tz1ktAg+68paKJykEmL7kKXmZ35a8KtKO
XNh+GxW976vVKG1C0ku/j9EMGtVriKhX/AhsBEjeYObV6hN0sO3BUQHCMNZlsgfS
Rr/SNk6TAk255PRbyslk/w==
`protect END_PROTECTED
