`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8fueL3L/VdyCZppySkxkd5pxOUahnLQQyNo5dTV6Al6TV3QI1tMGibZ99eIXSW6/
fvqmzvJrqgStL8yXIVtFKANkmxkHRRx4NVWlhid8NuFkf3o7znJjZbE06cTm2XPn
Fd9k9uiMiluXTMmTaZ6QaAuQ5KpqgP1AMgft0xtCmivcp2CnOU8NWbnBBfLLJI5W
qldCNkkvj4CLvoumlxvIZt9uLBmR4agWoUxoPjwz/jhv9DZW3CMN1I+sA1q6CAOO
ughF4bR0Lp+JVKR7KyR4sA6aDKSkUsD5iySUN/Nf7zTdpogoZXNijLWgyKfiT+2Q
FgNHrmF4wThLAPCkdeB3hRZbw+sBtV67bxSoa74hY9gF4vGW984c5ljQpp3Ym6cQ
WiFLcynB5As1oV7hxtnLEdWyAXedLbvZOgkSD9UpGVjd8jAM8Zr/LKScSOHxMr9Q
pKTlIp3gKRaQ9JzFu39j4I/RrEvJ/rf/VbSAloEbMXJDVfQ8mpipKBky3X6twF29
N2lqLwhq25uaMLwZEwqbSJmZYpOaOSWWbk9Y4SnaHXiNowc9QAihTs9jnM65JxFP
gXKeF7VweeGgtUa7zKkPE5HhAMQCAeWUGF2j4/vn6Hs=
`protect END_PROTECTED
