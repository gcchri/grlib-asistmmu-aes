`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lL05ayKDgG2kSMqfolF4bsqBBBDgN4+JwRSqv5+qUFxdY4O1UFcY/mi8y2nI4y46
1gXMpkF7O6eioF7++F5An/tN7PytSowynQlr+EmOXdP3z8p5hZAtx4oPhRUAvifv
4y4HecQSn3F1IAOO6Q4+LG6tZ7i4Vv6z9S2DPS2+k6ijOeZcHSdMVceaJmgpF+53
JM0ytk9723Rr8h8FAJKjRnaIs7coYye5c4z3/xrVnwtJ86b9vSwaIogP0wV9wlqe
O1NeLenzOIL1kkCNY8RK7SpvB04O0kG8v3Lrgi0XMmkxgXBulxQOtHE9np8f+76u
9m1RFnvxNCM8rB8J6xa8XSplV1q5p7fGplpKu/jhU9nvtpoSY6esMI2QtOjKyxHE
oMbkflJ8w4UapDZjTOkEVA==
`protect END_PROTECTED
