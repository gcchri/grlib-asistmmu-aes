`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3SG6GXk9r5wBscr08ZlILpiAbe4+IBrhlZGqXoj5sA4Qai8LDPNC4k0gS9OBZv6k
wsdEbOOLGhLE4DzvoP17ThvpufBKEYejD8LJ2d11ocHWuZ9mOcDOLeN45Z2RtHE5
THsaI+GZ1p1G+JLT6E1LcFIF0WhajM+4Ekrds1DUwZNvBX/HcX/Ux39Y2KFkjvrL
DgA5CgrzSZYFwR0Fjf8B1/hQAmRPxS2MgBOyZIyiM7H5MHi+38NB4KcD/+ml4N9N
v3TF6rPl0evBnBpjI1K9Pa+1e4QCHi8m3WwydlizgS6fE/VB6KRT30ugSUZ2Qqcv
UVpPQy4zjpAiY/9UZpeT7Ut8Gls4Za+iZZvpV6zc3FSeRC6O2/oLipAFNtHpYFtU
9g4wVohVV/tD8ot1qT9dWRdR0vqeSpGXME2qlXnMA6ukZiS9pKlPo7KASHXHvodX
MYfHM43obeGDWqFrc6HDIXF01Vhjjx5exI/ui00Ai9EbDVZmoUWInczXIUB5qPK2
0Is3TUh7RC7npOFk+J1YOn/9uLncfkFk/qK7l6pT2bYqxIkXuxFXGb4STndictf2
SOUGzv6JAN2rs5OjoI1CAav47i34VNp9URBG8ieb6m8BbDS2IBDygINdlFHS4rGv
SSLZMJY9qx64tpMg0hoe7PAwcoQndzj2UTmxz3E7OmmtKHhdvi5iqpXcpAxL2dAE
ctF78H7m5nXwSbyIJL02dwF679/PtCiIwxme+w6KhSXw1Q4KIkGKEz9MddwmKzSu
SgYMCDYU8BFjfOrGbpxt1w==
`protect END_PROTECTED
