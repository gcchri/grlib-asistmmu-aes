`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8s/ER/LLFYOjDv8a8K7dkPePE+dK7Gwm4RrKqi4w6yoMmidjwPrjm6QQqkHwIT4/
w3yvfZHD5nwZsYDA7+R9HUYRUiTNQP8yuC3gEd27Nmfw7aqOK3VhW5yuX1c0DxZX
4UF0YYE2FELtP225a0j3/gC1sXThUwOxcRKFOqzy6z80PaBW7in+rsTOloKCpVCe
AhFJl0cPIKBex2qaiGHdXje+USnNfzlFd4X2+uUNs5I1zu/GMBRxTtqnN/8rste6
PArmGuHMjzKLzXmE6vjVpN0tlnaOo7WcpDDOyP8lniCUHl8QBs503CeYHpGF49wp
nNiK9OUSAryrohgWjPgXa6utRpKeOVMp+sZHh3YES8ZonjfEUlPcVrgqwISKWtSF
tNQRdCnSmm0H7yuNQINCmQ==
`protect END_PROTECTED
