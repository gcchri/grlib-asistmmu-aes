`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e7LnP89ALKRYTtEsNOWu5YhU0eZIgYMxb3s1Ag4VFA0bJtAWRvQ9aknxnofLLEkS
bCNFlUkYbcXC9KwoXobbN5uu4FHIEIH29fwyuca1Abu8gIS8zEtttFBJj5BwRoN0
7HZJUPfP6gOXiaCkET0nqk43d+wD7AAy1RZelj0rc2ijeHIpCDyt/gvhAXzgvgEv
til51Zfe5gYLEPXI9N+6eO/6HyyC0J1ZBAR16qMxK6uUBq8aCZ+irbrBmjpMVzCS
+tErRXLMNQUUOEb3zaytoM7kDc2yv9STn6IXGswf0zuFX+iUuE025ik3O+GUumuA
zHrtv7hG4eT1g5+tRnYi4+Agx5ZI2qBG8BL61PBJmSmN54ukmmHmkVozjALgFKax
DBAZ387wEppFobjzbGkOenBIm+f56qMZNNktVcEtm+6YMNXnejEw0m1OZNffQMmt
D8y+uuFhnGJXqdVOBhFhHdWSm6qUiEHZbF0ayn6Di0SMj+oyy1hQghF/brNZpo/R
tHhiFMeU21Gj/oxCGrQo/0bocL7Kciyg9kYgG4JxFcwLlKYHTjbGSVOgK5B3HDFc
WK0EtSFIQMI8GWmGOXHDFLANLUPiGwBY+Di1SFTRPlUTb5dNiKuYhbGot4ScnVal
/p1J4yUd7QJUjZW6h++6mEvTlvd/ahFd5ZGpvJgOmQqB3JWFR3BvfwiOL2UQQrTu
/yKreCHedXGfJknfJNLYXww/7MNuyZNWpAmOocFPXJHlJGQeFy6eNfb4iXfFt/tR
D6ThPeF1FM76DiPnu6oYgECtb4EfxPTSPIygd8GRzZKjxR3gDI6n/CU7kYEOTWOp
UgbZgVpzkhMOuhQLrM8zc9kaCYuktwOqlpA0TB/U8Y7zn1fRTKAkV+3dUqQUiXa9
tvn6FEsi8ylbJ+1DK6S2fEBseSON51B1gt+grDO/dsc+qw/b22B1UmBNjfwA3ovb
A6TUbNSdpiETZ0BlvTUVghN0+KjA/FfALboIm67QPkZPxTHtKphf6gzMt29vl97S
JMFm0dDz1PFiHRrVLtCJRo9fe9TD87WflMW7viakFDdfRpiUwLLR3mFJZcbY1X+n
TpfegcRGhlfb8kJBOVB4L36o8zcfNoHht5VrdbUc3we2B2Tif8l7z90rGKUngsbZ
Il92CF7ya5gNKsvKg1MaRN4rPlB33/WgRirW2/7NhRpeZVLxv1KzonMXXXJxEHa4
o8ulqQF7bk3sYYLs1fUSGO2LH2lxz8txd1IEbBN6P2aHP2hAGm+1P17DHNu40wDg
Uo1edQjZkDPsDMgEGmN33CDaDbl+eKE6Da8Ay9dMbYVf9/YsByEkaQ+DnzJIObr1
RM1G3MH/mhkkoHJ40bu+XWuAzN+lpBPlza3z3eCwnddnyuvZIC8iinvmSfOpv3pi
mApkEvBXsg+nTBlUHXXS1snieM+SNkY5C82eDa4pKjxYcbRiW21uIjqkUu7K5iWG
4RWS61vUpcsh8ruvFv/YwRSx7kTn/+sPPKnQei9ftd9o6wCzEDgz5nvqXrpmLNkp
ZdC7f6L78bNdhfapsAWXxKxTjkdOWKzFRQY4M1pWIRHy9SQWskT6zqmOj2qvBA9g
PcDROnby8Qo3S/7GQ446yezAzIdajVs7n21Z8XJrOp4pwH+O/lnoEVqU4VfNb4Xm
oSLX1HmuWfTdMC7CINDbaPWMSTOShBqaNWo2mjjzA7WqZFRs0ckTHlesZOpQKbkf
DBvwctNCZ8oFQAyqBoZ4fUrL7sIOgfJVnTTgbxrc/0Lz/b3ET6ANuZz3zgntjTdA
VuVAb3mCeBQtv2y5T1xK6Jb6ANiQyCZOTxanpt3RvTmrAwiY7/MYi5dCCiTf7aw2
oTBMzruTyvS/mTJ29PMKwjylN4DbRkaXmIuRp2sGfe8nLTe0gSCoz5Odap7f0FSc
iik2HePa9HRdj/RDo95ZaptVEQJxbEFKQSrg4eLrdHlXyJPNU0re3l1jaKwz2IrR
t7N3RFbQtuzkVtZhBU0W29T1zZq6GMNoLk1XQeYQS+YBnAKLHhh5cxgOXCs09tXP
FCCkGugxaJbgS53vH9IkkuSGsXwJdIs8JbeRZzz1naXRc9llTntGef1v+XqL82iY
6GwBqinvBuGgDLkCT1uUsCuhRGDm0B9bdcZdOmZsVVoHzRPw3vohSLMh9ns0Eskv
hQG2PywZCw5MRktxoPzVuifG1BBdUJ4PYvk4wKShOzCch5Cxo/HL4fz14kLKX0M0
RTfwvRuJ+8nXUx3NZxQTstvL/jMunxlgw0JRGhVAMcfUYjJh3KZAzKHZmDvSvztv
im0NYi+XQyImB+3aQ+i1b4NSO4Ubezn1nimyrD2ERYgn9QSAqG+8Vb1lgsdaVfMG
B9XmMj24XshqEtcRj//35VLdd8Nkz4YZdoTAV+XUgWwbUGOfAQCCAYq289eAX4Hz
GgXVjsKR1+TusfJeYf2cZdghiGeYnOKhFKMzAwJuazk3GAXkP2x8oLQQX1/fs+o2
fJcNM4ebqs6ufIN3fdbQJlTcbPIeHx/r2mQJcAw5ik+epfIuzxgBQUxJLuNNULVp
99DNh1aiGXRNJK4V1bHQOG35WeypsTF9DY5SBgsLBuWWJ5dCfRJJliHyUNqBdMcw
OnGrd92XED6x3NcmD1REVnOxJEgMK1FMQdGYCDMXJzsLFgi+M3rUbnEmV96OS/pN
6d6bCCiR5+6J+9waw/+eW0E5fuA68h8CHU8a27ccAM++U8Z3HtPZPFsvWtgcHa6e
44ZAlTJjfz5zeHJrBRtCgPR1Ree6HIpueVDAOL4speDjDcgI3WfTb1nVKRxzuyQb
kHVQX4trpYP1tdTmU7ujF3IgkLOk5pKn+5ZALhffafoKCPdvsq2HN9vOLtAUddc3
omVhuO1ua6z19V8VklxUb9g0iRlNwLdDOZZ/wG5UzLs37CGP/qwULMH8ya88hh56
HMvlz0HTWwhpLj1hs3Kez0CH6THQye43a4JC9ZoV2w3GeBwY8hKFFc8e9UjyZAlz
VE+tZxrlMvS4R3wl4gFeXUPLYFDN5mBhC+rj5xdwy3vSc3mx4RBO1hKpkCQj3CP3
IsQox1mpqoHL6sHmz2L3XzccsVzcluVmeBESmQdVDvQzxZ2qHn5oYSiJwXNdn5+p
nKckPdJgfJmu8BZCtBSA+c4yKiUeRfre1M5I90e5chIDzj78jc/NuYDnfyiym6z7
FK8x2x09Z0KLYDs1WWPF6HOxL70KyhQzy8ufzdHDFsRzj3334cZaUqh7JaN7eHAm
u1paJU9AmKwNAChSxGiJHlbldXnPKQP+tDHfAQ9NV13h5j/7+TQRHgn3tkGw5htY
/wRy+vM63KmrGcmb7p677wWHPEpypbPe5sjHcfuM5HatS3BFx2QnbFUf4Vm8u0S8
PeAhbe6cMVCp9leOQZ9BliUizwQGBhnoa2N36xtzeMW5hv+iPxGBydkDGDnJonI9
vKEGSu2uw8hHa2H84TjvDvEU67xulOU62EtJ1ZcuRrk9MjHHHFcHxDokvLN5fTnq
xt/RzXa1BdGELdWAS5HPEaBcQuA6V13hs28iV+qB0l/cpHYVaOuYv8sqQi/Kdb5C
pFXpdvFN3Nxzd8L2IwY91yFbehzQtVRaTnc2rQlLhqL9eENeK/r5gXD5kBn80ekf
z/W7j4RzjTBGqilmNmb/cz5xpk9KsQupqko9m7JCjlTVw00FfhAc/XF2x85GEHPP
uyjibXXYisBd9JP4S5iVX59UH+hk0PbIT+qEHIaOjLd2OYkVGfLSMwfwjCw26vS9
/zsNi1I0pgkHLolSRRKSmR8zrxBGXfmk+kLfi0k1F1BErUTzRKlhe1zecJYE1zG8
deHW731ETxk9lCggg87WoPnqKSZltcUKa1s+0yg21r2cIvamJC+klKswVgy9jsK2
t/Kel/tU2a/BRdpiQbeY+/ThHz06bT+5v2IDDxXgslc43uoDlXXTLjfv/xQCq+YX
LcpVZDzedby0NSJXYkDMekQat1OUUgetlLCX1pSiQV/3EXNpqeDSr7ZU5QQWhuX6
PDzYBXx3cuqFy3z2nGLIqfFoQVPoksUOYK1PcS8GQgEPVnqyKEqeOdVJxmNw1JVH
iIXQOadEH+d7iQWq0N6ZRKpPV/ty2wY1LohVSHDmlWrMUKJtSV2sGI7PRS9t0oHo
MXekCqmPoNOlFXsOu9XvvhHJprAKc/yjwz/pDSzudIZm1PCxxnXEE6nRrLIlY3WX
o4Tup8lsJ/F/TFpVIXaO9ucsUd3mt54wtV2I7ozpP8++fnRiWSugbJ1aD/TqChM2
qyXo5RwXGzQTBzcJszELRihQkDp5wC/lJFTnSeBG8by3mdkcaVACV9dGfyJoIXB4
JijtO9tsMPCfg9okE47FKHVK6KW2xKAWPPhzpfW08sSc/RVj0XMd6HpuG14BGMPT
7loueH8tb+//MyjBP7rrQu91jEc1uhLjsICZ9LkBAfMthF2bLwQfkfjndciEASXP
NnlMcOWPGxHmXvjz/1DEhEKu5GhLcS/Ixs21XIV45F0YxLBLYB1kz+IfyJso1Stp
tR9J+/eLbtsgsADdojFCTMk87jm5XPN8QuXD34/zp9fjnOJyheSHCH/bNWjEs9FT
OWglMZWn62OU/5p10/xqUO4tg0TZdv60VkVvwtjx91vy7sizAE4uy7DhzvjCGLYK
w157hTxOEJOitjVRqIzeJaXGA6uUCjX3+Zn+i2TB+cX0aNtzRzWCaIndv2v6FZlr
APOPgq4WVqqx/Uq8KUL21GJFusz3HKbUAzhVjlM0S9wzdsed94vj87t6QbqhqBoz
5QOw6+NWNFnbRKgIVe3uTh/759wwwgC1ucDD83yYdvAwjQmCF2w1Hlm4+1U2jm8Q
mREPunkBZsbteARIkvZiys/BiHAsf0m/g4Kb2lmXQmRns8S7uHu5MaEzbYFF932+
kHD0dF9N917BQP418XjcTKLnXGtbu90FR15+PBoNnZpY5z+qLdeK4s9itq9nF83R
zKJu6eTGDwvUgBwXKKkxlYXJOXy0yPTmWJYQgkYVDGjsSUFYau7/Ih//up7D7dMN
x3/jgA2vq34Y0ySM46ZPPQI/4YDX9dkyOfTLxkUCOkHmixyvWxRTDIvFyM4zC4fz
7WrKJyo1Q+7TR/dtx3B/K3nDahU6jU54HuzOKWYHL1rMBoR1qN4rgeDMwCt+nfXA
vHZjY4UEfetGr28DgO9eET4hsnZ+nfg6W6dfqdutNV++FHkt5O8A3I+nT9vX8AOO
eahR2dTeSJ64A/DoDsP+VaOTreKVnxgfCifkryEoaH8O963DnIx/za3JSgjPYGRg
+Fp3GPg5fM7IugwrGYnFaJqOR1aVSmykbMrvFlRyCSvY080EbmHsuKpdiUTMC0la
mz3SD/jZPwE+Z1D2MZTosoqgpwRSLOt5qKfoxJBeAWau58TZMLlqGonZL7lHsoUy
Ef16/3cNbl6UsiVMhwPp8ehoabhAOnWYi/Z1gb9ChXYesgxJSWJb13CVieV99T9f
65rs7LfnBvrmy5h9HlrAC84/N6N4CgY3IJdbFR6t1v5qXv95V3Zx9Xvcm+/Ebog0
L+F82QbYm+oxsmHbHp/W162+NqtA9RO/TckdbqS+1QVaO2AqC6kHzJa0NyHtS3gW
X9kdPc1oC6cHxtxDPBfz08Ie54z3tqJ3vkS0qyv2y3cGhX/rzzQpkRrCtb9YEI9g
eyMDbsICqDOgpb/rrgmzDAKIIAF+JB4zQZ95/ogXqUPYDNEbaip2qbyy9kur0/1W
VIL2pjbg5cQuICRqbLaT3WMRZQhdHT4pRkr4T+TgJz5HrDs/B6b69OdH3oohSH+1
sz9hvdRpNqm8nkTcdJi1cZbls8MVRCT0u06ke6Hczi1qAIOCWdaGMSmsUl5wPSKb
UTs9uikadIhWQ3QAmuDD/e2FWrb9rS6SEUQokrJojyN6fKwuL6ZAKBQXa5Y48GBQ
PF1GrPjDKmsmh56rxCC5mAoQrT/+jpebW9k6CWrY8sZ00tOd7sumuPn+ZElWp7CN
MiDBeN/pONopPoiUHKB0Uj3ajO86pxhzHsnJQZvSPRW3RQWjz+zIoU/0RLfVWrC+
74DmiTlOdT+I61FP+xiR3iaVdWfIEUbWvqdESB+OeovsKEhm0dOAmfgNP83XE62B
wm+SO3nPfmXs73KrYGWdJEZuWhHAvjx6uqOqqyMYZjLa+kGHS1r8boyAkmAKBKb2
YaC54hnHQn45dxdwGRZfJwjLDMXY9y1HZDlB0cKfMGSMP8MeTOLTtwMHe0BqKJZa
oDLRLqMq6LJpO60IyHf3pxBZ2FVtM0uQAgTh08L41HNDs/SSXfTbqjInVgyCO9YC
53ss9qQm29vaLaISvu8cztUkCq6SPPg2FG7xjXOiI+0rS52VnMgTxZyIF6KEfmeB
Spr2AjCMhxESOOS5zr0rSnqqrBrgEWbVLrG0wpSxf4xTsY34QPrHlHlbddo+VjOv
vHjr/LnQ9srz5APnw2xcivtx3xZ47MJsaqnu819iPfJP4jRF/++RFznFCYMmqrPv
NC5tZucL8IsdG1YSANdFmGKO+G2HYAXHWmbPr6hRPcPqk8WEDimmxOxfr/xql1ts
CM65o9I/hQqvQ7M80gLHkbIULB80kU11EgopMM01/t7AhsTYqF69GS/65sTglTzH
4tEPslxtXtyTRASZtwx30GMVyazzIuJo+5zOAH9vLJhPg/sz2MZ4dmH0cLIQAs3y
ib2kLP1Ik8DtdJgzxNVG7z9k0htXVqrAxGaHisQYOr7dt1oLOorzLveWAS3r1/xo
SjNJi0Qg6OD8t3YNGS/ovHeIZfnE4mJ1jOIMqvZJHtzsZMHLZkUvVEeBi6Xr1axv
9XdsffNfkaqNIzIVWXEk8akJlCG8nFXsGxzLisAqyn0G7RG+Mf0d4b2jhefOsoCH
iRpOCCi5eZUEWGzbs60+OS6IKeOt6G0t8kvXeym94f7NGXcFa93cOh3j1AYCPg7N
I9Rxfe2EW0WUEFwz+Bq+l4NX6P4qhHku9OYPl71ILeoeZe4w6NqbdiIUtO3pEDi/
65aUNJouhS5X53CfBIJsmHpgOgzwFFn1LOfhyrhmK+Q78q5JJgylCBgvBAzk80Qb
oAnwH/4M7ubmmwL8OzgfgZ3Y3y7CyjFhAw/m4XMQHhBwabAjQzuQrWCQV8VK2eN1
tsqPvDBuEu4Pf+L0KORF6susuP+oJGmd/V+mh+QXTA6mMHOFtMib+bIaxnjBtL/f
+uf1h+iFJ+guh+mmF2k3XvWSGRZiI5u4RL3KM11MW6SvobR7o/lsjCwnrqlmIwaO
st/gyq24dnbRCTa+o7Qcgh8rWhHqMEeV7P+I6WCLuCCJEOKnQetHHlQJaluA12wx
DPEtNu4T+wW0H6N+BL0UPiVEZuVryIqkdpfjJ4ezE0XzfIVSHv4x6IZJpejd4Fm3
85oItYHHKDyjCiydh/Ifer83sdLfIGnq6iuE3rbTrZU46SlHE+cOKNBT6mveI9UU
oStpULmrOvcvwoMYpLR5hHC1JfXECx2U9o6FcJcmHlR0ZeI0ErXwFv4TjnQH+RZb
aOWkuccjfFjHWJGBuiMpgKMXJCiXBS3yxnaBiRdlD2hlBh8hPhsr4CJdD93RVit7
gOxPsaMpRKX7FSomrJK7hKGah/SOAwFY8/0b7fWO1eYLWYS+XiE460xB8/iAiyau
1acr6Wm918XvNAYuTZar+S1HXykDYrvDbTDW9PircNrpp9AweOvd2GxdmHIsZtEP
L5fpUtD+IwMQmtnopwLHq7mGqYMBJOIAlJ3/4BE/a+Lm3cn/f1Y11hPgnaaADYYR
+vmKhVADjNAy1uSWapGsBCHcbIIRTL7OnDQu3R/Lkk78Pe+2e0ZC587PhBlFGfGO
HNRXaSzdSg05Yha4Sv03+EWNEEPcMD6bNdPkavEw3Y6vJgOCwUBPMyu6dJmasAy4
Vh4Tbx71pD1Z4mknHItOtJD4Z2qSe5hl9NHRAIRPVf1XTMFi0npUAPbNnMZXOreD
T703DP+taeFY1HMvVhA0ksePXt6LG4MBsPROj0BVYp9rtSH3eReKxlpd0agwZq6r
rHJ8ujpxKbSeznXiFE3KGmTqEzgzd5GS81DNpxZiU8D7BoCocbL7nSZlqk+CeX5Q
dxboz5mAcpBTzcebNUCEpNBK0I4jaa+1t07KLTdrm4KUo0VxVixoND+Y3uTldcj9
9DEZFRUF2iOnhdirAp5kqFJ0uajIOyJ6dvkJNPnWuzLrOW5P/aJ+9R6CNyLM4LX2
wgG9lm+zoNNS/l3nb1d/1ELIqypk8+Mg1+Od2n//wN96YBYcx17syfc3P7mZZ2MR
dTCM3wAY0j81zsAuaYw83zedFsv/0Bi0qk8R/+o0KgIQCHEPCITEgbzZism4PmZS
zCVJdfY3lpOj6v5gRcund9Bgw1NQ0SzL9AgltWNl4cq7iGo9UIsuz0nDjP2nGoDo
owIlfFFv7ACQmKfpLJVbhi43GMNUh7jHdjQNRosuc2+6qLhr74qBCns/O3/eJDC9
+NEnmBCCwh5fX0tAmm9fs4+w0U7ImHRoPmHUq+IMaP2NWzGHYrHREFuYUyP8KuY5
qB9kchIp2ivaZEzcN9AI31+iHYIrkNmQCnNgUYrsv41m0Tk3fm/Lozabaf+Ceego
EwJAo3Ec2cndD4Jq4eDliT/Eweql9JBVyB0LizIOPPv7WT2POnm6e//mrtXQXg12
Qf9DdY5jU+zQhwzQnGha4wnPREvIZam9pFA9T+N4vngtKND8FZACL5d3FNNhYCgU
SQCq0BW33PD6kv4QvH7xqg1WLNFNBu8yhHbWxXhOZh3wSOlxTsAeG8ednTE+A313
0NX46ldVhBf++ZSj5amXCMZtQRWf6238ubNSMvAkxdJLbdqAD1EduC2hS//MC/50
G9gNGejfoc9lebA6otjP2im+jov7u7jQc0vd2ouCmLLB2MN+XDACDVCu7UCTk0v0
tKEDgfLAKhATSPozXqp+gXlIk4d8tmAV8KCw4ouqjTIS5imjKVFd87tGPR6ynBwv
2fJBjabIPplU3c/+UeAzi5hpsgVwbV2AlJZCXROd8IDYg6IDjZwDAFukY8mKvH7q
+gnbMMeegPLJZmEGuxBJRdNqRz8JvvnnB97AAZSmx1G3jLvYA1GevTUO498vP6dT
RGykJBdRQPvqzI60C6wgW0zYA7RWuC6fXYbPBlSFs7kXmW+VaUgnj8YgLPjEFLz9
wqBw6T19fZAuPhgasoSGArWKv+3Inr6IGdJhn1Ay1RH5Xe6n8aGrnCW5IvtU9GuA
SOpSjtACOwuvNiU9QrtcQTVREVpAN/8Px+cc096hoa2WSVE45wfmaKZlt2hOeHny
DpjOcgQpAX7EfRKi705s/7VaSiCbCf85Ztpgb0Po3WEaGMwaaJnyfX13CqaONElA
tCYMXEI9aKCCX/CroANZ5VvUkFS+aaOMI8PNx5LdL5JsHUGf6E3zvYO2YEYymmim
MomdpLbZzJYvcDVGOs3CqPwqB35TO26UJIGn0JLkQxy4dJpQA2EYBFpY92OQsgOr
2t6g+8qozuEWXsQPon+yQKn3xI8v3tePA9vhH1kIUqz4V/h8lOHRbwXb9wmuQi8C
YaFt8wSJeMPh6sJgLTjrlk1rG+e9t4xWMn81ZSeX6L6vL4G0WzhOSO6vbpfB4GTO
ZU+s075CS8yNqfA/1C8/2tTv80Dy61v+QLSEYcR9jn8iuSeFdoKzUxr9pLzbc6Il
XAW38VU+NYuF979qqj53f1qjRwYtMGX55ahjng5BU6a7HtELBxBkxQZzX38KwbQG
+vlXRqdPCeITQ0FAyQQlYVmVl7nfHUIK7RXCJXS+gkGdiOBnwqTOQoHyKKsAfvLJ
Dc/jYnNQyamj3ExLXj8nzN7cpleUEVQnYtl1h7SMevyGwJw6b4EoBOEl3/mpOumr
jiJgIsPBlE/S2bb4OtwwSZLFDScNIWUQtKPzBbdCi5caKvcLtFW44p4PtnhiiYnM
pDuNYAMvWbrYmi41iGuaRSHuUNBXH4jFyuVixTUd3ubfn1HeDGF0mtvVBgnTXsJ0
JN71rwmg1UIN3f3TFpPbDOVMdU75vT9Ruow0SEP6qYcGig+2srw66xqEx+WoSypy
w2+IEygs1pxEtFssGdHXvklQ8osV3Qp8K+gZICakjFQNq4k+oUrLhKfg8NoHi0SG
/6yMACvmSmTE3fuMkhDxy+5jOLI02kiDbuG23bdskTYcoWC/YmTh+qLm8LI0Ioir
/twLX3nT/RazkrDuKyhggPcdID3Qb3rRN/XeDAqZrFVz5EbsytpTw0uY9TNH6aNl
4Kzit831HhXXWho5qPUG9jF9TC5oMp2cKwX1/BRLqHvwrXouVFatqW4/5sx+Dm0W
A3Rz+iCHO07JtLitzduhZrxZS+dd9vjqmafac0oNNMWxlC60eWsezbAvgAqRTd5Y
CI7l2ZLjSwR4omPX4mEbPNopVed8fEKAnxEY9ibMs3jqcfYhxQfJD/kTGXS0AjXL
2aYCN8PFuOkT+QiuaSoDEA2TZQVjbXpioSQhqO3s3F/e/D0F9IgRN5vOtPZY1c8y
/vAFqZvOppT/nJSWavRq2LCtOxCjj7viILhufwhF6FJmU3Og+XEQmf5QsMjpXo2j
inoI4LX4Nc1S7Ai6bp5cbgAK60dFI5iGoEua4JX3cctW7NCedHDkzyrDLrknR7jy
3D9/UmfHMmHc9B8b7oy5IGCrs1gRFrCFPPGk4GeEMSQs5UO9Im5EFiTKzt3YFLLZ
yuk07GJ/S3xYcTdt7ygKa6VLdV0H3eb5qtxvtvNqy7fWvTaf8CscK+DQ2jfV6hpe
wkfaqD7lh0TyTyWVRjVL9cf5B7n8fAbiVNpPdo1wHaGsoylKe2xNZv9cnnjru4cx
KFx4sjHt0q51UrA5JGVDLFCmzWIe79/r/5fZe4sDOhUN8cdld9aMPFdx1RLk3MBq
KXHPxlHbKADFHC02eCHTDxHeTk4oJn7GVX0/RQoiaahafpSOrGKTeAeLG+386iNT
1wrI8dPzYzAMnlvdrSMvw56VOXqNTqJziXr7q56WIsakTv3BAJ7Dh7O8ik7E1Th7
bgur4NLtGeI4bljgZrSXSj34oRWC9HDqGyuVOx86swSnj2dK/ZRMMzykaPU+RS/Q
uowhHjaoODy+YNQo8ZaL0VRuPXWBxU6vozzHIgiaDsDXsFj5odeItLPtebxt6KmJ
QXHqzuAM/SQggzQYP8JE6NJj8ozzgFoAeT0TbObOhXG7/bPJxG6v2RRbvAxmdFpQ
8xGLWc/YPYJ430COwOdEGb9gZ3R6KVq5aHjg0qg/kKLugF2/5x3S6wBn7e0fH5A2
7f/P/FPiwLJ89Fjkf9JSYfKAPf5vvoBqf+lRzVopsaBofI3VB5oz5WXahY/sXDaY
Gab9kP9pA232KqTs44qCdxcY69UalB223NKdbJzjCek9xZK8OXpT4PJusotV3LR1
7yDrKGcDWePrzO9UIMDjBHjOKE/RTnEXxSwJTJ2GMgR7o8yx+fowr+RYWq2xuTTj
UIq2HmhzsjCi20qRvSBFpnzxKtLb7lI8H+jqDmvGv6sjIc/ZwI4nVhfl92J6j9Fb
U4xPMD5GBxrnPACRimV4DPiaTVpVfew6t7KgGqWX1vdBRea6ObNLyRcN/lPpd59J
IHqGOrVXHrrcAjN6t1a0vHvnpojDIK3KG6G96ABlYP/01Mz0g5mQpURZZVzoE9ag
3YwkEU6xboxKAyaaWCQaDU/oARRi8V6hCBnqfNFUJ1T/z+uMs42oADdt6FQBr3ye
JuZxCsmKoXynnvLGnQOfHlwE8bGHZwYafjbic4QUMR67EEH7T4w9BaNCn9QyaCOW
+YeGqFXp4Po1pcg4oYnpoB73BNT7pNiD1kZGT46OG+vJUdHtQRhXi5QucBpB+hY+
ZahbQKs88AVvnDdyRI62LNqdmCp4ExeOZXvf7og9OfMQ2d8TaIg+NdLcbRLuFbNk
K2s8P2ivnNPO/em+GsFcoD8gWdr4DipW9+MCLb5nsamFFV2ao9OHTXpwrF9tuvjq
97nHdF9umQX/FkmxYXFR5ZawPLEZndsZCy4S4PCJp/PcCu0PXgRVBhYYyeWx8Xjm
QzSOWY+A5/YSnM1RYvRGt6xY35RKzBCAuw8fYeVPH6yizkd7PLF2Sq70zc2pl8cG
XDgya4dI2Fxeq96LCs74PHUlqwbY5Wtt9l0C7xYR2M1XLAMefX7tpeB9mqKEFk2s
7NoeKl8Z350AOeMHQIp07b9ArMVfHO44wzyyyNJRaHVRMMO4SpVpooH8U/d9YhlK
KXSkKV3IYO/MqKRlvBDdih8PkroiOtqy63fckR1JOgGTu2C41Wrm7e0xnG8gZAl5
Rv2n85KAHtRze5gR6PdSkyMviruEw0LFFP7AU1d05c8SqEgH+RGXJ9+WAz9QQ3Ip
/7uVkentsd4fc4EoEgntM2YWle6gC1uU3ry0V7yW4mSQfRfDNPDBQNnTmKv55y9v
B83nK4PCZNHgNxqk0eliXfVuwVjxIpzq9NyXaLyRgb4vNCwimRKsm65kmQaYQGHe
9ipp/Dli4lNLh1jecvuAQAIvRlzThNmE6xmz+DxGuld+F8igFZLhHV39Lu/k67ZN
T3/ftFCWhRML5rC2PcoVyZc48hC3qjRXRLYCy84gzVI/ji+nj+UN+p8dsAyOit0W
Gkow3FHrPYXAHMsaaSlF75jUz9EHevwgoknnpzudV26SVFl8kjlRsJ0uTJKQ6C+x
NcwRsnRviOR3whVS3f2di+zbBFqojHF/p+/J0jry8nyqTMl2G4oaZGz3ZjH5cst1
UtwTWc7QCkKHk0Ow0u/DURJm7isrHTfMMwHbF7sHB6MK4NsDNKKVeYhj0qCOh/vT
L+GVuTIzyR2cQojJlht4ioSLABYc675z/sN3uAlUD4zK9+A+oFp9vC51rCLSBr2O
OOgTjAph1N171nhVY6R902Xyl5ScFMVlmwkcpj7KXklbT5aTWFUUsm6HnoIc0y65
jV2RGNij04S/C3z6YLUgXod/rXXeGCPH5+gmrb4malr90f7sY7I2DFZrCG+xDxm+
EiDPF0DXEwgoo0IsJo6m7BDMxxISClq+HDzE8A1jne1D6dhlSuUhjcYFjz5SiXKi
0YqrugHP/75+9bL8JcTWRGvrYAbtKMEh/6GxaME9MYPcKjG6kAjDsycVG/dDZL9m
AIgpiq+RRTsp7MMXirHs+vtRgR1broHSdioYClo2y2qS+OeRNzgUf7aSXk1bemu+
eTtSCHWqrm1mPHE2q0pZrSQFteZI0BsAMKBLHZ0HJSAZ5+EE4JeoYecAYAcUwMms
ryqA0XoYW8wJOnJLP4nNCtbyyKQlUULvcTBcp6vMwB4OqXPlyDXeJyblNXgf9LQF
6fDZs5oQE95VoPnGsCr4sdqD6ZXFg0kZLEAVGOHEvT8e9l8YS/gFMvwi4YDKrx23
XeGvFotJPQms2YkpMkMMVaN81chLBVMehZToSC7t1SQAhKkChtQNFAydYypBvppF
Y4tRNADsl7BWfVS4jKfx7YswVjHNICmC3/yLWWD6P/6r1pVg+yfop5huOx0si0Em
i0W+1Iz0MekVsjTgyl4IAVN7vyIbYp1Rm9vIrocPF7VBdGZ7/0qobtFwbDx8AqbB
eyKN9UI1jK6R7oMMRZUp0uf9tlluTdzZUSmu0A2OYTZg3QTi19YvcXNSfNsmdGk/
9xnq6j/3ofe7UJSAcHARbX5hGMlLdy6jJFa3ywAkKEb2hmcVGQrz2AEDSouD/0/y
bzFvvy537oeLQdLrDZ1eTdUKAQuu8Wh3FUHtAkcZpTXMEVE07xWCmIp9iFBhOxhj
J1aJbvBjxB7S5DxvDRA7bbBSMbNWkEBvtParKKWz2XuVti3EUAioQT+LmZlVZQ7x
Oc4qUWnPPsx1F7Yj8QkVEFAz+NkURDeVUY1imEtxo8foEs4IMjS9fdPtN6iZQYjO
ysvR3Q1impdsF1dMPpRjN1nHABMkEd+ro0CbpQsVkkQ+mU8wM6yjUsrdixSNU4Yy
iPdaaA0xBYeKb70342yzusmtBSs02msnTD/YK/gUs4SqT+i1NgWXMleyAMPiCZqK
BHHEkXRgql+AGTiyL827lKz2biTiljbn+4etC63g88rEhaujll2DJKYk9erWMiBF
dAOgicgY34LsiAWIY8Cg4fFgcSm9pTKhuqU1i0TEXVy3Lzsn8iIqbQHqvulKks9x
HkAakwSUuTqIXIJFQwztwJj2a3QjTl02SYBNJjyx32QlosYc8+rU0ZcJKSKdaCTW
B25XhdUPjDeJgGvVi106TQxaossz7oOO6kQmhFdnRC6/Vib9zD5Q+xrbq62BzbRR
+7CpfmN7KIsLanRPi8Mdh3S5Wzw8PG9nR4kMzSOFrBhmdNYHc0XZL622wFJAhb4Y
3njPi8FAKziDn6FVFmZVtY9XPCUFZfK9H/a7GMqpDbVy0h84UHxXhzIvW30LwwgD
8WIkC01J82BPOFoY5pl/0Veb+KZd7SmJ7eItRyrIMHA/dBkRYTwPnvxRzDlRTzIY
VcmCLt8Md6oQ6kGBWCwrZ7z6/GsYNcp+qej2VS7xIywrZY0uqxBph42vfIephKB2
qFBUT2HBpRvAyLDtds3NwTDTevKymxxEzQad0evB7PIJpv79LlD3knn2neTWQmy+
NxBZzzJgN/7VdmSijwHhTzTTuOq2XGr3wuVYltNwroc38oNA2ckDQhXD9dXPw2/F
e0pEmTVvIR5fHfIIWMNaJdYmIKDR/qqsJXmhEUefWs/64qSEBI7oysoUib9Mliwd
TXn52hoRsOzwObriBEtR5oohL0KrFHAPR7gFV7onf7EtnQvNDWSUf7T1PDSEFp/F
J3FQeS5h0TAx/2diG214J0CUsRHed1xj+C5dgOfvPgJkhuwC+tdVOg2N92V+8y0q
nfv5oVpIh7UNiIkC7lbtnBo4RMQbyrYAKhC/yav/O5iHNxAOsnI8trBilHR9zyuD
PzVDvqDPFkr9AB0dqzMEKPMj5byUwaSiUBVmQIAcFDJKnVz9yvm8fAekcvRrpNhJ
/FF+d4cC7PZYNZ8LYy+31zYkgc/zu5hu8te+/IT+EoPJrjUslEN485Svq2eSwg0A
jgeWJZVJtOSIprpMHW289RdLGzFZlXAhuxKVQBd3A9NATQThFDzBInYUN96mm+dL
sjfhRvoBRFsv0/KXZ3lGUoTgXmRp+jWaR5ui9WFqh4cPmQG8h1TMWui2eWDbW5W/
LBWVrS3Xqis6PcH/9Yb5WxuLtxDwwX+6otDyg8zYjCJOSfQx+3aIKCBzJiN6/4Pa
cP/27ZFwq0dajQzjxY2qKDfdsOl2CSMl5vzP9XrCAQeNzCAQl7Y9F03JanB8K9qo
6lf6XUWQ0pJHW9UNZLao+/xlL2XUSOO3eRCDGtXxRAZssbn0c0RMpoIJ8Fc0Tj+k
BFzPBpe5Zar7NHdMkuB48pZpBmvTHJwf+BsnHhQuQZRHnVMIRUuxUqGnreGR67Nl
PWeTqOQc4TnbN8aWuiXH6EyIMUxDnVVeWNkM+Q8KXNh95ZR5qTUGdUU5BWr4HoUr
9cXKlwjWECVgupskcZceYyZfA7Kz6XDhnRGpxYTdXMaa3WTIgTX9XSP683iOhYzi
vfbt3Xh/VVKmj6luQOBowO85nN5PKhOIoIbdH2v5LjTo84qDmwQmV55dWWx5WjtC
4Q2FAK572TiXbx3hl0qsnQmxjMUE9rWCYzkmZhAUZka+iGedaOrESfqHDDF3tPUH
AGfjGwuWg0RdJ+OFpEPlhjHIaSvnQvd8dcZb+NRssSZSf6rBmxr7SvSiq0XW0tVw
AJoYP9UQ5wZvfVuLTypfqN3uAw0ET/5VTFEVvBOBg1dY7lL17O73sAMMSAaqYX06
vSBI1v7dle/yptE4lt2aiZU/jj1jO9ys22n6JFf0U55KraTI+ylgBo15CWHq4FqX
wsmz2BxglurVDwMuU2ZlXqCSs2a0Kaj4jtzjhbpkUuF9rNZjk/4+VKZVCvun4/Lw
1fXVbhaBGOEcZWj7XBxuJ1zH5U93foJiXX1zi6sC2O49HDB7xg8DSeUXNhVeobEe
zhFWqOiADQYWQGBhVZexF804/NMlBDrX2ZaK8ZbRstQB9VU/z4nCSQpUv5GDFGvK
lydp73VBlwXBa3LqIFyLgKOfTdu+RTDGm7FFWOR2q06rcyMWcka0nZ8b85cssQ0Y
9o7taP/qIyI+u1mG1ULfKaRi3+YbkKSmSuUqPlCjE0JqQ8rB1y3WhFoxksaIpMUZ
Egw8J/SzJIr6sIdiWdwrvw985dxtlcrhQfTAKvcBV/awhoVSldC1jSfDKdbqt6Fi
EagxpMm9ohM1qiXwmAuTjcCbH7/5ZZa0v9NcSjSXNpUL7PhfV9sBBfur3MpxVLaf
zg+duYUFtYbLPba1s+qw46PkZFnKWK3txbkdIYVZFSrs59WqJg1emY4Y2A71l68e
2pl7GwZNk8KvZElbrc1PfNghMTHgx14DdM/QTpJp32zQ+gahAk2VC9fTitpy6qYt
4GlVDeOvxZnh1XR4DgEgISFlBdOSw0wWvofiQlaiUYcxAmqnoURjcoLxBlMhlMMI
IF0qUykkgf2YnkgGJRj3NMx65/NwtPqi+h+K7yMnN7p9Bkj2oMmMg056iuiZTF/E
cwLYlXFeZ04DrUpq7JlPQecQm2XT8Rg+O6FPzz4AN3DXsyZbFHhUlizssALxY0q6
vlBdnKD26FV2R+ub2gPuqna0mo560gkgkMrC9n6eY/m+fzwgzOtw8zXWo80fpNuv
qoI6VIc/JP8VelMibjvloIzK/8L1JBeIwLiEJSlq4Fp7Dm1I8AaIxB5Tvvf4fgQI
Gg5S+Biv9KRqmDgioqzfU+IhLRg+C5hY3Rbv5FbergnL73+Y3LBHnQm5z+zPQnWN
l/lNI0RnmShNIj+7Sxs/loXzgvGpO4QUoa+xBuUvBdc+u5n7uUqjQSHBEsNmBpjW
SbMCoBEIhabWvUQr9UlRPu8rj7BUE6cpYGJ1qxgQFJj53OgfS0l0MmAcILe6n63t
Qq49g0YJrziLKwAl0CXuOCviY+UdGVTUscoBqfLn2sjCkgxdbToyBqxJMJGfffes
YAyaQr/jKjMzdotWkivJe/rHkVp5xRZFcXt4NayD1OFjmeymGu0MIxhtvjuCzswR
o10c5BdKdZM4NdjWmM4+PtU2DU2KjzVMZ82J5IFcmvXdvSmmQeVv+nQyQ8vzKYVB
qYIG9+EXmpxKHnlRD4fDlq1LqsJlEUk5GzKzBlLm4SZae6nVoHN12JencDZvt3qr
92r3JZ1VbDSTs7m5maWhgP5gsn/Qu/4uNQBa3MLbAHeMxGI8yacJTZWu+WTAOtoZ
tiAtijn8hxL40jdqsx1qyt7/+JmC2hWfv9tJEJeXGQx/B2jJbVD51yL+LXffDHXw
JricLyvjpghXQNARbieksvI0dtOJ3fCU1yXinrTSpqFhb0V5Ns/X2OD/hEApVniv
HbLlLl+LB0ovxm+lbxUeRWNH+T0KAU3iJvzL7vsfJ9Xms9eWs9nSRR2WWrObj8i/
aKBwxj/WJTNiptuAfTezXxQnucjxeX1+9e8vcBHNzbSme2l69D2PhvY/szDvo5Tn
GhytVQxBwuPPjbHbyE+Tv7mjJrmNBBl2Cr4V1ljQtEacAECODX8ffkis/514SFVB
5gdJ5coY2wv6J+zqsu7PI62nLQ52YYPW53LtQfcbOodo23PRc5epbtqWes6dv/vV
2umCP6hgiGJ0x4TldWLy84/oZqkY2rEOs/1xTNQkxpX1h+R2XKL05xS5YVpM2KYt
H/M6+BzYjp08IGKx6gFWoj3xWxOd9248U4JkWiXMkFtsDvfETmSv5Ss7iiw26JLV
dpse4uMXQ0gVRRyy+dwbkZI3IoN8RN5DFvNCKgDwBQVv3MCcPEuIJh4Hz+THhKDs
Z/4h9/n7FVvKtJkI69R1t7uOoFHxf75K7vIim1vKVrtuUoIOcZ/Z9eP0S8JckJDx
okXLnkm622h7dh/G0h9G3jyI5XBgA6eUHDUIUqekvgG2ChBGoFX1ZmGYVPZGAP1z
`protect END_PROTECTED
