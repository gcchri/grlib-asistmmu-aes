`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
orXuZxphDuXn18hqaMrKqjgIuuPfv41zlnlYa/qqWxlu8k5P+7bTRK1yUCLIdywf
SBoshqIPduuw7NxEMaTi2s+RFr5Di0aeuMavX3iGX3mGXOohLD6mcLswwBGy0huM
Ufg7yWSiNOTX4X/ZzE04CBpdUgpeimNz00QNTZGO5tcsc9oPHXr7pJ6LMqCGU4NH
HU72PJlCtsjFNLiXBekkGQEk/AKsoq+AC3fd75cvIJMYX6ApDT3F+vZKPvj3uvgc
fVzDYiZETHheU6l4L022rXje9JhPbjJ434cfo4iCiEGKpGLUmGdJ3GxFWWg8Nhpc
YhgJtPPzPoCnDAL9D0MarvU3uWbKLnN7GIMYxcOeaMALdWVNGOeLdRA/+Klbw6Pc
5Pl3yIoH7IKHyHCKR2JRkRp86V0/9j03m9TaMOWMotNpFS2NDV45G1MQFuBBRZGg
5NzT0Pwt0VZj9ejXsVOpwXC3L6XSow8YSltW0kVmfKBBpnSp2uBgSXpJHq0ArC21
sZ2dX/7d/lCZsADf2GXA+bDcw5HCrHWmdi3VjC+jypiQAN+JcGHK4jStillHn1Sg
KGEHnmzqrz40l3oFYg9IGrmcNp+TTsyHr2VgnQoSuM+/bC8tejUdvPc6st5lIcIf
mPVKiT1siTuJp8g9zG4gi7mBB4m9Z2J5Oiztro1s/ZXelbAnnolORgtFWCpqOX+F
vj3VeGf8wylbld4F3RM1Vk6GsV4Q+nioNEiQ7RXbk+k=
`protect END_PROTECTED
