`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MWhpJrTm0FNLGoNwyiqonte2Qvk49RhBd1pwaDTw283C371Nb0cb7wMoUAzyq13y
eVFxIuMamySGDnFkkn0FFOClgAaEh9HLJ9/y5ewzydWSk+6gCj9Xab/As8jC20MA
sJPFM6bTAPhxQ7P0UDck//mP86qMso/HzySTPA7mujPoJ+uL+gIMUTWoXg53vPOH
0vQF0AwZBuxKUiU+8EVagtLQ/CXWXah2g76DAXLFPB0TNMaBRUh2SGAEond8djPn
kOlrBtw5TNh2TO+TmnD43FYwM4cnbDwX4DJ9JdPqt+gWwvUQFuqoxkGjrK3F77IS
vu4fMSvMpdXtd82AmP/DNTOSSS+pw+bpg+F7vJ+cY72bOaf8tVl0scXyFPSev63a
lKQjfyYfX/YuhzmQWyyRmkdbdCa7uSkdZ7STmuhoRIwiN5qYuT2NiAB7TZ/WYLmy
YnQ2xEQ4XGVAlweK1c2CNPckqTlnBcyDgvWj65MKnIg12MmYftH9yH57lHMAg3K/
Rl5QChifN2FAF2UhXGk/fIY7Ix2NberKTjrJ16DVzVvYstK7I1BV9a8fpZSm1UN6
+FMVfKu/Qwzjqr6P4EJoXTeINM+GSi56Mtyy2wamDJyp4F0a5EaoTy84oZ55q6+X
cDehJsPpb9oLifRLWoPLvMEbVzut0fvnOSqIUOa4FSEb0QiU7INdYloGMyNext9N
CxNVaCtPHIL78TvC4XZv/nzIRl3P+DlPvRwxYyMZDkGiDGLln21kkAgLCju1B+L5
PBZgCPLjo+3RUHiMaUUcn0NUPIEcibGxsmzTtGwxe0CI0/32/EfoJJGWxwrfhRsX
AEKPfEowGOQPK9RmZEAOlgDmN3nT008ejOypws8EzvwyYxeMAGafALjzD6Q/bD1I
jpFUmvoYsP5nA38rS6qv4CAcitU7pXuiu5kuTN5EHGUNdroSK7t8PeTXG7QThwCf
jO3+9XsLoMiloS9YbrSuR6JdzrTPqinnIyFnVxcrc34=
`protect END_PROTECTED
