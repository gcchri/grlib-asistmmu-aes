`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A+PErLH1T7UcUO0G5RWFymOps9RkZouazxCw62r8znF/Kpn57FdcmqaXIRMXhmBU
vIBMuohlof71uxwQ9eGv5A+rd+dYOWsqSVTCUpDWeYOs/aP3wTicyTYNCN1giD4l
204SWkrvaBhByuTL++zwSk8guNZ6SMgp6m7BOVOB0WZnu61NoxVuqtorKKZ7EXq3
ueOM7JNkLsAey3ELLH2VITEWOBgqnfbzYSep2RGXRWtU7koDT8CoCCtnFOA5G/Tb
hoE+ztBylv4/FbRsFfT4IYFyXkpTAboixExykrGVPrE=
`protect END_PROTECTED
