`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vPa3Ly/4/l9VFKfo7zJF+NPFJVqydIhjAa7TNGbJUSMZPJrnLjGr8GVXVfMJS/VV
BzkUeXcdoQS21+30ub3xZK1qEVYrxWJofvsDXxRmo3mLTFhF3hZdJEIcIudmjBHY
n99oEyr1um910FQD88ZhIpP2b49fYSDpl4EralBJsKLmVghieKal0RYnL7psNVpx
BrvUtkHbwgmNe1qbEr9q6yVKPKmj0UYx4ub4KiWFNtJtCHp4xCPNCznRFDOhadko
wJ5aGNxS4MT5QFOBOOhA/uurnoUvYz2lhAMtJlGlnl6HLuotdt5CfjqwTqDH8y+5
3d/wEX85WJyFNJwSD/rye5aQi0McHcVI084lILVZ0GEKyAl0Wm6d6Bl55ZDcitNT
k6hGX6zEtkMGjGMGpkw9z9+Sf80kWPwNZEIAz8gYVuyfweMLRcb9o8vdkmFP4lnh
SJFY/+8yepFVoyLytACJpZZ/7gvBslwRrVPMf2jTcOlrTnpoOZgdjDmQU5U4rjAp
l/I/6BmUycjT6IQc32a/l5ALwZPT1DqZ6duhoB7A4qpAhrCDSelTJ4sxB8pEjXsd
3unHx31/nNTv8OW/BVw9WyN7nzEDLxc+Ef1eKMATY8IxEmExkUkTzLuTFypMgXwT
7cuQd3hFii6N4ZLlGI8fNkqgbGyV66Wj92UFKtaZ/ebQ4aS0sG4LS4R+GqAFqVKl
XZMfpMzLAlfP5kv7YmJbC9uhGYUt6X47178WBPgxMUsnXFogDA50IMSWP/AgWlaD
`protect END_PROTECTED
