`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zqfDGvj6i/kh1q1nC+/HWPmvfAd43XGSNhpq+gDSW5KwnQGh6i3MvgqosbFhN7sg
byf7ZxDeRiltERd3jZvOeHkJH4kLq9b6irOZ0JLrD5tA4De9WeZ08eulchfg2YO4
sNm3LJ9JixaRcSiNOmEeYsBGhPCJ1hLk9zE0bw0xee+KC/KXI7zQBrFZd9LEQ8qj
OtSeVkcq/tn4uhnBkjD10lrvfWMX9ILJd5g5H5XKj4fZGWD/gl2KUZTRpjbrdeGa
HmTAV8MJ8kGqAImaomntxgwo7OZ8L87jdjPxjmdy0U+QxkWshAh3UjTzscJ0aH3y
WubrqYOnEJX/HDHbTei8LNlmNXlmyhFucd8ixYGEz8sRfcgq0jOYBC1Fr7k3+dkq
hyaa31PdeHfQOUe4iE0Fbg==
`protect END_PROTECTED
