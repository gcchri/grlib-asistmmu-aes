`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pPWbXFgPsSNFeQao/2lkFvCiOa6weBm7tdItBRSvQO84jgVakXvzqQBG/pG3swMQ
qL7DU/2GQnucPU1JznBCcpkoa0ZdvvOK85FdGRlxzIuOia5DeeO2DM641K9KJycC
kxJ1JeTqrsefvbBdTxpgiJedzR4xiJDBLF4aYj7xmqo4uwwYq0XPkkFwcsBVnHwa
Fhy5cYn4z/PVcdUeCxM2bOfLyVlVH7oZ+8cCyQ3eZF8UktxuQlk5ae3WBm4YtXOg
yMI6qZdJvT4TVa4F7uEGPGlypu4RnqRLvPW0AiFfGb9njymGQE4S6jH7IXKu5mAd
UyvJwMYF72VaIHW/JfwISfpbrCPchpam9Xp1puLzZFWlFYRmOSqqw4wBeUUzFMtC
8FAKFQ9osjtofjdxXIWwfmWOzXutWAwHWcZv8ASYLqAXXJOYV+PPwcbeWxf/TIht
yFkp0Xdeg1FhTWt4JJjM+xHvGP+uSN92lHdj0TuhFEGBYAOtJMZDUvBoacAGRGff
DO62C+ffYS9h8EF54MH2AzfxyQa7QU2WLJ0TF2FnJ5M+gr0CHzuerl44JSX1QkK1
dOc4AgV+VWs0EPTF2VHJfyYBraheAvS0RtH8Lcz6ezV+DjauiQhopehzKLnxY4QJ
nGWU4oUEY/6YQjnY/DT4f/sDNN8LphueGsw6m21nHFmQ/tOK2vXwXLXVxFqC3nn8
apLrE6Dndf7bTvx2DbsTas+3Mn1LBIZKWRy0x3sEMOml/2jxkZJv0CDhbrmFEUJJ
353gxjZw6DHpe8gkbjPAwcC8hOVdjVBv/MGHiMCTw8vd57rM6fdSgyj8As0oHGSa
EBP4b/z0sLzUT5ZaTQhpuSRjZAvEQtu6sDpE25Vso5jiF2iItV2VWJdjr/39EXlp
qNLqkhTH3/gnKYhDHUzF2A==
`protect END_PROTECTED
