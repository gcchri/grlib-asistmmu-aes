`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
StxPlOdYbj/OKcwDn+jWEhFecZ96qQiZ5uUu9m60yyJk19cYr9T/cF6UsjAJfF4r
Eg4qytsS8RmAr1mmkYodOQqCFbyObh8bk84ny/qp8fb+MT7RvHg4Azz+SuT9JEzy
YKCPjn0m8ek8qNkTz1phaBTfT+PoGEe15l1TPeXiVXSCgOfKyOyIZbAm7p6o/I7s
lfi5mg2I40eUJI4z3Ae582pT9q45pUQH2WdCheMUoe/Mg10y9n5q43y/yeyKUdS1
t43cPytUgkCqP6LZoHfxPB3gc2W13qRUVIGIGGf+F7c+pveEZoZY4PdqO2bK7wm3
5lnTP4x72SJO63UFLzUXO+qkEyUy2CvH6WEwOnI2DECzyxU4NiHIY6o1y4fF2vuG
Ud97x/11UGcH+oNRgSkxgizxrQjezGrN5vRbyomKC5rrQzH4HRvkvUHeSXExN0Pl
U7Ao52dv3H4eaJH/pr+7x+1NWKoButs/MW4chGwndYbDB1uUsFUwerLn8sWLQdXI
oqLR1v28d7+InG4d5JGDdNMNEubkcGiAfetsETT8DSn0GWcN9YhHmkjhw2+yA/z1
XE0TEvsih0tYTF4Lrxs56atElKLPRD6IHMONeMLLuD6SNwUJ4E00mLNQ76O+1ZLC
ESMHsbqA0Jr+LO45y03JHiWPZj0qDYJOoKNyzYqa1MHSCjbGCinl1jjLh6NQdo2A
yKnZQAPxBtcu5qc8AdqvZQuXG1l7b3sGGSivwcVYB5LJIJxXSVEZ4AMwnZ92KtNT
bXrqMgO7Jt9DGPBb21+eM8hGyJFzKxvA7+1yOwFIkfrtopBfSWC/iJ2sxeVptYry
fQE8PoLXutdXkYrboC8AzAjkclvLt4FhxX8rzJjuRnU5Vg+tG/A/duU2fa5bgIUw
JJ75a+OIkzlTaHDy05D3su5fy+nNAxf41YF+CZTdWPxw6IJm3KXdVzEyf3/k8HL5
viBdOB+meVA0DLkVayzBWzXcCnwF961bOrMuG2bsFY2dKDw8Aq3lslLYD9E8FKiF
YjgYKIcZDj93Onegmh9iAA==
`protect END_PROTECTED
