`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wBt1NZOZ4PsFzgWAQq4ZvLCDnH1H+3pshwhnNeMMUGpyEnzeaxh1Q4/saqaeSTvY
bK0RWP6vU5ZZtD57feDVe1qi3B5u+DmNG/FpiFJ7JdE+5qWfnxGKL4Gty2P48GYJ
jAvidVxUs8HJ1B54J1krZSBwAv5ESaus8MGIOncEAn8xwjSXid36amcinkTyNx+5
tUIg18ZIHW372NjChGz810FSB7d3eshkhi7qP65Pq968Bpb6gWXr5z13jTroQ2rO
9Jdv1f549ACM224gDIika/0cl3gplTTpzaVh5hIMpUQ=
`protect END_PROTECTED
