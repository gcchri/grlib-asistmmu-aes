`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8QtDyqZO/+trrsyrXHBrE06nY9At19ofnkwEA3s+UZrMjTVPp7LH5NirQOaU+aqI
52MxTO6zJQeEFvs11WuSoz1wI7fwuQoiGKneCWhcz/U7Ja2VfSiDEz9eHE+dRzmw
VInkLACOQgwiM4ewZloYVTpV8RAfHVFv0Y4aFtbqt5gkN2XJyzwU++m4k89EW/U6
2EJi4hxDpdUfIl7HscrT47q47O00qrfdXn53j56jyzaXnExG6T6iCBri5VA2uReZ
RPVEK5ijwRMzhQRQ/iX9iwCM120wsR/noSSdyNbDNuWcjlsPZun6Pnv2N1Rgkejs
N5Ju/d/O4lnffNCEGy/mDqs6QB2DrhtZK0YbRDe4NEcHvYGkQ3ZXoR64QZsb4Yom
6RqvKwk6NXBRGBKgZw5sfDn2ANm7EEsPlnX0Ayx5+d+J1iszoXWD7tj/FPXx5Ciw
8xs+kTJzy7Qt1D7YCoe+ovzxZQjsBS91xlllmnU1+LBaqEYqnq5ETsTGxf83lLDr
N3+m6lmu0dK3/gZlhBA15BxonQinisq++HAaQT766Aw49VOsJjPAu7d/8KILthtw
i9VV2z8lb3E4G/R6u8hyZJ+D+j0umhOlrUaue6vekmilj5R4TPJJJtxFigQQZ9IP
lhHdhnCI4H8aNUzTYz4hNavfCC/mSlxCXZMTOJ9uFUWrANcHmn078mixFvG4Zqff
H2RStHeqjtxFmbG1v0Ul0Z42Wqlz33R72+FPD/wIhq28FE4Lgey4i2gQNd896nWT
nDs4kNWJwIEW19pedjsMdjY/cLUhARhDwAz6FIdz6E5z57leNpY++prFsY4CY557
WTvkMJaKW68qrupCFq/BQEG3KB0kZ3dFebuqbSR/O777A3yhTZyghU+2Qts6Rdfm
MwnENzdfE06H85AV0wf0762zmucTqYQJLAjcBuVdYz8ooaBOwMpjAjpJm+ZHuVR+
ia+EjPGamVSPLgCLxgSLly0RuBd0TvnOeag8LhxQCXLoLbQvUse02eRx0S/97iEv
kuBSkQV5Y9CMEQT0yftXmgAO+DJh46SGTkYUL9tammztgTvpYKN4p1PYThqYQA/1
QEpiYrlykgNj/4zTCOv7PfbIJoyPBBqU33QN7400zaLFNx7T+2ImdrlLYk3azQu1
zlvsT/c5YrlUGnil6Vg/1Xla25pSLVAYxHaz30F0D9fq9unMG0WKNrpBcxnZeFOD
nkwC+XmXyLIitURBkKbSz4155d63Yg41d4WLE31RvA3lfATj1mU9nGfU3kPxcOjj
J1NK81mvrWA4BqFU/6rvl0SGTbrb78LoBVZIJ8dRkzceqRWohOA24QbuU210n5Wr
VwFqUo0MPePs4wNvDtJDkiTo/hnngm13yh20qNNlsBTh9xoUGL625A59IdZ0VvuA
yf8T1yDq9VcKcusy+HKPvV9Izujf+zd+lw68R8DjMXEmMGpZQNcQ7HeVc1E8z3A/
izjC1jaoPpE9QvIT8aW24o5LIds4PgNG3f8cMIYPiS/G6sB0uJ2lNhkDRWvJP6V4
X+XIgHUO9vSe8QBomACinbprSYJQamGDfJYfYmrH7cGR+8h4ASGx2j0PtZmzfX/N
Unyb0SvT9Q3dcC6Pw5LKgA==
`protect END_PROTECTED
