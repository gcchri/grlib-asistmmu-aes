`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
phaH9GCgcdVbVQ88FE3H3aweY+6TfFGKc5ONBU7rsriwhjhpEXq/dpyXocHIO+aH
z9l8/v5RuiEDjVQ2QdC3BMILWQCUI2ysAe97/8zSjSiFV0/JowDEOpiN4xM6Tptc
JSgk68dAcLl+ewa6Jj+L8mDw3C2djyNVPdkaWSLzVgAIeoH3StPwZ67ppsmji1qG
Bdg1aCQXmnnZoMzv76Nx1ougjSvPcayde9loUCe95CjktVs97BsttTzgAJrVVaMW
Cl6r0CiMIRLmCpsFfwuHB3RV87SfEjjX9wTrKZtedd6X0wMvT2vQZRYhyw9vUK4s
vGvYvWNhd94hGwiD/WODBg==
`protect END_PROTECTED
