`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u7Et8e9vpN69vxZILH/xIATBISLbD8DDUaGaGEjc3YvnR3NhbKwDG+4mChSzHQvo
lOXIviR4w76Ye6so44Zzjdo/ZBQAAXKu2lKucKd8S5ct2iwiHSwIlAjAyjVYTkqA
Lxr3K24EyN8FaKssSd6a4+HtbvAw+z/tScDLVYhZrvT9+AVAMysei4AQd+2N2R9w
3YWJFDREdXR1/3vfKfUWTDjxxNW8Wa2uGRUfL5Yn2k4aYmXvNTghlOKOk2y0g7Mg
XTTHLj8v+L6UIkkGQEf9kgTPMLFAjIJ6to0nyStgt7aob8oXdID5sfEG9NSe6CC8
6UJOXKwmTsnfam4wLq7f/HUNXF0KPZkvlFI7/p2rjVVfLsa9QBTnOCvp2u/QMcKZ
EpUqxBfRDC3+k/v3+a/t7VmONe0mw3nlur6H+hWliCHknPYxdEeqrMmuz5docj6G
DU1Wt/VGQM82XDHAUvcN642YWFKtWs0B5OhrtaaDTIQCbC63fn+F4P5tZU+r4BbB
tPSgcGw+aeNOazXmd9K6H0K3sbtA0GDo5Nn4bDZx4oaBgditJj0gYDxFRNjYalvT
oMGanaW9Y/mtazJcAr9jbNOe7CubHO3qCJcWRAiSWHAiRWEl6b9UwuxehecrZ6sl
7SxLu8GoSiq+U7m7vIa4q61+KBVXIdKL6uN2bxwZtRKB4z+GgjiOsXSJHyVFeVz6
+IbTwGf6XxDQEBkeEhBYpxudLa3bW4WJ5TmNwMExJkEScZUj88tuGVqsJIUaKoWj
+gBhIDO46rKltgCLk5LLT/Pt7S5bQiOn9LwWEtSjN+Q=
`protect END_PROTECTED
