`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ICiEHtQ8H2l/xVVy+kPvqqjafQMCErBMajXRm2QP4yrsF3OHPfR4iROw1AsbYRA/
LOPKoB8pv/O7gpfbwe1absIX7F7siMkZEBu+MFBRvF0+2rJkh4PNi7RHSg0Hz7AB
nDBkuZ4p1+XkcS3QBUeMDraaa7yP94zEQWMje6fFbCarXEk4QmyRFitnoysaWPWz
dDNchHubVAxD4I2bjLTJ/bIh4hPfLM6CZkSL1ulWqdRiYnw0gCNab/Ad3jXhjXt1
1dK71QUp20UgjKhuP2CRCkSE6stwKj83rh8U/9OJszbDvdA8geAAT5YFtrVRF7oX
lNPkxHGjcO2nQ/JdeUlM2do0d3qRxM6736u28crRapjKwCx/JSjBSXYttw9+EBZA
r4cs4H/F1BllRSn0/TwtIA+G7lirHRS/i1C2tsUcEPZQUyZWEEkGgBJtf7DRY8t9
8v9hwJoUmVv/IBaW93SylxH3MD2MQK0YYYdSU82lSbuwUbRwAlO/9XMYOy/r5ZWX
jnU8EzcH/k6jPSBznWmu3vwBVhhgMZUaaUoXs6MSwgeYIxpXC+ywYvEFdf3JFasp
/EKBgNloQWCKwosTR9u7BIAkalwI1cyVrCHhHCXbwg0I6oJZHEbhfcgxzh2cixuL
2U/qbaC+RdOIdPyh1Myw+lvQvb6a/cyoF/UqguumuB4sXnqqO87FrJd65DZ2sqgR
GgeJLDK/LQi7B/w/87NgAuMmzhPDCf7hQ/vXK/fIe8FU8U597bM7fuscttITllys
tSXEd19RL33crc41RS8MmqMvuyEIJ7Jd9G8LU/Hx3IV7AVYY81YptajRV6TMBUEF
KzN+oCXpfXuZ8lNFxEvyGZgztk8XqYlyMBiY1E3DmaFZKmgDACvFx88H/RpiNqBP
6leXDWtAdWbmaEiZZKVsROx4w8pcuekOWXAGin6a0gBGGBzLqN2GvIdWCJehD0VD
`protect END_PROTECTED
