`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N50r3u3K24/UfuTt+0pRFUDAaabk8LpdzNLTGnuTTvvN7mYiDn0fbHj4Z37JWtGm
pTHaqd40A1MfouyH9MdBQTiTs15KFP8fH8CNi1U2E65yfpTWB8FABBtZEbDGHIfg
D6IboNKpqoa7HcdoW8cEemNDQrXR4zZpB1q7RaWfT+FxxwnX8y6l9wa6s1BaaWT6
2MBEmTrQ9yyEevMMbGqsaKYrKukJj7J5PPzVH0xLY+W9VR6/8qaCRJPXQRdUo0f/
xcHSAJKqqoMFMs/UTihAOcO5JSSeG508ffe9z1dl/0CXEC/Vkt0rhyQFo20IS8H4
aUZa2zh/ykPKXKkN53OuX/vbCleY6F0BEIAP6j5O09T5I4fCJPGxWNn+uXQyXGiA
qWxNcyaL8yXDH0pVwQYyWghqHGpNc4N1P2pPuisskTd3WKQ2rUT5C25fqMJA0Xc4
II6vQ6H1oUzcJu1Tv8Nl1gCVWJn/6/r7h5Oxkju+Fnnrs/zQ6ko+KcHFbNt4l/h2
LWAvrLS2d1EBbHdvHINJM7dBS93TvHwNv47+1NKZqo7G02BAcinSuUHFQiDwfcDw
GuuQIvtl7S8PP3ZjbLczR+DnnRdcuk2WvZUjn7/GZLvnPaQ82kjK2ccg2SpDRGiG
pm1m6P3d2+Y8N96RDi7R/nwVTlD+V335buJ5pfeBmxGgpDdPff7dSgaT0ltu9H7v
6kbIHn/GXLKRjnxMWN26FAK7s9KiB1aZgiEoygsobzFuBRr8Xh+NljpAOTXI1cF8
`protect END_PROTECTED
