`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
78tuXUZlMdeXcM43hT4fFDFmBsuo7FWSCwP2UByAgKkMTihWAefzg5+F1Bqjm0iz
2hIByHi0dpvWpDdxyIlLsV7wWw4X0NdapiowIO4oeObzxcuoFLLmX30sDmlPqKto
g/9L15okDCV6Df+K9G/W6ThYAmO3+L+HHOzIUhKT8NCPPlTGoDFjSliEZMSOVL3/
t/fhvBvvw7yvjbcTsLPPxtCnk5LiKt4JWeiy6db7a+hRQ/SqzmcwgqFd/lwocBLh
84JcyKTi2Swl/K3IgN5XFltBsdfSfr7LfDlRtu3h/7IeGPYQg6XhwCoSbPg15xil
Omlp2YHnyN0fkfsie3rQMsrUAZ/E0XerBsUes9OSr5WA18TiWu0nUso3DjbpWaYf
Tr+GKd/2r9AwWyiAmBdr9Xw9walKBShShTo/BBaUWdYnyZ8b0GWyLfF5luszdhES
oQnbNN6yUCvhn6Vr7V5ZrraQia4mkYOdS5iUZss0/7voymWCOaxBXnKz1RTpk48p
vQdFeHcgihi3RuVuP2KpV92+U4VKSREZEEmahi8BvBcOqkW5uRozBGNyrectGjGl
hAs49ie+tiFBK35kgFG8kaTJNCSwRM8BhYx5hBucKGc=
`protect END_PROTECTED
