`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZoRF0/CV+B/slgArW+MyhlU0u8/YpA0HzN+wr44eQIT9CEqX/PsvlTgPzwcoeQPl
fFmJ6mGiiWsXrYAro1mvSiNyx4h1BtJ4PNnMzAObEDvbyLUWPaxXF7iW6++40WB4
K0GeJ5Y23kkkCCGP6HtRwdP+rFhLfSGQSsCHbpY1Z8CXwMf7D95wt9y/E/I2mO03
vzrAwenoS377SYzHNZpw5Ya8U3R8m2nuaBg1+kWfYmJ3ReZ984HeNPdWV0uO1xWV
iEGb3UJVXUdwJKhyGo8ZiMyyMgexBM2H0WtHQKgVCGY06069rqtajoRzQKJ0aq6D
Q7wEprBIPPaPNspPkhVNbnl9/uivW5mYawkutnYqAK59JkQkf5dq3G1vOEFQaVH0
2eGo43tnzF2CxIFTe9tfRzsnNBjGdqwsWDBJo5um5mlExBdDAW1ARJYv5COdMKRj
3XjleMyOTMKXe0IHYOJWYh9w2SesiXqaho+EpcCPK8t+KYw3vO7R2NlJOnhNeW2V
e2uGOkT5Ta/B2Np1yTJ5LtzM8dNhCYlXZTpI+YVYTri0oEJso+Ib1ZsJkwpRixul
CDztcf3O+wLetrc6bIQySdUileI+DOkm0DUAfGM7nAaOPkpcLdC3opowSfDrG+4o
HuhB6R2AAN6y2X5lqIOFTW+Ci2UjW9PWcwa6ETeKBs2Pdcz0pbGnds/iMloSzbQq
lztblG13XvFCfIsxeivyDG/X884cn1NiTEkdnuq1UudOHuJFBCSzZoW4wV48K9Kg
d+7sPk5gS0KXy5vatmpRZRc3qVIQi1gF7iqDJME0X3DBGCKydL/vgEe0DNIodYga
gEeLeRhs7bWZdKJvYFhFgWfyN1rvwva+S3iqK2xvoW0S0fnplun1dqwKwNX0Fdoo
HAiEIvX5+ha1Na2VGxvrpruwt0HpUfoaY4TIA0lsSAJAK6Kr6Jhe9fqE+Rlj60B4
CCVf/uD3AFku24otg5dh7SIJi8pSjqTj5c8Bli0Fx/8CncTSWECTXC5u1Bt05fr6
EMq5y5K2HJBg3oNtbC+xxilTWD6xVGhxKsS/XABFHkhFWcbtc0GsIqunGZeJ9Cam
`protect END_PROTECTED
