`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4O97bLMUQB7OmUsr378IYm4JySCuE2ooTq9gXmvmTEVK7DsPMU8LnKKym6hvOmPS
sW4tSvRXOHIqh61i5RQy0PB7GLpRA80kMwyX3LZZJWSoP2aCRaG+eEEP9E5fhChq
CQi1NXgL8jjjfpDFnkYEKPvMctDVFcbP1Eu/5tRJsJ6bIinz1hrma9URyLlGwa3s
Le69f8KOvoavF2DN4YSqxvQeYzOVEB1FgwzkPh7scYI5PgiWBMCv5Oy7j4S/L29o
/YSMc8LDef0Kw2cEc10veMPwM4DAV8TAR06fhsk5Wz5dPnu7ciTNyb79UIySFef7
98WyY/+QZ3tBgFZlccTWvGzSTJw7IUybqrd1U1nUthrEdOgaCvNYey4hJJ3WEHHV
nKdUGagjGTwVUPmwew8jj9LrOOQOvaN3ffBevk6gnXtg54pUFTDUZsrtDgpdoukS
ym9WuJnmV8rSF1DN2BhHhdHvOlgauRWXKxpDmPgsIM5lJtSgeADuZAAT+tEfDIVN
y2Ug2P6/SjPNG2l2XtESXbgV11SQXiKieRwNNY8qsL9hcLiM+XNeVlF21mAKyTCZ
OiNq6PQJfsTj+PmgN8+4VpySvyQWdrd/gXUqLPBwAXE=
`protect END_PROTECTED
