`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
prKtQaS3WrM1ScDqXlIrzZlZQT0KaGdPmEK0lTE7Qf/TkJ/0VroWddiy+1BSEmmz
WzMtDCmN6U4naCD+dKT+HQonO+Q+pcTzB6CxOplxQZjJgg7iHolhxrZbmK6mmwja
H/KCOKfR+xcK2j+mTQxpnPwL9QWna5TrTyHPbhTqYLC6JHqlHJTpjRNZ422Piu0u
cNDLapPziFtylB5unxCSwWX1/7xScjWj+FvsXT1NAw1pTaGQFjrG76fBq5oOmZn9
5z4kMZVsV+dnHYLIXsXlulhg8GPFrg+B9veO3FI+bfRyko/PypOQmwWu5ILRKCF/
o0bJ5L1GoksgUJcAwQ1Q5fa8074fq0fDD1n5e1HVfmycImSBN+0kX5cmovwFSghH
3Lh9n+qj39JoA7fD02KpVi5KrkEz3eCdQYzMVE8aabYlqEoiorwICYRUtyYiaIc8
HAnslfJ6Nc4UFDg507tZ7yhpxhLtDunbowOI2E+oxzP63HTkkf3/Dz0UMe1nqO8Q
lzyb133NYxQsLZDbVe5RAL7yhRwusrAGyoUfm/seqo89sUSdomXbvusq86Yf+ptD
SYTfpD7oZ0SUKi6XJNI6dmHHMQWat+ZgyY0b/SsPrsfmqODaaX0Wte/a1vZ3P9LP
o10XSTlMZ6d6pSg2m3Xt3htn2LeGZxxAKfBjXgvzhXcP+pDjKdaQbwta1Faz5HNT
Ls9XgXroup2CTSNjW7uA8JBdyE63OfPauO2mGjP9x6vexOueCs3F7Yblhvfzlnav
2Rrqq7Sx6WMTFGQfouISSdocNhnTGz2w1ZEzmB1ITh7N9KvZ/z05LlrhKZKAFyga
BMg1o4Ox3VXgLWkHSzv1713Y6PWnhtocsigZQ/R7SVftbVMYfdAscNSXNlkG3+mr
N1Tn6X2zf3VD7U/x48igM1kRevKsR7tGz0NsYc+ZKjTr2CXOkPHeGTVjCbZtKXhv
r854YtF+p0PhuGSvhZaLPzS47n+kDna4C80a6XvrEJSIPZy6gbZq9YIygUxvWMeS
iJ7NNruEv4TO5mFp0vPtumR6ihhgER2SyUztnNPnnGonTa85C1XOulacC4wbVbi6
iiaz/J1dem+0rzc5wsfaUwgYw94lgmmAD2esWIVD1nusC8eixdgQYIjTAImmrWIA
MISbJ5+IrXPkFW3WXtaXRG0tRCnVhg1CH48VfzkJTxQjZ803Daok7UCgZKULIXnO
1mFzNxyub+D4yAWsn2xeOBwJ0V2a1piR1nGt3EHZjFnpSlsKTbTsjYUEXVfRToh6
eldUb+lIQGtNu4nFXZlmiUTwj8Lz25z6pVPPqzE8mfNNskT7Q4DhuCTe7FIyoA+T
3Jrjy9skRUVB6yemC/pJoltHO7j0zQapW2oa2JRLwvklzTHsrJ3ONAaNVD/8o0cW
P4eA8oZTTlzxG87SMYtzJ837iPOOrV4GZbwwJqXAKMPl7+dGXLKnftNnRIz2vhm1
3QqOA2tN8Njct7t5nArC98EaSBLYqI+0R1M5WB+8A8WB6kEfJ7dyeyyROtk5+gRL
AFRCljrrp2uRIB9uqg5NkWmDolO/3R7pQmWXTZOAmh0Kr+gZdr8lYI7rMonfxtDg
hmRDKbk8/d9pjEnokVZZp5tCVxcdfj56+yMZOMxcD+FmyuLwfWPyIx8aFjqTfhzb
3fnoMtF/zJ4izj4GktkfqHALUvrbid4go8zeJvdeKDBflSpNZ94p4Q0kQbKj9inU
bKYDZgV3IFvAJF9XXfJF3DOn382cje6ZtvhuFtWQd/pik89i3LdLpytXFL+NN/M8
evwv6CSHyVulnjcZyhU28qL+uz95QKby/OMbma4e1ozDVTeW/rW2pieh/zNd3FPe
GTsBNaI9MCrFnUYrMKhdO973BEEkIpy+1fcajisd0gfs+E1Df5cARCtLT66zV/Ia
JI7IWo84rf04myMCbfu8LtCoqhjcZTtCpD7CQxglNGYp9/M9V9jT2bu69/9yVh9C
Xr1d65nfgS9I7osceNqIX87D1uGX47QTnYNKQx7k8Kz79tEdOh8rCcn1pXLJeN31
7oFZqx/GdXnTTQyf8Yp637ov92E7Kb9TlPO7UKR5St0pAG8baImRDXvzatO4ifh4
RKe1K4I93loULC00ZgywkiNbWyK3vZc+cRbNoxTuwx4Zz+ewOhF9A+IeSSbmSUFc
HVrWTkpS2Klk22lYcyY/eQKLto0xirfBihPnKa8MXMifdAEQTAlLdRN6QudbMMtH
zc/8VAxL/twew/+zHCJP28DjeIlZeFaZik/b6dv+97L2Odk2/gOHFicV0NgfcJcv
KcitFmn5DPkyZkbuuvVp0DOZWmXgwNUD7VZnx3ji8KuHLCGXMOATi62YRimvmE9F
UGcCqsrdIvlBCTqPTOjt0BcmP3LpNTNIV0ek31vzCHetUeh0pdOQdzr+DOTgy2pr
mTS9vp8uoh4V7gT5BLSM4Cghs3agEjgcfyBTcpQGsjEAEToMERnTZdvLQO/+mLCC
JH+NvJo01/K1HPYeb5ak4AQcDEXwPZ0K3GMnVTbBj4aCRmFv6BZU2bpFEoAG6NMB
hlDF26VJ0gaJTuN7y2VJPKMPm0wm0pPjhlikGKjecqfnisSXgYEO3z0P19vdVAZL
MeXjV3k4aih2mMyspbvVp2nzfjQdhYZ+iaFqpRfZzioeMgMKixCOvRdoHCbtEVOs
29pFpN8D1AXVWGXkv/UBBAFcKdI1VcBEX7SzfQ7nCIIgODzaYh5wuya1EHjOAv4d
y2k26x7aYoxc2i0HHjJ+XYOijpn1oaCn5sJXWFJPTebTpl735KHMGPM0NcnjJ2cq
aXr+fbfda4OJYxN+4IlvVmzjiVpOmrZvHx7zycpngMn6pW1QtZ9naovDWMNwL2y7
W4OktDOkH7ODkA7D0OewPrkWZh1X9Zv3r6b6E0+10W1WBxJZmLYYCJ114uqbvDAJ
Kb9TTQDSZDo4dT+GAQXzPJ92rgbOKV7e1QFXNJNdRlxv3Hs4SE5JfTf7DIxedy/x
3Ix+nr5gNgQbHcwRyOVtKtYmRPa6Gg4kPWUpLnZcTpxe2nV8ZK3Tdp2LweN7Q7VM
77xizL7r23ct5/57WBzwW9uRxY5QwM3IuQXkGZBjOD3K95WFjGnhhxY8pe0L06zj
/fPIs6tdAg3VZdfPWnbu41LggVLpkT0DhtQp45Ax+Er0APZKKcanZL+OByVkDXsF
uun3qwzvV+2AiFu2DvBf9DzckviXgUyzgQ35wSLcs+cL+sH1pT3ssd4DQqeUdMvy
zbwpRHo3EgdYI5+HeS4KYc+aVS2AJ2LEbUkzkXqchCHTZ+bKmOK9riQ6bKyZX5/O
k8B6cEhe0JDx12kx/Bw7hpLA+k8LVqBBXGiyftZ8ORWUSwuKgL1TIzM39X7uewJz
lq1IIFntfnHqW1hWeMQe989hQ5+hp0uc1vXQqX6YUadHvFFunY9DFDEZcxehhYsc
F6IDmH+xLbSrYU1A2jQdAElzTr8jDp3dcwHW4uxmykVVJ8PXHkBGvFfUjsx5D+Ve
liv3Kf0npvjs7zsGZcoSFDX3FXhMjby4z/+UJxrTyeJ9iNRVaBOnheLq/dqn/NL4
4RAgf0icnnAtLF0e4WohXFj8zL3dx+2CptJsCMB/I/JOTsDEBp6AW9ybB9DBAoyi
EEcLfDkyWWzoldgkKCOJbZ6Z2ZIGIgvkBxq1ZmjnXHuhzHuLT0CBvREadMVquGu+
cgsaNdqoroeV6DN5wJmTXFcSwnJ6IXsy8QhBgFD3zB6MTaHd+L2mOezVv8p9ZuCP
BHCcofq+AIyiytp8CczAtdldJg5Rp37FzWercHChfO2rBHy1sdgDphkFnLkeevs/
nakoKrff0rFsmeLspATUqvhqHzT8Ya0gSPZj2ywvPY3eOzNkIaIvQixKN9anXNpd
XHh411/rlHAPxYa8/TsX9nM5nMWIlAuJgxKKMSadWzMKpfFGdqpMdAx39XS9eh2F
c8ZCbYDd6Qmwiph5TQaXgeLIpoAAuEqEu1y5wDGrXK8+5Z7eHJDBihsev3Mkl+4o
1uMvjUnslptR1lgXsbD/OUOGNX9tjOb5DBTAnJMse6ZOUguyLNRWvEwXpb3Y9PkT
NcVw4PCa3bg/c3/W0hsTghJjhifid0sUh3JpvFYt57x9xStAlFS/AcVwZfNzI9W+
ngR3flfnmlJKSw1datmjp2dlEVRi+wV2YYLJ2jt6aYMhLGVulBCcNioOoCdskWrj
9nBTxJq56Lm5yRdq7Z+OuWstOZjHKQlzEqOryauY5HuQZgkwgTtmjW6obOnS80jf
9G/kWDziMHjyToEFbx4cEbnGQZrrrqTfKMU8JCmiqg3Y3sthEMk0wmYdHY/ADTXS
YLqqUD5cogLZ3JGSAVCU84uFdWbo+kcW/wIJBCOTT+8wgAOON7KyJP1aNILK5Z6I
XrR9BwII/b8sUtkW74qXUURJNVNQH3IVYB50T894kBpjqCtOEIbGq13ypHM0Uy2W
3gh81yDaRDvAGV348ttOpxNh4XxWjsOyYAdS5WCMe6x7yXoA9CdYa7vOZ3N3DwFg
UjeSatC0n6ZoukenuFeUm8ervwy/kEHzhY6NosExzNoM4+S2+Ll4E32UQXXXJVyt
IV/YzsJilZdwzV8lVxCa8NLnSCZhn5yu+AJ1MDwQi90NxQhBbi/UN6ANH3ue0clv
085BilrJD+vDascLdQ7RwYg+K7F0sV6YiM60vjvBybJv2u9uxstlH71raajiuupJ
u8apID9HY/rbuDoclWHXZ/1LM527C8dcDeKRgLDnSy+bwpDCoxNdLs5w1MK6uC9g
gklTsfZm+1+v2SL6ay1Fd5bHNa+IZtt0G2E4yWKZdE1HBoq1YOW9qvGMUvqZhUgZ
7k7pZqbKNYEKG75IfaOfIkUMx7vYBEpR2zJgsZTE9m02HcF9fzmyuyVCuk6kKIsx
Y67PRIVIeojHXhd3wAitX+GutZIXhVAOcTBOEXotvqt04hHE7ofXN6pn0cI+2o7q
02OuF31x1fF9FhEy+MaXJVF3QM+MmfS8l9hHaO/wIUCx0/Y+idbn0pSYGUGuVZ9K
uKPheD2UJgfzr04pqZkqHRGZlqW+S4Fsa6PpVqCuJOiT6Q9OtxNhx0rcnU3LX0V4
+3yCTMBRAHCE93/BUTtQWoEfjBXrHiHcH5xshBvMnUDe53GDR60Nbtj2m0WUL/sO
3lX9gP8kniZufrLVp4gqds317ZTtSl6ztP5rcagE5hL1xxKK4p4Hi9agIrSiDpzT
o4diAWUhbXDM/yg1OZO1IxlS75mYEuyzHrKD83EKpQXivGap06q29YOI8QZGJcOI
ja6qFzXF+2fXMfqTDhI7vTNd1ZNCAitkdb5053HB2+0SABBPKRRgwql9NTStfiw6
yARozuFPXIC/7IsRXEYqQUjdZeOI+32HrAddqjTmr5TMCJL8zvaFI11tMpMpvd/d
/M/54tEdJrYoqrXbJHtaMWdHafuki+7Tg3ud3FUWsngNNFU3uCDUvKrJRGKENWyg
xNrCKO+3w6KPiTjZGIPz8tvkkqrxmXkVyu3bFgsAr53EYdtszoVeKNKV/gcAvYcv
Pl34dUZrdY6DdNP/dU0puNR83ksNrZny3pE1l3yFk22825YcYIuPgBL4xKjdcnel
`protect END_PROTECTED
