`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wQhQ8cEfYkGZbV+L0SRijjReUB6IZFMKCl8goe/EGG53SaWF9524XGpsq6KEsliM
oOAlgpJaDKRzTuw63G44uJw6yxZV6BPLQaQIdMMsDidCkD22hcoQqlVB+fcNqU1t
5qMA4hSPdz0ER2Axzc0vkqswfON8YDS5QoxXytGffAU0nG3tXhtqDOucFSLCiVe9
j4he35n7/u5x8oMlx1z3AWhtiHMPKAcATViv36dRfJR9HJar4mGFHmx7Vnb2AJgm
ID7GZRq5cgUPJ2IHpsl8WyJL5dqbOMmfLuylZhDKmKYvhT/0nQTGTqOWwvJChry5
CHVKNtGuBlLxuZjBFCaaRREjtd0SN6wLKjA37RjtM5FkSlTTkLZPrabQErLtiMa0
9oZifEqABtiXlY6ZsxQgl8Axeur0udl6VdBpwcQGdJgIIhkZvQ0GN2cRAzDYWDHZ
Ut7m8pGJCYHwwzTFOEc/fcAVi/5un5EMPM1Pa53TGQWk2CK+pd2bF43X7hB3/s64
mPJb2UHqMfMB35FwzKaFnQ==
`protect END_PROTECTED
