`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sX1JA1aijAp7MxGttdUKoHCTWelR/zBFRFxtaweW2HwHygEI3azs20XYYO/hsCKR
tPi0SYfAvHAQR+q+B/ySaNVfODUtk17CBMh9x9xAubRwRxlgCLxmA5Vy3HuJZg4v
dPf5EqGbCfmGhlx2iXsZcoWJ9+Jk8kXwH+nWSNY/d2NbB6gtpiYi9VV/JvI7Zxgo
GNBhiBlORsyiZQXuIuaMZWSR14zxZeLhDoUSKbNr3kqY/ElvIsQ7zoG6hAAcmvg5
toJEDTxHMnyA/bp4bbyfhsZt5tWPHWWKyLytuU4rq1/8GJLf9lof5EqwsQJOsotO
IHZvnNn73e3tG+Kgzu6OT1P/CXyoFpbiynvISCkKi/yWE6Bw4aF21wKcYOqEZuXw
Nq49SjQ8CxCw+bW9SzrA7kp4ZQIv9y8gGYF2GdSVLlq92/8s3InSw3BNXpi2+NIk
MgH0rOgGRNEUHIEGZJKenE7KxOVCULtAYeP9H2caiHNxy+IvlKdOoxZRSCGiI4Pq
3MdPDZ5E6RW08gTF9K9DxQvfBXHlyvB9vg2RFlBzWHii+JWDpmvfi7S2K1JdiNMU
KjPzhAvy+uTvcAHqtgnGVYVHq1Tz46fUrdmx8FEAHH8m6mAn88QbfgIuKwgtKyAG
djdSMoAY01glh6KHN9PclQ==
`protect END_PROTECTED
