`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5iKFycYJfKVCAH8C6vBsyGrCMkD6rjfXZNfM5yBNBxVghOIOjKvuaKasZzhADgzi
VrFTmBAQ67d5EK8kSYH26yJhPCKaB94ykmfB22baS2t4m+Ikuf0Le3yXi1tsPTLJ
ZzdW4SMALMS5JkyQpgPKh99Fr5YJI/S7nBdnQd+MI/h/W9uHgezwYlY/XQvX7vyW
S1NszgqtcLnlR383KamfjjOleymnWVkybL/IoERQCLhL/vjP7+DdfO3q/4vIodII
A8+9MgCSD3WE7y4WEV1FUqUGXJOD1lj9m5rQCr2W9EsfdQxi7E06YnIh89fhN0hp
HO5bDigel+W3VjJvI0EibA+g/gZwojjYE5czhsQNcNoqyGagVKcsZTo0RoEKm+13
`protect END_PROTECTED
