`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0zVxvQLiXmC21qgPHu1iWIhqIVH91Cx0GFnilcNoNiH8X7t25jilV5hdDsCanOd6
RlrgdI0fO2ZB7J4jdRm6sM39/HiZlHhwpehhZMDYy2cC2djnV/BT7ufC3sZXFY+n
tWNOBpKc3NyLMNSQmmVPsI9WgHQeTKwVWqx5K6khphSRkWqED5F6h/l6wR6w++UB
pm5WOZsqaW4nzuruVhmkJNszfyD6WMYNNJX9HXT/35L9BfTsn6HTC8IvqB5kIQif
lNQIg0ZSrq8nensoU56WjCk0n5XCqeVqUJMG5phTy4M=
`protect END_PROTECTED
