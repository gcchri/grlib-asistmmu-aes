`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yye2Wg1ICkks46Vga0YPDb/EZVrLIT+K9Vf9+PQDSDZ9J1ZeB2U8gR9yD9QwOGUN
jPlCj3HZ4O5ewsfy9sFj30fcVEra8yUFGeIz1pBjYCM51CiMCfZV7Uopw3/RIpUf
GbJYiaz6kiTBwen1aw097FeomczaQQeEPATbmZefSHN8ycxVFNS9s2YiNZkKunS5
GAiviyLMgcOtpYkShjE4h10VpDwK7AumDWHr/iJruWWQsoBh/IkyOp8KlfOL4sg3
9x4kOFW6JZaaX9TZc/fkP475JwWGOVOVKxLsZOZJyWc/8BUmCUB0ij4Y74cdl8LZ
0/AfTlEzDuwtswv/kUr6Bhgnf7Su8sfYG3ODkdUuXr0qMxUhbKs2JyMR1SjzB2P6
eellOwyFYMmp8qpSYfe09vk3uRtkGSIkdt2ViSTShgMRZ6Vl/jy/1SxEsWd0YqRi
`protect END_PROTECTED
