`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mJ4A1NZE6bznrcc+vkN+Lh492HafUPChF7BiS7Tn+4oGD3yl5tT1EKpcjc2HayLE
d4RLyq/xymp0gj7STg21nonUMLGw0rIsWGejgtYoc7+OGKk/o2Ltb7tWwUFuMBln
8aM3Cbue0NEwsGGz18IMBxrQ5tcgCSCxyr267CBBSO9ycYaon8Bfw/qrugLvsAmj
lesOaeT/skyLjnEV8RXwqeFpywJsr2pzWxmGHFEnDTbeNh0GVuGIyGtA6gW6P3HC
AGGxnCeUfKuzv5N4tkjXeZv1jVXkF1knkBVW/vO1ne4MeYD/dZEQGFW0JW8GLVa8
XDHddeGUWCryGi/fMoIzGSV0r2RuUVOj6xwF/K+kXOT6m6ab7n9+MSo2fzN5Ke1W
0aH0WHrvLHitEPBkSSoYa4kjovJgEy4csBOCpZbRrQ3K1Iwb0tGUQWnbxh21ubcP
D8uD8Yk4iSxjD+hnYDh4/fopB/ySKPshDIFLUxjVYyDy0clPb5Jaal0uRDTS5F+t
`protect END_PROTECTED
