`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CEfWTnovcNUCG+Y8acDwMjbUXXmQJEvu2/L3w8tfvNwT7F7l3pbAlAvsiEUIPu9X
QKHhpWPsQpX42V5YkH5Vqc+Q8AflDbVlv1MlCh3yMHibJozi+PDvWUJQOP7j9QXX
LihBgxDdeDLLqbUYIX9N5+1RpDTfS9pRB7CbKWPi1h9UQGwuDAAiNyzFCB6GLyG/
htAKvIyYWNEzC+KtbmWzqQcI6guNKfFnstmooGLUD9x7BUCT6nE3b5i5JXYcs40+
5ONTZ/aCgJFYWXj+nKtIUYw0umKNQgYxyR3cM5vfafHB/13DxLJhjPHo8Da0hJWV
PLsNFbvoStW+E6YCBNUTlbMFFI9E10vJgYkWQQLd3UsVhAM6ijFSUJbA1Njk8a1g
mvl/UohQ2CjziiR5JAs0en+DHIKS5qua4M8c0MDrB+E=
`protect END_PROTECTED
