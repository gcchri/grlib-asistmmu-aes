`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YoaCYar+8LcQaNSlDCFyQpAmf3gSGqEAHNJQN5CUHJ/kUAfYNku+JqscYuFtM2JZ
R7MIilsB7iG1QlZlPCVHlwyL65QkHInFEP6b23kUkY1gSGh4A7lf1i+/KPIo/HM6
8EiV0pgJrBaqgkrMg9EYWZjv05PgRYHf4uivC9XshiM+EoYX5KbK+lkhxvMMfPag
+y03XQOKq61CagakzWibhPFDYbvgfljtsq9RtS2H1X+qJRh4JxNKa1oYcfcjG4oX
ZQKCfJHbl6b2vT7xz8wX5w==
`protect END_PROTECTED
