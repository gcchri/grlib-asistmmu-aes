`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dPq2DBOy9NOR2w2EkmQF+rcfQ5DghvCworJ8Dt+D+QyscIU5+9veHjGQf3+LQJ3T
6oZ2OOFtoTh2RTy+8R2d44cKUa/etB2ZFBwcJyh/b31XriNv2/IJMM+ks82hDfLw
13IXsY3WJ6590O4/aWbPYVZshuSuW63pTbj2CTuqFk3q9Rp+OPMo1SG7CCvUNfEN
Q1R0GmGVKmO9YXpayyDDsB8anfdQECv0LKisxuW/gjQkiWqrgE7g2NQta7gh+UDt
B9ytNdwIl2eBYe6FVFoEoWmu2Ec28zKwIKlKsFiddrGgjOWF2Ae251C3qqn7bz9q
DbTQ2GV6WusZSce//zz7eq0rmCdl4D4OVVGEaxERr+cbUqGMWAXsZGBhvOXIIMkg
+5fjYfOCnGdpLZ4JSTWHUOOztro8cvXtxAfdmG123Zg=
`protect END_PROTECTED
