`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bbd0qkOS7eOguZomLMuvG/S/tt6cKmHsAhLaJx9AI6P49HmEJMo09mFfnalt5YtF
XGUfbl7SA7Eu2lzvkxWDZ0DuK/cxOtAyl1IFc2GSZUbEta+ccJUXWc+cssdxRG6U
ZHWpDkzognxpMSWoMDyNL6CBCCgxWRvlNuz/IlzzXyvGIPmGYQbcb6WYGD8ZKNs6
ER5XWVqQR1arVtrV/bCe6AD4TOFTmIJ0rMlXGUdTz/UqXtlUHPxBJ4W3ZL8xHYqj
qt9XEUA02Dnabfu+bT8OJjOGTAj+jTqVZ+Cu1fcEG8sWtdDLoM3S1d/0/JpTMFwq
TPtwd6S2i6WL/H/aksTT4ZwhlYRUHHzebGXS4Ck5NuNEEi8l+//+MwBeCHzqL/6+
Ev/+7rUK/N5SLtqjealDENXZyWvZ92jDzUy5g0yo6K1THStxinZKyoJ+gXMO7jAG
/TpuJRQkdioyzN2ZoZ+CLJ+pzrK4ykkGLpj7a5HfESZ+3LFIhtIjRQ2u0zdePCzp
yZq1Km112vxDnUsXYCKVibbXbVCcTxsAzXQqVRBfKZEo1r06T4EQCegHvhLAyWjq
Tq4daEsPKnyWHj9xsKMALGe8px8l+cJMA3aiQ+CutHguvgjym1R0D9r71RIZiLmJ
f2lpbI/QpbOkze5H3uhTDemfIay8j15A7rW3U97jnDEmiqCEHYm7vLb9FtHicB+x
VvISV8L4UdWASqwU8PdXTwP2E3Qv483G76BAujh5iH3wUqnFhu9JlnSifBWcXJCq
j5VcwCyhSUSFBMNNCGI0FJYn/EHZm+Hkh1bzb/jTtY5NDYq1N32ZkMTWsaBl0j+M
JBoIL8URFWXMilvLc8P5EbyKbaG6+FD4x95Y+8WXjqLZVXoIrNxjvBE7gZglGKQd
I3CymIwKFN4h9o9+JEXy0J3hDn4dmup95pX9gOZxS+XoULaiRKxEUSe4GfFBaoOs
ca1puG1VDwzNdYMj4C7raAAI8b2pR19lHSV3TfDYfAuHeeqGwjZxe026aRe73JEq
0sJzCODvUqT2gf5IdwxHvWhgFZXdsmZ7Q+4OBmkxPxollI+D/PcyXIDswQDP5lOQ
UsBtWKK2j+BR9fMUzNLHEk+spH9QXKOqbqttADpfLt13hPWBKZ9qNhjwBIn1R4sm
hSVbxjQ0eoq4Zd6PltKAOK5nygRh85R/0wPeRn1Bdvz84PJfOybUAmGowPELWEWZ
jhzoFEB5bWAQqm+xScu5Z7pNgOONyajg4oAMZTnyOerRYzmIjZcNhU97pStPl3La
lYqt1NBwAqwDPIe/MRtJ7VuYjhheYqQWmy4MCKF1VaomkVhc0VmcnW6v2TjwC6dy
i0aAOgWZXrN1Pv5k0AGdUE/DB0uYsyZt38w/mM3e/J3vYB5AB3SIAWuvBcDaoRRF
lisKTDWAS/7HXKTL1KhNl6sftTs8CFLbVziRYVIGVnj/gqoHeFyTjxR+DBQgV2hs
3hAVleGMW4HH9OJlWxT73MBxMCl4Xu4V6CI8HpJP6nGpJJZ79R87UFoAYqUk+YWa
vxhLhRL2iBrsN8KExgRZ2xqV7vf8gMNoazpRXsEV3Ms8FI0iY8sgymyOwvy/NJVT
GwCZWC1AnO7nw30YFmJhKvI+YR+SUZabSAv0JNyXrphF3HVyeA3sT3HFOrubSX4m
T6qvro7Uyv0+4GLhNSgT5JMRZhHyYk/AlbxWZRyxnh/nn4WN2UbB+NNn/zqGyxs1
hR4y8wjXuiSlhitpWvmqRptJWv6IM4tIgxlHNvILPnLyoBI44qMv0m/xjyS6Anlt
3kylxLPtOHrJzJoXYrcJy4503KMs5P5kWqXACoWIgTaKMU2ZuX7AODtWs2Sfg1V4
tOH9335K6Roe755c1nHPSPSGUl/nouZH+Yb0JLUDfegdy4ygKxmixmSMZHljE+3K
eLbTaBIQd+PzDIpEcKl1xYE37Fxj61Z7mtRllgTY42JBKovOqChBCzAuuy5LMOLD
GnaNenZf/AM9KYpPNzzbN7WJH/QeJsb7f1NUXML5rSn/zSxVvDPE8El4Ue5gWWgk
wAvjoCU91ioy7y+xQjGsF2LLuNwZLszWbzx0sY06RMSfPsDmZNPop08erapr7uuy
ZzxEr6BmqD7yKA8AFMBL6HBiaZgUrJz7Zz0/v+n+XMFAhwzLT3Lw1nVUEFrLrjny
Cafmoyno6GM4/JeiYpmItu2S6Pf1/62msVMmTaaipytLcF43VqQ3em/d81gTMSd5
ZRSX3u8UOiuHdgp2ApeJUK4M22iX5c4aREPtF2X43Dma9o00X8peAGPm3U2W6igH
eJyVb4wdY307vdVUwc6+YZUsOhH6q/5yAM2OrNAW+wwmpEbMTgj1k5Eo+RV8xfar
VT/nxH7l9mS0BVFN24ppQZAD8Ay/BpCJ5nTZOWSXMy+aEV8g56nDsf6WtZhkROAv
i6UsqTOr8aFWkmU2draELV/cs6RvYHjqpk262frbh2Ho0zttYlfH44Sjfjm97iK1
jizaNLT/dUqqeBopkRO2WjCIbq/K4bCFgoFxsDplqWURvKqxAfp0UwwuEwX9Y6+a
wjotXvVqDAyyeucqdOIEXjdGiUAt/pbKOey2cCsBKBui4n22EdYXAXfD8maStIvb
R+Jy/t7spqwu2tKGjfts1wT+uUn2BpHQNXgyWirmPfY=
`protect END_PROTECTED
