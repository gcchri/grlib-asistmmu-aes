`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BI5PXRj2tB+Oxi16Q1kJEHT5truB3oJspOIxR8a+EhGvdWV6iKyMkD9E0tI9A1SB
ZPdjWG4lme7dzlCD4Gv+dxE6t08I/7/57B200gyrwv4PYfkNVuIoIQbM/yX64XPR
ARjr0jiDQFo/xEExxWKkHStYuG0HPZNq4ECzRzsaOebcUHv/RYCWI3E6gJLSYeBY
erKBqdYdaalXZm4aKcVMa/w+GmfWMNEgaCAiUG1MxmwBVuD2b3slXpVURJCmV/ur
smd5WjZRqsp5BbaxvDQwptQz2Zj+T5YK1Ew9xss4/DlV8JZkx9UbpxD0Zfn2RoO7
iC4o3YS6bUcfXQ/sog+9A6sVGVdoUuKYzY03fGzaXRUikueaDcuOfOOZP8KMf63Y
oF2H6fePN7SOoDi5eP33f4truCfPP/xxksOsrFLREjud69bqcckEQRSch4PpnrDa
ggW3SaUC2k+wHrtMYvQiU2e1FpXjcaPAWr8KKL8r84mHt5tdVLWMrUNiB3+lYY7l
/9F/iOVbQ6A7ngW3z5jzkc8+egwI9jH9wwo7Ln39Eh+5FmutPAqO+YVHXT5CjevD
+6PwDpJ74thsSyjakrNPqg==
`protect END_PROTECTED
