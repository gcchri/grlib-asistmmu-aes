`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z8ZLjZr/WVkaaUcyRfLiUk1jrGzwLgLZYtQe/0s8K3Q66aXGeW7OCVGGIyRpY9LP
Unaj4QPyHsiAONCZ+GLHAqb5sGdPAn9/8LkaiOMaSGv5yVF8DNBBPsuFnfWxTSIy
C67bedv7wN/r41GOO+9HjPeMXJnBq04wbWbPbYez+UyUPWDqxT4sl2+SmH8bnlvo
X5vYOoxUU8GcIkCYO8gtU0OVJ3/GYUQdUMoglpPUi+BXe1aA0QBThxNGJUoNeFbl
5BBg/DLwKZuaDHPqyDATJaDwq7nq60TZdQ0hbKrhHkggeXEkkrB2m+Wy6B8F6C+N
Fy2e5H7hvycKGignRzhbMMn8mPOYwfgMWg3PQ8kOZu7YVpr2BmSgZVlhdHX1zgBq
`protect END_PROTECTED
