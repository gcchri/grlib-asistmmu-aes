`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cDCRHu6hvxKUFb/w7N0PLFLiAK6wZKcNgLCeFDsJjJQVRTMRqM8G63Rz0tPSoa8X
PIvYCrBDYrtwJqoHZtkEeSV248WAeQi0Qdo+qKmlmpznPDY+kE0lAfvmldWuYj7t
E85ImEpDuWNvKJ+JNJsuMSMQKf/I4OTBzsCpA6rq3g4s2aBtAg7kjEYR+5P/stAH
Y9irrCYojeGyDwKieqvADpTT1sSlEDHrs4TdawJoSN8yEgakVRvVtWeGSA1FFHiv
0JhEpUEfgr+4qa6cGRnespk6vWKYFxDp/YNNY9uFCjOB1nTd3OvCYvsMuEAOElp2
Oq3gkNY6pVkKONCtBqGyZ7RtOL/9tJPqG3muYPjDGg5ClkMfu/V1xudED4cwQ2rX
bXcR19f2Ri1JiGoE7i7O390oEoEHz5fBnwCNATE5yQ3absnGGI+7IkkDdCLtTvIP
`protect END_PROTECTED
