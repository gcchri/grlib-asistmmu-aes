`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
71IJmf4UzzZ+BbErcz0U6pnEkWa7OQ/9iINhqth/Gep77AQ3UXPWzPJP7dIJk8n/
gAIe8VQClQ90SQCgLkzSZ1vMb7sZNcWedK8QVQSzcj/MD9O05uACJvkQ9CbZWZHo
3PnZOE6/VCvElLodY6l1kxxXrToTJtuCBql5n+G0KfgSrBLJqvuCQKLpl53rnu07
G6HVcB6Vnh7vbXtD9SxaszJQUfbkgJKZq3ptpjNgDBpUHO5+RZUtZ/SDMkTRFVMj
H+OzYe/PnZ0ULo+ihBrHp/0IxTXlvQbM/Qk9w5nne1uHNUeyIPZyWLnpCOMaZK6I
ExRGy4IGT9IaVugvLagBdwMuK1+uRxHxFifSzSVa7lY0wIbeIO4PedRg4pOgnCvF
g35BPntN0wH+NZ3u5S5QSaS8Q8k9e0UtLNGp/xABIHE=
`protect END_PROTECTED
