`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
luV2bMDKGpBFh58XWXxFzzyI7gkUu82yzQB7eyEG8LjonVsnKOfwQQJhOLIzXNvT
epi9VuXpoy/sjiFF7LowdaOClpblh9bHQLVcJsehPCwetvo8ztcGl1D8VwImCKuh
cat+h2RUxHojc6Se4+Csg9SINXCoNTu3yn2Qf8zO7Y7wNXWjNdIgqbXtES9hbBa3
er4yTa1BWvP0GzD7+2WTR8eGgH0qcPFwtk+o3AADUUuSzbWPKKKs3ekGncvz/k5d
B9SraAI6weRGuRVRsO4sZtYtaqCpvjbaPXhpm7szl8j5qY+7MpYqhN2g8NKucpVF
jC03cZOuidtXW76kW39uHA7siACeQfFEk0fM6TkXGw9MiE5F5B5M2bGlYuFezfXl
gifOARDTxDyAOyMXuV4ajc579euQs8VB8hHpS9edGqRTNNmjEoLlloDVMSn4DvAR
raPneWkpSOXWJcNZQ1urCpGY4s3fvRUUPOV/fwXYKGz7/brR/D/4c6BCWa11Hq7x
vQ2B61SINPlo0lJf/iVD+JyBhTt6YV/yghcoQEFOoPSVW7rnmXWts+DtN5KdYo72
W5CZS2EPqmxAsSEHdlV3o2/usVDmGaoPIZtNCdBTVzdKwUVjIa9Rz3SpwALd/XbL
X0+Q0cV8usNaXkrf9wyP3bh06EWOOo52PLV2+M7XjrfG8M0NLZYvYyNnQfmCSwcT
jQm7IjLsB0qOsMIo9Y+1ZTXqW6WdFXF5OjpMcFdL/Ar2Js7nqS1UMYQt1kE2Wcqg
T4/XooyvFkDc3ptDTvOzyHKd6FPuAIE9QOuToOnpAFDqOONXtBlJ7lP6dtkUnnQ5
yNNhAmMhTjj7VFv/nLYcFezWebCay21rIHd+AlVD1WnRqyjGUozLAv3B1L8nDuYP
ZvQrzSd20CKRMvH8q5LQ8KTyFJFTLkgTjIZXAn7qMGQorLefMl2+YyogmHYDLBwN
DwKUUgLc8dzo4sWRIo08KqxMqTq2vK7JDBj6564LwA4vrsJPMbw02R/abvLg5Fwq
dLYCXmW6QvZCkVYyNLJvh4ySlBr//HJ9Qnq92YVlKvtNS3s5AKY+NuJYWztvokqr
`protect END_PROTECTED
