`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tc95fAAVycz9Xl6Plb94P6c30KNdpBuBlLadB2bUL45xhulAdTVYFXiRmWUAQ11r
l9XfgqdLIXw8cpQjoXCtCOQ3XkTKPqLITArt9+pYtgx0Jc5i1ChZ70fuzBYQNsrz
Y6PQjBNOAjeUGtZsWJzRurSD7Sit7oFNsx0cm4PsezPTO972vP6uy2AtgFbFZSFs
Ji4g+RmZiM0pevu78cBJXqp9DkPF7AB07rOWDDPgY1xjWCkz1O/5lsy5xbOJkZLh
xUSMbWALAYVqMrkVfpd1f3yXaYCZnZSMcU1RztEsMRs5Gsn1zOiFkf/pqAX3Djp3
EgBbhW114FB/72ZYid6jhUeoqOQ5cMmGrjF/jwAysxa5z1muV8CUy+6h5XAkjeEV
WpfVo9SSkLiCTEFpzUhgkYKsJ7ff9f00lHaYaw0QwQx0lvPfptCkCnEigi/jKl2D
mWrvtXeWKmvfIIHQWYzaJxLtOxFhMSR204PROJny2FU=
`protect END_PROTECTED
