`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h+QPWlEOYEp5DwkFWW03myEtlGuG+6cFs+do6iIQH8LMRScoVZZP/2khLbWXmIY+
ca9LrAzla6wy01Amw0uWl/zoQV75wZK2koBRhyj83gJzUIKWzOudFDnkrzRu3w+d
O8Xq/BI6uaQteZiRGIZX7w7aLwHES4bNAJLMEnVFrywJgm261SPG54EuuKc1rC2m
2x3IRtMpkI4vBU70cxRl4m2eeDRGzlRB7vRs5MBkBBrcXLjaPqWWiGqAmcgyxdEP
`protect END_PROTECTED
