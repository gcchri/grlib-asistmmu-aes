`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xx+rfQHHmLloEt4Z6HNeLRK5Kc5mBQXJLiwyc5qjDNbTcnlWtRFRUQ75V4tW9b0a
VbQrciiC+PB4BJ0Iej1/qwibSvpbuJ6C67VpNxJsa9Y0MYQqWRlo3aIcBVy4bHLX
FtYX/2xCBCAzfCM/hUwmzrBcK//Q8VhtMdXMPG62rfBHVouwH+z4hdTkJ2jV2jC5
BfgO5yYJ04YXUN+NptqUR6B9f6ipzSSGDHB0xFs82UNY2FbTYCSvPAWKP5Wnmp3a
j0FgyZtuVWXxQ7g3RM2NWTsmxiu5IIM2yYuDXafusEHBrQfSd1C/RbU6MOCc0dva
qb5QF9D1Z8hIiUK3GuDUykfFLpupn8hcORJm1eG9Ya1Y1s3p/noVxQClTtOpRWI1
slDzDXq6MAP/92gafVrhJEdDNlbOBNeAc5e5oeKEQTx3VYGi2EiVVejkjg/XMW7d
4ZJBHQS7Mrv/p45zX86M5w0l1vKgdcNcNTRiU9JQRUBMqMQyyL86UrXeNnP4KU+I
Jx3953BOQyqQ/QomQHedHZeZx/mnQoFEyCeBKCkqmICGdZHzBkrMnrroOHvXjEtS
XlrBvJwcQ0MVKyxSa2qCR3o1O7iFQ9LQQ+GZHNzFBtawSkIXFWQpML2fZXA4dmlb
hWmh3M1leuF/RLAf4WkQIP7ewwBiCKNmefzf/2xO9QEcIsmrsjutwj6VG/s7kvJL
9JJAW1Gp5CcjWjmedGL6q0BsFNBZgolPINvuxLlYQ22eR82m1XK22ivRV9NwXkQD
DRbXwHznw/5PS8ShIKpUwbIO1UJOaEH51dfmup1Vf775/a/ZDEw+nyg1LZEPQYKG
tJBnVvz1yL4NrGRsat9h/ADRaG7KqvSpDqIsYGEDe1AAE9F13lz5vYqjrQTuBmBW
A+4GKWPn4yOkNOv51KvHwHrI0WLE+lLT9kPy/+DXWBnL04B1Ldxug+Ldgk3UE9pn
dSBtXQiXjysKu/EqxRT/rLOf6eHSnjIt+kP5pbzb7KmdJ4Z2EWNis14gJ2dLOpxU
JYAtAN2NJMNWBXDrnjPlsdQEbpcMNcG15SbQltLY8cTPYzphBtHsrrmqgorxVGo+
G2+8buWh0zukAbVrYbh9LgPObWNTuiIg5vx2tprnOOfjonODjf0Y7SqkVBMFHG5n
l4vrMVH3N0bAIM5XVigixktMxWKFL5jjNcm3D1lzYFPsx6Zo1aosYQlTWmN/PteP
AFWUQ/Jp9c1/pdld1kwMOqJri8L+GqPiC7JfdJHUqR+D+JKBkoAZI1F1f1yN8+Yw
wnoorswaEX/UcIE+YPcys3+BRVwYeRC9w6lzM4DC2SyVnvhIBBhX4b45CMBb+fxZ
/REs4a7rl5lT9RLhSfODeRMqvCNMkrzd4DN84mUPCHB0BYy8S1i8D34jeky+fBgE
r3lS7Bdyf6m2k2Ks3De1Rw0DOpq+qyBCrYOMisOKIEinUOUaPol800vL/0jRRBHF
n58JCHaJMXTZLS3kT40WOsZEplgFWBIQiK61Xh6JMaGcmC1lQVxnaSNBik/GRU0a
iuHBPGKgVnyOaeFT+Jbk8eYhQIvrTfRzFvogo7LyG+ssu47mGydhCVQI7/2L21dI
SS9rPoGWMfINfgIjCXgSjLBectCHUw7iUb8LKOESeeYAhkM4KYNw/oLaV3zDdVIm
AkHeICcQKhOGDbv66PSdkkfaRARO/uP64x1rrKO30NmRP3bsa12fH5Gz9oC+f/Xn
LMWCoURj1PFQ9zzLmUZiN5cacGqlOBlup7gDAkX/auS/zFDt93JDgOVWSebACvai
yEXGKeI9aYLFzrz6xkSlz6KRfOsb+KI5W1DHI8hOAd8doUR+i4dCp68qQeYY+d04
TtZj1svF8WLo7YO9PHFqAViNgis02Fq6DYEGz1mNqiCqghWB6WcvnAqB0YhVWz/Q
ALUVe7RD7feMp5S7yy/NY8I98RcR1M6XFd8u2dyK2qaWX3ux3bOyXzOT3CaBHy3Q
dVI5Lm6wufPhkIJhdiP6EqylHLHRRNOqYLXi4mVHhnL63PLN1hkfI24K/3L7a26l
kw9ZwyYXa2QYzQucazsUUjSH2C9R+v0qfScOiBcTjR4vURmxeGRC1bmehG8Q4j6j
KfLhoEJeaxYcT6hsdW0HZK6ARHR0RgbZSmkrs6gWD+I5k6F1N+bciu27yyJVmajv
jjYVDhptIUMJT0Z4pGnfecNWwSQaWm0QopOgqxrlqt35+aXCqovMMOXERCS90VSW
UdI7M1YSoopomC7v88nAztsxddrJsuBOz4oJuazUdtlnNKM3T+M+V1GC/eZ9qILW
9kcGrnMMDQ98R8WxePsr6AtKD4AgdZ8QHea8J8S5Z6GhqjwXKuK7k8gWxTps2+lM
V2OfCa0cDSkDWL/1RctiCdvSzOHyI0azz2MCdwPzGXQ0hUbKjmoUEu5JWlJs3L9N
3EcRBzlZF5OtqapsxAUrd991QWheUseF2CWS+b0D3WA26NXpG7+V9nXpKqXC6t37
a6iRnOY5t6h2jg8W6iwW2kR3YX3kvZe1Q70pHFc/fkQ2eRgWjloedPYv8vKvsCdx
pLyT4qHzDhqhhQgSZbtt6oJwIJE86UWV8Du0KhqeSO4dYh3DhoncnKb9c57L894M
Z8PKbhf8rliSJWU4G7db8oDLL8ERXPPwN6bGgRW0DIw=
`protect END_PROTECTED
