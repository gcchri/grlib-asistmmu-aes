`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J0j83z45qedfU8DrLZ0i4EPPEv8p4dkiYaDa8uy3wf0jxaI3CFupUNkasBJn4Xcv
vnuY6B6vFeZRg9n/QjeCy26sQW0wsLGGcpUlDNbBSLBIX9QCQtFzXLitSKha8Ye/
7PrWeHwq/gkj4ZofkLpMJa+RqduYlDBqf9Ijie7tsDBLspqKUylk+5l6cf80GZbv
5RZlz7wC3MrWYXQbWqLTil7XF8yMp4L135HdfJKzE5g30MEcXav92FG7z/nm4UWl
7cWjEnLoTmY36OyWLBid6T8nru+gCj4E07iQXEylvBKjpbkJ1gMl9vcHR5w+0p9M
zRLcRKQTQFgNeWIf2q3cHygqAX6K/CSvruuXoHpK1RHFmOwZ8JDnk8/j0XOrGSK+
`protect END_PROTECTED
