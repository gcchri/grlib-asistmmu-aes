`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PGSXydjNVxUG/wJ/0DScoiBwp9zNV/wil/TMmCF83osHat1V6X6mYGG0aVYUAoJJ
4xpB7yxzlssQUUoHXxlmYmqpluLYNn+nh9xJYmpOdlaw4dh4uWfZg1gavEVOx3ED
GBVHA4rI7Q6YH4pcWLpaxXLzHG++M6mNS40ZjX7dxTJsfIp/uudgwPrNUPwdWdzD
ARzjZiEJ9g+z1oY/xHKnuUbq//MDKLDJQ/Pp8ANcc2SCcN/xdNoDT1aOYuglYYA1
3D6gWuf6BTcKXkAC+N359g==
`protect END_PROTECTED
