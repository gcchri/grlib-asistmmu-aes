`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YfgNQNIy4ynwhoalrcB1ehX081MXGvdUs+EEz0mM4rMJFKH4zCG6/4Uhx2Y9Mv/r
8GrISXCqVXemZkGGJiBo6DbZbL3WCMeHUKm0FmXCm30NfLXo1p9bNO7qenrrd4i+
xZrgb4LJTWAJOJSSuHfFeoAN5BGbpi31BVFUvYZ9RC4Q5PNJVmcEL2eZz0ncsMMe
MeAO17cxQNQiLv60zVx4cT2MHOzaJ80JbTa77HEJgZ5DAKDbS0JE9R3eBg045F8z
zLjoNpDdzUbEn/zEP+zv5pXDmsCXo3VmeAVf6K6DQPKjZsdYZav1XSrkZ0QSWstr
`protect END_PROTECTED
