`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
efSSLd3xAB5/yb6vdWKcx5TubB3HifytcZuHDJUdLthLxGhQMHWlLuw1yJfAdUxc
madURz432J6jl0oOKZ81cBjVJL2xc40Ey8jMbNQGf0Jx/RKIRH6w2JWwJVHIXeuK
Z2xuw0xXbMFcBhivpZK9E1kj2dheGlKEPkjRAZSKACSej9H003WsaddrRayhsvD1
OAFOil5csWdEw/YEg/tu5ezQQjf6XLHT/bT9Ft7RxlNWZxiVaCBf0cpp4nxoYWWg
/uoz03iTqiUnADg9NIJ84w==
`protect END_PROTECTED
