`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
urkjiVnzOXIzZ9194x7srEkfq9OGlT8YKE+/BU5FuBkHjJLsbEK5qTWjM7jYCtw8
Vo2l3F91sMjuzQ4XJTRlk3YJnJWglwlYCHH2PGzoAtEBHUiQU8jaKxCgMch/lrOF
MHO8gmQ1TXrAV8C1zD5m2FePqj7hRd13vtMQaCdKjC02ARoy1UNKvRUkJMCp8v+r
/TseLFN1VKfuTPaTeEeLcHTVTavZJxNulwFOWqThE6DNKzlX6r5DiBwfqN+p8Rza
AC5b71GEDZEOOD+OJ9E8OnR7xSQK7v45KgQLgZkiQ8acQow79uhqlNRbbJvB+SeZ
X0ZtXCXVpKIEiodrgfP+jV3zqJQVHARbRBBiBpmmk8klO83bkIT4a6fbefTyc0nc
QtLvFSVyKLi+YRC1Q/c0AM7kLjlnC4s3WQkLJJBWoswJj8BvPDLRlLhPGGrFufBG
NZygVbRWJ1cciIc6I4Ie0/gXXqR8JyBKsKFiw8UVhvhZb8ZNyQYkrgAzyn9loy7x
2cNeppNPfpI3P9aUDQqFkvuDfETZkgbakZXkoitOglrC0J9n1Le208aZCKnUFFkK
mTmE8cutAB8kQ2IGVNYgLdcsmTeB8KZ2RS7ainwZ+1t4A6GYXjfr+iXaZh2G8cW7
Y14+9ftCTsKRUkoM471QXw==
`protect END_PROTECTED
