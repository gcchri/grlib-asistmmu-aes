`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7iPnFZpVvJFuWzC5Fi025hoyYZAv/RirZ7Dhhu72gNQXWmIvUbbvK4U47W8djAVt
B3kOWdwIzShbW4no2BdZbMgeacQfUapjyOhdw66yAMlXmIsSjVphpmtPxERPFT+f
RBmOlLZcjVzMlOlTQKoeXIkuk7MtbogSLJyZSVaBZVk9lEy5Y3g5/QpVbIY1xwKn
W0Th0vbOx1Zsb4pftSiXzySaw76c03qpJ01lqe5QxwUlRBnBFW1IG1YW5jkNnrjM
629oIofqmBQ4iH2c+l6gfdUPGT67IYJqtAnuN4Uz7tAI0w/ps375lKemDPXAH1Oo
`protect END_PROTECTED
