`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rh53888LafW3Dt88Z0yoq1mBEHnJVnOlfj/YrHMollN6AXd34ebxhWBqaRXwnnET
knMYJ9gbAhS7rl1TQwDMq7uboxfumx7IZOWQZFK0jtBBgi7311lFkK72K3sSFiVy
N+Bg2TU3m0LQDTW6tKk/2rtvI74Qs5GuoAQICVvzFO1OQ0QVbn2KCv1EmJMdGVPq
w9h5R7fL4Ht+WSpYTrW2xpqLGgtf6pzhDQMZwy3hdySPk8zAIbB0/jwWFisgK+s+
aDOJUE4HGdAPd7QiqYIuFZSIBxJIBawjYvgEKuvGiovmkrG5goL9kDRjsXYUy4ax
3AKjd4RHm7viJhdrBOBgbk5W6TY/kCIZA70AK8c0VYj1Lb8ZYRPRs5z0qc7dWDZp
BOsZk+Edo6yvsPn526Z/Nk1rIxZmNe8nL6/cxtSMudj9+TWgzbI/O9VFlhGMo3Od
VqkQy/vyb43mz8erGeZiR/iYmwImbYoLMy+DDA6VOs9PVVtn3Vt+90h9nqDBtFLx
C3VaTJpU+nPfOOiDKiEkHq+jAv6wCvW0b5bje0QglkalUo2deHBtn4PLam5MG8fd
aMbM5u+fjIF397FeRf7Xfbhe+xEBBAVYJSXZVNI4x+/ifiwEfr+IYOqUyIjC/QFW
v0aIJPkln2rwtgerJd6DxG5LU9SmpWWAEXsLJGKa7AxEWqhKGjDlJtkuMLsVeZ3K
aexi3Ha2PHne4XpMrbo1K+L3u9hhJzw0cXoskEGH7SfTU+Amta1yHrGn5xKKe5tk
z1cAe1G0oM3cXeTYlyA3kHMTIWBfcLq37PO1ssThW1w+PhCJRsRurG3j9bCoZBlZ
B+UHOLTUBqx1vcgTW04KEd/JtJw4swNNslxu+0E7kbrm9vVYKwBxlhDjVYaXaq6x
ikTHD/dibHT0kdKL+y4Z/e1ybcvAdgTsVeVaCZgYKfltQ2/Wxa0mnbmhXgfOYgVt
VuI2S7DthYZ1XnyzmgmUqK1y3aerpgW0/1WJHKAcF8HjkMGPin6OxmqoaStY0yWy
3mLmCOdi4rcDOjb2nvez0s2S2mN1iMVj0/rW5YQSTwhYzUgn1vtAa9cKw5++cf8z
3lCTpXu7wstt/ys9fP0mADw9UOVE7in8JwALmdkuSnWQUJWCnTr0CHWBc1XzaT69
ShrhBHiOdMnZKn6rUtqXbKomuLqNG0GkKwrvmpay9EMdxnfzAFHfWTu3kbQDwega
XauBDQpoTsvHh4X+HPAGpgH0GMTl09I8AwgLpV3FuwZeJuMxOBFEpYSbuhblkGVv
AowMhmkrTKDuIm+s+IgQMvIOny26T3MAXJlD0T7pcKMjTx2CJZ9nX7xFVV7JluQ0
0GYnvGH0Iz8dZgu2+dACpb0uDRnDCVWy7gsrEUBOHjhajvjHgGNq4DO3ZPFKFrrG
pCHonk7XakQLwa+9y1+cmA==
`protect END_PROTECTED
