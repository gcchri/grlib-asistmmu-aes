`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L6VwJw/9/xaUi4F31xTBnigkWLEnG2QHyu6QFMz+Pb9sLOSAQP79PpMDvjGa33gG
FzMitmZay/82fmtuqHeXfivoV85lmBLgNmbMFCoFB5li26u3MddtzF6nz9i1Zd/b
Z6YOnC9W2oPnznLmR7dF32WwZnCE+qi6yvlNiW+iAGLQpLiByYydTptW9uzlMbUw
73nhWMkmHf0W3KObj7bT0410I5eJJglid8qUTaISeMOstjqK8Vckrqje/+jx3KaC
eCbvnQpE58DwMEkQSwREtmv6+gADYe+iSkBzeetl5fMEtyInKMuPhnLQz3V4z1SW
23ZGqBjOSP/tkfgmc/S+wxK0q81TqAhbuY0qu8qB4ubG2jGs3jZ5SnS9QPjaDVzs
`protect END_PROTECTED
