`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
awVOXYn1KVn+vUr41JtQqKNLrz3hk6pO37k+YCa1EU1iaLdRxViLjpPmVi8k/P4u
qs7r1+ul/mRdTD2f3RFvpj67YOD0vhTUiNtx9JBqW3+MHg0I59ivoFs68KXs+Igy
07cGklEZ2aoyag6WAPX1gtwvVHfa43J6lypu07dDvLlZfxrmgZ/57H/G1epwZkW6
ZeErkgxbUv7pbpnQOEk63D2k54rSSUpp+soIsmvs38m17XqmBpBmMZ2upt5WmKhY
DOF0JhVoyNrsyuO4kxBaQ4IVPwHcoU+1VDGW/pY5XtNhEzeBT/qSa6Sre6iZGcTS
oHK8FY3NkDQEsmtHOgcrs6WwZzVTfMoo85WaC7Ip0YAogre3hZgsiScTAskZO1Q5
igzm0h2oYRnV3NikDdZuhF1JBOplolmAfCdRWbTfEZhSmdL9v1lUUzUxj+e9zLwn
9GKClmPbFl/U0waN5yII/rGU/W0kgGUOWTr8LboiVtiJwp76EyeP64mycsTtksLb
fpnuleAcwGpI5T/6FUdhNUhelmfN91xhAagrTdDBuRby34c/4B1bP9kSne8TbBzn
7QOXeHe7YBqlH+FcURyWKFieEo6st0qWZvn40g+9wSwTDrm2WnFvAC7cDxJwpWkY
dc1Otdgxf1bSmYnqXlSv6CTWbtXvo6osGIiXIWpP4xjP4i16Q4TZjOciAPnIzmLd
4ACrN08iEBnnfxNps/YymtKTFA0iGcjY+HIiYnBrC/1oQReZe7XdDb/JRUh/tPxg
T1y2YiouhNUaIJtslFkW1vdZ624sj6XrYX7I4XpD+aftZjQnGIa36MjcoOY5ou6M
KFzWA+aawgBn5O57CDILKgYrhy/dgYbZ4XbXfjBoVVnSAw4pSjHSnokzLJiUcJCg
iWfgG22o2EKHY2uxAaRzxpB5qNYWTQul5yUCPOCuf2XTDR/9ZDZNh7o5mSBRyKNk
90w1osCwM9+cWPty2KRqHEQxUOlgCAiAvs17Hc3dUuuPvWXsPMgtjJuzKrqO/AIJ
LiJX1p/sUInm+Ul2YOVmvszBx5yaqG2BHEzTVGgTYSHdcwVMJfjORawB6LzRS4lm
306BvMO6uN7/vlk2fEIbmf1Ao+3RZ0FEtv73fp5NY5D/qOxAzN/cIAW7TlDb6VoQ
hWpefwOBTKeV79RRQmMnJj/VP18G6E4M4yfZn2o5pVZ7Y7Q2dUC03EArrhSJbQIH
QcK4b5LQcH/ceYh94Ge+DFdgJq30VdZLM86N0vWBmjI7frt6VzVnOIhYjnPolde8
pnND9Xv2Oa7vI8qsHZQpGG8Q4H7qIyg1xKFPqbcvvoXxAYJUznvOXT0YhhfJ1RMT
PKUfNtOaKZjt9CZGraHIgfEdyK9wyFHE3ixfmolWq99Om3XyZrhvZUDBaT/L91Bq
DXevU4gMnKH3c6xvp+4E6HvBj1VF8sOO22LyxGG6+Pny2D9EQb8R4S8lmMJwL87r
lO2jfp9CXciVjnMD5wlCfiDjtk7emO6fDfjsCHdgOzLre/TomFBun88HACdFIyAX
tXHU1EGmBvgCXxoIwdjtJ0RBuf3PBHz8Hp6bJepG+2IOtnypPpJr7K/YyzeucDT9
UfPbXdc6lTKmwPKOAsjxhZ4qNkf79m5M6kWCL1MgTzcv6TXVfAjB3CF1bPRWJ6VW
kJ5i9pUrIcpdlU9e8YGOnoaFotf3J+Xh17ZujjAj9FKFYnVsZfwGpIsKRCBqcPuD
FKCNTu23DyUi/Pnqzz6VBqDUpnOpL5qrw4vvitGYsDw8lPZ4keMF/PLtiIhgm1aZ
ydQQkyK6qPWHyrv+vRze7OOXoNV+/rhJCJqJL2yNrtvL2Y91tLIlFGztHlH3rDd3
`protect END_PROTECTED
