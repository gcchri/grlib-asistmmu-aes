`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XCQ87wLrI0BC6dyS2pEYjgSCpFjZnitaMwNlf9eJ6uEYLKf8KroqoKOk/l4ucsZm
2k8i+pkVg89pPnbHfvVwBjEL5Eh3UqRd5C093Rz2r8DEE/dNBi2i3V0eu3riWC5s
goxtynf2MGPaOk2y+yuDg4M4sHpnUrEf2dtMLWTzZG/gjBz5J80XAQNc8Gc2lThb
xFyysXVwN+iOlf8UpBFUkgRQM5FZFg+gmWrzeY5glkL+18WSti4hEUpe8JlLM70c
LtGmYRI+WPiTJK6s8v7rVc4X+d+oHixZT+bIRLMM/ph3U185HDa09zNi5xvgsrI6
DWaWHkVeZwHiIqUsgCaD9AAmg4mgfqiUt7PZ5SXwTbb6aLRBuN740GLttwu6SZI6
MckbpNLx+HP5jcFuDQv0DJ9E0JvE8wsVIN7v90lD8VFlnDKPmhJyI+FLXq7SY+EE
uwUNKfXL2z6iqOx8PAqM+2MZ4tQkxdioHjoLNxL/3HE=
`protect END_PROTECTED
