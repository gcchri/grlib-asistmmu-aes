`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d/APLtvcTeJOH+TpwA5ysPnU3UuWtt9QxuAyM/mrtM5NlQv0W0bf9vUUq0EaiaGd
hPDIlQrLIDNDdOxQ+xLag00zi7fOhDk428z3vjvqIvW7ucHEWLdI+sDFQtgDsLOa
OGvXYhEJZE61DN0IuNf29cHOpsUkt9hGS2lCbVmLLhH4Df+KvZ+IvvZf0mToXDwd
gHXdgDQkyfn/D3FG0WONDAJvdaBsT2YvXh9mY21aat038J88qGYyGvbtK4+jladO
nrrblzf9z6iReffSZsFD9WUig948mhNGvng2VpkO+xQkUJ/bc65zgXC5qJFaM95q
1wnALpql0rj1upFQFBNP9wpopTN0HPr+FKMA+fR34FncPMLXfzqvTWrIMROCDS2e
lGqg2y98tB5/Eiyq2Yz7Cm1tP5NkNxTkZOAtaaWEFPf6DpY8vi5Eq5Oe8fzeTPHg
`protect END_PROTECTED
