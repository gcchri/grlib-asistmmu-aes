`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G8JnI2jX46PYfOPP2Mo8/cgQ5a6cqgYY2/I2yVLY0D88iEq7c+QoWOvQU9Sr3HEb
e4NRMw7FXkqXkd+o8dmsKat23/g9NB6Y5ei3mBWHNS2plSIJ8uaAQsYEnkliFLIh
3d8MxWNZWUk1t/KoeVlRyJm4TnuL3U5gCNLPHLUwZSFtAwRWsDcKx1DyZ2Fe1295
N+bXCv3kh2sjxkQRpTZgfCvs9CkLU2g8y+Y8ldBIytvI97tCVfnTn6miktbrnBD4
i9gXcN53Cl5tPMVN3Lu48EVugjKc1P+GhKCbTZp8gJRjV2pUHFfAixTJh6Btby6H
zk2VD6579zRlMGrZnewqBA==
`protect END_PROTECTED
