`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w2GQ8ZJOP6DtT607AaLTPphWcSHB7KoEt4QcfREDWtmWIm4PlsiLLcmWO6cqZTmJ
MjzVf4c1TEWWPqCR7NTX1oGSI0JleqxbqNoACB6Ru2MmZBccUVzpaLI5yBwcl3mv
Qv/LtJ588Y0/XhM/5dHprDdmqTwDmfJvHMVAeuUdwv1kKmbotEERm9F0eYeSwCBX
tPXNOs7Jr+aJ6Df5ODavIwKYGpgxLX/YWtcfPOmdckbKUKxEb12TaBtQRItwyqWc
w4+vv7L0G8KkFZTyHxu6xU4kVXyGLOac9PX27b/4VKU6CanyVT7vJcsRGlQ64Ws0
z617gTEiOy1Q560ViQkd1FrMAF2KgcnrGLWk1H91R0CCnJQDB0qsnE2lMkG5fwH8
OssaDYYOBxtvXyIEl+LAOwwFT7+s3tr3h72oMYbnSJVT8Z6TvWKDBC1xLgXQOm7L
6id6lZFmiQzH+wFAVoPH9WpeUZpLmJYqzFN1jMPUzI0=
`protect END_PROTECTED
