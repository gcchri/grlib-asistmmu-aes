`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1fMhANIRg2H5IKgDgEeRztNhSbp/XktcjNYMh/f3zuUdE0rZBGJiMBrdUg5D34xW
tthJ9ZXjjgysMhKNGHQd/udsoAgZ2dva37yJjkbaW+Kc46EumoiZ0PEK5h5Z8H6g
xSX6/Qu59xbxQApefnGFQe5yLGocbaxfhUQOxj1t6veWI/UOeYtE+5UpoVaaj5TW
TWEXgsLv7Ij08Yl7sTMT1irdyxD7Y2KQNeK9EwPQCP2YXisO3gzuICqsfNcFlR7x
cfabve4Jsa/cEAZA9sQTvXkyCsZpKsiJBnM5UojbutA=
`protect END_PROTECTED
