`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PldMbZzJWes8vgksuM7Crg7N1nLYsWjVJVt6RPP6G8EYE5DyPFw6bhT1GF5voEaa
yeNJ7uE8J7dF2uDzqpBrZYZk23Wf4va9RpTESkajYl5eSMMOago/9kZsDcAlwypd
LbuT7MhusZ1lr9kV8LCzvY4RFXK0oI1j92ws0Msc/UEUM+RnxpoLXht2tWH/936l
8fqk+syXs3BwlaltGe0NMK6HCyyqPrbiBpOhOZnU4fmDEdriVHJChzsLe7p7oBPw
5T8EIenBd9ARbG5cSmycXjkGlkwNKp14ryAKeTwk6qsniIJOkxes+vY/NRa3UhaV
pJ347qFaQ7DvuaweSgOdsNWT0LgZuDghlB++f3B8qe7Vqjpcc9ZSIchLgilzzQkf
H2dOVBY4dv6OkiRaKzkTpPd1envkyvKEg1534STg217uybOwik24T7ZSvHEcTliI
o/1d2cxF9emV6lj0nvPzbHda5R/8OeBSBuwind1ajl7l4QGNgtt6hMAiYSpTn0ZG
BhL9eyRL64QLuyj6eAeslYTqf+EshLGso85a6m4Fshzj5j6br9XK90n17CLzksBk
`protect END_PROTECTED
