`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pHrXIoJ8WPSYjVErGII18QcpSLCAY3QMEeKAHzGxUcFWiLW8jaFALavCT1221gtz
Odrsvm8HgS72W54/8pm/k3t690tNMz7YtPhB+f7Pyw3xQU8B/4S2TprojgFxz8mH
wAlvNse4QLvixa3scI56o+oFY/WQgqAfX8+vmFecIZOcvyR8wYTMKUuQGXBtMc3y
nD9S4WyDX7mKdEPXe6lE6/XzGnHM1SseAGopRjHgbJ6ptL1e4bgB1ukoceIyQQYx
HqtX2nIcsfqtpw0xRkVJFnPpEZtLYXpzd6UuBKqYKCUIPO4KXIi6+iZY80aSJBAe
Ol9jUFR9tTwhBMqd7RS5tA==
`protect END_PROTECTED
