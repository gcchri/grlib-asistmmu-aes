`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3IspfoX4JVxp2fFeH+8zW2kuRDcUucBfjR3RZSkBIkuYfCFdsl3bWjhleyN5XEs1
GmmUFBZuDh+mmlxz+uRQNwRXU7VwgnN9lyS5hJeZ4DPu4pzj3nEdktT7bOAIxypU
DOMnkvrFSrbhxb1JdV0QIPBpGgtaBqHvJDqF+W1t6fMy5p7pva3bCYc95X/a9Qsy
WiOed1le4IfBDK994X1yen7IjLKyCV4TGbL3ThVvVwafeH8z7L74ScZDJcFcWXib
lcv9m5Efbi/i7GnxQenosC1G8MSx4+CmvbUf/6MmQL8FngyqnFDZ9Ch4q1tOAYNe
xO3eo9XYQoMzt49mBnq0BqEYVSr5L4iUh26lpZb1SprTqEnXyOnw/JwhrjGtLTor
sO5RZRa5xz1lrqPMxCVkYtt4q0NBfwEf/5pZz4ztoflJWpG0rF4MoEAzRjDVsxH4
lUlge47Rf79yWGsehNKB9mEjTs0hBIIPD+DhOz31uvrcQCM0UDLJnDJ+Je9oRFZD
1jpmHOGJqJpW0+r3hJK5VCxGfp4N9HJiSUJD+HKGNiMfuCKjG8wwRo88ZYckfnqc
`protect END_PROTECTED
