`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
giXcAkiUJnIF9DEGTObxwdh1NI50glTMCiCGZ2azIbxAjC5jUqZu8AgBKYWmm9gV
h+KiKcG/WCeRx0ggPW3JAMYowHVKCjAaw2t+lHhWbRAQE9/5nVqD/4IHQxOfg6he
0a28G/217sE1lBA8qK3Q1GcpcOYLR4OU0c5GUguPAeLAlea/IE5IjOl41DsLw9hQ
6PtOa1WvEQ/cT62AoaAfuMrRSuvuW36Nmnl7aFHx8vkxgA2IchTs6AyRhuJMGWAh
duDJrzUE5ZN3hrzEkubNq/2DGMgFXYxAY5/kTYGQpIAWJSklals0SRDbD7MHBGd7
jQebYPSxLFVTBanOIbuaIoMqiKnvzEkPodwnKDgJ3kgHO/wWTrrGt5g4LhvW8iwo
VL5kr7HLssBILoJyu7s+vE54bkP2nsR7jVbw34PljwNwlgTyxxPjPRoLBM6v5fMv
ukaxlBrsIzAanlIbDuNCybutyF9hC0YfCq1H49ciXKU62dXyVqI7AiFpj8zeYslI
le0aPAF8pr432XBEsOIMWpDw/JMdKIMHhuvLBW9hDfx0BHo5UMU9nExeJfc865ab
7gSnOUDrrCuv23Cski+s/+dHLGzv85IiouKemXhJzQs=
`protect END_PROTECTED
