`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AIwDLEO2G+ErUELhEPsDI2eKUEcJBIz16poN01DJ4i7LHuOOi7NgY1JTATuE4PpM
IAit2N+aBiz8wHpFFUGjzkJ95lqYvUPmNbIu8p95uzjrINXfqV+Qedb2euX2gqRj
G5JOFfdNvRhVASWBMGdJbarbKKF7cISbbdM5QwIL+hc9wO7cp2zGucQrSps8v2sb
ChEyJlFTNq5e2VUavU46LsSRDFGU7EfyR9+3ZkcbyCL94i6DUib+V5Cp/KSn7otw
EdHnm/vvMKAwQ0ZB1GQnhkpiaHB+1N/T10Si6dU5dWmGoQMeKO3cQ8pZZizS2Ztv
t8cKVHapbBo2dVRD/XAPNrZTk4wV0vMJUdmBJsIn+jtsmPDnQoUl3jAVe+J9MAC1
pKmkQX4KrTnSUE9opyir+GE8N9TWnzMy/pp+whcZjTWc/Io4gOz9zh6G9xxloAyt
b1cQM6OCKrQyx+dz3PnUPYhNjVDUKQK5VttBv32VXt/kDW/Aqbg3tYbEfG6u0+0C
tTs/rwXnJmdABwf8VbA3nHOa9HgMLlqFdYf8ORShTd/aCULAQEBrUvO2fotTaA+S
vDradSdKVgbXYqQrD4d5tTu1XJ0zU1ojfIaoOp7YkqjH/FSHDIxPrzK6xsvjkvqk
P+FQAI1X5TzjnbMLwGuBVQ==
`protect END_PROTECTED
