`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5AuCdzU7RWv3Gcqq7ryIDFoNEZcJSHhXcF5uTciOOc8YvuP6aMIjWhmGI44hmpyt
VGrETCFwTh5Y5Nx2S5TfbEXeFKMgYSP8TOiMfWiuvsAEwsPbJSGVGIb77Cw6h8Kt
Vbq3Effdf4lqgI4R4F5zH7qhv9CbE+O2xx+gzQ4IRPDNsKYozzqfzWDy+BH+nRE4
ZXtUzrz7Awgo2o6SM4J2MYBA0rXsGnPMFaI5wcdi0VZdbEIhrNzvjUhZVc74S+sC
59mY1VTAZp/fT+sMB3g37PvgJsj6qrtM5lOWjC4D3Ihp3br4wyJJrhcVLxUNzjv4
BmYJ8d4C5FxZH7LcwH5xSeK3kdzZXETUmfj5NVu9dg0Hrto46hR6mX8uK+QILoPb
Nf43Nxc0urXl2iVf82i/wA==
`protect END_PROTECTED
