`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QkYuk5Ftc/p8HcYaXGG8n1mmRyVk6tia9wheKbIYcdIIN7+N5jebzzVDDjcboYVd
c4KhGmS0bCwSj4tY/xu8RBtLItlu32ckeyf7dj38cD/jAVQxDpXzHxosXy6ICQoG
YezI3cRL7dpTkD69LLzjK26uCLCoxWlXhyfloeCAt/nPQqD3FaGaG7NR6qNDpL5s
rkNGEtB+leeNlNq4lQLfu9g5bZykFMt3nRKjF+hhK5Ir6bVupiOmgWHHB8Ocheoj
s1S+axUh907D2rzK8KGqN8SWfmMGmPv6mkEmPh5goSyP+BC+Q7lXXdhqGNSugUJ1
68z5PCljb8GtwhwyZ4bYp73AOMQdjEJ1OPgSPNdsP58=
`protect END_PROTECTED
