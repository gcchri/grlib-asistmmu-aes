`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ap5VfyCniYj7M/0sD/tP04MyacVAV7gJO8q1jU4oGfL2lUL9tGb39EeSgy2qCdqP
wFiQfR3y0kLv3FLuPYNtr8BZ/eC1LIRk/FNc4vl8QnRN7Po50qYKotIdEzNCeigF
lOZ0oqfsSHAbxoBYyVYgoCIYlvWfG99aR3aTVYxPBVif2u/cTEHCHQKEAL1UBeQV
NbMxM/Vgkx6JHyWFjdsKxNM8P/1Pkzd8azKfHgpR/cXegs9Wl0YmEeUVqrn5vEi5
N3KYAOcxfX3Hhsp6F9b75XzFB8agJhiAzKIVhyyldQz/5Y7WfB4C0bSnb86ob1xc
xKlzsX21GuqM18ZcCrKFZJQR3D7ie2qE9NPkmKiZYx+YCed6CAQu8q4dVzzSUHML
ymomUzmTGctPJj7zV308vLgK560Ukp7/YTLFEbFVXDPAqtiQUGVeRm7DRST8Bg9O
ykJKsA18gd1MZWcRayvgdeWkFwWBFwv5yRIJ3lKHujxf+QtKWXwV/KboZkNzENL+
b6+0vS+COHALwGXKv0zkpfc381mDYueRcTmcKIQDFaJe82d2YspWS28z9jiwEe76
wLkPrCsyaS7om/dQV98CGp6y7IymthYfq23vUzFTCLdHs/iSW67zbxUU0HLd7Ju8
LAf5uTjkKdmqVbsEceteImRwLJuJsHmjaj3YRLHJFUdhpvOOs5MAnWUYOdc7FpqD
r250lWB26Jz2jRWs5qrnM/DFWXM45oEQczY30Vm0iNQ9hUk+OrfZAYNKE4q+MdlJ
Qb5abaXmLQb9QsE24IRUeToScpUW0xVgvSPF/LHRYsSle2qw7iNuOFvyEA2yiBa0
b1Vh0eVUzSAOqasTIdHp/5v/EJ2EGh7A354NQwboVZmO2432YPv9tNcI1F+UfdFS
TOCKG+nfIfzklm/Ztl9OEQlpb99UnhdlWByNZUiFAJmEqZvorXO1iHRiGEemIKjw
eZfuNI+btTyxA6c+BHoRv0mWZQR8iD8i/Z4M/sJq9iBO+wpp9+NfqeHvnLBoJKAm
LRVMJpD4tEthJztZnISaZ1H8FSw9C2PLEaLWZQcgOm9JGJWY8F1r6SKetxv8aIM9
V+rlHXj+5bUJUrx1Gk/hamRk17kei7WNI+Sy6xK/UWzXbZLtICZU/HJ7fMe/j3Qz
h7RrRmbiRcyMDNJN3enBpIkpE54mHTL6ph+t5Q4sf1jV1nDjbpZUkMOE7YlKfZrp
fcwp36bC+GctspY03vPCONBF602F6lA5ep8oXFWrOd4SVtQGSgX/mf5Ftv5IAxRL
vI8z9+c9x7O1sX0iT1po5KYejdD2hhuB3v4SaeGnkfxapdGqzsxBBxagOrPwFCVv
XrSLl/+WPV1xSl3v5+uYzUSLKoGtPtzr14ezAh1AS/eYz0DRfIdQfX97jkbsIZig
LDhV4tCi/gDSSZB4yIo8yiYtdkuEKqHPddWn0KC71IegOT7PnXc5PQl9RFCxMjDS
cBN5tfuQkMimdmU5PpYTOiN9pptdtKFaV1Oyloz34+5H7mq0lHSobuJrLKrZ4yBX
Upp4GFmYRjQNYUzRidMBrWlWUgRNZF/dy5GjNCie3UoqZW5sW7f/5KwIvjEzzXJu
Ms70ocp3ZhCb8MdWlhqjDPcCZ3ZLSbpE5I4VTP+3dHTnpuLPM3znG8jvV56a6dL0
0lzrmJnfIXTvWcNCQKFGS2wM+8aFCNKOY2jG7/51+zA5H/gFDiu3M3eWuZQ/J2RM
NsHzBZJhhAwAPpVupw6UAf/AhYJ9Lg8dY4T9zzVW+oi0FwcOCH7B3b3EFoYy+KIx
Y3gLQziiPlX3E1UplwmxEgU7CJ1jhoVsU3Whp1hZkF24ak6Nq7C5X6bYC/x/68Dz
ILMS4mEmvR5cN+TqO252VREHyIcSsWKmy4AstL8FpYE5BjQY2OMOds9ywQM/KF6I
VjRw0vmMcoka5ifUQkqSf7TAEF5MWy8tytPx0snrjpnsdkndCP12Y/39HGnaVChU
eKj2RBFA7LSl2F6W96QvrrofevEP5DukK/R1D8TSlH3+UQQRmzDAJVBMNkSmUMGP
MG11TWhtmQHqFx6m935RTVjG0ithLrSqRW8TzLlRHkmWPubGlXU7kn8Zl1+5EKsY
DUXqf5Dpfyl3lg5YQa1808qevEAIL/Nv6z4nhKUwD+99EBPGE6Mn2jTIm5YKZG9j
hGrMEjC0do4OC0A5Hk1TtYiBm+49Tif6iggwFCKu7Kn62M4SgJPiBnePS7L7kSDm
XFkgZ6mGEwRRLbJlDna5jj9byppD0TTW1/VAPXnpJAKEWuLj8o5wpjVSLPh7g8WN
lA+XjYcqY2e5ArxjgJxSN2GKfImSMyDVAlL77Fkfr5842QGpV6s06DXHh0h5Sf8T
oPwSakqyfSqBA9IdnT6bStkSkURvS+X3sMnIsQwkP5kvmz0Xrb2lyNPHrVLRfwjg
Jqvn222s2qXWTO8vdXVALwC9R/BM08mfEPYubOTt/ca+OEod4FS+QGYhL9TG+QnS
Owdjnki4hkZsJQe2Up/oUQLCHVZ/VabXRVB9tXhyV0iDwepvhEN8hQkOZYA7Qy4A
3e5cBA26jPepge4Avk/JoVtJDiimLfw435d/VUoBw6Nwwuy6S8eF0OqpSLD4hx8U
Xyd8Qe7cCNSsHFgy7arIYtAnv04BXbqlYdmaYclEJ3oCnQkfbPb8nj3wMKJ+ih+O
YJI3/XdX1MWWDG3C4sYE6xXqGdNlaP8HoA2Q0MqrPS8iPLoSE7fRiDU36hmhAhmS
69sQ1w1gJThQVrcuD6SNk2K0dRXAKj3Iqc84hZ1fL77SRAPGwah3PHlcSKC5JVWe
4YcnY8z1UivIk4yRFJbOJ/cjgJmm14VNZW1crzXBwR/TsNU+m6CBin4WO4HR37PM
1Nt98UQmRs1OOdDGeAl8RD0Alj8zNXS7Tw0TD2yVw3QXmU3C7tUyaHAKnoxI1ZFP
qmvY4j2pK6i57TpkSEj2zILiAO8z39lpSNtkTYi7KOjYF/xWeBYiRMtPn2mQ0AT2
ipyNgG5R87+xW5Y1qizeWMnov+Q2keN0Ef/KY+E1ruSoZFXG8D59GV4Veog+m/Yc
7HqwGAlBO0wc3OBcqRNqyNILB48EZI5EgNq0nidVYx/+4OGNJzVEl4/oO/kB7YKX
cOV1BShDSQikTsSqo8SyyP+d6HUaRb4sjxhzfvzEugD/VAXll6kUxiHjW3eU8wZ3
Pi74INmU0ZrpxqGRqP+j/uiV+bJp51oikuKbchYJsEGQVT1sEZ1IG1Wbcx65OIyH
`protect END_PROTECTED
