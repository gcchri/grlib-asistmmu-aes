`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pvpxKvLK1m1pcDCIEuibz0/zP5isUjYdKbTtIW41FL7cvgvXuzYiOs2M0hliN70I
kv3kLmuFtA3X0tzZA5AMthGPTcPLozCXDigwtkALZS0ttJ5JAfCbvFQXpDmLqYYJ
PsobPJk5vDjC1QKHRIHL9p6k137FAVaqD3WD11T0X8DuAYPtMdwaXhaNvO+p0hfK
KeS7pxgE+m4wlPK5g/JiNtpme/cKxqLbmkPlPEsoqvhcpfsU2ifP7IfNAurlX3bt
HY0KgsUB1bw+v6hQwiQWUiHsoW7UT4KV6rignD7yn6A4q4XwtuwgSEAhJxOUhc8G
LwyLLhib6zzYlUZ/GK48u9P/cWZhW15jHJHJwPNL3ItSIMXuJIRrpn+/XXfdeVSQ
X7kfONwonPIosFU8+4Rm9KfF0Dajhnq09R5dNF2CrD8+liBwkFqiwlT1OT5c8K35
2qpfEtu0hugKB9XjL5EJ7BfED/biSAlC+kDd6MGpB8ELJHCCJu+I0PxpRHrt4JKB
`protect END_PROTECTED
