`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lmuaxlYIbeaGV2AR6OL2zq10j9h5ubib3wP25VNk0ia/2UrBO2q3GkA/bE62aUCh
GCaTY4qNt9qZD7dQyeEsf0ichT83B19h9+OmqTBiHBK0m5Fq4zIqvcqwZteX6eZP
0G64bkFu9dsb3MAFKAIKtVhs4UxiVEGC5cmYIVPWd62cVHPDxqHpXpjbVxNR8kph
eLEN5NCucfQQgdOQ4hjL/L8l5KqTm2ig8liFsS6DswHbSwfyY/ucVHP9qtF61127
WsBzEl8nY/B68wYcYUwXORrv67/Db8yj9ebCYtvHEhgbvgg842ue1baAq9KFxDjC
P4ZnE4KEsCVHHa4w/dPjng8h/Sx13q5dk15dqqWqaolPfYPfkQ4qby70NF9MuYQN
Oi4IqpnUl+miS7ZVHVB/rQ0aHDROLj6iDjrxEbohgS51ViMI+zOzc9oLLVBit2VL
GrNfE8ZoSACCy5ewT/juISQ7lTa9I8PMnlQFCbAMKciKt/jt7xRrXckVsS71u9Ud
VJC/t+jMv0fMDnYWI2m6BWNmjnieimaQInV5pkd9TCa4nVMi6WVrEjzEXBrHhJre
oimHD0lGRTBf0OkklyXrv+HAwUJORYJ4/J1xuwZHO7s6fB3Tz8jhV4Ikef8m3PZ3
/ABQ34ezWi6VuXQWiSfOeoH8RdZt50ajEqC9m7gsFiO4n3vI04EzFGMhax8Jtuf8
cvuuyrp5uNu1u22caHG2cVwU1VIbUZPggRx2AAqOxn3gmrg3DhwXOdg/egwB+Xnc
S8Jid4jlaVsI2GVmjKFhXz4aob1L90O3eMMdiKa33Hr+DD8XXF6UOjlPg1nEIInT
7FfJt9vmcFOuLMfj9gKaabS8K357WG4xtM7YD1BD1gqpBVXvCzzHFsyG7LeDFVnJ
s4WbHRkuLUXEmv1VEAtnVb0mJsBDbYScoq7ehJXb8JOcBmMQzCSw0lgD297vEJn+
VcFxlxk+1oP9VCoYNVZfXdue7hGIrH8zoe/optNAOZhHJ4DkQyOJ3IMNPqdcOMjH
3/JjUNUbpaZYPQC6mW1FKA==
`protect END_PROTECTED
