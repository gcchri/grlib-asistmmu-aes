`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MaQjG319R8xRCvzSY/ErQV3tNMyRP89DgGfYJXB5VLXDffqf6udv262Bw58Pou+J
0EjaUGdI0Xvon2sJFoRmnKnVVHpHs5dJ+kxk7q9rHTPEEgBdrIDOnJHluZm7c/Aq
KtK4ugrI9gLj/h7u7LOoRlM0trhnWhM8ouMtffheG1N4K/85B/Y4ablhDCm+BnAx
DG4VeWiMXFlGaNmIottkv7eZnbQ0DeDoTWkA1/dnCY3h1QZowQILkjv6PwpKn8t/
uk7rGuOst09GvcxokSNmjf2llkAkqVHdYpbtU8/wlS+3BbD/glDRcygaOpE0z+fj
gLdkGEqesbbYHd/VmGcvrhaAU56fdTZIpsO4rQvSqUiOotb/E8Pgl3yC+Un+sOVN
FoTvGpeQ8Yss7Vp6qCywdTA09JNYVKsMd/iJL7SE4vUq3+PoSPdWNdS2N3DwMPwa
zdejTXzylrTuk6dHDSJa4UdhCYLLHEuaky0N/PTEJu+dOjNApFojbFggZbadQQe2
FrIhfwQotpAPx77KV8LZ5lonGe/+erwDSR/91pMPZIVisOonW3CaNr1m0y8KIqdf
lns47UZmNO50e1vP4dXhra/LDjGPCluZPkg9OTojtmnU9UcAkp/Eky2zaiG6z7Bo
8PoCTWJeGlw+piRt2DTe9TKAltzyV7Z3X1ClrpX2aHlpqB2U2OyIzzKuFyskqyKI
cMG9Fsyktw9DiAcZS+soks7mQbObYci4+BydP41F8bPEHw1mqwWBjkaOC070HQx/
Gt73YsFjpWlaldbsrkRXcprVkdwZJOu0bG5QVMQ+lzN4NVRbFftTdz5irV9+cYsR
XyTu5xL5LOq5OeDOMpsVT0rRFnaqD3YEI6zYxx5OrWKv7zbI5xyrZut5XPXHRI3Z
K6DQlr38E18MgXw/270RgURWAClm0kM5ENStypZfHsBgfHuYa8uDqoMTx6LDxbCN
Um/4pH1BSTJJOoISxXtj9zMR+UihFkEJdb3WQPECnEwn9RXTthbNKKzZyVerx62c
mrWehAl1823+2smKJLM7gVdu2/Tf9+n4BHxQeawzyXzswfylELGKe9Z5tvj9ynPo
wJ2F9e52EGqmcJG/G7xAMACV87rfV4FynHAa+G3I9CWTlNali6/bet1lw3ehI1qE
Dh9ZUEpyh6kykI+wt0KcOHmilSDuNmjPckbnUY4MRD7WGon4sgeuET0WrHOu+qtK
T/9mIj5l815OCHgUu9bba7LVuk+xReGEHyJnxl3nzpUTuIPYzNlWxreT8pMVs3vg
FYl1UKZAp1czkHSHCsOg3z8e0ckh8HCsSvHGubPLN+vBo5AtFW1YYjjNVJ8ea6/A
OqBp/QMKqNuq6VMu2yJxzKKTnviLhQAzQ34Su6xb4acXE3RgCJLcy0rrCDoMLLf+
6vHi2YfXdaXgO/2TVTJl4NWOpRviuLY0zmYt0OmoxBeHd07wt1CCMgFb67LW55GR
Yd2XhKf8a58DtRJi/RTpQVImTg52UC0yzG8hYa5mp2J7ioafHmHa3hpSOzNrHcBk
jlyQyykx91Oo6hKU+cBb47De9S/xjJXlRA8cWRjEygpmM1baW16uxNVWrYCTo4No
FNpdgNFAOgx2Q3wm8ZM7pSir7RcJ0O3oxhLJDwhkbHFlhyVn3w9EORTorb3tWiLf
H8F0hjtwweDyRXK3VYStPhnAtS9lBFSephvABqLDIqVUcZI5u0RkL8KF5pXu2jD/
Uk8gWM/TOC13GTD6Sl7o8A8PaOwmJ3cK+l3jXo9CTTg3ct0561D4o3pCRNDVNDii
tuwh5whlfNBbyg2uIuleJ8UfTURVTGk1nt4lNQWh3f7MFY9iJezVATSCgGLT2/p0
qb4I8oVJ3jY1KlQW1rWpErnyz64kkkIlFsxzJ5IgJe6cwQv06bj4FH+5nAJTKXCp
dExEHyXVQ6cHDvW2NN7iHk06Dyn/uqDCxtM1BcQCo3oxZYdBzLKWYUoP+QekXRsS
`protect END_PROTECTED
