`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gcpzxD5GwPtRgthKPLtKxVSnL6SOWMtQtRxMkwKUS/0BmuzDYvVcdKx3p7KPr386
I2ECrPh17GB6g7SXC3TOGp7McEp02LvbRupCTDIHr1lPsn2ZMn/8Syfsngk7x7tF
2de5PUpyIw7BOPxSp5i6JarZNUN55nKF135JEPSerWUT9uZc3GYfiYqfMCe+zzgh
ZZOOOdIBSM4eyIADuMj7bsv9wy1WJ2bqtWxCenLR4OeKC8fmw3FfCY/lQF1oVcPl
H26/4bPjzRHOZCvg73lx0xZf5I3hax8nxU948JrdGyKAaisk+etKQosdCdw5fMdR
6dF1OtVT6mFrU64pq2ViAGZmCdG7SELYXHEEaYA1QiQt9u+sK5BcTR74yqGHc3Eq
Aaq9GkFrzt2Gapwa+6qnB2LhRwV06BHwtNFQX1U+N/C1gbR5hajoAJRqROKxKCCs
ko1ptyHq87bpWd0bRPEwaHhTF7AWhFHm/Y1Wg3VMyzg105a3NK8epI1m/kw/dX6N
9s3hdGH1RHR1h0cBwNkk9LdrvzpEdTgDt3fuM0xlVS1wvFwRMT5UHiyVP3LZdPP9
ctI9RE9pWvpG5om8+hJpbkENHk+Osf+O1DJjZwLOwE0=
`protect END_PROTECTED
