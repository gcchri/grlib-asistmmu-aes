`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FPeQI2msJEuM8LmcKH4sJkZVb0XHXryGMQ3x/5mDDnt8mrqks6g22+rML6RhxxSj
REjS5Mhy8Q/JvSJdAwVOoTm7cViu/0PnwcZab2gjIiWLTiRx1IGTn4MMqcJ/JqMW
H55Oh+VHi3CKeTbj3OomJxZn/dZbPT5Er/1P738qYaHf01h8qjX14lITTKWaH0wz
LyLWLBzXVOi67VEH7vRqBspMH1PViYRo+xdVx00XazJ8ZOUepoYraT6oh3tXCqiD
+ZeBC52SLH8k8RwNHZ4bgLZ/uYAmgHnQMF1BAI8RXrHipr+XdFdmYby/1rd3Rq8T
rudPrMqWsVY86MACsZ4fnIrkAvabjLpdRaY+mmyNrVp6+NS8lNo8olJ3hcPA4Isp
YjI/fFly2DnL7qy6kRC8nxDCi1QAZRqIpiXx1gBDW8CPgdULr862Mov8ZS5jPY08
f/bwliLJm1z3LSZZJnS7ZvLG/ZFe7pk7x6Lj2lF7OZ5nSYe3e1tOIcVYk7119LAd
uWctaJgmt/olaVQRk3Ne9WA3kXNFu6PuUXcSZRJFaYRY6Vd2pkxUH6ayGMPkIBy5
`protect END_PROTECTED
