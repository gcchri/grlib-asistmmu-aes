`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oSCTuXKsD7hgFw+/fz6fDr+WRS0O57SpuR1Xwtgo3araxlo+rctIzz4lTxzCR1ef
aZ4n7JA8Z3LsmqfGZPdsTY6hKstGUe06PozdETcwo4kvw5ySOVW5fF4DPwDLVJtw
Rxj6M6uTcyx6udo9+SpaHLrm7mU+61f7MNzYMbN+OeiSeiduloKDLvVLmyY+XJE/
4D4my5AbdxCVRTEBE55ZGGVBsp5BCRBeqneHGSg5L1rUyukn+w6KkIAwz7dXL9qC
ZHzvP1Z0LoIV8sr/s/SVm63lsmxERBK1pCgGf9fsNgQ=
`protect END_PROTECTED
