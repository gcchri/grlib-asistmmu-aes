`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z1k5YiuM8Ck3TmYlbhPqmsIeL4QcO6qdsKJ01gP5Mk34lcjUZOL6ZCgE/fje1hLJ
IZYiWD8FRqWd1DD5VWu7CRAnQ+FfvOvLhtN/to/1ZunUTSxZ4HTrJuC8ziVxvvDQ
G2pvhY3TipzT4uZ/k7zRfAqdWS2lBu5jsCcSVcjR08Wf00vxYgLI1jXnxJmwgWqG
+Mm1HY2kgJdvaABf6LlWl0p/w6t1r7MLrQOZPRFo/ndWaJeYSNLuxl10KC23Z0Tr
hJeViyQqNjGXMGFgg6wzROwsEOW5IaDPQMa+qMgkoe5psqak955f1h10GndoqR52
Z3VvReNTYl5XsTAlfrLug2Wf3Rfbvjna0kV33Nrd8qyN0aZFrOGf3+8P/y2pPtkc
qYkG8k2CUqa3wQ1x7rqSE13c/HEy2vKA6WrGDkf+kzFpycr0ZO5oPeFFG8Vn84n+
rgOn8QEwgNvWrfGJkFucrxrbUQk5sEazNz8PgtM8PrygVmqUNKccmcFPt7KFWZyO
o50oIpqt+Z+a5c9xzA166ZP3oMIKmmhon67ISaUHwamRgqFJvql04weaG9i0na+F
R+8SH4pGUOlM1DOejkb1muVcdjo87dR18oe8WZDw/ZvMeSBWYfrl684pub1jyExA
UYOHkEltg86zrTTg+lzUxJ3lMzulL/vSeJsibd6SO+BZiiRxnr6BRSlDmn8wcbce
`protect END_PROTECTED
