`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rUglG2os53NSPSs038oCnCIo+BvX8MfyDvgbzuWllBHxu+6K1mDUJi/hWlN1s7hZ
vfumO5sEOjtiDwI8weUlGU2SVLVuyPlTUmQVVEH0swDHZg7iN2qHhKrw4wgLoFs7
DhJ8yVZWzYv/86F89cxwJBxQ9G6x3uPAscOsupGoG2M+kbOl1YWxsgpTnxMtslMS
QI5bamzVxt5dTOcVncoPhVSyLmfwkF9hPVQPlgNv7veOZJalhkUSSlnFfCxLoYSf
mIjY5KElIWYV7Ot9lhQkIwn3HTVf4SnWLvBdW/Wqy9r4jrE+JNudJHzxZQiPDmjj
uIt1Nt1JQgXc5vTa+g98lbuqOOyyPLq3E48eOKDSrpy1lfqxI0Tz4Ayv2Oa4xjAy
nSf8TwEve4W1eHMogNhEWK2ZrTjb0PYM628sHkxF6hOJYg0OSpN6M+HhPHiDL197
`protect END_PROTECTED
