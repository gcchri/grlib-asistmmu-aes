`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NbIET1eKkUQOf6eXpA9RCk25VHCSpwpxerwMLcqL32QQM1xR6CHa62h6Z3Ab0Sqk
YeHv0X9BNOCmR01JxtFk3GigSAr3iFXJDZpaIFvWD00Q3kjD8DJKi3QFS8g/sXJP
2/0r3cOtS+UPF9ljAOC8CPdRwk47f4cX9t4dTsfrIq/wjmvPv7WFxd0zqhKQj7LN
h8kyGbF+4658qzeKTqsswnlE2SeuSWEQ0tgI4KngnbjfQcJEaPcyvtSJVwSn28NC
aukC2CxGjBeRnAHKE2sOIblZUk7YdeB22KWIwDGtY7FDX15iDCleOWp5/hrvX8Zz
OsiaaEvYD3ma3onw/jxKM3+oHcc8l+rCK2yqGpAPaeF3zD5lJFdhlteHwh1sesWz
t27FCI9mejiHCEMqDfnc8gQbKb53IgJWuRUEUvc5HkbhqJEQOR4MCRvKentaQUyt
J5/oXxpST4KSVxdQjAAxn/ahORZCgyYTWkI1ylNYrA11mrFX9443CFnZZ6T6u6Ls
`protect END_PROTECTED
