`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3NCZ6kmW4zX1tgvG+3j6pRBjjoDoKW8JlABsOFNz69NnR7FbJRzhgUi8ltTU07H+
/Jlrx9hdcfFRHY9XhK8nRopMfZ4sXeD6/fTZ/4eUjRt3fk8s2cauS2dwTtIY/F3W
rOcHH3BTC8Iqt4kHszA+htPp7NNkUrt1DYY3LIgG6Z2psDAkV4eM9bp6lM1FoF9i
3ZAPJJkMPpgLNAGwpUFds/X6C/Jdpo4CpswntZzmWxh3+zVCPsICF3pOISAea8DP
f+e1GqnD6SiZY1GnOZvCE5qWSfH0atSmkEfnVn41QhjJFpAM46VzA30ujegrjGMy
Unu2YXFBDfHhFlbFmsGTkJxPOswK+Skl/sqRFAy4lavmExl/+O2552GNXwZEaiJG
/Ql8g/gQMcTtAQNuwZmW5oygVMmVpynef1v5F2EsXTx2rv0dgr14trPSuoUSIk6W
`protect END_PROTECTED
