`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5WseMfvpqkl57O5tY/fpr+q8B/bihO6rmijNmvmZ7WUsaaNgWcemYbPe7BLsHp2c
IDG3MQ184ktd226WfuHwbwi74enszlxKQE8nia6GICJ3q2TQGOvDwapO3xjHLUaq
Hhhy0TPbIjO+EGg6CCQjuyak2H9+skwKn5AjqrXDwzhKG8I9gAqzA2pcV0wpYj6F
kCbw7idI2aT+3Bv5ZwUe5zGsTPPsVQ1JqWyKMl9N4WGzslwRrgCTrxAw7kaAzSVo
QTcNlfsyKRgTtuvjsv3YIKFfCYgFwkMTWfo1y33m7Q5x8RjLIWdeg+TfnYwxYEos
`protect END_PROTECTED
