`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eN8ttxRViRgWoO/TWd/9Wlh0pjOeGNe9fS3wDOjcNWdnAwb9GKP8lSNteP5HU/VU
etfQj2hZsx9XCuLYGwV+tZHyf53OesgdpjZGvfeINDPGlkchmK/t90DnVvYFykCH
ok9oRWvhhsoIQnmhiASrx3n3pZbgVvdd583dxZV2yzZgMo1YsU/DVURtaWhFfcCx
9g2ei+6gAvEKYPy1ldm1SVYZ6d0zrwVs+rckIsB6IPItH1JvZ1WecvCes2fTdrGZ
/nqT0aeKt+x6aDTV9NOWmVXREgXo8bGwYcUFpDJA+AGtvWJo2f56UamLFeGurzd2
6BLcYTFxTFPvbLr0l2VDcGcGXFUx3LoTaIwPbp1JkEr2EVSOorPKwjSHVVeUSDmj
T9Jtf7nEljAy1InjmOuhojVWLAbWAVDwgpoFO4BEfx5rCjFfGmaTu1vmoNOmLEDm
Q9JRxngLMo2YUXEKke2RNc+8vvhN08mM5QqcUioPGOArTWlE88INumxheknyWJqm
V9mpvK9OXz9oJNB76kCAyt/PYNKEz3VXP5rRySt1qEkkKsHCBy4ePoMh6iHfr+i8
VwHP0eewMhmAbVRlsNSpAiZbddHhDxjtYuYWtkMSTPomBBluwuEah1LziaWA+VI7
sUdeqZsN5qh3ihsDaAhPYPh20jSBXWVToUkDBuTLqn6BFNpEhboAoYG0QcVRwlpm
SGcfAl7rbCOYpd4rOCmo7nJ097L8/IRPAnf31aGF+A9liRgFP5duu1pcACVzPjX0
infOu0NATsxKInVjttu93BbZbzIuiVs5JmQDrUpxp213v8hS0/6nkCe5ndvZ+DwW
9uuSNrmZuHLtY7BA8gbFF8/4vg5Ok8cTF1fYw16S6gsyi39YZY1jsiR0jyfNUUrJ
lZGvsH00+LeSpUOirJkx58Zpk7hLzaU5mMd6pJbB2Rpyfp/dqMlAnEOfXxmhzcsy
fb6B7H0YkVZL59UaohHST9qFDYMDxzRDqQ4gcXpTazAfMlDiH44wlGFCfo2DX/Nk
3hCsfgHQWphlEEDKWp8qgNVmVFYcrOHW7IZlzqmOebBK0/H7OTeJ8lHF3Puh5qFu
iwzKQ+6d3lVGntQZRh54L1gaKWZpjylOcb6J93l/Gmybc11Nzb1TlUjGUn5QNNYl
ld5bbT8ByjLdy12Hmq3VsrNoV4gIueTtXtLqsu4C049mwK1FIuqDmpbO9FaL3Ky5
xlKTh1n8Yp2ng1TnknJOWPLNjmac911uQ8SNuwXK1O5+zpby71xHxBkE20Rl4KGI
hnhWJdaw9pQFRogb+NaIzUHgUy8EpqMfiwcxyQEnmCl5r14IfHOl3jvxSGRJsZr8
AyYs7gjXozbytS05Ijc6ziQPviI2CjygXDCUdpKgT6MPtPYxQDAbwo6H3+a0hxtG
g2Odm2Ez7X+61UfwMqGCqqalax7lkcHVNe8MS2RwXGytXleU4Prcj7Ls3nNVU5kS
3sjDXMLOIp855SvmR+/Ik/6cJIsGaVs4sTkxcQL1nlgAv1Nhn6SS3ZuhCuKdYYsJ
m7cH4LzTGhkgifoWrxNi5b97mEhFWkyZ4gYko+K7xBf8dplK6AzokUEX4/dPXFSV
4WSTpO19SFs+UzzzMOyGqjQwiA/5YTYgyTa5YgwL+KYxpUO/lVQJ/BrRrWaty6fC
K11TTUJDvC2nzPf3tL+o1jeHodwckW3xnHdz2sAQjxv76uLZAydid0sHAMebcveK
o+Ql419P0V+u6Rt3S1CiE5enXDSLnX2bJbTRSOYjty91PqhjbhXwmMZ7h8XGsHTA
PhhA8PQWztyTLPs47dxb70e7Fd4WxILyOoehXyYjo5m6ORekdBymZ+3xYdASCVWl
mZHYRL70PXGIrz8u6dOC84GdSySsmRtXu7MhoWZ0+ffP3d4SPqhzcc4HZ7x49kzj
71WcBVaXYRUvbV9Dnxqf5ZwI7ea4RCdtHi+5eYaueYof1MEDe2sc02iFOhDKEOeD
Un3TsdbTYQU3DUrKMqmLifK3VJBvDHlAq7Dp/bij1Y2aM1CCeqUL1nZX462UNhvA
lR18WvU5/pfpmTjLtTsyAIlKIKQHu9kKlXiTuNq0MoRKeYqmdsRUSN/ZzdhZAjCq
YCRNZg+BS3m08HDGepojZOqoa3XyxTCrfy1MWXNe/z5H95yZu6O7eBSMdJksKKHM
gnhcOfusrm9VvfjMlQ8oyGuXJtbVlusPazBobwXbvIX9g8n3Qd3TZ0MYAXVlB0Q5
oE/NHFxywa5DI461Kvdp0g==
`protect END_PROTECTED
