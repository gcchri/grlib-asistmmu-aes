`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dxT2iS1X5LBr/Sa0RxcN/idhAqrtga0IfCTGjMrtkrIbSREOtMxCNCwlBClejZbv
cHkDMmpvmec+hqI6u1bn3/OAEHkbxz450Mo1BMO4xXcbRsnENT8mXBC6vIikgBeS
801RpooKtvOTM856S214a58h1efKERB6a4kmkbblgLigMOJCYJgJgmcngwFtOXlr
dkYOwwRl88pUh2Bi6uKGKPtIjtmJ4JyvHqSbn76qGoviMjj3sbhL6ouWCYODjiQu
TNGY2oyUlvhmQlXybYtXY3GYeTJDtJTvpCBT3jlZ9O3xbw64PiL2V68ibWTvUxg1
MLWeXrznmdDzPsZUcUsNDz9izsoxiBGGBUkO0BZDT70S9DL0/EVmD6sXjpQT+ywf
8dO9qVEM/lgji5zx0wz+OaexslTCjaWWpvEZsfrTSjLvUFsYHZzvsfWwxVBdnKGx
XI1NpLQvZh6xCyWDW7QyKQeeKBqaobvlwYR9yE4mKlzLKibJOkhCd59gh7513q4a
2b1x/yBajJCA97gWFL05bTJBd1N1JHxIdBNNatOT0mMrdXEEcs0y1C1YAGRdNcFZ
Li+e7AU+gDyvwCHf2/6YzgApVqBNolnK805Jq4lP3lClIOZguFURIATgWBryATNx
hIgw/K3EfyFyVOa6eKqP/T102He8Gg6xDeD16qIRQ74g3PSaaDgiktKj/sEQS5yy
14NpDriYMH42fdW5RN84z6QV/PQg5EQwmjj+wNcHiTYC07/97CSnA8LBcP4CMhfl
jFooqbqxz4S2/IWf8FdW2h0NOc30eYQ3YO7+HAR1bbvsX2Xk9QaCUorO98J//11V
CZcLhMeh2crgS87ZXBOKuV2BRzV/88JXUpsIQpNpxCS9e0lXrKZwhzZ84U4qUjNZ
hJ6qCbP/pgwrWrExB7DTDJzFqEsUiTusJOk2QIKl7EHgDouR/IMsEwq4jIP3VWJt
lGNt0G4wY3tmkuC9eOBX1xuRCADvst1WBli6pb1h1Z3pLMfo4Bd/Qpu3TFecz+lL
WveLBHUvLHDcsZPQIvsiPdWO8kg1sV4cd72MDXx4yy/BnxTLa27lD6FKfQ5olOgw
q9o3gV7rVcDRtFV5EfIf07c/sCdtud6yDXBOPCLNHd2roJicltV7oDsZ7ddl7N6z
nJIb1l9KGXp89sztJ1Hqd5LWp2TPmM/ybFG4kXnGQCcx5kjo1pggdLglCCyLLVt9
B0mS+0gpbM9ZFsd/rc9KYZTb7HSILdeONgSsDq3EdzmnWogREId7yWAwwoz6HJFw
lsRNxKWSsPbD3pLImj3YQBMbZQjIURofPHkmr5Eitg+j7BHGyptJcmRiQiZU2hhu
Vr3a/hCOayh9Cgq8bPZRZ0NabVROOrgv6FG53e3QeEQuNbWpzcAADoBQbVE7qXL2
T1I0g/mho+ZfqZV5xDbhANvzCuXnJj8jipNQU8Mu7F4SimwHTDgd9/zdxTCCKFJn
R4lnj4VdLPcQShWw0ultzTYAzW7sxskD/NsIqq5FC4C8eXe8wAQiHNr/h0w0IAZV
mCi7pMxWT9aFClqZd8t4/1anvSXdWFmvVv6bbQ6W1yckui23647/5R9a4W9eY1+S
iL9lCdVC+5yJL76COLKzmKYLtYuxmHa1q2/yt/oPGm1PmJodzcTki84h/wMCCXEJ
K3IB9xHdKf5qEzrtQEunKps6mo2iSvy6iTEpDGZ9P+Jovn+b4a+Q/7MJvtVtKeH1
g7XOZQ4p1JiS43NgmAQnJohxphnDhoND4hw2v7LviX97kbBNwUVkztK2myLltpxo
hPfABnJXh0VHDJGGDaEjG+5FOqN0gMOc4hRE49BGlDp9CYCXiSzgtz/BpkX0vFpO
IPgwUGeh4qDVW23YdDaoT76LZQwrexL/TOr1bOZMJgBsams7wj0fstgqP89u9l0z
iaZV5DeB7KMssqm9a4JvYj5QYPA1TPcrQz2FqVqHYC31QSPFOm9vrQFCJdw0KGpm
Cv3Hr9Oc21+RZE42+yWANRVoR02T7+D6s2E50nOr7iCOixocQKRt75Xo5cbhjwYT
6gU79KVG7s0uRrDfQJ3HKM6WGLrGbQLs2ZVK09hVV3GWTD+xsbxUFkoBelxIcQwX
yuRhARevQFzNkVU9+ZsWmw==
`protect END_PROTECTED
