`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9wABkLBGowQGG2jmh7JOqZyeaI8QQ4LSiZKpwT2OT2EWHtrR5R1HXrrCC4B5A3g7
ilGeLDesofGcKnvkVDmqniQZDVnqwgvwg3zZfL/jXBW2PpP9zXMowXSnFJzRfvxy
uFo/8GAxcvyjnIU8iLPD//aRYjWBjbCHsmSSB/wsm5h3v1phwlnsU6cwXOHp45Iv
uudGhe4a4m0tOF2LC7cIJ20rAOZ9UYbMxFL81PDDBDN+G8vpUJvhUStHU/VMvx+d
dI0wdzo0YZiYPvXdiHwq8QgJxHBqmn0cZrleKXmiK/WrWFKtd0eJlty8iSmxG+xr
3k618P+36l1km4ykosJKS3hXHG7hMuyGsRe/RDOazBLq55NJEuc2Yqjp51yhfem7
S9jX8jpUifDU4cLhkIH0mpc0kBDHsNDCpCjqpHyGavxIgRWJ12Y8YcPOD6goEltK
xZGveUavDUxa3cg1loo7NhSDB58VvMcL8D+vFPHo6TSGd98ACB1HDETm2Uwb7KfP
I/xjHj0DBQMXH4kgrPSZz5dwuikFXY7Pf1lPIQPYURf3tGQvsm4Mym2X4DknPEvL
VdFPkAGZvdBHDgojmg9SfFZPUh/1cEvO/OCzxjFf/5xvRRyCvGwZdZkG3SF4lSF4
XhN0esumAvbu53QDOy8fDGpAatB8Q1QUg22MQq/NjSgisN5tIBFW1JvU1VdPLZlO
t+4+BsXlucoWo0ggafmJaeMN+wZDPFuJufisBB0tuyaW9dSTu4GT9yHrDumFOtMI
JT3xVfSDh4d6xpc4JqEs0mFIiYxQAbrlCMv9CmyUCyA=
`protect END_PROTECTED
