`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9NJZPmv3ZAL06ewyKkJthkpGMb6XchbzN3fk8E0u6/S6Hm389sf44BWS1hCbRY/h
OIaEk2fNSbij7yx9OeZKE1vSXr8w29wuDbsLHAOQPpzd2yUUR0/5866JJ6lm4vYF
8aUq/msOKL9gmYHpUfuVE18CLtqhDmfZJbTKtsc9QflHxiQ2MAzt6dyPia41OnC0
/v3GJdDH2AZojiXL8B5EoAkktx4z32ka/C6KVH8Wm+RMo5sTP9iet9+kn6/IlUDA
JEvLl/C0FaI0U2Pu6nHxlIyzlld5nLySX7VgiYTvKO/xjwdPmfws64Rq91/zH0JT
AIPhrOBwcFD5m4IG8weLgPrv3nY4Yb6D2Z1IA81scWP22/1BKyNiLA0N0ksYS+LG
rfFzMWoa2V0rgksBSbJT1E/c1joJjjP4ZnqU8U0uK/ocoij1PeEcM0/Ags4fU6SB
A+smQ4teGjqEUH5cwMigXVHX7Qwa8iGwO3a9omyBCw/cSIzPuQRs7j/0JBYC2veI
XQoqvOMyK3kmmTLqQJwQtT5je8aBLnMSOmqKReBfUO66CAflMMEZ59pPk6Ugwqbm
Ohtu4d+h+pceaCzQ5ywrOG0/a/cGwqlilAPWHoXRJToBMSULew8+GZR9h+nDkeXy
M3gvuUj0L3fWQUOe81+kOkBfCJTyvwg+ukm2GpyfBGnUCA+p6iZj8ay6f8Ei3lI3
O+lmmQNdgMOZ07vNH5oTIK7ZibVPV50emkAp48ks06wevGtNE+4B8yvo/H8cXy95
dVaB9Sk+qVCMeEIYOns7Zn4OG/SBhEjFOmzpfTkQzh3b0OOvy4EhUY4xZgHf6Dvi
9Ep19rHqeHSRSSMt0VxPYHW8EWRsdNxggAy8PjzLl3XWQtSzaGATQWU4MSVRvlAK
1wTUtNTuZrg9MZUhaiScsUB8yPSUq3o8HVUVu6I+mYgtzQ9cgWC16PsLwhUsIoYS
JCql+3N42CbiHe5SpcRG+Q==
`protect END_PROTECTED
