`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mHOKM4Yn1OG8I5fnDxIoJq289Upw08lgZ3z6INSw60aS0YplyHbUt501zPFbfDdq
ZHQRdzQQTZ/Bu2cvB8hPr0pYBC7FDX2h3J2Y2D/YKS1XQ93zKnVw333PHtMP7mca
AJ4ptmSY4cEJl68KbNX8a0flihx0K3zeKGmY9T840AtxHaMWIzSS/2XNPlvkYzdo
oSddmo9x6MoOpD6nUGUHpmWgIio9NXkWnz/7uDmDFLDj+XD/6nIVINVFljcf5ryA
CD6S07SnnD+3icYxPgkdp8/8xSUMshiZn3FMw6zZeOGKyk90ergVSfbMDz/+UdV3
UftF1otK42yTbRWVLD7NPKaezYusnYd3dhV1HhGZjKJTsWbyvyHpdjz7i9PpsY4g
H1F9xSmZT+CMcqYhEztH2Qu1iTSK57bX/48mBObXeWLQ+5aPjV1K8Iv0bPJrolQH
l1mzUviX9202Cx1cqECVOTIvroOREerSBuBJjF1TzRNCGhpZYSEjWXHbqruQ7kxd
AUBbWSq8fIg0skiLbeV1Omn3bhMNqmh2L2t+2IfGykpyx3OJJMD47Edgbr2IAh8k
S4X+SvVs6WzFmPb6Ku3kFhQmHSDaOR8Px40KMtx5uBut8lEYck+m7wIJI9TbUeua
eFfS3tjReLfbf0goBUm4sVJjrLOH6G+zl8ffzArwB1NdgBcaLxVnRDDp+dNZKD6j
X/qbsm7jMWAyOtu+wszRyCtjt+R9n0Ao7ums++2WT5r9kEMW7gZhejjYpT0ppoWd
97APg2WTcd0TYot6Yn9ryIeRnEhazG5anJliZQT83HgbjiFAEpKqlRUo7oPZpbPC
j8XhxL70XnowIzdrQ3AOXtGMbgbhUSg29apfqjclo3d3wW+5ZE3wza/mNgyDx9AY
quoWThLLuB+4p4+0FX6poGPU4Iqk5Z5GQVsRsw1W2aG066hTNR199ngNGeAUvTVj
6+wSF3fE6xMVz7iyLjXqkMO/nZKCAImB2wvwUqBMRY0ERuza4X06JdygPo+YLJqM
oubRaWD7yiEaxyk3G9F2cFSbSHtBMt29yFzOEKjXmH6mhxRnj6BtISecxCmEN4vG
g9EA9pXdr/xVxOJC3F6tYizXtk9BfpSbnW3B/TBcJkH9S5HjrED55gYup450PqDb
Tp0W2YO3nJ4qBqRZsvkyVkZrywS41saCT5YJMP5yFVhTfROZfVDs9C48HLypmCjY
gMrZQQ0RoVDlJ6WBCohVr3O/F8f0nlxwsdEXnPEc3upTjI3z7ADHnA6blXMIuU9/
ZtiCRivlHlE33oWgo3wrIEImBo/nlOTyeG5UFv2K4kEn21ZgKyMggNwtEEi0rm+I
u5tVrIqyaors0ULM78SQjAQToxuOaAYNUd0Du/n8Cu6TpnXQ6boYweotbbKHY1LN
qxav6jdPjW1cSV2mHMzX6739DBMgpiIn/hXXCKHkYRmDfG+Yn26hQDh8dJw1f0S+
xqnWHs4gnQmdyg6rcxQYHJIR7ZaJWhEfdJRugS/xmNQ8Ib7tSodxeLvY64GXnsXX
Ya+YvPlr6lXLUvl1N3VJbVeVEhRwQ0KLc1TXkcpAzbIpzCnxZeuPZNFkE3n+4sRA
BgK68DWLcchpAGaSi+lKlVsIaLDnNTCz/fMDFsBe032/XD6m6QvOsAm93cR1zkSu
plqx0GYWKkcXzBftv/t3Cz60QROmb81+Mvfgi662A5KG+cjGwyn8a4uk44mqLAq8
s88H7frjtywWc+5BRYM3SyFMEISYwHqltJ3G4KKGLbxuwvnuMA6oywh2AOwHEfUE
QxVmAiSMjFoTy+eHdRWmyH92MBr436BI1attK9rTZI4xkaJH1ouLdXLb36u7hFbk
9Cs4U++Rt/GQk4zBNxSoizSgNxySsGCBMzPbZIP21Ptvd7dugDLXjua6CnNpkVD6
Owzah4NeNHbo1NWesW6RpMj5oGM+3163LtSuZoWwMB69IjsdQO0nByUVmzVZUk1h
AjTvBXTf0A7GIkdy8FyQO27IOmTSZV/kOWUq7F8tPQzxeTKTbR1UANwX4nteVssA
RkV/Y7OOWpVHThSTLLETyc5b1qoFEu0vH/66Ip0A2SvMBYoLoKcEBz7xqtX1JJTr
MmH4KOViQEhK1c7/CnZM0ElHBvav6ro+CJDtNxLrXLke1gXiVKtNxUHzKU+WLHQU
W6mpBNFRNUlxq+7Tr/nsQJJ1D5kXjRDJx02eN2UTzv4/MxVmmTTpxqVHyBnIu67U
IS1JkeMMKe7tnGJ85kf3I26z9Q2oiH1UnyoQdRbdKHY3IoAZHe90jGMPB504HtWL
UyhUK3WTmMaueijbJLHhmYbUBtoTcpUikYGf6bM0FXQRbk/5U+mJqqefV+gMbr5H
dH33dyFTKNK9r1zj74FIhk4OQ0kQJMQn6/sQIlh0D/HoHT+WDIzKlqZzQJ2qTvnK
ZYo6dLSlwj0Gl5SjCb95v7LNrgSYRTuhW2mZUxGPa3NDt3BEgoAc+T3prfCBqVdu
RR8hc0Ah/qT/ha2ahcmAQILrGfPgImjmht/zCYRxW5pcoxKBbln8xsbIhnJZYf63
furcA7KxkT+k+JFms7g/4TAb9N422Q+Pl21DggPKg1tpi6octgVXVq4lV3jxyXnN
Oc72gaFSDdC+6mHXzXi/dVgyk03bokxyt50tz1kE3PEjiXsLQIVUio+A8erI9RoB
F3dpLxTwIr59ipyGsZ8K8iCGJw5gvWke9LQaFjqa9l3BogpEvP6jJKdCIQSy59hV
skfSeoPe14iZdPiHDVWHyb7yuRn7k5cuDfssSnwzmA3gmNP13LKLyRROcUTGhpY+
7S8aLC4K7ryASYDoigJygNdnWk7Og7J/FKQVdOe7XyIyZNL7tQus0i7uF4EKBub8
6Gs6DOrInmuc+Km88GZ2TF/HFhcEIM+S2egQgtnhuNIPU2EII+YNS2ddz2Z8tDEB
4zp5ERrndqzOGcBtIQ93MI8GVcbl9clAE7/gUrsEJna3z13zRoFeqfeiAg2eq8xz
YlNJ3b4SzR3OiYNpOAvbzxH32fFACWqOOuGyz+RBuINTfoZbVvKEBD1xv85P1r4l
H8b12GmjkS/paOKanqOrTJCULxxzmtnornNFnpt2mTH+Sr0Iw88MZK9Qd7mS7R0C
J4Alnz8fRQ/NS0wYQLPkhw8bFH0WAlSSWko2AqdEzoiewN+MhHU46Da8SpgdYC4C
SSK6qjvSNfOd27BmoKIZrwUrT0SrWZ4uLzNO9Kyep0CbgHc9TbBYqnLQrXFeRLvl
Z0uO/Epa5Leh+N6VIRU94OfIj78wDfysoegCRgRw7xI9ecsO7pxjrzTH/OkAvLyR
Ua68Jsy8/3ch3QkXAp2nRGvS4hUxEyMtXbo2/MUdmB5u2a33hq4I+/IMQvzQq4il
X/S3hV0sRvd+DSTfPCBlynoHP1iHjSNhgXqv8qPU3x2mtWVo///62ZvrLoZ0kmHh
YCy3Fx/OsFNN2Ou6UtGGrPBpjNmDHaCEji995I+1QaIKxF8mBnRwtBMyM+eW7PMj
E99MoEf1rIQRj9SEcI1NHcYMIOwpssmoIU4FvErU5NrHqj+XbA9tg7blgQgA1M8Q
7h8LbOOXb3nFg5OsUS7miRAkFhMhRyRRVdNj2mE+554Jv7HgWQc4YMj4HYsIXkHd
jkJhBvjOspZeZchJziX0fisQZRkiiR1/WGqeXgSqOZY1SoZp/vshZYsFaa86+k6S
IW0jbE3/1t7Wha9KksuKnzdJdUoSRotOGh+YOqRwxDbD4A7YpCXcXradRFxNC2/D
TNfHEBJLzryYnxB8YxPsS0yz0ruAUQvhTVPGgyRT3MhnRQG2wjbznMVFexa2e2PX
aOcHjuKW68S/YxBxzXaEt0M/BzNdMNo1IXz9EgrH4lsCru5MDTvX8jU9qeYPRjE1
Sdk12J+uSM9sMB0KuOXyHUnoCOEDB3EpaKTeNDTI322mWdllU3Su6OxLkTjT2f3r
jGARhVIh8H76CGvz17L56iCCSbGKvvxe579zvdR8dIIGhjBefovpiUxq3ct48Zc2
5Vjh94ymWudQRaQpsU9Uz/yD9XiH2IF3IbIRQzfs2gAbZ0Bdqh2BMXR/JosxShCK
9tOdRHuf0U/b0kqQAKYfCJ3SdQV9hCW0ebhmUc0QTSJt5IuhsdXDJEQS9dr0tmC7
nKgaAThwiX2Z76y0G5jt4RVf9otkV0gtteZg2ge1kVr6oro62iE3QUznj4dJ7sZH
FtVPgPA3rtap2EZ6kk5XMZobqW0cuoiulzhfUIacAdsb2YfZWJ/633uKGIRN1YGR
iois4rTIK13eE1pMh/btbUgb96T8Of3qhaGoDu/cHgG+uBMtxSVmh+FBWak1pFix
XaIJYu0BZXpQIvw+FudGJEPgy5JbDUyOra9jhYjnYXU+8Kij5D4nXcYA1zMr0QpR
MaK2vw/wAZkbbnhyC9L2FAnhWUcjVlkYL6n2zAhA8n5rUhoP1hqL9h2UWMog528e
AoXp41F4/eKO+OwOAiVz3c7KpSnr7NorpiWu6Rnp/XogOoRHInLdJP8FhEchKfRK
gf10Ykqum9XRzEa+B2A2N/6MIE1OUg6jUdBShxG6/VMDOWNL91wruC6toTnQwbLX
vOb3I+4xQswpaFXCWJtJFLKlkiEkFuG8Kb7mSXEONKxdic9iga9XG8AwoiF3FQJl
u5xHOUjc81nrbWnfkQPDi6rnVya7xqkXDIKG4sUv2ro0wOa4tmyGB1N7HHyOf/yL
IvQoSYbMbHoOK6gV5ytVfWZhcHooi465fi2F5OMK/RDaB4F5E4LR+AkD9iApi4ra
8KqDCYNWbvF+4m/5otWn99f0VsT/iUmEHuEF+KZ/2dfE+l+u6wq2+X/k72I5omCu
jzYn1QmtJJiJhrzwoDfobRefQzxNQRXi/mnOtHA/7jv+EEHW6EklN73G2dVnKITF
+kkjtzPRRLGecwW089XGuFqfwwzX+IVqbF0J9pElhrgbnyUQePBR6bIc43ypeWQN
fXBKBq7p1/k/jc9C2WLZfXCxyypez4/2dVvSpi+LNuaj8EvrB34VbfzZHm46VSkf
NGIxnP88Vq8Xnf//cvWgao40axyTxfYkqmfLq14OlUZ4WYRprhDFjQtuZ5yCOkKd
7hWwlHd8htEHcQO1ORfqPnIs18n6n+ad1VOrJbmVqwHhg6kuVFQmgWUnCrhhCsEK
Y1NMyXCouAUZTz2eHwziNeJ+kN6umZPPFYp4qHKei9t0iAfLDpBGmeMmgu43ofFB
1httEA2PfKV45LtHAOY5LiOlTb2q6mqm1OfLvV3wQdfmfjEj9SKNVITH7UfknSOU
gxJWCzTFws1aIlSwdyF0MFSyT6CVGACzmL+tiKvSeetIAZZG4YuptRHMkDUWy0iK
NSxu2rzU0cv/9A28h5P2rYVIXCmsmwcLQQu6xknkuCoxkP3yKb1ncBGUiPF1PNKL
ZF3HExhSR/L6TftiPsVOe9D11/fp0MaptUZKt09kEZMZCpfvQLQsqNQCvOIS/AMe
jvahKTS80e8s7ffPobheoPwmzZ2d1IfuWZC+xUaPJPfL/CbbNcfxBF9scA85Dniv
tj4wQFVpUvCW1QXMPVHF0dY7mC0xtl8MbIB2s/u/q66JTCJim3RJpJIJQl7qoX1P
p07TkaAGto2FoKjNjpGF0CArjffjddZF4JjOvPqtuQDSrNhghATKz5gQWbSbMBiE
e2QiP4hCEHlV4fOisTzmpomoEDwHyh2I2hxQ8PHsxXqKGER6qoJ57t11vt5Xb8A8
dH1HNKXDuWWVXtR6vpBdvT0Hao/Y6TY9QBQc1Xyl17CpRgOGwM5rpi/T4Y2qctnR
OgDNWW4koLsrLc6ZxMrGLg9K1BtPMqtxrHodVoPl7Tkpq8rikGG/kkc2Qq4Zgp+i
99QanGjhNVWcwfHRQgNheFVoCKGxUq0ZM53ZwwhJpjjsHW3bFEBxdz9TtrJ9yduK
BpQwjUghM1VbVMCEHLeTk6AYofexLYI1lzhyW1nnwCER/R1qLEtRWF9cX5UtCf89
boygEphpQZXW2PaDFcIOowo1f7JVIJUpnISLFJVLWETGCG+bMj6pW2UHudWB+5tr
Y0ksgfu7z4FLwds3XAe1u8SwshvhjA1qglEssk5CjuqaFxIunGbL3VquIiXjVGig
K69Yt4uqQp+tT8LrtoYYxDzqE2EbGRjwYI2F5on6B1azxpWE/yMgcDWfNsdohzp2
hoajCb9pSlQwZ5j68phFyMwz5OsVHRHRJ0LVY7LodOdmQ2vgY3BX4zv1jtKG550+
r/qYsOyG7X+/ts6eZcioIhCrSa23vAETGHhFUgDQn4iEKmc/7+KYYutQf9TA55vS
+VXGG5TfxZpeWPlQngyY9Z8PHs9UqgVVDaude8lEnl95T3mQCbe5pC0svJWrof6n
xM51LAD+WH0bqX+dzzEOcLK22OIdwV77Apoan8hZG3xlN4uW4zZDnvVnunTUvtbo
JGoKpHG+SzgVyNZ/Qzr13Zj+gde8RPiL+tIaCCk3Mo95HmJWzQG+2tujjxWnlzUd
ocVZ8edrIM7u+jNbzraswZ071m3+dV5VOxCeGfA/PaXNKULr30EmdF8/1jaIByoz
9W5ZIL59+GPyCRi4g5sfo9sx7RHBPtYS8S3CLYz7w8/AQszfq+3Q+C/Pc4fJbpQc
D2kxJIcBdNiTTPxCpzfjersCQrKuP0dhYHFIAJQWpPerZZn+gtua1vXu5KcrSkCg
kPoqpHxTsOBIoT9gxWxzk5EW5Rn5Fd+57KL6ZCWdBKyx+quxjk5kvnTYl3pbH6Wd
4uHWiEG9QpPBu3h03l267g2hzkYxlJ/gQRBcvewbaekRl0XmhBKq4xzboTGxr8C0
AShuDVdgKR+T6BamqCn1rgLctIEbEzXx7/4A3ji3NrANaioXnZFeB8/CzpLh1u4L
DaRwFGZlkp92EdWDQ5T8VDjNuORJB20P+c3IsAGRHysyAmy5b9YcdyatSI4qCH2+
jaBUcwygGf/qiTzFRtibCyqj9eH4x6ENP/TU18cMv76UL1WLNHC7qHbqyW4JFOhj
mrYWIqNT0Es18waW2LDjBu5VKHN77lyhTuxXkGRWRvv3GNC3L2kxFcFqNQqHb8gJ
+HFT9gtiUvpqUtzWlalxP1c/JuOq2umXythby8dsI0QM/l99SyyP7VDD2/2T6xYM
IKMKaLBMYaajqZvGDNl0aW562JHp5r3gVPvEEQFEXs7LG8Wefm/mfrb6s8xHJay5
/fPvxsE1OOVxCf18WUg5+DoTylaXh6XqmgURpjrr5W+3cRoxb1TnwYUaN+/lY3Sk
ImlYD0mFP7Yj9UOeWp9Xioh78LwQn7bgCnmJTOWfdUIiPTajzsXfLxaUuTXZO33m
N8LC/oQyYATn8GH+w7vblI9OLasUgptFfh0GmY2bUAth8Ro8UrIAiztbu7372GTJ
8irtuXDiwltjiNJMw4heT3bgrpDVu4z9jbnyMdwfHJYD1lqrsIvqW8EutaooYqAR
naC4ZHPuyFpE/0ndf4UlG/g2Va7i1H54CwOS6UL0Ntu2HKDXLOu7lorcpVet2Bn1
k7QdNEHLMUxPew0ZjD00nmAgqH/vbbXzM6pB7EtHDwl4KmeOUMQ1IM8uCu5JR1rl
NpJuHb7KdvcN21Jet59CuIi5suZ0HdKuUBYzI7Foh/Vaynj7fOpgX9LBtcDnHd5h
g/SFrtOkqVzicm1I/4vrMezx9HKrSKbaOPEo5yNq4OiMaKnqJ/P9zFnBUwClGSY0
rrvlQ+qZyJFZLFQcI31SWfNcWBck9ctLHSqmkbsJAEcZ3Srzwv1yKmmQT0EMe/H7
pRJaW4jb5xscqTnoUIx0CJN4cIAeMgBHCLImkMv9p/UajMRePCw/jacmGDO9P50S
Mp2iI3flezw/WrizJs5w9vFHgVO0FGDL68L0YT4Ga1M3VRzA9HryeabxjFir4QCE
v7WCUKb95U8nFx9XGc+KwHKGuJDhYUFlDczw+nyNBS5S/lQeDRPw0QucwmfAIWyy
6FE09Xh5xwlEclJLTSLxHO/OU8qDXEPG4rgRmNxRL+B6td+H+10KopgFqaHISAz4
c/qcGaA3/z1dbQFUid8+ECU3rdRR94CCTpVsS9SZL4GGj6Z7tIc74U7oO60uJZtu
r2uucpcCCmMORT1JbSnXbxudv707s1TjadO0Rrj/9YImompCfBruD0dipis+ry2X
vNsHClCt3de0jEJcUiC8aFyduQL6f2MZdsqlsJm6mRepJ7hxLkN6fg7iKy9NfDDB
srw0h03IaAgvFjBAjTtv3yheqnjav9vmYijp5RzsVgJVFmwkgvQxNtrdWp9Oz3cg
SKz1CxzDVmScIYeInMdd9L/ka6PCG5nRheG1uBQgKP+9erPOPUTM1WcGgZHzO1hD
MA5NGYjOBvuTMD8H5/0+Orq3sIvf38QfMydEOwJw4iCNPwtwmblYpKql2n6zT+0Q
aB6h9B+eveGCcvj6Wko6mOICbR0YQGT5Iush5xxpsb8wAVNl2AGQlQtG41fhQpyf
kvnL+hWxDuMDhtoGqa8VIuD72Tm9waj72AlrnDUblYJzbD8aUP7w9W6rSsu1SeTH
woQdfbCcu7e+2aNtHlXucV6sm8MqleL9hq3sXnCY9A2Pr72oOuR8Beto0B/e9esB
e0npizx3ot1JZuxQ2nFReB7IBwyYluEuV3aoqrQlHfLiX4M1lNr+56FxPrCU7GgM
F3WFCtMcroysCBOH6JaCmZRAqLwGeRHNX2Ka1awcpE5k7+WqPJQu05M0l7hOU4RJ
MNiRQLH6MT7OrkaJPU4o16N+pg/nRl0cHwOBqwXYcoF67Lv/c27MCA/CxoDkLjVX
m9wTYXaGNrYyExSoAvOu9/m9y/aUEH0Lj00LVTkKXoxcZ12F7MOgDIceNf4wWkTY
2t/fOEGEr5RwW3bMi4d+r3otSvYei/WjKNlgOy3oQ/wmIatDDNQq39VfFJJizvUa
RAZwwL3/dfQSu4N2MUleSYrwaVEbWh2iTm/AYhF/7Rir6j+zLXwxrKzvvWNipWhc
TVI1ODex5ZAo20cBo7JwO5usR0pcTmHc9ZvkXieibrSCds3CcLHufmGIwY82iXTv
5rHk04gQNem7jr8vk8h/qNY+EvdbcqwI0Ymupn6O6QpGrfWOEGvr2Re741QHV/jM
gsjFO1L2dJtPMdqmn80EDv/4wEvfWshAmDcLCWvYPIqxzGmTvJy4MCa0ArBH6fbR
U1F9PuyFZ62cA+vRBJAvPT/HG+ZYhlmViil2b1yANFvHaHfiRERJBbtqsIX9BKIO
mUJM0ooSX7bzNrUH3V4Z2GZkOXmXw52CMlA71DGs9CeVj89pnSVj6EeGCL/D2fId
wPwxhtPlySbBN4lp/ZBqYVSpaQyV524pbq6GkTctpTlp3zPT1Dy9Cb93NUExR966
dGfQTi22MimUrt/4N+AUO6L2BIRBbziwb6/c7EfAxOZtlA6/ztPa5v9Z/tjbbm+t
zcsRJ3gi7o71prLJRzfN6jqcItCU/kMt2rSYs9O4M+cn9rBHBO7Far+5qAxK7UmN
x3HhcQtFh2NWGQUSpvIUEyrg9ETQcH6PHqkDO9VPdCVQ8j0toG3Z977ECoKk48Q/
PAZPwRP0r+lwivgyqE5SGhjgTF8bzMGeEdz7cJNvMLajbbqGXU3f93JgAs9bDEqu
/y+3+S6r8o+Cf3DNfOAXcQd5JAzVXejUDP0G8htaBxDCOXS9wUzXqYMtbzuw/O2e
E9Q36g+I4+diqsGQvWYDHn7MV4oVrckOXJBs9RY8Up0PtKncR0IZcw4REU6Kijjt
Y2MXybusfYTNP4z+E3qSYe5iLf2hT4SGCaFIRLEPu2HV0Sn6GIK/tABJvahDSvxm
g46IbtsWrgM9Ty+up7JH5XBlnfE4sMDFyApW/uBbyeyuBs2nmb6gOFGwBirMaWMt
9AaF+5W2R2ZpgXyjPKmW+0nE+ObMr1xN3UG0I2uXCeR2u0B8AsPPpnFLGaY0Kzv9
bvZnMGxkbaQwXYfIE53w+xUH8sx9s6Q3mfJaObhfGeaw6M0IJjxUVOnhHTCtr2CV
qeGZMqJgF8W3/Tn0Zc+v6DzEVN5dHfSfKEKQG5pebhq1EJbq7Of7iFSC+sFNpw+L
HTw0WZl34i+CbnXAuG+Dl5YAOCjlrjfvbEP8WVB7SeyHsg9X47np43i2BxZiN23m
GgSym8IYHDH9pQr1FDm3BUWgdd4wfDXOX2bPc7Z15ef26Q4u3FfTJdRiSOMlj4Hl
+6dJXVQqyzZ9fvYt2NaD8hKYsI0/oQ+vvTyr7afnlIVj5sVTRI/NFNgtsB4yVqwa
VDeOqE1aR9A5zasb8DfE5ZcNB8ReCnnQH7fbfqIzTTlc2xTXTFc6p09mbKzYp3ci
OLYiqZsHu2gNoW+6ayvEO3kIgNO2pPqrN5QkgpEM2+ALjkxM6G3qxCyFD+vYUIN0
rtK0rwbpLB2hFVQl14xVFUTCuWW5aPC8V8L2rkD0Jrb9j0Sh/en3HpB1zS374eI0
VZz9Ui38qUzpYJFLar0lE2hNqF5nQSIcl/+uBTIFdwdQRWGtocYLkiui+agPqQ8I
wQAUXUb7EDY6ye9aZCRZaD6kxvZUFJDxobUGE5oWs2z3vgTz60r2sYEcWTePAAAH
2nCx+IzN86YW+D+u/Bei9iBF1rfr0m4Ogsr1ONefSTfoLUBduNEqIumeO0Y0/nzr
7WpclhOTBUgNj09QVFRos/dfjSxcbTnTItQv/4mFyQRCfOHwny9b2qwDP7KRhyiK
qfJvFJ64S7kbikBZol8Wt/c0sLDsnBaNhwHt4NQ7eaDn4Aus3aaohh44BiBzAd/M
ilwbuAqgCFoH08dLfXt1RjmJ9XdK8BAyXMHX/V1CBOlPyqGQ0zBQMApWnAPd9NZW
EFhjHmhhsm5+SXzbqCR2FxtJgDFJyZL1ofrOozQJGzQuh202u8FrOFf+H2X2x7Ls
s3QpSvMkdogEoYwbru2TgYub6GdBuri3vQ+ltNhKPWSNII/XlBz5XUP52LC51iK3
y1FtHqfxKLEj1ZAsb3oAtpeYau/XbcXE6RscXVNGubuo32dcXuUjFxd+4b0N3Q/i
7+b2qvbYeNMwH3A4V/FyTq1/4zcbiLKRn3oaRnsXweohzCypIphQVLsXQLY0iGH8
EycqsuNSUXfvJ3N7FoV2j2PkIog2q/2FZRVziMtwXqOpfRoYkZ68VACc4NwqeBNR
5QesSBP3oanirqTZFa87anxHQjCkH1PJ9jTBHPHcq7p91V3naPyZCfFCmMpW71by
eFmN2jmlruNs77qmOpWCvam4SRFfZp0hW4Eg+mXv6ko0cEWumIVgo+oK2ZyNI9GT
EVDB0oLOID8G56eEiAuTeLbZHeLokqZLVY3uTsrvNyKRpcVKNFjYiOc7UFdaIix3
ZLIC9/VlKV2qaCzM3hQNrdrdqf9sQptNNmVXkru1eL4LZ4gLHiQALLUdhIf7elfM
IHp3LTeWROGBgn5gArwrhv+hT8V2bwqhGNnRFWq/kW2vdpKSFzEhcox28Fv/0ozj
L2j1K/a2kNDuzHgRjHg0qsJFD7FrVgUQabnPRIIsol7w2XOdfvY3Mvqi6GhvROlP
xfoz2/stdHQH+lbp0zmQT6wIf2OwxWYq3DDUCLIM5KhYBk9y2cP2te/LpvYMta4U
x0BN0j17/Ksg5wyRcWGwuT/3tiQQKAxYCOKnUDCoH4IiqQzgOdzepxBtd7L3hT9R
A3y8mMAIaxKAM8C6bkqRLJeQQt5KulG5KKBqKKZ9tNSjVf8PpN96J9VkUf79FdkM
S1q4Vr0u35b+t1zCJ7A+/ZLCpclGMGgewemV7UayY4WeMk9+CVatRSARGVBwV7ni
QBUoooObOIbamjKmrChE9DCwohz7Fk2QEZqhG7+LTS0NTdkG6JqxS0/7plNTRhPp
Qpms3wD+1TJlj6Qf2tWSrGYeq0OtZrEig6Csa0+qluz+B4L7FCDoZPu5+ZZr6pMA
cFNXz2EjaAC5DBrcwlWM+bjupAXM0Hu5Ruwe2M/jS2FjLBZaK7/C2O85nbQuwssq
Zzmk/vVZYUpo/h3EoRBpQMR80SA2QkSTLhU4sOZ19pU3Y7DRdOpDimJyGV8UraCl
QPkqocV2OnMpZqvGPkmbyb/57iBMo7Cq7zVFR5I2zjZ3Yl3n40VwnoYBhdWj6khn
oUSDdJ7zNjcgE58JCAplw2RG0dLZLNgXvuGlSl4YMOyiAF0NOuK3+bup4lcfZps2
uG93/UHfBW+HHLhRl8OsLifOwyeEmi4zb+iEFLgMhTntTfrC7B8PkeyEI6fIcXUs
l+atVGt/zAg9WnfYJ5KrBphLRETURiGBhMG7iHLtSG/WB5Cy+bPC8O06ylO5gORW
dzBoo37VewSaaaU5OiIYi1qSMgSvBjt3jwuIGIgYrqaWf8Qa4C87fR/BdUQMxDIh
P9GQCiTSSN2Y8oMceM/iYEOekFHTkZP28R+kFP2IcsRt5yhCd+J+2cWwF69prqQt
+oxULyF1Z1Ge9OowuBlA08r5XuEoUGqO5NUifYMm2vlplWkqoZ41SUabjc48qAUA
1dKrfNsEhLtHTH3in86btQE7wCCvZ+O/vLe1DrzsRRsH/bFzgyK/Qb+4JZbxwJks
+KMCNDySt3T54darto6LI+3m1V3r+pIc6+w0nqxRgBWsPkTogZGbuC//3g81/a0+
el2i/QqaDNpy0hE//JlaO9Q35YXG+WjgiYsoTaD6mGyPeCMNjSEyvS/WQVHl3dAz
uqbg1ADAfeSE1lg4o8jbVyDv5eLF8bsLEGZFlUlsvc+y8+pYgy/HMCCTuKf7qULE
+6SCabzHKWpNd/vXn0O7wryHs/jP2BbzJbc620qN98Pj7Rh2r/wtFlEh9lM+9VbD
ou0xsvraL9SpizT10xfHImA17f8o8RYENhtQDjDSBCdWNzvH4Ci0DnJikNrFll2s
kvIdmZdMAP8EDomFZHaED0sFXX53mvsLeb1nLajGKLi9rlgRaLHmvV5L7uNIN9Tk
VUFMHyS7W/RtF46VWzl2I+B//yPb6Qf6VIgu4TXwndZ27EPmBDNDvIlo2iPK8Awy
XluEBxOsTRDUqaOrWj+YoxKs0xQnBOzt4uxpscOq19KXQo/H20rw/a6/eMzlcf/W
ZTUOgcSvI7WfzrBr0SauhYEfKj35yv6A280iO4VsBnnZgMpIGDoX1NPU1Q4sBN6b
x3N/QmGWzdc6sQ7XU99aHTqSBGnlz8PLkHUrh24uzAa/YdpIoW38p8xLBtQ+Xg53
rzgMZDvz1IkxHdJw2Mwbq7GnK1+5sLClK0MJfb7JmR6XwREbmBHF9fImwqy/d+Li
0xtsMIcxcHqvX+ndE+4ntTCL6NwDDIQl4OcbSAsMdhbmjzLGjW+fdAafIDcOQp/U
jONgY7PHDYbNd/ZoLFuhBLbo6+6UEQkDlhdQ8noWaidSh7QS1J5860ShYSvzP8TR
Ov1g2PTA7+TgDriia2Fq2rPnSOmOUkMF/gUn3PN2wzyHKwx5VDcQ6Vy7CDASI/Y9
ZOt+yC+cFVcdICsS0Xao1Vkmcd1aj40+PYBuis8xmWdoq/kMMqEfisO9I5Y4nl77
i/dDLpMzpBzWZrpeMU+quiRIFBql/hwALZcWPSr1jByBsI54kerB0eSfj8GRXhus
+7DE5BdOmOnF4v/VCwumQ+6b5tu3JdZVzxjOL/GfbtPOz6nfs4KXHJX69wotMlrg
gtFVKDLx48/WUcxHLgCm6+IDNeY20mHeC43iaijnu9nVMM9e9amzNIXtVAG+3dMw
eKXqYA5ak5E8eYGR8RyP5qhMWYwM6zEwW19R58OWfsCRk8fS2+Wr6RSi7Scgrsd2
t0BtLbcYzzj7UztiBqDNt3iThShkQbmjQyPSExiT2aY5E0loKZaWvVgHdWwha4m2
y9Kyt7sIJWDlCU1TwHLlf1H1R8GTra1HbNg1f6WSf1R+E11YPmCimfVtTpEVuSZ6
Wwvh+B7EsOrjx9pPBVAm4l0qZDbB3RDp/DIyqF8d3ib51GsXaEz0TmCDJUJA/YcZ
8dfklyT5WifSNI50ph986nVrNAbf0Ng/VpxWvnMSEFpcUXQbAzU9pjSWCVh38vcp
D3DX2aTBR5lFi1to7IcRzhTKMsxF24vFQ9DRdERF8J97DefbGs2xWkcoZtB5RGjP
ArF235uGHacUgycuYY7Hudxvk1G86iETHRr775ynd+zKXNO/EQuUot12ITxeDgTM
voHFONgrEQK/FQHd2XNqBn9c+W5zDu/e2YdgtUHL9e3aNADL1V1UpC4P2pgTouyF
pW0xHpn0RFYgolt1gOnNiGPMsz8QYXTmg3ZIIILCwiGWfk43dNAOH2mt+D+wcPdU
6H4nXspyclIMvJKBSUVcqlq531qE5sPJwHdSBcTGIfSzL0heKXSh9QPP1aDVVJMr
AvXm+teO+QP9PSaD2BD1yRbsGW9gUQPLDpmyKceaVvKBhpyo3vmcUqrAsqaXRvdk
6A+xvhTVbwyQYPN+DNKsEkkrtXiKxbdySGLssdqm4CkHLRW+DBI5kop6yvuUpq0V
NaEmXH59etsbkYCSfBLqqpdC2cUC5/4jLGeW7ZvD8A5fIvYBljO49m7+VZt3kw9Y
KZI+QSyf9Lns48C5hnHaVrmMqqau1/pe1PK8cE8YSrPaEXelvXFs0P8pvHZSB9Nj
dmG/ghUjZlJnFQ/EzSm/FV5VfWky0OKx08k++IXzUy4vmOxL+ZLzjX3MjuzASCj0
RuN9KCstc0M9NUnDRnhB9q1dZKpXHh7U4t0oLXa5woMG6wxFMNgm0a4J1Sdf0d+o
XyfvwKpnnXKG1hKmGpyrxn6P1DV+9S1BxPZZB77prxsPoOJcYJB2fBWmUtvR1N+6
0lh/5GTkmLyQvWbjVFZjHA1QCRFzU3Ur9FGxY2nDt4X9lMf2VOOvsxPBCvoFk0WI
zrI5Wx/oBWuPUlu5wvjr1ypE5/MAKIA44cELmV9pqjF8TfmsR9A2O6vrzxqjDTY/
2nwt9d0+RwPUJQlLWJk7JIjvCm+q2wSLJKF2AlUjbmQq7ZMV/sn8rMGYkMf5KXpx
GjabuHo+479duA8fGXEgRmni0WPA02jJLbR7qA/M/WkXZPhd3nPO5QabwfL7h63C
s/ILAzV64gV9FziVFbE9VC0wWZCeHopMNcaLYZt4Y/TjJxyVdMdb33Gb+i4EQQdL
x0xuX35b0ytNct33ec3pqB6uU5ebF4crD2+rhLOC0ifdDfJgeZTBrMvherlzFB5m
iRGeIwkIyOnFv7JXAgMt8C/4IH7NtMIwElcnr30oS3xIPe5/hkY7v1x2reeCNXXb
xoZEnEXSRCocip7d/6daWaOkzgwWUYxPvDJCGMJ9urEFLFViJ624cBIQnKzih/jD
bJX/pN1/wdbufbDCWDyuTprA45N8U1eDDtU9ndMVxpebThQjKlhxis17jlc+WJBF
LritgCq/mvA1/pXJvO1Bkz5Mx60xmG4x4TbAWARYU8o5/B6sfoNjh9xPTIex72ff
t6h3TonL7JqrcQE1QGdHKE18gUT8qOhwnR9NAWTp9JMbU+Str7iVwfUVtLbtvB8P
GhhLm28i426BGh2PoxTIrD72dRgJQMR08EUsTLu5xD+xSws4VOG1htL0LsYNsnvO
6y4uvSaEbahYouV2ESM0M5F/2thT0SdYLjZO0fzmrsWSUFvZT6GZNwtYPAktIqkA
P7AlWQMsKUZ04e2AS9kuXjh+H7wMvQuPncJ8uLpSAQnn/HHSKwPOOXMvh9VfPYal
18cI/zp2NjugZ5fkGMufXpHY2nRUhVwI9efh3jHn/C6l3s+FZutIN+6ZwkLbzUOz
tUsmN4lEMvxY03AyaVlnjrjGs/CC2gBgVc5G9AK2iNqtMIL4lcrkgtQ0I9fx6CsM
CqfA1nT3CB/vLhizhgco4GdaQGuJ5Vy4k1UHCEQ0LQQ8WYtIgqPrIf0lOIJny7hB
5Ol0lJptAaeJZuWC6nf7dSJ432x5qbevu8oBcOmUyctJpghKMN84Qxe198ZRxXgD
U9EHoQc+kPgBKytG7SoigJWFOHn8Iw6IPt8tlKlO1uQPHqodlGtXrjjYEq8yeKRY
3vuHcmxR+uzUdKQeAdW5vUqMhEeW48toXXQHdWc9SayNITOXSzaa+tTOZ8MBSviq
lEVXUcUst1j4NYF1S60TM2a9WHpV7anPEfyRv7w8x4TIldDjOBn0WdfBYbsf7SxZ
056PuhWuyG2zmA5RXai/NtbwFDcp77tukEHP15jRzLDiFSxtXZtYXh0C8fOSk/Fq
7x0FSugVXTVF6lcqD7PboJtLt6PmBPs5je6sRjEbQ+dlk8WO5M20Eq7/SS6YrEXb
/LVdQunmLIGwKbAD8GRjZ6XNVuHr6sFWeWQuVPvWrjNX12/FSXxyyDIry7pWIJxl
96QwKtay4xYF3ruw/a1NXnigmeJqOgwyRYj2P03KUu51GyaZR3mOlszZwvE0tdF9
QGB8l5eXSRMVSVf7L3yZw3+xO5nQz1ab1o+ZXt21cp4IkOShoVeadUV/yqTXlCPN
xsjY98HcAm1MdJ5PMG5JOuT91+mbYrGvF+HCBrNfA82q3ylHavQy0xqPr2Z5f9Go
VsxcuowyjJcmHtAXaFAW5pzSiWJ2WGetENgQNhQHTpfA0/n0xW+vpwB1mJTeOHOt
FoqcDGLUSw3Nh7Q6gbQmsgyWnOVMYAF8FB66rQVT24CzP8d5HrqMw3D9OCWoxgju
CdEpwBSqjAbSAV0MBE2/Nqmb4OcJhg4EocsaJzizBCvfPoAQ4vEszQMmj+khYXk3
Oo0GxeAGcxKpOUlF1XALzdqUSe27L8aAYwcaTA/q6w+jJfqNpn5S7e3lDXGDuCSF
znRu3dv1kqVqFvYGfw90Ksc1ExC69y6n0URDa3ycBWP540IwUKqwzzq9nqD0ujHA
QOu+afDDaTKixMAnm6o2kmw5k9ITgurLgnD62r3VSbCGZ8VScATMiJte2xvJsbhf
sbwVvsPoUF+jEL8pn/YBTPRgx8jj3Nntx8i9DAFgyvRmJWcqbjyN0vWi98y2quhF
tOJDIAZbfNExgAXFFJ5yV3NaJPSNDfVT4WVN9VskafZYZHbmtn5H8x+syBVKO+0f
/DH9pZNMUCL85eSXpr7N8u99Suq+LiyzInyncalxsXe+KmZZvMroJ9pK0HzgDPUz
y+iewy0RmWNbjDAoqhi7lN9L6QyEFuaRDvUDJMsRLHcjj3T/CusATY+O0K8T7POH
9JFXKptpntPr+9Rq2KVybeVXSypRhDMYSH7eKL1i+kojaoNdRuZSut3NjTLONF6r
7Vkpn0k3KwHEY411FrpIyhWFP6E4M+yMA2M6XXCjNBIjz0RlIzboFMWJecOQHlXX
zt4dDmFNlsHVO8Av51Rspk+Ckf6/4Q61oTELItLAt3XKdH/qRrT7dAZ8lqo706gO
mucm3j8DcZiBeWV1WrsCYFp3YsCETLCBKdwionlRpJB2CH5LV0XGigv/CoU0srpa
vjgUHaUweox2zPpgNWKyMsMe8g5+ZvT0Dw7IoUmIaWlXS34mS3JC9VkzQqpa1vG0
PjowMrgrX0aSYrzc8KqPybwFKgQd/4uJ/d8hlvoPgL5lEajvfYEtMKsfqXdP3vAx
TvImWDTfXeihHjz5cN/7lh0bi0XjYGdWm/UA76Vg0qikCSr5dvPukQ3nNiMth3bc
76KC3zkCD4S5xmrHDQhCcR/tVbA1DYG5y476/8SMjDlV+ndalwrjQuU008TFH6wU
nMDrC6InyT0O9rhgAboc5et7fbMuOKIukefCj4GZDOtyZIRR4+QOKjLd0vZXhp4W
VyifDfbgLj1M7aN22P97Mdp1l0bli8auuK90l8UWM+uOX+O9udGtSmun2hocfpbG
WF6ws2fJ0AFt3K1iQxw1+lcgT5F5B0LdPrVwdoqIOz5ytfn2DxU2828Wn+byWKVa
RhYZLGW2pFq9ScYgxxeINv5w+OuVOBD9n8XLw/PvxD6xhi/iLT1nyWdjKAhdRWMp
qnFG4531N5hKXm0/E7Y3vJJwKZ6wXRMGt0ao8qxdlU/h7ndC6/KoxVmqO0z0SV8S
TwrbMsSAPGOkmKDdSnKGau1HNrmP8D4qRHJ+NAqysSzBeg8uDibd+Oodu4xBNoS8
YZ+gKcF32whDLVK6YEsIVLjXKERu/L95ddudfWcF5ppfyPGDlvE1LVLJUgkgKqU3
fQbUU50GhxWXvG0I521sdV45VhjMRXwXCOaAA62U8ZZw+bCHSU8GCZcmbWvGZqjp
d9iNzqHHgmw6wvWmp04ySVnbfs/GomiEScgythJZqPPGe956TwvA3bEO7YJcBRbv
ZU1Ekin5fpe6bf+jJ+vJIgruiQqiybL4uICZO00ikEwJeRZyI7DNQBMUh/SWnznj
EbWrL+k7Ltk/+yhqQsz4RyHlVoOZHMjguJ1Nk+k8qZgM9SZtnTgYpK5FNVnftJJD
WXajuZSRlWeh54/yCejDACUMtND45U4zDxGIX+VPvcIyvYjiiiif3LGoxxO+Xafa
gXkXWm0H0liybysh9hTCQILLEmhCLAFA+Z0F9qMQZ2VstfwYV0+e1EXqRWaf6Irl
tD3p+k5tgNzMFiYs/bICFw7Zg9sgzGZz7rYEh4r8IqJY0CD1ajBTE/b0QmF6ALeF
9ZF22BcKTGiWW1gR2OlDvWD3B9nIIU2pWVOD5Qd17pSbxTFJlHDcTpefyERXqTJ+
vQRU+Urhxag9h5E6ZZYSXhhPM2kV7XX31K+/Ml7E80WBQN8H/yz5dCZdvPGsJWlI
ziwTygyNRK9r52RPuoJFlRAalo84l/t1/dpGMjZ3aC90DFg/olpHlu5WDijwkFQM
m8Ahhy4hw64vnqBofAiUmd4D4OqXRYTgLJrfbPc7Z2rWEipKojhhPqzL18DfJGUH
P4U3w1akKG01FCA//c2Rf0R48Vo/QMLvKyetsLPMtuoV9+vKIDxrrYOcHQwtyu/O
j9jL6hTOwqrzcndsvzPdSXzAODP1wdrw5bxCgtnOeNt2xUBlGzyHIwyEBDRqB1qh
WdNe02sf8zuNyoNLMhiR6DBC3d/037KG2OPVouVQh+sfBZOGrJZfm04f8RqD83Mx
sE9rtofz2EqMV50hEXJuJTiYB0KmeIhzm8qXK/2YCz4pcKx2IMAcxOZ45jlf5zxF
yMd1xVesrIQMD9V/X6G3FABZv7PHhk48lwIuFlX/lH/VTOrIGPk3XrGx46nHOpV3
zjHYZ9BnZEUV8QKW8ushLNLInzFQM8so85U0bGWNL0V1Kt+IZVV59BWnki4l+0w2
0oarG2pEzkAvqZR1MVv44gbMEDykRRCbunrmDYzDOix5Maq01L3FQbcpob5Xipn2
6wuD0lOwmc1zq5dk3QFmRRqQLMN2+CdgOirdSp89jksnPQ0QgPywHYSm6zQIqQAD
h6flh9qH4gK8gpmcaVAFx3IvMH+sGyEe+LN2SItxpDjYRnM7PseyrYlc8bivmgIi
Y+2BlybPDZhfCYrLmJ2rRIBodYr1BQ6EQWCI9Anz9CToV9Z3rDR3EKniw3Lk3B31
b2viqbYLAw84lI+w7pD/cFXSi1WmJIdJOVClAiz5wDPEX9o0fG+jnFcXFn+wIAzh
ZSVU+vW3jQXoVyD2wxPFZIdeleNARWDgKA7rxnGyNs5QsbK5ASMsf41lVITzdL+J
LNcalfXohl4jAoxB80tXWMrVVcWsTc4Z4vY0/Wn/mdM/LIWOz5mO1JAUvIp6pEqX
FZb5+N/U3723Gi7y6iW3Vht2XyZ2FqlF2QgQivsvVEeOK8xadxuEOXQllrNr8o7h
DzxFd5pd9bIghkgbBBWQ82h9TcmdujX2c/ZraxhOrFn74F7FgvrOBHfePSwWdYFd
uS5OL0d12WAapGDJ39+gCSAKcXYBW1VgFweRZyuUOFs7jYCUPIug5cRgDPMTwUma
j3MIdWiJUKZ7qnFhia3dt9mO4T83tCQ0zH2+U6an7fDG14jZ3qxxC9gre558IduS
nVTvGgSX+Xaol3ZVXKjNe/oFtVTdacJ0NJHGLsXHNBNslI1ClcZ8n+By/bdzGWPZ
u7G+ugV3uOuXFzDzEJb4mZUl0B8PMUQhlRfm4fvRXZLTZ7wfWH/7kirleLoVKutm
NrcPAC/K74sBUaHF3RJZaYV1fvSUZG0EZQnWfinuXA4JkiYmDpBbaR8BHGQaN2RS
O9H32LIKThApxbw/HZjdsh8eA3Rcpf/l/sib2X5DY7O2rLTKT2FHEZGovUp8g3C4
awsGFUDs3VjmDr88taYXCzvSL1t0ZqXJzId5dNCjgQ52Qg7uTbKL/6SSEiDTxDYw
BMhq4WeeT4WKBzZDH00/qJnmqOOLXlE4p7nUTktELBVyZ6rNjzkJCvZhZk6Ev+rB
2iLnDEMqxALRio8gfHNbAKwo74DHj/n0hARoJPMR3BGC8Opjme+hiUaTqeRLliLX
kwVb2MOFFYd4HJpgjnLF2YhHLrceGjs4dLUbwjMxPnsECBioHl2rtImw7wlmmQvU
eqL0cMKtaqsTU3T7uf/RABHSssiTZSdvOQNWQUYNZqxfLI4D3T2W4pX84419kkYv
a6XLBO1nLUrqmxYooz//4xwPczDL0RhaCyyuPcjfnAhquEYLb2a/+jX1z7+LWMxC
AbU7vE4NIdqLhM4K50qityhKvDYvyjB7x/yqJjJQaWGQ9Hh0RaceE5avUN7M8iti
q3Nbb+x19TdaahFee/jtcBuOGJY9XsQYhsri/vaBUibY1RGHDD50WKxKwzSxsEBO
mnUG9c/Xk8i7TXc+vGDVneRWQzNGp8aKXxrjM7IbyYG3PCGg1MN4eJYPLPv2VGJ2
Ph4dhGNxT3MH78DVjZsyC1yLwuUd5xCf7AIdj53zLVAYB9qmB174IXw/CGJynMDp
J13k02qyvq1yuwkBO3NBVGq7szEWTGjlYZXM7JWxaeQvKiQhSPn2KI3mszECC82Q
sjFAR8MLGW6pR/a0Y+6HCEjJdIiLvbg5NpJBG88LYcKdXt/4Vy23Qm/O+zhhXqBh
bmiEc1AKrkbHiuKVMPw7PVqpzV1+ZmivvrB+2IiUbMigGgLkEIH8QPYkjiy1hywy
UJXZmbSQ2TU35zXSVmNi21+fxoVFm1/iNJtRlyL8Th0rGgrQEUjVHYvr0Wr4Xy36
ASIJJ6E2PiXVS4eZF57YcrAw967nlcHAHS7WAxO3eQr4ehFocxENLcInnIoFgvlQ
D9plMRB71lRsh/mMgf2joC9oe3IfOEkVG21xUiNXWvrpkBCAKjR+XR6dbmbFbCt8
jgCyqb3scGFKjRBa5vM3tCW4HZwVUwQsvSwTmaAe1Nn0mPpyWDKsvEkvLjfqfhig
5vPt1yRVNwVt8JvNE9AWCD/ubnFelWxKYvTUWcxXBaEjn/z6LZYY8F1AiAphMSoS
+fmheS5JIm6uQfpmam56/XfvBKYthfA7ii+jSapg9bG9/HN7T8Y2XCCP+ZX3ZLI/
kZhxzk27NV2H6XxuMF64DgFL6J5jH/nYe/hzrHLHqXqQIas9EswHKwdv52+HK92p
h2RZ1Ru//YnOJ4gK9h/t26e4cg5wiqow/Oolq1EZ+oYKnUiJloJMzBj/BEP5hmbZ
XW1uR2uIt7HORQv6u45i/7cpqPJensIKScqdzFaWxfqE3oV9eekvJN/8/2xXhNtC
jJlTlb+yGw+wzGGh+AohzKzy5UuxthlRj7ALubWYng1+u6yNamkRU3xnaMYuUH7G
AFLlULkqQU+6yDTyn1skkE7B+yp0JeFV9jNufEdgZrHUHDL98cNb0VGkiLKy6SId
rhI4rSr4stI7oRmWv+46zDBy4EUjXnDumYNHvax97dEp26XJv+IRf9b7O1f3804W
XqT8BtmbdnrNp93k8z1jg6ymGRBzYo7fOQG4kPWS7PzqAiNW5iSuMtvruksGkHXS
DpWsS+Pq5XMo1i8HwyIkhoD/g4G/fVvsON7sGaa9eWPqxylTnyoT3FjyX+y9n+88
vhw6ONRiyiywOCLnnYGAc9q1zMoVxulU1PovNRAt+HQ404Il/yY0ZU5/RSSdUl40
DiEBiCa7m4tBE+oOuK0dnGh5NLQVVyKKBjFpWwRy0gx0jtLERWpVfG+JmHXgR2rK
REmMyKT7NSb51FXfhuLlXrcBOprrTCwEfKn4lby1vv5Urs3/i3bPbkCAjeNT0dMw
QBNZ5VIdWGK6qv1eXSLSm6pvVYZq0xidaIg+d5LnblP8aMzVQatcf71jqSSp9r5t
0XG75qR3sAVp+H9IqM2CoDq6fB+4SnII24f99uGnDvYZKWs+68pNVPJC38U5G3RK
bZhTPWH971LYImTDvyvJFMzfJf0rQGm8+ATuhrNgFtKb+QwbVOmFy5/CTsYh59xx
t0NXs97eEzLgwY6YFHzt4+SfZsyAFmawKfX6gmnp8sBroBQWYSfxO241RjYUkVHq
+Uv3JC9ItaCIQz+IS3Rf/lVTouhw6toTSJHwTrzpdt+CuNvIkfYScfuEiBFazI2x
ePvJK9ote905Vbs4uGEcbNn24l9W06zzd8ev35Q8M14mcwjYeohSK0SFNU4vuROJ
ykym9siUvPYLfemv6A63f+uaGwy49mD2DCG5TB0JLggLWlZdVBccsDI39mh4u4cP
2C6EsifuYM0lBKWF0srVDbDdgRq4dtWnNtOCUKjeEQx4tX08o1fG8pNstoU1Vy7r
Y+tPGESfxHVsjVFSALmdckaNlPGuDKfGOSnpJ6SLeLGa8ENwWeJ+e60SCZ47kLpY
0NM9OO5BQwOl7AfDhacgwajgqzSbeNzODxoYGi65qyiTcNeIN5kzJU0n1AJcDJjF
Y7YqGN/+Y07Pk223GHWQmrwVZ+fhYvXU8dsL5dtb4iVbHZXjzforfby7ccwJiorW
CBk2L3WTms4Tv4PV50fRBXu2vol/sqtt5yAE+XPQyuZGcra+irO2QnoDgMl8fF3n
Fe+rCjUF0mrc06q1Z1c0hDVW++Fxun2qcNgGCTnpOdDQf091T1ZcVY3LQR6+Oq2n
e0p29Hpx9rPZdyzXD4mllCBO/FEFCvu7W0rYIUwLjs2Irlib18QK/j/NMP8TELEC
LpahKlrBcdz2mc07aYjch4DXeYHTI1zTUbENC2/5Ah6bt6ozc3fceig26afXDeXi
qKvJYGLhI4MRjABfJjINk4C/36QiyRZMarW33itySwOq+itdjzlpx60XwCHA2DUT
BQJO+rZa1ATKAJwGnW/j4Qavsq4Nhd4b7Mw9s1qju0RWUflOG6bnEAZbM4E4mYjg
y98dm2GvcyZgq1HWEjQUni0839TJP4CEKUnB56Kpl+ZLsm10APEzyFuNGSGXsDyW
CntJRC+ZxzjbwcjcIsIBdPGbLoupVo1sL/iIlovTxsQXlrucqSpUHZSgxweMlQ7/
BCCsqKEcATOTCdpPhb/Z4IzJTdKOn/PndiPF61Y2Qrgem54RTaYnoGLIQ481sjkb
tv2PHZK4ripNJNupRBC1PKqAyy9X3pDo+PF42Zre0TDXzGkM9hMe3627vws7oVSy
44U4NdVTQaYbKnQER0AGqHd/+5haL3Jbg0Gcclkx/X0K2H6HbOGwatgMkAKrTg/v
dbS2oClim0vvE+luDtXIx9OVFEyaRKb66pA2BhBfqfhGrH7S0UFGhZB7O0NJY/02
8JyWA8Zx+hhXNpHXrmP8kl9YR5mghAaWKpsFMPRk+RKbSRWPld7bn+acdzZ/18n7
chBH0LTS2xG3h+kX5zu+FoTyhognK2Yo5VN0+zwiAku8taxPqfqoz70jjoQTrjvp
crwTPs4KYWD4SRarqbdtq59h9fdxl9r9Z2GtV8MLnyCCmQPgQHWvxqJAi9Mrcs0f
x/6hEBoBltdqt0F5AiavbWv83At23BjYoDtwTQ0rcZon8zkFVqIYZ7akmkJ67qu+
yGj5ZHbhzV0QjNddIIBoSceUKsAKE1923ULAzPSP957OU1Aoliih46vmyqH82qeu
wZaK3LUwk3XQEr5Og6/j4qdzN8xXojd+F3UH/4eEHqJc8ka1cyORSemn2Ne4Sa45
Q2FA/De7/TdZQdIWfAgbZE6R0EVXFMQFihb+kpWxP3zThYBhrwNR42FqDhnZJEhO
MYW034gD766IDHqr7wPyabPabFa344wX//kiX8D9nRCMXyjAS5ceRiAe5mWJpTuT
lQpWwF6z7NX0N64nIp1wIz5Q6SdTyGgG+hbhgdTzfF736W7J1z9bW3dzrTvVVipU
H58uOpKWc8M2li1XhVgnLZnQFyJ4BVZiLj9hH3GthQ4iLU5XD6H8+nKE67UZzUUx
8eGjpdscLfh2nH/3xRP2lZqwkWRQGB/wlRcs9i6nieTP54ZaNx0JLVBg1L9QZ/V9
vjicqLqBbbOznphjDHVFw/rPGQTREyN4PYXTRNdM8CdQbEOe6bytj4U2cXLodiC9
y+iDqJXTCv4spWdIPUXZFV2JgdNxEHgb4MYy3xvb6yQw71ZMLpQQsOrnpKfc1BTU
JY3bv+7gOpkTNSEH1CMLHt7fM681D7u9P0cx+oJ1lKX14UKJsUa3R3jWTnAuFBlR
qjxC72A4Q3JGtJtAs2DLcTKUCHeuld09OZY64ULEMSzhjiLt3qIGz5Zq15mhEhuA
rM1xNK1IBrd34fZ5lK0jAoZeOJ40hsXbVtsYmPqn87uUl9y2dPIxqi/2HB4r8nGv
QG/usK6J2tzFwIXVv7eDah1qRYYoHacx7uhp18iLIjKerfpDUeH098Gvk3LAkqSn
hQVP979enBj0MEe7XRxaODUJ9w+SNUiEtBF57DmN/03S2VzfEC94hTTYajz9vvaA
bFunSk5D/7Hfml/fCG8IdpYzTME5Sew2pT8cvkwUa8bHIkcqpkqir7/zMNaLTbzp
W0d1U13j797OvhVEHK53C2ITJ9glQZ5JlBg2i6JNky7E896oeEUQHRGKwBGWrWh5
ROdD0IAoUk3kjVsNumeinoY2hw6jLlWEX/I/HzRAmDAX/i98DoQeNPeAvT88eWyc
/KZ83f5bSWFS4bvqtW1vns8FcOZNPJ4DyqJSQufIsY3hcGypIBNiw0f1xuaIQHk3
snLL0dMICliZynTc4pLO4a/5znnuSn70irRa/5KcdhmbNFCKslriXZ6+8zbcpg9B
EWidwikwzf1fShxub/uTo3s7IsDDz/Gd8jVGXmEgtX9TkCB1eOiW5VnmS2u9t7sG
KIoEP0GTr+QnmfGxOGalbQ0OECAbZTPj8a8M00JvI66QgtmaLLM4fhzVvsZ0BP71
vxC6D/ZIxBUgqmSP8UAvRoKU/EgOnBMWfrasBvVGrasbB6XUU2KE0R83lXyz4Ees
sBufVL7P4eT288cOMDXpo9xtIeaOh7uWraKULPGGivyWu8m+68aHTxA/5EjqmOlE
KoofWNqtjFxi15OUMige/bCuPBQvszWNzpl64rTbIy1gHCUsmlDQ4MeF2907ZtUW
84MllfVLEkueejnKX3LIOr6itPMd8xUbZny45Fl3L8gBE/8kLbbG16dVXB95bCWY
r6eOqo9DTECu+uV3g6pbKhHFBxlTZ9GZMfv9PiDJO0Y7K0wly62Q7UqDlbYsl1Pt
pvVZrBt+OqSe1zzKpR28nUhz57KklcqZNqC1mjg+bGz3spFLsOrPYvFi+N08nxkB
MnQwAB4ZQdEi4skm0Ii48Ty2ndE1P/oB8zVr4mz8Gm4/lhK8halVpVr2CEBYwSQs
ySCLt5lpe6HrNw5Wsh9Obgpc4qKUrb+lbe+YSgjh94hSZCuiS1VR8FVhhOcHGz6w
SHBGq1wedHdVhY8/bmDu57Op6MaPtqliqrUrF19ykIBPeun5NkO/fi7DPwWlSS58
8rzcraC+PAdeHEEXnjykVWTbx7TqnVeu/Zfy5jaVnxnslwYfxCOlilW3NBVIU1UM
cPTIE7OEjlvVo016OIn2FPRjis4CnkLzrUTXde6deN2ePXncFBWUApxBwVvrUgAV
5zpiv4zXu4scror+QLIQVayOXtzHbveswiQ3fI5JpslvgO5yT9egxVuUbQ9dvOFm
ecEDF4+DWRVjV9FA3TC8AU/tS3sJH/zK228tuSTeOxXM+rFK8gmzA6U6efUezEN9
EHKHk2rYdRsmQRF9ir0IrbRgYP4Cc7et6pKipm7IpKbelVaOih/E/aEb0M9s/YSa
QkZ6V8myTmd9fuxGIkY3oxQs799dyWjkme0QuaLIi+BTdF6Tff+yyusblP7011n6
p4VWobwAtQ3Ns5THuTBTX3xcKVwZExKedPP7arJso8bN19Q571EGOQtIv7n5SQqf
UrI6EnsXKBLPJBCFx4pNYHSvl6no5T/o7Hw+41H8Ks24XnEKrFbNhX9XLRUD5C/X
XX5u+g9oKKTIw91+Z+/QS2Sg6BMPNLu+v4ghb3mtVBs0MyXNfogc5spBhv22lLyQ
OU3huYhF9FIbWb5syGjJuc2iEN6angelccEkP+s83TC98gqnwje10wDSrlasrl99
I9FUpsOE9npBoVYSrOS1o6qjWp3yyqIfz1gBPOYwLwqD73UDi5mowkPBsZexBb5K
J2T7MEwEaflLdyJL8IxFo7i2yvGZ1mQ7Akr94TDIhnCaLHJgqOR92NHI9bGqGpWI
a1+XQxY7c4PtuhVZqoinEe2VwnHDQjj3ZGNdy/swJAtDQY++0XKm2RAOYgViUrrI
uNAEx/7Yvp/UoV9peW7RTvHSLgwBEhpdElf+p2CnJMvAAhhn6nuZ0NxVSXZGRHDQ
Y67cpRlpBGAlz2s5tI3JHmXLKWYTozhz0j6KCfCIdbdNriD75zrPRMXdGTCmCM21
1gm2G/amcDsU+4CGYAHubiB/ZPVSO/eCJEA2H52+ZBt2aUnKE5JFvGyssr0SOhV6
fhmn3/HK26hm4lWA34aJaL0x+kyT1biIFszQn0yK+R90mLCV3bVw8wTY3GONt7I5
ldC8WmUMheCKMCDh3fG1lgYxZKRr4hRlIdR5iT/lFGklvgv7DGGrTUfJqOvbLJ6M
yrUMtfLZOLgwl6CI/6BsOpTiHhUVxtdwySM0gB4T0vswoN7InCdrHaGCqOvtIuc0
1/ynTNIw13WTsuyVSOrINm7UReeLVYcmHWqDuBLoushOc2AXGKid0Ljdu97AMKjW
5GYnL1DPPBVCvXcJqmZyD+vVkMRJhB2/cjb+0br/a4wi48P9JAWS/6Rx7wdvZMO9
ZZmbOuCrlKlzup/tXNb8mu1SAkJ41gLzQVs4ccxCc+9Fk6OBmXTz1C1gZU9goEtV
lq4Rz4pBdeOBcr5LKg91cdqVssFWbjdFcZCzxr+UexILJXZiZR5h8LTgQGdYARXK
ry4PJPVhhuGn0nYRp68zSmua7Pskc5zYdh6wf9X/wbUrfB5f0fjMU6cvzeoVqBOv
4j6b2ekgy7iTETHT2XqCMCRNsmOQkgH1YGs/lH9VCLQPJ84ibHmiX6EudruxIAiM
/7Vw5dWhD66urXH5gSIzbQAuMPc5PNb0H7kWkU9HSRdkCKoRfEzCoCbWKJBjDPeY
YnAHpirc9n0asXY6ZX301fU8O9unHyBdT13DQEClMVP6lCdKsO4eGj/oa4U+mFBU
IBhGmZK9eFVTBsv5xNs2qNA5ZRHXF1CzSCqr6mDsxrn5yuEMHmVohqat6kA+JaXE
A8d1AB/o+J28koqk4XNn89x+L6lAhF3tfdG37SOD8/qhQlJ5iL0RJCHOaaOm1Fxf
x2eozMvausqJSfrG53NzbOWFOrQ+qE+ylrwli2Fx0CrXuRZ2ly5yivvv/x0ILaj1
Uh5Fxv/ERvBQdMEavV5k9ARG1bfv8Yij6CBShd0ovSnDuGY5PqHqS8RvCwnk42Tu
iOiFEL5LIBpF4P/K/b/yc3aQRytRJPuMMTeQJpnbe1SMoYAon3s2fV1TOmvBr9YK
sBbtjp90GcMwu/B4x5RnbJy7cYhpt0rGv9wXru3c4+cW9Ije4v4Gh+2u9ekyUk2M
7/7yECTS5UxZ2CpngCoqJtOn6eCrhtgyiJ7lg1HMfsRO5yvQcyjSztK9oCdeid5p
4XZE4+j3EIAfp4/kl4wltTcFNMYXrX/JrF9n8zcWorTSR45GvrlgTpa7DQAaSYXq
pEiyv77cfLoY/2AGgKaQ+FaASpF71af1hqssPMC8H2UFUCuBKhV9ePDUm7HJKofA
qc6QLFlKMd1WK4Y046PoZdrbeJIVMF3mzrhNPNXqLIyV91pQ9lbvcB/VOHTqgsID
izEJBvTVknp8fCt2MKnPz6f6XmOJbDYqBQOQtMEJEoUSsO9KFXYWaqiNpDL2QwxZ
4F/QOejxi7ElH739lxFzUaHskaExodWGP74moEYaPT2pHNYtcK7oICPmCGJ2wjPp
rcaI29rOS6+QS/U7JcT7/tXIRivB/5/rURSJwHWYwVHm1OiEUQf8RoO41YyX+l1D
0Zhn/W7VscTZx8fmoIZj9VUzPxJEee/Zmt9aWVsochUN18QQCuRauP9tHb4x66yW
otYNbpc+9MgT3f7wdeFxauo0O8ypTQrneWe4vVZuCAFvkLomw5TGUWeFNiYx/S1V
6mwl71712jDJubf2DdvFDV4tPUZC2KgAcf+fIrKu85+jeydfsBtdyAlsihOD4njj
yQ6GdfhaHaJl/v2qJ/6ptNIIvbcsLMF0RtHK3xDkyTebgkReiHdUuFhWkuoQ8Cby
DdMyXvBa2Pr13xAZ6bCjfu1H7GmfqEnJZ0BCmWLV0Ka/Iic4CWGjUyakmDmHqnFZ
QhCu2JyrUqdSrm1gtVB5B8DH9p1jAQAEx2QO4QfTxpcYC727mHVk3sUK3LsF4NAa
7XguHAl8yzeNjGeZEJj0Ov2xiA651aJhTo7dGbvYZcmcNxqQVoXpj8FvfoaWslF5
w1zPAUcJ1TU0JgGR5pZpPTu95h5A4CKJqRFlhc9ooxBov2wA0t66BQKLfatg51sN
CrRx1L8AzWDLVTgqAPvQ3aT/2t+i1W59d0TqaAWGfA8CbYqknL8RQTAoZ9O+mfGb
qGpbW4R/AVbAlseWJ3GtWmd9yjUvJVHRFGkmt9XIOjLvISpJrUlHgUUwEslP7Jd3
ZuT5cWYgL5BNy3UxcV7OUiw/Bc4LiAKMVvqcEYg0EZuBpSVM5Oy+VFASQgnVePud
yJMFkmTNvAGuwcUz5A+kKZBrbOlcRV41/OI1bA9tM5Zu9BV21LzdTJRJBVt8pksG
eWOrNyV+t00xvJLVp7kom3kkY6HR33Kll7bgRRjbrvM15V7SinjCwyG7qOfANKEg
mLSld375PrBIBUcKCFcm2FZ9XVWqyF0m3x18TL/i4ZkwbnL2cUaXO13ug9ExM7js
/cG5vFJSf1GuvhHtb+KUS134ZQKvzAJRfJAtvXax6vXQlK5bf3KdYIR78iBozENZ
T/1UH3CoqzrVuBf6rN9TT0tow6NWwJEJ1vZXUdsC6vWR/rkhFTXRUx/0GPNnd5OW
UhEpQhTm5ceQYWOQ4C7nPV6iDAiOZ3c1WMoyHgVxyPvZc4VcopccnylfGhwPJXI/
EmsTy3ali+il16lX/zg1huprjexcLxBirGsqVUGTgaebE8RrLWsW8+2zvUG01uTs
zjmZFzY0QmWyAZYqzhNF5ENp4ewOBFteQHrDdP2W5vTKy2B4xypBux8663xEJLD8
F8gagl/b2zMQN6wb6ppQEFi6tKDSEB1SqbuNK1IE/yiNeWWNjFoUC9UTjvkbM/oj
/LNiAJk9F4Tt03d8zK299aFJdI+7jy+U2HrUwjHPXRoeckelTz1qLLVHn9BM7ZKP
OKRuwNQDAlyLQ+qUydBwr5oY/AlzcF/SCC+ebCJvYzN/dArZ8yIxn6VlXqTmadMZ
pr8TKahZaIco9NZ0aS2vzbh/IecbyT/Z7iSHKVyo929UWjNFke0q9AHYRGUUbcrK
tsgK0YT9aILQpFJYFMCYGBrc89SjDaMMzTqZup0iDanxNYARF82YVgF1bhEDzsFN
/o8KapxHzgnh2n8DtJIdylCC17i1ifW5Xd58Z3bvUNmvh+HZaa+21xyM075QF3Jk
iBV2PsDbugqkOzdwTioqrQ53B16kOHJhNtoZZTgWQvHmOdCtd4+9YLzNYv5CXxml
M27oH4e10EiTcx8K+mltmbmqu5o5rC0dwhHHhejbZCrQ0gbFaYJLG96bM10TJE78
Mv2cLcBXe0Xlkem9U1q3k5lqN+DHcTdXF1zUUmR1Rhc3rKGzYvTdaiSfW6Heo253
bm+CwFwscOrsMJXtFb0DRyUQbldeAa2hhn4oKG5DiUnHE7fpiBJvGNiMu4zxjumm
eVDseb7gQiZphO+xkU4Vs/yoYKHOkXOucxRgfx8FT6SFPPTwPi+YIjrkB6a6p3J6
DBZCM4KCL5kEIV8TWTBmK54Jfh1vPMKPkQ9Rt1OHs9CYmWInde2xY83qWygLLZxf
9lTEcbwcKGumT08bc5FxNHTlxsm+N7cmi+2lrHv9UO4krux1KEg0PRhHY3k43Irk
FJwjFm9zNG9bz6pAe5CbHUZ70FQLxSAIQIbw44kj3aSr7tRbB4UclqSRb4GgmW5Z
XZ+JUeSf1ryYNP7o8riUkQT4RhxT1IDs94eBBDdL07WJuIoqSAHPg4W9l2myXcgk
ElemOZCEKi9bvFlNWSvmMcVf8xXxDCn0v/pcVHifrA50umwn9bwSjqU7qmQFssJ5
xkCBFbJgJ8u5UXkU6crY+P5Jv2sWV43XV7Abc7p04PV5BZQA/6gCu2pQaWE1QpVA
HfWHBbpp2oDpOAnB9SUTULUl3xMrD3erwHowg44g6QX8nFEmET9t/LQoJsT35hda
HxtZwQc3YnevZe013I9WtYV/YBNebsAt8wNTrwD2XuQEHg/5/U7kadEy5EqmX9le
b4lEgNnFILJt/VuzCdFTzg/EumoK1KqPdpR9cqiLHam/qa2QkXoQu0TMT4bgUvmp
Dxsu1jbm77us99uD6dNE9JZ/WGPgZeGGonwRsJ360RY4BCc9E1MO9iHb89kMYTaD
dPSCozphzvyz4jOaYGXnYYbswB0bVdTpbBCA35aRyy8qxZUo94cPUZ3MXV+vRmCx
G+v1BgCaK0Cq0vJNP0Vs6jmgMKNYK/RTsB41j2u+LY+LoWrZ73WiflwkWlIUpyWX
vL4Jd/7dZNDy29JL6Z/8Fxn8Bqw45w49YKfc/gehzOV6UEUssJ6HawjiHiRsAl0+
ilSXYvEDcybLzFzBvBFJcPtJbaPXpiKrVR8BtV4OpiNcWtv4nuENThfVd+KutvKM
6EVUsr0YWmvhD50sgMuBhiDeFOBTeD+NmGSa+mxRMQLoSBbLC9MHdyq6DYr9d4IO
ob7naVkdyU4y9SYAVzV0ABoFi8TSDyFps7PtpdX7yRoZE7WMhgGYz7paFeKkdrKq
VHSQ/jw5yFEVR7BmOSrOsVhmQRIcCoIJgFP0XrF+zkqlYlThmtHOAPoc/J1BDToG
60Tm8/kjxKnSqiFnckHskrECFnmNBxAmYrkbR0+wl5s7ROxlylo39Q1rwZmYpVPf
JBx48E3W+T9pN3J575/Vy5q2mCYXdTFnqIQHbE5u/mO3DbnPJhaV/FlagGtgLpGk
U1PvSgZP3+AlTtmVRFhJQNJqsnWBC202/5DYYLBsexeaheQhqjALdskkLKdYWtFD
SdyoX71DXcBLQIGd7TEsrUDqgF1ove1QJRTkJgnTFkuPqmLbNTnrgzKuGcQ9xIfY
50STf02XCKKp7nnKHMIbwxYQy3r91MZeWgF26AIrZ+8kzuMWj8xEtrelxlrq3DVJ
IzSfsTwQPOQbDl5NLnFePu1liN8hvfxXbdzpcQ3fYRurVeWZUqhDlmph5EH8aU2t
oGKUAtkmAPg1O8zayrGnI2w3YLKRG/H1JPBZkPKY8KKcMAu7P+Y7XGWgtgSkkdGt
e7q5LKmyjL65xXYS/9r55WAESH9Ma6E41/qt2VGZrloTmVf18nHD82hKpanNwmiJ
CtAx9hUOK1MGHCygHzQVTYwwDZKQ6MedauAwHAbtnWFOdw3WOR4uIcThACB+vXWP
cdRk/P1C8ztIb5P4Xtv4RjS/ExwqU0hk+KPiu9xBV99fu4TI/Ln/D8ISlVfaPUOD
HhiKcwFHqKwB8DgQ1kiR0k/zMTbgmq1ZxJjgaJVqUMqsRuiiXDA8n7egMunYx9bf
YZR+qm31qCXuHRulybIbldjAThB+NHrjvbx17I4W4EJ8/WTlTxDcmv5I6/sDPqpu
DrQ5IzbhwR0AbdYJF/r8ptPxyi4nFpgpVMBYmwbtAWLbC1JAmHs9x1SIgN3puQ57
dOFBl4Nf8alNAPGMEZN6QtajiM8f0Z31jMXV8PYwDTbRZC4gnztqpcr1OKdgCEqy
UXh8j7kWxHGr/LZpQeI6TSunBkEhCwUv2ttZ0wHmTUMjbzc/sfn3wp5xQJ3oY9+g
a1SCUFa75wP6pzR4iZwTlUk0FQx10Yh9gPuDF/M7xUufQZjujHLbAK3GakrPL4AH
SN0idTcKr4+udoa1gIF95pWf7PfOlFa8ZzptvlDxyc+uPI41s2joH8TkxIZXtMFv
324vhdZVFo4JID6H2d2xjDqNtA5YFZAfxwJLt3jJ3E/GybnE5BULx6u2nGofTVos
AaGNByz7yW6N8Jf7ENaPwXvj4xvBMeQoqCi/swC+BDU8m3+afiS9a9rqIU+N8yPc
LzeZCSFHnRtD4f+QAt65ic0WJwx19uHUdhMgihiqS9BqwNLBVnr4NbjmDWEILjpA
gnnQjieF9T4drudgOSCkAiXQP9ok45Fn3qLjdDuU4Al8ZDJb4VZ4kBupDXu2KAxO
Isrm+oy/vuU4NpWgAGTfDS+c16IudmWA6l7/kbCuUvdpKrmkQTPUouvD/zhY9vfd
okdYkDmkcBjPI6+1JsFqAzCt1FwqNu7pipOx7/aVMqfHrapLZBD8Gm8xh1gvmhRx
EzbMCYsgBpb5dYFf+ixuIrQ4u8wefkNmouQI7fdPJGepz9AlLiOUSrrBHfMz0zfb
zT9s9aonVLk1I2duQwNX+12+zwoOI/uVATJdWj6+OrGiPm53MehUpL84a+6Gs0u2
zoLE4/bhqIUg+R0AtsTTq/WlS0r5404tQqFuxdedDMJ+2IAcV4L5kdZmdJI51L58
u+OPmgbaaZ0RJ1rMa0QDFbZg9cVWax7T5xY5UbRkEW98o24fNu+v47p2vPYXMMcp
VGqi3KUPVWo51c8YDYEsmwEgFqcbaZcTvm01o6P3xqjzO2S3G2P5asl2Mh8J3Zjo
obm5qy104I7pSNi0LSfw/A8VTpLBihWRKq/x0nu3WyVC36Wf1jBow9b9TLULgDux
UP2lu67Zhan6Q0dqcYXKOPBDE+pRY8g3uMvaO3E/g6FDJqzj8nnNAwH1e3Zfso0m
Wxq4GrrhGPy39czoqFbfEZjTM1KRwnJZT1kx/hRapUWYm/wpW9hdzj005zC2cMWI
wRWxKEutpyoG8eEkXevd47Jw1EkcbB9gKPQhZH1T+wNAQ/BegL8LyU1/kj3Pbt61
Xv0qjtqtbCUjADfcpjRquF3FC5jGrl9YY8ufpC6W1ysbYdtuK5O+M5XwZq9HMn7u
LYf8C0MQZwWR/VRA1gwQ3T9d8DXQKLcBKAWUSjdmGG3ycOz5lxewLrpMlUYPZt0E
VdDXJoj14xBPIeplgXPuuu+Zg5jkJvnO999+W1aOfS6e4JP0tl342GzLEm+7BJ+F
kpIkWku2Z0dXdp875PBNLZKKpAe0HB3WgLaCbmb3IDE/COSaKlg2SLzMwnrxhMEf
Ug3osdsTuoRp0jAOqpSB4HaF8ZHhX6P5PDci32/H2mo0Lc3deC4Q/tiCi7zwQhNe
4VQ15nwUZXeZ4gFIjher8k2gvjrOkEKoY504Kw6RYXYUbH1xBk5rdWF/ovjCSR1k
z8LfizK7WyFEj1YLc0ezSaT2/msQgtLFc/sizqXInm1Sjo0dUytYo8L1B5FEGNpu
Nm2IBD4NbO5zxobq9QgtbzvKsTDROdxKJ8xkxlVuIyetv/O0N27oWPmxajI4COL5
mQabOBXH3CY2swwKQB4a3f42/+aUZb20VZEdNdTAp/arZdZ8qQWwXXAZzcQVe1IV
ndyZcYvJe2YGEYSciiyCh1EPxkQNPu4oAgkcF2kWE82TZyzJ7ZBrVOS1SWiC+RpJ
i2EsrONbUfBe7rMch8YXjumpGo2A6W7Kl4qHnhyItJUUereg54wCTpKW3FZtrvfc
KzKjrxNIVTPCuz1BKJMeMYS5I5BWeG9n5U588GBd/nGsiTSMOOen1PD8GSOF5L5O
SjBOCvmF3Nvb22KfRPT14L00tBHhjdQAGC/zuRsRl0eFHjLyusHOa311ZBx7Iat3
AA8sEz9EbUvhIYCLoPGXsebh5abv9xQRBQGjEzmoOHPaibdCyPf7s9PvyAIkayKI
ekq1Tsk8+Gv6SHiLGeaqOMujQXzLSwNWcTv/+H7UZgO+N2FEo4HnY/oZlLO8K9bb
VssOJ8zm3byhjVRuvATK5SnlwfGrGyP7RSQVvzQY2YilGtp7C793xcAEzuZHNTax
Cxm223t1nzubBAIU1nXgsmHjPNNWq12w3CudcnMZXQ0QXS6RT+4GVToZCDbNQwTM
ytpVwy9Dys3wb4TaJLhTl2OQrbJKdXWDlcWBHyUIIJjUa0ZxOaPMxc0aA5JUcEF0
zpBbqfg812ULeEvOCfxWL6d5Lbvaaac+9TOtciONSWd6XMhjDTM5Gx/y/1VYmT2n
g8DiUbfjWeXbM6dES23QApl8MNG4D46dbq9Xil8Wy9rAZCh0xUBnds0M/LCEqpp3
Eg/jSzHVkP5bp2ff/+u/O7YGCNnuBELDUq6nZ3xF03Enz8slDKnkhBccf5NkigrN
I8F/tWNoPqfhc0eMSAF12ZCK06aDyY6NCkaVv4QTnIP5p6FNhcrpPHk+3Dxdj3Ir
fabiLB3ewMrCByHTFWIRhw4wRLCAAAR4CX5DkpzFcMHcSvXWeYDmjSsQnwTwdOYf
Tw651nCxnwidpq6EvJvRGMdzLd7tF6g4l9xADyB9T8ExqXwbsJ2Xp/Zl94qvMJyI
qGudXeqKyAi8eipFVxbnOYIvhNqE8WTXvnPBInYg4Fl1S8uOD277He3h+U5uGJNN
R9zni3gkUdKMWHeZ3DIWKmSaHbSqpUv0nCcV2Gar8V2iBhHrucQUGm2gy5UzbJFv
zh7oi+1JTT5/YbJnZjxMgdEdzAadhX+0AKdGQeRTTNu3WohtasMKu/8Ppg4WQvRE
0mbtOqxcL0rWwP29FdEvTZ9Ehxs5q7Cts5XPngv1L85Ss/o8GKzPoHYD2O7wdn35
Y2LRW9Mgk33cpZVw8OXvZt8cEIUqMsQito/N1xmU6BXwueeGRA2e5L0n2YwzcXWW
833ZX8RLp7azXPBhRpOYDhkmoPf093HtWxh/KMaX415gZ9WfCGSnR5N/EmeGVrc9
AhSGz52+E0btWTNHUYMZkzDaTRunAffp+juBkuE6a5+UCdFFIWzOMEKxRnPpxRVl
4IJ5yDbL2PFhP9GKP1irwoigg3c4aehRcDstBr1fHSXpsIedcTW0GmB8P8Wwx934
LHddSASw7gsMZ1m2bAYRDwfM1gPLtwgWK3uNwEF05ZYzAA/EWbTT10F+Mxqq8izG
ol7NJleYdL1JEdHD+zB2ugZWrqyxilr7RwBB+gj1iYdXxQTE2ky13i9LujgDyJNd
4INKbZ2RKenUwz+uuqctJkpxAHd68Ozb75rSX1pTRiTgVR81AJpPKwxgdJ5/l7Ir
ka4lmgJz2W43h37DCp0mbKnghYzdjE1/E+8aFHIgaewacqop/aLMUD3n1chMTH7k
iG9ROoi6XE2VmsgsvIJsqvdYKGYnwRRBoafk1nu99d/9aYcHzMQkabgYiECq4flw
iELbaXtln0lE4VFfvPy8ZN5hzxT2CkQhJQ8zm4bFnL146xMMP0N/Gl5cQ/2uNANB
NmvNMBWCJ28+lEntyc5GO3s7w20aC2/U53GYA3pAZ4+88qYiU9rntgQD+wJ6jYKg
p3FG7xqFVuBT4EfyqJOTqjdPXi0G5LQcCXdGeS0ggR+mcAdkRFEs663sQuRwClp9
5jhCBk4Qyn3/cK+BwBIXpvBuopfwoFz7Yz9gEjlcwvCF4hMEjBuTVlQvSA607jJ9
ytuJmCALypz3DQkKG1U40RFoIhD6Qcro1Nmg6lRXY24TqmMI6YlHOaDuuIHgMZbv
TiS8a2wK77BSnPuy7WPS1NRSW7epVMwbVBJ049eRBynuS/+muaePvQKcN+Lvzk8x
dBUdKYVJlg1OCJSykpYmqPDydi8KdiISGfcUrQbjUML3WKyZt78ZpI6MzLtRflYZ
dmS2twJ66ql808L5uSRENy+QaXqI7h41UFJ1wBcya0H67NAy6lQEm343fUdjsdBE
OeEGVAzX+XFFwFkRIYqbz6HzCde921Zb1b+tN+u97v9eoAXkMUjqdBA27U5JVERZ
9wR7OO3/0SAavSQe/ORCDLyE5vu/1/bVEjdoAJipoz85a5XNWbbVrKGCWpupYlqt
zqRUFHgwbkFIKCaYzQzxRQyUoUOCqkflzw47Cm3C7Ow9WFHN8F/K/1UtawMr9LVI
/Ojan4NIoEwhDS6cLG337a9A5H2J4y2mHvI8Z5Gyi8eimsMtTNS1FgmZJ1gOCHpy
MoE96iFvFbvAcGcCyO9mMLVegMlbFo8rzYX/nLi5EY/lKbwv7rW5lCbfvuuQs+85
UaPmJ/e+O1pX/HMR9wIx1KiBQ/ekwFtIr0U1AAchw57kq7LnlhHcuivvBwy6CGZe
Ugv1ddr6OW5nmjE7+QhWTh9Ii16imWwFXGPFxcdmzC65IBHf58vh4m2p6jQRiUdZ
v2bX8ouS8LVvMluRDSduVFC0X3kLAeigcpsB9ZpHce4daKKjDrte99KI6DQIa9xs
NaDGttkSAqc4HPenGV87o+XXF2hnzKwKJc7ln+2p+NTBfdEHtQDyIVsY2eVB80bb
FLhtNWHmMEX8rUSeiUIimieqIBOAI1jFS7YgZhy9LLvn4ZjWhAKIdSko23IlBF7n
S78yc4T9ekyd3SYb5XUT+2LNWGslx4RIjCtjs32tK5i/FO0Jf+HxBBxw8mEu7+1V
83p2lHy21p2t0sEimO0C6L/+wHyKi4m2iWWNGQNQb1CMmmNSymutGcqwzShhP1Ei
/jnyX59Y8X6JC6BkxJXRR5nD2janY58sPFJ7n6k1G2ZpNrynDFAoGMvaGBMdTRC/
w83gG0hN0gldP0tRg8AvJ9utf5GrfoHNmota4lZA/uD5SsYzmdoItQSFlWJQ3JQS
a/8n9cX93lOfCGQy6hbWlrpM0NIhZlO1RaYz+ZjnQWILbh7GD4aEqnpXFGQGAyuX
vNrgKl+5rC1FEOU56o1LQ84kOArlPp778lxGUBvVp5+RdO7lkkjDzCFdY63UofLz
xATN0AKbSwq++PW4EC8xpEuP0dQGyGYru/K+J3be5syDzL/hDrrzyFlw5Jt1HfJ+
BemB8T+rbsrMAK2y71OBFC90tjD5u+JdHPixDY2wSxDxJ5xEp8wIcH0zMesnDve5
JAq/9v4/hVuCaP7bRsffA8nr5HZcc6KRLlTezxk4Ne63jgsUa2q+EL+6/kI3Dem9
LbUtl7xAm4GIFDgNay9VMs4tqyCot4uz9zoOijuSC0EIzrsJJ5eUshasMbusT/5u
vV+Md36nmBCRP/8sYpRQldXMHbxatQ71+Xj0GGMx8AX8iPc4Ou0gDLBl0qWotNuc
nW3x3mbFEB1NdYj2CuU61/6VP4stimmlCMDTh4PCkv2d+emBlRmQofNHAMXLHe5U
QUnnHBSW1Det0VcKh319ngq9J9b6Pr0SWjlTNlmBFRK6nzvK3NrwpNGh4WHItcEG
w5bf42hn6UBNABZQ9fSyfLk3qsqJdR2nkJij4qF3ezGxMlIYQrf8fMRkwZ644Rmb
3J61TSA9YaOvaVphmYjfxptH3fmRd4iKaC50XrUGR5hVHdcPexH6OZBbcxvcGDlj
79fg//116DCW316uA91DaHnHP7LZyBiISVSrhLxt4wWcw3XgfgfcGeMq/hy3/HcW
BQsEk92sPjmgRMaVLgehJP2Qf84t1svLDRx7Ge8Jx2wItENLRis6knHK5xPpqJOi
xi2YoafLo78H2wFl19+xQlwEijgOp3/VF+B980VzQFpnQxnpRoHRyADzajSDikIT
fbT7Fhs5CERDzOC+H4L6h1v246Q937lFoi62QoIgaStBuWocQEjw/gNiWtxtFUJm
4X7eDXNX0ehfORnwygpJuJqe5Vj9PTJiHej96DQZDFIpM9WzztXd5g/S2gYGr/Rr
NKUr2BOQPIpSSjdP+IMo0AdHgbcebJFPdpKZAGDL3KLavy83LyngL9KCJWEKGkf1
7x6lKrUy53eLuWC8mOkSGJSAcXj5FSiIfyBHzo1F/AFvevLt1MP2CQDkD3jTIs9g
UlRD25vd1r3WGA8+4y9p/7MF3YTkP8aOzaC9ABzIyzo5jPvmAORRzs8lw7MeRX8z
AtDY5RNds+qawSHO6j5+lnA1nU7gZ64g7yp9YMoJgYKDHV7KrNAhcC4IIP6uYHIu
VJKTa2msW8QYnn9Ag1q18E0ThqyINV83Kq6ZKrCQnVe5qJ/SYQkHb2AdwTITPNmj
jPxdsEh8OjdlybXdGtW6P36S+866B+RAw2hVkWp+ZbvhjjDO1PnVVX6StAMFQIJL
+Jzno9qsubUG9dgqr4xsRHmM6MitnzagSLkmOJg1tk70kmRlz0V81yL3WuiRjYwJ
6MLPnqutdKkQquZUTotZM9lZpbYgG5204Io5CHx34iGQM9pIR07yn/YpPvkX4IHM
bsPRStDl4ZOTtHY9MtAIBX6T/ih+a8ZOXFeHVMQ2tjalw3A0Zp/KEynM7J2iJLYq
UKy/NY5oby+gVLdclOaAGD6FlHlrMDxsTRbk+TtKcXljcDbZ2Zzg5YC8eR44d22X
dbgtQ2nYNSg8elwaG2I9lFuNmCbq9aKp7nfuXcu3YlB01Wq/dDB/8X7y7imYic74
hcyJJ2PcEreF/zFoMtrWstgp4uuwVsV6Tidqed15QTE/zgWHRUM4jN94so1WiNBL
on+/u9J8WGyFsKbSRM20B3PxOQwbKx7IwYGGDiyK5M8WW6ML2b0roW22fSAsEX94
32MLjKiAzM4tmYQq0PxD+Am5KuoZTBbMEmaUUHu/LuYwXN7rzWtIG8FxwiT+Xd3B
mY9V8BfwhDxeOpTbAqa9L1ktzqbWvCB3yhh0X1YBaGgSe7QjVZt/LSPnKB0ZXwzZ
lt9+zVLA6ntv79NPzNHvrRxdUSEu1906kYNgccA25cYkAGEsJcvU9Lx3TTxC/4LL
tCNYg3jbWaza1WzBukepcTA1LtDc6NhT6yF01DuFaeqdU8kSR1AKhqqrMCPrLqn5
WrqP9mjjlZaXMUzfRHjSbuR019i0UgjZTjINxWF2Qptf/uFhlGrePDVer3JnvotR
lw4gSA6jeVNpcobjzEM8/jf7EOvm6knTjeLeKoHAndHYZj6NICBqegeEN2GMjFPW
w8YmeIqEIkyAgU7Wea362D3g+eb0MVQoPNXJtjYVDITt/jONggLXz4EtNuc8Q6AV
ZCA3vbqGxBAS6f1xFh5iAuoQXRwEpNxx5JeO/ykI3ixGtOWEkRd1WEADHl8Ou0C3
C8o1xTiNT+IvSelAgohorD8E+JlO9Zo9z48tXDTygpHvirNcnHVocX4+sLSb7GaF
ab7bIOGxZaptVm+YxN19m1r2mouf0j0TC4uZOgTz3jfdcl5NjgR/CA2Pt6PB+sJK
I0V4WG7dova3MKEwAdTvO2jwa5Gb/cb/lQfL115onEq2vWL+6MUyZZqeRS5QeRVg
v4C67OWnEFgAwJMtcSspJHkuMPCcjVWPHJdrfWuUQz8HSPrf2oRj5U+fo9qwhHbq
0BFW5Xnx2xkHXiDTOJEeJqp2rRy+lO/nw+f+0d1FXh033oz2h5g7ocEfATXO2G8E
oSHPrsAd7YHKRRAcyg3sCmaLZANHefXDvZShzyulp8HUtCR+hcOttqKKg6+mjCAZ
k6S5m+WeXCmmPeygx+cd3QdJlB8UroSgOR84IJWcC9C+xmkF3NpwL+IwcQv2NKOS
2AiyYxDpM+fQ5W4l1FpcUfF5BUeX71yFwsCLTS0705rycDImlcB5xx9a9CSLsA5P
B4lRJNNB65NBVQHblTgw/M7YJ1qfFwKX9EM/2i8nF22xJ8Znuidr54S534/Za2MJ
IJaaKxF3aCoGG10KEyld1u5bpc/pD5+Z7fhSiQWdeb+fA+PBWQMGfk9nnR4qkQX7
+TmujBNcNqZqSBW8nCTSQ4Tn25IeFMOSMP32r40gG0lXMjKR+reQiiGrzVjJZtMS
rcZJ2xOXpU8nYW2XbujJXn1VFVkqNvBQczPExTB4wVZBTHFFipjJaSbNfJRL4Euf
scLfqTgUSHu+tpdDVv1/B0Drnolw5cdNCMamIcyUcUd843POrrZl/OIof4B3YHLm
RYrqduC4JXX1e4PL1Br99CM877nkYdjUyK3P1KLkoE8AZPEN2V7+W/ZWBa3w2ODM
EFOvJ+H2ty2mIrX+Xob3/2M/LXUbxF1Ang412/C6+AXDv9DEpuEmwXBZlpTOBi5l
8MS61KCgnC4xh8IjlpbQVPS3XXflxY/Sg22xSJwcAIytSEGKcKlQ+zem9Kji65Dx
W/uv30MWv7aaZoYYLNg+c3YdyykvpNgWaxGSBRAsEo8hrOXOuVn/lGbGFDBJnSCB
BSRPgzRHnsVCmZjM2Mz0+O03AzWUHRhwwcqKWh/1fnySVLti6PBLfqqK+dbqwtVr
duLxRxjd3piZo2/rgYWhr4R4Yqn4APrs7/pyMcbK+n76uqjRvx3FPTMBpDjPm/Lc
+MShzcFackQsg41fjIVk31LFbLFRWgzsBbhP9kML8NAfbcCgPIVHK7g5uyq4+1K2
b5OlDphaw6NAw+88psS7rgUTOOy8g/L415VZCjsfHqHoXX0QaUppJ5RmafXpSbta
8KcIpZQUM3wORmc6j4xQO+FTY9nHuIA3nNCP+Zjpo+5XNw2boXWGzx0UGlk+VwpJ
WQ27JosSwKj98FN7fMzPO4SZzWzEo5nCbm013YyQDfo17F4A69cClqQeypYIb2Dk
56LOVMFhJB0UkFEk0F5Ytm/geTQyCyTempXYaI2QmHUWhs8xJtKSCIjYoQcvKJ9e
74Y70QJn0CJvrTZLwW8OH0EtOHeOSAnROCVKIbD3qrgnumfR2g3zYZ9tC4u16K/7
4d1y40SwdoE9XpHJS9AEEDS0TUQ4AmZcIMVrual7ohFrOUPJKmVwYzR961x7nRJh
/j4B4/m/+URQ/nAQyGZ2AWaTbSF6d62zdiUsoCXAS2mhRGun5+KiwsH06QyuqJvI
ep4MmKVLNJJrDcWGdA9PXNBRC5Q0px6Ye1+ZNJZWLziU2cNmfxDDr/4T3EcQk55K
nDYDv6Zk6tSaAgmb2m8+aUC0xu0pfqSDYDUjM3wNb2XVMRAv2pnvzn35gx6FoquZ
vIG+b/dBxoaKvgW6USLH2GS9AlSLjjSv4PotFuBpVzsRdA1O4+MNU5H9dU//UKwu
fIm2HwuAkCO9VjDxrmYNyqCrugn4+DCSuqjHoD+C/oea1bEWKgC1Ce7nZ9O4RoeB
eB8nws1wteRgudsebMgtZBIvsnD0QAsLjXbDqiSSeqBERWMCmKDBwWq8a4Nar6KI
f6GBN0ahR6XC+zmPFhAAbv2RmQxVUcoI9Yebh57BKdmDynaVIH9q+mkpL3biQWoD
bK+RJoQUBnnG1GIuN+oeBYHBJN877pof9+yUInme/QH6SfiECksG19LZYKowisbv
I7nS2dbbjoFmVHViQtzRukvgSCQEVhR2jURaz2iIe6X591JfVLmblWFD8SmnVnnm
aAEOkYKsmkAxZz+i87Oxnp8vO5TcZyfhpb0cAAZgKTI8q+40dwRm2BSKBC3CpxVt
zUhhhxfYCIC3NfyYYVHOXw+hnasVa6aJQ8a7ci+/Udif4jK14eru0WEH+X40kTET
b7JmYGx52Cq7Qqvzv+2fU8pYVbKFw6aXKTX0KFX1cGEsAWBguC2eAwtVEArYqEul
ursThlQ1w3NRjBg/+PCEpOTMn23gahpd6GlCOIfZC9Ay6ubALHyYKlwc9fBp20wR
O168rEutk1kPiUqVRTeixhvVedGh0ChGEVkJkJ2dt4FGoSocpvRIk1tIsIK1HpZP
AHxhZTT4mFc6ynJA2jY7fVVss8tSRtbq6Hw4ZKQSeoDVlR9fTvgvB/Tq/gBwiHOT
OuZlIL2XyuONxnr0LpzChEA3nBdRMG15mb4ft+9kGFe8InQ12TdBMkqY/YGhA+Di
mrPJMaJ7Gc5Jrv1jX1Wk54iOXLCp0mHvsOd6JwyTMKUSpkH9eg9cUt8sx99lI8ue
etJB844qSD+J2Q2CgtrwNRULvVwLj332toW1J7R0XaAXiWkolBiOZtF2GZCX9Mkd
shZ9bfkEeKQxU1/HLXYh7MSmq52HVp7Egzy1Wd3y1yTbPTuYDNDodtPEvud2Qhus
MLPaybMqaWzCpPXtIcZWt5Ij/06NZfP4Y/eLIKfY/PwjVid12EFvhOj9qfWVlZvW
va4JpzSbJIibopekt5VONBsK9rpKiMmwQSuHOvMmd60XXtiNR0/FsC0jbHfTWmZf
yZR2RVYhi0I5socvVXR1buhFfcqRhd1gnM2/VNL7Mg30SjDYwouoKd+ENlALy22f
yAsJJgAx7oA4BSYQh/suvqk6SemWk5SzROcaQ1HIlnJ3iLfNoeBCNI+DMqIDyPjg
BqH7tuhh77RqBgqKEFxOhc31P8IY0u5HqFB7SehWWSw5IWrnwBi/1CGBXlD7FYVj
rpzEdljPWiC5VvflHM28zMg/lZgm21VTSNRm1pcCn1l6iIR35m6NtxivMNeQ3B5J
rM6ezdvQcMABpa0Wyi9DF1FOAXaMs37q1G+5C8Ihu0vgoXR3UgQxZqKcavCrcuIQ
fxUNnz66RvG5+Ax9icwai1Mk4A2YXtQvOoffOB56CsJbUTru8kx7NGP4DAlA6s1t
3MBXQgdtmGbMfTvkOIo8sP3KTs05TFF1rezSAV5gGypUxhwyDckQMRBawUqD2kgq
/BJ/3WeLVJd0w5XH+hx+sxNpXcB0HOieFF6T6bBJrHgv5Pie/6fh36vbLYYkuH9Y
k0y4zPoA0AW3+iv++1jBrg5aT0Vtd/biSjNm2WpAD1jeqfXBNj4fX+dfZCyNoST2
SQ8BY4nLK3AgitlCOzInPPvmePEJ1dC9UL74N22D2NpVJpfeezvX8PZy+zwh1UeM
e5Z6m+inT6/cCs85Hg8NRkS+Flr+p9QYqpJk4q5FwS2NXLCQz2OHsonQfv57WHPC
A+QjkBqSTUhl0GtnVNK8eJYLL1b+40oR0eyHbIRpVyO2ri9KafV2XO337qP5MuDa
Nui6e2BbjmwTLIywn+HFRf4nPyUa4runnrEptPi2T5Ip6sQnOUFTVffH6jAAH/Ih
1dDP7p6pkmCqcF3eEMurfZblV0fSH5SaJOFC5O7dfeYtSp+x51Rel0WTj87B5hN2
vskupNxqi0BiM34j5bfQA5XSdXlZm6ovrx/xgMrFmrT/edp79dMVFgDjVpqAJz/U
gxczhLZ7QEi7ZNQvMmg8dmMctITTpfDMne1JWOn9+tP1qXsGwSs2OZ+JiuxEg0Qw
JDt/nkDdsJ4ZEeS3NpN/xEHZ64NwJ/nvmUD3wj0NccEfWFVbox1CsTyXNBifSBZI
FVDzefb+sTTG3xz6wjTSvJkTvfTQ2m4gozvTqjPtaviDGwsCigPgYcF/qSjLf/z1
dkioJ/2Reidj/6HsLw6AfuHvHCEbtkAeZYUeUgja5OtK/6/1oyKQgXT8Mz+KfRcA
Pr9gscgQAkc5AN+9oIchLL0GKAUBde3fzU/c+wTJu2IAIxF71AMb+FG9qPsNygmE
fic7sx++UefkhMCunH0dOqPjPsR/cpFhzGhXROzWQ6il7S6MyF2IRK92ys1Ju91C
9n+qb8OWN9It4LI12cJ7uAacrTBFc+074tCzdzOoP00thVmHXtdJlfcR8wTi1HMY
l27XQEZoXfSmdOgCLOeawKvfiEYrTzw7Rau1e0SWAjqjKPWdugfv3psgN1zfXMSF
tnCxNXPLSRHPAvpz99ESaosl4n7lJXHCtaOphCLWtZqlqBVuiBC1IBBUdWNpSML4
kvSl/KhQEfU67oMMcgBHS3srQ52IPzKsuKJdeVLnRmZNGYpcAClQ19ofDJreQDge
tNDEKb44Y16CaQJj8NJK7VkfEpCTwKPTrswyltwvNmV+4u07BZ1faAMgCrc5D4jE
/8ddy1CAG60KyYqhp9agFUl9NewiD0wSM0SPJoMx8sP9AVJ1UbF6cKPHV34Vlw4F
hy2tahNoy6NxgDGYxlvv2DzkCxPUTRW/5nnp9COQ8GwJ4OF0fTlJwUsXiJUaoWlL
c73oMhayjs4JekzKRTJ7I+uzlnW0RMvbkLTlccSiwo0CeDv5MHWjh1V3sdKxn3Et
8qbiSWU+9h4tqOeDx6dKKcRQBJiVU6AMWP2kUBVhbqknPo2cZx3+1yjCPLtmwXtX
k2tA9hZEyxc5bVQ8NfpuVsDG+WFG3RgpecibT/bI4GvXdT4a4dhoCaoUGLMGz7+w
qNx6StRke1wbgAk0JdAVXwFDxKvolB3rCscxuW5rz3EJXcuGiLxHFSzmmoijRvN8
NvomMizcYZ4lRZhSKtyV2Td8LmX+oTgTFUwYHuvOnAWRGZDNmOFte0u4o5seE5NC
rKYe51T9MeG6jNUYyo86iqrwR0istyQvqPEIvucAZMfLnMd+2p5ODjeMNbBd3rPj
Nn9C5ocX6jH+UBlpV66q1XXXrkONrs1ozp/ps62zm7KmJvAqcXwHGhjNgKYzoH3V
v6BnAfHGQIOGSDynnCFxhcLA73mpi8cufMxRk5hT+X1dcNKKvxtuYcPm8/HyJHAR
sIU3vVqadhsv+Zdxe3SRg9lotclOPIuNU5w0NPO1bqJlsShvKbQ+VKmPUcgnAmnX
4HzLKnwOk/Xsl0YpjEZRBpjKdF5V/hDG7DGzKxH8VE7wEW8gIy4AGys9PK8ofX8W
8yaT9qo/nzyAQVScGdvRtR+efVe/c4FidYulTP4mfjWduDBE6vx4K2mEzCgvjKO2
T39UkvA+so/eTz8FwenBjvpBOFgVi+d5jWJSuTrstfYCk3Scg6vWCIczmX6b2gDq
TAteZwtUYsQq/albmCPfAFNbuT5WDq9caDJPt+bX4EGky9axm2TDZ9M/lSdwlRIV
w/pF0gtvy70ViJTJaTNILjcYTbJY5ZHVgnleIZBA7OZHJbCZGWPhpy8j5JX68cN1
RnzySDSLcl5bmRh1uF8UjgozAcd9/vMCjSJtsQE90QaE2lk7TObazvfgHlQfwRzt
srRsFvBtkB+/jX4Y3C2MqyC0+MJu882xSyEHLR40RT5LFOngH99JC2TNy0cHLIm5
JYlnO5dssHtcPTv+hiEJGFgh25WWXsPFv/x7bDL1oRITO6Ca2yYiYI8xCsL8hD0O
jDDlGNfK9ycaZdvXh34wlPOyvPU0CRuMZ1s9Y8oMvIAWg5+CaIFrfzGYstr1nUMj
czQiTOEf4HPmd6Ksw/h4JVQwvm92LpJ57dfmemtOBlPsiYvu3SoFGFr85MJ2LOHh
7PHJUUqS9iofcaQzFS/FekXewX3EdSOy9fHxYnKSeP5crDkOBHeg63QLkZoxpYaB
vtOGbtD3i6nPLP/yHjs41Mk9KXAVYcEh/Abyk5PH28tUOwW93PFAGyuxKZ5ppJBx
TxvjLdT33X9RVuDMdJU4OutLceGiEKidUzruDDbLXdgD7LkNL1PxfOoWF7XRQpnK
eg8zD0BnhHW8DWSK0UH6SuZBbGeLfe+r3ubCOsp2IvEeOYBT59Hd5dySOByO3qbE
w5gMkSUt+RQBI1kdTEeOcXed5JQaYhgOXXOSsD8LjMvtN07+J/6wBKMzv7JQGHsd
/zWflHic+MdC8TXIDuDYfroQfkLzwoqEUBoRPuyuzORpJpNe+ZHN97N8p0/SBSwe
Yl85Z4RiP0wE82UVEBHTnBu5IdUBsfp0u5FTRXu1J0ENGxVdzYdCeWP4TVRyhEOx
NCBWnmJo5FN4AWfXFShzwI/whm/dZ0eP+7d2koeWuPk0Jr2Y1jTkYUd8Uv9/pBHA
K3t6CzlmFCE3PHB9CaoGZ/ir/tjG3fLlGAaflUBSE1J+CvdCV24h1Mj4t9TqiIyC
xmSpMD46K4CwuvPPEOHkbIaATwNW1BUaFwyQBCshXstU14YKEBY1QfgUTinXcj9Z
H8odspLnhhbTtImh2MeHmPTDauC4Vtt4UDBYMqSCTbRD+AlLOSPlAaLV/xHEdYaY
nAwBeQ/25CejrJD//4i8pyPQPH1kR5Nh08CUSuZ+xPiCAGsbTgFKzXclqdYsqTGj
XjWx6/2g41bijwS8f7Cj54XtHZXPMXQHUswSP8jHUnDGCK8tpD5OkivDu8/Egd7+
tQjT5qp3z8EKJA1WLlclnu5KIN3D+6Ps+Tx46FzE30vDIkDfvFl9Y44zKPbY2kBI
WfQv6q6L5XV/zhkXyRSXNFixhdFsFfeoyE5GRh0y9Qy4R8OSpYdk9g6mnJ90kq6k
8+9BhU3vW1QTSVvjY88kO8AJl5pO5lPsDzZfIQmiD9ElIwqa1U+BrVP8TBwh4flF
SsI7q0t4cco0l8Ils/o5yYCMZle9ynzSeFR53ECDqB7msSjv1UNOsosQMv7qts1D
jdeFY80EbIyM9SX1m1bDtdv7U9ojuBXV6c3aIWgQ79YEl26e5BX+ZhOJER+AcxoL
iFEnbjFLYtWOz4gWvnHHrIUL3F0cPl1vZoYT5M9xMQ+hd6gN3P96voQOgDRCRgmQ
gXV70YRCoezYTy8JTsrdVyPl5510wj2J6uu7sw51F2Ff0rNcM8xzS66bNVon8gKs
EvQydee44UQB2VahpUrQJlAxxud9yBMEV0YpSCT9XZAQwCOXYel8+87jC5Mhb1md
COGOowHa1ulhG1LhuvhkehYsOmLBiCglLP0F7yhfbqcUWy36rTSF9iJpLwbVUGqa
d3fEWPWZWMKscTOFyRMw9iLhIr6XNVVTUaSbw8rg939XEvlm5nvRgu9hboUUW7wH
EGrf9hfqamZdSBzTyKc+0PWXCR7QFcx8syYku0zrBi9XXR+OZkfQWEgmA+0cMk/F
5J2zThG6GH/9jC/phC42VhjeoB0YnA/BXYBueVJBZWYALcrtWEAXB8TVETf2gaNo
uUwthDKyNRntO9lF526ZDkQdDrqio+GOsZdEdLKhIJ9G7Xzd92bFrEKXcVgYQfvM
O/Z3R86IjNnD74l4t2vTwC3zqJRZkdqUzSMAOeBi8O71Mch3YIy9SwN7MYHP9f89
OZYfnVjrYQIc34ZH1Vb3NyTcwtfOTYOOx4wLgy8IUrmH2pn/SoVUh+mCo7SjlFXj
EIPzJslUcNRRq8QseWXuFuSWgNOt3Msmp8sNd9jbiz8KUoySheDcHy1GQpWu3nqQ
0XvnSahAzAAx7Qmn2f2ZtlbYmpHQQ4ilGuR+YX11e2eeNeNhOI0SEiW19KizA2bu
ce1vSaEZu50iwnVGZYkaXgP5b9p4oajl/qlnkZ49KZ5iv+hRFKWn2Ihwgb+fBlY2
k/LL+9f8lDfghCQbJL9qLqg6K1h4GxcizJwwo5jr81nYAd7awFJZSAYlEH19Y4Ib
r3uDX3m+GZWHc5jXHT1Yzf5b+4DxK3hdRVZxDTfGaN6XC+yfNRALP1DCKxTpR9Ak
sRlW3adj8YngoMppuWdxXzYvu6SUUFTX+WBPJ9S0hcgkm7m4BxIReKFanTHiD/5q
80MUlF6JyrDsKVcQ0qOME4n73GU4YVed8hiRQXAMvFKk6PbVWg1jnlNxQ2N5GG+C
DEjU/0LiYR+Zs0TiHFuv2b4O99mj8Q2q6MLaa2pOPhzX5shPimsAd22yWh9QCwfr
aqT7j0IWQJmaMAmRc8DWYaW2aU+bkP4c/CENEsPe8qZ5h/L1rcXlle95RAK++mY6
uE6vFEUD66IhLjDLetd+hBCUPz9IW0MMXcoUcjc2gKCjEH5HGQUZgOPpt0AfaXRf
WYkQ1oeTutgy7O7TmPy0IF4722zlzvPE2M+dWNi6EqYW+KmLLhwg/1EwBPKdn9JV
7bmtzyKaJ+CidrMY21KRLYmaUgIYZywY2q/5iFdolkY967oL9WPwrTsmDdD5YTKr
lgIlVFjOmPzAatXU1Y7VuxRt9rE+MoVskXx6p2wacmCROqOHdob2YN+sjT9M5Wv0
XkJIihPAsGy4r4AJvOsenR/R+I8Jy/ruEkG5/zW3zLclS9FtsCbDXRjpsujDmz/c
1WpbWjZwb6K8sxoKxRCObkl9VImrE/sebu95QyAK/PZVt/97Ci2lCb+s7Bekwv6S
86b4XCDxRM80KqvWD65lrEL6yxii9IuJTiYhsf5G93tCtp/YAJ3y/LgHu94U/pdm
jqzR5P/5D+ldBQHYyV1L7DJgt56uaVcz1EqbCi+gGQvFxMhszNk5yGkESNKaTsCp
ODyUUWJ+PXpnujrhZ7PWfTUR9GwWVAo6MA/XAKMUhsQxDibp/v4c6yi+kTT6ZWuU
3Jk7YrVJV9+Sy6dWB/LpPLxba1e+z8p8peda5m3mUUgBHep326FevdhqPSRX4YBw
ufptTxXR1+WKpTK5feUBptQ084ecsAAFTS+FltOBlh3M89HjyH7qtFhTfSro7MyW
1kfNs++6X7dRz0BAUGGmfzFHX3H1gJrY/rH98SV4+0kbSlrvXOzHS38A+lGTKcFf
eTQ094guyHy+CcgYCDc7F22sjzrGiXy8hylbZMcM7J3fvH4B0go7mAMnCMD53OZQ
EWUfW8LC/cqyaX2onmDcj62svQs3IRNrmCTg7tccJLvbe6+TunVBOOWOIcbvTkol
Er8Qlo8IsyVcgOOc7hFx3EASm9X4kQ5dkELnu4qblJL8jMwhyG3uy1x7U31QG6tT
JaBg0xPiwf4ld0aNhVVm4F3uWsystH8bbkI/ZXDZ/BimGVZ/QnUJ0HPOBKFb4ZjW
mNMVckOyfwLMV+rB0fh/dsa9X7Ze2B9ch07NuLBvyZw/OfBze6q+PXHNTC3l6DDD
92lk/r5uwcL6v++1HOPaaVweWRrSnhvXILIn35Ly9MKVlX8+mUyUz4SCZWRqdrI9
PoC1zrUnYgaarvx28fpiuDjMYgFdIYHDNIgsGnVEG5ac/sNyFd2dPRmw3KtBQJlR
+xyx4PDU9C8WXG+Z9ZttXH4c7cx4+yMTGv7QsjJXXJfJQaXCtBlOh98GL7rpuevW
XGY20buJQFynStY/eDsFUrIrTMi5DTe2s+JUrY51eBnyx7GZDmVXBaTJmIT6R57O
Me5vRbQECL5mN4nCwG1ObpMiO2bIcwUwx9VFRN3RZay6aIrmZR3i04tBQtNB07PM
RUgPhcA0sAkIL1a5PuCAS8CZ9/2/Wg92DPYe2jEbA6SZr1aI2R9hIyzv8xkv9OzY
bgdgGkonakj7teta5hG3U3HE/QOK7W3mac60mKvuqTdL2JqtAHiX4uyjyTyHlejx
1fdgU9YlRc5YYtSrHe2zr3C96aIWFYlQBbcYqI7DqupeHQ1+5UxQqBlq9akVIRVz
eooe3FfaJH8Eh60a8wMC3+/FCWkprf5ck/cxB7BAGQMkfKVQYUlN2VwoFfXjk9tK
Ttl42iDfjf0t86GeJk0sU4gsbt3C0ujsHzP/ASKKAyqAmSvPwnqqM44NStmIdjnE
mIs8xRPXEbXOOdZIYh9f4Isy2/GTzB1BfLxvCkLtuU/LVES5XsrxVOoat1oo5mtn
qXHcNVRhcudOq6lSyaOJNiDoQhPTK5yW/Yl+vQ570n2Tn5yu1QN8g5ujjZQopiMA
aiIu6ubq0Om9ZDq7HVzUgL5BAlNusKxLRXfEw1Cx6rBJ0lDlxTHKFR9Qp/gAccvQ
DGubotoHt2yR9cGOUoRUGQpmk8FPulGbugVR4LKvTnUnCkvJV3f2YPZmOM0ZmhPq
K5x43MZdbXs4Cg3BxVPKnGVDiLjU4qYeOYUJqdNK2+Kts7zMuXPH2jo3N5M9voN8
ZydciSP//V/hHWV4tVY1LwvPVYHuS4vw8fWVZXqwtFFufgPnr0GxcMeeW/yW8BDJ
4ELgOnNxxKv1RViAJ8vmjxtMZz57q5wlZBIiNpGt9YC5LeZSTpJvBjna/hT69A9K
TrD1GJ77VCxQ1Xknz45Be7Hij5i46ofLZm4GfpI0A7dDYtA6D5TTzxxD0VvL5PKk
YHtz4NZHudnj96naTZsQPBUEkzefU0bjlNQkFEjvLnWAeUhs6NccgBqeaBUQLZ00
G4UDZ+qBj+Y7wuqNdYznCZLoyvg0YhFpMtl+nwtv/kzagm6tUTalHwukV1p3a5JJ
Z+06YaEipNqItgAAK4z4ZAHyelYSl5rkj2oCIuh9c3Q2bPo9m47KmGdRrTNMCd4M
CnsxqCQ+dznttMHRyNsJd5jCkfS4lbAhhNG5qrsbX/IubROvqidpnilHrliM6V3X
XeIvKmomTDh4YPWRghJQdb87hiVOdtmCOs1upxLHHvd+F60NHbyv1np0uR6xrtOo
sDm7JqRFZPTlbx7CKSRLi5Xeqn1AMLtZ1orFemsscRf5LDCrZVkaKuj1K41857Ge
gGfRVZnOfYQ6rAhDWYxh92if63O6dq0Zd9bz8MYAo/id8HLKPpjuiLE+kF87DawS
BKTRwmCRPUkK/KCxD3Os7DNAVwZajiHyCKIeWdJ4k+5grlDPXN14GgTWb/WPpeyJ
1NEcZd+xHecaFhhadDRj1SKVk3paWq8l7yZZcvfDsgJA/EprvsCMmLep16CcBYYS
DPjCg7n+nYuFcjY9rv9XJAMcGt39UyR9p4DdpjVSkvXRP7xsU9s898yuIAGvx2q0
xZE5TYUqjKEwl5FNEKfFe5zeoP6dkBPgYQYEVFDHIdRxqaAAhY6noa4nx1e29VQ6
T9/wUvXATKClQtLVZ449sdHbJwb+YpRhIkrUFqfAN1wFgVvijCbBIJqbKLC/rjZX
SEwYem+ewkbM97USYVXdUHifGEKv/S8aG+M17ywhfks8lcCvaFWveQpp8TDf4DHd
kTOZZEWnPKK8ZikyzGIY0AU2St73KhMV/G6Q+5PYgvPIMqnXhEWLdLMUB7a0NMtu
2ks9o4HpBL2PIRhNM4dxI2pqarUWcLcLwzWgY036ilItGh7fmaEZQTDN3XnrAp94
sTCMlOXTn8+vdxekJDtvG3FiD7XejTh1PCkR4bW6eChRvApIaO56x3kiHUudlhuJ
71WdtmBBB8GkoBGJ2UN8gv+KinZB2PBjdM8HevNggsQ6SARlijR019XeFkI7YYVp
5/u0bs5ZLJpb5QSNohHbeMw6bssv3rBSUpD8GoSsQ5bZZArDeUH2TJ7Clg9M5Jvy
Rv0YgtrrmSSU9YEILd4558jR6YI3IErQ7zzOn1rCsXkHfxZLuJPCF9rLxlv52TTZ
lIlf31EKgJBSWfy5Db+TBiKiberG2kYQ2RopUZSHGw+7SJPomZgMxnoquDL+LtR+
l6k8ecEL9O1vmGdWqF899lBavFl4bXNRNowmIKN9NUWo3620nFDCS8Mc8AuiG4Jw
2o9ovVqlUoD6DWyWdsinplI0GjnmxTtHaT3MuiEd7iZs4C8zEzXd3r7jNFaKTftI
ZDCK7U3l+sppz6yVlART94whYOJR/J3d1agLrTFTjNUawp0269u4FJqYjualSVm8
e00Zqra0k/sOStWol9xdRo05/aVrWxvwW/UAL5e7GMBYOtQj0g9hnjjHSBQlW1/I
dP87Qiw5qGSftp6n0Ycau94nH9pvi9JIFy4m368io16aSWtPQuxKKmnEdoMCpUv7
EVMeOQvbYeEC0JkwOaPzozYoHT/Cg1oEQWT2YO/EYCLzHb4ffRZEWE/r8X7fqLNJ
oVe8AHAhqOT7M91jwzm3uO62nhHF6clkQpIZl2MfLA8PQjnk6sVBioqbrIarApMt
GkEAI9yg2fwFoVvQZWyy3/kzDVLuPlMZ0Lbk9bQMeVItmX43vAC1A7CV42LEh9hu
Ym9RlYtQ/U8fruBINyPIGb4Hsj3LwKBGRrCwItVBP/7vCtfOZrBR5bQ5tvmu7Sbg
+RjYE/Y46vgp8gqyAisYHIoVrg+8+Yjn3eKiihXaXjgYlp8oK35jqOESPo8LJ/O2
b8XNcwlc7EryuhC2ogiOedqVTwghy9nvnKf2EKOLE6L1z2l0wSR8jdoB0POkqYd1
WjePc454T+sDQZpLzy7wfm+VW7tVY0BY5BHgkTIc+E7l8a3Vk1uqFHbVVZVO4imN
hWvjXyIJcmn8CzKWhJWZTn6br1s+7qhc+Gy0/HgiVPDVvJ6yD4QDG2AXU77ntJkg
FObe/SQc0pE192qFJgV1IkhGcdxBQyy9F5ZB0d/0NzfOMAU9hjr1YpKLEkyzbPv7
j3elL6pGb6YE4LRpmw3/Qa+b0UJkYWjV+2fa1Wb0LRrPOVcdr0FgabMq6FiJtYCR
JFw29Zs69tQ289CATG6PYapnAzfMziLLiYz7KGvPn11MR30kvcexfUOVv1891KXx
uT6X5toMXV+2RW6zHN1dRtWrvjG0dU53zO40K+QP5I9/qMJQDWZkFP2oyItrlFzk
M0WJJFz2q31mMlHf2TImmWzH3GwF/cde164pfNySI5IS3lNVdRWpUopSBf1uigch
CXox03UyksztKO/2qc23AQrCMzrv5RI03drkEuws8KQseWqDHUlt9lU3H3/4q4UT
skDDYcVQh0QHBntB1zz8gF/XASOOW4bsU0PtEOvt0w48PUgOU5DcuCX0CzoHjyzs
BrQ2tN5zs6H1g7EWJzjQh3elNFRRdyyPdwrkmKYqCPV15VvpHjbWJah6EZbkTdaN
7gYMtPykzMrrE4l/KKIuiLjTdAIr4bi+6wtfSU8A8YRC9ax5yv3hh8uz6ALdiiYo
ZnEq1W4sP4ZzB4gk5jRQrb1KoO9CcOwCTDUMBZlShO+ZIVI2N0u+nX94vwHPNDBx
JRtqxtjxTJazN6czAkZQWDS1s6ENRaN3H/8Q+nL4fhtsjujSbzicSLHjgC3HJbnY
xazVWfxP+btvZeA47nUD38HIkJLsxgqXuKtl3pOaSgy6kQzSkoY0YWsEtWrdJIWT
+UcmeOlB/JjKxkRAqhGDnEO8BTxexqIFS6ZQCCwOFZTcwSlIpl8GhydIDCrG2iJP
V+k5Q+jJzIJ88jd6er7uffqLr+TEuLG2Jd6o2brvXoJyEYgWu35W9M6QLCs9H1V9
6Sfkg3mPBPjjM6zb1KjWTttXQq2ToZGbZMpPMxukd9rdYJ08PeKa5ELhChWm+0ee
p4eyQCzv2ue7GCYB9t1wLABfJzNxJzhDZr9YS3zqbXcbDlacRoV9/2vFKz/wVJfQ
RLWHa7FMvTdMFypPtSWx7K5HBr1DbooTYQrXZsgt3HbLuL+2cif997Z4EYDlVA2W
8Q1w/aHJ52OJH13IZXCyIEkmZRRj7iE0G1qI2kssHRhqsUbDrvoYytSSJa7MQw7W
LpFZ6JzYInDI72qGTJ72nAJQoOKCwGN5Hs+1fB7BzBxrE9+oEoIVkdxd1yzzInBV
Goyr+alngSK7e6z4/bWyHd4sxD/5FVextOIu4YVIyTk/so/zgRDNybGpqX/u6haz
SoELKKP/v+NB7St9LJxblPMOCeK2el2AcGfVakMjx8mBLS0dEQWeqIPxNITIBbJL
Zwq3Uhw/WhHEhnAMxUWCiQykWFQQw9xq8srdwe5n6e+IABieQxMHKtH2r3G2K0bI
nGHRldfsMzqwAmQYeULToXRLoA4qyuD5ULHcCYcFOkf36x53PHOD0xbbEouJ13S0
ek5GoWh8G/ZXMV1w6yPet82HCEAXX8dtVvTGbLQc2wupkGJhNTPtT1gy4mqVpUVh
eKewitO12ZxI3+nB2p5ruHGhUOmh9AqqAdzuScIzCfgjvmzUG610KQo72xO5rbd9
xCC3YgBiJax0KBMlUSSwbJPtJrBnVvPSV2yaEIaVtHe1iNY+qyprY1mDRdwAs7Uk
inu80n1Yaw8u38wwJouCRFDe89pOFjk6qVVkbwg81IotdOOncUOYOW+fJNAGIRBV
V3aol0+rdI5OR9raeb3GzHqcWBKH9aHZOA3ZQndHwV0Fzz2nABjYwnZZn9ZpADTU
mCt1Ij4alnRqzZ8p/lfzspLUTA0vPOJSOOgow2Msys5ILDyS3yynmDNgW/OZvdHs
sS2w8q89DUTaA7GQz8sJDo18nsDbQXZwiq5tKo4EWpWmqw2cxP//9jkGOlkknWF7
UjaIaXFZtUbK97L433beqKg5AoWp4LnT8YFTCYUqLrdVY8JNhuKfAWlBDQXT0J6D
x6L3a5Bmfubu5c6xz5Q8OGUjUQhrECS0PAVKJOjxIJXrbPRRcH8woNoI4A3KyLV7
sTovV4GZW0SJmjAkjEg2dqsIZ3Zet7yfqUpHgszHXFq1GwC4RSEo2jRyT4kQoV/s
Y4NT8UlKzPSUOLUqNaoocZU861/F1bsW6rzP7lKc82zX9BSxvorseTl2HsLO+d3y
a5IiRmFTXuIOMv6w8ebdndfUZaes1SN4cxEaVvEf+ziDHVPlMgyZphbzZvj3zlwX
QoBeZUDUIyPmL3qZEdXpynp9nhAcHROUyuFMJ3eZXjYOYO97xE8dcb8b+liy8jHi
zSEE4GPjFbElgeqpjBSGX7mOdIc5HtcE1p0jEQ8z9go73BMwzTP2fL0oZAvSSUSA
ibtED2EQ2YRmalMrteOAcgMEe+6mR1sgFyr6LkzIRCk1maOfySI89d8S7bcU3/tR
EqN1S4opb2bpsknpv2Ng0KIyDiOlMpJU86z7/3ehCRTLuKR4pNTaIwadL0lJwQP5
FDvR1sCxWoPtLrem07XeOtuWo1bh6Rkw4l9DqsFdSZhAOXn5wKM9Bj317GS88mwx
oxe5bJ18waDsKDdOWZXfwWJH6RxOQEmex3a1ByAzSFxHJ4zNg4ZanCx2CoVB27dx
wTO0Buch+YSy8PdTNPQ2CqP6LZu/jpDjQezBpBocGWy5OwB5OhTqZDAKDvilES7w
u+tQhTVfZX8S6vwJFrLTjLqLkKtvXgHt2BmJBQTxiAH3HxXXWMnpj95PKTPNPbpo
djJUW4DNsYnt+JtZDp+KmPFmJLaVRMj/ZvkXOK7q9qG/4ZstD0U0FIVVLadD6/Er
t16N4po+6Hdgmq/5yT5JfgUJvdbaIrks5yCtQ1wT69YknbtRriXUoiRsbpfe2IQ7
MOZWzVTb2bE0dDKGq+Dkm5qDlMYxiA8SBZHhjIZrmyGqtF92RUApTRid3D4NLdz9
rbZ5qlwhOxlT6KnDXgXGvAFba6hWBzibclSv7xTWhHIUW+v5wAFK+sWXBoJ4EVi2
E2DRcyotCnRzHVVW2zVzFf+JFrbg1hGUeSu32nwQ5VoyVeaOzv5KL7PaLkdBHKqs
YOR5D/uaL24+uOdkQtrdRVi58y7Yd3aMBLkFU20OWeJ52wjvhTOw6M071g5KXeg/
lqaN7HfvarESL6qSAhJC6FbeA/cFHU4W40oZx3MfKqyrwMnARr2VqJ0Ak/GPVQLH
PVjJvP5JNIqeuL0nVMkdyMIevk06Mj8yE0/gd/bAJSPXaKsNBm7wGObN9LmN40Dq
nlu36jfIA/uFmgj6CUCGHFLFm2GZ9yzbruwsulQ0k1IWifyYhh/Y2H9c1HJvedn/
zl1vepSzjts/ElUseqc5uSrk9zzvmySxUAhNaSEy0spE31SWDKQIFtWM6rSizpie
4FJNrUak0nyqo3pQGoqRTFbD8Rn8OILgS/R042lbjZGEMnmhMZY+CGZBOyxY43n6
TvlHVVOedG6GwAog6cJMnFFgo7S0E+MQxGpN7U42J8Ojl2md+2gpaRvUAfPo8j4S
3CH+Bbd5VE1ZwDknIxYq/ukZKSAjpRYOFOijMJpw34tpdfr1p47RsHlkZq42ima7
TwBGttzK13RvtL1HxFsFGMoXizp+BzsiawMi/6saX9VACIfCI/Njcp3TNUovJIAz
AiPmGopkiIDPq7AjwP9E1ssTnqxcbJjImv3NpRccQw7i3bSRHjmiqf33wwQN5UeI
bPGNwFe4sPTctkT9eN3eZPYltvFmwTC+TGD4BZGfZH6u/QkpG5qakMPTDQyqeW5H
KjgJkWFpmBU9T+4qN+FHIrelQiItXnc44N17Zi8u9N9uAWOWKBQivNrtsbtqdPYy
JrKK0TFLUOkqj/fmdcGOGrmwx0OA7AVI4e3JlnHPz/+ZjZDz3xi0EKOzfQek6dYv
SM6OKfUKi8I0GsFfuJKI3iv5lXh9+3xf1PV7R47AfcbYSftMupVf/mROsEbt31FQ
YkAt43641Ax7UqrM9j8egBeXorgwEzgHiprBnDfnsg445i/ByzkHWNcMySdpOHHT
OaR1xbaYvOdi0sbUaEkGOlg9/On/gUcb5dY1JBK5AxCTIFLIJRJLhSc32bH4dg06
PnnyswiKBt6MZC83sDhzoERCITeXxHhsyMpnoPkeU+I7KSJFMwkXc6xxcPTxK53W
e5qX/esMm71DNqMDppCe+zxiItPUUIi+lsOx1p8lxeb3iU0AYSD3YmioFJ9vohBc
s98QCT8MWA40ysW9gnMHlEX9wKjusbBu1nxO+7bI3G1F+yP5awczCmiWyzXMuOBZ
d3RDzHR25oAqalp1f7aWnRg4eYlTibJUrERy7Q7IY6D/rB2T4NB4h3YmncbUqeY1
79HZ2Ui0pQHCD8CLFj0sBM/bdr8bziClL36q7I8NRluNZj38ZU1sY8h2iQGTRiRF
jjsrVjrmW6/7drNEiOPVkpfxU8OagWJsrVOJsXOLQnXSv9ZkjMDgT6lSKeMBYZxg
yWqpAgaq/CLSRMvGVh4nUY5aF/hk2IGkvA/aAjz0I96oGZX8HXiKV9zXVVv1BPfJ
bHZMlI75OPwMuTgdrIP1dW9YJurswZdf6KcWcBbx+3z86IaLNkIACSeEOPKg6XAI
O7dofDXZdEvs0Pqib+B0AWlUmo0BJ/RFW+ULith8ts6wYwSRfwMNv5dHdNdlCkRi
USTp9fZxT73Za/LNIIOycQVJ1oAOEDn7HGQed6+TQitkHX9osngZDkMlFlbOuwgl
rf3Y+Jwdw7M5lZRSaKj54/zLC4WC8Ywdn6xv0d9XcuCK2WmP4akmom6QVbUDRYz0
ohemXSWtOF5xLp/4bj2RZ/K7hg3KU1vpAuoyeOBiO/Kc/7guB7a1vr1Du3FYP7Zd
V0a84JNi2KTw5sh0v7CuQqASMiojjoL8DrFZnzs5tiA2aZop6BJiak6hj2yxtqo6
NvHgWOSPEW6GlTM8mdrsmtQsrUKsNq0zndydqOQodtrLyOK16XYKUUnSpSM67XMm
PqOxHbViGei9M+2vkXA+fBW9iwFpujKfgKcXADFCQnS1CAw9dNivp8SzabktXHbE
GNfw2jE0jdr1UWCOyFkrR7iQAt28a8V8DJ+7f9QFaJFNlhtkpXkVEOrH4YcsSd/r
E6FdLt1/X4am1DsG6fKm3aB3LRn1n+5DNJp+BO2f2QuBMQw32jrevy/T2zqah8lb
CfwiwrxsWl9LnvJ+3eNcJx+qyZDW49gGTt7o3/+QO6c9KepIRykObYUekMx0F0AU
JoxKQFd5Xt341ZbrajEs5G4nvI9gI4YK1oFiVnK52mUwHKIkIxWmjdnrxtEFh5vx
fovcg7RVco6W1hXj7XIs2OlSXlo9W8Igmhf+jUkkuSeRDYz3vfxJk8IVWVotBHMw
bYIgKRI+4cfgatG233F2XO6l3YL1vPGwcgwTXSMq0w55NmynZfWCylG8eS5S1ys5
MpBuvTLNGCdc+PsD/rWoCd1jXelSdiTKhcXWLqoRb0QnSGZ1Co2C9XU36xCtCTc1
YhJx82UKmfRRo6CoP/kdskAayIL38xlBkX47sDCNWMvXpU0SQzoM5Bvw2+dZnZcZ
MqHfaboWol+G7Rzr7+jKpu/I2Ugof4LxmVRCx88LzyfkNCVrHEnu0trpUVRhaHYu
Ei9wibVmNEQGDPjrxuEmSEekFzgXekuCMRNwM2BefABag4RsSFizVwMNDrWMga3V
STpQ+s3wvFVvKIYyjaacWxQ/E89cQWkl4GNelzSWIQIFYrajwsjd2cLqFZiYfWAu
bAIU2az4n9WB4jlpD/VKmM8S6z9Cjj/Z7D00W6F0hY2GNQHEHgpTq4eqpejdg1jf
rdJRkDxUsE1vWS8Gl8KXN7hzsqQQCpftP9WrFIip0byd73Ty1uJ9nYCNznZRE5hh
Ik36B0b1lh1gUUs90L7mUTgiquAT0SrFpk9BICm9MUUBq6/DQB1uZnCIG2UhXkfp
LGlwmx7rcX353Ua+EMWVY/QnDn1H5Fd9c3IyNJ/Miy5R5JpGaqE8eLpLFPzvMGQP
akAwGVoS8DiRK5bn6WJgMR1YxNrSG2LCHhXXhIfQyY6OTTQgROkUa0BCD0eTbwYu
Af0hy1h1V0vSVNk2/FysWA96L6QZTjuaNBKE4BMlo38xf2l6RNGfYcQYfi1XIWAC
q8PLaWrf/SdLPgy7bcKUaiCEVvaA8SxxN6S6Q6rKR7a4tCCK+vZ3pOA5YRAdxA5S
xLnNrcFnRmE0E7mOQQV+ISMvRtOVQhQGlBCbNSWTRnreQNKstvfWdSvxSLSa/mKB
Vqhn9va7k3e+/1siugrvqO5MJ4P/F3Pq/uVm5nMIi3GYtlGwftGJ1H8SIoBGYvlK
5bcMtpWozsJKXzwSSOB3q9voDAWO+1/04lS7IMM1QP4pfBf9OEMl2x0AqouElU9D
YEYaWQf0+ZK5gCcKedbIhIPS+AuqBKi1j0H2kEB5//mI/GMbRV2rjuFSoltaQOnQ
dD5NXD0woXycjWAwt6Umk4U0kgwnwUy1IS/5qWOYL2aj/V5ruGLsA7fgUQDLvqZ4
isqYdigxx6nqGEl9rSs7hdsnHjTCKEZd49BF9UCfTExdd9RHLKU3mT4UeO3Xiuyj
80+NkSByXf23fQN+5IW55z24v7k3QZSG+pxSwqSHWElumlYgD8gdq4zDCO85YUZC
u2x2v8oh3gJz4xbf9/dVCd/AY9Ht6YDPOjIa1RpUENd7hlvWM5S2ISkYE8ngk5o+
w/IdoJ+sfzI6OHFDTSKjREIIgk7kR575M1hGK0iFgI4DozmVTb25nBPpS7hzP5MI
gU6S3QZZZznmaxOrcmJey2NI7TZ5ob/chF2kY0GhvHdftNVqxeNqkRKX3fTyJ0Aw
MmuBJAG46h8muEcRYnPgAsA8GdIcXeH0KdF6DZ31GaOATlqanG92yvfocqxJByq8
oUUv9P0CR2wmR21zRZowi3gn9nxTC1uY/kxERpqCLvj5Ec6CrUESaeUZU3sYwKnT
eXeUURTu3XrTMa97RmSAYCV5aBZwuzjK9WNFGSKq33nPGvEzXVITZZ6qnTz+IS+Z
aF1UBnMYj9tqiOTGwZuL6Z9qePlq/Jiy2m8jqlzNieEQlx6Nrbot89ghIXphklh+
yAMdLzt5g+0xABeY5SwjIgA73dl7REpJ+ZvBdQ/jdmX4HoF3Gj0z2w4PQGPHsET5
CTCGa7PcjqYFjVl7skeiGnM3kiOhXNcM0W1Ugl1WA0etI2Cmv+092JlIFYb7gVA9
Q2Phx95sFIbVYlgzmsCgh6A1zIHpTrJlZQTohIG/Tltt9lyfGJLLcF1ZIbUP7hZq
hczH6l1gNPz12AOoxyCN1H2GvmlPlPHcUWP0Nc/k0xarRsIXEKWNFF6O/GLPzlti
4AUUsEvNxB2nzPhj3AJkU6iXfXdXPAheufF0zBpxx2lcp6v41aIlVyd20vTlf2hk
9PbChZZqL/+QWaYd45sfrw5b1bsp5C57HI11E/+jLfcM5L+7As+zkExy7QLE7GiI
SRed0BOLeOIds9hm10aTwI8AYTih0kR2nKKDp7syjmPfjdOUC9hGWXgfoGP0zEVI
lCsinzRkGRA48uN7EdTmo6kBNDvsHpW0MF+Q6AYctsLNWgAuvw3cX74nzRWPPbGn
UN6lqPojfw3aJrW7SCBuh+2PzVpcgJf4RMkzZbRZZvqSE8GuPpFy8PE4Bf0Ywqyt
AAjIb9lFLgBqFxRjmjzkwlGTCJnBE093gIlWQY9VjzevGlPjxQyzEZpbbKHM9DOb
qBZFIVogfse0JhpZ5mhh4KeWWJpUtd0wdYvRt1bpUnGuVACxMZWQ5dcL9NSCdoaG
Vs9TW8GsGngJORap9hdQbYWwQ7n3k/4M5Qh+WnVQSeI82bQVG55UDyXxLGF0mW8g
Spbk9BLUcLQLOHeDUnY05aOJtE1iQtdKPqcGHjbD6bPrE7uUXZ7XWqx/xbIdpzKt
MuOQkhQE1TxIFnXcYO+k+YXQO4rA9axDgBJ3EHLVWrHJ8SgylZ5aHooNn2wmLx+v
Lk6rHCzgaO0AnkZ1j6DDSmTw997XSKhgYcCmMVktsih5kNyBfplFVQPYTDwdvRn4
4v1AGj6mecBPzXXOXW1J82nnXfwvngHYYnQi8+GWs64tZj/dPe/Mj6y7z18DfDuH
1A1H/KqUW/64oZoMf5MfdcGmyFnusDBJU4tjuz1iIxlMz8uvRu+lgLCzgUHd5Chy
i/IoV9q4lez9LQz6JAAJKVPS3Pw7eRyDJkok3v6R63rFyJ0gEvXUjXwNxF+IkXop
ZXrbmQppP+Ai4LpGcoH8CtASXEczXwejJgt0TOVe6k2dfhzVeqvG8AkT6NWMwVzQ
ERm21FI3uDM/JVrdL4DVRdeulZ7JzE2nPaamFwjGnokIlksZKppRJuMxYbc/BHYE
mGvyVknibp7q7A919Op9jiwp8U4j7zCbnPjqwmv6WmV55y5qiCWNxhf37IlJTHZg
i88QrClY52cMQZkq951sULvwaXF+qHAoBOTuefWHVlxJFgeMDGXPAfVdzcjM8pnU
h4TNmvaaquPIMiTw0NsqlASE2ESG66mNuSnmkRS50xZoCTPDQcBSmQl0SXkY/OLG
ZknnTlZF+cMY7/zQENhsKfWezJwbWMSWdC+7fU1dLrEam6JmYWtkjl3RPEY/IFzl
o4QPxZhc2sfnQxg27D8MD+corFKTK4yW535yY4a/xXIW9cLOTVA4Yqidsw+OTbhL
5tX/eDpeq+HQpfMOcd5zg/3kFUgrUDJ3UULTOYYvlGFfUzi3/GnuZsQk7Z+3xyfN
iE6f5X5vDB/ExT4ffXKg46xe25RDhN6pRNcMB+w+sz/GRqALUFC04tbQcUHwTCrc
SE/c7YvBqhmMpo7WaJwSrSORV4JI4H+8uazwE310MhYPW8akuRvWnn99XmdGJ1NT
SuugE3W3uaw2njnUe/FBwwcDrj7q24qRKqJS0/DI7C2W7Ijcou2ofDmP0vrgA1QY
LHmiGRBtMQxx3gRTJZkJO1+RNBRRRmwiawi1BfI5QhBg4qT2tfWIGZy3FArrv1LR
2lkwLEHC15mgkcc/YjLdR+usEIhPPlf74cOsxBfW634j1gFmgBxHvQFjukapvOuu
7AWdjNjM93BDu7jtd2FJU42YHfK/0Tr0TS7OVt3K3AmaGezO8Ajt63FC4IzfZRJN
y/hckXVkXfhQfHYhE0VY8qvMoAsZN2zA0cdQh80Xjsyo5FFv6ZIGsa+0GG7H22wB
J3J/CDdRA2fxZNddsyyK5FQRD9YXuuis/ERFAzL4quihJviq+NpI5Sd13ZYJE5E2
JwIzO5Yvrzrwd+MR8TvBNyYzRvx4BgA5rExgF0m9vgQMul51FWfXEOnCyPqIfLZE
khqfzFdzt7jbmGLbOCECJf8t6dzBrrOPfFUMiHvugCLaugQOFnI3QDrudfNqidbb
3BHLxjwO//PSOL/mkGy675FRC4SAPriM7dpA+c41vM4ZywiVX4dWan4kQ8dy412E
IZpI0cRviZY6xBxk251Ub2/AxrIu6ZI+/NDpmmXU9AleZ3Zo20EIJk08i4u6aRJw
mXlRLR8Cox461wJmBFXcHahBRnZ4wlvCLR3AketQnU0sHYv0flflCxSCnyNYwDij
eiQQ/2zRWy9t6MYeS43OlfkO/Cy56ZC+4r6+Ckp23s15iYBvOk7qoAQwaKN9NmhT
MFnSKBEO4aHdVP2YLIiu2zCpqMaI1ENthohclJe7T0vuFOuLRpRTALpFOJ4cRJbi
Mpf9tjP08w3uiCRJG0U9Q811u5ornj30sxPUdLOVchMXavIHoYi+gbdrGdj8eO4w
Zo8L0bN+G75sqRkHdyq8dqfgfL6DInW9si7Bz28JXvsjGKRnztL+BCWQkCjDaCat
VrmDaqsxGkleWSDFMbBRvlpDH6cNSIKcHJ47nvIrOUHCY2ibcHgH5oxz44RQ6p19
Izns3o2vyjJnwZ3wUM9zB7i2VOo+FCZ7q3c0BLieL9jhENWwuVf5LaL5pXDKDbwv
bKl2UoSO3YuPJ8e+H7XyEeOFm/R7k3rY9uyhhFGPZfwVszDbHp8Ri1xILBTV7huw
qTHMoeRRXbhUiJKy9tU6LH5Vc61dTuyyLl8+y3/02FMQtNLNVgOLAk2l3n0Jpx7u
zKxEE2Rb6nqde40/N5r2KvSvu7j4p8pnpqxsUVXwZ0qCQAh1wb4YcRfSbbeXGNKk
1ya/gLEuNgECopjPrM69ETqMkvYEqHr7Cse05GBN8AmhfneV1AL9GkqiXN5RWICz
olsmr9PYYg10vTy9fERjwJmlIHP7KWnJR5xTFpja2zPxJSe8GelticcZvopMydKf
ZNH6eAuPx86/jdMJmxQsz10MngfXuu4oT754WT/gWtKgW7E9EINvJIeY631ZTNWu
buvmxoVRo1b/+c9VO+VLI3UyRCgkwJKMj8VrivXZGZ5oTEu2Rw8F31bBCIkzc7zK
HSPXUfBkGhNmensLCEuaeAxSA6NKuIaVF6x3+1M9WSByx9D4jIDMBK7WGpsZJh8k
06y7snH+uHC1nAoTWyUUJ37k1Caz2ncyVR1uz/vCDNVjoctEIqz/YZFw+bs6kB3m
oNZUu3ECGYYOkMVYbEkHMO7+Sj/Hn46KmIZXiNFhxNk0GKQwftuO4+UW1WuzOBSf
PXUNa9HROSHzceiZqEWamT5z+aVDb9kXn+KmuCP1le4KHfR6zpOOGRbVKoqokJmi
VuOP1J3RqNx9CR5iTlPLdXtHXIh8KnHySGaVrHsj92/2ol/NfYVA4avqhcZf8tvM
j0wKyeK+oA7XzulXk/dCe/uedn5oN9zVFrY7KMocjd+9matlu3keCN5E7YJ3NoBU
eA1FlT0vam9bGj4BWFfP3LKl0wJAPG88ULhnOeRrGiDaJMi3d7L64gd/BB6w5a1x
9NyCln2kYJ4Pl2ADZFjdt4ZUgnZGMEDIi+qtLjGclPS0iMFoTAxLAcOgbjNWdmFt
CL8zwi2x/Tw07e3ZTPjv3tk3XI2ChNztfvajmFOSumcm3dYy0UUyDgFZsBOg/R2m
Ke+d8zmBczRSUuvvqNpwoUM/2iVgBdTIqsBKLqUJXqqOmcd8ASdPCUQ8TlXFHXao
2BFnhzqApyk0++Bn6/e6GkSyp/Iq5S0Lf2nKF++AInlIf9dY2Y16nUK39hP6Vhlx
mlu/8uBQZj8kVBCZ7mVtMXSogfGt4U/T4R9zAsyTiHIqAdP+FEFIWaiXjmjppvb6
3yxEyjGCKWWaKVN4V7Vy3jCY4HEQzqe0wMiAH67B8BToEBHK/zppO4i6MekXrpIl
ieGawu+TrAcsfzGpWH1KnVUjpDkMPs/bS3hzvxgXqIgum7Ij9Q8+w2FAoEIEm9Bk
xp8o2Bpw1jO6SLqhT8RjLq2v8rUQyNuZwKc4Dw43Jlh651FF9dnOM+F/p7jWp3/f
D6YB45yMLbPicZ+Tgo+Yci2s+jATTSoq60qtQJTYdXh5Gxj8U5aQycB5LII2c11B
Cdo6TQsR2S1xSoNtWz+AZO7Sogr0amN2SsAdX8V+FhTTjVSObch6cmPbEUDtuic8
g3ivCLBCva+R7LvE/Ex65GpyuMkO7phl8Q1wrETFIKIR9vTDBowjTJw6sKk43MQN
liKnxI4noFlpbdkZUFBePFcmm/tbKbe7JiqntkD065gd4va8WrrYcmEoIC+zCdka
LCmF51bzR/28eVY+rAzTAz01Aij6dOf2pss5hQEQ0+UZIzuACpf+tiUgYOh9UV7B
BY5nYSmAI7bmDYt4JIBWqxjzJ8/BFMZGgnCg4VItQCF7GcmWL1qili73/xv2OMfT
LzZRTVKw+7j8a/1NZy7bFbvg+FRZpAJpSXZsBYPwIwRFNhzuFgnhYT30e/hMG1ca
U1UPosV1B2S4dOGJwrzGwp9wUKK/R0uqUsV5meuoQ2S+srTVtKpesaOLzPk20ypm
WggzBgS16qkGi+dyO8e4Hj/jFbo8laKuiIy7mQJ6w7z2kzEHsfT1u+vMljTVa2oV
yHXeWkmj9jdyZ1Dzxh2LsxK7AB90lAQQhyniMfooDpZEQefTwclFIHwB79VdnOUE
zlZRSwGJVzDezUra80N9OmlTfahJUh2iCIde5xJt+vAbrxMkr0hm5eGKqcpf8QOH
JbKGBpeamFhhTtYkuzlvIXH+WiV2PZiQ4L6GhH/yAFVhSFtmuuz9InT4Csf2IzMA
avdQ5ww3JIIoqlPnye6H7i83+xJei8qN8eUCzyPK40ld8/I/+gSdFUcR6+fFAHLM
0y+8PQkFXwkZaKjI0+AZxZ+ZK6UjRfvYSh7ET9mqk4utFtMKFlR/cK3ROFimojtj
veTDCW4LfRWWDdRTOzbfNRoMB84Bi55nW+dyFMQsK4sjiY3S+aXdMAwyawtRsoyC
0T8h7X+loIHzu5kx3X3k9MCjeKGTlGsTbH5WBzIloh6KEB88EJvUQTEHdpHzgfxB
j5Z0In3F8uhL/R5q29k0SP4y040qPylTTQZiCm2mNMujILl5ummuCc2GB8/OqVb+
hcK4sXiA+Jei1kwsMw424TXnnKzn98+XZ7f5bT81pxMapCsQQ2Lel3aa+QeBqfSR
1lxe5T9VsorKynyZkmKO+ll2HMCzjeJUk39OTVaYtUAi1hT60xNJFJeDmGTWKX70
WxLGnoPps+4j51FcG6b3rfA7Mo0HjcsOAtRLHPPj2Er1630hjMTPRu7z57azOwiB
FxCRcHR2W5E2VZzw4s3f2FyKvYt95PKGC7d/wN0gWBXF3QFWYw7dQOnWjLH8Lc2o
bgzcFR8AoaWJs9OF8c/MO5MR0CN2e977Fqa2P/sq1E9WgHsr020PUB0QdK4YKKUF
xSEpw7EQCtsHe2q3ozcuxghZYh+Ul6Foa8Lu0SZbdEo/hXYhHj//4ll+viszsaIm
n7JrMgLaL/kx3nRSEOvaP2QbeXylRtMFMy4P2zOe3XQ0H8Vgg5vFX6Ri+vmsKsFy
u24NdPcaHBhHR+jWcpsJdkFozV01v1yaTONZV+kM4OuvRFGBP+10TZJEbhKzUZw6
20mdWz8FjcPsZnTxX5idF2VhTwy7MUURvz3MUStUGijDINJqOPpnFErhaWyecZw7
lIX1/xBMvGXyRpfEZQ5T14Rx/AT1rIOnJdk603U7d+vlyj+VGXsje4Oj38Pa0/4P
IIv0IRpPKE+KTy7Qk3HHTmMLYCA0N6MaBdTB1vKBlKpD1ZvDTmMEPu+vrZfrc0Is
wmckb2iPsdlM5QSqKGkfAK+3O25BoVkUOZDoTAjoZanadFc159ifIe2VNnnS2/mU
5zKU2bbT+c3tW2xK6IcfY4nW+rH45mD3Xnbk/IQ3YFp0q/rY2xRqWgL7WRABAkOC
wsW+f9WTNaysehAKugr6KQHaNs6+1zgnck5NcmwzZv59dLuNct7HZbX7g8inMz9p
n6gzJqZy1xlSRwybomu65SoiqQK8J+8ffGtrXRK3gjt40WcUTbCnJxg9U98NZQkn
R6JBw2/1PSn/+kY4xh5qjqKaIgnOUU8f3a6pgyz6DPllPJKMKyYWKOGKyZ9gaFIb
gcXaRXE95anZjc6O6/8gBRo/Kh9GckSxSrysqhDzt7iBZGi12EviIfVfvxhvWTVA
omhahFCDE6/ARhrSgcDYdes8i1bSfaAdegel7zpjYsjgakVUkfjY1rWbj7lKRFdt
Xv64nD+aI7L7Wr9Oq0mXmk0Hln5LQPpj8ABC6hJ8PKzzwA+ER01IHOh7e93HVzdt
IuntEv5mSz9blzZfH4Qkwf4JKI9jvWAVHdBMsXuNYqanL4fDKQQZ0Urp9XxAdwja
dLZujQKXVCrMIsL4rOz3ASxRrgaZCXaiqDWziMg68t6XvOS7QcPSK5xdeuOkHt60
21Gw2NK639QDFdqWycNpDN1nBjb7HsnP1/U0VlFu5UgTEfiooKjTf/+oblHit3FV
UCyt837+NBUGiXc/9TGnZp0Hf+yHcWrA+vMyJFODsqjxcaPDgxz4oLW/9ql3iQwm
riKvbcOFAV+GVAEtbuv2Bl3PTDtq+8sdZRLnOJEtE6Rvuzk1SGz6QTF+TU/9eIzZ
8iHtrMNAnTQ77bE5YN3gXI9OuvSb6jAPd6P3X2EFkbi6jUi3GLzJ/uBd9+3DuR2U
FPU6H14BBwsVyQr5pAqa+2KU9dpZDRXxy9GekOuOSmuJIjc+RgSEWkQWEPecEqwR
Y0ilyNxuPA2RoMqPHEpOCKtI0rvGA44sc98MhFLKgzdN1fMU0EeNOilP9ssb1Z5r
I/REvp65wMN9UZ9WqU/zNcmjkLjZORU2OndQCMXcff3mCvQWifj0kUCuJdNPODSl
sS1Q7O4YB2T14lj5xexhvK3WhjHGW5pozyegDERk98vve68C3QRwq1ia66bOdGc7
DV7BcS+9r9GKhdBiAk6AnrEjAee8NT4Rso+z6OhHrqfLncwgAFqr6uFUik3mLiMx
QSkFIcs/LnxDCMOKYPRooefoSaChcMtoPgMMCjlRcLgV8pmQtrg9f23Ah3ZaJfFx
jmt+K4BGsjQ+rk1sQGZgglVJEfJGYNRaIuh10PfaCex0U4iTZ+fr14rfnuKeJdGz
aFZozR8YL7udKmhTXEZCcZJ81Z6rRuWp/SVOzFDAMjORYwx3vsgwtfx250w2qlXR
5nQdLsDDWQUKLLCfOH0TFLCCgG1zbg6CM7dSzLSAal55AVIotse1gxf0+2n/tPNf
ddr26L9CjJYJr/WjVzRhoRl9fwVlU95bDCdJC7mVp23VlbdAzCfxNifFHGielDFW
Q+u7ZYt1SDk7bzZR5BesYsocGbdGiE2lEIHOBXx4dlEyaFoa+LHhQWfOOJQ3w/TO
0kntrUPWzueWB/Bmkm3ob6bWlgRukWcPkFwn/ZETeArwI0RQTys4z9Rk+099bA3N
Cc+1L3qF5H568LDyCvu2QCMVTwT1SL/3Hhg3AhRh0a98798hQNzm3NNE/kSslk1o
4JM+vqwqUBH5jqk6XHTqe5wkeN40LumUUHV9phZArqYHg9e99iUgeVMJPpCQ3bG3
t6buXOUA/5Z9fz8hwmRK4zJdNTUCElL0odaN/4hQJonXReshlnx7n/bNEashMczD
UVeafgzsMumNhM+bopMqPhgUyk4lMfsDOPmgL997wenTgZYEIe8soaHaVRVSSFqj
e4tcYk219aaIowtSii9uGyJhpDk16AGTdFwExlpmfoGuX9uBfc3563FeBzmnUl5f
YkDXhAKUVJLtfYyfHi8YX7nyqwqtzcGS2/C7RbBAJqIxScYbbAPeLC71jwJDEQcR
y3YTvFbENy3rhyjSe17wyx9t5cN+isz4P+Y+LNBmw7WAsszUAfL3S+P1K1c2SXqH
lfdOdLC8QZ8l92UCUckpzJaRzpKuvFWypJA2dY00smH6xs5TGtlWYlPfi3fyZXI7
yqOVtMHu8tbc7A8kBKo51OKmwIxdbLuE4yBxZQuLjU+1YbcMP/6ykXEcsL52fOGb
TCkRl8IYFj0lh23i80c5KFU73QIN72C0z7YpIEGhdEjanbC0EG0JdmsKGeK0Aq0J
uz11Xx1UTU1Q47Hl+QYXh0wUXe4w8ExM3eeKQ6S6J9eUUiuUolV/ROzT/MNz0vmf
91r+X4T48/lOIqmC4/Qsxxy2eMSDkuseiEX04EElvbEE9/HGs8BFkpCBV/f6vLrU
Eg4dR5WqOYkNCIbjc1xR3tC2pyJ2T9BLL4DHnMv9LtLQR4GowAjYtFbqpUgchVwh
OOTfvG0iQfAuycai6PD+jgOCgOBesp4hdHSHiBNUQY51c59IbzD8RX/PnByZmwhT
oocZs8yCYlMVuvRfliVbwLgu4qRWjLwZ4ieI+FTqPEJJj1sopolW8s+Sps0gf2LO
jAVW+gByL1PYPZLvi1h3luffVnCvJb4RXKN2+mVuBen3xES87MUEgJfYEMHeXOjA
xpUuOgQBjg1Ry2k7yvXPzCeJ4RFLZU6+K2WdnpGBwN8g04HsWKUAj11WYE8A+9iX
RrccVKJg/x5g9cwvsBqsBbjHevmWFWAH/MEwRrYa+S/lpFVe/eDlFGtXJ9Rtirex
cdSBDpcWywQjbD9CrbfzkYlawTj/Mf7VJGl6dZAQ6/5ydVKqJG+9Uxoaz4lKG41d
gQzq3Ub1yrv9tgHt1jJrlstKMSN7xQaahLqeojsORWZWtKHFvS83BKSxDY5vb/6E
8uiZzGLA5n5vvqLdx9J3ha4SE4wlapNvihYufmQx4pGgz+IAh+6JFyRwd8eLyMla
iPCr+uwtXFsUA7d2NxcSGw0zdzumCtjFmcjfymdGvWitFmqSfhNoHrdAmtZykx28
Jm+fOB35gnA4yUrmwqZZXkRqZVwN7gUAOin9KGApMUvK8GqXwjpg8rx71Ufg93F5
Z0G6Ptzb5Twc9eN859HhSttfPhrj8ASt2vbj9lSppearuWCNg+wl+sTXh6/XZEuV
2BQ35q8mnkjKsxJRRc12c62JrO2ADEehfGHF+kvYCvrc9LAvnHLzBPUQidboIfcb
mfMOcdIdobIKzGsOTERizqIiLmtllIz3CWba+0mcOtK3cNFpYvj0eB2HkUU/E74H
TzrFL/P8+QilVJBHqAwSf0oL+VJeZdtIeaH5V3YIcVpGrlVfV2icu51Zjbp88nbQ
vfQuY/yhmaiFvUbshmnSb+fSSmJjruJs6Ct8lokkLsW31v5WHG0bGQLOyMTVZW/+
ZXwpUo6dM3DnDl32f8qUm5JcLNn4NNTBjOLKtfvVpgbqoMQiD9eZ0cfMmifAmxqD
6J65fwp+EGOBVR63Hli+qjSZgykg7EGOgbauWMVjs7QVBWZjz7qdtXOqUdLzlUEq
HiVeQd7E4Br4HMwCOZCLfIOX0L8R2oraNhfeae2fbE2YuCMdepT5WqQ/Uue7IEv6
MU2I3cdb1hNjnCPbbd2M3V3NnQ6MNcv7u2CAV3+jiYWXPzDCDQpPepB4H42NiPhy
E+9vB5CVMrkGxZ53c53dFL2yFDQB+I7+83D/gBd+pnf7VXrCoa6Elj0gVSRYUGLN
KXsUBzpQZk2vhTI+mD74TOGuqxM+k9PhBohxokUxBOuATpGRHyoNI+hcdsDGMDw3
7m6kehmA+TGQVTCiRvPSMr+UsGBq+ksatwEd6Onv3VW84XBbyN+hPruqkQwcZ08x
vYHVZvQMSqgh1mTxgbSFeGMQbmpiJIYVlxwYg6IF5g6OTdW3N2GPWkm0ELu71tSA
HysqXBgud4Cq3GeDic5shZIVyqURknFzK839QBwNHSNvWhQ0LrD8RIEQLABy7ZW0
TCrfQK8DZKapUTf0eMqDlQeSNob8EoQaIjbRD3Ao7Bz5VB3rJkCvat/VOp/kH9zA
70hL9VgYYOQZodvIXJHwDSwgkabOyFhleSeTyKUu76HpE0N32h1EXbq6VXKfV9Zp
7WqLWyO/3cKmR//UpTuO30Hv48RI7N1tEi3kMMM8u2oY3L+swUHDGG+wFoTPHNOI
L0w30A24HDrK6FdIkMwgmA22xyujzc/1miwMQH49NR6s0iPeEZYWWynYPNOyFInO
9ehKJ2L7EP4wGsdEpooAUF0SM7CJPpTtsuvb0tJim92wUkUIz6FGn0rl9KG9kZnv
4qIu6VH7JJ2a/RKJVdkI/Cv1EUKDX6DFUg3xIaB2aRmjKTyMduRGhCDf1cfYm6te
2aYfLbVnsZM1YbivKu8tJ1Y+l+UtnfMHCTpV6tZ//DsvLf0q+KmnjFrQGgiKhBk0
Q42p1p8BjqZQovLELkJUN7eT0HZlH/gYqRPYPV1pHmUvewrsNgQknDEJC8I1b6Mv
FeUP1LOTCJjDxEEcAo0xUCoU76kcnkCH8+gxSrlFmP2s70Q5tMiAfl7oC4U2EFZk
vi3cYK2jdmWM/X13g5NXUpObcUWGyxf1QXwKn3IMFvBLEZNU2vUcQKgAfcXFOlfG
S0kpxZ+R0ajIqM1/3q5PzdG9WZ2+cU44Nlq5SaW5C4qM+GzMaDkBsjotU6XzDRCp
QltUmAXtHjwFIyvAHvuLL2p1Cct4pCjxLgRPmhWlrPSHLODbbNlFO20bCi6TtPwy
63v89DZeZnG4wWdm++JgjDXznERNGbF8mGPKs0LQ/OK52L+OF2D5tJU690ed9rQk
jfe+tUgnFTLtGhkPaaiAJCRzcFeq07C09b/EE46WXijlW8sU0JI+OBlzEjpI0wQH
jS9UJKdHVauj9iobounVC0NAG239O4LGDzMNgOeOp9gQpTD5eJgTZfiqiWmKP70p
r76rkxLMbtqgMfhIiF375GKLPrYCMf3897ZEJFFkYQuVPKmN5Kt1EdVuqQiVmrkh
2rcG/48SIPENPfU3ycc9pjgYtwC3wj+sJ4YdxhmcA+m2WLFtsU0Pe3ICijfO6rzT
DCbf2ANSQEAAmk5OXZ8gf7+E0h3VdjSRICOY3PrGI2OvxLjKowUkJoBBlIPdjfxx
md3po+1ETUNvxWkHrhgZvr7MIO3TL2Gex1o17QpYHhYrpSKXnguJZcrlm7WTwT1T
yIha2tOh3dKxhz2ZT9G+x/ngEzPLSiuEt4UZOKDGUgq88MkhAxE645pvOm8iGuBd
Ph26fsUcg4BA/8S0NCBp+KnZMBBHUyMxFGg78ctOrQWIHc0WBCF6iFei1NwoIjkH
Wp9FbP9BRvVraeLXRpHQ5I9GgMzeo/sE4EA1k0qxeY2sTQqzSwPtIdCCie2izaJr
et6PhQDXPXcBe6p0wzdPHDn8whbjv7EAcHpoKhCSvZyAUToY5ocrOFwS34oEnCzU
uoe+DJ/PfRw5eclonB38QY9iVCf4hrmWqrS6+5+nuGLgZOINhONSfMruO6eZe9Vf
BC6/N+/sNUhkGXpt+fIb+rHOLs+twxemMtP28exp0MWK0JmQabiZML9lUmMx3HEC
Q5qJf9yZRBUZpk58cnrBAuDfIDVfP6g45iHE5JgKVaH8UsDTNOWRa+2oA6Prco0C
p3cQhMeCMWvoz3A8OZnrJ1hesk146gGBT0ITn6ccLcKnMgxcTIsyI1YlFvAL3dDL
6GJ8FZuK4d44H10k2gQDIN0lLso86yxvPiZXWk552Wpfm3OEIjO5rVPeC9kbnBHP
45vtny/R8W1nXl+UbUYqzMowsmRJnB36w2uhLXxm6/S5YUdP2RMmPFtQJKuxmFwp
EJwcB+RoP8OXtVT5VsXUG1j+drSdRXfOZ/zqLlX7ZgWzRqh3Vg26G0MdlXBjjORv
MFGwpy8jNWiCcWd/t8sTN3Hn1fB2pR3fHjhQIt2rvq+hE/VLlCQd9dhibFHY7npi
TXRvA48/+Lv+2Nq6WESQduxlKdk21ZvH29WNJh/Ytke0AMXeSBPk7VpSOEwj70pn
6RSSE83SOlN9zI7Fa4UmxXYs0PrX8rac0FO9oaFXod9dWMjrP3i2ypARB8LOpFun
wBa537VE8Jv0mYOgiDH4BOSv2bwBDolSFUxooWKxSrmEl146pyJ8tWGKHnwaboIs
qiYRVb2e0qkTclNgNqr8ANB5OqE2Rt4hRVpBfcO9Fsb8G2qFDfhnm9Sfnapz2m+s
XnBUP9lWyhmUC7cwXNGZk11aonVfCd/unn4CqT7lHN1ctL7UHUnWzf8wcDgyIR4E
97LbGAer6kwaKbc0XNPNIhnL9G1I8ZHdbtCwKGAu/K7IXW6IHZABZENzWwoi3H9p
Fja5pbHWL0dJoS2JHvFsxP5TVZuook+SDQcEbMQc8XhzCCRKnNLcpYxKMaSglOs5
CeSiAHEYwBpDcIOCG7ZKcKlQ77D+sjiJEj1lBBFG/AYiBTNcKi7SZD6evB7KMXKj
ljP+3M/e+Dyw2PqcbY2aWHm7/jU1TgLtpho8WKEL5QPoVMsCIguezEzi5YmCFAYi
FDl6CSwL3ECHlnqsWG5wriNkbTJZqaEq5pRpMN8xvJn6iToQEXTuxxrWQvb1xXYm
6HSRhw8pyxwuwDuMHtL8k4nJCa8zk2XsUYth4r+xnh83BcvA3okFUtDeMbMBg5xy
PxP13hGWJlKjcJCUoVQiLXaApQTWi2+eeSWFX6DuCP3v/p3/eAwzDfxjwukOGL7I
uoCE9wLi9eE4QCRE6/86E4B832w+cntumxlVKjQQmIOnfpyFCo7B+hbkpx8kTo1l
+J4/JhSjKh57MSZAA2hToWS+UYclTwZu98jf4LvNCbLSVy2Q4LcCMJtCjujS+W0C
xDBZu3eaREZMti9KOl1vhND+0arxplHCzTTRmQJpMU4CDVWVYlVNPRgY58RQpVP7
UnpcFXdMzBN0+H40wLsgAWIKZPlXHxTtTL3zmIWNmlcbyoZX7SkGnYseUNvX128n
Ar6GpAuIfoB1VPiU3aKsh8ALPC/lHdUnoFx4i6XnTuKRhNngZPgdAwXWI1ywuh/O
La+udnl97DZJQpGXzgAQYRPXkTHnt+BbVP13adeRZ9Ixu0m/9OT3YbL0nEa07Jna
8LnrivyKqCubNIU8DxNfHakVnPze4DgxaYbaFdB/uRoNGFltdYcSdAv7tIpYPsPi
8uVJvMZ1H8FxPLgphvb2XW0wKBjZ6ddlaL8wAhuTm4F8YIJBrPDHPayZ3N6bPSUK
3mOChgUIvbmYBABES0VHMTRUpuB74ExLyJT5HZu2FJD1BhWqBpU79X8m0ZQb5RV7
wQktCHXfamK/xUcTqxgM4YgEvrNTjr2SZxIM2SjsJzgQ/GuInX25/5FNNmLR1hKp
aVx0xLYL+qzsSLd+2eC9Utrc9ArVlQfHhHwUYjxoUeONeD0xaUX0jkxROgNroL/T
s3q6+ee1JUCt7g+mYvonaLX8uuQJuzqk5vH/SCxl8vptRnVdOnFwEmSuWep4mpu9
fFM8lg7G6Vp5CwDVEBoYa2Xv9bHxS/fW3z0421mpJLhU0Sa4Ss9HsSWwRVZgQ1Xp
SHCqE4h4HcRDEmrPyrSA5vJPLslIU9GwgFbSqU/ytv1tozJG6hr1NVUVzR/tqYub
ug37M+6Dnz/HLTR1eO7Ln2aVih1avRW/vXH3Rv/tqjfHhU2P3QZW9Kdfe9jAlB3g
/bo1HQxKpi1iuzBBS5AF4JFmFSLcO/r/2K30+AfVQp+mJ7XZ012Pyf7QHHCZx94g
7Wt64GYU3EII9APbPQivu2wOV1n3/PKwru/4tyHmXtJ+YpajyRw7veyCnhaJM0PT
idqJpdeij7/U7FWtqmn3PZsUwsiXVBUgaXu1orXBn5Ils49osmkAruN0vkvGYCAE
74t3JqPPWS7z1TOD1ksIeHZnTkyT9utvef/GNLgxyxTXPPd/OVuC7Q+syTi+a0Il
3QtXsUYJ/zUl7QWBJ31qaQldOVmFs9xwkfdXcwFWMQrR4j4oahNH0fMLgTMOrWfB
tWTcwK60YUXIVf0RHUtrByZ9TwGnpW4TjsNDrlISEDSj1msKWqnGGMlfzTbDOKm0
+4WfkfcYj6yp1x3Pt30QSN7RYgxg8QBalHDkbUUnxcpDFbX0s3Qe7LM0u0w7FJXC
xJCXlWOg0EDkxmb/46mUz5zei5szrn2scSB28uUH45DmnZsb/8sKoTFhf+PJ8oG3
gBrUOMyo+KtDbMGuSBd5k8pdewpiwXjPXb4xxfAJWFnBlWVVFAjNvdcTLbt98Zp9
OYtuL7SVjjNdoG/j7IY6j9SjyHm4igmLj3WDeeTy6z3u9QUjuBmPXBvP+UBJLZ2m
nPyCS2WaG4nZUGOo/JRCR6MZ4jvVQFN7NfpMii+7pB/CdBKijMkEWTp6mGbBuqO6
6vMc5RtHT2jgNUJklXWKg44gPhl0yJISAAOZ9TE34KRA7rULsTIkS5/Kpe0+xW/J
9LpPP8V++5LcB/2NuwBfQ6nBkYR/2z+7pgEq8mbRa88ADNtUpOmgBJtiOXdAvTQx
AkeBuJ9h8mArz/fwfHJkdpXNE9FoE+mmlcClJxtZXj8XdffhRiTawpoa/pgq3z7c
PaIyOzwkTpn+wFJLiRet0ETogQ0iZny+pM4axcG6eqAJxYm1vx3/ITccjSqf7Wb7
1Y3VT6kgqTVnq7Smejgg9RgFinQSqdCKHLo8BY3r9bhQAsVOGIrXMwHhI/KHjDok
800YmY7HyHbJU9BYO8//7TkAE/SwT+cHRPjcI+szOEndqZh0MbvA3+yW82tsQPj6
OU4D2bNNg4xmC4F8xigLm00+vVJoAybK8wnD+RjCp5H5l0cxtixvCYgeNwhfvz5Y
OK4TikqBbmmV1lcNBMCmPxEgW4V9F7TgWIzbSftUnc5ZATE0Hy4ZBHLfFhYTmSqz
yf2nJB5j86yupWC0xEuiIEtTE8iCqHpH2qTTikRrUpL+bGKv924+E08wLk28/dM8
LI2LeDpuKMI7SQDI5E+Y2mI44KRuSpTfj+gVwts/krerT0n+W+n4M6DHijeDkGNC
th0a4WtiVlLv38UaxnA5AcYjqoR0LWcuLo5+8b0kLd0uOgPWqBian5//Fc/uu40X
SvykH8nWv1oitoD76JLyPu9VqfBYrcyLsKGV6dCc+unDCg+dBj55Igy8k+viZ7HQ
Munr/5lFIU7pU7zuV3FhHgoW05HCIEWO+3EO4yBvEaX1eKu0G7b0kPUMA+uBIWZT
7uDuldLrpns3ajfHeSm/1W6mXELup0nggos4j2LBHYJjOQvobtsbcLIrEc7XiPFX
keADpG9XOw7rszi9Tm+DzbmZ8zgVEXgUOf2jwL/wR8cpyPsPw724kw2WEbuBDq0Y
BnT/DVnxdf6cDgRXQnOuTCalSg5Qijg031/vAEB8sVCWj0kXAbGaRFQT9BN6w6mb
QF0o9cWZ4B58bkGSlcgA2avdLoiBizbdNW9wyFEbBPZSjXRC4b2ANXWL5j9am9bd
LoW9AXxM4/xkt57u/Qqd6bDS/AbuioAptaVDRQuDHz9fsFjeyxiKcNKd0M3fzPdd
RWUk4r4eVm1OpIWet92vVnGV9gjqHnnbA5jIzf9tZJiKplXDr5Q5TkmaoV/IRk+A
QjXLSuxGFptfvUMabdLzf6FINPRTSEGL3JzJDuZeGCk0Sl5EBGZ5pubmvCd732Kx
mfPp5VTaa1lF1DmrXGBF0UPXh+bSNV3KNoXwSna0TD5LllT/tL4/jAAFS0lHYWvv
1zVDhFVKXv6Fmq3Eidi0p8ZHn8zQFbdE7CZZYXz/eHTicSVyGNYhUG5YOv2ejF4x
ahfq9HBqhETMOsO5HxBwS6zz3tFHbtmWBThXReH88N8/8bsGGN409TESoLbOUOwh
bSqXtOTLiLDLsfAh8rw9CtJKth1izhN+8viJc3I2sZWK3E+v4rpPkYscjgacqWzf
2FCZp4JrZv62sIix1b+aEZUe3m6gOCXwzTPELHmy9fWilBU45/7A3tOYWBqY/DqU
dBtV9Q7OOlssys22B8IM/+SzQv0TJ3yJDzt2jcx8WejKu3H+46mtuia0sGsKAZJ0
D/JKeTsLPjw2PKJdFcLlxsLRK7fuEmULa4iCLp6vgYISuWCSvCTD/L5PohFNFvfP
0E2mCF1SZL6oVaGGGtLm5ykpHdeSjzgCVYr/WqwpwVWCb32Q9uIOvkA1hLbkHczs
UfW60a1yDNvE93OGiNBa/3bWDAm7/nYkOM1cV1giGRNqhzVwglybiPOHnhaIdF8B
91DhAtee5KWnQ3auBZEuC/ihwqynuBlptZ6RIEqe4IqKwz04lA7jzfiyNnEWBAm1
H7Ah/RcRE6cyiazSEERfdKm44bFcFPItRlAy8ZBtJR2JekwaE34ymiH3P2ugvOow
oJP+iJmmWXa2toylFQbxSHDy7yIr1QId0be/6gsLNzJQGSBkyTBgkELyajUAwmIO
Ioe59wM2LETiYa07qy+jWYYMv2+UrErMP4Zwh5i9O3cTOXMdC4858EDSJgDrByf/
ILSK+Ps+kCQO9pHEMUqx0wMTpmbJvPg44VFw4Hwz00hNSv7BRPb0zTZcIqmeF/Ot
MAchrTchTtOnyW4jOChKdZyl3rqro9howOF3QGH1547cI4ZqKDfmGFqIOP17r1+k
`protect END_PROTECTED
