`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ookqYF61rJy6tAFRZ6dH7CpT2o8hHufJc5eOe1VSQPLwl+6TwDyItrCQFBnS5cH
4FkiVQMJKxiy0S53dvsYd5lj8BjQ62J/fpTLe2TayAG9DJjz9yQYgqlCQlfVkmyU
qgNml95XGcvpOtw9kCQXvTZwd4DMZo3141N+ptpKGW46z/mu/fzy8Ncve5GceKff
Hi6gyYrvK+li7EvIFmwrh9IqaHANBgsAaPKMeEwRLiQloA0oMStu/6FISe2vZy/m
YQfNapuNpgqImV/aNkWa9Adwye6wvTkReubaTkbHjCBsyHnXvLOwHJo6BLTbzM5R
/Fe/NQDbZztYEu/Pc/ze02jtTTsmI8WZ0IehWnhuYFo2uCPHXFwgMottPKSAUeU7
dslHsdFvcGErVgsZM4gaPt0LKSzmJ3y21vCx3XBP7WAKMVd7B7HP+FU0gPdAbemS
IbrzScCqofizcLMqMEI1GJtUw/L0S0i73X66p4MjyAWI7VBXA9Dm/Apr1izvntro
HjxGhbkJ6FiwaxZ1+rRPocOeNGae7jSYTZhN6d3Uh3MaqKJTGPZWxTVWGhK8hK4S
/oGB49E95eETu6EvnVdmOQMFu4ivS790+mm45RHqRW8jvchCQsOq3ujAHShJeKxj
NWMWCBV28jKywRcXmGgL17Uic06gWxN4uecExulm1Fu26l/y2XstXUokgtYb6Y0J
QFde9/bgk4awHZscieytIhj8fG34M6A53SDB5uwEwGjNLBJI/yrf7ckA0k6JdBYp
Q9PkupGhV06HuyRvR89iDbBCpLhzxQK//K1tMsDc/G5Nd0RmwfQzsFP7urBtIy2k
UlD4mhRP6YBDA3qVJC0sSIdK1yVtvJd+GBfjJ3MElBZ/Qz4Sf9+k/Vzxvrjbj7/P
8mj5Lo7v3tAoJHZr4JsdPx1OPKzSUd88meUNC4BqIrBMpD3GWbfoWWlugjq05y3l
HrqrnKoFsFcu+uxOk52qMbhQiT/XXdekgWN2M4RwZsmWMJIYKo9tpepJY4yUrll2
35JKep+gFro2POX9PRQBFVN2wCkQQSAVCpYzfQXuOCOJYQU+2fgvnj6/BaQfKy5U
X3rJdWKcjbfXJ4I53Lc5SNZ1M+UrALD3LJ/Mi/2fXy+GZCaY7iqDiIJw2HzLMwaa
Rq0JzCjg6wJzc073iwSpMIG5BnnfbZv9/hfJDM+3nRcsnvLDZFU9J0fIq8F78zOG
DpzOkPzkDfPk3M8FUtnCxg==
`protect END_PROTECTED
