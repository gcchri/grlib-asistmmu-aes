`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1arvaLVuoLLPjZv74ZTD4J1HfIqB7lNS1xi4gin1DstNTiSNoyMS37QnehLW/s91
ajgiXd9f2bYymteKCWsvsW6dIZulM03zjxfOhgrWVAUFKl2AEBMDySEeVaQ02WkZ
Upv5PgNdLoXiQb1A7K4XrtY0bKf7d3z4NKudkFWEEWZ5sjIpzLyNpnHyfq7o1L/H
7+eKDtJaRsClTnyAqt9KmwQkbSuf9lKVrVGPOfG7VgGyPPQCuMbMrt7jQS+5DtC5
6txmY03DMPgTU5+atrwDEA4/fIp+76ntsfDx1t7Tcn+dMACt+CmawDC4rXM30DwL
gZGzTmFZiHsPQcHbz3aE+5JsSnBVC3iDdBTmIe5q8+e04aOwnmEHjajFdpX2x08Z
9hhuC0iBRP7KriBOHBTXtn548CcA4CVpqqTXfZ1mQ8e3Y6A3YauZjU3c6GJ8z6d5
+nWGWumPw5yJul8qqMztsGsgp8O9tpi0rKODqL4tRH6Td1SrBI6vg69H9L/3oHt9
vWY1ZuDkjK+Gc6vGrb+lJz1k8RaQe6C1BAhztkWoP+SFFu5pjv6pInuXr86qFZJs
`protect END_PROTECTED
