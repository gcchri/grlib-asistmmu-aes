`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kU1Jkjc0jIiZ+s2hHlb16NSLjkLP7PFxLFFZAPskQnl+TfI2mpPtg5vV9wrQbbMg
9Ta45cLm5WizXTANkzdAxkDuixXsn6xjVdgJA3YCTGTCeQ9BYxJbbanNOsxXJdYr
KGtxs8TWjruB+cHPunftHs6E12AbwMtzUB36GJWe3XcYPqBinD1rrNUe9Ydus0t8
ECsVAA5rJwTsd05KZmu5mrVKe0A+YFr4W86MMbhkGz8NdADsEiB+ABSZ1TVY9EqR
Zvusw5fkH5MaR5kiG7WIKJ/Vyfija7cQOn2zmTcH2W1QmcJpZ6o9Lo6ihEYJyLa9
g6sCGh8ZdlbWxDqjgct75WsZ1tfr/yWHkJOUCzGBuCx6fbufcIICRLNyuqhH9iBr
5bgp+NwJk/VHk5a8LQFJXtH0TkStuJSevECaA+pBv4Q=
`protect END_PROTECTED
