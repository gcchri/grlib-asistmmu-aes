`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C6rkgNERUYMRosYu1pqvtsJmujL+2+5ekys61+srAU8iFb95vmSCiHUQY1BOJHG4
5uy4sNklK+Au6VEsZFncyE/iLlchjLV4X5IgVWMBiXZOpXmhG32U1gIgaknkrP7N
w/10l4rpgONT3ORXKUXxKGZBNZZ2ym04X0EjC3hxTR/0JOYA+bX5+HHbERtiAkKB
TvIVa7GWUSaScC+1o88gjuYSp2jheHBiobz1hALYG6QRwqsRSdWaXfWk015FRvaL
/NV/d+yvmDO/4UJXeF3vOozGwJYXGIPVLYd9E7MFdeRcwVBBUSdfOGhnQskoPa2M
x62gDNDNGVwxGphFpEAJ58SYL/fqSmtc11zZI8kDNY11Y8YFzl0N0921uwtBk/p/
luc9RNaum45AN/yOGye6hoJkSNgrPZlw8iVO5oBJih/cShxT94kD88NNyqM7X5L+
nE+XkumvlKOFQLeN/YRX6vW4G1/tR0GGRbfNmNy4bvCMVsMgQQnfkw0FyqVPROLz
Y45BBGfnam/Lx1k9U2fL8m1//RopofhwFYj/U0EOBIr4P+dKwm3xlDrtmQJm69DO
IYJhHmwRCmMQi6IOMEqff5vBxaWrdGJBu7kwYnn/lwMVKdDy4SxQfbyltp7K7m9H
0/ICZy2afTXm9KwReWEoKH9gw04JOY7yWktPCEgJ1jn2a+1XIHYbUgD6u+X4JKcH
gqjZJdW/cxX4zDbNYpq6G91hgCGCfHBS3u39CfDojbwIXVZxMReYLO7jONx9z+iI
WB27V4Y+AaCRgQGkVI4gqtYOniS+URn1VnHwizvx3fHzqlAyGckcAAExOgwCEe1K
5K3T68Ah2P7c6vGXTc8WtCGEDt1EWyFmxn/7w2YCK6f4nDwz4lPxl0LWX7Xs8O+i
e+yOAdEDE6O0GcYbsCFPyUPqvXrc4EA5Zo1jxQLRko8Vg81BXRNd3ojO8dSo9h1E
twMwZr9tesbdxHfCeIQvbu8STtzK/sr9YsvHmLOEhA9f5Ew2GtTHQ1QCZwhjsVNo
dKlCyfK23piqua7KUBRCSLZFv0SxqDv06PurhNF/yQGt8JWyPCr9mB5hWbUfyozm
HLnUhau5I3VqABwRlAogPDUr88DvsvP2lgGTp71qk+KJL7fiWSUXqrpCbtDfZaFo
xalAqqkA0k8/2Tlb8n48EBBPhUyQZY7GzLWGDmVLKohtV35nHjd0WfxpCLURg0lq
ddCu/jaFWbuexs3d6J43mUODw0iGTpD6FkntHuEjEo299eAYkjxaNNBRblH0jGLJ
mDC0agJeFhemS/x9PsQg/37hP65L8YXT6NNx1rI74Dapo0g2rjU3hVvf35JwCaoc
ajd1mXTyL+8wZ96ICpEC98IyHCQ8mEV7YwGNcj38R1DD1NM5EdLRbWzT0r0PBjr1
43X2/uehDyZf0/EMSAAKLShFrAWelXrVk7naARygNckLwRhHTU3jbAYiPBfu5IMe
`protect END_PROTECTED
