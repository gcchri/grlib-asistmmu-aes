`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rkUVCbO7BZK/I0LpF0VBhDkZiXjZofs3aoLRpJstjZahb1Sc4FgEeIgvAX03reqq
gzRdDNvD692MNSAe37eX/DMJtNM7OEPAqtheKzDjBcS6jrJV+jC+4AUGMFLL0bOk
cSm9fAWrlhh+kITgMb3worcZhzFXBXDVe1x5zgb8Q/DIiEoD2h7IDbXWt4Xg2hX4
djMlZ8VxwP0TUusj7ZcX/NSSoYguuhQ5m30KIkeI1bpV9q8oi/GRqy8qigge9B/H
HGlr6stODb0rAvGZw1ngH54J1CW+elTwATM/7p3M+ILzz/AaMPR7IXDIhF72EDyy
`protect END_PROTECTED
