`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tdzxUYIaCCA92OlRi2X0/6W7EWBz30Z4DvYqD8LNVb/BxwQlEPWJEzqmc5rGspxk
FD6ewgnUpqF1N28plB0OQkYDwxUZ5GXgyVglNlOcd0OO5k0wRW1G/cKXlUJls4sv
uATjbyPWAiWea8JoGREWzvBfWvginKHUXM+aSakg4RmqIMVyCxnz/MFSiCfYCtbk
uRVjJrxNhH/g749Zri1EFzpBlk7mnQE6DrkaP+A+AjGVqpG//se00pT/es81A5Uc
yJVYauWi32i7YTeIXQGMvFyxmP7GpvWekP+7gvNYC8ClzkalOdaqMrYBBDYMQrPd
73zJVtxoFqr30DDctgWk0inG8umhtlVNdid0etsCm95Gt8M3yfXW1OHfKlNgILiO
tdSbJ0t/rX7zSjMj8JcEI8hsoFO0Rxgq/K7vNO9pGlYGaCwhp5lu8BjJUNoTQVDZ
XAeahMHNfeDSnp8DbVGNLHEoACuNl7g/HpyJY2FqOVvXHwGK7OZgDlnO3vA+RxcG
88n8roUK+vWFVPVI4O21bMOV/lxiW1h3CwoaDfPSk3VCz/zrX6VcVOlGdK/faBlB
IRk/KgvihPNoya1GstRpm1IaSDVCIGn2S+5sHvIg1b6A9JnwJMgrAZy78GjtHMbH
y6BzYNGSsBHtLJlIKOb/3AmW09e+pxjfr/L174sbHBJMeyGdKBECTehrZG0ZI1O1
THiSF5pJWqzUB1zCzZsg2yARmaY19XiTLTMIZatz2iEP6i9Vny4KXXyIQHoujj+m
dKL08RITM2wBaFRFjdWZfEbn5v4zIDfJZCU/h+9xFPi8gVgYmw6W4z9c3C8JNCef
bVsoENo6vKjPYdM2XPWe10cZePIfdAF2G3JB6jLqsyrTEntmVIeZBavpYA2ZPzPd
wQAnFR+763sBL0Xroq9XCQYR/iBSmejvZNyEaOuwr+8=
`protect END_PROTECTED
