`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TVaUqV8a3DkI4aeAjRJtOpLKky+EHFoE/oY0oCU4QocjqRHv8zeAU5xZEhaYYLRN
vebBkP+wYVpgw07iEtCmW6KpZY5w8ied7dnQnh3JrZe3UP86p7a/6zyCxZ/WIUEc
UXospKxXDzgc8M5jzZGivuG9YZY52QftJdTqc4RYsRzkKgWExqJRfzV4c7anb9B5
okM7KkYbEmrIM+GtPPsO/K8nYWyDBl7OiANOOzJOTGs8hfJ8iFgM8IMYWqaswyyD
qh0idibpyIvrg66SlSihfexEstNK11PHXI1xDGhEGdm3XP6T0jSZRUDziY/xV781
WwdYgq5eWnhBVrXY3QVlMMGZ8C4IPhfar1GViSbr7t8V/wrXrVq2z8wYHrXXVnq9
2ao8x/PwX6BMlpj4DVm59pWF3hIlCXElHQy0hD5yt68IiosEHvE5mPMJr8QXQ8Ld
XNNhlMOyQZndkdNRER4TPc6HMJIrJtCndjp65xo5132+CnyCdR01ORNobT64fVIS
zC9u9LUgkAyY7Mw6NTgTu2gC3bRRtnQjEriqHt+bBgI0TMSTiJWfxWFhlfVUxp5T
toXJuWHhquF37PI6ktaF/XYl9Z/9F+Uzt9IZqMwcbPiUZj3dJ6FjggngwGEketGi
WRpU0KPu27I1Li3pVIFecdHI5/5H3Su1BOUJF3NrA3PeQq/+PNVWevgBrN4/04K6
qV/oOjXDM5Kjty8/iJ2IcFDx+QGamFc+mpF529ki+ADLYBZan6IFU60A8bcpm0T5
Ghers4NU22oKs3aqyS2grkt3GqPqewPvFcdMPlOLURywaLIy/1xbCPgAuKUMSXLK
r76/XhjFDIU3wM/DigGGYft16CuR2k1E9DbopJicwYYGDaec9e/ipih2F3WGbAWz
r8bjqF+DapObjdsU9tRYiUadsn8K6p9RzJVa7RAA3GNVxIFDq2JSPDP2GnQa3Vo/
iLzZoo53G1p54uEiUr0gi4C4MtAU1le2v2qjLnlftlR/QvqPY3HPzYRBykKPeHkR
9V/5bi3hKnd+jEPw0qN8sXKaMXuSz+gu4B/xO5KXEGYtoXg6Nnj/oHtTSIPdmdUu
AUUKQt+y+wiZLTTzDu/UNNMa/lZ4l72YXp8EC60s9jWFnu9K/vyG/6ijmQUzY4jm
HY+E4Vzt9HDnC/mVxrqT5WPr9CvjDn8lSVPHVJbog8pHQbCXqq4k9GUdNuTL/Nvz
GRSyzJ6t2IvQOPqCpbOBCAgNhnaK9pxET4hANAXX0maGFu4Czn88aIIEgq/Kta3Y
xzaRnDFxW+E1fSJdRsxYLQBsbbyS5azmtpLnLEGvBChuaQ6aMAGzLWEMKISXk1aE
6A7Vx4jLt7D6fiHU2k5ceCJYNfGQEr4MzJ5yZacccNx4JoyjjdncfzABevCu1Ngf
soFVRYAgrOXAeInkeXLUGpS8XzwS4/tzkyWKy2ZMH+xYfeklWWTf7TciHY/77cNk
FlpB4RzffhuhIrtt6MDcsg==
`protect END_PROTECTED
