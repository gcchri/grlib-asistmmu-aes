`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nENqJ1xyU0d70L4nvlKjHX5dKOAOf/p8nG+87c71db8Qn7MZserfZLnIxMZKppzm
nFCwxK1OzN7WKJVHSgZzFNezTE45LCebfiHNassg3ote28UQPdeL/rSQiOTmeI9e
gt13gexD93+2ThpaD1CA1TFYZaPKQUmWSAClfQYHQZqfIo3SU7TNLkY7FHh+TN3g
2IYX6ee2lyzwzByTppXI+8wsf+pcZRFNwflqVHrOeKx2OQ0pb1bKgC3RUJvNcLZf
0ImOZ+DC5iTGPDiwPnobZ8cPhNOVX4gv4kap6kD4ERaeF878MYbuzG7SZAYlVcUl
JK7oGx5Np5W0JDT+e16ejVgNpNCD7jC3q76V7pOUpxeLyd5QKW+Eq73GTJsW0Ohi
Ha0boE1SFAyjBCnTgYE9aJ7mCsFghkl+UJdGPPZAU9o=
`protect END_PROTECTED
