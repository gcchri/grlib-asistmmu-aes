`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BdyL9fYzyQnZ+6nEkokqAOMt5PtIMZn2m7rm6SfDAJZs2uIQ60KALafahRXssoaP
7aisHE/FYb6B+3YnwfTZW6NfN+yG+t1hAeYqaNaxu7roTD89eXjtiMsqX8JNzxWk
mqLYxaba6HVY7KyFFnAYa8SxiU+RObGuX3l++3Vn10DHHEyDmJFBtukHMbbDl/eR
RERE0jhW0MAUMMl/0HGVtSX3indpEi1YINwziKe1U0XG3NEYFURzMPjmv+7pKU9T
`protect END_PROTECTED
