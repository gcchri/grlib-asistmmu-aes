`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TGAdpzAIyZwj4/ka5iCPxvl3EDO0FDjzkoZcXROPguyhvsoEBAhWXno7PCAhLVGf
RqXJSCxd9HJcYxNmIzDewz5vQZOgRblSCNT8aWg7k+zDlwik34gdht06iCfFqDoY
HxTSP70yoa8pDO3VtiWoxpxECmMkWiO3KXxzQzGIvIZYEpCMciQJQE5WuOeoWoig
ErKxNYCDGGKtyPxvqDQCyMc7xpdjs/I3sV6GkmgLw4hc6N+DLjyOpIpn/ysn/FaD
Wo8hou6FoJPTeOJ1PkEXaz/M/y2kyjUpcy56kcP4Zm4yfNBWBFXy7bYdTMUXDvZJ
t5lyQ7k/ydiru8uwRZrzgiaqKjTls4l5rdkGYr/S4cBYaRPOlYIzQKYA2Rw4rXrV
uFCO+r6mhWPQVlGA2X+mNvuQLEJg7W4+09o8W0DxnzDwmlYgYvXw8ihX/Ys7ZKEb
6aKxgTBIWklHqc/JfsmbomMP2FXkRvr+PJr9RU8fiZXhFGFOTRZ8kWz1lNpMpiFA
iAVTYQjxtIv2BWXMsm7JGmGTzQ6QGfJiYSkysRyzWd7NuwDV+4pTQyEj8P1mOFvM
YT/lnYTFFPoshoA8kZZly+IYL2OQl5/dkLY0dBtrQhTRyDyIHAc6w+5OCdVdG1kz
crhtLDdY3OOtna4Wq7lYKXanET1b1U984/WFnDBJon0cjqHX4MIHopG0c3RObRTL
SooB+yyCjGoh4Dy9HfFQVWdEgDxkLR2suH8bSqnXVrsvu/dYSA+XqXzVEDuB+QOG
+8UU61/7+Q5Gy6bPYiM19z4rQd33TrsMi1+yBfF95gY1bMgDJKA5O7eS+5iZUjcj
SI4iaqDuFCedq09IH5ZO+Q==
`protect END_PROTECTED
