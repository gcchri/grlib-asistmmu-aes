`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q/MwFnVkgY4I/sSZI6L0JYG473lzSATKmFGw1kheKqx9DnpwHdIF1U0ITDGSap6D
ixNNrrO3hMRkvTEgqPfkaK9opt7mWeIkrsGfGjaBlbker4H0eTtEVECsPBcE5xU3
ueQONNQmb0LHZ27ftoMpV4dnBQTLozqxENy6222dA7/g8tv88vWHA6v4l5ZUPdIr
xED/gHoGWzgjgX7Ma/+zHwAVqiKNkNIHOvWRyv9w3yEjbAVeG/6J0rPK8qVDu6f4
MoXw7hVYNnVmkdE9k1nOiOsvU+wNoJF4oiGOUil9w5Y6jpPqP5S7lIby+Fu7npzd
U9KU3+cQ6CPf8oOT+YfjUi48NrQca3AEO/FUFcpUHGKGFlK9mEt/xCc5VUc97wva
OXVcdmeT0j61R5Ww1WIscomcus2yBeksCzdGU+twmsAAeoxQOGkVo4SKOdyIzg3C
8/RdigO4fa4BhVKNiKi6hyPgiC5uzwDwiQA0gRu0asKkHgKqP6p74LO2L6wY9jur
xjWV6prXmxskI+FbJmwUpieZMQeSapZjbMv/W8Q0DgDvV6xANMKI11pbbxAi4NIS
vfbf0Dw2mvyu3KbE05Klf/R44JYMjU+JZbpvMH+gdBCHqU7Z3W1rzrnVqaSGtCJ0
ijvT7xtcyBE9uGt2aWB9PEu5yprRivGwaQwXwCQGtJA2MKa5QI8n+bOzWUeh00Ls
SVN/1ogt9o0mFDbTEE/J5/DtSz6RPbtvqhvoONrUh5bjvVQZWnZH8TS6i8qNqojC
E6frxq82n6BPIQsqKBP9+bsQRggs/Fws/6O1eyxE6ktrWszSW00W26jVeMY3yUS4
4qVxYqNLw9zA0zZFwRTWWKyyinEFOhDrvQg9e2OyMjKnY5Xw0wnPss1K5udHoOp4
W/4V+feJMuIBN+L4G9vGB6skYkICsBVPHAJqRtMACY5KBUbYHKblhFarCj6RNuF7
kcYCIXYBn9rnWbtIDUFtsgxhm7jwwwRyxdZSUduaquMwJa7lx1UQjhE0O3H/hSk8
HtSUb3VEHQG8zszzLPseBGt55z0lkh8/KCkHrqrh91zYSjVcwFJi10DlU9RLFrr7
n7XUqOjGPexKV07YQc2QQwEDOgn8SjeVAAdH3IJEpTNWsy8VmM7zTEnrLDU7SOl5
i9oT5yQrGeBaBc1QP880dh8xE+7KJg3T2/eTRuBqyXrPzeEWPiNFr4i7VLktZ435
ybo+qrcfOK7O0zzVqEqPIW8ag0ch+dXng3OBVpWkID1u42CP+hgzvn0yN4vdJ0O8
WAKBfxSx2Zrd7bAlnbeH331LJwSSy38xlUg5Q8G5aDcnOi4jkFF+B+dXphwDemjg
sJwQseQq14c3ngMJKzT+zPI+zDFG474LOWlcWnvToqiz4SFkU1h4dpU0dtNb0t/W
WEkC0ealcrZ1pNaWi9XtZ9wDF1+bSIuXHJWOgif7jGlgWRuJP5avuOVkD+yGlbGP
8bEw5K+bCQ0ZMAHpRpDGUVeX7Uda3Vf6Di4qZnklvX9ARfR51Wr4k4Dn9ZWmB0gY
eO9XVsKhP9QinG5QMnvyNJSYoIkf0APs4zPHEuXVpU58TsUbY9FLrgbuqTeQyz3F
vcpSpSbgMFNCzuMzsWDuMkmLStFavdnCHd3PxU33jgP76D8LjVSEw5GHoJfOe9Zm
gnXZR7sd3nVF42GB2Q0Iw48LOXrdX4GT+ztkohy163S3BtUZV+YdI3T3CkvodNdX
HmS7wVRYfW3RX75vZmWoH/GPoV88nGK873olWqPP1qAh3c90wW40OaIsFrQa5peJ
aYPIoyaNo3t5pKiE0UGnx+vmHeiaml2bq9bpsYH0akdIvWgZPHIZEbECpEfQfG3I
ClS7WO4QxKmqgDREIWnyLLMjp3KbMCg25S8BqWiD8GLNJtfnpkEi8FUjdvT0VF3D
bqI9qHkEbX1lQ4hg9gwv2WXuCED33DFs2W/inEsPH4r+8YObwW1RLY5oa1GO4Yrz
DuS2HkMYrU7h44yWsrHzBiwGb5hmngEQ5zbiiTEmqb8ujp2DgSwam2sj/by6bKjq
k5HPkbTu640S1SvKJfwqmkY2Mu2WMlAnewzdOd+0s9a5NtFK1qoclVmN7TwttNpr
z/1ut1jrYG5YRk08Svf84bITgh5gQmuIvRVBXisVxt3w4kmuaRsZ27UlCBvcRpV9
W9vIbz8L+uRQSmhlqBdj4iP4C8VGwHZkxDJXOJR1iqiWWPGhHNUd8lJhav6eWxH8
dOLDQjAHvKKyy3iy+qrmpyLOAzUBlSJKz00Rre594oC++KS8h2z941PbjiQy0iNP
qI40+kzXbYDDvnamWMrGZqbhWoBygdL1bmZq850PBil/INq79UVhloKMdWeWE24M
RPwwba4I1Zp5Qp1Qa5yxwK902i+Q3hm4Wmslx7hhAmvLiRfC5FrFqdVQrwz8EA5C
OQo/pfKATw+2NsCtIpO2dVwGLZqHaTfREsH5SpID3jDjTMzI+aJagqK10FCUb+Rs
yNy7qY9V+0cCASwD1LrjYb8ZPQM8y8N1MPlHUAnQryM7iK5LiqnUhXHsGLqDW802
`protect END_PROTECTED
