`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gBtDzn/GeCPr1zP3Bo/ur+jPa6LJ54P4bdoh27kN3au98sC4+F4QOlPwdIb3csGS
rT9yYWPZQoVmYK7jg3pH3qknOoovKBDvznkgITnxmvp6r7lABHsOEbOy5wpgUzOc
VIauk1Jw8T2o0CK/dDoxbkj8KoYwhZy2dIDdY1AvWCwSp8QWRf1e2h7tPDwhGrD8
oZm5aYIFrnttoz0rscAr9D6fAD3Up/IKHCzuhEqRqHxQk+J2g7yZuoJgsaBnCMlN
ske53KUDra8jf8DdOkJ8vY4KkV3QEzXnmUTy4K6SrGRkBhO3yihBM48tEAo0U2ir
+pfX0UX/LSp2utKQBEH9qF4K+ZOzhYA4mfVbteD8KINpt5IlXYWgJDaAbdr/ncw4
iGpikUVrcqtriTfh6lhEjQ==
`protect END_PROTECTED
