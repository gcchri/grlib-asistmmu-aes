`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f9OM9MRpGxvX2UC9LTBsxNufUAp9AEAmBWhn2Ey3p9FFieGNelTRSHe4WhnWZcsV
/WXW4OGjvnk6CT2kovO5qqN49PByREeofvQ08NuJObL51mcTRJmTY6YwUcfTQudZ
LCYI86PpOMSf3WP1LdalQxyOlZQq3usNp57KFI+eT0vEzL9BYxkzCKNvu/ATvkvz
AzBQJA1dY/SNcJYnsA3T+jl4vrYkJa/BDv4lZ7W6u+uaepivPVLVmUXH8ap/X347
JAGuKO3G4EE4zdH5Fhq/zNWCYEEgx7P1zsKlscen2pA39DQV2GP3obvpbAtqpn7N
V59wvoGvvNzVUn70u/tQJhtDSdUzTVe8Z3D9C0FXfaiSfreU8+cFFNe3xshaVmZB
nGHX47rn/HQXlwEbqmUU4rC3crp4awE3ledfEwyt+06T2kTtHhGUhbz3Z3Z0QTcM
M/cKBD/hYOZt7S4V1DkJvT+vimsHVT8xD5ZJ6Wmx1erpBMsn1/ZAuGm2OGmIT9iY
YVu+2DBqUNCfYg1zPUQzc/Woe4nA78t5ZqxsvPsI67Iv2gpzVahoHsIgw2FTUeHf
afUhwA645yMs8QtknisKz1t3QL8Zl0Ksw4YQ8uqbd2WE/Pbasy/W5e8vDhK1H2Xq
XYd2gu0bAzZs4c1pUKvJvEaklRnyGhbUbqeOlsVY8fLSXjFiifvOSXLSgazaRvzm
EWQiO7HBBIIL8P6IuKkg32TOsDYwV7u7Ezn58obiXQCmjTBWt4M0OKq5x+1zoXce
8HxaZhG2ITz4NnutdhP+rpMZklUb4nIpSNLhtLrWivkdPWM7RnyB7n+REpVKWnb1
o9nev0smajI7lU0rZJdSoVu8pcNrfS4nIOccRg0sAM1wL0dufxu/D4QZTv44imDL
ZOrLYDGGA3KGbNwpBPCK4GkEFNW34KVyiZiO+YzPBOKmyZqNjLk9pEXzBmdDJYj/
NmbVFU9KOqmRLHyasSbKPiRyCyowM1Z/zgNaQJHyVxWrMhZSgJk343ldoFVhlwTS
5SJvTDPfXXuGsQlZ7GhVKiq3YimFA5HIE7b9XLY5De+KfN8GcM5AnaoOiofEji5D
h+cAhYk8SQ0+XO5zVpMu02Yyf80uzZcpmQS+b+S2mjZAzMNb20Q8i0Lwls+nGqO2
I+AWOunTpcR/ByUJPvYnHkBCC20mZeMUZO8EioRzpL7fJDqGn+lgVT3hipNzdxOT
Y4lvde+q8ZsgXgw0A1XNH0WSIqkYC6z72xBo0nlde6S7Aolol4xHQILZ67o3EG0o
HlhmVUd39FZozGLhF4Gro7/4H/X5hA4Q10T8ub0RPdiJTacoMqCb3ZlNcPkxPrXv
JF+Rk4R9igtGWvDnYiqmWdN6narufRXGYaImttK3hXaniqH1TnbBfmvTS3ivAhHA
bjaKBpO4JIr4RlA+WFbQeOBqQj2z0J6nqT1XUe4aS1QfeL1ACIa9rBxlhlNKsDZA
PjDNH5h5BehvlXiKQhm7yTGAY0u3+C91Mhdzsok3aw2SQ+zq9Jpu2mbuJ1Yf7Nlj
Fg0mYix+BkCmb5GZ2mEJW7O4sXMXTumoPLYlN2wEmHPJ0TYHle8brq07VMT0LbtJ
nNU0qZm6mSo2H3tf7NAxGVUxXtvDOfpCPhVDEO2VnZEytu0V6uM0TVqwA7JVqdfa
hsmWH0HbcT9iQDOuadUlWFsajLVGDaPbEaNQ3OL2BiclEIR/g5ozPeIfkm263j9i
Au28aR8QZahGDcOQS66z1QNPtfYoJ1Ob51L+R4pNYcRlvZhIyzPrOWJzdcCvdbK5
qAjQ0FjJYd6ypFin8cnrXqS2nfMKaN8Ud2T/8e3+POAOXWo8vwkhW3NAF/A/A0ej
zWRY03n2/eyOqGXwHbhWfvrJr4yLjhbe7GzBkai5VZ1U9Dyeyk/fMyhft9wOv22r
jAUVsYPAd+o6utH8E21si+TDOES0D0kj0z/ILnRsK1pevwlcbbEwXC6tIvdIdK6D
E6jOXCC6DCIL1X2GkaKGjTyCJ/i6icDDi5hVWUEyri7uXnfSf0ZWL/qWt+tqj3DW
+ag+XZ3/P0/GjuftouXyxQGPyZjznbVAhSFwkg/rASx0locoqEE4HXoEifjsMi1F
Wo92eJgZ0Q3TZ6tEAEIvIW4zMqyQSuh2vDKtOc/WyqymqGnnHfpT9rTOSIgnD81R
Zz5K/5CWk2rYPndaXttWSKuU6oiySLZLUqomxjf32JwKcLJIGfi2ABRBrm3RYTOx
w6WYtKyFfn/mW/bfpXjYasat6Q66wtfTy2YgLpnWbtRd3nrzwG0nUZdCyiPyq8Us
fccKfRMneNjjbDhFwKPrfbG/48fDKR71lbLqqmq1Xho45qIU2fNztJZftRJddl7N
6xyVrW6gDpmtkrZNZ3pvtWXsVrQSNtj9WOI0ogbHVFk=
`protect END_PROTECTED
