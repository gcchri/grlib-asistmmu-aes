`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iABOxbrK/eGZ6xilMU8g/xqGjlfzy9IDsQuJ0HJ7vGZ/ruiydTy8BMvzDZDLmr2i
EoDpAulCaMwjgpiKT7tWw28FG56waKFY2/5vyHXhHKGkui1g/TvlTMOVLlMPcpGF
M5/EEsTBmbFJGT1WMfYRCpWFh8JPdF5bOn0zFknzQ48HmwpC8uaxV/ecoyo7f6y+
4OAgMb0fZ+F3qjitqPzN0VoA27aSt8ijvMQie0f9KOgzqSkvHMzyn0+eMJyWpGzF
VE0njtyPuM6sL09TpDbJI1v+fIVW9Q5JPXXDz2/7fLXHq0hQ/g9eJiM9vUZ1Olrq
9r7EqGSklKWy8DDigW6Z0pFjKEULuSFjIKyvDU63Dfm/EcCa8JhtWPFbzkOsNl3q
VtdoVNzzFkFJbrBUWO0FIg+DsZssaCHEKtLFZsp82dE=
`protect END_PROTECTED
