`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
weu01+YXMcbmzICTTwWryAbSI/k5ZQy6APTkkeGjiGty2ySlhY+a2djWNuLtc9Sj
3MVb2QzS2T79uS6VIH/ZBtWKurjeXq8YetGs+kmP8EKavaAUC8YQWAVRIyqEMUto
0KAiXwvUYEc83OPQeFNkJsulTfADBQSKp6L3S3LNPdhxmWz4lzTnT1on0a4hNcuB
JgQadIf/YSbfyJmBp31mbiTP7GLlzbPcNqdqjhpDKpsG+OiCg2U2IJuqLdamgVjE
6J8puDQunphMyhYywwNT3U6PLryNnLF+hKKqRiopz9CjWAxhGfJKd03EtcpVqOiY
uKYp6sbLIMgNzcwc5xJC1g==
`protect END_PROTECTED
