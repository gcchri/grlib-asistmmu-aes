`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bhumSX7S0OolL2+BKTFEU5F0uRXebrlGzY2HVfR4b054Ep7Un3jcwKLuIOZsYiiU
O/x2HobpZktM+YOfC/MqKiG+REMmtHTsE/PJ+AT3KABxOvO+9Yoj1KmLn5M6PW7P
vzRVCceB4hVnvHzQSMlbGDe3zp9LYLJ5ZCyE/Tb/hejfUGsMw6GFp+/SIrcGlRBl
CyCTa7510EFqc8XRNnNCPQg3c610SsilQylGF7gW62U7K7KUmoYWrwLnYiURojaw
EpQ0+Z2PRyKQKgUJqNCm/GuH7kKmbgXszQ6lAQh3LYDNhyYgvQe1G5tsDErhy0ag
IILGWS0iSRAaK3Ok1pBiEes4e+y82zw4vJn41SIgcIel2JaW62K5jSDA4vK7a933
t7WWUemqUzgY2PVYXhEhgbkLZwVLY9kpZffhQY2EpZl2P3V9gnAn55oX/f+pWmkV
9FA46dktam/WcOTn6xi2tdR0fiD7NFBHdrlUmlOeg+kmzrNpstqKTEmUTEn+v0BG
`protect END_PROTECTED
