`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5rzcMzl7U8YM4UHe27LBeZpZPC5AKmrM54rBROglRvAlPlHXHKMUQ9ucdcSxgxm3
ACxoGtBFnV1BtDJOsTHnm8pzaERlheRa27rDKAt3ho+iutami/0SN/LWxVDTvVi5
epvcDMURnTEFbWWNIcTL9Ixntw429oKwXFa0aVdezFkCgtNVW/KUgl5q5+y41G+Y
UGCVFh7UgQ2EV+glG4nI6DAG/dcy3afCkCplvRVzq05kxAxh6iYLn9xPCUoZgzqM
CYZF41DcdNGoNQOKjZ1rcBfLeRb8v+xsag19RsD0j64=
`protect END_PROTECTED
