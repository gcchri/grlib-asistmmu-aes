`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c3Kzmrrde1v6kgKXu/AFD+LTtWv1ygB/RzvY76LuWviaMlZdqZ4a0KvMbatBnWVj
GHsgo6pZ9zKYl/BvsEGNhwj9mWm5xfEw4kaGMnjuoR9xgwMKB0rb4VIDKC/05V++
lE6i9fLCbN8wP6hzLpZLchrknnNhdx78Hcxa+Mxzdh/lSyFmRioP2GCtIBmtF32z
QxsBky4o+hQES4n5/qr1sB466BMA6AjUAB7QVF2wk2WpuNN5y+gyHX85oPM4ICyF
52RIjTgBF99ie9Dz8xtrq0YDQEi1iHUNaqBmdfYnn3eXe4Bu6Wgjlzg5erOQBsl8
9yh4nVRoUyaCyPn0lIsSHyAHLzeYUEJoS3OjAJfV8KLWk2blQVwMngtFVBDaQkjD
knA76xcyI43NIVglyOiJNW80RWQltwuDCemjGn1DDC5mv4H2/d/UZQ3rMnzBb30I
QPA3TB00qlFOIgdfG/dtsjqQAvS+Sq2GnWxhxVlXZdKy7GguWJyZdnGFsbpRfPtb
1g5GCsBHPR9Yv5lXBz8ITQvIxKJibO6bWKRDdFsdMN9R0cu42Q3OAfls/c5llDYk
jY+L4xi0HHWk65F8fQ4QVrGKMRL3HJv0QbDg1t6FK/T8wQ5fyyTBdTw+Xqe7O5Jd
`protect END_PROTECTED
