`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PBchN0yvI55mhNeA699zqM8HssbUsB7JUXNpDzEuBHPbLIyHIlV0fThvZUDkHjam
Ld9jl215wfTL/ailuS4X9WTWd1LFiZ7OE7M1AFhVsHe7lbW9Ah6st+xy3r/RSC2E
vpUiVuJnPDDPOkYiE75plRMtU1fMonITtHpf26R1C2g5gAJaWBogXTEvxJhuKjy1
p87jsdv03MmGFQxdYIY2P+qCUOAV4phracgoIc+9vq76HnmCYDkOpLeGCFuRTnEO
qoVAygI/ncEQdEIrCbuAYVOaRyVayGcrGW+G6OCZi/oJvy8/2PcnUWmW2ttAlcqz
TTCCeJkAwLxnvfrclcwP73lUZgt1XNZQGpKiFlF55R3xs8yv6ga3ajMCNYtwfpel
4b1WylljDgKT1uaL/yMpW7h4Av+7suSgg52mI0FN9r4Awmt0JARkRt+sgn8ZXojS
z0bHGkJ4kQfaSStZlwQXoBskgI+vOf/L3YD7UXdwlChUE1B3n6K2f8+1nkwEUEk5
fcovdMHRy5k0Hw/QwUwQZC91f1Fa9z4D1TGG4Q/A8nvfATmhr45WOrXn8l344m5X
DlfrGpI9tngm7qAyiIQLPNexbetE8peGhFb3kIG9mI3ZDU+7cwASPK/AvolcQCxO
d/bTsraT7VTM5mgtu91sgMfHxwxfQM/1V7EsupK+gQBzfiaD0BMXAbWOg4x6AlLz
BPQAAS89bb43u932nLDyxBBbDWVTkhhlfvs1MaYq1987U+yh0Z5fVLu8cKBRroPn
ZNMJBZR610kzf7mIeNq6kVWakMEtO/Gang6pyo/kzoKtS5CMqZln8m1i6vil5D8+
x0ZlB8caI+vuf8t/S1Y/fuUslM84yYtAMtFHqtMJNG+SY4lPt2Wl9RmrUkr9SgMA
sAjcHDT6TYZkD0Fdqg2SfzjD91dlRQdaCSN0QDIi5QCkhZQj+iUxE6ylRKtpM8Dd
lOCOe+uOrTyAmrglFE4TjMLmJOLueYubBBCSNAGDNW4L1toEddt9uzwi7DCoyQIs
CqMTG9XAs0G6x9SobZPrC0EsB96QFJWVfHJgSojonCO0CWUDHqmlEnTThHP+QFsX
Pa7MTieTSi8Q1ZZBxRA4OKTJkv4qTdJNqi38cEU+PKSR/GLvzNwR1+nt2ZVeTsmt
`protect END_PROTECTED
