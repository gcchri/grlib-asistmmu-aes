`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rRMD6OCJNBbLKseM/Q9JlIDkbzmDLIlPs1ktQi8n5TrWNrLqdgbrdGvtuzk4RhWZ
MV3wuGE97wLvAmkRKG7V8SASdEvc8zvRFYY8Ud3cbIg2IU1ECb0SVn0HL/p9oNh5
ixTnFoFOflS7TVvwtaWpML+ned9KYmsi0oRiorl8lC8yEV8i2tcJwBFwQHurOATC
llbm9wLn5c/Av+Ylcmee4PgNN+3my4TC86gvz8Akau3L0yiMorgvRfg4up4KFYs+
0HxQBHz4/hXEjvpsEtYYCIzOnXDAH2bZPNsF7f0sGGYXb7ANMTF2FyS1Ci1q1Hlu
lMKooDoiekGhcCjtZB3e1QfzevSdUVRqkJVkBB9UkXuXUfxrgsjG1CVsS2uFZWho
nNQ9SEGeLN8XKK0ZuDVDYQX8YAtKwRQed9hYi3UngcEDf5ofkOm/v4fuSOZfIQJV
`protect END_PROTECTED
