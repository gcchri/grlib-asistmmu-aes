`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gmw649oDJRTPD2H2wnjmyOu14AOFDC/uoZ8eB9nln0pFp421/UuzQ8T/Dxb2QJ9p
55KsIKbsvwCB9+bnNXMc+evA80DrBd3in9Afit/YNRW4f6+sAjmwvwIBIZC9xF/a
pYSFDUw9enR7inJ1vckEnitR1232METvRwQK3b2Bq+IwcP4CRVT14t1fHme7vj91
83o8Sxo2LOGw24E/v3rij4IlxGctISQUrvtngEGgstB4hWldIfOXEhSNlXrTGMCv
y0LFfzXnSslLiJgK7Dmt/FyBwKBo7hOJpeK+Lq1kldR8wlLUNFeDnaBNfV2Vt+FC
qAFjWZK79qOCFsjilohlg4IxwwLJyML5XU6aqbnXIM2aJCshH3M8Fkfm+NVTctf0
1/aT25m7PtYzlUYCZpRz50jhWqmSF6Q9Vxj0JMkzyK1LRJjqUBHIT7N6MpOwpT0r
6+OFojmCB9aRUNSoFdlsDCtf5QCnOVYWy4wb1GZZ13fNRpdtsRzqeqYZ5EMhHddu
NN11tWcbszIhYRSXzS6suFm/eXAA/k0+kfstkQBxQXXaFEsCW2j7RKmQQpPh6MHi
Us8VmnGLkjKOI8H9/DF7EMC/o4awAOi7Aq8EbJnnqz/6D/04QSZ+QkHoor8PM9lU
WENxTVdghgDQdTgN7PuFPgjnEDSR8i54bmUZsTZQln8I5bsEax4GyshetgO+nDAS
zT+m9d2aoqhgGO9voWzCDsUKuleLslJwEbjQQgr6hN1jTrrQwHxnIZc1kYQOpyho
kjDIvZSUWqPy2u0hP95RAAbJlK1kqEC3pczxq5fhgCF0PEFWD+/c4YyYzbejN5jv
Acssn0zNgBq6CrVetr3Xf7/Us9XMquTdkI+qesYxCxd1NaTgfds1AnFtXxt9r+ij
iX6fRhwA4IKif3+3B/OXcTEtp17KndZ24nTr3SCTIBn3eRaY1IRJEj+IyMCiHpET
SmPJJwIZXzt3Yiq7glynEpyvSekyQpA09aC/98del5ZXAIUZotBLvxPatVIXbaK3
jMG2cDffN/Y4EjAk08SGfx2q7vujySxD89NE908EAI3inM1mv4RKX2hzUCPj+TGx
yVttQESLA6HECUXTes/DSLi73xdQpBZDtuUBoFEJ9a9HX9YT2yYVmNLoes8pJwCj
EaEnSbl2zW1+sstgWMck/SJ+kXZV/g4JizCK1eYB8qGGaAZgmdeyvuvs0j1BIfMX
HGDxnbXtsAqQYrj8n6EYZQb8guNNHjgcSto57MMYoCwF8CdwGHZyY2J10aXIajdo
NWX79Vjb4VoaJA2fF6u5xkyr6xmBmzFC3yGPaR9zbHxbw1urMcYcPum1OrrfALik
1XkAVCIVHbtBlav128qdtbR834U5Y4BZD9t7nCvCeQYx3EUQmGbjHEGL7fyFhRvc
xp3GNeZ3CToqOV4GLoLJs2o3dvRLKBvVfZY9Wi7pkXrxmBpwyanUrRaRXY5F1K60
3P8PMCBEaUDTPRfMkpCASKbde6fx8op8yNyskOfijocKNIVxF7WRcMh3CrOnFZ6a
QVtn2tW4NaGOevGOPBPSS5IMPUi6ne/3PIJwY7KpZHkfvjGvZNTmiSmunnscZlmH
IZcfGfZvo7qqyqqBwO23AJLavjqlNXlUIKjW/6nxasFcTJunRqJS559Hht6R3a06
tXd7N30HUx6fwiGt4l1hn3A0QQCDju0aFByq4q/+tChEdaO570lFn3JnJ3W6YLA2
qce5lVyr65/p5yCvfvks7+aROuFV9BCzuQPeWmmyB3RjjV4z9Yc0Sd2UTRIqlfeG
cbAzrRHU8v2nnE+65VSkm4m/ZOsXoxhFVWYyD4JMNOZRPDsbN4XL6P/IJ5rkJvHd
EfFq67de5tGJpqLuRj7dKTtBbOj82raqqHk6Ba4BR1PtyttXih2Jo+Z+jH719XJY
03GPQLpi0FmSriHwaTafmrN4iUYxvUra2a4g6DCWLwaF2YJ2a1ocU28/ibcqCNO4
MwIgdWfBvikGnIlyRRW/fk4dpEcwyK41Rfzr5p3uNmN59XB50lfNu9B0BV6+aIpC
OxHBU61UPkXIg+IKdk/+X5dhv2yx2iy4mrPf7g04YYm75oVy2i53HFE99wngUt+3
dO59rKmFYtBeuM0NMcQHgS6NBGMT7DhGZqlgGIDbrZPKKlleaY1Rh9ii118ICKI/
SoLWK3G7lj84GFXdT+gMn1kqyybcUWZPmRrG3M42e2hZHH9ZSPWu2YYU17G9jjHl
WwtKzmJ0xJhWvhPKV69j/glt/N4ZqbdGr99juIxu4qpXa3oqMKSlN6T4xtT0eaTx
2jFH4MlDRIvHUPB6BNn4mAi6WZT0iLlw89e/phnpv11g7HIMWZVgjxTh7zKIZ5gm
gWu+EDszbW6YlKPFS3xXYdWAAiGxSbNTIeGP+SXHXiNxSbcgtdO7Ro6HGFsMcQeT
QqTbJxsjamGrAuYMx+Lo7aAJ0WT4Fxwyg4q/LB7dhlehGa1ufv+fOWKka49zctBq
WIGSdjEcGSv1L2wA18GWOQjVnluVc9m0H/LKQONDzr6xB83sR06elJQSW6iL8PW5
adgqXdRJvrV2h1mCnb9yxKM+3uPiTH3Uxp2B9wH0udZXOzwYgUEVzYno8cmkQ1qM
1A+hWZei/o8OLNkTVEgHaxnrjxk8nTgmczPNMUODZaf/hfyvS4TqaIF5W2+cpMPZ
EXz7hmYdpFm9CuN3m9m3Qpmrhevq/NxRfsHQuctWu+luEpLRzbQZnkVb6msbHvKS
nxqhiYZA3sV0bFT32GSaKNlmCykjP5KdVHRZgs9xRw2Kj9rm1b0AmiSy4zQg1900
eE1oLj/TqdxZUnzyO/uLS/kJ+P4vva19EqQ6Amtuo8M1MsJsjhwBPD4uAt33fWRb
bwFqalOJfcS98I8rTkyqlRhRGD9n29Woc935imzZKrBCYTTFFRhXcpHqQLRym/2A
U1LR9mVj8yqslKaDIK4gcFXL0fdN3GCLkW4UAH9Zk4yGSwv8b0MNwSFdMPAL85qS
Fs7FYvpDd+bbB1nvds2v0STsMd6s9Y6PGcCrcubyTKk=
`protect END_PROTECTED
