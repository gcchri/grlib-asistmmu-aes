`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4iEBnJYmW6/XIQKPa8cT1U9LvNcL23ee/25PZ9VhZXF70p6LEHYoat0d2xOq9o7F
4xxd7RyCmR25DEkPoMRJYlvt83qwvTbxkV1lllxZkAPg8yNcev/8OSmLrBoqONm6
mFTh2Cyo02yaVijHaF5lLJ9AWf1xDVT+yleFET+3fBP+NpzRYKwYlMAOjaWED5zm
ATfIgAw9XHM5dPDFAzEXaYz42A/DRo+FpELbtg9CVKPCKmcGIvoVVm7nhClaSz68
92P98DXV7gPfKQC/AfpvrjY4qpJk+JOkNtR4rA1We65bzuMjIN6lC+ms63QFGXTA
Am7dNooi0aH1uJHILpCLwfjbzS81V1AdVf8IL6+LvGFcnFJfyJTaQ9o62glnV7Lm
J+WpcMJepTg1x4FAVrWZtDAXc75Vm9z8gGdCiOnxWiMFcr8SHv2ZNOZmxl3lVsbK
wj/kZiHm8XFJ/1jSfIv6Gg==
`protect END_PROTECTED
