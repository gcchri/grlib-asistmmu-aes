`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HmiGeSRyXssObLVdFsMsveqB9rk2JZ5PGB1hYnOCQPmeXkOe8bviyoL4tzhPfhU6
HrazLSH4Y/zkJqJDLPiKZWIWCQ3Bf+bEIp0CQ6RjScyoPuZiAxD9/6IqqkWPMTWo
frSUC74fx2rqYkhJSQPvoFvP4wakxjegldSKIOOYu7NqAkNiUyu8Lx3tIcJPimC5
d+ubWWdCzQzrkGfW0300zXVNYA0fMefLqttN/2Tld5Y2FDlxc/SjszxLOo8WpN6y
lGiaoN8tUqD05248onFtx5aGOmV6iOA8p5BBlDhqzo9LdBtOTyEaT2YSSC1Xkd1B
LHmEwjz0JDoqDFnTR+q6h+zzKRocpzjRORmZ+NluGHIRrShhwwWI/OwGgnQIkZze
GlKzRnA2eGEMGHxuLlkDHMA8kBwtDyS2jFbuCPwn0mS7wZmTdeL/dmcmh6cUJzy6
TEtecIQKgAlKFcKUrXn5Bciu12o3VM+UJ3D8Gx8NFrL8Q46QD7symuQKvT1inam7
nioHZBJ6kMXm9JhlzKFjco3Rez0isHJo9oybJaFuXM1vlUW+ruzfVUUEGtQmI2sc
wqZIsqKLKwAV15AOwfxa/uRdpDbK70f7czjjFTdF5Q4GcviD8h4HrZoA9MrtLe18
9Mkl1kJ1XsYdqS+ynNmysYOknVLC9MSMxm1Qu0A4B79mOMhqTfIlEVTj9WynVNie
bLJ1E3NY2ugoHsB87akgk9mrzI1uJBhYIb1D+qccVbsMFnPo0cmWpXDvEG/ySyJZ
f1cip0QbcF4oO1f3s3CR4skFQG/z7bI+LYpRBDv2NwHUBs5tFo8AkCEMNwJRN5uf
WhhozymdM0bTRQsK9GV73UnkRr6fqrVNbYGoq2ruUpTfsNhza7RBEaewm9VovznF
KR4IylZ0taG6AZ9AJh1Gl2hJNE2mSQy19Zl4TYOePV8LcIXjgH3uBVA3dbReMtYp
TrAeR637STuzjxSKDjW2M9d4CIZBfwVeSRnPj71eNVvAc/o4o2nMqHVcl4m5mWrV
kwa3d+v2ZXArNzkSFMTqme0ow0rrCmLHXfC9ZECsDkh6JmnrUVuS3PjyQRCh1US5
SIQA7S5hdBP3iQMBpBpjU505qQqLQfHVr+wjVckI/Dfo0ZY8AkCsmAQfaPvXZemh
EX/ysNjWZp5M40loXVQyAzjlTmMwXlCer4tRzfmPnVZJ8kT68MUgkN/tRmkA0xvs
LTDwaPrXpd1svfBkmC6+uVVdUh7BYV0PZ1pSreucav0RLIUyiPi4ttuKqvcx2+Bs
Vl6kifhVqEVh+DR7cIt+cnqMOlq6v1gdZ0JF/mFmsVODuO6k7x3BPsjDqT+nRKnv
lLa5iaNNbvlcyxg9A66Ohim52Ux8htJW9iKD6jZAthR+0VkRdo2bECHd+aIfNqU5
`protect END_PROTECTED
