`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FThpicRyouIImUDDfyU4Nis5z782WW5eKyMhdDk5+68TOjBSVhgi18IYJ5W1Ggxg
VyOwOGzjVOHOXXaelNlBT2nAYdgqR5yQJbwcfpTDO7gWBeb7+bKt38mfxvEoHRGi
NU2qYU9jNY6Q6qeIlkLtOCe2rHiCGhRI7EnD/9TnFhP9thOZlVTagC41UJuqHHLq
ctSmDvSNJQqwDwxtL5kWb5hpjCgUdXOzydbQfBMD32ApcdOj4LL1l43C3mtL3LVB
ASsOTsl4rpIHRFSpWOxM5Whm/LRQmC0xo//mLCJr/t0=
`protect END_PROTECTED
