`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5RA3K4b1blPP+rDspnU9SWAke6eECB9w75B4oFb0rRiPINOD79lAWt01b12p08i6
L0FW+yXcmEg/AIx4jjmhdS+F+GJ6ZhYxOYhM/STNVbZSxNFWxA3P9mWjwDruSwq4
K/RKoRZAcu+gDxDNz9Eu/0gP9ierkbJifxA5qPOmHphHldWn24bfhlVRYZFpizDX
pjuTdMVCMqozJk05O6ns6UTWFZxZkPrSOEJiepmG1o73uZzq/6HsdY+665SCfl7+
/qu16SHme+w+uhG3zfbr13A/t4YMHrZjQUDl+7ShB7Cqk6Mic/JbhEmyry+SyKGz
a8JU+fwZhPJDDeekvo2z7sP3jk0DqBvlbrOSvQwmp4sFLKCSMC6aL8O/ByG+578U
Vn4799pLtdTK2nj4SuRK6DAHVknN52Yi+V+G375fIXU=
`protect END_PROTECTED
