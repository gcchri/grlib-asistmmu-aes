`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b1f/KbafOToaqxns9b6c0rMtk/KIn9PtzsrbQENFqXcHi3l2I6TlMI561Qy18DT3
MaMyH+CDGlRKhDUg1oHcviHpWLRmhdg2ihflLASsA4EI0P/7cR583VYpHZxd6SSG
nZeOH+c24mJv4MOaE4zbAv/M4ZJOwnLCBCZ2rDHuYGqAthSDHEZiwwoG06AON2NS
UXn4emZ6yjTY3gL4QdbnRSMKevRNajAX36tWTxBnIHwPKffCn14T1/bBh8ID8ni8
B24C0HYVUFS+e9RXerftv2NZwDhFDnA+NaZUCDkFPpqr145bGzM+j6UvJW2YN/Je
aKD+wzxt4O1h1RiH+dmMFm74MjwsTm7opO79kCGt8mSfwinHDsDX50q6qWViQc+d
jTZGDf7V37LF5OecUJSS3TQTSaQR+GUOrbA/875Dgu9nL/8c3nU4nquxMsWeuUNK
qeYu24j4B/FNu5m4lQaIgtPRNz9dK03GmJpoAl6MBXwIrBhfJrpvpi9aoPWhWl/H
ZmEf5hZs9jPUlq9uSaI/MXDzsk3X3GyYkojpWzSSnL4sDomxITPoaJgXfG5DuXOJ
rtWxTX5utGNWPZYZnbs/X2w8tDAU8p+/WPKg2Es2BNHE2KjvZ4xIc0L2D2mDTbsE
7x2uSImvhE/VcXFWOehIgxo1IJkfXm3Ogi+pe/1mOlUqAdkJiXSAnz5EPGUsyrAC
CgktDwlxZArjLZc+wxloUQ+YCPrjVbLUFuxHSWiFsJUZpsyxRsLYlmU6Vj7TKYO9
Aecdio2fdIDK5fPoNMhFIl5ddg0I5EMMwOGhUJjGTPmND79oQleOb8U2nPMo986J
oQk7YR93aG8FajhCuT5S0tYc/kJMMj/viQiN8qUpLoyaQ/5/P5eqFfmD0lpdrdfZ
TWCqBMZGUtcexkIBowgcEbbGc6hdd66bmQ0jAEs4yqpr9E4b4kL0p0zQpM6dqsZz
fj+5hVgYaIeBjx6hl04B8w0UJf5fsM1zQu0XYkdEUk695vG5D+elatUQTESlybTi
1VxlgYtdm1/kLDNnxUg/YcmyrZT0zrzgWOOyUsYP2+A6ooq6Hp2ANsj4lgurr0qf
oVjXlA0gf0YsslCPyg8wEA8YC/BVNxFXhZiylCzZAdMXDeUtFmMgHtUK/ozbIXxj
Lo4L9qdrpHQpUutYCWYNMfHYh3k0vZU386ZbfXpDqzc0jiejpF3EQSGFMUx4rEy1
QXkQkxglhcvH2LqSj8P6p4v20u1PbNq8uHkzWY53lJDedO2gNAj8zbkSV38yOwJJ
+zgrGa5TnpyQR/eyrNvoYMvIVN3wmZ8wUhyKmrvHs2gWFO2cuse5cqlLwg0ZqgH6
/XwU//58oVs5QfFx8HaSOUABXx++AF5SKsFjCPAyGLSSggA9wlLurjmpFOXEeBa4
ZH09rb5eub8n5ukK93IMIEZsEH0gc5l1kw/8mh4RuEakfevgkMkFXaSZVntzwdmk
LA9UK1uw0ndWEwB6JvZZXtVVfVUHyhcPKIG5oNjnhl8gtDaIL2ELD/uXz4gHyeWQ
iHQLKVbelX844jjQ2FGhDWnQrnmHsX+KpQv3TwjUv/uwGoiVjTfguffCVNvcMwRR
2x6abpQITBgYLotRM2IFY+FigFTZ0NhGXxgIF6rGxo/cqT54Qw8utg2MvqVLoK4S
iKaIv6iTDozIVRA+bpD2rEH3qS4JwlVYTzid35zsQp7iDisQQV5mkIyqVwi7mfCf
ttbbf/QEITgpQdX5xqNMEMmeRcewkUDjlOw5/SqeuIMxd3z4MRgD92QJqmqejDrI
GHLVdR4pDwUmvlxUGSFbOONjZAudleD+8RueBHZOL8Mj/u6Bz19DBqsylztYdP9q
oLwxLkFYMcKhXrrNUOn6FkjGlS+ZqWbrxvVA4qQAUTomTbleRyeMzhC1hYksXyqp
GlSUxPPUHMEykaqlSH65dWABjiGHky5XR6Sycj/Q3F0vSGHG/q/1dNJYfc3+nXc4
dxSQ1ZD28L6Xy6GXjHlvmnv405bO83SjDR1xdxCj/NeMEkmXEAytTzR4SqisFExK
fz/Xyvp3FRl7Ioq9XAqLm9Q+GjrUzgRQm6vomUyulXhvaFmknzfI7B6UujGVy6Z8
GNVgNXI9kBfD6Xuc0yf5HnASYHPgPE/8xnzhmoSy2IQuxR/tL8/i3DnKhIJ9ksYs
yHFAK5ItULmGpz0eD0qiP42JbaXWOeLpigEUUB3t/AMWHoUQG8MqNG/OghjDZq5l
YMahJKzjJv7lX8x+e4RWmfKUIjd9leLScK2kmvLp2mvA9J3qB6tq+n/uxjHWlLfS
aomYxSVcYiot+3S+9h0QZFG5D5KTYuddE5mnLhdNZS1vxc91e91xO3NOwQ8+LLKX
f6PCH6jea1uGzgLyRajdxn3/uu+VlZHQjLZECaJmKMH0o1yg7BSo5/kglYjtO95n
rjHRRkm2dG97BxfeN2Q/sc2srbC4h65YD8xoMymTzpcLluf+ucu7DEliuvfNgnuu
7VZ94R5Q5nI4MN1uKlWHdq+qk0bdf2NGa7ber4L3ZQr1bW1G7LcVLOnyUk44cqep
EQ04wW5ad4H8QlMHp9NKuJXNNnWwOvxJhpxb6ZA5wFsldlNurUI6gij/eb3GC3kt
kd1sOewd76Rn3BAtJDKVvyDHOJzqEkVIUzXR4VfphjbhH9/2ArVWwmlcuBAvywyH
+gkoDZe8rT2zaQjt8hnwn2hv+E30EUWvtvUf5sV5tOSHyV9kfG8oG5OmfycINCk6
AQmWfazpev1v6e2qBKiI4t0N6U0G5+lDQdKRnjLBlp/nIRO7CAXnqZjVwgYNsWEL
CBROxSsHLjTSLfRy4Cj59uEd7d0Fp8F4RqKDCo9ShwG4HVrFaBhMIYIJs6lnlV/Y
B50EyvB0I3bB0koyjtUzxv4w1ltNBdgvP+TgStn+DPV+4qDDGrB4bxnGQBS2sKrQ
1MA8GQqc+OaAmHJuGaDSDJxpC0rTIFS7WueDCLbbWDDzT+0ExZl2LJpFQzysWPnW
YgrX8DSN8B37VDyN0SQQtmqrpzkmHxV8kzQBE4uS1g4otuvVRFgT/cSCm9YK8dUz
yo4tF+rB4KczsgySi4yRh3UjQC4zDnsCJxYzzU3AV2QzMwN7QVlPVKoswi3cOUvl
9qMbpxibbI4o0VduLAMVuFMo3wVwn3kI8517Q3uYCH5Fd+teaXe1gJYvgWs6Zgh1
OW+/liopK4vc7Gb9E2k4ikUAS+ZGZrwde9kr+RjBzJ36Guy4LEoqpnhX9Ah6n1RE
Hh6ZEuDSLuWdKbHB3cWfSRgDz8TaaQ/pmcOb3zXDohc+gPyaF4dTgQAbPFIOD04V
xh7hKiye3K1UixSPSItfg4sl6JmTqYcQQtY09eLrt0BvPVbjMj1SKkWd8a7e32Zy
rXewam3xg1uO0PFYM8UINzPBuviQGOBJGVugN8f75Uy+YAFh8NH6Gh+Cq9xzzPu6
UmLCNvTCOpBkkvMlCo6TemXl61yHVTX1C+x1Fnj2tgU=
`protect END_PROTECTED
