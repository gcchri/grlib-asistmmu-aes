`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H6zqaWdRb4BwEkM7WIOtwQq/NWBHkeoJQYWikn5dcHOO0lKEF+BSh6x6tgCXd1Jc
87VFkSwda9T4Ga9VzlGT6xicE08+Y/wkeHZiTXQ4l5FDEAGX3plTVKLBYvQwveUk
ihnxmGOtssQKuV+z1PAm2QRZYDZkavkC0J5Evn6Eocblk/Vju1g5ov+xVuKAn1IT
Pj765fYAJIas/LWnDQg5ojLq/NHN4ndeDDqtLeBBkPMGaTb9dHd/XpzCtcowZ8zY
vqhSKrk2sanYdMf+8drOlu3tCJ0py5m0u93vvFpIpR/K5pVxVwuWMRCMQwyYk0Ya
I4CdhZ2Awry+fNa1e4+fmdaYDBSZQzp2HJFemYXsN8rcB2wlDU18YF1gJ+uF68zN
ME9LATiXvZ3KXwr7fay6rWMk96ZkN76bkHGqvI01q6rNQQ/ZLXvZ6woY83jYLtBt
1JNqbkANoh2byyFX+YIWSoJKyf1kG9BxRbtt8YHzDoHjNPZhxs4LLEjC05cqP8NE
tG76Ca4/8eGw7OpbBpFzOkcUgVq2pquMHcZHefhWjv3dfo/CLoMtCtpBQYXYzPrv
rtnx8NXhHNMP2RVgEwsAUdh/GusiGM8UAcd448DUAoFSoCA+i/3ri59BiP1r0MjU
z7cJPW1DPVq4M9u/gK6itzkBEurDHyBMugqCBgrUE2NMqXGKer84D1szkPFIGqyk
MviYrxk0fxc+c5mF3CowHN7+PChibrRRNgwsPvqJjI5555FEcnXOEnUhiVi/KwGE
/8L+eYcZTsKwhk7ciR6cSQVy/kCmlKjadGK+/iI6KxpJIiOdvFzoWoiZaHjrCqum
00+L8lHxDwYjkAhvM0a/89ngw5P5hjR9sFlbLABG/hbXqalPvrdaJTot8Ityy27a
62kszrGrf2aClW7CXtTM4XmS6+n3TLEs1RJ4zhKR7+IajBMQKO9/ap8nkuXO5pJO
KtC94cSOYlinrM1ySrcOwFpIJQ5xOOx6J7IIwFMSwjwP3QMeSUDbe5WvHpX19vFO
keBjIfM41ZRJEuIQT9FbmrH7BLpii1kVS6yRW3bN0k8pGjmJCqsUy5eCo2lZ4PkX
2dcMonUoFmXzgm90zt6rHbZJFKpl3vzCJvX8SoOoKG6TQw0Mq8Y+ZeWMwdDtLAmI
f0K/R8pst8adlPkVuryrcvz3Qf+Ax8X7ZlIWnSxtQRdV9ZKnTRJt5BzoU5LeYJGx
SLXjPJ8DPqkFmnmS6ba6BVy3oQhdYoxx5PDq5PMKL6XuzvlSqm5O5XJpG1+nlCUF
wy3Fcz6iVlMOgw4izednA18eeC0FAQMtEiUFcS2CSerg6y49J/Q1xjE4Ni1tFqKD
KLqtifVDP7ggSLpna+szJmpfmqysVYa+mTVC3QBiw+JauJx9UVWXfF2X9dtZP3xl
9qz33L1iefCd5Esv2KT536Qno0U/69ckYzwZdm348HtJXQGPlJ1ht122OoG2QxK9
yaybhENWpAO8ejw19N/NQ77sFDy/s8iMIWPeXezlcLBGEaWVXXaKnREirSwKlmoL
ASIr9p9pN2PBvepKc1W7UgrCzlozBAbsUJyR0Ak0YkJr7HuR7YMalRfIx4VlY7SR
mz+WnhufIArTMXCcmJinp+1jITOhej8I0qGY+Kg1Tu2G4HTYkXovhe05811ka1is
FyuF96skIOhwLxYkMMeXRcVGgnmV9uT2QyraHok4fVtf5ncZf1Ktvgo0aJJY43d5
uOf0xZoNMo9C5xpUXGb3wb53pNc+LtqZHlGhDBvEupWFoMpKeEkJCWl7+/36f82o
5ETuVooVayNYKXbdj1gIU7FDq2U+ohHqBzCPviV5mVJyCfQFSjvFHc97py7rE+D1
9g9cupLqoqZD/W4hrroc4inyU8dF7iYPinsgYh3zE2wTyVCnrSdImPZnrDaK3rP4
bPdaSd8L/kao1kQkFTK15BeBoWZxOUOYbudwIhtzpK30D+r4+OZsb3H0lKEhe20z
oVDhqzPATkvn9zmig9UHiGjZkKBHxqfbahCVMPlTLmvPWstWPuUHGNRY1YrR3Odf
pux3vKwws0UTE3/q+ZJWBILRurUvYVWkTVqh5Tez6anodP2STBFBTPvrllZkvdMI
NPSP+2LyoUqCwssXHOCB745ZKM9YBaQ+gKtUprNS/dY=
`protect END_PROTECTED
