`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f+MDg8wUDppWJw89ny6QkUoWgNqM6ddYrQYcAQbFmA4a3zAXeYC+0ouqf8FoNpMz
6Tp3diujDmI2OBFqPV6qnPqd9ALDbyBCBCVn+qYweUn3/R0hr+KiSr6Z+ZvKL7Mk
XhDLIze16KpUx0KwBiI5CwGJ81lucYwkd5GvMEYwGU0Dw2/rPJIq4qiBNHVtVw6s
Zt7hYsRe4pf2+P6e5J6lDH2CNnA8FfhwCwqSZFOagbl86XqUwVc0ppkixht7bwAa
MhACDOMeJbml8ozjBsI4LdhPczLktdtEtm8RCB50LVdM6NREnZ3YhWPLXHLd4UhG
O8OgdR+AZaTKQyLIa7PVHQ==
`protect END_PROTECTED
