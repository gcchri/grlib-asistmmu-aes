`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8mntKOXv47SYX6wwWa8xpZDH85KN8TrBExKI3yAgUPAWyIWziZdTHcAHEiQX5rg/
pqvgmXmGZf1IMfc/LWBm4sFXgRJOOxXWhDp/9F/b0pWN5UHKODOTmsKNbEXFTMeX
eDF4SXeM/F4SfZPoa/1XiTcvHoUhnbmkIWLusYhVm9nzdgqxRgWm1tvJNzsIn9hR
WESi2mkuCFnasE4a62bkoIzsEWRZUL00fErzuoLoWE30W4ghGWNU7tbiggRxTIQA
wFqsgR6WH6t8HjcWCe2t3CinfQRgZlu0ae+olGnNPw8fpbZo48MC8UPdaNx/PgL8
jWKdl0eUusc0bbkmP7W9ppm0XlEIkbu9Ay2GUtgarJtR4nDJ1CJMzRUnmvmXud6G
80rXZ4heizGkh3svNB5gyw==
`protect END_PROTECTED
