`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+34Rh7e2zbTm0TaPO2rPtHlv58kqAKe0ZYU9gdl2BsgzXvB9kcYrBzaCDevvBE55
w9bU0mwd4EJ8+Fez9KIEs/Aiuk/iiGkk9U4haYTJoA5zUZ48sD0+yPI5Jhp33cK/
nuCPWKwSR0iD9q6xjDNPRr2JI7LV7N+0A3EVs8DxKrvvAbepwYo5KatDCgqabtqP
m2RaD/GxsyI4VloCwL5J3B7I4Egdhcc9BX3lS7gUqeOerfXSmhY6Z1fdP+msPtYD
CqZnTUIAVDplaqjTKggr1ZH+6t6FWySkjOCbKnyTqt0ZK/ZvCJh8Aq3O5QBYnFgw
ormcxLs1i9l9LDWsIawzPg==
`protect END_PROTECTED
