`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qKupTGs1EDEI4/tEo9KEGWb+RxzRpjv5EJEbx5Ps4ReMwA8POIKg5f0joQzHlUOA
NHIvuSNXnK/lDR6Z2AdsTuWAx/pt7LOAw5DElFPPXwyNeBrhux8dwGZQeBk73T+J
Sbb4Y1fZBvdW/bNoAnzlCgzpP7k7RpuEYhvHr3BKw7Lwoqrs9RQKuWMPGG7D8RqI
bnPQ8iDSucNhybnpJl5Buj1DvupPUb9f4o5NhNuo57KfSC58dIXjYgmrPdRjkypi
HiOMFqZgnwUM4N9kkGeNeclihBHb8Y0ROxQLfNrmeIWWIh59isX6yqqs10IcMoAq
HYSj9gcjR+i/YCPkW22iqgqqxaDtqaa9A8ghhrZEbvc+fGbkJG6PL/2PnHqa15Q4
P1h3+4mZsmys01v+O8jJgG98WPUq4Q495S5LZT9uvnOCxolqI92Em8UjMSHRZPS0
apJQOZa8fgHjPk9Ln7KmEUtC7PeV/wsuVE+4LbCwaDjNriMzRGu8PZvgUdCPaACk
`protect END_PROTECTED
