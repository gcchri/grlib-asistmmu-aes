`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sY7hTyAemH+x2ZPb3uDeE0qUQCo/TfZM1VSOHPCslsZ33RAu+VRd5ksDfkK9b0/X
sgNXRugtUZ36bziC3Frm8XDO04h1YlsX+dSWQLx5wHq64jfEYHBpQP3hil+Q4qZJ
VoMU+OM1qyZvh92O8Z17VlqwsqDGtDoS3mSiKtalheH4hTc8CNCyXj32s5y20WEO
VMqky1wKhx0KVFboL/iZmcUhITCd636QgEmPcMA2n6FVNZ/4rF5gea/91pgNGleY
YtOyX5PTQ0RwRSOKWMi5+LSz+TLkU4C3v9Nti7Bj65YtHAFO9SNuNP3ImzFK4cgd
ps4MDnpjPnVEN6/5VgdDIvM2BpcBlzQwGp3O5BKTyGDWJwcA+V32nUaHKe7S13NJ
camFiwWrzZ/38cw9Hg0oRPKBUaoo3+OqDSTWLkkRiJT9K3e20NdiJFMX9eCW79g6
20qwQaoB6vVXB8E3pFvMZhBb811EQmpOS93Sr/KQQANaBF/GcEqxSwd06GWwU8Ud
x1TYc9hDkeF78sOj9itYhxb+tCVHpNh4O3tbCI8Th9nee5zhaqD0/QAKdtECbp5N
VIs5BL1aNIf7XuWC+PlKS5bLyDZgq5fn0ar8sIffDRE8PifMYwEGZiX9A6dmSxtZ
IX38kn8ipPjnIu4xNTDENTlHaC3xJg0s3102iqNlOU+czFbdLXBKGiQ005De48yJ
ZrpySHCGvkQW7kb089nDmk1UpXH6M7y53bhWjFPjVwaIWXgU2SbDEuBaVBcoma8z
Ip/qFXF6hPBwJ+DYqRHiRFpY+6V3iBMmI7A8KvEBUUNlhsczxScSThgdsmQiyjbC
3Ir3eUeqydpn+mK58rNHGa009QwMCT7qSIb4ZQ2sRLd/Q5Il036IB/fMjH8wR7ED
OnA/nYxrRdXeEcnXbP2u29AZa0fS5KLEArYYyUJhEvAAuoWugLeuWWYJyGPA8fHK
Hnpq5ciB5gE+X1wzXPekGuyPRqUxjX4523sLSSYO80b/ioD6jfCufz9tozBuf9Sn
G0Y0xM/zj2b31MVcgQy0KjZxdyllH0cetkfYXGH8iGmivCBL54tkN/vuTRr3cO+9
lpuJ3tO3z0P4XaeMBy2DLn7nIrtHwjojGm+odo1TtEExzbhyzWQEBX5HzJBiju8k
kfsHhJR9bKrs7jZYJGsyIuZ+VWXc4wGpSblYYRWmPDOdw/Zl2KxeXnMWu9MgpxrU
hpCqiYfwkwiTtuSEhIKcDmaYhBCjugIu4YLX9nm6lYuzBvMBCTjH90ZBEVQdft01
mQ/e2YmN+z1dWAr5QQ/F0dwHZNVzI0KPHktHWr/SALko94zgWxBpuRE0rATzdivr
lo3jQJBqezhuplbSECwHhkPgOsjjWajdwuULY6N+TFq/clsNHQopESKgqdQUmwCU
hKVAQEamfZBckUvHPsMUNUIg27vnGrGj+ZlhRFPLmzVE9p87GwaGQCfh9Ll0pxKn
AGFrcACUWX4zYMFgLXJUA+2yNnenkWD3WzcRSYqQgs8Ct/NKlCGlUAvzCo4lwTJn
DbEscoWbgi3xjDp2ZVAHBrp0boHt4PYA4nnAdta9AJoE165zAolNK+wZxKUjUXZs
DuBT8r/pV1KF9c9jsXSGXTXbE4sd5TKay2ITQKrW1S8040edlEhvsKrhcTSk8o2X
VIOAqkISpGbdLZPY4t+s//QPgXSoEN31XlVi/NNkicF1VVk/NU3OAYa2ZGgLf9qL
`protect END_PROTECTED
