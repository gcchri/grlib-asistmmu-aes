`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G15Z8ULPulyJDdZoh71Io+Whg+bmyk1UERToPguUwnWOt9GVuLkWoQOyowsDgNat
W5SlTH+HCRGjxJ9YMzsdOPh+jILSQkOEej4ajj0JebAVrewZiPPLJqak4hdnBPpd
WmI6t1Slz64G3m8akPCG32mejPIP7OiktbmYL1alurpJkXuaIo1yLXSxkaAEM7sq
tJsKCr3qoFYfLYQqtnDaN7JK5cGcypZ0g4hWLjeiLPLmq8rABSN6/3c+VFM6C9a4
2iziyG19mDNsQifbtvIwjPrKzMD5rIMHMB/4K0Wk4RL0J1qSsynDT2m8r2WjneDL
tX2+jmAu2vOqR7FrlIiwYFcyHW2Ch7wa+F18mThKGzDmWFS2Rhr8t3I/zWPQYwa5
`protect END_PROTECTED
