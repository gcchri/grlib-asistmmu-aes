`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UZoFXn8J56Q3aQIxGpRoFM057LcgNU7pD7s8eqbfSpFzXjkiZ5V810/i2DotI8sh
Pu7vf/39c2NB2Xoq9xGZtyn7sIoZ8yp9FA4HdKzlnl06+Ms9gE4g+dE94XfMyJxh
mBzPQL+YJnylgWCLpptypSpFGxtFcCd/h6ophvQGYV8piPSLIV5BmPrN9voxmRKS
leoPcamZgzY78i60Vi1WAveoPUUWrNzgmvrmd2ueCdxvFjgDYZPcOsGgprJQos8M
PUXxRv2IL6jJJmQ/RXQXsNCerU3c1WVeD90BJwKZAWxlkq7BlZFHsGKor0Y0+aKH
fYICU0V1C5fPbbARsp3IkrURbap4bWxsGMm6EHjf4gWXj9PabuU+SN4EtqMQVowv
FZFQp+asPKY/SErhe/w99E9NCuoxxvw1vLe3b9MPLdgA7Lqw7P5VxNGjI0cArUdf
`protect END_PROTECTED
