`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iw+5VCv/UbfDTPminBdZbQyoA/w4lhsh/tW66XaGlrvl5/jBTCWrzkRImUYlMXo1
thsIazdBOsIUtrVolawu0zj3VDOpbRQR7cj1hP2Lj1XEDHw8n6/OzhilbV6eBkVk
hyCaTeDoSBvp4whD5ORRPKKgdO1rDdhAyq1xnhYARIUD4GurHyYMGv/9vje3gfC4
jrc83c2/bywnjbbkk/fLEShdyOQDVyomTvL+Xag9ejizQNbLIN0m83ZL+TcTbWHr
e2DoQHXGCmdIlYRFXmHWEdekxIvbVNQOeeZW236qNaJcCsXwtCgPoLWFPES3e8Ro
R9TnVcQyg/77u81Io2sfJnBDRq1+ZmHTEETbF1cu03iXvLEkBDhmMVujK/1OcfjM
P5yr2tbM0dGvbX2drs0ixUz+foD1Np73CcT46MmFn/86nBxl6VuEGhy5N1c9RWGR
Vhm/S83HjjKmtIpr+7l0R1f/D4ApWxtSHuPmeiRBxGR9k2h+xqxwbNK90w3Vsywx
ECeGmQQNaYM2DjJ5+x2Cr/UGRV6Z0nFbbMN3F2VGad/Kwf9at/w7j6V3nK9y24g5
SqUdDN10n8wg/GbAtW9lJRDyp/gfXTfaE8RvrdO4zbNLHpI4szZX6KtSJqsqQc0a
SJb0dVKJQ8GxFzSvld4z9PkhGsUYR7iHOgNYXQHEgE4=
`protect END_PROTECTED
