`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
obUI+PhzlwiYjVzfuRmsuS/msskbFBwxOedGgQzPmxqM2SZAgUlgwVJIC3ckPVn6
EwNKUHdqImxmSpCC9xU3MgI1OVpgh0BsWuamX8+4Y++iKZKIalsQipRNe6CDPjN2
yDIj9238Dt9Jp1G3JElSsGJeeu6nHGlbdqKYiHcK9m+5HbwZR+mLUglK54gxwV3Q
DJjE4J4IiT1nVEjjYRonHhaWnwVrK46qfu1Bh8Dk6dHUepNwDAvqTjlTZiqxorFh
LXT0ZbkTEMD96qJ0RsEZwSDsyMJjgYvEklvah3DTPcgP5UtJ8g3Qxt+L9XYImCbC
plJbw96BFb6bhYRtf5K53BjRX4wxjy+9kZ5i4djw9wlWYURemNSnf1iypoO1Rn6H
mKidTtm4wJKMDBN/tZFQYqENeIzmwdIwwwwKuh65yzuPePGv0YdLNNGV8SERjLfb
1eW4YMR4cYfmlRsMPyOCsSJC4hz/Xad792wuGBhSHUJbdRbJufHmcOurdblPdqRE
FV+dYv9EGi/hSZuteHt0upIfttcz3VCOg4BEznPgH6EAXIIDkrkwPSrDYGRLeVAI
`protect END_PROTECTED
