`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O2LMKp4xZq/An0mA+RHVYJf8OYlJFfVB6xd3tvJAj3juEZ4stIZZzhfRJccJSW1y
VmOrBGSpnNKb4zL+KVze+psFsTY3WOf5SAg6ibE2z8AUvenE7F5YQDNZHJx7veLh
ggiYV0eanvF35Fv4sy2tvMFd8rS7XsIsAse0DRRJ7Tdg2msibOncxli/f5VU5vwH
MQxEI8A49cE7JOmk6F8aeV4Bk2a0BIKHLihLwP4M82lC6LLmSorNlxYggqF9+VGc
tdr2jb8GNcMmwTiIG7Hlf3QT9iSC0QhA6DOtJMBIl7ipLQ2X9c9rsEir+2G9bQL/
ERLh+k2oK1qLlwlW0+HDHn79ZIrEI5GXm1N0j+LQMi0+NlObwj0KjCqKxDQ3C04J
vIhLtjmS18y7gcbC3ISuvsh03iRf7tjVWD+IqYrI1pGQlDbwg4Fk2t8nIo3XDXdk
Q152MUXRP+gCg1HMO8MYOsTo7dERSvMOd3ms1MKCriYf4X6ZPzTm2RGEq6WhXU8H
bi2NbXHDz9WMdO4R9XA5os0+mQgHMNpO2YHSU3l4FLXN3W934w5DGeFxyEz3rGO5
NWnrY2arwTHECzPYgMnewCuC7oUp/Hj8IVuSMs7eKO5TElu5TEHAI0M8ZJL5ohkP
iZx6tls5LKGAiO8oT51Nmnm7+kZwCfU/nCLKpuko4zOgtOSFgZlGp/PZ3IEmoWg0
`protect END_PROTECTED
