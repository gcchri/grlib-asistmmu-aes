`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ackU1ClPsmDDmegctq/XQj2X0RAikMdCNNbiSqgOiA3W74u9+LI+KgxHS/uuH1d4
x/ws7xGpoBZkOdDjNlWZ9PqSJNbMULv6zrqYXE7Dv7ad/uF4Fib/NA69jWNndN1n
bOzO4pW0VFfa/e1kSz3t7u5f5xr2qUO9km1VqFXBpMMgqCNNGk9ht9M/shg/t5I3
lQpIniqt9ExSF96qkiTmlmqIaMSqCnn8njb0GlFzWdpY5LJLamk6PLXBRmU1WE2+
2nfCQJbOakANdTUWZKXO/f7qpA05RxH2CK64KoUOZlLPFShIsfq+I0RJOsr7fHYZ
8QUO3j5rmnAV14ZXKkJrWmCjVLc86bxXWqFpwCjX6COjhz6iobv6caM3es3Bb6y6
8pOPSVA+b+26vJZ7e8POLIsMXSmcftjFhN5aEisV9Stb3sPPo4Y373LHxqob69tn
Og99+6dqGvZjHlXvyAvoSm/EA/F6R228EL+LwOj6mXMAF/K65AszkEBXqfvMKNd9
TIcUCa6TMV4yx90Ovz+nSEPIQQxR1wqQObM/cjL9cfDdFv2Ov7RjVBN60InHp+u3
noISUmxG9HOOGTJIWDv5cmVGw4wqWmqKu04yUr8M+pjVHdugqUisqR/tWTPeuf1/
+DLAcATWYPLccxh1asl2xp8EQOOat6+fRCmljEP4i2rrjAdpmkH/55XM2u0I/6xA
XIErJqjxqH5oPT8or1XHJoO2kAV+C9/H/3pj9Wjp0vyfGnCcE7bIcukpo/Lvx1wF
qJA9q5Z9pvNwW7GK+aUBGQvTLZwcUZSHHwjhHgtMqKKlp5mKEAvH0ncwRbg471m4
4aIcCznkGABjp4pLMmldv+zbyt5CLWSRULjHetHVzUoNFUt3+Sc+Gtk4httR5P6h
ZOy6eklRkOaSjG83Txt8yiWwmT3x3wrqmqlMGGOarQ38a7yHBg/sRG0/mS0vmg+X
v9Xk0ICt4TcsqBLKPGOtNGc0vo4225h9DS5IoAPb2m5ygn94PNhXF+7UjfRegpHu
TfZ7YBYdrJJXYrrxyv3/WgR7zDwJsgcQObg/b70XOs0M6NTJ5tk8dRh8UYHziXju
poCWyhhntUVHj/+ZcuevEj1syghkMv/ELUOw7vxn47ILs3xaBvgpYFpht5SeYUXz
RazQspAdOrX9ZcRul+HcMA==
`protect END_PROTECTED
