`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9KyvkUpiKzzP9R/zrzb6Zpof8yVpzZhvI3HO2xIgNxS/RwcHaH/2caH038lVzbX8
CHxZeYb3yu1Pg4JNqppCYuak2D7UNTpHYXNLTCkut+WJNtAgpPeDn1nvkjedFLbo
T0N8dySBRvCCbiAsROCCwdIZKLFLvDZkRhx5HjSuEilToSP6ciIAcI0Du9jkHZ7i
dztYUm93LrUkV6ARlFqeZOuMLbyUavW5h10iEpgwQR5sbXSldsx5IeEREX7czBLe
ZWtdHPIV2+I3ZjAWfK9M1t1DmGz1KnrensLJKb8a6VsTpAjf56pLfm6IT3HLQDhy
tE/GbQxtrN6hKQoU6RFe26GZm9e5m3X99EWB5O95FzmkdzOKGQ1p8bTk7P43ndkw
plndO1XpLFz1YWWPCZTJonxukIzzVC0xEDFlJL1N9nI=
`protect END_PROTECTED
