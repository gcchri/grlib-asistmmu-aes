`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
svW+mw0W7u7b9avUq9dvIwVLj9KZQjbsbiqlkJOeeOfPL40OfbJvDjbjBd8muQgY
55bQY8ODHXh69wuC7QBAP+9Gxgvf30/6FbTOjbBr1L5MxtXvczIq7jRM6TmGeqDm
axz2XaaFPJJa03YRw923qd4Zq9BGsj/tcTCd9lM2XSu6LtYi53nKAO8M4FxdYIQx
t05K2+R2VcfCEVb17l/3LEof1Wqe/IIG61OO/d8LbOEXWZcedRcRw+DY/NkmogGQ
6oQcTMk8YzJQJeYAiu4kgxxYPAXU65wfobJor/+6zpMGLQEzShl8x3p78217HdvK
mlXlg2tOIKzrghe8rcFNC0rIn/MGptaFBharT1opYeKm9DNjN8bDQrHhwy6nnRU6
0pruy+RHpcn2yA4CWoCEnOBBDXfZsmDxpt+a+cYxzsU=
`protect END_PROTECTED
