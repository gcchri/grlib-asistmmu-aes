`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tWwiCF/Mo9YFd8x5E8IYAZdciZTqSFUFym4w2PWq5Pb5ArK7ofZb4P3LJstqFghz
Fu466WrlnkJWqyGuQgxY2ed+uYBXuuoNvKp8VLZR+/6orbjwLJgLt5iW4NNwC0i1
TI8NA75WcdJyhlkQ9liRooQV5vwO0SHrM/UvJ/YjNn7kQfvPExkkU21pEz+1g5FB
QfDoTWblGPyeU9QMNT0AMEWT+caqOC9ng8tMAuXg9LTDoJ3SkgTtUE7aRZPHyWzZ
uhrpxYppFb3HZkrq2MJs2Zs8zmHhRlKgjpNy5mWJICk/bqXxlQWgxI3cP4wIQ5Aa
TDFjbktk3XN3DkH2sMyoO1ZKHHBweYNnK/Y9/yLCJrQjonn8SindTQSplR4roJhp
jfC1wPc3IDOYkDOri5m34cV+8jqcL0LMqTOALvYIlRbXwcMFcWGCe/y8mBcMWTZr
K3/bCqW7Z4eq+AXyivPRkQalT1cBpzMJ78gN+1lduWPEHEsUzExLIAx3bDldu7jJ
HLqUqZKZcFieEIF4v/MP4w==
`protect END_PROTECTED
