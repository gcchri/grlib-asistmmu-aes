`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x/xZ7Cesd1g8z9uyyAQZtC+vUO9Ni6UR9fG92rcHZ4BCAJo4zttOzNfLPYDifeHn
WKIbOYInDMo6IT708af9fgyUtQ1yie7hXSOoi0ic6xjTZtjH1tgU0UBel/DegTrS
F/CDr2NPE6kTUUTBt2S8PZalGmWyx26xkWURUOiVKr8m2HTTb7eyaT4ppIQd3Fzn
vtfo0XL8WxnEqQkE5uCLYqEX0e1ZEZktvuoSZiWhuRrlgfrlKdw/1c/UBxl6FS4m
IWN6RyIjE54xZ4XJceHG7nfFkkbrH5oGU71CbCA+1a7fwzkZOQtP9jSndZKJz66j
WsFJsrmE9nSyJsU7dGueH5jZaTkP4g2Z5Ho7Czv5EVn7Lan97fPAdGROpJx6cEsF
oqhH01cq/a+yrIk/Brrai/N6aaQ7q0TQWOK5u1qwVKJo9gNh4BJIHAuUZcWKFEEK
yjBE6o7QnYh6g2wqt2Y7yd84IBFIZGvg6hjuKBLb73s8iWpn4gzYJd+8sBT3u+kD
wrQQirWmMoLwqith+LNW6CWUGCMFhh6eqHA0lArBr2pw67Ht0Do9x940+HgZIJH8
9PA/vJBMq9Uz7vbs5mA0e4e/lhNinD7meCTNKCWLXUq9/eXFsBEHMWG3l3WtyElU
ReLGeuiGZOwUhbkKFQ2wa9UTVYu5achjS3xHcurFfNv+q6ilgmFk5F7CIfYAviH4
HWapFVWlXGlBZtnXgytf3rSXmYXIVpIr8Mwaq2X9DYp98Jf8M+TUrOa/7sYwcwqG
ajM3P3G3PZhppsm5Rwr2HBL+VI160Q0tUGsMJVNcUIZJPPU+oehSvClP/JQV39Zw
h6Hs79CG4LsWUQ8EJYLVQh+1sCDE+ZmNQ8cwpKj/UN2VXZtJ7vXhFy90gLOT5Z42
niUjAb11fD6RAsQQQAu+l+/irElEbTpylzYx/H/5AeDPCfNAi8WrASwTckw3fjj4
nF/9I+KxLuu09wsgnpnN3C/SJAj6c3uQmLIMX1FwYqTqK2tqa4rEAgWfQf3qnrCE
7OhnvL6ywe9dJBZB9sO1W+QOd5mYGN5CQ+CEqXgFSpUrlZrVcyu8v62g05RLBcSn
zC9qDZS9AFHrP+Rr2WMEByzqzqyjwsWWY+RI44s65aa1L9pvQGjgzYwT5kQPKlMt
fgnB0VrotIQBn+RI1QCnnnOQzFbpN30p3+mu7JtzC/J3h6wu0vFgb36QOY3LjpUg
MDJ0mIpqIgMT0pe7MwqdZ2OB1Uxi8K/QZCMGAcHQ1/Fmme2fHih2PF0UXF95A/ZJ
kVc3CsJr12fzvH2n+YMGwi6PI4zvNG0tPneOIfYFOGxXCPfA/2BBeU7Z3WiVivtK
dmYmTi/ynPdikt4O4C0uxPDlZPm6AYBo9re6h73xXKgJ/RxeRyYljxclalygWfut
7vzdqfjEikK7Gt2kzG036Q7HLh03/vtbLQqU/FBypGt9s42ueNQ7GW3EpYwPE0HC
7QQjIRvaPOVquMdIeJ7k9DcP7FJiH2/Exc3pol0Cdg/K5LjDhGWxky//kbG0hEw2
0RknNofGfAQG4emux19Y5JHVaHK8wJ4rXbXj7Ic9FNYCebbBPd7NKwabf5tRjsa+
MMocicRBoPxa4HNAq16/bJJ8aRwKr/3o/SyVW9aaQw9R19qiEUQMuxuZaVjFwxSq
lK2PhQ6Z1/YnBL60UD1IvYo5sDUNBUVrCPueqzRGn4TQmnNsFXLoY3Ea3ABtBSLZ
issmXF7liBxOD0Nsr/3IaM+Umser92BlGdVr+GqKdTHyMOrdwzWUTpaUl6eAbrhl
TaDMGgz/hAP2dCA+3Rpp1NCgNf2L5EBM2gHSj3e7w4EnBBOxrvxj3kj0iCgV+TXh
yl5SV9+n9RssLHPX8HRRPSLenrHYJMczdeo6EUGZqPhRkYYx9+J3zDN82w7cbnm5
wVrKstNiXQ8cJ8g2eOmVm2s0T0px1UqBKWXdSwbKCwOc0vPGtlQkn2uFNESWC4rU
FIiQ5yyOgIxPwDbKo1Ftoy/U4RVELB42lKlm5xccIR18eB67NG5LKGEUH+PeS55E
JOYWEBkR7sqr6UNAe/bbRhiVsyq9hPKT9a3HzvrhiEytjEBChsxu6Mua6vanLTqq
OLWKT++dRuEHemDmdyjtXcnXjGbz5P0JAMzeb+rnBVzsEzIgpxautjrd3EXCv6IX
7Q4hW1OHyMdCV8+mfYzq+haWWGd7QgWqO9Bqxw8Y/glEfpvlvZIqGXIRVCKL+NOe
SCukjCY69vbT4/L3+uPA0t58E3rBR8S0iqeZ1BQl6Des2QdgGDux9wvEWK3zxIWI
RI1TYBdQpJHRJQaCdudNurjmYYP9HpsVCFj6/IeHLUQnuLOwQE40GVIrYchJowpH
mKuX37hm1kkUVrrUWVnje0uCUcmLvT3vmSurVRSLw03rmrS8iuaebvitA1IGqc+q
W9nquetoOykA1owR43VbJHupXHpCWtcMwCaYmQPytIOtQLA5cBBEvM0+gIw73SuM
cYV89C/JtjIXVfGwOuvmdgHo6jdKhPkugO7W3GA0ZiR+VuPsWxw4MXk+ROnr0kGR
YQNI68KXFd2opRSNwAhaUNfGGklgpcE2yKksjMcF78ReTqr/svlLLUQr+CJrtPCU
XiJL/j/EQqwL7cKZtry9MFYsvJ1yfwVziOT/2gZ0nV3wXz7iO56lWZZamjbG5vVM
hTg2vlsEt9u9RC4vpMZj2NLR3eb6pb5imxN7GZJXijHOw3uwpTsxq+BgUHa4TYxn
hgsMvtUxQy9wGcJ6UyoOlYSbRBmT+yL2ZEeeU+672fbLVFZL0MpHlCSIG9RNnaON
sKf+Ba/byeVMgDvLH/Bg0Z9lPxn5KJs83Ph4n8L2omWxcHWFZQq7P0rqQ4hV1tAE
VYyo+Sks6kfgMlhkyCJNOkEFWiJpmj8ypcfUUgrPzqb4Xr5hOCcRa/cZtEwrju/I
jFYLRARP5uKnCTKEnGRnMUrZSP+17eMRJ6ipoOANZXLI4G2yFzHv9E0QGtSX9DDd
Te2aHjLePfTaprAo2GEVASGWT0ptkSmmmyYiMAQnVEONP+OrjvZvQFt533pSPb0i
3JZgfORy232WsK6bdA0PLuzKVROqXWu/Wr8Zmgq16kRLoC90WjmnljoK9i85d5qe
KMbBTv/JdrO7TvcarOD9tlE14gR8U6wVj2EQMbe7Wmr3GIY6+XdUec/F/wb+AoOp
CL5poDattZjKtSSRYB0bxD8iffQWMclhEBxsOOdkr3LZanyclpezK5gPo/bhX6sG
ATNqDL6qytSwoDwt+zJLAj/oGrvZhLH5/FIIxLzXMp3saHnYbzWzncGFQhcUtqvY
S5cALgC4h4L7wvFmyvEXt49JMEVKo0y1KCovylW+ghWFCNoHjXC2XKDysmvZ4U6m
sZK0+GL1NljjYUN4EU4RR5P4g7SBpFStoU0rlWYkz7BO9wj0YugwSn95EljaSp/R
xahOAk5tpQuk4l7ZoXhe4loXPjSwY2XZvob/FsNZPproHu19T8sTLsFvWBK1nF3u
ikZEDBbiNVWzjrOEMFZxXf9crVlCicmkUnDoNhb6wlsSQJcxTU936lhVdlnxFlQ4
cd3efrm3/xAjJVLPjhaf7d6FskXaYmxrc11EJvwDsLgGEou+bNEwELi8+Kc9JGit
FThoWFnu1+vF8ssctXsueAEQj89rzEt34sMo3c9Myp/SIxi5MYHBumdqdjgP7rb/
RjKsEP3kPdi5Ur9mcfxQodsdxWqd5jp1DeoVewB8CuhZx0CBhZOpova4nGaTw51W
LTYZflx606FjofC0vCnq1REoF2OWGvkb7gxOVVM6Ol1SuQKETv6cZWJapaKecjt8
XhYpaKxfvgo0dktEADDxAJSlUokV8tauGtcXhUiKXe25EMwiZPrNMWuzW7CCARzw
NkbUT2sc2eqwSPca0/MWJk78rbAdnTmjBRIqyytTrIb6K0FfCLQHvUOsYIAp+BBg
0vqVCAnNmHeOVDkOfv1xqWp2Aq5UuQkCeOOgo1R32w5SRhDXh5MZVYSyt/Fvz8zJ
UI/Q7Ey5f9wEYEZOIFm7bT8X0R0XaF1BA7M5vP8GBjmzbPO0dK95D9nOFXt3ECFn
/CZKgvUlzxAKVlPwkqQFBeCV+WgVvJeMgqnv2iO2CSvVhNnZtlKchaDffCOqmxpq
/IRlmpkeTbpszmavTf8xU7MfA/PFYEqidKaxKn90Jyq5/Bru4rlP7FyKoHFUnyic
7iV3vbDvh1/8Rr01KxZLrKssZJtfjKx7JTT2i6F+XuUZntOessVzgp14hz+HnS7y
ojAaOIDszlprS1Kb1Lf9DEAPrlNUuimX8ioheSaTWLhJJqxSWycrmeHB1pwGMCrA
xc5QLP6MflImEYVHZRTkrK+PEBazhTrmY2AWeQXvCMPN8ms5Mu+kQjMikIE/76VF
mhsqv0Zntn4/jPddvak6SY0bVWc+N+AwztJ6LXX52bzoKkNXSI8Y4OCMSq5cGbcT
Mzy3ZZSLHbGY2U5aFSE5MIfDGnRRqS8F1mVDWiQs1Er9FJgnsxx7CgCWWbfaSX69
dHTKjT2l/OU50rDk8G62ayP5Qc6QXcd5No5j74aC/Lod5FFd4gT1AnUPWh6fF3uZ
8I1SQbGqgMes9CV8cDIHbOH0kXqlBOzo3IoXFXNFGORTm2ccq86iflWtvzPS38Qv
3P9s3g0WxjXev5CikI3e+357qVR4Wo47NHhsCzsXXASM67vzL6t1sl0tQOCt6Ee/
7KwPTsu8DNxGRy8QY2/B8TeLKQYBmXVTsqQLdz5w3HLcxV7IyOGncYx3koqrSIUy
ZZaQO+XSMpIMrW0ThHt4zUgpsjS/AF2OSwjzhogT7Q+bpE2NtBsnAenKFWv/IekL
uimRXTc9i32OSxr62iaP8vTcL2SrhYtc6yrxBTtOceG9W5RJ533c9idDZjIv/28u
qDAtUTL5WBvWSWNa/6SJfAbd7k2b/Qb4XJc6ucJSjtxt3+w7FJQLfhvJ1Ni8gUfd
vsLzCtgaipJsi2l0UMTWOhoNwupNoUDHSCZtcnuri+RR9mG9jpnpfxZWmUFEbmEv
pv62q6CHkFA175Q9gV5s8q4ALApeHSt2T2ESdGc3sniZQwNtydmmLLwKLL2gWH9j
/WGfbRrpWeheic4RX2E5ht+BkzNkh8H8+nnhE1Adx+MVGaAI1bGWojIcm/kTMHLh
3ut8mgkBs2g3MrdUQ48o1Mg/ObVHMp6v/ZAmcCLCqAdNdbnPxmVoQgV8mfBCwAMG
AQrMxvDj+2KTomN2pTMa1YNxaJ7F6DmLdrMXp0NANHL74hVVNNtrjOw4vEM/SaHw
LkQ31a1GzT0iemlowSYj3shGYvBC3OIGA5NGmb3k5lbI9NAXsemllUQjzhMvxrPi
+KlMKnZit0MkCssMFeGCLwqTJHZMglU0DHWctGe/+ljyvfvKHVrITSdDOlLtSfhm
Q1mtD0+yiHjASdTLUbmU1kVKFX/9KDjxIOc7I28aZTmTL5+XUWUwBUeYVVlAxaHg
NSLyiKbq4mW/T9TwXL+DdZAfgHEaf8UKdI8LG7mhV2maoXKeP6v7iwp6kRg8VEAn
ySjI6nSLJilkE12bdSYQKN4FIP3OC9xp9Y46YrVNPnVT9WoIILmJ89j6Qf7alHHF
IbtO0qd4+SXFJkbiX57MH9Q48LpVdre1PB3wiTjtSaHh+5wvUD20vbGqNh9J2MdD
ZUuYs94GEuXnBDH6bpTejpNu3jXtxWLQ4m1GV/EJAh1DdYWz86nHP/PzAMYDU2A+
f9ZG6o/LoUyAyw6P3Ymo+y036ROImzcEkbQobJu2HBuvimU9eIfN7rEOIwvYImOf
cXTrUAtA7SlXLWD3lCCq69emsTrp8ll1ZfnpbM7eDHgsr8fronA3e5oSRgG2vmzR
MT3FK+qURb1J5aVzMjSur2eqUF/ioDNfXkSvLKWRvhqLw+TRgVt8ad88SmBpsS1l
oDF5hrt3rVESlCVsFd7v3C4njYAg2xV9l3Je4U5cz5zyv+hw3NXiSno/HbeE6kUZ
SjsJTa3f8XluHk+5urOnnmWwWj+uemslVQOLdrhM1ebl6EyrEg4xt5tjh3pHycGN
OWLNX+V2HtpMizLgoQPPAvDnY5UsaQfCR9/HDnNDuu4g4dUESyparIGMb3cuuEQi
k2oqy4Fg2mLXAUfSiejbi4s/LF4v4/zxdpgd0PY7jibsuTtIpyexJ1H3//NyGU2u
xrLg56Fj0bBmqG0ubFAbqT4hNtPmsxo3aT+pzEwom6L4SCbiOXlyXoK642XlcKm3
uzoRzi2QaJNs3UgIdlkutiFv3z6VPqWWVe79MFbJuCosghLdJpiojbC48wkfRhIv
3irH4+zx03TO645SU+p0pW8aviVm0byoeAHMrByj0aMOsvStbMWS6qlzP/IKAlxY
UB4CKDGmjJd+RCy2e0ixP2XIl1BMrTqWNL2yesmSOe1ORB6sYo3Z0796husTB3LN
EWCfQmr9CmLvr/a7ZwbUCQvpxSq99HayUOGvUN/3xK9C/bjPXPT5qRMPhdg/PRIS
05vsTEitCNqXoesADh5Yvu7XFm6Y2OUJdPAkS4aZ+2evrnT4n/tyT7f3cRqJqJP7
0fSNWVDz4B7GtCxZKVO7vDl4sfdxLeHznWzDwBfjqCmOML88+1r0JsHRX2yjRlW5
9mPIGA60/XOKBGaDA30Xf25U54OcYVJPvCMLpp3lW3gx7yE6ab9BNkU1B0tL8aad
rTVcjOXZOhcNrPmc/FrGbOcnZlnzSvin6+ftZSD0ZfI9k5GNdsi00twdCKnvR9T+
6ulDcd5vs1rk7Q9R6RJjOSlP3GEywr98Pnpj2xOpsobOPmByK/xd7f0i816lhzCK
+PJP8lsnWW6AGNsauZ5y3Vk1eF7Egt5ip5KxXl39x6iq3tJ9054w8+FJuHi/QLJb
L9SMlAUOUeNoJRl9Bbj5p+CIu/qIxY+fKwbi7tb7MSa7v6ro8jTiUi7owbq0ev2h
qQc2WCSjMO2OS15XY9yc/xiah46KTnDjS0IvX/GJ9VPK5qN4d82HB0w6Pf2AT6kh
jUvLKwvkJPZ6St2Hzdp0y6ZMkRJhMcs9PLrV+GyCEHuYTOJcRpHvcufsoYfBWGv/
mWg2j77w0zDptXXT0dZsA5Ik/iXaOmd7P8nk8/7idy9MPi5c/AXwaYoPYl1vBeBz
bV/7tSxAONN3dwAG7jKIxYqG8yRTuV+dWk39UUr9ejDARrWcnViwIdSnBwVJCWe/
EBqFrcP31XisTluwLytgvbmnjPGJdaCmq14mb3SAyX2QpuQN1UwKxunWBqZPYGYE
PXEjhOmSYbhc4ViXJ19J2i1WOScbEZQWCOFKF0ltxieSCfGEW9zMHCqVhSJd8WLI
VKvO0XZSPsHABPpwrvKrXHobp9oCpWghIuoGd8mRjAbcW48witvzY6qFd56EBKEV
Ixm/9K16tFvCTRqoc1O0KO11SgNLuQX4JNEz47g+dOc53KXF8z2JwoSa9SDkQmnK
Rdh0kuyd377d/KX56ReLM+GH8eSlQSzXmIbgzgpYgEAK8/Q/UeqLWaSVfms1YJDK
oqT6+3JYjycDOUulwvCmOxYyCMgmeQL1v7CpROAqSqLTbWE8gxFgRWYnZK7c8rZa
0T3jlYnDvcy/qgOwSpedfvg6kg6wSRNxIJveV8SlaIHKweSbfGrPkVhaU/gjMPek
IcJ4ottzq5dOluOySoRx03DhQJvKH7GbyhzMy8nYM8mtWZkeClmPO2su2QC2NP5K
H/MlbNUuq44cYR0hVhhgzekW+8VpUsQoJ8ea6hYQEIaRDHL0xmgv08b9uvtHMvh5
qrCSnXd7n4GqhwhATZdRG2W0cvNbDAXtDU1w7cO9Wfy7zlEv18WhBNmLfHGa1okZ
2siytQOPoGLV3AH6bHKcYwyV1MdsHDe2pjGFS5MJuS5Np67Iuaa89u/SqgLq2UDv
ZKjYeKJDliGmt9/pTF0Y2KvmGVbcw38mzGi61st+tzYUONvyoWkMOtG/sjz/KnAL
RvdzmyzhsD25e4v2GVZczfhWvW4B54JmEj7qzJYn3FfclWaoX7+38dE9Aai59X7Z
QQ6ja7NY4R1XMJPXcO6MPhzDbMrBrmoi+BL0ZapmEZ1TbULeh4J/vz8B5CCmtABI
RtFu7CmdFNU7FBalrzodZqdRt4ocd9AlvvuvW8tGl+WwHrNsfm/ySsESa9zsyJ1w
NvJIWK9Cx2C0kkmmG7REx9KVfbXsBJAf7OQtiYlA6x4r5C4wMB9yyfTjhvN+bvcI
aq/m92UeFhmo/KCeXRZfOqc0NXfRYwjeXno45day/wXYUcSSZH//uLmLHkWb8ku1
h1ZMTD8IJgL6saRQJkDaNYj+38Btfrg8SdFLRwDrAYcdgF/HvXxntfgZr9pA284o
p5mReIKY2c2jhLxcZyWykJ/5R2DIPDfy3KFXqKFYmZw6Z0t76TwXvuJzIesCX5+Y
NHJkZP624yNYtwSjPxwqwPGcjxrAtdRfiUhH/aauEtbfOnuBo20VJ5SMvjLLO6bc
7+nFPnnpIQFjww3vfCaAdswyFDpqs7EtzvH0BWZrKCzsPflLerVXCOJaDCUFpfyS
vMTwg08wHkOw2VWLKzlfsLJ9u/O3VyWU71Z4e9QKmnRspSviT2iKWMihfySBMJiL
71mSnFeOSQn7RZWeeHyo4aa/FqxauQ0Uq6n4L+MEPRidm3TJ+Ve8ERKd77AGHp1A
z4bNV7t/47s9s9tmV52dikCJkQ506csuod16oE3hhZPoNhjkqZY+vSsHRsMGxVCk
SJVFqsrZHZiYE7VNI0G/wyLTgerIjYM1LdTqwXlVBvBfBQ+Cb8PoDsX2WR+mniyO
t/Us26rVYR3R7YfigLwtPrr1viV79/XzUmRPcfWAHQWHowBJm8AaIpKNqYmpOFZ9
3jAwZ0cA+/obo2ICFElrDqbKEMvtVGqrOvfvc/Z9pd0LCNmlO6bSI/p6T23mpfFo
IG/R6TZwXdmqmq7BTGvGjtF+ma4xdmmyom4M7GQZXVAFuD9AZhqKH8xT2Vl1dMD4
aXzuidh4icinjQzF1Gm7i5oXSquScNyIdQ3JAh8Md39ZTJ0uo4zQo+hI4i3RpUvi
KZn5fmTi6zyPuaXFgsoEeeiKnlfT4mzYtbZm7DYIx+n4pYrl3FpmeGfbE9uw8djN
XArPcv9aMHll54zDyUZh/VPmZaNDROexOP9/8CkMUN31xGN2HiO/k4xsfDcS1D6m
z0hdXWDIBXziP/9vYpbxIHxjkuOy56A5qx2tfHEw8JCTLlO5YaacojQ01U8s/Lvs
S0p+Gwo6QruBpTHUlZbw73AkAxZktnD8Xu/TWRhWLZ7Llm7RaM4aU0SDIS/vi337
cbMLcSD6HXmRYDQ89S8Uzg6asL6buuCkwbAiC8Bsj6EKTPBWIxmbKIKE0kAEqqXw
DJwHmLiOfLeRjXXumv5tIO74Bw1V52J/IaWMIOfUcApxqnVbxSn2mmsCNqQKbMfg
iqwc6gVxytyneoZjb9RxIITa+W/eMGZ2km9r/Rd8chqPPrskLBMhdJIVQ7wGJZTJ
1zgjqoV9JENm4sdc0bO6XzWCGbEF+rV6btwijYxiDLZ80OAhy6TAtXd602W/czF4
DbJfdngmauQGoGLQWAGaA3EcxalSkgjba69+tzDgZpXvbaiS2qRQLjT6ZdQyWPD0
0Z4zCqSoIICaVz40f/p2EOQAU7/dKjprp732XyUsxyj3MqN9LNbMoSdvcCuOtO0S
jmflgaByal5HcvRs2KWgu9IQvYnY3980SBDsz9s0HCqwAa5asdUS1aS9YG/EG1wT
xysGbSMjvXxNxBuH8Gn976NUUD6cqMIMXNyt0JVBDt4RunLuWBZD98+KUjTbUJ9B
EK9h4wxseoA5urBzh9fp0D6F1LaCfHxdTewjm8lhsE5gTF2f2J8pYESJzOBaIfIB
80c+D19b+DFcG37yqaAsOg2QTmTQeuHTtN7kIey69yFpYMINBc4XBSVAHLgckhjk
sqt/zrsVrFmz3GdzMS7YdpUHLYGQEA1F/gn0UPas5DNvclX+8vkx6l3hnrgAu+jo
pqwKof2TZOl8vSxJvS1h/qS3fP2bWIYgF3+g5EBIfdoRDo+CzagIyJFwPTqsqz5d
OPTUoboyDyJgzjYBetxpYUfFlUfRtjPY0q2jWA1pZ+7/bXpdcS6D1Ag6++Zw38Ss
OzAfRZG61EEuUp+aOgQGw7miQ4BJLAHOpmy12rkoNoII5IIGWjjawvz4K3hRSJt6
nQn7KOD6DHViFQM/H3TYJKR7akh9Os4eLz0OXzqFH8nbWxLfbRDPTIIi1WpoTHTx
47vQwjg0DhEQNv0IkVJ84KBWdqMGS/OtCEFy4M1g2SkgkJ8udLhsnKMM+aVHpZDR
hJEXuOe51UAubKUf7cq1e8vF1ssxuVv89kEuxkoC78PvA3oQ8Z8d9inBh+yjJUlf
u7ohcWHiKgEHqjPRfumHnGJ44ePbR5W3ZywLFDkJcLrGmlX5V4nDxRwlu//shwvT
FFzVNsYUFSC6oukjeQlDGPHTJbPeWuhPUmv8IiKz3dap4pZl1D4hUGTzj1Uwwwa6
GkIuECLKfkOj+smo9GufZD1ditLY47+DlQ5Fz01SZ55LGtQrpn06QPKKkh4ZMWbk
GkIQFp4MsxlobVIWYHj9xFOmdO61PD0/8EEVYt9LiVd7TBMLez91y9bJS9Kw1j70
zNcWlAOziTQlAJMsRm6hJcDRnJWbfyxzt3aKtsqPGY1JVP5UhanYa/fvjGt/x6Rj
34MIlZhGY86irsVYXNwW5jchasPlTn9leZ06f1zhsTM/OmXtSkynXgDfCpt8Rb3T
4lgh1LY76QDYU0qY226PmIiP9KWAU7ix/w7G898ZXuD8iVpCqGv+vGvpcUqXx3Xs
SU/tyw9RjkEy82Ru2Qkv+8+K11rjM7Ea2f+ENT+e7Ap8gyDkkFeUJ7SyZ0uce5u5
OjEDnZXHIq5lfseoxIxMtXOmMs67hRz7r3W18bVQJwx0iXvzwgZt9fqOEPvQCeqY
8x2HCdyxTNE9xJkdOPgkK1EpqFc2xJ5UUcMuPQKLoX9pP2drZQflXkvMAkNsysxI
76SjRvYQpCsnVvBNP7ddihkLL7yS8FDbSTwdS7LL9MkkDmcJRhk93nftX9rbYzEG
NeSQOg8MQAtVdIlzTmSqH+qW/iqX8FdV96ng1DPpQ3QzM+MvGJUY6vH7brLPBK2F
VFWah2cddjBE1Zz+UMJlrzr0afF5NYIVDAyLsbFKtkRfh0JNky3cYOZgIjuABsHx
V7IJCryyE6kcj0KBSGv0sFt0mNkpb/pqVdyYDZtzZY+Zy6FQOrGSEVYxvshm6RBi
8x1vOGPPWH9CXkgmEF/zSpr2C/MnFUPChFn+gEprNF0dHGGxfChYgoy5Lb3vCCEa
G4rV7VT3AuzWUD9g7IsXDtZ2Zrb1ve0r9OYNbcQ9w1RioLlZIJT/6wBR/K1fpD9l
V0yfxJcCtycoI15rNb6kEIm9oj7Xfno2V/5G91nJAO73cHB1ReuWpTxOdd0YG+mE
tB1JGmRGJFyshcpdizuHlh38uWS+y7r8pI49p2Po8u5LnEHm229sTHBy2RNWQEgv
GK89pfSIj5SQHGvPO1WpedObJBu+1ZN+Twvyw29NKBzENDrSW7uYwmapsmsH8fB2
IxWyUmgJXtTl5ImSwNg4zOmaSFLccnnhlrIO+1s4Uv5PWpmFPXLZsoIv6WC1z/H+
rAhUQsTmaLK4QgJOHEL4pRSRven5oPJD0KBy5jHPVheZN2GW0mxK8zQ6nJcpvUct
SbpGZUs/oBcUQO+p3LKlCGq+zQR8CzV8SbPvIJzjlJHOmcJQFWx3uMw7Z5ixkRXM
0ZSZ+ZUSDkSgCFxmhAaDLCHOEDR1KCOyU8EAqgkiQALRmJVZVMbYN/RKxcTABatJ
6SikU1bfZTjdp7lSbjkzgjv9FZfI6ARDbKIH07586GGsU3Zgm8nfQnAo65f5VApU
uDGrRri57aF6DB9NxcbGSYbjOElMtkFlCpXRFK7dagzCZbxuoBvYzqugDfNyKeSU
ZCkz7Ja9V30tQ6S3fc5GKD2hpETnv5t0s3oK/FK7M6JSfbB4xVUm+yw89f+VteAk
urIe4Ps4zFhRgMus4uyONcnNQGN+j2wrHpBev8xhoTz/wWojUUesix/Cq5GrlmT5
QWm4r/bxYtetv0JjCMHYaVsH0besrKOWY7EUi1SNsmEnAv+pxiyuHJCIECglAwMA
I3cK146rdzc8Mj0ChUx82t0RIRQLgd3hJ+bom38IJO39iSP6XJqLIrHMtNCdQxRl
3dOWlE0rrqe+RJ9zQQagBHNRO4Rjft0o3ZNJfoG4NHsVkrv86aq9mNYCcoAwyiyI
h8TmEuyRGvzs4Pw/lirVb+J8qghrKsH64E4hYsuFF/EPkqeP1Yc7aTIfXGYj1wZ/
uWWcr6hNnFO5PjrvqmNjv1+mHWjHbFvxfWfHZ9kcF5P+Cg0GBDA5lpFjajJ19di6
sJ19SOwud28s5p0Fc5jq/yED3XgJOVE6kHrY57WIywXIKIH5hdk/KKEQ/rFr2w9D
862rqUTZpFUO201cljiYeqemvNM6YAsU1m0SFzf7BXyGTCJMKaP9sA9u/EWNWvd4
8WHwtRfWHH6S7oWr/APjFkFtiKAu4sgYzdZv2LCtuWvvCSUhsom1Yu0KweV4SRSt
Jlmst4FlhD4rEevKxmucOo92FjLiXN3eJXwCEJ+uIjC/VPlY7UqD2sPcX4w26+YZ
xoDPiQBoI6f8e6Fzs45RyM4cXw/JWDX1QIviiEZiATHN9CHT5b5Pl9214ZSPI6tY
gTHfzxUFZRJe+vp3uEwEnRI7AVjmIWsiFp9PWmjm3fKqAvXD15AwxRCrnYti4KA1
9Cu1BBlzmxP85hANHNlBGDEYVWeia1U9hLctS0WSVSj9ZqKFusYL2I1Q/bWFEqBK
Luxvf5nq7+Rpx3MoI7vEwPm0JQWFVSHo46S/HdxfUGbbwXDEMN0EnXCbWSQCOf5s
tZh3s3+/brULFx8WoyfsXdrDuMlaLHE7XkQJY8rL4EKc/S6REd7X6JfBiGSomIXi
BgBxPZ0c5Rp8F9hldpVDRWEuAMDwESt8jjeE+1npsTG/CS0HXmqDa5OuDs87Eus8
YzetWSbQf3meu6og63FUBtRU4eY6QXjN5UCNtVw2Yxb2xIklymD/p5bHedezHm9k
klwowXXw7MEo7MgiUyc9pJi1okDVShweb0x2555lq9XX4Hnsy9LtWXGBcna/XFJz
BCAeJ/FtWzfX70w4eAvdUlHE9c5A1nO1K+Fhg3MVcBjnQg54DK/rnKUI7kAb0kAH
Jw80ESfKSW6OJw7kqKKCVIG4GJFRF7OfaA4kX+KMqt7zjRDdXnLTrwIZDi4zOTx8
PAIIUoVp61JmzqZ+NsWgz3rPWUgt1wTXzviS7aauDuNusX9JsFiDe+5GUvkczLnH
wACMbtIO/wc26DvFT6vWDwe2vdFveSb6hgciIcO3D8rQDZyYR8rvicin94vTXXmt
F+W1CE+asloZEuFsV5mLD8yYfIG1zLgQUDE3SNWR+6++sSan4/1UafLk/N869Jsh
XuayznuJsWfq0FpEzzBZCqT24tn8rbAPSzDNE07VVLDVIKzLPJygWAPrJ5Gkxxrl
hme2BiyfCj8JVGV+OHvB8LNNG+RfkHedFaNtcK8jm34g8AGnsIFIrvvnkjxwmi88
5i1P+AiZv2HguYLB47Mwmf6tn9y2UMy5Yzj4z0exLM5bO353brVyeELaiF7JTGw2
WWCLW3cikCYvhhHZGXefy3ca9qdsLaBlvPPP3Ck9Nu5+BzPKV3UucXIAhNDYoRqS
rXgLgikHAQMhdj14pAIroBFJiYOp6q99rMwYPoD9zZtkZjlGHfETDKuSLZgyhYAH
no4SjzdhY4ahJgX/Uqfyc5WvEM4spzcdYpAf3paAZMFU4IzEUas3rjiNbWPqEAHx
H0cviJpDzbBILKXuezmlr7UusB91f7Jk+4wQNsWRSMEANiUsNX2cB+OXl8wDFXgo
M60u+bzTIS+pmJTp951kuHRDASujOR/IFspiILVgh7Fwqpc18lPMORxf071lq+Ct
jklhKLh0eu1xNf0/ex80wpqsFlrVWOP2I2rimeS+8bljJSaNf8pw78uPXO64vR3S
PiD7uhRsxlEAZ75gg+7hPqzZTNAljiEvmuiKPDe3yzdvNKINuLQtLPJ3J18MiAoi
8LtlV3yy/wJUrvVB8wEAsDvtCbVd7pxW9L/RK4sBIWHiNz8wYsy21uSDbqgySgsO
yLY4akjhIvxjGXbMtesUWAhiQpFKvok934eZukFurLyK6XCwmu4h/wnL2nUGnfLV
8bk1aNbYQ8YzSMSzzGkbYXuoBsui5fxR2X2wZacwL1kNW8qx50iVFPhI2Y5yEG82
w0tP3xbcPhsjTJ0jOSkl+WV29LQg5/Tx1j/fjwlZR3y4jpPnLCsHXiI7ATZ9ePBV
r5rRuxhkuVDqpIV3uxNEp+yD+vOY5eIDn3xBwXmsRQFZNCiZy5gBlK4QCQQkDwqU
VVCMu3BK1tssiKUF99f9bMdX1e6Wb/6x3UPIZ1+Xr3ijl+ScIzl4herBrrasV16k
1yM1vnxYzvAwWi2EqaP1A5QffzTuNeMxBehraeA8KnCRv6ZPJmE2Q8nDn5Irc+HI
F4tllnjP1Tp2z1GTlc2Eq1zC9xU2Fhtl5Zhxe6J3nIMC7UC9WqZE/6M4lw+qeDGY
KBd7O9vwv8VZ6BXOrpOJ6EfxHwKd8uhsmBixsgIS1S2D+jPMluxSGBl2Qyop8mTV
KoBHiYoUE/AvDdSrZYP5y/qU5XmPS4ZoLhaZujdAncL1vkg9O62VUWG2XWrDFR0c
VOfTqyJ8AkJ9bLt+4OcEE3tXnR1ygLj8XGz5TTFg5/bD982SKo8e0eszdgmJiU8f
zFsKMbqjUcjohycsGyty201cRsjVzJ5yxCmAgSx8a2Zxgpjde/85rY3ZfTDQa/gJ
WIqYaihBoy39I0Ii1fcLYwxXAqndGpduruXBtPgW0XRmAi6nJj1HK42Q/dDyimjl
eKxGWGULYsKPgqZvo7enzxn2AW50pyr9M3LOXRss17gbM4qgiwrJbRWvvzGqAi98
R0/ya0F+N4MKGVairEUQwg2OAz6/htjmQXk3aTEOKb5P8GKAGQNC68nm+IcIbGk7
VVmyT21NsSOVVbzResdZXyXhWOeXWEx191em1dHyyDRoR20zQa/suulwIwPduRrC
0zi13AalH41BP+jgBFBSILC5G7q6qwzLGyQp3PRH6RbcroF481HvUC18MWa9ogOM
92N0RCW1IMu3+NZbI93+Po7NN0Hax3pgGXiO4i2d3cv7AKKS4337uxOFB8aI8N26
X/y28q3Ak1iLuMWEcTkMcRUZXKt8R1eAzgSGyP0RSs/asoYX4rkzoCRxWnCs8Cnx
dlhprCSLzp3rKzETOZ2sQKCgQocqNHMax3y/XP//3BvbY9tMI+Al5e7Qtrj4asPu
r/zuUeXTUBjp0v7ur+W7d8xvU13BqsOL28aQ48iXzkOK+8JRhBSZSC+lxXFyyLJp
4W0eF1ihY0mkDxfYeFTbcAFRv7yYe9mFBFd+NwJrqThbMEdEMlBgHfRrEaacHI2x
l0DEM1jGkWBsaoNvLf+AnmEWWkOcMr3qmoWmsYi2t84OC/7SGTv0hVuZrfw7Y2Rh
hkA3ApdjzIa0LnCnMRbKQJdgqMCQrW8PCYL+EdQZDdg+2U2A8jvAWco5DLY0LJpY
fzfP5e59SDo97ULJk1uI0ekSFJ9hJOn/FMk2bIUf5egc27uuUTgzTHNmmzg7haku
1ejupBCptauWucQCVQhcS1ZoA1IwimVDF1/zjj82/3Md/PvThfFuGCTElnRZbAr3
W4qqxsx3CK8zI2B8ee45pmLrT6+CTuZfafXU5d9C5ZkJ2+ME52cXIGxzE28IQKAO
W2iN17S/2JBIYL4pQ8H9VzxmB/tgi379vXgeWaRMzoTk2Uw5jCH28H7TivgV7qF4
ev+emP0dB+J5F1Zll1E8xkuWT0eszKykwaIYLJZi4+EsXRILt49qjIvWBFE6A7w2
IQ7kNGMeJ3qQ8xtvi1jxfJkJeNWdRbO4lTX4FYInJNXH+jDaEDRCV5q9N+ukPRx1
NuXL67fDptNzbj3kCnazyrZpV6/7/1v37Xu15ZFAjDHOAHyK+smgNMGmerGMIlrw
BjrfwHA5ChWcaL2QCMcfaglcOrYlMgmExyvG60MJ3XNbVXlvBaCm5EQ7Kt0BVuv2
zSom26WjtjQBnbijOzqfvSKTnbfzpnfmGgRcDm3E/+MY5PmeKKsVfrnfRUxhBc3k
sgd6GZfyWAkvovizJAIfi+GDAU6c0vlM0soHZ1z5mtSz/1rkO6J5JopPK+kkytMq
wj/oMy0w3FAB3dB1wsiZ9od1BWLS4SkMZ/Hs8vaYK2MV9DiK1ILvgY2poxQ9r4TG
UYf5JX5IGC77u7/dsRSqeYYlxfOrezXkBg7eLxzF6fix04aV9VppLw3PnZY7Wv4L
WdeCBTbH45UBbthrxql6SxCfhJDlpkuAtZJgcy+s7agHIqjHGWz7hyIhSjPvMF15
a3JM53eebVgdH5fZQGtI6Y/JVnJsryUa+F2ErbL48tyGf2uP8lTuSsjTV5F145Wq
LtVNpPcASOGaoi23mSRfSfh8WqdsldhQn3tyJOyKsvKbL8YL7Nl8ToIreufkKm0Z
j8kuOCOu/w2q4YZUvl1hpNNVHn1OlP9eC+se3eE6tWx+JgF3Iw5pMHpUvzMXAjXU
aO/yIPihRjPK8fWC9LFSpan8x/bTBsmH4cT8KhBHbrzJegESwoBAVi2L/i43kryx
E3k9mNx3+fNMtnClrtKj1zXiSXjGruuxlPMkL/prBS9xA9hLxnGwWaDcNk2YdrBf
OipgVeO6zicAzkKVwRRuwRJrOe3l9XkpSFjv2FbagUrmN1ahjIA+X90SxEexBEAD
To5WvaAHFdxd+KwJvhsWSmdpC5USpbNecYgjJkhWvuon96Lx5lyFI5aFS0g9VUR3
e1LBPh6A3pTZxKH8FmZ3Zc5BlRHy55FPOc/bChxEpDTcT0b9fZ+5erfOmZGjlWEJ
/ciH20Zrr/eD84vQLGvBh+IWEbJOUHfaLIJVgpj9H6TWD9U5ZqPk2q8kgIpBA31j
hICEPqtqUGBSG64SatXz3sMQfw57ZYBey7p4ZtEvafATzastt+724y9wYw1lC1e/
USuhzt6/KpaLDER3y46vgaUrzi4zOugi+JWw8zqV7nVT+f964fLOyQOXAl8JjRyU
Ym9jQ4hf0KX/kx2Tlyp6Ezgr6ZIPTj8jNxkYFw89q5+gVCT6sl/Z+xxE+6mOg03j
RT1Xsq+Wb72+D4kPbwvUbFhCGrbOUpKDxdo8K6mhG9ATZzF+lvCBeu08xl+8p9nn
0UDaN1M5aIh/Iyk1Rjig6+/FYiACw4nqCezXljiO1k6/nGaHAVfPflie1cQVa9sT
E51qDOOz6t/cnRQB7iR+kY2rijm0UboFWpygyjTIo3D9Sp5CV61ZrEWlc8FYLzQb
PB1q4IXrLTAzvqs7CIYmvfCVDaJgfhNhZvoeO8TAYic82rP4zQMtDFRdOikC9naV
8ygp7IBxYFOp4UY3+BZ0C4DfqYJqt81IL7U6YmMJv13sht9lZR1EhLO8UnOHZ61S
QRRbD1lR3KgOfQA2uwAP7+rDT0S65oS4Ch+8xNc82Lut8PmtesJ7bdq25UCddCU3
m7FR2SPY5Pbqf490OIj7ivQ2fD3XcZvLgecjrAH0qJbQvrZ9+WJ9CgJL3k9Kk3jC
Vp14Rh9xdn911bz01X0mc6H3Hn3EvLVwwNySarwacpNFRk6YDJ5uHCI2Ma1yKISk
xNqDbEkGg+zKmMlUYaqBS87mMj47auChLus0/gE8tzZkGWjh6JIDIezqKY+OXihA
FRQ5GABNDWmOAw3SEgf/6MRyKi7lY2h5NjJg9kKhBXlFip0RXWczFZfgYbt05ahm
uquoU8+GpvOIdczeOE6ockDqKA7noiY4/X3V8VUmfnwRJuJz8n8xnvRkxq7hbN8h
vn95INyPEYU9870vdhB2+xPPYGRCCWSWJfR/ixDUDfhl6UpfJHQbp+GRNmCQ0S7e
/XUO7A8FZXYTibo9LxCcZo/XieijPMS8bozSjUbrMawSyNI4yP6UL0VQmaN1oiEc
idjMoec1cFGLXOq4KNrRYZpniQj6vekbGxQWdrME3pm7b3NZXwlL7aqq9/r3Uf0y
`protect END_PROTECTED
