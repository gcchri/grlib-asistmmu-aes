`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6AJOto0VX8qcRNjfx2psOOdsgcP40eti2HChZW4dOLN/GxVXijZfXTf9dJ7f6oSN
fTN8KCuQ2rO9Xx0jvE0sKASEET+IfNOt8xviWerVzAD8XLH7scbbIZY24GN07FCm
PjvReeBMjNLGSl3pvScbaOE5+Sj/xas5STYgkkrRM/52sJtZ26dhUlt10C/op0mv
wPGGiGBs2GEIGtMrFoK9ZYuxKbM1h1mKYx77rEJ8+G+vWupANXBPjMK6p90nY8GA
DjfVsbxACl9pHZSWpqxN+G0AcvyNTYtKhtJXjyU9emS+UVicKdJQd/9w9h+efRh4
XShBNOiPKBt7wc/iNk1r+K1eBFd8ye5UfFai51KPEQDrRIj3ks1vOUzjMpnq1X4A
4ruDqoFZ1YcfeaSBuXGL7ytLO+hISiVHMeRVDRirqiLV5d1NFj0hI4PJBN2sLoy/
kWTt5HjJXa7XSgS/qdTlSLR7poks/WPpaAw8uFm5f1vmpdSIKQJ7B0yALCX/Z9Ch
6fcx4C/uMRyg6XmyvFZGxys+zpUP72SvXbzvH+WKUytgNKgEX0OSnojszEiXRtYx
/z81HSkBQ56SWLldtQBh/EzYz5nIw64a/T/EGPb64JSCjkxbzmHLMOYooNZhGJBr
rKEwXUJE44T+k7APMJn4pD2THtfZAqd+FVML/XBj0FlGWyHNFbVZu4VQYzvHHyyv
Gg1wjVmyeGOrMA23zccqYwo69UVLoyiPLWNfgYo7T5CYYQX1U53YUcCjYXX0g694
lHKzn+l01Q0mXxnO8HkVOt42hlbuhHaulk3o2+6mLBVWun/eYrN7i+LNfrS2gFeJ
Bda9ollhpvivJ1qPEl0+4nbmUwjtNwCzgkCjmA9Z+F2sRIkZe0Sce4wUveyMo3dP
`protect END_PROTECTED
