`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d5CXGYS/ZKXxz7a7NDc4RWtJaTB2UyU8p4aVHnp47pcQVcjLPRI1Jp/Ckj14xb7O
/mz+ILZE5mMs5EyCN569ytL/mUnfl2tZwRzuiKlsX/VRLtP3LgnuFv83BNPKXPdb
ouHG+k8zvUfLBAYh9sxigkYjokWpiVhzBkTM0nJsoiAUXIawYfJuqru72iyN+DWZ
imdk2QWhHfZmAwWmbEWspCuOFycDkuREZEZ+Lw6HgPfi02yYO2L/9s9LLofZuOJE
j6/kR1lKt7gUHKvIrus39idWGvE8WH3dmlo6UCyYMC+I8xQ35lwtAtklRFkiRVS3
4tAKHmQwiNtOeilLRqxYHyBESvZSBoNgB5htpsEOt7duqH5PGzLyA6eQhJ+npTGZ
FuMUyyczdaAncGI3d+aqVGfI/sjMa7/3riE5NagVCHcCZz1O1kUO4qc0LAhspJkA
ahKJK93ComUFnUMEtZKD6Uk7PiKZrz/D6JgAKvzvRTBX7D7vVGP8G5v0sLivVd/X
6utuOuvRZynlR15+9OhsKHy5kx9y+p8d2s3m2DhrqHr7XY7z8UsDvozZ6AKl40tE
KZw6xJynj+e8Q9IaqTTG2L555C+/rXVycEfmjbB3PqReu0ZygVILFQFaKQH7Utn/
`protect END_PROTECTED
