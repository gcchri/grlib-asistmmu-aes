`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sNNW3lrvG8PX0TDWd7o6E1wxqZROKKr/U3dvkNnuFTyiz8JxxmKMebG0CaAKoAau
j7tG4Kl1kJmCofMRIx2HFP6+480bEMheRB7c0Qs7/BcZoxYC9KpQDerHdmefDd2I
gD1sZ1oSHGvC5sFrFLuQQ/NFi2hXvFlq/G0uJksxfuPGoj6iHVWk0EBvWe6pU1mO
sARF8l0RA00Jzuvk18l1lAGaHn3ihaZXci48+zVucFbjLXH3qlCIAISJUiYzwT6n
W1fvz8SDnhBRal2R3KsFRXyLvgbubu97zE6dVlNGrRMHab5V6YnxD5gGJsp0SeJu
+Eo2mJLwIUB3iBZHcw+bZ6qB8EUcvmOhmWx4IHC4pGYaf1D1bG61Sh79t9hYX4PE
ghL9qUHJiuvkU3ONdHdhjx7CqnjwmM5DoBc6MdbS+IqDSABNtY60zQihpUEKf0JN
tYE5Y6JHzZQsOda1IILlLD2E0xKZiHBSYKqfIxsruiU50JeWKQPGnWBgOwgRhq5u
9xFMbJfdq7ZRJyAEgh5bqPzROuvq/aU+2O3fxtWfjp9xU/HdhGKSX3PMm+aaf1JY
2vjGLKdhs8zjmFUDkNPcAzEm8nYB/aVDLXMzDgqS7d6MZWnU/t7Y25ntEedMQ4Q0
p4FZaYpqMnR6rBV4Phu6U4H3dqs07LHd7DrMn8Qf0OzIzmAvScNyWI+Xv7F98x99
GSK6oaI3RykSvGyupibdV9UwVRCdqHbecxrhwhcGexRQAtqAK3S32Ma4uoljEKO3
eNmqLKSORJd/xOmES5u5qpiPOLTyUXWi/m2XU1/I9IwS6LHCH6C7QrDiSJ2476gj
8FfNPr3nT55A6OahbOk1zyEsdwtYtyMSqOXJvKCb5V05EQAmpCcQrLXcF3deH4Ox
jxki/+2Z9Kaw7Brq3ei2C+1hxLIgAyREdkyMrtMD8t3cGhjuo23edH/ZOyLAEgcl
Sub5n2f4+G7rZVnq0wflyfLB0lrSJ2UGQpA5AKGibtCSFeD4pjuzDm14xAObK8QK
FsfzCDbMzFYcWLNOzRKzznkD5HGE0UjFiGQqFeQ4FA9l33YhpPSsqLLg/mmlq43z
BN4Tjq978B1ZiKtGddXTU5ZSDqqpyUvx1AOLBLQ6OPrPcgSEbgV/OZXlbUCAD+Bw
G8MjVtTtXtcXsCw9NF3eMtVsSldp19rWS38wZYteXCze3I+SuiK97+hUU1ViClcL
8+Vq40//E00gkHPy3HTR9jXw5gr9uCxVZPXB3Ymoz432PlZChR6W2ttMRRH+XgRS
LL4HYl4DwOuz3k/aDr+aRdte7jdAUQeetD8XkgT6w7K6UAJ+1m3tyDMhxaZ2gYwK
Z4uzpEI/2hdJryMhax4ucXqi4CFXEdpoczVL0RjFyZ3hDkkPrqpnzkNTMHp9u53l
tBNRx39SbRh4Xz1le66LOXxA4Wy8oTcrwnq0PpZJn0WQhpp26jcPL38rsTqYP6On
S0i5TGGeaCH3Jsa9R3Nrs7Tu6oZg+y4K8hN7r5Nc0+Iwug4FipGOAS0RR9sB1Uas
YhtPKHcEeyQGN+2/Zah3sGefgbiccLx+tLuDaBqz6THLC6ECPpomUI5yIzqCvcIj
G3mNTdw9hgatVYL4b0TMDpYVAZrknxHhdNwSUVaACwX1Y7Mqlo4YwxboYlRDlcSV
sIkabEzFbrJmSnAqBXamPO2ZVaO9ew77gdeSYNrMehNJB7GpBDE7iS91enan7y9w
ZLHKkA8VtNWbfr8EYQgo3fQ9OYOtbTYZO+ZA2+NjnmbJjc2ccNTZq1O9liAzuS0s
css6N7KXHbCmb4ZCIiCfrY84FL3yTw2Zp72EgEnrYWqfBExUSCGpnkd5uLg0UzOf
lzM0/GmGrLuoeOrtNdm/GFTc6ztDPOOTyQRKw6APk0+7E8IMC1/CBlpwpZ3X4pb1
ZAKY12ohKUAHNDCfbQr0Kc+s1ymanq/VoDGL2pywb398P1urfofUPI4J0Byj+8U+
r9MwBmn4AJ4s5AMzE3hdkC7h3I4tv62TWu8TmGPAtlt3BA5MJR6xVZT/OdH+LR7w
pLLDFG/ipW1n/Lm+0bHQd1N1f16gVt15itiwU/skBgGTDZI2WecY+4Exsd/1bh/j
MgAhRmGnRkXR0WenwKDMnxHuqkQQZwVic4jkrXmIRgaXkJYTnxQezAYOfmVYSiQj
mW+ulrbpFGwPxnnxi4N4QjQZN5hiCmVSJXwZUUEzfYmuGVWOi0ZHJbNEsFnZfAdT
mzx6Ox8ZJZMeEMJkVaizzAp2NI11WNSi7xK40hn+zVIOl5hA35Qk5KGZO6/wVl3P
5JdUddP8PnoYiQ4zoauwU9/WnL7srxZcZ1fG9wCchIWLiL8L4e3J6OlugtGJKC5G
aj/+wjEFnOvKFG5zz76+YblJVNzlwT9pAig5k9MAyli5//bVT1dPzr1QKypy+GAY
dnefLtdJDQKyJboVtPWS+boPnkWCRNXQszdq2DdJ3L9EH0Ikujw/eoblRIFDkrlh
//vXlaICUx0MfXuZoj1obhtdUUByoUnkZzXRXbxTbyOxihsEcphtS+g7lCkjhqQc
fw96w3N5RLNQUDY9QUVOZp1hCaJTr1XcL7t7OK7t3M0jd7fXjmYrBekgo842P9+k
/AVbr0hF+RVqTzpVVHCkezwVoS2AHOXVGa6t7g+hzquHM63vE5gfYaLJ4gnsg8we
lILSF2xkc7B3H/DIoTrkWpqsiS+P/JQc/srs559qy032XfKMORJYN15KYlRAG6ze
NXS8t0ZsIvS3gHr/s+oHEQ==
`protect END_PROTECTED
