`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X/ticL9y9OPl2jpPjClq+ZVt+lR2QstdDUnISQozJXCVpLv37UhUslYR1fj7qV4F
M3qogWKM3n/bj1P/9dgHwKfYZ2ISaAFTm9hdtjytIzMWyo7uwlwdab5gxMe5y0ff
/zXFFUXnM2PRAQOKXsUZTW0LK821yPHWTkb3ban6VsxecmAzL/bHR1f+uGWCJxYG
LvAG7Psae6Z325FyADv4hTwxnU76vidq1kPeS+3iGaDvJYpKnbz1Hn2RiaReSkBb
PQGEYtTpFI1R4iw7ZwRP6iuWTIl4tufFcArFNAyzOoj3+cMkWgYfzwHQ9ohIeCeN
HTExmcw499ReAVhL7iIpT2VELdeWjL4vIMn4IazRbBEiAVImPa8V0ThGs5SJMGoU
+ZHRXtLnRvvspvU46mqXvg==
`protect END_PROTECTED
