`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NWoPDhJQtVh6kTNITbKaAv6WPrIQAmwW4ayk+GGAjXv/PtwPDL6fjy5RTiVEKlGy
WLCG9WQ7sj+XYQtkYNArcdog4kOPRziyfI0fbNTnu1YchmrbDPfyjMEg/DBZiNU/
huaikx0vCJdC3iE705L6SQwv5vrT1RbwLQCYtf75b4PFHFke9LfH7RaAX8BxIA7x
OFkx3HFzcwUR1MRzygNRzYZpJlYUkVyVgKbQbU9QFZefeo4qjiOG5E/tWSEl1ozQ
T2i3wo/aR5klet716eY/M0D72O2F7cugH2Nr5F55yYYU5bBmB2tunGCNJWXyCk4b
NO57oyrnkzRLOO+D57paevCZza9CVzMkzDQTKIyiELlCP0bjFGFew5lMRF0qtKUk
rPr/MTPUTC7GkKwfkxsNGPJV1vhUa59N/G9X4RaxpPv8NfVJc/I98gK24wTf5XYm
Onzp/kT5qqZwnXlbMbdk/zapHzLLUZ/Re1o9yX3JI/UdPAMC5j/il3YUev+M6Fyj
Z7HBdO4rykb6x7WtFTgSpTuUTuUtqIh+AFgeAf1Q6B8=
`protect END_PROTECTED
