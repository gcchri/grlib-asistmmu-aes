`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
70MWmnX4C7o+ouIxx+OyKdO+T9K/LTmyot97Zw5nzKIqjz5RU/ecQ3U5MDFk0eXm
cm5LZ2k3+KADGJrBhgjp79ppuXUVbCf2boTAbRSCfXrAUmt7qppSipAd52uzC/Ri
QjQCZ5FS4T919jpAMBXtItxVeB8oRmqlX7PKWTduSdmSS5ArtvRDBqRpbwQvyzot
UDul+kFS/vaiiRQeggguJqjTOeDexWV2FqSdVst5Udk7q/TTqvqCTGxjnfNzy8Xg
Dj1hg4JuGA9qRtO/vrlF9GEENmATGKLAZm/rr7ZfL7KARueKbtcU3pGyOdHNUwQ0
fLKRXPelPf6GEnMefNdaRcZXHEjPRMC2vVFd02oZv3VkMlPtE9LGYSITEUTuYG7V
`protect END_PROTECTED
