`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
41pqTeVmwpnApRWkIwV5jTCw/sB9vnmIVLdnjuf8/oBUkL/o5HhxeCH4zdA4ztBo
OAerk2/JWQkSZA0k3vgGcx2BZetVXcEMjL3JZJvxYN406wUSC2u/g3Au+qUNhEiL
cfMZ4UH3JXD9R6YF/wV0XpBTq/NzL0WHYyR1VYYJuwW1eMIr5zKcwU3SlO0AfTKF
YYQETFB9pJPq4L3aXApnp9RbKzred4bKBi7lePjCPqx2Wz03VlB/psHT9YC6Ve8C
DD7EfgF6o0B2EgBZEyOSCTvnPeHHP8jrZ/N/32K5C0KM3YH9W22iu4HHCrLooIYQ
6+HUFtPl+6clgVkqr8o8gCr2dJvqO9cAzcm9DSCokrLJCX/oS9bQCKR5OVqUlHWc
fMnQb49jnZvh0ZyqvIlcrQyR/6t0QesW9+6BeyNIkp6rnhoyhmvJMbf2OhCtzq8e
g1imSxRZUjQvCc1QgnmYIvcHvwcQ4R/ephjD384YlYNib1gML2Y6keObfG/4KbZM
FrKTsHtDopfZw2HKdYNbXSWQRErna2WMYUg5DhUe1/Xep+hQLAzY5KSR41l9rNEz
c7VlfaQZQkl/fyBapKDWmHmQa6ljt7hgKWI/QBu5ExwwvXkym9G5kNs3AWcn4Re1
CvnQq5aHj2LivAY5N662Xg==
`protect END_PROTECTED
