`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X9ENEYr2+3GeLMQtoRkyptbgwHboPeKS7M8nqn3eqMNsupWy6HYEikEU5X7gDXTt
mHlqyGPH4g0oNJW3tNM11INPRkE3TCX+f1/rFeRHxomCMNxERZIwAmvTHqoN4ANb
5ZC+wL6hd7TVRNXCG3EEl+M4vDnzih9sT+ELOwg2Aig+kzCqUZYrPG6F2wdfsf9b
bndkJa04hRYkgA034IfO44EI/bjX1p61fUz0bDbzrbIaVoD4HHJLBknR5ftUuPFF
HVPNkwO/hbEDYzZZ9vqOdLh4NSLcPzdSB5pUArzFM4EUdC7TNikLBTOYwCd+oTN/
WVmoVViE71Mvdgt7u5WGvwS3qkaL7RoSejtU2A62dKKzAN6nUjy+Irzl1VKd9Zvt
Ao0vMMm+iJFJftAyIzF/WGJKFiFdMJ08gQLK+tMuPze7MVWraxDXNSt7yOb7cgPN
BV5hlBFWIGwlDJiwW/BTJl/71eWz163Ep2ZkGhudAijm0dBsbfX1vjVpf1+qwKEt
C5EItyw/3Dha0xdFW5YGaVS/CWKu+6ETSUL1mSx0sBTDedYn3N5QwCXl2nsYZDJl
Ls+WzjChmzmU7QO8k0VJjgzAX+drftyuowyfb+EmeSVan4fOsBdT1dehW31ifZ1C
0K93GPZrl/ewog/U6bRan6IDESpqHezPP4Hqn8rTIgq/f2ypcd351oMNGlaD54Vg
d2NxDveqmmNlhFBzylfXlVq6fk3+ajN4CrfCLkQPjA8askc6SsxWLgUPrfD2hNZB
4W5UCsEnB5zVsQ6FZH/MA8viMxcPbHhZCsJ92byRL6zg7pfCuPK8MsADQ+plIuh/
rlbTckiuoN+ubU4k4ryVqAOTYP7VVrHUxxQOW838q3LLytGk+iNch3DbM7G2KuKd
2tPks+ZAeqeP/B12IxkQmeTnPORDmmMZVvdieDXhf2+I8vuMFp7C+NLz7mlQhUka
meYeGJn/ZUqf6FmYWr8m89i6IhL5NMHOM0YbMbFKBA12EHxXiMUaxl8sAkiKLkLs
y9/GXK4ML86psv6cLDewdtDwWNVWetJgJ6kjcSnKje2T+bTXFzh9ayTX98FHpF4p
f1X8roe4kKSaGdjr0Lp9A/jFeRh3GWdTs6hYvhJd7XNqAWilRm4PpSTd0qKoUZI6
kDiYJ1cFDYtGDSE9ZGup/5+6d0QYeBHTck7nV1nV0mdb0biiACcaFhx7MTF/HiHU
rSyOZFZMiuhxKLaa0EcLjuy3ddmC0QPNDY4fCUY7sa9iynDU+t4mkVvOT57+lYNq
oGA4gdaL87JI/YVVGZNtUBxRJe8kBFWx+qyQAeq92H9CcsI/VTT6nhBTm7uv/FiT
9cXlHnzYJLigKSnOQYkBLwPVM0CXflbYHyOjYZf94skj5rK6PNrJlh8trPBNWe+Z
Fwf8DyC4b2yrNrftSruo6JVwdZwCh8fQ2bxh5HhCTvhkc3EOfwffEMrwnf0Q+AZx
sYUomGBbohRhWkKnXyJfgJOuGuhPC0tAOHh8ck0+w/xfOF7GCXc8C7BJBiosOoDo
oTobcPF8wqmm8f9bEKp1ZrgbgVqJZ413vK+UebM2th/e1DCqzqwIB3tyNlq5htu8
aXsWp0N8EMTqOeDZBGTXlXciFzsA8fu1NOyeXgccQpap+LKfkuWgDLzKZG3DrjmH
d/25Aodk5QU2y2xqa0sDTzkHeGs5ggWSj7NBK9q0hVX3Wu63aBnqIhSOQX2QXshH
aj7qEbSifyPL1LzTEMSC8ZdQ6z6iAattlwb9eZWkeaQLT6H61LwWS71pz1n2Cs3w
2slH3q3JUB0vgXY2QhZrfW9bcVWNGygxPFqP21eeRLb7XSTZR7rIj5vuw+h2wuq/
D/NaJrAsWBPm7YIo5YR8mzw4Z6JUObq6PCSDpO0CPL2JS4cOvjlq48+36m5SAI/S
hdoodMi2Y39OJuVYIiRBzmviyLdugy4rjthDfc+Q2m5GoD0DEWwgEWsweJS+3RS+
9l5PCWt4N3vhQPMBb4eocfEOsGuUdEPgnsQKkgowVkgSeLqN81tc7m8hATZgjzWU
IW9j66Wuy8osF+RN6q/gm+m/I4pMi8vb08/gurei/1SNd0HklE9u17Q0foC72JMl
eWcVaWAAI6dxESUF+jtl2g==
`protect END_PROTECTED
