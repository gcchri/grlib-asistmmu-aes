`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QZTG3pa0GjuE9KYStZH1VlMJ8b5CeL4PFeaPe4NObO0mPgkHrghBtC9BHdOBeeeV
KIWEXRdKQIkCuj4XPNkEB29J8jWw8MTlPw9zj1Lv++v9ERNH2oSvxR5pEqKYBTCw
f9vGUF9p7eX0LKEh1bHtkrztww3habNtL70FjswNSK9JxkUSaCr6paFGINmQpDLe
U+8zLWkvgk1kXTRGUgTYUJgfKMp1nvjF675bIb5W4l+2rilfUAmPT9Cqv+8/CVui
PatkvjIsDqdGfVxpvzV7RT0Z4A3mqZ7Na68UyAp/TZ3WsEAMYNOC9+Je3BiepcwM
/khNCsC/f7p7wGAuldVn+w==
`protect END_PROTECTED
