`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uyX0/Ik46wy060ky7n2tx/OLIq8/ECwcL1i24WexnWsQbWiC0Jj007IASX9ezLdl
+0utGfGERKMG51fx75GEpLUmFmkb8LyQPXxaegi240klav5kbtShSD4MH1y16jtZ
1bvgBtA+ygQj5eoj7qvnM4ElvpS3LEhOG0gxK5fK8KiHl6A7Isc56yBKNnXhcv9O
p+UDV3SEc1vUlY2oylSnBx+d2Y77JyRRLMu9kBbqDGK/QugatEHZKNyvg4jo8Dgv
V807p6dHmb7SIMxOcXyNz7dtFbsiDDfSwv91LTpoGLN4r4KdutCGrj8KYPn9bSsl
OBDXMzWUwOLvgZKXUy0vN+4MBLXsh2ACTr830KFog1qjwWOF3zykv7u6pzlZu8yd
W3IDmM/U/orMtnbL4N+rDXT3OqAbkc/m+GGCkGHZZfkMjH9mFemTID8jyj01dzUU
2tnUnuQQ8a8RVXQI03mxS8JwP5Yu0mSrNxS/9kzdtYY75w8Nya3EU/yyPdAXetdG
UvUAsE8o5nrGuT2WbZ201Rae+s9g2Gr6PaS+LLK+j6EKsl7tcOfaYkQIaldKjbs3
zEpmcYCHJ8Z9ZGUUKUH5aCoNxktlNW+kgdULv4jYKBYrLFKATktCw/IigvbeoSed
z+PxO9mvmYpKa41R8DadJ5B8dlGSOed2QL4Lf3GCTzq18Ga9ks6OzWKyvklsTLwG
o2xaXCZdIRlr+sZH2OSROtFtL8J6Cy76OQDblcsdSLlENVe5Rr3/w9WmaN4a0K61
oogUru+3zuvtu4lgz4GOwjoS92fDY57E7pEogPsrzBjcG5W0uxHXMdPZVuhFQKMA
T0xO9AUTxSCWI5/LkyhXBCdK3DdlX8hE6+qxJB8gE4F3WTl3p3LLfCoKU+7aob5P
TfrdtPXItO+azmVq+BL/dQ==
`protect END_PROTECTED
