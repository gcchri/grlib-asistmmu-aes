`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UWOjTfNmJguNmNAkGtFD/+ED3kaPcFuoMGprilFq1A7x2p4pBRgdlhFq7vDPVQz3
aY6ZXDmxs6q/ckqdwp2kGU3EyqqEn7iYi4Uf2qX0azuhqI8LdNiacRKZjNwlwOa7
kauMEQ7vuG7HYfqYMd2kWQgtRWe0cwah5RpTU5ZiS1Od2q9dkdJCos/ygJqL8sTj
UqtYQlyNkuox0wX/13keTV/oFvrm1MRRcfHFHMT2Hcds7nXZk8QQiQfRHgh3zA4d
FdL9j3ky5hQSvVQ6EuyKh4DV/oqPM9m8COXWwHU5vWqdI/8rRPQ/HDYXlWQoLjwO
XMJXdf0qsMbsQiXN0t7InL81stpdYHrdhlK3/lAF5i8MrZY9dlTS3ib2x040tEE1
/anQTubMQmWaglVXdkNl1eUSd5CfgtH+e0zUu8W/vThyxnSC5ktZMwQmErJpcmop
`protect END_PROTECTED
