`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qvLRKqYxAPCwbfPR6K1zEqOA+um42NSThTb5jUn3fmc4/HJBTri6TER3wX58T/l7
UvUK+0gyQDrARi3Kfn/Xg+jfNTJYISFlNM+Kl3Tg1FwxC5fOuM41ePOlLnSFeyfl
+yGt8vytEluqx7KgEleznVJLiKhKXUDb1rl1m65s4cagHn4cjdo5nw10FPMu2Yh7
CQyqhwXLJ5W9tV8g/2Izeppxona5hV3UrsDv/em6GWX0q91zvhqM4dCjRDMPQVzw
P7Q1bICRBltGigqLIiu9afEl0w0P08C/Zat5mAu/zlncUX2UMT5VkD0vlQwqfHNc
UBVqRIkbiGQlx7uhrlpcgnQu0/do66f1izI0xpKJbfML5ru4tIJcqMQceaoBnYc7
kfJz8iH7wVmpwLMx9zCoNNCJVv22Ebkypl6fAKHSIGe3QddHYKuJkq6czv7GXDC7
Jknr5Qtg9OaXy5bpzzFxO3bJDxJ9B6anMItY8QqMN5addDcUFHB+NVW8770E2j88
DxE3JfUAFNP1DPBLnDNpQZBFpZa+OchShLRf7GbFtJINSUdHlWCrXeiYGA5YLSNl
XvDLuM1cqFV3eHiUCHUpwa65UA0/AhwpdIgbqZ/CVu4BF3IhWj4lfnbR3qqRUvLr
V2MuCCz+lW2ve+D4NQtoPOjExFGTLQBGLNAEkaJ/f5CFAdAECW5J0zvVDTXI4Efe
5p6kSWzU/uSclLeZhs9/21CB9KQz+8Fn8CqL4noBHDipeQkjJ7oq2A288XT5EDCX
NHP63ELr+LrIz104WMNCltE2Sj37N1ZBBJrq1678CdHFROc59cgdpJ8nIjQOULF3
RRPY/pbob1/l8UHAlYfhBqG74crK0OFuC8Suk4/IUEsqInDIx4mJ9S86r95z6hbj
uv4VpefTxO6dplqmpCT6ESgzbiK0yNRB4piIntEYkgF2ZaMfvls0qAzcYE89pyJ9
OdwA0Hi7AvGIVvKZiKNhWPHhbMNg9nU0SJ0KHGNz2rDvQAfk8dPJZPyeJEir3lKz
j/VQ2RlBt7f8TeySp9UEwHQoUecl+VdaHthw4dGggWTPR3Bkf3iuS1VkVZYUZJpn
OFrI3WzLca5qAZB6LCT79ppFVt5mxOfo3h6sSUOpmybudoKx0BfFzf8ynIiASpXs
+OKhJ/7kixcmaOA5Leg3wdD29g/+Q353KBIImODH1Iuxx29oCQaA7oCNtVLMttPB
gPoQ9UIE8moLGKKcUhHbU9ob5FnGj3ur8jz46U7UEVzYp4wKj2MV/laKz3tPv1yT
h6dvEdf8OD0Juub7pUBPbTuM90ysikgZJJ1SHDtq2EYIo0yWjRYQLyY2TU+M3mjX
rvUH+Mzcu36KoEgxPJOf+zIfOZfIv5h0cayBac65+g2S+YLTmMATNPM7iGh5+5Ck
Q6RRjk+1TN+RqG2UuAMvEhGEDneKK/lX+BerzwoY39t2ViHR92iP1W9zIMGZOu/G
Jdl4IXpDtHK6s7BRmeJaoqIlZganz2m+1SZlBpoJIXV6C11KhgzDP2UM4AMr9Lso
q9H/VhP/frZFRS1IhrC7YofRqOsYuI11I1CHp/KATg4FXGU5tGDJb3khp3zHDlPk
a5yTFnqf6bGIrF3pGXmz8nYLtojQzfu4nSu58RHntXTC7ULwssB90tZN7Nrp9Pwl
dbw3+StefElBy02JMNg3mMyP0BHZmMv7pvg1D6nN4mDroKx09u/gVdZKVlFzXtxf
K4HiL7W5MewmbYCUjT/HuMY1/Jdf9EnEWHDnX+GOom/9Ps6yvSbxM++8OrV1yzvs
FuRksj8rINLi2ffbtXDlEAcHlA8WFAyIuErexgoreeVDSRjjHTc5CvAJZ06pP3sz
YJkkUHT7ysJl0nWD4rt6neM6fObZXuXzvhF70NxdsQ8xkMlGVToBAMOitREArygX
92bspNGkcQV/8lyPbSEMu0e+1Om17J5xJDLS9vtjIu+tW2R8r+bO2DfJ423N9sD0
qKnKjYwaFNUreoSznaoF8fWHm4E8kblL4Mq7B1wOLefZbc7ATnkxwbOsGtqs6DB2
KbnvN30ZkkrFdiU2Z6JrIp7d9k4cCPVvWdZwQ3CeMZXfXPhwL6HpdoCjkNNCvoe5
ocrgTkoUTFCJw0uDYbiGXpFyRkqtgTaTWdU6txt4rFcZm6NXqxmt56KAgLS7srvS
ecQjcLEXIoOIJE5Mu1knLSMQ8dX1pNoqScJG6+qT+xWaboFmGxToQs7snlRzJbMM
wkK6d6ouqIM5kopvqRQfiralT9qU+GYQoZCuuOQE2+U0rSrYYrrFx1A1vJRmtmaM
axgkzhjxjIA/M/e65GDHQk9ZkhDiMVO0rA6JJEer/dFTUhbSY5dhmFqvaEbwF3Fr
QmBz8thqwuDxuzirS++AugMHdIDsZXWhAUVX7XRiXKUe7I7GBEK3uydUsm+quy3S
GNxHqJnRguHBq+3ZZntBp7EiV9erziLtvtfp8zKaTbdIx57pMvfN1at3HiY0fVRR
eZXjbzFyIuI8WMu2IX6TWqDL11eAG7EC/OIoQzc6/o1CgYcKjfKCxT3D2XWbB6Wj
TrEabNlRxenGSnQmz89zil59TJOw+3B9NVI95fyjeiyBDW36jp7rS3lcJcJsY9EM
oScH/t3/1d9IPu1d++NgVMS5Z9qga8ooeL7eL/tTpAD3t/8Ahs1+zEeTwV6uQGdk
GjrEqt0VjbTe9h0NA9vA8SfNW0YnGmuZNlu/faOGfltURkl9WsiUhBHgOOV3gR82
EAWhmbgGIYtag2lfQyeACMQ0SjtDE0ilSQqKgvFyTL0a2ZWaJg5piHJrRNvFyQCA
B/2xFAHAwsSURajTJkfUsY6zJcRSSsTn5hvtlBj6AmxQPA0gNygZtYAllES9ijqR
rptz9edNEKHszNeWElpcYjRScUoMCx7iEjiMVpdgDtJm8l2yFvfKdWJWkdnFNF+9
dRFnmSKvxXs3WvjP34BKgMsUcZSMjnyJa1leaIVXofv2AtSNthl+KRfSDFHj4ZUe
8jW4KWR/mYjuDpTOlXm1a1Vk3KesDjVNLOdX2yNRZ2JGPlVG/vzVgrUOcxo3lpxG
YLINu7KjQHwWFfq3eVbye8E7+XcwZE9apm6DNMnrztlRmOtiGPUxGvaSOzWTXViq
o6KYlxqdVNyOnJfp4jHdvDn1lGn/B5LFZVukugr6yjZ9P8l750OT9oEcRhTLhDHp
gdUd1GsHYjiL9enaOrIBeH2URZrh8wjFdEduzjZzGhqnKi9qYpATkGZ1SeXYfs75
+EVYdZ9LPljZvhOtGwtcJFpuddpao2CRdaUH0COzabDhObPpZ4QbX1XfIMD5Ga37
fOhnJIcGqVqPF5MwFFkz2kXHHIN2t6WS1j2cY8LJXxWuF8iDFlnXd9yxwskDGRBz
5hS9TxbsOKWI+hvArm0+QlPJXeYp/Btj9DLzhDBCh4rrpPE7mXeKIFL+Yrbmlk5l
9LcMHrjR3WJvQnq4eR57YQbj94tcPCiWewEZABK2fe4OCi4ivmV1MA6hQ9ytaosC
mmZG7GWwxOQ8QU4TOu7iftZAFPqOAfxKwC1EaVr+cvyvCZ2iVlddravnIpiPidLY
VaCf97ReFIBTpNEDG7f6o6nHdCUozxyf8O6nXQvY3ZfuCVuqkAj3ChHHeHg1iyf4
lpXfjoCY4PgEsCRTEYnpEvWqOOuKFpcxG3T8c79nA+HVcPnKqnNaqq2XkVWS7IM6
zyVGc4Eu7ee8XZ0l4DOtEHbAxdMniro1PtxTsBrD693In5dmyZuE/hBuWG2QofWP
SdbY8lhHlEyC4o5lC9rIIowNP7BiiYFL4bluch5H8Q2tVhmjce0zCKTOuaFozxU5
dfCSJPraBtIlOluFirxwbCqWzQmbiC4MCZu2rHtrBwwXZ7zOEB8/Mo7gxJHKLz8M
2ph/4nW3/HB8hSmKa9Byl3kvO7L9rPnx0M+vMA5sohhmhJAvK1qKque1mYB3r44q
BvqDcOmY/No36pWQ+DSnEC3I96qbdOkNBTgssNa7BMYqyspNWv8BY3LTo0MLLe8Z
StvSg+jfGQWCe9d1Za1pEJYtdNIC2fjBYb4Xx69rqZIrb8CR15lriV3hxaE8i25U
33z/zhkVp4AIpefkYiIADOOzcShnRNPmSFaUTBVMxMcPHPV9T4GFnvhvdkAyDXxh
ZDSnB0VpVaqequThdcL/fuYPEtFM+RruiRurI41j0J+cXMLxu4GzJWZjDVWBbodE
zNqy1WwZziTqqwBA/8hXx5WLDeJwI07VRGi6Q1MvDjxYsUX2mbuYR8SkU+j/7oZU
WuG3SmywLxJ6UneqpV+qDbgRGSc6fUyw5eOzo/fmw2tgXQUwoXhxrqXdJ5FjiJxB
Zdvr0cJFLaRvBc7LjIhK4vaQUEWfokWVts7+ElykGLgl9DfIkqL+bUcQ5IU9P9W7
8HmUeF2fibIa52nrbm1p+rzfO/RBi8D12krL9Ix5m+iD+NfSi1L0qUkj5JCOFA0b
fvyLsCdMRu+P/0icD5WRptUauyR1xfgk8b99PrSFDHakOaUvlbbx2r3VBhLHbFpJ
5ByOq2WZjlvoovdETGRIS9GNaHIKMQmboDXU18D3/BhPwXjVYdSebxKjZIAkGHwC
AnLmdOSvvF5Gh8E1wHD2Iw5+Ct7IfZyhHXwGmTeci7QT29CVSqlS2DujLUzGaneT
CY+NIf+lmqAmnW0FXIU2mIft14t3ZwrqoN0TZxjxZV+ReNG4KZZ5ynV61Y5qOxFZ
0cxKilmklWKfFbqpVWt8xBPTaflUe6siWMBXXJdNQZ4n5PAoNQLcbfGj/Kue+nFQ
IySf6p3EHbB8PgffjOS5EOXy0xH9SZXM5XsYiFLcMsv3S4cgAvgLbksF/sD2MWvV
CCuFib+5KXic30zxfHVjZS9+fX6wFf2kjC3Lt3nzQDK2vZT5jyIgM4QScbnfoTZf
Ba+m4xe9UQB3/4mA7cglu5vqF9j2/nSJf4fdqR7kaEKz0zIZ26iplP1OCuXK8k7b
IK+YVXsbbXykkO1kYICLCzuNtyI8VflEG9+fQ7etsUmECHoUcyxM7CvKUEp7aPqa
UcsUI4WKztMOC2NlB84R966sImvAaeMAc3XcFpaqJWOSnYFUhlizmSzhAn8SlXqx
z4zzCQ2iBhL6g3EjimiWAhS6LxOOKb5MDlfQTCHlYWf1jrvoqgjJMbiseeWg/YdG
ZS8OuRZK+x4p5OcVmMYtWi158l8tj89VJhAldU55dShst9WxhqcedOAZt+021u5c
vLnhRmLKU2rm1KOnPNSKJ21/l2UdRF6vwM5ekCXkVbkzs6/noHSrPgsql1mxbpZ8
9171zg5B3R+vR8+JaLBSR3Dchz8950NWwzI3H2IKdE4R4MlkUe4bpQynlXT0Pu78
+IqTfLdc0QEsANgNoU9WiCrV9qXgOcWy1+UKSKPRtf/z5DqrnFIuA78ei2pQOzlA
5xFKbjMKxdlVIqpPx6Nesi8qSIju1FGkpyalTcDmeA5wbtj8r0/ziIjc09Db6p9e
NuFhsq3ZEp0+B2k3ulQWb8kKdvEr9dMErsaIo3ifi+R4Olcp9FVVeB3rSRYVo8UP
IQ1RRaui4HVnz74dlkZbwcgn0iIZHtWXFFIxA3y2BohX5mt9qGXiHKx6hKUnRyQx
elthpH7TriHqQvQ8f3iXQjr+JDyBqyrLn5qzHGdjGvd1VmqmRiQPQCTptUCP0uBQ
63eFAg9xz120SRkLGYSdqmhHtewFbrHqWz4HZ5PScM1Gd7mJy18JzXDf2HcsfDhn
FNeo/SBR/BgIm3bMELCNlej2mDxj+1OrkDa8DpXBtcVjlBIXrKI4WMSZtJ0kTjxp
duZ3g94zf/a4YvRmERhXApx3BmUXxpOYe2fI1B1GipxF2H+iYVYaP8+XEj5Xpk26
GryN9gtHHMKJLfzvqpKyYY87Xqy3tjLby5yHEYW8Vi9Qs1d6eiLYKrcE6JgrGImu
Mq1w/dzy4Glf0q7seGQLg9V2S23Na9GixjOJxQ69U5z0ECn9+tFj5uJ9BoVQN2vy
AS/ff0ZSQX2GlMICS9DJG+rSykAF3y1tXCleY80O9d4fbf4I5qYBn0UUKwv5CR7n
m+FrqUJnLGXobuVs/jJLZHxGQh4eIx/K2XIaoWkeIETr3oY02HxTUFIPqC6xtKQZ
I23tNPQojLTzytNG+isD3FXJ/y+pqXzoiJCjbiF5Xd2I+GoulbaVIWGcUi2L4hjm
ssLpqj1ypnptj8lBAwfI4yVETtZGwhSDPQPk5cyuXmSymnyH6isBKh33YEICk0WL
JGTyFX5q6qGZhnxT0j4KdIo0uP5tiP9/hXcHkeRMYW7eg4JDcgXGZ2vzZbYx2LHc
BWhjz8OHlSKZKZabqL9FeMmM/qPez2ZR/6h1aSz9zXYl2ZAXsgPSeE6eqKfe9rOm
svsKvtlDdjCLf50pQ3dy2+50na3q3RWoVTcN9ktf5yQh1j5GhvCZwk0TNJonNUGd
4MDUgR0JzXbC1I0YLdUgjPCgB/uuLIW20rxa/3gBd0ycfhy6G8N2JkolSZARQJNN
2ym2SZIU3FKxU+rdIJuEf+Xp8uhjlLHG4LqEFfHN0UC1jHe6nUHZdmkpDeuYs36a
7++qClYMk8xKE+qgxsCqB9+6KNPssNfHpGyUpGtenRE2kCTmZHjfos6GdlT0aNyc
llNMlRLtLRMFuAe0zVj3H/76aDwawx+x7LikuXyp7PTOOWc5g5bWmtkyN5s00aLX
XnygAEoUhIaniVzMzLBJWMyqvaulpHcqS8rc7XyQHkeVUNGRNcaojO3fPTwWkK9D
vkmS0BwamWoMsdmeuVx8eRvaLg4ai0LBXoWI9woDUTUF41zCQDWrD8KkST1Lz5Jq
We13Edagrg65krt3+y5bonrxszWLT+oSPj9VAkMZzphI53z7T/NqRhVcdICR/FDQ
eBDDTZ6XfdJfBVxXd0UG4KPiolv717XPIJQhQOK5wYcnuYG8Yr2RWUo3sjujz8GT
pKX9O20QuGNAG2ZYI2UvKMVjb60PUBFsANCP2tiqpCwjAow7ZjbJQvSKFHY2n+0g
SDFAbP6ZWEc6AnkyGv7WJ0hN/SsVgpAD4SDSS9qd3gFYiwQmb2luFm7+R82f+oQK
gvpqJrHXqFkUslbtwqsgMBoJuQ2Dg9E8pUOBQxRAWRxmfrfsw5se0TF1NhsQgIzu
HbZFmmU15ugUCJpcL+LLThp0XOx/LuqHuBtkoum7tkOZX2RqU2E4+zr/b1fazYE3
Neb1xlITS/cTXXSU68pwTOCtngGm/WBkWOmLKgM+e6+zJHwrUTJae9MPyM7w7Gx5
qwVXTuc1BQi4dJ/nu8+0spL53uF+eGzWRaj0K/4kOAWv8sfzt+UyAa4tH9BP68rT
8vWPrE1FOUGYHve2d19gBi0xQrbrZVzip5lyrqUd2lUfSD0/obw6Jiu4DW8xpZBJ
lWnYlfXDdAm5AvAaDCEasAc/7z9gV+D+r3MEutKIqbi/XlOm/rlJOx9xLZ+3ksRw
tlOqV03wt4OcJxfNYwnUKZixRdV5KGA4X/jZcN/l/b6SQFryfUlSNbotWAeXSRwp
HiC0LdlUvAqe8UozghGjTzSMR7qYn2LXkKS58JKRd9+FYuSLPMVClVWgh8yGSdw7
WmTvAKRh3WQkK8oZ8G1dzFZ0RHo7JjL98cqBiXiATs+THFgqooNP3HC2ePXYGIIP
5tYvEU+fVhIIEFBjI/leZonHLF3Si4hro28vUzFUEzGbcz7sTR/R+26FY8zeuEk4
BEeBjXyNxj8cRu2GDRYmjuF7qlJgmQuOB3Be16PNILjvR84nMt4azRn7cdt30kDg
v7xHEn2hRNXSbmCwmZMfgucuCPGPhAhKeKr1EI/e3TRrZMYc/hSGYvy/pFEZnx4V
ofUN1vP8Z8M/7pX8YQe/gQ3jXK6Flp0mY0R9bmg+JcaQcMsQYNhrFEf8DnqbroOQ
gEkhdIPLdW9cjy9slIk7QzQJxkNYakePujIuKc2nhrCiPrXJO+BYBhViTz4RGQmx
hCFRXZeieXX/DdEGKCDrQ+CrCx3/nVUWgvyJXKXv0sJ/cmZ77xdvMMpL71ceUe7/
bGikRRWQkkYYnzGARv3ZZdjqHFYqIrK/XrjfXkbd7DyGxl8yksYIMMuzZd6IoxXz
HWJxSc71X2f/CrXBJpVit8cTsjggLvLfbqBfX6ixxaLoXdKH8ejlfyJlM9EVJfw6
eqPp7KPTxDrql1Je7Nlh7KsoboNCQwHVnOtILk1c+baeH9ISgIChbSeGUjSCPvcn
`protect END_PROTECTED
