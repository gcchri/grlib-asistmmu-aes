`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9J/7jjyrDWpzMBSZRtyweYDTcjZ0ReV5DFu9Ygk8K4AGQCzTd2WC7Q4WjnQze8kl
sHRaaZyAx4tHgFDUllbqN/pbzxb7ReiYHM7eomVfADNvZKspShS4rGHVTqukzpWB
RezfBmulvFq4TvpixI/xPLerPg666ealoQpWsVJXxVGZxd1tRh9GrFrKVM8JW87P
KhNLs4M9bv31bqj+aXh6PUqEPc5fNR0oV0cw+Icn9ASxCQM5zF59I02/r/I04kzV
B6Q9W8gMX6nRnrTdPWy8DASns9K1BT9dn9WMo0AUdr+U+IaYwRrfMUQxs+EWEWoV
eEh5yv+Vp1Gqsm4AbMp9Q2kCFKIW4HntVY0tjUeaAXJCUIYvXgEv39hnSdSRDx0D
Ye09rO66P3V3s6wUJL8LNOM96VXHxGjeoB7pDCYb6lM=
`protect END_PROTECTED
