`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LpW1rwK774XPr3UPd5Y3ZsdLaZuZYpvSHD6WsYg8Ym0wKcJlTBw7Y6FO95rhJsOz
Oq65vxtSMr4BPfi1HAYAUUHA62G/DsAAJQGxMJtIbeax5/HzPLExuV8Xt1FfsUum
j9VzoDH6AjS8dqXaGCMIPVS/7aoGUpBokADEe7S5sNMTrCHGjRDaPOzdN4wbg1SX
alJVSkQsx1lAEg6vR4iA0caiOH9FFjfAZlATp2Y1vlqlV00cJPufDOI9B+CVAgr0
hkFt0oWbJ7AHIKgKwYIrkjDZUCLmeahg+ooQmgH3stF7gjDFP2cux0sm7VrdKVXf
Bjfu14YWyp/XMVknkWeKeCyOYCfVlPMPdNicgjgkfyxJGeFYlH2XqyDFqhhk1uTo
eDCcZIuxQogqZPCUauYlqBrh2NVt8U/had+hCpolXuKamI7HAkhMj1Wq3NZShQpA
6vKi5mGywfzqA/goZXtaVN4tDr6ROYbLHacg/3wgtnd6EeODh+KKHzCV00aS4obf
9BouKi6lfAf9o9IWMAdChnyDPlCx/AImYExHESuqpubLA1+7c3nysRY8+mpwe4rA
p0pANL4CZ4PuQJAam6/z/97yOgnyPaoFrKEAZHtVcp8TLgT/8baLAMNwp5fIjyeL
lfMjwEpD3RxS2zIUrAn8/Hjt3omXPtW7NbzkWsVugkS1z9mW3R9swITs3YWq+3qe
JBg3O3vQ6BrewhJig5yiraEoOmjeY9/UXXynHQlonmDqCkPLP5xOiKu/jltjqOt1
7i6r+Z+VtXoc+t8aJpUZA0PaYGwfCjkL+6dHjnZy+UkvxxcTjIKwXYVVKgoYHhfq
2QM7fTbE2KBaDnm6bQhjBYoUKRGl7fpHWDJJazctcefZk6cEZb2Sa8r3h3Rx+j71
pbkqLfz7XemC9QSjCfcoXuf0Pn/BUZMzr2sIRVpx99Wx4/E8fr7/Vn7YGcmknhFw
+jVMwH2YCfRDFpJw4gt8s+SNjM91TjnSjXqhItMf1Wg6oqk7jAyOYZAOWrNf2gCn
xQa1R39KzXFvOc7AL/qO9BduofHstGCGH0KXIVShlaOtWEhiKRfN7RghC24IU3of
ZmM1M0Kz0+1AIXwXSx/mnilSlBRkFFE726JIKQopoII=
`protect END_PROTECTED
