`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4ksvraQVrZAxEy4CV57Y4QLEYS3ZTO2CxABxwfwtKKgS4CVpS7b/CIbPAqyBXFYH
vXsRUvtd7e+fYXZdDMmhsxz68kBd2fufpJhVpJU29XW2rVcxJ+s4t3aH4rRncZ0Y
Gg8pOwGap+kbD8aZ3cTS0OKZccsQGVgfrNNDpM207wbvYE5ddL78nZRIC3e5QGxe
y7MREFGadDZaI5WYkvrTs7YEHh6PRTpvZhQns9ceJnR1FHGbENtVfWJgpHB7mU87
wXOmdDauyhq+9jdkb6YskWjs6JvZbyXoFuSVMweyzSlvq/GeBaGfceGhUBe/zJ3O
NIl1t4QhvXgqbvmknbeRuk9oy01ug4xjiUUQpH0ja4meokvXMvZmM5LYwHtG+J33
BEe3kBOziGjwLMp5fMzvORINK0v/xGDk5LmzUX3446h/YAS9M/+ntkgcvzliqD1x
Fn4Vc8ipM2lP9ZgVn+Ynkw==
`protect END_PROTECTED
