`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zTA0YWPTqCgVnDh2d/h+jQ9gMT/0FgAx7LzM/TuavxLNrnae0eiN9aF8dTQlifhC
pJCgzYlyHoWY4SAwgVE5w5jg0C+kZKh3FIzGrgMMLDda78Z260ISM9cCivEtS118
ET8HakybRxsWi/YdSDmT5d+hl8YE10NKrLJ7ZUVOE3s8OlcE0o245RTR/YFIZIX+
AypZXiqEEJhoOtgbgByQneh6ywljjOCJEiwA9P2/JF6LXljM4zq/QU/SUtFBQEQb
bJHUbFz1yrFFZq3ebmbZ3g5NLAw9ZVpMACKNjgRjzNY=
`protect END_PROTECTED
