`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LdNzA7j99lWZJ3MRsOeBxWvU6B4khtexuDHl8A03nNLZjSFhcI9tDi+U7dIRTnaP
Hs+dse8CMJQbu/ku6kWFxqFnJZVc/vsIQibJU2Woq17e5Y4VjzjBqF/NAcAh1IMT
B13M5Xpi4Td1LGrLYV6EUAcHn74/Fqp5CsieK9gnQwbcs1d8bx82QyTFB/mGqmeq
6VBOMcuLvyDiKwSDQvXdgFqNMORVOHLuTHtvkGR31uMGdJuRi0YRS5053tzjdO+b
13CeEUuZ84NvW3va4ygUgWA3gVDWIabIxJihINA/zBfzTQabo6IPsO/NTKMnB6Zf
Pp+eDfbW9hx70JiQKP5EDKtD1pTtZaLGHOdCI19Y7XYzUNbLyLdZZQ51AXtSWaED
yrNZ4dwT4JyiDhBvKZp3pi2ohwIO84MBLZ2swQ0zsOoiuy9Yh+z+YorVOqWfiJAr
KkKuf1Z7XOtyg3oAPSL9WH4b7+O+sFoPgQT042CG9NOQPhb5Mh8TXFzlr0Dy0OGK
klYdvaJFoC4Jv8AQ4Ueb88woUNXl5hoU5uhGzvySu4RCbljnf3+mNib1oI3Hs0az
KdRmDvGhZUilNzH3gw0Joro3urf3/SHJFrSj+DMHJq0trDmlYPwOUSjJGitoBkg5
VzXZ1v8FyO6VDS+S/BsWlhHE1NP0bPdqzABcz8O1HUFZcY+ssp/mzFABVlkzark/
mHfoiTcLKsYWBa1/L09KOPJ9uziD2lf7u/NuOsvE6CW3Wov3wUD+bWIbYhhokfHF
SSSb/eH1HB2gfrvYRjImQO22oQE5XYuhQDsYsOLkLRYq06S/CeTpMMftr59DNo/9
Ka8cYGvYbKYXF7/mHpaO6BMiSFU1mznueVg2lVoyQI1sBEE/vwLN0t3+x9NXwZaY
cYkI12I3KaPcHF13eO3XWgeXZmwo6hiBOP5Ihh+3trwkfAqQ4eUnUsw3aLuWxz1R
jLY+AjDmDt2KtyaFgkLrZQt2KlJ09KubYiLO/6TSkNNTsWoP6bi9YlYV0nPDtYzS
b97UDMZd/9zJLg89IhPgZuC1vf1EtFovwf809EpwsYy4FKpkuH92zwIDdZyS87eD
ZFOHeauVqGNogcwYVjJv2X0nuPNTLCgZay1HWcH08cG8p8jNCtrJBiTJynt46Rbv
i//mQIS95gWjWiV60UbTSKOVRCIcyIasRHaz6csHvV2RY6g0vMg8Fi3ZiBSViIlg
pGn5x9U8W3OQHusAvUxqlcCDc6RVIopG+MZyswwFbfhuHRPM+PRY25lgoxeH1FfY
QJeP7uiSLtoM+IUVFpI+NEgKuht5WDg9JP4OOsx05jkQCp21WSwEpPGhUCLOqLaa
ZlqzDdSEmZXueUAi0JaZ2O6x83OwTRuERH+yPE3rNaOGOTJYkBR6/NRMGWSF9cn5
XPylx+iKQCh+59Nmkg42tofhqZRw488QeRZk6eervL9zXTmziG9W23pZHq5s/0Zd
0bOQQ5CvJs4ccFqLdA+YbeqQTCSdYGpRw+D9naPW9bs5aSgxwItrat2figFyiCQw
pFoOjS1Tbs4ocKOu9v8mV3hRJ4uYezw0eTyuM5lwuy/MgOYQZqaV7tbwOAehphEK
Wnznq+gK7Vmya3RxzxRaRTCB65bT1GHse5xGQ7HayASEmadRZM5sU0OtoNdvHfNq
qWEk/Wdh5j8R5BZfRAQvCGA6qQxbYApIJz11AB+Eu7hcrnh2NpdxGHvg9/yAbsq/
EHdtW9lWVx6hv1nIIMzYYP+d3qyqh8LNkEU5/ZD5ybE6QRl2ZgXp9GnAJLMVHK65
JqUlkeAR3V5rbFdbOVrwbQ==
`protect END_PROTECTED
