`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tIlQcGCbuYSQHL6/u1lMm7Yf3n0G6zcbRWIYpLuPvTYbMfrZUp1pnHBD+Qe3z+Hd
/IHUEuOl17na3hu07RdKV3uiK5VmXfUonZkj3Tsd5V1WqIbwTyPZA0YC0TIrIC/A
EDHEK/MlnC9kfwzWaeANk2X+hpNVpgKruZ50kP0l6GZ8nwfm+BdGYf9jOvqBYMsx
07mozRE8pTOOtefletd9BxXN7j4SHwKwrF7NavkWuY/ttXlo2ukRIq81NWt8Vj3R
V+eTCwpeSNtkyJ6fcrjpblUIBIBvcN7BF6yl2Wz/bNvi+QbaYhA9gNDixVNq43aO
S7wg7ZTLcl4jS04AXe4uwkXmO+VvW5lC0ekSlc8CcgWUacTUCfC+lodJpkuKdM/5
MYesTfyjF4cNkfUnoQapD77O1n0CdtblxTjIWuhTTcI/xcVJ7CEgGDDzHAK74l3K
Ltw9IUNHLLAJ/K+9InMAFaGadCLMvGBpi0yYXqgXlPNobCFKXzt/ap/U8SapCf9/
rAAgQJ954b8us9rND+JsC6N8sQSI5sU1HSFW1uwJut368pdI2svWVI5FbWUOMFif
ZbVPbtiwagti/NEG/MHCRr6c2n7UdL5dfSJJIJDjh+14sS8ArhcUbzkrYkotEC4A
iZWbSlTvrRwEUimVdJmEKx30sF4NFUSiye+verx1GOpSURVu4NMOoe3tKLrWTzRT
Ogdw/ElYIp1LF7RvzHWF/1a9diRJSKQJk9zkhAzZxIu8Dh1iHI2AyccTVhpjbaR0
jBTgEqT+MEJlukiwrnw8cRI5X8dfVpsfSzWDWdbiwMOTKIWW1bIecCqHTnC8Vj9X
hN/aB+0+kZlZMj7gcVShePOVmfp5HrYG2Gqn5yXfg1sZwwIcTl7Q5ouZUirNFlsI
77R+XV/wO99Z2MLD7MOMd6Hi/H9CbwSJOeggLSGGFb0vaD5gtkGdaoWQE/IUXYwR
`protect END_PROTECTED
