`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
06bTAeI9++ABhkKdy76dKGqYhbR1mQj02m3KrprdXbU8QaRjn0cMYMIYqePiqzF3
XUBUofns4lWv1TevqeFSZvSCLh4iILFANQONauNxCtpPlLaAGLL8cVpMs/JKQQfe
lfGdYDmr+JJf5zvOvUjEJxN2ntE9PTBcfRSv030vicBvxXBCSd7bYi7QZQy5YIo/
Futn/k+0rajxSYUFZL6n/QKySkO1vOKtQw89rw0EdaCWXGW9Ve8oRI70f1se0X8r
AWBuIkuWQSQ+HTuMD657GKuR4SGqusTIeP0s/jhXJgqr7TpHChkRpgmv+8jzYP5M
8WXjwh2iCZWFJh75lAatnrIFFsUcvZosE6S6fd1ezaa212KHwjAAf5XQlE4E6Da1
+kLv5oGvlWm63B5RSR1yLbMfuV5SuYRY/QZLaQQGv2+VOZea74zetY2DBXv0jAdL
avpWs7k07A3uWs2mKXNyHOEfAZWz26N3OR76b9yWtzjddUxKzPHvJUe364tkiSpj
mfhZ5LSNMJYuNj9OdBnSL5AtPeGDEfX3SxRzVbKALMCIca0pKlhHlWKbvDwde76h
yFM9Es2//L9m02PFJNm02NhsNuVvs5NPx37URYyFvksk3aaeOCPUHrqZnACcInQ+
EGQgdxNfxdhkT0EF6VZcWXFnwWl6pyCq1KzZIrAOUMa/L1s5lda4sv0wdNyWBbZ0
m71qWrp3irf2bO2Bij21eb48XUbxNngbo6SgcI47Zmh2/SdZtH0GKW4MjAVUSZL2
GqrT/Dg/jHVLSOpnBkVN42nJAagIo1P3C9r6kqgzyYfDM7M8QC+jTXAA3Mg4VOA3
Yei1Na6/gKciMTzAHsK4R/aFKy0SJ9fMThZ1kXe4LQMgO/bBaDFM4gzp/G2NGTWh
y2Z8QbBuvgPAiKOQ/PMzoEQ1tAAJi3jSJdqq/nxurfP/gMLkdhcmdXf0heZKBn4C
HWN9QiZ3QgOfVHLJqym6B7gbdnGyD8xsE4f/VWrl1WCX+T30gplfKlkaVpEqQJvr
qCXMjt16rE79nWrgmn9irE2FxSRDcrF9hVMX1FELEWgrgmzVPjyxMeoMJJXOT0u8
uajy6Q+SABGcOOFix0fab6757f0P65urmjfRJQGc26O272LapPoBmrsiokV9KDSE
Tv/rCKCqIQ8HvaqSt3c8AVR93dvfGNYYHHT5SGEPIYYrgWifIaQgipvo55hjEgMj
ZgFM1RyZFULe2p0JtPByo9zDIFNsyJlVaW8m8B2dVoHqPfNRau7EUDoyaQ2ANwMT
5jhrANB/gxu7hnNcCbJ2qgyNfF00uWleBe0bdwf6a3ZMFz0ntejPMzwwfnl0WPDl
Ug8DU8ObnFtUge0ueauZ20R5jmOt8Hgjah/vNqCAd2MUX65WZh9+i4nDCzYBuZ5D
G41VZ5Ue3qumqKLbBr7LQM9rnIzbtwers5j/rkIvFQYJSUZs11rwtdDwEJ8yuGI3
TfNO/1TCJxN2P9E/QdNJyBSNr4K4frGBeb2iRe2/U06v5ikHP1zInvMMiGj0Th6x
ZP49/y6CtqRBWgVwuoopzRJ1Du5rvm0g0cq8R+GeBXXKjyN7W6WoU8exSOr8YPwb
bkMDy12HO8WWJU68p9leOwVSdlU6I3LkMoYEueAawi+xR2qLTo6NzQxPME+3KgmI
XDQIUv5QjGDbaX0RQLGjL+X8GGrlqP0zGRwNmGUpKQNfh7BMiG9vGrJNHFPOd3kM
paQ4g1n2+UMY9dpk2BB9i4lPsua13MfAKCD2BTPGswLEdkiPB1sFi/GIYD1XtD4l
dyKyx+PKi2aqbmFHKob652inri6TqD3qhG7KWTwTJrZYdfp8lhPjoPrzWXYQ4lb0
2khf6WxXgqrx9VgjXVtVzkG8i0MEQMZKuCEBh9VUiJhXK+1EYzWQoF3bINGADkTG
4ePhEbwsRAd/94XoxEiLv9e2G5rsHJb1B//Eygji76ESKQXJv3o39xxSCz9ozVsY
gIo1oI00/vhaSYdrkwnPyrua7MmuG+yAr+BuHxqvjOe5QnMnZTQ4bem0MqwY4ZHX
UlknX/ukYXKaEJba0mZpGtoX9aRU5esiZO6qK808AIp1ByVGa0bn83eUjdt05HNX
lx0C7i0GBMZ0e07MyzRz/3NQGlP+nobFrGWTz3o0GP5lVcNcSrHkRGIgITaSBqyK
kX4iStPUY56/PvBAPaqlMCBuaSvXYuo6Edv/yN/jBSIzuzlA74QeGJiS8E51tVAJ
U9XjNRcXuhWzIqfE5ELtgAyxxYUw4AXwgIn32m8BtQXYWFrIHrvhgDJH86FMg4L/
x5h2uqhijLVNCFc/nN1LPEsPFHw/gqE0moX+BqQt4bXLcXqhHNBb08A82M/AuTTk
pvPg2dzps1RSZemJxCK6AII0WLQNG/OWz95PkOTwm0Vxh2sVSD/FXEMb5skX3wX8
Y9sFLFFHevxvObcqk+9MISG28Qr9ZvedGRx5jM5s9iQlMQbKcIqdzbIGGH2RBKCQ
3o4PIcCUU3xGk7DaXSBvrPtPL+RvMgJw2cMvp6qp58pm71jxH8VLg3mB4Kx6QJqN
ud2cVhqTvvL3EMK0DMNXZthTzfQt1RYhtbDNxWOvmbrlA/mgF4QcNIOQlAK6CIxp
npXkKa7SnO21FsGBiIiMGCqHsrJum0J4uJg0XNotudBK+OWTUI26HvidbzfDRVq7
b39SWeJeP6FwTAx/MgO0YEASdYaxoko1arwJgIFvfqPyk6gSWMxS85HUNh3DaVWk
F7FXorHTOPeg/UcRFhoaYo8hoNzJ/2Vsco4M6E5QIy/eBfl2q1sQhpzsMx/yG90b
FnR2A7nxeW1O08XJ5ZocQc6nfrJx9h+QFAyPQOjSvqPKB79mCLarrJ9FHrKImeoE
WwzclWHzY92NqeMEK6IjiPvw0zfoYMwPRe1pFwPP9FCeLODB/jnqFuFkQocXPN1c
dQ2t0uNHOsJCDiHtnDULace3BNiA+52p8fUz+CeeJFyk4wDH67k8LEh4yULICjAx
MEO/RXwK5ENvs3l8x3flOhAl5jubf70meAVSpvrLy4iiMBK8IEV3utM6oxY08gKi
yY4/wK5m9McqmnHFPwE3PBtWldgrhw6HhGjmcb2VcbIyulfM0Xak/2mrVyHUx6O7
NRa2YnpLzguDIKUxUSy41Jmj9NNQmNGZt0dwkmah0xLVDPCz/f3xf+kVTLP1noxE
IKSy3u1SDpbQdXzsCWvB7lTToaCQ0FT9gGaKMcU+jt/w0qZLTBj4r6jzc4XWkPWK
PumQg61FWja6YjT1X94/umnNopOmRc1NqQVQufntFQ6e4S5wtq5XSAggPh36C2tE
QetdI3Sn03u47T1HfDS1pWc3XpA5M3+1DHkUlxi5lFFru/euh79oqLfrPHIOTtG7
KKowreRyJEr7hWZWEW1/8TrhTz+LyBmJfM/PVOhjVob0qsOWNBKY2XUZFq82TMSi
U6WV7ZNQPxuWqJ0N6Lg+gxnKui2peEY1/f0Z3ljzP0MC9AfcoCaZ4/E640faDEgT
LFj0Zyo/fju3Ga+os9Ma1ocOGZt3X4rY6mKcc+EDV0lP+KRCnHR4ZXm0YaTZUfY3
0+pS6P9IFgcojd1b+ndGaR5/6TRGqkVi/yKO/ucOJjz9wVuidIpNnVwSejkIc8BY
cnezYNby5HdbIIGtyT3QfOVw6SZbx9vkKD8AA8Vam6rBIXFR2fNcdtLdpuzigKW6
bVrRa8aRk396jakAcKOUkDi2k3q0+1Kk7smx84objRPEGbBM6spK3ySEp4JC7lkN
cNQHRgcga25wite6HfbyiNGDZephUTzPvbEKh4S5/5Jmi9ShRBlBBAmTaaaQC4f6
OtgAvrk94V9zJ6qHpOZVz4jZGh+0M4KWPwlYnDq7GBFAOSHFNiVUgzGu8p1A2puV
+AFXDEiYcXk43JC5eSZpyEPFkFHCwF9HonjXGAyDCv8xOgnGQMl1EUHY2fbKG0Vx
4qI7lusmrsxWP59kzOgYCFziKiu+Bra+7/c4hUIpNSo0FQw5p/LRwI83IxCnNezv
Gu5J28dNeK/+zeOtRbARHOwv0xkXxzGuuMJlUSzTYw/0KGhgk6FTxh7rw2I7kQBl
WfuMBrXmRP+OEttaZSTsS0i1Hg0perJ/ZwnjgFCrsr30a5kB/qfUe4OpTWcEI5AL
5AJwwF0kJkLOiUFsjNfr9uPKr0hCDZdhfXIvqIBcyyEvLis0bNFqRRBVm90Udsw2
pXLNYEJZX0bhhj4tpV2lxic3XnDggBkK8tnwoN1ue1wkX5AskBXAXzcgWlYALbQO
ywBDqnC4h8rrg1kRBHicmC2MUGC2WPjVGdmIWr5mgMWGw7XfQAaCTfj/kuwFvrD2
lriuWBoI+xv0FOReIeQkmW4/BC+Ct14WHnndQ6y0qoeFppCdcWls5hFYrwqq/zk1
m0oOixHU1Ob/PfRIsWX1Lpwqpye3/r0/eU+sAdZSW2w5T30nYIe7dpG2XouEAw9m
IC/AZqpSaBw/0RH9KST0z2oS1jq6/7TMSCVLON/njFgiqOcJKX1eQf6Yukv+WC/A
zPxipFkjO600B26uOkWWVgGcN8wG5J1vpjJCTWjzz1Vxmvk12SUv39S7kGSIentV
psLyV9A3UOlm3FoYnnQRxH3mEaii5HVwRtJSIKB5c8q/Tw1tQPFc/6JOuziB6MP1
jWnUCtp22n2gveh2VP2EUklSaBphoFRZAfuniLNoGSgeFzYK19RMBuWxsmQTwQNF
5wUWtUbg056hcyT69zpXepJ/x2LEuTsYCFLsCAIyC4TRIrWWTFGPbIhhw4q4kZEd
pf61asolw4S1KbrHFblFIegwydDtcpnPT0RBFtqkcrj8nDay2v5sjoX/zR+Bl024
CNau6Mn6BT6Nxy+maI0IwsI8Ixwdfunq9/H8zKQucSWVpvEI9n2jfieiyNqhiMpS
z9YB0y2WZ2osSII90mkgHBUQ76bkx/Bf9dB8+cnXwZqCEzo8FAgJIxAaSTbT9vnS
1L9Y79gztBQCo8JNMZ/js0+5NgVCwsOHz3iuSREkMONEwsswOLqk8CkJ3Ua6WTRq
3cu6z1RDNKgQhPmSFnSIXLWyObwFAumWuY+ANy3eN5CRspMo382WkmevC9l+I8wH
IcdfcPIGCT0V59HK6s2DF41x+fTry4wbJP59tdtJcvj/Unth4nOTftcdV/tdWJuU
Vz/yPA4PAy/trCpsZ/jlEqfZZUtM+fRA6FdL5BEzWXZlL95W3ItD5skvLbgDLE6R
eZeX6MbJx6mAa2e+QvIuh1d2B2vP0OHrMHYyrawe+IUrN9AqqCBBOH0eK//jkYI1
3GmOxJWOpOf95OD0BadAq2iqgtdV/G1KL+nZd4US+nXbCHthnTN59LxYnbbjI9n+
BvMZ67dSC1fQUyiPQY8rxdwYyG+MnePnIXhe8osgtw/b00jMVDWiIXFFeb2fsJS0
zwcL3L6DI6OUYvk5bz+LmTTML9VC2Yf9NhWeqXSvqghwb7umCZwN1OMK8MxG37Z7
g14wbLaIoZP9nN8w9L2Gl0iALfUEAWUhPKYHhJASaq72uxi7fy9lMdm/hiQRixul
5EotD4/RqUJhGsjIlrNruKOUGARuue9n/YGKajppO+wWCq1tDvrmPloZT3aHsWg3
10JQDO33NdcBdgAAAPE5QTcx3Vl5d7Bi3rH2szpXxaGyzdkfuC6CedlEw/KKTnbH
mJ1GVmKlmCDA0gP/qHEumHdfNWNCVICByvozJXpRx6Fu/g4zSs/l/jqI+2Y0Ve/5
41La2Ui0sbB051oM8kzA8RZhVz6ejUjRCzWmUp9yYwQ1Ch0fEl9+bpWToY0Wo12n
Z3zKvytBq7PTxufM0UP/6MfIO/gXn+XbMbQZDKKAuuNqDd+L9J0nhH7FeNcgOyEe
FHD9jMx09EQbE71dZOXba0hsHKu6lyrsYOI7paJiPaDD1kxyHQ5vXDrJjApixSn4
Z8eQ7o07GPEJLE2G8M5gnaWi0ns8sppKWA72Whbf0Vy2b7LmE6bprhOUng37crUI
6TdgkO+orSDGPUV8JPgIH47D3ryg4UpTCWhG/lsLhuIM67qV3K4AGJvh90P6jule
ieptRflYAtotkaZ5BnyH/11Sv4gQJXEoKIeGLcp/Xb84tmYcQCH7gda4rwDJHR6s
gq4SZJfjLRY0haYRfrVSjfEgxA5VaPTnc/am3nUnmzQWXgULd6/8i3c0aqjBT9tO
l9erAk3YGWi5PURyq7q9OP/CtiZjfmozEpBshBaZQZc6FBqGxOVsicwBfXOCNO3T
XxLGlzAAjFN089ek5qCO1hiXSehTGIUMNZ1j5gG509yzxhpv6Q7cPyQ3hQNwOz0y
/I3QUXiaywg1Tnt/QDaBz/USSq8h6nOwsG3+8zIZBKvtxFTf93hCgJkjrnxXcnfG
ErbfjEWjPv3DxdujBj8YaaIKhvsHvnEvKNGUWykXHGsl6VQLkKOV9XTbubPawWNc
VQXaNAJzrMo8pNWykO06BBn4RroT5loZlqCvZmQApTfuGDzveiFNuJir0v2bOd5Z
iT8pqzwV2O8EQnLL3Z+QjdjjagTtQutr0vsMSsCG5w9JZRr7+k4NXVYj/zd2k4ZE
Rjrt0tKjain/COv45SD1GaNmjwVCGWwvb06j4PQdNiwftgMYI7TzRsEdXNdj4KdW
f87BuOiI4ybIU0j3IcmI57dJ6XBJOFkAEQHUeX+BjTbzC6niP8n5l8JNcjFP6ZUM
Wk/QUTT2kj5YPUFJXsKYSVfduInyqrLb+3E1Wl9MV3q3ejodJ3JVqJYhAbrwJnP3
xo5aDmmlZFcyMzwIxsR1T5F4JZ1zqi1+pD1UPyTu/Cq8CUDtnU1usT8fZjtZaUqO
jAbDeB0JRgOmmq5JKLv06l74GP89KyLtok+9EPpCYI7L1SfmbT3HVEL7O0T3NAj5
3to3KVLdw0Nt0XhIPA8KEUagUa+sKwYt4k1JnAx7hXJz9ckBSbZtFoW2+FAcC9VC
ENNnvzBa6IIBBOZjuBYLGr/Q782rqYOFa67TdMoPqGZCUXdsiX/r3CIptye9OzJj
e7IlCaX7pNM2XlbXhWV94QILdQP82/uZzZ8n3tmZbmr7YGDtX3nmiiHm6/7D62eH
`protect END_PROTECTED
