`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YeJu0Wgj5p6OruQMmoS3OsDt1bKjOugULUW/N4qY+KbeCJbJ4nSVLqlvVMn6chZq
mDkpscuXTzXYV4VAh9YCFPd+OyFw/FuXoitDa6vmByvnIx0ercTujdS7euhH1yFZ
dpfyxt6rgpW7qHqUudttsk+XDP2fgs46YWoPbObRf8dk+MFQxNypPrQ4dmzZwEfL
rFASz3DwJ8WPSI68iEE35bFEnzOfeuGLGkWzDEv2kqkuf1DyL6FHEoFtPjS1tb4Q
JZP0pQJ92miEYW6Fdmioa1wHYZuK9h1RXSz8nAx/KraYRYIn3joFvarWwhu5o8/s
kTKDTN9YwhypTuv3+0Fcv4sK+b29wXbNPJVqcbo0UDARcIzI5zYGD7GaNdKBhV9A
6hjRR7ISDA4Gq005gTkmGk0+EIhgRDzy4gDzy6q8b78Y6mg3VAYX+A552VjoWReX
P90jxJ19UoGGZAmxkcC7O03RtMeJk0j6SsZHfLZX2tZpGhWFwuWuRaSunivTRbsf
JRBValX6KGux11x3Ri6VueyDZYIXA/vQgWLDIndTZGH+DpyCo4vY0zs1UxCJij+h
bkWrREl6iRDK7JQtzBwdFA==
`protect END_PROTECTED
