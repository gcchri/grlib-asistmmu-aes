`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c3Bh75ARVVoSXFUqwuNzenjGJ0FkAeZnfq6/WL/DgAO4iOeKCi42RsLQVpaT45h6
Ih9geny56hrbk/mUfuMojdVnT76IInkdIbHEzw2KwfoeLlmiwHqdjvjih4N09kH0
H1vsjOmXjqd3ml9BXZ69GaML5noqeiSMUllMsjiLncYIg+yPZhzyz/RrQZdnaiPJ
PATTJ9VmqVrpLPgFG5/0+bFaaffebOpXG99o6r7MF4mvlNnPzfPdyu5rWxG6eIx6
5MAOJluvqmDRFjACJyMKj9P0Td72sG3qlHHkl8YAwTzBsAwjMiyilEpwopaTN+BL
BRXcOgVez6yXSG+BkHynJjru/ugSHbhpRbkkJkpK02WxHAqBRHw96mx/KXtHbaJ8
Tcr8ojDxwPD1onnp7Hvli0lAGE25kmeNWjdki6fvEwXojrWEdHXW+PjozCJHTeIZ
0tcQpTlZWYuyE+b7agJCpEFH4jlTq5+OPGDLP0PuNhRBUEflltAc0JLvLUzGkpmS
wa2sNmvPdVMQBtWUYQiJDOmPjguW7xs8f7Z3BdPKgFvLZvdaHlRPMUnadB64ZZKI
uU0h7p8aDH3D6DqQ8vbdpXOOQWdehBf1rD86QMQjhpJWkksTsas6ImWRvgc1GZZR
f52BbeDAgIw9eJSI+04W+LKOq44iUOdPTABfuMFjHkyhgKH7PKDrFL9EtcHCYyuq
e6L6R8y8T0WS5FptpKQS34Le2fspkVeKkWkWPl251c/GDCdOELokoaIGeJrxC5VD
Qn+DIeRFqHz+I7e168bJAf0pRXKusqBBFo3s/vYVyZoElcxGDSwWj4saeM5/c/Ea
Afnq3J4E0l+PpJA2LusXuup7Fxd1jedEIc+O8UO5HWtJ9eqRVq+HFgPjq5IVE/ys
7yObtwVtWvqcN7FN/2w1M9Wq2e9dypS0g2Ec44sOUQZYBQ5QfqjdkQZ9acJ+/vhz
PyhXYcv3e3sFgHawKg0dvvY+EF127++Q6pJhub0x7EtCZgRzN8vmcBhjJpUmTcEA
uYuhl9A8vkidHIPR8qrQbFXEmc/EwTPAjdFxiSINUQExR+AFtP4Y7k+zBMYj4zMX
ZNfelu+D9+cC97eE+7Qeabp8rJYjf+a4azA1D1YhCC9QSD6tUtj36Lnc/8WTIBzO
OK7IBCONSnIS7zL3ICjzm1ke51lckkxTTho6Ukx9x+5W1pkj9pfthVZUTJbJX+gH
mLF3KNjh0INJ14aEEXOnzUP0h6+FwEPvFRE16xNs4XKK4bcQMuQ4CIastbquskXi
rQvxeVkI3yBQ2jHFKgHEQ/0DtroKZcHRrhwaj6wJI+rfVhB8MIRFCf4PYuhdBN+a
xvI7Wd2/vOnQWfReGu9FEuwayPc5nOCJjOEb7jmKuKRO79rZ1zwefZQMJK+yw7vX
dw9kgm6x3kINCLQfzEIDdkr/9z7/PfLME7yiuxvHxJimZIVnQCB8h796p9mDRVgQ
p9Unwv+T7MNHHZRXldIs8VKGE55Szn4NZoljO+oaT0Y4ClYLHobzlZN+BmuGGH1j
yEKPbSdBGk/ObbMGcwcW57BFqppZ3DVLfCX6cms8Pq+bqCR1s135zAtIBnvAHFCn
0JxaKDK7JWWhF0VlcgozMzjuWj0fjx4mdIE+R9+Xw/Xui3Gj+9hf6kP4sYYAFZC2
j3KLDliZVxuIrxUrAmM2/7Ya4QPAY3pslTdAwhVxuq8xcuMx8DS+zzHaWkHJ5yk8
LieG4R66INjCOsmy/z1UEw4ZfsvnaTRzQbFZkTIe7m2Hkn1/Hp9/223tw7luhY6g
VYoqQNHGOYdEUZwR/G5FcUBSG0K1PwiTRsgkz2NJVYtl8Pvh24bb2sEV/Z0kKa1r
FLcvHkhOVbZXwsmEqxXG8RLAuetXnBsPeGHqztRbEux4YE+OWuJFUJrjR+DQS5C/
b9QYAxdQ3ymNfnRb0PZzGO4UVJrDjt83gC8EAHWfD96JsBoDJsHnv1IVn2Wn1zUy
xFpSXXNqP3M+WrrXL9uGWgvTmpHO2e30VdMWOY5/fQl+LrKZqMEQyjmK0p3jSRFd
kjtgEqZBh8J811fmHQKz0pGKGvbqs3hnoJyJduj6zY8=
`protect END_PROTECTED
