`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tJVUXyuuv++36rIqcE1KGcPazNjfa1ZNnd2tQKbrct5z2MdyjE+EJEc91AIPNZ39
geT4+zSwDWobUXXTv4AAl/sKkWdMHgpJBEULKZKuRdGyqDmwa8sY3m0SvZVnFyLR
1SpoWpJSX3QFHmBmCEHGZ/MpbKZwHQ3KlAXJIMvCPm/CR3ZHPkQg0kFR68vTPlwF
rhRWo5XRj0wPTQlTJG1zKx3Vmu6/H4U4GWYPe6GzEwVkqpeBZS+ldPVn6s+S/hmu
EpnerN+SoUOwZmeVBGm7as6VQFxuR/tbmV5wbAd8igCQ/zRbiGBUhXkv9ZvXcntE
Z+e/ONBj7QIdh6NQJZmzpV1/O2R7ej6aah2OAIGfBx2lMmuz5cwsytTQOr7+USkj
YtDZZOpaRrSnhDtPVUW7M2rv4Ktkt5Nt5KgJfckBqEZSS3q4Evj6GQ7yPmc7bays
T71+wg+XAwazaXm0o8mB3VSEFlAZeVkoAVetQEeasOw1SGdrs6dUpidGRxYIwbQz
DQanw02sp43OmEfOuvIrpUB2+JlAQe5mBvUtteBhKUfydvMS/E1LYd2hrh5KaMWX
EqFWeK1DcGjEPEboPO0FfDnfZpfC8n6wiJ+GlQCHk8zqglPxjxWw+LyE+5E+cCIG
Ev0GMDlOUoz9Z6IPuFZFhYJU2ryl5nJLE+4Dxje3t7EoqidFnthxv4zqBZnEIC6j
F2M9mAUyG+/Mim8fLytrHg==
`protect END_PROTECTED
