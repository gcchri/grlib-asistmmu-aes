`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sns0tCw6A02uU5THHf8Ct2XZDOtnH5WV/Nnht+C4OPCsrFgl6Nn6+UT+SqCakD/P
6Qm2JT9Y22cCpxMZTta8eR0eVgVpSliAY/UFLGRwTyXah9/PQSx7ed9oLS7lR5Gd
lZZWMf0zVoEKlNQmyacTGm+IJ+37HGfNhBYROIIP/PBNwrLcJ/JEhUTpVSizzdiQ
aRKVmWq5tP2TtFFt5UrxWO1QeB3cxlaO/W38FWZ22jOAEN3oRYRHYFref65oILSn
1bpM8oXWFzV1Y99ArSqGbBxGzv76fwdEFchsH3LhCg4MflcEvl/c0YO5xC96qJRE
jHvdQYhBsCzSrWwJwBzVrA==
`protect END_PROTECTED
