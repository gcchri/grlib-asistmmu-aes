`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sut0vLqc4Sbk9x5EKLrYOqnpbnYaXQeLSxzx/8iH8HMNYYvLzcU1cBD4wGqrSTt1
4haxQuz/3SudOKee7hsWol3a7YpwZkauQxVc73hL7IlgVsQOnR7ZTo0qf3U2MfeA
kOJNeWdFXeydylROjC7Db4T7MBefqIJIcSQZe/wMyCek2OPBi9mFUhWUl5Jv5Gsb
UKxqTN2ShICn27j/JldhJo2phHaLADVAa9sz8MCpOj0O7vhc4KZeQ1X2eGXWzB5u
uJpmt+0sh95g0Y55UQ+uxO0qDupYsguXPXzjovG4N7AsLg4l1faxVLk3FfhyYZQE
KEeCa2U4ilxxDFdbdLhVK2EXSNv7VOmMQ+ESZoewpZr86EuvHiPhJUAcTbiEG0uc
+eeQ6zm4KZDzGb/TtLy3nP1S3Dw+7RVIiA2P8+wthBnKpS13MALviRcfx77HcX7/
06Y7ZOWOIM0E6s/svWct/dAAXypLdntyCQh02962ORyfyBNsU59ud8YodQiXfec9
+FPfWgWvsXwMgjEOcoc5i86lcyWL6v/iLXh8QLud5K7YRzdeUODWvXEYjswmPr9k
obNsfY7aDghjUd0QLb4c++afh0e5QaG2q9BcI1AfD1yFR8wIPmSta4NYRTtyrBa1
rA5KldnNLFjZu5X9yg1OleLkkFHkXaxncHjVHoMCCucFD98UlPiAcOCL2WDfzN47
ajpQQWUFoRveBwcHu8Ufabab5wRMVAIFyGv3dZXgcgi+iZbmbA9+v7T2WiTX7w+J
AVBkPp0Nc4X9PHh0di1N3rSczt2r5EsnrHeCf/ZI/jHIV+UgVwtTJMg+CyGV03uf
GAd9RSLyhU/og1S28hStjBAvo+nI3GZXpUnvCRfxDWWUHPkOtj+GXDfkAy1Zq1Uw
FoBgXXvY/PiaM1WgQdLXgSTmQa1dCYWaur2qqdCBGbMcB1aDw6zZXjPkIvqs7xVE
bBwNDcB9gQIKn46zfewX2dphVg34m8Lb7Zpe4Wauq0MEOoP6D/7HQzUvXiTCMOO/
Nd5P7flScW7kOkennjWowzhDMIx2iVA6eAKzSRWejz3AmEqRIvUTIUWBSC0BJJG8
T9wNusGcI53HueePnpV57z2MBg/GghpX3vwoqLHh9vdDoEGenuxzc4j1OAqM2aFW
6z9B1mWvbeRf7FRD7vytpAYC0V39bzaP49Bf2Gyn8SI8spYQN8nQkOZInw6dPhfR
F7g2aAdaqABfiT/NVQ/I+XE5q0AL5Ta0OFxr58XJmKbCa6IZbgEfuFUYsRlL5fck
B3vV6v+kyvb2OTZGIKtEQmk7qwdTZendUkUbduXi8dMxNgOtIW8ITXBYMGs1zEn6
hBx3U3+hMgpnngN2eKVafkH7nudN+XlcrSRSQezel/0yv+CgqALE/2ytMdVA9Bsu
HaEm06p0fkYBUURHmZg/VZAB3qg0wH8IyMFz0v41GC+advuykLgebj4fAClfJRdu
8QlW374sI2HZtz8HQvrFDi1TyjEo1y+CkMWb6oXp3SnevK7BPMFXjeMd/zen+lVU
z0gTSdESrvBPtwEHM/wykq/DbZmfYyQK8S56TL0pprRYw3igd2X0AxTMDfVOn/es
Zg36Gm4YRHttGuY3PAqpdqONd2dMGccz3j7sFYyPHmSclBIXt2l7mMJadoDj6WHm
fhrURbXTI4ZtlVwhf77iYiPpfVU+ITIoxksUiRQi8gM4+Qylqge/fk0ykgZgzBnR
NwVcoDeLuwpB9PR0d37+orGQ8ejHoFVNSLydK+u/K9AcbWRNJ4vrAZ4TglXDWHaA
fdol1GKmnX6pdulLQkVHACCn0R3M9ABO0n3KnV/J/GQ+Q1Z87BHQEuo4HCvluf/w
mG5011q/xhsIBDdXvLndwhXhxA6Q6g8SApfLo2S4FHQHfVOhKsSgTZU+L12J21SF
vf5E0PB3wpQkWP3EZF8Z5kj2Np5oS3dfo+7n4csZgKwGcmD9wYkUgewdhLnfjAZh
1Nn/aKUBd1R3s5B4bRQZM8vmdj2h6vqGhB4L5OeY7sV1/35/Kb6u1rO6SQZuVYW6
8pmbx8ZgNzS6UmP0Pltlats+vqGzHY2koilTzvePxdg7QQ4GWERBi3DBN/Zljsi1
`protect END_PROTECTED
