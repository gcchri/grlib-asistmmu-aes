`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kK9MLeRbktDZrswKwCJNJpNTwd9Wlv6V99AToDdH1rqgNFRiBZBG8vptH+0vivVy
azkoN5qSsAGk4TCKSTzpuMOVR2Je2l2HeySrtk0NslOP4VvPuR5I6JMfXjZeIwr5
ARo9RI2NcUi3jPi8tSVfMBTzeLZD7huf2+q6OcoLlT30fmGHUpNd3nvfqqETGj0T
xWEXaYg/ym3pTXeA6C8PtPFpiNTixqnVynJkAWBfNK4MW7KsAr3QHMO9ISXF6Lap
W4viWDyr1sm+MSfAVvqf6YAgDEnNrdOPcYuLPkRpkz3RhqzZGc7iRzeV9AVeWilY
SwjsbVN8R9sUDU8tXGfIpr3SRkZ+KKfX6XCcvDuDFTJKH0xqdYuW+PYCPgKSN2K5
C5H+X3hkWcW6SVe/Y8J+EFH4dMlB9FiYmDYUVp/wkyJpV/AqwdKdr3MGAAsO8hXZ
B2AJrScRX21Fo5n+EHEO/kK7NMf8sO69yduK1WiNpjvbOnHlK+6wg55nPngpbzg2
`protect END_PROTECTED
