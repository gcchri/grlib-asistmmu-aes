`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RGIO0N3YaK25+VVhPpx6TD+UhIvhGm4hQudARbP0pP7MydsEQ1bEi628LxW1a8kT
EjjGBdC38df+nf2TSjOHNDLBIx0DzujxOmyYrgiXYy8hvKBE4nC1iUp4JqpIFTTY
54qW9+Dg5zJjgWKvoZiugyr0MLwIgMUkQXXGc9m/BZPUgVxx759v7BZsdFEe++Xu
X9k4yp1dQG3Op1dbtau06npvN2V25HAxWxVflnLDf0ccjmVm22kvtkVi6yB09lgF
JQUN4+XFKAN6vPWIer+fGYJdeJysjnLKZKu7Kd4U+dPe+vnsLuaXO3RYhQdAEqje
x1RK6PlDmZ0bjVshb4TbwgEJE+Y2Eg7PynfUxl/yNkpBtYrulZ4EsEBGe1POOreO
elk9ocmupemfsub4uHoNNSlkzJeLXUeVnAMR41cjYuPpF44rkqpG6Ifirk/MFiP4
0yadpP8AhtKTd/57I/IDhlVytQAloW/ve+lgRZC+1ssbGNq/vKkC1yWoWd7H0Ko5
sjm3wdic+54d7wOsR646g1oVZmCMMnftmj7CJGgM/wtjkKvgap5b0/CMrGIfSGp0
KJExtvwcWEgy4q/FkDfjYwny5em4lBAg6XkupN8b+Kob5igK8tCjS/R90Mz0aCbG
rZps+RRt93Y+AGxHfdMA3CcZKXWcqj2U7bVFbYbSo7YNg3Yxdp2FB0nxFEqyy14e
idzipNEth6l8qz1KV/SrKpkIY4lJKZvttQbF2YE1KJP/lu7DNPb33p5ajDnE3HVV
kgxR06fjxj9dQ4Ib/zjEmQ==
`protect END_PROTECTED
