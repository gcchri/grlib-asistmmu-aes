`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
afb8K+7krK2elYmsqeb0gLga86kmHolJgGkAnAkwygymiDJX0Y6e5Qw543z/ahez
8d+zU1o8Eq9LCb2vC9TVqL5G/jN2ZiG7Jy7P3dCi928C3UlgQeZrj8CvIB6Q/VPp
hl3mPjHyoDbXwb9bHJ3PETdhfO1+1iPZWmmR/mjoo5nhVfnsyVz6l3R+8VA9MskD
moRZkLjdyKjVWZCrqeMFMstrtuH7d/hEPo5fEIs5E06jKzNftw/sQnI6kg8scrQd
uRmB1DbtMY9w8Rk9MtNKcQ==
`protect END_PROTECTED
