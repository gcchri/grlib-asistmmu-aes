`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XUTuP1OOkUKoTCQw8/xiPwjbWxUhbe1HNM/WI71K8Kv1xioVwYwZQjj8Fpgyg9ye
sYxDG4Y54++aafhyZel2gc7qmcZIEhij0X+d/Vycur50EP4yQ9Xa9CiDEPENY8HR
/kv8FXE0ILN2IprHz/qNBBfItLFnx5cQqvZQKNgFDAqHIJbLBAarVVMfOe+y3ped
idkRc7IejtZPk5rDAgyk2Kh7KCxIkAGzDb0Eu9v7bQbz9B4230a0Op/ZHKOTMq/f
FHOtXKNwfk5tkUhSbHe70Q9xlmFx5xTWOCpZ/8XYsbMDXYBnDQ8hv1dHUFTAkgq8
lDVvKBG88bN32jmBspcQnsluvVmtdHXD/cOLJiWRIvOmJmxZAQqHjkMcw5Sd4cVK
1UquQ0BYUSvfw4N5RVZEwrGcqBtsKG4q+9doRQGXEebbXmFe1idMFmCYRliEOyhH
`protect END_PROTECTED
