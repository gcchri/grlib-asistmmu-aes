`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xgOvZoYqoo6y10VzjmpkLL4c9TBVnQKD60HskyQKDGx6rmckNctXNQVAJyxXewq3
NFQWzEmadY4fVJUl3zV0OAgX0PT6tm5jrrdrXH9B2Md91XPn3k0ftq8vTPhiQ0zn
151dAtx2HgmwauGLe/1FRqnkMo1/F1ncc/JHFE0XpfaUBD289kItqzoQE+qj3mT9
5Rd8QqskLu34i/QPjSbe8Jgng0mMi10WQSozTyybCq15hgH99e3Su2i9iTWeND/K
Azol1xgeuTAsj+u57AYJ7UyG6HdDZhRvKIM4LOnnZkdPycG08LavZtSAEqwUMhpx
mImW+S7XeJO1jUbI+nHMVZlyPKFCXU3tV+Kdz2jJ+Ia1cLyv6b/Go8DHBk6kD83S
EOsV3OozSUENYiqu44V6Juwmap/OUDPv1DEysfzcduRjUhiQdMMIaXcoGRhYXJ2p
RZhtQhsBkKnKI2VuHIZAxvKsKEaZ3J6eSy0y/uiOLKKMbVW8A6Jffrk6f9E9pxK+
d1wXO+mFK4RdbiE+BtGArlcO1jHrj5JP3BqS0SZfVzsUHSeucQxn7VAie/2ixLhV
rpvS0pJNoNl+4lzybWN5TNAaBlxWQjY/dF883rCuY1XbjdbniR9eypTg6EoeAMuz
eTph8hKeVkY2PkuCl2rd2XBiTljlRuy1C0MGStW5rL0=
`protect END_PROTECTED
