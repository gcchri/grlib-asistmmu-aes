`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tdXRJP2Eckyz+Zz0gk4t+9hN2pdIOuACFa0fpQxrBTjLYFMPfMM59klmn2HJoUUd
lhg/2tT5AzGQXOiOTFYX67v7cFjx2dGL6k6DobFxs4wt8rc1zuNX1cCmWX5IEfxG
rNhoJA1kmAd4qqCd9wxrFPhxwxpZc/YrtyckdGyd1x9ZmGQC59CbSTtMGjQYwjPx
ryaGGAlyHgyR5NqCrK+DCy+aLDXYut8gUvao5PZabXX9QZ7ue4rbWpqF8jXbI8q3
Gz2yO9/C6PKQnY9Ka4t+Xg==
`protect END_PROTECTED
