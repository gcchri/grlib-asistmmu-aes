`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AOJj+PBAclQhlungDTYYHuzgdakjgCK0lS+/mRKz0DyVzObJHe3KoyGIAHqKyDJ2
D3FuZPzBQTnPW8H6eZR9+DQEqreXbvUEXp2de6AOrObnOEqXkmCbiwj25sveJVw2
cd5t55aBEDmPnN2jpdAqu6Ze+ssanCzhd7mZINDVnJ0M2f+RSCWgOcaIzoHbg5Fu
/AoZkPURLorcmKAqRz0DyM/hiq6Ve1q5G7RiF+fAGOPC/jtyI9/5kZc8HiYU1xkw
`protect END_PROTECTED
