`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vn8UQwbsRI1wYE/dQsH0/lnZV9eeBrJ+oA3cSQ6fuERiohSvc0qI82O52at8wa+i
qA5Pzoq04zvxU1+xgCEd4qOoGNMFm1u3kkdYlH/rYdS9qebUHIN1nvxrO8HiSw2I
NJCuFq9el7RSzH+wiOCqlOl2uwfmGVagm7vyobeoU4YEbalhfvJBIQ2Cqypie5XF
Cyw3MFmxtSJApFT72uJnXEULSLHvya8vugqk+YmllfGtRdoRcufPhqiSMuj0WUQp
J2dkzEjVYL70t5fBmR/m4eKf5pCvlDiId72XWFKvn/6tM2Vhbg3NQwCWE36nSetP
IYQlGy3Ovq0/24LTd4zRWg/L7G8eyFfCnlUIeU4RJdhpMAj+lH4g+7O6Pt75kD/6
xsLTRuVdKgNhNb+vMUuZSpcdjTiqCBUcGUiuQ90CIW4XF2E9ZWfQttf2I+0MNTVw
aAwE3E25vW+wuLS7ggdUQokj4kS5qES9fYtJCligUCIwhBKdxMlWGxNjxDIIbKM9
Uz4NCXgXCqWR4oPzT/ITUoC25NpivFCNe3jb5EOu2k4pIDb9NyBpsfVPM8uKuEcv
CINRjEGjnvaQbkZ/ycpMo6d/1SRgLwUJwVF32wkQbBDKqda3DKmWzi1v2vcJ/VtL
s1lIk1iWeC0QXzfNIVlrh2lF6/rWmsQMjCKKfWMuZb95pK4kbiesa0odKsQwUn4Y
e7B0IMgABmSXGT4XmxkKbDdqqBAEa5B0IJ80eJQYwV4up6LEUwSaVG6s8IxAQ6YX
mfSMT6PRCMRffHl9I/ePzDV6gyQjPCdFY1KN/N2Df4qQgNqSIVJ7o1C0gmolzU7u
sfJFGeEOXUGZK6zRcjFzK5pzd8gMVqhjuZlSV0JZjn0FUM87LzYbYXSK2tNn5j+s
AXlWuCaoyH7XXwvp399SwgM4GZ5bfPw4bO37XX5JK0eBwkOM/r/tMi2QiMQ2gcws
YXAVzapBOvNJLSheOmG42e4km1PIQB35ful0nJVVMOs=
`protect END_PROTECTED
