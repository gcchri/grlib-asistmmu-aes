`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aZBAO9GpmV8tZz53jpHOxkDbqyJr6TBQAqu/ohDpAyiGU05CPn30TEXQuMKDhCUp
DsKjp1u/6cOnlYrsjpBiOeipR9hgrbNqY+BFxGyDbQkZwpPzWkhJFT2d8Wctr8se
LRAoJsIleEUMGCNPFs5eplGSX+tiS6UXes89MQW+e32BQTEXUP4oexoSn8oz3k4F
+ft0a8R44TovCmwJEsqZGpeWtmr/y5cLzNq8UK3tHDUwJBZedBAqMTUTyZgsHO1a
wKPSIL6xeyDGhHvccJaB258PnvIOsL54uPUbIUeLaNhz8QkhyNwUMwU6pz5va+Qv
um/IWrbd3fImz9ET1Hv4hLJDGaVfwX9Pr1LRcstc0EnuhAw4hMlUfu+sWRJ0XlAv
FNMrVIAxJ/0V+Tyjn61PqniIjlx41LOeX5B8w8PhKHuVsAEFsl1zantYVqumuLFr
RjLpex2xBJS6RayqOk2a6u+155RrRmh9HwOB4oCdWwcshAG9wzdsNQa/ORR41BX/
`protect END_PROTECTED
