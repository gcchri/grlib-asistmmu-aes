`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xJnayXJAPUlAHk/7OokOFfnpXJxJGySvckttcZnS4J5V6lCb66xcmSmOuErUu50n
7zm/kQt8CPYcLqm/Y6nO05kcTKiIQi7fW8ryf5mqhWSMSiOlQUoFV1dQxtOGDre+
SSE/uQ6aS/C/gtubbO/al6Mwr/7O3zWpv+sHzsB4N5/+a4r0RmKQ7XXeR5oaucQO
j6Le+axQJQKemzztUImDBCCM0ZuZu3W85+f5jUcCvKeA1yy+Q1WC2iqWWWj0hsn0
4z7Oie15OYfwiD5A5ESNV1e7NcZsmIheuU6YFpTY7ifimSzKTp2j2sheC+3jHxoC
LbUJIzK9A5dcGIO7XgXeBPPzH5pwI/Y6rz3aGD5McZd0KG6cRWc4OqwqleA9UQYR
RgzAQ1xjlzzuuJp4iMKCeQaOG8SVJdYWgFuAMDQbRtoFTNsgLSsl7yybFQIxFcG5
IhyXTv2tnDi1ppQ13baedz+ED5BWGPeLzN6OUGNOq1rscUyHlvl5X5L5Il+3sBDW
PVvjtHkgyRZHnpfxAQNNLe6SxgLfdgDrpCJjmd6OA4ivRRJnz2C2PUMw2d588UXh
FbayxSBVRiUHiiOGkrUCnAyErEYijY8nJQ9hhaYFC5TiyPMY4GbmqrzBI2RqVaMS
`protect END_PROTECTED
