`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OI1KAot1/ut5H9/ntOfyPTYzck/YU6WC6NjJj61oKmmnsvP3WN0iLYDacAwMFalO
kiT7qPPZizhNzgR5xVzTdrEJIWusb2/0EFCNUh8cYcboEA9T1Ds3g7ezzulAnHXh
r0E4wR7Aft6Y6dlQVMZlshHjCTHrASGEbY8+WOImpzVc8uy4RlYMxMwalFrI72pm
JIFCmC/d1Y5VL/zVnR5KtQY8PUlcTo4KaaZEJI8ap1FsuNyJeEfmUsh9i2F4vnil
CmbI3KoYa79SYFRybzQ1Rdpkp6D/B9p0wZym/itDPhFR5I0cQ+L1o1/K0ckpOeVf
7HxxhFWjcxfu13G32mOoqVHughW3pTx9Q8GB0RGy90zlgheNKiGhlTJFeRMRcNco
asE5pc9U8lStc2Zrja3hcC2Ny4GS3OwMs3O095CSFioamwelbk2Qtj1uCCpNkJEf
1MaI2zw/pahD0UolQw++VISI1Hr1R4Wo+M1wrNR0wsBgJXcRW+0R8Augcz9l3bdG
EkNX2QYRK7AssECSlwcRqMPun2dCrxnP7diQxRIdCmx4nu7sVzGZHFOZqg2KD9ub
1qQTJv8+BBUMNm+0YgeiABi9gMiFrJ9AXp/VC+peugmJzoLHcIflZGsUj2rciZiw
RW0kt6Lh8obesZ0WF6/sOtgOV3R/uxXDY0GdqoWUUwZLEDEZpe37CEIN6yQYswI2
2B1+AMDcfDf/biWzHf1ScscCRQ6THuhDzTlZXWFFB6F578NKK0wZPItyzKl7QSgC
B5jOprtkEM70yTrqRHi4fCxTsXHMRUPAPJDJYgMcXF4SgEV+Y3nRtCnUwoaiNJcl
pTWmW0R/nfDXsSSLYHODqUw3CVhlantG6OXEY+kbyLLYBfOIkdi00smC6mJxhRpZ
qj6+9Xv2u12psMepFHTcbciKVQ+reFgazj2Her0Li8AmoMbDX7YZW1UAnDFQYT3n
7rTzYV9QC8bglUQlQfaS3A==
`protect END_PROTECTED
