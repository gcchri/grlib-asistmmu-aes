`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L7gxJ8JieYCtZxPzac1N2GTVfYsWUCWJjMjQECAtjo14VJ2fehciK1EhLJHYKbUB
m4oVK9NBl0Fj1yF19L4hfn0JWuwxLYQvMVAOMDd0l3Yt4MahJFVmRFV/okNNfpAt
AZY9/0PYVS/lfUVK3tyq8OuFl7nAQnjtD6ONmGmSIKxX8uiA5UVRWTVRWJaVr/L2
cYah8vO5WUKG6sXBSLKNgni6f3ZQCLHiYBpVZEADrsl4sbVo1SR8rLTFyspEPqoQ
xZyYtkvmmo8MLhNkv0eFwAVe/jT99/zEI/0s1hFrnLaXSxH6E6ovWwX5v1EIS0fC
lw4LLxJu93NlDgh2PrWU0QHMIzvAkUxq6DRI2mn48jaUeyU5HQV27z87KUhv6xaM
S79xTCoaLKPW46pB0ScFNUqgwlRo+HliF5TjrYkCAU+7KAoBnLb27fSoexso5uIy
rNJ71vpeY/Sznxy5ikBYamQT/R5Nyg7z1D4dzkJKAW/c9MpMgOIOMUu0MpC+7Mzi
HyHlKXHv1dSZMhKoxCcsXV/rl/na+bfZtFSA/kIRA8tbYoDU3SKoxsufgxyWxSKp
kh8ivMv4TTs/BNZBeWoDW/2IamuYmQGAEaoeKs/wj3qibVnl++Atp5C+12n/nm7P
42fNep8+mc0U8/TVuq2tvpjojgCVC5tEDqg5HjxL68Eg24Z3r8BAed7JXK3cZd5Q
8Doksr4B1lZaTiuasrurQrifU6BzTSRCbU7uoWm+GPDWnuT5ud8sMQW2hveF75nE
t2IXrWh4SwOKKcl+/iE3zQZb6JNWGDn9s03XVjEPLWUjsa8JtOy7aHuUKt3mDwNs
flGPEVHcpTSW/9p79r+N0XRkpANTtLX55+CYXGTOQwMrIYmXoXOpBtweRgmHbi9m
XPsXuGa2aibaqSgpu8/HSY5GDY4X94UWfqP05z7ZwDQZXEuZWMQN/K2ObD20nMrJ
yYSpmkeLp6nKyt3DSF4OgMFWHw2kDm3Lq6iJy+/6TwgPtkhe1ampSBPWZrrun1gG
wgBRk3pVo721rU6wknAil957VdT4VHWbspxkKpRY6MzlYb7APv/PlO+CK1qtuoUF
p65olz92PKbfLkvo3wE8JtKf0NYIt7XL2dBRC1a4dw3hTpAjeVwtCd8jO0YJRkni
`protect END_PROTECTED
