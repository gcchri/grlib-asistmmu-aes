`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9QesjJX4xwmoaqeSBV1giLLihpsrZs5w5/xKb5HZ+GJ6yFq9nPNh3daQtdAm0/Vk
8vzPe/dLfVvCwDv7qe66sXgnG7SoNrlA0g158Dm0e3Ux9XbFZGG/26iZgi4MNUkO
Uru+urhiyx+8xj2v2WCoqB/ml60P/5ZnKPyCcwDHxt6G/RV9d8YFDKlPaherx/97
YAW9/gAFzGyGvIvC5+ytuNjWuq2oCdhDPqu4yzbS+ottWa6s7IXk9fB3aDo/LJsr
yudOdvIL/VWxoPdHQrPvCcW/Dxs3Rg5zSdAiixxB17Zee1Gg+9s7zauH5qB49Jxu
nZD0BbIJvyold1MLCAalugIxJ1erdseryshOOfIgwOC796nm6jgs86EyIIuMAGH1
kjmacVA7fwLyUjEgoB6ysBStrDEoL0uBnZm6Ox753mhEe9VrQCSjhQJoWcpgbdmj
XrCrIJ0jBr2pxTbloMEpKHuHx04iz0ZGKpvuyog51C05amXqTbDk268pSUvA7fw+
Z0SQGpU5ZXnhBU7pveFlJ40mrajTWwd7NaN4E2h38WuyhK/Mq+v0DyyK29YLqs3J
Xr+03MMK5NLdcfMUS4h+c42JSlTw9GvPPd9EizZUa75GxsS/AzyzBpUZbL9EuNTp
BXlDk6tLpJbSybX1hrQmVyyyRWzHv9aTFCqUcmA/9zw=
`protect END_PROTECTED
