`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jB6ZpWucGqU35hObQjxYHiUhqVpUHALP15B1lRU8FCJQEWbzYdPr0cjT2vkuGlGB
fuTsVplRAPXGROQAmo6VPILX+kHQVc+AAZkUVqyXqGXbSGr/8dCbwss+MhodxLe9
nkNDf2dcqYVcY1g6mo+0brU1xr9ZzLAGxdCXqwYyTUj+Ao0dLdoxC1JgEdFeYMsF
tYnjow82q8zgJ3Arh6HpEYhUDPXsdoLAKY2Yfwf3aJFLjdCHdwCK+6xXZaGpwdn6
ZxhoSh5cz3ALwdbjr1iAnx++W3o7xUX3NhVv1rQegz1GPdMoftZPaPkXFhoBmj3u
ANZ8m88H5huUGEVqvDMgK1gkTDkJuBZHHHe/AlkGH6K61cUNDK3NfbuzjGK6bIV5
cgBA+ClphqLq23kspSMLmXwZkS7nIpIzsYRKy+tsUfp1zHBcG22+Jo0nJVlj4q8W
2yQcXjngGtcHcBapNfDDE7G6FQfBZDwNPCPifBfxodcWRaI3bOPRuR/9e2X65GSN
GjH/EDnTrIv4bRhjiKaC0cv9WxcY4FiP386LCgMtiRYG8JrJu6z/y4pToogNfVQv
wKGL5JXK+HIMWt3o0HF6QoyBe0cxD2rlo6iY3cStk/DIoIE91JNGc6Du0DxuRXwD
1DAz31SwOjl9TZzPqCSMTKNz/xTILTvcfBkKaXDEqzZajxg4/y/dBcPwMloIWOM+
2y9iU7FD1P+Dvw+deMnlfxz1cwLA/8UXm0AyxKHidUvEbpBzQJZrsd+pQ5r1VzMo
Qkkz5qClg9q4HkEtBwKdPQ==
`protect END_PROTECTED
