`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9k2kjEZ6hJXztvVbJ8utVJL9R1K8Tug9UkTMLpqbO1OVd1dTnv/NGOEEoD7wJK6q
BbRzsK/BgynVehX4N68WZoFZ3y2RHcZVEijGH1Xgx7QS53ZgasjybmHc5JQqWBZe
wE/wN/spWg6J2BeuJuQqwAi4W96/c7GWYvPdRjIS9lkzJAG6Syg3wejKTt7Dh6Uu
HD1MM8+4C9PO837NmG4HouAoyPBF4L+3JvwG0bYpyjmvkS2S14PtdefpUecXL/Ig
chE+ePBhASQsMDZQZiqKLrngmNMJLG7BwzLJj15JbezfmrCi5TTYqrloUQwH0Uy0
smLauwNAorCUKwI08MaxlQ==
`protect END_PROTECTED
