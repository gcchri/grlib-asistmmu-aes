`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OHYTrnm/B21ebfeMNCvysB/8UUUupPrg7qevy3IyX12VDVjK28k0Tk89FlJPXOsY
qDCM0kkNXujwKIBJ1LOyvnObjO68ATmBe1Odo/EgI6xtdBdqLMTQwcZ7cB7qx4hD
VmGD6eps4GEIBoau22u/Bczro4ZdJUtJ0FGqLTaX8IQM6ulX6ukYpbR1J1WuW6LD
d913snc0ABqpOiucjQBVd+mJd44TfF3eisA3MlE0ESKeSrbnshckraqxJks07hqo
DVAnA4kCO3vlox6t7AC/R3nfBGCUZFu11RJwyhbDJY0/21/N5ToFXIMh486Vtlwm
PDjaQMMdt7lt//mb4wxLiDZR7mfUZ/h5ctjS4l5dhGOT0pGicYkAN1992F+gvETV
t3BVNl92ciAMaZ1ShPCbDWjSnIPlXlbPtExqCySls+MuFdaMSX6p5DvHeDvBRuwn
2PC8V70EKqUlKDoLM5PsQF8t8Jdl72e8DpZh8kCnq+Rgjl1oDxoFvkKYWU/0QnMb
CYMd4iEe3h2P8EWxEHQsx7j/9Y3/xZJZBQQPS+wuBmMAczsVlK82aXLyI+Q+docH
OW3pehUCR+WC8GdZkEt7kyUMfyZTLZsKIwZPNWEzP0A=
`protect END_PROTECTED
