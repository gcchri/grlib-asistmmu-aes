`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dlPZtBKnFTUQg9KBxiO0sRLvOfuP8fQTnRTwWr5tjIuXx1usyQAxSplTBqjiOawd
7OjyHAntM3EoOkXt6kgr+rXT66A7qk5BUzpGVgrH1nkBzBLUbFaAen4QPyaTwC5v
XS8B4oVFoRXgxiS6NJ3Hrtdi4Suie9OpOJpLvNIcl2UX/fwRKxiO4F3xtOHX3h4E
tILg5lsrShHRRVHatoVVm7grYboljKOZFlf+iYRIPqSpJedAK4szLMYNhjrBL07W
25eCEnaji5aFjSWkn5v2nz4Bt/tWdY24VKpwsFvlrTs0b1I7eFUTfCJXIHUWSCbD
yBEcQTNBG/r9faGQbjNbCn9OU0koRPLFWT9qCHFYg08fb8cwq1kNdWrYbrc+CuLD
Nc6imuT4CrLBNAKP5KqW+AKkXguv7mlyUmjBl/NtxIi/L/4RjNAMwkYqkPSkZLSL
5//WFV4I1jCsZbUjQqG0wm7uWQb/wQ59sa8eK9DKKUyBs6HY44SSzwb63m0J9J4G
3uKB9yaEoOwFl4CJfSCcaKGk9Z32FWx4zkc1WENBZ+Z2EuhG38EHRQddgxFC0tML
GoRxUofSM4ys94kLJHT1788NyOsz3/sTrF3ulNgUf8xRA0o0XvEbg9ncCAZVBNnL
GAOnAamH6nIvi3UcGAFEQ5H1aqsZKtWxdwmSLuFStdIs6v720AKlCxg6+nIdX/3v
M11Q6Hrs15e1dE/YDtC0KWbQesF60vujybG/rMhm2wwPgFOmSunJPQ9poXtq9IbG
OnOP9W93HEuijwtfUDDO94L3v4+qBp9isSl0UKLImfQLTURwa1j3IxSs8WTCS7VG
oFppHwKnFZOisIGAQdetU3SmB4IB3OzhMAsp4k2tn1RzSiMsIOkDOnzBY1Mza+6f
lYusAIEGaUmdJ2Acv/meyRv+N4uyz4XvV2aRa5XcTjfl+b4WgVLE20h6FDvWTU6a
VqkGxKVxh9LQvg0aa/x63VuuXm1Q+ygn/hYGSX6iMzm9gURrA4KUhYTRHnhiLhdb
lgvpE+ZG7w6QFH4B+WgI/RJY2OKunk3fjYaLjGnFCm+DyLYtBoNyi7aBEAlCrn4v
caNFP7LEh77NMjGgSY+H/TkAVz72YGrc0O9qzlHagxvAHj3R1+oohQVDGWye081T
NKBj5RJkP+JCHECAa60fpyyz8sWZYojQhqs63Ak20H4k554DWgEMY0xaGh6VBFyc
PWa1GJZEYcq2yhrzWA01TthsFp6TKG57EEnCHeJ3zOWtASmj97y1d11jyXiR2J+G
obQYDZA3DCPqWYZtu8IZKR+raRV8We90tK0uY0nu0LPPW9oWNR0xiMQ7u536zHLY
t49GHHbkGjXK+UeMgd+2eGrHNRNRmwmNHayJLkfeGIEDgfYoyGh/b310rSVLTHE6
2a3I7gXM+l/BrZTF+PeZwwAK0nHU3BOsFrS4d/an4tsPJ4CLjZQxIZUgd9judfUL
p04UZpKP9dlueZRUPZNOHgtmHvBIWjkwTJABtSVigvIAzUf6wdC9V9QcIDcj+mnG
O86YghC5u4tGGpflXqg/RUFd/9QvVZ4eKUMntmgsX5TubzQdmizbaC+jGJ+itM6T
Gm/XDa0hpM0lhWj+BwcU07mOBxT4y3nfc8TK/mpHvwB5nZ8WYXe0xtABkmiP5QHw
vHpTDubqojizmmfev/v15cm3wd3zqj0vq8QOxBUYbSoUTyqTqVzIoWseTIJ3LaG7
PK+Xl+7MNVAA80vngHK0nO4E268s/5v3EkOlrkIZUIvXCLC4iSIDfYwcgWgnoYYN
0cIvwI+s7CysZ6GIiflhQ9GKD+UUv7LXqc/TNPQFufKiveWqm0kGWVJH6/0hVBmn
S9eisOMCqmMmKpRXYlimwtvU1dTulnitcO34z/IMq7RBSxIyaPrDvn/sksES1wRv
4aAVhJNgfRPnC1fLBlgzsdXA+jO1u+Szwg9eO2yyijksvKutJEDlM7D9L4wKR07V
igf8iaYIdHl3x8GGu4q5/ErSLvDv6lalyLP3wCHiD77FT82AqFEIFUNWawm3sKGM
sfMWbBJ53uaCWBbyNSjRDa4OxIgffkztaTxwhpxZpWSZPK7aSzeoi1zhrejyH7I+
JNdlR7PpVSusVE8jrXsiuOxOf9rI0S3JnWyQoDthvpHo6Kx7nSqWuXhDMml76bHH
bpA9FZtdxSFrKaKZ/kFaNKRhTn/LzKP3sL25rVvHVULQwVLMcYxvb/cRfGFZ6ILS
rlVgzr6LSBdkKsQMTnFKkoeOI3/iemw4B/+/S/tHJ/qDU7zOvNJHWawLQzXBwhZT
nCNdzzdh9csCEnsrLSPlVuKF351kGyLH5N3cFu4gI6Dl7RDw6SNB70T3Mmzw+ONf
pqgPCtHnC9Fr6X6dG9CBTnkKTNoVdQQAceNaYgE5L5IgPcFdnrKsa5UsVRxU28Mz
FypOk49xf49Qo8mKiu5Gl3BzLWltVdBvzIJj90RRR4zaZWt7RKBRmJyu9xvmJnBW
fWA+Y5LaLZPySirLFragl9vaIjyKsf7jnL9eiTdZl8W7+sBvgXRkLnKHsXECTVVX
OgapRU4KQGPBaT0qoXr52HZcMsKwqxjBMV3bS/atF4U/u2YHa1vchX98Q78A/IG+
wYonH/pJdetwCXzl6xyUsFlNnC+X/WewOT7+Dw64BDccLgONbMLMZskHJWqj1nny
FSr9tsXbXW7Q/JqvmEJL4sgF9mg5gsSoLNH/VUTZpSqVVlX33oYo8ZFNyIsRu/rV
JMLH5u4GZFVhOe9cFHqEcPvjAjo7QQuXou4gZg7BNTzEUMADEdotr90P8DBmf4s8
AxDrnODIcEy6gJO27/Bku977M5+PocB+Hcb2zBFlWYO3qP3mIjySOjfBFfzVZCqJ
dCcW78v/Ihs7URejiE+Fo2s26Ce0O60xxymodt99ewk=
`protect END_PROTECTED
