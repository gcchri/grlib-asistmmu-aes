`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GlukzGgeEE1blh073XDXr18RAY3ZkexlvIVfj+IjQFcAFv4iIWzR2tNi17gd9R/d
3TDj3r9lUlRASAVpSVy+RfJ8ulQzmUlgH1W665bqJ2nk+L69QEeg4joqw8haIdOM
JmKP83MNs757/AErQdk+NZASzJi13/HDKDecFX+N+Lf5dU2JIBI8RFpmHAP8NzUE
5abOQokvcoALh+3TZ9FojUMhJnNUTLX1pfcLBD0+4TUFrx7HaOstzEatIKU8tSwN
jxuyDuN4c2oZCz7lc7oMbpG7paKUL7UNlhgLB0mtHimH1UMaepK2dPxz2MLqDGSv
glwsXvrP5bpGwVWWAdrZOA==
`protect END_PROTECTED
