`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cg2aKlq7rZRxg5E5C8B613m8CPSlEICrd+vP93UADVPekvznBltfj79NCJRvQZ/o
7Wa+QJTp7YbU080T4xzXkG7sfk+mnjnV8ZgSY6GVl31vGsXbblURb9apvZEPI4Ht
05JhF/pqlMHQHWjvoIMn+2XdLSunzmNMIjLuVA380OY9aMxw/FUrbH+JbehUGea7
xHX8UElSt1Lj30IW8GlLxYLyNNnPomU6beOskaET83673jATvGt6yMk5NGrkipgE
Suh4KhNLxaJM3ir1ukXnDqHI20BS+CLSJNawQIusVi1feCSUm3WxDHORAiIKdN6s
/v57uiuYDGZkjC7ziUB8Ug==
`protect END_PROTECTED
