`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7he0rnA3/fnzhAzHhrT+p4bL1cyUnJY0Pvz4DMAZCJlZm91tzSkIfK6e7mg5/MWN
bVHuqkvEJXG0123iHuLUEOjolKzcuu7DPoETJXj8jR0l6KZ9zFSFiIm94jtkjT34
m5CjQlmKrZiT3zCm8TkBRa+6IEmpEY+z0M8/7hOPcZomZMCogrV1CN1bwdBhhnEj
QlzamWlWheT2/10hcdwZ4ALcH3NIVwmg0RhYOyU3QEKGyE459g1rjTvQvHJr+5zx
N6D4zTc4Wwbd2qsPnldFaCh0pWzZULBG0mbY3ZyYtvhKgUHvGWL2y7dH0TltmHyu
XLY9ReB9SlmI7lZv0M/zAdzCMrgy1ob6Q2l/mzrfHl6YY5G+k5NbcIRI9Xf6EJHk
ZAJYRI9MZQgV4GUUkVWweFvMRw71D2LpDBKJ8K9X7Vpq3E8cKDUEZpIhejuQ54zG
Kl/LcxCjqc8HNqt3HbaYbK8I9qNIUp2OZXX0u09i2PbCeMbhYM3pXeHsHhlQismu
wKE/hb3GNQAs7ATj39gdyhFSpfQeQAAsJVVuSYsM9EC8jn5UFEjC25buay6X0ffq
kxyFfp0mLzqPjJWkqMqjaQxCz3e13t9GGeo1DSggGj3kK42mGyrnZVMSr9PvTeFZ
f+Y3QzpT23SCpmWPotMxPwlBJDDWlarOoXKnO8/KiqQKXIEohPs4W8M1aeVLRFLg
ahgORGKEKaN8wWuY7IG786VbqN5PHgCIUYgkyuoaEbHMsesdXrqbQotgbU0nXLTV
kHTYieYOLcKVDc6iLfVA/Wae1UnESCK7o3wHvMqLoxziHz37ezFFklVrhAjQ0Rou
Kdt/nXaPLLeTiR+cbLYUkRtzuyXaDron2vO7n7epNH8=
`protect END_PROTECTED
