`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wSK7VGz1OewEbKY3FKsRZP+NL1rclZRXXKWl5pDqYV2AbGbvO0h2QWSFMGwEyR3e
UjX/GR52y4HhEimD9XZR/TjHLWnoMxTDp0gXxSw/Y0HETUBOknR3Xq6Pjez6KyEa
ClzgPdhYN5cETFSrsWHAprER1Rta0fNGO7fd8JX4jt3gYv0ETNeTUVrbQnC9uobR
YSbTthklPp6E+rHAXNJMs0WW3dYSxf3GbYH4wlVIT59xuVGtnYr9Fqy83lKiu7kK
Vn0UlNzzdUMyqTWFZht07izFVuEh54/kRAFcEdr3uRYI7IgfMcS1c8aSjSyKxfZW
wzC2QM0OTHj8etSGanD7KU7skFzCVc84umMX7kxrxl7BgZwQG38dxUJytIEJRUnK
WbnOPXC2FCp5jQ4HQwr+gNj0O8zTtlkP0Q4vxl2ZlR/9l3MKFjWO65uZ5WTEEqns
Kcq8RafmyZWVdsB0At5TkcAz6wH7UZ6k9EcNSzUfOQxIs4xPC/ceUnuthdTJLuiV
Qi/5wi2nk50YoKuJKR+YwVxjWquc80iJZ8RyN8O1mnA9SnI4AbRf4KlYWAWhTLrQ
oDq+B8BCCza2mFD3B0pESDQPnpC18vMTPG6pbrxjU9wtNQ+T8EEb+e1T4SbrONR0
WWOFvcnWF+iAD+bk6ZYSnXCUwFQA7ZF6hFcH9yEToP3Pku4SK26uUzrqzFMP2Hyp
v+hOD0sNUZEzZWKXMIZiKnJItu/jSmJHaXQ/UgUiduS4VP3v+Zq/fgNdLOanrQyz
o7FPKef4iQyDKLJU9DCOtbcn+x/W7uIoxN2H9yKgMUpzOM7lnT/N3aA2JHhFKU65
5j2wj7t/NFH8xZHkVAykdel1ApJoXD+XNGHPkUk/o2ttPyz2rgb4bOFDPnIUuCam
juBFsvfwmjBmwfav/mV107a7J20oUei20jmWbHjhLqQ5CP7MN847B2BIFjgrOY9w
08xz5H9e0pOAJXOVrcT5vx6f5xsBvq3aFUOQCl9GNa4bp0er8k24D7ajPB4HTA2B
qFZHPBin3lEDOO5VXKMNW0YVeVqbK9Gn6zsomQ6waf3DVNyFO2q1eN5Oc88FuXNI
w9H3LHMR0bsBwy4OIUKl49+iBfPECuFTj5LclfZmnhSi/+WSE0h5CaDaGK2rClXF
5VGmSvMaX4vTXnow1+UqGS7TdVnvcmEm0CO+Uu46HLbhkPVtsf2j9AvoBg1k3OTO
uq3aeqQIWQzS6ipkUX3VofJFoBcyvb7aunPpsOki1+z3PvgOeXLNjFHm/pI3PZVw
V0cs4cMzdgLLy1e7Z/SlPKgAjKA/xQwBQE+xFsijTJhQj1iYRBntqxv1AcaPqUhU
V3WsNFtiNRPCRr1DjNj5Rx4zUNkJB8o2QWxHS9HWcoPK/Pwfz4oblOz82tOe+Dad
iGD3vO+0mwIxSRhKmhxrCk3hAEEQgQb2SERn7htTlEFEUSBeERkGG33Qphumln0k
y+tQg9HA57YthR9AW+72va6P0iJKdOeYL/5l9PCSlxbUH5MF1BHtbpaHpQ7wYtMr
0z4ENJyTK1RJ1DIh5oqgKzqkrWs8C9fvFeT25O1KqpeleHcNFIGzbamIwTT3DW8o
0iO4hzJ3m/VJXC6heb+WiSOC0kuhl/kN8LVvkVu3dvfy3wvR66O0gTrpPEmCNJpW
HQDmjK1Xxbc9jByJUcDz2TT9W7hVtDiDlgsJOpbNGX4Jy+MHSuD2Aow+rVofzVyF
7ZMhNJAI39Jvt+cwQHzONdxDnErL1DfnO5fT+F8dX0eSyNUrcc/QFrd+7b+tvfRc
FzbGmC+fkzCNL9t12xpxSbLog3nyEoI5T4RtBKrDO68cj3rtDzoLmJHUB+sMayKr
LqRHag3IaEMBLCwML/ZRXfZZPSAWWaHm6DWVksJcFdwm/Ml0ukHJTsBAWOxcpW2y
GqRRJ87LQdSosURwqms+60tlrmZ2qgO31Jz2nvdVBgpGBBgoGlv4YFdckTpjDIQC
PnNUSm+03NRvfvVPBdNH5ogK3IxTvCZ+D/jyf9IVwdX7nYuzCrhOnllO6R7PJr5i
6PcLXwcRsx0QS+y+6V5ilmVQAgVfCzvTgIsAhIlQwGMaRCc7a0zJwH813/PRHxFw
jiNTIdAOlLyC4ufPexBN9GsXvj9eR7YsMEKbAGurFTHwWkve4X8hzpZtx2Wxg+sf
zKMVQ4WbI3JW+qKdSYdD4+S0lHGwSPs/ZmWfx57+i9g=
`protect END_PROTECTED
