`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cUbA9RttrPJ3kL8UUFti4ovz1rsapVYZfCc5IRdoxuIyBhZ/0fZ7/qY1GG3sTuS2
5JzEWkt72noq42cmoVUIaPjMQ+ITaRKsOpKkbGMIeumioomXjzlNV3UAp4R6th0x
E3HdBzXlARRkjgZt2S6d/pCGzbIEDbbIyqhOlTINxH++Vj5bSzukrHP+0fOpOOLo
0l2+ohixr2tImPOe3tXKbSFY3SNhnREoVy/c/+q18AljXdsm5Kl5K68zXmduAcPU
IbPmqEloowfkC309+WgjBUht+3reZIwKHHR8aWr3hbQs14xcmoyiKhsxT/PQFyHx
N218WDdVgplwuc+VSq+iKu/TigF75MK4mM6UwAC1c/HChlxc8HGanAJ1H48jUx9p
mbtgfky+TkHH5ktgZoMEESfr8ngbIH0B4iFL5a3xhImv2DG7JuX5IdWFCGH5lmmC
TM3qRF18kqoSmq+aKS8Bop1usrXOrVYSrlF4J6fGBJc=
`protect END_PROTECTED
