`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lxy0C+S5cHfIZJ3gfZKOMl86ZU4TUfz4S27rQE44796Za9olN93Co4fMGgPQ09Fv
Do9Qi701d8KaH+TW9MtFq26lVgpOBZW10ti1Q6NUragvhnL4tpbkhyTPeTejMya5
cY8htXgBDwIFOgteYzLsintHpY4UWqbp5x8gGYPS0FqK3AqCgIWsD2k89322FZCa
yGohrQ2hWCn5Pv58v0TZSCFCm9MX3KB3oxqrMZ0KXzoVBE3nAfwsUnxypPZ1z/m3
GBl6M+glKmc7oQ3niVLKk1WzNR5vgFEfMTez4V5Tsa2kxbpH6tVdxvNusZFEmpRy
EYOQs4SYMuadn+kEdRxsks8BSJBMCpck4x2vYA5UERUz/FYwMLVhUdIxBFA9pRiP
gNry/DJzCFUv9cpkHGUrEBc0kyx40rhNmtHBu1jSwgHMSC6vXXgw5XIDfM6Ogfn+
WNsJEcHyqkTceiYATsKYAQ==
`protect END_PROTECTED
