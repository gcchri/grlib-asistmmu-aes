`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R+jWtJm5j9pxI5+iFnwQRchs0GWia9xUu/pMAHPoJ8sYVa/HVyy1uxPKGrho9e9c
eWBAGwgzorr/iolY8rlS593Fq9t6LIJMnc7Nql/nI2/IDqPo1ez6BjTtePs/95j1
Y3boc3BZzgrtjZ7LmtDI777Ov/+DyEsKpylm5muPfYSgHWOnfwAhVP7yN8AcCVYD
DUEdQNMQOexvrZpZRItLRZkLWLmJEjbwQWKT9+wb61vFa7xfEazeV2/Q5cr1YHwO
YmDDakAbDaxAZ2Hl1OmdmQ==
`protect END_PROTECTED
