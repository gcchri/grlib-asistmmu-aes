`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RZGUYKeH0JWFp4IcLkJ/b4T1QOHAJ6/Bozbq37a7yg0/jqpETb06oeMiSgLgqXQ9
01QqFA4p6Lkv3WxFERLfB2+ORnPfUXWy4TT8goHwGMyPm6OeA+0/n3vmdNxNi2wi
Ke6EzjZhKfxCXngCDzj8bj32y1b+/0S9O9e9TvJST9mIrxZlPGFhNOSi1KOSRv/8
sryX2Oin2x7saywUzb1ijlh2PrG++neAMlCDMNLnPqnHt/12HNhxjwhI5AC40vGx
G8etyr5wBOBhEhi7aVkJTGsQO6M5M5KMOgIZtd7BaiVayCb+4YlRRbnNw/8bRqp+
aunMH7o72M4DxPigYwWyFXxNIqTeUea0QXslMr0YgmIoGlXMOdHANYcju17Imv7H
8lu5DCFDwpWXjPqegCn9frOn8IaRMv0VO2C3zGVsa7g=
`protect END_PROTECTED
