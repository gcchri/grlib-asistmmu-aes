`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2F9uiluKGWgdGg+0vX4OQWmlNCQ8T88rwkpOefj5IAVpXYoM63q7WYGBIusmkgwj
K+PjxQz/ELT1UXrBW4c1qPK3VEJYgu7rMxko3siLAIRJsyx0cUB5jKB8erNU1SJy
wBnbyXMFmMZxPrRJmnZOL0RR2TjQWNtqYSlsHhWXUPoRSHwWLREgZ2nrDUZ/kCGk
23YWvMHBZY5Z2/evI9w7BIXohx9+zVhyMvRHzP69fRQolcuWCVgFX5HjZogbkjad
u/ln5+IPWIz3ZX+bZ8qGoLVNEXQ9+KLZr47LNtQg7iRqaIRGUeEGlxJ/O5DJobwP
ZxQa+WvFjnMl9ONE4GhsRyAu75fDSkiB6W/4B1f0ZoF6ze5ZKgTlFL7uB551lBY2
nS7tV70DExfgPmMrBf6MhucPGu3kBDkpvKs1zTTbW5WbPifsJywRYqxXCm0ZZ9Am
Y9VkS5NIjJryp+Ocw00Adkn9FdlB3DWGw+SyMO77PwOE0xALpxSeEBjNLFocGM9p
yBR+0XaSa1tliOUg6jqAJk8sMkjedhcKnJvMD8KWwcdkYZBde/U3rE7hAah0CdML
`protect END_PROTECTED
