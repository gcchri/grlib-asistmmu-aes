`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o6dH3mBPOpaL0OhbUlYS/YOWeoBUjFM0XmWFvCes1rvGy3qS2TjYu+DkYBtOC7ol
TjSJa2xMH0HhH9Uqvngd2zSpmA5lN7dYR2JEBK7pugoZno8syNQpMdiELxb1ccoa
aclxnxTAUPtAIt4V7Z2kWQkoUU0EoDwdMDl1plVU2kc0k2TioG545qKmfkDt5pLK
6y/0cqA9U1vPaqxLzNDBN1Mupja0u6b+FSN2Wi5NY9T0ueShrSMebeXC3fYP8kV4
0o+1aGFHN2JUbvmMlaTgXApRl6e8FRrmE6DLcp5bthgV85VpEoqziMW+hyIrKaLv
1CyCgcvyT+b3wDRj8YuTgM5OMEsCoPF3FlK35nJ+Wh0SMHfkPL8weBOctm2YqY8Q
2zqxFfVkOXlvpx5DR47T0lcuOrp500joyXq5N0iLZm/3V/3RV+Nklv9hu81xO8bM
`protect END_PROTECTED
