`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ujob+nE+qoiVNDFFlZW/UJrLr7kE4y/gW6jenmIfyBiaA4E0aFW9SRwjwA5aTTkP
uJXOL2EF9RpC8M8WH65AqyUeVIagXJWwdniLUDWjjY53mnbSpGTO120EJKnwHkIT
qRYAyWoN2fkTwuUoW1AbE8YaJshXjg7pDz4KWrBBmNHvxcQ2ZekFgrwjDIRHK7jA
hu3KLTRnlkqoUKA+mBWe3hbV5k+rDHiLDvRnYzzaONT0TaWJ6p2HZLSBBW/jiBn6
8yxfjDXIxKsoN69i6b75a3IX5IQ8QtkHJ5T7YVlWyWS5ZAbmHuWsMK9OK/I+j7zm
wRKn1HarqUkHjdrsb5Bw6Fsd/kRZL+lsP9QYYy/kPxpjJfNE9WzA/eGeq5TUPN6N
UX2pify+i9ZyLrw7IYxa9G/Nd5L4exQY9FglEkW3OS83bI03WmqYxKHOueen57je
uutxS+AVrQhOoJAu2QTA0bhTJZWJTDuFjByVIPqVbOQMevDCs3I8HSDOm/o8iEqO
`protect END_PROTECTED
