`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Em+rvLCP2qknNIaqu0PZTuKHNpp5Sgd84kaOC5gKBeiQ07aZILx77JuQedoCGGN7
i1+VcwCTlmcScm1YUkknFeWq6kvO9kwebBsiyrpVX7AKsRckRI3VeOPKPvrLhAoz
iaz+cBqmLZCsRWWDJ3H6mzglSmhTQnweHXgzJagIH3k0yS3eEOIiTcME9kPw+sv3
Xn6QtGCk5MK++u8jLYpngDpcV4W47CdeUEC7XJ2wSpjshATp4zCEY+am9FAxjzmP
NGkeDs+uLSyZbtznIBJMKr7B5NNbQQkh8pGWxkU4wNU/FahDraSNu0uJ4lJtxeeX
9JsL9myOw9FvCyS8R+Cc5Q==
`protect END_PROTECTED
