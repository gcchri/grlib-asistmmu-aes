`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tu1agkk6o8ZRtKQQn2ZssaMgFFhK8v8An6D/U0X9HVlPJfHd75/WIGJ6shSK2ExN
Pnd8TBAhDq7/6gXiJFyIiCoKoa4qBrbCBJQHh23uR7AFYZ+AMCBU9FkRrkOcCw0P
vCk/rhid9chZdwJ3yL4GSYJ0NpDcxRjIMJ8cM78OprTtslN3X1nheXr61QA8QWU8
+owniYsmnCefbyXP197yjZvrXOKMrC77ZyH9T62LtgVIQ9sKzHuSigoi6SngEU5B
tmRsej/Bz/dAPneW+pPRvjXsAgrNM+KZE5vLycTx1nT2bmfJgHGRDPAh1zcwvfIv
K1y1ts2eWqQkcs6AV0+M+pYDTTR9zM9MTFvtwlq4hpKUx54zK88cLvwppQMC3wrI
Idh8OfqfT1IpG11i/iztRAQs6onthaPAQwtCikDp2FOK4JwGJC2On6XWaIFilc40
`protect END_PROTECTED
